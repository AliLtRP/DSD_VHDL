// (C) 2001-2013 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License Subscription 
// Agreement, Altera MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


// megafunction wizard: %Arria 10 Transceiver Native PHY v13.1%
// GENERATION: XML
// native_gige_1588.v

// Generated using ACDS version 13.0 0 at 2013.04.23.16:54:25

`timescale 1 ps / 1 ps
module native_gige_1588 (
		input  wire [0:0]   tx_analogreset,            //            tx_analogreset.tx_analogreset
		input  wire [0:0]   tx_digitalreset,           //           tx_digitalreset.tx_digitalreset
		input  wire [0:0]   rx_analogreset,            //            rx_analogreset.rx_analogreset
		input  wire [0:0]   rx_digitalreset,           //           rx_digitalreset.rx_digitalreset
		output wire [0:0]   tx_cal_busy,               //               tx_cal_busy.tx_cal_busy
		output wire [0:0]   rx_cal_busy,               //               rx_cal_busy.rx_cal_busy
		input  wire [0:0]   tx_serial_clk0,            //            tx_serial_clk0.clk
		input  wire [0:0]   tx_serial_clk1,            //            tx_serial_clk1.clk
		input  wire         rx_cdr_refclk0,            //            rx_cdr_refclk0.clk
		input  wire         rx_cdr_refclk1,            //            rx_cdr_refclk1.clk
		output wire [0:0]   tx_serial_data,            //            tx_serial_data.tx_serial_data
		input  wire [0:0]   rx_serial_data,            //            rx_serial_data.rx_serial_data
		input  wire [0:0]   rx_pma_clkslip,            //            rx_pma_clkslip.rx_pma_clkslip
		input  wire [0:0]   rx_seriallpbken,           //           rx_seriallpbken.rx_seriallpbken
		input  wire [0:0]   rx_set_locktodata,         //         rx_set_locktodata.rx_set_locktodata
		input  wire [0:0]   rx_set_locktoref,          //          rx_set_locktoref.rx_set_locktoref
		output wire [0:0]   rx_is_lockedtoref,         //         rx_is_lockedtoref.rx_is_lockedtoref
		output wire [0:0]   rx_is_lockedtodata,        //        rx_is_lockedtodata.rx_is_lockedtodata
		input  wire [0:0]   tx_coreclkin,              //              tx_coreclkin.clk
		input  wire [0:0]   rx_coreclkin,              //              rx_coreclkin.clk
		output wire [0:0]   tx_clkout,                 //                 tx_clkout.clk
		output wire [0:0]   rx_clkout,                 //                 rx_clkout.clk
		output wire [0:0]   tx_pma_clkout,             //             tx_pma_clkout.clk
		output wire [0:0]   tx_pma_div_clkout,         //         tx_pma_div_clkout.clk
		output wire [0:0]   rx_pma_clkout,             //             rx_pma_clkout.clk
		output wire [0:0]   rx_pma_div_clkout,         //         rx_pma_div_clkout.clk
		input  wire [127:0] tx_parallel_data,          //          tx_parallel_data.tx_parallel_data
		input  wire [17:0]  tx_control,                //                tx_control.tx_control
		output wire [127:0] rx_parallel_data,          //          rx_parallel_data.rx_parallel_data
		output wire [19:0]  rx_control,                //                rx_control.rx_control
		input  wire [0:0]   rx_bitslip,                //                rx_bitslip.rx_bitslip
		output wire [0:0]   tx_std_pcfifo_full,        //        tx_std_pcfifo_full.tx_std_pcfifo_full
		output wire [0:0]   tx_std_pcfifo_empty,       //       tx_std_pcfifo_empty.tx_std_pcfifo_empty
		output wire [0:0]   rx_std_pcfifo_full,        //        rx_std_pcfifo_full.rx_std_pcfifo_full
		output wire [0:0]   rx_std_pcfifo_empty,       //       rx_std_pcfifo_empty.rx_std_pcfifo_empty
		input  wire [0:0]   rx_std_bitrev_ena,         //         rx_std_bitrev_ena.rx_std_bitrev_ena
		input  wire [0:0]   tx_polinv,                 //                 tx_polinv.tx_polinv
		input  wire [0:0]   rx_polinv,                 //                 rx_polinv.rx_polinv
		output wire [4:0]   rx_std_bitslipboundarysel, // rx_std_bitslipboundarysel.rx_std_bitslipboundarysel
		input  wire [0:0]   tx_std_elecidle,           //           tx_std_elecidle.tx_std_elecidle
		input  wire [0:0]   tx_enh_data_valid,         //         tx_enh_data_valid.tx_enh_data_valid
		output wire [0:0]   tx_enh_fifo_full,          //          tx_enh_fifo_full.tx_enh_fifo_full
		output wire [3:0]   tx_enh_fifo_cnt,           //           tx_enh_fifo_cnt.tx_enh_fifo_cnt
		output wire [0:0]   rx_enh_data_valid,         //         rx_enh_data_valid.rx_enh_data_valid
		output wire [0:0]   rx_enh_fifo_full,          //          rx_enh_fifo_full.rx_enh_fifo_full
		output wire [0:0]   rx_enh_fifo_del,           //           rx_enh_fifo_del.rx_enh_fifo_del
		output wire [0:0]   rx_enh_fifo_insert,        //        rx_enh_fifo_insert.rx_enh_fifo_insert
		output wire [4:0]   rx_enh_fifo_cnt,           //           rx_enh_fifo_cnt.rx_enh_fifo_cnt
		output wire [0:0]   rx_enh_highber,            //            rx_enh_highber.rx_enh_highber
		input  wire [0:0]   rx_enh_highber_clr_cnt,    //    rx_enh_highber_clr_cnt.rx_enh_highber_clr_cnt
		input  wire [0:0]   rx_enh_clr_errblk_count,   //   rx_enh_clr_errblk_count.rx_enh_clr_errblk_count
		output wire [0:0]   rx_enh_blk_lock,           //           rx_enh_blk_lock.rx_enh_blk_lock
		input  wire [0:0]   reconfig_clk,              //              reconfig_clk.clk
		input  wire [0:0]   reconfig_reset,            //            reconfig_reset.reset
		input  wire [0:0]   reconfig_write,            //             reconfig_avmm.write
		input  wire [0:0]   reconfig_read,             //                          .read
		input  wire [8:0]   reconfig_address,          //                          .address
		input  wire [31:0]  reconfig_writedata,        //                          .writedata
		output wire [31:0]  reconfig_readdata,         //                          .readdata
		output wire [0:0]   reconfig_waitrequest       //                          .waitrequest
	);

	altera_xcvr_native_vi #(
		.duplex_mode                                             ("duplex"),
		.channels                                                (1),
		.data_rate                                               ("1250 Mbps"),
		.bonded_mode                                             ("not_bonded"),
		.pcs_bonding_master                                      (0),
		.enable_hip                                              (0),
		.rcfg_enable                                             (1),
		.rcfg_shared                                             (0),
		.rcfg_jtag_enable                                        (0),
		.hssi_gen3_rx_pcs_block_sync                             ("bypass_block_sync"),
		.hssi_gen3_rx_pcs_block_sync_sm                          ("disable_blk_sync_sm"),
		.hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn                  ("disable"),
		.hssi_gen3_rx_pcs_lpbk_force                             ("lpbk_frce_dis"),
		.hssi_gen3_rx_pcs_mode                                   ("disable_pcs"),
		.hssi_gen3_rx_pcs_rate_match_fifo                        ("bypass_rm_fifo"),
		.hssi_gen3_rx_pcs_rate_match_fifo_latency                ("low_latency"),
		.hssi_gen3_rx_pcs_reverse_lpbk                           ("rev_lpbk_dis"),
		.hssi_gen3_rx_pcs_rx_b4gb_par_lpbk                       ("b4gb_par_lpbk_dis"),
		.hssi_gen3_rx_pcs_rx_force_balign                        ("dis_force_balign"),
		.hssi_gen3_rx_pcs_rx_ins_del_one_skip                    ("ins_del_one_skip_dis"),
		.hssi_gen3_rx_pcs_rx_num_fixed_pat                       (4'b0000),
		.hssi_gen3_rx_pcs_rx_test_out_sel                        ("rx_test_out0"),
		.hssi_gen3_rx_pcs_sup_mode                               ("user_mode"),
		.hssi_gen3_rx_pcs_silicon_rev                            ("es"),
		.hssi_gen3_tx_pcs_mode                                   ("disable_pcs"),
		.hssi_gen3_tx_pcs_reverse_lpbk                           ("rev_lpbk_dis"),
		.hssi_gen3_tx_pcs_sup_mode                               ("user_mode"),
		.hssi_gen3_tx_pcs_tx_bitslip                             (5'b00000),
		.hssi_gen3_tx_pcs_tx_gbox_byp                            ("bypass_gbox"),
		.hssi_gen3_tx_pcs_silicon_rev                            ("es"),
		.hssi_krfec_rx_pcs_blksync_cor_en                        ("detect"),
		.hssi_krfec_rx_pcs_bypass_gb                             ("bypass_dis"),
		.hssi_krfec_rx_pcs_clr_ctrl                              ("both_enabled"),
		.hssi_krfec_rx_pcs_ctrl_bit_reverse                      ("ctrl_bit_reverse_en"),
		.hssi_krfec_rx_pcs_data_bit_reverse                      ("data_bit_reverse_dis"),
		.hssi_krfec_rx_pcs_dv_start                              ("with_blklock"),
		.hssi_krfec_rx_pcs_err_mark_type                         ("err_mark_10g"),
		.hssi_krfec_rx_pcs_error_marking_en                      ("err_mark_dis"),
		.hssi_krfec_rx_pcs_fast_search_en                        ("fast"),
		.hssi_krfec_rx_pcs_lpbk_mode                             ("lpbk_dis"),
		.hssi_krfec_rx_pcs_silicon_rev                           ("es"),
		.hssi_krfec_rx_pcs_parity_invalid_enum                   (8'b00001000),
		.hssi_krfec_rx_pcs_parity_valid_num                      (4'b0100),
		.hssi_krfec_rx_pcs_prot_mode                             ("disable_mode"),
		.hssi_krfec_rx_pcs_receive_order                         ("receive_lsb"),
		.hssi_krfec_rx_pcs_rx_testbus_sel                        ("overall"),
		.hssi_krfec_rx_pcs_signal_ok_en                          ("sig_ok_en"),
		.hssi_krfec_rx_pcs_sup_mode                              ("user_mode"),
		.hssi_krfec_tx_pcs_burst_err                             ("burst_err_dis"),
		.hssi_krfec_tx_pcs_burst_err_len                         ("burst_err_len1"),
		.hssi_krfec_tx_pcs_ctrl_bit_reverse                      ("ctrl_bit_reverse_en"),
		.hssi_krfec_tx_pcs_data_bit_reverse                      ("data_bit_reverse_dis"),
		.hssi_krfec_tx_pcs_enc_frame_query                       ("enc_query_dis"),
		.hssi_krfec_tx_pcs_silicon_rev                           ("es"),
		.hssi_krfec_tx_pcs_prot_mode                             ("disable_mode"),
		.hssi_krfec_tx_pcs_sup_mode                              ("user_mode"),
		.hssi_krfec_tx_pcs_transcode_err                         ("trans_err_dis"),
		.hssi_krfec_tx_pcs_transmit_order                        ("transmit_lsb"),
		.hssi_krfec_tx_pcs_tx_testbus_sel                        ("overall"),
		.hssi_10g_rx_pcs_align_del                               ("align_del_dis"),
		.hssi_10g_rx_pcs_ber_bit_err_total_cnt                   ("bit_err_total_cnt_10g"),
		.hssi_10g_rx_pcs_ber_clken                               ("ber_clk_en"),
		.hssi_10g_rx_pcs_ber_xus_timer_window                    (21'b000000100110001001010),
		.hssi_10g_rx_pcs_bitslip_mode                            ("bitslip_dis"),
		.hssi_10g_rx_pcs_blksync_bitslip_type                    ("bitslip_comb"),
		.hssi_10g_rx_pcs_blksync_bitslip_wait_cnt                (3'b001),
		.hssi_10g_rx_pcs_blksync_bitslip_wait_type               ("bitslip_cnt"),
		.hssi_10g_rx_pcs_blksync_bypass                          ("blksync_bypass_dis"),
		.hssi_10g_rx_pcs_blksync_clken                           ("blksync_clk_en"),
		.hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt             ("enum_invalid_sh_cnt_10g"),
		.hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock            ("knum_sh_cnt_postlock_10g"),
		.hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock             ("knum_sh_cnt_prelock_10g"),
		.hssi_10g_rx_pcs_blksync_pipeln                          ("blksync_pipeln_dis"),
		.hssi_10g_rx_pcs_control_del                             ("control_del_none"),
		.hssi_10g_rx_pcs_crcchk_bypass                           ("crcchk_bypass_en"),
		.hssi_10g_rx_pcs_crcchk_clken                            ("crcchk_clk_dis"),
		.hssi_10g_rx_pcs_crcchk_inv                              ("crcchk_inv_en"),
		.hssi_10g_rx_pcs_crcchk_pipeln                           ("crcchk_pipeln_en"),
		.hssi_10g_rx_pcs_crcflag_pipeln                          ("crcflag_pipeln_en"),
		.hssi_10g_rx_pcs_ctrl_bit_reverse                        ("ctrl_bit_reverse_en"),
		.hssi_10g_rx_pcs_data_bit_reverse                        ("data_bit_reverse_dis"),
		.hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass                  ("dec_64b66b_rxsm_bypass_dis"),
		.hssi_10g_rx_pcs_dec64b66b_clken                         ("dec64b66b_clk_en"),
		.hssi_10g_rx_pcs_descrm_bypass                           ("descrm_bypass_dis"),
		.hssi_10g_rx_pcs_descrm_clken                            ("descrm_clk_en"),
		.hssi_10g_rx_pcs_descrm_mode                             ("async"),
		.hssi_10g_rx_pcs_descrm_pipeln                           ("enable"),
		.hssi_10g_rx_pcs_dis_signal_ok                           ("dis_signal_ok_dis"),
		.hssi_10g_rx_pcs_dispchk_bypass                          ("dispchk_bypass_en"),
		.hssi_10g_rx_pcs_empty_flag_type                         ("empty_rd_side"),
		.hssi_10g_rx_pcs_fast_path                               ("fast_path_dis"),
		.hssi_10g_rx_pcs_fec_clken                               ("fec_clk_dis"),
		.hssi_10g_rx_pcs_fec_enable                              ("fec_dis"),
		.hssi_10g_rx_pcs_fifo_double_read                        ("fifo_double_read_dis"),
		.hssi_10g_rx_pcs_fifo_stop_rd                            ("n_rd_empty"),
		.hssi_10g_rx_pcs_fifo_stop_wr                            ("n_wr_full"),
		.hssi_10g_rx_pcs_force_align                             ("force_align_dis"),
		.hssi_10g_rx_pcs_framesync_skip_none                     ("disable"),
		.hssi_10g_rx_pcs_frmsync_bypass                          ("frmsync_bypass_en"),
		.hssi_10g_rx_pcs_frmsync_clken                           ("frmsync_clk_dis"),
		.hssi_10g_rx_pcs_frmsync_enum_scrm                       ("enum_scrm_default"),
		.hssi_10g_rx_pcs_frmsync_enum_sync                       ("enum_sync_default"),
		.hssi_10g_rx_pcs_frmsync_flag_type                       ("location_only"),
		.hssi_10g_rx_pcs_frmsync_knum_sync                       ("knum_sync_default"),
		.hssi_10g_rx_pcs_frmsync_mfrm_length                     (16'b0000100000000000),
		.hssi_10g_rx_pcs_frmsync_pipeln                          ("frmsync_pipeln_en"),
		.hssi_10g_rx_pcs_full_flag_type                          ("full_wr_side"),
		.hssi_10g_rx_pcs_gb_rx_idwidth                           ("width_40"),
		.hssi_10g_rx_pcs_gb_rx_odwidth                           ("width_66"),
		.hssi_10g_rx_pcs_gbexp_clken                             ("gbexp_clk_en"),
		.hssi_10g_rx_pcs_low_latency_en                          ("disable"),
		.hssi_10g_rx_pcs_lpbk_mode                               ("lpbk_dis"),
		.hssi_10g_rx_pcs_master_clk_sel                          ("master_rx_pma_clk"),
		.hssi_10g_rx_pcs_silicon_rev                             ("es"),
		.hssi_10g_rx_pcs_pempty_flag_type                        ("pempty_rd_side"),
		.hssi_10g_rx_pcs_pfull_flag_type                         ("pfull_wr_side"),
		.hssi_10g_rx_pcs_phcomp_rd_del                           ("phcomp_rd_del2"),
		.hssi_10g_rx_pcs_pld_if_type                             ("reg"),
		.hssi_10g_rx_pcs_prot_mode                               ("teng_1588_mode"),
		.hssi_10g_rx_pcs_rand_clken                              ("rand_clk_en"),
		.hssi_10g_rx_pcs_rd_clk_sel                              ("rd_rx_pma_clk"),
		.hssi_10g_rx_pcs_rdfifo_clken                            ("rdfifo_clk_en"),
		.hssi_10g_rx_pcs_rx_fifo_write_ctrl                      ("blklock_stops"),
		.hssi_10g_rx_pcs_rx_scrm_width                           ("bit64"),
		.hssi_10g_rx_pcs_rx_sh_location                          ("lsb"),
		.hssi_10g_rx_pcs_rx_signal_ok_sel                        ("synchronized_ver"),
		.hssi_10g_rx_pcs_rx_sm_bypass                            ("rx_sm_bypass_dis"),
		.hssi_10g_rx_pcs_rx_sm_hiber                             ("rx_sm_hiber_en"),
		.hssi_10g_rx_pcs_rx_sm_pipeln                            ("rx_sm_pipeln_en"),
		.hssi_10g_rx_pcs_rx_testbus_sel                          ("blank_testbus"),
		.hssi_10g_rx_pcs_rx_true_b2b                             ("b2b"),
		.hssi_10g_rx_pcs_rxfifo_empty                            ("empty_default"),
		.hssi_10g_rx_pcs_rxfifo_full                             ("full_default"),
		.hssi_10g_rx_pcs_rxfifo_mode                             ("register_mode"),
		.hssi_10g_rx_pcs_rxfifo_pempty                           ("pempty2"),
		.hssi_10g_rx_pcs_rxfifo_pfull                            ("pfull23"),
		.hssi_10g_rx_pcs_stretch_num_stages                      ("one_stage"),
		.hssi_10g_rx_pcs_sup_mode                                ("user_mode"),
		.hssi_10g_rx_pcs_test_mode                               ("test_off"),
		.hssi_10g_rx_pcs_wrfifo_clken                            ("wrfifo_clk_en"),
		.hssi_10g_tx_pcs_bitslip_en                              ("bitslip_dis"),
		.hssi_10g_tx_pcs_bonding_dft_en                          ("dft_dis"),
		.hssi_10g_tx_pcs_bonding_dft_val                         ("dft_0"),
		.hssi_10g_tx_pcs_crcgen_bypass                           ("crcgen_bypass_en"),
		.hssi_10g_tx_pcs_crcgen_clken                            ("crcgen_clk_dis"),
		.hssi_10g_tx_pcs_crcgen_err                              ("crcgen_err_dis"),
		.hssi_10g_tx_pcs_crcgen_inv                              ("crcgen_inv_en"),
		.hssi_10g_tx_pcs_ctrl_bit_reverse                        ("ctrl_bit_reverse_en"),
		.hssi_10g_tx_pcs_data_bit_reverse                        ("data_bit_reverse_dis"),
		.hssi_10g_tx_pcs_dispgen_bypass                          ("dispgen_bypass_en"),
		.hssi_10g_tx_pcs_dispgen_clken                           ("dispgen_clk_dis"),
		.hssi_10g_tx_pcs_dispgen_err                             ("dispgen_err_dis"),
		.hssi_10g_tx_pcs_dispgen_pipeln                          ("dispgen_pipeln_dis"),
		.hssi_10g_tx_pcs_distdwn_bypass_pipeln                   ("distdwn_bypass_pipeln_dis"),
		.hssi_10g_tx_pcs_distdwn_master                          ("distdwn_master_en"),
		.hssi_10g_tx_pcs_distup_bypass_pipeln                    ("distup_bypass_pipeln_dis"),
		.hssi_10g_tx_pcs_distup_master                           ("distup_master_en"),
		.hssi_10g_tx_pcs_dv_bond                                 ("dv_bond_dis"),
		.hssi_10g_tx_pcs_empty_flag_type                         ("empty_rd_side"),
		.hssi_10g_tx_pcs_enc_64b66b_txsm_bypass                  ("enc_64b66b_txsm_bypass_dis"),
		.hssi_10g_tx_pcs_enc64b66b_txsm_clken                    ("enc64b66b_txsm_clk_en"),
		.hssi_10g_tx_pcs_fastpath                                ("fastpath_dis"),
		.hssi_10g_tx_pcs_fec_clken                               ("fec_clk_dis"),
		.hssi_10g_tx_pcs_fec_enable                              ("fec_dis"),
		.hssi_10g_tx_pcs_fifo_double_write                       ("fifo_double_write_dis"),
		.hssi_10g_tx_pcs_fifo_reg_fast                           ("fifo_reg_fast_dis"),
		.hssi_10g_tx_pcs_fifo_stop_rd                            ("n_rd_empty"),
		.hssi_10g_tx_pcs_fifo_stop_wr                            ("n_wr_full"),
		.hssi_10g_tx_pcs_framegen_skip_none                      ("disable"),
		.hssi_10g_tx_pcs_frmgen_burst                            ("frmgen_burst_dis"),
		.hssi_10g_tx_pcs_frmgen_bypass                           ("frmgen_bypass_en"),
		.hssi_10g_tx_pcs_frmgen_clken                            ("frmgen_clk_dis"),
		.hssi_10g_tx_pcs_frmgen_mfrm_length                      (16'b0000100000000000),
		.hssi_10g_tx_pcs_frmgen_pipeln                           ("frmgen_pipeln_en"),
		.hssi_10g_tx_pcs_frmgen_pyld_ins                         ("frmgen_pyld_ins_dis"),
		.hssi_10g_tx_pcs_frmgen_wordslip                         ("frmgen_wordslip_dis"),
		.hssi_10g_tx_pcs_full_flag_type                          ("full_wr_side"),
		.hssi_10g_tx_pcs_gb_pipeln_bypass                        ("disable"),
		.hssi_10g_tx_pcs_gb_tx_idwidth                           ("width_66"),
		.hssi_10g_tx_pcs_gb_tx_odwidth                           ("width_40"),
		.hssi_10g_tx_pcs_gbred_clken                             ("gbred_clk_en"),
		.hssi_10g_tx_pcs_indv                                    ("indv_en"),
		.hssi_10g_tx_pcs_low_latency_en                          ("disable"),
		.hssi_10g_tx_pcs_master_clk_sel                          ("master_tx_pma_clk"),
		.hssi_10g_tx_pcs_silicon_rev                             ("es"),
		.hssi_10g_tx_pcs_pempty_flag_type                        ("pempty_rd_side"),
		.hssi_10g_tx_pcs_pfull_flag_type                         ("pfull_wr_side"),
		.hssi_10g_tx_pcs_phcomp_rd_del                           ("phcomp_rd_del2"),
		.hssi_10g_tx_pcs_pld_if_type                             ("reg"),
		.hssi_10g_tx_pcs_prot_mode                               ("teng_1588_mode"),
		.hssi_10g_tx_pcs_pseudo_random                           ("all_0"),
		.hssi_10g_tx_pcs_pseudo_seed_a                           (58'b1111111111111111111111111111111111111111111111111111111111),
		.hssi_10g_tx_pcs_pseudo_seed_b                           (58'b1111111111111111111111111111111111111111111111111111111111),
		.hssi_10g_tx_pcs_random_disp                             ("disable"),
		.hssi_10g_tx_pcs_rdfifo_clken                            ("rdfifo_clk_en"),
		.hssi_10g_tx_pcs_scrm_bypass                             ("scrm_bypass_dis"),
		.hssi_10g_tx_pcs_scrm_clken                              ("scrm_clk_en"),
		.hssi_10g_tx_pcs_scrm_mode                               ("async"),
		.hssi_10g_tx_pcs_scrm_pipeln                             ("enable"),
		.hssi_10g_tx_pcs_sh_err                                  ("sh_err_dis"),
		.hssi_10g_tx_pcs_sop_mark                                ("sop_mark_dis"),
		.hssi_10g_tx_pcs_stretch_num_stages                      ("one_stage"),
		.hssi_10g_tx_pcs_sup_mode                                ("user_mode"),
		.hssi_10g_tx_pcs_test_mode                               ("test_off"),
		.hssi_10g_tx_pcs_tx_scrm_err                             ("scrm_err_dis"),
		.hssi_10g_tx_pcs_tx_scrm_width                           ("bit64"),
		.hssi_10g_tx_pcs_tx_sh_location                          ("lsb"),
		.hssi_10g_tx_pcs_tx_sm_bypass                            ("tx_sm_bypass_dis"),
		.hssi_10g_tx_pcs_tx_sm_pipeln                            ("tx_sm_pipeln_en"),
		.hssi_10g_tx_pcs_tx_testbus_sel                          ("blank_testbus"),
		.hssi_10g_tx_pcs_txfifo_empty                            ("empty_default"),
		.hssi_10g_tx_pcs_txfifo_full                             ("full_default"),
		.hssi_10g_tx_pcs_txfifo_mode                             ("register_mode"),
		.hssi_10g_tx_pcs_txfifo_pempty                           ("pempty2"),
		.hssi_10g_tx_pcs_txfifo_pfull                            ("pfull13"),
		.hssi_10g_tx_pcs_wr_clk_sel                              ("wr_tx_pma_clk"),
		.hssi_10g_tx_pcs_wrfifo_clken                            ("wrfifo_clk_en"),
		.hssi_8g_rx_pcs_auto_error_replacement                   ("dis_err_replace"),
		.hssi_8g_rx_pcs_auto_speed_nego                          ("dis_asn"),
		.hssi_8g_rx_pcs_bit_reversal                             ("dis_bit_reversal"),
		.hssi_8g_rx_pcs_bonding_dft_en                           ("dft_dis"),
		.hssi_8g_rx_pcs_bonding_dft_val                          ("dft_0"),
		.hssi_8g_rx_pcs_bypass_pipeline_reg                      ("dis_bypass_pipeline"),
		.hssi_8g_rx_pcs_byte_deserializer                        ("dis_bds"),
		.hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask                    ("dis_rxvalid_mask"),
		.hssi_8g_rx_pcs_clkcmp_pattern_n                         (20'b00000000000000000000),
		.hssi_8g_rx_pcs_clkcmp_pattern_p                         (20'b00000000000000000000),
		.hssi_8g_rx_pcs_clock_gate_bds_dec_asn                   ("dis_bds_dec_asn_clk_gating"),
		.hssi_8g_rx_pcs_clock_gate_cdr_eidle                     ("en_cdr_eidle_clk_gating"),
		.hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk                   ("en_dw_pc_wrclk_gating"),
		.hssi_8g_rx_pcs_clock_gate_dw_rm_rd                      ("en_dw_rm_rdclk_gating"),
		.hssi_8g_rx_pcs_clock_gate_dw_rm_wr                      ("en_dw_rm_wrclk_gating"),
		.hssi_8g_rx_pcs_clock_gate_dw_wa                         ("en_dw_wa_clk_gating"),
		.hssi_8g_rx_pcs_clock_gate_pc_rdclk                      ("dis_pc_rdclk_gating"),
		.hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk                   ("dis_sw_pc_wrclk_gating"),
		.hssi_8g_rx_pcs_clock_gate_sw_rm_rd                      ("en_sw_rm_rdclk_gating"),
		.hssi_8g_rx_pcs_clock_gate_sw_rm_wr                      ("en_sw_rm_wrclk_gating"),
		.hssi_8g_rx_pcs_clock_gate_sw_wa                         ("dis_sw_wa_clk_gating"),
		.hssi_8g_rx_pcs_eidle_entry_eios                         ("dis_eidle_eios"),
		.hssi_8g_rx_pcs_eidle_entry_iei                          ("dis_eidle_iei"),
		.hssi_8g_rx_pcs_eidle_entry_sd                           ("dis_eidle_sd"),
		.hssi_8g_rx_pcs_eightb_tenb_decoder                      ("en_8b10b_ibm"),
		.hssi_8g_rx_pcs_err_flags_sel                            ("err_flags_wa"),
		.hssi_8g_rx_pcs_fixed_pat_det                            ("dis_fixed_patdet"),
		.hssi_8g_rx_pcs_fixed_pat_num                            (4'b0000),
		.hssi_8g_rx_pcs_force_signal_detect                      ("en_force_signal_detect"),
		.hssi_8g_rx_pcs_gen3_clk_en                              ("disable_clk"),
		.hssi_8g_rx_pcs_gen3_rx_clk_sel                          ("rcvd_clk"),
		.hssi_8g_rx_pcs_gen3_tx_clk_sel                          ("tx_pma_clk"),
		.hssi_8g_rx_pcs_hip_mode                                 ("dis_hip"),
		.hssi_8g_rx_pcs_ibm_invalid_code                         ("dis_ibm_invalid_code"),
		.hssi_8g_rx_pcs_invalid_code_flag_only                   ("dis_invalid_code_only"),
		.hssi_8g_rx_pcs_pad_or_edb_error_replace                 ("replace_edb"),
		.hssi_8g_rx_pcs_pcs_bypass                               ("dis_pcs_bypass"),
		.hssi_8g_rx_pcs_phase_comp_rdptr                         ("enable_rdptr"),
		.hssi_8g_rx_pcs_phase_compensation_fifo                  ("register_fifo"),
		.hssi_8g_rx_pcs_pipe_if_enable                           ("dis_pipe_rx"),
		.hssi_8g_rx_pcs_pma_dw                                   ("ten_bit"),
		.hssi_8g_rx_pcs_polinv_8b10b_dec                         ("dis_polinv_8b10b_dec"),
		.hssi_8g_rx_pcs_prot_mode                                ("gige_1588"),
		.hssi_8g_rx_pcs_rate_match                               ("dis_rm"),
		.hssi_8g_rx_pcs_rate_match_del_thres                     ("dis_rm_del_thres"),
		.hssi_8g_rx_pcs_rate_match_empty_thres                   ("dis_rm_empty_thres"),
		.hssi_8g_rx_pcs_rate_match_full_thres                    ("dis_rm_full_thres"),
		.hssi_8g_rx_pcs_rate_match_ins_thres                     ("dis_rm_ins_thres"),
		.hssi_8g_rx_pcs_rate_match_start_thres                   ("dis_rm_start_thres"),
		.hssi_8g_rx_pcs_rx_clk_free_running                      ("en_rx_clk_free_run"),
		.hssi_8g_rx_pcs_rx_clk2                                  ("rcvd_clk_clk2"),
		.hssi_8g_rx_pcs_rx_pcs_urst                              ("en_rx_pcs_urst"),
		.hssi_8g_rx_pcs_rx_rcvd_clk                              ("rcvd_clk_rcvd_clk"),
		.hssi_8g_rx_pcs_rx_rd_clk                                ("rx_clk"),
		.hssi_8g_rx_pcs_rx_refclk                                ("dis_refclk_sel"),
		.hssi_8g_rx_pcs_rx_wr_clk                                ("rx_clk2_div_1_2_4"),
		.hssi_8g_rx_pcs_sup_mode                                 ("user_mode"),
		.hssi_8g_rx_pcs_symbol_swap                              ("dis_symbol_swap"),
		.hssi_8g_rx_pcs_sync_sm_idle_eios                        ("dis_syncsm_idle"),
		.hssi_8g_rx_pcs_test_bus_sel                             ("tx_testbus"),
		.hssi_8g_rx_pcs_tx_rx_parallel_loopback                  ("dis_plpbk"),
		.hssi_8g_rx_pcs_wa_boundary_lock_ctrl                    ("sync_sm"),
		.hssi_8g_rx_pcs_wa_clk_slip_spacing                      (10'b0000010000),
		.hssi_8g_rx_pcs_wa_det_latency_sync_status_beh           ("dont_care_assert_sync"),
		.hssi_8g_rx_pcs_wa_disp_err_flag                         ("en_disp_err_flag"),
		.hssi_8g_rx_pcs_wa_kchar                                 ("dis_kchar"),
		.hssi_8g_rx_pcs_wa_pd                                    ("wa_pd_10"),
		.hssi_8g_rx_pcs_wa_pd_data                               (40'b0000000000000000000000000000000101111100),
		.hssi_8g_rx_pcs_wa_pd_polarity                           ("dont_care_both_pol"),
		.hssi_8g_rx_pcs_wa_pld_controlled                        ("dis_pld_ctrl"),
		.hssi_8g_rx_pcs_wa_renumber_data                         (6'b000011),
		.hssi_8g_rx_pcs_wa_rgnumber_data                         (8'b00000011),
		.hssi_8g_rx_pcs_wa_rknumber_data                         (8'b00000011),
		.hssi_8g_rx_pcs_wa_rosnumber_data                        (2'b01),
		.hssi_8g_rx_pcs_wa_rvnumber_data                         (13'b0000000000000),
		.hssi_8g_rx_pcs_wa_sync_sm_ctrl                          ("gige_sync_sm"),
		.hssi_8g_rx_pcs_wait_cnt                                 (12'b000000000000),
		.hssi_8g_rx_pcs_silicon_rev                              ("es"),
		.hssi_8g_tx_pcs_auto_speed_nego_gen2                     ("dis_asn_g2"),
		.hssi_8g_tx_pcs_bit_reversal                             ("dis_bit_reversal"),
		.hssi_8g_tx_pcs_bonding_dft_en                           ("dft_dis"),
		.hssi_8g_tx_pcs_bonding_dft_val                          ("dft_0"),
		.hssi_8g_tx_pcs_bypass_pipeline_reg                      ("dis_bypass_pipeline"),
		.hssi_8g_tx_pcs_byte_serializer                          ("dis_bs"),
		.hssi_8g_tx_pcs_clock_gate_bs_enc                        ("dis_bs_enc_clk_gating"),
		.hssi_8g_tx_pcs_clock_gate_dw_fifowr                     ("en_dw_fifowr_clk_gating"),
		.hssi_8g_tx_pcs_clock_gate_fiford                        ("dis_fiford_clk_gating"),
		.hssi_8g_tx_pcs_clock_gate_sw_fifowr                     ("dis_sw_fifowr_clk_gating"),
		.hssi_8g_tx_pcs_data_selection_8b10b_encoder_input       ("gige_idle_conversion"),
		.hssi_8g_tx_pcs_dynamic_clk_switch                       ("dis_dyn_clk_switch"),
		.hssi_8g_tx_pcs_eightb_tenb_disp_ctrl                    ("dis_disp_ctrl"),
		.hssi_8g_tx_pcs_eightb_tenb_encoder                      ("en_8b10b_ibm"),
		.hssi_8g_tx_pcs_force_echar                              ("dis_force_echar"),
		.hssi_8g_tx_pcs_force_kchar                              ("dis_force_kchar"),
		.hssi_8g_tx_pcs_gen3_dynclk_by16                         ("disable_gen3_by16"),
		.hssi_8g_tx_pcs_gen3_tx_clk_sel                          ("dis_tx_clk"),
		.hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel                     ("dis_tx_pipe_clk"),
		.hssi_8g_tx_pcs_hip_mode                                 ("dis_hip"),
		.hssi_8g_tx_pcs_pcs_bypass                               ("dis_pcs_bypass"),
		.hssi_8g_tx_pcs_phase_comp_rdptr                         ("enable_rdptr"),
		.hssi_8g_tx_pcs_phase_compensation_fifo                  ("register_fifo"),
		.hssi_8g_tx_pcs_phfifo_write_clk_sel                     ("tx_clk"),
		.hssi_8g_tx_pcs_pma_dw                                   ("ten_bit"),
		.hssi_8g_tx_pcs_prot_mode                                ("gige_1588"),
		.hssi_8g_tx_pcs_refclk_b_clk_sel                         ("tx_pma_clock"),
		.hssi_8g_tx_pcs_revloop_back_rm                          ("dis_rev_loopback_rx_rm"),
		.hssi_8g_tx_pcs_sup_mode                                 ("user_mode"),
		.hssi_8g_tx_pcs_symbol_swap                              ("dis_symbol_swap"),
		.hssi_8g_tx_pcs_tx_bitslip                               ("dis_tx_bitslip"),
		.hssi_8g_tx_pcs_tx_compliance_controlled_disparity       ("dis_txcompliance"),
		.hssi_8g_tx_pcs_tx_fast_pld_reg                          ("dis_tx_fast_pld_reg"),
		.hssi_8g_tx_pcs_txclk_freerun                            ("en_freerun_tx"),
		.hssi_8g_tx_pcs_txpcs_urst                               ("en_txpcs_urst"),
		.hssi_8g_tx_pcs_silicon_rev                              ("es"),
		.hssi_tx_pld_pcs_interface_silicon_rev                   ("es"),
		.hssi_tx_pld_pcs_interface_pcs_tx_clk_source             ("eightg"),
		.hssi_tx_pld_pcs_interface_pcs_tx_data_source            ("hip_disable"),
		.hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en          ("delay1_clk_disable"),
		.hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel         ("pcs_tx_clk"),
		.hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl            ("delay1_path0"),
		.hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel        ("no_delay"),
		.hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en          ("delay2_clk_disable"),
		.hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl            ("delay2_path0"),
		.hssi_tx_pld_pcs_interface_pcs_tx_output_sel             ("teng_output"),
		.hssi_rx_pld_pcs_interface_silicon_rev                   ("es"),
		.hssi_rx_pld_pcs_interface_pcs_rx_block_sel              ("eightg"),
		.hssi_rx_pld_pcs_interface_pcs_rx_clk_sel                ("pld_rx_clk"),
		.hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en             ("hip_rx_disable"),
		.hssi_rx_pld_pcs_interface_pcs_rx_output_sel             ("teng_output"),
		.hssi_rx_pld_pcs_interface_pcs_rx_pld_clk_en             ("pcs_pld_rx_enable"),
		.hssi_common_pld_pcs_interface_hrdrstctrl_en             ("hrst_dis"),
		.hssi_common_pld_pcs_interface_silicon_rev               ("es"),
		.hssi_common_pld_pcs_interface_pcs_testbus_block_sel     ("eightg"),
		.hssi_rx_pcs_pma_interface_block_sel                     ("eight_g_pcs"),
		.hssi_rx_pcs_pma_interface_channel_operation_mode        ("tx_rx_pair_enabled"),
		.hssi_rx_pcs_pma_interface_clkslip_sel                   ("pld"),
		.hssi_rx_pcs_pma_interface_lpbk_en                       ("disable"),
		.hssi_rx_pcs_pma_interface_master_clk_sel                ("master_rx_pma_clk"),
		.hssi_rx_pcs_pma_interface_silicon_rev                   ("es"),
		.hssi_rx_pcs_pma_interface_pldif_datawidth_mode          ("pldif_data_10bit"),
		.hssi_rx_pcs_pma_interface_pma_dw_rx                     ("pma_10b_rx"),
		.hssi_rx_pcs_pma_interface_pma_if_dft_en                 ("dft_dis"),
		.hssi_rx_pcs_pma_interface_pma_if_dft_val                ("dft_0"),
		.hssi_rx_pcs_pma_interface_prbs_clken                    ("prbs_clk_dis"),
		.hssi_rx_pcs_pma_interface_prbs_ver                      ("prbs_off"),
		.hssi_rx_pcs_pma_interface_prbs9_dwidth                  ("prbs9_64b"),
		.hssi_rx_pcs_pma_interface_prot_mode_rx                  ("eightg_only_pld_mode_rx"),
		.hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion     ("rx_dyn_polinv_dis"),
		.hssi_rx_pcs_pma_interface_rx_lpbk_en                    ("lpbk_dis"),
		.hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok       ("force_sig_ok"),
		.hssi_rx_pcs_pma_interface_rx_prbs_mask                  ("prbsmask128"),
		.hssi_rx_pcs_pma_interface_rx_prbs_mode                  ("teng_mode"),
		.hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel     ("sel_sig_det"),
		.hssi_rx_pcs_pma_interface_rx_static_polarity_inversion  ("rx_stat_polinv_dis"),
		.hssi_rx_pcs_pma_interface_sup_mode                      ("user_mode"),
		.hssi_tx_pcs_pma_interface_bypass_pma_txelecidle         ("true"),
		.hssi_tx_pcs_pma_interface_channel_operation_mode        ("tx_rx_pair_enabled"),
		.hssi_tx_pcs_pma_interface_lpbk_en                       ("disable"),
		.hssi_tx_pcs_pma_interface_master_clk_sel                ("master_tx_pma_clk"),
		.hssi_tx_pcs_pma_interface_silicon_rev                   ("es"),
		.hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx         ("other_prot_mode"),
		.hssi_tx_pcs_pma_interface_pldif_datawidth_mode          ("pldif_data_10bit"),
		.hssi_tx_pcs_pma_interface_pma_dw_tx                     ("pma_10b_tx"),
		.hssi_tx_pcs_pma_interface_pmagate_en                    ("pmagate_dis"),
		.hssi_tx_pcs_pma_interface_prbs_clken                    ("prbs_clk_dis"),
		.hssi_tx_pcs_pma_interface_prbs_gen_pat                  ("prbs_gen_dis"),
		.hssi_tx_pcs_pma_interface_prbs9_dwidth                  ("prbs9_64b"),
		.hssi_tx_pcs_pma_interface_prot_mode_tx                  ("eightg_only_pld_mode_tx"),
		.hssi_tx_pcs_pma_interface_sq_wave_num                   ("sq_wave_default"),
		.hssi_tx_pcs_pma_interface_sqwgen_clken                  ("sqwgen_clk_dis"),
		.hssi_tx_pcs_pma_interface_sup_mode                      ("user_mode"),
		.hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion     ("tx_dyn_polinv_dis"),
		.hssi_tx_pcs_pma_interface_tx_pma_data_sel               ("eight_g_pcs"),
		.hssi_tx_pcs_pma_interface_tx_static_polarity_inversion  ("tx_stat_polinv_dis"),
		.hssi_tx_pcs_pma_interface_uhsif_enable                  ("uhsif_disable"),
		.hssi_tx_pcs_pma_interface_uhsif_index_selection         ("uhsif_index_cram"),
		.hssi_tx_pcs_pma_interface_uhsif_linear_pld_delay_value  (3'b000),
		.hssi_tx_pcs_pma_interface_uhsif_linear_pma_delay_value  (3'b000),
		.hssi_tx_pcs_pma_interface_uhsif_lock_counter_value      (4'b0000),
		.hssi_tx_pcs_pma_interface_uhsif_lock_segment_size       (2'b00),
		.hssi_tx_pcs_pma_interface_uhsif_lock_threshold_value    (4'b0000),
		.hssi_tx_pcs_pma_interface_uhsif_static_index_value      (9'b000000000),
		.hssi_tx_pcs_pma_interface_uhsif_unlock_counter_value    (4'b0000),
		.hssi_tx_pcs_pma_interface_uhsif_unlock_threshold_value  (4'b0000),
		.hssi_common_pcs_pma_interface_asn_clk_enable            ("false"),
		.hssi_common_pcs_pma_interface_asn_enable                ("dis_asn"),
		.hssi_common_pcs_pma_interface_block_sel                 ("eight_g_pcs"),
		.hssi_common_pcs_pma_interface_bypass_early_eios         ("true"),
		.hssi_common_pcs_pma_interface_bypass_pcie_switch        ("true"),
		.hssi_common_pcs_pma_interface_bypass_pma_ltr            ("true"),
		.hssi_common_pcs_pma_interface_bypass_pma_sw_done        ("false"),
		.hssi_common_pcs_pma_interface_bypass_ppm_lock           ("true"),
		.hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp    ("true"),
		.hssi_common_pcs_pma_interface_bypass_txdetectrx         ("true"),
		.hssi_common_pcs_pma_interface_cdr_control               ("dis_cdr_ctrl"),
		.hssi_common_pcs_pma_interface_cid_enable                ("dis_cid_mode"),
		.hssi_common_pcs_pma_interface_data_mask_count           (16'b0000000000000000),
		.hssi_common_pcs_pma_interface_data_mask_count_multi     (3'b000),
		.hssi_common_pcs_pma_interface_early_eios_counter        (8'b00000000),
		.hssi_common_pcs_pma_interface_force_freqdet             ("force_freqdet_dis"),
		.hssi_common_pcs_pma_interface_free_run_clk_enable       ("false"),
		.hssi_common_pcs_pma_interface_ignore_sigdet_g23         ("false"),
		.hssi_common_pcs_pma_interface_silicon_rev               ("es"),
		.hssi_common_pcs_pma_interface_pc_en_counter             (7'b0000000),
		.hssi_common_pcs_pma_interface_pc_rst_counter            (5'b00000),
		.hssi_common_pcs_pma_interface_pcie_hip_mode             ("hip_disable"),
		.hssi_common_pcs_pma_interface_ph_fifo_reg_mode          ("phfifo_reg_mode_dis"),
		.hssi_common_pcs_pma_interface_phfifo_flush_wait         (6'b000000),
		.hssi_common_pcs_pma_interface_pipe_if_g3pcs             ("pipe_if_8gpcs"),
		.hssi_common_pcs_pma_interface_pma_done_counter          (18'b000000000000000000),
		.hssi_common_pcs_pma_interface_pma_if_dft_en             ("dft_dis"),
		.hssi_common_pcs_pma_interface_pma_if_dft_val            ("dft_0"),
		.hssi_common_pcs_pma_interface_ppm_cnt_rst               ("ppm_cnt_rst_dis"),
		.hssi_common_pcs_pma_interface_ppm_deassert_early        ("deassert_early_dis"),
		.hssi_common_pcs_pma_interface_ppm_gen1_2_cnt            ("cnt_32k"),
		.hssi_common_pcs_pma_interface_ppm_post_eidle_delay      ("cnt_400_cycles"),
		.hssi_common_pcs_pma_interface_ppmsel                    ("ppmsel_1000"),
		.hssi_common_pcs_pma_interface_prot_mode                 ("other_protocols"),
		.hssi_common_pcs_pma_interface_rxvalid_mask              ("rxvalid_mask_dis"),
		.hssi_common_pcs_pma_interface_sigdet_wait_counter       (12'b000000000000),
		.hssi_common_pcs_pma_interface_sigdet_wait_counter_multi (3'b000),
		.hssi_common_pcs_pma_interface_sim_mode                  ("disable"),
		.hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en   ("false"),
		.hssi_common_pcs_pma_interface_sup_mode                  ("user_mode"),
		.hssi_common_pcs_pma_interface_testout_sel               ("ppm_det_test"),
		.hssi_common_pcs_pma_interface_wait_clk_on_off_timer     (4'b0000),
		.hssi_common_pcs_pma_interface_wait_pipe_synchronizing   (5'b00000),
		.hssi_common_pcs_pma_interface_wait_send_syncp_fbkp      (11'b00000000000),
		.hssi_fifo_rx_pcs_double_read_mode                       ("double_read_dis"),
		.hssi_fifo_rx_pcs_prot_mode                              ("non_teng_mode"),
		.hssi_fifo_rx_pcs_silicon_rev                            ("es"),
		.hssi_fifo_tx_pcs_double_write_mode                      ("double_write_dis"),
		.hssi_fifo_tx_pcs_prot_mode                              ("non_teng_mode"),
		.hssi_fifo_tx_pcs_silicon_rev                            ("es"),
		.hssi_pipe_gen3_bypass_rx_detection_enable               ("false"),
		.hssi_pipe_gen3_bypass_rx_preset                         (3'b000),
		.hssi_pipe_gen3_bypass_rx_preset_enable                  ("false"),
		.hssi_pipe_gen3_bypass_tx_coefficent                     (18'b000000000000000000),
		.hssi_pipe_gen3_bypass_tx_coefficent_enable              ("false"),
		.hssi_pipe_gen3_elecidle_delay_g3                        (3'b000),
		.hssi_pipe_gen3_ind_error_reporting                      ("dis_ind_error_reporting"),
		.hssi_pipe_gen3_mode                                     ("disable_pcs"),
		.hssi_pipe_gen3_phy_status_delay_g12                     (3'b000),
		.hssi_pipe_gen3_phy_status_delay_g3                      (3'b000),
		.hssi_pipe_gen3_phystatus_rst_toggle_g12                 ("en_phystatus_rst_toggle"),
		.hssi_pipe_gen3_phystatus_rst_toggle_g3                  ("dis_phystatus_rst_toggle_g3"),
		.hssi_pipe_gen3_rate_match_pad_insertion                 ("en_rm_fifo_pad_ins"),
		.hssi_pipe_gen3_sup_mode                                 ("user_mode"),
		.hssi_pipe_gen3_test_out_sel                             ("disable_test_out"),
		.hssi_pipe_gen3_silicon_rev                              ("es"),
		.hssi_pipe_gen1_2_elec_idle_delay_val                    (3'b000),
		.hssi_pipe_gen1_2_error_replace_pad                      ("replace_edb"),
		.hssi_pipe_gen1_2_hip_mode                               ("dis_hip"),
		.hssi_pipe_gen1_2_ind_error_reporting                    ("dis_ind_error_reporting"),
		.hssi_pipe_gen1_2_phystatus_delay_val                    (3'b000),
		.hssi_pipe_gen1_2_phystatus_rst_toggle                   ("dis_phystatus_rst_toggle"),
		.hssi_pipe_gen1_2_pipe_byte_de_serializer_en             ("dont_care_bds"),
		.hssi_pipe_gen1_2_prot_mode                              ("disabled_prot_mode"),
		.hssi_pipe_gen1_2_rpre_emph_a_val                        (6'b000000),
		.hssi_pipe_gen1_2_rpre_emph_b_val                        (6'b000000),
		.hssi_pipe_gen1_2_rpre_emph_c_val                        (6'b000000),
		.hssi_pipe_gen1_2_rpre_emph_d_val                        (6'b000000),
		.hssi_pipe_gen1_2_rpre_emph_e_val                        (6'b000000),
		.hssi_pipe_gen1_2_rvod_sel_a_val                         (6'b000000),
		.hssi_pipe_gen1_2_rvod_sel_b_val                         (6'b000000),
		.hssi_pipe_gen1_2_rvod_sel_c_val                         (6'b000000),
		.hssi_pipe_gen1_2_rvod_sel_d_val                         (6'b000000),
		.hssi_pipe_gen1_2_rvod_sel_e_val                         (6'b000000),
		.hssi_pipe_gen1_2_rx_pipe_enable                         ("dis_pipe_rx"),
		.hssi_pipe_gen1_2_rxdetect_bypass                        ("dis_rxdetect_bypass"),
		.hssi_pipe_gen1_2_sup_mode                               ("user_mode"),
		.hssi_pipe_gen1_2_tx_pipe_enable                         ("dis_pipe_tx"),
		.hssi_pipe_gen1_2_txswing                                ("dis_txswing"),
		.hssi_pipe_gen1_2_silicon_rev                            ("es"),
		.cdr_pll_bw_sel                                          ("low"),
		.cdr_pll_cdr_cmu_mode                                    ("cdr_mode"),
		.cdr_pll_clklow_mux_select                               ("clklow_mux_cdr_fbclk"),
		.cdr_pll_disable_up_dn                                   ("true"),
		.cdr_pll_fref_clklow_div                                 (1),
		.cdr_pll_fref_mux_select                                 ("fref_mux_cdr_refclk"),
		.cdr_pll_gpon_lck2ref_control                            ("gpon_lck2ref_off"),
		.cdr_pll_loopback_mode                                   ("loopback_recovered_data"),
		.cdr_pll_ltd_ltr_micro_controller_select                 ("ltd_ltr_pcs"),
		.cdr_pll_m_counter                                       (5),
		.cdr_pll_n_counter                                       (1),
		.cdr_pll_op_mode                                         ("normal"),
		.cdr_pll_pcie_gen                                        ("non_pcie"),
		.cdr_pll_pd_fastlock_mode                                ("false"),
		.cdr_pll_pd_l_counter                                    (4),
		.cdr_pll_pfd_l_counter                                   (4),
		.cdr_pll_prot_mode                                       ("basic"),
		.cdr_pll_reverse_serial_loopback                         ("no_loopback"),
		.cdr_pll_txpll_hclk_driver_enable                        ("false"),
		.cdr_pll_fb_select                                       ("direct_fb"),
		.cdr_pll_iqclk_mux_sel                                   ("power_down"),
		.cdr_pll_datarate                                        ("1250 Mbps"),
		.cdr_pll_reference_clock_frequency                       ("125.000000 MHz"),
		.cdr_pll_silicon_rev                                     ("es"),
		.cdr_pll_output_clock_frequency                          ("625 MHz"),
		.cdr_pll_pma_width                                       (10),
		.cdr_pll_cgb_div                                         (1),
		.cdr_pll_is_cascaded_pll                                 ("false"),
		.pma_cdr_refclk_receiver_detect_src                      ("iqclk_src"),
		.pma_cdr_refclk_xmux_refclk_src                          ("refclk_iqclk"),
		.pma_cdr_refclk_xpm_iqref_mux_iqclk_sel                  ("power_down"),
		.pma_cdr_refclk_refclk_select                            ("ref_iqclk1"),
		.pma_cdr_refclk_silicon_rev                              ("es"),
		.pma_cgb_bonding_mode                                    ("x1_non_bonded"),
		.pma_cgb_bonding_reset_enable                            ("disallow_bonding_reset"),
		.pma_cgb_cgb_enable_iqtxrxclk                            ("disable_iqtxrxclk"),
		.pma_cgb_pcie_gen3_bitwidth                              ("pciegen3_wide"),
		.pma_cgb_proc_mode                                       ("basic"),
		.pma_cgb_select_done_master_or_slave                     ("choose_slave_pcie_sw_done"),
		.pma_cgb_ser_mode                                        ("ten_bit"),
		.pma_cgb_tx_ucontrol_reset_pcie                          ("pcscorehip_controls_tx"),
		.pma_cgb_x1_div_m_sel                                    ("divbypass"),
		.pma_cgb_data_rate                                       ("1250 Mbps"),
		.pma_cgb_silicon_rev                                     ("es"),
		.pma_cgb_input_select_x1                                 ("lcpll_bot"),
		.pma_cgb_input_select_gen3                               ("unused"),
		.pma_cgb_input_select_xn                                 ("unused"),
		.pma_rx_deser_pcie_gen                                   ("non_pcie"),
		.pma_rx_deser_clk_user                                   ("clk_user_33"),
		.pma_rx_deser_clkdiv_source                              ("vco_bypass_normal"),
		.pma_rx_deser_clkdivrx_user_mode                         ("clkdivrx_user_div33"),
		.pma_rx_deser_datawidth                                  ("dwidth_10"),
		.pma_rx_deser_deser_factor                               (10),
		.pma_rx_deser_deser_powerdown                            ("deser_power_up"),
		.pma_rx_deser_op_mode                                    ("enabled"),
		.pma_rx_deser_sdclk_enable                               ("true"),
		.pma_rx_deser_silicon_rev                                ("es"),
		.pma_rx_dfe_atb_select                                   ("atb_disable"),
		.pma_rx_dfe_datarate_mode                                ("low_datarate"),
		.pma_rx_dfe_dft_en                                       ("dft_disable"),
		.pma_rx_dfe_op_mode                                      ("cdr_mode"),
		.pma_rx_dfe_pdb                                          ("dfe_powerdown"),
		.pma_rx_dfe_pdb_fixedtap                                 ("fixtap_dfe_powerdown"),
		.pma_rx_dfe_pdb_floattap                                 ("floattap_dfe_powerdown"),
		.pma_rx_dfe_uc_rx_dfe_cal                                ("uc_rx_dfe_cal_off"),
		.pma_rx_dfe_uc_rx_dfe_cal_status                         ("uc_rx_dfe_cal_notdone"),
		.pma_rx_dfe_silicon_rev                                  ("es"),
		.pma_rx_odi_silicon_rev                                  ("es"),
		.pma_rx_buf_bypass_eqz_stages_234                        ("bypass_off"),
		.pma_rx_buf_cdrclk_to_cgb                                ("cdrclk_2cgb_dis"),
		.pma_rx_buf_op_mode                                      ("normal"),
		.pma_rx_buf_pdb_rx                                       ("normal_rx_on"),
		.pma_rx_buf_proc_mode                                    ("basic"),
		.pma_rx_buf_qpi_enable                                   ("non_qpi_mode"),
		.pma_rx_buf_rx_refclk_divider                            ("bypass_divider"),
		.pma_rx_buf_rx_refclk_en                                 ("refclk_dis"),
		.pma_rx_buf_uc_cal_enable                                ("rx_cal_off"),
		.pma_rx_buf_uc_rx_rstb                                   ("rx_reset_on"),
		.pma_rx_buf_silicon_rev                                  ("es"),
		.pma_rx_sd_op_mode                                       ("pwr_down"),
		.pma_rx_sd_optimal_setting                               ("true"),
		.pma_rx_sd_proc_mode                                     ("pcie_gen1"),
		.pma_rx_sd_sd_output_off                                 (1),
		.pma_rx_sd_sd_output_on                                  (15),
		.pma_rx_sd_sd_pdb                                        ("false"),
		.pma_rx_sd_sd_threshold                                  (3),
		.pma_rx_sd_silicon_rev                                   ("es"),
		.pma_tx_ser_ser_clk_divtx_user_sel                       ("divtx_user_33"),
		.pma_tx_ser_silicon_rev                                  ("es"),
		.pma_tx_buf_proc_mode                                    ("basic"),
		.pma_tx_buf_rx_det                                       ("mode_1"),
		.pma_tx_buf_rx_det_output_sel                            ("rx_det_qpi_out"),
		.pma_tx_buf_rx_det_pdb                                   ("rx_det_off"),
		.pma_tx_buf_uc_gen3                                      ("gen3_off"),
		.pma_tx_buf_uc_gen4                                      ("gen4_off"),
		.pma_tx_buf_uc_txvod_cal                                 ("uc_tx_vod_cal_off"),
		.pma_tx_buf_uc_txvod_cal_status                          ("uc_tx_vod_cal_notdone"),
		.pma_tx_buf_silicon_rev                                  ("es")
	) native_gige_1588_inst (
		.tx_analogreset            (tx_analogreset),                                                       //            tx_analogreset.tx_analogreset
		.tx_digitalreset           (tx_digitalreset),                                                      //           tx_digitalreset.tx_digitalreset
		.rx_analogreset            (rx_analogreset),                                                       //            rx_analogreset.rx_analogreset
		.rx_digitalreset           (rx_digitalreset),                                                      //           rx_digitalreset.rx_digitalreset
		.tx_cal_busy               (tx_cal_busy),                                                          //               tx_cal_busy.tx_cal_busy
		.rx_cal_busy               (rx_cal_busy),                                                          //               rx_cal_busy.rx_cal_busy
		.tx_serial_clk0            (tx_serial_clk0),                                                       //            tx_serial_clk0.clk
		.tx_serial_clk1            (tx_serial_clk1),                                                       //            tx_serial_clk1.clk
		.rx_cdr_refclk0            (rx_cdr_refclk0),                                                       //            rx_cdr_refclk0.clk
		.rx_cdr_refclk1            (rx_cdr_refclk1),                                                       //            rx_cdr_refclk1.clk
		.tx_serial_data            (tx_serial_data),                                                       //            tx_serial_data.tx_serial_data
		.rx_serial_data            (rx_serial_data),                                                       //            rx_serial_data.rx_serial_data
		.rx_pma_clkslip            (rx_pma_clkslip),                                                       //            rx_pma_clkslip.rx_pma_clkslip
		.rx_seriallpbken           (rx_seriallpbken),                                                      //           rx_seriallpbken.rx_seriallpbken
		.rx_set_locktodata         (rx_set_locktodata),                                                    //         rx_set_locktodata.rx_set_locktodata
		.rx_set_locktoref          (rx_set_locktoref),                                                     //          rx_set_locktoref.rx_set_locktoref
		.rx_is_lockedtoref         (rx_is_lockedtoref),                                                    //         rx_is_lockedtoref.rx_is_lockedtoref
		.rx_is_lockedtodata        (rx_is_lockedtodata),                                                   //        rx_is_lockedtodata.rx_is_lockedtodata
		.tx_coreclkin              (tx_coreclkin),                                                         //              tx_coreclkin.clk
		.rx_coreclkin              (rx_coreclkin),                                                         //              rx_coreclkin.clk
		.tx_clkout                 (tx_clkout),                                                            //                 tx_clkout.clk
		.rx_clkout                 (rx_clkout),                                                            //                 rx_clkout.clk
		.tx_pma_clkout             (tx_pma_clkout),                                                        //             tx_pma_clkout.clk
		.tx_pma_div_clkout         (tx_pma_div_clkout),                                                    //         tx_pma_div_clkout.clk
		.rx_pma_clkout             (rx_pma_clkout),                                                        //             rx_pma_clkout.clk
		.rx_pma_div_clkout         (rx_pma_div_clkout),                                                    //         rx_pma_div_clkout.clk
		.tx_parallel_data          (tx_parallel_data),                                                     //          tx_parallel_data.tx_parallel_data
		.tx_control                (tx_control),                                                           //                tx_control.tx_control
		.rx_parallel_data          (rx_parallel_data),                                                     //          rx_parallel_data.rx_parallel_data
		.rx_control                (rx_control),                                                           //                rx_control.rx_control
		.rx_bitslip                (rx_bitslip),                                                           //                rx_bitslip.rx_bitslip
		.tx_std_pcfifo_full        (tx_std_pcfifo_full),                                                   //        tx_std_pcfifo_full.tx_std_pcfifo_full
		.tx_std_pcfifo_empty       (tx_std_pcfifo_empty),                                                  //       tx_std_pcfifo_empty.tx_std_pcfifo_empty
		.rx_std_pcfifo_full        (rx_std_pcfifo_full),                                                   //        rx_std_pcfifo_full.rx_std_pcfifo_full
		.rx_std_pcfifo_empty       (rx_std_pcfifo_empty),                                                  //       rx_std_pcfifo_empty.rx_std_pcfifo_empty
		.rx_std_bitrev_ena         (rx_std_bitrev_ena),                                                    //         rx_std_bitrev_ena.rx_std_bitrev_ena
		.tx_polinv                 (tx_polinv),                                                            //                 tx_polinv.tx_polinv
		.rx_polinv                 (rx_polinv),                                                            //                 rx_polinv.rx_polinv
		.rx_std_bitslipboundarysel (rx_std_bitslipboundarysel),                                            // rx_std_bitslipboundarysel.rx_std_bitslipboundarysel
		.tx_std_elecidle           (tx_std_elecidle),                                                      //           tx_std_elecidle.tx_std_elecidle
		.tx_enh_data_valid         (tx_enh_data_valid),                                                    //         tx_enh_data_valid.tx_enh_data_valid
		.tx_enh_fifo_full          (tx_enh_fifo_full),                                                     //          tx_enh_fifo_full.tx_enh_fifo_full
		.tx_enh_fifo_cnt           (tx_enh_fifo_cnt),                                                      //           tx_enh_fifo_cnt.tx_enh_fifo_cnt
		.rx_enh_data_valid         (rx_enh_data_valid),                                                    //         rx_enh_data_valid.rx_enh_data_valid
		.rx_enh_fifo_full          (rx_enh_fifo_full),                                                     //          rx_enh_fifo_full.rx_enh_fifo_full
		.rx_enh_fifo_del           (rx_enh_fifo_del),                                                      //           rx_enh_fifo_del.rx_enh_fifo_del
		.rx_enh_fifo_insert        (rx_enh_fifo_insert),                                                   //        rx_enh_fifo_insert.rx_enh_fifo_insert
		.rx_enh_fifo_cnt           (rx_enh_fifo_cnt),                                                      //           rx_enh_fifo_cnt.rx_enh_fifo_cnt
		.rx_enh_highber            (rx_enh_highber),                                                       //            rx_enh_highber.rx_enh_highber
		.rx_enh_highber_clr_cnt    (rx_enh_highber_clr_cnt),                                               //    rx_enh_highber_clr_cnt.rx_enh_highber_clr_cnt
		.rx_enh_clr_errblk_count   (rx_enh_clr_errblk_count),                                              //   rx_enh_clr_errblk_count.rx_enh_clr_errblk_count
		.rx_enh_blk_lock           (rx_enh_blk_lock),                                                      //           rx_enh_blk_lock.rx_enh_blk_lock
		.reconfig_clk              (reconfig_clk),                                                         //              reconfig_clk.clk
		.reconfig_reset            (reconfig_reset),                                                       //            reconfig_reset.reset
		.reconfig_write            (reconfig_write),                                                       //             reconfig_avmm.write
		.reconfig_read             (reconfig_read),                                                        //                          .read
		.reconfig_address          (reconfig_address),                                                     //                          .address
		.reconfig_writedata        (reconfig_writedata),                                                   //                          .writedata
		.reconfig_readdata         (reconfig_readdata),                                                    //                          .readdata
		.reconfig_waitrequest      (reconfig_waitrequest),                                                 //                          .waitrequest
		.tx_serial_clk2            (1'b0),                                                                 //               (terminated)
		.tx_serial_clk3            (1'b0),                                                                 //               (terminated)
		.tx_bonding_clocks         (6'b000000),                                                            //               (terminated)
		.rx_cdr_refclk2            (1'b0),                                                                 //               (terminated)
		.rx_cdr_refclk3            (1'b0),                                                                 //               (terminated)
		.rx_cdr_refclk4            (1'b0),                                                                 //               (terminated)
		.tx_pma_clkslip            (1'b0),                                                                 //               (terminated)
		.rx_pma_qpipullup          (1'b0),                                                                 //               (terminated)
		.tx_pma_qpipulldn          (1'b0),                                                                 //               (terminated)
		.tx_pma_qpipullup          (1'b0),                                                                 //               (terminated)
		.tx_pma_txdetectrx         (1'b0),                                                                 //               (terminated)
		.tx_pma_rxfound            (),                                                                     //               (terminated)
		.rx_clklow                 (),                                                                     //               (terminated)
		.rx_fref                   (),                                                                     //               (terminated)
		.rx_prbs_err_clr           (1'b0),                                                                 //               (terminated)
		.rx_prbs_done              (),                                                                     //               (terminated)
		.rx_prbs_err               (),                                                                     //               (terminated)
		.tx_uhsif_clk              (1'b0),                                                                 //               (terminated)
		.tx_uhsif_clkout           (),                                                                     //               (terminated)
		.tx_uhsif_ctrl             (3'b000),                                                               //               (terminated)
		.tx_uhsif_status           (),                                                                     //               (terminated)
		.rx_std_byterev_ena        (1'b0),                                                                 //               (terminated)
		.tx_std_bitslipboundarysel (5'b00000),                                                             //               (terminated)
		.rx_std_wa_patternalign    (1'b0),                                                                 //               (terminated)
		.rx_std_wa_a1a2size        (1'b0),                                                                 //               (terminated)
		.rx_std_rmfifo_full        (),                                                                     //               (terminated)
		.rx_std_rmfifo_empty       (),                                                                     //               (terminated)
		.rx_std_signaldetect       (),                                                                     //               (terminated)
		.tx_enh_fifo_pfull         (),                                                                     //               (terminated)
		.tx_enh_fifo_empty         (),                                                                     //               (terminated)
		.tx_enh_fifo_pempty        (),                                                                     //               (terminated)
		.rx_enh_fifo_rd_en         (1'b0),                                                                 //               (terminated)
		.rx_enh_fifo_pfull         (),                                                                     //               (terminated)
		.rx_enh_fifo_empty         (),                                                                     //               (terminated)
		.rx_enh_fifo_pempty        (),                                                                     //               (terminated)
		.rx_enh_fifo_align_val     (),                                                                     //               (terminated)
		.rx_enh_fifo_align_clr     (1'b0),                                                                 //               (terminated)
		.tx_enh_frame              (),                                                                     //               (terminated)
		.tx_enh_frame_burst_en     (1'b0),                                                                 //               (terminated)
		.tx_enh_frame_diag_status  (2'b00),                                                                //               (terminated)
		.rx_enh_frame              (),                                                                     //               (terminated)
		.rx_enh_frame_lock         (),                                                                     //               (terminated)
		.rx_enh_frame_diag_status  (),                                                                     //               (terminated)
		.rx_enh_crc32_err          (),                                                                     //               (terminated)
		.tx_enh_bitslip            (7'b0000000),                                                           //               (terminated)
		.tx_hip_data               (64'b0000000000000000000000000000000000000000000000000000000000000000), //               (terminated)
		.rx_hip_data               (),                                                                     //               (terminated)
		.hip_pipe_pclk             (),                                                                     //               (terminated)
		.hip_fixedclk              (),                                                                     //               (terminated)
		.hip_frefclk               (),                                                                     //               (terminated)
		.hip_ctrl                  (),                                                                     //               (terminated)
		.hip_cal_done              (),                                                                     //               (terminated)
		.pipe_rate                 (2'b00),                                                                //               (terminated)
		.pipe_sw_done              (2'b00),                                                                //               (terminated)
		.pipe_sw                   (),                                                                     //               (terminated)
		.pipe_hclk_in              (1'b0),                                                                 //               (terminated)
		.pipe_hclk_out             (),                                                                     //               (terminated)
		.pipe_g3_txdeemph          (18'b000000000000000000),                                               //               (terminated)
		.pipe_g3_rxpresethint      (3'b000),                                                               //               (terminated)
		.pipe_rx_eidleinfersel     (3'b000),                                                               //               (terminated)
		.pipe_rx_elecidle          (),                                                                     //               (terminated)
		.pipe_rx_polarity          (1'b0)                                                                  //               (terminated)
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2013 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_xcvr_native_vi" version="13.1" >
// Retrieval info: 	<generic name="device_family" value="Arria 10" />
// Retrieval info: 	<generic name="device_speedgrade" value="fastest" />
// Retrieval info: 	<generic name="message_level" value="error" />
// Retrieval info: 	<generic name="support_mode" value="user_mode" />
// Retrieval info: 	<generic name="duplex_mode" value="duplex" />
// Retrieval info: 	<generic name="datapath_select" value="Standard" />
// Retrieval info: 	<generic name="channels" value="1" />
// Retrieval info: 	<generic name="set_data_rate" value="1250" />
// Retrieval info: 	<generic name="rcfg_iface_enable" value="1" />
// Retrieval info: 	<generic name="enable_simple_interface" value="0" />
// Retrieval info: 	<generic name="enable_split_interface" value="0" />
// Retrieval info: 	<generic name="bonded_mode" value="not_bonded" />
// Retrieval info: 	<generic name="set_pcs_bonding_master" value="Auto" />
// Retrieval info: 	<generic name="tx_pma_clk_div" value="1" />
// Retrieval info: 	<generic name="plls" value="2" />
// Retrieval info: 	<generic name="pll_select" value="1" />
// Retrieval info: 	<generic name="enable_port_tx_pma_clkout" value="1" />
// Retrieval info: 	<generic name="enable_port_tx_pma_div_clkout" value="1" />
// Retrieval info: 	<generic name="tx_pma_div_clkout_divider" value="33" />
// Retrieval info: 	<generic name="enable_port_tx_pma_clkslip" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_pma_qpipullup" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_pma_qpipulldn" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_pma_txdetectrx" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_pma_rxfound" value="0" />
// Retrieval info: 	<generic name="cdr_refclk_cnt" value="2" />
// Retrieval info: 	<generic name="cdr_refclk_select" value="1" />
// Retrieval info: 	<generic name="set_cdr_refclk_freq" value="125.000000" />
// Retrieval info: 	<generic name="rx_ppm_detect_threshold" value="1000" />
// Retrieval info: 	<generic name="rx_pma_dfe_mode" value="Disabled" />
// Retrieval info: 	<generic name="enable_port_rx_pma_clkout" value="1" />
// Retrieval info: 	<generic name="enable_port_rx_pma_div_clkout" value="1" />
// Retrieval info: 	<generic name="rx_pma_div_clkout_divider" value="33" />
// Retrieval info: 	<generic name="enable_port_rx_pma_clkslip" value="1" />
// Retrieval info: 	<generic name="enable_port_rx_pma_qpipullup" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_is_lockedtodata" value="1" />
// Retrieval info: 	<generic name="enable_port_rx_is_lockedtoref" value="1" />
// Retrieval info: 	<generic name="enable_ports_rx_manual_cdr_mode" value="1" />
// Retrieval info: 	<generic name="enable_port_rx_signaldetect" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_seriallpbken" value="1" />
// Retrieval info: 	<generic name="enable_ports_rx_prbs" value="0" />
// Retrieval info: 	<generic name="std_protocol_mode" value="gige_1588" />
// Retrieval info: 	<generic name="std_pcs_pma_width" value="10" />
// Retrieval info: 	<generic name="std_low_latency_bypass_enable" value="0" />
// Retrieval info: 	<generic name="enable_hip" value="0" />
// Retrieval info: 	<generic name="enable_hard_reset" value="0" />
// Retrieval info: 	<generic name="std_tx_pcfifo_mode" value="register_fifo" />
// Retrieval info: 	<generic name="std_tx_pcfifo_fast" value="0" />
// Retrieval info: 	<generic name="std_rx_pcfifo_mode" value="register_fifo" />
// Retrieval info: 	<generic name="enable_port_tx_std_pcfifo_full" value="1" />
// Retrieval info: 	<generic name="enable_port_tx_std_pcfifo_empty" value="1" />
// Retrieval info: 	<generic name="enable_port_rx_std_pcfifo_full" value="1" />
// Retrieval info: 	<generic name="enable_port_rx_std_pcfifo_empty" value="1" />
// Retrieval info: 	<generic name="std_tx_byte_ser_mode" value="Disabled" />
// Retrieval info: 	<generic name="std_rx_byte_deser_mode" value="Disabled" />
// Retrieval info: 	<generic name="std_tx_8b10b_enable" value="1" />
// Retrieval info: 	<generic name="std_tx_8b10b_disp_ctrl_enable" value="0" />
// Retrieval info: 	<generic name="std_rx_8b10b_enable" value="1" />
// Retrieval info: 	<generic name="std_rx_rmfifo_mode" value="disabled" />
// Retrieval info: 	<generic name="std_rx_rmfifo_pattern_n" value="0" />
// Retrieval info: 	<generic name="std_rx_rmfifo_pattern_p" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_std_rmfifo_full" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_std_rmfifo_empty" value="0" />
// Retrieval info: 	<generic name="pcie_rate_match" value="Bypass" />
// Retrieval info: 	<generic name="std_tx_bitslip_enable" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_std_bitslipboundarysel" value="0" />
// Retrieval info: 	<generic name="std_rx_word_aligner_mode" value="synchronous state machine" />
// Retrieval info: 	<generic name="std_rx_word_aligner_pattern_len" value="10" />
// Retrieval info: 	<generic name="std_rx_word_aligner_pattern" value="380" />
// Retrieval info: 	<generic name="std_rx_word_aligner_rknumber" value="3" />
// Retrieval info: 	<generic name="std_rx_word_aligner_renumber" value="3" />
// Retrieval info: 	<generic name="std_rx_word_aligner_rgnumber" value="3" />
// Retrieval info: 	<generic name="enable_port_rx_std_wa_patternalign" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_std_wa_a1a2size" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_std_bitslipboundarysel" value="1" />
// Retrieval info: 	<generic name="enable_port_rx_std_bitslip" value="0" />
// Retrieval info: 	<generic name="std_tx_bitrev_enable" value="0" />
// Retrieval info: 	<generic name="std_tx_byterev_enable" value="0" />
// Retrieval info: 	<generic name="std_tx_polinv_enable" value="0" />
// Retrieval info: 	<generic name="std_rx_bitrev_enable" value="0" />
// Retrieval info: 	<generic name="std_rx_byterev_enable" value="0" />
// Retrieval info: 	<generic name="std_rx_polinv_enable" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_polinv" value="1" />
// Retrieval info: 	<generic name="enable_port_rx_std_bitrev_ena" value="1" />
// Retrieval info: 	<generic name="enable_port_rx_std_byterev_ena" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_polinv" value="1" />
// Retrieval info: 	<generic name="enable_port_tx_std_elecidle" value="1" />
// Retrieval info: 	<generic name="enable_port_rx_std_signaldetect" value="0" />
// Retrieval info: 	<generic name="enable_ports_pipe_sw" value="0" />
// Retrieval info: 	<generic name="enable_ports_pipe_hclk" value="0" />
// Retrieval info: 	<generic name="enable_ports_pipe_g3_analog" value="0" />
// Retrieval info: 	<generic name="enable_ports_pipe_rx_elecidle" value="0" />
// Retrieval info: 	<generic name="enable_port_pipe_rx_polarity" value="0" />
// Retrieval info: 	<generic name="enh_protocol_mode" value="teng_1588_mode" />
// Retrieval info: 	<generic name="enh_pcs_pma_width" value="40" />
// Retrieval info: 	<generic name="enh_pld_pcs_width" value="66" />
// Retrieval info: 	<generic name="enh_txfifo_mode" value="Register" />
// Retrieval info: 	<generic name="enh_txfifo_full" value="15" />
// Retrieval info: 	<generic name="enh_txfifo_empty" value="0" />
// Retrieval info: 	<generic name="enh_txfifo_pfull" value="13" />
// Retrieval info: 	<generic name="enh_txfifo_pempty" value="2" />
// Retrieval info: 	<generic name="enable_port_tx_enh_fifo_full" value="1" />
// Retrieval info: 	<generic name="enable_port_tx_enh_fifo_pfull" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_enh_fifo_empty" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_enh_fifo_pempty" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_enh_fifo_cnt" value="1" />
// Retrieval info: 	<generic name="enh_rxfifo_mode" value="Register" />
// Retrieval info: 	<generic name="enh_rxfifo_full" value="31" />
// Retrieval info: 	<generic name="enh_rxfifo_empty" value="0" />
// Retrieval info: 	<generic name="enh_rxfifo_pfull" value="23" />
// Retrieval info: 	<generic name="enh_rxfifo_pempty" value="2" />
// Retrieval info: 	<generic name="enh_rxfifo_align_del" value="0" />
// Retrieval info: 	<generic name="enh_rxfifo_control_del" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_enh_data_valid" value="1" />
// Retrieval info: 	<generic name="enable_port_rx_enh_fifo_full" value="1" />
// Retrieval info: 	<generic name="enable_port_rx_enh_fifo_pfull" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_enh_fifo_empty" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_enh_fifo_pempty" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_enh_fifo_cnt" value="1" />
// Retrieval info: 	<generic name="enable_port_rx_enh_fifo_del" value="1" />
// Retrieval info: 	<generic name="enable_port_rx_enh_fifo_insert" value="1" />
// Retrieval info: 	<generic name="enable_port_rx_enh_fifo_rd_en" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_enh_fifo_align_val" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_enh_fifo_align_clr" value="0" />
// Retrieval info: 	<generic name="enh_tx_frmgen_enable" value="0" />
// Retrieval info: 	<generic name="enh_tx_frmgen_mfrm_length" value="2048" />
// Retrieval info: 	<generic name="enh_tx_frmgen_burst_enable" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_enh_frame" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_enh_frame_diag_status" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_enh_frame_burst_en" value="0" />
// Retrieval info: 	<generic name="enh_rx_frmsync_enable" value="0" />
// Retrieval info: 	<generic name="enh_rx_frmsync_mfrm_length" value="2048" />
// Retrieval info: 	<generic name="enable_port_rx_enh_frame" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_enh_frame_lock" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_enh_frame_diag_status" value="0" />
// Retrieval info: 	<generic name="enh_tx_crcgen_enable" value="0" />
// Retrieval info: 	<generic name="enh_rx_crcchk_enable" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_enh_crc32_err" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_enh_highber" value="1" />
// Retrieval info: 	<generic name="enable_port_rx_enh_highber_clr_cnt" value="1" />
// Retrieval info: 	<generic name="enable_port_rx_enh_clr_errblk_count" value="1" />
// Retrieval info: 	<generic name="enh_tx_64b66b_enable" value="1" />
// Retrieval info: 	<generic name="enh_rx_64b66b_enable" value="1" />
// Retrieval info: 	<generic name="enh_tx_sh_err" value="0" />
// Retrieval info: 	<generic name="enh_tx_scram_enable" value="1" />
// Retrieval info: 	<generic name="enh_tx_scram_seed" value="288230376151711743" />
// Retrieval info: 	<generic name="enh_rx_descram_enable" value="1" />
// Retrieval info: 	<generic name="enh_tx_dispgen_enable" value="0" />
// Retrieval info: 	<generic name="enh_rx_dispchk_enable" value="0" />
// Retrieval info: 	<generic name="enh_rx_blksync_enable" value="1" />
// Retrieval info: 	<generic name="enable_port_rx_enh_blk_lock" value="1" />
// Retrieval info: 	<generic name="enh_tx_bitslip_enable" value="0" />
// Retrieval info: 	<generic name="enh_tx_polinv_enable" value="0" />
// Retrieval info: 	<generic name="enh_rx_bitslip_enable" value="0" />
// Retrieval info: 	<generic name="enh_rx_polinv_enable" value="0" />
// Retrieval info: 	<generic name="enable_port_tx_enh_bitslip" value="0" />
// Retrieval info: 	<generic name="enable_port_rx_enh_bitslip" value="1" />
// Retrieval info: 	<generic name="generate_docs" value="1" />
// Retrieval info: 	<generic name="generate_add_hdl_instance_example" value="0" />
// Retrieval info: 	<generic name="rcfg_enable" value="1" />
// Retrieval info: 	<generic name="rcfg_shared" value="0" />
// Retrieval info: 	<generic name="rcfg_jtag_enable" value="0" />
// Retrieval info: 	<generic name="rcfg_file_prefix" value="gige_1588" />
// Retrieval info: 	<generic name="rcfg_sv_file_enable" value="1" />
// Retrieval info: 	<generic name="rcfg_h_file_enable" value="1" />
// Retrieval info: 	<generic name="rcfg_txt_file_enable" value="0" />
// Retrieval info: 	<generic name="rcfg_mif_file_enable" value="1" />
// Retrieval info: 	<generic name="rcfg_multi_enable" value="0" />
// Retrieval info: 	<generic name="rcfg_profile_cnt" value="2" />
// Retrieval info: 	<generic name="rcfg_profile_select" value="1" />
// Retrieval info: 	<generic name="rcfg_param_vals1" value="" />
// Retrieval info: 	<generic name="rcfg_param_vals2" value="" />
// Retrieval info: 	<generic name="rcfg_param_vals3" value="" />
// Retrieval info: 	<generic name="rcfg_param_vals4" value="" />
// Retrieval info: 	<generic name="rcfg_param_vals5" value="" />
// Retrieval info: 	<generic name="rcfg_param_vals6" value="" />
// Retrieval info: 	<generic name="rcfg_param_vals7" value="" />
// Retrieval info: 	<generic name="AUTO_TX_SERIAL_CLK0_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_TX_SERIAL_CLK1_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_TX_SERIAL_CLK2_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_TX_SERIAL_CLK3_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_RX_CDR_REFCLK0_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_RX_CDR_REFCLK1_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_RX_CDR_REFCLK2_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_RX_CDR_REFCLK3_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_RX_CDR_REFCLK4_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_TX_CORECLKIN_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_RX_CORECLKIN_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_TX_UHSIF_CLK_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_PIPE_HCLK_IN_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_RECONFIG_CLK_CLOCK_RATE" value="-1" />
// Retrieval info: </instance>
// IPFS_FILES : native_gige_1588.vo
// RELATED_FILES: native_gige_1588.v, altera_xcvr_functions.sv, alt_xcvr_resync.sv, twentynm_pcs.sv, twentynm_pcs_ch.sv, twentynm_pma.sv, twentynm_pma_ch.sv, twentynm_xcvr_avmm.sv, twentynm_xcvr_native.sv, twentynm_hssi_10g_rx_pcs_rbc.sv, twentynm_hssi_10g_tx_pcs_rbc.sv, twentynm_hssi_8g_rx_pcs_rbc.sv, twentynm_hssi_8g_tx_pcs_rbc.sv, twentynm_hssi_common_pcs_pma_interface_rbc.sv, twentynm_hssi_common_pld_pcs_interface_rbc.sv, twentynm_hssi_fifo_rx_pcs_rbc.sv, twentynm_hssi_fifo_tx_pcs_rbc.sv, twentynm_hssi_gen3_rx_pcs_rbc.sv, twentynm_hssi_gen3_tx_pcs_rbc.sv, twentynm_hssi_krfec_rx_pcs_rbc.sv, twentynm_hssi_krfec_tx_pcs_rbc.sv, twentynm_hssi_pipe_gen1_2_rbc.sv, twentynm_hssi_pipe_gen3_rbc.sv, twentynm_hssi_pma_rx_dfe_rbc.sv, twentynm_hssi_pma_rx_odi_rbc.sv, twentynm_hssi_pma_rx_sd_rbc.sv, twentynm_hssi_pma_tx_buf_rbc.sv, twentynm_hssi_pma_tx_cgb_rbc.sv, twentynm_hssi_pma_tx_ser_rbc.sv, twentynm_hssi_rx_pcs_pma_interface_rbc.sv, twentynm_hssi_rx_pld_pcs_interface_rbc.sv, twentynm_hssi_tx_pcs_pma_interface_rbc.sv, twentynm_hssi_tx_pld_pcs_interface_rbc.sv, altera_xcvr_native_vi.sv, alt_xcvr_native_avmm_nf.sv
