// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:01 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rnwb16/XFt+qdowj1HDxd7VoxNR2xTm6NBM4T2M1VABANjWGLrVUa5N8jd4vfGUQ
oS/1vDIi6ZOhXjQUY3uHBVykkLa9GSLyJ+N+2xn4FLobItpH5ielhT+Uc2jv7HB5
ntVxqDWNgud9NlXOoPNSKzgCOHlp2Ud8SnHDVHidb9o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19808)
9udYvoxENkGXu5xErpxzx/HBCejO/vwbOknE7yMgmOoDKGICN3rVezAu5o7wwPDB
Ek63QqwJB7XsA99ZF3PRX2GdC+uTBS+XGqJ0a0RtErfCe2cou9LckW/uQwUMWYQa
wiMtMEDg07JiWcuSeQDVI/D3MDfHlb6RofpoqY0ehX5k6GxAiVu6A4RKPdk8xpQO
k3f4y0s9VoEXjNkPQKkzyK4czeSTQ8kmP7yMsOr1wArSagvtTWB3+tYUjPEuH6eL
Ugq7/7MVrhqGdmhMg5KwPrmMM1WWeb/pZDYFX9Sb+tXMQceVlYzwa1KFiiCTn5da
jOrmrf/KW1Qw1ZnpJqLUoh7QRYxxxtNO0lhL83oQRjiqalQcJAlUJx4t4kBU9iLA
qmEqsdNiAmdxsQqiKiSR1BE/GVy/jOE0hT9uECGjyQwFj8W8D4S2ncsD/UxcfeNH
TciOcoOtDWMYPI8gfSYWXTKkmIRgzxCKTmONU0i/5PpH4D9xXdKkr2+OtsKu7te1
77e/l8SxnwBetL14x4vxL8bYN0ZZtEoqbE+nKlxOqloF3Sizx37cZ6YdTsrfTSZB
/HftpWW2Lnl1UVMHfQGl2IrY27PlBOVYG4ymBKYcE1LNOwRNmZjaxTdUx0J2X1UV
a+B3t4mHUMgCvifjGMJQJY38z+jHsb+VR1XqM7c3kA0IfI+35jVNwF8yIWR1Mgol
XPy2VdKvvlGxGjs6SSG29OdR2I4l5Y/AJ2arBxwzy9OQU/WIzTKaWxpUpAqx9q1w
REMJVXrR9jJUSlfL9Tvj9NftBekpOn9uYmg22u/8G9g3cUr1LFHktXGOCCI9MS8a
sCbHQRtOfp45JTBy0F8S/WV9EVS+JmrW+DQnLNvvfTWn/x+5VRVQZw5pdfIX6eLj
m+FzS2DMUd0DiUS0qL/xqSHUWRXkOa6WAl8i7pmJ2lAC34KzLbwgQmLfoBHrWDnX
AJbvgEzFTu+m/mii6xLTqjXsVEX72rthKz3778UqKycXKAbyq/FiTcnRi83MTTRA
VWhbHpOw9yIIB+lEcucd5ovaxh9eyiev4Zq+/WIsjiTfiEgs8KWqKI9iINxyGqOF
zC/Oh0JoLjxh+xig23I0DFSpQyFW6cIYounrX+9+/5bUm/z72YiyhI7Q7GR3Nhnm
WVRLsS7YXHYWlUORe6ztaLYv54HyDNeeFWHt4wroTEeGUk5tuZbp8JqGFMYHoU4V
AAK/19rmPm9TBnPYdsB2LS1dG4R5Lp5br9wbyn9rwuzAH6UFV5pZYMFPwrRu2SuR
LTCNksiGBRCIAiCp18BdIdNfdhqp1/YM5EYh5s9PJhnk3vW17AnNp3kwpVPFNDGE
cazeOOL4xlvP5JVXjkUm9p1KKhlrrpPoDAzJDRBttUD4BsT3xVQTamYksF4FZXy3
L3aFhvPDiXC88rtg5rNXBIHAzE3LLoe48RfledF4wHzclrbPc6fzpxUhdRz9ABWX
dt+Limy0nq1HYuywnt0CAIltaSv5R/AzMMV+pSDOriuQRDDmgrZ1+h/wdQ4gsSAd
W45i+tJsZHhkZCgBLNf3LVgnm8NqChA8A3vhGXqkJ9yKyaQ+zPAyCapZoURwvYqk
5Z6zQm1NqT0ck/cbmR5wSFFqdulXAp21Z+v1H+WTlO+BS4xhqcTdZWS79TvG028Z
wacoHMTzaBwVMzGppG86Pazogfu/1ipdYWArMH//F+5WzKlmArQTjdGlpS4Hr7I8
0jmZM2cgCXp50WU+4uk8MU9eagnWi/7e9wnYUbbRFrqBLb0nGt00uuRDVUW3NRry
+uPEUG3okpP4qITw/sBVLmXh+P/iLSyyEUTw/O/Yw9qExSKhuXwtlAmYClrOF7DQ
vXwA7pyVOTpKoPkRXaKLaQXjEWy2tXytdd/T+RY+GXY0X/x4ilV87Uo/vDD6ls3F
lWGyqaTpamK1mnWM03NPXhQDLgYQ61c6GszAO16XObPKuJib0CxCO3kF6bxkPUoD
jR5X1uM5tbJt86MYl5wJmVrqEzQsIsDUIF8wKR+kxnC8HOBEI5xVLitGwGHwJLV3
cZP58q0tpC5oXMBsNfEk71Je8Z66AD9zHjvzKzSJ446MDm4uCtxNy9XNfeososCw
qTpJCaT2kCApxJ0zLFSKPAeFaSkSvg7lKKSmpn3LZUMlL6lWrwdrXAkS8vdXbydo
Zir/t+DcXSV2y2HFsGGgR89guchyYitZpcOCKBIZ5+912Yzh/K7loqZ8giY9ZaSz
xikC0QFFg6grXqmO2KxmihPGMS9bl9pWEJZCH/4W96zIEhOWGtM6zTGiqJKuUmiB
WjFKWKnHB31Fl2R+eAgg/J5aZgHLAAhlYx/ncGe3sa20tSiuWB5rM6oKpGNrGEoE
edOTJCRI7Ypo+ZPtU70cSDX1tXII84Qqs3t7HcAftgKaiiRs+qrSU2FStLAfJf8p
YNMcF+f7CrWwhPrBVBcnTJvHHucndiAJQOgYi73f0MxqyOOLipMbYWIie0dNnFUq
W2G/OITkv6gclPUi6E89I8THP91UlTtsnXjjxnNl8jIcDodtWdRWiuhnYSITksgS
k0pFjAtjvKXx0NsAXWV0+GevCgb2v75v5SZHFdZ+0Ks81IAmX9LA38f2r5LmnwW4
fV4l5juxzbJhG0ZMa6NWk92T8pzTvHt3TKUTK/fU9FGZ76C0XBNb01NjxdhMHP1s
MEJdN/1ugceU1H9Om+CULhRdoZQRnpB/0lnSDwPBJdSyDtEosRbTUMIfHLH02yFy
Ge7nUKXOyrAoEn7D7CAzgXqiJIs9a8hEoWTiuwMxNTgdrBJyx0iaospt6D85HqHW
poEmEiR+mSbhhMDintOXL8Kan1dhOFMEsD30eLcw+iEeift2YJ0mGmJysVrjglx1
1uwLqgcGCW8RSJXR4BMnrrKFZ3D3IjX1D+ogENQFrTGc3enPek/hCsxBrnH4U9Kd
vkXCcC4UXrCi1z1xWvbZKDSjuf6PWreXGuaymOppbiSLaMXrZe2GqR2P1NHYJl3s
BHW6ogtJ6gbCF90i9rYh6cOLYJPCjN9sv2QJ3CvQYDpQqGF7qn+RosW85DvxN7cF
1dlJRrKJfH2qXTqE5oHt3MUfjBFPeRU/SRkAHCuR8E4XeMIXJmw60k9vczPiUj3K
OT0M8YIK9RC4Y9YT2gpft3vYm5vMN6/ye9WqC7lGyrB+aa4EgOsY2dPALvqcfFTM
UtkjYwuztDiQmXfhuVq3HM8u7jNBJgwPMcg7E4M0vbQ7XoYbT592f+AgSs+UZwIS
1ayNoPpQY9qpkgmucSZZytBBtkQU4NbSMYn48lEtESkWVKl6mgMbr/QeLgiaswes
FkNMEyfHiCCv+w9N/ucJRbF37vWZmlik89b4toH08j+DpOGKvDzBNxZIxKi2PQaD
Ho4QFNf4mEp/UnSrrPKsyuhWPUAyLRqzeaFpFOODiLR22ni7/Wa4vqth4AkNGzZG
g4OuQICuUriemtxguaT9W8iD557CwfmWA/Ufpfssx2WD8xVdYn5BFSpEIhgP8Rex
z1Ks32TVfPNbx9k3+edsleOSXLTXkxlg5lk3WmDiYgv3mcCeMsawHOn74CKyyK8k
9r+07My8QFY37e6Gf5OlhqVIFFXKpzdYE6YTICw/qC0l8lMlMs3pdRTmCIYq7/SF
ykjw1h0be1UheeYEAx1xhojgCT/3eWbrGZhL4OtUo+Erc8HSp3JNYgwyGT8K9AeI
oHhJhSA2D1+ltV7d2u+346GyCf8MHTOz5VXdl2zTRnPtiPYgFn1WSv2yLeMg3iyr
Caqtd2AHEQIFwEfiptL9rLI9HDg/zOktZzR9W4JKWj23KXMV56FnAQ/gfXq/npjd
4uh9fKTkSBGuGIEkQ1XkABX/KsRbdgNHI86eySWUPw3JI+vjqECeztJTzHlvqGSt
tAIxGvr3dV2nmUyr0EEeh/4NnbSz+J08h8zOFe9LWwJTBtIi0cGrmsGBKE9CkxZH
SlPz8/AE0QMl6HDlCYegDYSEh10q7u4HQwzB6KwThJaqIjWVAHxt1qc0rVzrYUJO
aA9pglRaqKyoD46RXT2Gc4lDtCFxcup4DN8KQKjHcI4IXdC0Mzz2UlBkM9dv1EC0
S6qg9ft4YnfNZhV5cJl+yxVC23Ba6Gkz/sBNhlnSq5fq6VSGQUwg7PmpEbEp7jyx
LLNqmdwbe7t9kGhYvk7MBku/r1HXk/IAKJ5+DfcG8onG9EKAgdSkiPgTeIYjrtQo
5qBIBGLIWgg7WZ4a4hUrjqzb1GIt97iSUzySWbD4gvhbpdXdNGNdL2XnrK1gzbuJ
JqDPzwwYvAC/HdxmsHhb5bdox2jZ/4/P+zEVXVJOxrrTTDU3Uc8leWGsEkjph6DH
CQ0kyDZmveTfQ9DMK563wE5rxZRGqoaaxIAD4iH5rNePoitodh1p6DijkzuiuG1v
xx7tOo25HK2VjSDut0mxu9JjBY8lIDU4Z96UztF75/5r5YHXTYETzgHFFTS7fZjO
/SqC4KX14FAoQgiAuOUg0be3JTVNLPdZRQdHlkGoC5qsn2zV3uLrZYsRL2KRWBqV
TKlqoGDj6qUZz9fDKLESIA00JSsLrKmg3U4WQvDkRLXM/bc74OciPjC7ubWalrdm
QVoZd5CFLYLLZ4UBDtIUUdkTshO4l7A4RoAz+coBMrhMgMtJfhmVHWHYUU97xr6S
03z9aTOT03k/nXZP5aVVVHcuJroWW4VydsuCsLnYm6FIenk1MLwDqtNum1ZLLTbi
Nb/XAWTU/B/xmDkCuxKjxA1onfbRCPKxKoWtmjLpDch2z5swckpl3nIwjQUMHrqZ
vzBedpELqpvSqkLGU2AbvPiVFQ84kwCjLbLR7yR8uHiPa31jzbr5Owac/Y1k6O5V
+D9LjSnr6tUGNa+FAD/mTCdkobLe7jbDc1Vg5WmAT88cSV/K7PGMEH26OulRhBuW
QrNjmav8B9rtx0qObhZHiQ4OGCanXYg4U55mAk/Idlx1fQYydYB50NDGTP3MM09C
hVIFJKSzqrYi3xwazEaZbv6ijKJHZCG9D15fK0CSa4+uccGclf7AbkFkP15R/lHc
henJ+D7ZTceMEbhsfzohp7xRSh3GRnO5WWYw9xAu3zTf1eXyyfUIyyLG5sR5SZvH
3Vj4JKxDG8yxYzV03oQBItTX6d5wEsqvhDO+15Ntw+ko2IvYvB8r5rw55Ws+3VIk
UlLrmY3LGjPFuLAR2lbeVo6rkDjeF5OGPurbnHuvSkOjdlDiSgu2u75R4JDq2vzL
LC6u5yrOgwynsIXn7FqCDezLJpoZYhtWd0OFaupHu3AGEVZJwZr8rU7YfeFr8anS
P+udrv1JxVHu0nPfSTnooMEhLP9iQzxtnPEDCXhVFcMSHpiPvlOAjwQaEdShpq3h
4ke3SfoSt+cZrqW2qUyp0+b6wV2KcRBmtcDP76ofRjRg77JuhL1Rt4xb5mEJOdCc
ObfjsaZfDCMzU6LWPmm9eYtKPH9i7CqTNtsVHHhkkct5i12HMtql8sqrWkLb9pMj
KJDCienpOGfoWpgVjFfk8QlYODeb4sEJTVLM7X4avGt51hrfM4yfpLTrNmHzvnNn
Ulv2Dt8KmO2EV82WRrAsaPjtGGh2Wm4mc9OP2zvOCUYBeEid+f23d7fNX/ZYOe/7
dkG38NE9Hx76IKdmQ6rZWBmIJIrA/hrpz66j16IJgtogqHcldI8aAcrA0d9srZxO
3fBT42dmeEdmW2qAOykOnKwrXON5TjKOk+FI9PZAuOOrq3gP1du4KVBL7+wMOT/8
cl6Iprz/RIygwjqEMOn1iNGxtl4BostO/kN7yd2vBA3yRli4DtB8su2HsuDih23c
rbVK7YzOKK6vik1hn6jWh2OGRxFc/AhbqQswEr2Ghz2Oi6RAEPdvWH63gyRNpaoI
ic4eyP5JLprP+iMgFneCdOmben3PF808373Ti/sG3iy2mGtluQaoWMItXMPbIPOB
Rh9cIhgCgBlSqf257UjxHE+suUH7kmxU4QHEL5kudz6Gm+4UDk2W4YUso0qoy4z3
HEvQtYySu3YCD8VAxaKemRG2qw9FZHCPjFDBzCuePRdWsPROObxEgr6tbddYLlNw
TSf4qCfr41MR5cTZJVtP6305TJiXT6kPCgF667ukdo9YidKjbtIZITbIucBMxkmB
7dNz1+L9zDIYQRMxLk4aEZvF03wBLN1IFrV9wA8IYGi/JCxdH+v5sU+nLmAOgPxz
oUY/M+33HrPjb2dZK4CUqfaVgVgCLD7woTMSJBRCpI3wmAumTJw54bMOXileejfB
AARyZI3LTOZ5a/nudtOAUYMpNAeRn3bRkQ6e1jfuX3KlxqNdhO5lfHXJEd3K1XH1
y9i2aIYc2Int/mvhpSrhs598tXJ85OAruGrvE34nJoAhbAds1636VC41Tq94d0ZA
inD+3v15LY15nBKUfuji9vAlKo/UMcjfTQZ07Yqcf770XOtPlYaugtEI0qD63eD8
DrK5wQrAWy4BaSraFMNqn96XUJBnyeJ7+AtlqdaycNUx3fF1ZqQWfczgBXsZJ6vj
ylim3+0XeK0a9F1MJi9KdDbFvD7dLCzBF6NLDX2G4xgz8ze+PPyDlJwjZvDzLSYM
L7XvOlK6gaO4ammgslblaZyPixj5SE8lSRAV6s6FgD1hFjPwUrkikIob8yCnmb+g
ppypr8S6WMlcsLt820cD/Rkga0etJj0dW00bGBNT9SWmA6zb+Y5EhkvtCb2N/az0
0OH4AzYR/XDPCdQs3YNXuDSFIWKeSI6NZpiLE2MGwEZApValboJCY0qwkufMN/D9
t/VxWvBbWKsdiAjn3YwjQ7wCoIvIvocgjBRePmvTKfyyQhD999S1rd4BCg7cPXhj
Hr/lxDCLVyG5Shhkw4LPwx1Wyr0gpwF6KmpyfobgmtJYGmITe6YN9wTBdVmvDa7F
UJynGVZggq1SPJbA92+GAY3tJBDpWt4tAco4wYcB9RQ+INx8FiVI+/hfezbPH+rj
b9B1A8up9zXh/jNPQNcO26OqmOT4XNH+MA9aXD6y5rC0LWv25wfQcGaMR0/gkITV
cjsqoDi03nzsvYAGpUsNXOoanpUsMZHRP89mpUXkY22jwhB3gYTfSYDEcx6wRCEc
tvNlyqsQsbGv6aa3nPCR7fX1FJLBCf+moesrxKA1+r7WZAxHzJ2XvdItvx//msBh
N7Umzi6D3mv+eVZJMz1oQ7sv+Af5SGNsoJ8RxMGN0gGuYQe1dhNRfVQN1okSBgpl
1WGxLAFexpSp5SKz7Kt2hqEaKgTfzBA1rwC+/WoIzAePmCkJDtksPf4/v6tRl4yH
zypRvcYENt5eUOaf3Ay/DQnap6aHhYhAopkUAHY3vsVAHkiG+0k0Wuwu+7guXtKY
FpQW+nouyjkNeFPuxyVIGWisX9+3fSrLBUVQ4gBWuMZGefrwRONZJffQiGnv/2h8
urG8Qx+EO4DLZZvh+QOI+pMEXWdVwl+ObTRLjbJHiLHLzqjq9tdC/BWGPLAiK8kB
4ICUHN60i6QVJWHBmL2ByVhH75bOf4sIU7kfm67ZBHUSUl/kpM29dfmEnQe57Yly
fEG/BtE9ClZz3Z1DzCSPg2cmrqLsaUB9NqE5OcUL4+DITBM+iUMZWix6SS5EuWrU
Oqn+whYrBhLtoI36HvEp/rNZnrnVsgi4MUzG3QTQO9q2ARO21QWbeKqN2rBdoQem
wO0D2EySsvFyMGB1pEDF6TINxDktrZTRwEKQLjh7hk1/F94mU3faqzAgKucZ2kzn
uswkeXh+k+8Ov5/Cwf8/9augLfYzS2MbcLDmCAvArlXAiOBMBvhkhKvhSey6QpBR
GY2GBZoajUR9fjyGhgyjfzQTvMtLdzNN/s2VA9nSQW/Mm0YJu2ghQ5j1+er3ZVcF
a+N7+eFOQie7DcMf1Fk6h4Mn+DoRsX+kx028mfOHTbrLD0vzHzSxzEh09LnyrLBE
E8oDkBGRU1MOmecFwZf69btJkSyybIJ71QKk/fYUP5Uzy6IPPZSRxPDEPPZj7a5Y
blYmJ2JB0Iobxa2PTrh/Q8vG2u+f8A6ApCzU3PlK4/98DhMlhwPI66wq8VeiIeAv
mFLIlMgumb3jnlU13zbFlQzSNbUMEGoIRvI8+w6NGABifZXJfAT0aKMgewEp4s2T
nb1ct3Iw3kmNB38+7FH2rBWeq2AIY0nvlO8prYhXI5SVcxANqAjkmkisgb6ndfp9
esY7TXSEkUiOMUGKEk+cVEBv9UKfOYJ7uniqA0hnxl2L0pppyzsFN7kH3bz9RLnA
9WpA02ySPivVOx3ASpR1loD30jSIXcsCZj+RWBcJCzxYC7cwwiImd3Eha3dfGHmn
B+Sfpmb1pGkVHsXj/TqeiGMe/wse+lOjKJCve770o3ijGHbFrdYpmFbx6Z5KmMiH
Dt7PbzsbaSjuYG+lDuBpLcMkKAj0HSgXtD0rvqz+MBSYALa8SY5j4xIvDMjGAfUu
ViYqIPvuBdNRwzqxAhqIMZZfj/ftx/Nstmb9TXszzhbytyJ3eQqsUixBm6O+PlWg
cl5qjum9xc4nuFlvrJNqd01sNvTTLNCuiKP0VYWShrdWb2ghEgHcaogWbSrHJfHV
L5lfxq1W9j1HV5zV4D0kr2kHlZqzQEudnmfnFaFNj4ZT7ItM9+Up7SckOXGKiLjf
sO6SGecoLJNRNlW5pBsjxr8uFPVuENmp3GevdUZ13oO2Iym+nYlKJTP6GytAHKOm
Oxzoex5gg9c17bavrUq/eCXhqjDQk7R8xF0UrZoiTYj6yT7TysH74g8iloqUJLVH
Ath0jxgZJhzQT1lY+fSiVLmsPqpeXBCS8Cg4UPhxKPu9UugUKYw0crzW2AqKmHjz
80R9Gmym7ZcPSljbj78VlXgQHSkcELHUk3ArHx3R1xEZONMvg4jhip/7GcAtTTvZ
5yySHNsbwhSmB3Q0OP2V2m3aUtufYTFrqNkE0SoiiGOuUiaTQYh4SuVhRcRTFczU
L1OuaV/vItFYOGD0wIra+StQ6bCWBW69FRqM3HME52jN98Mozzu6unXi2/Zj7uMM
a8AYTuOSomdKOvACigAuE/3OTjTR/uhS8cf4hjXdN++PwqNUaKBJubudLqhQiJI2
Hn/ky+8PoUHMMjnE95+BI7zWPo+YegUBOZuh7tbTBsXbt9l9LbQW5Oe1rt7N6i5e
eirPAJksAdZoBCuevAEUjg21LU/pnQr1cbdiK+9KSZNpZcSz+eMHkIqmACCQW+/q
YRtC3tatGGwhvNvUPZ86AqIiwT2/H0TY7xpbYnkMJAUx8uftprrRcuv0yZI8OpRA
yUXk4LMHXxH2FPgIEbiJbIUz6t7ioHbNXq7zzw9Wb0KM4pSheb/r8yP5NPTo0NGb
Y2kvzzV1skvvLowzEXEGfsJrhHWo5OpwF042slc0fHmo9YOJ9RUn1mpQRCwZfKBh
w+fSC+50uxZJq+yGFFmv2wHSfgZiK/XTot6ian+E0UeKwcSkdLVxvsPNWPniijU7
aY9enfHIPZfYMy9YBUqFgPBTBuIsur3SwD2oUauWoOr8w/I7nVOJdfLPRBF9iFFC
E1v4NPiaYE/JW7LETVgumEZSmqXuTkgpu7157QRWtjAhadQTqgbUZlsHxhfnlh5w
SIohpnJUuMDgkZlxOtOnIfcjtMar5x1+iCI0wPCpORJ5FDeDUaRYA3KkiTU/YxBG
BZ66HZYXCczESGMiNf0Q7KX8NuUe6v9jA1ePxpKz0LxUbuz+ocSYJ51LAcshOg1w
/qsex3oZrqyBByXdjyeaXb+BWa+2UwbnxThtCFg5Q6DxzfPhHWYgs6lyG+qMl0HB
lLlrX0e7Rz8KBWQlMRhDEzwbLkU7wLBhH2qbTCL6xHbORZoE9VZqE5yjJ7p7YcLS
ahm2ga8MyhxuUgdjdCwX0RLgswODqIWX1+fuASAixggWt3ijXOfFDGukwEMtush/
lDMp8ehxiNZYuDiLbTsj9lrXolTR9kppetb7aXwkJK7wbA4P7Y1QpKC6RnjHNv9u
iLbRq6ky6h7Kfdg2sD5UDxTs3nIArhkZMouRCgjbYxFnO/kH3JjNpJ6a0xmbyOJD
B2yggFxdaf8MLbW93CjwuRLfyDGgstqbx4dJR4tiDvolAavoVyADhGxlXI8BHq5d
BkkXpgP5rnOgz6El7v43lKszw9z3BePX0QI55rF9ohXovC5F7GKFJGw12r2aylsl
PpfsZEaAaYFqcjl9GAwEGGb2kLQIuw5AhQ5JjY02eCq5mZGZjyaUEJkFHMdFwkL7
5q1yWmPaxdz/uzQD9QQtWmUtnEsj4rvRmWTJ1PV1ttuxxnJ7zVTOvzYPNZUF1luM
It6xGsvm/MgrJylz2iwEpBOGLiUgGkkX3bmN5c+BGBCFyUrPhYrGmDAU7kAOIfub
wY4qDL4cQMfkdLbkhwz0LvqoqITJKWsDuCnIfV6+hOynE4aH3OX94vMgIRUGL7Fu
h7+7x38019JxIGVuuryIQ5aghzEs5l/f7o6Hlk0W1ctUecc8yh11aOAYFjTHUeeZ
NeDo88Q9EJ78Pbc8s9HF8m7YOVJRRNmvmFh5NqmAdt9w/hY0xYmXMfolCMd6v4k0
z+fB6Q9JJR8gAnyaU1JqZ8y7TGU9txht0WNAAmsAwxC5moXWF6q5kDg7G6ak2VPL
5OJ5CAz2B9Imkelbfr8Ej0hNfmaCDEgrTmB1BpE6S2XAorrKmm2qfDJzB56uRZZT
3Q4IMRJM52u9pfECySABcjHKIlHVa9UsQmkxcfc4ksVN7gZGRZ3cNzckwR9kHYee
gLwQL2LVfz8ch1PWWt1Fha8iYB+ccKhuRVQoYuOYN9zjf+cCZnTGRPPaqRO7QsP0
MY095gbV4u2i6zPFv5rZW9HcDI+aByumRqHdVCuzzrHcDwqTpVtU5FCcHL4VzZ/E
LbXv1OAJUZY2TZ/NnvyTpQNgq87EMIsPXYr/VtoqG+T3hv/MYEdjbgaJ54waZCuI
qzJgQrCvBlbyRN7fSTmQHB2+0F4RerR6YJyTeCw0DpW6b3RnaAYQtzXTjMXXefp9
piwBT+ZLuRHXw1KIqcoUMLOy5ICrTJ+s9SE0jAXzNmGmHlcgG+bgyz6rI7j+gdBP
YY2LZjHtYUhWpzrGJRvy+Wb+ULmS3evcEbOkA2qaiyyOHo6aJKMy9EwmWZ4JQxom
KY7ig+m3Rl0pafvoX4FLUecuMLdd7OBCDEpUKtGBKiYCryaulpuSFaYXezz9vX9D
jXv8Tlb5UlkHyfJ72WPdFEVCo385yyQuxVT4XiGBeG62m43DWm8/SgTMMNw7aW+w
aslppmHSum5o9zK5ZG1vtV/tlb9zuoAH8ANa2apopJRtpZmq13r1eUUdRRMoZ70b
d4wAmqrKJleBq3ZSHqk0eBGbvFhHtbqC1MBQ4kxbl1sh0HzYYM25LN/s0hjM7grX
091SIxlY1KrJsSayPckxp3G6+7sAb3PAvLkxJ0ZATHa/qGaj10H8CGl5P0qBWNER
mwWQP5ciFv8fNPktxaXVeXK9zb+CemMBkb+IzutYoh2zv6bpOxTPFJQrsfxuHH3Q
6i9LqU9x3JM8h5vV4TRjHDbS/qjx5WuuqcOc8et1rYk9Af5MyKnts/3lTEs+xZ6N
CNR4d6evG35x2Akvq27xTN8LLoOk8+oX//OPdAMjwlVMPrzoNW89FmOSd7I8BBUa
2bFGlRy+MMxFGfKhnfX+b8TvqLEbpMxe2f0IclewslBWYW/XhHGK7oF7TkUzGFZc
N2I6s/X0eL/2ZrR3KklKtJOciHA2zjVSO7E/za0/bTGNFJnjt8f5GIcasKWbHarH
8lN01UffZyihzycWslZHYUag4wRuwMfOz83pLMmvQE28vkOPOrBm5Mz+Ua74D8rI
ta8Kjq1HNLnAnOvmV62QyRxibrH/HDA0p+SgLqOjyK9IFQ+r2U+y3w+1kQsLCWFL
hkLgtTSKXAo01hoSczQNuuQqPj3rY4rRonsZKFEP2oUra4aMJv5d8yVBpwVk6Kef
EqDk159F46+o0ZHV7U3bWxFpatySmI2LFGzSI2VU4Y5fJmPgiZwQ2bVEygvwEboP
KfFfXytHaFqadVaSDIAFN4ZEuPpy5hSYSaMKYlJW49PqOCCNAv67zcgAYm76/Bu5
ISpfZG1F56RDr1oSra4nt1jt4Ak8gLI2NmwZLjkQv2ucQ9r4mblpEVS04tVfzMCl
jKLmq+n7fkz7JiGLrErSnRHCNgz0pT/RQ0rIfps71ewvjREAuiMMoLPDaRqBflO0
R78f3oZkK5egrO/LXXVKLNOeAax2Rk/a0wsoMJ74ZKKgcqTytHXk7rGLTijdsFZz
bwzGjsF85QWi/KFe24aZbT24YB8kORDv7WcczkZeqtCk02IX6PTQ9KbzWiG3pi3S
EdOUwELaFJRMvrerFI46PgzBQ6mZqwBvFgi1F/g2wtlEiAari7wxcg91L1ToVrYh
24reWj9Wnu+Jf4Ru42GMOwMb6SoL3a31AcY+zokVUtJrWxN6RjvQlOmst3y4LHUt
On4gt6imvId35N5DHBoEKWI3x8TzG+mR3nQb4utArrNfXEwL02MPtLj8iDYe4tpB
08R5ptujDxL63PKVF0Ep+qZQi0hZE3MUdpF7D/ZKVIbF9UYNep0d8RSU0SoMohHR
q5vejL8iM0JZPll9ytDsubTNGlnbZ2qAdYPGNznDORIWaoiFnD00DWnaO76ZwXRW
ZJIaU/iAjxOCBEWVJz9A/2EYX5EklGeHwZHgaamzsbZAkrNMQpfcZr4Kdd0iDkW/
5EbPumgevPaVQ4qNF1yuDs1P/zDEKVOQ0R1O1VpHAHwMRdxFU+5oBlNQEbTbwrLS
o5AD86YWr56KQRwVh2YP840IfbOW5Swn2eFwO9hH7WSnwQtdPHTke6nW8AUTnkeN
IGYrkTI43KC9jqp6wxikxZvVapCgKnSymm+AmjL5JoXVngjpytwJsBdENW7aO9WL
empuIxlaEgCscwZ814a0ja9Gr2wSQTMPVCGl1NAtF4ahoygHXtccC9zyQGIB5xvj
8Gr5kmrCvgj7SK9RkHfRZe6q6yqfdcNcT/Xc4kev4GvaZOC8Hrb8KIR28Z9Ji1J2
vXv0EI0cjdUmggK5ozJ1MlQjmbYOhBaKIH03u7SjrdMRfKfzbWXUpcWoKj80RkGS
/2ocMatpxokcIflxkUCiy5hOunzRyzx1GTXkBdnhM5kV1+Zwy5LAi/wAQKxUqiFG
0fxRlm+8rW1IvZ6ubsV5GC2cuLhOU7D5MsP0c9OVIiruYBiKLLSadVQ0qVXAswj1
OM2Wj9cHWtazCa+wsF/6wTlZDdao+a9jkIuOETpG2Q1RxROXVjpnghs5pjNqj9TB
9uXXHmCv/C85lMUvlppjmVl2yHO78JLn0qrEXL06csZjE3NWw9bJRq7VQ5VyrxNv
sWIB6RIisq16pd2EWxmh+8B4LyOAVb/jaqrjKi5gY+5zE8TwQY9gYT4jliwQbU4U
DzQZzJB5MNGTWCA7tlWl+vX6S2MU+9k4Mo2dBIhhFvfqiThtlsbOWNkWU4p1s5Q8
6CvZMX0AqbujQDxw3LqgsSWZmeclmVCJzSPpRmmvSbXufSOpD/e3VlpT8l7PRNOT
aNuNMWX8oKJUSMLUz1CS5tEveLIm/HiTIlJk+onzq2QYu8AtSjemrjh3nRgvfXhE
WquMEv8wXajI9KR/Mk0GGqaraoRz8LnxJ9u0rbljPye+KQ5e5EAHmT6T51u0dbV+
fvJnkKWOhiVLzqJJaO3eCi9a4IUTaANi2gF7R/9NxQ3RA4oROhUu46E+XyFRZuOC
zvyg3hET2J3A6xpDm2O0L+RmPB1VCpZM/HfeIUu3ejTBgnq6aMUUHNY+wSWZeQje
DFK5tGwWD0AG1xYLlWpEoXYOt/RMHPu9jeGpznQJongXur7XbTNxc6I7uNieEnSh
PdV2Bxyxj6basMiCOugDm5Cw0a7b8Q5xUiqihlIES+3DKVBON1NmCARc5wdBTpOG
OWSWnOAowXfzXMjGyAeUavrHyvlRev3omwcfQvcSAzpCP8OEgKBDGco01KpfYUQl
7oE14JZJFbTLTUX+/V8H4NQk884JEBkjAvVmHBrqvh5eeQWCC7DqSlx9rVmA9MBj
nmc42sPebIfvY2GvL7MFNlr07Kj1m5nfadOdshYqL/BhtxwWV5+YY6jlqH5uExPc
0v8T2Aen7w/hxmtYf2B/UoDFBQchE2AFk5RK4cpfCzRg1+0n1+AcUF33GBb+asPm
QOLAlG6m5jSO4koert1HPxYJszv8tXegf0yDCvA7DwzqxrSWerLSpKUeIfu2t04/
HTZycvxYLbo4Ta5jul6bphi3snACl+N4AvgABnv5BABJD2kHhawJfx6m62/qPLZB
vVFVY8JUlGosz6QldjIvvuKlDAjyIBgYtovwrUPDoB9k5NJQgPuYUZH4jy7mnqNn
MnYjT2aupLVDKSlTiLgTzpHhrHoSfQyxyIcwgp5AavNdkjtu9W3o4zDoo3pK7flL
PQy0Spiu6dDIhm7actPyApKc+zrwOCL3c8/kLFT+u+/b2pxl3xnWU8p67xCRY6Xa
dzHSDtpm0yEb1/k6h2od0NjR55rY8qTZtOT3PEPIypzBNAW4KAGlq/dx+psyRDWL
87SJbU2o/tw20qEVRvvjCYZrHvfgGmf4JkhyrZYXPhhzdnaHeHRvElaxlXjcJ+4c
4koTZ2zqZO04waAzFxQt+RaGXtymgKPAjS1mOuTn56kqGqDSpAaJnmX0hr8YF9OY
WOtx/EYNyx1cqMs1BtXUU4m2V7d289+X+nrWa/XB39y02pmuVsX0mlnW7/8nR1X+
Mk0ofNtxrhh6h6an3teLija/R2z/giIrE14pILkNDOhVRAvq+EfBFtb4wOXLfuvJ
S7bu1rywA9v+/N+ZjkBlEtdBXn4hsnfJieeadFazVaeJtY9/Odklofl55lWeX4TK
KUWyFs41gywSCU/QezrQ7p8SnW/CpJ+6AdPubD9mSWoudq2+COHToFeykLwoZL6l
c5eDROpHowSHWAWORbyEJabEsHQIGl8nNyPJQw7yuZQpHf5dx0dE78wvre+Ko8XE
YARxfIh8BqsorUQ1pV/LfPCFm5MQaSSX3gX39JkZQaoybk8TQAra8jnIvUgmPIxR
x5wqAmAEtEOZ3OgmcP02KvQJ/Inpz/Fcw//8ILa+3Kg20GQXrMfm94aCu3YrfGv/
cujP1XOIZ/DSZsoFbo8G0SnQFSwGhZ29TTt5uagx+qYVwXAg8cQ2Nk2cMgu+0eO8
39aTpdKUSv248fsT9llxTJxRpiWFj/znKtsI9CkoDruErRkowVCusw+enJl2TNGG
ZLBJkBlUg+DV41rmnWoaccNqTYv7XwaZO/mTdKioU9f4IIZbDjDhgKmo5wfbOzis
fzZNalqi80oakloyPJ9xJZ2a80bWuFBdK1w2rj5jb+YBvubVjjjmizRxTyEwyuJ/
okA/JuziqgHeEZMRhdnJ8mArN/ByOz8XjY5vJGvLVHBHuoxPFsO3K8npfFrerqLM
fsW/cYRc0LApvRUOOHpggtZIQZe0huuJZnqkDc+QCKbuZDTCAQgqNP3C6QJtR0D1
efVfLX537cuE+6OjMYa/0brduGFMSnkZDcS3HqsJxt1SuL5P6YfX8Ead1iPZPXMJ
irk2O939XAmkNH0klrqraO1G8GhINBd1+T8GM122QOtq1YtZyb3p0WRAjm01T9Ym
GA0M5I2OJ4BwAh7shrzaW/9UeRtRAzKKR68D8sH/GqDmKj+xd5ajSSxOW8JPqDUP
w2JEBwCLM7fa6omhZSqFdIDeCV/fKPi5JJCdUfLjOcBD18iK0/uemRBUStmZ/5jm
vKk2Xemwi4pf1MdyQL+PQY2yCj+KKOGRYj3LtEkWi85S926jnIjznVaSfxQkGaT2
txflLoFcckQo4N1wp2FYHra7EeSU1vwMIqbyT4Aa9byZSaBfn5EggN1mte7cUfNt
y/2xcJkz28ZH8f4fIJKPA9RpA/CUehXhse6Tu1hr/Vnnr32j0ALJzpIYjZ5BQFa4
IDGpfYPrYlw3OxjywQWBkYuCqshjNUAf5lAwOO/6994UiJK/oLJpgB4CgGTDCjKo
ziiIVW7S4YmHFKuV9oCvqFePMnXzTIRre3r1KzchuzzJNxt6bS33u4VUsIStZpl1
YXcgYeGFQ8oRglXRSIamjyqsYfRCMvgquhWFqgl8CFS2YPfA/dLRii4BDQnmhg6s
FXrEXmMgMi1A8hcqXtVMZO2h+gY+axXmwTqt17+LE1Lr9X2OaO2MwstHOi5UVlWq
p+0FV1Sli9VbQWEYkIqP1cYE17VKJvOxKFMqzzOGWBImk3c2wo9shEDfopRTWOno
EKiKUDi6S1N5jj6yXZdX5hu6U9ztEpC8N9jy9Knkaz1xGOESdPc7tetnVcBa2eqH
djuLL8ZQQ7YlQiV9ZR8Emqyut7Nh80TnND62iEBkyyl3ir6jWeTOh8bKv29Qs+sk
ZZHvWdkECufOvsSwAwkl9ukOh6TeViHiPwureMjS2lFO1uwKvSf9pATpKiHDvFFg
cjLz6iwixBgdhXO8SXyJvEK0B4YFAfvqkUkYVcJIOuIpx7UJ2WiYCyfyobjac2BQ
xIxvLKynhG8Wk8JdxG9f74OfilFZJ/saWeLg1LGowvmo13MobCqv+ErfMHI29JDb
90onAIDRb2HQxAWM02YezxWNgJLJTcLEkmv9RuXM/jIIDcipPm19yMJx7zsLzov0
zbrnZYTDofaKZq+anCo6n1W2SR0tVhKS7zkPhDWB3Sa5JZ4fdzDnWI5Z7WmOYjzf
010RmyLXx3MEE3PoBE4cWogJfW8m33AjuAVHFNVS95263mTkvDkdQBZV3Z867F+q
yoABB8OYpGU4FKnejqb6FSVjiQEpjZPwZCqme6KFhJxO3hOWQwCtevtwuk1nMHpr
lBB8VTX8rakuI9SWFAfTf++MUISESB8OkYy7PlZp3o7iqXqr8wJvKAYvbVg2ow78
Nwfjh4MDmN1BoqO1m7ees/DDu19Z/oI/qca099oYOmg4DdLAX4qJre1L5IXvuqCK
F0yFK3huGbhbztPnBycoLCTAErTvjcQxQngGCw50HQEscrgRf9jCNi6FkomABYLd
AqVBLnLLGx7wgq3Y5OkSdyFXtQ3fFc+1+qSeENI4Ta2zrNMXAwqF97qANvYgSOSB
GeHOhtJWivK/NFX9JiwqkMMm3LI00uU24z3wnGPL14SQNNAWeSlp2VXI8xyp4DRi
W9zkR7lWmz+8u5w02De4IEGkhz5bwyL892JgKrQkW+QnBuLkiiQdWooo6u9CDx83
ZPHGeMXUxVXNCKpFaHGWvj6O41rLSO6NKmh793OKNAGkDSaK53Vl45VHi2BO84dQ
3o8DT1Vx2VcV6hcpQJA5FxZhnRX8zlszkY54yWFzc2j91Iu2BrlvjS2+D7vSJ5MY
ueOgVl18LZSywyot8hbw/OGsDy5EX1Mak3S3DR2LdHxeF4ySJbWN+N3lVgVbzGXW
pQlwVC8hlUQQzhfJa4G4ln6X1nIfsk6BgECN/Hdc1f1frWF3uDd2rkSlA5ZXzB3n
ZFyIbRVhoEEvxYhiUWMPgA1tXGcXo80ZtXG228hXzJJ0zlHxwHhVz4j6DEYCahMI
rSuaYKcOK268Yw1N9Tc4wLzPb/1QMFFg9kbqAn0Fs/g0nHoCKx3lZOn1N7kRMqmU
yN5KsQ+/No7667JgtMxcZDvRltE1btDR104ucRWTH1Fc3wD9vyp3UK2Zvw8on6zn
UJw1oLhGxfOArfDQGO3LfI1wdv6d6XjNIXo8tn9Mej+aELMghDdZIbGJF8TVFoTQ
6t4TPU4/wLf/7Yzxi8oZEHhfcKhGt2JXITRZMayLgXMaC2aX1XBdh1q+aHIeWen4
LYo831lnXW/vD3nlSmvdMTXs/iQNz6XJJn1OK0tdD/rkOOTUYH4xT7MSmp8B4n6N
RNrxYROmBowbbo/J0dkbEy6Bkuh8EjyrrdbhjEneBrlCYIOTGvJT8IWK8o9zjpsR
6BU7xQKsubC5aSlq6BFBI+y2F81e+GLqCOLZAIPvKQyXKZ+QaUZ5ga0zcombqHv7
Und0IXwrhcpGt0HbK49HTTi3Iqu/VGopnZJvkbHpbSS3j3O+GD6p34M9M3zMBvP4
1WXyhQdKJ55KydsrfZ4CD4EjdBQoOfx44LZvqziMMFrhtRpTPj2Zle9VLLnOv5V/
zof3PERFynJUd47keDw15VJv1bkAWC2FxZyKaiZhIKAhHGo1YyhKzB1eYnWTPXCY
Om4AnPLw74xdLUid7moA6UV5ZcmbfYCaRtYJv0FB6vAOmH6Iu59gw1Ww9G6lTgVG
K2I/7OKIKz7NY7/ZHC9k+Qnnjlv+KYvi0jntU67MSEzzh2p17P5jwlyfCF19TRQx
KfwNrwpkaQad7fNzD9mISMsPbKBJ2m15tH9W+tq7Csc0ok1NdI0tUU5Bs4DBXkj5
rn5DiUjFUftpAV6/pTOPpOGotUIz+A6DAIXDBuyYRjrUt592YNQQTI+bX/1ZXEKd
o4gJcq5dW9n7mkAD72RKXCvjPaEeMnY6/dSKIjcn+h+xwKvn3Gu158v+iLhZhDeH
/5w2FkPXW1CvXkc8tdb2B4IjTR2AWfjDFn82YRObbzGQKzCmHNbxnJ2Kn3UhBWCS
a4MtTH46jQaOjjFuRghnv984LG5mwR+zCfArhLc0TFLTfZNXHFQMXU2Usvd5dyir
lqYIXhczmipZVym9PRmhxGDMktsHM+LJM8F15vshceO8heEmSDQkAiNJ7FYhb791
6GNyH6UANIBfeL5klfY6UEY7GoGMWAmQguzv36iFY0hEKQUUGFgqXJphQp9yTZnD
Ym9GxGqsdTJv8ONLZKaEh6kKIw7sZeSPTh0UxmkEEUv2x9k/FGgjaq421QMOmsO/
fF8frA7nQyfo5yxeD0q+RMVZuJJWyxxyXuxRVT9BzNYRUKZs3fFf3VpZB18osyCa
jfS9hQlDWcYZ7iweIuO532uHnqwOpR3fgDIiXhQ6Pu06QetbPZzQ7Q++kGKkxd2T
k2Jj9QTb4r8gKlXZ1i6OfZ28JOFBxABtCBTSbC9H5aefDIwyW5HjL7YAi8sQtmQ0
OM3L/Qvp5GvmHkbZG24HZCnwyHk5KsRduHZzRCIH8yek6vun8y86kGTzXmvYcFI8
e2OzWlSS3hXj7DvVUmsPcbTsOm4FMoVc13QePnGOSavF0+GiDcmlZwKk79AGEv55
vayVmlySscXGkEJvHfuyAoGCkg090yA+/zkJlvq8+CkqDA6sHL8/zR8RXQdqdX7M
ByAjMAAyQe7sH9QULOnIPpwaQuZbgaj3iZQMu0cCXd/syIXGdKoaNzUX2gFls5XI
N+h9imPm0d3Ef2JTh27PEHyUJeHA0RE/T4u214I1I3++XvGUg2ugla0Uwpa/GqiR
YJIW98cxMGnnMEtnOBpRLC3+00zkEPWT4G7KuuODOIdkN0wKFDc/j5dou2m22bM0
p/gr9JPSAUd1JIOaSIHWbNRIsQCiqRjTi+nu+W96PlqBl/354RIEJgkHYQOQjUxR
XYDy6Jqcs97tJCIxcSysZSLu8SNNTiVaZW0nvgAbJ1lbvRoOAU9auPTqUvqr/Wnr
zKQSGBlrNOmmnOzmM5QU9iZP7iOgc/ADUxKYqeD/Lfqqbgv5zUjGdCTYrYNy/VDh
ut5CnBaGC2LKhtD1Qy2O/7mQwf8rK3oMdu6NKipWjNGidBorcDEbHPtW3c3woaFa
xBVsHtCpRun/et981eCqbJLlvDozjG5FO4rcnCh0RAuLSeTMx24b0ZjbEFJSaTzQ
wjq2kUbXb0icpmUVoJH3r87SmJCFaRM40l0tUX4V3GHzgSlGmtlzIa9wE91JfZtk
8uHAX2O7sVW0EB66Oqpd46amucNM0Yzks5KXvIb1+2uvNOk2e9TExyo6Ahe/tuK7
9fPDpHkt1eqRAMeyegiBkdcinNwkOYK2fyQRcHcEtMG4mRjCuT9kZBkBMULjmYWP
jVoiYQmJ4FraC/ujrkMgbmi9Z8g/0nwl+WJB6VI6gaDlKZlE9OTdPsAcDHx6kp07
VVTYHLBA8AY5pnTydz/Lg9rmYJ/Ofmwqrjkh+d5wINjDKUxoAxV1NkA/zfELC7eD
NVXYJOm+16cLRMC8OkG8z8MzPTkf3n5CA+gXVhnpuQsbCrxhc8JG+CpDkjzgc/Uc
bl+cCIdnMlE10O7MXxF/1ri9JyS+OCBqcIuJJdacD0SzCOOi729DtVj/LDgOQFQg
+uS+LLOKDZJLHrAOzFnbP5rF4qztu2/Sk2GnojspKLFU5gjtcIksBq+p8gFSVBqy
QZ3zCQck15K64ub1zogZa+TtWoFYj25K4ucpOeMkXGXtACezs8+uab1+M1utSK8R
OVOi6Q5Rzb0B6UIZ2LRAFk3WnEaqvyE4TiEs5zSxgCAowBpvDIxkSvahXfn+Byr0
h1AyUk8kOy+QvGX7pzdS/Mwmiz1F2FCUTOkInLzLdWAMKryiUi5ALp8yPdKI2DaB
1vautdSSmerhHnUCS9yhIxxpPxGpfkvY50FLa9vG13tYNt92r4MiAy556oHbdL55
HRq82yHzG5rt+j0/nxN6mKzsbTnCn4ezbQBwfOqrrN3zgLgrrGVvreD+E5XRZ/5B
zSevEBeYeERaSMC34gBVLF0RC/lR0XZMSgoZoNKHagpkqF4zcYz0NJblwlOlqrhV
hTGzXkh1DhDLIxkk+U4WEPxY46fLiaTzmfO2me5NQ+sIVQ98u/3qgiBz+rTCj9Jm
2f9sz4dC0bYNQh4CO5T9IvB+XSR2kC9Wp9J5wpRqdA7PLkUpgodcuVGdYEAikRIX
cxRtlRjjNEu9tVZsqsfZKGN2f9Skgg/w4mMqbUkdj9kvdJ/h07SfGNpz1fM/1+9f
GCCN9cq7YXl6nMalA+fmrh3A1NgCcMRbUFBWiaMqkZA51a7TJ04m2wowTWg+3S4m
BCENORGqVvpFuh5FJLBYz5cLvqPzkSi/DWXrOH/u35cc7eBfXIWtXApww5BPU26r
6DJ5OufiBC4rvZgabLhlkhZUcHGAV2x+PoGsTfyMKrzFGGJ5Yqbgem/c3SH8HF7/
SmRoBXed3yR84tbeuc/oPPqgUMyVd1c6Yodu/qnlzVJl1rvknekGf3N/nQTqg7i7
bxyoFFVKAa9Z8OU3an9zVEBR1lvPEQOPEjSAkRSWkHSM/qDoW7MUxEIQzwR4iICW
ezeXp8uR6KPXD+43aqRLwEMqncy98ZLraE7bJXnc3Vw6a8Oma1ITWXkE9Fv+45jH
u/n8bcF6kkCJdeyFv+q5qf6BSq0lsmvcTg+MSNgcM+Q6K1ztmlkn9JyhlWlkepx+
bns5sXSaF+4QvyRwuT1oY95IKtymZvAus1uo9Fv14CdlvxI9/wbX0YZ7Q/UTUAb/
e5DdIKRLdPSXn9KqgMptsuvgVpmAAClSe2W5eXAAR0dIpjkXHXqOAWHAdxA/o19m
SXLa5WGP2S6iLuboPUVof7XPVkwUUUZxiPMSRZbTKE91I1BSaL9BMnmr84/Xwp7a
9iLghppyGTW3Pny84SGXOg7sCjGIpGeh7w7QZTz0UhCKwy8qw4+g1TC+FH9TdIJB
MLuW2IweskQFviF/htyq5ggtS4+1O1Xz83+e/TSAQGIk/HMbTyPXJQYLvg5jcxlT
SIRXtXxfI7JciMJwKdwqvJBi97RSgxzPYU0RpuDbqKO81ga863mviymgm4IOSwKM
0TGXiOLUI+dMTNas/rua0C1kQNGYP1uDQJ5k80IF7U9XZ2gLvv7rGQtG1O1rVi6F
87sQDMfqRfz91ymQWu7pYIxIE2Xg0bPOo2Pl6lT1Vb0moo6NU0kn6eIurXd3ZJJO
tTMOGYdq2LW1dliNZs+TkiYPH9aXDpXR78rmTdkAYXy/nMD9qIMDiZUmrGBqPrCY
ASqtWRcL64PH7o2wqxX4iXL9FJpDn2Jsj1lkr1Fr2yu0xcf8KfBG9HDRVWPPaChr
oE12GZk8bM6ZeQVwnlDCnRf/ndcRERX73sTDwdXZkZQmRYD90C1RmZT+iW7OXXDx
XAiRA1jvN2Ox5M+wwrmRQJ61zEtUBbto+V3VX00MlHaelpe5CFYFnrklSZegaAo/
fGT8LwJ5/nOsqqnz5RFMlfefIEk3izFO6br+FXfH3ydhSVTkxybpVmGDMyrWxzgg
eL/FfiKQ76zZSAWc7QoQBfpeUG01pOXLbBCDwzay8Tp1Je/DEfT5ctDpV+G4MLSo
/Oa9iyFudTGebnIsxgJLKHdr0W4c9f+R+whWywSoksPomrNQYBCIky9KaeYOWqLy
2vFG51ovf5MtxKEFUQN3fb4ih5UTcGqQzxrSSVGILUKNpKnQv8iw0leo4WYTsoaE
m9icH2PHzWNvlZVFeH941lUtj7Ky52VmyjAEbGC/WBXsjUomHIcWXLgobszpu2bk
6qNjWHN37NhPhFkYaBpEi4T9lzRFLjypiEgwBir3sBn0Z7be49Q2itCZOT56QLMd
DBlh4B/l3GzMrpBICl7ABcMJbWiUiISyal7nOntcLa0P0r5fWRqUjnydAGEUVx5V
4m9jFsSy9GKImTyUgkb384M+3J+DKe9/M9amh5+ig6CweQ8qvqrcyerPua5i3kF5
09iBHk69vPk899jDEXF7PqRwVeY1uPvq4QAER41G3hCXEiVlFyAt3U0LpV33wCbJ
Me9h9KUfeWZd7v/FIOEbm/KAgdbyJI/kmPDMCitNuEi3N3cOMjQQml4om03t+Ilx
tFyTfrpFApwbgDU+g/8q+pxry7UYzl4xzjkbkd0AgIwiDhTR0M61CKtVHsrVyqBa
wkeSUJeRUvAVP9V81OQI+VhElUSWIFSiHA+hOOlw9AcwjezZZLLF/yetAReC6URJ
2/SUSmXG83MeqYh/L94tmau6rH0cgfwbfXiGf9vHTg4TT5cXc8CMZNMV2i3OgNb2
dEefkshKY/bLWwxJ/I68+dvT/0KEG+a1omLJZxxPYdc39UIYxl4otX0N3CZQzybq
2RhA1wR+xfQgyeiBA6JuuBFCbCflfJFrVxU1u7uIhkO+oCla5zjVwiJwU/n4MzlL
H5K3Grb+P3dY99JiEzkCSsNeh0ohNm29IOOvbVFAIeRV9Z9UIanTSzjAQz+nJ9LZ
Vrc7qoDYaSnmayBBE2NBROYSjFGbHgFKK+1OG1FJG1YfBkCWX2Vh1+99TUIPv1D0
RVCy/0hdW82h4JdrnPT1TL0fpI574ohBPfmJtaNwR7sBQ2IPBTAZ8Bx9cO3gZmDn
PK6RGyq3yB0qDMaqApksFS7jid4JAhdMmS7b28krwqWyyC0yHr9OCLZLWg3GECtl
IEwy0mO3Sj8q6MA89iA3icexqUH6l6Q3/LDhpwDRjAkPLsQhhVMuK6jFIHJgHYEB
ODYhUr45+lFqan2ppraLKhkb8E7jyPgt5Ie8Uxt+0lrY0UM09uoCBpaPzCUYk+gc
E2kqqJkf7zdMKe+Lgv/QEsCbqDUTQP47cuacCUq0BsDwHvhyroJjVwvlvLu1+T5o
udQL/F41/+QaQJZ63JsN+wjUbYaA9F4eEuFFsXCZmlLbTnZs7DuoASWrnqrfrJC1
SJJe1udexlHYsYIrCohxQlRDCBBbEqDU1W4aS6pxKc0nLFo+ELVhVpk8/jjhNt/F
B4mGi6hlDifzvvS3XHX1JNE+jCiiIyT6Hc3se5CKLRViB/NeYFo6GvxGPLcabQdR
nKlmkvGDM96zxRcxcprsIngyQG1JzvR/scnizFSAASGW3FYAk/NsOqeTrtpfKMZO
Qe1yTKBCvKe5j2nD59sVQv60jgCKOdB9vvME9UeudBXwZpAuxu+g0BZU0mXoY5tv
oz0fm5jWT+vsExt5f+KvoOIdGSG6dJihXYiJYOJmg7AlddFFeSI4s9vsUQGu0ATd
6TNul0YuU/5FuyhjJ9c/h4TujIYaztsl/uUcOebnW6AoH80CDgDvkkR3V90dBpR5
yqXuBjZPHg9LFq2I72MeHrBRm8ag9oWM34nf3978WxO5PK4qyEnBfBdxs2jOOK2m
DAO1gvbcWPvD4VNPRJxjkEPtUg4X0ToDz9TA5kAL7Kjv9vzZd/jmEBkJacdWaKN9
ud+v3wjuQ4iIw0C5fmVE0qEq5kbbVdFgCM2l40dM0BYOSLBnlcZ0SgbYtYH5zOcE
306JFFlPn4iSZK6/12L5+OxGJSApkdqdzA/RWrOOtfXbjIhLYFJ3VZItLbvbD5WA
67TXtSwDIXU2FBbNvgorVRvADbkTMoFLPpdwvhj9ovmRGl+lWYRTEC9s3+4MnwRo
MwCZACFfMf5sREb+S9xwu3rz1HyxAGALwHIcraIwyWKQKf9cTNmE/DFuLYb8eYzD
Sh8111ndORrwKzeiNpEwLOnTj6z0YznUAHC0k9TzQBWTlHmkPPDm2ivrBszDUHSn
c9c/F7QMvxhfIih789Z+AIfA9VBVwttwpQFuxzDX2tvmVEmDG1Jkdl99zdFs4KvS
Qifp3DmwE5i6Ar2nBXHuxqaiFLtjAs50Yj8+JT+aYTl4XMGTtHsO0eOJdTAbQQm1
hHEgddXaW2t+4MNwrdH5ddRiz+EHkwhIdCWBPL7Par8AjNi6iOp26YgvznawDjQ5
++YWj86QKoDsQ7ZwIVycgQia5WyT/y7SRJdC5XgfsOwDY+rijY4atxSeG0K6an1g
4MSDKGt4fiP3YOeJ1uF4PDp7ccwtPS0c4ek7RhNbN53KJvYT7+kmjjogKZgYmb6y
0yrHlboEXtKYgF4x6eXaBqchz3ppv+LKUwRmwyO/3M6qttA40PbT+0queEN/LmC9
hGp+15lJIjG4ghCBXLIqUIlwOjdtAKcgM8ISzOSRNUMeJ9Yp+XrwplVuTGgGel/N
JtaT9ucMYJ6obkCF7HUu5H+TydBVHg16taCT/CqgOmcqMrnLn2WwteB47BtCN1ti
/QzbtaLQc34oNTgZySrR6GCWM/3DV7RUCjsfVDGC/d0I+/k4PnqAuiv4feeZtCgo
cvqZNtQkexZTURcGybgVkG0IHP/pprhIwcoieUDWK0Z/UcqRzyWWDU+k2iynjFor
dLKy3/a42xvm/xI+W2VU4EC2FD6lrSc3zcSk28vrpmUkw/+f9kAR45QhDTiBztOj
6Eh6HYVR+Rq8Bw3urMo9t4xadRJJUUMYSqK8aXQj6R0w+ApIvYv8Tfyu978ucoqn
NCDGrbGsXBx0kTqZ1aSru/GpF9wN+N4vi7+wOlx3SeUZv6gkQ/XLFMS6xmSN6BRv
jJGeTB8oX5lhV4iI0DvkVfkn25VHUjjLPkX0iyuNLGTCtZJrfE+Vjddu7oBQRBLV
Uv0egp3rSVGWefBMPHxQI8P6Ucicc2h+F/q7kG2eTrHMmcTxmlIldKyZExxk4Dh4
tDJhji5772pbmt+1JDiUFMsiNVXYmy8PKjojdvNsCQwNbstS+RPvZrFOTFbw6kIk
p/xWAPheeP9mzzhbFahG/h4rs0nAbEz0uHVADDM65y5bXEQhwttljcfePZASkFh1
76AFmEq8cuyuuTyAdscck9y2FRsuREPrsDDdK2P6TP3o56ZgkyxrQwJGH0OwzcZV
su/1+S2fYgExHQ9fYbW7G4PlwZY00DBgZXXkE8yUJ7A080MRIVxE3jfmoVsGEy5D
bJULoS5YGvm7C6ab4K6sYZsL2v49WJHtIrOUjqCDEnG0TFwxVQsmCryksHtURwVc
wvCfN9OxwE0vLextzGjXL7oSKQzlB2nlN1ypBTuDpo5aliXDiWQAghyQK9unak2L
xrXUS0AqfQzuz8ZUhEewuF5qwmrZ9Swry7fqtW5zONOPB9RrMWqvsNjzJsNcARlN
agFF7C/MvBGN24RJVPL6JlZ33xBz2n0RV3oEyepSWYKqBRcxkZx3KuhElcREWSjb
8nPgmaEI6eXz05FbO7nfosCwlRhL0B7EUDmpuy67Oq/VVkMiEN1FtIyl+DFT1LWS
2ljSaXqz9kMw/F0qibcUvCnasQOQqjy6IxepSh3RxbBqUaeQ4bGDxvZyXrxNg5dP
57kZyvpAJALKV1Xx+Oy236MtyM+Z78pbg61ELltaVlwh1HFo9hNsAF6oHYoKQeEE
eK71FXipQYAWaQT5OECCuK1o7ngWfu3WRp17wrUiFLt21YFJyEnN9CI6kpDIh86e
VQvw/SUiVpislCyjXDbeMcCJ53W7rcdd+PbquC3SsAyJrcLS7Cr5DZadlCDgVqa2
VjY+XRCOJzgDJ4/Cq4IMfeEUAEqV02CIC0MCsDLHhEix6vhTm9PwKVxF1V4GwpTF
6P30P9Esd5euMUWREGUeUn8p5CVvFzp3XV+V8FpLjQhZnLpXLWQAvvMLNZ444g+X
x6T0upFC3B6P2yhCjqfwL2MPSH6544bKSzn6D8vmTtToDo8u9WWBm12jBSbYjfZC
3n+lDqs4DGpfYW4dYk+6R145b0w6ZmIt8zFULI/axSk=
`pragma protect end_protected
