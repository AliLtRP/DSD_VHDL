// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WG0nK84nacPUEVllOoTqPw99wvKlA2JBGqIEAbxOrA5IFhp/ogInSVOd9jbSPDjz
/Jyd+AawBcXiJ2QrhYS0Xd7iartsmFnJbbho2u3aP7CvYOMparPT0h0Tn/287Wk9
tsPCp6LQd7B6VoYLiWWujpSxAwO0cWbPo5ENteJIBg0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 40272)
lxhTy2OV/clEMm4lfinHA16k3d0+Yu5IO4sdikXgQr/VbK7uFx2ttNBmyrN28r90
zIsk38AATbmct6gFhAgcN9pbYe20Uqwwwl72OEGHqU3IGGkHxVRMMycH5BQsQ/pn
ixjcYXK/hf4eR0zMTl8hsfB3VsSm516NL0HMENj5G4F5g3Xi+SyvaF3oEKZSmeVY
nQLkou/ufUc4A3AQpdpHX2NyHQEjHWW2wNs+W29d04WNF2oiA6H05fkGXmbYzhzR
flVpF3ZH1xagQCg7pcCTZ4/LRxAMJl/Oj/k/dENXybRsc9p/ujuQ5YqsspFWwK5z
UTImKBBKB1BrYY5t8Dw/mF/Kjt+t8VUihh6wcevG4nf6xcx+Jy8O3dUeihXKoqQZ
fbunFX78kvl5rraFqF6FgctEiFdLcU+DWy5jI1KPOfwFF/VoMa45zWuXNJnIhVJq
RWppA0pFl3uLPB1IB8uiatCBY+9Yj9zZwRIbPK+ikBYVPlLnN9grhXaMAvmz7axF
c+VzY0FVkDcDEdTjBm/ZfochP+9zpu4LSQ28/tFtPn5FVKQIp/B5x6eWRYsxsgOp
Z3rAsXAKPulSEcAyDhMTGSQuwXFizKwAN6t3KTxmvOnXuHuQubuTGkUWJrQ0OfTy
46Ita2+adRrfcMJaN0CUZVutzEn89yDBz19imNHISGTlu70jcbjyiNpdk5y4VSgL
VBPKoEIIkngxmbFIWkrGD7D8vFOmUQ6OlAw3h6pFVWVuQFyJ2j7p8lBXpsVfDYlb
XP9nIEu6+ZInzB7dwz75hWzWjiK5flEKmE5c8M7fxTn1fFPt4qaflZ9s4BLvOfWM
5W1ehMJBHiJkkNA066VNsEAaj6gw8eCXjWglWaLucToVrPogY4JE/qY2hDgLZVtA
6E64lRBMz63TTPFqbpIO/ZFtop7CY9hRGn1MG9Ld1Ce9m3wkKfQ5GuAKpK50kcJF
qDB1Bsf9HRNhq12kR9U814Xs8vbVe1/FBitfzOt2dRYwzl56B322X1GUDiYad/7F
FZqdSy0SNjDUMoFKhehJFoxKl5u+EYdQVig/R3BPNdQDJwpOnaEJ8ZaItNdDLsC8
Y5KQBReaMUo/bPkcw2oCpBJZ3zbVhTNU7kkqJaggR3+aUn3Xfhp5o+jGVunnlVtB
FgCpHYfTp3LoQujwKDXTumAAe2yEsQyZH+gejcDOafpwOoSPyG/GybSgFDWGnT2z
qY7vlp/aEo9myKB9YQqxqgfZTA0o+EOAhLPomhsywoSQ9OiNxl4kZTVGjVuY5w5p
hSZrfUnE15PK0yAhUvsP7MT1XsF2crgWS9GS4ab3PuJFYiUFhISxclfcp3uvDRRn
Zs9xvQR9lmLC68MNNzN6sOiQ7zRQeDdbNk3DElGd5EkPwV6FdX4WTGqHLeOELVay
PZqBQ1HYRXu1lY8LEuSUBEa1eiQLBfk5iaKQespDKBBZzssZZskineDKdt+eUqHM
Dg3C+g+e/v6ftimkS5zg2lAJoK1RdU+TyJHxG+oAIoaizTsMZdOEtnH1S+79vN4g
HL1MtJ4fmQdfBOMmU683FtpEa68/1R7Li0UGH0jnCFjjO+wErFx16V2CgHwKrkyY
sm6g6UKbzWPhUiIKvhBy33CoO1jg782dsmSHOaHa4EvRx8obCJTfGhlVdtSTGj33
Qsd4hf2IROKTTMAiaNgPgFwNzs31/T+cOgXV6K+y9EaF+R4fdiFZc7rOkpsXdypM
oWGbEFP//syg937GVmAiTSC48sAP71SSocX4f4e5An531PXBmx4X93h0cLs0TLKo
S3pqjwyB41hLKkgxnmMvvtGpRqdyZIos7Nszpd+EESCM5MLKBX8JWM0dVyuVNw6U
TNaiHKT7eGAh9ppW1xZtlZv3ocjDBEBtzvtwc3iyKohtwbDnBfor4uLVBtuA0FtT
anZpksk8EHEQk2X3RlKGN9dCJh4YFdaAROylYGlItT48tKZ05KW7+7mFYsyu/VaD
w0JUsKklbyTmYj4N39fcFarEQPIhOqLnoxTUqQixX+KZ9OZfYYj54zz6oPlIfH6E
4BBEjGkmSe/y9xCxB2gJi8xGZTfVvRWFaKT9J2vCwuW5RcDaeENrumOOvSvnpX/m
mtbTRFjf5X/yIEWaonZq7NEnlIO/FDjGgkgu0JxnLLwaT2U/pAOBZj+M+SIwbtED
hhb8Lj0bFdAzwcbI0tZizDaFjJScmN0LbKADiBCfnuLHFT9l531TSgrA++DFdCrc
sUlqeeU7M8PLgKwiWfHCtTV5mWsmY7fO8WoIJn0gjkgWEWsdL6+I0nr3n3W2LoTq
sZW1afOmx/D8DbMLxwS4lIiH5AfLj5pXVswmsTYOl4S9OdrS1gJ8LilbF+mKIbns
Dvs4EMP5wMxnSGnORP9PxGUfOdNjku/28WMJmtTsvzi+JZbpgy56gx7UT20BMVXo
G6wGzwm0SOUgHtWuqTcLBwMFNKbzbadJ72QTCn2mk664RPWosFHy1CWEdVTW/6Ro
GKLSZuwTFpdKfF/lMVY2DrGcDyi5m+p6wmW5RYb/4OydlmsYjbitmRlx0tHFaZOy
rzygO69JAZvpHkd6XjuCl1+17d7t9ulFeHWqDfcxAJz3cgsXc+EUn29usVPglwTT
BnHkGMIhN2zu0CJZEAw+2JV1L5L5ki+W/E7nwAb8AiQhWGo0e1a3cQ29L0BlPmJ+
2CUOIYvsTD1vgcCEYGOQcHD1Bbq8ixPMvgq995mM3Fazf67m1V6ahAt3GavxzFni
XgPMoh6DXk3Qez2oAc1zclsDBFkXUoLhtZ1TZ/VWMPWiUdn1S9fLQbGO1JjD70HL
uXJAwSe7sxcDkU8BYUkj8xpipXY/ZwlOUXJ99YljO32zFvt7O4OMr2ma6d/7Ewav
8kdZPZQ09CR/eSXLc5LOp9I474YkcZCjgAOucsXY16mYvKeCDvdI79UyoRnPZLhJ
9FMUD+7PfVk1ZZwObVSVB002V7e/Ii3MlmcUe8rbo10Gk6IruKCFS5/i/D5E6F6t
ltSf4BtF0irC+BywmyGle143lpds5ZJl6gzYu+hUZ2KESpCqbH8rKXx98motH0xQ
JD3c+1+SFmQQIdRN2eH3RJhISNeXsiTkfgPwJlJAhGUuS9oHkM4sbORXio4EWW3m
pCKtKzuIQ58SFTWNUGlGVqckKnFdUW3PwI2pMKqpDe5PGdQ5+dfCeg5Uwx/MmWcR
9156VgLjV4W1BxD5qaQ5GEEj6WimjBRnSBcoTxxLTzThBDybj8eu3jc4mM1FyzqU
KYqI1MIISdX/1hi7rOcfTvTiC4BdfnMezHvug4/zZGhi9H4qc1MEFxyxE0LlKg8b
Diu615l+/00QhxZb9YLgXPPC0Mf6t/GmkguaJ0VJAlPOe+gepklvWPG7psuYNzDr
2VATIsc46YkoRAUVx1Qx4TBPyYGz1QZi/zw7POa2la6tQwKTBAygT3xO/1zUD9WI
Qqk/ER0T9XPBbt2YuozVIcEmDeyIgULZ88fdMS6iQHjGGpdo20TxnHLmml1IIddC
6icOc81fz0Yu/XyMN2gbUtHaibaYy5yFS1h9gfVuoo7TtOQgDkr++vUF1tq2UGBU
/5JEEsyOaurONIZP0zRmAOKRJLtdBnz05S3b7ohLhkARVyLWzdoTWjWpd95FF9Ew
n0zL8sigOoAXwW1Mfi3j7w46ENB4tfIm9TaKmRPuzrtlh7oi4nCb8zqhkd7r2xuI
mfc7eTJVIF4HDFrLLXs6i/F44l8HUTBsWgKHThXRHs+7PjxKO21+DFj7Y1VETMss
h3hSAjLHh9/fxHKSpHs2iSyftBEsWapivH0z0Fo70+bvavYhdG7LW+gnw9X0MwMT
Piob1HQTBrH8hMW2giVUxr0+RTLH/igyRb58CWjwyFg+Tr8v6AZVDD+CSglwG+h0
6Ha2dsp1B2fjZjKY6r2v+61B+aUlZq5bj1u8AFoMpjfqDIuXaLuvcuiTmmSKAO8c
AxksPbYnp+VAZ72Rlw3M+23LAN03OXqYy3mGpsFEEymymLmsWNeXrPtmIqqfMeDf
X49KNojIYECn+EYzGQcZRB4gkBXVtoHvQCiXshXq8KuOi6mKR/AexIXeLqnjmDLg
SPxsQFan9oCYX1CgKWytpc+6Y9EbYzeKUznoc41XQbU2PJHRwfadgKnoFXjejd0A
qN6IWPn1spOkqjDO8K2nm87T0CLQZ6eRET04P5ENKs3Z+2ac419YHA/qp3J2hfxB
oSZU2kmpF85qRaJOx5qq2yVSsGCt77tu/r9mbxc5mxsMHrdxaSaUdk7bUOC3m2d/
Y/07FM4EefCIExu01658kVG46qD7TJ/y5OIp3bdpTakJ8BTXazYcKifErPa62bCc
EIrPvfHDfIu8QlbEAX1OiTB7NISt4oEerlvBxbOfuWc6V2HJ2+CzgfT9eDe64cVJ
Cpc3V1w4Rs94tX7TDDcWwpP7CgseiO/+JewSCQgjmedCTlMo3yzcBNtoad8M0i3J
KTwIgtbdq7hqXnxWm7LeCuyF5ExJTJo5TUJZR9Jv8C3OVe6Y523AvyR1Uituy+Vl
0BfflpBUIQrXJCJwpw3LR9K97CNiWiN1z/cc87E4CTf7d3TaHtXs380ukc2QKs2C
KrhMeDOqCZgwf76soYMC0vh7vdFtAjMzEJjcI4UZUv9iG3OUHAIXlHP088SSNEnN
oYLetwMFFxT/j5ry7FWjqEDQ4AT4fsAGc7PDpJzY6DVkPOjKEixFzq2CTMSt1MUy
Bdwo8pGoSoLKUQvDckqYQxo4c0AaxZTceoVPoZQN79hnQOg1jkK0cRqGX/6DrE1L
k/Y8gslMiVoaFdd8EVEDQUkDv4JTtgVXVbmAz3IydjvkDbfAzDaN2Dpvzr97W69V
kbynnaB/O4809/CT38kHyF3P/vCaa1h6T1H7Z70D2pJU8vN5vsePV2F5+UFOkjT6
NBFoyTqmcoRBBNqc/3mAtg5pvkUO/VeR9mxoKvm/9gRtXeh/GHXEwZZ4wFqOc1HD
K8Xf0utg6zAbyvYnTzUzIPyY+Pi77zkMLVD0cwtdz6n2dI7Kc1MGD2UAXERqTL2+
kfzziy+IbYGWWk5NfhknYmrQ1KptU7xFvH1kBwrT+/TfWlnmqLRYoyb1ZAo0Vy6p
44nvXlOwecvOoNvXkVJ8icU0Zmzu0USZzE1TIBaGZ7kHU4QYbug9cM/PwHXmWPe5
c8OqslRsRzV5vjhARvXLx/R6ZRVe1eOHTyVUvJWO1lTt+6RLLQNCzR29Ay/xv4x4
6+dG9cFGdYDyX6NGqlKp3A3Ue7PzbltLSmkqw4/zDjkw9oHqo0d0ZNc5vAW+xnl5
moZjMRtXkT1TUTk4G5ZXmz1RBN0l+czd241G/mzRYWsygALTEK4rh9kktL6lPM5W
U6ttM1SX0/BrWJmFyliHwqyLpjTl3VULhyfrcQb10K1v8dk1DJjcY27CBlE5isrf
BI6puPszRzONsT9Cg0OgUBWIaesow0TaMlB4M6CiHQvjLw+n951JW0Tnx0ZridM0
zzqHzOl51QnXeclOC3untOnhdUpF9lSNDvn7huYRiCZKUkuAVqi2rfHiQuaDX7sV
QQCEhIC00NeMtkCc2OGs38BFGp37pBqC0BUvqEbl71OsSyhARJesxp5uUmL/XSTS
uQdXqU7pJXQ7HfdM5w7pQnPc5VWg4xIaMZs6JuiE4CPA5LfePjNMvFcJSlDYKz6v
ExhL7WFsXegWQHDzAbYjFyOSQ6rfUq8kr8wMbOHipK7+G5B+hPdKPBTUnLNfzKQp
njC2PApYO8lNpTjmY78EjioFX2X36/FiS+2/ZOQXO7+UY5+6A3uPwNHpWPqGKzxu
flGqm0nG3TAptdDItVxl6xKEHdH4Hu2jyj5TSNpMCz9OZGqeEGXXXBVo3VqS+8JJ
Zmh0yuHUbkR38OwC8eRXJ9Ix2nrBQV2+i7NdufkXh4i/Nq2fBc3WsxWzEijVGiKt
WzmBWn0ncoE27SyqLk4jVDX9DSHQjlppuf57FgdlwWxfsKdz17GqvPnYilGmOyLq
mMLoyvZsJY5B/zIpkCecPPcMy+KIz5pXIA2N5NpKvV0IQ+yYEJ4/p0hDE3xp3Nml
iF9b18q9IwbRj1ZUHX9akXnhfZYllklRVFrl1kUtmFF6PASleCgvQkM0WW5A3uOK
TqzXYs4JzkBw0nAMR5EqYiFQdZmZSsjPrjBZRO2YEOTSISYNGBpthqWnGqZY1T/8
BCMMX7FkfcjGwxBzMbyAIp8PYTTRBvJz06DR88th2ia8FDgNi3wMbxlO4AZ3cfCp
zaLELSmpfoGs5pk8zFqPRwagJj7FSaMwiFj4T3Y2MBL5q2v2XbN+InXvbG8zZhCu
Rz9Av11TlugP1j6qq/Cg/+EVTEpx7Eb8hSUrBnqPAcQ31a1+nJtlGVaLwjPLWRF3
CRnTPcHRXM/ks7KQAPgzcK4GfzfwkpCtoZ4vrZSweumOgLquKQML/w0vt3oZdzhm
C3wKyBkIqmmPYWDBZRfnWaUoSQ16ZjmHP/mWwC6yMnYly4oGrKhylufrZYVjFUFo
wUHezZcVP8aqn7Rx/gcAPKGLoj7DJsdJXVnEhfIfIAhiXVynBOzJM1/IAfCLQbVy
aNQsPDL/K2ykMJw7XW9xT/dJc3/TOMklq4rikpUlxClgSCCfnzRV95VeObGQC9Y4
BKtpwH/rXyO5Pb/aSewfadyzjwIgKk7xIT6UD00r9pinOtDjNyPNJwXOUzszjGUO
k2S7eJaf7an3qviw+Rn1tpy3OjW6xBicTuHKs5dH2YxI+BcCB+E25GiSo5khm4YH
ZaFZqlxvo2ro2BMtdQiC2QySjtOn+YlRij979OChcSEVuwa/po7UdcbWEXfiEM1X
CUEfRu7CoAp7sFtyeMxWi5LErvOzsj1HzHccSyi5IR9StzshJaogQRTycLOrdjEv
DO0X2pZRcKdBCwzk+oOCytswjp4yRdGB9BDpGvPu6BdUxPINZ0V5KfOdSd2HHuGG
qxTnh8D54gt/BYlxoCU42LU+AEdeJ2cHqqJ6Lqhn5eFXevIaqnA/XfNiFpfA/ss9
ilkDUR6zfJxm8x+Og6wfy77BjLCRW31gkcjElJo6mvP3E/pWzhme4yYl7GWj1Bs/
KYpFf6gPNbzQIRpZt7c6E7jd4FxpKxo6BCl1MtYF68TQaY8Xi3X5puGtV9UNm/iL
gzBH7IIdN1DLJb8LBnuqKHKVilsQqrJsdf1s1vNtaeCVGWBVF7Y+fLboN+BDlrWP
HioU0jmBWCSOaY7MomrQ5STVQVWhocKIN6jLdGa9gpRDiL+YwyTs+tiMWU5CQkZe
/FjgXuV3s+QW0paAaeBA7USz/NhASHlEXOGqhDwRk8zjgFfNMDkaHgcM+SUAnCDK
5+oe77vS0+FgoxHjntjvLglHNBBvrnRNsNh3W/IZbp2XDcEO7aG6scyGv44hC2JF
Md/pJCrRsre4oVKSVKz9DQUqr+WpHl5BJQUX08WHQY2s4tlxtUqiPEAa1T7fT8e6
LP5WA7sYO93EPLcp3TA7ll4TmrNfynCEYtzWuN/13s1q0NLaNbbR+XpsFQlRLxAN
EumBeIoStiExChuUFPxQIA+NKDyoWrioa6DhJpWUof4ca3yz+f8oJmGVlsMDOuZ2
tM8JOQqy4qmiq4f8W2xsNQ/PO1ikGc6nUY7Zqm5QU5oOpIMu5r911nLAMW5qAmcy
QlgJqCNKSwe9KjztKqiUPJUeG3FlGlqY3TN0C7RfIVRN9zDPNl0hfcQmpRQ4sRod
mSYFki4PXE3vTKEAMCKmins/i6ZG8efsyqqfuICEY8RMBQnFUTodRuqNyFYXPSOa
oJ1gZaT7opX+ugrayjIpeyElo+//QvqHYqhcdU/NXJKkp2udNcuVwbpfInhmScBY
TJrLSYf0cancod4dsHTTlzJnkcnUg97w7ABWj2txNX2kSriD7rYBaGSkey+XyE8r
F+hkjq46fxShLk2gjM85TyFckBxe5xMJ82YoYGkFuK9MRU0DvZcLRo4fW5n3uqIL
olKg7Y/Zd0NiHSlbTL+Uhh4HAnMkVLlbWMRVlNizt+CZhEreSieV8i+kxlkDHsFL
9QvOu/bnTVolu29Hdk2Cct99liI8gKNhZwgaVndN8v3pTOsAVyAvR7NaH8VA5oGw
c5s7lFRmTyT08lknHt+58bL/JTjJ5W3y0piEEbvMtaSug6GkG5A/B77NSo+wA89m
/uHJa6f6mObv1lTrEIIlDP049bE68RSrYGwGnua5KYWRnqXG3eoze8wKSLK79ec8
hSZsVT454iTwycefx4HzQb1wzvgULm3001+3GpGGjM7Nuz7kLIcL3aCWss/gWDaM
ZIet31B/d8+CuYzmu37oSwYi6xR3gXUbN/N1OJeJmPIlwYgJfm8rrO3JZIxoioqE
dYWae5yzbKr10XThCEkvGME7zG/4Mkk+wWE+WmN57gHQkj9NtYjnbKq+oSsTuLkd
OfKz61GZaRa2i6jR8Sf6veVKbpaITCuwfZKFMforLllDWkhhyMfvFm4JaGm6gHkl
OII+doqo4wV0Aah5ErnnqFSDTNot7uDKL7Vfi0I0DVLvZn/ZzhSEWxb7vx9loRjI
MrehVzgO9BwHC0+IDRD94ojGuo04Mh4JRVB1XHe3p/QDp7rFQuCrJ+8JC7aYTi8w
CTVTLPwovaZz6jh//ocvvskWLUqLtE3L7CdUNFXkqDGvaiNozY0HsRD40Uay6Obo
0A/VMOp2y9+BkpFyLXwophs5zKf5ncxMxscbC61ZveqSn1P5yr1kF6jYNB4k9EZo
pZSeKqOyDPZmv4CNuJbKwslkmKv+x3rAyhcRU4PnCmIPtAgS2ItxNZJxeGLzihdS
ssD3po4sYjeUxmh2z6HuHHygEuUGimscYJBA18VaYLzc+k4HuyUdhFkm1TumTfQu
C31lPfRWOlX4ee4paOX4ZZohe0zvHsTkk5sWCObYOvU45NZHFEQWVPotPb+G+BBo
ao9N20/pqpa2J5b5pOJ/jP2qU/NNHFdA43s/ZQXPWDBBZ3srhbOLYCxVHBgKLMF+
ylYMxLlbncD+euZLSn6YrQO5Pe5XEhELhxNgKrGR+QcgvEWC09BOUF703ufAWQlF
ehc3SUaKKBoxE3sXuUo7r3y72UZtpydZhL1htc4xCJbKOUV7gqqvxllxhu709hNY
rIYkmlmDDE8NBon+tmKXpCcp5aUhUJPgbJuQ9k/Onhof2CHoWXs8f7Un7YPbBXwM
3Q45VBRccT8iTbhadJl11bJhc2CFzBvJ2ER4g1DGrIBTmqV1mUeqr7kFpWg11XFZ
5y2VziE9k4M3lrtzFR3z57DptcYZTFkDnxpOGVi9HzkbxLpZeIahtsuL1wECsm26
EqigjHi8egAhMxQtpQ0BRSqXlQ4KXbfIER92EwTG6ZeJ/Fj0z4hYYny1O9p399ce
90vgUomvWuwIbpTmdduAwRO9pnSnqo2nhxB5KLtyHYhg2GkmY7JIslbkbjv2njPt
INBB0Jmcz25+o9QKH/mh4zD4DCcA37YZM4B2/U6/lpLXAthinlFhMw/jk1axZTWq
VveLwo6YdRH7Ec9S02u8//cy8frGWROMSAdXDOelV2JZRQb66G1z7liG3yCWAaof
4DHDgEdoS5RWtRLdU2EQGc6cPKF+jBRnNPq1Cy02QT8oQdZoAT2LTwnHT7zP91YK
NuLrhEghxX9qRSO40PFhy+wZ/FnL7qFJh6nzqlMzcgRNMeSKqic+O4PeNpPBoPN9
Y+9XbYqYtP2lfeib8zSL05/4IcrxDjDAJdD3qJrQlV+Sw/7mx8wW18uPBuaNj2Kr
YI46AuiRnm1+MaEyr8t7/aBX2/jyjY6B/1MdgCZUJJac5wmH4nFDRRm8RI0ooOMo
WbM2QNXcvZyuOnW6HfROdw0cDowvyL/57EavScVwKyelS5DReDeUoRAyFrYYbNN6
QHuhOtbyarfsjXq3lHr9w6edx87jbr33d0Ts7Pm187DIPiBXroRuJhLTbo/LIDva
qU5dDbd7bUK1VJyCGLzgdr2HLCT3fiIM48sGiybVJwmLnG/FcxO/gX/JL6uB12IF
v2ryKLGA3/ozQZ/rhcAbNeFgevOuD2HhHIW2OsjUTSSRQ4Qn+yUWk95AzY51mWl/
OxEASKB7gSbzaxA2gD6sgtzHSBinH6J1QsLdfh2WSa1nq1cbLe7Nn5K3pl5UaRaq
w3LsqZ4QwADMQJAmiriRStXQbVFjHyfTjY5PD7yDWMNxR/IsU9aa94l7PrGwkvXO
chjDgyulfDzHWbgJx9PdCm3YlSkURJ9+4N+t/iv3qy/OvC14if+6SlDdhhsFWCRl
Er51hHYsWvRZCkLNCr1F3rnqfjHa64NHe1DoUDWuhsZzaIRhsoA/UxtsPk3gNZ91
7RDoCSSI0s0QYNjt1X3lEcF7bDk3xV8TCwnodKuonRoNFbcOG+2aT6UoVoE72ynK
ZbT5MPInUGtpWLLw4IG6VbZ2vt7nJwbt+gqwnZiP1w0/JNpqQLIcWMvngAal26+e
7Aj8a6jUz11uHjyhiSRHsfuCkvKLlrjQsRf3i6Jpef7k/TSXAhfamm5pjcltF6/x
+njj1GpiyOWuZoFs+ZNiwH6xlNnMJ3G/02gyqlWkGwZbklk4Pmhfyt86gr5aev2i
Srd6TE88xfikp5ISnvyofXbRiDyqnb6y8SDf96orw5PAx9y9dpv9u2eNYqWt3d43
712UG40csisrB6wO1dW7BuF89wGoDt/vKL8r/ZE8OS+b0aF/foPg4RlOiQZ4a1Rm
GEFzIttmq5fEdUyhWb+0atqST6TrHwtE04uwen+4wIErwLzXgbATPQty/uL3kPPk
RRGwzcOEB0dKnZOFWH1Md5mC1FUECpimhSmipL79+KjYj6/ix1jAAogesWBMhLn+
20tM4otaYLX5RW5hxw6U7C74BTgb7Lvw7A1za+41Shk5utUG2dGAkbyexcaB/jal
tzlokXzFTvjrn/Kqb2MIPGv59pEorph5oAMORqO6BBuwXz6sM5VC6LbjhnTTNDvI
wE8DAAs/f0ir98TRkhR+7kIEsPNOhSezylVpqI2wrBqmfzAvTR2aiIyzE7q/RcUB
tRfIR7JBLKwgUkUJvos49zV5HxMjX/a+5Es6XLP5QxAzLXkL5RG0j9vSfe3upDs6
ZKtb0Ob9Iv2nocG8+Gj8u0w/33T9igwikW44PsdwqTQC3moVY5AEgiSZ8a5Ht4GC
mwhy8pw6ZJ+fgwO7ViISgx0vsgll90QnG11HsOxCcPHKydJ2q03XWTkDzv9fIF7U
/TEMagbt+WUpGol0YMDmY/6zTpNp+5YWbSuSV9m4MfDhgjeZfBRrvZwGCEH0QIyM
bGdX2KXVCMScPUvFBpC1uM+3yI/hLddUlk0btBu0saofSZlPYEBlgTnc2283XUsD
P/2/upMpdy3RMqfCxdP+/uNSLm13pdcY9WEK2gJKazGttCtgg1uHDZkYJsj6XEUq
wKUfabagf9IlomJtAqavYbAJFyr/v1GhupMGo/5rxDgIg9mMh60ahQ4NVsS6TfFs
7IFP/UKiSnnZBPdv/4eAw7AMoyV9uRfeCEXEHHyPqbmuOZRaZhtxVX8spFgP+v3i
d7FX2Gn8ipt1yM1xPYrEKVasLePyV4le5Uv9ntft/l2l+Rov2KN5pA4+SRRIJY5c
4ZM11DuRUlf+C4xM+zWaUSGeT+7x+X2VffuEKrtuuuKd0wyGjsPrV2Xc/1K6atWj
jxNWzZgdhmliY/1POTVLavzDc86u9Wi8/3noIXc/OrPnjQY34GNCFdz6Cv6tDc/1
hEOXCExoyVlwMt16G1pzszkmpK1fHhIyimXjgEh9jC6t9R5pfbLRhG2reEwhXSTG
xsrFKxThGEoJZoXhMj28hHkjxpRvQrwwdntrJLorxhJ50uthy5lCcV79EcUtTUIf
xBhXC/2G+Hw7i6uQyxZnC2FiJiUtvqKiZD/o7J0YZq31RdaLhNEjd8rUrF4POedi
F9cl5B3NPv/Hf/aSh3du2KvHNMY9TlV0Lr7GZDVwXJKO9DCNxDOtgG/G9044zbjn
nBPir007j5RvLq4vkpRQ4TBCFWLKlNDmnvip6j96KwSUK6StZk8Yx25sujcythy8
aFsxjOAA+N7i45keresvzJQT+lTiiiwaUtkN4sHZRJRWhJERbvohNhVcENqHtMe8
QD/OoJUpYfyLHZf0v4uAuKPYx6bl44pj/grEocK5JwNGj52YnUoY3sK4QsOSsXAH
kBPPAsedfWv7tUM5YkOJoVpxsXqU2xQYmf4cftU56WoraV7Adins7uGDFGCXWyOQ
ridYMQZMBA2wwHtho5O5Igw8OA4spDHc0myONTH3OCz+4kwp66dYnBN+ZEgU2d75
nNn55oOw1Zo/xOX8t6Gh5y8Nwwjv/Xoyu/MGmZ2segHExmSL0vlDIeVS6kv8aqpl
pGB/hCxLXlry4VW9ksiWsGouqUuHa71RSV83tSziWed6QKMcTlLJSSeNV81XJzWQ
zuciFpX9uCfN05szOYhj1KK9nxmRXR57EINBupt72eQb3+hBPSG+K0mLbfZouiIP
gV88QeON/ThO9UhStQaMpTXOKIclRNFF+csCU3h4QDyN4OgDIPAbLhEG0h+5+Av2
mKpYVtGdYTejyO48RSvFbj7ujQp+zflbbkjS8ZJiSaeiupMEFEoMnh9Ie/mLvvrP
efUcmLo6amhHJPPHedvXwWB1cXc8Cjqe84L7RC50JXqj+wrsDqvRyr1I0cSi4Y9c
0NirExwQOz+Spmj3mnDOWBG2nESQ/Jaofjj/MqCnYyJrLj3UDDDJEJo8yv2wktBS
ti7btUBtHhHvPVK8h4NM1IbCaiR3v9t30zap8QQqSMBgLg3RU45lYC927X6TEaEe
5MzhGElbFcsxMc9y9395bseQuVRAJnRikIq6ScLbK7mlSI6SlF/5yPUlaWWl+he7
esiZuqVc+M81q1oB5ERru+f1u4zm4vHVwvcQqoGajB1gCXs4LgSGJX6V2DL+NdY6
DLihhiZnRnzPGqAliwByw0rk48cfwkNekVpp5JyUJ/iMX7KHmVJYeSUbZnyaBBUo
ELpI4601tUdltjZXx2snuV+C4yqZmOkRY4eBt7CULS9MsBpR6bciMHpwdcx89h0d
FCnZtJP9CGm8580LgB3bVutzuK3uxH7rM/y4lSLSMWQ2v3hBnUpRleQbXPJDuMyF
HfBZVTnTdPYrM0yDoGELJ+5SgxkDhfAUBoBp/ecouCYAU1nREmLYTyMe6S9NR3SQ
IpBQG8OZd34geSbjSWlvEXI3vNCdZZyPC/3jIi2KHd+TS45rqp4iEyD30NRfudKR
H0MZ5TkGINn4Hk5/qHBEG2mySfSN9Io7xyEVgxikYnuKlc5aLu5EQCyABPcW8/PS
ZnHPIyEc4VgIYcNRotltviZIp/ZjRErJYZ29t2yGzOgDQ+OLGfunOR1tGi+TnDwC
rXTwdTPQzrfGHkMdqOMw3KSk5avAkl5UCLnIVzl5pnEqfMQ1+EOfLWLEZlM9FYRW
gJ9QCEbPCqoeWOe6Ut8JqM6kq5AAoqyl1QM3IKDviFwTLvQ3sHqxgQjgDnH2Cmmy
coJ24hs/c8pxcXpAi4sSa+j9iDCrQ9Qd7s4w2jAb+oLwnajoiNPG0l4WEqviCn0q
r3jtiSBeK92Mj+fjO9cTAIZ0xTjhv9unwqhR28zv218iXoeGlBh64bfPsHGUghJc
vqI18gGp3yUFlwmoKh88FbGJrT2ot7gF2U07VaHouiKS2N2F0YgZNH9ccOTS9lxp
yC1AwUWGeyUcCKgmczsdoQDBXB9O5h1JBgSZ5ZhLq/kGVGTVy3ptpmclUANjjI0g
AafzyUThIamjB23TQgl92U7tQyDOXM9+zh66jahi6meIVo37MYLCZaBEcsei0IBy
IkPZVmKuKDqFmfqRz1OYB33z3e+xsyngdTm9ka35777DjI2Tr1v0+ebci20ISsDF
zU5EI92bE9PIynXVWT9flmM+sW+ag4WcUDEx0souMQVtFrIex2EejWWfrmnlPKSM
FxHHna2SkBnaShh+B54jYz7OtX9HU1a7PL5yZH5vcYXIlcc5L7bcC0R+iABAqyXc
szBBnwVSANYM/GpxSJTczzbpJDEE+gaRuIvUzGcZtxr73LQaWP7UK7qACQvtFDj2
blVg9+TyQ7gfJgWw3oS7vieHeCz5JIW63AB1pv4hjtdBbxzXX8qQP7V2Z6qwWpoE
A+wDJ3fY0vKOXAm+DW8t42YLIaB2x07QGbkySKdFxSX1RPoAUbSy5CV+Cni/q5vp
aLYPEdEZ3gkOfEA4ZrhhOGPY9BudmFZPga4Ae6Rb+hhV4b3Vjcp1kIFoTC/hlfcW
avSbP5rhaeWG/dXbcslGy4gGPWQfDcSE8krvlOeIj3SMfheWrO5vWrnxgwCwawi/
Mo2EuEAOpnoVzSmR1YqMUxnwKkGrtMsSFbzbgm9MCrD60HK74hDjg1duhmnT5HLM
1fGxdNvJlTzOpAg+ql6JSpbWAZ0glrOly4RbwMh/VreXA8flMMgs6bsLwT7T5k+5
KN+amvlcTa5unrHGyY0TVX55B4CFCHZyUW0U8nEliFw2ZHxyUsbwlsbsmaqAd1C9
ldMCV9Y+f4Q4Cw3b/NzRzv6iUcPAJk9xEnLNZ6BUc6CvVBUiPU5rcRMBeInCYgEo
0nVSlMbVwTt4rETcWoi2Zt4FO9dr4NXwUYihiN91hPzT3V++l2H3OaFWsgnYA27v
wtWEdL2Ime9BWKsqsp/ulXPEXl1ts0pxUaVZsOfJrGdHlYIIUTDA+4811DQhi7zi
PQkT3czzcnI5RPRMruO7mOvefOC+e8RKJxUSwC7TJKbggDP+8+3eO8FxTydwPrgY
TPuc5Xv2QeEsWbMbQIVT8l98z1CwAcOs0bf8KJvG3d6K3OEpjiV4P/doJNg/JLCF
nW2dDi0tMJL4t2A5naNJffKt+tPYPJCTdJlC5RcMteZRbYiaHok31LuchxkMoyvt
tVL6DexjxTV+yOAEmu5uiJmnnw9Qslm9T0cCMJALZAiYDp1Xco8q2qvfMJ0O8+eP
5kDdM6QyuyytrV3nrhodpvHka+oqiKdbDxnlPUrK/kUH8O1mVC4wVT0P8OeMehed
1cosGL4spxmAKVkoWAxxvhqG5ED7/TQ0Z9MnQ3HmP/au4tPRVoIVDE4MST2Z1e94
uEQlM7vQVc83GKMXbnYtzSKOSfafBRKQ+wrPLhbkgGUggX/Qf2DoTY+xWrAJld+G
PQAZXN+BXFsh+jQFydL6/lsFlJ/IcGsnQRj89Qk8r2f1W+Bzt3NukZSsEPXj/z9i
dFHYhOVlAPFGtab/f4ya5ejp9bIDI6+HpX5ynxS1yk85ygZTLtyjTxfrxDPVbQ93
QzNxkad11OOQTtBkT16GVfjAzf5U7QuUOd8pvg9H61mmwqsR1gWzpavv6sDoTri5
m4LQIbALRuKsu6/jHA5qq+Xd3g+jXOIhkjEhSfSKT/vF1gmDfhx35VnPvEyuwhtW
NMQnUpe1FlTGXX1Z62pM/SAZTqoYAlWjFsZzoEyOaj2dDd0cvK6bnqz5XJjZ2tqh
puz4GWqMPOQ3YjRlbArdqR3SLxgd/Vm1RA5cE4dEU/tFF2QjrYn7ktkrkLbfq5wA
h7Z6X9hoO+gidrlm2pkQEf/dQN+z37vuxSIKBuP1C7ZPC1CuWVtfTq2aIEjutLRE
agcOjpZO0Es9ZvbAMWvrNHDaT03UIlcrxLOxy7Da0qwBGIzEqlL33SyJhoBR6BxJ
R6tt1Ni86newskPdkawpYACRCadq1yFygvWoWotRi9ix8Gwg6veAg4o3xTOS9+3F
RWcFuJj8ghTSdF48xN7J+3OLvs95JKr5UkbnQeJOFEfJivx7MGbnRoKNsdObhfml
P8oWXTA7twiS3Tc2KFl9jJT1FpXzc3vgAdHBdrWnKeWSRsb2pXJE/tqmZDjfA++U
XmNrY63zHG13QwMEXFYFq+NjDRws2HdzysreKrdliQxnvdOaknBY4/hgUnduvCgE
6vXWAoNBkIdca9xRc5GJrPyiY4FvY8iVL/tAHzjkwmw9qqyPcu9kmSX5BZERvvp5
15VOr9jXysFpBZ8euFrWKoiIZ6lS5MyfpHwOUWbfW7ErEWDvNJ+9DHpjoO1F23V2
wXccGOppbttrdjBe/eoWLi0b5JKk7v2JwK8fFeySq3HvnxLoSeNtwzIlIA9+/YGH
WkstLsPKbv605QZmgOoeHULwByPQRdXjMxaQnXNWraJASu7KcBqyLbzPZ7TgUVbi
OBuOc0EkMSm5JFhNPqCMxPTZERqWE3OX1mpOnzb+l6ndvPnfRo4US+RpIqQk0r89
9/e/iaiMqa8h+vW8RZg1hOiTHNPGDp0TQNkzQFKrPSs4fYqMbpdKxUix+AB8VnoP
Mi3rGsTaq6Rpevgz5geUKu/GWzOwOsnl3iJkO5tC7b8aWVnjinzf6h3n54mwI5CQ
p5S+60dVFqEYwDkAcvBgoPffSmPDacob4p8KHvEvLPbQBn+PAR498awcrADg4D07
C1pn/bJCf27pTWUovr2A7dCh7OT2fyaqmX0hkHY7zsX20/AURG19+HVCYgdzabI0
/P4/l6XHT16nm7e/cjWK3psheFwZGlfFEja4Yq4M1cqsg+iKaNpa/ea0P9X/OVst
/2IrBf3LQEb1Lh2mUv9TVQdWq/fGFm0kFVNdTSQRi+HK0NGkb2eJHWKzcR+39ira
gFYJLFnEZTwrxjR9Ed0XpidRMmXjEH3Kfn9TI6HuDM9c7Nq8KtAyMsf5OhwuIMfA
4HSuSuTdHkYln5FM6egnmJrUYkMMwmXG48H0f2xfMDWOdMWUT0fVtFYY/rO53sKS
4MwVLE/EgE6JBEbSebgIRYxAxWVfQMOLSUno1EY0BX+cuZ4nuNPHrcM2DpssoJMF
Q50eJqULe6XsSArNdrTYsfyGcvEtqbSqQtHz3lt6ZwFJ2X6vxW5tYVsOy6zNVw/4
7p8sDeObXUBbOBty8F2joq6AjG0VQFL26/E+LOjG7GiCwMgWXG0by9RxjjbTX1sW
uFsqgmo/vJnlBH3/laaFmTpC7KTQWxs5i8r6cVvU8s7LeqsPq5TR3Zk6v7hO79yS
hdhJEbW/ROIKo3sR+yLqLZgm92SdLLUog5npU+vZQrI6UqNWS3axj/5XugD7lCpn
wix6xtgfQ4hTKD1ja5K7Ls5Gt0L6NNVozd4OGdarjan/KxyLQGOJYqWlaSjJD6hp
tZBGn7McrIyijCls3qj83mOwdI6CIx3NV8H5J1w0YVfi+KwtXqytzWlWqI/zeYBj
2B1DMIzbuRm7tXX5YKIHX7KazR7Ox+NHOrbFJGOe+RsWZCUpIvQUyyDVG8RGP15B
TbKnHHlF1SZa64uWdGuPiZI21x2PweJtl+owinj1eIGhsAccTzLaJJHfk7uLTngF
bnLG8bGhhZ2r8MuX7OX/ZHmBRpZ18r0XLx1mTjf/T8/rpsdQE0TZFrpXF6QwjJKF
jMtSvpwE0RjNNkA7BhByPrzhsEZfHfiL0kAbhhVJKSUS2VCFGaZUWlOdI3fa/WOo
Pa60Q0pqZZEDPYAZ5x1cSYaR82U9mtWZsXFjO+JX03jKyxL4TaJAA0FDJ/Sy+kUI
+2OtK5o73ouC8bGxXcpsBsO0TYkv6uxGK/Nhkf82+LpqjGs9ZjQ6s+Wbv7SHZXMZ
78UKlDxzq2EEOMVMNa5t/pMXf8d0RLj47kkAxjNZque1xzyy5jttImbK3WEyBsT1
tgEEKVksKlCMDl0um/4ic6fl9YPbXBA7Pe4KmeDFG46goxHXMsVGJRGJyUdcsqOC
lkjei/hG+1NJr8hZnm2QhvSakcbFf/yRKNWCZeSirlChaSzQzUEv4k0vGWEesDDH
jjhCzhvBRxPyVn13A9io0N/NIwBBbfDpJM86Pn+i2vFKknKecrAeGCf5yNXvK0Ke
XMfYuckgP3uBkomC2qhgL7gkjtQanSYVYi5uoG2BD0FFQMquU67Ga8EKbS+f+YrJ
eujjyy3+11CrizpJsZjO5gWCYPkqZqSiEaffoGkbATZFP/l/r4+/+3MUYjvmH7uJ
bpYBQkX0npBndFQHqwednXpa0aD1tivDgaa/PlqMZy8oajNxBvnEPdOwQ6cMrSoc
ufCO1ouiqzFXmGOg19bgtwUd5WsAV5ZkTg0OAODZ5aN5H4/Nv6gAexclZtRle0SJ
8Ej3HevPVoTLOkSVrRXeAXP27iyFv6Nc8jkMU2WPJRw/tMxcmQApm60Ipc9tYDk8
3ieE0kUTwUdQDHlfj+PE8UjZChJGOGbV/tCrvr1x/tlH4yVp4uxCV7CX45W31uUl
6YVESIMRCbnFM6t0VhfDfZfb6L9E5qRzPvky8tHpQPwsJ8686s0lLgWa46QVGpQQ
3nqFhnrpmgcO7bTu7dPbXeg6wydDE/v1Oh2s1QmzfDvHSnowVdLyzIeFtcR9VVzq
DWOaomR8PmG8xxNKvhn7XA7JhaFIoi3im7FsGSMHpEgf8iPd7ajNJajPgpkv0CkU
usXNuYFa08SwdujY+kcMO2z4t5KKD/R/B9BEfwJE71P6/OE9CP3EGUSTVhj5id3v
ZsuZMEFAPujE7CJUQxK3K+zAyDiK4XS0IHF+k44mk2BzDLN5AfRcXQhoIzzAR7gF
qES9JUjeQTMfsDOAajGa/8egXyhJ/GufCa6jYZvHMQwNlsXsGkbhvks5n2WNuKr2
zJ6QAiagsgvIFniMfNlyWxWAykOzCNR2E5kFnb7ZcSR9+hRuW+jNEF8ewFuVewQR
guA9whOs7Ps5/z28707h6n5qv5/slGlvbppDEng6DrsacPVppL3Xnt/GiVkeAznV
vApdvNhCFYbBNb876bRdbw/tXXpxieveFynIKSgKbd4dYeGAUfmjur5g5HQwYcaD
iXSsRYw/zRJuZPHMmMFyE03jt/+L6J3ukUsrsf+Nr7Z/XgZalCSgIyu51Do9NoNJ
srD+2Gq1fKNFXJFPyHcVqvVpYDjJMeHlW/URDh0Q0A9q6qmT2z9/1dGH1kT0eNWe
+aBvUWuwgcKmkmC/TPXAeZyjFygmtzjBJIBYmbj4pHefcjTx1uxTjW25my6oLfOC
tZuE0TV4b5sEI0LApeZwyF2pH/+nDVJbrbVZ3ULcmTRXAkOvtW4X4Cpd9pS9ufXr
EyXrJXqh2/5PabIXeAz8RO2VGSiZ6VpUoZ21LVnKy5OMg2MA9Y24u5n8eyU2EqWf
a6yWzl0+B8zzSyYiY75uRhHjegwwZ098uFrs9z/xPEscfV5MPTbhU/oBwUIp7f9x
Mi2O/VUMQSX6Xn8NxsyGn48adfg3uLqXy8Xd71eUe1mE89NvT9tJ3WeXIGJ3P+Fs
B+YoIJ6Jf9DjYh65zhFNns7LKj/twGwxTTeuSQFeWSxgiJICY2zdqcAy1qGa94KL
SbJN8qsnnv1nMifXKivZApDHA16Zoqz5oGBIJdh+hKcMSyZUnlBoa9I/kE4qux1J
6K1vrPZ78djDXz6qwFD2FSvVNCVK67iNhnBRHT/ekFn6jYDSx9uo6UlZJM3kIGpI
jcu+SxAGXXJYU6wK4yD7r6QbQVvNgeUyAHbcF9Q+Y+m+9S7Vl+vVDQpwE1WIMF6r
px1tDGvbGvTerYwAlZbJUHtHG4lDflJlRb+7LInLrlNCs+XCbIKL0edxDYz4ppyu
FjMOfGfPowVToqiPLuaXkDCEH4ygbFcHGdoTmxICTjmXtABN1J94QR0PbyCYBe1J
fU9dLx8Hx2nQY7mDbrjF1NKP/5elVR7GWMpmJsplXbIHuUMKwZxpeJLwi5d45g4g
lMOwlZjweIr5wHkx97FJQ8xN+4atv0lG7Gv3SSPz8zGMlK4ME87Z1tccC7pRL2sJ
wfhgj1yIlE/KGw6avGH0JDfuiB9x+UIVpgZlQFlj13GsBYTsIXic1SHxDiGn1HYW
4kkxaXgU214oPKB5IkycZ7PQemuNmEtYSM8gAeXmWdqHQunFFdiikMbHzn4mKdf5
kp8qdO9MIhWOe4oZ3KsCUA3gLRFShiNI/Ai6Drg/lc3DXVqSI+ZaaoaFV4ie7yxr
a164H2urupmTsnEeFmZ3b2/tWpckLiUJiivf/Bv9NN1KsSGTwedX9/NipULeInq+
rV0GYoFvYIjcWKbngIyN/1EV4TMIklh9X2xdhA4TweqwXbeFxBs/f2kxkjqIE4dM
I1QTdFFU4abxXgN9dzNc3iTUVmRvZkDxKNYPerQdtZc3jEEK/iw+Z452D1DFqSdG
lsxMPq2Wzk6m9R04Gn5cX5LVEl1EfBIZWmd0NeSIEvpItPjDk6PCUZIsgORUuNKv
U7OnvG0JPkB9O+pDbkMKVCe+oAe2bH9JX/CfvJTdRnrMg56hWYcvefxJQE/qNMWk
pIhu8wp2QDpP6yfmAY7tGiWMRI+1DlMAQSSVo7fcpoUyWrC6vSxhS4nJ4BaZsWux
3++fpVn3jbFUnRFfusPoFpXCAjNoTq0SHJIDmC6v5BJYHISqTB+GdmAXXL9qVyy5
S4IZAwXbyMWyTJVw0Lx8RG+5gepA9gS+HHM/lwXnhEZuDhkb3nbNpN2srr7H0m1L
RmkjSb2eHmnJLFTZluW1BPp5T8fVtaGUq0peDCjLDL5VmH7jlr0soD3havv3HHVz
1b/1fKy57tIweC8RrcYUBaCca0aUvaQU+sG5+hcZbcpCYRKw8r04ICnAr6MtFyzk
j1WBNYHNjMS6XN5DTVk5CynBoiwlCzH2QX+Y7y3YPhhj0hPeKUdDi1OKj2aGO87T
0bX1cmn7+kYCZddNti1KaiG6HFsK2sbZ8cpwViutwMhQmfh3UFq7+xATagrTXat0
pFaXNjvx4As/K1Fby61eQRx6p4Vn/rzUj0e79CEqvsQ6gRqrR6pyaPU8fgH6aXiU
YArcn/6WythK4Ioq8hf+2tiIX+nQEVyscIuhYm6gdMHMaS3+CGxyh7g3foeYLUQg
KYnrdIdWFf77cc80nt2p/eKhmPFt2/dMC+OYxUxGn0W7GXR7a7h19eSHN2vPEEm0
+8OH8F6iW8akE0r2PRo8lck5RV9TCnJ2Shm2G//S/Kx33ajLNffDIidp00aS9W+Z
QkAQeMl2Ac+sMVsCdyHbuKKycf/O/RS1pyK2Hd9HbnkHkxYNdwefC63V8+GBGiK/
gVr539umDIt9siQLCSNac7PFPvk2uMmYW0g1tzE5vxtEd1zvotB4qNDbbDpB9bKp
c1sADhQVT2gw93js4VMCTqXXWR69+k6qGmuEavAn7XaY/FQGIzUxhSwBTe8myn8G
Tm8iHdp7iOpZSk/gyHbE4I2sgjwfJZGCYqsCx0EgBr2HQkQwo1ecf8qaQKJ2phwL
zpHgejYDFiU0OTF0Qxguf1zQjXfOXdODTcNfDjUCzb13mYRrSSKtMSSACWNvfpq3
HkeKzU2xAR5PwjgLL8+1YtzgWWEKL5jI7BXUoFkcikyFjSPS2o44HEkej/eMOOm9
nlfQOCVxPQnI40mqcNeROlAmDlwJtU2EijPsfDY1kc9oWBgJHFSMKg+jwu4cp18P
TPnW/wO5AR0NmeVdL8MLKC8qpGY0Z9aIyglXrXOJNMFOfo6kePxD0v/UEuOfuB//
6aZZlm6HnCSpCZ815cMjoltK3aPEYHFpiJNPhYBr61fXmnts5G8gniaFJ4wO5a1E
V8WuYfxM3sedFq1ox+oXF0YdGcro5LwEg36tzBzKvab06HVTaa/AMau9nCcVUEIV
XwYtPMFlY4gbHDPLcpVMfx4LCUyh2SJygGHTBIceOoz7Y+kT+bk8krNoA3eU3C4K
wDfAUWnDCfvDJrrzv9MHKGESnrJUHdXAbpFrSh2fP9lPOga79gXkIdp7qJ4VoqbH
stYcfRtR8rAYcp//VdqDjctgqZ4fWwfxBlCSdSgNE8AJR1utghSDoLNEj1rA8bqN
vzQJcR/a5q9ZwKl0jYdCFGzbTCCNdwYLbrcHFeq3miWIm8OjYjHY0J93O2CbanM+
S/iYlDmz8/5IepI7tuTpF3qOVFQHoOKF2bd8kV1UoQba+XGAXPn7XMbjKTHFPc3x
WpDhADBCt5t9uBpcV+4NpU44CLAFJXSRbEkrpBtAArPEoHM7CX69qw9FZMS6f2gY
7XltKJqeH+mgOg2d9YZzP4O+hPx4wZTVKvQyeg/VwKVeUKyhtBQW931gd8c0iX4K
hYtheOaHEZnArRjnZUwLesOutdrjOvq24aGwssw3wyeT5g6e+tcaC7WNvAcTaNv9
H0fWha6gA1CBTFnGSQZt9dMW469/Dy+LBNO2fKpirCflRuzOfI8tk4dhIQmhPX0w
bf5HuPpKat1Buqj4QhbmmF0qpP2xrNoxNu9c2jNyYLm5RwcUkdtAVm1ZecYWHylo
6rt/sSzWBUUCx4ksOB2y+DRdzCVMBOL1jyBi7gycWi0uXWri1Kr2o07klFvN9Wwu
Ow4A1MvqEYn+dWu1yn36Lhkg3aldaji92yOq+fqTsDtVZRdrCF1OQXdViw2GAbtA
CjzOYbIVHNtUy6fXf1UnshW7Xej9GatHT+qSTnLlRqgrGtiek/djeyqfn7ujLjsl
XKROwcmQUrA/xL61UXopFDJ81YMriUvKfgxrlcptoHBH7bI/cYkUpFTFUuKbKAZY
Tpzl7HsOBgPRKjbobvj90IvWDuwvJwBeqCm49Z99/YpNrWfi+FJBEAAMTAGHBzIy
ebGJmOF8oPjsGzNZmGPCV5DG4Bv76/zVJ/g8ZhVEQ02j+vjlj2u9C6Vtism9OX6Z
KcLFq4nJhsiXiAWSBYYcz0jjZGuPK7pnFcXWbLauLFCorEXU1EaOuTmi6YvUt0CT
V2E+GORjAf3MCqzGln0B6GxzlyDSVpUKJa7E6Fqw4ss9MwET2jAi25Hda6Mpjp58
gOGKyWVs2Eo1iR2kOc+LXMh46k4feNqxuyK67YQciY8pKWulTUcwXZkmUu+QkZXA
e1TtcTNNASXaT0YSjBli4WcfSEpeLvXXcHOZl22ojF6VJAVwxdCjnveY3QoxYOpK
ui+dMl1DZ5vjoaH5hH9CVVBnWyxzKuWMs3qRmQD6kiHpBMt4JirfEakVLEd9Pju1
o/CoW2nTCs3jC1+h7sbzHIozG5CSksrlkfdbsWVxLt7QLAOC1ftB8a9LYbewQb2A
TkzW9xPNAKyqgugmYQ6OSjiD3SWx6DsBFonCtdxeA9hmP0VuadtnWUWIJnVRP6Yz
J3dkhd8PcQ2n33ccUqWo4+o7A5wyfqnq2+hy8XFpT+SDYmswCGWpyWqT15sRqUUw
onsmVjVFWH0P2qHfRm2yKAa19d+N+dnP6XeyrueogK+L4FcVIFWz8Kt9V/bYhAx/
+2WOz6UuHJr0TI38xJzWfYKgZsxW7maadkO0p5Wbw7HYxgUqaOLOkyaYLa1BRIxw
I5cKkfiP54oXp0BLEJPuxmNdHzQ5Y26N2uugnBVf+uv3xy5U62XGr+ZhyyvmUvmV
yebqk9sHFZiTU8Vd653Thz2YVyrmPTtNOdhH/sjMI/iniVlFR5zRaEG+Vsptzhbx
dIlWD9tjzJtDwxvT+35wl6vxMtBmTDvvrCtRQJ0X9TI7CHbsjPVEfl7zMC8LqXy4
ayhacFmSjUOxLMzqBCaYufWzIHgFwElSUX80xX9w2eGWZJ6j2hZXNY+clUQBAPXM
+3sPDWeXFfOyH91t8INGU/uvY73FVUL6PAdSqPY+0A19D35vNiafdB+kYsP6/LuG
7lDlvSfPTPyDE3sctZ+OyHWz6Pp4+QAT2n9e0EyI+IwVg6bkErwP1lhPvEUX9NfD
YkgO6zHIV8sR86CYYA6XbZHc5F8MO8nOgOCAHn9xEgQK+Xhfiex/A3iLA74iKUzk
Ikh1yBBpAbnBSIMp9kvLY4TF/NXB8tfKL/8faqcfLmOrk58V0tP1BVxXbahfbkBY
ZCXc1JU/v1xaiS6exdVzq5c+D4KbDvEYZoOZUHHrv9+/VvkPAlvVrCDknkhElNjG
Da9AREfTEAcLM89i1vRcP4R9CIyliR6XeAwVPayP4dzFJ8nIZ2hUXlzEC1takld+
UlrJTwdLIv3KEFWDpJ/aNg/dwXgEJxtuxCDXI0dfPdn35T8ZYho76mn7JS/Vt1AL
vdRzuKe1E7LWmGXmexxcLMPlKakkAUJG317mRnrtp6IOY+lNRmt16exXtJ2Mb8XQ
Kga+UBXlFVdiZ7nd+9jsU50XpQ0G3CuhO+D3FGB6IG6XCvZsw95ulz5LTrhNl3Ng
9oMhvyN63jk4UYhsJBhWP9ptqOt4uFQWlh9FeqDNRih2ius8WFJoujpZvHvfkrKr
d5EeEhbIS6zktSXAPw0vQlWcMq6uwD68eC1hyvtYUhmq7VBkUZLn9L0TaVMpoIxq
9aSUuxHkUqNpdc7Gomu3sNRgvHV0xVz+yW5zSg0xToks1SB0w/n82yvpkOXFnT/b
ZxuNjLiSguts5dBxkpXOmseUWbLiXPTEP6fCbSHdY5rI+LMqsRLrfXARxen5yFbt
6j1PRvAqQfDcEVw+F5QR/3D9nie2FgqA1M0OwPD+aysYiNl7UuRV5fvyn4XP7vs8
jz+xbHQw4ik2DZAmUb4z95M3lnjxfajk6wV2Q46kJ6dMCob8zbabNBkI6Zf7sTTp
23S9ThFb2xDms5HV3HMgoQ/H4rsGM1pkxiWmVqH/9/cD+Md0EKe2yfTM+v2VIC8g
4SgW+lh9hJEQVQ+2LnJq0GkU8Mey8sSkP/Of4T43h5Q8WwkcpfAbeX15D8vr5Syu
gEQEkagzI+SbpOHMDERQ9APGZ/fGxUYsAO7G8HEAvf2ZLyvqeaYT+U73GidC+Z4Y
RiLbwpxZ+/EMPnmWgjmeSziH5JjcU+SA+6orBmXIrREXHTTXP+LWYb1dRP0Le5iY
Dcp3scsK9nPqs9VSXuD+kRwf655WUOtD1u4ziF3CWRGRzt6yKl8UHwoQacg2LuUa
RGKLKKPFsfFG5Z6mCgR0qhDDbt4XOAnGL/uOotc/tKCKeJAhXs+DerX7F8jGFQ7U
QwvmMfQ7umDVw2m/OlpeEdTgIU/feJi26KkJaEOT6jW/yAaECx+OtCNxoo5zT5fX
rWMh9yBEMTxlrfbFqmPFFpMitSg6Sv2zDrzbveNBjJ8+H9WkZTpAW0yqjktdq84Q
O8o8logFVc3sxpAFc4Ce5x2LJtnrp5WZFHdrqoGMpbg3dhTwjcJtCiWeJAx8r36T
dM4EUpG0Gi+q8f1GNUW/6NoWBhc25JUgkcFXq1XUz1NqMza689gVnSAPG0kMm6KS
j57+xKoNVmhO5QSWzQ69fq1Q2T+mfKvjLG2Fsuau6dtNg6TgMy+ZD+LxeS0vGIe/
HH3cuitUyT4Um+ZxbtoB2Jr+ryRwZ0xbdDhFMHmqF4L//Aor6/3XnpBPyjKKtRpI
gmQllmwJOOB1xqFhAsi7SO9YiRSRfU23mxL592qJx9MXqL630MlsUlwkbfzE1BLj
Cx/VGbWGgtEjvjR6HIRitbZtEtfR2rR0fpay1ccEezlMWstzph0pmsT4Ahw1nyTP
6Fxflrgr0Py35+sMZ6IvToho4zs1zxXPJdfJBU9SdTDJFvFSQxppH6uH41overO3
ISA/3Idz2aSoKcUFiQLAgP089bpW1CLdoBtNXNvd5MJsyfgezgrB24t6bV7iatc9
UkTENQ6OZ4f4GvbNuFPwR6bCDMXc+b7p4ZImqLkr7X9w972dEBLPdnl9yJoNr/Ih
hHUr50uRoa4dNU5IgMOhl1XUNg3zCHggjZri++oaHMKRO9ZDMbWfnxXbPkfAfsf0
KV+S4UaKDJ365VLcPDLZvjt5m4AaUbR6f7GFFhhRTF0bfDRb4pKjiRhoxhGBRw6C
IDv2HlmX6501dJDLlqNoA1ShNTvtFzIe65F6I7FOcL1E2UBEKyGL6VCr7Vr6Ctnt
QO841sNM0k7NSZhZ1SCQeOOSzZ4tVY/w4v/NXmBSMA8oTJIptDR5H3Eeboa3Q5Tl
AvWSQCOFXIVSnfVhENB/QGEtpGAPnI+6Z5rze7NdxFNXVKb57yAGjkK6Pbxg2xid
yrH5d2XUleaA3NM9DusvX5hGoGSuz7Bc/mIoTdoiHCIPOMY+p6hExJIihUx1sCmp
czsQEflLIG0esXKMxeTzDjNbC75VSuc7OdhLov22QlpmVdT3nzVjVFcDtO1L4Nem
VcykAky/yJhWDKfVbAaokY1dviM32E2a7TKu/lzqW6IFkw3k5f3VkRuIh+MWtJ6p
tiYpEN55LIxRe+pzLb/OEJXeUg/Q8oBQqSnCzswkN+Ll4nRLTCrbmQSTB2oL3Jcc
NovOjTSTKkzfAYVSDyQjnlN26rze84ZTj3sNPR+sBr+EKgr+QoqO+WhZBl/jAEgz
otv97QKQT9JFl96EmiHR8qRQJ1ND0m/4ApHakdS9h+iD45w6cQl0SogcJZ481t7Q
hLLt4iXoo+jEzgg2OC/XLV+a1Sgp/oqWXZFuHl9PTV3O+PmGrVUjNTcSJljaHnl5
gjDvcvurbTjonFHgF4Ffe774vshYS+W4xb7WxCCOv/N8OBYktT/dZ56eJcG6UAy3
iy4hXvBIaWk0LaDcTuD64ryh5nbNSZQHS1CtleiceITPQ7RgYM+latNXxocNiV4Q
EDwZojsCwpT17+cF4JHXTHpVO/tAVZGeZ5DMXDRXaw6pzn7YKRVrQw5kAXtJ8rZw
P86wxCw2YFb4uoiNvw6UW0klrs++JTC/C1a1kd/RpQF6KLT3JfgSA5SBDlXPSMCh
3p2vuW8G3eIC2H3ePHPhqZFqCKFaY60iMqYQ36e1QdtJ/IGV5vSBHhZREaB3q+mV
5GLgrS3UN4KjmO3XkTWuA0G9Nx1fqr2tZCBx3QN0j+tgb9VQim60QyWzBa2rLdyr
rMrkPXR/HBML6Ifv53p0qNv3vHZbim41Null0oQvBAK1ev3JxoxiGJBDK7iC4SIk
sx9+GnRKc6Rhhdu91UwNG4QXAGwiIvvCbP6kM/4gF7W+JXfuVozyWfVzEAjkPWGs
Ids4A7VL9h6yu5/tcspdgXfcnHmvrgRxRMspDVs3n9CWD7YGwIdkdGJlrKUZH493
DqPXUdIr0Fry1NjwsC0JZL6fJmU9qISKIk/esLVWBll9YJGSXAhhV4CBQRzWHQlo
VftRXBZNbXuVrURHL38FYJt4HGOwRfS54zaEZmM+rtXyW186wLqxWuDY5HJ0eYM9
uVb5BZSRbpPsevuGsMehVK95axF0KgrllsPE0tHhiLSjxYR/t8QBrF4v38SHq8A3
ZKjn0YTi7vFfUWQuF30QZmK/gcqee6ZSDB0sAjmBjpw6iUamYG+vRrJhQBkG77XI
4d9jYwf9gy+4oQ1pFqoig+EkZK9N71HPubaZE05Fl/CrtN10OaUSdyPFfx4M9SAY
pAQ/VyvrbnBNPn8KZSk91EtDo97gp7ID25PLRbDKCPjQed0QwdMEU678kplq92+b
jmHD79nZUrG7+DOoykxd8tCw2a66Ogf+YRKzHXTP4kQHkb9v1Pchw3fDSccsxJ8b
WRyy8otpp8PzjS1VZoKAQPqYmNiPoaa7+tyAF3UJFhWvdY8GpN7pxZwI5Fs4S3Y0
B2Dqh7l3x1jvTKNXOpWGpmYMcxUK5kN4dMNBPoEB6YrQ0NxBznKivTVQLmL/Tl2C
iSoR59KqFEuPp3UPqUCxLngMSAv91xta0MYKjs4zxBi7rpLrRuyLcljYK4ICAw1d
SSnwGP5wwXCpQQngQYZpLTeRPG7513mgGQgfmadt9gvmZEz1xpX4dAFy67PHNgpa
KcSt/vB6bHd4sljcemylyN7BIBitZ6kU9gpEqev6gRzaSiGJWiHWKcnatuQXZbPg
UCdiiRxRlpdXF18h957yV35HSvzwdlJ6FRJ7db6BLzj3znMWjPauhfiMRgjtyaRf
1CMrRNo5fQ2vVxhSUWhL+Ss5T23eYwnP9RoTgAnuJsOWkaYwOtIqg6PiBd9ZSPGr
fvyT/6URrWniZb2vffjK9rPfhzyL9pbZxARsPuk1w9QotR7NDIUjiuaKvPOyiHlk
y8btgZXfAc4+2rhv1LRcjo5fO6LmYdGYYST8AFW4uNnM+ptpK+bvLE3sU4tqKglW
pKvGkjqApTiaLLkMXiKeigAkwRA6IN8t4RBQLtfxIxymgK6+GAPgR58lEdQ5eMKK
Q8xVRZ7TrkUT0fKzmYoIs9nvA60oliUAyiF4mq95nPDYI4iSipZrvKNqMShkeuVG
SyKeR+6qiYCn4E2hgVA1P/pJJy1pxzNpqm0n4hR8kyfvHY9qtAx5aCVutAGLHm0h
xIxWz5htHHNtUuwFEcXTaLLKP7HNWNkcXKNwGdOqRq1Ev0r/Q8bVABBMiukeoD2r
FwA3epkDJo3XB4OoeXDSe1cirF5jlnj6AVrbiS+CMpJFt24Dn2xeuZrRCF8uNh/w
Kih88JyXIsxlTK1XjSo3gbyQh8AkRqKzt1nnvkWClmsPsb11QQ3cUMTjPxXVD+sb
rEONOlvDhP3gCcuH+6rzY7uFjAkCAxlEObBN7kcuHlAEDzCeLQz2ZcaLBGR3Bb0i
dA9KWj9Jb03PpFdPArfA0Te45t1lcXOJpdwGY2pCytyqF1yw6z+RZBJipj/e//Xq
vPf5WGEszkC4AI0BBPR02aAuxr3qWdY+Mk55LemV4fhmGiuOaWlx9kI22oFM3rJd
VfhRQvblv5Egnoj5kQrpdkWTxiJ5Hay5jmW/VsT59/7HeAQXbXdAjjC44G8BYUfT
m++YAsimFY7xB8ad5HHo+CsgiSMNuzKSSapZP9DoVGr4rl+TmhJdy6ZlVYllJHN7
H3mG2o7/Ry+0o76NHC3oKRCGNAp3CBm16F4Mb+YYAquxzR+ghTmvNrwiwGEpTZO5
aaU0Ke0373/aS1NDyC2aa8GJAg6j2ZEdCzTF1CTQhByKXpack7gbWpSqSgG6hLyJ
Jjrl7AM1iH44e0cQnSANShV2SyW/C9k2K1FOcoakIMClU5px7s7wogixaVi7T21S
j650YlSIFw+BJwTejyZOfw37CYO7VFQnvMUenahi+WwTcRn8s/u6Im9qaavEFS6G
HDK/is4wJ3gLnPQv1HsVzxSxhxrpF0dxJPGlilgJHZZhobZEBsK22kHnWxPnkTrX
YbrfjJRBX0Yrwsv7xVxBE/v7Nkcv0FI0Wl0hpw1VcAZX6ygHMbB8kv6yulmCbf/T
3EO9ameLGHv/n22v8xYtOpqN+9QmyDCq0ge+sUZheJQd14+DnJMaBzlhpQdVTX4a
awObMZL6HAvr+pNxbx18MqxWlcbalpruoa4Z/+5swTKxY+TZsEuZEy4WPw9CEJHf
gl9fsf9ZMsZptEplIYAmVsqQs/J/mW8eimLUYl0ldfAhk4HJrvUkkcZiZj3DP8Sj
dY4bSsSZPf9h+XMSAAoThuLlK1u+0mTNR/lOGyIgPbQzrE2Ygobe2C1J0krCU6eq
GKekQCcv1dH0/3CUGOKSjxaqZx5smNYAiHsikfIapBlWIyiQJ3+KoJCw3KrNEdyB
Nj5XlXkNor9wAPh7ytRF1H56bNx0qlYmnwhrVKnXeblUSAJ0r5zxMSSOsBCr2PnJ
H8G1+8LQQ+Gtd/SA7Vv71E1aEmo93KxkWqQ4zo3gPLz6h7Y/XhHlRlRcVNzUJAM4
bLDzdMVWwj+xqyxz/DGAJCjK0t3EPP9oj9bcQR/cJNghQxvFHl8L6Skt0Z1Cxi4V
W0drW/VnHoYzg/iKVqlWtfLwwYvl8PI1eI7U+UqZbBZQ9hvlmEa/iuvPDcQe7znB
4hyrUtFgTGz97raj8l/xF0QxIhqoWkwlNhpjclIyKDfDZ8FPXcnZ0AJtbcuVd374
31/Sofr+4Zp/uURZ6AW7fSWUqfFEYh+UKfZpqEnqtk+IiRedKB0rzg6xlZ3D/Sz9
kF4z8juWC0vFdfhhWTyjIX5gHR1yZkU7XQnz8i7xoTCpQ7NgHllIoC+Z5cfBh0Ip
mMZ/OZfm0N8DuMfif9paAWTQYMtYagsiXaSWf7DsevsAKW/H37dcWDO4g//i6iLv
FNAwS0iomEnkGXR22kOeiQb5DhbHZF3yTrR95+lUQQy00xaQlvwVJpy3+iT6ew9J
ej8ePLIlk716WENsS7ej3ZJ1x8XZtCT1LR4Fr8gV6dj5nJlg+XMgIZilIovBYLBW
Z/zIXXTv0kg7Wcy2fEjWh82WZwvcWfVGC1Ixr4HKL0leYAVPYkwFoQlxfBCuw9Y0
UwpqZBuQfkBWGjE3iLlm0z/NXDlcfPDC8euXwp8zh1ZXqPASzvQ3wwdcyoG8tMGm
cltWx1DQAykW4U1E+mZbbek9s3tpd5E2xjcN1JprAIOxkpn2sXSCjHV6NKMqlFxS
jRbvLwrlyQLKCoMEnXdUmbTR0JJHBRfTjQMfDmou/ZF/V6/lUf+tLQ5c+LHQ9ga1
oHUj6F/7cJHbcYap115Db8Fcgs8tZx3WK+Alzrb6xiW/5Jvg53nm84Pt2r30kBAT
yTM4w991og2pTJJf8I7fWLj9mfh36x6qkIAxJBEvQhWSQRpknzSwXZcCpfhalwBX
Ku55iDjlEsScPAAMEkljvmdfvqtT+LXc2Iy1L9/naEZmk59BiLbYQlwO94s366sp
zFUhq3/2gPT9TdilcaVWwEnMVidap/Gq41HZ7n/mMDg8YB5b2z9mhtcjBIwXxV3A
1uyTcnwj226T5hdv3VxXw8ZOoyno4oJMCJAqJEPJyQDKVdeXDvTYqUmcb/NJ6frD
bVZNwrIEAHa5Ta+OCJtvzQYDRHyCYS4De6LLqhKArHSNwj9LQnpty8MH1tWSVj88
QiMpyLnqfDSTGupeAPWhzNmPFIaCb4i1CDj2DZz/Rco6uo6KiR9bg6BIz66VpX5S
JTu1EFdiZkLeiFWa/sB6fajEAI9wLdoLV4C9bQHu/4HNt72CyZCuSJRvxa0NZHJ3
JDyp+hbr1i3FafdG9H6Hj4jPsFko2xb39if4fDB8fCpjVycBwdXyZQFMIN2MmTxO
s9M3y9IbzXNUL2TDCK1mR5JA7Aq9Y4FqjVwwXTtaMcm9evZEcpfQuy2QgKF9VNVZ
Sh/eRSFRZrvhcbaTvTT24YYxSfaqp0Maafg6Pu1IuAQwl2asb25VnSWHw5x8ZC+N
2o0XHKl7mzreOl1ImITaJE3q62DKR29benFJOWaT+QRDo9KFZdp2ojQz2x93NZHb
dAo8GDh9EsklCErBiWLvqgziAM8CGuRlSTAwCBtd/sdo4mFoztKOt/pF+ymAnS5k
gSnTcj8+e0kJ7Kpgf0l81dLaLmSC95HsrIbYg6v+ZLjQyrYTnwBqp3hmJNSSnMxE
DXRd/I7EI4J5HEWsM53KwZAe3Q9hVm2eFtNGlfvpS0Q48ihxQE1B4ZZndQe2SxGp
TrxJfQDGhYAQpX/YVsbHY8ieN0jHJzdqy6T5TOaEPvdw15CLTHMt9e0Zy4ZvEba4
F4csqgj6l07SrSTx4nA7PZ0LglAhs58by7z0kZAqrw4pygdJuPntCjBKAmgtCz4a
cSoeJOrPyZI/+u1QRjZXHdIvnX793y4AjmmlN3VI9i4g0N2LD7fiKQshVzv75Uv9
tjjwaJZBFyf0yi/taSUtx/4JBaf0nzy4tK0K0vCXBpkCtF71v6v1jR9q6eRK98N2
H2slVXVNqRgNATCqHZ5n5qcplkqDY/3hinz7u3MAefSGLQXY1Jit0XdjpiDkzDB7
L8eNBT5EuCuCXoLbbLDo+yJLWYdC/2id6uUP4VCUMA6zz8u7Evu5aQ4U4W7KC5Dn
0ofQg6KF9PBEUxJfqr6cLbyRKBWHJOX54OJ666sv9pfFaVWNvOYmpzxaTH8fSz14
oxJyzwIv08SXfovuVhnHDzfKuUYOAfzOqCAdLpS+22o7MWKLD6GPJ3A9Imlp1oAL
mpDkRsEtky9osj6aw7grY9b1iKscHjKKG8TOJx1TCeNK7+3t9zcOCwNpIVFLI/jm
YyMBKurTECS6i8v6C4h9M2yFMGrHfuCgs3WxVMz4LKf8qAoy71wdO0zfRSNSdK5A
xfmBXHgnJAdbr6M55JyGx7vDloG9+N3spFLZ4IOGdbSh37R+XuTR7pGFApv87C2D
Mv+SNYSsAyMho7AuT1UBcVDNdOl1KqdxuMFf5mH3LruEMhOsRmokn7qhZwJyhZG1
WcqTFlqduW/WmTkROeQgb4WWvcV3KHljkwqtxDOqDaBVybn0ElV/N9mAtWIOfs9t
3IxwhgllTJ/4hPissVyE+eRnVMqQUY/B/Rf2LplJuXampaTW9Q2nTCU7hLoTFLKA
CnDYSeC8l+SdCIRrDwsOqBgJiv22k9pebQlO2gfB908AIH+QGrZFWURAmWAKb3uF
GKra8C8/+OLvH3LttjHK5vaKRvob5E7Q4j80Niz83A2lCaaNCP/gniYqn2zmCS2+
GQ7VkEPe8uNEf9WXotvPyR0KZrve9mt90gjN5gXCSCp2KQhAiIqffO1stUFh4Mrn
XeT6DtlryUV3xtBkfaxnUlysqHzgnJnBOPc/6dJxbZHuOeOtMTAvyCmkjqm/j7nP
oslftGkOJPvEbltNfhJLcN2/rZxepQLJAtM3z1epb908275W6Gxa3XX4gG/WNoU7
D0vt/76fBeA73pc1rdNjT8MqyzbXCyWoHBFrBZlSugbSfVSf0BKLfV1uzCVwpNhe
NQgMGVP6124nWV3TdEu8mWwIfLLyRwOgacTF6OFDH0YeI2eAxubgh79cL0fDXq5e
zCSFjqn4MDzxoVzZjK95WNo1WpNsmdKxZxfzoY1oMgLgCbUp2olOJFpLog/8qLqb
TsE+leAlOSkNExchnE3NSULD+nnjydJmu30NB1FHicUQtjmLWUwyEjg4QbnvQRa5
XmsC/7++Y1sG3j69MBDil5fkIOW5MtWWZ4SyydCnCkc6FdVOfapeGEOuAnT7DXsz
fkMe33y5XDOxIrpTEw11wrfhNhmdnChNsQ8ZG5K9yr64lLl4eZcDGS8bBhtdp11h
wvvxc7yNIfCv4NJz6XaKS7I4G59azaq2lj/FBsig8Ccs2VM+VY7qGKll2mmFzArU
fgnoVVLYdxx8DdKLbfEP487+5KgV3SUZvjV3HZRApYHj9q5qtrEREYX9+UFA3X1r
3GXWtAqf6q4IvOoT89eUfk+mUbc7ICH8zrffqFXAiSFvy3r+aLoBkyf+3EKlGWum
rVJXqZTUgGOSHkI1im+IPQY+MJbpFiAWhINgNO++w6jdNzIUz73qFn37CIcF3mxt
YR92igm+v37rVVqJwOzM2pSI4BSleuCIuG2dhjPa/zfFb4ylHElbvTveTT6L6Kx4
/B1gl8kVyJSuo8yMxddphmF+Q4m/mkCludBJVGQlAEAJp394PujXgPIBfbAEpLi7
Jec4GtyQaglW/sPXxpGau/cz+i9J1pOyB6jT5D3b7lSJi9HIn3T7RSa8ATRbKxFH
Avrq/Ss6Xn/SfOyWmwDwZwVaTPQ5PsucfJA85q1j3JUPsjWtPHA0Ed4wZNsu95vV
TlTHSWhSX2LzWhj22gH/zpf9xNCnfi+WA+Z8yZiBiJ74oQ2iaE2xuT+hIWP7mDHN
8KPWEUX/B6EpRDRW7giIBTWvm5rJlL3Nuw0qRWb+wziEw5OW6SFwq4DuTUIVGS0m
vEtWvzXLAC3vdbmnYe4f4l/sT1MYPWXIlahS5Jb0Ot3w4R5DkhC3OziJ+2FkcpDT
SDrCsbOwDXZpFz2eoF+mmFo6zOBf3u+JqnyYy8v/92GJHzOiERXWo/EIDh3xyqR8
t+vA+Cy0RwlvHdPO/4pQRPfV2g1gGtnZbQ9xzvJijxcXjQOBsn+Mc84CJY70kBw2
Oalkh468n0l4H4x3MHb2qrHsNlQAuUmcU/wHg9oO+h6cXUpHXgAgnd1tbxjR2R3R
BKQspOxPM/vQamPS7DnXXYTx+eKXPtzzpLts0j14GMEAC5/L7t71MrybGPC4zHdM
e2OvGbWa1re1iA9LrCxwdUrFj5gIBt8nCPwfmToar0un2gzzDxZJkg576d6GWQYa
0j/Y/ygyHKsCPLZmyuaGanMUzE6nQ9QFC6druxl6EjsWLJ21jixoMAKY8SRvq+1g
bK0YxiOou4/x8dFWBZboE8wmMzb2uL5LUZAcy/cR2N9x4pYhdCWE5IY3uq8m3gD9
Cb1+HIm7YL1SotedI8x5cO7bZ2p5IpsVXfM+yO/Q9TLfCJ9iLeS4+ONOusSl5vhJ
tOH/8rMoY+WC4Vjp7EQ+fjMyJNlzeoCh14vE8nKHG+vEQkp7UFy8DEeCQzrQxw4z
CuTdB/23fpDQ/RPMi5pgwCGedbktQ1xRS6mNAdZHFwHnsfvPoCDtVikCADo9YqoZ
cB+9uUSh5+vh3hI4ifDHeannLLYVtlH3LyA/gEVey4+9+vIKVByy/BzoFajVNR7A
iJSHumbx0ZLeheqDewPF4WVYBrzRXeux7fKpye92RHc+e+mB9nmu4MMrouyLcmt7
qB0eh0V7Yf8pQQLwI1mU6CruxcjuBeKOo5qwTVNeAPDPPzz6qSvEEVjSYb9N+W72
Jzd68u4ETKgzLpVd8HIhGrHeUypd4Y6g3B6TMHmzoDK7KVTJzkNJg1WPFYhTl1uJ
lH0A2SWh5FnK3e2p/G7/uHd9HpSbnxRZVwzOYw+C+YNlC/3M+FlnFtP65OFmN9GW
tevT2btgHb3tvBAkXK3aE6toSSmzZ0rbSjhXrGD3rjIiCwhGzLGfgHW5LAuUmPYO
MNo2VLFVzB7Awjx7CXfcJvsLLITyoAyj/cPu0gUQ3jijZPZrc7EEHo3Do4RFMFA7
h9n9TkV8DQXtmCWX2lZyetNkMJEa/UG3iB8eVQyuyqY9l2tuD3yejQxx7r+/HkF8
IB2q7rXgCvGnxWgpx/ov53L3MGCXwMW5KbgD6xCX5WFqw+fuDEGBLJPAXZup+Rcl
e1/oi1SVY9Mb2uQoBrfa0TKhTAGSQayOTh26+x5Wp0gJbpGyhq/Mm53VtYsKol9i
dzKAdrYRhbzI9t7TtDAATn3kknLMHM7D1SLemtjDpXwGrGXo8BZoBKp+uGlIDpx6
MBb+eXGV1oah4M2vLNL3LmPwtwPQ3h25cjEZZW9QuYahr/JwC4ofLbNHc+1/TNr5
mhduzPATuHCUZ1jt6uw8CksYg76+eeULvp9Cz0bLYdvB22oQrI47a6DnYyfMy3Wq
NCtQlQdXAy4B+Mu+edf9mPV4ZZRwjC80d69OIlWdmt/x3A9so40ejYVyiXOvT46s
jRbFGfLLZ9wsJILZJziNE921nCliNadyH1T/87swZ+V0PKJZrHCxOSDNzu9qen4C
KhT9V3hEscUwST5e8hQwISQFqgpvcFTKoF6wOStD0iJX+UILk5rMBz6zqtxXmFsc
1nN+NwOtTbk7ootGoaTSF3XALqFbgA7XjQxoQcfuJFkFUad4U+E9YLEN6qlRsKmB
R6lTSzpZH9SlWyvwkUB8Mqd5/t9LS+QFv1L5vf+3D/LrkOZyJb72dVnIQ/lPFbqa
iTp+GGXB5in11BNoaVPl3fJBfA/+07sZtNO9yPsUxpBNPpKvmzfqzHniF+8dP30m
mt0ahfXWS6J2gLGHw5U6rAryGfcnlucLdUpgiGYBaU2x4QpuMloevwM+wjZtEXZl
jl3jBe4Q6Di5hu/0xdLCqGu+RlW8r3kH06rEqw8K/OQLewDXOrJE3iIYZ98oj67m
jTOckn7ikqjW9LjP9W/rUfW5s2owVIX94slgultBeIAlzdYaySbf/vPPgHXQ/W3A
7LTZlKmVDyfV6HEagxdLJfNo+QRn2YQlJMaZjHJNLWkWxfEcJ2WmmlkqFVVOiysw
nZsQJeaaxSMy6rRq0BRHmn5H7HOVmsczCGGvfKBJc0QiH08EfivsCAeTbcdd2IVH
5gTC5B2HpKViB+jZjTRars7x1T7ThdLzBp87MseHeCchYwAF18N2ruGGUaGDKQDB
TQPVS/lbV3qIAVUrJmdwyxe7zbHPQbFAjD5ad9hEouLa0AjFC3BBX7Nx0M/Ks0sM
sY0QqiJmMaQQJudJucsxwvyu6k3l4kILnbqycMEIUZcMOf46/f0IJIAeendMR12w
odq/tuPPWS7HjuGA/e8HutMNz871LydCHWcg/9HAuEuxECot1Rrw0AAl3l3L7oXn
DQeVN96p/Y9pocjyN6GomzXXHawXOl5cb7w7erp99TeIfVF0fzaz/6OPvP0WJHof
A5TU1MhUTxEy8TOVJIoZKxkwDA64CFEUN0mjMN+za8cjR8YVmpIVdNC2Nb5KcHX0
LGjzdC8RL13/zovx4pT+4hxdcyRA8Y6NAA519hCpAIEh69vfOGszlWXiKn+4B9GB
nWZeTQzEbT6rM/Afe8TCJhUOaitjH7Sfssl2ZkbKR49F5rBXbYpqieEkfoIqxgr9
UET5TvUXewrORJFJmyaoOswMKgnm9AyHa2WKPrkQhm8mSvCTKidKXDL2xzwbFBuc
n6XjrsrnxNHD7Ee/8snOk9ahM48oHWxzePwyw/LdTUrOkE3V5AXaUXtPXyhHGxiQ
nOkAtZcqoGtJa4YKwCcqUSMZj0tcRQGuOiJiiVhB6Ux9ij8bhblcR6j46VatzUaI
0nN24KhqvtiSbuoWNGk2r0BAGiagoeapxinGOjdxwEeS4HHIsyPaVH650nix27Z3
HONnOD0hcg+8ECXJk/dWJLiOPR9Ew9VwyE91kH/KtGz59HC0NNYBOG77T9Dsjyzm
E7fRhfsMx7cAFl0sj0QKhze+ygCbnWSn8UXR7xr3rOxiFJeybl/wve3G8/RRWYWx
VECkIjYeFlNurLXYBSrEYfBXCdxpF/Kjn87iRUG7eyYLqKqoFT7g2H692ejg/lDK
s5hcy4uTnpP0lAJGGueuw+fekm5gbq5xbAPg7YmzNw//2IQbldqW/NB0V+VKGPAn
T4sCj4qcvW8vSHhmBUK2FXKMByWjaxpgMVP81fdESCa5gHGah0DWvSL9LzzRe8df
eyy40F7W6p/MKbHIz7LBpz1JcrDbfYKKjewKI7czXnNoGgkQ/yCTvliv4vAlErfo
hxn9TsCVieU8/0DXrN7n6Hmu3wFUG7nPC+AmEmM3EsZUm/qC3r1LbBEfsXeYiBCE
Y0uGz8Z29UTXAQqgxswIg1EpDXPak28akUOXTwqhdjLhFcTv36H7WWEQsx9TCdE+
njgL4yYjVvGcvdJOkikc5nl3qZV0fznlFtQ6t/ID1nFMyKoWMBcPYx28LOH5iPuh
Wyj0l+rDgJmeEp0VALlzNNYS5BRuZXvOhdn/OTUr9I9q+Hbat9r7TPTRTdj0Q3xe
W6BSqClPU3U3ep1i3TmpAb6yxd72pxKxuhMwFDJmCCVu2oLnqLig5WvM2rRvGrUc
vdqtltfdBrWaVxAawFhyM2lu0x998KENfQTdGaOGx/xPjdn6+X2pTiTVoFgbSNhx
Gg1/tYYbQty4OVWsB/RMfVavKIzphRKoWEpyBcRUYN87421Txqxzs2++nvQa34J9
hlXNsr15HjkcEDjnhZ6GalksTtHOh86BKktRcDj/WgYnBQF/nr31B17UnAwskMYM
WH1iQMgbqgfa2qfbtUhZAmDdmyKlXJBawpEtz8UPo1ppA/i9rT//2RfDKq1FPnS+
Qnlcb5PiWOzap3t5TCj62DfnVN+xQnXk6HA26jC8wRCCZJwYnYQm41yeyUGWKCaA
K7QEzlyx8QtJTrNiL/AnWrEMSI/VtHF7zpU197VDUk6kC1b5Dwf9HrQTvU3qoXpO
W3BySO4UZ1zJ7aIly01iJ/o3V7WVCoLNb3qRM77u0a/40CMaG+6fo/RxnXVm6GhK
yh4I0AMlHbLhoEgaoVpw+Ugys5K18BVxmKcsuCSvEGi5cjB/mVMFjKXGYp0NZK8m
2fiaWjsnB2y4+Ki/yA3WLvpoQbuQSl782ZZvM/RxmuN1ApmfaV11FTsvXOcHKz07
uBE/0guQj81ldf87x+ryh0QoLX2Z0pjr7mdvB4pnuEPgzJSbA6HeZmRKTXKWTMzo
BNC/jFmCHzGK+MLD/vTfFbvv0k3OYPtciMDQhM4QA21bo2iQV81eHJKcgI+Tq7jF
4pFbFxlnOJcJe1Ei9j6KEd6FMlrnFTArofAOVrUwXN0weMx1EQSG/d026RBEQKBG
hpnmsz+xV2iMBNB61IAn619oTRi9nZI2MbfW3Sf4XzR5iJVSxFwqmIHEi9teJ9sQ
qxESVwp5eqL73EGKWVefm4HdzTua9+9ulfbxYWL+QItwWP93YYhD8OP90H8mLD1+
W4eQ1VrTjD+pWOJ0fGsYhJCLxZKlLNHWUYvAZYI5aAI+nj5exIqaLt/JflrveOTY
iAWpS1NxkqpRLaam3rs2xUgPrMKU3XL/xAoovlq92651Bslc5gSspdEE2BJ4E1L6
vnu13FF7onBAo3O6GlGxRovM0G48AVbGYUaTnbi4/gbtsIu89O7uYVV9+3szLkYC
W89pzYoqns83KVcCedsZQaoLZfHIQVo351FmkPBmKfx9bDNZDbmuwzqLO72H5W/n
BDS7xsLo0ZICRKDO6KwXyfcxIYi8zkTncEqc8DHUU890NbtNgMX8oFGVtUKUztPw
33whacjtaPE5Fg3+OrNAk2Jf7sxKvrCu16yuzoO7yYG8U5l3KW5i+1uBfm9n9uxA
ZKrAakr2ueBctCIzLVmKG072vU4Tt1EANQ5a7jsSRbz0BCIZtgdI9hcDaJU4sEKt
u3ftecmSwP8tH+S8bmNuraY/CR+6u8arP92BQwmDPUUOi94JO+zkEgLbS/jYXYnR
NlwvV4wxAoEtmzsCW5eqDSt+uK4TU0BJ6MXcfHipJI747RCvbkDHZM3RhB9l8WWQ
k4kAAOgyLUOIyn1XzcwSxbcLcZWiLoNgzlxPybKRfFCMuAnP/u379gZxXaHQ0dvq
7Cmedm9HJ9f+6MD1i4SLIFSXYBxbLjQTSOjgUtu0smn4H4ruY+qDgxopOKteIR+N
6Re2HKEvjbaxyWFh7V1mA06bzRlbGxHby4CVj7tKp27AzjxT5FKCNv845Ggl2iUb
rLo3eTLOi1fvqX5G1m141c29k59fsPZC2f4iI5G6n9RSmDAoKYklYhRGhpDLdP+1
KpaRPgwRD6ErjaC533gS1xzvkK1v8GFxaFcs6yl4w9VK1ApW7lGaAdjOQZb6GZ1J
duK5PbvE0e+St1Viz8o2YqJc/o4TQQ8m4yj9z2+ZsJLZvQBq9I4CEYH7P2Gak3JJ
Ae9Hu2zW97Lj4tEROYj0zvg5TQS9O8SK6ihHBrH7cq1Wh4Q+SjcOtZ7XNzK0RHQw
9soJ8wTqXt9o3Axabc0GF3uqB9IuwXSpWCfbIdvkTS3VpkzWQ2t25vXNK7QKkfKa
HMc2w3+fZ1DqsxEsVCpQhfKheWvCuIvjKluIOwNzjKpWZbX0ALHvOqXI3C54xSJZ
vQ57bjNS8atYOiVHekfSvvK3wetvFQy+5rmAbfXCDN2wtxR9/4YKMwzzbsW/h9JE
Cya73QMkFX1fj4VIRm+y0TDjmDJBZuzIdOatex9er80j3ilxOuODZbBDlw4mpTH/
kzQrg7Dv4T94jgLDqZVA+a4tLK6HohGM11YWKbuT08CTHqKtzfVMHD5skgouLRXw
m1iY20h5l7urxBiiizyMqk2Ey+IbcfDnMxz/e0rwDHiR9lTz6yBM9LyyHkWF5zey
E0s2cYdAMEDU+t/oTOEnAE1teQrrp35S/024frUlEhkwblzJSaQ63h9QWe5yh4kd
+Q6FOLMzq1T5XH/b+L33x5baEFAAiQ6S3/FKsS4vBnsgI0XI7S4gmRvgQBqYXTKD
dEP1/uHQGbPRjMI7xMReb7DwgIFw29YN471eFcdjw8RJ5YmFcayfH0iAVPEttRNO
f1VDBsVcdhmSQ4vDWpPD1dMRxstV4hTFVwewEO1FuZo4pwPcFY2XD2gdPLwUwwtp
MN47ATrC7eQ9KH55JFgW5iTzdDu0vHMYc3JSqs72mK8ih842kcTJUQWz5tH7dDQm
T59aYzr2Hm38xbK6IH9FmXw/FPDsJQ+g9zJlDy4kCdv2yPlsxIHAgkMCsAhcB3gn
JGtTzOYNs3bTovajBq9k7Zx9keCcnuBnfcTrBIi3SSQeGV8rTpyggYyL1eAAFwzi
sp6yP4/X1gmOpFn+crm1Mm96/OPXT29Vmkh40jK25GdDunPVJs1kFbOkqM7RWM1A
YkxY3TxDpQa+/DVGbWljZqQBDv22SkWfjyVZr3RhF/r/2/5W2bYfYkpdPtfEHntv
0GT+pnMSsObEQ+DU274RO+ocy+UNSCcQqHUITVSccVXB+KyiZ+W6gZFvvE9K3blp
H6X+BkJ4qcrpwi1zJdgLy72+vc2CjV9yfyLCDCJA/usAEpdMHz4XM4Ze1ruF4e38
iTvbK3YWhDGWWrKOmkrpNGbVmpH8d/RONw8fUv0Ele4N68ePVkdVXjq4sEzSS+/9
MNbWrDfVfomtem3VQzawm4JwpqFFwenn+GjDtGFEi9X91oZK5nq6W2W0tpez+QKM
gxsfTGMh9zNTg6wxWtQ6EpQVRZ1EfEZoPazM0KRdPQK0lFdBW034jZ/lm0Nj+tNG
p9gui3pHzETgwcsCvPCu1Fax+Fu/9KIcIi2URO35RGvz8HzkApIt+cYMWAoqST/p
Sst4uycgW6r4HBDVt4rKgvSMSU27/CKqwMctcgH75fY5jEW9/R+LbwAU4y5I5hRW
pFE1vuPMdyx/5OXWRqd0IM/oi+2pUjtjGajzNBZsA0bIX1J0ankJLzls8Ay8Artv
eRZMOHqr+5k4qW45Qb748H6gXC5QDW6m9TRzQOJ4y62TD2biLbyv2yxA24ZCXrqf
iFs1ReWudxceOH/1cgbZMA+kyYzP1t42rMmHHOwBpyYQ1tbH1R13FT5n6HKcXQx5
Xzway9fvNtkDQjZrF69hoK9hr+iwsOja5TnOIQ547eBX2l/a210n9LZRkilWmuzT
d2NmO/vGxOX7msdCM1+TeEGq75EUUUcMlrv9P5VsId9rO6rQIJ+KdLqdQv9w4Pa5
IBwbtY6/9EMxhzbXBe21G0bexUt5fm0PhPwS4sovghRfgy2Li5tcujvpdDChlvog
/gmUg6/KLJxrqcPqyr/Qwan146R6M2YlVaBcp6MkcxzTjxtAKWrM7aWMUan/wcMb
zbeOO2pd4WOvJ2B7Vb0ZivjatugwnTAk+ue0Ipw7vl0rB+1p/CKiYQehsrfYddgO
OiS5Yw+w1wRw36YRC3aNJ57TZiQvDNxW9H8KDwyy8l0M6Xpfw6HNFUJ2kAUuUQ54
03HEE/e8DUvy6Ggqg3Wh20eiaCRWzL9ZAQs7n3M+QWiP5JDkdR88nzRbWmxQrTUO
fvh4jbI1h/joAIQlDSE6WRwea04KSg2NGlqF5nUaUMkWHJvORzi8ZnFxhnOfHqXs
Ls694vyzZeohRUIBzWPd/PVVibeZg+ipjrwmS9ZAGBFKNjRgcW7kUaiDSM8QXVX6
UCHnjLLo043nceGF5saigCW5WOTXS6thFLWrPEb0oe/vJcNPKDwm8T5mvx2jkRYx
wcJPe0khtuz3OJWOxfhcSMJGDXAtlO7U7t/WF0izS0NVMDUGba2smYawZxa3z3+p
Rfyqm6j/vT1GZvduORGRp3NYwydx9SBskdC25+k+y22je6EQAAQcPl2Te9tDGlh/
CJlD9R/BdEmXleRn8K8X+Jz5LZQkwXA6uECf7zZfMRDJnJhSkLqGnthvYQfFwP4V
v8LR7y+6W9cQm7+t1CZm3NLm7rJ2pJFhmlEXTfBY+04p+Y8Yk1WI1Get52M5yJsn
sj99sw/IAPBI8l9ZzoCdMOdoBtdtQ6c9wkfttTPB9aH76ixhv50rPRQY0GT9VSBU
oNKtcwJNtVdl822PzYDo0yGju/7yFYF6bBf6BiwCdu3tg2xYD/dWv6oWxNatH3If
hURes+Rasr2VD0WQqdA5Hu9CkO/uottf8Wjtj5WmBehbHfz3w0HHlIwXZUBLYzW5
mMBD+0rrtmHzxevtfXzZz0I6sBXD87AE6qcwO6jup36NjMh+Do304ShkPm8X1Uun
QtnaYQIC5/yQwhvadQBeofLqWMj4KRUfNC9zyzS+ynFBT5n/4iVUxKLRAcQTba5O
1TLYmNbTtaWSReyVFzAfaSwhIa87ikQEnrzAdgDyfYuFcWSUaj5MyWq5QH2jCZZ6
OhmvAk28TXpTauGohBofgZaIItJ7GG42ZtIzRE0R31c+BbUcE6EArA+aLUBBskEI
ZDg9U/lTosT3lI+9/Sn8SEiGWpFh3zVMc7OBr8kuqc173Kj6E2gePjXLOa4AV+79
52Q1/xpsCBk1caRunU5zxHOUKdOvvOjclRmT2ISd8l1YHZG3Buy+A+8PNFjXr7Ry
NvTKFd+WMxD8/rPemQpRp4PSo78k8l1ryGujmy4oyGW7NciC1ym2ag5hoc9FMUjY
dxy8gPYDpMn2JJzThsWB5UjslTe9aha0eU5HKgHW0RKmIBOH77V6f0yGQ7Q2LiLF
ZmmVd8pKLvQJAfU29b53zPsUe4sf/pkhN2sLmnplY8EUnbABaH/mwWXe1TuAofHR
NshopMLNxpibjUGNnZz50K3gt0n9BYC1GC0es174MdgqX8pmYnuJEOa2ERcxpb9z
eGa1CXOnHPwUUGQTDllL0AJt1lqGpq2ppJ/NoAnH/FGyPb8bWMXZp2S3EPNAJwqS
uHJtm93myKOmTok5HO76IlIXZF+YhMEi+PtAUsfb+4ePm+mX/kPCQ1QDUergPEx2
ZPzSIzuMgySVbvT/srPHzcfWGU2gDbi4VEMKg6wO++sXIEV7f3pCHJX2N29xnSb3
ihCNmzu6WyZEWKH0fjwTmJP7zePHV0ZyCnySlECZwDmHzfGerVyj45h3t67M7mWZ
A7HrWQryfe1m7yXlV+RH7ABjubEZtqOaLS0tk5R3fCCtcYJvgRcQ0c0WGMi3eJZ4
L1I5/NhcMdXXTkNRY4GoUDLTKEev/CxLTA+0E8VIm0HSDZsH8hD1ceORH5Qglx2J
d/fKP2zevIscQZAWiWnPnRTX36H66RV4OQejZIarKzo42TpRJcK3+krWugK/QhgK
bOQVE3Cxqr9mT0ASyJOWtvdXdtXyvUk+XcIQHYGeqTO7+Q3iIjqqeGgWOWRoBCrD
GQDMfeRGLqbiqwwX+Znq8IuLbwDG10UMxY5D7keK742QOy25xY5WAw4Om7rvshyT
M7RGTpUlHC5L27BhZtFGw52CtsnKTy6iNN4MVrZyRmLstHWdXjhFGC1PpIs0q7JC
4C0vMvFOVpjGi5TNjCfFI+3gVABARpRO9cgJoX+vf+yoKQLdtrp3uLSCog8yXXmI
KX3eXg6OsC7kh0ZFMHyurxy4tEY2tb4zJ0es9+XFu/r/lbcuSW01+nLaWGnME2vE
V01XszBoqfN1rjPDgC5s9hfWUYnJvgv6FyDTnfAGiyuwXCEebVMygEPAzsQHc0uJ
02h3eT1gBy/5Px+FWE6H1oSHAG7q13sLapZbSiPcMGb37VLxlBdSNrzSnmSWRura
k9bhh2X+UG34kHmZRGKFAANr/9W31N9L1tNRJ4MTxLrP3O4Bp8Nbz8UgbysDy1gb
1y90T0xCMCYUlZDgSEnhHOIdABji1J6zE0b9Hcu6Mfe92f81szociunNmYCcTQgV
CDk06EKAZpSO9FZPtfzDl8sQI1TEP6+ewShcpFodX62fMRBdRYoNyXGxWnpHsX5v
QpTwkRTi70xWx0rnUj2A16ZuhcHwctvf58Ma5OWdG3n5XrhyBuOBW3cS/NWCUWHT
6yY48MpNKYgm/zwQxa1k4I3gN35VOJR+JnhwAxC4+OvgABict8gQMh1Tv8FXaD0q
hyPJY8i5x0ewqLQ+FYKZDVptXEg+aL/770ABEi4cseLUJbMXwvpJLuhMEdYYdUxZ
mNdu5PXBfx/2Vg8pU3YJRQAen5rkOVXWunp8O7sEA3NGpUHpuvhWl0E3HMQO5Gn1
Va6LS7IzgYvWm1hpfRWWjy3TyyhF1U5rkV6eWc9Xj7PYUkncO6kjKSNY18gqE4Br
65Ii+diFsc8PlhUa/7vqIVS6rmDz5/VOU9dJ4XRLY/4fhi0IuCO6CGVgsRBVtiE8
Vr4BDYzm3pye9TQAjHtEHoSwGwIqDzElj++X6Pq5Bro3CYgtlTPOCKjryIvL8ekc
64yf0mZxJY/Y8tp2jmh5XRtML05npR8fdH3yWRiUQVUVGUwv4LpHa0vm6/ysI0JX
oWMU2HxsQudEZTWsoAxzI12jhMj9vcXxxaFVhqLeYr5Gs2guqDvyWqi8CvOJ1AnD
SjDpWA80ZcWv4Z4uvHbNoim9lNmdJbUNMjsCHMs/VmY0X2AosH7WHOkWUwOaX69W
OTxjUg/O64Rrx+cV6BtKG8/Xsb6xUZkBmbw5W3hD9ms66qYgoeVuZ1NciRDJxN6X
9N8kgoDqBDKtaxfedfrJrBdLeSK0KIdymmLyQjB5gNMXXNAqMD83NSH065DpZSrC
H/PmvMu/wNwikQQfDKU0nZ+8HGqZzaXMAydM2kEPXLqyz/3RYTHwhgcjKWmG6EFk
isLo2g4iyM+ILwt3QSp/P441rfLWxlAP53/VFeqJIZKwsLGyFPeh+i5JZgo04ihl
k6UVj5W+ejbIcNyIXKOUh8y27nOGWoTLRrSJ9sfhiRyTW2NbWXw8oQIkKOBfL0cD
oRxVxnyl9PazUU380GzsQuPEXH/IiHrcpNmwXK2qatgkFolKFcCyr0Gf0jdI7/2k
V1nSRiVdI1oRr7IrUiMdfoEsS0FdA/moarOq6uY8HzQrFizJ9IhqTS4otp6LkDKN
U3X5aHwbXpZnuDqvqG/9JkEQSgoZsKKa1Ic22N5C2iW6y5DF0HHMs6HLgrVWxaEK
z7DepIh5mHRZtbPwyZa+FcF+jkGXGR9c5jTA1Ti0/RFovafH6JgPF7xKb1LzFfyh
oYfvgcZqPoXlO8jIZROEPmq11f/Vt3MuBfVUk/uCGe06cW4+//AbHAZQpjWXgjnc
m0DplvaALms5qbz4MD5MbTPc64wGkgT09NE0dTLaxMOxxe9VpdVzoPoB0X+gYNlb
R4XnHkokGttO0vsqa0KuvWDtxO9ZE/ytbA68I3eUeUOpJEsBVDTRT5ijy2/CMVvw
e+a6vdxJbn7UvqjMZTj4rSjOF7gWPcdRcVLCw+5x+i9Vm7SWA4zveDbQ1PJm6MD+
nXe0+AgXbdd1/GXpdNGMjAr0GmArVlW+URm4iUY9KKPPYCJeDJMGwEgKtjClA2z8
4I1Oa+K45BsGV1Q+E9nIg4z3AXw4Gk1AXCg2a9Z8qz6J1E9eWWUMex5oo/pdEd1+
Z62+P+JdFjkn/awM0+oI22gvdpmwx8og8Z1yfjGeCoTWSFRIV2K+uYsYLB2lXEK1
cfK4nLips0HXVo4809cC3PcCglMJEkundvSNzY90lwsQ9E58r/lnqnvem3wvz+Aj
gQApApevO1WItmOlX3X2geP49ANP23g3X672/q7+ZPvtQHK9TjTRk4D/vSYdiVcs
kew2FMUQ3BcuNzRTedLBYArqmX63yAPFeEYz+QUrRxkJ/ODoyiifk3EmlY5NpnVB
BlNeo+7WxeEaN4ZTbMcuc3xB7S8fmJakmCeU6C6J9dpC32KrZr06sXS3BiYWCt1u
kxXDGBVOH/wzv8EDHiYVqB5TjAM8Y5Dg6LMqmN4vnXXgbfhJ9WQdwyzW4I8N/EA5
nYDkJ0LiMmlvPycfdryDB8l8DxenJJ5YtFooH0yV5jA5Zgs8lcPnTzGZu8lOyJnT
YUC4NZeASSDlkCc97lE6IW7MSSNKCliL1vC3v2zWV3h/S2ubrhkUoPKXmpRGqfAS
PSD/Pt6Reyu+txeXLc9e4XOQBJ+eZ3Nq+u60WELLw+uLGb7gA9CkUUUmkl3wAFsI
fAKDzIfHqsr5hj3rOws1l0hbv/mvusSGdY12YtpXO6copDO4CabrJS0CGBCzvpef
fuggdTsh1koRcDlfx2EGed3doa55/JJ0/+k2TfPn2/gY2Mh1D+I+x1O6cGpMAH37
QVMCxDI//HcpK67W9Ozg/eZuGQqt01q4vtRKZVbUcGFOvryCKds9cvGjc3kEAyr7
RVt9owtw1m6M8C+oh7e5NlXngiiTey46IGlFkxmhvBplGpx46rYzGgCF+u4y0Huq
hXcrA8GNXuCoLPNIGmLHoXBXI/BeAFN1YDHKw4odFUNLk71nxCCstndpsE9o4tqI
WHr2W0bPleQpK3UTm5fT8muh8zDaUeVByImkvBB8WGxh/ptKVS/aUQZ/hf9f+h2P
v8TuiHg9s9uOAdLsPnLjT8WUeLTyZfAVzaFSbutTVtCJjA29L7z+d5PZV8bX84Ai
LmS3+yCYKzFFzd53BiQXubzlRb6MSvhVZ2d0vjnBIgCCiVRCYZH5Emaf+owouyX2
sBKkPQeWodJEIBZgHaZHAsOiu1qFigErNNX6WAHhoidkc6Z11RRnnsY3382cakJh
wDFVg0btgiWXFTwFln0DZDuoZfANVkfErZrAVOe92Xl5u2hcrVy7FjKAHJ61wsMH
46HtleX+PIh+54G4gSmSLT3X2Cz05GgHq8ke6xngRcJm6uEjpPW1TEvkzycpuOI9
YzBP0ItOQ2qImiiLTmMkFlR8gZz956bRhu6FqJXXfEQZxKvbLOb2GKwitcjMJUlU
eR6EszIrl1JNSVbejSi/OznOE3jszOIy5qqKkoKR31HsuKo+dQ1XW4auEWetNhi+
cLxvewzC5MO128v380EWPHB1S8PXik6Ik8oFAz/23izFW/IaYuwL76KIq/Q2MjUU
WajoA9w82387tDOGnjrnBxixWjxxwrpr3GDsVydNWCPu//nEfOxNxMrUg2TyX5lS
2cK5fGOumonYdGlgBsOarJoxoNqcgOsypJndxfXdudIdVnTGH+lLynu+Hm2RzdNB
qFrfy0VjNphsZJYAwXxt6SCj2uIX+Efc5gyx6u2l7dsoRBkRIrzRqnseEVenP2Mc
0huJAz+Qpti13Xad0JYPIt+ghYGfnLc+AGfLtR1J2B+BHTYtjLw+kvH3xixyKuKw
Cj1da6pSuRlLUWjbEad0uOXp6Bvept0T9EupuhTdk2UiZ7C/wHjH0UAIqiSHcFsH
CMXMTLUd0IQgMu16wmCuu5WEoNYqulDUL/R5DqC5TlVShT26XogwURCNbl4doudw
GurSw7HytRtiwAIgr9Ax/fc8FarOu3j0WYq9wYUu+bOsll25LYDzXU8Wd9jEOYLF
7lYu86hvmTOfTwA23Ly6I5JbTY2Gb8AphW8G/lzb3UoPqKmQ0M1oPKA24u2lrpqR
vUaF/6YG7JCSpfmshVBTvXD1b6LJmcS/P4N7+oL7kpOsWfgWroY3voLeHEDqo0Xs
21uyUFRVavbbRd8riJ9HQJaUttZmt/0XhRpzRpYXUTs4v3d8fVyR2MMoWFcE6WXU
a9LfoUsze6iR8K547EY9l0UYOJygAJeBslXJyeVcYDVnPw7di+Pex2C0AKI7Gp4/
u+BBzGO5mpF3jsp9X2x93lChvtTKxnfpVHrFYwWCGM9wOCCQcwyVE94s3EQWXDia
Fta2Z4rKoWz4W7dXK7L3IpgLra4Fv1UAosO3T3PZ+uNYX4lzFxBcw91Gr5xuSEc4
qCe6fFsHARok7m8Tu52tnrV2al7LD/u5RZ48bLtj4Pw/sDUGSHGMJFTu55lIohcK
SUvXV4qr5ptpm0cGu6tlwff2F47/Pk7qeYjTSPPdjOKcQfRrOsqZSgYBPEb7PW6X
eYqWLcs/p77llB+KOpLvAaYxFeaHLiJj+Wvo1wsg4RAKgbYTr12DvCXX7rLfqqVc
tzED88HQqZczLp3LFhzRB9RRKwi23BktGvDbLE92nMfOi+SjGYaFYCwdfPL4gooz
4rYtMvflQkDsufjlyYyWJuQXA/2VfA8DPnGJzwTFLA/Msm7dpPgxum95I+ABBNsR
cmujQGnTKhjijjgz5Upg1ZRReVELLzTIwr9OKZCR/ip8dTz4HbYE3KUuousTQgMO
vZ//MLkQGY/MeGGOIwK1uKCA01mwtzQor+Eg68hJJqkKvJdTqalkUSAqN2o950nC
UKEMHz6s/JxrVTMPqEfjLKMfBsLy6y3LDMo+V2KIatmbn89TFyuHGtmCTUtxNB0Y
3BpiwL9+0USEHZu+UYjPu1JroTz/wbZPJw/a6a4xT3SGp+OSg5eVgD/1pg/c9cTm
5FcS6EahTVrMPjj7uMTQ2HRY9nm5dNzqTdg1EiensUqEAaJUv6dG7z50RvYX9Wow
GW0FCNJlkF74ZQPywLaMa7Z2xt4dS5jn7qXSBnIc9AiXzQ78FlyMa2JVG55U0T8e
BeQ8MQgCEKmPlv7fLYak4L8Rwum10sEPcYhcQx6o7YKAGopp9r9ixksgFvEUvgLa
9Cgsyp6InqaBTqBIRO75r64ci3jz8563wH0KkOGobXinrI7W7+5Xs3FM8+OEF7kd
LHkpqzA+nEfNX022kdoDNGlCrP3e6ENA6Euw6pKIJF0n+jzVNq+1MuDL1Pfm2Uo/
GIGM7ygZae1f/XiCbshmOMnZ9ZL4pFo2FWXVQpyY5RSb4c3xBtg+W1ojGlWLMca5
xvodlhZF+xL3L0gDuwW/8r28Fi3S9jbOp35jfdDV/LvPr38oSmHk0r7W/gdfauq2
0mQk8cgMU2LxFVTY38Qajq314ENv/ypN0Nuefuc9Ig2/6mf2W17+NesOjloMJBSj
LBhBbLlpr7E+5uGWrgpJST+8MtVIiN72/o2Kk0siOcx/8pr3lOwMm65Avn4JRp1E
im+KNQz4KIP07tuFm1SZIkaQC07jUndu0z2mQ8I2u3pY1sOebmLP+asp0eBDGKe8
J/TIVhQcV/x0Qo2xSI+3ItIDXa2ldvXSarNxICC191jmkezKDDQ2xTnFgUnVjhh9
VHOc2qQ0o6vyQJtpJZWcaNZ5P98YK3pnna3QQivk/WhHp2hLjq9JShLdRGYSejWO
qyGjDOseWA/4wk7JcS1PedLBQGEUBmZ7Oaj4V/YgyrRqj4EvAPUNju4WdQ10Fw2I
S/Yfo5tMZoySiiNSaXZ3FKO/BX/VPHMU+YNZjUK1ZpR/7CN6pvA1pvuIxJxDXaLL
Xqupw/AkpDOuyBT9/CHRo+de03qFcCpGCi2EBE+OX5RfrllEnnyhib79iqJApDx7
nlXnduKVtCs6gVNJ9gNbhVM6LR6eDtZlhvUODkZskBQL8KvkxjFd6U+URC+JShyl
LK3kTdC1HWxlLJhaSU49e35hwxKnFkeUbBgYKKkRuxTd0j6wthyrcZTCEgKeYiaU
lop3J39Ef258vJ+dirSb96QOPegMvp2hzwmKSN0JuuTW5viKQpCaaaHZypcmg5Pk
98cOW172845b+GOe9vUlC89kiAqKKZKkccLpXqbA8GIGEXX/mF+LTPRmtUsLzaLu
DC1MA/ltNCiUzCLy8ULsjeVdYKmTwSRYhRvFzlPL8JHehiEL7yUU9FUjj/MxNBiy
Z/GO3HlyKrPa8iZbws2lTbYWASxYdgBWdU8j9J4PG5+kcrq6XvwQ5fpaU7MJHoQ5
Ai+KFmQgt2NDpPjeIzhyeO9BVAc1vUiJK6scQoMBa37g7Po1MLtPFpcHvzyrJsnU
ryAC/ZMMGFxQvOeaSt2VM+TruGdElI752lT8PwbafMHYYeVAiifjPzPPHkM7nU9U
VeH5enHkYq3VQ/W4KnOPOytkoIXTAPFq4FUwFhRKD6D7azRuc/6LfP/+4B33fRv9
2ASDbmcGcR5eyW0WH4rrYYER0fU9JfmAjITsifsNAlH1S47tti03YU84IL7WhuRa
fZgzXbfdd+UmTk8i9pwe4SfIPSHNOdyssuOl+ZUZjxWX2lYVnk1FYI4z91aRx3eF
LRPyMzXEX7WAouLiCIeunBjyUiraLWQ19lZXLS83Dg+KQRQ4K8eL5kZqUxb4gj2k
Ar0q50m/Ebfbz2GHNXBbDb6lXbjh6r++Ni/pb/o/bjB4Ai30O7nQ9TZ5FOdeO3LM
7nVfrX8PHX+QGZ6quWzE2ZCkI9MP91yD16T0f8zb5dzoVnOnf7FiGa5ihwYbrsVS
ORnxBTaB8RzR49DjvQvmtyPpj1g6L+BLmg2k8VrrSs/RHHJxGAnhq0TtQrlwdYu2
BoLnW+HCMkN3htsS4PRLgDG3gWw3rz3DweNmS1jr03pNcQAiv5m91UzwHLAARYee
O/aCweAoQ8FuaMsyjpYc7RdzJc6HLurdO86mOX72JJ+DLoFTMdz1ShT/Ko7Hn3DB
8MUrMKzLuNy+2trIS2ar73yNMEMcy6PNRGfosJkPlT0Zu+lYrN0RlJzgXwrRHJUI
pmw0E3I8P0nK+j4TiwAFZWZR/kjvxriRAOu2UZm1ufjQstIE7c3QT6DVUBdS+aS1
Sl64RcCqzeh2BRo8+Lkfxchwq5BLo6IxzDp06CJmZjgC8yRQXmhJun6HuwENrpsf
OHNBUNbBP12DYhs9zGos94jYIDaaMNSmxlkpQ5D4N0l/7VFD+8/O7cmuX4+3GoPZ
HaV+5+44aMNuCZAGTG0kQIDh6uhQY1kxMDK+OJE0+KeosVseNdp558al2XfgZsvt
6P0m+YtGitqNgiicuULuwb0dKj374WMyKi5Y9I68RaNcvMVvOkqs+v8MFwQLHk02
DP7kHL0575tA4Kg7kvR7PGsXsog/mGsSrjzFx0i6LCs3b86uKiOp81gahIgbQbmt
bbxB4rQnVnct7EFbv6bz8WF6ieuyaGLwgCpiZR8aqadaw9Zw4nHGL691If2olPdS
fGDdNA7by9IXolXj4R67HWynPwWIulvXFBXNH9iClRdWIfp8zaoq2ZGIgUoyeDo7
UJ16tcnH+0y7qtPIH9QtRPH3MxyUvoQyVMF1M+VrDEXeh6lCfBeQeGI0gHBxy55K
dUZw0E8KNsr+CU7Fh65MSgvW968IAYpC/ad+rGAiGfit4rSXbeyIdkwEJhy2HK+M
D/XMj42XU23GAcJaBdv38KJQpipHeR73qm7+kJ9NQpgdlS8QRaLfi7sFQbKSH47D
j89hzVShv0ViY//2PTs1dRukfvKtZDbzrdqobdsu1N975/15J7o79U5ZYRGQX4KU
DS0eiEK8kzvokBYWRlNmzHuKcmnwJwiaUUBiaetGwR5w2U/Yf7fggNy9w9QzWCxN
lvU1wknepKqiW2Yznh9LOJZ1GoGAGx27gSY35nzH28eF6dylcHh56l/1Kk1jX13E
4x0iYtFlL49mgwM+u9oZ8zPfQB5p5jMrJN4f6mCbXEBS4E5GZxyGHiGTEjVdK1uq
Qww6B/72aSeETXjYQcxmwOd2tCL1m5hcRMKDqh9kiS3qiLFfV3bf7BhXVmQaRMqx
6ihfaP3VI7FnlIrImIrjatIzIweCUFju3Qslam9rXo/hZ/XJqk479wWZ3QTVXQed
XW/vuwgqODbKsrBBk4IAYx6g8fij5UQXak+TJhTs7rTAxTS3pM3hV3zJjG+3kcrX
Bxe6IEBx6Ba1Lw25J3Bgrf3pSgw6H9h9dIBPu6QDpBIiFHgdWuN033pCjOmVHiEm
RmD6mrXZcLH+SRLiZQEaVd3hygcrPNkYsgLOK2StJ7ZumXCIvmj18MeiBdgO7kno
wleo+RGoWpMSuWnhCtQWq9Q7cBIA0U9TS/xcnPDUcnLlm0zO71rC0FMNGScVvk7q
jh6aSoVP0hT9CayCbTroKasj8xG8waFE1r64A3BI1QQuGPkycPKK7U0Dxq33A6Ou
TfBrK98sEmYgxvVr1RFWMacT11fgIFvB6Dd9lkEbVvPiEs0SCgVYX3sBYQTca/R9
ozG1tR7Rhgt7C6b460FXTNt2FSldK9pR2aDLp7PIsay44qL9aA7tBXeRbRNpaWfm
1kvjqTVB/Ta71rKYS4BhLW/Sfcqe2AdfAP0BowHyZRck6psIReVqPzrpTbfJfGfA
0Lm+/OGyNDkIl0701SdrOi2dl3FvrjAR4gOvj8V3ThRRYLDVm/A/688ahwcqTEOU
SpNQIPkK+U+KpELvuJnGUFaCdnJOwQLOEbcHi8LgQ5WYZSP+3HJHq0skLZb4SpOD
MkqUhunPsp6dRTVt6tdGBzRMvbC9cPJmLALfD26bkXVW3dvf93hdrCXYTslMwNsP
GzJuKvbQE0tM1dAcY5vFuyoPlwX8jvWf8gHMseS5AyTOnY9kRXaPyMMvnLnK+W1D
KZ+k8B8Ww/yWFVDmbevCPpUjXZyqe1zT1Y6jlGW9zUHmPlFNLkS4g0698USyj0CU
o7tBlTQ5CwNqySUnl5QEmqyW4pfXxlbg2idan/L+nqR2bOpvxFtwE5Nlm3tfEAZd
dstvD2IufwvIDFrESLwg1JTA+6pGQmjXCWHatcolSlqRFgLTPvtucoNsJR1GIPu8
rWMpWp4eJzgHN2IbJDMqQmcebSIEoJd0SvCQsO6dLgDVX/NVqIyA3BTItXg27ggW
QXgkMTCvGk7eQD7RhqSrpAzWQ3sB3y+MSC6IoEPDXsDecpoOWn9vJC4zC1tbIvx+
T0o/djov8+Ue8yZGaAp5Ff3bAB/9lVnO1tufqmshemc9SRVjr8StvKGZZzi7P2RU
jMi/WwZlZ3qijsTiBtXC02WpY4tzy3HB/ss/zugvVae5kh1AWn26c2Kio61jDkLH
/uMj6NGGiICDwYgBdHwQZfrNdz2smMSvccSHUVvUQJFj+4/oN8e+tP8tahSlYj5E
JVBFlCtq+R8WplUxBk0nZKqzi08gzgAfw7quLUXmFqj+kXw+xDun1EnwEugfRwec
Ih+hGPnlctUkCKF3FrRsdNZLrguf5U3MW/xHy/VkjgcBgBQpvxt1E+0tAqH9c9cm
UWGcNWrDDICTYvlikAccUWSGir9MFB8M86tQSCb+Lp52tt0MfTQjcqFbk+Vz0Gd6
3e9Ris9kFL9aSVqliqbvfR7aZqKn8aj3TeOgi/Qq6t/Ugyee3jlty69L7miLOtTD
z8I/jAKiYwEWrWp8TzLOQCC1ALfcy9AZe2Cp2R6uySTLu3I2QH9M4t1Vw0PefkHN
+UkJ0X2u1ErgTcT0/QZGCZduhxtzOOBHJsBEAJFFqcM8ZDUaEzmJ4wOzanxfqOAv
FC5zx+ZW+TUsuybmbJ4x2lJcYUVgIB6/VU6f+fFxYIQ01TBxMkxDTHac/h/rYZK4
ELKIbsN/1khLdFTyNk+qXXmALafOjEDfH6RQi0x5S19teg3H8UeAruQygyWEZd4V
ZItFz68EEQIQOpWLoxDgb4CdXvyOJlB02m2wR74OzQfK3hilYH5DXdb0msyhJHyk
U+EEZvxzxRngCbEEno/QGFs+OF/3871E57j5wser89jf3lqWabDjCM72YwyvXi2V
v1p/yw9U7LA1xwSeM2Tq3iO05WkGfaWSe8Zyl2y5dyzSBPB9ja2gUURG3V6/agn/
IVK9pP1AnGf4KAOXAIkt/gdb0loBjNrxPuqaxXcbY7H0JgFUbYm14sVh5IrxsCz0
AGKQbr5RhgehOMp7v1ZLO9nLgeRYPMiDElrZ3zdrlr02gGu1951LX24nsP9kgpfQ
VW9h+f3oae+B0nVf2/WAbDhX5S2AlJW9EZT49F9e/UBOUOM5aDm2KxeuxqioS6Zb
+f2cxc9TtbXdOFdxBQ5Z+m4zIn9X4pofTDd7vElm3LDNcPckDZSKgl6gcWUKRDOW
6jLk+BaGaB7HdCmJfeUdmvfTU3aGiifOg4zQ/iZYnhVPipOn7d+yDQEgxBo74TWf
xosC3au+DcCY61zpZnS41+6WRRqePXjBBtnk07mL64l5uaTfMVBUO/gHRWUJ7DbV
PHH8dTDgAYA7rImeXuLDQW9jJS/hmlVT4HaB5pH66LCJh+qo5bGM7sPlFIZTY5Q/
`pragma protect end_protected
