// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IvzCOFmQBhE9lGZi2gvR4UVN2wXgOAIt39UhQd+QIKXJjulyeC7cffLVVt5zNr3f
sz/vBXhSMXIhzgeoEFogVhEjLULEeNv+LMqCrdeSYamoW/m0I6kjFGHLzSjh0m9g
8uqTjpF1hgpVHxXWy9rP1t0b/DG+VApbb0+u8kvrg94=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19184)
kLbLfLziBG6ed1UJkzxu1WvieZ0hZ1d6eMH7vfwYEIub+5ERv6v0qWeXbO04CUoc
K+yEtm9rQoJCMnvK/Eh3adtEaeJFxC5t+riJp6XVORUj6mWCyPhmZdXCUw3ggLOk
MDdJyGf5H9qY4XIxpmIPqDlJ2ndw/+WSbeu/lcRWTFk3LUHtnO6SFEukDgKUNvab
4fykz1f9coSG5xoD1mIX/I0Q3wMinXQh2SvWei+2JBYMvIxN1F7fhSSEhXCLRXVi
xhV8H3w2RpEfOQ1A72qketDikm5nezVLZwUP1qCdogQzcAbpc11DOyB6ItaJ+nqj
KmBE6VDASQV3B1NwbbUy+kFLJlIe0lsSXAhhKdyrQK71daNKrTwHYn9EhbKCID2L
z7LLpGLFW3DJJGMDy7pSlR7ViJMqoIUzSnpj+7v38SDs8dIlkT56nt2/B9VAVxjz
hSP1PFDSqQTBLObAtdAqE9NCEYrBS3bQwNolbZ6INmYgqaoBVXxGS5fxbHABVgKk
fKRL0yuq7zLyoDEFWCP4Hh16Qe6A1IDkBx1b1vC9xVDIoXYIY3aMzRaxuQO0ftoB
c0twLGWYkF6kSp4F5IyiqAKhMRQgc58bIyhiOVwJBLFmEpB7C/HPnababq+vs9mF
jIADTpTlRcmdbM8HUtO1B8j6Vw4xgyrBnBOG3izj/oZ/f9QACQSheSaNdNldeM+b
OA3LUPC//T2W+wSG7x5szDwGOqfb5T94jOz3t3gmCLhxkfsEzw8wQB1CLLyKV2mF
dteKIKFFsE9JRgMdtV+ZJMkdSdwdPV7QlDcGeyllbwmpfKt96fdaKeP/GCCuC5DS
Wob4Lc5av4zHogT8i/lxn5zgOze4sn9otznIDilUIM/ZmeHAhQl87uHqY48UW/eM
sR5O/GDzXtBOademLk9SbxT6nD33L2qLUoN7Dn6hCfWJucs3Qm7pLaUnrrePULsC
J+pnsVlA5YgPzzrLAxWf6WGCL5Sev+juRoLSr9Bj5R325/KWMJMpVNRJC/csRqIk
ajE0tFXG1Ps9NmPG1J5Lw6znCg0eMO0tZyLdAzO3X+RpI67kwWyN/vTJnvGr78Ut
H5gsrvB0QtcCWRfAE0BhBIZjPmj7i/l8veJIxJS0RbNVIqPEJccP9D1wowOoy8qj
8OyKuO6Na2gN88hT9akZ9YPJAdVIJc7xAiqWqIf+117EmdUF7Hal0FyxALxEGXu9
4dZ15pH/zeYahbSewjfofTMzCh9hv3NEyx3aO6+IuKfzewGNOk00nl+mGKNq5Y63
wDbQHCOJztt2YdjUPYOnmX7Ze7V5AAIxOLTmqAg9O20W+yPxLsAbUsV+kFMjYcWc
bpdC8A6Q6looqQzOw3vQzjQdU9mnJAW+NDE5DSiS5S5d366KTiqdKFSiN3RVlAla
mZCcHfM1fEPjKE9ivj/Vtq4Dni9KseThdHljwqU6lpAPPtWKRVNKbtVFGvB4KBGF
WAEWTNY5Fwt8NRl1nZ5Lc0tMNA3IPWsJnJT+XWm/jVVd6ZAmofiiWQfQq+jyi3Ub
aXot68FAD4VIudpJTsxiqXad8Q1zs+npFN54ypz0GSqtJZQGR/Gt/nEN+emaWBLu
+ksRP7AlN47Ns40LuBgDdL7JlHLUcPwXz9xr183BAN45AWbr1h99+bDV6bA1rymN
qmbXSSjLb2V0Hjg6lSQrdECpaI/JG3dRCVLjpOzAD4LN4m9DjihHDU4d+iI+Wmm4
TF6D+630DjHQC4+GLm7R3Bt9q2/da0iAXYL6pnYySJz58zTyjqp+Eb5s/6/VWNpk
H4jIj3pzdxOBiv+RHRb7MXTsYRnZRIW2BvpP2nSccqWhZ37zyr7TC/63TwiPhDlO
79zaZ1ofaI6XeKlSm9z38m/NLKmnY16BzRdmjZ+05wjfLl5ngIv3FaeYoPNlW6iq
h+xbvJ6uzU83FP+LIURiWH0zwXNs7+mM81hix+1FLaMjTNQLunnfQYoX0IpyVhir
+AakV0OJjWSDLaF/g5IsRDSMyCe/Z0LYwArYdHPZTps49XbTOngFdE+fMNjsox+L
9qA7Y/87FrMGAVbVwgR4on186x7HxCBsvcZmN0licTI5kP4C0Mv2TB1c2BsmFKpP
/kMiZobRw16fY5On5yYu39Z4vrFyzxWaPecobJjF73k0KW1+Q3mw3Nbjy1c43iYP
v40f93a9/rzb2sc2DWPLiH/EXNg8D/t4rcP/8WWw1DIsOs8yPKCojRuBPMkVhn6Z
6l+UcqMrM85H124NqQOOnqihNNSGnrEmOZE3mt9PMqtN/poOmr6DWreTVJVesW+P
5bUfmmLVvmemWWBeOmPS5t8rVlrymtWF8GHkJPbsdxgU0sDHi8VA6T8RcES+6lwb
UY1iA2E/FS9BBRKFucwqfWBA3e1qCIIY7KkDPuSDMCNARBUEPExcwsOQMMyUAlhz
cU1Ekk70RavyMvJogsWH79pdtkndhlP+PLUgf9lNvg2nqKVqd3cSDd0BtzwI3/FE
tOatgigcCUeuABVQ033CtsEgT+7V9lfib5EkPH3NjteGiiT0wP5bH1PQRRtZ7MSS
fQARClGAGcHQmw1a+mdbjMygKqJR7KpmFQJbW6HMtlj8mG5Ajox8Wcg3VXnXeVyF
5Z3EuLcpwKy0BWWUBvBxJ1hBiscyvqiWdnWts6pIEuA22v+lSHHNRlO5XNu084iS
hONHfG0/vAzIdRKoj/ZLEPHd3YHdRjdIfBQE03pFnVb2zaUosMJm1ejrOw61I7hF
yfBD/0AhOjjRlTRCVhRSeQCuBsgSf+7R1NKBdaBxNLDj5Xem68QFGEUI4l1lz5wM
j1k2SDjOYcYhxSYAScZkcsahTBNV7idB0Ixg7IUUf+mXqG7gdxmacpIRaBvpAIR+
y7Z/U4eZVLLieByyFJgL73Gqo9sIXVYkQd2gVjjBiM3gEWuO9reT4kFDYbDc1eTU
B39OBtTQITINQnpCNlyi7YcqXqOBkZR2jekDi5Aq6UKQPrbQ8GkbIW6DHuigoKrh
5gFWD/d/N+5ny4DA7A0YxRRZMH/QrGt9zFNSJ535oU9M7qLvy6bYwG5Q0m79ZtBW
k1KjbQ3mtv8giKUAxdUk2i9e9GrRX1G/7D7L6mElbyhq2LLGCXG/Y4xn+NRB3Hzd
c4exNlDMTtVNX4YJAs/RDEvVPqQjhr/awR3OU5BAH8muABiQQ5/43Sq0P7LWxyqM
fsJcuSrgXyrUbG2jT7y7RYN/A1dL+hCbY6OnwAw8HJfDHG+Wcxqg7zhPR/jHJ5s0
uuEgYqBwZpaYTjuip/8YD95Y9Zw7eDrBn/oG+EOzb7uuTFVDkcDQqFu6A/Aca9Vh
4UxjEP8dawyMCjYdWLRW9cqlNgi5ERGpJkdMsZOXhFRu1ZuwYJFkjfWV/GxGy7zy
NE49HNdoqtS7Ko4/3EgjpNvBbK4/ttwFIP/Wg0SkZEv2odNvZ16rpQdBmMWrs7qg
9Fg+TCgcmcZh+PdLKmvyvwB4DmtFOang6cyQeji/l0I9/Ega35uvnApYooV3cFQB
Se/Xao/BB0YveeaN0kapiN/tgHvdgfsn3xkhpIc0T8ZekGTpp3fk8M1fBFsxGwHL
+hR+deVO9nDj8Hirk94M9mLgXoeab+wjYan+MKIUGJI3W2fGudf29YmXKMda9M5B
4S0NeSwUjG9uvq3vFrPvGeunmZgsRPrZGbqX6B4e0q1g5k3gU1FrFPsS57O4AORC
KQZhMKnXzzGoFIydvIHCcf/x54VDANaup2CstUamrjxyIgyAPfWOucU1DFLZwRkj
zlMfBbEVbVYs8Lpv8X4X16Li74/t2Ihmfsn8kDdHU65xBBYIcdbhAyI7tE9ti4Ql
+nJbpF8yyi7SxXBKKLmEynX7pnGwDqdkXUH/mpG7z2w1ywc+ADAm1wQFpNwim6bW
trFYyTsENb1qOJxlHxfJjhsW1FkjMjTcxVwDw34XOwpIEZPxcENHps5prLOCDd2j
oqml9kt4h+I4FHa8ypCXzlA6Kr+wvGfhT/L17zmZD1tW3sysfNTdDAEJGa/AbUc7
QoZhWdJta0UP9isBV5G0PGrrQWN54ylcHJvuqY5gnxCuBP55/5m/m9YqRWr/PXoO
BH7PCWK0q4QkGKnG0JzN3Pk8fPplJ2Sx57T5Efbp619o1qMPRbHkHy1f/qeNwHO1
i9OTv5D/we0TYsqZTQwDAL7ZE7Y3YROie79wwcoyGRUglTv8D16mMGC90OcDN5qu
1vAl2cMf1nV4A529hxcUIXeTKeAunKWw9v6uBptEAbrm++GJyNUx/1NiXVGVNKZO
FLZ0YlmQYATqOeIVYwcW7XtKOGBxy3+R7vDvMdH88AOPIGKjfbVIv9wX9IG55Yoz
qwkQq8tuatDDeAxdS4Xff/ti9r6Z/M+2jGVealW0l8W4rdn8p+m4EOG5FbwRvJxn
ihe6CBf26P4ubFTV0R9fzWrg/Yq4lJbM7XONn1dhe/PeyzPu/SAX3/ZbftTZZh9R
bd0UaKEalqGGFDqzFwz4e+00vSgSkW6hVCGgRH0LlL4LICPCP5LBTWnGi9oOXjN6
uBuKt7KaZTd6kjZoXdjGJhyVUA0X9lvamTfm02nmyqNzjDLogWtuS7xQTgar2VHr
RLaGUTgIgchcJNBEl+eG5sDCS7sURM2EhEyo1khqBfw5pKGYSOpuADqehBIOuosS
Yzne0kabCCxr5tpCCun2C/TnYaih7e/TtEVW4sIetjsmluEGd8ngQo4fzCS80BhK
A5sNT5LHZMkJK+TkMXMOl8cXncdU0SdfxRnvRaO9+Bc817tRT+Yzon9xrXOuCy2q
Edpjt7Ah58iDs+aVl7ahRsQmkhkA/QXe9K99XWWD2s2twCPViVfgcqWblEWNYVac
Gd9hjO0NvDL6+AcP89QlaTl12NuUj48pt+eDB7OkDSSk9J0orNU9vggxl4qQGjdq
AI3N6IU5m8z++rzxsNFHiXXZmIN43D6TqDoO9ksiybsdBTodWAJljjDrBcbnMb0/
1IFy+pFHhY4sXLBpayTuiogY2CHHEB6NZBccCQCbgsqmXZN66Eu9UbUB5B989lg4
I4RH03bO9LYVdie/JDA+6KqoSEXky3irYtHdJfyfvGkltGxQWB8JCweAR6TUF50Q
kzGmUmvbhdswGGOgSnSOWTCt7VNgQwoxUXHXH9Woy953rkZ0rngsS2yY/DNc6YWX
TGxGwRVw5wF6yHFY7pGnNfNclUpNdW4GAp+N+nqPT9LfuMzNXXJOtYR7rN//zc5g
dBWvBdEo/pgDULKtZeU1n2KeP46tu3v+zNL7ySqIsqwG5CbkGeZ/5Jm+KgTlD7tP
u9tHhYkYeSixTOktCQtKLKx82urKuZh8acv83IWLxZp+6vcAS1hVp/ALRnOSvBMw
c+IgX797akGQZIL+iW3C1T8U1Ys4OjpeTiNcQYbZPl4OIQtwT8dKQRTLQCtVYixp
tQLnGl/sRAy5vbRihl6L3MTAiyQulWM3+Pf/ugc15XrbNQvRRgI3UI2zALaTI5E/
FlBRwgxlIRfBRhTYhHvP6p7sswToppDXtRjD6R7efi3270jNLQ+DTGaoBRyAVHw1
q8AXVgADF5DoYgwttnx2sQ+jExIBmtjZTo5/wJ8+1fS6n7imqOkrhVTP4ES4PMd3
MtTruBo+ytd2nptbBLhFGzR1J8Gd8r904JPKAfSZLOyWCAi5/M5EdIgsdo6X0CbV
hP6Sy0xbfz5MUF3rvrxnJayau2adcJwBpmr+WOuif5DROdnfGWqno30IqSEKs11j
mf+sCtUqL19564fji9drwUFK/6DxUibIV7t/0rAc9YduKLIk7j5fXmtZ2SLQTLN2
1Nrkcxx9x4Ht4h7PyPHE4QK0HZ7k7XYg5QTD9Br5Ig4p+Q9+ykonB/ugkm+5GXnJ
Q9Gu3SJvbOOnU3ZafeST8Emfz0O18M8qINq76Cn9FMuBqxSbxY9a3AkvMWpllr5D
7cqSz8rsqBNpZlGzpOaXOfDkOm1lEC2JHyD0iE6hz004nNj3A5y/NG5B5r+GMjRC
Kz4XiIXIIAoKYPtTVKoOS2tqD9pUkddCh3/sgbC1NrZTDzrLsB0B4iA6eTdBwLLI
IdE5MwgcllYUU/KJbYVdPHsVG+DBCk4dwJ8N+k+L038RhyAfDldiMZlLfN3ophxx
LWfgJCjZusvZzDDqF/ecokVgk53LtDzi7LqZOJtFRC+TUO2Nxv7YWpEp6+eOfXZJ
Mehqouool4DzXhsdFq3pOlzz84GWgOcjkxVvYGgbzO+/F6iZenn4nhm2TtMguz80
1kUCI86utbq/2/vEYraHUQo9Xir9bq2pQrPhFxPxLWzdANREM0xvbkaYwVAnxW7o
hSkPmZCjlSmIc6QrJlq9hUzb5GpY7a7dOc9xWngc00kGxltlx6Qw5QJuUdUeeDef
efJ4mGTO3a/x30iL2S+1rZED36aWsZuwYXDJwfJPSaAa1qLrq6yoiNMT9l/N9+1i
ELvWcL+kVhcdO8qodNJ05fVr+wzondy50LBmOd8J9Hj2PmZM+BK87PphIzOrzazM
eOWr3eY0Bc+4DWrPnz2slOcslv+2h4dTf3FL26+Fr0NrHLrgXsC4xlSZvR2+dHN2
G6sUudrDncQSfQuTTjlF0cGgBqDl22gILhoA9Q9B/X1Q+b4Lw8A4PsPRWSsPFTmD
6TG9DHUR0kUDzhknNIk1vre7hVJV0nauqfeysGdx4eVsJlvrmI/D6UWl7h6MA2sM
qmE+sPZUIwmn+3NZ3oe3kjS3u7M+nRLIi9DChOIrtzGxvvEi+2gMwDgsYJHjgmTB
OGAPSQAciQItxJxdQJYYnLo1SELuK3UVf2fHEfCAhKD10XJ86VbagiWwfdXMgH0q
txSVsa5P9DCJ16SacsEi00kS4OCS/jnXp7ZN+THUgSvwmYBAYJF6D0t1Si5AYsuc
z5hBxAw8Zd4tSG5IYsJzUfVgGuvdJo70+d58vT4l7iLZCchN8fc7qZw5CeU/kiCI
wct6I7yfqQICJK3BzaGATuVSeOFi9FGogvTYcXTrBXncVu0BzjjL3ffe2GWp1Tda
t6TxlDGkFC61bmD12J+sMII1pWRuaOF8NbKia7rd1j9XmATu929KjVJcn/LP4BAg
AX+G40HIOlNZ86tDZCnc4xUd3/VuRcyeaclL9ltawkTSErPoDRJTNF/k8d5pWbcj
yNpkKakxCRYeS+PIwWHjTmtryxWmgOBdsT78R2dTn3yqwcpmIBOowRZE5BsUX/21
cJToBkTpvvC1ZZLNXMnfFy8NBqW0mHFbWrvpDSr6ektnhbPGcgfDz111VTgTXmOB
Mm/43Yvcwb4wgyGt667rmaVxwubfD6CPVFHUsoidTpS43CPAaIWGxwTOo19+CN5F
7uvX75vPSyxnPFrX7M6tIJKdkXaIRlsuqswAOgdqHy+l49m5lw5OHIONka2AK1Pd
eVUZUvpMt+kHix5llCcCYMGJkVgnF5WHhaxUVQRg+gBOfv61K3dRZE2pY1GHaKvI
64M0xjMTrTBagZC4+ZKacwnmJOnHjlYWhGUs/5m0NktQTBgYOIAy8BckfX1y5h9t
itKqGeF2msSkd2ARl7pVII6ob5OevZNGUjNbml08hQpHcwGMZokeN3Pa+bBWFu1+
/R6SqJGQgW5dq2ZisKjfCFSQ40MXlnl0LmUFrJ9SmJpiEqbULf+NGbBfB1qmI8kH
f8xWEv0sj5RFyBAf7MKahMpEBkyE/N3aIrDJ2AFmu8gpGd4rA55Y6Gb+00MlqQzW
PAGIa10zDNopMB440ugth8SV8oerBXEPh6ulosfhYyoy4Nc6gm1+YOiC8HunIr5B
yRvQYtpzCWoldFpsJOM716mmb/XRlvyTsb3jFcfpdj3JnVA7PVi7p9vpGU/t+N0q
hDd4SOSjnWITgbql1eXppESohDNyK3DWGroeYI7e2ABon3XolNvXZ+u7p18yAkSr
ewybep2XCah+r3ZHDJhmhaZfdZvmcLfQf/qCH1Sm9AiwyObXNcccDKRh8pubL6YM
chl1pQX7ZSwsNO7M+LQlFcuj7TX0sUWYSSGtvST79JkDQrYVJHoM++3zKdD+B098
ye6wJHCw+eJalPYtTP5iP2oPohvT/dvmhcuFppK0aWk0mXEtM/T7DCStyWATdeUg
jNKnvbyVNfT9RL//GLl2fClTgqk4T6ryibyQXQ3ClaVbRssycKrqdmQa7l7sncfp
FDhvptebUGe7iQX/Kh/qMPGnYMbbHwRnsWGL80TzehGmwG0M+GTXVXY/1A7L5w8c
U5p7qo+5A7Nka07IF97rOcWRR/0dJUNjxSEPolKolmLy8/M+ZQjtbs5K8nkokAp6
kHL6NOgPDdij6Q/j/64Vp9Zu0t1gT4Xd+dtIzvcCw6zOFinM+FjvCV1nz8FD0WF5
uOunGW3i5izw4jDFTcZoWP4i+weSKjg0BK+9OkeESkmvMXrIpOkkbZErHMnvrVad
WBq+LRO1DErJx2vvOxfV4SzNJxI4qOcVDEKylQPniPrWLp5cS/NZePGVoTKDjQZ2
BMc0ZPcw694LMJSuXDLjkVbQiTGo/FosJKJloN3mwn8mx6WhCzlMBcOFcU7huTAn
oSyrpGBdM120p+a31+dyXKK83UrO4PZYwhqmRIry/Bmsh1B5L+rwi1uWF9wfyC61
mvJNlT46GHpkMJ3iCRHs05IhxqQzz/9UN+VMBnFqmjdfyyQCBQjHFHshIJOkM5Aw
ckDz1O9WyqTT6yXYOQulvoC8ow8IwxQqROe4Rh49K/WaEfCHZQgVkiZQQogdk/Si
soS16ncyVwfS2RaCVWgeZnzZFAUXcLme/ToDZ+afDX6tQPe8TZsZehQ66eclfrh8
1sPYue/BpJR1QM7EVu8pOLSjiIfXH8j6R1poCXGgO9EcK1pPvYShfhUO5tknutIc
dIT3RjQD3xEZ56HnOmP0U4ISMcoA2dtzDTgvS2eyhEJDD+vOwb031hNY97PErGWk
4CZPaV5Qa44VWNPj9pwd2wPai1/KfCTHi9nXfHVmZ9HahY05XNASigCEh+7cBKaz
znIV/l+emCZtGtipBP8V6lPhVhdYMBzbajiKNBZeInwMmM49jdkJQVJcWAU3vFq0
2/WIhJYRWwk5urn6aYijiklPmOHGDAz7Jo+0YZFl3riaek4wUxBHbfNzy2JGq6Du
1Ya3eZm+P4wBE7txMrEFQs4Xcd/uOprxxqaKgKa/Z9hstpLIvPeHbMrTX4aDy02u
lqWU1wqwqQAJh3+BOm34RssUoXF9wcUJhBtrRk+vswzeZUUuXf0f+ouaiDiMS0LM
xEi5iWMKiETzNtD4/RAvYUcGduwlnVx4CTizrimowuaVWnZMnYJifer8hk4YjVT7
YZyfd6OAzX4x7mNiHprvoHMZkw+ffBcmJa5t4zpzBJEvhdzCyqgpo7SKcA4MuMqi
cOh78i/Ov48U+Iziv0IeAAv+4SU9rNhT+0scg/SQX4BtOj1JK80UaAldxc5aC4SA
ThC3eCvsvZ7K9p+3zhzeoGd9cuAd3iB1ihQhwJQQEBtYxXiWFIUX0ZX9gcNDcDOV
6eb6ycf6y4p64mJ7t8z54PbYM/sZpdxdiNUWpS02Bjntdt/jvnLfI6EXOmFNXUx5
RABaNXNBIvwiZYzLv0D3uvZyzjSLXZuR1wmT9zbeGwYz2C0MrR1Ai+FLIFugKoFx
U1njDiIKJeMsEoEq8syr5reVVQ5T1KWpbb1KTqTJau7jabw2IxF12YcSX3lxNU1f
9VGtWSfxgUaNRz/uDx8GhMfmzW7IPb2cbhW3JqtsZBmFCy8X/ZYy+pKZpbddjNAp
zI1flGxdZ++jOjlnPDIlc/6W13KKbRD+xsr+VP41qPUIB30Ltoi1wChz6xET6Xpo
yaPUY0BdNo4cAT+3nUSBGcxY2tzZ16tS2SLGzCTe4rVfYiA1QwaBeazBLTOVt8VJ
LOqfB8tGdvUBivXNvSE0S556WkI8USI1HvPJEg/DNxKhLq0pauJLY836i41kyZvT
KknyK/0KoEL6HpqFxSdwAy9bwmY5l8LfdGLULAXBx+bIxqRn1Dgu5QCZ1UfoWhnB
InnSq7TA296c1rKTMp/8MsTl4kf9OyzrUZCkflcK5pqdTqlCA3Q0NeHFPjIPWrUY
Y55FhzIyPRQtxWlaw09f0voXNmzdBi1DKw9xboqokfNwRiPj757GwuY8vGC2tlY0
owXGNIyh/YV2IWK7kex+pabtaSleGW1JG9Orvex9sA6wmrv2YI2Q9Gw0z7jCtgk6
JlpxWRsdiKdB9HjAsBMi6eil+c0jmu5V9csAJENpMlzJAypJHIuQtNRaa4l5c9i1
2yffb6jCqu7FQf+IC4G8UgNxamVzAFfouq2UKnssf4TnFFfwvcbbFcrkv/El6Fxi
mV0UxbRa0buBQC2c7BR/hv7fNaWDzuDb0k1Kaft2sZgkwV5RcWiHqyrGN4sTFtUr
oPTLdSFioduIoWZo9qg5c0niZpu2O7o03hk1YXcGEVcA59hPo9OaB06aOd3+UNLK
pss+L85ZBV18tftTGu0pygUg0Pt8VcdYmSMd3vHMALNWZN945wV44wmVfEizJ4cp
lPR6UGI/eQE25D2EjqHikMsuNcU2ZQrZsgNHcrIuo5ACQOqwRTF7QRMSHOe+oVfP
p/VotCsxzKkpsmVm1nr8fGMemfXmfrh3hhlgiWh67HtLxdUfj4l8yiOZR5iR9mRf
f2sHmJnaOx4Zxr4HB0Jwv5bPEgYB7Lv2MGvd3xEGRudbrGQvt09e6qybyJ/tCtcf
bbZcp7Oy1xuFwgFJrH4mxstv6bAlTzaweZjkOUG3E44mu1Uu/Y0yCbzBfoRt5Uui
/9cC8rgE7L8L3GXfC0i/v96pvGuY9pyFGMc/4UFEFymPxL1wVwpwW7gUYbYIgaJ4
ZMk0Ffov0OzZZJhrg1K4ciO+tHsr54+xJkvGj9NzzJD3hpubsJSPEohuEyz71dDl
RR32RTutD6oeMND9UF2gX2W40H4TBWkisaN2beP7XH0U5aRv19gw+71pW3nnthVj
oEjZvgXjIYlUcHFyMXxuYAE2PRPwrxwp8nrFGnxTwX2RXc59nO3fqXqskYh/ab7p
j/kmR069xQkE/a0w3p0QxN91WfMM+KUtzKzGYENlCwb9AV9o15qQhnZd6GnGINXo
d1nZrf7TIlDVjGQlL3K5wcmgIHPUxwAGhjvriQron+7ft4J+h8ryBAb8Q4EAAhcs
WDEWPy/a2x+SndmGRRws/MXRjiphy0ZYiUGlfItsXpbyrEOCNHrx6ql3Nw8mFqg3
D3G7hqTQMZUJN9A/UXOJ1p0lhEyC+JEaLynMsMZeyaMN3Fo7t9HYHhF1nrLpMrZ9
oE9l/W+nuoh6U6qTq2+r3A1iHKeTmO5WWOpawvfVjH+q6d+6pf3RSlbbAqWz1me3
Bxqr2edRS/9nZEvpjbz1KL7c52B6othbve1Uz5lc1bBHOagd0fNcrYj7P9BKdise
qi12pjw5F757BPLAwKd9tQzM5mq7OvDOrdze7kdNZ/jHtgEhz3h3QgpT3e+Tc4ya
Xr7vGeuwQcJKucB5Lt1D4GipBrYeAP/4yMS1utOYyC86d+3Fx3AwvcTfvy+C87/u
B+R4fGPmNyI4RKiAZwWkAqk2tE/RteO9qL2XHYohA9M/EJ/4IE7d+liEJEjsWD1f
+pBaHSvEKZYpQ6iVfBdkAJMct+hDC4m6ylFLU+8wBGnvb5Crs70iiqXtNiULz+Lb
ATKVM/N5fo2d1CiT9sHB2rAtz97rCMjZHJuJvg5emPrl8t6i7kJvHZnKlezzr5eG
L1PrSfgHDUxcmy4UmzkEnlevBSzOAQbW4iRMJzaKN2UxNCRDKZm12zFKQcyRLDoO
jj1E/+ct3pUmj7lRAnN7BkpW6fiTY061QFAkVypPeH8UJj2wgCJTWTrKo2xIMsf9
39y59TPUfyq43KTdQNWXEdwKfjJHl3kczUXf6vNpParWN6OlTNXWvuTGCpOtyNxJ
qxuJVVBUcu6WbrHf7QNuz0NGz+niLHXXFN9r9JHhyp24IzZ+Q9y6NzgOBYQWEv1d
yfP7/Hj89d8WDnp3NrbvfpfPk76M6LDh9UmGd0k06PgYVbgAF3pwzmDbbQT7abCW
JksG+L1IgICFKijuj8K46TVZvo8KjUhWOmn9yYyN8IuKQFd35o5xrh1RxgRWGtza
CEoEfXnpGnUo/vLPiFbg+r6AyB9OoXbqnRDS9X9eBtQvVfkEL5vG5/JeVYSGGwCh
ggC1MX2mOMJxpWicz+09VuAb2Sp4CLQ5qEBZKFR0OYwJRuA0agVIUx7/k9ygkO+d
1YvAo7o8+TAfcmw4NUnfXq4PYfVp9odVrlxxUHhNyFKlt3ZDO0b1LBN8QsOd9tRc
S9+PAdSw5nEZNp9KQDE9tpoOdmrkw/MYGpcOt/8jWUovYQE7u3ALbw2oAhqXYa3O
FQOVDTq3qvoUuU5PMbL7iS+POzLN1DY95b2zjZ2IMlEjEVKV6yf5SFfxWOuPOpVW
9C5wetsfCLnD9NjIOq0AqkyNenkkdruz/etQePYZyA6sj8AiV6vCkkj18SZwZQQl
1ckHUMSmtfamvNa+CXs/rmUB4RPiPHY79BAWKFryjWZRX/aV7KD+y7/aZpTIdB/z
y9EDNQ9yc+gkw1el7fETbW2h2h00l9W0E3g83+Jn0nRMoKQtiNAgMCyEMXgF22+e
AXGRPJhESMLECDHucSKNlT09Sj8mSNmkNlxJbNiDD8hbsaiDxDi3Jc9U8l/DzgDe
2oeNWT6vkoq8+MFkVXrx5040WwuPiZ7k1U1hwt3IywOzJI0jO/BW7gv0l4I0mDCt
p7SithxaCm//cGkUyTz7scjLGLMybdDfgz4EqHk0sTX0hMo3o85xXKg0hECBnzcQ
XjZaWY4v/J09BMuwVXVSw6qozs7RpvMBV1OG1xilYPCEB98NuCn5n5N836XjgswK
UOSHyNQRWmdjYF0libTmlduoZXo9poDUrvsm95Gk2B14gSx5WJmuobxK0ntQBEKS
tQiLLkrBW68iqeUvPtUDbdmavcLE1Ca7dyfZKg5OpKIL+Dg+0EWSDA1bY0A/PKi6
u1rIBh/vuw6gWayg+CoLWufnooUylAotQaEkmM11rFxviIt+qN14X574kGHRaADw
OI/RjOo4/mt8pZQdSEcfT0xABNFzWybbZdKM/NrW2R1eNAX+Zd1cIDXSxe0aMH3C
hR12n6eY7J+jC8cASYBlf7B37u/+p1VaozHerj5khBSY9NG5VZX8HEDk12kGwV8f
ccqy0ApBMDbsiMxzpQtulgeQILZFxUIayy58T+NYG7K/0e3hh4h1oLo+FOMd3VfP
egM1M09RL3GARw190hZgRRtoIzmI7RNzWLy9aowDFZA2jLA2WXJoWFMcBrT3Nutc
Q7bB4akDOmy4yc/lM0VE7zQ/LxDsfM8Yfy2IB417Ja+mqIlcrdtMD6k58EJjvAGy
l9G1MIuKhr9VRkvkCNM1RvlgDFuh4o54OXZC1FG3tFk/SiWp7cVhe1jWygghVYIN
oxGcGeM0YP8rBbCfUcL2LSMH6Rx2m6+EWLhl5lR9+sMWGCJ9f4j/4JmMRhNm1gf9
x6Drw9cqriw9mui5xOJr9dzNxNO4OKvZP2qsNi7WNwUecuPN2tcTZC9+ByMjg74F
SX279HuxQcxM0ify/dNV5wLS9JC3oA+ad0pdCZqlSBUwdsNVhDka2uw526fusjTL
uRgR+yi++v01yiItdnw4cMhNFkQS2zqLdIfltxBkhWD2CpTepFbLWGCVMpJLjkrK
QSvujH5Fzw55dDQTH5UW0DsqlRESkVw9b8mtKbctpQHMCgwhIfDPjFd6jIEEESB0
aD2Bl/9K2OnrRKAxIp5sGzQ+73AZmf1vbH4W+evrbTA5cOU0I9xRE9SPq47iDMBW
eqTSGAILpyORxfvupStNsiaPsZbpNZduFYqnlVrqg3iT3aUbajl6KKURcDoHTnnT
LXz/roC1BiYpX38h9b7GDGRVX3zjz158XM/UDGh+no+iOGkH8l4kgM12TO21Owr0
prunoKEcd16MRgFfB5+LRVSlE/VLSVBUr8nFbfDXU+9DM+pyo1yURhQhXHkswbQm
sXfMkOawpNvo7l90LR3Z9mUnc4ebOuak68BQ8YSVQU1pjhIxOT482fYdx2oEesqO
weK90OkjqfREupq/IQINA1keV4zSNTqsk/Buv2Lg92nTwhr5xmumwuufgDIqw5th
lvqkWNd9g1EWHa/bwX+ZOH33r5h8dEunh2Wx8icpjpEFT6C5SyZD24mko4dv+Jnq
uR90iIaPdHdtIXAk10V5AbgLpeH02vWI9x8Y4qPo62lXPHBb5EpbmSaLmgqTCbgK
62jzrNSKXoZWjB3MXGWpT9fVIn2e7eH4guM7KXumua3sp1f6ghXM1/CK77fRlupJ
ghgX5r9OZXQJnph55//tie4oeQB5aqCo1PJyDpqYJ9zVPkVPsoBz5GFOxNolF+tK
hl58N8xRKK6lXzqEhkdIc2VUkTGUVBJJz9VfJzAZA362PX1HwUkXvohtc0abmrUW
Gw1ViISs2dhvqOlM37tAQhEELSNjg++N7kqkJAA6MBduN0H29Dc0Wdh1i68LAoWF
3exZeS6rsDuhOvOFoZYkCkIElttMYgUEHhpWMqJvficeNbpGHRkDoAYpDyPrazeD
qWzNBVFwC5yCTQFOVfRU4yRXQwGhFZnKZnfXdPv7Ff5bFFa7wjDpzO0NNvsHx89I
cUM8oZgw3KZoZETbfHDwMngpYsFkLX/t6KMvUY5D8J4HFEnR3lUOsFLn3EH1GyFB
Zzx+zakis5VSxIMlzhX2csm6/8a+xE2HS5vP8cAzJcQ3mVCRnZgX6sSfAnbw2JWw
hrjdq8u6Nzzvqt9ffRSoQuxsnH/NeqRERhsDJv5WHlpF90+AhowhcAFBiAzVAaN+
ZbYuxHIjQK1sbOifEtziZmx4Z4LhJbisSbLpRQnFNONyQcHZvjhZRu+4tlITdYer
029mEwUD5UgfO/QBWSZneSTNC+FJ3YKc0bxSjjEdLxMHCxrmc3H+jglmP1m69Pl+
IT0fxJZPfq/V9N5CEaANmkpIxB6WlGIQvOn27RG1AUqWKwXJXxGr5gPXvZtUVLdN
PqCAGHhM0WsUpzlA7RedrZtF31oS4JHeSRO7APFO/qzKJVqx9en4uFTSDhvlofUV
PSRXnmwuxN1nZUFUQ71fX1Z+rC5bhgSM1NOqoIZYsSjx/MvOipElrk8HJ+27jfhC
8SyyNPteWa2lYECdSFjZLZHK/A5+4UcpUXbEhUISCA3aupqstXohbyE0OH0ZPOsB
/sBuNllJjXWCB72Z3dE8H8YSGPasA4ar2un+1sdqfSzozSp9mMW6M3GU93eJzlLe
x/BmNHjMK1MLGfanw9UeayE0ToLMBfGuWwEZLCAl5LcusmMzIepGvR5NkiEjgKxQ
MwFXfvwXjRilDq5oSlKMHhwSb5cegmg5XE91V27vPw3p3+mvJccBkxE589wh6GZA
rE+1WRLAh1JYR6YXWFx4L9nWavfgibnH0Bezt0HKWtZMsr4OYd/K3uUFuLKn729W
V+1fka0cetY8UtJD9ZK7MDLjaLGKm1EN/v4g33qKZkGK0iniAzaXCh2oxmWx+Y2p
VXlmCNCck8zfbPtaxgoaOUpzw6NKj19i48PnNZ2p09PyMd7cRHptPxtmp+VNrZla
pYxZUDz2FYWzh8qRFEo14fv2V8jVPRdAnQNjCu9nZHnW7ESiZL8qCqImgkSxNnn9
UAhEyf3lLNmi82gqgTjsmKVUsJmNpUv7Ll9PrvxRyDicf9luh0yie+IFnpH4Naht
29fg8al6SYR1K5gDAOqnnmRe5HUkCRbiJP+3QibSHE6IBUddUe43bp6UXEGeyCA/
gM9ibylpM9v/gqOSinX19BMTdN61x7/PUyYL9rR1ZP/GfeU+ZQYLgfAzgZGB5I/b
bvL62+lVmlhdsypJgiDH73GFUPuq4y0MoIHnH2dOg4bgCFcaVdYKVjnzLJ3eGnEf
WA6S1fOZ9fYHusSq5sPKPC8wrmyqRBuiW3BQaxY1fWPozObjlqq4eSlhV964/0cp
0G60jwHM0DDFj3Ix9Zn3FwIzfVvzcJOSB/aPEbJI49AehpigzvBVru7/uK/5InrP
3SDl6SJXarLABK/Yb4jvZPiqVs29XMq2/Sdt2LGZIA/A0b4yeDs6rnosbQ6+oAjO
IIZYIO8d0zq7FQSnxpxVWiBAcBqHMdTeosnAKxsIX7juC1mbiQGEjg0u9XLckjHT
yjdqParY8nz+Pa/+CbNHOt2EuyEmNxHLSeWcCmTd9Wel5uePLYwlyeB71IVM4t0g
pSTXnWlBpuKIJVComXpplmm93Z+oODhiwywloIjzXsksJfOEQaoFVGqcZONKdo8X
CnbjdlBz7NIrFpRbFc5nABLInw0acQHsxIIkgrTSDrKivPotW/J1leJ0XHHZ24+u
ykMPnQRt2mrlquXlkCVSp6zQleuTCJPtZtZmXJmFwYNcy51MpbXHbnOD2VYuU5n4
HAJFx1hxiomIGIpcgGDUtRmdPfLcJcINqapFXigJg98q+w3G+XjpUlS0KXh5goPR
o+TKFyB82L5xNJM961dV+Pasba1tegoYzS/SLxOdeOHYSasKwRseV1oqKjN00I9s
4mK7uR1t85q7ZITBeKgXZhNLUPvjL5ItDsjMLdGR9jzp9r2xGwpRb+7Zr8Ri5zCw
E2vKJULBDq11OUp37B+7k3Z8A8KOWg0BPrtdmEJx78wLg0rYKldm2KSKZYF6Uj+v
tNvkp6Zq2MzhsJneYy70ITwzGm+jKqMetCnGDW303uJaOXVB1S2T78j7gkx+BfxU
Nwyv0Fz4GGukC4BBs+zuk7nbl0lPmh+/StamYO+jZCRDxnAOG9Pi43GM3a/FkXxQ
FogVDrzFoY3DPrHQbFw0k8usnf3rUNAIG36Tet+6rqSoTp9pZEMAbdllPLRyCBWv
hjbWo7JNxXSDHNT6xo/+866+kywvR7cvPijheD+X53Ach/vgu4lNmvrCnAUHbxev
wtBDldS1tuWcdVy3TQ4eXJp4WAxCMh8hT1DeR3TVrWDNQC4718gItsgYLXZQHTIf
LM47sNXMfbwMIQn0DPI6dTxR9XtoYiCZMrz0Y0pvC9eWAv7foCGYRjIxxDtZnBIZ
1X3o2OhQCvxyunIQtRt24F/IWnx5FgDN6urzPW3ndarAPk/WcVT38rvLGQNsf+sq
ImG36iJGQuHXY71kntdy0/BDxZhWMnGwPdrZi4eskdmHqvXc+JQPIxJaQDOeOEpW
a6GHSfUlro9/N0jm997R3bMlLDW7bp047W3RswHY+Bebk3/rP3/OcybOvUXuqmWq
4Fu4wOW8eMtHDMkSL3o1lNMxGbqmn4NWmgSMzCwMqcQWAKnHRfR5R3b8f7iRNyC8
BcNOwFgPfUFzCVHwEFV+6wZInCAyqyygkykDrzbE5VlCVZg9jedAM9lpVzddBY3E
jH/7Os15s+JBgGZvDsjMTpZbhLKHWLiHRc1f74VFTsp1YNCXULHcQDmHYdtN6BeY
JbYlp8+y+nzxvw1ktcXkw6w1mPsSIq0mO0j82LLonh7gUH9ViXjXSOFaJYIgvNDJ
P6QZdvMjxHYnWaRA5tIEjhhxgLAL5enXwlUAApqvxQlCjItoNnLdldD8DtkLfsjS
BGj9GEfNP3bcCbWcp6gPFQN+PbyJ8tff/wgC2Wn+SKBGnZPZvBhsdfVtQUXWEbHN
OXMvR6O4+K83/5hctI4i1ofOulfK5brmIWa6Iqya24N+kZfWS38ZAIIPr3yNO2x3
TyDSZ1TVtFUdLXFzUHuIy+iauBMtWXWfYqVkYaLfKKyF+ItWCJwuvf1Wg9RWh8iV
Dc3D7PgIQoN8fhqrfKpVWKbxN6kSohdudtbzw5AVL+Oja6HSkOLGblejSvkZaJkl
gZXB+O6Zj/c130Zd6WdutIJt/1G7rBFboVgPfWehH2MSKRTe/kx7O7su9DgUds0N
Puvo+q7dqRxIkkTWBfWJoJSR3Gd0NfbMLEHHSoM/n/aENN/xon5QRjwI9G89QRw0
pHiUSVb8ql1Jw6ikkM8N7N3rPjWDkE7eTdmAjAVmDszCd5s5YspdOlT8AfAsJFYP
UeYWqTxQpjbdJfDzrPiEBNehG8Fh1xsDAH7CdIE0VuW19gDH3ATTq7WhcEjP6cdj
PV0Pudk88WuxZwEBWg2flY/Qlr3qROjXFW+rrV/9mGnkPY5P/IF/UMX+ruOeDI7X
3hdGAmO3srmkbnXTzK+w//azyl6wwrI090br3HcoGFVGoiw6e8O5deUaW50+VX6K
c+/bQ0lDKpy1hD5tvq0O9hlmKD1AVFpPbGYo4kxFJXVbS6EyuKFwnx88l3uNDUKW
/tzHO7TQI6rHWY5Edgx4RwlEyVGbH89JzebNRe3AS1zuuoHGVbhCSOuwm3/nxkis
qF3tL2L8+hHibl+leHNxZbzF+ry53y7HTdUgu6xcDxAq7fUeZ4kSDsWjsK9ugKcn
WTOIauZ0sbQ6V28r1neHN5lJiOw93/ClqfY8mN3+eXY5QlXz7K06dpfP8Xp9E5cb
J0EKy7a6W8t4hsFr3VA8jMUNRhT/Cbax6Kz+0WkVL8dOvVn4/4Zq36GP3Zfnx3Zf
JaBcf14y7XlVhVT2/pZCeXyEllUIZBX6oWswLwHHWy6DxrccZDuUrThvGXtub7GS
pfk31wwB/euyUgWY+u3oRr6RSh70UZRudNpiyyLM7gbGItx0VQ/m4ZO6NHWyEats
HzE/lTstKV1yfLk1HkJfD3I1D2GmyaRSLHIVJM97Kq1Hs/d43VrBzLiICDcA7rk2
/dHexLiz3+ggaZYcSBd0UC1bEhkar9+xFp5uEMi24ehlGgd+K+ned+9/USvQbgfM
6W7FDJeio9Js9PURpk/mTe0MAJ+DMfiliPVIAJlHpwNU/y5aUHXc8wQ5FbwAT5YY
+XncDdpu+tOajY4Aqh7nDeEGlj6qrgkPc3zXc2xHtLzSsBKyfpDw9nkOSCLWylQf
/7yoh7OQ15zKiEj8h99Gin84dWEoqisDiCUMu0yHPCxl9FP1luk3Oot9chaomP48
9J6/zlTYxhtllmNobve4/NPvuUp2erfBPeqAc83TppIch7lGEzmG0GinzboZLKhq
dpC2L5vIXO1YwkD+yPkMJOalgqMo+g9K9/hgezg6hYp3OAX92uJzu0Ig6an1VyAt
eg5t5EczI4xtQkU3QX6SnJWBj09gPjA0QfNxicEprwnVb2qeKRbcUHALh+pgh5gC
WagkMVKzdqXrtxL2L4qA9yWQawo91egmTKop3ZAzmIvhYrmbg8zt+yG7BBKnHTCh
s1vXRCRlHic7JPvY8PIECPeozZgC5pyqIxGTd4OUn/er8S/u6P4TCKIhjdQyx1vM
TFOx6GamiH+DvzOb0JCIKFXwucG8gNOegF8y4y46U1MxkxI7wVBbfI8FPNNuq59b
qy0cpj54QDwXTBHXr52lFV1QKLm7XoPBsGJ3I1/XZtTJ5RIfOs7AWgHPLT3t0e6X
k2BXN8s7VaJKavdRJT+Q0g9z4oXazes9/MOmxIIK6U7z/LoQLEpVVDiSMyhHC0uP
3sgONTrgdlp/2iLTKTbAy/fpwb/bnKT71hFVV1x3ITtlhNQrW81hnnajsfgvbmRX
Da70GcdRUMwDQTNd6I9f1dgYWfipis17RwUWxwnhzBtELXdtlUPY681Jw9a8XOw6
lMG6wg475FMg5+xiGpfrKTQN6iDsFxukcFuYev1tDzLwzbQmZTpmsfFOweblZRt2
Y/ctZk1adkMbKYkS/aaeiFCEQi7UjTCpA5rgDgYkFYAqaCvX4dzNZ2u39Q/7X4mi
0xscpG9rcXVGUZNjgs3g/wrS2qoIDDD6sN+c0Ewz5uD+NR0T7Eu/IUxY57QYoQYt
YomTaYi6YkUu7XRN5jlvBDT4nziqUHVbW0+9uu6XjYJrVlfB6iFCEFikoxDstfwB
roAPhvaqVcTzlKcyrHpE7HYJxpPFw7fBpSP0TvJ3CO6JawGu84mOO2IvF4KYJs0x
EBm22qFairKZFaGyrxGHahxx1NPiJG4m/93evU2mxEYZkQYz4kwLP4sj+2TkKMmO
4kPgWwjXoHcd8MK0yl78C8bu3rGMhGB74t36S8LqeKzyl6p9afo8GR04oIbDOFKV
I+diRUwv/Wzyed5XqZogcFcA1bvI4RxjxkrGUQ5f020x7UUzd7o2xhKDXZvPTOiZ
5retcRdk/9WGxN7SEoacxNIOHiRNox3tLjjq4hj41iv7AyeKHvQq4qIz4HcG2MhC
Z9L48O6FV/SvlJ4ijkWqJ44B71uTjL6WUIhmwgIfYvjz4Xzj1bmfVxxheoXL7AF6
OBKgtMmauWSc59T+Y1Y7USfFLuGuJOYtudeS6uST8B1zJedvdFgSunh3aKEjf4YV
ajKV0Xj6RVwO0I3ZGtpGt5ftR18L1jOcYvg9+T4Cjuzmaq+ZZTAc2N9H4pdh7zho
mY3I1pidmN4LHCm56O2XSw+vCfrmdZw7GRec61l/pQttbqS1SxTgXIoeeUVH9XPX
LYtB5qANRXrQYkm1Q0fwoRk7LLUovmU3hi52wZgxFyq1jIy7CHkx0rLHF7mDLR6S
ol7xv8abreEiyNzIg9ZettTAj3lxQsc423OZKseeURm4rv5/Jox6GlZNaA5b9Nqi
U0F8J7f4FSb3iKqxRM/+P6OKP8RXjETLHYjx+UZuXv9Pe8TLInX3PYJBIyVct5k/
UknGvScABIdlMGnclPC+LHfmamsOjT/SnGN/6mCRUzXfdQGXu54Qnf8GGiZmSEHU
YUv/f4pNUA7GtzFdjtBS+CPVOZa7YxCJY4egOpHdecxsU08LqzuQ2RRCIzG3FnI1
Vr7a5+HLeg/hCbazl6d28EDzLXugzFkGyr1/Ul2AkdcGs496mJEh6woOz9O+VKzO
ot4oTg7JOkf+fttois90skpJ7IxVKTBqlfhplFi7/BLW5hkOAqs0hTyQtL3qMmZ0
PhF/6ec+/JF7Pmz/C9FTYjLZfhzmPRKdWMNZJN3RTRR8qZUR6DsODQTLnyB8i87T
zjk4oOAWDTDORB03U2ELSNj4Xv3fameMufK3AIkxLTGtsvM5ItZElbzhKDclv4GT
WYoGWj4xH7BhUOeHGeodPXpUeTm2pGIpQZCw0/REJj4wAyKXu+pdxMei4RT+R0ME
17DRmdIcGIO5jfUJnQEBV6321WFaKqNRwjj1L+MnC1hDArwC8eUQxRhz4Z68DNGl
9F8SW6fyutipzpjlnPt8qzOvDNZ02nDwe50HCv0Th2bz6Iqpyed3SwHDKDSgEc9Z
x87vfFMwhCiaNkR/o84ZwFGccaF43wPTwaLhlaeXpkCIJYhn3BBr2/dViJG9NUw0
AJDAv3B+3PbsheMfhJnZqIQv2ij6aJsMuZkof4mlvwF6gx+sVFQj3TnSPzdIOC47
aagYCzXIycMxWs8MHMQ8AxYB1dYVmkVWMAb0PW8o2OchtB2R7PR+ndhLJh06SNiY
NaRGdKenrW4rAgVi5pIDNO5PfFx/cFsi4QOslhKBuV2ud0TqnaglCE1yokm4gFDN
OSXvh6mH/oG6kUziBxhSQZH1Wj9ACoaVEMOn05Hw1NllDjYiB++gE8kBs/wp5zOP
MfkvongFkwY55spcELfBVo5cLDFe2GdVbvggor2IVT3nMMSvm9E4dfhq1TYXJsF1
EVRkZzSk3m+6I40gPQpN5ztGNUOGO4uBvnOSDfxwWRXxst8bmM2K/dPHnzrQIfaB
SLfq3TH4vUfd7z4SpkNNMRfLP0Ww7fF2ZAQeP1dFZpYXaK94O1ZLalg0GtIA0Yk8
WaXY83BjcG6XG07vFw2HPQML57mvV7UhmlQTG5lgEoa8qPhhclJbrozFGMvNdWf6
zWfR43CFUh14oRzRGCZeGF7QO9jaOodCkIFh8F6Zor3Uvn03KVRieEIXZWwQeIG3
1TIHdVx2Gbo5Au6uIu5/AlPNiJ1ighNkaxQqVZU8T+mzsmPR3kq30cF0XzE4OG5M
2rTP06Uu12q/rRw85DJEn7Y3TC0+Vz2N0IaS+JrI7ibwX74PEvjWncFgM9JzIbFB
7LAvAMp7WpPDSgkYFm+neRoRlP7qyeMOouQsTgEKZvJ/42ebAGz6K83DhXbTpiJs
ld323iXED47zac+BmS5lzPRNHNCi14ngiQGjm9HglhpH7AOz5EW48rQfvUkAMNt+
Q8D4lxi9c6kzR3O96ZNOvmenZRGeky4AUIwPofEvl3gN7W/kUQx9HBefq6+wz5js
KZPOUCMoUxVy2lkskz3XJRWw5CtYxhl12G92yIJY/SIPi0RFWFiQO8AddYCHA1vh
EI5S05SThuQkISVGSlWCfX93FdSc69VyTcpuxaO1t5kKcSQUu0jObWvXfLKbR7Ag
d8yn+WI8n5GgVLR+7KGhrnZQezsIeVXGuR1wgYmwuC2zCBM88x9ahh/kfk7dW+0h
S4GQ3CzzZpNRA1R48YSjxxxBCc+8WY69NVsOlSzU6sqcKq2QfN3+mUA/QlwtVcVS
xPHayyYZUxK6euf5nDTGrlHp8a/YMg0cbyEhax9YfNq7NVwcPQFiTF2K6sECcl4t
CJANDl7uw2cRmsRlWsbuUco8PQQI0ljoxxU7IFSzrc1QPvAz4loimqmOJAzaQTxY
EhqbrATcZl1K6YZVyTNfh/GK2zox1PLqWM/+V6VMAV7yFaZLyIeTUhINianrhl/g
GxcrZjHCAZYHSpyz+d77X+kSSNpULYO/ItNSb3+m3cmjrRVy/Ke2Q/McSjTNfHHK
6fgpfuT9dgmJLF7c8NMQKoRnd35zG0M9foiO+MprCR69lpAoZK4hn4yocb7m4IuI
ztOO8KtAwEdvXgepV306w6gZz61TmyciwyFWnltxd3XHIxUhySEja5Hyr8mqpvSq
tP7GA57Qc8SuLteUN6QLA84PIGEjJmfrxR4pwIBjVrHW+aUzUDD/IpAMND1ireT8
ZYfwRkGqahDNFeSxtFnMnwtTlOZRcWFinhJ/iTGOKr2wSQCo92auISKBOAZ/ZTaA
YnXpsRElWGGvvHcmvlPdxvoT4Bk7IaLlT+yhLu3Vz0Q/U6bT9Dua2atnmoIn1Znv
b+DsLDRF244BEL8hobQ/KDilgo2tMZJbKnVJpbUvxV86K01TTo033FDNbH/efis6
t3ARDsnvRCRwb+oV4TFYJkec/kDHoOHb0wPYBqw6km1c77eAlArKDUIV+PeqalDS
l6C3FSp5zXJNqC/QVVGvoD5HJFAXUdxzkC9yEeikBQUzdfG7bW6cD1qDIgM8isX7
j11ULjM63I/miMibMIDmz8182nRb4p5Y2glsI877K+dupdZecm/j3gL+vzoWj16q
rRkCsu1oySY/2Msa8A8N/AEvr/u7Bkwf3NNpwC3xhJxSWLr9NaoYn8NhB0vtGYZ2
ZY3HEsSWqWJ0ncuDIw7oZxXJeGskNKnyERfhyPu6J6xG2E/vvIrBuyfKbCrZQ9hC
vsUGWvhmFl0LuVOfUBvak2RvxOeozKYkkoDa5dA0z/lXxq254iZDuw/odd6iIkz0
eRWEY0wsuG9fiYIfWQJan4oLoVkImC+9jke+vMPT2Br9dgr+ix4H3NgnyABSImSq
+c6XgjrIoakAMfzO2sWvFhAP4JJ/XFFeqAtxmTfIC1rHYcJtUgj/PSGaHRHw7Rfj
+yZHX4+CCi8c1+ZKYbetbzyRh9dBiufC3fTmp6ddEZRihzeRcx/6Enp79xPk2L0x
YgazQxz6wgGrC/dQiImKp0mtGGxOlrqwYqWhJI180aRthI3ot2vbwZHrcclhLDK1
AG8q219dmlYlkQfcH/n6kEJTjIQfk/ZzujHUTNKxdCV0o2065j0VCnOttFbLaxp4
0Ea5g6Bk4+hH3Rz8MtkaeKDPVLxaSbuDwZeDrDXHzxFZrjLzvL6Te/qRAPA3IhyF
0/0PutHO1WLq1mU+Xl+bDdB08mwgzT0kYc+f++F6hRA4CbWf6jF48zH993WahCEG
0hCHTglcxx5htkBjqjk43BSbZqXWqIOIhhnSwuaEMSdGbxc6vFhLCfEE/k1hkNOR
tqUBfnBZZj9/bhA1+B97bReGVIQjHDdMJaPTeSVm9Y44VhjJFL9pNCX5mkBt5yZO
uO6x6mJQxAl+U2mA922af3Debfke0rD62JW627fTzxgTj+uYVwg51SEB0tebiXz/
fRHdhE4WHyP0+/zDyWY3H+Ep06zxb3D2QLC2UOsBtKvV18hWax2mTCFn4Bs7+fOA
DkE9hAiqc9q/jcKDSL2QNKmdv8tit8+edciDt7LVBrpFgptjmKasYHN5mqM6m9NF
zPjcexcjDdL4oF6BYLzPsAZpNMVcdSaFu8QHBF3nXSr3zqRKMplm49mLg6fl5b4c
Gr/LssSAPLC786f2dPRJwG/bxuyWY/xvkhkrZ6HTOZe1SE7VBeWZrHBVsxc40ujA
6j32qDOxjm1AkwL4GpV/F/w1WftpTakdJvFXNt25ySKCGUlK4wtacfS54mXXagsi
PZv5u6x120xDx4+mOP8jTo0GRzpOS7b0hqwz0gL34k6LOH1v0YTcqv/AtF/ugAf6
YRojLboABED9OSP+O31thBqrZHnt/DkwvmQ9aBrft4zy4UtMTaFWqUTr9ObHv029
Tm0B19ZPE4yq4JgjvE6jnGSMamkiYPg29b0wy6xToe1GqxrCMhD4OYa//C05cYtg
Y4yLIBbSbXuEGk8q4X0fRotDyH7E9dBKy48ATwUvjmurTW5HuEHEZ/UmmIfbUm2d
RqLLo5rw0OxnytqHijfK/epd2HqVSIWGWW+asr7lyRSgNpSsf/jDzJ9kwYjvSVo0
DZ4CKUpprA5MhUqnHg2EgRPDc6ktkENxv1jZNqwTKUFzymweIJ6cuPjtaCEafrDP
iABj1F5u8Biw8IYfNwQ/zXw6Gb24WeXOu3qT6Qhnu5S9mugO7Em/69tK8qXafJQ+
sU1k7iOGERafafzKuHao9q135931FC3Z9usDJtJ/v2WI3FR3hC+jWl2PGUhogG9U
/dpKqZT5Lyg57hni9WlzIicSRSM12VITTZsoEVrw67XUDWiwRcCG6XjSHL8inqwc
fr6DfpvedDWtOqOEDzAZRjWOjv6lAucCApd1YG3o2TnBsSpP2osakohhCbYa1QZC
tJWEX32cCIG9fPr3rWs9+Y0xowxBeQONOtEmgY/yll1CFUEgJD2G9ykUPptAfYcw
4VGyTUsIZThwk3nG0MOrHjwL/kqTyxL+ejg10y/6x+nWZ+nJyClJLWQXYXxLjuFZ
Ud2Ng3ilszQB/JQpfl0JyvaCCBUAd0DwL9IBEmRwUTiR730u089yyO7WY612LoFK
7Wy4iLp/Yusp/jrvkzbZgDCjay7GK8WsJPyrRLXimJVQzdav3PQDJm9jHg2EZk6d
1Ce/4gudC9isWB/TR5oTaIYcKHgdWLQU4hD/+xo9iKTxnDLWCKaA9+c4G6aLv08k
fb9eA9gbbskxxto7A1eQKWXECb5Q1fOH27H2kT7oQi5s0lJl6Ulm0JgNGYn1Bz0r
SDR7pMbkwHGDyYgSjmZoSljQkyF5nbCm3/nKamCQ8lU=
`pragma protect end_protected
