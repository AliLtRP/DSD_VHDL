// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:27 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EMC1F7I15BK8DFWKsbIoHSowgv06N6CKKUGKCAXeZW7fjPkBniQR1Yq8OHhyH7AO
U3rltp6N4Ok8O9oDaLRtCZ73IYqQvsvN/9xKy+vttcnH7sZgOA3nwHPsAWLSoucY
quKUkNyAUf08jrhMXDNdqIx/pgiEbJG+2w5Iv3F+3Xk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 52880)
cyULvM2h7JJKQEw9D8IjnG+7R/YiKjmTtKd+ovajqw86Ul60RAQtST1OHqzFnFKc
FyEIDaUUBDcRTGH+rv6g66E73h2zwsLZnfyKafMrBFOdGtIRpgwWCtNvBDMgS9mJ
G8hUyfISB3WHsq18cVG5XaERvNsXlYXPOAmnqPO75YBK8pM9aS+lj6NjgUbMHNgL
7Xz33gw23Y+Q5eDfANIFTslXA2wfyJz0HpR9c0Tvl2bYrF9fjJz1vyCnpVhBPwLH
AlM6poIrz/LGcuyP+z40lXpL/SnvzPgm09vzu2kUKiHeAd7CKgptH5XI0G74fr1v
UkdUd0JhASyaQVvKdOLDAH8tNK3M22n+CtRn8zmxQ7Q24RxQTl9qD39yrOYXPbgi
i5H6sKoLs7JoEQSVNccMMhd0jWp4F5mxMg1rUyJay3NzhdVfW979IIpQY5OtpRBf
PI58mn6TOTwcE4FhzUUMa8vOx77lxV41xocqz11c8yEiigmMA2mvjcYMqI6pft3D
u0iRulHaEG7DXDi/uMgfMeH63yJROkWWthfeBMRqVSjQqZnYICVfezXhidAL7aq9
yN1wrky+UpEuDS9PoUGYhE/nwRBDhxxi6zWPJdvdzOp/mZ5QpYdLMLpniaYQirRR
kQWQhZGhIDSUqvQSxYwIXoK2BF5NuHeUWODxFmQCvNmvXqrBEj+GkTgxW9yGrarg
Rrzl2NwqcSzrHBtu0FvAyEuLKXP2oO4kaZrGrYfVNrcYABX73LWONAF0rqeqvelu
cIJAaFzzwGmPB8reoDpnEiPCBt/fQV0aV5txGltt1+TWG3/rr6zZRLc1eq7MYSmk
UbcX/rhQdi+anKr8I3OUv5VELtOIDscfyYq4eoJHwcX8EBH0kc+YS87af6ViLI6y
SFCUAWdpW5FZXeEpv4nsxIfdrP3MZCboe7tztxOOt1OvMFjnPBtplCotn8yYos5Y
o6b3Ch143vx89GmRDlXyHnj7qpsr3GcqmbH3NXctDKj93olH6br1dkAdHyqk6WWo
//RwGV16m69f++d3CSVcnZ2SGgGB3n93aiaxPfGaD3wdzn+zGN4xGiWP0qxdq/KA
eJEx7PynD1BtWC+CNjOxc2tj41xp8yDde3cuycu9FYc7q9MRBsEVFIc7Eps681yp
bLD7yeFuSOV3Oi7PIrDcXfmGp7wBB8n+jNq4J1cVP+14YPkQ3/X403P+prGpN3Dy
NMgfZU5Ejju1igMV5LZqcVCs+1JGLa2QzPKhugioW5J65NgfQsy6mHcR4QLWGVN8
P8DLogSPpRwc5L7W9+HH0b6dAFbYcslYSOqZf4wc+GcTP2ww/bbg7CsmPFv7M8r9
51+lEAzYr0oufi4nI3l7E+sT198BWX0c0komPZ6Jfh+cdSTLuWeHbJUmI5xQYUg9
4zIeGBQyBv3FvyauaNA0sonyw/rRzMHGPVZKRD3rKZNqQtKFq9UOKvyY9w4fC50z
4MeX7y5mGVvbsKzRnyqoC02uJvN6cLeWUhxGiaZPH7AMTCp9DrtbD7kj1tXwqGn/
uX8qN20QTzG1Jwuc0SxWPlbRmnwAfTJJcTsu4gbcGNeweuj8Wl0n8mD4B+/qQVWH
TojV5mHku0ZEzpGfS29IY4C9pYaf1AKe2A2WbbnijWVACmEYOBOWFgX26OJaTfgR
bGBCTIKkwLQcok66ar6q3Cs3lgqc5+s/xN0Ff5/nNa+dh2uEg8TRzDFiqrf0arF1
VlYsDFfSRZvos07JsNQDLlPdT8+JDLogBXp5a07n2m5ZAAixz4UYRgQhL8uYO/3J
480ayc/rrnIyaO3FL2GDDI1ZuQ96F8abS5K1HUCP9b14Ry8LSLYj2X1JQlczja8x
74wipBAP4Xlm0vZr66pKNHOe0+vdewCo8A6a4SOtiTKkx4cGo3H6VPQlu3FQu+l0
k4266R54iOQf9MbBbDJB8WuvBvfQ5bWxCsgD90XQioEpMrWX3IwecWehXg4ramU/
cDRFSeYr3ZUTQZHvqltWe3KhXLZ71UdFuyxqkMrG5PbUBB8Z+D6SS4FOIh6pr+EC
ew3Ejehml9UI1Fxoy9Cp0aLKQiRQ0kXXZqMQwlYlXfX+BIdSt7gAeghyoQvM2Jrz
+5H1vJZI+5agN+b6Q8nkrKwxrFgkd2n13OG9atzg+SZY/1ckuNjOV0k5bqYBTpfx
5kQzB1fPryrdexkbjSLt00GjLoy3wxSc4zo3qXNOIjOwxxIrAOCJM/TSMsZi2T33
4hWbv0rfgmsKykbVeH6W60iXjBTFRFU5vtBDN7dt4sA6cmEHCzhJLGrpb8ZUh2Kw
NDyDPvqKB7RP7OwezIlaB3G62Q4kDVcbVlr9l3AWqVvkF/1nIwUEAmx/lROZ8fgk
HIraSMqwDnjg3MZsYopdpCEokbFf0qhk/DcpW+q1aAfgcu39h3uKPXg9X6043RYN
nAMn5NpVtyBv/q+6e3MQ4laTbRwkiGw7te4vUJSiK4bOyCy1OJ3aCJP6Tx3+wGlN
9C0h47JPI//XUUy8Su2flu388ridn1kAe9OTV/9Z4MxdgRjtYg5kdqOLlwa0w+rc
mwMDrWobD0eymd+85qL8CJMnSpr3wcw5S4bIzvvRVNFFYtsPTp5JzER2CWDE68Lv
d0vaf74QjPXiIEGFcBJ51ZIzZJHokjUEhKTdH7U3hJbOR3n9d6OQ0BfKDHjfKGpK
lluUc9hSXo5Al4uIDBPvR4e2geDKoGcrlxiZzZm8Ra5KfXZ1CFRVZupW9JmVBZUe
HVyjAeik9RGr+yOdLzyszhqGBq0yMCeG1+DpLf5dEwSr4yexSiKkyp1MMAsEXUlU
zgNXv2sdbBsuYYB133WgJNefgpzaj5dTVcAKC99OUMkjrcSXKryuJNQP8Y7y88hh
bCFG0MgB6lAKC69TY+PPrA9DM0gdM6r2dVKvJKjXofUCQlNBhe0qibfwZ8miUeaL
Kspc2f5EXDxt1TfSN9V697RgkyQ23jUZmbfHZ0V9p0o2TcErEGQZ1E2c9IgIWqK0
Rm7LzWDIBwGo9kJi6DHvXDUmY0DKYFxDQUrBt+nfjT7XrJfwBzpEUkmi4PrMDZRQ
+TYbe2rOrA8ZuLvqr8xnKQ+OsEzMXJFBBSwFGT2r7d+2fj2uu8y65ykibX+Aegkj
hxukqPlDJKU+WmMwCIG205S+NQ5kJWsyL8FSG3q9bTratKEXHV5oONBhMldohl+d
T97W4W6NyFvF0fQJmAt5acD9MhAsxzhUELyakonq2MvE8adTTiLHnobRmFLT5JtN
nbF/gJiQSWwezk1f4OGnmJ3ojIWObZiAp+03AnJgPVsbTjAixhxkEffbe9JPdt7X
ze1h0Aktb1evwA1/1Fn7CJezT2dJSCujRqkmP5xot6bKh3dlkOHjoypYS94bPkDc
O8kDBgpuXy2lWcLQOZhUpfN1ZTiClUbG450d9xjtODP5lrGIavwHE+CcITHzMps/
+OL5vTI1XwYadmga7aOQVDoe0tcaQ/Qm48KWBPKJW5NfcOoCO91hBab5RYA/SsC5
6Q4yLostcA5sokaH+dqrST1md7ySNEoiBbYqs+pn8RaC1N/mLHBYvdxJPD9m7Ma8
P+2BaBeNN5VqrWVTyhyTsKi9QR3ajvUDM+WeCYl6vPKWrKfiPArBX/gamLAQn2LL
ElTn7DeqCZ0Ii3i9E2EiOXRZFoNbacPyr7G1l+v6bmIzdH6r9vUtGJyiCHEU96cc
iLBdqfPMV6H8eJDx51YV17XaZELuTXyf1FhPSooAsWFcXoZLnyjZaXAyDbsYJbdQ
5eV+4hFConZGrxV4I1aJgYL1o2jPT22achEWjCxE3iBThme1DC0ajLO+CWu8gGJD
T9XoSPghZA40qrgWdHM6yfQ8khMt29adH1q46tAhyTlLu2QX4Xt53VwXNanfrTqc
rG1FbEc410m3RNABtflZRpiSKjq6IV3lrfdqlYwzOue1vIz+RiZWjg1zSixgS58c
wLlToEft8zwfZ8cV0l8tFBGkgGiclWyuZqSdyIKt8UCGJRW1DAG4VBaZqziK8CQv
NuvGxmOyFF8baUsK8rffO9+sIXuL1pW4ViTTGDcWi6PA9tMsY1dm4Rbcyz7JkN6L
pCPmxaym1fjVxA7oqDgfzCQEKvWvig54psuFLhQEkAT/+YwLI7/BKWqeqkQ1Mfl6
evj8KdxXm9cEQ6L6d49EtuZ0nFNKYsBg0sFtQZhARr/M2euLmk586qLoPTthi4/Y
jbhZ45JSfJ8L9CWc0I0KOAsqVVjXGHd5RtkJmoVp4tkpxR8Hpl5CBv9e0SKLNkYv
jPjPhxBhtm1xT6/fj61TL+cw1FECoka7XHmzgVagOroYk3mhyQqMVVWESSi9Pwib
w6SyVr7hYX7kxJCHHk92FEY79FbuDpgI62xP09CXHtjfZkgmrHUJhd1Ovq/rrkKE
ZLMdB6TPuI3JHzbSdxHCgLuhRlM702lqQg5SVsokwBSVO8GpsJmQRJYhFwAzMV7T
ZX0pXNWKEMbhChstrVt66BCtTgtqV235XpNY23Q3hF1CNIzaTyfqdeB1ZMTm14ew
da1ycFhw3hkOZGWwidK3NKdFLY7C5HeAo89mwTDPcWtXyK4oI1TAl9OMWSgKLnAQ
yS4LjDT2mop+OOsdH3ox6DYSYp30MfmKr9SnPi9xIIXi72zieH5iVJEudpE69+93
vlnCQgebpMKWCMdcbBuqSCPXswIDfbaEh0DznzNc5fl2NuhKZk1xwPiObD4zlKY8
yzk4yrENkAG29ugPBMeHZPKT9SFq/wR3IDrgKqi/2AIGeMiLXNGEwY1LTP1gEeD+
iew+Pct6Y7nb5NCRe5NBMNhDvXKYQjFZOUwStrNx8ybjXQigQ18/8ZDoeTe0IzQN
zfkWjWj7/rCadK9J4rIC2arLcl6bpnFCQB+XUbvhVUd2zPFMBy62Ac7yjmd3twcj
3OFUeYVvHDX0H82yX/478ynTRyGoVE5lqDj3zu9RRtCkSQeNZToRzFssCQ2xipgw
wXetNtrFAx3vF86RJ3WgLb/FmZR7AvwNxjSb2Mi0q3CQ0VjGOWLJj8Db5LEC+Hmm
ExWpuCP0/hde5kCY00/NonKvQ7MpvvA22PVHBF3BYAyqMQ4KwtlHXPDDm8OINuvM
N9onqJjlypNh+6GB4YfYRJOztfzsbobbb5nFrqmyKzZ8Xtvs2r3yeVrtrvhO3gm2
zZkdmGf8uZva7938qTsY4vMUlm16lL0VMJXTOEjxo+X/k1J3IWnQQofT/iw90OK5
lAkA5sUbJpYQ4yTnXa8lHP9xYewBRzvMm3zl54b1AdAwqLGXKyjC5OiMg6XeiFGn
IEIO3qHfwMVdX0FVmzZDPudRiBXF793ibxA8X5aMcEDHDlKsAgDQ4dMreYx/9tB6
T7JMhqfvcQZB9AdTud1FWYrHv13mzwawM/AEEJ9RAUt/4r0I2/xxQ6ZORYk7tbGg
2kuxSt9LsoOziNMzmC6EB8nDE5YP+9mNz0Lbp3dJa9lUHxepUTpm1a97C+1Ha0ME
NBUAL/y/dABNeIWFgQGcKr0Z7MnP4m18aVqi2HDiRMKX7ar7CoJbPfAAIeTVEj3Q
gj2Rop6tVR+IJ/xA/sXb/Cx8dxG/6ooUhSyuY3cD+EY0sA5Jz15s43ln5YOyZKgi
CJ1c+mx2Z+2aPaqxayloFXPLMaZJN/0pZZcj3iSLqvohL1D/xMCfojMCyiQDlqGc
gwwgCqm9KPRIxUoepVWB8tFEQypRn+/wBT5aFyhcKegPDZTI+STqxNhiw8YZkGaH
m5+Fy0E5NWR7E0ehoL6tbr5D/h5l0yG2v8At70MeKMQTcggUuOua3zyDne7LUz9P
D02DR+CXbiwy6LECAlgRZvwpxKSAdFJ+NoVE+EJK7dxwM5hU+vNNqyEDK6c6y4YA
BRf493VvOcPoRRVUmeJzRVcdroFKzJZfJWh2tYanq7ZTz57XjxoaBCkeHFUdDRhi
vDJxavfPI+z2sCbFMXaL3PtXBQiHzcGqsvJtxISFdohR4CME5CZFg/Rgawf2eZKV
1MatgoLBmXjKcDbrBkc4s6yrNlXqSsir0QB2LJdYiDv6LAOsB07wIZUa7cmQ98N3
KA8lLb0YQCHQY3X4ApMvjMmdAxYJfDtqf2q/Otkv5RgPt1diQlqJLqYT3uJQXyeP
G78rMz2B+3tK+SZ5c9YXfa5GGJ4HaruaB1c0R0z/gSeY8J0xLRhAqlUdwpa2lBN6
pFS8l7dmbrxjJ6BmNO06TQlv61sANpE+cJHtykwRkGew09hq8EqDg8dB6dT1P0uZ
6sW2HE3ttFqi/dSp37pl2MZKZnrh5odFRFKFLMIyjlyQg7b2oWec4+45JJ77ikg/
VxMS66oldM0jgzQlPhs7IaXECuavf/EsklOkSf/u+lYR3O4MzIuyGn9vvt7UJP7W
tDnRuvOLRb5cDfHx3XcecJlX71h1flhYGlevTGsvRrp2By0w+uKV2bsM+IB/0QtJ
5yna/HAS+aqLTba0+0gPtus7vr5/tHviJmD8l3ESZWiw6bLpmayTAOVEw/gE+W6Y
rFW/O7KuGmiLZ9L9ywUgQ6lIPx/+zGQD5aGBAWR/82tokF/xWiTZp3/RXMaYGXGk
vtGTvfT233SsYtCYPSubwuxKtp+JoR8QEVVoDQJmrOOUnly89/pIBmE0DtDFsUjx
lmBK+eyau2Q+whrXiIVPkagFral9d75pYo+Z0wLF/9Qx9d1JxJFXw7fcBDOFGa+0
FZRHTDgM5h3KF6Nuh4ZjQDOjbm0BDO/yclXA4pZXTlmR54CrmY7wvpCUN3UmKDhW
EAM0cBtpnMBPOs21oogdNCq9rFTOKpDrFZPokiy6ENDZGmiOTIpaW69JSoejgxCc
0jXoEuMkD2hvLZr6+NsrYcGhjZgaIXYa3Ait+cfMRcSoNH1mFO4T4C5VU8lmQbEW
pOc+BVPeALB3BEjLS1vi9s25jF3oxTimtZsf+ylpPK6V5F4lYBt0ScDdr6N27GbT
uiO+D8Xb/t1KoBPmczp4Ra+eHIS+v9V6X8ffhBhZf4OYcu1BfJRX6nZ1D4FQDFeG
AkzywDl3BjeNXR2eUemgZTabWZHgizGcnDLt1nXC++oJ0rB8dlf/9cqeVLYeCDjD
xI0N87TkiwUAhp7uWyb4or7VeC84sd2dWxdnRVTG8wV8OSBDuBAfKVCg+WuDdsZP
xYDnEOkXAvtbQZjvKqF+d1FZ2Jm4oqumNZR9+fKBm/ZCI7s6OCebQ9zhuSUEdqRK
0Yvi79+Zuc7uoA9llKNIrCLigz+IV+/hO+nP97AUOT7oOnR6iUTJ6Mn3Bt87ZFQr
dBDp/QwiED6CUjLy1/B0FKJ9BNJmBVVwaC8Kr3dIESxEdcLzeoebO7ikZM1o/umb
m+VMqjRwAGf0frSMMM82lfYwsZq2IdQEZba//hUw6k8zExPGkLpyjue0tPVlh61Q
jg1KCYn0D/cwoJlAOqVkybxDLtshYkXqUXECQDfiPGJBubgyin3JvQfxYQdoQhA6
IYmoBwaJoldUsoKlENsYUD3IrDJMbnqtdQfszDp5EON6sP19YNNEMq8zr3c6kTg+
DTCgM8hQnKv3tn0jDnCvhP5maC19XkJ7VqFyR1n3pPRyYdn6uHAHZ8W2cSRSLvu1
tcxnmlr5WCztwXI/nn8k4QrLkw5xt1Z08CYu/Uttx1uYZH/Pxd5PjX0tWfgQdtM9
/EAGZ2+IoUQdrOXJZH1QXui1mTxihWx5Gkf9qJ/xOEqz/VNwVJdYPOO5HP3FPcfx
GrYGBy8ZFnHTH1IB2+orT8NoFmQaNPXsJKRI9aIpoiu8Yl73DdDCsvzZyP+HWw58
TmMqLBeu0jy30sn8eKslzdw+ZWsOM3ayYu+Kpl+AoUp9sNHmbmboEMcW4qno9n4V
EBluasoFh0XbiIiRGTmNEqiefW61ky+l239W0DWtzTTOsvBl92WzZ8eOnFHneINX
/tCu8caqopCX0VGRZ9OJndN140t/i/4gEmsJdVMY1MmcYXYq+MTkMQrTDvs0s4io
q5jlLraApob17n8M37FM49LVO0poJ8GgSsdl8L5TBJcUAYFcPr0A3F1ZC0bcgzOa
WCgdPo++18HyKkdeTZebh9NQQl8jKqzF3w6FZgJsdPNqLePRnYinaTqiW+YlGTHe
SfkIynX5iFWOgv7S7WV8DpTOBHzshnRwF8DABkSDSufKJ+mCNpSC+YJ/ePKl44bZ
9clV2x4BKtBjNEP4OBrr+p3TKfLtHjTRIUxCA9GgwRal7kIX+6mEKMJd1ZgjHtkc
LC6xY4Qu6cMkvCbtgVvYxsRS+i3DmuZ9YDqm9hu7Bahi3JwJmvq4c500x6wryeHI
U4fli7WyPGjDJoHrRD/awGnWYnvMbDWBqfXiIfSQxJPZuv+m6wc0rxHZSbTgZ0HH
4k5okon3b8QoHPn68n7CJa1wiphiyuIUQIotrYHf9Cxys1z2mv0hs46e05JLnpdb
Ik61GL+DXrKau9+rqMDPqFbocyZDy9sYZfFssFM0UmalRETDCuWCs2ngVKwHx1mR
ZacP5isM/5Ualu885mmAcMNHSUyzElWNp41yGau3Pkj4U4GDYVxI1L+5bJ18Dgza
8Th0CgiB4CKeNFaDSmWLmH75K0lZFcJAbINs7otGmA/lot7hRJaPJPCaP/xCszXe
y0mRohOXMg0Pq9RTNSNfzVt7nOg0n9Vkzh/7Gkyc+LR5q+xBytlIDb1eywoHupY6
zA011dGkdZAfQh07Itwve0teGygrVZactYPDaw5m0DnQQrRE26rk24GTa1sh9Vpw
NRpFSayzDSg2zpRY5zgLRQ4YH3hVcEAxK5Jp6G9U3TBeh3rSMnshiNwb4Gk4v3/W
u7Kxr7ZDc911CnBTJSIqQ0RR/WplxtdlrCFGIG6rDa2QRLcBgt/Jh3mgXdH6r62g
ERulRgF3dGEKdW1dV89TbeMsvkCicgl9q2Otrmtndj+ztvMhgla/NKBxmxUB+Iqa
bbUrAHB9SInXE4Of7/AnaEJ6yBjSbUw6TgQQEZI0uvYQx90/tHgvT0A5WfnhT4yV
0udkmAsnB2XL5kiqIXeXhWNfHJJc+H1jdSKNzgSKCsK4V1PWzBsCp/b18Yq6g7kL
erMRoLblSAQGgXxUf4W/fiWlGNixbpCvl+CClQ6dGjg72CEcwt2Yq87qvsk/oafA
1Uzfas6FzpMq6sFjGIcB3czCc2/QKIhyrP3GUtvUYbdkk8JuGXYxdq/OU2Ik2Os7
EwA9mOAyUpI5tjZN+LMchdb63GTWNU1yjzx4QfE6HGxlQzWQOcLuVDjZA/HtNYiR
TWSXd2dgoRjNFKvi56RyaJg6N1qPL7lMx4bdF2ZyRlOszmln6V48p3avnTOnt0tO
IEWW1OzqfePhxN4QTu9GxXajJKZFC5+zV7o6qIMAjpEE1vyC2IpNk9vj+2ROOFke
p+ZafvngwuVWdJtfnxT44ZsN1xNuu+2JFEvFBdTzswCEpoTV272xwETfUOtUkY/N
54193bFg2Wk7t7aKFJxnfkQ/byKkKi/XbmYQL3kEoWuw8cN9UZbJMTfTeppWOhqc
qH0NwtTOsBv8dGYRwfgb4RgA37Jp7RKl8W6UiulESP6Qb7Gq2YdDpBj2fQ70A/hx
u+kTDstoE5ec/EVzBKl3fkYOI71ofFyW0E9YF/NZfVBuhXIQ7Pzb5duDHYXJDvP8
kjucC1DKC4SnaItZ959frtDy1A85AQb9hPYNH22vTKUV4sFSGVc1izf16KLH3MgE
GBXfCE1RKXVz/JhkdvctyevOJIq77lBzSJ5Ct6144rOxH3Y72caRkm6xZ3yQcFI6
+8G+u10PRwZoDhrGuU8vW1s17YMfu3S+E2ZdrqHBbfr5jX5RjpuE4qBwGxEWeKvV
mtsFnDW2du1Z8jL0UqNk2J0PPAMDTsSiQGUanU2r9RqqJG+OsjpIZLVsMZ9e1waE
Hnm8en6gmwcsIuNvO5FVUQBaMxYt8N9WlE6Ies/WF/TEPv5WlPiKRd54yJ0V93om
qNZPdE3IwoD7PH0rTIu3mLi0CipFFjLwfvNC85FxfEo+2rIHysZNisRUEvDoytJB
8boN6TQkc38S4Ug+/Q5aqq0uOj4RMH04eR1W4RDTMHuZlwJ6F3WM7xRU38zDLqNd
p4Fi4hV41BsnKAOm878ZNm490GFz/zvfNwB+bKE3XomxIJ7xYRqrlEhkmoJW2z/j
IoIlRTem2A5RHeCEv+ruMg80zWcF2VpRPx9t32D+RvWc2xgNp4SqunWNJ+gUqGJI
j+kP276GpbeXKA3WPzvDMLSi/KPBSP6qHwTZ0bJdFv2/HuL/63SBD6HTz9RvAD4d
QqjLiCWl7DzBSthc9AFUZ1wYKz/Yqpr7sXX8NWKcdjQFmYZnhWR0vp6dX19GOatn
V6LZ5nFWx4h4ZNC346d0FQMcksNAe7lZuEdqQn3v7MX+BbixJX+8cMDhuk0B2U27
zBttYy/8qFxC773YP5ZWhVbZ0N3Z6/zI7w1VC/Gjju62n/CG5n4by3m4WIIuE08W
33LkiguT3c9dPgROsN3n5XLwY9lG2fwZUpG3rnC7IMeDwK+D8bnzomI2Pj2mBoaE
81AE5bjxfjW7k8yTQobgOfk3HBI49VYXugaV0OtZzlV450vJDiL7UmaOS34/rD20
mvCRZab2ZTD1F3tsGrruiiXIaya3a6kyQM4Y9Xku430+CgxCrCjjWU2AhZktAxoh
zx//n82b9ar+cJxdUcnLRfvtilb8ZWq/47sodOrEmyUv4vR/VDT0uoki5jQQjaIE
ARo4G1whfHID805+UI0/YS7C659KcsoDSXODjez23/VahHJ/cKy0Snz238mW4M1r
cIdeGp0knLZS3IpDV87mjt/h+/S5pfsyUKuLurGZGrNHMEd/9ZqbwyZgDe0pfX9E
Q1VA6q3WRvFtCunLkWt6XYC7Q5QD/FJRjxvVDx8XOtobxJ1YQvlYkZEgqmBgZhTU
oCXwQjF6uNCiRyzhLsfTU+L1i+OsEoxEWDUyCyVp+7szjl8R8KN26CPdeYplCuLu
WLVvTAYsRjCsM9mTtYZPiTKNAtvdQpO/NlJuh5a40n1OIblAudHfArXjCxcMNiQB
er2P9tsMF1IbmmdwzcWJsT8M8BsMyti0q9VSqgpvrrWwxX1dTuGQQDfzuI7JwBva
SSdjhEZ/7DhpOOPTtFJyXM7+LToZ74xnj7HBlFRe+dXLuXekCLszLqAJLVnitka/
sL7yzW/9KwRD60WbB9/2QXomutNliQZpMLHqJl+qF//GmDUKmUnvbbWYfPOBZLet
ZsXxeEiB52/bF1ABg4zg/7aMwLjPbKP2fJoD6Mp9uDlPWKWzOpEavcHjN/dcAZLJ
Yw0AVssjuCIevtuU7eiwnJ+1CluUZ6rfsmXYmwahsBkllicletGWuAtJmeFRAd9u
pjMMGuRvYIqzExzAuuPo83soQNhX3nbspIa5jvzxEKgqsl8HAR8MfMOfTmcb80SX
viCpeGptNtBziCLw8cA4uYwfUnRnCLrzshI8sivKZsm9M8M7QV0qz3txmIIyy73y
YTHl1MVLGpodrVC29rgSvtQrqXU20ewvtTB/QbeUXH37PwZMw/aWpbtO6xys0ynW
6hf26nO01HDYobH2Lbn5KI6XHgY5JEXmAKznbNkz10VQ9ZJFyiodwodwwI7dRrm7
KAhC7LHakNV9e6hRJ/jSlEZb65f9Pgr9yA/IiqGnVl24jOEud88yRyXYen6YTnef
ykR/vG/GqY/P27ZyFT8TdrTLot51dq3krQTV0o7ZpY5ThzHcxeE7M5YoJwouvnFT
Jjpy+kzR8Q5hOy3eASWdlmW9RA/1XHeR95Q4WuTkimiwnng1sxcGri54KAVGtyP8
JGuP7bZljVN8vaKECNN54gx6KhGtODwuj5w4NP9XJE36iMRgN00D12cB+0cRYD4s
vnEuifRUvcTQDplj4Exb+x2Jwpw31sa5jV9oXKB8V1o8IAe6eKG+YI+mGkd0s2zE
LFE0aSoXyUfPpVdG88oxJA0YkjTmZGaN92PayhrzsoXj0Up/X53zWTYF4++FyFHK
EjeqVH+Ciy+63gdj2bOP109iVdJOriSqbfLHnAxRtoFe1gsz3L5FhjlGjn3JV69+
g5SficOIwwhomO4SEaLMxxQAIr9ZuUU/XRx5bmtpWR6LQj6YAoE4gxzYJgbV7pxQ
y8pRqge4hZTsxX4EJTk8rJfkOaBaEdWaWy9+RwfBPA5RgNkgGIM6EqLHRVvTXQOh
asCVqjZiffg2N/NmG3k+8iLLR9uNboPw23QJuwnp4Q53hjwRaupKBT4l+QkyR0kE
5LcOOBsCRKtv9qVOxuc5rCAPD5YRz+xoqbbYvONqRttF05IcWmWUGFL54WVQ57y4
ED1qSbz9cdV4KUH75Cp3iAu3Ykl8c+/TjZfwO6rbyNMAT+TFcSY9re+bMh+7k/9D
qpXrSqGJvWgsSaGgiQK3Q6UNrQeC5lgvBbw9t9RE53WQNROy3+hMKsWCxa+FIO5Z
NZFJa91YqFgHfBtm/Uqltc8NfnSjZLO5QVs8+92M+eiANXaEkFKQgSK8oD8wWTg8
mqKm/QGiIj6nkBCVJ4NszNTsUpJZPLa08s29sm2XOQXJGa+1aGRQQc57zjTfHeIV
obRPb80qatKqEjkVDGk+xdM+drFjUoTyx9cIbeScqj4rhePlx3YA2XxubFCfohPj
9um9aIJHT95O7w5nsV420nEf1HjEBGm/++GBFC09MXLEBZsCV2jB7eYOJPch34Kq
ylalpnYAvn2wmtM7dcfvtnrz8xDgy3lgoW2On7/6P8vXWhgFqR5teSADszaEe7mI
4+fCTYMFl2ivRrXfpy+ek5nJJAsb1avNBUNvmWahh4t1PtIYcChQiCF7COs/31nf
bHfZWZIYmhBc/5GehXs5yc9hCLn6SgOWbEa2YUTRORlZdlwCxNdR8nHSS2gXGdPL
hHdQDrw9iRXemnJQx6qy5Zu0SQNaNGkvua/ArG6uyzdBS0u9IPjOifjX6qnDdIB3
k1uyYJTYpNwA4yOIogEctLV/My4M+khS49Syl0MAWlShhq+gwQREC3NF5hL0/lzC
nlfXIbFG5/rzdUnAqir8onSc1nDH9Qz72ycHWvTZo61uhdxbNV7BGMkYq3ydsund
9bzdFw+OQTAX6BbGsoZ69taShpk13UEEVc/gKOcWIhhqJfXCzmY1itoDazAgcRZp
XkgR48rclwb1CEkGKl+gZxPeOrXfDZBDuXEYYtv0g4PlnJGVnx1e5lPTKsyQAu1F
TVRZNOk3RGwdfe9BfyfysKnYP5O+nkj8sju4H0z4F1GpvyJZmZHIDW5veDuZNwTA
V/2Lu1nDzfSQffum2HMEnvg8UbY8not6Gr4RVMnVvbCDEDkAWBgnMgmDm6C5IspE
3zydLph/RD1YA/D6eywD40z+xKH48x5qN/pBv1WANztRN7no9GpZzlVW7eadQYql
dAqqp5XRfLwxHJKfoa8DHDVusEM1WsinLRcmGMReP/uR1OotZ5HnzQoDk2Tk5qaq
bjyFGqyKD97+ebm1EUWdUYxB5XRS7tqkmrM9xExAVlCRDymE/hflH1jFvY5K2jk1
zHXH30A3b5g/ho9V566jp0nHN8m5U6HHpjlyWqobEJoFT4k/0HQ0UGdA7E1IzyFj
0aIFIFCX9LZsXCwz7KSVtrFVrC/oBwoef6pjP1TuTyQ/SM1C381SWEpNUn2+zSA6
Jva73S58QwTexzrYvletwNGtNrL/g+QgT8T/SpVKcmNDhvsyT5mQct7DIsRM1RLT
7qkx+mG1RTfJkOUVT8CivC+pQp0wNZkaB9HKqNT5kkoT5rEJecAGLEDMxtE6nJ8C
02wYvMppGByOB+NgI3yK52gwJ6qVKZHSv/1NVBQYFrOkvWL+BV3t6T7pXNzNSpWl
l84NnjKybICMf+Mg4egZH6SuIgpcA803h+wOQrEUwvfilT/rqZV+zqEwX6fQ1rOS
VCny01rFC0jICNjuXuwLOG6U+uE4qepzdwj+BW8LEazSGNv+3rL1SM3HVhK8UN+U
OVG9BhinRkiTb9CrITSmGYQMwS3UCDNAlwFMtnWYn8SEislOI4IdNEy6maQPgHB3
C4wKtKUp4vmo1a/IWN99nGzEMo42mYMhJ+oScgBZO3m4yoWvhHIMxsFfH/ipVo1S
t6S901PzY7MXpPnffxEBxH0uCSjeHFkJRh5QaJLw4jiN2DZBpg9opLK+MliQe6J+
BwYiNqYII6xlioIbmQ8Gk6GuV4BGTDte8K19G4MbYnsHPXGcR4y65aEJdOA2//72
IEIGfuKaYUQOVCrMdbmFCAJ0sy+tokD1t3kvdaPlkk/IpNS1SQDuZIXE+hFDGjj6
GeZ9tq2Zh+vqgo1Tc9jWn3nId1K/zD6DCxXR7iFOFIm0fb7LeNck7qW1JS76Wc0N
yk2bwQtpl3y8bXDxZh5rc55YkEu3ugjglnYmJSkHmUT/EEDy+/4WRofr6PJr5rLS
Hdia2qy3lHczKY7WUmL6HC6GbDFIDtB+1/OtalJTO2no7cTYVuEXWT945rf5dFTw
zxytzqvk3OkEw8q7DSV9cWQ/cxCt7QF2r9XfQYi0GckOfkvtGzesMcI5R/ANROfr
bRLcNpYsNhFfgPjNKMS1ssnb/KF9DtWoNjh/JZ4G+8lm2NF913PDFhIvotjUyyEJ
OePeEMYyOFaWt7/d6EIResc0z/n8F2AnXdwp2hR3dNY8mJ3xzATjooMykahXDofw
YEVtxv3nYPzkpUL6j8lshCWs1jN27o+9mbfFsy4VW9/1O83/z1If9dtnWi/t+W6T
YiA5RYdqZ+LsEjcWsmS5XdLU81yR28gbuuo0ZXLIrvpxdvp9+h9Iq9aweocYyv23
p6V2iJECGb+GhdQB3wNXsDDObormvE4Hl4j0l2KC7UA0n8+LnyZCfA81QO/CozCU
FCgQcTXN4xmdZIQVQriDMgVcxUNv7LU6crTnrxhWYdDR+7jxuhSEJGUyvv0dnaGJ
mYrJcP22cGSxw02APHiwY+JLZwakqwNSyjX3YE2Ifs+dzypq8iMg9B4O/Ut2qR8S
VjOJS/1A3s1CRa2tN+WAfVQIJpG6eyiKMgfS/YNtQKLHEnSWAr8W11yJmdSZOwDS
1/540fSiBRdn4dOaJfVAPyHa/8hFDy3jWajTz1Tg4Uw0lWlFp0qo8LtLMB2Q63v/
g41szqXwll1zB1UAI3F1uickroBOa6i69hWqgqc0Fs0kXdZT+2Li7IA6BOt7KPAj
ir9KCqT8BmpXXqsWcpgJ0yznUkxsq2loHFU/BVyWQ1gl6bgA5169Gtv+UvoP++Xl
dN5qjFMD9DAZJMcrpBuVPtfHzf1/RnWTwIgrIDRUO/+Uya4/p4699ufwXWpry+bf
EpyhwODIwFsFkZShyTDrGjIaIwnSyYDOfeOsWNH365y+AG76Ufu/R79jQQTc1CMo
EgtnwDORs41j6aejgdCItX0WIYXzpudqjjXG6HIzRIKxnqd48ELzQDjey/tIQqim
VENr0eeLyF6NT2Uho3x2F8y4qYKhU2Cmm7b+8xCEGXi1mqbEnHKP7fB4cqOaFSir
TKCKqIORsqjAZvAIthPvELus1p7KNNMg/9LYIHNP89P8RIA1ym1WFfg5XziiPIvf
BFGiJLSDbGUlObDNRu4bs55LmyOwpU/KnO9YmhpWiAg3ICiRRL+XnWXT9d0g6nGI
0YquzeiVN1/fasW3irfKingAnpIcJi6BXnaXgbcHs5OI1rw5cZtFfLgN/2Ad2/0K
ctXU64dFPXySTSUSNQa58tyC2+MGMZKW7vNSmtXSTEypxb0nAKPmWgoqScGGoxnL
1a6dntUj2CBXEeF6W1DUnLOeRA181doQ6aljKAwh6DBT5YKMZkT08TMsWmQ+DwoK
u9sFSf59dk3hHvd+BE1EpVSzd48qx6u6KYfIePI+mKK9PJhSEQ3uyEK5Z4OSS3Yi
SjULWAg3ppJslBotRHboAsn1NFDRnYsg1Sf+uFKtyJ/Rl6abrGVrv5OUUJgPACjY
QdngQJH/J0h/omXlmMmWkPBTS4ImijDtH8Q4jjWvE4RfBVR6lVbDJrWLHXmyiwrb
NxTqiRSNLpdG26ae+NOiIHPsnxvP2rDQ6ygAylYDMpUWraxv2Lv0iXS/Fbsv9eZr
bUDSHPWbtI689S21I9QwQ/N+vPkIk6MCJrxoVVs0FyKKQXZw5FRV/tQZjGpVoXVW
Yc3OwOG435oaDIVzujHRwKVG2qbsG6SUZVVvUwitTmGtk/44NXQS2OJZlrSdaJXi
85EGLHNf0NGSVJPjs2ltwm6fa6Zt5QYQJe8V/t/hBtKDk9BqFjsVIm3I8AlkFamK
uB0mDU0Ao/0n1dYZNgv2Y0YroOOWt+SXr6fZ+0+4j1mhlktbyQGlBgfPkvla/Urc
HTnBUm6x5CghiFs7L0TjQywmh8NAW4N/fGq3r7ABkTG1MgvNm2/3RWgoaS7jMo44
LvTyBJX9d4wly70SYIEW8YOd4gvjhBtKAppyh3jgZ4kp7aaN8yxAvak9EPIEm7Tx
3itxr/pwGf+WSnWpbu3XPc9RiJQYUjdehvqCCFA4mdBIx9P8ZkRm47mrJME5eWXr
DZF0hdRyE/0s4aMycKxQu+cLyVak7PHMfAO7dkHv3suyKsiVERuP9njP1CubMWf0
WtKhjbyodWwOa+UskIIglhLyHP3MpQV/5JTf7gXxz+tchhH8lbPkLnxiYEnKicbI
Fomb5LiFgUV4mG8a3sVvaNOsFgkIm4/jx6fvTG2Li+VCuJUItIBNDdlLJgjHL9GV
UaJFmETUfXhxRFX+Vy2GersKLZNdBCcYreEZlddzWrllq4wkJX0O/gwLppyfCKma
5nDOsoJJxw1V6xv5mRv87flxiHWXXhT4uxhclIniTKsVcP3/4PQ4fZhAqeuUvCl3
Tt0IUyQWvy1rrNuDdqHNLN/n/G4WoA8I5dYXZ5Y+uzXeJIc71Gb+Ai/8Tgvz73IN
QCl7YYJIebqUTLwdJm9iA13mUn7MscYnJSJyLECORjVkGtx3Uf0atuaj6PEFsOtS
RpyI5s96QZtGJYtrNCoaPk5A7LbxC4YASTb+PG2KDLXFo0jy+S8rKzSQymAot/t5
3L0/BSVG+JP82kDm/2tV08J8eZUj/217FkwRznLxMcR0hnENnZkBN7xsKDVLiBb6
Okr/0Z5azlha4ogOgOeoHmqoNe+dPiuYQSE0JdOl5Iyh0dEzLrG7O2Mcf47VWhKU
kRC/luKfmOr1oeefBh789V9BA1A3vfoZUmad2xeP4Z6QlvISuIUUaU3M7S3DZaTs
DR2l+olHewy1JcaKFBNekNJdDWG9lWqwovT9wrKFDOizDbbmEJ1jt3r7PieZFsUj
VktURcmxgqSeGjRh1wxtyJF1YXihlhwomOwDzrqaQFXMVMAoNlAEdMfgp/i2wmlZ
L2Q1PK2p2JmGAO8nDAGBuf9IsnEJbzGSf5gMngVqFcF1Q9lbDZhNMpfVz2z4+FfN
AGLGlr03aYWEjdJzEWfd1lir5Jvk9QQfyZYfsvoiFhmKxIYhTYuPgr5Ir4Ba07X7
VlLwgE+LskRLyMI3FYqyrZvxonr343VuPJSwCnWrL+prtTCucCWh155y3YxxJYqv
SeJQTE/gc/rWMCMSAT8zKs8KtPpbkxTV61PR/VpdXUhseoGAJA43WdJ9zbBi/W1u
pWagKOz1M+JvNbrTWX+s2C4fxIwsiW82m6Jgq3nNJTJBGRfYiIXAbGu3qx4xylmD
y3exwKNlYSUrXJZwkJdl0znopmrZj72W4sUJRa+mg6BpWrAtE+7sbUwT4NMEhhKD
S1r8YCmnfPX3rBJrfaQVzoMvtxrBSDyVk69EjgQOiG7ZSJgN1v5j103CtpsrQcgI
heRtQhxg2lV2C4BQMXWIBznFHNq0UFcbDYtF5pKF0W1MCmjvuEccggpBI02Bg4qX
FZdMoOQBWC6wjNMWPxk+5eZLYI64g3X9zAnfdppyciL+ug3locLd1GdEWB6PJJAU
ghuCpv11GOXu8jDxcFnR0+S8MeXG174AifJZlWKUohmt7yHSBnWKgZnjPOF/hwRM
S7/hRkHN18CYo1dEXrB/dUNqXKjEnFaxayUrJlHm5eSSlmELP42HH1FJAS9TpEhW
r+CyILOLvsnWkmIb5nMRpznsfusKWH1yODKKmIa2zY7d5G6HQfqBfHUBArEHqQc0
7Lmxm3nEfgYy1k9WUn1meZ5rAS6l2X8f8KKXbKKtFQl9C8oeGFp6qRoNHApCE5mC
egCIP0rK4xYsQCd3tBkJTQ5xqb34lM2aETbCTXvPX5xut9oQZ3qyn1ATbn42bso+
AW0ybub9YMUEs8KBuJJJ19f5GdhbrMfm9+RzxFWDi8baR3ggK3EDIigpiPFbLHRG
73ilZ4xCY5gooCCsKC9GhMnSayAwlMEZrKzs/aX7zVFsC03TrLlZlgW4R4s2wcnS
Gpy0dKjnspIsP5fgNXckdl2Qh+H5VwGSnq5VKjfdIg8BSh1/Ks41D9Lbo/f9ddyo
GcWUkYxI2ML9gU8xNXnYARW2VaCOvZNNL0oKeTjT+YLr4N1XB7tL4ZYhJeUVj/HW
a8o0wWDJ0M7VIGpFr4jYEmJGMp5RzV3Quty4D4pvCRU0nqf9wUx3Juw1LGKTdNh9
U/Dihl5Y+oUjVAbrHWkChFe4oqgCdgPl+bLUWPlgeTaua/eUVEDBU3u6Sp0Xpiz0
GhaLpQ2d1BW49crzKrSO+LYgqTdQ1PPouHF1WRu3CdpAeUB+kHH4T+NYP7uUpvoQ
yffYa/ZUhNkeqNce02wWPwVw10o3KrNr0+9AvRAhGaXC1KoLG4GO7Vba/o1g+Nqk
c4+xy0IW3unSisAB6PXekWySUjixU10ZDv5EBaV94Z/q8/xLk6UnIxygnb735lCd
CvlwSthjDZH43/qAR+fDyn4LYb1DeX4srXt5YaOv0Va7NCfAkLegePMTgxMmuELg
2hohvJ8JL3z/abUc82cBWx7n/DJaChu9bi77lKutntmpRJoKsxjurA5KuS9OdvBZ
7n+jUGWeh0LChYkSHUu0ggQNvyi4x2w/F0OaQktT5NV68VpcT1ateotI51iMhh94
WC/DlRMK/MA03kn9xuoC8d09c7LoSQ7HRvKjxsbFY10a4qczR05jeHJnQRCfv/F6
1y9umLDpA/w9HVc18gfpAZaYE+s674S9bF+ckHzYLESctW+UIoVlCnpcAmUAH8CG
4f/vuMI7Y4fZDZXmL/5e5tTSY7iHd/NHc5DfiXT7RTOkd4rdVZ9n0/qbNnM6LVmw
4b/HtbqkOWlWa2m20+GGXz2MGGICCzuxuzJWkCDLu3t9+a2uNiqD/BNUD4Z4pc42
xKN9ZtkBXK/l7djm1HN+ynBxQ+T0GDHX7y/at3AssqRWdT8fRpAc6aENQDvyPMZZ
TtzbmemmVKNEvyfE33fvqYr+IJC0W+NnG24W2VKQdwqPmJHqJKj0mNsW+WpQ0Tvs
rMshxg47+TTocfu4zUiix+KA1IKZ6kyNaFfAbLXvj3PSvn8cIuoiKnKzu8Kfr0RA
2qfMHfLxqeejPlic10fxTwy3bSVj4qpo42hpKWvcbpdsArfl0m152pbzGfT8nUq+
d/Yo/VUo0/sfBbi//wJlkJ3XCVsksvEkYtM5DGf1UNV2Tz9OwM5q2n3uPYOZC6ip
doJWHicD0uaq62n48XeVhZLTLqWhsvVHk5qbQ5UBzCBqjkLOJCMkzfzvFHM84q06
ebTPiIKkyVM+3jpQrDF4xcRYGF7R3SvagxYsJe+47UXGgcwDeKkdBgLiP37fbLmO
m7kspqaqAaOPeuA4hPtdoQt9l+0dPpANcZbb1rFosJHvuFw7aaWvt8syEQ9Cm+jj
PYQQAhTH+gcpxUs+0ngJSTzfJzpzyZwUyFW1sQYKjNJcsnCMI0FYW5T+O2EDbNgE
hZXLJOfEg+cIW9gHN7aCEniEUUUJVnjKm0/8sQJBXP4IUgObmr60V/eCHolvsFCi
XRg70g//568SOgyPSUyNMuVUYIT7dLwKdsuEvjKhu43da15BRgXSOXI934e7XC7F
gnoim4IdylcBDSnX3yp9j/Y2NoremD9Ro1vOuZPv5FUkRX8MnHlAfHnoa+YDcrCQ
heO8IMs9QwJJhgXKKBXik7roFo8WzC2rrhr5hCD6SHL0hWhbb+h9KjQfDPWBlN8H
xPD0hlcz3RA1NqJgl4Q29uL0qhBdGNPWraBRFnh0/Khst6/Wss7UIJSA5cYF7lha
zOXjLVPiyrSaV5tdmApqeCAGw4tio0tVIFXkggBUTmeZZ2itzWV2ihEeXZpQkSU6
qYR8bbXlaV1bmMQsZmfOpf1CktqXK8AhIXxYJ8FSnG0dw0TBVYJwaKhUsMjpgo9/
k5QAAHrH/6jeit0gOECjL7c+LwkaurOYBIQmO5BTSCLM/VTj/kpWiUptCTdbehoJ
o1v8ErcNnvkHOsbXP/lDYRfd+TJhEr7WV9GN2VQhkdAmlXPatW7YdvechI25tu8d
YQ9ay7UK7wgn1eopPYF7ugu5eGD3GQ101+nCXMVV+oZi3NsDiiEgHs0Zd823Ouoy
BRlt32Kux7L+KEcX4fz6EiCcZRKNyXF2kfU7WIFO4IGJD+hY/7LAb43FkO1yBzZF
IEKWgkbYD/3RB4NPYcf65ZXn4MazgqkET0FUvvWcEtBzfCrzfx0mowGANe2KEhQ0
DdOJvb9b4CvW8gNyCry3IVey5G10K9EvQtlb0o43ZNstUr0VMXokNQcsLZ4gT1Lg
VaKquupSECxZaQn6ev6anPIa0g/h182OrSeG7Y21e7U77Xxs/R4W5UXhXnxlJu44
Hn3tIQHrKOWMX72aYpvOBrDPl8dJ00FbbaVJUZO5yeBL4ggUAJRq+SQw6+XLZ+au
epnwvOrdFtVvX2EJmpTYjRiIlftd4KX4GY3sRn6dk1J7AQm9Z2vLR/PbmkZSMh6w
8ZFsKfEnj3b9w7LSCQzMHsC5ffdF+Ob2V00vSiF9N21+EzOhdN9jJr7KmkQqfhlC
H0nyG8TElvYr2C6inbIrXr8+jizBbOtPifDIngTylwo+zhvPM6pcSBUww5zbM5W4
O7VCIMW9RW3zUc8ILUW2yTx2Y7/altulDyPGF62cKxwF21rgBKBp8qHawJnqwXfT
O5WTMeZQ9TMV2iL/4+U5lmRcX5J2rvCrz3qL1cXa0lXa0/1RWZEUopJBHmsBQbsT
ik+LOd3XMxov3D8h5UHGiyXXOVQlZ+AWzBuSx+NgneSiqOVmBEgZ9oU25MIJ9Ogd
UubALeO4KfLEp6TX0TpWdXfIUXzMPA8Yg/AUYgnunVGsAmaJthSnqGZRpLt9o+2y
Xnnx0ZAkgR4EqofFRmtMxCStOWWv8idcmJm6N0gIs1mqbKTzqqLIsu6nfXp8HdY3
xuMgBZdgnWooOyesb9Nf6a4lCB9b/eLA2iXcI47X5iUVDM/HvnN7cyQoyv6OWX5y
ER6okMhwvbhliNeXi+3X9nQzP0ibfetj5AfxQUx0AGAVlWnTof51qQ5EGTYVyaLn
XDG7mdkIliu7kBmyzdzBZK3hOb+pkCendvABagI3tX/V+JRYBV+SnhKYYXLR1Q9Z
E66JmhP6wiF2+a28bwtkTYrzP+Zkqzr5DS/tuBF4B6SvJBz6dCvKEwk+Cf2lEoGa
VbQf8fohNbWSkVU4gLG/pE11S2MQSe8z3Ve+bEAsfPdKG7T2ETnQI6yqd7Sgtw51
ds/jXNGUtGe6SzzW7RHEhiWIM18Jn967VZqEAVM19V5egeimkAMKCWmBtaI6bsQa
eb7PzGvgni/827s6CV0pTSgAjgReYX+TuGk5MIaOMWpwiwLsCdXyKNCAiDXCAyAi
xCvGakz0KuVKuBJCNNiDhE9cwbBgOJLzT71/YwO2MbVKRqDZW3jY+akkMx/sVGVr
jhuhlxY5aGP3LsxQHP5QFHsMDGUUGMiPyTceJuXaegKNcXWZrYOUiRWu+0isz0Ru
TSAyOSbywWN69/8HQT0YOihVrIEck6H6YF2ZXwOWJOiWSQDbzy9Fzn9zW0y1wken
y+KPh6ituSJPYEvET6I2ebvD4RV8nifogNjUgigim609j+YSG/dLN6slqwlQRfGJ
4cr33vIIc7I7BB8B2ltpefI99usSD/gsclpwk5+Z4PwbLC6m0Y2qpyPoayYlFstl
HCnwU2pgEOYlQwAGRN0S4ZM50FPqWwq3BmIFqR2OlN3TYZcKS1MVo/HkL/ytNA9f
9c+/fdn62f1A2qXDOvGO4Df7KaVOaqvtwZMbCwEFqZ3u109gagSTeSvbBl8qEruw
/4uHxDb66BRPHgrKHC05hpjGsRhjPjRqfHtSKENqjYanSLiXiu00ZEFWm5sWOF7X
V3w4YOEuOMzpyizM6b7NBo57LPpqEoiLZaclogeEcSiKfxH6utIhTpt2ZiRVL8Ai
ZKGt08ihfLaTnn+rvCAKUOKkqOP7c8Yw9OH7bKvlGX/A1TuaC+gWjiBIJxd5A4yD
vAJ8RqW47kEolPNpVptI/Yk/s7dFXQFb7yse0btz3q/quRxZRiJME37gDkEjN5D6
xlYvUuJkduVxI0cjT4BOLlCnGh7kqJ5eKEGVBh52tzVEO8Zt5Ib+2VVYJhyVMzDO
JvJCriB0VQUnJuikzcXe6BchDQiT+BM9pMxtBNRXDgU2OD35eVRmcT27A19Zf3Oj
je80KTac6mqRIc6FEq8jxpNg/V5mGC/fpAgSFbpT7Ecbqd4tlDQq4076eMqMkxUE
B8A98XqP3WlQSZFnl+kLV1YYyYyuJkkwKnaHqJzSJDEHMyN5UjyAHXetg6Ql+Nxu
HajrzCkEgweaTFOo+1t/LeY+px59atgQDMbNcNrdJSn7nmR1KKJphD9qtSFvQHlQ
KtaJixVc4fK+i8DNbaDz8KCgmxnu/cbAXUkK3bqSdwMjcr0iY+Mpk39kh0belfWD
HNdZazWA2ahAstSDJRWZpr2JCc532GFGPDZ2bLJ/Tn3HYKHdbUhyRCyXqhItPH0s
xuyXymHfgS+SPPjMGLE4C20yJ5ZvvmHrJFVJPeIRvduHmfGAr5prh1AWc0VjJwOS
3Gf8/RTYUk0GM6Vw1r43u72rKYAZqSBSchv8lOyQOzaLhZXT4yALrm6X+vlh7reW
rgtD533pfOuhZD8z5fZdU6mJEsWo1CaT25DAvsNTdblPlqW/OC1Bbo5IyHQw6TbA
wR9EhLgoVn1u9Y78O8ng+Mj9blQzK7kXkRiow81trx9mckRFcQXPkpVQrprILd9b
hZJlYDvXF4U0mpJMIU44pqCj6YQhXYiArjasdZd3QjQ0/VfCG9WNkUcKXxd1VFrY
d2o9rRImImpVq39ssStQueZ+V5Bn2n1CEtEovqnCEnVVGzCybNOWA6iWkSEA285g
9/D6V0oB9QFS4jnMXgZcsfhPfynlJ4FqK3P+57Vv/KyWWTRTLI81st3gohYHCfBz
xr2TOP6iF5YB2Zj+5wE8RE2w/9vlgkEziREMSHviuhLsApu93SK7vWIzfOJg3pEs
7ITRygmIDIvH7TqM8L59uXnLskCCX8GhXufvM/dkVZKsTst2sWR6epzVmuLUzlUS
Z+VmDZDpIM1usOw4q7ovcXpgYFS1TOIgSk4aetlvcv/Lhak0qmv30WcyiiV3x/br
9kxt8OHSsyfk+R+YTsV5thAvLx7rP72dZooGjc5gjLqjjbbboUKdmZ6xdu3jNQjn
nq5xUadHXn2OdyYjzlLLnMEDdHHBSXa3LN/80L4h1LfC45Us07WiVow+pn9ntIcw
CS65sI/OCEuZqOAmtX5nKDR5qL03wEfIx+esZEytBZCiYG+hgyOyTxM3sfXKB2gw
QQfmue1KcPci0/7nysGDN/RtqvLtkwoTg7uTtF6abCuclWpNvPWHvoEkSm6qSFyG
JMfzxiodiHnaPGf4h6ia0BYOn//XiF6sl7jJRpvO6kKgAad7LA0742seBJ/SgCfZ
C1ib6ppIy5nxpZFKt5E21ldGfHpf6oVkQPwivYyNB4V5hiNy4VaRaw9dc4gmIned
jKEbmoa3Q7BObwSzbp1IaRhaqzJUAzWgS7C+9rsT/q6SN8Q9GY+6xtQiVPwRa5ZZ
s2ip++oiH3Ppn/co9eXkgfJ6N9PChusk72TyWoC3rMJ2DbBFwAM5NTzBdFZ8GHnW
fyIl/oMUKt+ILGz4tRcwuF9e8hL0MTeb1CH6oi/mkRpbsai3i8J56cogx0kRfrz6
WoTVPCvj6+odzcOgQS+vKzqQSXhCoOYrAomhVOlQUhcDI77/qZCuwsurAYAqZkFh
/IOrDk5C5CsJxltSI2y+8P4SxD6iqi0TrclZqIHzWy0llHmZBh/q+97aKQjw4jI6
5JikKjXT0gz6EhBNjGZUGF8yBNcdZkrPJQDTcQpgjLJYEjrPbXIaMWt0iYXMmL58
wbnsc5u1ZY+u5kQKxlNuzIMU10Y1wm5VrDSf5Y2J/TcTyMk+fF3z4QD7xQce1vAN
FffGbRb3Z7clf6dnbHGRUe1bOspO259ct4KFl2PeXreeXGqUYe3WZLkOlo34w49c
rLv1zmgvhPuQK1XDi+UOT3ImY1eS2lyf5ynhemxtuq/cdz8UVMTKsMtCRjRb/TQE
i8dTf+SwQJorlOC0lE938hX2ciNHV0w4+uDzPL44OEBgz8eQ5/jq0qZW2QaIj4fl
6MuLKB97niJaOIcjL6jIxgMtAkKqlfvk1oFfs6Xgs8GvJa7GLoBGLOaqQCNyFsw3
dV0xOfIJd4YIyyTxj635ppCxZwKWEDG+Vtqt6BJQcBFT2vFcfGf89rAE60RQQ2Vd
LKJaUl5EbR90uRkfmhAxkC0c7nW1NEzokO3iR+NZ1kyQrJ/mob9qxasFPXRxCsee
7pII4MSlI5prV0WsaMn9Vy1OJraMq9CG0eK5y2NP/TU54Dc7et4EbWJ6IhN2BPCN
wF9/9nXb5U4sojRpUaVgHgQCoCUw4umoRxhG9sWxAwn7rGqXUcf+2ozMJPW9iJjS
rq5CRsW9c8uNkE6Lm7bdSQL5DqE0HMNf6Aqo8v25FlD//9ZxTVUmy+Hp6pzn4xsN
gafDcgb1uXysjzNIvB9jLE/JGeu3bpnI6Pd4WCQm1qj6GAXAdli04mREf2zcV5j+
AOoyvl21bUnidt7oiPkNBZ2MsFOVekd4sRctYoddrZosSLnKVCcPTXYu1VbKJVL1
Npv7m4SIyB6D+iI1ndMfWsYbFWQV7gHE6eERc1z+Ik4D4X6wmrDeyJg2IZWLcqaO
TvWR8zRD5ORjxp9/ftCyTiAlU0Q2yz+qC6eO0EPWiDfFj3OHiKSOv/bvvdcBKBO7
W/FxM6XHw6HY3nQ4bWtns5FdCGIJ8Hu/rKKn4wNyNdjLhZbPWaAD9yfRPNjGUnnm
teralTg5/AGXP0eT4vZpIDQtmFXrU6rGhi6M3vM0qUvuqoTOTlCNYTvu12P1Lcj2
ZLRIYrM19ElxFBeNi84ftd8PjThnOZxlfdt58j05on8veszLaaOzpDH/zHQqGffZ
HZv0s3zYIMNE0SZ4Eseaklf00xZLhWJvPoBbc3EKnGkKD2/qu+vLmXY5Dz2mPxrj
I5Tr0Gfs8WO/0wfueXUUjkfwLth79X93D21riB1R7lZl17yx/1EFEhqYpTv8JOAb
uj8n9WhIKJmUJHowt5jdvFol2eSNqagdXS97svAxUG6EUN5aN+x/svAfDnGrJCPa
YbuqADh7hvo0vUmcSuVBCnpx92vaOFESfZ0fxZe/fVYWJZKVP7in3Ptoqfj3CfDw
oMhIAuc3nK6kANWPbDifFnN6VgqO4I8luJwYp+GQtoAYfPlXzxyO4Vj7fptEnB0h
F6rFruu7+ADxaLbNmENfA4Rkl6tR01dnajCJTklq/oTAw51ORQogHOSkLTgYipWt
hf8Ne1O5D4f0xWi5id5xMbZKrfg/pyL2ifLGnRBaW0GA+TmPgPoJCKAgrw3zGP3X
PO3N/fxAe9/ArQ7h4Pt1/qDLKtx94ealuV3+pyWqcUOLKMnsRJjdZPE5iICV2Hn7
qovAfE9xjVse1LkTBmyA1DYOEd5+tqk45DJVI2L98tZmCHW63fJ5UkUoFAEo/T9j
CXWqPVVG0qHLc7+gNWeqnGl8JtWADhGKkCXmjc986LQsKAHNYv/tQZBAkiLXhH3T
pmjaRvQcZoFUCQdzLsMxHXtFJXvj0dQq9NLbPHaQIDKge4Bh8zWX+zotC9kgOuUF
FxbWqFYul+Z7QbEF8tdFgIJfpPIrdwgYpBUgmPCuNBMVx9E2Vrq1rt7aHy9oX1A0
/thZnF+O4KdJAte0AiNDYesPhqvEFYU6QuA0FooRH8RMJUaUZjoziFYhx3f726BZ
SsuNfCVMrQpBNgMvpSZmRaouQgSTNNjBQEAyQo4JbFiFBJfC8Ypa/6DD3tajwyhg
r0k4BVkP+MzFbMqDrrCI71OmTxVjkIE46Lbq0Ww2LhE8yDU/bKpnUva+yLTLh3jM
pigyBZeAmOWkNV4lfaIIyy6g23ZXd0nLXreZ8Kv1PYcOzOSvWV6/wW+C9Ibs+49l
vtxtFO1jAiIIO69lRxWeWanbRt6jU3sVSIBlxuc0t67oc78H6nXvdQqkzsp78X4l
pcY5Nr2gjqPr5jJIfkPvaADAF5zi05SLM37OasR9ne49itYD229bsI3RcNazY2Fm
7dwWaicikM+aM52tdFqZr3DZASgfsXu5qN9LWyhthd2iBwbvSxVo0pLQjHEp9kmw
q4GBuIBIHU2NWMarEMyYSmj8d2M0v/MDKUj2/cT6F34kEhq7XkCXAiT4fjFrnfy0
ucQ+Rb1ppapJzbVhUoTK1aAmhtfD56YRk+la4qxVFDdiKGqlOZqnCTJzMpIeAZVX
fZy8Ua/gpilof0ilXqudA0uLrys4OB5Wo9+qaKJYpCQO1jKMOdATuwNBubMoHlo0
oqEXwMJJcVipTF77n/XPw3eqHbk4bm4SFAdP3eDC8JAsKcz6875J97e11fLeQe8A
fnfxDfwkM45NDfom09B5XvlhCxxXKQ8RmjxKmLOqYG+44mHr0CMhd+GMjibWpv6N
4VtqAvBRw/5ImvxZ37Mojlm938WA9c6HuCjPRxxez2ShQJM/k93uKmX+76rAGXP4
IRRgnq3akEQ8B4sruGJTIBaVo2zyomat/CWPKDbQC++OgesfjcrFpfepSiLW+Qy0
YFy6FCU5Acw0bn5Tk87lsx8nygv81e8lRInleU37X3e34vZ2W+VR9EpoIGT9j/0n
dTIOjCh+Rd59Mve4wYGCN/LbL25X0fYWMujnhj6ToKrIzR96lsKLuLRB/5JSOFHz
aPaJkjSCAkyNB1AuPOvjCv19qhX5BvUw2vwS7Pe0NIZIEg611tXSgXdkIYsY3TO8
auivQepKgDtZxg3aLaBcsp9CborDs0e+PFRLM5KWedfZodAMaLEeQ/SrCS3IShrd
mv0EmOxwxHZ0o6tZLllIDEAFqBQxXu7/i5T0IGwzuj7MM45bD/qtfhLJjK++f317
ak5Njg2ZDYq5CJ8l1tF4ugdyI8Hzc/x71COFhX7kGY35ACVA4jWfB6Yd49mm80RB
FVs3VeIPE9pISf7FoERzEQjERO2xdp89FlSj8/ymOhkQ85DfX7gKMuLVRCl+cvF7
x8Yg8rvf0rZet/bKtTagqlaI3yxRCwL5Dbzjyq4KFqLU86iG/T3/OIm2FuHX9xXY
AZyqwLObTguspBM8BaEJO03vNTTOuYpjtlQkmwCrCgn6eWLEGmxgflusUxD5cQZs
sw73N4p0M6eLQOlYngP/6m+daJ4n+mhywAwVBIzJxasarTppB01xTpxAELQ0AeJS
7rIST4tJqSxoZnzT5XgjMHJkUhFmF+2F/hbFQM7zpPIdS32IKk81BeQXl8onluMc
cHxEth/warKDQqkDhXhkWJh5lYQTTs21cIq99Wqepl9viZI+PfWNAxWm5l8tgTUd
tLm1f/51lzTSFaW53Dxib1K+FkQljFrsK87q6XfnR4udR622+LBYA33gG2A9C9ve
DTNIWU9XdsuD1n15eXk14Zooc7vZQ23COXBTwqXWowOZLR94j38dvNPZBwk29X9S
kepvMX4/tsL4r5+d7a6Fb/pJqDvVct8dvmoq2LvuQaUqL3NyM7NcFX5BkEe6hUiq
bvYEQqmXxyuUIo5m3XSsxPOHEDfEmnRFg7yb2p4LIQbYYrn4KWWXGF3GJ0n3h9WR
wIQ5IX6y0zcrI54gpiZSHZdeJadUfXrYhgZXzLon2TJaNmvAjtBI1vTrO8ORkbUT
uoMehOBXnXbDunSn5y60D0tiiWnJaBBl3Q52iJODpWghsIaqk+KgTDfXeXqKnAF2
qhY6Mybbt+iYc4q0QKinha4yWOLu/Uyu8WPkAW4GXHXo2RO/MJvTf473RGRqWfBF
ilO8B0FUSWiKX8H3M3xKm9GorahcvEDMXZux8oI1dpIwjNxBURky+sifncaP6j3I
aAMdBpxl21kIMlNvbCBEgIoCrdKBqYK1iTJFUh+jMPX+eu74L+1DkI/6gC8mKqF1
UQxDmRweaRaPFg9wvcVPkNsDscMi5ZTMucwm/6wHRTzPYv3EkDp8JhTBf2o5GgzO
Sm01rj38j9B9LqkQE/kVecIXCdNTspHSP2u8stEfXyBFFStgeqUJu9Cu/SEWH6t8
tnekfnL/3kfS7oKGRoqbRhjzUXjEdm60Z4CjkTFk7lBtbUfInwbx4y8Ln/cuDYI6
IvPjL/o6bQSHGJgE0ix2c9AeaMKJhXMLQt8cpGL2RsSC4qpLdDt/2tkGvrUkKgRX
xXucdF2RszXnRlAp5Ii/IDhk0hOm4BGb9yD0MKnPuyPujxShrIkro5bXhorbm3tJ
j6YhYCMAF5TZn2QzGdcOZ6ANlhohmw3bO1cgFAjj2t7RtefCe19XPm2qt5Ro+yEP
+/+V0+c6UxI2zgoBVTJur0jxbiv7auD4q9dTdsVYNLN6uxk2NwrhzjTq9UEqoV9W
kWeaTNRxccOjSsxpaEDgH1zDNzTzgbFcdiMeUMcG/U4+8QyJ5Pu8Jr0h+cvauiyt
gI8Yo84DtAolCUqtYGzA2tW4riVt/lePA9vdQyo2WoXmxhmWezAwv3ViCAWsZl3q
9D6ZSE1W0wGO+5F8cMPx1AbdQ91yyMLHrV8RnLfHiq/BaTnku7MCQAx2N3mKYYsd
1Nna4beEvzBC5DxfRRn0LzPhKfW2RzbjrhU0mLf4nU+F3Mn69hhHxSDoikITnzDr
tM3AAWI5vayMdRuuhevR76/5QkfWqfzhJrdhqldo35tz3eQs7ToikAUS4MAto9sx
pbVDzXFDGFwIBuS2TIcjWzZ1Z1tT0/x5cO72igCGUb7/Pfs+LjGAWMNQQgnB3QSa
CTAuhobrsrVuIoWTvd6p4a3oGWQV3NdbV0K9X4544F9/khOwEQNH9jglDEQ+HteG
Ynaz4e8hgMphQwDTlXwbU3BGbB5b3t8Jd0RrhA3MlsZjWFbZVt6iYrdhWXfbA4nl
ceh1CZMXHx3W0binamEPcWKtK4MMc9NirNZdSGxVY6g5gWOD3IP5v+wqzziSkjQt
+Z2eytaWcUFVH3OvmbA96RTil4nvlDN6V8rLHhJqGF27ttoY7PnQ/D1PvMzSUOV1
SDfKgtLSjcgqtAbCvR4nvLAov8bitv6Baj3UP2naMrooih3l/FALP18ODiu+t59N
8jlOzWe24jAns6U10CRho8QeCgEVrO+M9DC1Hkyy0m4oP72XNZ3jDnQljq15BObI
QAQOtHQ63LyPwjvlAj0995puIsp4e7TdrEJE0nCGk5SsaxWLfHhTuwXFhRFexacQ
adWfSj5HAt/ePnZRtuaheQ7JwSqrME8Rk6zDiKrLGWnyr2v+SYSGTj2hlA3I74N2
k2alFMYhCOaGDPQye5EQt5C1x2AuM9ULn4mW32FNjR2qBYOIqy9pMZlFFgakuK9X
b4Xox076+iThmSxy3W1PuKUpXzx1H37xtKvrFRWOhRjEs2NpPulymOG1sGaJmbEv
Y07k9eMAwnrEpYDbxQAZzsM9n97zfDkPoiT6oTDEh04/+L3IpwYV6tS/e/86X7xd
OzGvGtG9CmNpzF/0vPHyN+MITBJJ0tmxBmUlpg6US+0lctVt9gT2t4Arjar4F2D3
4NMAx4rws19lO6/znfLX6kIvb0xNUVCYYNlZ07e9iJkyVi+WHK4g+TifnfUGPb1+
qpT4BXLbthG76VdSOshDNAg0fhPJfmRswlDA+Q8Q4RRDrewly8kK0E7dh6KgQmtE
zSV6+o6WTawVZxpIKUC0Q7jrK1A+YkjRMN2gr4dLUw7o1x8JAuyqHTUl5niAditQ
ViXsUywXmjIcxF42Zyc4xdYK5M+WsTIWh8/rzV8Ymz9K5qucV08vUH9aztZzKB+o
B3LkOXZrM0xkbnJc8uqu3hee+4HSVto5MdionYSlT5BaNnstQFgUg3hNy6hJShdB
ORrzzK5Xk/5d0oSAcYgkIx4tK3knpek9VLPbzU6JrpYWlz+ozmX43M32a2UnDY0I
HIm4392c9Lc42uOvyuhnotgtJbb9cbqhbWKAcOXk7Ns8/S8PX6pV6NQmD0CQnbzo
YjnzslPt4hb1Ia4twN6lWSfXmlKzQ7+gChKAGxEkYDYM0UyXjHn0i/X2GsG4H2m2
2dm8gP27ROwIyw4wieGM93lHUepbUheyJpZ64rR/ZACn+x13fBqUD2ENHTpt/ZOh
wLk/eBkPKCrBWgvQIEx7bsZ7ONNbordf/DfB/sPny6R1RQk2jtKjtDV4gKjCrC15
UPFUf0V3EnkpN9EfUlRQkbfyKRqulTv3uQtGSCiJ7qtZcrtXLpVZPqX76zMt7WBs
TwsiFLnkU4ZG+Qv8siLqjS5uG6zsdXePuuXj7KKjVfuiiymCSZwt60k+5FhsIm6N
tSZ/g4plGilo8JjVWf++odEUnUImGtfbBStT2O6ZdzM72RT6nXMB5llRCV9w3Y10
rOpXILChgi3guKmdBvDPDlrzYJ4XPpAR/4Lnn7qjrgxdhLQ6tNAk1pBdyJ9QZN0U
tOk+f+d9jRdAYpHfKvJWTmiAT+fOJ7zw+AfWb2dxP/oUQVrSGArqbu4J/wZrQt0l
QPw4dt1Fmu+5iKNwPFjWjQ4rZg+mZBsSkus56VS8msVxMVpxnoSw7DNR7YjoZn6W
9NmCcBJHuH40E+4b1rXptC/oZFiPeRhSQ5yr//GZ1IHWdGfQZDIf0vVQoQUHltyS
oF199kLl3YB0DNWSwOKPMlVYtzdR6OYvU3Mw3fpxXO7uOoC4gUFoYfN2jHzKK7FB
HRxN9dF14CdPiWOdMZOM5S2ocj5oeLSpqlz/nCNWIxGkRSHsUnl4C1bl9G08mZpx
DdI98JjRqI+axnMxbtAKPCOPBEQTaeldREraVH+siuuK8CO/Pt5x0i86yZ+nGedg
ej5HWNsIKYLdRi6MViz1y6/HThagvNBAt8YA/lWTYrf8z2TSQIlnanpR6VMi8EPO
nvTytr2W83wbh0tG6FAgpzkTiiBSQklTXmVICx1CYs6qldGAe52NHB6iysoJDXor
6g6fvmVNo4nKpEY7UrVTFOn7FN8c3F9KLWwpMK/+jbc4xIkYhtdzjvCBILWgmo7x
KpBHVbzpEUL2L7yjzJWmTHsiENU9XGUZuMjN6Am1+bBfkf6QdwNif04uLbft5DoU
udPpmGdDD42SzWT4kN8sZdAJxckrQAjJLReJEwc+vpTG72XboWvnJgkYywxyQDVu
vKKoiLdcXv0EDOUpoFKAzodfBB2iorNEXxzDlQak35YI9k9ysI36AcP2/oHXLFwE
rPW4Drcvro2wrRMbsfhLobluecJUuDtiB9EXtlBINZifsoWpNSa97npcdkoWe2ZU
RSYxkFJyUTLnjjMQHCTePGx5xmboSn2Psq6zORP6qWfkjG+S7F8cZDJJ3kJouT0d
Kx4tNRKE534XXEnt+GyJP2+X1tASVVd2aKO5KBn7PPF3AJdDVQgRl21CHYZVBSTt
InCwMHWGBw3akFBmJcDr55m9+40eNpLd+Bei1ff75i44Yt9V3KfIN3MNk2ThP2Hc
JJSwajwXglaBiCXz/gqNG5AccrTdtSINir7UMdZsc58lZMjQsO6RNli6lot7enLx
Kzd2OSo29VDwZXAPnUPLqAHxRwowXhQXACLsI0CVMQWMIrZNqG2V0g5hmjg3yLln
P7PdjZIu9sAiDmGf+doD02N9wcNeZBYPt5/ijfu8RaRXXom8KxHZWyAiQUi+EoU4
JGZofFhrDx9eQQ9lECjz692oyhxrqrWKUvBg6Iw6HbfwpUIdmO4C+P7QJ4tErAdS
UdUUSvHGbz5zbtJCeg9qveV3QYUUT3snsIkJQVvf9mjJtGpsh82hxuiassVwhSoU
zvXrpg2yPFv7nOimVunZh5ZJysL+zXN0HNqr/bgoCcKy7RzzQGEuU/XwZM8K+Jdl
ZHFVYOrM8V+OshZw3b1iU68DsIyBwbvMDO54ty6x0E3ewQO6K0aUjklIgYBRP+bG
0Uk3BqhHqNZw/HjjLUE1pQ1QiRu6rPESFt/O7gxowrwIRMJliLHoVSbmlbZPr4rp
vmFB17rcigNIXl8FvbKO69vpsjZib8oCl5eCjcXZGCZXXmWqyipDkgqPIrwoI9ql
E9RfUYs1BuMTF1f0LgFt2pBWysF/2tZpseY9oE342KNXcIRfBxa2KV6PuRUOswpk
K8/W1iE1tVco5yhGkLLa2htWMlPuTgtnetibTLoBZR7YaLmfNK+m6KRnkbx3mPWc
1KU8UpKtl5M9eTQYxvP/QPlBASmq6bPsiVtOS0Ns+DnvejioXSe3tkHJufZA3K1o
1dv6JnWmagLq1MbDJcqFWlgyABmNoLJTWZaxSfiMdTYwImbC4kClrIyhv4YOxnZx
ra/Z2d3FB/ENfZZlugswxiEiGxdER8hQgERxydeHrisHvjg78dfxhtgDFfxlaT16
5WHkCLHACnmHqT1lvHSeWG0H2FPE7+mHaTQyuqmNEnLD1IbFtnIgNiTQdrmoxUIK
QBWQzad0tpJNzcaX0oa9IWpwFm7x/8qgIU9XAGd/jCuahXyZqDarM639qf1HR26s
uE79FGcEb1knxMaQRi0Y1EbblcXZEFtX8fYUfJJxI5mvrw1EzGp9c0gtXpzmwsA7
ddYkwqgu3OyP1qUbqJDbU2yjKzS81Kdie0YcXz6O9VP2pASosbrkOuXzwUgte4sN
k2IxKANTXKidmrob8s3aJKcRYhL+qfCVCDF73UIjUugEKJtnSDN9OabMbA2QADjE
OBbos8VrMmYQd74SNASG3FCJoSCD1Nr88bKVB7Y1dy/dTO/EVh9V8Qk/ltGIeJlS
Vzv+KHsbPNecmMuloq/nFvLK7jfI2bcEA6bVxWFZy2aX0fBr+n0ZMB5HOXJd61VR
LSq0fMZubkYtNpG2rgKUJntm18G/I8hBYFXTzvFZBZDWJlFNU/XdCTqI46dcCl2d
oCDkLEUWFrrniY2uQYcv1TMSuRGKAKHdUah3s7UQdikqTKBoK35Qu3CZDeTX3ydh
IEkkPxJCH6KTKF7RLL1PFtP8CJkYLtQntTyoHl0BtFwKCIrQJbkrRTbNvXjw/KZh
0S/moiRHd0EmMrIMoPDhq2LgDTZ1zT5mxIRhN3ZwhHjMa3PrdGdJDou6ROumiZDI
0ExtrYsM8f3y+MyjzKlfsou23xLrFfTJRWjuDPy6QL3jkMjnBSH51G+AKK6pDULM
NRPxZkbHAjMTKNX1izOlWr4ZbzTJdvq806/d4RfATl2ihfg6ysKjLa3kPw9fJGbm
ghdaXJQuQhkTvuINHPYH+gbo6zzhGVRiXVUfGG1rdrgvzrNX9UQm+M3z9l6MBg7z
eHFAJNpW/dFtCpADNqx4nLyr1dmduc84Rw5w8vEXYJUuQRbyxlBmEJj42oDyMNYe
TfPl5X07i552l3zVnnVkvWYgzQqv9tB+z99V3JyZjzZXOSE9FUuxbniLXsAy4WXy
9oGDOh+eCjHk+x7rcPD+akvvBlzyi+RoP8W0D8rofPjCTHgF+2mP2L86juhCIX2a
aqoaKNRVmK7K8L+CTcyxLWdnucfRvjL7ttqDTBh8K9Mhp0zNgj/ruiFnQNh0dh8P
AAkq2kWKsa1ENlnC3bKajmEW/EFwdXLUHxK4qZq3bipv+Eka1rGmIbZnsdK9foeO
ZaDO6zELGtoo+0JI5sekay1RQEqh0O/tLMVoPTGlBrDChjVMAnVrcYLeJalopItm
GkbvjR/Yb29/2w10KB4gdtqLey/V8lRlhyPQvm2jTV1UandHDYfRjMoNMLQKSnW4
+ZhUhpUqlCpTZNUD1J/9HRwGWdwJ0z+TK2qx6OZi+aL/wTGdT2gySQx4wvHqGF9B
+X+bVnPis+KNHu26ENkeUeFhEk7PM+D+z3u5tYptcJwiQTq68l5ZBgHTuFZRPM6W
RZxRQtLJAM5ERvIZZt5wz0gxNjG9dRcnVogMEx2gXSQHl25E74Hx5q+s6OG1a1ce
mYeTCVfz3/ncPAbbomnEc0R5sqqsEqrf3fYSPw2n2B+wN3Df1H1fUoeWbViokPjI
8MzT2V9vnUQb8l48qTglEjBlJcXXvdHsAHKpyCApFeIN4V1HyEDYfDCluys5iTBf
vCuniU97nP50486fWHszzs7cpmZq5CNweJs8fAm07sLKe9/ErONQ0uzbpAyTSdSL
olX3kp8knHZsVxVToI9BXCag1DMqqKW0OLFdDlsLAO2si0Arn2inS+ogcUDVu3c5
Du6k8DDtDCdwHHEG2k9mezNQpoRMrYQfUtVl+48BrBLqS8niyGDZCqZGnZmQ+ZFa
L787VqnJe/Gy1tuiq0mHds91bK57XCFbfCTTU08AK3s+9FY4rHRvn0bV/nm7oADr
774KXm9suZHjRyMux8dCMHEWohPDFJ2eLvuGPMXXub2AHnovka5akz5qY1tkzcmo
CT3EjeWMQWqU2VXqfdVt7KJ7AmYg2CAoFg8pyR0ay7FfNmcsFokJV2eK9nv4fdwf
liAVayZDxH/sd6rHJq5cueCWdNh6O/Daji/HQj1e5mxbHExQnuKCHXD7dg8ZMT05
Rr7/0LZRcG96igTpBAjmACl2xG16pTx6JOxg5Ph8o+NTpkKeaa9t4S3vqMyvMzN0
6ptRkTwzRT2soyUka3NfKJphlkJbWXxfCLXJXQ+LPWSZ966Ro69HcGajPTJ/chud
QeBdj1lZh8ru2+uxagkelQ9lL/toeZljBUhKmRDr/GBtiQ3Cuq2a5ZDVakn5VbJ1
4+yEcsIYRubvYvAnV0Aov5VacAef5LFqSEAhTDdVjYXeI8G2Mv1bb4A0w8pSgG5E
oh6MM6htC1UjDigAej7a+fElSB1vK82OA+SgMghFC3Sir7Qm9e9BU+CSDMkwR/Ox
oRZLj1kZxcF9k0+jjgPJ6L/0Kt9/fqZ/3NkvW+5ziEq50tBFFlu6PlNgdk9h/H/F
MOmo9kW05CyAgaoii6ptnHlZ2S143Gshdeww4gyZzLFNu6k72YHk/ilJYRph58Bp
dq8D5kQ52BpCy5A98ReGQZ3qppP0oydXNjUgGFAD73fDGuFL9EK5yyTeOC9VbGGp
H5+ap6YY+D6McVEBSOLqLTdiryGToJq8PYpWHZmVlc5aGXWR6aPbtjmc25vwIu9j
NlkZc05yV3ld+QZnl+fxVsrH98hbjfLgZG/hVs35lx1dMSBPzZOXmM+YKStvA5zr
5H4CuJg7d3Kty0dKzk4iNlnIQKKmzYaHnR/pbX3tTfzrkkshWatJM4MxnHXBF7lq
1b1NRvmJhMKoqoDEub6DQhB1wcBgVWNuAty4qnPMTTfMqmc8N7UwrLXelGaUm1ct
+8dXqZ8/ixyhNmr273ESvZxx62HnlkLu4Hs303VpOILUkut6t6gVnJRnCM+ZWIsf
c3CYaLlCQF3ntLlBJVkKTxoezoOLUQtx5Jp0csFcXOOURiDGcntdrXzLeYCjNUeP
QoKqejQQac5+v+q3bDfLfCVWQs0vFskf3+xrXL9zWLsA0XH1AOiYtzFI1f0OEv8O
XYVxHOdyaEwD3ynstKkXuFKuDQKgatLr8jaMx1kVbSs89yNZkayVytRhox1u3e26
ANLwQwc5b/shwyw75o/G4JDjrX3lN+yNb73HTkZs55IR0Ct5K0TucFIAP1zmYiKE
BQmvOphY06vZFP1WuZ/fp1w76uDKifLnAv/B1JH2tr6mBJCq77+lShwwo1MwqUfH
NQatrNiwncbL04AfAHsBj9VKku6To3h9cOU6tOXhC9cJ5eYV1CBHp33I1H+b+Uwa
vm/U/EyLdzO5IVgeqNTWq+VASzs+hzkTopSsKz8gAFfN6lLM68YyLNP1hkoMqaQU
39nIRhITcGIAMcH+pblU09RoVDykdOfSdbRqdYYf08yD4NhTECnp+xWwdIQQyQNt
46o5/kQzAgGqHRuZMqStXVIZcTHZpW/mMvudoUTFn7jX0CqWnB/akUlSvz9JGsbX
6vknP8uEFfLUxMgU+bVdZyOjCJ2HKA1arWNjeioiBJ7qDAe/dlsBve/G2VxD2vfj
bswU5P3GwhT0Roukn6jhaYkmoIQADxZahqVZhKD0QIJUNpm/51Q8aesTfPxe7rTH
GFa8ONHb8NmdUPufRPm2ftjdwqDwvi1eXqdWLtjaVxhWvOHKBEcJCh6NvfQczLsv
MbVkg/jxJjtX02e2Rg2pYEmIRPqUxBHi9duTtct3kTcPkbC/kk3of5Q/BSNYOGEB
xxpgcP25y//XtrJ6FlULn9DnbZzQfkMQG9UmHIl+vl+wiAzcB7UVAIincgpSmJpr
DSzmybLmh+2UHWYiKO8zsRBmWywcZl7xXFUGYfZV+E1SEJWAW7bm44w0o0SbZs96
GAAHOEAg88ep/jzeNd5Dje9eiBzEEOgavd9G/ZPcX4gfBuLwDaPhhnO/5MlhyYHa
YA8G06N2H9gKGfK0obotsJ+Jp3DQ3ZBmYDaujE2VldA96h2Gq0xxHxR/qqn7TZFJ
YAzVPd01rYrQf7BG5tx2FrfAYAoTS7VCmzKHpgJT2ND3xSt3RPRb+XQNPuZdF6kZ
18NTjG7E9xSR9t04PdxZwVJYv2zzuLjC421ECPba5cPowY6BOOIqwZYTS/FHJz5n
PmZ3dz7Yg8D4G1D2YuHIl32yIvEATHsce4USUJTz/IAJZYHdPp7KEIrLbJgN8p0H
IHvttc43650cgqK6wW4utwS3Phw2XWSKbj5hjztppk+j/I7G/TXh78y++tN4XvYA
B0cdYZ0ir56zTCAhG6/4PnAVDl92zATLvt24BG9WpQU8GbQLVcOIYVJwz4t3x3xV
hqBtIrjEzVXaMCtekaEyVR3NUN3GZlGGymGJtC00l7PsYFI6pISazqssnCTUott1
iGGxK8GvooY4W6UzGCpts8O8KqgNRvhpJfh8ClqD7DGn0XmXyjqvTVIUYjjqKKfo
GblbS9ZecvErKgKgTWjAYShn0jqHzgvpTPVi14jDJNgvYrUvqb5prkDODkGozENm
IeEEzyB5Hk6yUCw67b2CZs/+xpjcCRiLWeGXCSs1cbX2uYPWJ4vJZPJNerRaHmER
TN2XhYGOnyLxHPPgQklPtbrchE7RKkY68/IsKzpftnvGlN40XwfHuVHYWrywLaFy
LKjxHTg3+VoMruZKv+rFZBKFwaxLI+OfuQDgX3Kd/dg1x2NI4KwrDmt98xR8WXC7
WtMeRw7K8pOXYxp5pyGEq5KdDaVH1n0dkEZ18OC8+lSwJUOd5rNhqi/CeYIz+xut
Z0mcyG+ct8w6x43S0XdmfizgE8OZBjeZP9PNBIvHoVypmiUPT6vfWgp4a80MTq4N
qfBosduugU269pYutxf/aipKJcOtNRlV/Qm4AQWBiy1JslkCDuhmeX4y9Vu2jjou
qVvvDHp6epRDk2FAZvS0RDxEIC0kS48ATiUzbM1r6+kmdyz0uFDxFDW96jxoOvDn
AB4WNN7UxbeJMCjsykywc0htmtaquEGC6+UdhFIg4vmjPDTNX65Y5nVELVSz2ndB
y92ChCfCS7tu6axd/oYhIaCqLYdYqALfmQf9rbENTmWLFifOaMhcVntCS3JXjTZJ
WJUTsWykO2Lb2Zs11+lD0Pnefq8O9STjVO0b4UNEFBRP48d2F2e0oO6uYbFAImUg
4vZuOc/++9xijfv+KvFLJCgQXpky0U1jSkOZiquOvoOJFAjozgSYJwOTS3FOoa3t
twADdpCSWAGjyDk7efv0zQ+k8vV3VW7q9iDdp1Ogy0t1WrAqvQYBsWBqEX9GBuqo
fVNGpIi1PaDUkwWwBYGd4fgPnZ8rR1hYEZ61hsyaAkwpg4q5PED4jsLU6TVsh2/X
13HZGjplYDPPisbzzSEpOyxq+rh+7z0dX2Ysw020X9EOQClbdqkFUQasC0hRcn1+
y2oS+hpYbs6MI+qKw2t2osNeMQtWCU2R+03ay/mtrdAQAMxOsX4wikDiSt4+dcXH
5mUsoblI4QY5X/NbP6Y20hE1QJEs2otXeFYmnfVjBDffdSlmWbkvHMxIKVxZqwGi
FTTa6NBpsQUga8HLXrHsFrbw5YxMojT46Aj7vQHuvtQo3MyClcFkwCSpZ367tb0K
KrJYq1uEqjrxDDTov7F0qvf9SaPbWhLxTMi21Q2YQ9T3hFIU6oWwbFG+Tkn0R5Fs
8jZ6qkGxm2Jb93FX8qrTpRBe8hA+wongCbMjkLo+rjIpiV5YYp48gFm37K5wGezz
Z9+jwj0/wELM7Q9/iBcL5bDlacqMQ/VnyUN50liwLh3O2xCo5zMMDFuUNlP64MpD
sH1n0xgN6TBdCaAnvF16h67f4V+z2nbuQHBHUzjNqAsfoGSRNbNHMoHmpQvQp6VM
pau31FjYT6oobGdABezEZ3xuCOZUU28BxWTS44sm9emh8zgl2UC5kJuhGyWFLzs1
mUaIUUjONBYGKnX7so9jWTg29SFLkuG0oemIwSvlksoh2t2kvVh+DoR5iwAT+NUB
RKLwiQUUcLBoe6gLI6QN3fUWZIWjWM4FzdUX403m+o7nd+r/DGdKt30cEjNvlKAL
4jOupVuctPZb5ZWtfR/IQ8mPegoexwBtDEa5J+dAQBws8o9nSg/xvceC2xDY8K8R
KOw3eJajIQvcprcNX/3m0LnwtWAIgR+eeqU4M4sWp1ajrr3qhTEyVJg/vcocHaxe
3ckfNterd9f2+thSeUWWnmbxd3yJK5Mqe9Lvy96FWB9IonOWehppXh33TZbO4Nve
gM0MyPttVeAGs0/3LlUF7UVzPzVRQFILUDLEDRB0iF2ZkPPFIDANf753JWU6Fehd
OIJE5x6X6ibnayYKtwAz/gZ/9mHalS+WyO4/pmJDmGBnTGaCJsYZr8EaLL5X/Q73
Qf2WOJrgnZZvcU9WEwPWNCcoBFQKpE+VSF+zZmsMmNscXKJI0lYtxAZH/OEfoK9G
zCXxNbxPr9/I/+fbGasjCoTzytMlxVzH1gZ3mFApqjvtOSofADwGcpPr6amxlYpb
4nyvsi5BEtuIXbZ7I1KEN7XImCRJiU7gsFkfQzyW0j+T0wGGcSBVFwrTWYRrOL5H
38rQJLFVc05uSf7/oTdeqMLYuoVWPyDYS4EdO3aBfijAiM1iKf5Kwf47W5aaYMT5
BlkUO6JWzM0h9sHXfRbRXCbM9Vpnfc/XpXSxDk8zd2TTX5lfMMYiU+rs1nKOlqel
Hb2GYDWLrtb6yLWLNewGL7OArOqOxaYvNLwu32+I2TGiBs/BAyOBwUCgNHXTGb4F
FayDppsLYFzC1olE/oTCoR+5mY67ZX8rptjfdxlSSyHDe8m811Y7AZlnDdZC3HDw
jO6zGKDJztpGJClxNGq6tgd4swyhOet48Cr8JpoWesrpVMgnZhzmBhpcbnQQStov
cglEfpk4vuX7tSMC+tMjmk88S9NLZweMPdbh2A6UBwmaxqplw3P+0nfs1BCfCb3m
oEUkiTJcZ4PSDTyNJj8xQWaBaT7fRBmMaZIIWMA7CZr1lVFmsi9JpYYsx4dHyEWS
3LK2gQ8S/qJer1KJEGSl4ihNfYXNi2Q5Hkk2C72hCbeHjHBCJdhZfQp9F/rH59cg
zBkCgoJB/IeRE3JnAZ3GO5qCL0SnLKUAAhj9l+W7FgjJ0Ys39QDYnMJsNEdSvMQV
0YGBIaFxjz7lI+yh/AOAupqdkb4vDQpizlnKiSweIbXlkULgAtpacZuYiPM/fuVK
WgbuSKJWwl8ROWzWuWVwDs0ukYARKBp5lFHQCoqD4+HnVjokKZY5hVitSyXwT+Tm
LwEga4WFqOF657tmY8oiL3wEY6G4yyeLDpWR96rqdw/ru/bDEfCOHiCV0PuX9c+q
gMOaHdnoAu68PEx9JLJVd2cNB7QzgMqzZgj2EoFEILn6d1v1M+TkMNWNwGkUuNmp
26jXBRgHwT3INAEIF8fPsXT3l9WjtnXZB6UbFKXZpG1q2J1wQl3b+Zz9108eKi7u
m9XaPezVp8xBYnBlVr2m8hS7a5YMJxlLJZZVh/fvfUrd8I2yDh1sbfqeT/8b4s7a
riJHEDk4sKlOKMo6mNBa3JJekLxJMK4eVG092A81SEccE3d4IX+VUQvxHflglGrQ
QKN9++Studlbp2tVmjPyjUJhI7n4u6wZmsQc2RR9Vd/ZdFrKfIzJg1QPxW3OIrpe
wWfKgnUYe7Dyhi3MDwzF8qeAVLaSx8Jrw3hoBj2T80VvaV87Rl4kllYghaeXVlx+
6xUPD6BreHfJPzCjAlkwp75Qyeihq6dSxl9LGIt8VPHcZDDb4T4jyasVU8AtmZD5
7bkR1U9VKlXlDgktafKIq8537BsD/Kjk36yyHDO//f2AkRTQewJKJSgsVwqZtu1R
8/DDM3eTTTE5ByVnx/Ows5S0rxj0XO77c+aYM7Xkdha+Pb9sSTg7v9qaH7kROMcR
lofi9vf1uASR8rPXZWf1bBNqjij1ABlLmeq6O34ixtvvpo61hQjfQRS9dU3uX3IH
dibivoo825i8qWJSypxxd0oaxPtjvlaHbgRsL/flvS/SyA+MeE8NBK94JNrSpSHW
4JqpdGCLBfUqjtYWulFijhCyOa8Z5w5eSL21v88WlyDg0PApgQmHCb1d5XSC5cz5
EgHA2s2QQ8Ji2lg4OmdRyfMxhRtQNXS1HbObloC8q//dNj9bIJiAI4VQyatA1ayG
9/dqYqskLl5C4w6RQUFbKAectwQbQrnrKKi2b2aA9b2sXehQBfoXuhjzZqF/yzIc
Y0udSvWOft4LaQDtmB/RTlS9JI0xaaXrlJ0DsZ87aOjGiuO2ClI75z/DSxWsHeW+
9cz847ya7M6DUJ6TfOPlu0+0Hn/Vhaaqcp3c0/AH2cAQuXkxOLbzH+hl+uJhVBOD
dwm5CTCiHs8UdmEvh3GTHihOfE5itDSWlNhNFq+AwIXdAfhJItK4UQBjb90+DlYl
UjgzZRdZHostz+h+sC+SgI2TBtJYQ6wg8IMOfUu1qimBbst8yJze62IM1zUoqyFw
HxkzqES4o72Xo1f4ewnTRB0nYICxlg9Yr5vGQKwA8gB1pfyH6r//F8htGHzR7Flh
lIUI5P+fC+RgGUo8Q6ykoR5qktp1XZyE31L8MUdvtC4qpY+kqeguMe31uZWfGF4F
zIzZ4XdRzGzdOy3nDwRTbi4pYQPtNxXYjBqtNLUk69bnwXEamBAhFTW77bbpZ4JN
PrniSaK5KXCYTknm3ndTjwNSI+hjVcIVeQnl9cuzPKXxOx7D+xaKA6axK8XPRLOv
FF81JLzLXLP4XQ+oHxSajgKGCfc4jPVG082PTU4ywzYNjbeEoY3obj1TuijUbN9m
9aU4l/KGSUyTP6FLQ4HY7bbwpVgDwzvi2B0+EApU++eF9LMr/kjyPUvMhn0hTcVK
DDE+C36ff82dYNbwaDOFzaKrsENIlZs15s3K3RHAYlvu6JzTqZem6yKLtRUOChWE
Vdftw3jNn7fH8Tx0MissOs9PoXY3BvbAxXbGSsSys46bfgVrt6uqZDVt7qFZzcUr
j54LmtHPFrKobGeaBxgsHzYtC4or4n3suHmvncaa2SY26T7YcTY5rzgtpxqlb+Dv
MvdPZcddKBtDQP74pIr1/KQayMvXnyCKb18YfZk2kb3yOAhWceIw/j7qTL7+DbR5
rlllJvQghd0bUttohJqTn6MtBpJAwhcg6xy88eUtSSChCieVNdC35067tWl2SiOv
5vHCPVAf02PIARwTd0ov73tTT+oMAEul8VjX6o2hnN8V0mEYFHHIKfmiwYcdoQY3
O8yssaTmR3fosIsZly7CvXBKN8uhO9Q3T8x+pSnHjQLblQPB/noFGjFrmoEBgBZs
oLIBikT0iI6DLj7V3Kz+Gq1VP/jnbaVFNIG+7V9IBihPEkI2z6aeTlnqWTBrq9eO
CuH1F2tFa9QTr+oTUtcMlvKvwiA+tIazYw+/fKaJWCz/DBj/LieVLmdpnMJsC3Bk
au7DYTnSGHXz17z7R+WIzOSlNEUEKUTpX4vVLX1HTuqKQFIJ/omSwog/MFcqH4qA
eas6Fal+iRAUMXXhBAVHFVMQ2TuMNWV1YyzbhuSklGX4MoKcggQhOo1C/K7eqWXf
SWlWnBtN13hqYe/F2Xj42wWV8Y6GBQiEW9SozWo9RoFYnIqvSmXDqSZgMKOLrLmL
ra7JGvEJq1IKixQUkY3fW2tsH2i3SlyZqjZy73LUBIyh60KHuiPsDG3ayv9Wfody
i8ZCV0k/sFssT2nVdUGOArsfbXuMWmehNjHIQYyR+tN+Z4oLACslpm0cznA/Xr+t
46JVPsjLTsG2VZowYejTmWbIlsR1Rx1o1mNahrtc8EAC2ZByn0I4tgCM9kcDyU0O
QauKMmENGb1N1xntlf/2E/nx2mqaYbjMIBUl1i6dtWP/Gxva615wihVjfS4qgRKS
dISDic13AtFp5ivGWeMNNRoI/ylxGLTv0hOC0TNfD4l9KHf3WSydbM7T35MxO57M
WbJB5Sxw5B0uqmxOtpBsIZ+HGtJKNaqSrpKqQUMJRDNYLI2HRnUO1ZIE79Vg5LZH
EPyHWRL0AiryVGYwDhG3o66FwfUghxXFfwys9NHzcbKCELDbwuz7tKTv9GUIzzTb
y3GUm4Z+VyCysW5hrze0+qozTKojIfXPBhjXGMnxIdPcJ5DvUWZ3CV2Y3dos0a2A
bk/NAh9N3Un23hfjBD/3gOll+mhXGyGARi3PfepOzTSpeT4qic/7F88Yu1dxvnU4
SZrpCHRTaH/BlbBzEsCcfSNfthGHqEe/RGuuIGAm9eqV0XegvA72PoPATijkJDBE
W8k7xbjzqUr7PkxKTX4oAlGIlMhDcvvSImDPyLrvn2Grt41U5Au+GI9QUzdkXxPj
UTcC7F5Z/N5ZLnetuJm5mBzpjh4nexyryWxggS4jh4jwlplWwEtHsUdhNfVzANHH
/rXUYO/kwJFDX2CJ7L6vaW2hJAepcIaZ1YkwkRfiQBvdhQYJait9eW/J6RwW1k7c
hlHRaj8qSw5a60qQxPfPePX9l43FZBtrtD2znkL1nNf9GKBlXJ2R2YK2CRBBjY7j
TmpZwWBWxBNPiPzRAmj3eAKpDh5vamuyT1MrcURNJ0HGbNLluQG87DIeYFzs76Ns
Gn79+0wxJHLpWFBryhVaIp4ZdgJowGKZlHVjREXyeUP5F8Y/D1q2Ms3no5PFpPlN
3ccTY9GBfK+XM/fUJDi8xuxjNHqV0Y/vdHn/bpJOqfFepIAqxftMBFn0lOZ+VNbS
MZ6LeXN/4WrpIJ6S+JVe/nsn2rZDs/9fRM67qwn5TSggHbQ0Eh4U5sQrcufxHhlg
7DqRKD+CO/4ZRtyu35B6liV29/QtwT3HDGb8GwPvrulACLN4j6He0hM2yPA1TzzI
KO1fwRQfuDvudOnvrZQMi5toPmQ1yTpHIFLGE/74kiJmvjGMt0Kaw0f9r8/i5fjB
Nk5Vu43gJbmMILNNxm2jXBTkH2KaVxlVrDeCAxDWG1BwV2eNNOK73ZFTH6ETtXcn
Ie9T68+hrF40GANR68aWD7V4btTZ58noU5REfXMCjocQU6IZdXOZ/yglnoZMgisO
MS6zq2UTOYBSztGiYdm4AO9s8ZslsSOB0zZfYuUGkb4fwCQwQzAg52FTvSuaCufU
po+q/Ye3mmJI+7J1EN94RDMObyWu6HBzob9G5eUPRh8Cl36xe33QwbPDq9f9ZWYf
wF0bhfQh+7286uvTMND6oBtMRn/MxxddgetqjAUAlfwtvWq5vGdKbBZHTFm45UTY
ODY6hm3IuKZQSvgiGlEzDMoiW1aGF09FMnpYCAvqQ43fmX/Igv4zAhQVe2ixqaci
dx/FscNtgIySdXpwX1WZNpzLJh12Rn1Mgsdg8Zo60kv9SNiiQwG/iKF/ywvatdXF
ULxWU6EyZpcqzYPuv/jD+HKofGSSbfs4Rf8AiB6WYHNO2vxF8Ps/VDXaXFPbmHUZ
m7hu5PVzvK900eG97un4SFrdZvOVkpz8lmRDFgK8XmtINluft7wY5tKzw8+95Lnc
0Xt5yYBS4s3AFhoRPJjoUNsricVLapJg1cfC3wF7rn8LjfA6YTivJHIHscVAjGH6
I81ed/Y9UJXSwstgyfkzw2uYVw8wJQMbBk/7kNY0bKPQ4k0Wy5g6KpgHxAcOAXQv
YzRnz7OhwZ89KA1i5SYjGMqMDz1zc0Bb5AjHqjppwwRolJCIstKWFvbPcMnBDgAU
KOB8Vc4XwRb2UgT7qdgj0bnf4Yx/XIcru2Krkls3+KAf5OZLcTXrC3+f6r80zb22
BBChRCMt5rnzPvY5z7tPRRfYqSNW2GqJt9cf69tcGZYUmHh+4Ax8g8Zi7pxKMnq4
ftn9nGSyoz5jZE5TBicwq22hk12MfRJzUdoL79TL3iQIJNjjTMMWQ54tfcqWwgC+
H/ZcmdAWL3DBRhV4OPyQ6IaTjs9k+CP9EmlUct31XZV/11cJLMLc0BDI1mWksM/W
9hJRnKv/OoEO/iCGW4NoXtf2hqqzH2Xdnmi9f6mFGBS/ZeZfVgGXDDk1mnVa9L4V
DCbi9TfKUsbTLaS+0+NjVAyL5TSQR5lm3/OMAevoaO3pzAQfWQ+pdx1x/fH5FPdh
6rdiHZiGn6OlO3OHiatiHHQ4a7f3q9Iztw00iyn3qKWqQZ87LxobPBLoMppp7SXa
OafTO0nMyldbW8+zq6eUgqXcCoRr3WfWfA0M0NznX1si1YAclrjxtvwQWnrRgyGs
q2w6scq0kYtQPJbe5XpVkFPYPAGl8Jwgq1kxkDZO7yOKbC3QjzdDHLS6JrD/KJlR
S+x5Nh4pUKc4aXOli+DEaka0RDZTk0sIA1iVDogMyoDUHh1/ccOx5J2wpwiSci4C
hw2QJoGZgCgOkOas+7afJrnoZPoujj7eqt8h/AZcLUylIocWX9ek3AYxgpB6+NOb
I2mknMwuigXeeODF6s2TD0Od1bBHb3m5ytmV6b8RgLZbM3sfbiw7UIuP87jKTi3d
Pnxg7T4XW40leUgmuJ8vharfiFtZXF7NM7+DptyQkwhPGRHqE9v/0dPPwXWlJ99D
hr+3o/hR30DfmX4ZK4yh29mCdQ4scAKId8xBlKAuH+tPH3fLh5LwcSi/u2FLB4WB
qOdc7s3k7gZnFCAeWWF9romRaJop7SSSNTYki+bDcPMzUOaUX4MFAsxR7WuockWR
ImfQAELWGmg8ojy830RTaIXP9QrAE3FgtZBGUCzOLqUAhao93NPdhC9Xog7H3R9L
TOKCDqfMGUuNo45h+KW2VHlkU9LhamjV5cwlZDXG09HuwWNQ4jYVBNwRoxzyAtDp
N14JRhLUOgn5n4LhatL0007wgaOIPAEquXvitepYjO6wbAQwI1/Lu/fh74STzIXW
VNKoJ2HOAzw+T6ihiF62irDEeLbtXN9TtsDsRt8iGAWMxxrtAN67E3kp0vlLA1Oa
exJnraAEnBD9k9KaHvUYr+N0TTZ9qwm/RmLrs0vw5aS4r/1EiqOy3sWDjJTZ78qK
ShOP0K2oZ6ss50K9QWTJ8Bc7EGwbrttfRnA6Jr8dg2TO7HOWy9zq5DepXATXVmhE
uPCM0xS6OrtgzaHced36uF+gZoEfeYua9mSmuR8MkZhkbLtc0JiyU0MtgURaWTZo
P7Q63wkej5TxplhuGz8w8hlVya1LszLPsa/YWvqfzCMH7q8SEMWhP1x9HIDcwB3Q
38Z0Ith5EsqfQ5BE1MbBX6mLPp9jRxeKmliKAiw8gwlG2YkGIYxUjedf9g0yCDEa
m1j7ckL1lCgsYLldooKU+gZPnmOokIQhtNEFbvGUPBzosRmJqhwQ4nQKTUmwN27Z
waZWCdp+GdouhA4nMxVygXsN9ZO+5p7sNGKPVcQs5os+7JL76ESOC4oKBv5pFYpo
xy4Anc9f8q7wcuEZaHvmZQdUa0prLvfnbvFgylJ7P419LClED50nDmi6B+zZK9FY
TkKnKrg6tJmIoAM2nr4FYRb/F8qPMagfIBeMJRD/j7dOa7zEZPcluklSRMfHcHWr
8xGZ7gPZNmh25uGW6wWyYLf6uPtOtvsgxc4cV/sneHVBTxlV37ZW1uTorTIxEwbk
tNfJ+isQTzluj5ByIdE5rR0gZD16Ms4G5q5PTyoso76DqpS94QbT9CNYkVN2ghnz
B0pdIGINt/9hL/gfdM6693dT51hBh9ZRdatbsHxdxoMUZlrRCua5j+KUl46xT3s/
LqhIlempUa7hL1wXNqHURpoHkx4h+vVQCXezDpjEz04Lrs4k+mJoDb9H89YGpN/j
e6lLDXIe5w5db5MFW4WVqrO9cotSdnUDDujqUvl4Z/QeZnvwlKEvs3vlp3dB7jk1
Cl5znb0hC3A25yNuy8/Zb2heJYSC3TZp5pK44XxcWzUN+aNEN/AlADrHv9YY+JuN
swz0K3xKLur4HqUcu21uV86+9txeYD9MW5p7OZuC0ftrzLLdtxcS1HdjrbmnqrtD
kfQt6YoKJPSOzFd0/833HuRv0YaXPYSab+HcQvkw2rgGYcAsVJzZviFfL4C3/f4e
dRawPOEtpErtb7xkizVzJYJ97XD2e/RKxfdpzT5C5X8KYKMn1WCb8cJiJpFky6uE
yvJG/qgIlobjrm5MzMYLsk7dkp6EwIQJUZttjSPWD7v5afkFqooIWsT2WsIIhiDT
G9X8zFkleUQkgYRnp3z08u7fKNwDXFhkRnFdwJxUT71gY60xyvH7yVUvp84FZA95
i49DF7Z9yv0dt78MM9ADKoj02/5e/nD0AWfkLlcz3qQ7Jz6sAIMLMRm+CH9On3s7
49vgRjoXqR6+F33VZZcJSUsoXERP9f5MTVGe1UG0X+1ukTGmyKyF8NFhEIzbYBil
/rDosArusQTf1BNcX8gl4ymrj1nP/DMVfhkeXsfAOU2Zwix5gCl94lz4m5P+w979
46ivfcvwVnINtGxAEPlQvLxgfmuvkKzsp95AoxqO8cbUpv40uLSD0NbVWXes6rJy
UfX8oHORFfDg0ZFRly5JW741JrAJxOwUMUweH8O6RdX/8L74Enr3kuWIvs7Op4If
RTnTixrNa9YAVTWM4dmHNRaq6DKuDJ7qdiJ2pX6dKGPY6tD57+EeXe+sgFFxSAtt
WjrCUr417edaIV718zAf27tqhoruwI8LhPHk2oYVOq2eq7MROHBTonjcIi0kFnhY
H0G+EpSV7OMZ/tOmWB+ymo+PC01TLs3onWwqAXZZXx852yst6JZUwiEktTUnGjiN
GvY5I97amIlcyc7hRrKLX9hzuvVOTbjWRTiBX6aUh/ivOMSKNNEVlh7X93ZVAQ/Q
/b2ayvN3iP7QYOWFncpBANHwE+iJkSJ/SYq0Bj7dK4ztkseHSj//hFk9vtsXXUXT
wxQOuaX6bS9bxI9XdPfEysFoCOxp0RxNL5IqEgevaTYM3Z9tSKLDFJPvfos75F1t
Ib/g7xaat/AcNT9GcsdR5NJLPl6Up5zvmNHbIkj/aQUn9lZr4L5mff5atnxeh5wr
aGhldoRjRNTAdaQNZQ8zAPeWkqVa0HnSUjGScJaXO87bp7lQFUbzNyQY9YzHIf3w
OwQNjRgsyHysLVg/tvgkVuk8WzEeRUlmtnFM5CkJ8Y8zePq/o5AuDHCZLv8Dl2mp
WY49TPPgIevQ+aD1Z5TYWQKAl46qmibdO+ETfP4hwdD+uAuneHxmYYDE4Zx/i1/G
mhJCaqqw/QzYQzU++lXeccipHOQV1GOW+HpSZSDbALgVt/nBHtbwuGMgACkuFxwW
UZvIrjkWpdQ25DdHU36l/sH/o8U1MQSqjzXtuLhJ7ayfcJBIemk8sqjHetv/VNYp
2JLCDtoEPKtgO02Y3lhy3QJ8BYgAshA1H6XkLm3q75sm26wolHVje+AjLdJX+I8R
PQ27de8tuRo6W3k7Xq6RhFrzffoVd1/USF2fB5iupfTt83BpWhm7HU2dReXOhvdy
wdvtapt+3+Oqkl7vK0tVdfj+SqL3FXI1BA7MK1qPUHlD50xP5BE47GnsBxrLqSpA
e2fhEN6EYCmywz4hlQqiscijBrQdch9SrCE0ORaEuvdpWqT4/gBTOfEN3BH4PqDF
QzUYwXHrRn9qjAPmUbnanR4Npx6FhBbDkV/qhjo4dZI8VE1NSzUCGhvio1jMKZiH
Tg5p0KKQolTvzNpTtKqrA4Dgs7LoLXYPcgyGoX+QVWYGz3M9lCLBjZXiI5KrngqZ
/1ObH9VZKhmFSXsCEq9rXzLL2nUhywN8Gw839p2DDNi1xOIqvLkPdocFssmDDlfv
0QDtJwrZE1gTeKlNE9+w14HA3uMbnN36F6yLhQn1PmQ00MdTXzrBe5rSTFne3AvF
S4P5GH8NvHvFxlUtWP58QeBx0tUIQxgwPKOFO7lp9mgNZjbLeVUDk9fqC6Cpu7Yc
Gwamdtv/yUxWzseZUOcHDKAUGUxyyAYKUabOx9PNdNSpD+qe6FGQ7HJHffvxX6gC
1ZiiCIvfnCXV0JuPNCao8u5jwTYTseXZd2oz5ISw+n9tbqpOt775/JHNMR6NyjLH
hQA9myJ8SHNTZnsF7z5Y173nE0EDrqX061bselPLZgk4RdK3UoVjHDK1wyQMzHe3
JFwmfiNE1B4kzvY4i8IGkV5kRUtxZdNe6EOl3ATxOc6EIFRAP072MTNZY/5rO+3t
zhkAYow/uyGiUuf41+3FKtrkXH1Ckd2WRuMvBEzfiU91/0KIeDzbv+1nc4phvP79
P/gVf3A782SfoOcOyy4yczZuTrrUubbAJmUQz3x4JdtFW1TO2RiCgLg/z7wVNrga
HCYjwY4RuuS6byJRU6ipEjkac1mZHkjcYe3GF95pQnrt0+gp50U6IKx+qE9IH5In
+zIw4wXOsD0VibxI213hfQt3QXJaxTdzkYJt8ujShaLgner65WHNCwC/YBDs06PA
LgV13qdIQLpO052IVoMzW0nV4jk7SGOfMnwW0/bxauy3mXJwY7vlXXOftDEFx1Kt
TX8JNqWp+qfz2C5s3SHx9VQoKxQw2WvtXE2YownQbuDSl5Inu7rwxuLZySEIFyCq
cQtw5BBrtQN4n5hBDtS+BFhQYyAPXLAYEQItki+o6uLfiV1ln2mp+/zmIK25LCtI
LoShzGFJrfKu9NJ9/cYcLLaH2ourWaKXYm1gRlLTli9A7Vdo8gyh7y4J3O9nhyrY
3MYooAEj+HGf7tSfKriTG0Hjz0XoLyN55e8zQSRgxyvNtOaIdymLsE1ckwQPosVp
0mvaiLe6O3I5mKTY8uRcSmHF+AuafySxtXwVgk+eK+hDrozoHMhwHm5JOs2dFIVV
0UcO5g3G5gYe85JMmGv81Vk+r0U0YLZlzGBaVI64Ed4xiMsVs9pz9y5kv+/Fd49T
rclYHxByTHwFWH5r0pCS0fzP+l2UwCex0eXWJ9LiYx9gfXz+MIKsl79gl9XCQpxk
6oUPdOTp2RAb8no2rB/Pv7eR7g0YxhWuutOj3FdPFqRxVMIccxT4IIDraGv903kO
GFQFpKVfPWhyh8uvd+E1bGqY6Be+blM9MQSQgLb0prBQjJMQisNALFj1otUr5ZqW
ILvuMa+W6+L3lUaMPTJ0sdWeH/rGwYxki3FdFq4T7t09aNIucSXmu7qHjlUxBpME
qsSIsvidJjlBBac+2UUNxXYAHY4//IsMG46Mnf+IhhZH3k7sypEc/yKF7rT7TDSk
bt7M8jL7Hf9DAGiHsAxV9jPypzqXhuceebrOAV93Rbe+Wwj4AEVgVrEhmpp6V/wo
1cRFa0g0zgxnhGXyTIE0AFklzUQ7Xp96xaGCdmOzk87UaFQ/Xw/sMre40vK6RM8D
QaXvZLFufVXNOdLv/tzTjuvmD2VnELFq6lk465TWyOMEeBwTSU0tZhiuJ6fhRi6B
2W1Jid551ELA65ecYhywKXf4ZrtdFV3/WTShucy7tkTOkJQSu+PW1KRfIIdvM9rv
TikwBxlYUZGVFaKKa0cYrrZoRHs1c6qIc1Y8rG6wGT4xM6muQ/mbktukp8VD/+p0
YAviihKij4vsu2OJEVXRQmL6dlU+F4xTTThLnUXqRaBhTqbzqOUy0wuF7S0ZGkBg
eAXBCmwEaX4bJySGvK9IZ3ppYHdp0Ul/PEJeKgUwbdvGl9bp72r6OEftjsqhX3+2
i+QesQdEr7Zuso3thhfx8NYoCOu3HAWVZ+d/kUaRI52pQAgHh/eAiP1HPVry5S9U
TW5dlZZcpbMvsYQGsXT6w1lfnUi0urrhvo2wnxEiVOWubYXMATO5y2kr3Y2+Mrca
HQjcbQQwcU/APAKKB/M0DgnB2xl+uyDyzujImeXCT8pxryE58YrqnZl4ss8k99xU
/XNG5/Ln7g//JttgabYIvFSENZEylTqvt/m/aaXwISOSE4OzgeCLHBTxEz6gZ/f1
HhdkCD4LsdRRDLUILduOmuhaLS6oUYS/POldXNxsekPRuykaBwWxLtpWKOEAEyA7
LbI8/HOH9Q4jtfWPYJXq5+fzxlG6XB+9feX+yGy/iU9fQF8NcRFvxSmvzaJkS8qc
J6VHI+ImV00jAT9er+kyVkfV4u4PCwpTpFjMYhqBkYJzROUX0JxlbjsSz0BPT5D0
lpH+mDq4K8u/7M106pRpaPl5brttfoCwyD2TQT7zlfMRR/+39v0yeAOtaM5h8Y9K
49S5UPBAPkMPUU3m4s9RIskZsrDFn5XZCqbFASkFMpr8O70CBp74UGuHfh6lqopX
xK/GmE07zWVcjonhJ69wdG+Xe2pyHPeWI/30NJGbAIlN2lqklG8BnRz+/m0csQV+
f6qCpiZCh/DtnpRV2BRYhjokXW0IoiWeVqC10xjDjwK8KGb22wJB/6fI+di/NmVY
zGaiTgCc76ANQnbtbg8hPHNPyyGtEYniffn44asfdngwNXxfNevgPjVame2IspSm
2u9EiIx6fRgeTdUg+h0LQupgTnT1zFIpDLiGTD9Fv7XfExjqICIIoaGtnP5n+y2Q
NxsUEfGBcg6jCWwurU6LNOmrSP5uIS60Ku2NmsYPrXM106J21cY0kNeAEqlQUQmW
tiG25ykBxnBFGgX2jev6pu1aMsQG2VB7w+jbYCklPyeOfxL9C1w7UwsYS69IdgV/
uxuGjEHAheHJxp/zPJNRkHvQyohP3CQBMGjEgB5DKeBNK66R3zH0R34FALB44+HF
spu5bdEcNRgM0IF1OxkMjDgwHHEbnPXOJv/fDcCbqdphuWeMb64XOoV1znUdMSZD
tSCB6M/bNpqalBis/IZ7ALfBoTE67YcRndP5+OcVFNX0uw989pbZQbVxqAY+EhvT
lwKcxGV6GerFZIq+eMQD8+T93BbYRho1iAVV7okIvpTvpsqDfmpljdmyZzLmgch4
2fhKSwyZg+PVTf39fnvyJiPxrN+3EdXVsF20kK2MeSCCmHwqNaKl0I6SSLcSlR7C
nVpHbFn1HIczrZ/J57sx2Oj0nyhwwAfmp07ffniQ4mZ3RJZntvUumyS6bpq9Hop8
z1xqFslyz7D/T+f0a8fL05isuAXq6HKATqWtCPreB1aAtfDIEKuln8IOGwLFfCfO
dxxmri4Tf1meGMHjh2XR4uqSDzdEllmS+8inTF3V8MuGmas72svXY5Hke8Oa6ApP
LJkcQdGoYNuoJqUBLIcNvBREGBpCr7oOCvQrZyLdnoQ1oqKhRrgNtoB0JyTB8/9z
mLHhS7+7bVCcvl06eOIyGTx4KjfGL/fGc+MeXR8Dv/Neq93wEKdf2RyUNpywiTvf
q5SRNKjDT7AFnApU1vSf8ckzs1IudD0mAq3t4ZpMXHBTR9wCvtHKYDFAwXTI7Bsp
YX9S8JQksSKab5pqMv5Uq3cJrZxFwZFuYib6A9RzJy6KEtKfJjxQhdGe5L1KzAS0
KELuQDYnr/UcI//7rlX+KjZvLiHSTJ0d2TqwOaXUpvcbpGvs7B2XrRpuTOqBIcHJ
AbOTzIPDxvWxTPijaCZ2IOQ2GuYGVFiQFoVPqb4wRizpcCRqPqMAkCNsRn6WRLmV
c4NKWqy54nttXJYBi5EdHyxdJH06xnMhb0WmMl8a7h8z8RIeF+MHYvPVQ3B+Dw9T
5+P79eIv58G9MV7NI3VOeZObNnbMm+du4+KscDehFMgHI82ZaMF9rrwEt1gZWKTl
nPd1TpR/DNcCnqxTRVplS1olerc/PuHuE366In5yHRRZL7KNJbqpAj1DHtdTDNhG
vna01uH9BaqgqK1DfTrQ0OSkl7iPmrCSKUK3RbfDlevZCyo1mEZ9KnXJr7xjlLOv
SoMb9akUMmx8f7QMr3WwMIGi+5sRslpAF1gOPH3K/GAWE8A0jhfuLKfJNKhjIALJ
d0XIBJXNZbCnC+7QzSBl9nSR54xCImF7KGVd+/OxDCZmAroQ599tSgBnNmdGLKPE
81t4VVmC263G+voDX2pkYb3fi27RrBR06QVpxFMj8YfC2h1HnAe0gT7UPMUkFotS
swoDygfyqUNDNGZo1KQDTkQy4nvKqEV/dPNUmekxBS3zg14FFx0WqHFsmv78CpOi
bH8pErLof3Wr98/2QMTyl0HF4gz7wJ0dXS5cyyXTTcah7SsrX+IHtvtrn3RqAryl
syOKex9yf+UhghlusqagFG0XEqNlUWCo3c5xezo74DZujzR6BO42OW0X8cowpDU6
Hn46uxLDqT0FvKiETvCyjZcrBUyUrwOmOcFttqewwbkJsIiW7TCJVqa5rv1Ow7xQ
xe9tTTHaxIiLvUNga9diYslPBulOVj2XneISBsLOvw6ScAJMXG2w24swLtwR5YA1
IKMpcj7eLaJP26Vgf+TzENI0UVHXDoshmA3ybEmPnnUdms368sdSbP2Wa/PYTBsb
y3DwJMlqE/ykoBzp/TEmIvJOgP8mqgDpPzu10ATQXj6xJmt3vc0BWlpPUEsqb55a
ses/uoKCrQDO3jpMQkSh1QtbUpehbiO9Ze3Da7zH76Uwl8vpGkTtyQw1hBcADyv2
HYw/q6fYDEfwd1/7H1V44fPztt70r8Z5fcFfFQmgbeweQH29bAO4F+j79KHIN0xI
vEUUTEAYrt9iw/p3EfIY0LdD8N4JxNdkvmhfgfbCa3x5II3WwyRr59CFK8UDZnw+
fK8VIBUr4CmVA81ZlOzYuDJXM2MGh0CuqQ2M+UwIjhetCU2kokL1CuNuyhEe+FJ+
b0no6oJwWmI1nuHhEUFt2nGNyz3soKH5FRuDJgVb2+J3ajGIZ0OuzIYLFu/GBUlE
GzRRItrViVdK+arl1mpqJSqjFnJtXijAIkM1exz2Jp5FsDxzOaDjumEp+Yo0YoAO
b4ztrRTy7K1+WfeCHv0Aon5yN/VALBZJCzpbbxD2engsHEEiuoWQXa9JckpRGCWM
TXYYDaqc+ewzaTsWKzgt2kb6OMMvYJ8xqqW5ZWCaliw74WS9sgD0is3C6ddSln3S
M38bxpovi54q8r85bYjujX+vMU6bKZ852tfjXMNIn/MLSkvxIXOhZCsZjFULlPy9
CkcGc1OnKMYzPUAVZvPz4l3IQ6cUiB7Fu6IVzSOtVSJLwV2bxZoWKsh9KPcn6rNe
KTRzVKBHP1DwCy5PlSqbdTDLk2Vu/u0TeHAmLWs/vhRVSC7QO9IiR7Thm3t89ADp
U0YUB3MDHWS53pVhF+/3jWF9Ux5jA5wGHCZBUF499sqGu521NdadNdL5bhe0AIuH
BpwACaRovV57F3QpQlxVrjFmYM6V3reXh7c5BubHgeoiIvbXpPgo0LfDrOmFfDhc
6g+uz3DLMtoQBTSDo+L8SSENpkXTmF7ugoi7tV6yP82PE9kTS1tyis/1KsxdV+Yr
dbWr8uprcVy8Xda9Y11jdqIWyHMrJAB0h8sESUM0i2FsFTJOy1RvgiBixC57HZ5N
KfwUro/MFit80NBx1H+DiUq7Gjuj2HvGYp/KlG4sf9RxnlcIgeMht+mjle14c5FR
P8cFtAqiRwEq+eH1CNP+JF/jcM1kobjXjE1HQACuGzzo6cbhCsr70GyPxqmgIZ8p
MKo2klKTVm7ab7Zs3ZPu35X+aHCG8AkQec42gJU4jzX1yO9VexNkaCZALfgYnyp9
wF+/IGMQukh95V3x8QnK5JbDCmTKhOCHJYj3Cie6OTpFcybvzqdb4xT2n0ZYVsNH
bfgUWnO17ZsZIiS6be0mOMlqmR+hvla4Oanu/MZHt3mlgyImBPWrFEzutu+1Y7r5
rH57er3gKZiYAev5oJIQ98Egw7L6QoacRRVdwGvsKjmmPtqLDzIvBAUdKEsp53k/
ol+IhvniQ5+MW/iSnz8X63XQOyxAksDucp3CpeH+Cng7G4+49z9/Ss2SnAHCGuEc
RjhGOhtO5HpYlBjRIk4sUYCQlfgOjkttQGEtfB3+M68d7xCPsv9C5NUqdgZIpdNa
dTHqNHLjNI/awGo75aHOP/CAgKVagjejjiozZfl1a3tRWbB5YVL6o07mXRII2XgK
wVwce0R+Gl8FgYShyLx2uGSBGNpuLtLOOUcVjHNk+nc2ztAF9/vPqRseUn9TmIiO
K6DjRqXpCHA2MMmd6FpKQPWZaR+bFVZH9RwWoNGu2Fnxd9e/5TCxF1d/ebidWWrx
gz93KzGa7rs3276EhQ5i4JbXzetYKqwUIQdfigJ4tQ6vshgoETuiw4gGW7EnAEjl
uhjKPalacf4byBTxQJzYzwEnAUDtJ7t0Z4TRHM8j6Z9lPVJwBffVxDn84eeBdO7d
ecEEojmB3qqtbrbZ74JzxGstn9GFCuLY82oIQL1ZK93HMP1+yUZfoU64TSQ9BMaP
c4WndBauU+Kzt/fXXAcckaGL+/98BSzmoWZhwkfSd1li2B4iT2Lk+Gb1y+NW4s4b
tG+y8ReD+N4QfKkOcCKsrnOXskqWlrxn3MGH1t0CHG0oV4XQ8IErteyWuAE4Gja7
wxDUd2+5xtloIBQOZAWpqf9e0SLAM/0BPF1hce0W/M0NlQFwpN4mLZpFQkDKtLZd
nkw4zdGrtDwS+0o6MK7Eg1eegMy3zwxHIUbtJ7TeeSbiNaSiKfvsyHCMKj2qjX2D
Rp1nuflY1UgY4QC6zgaNlXNpSqtc3+D0jf40lOM59UUxkvQWcX7aTv9B/dtxH6NS
AucGisdZGOpDnX0DUJAls30zdGbY8xTzWAN1JAJXLfcLf8EBhAx4EN53eG3QQx5z
57AQ4vKue2rkSnEF5Kaau62aVdG9aZA/QMnnGTP8AsmChoNrwmMfNJBtqgE0oFq7
lCKJZog9NUDmqTWVp81zCkAEjxGVTU3DZvRItFVAvwCXcJ4Zw5xc9sHdJTEwISJM
0NYXQe35k3Pwrc9HPvAYfFmYQv5DcXTRwTPPYh4HUq68FM1rcdpOuWmiU9JBu9Z3
MwX6wtNKLrMHu6hASR9vYPD8efK0122MmcIIMqPf2wriegWLJ2hUjJRPT6ownI5x
WFZSC1fzSt0j553CxqDQjq2KsKB/n0TQDJjn1BkCb+ibxSCMT/V/EusW6r86ey7W
56xI/ltMxe//oVabpr9WoIO31Iulwuqdj4vQJcYyp44a1h8HO1CIstEv0ky5Vlsk
/SXEFSIv95Y7nkPVOgfcwLTypU7zzrhMsyHfEEuEDmzM9UIuozseLIdms6qbxKsy
+ZMMkTjNrhoJP29PLXEDXmSga4BRF9kQpaQe4UbhYRzN8E+FN12/rFh3lHajMZb0
CyoVb7Bw3OtekvNdSwKScLzll/QE09M6dCM05BE+7d1GEMNGZTkFduLbgE3TRBhp
ig3dtBJJEdhbFVakhY7FV+7qoVfZpOi2cxxzGQCDxC3M/qHsvXvWhZpXyD1N34oj
dBjCJu+LlTUvXVfarMz+dJ299z1ECcxF4YVPAmVgX6W9POlAGWFED0X9OnbSGCkh
f3m1dXRrmW9z0JZvB8aRPGO+dG9YVEEKS1DLOJfT2a4vVn4J6UjwysOJhSOFJuRI
fSr+OZa6hY9SsrFKE1Pllb9i4Z3l8mcO9Jo29Mv/8olOOixEd+BPeQA16ZHKQhNB
BwUEHA134NInT4jou1aopXhWg9elLHre6TFzYCjiwLcl4dqD1uBod6reS2Srl8AW
i/t2BeGC2tnBMY+KsZjm7DcPfgqsp1TW10swM7L+YJXeEBPPLB4zx5gNy0I1mrVJ
0f00pbPZLOkm+sgYxABsfsPJPxgnutcTU+9xJRSnFcX8Mtui96gmpmP+PYLntNAg
E67QqpffLQ7r1jBA+gL9x+tt9TC6KrV3N2OFLF4HNiaSnQUUmV2RkVrbjatwjpZB
o+divk9sTufO9GmuEO5EIy9wOsZvMf3HSpdvzUtvTxtj89feR9NvIOb1hnVwzO+k
8cZNV8j+W0WelGLnrbwU07/hQkohQxbzlh0q5ZBnAyl3QYxVUewYHPLuqqBUejnG
z4ur0uK5DViv1LQbaL5ISwfA/I/b7sG4N6uPphd6HcoYPhE7zEjgR0xlegw+rjfK
kJ3AqkBjdcBfhCLEI0fgPSOyZnStknq91R+OhXEVLolnQRFigUs4jabWaMSj8kjv
wa3+fs8rylHB65u7fm2uLddKwszcico7SRoxCMFJW1EsfkGy1e10lF8XjfRrpL9n
5Y8TOgubK1Mp8C8EzCckUMcEBhrfkYkI7mgtHWrhu2JXN2nB9uG1nYKBSZlO8FpK
gTHXhG79tzhJx1OY9ogmqJuHMjpsWf/3/dVT9CYH2VjYwSWF/XgfNDmOB7TQG2BN
40gT58nJ2fPzaWN0d0ubeCTv6Y3J+Gm1nDHa5BAKTItUWvxlctCe3IR5haEgg4Tk
AS2bTyOD5RELG/IWQRzp7jU7vSLtz8sqJKTop/sYGZRNXe1106fapir9lEFsf5qX
XFTOuBggWo4liLpbkVKvYV4UE3v14DyRVvwh0vmYYfjdLbQ0//i+utzW/d3KffWN
BqIEvSY42GaZUssO/cla2/NSkbec0gl74XCwhv8CuVZM3a1AohMAj3gVRdqsMRAu
R3CBBP4dXpNbO2tLPcD+wwJwmK6Of2iDTaFYhISe3NZaM0aRw1AKj131HPQfQ8Rq
1qKJlEQiaJC4mO3x1cwd6nXs4LJXYJh4mwlqCEsxy1sO2RknGssf626Q2exMRsBQ
37tlyAWp2GJMG2qZXXFqLICrG4ch0vioylMvpVsjCwa05oEAfvElBeH8HE3zRd08
wZdFnaiVeWWb+Chpny31H3wm12t6EFhNm525uqP/2BxdoG70wITDmRAM8NAToO2V
ZBVY2fiGfbfSH2Ixq7qwk5Y1XPB24KDzmLhFdInyKPeV4JqH5SXXgwdtSsN4Xomr
rZfTXJmmp3Zm/bBWCMJlM3v7eSIiX5U2aBeXEyUH0jWOqZUeudRwI07WOiJy/u0Q
GaK2/vq9QUXL/1ru7MuodHTPPgxUhHHasnNZu4cg4mXh5M8Wt4PtdgiY9ngbtZ0S
zjxp+Av/HPj4H/91TQ/EKWIPr43CybLdhvMhlKxmd7Vn2AKB3OyrUquwV6cs15Ox
kMASF0YbbvkR9a520JBgnSKMmje6/uvn3sun0vG2fiJZ/PCvrB1VDKUB85/DSGS8
Km5Qj9IolaVfiXRphXTzMWhdU3YuC+LwxuuYScAiiBpVLmoohsOwIaSEh51IIpI/
tIVMgj9J6daXZPzLOCeYDVTvnwOUG9RfIKuDd2fclVr1+6iLzMB7Kqxt7HU3N9Hi
mtyobWh4UDfsARxB2YlJtecAleFhswOKzUAc9TXDrREzgEQQwaW8163Q8uUgh+ft
TzEYCRocRTw996QZ4aNfk5Xa2FNVSSbVAjbjHrtut5gri0ZEwiWYbMiMTkuR1xom
JaweikAi9kcaGhz9ZpXU6CW+OvDeiO1qJiPFRbmLVufYnEP6Pw1wVs9w6DN0E1Mx
sODT6linWhbpGhBp/kKjTm1y2yRoKFIsgpfFna3c2bJgL1dWbJAd0NEbuXMowE8D
b/5YCgtLmPN+XckOQBqbU38be/OrZdWyaiQDAV1+5MoDNfZs1UyslIdiiJT/+cg9
LSMRMqiAjD/GJ80F5MsVXqsFcHFekBLmreGII94lfXKSuU78vmEKnJ3srQhohf/L
92tNt/mNJP+dsCPyeSvg9pR05k6lOoZmDUH3wzxN33jZNfWr78lcM/SgPX2vWBCH
+Oho2J07M2u9kejGu7b6A604yEivkWUnKQ0lRrq/o48hHvxWnSvDjMwoZJ7V4zhj
QnZqf8MKr2LPlJJRHhpyNvk+BRdt3CeZj4ADFURjbIhmUb/l/BbI+72rzpHVP0Pm
0dTS1vZbfPBq8NPdF0P/wQyuINlLLlwX/Kk8h191AEuVDfXpBZto8vxwHaInZPwH
B4QAHUbDHknKqGTMg2mdv1NFU1CaRdz5lmEcHqfPmzZmaM0tEVS2K1MInx98HRfZ
ZcSYhKNoVbiM7XeIExxB617innChF1qjbsSWMlsYVD4WbTnpqRQvVuxoHMum9uox
cuXPoQuCUFLF4dTQuxx11Uc/zkpOZcvsCAWVwzqkNe3uDbrxeojCjnWQ7kWN7T6h
UltzNTg3AQAyn05lQZL/gjVThM6nz52zTPZEZdBH8+o/0GLzQMjISas5nS6Yzbsj
gGFh3xjjLH7/5BaBXaaJ21XFaWFL0vWseHAmW4q94PgxSi4eSwBPPg/vfvolhSQT
x9rQbBU1U+USNvzSSRjytptIK4RLIp3IFs4C8skwNlnmtHZvWY4gU68Zcfoyb24/
QJXJGggQp2PiO7pYxgh89He1tBNX1gc2gZ0QFq+r87J7OlssX84hDD2GiAam2Sa+
/qLOB506uG8Z/QCu332YDX1XU4LxaLJK9TJRGC+I3qFmgzKWbro6zXJdHFTa+jFn
zVK9g3BY71R804A5OCQBN4bltrfAIJVxRL5dG/1chwhAhAro2sy9ZEYXB3XdIS36
KUibaaMLGrSmp1+mCIn0Spdwpc+MbFUfUJdjfx8ua4ZxiLPR/5hL0IcIRfiVT24F
UKo06Onqf4dgDOIjTjNcH7lT93HdrU3bnWr/049BcLxOGtbPNc+IcnpDMTR68oK+
sAINFWIkmAVxr2Hf3FzjhaRb4sCtjxgGh0AvCQ1MHOaA8UOy8neGxBJAsZNPEeEQ
rs9+KXsxNpT5kKbxBR+UnOpzoBy/k8wVDyx2bc+TaRHSPRC2FHSoemnuYt1NvbE1
/aepO3hApjPtEsRLc7s3behTt1NI2xdMC2q6ShZr7Sa+NbjcXYqAeYQ6E8uXzBdE
zVEsqRMv7vt4TEcxXSQKUAFpHI61PkvsrjP52zUV9B0FLu4qbbl1LXOKgtbUvuC9
cX3b3iY0RjvA1ut5XkxSQiBgWTOkriewihYl/giFOtpbwx8WbpGpMAoABSaasJSZ
qCO1D9wCXOzDT5fJ4Gbu5VU06WckLUDjykAgMtXxGBjzt3Ciyp068eMfE6/cx8yK
/J3f9n4YJuqfavvD4+qR4q5BL4UhMjXr5qACLG2isguu5iBKTeR4WUvH8OPWQv2H
0+BeHqiPJSpq/P+nZrpEgG14G83ygxt7rMm1mVgGSw2vSI+907lup9lI5vZmuea3
rVBYAnH/mxCg4LQwELh61oIjADYyGq4JDjtlF11eGryNcKWjQSNWBYQApoDgg31v
OFgci75lhwuvxZUiEAjGbkBrt9A/gbJ8diKfkvFvtzE/FYHLCmTpILEkMW7chYeG
QIuwGJw/Vr7j9PGBkavG39zdEssumjyT0ECzZCt/LjwbJIq5tI8EZZWoKg++RT3X
s3EVl2CCkFH0gz/jq5HeHinYryP2FxkOWCVPzoSrXGBb6gqml7vPiYdquyHs24P/
IneFsT736/cf+YmkcEWym+aqqhrrWsdoq6YMC7/G7fL9kgIVcmVy1885GZPvxFXo
xHkZIgpRFi57Okdenrt3fBILmLzjqAnWVgX08c7c1wtNCpzwgbxPCwwlaCQlme9l
GhFlIWFy7bU0AZchw9QsAXSEMWMRJ8a2aFNzsRUI5gRyGdJNLAeg0QlVCfltylRf
b4U264b0MliAHRjThwL//4vv7ET6LOoUSFNkux2ZR74XblPrFeGFnhD+Gj+Z0Bz7
7b94tocBO3+LnKyNO09mDpPjfbk3bnY0jPUI9pTOh6KvohThNXzlLxtjX0ChtAC4
xE1pSNzu8BVVHO2ovfKmzIeXa2UgNiySJ//+RELMfkwk7ZvG9cFRVbVqOTMr710m
inf0vLUJMHvGszMjgkG7AV/T0A07k6rJT3wglYwWSzkMlpyPadOBu085+EuV1Gzl
YnmOTeLcCHckTFcvLwXpRubRJOOpUtLh/yv4JQJyP62/y7eO/LbyqXkkU9dNp+Rf
iKA8DI+ylV2aZtmvy7EanCiax2yVpoIvZ3sNnBwmciWONsv2StjBUVUnvhyxo9ql
Q5hOr+1/blkwPA0MqMVYBwhp/tTwYmTA5DJEILdyM9Lh3+CNe9cMIoGFBH/YiWSL
WVkwChR5TqWiwaevNwgb3pYsl0gqx/XW6CaeP+6wFzNXAClWeD7iLJhoam+TGPhC
eC8JLW1mzfSbOIYDTMKgZWoGvVfUvnPW1oK5GRyuh+uIpdak60TnCNy+2ekv6S49
qLo1u3cd/MnIzumqVOLVcKkl+C23Jd3RA4PGhcvkwdvroeRe0DWzwEHXVFR3+SwG
Tyxyx0QmlGJshb8J/3IaSL2rdK81VzXlHTweG42f5PVGUehsddAO3sHW+bZtVT5T
IJhm56NtnVg+PbkLOTa+hgv9XzE6py5rXXcATQk6alrBDCXQW+X66Su3ecuOIKi1
6fE4tLJjpdeIea5j279X8Io5qt20dqmF3dRyXrEle0dhbm1x6WNdc/GKk8F2fonn
IN5j0Zoas7x1Mb76JQdVoEFDIM/ST2E0UQZc71EgIUNHbZZdasiHQ9ou1glgRmyP
PA6RC9P63tVsCDdHyjp2tdeaNMtpESqDhGDVOKmr/UIEYp8Un2zTNUOqaS19AajD
2urk0V1noWYrRyeRF2SoEIdlQvnrSHyTt8ocm6LOmUWbcDLT3Oc2au6x2AkmLKvw
5yIpl2vyZi4FAZZGmHEi7O4D/VfqRA+ldMCQhHwt5uVeRz2xFn+Ty1dBP5Z3M2Zf
HYOkyT0kEvfYz4tKbhAMS6vA5pzhQrX1unrbm5slRM4xI//6wYinMqSM2RZKqfe8
01sND2RSAeS+yjUjYNzJzfeglyywvX5X3cqDGimAWD+NhGpyC0Qttf4iPz3PtSrR
3zDdKOhQoRxYWAFx5hfG0PJi40bEoWi4YxVeXhitDQqBCnnhDG4KSf5xmnIJrnZ+
/Y5hI/9dH8MaNU7pUj7HTQw3sBj7aBFpfEu4JA5EIXh/KBYGFtGPAejH4e8rmtyW
dzW2C6Azrv7bKnUugK7AVheonwzAjnLRN5qz07uOq91ZdpS6B92x1cdMbjE5MBks
MximxvonnzqHvl/P10soOV6nFgdlj96GlISukxne55lPC6aNvPmgLgsIiDSIwdTv
OY48mT7EcqBg9+vJZYPl166/OtSWyMR4RV4p44+6zsGhPrYiHz9DT8JDRk6p28Sh
jT5tARf3CngoIBEsVBQmmpKdBZx3OldHoWliyEruuetdMi72SmZKXj/2iOLJmzmT
/Y2qNsnz6zUgbglUVDjRkjaKDtkGbes0EY4cKejCjXvpTqBlCwIBoNjWfq0vOdQM
NGmT1J6sGldS6VHT5li3RQanDS7bgLEAFhsIinXYrl4p3woF3gmB/g2+nYOr0CqG
h1RaE4bS1CdemGKy1BNR2ZoCSPgUneIWjNm2bhMQEMKVYuzFxGRnsfEuO4i6m4KG
hgvppmhRVov9K85qKs4kNPjvMU78C/MKQBAAjdBNCWJfXzjK9NOh4hJBaC8oN6Rz
cZtw5Qzt0/c6KVhJmFF+qJytHuNeqwIKKB1zpWeDOGx/tbslZkljdVfUxq9yl+Tp
8NFhJPk0pSgzqlBDmNmGfLpd9KJOT/ZrgH805gur1j5lIBUQ4uN9nXvZysEHSN6G
bJErQNtfu9j79rqyXh6F6ox1Lkqit6ZSfuqc+US5NiQ3GJBnBvGmUBVeoSBKmP3l
Tu+f+DE/479SQTCyS4Q1TXabswd8FN4gEoOl2ENefVuFN+trotyeqvIxaa630rxZ
4JPH6A0i7eRN/v0sa8lje5vb9GOjemha7pJZvAHa1Qy43CNvFRBHOp2I2VV3u7Vv
uUfH5GHE7Zep03v5bDfsMru1pqHEH7gfAY5OvX3D1qEUk91BVJ2a0tDCJsEP8I6F
fLcPjq4k5ccR61ZA9PSqM6G7xoPGVup6F0AA6gV/k/FJPyF5CG/T1Hkxsx/MsY/Z
s4V42WzwB48E3o0ewSGwpE4lkx/MlWMleJqruYfMpOgRkVaxG0UjC+rQoXoGU3wj
CGoaW9QHXoGEftsLBT4Hwd7OewXaSyAG3+GSr6IY7PcLY3nlCHz2uJmWmzTlD/Fv
IyFSqocPo28AA12GghvkvuuPLJ3HBBFr3GF36Z/+9stu9jP14bJWH8ZP4+7Uc6K+
Yl8MZkasc04NmHLrtZFmLT1OxIWNos2bxnsMMVwLRie2z4d0eSVAX8M4AVQX2s5C
NUZeSeBN2NvMg1PT7FLIH5nFVjntWPoMFTN7dPEp8nTThBdbOn/GLKKkvRq4a4I+
6buAe9gJeBDPqTmJa4T6/+1nMKmLEqokFFMQrBxZmyuawcrfp4ZIxBbSooLggcZZ
b194vdw8oMYRYoITjsNB8OqYn1pYsHefAezt9shmLUQtrRj8rSKRI71q+F/YCBoY
LdpQKu02RAKud0gpqr2eqgBYJWhV101gUvsk1r6RfMYjfci6jQNQa3pQsSn+LIGs
+MFLDJRRTm3axq/WPvk3IS86LQXbarLj185B6bUrYkF5pLwUkEv78DPVmhQxh4zg
omKfMf/MossTrZ2IjiOF8qoi5qzsY9K6yVKWCrj4duBZqhME+P49iOFBBJxSdpDF
bBI0s3nKNsq6z4NPReft2pI4LfK58WQ3Pcqm22S0QZM0g2eVA81HQ6etxJN+1Th4
fn5CSGstrCp9ALzlLGMDRyW8p851+/g2pnT+dFNQ+dE6bsNYlnKWJTSmOE3ymOGu
6713XhRK/ZK4yCvL8efUWJwTEYSPrmRyV+3SroiUaXPOEpllmJikH29PxZzrZ5KR
AsD5ENJyrFvd2uTPTDV+MxGFnyBv17IB6gmVp1snWE2wjnqsXrFGAdlFmcuOb4WG
VAtITGStvaAzn9zt2XPt3FffPFbsXK0qO0ue9OZbh3ngiign9cyOdNfeLDykJ/Gs
ja4kpd2neuPc3qamd6wPQe71raIMYFVaO8zWchwb1V/rHkt6boqzffdZ5kQ+se1h
r/RGT8pGU6z8pn0Du8xvK8uRyFJVKQ3+0GEGNDUjEKIXNzsc0gC0gMKSqo2Tc5Dl
n0ycb6ZW48NhfNesOP6hyzbP5jebgX06zJkGHqXuVx8tHPtrla2YJGgvOEaYmVBK
8D4OVSIKjXAP87Kp+JZtDi+oh6lwDwwElZdMAtVwTAkl16OROajiICI999REoEQ+
Mjbdp1MR/4lVZEbK3omlJD0d7yXE7a5EktWlkFiIAKJu5ZfU4X1kpsoaoP0OWruD
8eytBWsSmY+r/fpYUGJJ5Kka0E4/SPox5SDNXuVFzjQMFIS45B37nJVuvNrmHt4u
kV9sYZpCYxSVkEpo477mcAp7iAF7ckTo6hsPsrYX/Dw4T+2BGaftNENzvRzSluCo
iMYXuZsOh8jHxFnLpmMyShc48hkZmXCXqmUzYkP5bRqo3hWP4a0SKLINMLasEKZX
Hf33uO+4Kfq9qBHOgBvG7KbJDIYpVybCeEJic6aj8av4jhTSANPl66MkxG6+bePq
h10u0XHS1tgd3pIrK1Qo6zAAI4Nwj97YgfXtY/4NpvqbQTTqnYROQ1pU48XGd2Jw
5llGJYndue0iFUH3hTnUTBd/OFOysXiC3fMqoudIPOhDQoxWkio/zgVvZiflc8+r
wHi5xw91DB1EbejnuZyJZrVdXJ5kwoDDQ0zpKepgddenvoKU2nCpcK5gQKoGcCHI
C9sd6hYppnPbPuAmQMxc2ZHpUnkb6bAs00jYd3zs81/FLf4vhXWxV1f4Htw4n9mq
+eHejlhnztQ87xniaJ8iWcmZv7HO1GJ1ciYu8FAFbckQ19b2Dra0ybknSp/o+DUg
eEd7H58vEt3e0+k7R8NW11OSLCx1C/7sKDh4zhxrdaKw/x6H9WXcELAV0Q89xG3q
KaEb1CFxXYAfOwHUDq8IsyTZkqdwvJsfkuTxUjiYafmSa/LrISuy6DfKKO8nto2Z
FpehUKn7dkf/ktLtA26MpelCZ67+HG1WD/yewYLtA9P0IlLiL/7MMpY8VxedyN1m
gsxJwor08rL1YYpzGzuLidqL5T//u0HAu1MoGdjBxGw/oa+z1cNlmpu9DhOLLVx1
zYVXrgO2C7rcYa+QJXXmqxztBjeXSiY/vrOimTkbcvA6m8/B/aHQpALLJGTcz+Lj
sBtwJlggLk6RYrisNamORVgfTJIXj6MYuMrYGBpVO3bmfmIEqGsij+nn618Y/ZSF
tpW7GbOvU28XLMKvBo0pm5E+ya/O7GJGVG8vu0t+fDaMD+Ze+nuA7o4UVKACwyFE
tGexZEz7EaID0wsJUaNEnJVqs9+vPccqIDzyztg6cwVgLx2VIsMi/Pbw6ABlB2yy
hLBHriWncnCaIld6TFy3TxJgl0y8xmWYB5t8F4cCkVCMwO6crmHwPv7M6oenLa2W
YUlWbm581WExI7LnR5+M9zZo5bG9ldacY6oFNcuLjygp2FAfJiP2uiqnxl0X/NWR
v856RHbE0m7FU3jXSO916b8XILCr388xtSuf/gLe5AVEMY+z+HHkv8IvpicfZ57Y
gOwY10HUaqrSiEn/Ua9H2Nq40hiNThJ+Eqfxa45/6aJKJh4OHP52hrq7uNCupqdF
DnKLwJmgmbcholH2WdRVa9BHy+RosU8r5vfid1DAiG5hlYEPo6oWscvXGOd8NciR
uWGjbQacqqYx5eZz2JctbaTquT7SR6wX2XheuYyeQ32/yEeDjsC92DeLalMLs/nj
4x0FlcEWTQrl4oOhda1q13/EqpY9tMY7YxyUJqmMuoR/wv6JOMxCjdVkMPpFPJLG
U42ljX4CBrAqrjASxfpx6L7SyvJc60Kl49jBK8xpVSq//LyyK9gKCFm+tw6GlUvo
hShfzsGKz38Mu/YgZDfr8NZTwcFPKhWNdup5493X5eCPMGMrHrsmLFhvNuxq5fAW
qD7wp8utO7cCkKJu49u4igcoU7U8LURduH7ORKFNX/78tKIYAIa5FyCPrzEFR7Je
5ORVPK8PeBSdWYRZ1MlAv7FnHTQAAzFXfO6nxRbElw6llQrTNrp4D7gtxcPlY0nj
90q3zW5c+3CRD348lHzdz2+Fzm4OU+fJzePpgF0x9ZWP7svThCtf7x/b/uWhLQ6M
CI95EyRc+Ny0Ws8aHuCzzgg6HMdFK+PhKq1kicsaYxmYxbT5Y2fJKbOjJzCNMXfG
eD8WfnwKLvuZGMNXkQN6UVzfZXhaBxRgpfgDPSZjjK9/hkmMJ/nrhpTVZkRB2mL1
M6X5AuBvf4bMUNXVd+zK/I+cVbuRBD7mcQuRxpgFBl+tpds+Z6nLN8F4+NLaBxwF
n2ysgTg3ACnDMP9Cvwp1EIN2QtEYjre+1h05NG8OjVU78Hb4GU54/yrq7YdfPF9y
Tl8mcpN/STnayg/io7arAkfMbBVoEdqCtuLQLO+tKvwzKajiQkcebDQ7L4ykmRB5
nv+VYDzRHmGxaVs/ARUbPGDAoANT9IdUXsY09gc2+U9U4TXWs9+cSm9TeQsjwxKd
RnN8jw0LsbRtpzF0cx6yLoqwHIfvG+E7OXr2eTsj5ksif83slipTqCF3WaTttQqZ
wzafxWe4U7nxGtRS7k22lxXU4HDL/jAoNYMv1ym6/153ydnKmANYkgOqq0N5R1dq
6NEvyOxKCCHQboiarLXzsH02H6oT2lL9mCbZkPDo58c97Fq1iMkRgXTRf1jOeOR6
cgkxMyRYRhaqp6xW0FJgPKsUo5uvpaXRp8dcHWMkl5jZYiubBmanx8MmeBilKzr+
L+/0rD5LDbxAP5F3WzackAj+c8rOShyif6ON7Vw4XYXRMaD8Y6BQFzxn9YMzt6qk
IzPbG71J3xAjjrFR3yocGmBP829xQMop+i1ZpT+xl66TyOfZpcmmmJPMBEBF3JsW
lmi/OAkGL81+xlO6uClgm8i9ZKu4TU7U59ztiMOZsP3d2HkwUkjAb5BbiQJtMrQK
beQM/qVqgxaoD9TDCjCPnTyGHfqq9aKyW7s+unQyYtv7qpclxTZOlTArOwUkIfkm
2dvddLhXNz2w5zdON82YP0Zed5KT1erGgrwsoIniF7Kr7Rz2VyyC1e0NAkoDjJS9
i39MPQKT+LOWIpHXL+C4+265+cWcDE+RAfjpr7R+wovDKGXDmF4drbdUcoeGJ5nK
4DMymCnDw1Werpi3E3jbEBl9ffnuArJXLjxXPzJ/9RDpUMOlM6x+3MB+nZvq9mS0
5JSDG9A69ElB43iUA4KjVkDpZfcxHN0SlppMbZ1C3mrX5usMhILQOzwR7kAg8V+O
gTNsZsiWHqHeSkmoI8E9RvotKoRFUNVGjQ+uDg1WisSPMMPT9bATJeFOgLlxPkMV
hYlWrOtfnJ3tz7/GY7djy9gjnqfNH/b4ZeLe1pJwAGPuMEU6/DjWgCEq/VC3YvAL
fue2qf4plT4WnzZx67+L4+CzjthPE8CJYUNfXqdJaVZJ+C6SaRnYh0lWAmWIkrbU
w2PRC6QctUPZadBlbUpggXTDyY7surEOltBTjZa8SeqC13vqZUHaO45la7JkVlmO
4oh5KBa5ykI3961giNj90pSDb0WYBtE6GOppI7mlmC6FYAL08sE7kt+MoEpJA6L/
ZyseBAfKJYW+QAVQ9OrD8KGY7hBVRWF4R1JssL2mkaQ31ZErcxYU78nZazBd/eW7
iCX34JXFLvauUKfiApefRV8f715e0+8J3Uswl88kQaIS7Ecs8kwXbmrn3XAYNb2C
UchZAdAK7eUwAzfIc6CMplNJ5+NX3fpkRFn0iBh2b40n1kSsvTAFcJJnrMgHxhxL
Ne6lTODEh6baZOPL204UK01KCb2DsDd4uivZXyvSBpzyxdINYuqEy8omgifmpaHb
Uk6VQ544JqFWe4ysOqdw6iL+aOCb0ZJrJ17H16WpZlWBrmeRFbJiUU1901KX+iwd
TXguOLJFkSNzZle+IAy0RNRbYUcUD8cOYu9P45/EwjxDoHYVgdZdswQH+qUQNjyR
c1c7waTY21uHVwqrh6wvIuk54Vq+Age42P3KIOI8GCR42WZHDwKZSlmJY/FQkVxe
KsBRSj6YFs5RpZkKhJa1MvuAhX0Xpsg4Ok+15WZIkiJnQ/9ous1LMEGsrM/YvY5F
3B+GngliieJFSIixSPbxNr+kA7v58ZNOg3kOcPcR5UZo2gLRqS7rfZSH2CdWVsuP
B6gGuDzkVSqlUvjcq4NNzMrQh8Z6zhX2HkjFNmUKVNr7mZEnsr6sO8pifUPZtTjb
r1FThbUSc8VZPZtZJz/KwVtn1J41AvFDCXSBFxSBYh8qxxM2YdCpBNZ9dJs1Zkf/
CINjLoceEsHWdsYLWZGwRQXCcMwL76GRs9axgzTn61X/kdKTt0qxdRfw22GH8LGR
kFjJJ0h/JYQP25GXBpOaJw4XPXLsNTAn2uiAKg+ntD01HSq4y0Zjvkgh9w5d9bef
tnhvpWa8p0g34/s9mqwiTRCnwIJf/f3fg70p52pvGv+652/8bOIIJtvltJH85ZpZ
Wl9EnatrtFA3UdAztBuf3Zu2LLfi12BE9EIOa0NDlQTaxff/m+im+WA/2Ju251rs
mkQQS1BqJUubbCIu24CbcV8xK/n+NAEgyUHARiVEtljRglYaklKpdRgZbe73lS7n
8IIlmGrzT3TzanJ18YolAGffM4PUS6NH//3jdZs1+M52a51dUxq0daFw6yPcwQaB
YxiuLia/EhJXzJHO3mehBrGvJBd7AMoIBttWkYd3WvbpkBm3OW326+k8aOJ4gNLZ
JRnm901vfDIwtVLKcxRzs5y7WnnDtjSjN9IFNMZ3Bn3zNVLD88tZ8Cr2Q+j1Co/P
5guaqb0KBxB1TdJRCTm08sstM4WYYOL1+SQAZDkcnXjLjTuC0FUl7MQioT8J7INp
jIlNqnzrZpGaxu9pwwNcn/40T9RPSGCO97Q0bcYQ748YpjoqcFCsvirCVutN7qQ3
2p8Qsh9bvB6MLDT+mXFwEuiR4DMD2G6AD4k/3dZsOnEHt7vfuDCdaHsI4Rgre6TL
rxkoaIUjmT2CyK/HdG3tSGAzKbO1p/mYQ5Y8vS/Uy2wv8ELywsFmsxqIDlXgPdrq
ULijrpYA76c9lY0aBI9p+AghkkGJtsNRg8xP5oIo/4pOjl43mPDvFDJ8CWGbOJGp
BDlNb5PAbw+Bkn2A6IaMtF7JL94RV7jaFYP66Ro/OvHaGYfyn3v/3QJboHjjlU6f
deCS/jFMAX/PZGXQwL/GZJqAUfvOJDwRP7iaP+SX8qXJgclWJttIvCxknGQUdvqs
0aQUyrOtchIcKD7srGcOJlQjP71VJ9IhTl86OJS/DW34JthRCV8c/RonKHjJC3aw
XKIQYm3VClLxG5mylcGwmaK5yZNoD715fu0S09nnnouV+opuS+1hAvowQ7iIaODG
2CV3W+FtzrSjdWhrWIEzqnsLs3c2H6XR5tBuEBkX11L55ZpZ9nlHxCk69ZoIbfbU
EusYUOm2ezrvs/fjWbzG7SAP2/6w0E9pnnvmRkjqG2wRWPo/4P7oztP5HZzNTK8I
Z8wVtUNQI+KalJ4G5o9VtdjGl8LgwKutIVp5x78ytViXvUYT1ePu/FNzWVLwQZoF
QAG28h5fzNTZlOvlrU9lSOq5lWxz6bIB1LEHH40/uXq6lXyPG7dNe8JRnYBSlUj1
JXOJL3vt9NvvZB4UlMQAoZCvH6wDBpKLQ5mDpx/zoErprFvQ2brHYI3sJJa4eaP1
IT9I1Ecx5t2OBnnbexFiKB+8+d9wFTf9s/5Gn5DeoTgz6k3f1fVdTUSWy147lCnm
Dso67wcj/cWIbem+y+j8WRNthnaRHG/+1NWlchKxgGlYsp6Ir+bZGVS8QyjQhRg+
9CVvVNvwYwOcxGrj8jARfg/Nq3FwcqKM4dv3dd7TGu/lQUpenTN+6bsrlXsX5F5e
CbOJiKvLci3JyPvjq8EkJ5KKAK+dJJoRhA0n3nUPadKbCx+93126fDqhQaeRG75d
uIZ6cMbjp7nx9GkS9IKqo1EqBDOyt7SKPvm37ASDUp3U50MfPPdYmbWQIX9bCh8r
2MmORmDLaiunSIXQit/zgUPel7lNEmRZQTXaDpQLUcat5ud/QvxTqsX38n9ar/WH
HcWNH2WNxjXtByFbAKZ1HvwfLQmgG8Fw6SdQxhmGbSdT/ZEZ1gvEZmtDCFFnmoeQ
Rp8JTcpnWt+Fhmorfe0Tk0yaQt6D0T+zJ/qH2YYxMSYo6G8SXBwoK5PZIx2Z4YbH
W67rJqwWOFuJqroKvIIyfI75hQFUg908vc+pi1MtZqvVdesyU6ZqrRXHHFmJIFbS
OYUkPeI6XisBKam+iEId6HXgSr8y3nIyh4vCHM+ZBYXVnvyJ1phUDtHVxKi3tY1e
VqOn+R4LZzHrqAQL5dZ7Mb67p3HBaf1Vl2C5flCoD3UJVs+MZadg1u3ZmMcuwxM1
B3pNci/GnnHdt1F9TMZxaflc4m3fJcoHq5IkUxSbKpUxBTORw7N0WzKGMaMFGWED
vYgBgkjFg/58rzLcjerspGGvsc1qByD38LM86KsO0m+ACVIeZkUYpgmf9MiMa8W0
oWCXg2tYkwnFBVwxsjtNzp0Tcf2KZjUaebb5nubOuTwUBq+28jli5SJhTSfrBdkY
YJA2VY3Zlm20Ei+1WNbY/77wjMQRb3hm9LGRm5oTYSlVYd3VuyOR7ax8XHgDa7uW
WRm9BOOWvrW2UcMLhI4xGI4InDCNGHg6bhHRiPndcVhCkoZfVdVkWiu9UZSuSOLX
sd9pI/aInGwE8WgDc1aV0PHsM3Kywa3TM1znH4WSNcedu903x0tAIj7j/xaSCXiX
/FLTScPhE5FDImhVbC6bxnNpWOGL5HfQh4CgjxAEyQMSiRdQofibyaNcisRX40ET
gG5FcfNkzec16f9j2ieTSmoQ2fudazwQpdGwPokdm28=
`pragma protect end_protected
