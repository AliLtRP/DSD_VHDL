// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ly3rKpCT7wEJCqCo2gvqEZbj955GH1F6YCMBewdJQFwuXj2bysnzDKeHfLxCXlV9
PU6oqhPUhUjO/fsFeHV7PEckYwxk/hB/oKXkWFuoGmO4dtlZVtMX0apWycdoimGg
z6A/diRJUFV6rXS4IciHYGEuFQ1mccB38/Pi36LIjTo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5344)
asyDBdrCTxoW9jPJzahRuSD9h0oz4vfTh3WtaqyRLenUozTTkx+2SRipz+wrub0S
Uqv6dopur28Q0qqAKPIu39gz4twY67O+plL8YkwROIC0nMgiKkbE4JDLDkn8h6kl
4+NVs5QbmB7KTP6JVeNepXsHT2S3AEM+PeFxLfEC5415HnL7K6sRoHTkuul5D72o
R1zsJ70CgvlSKM+tCoZHrmQnJlb3xmIh+mlcLYKeJDDveJcbU7K9qzWTn866k9zd
I9u238hZ9dwyOlBGks439BOEZDNlzB7k/qrC0LDkgXToBnmk9ACqSoQD/QjFPm4N
7wlsZLe2MJgOxpDslfjP2vlqlnic/wL1z/X0oaFX4vKOT2tQEsbFJ1UjNyi3A+9q
gxe49fcUXGrZOFtTk5+TjsCQf6Mr/joVs9W25L5rH8ASM5R5dtgqiTeXtVjnako6
V67Qn0PC9leEu4JtojyJSiqBJR09+8M4f9OGQRZED22KXXer7018bIFl3QHxJHec
9kK2qZW5vHZI0vB3YVg8YFfnP0jvnQ7o4bmcRXV9HSlKxEBDsNfCw6WNqOSBS4sX
8wrjHBX1BUyVF/z/2mG2X54GqN3TC74KPRWUdv7SSQzn5ZlYcNunxtkpy+nvzy3n
ubrsmXF+pnCkIk9/xkzRtViM7mLObl56u9aO2GPCGBQxZAYBH8uvatHKIBFB/lbK
16QapsdzpXlWv5AAaNm51Wfn9z0qPRBO0aMaWxpI7MtQgD03RiuXPo9hmEcdg7qe
+z7Kk+ayRpdxbUKs45vBZQdM7QHRdlvYGHKtIXPZiXeOuGts0Ow346pbv3QWzi+l
9qRWsfSSPRQeGXNelt0M8kksaxzu9EtK630kUlE5T4gJxhNxltqgOw8YIiY2viR3
UPMPKlWNPAClVC80rtzskUVWiGWpqOyuLBWauoLfn7ofGvxrUzdWSacHEEBbTVww
P81mxFAr8Pz261twPhrHQe10l8vu0XaTcttGEGfWtkxtPoL804UOJTlugAUKvPHp
XAkq3bJVgn0QpKM5hgA3J59+ZUpjNz/49xgopHv0/g4+AukTBMKs73CCm/vyiXvX
tEZ3Jw2S453r3xT8CWZoJdu+M8ZzFmjqoaJQW7nNhwyvO99KnPUQ1hHedlxhk1PX
Keqv9tx9ZZXh+ZKj3jsqSQwMnPv29l7kIy2QF+s03sJ0EQN+8LHLzldI24HhX4RX
H1qJQsCh38L79L+8Mm+AE1NsFxEW3De+KYHeOuRldjeqSepnRbGTlvxRujB1F6ak
jbWFHez6W/8kH7ci0pCbKyw8KDhWpiLoKunXyUtIF0Q24YJGtk6xtcu3b3GNL6er
3YH+ksKBmkIoTQIq/U5YzkN1IA+zFDnepKnB+MT9H2UbBdytAKOmlpwVsFDShd92
9TSzhswgmiVtkQGxLErYFtPs8BIpf8EkGSr7lpPfVo1/nvgx8Wl6yYPWosARzwIK
APG5cJK57syaihIM3QLPuHF2TEdbiqiQ9NDWd2pRnL2xn2uYWubW/Bb170vw0Wtk
RSp1sUx9EkGWEGsJueJQHf0K3fMBKzDLHwi0sul1v8hr8jqa87jChwTtM+t5Z/b1
CZgWMUmwhf6iItF7FQFuq7F0GXVDBxFmLN72BrtjqiBeY8VLYyWX4JDK9lKikcEV
Wn/OKhqQ31pKqCqyYpP1zwdQDIqLEJA8+B/OB1TT7iShKFqtn7n6YSzoEG3E4K2L
eOYBWfcr1R5CxcnCqQp8215PxnXZvSl2WbBkE/QpIBSk+E0BjMJFE4W1DwuZsIlX
suWikT1SK52hIkPmt82LRc6d7oXuzp0VIo7FYALAGxZBgSTvod/r/0bSE6fDTnrT
310f7AT9ahmfcoA8SCp9e/d+AQmBgOmBvAmhAmpI4Fo9QyWy6XUvY9XjnPc5yC2E
UqpD9+Pw2qwKX8jsZ/2t0ksH8HNO2ZR2Nf/7QBkb1vNX12K0Qo8AMWAhkpkYaD5c
4ODTH8M4vsUkeFUre6X0nbyuW1FUxLB1tnUSgE6YNiOO6HebZIQYtzBXJGJLPeDN
zPqAZpg8wWz/sGRl8ogWrh5UbsLhM+n91PK+shoZ3nsoJR+ENLnUB9kZIzyFA7NF
RYltuJNDuWVgefSP2eJU5oU36q3vUfnnRr3A7cREWJFp5iXH08MAFXXCpqV3znF4
9oS9VRs/pNSMIppIHhvRYza6VNaVLzC9NEhY9lhZboojEsdhkNd3th2ns8V2Kv38
VG3V/7Srw3X0hbwigy25rsU8vVuAnkLQrqA1mY2YBGyNjSFAGBr4H0JiEm6Q0IHv
DLYG+KNFZqWF2DulBCD+29lqj2LjTCB5/g3yaMzbwpqCpK9Kqe6gsuhvf1QkG1oH
RZM5mNENAHEdzBF6UNgpHud5U8WWtcIC5yDRKIts/0S7eDFiyQkYUuULxZFJoBxM
eXOiwA+TsYFBMmuohre2PYtgxw9Jr+V4Pb5WvV+bLeGR2AJTxUri4unTseiZwg+2
PPZd7260E5W57WbSOClzIacz80BEHMjoalPd9AxbBAvooZdn8o4JWJ3Yw6asn31V
mBmRkoShgtxtSsdDnGTC6DZ0TJUDvW3P/pTqEulVsrdXe5HPfLwSKpj7VXa01SHs
AFA3QaQZwr8BZsyemv4IEu7TYYSw6rqRYMy8Ghjx5wuLMolO1Cr17X9ZespYbnsO
MD48w0GIJlZ08u78X97KQRbvVT5HEqwI1OZN4jmMYS5AVlnA1sGAmuz8M6Hy4gYY
ZcXX82HupWJr9J/oifNkii0LgzT/+yC8tXGIOLeGEX5SkTpfzg5gVZWsB5BAJ9ae
x1navjtLiyH5mixFcYSXt14RzPHHg0nET5Izv3a73t0p2FD4+gUQWYg0+aXGWB2N
CgeMOqcXQJ3IihwRsl7hksF/5gfOlpZYOmYEYWp6AJf740BUM4NK4CezRLdbyGEW
UUKHZrgkut+QIX+5Y2H5GjJxke+LflX0dcRdGUdxgxhs8J6jnr8nZhRqv1t1X+yX
v9f0UJrvrDyKPEZhqrJ1YvzdSCyHjhhEyjqAOqGtA5Fq2uOt/V6Gu8gtuBAwV9OG
JSlMHpHVf7MfP74wCYk5SSkx5raba5gzkoYEoQjMAYPKzxhMvrFHhBPybgMsreU6
meFWAaDrDDseQC4StSqL36kZL1QZm1o5uPOh/06enhojPu8xrTfPLUnZ5RTAcW+1
GDyZHqDvaoB+lymGAagTpZ29eIYO2kPawd69WL19j/QK4FVT8t6xxHGbyyFdd3Ih
OqcNekqbqt8R01nwUFarkiCyASsdGMqYUvjw3hUfqFjQx4JVeh154Py7XHvmKq57
v/QLk0hvCN3d6NaIRKiANnxR3E5dxWSJ8jBfcQHfT7DFNXwMGwSSpmnp6yGf4eiO
PG9U6t0gy4NT/cL0Cw2ldmiX93ItYgQm5RgEUeg/7RoDZwMqWvM5vUnGBR1vll7k
rIhb2vbaklj/PrG1F9mSAB9dpWcohaOn5vZhq3xtrav/UhJuZdPaY4bwYZbwNvHk
X2qQ0xprZYoqroFHSfdlNh3NiUkYti8WD7RNTz1dMTWGPWClXXbdQxAabDlohyWO
vCZoe7LHVFpC47U2rY4xZZvVngkHB6ApTPZ2TDeKMzXTc9MC/ELU1Xqr8MonsBom
JnCI2YYF9FxdgfZLx6uiWPVo3bvKYCu06YstRY5vNltfBa3a7Emi28n6NiJxA0XK
BYhrLmQhe7+/17Owpu9MGkSPZsHhSe4Z8T1xRADcYueC59NkyCfPM5pHpv+HKAL3
HYPEi7xbbaNWcVpa458CVovVvOEW4WakGNjd0uT2TWnn/WnXtteapv4uVld52h6/
3Xv/+/iGTbpnI+0it8C+Xir2ESIdV6NRGmV+2UXoO9xhS+nzq1wpZ9eSjdVCdZ0l
igo/sOr7lMWRCrpMcSUX+JW+pbEIG8QQJQviVQXXov2IpTUzx8IwFBUrrxHN5UhA
N9uVAgYYcZVBOwIJkLYTVOP6UP+/yaPWZJmKs3UGMI5enNEBV9icsoPXSTwIpqMg
gMx1bt9BSK4+buRbIkvj9cwxpOAZqaVVAO3tprGp2AEI7bOLW/9hQF0Hwqjq8gLU
qCtwSiR4OYjG2vxV9KtVKIw5GiW1UPQH6vDJNl80R90OWXtUCCWRv9DDcCq3NY+m
dTGTD3WClB52nFT7tcx+BrEr2GaOCyGAo+J7EYOb+spuXJFYd25rlBmwXl9C9D+2
kRNa/1H27S4pMRvcNAbd/jsdTGX1fcs+JIEq8ziwZ1g2fd8f3r+UjufMQHln6I1x
wvFk6Lkk9lMu16SaTw//OYRwPDxAp7LKv2zJiu4UO4zyHfotYvR6aVImFDV1ulev
n8OXuGIOtcrGAvSqxZfL1F9hiDd5g5xFAbB996rXaBIQ7YZPFjGfW4FruinHvJEo
JR840p6w5GMyKfUq5ymKbbytyrtnxFKlzw+OYOb4eZ/puZQtawgUltgyWRgk+igY
ezbb/F+3ajVznLKQ6/IEDRGUBuJPhpkdVOY+WNsa++ee5n/Vmr8qcFIFdjhZq4S5
Ewd57xncmNiiQv09oQdAcCgomYzRLpr8cuJVlD1xaq0/1Sjoud7p3opQEP23/z57
itnPDt7fUli7BoV7sSTjPiBWzgJP3yY96PDTHRS9Ss68e/ljQZqEyhlWZMlQzBB7
K2I/4KGBiWTe5hct/l/iiOXA9IIZoA4EDI9HtRovuPwWdXHNWHo0VJOXPChd0RfA
nW6W1zC67CzeUZNlaFhEb0+Xvup51Osgqq6wMpBxXw59D8j48hZ+N1dJnwyJw1xc
TlO4sVWFtz7fY/irf+OAva7VCYmsyXybhw2Ps+WEZooelr/w68sjU8gJIpPRJ2Sk
Vf9Ly6kHVDvCmmihWMrdgHXOYDzdtMU9DozxL1pylEh/9dBKW5c1KzeY7dCWlbkn
2PNxQvmKHf9oLuEKeJlDadGtzEOBDwjQ7BVbNjzX9qb7aCj+hbaCdRCEVGfo5nDj
edRjOzqzp44rXiSb/qdEplAPCHsqdH4uGZVHKsljlyYswALAst5hvrtTB19ea9+o
aPUgBhkzbntgbeh4zfOKBGOsrNYFTZ4h449ykJLg0NUEcFsT09Y/9Xd1mxurMj2f
vGq6CjeK//Nm8P1rTA6k/gfPqkWWCypyT+Mj0rPrmWQZ1PG/uYNMgURQV8IsKpSE
+NgBliAxX2bDwiQGL0wNG/yt3BQ1VrDtt5s5r6qhnHz3lqbw2yqlPhLqNxU73Xg0
4SBlLdJeIaN4ijXRdi0fLZNVYI2XPJInsUcSq5rY1SrnNFaAFqBLHg5yhGQ3JhiE
hatrTt6mB1YxvNHwxx6bEd6JrTpybrB9VYbAahj56BQRVGo8IxU/FlfvsgbSJnFk
P8rcboN1cRdJmYC4yJATRwcKR1RQLLrgQgzle6Iom4M1FZSQHUeRN1JHoh1YHySj
jiwFklO/m5CvHNBQ83dBAmGvR7C/pcUwSvxaGg7mHeWKZyGXYNynOTiedjKt8MnP
zrNjNb7En1KVWO1qqR8qteo8ITWUHqt62Y47avzoRzhG3x8X6AuMmQKbSMjjAmd2
czzeaRINZBDOUUem3FbdnPIAYmUAS9J/x5OtjrNgRwVjmkk2IyoZVn0vITpmvBVc
kYyohZ+1qS+MtJUXeZOhjlENGvwdrgHVplf74e8EOuxF7AfdhV+10JrIcJMhWn1g
lJbqJr0aKHdIDbnDkgpJ7RvbbD2ghhkmAheeaakOanlCsd5T1VWcNDwS7aKvVh/y
88T9SNfo838CQz1g9gH8se8SkKfNyetIj9xcr53hi58iq0z/JrYPJzKrZjsboikE
5hDkpgsYlEUHJZqh65Ac2xywmYtEdJlTyUOYp8CPBxQ4z6xcO3vfAJN0eFfP0nW0
VGkwZFrlhGXL4fDGzn/zLnqGgFYt3a7wPfXjoY+FpDkN+DB1ds1AbtheBWaJyhQv
r2tuhH8elPlD7xV9HI4Nw3FKlgnzoaFvuv6dk4MNVHCt4J9kliUYHM/6tQj6v/5J
NvE/j+PJpntzMesP+dopgwkKgWkrOmvEgvizxJzuJBwUuA4t7A5ViaTvk3rGDLcQ
R/NJiJFSi6n2HUOLD3kyDkxvnf9qj6SwEewcFVnkzseerBmS5IPBU0AHx5CJjpn1
i2LDcqNqfqHWSty7gMfzXNTb3XDpr3zmiYz6Y0A4CVd3Y5YAxmo7zdR1T2nPVn9O
yy/eUptcnagL/1h0MSgfQWPxlSgpON2iNTcNiLivCEyIXweHbpv/0vCAEShIQn0o
WAxd7/J0nVDNEWk6qCaMJOVx/r/hjbKDeGtLAaForjseuYhhPzxg2QUQ5sgXfuJs
viaqfKJqo8z3KERTrvj/0L6YNPNJiqoajHoKdH+Khx1zLvagK4abXoM7ewsSSoNT
P5fBPRSpXu2Ou9NpejcupIUjeck1+Z3kVSbUocjVOcuBPAKAMTC3C5Oced0li7gr
fTOgdhvImKo7KT3toDA+H9CzQatGHCXWPJJbRM0JRe2NVcwTPSa0kzM6obxYI5tf
Lvohzyf6ntLY6axAjPPwMDf25jmIkM5rbpA8zTjRhOuG1080zcfzDrMB9usoEKWZ
9SvtmOgNKmuyVvqdxFa8n5zy/gozwS8/IN+FPAyYWRXJGlCmZugcP3N3j9iJDW/k
ZB3wsVUUZUBRGYFL0o9Wv6ofLOqG7Zzj754DTXYSx7dLJSMqXxemfw7EkcxQ+NY3
tD7fOguhyUusE9yto9buHiOKJXyW/nVIoPgNmigSEctxX3EQ8MxN0wSfBUVzWWgw
vaR5UCmC3xHzYsV0tkThL6sRAH6a1wRFtMpzk91wkoajuTx8WJEQGqwDZTooS3yk
g4QvgenXPBPvnozvojNaxSQLK2suPN4hCnzRBpKhBpRBldUC6XJG/slynBNRj/O8
I7m0OXQ+3q/eAFdhRjV6anYTJvjDwJtU31nyq764PdEHWL7LpUvIbfxUqaiwWoKI
/6jSUvJhGXrTQV+0xOFezBVZ/cr7Xe6VVfTastiHSP/9RDKCUFuP7Vex9SbEzJ/A
Hp+7K/DQJDVefS3cTNVxomYClseV/T0D6PHop5i7B3aw5hJ5FJTZHi1Tq/Y5B4jI
dDheM24f2V3CUXqKOZij6g==
`pragma protect end_protected
