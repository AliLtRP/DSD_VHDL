// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nAtBjQhkhv3SDEws3Ux5l0K3THsr8/0oW9RB7ccr68tgDEpKckGLpgJ/T0YNV1oX
9+ltE9MLU2h5g4tOrlRLSwrNfn2Q/c8rixWNtgE83Bdp6b+SDCDY5Nk8nacofEre
cs0tQyunpO56aA6enTYg+XVLdsFMFY2QMKLoKqU364Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17728)
+doBx7SLDEpT9W8n5tg2+flYA1STBl3CPU68BgRkkvp3LJtWWuvOqyAkpTJ22FQx
8Q+zhVR/cU8+sD7u0oCBpwBKj60fhyf4Gd93JBRNHcQFH9FnfEiHkVGCgMSsKkMJ
NlMkVeJrSqYWNQpXKfv3+PC5SCgonaIAi5NosMr4/IPzjZt+QbyO5Dt06pHMRTO/
J3TPXqnjFX9R44KgtlnrWTv+Y8gMaiBukMkpIXd+BG1Z75tnTkNVYtSg3EfFxYYm
iIDL68nHuOOvHCKI2lT3UO1YVchX7zQP54PuXIbznJHaxQtlfJaksahnleF2Iymm
WmyPyI3QOqM4ZWLkFvI0UsHtBmRUitigl5N/WySx6gPHDQkxhUID7ui3ochnclDj
NZqZlHe3Rhpvprj0jpIiPWyDytZpp3NHn0HXEdX93hBfjsVqtDkVISiR3DXUhiC9
PrLycEYRuhDluxdKRdfvRJ6RLX06I+ZqCqtT7rvw6/qVh7Rp9S0hhMOVvnp2XrhW
OaDLVyzq13acher9LKs8pQfny5Jnc987RrEx+RgMGwYY1nG/1MuWDIyrIu9IqX4A
qAqqSWCX7b30j343v8MiMn36RdVrQcLiIDwKN9HKELtppMUCGki/HFTFdEMmODy0
FR9L1AKgQREVCb4APb5scXwKHXtUUR9h3RJ84Xc8U2EuY4bRIUEh6wrtDMT2KRzP
fhbE2ZfQ6iNvFpdXCcqcpnT9/rd8/srVCB/HZowhogP8ZkY7oQ2o6wjFjMdLOO9T
+DhYpjJCGH/1yOAODZbfQhJvAWEx7qdLmiuBQnHsmUomd/7S0sHt2haYfuOw0ye9
v82ak0NeXOiyXBbEG0+oOmG0fuGhNyxQB1HFGtaaOGuNJIqqTbSQ5JVUitOYLt6P
SaamwcZaFD9S3P5sX4E+mm8sT4qxvxs7Lz0wMDOXlRhZ9xGCxaJz77yJcb0VPm74
u9/LSM5v6eeYkgnLYgjz4gfntWYZi4kFkEg0eOd15SKRBP0I9JZkI2RtGt/lf1Sw
al/GVnLu5XVPJpZwWR6oD0lMssXiu1SVkkcqlj+kEdgeC1uhQRXyqyfz28TMNkbx
8Cz5IXHKPcOEN9RnlOghpuphcO2Iqa4epwVkwBeSEHPTBf3uQjgYjyXDC7MB/Hjk
yfaqHZT9aZLioaWg7bAsTwDs2eKOO/tYdNARJoDLFnM8GWtxsG40sjG056raKBAO
fKnJnMD95E6l+KDaxehphYPVDUARGZNxFl3gzS9lOvksBGoMsJ/uNuaThSFMv3vu
8QO3dEZZlFyc2MrIQu3eX/27wDR80B0URnulcUDp9YA2WD6r0+RF5ZfAult1vKDI
5XoJzAXsGlo2mpEwJ7hRzeJoIknYnuaSEeA4APjlgaeHewbbWG3U9XPo7dy2DLTV
JxFJOwckaIVEaA0ZthfTFCqvYErHzQn9leHmnpXngYzxc3ns3m6Iahsq+RuR6rfL
OdU8R/kYu6GvE1YSsJyScHuXLQQfIoE3ukj4WPHrThjitu2z9TUIGDyj8uY3rbqh
Ur//mny8c2fW8aXt6IENbdqZPhOYx8E3eAFJ1J4pZmSdNloHqfbREi21UkIGCSSM
0EgVe/qeLZbsSd/7w4nXbFGTOmPkBRtyRdtl4OuD2qxM83J3J1M+mhOIBjpgt+qh
QjuIQ3DfQwW18OGCiMnjPUmtIQXxV/aZ/zdM/VrrIq7QMvvaOBEMZ+h6DCDB2EV/
qGi39KpzvX0iirj3QzEbeQKJYdAj24k+s6xrpbrmf7/XYv1DpfD7q830NbnZNXLu
ZOfy5uZXd3UElJ1qABFxej9gfLAeNFdJUFUZU4wXJ87NAIbASE/1CCygM8gtNPKM
h80w+Tx90TNGwL1yHv3VycjAKRfAoW5UtGcYFUgFcg396144eQ/nCfhRSnGIXqkM
KkG6db0ezbFpwE3Fuffr+UlPPhnAUiiydtqWbSqK9NOL8BwrBXv8MFa10c02XgjM
oyCZmmdPmmW8Q4CEdk9R/hi0QdLo/G5slUFE9+T1YMEB4BXLF3Jp2OQd3o3JOroS
gysXDZL5Yzqn01w2ptDl2UV0J9sexrPvzc9Tu9j9YE1gPilmvX7hPdRx/ny+KXbx
0lIcZmpfu8BkhCkIzFgMcLE7NIfRhJ+7uYN5Az3yBFhdKJL+x2VU7kI1BjtN0H/P
v7RklHPpSnXRbOCLnxtDoLPQ4GOjqhtS1+riYaNAgzg6aATX4MPipZS+Sy6IMwcA
+IB4BchFF4di6OxwLJzbqmL0bWeDMgTNM456Vn4yQWh0U3R9MxW+ln64wNs9yOuD
wZiUDjLcrn8tMGcAjNuuNjAw/kGnuE3lKqj/vjcT5uqilDvaKhXcgoJ+d08w2Z54
h9xVLSNxHaBsle+PNp8O3X7qsE46KlGI4f4m15IRZCURQuoUwYVYVwu4Bfpgf34i
t+Wp+UBdNm9txtM7zLU1jIKGw+v63uMhdBBK4cF4qkcKfjwAo3JLCy4KIOGLly9f
D306nWRfL2hPbqg84xdjaxoTEdL63T51yN4nmy4pW6hZGy5G00KdgfOOwvjBc1go
plX8+AXXMWt0FQaYyGqsQmt8L+2v+CpTyRfRLB9xD9WFPP39yrnViFiE8w+axwV9
iDXr8zsWPZ5th9GA+4vJkBJMhmeqPixGuISOYv7OQ7jyRyGR73iMp55vUmlkZNki
E9FM9XGBA3WvtDWpyhM8NBVUXbi23pScydLtG+r8KK7RDrOzzCAe1xGUHLGVT5Mx
+Pghdlu7XnwZE3PdeP1Rqdik5KDNXZbYo7H3q8a0lr8xT0r7Rxu5k7KmTx5R9Ahk
uecJxvZqA3fi1w6hvPmVlb5TfHX0RdYIGP9PNSsGE73Ydjahm6MxXR9scE/DZURW
NUyvXAAZrTP0ZiFdEjFzvO/2HT9t2kg6iyjBOrc/bDvNbV9e7ifdZeAaUpZ7y117
DH9lPGEEHx0spNEYZ/+St0VhqSt7bsOeO86YsP+JnyRCFTaF6pzDYg7/PomhjHwf
Cr336PvqJj0GvLaG8+d3cXwMRGO+Xy0h+VIjffcP/eAEmL9dckm7rf2wovOqqUw4
ssbpHMuKsguUMu7QRU5/cYvSsmHQamutiA2OcfAfLHs3MJwe0elQk3w/BjUOtGTz
aXBoq6O36sDdBYlk8yYJTwNRDLc9hmbgEpkIQTa8lh4BhGH7Ud/7qRHRVaqm5BiS
seiccVxWojcp3pK9S21AAzCy09HLcN6AKWfVWK9Rhh+tNwp6j+yLAHRRWG2nCaCZ
uYtnImLE25GaYw/KnzTgNV8A0W1DT5TmKRb687kCeNDR0jwN7uVQ2KCRDrf+o3dz
ankoVrwQYJM4JN1PCr1HycOf/ooicjCGSv8MhasmYSZfqjH8kRkWy6WogJm2clhH
o6I2tAWiuVL/8eqlA34aC4XvPov7qZlvweePVlQRjn2xVcnnTLgCOwofsxP6BWbe
9yRtnS0whwf/y/MvJC7/+I9M/k9Zha/ks2fMAFrnebxWjNUc4q6vuG5Y6G8JKVai
z04ruU5VsSlwVWiir0VBSE9iFe4OT0K0jc8m5+/K8chmmOyVvhtrv6MrLjyKmiGY
dIZmJeOmCY6F5Lm7kcnHSa1yE26SFH0c3t/jzKL4md1x48XjhH7T+34x+fIgOpk1
Y1R3A43Qh2e8yNdr+2bftFEl0IxPvHXgEwG9EHX0P+JeZPF8mrGFbETbBbxgP1Fc
Tp9KBk2AL2H6lOBE5ur6z/4Qlo3y+jniNJGgR9Q4zr8ronpazHWYMH5NfpWb0qXm
kAIdiBHiitvritfYSGyksUmn+9VcjWlfKKBMgWV/xPU+iKCqShQKVvxdVJAMQYGP
ipP4xO7tncjZTpC+C9Uv9dSpzccVA/I1Vq18m0xANrZPx7F/Mw0cOyBERtU/xf4N
7e/M8fQy14QlCsRyIGacqRg8uw2oBBQd/54AQpKHglxJbSVERondH/7v71Fr7rRC
BuiGr/xGYqzNy+su3bD8Ypyudrd2WXDHyNezZRNd+2Z7mEJFmVtlLRFWT8mMYe7X
gl5Y3S1pkdGMMdm3qx0YpCA6eNH6ofBPRiOo5w7ORxl1akA5JaV2Aidrh355OBoY
dp9Vf3t+4/yLEYnLkfoQaFBf6pWpbqk5L3JHbVyOq/z5KDywkA1ZdCOixin+NdRG
yO1zCc6FoAS+gjzIo9u5bSNzqmMdjntoTjswDUNNnnYN/i7B3B0D1QGsQzRYYoFW
rmAmLJTV5JWaaQtvNxzXeGYTg4SxWHp1hTAPSCMO3S6nbZ0PbgjywjWwnC6+z5el
i7D0rWAFqaa80yy4gMRTc9pFLLeUW+aKnCpxEqAj7MB2G9YX6Tl0BeuVocPpaVNO
61LsAPpyHmi2rbb77WR3iATwAyRbTBqEa8U86HDEMNGZmWeFUqX/usETR4srnigg
n1u60xZ/x/ZVZo5WDQ6fAHMlFh9VP5JS9VjEQugaIlXrdD1qrTq1kmVy+HOmmqR/
kK7d4ajVo0F9RUZHc9csGnoYC9Fymi+MIVaVkSfRsll41ijPX/5opruOid5Ho/Qr
mlWhJCELvDdxTnSx6DYlR0stZFjITXNwVoXdYIBuuBb44S09WyTp6F9N93x90zF8
LJ/hFwlet4K45+UOi8XEUMKgNfXbv834uiBy9m83iN+SLJs1lvqerPpNp4gE1ef3
oD/zRPM0tNx5CUgKs9BmuU0Sy9Ds5KPxHHErXO4gThmSDUFtwrUphtdgDAjQZIgW
f6eMyOyJ29OfPwy4b3UERuiKSAdsABctXrDxhL5lzrkspZp0vonBCpB9HDlSlXFf
shVHGTzTFMXQNe0MTJw9w5OEAG1YpyiLqjdl3nxjgvmfv+q7nkyb0Og4ZE4pwRYI
TM3NRX2LCDlbDxyxWvLrdInMelN0eXsXMalkQvF47VdCWcKmZ3HtpwbGAd7sM+6g
qvu05j9dT1sPA3de2QxqgBqxrcyiJ3iokvb5lN3/66UJn0Y7MkaA7RZcFB4HSAWT
V6Lb8LQUrg2Ci/aS6fo8+7gtVHg3hFhYW6J8Cju2pNCwrafxoJ1khDf7QHwwjqu/
tdedhMblkKaaUNDEdY7oB7W8rVHHWFN3teCLVyy4uC9AqYbC0ePvaD7hu30X0/F9
bQakwJ10fa+CSTPSwuAHXMKCf3CQ6sl2ap6pe+JKMP2UiW+nhJ3qSMRo2sR0oesl
seqhqx/9fJpXkuVUbJkeLYIz6nO7UUTzYyIi+YD1P7wx+j8w9KGq20kMXpdW6KoE
QbXDpnIohl3hEhph/uhRbwdGeHQLMr4ladOgzKV7oksm7ph5ictWevX9AMUo0s1J
qRHmUARfwhaoZhgLv/O04cVJcIvrJU3zlTCQpL+lyXkKOdfbBB1Zty6GrEYgiG1Y
8c9pVRGcNQYRjkfHnYDda8soNgNiGgs8mePeCC4jsPFPKi8435Ik1wMb0d1QHY72
cIf70UvhrGSq7x1CcxZoyBMaKrsdbHUbV8DVehkq6CnUay+VEVPD5KRsH8kUmXGh
8nkGls8OJvUcsvFgijtMNTrmBmRzDQoqcY63J3x/Iu5U7j/BV59cMhZ2zc3h2odl
GX3KEjqqSn3/dxG5ga6msvAnkBsXOmWLkoi1xHGMNuUCjxq8OjXbzMJx9NR3Glgu
0Jlt5Lubuua7xyAZuB2+l1j8mvfFsfBwHidjp6jzke5Spx9VtGAzI/9MOPA8qb6x
Vn4PZjxSBZdyEJVUXyUfsZLQkOZWzY7/5ihdFiyuTJ/4RdOKHDW36cvIagh6mzwo
IRY1F9L6Mg1aTRqgnsLCKbnjttCfnqMM8PbvNXXNe5E2o2lPebDcFUKDTfU/Gc/e
idGwNsVoEaXZFSXSMP+NKpHUVbgBk8DnYFC6anqN1aRQOiIUNRXE6C8kbVeL4Xi4
O+yAZs/jsOaLKzZkKAfJ99KZt95UD+NZ2vPp2GhJr53h+4DVP5G0M0pMYPGib/RL
BYZN5zsjNVuGIrzZ0r6IJ6RXsTWrXBZ96PR1bMOuFdqGxCPriPHACos/SO7RQFSb
zTO4G/nRwGKPm7ttxCRT7m3RVseosgGgNpFyFsjqyrbsy/JF+z2++YFf8Yz9JY9d
AWHc9dAe7WYRTnjXbRiYjZ0P5oFkBv8iUmJi756YCXeOg+rkLqZIK/VRj6AY4gep
FvRfjF33dImp/ECDAEmU2o9CUDQlh6LNrRHhmw4faIMXrPED8zFFoDV1tLezXykN
Axls+T53XWPeQMl5KIBnz9zjNwcifO8PJk63xsAaKBjO2ot3vZZM0c6q/JqxN21O
/k2ynfp4TCGTfAd1XEcUhsdsycwC8btkmIqLldxXPNxQQYipAbz/4EiYliUV68do
SUXfMiFjUefj4FOQAtoP4g9mrLjmP6A/VRD5axComi+7spqgUn8C4CtF+SWosNo3
aLeaBnSgwl2ribsTFlPsQj6Cylm9vLbIn6eLCw3MsyOAPX4bxQcM9s+lAIJHp0Dk
dhFbLX7dl2B7J19psixz1dAGVIUDmRzQWfQaJWVKLlugjlBEu2KuO48+qC/vjEpi
e+6piPJ1olJWgtuOzzlVIdTu0Wsk2++OCPS0SqtjsH7aeJx+is2TFuz/a6ESnptx
YrKoEPK7CBPRwx0jZ6Pynqi7Awl39snbxo5WmYGI02o/1sHsYfpCbG9W8sNkp6bg
jbFFodmDseDUyYgFmQGyRn1LslPGT1MkYpZwGUtBMFymVRT5EMV8gmR2qk7HMkOh
ausONY1ow0RMOX2K7gpmDypH+wpQQMOY2DvmXsyC1pxrPgg76Sw6iM8WOnG7XpM7
Pm0NfJ/22PhGb1PX4SMQneim63rYd29eEHjlJjDQQGT/LYJNXnH+yom+5Tzgdsnc
qir2mLregRkyuzVEvmlNoBxDcuRjzvCTuVIPUMH1QksGCBO3z77A+g3F1wxx4yh7
GuVLhpSa1oHnCztJhC4f+hr0LY9v2pD/E8vYzcuPLFkcJBb2Vidt9z7t+pbVrKRz
VaO002TjhduTMaMB76zyEmG/D1mY+E1cToaXpzn6GVOaqvNKltnlvvdsFNvozxr1
3YAFd10EddbIGahoJMZL4eGSrZLwojtcEl5qFwbqqkjHhLO31Kxqr4imBx/e8veQ
NR9CtbnDSZ7cpK4zT33FJHNS+8jaRBMfbjHCWnOU6fdk8WVt+iUUKRpbSzCanDC1
UnVb2qVo8Jse1FdlhXMy6V3vj7SQiiJeJ3hkphzYxMrmo2pnKtLILtl5G1q0yEZi
atEmo6EkauLUPSW9g0FQML12gXovsDdMLfHdCHn1yf5AsD4gS7k3yZYb3fqW5K+K
eo1t8EfLFKDpthl5lgoh55r+LDP9aEtxe+ye+eOk4XcHTVm9HGbACHkWhie+15M5
AvqeA4TMbyBe7Zzhj2XumTmxQMtqFY+lmXCsfkKEJSKLDn5mNKvASaHjus1LhIET
ScegLUhTJqzyIJKWBdLHy0VNaTVxQk2xRFbXBYoL9XV5+r1jjbwDkK3NTyDD+MCl
xdKaqRxYXYzOKMncav4+QPS+DIj2WIUZM6sP7kicxjeAkpOOD1xwM4fpep9sULPu
rbXDlE+UpudLh5O3aWoc8T0PB+noG28V2hsO6YMTlwPq1muk7+zanbhqdHyGlWrL
hPQ9xQeru//jGNur2LvaMoI5xUfu1WCYmoSUpXqsHVNVmy9yGvlpyFiw5zkM24Mw
guqLRBYphEEV4uPy1+7AIa3qteA+sgWCgsmrUr2mCh+xGxoOUrw4DghtauGQ3XiL
UzU2WI//MjOBvDCAiRC521PRw5DskdkhQre0pKx4IVesp/zIH1JNFO0HKsD3ibfn
55S9W9i/LS9mL2uPWsK5a6t5Z67qZXQSc1jPvN1VAPjlUgLFfdCxkoI1jLSh4ibh
6p5N8u/b+rAann/Bv+vP6jZ1JqziIDo/jWGTEB5WrDr4lCmjcKGIp/KFRgAsXdiE
p1LyxHIDc/7pxoVu3YgJ95I+mAD5tIJqrmhRihs9kOZOt8q5OkOLC6aUVmB0/g1K
XEMRjxG02tVIcG8lCw+4vyTXhp/TtvyGmQ+/SMnmssSIYsu9/JXDeQVJ7gvBv2Ws
b4AQE8mTwJzn0fEAtZewQxs/dSxkcnpDuhmIQFQonVGoFbh62TIM2f/9FlankoZo
rmyht5EoGlP7XmFFZjG4URYKiXUqpqMktgwzXPm+/eWru9O8PZ/dlukjJzH6ol8E
qeX3IatPBx6sdRgVd2FTDKM+ghSVdhJG9glSQHHTPpHoeQDtyhgT4irgQXtgsw+v
PcyuX/9UGjfJ7JHVwra2+OsTaRX2SiOCoaKjsP6oLur6GydtlyYaxe+DXKFcdNCw
WCszu78qxh6ip3Nnx+djS2+3+sBw/QyQ05B9d4zs38W1piht0MLNBZA/iAcbLVBh
M7J3KmXxNRetMM0LEhvcVePMtTkPhPjG4/NzNQSNDr7IRHP2lG3lsoKJNQo0QZWP
78u+Og76hL+/UKdFrsZa/1hmCiD9qQvPxzmDBih19h2ji263oipPcyzX8gAhgl6p
Yy7xSAEOs3BO/+fSMYyYwIzYj/9tnYZvNQcZ3rEAo37AUUOn3lG3Q9Lm1kT1GOYt
DRrGhpTfm147eXk20w9atUGtoa5+5Xolix4g45pBoPXaOloiiOTZ0xeKL7tVyIaZ
w6m+cY81iGGVDaRUgsOubUovW885DQo32bhZViqUP+0BjHiq84I/C49zO/mw66Tf
muKSpE/xihsPXCLN9lmBp1WXMwmJEgjQkj8y1+rmepza9h1r/5Q7RBb/2d75Bwns
gmFa4HKcJrS2vjDDNaF738TNVAmU2PrVb5Aeavh5faO2WtmoN2ieHfKpMIxqb5Q/
CdUfYUdJkdTgN/NlgHrmcftFdn6UJtbRqvqIp0BwWkR5yfUsj5YdgAP3ltfMXAZ1
gizODwI90FRfeZgOQT9VOPTuPyIVoZO65YrLASuUGU0t99HibviIzp7a7cbcei+k
7UnxVwS0BVwqiLsBtErKufHEdp1AVWvn0EWnx2sncaqgvj7h9ouBMKPtGuq8CsYu
V/0Ox5rG0tDpFK6ObmmULXDL2J8PIVhNuUd+ywX+EeMcYpwu5kLZTg8mZGkYN8vs
8CgrPa6oM07JVQPMa4680pRZtOdu2Tv3mE0eFHRQqMSocMuXLh9zgBPK27gKxfA7
ZPd9v7jYcf11lvk8NCNhRAnjaq9rpNDH9HPs//dF3l8MhJMh4aM7vYC6IxBzoiG2
I5KF1KUmO7Rwrso9cyH4hKz+I5n9NOjTvTfuDf2wbJLAGRD8vtuBj25JJ4BCJ/zb
xUh+O5pF1C7YDPvPcBKtbDQ3rUWXfNkz90W4mMhJDCMK8My7i3tbDKMYA/J02mJK
2FD3Wza9Xp821M116/iMdhAhMTOr6oB7m5RKUGD9/DCbFjTxk93BaMzyMwlGpASH
1uAX4Qsv5fmfK7c6b5wx1p3iNseh81KXpB4hcnOYn1nlKklp72OjwL/lnniDi0Iu
wevS+TVOO0HLVrL5Mc+F74i8Nzd6nSam74mHyusli/o4I3bvE60sdl4TDRofvV5j
EY60gJ4haEmjqlZNR2EOi4NMTfsSOLG72aGfEuaLkhu8xZC2+b5n7QQ8JWXgOA6a
BdJohpgVDhs5LR3+WOzuBws7j+hyGkYTN6uSXP4ITONfocU9yCvoxzWddrvdoXoR
Hv09TDcSoJsMlsJdmGNTlUuAn7b7i6iPawE4MnvFX3RWCBkpXDXatsnBu4ad8WI8
4HkqdhBS3T/p+l9vKd0kgVaQTaJY0WDdUOhlYe4wfmR+nRhRCFF7IRp2y8lo7Q3C
awe5CpD4bvlsh6aRkiQ9l1onY3DH0xv+Sxe/lzkytgchB2Ob88bZOSdlpbSxHDEd
VzlZx/lQzvCNG6SBWCSS74Hxo9RwVD4JzHGt+sMKXmPp2aL9U+XTpqd5LmyC8Rig
oFy1jlmRrY6Y/hO94T9kLItn0GvlG07NUVKGBfuhJ2ut6jKvHDBro1GSmka++CpZ
X5yDHMsre3k7J11mzyki9jk8y0bwQsXPN0TngaMxycv/+gtBbwqRN7G9OCyVX4PU
eSubAOESIMwxqp1OiJ/gpOqMQYP8luEtA73230OUZRjmGApt5irMAKEWTU9jAHmE
dQFwcTQ8Bt/R30sOcQQNyaJTABTlLh47sKTNQodyVXHcrW1dPacOygbDfnXQnyAp
eEH+EjUIBCKOz4s9ZbRz7NjkqG6csdBRgs/8eLhx2p7XKnD+PY9+QSNd8z4qv26j
QAWuBCIsyxTiSsEij75KDUdVhbkFwHlolJP2LVfPLV1WMBcyze9N0JiIWLBwiH8L
mjBq/sMA9Oauc6jeMeKDVgOggWe9VLOBpYXkc4FE+NceqYHJIGTMNnnWAK9azT3K
o5bUadgPHpgG3pRVQnxESUYyvBUPxWd6CtaSiSQGFFf778/1v27rFFsurOuoA1mO
P3CftULQz6UJN8RN9tk5ACsGXk/iPnr8xujPKIH1WtDD5UTkM0gSuj7Tw0l30xFi
mbxcH23UZaT8C+WCnW9VrQDg0YZtg4yh4E/FD4hcqzujbSEOC18uT8kTKtI4YQv9
kNX7keYN9YcEJw1JUBGG/cs0cXr86kql2mTrHSziZ71NzFzZuOcOfguCajqd0iYN
U52Z2Pu9Jge/vs0/Wn/VC1cbQ9t1eJv7iic09PIj3JN8CrdslaVD7GEEs6FszBje
iqQEttoslOE+LXQMQNZK3W4mk44eOBHZK3+NSD0Zx8pt19R+JBOpANZnT+yZNglg
osal3Q+IyiT1RU9fpF+rpTNi/u0fG0a4Nom5aSWwNNncs3LUEgY230jsdaKP3SHX
znZG0W0TpLgnb3ibbR7Ox8zQHMsPbcaaJ2XqzwIaxQx7PVpwoQJNBbltUqd4cD4n
u63vtqE/RsiRzZuMs9Mko6MpbvXmAe/2oLaRv3kiedcbms38A015XJGf0g1og61F
c8kcd0RuOvVjWlXrt3FIFUP0bZXpQiYxo3S98p+MDdnt9bPZe8Iu0zZcfplTWVqB
u10adYtrhrctTkr9w9AVtGyP1SVbL46LtxKqjppmpIjFvS5zhXGv3Nm/gxhFAycz
HOvmybGCDYdGd4/1rmj/QikDsTtpWlkCFxVcELeitm/NXG20RFnwM4Wyarc3Hyrp
3qAnMGRnRJ9r39PFMV/TpX76QzI1I3hqekdzs+Ns1VXzLUavYGtPXbGOI4vboedY
uJUvh0hVm1ojJAnEET10E7/TLbKEaotQQP7j/CyJea04QW0Uzb55IPvyq81hsWC1
R+eW23lgXl30XXjFGlQV/zl/PRrqey+GPRIgS2uO1gpHIsP4F9DmTrCl9csdViZQ
NdfUt2x5XcNEHvr9oYVrUuEF6R3rEDvRG7VxlhhcK2E8RHlmrT+Cn4QENd5zzRzf
YhrjLG2sfia/0F5QahSIDU+cX03uA5qiTT+FIVuvtcVRsjLhMJNJlevl2f0SroiA
FC9Zqfis0JTlR2XpTYP0HUIrjMPiOG8aKQFqF+aTXg6vZhoiA1JhGg424rOoyMha
+kTlRfk6rrXufUukbZ2Dt2xm3DPF6hwnE6zg473Lenj0By0sOWW9OUQUCt15Hl8w
Z5SJWErMfm0ztOXe3T/862e0mc0TyQJipnSrKeoWGqLzHsSFAFQOQZaq+2SqPHBp
RDxdj9s/QF5bhJo6LaFXM16Ymd6+iAxGrkVIYW/jRcg6R8iXq5ADQDn+p+FPIXsp
IAZf0EgR6k27fHhMsVKgk7ipwOTuDBlK6XIw/7q9nqSGxaOMSxvtpJZpJWf34vg/
gXsuxJIfyCxzJJu9gkvuaMlAJia5ObkJ0RZxdUt85tJ51cBFp4y7MPlqmM1Hv0yx
xi3ZTsk+V9oqgj0P02kb4CpZ1IF9243RZzWbfFP5sLdEUi8UvVrkAqTetrpRKbM8
Ik/A1yrJvaS/quRc+cahLp8oqzbjaTtP2hQBkrhihDpxbXDmXe7uJvFkUrxBIIZB
sUaAK9OPkDp3A26dmIaU71abRMn//oqHUWnbpm9rOh2I+EfpOldyS2T64sXExon7
uiD5YL+/Ceclchm9gmprQYPzlM4NCFp4sEjeHQmMJX31HtEAQUt+K8BBwzhBAxi2
epqYUPXu/kKo3YGK/AvPoWiDYofTQx83+3c9gEzzciXtDOhC7CYyP+vnZK3kPDCd
IqCcjllsaBS1RWmQ+PNIlQvW5Gt569x+cnvvp6Ky/MtNj/cw8fmDM6Ze5tCFubBc
PVoS2OUzLn9MyROiOZNT4vbwHwBzVXL3KHWd5vpgxhKFvLcwfTFNaj2f+OZ3mlRf
wGrSkY+nqALb5oaW19FpqzHLnMMufnqEbXQ+nc1FMlo/6spoU8vyxekGsBN6ttvy
a1rdIegwDh4Un2sF+dTE5il5QKyYFaEBVD9xW29aQrfJeMXVlP8T45CM1PE8QRr3
k/fdJggTLFc6n3V594Qn1332k8DoIiUKAKcSvwDf8NfUGTMRLww0kfKaPbklm9rq
icBM6elydfXfiX4VL4ad7HJdbws13usrJUSMoussPZidtAB9QK+iwtIEiaxePKMH
wkU+DGoG+rGuuvsELSFhY1Jy9fK6PUAEtbYA5ejAvWWFj/8YobU3kHHQzbmAhJjh
e1TwHRq/w0TaUf/Drwyp/Qx5JFzjXJ7feG6ng+7Cn+iMcb3zuxpYK3ZJu80jJbTR
yaDxd/Gt3aAmEe5fmpPCGyKgt9It1f+RTyD+ze67G9PhbTji4kUmESYB/9P9i9Mo
5elkDqjWqX/Ik7sWrZmYHEdY7APSvcRzHlNCEnA5bZofKfP3SjzvSP4xvPs4qjsh
HGwQKBh4ulSRFk+dfrazA51kf4ub5BdN4BBkD9K609IbA4afJ7Ky2HBj8gZyClR4
SCiyweyNtp6albS0UNNBlJi1s5PFIcAZ5MLOzEErkCQgLugjHRp6OPgsSHZ/HrFD
Pl7uHpYW0yekUSeMzgl3ZkbDmFCbjVt3JsottVk5YIef3MkCzj27UYd6PL9RDx3/
cP9KQF9g1ia6xPqXXjYRjXdFGkj1mV+KFQoPFBQpFiMmu3J/Jy+Z9X/NfAqwNpW5
DSdvQVByvJ5N5+N2bd9lDgSe6Ksn4jBe4s1JsxnpB35854I/er3QLEsmLmgwxtop
SSfHXz0m+LaTB1McVA2/ks0XeKynKzfrrMGifb1FipPH7ZPRDTxPVIr/0+yCzALI
bgZm4mBC+dnhnI5nEwSllbcMqggTEN/nYclHRK3b+wmgg0qTB2JmChYYVR2AkBv7
kfEt9RXJiu/qwOLsC5UXNZsWziwDoqWW0uem6NiN80+ZG2b+PXBREuM60bHPzo0q
WVTor/NZDCQTG9Y/zvN3k479Zzqa0ilaLACtRk625vAkqniEYb5Jwad7jhew/o9e
McB3CjDgRCNQ07+tOFbwVs03/8RT6YSQnSGCpew/69ZwL11DE+F1kTL/lVqHswt6
ryMavGHCRDQdIyZhQBAr8NGu8BzY3BPotrQ4vdRXObjJjTcZkjf9Ccs63e6NwwcB
I50TpzNbpfAsO+uOpyvPBZ4XYwRIM4tmYRN0C7O5Mzo0MB/d4sSZd6qQdKgUq3XB
MoqmbYQRk63FY/8Wtredmcz6La9iK7zq1k/jGECKLFihbcdCd2UlO8cIqOG1Jmn6
/RO1pS1VTnL+E0km3hTVp9rcLr2G7HtsEs+FUpzd6B1SMfpKgQf48tzmAWqmckO0
vLcmTu6JdPcTiMA78tiyaWpCtexYmqam/QfZI7ZKfG63tMexiEtCO7lWELtjWvGv
F4v/oFsgIXL5gKQlXNbLj98pQ8cZ+2Cp6jb9yoeqLHxGRlUOeAkHS8DrjpprUhVJ
T7J276OXsWJtjn8ziSQ4v5UnSnqxJAAB+gY2TkBf/thKyY1AIgu0NEOq/a9BQUxj
nBr39nK9nMiExVd4eow2xW5pCgarcQBw5BbDvhlp6QzYQfzl2+mReoA3fo3PQrtE
FdctR654lpCqBPBtz20dmMg7mwmVT671G7fgWMrLLPe6b21CnHMQqNRM/IyMaKd2
XG7wkvW5g0McErK3GQBDZQWDv4YtM+E2XFTRR4NZxqQ/ifoscQz2XYurjlWlYFql
jW4XnVVuM7hVlSczSgQ9IIPRmxlFkDy2xlBlTuc2vl+ZgjuJwl/FS5rfgRg/x8hx
Nvnkj6n/AX1+aiW1EZhXCJ31kJzzqb2qyxTKWzajrs/oEwKpqk50JHm2Yj8CnpxB
dtNUmDhV3nDw9lY0K4z5cnt/UzpYowfOjl4BPLAzuW2PRGc7pbgtcnfPnNnuC5CV
QPa9M9vZJezGChVlbTn/ha2s+tnLNhIg07X51/pFtbcIvgIdvD09p8zUV4idiW69
+2yIGlyV8+OEyvCA75wRDDh3tgGhCed1EnQnSt5eZ/YOZ1DqZDdDomFW73Uj8V36
XecyDIxszdtyqvQLUSn69OPo/FvvHWr/rDsljDFP2Rjo9klI0hhYTPZsvlma4DyF
0R1rjHMNXnDNEqC+0oKHHDeWU6I6OeW2bY6DAExNv4xcTXbso0zFUJNf5Y7dgdTc
cKALqk9X5SnrPJlruXmL7ANZIaPYfea0yO/bWarVfRC163YRKe0kZmT0ovMtswB/
XQk4F0iOYymswsvAXGyqPRSAK8kuSJJTfcAPW9ErRkzV/KtaeeZ47QeCWSj92DKG
vxuQ/MBktRqmgFQ3DzdHuefXjStdrXj6Y8apWBPjEsudK1A0PUS8zNIoPEBvrXLN
cw/To0AH6ovvQO1+1E/Mnh73o1LeLTvFjRRKIMBXQC3KgFfsFUoSTHSmEKlbm6N2
lZ8KU1rH1OICwqqgIZ+aOl63C7ajztblweWElhHJbfLb7nC4uPRrfDc6WpnVhVPD
W5eU0uFekPQOFtAg2QxEMWBzShMEeptWMaKv18nv8RkxCDtP22P4KmNHS3AAQfDN
QkO6CN/Q+2o+dTf2tTKgMksn4OeYFTo3prwezjbl4WvtJaFwCA6TqRllSneTH8F0
2hO95vHpJzpLXf/NW75fANfA/hg2NX2/3NBbqm5+35ajMrYtzcjURpo06MZK77RI
bNHCUOEVO5/HUkJJTXwdusOntc+YSO/uo58GqC1CHIoayqn1zyD8rr2sERjviTy4
x3DHMjvAYDr0UX6z/JrP8GyPVo+eSyrq5/Xkdp6exznRL4TN2+vPYpZUUeCVYlya
tv79iFTJvu+qdj9MDr0ydUj0sbPkLXcfPOj50hfn2+WMoGdGySu0rd9n0en5ETQ3
gXELqeebREigm+a2L9bq3y76u1EBXjvpt/AkTyZtAmkRX3nBAgRnbUKZMcBkEUAd
qsii/v4CQQrdWS+Pr6Bdwe8wZW7v01E9LDfvVD3c+WHnyRfBnrASPMJiL29e5NuB
y1pWTthEqWKKuf87MoFHRAxwmBglaRqLNHOL8sD11MkC0WbxxwZrRTaB1YHs9NKA
ekRnCvuZRGLEuVcOlvcqBC5gEhfhAswO+1jwdALpOrtbyv2NOuBMl/q+Nz89tm8P
k6n++j5bZNNYe0ZV0HX7zsDvyZh/n01QEBGhbWFDPBAvAbe7vP1oUqVbYFdfmVyU
886xXZDrhZESHuPECVr88opmn8SAi0dBpOAv/+ns2rYVOIAReuXFHi6QYgzMRmd/
M7rZ3965Lp9NwV4g7X9krXoQGZVsXopJGgM0UC6ZCL2VTBpc0mRHI77Xfpw4KjE/
gkwF5U9clE2Ukfdt5l/TssMg8F9fQYS1DEr9jMJdzD+We8LYvxMgH4kojbV0wyAe
RUkjCGLhlCY7Z8UKI6yVqQt4bpt91d5zsX5vdbbczE88Cc86SIlesayEKodfP2Q4
gRxXeFqkidWblfio+uvEdxaE6gEntgF/r9JWRy+TkiBOOtHZEgjMLg5QDSO4g1q8
49eAWDy61bw6efbfzf5M+a+CGrRumxp5UJ90wYCNIQUdMnNkMXFG1Sa2Dcj3Epau
CyvRIxRsJN2Ak6QkgU3xrvMhxZDawSP5mxndhfeWVYr5OE3JPPBzz14A/tHwvEkL
eE0XhaUR2hiXhPFPZr3g5qLFIzNtmSY14zZdgpuUusRQWmx5mfsrS6ZLfLF0+8ib
DJRfogotBz+LloCttpobcVwbQ1ABcEXLioXVWXnsEVquDwx8pqWIm0Dp3Hghc3m0
++jRUSzwhYz/i1rc5aHATRT+GyaH8gnsa6sbAj9EbP+XG3r/m2sZAgccbZH7KY+i
FyvH8Q5gTpuWzBJ2y06zq49SLNHxaz4NfrYAI6gixDCslltvYbGM6TGbsNQXGT4s
mE9qnhs84kNNmpK9d3R5INbS12FOZONvDIgI19xDxquu556YPy6LS157voKQaT6x
ija7/g+UUgY2pXE8Y4fETr2MIzuPQEUOGy7186OhMMUpa35247zEEAGQsqjkeogf
sBEMVb4d8G1BvfdMPUOKvrGr07BSHn9pJgI9it/K50LoEb4uHkEaD+uYBY2+VWKm
CUvBkhnBZwgEmi9H1m7pD13AbjdiVg8h+68jP+X8x6Q+OKI7Epffw6vl8ijTTDbv
lXBL8F2fM596qMYeycREF0sNWTRYalnIOx5FZOet2zWrbg4wlvsSuu+HTuh2Cihm
elq8/vmY6e8qhvSgjrlJGs1XQ/omX9gWiNESUSke8ZheA0+K92XglhhmjNQJUL8Q
NVovIK14KOTui1y209u9tmL+leQKnnuYfu+rG5zsKBeY7Xr84gn1bUnjLCDiGP2K
urYwG75u5rV/PlMf27RG97RLzrABF3CIAjtUJefswtGKW44nCoDKu4Zp0WLLAkGb
B8JnzbS3RRVp/PH8O1ckvQtYFDM46NxiwFTzJW5jrQTsnBQ4ji7lTl8APUiA5DQt
iSqCMaatVbXBksXm5alrI4rj6PA8LHBbqMDiXdj+L6rHxeY3KdoTMyNLCWcxX0VQ
A2+ID27q0lHHMnj42SM5cEQeJErJhuIttgdByesbRMgM0cridGsShaBvGBW8PICF
75v7/die3F0kPvFlfbRWcttu1PWr+xToTdpUMtRUY1P9i8LfrG7CFtft7X7Bk08O
jCB3qIWMwAvxKdKcS1dQ+17RGYfOXLxpiKzHchhU3CCqKI4kcV/SPSSp2bKtJGjz
1q3GVjjXGaoSGuPQ4UqieyjOwKO7V/LFy+B8PktiS9xO7G1F1Gm3FPTONhh1lrEa
ivcqNoeGxGPd6/Hp9Or4aZuwvSkllQllGq5XBQvCSjNIzut6xVhAX6IZG1mxtzSo
68zKa7uW9wPfCw3sfpSK/ZJt3LtwfS61koHkYEiV2qi1oIRyteuNjoRO8j0HaqOw
9ldsjcI6gJJHqYmkqPk0fQY798qEO6DSYL7ccSSMOHSxhyNocR1pVzUCUbo/L6f6
Y3BMrYfMVg0u02+nzMLdoiGtdsp0iue+7F/FqzSn6DCZuS46Bp50x4hyKwsA0GD5
3T+NLD6EXrjP9M/FbCwTE0Iok76bfGN0bMr1pyeXaBHpcx54VggTOvNq1wwIl2k2
EVHu8IMAxOsC5Ya4BN60QbWq9VyzIJnHBFgZqKZdjQe65hDnwcgTupKvxSCTsUjG
E/W4epTQpJHPSTvOrzeoxl06+2Q9dzqoV88vw7rNbbUaiJAZQVUsXDN9Kqxdgodc
esBP8bAIRSJBsHCfaOXciCxg7XHFEhHcC4W8jynmgza/Odc/keKu+dDNNr1wLkkn
z1zP9hWI5CO3XuaoOuWwRAIk8y+gJDsJB3p9ppsufUWAfvpWzQGm9rcHMmG9Iyrd
Kby1OBHW+WUiFw6IlH1sv2sSlmxTGcHsDYpDrGj5yDtr6voQHW3n1UmmQCGEOCmd
TqUMpX3MCNEykhCXbRxJubxB2hIB/ANXIjbCQv/TbkeLUMB7iFNG6RnNNco3/Cl4
vBeGDnkpG0LM3xgBiiNegV9ADtq8tRZnTh1qOI2BoZap5x5S2Ry8f5zMcPw0JKfB
gO2tyAjknDOQ+grxoIWe1NGYyA+qduzMKSqzyJXNbBSpJ1V8eokWJrDO0aU+nwqJ
mDTGlQxRRF0QW7rVj73AIwYgzZbSMOTlpfunJhvfAKOfNIpeU4kZOU8TqXDIIaEh
Wi+Kn/e9IloO9SwSX5u//Fk6ib62NQmvq58k/F9mnk8O8HoQCPzq+1FKqXSLJncP
dbEYN2TRGE38kZCqBooMGGzN33fk5jAhP/sLKN/5X9v/S1ZZsKKrEnbbthu2jmbC
/LLZO1RU4WPs2Z42q5xR6QRkfoejS7OTnUtl2tVDP+i10aUlBOmDQCG4bVHOvY/i
dqCI8PFOSXM3O9iUMpDUSgN+oNaGXNyRLoVocolWtq7bw+qYJ4c5tMitnRQMyLvU
IY6W3yPu8OsWtUtAklF6FlBe6xEfpfdu5U7XCEhlMhdd8frUzg2qAsEetikF/BXM
W2ILf84zKH6JDPen6ZWTG3xvb4djold4pm53AliVoQK2VHFqzt6r87p+WRYmIiYQ
b3lrP5m6kcXr+XcXVVSaouCp5ZMt8MLPURyIwfK7O8gNyix+VJlcAfnP/TlBErQ0
7WFDI1J04iyYcOvugEUj3kIB05bJvgJqEU5RGIs3SqRNyBia7yPfrLm+TcfpLN80
FeiI4vmHvbbZAS6OhEdwjT8wBoaHbDUQ/I3s2Dkifrf3+k0cTwicAzyH1fEfnFem
fw2lOBCODEbD/JRNbmmHF742G5rKHZFFHOLBZyyM2EYVgeYCOX5d4nhtt00ob4Py
yorlPXrimrhahRqTnndlNI3pF4Cd3Y4sNl1oW87AVJa53hilGgD+8I8jkqXfsL/3
M9i0cmtr/LndcZLM04teunDHqNCm0bWMm0mQitWlaYezZ70zlRbNlTQjrgov7FYc
Iax+vd1BvhWoROZ0tzU/iLRJvb1v0g81IdteD6OEfBjSrS8BW/mKnjNLmo1wxjYN
M3FCBY2cFVzC9wHbCf6S0dF7Vd78QtDQC7zBzy697xRjn+wumhR71NTTavIWwhCF
fBHYhZiUumrJV+LH6zfODEtJReVq5B3uPYsIaW8Shd6UV1hsS1zdm9ejJwniLC4T
FVQm27cN0YHzkxY8JtdsLMugHvGnJGK8ZfqoKi3wjJfrmTMnvnc+m+U8zXx10xEn
iFJ3K72YGYSdpQY7L2YbLsGxT1f9rXjH3tJVbZD0N1FKLq+TNHeWsn6uY6AQt2YN
stS2ThXU7YGfYmgL7uzquDtgFSHqSS1pJ8Wh4oxngEjUn7cAbFv79zmM0tX3XIgm
GGob3a/JyecU0d8YFi1eRVt4XLDIhAKA/HsIiMKxX5gwU4nG8S/Fz+Fu7a02DoFI
fPdO7HfauSwPh7K/t8oRwMl1eWs92tED3owzHEoZi0nfv31/2E+Ws0305T0KKiBo
Cryq1zOCQzpdn03ckPEu8VcT90Fx9Yj2uL6ZCidn7Noye7VWoAQmXRo6JfhNaQLZ
9pYqaivexWDfOtBGc4ARMV04JIXdZJvxKGEZSvxchUWczy2BVFiff2u04GYMt8nI
H4VOd9vbm2FrONhTLS1WlPRJ2bLrbK/iu0QhlE93BX4Loi/BNIbSQ5jXMSzC7ZKI
miMxGJe3RxBo6TBfuJoe2o7bxrZIuA7QNfLKqL6JLFEan23Noz9IQou9Dj+zsGK1
DhthVul2OERZX07mtI/H3mxMgGsEfTG+x8foSF7BUNm4CmTQ+e0MMinTj5BksBqY
VqyYPaMrfWFmt7J4n/snJtjY5IqtPqH9twLwObIQZJ3+EquPOlHkJ8udh9m1HNS2
1eEEuav+8ujPVuIPhY8jDVe1Yum+9CIzF7pHhHHtJmH9BGsTGqGfv0RFYUlur5HI
hEFxSWR+MbXeMnYi82BFEUF+5+ylvAAlEEptC5zOnlMcKENXbxiuQ7drsEVHSxK5
phbDxyCVwfhYl8YMhtcsMEDYRKUTHFD1f/WIZV/XvnLSamrsb36O+jeStRzQ7EzA
K+1Rlul1lQQQeEtrWwmLk1lSflq3SRqUPKAwlMz1X/pWosmZY0DXKORXCmNTYCen
XhOjPmthYewehA+M8dCoKM5xpROESa7aCRWIKAfKWNdstM9mdEd0ByPmBxRJGasM
CSvQFTOS38EESPHFMFHpyeEXrZYuMNfnsPrzVpvLQmJxCPlVUVjNbGpl4sSIX5QF
dwYnZ7XlNFwksrR3xwYXZe1NkGNX4UXESMcB6ZcveoimQvl0+HKqJqG7BgirJtPx
Kfg9486TQZiIoAibsaJgA0L4qF1t+++agasIyZ06twZFA0REKFhLv/hBpArf6NpF
ehSVlKhvsDWlHgxAK6b9yyGvwgQFf7jIZ3VJR9idmrJ/jgIi89iqpODrQnRC/tJb
294GQU19KBKnxS2+oTqahdIhkXQLTCKJK0pC7gGfgcngu7D2QHCGeUHq2Q/h279R
25pmmxD/Ax3/heXkW1F18bue/nMbnp94m7KMzAjGdLaSza4K8RjOPXp5ErT7DQMq
1oYMqlUHYmYlNmdipfuxezR9mRJM6vhxe0mtON/teBVbgYyNZh/vVXEQNbP4PDdt
iMSkqg7N2Qh24angBmKq7h3em7RKRv7/YC5vBr2rR8Vrivj/Tgk7ens4kWQlHO11
DhINk6bEqZi5AC8GHn18JSi5VJZAn1ZCP+mMEI/QKsJOebidJSRw/XeAZYDw84g/
BTgTKec0QT1vfv3/EyZpd6K3ONE+DiTeHIlRjMcnnuQZyKN1RtgKVXPY9Ia6Ca5o
WVdroYPhrhQn+u84yLXAIMwkMnVZoSdv6JPVa/+IzOmdCE37WjVkS5Q4k0KafOau
IQnl3D/+pcCHSZVwrrJqRFesBuAG/DutxaeL733YqKZblYKbkh8MtCZL+H+lhF6z
ItcaQRJOeaXBB+CmiuTXt3wiDn4VTcFZJmd7NsLXcWKEAA/Ap+BIg0ckdIO/g0vT
TN+4RqmlhGfFc4OwAKrVbe0WbbfdXsyPmGZQeeVpGOKu7q3pg/eBm4Kn5gOxss9Y
iTzeCs1ctfUbneCJvltiGWZ40b1kYHZ/CUGpQiFiDkQtqndbYmrHvVpr9fNvruXe
NbRF6UO/EgX5WzHl0PqKbCuN98Ltn0V4a65+Ds80Qd+sDqX+1X/mKqVpMXQWwNnR
G3WDUCPJcn8E/W9qgfKDAYmbJB7mOFVNbsdMqDx26UoKlwNMsSvvMUgl7R97qWe9
dpYyf1/CxDAE18ZcV2Y2qKADmCjQl8W0HBRZHWZrZxyPD9ObAQX3RouuiUpE2NQa
Eocyqy4spq1CJGUz/BxChgbhvWAqRxFjvZ7cypcbTY8qwPNUGfHnY5eslt4O6B7I
83ulJIRiZ9t2ZbsGbuGKcbDQkwLc2WrfZVzKBGiab3d8Iodp5b0JJOwaud9X32nK
HzYRbiK8z0TuVrtCNzLHXVnuLMjcUusxDz4+PtF+KSAG5PV+k81eeAFXYYqzswIy
jgwI0gQBDqDhzTHhQnrGmyFa6Lg0lgj+bDa6UOOwxvovJElsHJt/V5fT7Tv8+lsA
mY/fABs2iP4dZIrpoGgn1CNs6ucp3jBFLTFzqdJq5hgYXd3w08LrObTzaEhQDVN+
g62v9fPUhoKxFWePnu7hD7zWLM0mukdkudLjqOlVkNPIzyJqxdGN3oqnotgmIBeT
ZQ7BKF5UgyeTjFCMFYm9cLbWVLIvOFEE8Av0jmQKM6SbyQ7Xiot9gd3UGtO6HN7J
Ci5puVNl7/zg9pQ/mLLtAE0dxzUOKnM/K8NJG0m1wV2116M4icdYWll+A+borbmy
U7G/WvUmj1GQa4rOlmGioO5oHTeF3hMDEC+oKOIB6he+ySgx1w92SnfX3mVKQgKY
c0Xy2hNWR6acak7y4/ihkOJ5aagWn9u56jWIWznHRDKfZKhne3Cg3VSz2EivtXEo
hH3xvz3EeM/CTbV2d0AAPqzRqfQVycw63GH98Lxko4+d2Ko7EGIdxkuctTYs8O+N
xe3//ZWvFqZxG6wyiZDRNJJ0bXuu0/q/QZ9cIRrDjruiyA7jD9qzG/JKgDWtuefo
FA2PglmhhOHtf/QUIT6ZtfSfUdq1tyMt1agBhNNG7TXtezR2aHU7NVhipRHuGNMo
fRf3wyjSpQuYlxTf7y/UZaSxAx+tFUlZAhDdPN5rtBMRvxWp4iGbWQj22eYy8RqG
MbTHXjI68ydQ+VZAKWzab8s7H3qYgs98mFDexTFsMc5OLIkernFieYPepzaGECmR
K0FTLoF7BdHNTPOxwumtz+DxewLne95oO18DHiar+NzYZo8S0ONx6yAps7iWQXdT
Vyp5gY0Bm8kfUHm8bx7CSxxpvCpvcY6S1et9YCvkpaKcJIciqxlpjwKjulGZFD1h
ILy4efckXBalGGsmlQqUlaAhgW6DDr9aG3Cnfz0am+Wq3jsSPQq1Es/qmI9sXCOO
I6TCn1gJ0HjwOFcScXDrdtRYsbIwZtutKKoo8BQhx83cPFEWkbd3rq/5PMcO4+zd
O2Z3/i9nmd+5D8Exk1vtazZyxYo6LHRANluxJnUSTbGfQ1uwboPnEGAuMvDTtA+7
o0QtZ2n13oWuarNJy9T3q4mIc9tpFj3jkNyAyiKEv6LkAFfCwuZkCnAMwr48w5y6
39ZiGlVFRAqNREnCGMk4PvfPHVY1r8sPSFbD4sGbPZz7/WEaPxgIpLOWwXYgK8Fq
+bKaocmrRTslxoQGNmrEMvY5vP/M6l3ClS4htQbNWqBxgskEIHL7fv7n7KT2sQoq
RAkXsOCG4yzyvC8XbSHkFwTv/jcWZQdESzSwx4V/WcLZKc19GzlzrTMhxrfN6Kfa
wcLPPEYxPmsBzVJQg4uA1rO39DlQXeynR5ItIeS5ZY5vHsiKLODUwPMMJCiiAF+S
hlC0dfe1tOfBhWq8Fy7rQYs7A8b95lKye8t4foazPQSR+JioH/k/Vqj/e8lYBKrf
yISVjZMrR0dHEazTtzd2f3Z6pXguZFJzeyx0P71geVoMDoQuarD2NvJ1IOcUG1WE
ptsuwdR8JLQ86t/AIaSt5iOcC3MycaWxlRnCUqA+MVstMCUNjYxhu0HuzoFttUP5
8EZvf587NoWEKdiF6KxQ2ZqY8ZAmeflwNH8mPtfyhrWUwuDdbXVUyZa3G4rjRKjs
IsSsjffHgpRdU6nJdsBpnnIwnBjmQnGqS9sBpUG4Ex9h13UUgnpHubiU5sjsCt90
jidJ4vMFYILDooOJF4j8h8jleac15hSzQJVxws9dXeybEA2RDzF+pkhoyiuHSl/8
i/OXupYUm0myTCu7GQkkznglyhb24XFRyQXXkzc+kEBEos5NimIG/Iir6fJHAYzC
QNWmtatbP7bhpwv7oir0qCgeWbJBkVzRzchWYAc+/+Nu2b26wxUy0LrpycM57B7y
PTNLDIRDLsnRV020aoLWnPo5C/RlQd9axmbkEXPSifhugHLTDzfAU/vExDbZwllU
Pxv3SJvWQ27786SLEWDfYD9ON3iKET4lKsfuG0y4Ib2smGKr8UXVdBhlhWEHEjEC
fXhcBOffGoHnNzajRkgxsl4Vq1BUj6HPB5iARcx8Wh4coi/EmzqbQ7pbUtppbmdN
KZvjBnhf9rC4xdRYtWWNGwEt6Mj9w+rkytVwdVqDUgWtH55z5upyumRNVj4KJ8Xo
T2Celm4CooAatvWpqZLm4kZ/xB9BPwJwl7kqVtqTusrXMM4jqqNwAYYvYF3NOdQQ
86oPKFmY0Q+rw7sSvv3OjA==
`pragma protect end_protected
