// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
iRP5A6Lt5/wiK8gkn5vTaMqyHjdvwYgkHNr7ZLVzHrGozU+W8R3lAgu6Mkg3TY1s07lVISLXouT5
cylicl57VreVdBvd1JEfUj1Op/bhVCdknxChAT3O2XfbEFx7SBpkzK8dry+wFj2CyAuaIJrPFpy8
mSmmXBJ+c6EA3VYXvzf9NDW5B4kPNRhp8/vFhSEMjk+ZxByRfxp/jxLvA51Midxq4zLh9JXKWJki
20lyqBoaqR+FEBiQZsPuhreUyCRxq52rPprfgpY/TRh2de0HSg0vG2NWszxIxAO2u44Sc6yA70ei
k7F+IDoSI6KtvV7T+tE58iZ7PX7uijl0ZYK4mA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
GSeTbd96sY1WWKwST4LQFZ66Paw0PDPRlMVmLkYw/ZyG9KpvogjY0Kd6dWZJvTs762RpQy1gUblg
fDYRIRCQjCLX6r8mHaEpb1VD3+v3Ur7PqsTH2o1ybtkmm8/6gLmLWjZXUD1LN4AM2/be+FqjxcqD
K2EuQC59Vd+KZiC+wz6DdZ6V3gngctFdwsXLAcAZddT4vyAQWZTSn0WKyrsB6Cn7bG8I5QYUV63U
9KnjLKiZSMKhu4siBn34cWtQsGVkXDDto/qAQMb3CuzNP1BFS4t+HFhzVe0WYchEyX+aSyvSwarf
Qk+mRAt+Bc/hHJLKldHxYgxOqIfMq6ZYOk8N4XuT4Zt+SMDRJ59cA+hwzZAzYa0mhWwcz3S5dgt7
ukQ0W3vmCf4XBNQh+995u9pkDhCHkO8eC9KQ9/mL1F4VzwIPzaCk8mEEEdoNhC9td1Wh3eWJ8sHn
I7i1BKBcwfIT0WsdMMunp3BO5KTugWSXQImNH1UuhP33o9DOsepKQ5tSX8HbMnffThpibO6RZlmU
6m8ol3eP2lZ2HR1BXOxBwW7VY06ebTU7CibhKd5P7mXctpM1Hvr2HoMDibkyWqO83o7RCnmmYFgl
23pKUk31LKbmKV6AlOwv5fKEv85jR9fbe0HPsYyB7XpUAuys7nvZChdySB2qdy0Fwk5k3SwVb8Vi
KaHcLH4j/1NC+o8Q3wqb2CT7hgZjU+F/zpqlQrRDAFWOVomSJ7FGNtAeazSLgwWHHWqITo+ibBlZ
aplRGaVR2+xivU82YseJchq9Byph3th1g358TwXeWpoB7mdu36yuGyBOqi3ZPCrkg6WJ9WOvC6iD
1vu8wYTMiyrqA4JfkiUlcOA5MqDbfr6dHNjaZSnk209HEms9E3EbqaZs664NMHg+lRUP2OEOJEuf
XmjdoHiCp4TqmVG+wkkThLIR5wlyTbvEBGf+W5oU+HVGWXaQ+ojPQPvSwlWXuFUtLUa6/+VrCCzw
Hn4wvbox7sCjYp+z8H4xDef2yUWvAnwXU5hyqdr9eeGzuw7TMISAIhU4DG62yHroqzaXUHYA3ihL
OZc+10Byh6dB2cI7U7I2n2/w+FQopbDYNlW+dhbAjxCB5aWsEHJl0kk+YKnVGvrdGa8YttyumkmL
iGiWRAZWuSgitHfknh1d23LFKwZs0lyYkhhZ90QgXojZHl5AdQjr+KfomeXdTYI6MH6ermZmGMa8
br5d1Bb6BL8r99SqdNqbTMx9GKdPko1lJDbMJ+ZLbYPaaAG6jk1mQcub24g2Nl0MvKCqFcP+df+Q
4QxV7W0HBAp6voi2rvxjlB6PY+FiAxjNtD7TGrJpgtwLs5Gl73iTF0Y9Ow2ipb7SlY5P6fLc0oWZ
OuN8aAt68YBZGtziacPf130K2lu0L4v21XtFsAtvzH0NMX1Aq31eUnPuqkCHSTpN6UeO0OsDkpty
Trq9vlxeisIKtibxAEjh80u+ZVGmlFr2vTqKqwcW3IrTbY04IvDtKDjUwwkqpgURDA437saoS3oa
cOhuAHD2km6J+Zg67PXaINqyYhA4TZCr2MNNrkELJAhq7byHwmN6Meit4GyPzsOfej4K3Tj9KHwR
yTEngPxZVp2wv4Yqrp5sqopFroSGTotn5ZJT3lzOirVQH3Ey1OBMfd7WCvOE/1b2zdrK1rDgQO8R
bq+p5emnj0AmBKtX0CK5ZGSo+CeW+3XzGhQ2HvOdoTgvRVXs23qA10H6s96cUfUy8NJaAE+Yaez0
NKoJYXoZ184/AAb/VGsKIclKUADlOkgpnHV37WqNYhfmckx36+rqc8W3BhYpiMKUaPAAyY9qSBLJ
NDQldOBkrGztM78gGVcIyn095Oauimaxwc7QQo5ZhPmg7vb94u2pvKY6+UGXydqV/IxR2tjMkICV
8TwAtMA3n/6QrI499xbRFBXhH4c2xja00EP6f59bnNAgWzY+45fb+hrPejG4dKuYKQ7yYNTZG2uc
4fof+dKJ7DloXE4gO/Ec5XKj886HFhCeaLQYeZ0szLAXx4ObKRBuOV222VHMJ4p3/jqsDC+HIzoR
doM5FiD9f1OMPrCjdlGJjmlMMB8QsUXtXPwXbozoBqXCyn5r0eLqV/NcK6ylMmAdCypmbvDfNVJM
88hDsqu8JbmakBMmLtnUYl9JOl15rdhfdV7P26O7w1sHkvNYQuPIn88966MwOeaiZet3OUc+/1jb
RXIlzGjQHCA2sS4q+KNffvaOvr9ufZWVZrBu9S1AhZryx37y4U27nyF2TjP7rl4kVoUGSv8tkxxg
kIfR071Rc5trlRxeF86DLykUPYAJ4zGU3+2JD43+k7Pi+at0rEZGwQGE34Pw0KabZShO4GCu0XG7
GKe+SCJewmIvjKT14buEC8VHUx3ELF22vcqd0M2oTaGiKpHN2nok88UmbS3qBfHcg7H8aJktBVpA
cXBDQW51sGV27y9634xARUhX3nMjkIRPPxB+wsuUY9r7SEGHAcR9rGuMBFbqe0PVZOBbJKsx/TqR
s5vsAlEjluopdA1jUbaMFdPUOdYtr47DbSuOC3BLimLzcEgyTXqwLr+JH0C8VzdtlfwtbK4IHiQ3
QjUyvSgb9dUymdUvAT++jLgIq/e6Q44lAMVB2DgRXe92tbLurAQfWZ27WpsnoR2rHov0Nio32h1r
kmMKz1dC2Pom2RJ6+Q3+Z0ujBSxi6EJ/KlaNrBfuxN635j9fzF5Ci6Rj5IhwvNDjiAVrEUUH1yaB
rp2CmyrDeoPN/i9zXi6AZ0jA/9hSE4pRMmbzeGTbYCrFyXVTZxRTZLc/I4DtR78fe28m5jAEFQeT
bMuhKO+bv1CKrz1vN5a97/ZKTA8qPfbNDPmTs11ky326hPj6EJbfGJ+1s9MnTv/oCLwo5Nrfl3rw
OEUUK6LkFR7EY1BzdQPLy2tpZ5VZ8oIIIawTYnkql9o1vrwu+uJQ84CIJpq77BfhW4cAu2dftIPp
IGasqDgeKtdSB9KTg3klkw17ryUSpkg/5Fuhw9jeZ6jEDKDXGK5Rj7R2w0/zPLggXLjeI0hDD3+j
pYVwJXAxeWtufE6oo4J2J0P0V62FzsEop+WsVXO8XMKt240X9q5wJcX6GvjGVqUldoNG7K0MnWuY
h3u29i3/riCz4YUY54K6myIvRYN3tMg7Lp2fLSmPfA/LRGNF4Rc0oHYgJE2qSSdB/7+jNueDX+E1
3poNPY/4T+akjJWJkv/Z5Tw0o7iA5jM4VMRLtkrVYPpAe4GuWUTfA8nQMND6faeESsckVTYlRvA+
78mmyFO4l6Ya8ptfzkwrriKmFh5fWAeWk4uZoQaxoE9QXKsfWWUEKFqXS6Y21yt3KcWMnro9BG6F
FhpsfgvdtgMFPrcrePg9Y8RLNuzObtSC4I9wjYu1YVhw6dWu+5doV1DCGbXqfnepTUJf8XTK7i6g
hxV7mCqVwn2j3We1W+4Z/gUwxKcC31mX5owpu+VxpuaQIxzeTVuFZ2boH/iNVPL759bASRAGzpOu
1Q/8I3BTaouc7A6W/N986lc/K+8p9KBzIYESNSNDX2Gp7Fcp/FTn0PC7+OPILnTAtjKRtQ0K14rD
yAqEXC8FKoIPi0mpwTLbTtTl3Dt+Gn9E23hRHyehpC4jSLTs0+pDgNU6gvi3iKQW9y+L4EXm2NjZ
QFhtW4uhB0jjyKfm8OkrjO6Muubb+z1DmVZC7DUPyqY1CfBVElB4NWOrmmXsz1ZcqvwhT9Y55MBY
CxaB+L6sYkJjqfnJ024RXBGe3t3x9XJjqaplED8YMdGBIBivzTBU1LAzixvbqJ3KOW6OZ82Kylwj
pfD9lLdnK+/0zC1WBq5M3Qd1dmeWlkYKM1Pj6g8WWoUb1iBoqssXNGfqk32bBID1joFJHbHjByV2
1x7aZcU67/GELGG8sNDr8zfZCH0LMYM3+48efkFbWb/2GHbSHdWukqtAe6MFe8T6dlkK+VQXEWFV
nmhafUxVFG6au45JQGanwavbA71CmqUHNNSf3jNHKAI45ttfn3hQblLtBwK/9IAe8pY0YdWKDwAj
um5nmcSnr0P39Ps7LItoWwsmp6y3eFdprI/50qcbYJbVs1i6SwtY+RtFUahirub12tA9JqDsEUOP
j7+KI++F6kZLNbzNREFXUd+PhZGAb69O6q3+nwWR93x9UoOLuX95ELUavchJm8xYspX87zg3VUQi
NQ7vafR2Mz16ElAb6YMmG7FU8VmAH/7ZKEAcrd2y88gZUVG8RAdTdEp9mhNkYI09fXqHNsGjSxXm
6+d9EPjvY4Pxv/IdG/uez3NpLHgXJfifFfAe0GKrgUDkTlV2iWA1Zc3OYR4s3YrLWO5KB8Cr+LNy
iTjsIPWR+bJZv1hPk8hPICOcukcZBW9pyAX+kSakY59FhW3/aOrA09LFPotcVMr4gxVgx7ytQ2X6
y/uqQ95OvSuaTC7dkVCjvk70hzX918XYcL8FBtmIch3sK5JtExj98Dv7arucuYKOqI/Q01w1X4TF
Il2a5CbkJwfbhn25T7Zjzd+BZMbRL5d8zCRjQl8XsrAkb6Z+X8io+TdjugAmONOXkIMQyCWW+hbj
NZ+y+tB98+/wPViLh2MzLyVeX30HiQjJR0NaEXMJZjs13N6CgCRjxIlAV62YfUhF7G7vcHtc+HNO
5o1DTYlMblMrwVDdVgHDale8I9nGRD5JKyzdaa8+79AMo+fT8nIvrvIgsr85h5G6ssHbkq+97H3G
Zx7t31NqVXu1uj1JS3YYDQ6ctJYulL79fRDTSWMSoPvmpJCl+QMgGXIOE4dUZ8fofOb6Xf42GHKI
lj8Z8/1dv43SCP303KfC0Il7MW6X2XlRurypl6qZ9z+uoB68q9ce10Wzt+wx96nFI9tvzNae5DYk
hccP0l10+YqZ4m6mPUuEva9iXbpJX90iQUPLuyVe+EPKuYQXlFvE35ohIpk0Dc7cw+isWUAc/UE4
UeBnzbQ792eyiv02RFoz8Ow7z4TXC4Qpm46d7k7qn5KPlwvVYorHD6X7bK+esOTjeb5aM1s01xUg
0rcG98jnGDjUpLTkSNPk+E/b9EYZA6gD8q/kz4Q8+ParLyoLfMk9olZnnYwFYdVuP50vbb9/KV8u
1wl1HgCqqaBSCLkPGNnvDz+RfWSSCte40aAd/QXShfcZU84QB1YmcHdswBxDTWMWmGc6JpDb7VUX
ET60idYtQNSjKApGfExpyV07nIH3ufi3OHr11v3w5lvnhdHiB8GEVTJCw2n8wbnHpuO8SJsPvTnt
ESamQf6901ra9ZFscY46NdlF+VPeD3fb5b3p8BafVRvs87uyrKS4tFLgYPedJPaPHMRdceQZCCAe
1mcLqd6snU6vpd+/sklpu8fYfsXBVNn5r8iossSjrNV6QPJ1rTIE36Jp9UK41qlG8YQAnXOnioaf
arTyoHKtoEEh3j71l6sjAECxaNmsmkPMGSwYGua3ifSySo4zRV4SVsx8AjFJ00OErwm3Nhpu5V1o
OMHAN7eWTbBNR5c/Y0nM/Hz3LZ8S8g7CUeOYx5U8EfWtNiYesKDcgKfqvjBNionNBsqReP/uMjc5
JQCHjQxUm9kBfSzjt/DqGahmJhVBRZ1EkTpCzS9LzACYz8KgHbXCTW7QTeiuHt7ZhEyfzFLdqONP
dnGbrBsHc6QfVtPL8NZAMzGvqfTK0WBScypdvZMvHxdazBWXs+rZ2BSUmo+Clkl/VOl2oXeS5Vm8
Fn5cZLDnMp4OXAsBXDv2ERLbX4tstQft8m4X4kNVGpy27fkL8mdwYgnavLhqilY0KTllEWe7oWm8
2iKgPx5B33KJuNKjYyl1cRAOCLQc8U9wfQugxPqaRpV75IYbwq9stYttZV4XBO8jhysIh73moUhL
KJ1mscpoq7cE0JMrjWfYS//VwhdezUfEXGKP5Spk+Q0s0vWnsfgGJejXKbvj6iPB4fldENhW88WP
oP3jJZV3E2RIcAPQuZhvQT5FXAQUyEYeqdEgAyuBKO85BxKl1ByzJUzNigEBJQCsQzK6nOFJihXP
hxbRJlIbXLkZ4BOB0uCBZnXolT6EWMCVcUpz+xWtxxbr7fSNHPkC5w7SaUjIXt4to0N4uVjMAaqX
GzajiRSonScCsKlep1e0G8jk7L5GLpIIfAA+ytPNj7nMDinCp24igf1dgFP1NmoYGC89a5bS+iTK
jx/c0ABTjH5pAf4ks7zJAKyBfCfsVvOVnZC4T5MZmHkf/ntQPfSGCjo5tlSQl43qohj1nGXy7Zap
sT4gR86vdr/oz59g9F51xk78rRJ5Y6FUhcLEWx0nBMBj7V76t68bwj6X7p7ZJS9WcG/ZPl+xP0UO
RjuIgdF1vLDG9LU2NIw6ULIJQs+FifuMTZyL7Gj0QhayyRcwEhDpYPOCqaKM95XC0maSS15rHagf
IWBqHgYLvzpApzWwf4zj9Q8+eEuW6AkNkCXvId9rDJ+lHputIBFN+orUlvWy/3pk4E0+n4hLgBES
td0vBuLzI67G+nYXJS4P8Ph4NWJ/Ccuji8gegBN34z7jex0+onuNYU/y9JZZMLxK8H7mLXHpJ4DV
PrnPsjUuSDpDzFmCAGZc1XPJG1jgFr63j3uPUDJfJ0WhaxenVMPJcgHMMOzAWd0A7kHRtPSDwk0U
jAMoyA7c5p0MgAyRyt6SiWaJ1FciVTNwklh82hr2jVml+QleTWF2mSLWiTiaE8pzTonJafwyS+uf
L9TxiGRVMF0QWtGBKjVrunJuIA+aI49RSFZMMtiY2ywJ5WExSy5taEtySmPY6rrYiXf9l0gP+Clw
e/9B8CX03PYsUB1H2pqOThhwqdp/bN0lkPG7KHf2TpLBsuLRT0wKawd7AivweBq1flIZd4iV1aOk
+uw90GwV0Do+znocbimwzRQbv/WCgSPW19zpZjAsPM/f3mXiuqm2jgl1mesFmS4Gg5sjVeFUtXBQ
4GqNLqN0HJxr/2rxtSrjbZpC/M52VtDiJPfWP8SyBxPf3ETVDnwwVR4Fi81XdSvVzsoNKjx3umOP
U9rKZ2DY+NUKSLKpEGagv6VbD2vhZeotu+CrMu99UHChksJ/zprpCjab71DL1Y7++8HA7Upxtwjw
kS+YvTDm17iHj4y0Zjq7fE3kgvr5fnDFBl55eRQ92YuJACIn4b8Ide5qQFKOOho4Ubn6AIdEpGwQ
GxlXMYZX13E0YRicx1q7sygnDvr4PtCYRFXuUSX8SMoGHX4X5hYMH6y3KvW6hqVZ5GjX5t3PBIml
rBBesZHLuA4pL+toGeLfU/vAO6mm3EYiHLzXfPCpEfhJmQnbv8yf2NJHlHd+9KleaIKdhru/JJh7
wI/EHIXqTAIhqEYEjMUAsfy+gvHfuKCTmuLH5Z6ruIfyI2k0nZeCVgYaZUwNT26pX4se7PW+iN6i
q2jIf5vtk9eQvt1kkpe3R1NxGFtX5ittuerlQqVgiy7LDgj4YNGS4L3tVLKA5pDd+gVPgNbHQ6nk
N0MDlcWD3l2lvQs5ZvFbhIPs2BN5b6FLquZXBK+mY7W+xl3Cpe/6V7XIVjk0bC2FqLFZfLgNgl83
A2Awswc6lGP+G5MGZOJStM9LmG+44gYJjmRBf7KtRxigmAGjBzO+b3BmrgJXRRcy7fzoW/9hoXcj
Tgu12r4CHBpCk2BApZhLcSOscddL8aHT9V1qwFH5nGQRb9SyhONmpzZcKBXASoRCtgO9xTe8WiOH
UgsGzgX354OQPjCPiIYYTJ/LtbwnCZ/VF7C80qwrgwsszmQlqLFiSoYOp3rF2nd87T7HCxdFAe2x
SMZiPX5idEuJ7rV+drr7bMtK6mi2tolD/FBFAvXtjgsD99AD3U5GNoUtc1JIJ+hkQSPIRJV9U8fQ
ZZ86rfS5Pi6WnYq+TBzGGH2E4Srd4s29VbyFPF0Mu8ehOrOMapS7D4nDch/prZK2Sw45Y6klIAFT
GVYMuWnEQ1S5vmbL38/aKs0zZ29O5iusJp2Y+Ge5bFqaqIWdSTl2wKLeKMF+X9oYkj9dH4OEscmy
D4ttdaGZ0p6dz2yzx4BrkG/egFmCn3mdV8O/4UYVybsi0apqmBttXK4SNirJrO6blCKv+mL60cSW
cZk+S1rg67Z34MT31wYAeTRbkI3gMobaz6G6S2wQVAHgtBVRHKayi/JRTfebL10F+s1iZmT0TX3/
m8XhWLQSISgLNpse/dIE5iW6pAaMTfbA4wxrLaHHIpU6yFAooxviAMerqwxO7d9MRG1V9so0F28q
EWmAcIjB8EBZCR38zP0PqXQXfWU6gtzlwvn7Qt7kyZd+G4If3Bc/Wv02dq2XKwZJqI/LcN+B1TQD
eIHh3VQ6H5gYckDnmwLMir0uVVFFrfxh7cR45HIFEhuP8Q6i8fUItIuW+Kd6VSie4GMDFIuVpu/X
jvtCGlCDcDnosmkKylQ4C9i7LY1InmriwKsUiUUxBGsA60rUmGcNEFFJ4JPB/9mdvImV1LmKt+Bj
CrUUzw+qqKmGELKmq2h5kiSgyQQFOUi2jljAYRAfVaDHesrDPRrcygzpA9Z5ExOXOgb0/MszkHwc
5XliXHWgSzWDscp+mRJlAGUUNEMFHU9NzWsNYkIA+zGjly7FNjzCYusrb1Ud8EBh3HJhkpQ37f+p
5nZQHFEMbtYjeoB5ATHaVry+ykx7EX2WsMuJiiKCi7Br7I67G5Nr1khzRoe1/eJqctwQKWw66Sm8
BOq8oX4kQtyyoI8J5gDHCPj1K2mVWsaaxd0HHR4F4A5yB0cB1CAckIZhxVaiOB10kWh4jAGMfrbS
ZBwSDtHpWY9a2jPrwrnnk5RWojyWf9Au5XLdeau39L+2exfxe0EflaK5zoqMVj8iqzf8LESak6xW
YmwEy/GD60NzjFbPJSTNRw1pOORqI3gXF7bSzk/GS6CqyXP8iBZELdgxZx8sMd1wUtWIryt0QEQX
V74DakDUEneK4m0i/iKA4KCYVVZa88xhIKduZW+ijAUNcTCVwkNIGuyy27SOB+SU62i+lPrDKqWC
WbzU0M5GHTcBgoLfg+vy3PQQ0DqWPnwrVRi5p7u9PzMbu/ujYGoNPCx4STOg0166GFrspSHbsfaU
C6NeX+Kv3uQwRgmtRe50d32e0bw5wlJ3NnP8SKxp/bH7fEYY1yeW0zVq/G06u8GG5NYJBngMgwks
7yO1TxWqwTJZT4jZCzFr0XUi68yf8dpLLF0v1BB2pWiPzzgLumuzMYKJaJxetFeFXU87z85txTZg
95gr1Mz4p9d2u9unAMTNvsvKBIrLOgl312vIsl8ukCF7WOT4viJ0hp7qnG/E3g9u1oNFY32gUUSb
uhIDzeFy/C1F6gaeRCYiYLE5pqKTMpVQRDuhJXKv/FjTMXdVzxm3WBhVsJCdoegkrOjB/YhOPJEQ
UqSHPiSSEBmwv4iGq6h2P7UTKCcf/RNc3mXweWcOFjE6TFJSK2gWmBPDPaxAewFq0/4cYxY+3J5W
I6lKh1t7QaBoLd9xf/VSxQr/O7uKyQe4D2uqSjTR37lnXVRMCKAx6cftClXtkpNLQOabOI6WHA7p
0Ay/og0Oy0oaRa3e5hG3BN/9hWCq26vXx8rQamu0qpxMZ53l7oezFQgyYjFZ9u43jteGLmd4rS0v
s2YQObv5sg7TTuhVxHhmnhGGMdjwtLwPPzlF/l5G41FoPVuclx7KJch6zmtQiPwCDHs0tGuG2XMb
PXcmOITrCMPkySVwtsuyk0xovXQY+BcGPD52MkA0JCxT2BQDLv4trx+uocfpNXoDHleY3NLIIweZ
FkEPkc7cxmt+Vt0GOzyJNbHEf7ofI423Ek/KZ7FzGAHBzClAG5bdVSrCjfPrmll3tlu87humRUK1
npm3GPMjEAr3Lnwfco+URgY9qyMmQoBXldtsZsA9/AFJ0QjfrsxuKK+xE+mBWM5A6XyrR/Y7Jqit
XNXalLf1vjHdgNqTr/kcndMOBgvoKTeIxscERo8N8vdkG8HDfJNJnS5aXIhb9wTeDm7MjMtgwlH7
HD0UBUml6MPuwiS0ZnRJjEIBHUmVRPlDWL9JxwIlqUmmEKim3lH5OziIogezurq3LXK7lZaxPeGb
STU2ar0vMtGoV3KALGBSG51DzjFbxYjZBR1DDgkviuR8dOLxfnNIBbEfOT+ohKSvBTXh29v5ifzl
T1Y3w8/HrN50CpZqaynjP5g2dBhQsisa1bzsHxPxvUWEYh1zFWJDcMAvf9UZB0escJOdK3k8f2WT
ESJvEHeqb9fAylToc5hlMR7HgR0iOgxx9BFr5quVTTnduWfIZlU2CqqCZRfExaRzZSgqmnaSBFjO
uq0V/03XclXKcQsKrffw5+MHalFh/mf/lG1lMYCDScbrZJNo5EAet3nKt2jwqVhRFf2fKWuEe3GE
SxI5/iKWu55dkjAocVtXgHkvpS/sGqi9UdB8XOp4DGJhdSyPftZU/8zy70g9mI8yFiYoDcQZl4/E
JPCmW/+w8nmHIEKBD1alpG4ODAgNQJ/uwVuU6XSHTNWv6ZxKgLtkqiuMIoVCjohw5yEHt1S7lemP
6OIwobeGTI/mTimJL0o+B0SvZuBP9GX3gUsj0A26mN+Mvhb5v7PO+519ow6I4W4Hyh7JOwBu5N0/
1GLC6ZI//UEq+7qHOILBH1iCmFGQTZRlgSkzLjsaikSWH2M5B1YDBhGbztcu7doctSLgI+oLsUs9
VvkD1YtJfbd29481lMYDBqbQGNsGKbkaXbqRWK42AaHd62PDk8HFN19jMVqmjdHsnKQPzE1dFkIc
1t2acT42gq80PQ5uzOSKClf/uxOgt5cJzUVx713nugsWb+upcJ6TjFIe19tMEOTC3WEsa8yLj39V
hmZ7e00QDZDTZEXXLK6xe4C+2aZdc5npdQeqvw4E7a6EMahtCKTlrsDYhmlYly8sLq4iAUwG9QK8
rni0gPtvAIbpJpHayoQA3HHwHNLj3VE+VR4RBv2g5TZ4YAGZ+hTAdEgDAj8LJ6DWgq8+ZYIpi0mO
nbM43wx3uyYLfCOe3Cr0S3XHypTGTrDBlCsxNIBAu2Cq++ByADEXQ5+pnolGa+0K2i9eJwUV3qxf
HUnOZ7+WXQ3R3EOf8XycBhcVvEb6fr8kzoXxbnJMxWSdml0fferBo8PYS525z6Pnoxyxkpru30Xy
aOlB+1sS21WU/k6fSUeN5VdkjvrQcQ29WqXLldiTx+Cetm3DDdTKEXSi7t5mOzyXmk5rmOaO8SHr
6tMRQASgL98UayQ7k8sTzsxrFtJqDRZE+/duFLBOmP856qw9B2DGFJPLIf5ZwYo7x8KFZDIRJBKg
00bO+ES2clptlNxfqoJaV2ndxbVGL80WnYh37E0/PdcqXdYWmIaXd5K/p16F0Db8APfeWxLMArp4
KAkGcXtGCpXQy7uy0aeeKg+V1lPGrKrmuVHyWLnkr2UV4SReW0+llnA3qq/WkKE3aC25iiMVJhui
YKVMeTAts8eeNUBrNHBpstgRQQBo6OKo2BLRePJZ5/asvgT2NwND4zfgqydDfq5WypviX8gRvkfU
9sobmsMfxuFEDbZR+viCt/3laCcFp9RPy0Mj71AFe9opAhOc+h5LxTNDKbThTEg2aresIRvU1a0j
2R2CzPAg6Sb9cQqeKV/xYxmNouMvy62V5kaM/govmPDj3r6Q8T+Kuh3hIBLO7k6PQEivHcq6tHLJ
uTn+dN3DgHZq2jHa2bgl8mJPN+jhYZT5smfY3T2ZXLCf11E5Mtx4WbX72+ES3ZdakpsGnQU9CEVM
PhZos29XOKrWReaksS015Kn31BHbp+Ab95b4HqHw1Y7hJQZgiQfGP/41EZ6GM8EhA7YNLpYAZ6NK
22GydYVzv2NnGW0Dp4R5wI53q8Wi73b/rl3t25HNLjvkQRNPJGI8Vypv7NC2VBcKi5UmxrVhJM1c
YmNpe72qHpmWKGAU8iquUOVumaq7TonurXMDBtviF5qU6Fl+7v3/ltbx2htFqx7sh+Ok8CWkjHMB
Yis5QegW3yB0HPhJ2R8gB0NIWOqpGg0EAsi4I6s7AXesCy/gnmQlHN47uJyGOe6VMjcA4YuTTn8C
m9ILMnjX8xCpPvaM5hY6pAfUBlZ63sKFbpqRyJ8o+GDe5EKPu3qRitlErobNru1QWxZSDZnJI0Kd
jFK2NGdAYUFhwHSjmYYukNSFc8MegwN7Kj9gMpZOdDnnn68VXyt5h4fzcVqRuL6sZg9yflDz7zhR
Ih6Ys7byzDwlzBSTM9MJbiMU5VXy8hB+TRaKuC1mY3qyQyhs+wG29PqAg+r9pEvEuVXD1Ct4V0u7
r38F3eCgemZgByfgVyoS30EpAqnF+LWPCACStjcDvbnrCioZSOsxJ1OcIiJlhoMdYEmzkbSLG3i3
R5MMCT0fQsV3ROHZjOz7Vpuoqv+0PWA67aNN/tiN2aIcAfcbZ2iwZjEDlyk0kbWLbw2Pg+i8FbOY
C0ne9Z4DheBqE+gQ2Qk9zK7IjbvuKnnLlMpXL/KOsjJ6RdorWXqPsC2oG4vwzXEpxTeRW0sCyO5n
0bzu8n/ZQjmOkxs+2i5P04gl7z7xE5Yve4JVraW9nbA8LeGyDc0aCua4NGVhBwr3jPHrSnfe/D0s
S+kRTYZOdB23TK7V6+m3dAB66LqKFbR/qJCLIjKzToZ/wQCeLKsMizoBAWoTmNXspsyEhohRNSX+
3Nv2WKnfzT8hHczZd7RDi970IRPK5FVCsUqFYrk+8kM2CUyZQYyJM8FEF9Wa55i2XAeeTZd7aSZF
3nzrolWgBdLeRxLdQ6+8kApeTRX50AnFGut9cb9kf42AvAkBdU15RMRVEG4XXw24KVLTig81yU3E
IwunCfahiAkr86EFQPtrRW+6+7sFn2lr7g+DaJ9ECugLtXoQSpFsfA8Aws5O7CPb+Fq9du+adkkh
ONmgkZQDSPOhND7Vakk/vkhoAg0jvuQatuxslGyScsFZIzOybigO7v+yIczs6ycP5qF2eDeAywu8
+4kqEGS/Exn1QS4YEAVcvrs8e7HevVM2sha9ckrUFX1hYz9NmdyL3mINSd2WqOD2vko0Oi44Lg5Q
aWYr/x9gStyyrVlo1m3qa388VdZ4nNg6oe1ZsipwG4j297bPWip0wy03+tw7vUttgSsUhkja+u5m
SOpATKY4ENJuFG4DRGNzI7RQrJyODxkJ4uicCNbLNQJSRn0jHY8whEsZdkUgoAgA86NHtw5bsw+m
syw/Tk5gHwn7UqOpUWqCJ1bA8pBIFEVhvweVHUvN4smwybp8pGG5heZW9osJvMIQn/mfUWHlQUCz
ETvU73uwclVzFOA9FHSgrmt0ojmt3myQ7uOcvIxoUMEaYN1r0ifscNh76hx/3YpyfS4AOb4IeNSi
gKBcjHeiC5uwmk2ExgNc/R1glZaPoyXrYW88Hz/UiqyNgHS2f56+5feB2cwZe5VUsH0v4l2FTfEc
wdHlOXnJKK3Fv9xv3869mxq6c85lSUubXiZdTDaXhJQ3OYLsN8g48quF9IX4V18HOfzpKpClFuEZ
aXnWpuLthxnZZsspUBs/+LkQstDxFXNLEiUMTM1z4wVcx76lgLjM2c1dNrfLc/5HL06RseK3nHGs
7D3Xt616G9hiJ1gD7j2U+J9+RBzKYf/V56ZUtRmTxziVzlm3MhEDnMgGAJkYv50xNI2U/yQcHF/A
EzLbNUtknwNclyYu5qiL7pP8arD1wGTAqr4agoJufgxM1t8UqCyYU4Ya6bG1saw4Qidvbu2yN6qK
t8QJQC95wxPOBS64PhV7CSeAWImZ1pAq9zGBcB7cW7wgWud6tz6OFMCB+rCz5FRM5ZtYOrEr8/ZI
hKktpLKIYdWrTqt46/z33vbpTc0D9MV/wugOQbQVIIOKFXSaoSyMgklDcYf79/rMQAN3RzGXWG9i
4nFqjPS1ojiOGJ9jkAjhy9vNwt/lzk9YH2ZHxbobekfWsbsw3OqCrnMrDSfIttBvQPiynS+TS4aR
qpkKXDcbSIml1g+3P+hgA87Z1CfRMaczbJdHnYVBZpdS5f/XRiR6FLmBbZdlZoWjxGAv7m4ZxNo5
6VrizIykjhpfdqZl0vzudd2YOZiwghf+M7GVOSdZAGGyn0U2/vHEBNG+zm/fOWVScEZItHJx3yZ6
cmILV1TDetgEiDwTyGAwQB0VMJ16BRxvhVv+hYDwuie0CfPHku8jQJhKDf/shByYjfcpjZyDqpLp
dzeWtEXnDo1vEfo7xQN08aZxSmyPel7w5Y9U7jWq5NxznwrTyMhvS8wbuIz1ULCPgI7e9iNDymKN
28S2nOV7+yEn5PM2pxF5xmagOhQdqfz0dI6HGBY1UqxqC01tV4zkL+08o0A8y6ZE1qjin/X08S4z
LPBznI9VlxjPb7vtqBztdz0+u2OvaxzHxSoq+Fgt9u3zw1W6eVpwbyqAgz3AFQHtcCGe61HzAy7/
xmA2So70Ji2+IbpTYRkSiLFUQJOtQIZXx7y2z/q47Q+n23l4OqODOOR1hdKEMWH5p4B6isUjVKY1
docLIlNuC8oWCnEXqiSNCZ7v9I2felN97mlMkZhJNLvV48bfWU81CPt2eStF3VNsapSGdH+E5Lkc
a2+w1IaURYWCNZAjsevzF2Ync5CBH/tX5sE03GtG7ME8MJBxCtRiHmY3Tfc5ftcJdvzD/FWR0RSk
w2SMcXmzPI0M9x221VyIFWy9RDTLTvYsy4Hc2kfrYdQ9LOMqZuz5oCW6HncGo6DFUtnAIG7C9edG
ZkPVs9xV7kCVWlXKKvfUsyhzNLTq60cEwe99DNdgdx75HasiW9lMwJ90gbTpgm6kPxbrvjvFunRy
ff0JtcSRtVqVW9QkkglfiqDFG5V1oDjqXX9D7CpLWFo3mBhA0lPac5AvlRVHL0/5vWwcGZ951aof
iANmbsIOlmWsitnJJMvfVsr+SzBn/oHLpj5mFUO7ELRK/KpEXnay9F7GNESoYD5eYY6keIg8LExb
rGrYP2coySUs4B1+ZCkTEV7YxvGrTdT4hoZQhdGXvaY7voLOwS6yBiJxkf02jXh1RXsPrpIY0YNX
TNEOs9nrLW0fgULBSCemtb0UZoPcal9nxGxc3UPuIDslPza4obd36NY0s3YZnYkAlVaD3dNh0Qi1
DDbHloHXrg8Gm3r6VfldyQAUQYJYYhweQOoVhD/JmzPZj3dBfWYcC69VEsCsQiyfCaVhuGqKskXO
q1erT8h0ukQkbJbMt4J/xlRK1rkHphiP4IY+w5VnupP/ez2EMQtMUlj4WOABOATBRNTSF7a7+E14
n9QESoxfB25yf+fJ8DtcjgvZ1ZeAUcDXtROdcfE4KBduQ9A6h9cIkVkQggnGLQlzKlbXSyt/VmH6
fRRuFI9KFVq0lXt3WOJ0fX34vEGifmfoSeorkSnRiUyoKyGDdA4N4Ds9nWgQrtvb1ec1xntj0lsf
5cWAa9F8Qq8mkXgQLnmWfP6ul2Db1db7YyfD+4A9idJ+BKZOYNt0zNDfBkGmBSj69bvoUqh4YdGr
rg+gPk1eD5FwK/Y4cR04L64DzoDC5NXy9oSdXzNweRidn55ctG5FDch7DPXwrF9z8nwjty/5oeq0
xdfW+10Si9Wfih9Ld7IYlEGvYFee9XHAaGyDn0vfMjFmDhkFBKrsggUxljybEmwZiETfsFRyY4L2
qVRnaz0Vyw+vnLznm1b6fyHWhd7TNbJZLzvh1OwdBhmNYLdaEMMzLOcYdF9kMADjK+gQQeM9nne4
Yl+N4YwWSSUHceJDH6PAqxicq0Xk6d0uMvlDPyoj7Je3VSnFIICrmecmqFnfcDMPajRPfcaKeSDq
WSScPmqGbvw4EcHOerX94ZChKdSimdDnsGDDOGOQHnBwEy5KRNAOSA9GKQ3RwB34i3yuahtedk6G
TrRkbmca4gESpi+kM8371Gc4V4kk2tWbhJTIYEHOQg88G29Z/iOp+10asQEm7NiYWPet3q4DnMPL
i6eMGLnJvwzDNfqDEGzJidtlaNI4KogBo1u0VcsFlBeTyX4F8CYbPTsKA6LhGVKfzZFCOm0Gf7oh
EgY0/N05gZ8VhCo/xkct7e773QESYt6rl4nLZVEHrSHc6vvInO7Uw6Byt9NjdOI34/8I5maK2mFp
S8WiWNYcnkkGmkBJklTu1QKig11nt4IiGQoCvPaftKXrs5O8TC6EdXQN9CD3eHuquBPi8kVKP3vj
ugJQFuZcm65pX4m0YORwJ7n3+ZuWx22ODtTyGSnT3Y0i9XCSYmPxqAsfI52LQvgeGakQagdsmtJj
NBuy20tzhf8YUK4kLbNWLAqbKPnWEONBZsOIKGz5eReDv7a6Ge4decxrBf9EojwpgQscxasTz0yl
QhviJwnCmcu5/DjTXQ1hGAb9bLwSzhhpGxks3Bpcy86R6zuXfbTicAXeR1ga3Uz/3FZHMbvzNCiU
JU1Ii6QH8ABPTAQf9iLei9AZDw03kEFpkXiywahYs5JwHDi9TwJ4BmlzWwUsh3sg1TDISn/nPUqX
hprvOe4nCtD/qWSwsgBPExNdhU1ia2UcZzZ3+/aLMmtWx3O4lwLr1WR+ze4oASUjKnQREPwqj/+5
Fv5J6mDxyz+YC1CDppcOLrdzBMmujPwM2TOqeea/TngLTW55ALFNaqgnKgl3SpvB5M/LC1EhSKky
AUf0BgRMrA3BGAZMDlqztdDgGa/LFYHcSFfGgYGFJ5Np0zEoLA/fc1dzUW4F89roRYE8hyXYHXKh
cnY7tAMItqNXp/SmU3YkvWpbhHTME6wtGi2N7ww3feiyxrXCVJFcRlazocc98wyHwmGU3JQ2SR6n
RXj35+2KXdp1oRjHzvcp+hIMzz0hocSeFG3IAHuIAmZoVmgajlW9eQ1N0kJafeb8p6p3OxEo1iET
ASa/zB8tdL35J1Mzm9atGdKkXkKWelK3UhsZVZOJ8ToXCurRqD9txBnbvei9f3Ee/4ttMGRvM3Bz
iv9AuRSkwTIG3/0N1fwDna0x8Khr+aHuGEczvXlkguiK2LTg2uxEvqx912A1g4nD2e2pdPV1OYbI
pYCPiiw4o80F3SJffuGFsYJRxw9Ufnp6VxwjpOGKe6DNMs0+XYd76nCSxw3OH00mE/SpbfJBCvVa
4sZ/BbTp+zVQpdjpSA+F9QfHAPwIO3MGcX3x43qj770VhIVWEU11PSvgOcXKLz//1DNX/bC200//
lZB/5Zcew9ygBjZNTJVyLr5CyIx2kTabKfVp98qUeIY3as730bt9y3O7b/qp/guAHstZUtbfNEQ2
kUnHW/rIn4QTh0jSQILP89PV7/SSKG1XNrAiNxbkpyjB44X1bpSxfbh+iGfqA1OldkJl7MPfwQF4
rd+PBissMg4ohS8fPpdzsWpm+oc6/o4GnTS4gqMTiFS80Ntu7LG9pUF/+BZ2XYDHDYRHUvl8EalO
rKeG5ljZUPyDCxGECRemNPyFiPkd9IvvzHCngXurdMLfDfC07XlBIXkhw+AOIbaO55+3SlS1/hRP
blsACUR3nWBOfgFzkVbFm8+nQcaMAXuRSHwMVmAicuFTAwC7qP5+mBJqHKNKa7p/fuZo8Zu8Syc1
/YYqfOnCQXSCI9j9A+whpkTOneKOn24lfdXiko90txSVLXDfupoIVar0KYbTI+e8bDgAIt02ST08
Lr3bHSzNn0kkql3eRijHQwTcc8br2jKA/9PJvc5/TOM01LW5ZADdb12vVBa1N7f9FG2ImpT3Qmzl
tl5ZCCSLHI8JJ9BF5+0N4/1l7cT0E4US0cY7MWuWs9IQRqyq7cQ0THjJx5AyAhZkz/KuTJObW6Y1
yee9AL94EwKLDpHWwfITjnBYAjOZUnl+AFSJJSQ2ZPaOgwa4yJIzJ3NOwPiMi81B4URhwEQR3d3g
8zwn3Y0EDbdDtVSEWTDBNyqFDBPUcW/iD5iKMt49iA4DQ9VonNcnl3FN89kr8lCb0VCCTjdaSdNJ
eJm8oieC4GFATv+z4Fp/rW7icxx40nNAxNMeEcmez8LV9Fi3o05PIaEUUl2gwnNCQfsal9C0BQyG
5rbRz08Ae3S6IQkhInAWEJVUZrxkzQqiSlh0POg7HapiA1m0Srv7EY1LIq5aEpySvXgWnrnTrGro
3mfW8UHQWzMnQMzHyrvCODhtMwszSzsl2FhIRuYiRuKQOOwYDH7BY7nVf3YAK1o7c/W3666b4qEA
H9YcEXKJHWyqTtllioruxjL/UG3IZyZru/5tRlr2Z3MjYLSBBCnRIgHNW9i+jjdnPW4Koi3F0o/E
JfkI391dGQU0IvmiwIFlMktkj884gGT0GtuWu0CiPb5b06tTGrcrTMtVcskarw66Y1e9hv+luSeW
0zPXveazZkqEC2sh+JC1HGhHFtrJQD/CQy5KRcCPrFQuWsBpIZv1N1/cWeG03/dXGkuUlQJk1KCp
I19RPlz24EvgMVbWqh3rBpu9oGOWvAnZ0dWRxPwuekhFSfRzIFGSyYS2eHd6Z9rXvGk2/V0jfiyG
VL5zIvtRJgzuGRQgd4SrjTTAb/r2w/bJ6s3/owZUKCXRVtbu1KdC1jbhZkaMuPyV5vdy9WSP54mq
L5ZkhfZ9OFL54k2b34n4u9ftVCzC6WxeZXmDmqKVIwGKz43sdjdV3+E9paxKuys6y++2pzBjXhTC
vXfsEpjI986yJGmN8SsN46a/zDAknGxxHSgzLV0mthXsOzdJvrnjlJT1DdCyoM0QbxU1q+wlax5I
gzWP/Fwea+M7C/FBo9bpuN7XOfGnxUefMDZ+Y37TTN7TmQQt9ttJzK92MEIxEId3hECVhrS2CCvW
I/GgIV1Uk5QPnKjFIwMsoa0BZDf+CZ7jHY9glZdty+Fe1YAzHoNon11X2cRnZNJNXCdJSCB0u0ox
y96dY7y1IOuCGFxob/X5+mYREfwzDvYJmEyAjlMXtfa7PFQ2Nl5Q3DyJmVdwvHyAjLneXFlJ/XVP
gvyDvGtGxTywHCSFQk9h9a229akNmPmBQ41L1ldYwHnK5aA9rm96TpESZUwHlspYz6Lac3FioMAz
lTPR7npuoTtAnW/lqusNnIy2NUNL+ib2WDu5jvt08neEGTIiCgO/7NsrH5x+uz9MxdJNd3HYXTOQ
eCAQeBZoqj0hWPd/Y0lP7cZloz10+FZNvBfo0gmZIYsSSqnE7BBZbnjMNwN6tnaH+T8ev+bd7S61
loNEqUq71Hz+dyaUn5u4KneNwyArvPEgSOWjcSnf69SxvFr7rPGsTI1vBC0p+v6cE528S7XHOdIa
wqowh+4Uc55+9jYHaI+vtu97s6phbAWPEZRLOQygH7iuz3I/rR21MgoLTygQ/yLDcdm6Eyp4Fr9M
ZaEBMH+QhC5Y+iXf8pQh92MIfCszet4hOk7xuUq5nMkfn8mahPXoTnRjY331w9D01KD40ZCkmv0I
CACsdoEdLLcbLC4QNpIUFcVcla2bnmNrmvkhaTAB/xwkvb/04KJpJBqCriWprCRPEq3aEVOoCtFB
KTk0CRCWwqmrkuP0bD9FHsUWTzN4j6DZlBPDQ/O4oFw7tqbnYA5fYYwUn4iNhOHK4AWZXHPYG0LL
g5AC2bIk2mSvyYNWNj1YVIkg1UdqCc1XxbhbUYVUc5AjFWjqBHMDxqwbWxt5BQbKUd8gqoh8su/w
u1KD8aF9NoZyshELe1jmbmWMZOx2LmNEm5kKEge0ez1XLVWKu+/3lIu8omMTb/hSW36XWOOqVell
mpHmOLyW9sq6VVAF0koKMd45g1YnAdonwtrF0+qHrQxZmdVK96Bf22KJVMMrjoeayksrrZawGlQp
pt3l3WDTj6xvjaoUfXGYoJuRFhDnSCwg4ac1bHgR+YgIiN7SqTfmFv82QfGrtkWs7wdban5Msfcs
tO1Wlxl6K8yB4Moiuf9ZkQKMUnjvCY1I6Uc5HfDchg+www1PjqF7u+HPKSD4r1qHIt7lcxjYCIDv
ro3DR1SQLbC+a0RUMw2sMTiz1zGIGg7l5cCXk/thv6gUplSHWWScX44t4zQ3fJZVD10t/ujakQPK
C3ZtehufV822i8V1AWgABnUf72XOoY8XIw2S75iKpeX8FfH+NQJlfMzDm/pc0ve8jBeCYR+oE3b8
B41uN9oLIsdOAb6R+EEVF/3d49Y3pYt5meCW/HJQUbQIHpqrxRyI8KZatmBwbbqvIDmoOaOkabYK
YB4bVxA2rIWIaFARcjOkhOHWoQT9jmxlRJM/XMYakwWmiRIGClBgrfah+uncX9oGLYXu2vNFp1qG
++zjEsjZQQ1lzpgBYYoI/RBMlUKF3sV33XUsVji7NbZ6/+x8oo8F8gdsXF3u7dnIb4rnX/9/p2qu
0leBkbGR83DtXTXTKW5aJr2S8YxWTJHA02zoLYOMDpiUBfbUJ3mEtPVJCQvMkb2z2WMuPovYfRMQ
UYCcccJ3028/7UZZcT3BFAWvGV26bYxCfy0eFqO1O/8Tu2g6J4jwPVuQdMJjVVmjRPjdGNOQhUtp
Sun0JLFFcDNl8IDwK67Gv9ViNp464iIecTKY1990lhuN1mGxPOeMuejRtQIf+J7uTwMzWq070JmW
7vShQCM0Jy5uKMceBrITD1vP0nbpDXPYv2b+S4qDUYYHfpyZiRCmqFwR5yjf5y6KvgQ/p0xCcM5a
KN67EM3Qz99x7wJG/ZpEUngX8K78T6qc3Wiae8nwC82sgslq5f+jNa6y2+uX1Vbsj1IyV+9vrA7b
YArjO5ctWZcUs6pe1rbYGCX1pGkKcKE/MDGiOFZtGyaDWGpx5sKKaXoWyNrg9ANV3ofo3NbbI0Bq
CWEAuxrpS/fMjekydyLObo/3HAbrdcmCu22wghn59DxPcUvqBvBieXhvRUv0AxvnFk2KOzhixKzR
hHrIigyYDoJvm0PU5YNqUfav7JqvkJlZfrjRBdTz79Z7ZrOcRTcKz9U+KiXc2F4cOw0Ft2TCUiI/
zQJ9Ik83STxrNyT2x0WgKyahC51NTbBwkiuvWARiz0Edy3rZDmhYBb67ynj/yxHPgYYFiwDOvVgY
cTOFBAWLqYRDktTMQ6Efi4OzBpp96PtyKPVi8/y88Oi5M14f63G6x/z41KdDmRgBB1gJ2UIMIJoP
fYYD7TKqZVVJ4OEzJ0W4TzJUx/gWXKx5JNNfZvOFiTqcU3K2aX6ygWOm+wkdGkyOcWdvbQxEQRwW
eZSdjelrM9qQmTI8fCsVT0aieYJe5ekWrZvP+Lai0Wz7RiripqE7V68DjtxOkJMsiWrQ4L7+UFel
c2OhZh+RbLExWVZAcpAvA6R/uONMDl7DMREOJ+SgZMSigIuZBm2CBTVsJiR7eFCy4TcbAFgj95KM
lNzDrCt2C0jsYkZWEnIGGupH3jmtq1hX5OesyhXTLRJAO3060cvSpWzId1tb4iNm+OagCkqMfiIW
5zQOZYWdZBljMsHco8KGxpozI+OCJeHPrhsial+HjbPrGyzszVnauD1Uwm9uWF/5dgHDRdUHIVGn
/RcN7zUe1Ry49NzLouXdSzRQqC1MaTnhgqvEJI2KUdHW2EIJXVwXYb/91OHbc2IpB2utoH+tuqm7
DEKiul9haO87ZV5FONoR4Cksje1pYWeotsDRY/YnZH2JVfhO7yJ3tarhKvM0DAi68vXPSKn+wLlk
+yLztZqjmSgBzqbO6kgK+dqt9Qg68QHoxugqURlupY8z/VMbxV3AFGSq9UvM6CB3L86GoTuNBsnZ
bY8o2qTXUF62oZEm4ICVdWAAOl7A6o7XnsQfpkDClNuNHWQG0khFTgcY2NtXYEstE2MyWH5q7c9b
i4hXlRCqhBGtjuuIdKfeCPhdHUrZSZ70JiyHmJR8yHbW1ZRipwGjmXnPofZf+98CTmHLtNpOtc7L
NNrOFAbdIjgFvOJX104afDX8YBOODKwNUykwb8V93JgSSzIhVKwnuWUXNN+syU1iYXkpyGJXg4UV
OhEec5sy4ZMDu6NeWmdMwJCuapvej346mV1YZM1vYAvq5T6q0PzfUnPUmK5p8YddICc+i8s3cWZf
P/RQXbUuDvrZy9fVVFPgLEtmJBSfJMOhAfsSaALCl5OPU3/nWcXFzUR+l5847x/P/W5xg0e6Oy+k
RIFlcc8g/daamiqVbTQ7hxACGlzr4MqKkvPoN2Dz3VwoFPu4Z/Yg3XnHSKxGhYtKA8TyOT7VkdDN
42bVQjs+HqR+CVXB5TBogFrbnn2VmG/9Whmugn4thL0Q2ULVNyIBU9s6LS3eFQ8+vuaV9gFAm4e1
t17yP4AQ0srBkvjmBQah4qSGYlbNWbo8D0aggU4EErelyZAbqmz7dbZKvXmeDuVhTytuh2J9AaTI
66gQWTzfmib+VbiqZPxRh6x27uQjCO92tWitfev1VmvvWrgzCPN0TNS9fTE4ykDvhvpp03y4W+rx
kTsOf7y6MmmHibuEdCZ66XKVYuySO+knRwIB8+wTV+gZelMyjy0yzvjHa/j18BLLbQF3VdhaB3cG
CD/7vzvYqBIwkiNmvYDd6nBdLHCA3TmRAETA8/WYbgfJfRiT8yB230loJLF7XMSrTb4vOCDtZZqC
jF5aZX0hVYzccdiPdnrcKIpXGW+tVeYZ8jDeXS/0T8V/cu7y5vp4xR43WYK1wlysh4SpBNRXz74A
G6opmga90R6GJqrRcl6254v545bK8826eaKm2AvYakfgyMjOcx1gGotl9hnh2JeJgDNnusG0E4di
s8i1IXfDxhNZZ13CV7G7ghdIjgFPy9RVkFAfYH5zj3rdwroSg+CejxNkvEZzgbl4pKRpJuWO/ef2
7IJ1/WTT4AlknmoJLC0V/PYULRVvPIifv7Ey8Md0xII9oI7WI9FSLAY7wQ+RDUtY69YKmofagsli
cW0Ud5mHcP5HaAmwuh7mOzPC4nv2OznaxPnkD3vreNiSnyn73Hf8L0imtJS4RPEJs2Ak7njbOVqX
XmyTcBFlYbJQaqOVEBYeHt/xr2T2X0DH3yjVfxirMNBzqPLwhi0Zd03cqpKQFYGPkUavhHyEVdmf
Dy+1eotEdGNeTA3rTiO4Qi+mWFFHF6Wi7s+QCz8nvqVtMsrC2sWr8iEYvtoIHHIprw9bAWc2EPOi
8xDvbPlah/Yqlq+QY77imIb5R3zS7U/kddnE+8PDepBy7By4QzBB/YeIJYOO1W50aNt7IKuMfoHr
FDxOIw/j+P8xNlmbsvt+F4/AJ5Qz5D4mozojDEqmD6LCc9AUOifc6Of6plDj4acypeqyx837lrEt
RdqBweFTU7LYpeSPA0Q5fMPHYnZnznrhtJHjLHmLJSqpaV3NsGwSu843YQvAwZhvvbYfg4NtvLU/
J/S0Mw42RwnNY1TQzVuWYDeCdCKXh3ICZgzx8R51a/eOmwfTsYHPAWaB4A1iufA2dkBiRsipkW+y
WF6J48Y35PCw7Q6napiCqhGqkGG0APmQrpQ+607bG+v0NShIAkZCu1ZbcOr57UebToqSN+8E6BIq
IiMJ+y6rxeDbM/gsP5k53f/xWEiH31GnF46VCirOkBxgC3a8kMaJarAvnSHHFFzezKXC2wiUcXdH
LqawooMDkYY9Zs8MoHLseesrlGmup0NCqmkoWVPdrTz1kgznVMGOBAjpjbm8oMOxUaaKIrFzNh+a
EBig/tPVKZHPe4ySp5EeHsUB6fGzEjf2l0cyRFo/ktn89o1ch4bXnLAjSOPFpEbxJeOnPFxlv7+k
0M/07R1JBXV2AhVZBXsPT83P74vzxHVtbad4BFGsVxuo4Vo0sihdBbrROdCY7RT1KaBoPU6FyCaw
+0KsV9IItClHymf9483b+gnVwZW4u1jGRiNphA2ijUhp2/fxDtImUMMGeSBd7V0H62jdq6EMmxu3
uNmtOj3TXV7Vl7KShm/eUBOgyEzTmPM2VY/2QnDcgjZTnyUGo0+eXh1V+W2OpivYhhXiqSla+EhC
8+k7Qx7C9xhzqrNlO47xCrIXB8CV9SQO+qxCAuDkzJn5T3ixkL7K1y7qeOC3iJeANNczHyLxGNcG
mjoItB6Q9cCqPhsUOIBl/oqfMPkOPNmuU5NN/BxbRYGW3hEUmR5BGU9bI9SN+Yhuip9tQydqgWsh
oq2XfwMZZyV2aglbvryDJdyMM2BibpQadP77uqqv2TTOofQhcd+/OUwR2f7Ih3yyA9/OaqWz7E/Y
W72T9ear27L9dBpy5QiQXwLkL+xJpCbY1GxR83ihjMkWC579zMNrhspkpaJe7+dXjoOm1CKFKHKY
urlgNKg0Gx8+75xzhBOeeHTw/7pBHAPzI5NZmRojEQrCWFyMMQlk/GeFxNB4q8DQpJSyExzYg3UW
YAfaUsIuJtcpJ4b2VVrpjnwACFUzQYLVeFJXY0a8HfDoRzHAAnRz7h3p97h65TmKuRCVnQcXtjyl
u/cW2ecPCDHC1jXgRs6qbm3P5AAETzQxjtBq0NxPP7PajX75GTv8t7FahBhSOp1tPuBzsmku6Gl5
tBaQcv3LmAN/1xN4/uA7OrSZRaN8txHuebXtjREbVG8otsf8JDFMyVl4oQMnIZcS5rcfPbXRcwkW
SMG6H5hGqHHi4oXXh5iMnAvNST+zdKDC/f0uwO3jcKODRd2EI9QQiwq1RFb4vw1zH2CdFGxgUGLR
3CBhr8g1rXPFoUD1ZWtTUQWrdiCnEuxPdfdEbJx/X04Ifed9uCKUQ1je2WU1/x6WrylFj0FANxaU
H/ZQu+iH62JjdTY4R9PyTKnsPmgpkKlE3I44OhZXlKpq3D/KFC9Z8vqpXwg2SvrEBXfP7yHXJ5Dv
Nt/ns3HxElggc69cDg+fxLelftq4j+8iHKevPQ6gpNtHgZE4qV/v3wiWozxD8hWGrk34KJOqrmoG
kRNzL7VDfs+QfWIK8qKse5vMgHYcTIXsj9mHDeyaZDmyewyPAsKzaVgtNgdOAg2FtvZQBupk/8Ak
X4Kg+cPRq/B1bLBfd3hh91qwgUVLkmCR6bpi+qfIweCJbCD52OTR+xLVPGneE59zMQjS/Ohu3pzI
WyRFeZ0eThGbrHj5DoRddVVHu1g7p28VQhvaP6jul4mbmvWugrQe0zdHQ1sLZRSNY0ltxZZ304OC
hT0wcRYkKDmUujYfIurHPrrYmGJkzV5/lLk4POGEWb7fKWMKt9Dzv2V3WR3WuU78d9cdv84uO/4+
LQQVsMmrBaEhwomnH2wf5IClB+x08m5dS/px+1rSxg13eKyZHVMO4locUDFm3TU4X2xylpKv3GnL
On7NtmToYIGcPcZ8aDM1Z8GHU6V27JStYFjFvWXSUqcaldxREYkl4LHR1HXC6W0AJjc46MCHOsrx
pTh5436JhENpxMjoUiQjl/HCdw0g6GW1rgFsIIXyWpLdUgS+/EvGJ03bduuPuwLapaykmssnKRp9
VKEU4285SaunATaTz8C48ANrmWR+8lDDBh4/O2HrNxctZXADomBb7wQewThx3BKLa1IqqWZr2gYl
7tJm4V//B2AKUQWlHwdMHe+RzlbYBmfmjL6zGBuESPeKru3q44ga0Z2W6c5uy1+4AkdtcDT4PuZp
z+kOYLzNrnODE0+DaakTte3ugpN5Xd732NErzTUiGnzBMcfPnbL8cv5VVChabe32A8jknozPLFJ1
LvIi6LZwq51Nx3qOcV7xb2Qyp75VQg7WLRpJBGtmKoejUJYaPXXteILS3Rw0cBsx+H8fYg5vbsHS
vjLjPce5azJR2eWa4nMi8TPIUSUOFKLNM/yumY4WTvXDH/e+CnoJEBrPBNsxb/KDFotMdXMs9h6u
HWMLhLNAd9LLlXlO2E1KUpPMDl0UtHMVEW4sQrrGLSW+4eeLhxdbowNYJgUUxg085b7pzuQnburl
H91I58AKMtLrx3ajG4mKdVuuvZm2JWYSjk2EdFEiGtlqDPbiefUY+8htgpAI0xd2um8/ZQ3W+ORK
q2I7FoRwDe7zZ2dpgrHKpc4e5inYybTd9k/ae/PqUcxgwaSY13uOb4uH1sdTNZXTIhRS/KwSgq7i
/GGipMvsa8/3angHBqmIUs5a6noiAv48kYQvoiaxQJi0LAGeyU7uiowD7eMKaXlto7jpP5m8rsqY
FihgUY6sc2eo8q/6PUrxhgR7E2L+nBQ3/q/CQnalEUjB8S42SJbxRWrIyalUzqNfFQy3GHQHY1t2
JjCpcs4evh+PXbt8GfX1ioZtrG+1H1nmX9yT5nv/2b45ScezyuTWwtUBOQfeq0L2JKR7pPXAXjNP
Ri3NHJediMDUjr35+bzmuSfvt4ZZIwOQNdUKd/UjjoPHXDUukshTxdzn6tmi3QpZmVCg3AQciVNv
3E5qO7Fbgie5XvdaEujp003Yyon0h+lb8R9GtTn4wDQnYIGiVZ+JYJ7/8lJjEjurFWeqe1jt1Oeh
RwbyIy/JUa2w7C4liAa/F2E2vMKI315tBKg/0+IoZdSsT97pFjJcRbU7svWcOHvtvMBAwMmz49/I
Y7nJt0Mb4bZ5RnsLSRX7aRWOyJ3SIwpnxZm8osfyilK9c6uvgM+2WMNB/TFLDLrVAEKGAXQqDLuJ
Cvknw/0IvElfZ7YEvTjjX6BeHnrAhJzkc8fXPYuLAaoJCltIxwIK03gmpgZ9oTGGsxsyHo/T+EID
Svjxjtd+Tpo/cjEmhgCNB1uXCxR2PENnaAGX7N4TXm1NTM1sG1e0ipOryK0y8d8pH4p7DMJPV1mH
ZjszSn9Tymp8KsJOr+V7AERaNoP87qPurvmVAbadXJ1LG9XT041aF4/7SUHmPRhpqH+Y8mt4qrhO
pwMreoBTNkRqPpQnnc940vfUPHgqWCv7nnzz268Hhx+b6mozfLbySdK0brBStzVvkte9ZxiHcPB2
BTSs3VpWL+oRFNXZR9N+zaLwUhWMNHJIyiORaGXGT+y6ar+D8GRI5zfhuo8NmGuz/7vgEyN1tZYi
+FfTnu9ivHzfQRi+0g6r+3XrqGKSEw44cmm87voz28D49Xi7MeOPurK7WyMWhTL9p8oEuBtvgG7q
uY1Zl0s39w5Ir8NBGlNkd16scNQ5CUDhxjtr25jbMWJtLVjGjOdkddyqjT2TkTbZDuSzK+DGIoF/
65kJyELmknxZMC3qk6OxI7YSlBippmMO4L5rxBRzeMfZ6Rvx18ybCbOCDr5WNdrbWshZm/u1Zhom
4+howHwrD6spoyvF87t9T9h8+vroSmJmwgMX4DBzXMrzcJbizEWeVKEtuRXVO3D7wPeoVLhZvyJq
tpPOHITG73JhvNrnZknkgXudVc0deyfBrNNNeKlqlhy4l70ox1xHouzR55Mjnj2xzLsC6n9cGSpL
9+rbFhGh6Xm7MDyHjooSsGXLkUE23cazU5vG3Gh64K7V/NUJo/VnqlCweORGjso0TAiEfZ73tqr6
RjzbqUaVyIkuYC2/YMleickpZ1eXcX6ZujDWEzDJ+OX+TFy61WkyGvvPp8FAOhZOd7F49f/hXEO6
Hz/z2hSxXFAF2zocYXowaGLZdch6Rzo0EJgOZAtViQKGb3q18JISbjasL+Ct+p+7kCzMUvr3kAnb
yi+A0/mPGx5MecscnRs1aNr54ckEArqHt3a6QiwXnrkJPf8jiYqaMpqdkL2ayysl1oAbIQVAQd0a
nyy+p7cU+cSjxdpUyvA0EvtIqjI3jRwSjlZYRP50voKIHjrpCFPXHJLXUDFngCcBNpcUbCLEco5r
Oqme9GFYZyKy43TPv0P1JZBiuSCLXUAjRCh//YYPOANOx1yiKq4U3/f3+qmtnWd1iu4EUDwRE2MH
R4tH/qwgFv0AqYwOD0I00oApsVAIQVI+iXyssjMseDVBkAH2mJRS+nEbzO1dfknxwKTXXKeFBBaG
7qam6O0+88wgw7cUR6hPd6UvaKKsEhhZidUbwLTOgy1ItzBsFmOdsRu7ilB2TDautvuH+x8aC9Fl
q1MORfQi5XA55k7UkxLDag/bCPdYRQ2Dhg93/VxZQ4u+B5vB0cJOUbx4kq5m4oq4uMctRp8M4MP/
KrrHPDCXP2PxZrurK6PG+GV0G6G/eT7bJuLhq7zE1V882HB9T8JaPeXOh6CmWkIHwYcUUYz9KWfx
hMH+Tvcb2usLY6GxZw808YJXCg9rfUYzKFFrbSIbyshrKv7wiyGcGkrfZ68sVFb5B1xG99crHF0j
KA9sqFp6g3eCpN0Zs4fKj2G99+TOnfEuUc1/IgHnbBNFvKgV9lN0Nw9dkmuI1cJLrwQiBbAP2zGG
BCbeS9BNfuMrLpqbxuLA5YZfMLcLI0yLkOC2QkpuHbQgxsm6+MxL2p9++xMvPOdaIs+ikwW7fS7Q
edK4zyt5QzOjkYHAYu4UIoozGYOOQ52FMXADdH0AG+hnB9iB9i2OhS9xTpDQcUpBNNVU44NFiRCS
Uj8slf9zkOa8Yoag6UBq2anZwl5DtYQEpr8KMK7tKdlUCGcB/cwh1ep431EX1e2sOF/fooyDfJUV
pZ0+1r/PA/kTrmUTENyXtTaXOnO2WQro+y5Yz3iYM/1WDGdGVoK4Jy0DcEaRISIUCVt3o2oNBiFy
j6zpL/G+Ffl/cwlZcAb9Bgpx8x61IAWOp7u1Gscbt91fnzrtVwmN65dZLtjWvLA+V4nd/rtfB9V+
11ja6ncF8mQwzi8xABvdvHhnsTNStUjA6VRu2XcCB4Nu10bgBp+quQDxCUd9aMFkzAdF2ap4xcv2
ez6Jn/3dMSjZ3j1235F5sGIXPs5EkpCst/i9R1+XYwsRXLSRVr+LPAARftd3vTj3+gfRYuV7wPkk
Hf3CWKyYZA7rzmjn1GDKRf8Zo1zQIMV3WzOsuRh10IQo+9zT23u4TYeuDLT25/waBNpPqzR1/2CY
+Jql64HNNFknkJpWLlOXo+PZaKLSq2AX6P8IC8ILBeHras2G0XCaJq/umrMZY7zqjY3BoggfpA7/
4FCTe2lz+FzTbJoKK1D3elsdb3cZCnYAZ3/C+F3iZ1FrXU2Qt2PqYXzEFkMUAn0CUeILd3DzU52/
uxwvl/M4xAnyyhEAxPFlQfpq+YdP+3uyuYI8UzR7ZP07vODkV1n07q9IhnV9lK+vmTgRdYWUhFPB
pFfYLOdQM06vlvvWYUo7SgMRpwfUTkHsy1LS3FK7/8MJGHn5tfrO2uAYph3zdJpCsvbx4fABtC2G
6Ev+tyXQcM84Ur+hnQaVFrQkCyLglZONkp3rqSCWDbIJEPx7SYdRVUqboKv1W/OFC88TzVA1K2lo
b9adhMVZEVbE1CmX8DL0T1awKSIMS1eQdRfHSg0e1LnEYabCfZKxOeO0EOYbbwtmYyX5vPsZM99v
k6M24ZvsZImh06AIa+n4n+46JEXcdypEdVuUlc8psD43z6KKuiONWFPkAZV7ltYCO/YN3g3HfbUG
X9BBMayhb0jvJya1KKivCoWF5erMPizmOzxrKntBZN/+BawbqenZ85eDEi2pMl0zhxphsMhLdwqG
k+QWuFIlelND2iJABH/e0YizBIZGf+ry6UZV2UnrU9jgJCv07Bsg9pTB05wzap0gCxLb9GlTrELS
swBme42Fteh/werz3Nk0IeB++ctD9QzGrGUmENmGJXp1zmXpkzfbGwtVYHEtdIsb549JZLhXvrow
TJjg3/xpMJ6VdSbtv9XoA3ItkKp/dizlemEXT1z/KqtGnVKs/n7Rrf1v1T72+4H9+J3Iv0AO6GpM
yMnKp1QsHuC04y7bO6jTSEIBoUckKaxG0ZZ6FfA1paB1z403+I4u22GO9eFcpH/q+8gCp/Rw1qza
VlJu7I4Dw39LRK6ezoOM0DeQP+2pkK8YRsSr8L99FqL9q/CKsdcsJUkwSYt+6gPk9Tvs6Brxrs9d
klejq/eR2wZh4x9xFQpVFYu4QZER3KFQKe6bj/f/alUZ+KUhMzMsnQ/wVkN8r/ZyVNCQDhsi8QQZ
CnI/qnhpotteieUS7GWxHk0DbCnHDap4NGcKo4lT9o8nWlEjH16JQYnNOGW72hVSo1nc+lwoexoh
YZv8T3hX+8KH+JAP0cwt6L0Z7OfZcXt79HeTTCbBcB9bGulpWd/D5ienPdCxsH6uPQ0i5DmLnhc9
HEng2bKsr3qooQVB0QX2/s6f7wzEqIhVfHIBvYqTq0/tkSGnSLcO4SYtTh5I2ilZvmMIisgAUdlM
mxv0e3mPykHj6VogMl42MJYKjaMHX2sutowtBXYZzB7mvpnPh5tWczMWEUybsANey4MM6zbysa0k
8ksk38SxDWwAMot+cgQEMrOPENnea4gkZ7HgmtQ5XeUNeMjucj2GmS5X3UP/GFc3veFURblMMzRU
qX19GlPylBJjmXx8V85BoCPIF182/9bNrpYCHreYkZPWrkTlGs9xxZD7t/84LxhRAJJapnglH8T/
Ue6tCS8NRGGG+JulxuVybIjlnghabr7XbgT3kROVYLFg2Le0+pAdh+UK1NOh+y418kHaEoR/5X01
AvBkpbGF83abk8glVnZHuFacWraFPYs820u7Wv9xWLKXV2Ks+SA2IcOBnBREUIa7aP4ND3jA/o5o
5X1CbXKO2oVlFxNu6y/47GGP3Yh9KnftRio5f/MDpbhQJ/yPfZoa8KKTT4tt8+tBia//0fuTdqC2
kgpjDL2PCeSiAeqBsgowCD1Vpr8DV0VuTyQaDQz0b5ImEU6fblIjzC4hTWgECzvd5uB31uLepAOq
7c0dy+SRIT3pFkMO1gKpeTa3PWlunpdewA734kUCZVDe3rlF64sXG0753dKw56svqnNyRpqa+58v
a359XRoZcRVoZtdvskdBXROSe7Pd7MeR/jz81SwaHuaoEqvFtqXj4MH4nn2xfhXegIbNiaxR94aT
ObZ7espdTeFWRDhr6N2OimA/1MAMvkujM/V51/f+HANa6Ee9LKYXO0UwJ0Pmw7BKrb6KC67WWjnH
L3e4p3AproGYsM/eMWWxtt8OSC/t0LXmDiKS7zaQ31wF0V3GC0cq2H318SRidRPd65MDsZ9GHWiS
NP91xiRgIFWWDJ/kvMSGrwxV32nDOk2nek7Vl/v/THIrkEsCdnbN0WIqMfTuWlQF2VNEddisJzX/
kkf7UZjt4AefKiMW0AA49YRfmNjd1qLhNrYBODV4ZeLUYE6RZ0tyWmJWk6vdtvtOn9dKUPvfW3jF
4VN5eqp1r9c/tVDvPg304k0NqU+1HN2DPTALaDR9luHwHer0R9Mn5EO18yjls/d2zM8xnOuDJL3+
C22X00gNlCmtVcYn3Xfw+6msGS8s1cZ9rvGPsoUYoczkD1mtPfSbHF2uf0YylJhEnYcv4INiPP1t
hFzaBPB5I4KiTzWID83/NpPcJc3sxz80O37OYyyjx4QU6G6geJP1tbHvlNbq4E9cRrHXKnkZF70g
1KMRYHme+mJZXtXMxPm9xoqtlVwhwnXWzAY/NDYvRaZMQLLdjNVcl84g1N/JNRMvva68TAvUdbDz
IHv+esLXJNrH4NZzVI8raFqGsUq3VRTi+9ewcASWv6xjcgmsH+sJPRpRVf0NM70u5yT8IZhAVahJ
FDPKLQ1WFfo9FqcE+/JqFV/n2Ai93UuKshawr/4wa66abHWlh2OLYBJ5u9ZM7KLWXT7G60t435mK
ms/RDzuZOE1TUo9HUqN6e/E7qbLcOSEZ+Du78nV66Dgz4yZIqH1WJrCrynN/q3kwfDUkBQDSEddI
tsqBFDKe5I1IDJ/FFGXCW6EoqlJn49WISdei5HXs33cdjvQ4dK3jYbZp7fghgt0Jja6Zbn/rpKm+
v+oMedIkZqAfWzhvZYtwhsYsLZ3LanHXX3FvoQ5cN/mVxVEer4lxYxSsJwtvGeQOFNTS5IsEESPH
dxXnnfh/rGALAng2zZe+MtH76iEwN98v7WvdijcUcn2NHU2xqTuiod9hyVYpqjUmWOO5Y3bP4hk3
gmcEgMND5aj1//00oAYn8pSwQu3yWbjSmgAR7gb+MzlQoE3Gli0BGMwZpZ02+RiLC88Uue3DAZmZ
BhrI8q9jIM1qvChclQddTb+DGueZLu7ifgfA7JOGatrar46lVN49OrsljLZ15/KrKwrNK67PMHE0
zpWKdgoaSfnfSIeLd+rpxTqn1eRuNq2+YrvXySPyitaioafmPAMijkShNU7I58ySz52jgUSaJKzh
6+vJ9MoRVpPyCis9GTRW3ixhVbXP6JmVclHKd82JbIDyjD6jjfoOWzlbCl5Gj8DZkSPNE8jU3Ovw
rQ5tHKbG4KkaTxApkWxANBOD2Veodq+aI3bUiSFq6coLNqmrtQMAcEuE5R0QWTPm6FrBnLJ4OhmD
O3LuBlyCtzAgwzpMi+qnqFGzzO3n6Hmmo9fxZ0sDvGmpq190aUDLXUIFS0elwHfrV4kDpl/r2Sw1
ryyBnUgLzvmGtK3q76D5rJr0eaLa9sgTQpKa4s6Bd4WGTPYsQ6GGKlD5rQuBgoIPaLkfuQTC4VmD
dmXuxT1nWHtaH2JwjiGDxTDKNMzxfqXHAKSvOJ3DZOPR6m/npbeiFW92XkPcEtg1wPLClCtsY6Sb
f0tUah7HluxA7wlqYWH3p3KXKTZ1tzOZO2D2C3MrAk7JbLTynkXgEOIRof641V++X8L7KrPUQ/Xd
y0gDNatcTGIzgqECLWrW+rUPB4OzXsrGa7ZOkg6nPQYRTc/y9xFXbrJXwzTbPrB18fmlAfoan3lp
jOj9+GsoLP4Tfwn0bds4HgZRFOCL6Hak3bFdnkECFjqNoUs84rRXP0APMUdxt6vW1MQArDJIUK4h
EYWn5LrwRBkdgD3RHG8rjkEdCC26GszQLJuDdASC5OSP6RIlj0bIZP/joPtPZ2vHTsLl9MhxKAiN
1O3HopbZ6XzJycbdAfQ+oDK4dai8tMDXGoGfKZKHVv+0rB92fB/znFRSIzU/aQqZBXr8sGUeM7u+
zJj0WOlohtDie48JiuufIx4j4WneDqOTit+WheIMpBa2fMAKc66TUczz6yS72gZynUkEeWPdGmqK
ehxM2b59kDbtRZwg3yvKwnERDP5oxn2/rwbvvAWhDJBO6/+tmJ9mPVYbSkRHVs6zfWx46qEO2+gI
ciT0wmENZBSsNKzqN/Jst8ZR1cV/yN/Dg7ID4MAwUuIZH2kUrcOBL1eDycoTo9ApgPQ3nyiEuaEl
mBmNDlmUOLzPgLUl/9Ol1A+fy8MktZnT99NDciHRo6ZJQNEsyQTTQnqcKPlqS2rvFh8n3HlJT/UH
+h93R3vio9Uyci30wlaoxwi90VVRY488QsW4I23M4XHc/0U8I5xDUZl431lfSaWQQ4Egpya0Yk7i
aIOB/014WGw27R6tqddtVBnPRks9JxuKsFFSySmlpwhFQFxNr2JC8597D7JK+UaVqG3MmfHYZnAm
hM7aVZKt/tMoiMpP4JOaDf6S3xXXk/wJECfCXlHbe6mBQnX90tcDc9b9PXzW6sIn5J2uEmSCgxXR
F20wgREJEi1+CjG1Td8AAt1bhEhgAAxj9ZqCoeMYBdS1P/9AW6rKLwa719XYLZtMYrcf2XWZvSdH
MTpqUPkTcAwnqe5DvKywukKg7jSS5taAsM/TpDlt9C+U+K1Fr4vkL6efTrrBLywdbM0NRc3ulF8P
eX0B8rVvARJXOINECEe6qol7gTSrxlX2rUtpnFYDHZ5n6xlv7kGtu1/0zciDG6OX3OgHol74IeIQ
9a5hNP7pf5HnRM+QxeVXu5GTvJSUBgQkTtKoMEgVy9ZREtBwKNQBOqDsooQ1g68gRZJ7bIkmiLvG
fciRSTtAD5UyBR5wav6nlUkyh4eIPqc1VTPgNLzgPXwoIt469uY6OT+ssqvepWGoHeTQoi6P8pv2
wzRuTgjp1JrfrNhwazpQEHSb6zvBVaUP7Aze0v7lb+0KHLCJO0g0o8yupeea9JY/RGqCqeeCWJJH
8Z8YyycM84OdY0RpbeucdIwt7jvmq+YT66ltmGvvIczrycBzWl/DKOyADDB6aZF9a3mw93Nf73SZ
NJDiJvcUlCmselDH3Ty30/exYol3NKZSI/Bol4cMdiXrrYjRx5lO2W3zi4PSas4wiIU1VSF2EqJO
hoy6LUcPWdFPXrAH3zOrZI1hGM6AmsFqSOGkCWk1aC1120PL++pke3IzWEzwakr5lkZmqVSASbQU
jRP9NHoCfU7TBN2qE0SiT+QZnja1Am65VAHxwHrA5uKAoNUD/JAe3vwqopPXzuJNrO+GOSUWCX5m
TLO/mxfmW3D7N3fRcU8vsoErZ3fr6wwdjwlqEq2CIpiWgM0+BBFxXeI=
`pragma protect end_protected
