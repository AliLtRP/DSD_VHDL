// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:47 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
c6k99ZhCkCpFQdG2al7uZ3IWSWgLK9UEPdGvm6d89XJwxZnfeY7nolfe2Lgl5VZm
7l4nuPbJ41/DI4OF/BlpnBEucJPs0gXogKNwO+TmGRwpnCQrQ5KeOgTnIxT1dgmR
Gvoe1jmnirhD0HgLJaZe9FCG626g3R5LehRsY6IaHoI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13824)
AfEPECan9dOZ+mG1zlLrT2vSkZa3ABSKpY6/2DwlHi+sS/fBAwJs0Xxo/VwfG2ab
WDIJdnT1nLk5yTCGjnJ82IpkGARQUciYlAww3rJrrVldDjUujGB8soqoYZMdIoQ5
eop/PUJc8BOnvjYGnhf+p1wCEOpIMbcQC2C0jxkPYzUUVyN2pjuK7EmvDzwwHN9j
WUFkk+TcmmBTF7AIxiAcYSEs3cgBPV4guXqDMIFG0rT+haYXBnJqrNflb/oELWWY
doHNvr5spdzNceytifmiGNFBOhqXhPwCFOBirHHxJ4v7n0zuoVOoRIDJhimYR8aV
pJqc8tkqVeQeR5jqRjE1cBIM2iRMJF+pEbBf/7eM3YXKeldZC4DoyFjjwLfQABHT
BJvVI7rdNc91m+LjcHTsOkVAzMJTJZA9HMz9fhaQl4m0eOtmgQzuclsaF3hBCAgE
/lmkKVRIwjr00j2HK8dW48PTArptptjyISSQLKBCfOYdVM9UG9y5kb6sTGubz5sd
P61AWfgHbffws+BM0CSwf2KkQVNL7KkkVav7Idxg+SqgDiEVLtmT2hIL1Q4tX5Q4
L6BcGjNqSY817yKvzTu33krtnIw5cbzJ2YA11WIdSI9eO/RcYr44ORBc5noas2ti
KtBl6WX/9G6+Q4W184DO+NO6pnuYC0gk+8YE4j5BUTpntoUYzjcc57zqNpW+xjTz
EjbIYOhoQteXkBsoWtBDJFzaphivt1FHpGTm1lYvxLAJh48N+kI/1j6uMiAfaep6
AUT8DFGHw7m7vUvEMU9JHDLQR71po7FeY8clu5bto9A31B2wTzFMn3xUGH+83QmT
RYyPQtfjxApeXNuaUAmfBkDRgpN350PpxkQlFzoM43VwGb3FUSUUdVRkvXPbx+9E
4OlGF+ru1Neu68mBMl6M+2ukwHQR9r7vW/LGj7xcD9wH8A/JKJi+NRUiwGzIooEv
pk+gvkHnCSln3fs/Ls9igPbBJZav6oj/JmJwmkBsuDFnQhxD5MHj8ibpIzStS2pO
eqTw3O8+9mOGJwB48ZgtXeNECtSw9qTs8RHT7wKgqMAr4vE0mRyocA7eTlVWGHtH
+Qu9v3gGJHan1QblteLIhHDAHJY9jGtpPJ8HCXei+tf9VRxuZQYHonjyYL5Exnev
KJyEFe/XtaDWWM8pE4QsJ/Dw6P/0JeGT4gdR5Q3XSqX0ucJoNb0wLnHpa9alN0/G
VgxHv/NtPgjSi7hhKb2cX/YAYQKW4a+cfUAqRaY/1+/OL1GwkRWIk55eCcJ+Dr+d
yv7rRJemtWsxREAelQj/eqJ5Ce+0xpO19MgHM5MbLuNKJNJJUTN382PvN2JKX7c5
oYLUHKkyqgtAgaXZja/8e/sKa3cWnIygOOB0zjV0o/sBLPFsrxMFok+RHsShu82r
ODLIizuhHd2i6OJTblVBQNaxo7Nm/GJcme0oANhXoNHDM/bF/9muXp9mRtGSTzay
onQyXg4yL8YrGnaSgpk4MFY6UV7w4GXV2lXC0VK6Ca3uKtcpjov3XwJJc0KjBE73
MKOhC/hS3l/52zpVdrAxwC+5AF/ubNIxoQ7LMPJ3NUxTHACHPv+sdTpDYnueShB0
MMjGTZhsMjNY3ZMyJs2llYP7HbSTnAST+Q8nuLvUowjdJ4JKDYtSfbTcL9ciP1Y7
H8E8LL1kPUO+BX7JwDH2hkpsqbk/HnL1rhNIuQX2gk562jHduly+DiU8MSVlHQGi
BxmVv+feJ+RobF4RklnnLGeqrpK9H66g82MCeQTxI7qHPJnlwu6/FB24psFDh2er
FFxjDvKnL/82t088aMXYocNgaa8M57OqULxqUNeDQGsRX9sYEAuehIMr9FaU2/GD
f93TeCO3DJXGxmZr8U3LrTnZpYNKyxVck2nm+g/wfNdLNyU6f6Ut9mpYx0qmt1DB
NZ0d/tra8zZdDs0FeZK/hnytIFD1uuv2EfwBDzz/uRDqMePGRXHrSD6G1Z/Z7DbL
B+NDOR9NQPG0VHqVR2hOK0Yq4XLlUcx6iIguyiz7bB59mJ0IV60isgPnR9ZASjKw
oTewgNsX/kHjTGd5t4mEyN96JedqQiFNQCLJ6Cjxm1VHLw4doyUAvAb19+mbDWR3
vRdP+/ZnBOZ4SpjCG0kAo5YAxeMXpKV20Ot6HAgultprsKfUM+K+SCodN854wmlJ
+cLWJwGbv066Yb0qKOnBevqwXlbQi9DYMmdqqmwWaorzimUIiPlltAdiUp+gNgWQ
GRjuGyCey+B49cBDAjmuki4naIBsqL6kSKJtpvWcjAX7wuvvbNGAGTGQz0AxxgF/
uxF851ZTDQvHugXJ85Mm7O2haIhK6ENx8aZQDjdoiFUsgwujvnIG+bROq2WvWxBp
gqHEshke/EvBXZbiaj3zjSWkpB0wdoHshexBoKlV8sgZLx2G+ZSygduscbFkQygv
tQXZPe6F2Gkgqj3QN3epV+BElKTJbze3nRbEuKZ3Mt4WEVdaXng+raWbFZi4rmty
53KdFhR2fSKX7rJ+CG5D0XrmLJHVnuCmkG9NpaL3f2HD2nys8R/9tcQwyT1ILDSw
+jQr5A7Sge3NZTpS+cvfZrFRH3cBJ6pJmBsQ8EQsdGxihqmK0GpikVndRemoUO/Q
yUlwIvQSxEHxGAdwDab7wQaEJcIMiNUrB7syP3BA+XNEispMo3veJUUnSdv81z/i
6MV1FC6+BT6hS8mrgaBqA10f36Yncjhh2eMVUgyt3OzlnCz3zo+mvrqpkGZ2xv3S
UBkjtsKBW7t7J8biWsBOrsadvCIusl9Mx8aQsvAQBd2D/SW7aDBdw2Kj7Dmt0pJf
yWrkAKWhGFAV79PzVp2yuHn12/UAxNSveFWtW5uhLHquepuqRp6wVmq25pOYBXT1
oK9v3m07OFvYwdplcOxaXPA3qRy/ZPqwGaIHKSpeXrFprcYeLhBaIsCSWy+S2tGd
de8fCAl7Hb5utox5mAjA4pb+uAYi/vwuCDTk/Pgcd8+yW7RxpXLeNQu52pmV5/yc
hRBYEgUiXmrLDKOhUvv0rfify9GVgniZVBpdAolWQeW/qL0g+ZlxgJrWgSJAgIxD
GsgzlcrR82FRyXsuTh2TKzVq/FUn4BLfGxoN02w2Gp89wIlzQpu5t+nxcNiGeQZA
qjkkrtqOvHX/jeuhgm8qGjGSYJ5gS+xbgY+DEOCrgVFmvAzERebGllxpUR9c96rO
E/F01CXSPY6uqoONpC4VqFUGxcHto0/k3RJ8S13XaNC0fJrC1lGhywxhDbr5L3LX
TRwUjsRrsf6iF1siWkrAhMIYEn61phKlH9eWJrOJmQ3sgKHPKwnmuV4/BlQB/g5K
1ZLr2/1/oEnbwriinSGUtX3WiCCzVHoKVT53bbSaxwRMnWfPjEh87F1ER+rslmZK
+F+jQo0zto+wLUY9a/iYzgO5BQufIacL8mBBO17MztQ+x2vIzwrjm/ga5We1usOv
Gyvtx3XiIn/XzoIDM2KgsKZUHlTN47WH+C0eFNqDB+bao35rWxv+VoXo5mOHskZe
Ggog0sGGz4x9HqW7U6q6QItjTLtAfhdOmSi4Jx/vg6GHFa9QLA3P7Rl8Ve8gm6Zh
Kh9NdNa4CfeAmiEbhOFICtOrMEWl1pzgAbKKraqXQaQxAObymQVWPIardeZ+pdSp
WgHyhFBzm4bDNNynNM5EMgJmAlj3f/LDSNkLSu9T7oZdkatonYfIESF+TKJtbMKx
xdTEQnCLlO4bQWkY7qINkz9zjskOhu+3dcsNVQZHJ4u46Vro0ct9MEBE47kiPX/b
vGK882xeYzXbPuOtLjK45TH3dyR5E//MAvVTSVyT2Bs9UO9aAbNLDiiYzQt6gOD4
7IVZUAoN4wC1xEuKMYzen8ssWOl9Xtdo8DqMQv6eZje8RsyJoufWxD6YVN9e6KdJ
PXPz2s3NjT+PDRi9TWXEKwP9/fCBOarzSCwlnblOWUD7i7BTzlre/YYJJG7EHBtn
vjjcH399svokQdcgQKzSnA4zAK8ZzReN8GXaLuwavBg5yog//P3TGLE6WFZB27dT
7RqSIM1ga2Q24OQbBJO5pz5c0BBMiI2InNRnJPAquMNJ2W5fEBmKPFMNjek2fNjs
5Vfhj9+8+OSsuQQRXSwMZUZF0Xx5mdXv9Iic/AIGdb4M1oPp3FQ6DTkyWj1lXlD1
6Z6vBLvs8fvYpWarFOCUqMx7BCslyVIjjezBTdkvmpEuX1InN1avFKApdOIhD5UK
Z/DV45S1Ed6fbs3KeCE5TOx9gxnsOT4H7mdh37gtnuCtqQhHyewsYdr8lbKndbzO
yKeQfx+we7M+zpmhwIkna/0D2QwdU/kpfzzXZD5MZWr8BQNeUBwqszMtDoExAzMX
NZLhAULQI9ZaG3bo8SiD3wgHMrIEx0320JzS11zowI1ux48faoTuQSu22YkUya9z
SbMumTWTLuw68lrAAS2H6rViZ+fcUjuuWjVTcFbez6INh56mFSaGGgVka7/z1lJg
5eMpbr9RognO1C8gZAJjPlQiL3510pzJBQeml33SPHKSFfTSAyOUFiH1SyYBNpv1
ksxtr0Am/HwMq+TwvGNcxRB7fHXw6oxGaUrKFzf9mBT9xPew3hi0XvbSdNGbJSSe
/7moJLrnR+uJ7JD9PtYIe1SGux0Ax7kNo9EEKmu2zHY6oNdGeK7xY6W84rUK81Mo
yNYfeKpYhiBBukcS09h/bUFHnVWHh/M9qp4tMw/kVPEWjZ28CRN31szfLJ8SY37u
YVDF3r8hHFMcGkBmBrKIN73EMnFBES3DmeWunAe9AdxQBFVgvMWrokDI9/QmknuS
hYs3374HmGUY8/SCRy90GtCsjyWl7pVdhjDq1AcAF8zqTuQtroVE9XVmQ9XE5W1U
Hh+A9Gll9OZqC7YOwurUwjimMj9mUcqS4JytVJqSeXkVWXO/uSXK9AW1dRRU7Wqp
xUwPZ75cuzfctRmJ+ouvJp/o1M/sN7duwCfBsqKSxyr1XlibxBir2j9IyNQNSdd8
uNi+eCBOcyi/2kTSOmEpV1LHKCoEWZCk0lExipjiJuS8kR2jFXAIj6rOHrxu9eX4
vENnSW33zlnhA9uqal2Tm+w0gewJQ4sKnzBilOgH8ZMSZfHGSnucjZGEhpm33hp0
vdv8e3yv5YSsQgHDEz76DJ0ik0/rIZyrpZGnSvXXJYtlSk81cbHuMeY/RtvjTKQz
cIrTxfaj8We9lkGn7S0iOJhhVOH1ZFmyxYH/4u0wvQZi25MLwnNU/DmZ5Qekd9h4
8wb9LKLxSS7t5LzNKH8rvc23YnySKQ5qVLPBZWMD232e6bLjGMbI4krmJQFEx7v0
iPpu7A7cG6jevcGJKiDR2TcyJ2q0DEgR7NlbSFXMeKxvKB8wAYcu+RKm9xoKDJOU
lJWUhniIUjwezWl+3mO0WVD6LeXXhEr/JMj352JLeqQmkgmzL5h9bsLD8SAJcox5
XlKdDf/OQpNn/gIgr1FQHK/rGGp+DQdggJMQetqIde9VlIP6DK59l/J32jXPe9wX
uDKLQIxLV+vzDCDIGKvRbcfI2ajAXINL9zZLSwCcmrkN4O3MAujWt+dBE/hJsLvX
REBmBRYjEXVvqA35d1Ht+Djcr7sShwaUTUN4tq/yXiBUQncD73WZP2TOcoJ6liKr
nBbuRyqtigqbkJlXKw7rrC+eHN4+zgMRxU01QRAqZHEQqJlnGhYUklLeOfU4gPFb
GVkB8bgbY1z03KdvbehdctCYerJKtka/jpAeJNR4zx07Ez5YLrcVULwkAvD4pOkR
MUlp5fb/jsQ0CXeoyZOD2eQqCbWdZ/FpLUjJDZFkKSjmgBoOqpNXxExwGMcV9FWu
LMQge1UIUMjWqCm9dva7ar4BTA9gwm2DMpdx2ZytVH+ucfrpTPQVuWgxmPRptdP7
n9Ailg6/6LmEtfBTFj6lSdSkdnByRAaZbcQbVU4mzMaBSXc4Tm6fEnRX0a2Cajfa
Our/djNprWqzyQmvtP9b3pgiaXwVYdOmAjQ+DoJI/YjezZh/Op5CuMZKOQVDYpo+
wQPXyx20k8cn+0yjizN24rs3BrVAU/bVPMflnsMxbkPpdn+bIzB3vfy22qS7waK6
VpP+qztP6OKLJFpyo7dGsXyA9Hy08OhTqX1LU+iJvIjLlx6tK60PzjQd5/+Sx5Ry
JmooqIr5QhzVe0ot8HJqiVy/n2Y0B7p4cxHtRuy+CJOTqgQEF9IaOEynt9hoWOL0
I5NzGNRHglL3lh4gqsvGv/TS1qMlRzldY6t/wZouD7R/qPfB+tBMvpESA/xKewd+
b505QEyk5ON5tgE6k0uPkj0SVTmOLsdWK0mJXyg1zWm3U6MkFeicNi0r84oTr/r2
qjeTQBVuQXWKPXf7V/5jT/7XkfnXinFSugsxF8XlvIuldFLKu4A4MFM6dYn4mET0
SGGJSczcuBFaWABPpQz0xnaRfbIFMt9SU7tyIdVkxFAFjs/f8UsWaCpq5Y5mAuyn
Qt+rG6uCBqPXuUuqIyS+Fc/J4w12DgmnOP6TF85kAG0KKAqnCpflkB4hPL5ikmb2
uvGAyt/pBzXUKQILb7FX109zui5Y6xiPZ2xAj6qfDVGxmj/xsrbG8iq5VRnP8dLk
kdJadyj46Vr1L4LQTsRq5E/DUnxfscoEyjHryjh2Sc+q0uuqodJYcQSz3IxEvDi4
L8KkmRDl4EEWKhnKTHVjuKr/wpBEOuT5WrE1EAnqdV0jy6p7w1nIL8KDkgVeIMVY
eYLQ0cIRvW0W1/dRZrDY4HfJef3DL/EfthwmCxBUYqggpd59iDyjK/htba/Fg7JK
Qd3H88ofzSWtDOSII0pNZ4wQkvESbTZNqxptTmCZPKhGYwaF52RS7njQrgUiN4Xl
cae6E7QkKfo4ck4/piualFQPru0eN5E69/UzCimmYYVsqoR6ulU65wh6J9Mhr0WZ
3vaocA4ojPfN5N8/oXPFTg32ppiM3/GoLf1L7zFj8xi7dEb9SEem7zj2xavfh1ZF
okX8UAyeY3jBrO1dCyV5yw+cOgs/TgHbw+rZRCqQjWnTsUwPOk520oP67uoc3/7B
SKnBTDhBniwX61V/0mQjhCQuvKi/92au/Go3lc2xZExYeD9Nje9XrC9ME2SNr7JY
FFQ4rlZ7N/GiepwOunVCx7In2VVEBr/V3x8uHzEoSGsPRi5gYvVsW8JfsUDqcWp7
exfLxSVggmlB9GK992c7T2ZOXVSm7brQA+4byNcMC2yk4i/zS38Dz4RJpvrfkm7T
lTKuaUqxKhOMUOI3F+1BfVsmXaM4GF8egXXAXZpetlsm2uzC8wviHhpdQODuulC7
3MRNpGvknZVq/YcMpIKqrB/Ss+aD6AoddlwVU4ScDpHxFFCn9ccbYbOqv2KYvHX0
fpICH8Q5w/pPh8qecUfYun3y6lR/cj0LZ6jihNc6TgUP4aY6obzvLwhLRoL5Jk0m
s0rIHyXCfCIkYelpsZ8oYTOJKdHMhRNsDGrCBdYGIH6DXYdlvnPDDJMfISfZlmIx
G6ZYbNVBpXIX2yBFJHbtCLGWtl1BPO+Rr6OpYV41ea1eWo+rAEO5daf1Z2eu6wuZ
J1LI/x2N/LclHcdKieA1faSS//N2SsjQGswQMPxgwS7t4/nWs/1rGJH+DwY1Wzup
+bOP1EcevWJAYQhTtWef22XmLc1UNGlhV75bngh6wGUGq9OfMzDxy1TS+ATZ9KH4
5sCRPbbG7buMUyEPjRGEfKAS6+VoCviL8+UPl+FJ9/pcjLdxmvqUrWx67yfefPSK
fPz3NQAEQ5hOBedIdGDHd69sBV+HDhVJpFzvFk48OWvDd/ScHUssh+IpC3TVHlsO
gwrZarfIou2XbBwLe1VEo28UMr5dMQpuGgjwQW4ilU+vr+KJYo9QuTx8sWlN2r1f
CuBFh7cGi9g/lY38F6ccQnAW3AAas+q9l2NH6pTA0iAJ8lH1HH3NpUxbPVMPqlP/
2ronabON065HC+XG6vt3zSZltKTOna4AyJzCd7Uv05Rq2BGjHNqzXPvo5s54Tv9U
f/c5inKB1pQROPkzcu+xxQeFC9X8jAClwGMFV7oSas6Og5Xk9tl3fk6WI7YFVFHB
t7lTajCrEH6z/bi5ESeTaOclJqdReVRJFEDpvZk9PLqfYtVro4F/DoiPYycPE70k
Q1fj5e6bdcFROkIq37/pnupfgxKOV4xXi5tuLKYAAP/vqFHQiyeSypoCyHTswtL9
ccdpQDW7UYprqA0ddOs26hXB2nXPKwKeCulfVRlPFxq7RB5I+A7cZ5Oz/asovvS4
nSm5a19lgnpzqiGRa899QMFwmuyyIVxrRZxEil27CjkP+9IKYvo9Sa+pXHSzDnLT
9ZCUviABR9iRqRepiawftK1SUw+/BXjmAVg7KSGeGwTHbsXIL4pfIdyrS56i4NSq
s6voZCYBctSYdwvBAe07BAoFL1ALW+qi185yKjFvFqinf7loYRKMEF9cQ0D2XMO6
1sdmSW53OJzjy9LRxGv5GW6h0vqxTUfVL40YLgTBUboWjUSAE++77oU3hr0e7aVq
Uujk0W4WPpVhg0t9PDAzj2rpl2qDgK/VGri0weOFb5Aak0gwFCLR15IuWG8lhFx4
RCdjb/mVXxDeYv+Dm3mTCknOLaPoUp/bpzjNEvMv/lS7NtdpT0zN1ueisR9LKvT2
ri3OvvgMVOilhHiPCA2Nbi9llOQslsVya2JUaoiTGiLgT6YBcrd8KznG1A8oHO70
o7ixYays+Gud4NUQxOXQGR7TdSIxmjVaVhjsfU7UP5rrwLaIPulYvtRQfP3wgJgS
yDhw76YN67vvJtvVbXEmHPD9awM6D7gFKMzJIaJQNRv9FUVf7FE3tWo0Ixn9VsSP
qVi9LEIb86NdVg5Yo6I26BbRtNleqGFPhKaqeJHHjYuvrFoPoI5O91qTmDnDrYdZ
9teW5QyCbK3JfvZ1/XfnTRDHRuS7//Zqxj9iB+IsC3qlvG5JUUjXZlqeKWQbWGET
ItQTr4BFO1Bv1AfnS4rTpniad5Zr1HCKC//mQpapADSPaIW+W4Qj04adBbyddpio
+0zhx6jzxA6i17cgGQUt5W5qnWM81Lw18bgy/a+vUNlgvC8hSPr91MTNQPR6Ckuf
Dsitozi2mP3YV3IUl78T5R98oQMNfjU6/oPVT+y6xIurB6UKe3Qv1uhLThfkOSkd
jB6wo18bdlJGtt25MKWNETDNOFOk7PfqeEmx5zLlQLhh0MEXFSKgtbjHQkf+A+/I
EE9SZxz0Fvc6H3hOcOrPUQuFJmi7zdC6bBGfVdVaUTjtangDFQjgzdrlzkyh31/l
Itmkiy+h0Szp7qkeP3odGfVtoxiC03LKpYso59LxbTlWiWkVJGW4jMlolVLQKdlk
/cH7Qn17SBho58K/Gn0USWYBZZipzU6vq6O+rvfi3xNlDu1LPP0LYSzdZaSgPS1j
BpJcPeHriKlj7dry6gcmAkVMhNyl4KLs2rUeVI21HkPeWkhgBb5TBIMRgmT6Kj18
CXAQOQGrsTifFU5TrIJQ6lU6x0D9en+M3pa1Pv5jab8VRIANejMxdT4m7bvulKas
KBt0R0h9lWFE+DyFzAbKSCdCi+9Sg8qcMiWRUU1EqJtjsHmz62hPj+n7ToVSM+hg
RUy2yNYAwSeFB8uqdCRwZ8bVXj/hId3z2LUNh95WFMhhqj0nJRzh0492boXZacax
BizMT0EF//RuRwyGyVIejdccNPrHh9fZZDBI6by8v1gH7nVEP7NAFw6OzFnxxC67
Us7bnMn6dbjQUaq4aenByu8P0hoD0VtvwgRB3rOPiyLy6DMezD6GEi0e6d59qi7y
nSOjNWWJn5t8DC2/k/djQn5qEThrR6kpP1mRKwMup2K5LtrPeSNxGbgcAiNJ2YNj
Ds9eGG796U0GRCXomLZjXL5BkeLK3wxZCqzRWfle+SmuPkL/CrpKZlwF+EjSN34V
UtN3kcl98tvoIko+dwgBa6hAqRNN4oicNY/T3+i+V0lTjtVYf/clNqqenYDCsgdf
9gOjdAAre7Q85Z2NQcMaFoEOASJPdbqoAmtqanq+52+VQZ6ph9G69osivBDy1mgM
dMEv0oiDYx5YyDws3dAA9oMHTODHnzKSHwXHXWB7gsgIVBYZ57W8BAc2B2adO887
wEp77/AXXlO+hYkp2X5KiZ9fK6azjCkkjH2j55YhWWctPK5h+Rg5Gl1HMTiMziOo
TOqe0cx99dTWpLWR6NFieOGAz8bT8U+A36lQLdz3ZDG5WeTQ30PWZ+KB/sukLNy3
7fKs+VrE7YkG4HCbETglBvGtq8MM/WSfynxH7HeDiAG1kPCRJ8lpZWZl26dmAhZ6
aZqXzR9YcNVEM93Ughs7rwtt2LkFf44pNld4mDGN9vFSaJ4qv9pGsAZksac9CwQN
IguU5YdckGDPcp+f4PgWzsctNmUCE4/Hy+ghtFW7fDTyHLHo+L0ytatVbfTuI2P+
pYxUekluz18HQQwvV5QRTmSECIE7xcFah/7gAZxZc63RhqhWGI43Oh6ELGgiSEdu
TKQR8IDqOPIgQekDMOvRFcZseTU6wbmpBgdEKt2mIgNfKmC7MP11o8qBaY5zi157
aH9iDfeooc8UlMSRJP9854L9TJqnGScW8hEfBIKF7KULUUdsPCyI/5aBary7+QvE
QREjwdP/iVJ+XjIPIj2xqrROLjnHtvMN6n2EuH5hjFxwGExTfK0NmxW5zmbCJWS/
ONRxCXeUIGNkvooyTogMDpzhClWhSAiYiWIbruRIMuIqyj6B1KAQHgx68HV74znW
3Dlic0sDM763BC8unSQm1tFUFoJrfdNdYqtWsvmX8bQVryooAKOyCcq8OvC0M5O4
bgyLVted+STbNXil3D0WSrWbiKP3z7cAlMwpr1eugWtmNT6024qhhVoV8sAXj9Y3
SfM/n3SIBi+oIKmZBGAwDdThJeFkrYkurzbc+hH6+zvtJOf/FzvtHaj+ls/dU+vE
AsMWFgF558Z88I8c/9uiKy3Ylqom9REjblcCNvTTdfB5JoEQSUeaWulv9nkbUZRM
kicBIRRd0ARnqiBeRC5kUY9VUkxYOsAtCXAKufMLJgvbBEI2NglnWCKBYb0VK+HU
fGJ5UhioPru4YOzD/uHIdyL0OfABrY3NtkcmXZKjd06p0wDFYuSIBbbblmCk73NB
nQZHvja5s3tofc2i2+p4DgvmIpPXUvJhawCYoFEo+oDA7U0MYcfsUzmDZTkVrngK
LBXUq7kxOwykWuqi79tTjG76wW2BUeUv7RxEBPt7L7RimfVJnfcYAcQs7zE6CJ9f
lDDWZM+0w8/TaF2+wmmPNnBp+Oa+hd9VYj8JCYnSdcPx6v+DOEXOmH6KBWch/YPt
GoVheulrM1NWeuDDz9A/6liDOoJZta4l7K+g0rzRg9eM8QF+2P/pwwS5HNhUmkYU
SNzwMZnUOkRUl5Iisg3raxR9AJay0AK6Lh65fxVjzexQlhHRle5Pfs4/B4cZqq6N
zD3ffjIr9y12wPphZamvMUZdJuBMpIlBknwNo/8tTg1znrbNyNxlxWU/olvh93/p
no/pk7XSDjdXlH0Sqh/VhonmYUmWphjUod9yb4dTsNkZSIv4V+hQWVAeQKEXVsD/
HrV94quZ6+6zFv7GVUB7Tk1iFDv9qsq+y4yM0tygrpgMpFoQTf9m1XGWLB4hd9EO
8qqwS/rsghWEo4wDUZoRiIUFK44K7h11KqP3zH+wuQdmPHQY5tDQ6Fx886YlNkjA
C/sOpI7+MnlAT/wOsJiJK+W1+yQu3zpDQq5mNdf+dHU3IYlZxCCgsfxAl/wpH6ZR
A2qVxXVeJe8KAzt/5oZj2iKvADAEFY3bMiRWz7mIzLtJe1G7ByuDjpyglcxrxC/n
OWFDPbn6YHtJ5QEUL1YvXrgyzxjW+C4+kG37dVbyEmjqwKc5VE2m2DOhy06qAuEm
AsRQwUsdt/a2y6pJjSMG9E/p6BCqQ4FdvUBsQTH9iwNjDbiOqbuMbjqo40AnqvTD
plbbmB1q6eY1FwJwczO58QjxlAUdbkpKo2A23SrpjppeTV4Ta3DIrH2/1QGIXPPj
xFVNv6eNWIPy+5Dv8mmSBI1aWdZ3P+23BCEakI/DyHVdRRxvWfbFiO6WO6oIx3Pg
vGAaCUGPURbqExfupiXeLQRM1w5ypXlH6a/I5gn2R480C6KTtdvaKjs49HKIgYn1
oYpr39bb/yPNdZ2u1zeczeXtJbW6GqiEUuh2CZDJPKrMyP1fv2ihVyXoOKDse5vc
hz/fk10PnrXnHj5yEg1FQ8ozBGupxCOdzQa5+5K5LHjnmahI/SsHpw17z8DJXd/P
+EbxZ9vglY46y+PAN52BH5KhRNZip5VHO3tyZN3RmB6wrFDVtEJz5I6qkuFJwl7E
0Vdf6X4SiY3wEhXLPOOFuvAU/OqwenKxrFUD/gtCjhPZvRRL92CVGs96M1/w52d7
Ny8UjUjd8Vfttk17RK+exWjvqCtCzlx6WQMDEhVxeC9DwBgQDLNAQI+6DdOdzkXi
NbE81S/IkiQYe/ZV8fdvo5SeZR8FWmOhTegVC7io2YnlxLPuH/9UPR+A8hKgKSdu
3ZN9yiMCJZ4UAuxsNBlRUooXarzMrycQsxmTwoyvanfusXNo7oyo8Xrz9r697B6f
CRD9ORmfjHwyJpYOBL7VfjPJQcQeMyPtXPpY2p+CNYxe5XSvbleXbJt+ghXn+T4/
GYmJE/hDPhbX+j65QK/ywc43kDQaUl03K7r63rG8bhNrPtDGY7gR2JQfZAC2/wLW
z9xXnwiXNxR/T1QFJMpsZl+yq68BPmiOxkK80OCrlaxwx6Ror27RJtR5ikv8rn2o
qwR6uXCBGmwWjiBuQlVPgZmsLBglmb6Jr3wAeOurSEhXr8YzToJ11FWQ/IpVGMZD
5UuCyasW3nwpMtCxw4UBX0nU2Tni2hQN7+jl4ULONaYjZhUn5FOEsbGEmej163sR
5ZIOAukpbG4MAV4OsfpF5H6a/oEGYM2CQqgOtoUD65j+98T5akEZxyYdAdLc/u4f
VMy5njXMqMoDlIX89ha/DPbuMK1yXtL0YGoRlj+mFl6OuYdsU1LGqhQOXq4PjUvy
xpZzYlL6hbNEMoYh37ENbJMK+nnmWosdAWIQSwfjrEgr7KVCNYQA/q3WXmXBeg0m
nS+QCfVCSfd+gt9gITmxV8ty6EJQvs2mCXGGCTXiw8uZDRyErqEbgPEtGgd0+iz+
5OW6l9X3l/ryHiRbK4LgQi/jjK7vEL02Fkz6A4hkshFXYnzaJZudyC3RHOWKeOgQ
fqMkSPyah2wLI8JKbiuA9RitFfH/kB4UIOcwOGPKxZnK9wAAtzX7KmTtEqFXxQwj
fU3jd+0XGyIpM26R6zHp5bM1Uwcz7dvnZ7wSQ7axGsFXDhP9Xa5iBzEJfEb41YLe
qgctUh3TzgRvkpYT++GMpDCbnJzHahQ8upEbWmPxFfYUoLZU7tX43euFSIJ+gw/8
3BRZeHlxC4rf2kyour7XX5j5FdvYkw41ko5j6ZcB84kadEg6q4Xk3dbaVaBgHBMO
aQr4jnL9q/ryqj8LIUqdTd3di9Q76iaIVhCft/nDTuzUhtrOpD9ZwOyr4EMzIFT2
ZU9p2K+6GKYYmJmj8G8lCT1ulwIbHM3yGKDHfZ1pkY5cX09zOGMzILCmw3ytmYLb
ghiEplpWxIwVE1cAc8V7dlwXHcGCbXLMVGA2Y3VZYJVNjAwXDKYIBwelXA30olJ7
U1QbcfRTPlhKhR8sJGbMQzDb21iZPPAU16oDBhkQNgOvDBI58rO06hDHujs/iMFT
za1tcsROMOXsWmyZu1Wq71yar9Dkw1rCWMnE3ydHh8K7kHqamuSFf5nVJ5bvlyGf
xFVNLKNLQatcZBAE483lkfGAI1Vx7/x1yb/RFCgdvvICF870ujrVRAX/6gPsEwF3
p2/6tNU3TpXo7+nWvKzaD/dYsA+wCNFNJk3F5A2C1lLYoLyQWI/Z0bmGCKyhrzK5
xZ0U/uxcgn309103722OdRBZQb0jIcfCilGzlAPqSwC5nuJgnrW4UYNXgoLmm+UY
4qoL0hDVlSVdId0DiG7SEyVORSQcF7yWmaOrkSW8sFI/t4NKS3JMk2qe+GRVED/Z
f1Gkm9vG0+bO7cv95iuI2nchtfpwzzdFnTHJ7pIwOea9kMh3oFyH1MFfkAze/cHp
X2ooShuMIVqUx3VJbGdW1nrXQPK5DbLXgHuGgtPYmb031s+gKqa9nb1qcbi6Gn8D
vfnPjN6knvlozMcSshCLDEvjCV7a9FYCZZ/+22iuWV2LvLmgDA3U7F7Mx5O5l1pR
1AiAI8MPUp5JFkAWHinem4JsYnTVDZiUYmwrywbgdK2bAoVuYY3KMdkSt2OrpkuI
gvaTBfoNXhcgdzz8NJAz8Qrkz92ZGgDl9UmZbNN3QDRpEiC44gmugEeCEPdDe8At
zatfwwYAOQUMP2QjoLCgzp8lFaH35A/t4kyW8ZcpmtQo2VymYDWER7VESrYkyBrN
8m3gvXPCh5sTAUtnLN61mYZ+/ZaXrdnVGkbTQ8n+dLwAXowHK4it9dFBV8Oy9gZD
UnlKIO7xkMHqoDNJWX1iVGloT2fCePuk8iiowJfLmjx0fjB+cNpl+BgAO2wdpzxs
/Inuhm0ldJRhkwOfWxbnTqPdIDV8Y4RY1/lkAUzBgoIs2hPM8Z9mL+c4xloqgwZa
tQlqO7JrNSaIKnsso3qBHUEjp55UElSIyLvoUJZYBhNJLcGmEERCfxf7hHNNLLzB
G+5fwiAwrSYB4oi0N3JsLzqrC/NvO+qPKMAJRXLbeVjxypUT9QE2Ynfb92/yMKra
m53KOpLjvKlKNSDXZvetlY0k3Avk1PqLR1m42Z/JFbxwFz1WQViMRe8PbZmXAoXk
jiPPUj9JN631WfxjnwsFq9XKk7XezRdOAFPni3ikV55E/Waaf0zi/Avn8XdcQXW7
Z81geYj0+QuBCe78VWpc0CCRr8RN5yFB/eaBEZ5IbTEBBZ0hF0tKqY3Cq3Umlprw
CJdjq6ArgyVBpAoBtxPGIR1Z82osopsaQuLtMt72eI4cXnapQLlGkcDWBXbpOuBV
IjuofhQ5FHZ/BtaKKbMzPUu8k0gfZzNUGOP9Eah/11aBtxYh9h1b7KoTOaVzZ2Z4
VoBFoxfC20Ge3Qq40xPCdsCpxZT14KYw4qogehFCavYOGoCglu87PS9cInAjZlVU
Xx2Aoqwr+xHWYNbqcqe2JId+N3lTBT5/iA07tbYGdtYYGJAeGk+kL7LiaDKvF/Wf
ReKswXq0nhurPHRbgqY0NGIC5fKEl15J4MW9Q74Dn0ZXnPLjQ9oWK1RvgCgHqZ2B
cPinMOtw8GnFn1h+v+8Dlw3anSbRjzXiWG+ziPpvIIJdAUorkRbai0KwxqKijSJ1
Rrb6i4CotBJoodvyJkWM1iFuN+HQBGKs6FnFcV0pogZEVQQs7yFvX4kSfJ0Bb0yi
3nTseC3XzQMn4Jah2xQqWr8wChOB1yqQC+WolnbutdRYQ1b+5i8zWLd6JUcBqxh1
iZtnXCpSWaUkuUTudAJx97SVGjBPP8wexAKtoSkUJIu38MSbpi9RyzQYI+QIBVNx
0B1iP4KqunCMZDWSfyMZezTbVJXjbfanB/tKpFLx+DT2p8uj1QNewzDmRw1nUlbE
SkO3rytKPLFyoO7/DrXkhi0BCvXmmUhSjG0SVELBlsziUCqWYv/JfdIRqO37aB/H
5Gbtaa8Tqv0u2A3d7Ahfy+MZWQZCXe7G/dwdyhQmiW01ZSJc2oGuiL6hAVye2qW5
lqhnJW2qnhVpPkhN9Nt1pijHSTqKoTY3zbnTFl92Vnf/5Ek/SrYNzjyD/8giw5Ni
qvRVBfTg1NByow9oEOpza8T3++qBRDmRU96EQwGxyB7Q8R1bGpTfI0Jl3JmWoGxu
/iTXDc1vXOplTF7A8oV5i4Iu/MQrsJ/T4h6vL2FO7t11WxuqcI+0wgWvB9LDXbGL
Am/l3sVcZBKgJj8oUbpJEfzHEW/gtHR5J6OVqTyq0aAEfxURDqmQVdFWfvmQU2nL
V6qKCyn4UzHNbAGtCqRPkXQZ77SuncMoJV1c1OC8gsVOfPQsV+v5sTwT+LXq/ECL
yqPuZCot9sFZaZJ6R924TCVv9cx7PtasJjf27RmZTMIwdQ3kWmiqD2BIHGeBckXm
7mH6EaIuQKtI6ZNmSgdsNslRRjNx9Q9URi0tGkCr8Xvi1IA8mfI7BLpEF9NNBi5s
CvGZURZAthu1Hz8nxO9DQ7W20uEulcq+Y2D06hcjHVFOkGyyapovc0To1HQbRl2D
avX0vDaWXnsUxdDgkwnaNvN9Z1RXSddHkjhfvL5+8glwlv6O0PVeibqMLewEeK6E
40nToC4mSV9KfSClpm9kznfZQo0aIfKefEi2YCUWuv5vTJ+29z80Xg5Db4gLfiHz
NTq2Bfnz3xLiSEwH3ux3RCE2UarJTFOyoAMs1qloBAd00/9tyo4D1aOVFXY5Qh9S
ug2Iah+G1Ya3ZnNkmPIYcPkZsPU5iCFKmROqg09exZpNQI3e4TrV4eSCt2y/um0J
jl7ayw6Dg+XZiBnm5CKaQH/UQf+8HB7M6E4v9QCNmxOp87c3avPkgTvovalDyZVO
RfL+i4WEu9JuihatVGBal0BcuZ9zn4OfuXJ7V9L7YNJy7PaG+SjJSQBPCDROH2Ks
B6j1E3D5pjaJXOHNrDO/2WA41CWqHr7TOOsd8zOt+9re6Q+oo43vivVlZWM7M1NQ
vw9VSUwjW6F6BAZ76eqjtw8bPSjolOSLAXP/64PA8u9BetHjgyX+QZctnSPp4GIH
9Ulom8oCCdB/nXYwnqBJ1mnFbZRVgtsMDB9Jnx/0eUXtC6H0fblJaRqb2FAMofob
8ARDZ0gTpBtNOJpUQSWuqo8BuTKfeooAZD95J0w1b1JHKvMnyfYyM66j6txj23e2
3ZWTt7cXIrbp06+NjJL1OaFE0Mct1Vcy8a4Zs0TZ3CYwcMfK0D7SWovpdMl2qs/V
Y1duwl4Ga1rEuRyRVsdQyYj+QGtdzxrqfJXyLCuJQs54T22YMGAk5BcB3YXogPHI
iqwyTIzss+BO/mCvTeDvXvVRIL4gG5AiPTWXlfHQ6rJZ1G439Fv2HcBf7kG7AicI
bCdvq8HYn4m+JKdy3qTmSQ85Zjy9ZT8wkbj4E8fJGvBd++ojXqj/zCBfxOQWtYTu
huhR2xkV1HIMxwh+tmLyOxRMB2T9A0P/hERFf7tOoSXjR9FfeKbb/HbC1+vjZrP1
8BhVTo0SS2yQI8vFoFVRNNzjH5UrLjSv9c/HzvkPnuXy5g2zNwz6b1Gogl980SzO
/GT5tXw3RoX2vN2xJpk9pbflJtJrBcNTts+sjMiGtzWXCvHxxfAujZa4PLb3w5gz
pYuQNyqWfjf5MMQ8LcIZHfmBB3nXgGwwxAgtTEL5yb0EixiC2Oxm6YgMUAiFdRgf
Al5/nRas9u78IrLiBIfbNZdY/ZzagEqv3cy1Ubha3l4eyT9eLeMcJBuhVP4D1G5t
tvY5e6yNexwGracWZixOynh+RTleztjsQq/JZUKXKf/vjcAamszSPGOUb4+sU4E8
Gwr8vIUD+mtJfMlLPWhqRj+mcMFPtwPQbFIrP9FvTQCurPHjp7hztgab1ZO63ZhB
9lEOLTz54bPNG/yE4UJYN0y2wXKV2T+mn0DBFlLhUoIVLHEokBTZ9A9GbJRklP45
0yTNHxOEPt4aoL+QsLtjunpZJ36aXrjafo982BMGWcuN/d/xxUTIXP6pZ3jiPkb8
eVXkz1u+TN4Q4giHIfxuH6xX8aoJ1ufXpk94dvrQ10zY2aLIwJriumr6CAhGFbTA
13SuHifoUXcpVT5bzf12572gTQqxfv/nssJVzM0kYLL7aZK65n7C5JYzze5UE540
+zn8Nep8nsM1ApgYQD4Q7GXAvdHx7xyJvJCAzS9OzU+aj3oV8gHYvgMp2JFPaeBH
NG1Ur1oOVvvO8iec4WGqBPkGE2dZIm17ZjBO3yLDOiEQtMvkodwDWDbvOJDRNYm/
Hhx6+r+YUo3j47LEbdf1d2XB2+L4exdmAyY960RzOFc5CBR2ynx3GfWJe2CC3EAl
VDwrPRQ/SsKqIEwIZPTyWcua+yqU1K2iF9Ru1umEp9178x7gxhGVcYIf+fIT61Fx
gthnz35qHTaMpssFnaEI6yMm0aP7yeG64+LjqnhWMePV/EUmpZxcimFvnnCBHE1/
moA4xQlGr8Z9apGYPumsTWLTq3h8HCQVcgi8y1R1zft19xiK3gvrVNEpMwR0Npsz
gaBmAI+pNuwLjsnyqBSTTVfjHvax/WFoNp5irLSm42an71Zu5ww1h2/EXnjbLIzY
JDQG2hjqcVP3PRNYhsRUxredZyfN9m0Qq3cAVWQU+vK63f0oEAGIMMeVppzJ4OA6
B35LsrKF1UZ2YPMxJ+mVSrbtXb5b89ifingOH4dv8UrqAKAKopuLSHQH2IAREZ0a
`pragma protect end_protected
