// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jaLrlFHqIlyrCmN9to4S4viYgyQz1A2+w6n4Vhgr/RENT65upXA1L/SF+fRy0xi5
lD57EhOZe7nP2yrH7xxjX18lGv4P8CIkCgDKuPtQ82yKkgETXHeVttTZeN9uhUb+
fH9yLU/6n8GCAuVdR85mIEnX+VovXrIBaepj2ts1SB4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6432)
Euuvm9J0Z1RAbqm/TLShUSjvbXgtp7gwKUzWyd7tiRIMUTdtqcXkun0F/jXLZ4bp
c0ZYeM/Azuxh7EaXY5KfrOrdN18zs2inmo2K4IOu1cgqpP9AZP2FDhehxL7HErWQ
uQkWnuyM0NwJ+BOeZy6Nch9ayUNukI/muFs77rjDMif+kfJZtHux+CGiGecLH5hS
NnQFkyVPxiMYttb7BP86H0NMEzeV1Gnx8lDOU5h2dBQcMV3E6gdpBNZRl6GPgWBR
Qnoo3DkYFYgH7xekBVamncbqsfMGQuDBXq7XWgozWVUaLXm6gKrIA5TJVBv7Z7A3
KhwsWTHrfQlXir5gaLKExicMhSsRyXl5U3O4R0bGX4/MLewIx6C5nHDjGx7InmjP
+SwuSl7X+j8SsVHJz8CWwHNslgD1ZPEedNVGbhRtG3bmaX6n8bHdyiVE1ne82DU2
nj4g+uYqmddotbiEYjYW2JoMfxfhmCEJvwEzyjS//msTtpZxweTrP14+rnEBJ4D7
pzck37Ldpj31MxoS6wxE69LNe3WHsdFJ3dp8monQ3rYU3mqQl2WJ7bDmih9vTto9
0CxNJsN3NXpKR4lWeRHRZszIbmln+h8KZIYfRUptyjAs5OHUNJDXh/6+NxiPHkVA
OcgTK5vc1XAAHRuVPOywWJ9Y8PMRR7hzs2bpWuwMl/hj4Elz2JBUNzuzQlfsNRYY
QLMo0KcN/49UFMSH0XM8k3oGr90f6GK0bQRalIeXEFvUfyIPXaLgSSM8Yxlq1BEn
xQBiPzddzp+m5c/SMioKlRCNiDqfZ14brP2Bj2PMG04AcSIlbK44Qw4cb1E7x89v
C1vf2xg8dnH+c2CQ4YOPNmH3+lJg2qohnD8UUt7rJjvrBeqZjNnG5SpdrGrUlKfn
QbvgUhNbMbcVMdAfKWuLG8zP6+xp1j7wMqosWTrEKpPQJnRqy4mdqmKw5sulLo2K
Iy/pLP4ApHWl72NBU7sq5fYfS3PND45Od+2A9OQr/fHt63A1fKZSZMEyXu+gTJOH
f3IhGvlcwHkVnsThOW7zewH6/r/vKrg7q23Ru0NUuK7iBndbzl5YTp3uHr2WteHv
q3JNPsJ4JWYce3P2SGnuQ/cjPp6QyhwLLmorRgQE+e1Jefr7OqJN8Z7/xJ8D6GYf
VT1BbX2SA0sWDqrtKQ/ZX+34TxZXGuOi0o2JHxJn+Rv8ZhyI2KObvJqKPldrM+NZ
vK7pYFlDtIzgblsN6zRuG2PT9eXUFXwEYOvjkVX6/9VkmxvJ/ICw/zyPdH/jdA2C
SLtE9YxlyiYz51GG2+fQ4KR778IOB9PKeMr6h7/UtY9W/6JBxQ0tX7kzcbHGDaJN
hzca9+FsGy6R+uxpqO+Sfg7tARWOSdCxY/TpogLLexqIRq8VSg6Xexq/+RU/4Dk5
j48dNadqNbkGIAJRE7vay5S1/duJoH7KTg1at08MuD4RbqmR2loAO3bZRFc1G4AT
Ri7g7MpolWHWDg+BnJYywIvRrydeglVNc+TwUUrXL+le3HSiriawow31BTwtiT64
ARBAppEOHl8mrM8xw7dzuoCNY+wsfMUZWP7CBgZL8nGExJxYx6i6+aV1OtRJF2GB
5DNBoBB62+0RhTu8Qclvjv0Jr5fP2ULiXLBuc8PQ9fhhHiPFvRtPiqUFlhmnpYpv
P3Sz+1MLjAmVpzANYU04GIdvfjqyoy3Yong4me5BgcFZWFXdhh7Rkbm14zS8XNJh
8mZjvIiDdPnWOPUIvmPpAR+TXEB9eWGGTvtchStzuU0LD7OIP9MbAs9dXVHNaQno
ujNGyYtg/GeS3AhlsAuEAXN3quikesLRRUvey6aXsLDxYiUnHDk38bsMS7+l1mN0
oZl/tGYmrmRDY0lYnXmIsI/7Owl1blGUsKCccjzmDBSgxZeVd1n1VshRjKjGAWV4
hfhrhv4yNPLgsQkRDQHhgIR41l5Rh3cxtk8DLdk/v1NSihAcHMHk6DO5H83iFhvA
9MLcfHNSXyTA+N9GouylYp0fnGKxUFY9siq3ceMPjHJT/od0N7X3MT2HsI8AUDMh
X/9lb7Dtwr6WQp1Hyeh6G9CBjajkJXAnG/oxYcDKCm9L6f5e5v1yCtutbRGSjEsm
ICMIEKB7S+ytId3UKHJQUhQlYJc0bbG793cQQ9jFS/jCISXrybq0rQhY4xhbbQKG
l3M7xIpnMsEXPU1pPnKoEiLzXQSfymPoEHY72wEtYX5SOg6tWSRnIVPBf+htSBNP
uHULi+it+ayl+7Uh49fYYDXJN4Eg26nV3L1lZDtSEuz8LNeEVv5nlVceFvbqJFND
hkrYfsVRZdo3x5ccFp6V+wncu/4ugfiNlpvLki+XExiP5UXcIYmP4Y3hujr+bEsa
hhPjjrR+sm7yJpOcLQWVm1Dqr4QwWOUq8uEof0CNfFTxAGcXvjpjQa+3k9WEQ0RB
i3YvS/nKf8ImIprHnSpzn7S0xQ4qiusR12QL8rseQFgSih6aH6Duc23s9+dV+GDi
hEImn/DwReZtDrRSxmAGcZHWshz6K2XDkK0G64KFKcrJBVi5MtoKJNCJopQUdmGF
lTgBukkSViKb0Kd7Pg1D+/rQsq65snslJ7mH8t/cmm2X2T14KAlTsCXgDSQYqaTd
8Ewm6fqf4KPnKdetTa9hFNQzq2johzQYWxLxfUAWiwp9NZ4SCPBiw3jBB7NzaJLh
+PYLFUyd32xAjqM/aayAlA4+z/om0VqXZTHX5nz67E7OV3tUCvmVMpOXqAv/DhC5
GFSzVdtrE3Jm0r98dolWPP6uiI8wwCmCDZN8n6JZLOrYAu4CI3P/URKLVLSrCjBb
vK0UP7yoDk07Pnw/usWv82Wxc8HtUZTwFAQLomHBbUyVQyaE/eTSBs85yfuaSViT
ojij341Mnh4n0/fu6W8HKvnhb01KavNK9/hm+qJiDCVcfRDLfC+oVMDBkgkDZ038
al6zZSvMNmEsrGFJiDtgnF8PtjKgBN+OBWTv/MOTJ4QlwX0XGDc7pkNARk/MFl9/
PjwPziLpUVd5sQQTMagtvjFg8mylv2XVbSuLY4qy52B/+O5hGMm8QE1qxIvNSSMA
9hJvMDB12UBbJ6mvQSsIUnu0cj65pKzxJi36CFxTQUZIb70E6J6TUoJh5UCcuayt
hz4Oo7Tp4g2BYool+/qNwSrVjMSjdRGrFA2jI4IWCwMM7apvZzjdtN4LvpnPNFXr
PqE4Xl4s+bN3fenpgQxrbbb6KSk1I6sGi9RJsu+CPSw3u7FHU5o4Iwur6si55Wr7
619XM9/SwwQG1/cVE3mrhLbaw+u3X/mv9PcnSvsHyd8Hy/nEF0c10Dd8E37Xz0T5
C6eRGe0fOOL4y7SmWKt+SD1cZE7Uag9aCQb/Qnw6XC/XnCMEUeMC+KMPOVMQenfs
xlV9vMuxNH8jSPHv2+s31UHxYVtAbN3hWjV76c0xIkPoq/ZeiIfUD2x3XBY8LVs+
LJdPkL5VzG0KuVb6L9AsLGqKAYr2TGsiVQVzW46IYWAMYe5A3zGR+SECQ5ygU1lR
SnPq0CttLwJ3+3qyi/7TA3/Zl1jOkb8n0zp2ATEFwhS7YMrREKh864osFGPx6sra
klfsGAZlc8JNOCZZylNhtrc/8LkR286cYS343QG7cdwdy1LBotdxGZuhJNcMtWg7
IhZWVI7JWUJ/tu3SRNHsDGkzIzY/uh5pWiiyR8DfoBqTu5edb/cX4mNCr3+XtG8B
zR+AzSx0SQ5Tx+PDhjL1Q6iDWjPIP8I0NTIccVuD7ZL15sX6CfpP/+I5Rm0sgeIv
IAiZoPMKqZGMR7yaO1skJkZO7SnTGfOvHJtZT/45usZJuWQaCv59Ce1qsOORkqT9
kfhf9dBPTrCKStaK+UxtwwFby6fvNSWSs/bCUkzvcQlAqYWqJOWkjzHK3ULntDIM
EoCiB84nfRF4v+o1HKBfuM5nJoTfiO2kGGS8JnBtnLqhWbsT1FlsP/hzp96Wl2X4
/eVTzuVuOnAyNbM/d7flDNJY2Ex7NUrDIRAYoEQdPQApfjPSGM0mvVLyVAMBcdui
EJYhPdGlvCGM/CzeNBfI45/EBYkY15y6Oq0xJcAYtS83Uv8TBymSVBmwWsi2tZmn
DeGynf9Xl+7eVr7a15OR/7O1aTcoJErNLzDQk7UuUX25Ew+Vx8A4SCgkKpPNooMu
sKAAsbgcEBc798y0CfYyRf5YhI1+eZRLbXHCpEdsEsgcdAm0y5AoJvoTcASjhMeJ
Z0DnOPd+tEROX98+HnPebJdSYKgrc2cDeDn/uLznlJn9/ivSGLRFxdbzuV0mwV2n
uoPuhJGzH26xRgtRkR/765jaSLlVFO3Pfe/OUm8wl1ObauwVxlT37qEt16PsqYZx
ubadWHy9NigFCefzpzeZUuo9/V3mQICml6fZKogCEDvGyUd++garzoopXbVPjzHQ
lYTY3U6zJsMHDXOhtyeVl0Udw5DYFNuuckowr/fF3FSBfz11FuzRk+3rT663Nt85
7ns6ARdY3b/0mkfBueK9M9HmCyUmERXFYYmAeqKipZed8/9q6zQjp8j2lzNhM9Qj
DQ3BCtllN5qJ3lV+dg7BH4jBpECc9aWv/4Nt7D7RxCn7Voe+pKJY5zhxnmu3t5a5
9gMFMkEpvBDikynEftcxU3uUDg1DdzEvI9k9GZTBSNw1sFKRIqY7xvc8f6eF/Ou2
iALTHXTI93PBT8AHG6lJpcALPdkWMu5c7DFXznTmrawQsqOXOEseI8nGASyqUWKJ
ttkPEVsqeDCAFQkFcWSRwy+FePkXQunbi/q3hA1kq1KubLFf3SgYPedId5/Tm6Pd
2mHFRO21WHV8CKCG1v/75d5SZrk669G9ZFMbGCASCpQl3BRBE2ZxD4sKWCh+mLeO
/8iJ0Yvwnf+/z+XlzbcS9BNtecoGFCZyKhhyBsFjcRR9gKeGKWL0GnO+Q67CR0lx
weO9v8sUnGSCzoa4ePLBZVkdoGNHodxJMgWlAjh/DfR2V0eKGmTTPBhwrB5ybkWu
9sYqjNM5vH4VNsLggf7oBPRUFx3V5gmvVh0Dru9MFsrB2poefZxQGuWNTajo17T8
xG2ZQ6aivmdIofUpED620HFq7AgpXaVNbAvk726gzlpGgRaXoCIRrNJLdY9WhotA
xASUJJX83StcRLUMj8Ifedieptu7wwugIipBzz0AYo+BiRf3XegjhbEgp7Ik7Ycw
f2nfNYTALW5jBTpR7MKDbVpB1C2O4DJTJSMIa83WEVKtaV6MvFXbgkH7rIpCkvq6
gurYPRDZq0Qe+lcTSi498e1WcrNDTJ+ek1J0d2reYIe+XRfV0WygSmf9h7l98ZJd
xX50/B1go+EH60x1EZRDnkURjCzuMPGgCxiAenQsU+qJjSasA1NURJwWrdMxXFE3
lMOQQlFC93AnuZ99On8MbPWeQW49umipho0SUZUqOrpNFOMKj846i5Wonw/i3pC7
QHQmJBq1b1X00a/MdTJCyQUUGhqcdJ3PU9uqC4Osx9QYT5PdBKsF2ZMEWoYaxQHt
ZeqXznGUrkz+5HklkHzFFtyaa3+aF/65ctKB+0ImV1yZpXW9BOMCoNJKE3huPWrJ
Ci3z72xriLShjmi8ExdvSrYsHm8vvXlk/RjnIn2YDSpaYidqFAoUJqSdb/tk9y8N
YfMN7XXjtMMTluJMtbLXzInmgjSxvB/WuCzF4Q+tbDT81YRjh7yIHfluC+D+tfKQ
TfGR9CXDwczmJLRCR1fvMZn4ycakw79lCKu1EPpb/tA3bvY+28e5cYqtHQdRnBNf
MXCOUkxiyUlJ/xn/i2DwH0F8qL34LQiRlahvZDeJKaTFqnfa+tY+VEH2Y+vnIGUo
7sEc6xRfnBI6UHKA0EZXoytVZ8gynT5FrrHfg0SU88t/DNWU+/Iulzgsect+gDz9
zcI4ljgnYXaV1HcgKvSPlxPsM/7OIj1Ty8uxWfruXXtkJ4Rjg04LeIe30pIpoYk4
TfnGtQZuOX3ytXLwjpLaMAxmSdBwz0M6SzrehLE9wzJ65/9tbhm72hy0G95lj61x
lKe/9kSJBG1d5FEZB3f55P3rn4rIXleuP3TpxLhVbKEOvXQ9PBrIcUQzpBzhewox
h0xHX5ixZrJbfUYHCMiL27529ldHNAWJQBsz3k193EwRjQS0Fx6AtjvMRa5x8Kut
c3PgxgZt7utbWvBZT8T+8A4A/3IOT9bgeWwD4lEFwnBT0Bl5cb7sSMT+jGNCQVfS
95pqo3j5/MOuxtT8fq3QPE1WokkrcBandMK5V6XSEXeMf+D2uN9LMAMf0tW9iDid
XwH/3GhYJ8oKygGpiNEsS+6eybGVyPi0geCkeQANLqE84fQUCjG5iNo/T1Aypl3X
8ett3+GbiVGr7+Lr5PhrOGyoredzxro4oZBwB5dY5OnPMq0sFC+TdG0gIfVGMLKd
gesDwdBOeewQaHThqO1fP3o1tfAiXp3qTHA5bpjmXyDXjAKmk/73dvqCUfVrK2Q2
5+F06xuAtdnOzdrGSB5tQbNhN1AiQgQi2TDNz18UGQBYhhPhz/nEbTpm4hVETO8U
FK1C77gDCcVnU9wVJrrYhTP+nLHlKicnfXtQb7twSTs6DjvrRdx4pibE+YLjW1h8
qM8wOOFMDFr7QLYiKpC4xoSK04ETXSPU7t9vh1Emf9W9N2U/Vnqh+FlKBCHFU5U6
2606X8DyG0ksDLJXxkp6aul6dmvX8jBMGzdfbL7adsQolTX1+Wz26nz9nH9m8U1l
TAawdr+m1A5jUo54rEpjhJQrStwmvwyyVTKo/HUXa2tgsxz69UP4NeJ6NpZulCtm
R5mDyTz4uRC1zXJGfq4tdWCDu8J8lbYe7BRKQHv57LQ15gAy6MxCrMoDefbPEbAN
sLbfFFhufJh+LfAAaxKuRVxw3hFCbNaMT6FEcjNoIR5kj/37XoGqHxcUnJ57FtQH
HCIY6sNT1slDvTYHDkRdShX381p7Q/rnP/c40FZPWedzhum27qgVpFFyN76G4uo0
l46iQT1VLZNt0RsLZCYXoOZp8WqjaOFl5AkY+Lqi95JULB7Sh4fBxKp+6LXf9sod
ljA/OAMF/eKTDJjsJXasloxNthQSs9F2lLaYuzO3Ncwh4fFvjC4Rv8x9evN9dDFj
tNq/rgutMo1vNh+4EH0T3wWIyWWrZT3WWJkk+y9RpF8fc+UPcLqPPu0L0sBHmWFd
CzfMv8huDK/bMSp8fYqHSia8vhhVkDdahN2SMboygec9aSDmXu2Q52lDcViVl/5t
f5bqWXOJNi54O8QVmPUsVkWgkURlj3SmGDpO8Dg8pouiQx4XYJTI+8R5RcmA/c8b
ax8VNcofa9lg8YKWoQFBOoliInmamwY5+QKFM++Y5gb/Sx7trNZRom5S4qy3PFBo
JoJp/7CMAY7v/bkg9lf0vlnoKBo+e8MlYp2Zjh95Rhrce6fOTh3M7A4BlSZNMucq
FwNxWbXsHvn7/ORqsEGhuNS265eyUvh5SrueRSpPbEdzXMAv5Wrf2dUdn5v8jGsn
azntUIzEpNb6qKEdOnqU/ctuYWz+qPD0tRnHty5fsxqHJyrZBcpjaPUCeZHTaHm9
qyijb2RbeDZE03covaOVM0/87XsKxtXqg8UEkr8DRxhdrxBlOIzzh+9FiuNskDrb
dWHAHDMTZM+8iA7PBkMdOwnvvpXuvIid3wE0denJIjcHzM+jQ+p7Bbp1EYGDmjzp
YrxOEZOaBmzWmMwpsxY4bceCagFrt2z2T1qsQ0gXKdDd0LihiUsZrAOusY4k7ecY
wNpfOrIfC8obCkxR41Fc7aX/4Meko4LNs+QOV5oVD/ozY2I1b3gYXJSpFKyZ3c4K
pieXgH13R46w4dDKf601cjDvQztq8AKv/jDAWKleTSGeXMYaMMovpnuS28GgdG/1
lqjOWNohu2Ge0Z7iw2KiDF6CCyTq0n3EaYBhvG4Kjzf+oThqm0D4GTmqTEwNILaA
0iDP80pS0iPW6rXIWhu+MiLARCO1mOyFujpN5I4gso8ejNXQVZk66+AybJwzsAt/
eg1AW9vZzCuvt4uomLfckyAFYGeY7A83QNQkhbfxTwGWh57HElhwj36M+v57c+7F
XnCcLgLB3oBtUdafIyTYwFgPrzMUeN2oBG4IxN36QFmiG2JucOA1cLO+VMRJDKqU
3UQCVpZFZv450GJtcNg5d9KC8Mpa66bujkwYdozGAN0+wBCb9e5gwCnldFNkFOVu
XIC4Ib+XOUqf8vb4c54iAxmKfkxnlI5z8Irm5qaeSJhuAgelvyZqrfUp/fNNpVMO
SZQmwg1LjT/7gbBI64R8ShRyW6oX8G1hjR1nNZe5Tj/1vphjK/bjydklmhwAj2Lq
FebVGWiVFTjzRCgdZwaHR3ab33WO8QvuqsBvnD8Hn755OByPcRPURauS02Nyu22q
gBmnhBVb/VRQAdL565C3I/XbpHKD6u/SON0KwaHYxAYgOTM0q5wQLKJwSdof2urg
8Jm/eodLMwgrR2Zel7s1h20qHKMstPaAsUm/e4go4FZ/sqnMsqFatg01vG+BiQ5a
zKzDw3aB3fQ8WsVEooYpgGka7h/MGyepHm6QJmQ2/DuLd5/mZ1FDZMaRq20D6fhe
`pragma protect end_protected
