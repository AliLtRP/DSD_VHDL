// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EQJD20Pk0ln1GoEI4cejcbo50kOMqtQEbxMPEM8VKbJ1PJBowPIdr1tQTF0pWpfA
ynCf12dyJtNwPnPqq6XY8AJ6avDFy9h/Sdg3e5Bq3S83FTMDvTPCz7BrKSnrsaV1
jAqIf6uf20C9zLJTgrFolkoqLINjJ3jPHkwdnyBLk6E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3904)
65JAtiI4irluR5tvXFn6/Aa2d8MYz72ZeUmMsKtpOqPS7yE9mbpAuqOu57jnGx+l
+jdoYgddbe3laIIzMKbb598GsolaHYpJCNQTh3zuGPFfxP1vQjP+CXR3FDBQOna8
Cyj5PtLgeJne6QWpm8d5oVg7tYZ702x5FMY89Jwem6o18X4FsJ8ofoCLP8QLgwcA
aj4CVfwHcc5FgNcjD0XB7K7YIFtOGImjN9k6T2OzmW+62bjW8WpL8QjwHqWl9B9Y
5rN3MPb+kvK6dOgdE55ekR8g/c2H5+MM2hhvzoa93nvVsGj/8TDqlkJHX8hNtx1j
Ha/YK7ZAZEbydtvOfARVjEBVX7Tm12ZtKO8MFY3nsV7bOetmu2GlSxwwCq7hfCo9
tET22/DjSDVdfBl9jeo+d8+OUSlS5x3s+4jqfYtQcG2MQJUMD/AvMnlUz5FrNJeJ
Ch5GINz1+tQjpVxxyp7CSO6wPM8akYOAxM45Vlt1SLaHQ/dXgtHRCKszZU3iif65
LKg1bH0LNGVYu48Ebd3B2v04XiSjJit2i6rF9obcl5xIHFIrkpjQeJAfqCEUqzcI
JNxvkUOF9Is4rJpHQsI4r/N7xUB3vZk1tvcqyOTFThYRqitLzUnqvdNpzpL9y+Cr
tYvLKXGlHc/pVxRbNm9QyrzrCRIo8sXY4msUU4S7c5gY/ivGnNMjdN0LPR9ytRl6
JPb33Kg7PFqng+WIiiTVn4WZp/Kt4+Di7zZWCvkMY2NUBKl989aj8ShzeD1qJG6c
m+/ACOYeW+zgmwrhGUV6Br4j9hyFgKmj2nNpPCUejBX0pFlvTAF8N4/Mr7jcSuVG
9BcWowx2U1K6DUDaDhp5BnLxH1dKSMMAMpXuR8xVlQT4tx+3hKbG9YWnRD4TJ3L1
uDhlC62mlCbVjXrRDUWGcXQHqcLM+fNCpl9QamCdkdUPgIaCVlG7DeWT2SFOkcEM
HXeubuC3G1A4yjYJQVqHTbYVHLBfJTFIAQz7nhXwMb88vDgc8ZKQsyX2iWGpb0xY
lQnapVTKA0PMTrWRL5JxsBm5S1ry+FaKpc6La+QedLGN8szzhr5h3HlCFXVSWI3E
S/GfIn6Uc9n9lqgmynYQ4KRjivpjn/ofR0t+6CJh1HSk+TMQYyuxZWhwiNLAyrNj
2NHl7kckRyVC6SqmOE9losesX4SjVVHSP2odx2w/w4CEG6aWXZZ4ZIY5xFftzTkv
v+zYj6ulJIXKebNcBtSv4QoahlXl9aMN+D5nwTAkP7vQq6vH1bxKMBMCxJCYx7HH
/nyXQouao0ln+konr9kmbHrJQkS4jzp/jLwpz8Eqguwn+IEodQBH6ce50ebLTBwN
lfABMIlG3WD0CT/kepiTLFhqNa7b6WG10N3fHz2to4nFlygLXOh1h20LP7MOqK2Q
P6vQs9afzuJoxJGwdX1aEKlO1Vja40pUK/iU+Z3ij2EEr4387QCsaXg6sb0tnn/u
PRI2Vf5bJJs3YrAhxYJ4WI28PUGXyB9VgddH5oX49VMcUVIFcTul9ZF/lap8jeTF
tT+xQDiHBJGOs7+qWtduxX2lyO/gxES2SrmbSeYLjXPA2zyXkJ5MTCCItrJXxrPv
z+IaN94J8ikT6fbntVxSfDKsf9uHROQGQIUNNaxJWzIa8voOOGn5vanazwduUNeI
XD4iMLrxQkEKtHU7t9+5x/cQOoYQGNvgNcSnU4sRAnwjVfFbOlJiPXGkV7RCIgXC
5j45CtyBEcPYX7Ei1cguZW3AcQX4JN1rTrod4vQWHBP5IGd7dmzyIabe5TGsFlHY
zdyKicVWFmseeJgRPSCbD7EOX7JeRdXvcACIwFrCiiRHTM/zbltbfkH2PY18VtLB
eAp4kqb2ZwDzEE68xIq2MIDPoX8C2gzwwffL1wNeryrVs6crPNiSZY6DsmesNu4V
h1UY9XJ9boq65bYPouASaHcYiLbFKgW0F6+uAF82dxEZfivwnBEU4wDmto2h3n50
Jc12F7HIzYjv7PzAnquJv+e/DNj/B/4vftsnsT9CpL3DzXcBrhv7b6w7/7fY0xkb
1URaofqZvsb2r94PdOabmi9wOKo7gzy2Y7t6TrW1lRk9WcpAyekBUd53YdR6VdYa
fVcLgz8gZxPOcDGTVcFRSG3hlWnCCDeo7Vjq/Wtg4k3k4NpwPw3m4gQnqXjuEV9I
1f47I6aaRDM9ORwdI3uFFLt5mvBfrL42jPsPg7fgOW6PsOBfHtZVfl+6DE+dgQ5F
W2c450IKlv1/kfJIwasVpG+m84/kOnba9It7b01eQO1Zq9EvqBxgTM37m0uxCkjL
gEexGtUN+vBdjY5nilPrV9TaSXUFVRxbiC/ZgagIxODF8KKVwXCQdwRLfSpWSkww
hQ9mcdLc5HeKKXEsYN0hDMVGAZHfZWLXEyo8QYut80KlCjXABJvniAJRoraYgLml
mvBvDF8Ceur7oIzoMLXChNneRmopihAdwjV8Ztza5ByeElRXBNgwWJHnEBMZ6jHs
8IyHVzbtYwOXEzYLRdW2S7prdXxonHoYnGT82xgUwlqWhDaCpffWc8Or1UHsaUMj
K4sqCDQ1u3smYO0KBR0MB9xjnPFQf4TynCPbEL9ZpFr0LRHYE9Yq7bXRVY4OIK7r
H1VSAUboyK9e8H+cfNnpaLPzDD3El0DWeYYYofAQj4iauB8MulSFkJ6xuTWGFlay
H+hfdz1I+HsI3yktIF+uSWMZ0yDzgevSdXWj0Of0xloBKISaLohS1TMcW6RXbOmz
JclLratFRlaWVxG8r7kqjPJ2iMKwjq6uQuYuSAqb+efgRD464YkHUBL/MluxlS4e
3nvgZ2nSqKw9cibZ+H0nL1E+xD+n28O35NEfKuU0dMwggDeZs3xU3xo5G+bYOmdf
m/8awgFWtZUmuBMtadovhEYr6m9EKDtPdNm1XvXscMIWxB6yPp80JApIgtTGiR5K
goNBE3g3Tj5zfbc4MagK1ZKUiwzX05XN7c/rv5TMRsdkpJj6lQjkLSbBK/kOim6q
lCBjzo15iYbVKzYrDQWxWYHz339s5DXAChDmRH74TMHI56T23G67JxYvuoIwP90Q
zR09fGMvY1RWH+nV2cQDStC6fjHpOegbmGM0w8IWq1jYY24z6BkfFHmr4kzTk4bO
tPoiMM+Im1vC7GE9c3sJ0aVVVnjBDF+QAG8hKmf2yxitV70Knyp+Yu5MYzQ7TTQ7
OgXqIA0CvMQCYrRrc8VlGPDMdR36L6dyHX7a/fTFAVOvtZKA9wV5MuAHiT2XK/04
p5hdPc61EptkSlN3Nr06qfZmWq2qTeHrDDxH5My6op8VXW6yqS5wdMxhTVoARWN4
/16IWWJ4Vxo2qRN7ga6kOQNfgPqKsulsgc16onlbLM3HRqJc2Zz+GTx6NnswG2Zh
V/YnWEK3iiVLciDXCKfde3SjZLKEIYnjSrrCol1FxGQRqrX1nPVhDxORJfEbDNgH
lIvosJaUvoic39S9UiHCaNQRusP/yesHBrGSmQtzGtzNd9Ykus+XdASgtpku4o8y
SKRo69JVNzR7TcA1jNO8fJdxQTLM40aCZBdrUwRmgSMOFepM1rZq8cnWrOU2nrCl
2lB6TIIz0Ptx5RZwqHJTEB5GXF4uwEisssC15sY1tQcL5DRqtAk2zrrx8PDGTbFT
ogrD4tl0p0WWaQv5ZRL9QL/KmH+/lbnFsBUpjdcVLfdemSY0W287130X8t5OAqaJ
4TJU8/oa7/gPKzTLB53aHXvvu+qm5apZ5L9FSjnkJPB1j8XtQPgwgf+j1LOaEx6K
2Z47w1a82C0qTFX9z/PNP3HDBM/c2HW2K5PVJnI63oHUqckU593dMtG23Bl+7kjn
NgeJ6Vc2a0/KofVZZA+n2ROhOUOdJR2qsezhaBGz3rv8pYHs/DqujKeaPPSg5ubX
u0Os7/PBLKWENiyTcm1uzESKWOJNRI0t+s8rz3wkQj5/bD4Gh2VQTNTZS8AZ/Q3q
/edm/ZRIkpWhrEcEgvGACp72W44Hij9dV63XxJET8W3s5atLqCv0Ibe9hajrR0J4
v2JAS5MLwc/OXmSgMx1t2JaxDO0Bwr6AltnVHUtwMjIYlYRBOtppdJm8X87SRz4F
XqHBLzL6hXBHYgc52RnciAJZw5xoDG0ooKuJfnQAsnZypVM92DaZeYge1IcCXfFY
Z8kYBuGjAoFH7q0ARyXZQiEtCnC16+y9OXBVs817IgRf1rv8IHuXOdf5liAza30t
c5ZKfsiOkZSM+YZ14W9JrbNmoOc+2uKg8lfhCUc4X2D2SvL6fFK3hTm5CCWGDSwe
/BVm3zWKWRQYz5g/VFp+k+Z12rxzqdnF8ngE4JWbiO6iFYFn7PtfkD6LqwP3RZVq
+/i2iv64SAPw5drDdMIqNhTrejXiB8V5xe0pfx/B2wLd705DZ441FIlqTtCL7nNo
EgdQjAvPGFJCGdkvp9XixBKcSu8LCBMYAPnoeliuJ/Q3CkQXaLAZsaPZN+DxhqJs
aSYr7QzQVUVO6Dk/CQNT/pXXUeWfPDq4hlUUVBxQM0jluVMFND7snVLQqfu2o4ik
dDQVXGHFqL6MBYy3jSMTcSyu0/FDxxiqoXdLFP37m44mfIaeUXNvAXbDJpRln8Yq
3goWFB/r3Z09EIctH7K4Ul66E5spTmXhwjkmGynRSZRwCHP7FiSQOwjsdhJ+eKhy
hNXDPT8iwS4jm6+unhE42X36iIaNOA+0FPU3JKTOTA0HV30atbxMnkZUSlDHKQrw
xlP+pslat6K+8qORngHKANpx8Ypcx+pu8dQ/FlBsnlM6vFEO69zNn3XV1hJaSvl1
bKm022XrG5UOuBR9bWkAO/EU4Hgq8BqfHOlc0oMtzjWbDNBo7zvpnzPmWvFL0OCn
rarhrSifDlsfpyDl9rAG9kcRlFrGJEgFuuV1B8LyHnAmZIIh3esTqgSq/AzhPmwU
O6SUISHda9/wNcASrZ8402ccBpeoCaNRln7/jbU2Wo1J89nE1IOXcc1N5KuEZEvI
k/Z1qJiEOzbsgXnoE4eiUn9Awb+m6Zcysgw8+8bp/q6qCID32JeBGEtypzJ7FshQ
fkLz8G3/W+qkox7TQuQykOtlgqNRtuxlUFrFUrEe9qcowBrvEcik7a2Oo1UoYkXo
0xjSjPA5K3xUI+NVF6LCm6rSce0QIKyVzcTxQElXUSdsB9K115XALnoA8An4Bpe+
Md/Q425t3CasdzhkzSyEXg==
`pragma protect end_protected
