// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Q0IzNGRKyShLhJGbsI4TojHR/ATkiEZSQEgwX356eMwZu+AbV3YdkxuMAR1UsI4N
upwGa1wJTVaqCha4/Id8yPI53YlJqqqs4/F55JJKc0eq0kjzHOl8xw/BcLTHBfDw
y+ZqA8UJJsXawg415/OT1xWRs64iC+C5CafWzwbQEBw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12912)
QzIRtO7DS0EtP1emsro/nr7iN9YpqyMQREmB39yRR5E+1yS9UlymlfdmOZ3jK4XH
jTPf20KzH0wQmmx1WCgdc7cddmHXYqJwmrbSHGYrpsIA0cNv8FRbmAewPbletOEu
jypko23WSrK5pSt0fUCi/ncXlAWQrcMghkFHxdrwrZvI5UohbtWN+tmPML/l1kLg
KRI5s6L63LIbNAkMwnWCYXcKgWOeWFayZCtL/cOxmlZBy3kz+7/0JoU7BA5FFSb6
pUMU6fyJLYcgHVIEQeUck3KmTleXeHxFJJZgVcjAKlowq+CzcuxO6J8XGD3OgDNc
kWGyqokM6IJMUzU7Nsd+70J1Atyq6Yv7nIHWyig6m6Nrogf9rShsCSOyba5+1LHl
A4PmLbsNDWSIqG3kIYV9MIzTEzg4rSDzBfz1hKw8dFAi9tNn6BMTwTXD6vzkqJmY
kVjk+lxV1xFlLR5oRxHKSuMoTFlleMOTCaLD/Uy8k6B9eQT3G/J1bQ5OtqLAmCP/
7FIZ2B4NpPTfO8nVSSHTpp6Yj0bVRFjjalLqmbhRmxgDmvyClX6qCnvWmzfoJatT
9DVG1x/kcA2hBKHrzMWFNqUGQSm4Wl20DvHb52YuKsdNONW8w+otOW7xTNYMkYF3
oLKR+RVaenXErZBAnlgAqlRsdqbM+lq0L9KIZayjL2Y5Yexh+qqEFsoqdAsaAAnc
O15M0dKY7j8vZ/yrQinayVW2me0ikbyiQZK1CnBQTq2QRcS65X/Pu3OUBYC0K6X1
DeGBFkDMiQ3b7xo2a2HWocYvlwv3DWzczR2HIhFEQg2InBB9zbBeDjx/b/UmWgZX
fKZobbocQXqFMIyNHXvEpf+gIK9uVRYOyQxqEwZ54QzN+wlv35fzUYO+Jw3Yl7iw
DzyRG1XDp4cFovZ0/RdAburMTmaBCJ3MqMFNICGrI9bgSMOwClrWnMhpJOxkH72T
T4x+NZchzZVzsyNxpEoJqXe4G9z6f5A4ySi/sQP1BFsUnqY98CwlLg6GBjVlYxyG
0nJLenAiq6zXwM7oYKf0cB2v7jpw0f/O5mltxKM9Oc5KyrL6X1zH8b6WU8TwXmNG
ErOYrrlQYKyzrEcPHVgY91vNuFYWqcLSW3DDbZcBvZ0EQVOVvN3pA6BcXITre0Fu
qUaSTQspTd+155wyYMmDr4MN50KEF6DGvXInZPA4N9xNHJN7jtMDdM/rWR+GlOg0
QQxTSWG9yVb+FWMmo10ADT5xJCd+LErd2SuFrlQTCvBg2RB8SX8ZRAZjRhsAshva
iHnNJ97p9T7qgb6Cj3elMNHC666WSB0X+ltjpPeXJ48tO3mreTbNbbDQI8BpHOcu
e3y5LKA4EaWaeM9FszByotwLfkJ4YOJbx76na2aEzLNLYENexIjTxw6+AUiOZZNX
B3WQX4xuXrBgiqpSuPY9IlRZ8MVytpIaURcRl3n4D94J4Ho/frKkChagXNDhrHM6
1o88Uzz9hCvDY7kckpCrKZ6K+krPcCma4jiQboA3HQFX0uyaIZ0JaAHJnsOG26Fy
8KYpCdybcz8mk5nyQ6j3dblYikKLhOn2PP2az/W/i9xVSjqfATQbmO9LimeOTmUT
DHS1z/FKInnFClx7usbuGjV0RKG2qg3XeqJfgB4u9RMmyVF7/THcqdlRqHMH0wfE
b+OxXVjc0FZLc3n1XdzFxrpSd8wxo7vas7rKNDb6LQAQv5WiVVoDDIJr3/2vmAC2
wBghYngDDNkv8rdc4S5SVJnKYb4uVodyoK9uGx7vyXKr5FgJ8OnF+6F1Xhy6a466
wpzyCcV0iV/t6N9dOlLkunxJ1f+qcm36fgrpM9I1IRS0RTKNeR/MDAzqkakSzmLv
xdf7EuNyIqkmjOJdRT6nfEOpAbJEBjU1sE2+bJGfzXZ1/4nzzce74R9Y5UvBEudd
MXjScF5tiLRA10QKwVt7osUfDnpUpjmv3HYY1O2cViwqiw+N/X/pEPGY6rw7zBZG
m7rXIfw+oRggHB6un99S5vYaVxi66KG2rprUoewGOUwivz+yvQjNC7vqY5fQUIW3
kKg1ScCua54kBxPZhps5BAPQfkHIYViV/HVRjP28puAL6ODyahXXRGwIpkQipn2K
2gfdVJsJ1cec8ZOKgAE5Bkg7o0aMhqppiacnv/AaTFGAE3N3ZSxJDLKVoGLoDUkW
40lv67FwKsZ95qPXTtajH0E2gb9C3EsBWY9QbEiYBsE2nzqlQ57mBlY0r6XhuEx3
GPBngEJsuk+WC8ceub8dLshrf2Y8c+iiMa2703Ym/wXQ8M2iVcRti6q893yr/MvJ
bjITAHSfiDZbN3XGgaMhWMXsgp/zv4aPPMq/oDVV/50Uad8zy+R0FoMDzRGYlarr
1NzzX/IszaYAdU1PDc/aiGXHzVay7HgktvtlSJSpspbtsz0jVr3I9r577w4KUZez
Lfs1L+ZewSjQCat+qnnaezsLyspOzuURMBHDmsue8gY/Lp//eQyz/tBghuWzKLhV
wK+Z7YA7iFOlZwgeMyMENd2c60gEdeuheQ1PwD+xuML/dO208lO1tPTfciuI++Nm
vF6GuQPKJeuxeGUmFb40C+2rT4ARSbxNJYJVRR3Pl+ZO1MnrLTRrUo60RXOi5zfS
ifc0RkUxA0L5W2QGTPef2HY/YV3Ay77DyUtB9HH8/IH90Vo1Kfi78V39kMuGrNIL
krE/zooxIiYtP+Y+ngUeDhWW1+E1+F1PhKE0ouq+NJo1+2JvkgRfTtgfBiaO4nKe
wEwnat6wxNN3sQJ2qHv4r1BmINI3Am9lHJZyv6K9t5b2QDtkFzlkB9jAWi7MefmL
MypzhdClcbD0nP/uNJ3WQ9WT9FbYStwSa4t712mRCIyBhS0y//d/XqAaBOZyHwLu
x7axeWV2XZd95PfpXqFQ2GXQj5nqeYQj8IdzlLZAJCSu0T6N4j78hXK0ARxPajs7
jt0eWqD681wX5E/8wSUKiO8ol3FCorVuh9we4YnOBhrGt+qxoBHTy36FDsotyLJC
akrjF/dy8BZXS7M4Px+uLaqDPIEFaEvl3jnSoYsQiEeuSy7o0ojMKLIyY2FIxpZH
qeNoJm8rqVh9+kwHCaRXSkgeUynWvOxo851F9UDpuHjc1zDKO6IBKA508NTX1Nm+
KrtPpeoqpQQOlmkydzD875RstmbNdCbdGXrDhUko2C/VVvbk50psFNhskbcBNxU0
UqAkg5quYUthJNNGfKslmOJVgjR48BKaA5/D+ar0qdCMmppfqF79pIwP5YjvfKLk
cTVg1RNQ+7gPPImfuo8zgp3TroCQ/wdBelWHxOPaWcizcxM67rwqq51qZzWf5LjB
PCeE7mlEJLiEVQd9/DI79qTPDUu26jUHx6J3EkhWWvQOaDbP9Reh6vunQwwRiNob
bUSX+Ut6K+0xgwgqLrnASTHEijw/ks4IyOTUFsKsYj3ki0ylQKZizrut8NM4i2Ti
aUIyuYpnprYY92Mo/bCWV2DRKcCjK1O9oujfsPamONLpXyTzEAH/+wrcg/n1PK4l
uZKNaw5zs98Hyf+AwuUutaLa3ylivYZFi2UuSVmddjROGl7HPC7N/K44oBGAdcIL
3timOQOOaWWdghdyVOaKRWtv4yoWq4zGRTaoJ+1u2T7PYUZDbVTPIR2PjfiszGb7
o9USjNBBWum/najRDF8QsZWpWUqvG4RiVri1rpcT2+cq2j5ITeHPcQBvzguwBebJ
F/71uS4Hul9Hl1u22J5vVreyPo5oR8venOF6WYhQ6JCiCDJXyletOFFF/kF8A4Qp
9f6A/lMPW/HcXDN0hYetCN5DPlTKn5k+gHlxGeBRDy4TXfIlvB3N0DslmSddhi/r
8cXzmITAgiGGvxzx17c4WMrdCDOZbVnzHb4mQcyHaVBvq0yGni/+Q41rR6fyRSal
HUHuIWnKr4/0pLfWHlRpjo5nNO5IaJhavm/uLaAvozxOmtcLYaW9t+Dm2cvlsisx
o/eCPx7eGjgckY0v56VxVrt0p0lGflNbPazl0wOy5+x1rnfwNuD3ygpGB0cWGcH+
tDdU6FeLZe4ZJ7WEZffnYM2CoKyOtBGzXQodHGCrk55egksHyYW7PConCL8wuRFC
9OG3R+9qPFMta9JsVBfCN+NGY1ACIjfebCrvmhZUhomePsF7e58dzPXebJ/Zqi9T
CJfm6pUHTVZk6QW+LU4Lk48AV+vR2A4Snl5cCtXS4b9+KZOjtoi4fmULPwsa+s6m
rm0CpQmqxfiz9P8Lx+Qo+8KiN7PZTROq+1V+9Ufi72xHHnNoQiFSy1RAhywioUML
1M9u1FaagPjSqdahak1yjY8QgzEIn+HpvXkDYiVPzMod6bHiLRny9ap5H9/E3qBk
r8ELr0Yncp4QiImnw8rxOTRZE9XTBYw8DSEZ7TNMG1p6wSbsQ4OJscrPsTVXm7Qf
RrDj17gI/hHzcPCTNp0SLZGD6oDuNerPIsl4SXSOwe57ifEos0QxGdwyIb066NHj
6JcDN5G66x5CCvozelMyAuLNze7ciJrzOFbHSuozlTgP76wW9SGujBpbCcXbxHY9
Crq1Mq1hzjaJRWUMQmh7hkRQMPs2UD8tE3NLBXZ01M9wwrgO0xggIwRxzbo6hMRn
b3Mf7ouHJ511H74v9BR/S/DGuwD7S+Ar9v5A32rrSZOMcdtj7MRmMQnLHG1P2BDy
VxLdygi9WwjriE+AMe5f+1M/eiZPh05AcixV6bQ803IZEeVWbN+TPfK98Gg68/2P
gcouZaFXOPWzXJJSfnSkRaLQZpVFUplQWgIHsel4hrnF2gdorZD+5r/X58iHGLWf
WjPYTm0jI50ivNTKZmhe5Oqs8J5eqkm02zPSPJS6i44LR2+03CRyZAzI1sJ+1lX3
/qL2ENx99q4t/o8VNsDo+v6U4En68xI89Ab+mxznTDw0dDB7rAIG+EkCtI4aGcYk
VPXppM+WYAAX3fj/W+9ZuqUq+esBbX5/6GZBp1BEIIlwBfsoSKroRJhAcmEeoUSg
X4wEJgwKKgv0Y9zkM5uSbWrXxsQJgkGqZd9NOyiO8aEQYvVGnp3UeF/2npK5GzUq
VZxQr9AcU9bjtC9Vj04CDz69Kcw9kiLjvPMaLd1DofEdhQjjsr4OCKOV4JSavFts
61YxwsEemMlbRyiZYaFvvIQ82QrG8lRLBWDlJ7VFojzy5LVwhlaFoqrth1akEcRz
fxGQLG3G0RqCOc3wJUftKwJwnztOVLb+cTv6TNU/kBQx1XcssHfocgdBVrcFiEC7
uOWUy2NEPt51RjI8aj8v7Sm/9hmGl733cNv5YC01OXQbo1woq00Y6iQb2CCP4ONU
cj9E5QZzJNZ5I6NTmQYPiIM1VUP//YtxSkYLzDvKuNcCk/hXB/a5+XVdde1Q9mjD
CNuCXb6HnyQAixqsthBKodWKwkfkSJ0soHdy9X11MYTW2drimxOkKRrUr1+dCLg3
hTjz3gIXgi7RTatlApyNWBbVKl21ESl+qte9f/W5JW+e+6q/HlKAEBBxZbmuD9mu
MzZ0lCw5MS/lWs+leBzZWfzlxAgdpdaLln8hc/eIbVzJMjXim+OtsFHoXXt+OZ5e
vn7Mhf0ZlK5V/KOnRJ2AX5soBXuXG2Dqmj7/kGjBBghjwWFHLIFoEJcZtxNdbF82
qXaF3Fs3F/K2KJhrwgZPORTxbqf4OH83gKRy82IVvW7Y1vitH+qnbGHSua9X+d8m
Xzy22egkcE7YKUJmHOizfT9de94En7KAB8VhziWWJImz8f81YCCLFMqZXXwaJmH/
ofjuJcE0XI7TJ0gYcx6SR0DSRPCc5O//AsA/ED1QR9G2eZqlV62ED3NR3ky2ln/4
6I6NCItxYtXnBdLk2+DUtcD9i49+eTs6JPYdJusXQXPp6Ml5Bo2rOVFpnRl2hqbu
FTWOqwudoLZTIEF9SzvbsEURDTRRj/XCMIX7Cq9lzII/dcI+4XGxqKHgDeRMh4mp
8iYZ1gO4cFvSI/GMXhX2NRGv1mo+8uwpi6Qs5cBB7dbwARqVY7cCrN+CH2yfd15k
R95Qu2kGc0HLr+Twx7zSxHAjZJ1MdQqptUFVQxEhDRiKfbCRWQbZIvz+hZwaraGt
ZN+tdulIb2446eeHtE1KA6zBkwXC5PGj331xDL0ALvZP+NSBlbRKDtUoZBhrVnVW
xItY3vPxuW0UuEv5QTJZN//pMD/PzLLH2n8SLIIuVjOQEfvc0zuvixtDLAjbjNGo
yar+zOdUmXuwyuxzt8OEp4jy3jjf2NJ2KdpEogjNr26gAK8LcQScbPYvIw1uUrmZ
FV2wnlTfq7/RjA/A5LsA4BNGT21k/eXw0DaqDrfj1gQy4fL0xOUgrROy5/Bl3Qg6
TiYr7CMdfp5FE8y52kaVIIVuTUTg8QITYCAgVN+dN0moBRpgBomj4ExCWHJRbvop
s+cLNiLM0GE3i6txLrVB5qQH+0YnGcnM8Z50+DLW+Z39otThkO7RXtbg2S7eFY/Z
U+InJwCZ+hKjvP5hQLvNIymJf1RloK9dt5nN0h4g7uSMiRLFzsqgbuMnlyjsqd/q
ZpfWATXr3KbZ9nh7A1j508YgmsEc7GloN4IDPVT+sodJD/qa2RJRol6r6bPvBHn1
NbEI8imEUB+tabzppl9fMb0cZ+fRUOocq1tQ22RPBbLP3JUkF61fb4hMD19eqK1s
Xkb7PeMTBpP+jNpnbhGYy9GYsHKiJ6LBJzVQKxXAnDR5tPE2s5zoqYyTHJu7YrWl
d51bFAUxsJ/QNwWfgYtuPeq5JEOujzDI14AJYPHnCbrcWA6TPVs7oynk5LUecMlN
sXuV8cpd8rK0JHEfIJik0ujDTVtxVNaGKDkCz/h9gcvNqgUfhNYygYxqwL3IjJ0x
Ft/GOG5cipzSSQTE2HOJTzig6nPcJ7LEpJi3HbVUeJTVq3BpNtE8TvnS25OT8nTm
Q5//PhmReaFvKaz1fa2bTiwYJtJFbqqNmletnPvseZnPGrJtnKm4GvbIQrjbbI7F
MSKNmgOxD7fF14zPS2jiUQtOTeXMq9eANsBwZUbOkOyBmQRUxJrBJjDftLHyfne0
Nmn7dbEm/+KwEUa28poYO3+zTqdHnpgPKHsQJ++ZQCxXhZd2f5D/UoIm866+1vnZ
WhygZIFdSBOt1Hn8tw5W674T1GwTkd9moq7DXKOt2iOgZ+2nnc3+hpK7MbTwo6Xh
kaPyMTl2zWNliviJDNCDLqWUYodmJrNUfG55Euz4yUu5F2pIbuCf+5i9I1Wteu+q
bnGSINlg/K69lVnWzCC9Otj1NTNVOlKJcB6ydpMYWsIBhX6vs47Hc/s6Sz11424h
vOPgLLaRkWQxjMSEFn7DNlLEuHYbTS9CTXLm+qrRPd/e4NR9U3s0u9Cwd4ESgXTt
WIii7YkKacP+5cUNdpqrgpFfIklKM+RPyNjcArWznY7cG8lsWkC2tfo5UkbAsx5A
43anOY5B22WsFG2kVrZfyJUS7OFDYji1JpF9eeT2ZYYujmwYR3KJ69qes88fP4Qh
0EX6dpzyFXeGQXMfvXdMOzlUIzrNdp1q5WA2TZDLE5lsIpj3/ThSR7A3kbyKUgMv
Kq6ORxaHN6OHW/zUiZTcNpU2gcUcomVHB8q/vlOoVsUfD9UwRfo096/ZfSXxs+OL
OcQoFCMDjOD4dRp9tB9ZCsvXzh+aoMPJwqRukNHijqlOfxOuDtoSWNlN0tZIyjnf
NFD6pQ3EcQm5U4ZfFWvKqrzi1SseYTH9VsjLrWX1Srnd7wkaoRHHNnPdtwnuKiaI
PeaFlJ1uZYn5yjB5hxChB2RMYLcLALqSNZHAC+aMkFErrd0TZCl7wUjuvq294B52
TpvFJxHuxurFjsyWAP9KZIfg62sknxvJ2PX0K2EEs8mcStqp5ID2Kc9oXcIpTDLZ
X5DfoGCWJ3IwpRbLBw7XZ0oBaQWqVy4AAxTJzYetbUzHQMKHqOdXl9qQHGaVWuIa
gPRSub4hEjHhebbDEWNnBJ+eB961TxP0HgljcewvHb5V9Rp+ZjtLXpEce0+LLe3y
ixd6gE2ssOie5sinMlTdVnnHpcxlAude2qZeOoeJ43jmrV8BxYCMlDz6qqdeSWel
24SyYWJjK+TG+8oz+P5SAA32xliPKARWeZEjkR6MNDETwWt3bZwdQNkgd03eZzyb
U4SjdNJQ2c36/M0wmM48/aLIGAFmJGx+odmJ7NKDEcJqCvc0Uah05o0DcMNR5sux
uxGwvqUg8EgzJfG3B4Ql9bSKp5Hnnjm7uTb0H6KhgnobIfE4qUZkOr3cM8D+q/jI
eRpkyPqDhcKOu3309hpBLB9MMMK9rinUkcvP+yJQPwDAnV1WuAKphupHqflj7lhT
/WsAS/XCGc3wluocIKmZaNXL09Zq9qBPxW4jxGAxhvvYDiWXn5DIaHi/57OUSLeL
4WIgPCVMUDCC2L8d7eRJjwpNzVqaBR6igkgYIuLdd3frt23g8ZcMJqIabsD/0SdU
pfhXsQ3D02p2JsURG9RvVELIhhYX1wDWyWyeBEMTNMhhv+pqV+94TaFPD7aCx2kH
c9MkfjXQVHiNGv6Y/T4dxoOp+uFkc3kowQaNmJeqnNGFQWw4FD1ByIYQIV0d07ED
imw1e4io/5+SBTDVpKAFprOutGpvub7jmbiB9NuEFCP//QKqIFkX/8uqIsJB3c0L
s4e+qlUNaL2Umi1AGFWEdeiHU+aCpG2efLnIMIkHTdApR8Ct7srYL0PiXoKkO1AO
PZpKNKN1MeCM9EAmeK/I0njx+2gxnJTpoEaniKP6Gd/lLTqRPswJ9yZaolEropOt
I/SVceKOZZy14DAafGWxwVsYuUB5YqxdUj/ULjS4ijtms8upyh7PFwgvYB09uA+g
WRGW22p0RvDwexp875YsIfNk4herx4BraI5onN0ir+F0R4LFPVkMJP73C51alzeV
zG9fa2Sh5Myh4+HrqjUhjk7jxm2I/5lSBqtr5/1n85UGXla+kpXMVjZvy0pA76xq
Y/xD2x0Z/F3fANMBKtA4bklV6lwizncM3RwUzp8l3jl1MUr3uesXCwJ7F5OJI0sp
P0d3rcViUmQEq3ea9MUXhWLjNIoHP8Om0FwIy46FQPZoG+8dl79YZYrbZhD3Wq21
zSbUa8n4HWUZIDs0iD3wLVjfALzid7ZAJIEKe6S9ORuuLEUeAonGiDVAavHUeEnN
+CR+7e1sdhJdXHx1vn24wPZnbLxcoI+0Cj/V0urwDoIZQHrmtjTo4ZGXiKXRPVkg
7ZJ5nGxERwC08lpCVkoTCWdlfzcSk2cfHO/zXk956XlbiaX04sDwc/YIPH7/3gbX
1Irk0Fas4VGN5yCuzpPTnSU3e7RRAct97inM3UNcNCSIYFH+IpSu/RXwX+jglzpe
TRGbQcC4dgrp4gHV2Tgv9gEtlVMU5TEOt4EzuAM8N4N8SI39at/KmOrhF8pbj9Nk
vjEiQI/QKAo6eMzws1Zgk6+glN13C6AoVUTAX20iE8XEEKtb0nuIXADGkl1hOsdn
ddURfd/k2gDhri2FXxCzcK2s2vv+CL05WVtpjz3+K0AiDRHut6I4ALhEjG+uDomL
pHZZsbKJouhLZloodcyT5T3hYOoQbdIXdBYJ+cDcKduqv0LTP9Q/16v3qniAZs/h
/u6FieVYQYLkzDIJtTmfPU3b34btX+QhJU3VJUJwYVmnBVY5r9/dvIgOWrGjrJXZ
17EjyNqmzVXLzG0/hahyYnn87GyprwXYT41tP4mwfB/5BeavQsOp6Mzwt0DPoV98
eNdVyqik26vPecUkmFzVLpo6jVnuV5WXBnkof2uelySe6E2g+zAjkjFwWcbwM+KR
Quv91nnPosk2OurVihuPXgvQiXEDUMKpodQd3r+X8mtyjke671NDKF32c0fWFTNn
53YtMBunQ4v/t2UZXMeswHZf4p02HMjUuxfBcht3BDNjHRghaN33iwCUp/9toBqm
fWzoHE928ErDKM+YeMeBukA3EKoaoIRpU6aRdHHz2eFlKrXjplai4DQ/m5ianBuD
CUAOxNGxoR8FAv+TZhLB/KZMVySE2L3bo1QQDSPNZ8AwAZ8LlF3n/ZtIlJnu/7eF
o6AxV+rXWcIy0VB4ocFwuTUwhUNQoCo0PQdsau6SDMqON43FlziIRt5P68/qgFCD
qD7ZMM7qi9lDyYIjQahjGfHeOkORgsqn4a7yKpt/luMNvWRl4oeDi1M5/LB19QpF
SE9XXj1vgyy9bKevRn0RkGThQVgllgiRpPr+3z9OOuQhv02EzpvONLkEdftO4ciw
ZqVYAmPbc52+8wuu9ApnTQXK9PmrvRLxm69TJZXcJJJvnvbOtiUFdFUJcDkQxSGf
9pVY5ZwUrb929vuODR4dzxnTHKocJoXcsM1gEMZR+RpATXFEYJCTviAP1HfM+xAz
H7EyQ8TdAzRt/OxWD/Fa1vS3lvgf/82RCbvOAFHnRKVh0N/Hw+z6ddRzo6HB+mNA
G9AK9TT+TdimXkMUYs37Ni0F8+ON4SmuePjeCSu2x1oOb+HOm5KbXg/BkBKx3jQo
PQgRX5mWhC8pPyjLkt9O+dDM7VUET1Q/5GzJQg0Nv0wefv32/o5oUBABYG66t+Vc
yWxwqcHGFcldXmEbp9162/Bnc9dRrge1qppKslpYdkvgkdy6cE6vRAx5ZjUowXku
KIPHGPjMFKvG8A1U4/ikYq329A8EtC6RBBAvhuAyp+6I/c2ZsZ9qHXqlQWyBsbrR
pnPib2zxWA/K7ORRUcR83MSB4t5OFIRfisJrP+6q3mNybdTrPvWHvMGpmdSefhfZ
dvBJaOUyCxXSJBD0wpAp+A3rxXR/ZoxNRyDM+5VfhoSuaykUucsgci2C4uwy9tvw
lriMcIsfgmnLCrLq9hO7JYnEMP5Mfd6c3XTqtP5r5EKIWWADy7pXo1nsbSDKI/or
sxZr3huFOssNYExYt+gtQDUFi+p6UxPLpaif7J7+JFxGlSmphx02FkQBhp80m4Yb
1HELTaVd6IUNZUKLs0RGlcZDljUVpCEF+WuPqoHiHRwelPiovmLIrzDUEWpQfNo1
2DnHQCnbilAM9fNXMyHOZwwlS1PrsMpObEodtQ+A5Jfa8bBadxcIrxuwz1zQVK9+
He1lYfMi64pGuOVq1mPEpgnPiyPLnanEm53Ot92gPTO2pxsRlj8Q1YPoNG0Wv8Eg
AY/JODuibYoOO9iepSdJi1mgZIV4M1rkOS2hCe9Vona71bWgddaVqitRxMtrrp/v
ni4Bfen9bIF/9PqQ6x/OsNLl2k0pHlUkvFhLVbFRqWpV8EMwiBkbrrKUzCyNyyBq
1U8nMAywmNGDbLazgyF4cE5HBRk2VA+lwyfdiJGB8J5NbAAJQ8+T14gm0NHNerxX
nK5FIzmOwgGUXN7Vjv7aGlBJl6lhZDA6l2/hZOOmGmZmw5CptY0clJ3s09offE+O
y4y1kQAmsrg0nKSrfcbzDI0xhevfMwUP+YzSKOrc/gShJAxyZTslJW3SN3MvUHRm
WcUyrfSZJM9DBvawuY3vQNktWcE6i2Y6IJUPXLLPx/TsJCYPh3/OKY3z92JW+04B
r/ePj9deqtM0mpIzMgQEdxi8KYecpNOc1ov3mFPmXb5Lw0sAeVRM7WfkNXGFYsFe
r7qKRKwXwKvtYynY5gGXswruP7Vtpj0+zjSkG2JYI0OLMkEGxu4Hwk3D7sQ4vcfc
6Ah9EqoIT7CGg9NT043ShPJ02/c414wec9443oYjNSLrWdzg2CR51hViA3CwS01D
MY0+bmMGHqI0DERuRNutJKUYuSBgNo7Sl48V1CtN6DbvajEfGowlEP2lVmXQ9Az2
ZoCLiQSJvZs8yXX6Po7hmHGUiaw9uGaH3T4xNh09QJZ0B6HixMqSczbMppyjhrtT
XAiZoNcHc4pFbOJLJLaXVTbmupjtyrr/k4ybzTQBpZP3NUvtl75Fr/xLAjQoLuUQ
h9xd8lQSzocWo9ifzZZmH1ZczP3Fq1Fjuw4eGXlpOGclG+Cj9wz1rWUWgFdB/2LL
39dauSuKFYoFCk4DLRy/iF7Hvmk7hash7OP+Duby9I9M84LJ/Z+KPGfg5Nfe5Z5o
VJoczzUzVGnJho8FDvAF1dEsRdLCBs2fjH2jEnSqwqIrzx89iX0+5ZdDgYSv1eo+
9Y8Kvrk59pzgsu5rX4jj7s2DtbK0uJ9Iv2r4jVNd8sg0UsS1dzrAn9XErwthyV4a
HNpHiBaMarSUR/aIj0ircgvDNbKfuAUz2iLmmibyo4FwNf/o7NIK6arNqJfvlJvB
qWeQ4wzsg3AuqUy1PDYVrTtEJ1pVvUpXk6p64NGZqyBkXHa9EgSsWnevG7eB81e9
Ebl0CXedUAr0G6T3Z12fzHdUDTawW6M0GNuRQ1zaTxpqcUR6Ip1PMLKI54Y0H4n6
kWrofy1OO/6nBHh1d80IywUdhc0VeyYztHc6+6wdDM94p+Vt8zNcgCTX3fLmngsf
sLvqFF2RMGePSHwcRIwYpxUEw13+OPMkRVL4ExV1fqrLyg7hdesCcC/reNEoMFfc
ACHu0IXC0XE/qs5pim7EpSjRekcEArChyK3+DDG9yyMU3Z3cMGXH3RacxOJrUNBR
grNox6pBI2zfE1iK7tZIHdZFtCdrXKGsYazkK5Umunq04D8qjtJNBbsPtnGdF4D0
Xv7cylMjUw3V41FAqSknUtAPFkLQc3vLX6VXUQQsMJFhIW835IvQaL4tCda0vV+J
qjgKI6/Y9dtxLsecamAwMBTh+7HJkIL5RfoJXvAKOSfT+raVH0dq2mdy0z5AFq+K
uUvCfThjzd5iVV2f2v9MkEwz1cjksdHWQCWIVg2b5npaWDzlFlGY1L9vWkM0ZLwZ
JR0UsbwGnn9lBn2HXN3xfFUpsabSjffT7HXs8aXoV9yUZJlkVCyOP4sbbg8szYyP
3yBz2mqo6N+5qMCC64YfyFP8hSGj6XE5fM56b2XaAH3ksgXh0dGrRphq2By547nY
+cSHBIjLRG1MVYi4RCkEpq8/HlRv+0T09qcB3XyCaONpUN0fSgWFS2f7qXl6+FAU
NfJdZ0I06DutUnfbzidHsX2Cmrl+FkypfHsL3bGhBF5cdQrJ2TjDfqqtFXXEP9+l
Gwsq8xbaZYeuqm/KwdmU6TWPH+Hg70oky3GbVfNvUlIRDyP8HkiKEe1Uc5qK62nz
yynsQNiv3evzB6tlpLkJHEsoRbQurRrJZdArd/SSc4FMpWx2oyrbyU7usIeeqmYo
d1TPXOuwpDDmRN2XgL/U6r9fvqMN3STAwTDh/t0+nlNZ6pVstaEbWcvnbTcIPkRO
AUDcrmWIYMGtq0bVr2oUqt5PAQUoIz19847EbvWVccusVHxF22/b99ax1P5pyncY
LwfqG3tzZohkDwVuHg93REZpfiZIKtORH1XkH0rNi193UtPHOBOx+9BNj7tvOXWM
zb4lUO/zxuMiGYY9oAWe8VJyI06kqOM2iHJWYEUvKsVIJs5X7USKlc38JWjYwC+C
QgMVrovkoxQvg9NtdYnb07y+GsGUkG1et8CwdfpnH3qAOG5kS3qOSzxIlSP4iJy5
S0AMeJ4BfZ0R9K0Xap+gtdsF9NIR/Dn5AdcHf2fvvjwt1Ovu8IpQFheiBdfSTYwO
1dRdE0KWISLRXPvIL7uoBgL4mvFLKxEk8LmY+VG+uql15E9A5iB2zE6/UFP3qcPI
q7QDVCGOExgQgKTCp9kQCeyfCb+qJkZJWN4aRlz9qrH8vkHyPFL8SAZhWMTGbDHg
gsKWs3Sl3VOoA5TmNOtK1/t+P+IvaqTIGbI3ET2wtHfTZlhPgE+yHt/aCJJBADmf
vL7qIdnCQkGS+6n36CRMpVvoywINbJemwBfduVBXEuMt+c3Ul9tLwg04DWy6t9yQ
YTYx4ZwRianw13Jayzq8pt2LtD9kIcISU/xxOJPF5qSwN0Z3boowuykEH9deaAlu
zIsRyk6k4GixRP4RULbXPy/LJGrqwInoqwvRi5NFiGQca2BS3D+1FfxKNtMsg9yU
WtbXuqTqJXqjJ8zIxs4YDVnqOxEgqiC3jlMG4Eiv3AXLBBC0d0eI+6txf18syPHk
2daRbt+TmPytYxOFpXvRbYblJ7m03drftgztNNFI3rymxo3ZbBNu+DIXhQLQg6Qv
iVWAnn2LcnHBnHm7PYDtXrD//Oza1h9VEJ/+KAChYyF4uey4t8H66h3EYFOomueD
qn+uTg7SyVBdxxaSUGqH7JCr5VlweOV/32S0K2QKf1C/vaFA1JWSNil4qNfJPXVF
TEQLJD+j5dOIGntcEtYNY3s/Zsh+TSOp/wDo+wBJNQKQylq3ehh2gr7Pe3q8XZjY
6L3oJSPPZB3TxxoEjCk9Tg8KIHvRco9COKIcwqYHc7D9WO0Zdw8Vt674s2J+d9UM
R2b7aHZq4/+XjvSCrREF/MomYn+fWiHhbfudIkGaJPQf5KPWp7+Y+/gZ1eCXrfE7
CuS09f8sRodf2Il9QI6pJsuwFyj3mTHASNQEPSoastqZNBfOQx4PSGTm+yjt314K
3cyL09/yCIyIJyOU3NN9lG7GmknESVvYajH6bZfWVNGyCrQ9Cug1/KOK41XZHTHC
z5fKcm2YMpKbH2/k/qtQP9Hs+Kx8/A4CnYWa+l5UBi34T8X4wUj1c6bBS25DlToy
sCcjwn5cRL2mkjBlTb47SGe8xR7Z2SiBOgL7BXkUPTG8rnD4+uMOSvo/5wFpS6PB
WSH2KzG6KcfF92UXxomMrPEbqbeUW+tscdgvlAoHV5Q67R2SdyakEwL0w3ycCeRQ
aDJygZb+GsmQpuzZKS2Lu56QvA8APRLFfh8WGdJ4/92hhn0vCgVpKtjBzkGMuL+8
fpwuhOMXp+xa23dNi5xVZwEOzzOVL2ULuNFe3pcQx3CjgwnQIchrsZ0J+baptTYp
kUlJJwncxU/sVNfKqmY+bZIsoFDLURjsgTR2RTfhUy5QXLQMLry+GCWkQazeuE2p
5J/6Bbk7oksy8nP1GXvmiKaCN6qwFy8y0pJGAikDKZ1Weh0E0PcscQpE3D+cMk88
GdVzco4a1ZDhGdAFC6HqxwXK/wb1pVTBMpjAbdD0x9nCHxbqaom21lELOlSl88A6
b3pRojgJcRN9EEZmk25fXsq4JdUyQPOix04hFR64u7BVTnxATkMqqUwpBDS3a7dM
9+tt//IZHBUvfmlNcc/YjIFTXcSDFWDuXTMZuX8cSyhgmczCrl2AvkyQLpmOXJI5
KoPsYxmBsU2g3qFDIyYiIeI1AhXVjLfhY3q2SOo2kGMLqxI0E1IyShcyziGZFMdM
GfT6iAv+BCEW7YfeQlO0w4CTrvAV3iUG78EpS37C98mLnd7wTSP5cs3NyauXqMzQ
qls+dM+4//Y/gP17xirQjFO7NGlpNVp6dbT/bKMPG+oXhu4/75Z16vVswiR/ANXJ
tCvE7XmSfsFcyCynUPBLzOsbrolUZkzsqrbW1tZGguMcQT17WwELs7lV32wE/mrG
uaWtOwiZqGBfwYlVvlX8vy3RJoCq2xIsSiyky3iP020IRoH62kTGpVxexyj3iZY2
wClE/X3YKg5eSuj7VxE/fCp7frU4iZ+LeHEPGUTh3BEC4W/1nQL5o3TC/Q+fvx88
1oEmsMmxweBn9AUQUviq3L+ENZH1y9lte3ar3Ne+FpIh8MOqy8w85Cq3TEfct4sD
2lW02pZV4TWMyE1mWocJ9aHQR2aQZeifofe7AYxVQThhgUYIhI4j6J3XH3p24ryw
c3TOSdAslo75BKn/FxdkQpk5SEDsCqKULK5LhuVhALn25+g60krGlozp37UxtamR
BvLrneASpmj8eY5GvxFEAv45Jt/zPIe4HGMCvW8o8QTfBo3g0rLHhAp3EzpZf6xh
Ml+ivX4VElZ+3WVmfsjmHu7E5MoCvdDm1O+L9pEMJl4JxRNZBE/irce2prugzTLG
ALn9ZLqinM5cTok241kMcRERTqPns551Rw4uHyTbxIQjldFfIvi9UZbFid8OQ71f
Xg/77W/qozr9rn1D3iZAyLDniKlhhQ1eXm0t4dpnLHCNIntn6kIvhz60ZGo6XBiz
VlmAcl08GzKR8TaB+F6N/unzvU+Bhqp46qVnq+jHcLdY2TMJQL1hE7QhBsAqeJF6
u61QvJQxFByowUd9+HXBb7g3vzmX/g2evH3ZUrXgULHDgDWL/o6AWB2ia7GG71jz
PmNiOZtND1K7CudbIG4vBPnwy/8n6NcB+3F4OOH42dLGKWb3xCzEQCHe8Dr9LDib
yas2RMeiwea5NuSVZ0vzqnozFovPbZKdXDoGmpwcwLz5i8fh8fH451mImlt+FywM
xcvB6lAo5rhtHXWfsi2Bpu1BY5z9F1azb1kl64UxDB1upqsfQ/ia2166R9pcmeG8
+GoJ7TPJEQb/U19uGblrKP/yMNP+4d7762MQsN0iEyqASd5PzvqocwxHZjWmYZaD
VpaRcSGbsb9Z8gSOP6bGZysP2j/9mnbA91Ix/zEo1Ft/oH+XYXxXYvKfmjl7JV0t
b/lkenmsAVh50hVSjTWb5iKEx50pnyTbPtaiOdArQjEygUVd+pOPydCQZTdG7/vw
s7BjVjpcOK+ddCmBp9NEqwlb0AM2c5GaKd4rY7rpvQAmeLL5e2BLN9d+ilC11ycB
kkJEv5OETyvRCb+XQlyKZ+B6xFgKD0ai3+gHvJ+0l59AiXFdRZ4T41xc7Oo7Gurg
aSS/CktSyDLVwXnCDvVxuFEBzkCkhVEZan9sXwEBbGgzfmXG3yEkgyBaqAtlt367
H1WMoWdIi1Z/Tmg3dipjfB2hiGqa8c8eAgnrcLCHQNiS24DUHSXoHd0fRunu3uHJ
RjZURBpIKmRl4VS4oxoDcb8/CetBp8bwc8zvnYstS+9UUqSww41OaQuqPQ3OwaQ/
dVvqPXPRMtFRyc+s0bpnx940Y0x4sZy7Oh8Y7aefCZn19WPoCmOjvCkzbm8HLBiF
IHDBqpErIA1wqP4sE/VTdiLWln57J8PW1pvMRYJFcqf7Z2Y9enP23MaE+estf1io
jtfzKox7wQ3vXeuRnl4Bq/TKWCVPD3wdj8SFFRirurUDTiNGZdN8tYSS/JYXLWKg
dPkKyuaPtPQfIYzagb+avJgmvYvUhEvXF8Md9cYYl2kKHmzTzwovawJYeMJ0P3aX
8HV7BPPim/d28iQq1YeMGhm3HWXo4QW4Nb+Gk9+GcTw2u7ukcFe7SIxtJHyo7u+H
afa8tOuzwEQE6ZTINEi42FZZLHycQdROrtXhBvq8ezEq+yk+8Pym33AKrHqrFQuR
`pragma protect end_protected
