// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
IpXlHpUMEdy5rdeGkYTlug29icVb9MYiQlmPFwqp+aXrBcxxjmGMKgQpzcy7c3IGmbAAIf9IQxjK
GTQWjUKi9y2V51BWCGSPKvNKaejZ1y15GTsHyxDHtUyo5Vxvr5GlsEGtA0gisUeiXjvybpUOpTpx
JzhhmwGzg6G/UsBoeKekoPArBvdF6vmjIaBIWGeRa1DEANdjTXBmbIdT1AZRV3Q39+mwwsJh5x2b
/hbRqxw1cx0kiCV/eg90XmZaMnS++pMj/Zw9L3SV02XT/9visQJ7S+Sx6bh7nSVfvUF+stNF6dSN
smxcCwyOmbprJHNzSmrCnFE+mOWK6nxexzw9qg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
VfxwuLBl9fio/pWG2ooPXnzp81HB9V7mICL6bLpG0Ck/v4lks8A4i927Et4EbnWRRzE9TjDdLFny
R1D4OzvJvKqdRwyYChYSsC+7N/nlx1Ng54/lYWUGgKd1twJVz6pyCjtuvXHigVaF65ajQ+8HhRwd
RnogTzs5ZHWNY4SEeBVEFY0/iBFWKQsQZaMhDVDSMueS7b77g0hhgY7vP1miMArzHX7x0LMaHctD
uaIbDzZHchhLrq89/OjU9T/3ueLYDCrvOX7xDJUM+F8TVEw/V2riXAURB2PcGfVsJ6TbPFp7Pdyv
C6nbEY8LlryQ9Rov3vJaFbVHf+9erdAkJkDAdjyBlIk+ruL3nq7udKYrXtOko5DnlZOx4jPolQ0j
JXof1zmphcDhzq7mYQemIx3cxUkbYPhx0bXj2rZqde58uehQ9nsffPAoq4Bu26louM1truQKJiH9
wgFOyYvhOL48m3I1Hw53aDXCo0S0Rr0zRpPi4OfGuLtrXKVSddG5smuaadHUHZFLDbGt8Ue/ZWOD
C6eQbpdxXlTNrZYsnw/wvhTHnTWkyf8JwjObHW5LiA3ZSqrUO9xCABUCOC/mUGiKHBJbd1nAaPFn
zfcrtQnbr+z9Og7DpkIRG2QIGARE4npN/cmHLCCIDGRrIybww3cZBbtUfRP7io9fWTYS09wfHFNh
ac7LbWw8hVkOxuK/j478FP/sSCRKZqb3elsuTh/RYX6rf8ofAar7dkHYno4oNFnJoVKI23Fwv6Od
bjNGOD4uqLimPLVOfbmw96UE1uoZk+3sRfMdgrwBQpkhUhyjl7LJX+G/7EzcM6mYw4XZ/iyJMo2w
04UQk2WWWnep4QrEq4Ws4xMhmstjLxZegxZG3gScHyDksgoSBwKhJXdLIYatMFMv5+ZdeHUDHdLC
EHGsC1qTIChcAN4OMNjawnwHcIapc7UR/lvwbQL2K/K5l7bqG/na+sEa+eH6xkr1BpzmPWQuG2uW
zsLdvcjNPdaXP3j81FG/jkmzZYesdfs9iMu3Go7wP7O4l/d/VGHR2fy/H8B/v7DyqkKY0JZhIQpT
c9yYg8d1kCodooAkRoC2PI4SHsWvR6CwFz1dvOYl+z6T2BXAOVwEbNVN3qd/mfUeCHa2Xvmybjpv
/13hhcqUlQvKYfs+M9EwO/mmaPqBw3TorNEPH4Lo+3S80XerWRsSd8W+rfATMUoKUfHZWuA4ERqG
FMVcd2SlxUWzUs80cA6S6wFTx3XgK+iSMH2Z+qbfAn9uA7Jh6iji2hDU9QQtOFy/4h8DBBIRFQEE
w4OkNzsJpIXG11Y9ztSAFDR9iUdmVum7wdP/ho0//WI76NuZRY01A9AtpMy6ckid9ZW3p7sj2WNo
bc3nvIAquy69aaaihJmskupK0cAijrnx3l8V/HC65D3EaMNTnGlJUIt9o/MODjCCR/PL3flmsnRk
wB77mOejXHozk8nVPTzK6ocrD237O0D1w5HGF3O4vBNUo27dGajl2T0e2+bbH+joyOoHddU+o/1I
1/fJT22VlILb0978FUUhDz6i7qZChyjhS708TeqXj6JSdDVDJGqe742QklLFkl0LR5sxvNapBMpj
KdkOjFwTCsWA4GJ50Mpa3gNd8u8m68SnGui05uhlOYd1koN+d8LvZcP5PFP1CbPe0UpHoPkAHyrt
bNL9FHcdGhGCbet0zwwIqwdZ5JxY1Ev2ZZ8uwAUO5xupJ4E5208og+MH4ZSTu8o+xd6mA7q8jviY
ZMJ8l17JoHlWsgKoH7fngWd/kIYM/NQtPuhjUajx30S0RMAHrQVqHngvjgqf29cO84DN6xftelsp
tP8HfSreaii8J4ObLBRr6DJGbldbz5jOMbR/02AOp702B4chQ2NdKLRDJEJej1gXIWXrMYXgTX0o
zQ8GsVQdsbb6XmfMWgxVH3uhVdFsnl9Oj+QArPGeC7hwMBorQDrEEHlEbCYrCyHBGiv0RzZnj44G
SWJqnO6RpJFCBKBkgYRRWay1pYuKdRH29YX21xjBcmXZU1WAEzBMgr2WKKjpUL+ABvTVfBVbtTX8
D134yv0uNs5F3fGEYtn3Ngj5/l1W3F1sQUL1diaHfHokThGl4C05pakLAfznKf9vORzCMmDtrV+o
oNmvj8elIkQwGuyDNSXot5wlDh2xisrJUKuut+xOaDmS/6geP8hiL0ZXR9wK5GqhYUVnj3vjUrW/
44kuQq4FWZUp7w8nArJZ2d3eOhDzyh0jjkIvhk4ELiqJOfxrXvnzA0pn/ln+YpXmYtCTf491N3xF
AADWbkADPmN2eUPxws3UK+Qf/dnvlMrIfLexq+TvKdvWAv0Xi4WVnbmgk4vYYcvPzU5L8iOvuSG+
d2HwN2cWyQ3EKexZ1K+RFiK3h+eSsAUC/VeA0bez01tH4KFqfizdbpSn7Ga2TbGcy9ZUkwNUojon
80fcZjNhkw18AEC7DLZY1RNriKLi6F2Xh6ui1U197nDI7h/K1t1CbJbsb/YWZC3JP0IyLUSoXZw3
Eq2bbfmfO9qDllCBclQv0FKFPB4dJbb7sJsT0eO4Q91GmPr5/C5+qu1q1HND42jqUmRmRDBkeZKQ
kJMNMSdb9Rp6c75+zg5gSKKBix2bAf3YSle+F1t8k3QpBmS9P/HemqtbrYIWeMYu9Pt+QW/b2R/O
djRmeSkzUYQYegYNwin1mPdGGcvLe5JsDigT7o3LxZeNxSCbnrzPiwpF+ZhQoAqSguFDBUrWvPHJ
YhNs87tf29dKrMmOZFRCksuvQg9bn/CD3ASmP80jG1sQ6LjTdXJCeFuw9zLDYJ/eM7qK7Cnym+nE
ZhY51jjWbkgrQcMFjFGR3WgmNSVRP/KLqLaqC2zLcul/ynKc4sBfYbNHpkgx/G2ZYh+ibPlmh+kg
NZ/mVYqtFbXNEjdT96thuHeJAgA+k+RM0E5cb/YP5c9FF1KVJa5cGfGqV51JVUEweGf+L/HHB1GA
ATl2ONnZwDdZxOBJFTG6WsWfaJcXSBeRy8mugb8yChTY0mhbimSICSm5xktI29bEKY4QQf2HQin0
DDCU19DHrs35zupWY4Y/16mvTT8fnQLEYeSoydr1TvLyLd1NYK5D9suudGju2rS1oEyp+B1bwnIX
Na7L6wDRXkaukkqZDJLf+MqmxkR/7C4yfyiYRI/mx+L6bP4/IeWgUS0rK/wkM7HwWa3ScMu+q8pI
07q8xs2hQmVj14xURGkbBUOGYPJCmYBSqnxwAlhqul94jTArqBCH7Ne19d9+Iqg2X+1uHVOdOVfu
h+dH0mDUbj+hdV21bmsZycPfaqwKP9UlvngI4bs7xFK+slMtJcDz8051JK6aIvDmwgcBWX1quEH7
EoMWml1t9OIPJBVU9CAbX7eNjkr5ZBtDkh6r4Ovlch9ye8sBsWqTjTYF3w+qIhBtfuIVvffYiz/Z
GD0j09MdZTAc07et+Zy249tfowfWyJBOtXpuphPzQqc5ghFCf5QLDk5lH1QKqytdP4JTNgvwxIg0
Qs23/yz8aIGyuuX7i99kAQnm8LPLpDtgflViMjsvZZv8kHFFhspj7+hqsMkmyw9UCpM4SqiEU4JC
k0iybG20WaFpFd3h1DOiIaQvY1i0jXLYr0KwMU07mA0aJnf+k4v0tX1TPZKwcsYexx7wIEUZrpYE
weZ8VLDuj1aZ7EUw/LnlXALwPjqS4OfBye3+NzczWjl6VtQyJ+XDYBlransKhm/f9EmjKkH5xp1Z
K2cfPnl+3Sez99JDC61VfFIAmCnH9gueLUuC8oieQPl7VPmUml50Tfi5EjRXDwAvw+xpMw4ga+8J
OTzXQz+EFms3+kQSICGWwGMeq5LRrE/T00VJzXzPBiBkIr2Euxs0QxtxDyhgGT5Eg6KzIWtojzbR
F47ZZQ+s0CMr8sYyojAX3WNwItTrFdIsYm0ZEm4DV7GASrs3RU897Pgb+A2dfFOJbxuBA/Tbn/rr
uwj55HWtN/Z2tepUgYRzT5QBIC340k8LKyway14S6APeXxkCKojqRHhMbLCDUswkIiFFZTepnDie
+DafXcweazmO38z5YoNgs3zdTHsZAECOim0JcmS4R3KZy8gUqqaoP/Psf07AdDZRFsDM9BBkkP5f
cIzyeE7wG5A5CChJaWUVVOLOJz7wqM+WHtuoNFPii3AAhxGgAgOTNHU4LTFg/izgYrfcFy/gb6vt
+GqzIHfecbT1d8fbXr2SFuQQocD9X85+tO65/KFZqyRAkdGCqETb7EwIuBWMOY7GMksQ5OMxprfO
EmYXU1GjqupBwHzq2orALgh6RgIoNq8QhUY39Eet5N79xQLkQviU+l/wIhLCQX2lQ0SCPi4NuQOJ
y6owZUx3nBRUb/bakMaTRkgs2kYZaJ0sg0pSOfoP5HMGH3pcCVukIeUxsyVA8PnkIDMEVKhwkAYk
dhBvZooZc/ZpYzdb/qKeeqQfjAQxz4iRrwwzbreFNgBDNUKGK/E9EaaDsnr55msuTfCJh/xWFw4U
5KWBXv4gtv0N36bRgMy0U9VjjkWo4+B4eFEjlenVubJoytWxrOU2d0Ie2CHZ19z1t6bcd544o3Mu
itorGJ3yH8AMPUcBJX+aKg/L3X7Xmn874amPKf24bZmOm0qQlfN7jyKayIQlGFM9SUp4luT7vrTb
6oS/Dg6Yi90cLdKMTYOtTzcy9j16NdgQsP0Dzyp6RveM50EUFONM2wOD+1zpGZozWEu4F0Wwbd/m
68S8IlQ+xx6AL3y3gtCAO3pSKsx/3lkA0pD3SoWqL8CS1lJdy/M17CISDpO5omYBtVJcDPuti0s1
qVYakfs19FM3UEKMEvE32KrYU+8DBW3HojDe4cj4st+zToHKw4evTZHxwTbeVEU5zFdm8coL0N+d
4nre2IC40JoK97ZTMGjbU4/v8dZGtH1CTiH84zQ99vQr3AAdhsOnRi7V4zy1SftHcnPjo1zR/r/X
WPwMubt3BCwm2fYkan2Dh3fQDb+gofBkeJL5g52SNl7wp0aQxM7/21RQY5U4a+VKxyRCHuVJYnXA
/Ed4TxvfrgIWK8H5QwY3Hcq1QHxP2y5lK7C4oq0d+PYt+Pwuwdc+IRYI1kSqjZoG5e4zQCp7kqKB
5gGeIy7v/rAyAT5jT7K8mKBl5Ddqwd9NkqXyJw+SuKXQCoZ1E2JWWn1W/ZTX1OSi2pVbEzv4ee1m
Dv1Bjgwp3iQM79hfAvebaGglBcP1ZersPV8IpU0CKq9CCzQd5y0Cva5uhjnXlmb1HjfYZtBx5S/C
bG2p20d3XDXklCdY/MC/1uBLEoNvbBgyq5T6v076SHlsz04aaWaUdTWqKMxeg6VTvRgvGeAkQUD4
qEDR8hK6KSD/U49C53h61xGZNi0iIZQ8OfZHNBJTSUrNNJTsyVf9N3NBkcLiN+Mfr2IQFN6i0OX8
jtntCJE8OQeInvirupbejM9hEAGWIfqvRoKsEZpDQzA/71rMDE68WiXBwy0+ihgxV6yJmI1Rm8ka
J3zjCfTfcbbI73eLHb/TOgTGNgDNLcRn9mKUO1tcWfkUb+CUfm9KatABTqPt/f14lpxpNkXXAeTl
H0aBXzb/S8giGog9WpmXpArhq/tNtM+F7StqG6IwAWY8NH/Ip02R3i4nwCx7SQGt1jmcbfl4CQXT
aVvJMhL1dz0g0cOX7JybhfsCkMxvy7rscGdWfONQWpPPlE1siBeSRPuKEaiwDrg1TvbU7msY2+CO
NGibSCMMwrUXanDciJznqfKroNskAr6/LpdlXOZgM53IxG5hRtTRK7+TJHTG6xTLmM5zGghZ5VgL
TYw0DWYm4GW45P5qYyxq7LHnHY4VLL7mlUOKy6C6t5cP1KhgoDa7E37aw0QcAvtt0cvNkLTT73W9
4r3vYZZ5Y1Wm3n/C3ktT5OwJmr0m4LxfP1uGgABa44g6UVspt9V8Y1urHxCbZUaUwNi+kJkwqpqR
ru7DzIvvNQyTSVJp6KGro1oV6LuFBgVedgb8g0C5wcdaNj3StIZQu/ktji1yg/dc2CvcjU5QKyjJ
Y7Nsd5Dv0Y0LTzNl2zffKgwBBxQLFsG6GVQp4etiZN4FrmbrbrconIJHtR9aODqf9VUJjlz9dm+Q
PfpLR3g7taz7bil/P6AuCdG8J+kpM+UsOVoPAkpEQRTOmTMFHluL9SEoQLcSbMlzr5gFVVp8lI/4
g7XRKz7W0+uTd/jc1fXjUvaZUnNWgmmop6dUqgALfOm5aOc8aZBEEkc3nek4in24+k4K17KJclK3
2QvpjsAYugzHyGPh6mvYKd0Cn2t6PdQz4aBX+ia1c3hdUoa+u7bJgMqUzlOGnOKCnIRcG/rzBOAP
gPAbxZSV7Sbs7w1xF0nmKMNlxlcHYxN6vSnWBOuXDukR+Vo9w5QlYeBVo0xFkUild8eoU/kWZHlC
iYyghqkKLqnzI2rPiENvZlO/iYRrDjOhEpcmPQH+yIUS4lNjzFPFcIYtX2Hbr78riCNfPJK38ovm
q6HloLp3PphKLwLNd5sZd+2Ak7LDUDWcv7gMlL5BMBD6lWdChR9s3UJp+EOz87nUNFGf34zrHh1P
yvGZ+FQ/jTkQcFKYdy8OA/l0dmDbD6KwCHpLRbmEjdShAsv1LQZee/Lnn3mtTQ+ZQ2ck6AaNAWld
CyOMqQHjcTAZd24fY3cmOm6TC2ksVYZNtFTEVuDRQ/l+ciT3Yff8CLGVj7r2R/iEzLMV79GRQZ3h
LQl+jxYT6vZvWc3Dtn3OON+bp/WSdpF0hKgdPrsZHPvwN3XbKwpNtVPawTMf7AkV1NSp5E1nWP1D
lEfP7Mo6avovstscwYpK61PQKHOcg6tXyjHP6Zzp8U5NHCnay0Nm6yTvnGM0ugaQKt+CkweNbZmo
SXPqR0/rlzimYL6dsuaI5zHvd86rnTiGPMcucytTCWSW+fx9ntgoHPSQMGtBxhw5Mc7SVQqG+dUG
Ctbtv/krA+jbkSvKz76qO0jnqJkWdIkGfGMFG//r0rSbIvNObG1BO77tQMs8m06N2JTneiUvhf2w
JD18t1mek6rR0AkeOCShXQoB3aADnG5nsQmvxfnO3m5fudMlRJPBU65y/XWKN0MZO1xE9mqSjc3s
UyYisXUbRTKqDD+V+iSBXfeS6iDJq45qDij1IVlDG4U++l7dl355UGmMptfrMuiVLBFm3seG2ONn
fxatutSrT8sF/lJ0Ce2rt3RqjQSdW59K55uOw1j2tRrGwnqdbT9TC1At3nHpv0WbGsYZ9aVjD44E
lbCAgvWT5+Qy/QGIMQ7QzqnvMzEP0WtEy3h6i8eGT1adQCNB9/J3wy6vQ/XzMRmbmpy56Sal2Zja
vawIUJGfhZ4FXVMoKNKPY6Zqq8QxU8L8mMO0/H0Huf2Sy4b1fDYAA28yAZIsYCTcuuiLIj/kKnwl
B68mT5qNCX/L0s2ToOtUiNEzNEunaHyQN75UL+JnF3vjBGcE36hDWnkksK0La6+8/qQonInq/Du9
/za2VyBELyQP6oc/2C+hY9rmpZ0qI8gpe5eBHRraZkVnjqYT+Y4nu0mTKDaStq67PDSjFTzvh/wq
nQBIF+W7+DOb40qWxH8yrGWro8AsT+lJKc0X0o2sJ/nsOQCXHZrS3JyY5kxqNX23ZhuwnYaQr5Xb
jyNSM1de0xuYajGMvFo9EjPQDwra4vbLml/8lEWcycfi9/gIHC+8OByBK1HIVgq9SzOmFLlopfBm
H6zpEO6i+HnulX1EMrIApYPdLfmysts477jFDWin++3RNzy3N0Fip9BSezMP1TyQM2RYp5w5N1EK
tAtpBHx0G4L7t2EVeCxflOx0F54XxwMOg4mQGHTGOHFAsSr9H+Db7aZfl2hrJ3NGUM/yOQEUtQwl
wX31CCvZE9PxZYrZvYQ0AJkwzB0VQ2iXXuoE7UYi2Ey7QTWkYtN88D68kjD6bTnPh8ITsc6ib/zq
7zQZSEnCCO8yBj3mkt5nHagDNIIZggSLL6zy0hewp8vCZn1GB7Gu9+lwuFo/zxVcMvRy2Hvn3TyE
Ec67J3AK8Ed4eAb1NEmoP+Q019/rIUZahNAoYZWUemveoLoF9N8BF+avoEvfOIN72tHNGNy35k6m
B2Scj3/UYx0SZCVxhsdZgOs0eJEMxtKhSjurht0sg0+q8Q6bsIK103TtTbw+5p5dP4+uvEH6mNgv
rvS/dBD8in802LmCMG6syevOdDjI9DFaxTnTqzTUYnh4WI770mepLPWGoy+ts79+SqDDlxST9niT
xwCygVvV99Ph9ZGTym+tr2n0Sgfv/mSSaDOmMmExssXNyp1tpS5W9JL1LfBpbgNlTIaNJXBcCVM0
tXHI0nwPJ/AndnK74OcA6EE0iqph/a73nzB6bw3j7zGjbfAyi9f5u7dJsKbpD1uwCz7rMVJ5H85m
khv///b5rBMEa8UozosvNS6UHx3NwLB7bCar1QeE4G1n7tIVh683svpnN12R8sYiFFxj/K9S4koT
eRE7T8upWDMUXZPWYCir0QM7Ep8GmBJMhmrxEXpzDLRVRz7E1KAilvKnazkYgPGtUtZi+PlQ8R6u
JYMgzALfoD3trh/Px1QE6A+tA3T9IhFgyqpWQ2TiXtLQ09tkcWPTqSR8FTWvEXwMgX1JTNHz7JvI
ENM3jvT/OecEn+qFoA4nF4xIYdxeLUQaaGeQQZIor5B3o30f3lMFPjzyGbtNI+YlmYUI7kXRpkNy
GumAN2U4iiEAA8W1SrEtKmvaM02VP3zzIRg0j9P3Af7IWSUv+DSutHX8MA3N/mJ2DXTVroLg9y+U
ZcFHd9CwoBWaTuN2ovryv6Lnm8s/ZasM72nRE641LmvzVj2qqWN4I//NZXbQTbO5Pjv2U6ajZL8k
okE6GnwkgCd/OS6HjMqBO8MjU7kjewJK5lkm6IwR3o3ylY2AEZX+7sjXXfqParqcnJS4x6N2qVrx
Y2xn/fux7dN3nkdj5sg/Mido40bKAC7L6jf1Ip06m8wOzCaj0eul2Tbe3icgFTnzIlwBxXDZgjUg
1TOJTW+s4nRfcn/dkv++RLnRkG0RdmQ1bp8cDOArTIhP5ZWI5KmhEKArqatFvGbfmSDD/5qU8CDU
mLECuJsytAy2ZFgI7ILt5XBIWG/f3fiokWwSIYutSXdJOCIn8SsK9O5klBpjfKr17iq2/B1yLyQ0
6gYW/cXIuOoQxz9/4duPtYeTLmjLqvAe1sCaRS0FsRmRfvJyFHQAOac80kmzMGLP3RZdJxOHjKJ+
sgmAIMsnKfki9tTgPV12oD+fZoK/ps2AFXP2BBHQTKaxZrC9dZEtYaEWgx+mEUHeb+8CZrT/HssG
IoRbNAPKJ00jLFGCiji2CLeUbdro/J5xvFiBNCDt+R/UAOS2cWKPigDbjYBvVwfBAe6mRx0+GvO5
wjtrarCrL41H/exAkKcax8epPNPaetVjQ61wwK+wlKAa2369w7CP16bIhOox2dKePj6ORGdLmjbt
tgVZ0rNlCl4kfBi5ha6sdih5cSY/cz0yG6lBujwuFDZyXtGhf816W5ajhEnEDGigZvpFdJbs9DyN
tRga3lXJpWD/KxWaTSLvPVrkM8Gh/ZOSVU4vG8dCRKKTPHtRt1NSNpXUpYgrAb491eTzpACfxrmt
RR2xNyAe8KFXVVaqWdggAZh8iFXy+KmIH11l5sA8jkrkfLKMX+L/NTkM656k76D3AqpR5zdgTSJg
IyPPYkjNQl5/uTCW6/EcurYNbnG9WyKwpIR9QPj1IMj+v0+6E9wLeE+FUYcUULKw7VGGkaFDfL0b
Rs9qg2e/xU7c3soozAI6x0COQHgqtUxwzzZJVZhdFbYK847mj1uA2Jiekk2VvsO2oVNh7ZevysOK
PTn0VRuuGUKWJyFqiybQ27luqape/duiBBeuX+XdGBWt+vcLlRs5SSP9hNbVj5TtmJXax0WZi4ZH
ZmmG7pNeHok8DgZx0/qdgTGV9fR1AlC2nOVfHDMf9boEKRt6svPhZcyJdW3YTSJ4Zungt5zt1fQL
kvIAzfPtMxuq9yyDFE+yjO/E6k3c4YxLvHddF2skkC8MAxrkNQXWANj070k6qB/JnH5sMXdrmgx8
36P3F8kz1rqLDl92J5O9Nbm19/rauIC0rsbDnDH+ZqUOlI5RkJZ0vXC5tb7gZMoCtApHWxGJn3pK
2HhHuHx26OnMV19pNvpRtWdXqeKuRpPBUzoYeMg4Dw9hZ9QpHkz3QjqdWs3pmH6UpeCwFi4gKydD
a3uSxRPxOaAl8ezHxwh5+voYgXnymuJ5HrbB7IqATblxDIO3Z3fCPmG/zaZOiYD1BJBmriWFiPEB
cYEh59Skcr1Liwo5R6zRZ/BnYJGELgnY4Pfe6yMKqBMrwQJoAXHxJhh+NBf1TMnfFe86OSox2ka5
4XftOafr0CT004QBqmjtjumpMrPHi1yE5qFlYrZSZ6SNT6TmWDAak1tDC8V4gv7BtwVvajwEiXji
PunFBr+6WQ9pqjvLaOvrLCjaAlth5sYhlEZtCHm4NQpIOy61fFJ2RLooTazq+aIHfiILljCFiPuL
W43XCKV6+ECu9M/3EnCq6wx4rS56HM2G/wHYVAgynyncuNyF53lYI/gyHH4LwvpO/M3FcDNiJbKo
vt7D72uLTyZalWf/gX7YdznsvwcTjqWID/eBD/FxmNaVsZ5FSNtzMy1SIrQ7KKUJ2ErAR42Noa5O
gnWr9SbqLu0I604C9iuQsB9OSPQY0mckyAR3jjuG+boU3AZ2oUrAY9TNEfEr1M3gSRUaZ6PqyAm1
npJkG/AotgOUQSYslr8K7AcpQlhu9K2CxbpI35jLscIcvBMWhfqJQHphRzHLl6Iu/yhFdHQW8nDs
gSjFREChn+ShylA7q0qdHo6GNM2Amo54fHthBsyFzvNZBYA0jFd0hLx/Ffppok/CywrB6gT9eRti
1o8Dr6+bk+mampvXP78pAHp1eZcU2yu8RpLqy5RZr/6xesc4vm+jqQYxQfwUipfQXdpVvfIUfWln
QKpF+eO+oQiiZxgI0nAvAptsMbyywOX7y8BV/S0GvoJhdWxkpl4K1J337V1Zcug1kbljOeTnouPU
aEtQigch8mP9abxjdkBdVJVJpJ+ooaW2Yauqury0lcN0CtKwndahkJgfjslVK3J2Vh2hXeA2iyYW
YKPeiTnNL0L0wzamgKIc+t3BGVZJ47RL1xZo3COaFP0zUTD44zO1pN7CSFPbc1Ax0GxrH8NZR+ar
LohodLxH2b5I27YLsC31iGpdoOikZbagVO9UB3HWNdIlBiTJS87h0ah/crHy8JnFe/70/bDWEnZw
9nYYUbTmFnIsTUcP43hX3f5FZjjzq0HaCEjV8wc2aaJj9sqKIbsP6xnEGHNnKMA88N6MR76xM9rL
V3wR5taYEO/3kvqIzQNbNaPyJwpoyMISi/oA+h3MwCXP0oBKFxXmA0mZBkEMyhO2Dreg6fbk7K3P
FXCDnFx7jk1VLQnmSU8fPNfz6A0hETMhSI+UEfL/Jij/AG4s3g3HomH8sPQuBvXiem+3prMmAuc+
LYHfOTWB+sz6GO9LC08G1/cSgLKXI9FpSK4Kgh02xClIgknehbp+CdWk14Eu6wf4329eWc4cx2Lz
mze4CQf4DJNzvvh/k5EUyLyXCqhEkOtMlipPSnlGIGb2RaVVQd2yKp4hbIKdLtnjcyRHEe9XAkwH
r6bHJo8B++pMAxedU25l87WRLQrbNzJCZmG0L/S7Ah/ZBR8wpLetG4fVKCljvxEJ5MIaFNZSBT+v
rD5azGy2Lb2iABHzSBw2OeHh2RYSLrRRJR/b61DW+O/6yGzT6OjwS73Wi7lLgYgN7q379IQuh0oa
jYht+J9hx2Xh7y8wDZJopk1gZiOW9QEgDk1KxSU7Zg+eCAX48ZYubBOp6c87GJFBTJNWgTvCXmdu
GcRDvpTPkcY+fWo6l2HGqH+Jk5CdXbH7OQS0a3IAV5XMlA+v81kXQ7JuLivRPrtKTRiumQwImkx2
jURqWgQu0vqb9FTJxcoboD8ERZr3EgYJnZCfFTKJYDxi6N1G6Uzyt+ShDsf6C1PUt8vc3T7HZ27t
iJGD16tEd9UYcenxGdI7KHMMI47u8s49ifNmlpdrkyuioO4ou4pBZqyXRrgAkVFcVwUY1/VuRFpx
TqA4hvb8yVAdPs4roDn8hw3EyAAluCHE6XLvRX0Acvx6b4mEWl5G0acxl0DWlf+yFjYGFP62J2Un
kOpc0a+WdWvFMP+Ht5DSgx48TnqReAL8tsyWIqr24wHmoayI1yE5af3DMsSrJptFmPB5ZxUKjmwi
yZkyHNusrd3/x+7OFRfl3y7AiOTSwkj9Z+u7z8FOT3wMeDiZh46GPRl+piOFjl5xZS1BDCa5orvr
PJgkG5BJNQAlpC0DLG5pIHdGr6OvBqxYvxKj0ffM9U+b0ezS2bl9NIvAzltaXNp7qqs1Csb2KsBZ
Orpmdh8oOkoP63EmMHaMt2S6TAHx4Q0iJ6W7QdHyRzu6EEjiqSLLL4kyYc1YwuuhY+D8IdhhmIBp
YOUvMCjYO3J1dZ9p4wtOpe0dG/B1WHLlgKvJr5UB+2ZnykZwlEgrFo+H0Ej8JtlXq6zWwrveimoL
g+F/Qms7aFFf3vcXunKCDZUdnPFEg279lHvC+cGkc/w8/rAWwYSfu5/W/b83WEax3cEjtN12NYfN
ZwZBYfyXPa+fnFwQ11uHhOiNADKB/0FLS19frrx/zcfqIPMBVTq1gc8/nt6B3nHjYfK82ahbc8qH
xVKb9xnXqR//tHXqIvivYswdm+pxf0UtNdbWCSK8ga9xrwx70677vLxltrgg6LeCULVhZuu2s5Bi
53xNK9GlB9JF1l4fVKPdj83U9K5ikZHhdNPspmrI4KN7BPv50hJf8Eyu7QoO3Qd1X7aEupYbfRvP
/8Rq/60e9j+wUUzDpALiP1bgWDtvVp32n/YOVn5+C5/hxQViHSnsu+XJan52zEW5a2UBxKIEPF9G
5Kfm5tOAT7mZcBLoJ0EJUj7pU6dmet3SUJDCE1SGCYh+8A84y5fLc80UFAictq1fy9E09e1DTJ+4
Bz/hzFBuucyeCMoMZYXojh4ftxvCtwIF0LoX3DAhnAkliDVFIIMTpbV8zwuCN427NSHPJbNNRyF4
++1ojL3DG5tUOI56/sOMFc3+F8lZV4zDfQ+9QKhujABZ58/uyRWp0K/gM+Rfna9rZ4rrw9My0HCL
JT1UxQRTEoNu+AkNO71SRmGPLaYLNreeHGvUfc+sBjnnTizPP06mVMx5D9G8mWJDyXWwr1m2d5BL
Xw0XCXgiVIokAnJvRuHoiT8CTYxjKYp8NwS0qJilIHSZsU1bgrLHA0C1oeKnDxKwhebB/1hZPvWt
hBoB/dqbXbmEJCrIsdAxH8quOOetbby2Asp4r/2uJXqy9Es1z1u6qSHieo9s1YBO0O9RJxdhGlpH
jQQr2yJV67PLTB7M6F4WLf64nOFFefPwMI4FErcspDfItW4iTwCtI86cjsFVHwAoocW7KV0n9Bd7
ViAOz+4FJA/tIBF9zvjUWeW0+IMI5uGqp1TkXxY7QiXuIrVIqo8Mqa0UdyL7mrkuPD49mUC8vDgO
zSXs5tCWoyLsnxFYjYqNQQ+JAm27HRC6fWD5zgILzWD3TXj9N/B9YvRAV8PkonxvSTNrhrrjxfVW
HxEv7A8EbhpUminSGmGQs1lReJgs31e7uM32Ucspg+u1KBO28dmkAwvhIipR2MAIdaKsQ0NmPvC1
0Jkemw+7yAtqDO3lML2WiUwmEuJJtE6pujN4RC4snMW91LM+VJarIeIioAzCrQa+obVgIcCnP0id
UTmonL91b5JfN889qedhvhJyaNzsB9HbBhNinWvBQXD0jmGLhtZUPV0W0JwDpo1896VclGlsVgV6
sVZ2X2iFLUOR8XwcbFJhSr/tmTKQm5B8NcZJqOdcWgBPXd9cAGVtC1jH2UumQBVmLW4hMKkkKphL
Wu8cNrNGgscYz9nkI78FNhMDCpK8nMmVqWsS8pCe6Ijk1q9wxtmzMXUwzEqLyYRcYasCnKWT+hLO
a+WnnxLxMWrGtC8yWkBCquCG+CU5AoDoU6dqC9pVQ5ECJ1a31tfXH93RGVllDiaTNgjfh0FjDN7M
3j8LIGw3eVymqx5Y6lZIVVYVGhD8/8mA4KEFdPlwss17WOSEU+jB/rAgahsipip7etmil3guWEPT
Ea9LbRAjGEHM04fw3i+hvr2oXdTnkt42NDU0q6zzNY1nVJODOQ8mX3zRvsKtaDZWp6EYay7Fc3QB
YlNZV/3g9xCZYfZ29O5uCZfSxiWd7ZjseWIhtrHWs2xgs9nSfD/nF2QAOee5bJI+kUReOj3Pv1O0
ElBkxC28YoX6a5I7lmoirEQ3M4Ay7jdHl75wr8hQhyWIEpckkDQ2/Vh9CnV/gQFgOSMljBlY/9oR
1oALcq1PpCAb0025JB7qjWGEXltxv8FQdl4wngMx6Ap1ndJMRlKr10ldVXjKDIy2NTRF92KDOS6B
dBovVaoloV0dfHFuR8HCmqFhh/Nx3GVUGDDzz7DUO+Bf7WTDfd11w2jUmDg8P+3k5vHGMbh1nFT1
GnhmRge61hEPxpZf3YAIOxtqN6MuNMApS/LF1gE2UbHcqXgX4xpoE+6x0VsF3qpRgoQCN8B0vnHm
JsQwV3MCzg/hjgY4x7dH+hOW2O55aKuTMdS5KvlM79lzawwXSe0E206jrvQIvAsRDVhMI4yTypHs
a5YfTS52BKftO5xq82GxG8xTqN8w3Dten42xgvM6TKSob82OnFDvZbTDoAeqzDMa3+Z95jowvjXe
5cHRQ9EwwsTPJ57ql7tzqhAg4P/Jh6viPG7+mf6r4hrkcenKneEka3JCbHEEMoqJpUWkjlJTsFbU
pU2YMndR9NaEu7H3vmF4CGXugM1tSS7e0ZXNTj4QESecaK109ZLZp66rPRGLg9x40mWZn887C5Hu
oQnGcL0C5ust625YfBZqA1LUF0JzpCzPuV3oMcXH9V3+ouKcN2gcSbHuIUPSsJY7PztYrS0TWMt9
z3yeI6/4ZH61kYhY+2zXAHf+4H78JR1TWxz2Xnd0i+OqRUooWo2vLHVObQtHVWk5LwEBX/1gNGS2
CA9YuNWrRm8mjauiWMVEvkpHGmMg+OWaO5Giml6kV7p38cRw5BM4XmwWtWgPFdELQKnvC236aAah
1oI9zQXn1ewYJY9OTo6eJErZss2/dhEJkTEKeFUDy7LNybgQmG3UGzwcFBDqGN74SBjuGihk7OrW
sde5awrAWqbQgZGx0ktglNwveAUNZXJGH6+VR1Q4pjqLq+zS36T+UIOHEjI9Xzed9n5Psubt0FF+
5FJnp55yrUfNMMTexGVeShAgoxeBKC2dzJSMT5COqYvcdrzVovqBgm1VJFmtbuiiwR0QvmWTj+bS
3oAPFo4yTOiwBcPMXpHPMtBWboB+RKf/2AjpbgRW6NT6PCFXfxLVmj1Ys074aa2aHb5C1dQh2jA+
+rgn6ZVRp3snMH4iGeavTBZSLNcNK4L0BK0BzXcqwU5C7DlS3JpJ4KPC2Thb/+VdSY4Ut0H/vCNx
mpfTXyn4KpKH/DIL2Rybb+skYs7GpTsTF8vZIVgBIhj/dW6/QJuieMRPw96xxyNYFX7PJZEzmj13
BHQ3/HH4V9dv7TWTSkXNgLDqzCvWfvObvn4BzwDsSoEHe0m2iz1RGo3TS+DJhkQt4Uv1gfmIfnNi
IetkOx3X3zBP4veSzjPhnD49QYbejtmEBETdcWNZrTcK/hMt6KBnF8ibGTuqXfMvGIHLX/pRVKIC
qb0Q06X/A+NXanM9LGrnz28JuamDjpWWz1XRk2REeNarTgVEpq0xWcv9frNG8IP6nyRUw2S53gDG
ZPqAnwnNtihDzLMdkK7f9WMzS0sCm21GhTl5gieTniB5iPfb7d6YGM7E8Ha0q8/baySJBhMtIoUY
mfYnEJiXaURu+5L9P5L16o39PutX8+X23nXj6kcHtFPJN0eZli+IuhKx8nKaOSE+CcElu44Ms3CV
ju/SVDNmIVygYuKYWRAhjp9gk8p/tJ6FSK96gmWlK3nxUfiU+012opa6iOHv67zjTJ5tlYb5g9+z
bYldMJmRAyd2jMBRaUUaHDai4N7ZnrSVMyy1s/s2tRVQ/5bdN+1YrxfRWBc1ekN0LF0vH8TsnA40
xFav/NIxnpGYPVcQD6SMYkxd4mcByMBLOlU+xX6QRbdnciI5uPoZxikBOfpMISPMbIO15HPV6Wey
XE48oxRHTblngVoYyR0+giwGzt9Vzw+44SW4aZ+IGQTm1Y+jSTrmKuXjXqO4j9CwAg7Jv//7KOrx
E/iV43BlxamPUDYL/UMGZYg7aerulpripzWTyCZbUcb3e9aWd7/vfB6jOCGq3i7o7au37hVkfJ5h
35u+YbG+TXT3FTRyb5jKpp1tHLbnVEM2AachFCpP1MTt0EzgibZZwH4x2MrjjuQvNJR8rf0zeh0b
s6BkOwXbsO3UILRTux01qhbuBX1aqMffBcxC79YxvH1bG2oltjDwuV8n6ez+/t7ChovGNp4AjlvR
tcjnpg87PqBULZpFN/EJDTXrecrNpU509Ex0GgP+4xfElYJ/bRengPG5KGUuFGUEniT7ZA269jxn
PFhZX8PjmoCPscAtFN8NH9zz9f5oaiTocXYR0CNI1asX220bEHdX+RwYBWWJGnZeGC++nlXahr2T
0FW68c/Grmywp2gGWsImFCLVyEKq4ETeNz0oyMlEpeh83G/NT2TdNqCiSjL88vHmjz/fFlWVQLhq
hkW0JczVsuvehQ0qaHdJSdhMt612abiPuzhDdTuRqyIh0XuiS0Dznsw7yqXjMf1uzXsZ8b01Lrqd
n3Fps24vTmdbk06ocS4DPQiUnVyDbTRWo++2J6Aup0n7Zpxit3xFOftQRrWZKCkB3/voIW+4MQgw
/1KOSe3Q30hEKv1PLy02QseGK1IA7CWqH8qsrO7iD4BDVAgEIT/YHvrgEaYnt0X2QSqe0SLMglhW
N9wP75BMj0oYZ9EDPt8JQZO8idTjKSn0qd3JTthVz/SUlQmZPaOvEfzyTQUR/5YmN6rMLd3ORBtw
RQtlgJIzO+oaAYu7FVLfUUtESVoJKWhmupjoXPIhog10ExBy3tfEXmGCD4rF6N/NgC5FpJdOAZAq
5H7r7TqLU/vH2Cm69lLML9e5gxAwDAc8ygKJyG0ml5sHgnm30yIGOmlZsEzoTnOl3ruq826jsk4Y
vGalurtDoUlbNGuGPz/zNYmvSzjzz8puWm9FG+rKbbXypaZ88/KRoqe3ZGESgmUZB/hqxVjKxErX
OlHQ4YtsH4aoCR1IVQriK5Vo5lAO5xpoPBN83J4m6xV+R9ztBnNL+tQf7hidmsTFkdjmbKgrFspR
rvmO2X/mS8pLqMg+LfhoKoDqgS2U7eyBDAneRuIbMzHuT1R3qmjCH3EUjb/Iiob0rvZhu74CcBRr
NGArsld4hNUXxYokLfpIgXhIAafxdjOJqVVuCbYCx7NIYvkMomhw5iNRXh3pqhpCFt8JoNvwFVwI
a7+BEPfUXCaL80AWx0y2DS/hImWTyeqlt63warmWqI2cIiPieuBbEq+x/RKbj+WvGdJwsC0+3wZs
uuDvbAa2o09aZFP/xq2DLRRVv0hmRxmgJLgleGu8sgUmim/67GMrKAn1GIm0M7WBSTs8ChF0rQuM
BqLuCf+fVpxyq1OBGXV9at6b/FHJojrUAqbrhvH8vkr3to449BG7EOK4vmlb7bLWvU36o0o5kNb9
elXmtYUeWkOUaNU8Hy35zKhFG/0IZLIoALsJ+x4QV9C6gYgB5/VQvfj0efcLdIt1AnHirAq2ZN3e
m6AY0kRXLM7pGv9CpfvVTUjwVs3Y/uX3r9FcBL2cr12IOw8fTpSi3jErRM2wNyYfBmYvzL15aeCk
9Sb0IPMVMbMEhQ/bKKMZRj4Eba708BI3RqK1VKxzLZOjey+B9gKUczZJo+IS0gAY9rruMR0ZK126
5ZHzdfOH5ahnu2hRe7ElyMHoIxh9rmSxbuUPExQAwb2h020Xe84Fo9IOtZ7Gu+k3Xizad4SkcBH8
J7Iludkq1VPvOjXuegNsXBujcwgunyuT2t274YWsrEnRj2++/2WE+d6BHA3svuHEY6BOeAO+3blb
5NpE2u0Vsd3o+KFR5tKMLAkTqbHDdGhNqpYtpdOz9eQlDD4UTc68Nh1SeKbtRWgaq/8s8AjHqeH7
A6lmV6c7oUmnt0pjIET5U6psVg/d5Q+jcmRBYAZQZkuJ1lHf51/8m24cf2fO8JJj8TZxiPTYHkTY
IKV/uy2h9s5HRU+ULu/0mF9TetdmpK+8rh42mveu2ZSNBjiwC+0gmFx8ESFxh784bCKjl6ht9U+T
vCghzd/JOxqlqOK0OELzP7KIOyLgR1BFoCOjXgP75l8EUWxaqx3H62quFQkDwyBBPfqMUwep2cZR
aDhx8kRbfJ/RRLtK+NlW8TEadLzmVYJB6xW+RfgXIA1uoGE5xSHs8VIi0WXPcDQ7Y5WAfde/DHED
n83673fW5bYa9p6QgclmYFfQaqzIUagzXWZJ7nLrn46PRFgKQGAxLxi+d0OMSzHxfDCODJfqlIze
xECIqi4nxl3GxrQgPwbzumsICun6MJJSVAAfYZhFaqbllHaFU1v0R1OEh3O0aqV7PNmjH8o/quZC
EAEGokUXzDtZ1+9552giLuyd19VH8JyQ2qwyjJy9D8KzTRxFmp5pZFQHCyRO2TYWRM31PWJUicsX
zFppisS40d7vdo7TlJRpBas9j7CuzX2JJN9XsBomRMgYDqpnIxbdnFzB2VooI2lZxphOYUetJFwr
z345Ctc0amh/hcgJYThg4NZ+5YdKzZSFTIsPnH6rKUpRu2++mFqlmVLUNY9wNEqsEv42HLUcApiN
yvDLSQcu9VnhKLszlo4gymERKnobI+InlDO0PIvrs1EUfYjtWXKdGRSON5hbYmB/awffIcB1Jnjb
qxTOp9V/sbWb8WIQE5huh7xLTODS8dyUb6+gnBw3x+1YAc6i5VVzSgSOwhIqXKSajhc7RaDRxuYO
6T0nsLdNZ1e/7Otsu9wYdO2Fgr8XNfa2bvClHYSi028AlmNo7pFvZDwbTZEcPsSFx/oijLKDvE5t
uNv/xgZBIczUyj+q72fJw1O4FanHpZ9iFrufdvu+FnZYdjj5jm/O2xrmyMqzGIrUnv3Yv53l5nKb
jDPmqjHHN2yloL3FxZ5y3WVKSLYcK3rINK31xa+Xcz7n8UmsPBju8vUBKc4VIvIwLpl5VKyO9/pU
x1im6IC4s8qNlzul7Kcq+pzsCCb+UuhSsedaQnAkM0MNOE31M2c3Tr+6kQtLKaosteg3AB6CErSm
rcTJtv8ZZEyRopZXXLGkHfNGP3/1AjtWRf7Qj4t1j5/DoAdiM+mITgM+LM+xNnoSAoPcd6+lPXGp
3OZaQW3RJyYHp89RZbLaVohG0SkyZmKQ5Ty0kzaxVgZv5C9q2V20re5WVPoh3HHf6TN5XInKjnyl
T8lA1d6d6pPvQtQSyKhewEDYNvKaIH+3S2K8eNL6cmomkKxu9+fgXvMXIahMIuH2Y1VgCGNe9Uzi
4lfWcMVxEpaCnuFLRh9tb8YHEhRlNTouk2DmS+aqfA27EWMQOTXJmK55PVpUHNMdUm+/eWyau7r1
hl+H52RYwRHEwvAE/zQpO31YLDUgPQySYBjZ1ryCGYxIlR4ssFdy09/BA5DurAytmUVjZekgrpfN
aeP9WVhuEbug67FfvEAJGaK72HLj/9riIsyl2UK1CLSEZVLU0R6i1wn2LxjVbQvWpB76hJ7NXRWK
REPX+0Zjk8oLwucbmMajkR5BcT5MCQM+DnPG2sfc5LOuhTp9wHdXnmHaLOEteaoFqHmcdITJmao1
YZlMgMlqo9mfJIhpjqn1LySItthHxBA+4M6jbktWPXBuRhzAGEPi5kFu5jRb7xH3bLKSv/q2qvLD
VHvC7al9+uQkStDInKk72Sc7SQQjlbf4zhXxYhU1sc+R0SscHSKfS0ivbaFQzoaYMpgibxM18St1
xGWfKdyS0XR2pqq/sa2vyM6S+DjEphPzj6d5l6aTljnAsEufwC0pLXkRxV2icieialdrDFnYJPzO
e4XhdwOtpOnuK8FVoTashNZS38MTEUjsUEC2qAp7YjSzh0+/7MLTk5In8mbfIOIvON1tjXlYumCh
5SJ2mk1KsElVf1nZjbwxTPM6vh06bSo88DVYKsGzVakuQAiBlaWkagdL0jTa4IuIuPYi5Ka+NWUX
WINKPJ+xfQyVqrkJIrjB6F2kviACBbnNpoWSoecronWLe/6BSHRRFDMBbUpFTBoNwGwKdPuXQcHP
Vy46X2F5jivPKM97J3fbBSZBigUDTnpu8/WaI2Oz+N1dqiywRwsZpNXSqN0siTOw0iH55zo3rGS8
7hIeZc3EzBnisbmuYrTUn6lmHJajjFHukpmlrMBsHmwTD4ojLVTPPcLAL+ZE68I0rU+eNaD5kzhR
05tGwfbAZ9A7bvmjDmA5P4h0wJSrAp5GUVk8Ok94ACJxuSNbyWtQFH1GCKDBt1M9tGCN6hxtvGWH
n0b85YzjdOhUQowd1SM0yhDWZisxSj5OZHMPDdz6bdannO3okAdpwycJ4wtAuR1/fel/1uF4+Shj
H/DTdS6RLZh8wYM/LxTYOwHL5pQGsYy6ODPxEjFRCRjnOL6PaMigSF5fV6BuutqmAq3RF06B8dqX
s8oTpuuMMYbFN4DNiRtrbfjUSQOHM+d+0qaqt858u9Lxd8nQRL34ITE47N1h2HjyZvu+QxXhkTTX
2G18wXTcoIFYFHWCMPibu2vWdmDDf1MTyRxjrudrnvIVoXZhyh1aMdFyeF4gjFgbZnr+G24GNJeY
2wQLpR7rB+wPSGAxP6ePgV5ZVAcZiGbtmBRwVIi5Z9Cjv7EEFSmKrxOzGW4Ow5Hr7iuf+5Ak8ZUY
fGBpe8szNUuBU4YG1k2552qOzASA8AyqTPQqBviLtK1V03rrTgUtUZrTagihtr/hz27tvxoUI9O5
/y/HhABk8atmWHb+ZsBdDrHkytpy5BLPAyl6Zbn0yHGN9/abbiW1+NMR9fjX8AGIzi8dB8pH2gDl
ZdIbE9RiqRposakQvrLLY76QKwKOgWllnf7CuXJ2kh3taQMtnScxp4YaJohQmczuaXgDwiRbQ6/7
zXmxJccWItatkY5kN7AIgrADQB7VZdphTZsKc+VlZXwPmMTWIAvV8wHRY3HKY+sE7vBDleJ9oevM
JYFL7yvTKGUZEonCtHdM+0xLL6FLD/WC5OiKfqba9WYv2E09/lvLQeItldlphGpgQaZEHdRjr2Tj
eRlWJz+aehslg3btdA891bWY29jRXzeizu9g3aV7fBPUIEuRj75TemkIpR+sFB7Boxziqy66h3kW
zzjCsYEvaaHayhMcHk+zogFTg6Sn9dfPmL1kRytLFcVMP8AU95ohY0eE0Ydlts1nx6rXYQDg/P0H
7YmK4DI2aYr6et88oC3z3Ul0y2BIwsomkWbdY4TtZqmBJJxw99uIFTsaVUNK3clMgbozzygkP+tY
FA6ZUhTeOHFZtg/XZFPEH/AM1abVO19ZoGtyHDY/+WwqYQ8XlS894i94G5F1Hk1yNmY3Ba8WsbmB
bmb4VjMrOt1KazcAuDDSBwatBvUq6+QH760ilMxaNZEekiCi0df48bWp6bhwPcbXUGItGbyjhjcN
tTqGaBYK5DRawfiIvbsjM46Xck6xpcrjI7aeN12zWsUttEqhGECG860GmUuMhB1QdxcAtut1X+Xu
Ki6fzJhF+3oCnv0rwBJyyhjh5GntOr9c5MnBg1VXMAe5PIvU9T8df8eYT9+vUp1kQOjABGT7tpxi
cDR9N9eTCybRH9bPIzfciHtJNjZ1PRFRAAfi6f6hT/DKF3yi2hX2qbWGMkkATKZ5LetAQ5yfRZNZ
iU/+7D98jAvuZfTkqkh3AJfW5+i38LniHZHhKSmyhttT9DSS+PVh8Q3AcEf0l4TgJZoRbzrTOvbP
FFZ0Orsc/uYlDhGIY8R+Vyv4NGj8G6EgpnGEYVVCm0YVTTV03Cv3MXc9L9IzUEvjrJR1CYwR3riX
kkx2YPmseN1k39M9zS7iwvkag0POp6XSjlAJOl+mALJNP6LdetwIJ8XBgCVCFUYcwqBc7+kR6Qcc
mkNP7T0t5DAPdfMR5fDjEyvO+z+cDZv6DJyeudiYt1fKo3Ukp7H0eswzAOyz4h8l0bs/1jqRKvdh
ob+f6GuNBMUeQmea+l4qSPnqJwO4H1iam5e/Ex2fanlWdaPeReJ5LZd9qfGJWAI52Vt9O22hrrrl
wEo9QXcSCgJYAVj4r5eB8wbkYQYFwmRFNlf02LSdbQZmqpfB6PkcwetO7Wh1tmS/j3lTCNo2dGQn
EPjVmONV3wI9tjSEma0FDBr8thJxfECcmMQFCr+4ks0bpiOLoKGGsHpKVC7r7Q7lKNpJdmSPS3sA
DvEOBwuIwYA2skq/gaQ+WdZPAGICIPZBVkRBDvCJ+SdMtf9XjZ+VGaVNCmkrkO9syQeQXjjwwsSN
lEA9c7ZO0tWrOy1lxhv0RKqsblYxxsDaLZXEqnJNHXbP9JVR7YdzepzTrxhe7N+3gi8aYQlAnXD4
9pSGTYdCNJhMjgfaA115RLvp/3NxdeJdxTFrledlkdAGWLsRgJwRTwNNAORoSqEJEcgmuCcH8soG
+VNGwiny5kmhWsJR45gd+6duOFYbSyHqd+dFfPG+R9IoVa/p/zK9aRhSmV+F1KQIiJf8uyxgr2fm
67L7X2AcSljG6mLOkVu+cT4ioK4xNbY6IU1FL++Y6aNN6Rz6V1gmRa2ckpCklP9CvTWJD2p4Nh3f
9kE6sW9yrNnLngCDL9swV4jqAAGLR3NZTgBQvldH6ohh3+04Wi8t3iL7FbB+yZ7Dryib6CjUoX+W
RrBBWD8yn1KyCBxGXMmLY6BINU1OzjEU5OVIYSxpu7fpcHLfn4Gb7vh6AFxKyt/gK0Yy5ziU4DSW
riVjj7P4/VecC/w3Gs9yiFSSrUeKznGr/3EqHjB0FA24P5LaWCRkjrEDeT1vyEgTFWjPzrc8Uz1o
IE3r2eYdCTarm59KnbOk0meO6ibDmGJ+wa6t5qG+QRLsRpFFCnr81so0C3ccXtL/MxZGzmVkxPIY
P8mDjs0Ia6usdJ/732sCyaB4MDJfgMhGb781WcMuvUwcIxy13S+Pj8WsqvvELMZhYyOfSAGpHQ69
fM/LI9eY6EkEFmyZVWEHK+GUh0FakI8xGvF/MpwYafCVYmL4FM5TPM0mdxg03TpnIZjZ6lsp0mPF
k5dLr66bE/BCUGns8VzB0hRKFy/9A11sTnFv2jdq7x42Khq4aGTWEjVGvdf5suY7XsxASfczRlQR
pmhdFHciySP3xZ1gwuNUq0lRmuDQ0No5Ed7mxyfrXjPRQP10uDXZR+C7bPUoXu5QkRRuc4dfV1b5
dLDl+ohB7F47XwRqpLCo59f2X+3ohXDoJ+dFT2rjJRCagIqYsGIL02tuU5ufhDvbFB+rrNqYPKig
TGKAwVHRYJCeWCbt+qR1jHQ3TcHWpJZG9NO0sYYo04tBPJ+96wT+LEijO0cnhsRm6vbqWlcqttbT
P9gMEM36WbNjiKpecMHgOkA9ZRSef0/C/I4jAgKpoEjDxrNdyJQIeeXCGKINs+we0Pllob81IKlP
JQHf7hy/1lIU1prYjMfU+bRRYODZpHfz4oSfC8aHgbeC2JTw6nThbnKqfQZZGivcLOy/P3G6aPuZ
fX89LvA0vTPzPjbsvyAP/YbJrIyL27n4KpGGLwc0CofwnRhVh6yQvoYi8Y4in3tGnhUvaefkTWRd
ugCilqzXnomiImz2CVdUb6GkZA2oKWFEM446xNB8xY0YlwOTeB7vA073C30EBsC0WYb5Dkt5sk70
WgdMRceEqE5uDpYKSQvj3eG8sZiwbT4QUxAj758yH3icCPq83s9LTaOlDOdMkZ3lEeotWvJC/KnT
244pgiZrkUdNhNkpULEGzRdS//QScJuWZIbvZUJsmN0vsY70h2tDbvbdllHJyAzDmxoYvdEBsjlH
z5SczallQQEt0wyci+4l6nOwgvZTMxBvr/NCRIJpoA4h3Og+l/07pSU9TlcaQfAIos7RSML5i0A1
JH+3ZH/SFYteXFOFs6N8MYvPpbI5KXK6eI/VhYeH+yOjJSep6siCHcf++HmIeEcnkO60/zN+pID/
vWp1qABrm6w2+ZEUbLDBintlNn+ZUNi0+sUJok3Tn4a8JivUOOUDL5DexKRmBPf1E4GO4ruLzjBT
0LFRrZntaCMBTIYyLbhh6G3wsG/4PIS+JiSomeSGeHfKrzIHxUAxkVlqNRWkDS3DDGfBKL0kbCyq
lGxR756f6WtdcBiEetu4utNs6c4Liq/O0iElF/lwLlU/g11PWOve/5UqstC2fdqOnUM/6FfR099z
L2mNcSQBHatQrLgU2fqQVi+gf5AHhf935AuO3pb7h4q+JqStgjQCljCojUJF28fOXFrIsV2EGKL2
IpSN2uNhhJK7fGa7W4ILDcwTZYklRFcZeAqVx+T7BrQ2Iz+CevCam57cyIRCzp8kAcgS8uMtxpjQ
UOIthy8/LwKQZ3Zk4hEFg+5+yU/nI+BTZL80mYBpNgLXgf3cZ9qWgaE0ilDF8se87Dma1UZR5Q6c
477nCCz2gaYmYA/4ZQxpj5VWhOYA5ZQ6w/fV1q5IRcrOBRnXZaJoBVX9lZPNBeLj1PF1TnG6WGiY
ffQAHk57LG/ugo5Zqho4/sh8FR/fAXhAEL4QUB+bdIcRQSeTFdQSc1xDTwgge3osjudFj/mbavWx
S+rIXt7SeI80OQ43mGWZR7rryAgkO2wBfBF9T/gT9UiiOb0u0q4QZp2rNXM6rM3G1feC5B37jXn4
6cDcy+IZsXTDftFq2DLfMYURSZPYM1Zbvg8uZJwxCduIeXZYufxpF2bXTXke/vINExOgmv3JuD/D
2oPztbxluZNAXjJ2WdIyP0uJRPSc9LCRCey5DarYFLUPlZwu7SQKy1fRVGZ1/wLl4Mh4PvtLxezS
RXx5q2l8kkxg7ufmWk8qTwBuejigLwHgWuxgfdPztguO06PNz4uRt6U6sucfw1hrQSoznRgDusKn
ZaRSQ0kexV4KHeSyxLzhSOr+M3xPN/2I3H+faxre87y7oVpNQPhiUzQXV6sKDLURJh6It3tPB0dK
Wln6tWISnOA31TizM1EtRP2VBZf279CdgE3oiILy+6NzWVS6Lgh7+VDgbWRkogSYJzQg9oOc1vSO
QtTtEPmyskHBTB/LNtNjsokYpvIr79aMmw7rvqU/7pGwVe6iluQioS74o1jfWdsQO4FYs3ZGT1sg
xFIdvUc/AEplqwwGAEXFUEELBMNx+LVsfBCdMoNYVtULBj7u1fqzN1ZRen9WL+yKxlzipFOVmU6U
SUmPvxwJWq9RcvK+HenndbxO/GseSoTSWJ/rBNbbG/JQmPt8S724uL5ZEOjunax9qC/wU2kCo9Fn
ziILHZRrEpXzvzHCG7Ue8dnVqjwqvC0JRqOAmW2wIsWmo8glthFZ8L/aBSxQgml/c62COc7AjadJ
e8ofczxJrGHc4B4ZnNnVt965vPC5ibBfmp/ReYCAks7d/YSpmVQzjBAwA3N2eQd4MCBv9OVynGRe
s+mgG0vtMa2uoUTXgOKVYcfo5FST4hfSPf/tJOzgQNTuWRtiUDzojN1gPwEfPiOq5XPxbmMIOjOl
GXygqkhb+r+r6srHiOwtVIL0htSpkIt7hDwWrfy4YKWwlLsSfUmPOEpE814rGWsV2QgLKPxCA1N3
hgejo3LLqkzrD9vuW2uG+TxJrsgu0Pt7e2QUlTyeDnmDxYoHHgqUYedGRlM5gVlrg2H8ndp46V82
mkL2qygs8RY6ZBgUOYG6KmeyWat5yfPkFig3M5NxFOpFWdRpusMdSgaQNvV0ZTwk5B5uoyLkTc0N
jtIKGPODjd6xxEwW1v4nbT1p/o42p8bMEGapXVsy0VmC+V3ELlo15x6UOMV3YkJAF8uF6wuA+CXe
Qj19VK2T+EPe1bVTwVnfq1xYxWen+9k52x+B3+sMf1+OrFyoC1eQVZxJNnof7rSSx5E874kTSYRv
Nhh0Podz2xw3e9EADt+Q/UXnEI1VJsE/yRoF4S2HV2SvxgQG8l2Vd4mhsJO5WaQQF6CiBrkJ1mhD
W6FXFF0TN8qCSzO8krGxXBLlp+bbComrBdO6HRw7I+R1QLa8WUeLtXOe4rfYFziybxaS6twbmKV/
VsIO0kuXGoqDIjRYTvZGiNcMWTRNoc5W2sJxYnVfc5U/4B6tALzhscT0hx2cosYKK8D7/AQxlRnN
1fp928XJ5GyoTnvQiiZV04v5xMDwdKmAShWc3GBZla90qF2uYrTxsf+mhkEb+v9SnpvfxSYWskHh
npHv32RM+XPFlu0RhPk3z7sEpXbiUAa99JIP8wPlyeB38CWnCjedMe1b7GFTlfASPaF8lf4e0qpK
awvUg9dMK2SwawJ04qRHXRqKNKHiJnLyLlLfSSKdUp8zJ35e7do/95hGsKv6c3PcSY+ct0tU353S
D+RApFEmft/fnaal8VKmVvCodz6NfWxr/m/di6G6Lg4+uwuZWiZe4q4IfWK0Gz4X+LaqYE9rlc2W
CaZMvIMmghdR/lUNVFQL3Qh0xcJI7TDpPcMf7r/FK5kK2Lwi9acIasKaAbjprcJ1lVwU0pWMIiJz
FGIdshEN9UIOcZxtuXcnK+gpWz/ete/kpeIs0zrUp/lnh5pva6pwhN0UzOSVAegTyWcGlFDvCbnM
PT1FRhdxTSLRYTNWl/+JkyDOM+YlzuBqHca6c9/ZzOiLIE4SSc1Qf27LkUROEbgld92qGlAGk2a7
+jaODF0Hil48OjCupx4iTksQ9gzCCVMmRZWrAKfni9CbHG6NYdtAhpFu6iiM8yYzJ7MXNvptK2Po
xMHXLk64yZdej5Dr89Ub8Dzo9cekfhsE6tTnGQah1qwKEyS7tbNwABwSxoOsuUrNL/yBnAB1HB9W
D/jUELNo08JrQ8SQ25codJfCQwd8V3QPN3Oxytek+sf1m0R425W9CMrQwU4cnEZaz/M1YH3yj4IU
7x1ZyHh1ZTOr6Ce/4MhykLzpFMVd9WFaaoy4/VNabxRhI5M29w+BQ1saHRtX+jvAsakTgwRe8nGV
DSJvi9yI69Ca0JMkniQtJGqzcu1FCJx+8TYNWUvN+2bF03UL5Kc20qjtw9YFhDqghrTevEtHdLKh
wsYR1AwWmgC1Glkr98lbPmROS6wZIfcxrrpwb9Wk8m3E6M2+tT3fWA3MbAayvqyrhuL3mDvpoOQM
rupHWDu5PKUaNo6t3TjZQsGZKb6SJ68ixQ3APv17PGJjvH/64Hm0E9P3nkUiym7TZ4EjbVM5a4Vg
NlXPNn0N3q6dnB54znpPFtokTL0GhtM+kKPYhZ69bj2w+u2YX2xhv8AnGq0ULTXIsW3JB53a0Ptv
DF9iODFG9jWoq4vikJsRvRiV4CLCOdiF70jXEEm8lSxZa53PHHliwnhGzxTqR2b7T/UxPY5CCREk
/u/poz8M9IF2U9DQJ0SjwvWopY7ASB0dmCGbqv4kluI70smOp6YqNFapG5ksv+769MKW5EH6pfsE
ojpQ5C3JXCcZVfbBuGdOFGDjg0SPnZRvvYugv5+8NwXkUVHazZuADq4aS6mcvmlhpiyHjlKN/p++
nMzFx8Q4lxGC+xQVo4MHh6Fneat3QMAZir5GJSgKVewt9tha71PTssgijBBvwMUEO0+jA3vTrKOe
HDK6JdY8zL+ItlLZsOlgVWlLlyXJZnIkpE2N2RZBOXUSeW6sZNNED1bspRd4PfpTK/OWDn6bX+2n
dJVWXDvG3BPJYaVViO0PMo93yDiqXrALnPeZKiIHrzeP+Ui+sDcShrfFZ4DzTJCpXwoAplzs8xI1
wPC3zuuyd+wT27MN/aBIvjftP5xNlSsGcQxcGt+yVw7VfCN/9UIOhrL/aStdAd7+uObn+KT00q9S
zqPMvz4Y5Gm/d4AMcsNAjfm+SKfGRyOCUmgv+gW4vR5Q81OtFbijvB8fiMehDHanMyqjA6qrewnS
4XznWCjwSKruYy4HvJFXe/ewKhir84MLsj9xheDWegx31/EZvE3EKGlgcVH98ht908y5oi4z22GC
e3yZVUmoYrjXyc/tJoML2NlGf1qh6K+IvvbZgkt0jrh2f1LG8AOwa+N1ZosatKXEOmO++j8aUZS2
59bRFyPZfDS8NMZPTI2vKm4tcXFYYXxOyklGzLQ5u8oc2Aft8H9dgSAloJoLLcOuXsYOYFqiWMuQ
ZGvNdOWteNJwoBDkoi7hPjaAHFwAntltsc14p7fQ59ZJRTxyJlUIgBkbJhKzqPv2XM+GikaQ1DlJ
TppgAEktgU2/oxFaTQhpEenkXNZGcYHMmRng+e6Lq2hwxKZUml5v3apwmzLDDhLqCRKvYUR6BvE1
gm0pHTeS/2++h1rM+30ctviIdkWRtL1rxNXAsPcfxEmmfyfbHrdwVFJnLAY9QxhMV57+r7rP6ivR
Svtvn7Ra9bqpWzxXpEWVjVe1Ih/Zb+UrZfl2vEd2DmUmCC+O0ItzPxBKdni4SZLfW5pZpuLBmE3t
FguqupDnHmOQASYgS9qudmv9RH9eqQPNu8bBpOYDXjPaD/nhSWKdSo/ve3TQsg8PaFM8yd/r2yL6
6JM53/VHuYp6/qBzlGaNoONBRkRj4tYGEue6v+DGJyUbp32AJEMDWZkmeHfiPEFMd+viB8Cv4q9J
D2EBMfrSqqXD9qlL01i/7Ti+aHyYM3Vy3XzngWV3IIM3SbM4BwzO2YxDJylR0aHEXS14eHKdHk4n
P6JeXAVBiBlCNm7KcacVRb2w0ZprthjS43FDmTkCLswuxFL3OFg5EozGszUstDZ2/Lk4Xi25zZxI
etyAvNBgg7GuTuYlRA32huIVnLIfHtq7CuAsAM2ooIvbbQl3RZc6lUsfHiQwqZfaD0aMfxSPuAGl
sgu3nH5Z7aMQeyE94hcl7UmwmgJLPiFedq5Ofk3MFRc/XOXWavXJ+3sZbpN34C/2dgprJCZ274O1
FRYJ02JoeH/HGQbhi7rpaUypZ3I1o7bzRerieDIaA42GTtqdgVZkH7tLHp+aVt5yC7a0/4XJ57i6
/E5fVLDA3jUyJzJh2oyvFP/rqLrcc3KdAByZ2fWJglrtf9SToGgEKhnjy0uw3d3TdY4k+EO8ckYA
ncGvU8V5vwAW2vbW7A8jpx1wDDifQSrxsGhFrGkWKsl2nMQh4hylXRecdDIAjiGp44yThBKb1/4Y
JL3Cg0oFDru+EaYrE+D3DzW8foAQJtb8qtm3m8pgDn8J4hr9Yp1+SxYIwdfikeWgLs6gyyPYCQT3
djlQmGIf14a/3tJTHwWArK+WEvwjH52Xiu75KdvK2z/HCEnyQRAK68RkBRSpjNTSXvDHKXBVV9pv
lO03wnNodeN/0gROYlG/PdXirvs4bbE2yozqukoFA5ZJ+APJOWNyfwd1iBXfy5y9r/ImgNCYQhDQ
if+ypj73uNdvafDjho9RQSARFFryL9aS2OkNQwqJKUgV56O2LC61UJBs+TPQtTD1VCbBPlfh3gbK
kERKCKtnTBdXeo1i3da49LbrYGx0guwHE9u1Vxhw2Ok9PC9F2L34MKSGvrj23P9zGMdfagT3xWfG
8BRaCZBdmw0027B48mNcSvFnJgcw9ClZBTCl2sW72Q8Do901nAAvk5KjAX33mXEDPsdlHzw1XQnF
7MfpMf/Djk/SvLxkFHHQqrtetensSTVvCve8xIJBzMXIlSW5OGx+ETnprF0FaSLIBxkqxuTEyQwP
aqpdY8l92sg+hw38eAxFiD4cX4twtltA0ZUX7ylkbqrO6kdfB/HZg+sjWkUXqzXrcZFhkJVKQ2Ok
8hJc0SiQSDFMq/9J1vEPAEdFiP+2j1RhuOoSnEmfefoGxw+JLQR37If2I3POrNwjPm4FV1yYxB8s
pfhyNInLPQDoc171fzuInSBImq1K52AbFNs8r0wE05LmzmcLcGq3k0Fj0qqokLEB0Pna72Aa8skU
m7K8M3lBTgG0rRJRR1MHBc/0wZEagGN2Nijix9zPfPT7IHv3QjmqBGUH2rSCdwOfUP1zUYX0rE9/
kXYDC2YbuDDOIBtBbisDk6F7hU4YIXv+45dsSa33gtM/L6g3BMZ036Tg4uC/HajBngv0XHWBsYFe
+vfuBhrpYzcdOu7x4PXU/zYVoX7pVEmeHxJLMlXh7KyoJa9rZlQrSiU7s7Gzl3VdpRn2MFgGbgRw
uf9iIOIwMxYTX7zXsF0qhZ9YpwMRm1f0yzIlTz9D0OAsBfg8uQoDrhnPfwLrohT/eCdH2P16gsyX
ynXf3xwFOhbQmtV218m61jZNkOMlr8s2Eyt7b5ChifYmaXPTqAkLx765+76o+nAgvGa8FFoBGNg/
F8YfaYvxNBzQ4Px6zZCouDug4BkVQ2HuLwA4JWR8mTp3N6XMdcMBH+SP4HMBuZ3SD24cCYpvhRkW
MK/4Ut7lgP/qn54qv6pGLfGUfXM2nroYjiAOQ8SaH483OYh0qyuQIZFD9Z+T6+KuIAfVv39rdy44
mw1Ve0m6hnVpVr0cLoPiIw1vrCSKthhpZcQGzaIeef1my1qtgjsazDQo0THSCiqPByyM8xMUKhnn
cQUbCZDyxSTh7AkugHVyMVO3qyP3V9/vfy60d0Cl57HUMJyH6hc4eWfTuue7g8mpXhiIX+UhU+XC
Onc82GsoJGTWrmKMW07T3eE25o9EaIJaK35GeX9nUclLY5sUdqQCWp8+L6KssQShlf9uD8zlMdFi
rBFS6+SCVCGUWBKV5kb/cfIROTMkne5Pfah3RSB11nz0RIp2bKflbDG43WH81fuRAalgkKCOoB39
a37pAhWqWh8y93pEurwZaCzlC2WWlddDpXiazEAIo3SkmxZo68630Tp0
`pragma protect end_protected
