// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:14 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
a7X94168DzRE/oCn361sm6LBecU8BcrL6fZ0eWtHFfOyV3g+z4hJBFbnt6jH2MDJ
3xUtaifU0T8ln9L9MjkdAgd681tZjwF7XoNsxJcJ8f7s2Dx2uKmQFEVr6fj56WRI
fHrMZHTDg0F07xcuu9ica7IWGtl7530Pb341hf5DhHE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30400)
brK9g6dXIMqf75q5p4g+yJesFmkaCQStmJj+/JnoPaIsUzxJpRubBY7RTrhee6oh
C9v9IZCFdKPLGxxrbFpFjDE7ZkJr0H297bYqS7jXLfoGgGae67mD4ukQMUwXiJ9z
SBxQ34G0jlnOTh0Ot6Dd7EjqaRvIP8uSSrmM+QEVAl7+uoOjSGbVDLJvso19LYVn
yVMAQPKpkfI6KZNmkQkncXuehiJfKdQ9Xgj+51uvWFPEWUEHX3nEACTzIhbvORue
mRckN2NY0rInilWl/o/saJJqIwcdAZ3V4hStbx5itWBAm/0An+3KpRvRZdwzUn/F
YSnQ6VFfzg8cJUiM42RA8jAAVnJ0m1DFRjG6pcrbHh+dAFIlcK9Kh6kMozapUq9Z
T7XbCOzW7CaKbaq2wQf+TU5BOV2Yesnj/4pWkOjb5nY12g4Epl3otU8SU/+Fkd/4
VssehbBYCz9fEEyQOhar6M/sSYj4QaVEGyYNtPIjze1jXXpIoVoWGNYs11Gnnm1C
m+sRRkwY3Zd1qFoeVCowsQvkEYJv+H/2idrKWFobNwvlgb0tQ8Rx7qCaSMY7KKr8
L/wdFYaOlHjRedRttU6WI2XmbOHoB3LQBWVKJlLv9LKxtWVRHP34CumnOTxFt8w/
n/RXTmXtrCHqPYzeo1MfoD1CA4GXvHyh1+RIy6uho3dA3Q2Dqz84LHiPc8YwsO1s
qVT0uQfLoYMCRgi6uGd2vofLuO/5F/dhleqqqts9R79jtTXHHPRCJDN3IRUb1LsY
6KJz9Z2H8sdDPvW2pnq2gxAAL9Wq90MY4BTS291roaIEJzc/hGdiFXQlCJavvaO+
h844XRIgSlCBVpI9Y1QoGXhhvaA053/iP4DSCZ57yIA5dWQHA4ximxxn793vmT3F
y22kZRyJpaNm79QRKB6pUdhNvhuXdrFSKCRH9sjTzQe/cjDT6FNrCt6wgNj9LeMJ
AcuKM0xENRPZsSNHdvpOKnNVTZcWo31vsAfLMAiAKxjY22+alt4AhqsnbFnMYyhG
pWbc7cCqVIRgM6UazbfGs2lwGzuMaL32LHei8VU2dP2d5VyrAHNilAWkI4XV48cS
yWTGzntU+JCiACV7Kc3xzJiqSDxQE+oX80m6XDAW+ln3nHxWGKNFVUpL45dO+1yy
m5wSmTEdfTR9XBledVfgOFwEXBaBuQsOXEL1I4lL/EZutk1cdojLxNGTCmh0/cPN
DI/ebpehnoU6awqYP5uKVM76H+wzsnJYahdHQkxlVtg6coJnXQNw+JmKWMIGxehU
ARCGODXMoZcNBjfKcz7/oLciDfP1+WZ0Z/L01GlBMjZ3CG/aLo2MevLjpFmO4AAP
C6frvPF7qQPYrQiUccykA+bx632413axYDAC5oEXZWflB7mhiEw05AekOUg89tiE
ID8U/Cn+uWy0OFhuEzp80Ri6Rh5qpDy19AyWXS7vA7rcpATsJFK0Jo/4QQGrSEuw
8ilUSekpLPW+VdPYXeGUVkqs1mhfFlshggfriwA1trcv3jL4rXvWcyJivh9w5Fsf
j226Pb7InoU4e/s0YpEiRjQnv9/oUQaPYxa3LN9L9C3w+Pj7CH1KX1LM74V1Tvws
3igku8Ax4rk1Hv+Ud4egnqKCJzsSd1rJkT601Vmd0Dj+MEwoJpD9ccIZaZxGEjPL
+lwDS81it6xCNipKPI9ckkf0iPUNgmvYfxAqmQg4SzAWN7R4m39gRX8IDB7P/5t7
0Z/BHVyMTq/XUvx/XLbe2LCdfFJ7AXmQcedu4drYhCqtkNFNqshwt925NdCoN6pY
b1zJN9+TpKvzRV3uE/0wc/WqurlndNWii7owg/rcoB0D3cLgMdF7yFfRZXyiv6ie
r8TF8qFuUYAp8paN0BXmFS1TclaBVhdbcoKE8fRmpQHPv0fqMJVLdj9sjPkpHYp3
2xjdzrI74xBb4BOTDLNpRWJZzQD0mcDdQkOQ+9bqo3f1ffxrUcCJ08wj1Qf7GJEL
y4L6+nuV2e+BeOauM1Dc4dRHLuX2xgzbzgmc1yH9aYfRF0acsmu5jSv6a9+/qg8Q
hib9YH5HARePrm3SIGVWE2s3rX6Wa4rKEtT6c0UzLiTaR63uLC5n/KXo6AsOvcNm
YjS6vsuH+Nk7mFmhaH3mgf+WkngL1r+4TKKzSf13KY3kdhnBda6E+64cQlLQ7KSf
Py4OyCCM6P41kJukWWIlhTx7WLuQb99fwtsnceub6DZeFhs19Z6IeU7nrf7AQepk
6b7CAK+BwmMrQkzWMdA9LJjvHMCsRfajiiHArMklLTM519VNGXmhaMSPaOtBnXRp
kiUdzBwUkMljI8ZHVjFxeWFiMQUw98kqD1QjDZJwYE0bn8wRzwotWZ2kKk0MGkCP
9CjgBZgmrWcS0IqQlvbR9UmtjQgmXnAHvlMq7t0nOL4ikbEPXJ0LxVDggIOpMogT
MiEJUW0aRfBBeP0EdRgrtkH62xF9hana8gJ0OIDblsNwgsAo3nRRPQCgsT8swV6H
IZPKTP0hRXpLXrILs64Euzr0402tzAvDuQFsC8fyNqKLrM9RFB7UdK9pKDsq/ur4
SChOP8mRudx7tTocad2uB0JT0hm04h3YedyIIYf8A9LgtN4/rw1YCn8NusoW9WeN
PE+aNAOkDBbv/nFw3lXGBmQieVRtDK85VfdShWPr7JBBxzYfODTkh4PX0R7TJwE7
t4D89W0DJakmpkRKo0U7yc9Dup9+Anf2KOZ54dKK7S9PPc2nMx3uJamTC1rn7o3o
EP4tJl5N/8dQ3Xn6pn+JpesEm2yxJeAgNy3DsXfyQMtFA4yW9DayzOnp+hFelS2b
OmOv/tJW/6kG2D8Pg1jfLG0YyLoGi2iMPWeomQDtDgSYhpcsyL2g5lBB0NmjeFCC
Xw5kYqE/I+6tb07Y+YOAUkC6uXd/FHQMOb2uyyRIRcnHge4egYpFKD4m8ycGvyaB
LxPEbVW8AW5sOwKq0ffaxMLo+ryxgFFwsfKgAroG7Xmevo1ReJjXS/DDGVK6X3lz
oDaCEp5/GTtF+0cz6NXuG+AJLxK9piJTLU2DuW9q+QoFMYqf5wpTfGvaoFPvvqvD
N0p6PO4KIO6IQ3sKCCQEMLkiZlzW0OZVwgcQSX8twphUps7zbsq9fbhskh08yiUM
D725hM9zvEbFxunxGtocfi14oviohLO2xuEwiAPA6f37bL6bavVMxg4fGIY9o+AX
II14Z1KcsW83czBGfhUCOlD0mJ/KNSYXWcGpEoAqv18UzqotKIjN3t9ZuGZSXj/L
RaayHLGkDNpL4N3JS8TYJ6HuoZrL0S+Nua99X+kOHViYnDiqbqIc/xWDuxlCjkYO
WijDYKRSAHnv3ydjrSYNjQQzHEiK9dlQ4B2DJ+6e+gxwx+qXXK9eG8APWfFzlStd
DEC/7UeAo9OxMFnOQw+PvhZaKuQxd7TivYJQiDQqzmHpKxaFihDphvJwEMKuqZGG
dTbJAGKyAWz6SwBZGIG61HrhsxmQfW2le50ajQV9Bihw6K+CAmt2Ih7elnetdKVc
l7MbDjvJtgwRAAtvFSYIvJ2TcYN+H2VtjGAgmctam3HVZ65QKbv1rCQKuZpIjCSW
dXPL84iZr+sSCpoMPjZQ2JhDv11sXYrNDxbKSDhTb+gYxajbYrem8crLsxOTo1SP
mo8mojHxHohj+rjjtttMigB/U4v4tcF+x2YZ3uUkpqUtvgzWed1WU2dW0iniADu6
NI58MIUiefZDJSlN8zXu0nj8i1+bjzGcBdna3V9peaCfDGPA2qJyrqLrIolMJdy4
R5nep7gfgk6+klUGOdlqfj3M1iW+8XNOzcxr47GJvWonc9DJJF9s2V6x4khGWgEx
Ndqgy4piz5UONF7kamA9ZkDg3OEZSz/kHut0b4btXKaJPW1Tr3H2U3ZztlGVfES9
e0P1J/7PNAvBcfTy+mMyFG7wRAaR0iC8QAnjcZJVRXawUeqU5GXMmlW5cYXx6c2C
bnxbdxkr60DMucYL4Dk5lLwbqg8ehDILI9tFCg8KS2+5U/9lNxueWXiT/i3rL8CM
KViRWdB5yx+HvbsuU+SWsnhkUubIJdlTa/7jB59t2UA9OxMsnSvYd/FZEdiuq0OL
M2/Ik6xtPSwz1v/rBe/BhnCBkUjMj48STA83aSMQFzJ52x7ymSqv/ks3QRfG0LSm
h5FqahDMQ6/El8qCoCxUgg0/GdKj+HFs+EqcjcZSMHD0KF5VQAziI8SmGjykuntd
Q1f3Hf+3hfPecuhK/I4CCSfYH7zgHTzv12IafKG35svy3yHdMyP3lxQmoqmxhoVS
Mahi5uYycsQnt4sfMasjoiTEBw7WugBczGpzZt6LqJpr8uA6UI2fmmpvAkKJD593
DX20tNyl70j0leJbNYt5YhyHA4uOsuYoOhaBzgFSNy4ofTeKr97XrzQ/7Otx67f5
GS6i6Th7purcz5lIZQU7obcmQjnhYZi1+PUjeM8IakBZ2IqPtKTnUlhgcTrc2Ogl
9+x6Rv0+rEhABqNTqLmSYU+HR/VABw1tpe3yaDi6yL3pMimsQIZUWqXyCS1MZzTO
ESdiK36tBmdUG7oBVFzI4RaIf2E65vd1Wx4V6nIJs8NBTwdibNkVJvDAYYnYh26b
+PNSoLIzSsAAvToYUp9RGCy/PO9cCfkJw0Ct2KXlZdpO0oo3bu4uWnD+2u//tpfZ
yVgOeXs0sQXU3Xd9xDBBWL2Sckw5zwWtW4p6jEiXjMTT9XSSiORvfryMQt4SREQC
tCDR0r32g6pl+OR19Eu8oWb9aC9oXVEjzQSBOX1KlFUIPSZE4FrBoo8Yi7EHZZ4D
awIfVFwR+fFhUbi4QPMevIiL/26DckEzyWeFljWrZF8/9wtJ5wrPygE/xRESZvIg
4iWcZ/1dN1HMyyMQtPf+KsvhrvCO/70DkJ8iJFaXlHc5eOzsb1EjFuz+aRW0TMWK
E9TOgmOqBfgh0mZ4vBqIh/J43X+E6pkSpot41cZARr5xUo5u2Ir3qsef6+OegNXG
dyq3ayqY8/YpbMBWW3MYG0KbJHib0I1l3XrVe9mY0Fw2fkDWZYCqNEmcip99jroO
99iJeuD9MjFg2Ubro4AtY3qQ4zDkTHe1btLvQzmSZe4tOfpqZ1P33VHZxVCZvclD
xJ+eBPNxzOwLrkXbbYFNbYVL7tZR0SuEG/RVYrRN+Hqt2Y+U3gNAnAE+xkhLWdMJ
gqNBNypOzZqNCJSrwJF3ZR9eqyxDE7RGOgirGIsy+Qa+CGkFjw1Wiejw4Hq8/cSG
rM+chzHYyOOUD4wZKtDrCtPM9nSayvANkMqa/qUWcjfVjvdJCRjS3arubRpBknPV
Odv/iykM85U2g18vvvDq1eGkzvQsfk5LtI4xx6gzjzjJg/hX0zxScE0uNA+NDt/8
qEXeHS6ibDUY9PNpyfb47KiYBN57MGTkbCPvHEmiqRp3T106olH3cvC9URGT9dPd
nKwz1RZPHZP6p8n69CJMv/eCSMqPBLR9r/IQUwH+dv6heAdLYJP9XfGVsUrlx1Nt
mc0oVga5j3uJx8UUbREzYaQ2Kws3HcYETAc8euCXiYVeBpCoiBsQbqW2RyDe/W6O
55yZbRv1vTtTYNErocN8ntr35E56Xk+p34BqcPgXi7UxdkZCqURPZOHrdBoF7PBP
lecS1HrYkrI/aXdHz8bVhG0e0h92lFqgaWkbkeLWScDC16OPLot0/7a2KcklxS0R
bMXeuJmPu7nnLJoTjb3r1Mhji82ALnNsQ3T3P9t5Wjhg/Jl0kL39fDxpvPik1ot6
hi43+/uKMxOBwYFONhE6bPx3eSHtTfrO8ZSyD3Ng21tVE9DO/xM0fWMyNbLy197B
5doSt8ymXO0c2fr4bsasLKmxPWpNh7iaWuFyCP+T6XIDmiXap+rjPWy/jjuS/uYG
iAV/RudznbgKXSPYQDDU8I7wmQmc5aZUzCXAX+IbPcuNlzg9jxpDc45RUDxHR/WQ
CQE8qQ3Sj7VyHL4PuppWDhjU48BHX+TLFFVgJHy22Vq+ymeXfVmN+/CxNpC+zB8w
bZI6oTij9+xYBcEabcfIs/lAyMtsNU8pJovtbjIVd3zlKGvLfP/unqC5biQETLl3
k/s9+c4kEccbkbvJQjlgmo5B6iks2mUy/BJ54aQI4N/MyHDB8W3kXY2a+FLulr4K
ZCmKvW+r/d6FPdkConbQTn7Uc4DhcUmbGn+Z20lrza0SXoFer830RlgXkLhVVBs3
urkXbNfpqFndHij+QdS3M7sw80u3o98EnFneaJho0wG9ExrpNAHBbpNxAWjzdGeH
Q4BNTKJr3+roheaPAZiXzKLGHlBwy9rYLjNNJLVSmZURNtEm/FrwyNJh6hplzw8E
4f71JvM2uoj4UJ102VCbh60wHLE0xQp/BZOSxh3AWeNc6W8C5/n2OJfjQgE2i4q6
NplhsRSMgQeTxAnbtXkLck177PDcxu45d9yP51SMTy2xmmJWSDbNBdHokdTpKD7r
WReEa66vQMYCF5CxQcD0Hf594C5Nwy9bNT6O42sTygD0bfnEgVH3ij3d9c0hui8T
KaemDNcisFWxBf6WZN0OaoVqR6HcDQCAKFEHEl8d/mhdK3ZRsd6sZ1Tn/ZkSlejY
BgMefV0+hr8sdEjvCM7FWianElNUYHE4TKGRfF0cp+d/OOZI4LgQlGduVTzdmccG
a0n2kAqyCbTWQCUP5e+VFcTyz+/kDZev+tM70Ax9XIruqqzTSyRI/9c2LkzCGxVY
9dyCuqrXa9KT9fhAnLyydewv9Z9N9RDEnYLUSQ/lKYtM7X4FZRN0xsIQjHgtEkvx
usQAOOz37RLo9ANssnGSzFJM3ceqk3qNtjmK+dwWhOamfShLltWUKl96xXoFEoBB
lbIjpaDr+/W9XOjS1wQU832YjB+dcjIjqb1QmD6VJzoZ5UEhU60YEQOMGXyc37yo
RUtUQm/9lLy5SCPy1PDUfLDVCePXOOYnA6/m3tTaeTTRxdY+Bl2jxQ8MHpg4c8tt
ZlFBpsKnCpF55yj3a/1k8EI2G4t6B/vheXXl25feyjscE/rhgSfRWEZHdMMXhDm8
do1cTbn6HifHWDuQjQh6sZCm/54VeTrBnB9I9th1EmqcElplJWPyvTr87OfQaxLM
szW70L2qx8OykzzoNap4vznzPOz4U5xUn3h+2BsTVGel6sPeVV1EVY/f2vHx1HC4
B8zHj/aKgURROhJpx0qa/prsf9KgyZFrAVWzRbtFNdL1ejQ7YIwOkBG3fc4AN03c
AZvG0/u7kc7dBF5MtuMmGox8Kecrfn8z384MlQ7b7dijSeynQSoOIT6zxgbEmKMt
eKp+9vekZ3nME2yynd0tXLuJQDRnxf3pzVXQcDbrcTwaH6H5a/pdoqhOBpVjqfJS
TS6U/FXX7xvdXRRMZiF7Qjmqikwja4TvwiNoKLvQUadKSiVNae1vfXNP7c8AXLgK
+VPINJtNchDV7ucD3pl28kYNXLdzP2yq1BEh3fzZaz9CPYjbDptDEhP/Ghisyyx7
VAZVUZ50yt5z6E/2MDa+x8vWQWooJBDIHetRmnGKsj2hGKCHjbip87Cmxr1Wq2EB
dbfeZxe3Dzlr7hNkcsT3uphRpxsgUqlLKh7ODF/FFlMrCI44qlCqPIzSl+0GP8VM
Q1yaQLsyUZc/ZaQwR9i9s2RARzklgcgKJUUtoGYBKSB2/FfCXL7yKeRGzQvmqDmh
w0NGhD3IF7YlnWtKRHE1HxwjtQiHLw/v/M0B3GUnzanNyeqqw2MdC8NUY+E+CUs3
ZSxEiUUqZ0vizknWOEg0Oh3KoWE/QyV4OEth/IA9L3MaHJifcARSsxOLYI1HeZo2
sqnSND/P1f+oXpLjhX/XEKYc4+m+Tula0rXcOU2yQlNBRRF8iCdNGRk/aB2+oYky
feecG7RT13EYsYFMw6/ss0kJyc7M4DzVE0lmiqn6Oowi/5ae90yPRhFuKCz1BhcS
ShdHDPhyZseM6q2c1qjzCacL8LwQexecX3zaI33hYG+z5MNkniXBM9Su436wuG1Z
6dSrtk4gOBYBdlmGIbtmqnvwlBsAMp26OWEW3RL60mWDpFVCzGAHrKZefcllKdBx
lzEFhnyNkEBD0Pb4JU23H9c3+WHrIK6yy36zYHHUlhocQue+Msk+LJ+kKjAYim1O
PefiVuBHpOsdbSYE4hkcw1jZZoqGX51jCp0VC73Yfb2nMP5fX6LqRGzADJjPoyDO
vRada+pwJbSNAyzr/OFQF4rTpuRkicZRIEHp5f91hqNl6mGLsBVEsmq+JsCeKXfE
fl2EmkPJp2jz0dfjZEP+Knmt7JQ/OF4wBM7uSEryQBzm5acdPTq2B/UpttYF5k4r
uNrEfVckJykFuaHTSXX+ZnOCmz1mhcEBNnvJavCp2g01zYcbtqm7AVGilqBXlK0K
GaWRVdavw1DcAi9kNrWRHno6Go5d954A4QYFepeNlEYiFieHXK9VrsJGcR4TR88f
dNPIZq4XfoNTzTUdhhXSPTK20aJqDo03zKd4AacA7VD4XCfp7kHHFSgZOz8VMlBd
pZEhyAUZLyBbIM/GeEkOdJ+JUEJfvLFxamOMOrx0pb+LEwGCBRef1+sXgKx/UX28
69pHsZJXzJI7c3aD3Hl1WFq7iwOyZV+YUq0Z+Gx1Wcs1LtfOKwt3/eBSddVFBQhe
tmtesOtC73LajKBQTeCpboxI1BHCcP0llzuuy/N29/bFjHzWax5uj/HbecNmP00Q
/2H0WVJWehwi770BR5aGLHQb4sC+RGWltD860e/Q3ypVGUnORveHGunIgyLvKql1
Y2FeS2aI1de3qFh4fM5AdvKHEjGqrqk6yV+rfAHcpaGgXvfrwDaSEfFPdzOT0e9H
wO2KWu6jZm6vEz6a6OORHhicrJEcYBEip6/rVd4SQSceFefigSxZu6wH0QRI1rOW
e8B0v9bFHBtDtzQUua+n0JkE8lTPUwvuWjl7cRo3FaERvUXgnhb/LrzBJe+y9zom
+QLrNo6iOHKZnuJ0Mdm+HZ6HYJt8DluRvV5WEqoP56/VeLRaZZu88BdtDlbV/R4C
dVYU90lXvIlIUHqxdsBCLWptwFqsgyzFv2WrAjGIKSUgSW4u5BGbcE0MXWqFATKg
V8l5AAsLrnbKNHOdb+DQuxzGbDsjT/AltkIUhZodHytdnYTevScr1xg4h09cOfW5
oS7zgFG+3SJ0A2nmvvD3skIp8Zei2V5xraDcYjO7q79BLmOq8Egrp6vHgrfQ+VDS
DE8lO4MnTGN7uUB5Ur4R8tctfUc72y1pgtHFKgdu6EoVv/rFyYjQdttqyTkP3K8p
5DxI5EIsRBrV1cT40nMGGJTpcTP2dD52lWj7I9yC/T/SrDAnXzjAXImYM4ksWR76
xU1QGw+sSKBXejdafD54OER4cjatTwROO24f/lhMKLYpAzahQ/nEUlTuVQguhO4s
lKE79OFYIPPx6nEroFF8XH1iKXmwHPLKM9vSV9oNump7ouZvVKNt5m5g59a+6Stj
Zt99ywnbB8ecX+C95mg5Au2xtgZAQjFFa3pgxm85bKw8vfN8+5LUGeBTDFIcPK6V
9GCv3EksdQM3OqTxN+lEMSxIZFwi2xdQ3UO3ngdaAQ44UNC845kJszAV75JmOiFD
tU8sx8cO2j9A+6GzNNVu0ACX8fRPhuF4SSwW2+k2rP+gUzylXZKv5U8ulNObr3ra
wQdsyodXx/vRotHa2q2JvsUOhx6fMxusI2B+OUauAHis8tJh9ESRLQ5djJuWoLGa
LPdYTEHz0DZ1Yc1732K2LG2+NbfbGl/AILw2Gc3+awkdw+Lresf/azUyDZ0T+yAK
G/zrXr7Dr4ESrSRwv+eCgmH0l544nNZzj5g9rCxyTMVFArFJ8n+uLuKSJGwP/FkA
GrtPX0bEnyMCkpSccRay4RojH8OHQ5lRyw3OJkML4xHQv9ShpMs35nfmWAQGirFh
/QPBHFBNdh1Q9+wLgUCTrrI6fiLxWgNjOhuRaPU5cYkAmd8EL/Xft51YYT8KnNfh
3bvLfB7WkR0HiDnmo9X/290TkfNkhfSfq/NqmkTzV1FsHLnxFtL8J1vjHuilvPId
jLiwlG/1GhZSzYpXcw/hICO8JGEn38wN/IjNfpt57Qb1abC2pb2Fy4jRmkv+pfDW
/v/OvVe7IEVByPUYSIOjpQxfJdODKRNoL50gizkADC4saiMRHRksP/16JYqOuywY
X3nAyTK7TbcrYxA5Lzqf9DRKyYWaSKZX+SRn96D4dNKAhp4Ua9V2h6N2mJfH2z/a
VoVDql4O9N93xMaPIQj5++esIjO4IhO8mbkHSczN2lM089Uj44sCYnsOhL7O6Cqs
fueRgac26gaDqijsiKv0b6Ip6X152LXnaU7m+3G5oNXKMGgymMPxo5sMvKs8BrV5
glaQjWNbine8MMDvvj1hrlKxTLH92JG9pd1hYSMI4WZ7dqeWrm6h/SfLKA1ghNYz
wSBII2n5N1yTM0mGnSJvyWgkTeS7qfO90D7ix75Ys0COgu9yKGKNql1RYmwl2xaa
NbB8ubFDj1o7Ygbumc8q41H+G8mahCC/uuc0sg8zQAHidh6VN4j5AsgXqNlOU70h
7PtFXy1L/IPCuznf9zqxMgHsmVlDj4+cCkidfy2/C1lRMYwGAgjOBt2b5oIbjk2K
NegLbtVvJBiCASpHhO5K86UrZsTwuqUgrjnRJOVSdJMoW/Owke6cXH08Ec2DXoT/
2Mk7bpCEjzLr4FgcYYk0vp07c6J6dAOOhUsTvmYhwSuqkY4/lDLPaItGOjm5OIUE
1vAW8XVE05Zfvgc6AYZMDC0wOHH4t+y2PIyI4qITRarmCdvEvfLgrhC3j9BRSgWx
Hkgk1M6PJnymxHl4qe9sSaJAxga+W9H4iAMQpbYhsTzzQ43n2BW7SHXJ4drfnIA5
BtomxzyBiJ3caKPMFsekMPfWll4Qi9wbiD4DrGLymsgIR2Ox+FI1O5WVolXi6IYT
dapWXPxZqimBd80U3Z03II8AsedTnNld1XPBGMC/4NlOOyLS4M7LtKCSDcJQzwYA
p+1qhuGeRZofRV45l4cyNj80s+7yVYP+rV+97GR7Fot8/V1PF3Z6v+vOKs7NIaas
cRAVO/EIzr5Y5af+VsFtObvNHvYG39BxTRwFNtz94y/Q03+7G13/0T0TM4UTKsgm
FfENHeUt+62LEJPgMxvo5+mPpWSznvZmB3HZRYwNnOckyus8xutDPWjfLzQuAmy1
qdZgKRkJAQfAo35Rou6kxtz+YRx/TLFUYjSjzN33xWL/oMNmZmKCu5JP+Ot3FUtc
OxeKSLMVK+Q5LqWytvjZHBtXsvHM8yskTl9AK2U/mh9L9b+/ldBMPX6pV9l+d9a4
pMjFtchoKEQiIkk8DiZoGF+IaWDTkqkazaYKGubpZK90nMYa3W5ECbWObZKqVawj
ZAaUlVk7r8lfT5IECawwEtyuxmp5mU8xOzdCeH8b+oHTPWQ2bnfEOJ0C7+jHGPe7
QP7PnpuWFwVzuSgSDmHTGdC/hLNavIe+1C6Cpuq/UpV92SNdfYRb10Af3slIbWpf
VU5M56FwPqFeexRHFWRBXZmFWSfRuFk6sHI7mmE2O7L8NAAMQgRNj14Gi4QQH7Xl
y4JwzpPiBHMacRMIMHrtRrMFWZ+aSkokKh4ac+UaIOYniwlSiM5njb2RfkDpJA4C
L0+2FiJ7XNjivJvyZ71J4veUtE7fme+IbWgEQzQyAEJfATE96/s6XCcFUpK3OFMg
CQlO1noBxFujTVIVP/qccY05yTEdXQ27haFrGw0sQ8t9xnZdrpWn2wJbzjVeUyE7
80oV2X4v/UbS0wHW3kd7FyYcTux+/lQk1J6aXmbFVWA6o+dUwkPxq4BqHb7LWyIy
FySzYsrG3VOenQRddQCOCMPjXQS2/7V+WEppYYbrwZ/BNuNimQaydvlWTEOjXGDh
BmO6cHWnx/rZhDP8Xs/EAH5LfLcSoiJiy+O/6Xm6tePeVgqgYscR+ic+S/ySJpel
ZlpIO2SIN1ga0Lyr91k+Mqb1lASnc7V4VxbfFKGyty8jRN9H5amsbUz4NeNA/dIe
uJDx8EEGk6QL9HgdoFfaqynAYrXpCRHt/W422lqe1PQZUNiZR/sOnwRoXCl0BtFx
1t+H96bcYSmZGP5GL40rpgGTDSr1FvxlvhI+lKHh9oenIDqqHRRHYLI3LwZqLVQG
rzTGq6FoXqSODpn3sz0EaW3Iwse6JvQAWlyNBQAXPKy8uQFv3fQae0avibi0QVCv
F4GKW/80yTFTubY+QFwynjZKu6BMgBY54rgtLM5Hqw3AtN29X8bx+EsKHr9pmzz2
o79130UnCcRrLJ57ZvgLygqSZYy6kCXtD0I3/gTW6o3VkhSci9KRMS+mEiyUvZ6Q
vui2owwbXEPf0yVY8B7hkn2m0r8w0nwXlkHhPOqWCv+iO9TJ6Szf7bugclV6sa7o
sgxTrUehfFJLITGAJUEV6nDxJ3xY+x9ZJH2rB6RK0522KX/lt6nHM7f1TvXvITRM
hStMF+P41BaylzQVf5gGkB73fi1/rAn/QpGMMdR1wIWDl0JrbJ8RURCvpaJ1TSw0
XF6CXbLDg6AoL5VpdZLS+q7DAoBC+C8MerC3MURsTTYU/4AxWND05/djsrBo6xnO
Qk89MOq4olHvaaCq+ekfb/0jIwbebSepNSjlxDc79leEI4pqTrSOqWw0pOzR5cGR
Y2kb9JJy/iJ+dOYQX9fDN4DRVoYFMdweaCUBK5eguZDEvo6xKnnQeYSUxbUKkZ6w
wvzpEL6hwzLmBQybbx086rox4rbqL/k+XtAwojkh/RhiIpwPpDrE/FbaV2/wlPRM
2/+ct3V+CU/67dVU+po3q7FGp/7BxH+8nzVM9FLzCo4Hi1+b3eKb99wEIG3jFK7g
n1dYDp9ROJv0k7xB+/mp0B58ImiI4miNeb7ojYstu2WUfvQZZ5vuFxCBobg9qbJH
FYBV98r9RxZdGD+vt4cGTg5CknSkeLlJ7KZOyj7a990UeQK0KnCntf8TuQm/NkH2
GE+VEYHx+usAcaSwaCXMIv7JOXnloa2JRN7GZzaHQYD/op0PMfx6DVMTx8fZRYLp
qQiCtdj474XI7O0GZBV8pK1ORATCKoZ/WcwaiQkfSxSCNe6Y8icOEE50rtQHLBkd
wOzgZwxq9xfo3H0qb6nlgiXKCCDh57AFfI/TE5McP+8SDA3GuPZVSLHLazm+yXb+
4A1b1wVK4XkCv+nVzIBIxdS1UDabCJJ2USttooqAp8UVljN6l/zx3k3hi1Eu34by
0um7WNiD93Bq6LYn3f6/bHrWq7/ENkCukn/6blZEX1j3BLxsoH1A6ul3peNjfMZx
IW4BgkO7e5eD2kyCY9NyUUfs/PNBRd+C+S1Hid8Uwro3TGs1CaTvwAZN0AEV0Xlv
UJz0zVILuMlLRXjRsNBwxxHiT2FpyLdp6pKnRdHaXU5kxpz3wsQUSDbEO7J0z3aG
n/HvcONRpK2aSOpGN9osBWsZOMkRRNgXeH6OSucIdFGQ8IKOHqyrGvb8u4YQisDu
wgZHxyXT+rNU+IfUA0ordSs/SyIqw/CC2rBbCgMEONk5BApKKurD8HUSlvk9s5/t
P8ceGkjFoj2dXla9Y3DiDiUQHWYQjHrencGyuNsBcaaWRn6JyxlKeX47Y+KKCEG9
C5k0f2Xpx+tNNm7DodiujYfhl2zUWd1vRD3I9JAjsUX+NyTFhVitUUDrTM2glYp9
9umPHYOv/MIPSEEzyRqnorp5P1rvQiL72KFrbU/EO/iadO1QGGOGHC/G7cGveL2T
sr+Kb0UWj2OsJsDC52Np6kgXRHtFvlG4TWdzTdLChbICwfsmHvv6Fp6eRsXxWamX
yAwGMoV4BCTLwL+JRrOrxOuEiC1RLqemSpep6W9trIQ2AsMFGusGHE1VGzrhXhzN
Zv1vnTeWbT2OdnYYIlGPvkSo1IeSoTjnBwBIiMOn4bFZ4MZfb+7dmD1CZzRS3Mez
pl6bOoLHjxnDzAivq4iDl5Q37rfLvoHtf3KjhfH92i8q6vTNtEVvUMOf27njaA4y
DP8Abm3AlFt40NPeSXeyqVGW3Iv+4THR/VBNipxevSt4D7o5fMUf5kdHDuEUHgZ8
AU5Moa3sl1At5y5Hh2vJAds8VFTfIgEaGw29+eaMjTwPM5pxpyDnIiKhnn5QYNfw
wOm6ckfxOAmxqK6/WWNIvxzYlsa6imy0vzPDS/58PNufiGBbJIRPhW1m+nuQlYRi
01NuXanQZpinJQQdEzVl4hGd7Ws+Cth1tlVE7lsXC9o9S/AJ8pWQ90Rn1qU7JmFR
DscvXVAQ0/7HarQJoduNkv7GobrffbzkXUlqDjcgeSKGyTIs2QWPZM2PEX/6Zl9o
SfTjd+rwW/DmZdLbcaI8dUrNkUSpKE3dc5cQqLrerpxB36+Aw+5DnYh1bO/2ZwP9
uImvj5fpbMflok7e5fRp7VFbIRxjZ4d9Fnyg5drW1NJihknq4gBd+MUDsPf+2bty
E0UnroUOz5S0i/MXgVT7PImvPwydTRPYvVkSElObf+mdk537UyyyklP43l6Ud0U2
Q5Lj/skGM81+ds5J17DXoXoiSyYQKiTgVrGeWdudQsydQ/rm11CzRTAQVf0ik1DB
fRpVjaBsPkwrCTd58Pk+fKQ2YJtlIWB8EAjX/IN12P9/Nd0Ya8Dxi0cO9Qttn9wA
tVhz2GxD6vftoAtrgSoutsOPCVwUAaPNO1YP6+SM2uZvjkSSj2CM2EMdttR9LfQe
to1iI4XPXnQxCSRRzVtG5tmBicY4UPcEyzyaCCTpCM/UJnyNpI4WTqvlkf8qCnF3
C2sA6ovrR1QV6odMf+CWtnb+VNL2m/QF+1GeNooDifOvssGm2Jfx+E6TTVFtKnL/
+ryMpvVYLbvOJ3GMnpfHpgVOyGH5Z4knTCj6EHaDTA5TDswWw9j9hMI2OuzoMDI6
OmXmofRP7R7h/GZdB5xPGMyqo6Eggdoie8WLR7aVkMlnaUxm7hrqfs2U1oHwJXIa
F1zal5RDoOh65K8UYVHH5rYOg4WgiMuk3gKJK3iyhIT3hRdEGnABrN9h8OlYRCOY
0BTjDUAjJGPFikftCAIkko38A96B5PDV+GDxBCVL9US5MqjDdVTcBRI7kbvU205U
e5X56qijqCcG/hvIWuW7Eb2choYH+XK9f1FlWT4DxAiVYeONG1PHvqkzZ6k4EsA2
3gPMhBhX7d9Qtk541e6sWW7dpRBDjvQ6/fET5mJUw3icKWcEdLGgzGS/SY6ZyzeO
MRdlGuNc6+tbCcWfze/bcuaDVBdqX6EyMdQq08wAg1Y3f7RnKdUiYx8fSZYxjFi+
4jlhm1IHTcfF2WZreuraH8oZqU8Lro01lnnT+HLqSu8x/4YSH0Trmr+hZa0ZuQNJ
RRzlS+eHYbwTvKsQtTCty1zE5CYZvxiidgF+Em3qKsco6mlI4XJqsNW2UFpJryNo
uIl7nB7vjNIWJh9p6xfOmZ5hUaRfAG1zUxvPEE6qbPrMYkGsebyGcwNaq3YG8gtp
LwPcaIIEsUezjh+30NyBbjz0ncgRCx+3K7nEnPk3QDnpvaE4b3ghuLZyoesGiZEO
9MW5RHheiXBW7F+9kVWZ6HzT9Sx1e7yu99z/N+3SNbYzJta1PIHu4cszilxso7qe
wpMrTEBBtgJOsJ81HJy6ig9JUguOZHUEKkU6rVCOuvFxvz0GNZng2+m+3qsNOLAX
tFGF/F4mS8fdgKGf1SfTjxHZ+eCGeC1DUegE5/XWQTyfI8vZXzv08yiF7UUuFEtZ
AlgK+NgZIUER4siy0HGlWVAFKyE88W/XA/aqVHANclcRc2E5+oS+fj4Np6EMATqY
1ldcLrZ6PJ+snVS+bgsdNQ8dIMN8TewR5bU6DZaF+GAVkXuSSdC0ZG9fLKTyDhS+
ShI6R4kzPy+GQzc4UUO8DfqF2gacBcJd+Iri+fNVvxUC4Db9YpK4pbioObv/040w
H4nPi9SUNYbTupP+thNS2wGQfuG49ICo8w31HVq+lx17fALBOGtzrRQaZodx5akt
4AKOnstKeZaf6pEYOXVz/oBe/iGnv3I9uDaTmlX495t6DB+4uFB6sRR9rM/bsljy
HuMqNoCIgC+VU5Y9PhtigGOlDMDQU82WFJ0zxBDQ6MiMS9m2u2P0837lwpZMgsaT
n924DhhrTaXIdbSWPWPn49rUdKyz4hKmxJTFqBDnrT8c5udtE7Yfehf7BIhWq24+
TZI/x8fT6tBTvBuiguu2s4WMtC8HSYuxWQsZ1RLnvbP5W5k0ZPLHd+DqTvws9jBJ
GI8LoUVoWNW4QgLe6+owSVJnCnp2so45zacQjMepX7SbjGFryBolChmsollxA48v
azIpwo4mqxWe+Bp/U8Yc+keumx6/NaR5XgcB9bhwDvi40+whQ6tUwWDtEOqK05D4
FH9Sihud3sZwVpbyCdJm+Eiwf92CflpLemd29uTsLQBHu+mRiyHVZkrgji/n8Pxt
B4kjTaOgnnZ0cf/q64XFTtBaoriJOVdirFgTpmcEamgkyTzreTaUn+jK5ou0xUMS
GjxDVR3eTHRWPfxRUat1Hu+uyie2f3dy3jeGILA33CmOMkUA5RTxidtSHhJds1nx
+otJDQQ+mXnDMlY8ZJa4IlTt4g8bNyaJ+K4fYl7kiMpUZJP1iaYP/Bf1iTDo2/DK
sKm/DpLaSZ6DNvWJ9dKcGB0Zqopf3NOKkOHpsUqMgiVHwyBWP27/mWq1tyGrxoTa
1IpCAr9p/5dDV41iEGuGz5mPaIWOWN77hH3Kuu43VyDXUEvpPRCNaspuAptX8I3P
IZHMPfEFC0E9pSEape5KZfCmqjoC6qLTG2xgoShpNXlEyz/3G53ZdcFakUdZ6wkX
bzwSzhSWVlrggxtcoCRt/Baajeq41wec5KAL/PDPrgD3M/hGUIyFnccTJr81SgYq
RhAhqp4Xp/vgPpdJJk1TRq9xT/q4ChLuULLho5SmCikVVGiinVh2KeMxk98FsBeR
aJkPQ47qcOmOpek/G9iz+FXMSSBIv3o6L8Rejb0+C8zmdyGGDhfAXQt2C//3li/e
fWRd9GgNL2QQcLj/MUnWnz5i1cROF3+3T4xsLLYpqCfhFUNKVbkdHebOHyZ1S6qA
nOHd4MVXmiob4luViALms7om8T7IOXuhRGZ+5LaOwM4SKWZkiqFQV7GCBHYrn1Cw
BuNgenDYZCS+mBD7g1PwVdabkoI9EakpmtsUz8yqUh+V0KnaxsHXWDZ3ynSul7pe
F4H3DuJxDhGtEA5JvjK1B6AdDphGxxxPOAz7VUtyo0IqWSyfUjAdODQunh/rtHzD
zgkS5yf0uBF0lbcWAVl1KECAl3BjfX2km3833sug4JhjUbgTYhwuYvd7vo8acQjg
065lLD3oZu4fNE/TusNZZfJIRc5gmCNm6leaSA0VuWBQc5N8fofQNmOcvbuQrdci
nWbcoW3LUZpue7bJbHN+cmisj2EVqxjmgFV48nGCEZYx5brPm1cVxhBE02twiRY5
ex/xBDjuZIOJdAElYRcf7TbGpJS68MycJxgQEB+sZLU2FzVUjd5tqdqviFmP1nBV
vpAXdmH5p6wzIIr0TRY+8Tke2piUhz/t5wDH8XebtAQOQCLeh4751EXSaQV8bq6e
vjoOTJTpk5xELxQQRnsj5uRyKriFzdKAFvcnSy8fJ0I2Dv5r4eWgb5hGNuk+nCOP
Pne2uaLymX005MDWyitxM6M5PhuJJX1HvX02HOYlUkgyGPKk+LJkpu43jwEBFRQQ
v7lUEXjFoqSSaZMD+hDdXqMZb29/JJcWktaGeMINR0WLBA2tZIMPvqfxhieQMdLl
GXKbxZigj8KV5T6KvXutxc4kN7R4hv1+jTx4N3eUulzfzgqegIqKcxSGoJD9GmI/
fE8j8WOBZygdfI7USZJ4qr9IC2/lMNszEVDkwJPEluTtuAYbQWPelSQAnycAQOdN
ZvSY9/fCJOSmF9OcLqzQQrm4cEt02/Io/BwDpV1u/Y8SoFePbQG5mnPs4eMLP5MR
Bt3OR9L3gcYQ8Qv96uLL27ezBmRSnsA1BpIgiA6OOlNs9ytqpPdov77EF+q64Kcy
g35QPhuYc3HA8wfKTcE9veWXzhgUNJu5spdXO2d/Gbs6grk3TW748UuFpVKb08QA
Rx9eeVA52jpxLJqHDv+Ief5yfbqAdJklnJFDzqXa51ZbmLAQsOkRCzgo5L3aPFb3
jCE7KTq4ZCrShGYJhkWT/rnyNqsRM/nmG9z6qQuY6U7JfsFvo4R00oTFIdzYMifP
+mlPBLkvMUx3BY4v633Msi3HzeAMO7Tg3PwVz/pvwTCbsOBkuFQ2nKJjR52ROs6v
ng7FI12h4gvs9V1O9mkjKTRqbrX0r2LGpNAs0h22qLLQmCzU0MLSOFcVF4jvwuAq
8OvKcdD0okXZHwfkt16x+evMWkYpQhYhXIY3gbj9R2cxnojO2cgVdtw6Uh46Kzuk
YFBh+5P/RB9WBnMAP0KoiqthdHCpw7VjVwxcueK1G3udvlE1/4YAosShtsm4O2tC
wpXZJiXamZ0iWwE9yWcY5m5nNErTo1nBeufCqz3fsQ/dTiwxiOVOS0kd/qqoC0ev
slxVu9ENGuwUv41EFz379EgIOvK8fWDCuJsfaqr6wNbXKiiGXrScfuEZ02HS5lC5
pG49iF+4L/39eoqvtJN3HoKYQjp3+qvE3je7p4I0mCXhnq/FqCTyBkJRQvavryX0
dGZuzY5yMl7k123LrutRzAJ7IiJcxyrd8tqV2bL2Xl2WyVioB2jrILgNidJcUAyZ
ZRgmsCQ2vkNiSi6b+Y3WbIhh+wJzyypjRxAByuNfs1CqIOtzArWX7rVhERegK52u
nC2eriygwQ0SwZDh0R2gO9NgRw5MJW/8gUERaCjJOOzXEDbbfSvURR/BCZV9cZJv
Lwtu3YCnGlTf1r+xW9ZBJIjdVSRGTALvehz9I9j98i3gPsI4QFQA5AKHDqpjgKle
m7DnQaGiREE/q+7sR6VZeBzVN9SXj7HFgcMAjtuou6m4w+60L95iCjEBBzWOoU8b
OCLIJTN/oj7dfX6a4AWVxBHkW9OX+Mugf2SwjfWE0CybsHzWnJCkq1/x64NeO/lE
2QyRg16dVuUFMO3sn7JWR1+nNq1bet6E5iqlbKmpG9g4YcvpdUUDh326iCrB71Jo
pkLh0vrxhIYikKSjVa9a4P7F6GS+y20wOtgPm3u56QKCExMjHRVjrQqxJwpD0RKY
Pp9Szy5aPPlncMybPGWx/5rClQSD8sXb6OVHD+m1Qf2tPodC7P+M7e5l6QK/WsGm
zqgob3bWDBrnt52nzmrIN/PHZlEbtkD4HBwFmHvQPJxadhClUcicua185+d8KYDr
p9kvzXTGcKVvE1aQUVKPTQ+n9qol9AkiTun4+62GIi+Z0Fz3MLG8l3opb329WjgH
BvrCAYyCDXhJJ8BNk75mO41D1deFQoAxlamU5MCd7wHGNJxqduUDvI0Mmd5OrP6Z
LGMe5XBx/0T+6GJHbaErjnJi6iuw2/1Rm5Us6nzf1+1RGLal6v4jFh2FSZcUuKJo
q06/75KQyybcN94FqrZ32pFnejJrJKr+9NGwtfjp85d7iRkWmiyzFSAmj1OPkRyt
/XS70CsAyA4QAwr7w38hPtL8L+rTGeNjsw1d3fp5LtxGIoi+TbutH3S8SKookQWM
KjmXYTvzlXwM+TmG6QrFwW6qg3BR++uLwbrxdG6IsTissxyPgith/b39spDyO6Q2
2NqvmqYCZAMcfxEWe3LsUhegvRqbTcwnWECmWduxo5SM7yOsmLXPzPkFxBvV1j9R
B9Vo6OVyldilmnP+UbbkSawioHE1uxU7LoepZfWl2qPmxzeQwlFV3LGpuam3ypV9
IQJw5yO5LAVLY32M412WGhBlEffBsvu5UukBZdt75Do2NXYL7Ghe7qCw3DlRDZbg
xhsqQIxhEcpsxHJ2zcn/RWKKXq5YfGp8h1KcNPHGyNZyra2cXCkdBgz07+5oUBEQ
Vg4BkAMLEyjzCGji5Laie7xhoKeLNZ+G4sH2pWxM66JO+oH7e0DiENMCcqsg9lgK
Dxm6CTt+IZ8kmAUBFys4Zb5xqch/xCQYy+DkpU8keog+2QiL/OY5IxZsJJTbtLZK
JVpnRbmZEnaMyWQo+fqJuLM2f0ufW1vR4cxWa45AxJ53C76JfGNkFxo+J62umcHA
B4pTAFBsWf75kyuwEyx38QgNzfZKz7PJbacAwHEJfga6esNKsBDjf9k0mnlViAQk
jx8vfPceX2e0hNfkzG+YgTv0zqOyx3qec86Mj3tHtozpddnKAiasWZduB9PTDPCq
AlYQwIK0XbBOj/pkLbqlg3mTsUty0aTxPjhTd4TR3+9CGQ79gfPAEESQu4E868Y0
xiUvk+JuJ+XQvA2QXxUsYrgi1W3ppHq6ICaw8hhMrzs4uu/ttUuI55gjn+UF0b6y
7VQ16JhxBYM+OaXwA4d72ZlvmI8iDtsaav7tAkAbd1/0bR289xJbj+1IYuonNIju
hKDxYQQOFj7f8Ggau9XITQapzFbvRtqzJ0WNSByx14ft8DFsrBudu6lUSj4xurro
8csMn1WLR2DMBrOZnC/47pMKuSWyjiSmglo4CJRW9WiCiZEGa7mHk8KiEToNiqkq
5UXQFNFqRZcU7a3Z83Wo3qvR0GooBy4ljzDMYLTetxJ/lf52k2R9K5gdyrtFFztF
T8SxcfxJAkn5UUSQqJYs1INyqd/L49TzFnhUef+AIOIawlWF8ou9tZh+cjTqUmXg
LWpKILNYgYC7wGu1R4VmJKZOoicUiQs0qJfo6ghH2kApGYz1GNTM8jLO90nSYI2q
oOBirS6vLU0OzYqzf6KDmfSwJX4gWB80LuVeAYpGfuGW4DEsjVmMSNBz54L6EkoH
CMMpcATjZeHlfjKYkgzubRUV1vUGqDmmGT3JOy4q+sHYhbwulHK6bd/PCQYGpC7S
h5IOF0gfrpcfxDplDulgQcT3x1S02bYyMneaSigUIBZm47Lh517TVd2mMlM5E/nF
4AZXmaEzpOPLM/yFXcde3VGHikJJef5coddAsyCfbsAU8sYcSGKSHDh4cFD6JXXh
1uEzWv8Tr0kHRx2xjcKfAo0rjE8LkZsskfpQLMU/OaXIzCw2e+WM2SAHwxkBkKIY
xBr+TmiSUsl+gTwIdZ9I35CLvR041ginMIOLKYpXICWQxoQz70lae/G7lX95En8p
y8u6Y+JDo4K7jWZr8GVBMyjtzAKyBF7zhmhY0b1JfK5MINsXrliD6tSq6jmG2M4C
UsRw+0z1AjsfIsHHWf73IxqxqkEMbK8knafSE1h5VoF/h3rpoySzfWEybrocm95Z
PqSA7rqhZiBWIoGhnASG4oD+KoVbRN50CZixiRexfa1anB414LBF0PxdtEPurpNa
GP1dq6aHuPsGNdcaXSEFxBcHcFVzx1TLGuQ4tkgz9e83QFGzKy2DH4Mty+Hya9h3
x9HfOq/f4sIoaCdqsbCp3HSvF0SbCbraixW+VSVm4n2NALOHx6qia3QcAlV8+y9T
zpQp0G6fshZX1pTK/hHrqsixGapno0NeuzEyaUagXiEXF8kQuGjQms1KmboI8eF3
Z8/YSwxLNT39aEn+JE9R9XCI3sJY6Mo7V+PFcy83wGq/oYPWH7nsPSBHzt2IYEL1
3SzrDS+EOQwE0St/S0s7pIG8lnA6Q2Fl/MGYmncJjlS7nu9zms1hVRRviSP1J1pA
yWswV1Rw5diEPEEalzBMGiDwsHW+VonEv88E1UPaBhl8cUU/552IdsBt+5gI9DoM
ZrZx/jopf3tnANOpbAvA4D2U9IVFfudUv0KMZbhHSOSH5mu2DUDgtR90B1x4eSLp
icwhjGTUK3iWNpU7lX3p9WS9m3o5Vr4xHtM09Qskk0xfic6tpOBETDh6tzEWdXjM
ehF6El8d/OOoV3CXaFMpiqpN7tiXkpcmx1Pcu+7GL8aksF1jffvWGO9rQsFJvzX6
yMEHnF8bZ5ilAenWPunLBJfcRM/jjmT1CRR9HB/ZKJvps7AJlDzwtQ+z/3glso0A
w70tFg0OE7BEB1dRaVgcEz8/aks/QJmnyvkHUoA4Lhkxz0mPaHflDwGVDqHNAabS
vVbZAr8l4tLSh76D2ifxO++GHeVWmwS2k0qmVCzwTUfx1rx0rI2oE37xRwF8XYGD
PcKsqj0vFLQKox6F3JxEkSHqAYr1TZXBwkrfSjfl/5nsnHjs9mJc8ikFnY4vA/iY
AkXU1X3CAP4UhIQFu14Ieo5tAbrzqBtXiXWrPidm1rgB/udYVTYmBa1z5+qONoqQ
XF6I1PigIwffeYjsXc0YRz3xZnmRhqvQx4qxpLnkIKe8yZg3clXv6vrATGD9wDf1
3ZAtlCwZYweW7iTxanODhpG25rzauBuIEGTDV0fG73Rnj5KoCg2/y+AuwDAalehl
EeuaKBxyupQLU3ZK/EPOdsRrrU4xu1nZPTHwVogGKP2t+Gw8vDC5unhNZiFKhXoo
+sAbgECFMCtICBjnlwivYTDGlnDP3yeIyRgGDYLYmRzFS+4Non28bMNoXOnYmzlE
6nBpL8NNRkU2itW2BwzgEF5Glj4nae4KQ4/YMKoPmRVWHTyf+OwCGYoonWYUorVa
FeXV724XhroiJ+GK8UIZC3mm77g34YgOAYJF9fV1RN8KCsX5PbwZuFCQr0kugeWY
MBuAxVV4zZSgVAWdaaqIjfNODWsxxIDGz2H90QCiQh4VOeDpV3E30aFkqsf81VOT
8k3tYrWTI41HGxiRodC+pv2H6mGScx/bBITKSwHwIL1SUbaH7G3rT9ez/QkiII62
oe/KANSU0BafRsX5k94faqPXO10zH1huJ8sKcnWc46bKSjMf7Ygkn6nzofvSR2Up
wSBQo/qQa6agvgsRDgQ62i6g+URtwolshevqmtCSbwYTNr2RG5Q94B8yOyByi1je
R1Nq+zMQ/o3GRjG89mZW4Izz1fAWqjsgcYeaocDa2jJydEeG0QpA4Q4yR+blfxan
WwVp+T9er5Bf9vg0v2YpxEIadWkoje6HUyx4Z0w7LNh+tRbbOPU0aHvkiNbWI5Qf
eCngz2BlOPnR5csmnXnP1a52wokzckZQdECJYhNWWtVIyv39n5h+JxRo90EPinZr
t5HfCc4xl1zA4jP1wJgTmmJvjQse7d5HLVUI+1J18vq6F7gkhOzcXfKMaSzSAub7
K1zlqIo5sVypYekFsFtLA1ZJd6C8FtjoDs0e7v2gAM/THYpKgMKIidlozJTIq5n/
YdkS3RRShXgFl4v8UR73KuEC1Fe8b17F17h+9C9gRi/pfi34rtxxHlNB9uN89Ajc
e54LzrjhCrz4vy7tcgaEbUYtU/ghsLBPfe3P2voY1rpL49Iv+t8UCR7HewOC9oEO
2n2P363dOjWauM337T0APWQELJ0XIqXgngDjd9sgWhWQGqiAMUOfFbbpojZ19j6m
Gwd46O1oyBIaEdZQh9sp+nrF2Z6hSHBUgMU/C+pkK3fHwnsNPdvopBp7Jh1cpTvT
jITbD34Qm6blggWHw7/Zmjl1ILSxazHUxdMnTSo9VqxMHSuGrB6796q5n/5UlUJQ
a6EKE1K7puDMmqnqYBHa71OuB7EGnCu9UgpzzmABOyxiTHi8mqZ4oWfywZuDvV6J
p9D6y5NxVI1QyOg2CHu0RGc8Wc5fYdiqSlSJpfeeL1Cqt1yMRpYARcS9v2HRKSZw
dowaWQGo3yw6xps0jnc+xo0/u+BuqVrAH20ReGw0eyLqyeJ8+siIClz9UhVxzpE9
HalTBvRPRVc/RymAew4pEr4PgrFpc8DjKKJdYoGj+Lhn8AcxdMqExhdBTkVcJc3B
3mwoDx7Gl/STTp5X1++rr5knNLGvunRBAkDwgfan6N+NyrLQYL3hYGrM+GH1ubM9
NqgoibtL2bcsR/uRG9y3pquc5jXFiY3MG18reWR2mOr9MkLR1pQEmIT9NigcsYwN
oLU1Gdq4r61PBhCqClCq3HetjS11bvfwVaKDpxXG3dw3kOg5nsz/qoYzJZCWhm+P
qLauvtpmcxJY4+8ruIYWBkP/yWdrH1GU2XzQWRfUtSxpErXa7zll/RU0qMAhHPBO
CXevz40TjBfTnP4QpvObFiuNbwRmkI55eDcjrT077+ZQL8c8ws0Il6vYDIGrrOIO
HKUYbrxUroljGCg0C+Bd6ikgCCScXkdTQvrNkuc7ltP8E0qdCWnBRiEjMWVInZ/D
+tQNDkwY0YYjy+qy0qahH3bqZyVFBT2m/VC9hwInFhNUE9QQ/asJucpNrz8GNYmh
vQZydfCb689YpUt42/z0Er5wB6g5mx+FtK6qdQLrGxbzA0fiXSHxZc17woL03HZK
10LBNYWgTwdkmYtRH0yx2lIUTpPZh5nUK0cBXxwDgkFOyIAOHbuM7TazD5FNHFbt
GVktZXJmZLhtkI3sX0Fq1sJeDzewhCcoGBPzj59XpwZUeUXt7tEkG6daoj1eGFRu
ek1Eh48IqiuWV8Gvmsc2aGk9OgZYqSrhWuKjwSmWOjIDTb5Q7kU9ly0wxfEWn0TM
3g9Gi8veTzqoaJAKd/XX09bi1FlhzXgFZAMux3qVh7IbXy2Bqpw5vkgWRGCU2b9q
gqLOQOEPEJobNZY4kCvvjxehyfwNVJXn2eGTmAbgdRaE64UXe3/5cEQ9qhZtT78i
YQ+V82t5ErxecxWXR5hAvk2ix9B2R8G34mGLGdr4HoDD01ANrWueopYlPdjXAFO4
YZPt+cy34/s4IEqPEqrWlmZP+WZ0G1q3gx0npedkEwKvRqrskjLrpEvaGgq8Akw4
rxmNN5VNo8r2vYbrAuwfoyaor26lsMX2OIWO7nxygXnFURNCt6wuIjQlTaqNmeVD
EmvuZ/AxhpRXNGcfywXscJrDY+1Khygi0My1FtJxif6RHZiXTMlZH5YU9ZEuviPJ
5exHsc4GgsMjWW6ZNO1m6TceCQuNX9LTm8Jbf6l+OjGw9/FN8F57a6OdFBUAAXR8
31PqAVLxBz8Oc20WNKh9d2gBdwsGFr+IGOVBNP110DImriIukuT9pF5rIgx2j/kk
b/txHbIKJESKx1JN5bvDUQfmcL38O/D4NRPQWkCqMPPJErKy+32e+aSwD0Wxl+SW
zYx31xA20sSf1da218WWNCmwbKv1xaDWvxykWLxLKqyHsM/rUXO8212O4HyiU5rI
NIaKdRb6VZqxQeSaGYTRhvZCxHodhlP4IWEAFBU38N4HudjM5hK9xRIdWFZ069u2
B+wmPycJ8a1OfTNAocTUVQ6FPSUeVCssjs6HsAKkAsVLSqWImOIHBdCdDcIIuJ8b
SMgdFnWSWbAtQsdkDZDPlBVXjdOF1ODcS1Qyfi5I8vsF8/iYpjcDD4oAG9sa9G3U
+45OCic6DC6D2ZEg/RRBj+WI86rIEHV154RqeJGSAmMEF+jr4Jm1RdkGnWkiSg9S
sEIWM97DjlpXfSLR3BPpyaViHqUiSWz3PdDTWDo5ebxy3GE02KxWKtoPftaso4EJ
zeEQi89pHjKE3siFDvqScJcrrhSXFq4sCgL8wFljrLAXxXFBYSNru7Tmvke4klEN
Z0xbvPGaFps6O0VAI6Rzc9jpU0WW4tukDeYLNJVeweB3pE0xJSU4UcjJpKdtytrD
DwwY0z20s+JFMUNw4eeJhUcwtENjzI/W2k3LY4MLKjh9ZgcVTA+VQU8c3JuC3RLe
vujsRdxjf894UPtz2bqI6KzVtDeHnrRetc9wx7aiFQHGOu5nH29C/fnMXhAvi914
NoZiZzQ/3Y6kKj01FU5I4kFfB+RIXziEeZ/Mdx62jwsPb4qadUnaIZQtUBN15uqp
rNnCBFAFQEYIYw9uEMcZ4wLZidDdfR6u7mvnj50FtUfKemtBw/oifxR0CNjw+tKE
N+vMWvD+B3x/ba7/8mrXcyiKNAShT/5tFrEVpbwuGk0qM2k62DvgjL1UbEGVKSRw
M8wJq2stnYwY9490MZFLQVVeLqt9nR1GZZ2PMrLFI35eFNMaLs8IbX3pfTgd4GHL
8eK4Frl3xT5Zmz5KanJHfxtKpznhcxcb/TzOguS1h49XxIHaO66xR5zg3tOKbbxv
3I7YPMSzgSpQfEZu6m3KvXbOuf1qxd0M2pbZGG03idMrKoQhXw8fm2U4edmCY38X
2cw3hdR0qKgGeCBuZUUXuDJ6iiw5J8oowzV5LLCPxbdxW8AA3KF2/26GnMmpz19p
cl6f/dY7c7wd067BKREYnVLCGBpP2lhhg1Qi13iZP0ZZY15UsWmI2sqwFskn72cS
WCwWe9ygINQdDl4Mu5pKHSSntjtxXeS9pYtqKNnibcUek1DzIBcK+AQWeSDi+wbe
e8o1YXbHAB5+h/fp5u4xHYmajGtdIzu1AKSPPSkhbZIhnKz01GEC+hGZcrkxrghW
pm58sRq0OddIweUyxdab2OADyMuP6T+WXCWdazqWjqdSL+J7HTYMfoy+hO8gJiBm
MwJPiDHSk6ClaghRaXpf9Iva1G5H715KBSZbNiyTkkzEeoY2LAoVS4vivfScvD8Z
INsedOimr/L1lo2QQ3k51bSxc0gC7rCfod+U0tPZKIZ26bZj3XiputQBrXwFLF+B
e5GnlBqNW0p3Bmq3Ox2LEqsCcqMOxs4C3dbdXycMPTnrvx0nAi6zAVDKNKgrkcRh
ITjrP/duvOEobsxJ9ToPgtTpAd5T/30eUWBtxugX6/LILaZNMvRiJ+tleBiVnSW5
lKbnP6nDOJQgJ0MNhevLjAqnYwRiB/ZN6WbWrTBghYQJXYMS+o55GH4pIyiLEJT/
O7HVVqTamxyslPbnhGZKga8neTvB/HLGrCM5XrSEh4pVsHA/FEvoVZfChjldMMaQ
CeI48nwdzjqL/AYj1vPSeqsExpDQFEff915u3IKAw4oCMBIi60v6sfaQe5XFl+Bt
sYfCcUJ2sBH4HrdJ/i/y/tNVg8awzYb8EWL3V4f+MoPTpGNJnQLUADHZ18gw6THY
EcuqutQBqvFXT5nHCPpPKyNgVxNmv0ZcxHuzR2/K9NP+HQ2twlQDew6AWg27ONCF
ckTa3gBKKXH4Xx2udc/PW6mM81pYpAio2HXJzSju+VT/bTwXpOtq7Ap8lQcozJ3L
gRBWZnp6ofNjhMjdGpQlRZOP8dGDlNEgyNxn+ZnnSJ6Ja3uggSCj40GrgmHR8C8p
kDyEeBBhnK9hBUdBmqlkKBiE+A/DCZSPRr5fuT4qOkHXsEVwKv9xSnlkqdFD94Pd
rJ5fa3IsauVwg/DiGuPuYDApIPJrzO2QT8SZeXs6TpCwwBLzscF251Chcey7BkxR
QyQfA9444QMx3VTT6+DZ6fRk1XhhW/62UW4t9Poz3eR1FFn6WleOy86p2NPRCXd/
jS9tZn0ieW9MnvIYu6g3ygCRzPN7/Qhm6vrfjSGCjRnXyezjUQRZj9LoitkSsIRQ
HPrt62jGw54GVN6xgPU+xjs3TONTfLita5M+nyAyrLCYYIWX9b2Ab6zWmlxQfqRq
KfM5aPI5snVpVBv9Q3xHfoz9bQwq21SXECMagtUOsh68gflGmND9Jf+kXHA2Wf6f
vmCGkHNxc96Cm7sNvvuBxZNByv9RncZN/hFV7jEpQdrfTs86Wayec3ucwiObvrZP
9ig0Bbd36jotHxEgN0OwUloAWexQHk819E9aca/f58/9k/C90Uvec1NITytwAX1e
NLGINn+lAGUZ5k5eZ8mg4d7fYSDER+15Ckq/5qqR30GGFRBwXSFXL6xycFFU3s+7
Ae7F/92UwDgjbaDjg+hxmBncaFH3D3e7LVGHfm8j8ls8/Lgdo6zLoXpKhkKHEYPc
kvUfuQaBTYQIr8EV0uEzYdWwE2lsBQ2kMZiWhrhlEos5Q82M4KY7dW6PAFK5xvyk
PJTr/6UsvQ3aZP0Dz8AIpWDPAG5TFDJyz86Hyx4k1IFiqvh0fiKbPhXwPezlDDTo
oESZ7luVhB8BbAbxwGBvNrenX29MlKGXgltckYnwV8/w1z+yMDbj0WEm6ao3tQaE
xMwcNHmE+G36haBRvTxyy7Rd8wl5FczWYKONV4rvNlf54yCkhNF75IGOWPjJh2TU
ZfAq4Pu4U/NPq9BHINfXAgrDnTI9vT44kPF1aKDiSuhwSIOOEhVGYibBokTkz82w
fQkWGgxRb5hkfWN+aK383F2RjJLg8rVSmeV7sj39+y/prFNmEblkEVdAIvlEZTyi
fRbg97dcvqkg/ypAZ4EoF8zvw1tQ9AYuJqF36zhwqgoaWDNoYu7KFeKhqQsutHAp
xHZrQpft8dcLd2AUJ7inNNNsCasBf55rY4aMnQzo52kO0EJGaZToONuswwsNRyPC
U8G0m3mWqpnSibfqaDSx2tGfaVP82HNXuAoLuB9ZAEY11hBfd2NeJDLOn1mKG6cq
De7uDtHJNimFeDp0Gx3DuYiDZjThAmuReuz7ynuyNASLWPGL0q9VLaaqMFtfifgi
HJIXeHayBxV+y1QTcmSf/xe4xPC9oqCZf6yvU2WeeCvNlN9Pryu5EF9eeVsDvlvI
rWgdvjttDMi8RCJu5vW674n1cg+GY0XYdR9f/XBU3noeh3nISxaTwxTZ3jJccmu4
hPnhqI+b0vqfH5hZdNI16hKKZyR/qA0NncfN6LWxaGBW56wmI4FFE+NImGfQV3Qu
MQnVpVnLszxDep2uQdrIyznJYLgjQhPtrHnGTC3SruG2so4oEbIuO8k264FFB+xm
scNZ6+IfI+JS2cBwIQtcr7Ok/mCBUUrHV8+kr25fE3dEQUgelPbcWBEotwxCBMkc
x6ffN8B/W2h60//W6mI0P/OBLyAXvUEuF89vw2H+93FcGLY7jahJ6nO6t+a6BzFH
tPvHToWcRG0yi+a4tNdlK5dZw3ASM0I5Xm5P6Y0JDtU1lgZ2+B/yV0bpJGvSfhvN
EHcJfUNzRc663VOdZjtUxA7lb4SDdTaTtYM+2uEvBhsHwkryYq8nZFNLPMmfidZh
33vHHc04qQz+8UR5Qg4Bhva5UM9qyvYdCA4enWKreFOfjp6ApLy1PWgPYP62KDJ+
7ShSqNLROaEOPdRWKe0+8yOdZqz5NElK3tTREbV2IbJ9gK1pI6YbhbTDxxiUux+1
6NGhF+BEyysEGFQbg5boTUsu6MObLIYTzrCVlmFXRvtRgUC/NsAV1V3cyZ8gcpGJ
23M9jfaes+J6t67hWCK43BidQqKFaqDE7zuqpYLdGEiLmzZt54i7lATAeBHB3Tll
SwZGThtdy8kRNi/jowmdKzli6jdyPh5d6kITBXolL5XOtTtFi30KIPw6iUphUxWx
4bofl8zMVo+2gOfovCCrKB3C4Md1O48r5VnrSCU/0OBi0dyw/5oKs/enXGV13zjJ
reEknVL24YOgpf4ye+7bRXLX4zDypAPNi3ityTey9K0znP3oAhliTvHi6nFKyUrz
ibPv7ujwolefopMYvt8tvSy+0keX+r6POe7ATKbrKl8uWPiek+lJ36fZxnR88pf1
ufMqcSwWqkJJMF8Tl9eqZPxcoWGb8Sze1OmCOhqisvrTymd51V7SeyluTPJRifI7
9U4xNg3VBC6RY2TgaD9ZPSqb9RN67tvQ9MqN11Pjwr5uliFwMBsaY6F3pLixzk71
zM+qFkpt5O2zbhSwH/lk5ka1ZlfJrwaUpYms3IGd+qSemRsfhOLdMlR7fqJs/HXx
l/4sSeXOtYppJ+nhf3oKJzTjcupC5cOs3uVPp2Rlaz5H6kF0z6s/+H+NJk2woRTh
XHt2o3pH7b3wer4xYUEDVxn9BfSBXrOYFLwwXLJ+e2yViJLwP600xz8xVtgI5LuK
ibOTgykk4kkXcNgMQ9tvxhfWFFXd9mEsKQEe65Ni3e36x/RTgWxEwQY5/tRDUz8V
MRjyPJxUJ47TtrHAAm8X2fJGxDYbs765wxPnmGEpwflSce0ZuIa0SpJk58rufP3X
nKVCDtLKwjf5fwfZXqFrBlDPoAPuT+kQA1mEDk1Vz7JwSKTl70jl9rn0wHklLfNC
LbSWxZygL6+MyaUraLifqfcCmoXWSZbxZi0kt1rVMBbTRcmWUBNhY9iYFV6ywXMp
c2OMdEg64iad4MhUO9CjK+tIVc2b6sqVOcp3K0oUmaNrokMe67lpRQLxBN1vhzUl
/5Kl9uziVqxKvWWvCtlgBtRZarajUMZdNChK4R6G1bddsQwljXY3jCuCbBsvTNYP
wMUh3ZS9Rd6P8j6dB3zD3BlaGs09T3sjj1bTRW45OlE/gCBXcqqQ1sxQXaRU6aGj
UM1iM4W5Cnduzb9cLKDWMqxfYMe1CzjZeo98bGPQ55mA8Ut58oUkFf0t8JOCtJCw
7OGkFZvVDw1ViPJWF1DZk0gd9RKAOwY1eI7Rq6gvIcwHsQ/G1SlSSL+QQjJUuy9G
P7c7vd/LK+QvYeKCYF+eo066cjhSv9GCy+XMqo+mfhmhwP58BmUnUqRsmYs0isto
hshs4QrI9HxxzNUBO3Bi8irClaYUXplTATUQD4BpyiswFQ5ak14jytfMZkkAoRZH
hgfHryajsm+ZTg3417yaDYofFZXbwyiMqIbuarEjEhxQXFOwdhEXg47nc8CdZKzV
muknk4txThN3EfE+Wm/ybroyKxRW/g5K7vwatMlnUNcF3NmPJV3aYn5XZnEcVvCf
0INB/SUS0MRETe9I++YPsGCNx22iozHVUphcxHkd82DhxBol/xuzsrdx1BFLJPPd
1s34o6wt24JjNMm8NJcUnHmVG0GgB7wgSkaXA3ZAkFvae1DkO1hDSKI5jlre6Q3N
Or72JJYW9mHUiaWm2teraP+W84crufXlEhMonYGAdu/WFnsOo6LwtA5w0/hMYZe4
u2AFV3kd/+37k95TiUiTyKKnR96W/8LwVedBZJpioSxcZNF9oyBw53vQyy02uzee
NweXdYD/pV/f3UxeSUXxyxpJw7nT8rMlSpz59H+Mc0nUe5EjN8O6dG832BxFdOHq
7jchO5sjhvOGJYtPXDfXPSGfZlpp61okyQ/YtfZJwFrCMbYXX0Klv1bC20lfSqxJ
tEzOwMTDSzc+8E9yob+Uie6NxxtF3CZqoawwq6ZojsWgaM1859owHmlFXis15Ngf
VuFJoUf7U9lvdL8JUUkQMAAXNnxrqbsdERRup0syjkrXCuG5InQc37Ml+5kbsXFN
GPNHkhcysd+wRJTDM1o2zRv0MxiP3Iz9UZg+NMzggcMFMG52+v4BQJPHwxeizgnt
JtoOtzEnxWK84DbkV1T+QPWel45pYrMLwMCIraVs+g54rxYYgJlu6PEajwLzXrIi
kjdQ7THaeDm7tfOVvbT/mhrI3MzYrVLRXyG3wfRKLbBwux66JbRqnnBXPEfX1CQp
zImVXrfj40G+HH78iDOhXHeH6bqeNwHdx3M59H5jqHl3KJ1W4DgQu3nyFvWerC/o
bl3DgJ5fuqw3vNMbTdPS6Vub+AiIaEWU6PKGJ/hBAYry7u9OTPD/AOXCVJkbXeRC
2C9sC1MMIKaHNtcDHIz+lLkS1n/+q9+IvN6LFaAuD9gXLNe1R32qZVKKA5/3yYsP
Biqwex6SYkx355b0fOUFOP4rcvjhzY2DQH8HPmgzlVAld4W01cYdrefMfT9nrBPO
KOVCtCFfMyVZLyuzHHx5hKyR6kmG1q0s9UPsSm07h8szTtFZ6eORW3RIx+3DwwUI
KM2lPpEqIykl1gPBR2YYH2getxdCT/c6576hAlaKLdro6XML8jKWO+uk47u5kmm7
WWKlO8SrazlRbAPCMNnNdB2cLI/IMCF3JvoKoq1aQjdRSsM2PTfHA8Ke4h7j3OCN
VrDhKuMa4t2nqAo+AL7JQevc0ohHH7O4qu5+CenO//2ZWOCCgSZRYmWF2V4EO7T9
NIh6b4UrMTASOdVKZ/0YoAvN0QyTZfZY+QP7iAPmep+exxmpMZMiKBnKKIWmeMz9
xTrijnxA9T0Xu/z16TwaLy5MGWQ2Z7miYzxpWpBau/5ZsE6fvqmSG81jyeXn0Q+J
chIlNuRD9CbiU0imN9fSaUGF+sqMp9ObfJ1fmkef4CPLnIRqmOa4gs7e3/VDmNkX
pJcmiRo4uHqXeoJGEXkMh1GZfPt8TPV5M760Ojv9YXqU6VkKHjyo9raOqrTfL1iK
BoZSvQT6ehmvv2WmAfXErn54fKiKeI8Tgn78LBtDCKb6OsT8x/gAD4UKNaxPsuJw
+cZkZmOcEHrjyKbZFqhNrTsZHZiFgkM5NoWEwPndPRu0osVVKCH51GCaBPOC+iGW
yBrH+k0yW/hNgD4+3z9igegiT/TDhNTjWdEwyn8ANuph7snGUd9lbXXEqHmEK83U
eNZu2GCrcMDUOjKSlcB+sxBRz1goYqrY2taBhbHuF+LxXHiX0lZDxypUZ4VnhfKb
Rf2DV3IA/4z2HjcuTORzc9xEtVcPIZqD6B4bAv0kXRUdKp2JS2m0QKXg2mWzV/wx
ELgfipKLDKswYMT1orCiQIk2PySTcI29k44cSkJyWoXInWuKF6MhDv9ccQPL4tZZ
89CsTRUlO8HysFYnCMlQg0pq9VJlibUufZsrAd7OJ7aMBliqMQFSs+yHQlODG4a0
AXmEmfKleJpUIwI1C5Jsvlrw/LI7jgjEHGl072Cwv1JsDFsd8py2kLPp2I+fJBC+
iCOFCknbURKHAXn1HMSbadzVPfQuMi4egw/Kby2IgNE7PTae9XaBYzqWVC3fPqCu
fBFsmLlScK7dsVk/5On38OTvV8enFkJfYDCNdndymt8gG9gaGEtAkCga7RdJ5Twb
L47stWmnYlpq8IfABNVOd9N8hHsizU7JhJYGAXgL2ayEDEl4UhKYeLRgKEK6Eeva
M1hyQJ1hD+kAVB0PnnHNbYIsSOH3pPKe93v20o25sLbtHxQ7HB+14p6mZPSMvARc
iHGvsr4FcXCoKKW0DgizvUNgjpw9mi893m8uDhdAgVXhjK3BjyUShIArIDsFCrGQ
uY0a3e+DiPky72+FBgoZXbsfKgoOC4DAwNNysZl2C+L5b77symOKhkpFlkq5Fb6Y
9X+pRUJ5E3Po1Xqb5e/r+0MzJqLU4WdjkgNEGfvikNYw5KzT86R/aX5fNCBC8yrv
Ztrb7uXaNg6vdrIzu+Ih6p3h3GQZl1gNzbKSNIFDk5Ui8PPTGtZP+RoDO96sBQaH
0YjqCKr5c8DYhkNkYIkjKCzSnFVvPB8Ng/wGxhg4S8L+yNtdhMydk9KTPHOqvgvh
eAt10vXfWEjLHuVACj+L0IorRnN9SEmvtLg3pooAxUNrZuSSt1emem0OHS705WTd
Z/Zb4zVfnUxIQGpH0gcpJJkEq6CovPpk5/895nBajEz/sm2U3A8amrJlbTGq3ju8
ahCH8dre23aNkqTzo19uUxUNjUHgKvdDP+/7gKouKMhQjzjtq0Gd+thts5pytwbu
v3HrYRt/puRWBtDkKu2VOwJz626llFmrAt8anvn3XrEXgz3R/a3vw1z38sAphc1y
UphZbIOg89+u3Eg4kyRgb+ZxpuQfA9yT0L63xicmvuAjwLcGUr3kynb5Awy0exMm
BFSc9sDoRbk6iUgaGRGqCylRbaICeviPa00OCi+gFE0Wd/Mre4oeGzkXFMr0mxLB
k5mH46TufM1NOcBGrgGADCAoaTiJRxkEGw8sHG/bRBvLqwtzVhdV2MiCRVb+VOj8
+taMSv9+OBD+67ajmOEej9RcwE2tN2Jipqe6+XbfjzXvFHHc/joxNsRChyQLhUzP
d1kUgFmqma38ZbCP8FGLQQkwlcIWS5PkvGQR1RMsPuoPyBrQ7DQeGpk+h35JYS9e
7XiBW/JjbR4gO6kmPLGz6jmTR571/6d42UueBmvUYlT5OHuGGE+rcXIQmYJsBGQj
IEvCPjLVh+25ic79eamHo7DKeDvstyus8T+MHUW17U1HqmimF/E7xXK8pTQiABD0
+lCrhrSIPaX93HhFwfzttvdzaBAV8Xv5rPvMTRbFNZGaCR1Oe8vn9Zl2+zrXfulK
Py+qAr0eTq+cG5UMgjyFYbkkwBdbsRuQxkzdZRVWOcmUayTBz9tenKrz9hJcht8/
3F3RLPDYF3UJ+yTkTy0Q/4f0kjZOA10UKhms/qqTNyu14Cj9zvyQkdBMKYYj/ObJ
D2owSmhAXXlRjNNMhQDF463+HPO8FtVWXEOV/zXTp+R+mxA1vHhcz1w/Jpsk4tTm
mOBtqObU/4QWmpfLSFm8P1zXwU+b+tcl+vDA70qrkuRoJWk3iWfaZ5Ug+lX1Z0R0
tMPjoND/coFAAL6FyagjHZJZb91A4h4mW3aXyZXAkx0HLG1HXQ8Pl07IXVdur5i+
CWwgWQNCOpg4EwDB0xIpL7/cLgpBzc1CteGvrPmYYxjnTDyndfOtEWAF4LCO/hup
TJ3ttztu+izPCseYVFRvXzVpXsgiaUe+YcAeaqsF+uRTpyk/ZlviiOATVoLFGlbS
HIFQAhdJ6zJVOjpXzDZt0/hirTp7jOo2zD3SzGzxLYZMJ+U6gCSgFbBeXXJdkIT8
kr/leVOBqMMD0d3VBL9vAgjF5No+rSEgZdXFI/bvA7z1UeXf3wD6y6nlBhVNisiJ
qmj63BLVwE2h0vcMRbDOGjb7TKUExPiGYAs5ZKQT7zDgBA9ViyA1lvZkBFXobM5X
n0ByKHtWN3zuMSwWX9wtfPbTRjIRwgL/rGuWwfSKr8a+q3kjpyz8TCS8dfK76Tju
AoNLtCct/0rqqOnNvuqFfcvLRjExBZn29A2Avuhc/ETkkIG05xN/YYVZCst4x/wk
h/2m0ipF8PxYgx0ML54Zz0chwxxiTmWVIGv/rSI8xB4CQoIqMDh6pl0Minn+9bnq
f6OfdUnyLHxBsF58S0RTUPkeJBRQIhGAqJJwkooHWyu6nnuhWkP13bMV8ujAnKBO
Vvuh5T7ejL2Sne2tEFVa5IaxS6tVVwvgssjHFaqozZbDNdUDPjNusnttdik1bL78
B7yGofhZY+VotXl29stQLmJAQOVJ30lL44brMKlmtOuAtVvSDtif7UHCEkGrUO6q
t2fvcVEduLd5HiOYg4H/Edev9pMBSJfXprVKJWMRtxNp2vbzRG7OJISgMZxC3KJj
4oGwt5RehpvSwg4bdnGB40B5GmgaRiB4+fiSguLM4reoFhEL1aiXwUCwL4I0UEdf
0kubnogxXsJ9Fi0tHm7hLc/97aec2D9ItSCzBTk8AsWKKnuRJdfVxazBybFd+zcH
lb6na0xu6u2/92sCgf5IKBOyhGgxD3J/NcmWmia0utcrpDtEySECF/ayR58XD72L
09M5beOxbdJKbliKD/sq4ZEOwOGX6wiBsCpqG7hxYsn2pPOtu9k64Yq/HrpRLjg6
sG6ES7P1S0iFk5meVYP63EtHIsiEx7muUe8dWYhWktsV1pertRhFkpSDx9jl/QfG
JVV++Vyy2huI/iGdGCsccyj+HdPVlKM7L9KBwg8tWJJHCmQpkQwjKBIBtNr+Gkzz
tZL9Ntc/KWTPCVftz+bVGJFst5i7z7ienZjrP57DzfMP/a6mMOL37QIE6NDtzUQL
ox87LFRghFiAf2VdmE2+ZOr5Di0rAWaTSss+oFk/G6k/cMiZIFT9LBqZQ2NxykHT
b2xi5a6SrqHKz3Q3i+652WeH1FKB6uditquCM5rnsJ0CQxgR8dV/lgTFT5PxiwlF
UuVHi1oceHCUzAU80/fgVMxikT7cJ+yBFk78VS5IFGe/LcptuXGRCYIVRZyDK1O9
JACPp6HKYOebGzVb8A5kney0uWsxeY/JZzvClh8orq3sqaAKON5vS9hjF5XYxE3D
BAABNlp3L2lRx9SVdLWFw5bKMD7qLlW6MbaTlAvNu1VIuGLQ3T7De6m7Aabxpd2m
o+DxKbqjCYPWKQiFqF32tVWslvTpG7SATZOW0n2AhhYYI0+6gdA4/PDzuA4fIs8Z
fqSFUi+lX5Kq8q+K531JlNrds7UGDZoLMR2GcNnusccVMYYxOBXiBb0HnKbRkJMz
U70qm/3zAiHzxZJK8uIzrBS/9KwzI2c9fLZ+jt7XzGL5nDcrlcDjecSCaJ1Yk89t
jQk5AucDuRknQdLoOpHAN0R9BEoR4g/1dxxQcOwWxJkbE8VxMQnn4NsCEi9ZUi/i
JRE8tOsJ2g9DfmkAaoaeh9611oiV+I/TjrpvNcyNzPHPAsF18SrQ2pPqThDP6kkz
+SZFXtvFfrgwy4ygZPLqnWQy9DPhF64LVXCIRQNoZEyrMzsDTZE0DYfoGZ6kOlPu
cFOzunx85miotguf/dcF5bexAnILTr9TCj/CYsi/sh5vfhAmU14uD0cd8X3vpLrQ
cCuYLiSVBet0rLn/jM58bOKS3frUbZTqBspEg3YpBDrlCxYY5Nf1jOX1iEtkYYj+
Fw28H7bv7CYInDsY9n0JoR43S+YszVjJwPlxQWgiRM/m0GWI55LpimAu6VJVleGO
F9sgQuRIsRv0HiwacIu82Qq9nq/heRWnpRFimGN043BAeAYnDaBCJjb0Ve4wEMp4
Y6kATC7I5jlhrtWGbA79AhomzvyIg9/FS9hj54mQcNVJ29IwwelJ7ypZY2ifB/+O
OpvpjYyILGRnoPp9j7v8NhwMEACnqmTnzbo7Igg3v4Zw3vv6aph+OLIp5PY1B+j0
IFqKn1WgSQg2afjEz3FnDopu8Mkz7PlsGcK5XxoWVUCdqZYu4wc+gvGvmYn8cxSI
zS+sRGpRWHSsIucEPMLCvD5scqXjXBYQgMDKF0o1099MOz7BpAkWZOdwZxhIDoPt
F/x1OIlkWiHu5F3m4xpngpa8bTjQLhO4zs92zIKl/V8nl62OY/OjGaWKz5OwkHQ2
pjB/6hpWtJ/98MK4k8LpB8RPDBgIK42mF6w+PmazGo1FJ7/mwgmAtTy/0VsoWvpz
uGYuYK0Cf9okQkNkfZiQCuO1wY6zp4pSVOmzE9jSER2HvFW5kvoaG2KJOJGvnEkc
pBODpMG138Tj8DkaMJYA+bGs+ayXSt5vM7a/g3m3ISVyoKIUfam3ImPyjmxJnmWl
2Y0AuqUpu5kd9SKMc2GP1qVsw+taxNgwwilTVgidASBRpMvtUaVvLOAmLil+wlSR
it55YVl+bKexY83wADyZ93a/7YQWyJpmZTN7HqTFZW8ERmGZB8pPQkArDcjMeXx1
ElWZhn72sXw2QF/EQaDljk4ebK8HBmnFpYSnh+nnXj0wm1Hh8kQiDV1aDMV0UsLX
VsAvnLHmOkIFmroHTFQNyqYeF8bq7ShVSYHEqIW1gTauQ75atJQonnILKLNB3C2x
zSQUmQT/CSZkSkQPwwXUP00oONpMaKlHF4kZ2UiiOhKnzoL2AK/Z/VQybiMvUQO9
mqVaIfg0gAMM2zGoNCUO2zGPF81GLUhZzFIV+K30wQuPjGWOEhqS1gheiUatiy+N
HtiqW1FJPYjCODGN3Ts0HTCvYCL83qVG4lYP2Ig6ElAXz6QQqsi8bt00uFFiHfhl
pU4Oghght/lYKOyBsO6dnlrceiH7lm9dfc0KAmlofpSogYTOSrTSiLacd3dOqOgt
oBmSBSwI/Oi6P7PEP6cHX+aRHRxT49mLhIiIPbozUFtv9zT28pebADjohaGwGz8u
Y8ueQqh3vMAEqP3LAS10PNDGgkMl1QYBD6sikPonIX2+JZr7Xlet0HI691AddKhY
Y2K8t3ObsMXYRx4qBvaHEtIfSvD7iqmxs1ZwsYcIeuiwA2yLO3ocO7kGVROj90s0
i9nWYKxzPbk8WYXFQhBLIR2C1H28MDCmmlwkK0ipSBiEs0I4OBJqvktZVv90eSpX
n82zz8scubSKePBtnpTPoiuRow+5mDCz9zlTjJedlnDcE2XY906ZBZhFcCeTzXHs
6vcGiK33kxPOjfRoXwFOExo+K2Vqsr1FY6ktQtaf1YAtSNkw/J257vQPTFRG3NEA
TKkkzWmSqUuLarRpqv+w76pBkO67d+CwPQASpH5cWUXX24oDAl9uA9A1hBRGHV71
p+/TssPRVqJxBupduno7JY+F6ufhmV5bEFIvWFSKBIbOBuYU0bDFfWFJ/C/r1Ouy
bI9+3A7nqJbW7cfcvKrw1P/GxSpjNDvcaLBlHSIHJRdcfFLKma4cw7V2mxPUCagl
NYtSNX7EBAX0aaOKrgl4ef8pVnugOZjpyNO6Y1azBExVhlI3+tfQsLb5buo2CYFK
P8XOzJ+zxFQc76nkp1k4OZMfcoTQUk+TjMH4hUjMZ0d0qzHktNnSInMchBcwS1So
4uYeroAi0yPFTp/iL56dxvkOoRxx010OOkXt8VzJ+cfAPsmZjPiPuFqSOHYpx8je
YAMdjIe9AJ8tDcOxHIS413Vc27vqqNvwkB0VOQTug4FFvXxJ6rk/MrrAHjVefG8C
NEDgVTPzA4Lr+Em8gxcFNjQ3z5C1BonUuhtXA0QbGnAEKOsYr1bi2uq/UdBaTzbg
8Pfp6819dhrHB66qyhHKL41F59AjbMMecqTRkmss2hA8c7LK+AtyqmPeiW+5QLMJ
G0ZvqkP73va5A5DgmEo2TtAbjuUQ0pt9gyZqtiNKA9Fu0c1JtUpG+df3yMuU220B
xdNsKO/ohJQTJCR+Vhf4gjyMSjG40YjjW0VZdV6P+5PP85ZRPEfAyXw8mFkH8BsC
9zsmbAZ1oMYVgqiVdYuVa+YABks+bBS7K+nNTL+gU/qjA6H3ZsHMOiEDPwUGoqLq
ixDnbG77TQdVUsuyTpM774W1xci2rE79HUUq+ItyHJIfLxKlSWNCEo3mxTTYUmFA
UVNMSSXCybWByGoMLrEAZrkSzgTFqkWs3d1HHiWWPMMEa04MB2RZSWH1LWSvm3wH
c7wnPoK5yJm0h08aTW/TsgW1VG+7OpueltRZ2Ob9/X3JlwQU4uBlJYshDWhBHyki
NEcRN7khkfTvDus/HyALM/srkC7fO/hwnPEYuj86WklYUy4GldUU+QrbaySlyEDY
W/B16kzR/SYGBn9LljlWa/iYebmV0+Y4TRt2KnLcmQN040qy6+4rMP2fiCMCrf/w
dJ0aqcJeCyVTTrZPy5hesBkNtyzHvQRe9W47gTJjMxWosSmOkC8dKg/92Pfn8QCm
VsF6hGlYA7/aAVWk6OtZ4WziqwZmxNUHExft+UUmqqjqVzcmogyLHhBQdOENKzV1
T1C0DE7sZfLXDADqwDkYWN8FCNgQVlP6jTY0LJq+h4AmP2/6PfcZQRqZUv/fdsYA
vuZgSmWw7n9RD1VC7aTIvwaER3/oic7gRW+bvzrPPuhnDGKRWqNygUEGi7iBZRZD
q2Vudab5LmEeiogreqELVPLZOnPsdLY6lDhLpkOx8OqZ+vF6MedRmtjPnJpWKhKD
GRGDuHGpSSuUxlNEiluys1mfE+2sTAWHoN8eQkPHH0NG26vrZyP7dwY3BbZ1JeFH
lgx89UiXt920ieZu8GjB/zLMhW1vSpku/fdUylOFPpL+v//iizje5f3c6Dg/Blya
D5V84S2GQitnVDd9cIeUIhDUFl7GHPwKwhy+FDok1FYPD0I/BEOvXzRmwjTryz57
l+73M0mZn0kzcCXQ6JBN5ygtUQwWYt36B5sRpoX907QOXSpf8KCOBwnQbG+3MvH9
RE/0A5Uqaz/Jdkx/Q1S7HVbtqmISFlhGfmM97hUxjimccylOVHvb+SWD6iIMwRGX
PIn5g0hcieN5Sc8zUqda+fBkRd53vPeu4NAVib0bkGwyTUePiM3RYtflTwM7GjFQ
CAdPZLAJbJfIs5XJHJvDUmMy04CbYkItoSpPGxjymvSpbNbUJUoA/vlmPDftLZ10
WCNKqVNhBCo4A/3rrdt2DTXUFF+0PZGEuAxcfvE/en6JqfODt2NOfymckxD4qNXC
rwYCLioQjOzOA0zS66fRKG1tuQah0Pji2LwE1Vd+yGYq/zM3YUjlRLsUJFxn5NJD
RsYRhc6thbyVP7GW0RzQ8wnwThuJ8Ax5bocf7tepAeBS4rQIe1dPnfhPkc0vHgpR
G9moNrS9tAp7Lktnak1CuZAv+wdvGgrC11+W7HwcLjLZNkIEqIqM/uGhERI3DJFr
/layC0xk7GEZeLaQGbMgWtZkiezdvAhCUaA9IuR1MwOHJM3dQ00aymE2jbK27uR9
BbgVA+o+YQO+dyr/G0sJnStgDs4ZWTATzlkzof24waxBJJbqz7c9oaO/09pW2/wq
mI1aiGd5wvPh1AO2R1ZnDuZceOyHbAX6+TmSuQL+vCsdj9ad40kX1DU1/IyMVdmC
8+7h/IUQlwhvs5Ynx11ajLrXCpoGJv8w0YoiP0X/PoRptiRVzl5WQ7l28ZUcACdf
/BMf85KpXHYLkQExoTs8gkLrMY1ToyQuKOT2HorNU27fZRJgugxCXySM2Sm5/HIi
mnOGDUNRtvdQp+VS9Xf5r4p52yBCCMFwDHUMTUqkQxR9WrvwZ7+O8IPMKbgQhuSW
EAlf7PALlN4PnajxzXQlXPLRCpqFyyzndRgFT3LYIfXtRNdBt7eqvhi1yj9DwVoI
wX9w/PmGV2U+PR7eRiTj8HCDOhqGZZH9WJs3mS4PKUhDP9cHAUUEWDzLAFgCBpPB
2GHSLIPozZ8dJv7/3q0QG/Zja7F8srQFUsQyZFe7Amdr1ozTufTHZUHjVWboeYL8
/Bozy+2P+b07ssTI+zfvgw==
`pragma protect end_protected
