// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:27 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
r9nn31KFVi+LwB0oSzVSDyazg7YBjD++tPpCGrBWa1fpabV2QpDLGjG9mRuP5r6c
fJZ8yE6LeKCzc9CTaWUHKyQAUgAmbJvBTneaSlfBiNkoSR9f3e1jvHNVFL3cI1bo
kCr5Cny1FlcCbnqAZkciBpIb4uyiKOeikALJ3h9d+fI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24688)
xmVEbwT5qm6rZMCVssTUkFNLkeTOEF17fMZmjPlbe7DNeeruVWXapq++FFtL9uJp
Hg0yqBPX1kp9tkZD0SR3mvmn9AuMymACPXFpkWxCSlZ9MlFphSsv8ko2LXo/tund
mR9FJR463B0avofgI5Sblr6R2Nsr+KHbIBkqB4uJDDzaRrLlXiRcxq2W0LN/1mBG
Q4U5ivgtf9wnUIRt8aa2vVSM2F/q+vGvOLJDrqGz00ZYChHB9JgOF0+xGaykXo95
xFkL9p26z+U2nngNzrR+ZcL7GfxnAvP0qbVO7NVN0eRigLL1GliYr5jwK+pGV6tQ
V63/WMDnoCzzKziMPXLAXYAmveRgEk/Ckd9ERWLX07Wpfeg2Y9yxIVZgC0V2JR6q
cOqoc6XfsL4/UrsG9PFaYuOMN1ji+KqVuHh1Q1VHcBVxbYBbZ+CeRCqcDraLj6IX
nYFG7BXgSDGK5/6nRsLptaDzbnxqEzZiUSTzVvhfx+22RrSOqlbphuQs62X1dA+i
pTUc8avJKVp5hu0HDdBoSDa274q0KCTbFmLyh9zkAhl3wdK9SgSv0cOhxoivsjbi
5kxJRfSmoAgK8OTeQtp+RIwwmEqnw9h0kKEwjWEzWgZecvsMT+yTprX3cNrC2lPg
pE7Kf94v+ZZaqo/EQl3lAM19x7MccHjRttG2KcqJ08sSg10QEcr9oGhDoDX3mqNg
fKkKvOgKEjpuB2PxXD9Rqz99zP7UQhgcDMpotdA+a3aJSePsLuxyb7/af6QU+lUV
+YIglWRfDG8dPeERHWWYgVl1hn7jTMe0KIhoT8uqOxWsiqdy/kQ69E4jrlGjBQZ7
NtYKSjjdcnoyBj3nbfSP712xXPCBZMsQItiIiz9U998A3Gn2Rxeu8S4qhyusuwPo
cwVlJpF3cVs0ZXD8I0vvIk5MT+raa4tAxrIUe9ACNkB/26tunzRdn7+8n/XgG2nZ
DP+B6tqlcUcDhBaA88i9nH4P5MN+FfT/TCoCscr+IR25eZ3wU8i0VKRlTicVoAlP
lcGk2MQ+GQFRES4qONfih2Dyz9dE94C+drNScRkRO5tBrBJMCiWrIIo3CdVEZ7LZ
dpmNHvZJc7ZMWxulQxDxbGFY0vnlrrqen6PUWUQgwgHn/mxy+wnkgu+TQLhPBAmA
XIZuAebibPAJaGvC9bHdnQq6ImE9Wle8ZlkqXRT7fNTMw7UWbdS6vdLbgOzZLjnp
hq1GEcUlHk6m/zvtvYXais9I/3CTQOSxoUDgq6CWn28zisLPTPyGqN6edweA1EXH
6CNVD4MhKMtyWNxqBZixdhti+VKP1+UGvyEm3mwNvZn5dYsnIZ7I/yAoBTHyikcJ
GsJJDx4g+i0zhrIqx3GkXYdqaXwnMt1Cae/4RpcdAd5xJjCw4S7WQoxZsDMhjWcI
AvXKW2mI3GWiz647otug0nWqJhBWrgrj5Ea7mHgvGkTTrnKa7kxOe0jfnXuBN8u8
jmSWIwzMK30/Zl4G/J38dZt2y2xjLhQdia95ctQX5qE7l4p4aLB/yyTua0Ycr71G
j32DUmxKowMAMtQ89VL0hmcLPKh2rmsjAyaPXmpxh0jR2ECwDvP9oKsSPipU6xQS
fn62A+M41omOz3J8n0JfQCA1JLIP8B1o1+aOlXmGOAwPRadUu4qMqganbhuBvKrM
wcZqEt7tnHHFeRW3MBpxN0q4YU9eLHTxmsZf5uf7I0zgVhpifGab1AEt6XbXUvhD
rsxiFy0ujNdViO7SpP3MX5Rcs17mhN1Gkzqe0Px5YfA/mBsRBz3T0ULREO1tQItM
fb15tIYJIBHjgfuayLSBqVhk4GucVFlT1Oe40+MHYZoTFkHWJohBKpPGoX7TzG9i
7aMl1HDC2J8ouh1uAgRYlI/EQ7Mnx7PB/2Uh1TeE6lobWjrIwspGrEO9RH+RZL5O
7vMkiz3KbOZWXFcrFKTp1+3ck8xuY37D8yZrJivpvTIgADm/NnLkeuK0KW8B4tJj
rJNU4mkVqtdTwOcwrQadctYbmH7wGhbK8g4be5MB31EgzdwCLkIWyspNBguFxtz7
xuzUOyZ55D0bKUDcS4+MlW0GdNXwmx3RUb8j+03JPYPpeb6vbAAMD+QDnFM2sh0G
4gvEPxzp4NSSy7Kqtfo2FUnJsmB5dsbl6zNTeNHQ/43UoxXAmkz9i7RyW49rP9qb
NrkWx8aHZEFlf950jECy0ELF+hSmLCO6qVpnM6faahCszv6pHzHydsffczvy/XJt
4Scdmj9WW3q9e7iROGpVXPM29GzHThF7H1Eukfnf2Av2MKP3QdvJY2Rzub1ZQcfR
8zzfXS5bBuEiyC5fyz4eWAbHSJ2vM1sAMUvNTbeEQrhBNmYGF9LIpUfVF34gwPmf
VOvpLhsKCuiJ2/tCYa2q7ekKKY03PYRJExFFnUEpnBGAYuDVAmS+14qWV3hkMDzP
pXDwSY0YefyC2gPE9Nje23qeC5Dbkv0KlOChfRpm5UKO2JUrmZiIrj95mowQEP26
Hh72QlSWyKh4aSrtynWsyKS5+nnrJw77ccK8wm2vOnMNiy6hchDkRv6FkPFxhywv
e6KH1Q0P9oufT00JD1WMlYDjhZoBoPs/yvvQr/jcndgxNk2zWVBPO1rQVI24u+U0
+nFSoY8VhZjZ8J0L8avq/p0SvvvD1MVCbZJ0gBB/VevCDxcH0WVZs5VdNUi4X8r9
4YCneogwM4xGW5vZEH1wVCYiErkJh+79z3eO/6vO3ryzYVeKjTs7j8xXVtpsAFCV
lxyzGzz0Nd9ySTT9dlIyU0ubDkbY2+mFPosCNaQtBYZCDVva2Rw+r4T0trI7y7h9
naNSZvKqeEcHIjdISM8rHuSYTkojbzKsLaNRh15716Q7bC7P9ubBlFZyreS2lEnH
II3ZMUaSeF84EFvy+/W96BsiprYs3vRjZUtXWK7Dexa/VAdsKrPmTLGvSXlyQ5cS
go80uCc9yU3fWBVcRAr496e+hXaYeQxS8xB6FgxAWEZdoyailB0ax3Zi2mdrKFbU
bB5PRoEMCMAvm7uT3GIjM88mzHLW3EODabXWT9+9f0NpmSOzxkzJkLxbOvf8ipE7
srFTS2GtbPctw0jhjyDaEODsKHT60ZMCHcTQ37euk2iRQh6FMOBYh3ILkf/ZG93/
PspmADcRtSW4QX0BYBGan3T7tlXecxIoO1Og+hc5N+Om4zLwCWh6RAg3i8SwZNEt
kjmD7tsLIIAXrgYy6KQjXJQBgGAeKeuIo4pkGq5YHKUXNKFcGKDa6jJWSsStwvyo
3p7HdrII2n8rQbrXwQrHrMh/mQPZmh0pdv9iiZogXEdbZpQ/ELl9KRA9jzZSAkUo
1KeW6cdV/QiX/hNJ1rb3MUw8WqXf19zHL/2A6PzWI8rymoPNXisUr/Qz1pC3uj+K
geyUswQhL9XjnjogXMdvUax7MejOPh61imJRAP0Q+aukhwxggaqur+05hoQ2o2rt
w8Dc+aWGWpTM+l8wXxUDmmoBhOZwGPHFy4ZMrYVCAhzF7zQJizn6kHlcgg5wlHZL
CBTHuQDbOyHfWiGt52Wsx51ApgA6nheizJ0kQb3HoRBDRUnx5VT2KZFlmwboOLPY
Dk/l9BtGzCp3M04ypf7qnXdnrUIE6BpTPvtU00bSMhRtliB/PVm5ZGdr1RpL87FG
A/p7nbK8O+RzRJ2ow+6Mg3/1EGP0IRKT2PFI+j/hD7gm/BIq74dItAm6Gegr68VB
yn/tx4EMFgi2SOgJ+CGWig6s7zmTNJznS2YwXU1JLqa4MEgVi9j1CEeqCZXXFK8z
F3h5CFNaslxbMfLjLx6nV5henUtMz1hxFnLZMcLMwIEHR0F/QeZIi1Qo4LFPBYv2
lDM9umF5XB0iQdtKINE4bx0rDhEpdrIXzJs5S8DJEiUPWPokNVUQESRScYBHuHl/
BvspK8RuZmVvGaTOjo/iQnyvuVPXR6Rx3fVVfatBBF1U6elwC8Vx/MXUBN+lALXq
RztATdhLuNCip8qoW6etZUWf034/lrT31HAwujUC/RokM4UEjo8hiDSrtvVW5kO6
l/7oHa4PCem+WctWESknAz9oWdIo0ROctjw3TTrZTaXcmXJdD4BEf3c15nFGOa15
OQkKN9wgL/p38CO288KnIcDqqIAEoJeXQVvlhCtHapl+uwaPX82UHO9jQ5CNvBe9
K1eVMuTxqUG8thfdQh3BbFdHr0UugQQsVdcRCYCP3FULtv4kqs329ch5OjmLnhOJ
kuq/ylvwyEy3E7Jab6Mq3Q1Hjn1ooTw4cnhogCm5ray5weTkEyCirO90YW9xsblJ
JzRJhZN9RdDyuqC+pSp3ea0I1T8MHyT8XmQCoxFhqtjL8PkOZdZqHbQHr8uF+lr6
mO+01jvaFKGLhOryHWU+YlZyHPU45Lrdx2tRwNYpkqbv7QcUW69OS7SBbLzohpc7
dwlwxPZaWrJLV3KgsSRsrlBx6nk1MyxJizYWs3gKharMbiddcPFk8vDiom3Uevpf
/V/QVgEcXE59MvclwjJ+cYMTggpxQn/9Zo8ivGJXrjXiSXMxlTT2nWp2LOjz3YaT
rdmv218SgWmTBl33qAsEIOXGX6vm04FI73WGgrZ8G6B7RejaXX5la2yMj3H4m9NQ
kHeTlI9lulRlcJl8OOymvTmhzILHnUk8NPt7XXb+nePhT/tyS9wvKJH3wsyEV7iL
M30GGUd5eHy2pifjaKCLwaf+WEo+aZ14siSmtKhsaZwn8Y3bl9NM0qdJ2v8vcEpP
FCxnouNO1p3uRYxsyroait1Iw/16yU9aqUh4It1EIiyk7kA34F8Z3O1e6pIacbAh
aVqT83mZwvIiwaD+V+8jdh8Y6HlinnTmFVlG1WvBX2rAsQpLYTRAVuSyyTlcq38D
lo0Kb5tH78yxCVjMKtA5DvpmztfQ3BoxoWenurGEWVsCV46LL8LpJkIG/WH8vfoR
MHif3PG9rVesVxY8dMo4bI2SbvWIPnaUxVrbjeoHb1uS2tHgjeBlzgn8d4kvpCPj
5WkYAv1GU9jn/yWZXlUGpVfp70IFVOfLBbvzkbdZl1bKFlmckUFWvmhRWza/BmBO
ez3tB0JQrPXkll50L1NTjBxqQASEdYdXqepLSs7LAUIxsG816VcnvDSqYRElKvV5
4PaMFhTCZpZ+r13zyLlyxNv1mVfy9EMJQybfu3I8/f8Xghwa7ygIPU6E35gni8Rj
ZBMyQXCS44yBGZv5pMYIl2l/GdKOIoyin9uvqO7qD5WjPKEDkTbeUTUU+gL0sMPr
VD7p+Xq9GDQ3jNJWxaTZdsT5FECB9qV/XeWwqj2Nr5p+MZvirOxQOmqPE13FPokg
SCDMIlvyVyTZBEeG3o4urP0DKXKWlAJo9cMQgt5j3AX5LBY95b8n67DrqaBBC/+a
GtW/dvSTISqSbwVxqb3tGV3TZy0W32Ieeq3PCnNMNW0KN+PmvSYwP3isFDelK1S0
Q9ZdkAUV6sLs4andWiI30fVOQcPAjI2HvuzD76fy4HZrHCcMydhEsATGaPPbDKY2
OU6Yw6Z6bGV8ZvnSg0nBQi8e3OIutQw9iGcmEaaXpg7POE8bMkrh4HI1hQapaEK3
xW1FoIgrItzg2TaUGhCQQ7X2w1e5Awx4ttg2rCjIkhORCX8m5ap5T6HAGxFizkg2
kNeRvada7sHenlWoGakBUJ0Ot6HV2NSF5PUR/nqrrIwDOHUfasofH7CqTpjSBUYN
vkipYRv1PzQCzaLLpXsjVMLB+T2GK5NJh/mO9N97Px5b5YkMxPPbeBhZxytuqGE/
rF+u+tgELVQSNFqjRL0beo0B19a8RzDw4tvnw7D8qNkKXEO0wwtW3pjAFwUT5Yk8
5j/iwvNd+2tVwima78mkSP7VXtTefz7w9oKw/nCHaUX7Hd8HDhAHkViH4vlwctoO
xR2PSFLwdIa//TrQO/tfBplOJAmpPUy/PT1LR08hWVRLfNtx/hQ7iZHehc+Wcltp
4GfMFGlJpwlzVjlrn4Br7B3PPcbh4YhULbOOfbXLMkgDTaWGkWrZsmIUOX5SSJnb
iTj+GFwBXqOHPtqrhWwSwAxvBEalB7BaSu4o5dLqYnrf6goaGNoZPsbPERE0Ff/K
hg4g/qIH1iZaR22sLis85tKe1buAWcXupSd0caJw0/X9wwDdMdMsMorJ5x2DcUBc
P29hASH7XsQw+8rS8M11JppFMvCMdPDtp21N6SmL0YFFauQJlso7OLYJagu+0E7w
TqA36RA7yccFWNL/WOFgUSbpg03VulW2YG/T8uD2PcKAECWdDDEAfix52DoYnNyc
b+lV588G9/TvB2u61L//eO3Yj90g0VRyoeF/CFHY8lgR0BtGhw4OqZjCRseCVeD1
LF24T7Zg2LjZFoDdidkkQmfxHgMFJHM8EiYJuqHFNXlR0AGIl+ntpsxZhqSH1Nsd
jCJFV+s2LEZ8jWGupzf2zsoSCXvsIT5tk8+aa+ePVd8eWCh5U6UCLiSr3z5w0olf
ZCp9VwAnRnWYNImTdvzXIXIcUlOW0yRRZs9uC/yr7aWWh1uLwPzprt00BIUVfuD0
AP5VElldVEg+tJKNwPxVIw50dk/QV4MAJLGAquwWSSh2/JVBaH3WgdlYzRC0kdsO
KcJ9bLlVB2xk976s+WVIo3KLhfVsCHTGZBaUxcT1Kq5+AnrnP5xyN5unrZY3bDop
63TCINUC0MVXq9Gp1bQgZR0KKVqrlCYXPIv9pbKCe/qvqGOmbmAFV49lVtJ1bp0L
891JvsLUj3tJa2kPphLposnx4l5VYyTAk3vSdBMPK++3PfEjSP2ncqejLlLfFrqY
9ckOZKmmZ55VqDcByTymfGT9oscumzadGQ8CgHpR0Oncv75doyXoOJ2iTBW0jlmF
n6z2SJFpDquvVbZMbdidY81xRClN5qqqrSyMHn+mBQoeyfOzhJl7LqJ1i/NspVIi
loWA0MLinUSVjXqtAvXHuZt1kl+CHij9rocCE6fapCatpaCsgI9SkDl6IigAFof/
ziCFP59fIMm38+C1608oSVa3J/JmN5nkn7riGCm5FBEETv8ytqFLdIPEvVLJZBSN
h0OGsJmJkpybYyRlsl8WBupvM03w3EP8Q7t7JUw9TN+nYmwRODXthJoiUWjnN86M
SIgf5BIOzCVqkNSR7IPNNuJuZjAOZ9zVNS1sJt+gcA0ddT/LOXQy7ucBBnOMRmmK
fjD6xkHyxlGxK9RkcGVdKwVVfyxoVJMQWVYXhi/vCx8xhrr74yBlYjd1C82sfQwa
CgCvRT1sUSRbK7d78AOMFrugYJ4VVBHoysb6DsTQYWQlqljaajcD4MH56EbR7tdB
7cV+xDz5Jg6nMs7GispBkGNkICqACLiue8Ww6HiSldTgw2xnUmufS6gx8vIPG1Np
cGxC7hiT5wDp9mX/Y0sUrJ4/f4GiI2shzsDYdsSpOmCblR0fQc40WjMUQs7A64te
LgLiL1yfUafOykGHY1gy6FY8wA5YnboIQ0XcnP3K0WPdRqn5GXlB8GeAh/wdwYTt
wUizylD5rpFoXH49C6h0+U9L3kJsElIJVMiQiWFpRMCRlJu8CK+DQAY0jweExL9X
iSR0X5jOkTyMf3I3NbRsOt99ERojJGeXNh2u8omuW5sW4LIyvufLXdkYq++To+2f
mPCwRxz6431Nw2chprrCFg+hRNt0uq96db7A85t5mE3m0PRphHD3iCVo9mwS1g7n
8ofnVmd4GmajD7MqH8/XgfyMqsHsTtJ77SB3+xhKAB2rZ/J/l+d1nZTetLA9V97F
jH6jjInCskwSP4ZCpC+dMIFoS7cjpte2DSDJZfpdi8TebjaXcm7PTQRRWQ9JnyAs
CeUygUvvMbAt6yZPhdubaa0dlb3RqgVJii5EbPUewu/0y6dvXFtIBGhh/tM7CrTy
4ApoGMs8n6R7vfgVY5YNxu29mOors4EeOjbyDPwxMKKR6ji/PQQIDeiGLWoZMMM6
JSQQQLX+L4P2V1ve4Dwfk454nns9Wi4AhcFwsmuWQHYj4POf1gQ32AEfOsc9L54m
v3SX6FUzGRyGz2vftKYgeJxM1FafhNRqqxsOM2rbWvdtISEE3ANNDe7nsH2of0C6
4QgeIfvPcxFUdzTBGH+7DaaODwYqQCl7kzcl/a6+ms6SHI4MRKTDvTtjFXr4PmS8
AjfILyJE68p8SPo8++WUDjIkY5yp3RHbEI2PZrin/kKAt5xZzLxk5kEkt0D+x7up
gpOEs409q2ndUYBE8sxEysIDE8wTJkW24FPwOcoMoYaiPwsH4gMqeYOazwR6mn+j
cTBvSSwmpt9b5EmBBJvKiwvl5DvyC16LJ1ZXacQjEmWIBsTYnyDp2ZeMtYe55wTV
jXk2uSAhSh3whnJaiIiLwKt99xSoTR7q7BHzZAkuoRsIhZynq5NgZAuzP6p7+6fW
F3zBKW+COqk3RKD4U1beqcZdMaS+zG/yLEeAvHDAwolu3VJmZZQQsTNNOgljhUHw
RHzuPzUNx+lhQ7V9oBCV3z38Jyabtlli3V2EZWBz8CWSx/8AKNSt+doOLgxYqSVE
hSVzzYLcGX2s75LsUMLltO7K0xU1K2EbQod/LAjwEL1neg0FFTkSy8a4FO/KzMIy
yzx8Nz2QXwCYtiIys4tpg8tCavAyfiSfKJre3JVwWd8V2WIdjJkKRUZwhgU+BKJf
NzZuJqcqFS/c72MkqpkRJjug3pgF5eIyCKmg3VTIjN5qwPRdErfrtJcH1HEPx6fJ
nVJwYmMzbHrUWPDHL8FLORWQniFJO3NGC4rAqRkbGk9gu3NXdyGMUhlxuYGZulF8
/3xbSuWZ97p1ncLdqNSymGaHfCeiVOQsEtEV3zTU+0fiEyvw4cippG+XmtxMP+eo
yUakPPMqrGrbdGbC3x+dFPwtUTvmt7b142lOJqi6QV4RRaPbLp+0A7XdDlnZATUH
TbrghlFTHUwOOT/LleS5Zwk+Fu5GCg/Mz98AWCBUjSzklDc/wm/r85Xy3CXaDOrU
dynwqV6HXA5ywaRWLwP6NhnEI9eXtu0gCEAMIB4fCGgaPu4OawRjatZbm8TNCUkf
GBm+MRiwz09T7pJBciCsASWGLB6pTugymt+gTQZGQ4KnOVPgU+eyh0wNcxNpFpJD
aVo7wbUK2oNDiy5GZ6OvJEARpqcIxfIJ9vzr/h1/8iqNVw8GvOFoBMwOR5oyqDgZ
7SV1ecXFPsuYcAdi7GzU2JBltNDkQ66RfD2un0q724bs/5F1X1IJvJ+4nyK3f1H3
hc93rH2Pb4GEeYOAFjw2t735Y5o3XILNbXscwWpuWJ3v4MW1TgEa3WP83jj1RNeB
nVBGEpDMYVOpmI/E7Xqo1HQTZR4bFL+njczhQOqX/QxeuQYHzzJvblb3JPWBsg/n
KaqiLXrxggkkmxqk19SvIUqKIztTMxvlVa9QPPJgb1r0nXVewzZCh0Kv5bD/HaoB
aKwJWzPLSgzIdUWkGofstDatWCH3F76dKfSzOVo34OHBLm8P0l6QsxONTzU9R/+1
4jrwZ3ynOsXpsMBf6FgZZedd2U+n6YSKEypaZMsUfoeUwawGnyVok0wFxE1kL8Ci
HL5MmlKPicHdKXYH7eUhtuSww+3TOUc+H2z8HKZAeBWI2IymmDvvRcvwIgJfWxAu
i+cGXCV/BnP+/yTwHsk2GbjcVAv2AIfxkebmETrVZE6VrHxAToYAzPfy0ROZsiB9
iIVKo1Qv0jzCf2n++/sYioZ93lwZI1AAgh2O+3G/4rg/2MrPZjFCT3+U5K4DBX9B
6QcL84M4ccN+KC8GAtjaTKRIJM6g7SqbC4WdPoJzJAMyBoFGP72VuFhm/c0nAdsx
ofbx1AY9vjS2wzRJSY/KWxT7vxK/goENxqRQXmZmcSZGlADXs834miw1NxHKmrYk
pGDZWSDSt6dZTq12R2Y0Zz06Fea9IH++4XYXBoQqo4VGFENcMKRk0acHhu8R8ynh
4/m+dUSEAX5K5rtncMtyxNsXZ/nSTevNxAC2Lswff4buWJUYitUBwQHaSPv9kzhQ
bpmFzxBqD1B/vE63NRnc+peN5V/gU5OCwH4ZM5Z5QT4EC5cFnbBWIItJ+d8+RtSh
GZwriTcfytrtzbhpzJPBc0ybWlM+3pD+oLbATUf1cM1eZkUbkoZZmJC5PNM24zCj
1q2JDroQofHdf4NiC/HkC/3PmRvsHowi2uKJNTyEb2jlPr+Rf7NQFgOucqsucsTX
/Sw/y9FBDvrRy50OGk5TP7rOgHGBL0S8aNgdbZ9VyeUEjGJVox1QdwgfGErFNki7
gWJJTphG8B+ooyYbtzrVuvxIvuuuHjhy+T8NWz58ggkBF2o4t/MyuMHisH5Ht8CT
IYyTi9uQj5VypZ9lcDt6/mENUqNrVvi79qG3qHll29ijqX0HHuUF5AB85y4NsC09
ljaN3lj1tpPCmO/B9D+TlaNLc8YBlMbO7q0PpS1LeLoKmJ8ITSB6bOV/gvjRNoOs
iQkS3c+qzmd+hFBW88z1QxeQ5/rXd2nDKfI+R7yoYrJ4D9CKyKPfaropyRAhDkvw
Ioj9PM5AwIBu3svVC8b2VIT0LNcdzdy1AP69qLyVw3DEciGFJx0w2r8DuK4gscmo
lRtSHJT2YywjgTunzH0jy6gaOXfC7n7VeDouehIC45uv1WREOVjuAoSRvi0kRV7h
F3OHIrMnCrSfZOF52jBZ7yDbaSfPXJxvGTjkCNF6nw7e5wpffsZHDlKx1s53jmlb
0wR6Fu32kluUGt2+XM2TbK6bbfyZNz/Ldm4ZG2H0JWEczQYFZHEz3K9kZHEVWCjh
N6lL6QcOfU6FG8FR2+7MIptd4mn6U0Jy7Lb3n8EAqkoS82MBm//IfrRrgDEVkoyA
nfyV6s4kH5GFwoMMSeS6huCNkSKkFPuIMoNoG66EDlcDAcwdIh0sVsH43h8BsgxQ
LKtfVxU4h2aBv00OZDqSbXoZ6ezyQwrbKpFq+7bkT3n/JEgBVKw4w7vz9SMw5h1x
8pmMhNKBnrhm6Pw/3Ol4Fo2USQ+tdeeOcQjbEYhNDJbwfphCAUFsAIevgNKNx/Vp
zh5bb2evSRI/Pr8+6RKlrXIPav9A6LRsjDNvEJxJUw96zcJQ7GOm+WvBzTM9MH7t
YV23urMPchwI+XksoHn3WgiHBhqyrJfwQkNHaFSYyG79oZHPKOWP0WsWyh5YJtWy
RC2VhoFYXaYbbq0a1YfYByncpLRFd050gQMAeMyxDRvnxberpawRM28quZFAW/Ku
nfrWW2+stUx9yAZo/MVgX01/w7fol3SIQt8fEBNMxNe3liNvohWElL7e0VcYiOVr
SkUb9gCTfyR36j6wi+jq0x48/IYceZG3hWzGmo/K/mEeYKcP8e8BqWZ7jZx8syZ4
oczLGElw3NnHKWY3DRp0uKSl1wsR12aIWt4Rcga2TVA7RgHzbDaOEnYjmti/ir4l
exelRIZDgpkyDzuPWPS7nwDSB/l7YP5wan2K3B6Yp2e9fmmiWZ96FXCmKzJiuS2g
5ylTOTOqlccA2CKZ5vCwne5otodwDIzGcWu773yQk+PsU8S+k16Kqyd4cN4OQQoh
mXmMkRE/XGoo4Bp2G9Hjqvfa33tmL6CxqYsxs8r2B6ozqRbFOce4gqRhpgNNDoYi
NK2PS4+wvVHKrLyKw2NxUkotrnMRQrZudn2w507LySePqiuw6Dv13V6qbD6VRByY
eM/YWHPaz7Lund43M7ZqfAAePAjPszX2mvUKjKoA28RP6eh9p4YmuJE92CTrKStA
5yOVWOhnk66xR8G19V3zVy1CoCkHmcox625gs1y8RtWYz4zlbNgGVkWT90Ems5B9
aUrHsYJ1dxobvauZKuGv6kNnbXneoeZ5y+ydvLXKy71eccXYL2FDZHVHTIzxpPDa
mnflM7SjHBbpOYdJhVf7FOQv5ixWmzr5rsIXfSDWC/8OuK4RDXO/FkR9XG2GbCPE
NW6SK055HD1I/7jboBabE6R0Yi1aPBRz+O76Wm+/WMe3POe8KqtMPhRiCrTwoYFB
Vc8T4u/ieD7QYO/8nM7F4BFD4qLU9eB7XZkjjnouN/Bo42maRs/JhZtbqWmqHYKS
nfGem0cT+JUAL+xrHBgCyCcKyNC8hXZQ1p/ouGrF85KiRZ4hygJyAYtzn6vohD6W
5JTQrCs+zy8tZQL2l46J23fMScWjeuTmPPVbLtyueo68qCDHEaMjcSWYfCPZX5Q/
htqRTzTytYBA2SUPrKOEAhtCRhgQkkx7T3EwktLChufWOY7ubStMREFPcoOAdkoO
bfYK7SV6Tml6R9up3C2eku5w9Qabcq95SQTaNdO190NPo7XK/Xrbaq2BgoR0DuTL
BlcnpTWOjBSa+FGjszEiqJ7uV8P+lg1hulnoPpfmj9yjtmCQkkW5W6gpsgfZpIs6
WYPz8JwYyA35CrqYfR543XBazKC5f+TWA16EaT9LF6klOxeyhaRaRspYkamekfig
0DxmT1XsBe3coMcwiKWr2Dc+qL0nNSJlSMydQlpO76Bg07k7yo5WFFQTYc7umJe/
eutVgV3HIdtuaUZjMIGjsKlaF7SzbMO/BB2O/vI8C83wD2WGrCYnwYCLWFogGm8+
XqVPdT4lesQM2vs3je4epvDY2/yGlp0SmWufC9I/JND7EsSlGaOw0C1NjbTSDaVE
mjvEXVvP/ScjxrpvdXzMAHJlYEnnDSfxsDthWDMfMVByZAXBX8onKid6CDCKZdxt
FqzwFziaiIoizp+pHT0+lBiR3xScESxsXW6gLCjxcUNH4eZ+kHZtFQgn8RZ2bn5F
oHox3pRu6/H07XMH3R8WKgQ0bzY5hEkZb/spTagZUR8457nR67jzE12gdF6C9L4s
INYXLA5vUiIvolnAWXSQ5o7vh59Oejiy4VOkOfFAmvaXqnrpXYskDZn1dild9w1o
ZeqRsSyQq7izZ7+97UHPiIOVSmeyovWDPyQrAwdPb5g04eRN+PMwE/LwFzfjBlr4
YcuPJ6rwpDVRRak9wAXavFIqSX1Gx6p9+luVlLMGNpPJ95RAHclxsD4t3dchUX43
ogHYOR3sdIjoEjxb64K1iGSyLIwFagjeo85gNZDpvZNNBRs1ymIC8DsqAkCfrBgv
gWeVrQtXRg2+/ikD9a+MckFtxNeq/wKJSpHMVenxkiryx3TQe+sxrvDLIplhaL+7
JROBZnXQ3MCJIq0m9EaU998X4UTY5j0ktRPdbEreKxRHyGhkl+Qu2NDkVFKOFyA3
zc76afoWSTufRcDRSD1HEThn+fT9ikjGJyunQ1Id4lMs7wNhlHtge/5Y7nW+zjQM
IKJz+cCu6cTZBVa27MW7hPzqQJgptsKHN1F9e+Mq+eDhOkXxcVz2EOaLAXt+QU3U
rL4GU4aMoH2ENZMdxTOwGPpFPLWzf7oxkxr4C6pe71kBDirv6LNvXP3INrL+q5wu
npph3W61mnueaVXUg/vEEhxm9iDHumfFbYjTsDVSA9ohyxb/nDftwT+WZeAo8LDW
tjE/mnm+GI8y8UuN8GYWxB3Uf0u9XqQUi6isqJWn89dQVGTTl/lEtMaOMWrtpoRJ
KETgDJ46AaZlNXxyprbpKxd2z3Hiu0NAA9r8AEaGzsC99K+KjSxpyGnBSGuc0pig
OBtG0xqfBeawhii+IQW71kMW8RA3fYkThEH+NanT+tz7UibMV1t0v4q9A3Y3VP8t
yTs4WbxQLjPbxn36Ocn0RBiOfICTR+l9CGFgvL6Hb4kxXlRi4hm1krcsNYQbQ1Kw
b5VCA43HzVyNxwdwzQkiesye4DxIZ0A2CKKEZCQKFGVNZHZrd4h2P4OgInUTo3cs
cBoNethDccUjJKF2XC/As8wjAao3wxjkuux1MK5C0jRWapjbaDJ3zM4VZvgvELwA
WedkEG7otEiPMWgsPiW1oAiVh7MLZrma8SdHezb13yKaEGMzlMGs4L6plluOLmWO
CxSR9Du0brwBsXR8BMhpp+V4dPyV83Z2ddKiBG5vKRAognflmSD+eEE9Y9wqhnYZ
SX4hp0WN1Io9lO5UsuBh1YjoYK0HvHzVJnV93wmtrDmvwKWz+dO2U1fIHUgDEymW
YxBluCGYb+Do0T2YKatsmzR7w63q1DAigl6uXYWCy6KNGD0iWO7jwXyWNCveqMfB
MkBAEvEZ3xN6YU+dgIGM1U79fX9KKH3FDGBhFiHQX1TBV32e7OZRrBu+gyZsd56e
8RMBX81SMXBzJVaI/EGN6DYmyiCy34viGqjtaKm2levIYWwmvr+gIhu3xGVKt4rW
AW2Ph1c7NZxeNCyEOMgLwaBfNFNnqlKtcCegAJz2pQaa0Rc67fZwyS+kCyyOdErA
srunDi6AfegLdurFr59Jpbm1UpUw8cNGoBp9V9kFkUc/NxvnF884IVxdCU3n87ZD
hGTb04otkzYjAHc7VrvCI1t2TVRiIZbSZT/C6IuNdLc5OmIaLFgr2d9qelWU2vce
nWjaPOoB+lllFiC6bWwxAOj5LxX1e8FYvHkYpV28McB8VW9HFGI2r2rotL1VqZRp
6NU1Oxqqs7x8Rxz8A4VzakCFSFLnK3WUAt4DfJfz2uMXqAtIvTwV0nBpgBlJlAka
l1K74YzHAZMuwhaio5DCjrbqPNu//VBpgAoLPkKDqhUcG8H6L3hVgijgy4fz2sMW
9DvSTiTPd3EDTAFMU/Ok3OBZ9T7ry35LcFAxOp5wjKCL38R3YvGP70akgbWLRDpk
MpEX5wl0ZeXIGc0G25DSclMeZQGZQqkrYElVjvgYFYqV4NBKaC4kL41/uz2GqaGJ
NhZ/mL7a8oH5brQHUpJLPhFtWuLW3GR0M0yFJY7gYaLY72aWc5gl+dWqSC8INsgm
fqzkTHsQOtnKMnh1J1Ep7t5xqA31SMcXFDaf4QVwMgZt1posH3j4t8F0odqoNUd6
05ZsLPczUXuWx7/bMyVsAJoKFF65n1iB70/70pb6tmckIXXnCY8e6e4KusPguVPo
2jG4UzaPoXBPLa63cicJ86qLvYQnl6pZhkk9R4jO4OOfFdhikb8qsKLBul9zhFys
s2SNLnHSH9AfkFZwud9Z9F7GJFWXx5qYhn5X+PGGRcZFAyx+JfqHFhg6eoUzcSb0
7tgx8KMbhV1qAGM9ADucUBszRfsRpn7rzefZ6k0eaQ9zGSMhif2IcUh4Oqurt42f
qbKMe5en57Bkep76hSWziM+l5egoCcfUcU5sRDKGhpeb+ix1FYMDC2mDHBwxfksA
UCRbyD2EYaAOJIyir4fWCKq6sLMSLLyCsGP+IG1lINpsGW8nst6jIRy61ZjRaCYC
qU+d3Fxk3h1MzFWTR1gAr73NYT1zqPkw3/pB60uLNGLiwb3I/KkeH0UG5v01Qgwg
UX8VVFFvqquLU0CaP5LZddks94Djq/i79iYuzKw3iFbETw/5JI/V6wzxNKfhUTky
J1wCfsoI49eGGPXVB9fwR/XF8WCaqW4PUhMcGgVjmBKOyTV1ki1ILYUDxBPY+M+E
rxLNK+FWKjru/DExNUa9mWHN3GgwLURKXrLHugWY2YidfAfQBj/2n4LjBDBLVKDt
MKR6TLDf5Y+Mbn9P3q10SaKiMzTQPajCdSnwQVHn32uoa3PjL7czY5krSxS300yf
V0ytvMLhUJtkCj4EExjWdX0bPvrhGXC6qmaBlXsfgAJuN4Jn/NH4RHdnogVF62oG
dgQeY48yZ68lXd1rT98muLrCUIBJ3C6WPpodJyzjkj4x91WQ+9c/BiJxmnHmhfvm
iFugAwX4S1qarT2aKE2u+ItWBOZlYsIplTaQiRLsjjYMPsnrdyUI1amVnxvxW9fZ
f1GjhytFwxSmfrIq7v/1w5kIrVGn8PMAQwEGWwToVZXR/Vx9BOOK4+/BYw2mguHb
m3wU+MH8e2hJ0mtvPfwfRBTgpjX7sV44heVx+wwvnFTx2wcB4YxxCt8Uu26jcHHw
pyek6k0zAeUjzJtZF7Vuc4IaLZaAWnkwJ9vYHuwWs4idkbzcmu+2qpdBO8Gov7nj
T38BV0uFzJ16Av8FZTMsCjGGS9C2qV9pQgynB/kGTmu0Ho0LjW2TqKqg7Pu8JeAt
J3xonun2pgiHMI5nom7W2/DRZRCIsv+MVOY57mH8c+O3feetGCO+knXQK+V5QOwk
kNRreEqdSngXFcnfKiirAf6HiGsrzFlFAiPI7zi0oDT9u1mg2OpmPJuAMgliOnPc
g4BbuHQZ3hpLEgqxLOWV2NsY5YmuYDqoLKgIUaec99w3uqGNYNrjIOXB4ElCSReq
EvPZCcp7pX42J9mO4vTjFluu9L9SLs2f/GYVri9j8VzdVK8bGiEBQoCUWjr32KaO
VWBXXzKkyKVJPEcK7vleFRz5OsV1ikBKaPrX/mj59lO6yvFwsCwu/Kr62Nlt47Hq
yUNsB96AgMppgzr/uxvBD4TQETnue3fBXG484FJ2zxlj8iayaTodtfWd2XQOWNk3
HRV+MT/mvBGkv7StTab5qJ8IvmD9H0m8aJLQWHeopi5pkesAaXKnzc9y2sur7FGJ
MzzP50FNMA6QXpciJgC8pFlAQVPwRggU7w1UAx5jH9BJ2ROriZVhGR43ox+bHHzN
4Mo6ljYuvx+9tG1ZcnZcNL2lFovEb83GP0eJcyFya9rs5mWF1bsrUTmvFWTB1BL0
lm3sHQQaTvL53ge9RF/YAPitKIe96WjR0mnScWdeW0+Hmy5FyMqmzIsGEnVBz64A
H9SVTuI617XDC9+PR7B42NliU8g8Vvm9MPgM2f/OiaHkIc9bo2/n2oXT3RdhVKOk
PDz0N25ORfg9Xkx+xAbAXmx+ne3B3sEou+S6Db1eU7Um92gGFDEtOeZmLyeFaNNk
Y8StvmZds6naFgGjojv5MISh4jGkFUkaf4gCsEjVEiS2KzoUV4F1zvGT17vpxOPs
WRIVX81YPJUFWI73U4xHQWA6+jQWJirdNGirbb689tehv1hCPVoiKC8UnG6kcC3X
JpmR+ohX73WE0RnF8TK6qELw6A1TEZVmryj2OpNGn/WtptUe61jmPmEzIELgqmDz
OEw4xaEw5hplAzR7AAy/yUa9MJIYvVG+K7ZQb5anlu01J3hPPcn57OJnp/0SehLj
dEqWGmzpEsBoZJR96zIlZXVOmQEEedbT2G1G5qCkR5iR4Kt7Kpegmra6rxTMni+h
C4JfDxCknA6FI8P2Tqt0qL9hrhGMfZrM8RXjEiLWZfzpMNqLowF7TwLJMcjkC5gA
506yY0dKsUFVbKGrrooQ3sw6S8bNdLdcJXbkdMLbx/xcZTjzymgKxFRMqM243Kn9
EsnrH0uVvSEvG1trRQIx9zvSTJm1poSO44M5gjKfVlH1pIokPs+ifxeo/HVsfmIT
MIdLVVFXRfl1bmP2+DmEydJ6xVVV7cer0FhVIPhyw03nAnOIvE3Eqym2nDx0ijjE
GJE4iMqp6XeKEc1+pXuOWk1TOSr71QT/XO/K63R74xdZhxZyYzgUMgLJVmkqv8OF
6ARQLm0O+Td+Ac+Twol7pe1XKWqti8aT0/4RMbmfNPninYP4QKvpvkW7NfKMPeyQ
8SpXc92FsfiUkdMpahaHXVNO6IrNqCCK+AJx4DgnYhF7IhaJ4EwUFaa3TAcpMwww
DtBipI6EeTVgQrrbfr9rE6HfR/CI1yGtB9ZNxok+F3sTuHcQnSftWcy3WxxE24+3
IrBC/KSrsS06Sr18xwkscGBA5Bh0dVbnzWd3CV06v6Z540MHpC25Pr7WKHz9xqJv
xRYdQ6P1zwnXXYP2LEpbL+yw2WbB1ucLMzGfSPz6KVOJbA65PVweyBSSlcejFuvl
QKQQ/l9fFyd9PlACUW4Mjd5mIR7qedi7xJTK7q+zo63gC8NZMfiKAKmDflYrv4wk
X9590//jDIshhzi5KoASWzmsQ+uvK+iv3/5Ph4tu6addZqBR+CU3uhSj2HbrWKGw
0mD8Y2vrr1Vz4fOh0GoOA0ttV80jthStfHB7GE4l3E/Zw6De6SscQ0YUA3Mh0Otw
OTmeJJO2uoAXKhIVJXIsnXznLvBtyXiEMogXwrKB8rsXGcGRj8IWitoT71f3aJ94
HIJc3zUn5Dqy0280djl/vJOdUvUbq4Y/uOP2ScmN1FU8wY7+6R+uRbvJe5vetK7+
oCRvji61SCKHVxr1TErLqwxpPPzE35Jm3SQct2FcsKkASzJUAFQmM4+wrDYfydMF
jWv/0jC/KvfZYx3hkzHKeVrz1KPlez1NohHTxNXAOE3Nwe6CL9DELlNQsTA3+aPt
YxP0cA6mapL1+ActcvqSquqiLViD3e4MuwjkvstbjHhTFNQgyMI4bK7Szjy+CaLR
q7k/wf1TmUaHX2AE9XC6VReDmB3xDvfh2Cy/vdYZep2iIdh0Mvmb3Rx24jvsWKaS
iIbuSAUe3l38FiIfWPs3+6Dtor+5r2M1vKTJI3SKcwipiTKLZyRAwTtZiupKHCQB
C9sGAtwkripOiEwg3SAZoWIsD8rsjo8XRILg+kMxB7/X8ugnhGzHgfeq6MSmA1Lw
UsXUhQuAN/c/nkck8BGTYB+/G0nr+5g2rLN0o8dfKoHLs2GmOHlqA6rpj9ulFq3U
juj9eJ/xtoRhqHVmp+gzBoga8b6o/4IpRTcCKkbzVo8ndfC8sbYx0+bombt4KKV+
Bu6Mp6Mz064arwpe5kcyNZKJClgmMKmdLuzlIJ3qoVmAOo0ey1XyrDGuIu6vrlIc
l5aDlm1VUTnZQWbjEoga17v5vGzXk+B22wrZhOWIK65SQuSKCvAJufBrY4a75N8g
oErI73FmWw2PHUjPJQYIFPkG6VEzvNYWQWraBmTTbgLYET6s1Rq0AHQI2Pdzz9nw
4GTUO42dnUPx41918OlxJC6UEsWMI1eVuEidyckDa7AI7nyoRm0u0afQfvtm5f+v
YSm9Jv15TWTtjNunIFesw2LA/6pbcA4kXujnOGbmLj0ezVUJHNUYOG5vqCGB8E6p
UJc7nPA9hrJX5oYKudTUFoI2A+7SbEB3k+eaxBQtZAdDEIKA6WmIXfhuDWxLk51+
Shsb5A2wEonhalbVNR7HkPapePbOFSoygrh2hgY66kg06ZbiMDLaODiYoq0Vo93q
3ZBqkjZYp59P3A3zF0Qnin5Gh38Rv78xhd8lkk0goN/Kho+6WcnEOR7ypFxmmwdZ
KMQmbimoRsCtfLHaQ8wIr4YThLeaICbZGjuxi2AdNNd/WpJVmznoEp92S69Pr8wm
h+NQEPpM4PfE2QefkIJ1IGfSs1yllFF0IaBL8PNBnAkEkL0zxmi7Qxt+XuqAKfkS
swTtdTdpM2Es6h5m0VFbjJSAijfv3cDGcOvWiIdZYvOJrv2mRqJS4y43dnCIJsA+
gmIiQwzPIXp0lujfaPPRehcu7sWpS+bmSgzex8BY8+bCGC4VV1ALw/fLvFHPy4jY
XdsVIHu0M0Key4s2v9z9iengDIDhqWXEvaB2p7ZlM2JUITs3c7IsFcjWq0sWcJ4e
zi/a9LGVx3NqGwhcDbV6yZ9FFRyi4xvRQQorlznIEgpEuKEtzD/7b0mhow6cB8De
48cnGNWERL6DlVUm/GYavFkGEsuRopVtsGD9EPmHxsh3jPhamlLVCNgvkhj9XoHE
P7H658Yb6jGnUqOyxn6rkGXyqcaav4Y8E8zjF+qWm2ZmNmH+FfJz5CAAaAX08Iqm
bdTTKBLhKW52OYV9wIPDOT+LFWAwGoK4lUl3/FsTWw2ASBx4bSY4mbP9+qLl1ux9
ukhxdryzykaWSc9KaKrFiO+ZgnYC2LscYjVDocuQMsHLLG6iw/wrrSiy6hOpcdf3
jzj6CF+aZ4oDpqyhP5uS9kdNFDC916B3gJ9HU2vDPuFcQ68r1fZwosyz+BhC+yVT
xESBKohVdDeZPi6H4ffDyDjmPCvsCKKeGYLgpzxJKD2eqhJHChWOYCfN+xd8UAx0
J92qhYLKavxpfYGSI2rv2pZyEN3bQAe4dMaEXOOecEukLFzd4wFb/frH0KFa4RMa
KgEtLA5XGPA7Y+4LEzrD6BWn9w7gJZQc4Hk/fS6PYC9waUtK7AwyoqWTrwCHDj58
eAvWnEVmTiwQ20of93HxHrlfxWMCnHbUT1u9AxpJPbc5jKA8dPEvrs4Wa3NbFJiy
1PItXD/RvzbDTzd/k/X7MAzUphTQv8XJOafIujHAgCgM4KoFeJ8fYYihKi1efa0v
TEnEs2TuUF9Mi7A3/6kTiNi79LlXbCyVx0dLQ7pn3ejzvkYDwCAFC/LktqlVBLnU
xHUxDVGbuNwpmPkJrfnMAyuNhtKCEyK+PoSf/YjrTBc7dYNMdwIO/VycFENsOqh5
tUYhMCS7spRJzZm9IOM/4NckU7IlnSoEZ/Z4avYxxuoNrAkMxhjHziQ1xZFqfi0D
Af+/zb3k8JC7oMTz0CYz+nPdQDdZBkDuw3hteV1nJOkXwJaeRx6KN+NjMTbCUllX
UE/X2bzUWvXOyncRNjHMDZRCasUtaky5iIM1J0d40GqOQ+o0t4oJw9nWOQcbCIPY
w7RldL+BGgrfynB1VVAYFdfPD94k0eRFduDxUWE3tVfFmXPTCEfNfBk0/AOsfGr4
Ap+wCZry1DDmIAbs0iBQ1xhgt6IdXv8b86b/I75i1zL5g+FvLd7WoXr93iqeQAE7
qIV7pGU2bXIfrdaOT0k6WSUKbDq8a0ai+hmlFlC03vh5n7vt1u0NOCuZ/bj0CQ8Q
KeaSlEVwn0gB+UNQBSRXdfi5h+ofZzGHT4o74FoQj4fdR4hQlQUjBD2JZZA8Ohud
XaZg+m+qG40G642Ma0asNmZeEzx92li65OsAskehKxWW9idg3cIguZqhbtNfMCIR
4v8zoNfUhYSQyZ6cURufH07ftJ61N4TfEeu4pZRvzx8huqCCS7nnKB5BRhaIfOrx
Wk2xwuvI5UgtXCHxW+8iMzOe2BVxJeo/BXb5IYbIEQ4FLRM9bGVglPKjFsRHZNwH
aE/ZetFZpGbkiDAQmg7865KOYZwZS4jDWv/u+OuIYJ0PVIKWhur7QFPOt+JdDgKl
BRDG1sKrD4Kf6PB9ZGUm0OitX4zQC3qKm74S/0JBJFxbXy4lUzfmPliI7ipznSQx
qTNLm5+QaQtw2NMFpsSq0FK62DU2WAOgNWYpFVGdrcj4Fqizyn5CoTLehiVlQWKL
MyvDl6yVkdaly7dsbw1381Qj3wgUveMIzmmcoEcz5ZVrkR6sWe0gwT/3JXc402w3
DoJXC17kysiEvJPlgf+d8kPCI7xd953Wm5j2fWmAC+RwnsdfPnkKho2ERXKujWvx
oSBOmKclPoo44+MGEMyzFFcM4O7x0IWBwAyM/1EtHSC7Q0alrUScAg3X6C3fqQGQ
yp9XlAsDG4VNIZpwsmzXrcx0GkYeMXhCom9Woh7tXQSE/Ul7oK1uAJEYdaspRAoS
4dfUPRHDd+shZ6Srbk3Kd9GCp5UT+UIiL/iJmK55CCOUR92MUlIfGhtJLQLD5hCR
XyyQ8ysOYSUTaoqFcTWeDRFzEAk5GM+Ts8KX27CDZitJfR+SVvUhmg9037QVL+YX
vDZtpnBh7Ot2FRlNK7rqHD1Np9Tcf7z3+czkqk2Z1iblqCx8LcqNZQYeELcCsT3p
Vrnd4XsEq6oKhIm8XIV1FsBz9Ea/wPspwRewMS81YOHEd0955TNrf5jXunJpKq1O
4gMlzyHnpereHQOQGxnzrxpElzTTdLYVnxSjqjQpGvcfJxKI5jM0zvZINilk8A1E
W+c48z1h1zBMZkn4vjOTAKmiL/+r6Kn9v+uNLgAwL5etwb/fEVD7yk93A8GDGdQF
4FSh+Jo+u82D4lttmf9twY/zXa9nkQ0J/Rg+7hMyB3nVpdnfFhjxQMCTYdN2Uwi2
+KRQCfUDjJI5DpsJS9got81NK+nwwr/wGE83ej6v2DNme29USujq0S6ytup+74iU
l2Mquqka9kQjMFv+0gIMnHP/mKP5foyDYjFwyoNmJxgKG9G/Nq8iq2KVrKjJ2Dpc
xqm4S2HB08rx/pxXMXRPhaD9D3RMPt1VXkEhC0fwS+sCj6wXdFwi46O0xrd5wom4
k9SxzKq2sm2KJa9BIy1yLVe1ywCrPQpIA7KG7b/ixKe/EiFwaWprqsCcPb8sdqzP
4Dk5/VV2CKGoSyq7RA4o6UTllB838o+E6MP90r06khdy6Rp/WZ4j1nyCLaJGIfxB
Z5uvZo+E5mk4AAp+pzQrZL1r8/QBsh+bsI6QC7yESUh/FuGgPT7JgPYRoKLZpmaD
d2mWvufxD4zgqgloEziKQonmmQiEef6WiZE3u99ztG6yJPGOJviNiAMrybK6+eCo
UrEsT0R4qO99EHycdhu6kBDUvX3w8VJ0848eo3MsEs/pD5T4dMKgbZU18uabdW0L
aShPz8EntKo0dAf+OrWwJMZmsJx4j9q6nY6PP7bq7Q3BhCnem6RpfbAMMQ97UeVe
ezL4L8qW5nXMq1RWRa0I6aEZrOugTxYKMua0HRD8d2dTITx/oCCclH8+VoS2A+sX
4621BdVkhnAiLEYnr6CZQwQYQ2gG6CGiCNUQQYc0zAWHyxkg7fksS9dv40IFc1q1
A3V2CJyhPdLODzTv44bkXkI1QX7Uf/Ec9htZ3ktrNQ6h/kc3sVxv/v/fnala3Xiz
N3vWznu8PZjDlkgnU7Zf844r5fZVSbZKsi0kvP2tXW3oswHW1dV0RmBXJkoFB6uX
6xEYoJP8QntRyiNBQN+g+Ps8D7WgaprtT/QImJVc+YXhJwMAYOZ10RD/43WNVBIS
VjKQ//+gA8yWPFdqwhL3V2qBK2ehIPRR4GcCWSVpz8oi1AN/GVEen5fiY5n/wd/W
Y0YWmu51AJ4CwpH+3zz5B5tEgyDZYQ3j8Al0CydPuNYUlWieK7ItyPXatps90WOa
kgUhNEL0TpFvTeCpbzD6KWahr+EQkEe+xyOP7RvUszM+7cLZQVKXLUt6YTCs4cWq
iktsW6NH9Q52FR7DU79mlJsEXvsNLvqILIRk55W0LQvmTPjtSbsn1WIFjBdnZy2z
UDGMcsZ+NaT0KH2y5bDUggNCB6ip9k1jUf9g6ybYZmqQ2+E01wbAQ2KZPa7uFGlD
E37JqIb5o3j+PVoptMJ5RyguHrSgigmvGKpyKr7c+bYTvVHrNbOOY2s6P1Qz/Acq
Ihc00za5CcYg6QGKdVTMYRcWJp/8Sq+1+E38cPYZbtaWMeq16An+1UML1qN5/rzr
9M4Y/u4PJU57yua7RDYy0kWeqOlC4nlCijf2yTZSrFbo9tkEBEDCTLRC1an5q7lX
sK5mZUyRL4qLCm3E7kFGY1ysgvSnKAo3Rh8qJ5IfpA8OmEI9rJwwQOkN1cuoImFK
rWMcvHipXieIKldKSwhoM6+kxVkVT1SgF6YgpTVyovlOmg3zp4TcX07XjHcPF6s/
JHm12WBD2Bgoqp4gEkPRVXkFH8cQl1IQ7nOMlhJWtjoPsuhhR+SA/roRWlDpBmXn
K1+HppjEOOGJ+lt5jOt+6E0GgP0C2NF6vGGF6GjV29cd9HU0A7mxxZWZGMkxs6xF
WxsPrRmE5Hag1CVaS0I6PqQ31OZynYLvZUFGJbX17zQKAlroccgUKtI28vvxyys7
HVlpta1KCNpRZfXUOAEWngG72igqMV0cwMbXC5+H30rEEIIgUD7vAgSOrOpWL4cH
aCh3f7j2UFvzc/bTNH9Rgmym2rTAsCB8R3HLGzl1bvBYrAH4wkH8bKc7zcYtBkRK
4Y/uOsb800OVPiNzd+F84+CqVU5oET1d7doA4btAEnFg0hPp2AqZWQNuizByVAEC
9uY+I4BpUtdw6B4+53xsBVa6l6qMzF+ydD9bMwLJ+KOHWtz6yynEJCbUYcdxhpYo
ns8E07rKnMChJ1cIexbuqBV72nRV78YeZxDgFRfIFf4iibj0c3h/4X0FMfu4b9Qc
rNDbc0x3dnt+MhDtXO4vgpMClCHAZLy7IAnpkwW5BTzeMDCp3kHooqOsTwHKH1sD
Ivy2E2F0+pgI2cJK4HW/I59dQtwDU3lnSJ5q4J4E4693UKfBmxCRlWDETy1ukSps
Hc1bqRWmLAyEU97nDlBx4avKUgP4y8DMOF4RW07DKnLxxF2w55rdgxDcz5RxdvkN
yTWX2wPjAIIRQm1D9Wwj0IJBWwkZD8i1tul3f0iCiCPb4k3ZwV8CczDo/XeamRzN
b+jrbcpTUSM9CA188ErM9TTKDXLKj6Dv5Dt0cYXjVvKM9FugwxRjtan+s+m7b3rf
WzyKz/bM8TuM7FJtro4frdWEw/5O8gE19UZXg7rhoEX/dXXAIJ1Ig7Cd8ulaK+hs
CR8dUW0R+GQ8hu6il7iF8zPfcBrng9w2RSgsbqgRxeV3b3ekamiVIrutZHxgr10c
LzRZH+X1i56CipchE82Ku90xJB4fojjqvfoDoyj0f1shsxg3ud7jcJ0ssHR+m5Zc
UW5eC3UI84L9STcsH76Kb8hPMLDsgLgb56Gq2tA06bohlvKrXXDgujUanizQSASh
AjLbl+/buOxhHxLmlR06kq+AiS2ogBIMys2gLHDkOVfGmV2d5Q+3rUQCyiTkmyso
qnvj4AsYOiSefoEIFnH6+vA69UY9AinkgrckeFh+Vat19kGK72eKemlSEDgfmN7s
RzUMheeM7JfbfgbN3MOeGbevh+g6mnH5m1Nd5pRASp6o7QUYr8zTW1IZcX3Jxjjs
xyRwz3EkqFTNWKhb/ohRB8PsqRN7iVjguemLsa4YjCzBoriaKCQnpDabbOBjTD/y
5oodFEm9fUaNofM4BabSCrMyCvtQ2n28BeDMXNm01YMpL7LDkLMkrBtTNZBe6kII
Y8BCyW1a6UR+awD0ZGFQAgfO1Zfz5xZNEHqG2s5aMo0CtCVXhQk5DtReR6ZRpAUL
24X4v007PLDDhZhDMje5K/eiF8+E6aDi3/2KKWjkLWbf153Q/zbNFdA4DBHADRHL
dgStxwCABpXipwNZpfH1HuJnESUbyCF+k4JmhnmP59cFJekGx7TfJGtbWJ6v1iNF
DdR+wM4wOGLSHJJleiU93aalwodLZjzkZOAxF1XIzmFZuh8s97ARft/DqsGeRv3Y
72zZjBmvJxBBwVSJPagBI8wbezrJGpP+rF4w2P5VPWvfdB7yw7FFrqVz/q1dGR1t
oKXRDLIYQZlsdOAEI3thnK6oTPTBJRSJPUTuZcyHNleB12zDeEihB0/gwc10AUny
czUE/8cB5D1EPjaVVT0Qzw4CUjBhww21If/0X9h+hsaUgXTzD+fU77+SedU3Q9jl
ZsseuIw9RDJW1ZUpZYT5LYd23RoXdk4qmYUV1v9jAhqOdBn+cFrFKU8c/7juvFPt
s+gO8/TlmPdUF5Z1UlvoaAtKBKHyeW290dTziwJP7Ka9jTVCyPUGrAaM9Ywm+AMB
ypnhT6RUiWz5QHMSEQJ+QSYU30tQLKvus8OV2m8aYLWX0/EU4116nKSm8DfDRaSR
jVrkQorCI3nax8EMr6I/jWbZkxxAXQ95CqocJgsCXd+TyyUPqn/zi+mUjrzn5nkY
YgWxb0HTmqBDnYf/boU+qAKNy9YWlCkDbySYTDCIL+i/hy1ZVKMISKWbisgZsaCs
M6Dr12KwAT4zL2oXfXewy+wFqi0ur2VJ06dvNKxL0ii7ZKeduHrYP2iCCIe4d3wl
J6oYq7AzCdgXX+N1EtqwxgmZkuaycjKdicynQTWmjdAolrgfq7mLYWK8Xt7fiEnU
uk0y0zoc8JJU0f78vw0jS8VfvlYF0Aig+/DXoE2uv8urjlePuyBIhJaIbdCmw5b+
KNmb3PTViAXkSWXZrUaG4dlp4FGb/7Bl3V5SNpwtI2/k9xwqgnd2d435HYh4yDW1
dF7J+gWFyahZyUf8G+FuqVFOQ9EzY34mJ2V36ffyRk3tTyMyYMOtGNBf8vIe+AaE
4iLajtiDTIl3JQWk7XEZAcBwZS7rtjq/EhdMQpdrQclAclXdYGkSxgMdO6gvyPhN
1/VkmSqXuVI4EJHdVe81n/O8o2lxV49tL2prytBla/ItiYDZVIkQvNHOsu/1t1wp
CdKm2wqa9ulgRmdlPxJA9dvfM/8ru1SHb/bChmDgBeEUoT/vVJ1XtPXGWyCUx7VC
gVoxRROEEyyX8abmHg4U24NOdkmRvyvE9gigbwNNOn0GkS86nlzWgltVhjaWz3j8
7M4nK2RO4HHG//5BOePeOwduBSN+GLA5YppRv7nq6uZILSyyhjVGZP0MSL//nh3l
2xWPOZRPxg5GFaK8/gbKnP/FVkz2ZhhBVaxZ/zBlfkeRLPBm7FSz/ukf3+rQHd8F
B0LmudTlLuQrXr3QW+Kzc1CRGWKMiRfqQlBpCUI1I3fEEWPdhrPDkDJP75ghvkE/
oXaSONBJBNwy5TXQdUPRmX3QRAJbzLBBIefLsL4wiza7ubjjQ0pXEOlJRGD1u3aX
bxD1yPQqS3QZ++RcKHhCGdaRDuReAZc+d2BoVeL3gOAaAvvi8e/FQIneYLKBVbzO
/wyIXH9pws5zi4GfFNbphsFYUM4aLREXhbPIyg+zrSALqSxbII1WXI+h47bgUL5R
BsoS3pR7RYbW1w2pzlBBaodLrEs07GTuwEluM/zQF9qFevaHHdtWDRpz2mfmomsA
pIKc/9No3kAjzSARCc64IDTJGqQS/7HnKlW4C2uhUxXXOBrs3Cq4NYHdd0lSOgb4
AUzasLFNexzTZUPmQJkFGFt4QprEBOHfOMOpuE1NQe48cUJyFUaNqPkobRM6EdqS
DD6x7iwgZYPv40GObQT3F+BV+tlZhV+61/xM6m1w/6K+ozPRxPzvmLjqrMgi0cDv
SmIDCDtXlpUlV+6oeheBXJHh3BKTEeViq3EuLuz78eFWNIM210hRErxrTneQgLJx
eMAXW7pKEmz0ekIAoDpW3Y1k9JWBHiC1X4ECqsPctlqzH5VtWxYAJDy/qrErwMmL
AlPfylB8Dx7jK5qz73M5wn03QC3+MzZ7n99R6m9VybmVi110Xy2ta22s1iO0DyJc
sC9a1tpQdp77Bg5ax1T8nIvwBA+TVyfrXFeQ2ffq08gpCDSoRrPi5bck6GOBwX2Q
9zjiGUVMmJxXX5PWrNNR/G94dBeMVQffz+qdGni1n68i5/IqdvvPVIaF9cnWY64J
uX1DdlRHdSz0zifCuuoVQAskTdqgPTeqMVQegMU0a2ySyqlR+hHh/CARFe/+BVEG
v0zBRuJZ9VIzfXqXqfGnzk5s4l2fwz9DUYsfpv8gduepYx0q+hnEWgP5zYm8Megd
FcwxOKB5k5SPFUE4H2/nnzLQr3pNAVniNVRYaHS90GTCZwggfVkCVo7DBbdY35xT
wdOK3uPhUsAkfDtUKRQZxNUGjERe7EYfQea6VlRG8FFxb3mDKFOEN4VXwyXt6TKI
S8qscYXTJ3Ui9uwWU481LXPi1DAGBLsVf4SKSQ+CcB3uZskiUFFjD7MeMgk308yL
MwAAqLdahSU97JeUCnL0jJDzODHt4xtFSmPkwj8XkhPLwE1f71y+/zX5sN58JaPB
ub1XkQSe+HA04psXqTuY5Ib9sPvxMx0lL419FS7M/V37hUGdJxYdhqKHqEY/hXUy
EUJUAw29ZODxidTTVJb75d3gAiT0bu6YmOdcpCxOjIzr7ae5Yv9ljsCXF1vKwFy4
P8C9xQa2c9HAGlVBODdatkVLfLZ+9ISTJpsSsqV0SJy7aeD0Pa56h1h3G8iNmH/D
oNssyjn042oy+Egn/W4eSkWG4re0FaQOTuJPi6T6mNAYOJCJQSWum4OPX/aBDekz
wvcQ++ok68Lkocia94bWyhRUta0/68ampj64s/APMx1x0PhuPoV8gLtUxwPPEffY
nZOwul751Dlq5Wjg2eYmNNKu2TOc/4hw2PEdwx9ihDqVibmEV/ZjWE9kq3/p5bD3
fB2D5JONmPEhqe+HEd7paFOxsStwOrr+hHwswvXisO7MBmWqw4V80ua9sGPwsmeo
/Nq2dA4+0vg78cO7RutA0O9fKmMm4yXYBKvJtID43WLdVCsbooEc214xPa/S0/ei
KEPvkN0dwXBTBM5s8PQf7hXpipZA+wCkA2UkSj9cVy3cNgXNGe7keEzyOybHrWbS
tQ40tqsMGLJfRNkx17+gmkpZ7LTZR5BsboHbFy4/Rhq2zOTf0aI5dEtFgQkBJLZU
GYg/HcETRH9l15F1aupqtL3MqCWt7VNefg/P2v3kZDGFfOOuy1ek9grvEkCSd1lA
lLK4f7JJOk+u+EBxj5Kkymk9OSPkWeTAG+WwDY8ntXYylQQveVzNEFk/elnbueKt
gPCefFJ2EKeoXW2KSmQlF+rQS+r2aT0hPw1Xylg1couoVDWdiY5IBGZPXzcUEZs6
8tMANyDzLa4HnbkfhiMaiyxo9og1dpQlG/a4Ao6nCchae2r2PJmuQrmHlqLSCotS
GFXa6PSDOsHEdOjpFIW2TjNWfZGj04A7bwMbjPyWJQFJ9rPNrTfhnJMxIfAXPnUO
ileDF4tLWxph6v0p+ynJhSpPSjHAvkQyT+7U8n0B4XdunDIE0mJM+B8on3YbRxQn
3GYM6DOKQ+LVRj7OQjZyhLVEUnf5/wJWjXkjU6KiPYjsokaQAkmcIk9M868njUqj
mxg0XedUqUyJtzWlWRTr4nBTfAelG6oJE56AJpxJKfuyp5n18J1SdBcWrlybWbZn
UKfRUHaEgprOFh/gMQKxuF/WbGthSTHpSMk5tJ+OOcomsLBrzyCH7DA/XpemShc+
ObBzrLq85z9cWZpeqGMKH+dGGzyUU09J5xuOQkMzjbsGuoi6wNKy44UjZdOe3xiI
bfIawnbqUV66Jji0xJ8zvKJLnptYrDLsO0WVfrqNZHuL7HSq1J6/WnQTHoHMtaaW
g3A3KuOao5437L7Ct0GzpddauXzdN3NRu8A+S+yQG5JDmX7lqkl/0ExNasLai5n2
5uNWZrcwR1RQ9/PD+osT9GKXr3k88jyanuz684TqmxguviWuX/jE5/6YP0tCbHDF
dwz0hI+sVBCOIBT5qNJf0Hr0cIQaRn12hjPehoJoPnkuDfC8xcbsFeezqgAQWpWE
6yfh0nAPj87nqqZQwiDjG3/CV8012n1tFusWS1Ud2b2bLVVOCBRMtpjdmzSfV2d8
UNmfFa7PIBzeaAiy17o5P61KZlH50OF6bk/Qtt70tkvp3kxx+0jrRvg+Oj4uixwI
QeHRFmDGK33sAZnrZ8q/9OtBmM0O4FE02nRxKhwynjZeIe3+YCu9E1r1Ep/tBEgH
xqroyWgRWO4PW9pM99oq0k785lc6U8bwgnvJ1qEbXQDJxr86YidCyzTMTbRmtEPG
f8p9Gw/oCv/tESskJzORzNrSM01t9Arrt2TDeeaDhTptOLQuBnuRKPOsmrtyExIt
Cd2YMlADXTSdGlwO+I/oskb1DI9s8M+oJuplbbkk5GOjrkkRqotdzYNU339kXP8b
EI7lGYveX1iTgDXCWJITJ3oEHJyPzMF2ga1S7HQki4IBCH+YS7oU7zDNYreeN2Xa
PXlX1v+cfW9r9LNNXkhbfSmijBnukgJaNMZX08RKnWPoM1vh3ilhUDCiEHLUlQJU
GASq4OEsxy7INInzPPXTguuClPpuO79cek+xMVEAYs6uE69NSBWyy8x8+rhlL9ls
R0as1y4eN0bRD8DLP7h9xE4Lpbngb+KlhWRltKQsU7Qvb8aDobc15/xLkewPlxYJ
wnqUgJGiZird3WiVe416uGHbLQ8L2sHYcFRQH4lJwK048WYHQDH0zZkRRoI1rqU3
Qt6f8Hv3tMm2iXwmnxUDP76z0VqKCeok6rN0hXEWJZOy60JuuiOmW7yJZgDGYlCh
mKS3krD2zZn9Csa6+7IyBB0x+kVTiVq4GQQC4mZXSpAfKNpcv8evWptVl2w4R/5T
amx0IuhXTItamfhB0QN13qjna48eGl0cftYDeFtN1wOpskEc37X5fexs9i/KpUdn
pvpKx1E+sjdUNAryuA1gRZDhLIHz1XC3WKSuNMEvMULl4mjCVSmxEDGdK18rZF69
eiHNcfCeuv+L2wif4xMm+MJB89n0WptMMLEXTWii8oVjHXxXQgv0Myi5i7xpyELU
Wv4VRwoQq7tMsZ8m696c2XqPG2Dxumx3UytKF4UnzQMVCgdpHjKA0rKpVp0Qy2NV
84Zrflu4gqpVeWxdkiI6xVyWC5dWTx5HwT/ON+EO94ys3DVaaPcGT0EQQSDGOQh4
FkCb4kMgJ2aYlzZsOv0m+g2E/8mLsk1jjL5/C2Kmi+2f7B2dxBO7clLLarCr20hq
Hmq9f7g4VbgeofIDbIaEODV8jfzUj73jO0jEb3XyOOccPkf3ezfNlJZGP+E5/5Ck
8bupfo/wraWQLxT96Nw5zPC1faUA5vWcVQ/Jws16P+LOeV7dW7138fnxyrQSmHbe
py4hynjZuhOuwbZW7kP7NUsy5E6QtzMkAPISDoaYLnJcr9aGJzY6PaIxFawmWc+/
kBhKtwiRMu7fQ6pqZaf2kUbr0+kHI+Eb/bDSjECvi0+Er33slnz23TDDvd9VgWhR
5lql7Lo+ee7ATSfNsjBVTU6BzSPo1tEE+pPaMQ7tB/0xtomEH9lYwgbRhdamBMJ5
8WkcfEpIa+7dif9jSNaq7C6gmN7Pa7/aohcKpqHCp1QGugDvOOwT4tAwVoDVUcpN
IoeTva0dXbdLR3Rm1hcCMgpXH2SCTLCR1J+M//NDaPlihH2YT6dM+ILyLyOz6gg4
WwMjq/4vBubzLQIU83WQRnMhudGe1g8R1jxBpgTaCqtH4CM+v+8BUyJaakdrd9uY
Lm8Ze1iyzE2I0iVD1i/VRMIPKdiHDRu8nLkdYH9X8sotM+vPRZgGZ1pB9YGva1OW
FKAkxhZRzc5UjSF3Ajpkzk3iaJMquXf+YMA4vQFc6deDN/jRUvkhL+a/7EH+6GzG
n1I0s+62hD5WGNuXmxb8ltnyKVon8wS+HF8EL/XRND/9YuzVrf9WFlsKB811z5Bh
dOKvMSEqokaVgxoTq2j8Q2s8zUmHH/Vh7G81FJ43ialNLfIXa4T13f1kxadpJe3z
Y8g8ORI0mVrhcKskkxVrVwEaaVHLw6w8XIWZXpAW0XbIo10be7vAIhUsTbpMISus
IZvBlkmy0u/HPb+TrmhDUXUHr4MzDL+PzehXpj+OIlLEgzecIucXMrpIS5bimx/F
ZeHr2EqCB5pcvN04dtTE7FcrDGjFBJYHABMOg9Rr/K3aklz20O9FQwxjmDNzchMa
208YgZgJ9ktdrRw8dqE3xRUUbIRhrVTFa5FrNqPLmOMguJG/QcpzW3TNI6FgXW82
AjaJ/gKeymdbvd3UciidwBG9iN39ootI8bya79NL7bLzbV2o9vpKGyWuauILTw2q
1wc/2ehc+EB5RyVvbGbaEaoJFXBnM7zjQBPrMcYrrIyR6nbYsIb4p6N7ixaJ2qTi
nk8P0WGUktn3cJAOQL+1TJ+uFh+OcVqQFiUx8zgLHhuM37yq5uwJBb2qljKyaVN5
y76pT+lxoVPw6KGq+V8ndXhcybt++NAImjXXHHu5HTB9CClGHvHdde09U8JBNnHH
9Wxv7Mylyo3vKN8WCa406c3n1QwQkPrlEu3fi5cc/oYHOFo/wMIYfituYBj9hueR
65clI+NXP0wUS8rauO/6M/c2MznZRUki/H71PN2qmwXfUQiJIcmM0f3XuWL4gneB
kMaAW6Qfz5iPEjaUKokctssXHbHXnPUfbSCxbY8ZR8I5yCLYF31Fh4eshqiaz0dh
MPIySTvlCz90T6j89IAbeZheYfsRhzAGeeS4NGbooO5jN7UJuc/QCSMjTuweCQGd
EAIpDt0QsyYqTyos2vym0xuXRA4wukWn4SvcfKoGxJneB8O8eMddKK03uC5rPKTT
l48EiFYKuCKvW3jZ9sCs+CfHmXBoH3Blll5OW4m5WQ5DqBU+Aibt88Rxz0YVqLZJ
rVgA6gYDvHB/l1yKFHfnPCG/yYhiouo0imVhbWP1Pc8x37xhVzZs/HOxz5YlAowL
DJcwB3I8VrRoEaiMvbq2Sc7FZxzUCZWCRwb7Wbiqq8fx6UvkRyL02dhIifUiCFFU
jN2GmNHM8cZkPmguInmoebDC2kqWpY17+BH0AASLb+3Fs2cvaI60QfTZqC/ooMAV
JN8f71dTpnklb4ZQhUaE1yqRP6Tq3oen/KZkuB6VSE89MCuvztSmlxaFEE/GMy3m
xW6DlQsHIr1jUQmrsQ29HIMfHO0lhzgq9OileSq0Y7fhp74crnqbOyK8TycNdNLA
7RmkS5HMmrbTcFpaekEk97SsJ2OjssjF927w3J0ug+AQUqRxNbZ+n2ad6VrkjhBp
KsPlrxd508gXdou7/+c6XV4AWX2G/8kW7JHuKhRwEkUOrrz56+KdyDMvpAQbJK5u
6+UGlLvrptgvlbLR3RxCJ1EEiuampj33HN2PMUnCoID/8i7V2LhIErbct0nJvtHK
slPpc9ff2D/4VVlt0LlvlMIpa//YUG5WHh60GRXDLtR2IpuJNSmrQAFc9wWq/KLo
8mvi5ntoXef9d/cL7N0VF4MgYOZ6GIFg2ZCiF97JTt8B2akiqXRwxmLjc5LevsXB
ogk8bRedHtLUx0M9KWn+Hs1VdW5nCLt/KlqMFMrXu+Sy+sKl//2w3GrC8ABZ4m9T
PA8eD9BwV7VqOfKchevb7kciPHHH3a0AG+kqK4CMV0s8gLuofMtYQIuEGZpIPU79
TCsnMY0EXSjZBKujT6zTrKgHZVxK3m3X8KnZUxX3dL4YPLHVDt6zAKf9N/hB13Ex
rD2hWxNnGpm67MWCjn3nMTi4lL5BlNQ1BPtyhzzBana9RO1pGTe2fqoGnd1Xu7hI
q0eAzdOze8FZkegogpkMm/qG0ZNGbITaKt7+ABroNgTBXonmlF7xXCC3ss6L5dUH
L8p1dBe7DNdoaeOECjQby4gBwioq8YvOLYq3zeVE/m5Q4zDm/rxRhEPCMC5fKpBx
84e7EfZBj3GsSPkpX4P+1fqwVwn2jGs0oImz4qbjGdnn8o0MMWxj7KiWQi8/LYsI
Q8ovcTyxKyf6X83jbG4ItQ==
`pragma protect end_protected
