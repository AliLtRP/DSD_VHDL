// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
l75ahUCwJHV4fTBONsSTfetMC8boTHbvOF8qx6mmkWYi6SxwWfk1KAQU8CNYAcYb
SwMrZk9O2U7+DTKpLOSacN1saEGxf3ZA6UDVsmK0T0+FVZ0cRJZrz0wDcCWS0Leo
axtMiV32EAPH9pzPYtUoaJqe8lPMwSQPFOlUx4mqr54=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10112)
wKJMLOqacN7fjXLvDa0L3Tpk9v+iz21SoF2/DCKN1dJSavAkuJqpilxfpgC6M9mM
QrTzMf6qwt1LuZSI1YYEiYffdSoxX4gmZO9lqef2ct9mr2zB89drzWY0jlKrWgZz
CzimhYZArHd50US7d8mpipskvsd0Y8xOjC3qHJeLd2WAS5aXmbOczoIVACI3Q1MY
Up5Y7dD/IIMYdClqkCxYv73Ez+Pluy36tyXHYUQUhyGxv2hCvWeY/ZaTw9/NClyw
13tLPMHpsXxllp6qwnFXL1gC5ACJ2iqUNOxBsAI0+kmcBMCXtTrfvFMOfcwUt4Gg
/XPqsBROlH+LsWURu07IAlO9mLeM1fHae8lD8wPLqkxtV/X8Lj24DJUROQjyPk5A
zGNxKah+3VWYDJ2xV6GMnKBKAso55DiulEWhp01it/bEMBn04VQYPTA18q7UsSWU
qGaEDX1sTgozrXRsQQg3rrrAGzlCweIBSzWGcjtoAHRU1iwbzPR3M9xfIWtj5QEL
yV6l+KjdTZ2mjgYa8dTK2FUB5hACh6iMo6eHV0KopivWbRYilITP/k+FkZbRqKEZ
WRaayR/YzpTtfM2fyHXuerswgbTK34bADX0QKWJKUDT3xF0HvO4Ej1XOZaxeR5iI
IUAfb4sCoqReHQ0DMC6lOB26JtwMMIIh3mB3i7+jkpLgz4tougKHxGhyl8B8D/yI
F2usUWnL4iSvxkXhd+FOQO0lLpEO4oCgDYk637t4buIy80n5HMic4QKQB6Xcqc4Q
o3ExadADN/Mclu5ozu860mnvCX63xXy2iE0FqUmtwSjwxz9WdYi/vKreLl0YMNzo
6+uEdcu43AM+uMEyR/62jz+RpqOmCfqbfVJq7erwVKqCHAJTK2Cv3dMVwnHcvu7A
fWMjBqQYWFZnW9S+pEaP/KBiioYFNeY8JMzzhYAIjhHFIaHTbEfyqkTMVMG9+rEX
XtqKjTDwotczzPjFlLsOJTmwLSDGFiY81lyn7IW82fGyo7aUG+EM25tLPWw3n11N
LXAfGXMVdOXV2MlmcA70+08lC29nMJa6rXI9WxeI1NCE6FuEcufE4G81kQb5fqXF
k4ZMgsc473evTQA4J21/yvcxIlBTtUBbxK2v4BGGl02+wGKemVir1LJ5cBF5iKFj
bjoM+3179E7SjqIWciQoQFb1eYRkFYrpIU7CwJhlUdfWILtyZbbZ8jsrHXyoJSVM
QsTCHc7+vQmVazH8cWEoqfnDOM3/2lq1UdEM2vGbzxvxU4Ga+GclMp3mvOdrOWIf
ro4KIh7+3FDTdBtaHWD6L7xkTP1g3D8qNBv+mo0yBMBSYRrNxosop1RAuO8/JTld
+rbBQOj5NLHAZ0Uf9sgMK+/Ne4NBSSghnYcYFPD7ymgohIM5yZVRUh6qFnh14Bdu
MW4FIxLyFKbI0kkdgXC2/GjG9ALAk6HP4dEAwNv66gccqXWNGXSUoUavhcAVehnW
7Mty77kbQaYA9RgPVgG07FFUzVj2FY9xMxO0bMr/WaUM1WM84+tHIURwCYF9NUHM
z2bSUuzjHQ7FY/9phyCvkWU1AvcMW2STcubiXqQ+ttOiqHUcZQz5oBWgADCP8M2i
KI0eKvTFUcVyoPHG7y4oyRDTVMbxYCYWMqSP1n+Skvxf4cWQxLkgjr2RfyOE5LjD
HBDH2ZUO4uGV1mkPfNqWOSDh6Ruy12fQl6WTsG1jVE97Onss9DVPz2byqqoNbaqR
lMfxBrkyF2CbwjyuqswMKbbtqxTwHJ7G6sXPKIBVxC9MVm1wQuNjHUzuFuVGRTW6
yQpo2bjXzME4r8j7cJGAaeDzhpXheQ+3n+oLpzL8VM12v3F8abdjNTVORenYPSqf
nvy9JgMXfpPzK79IiqBabOsQy289GagY5mgKDpttPwnvqld+2E7h/a5QOjyO/nS6
r8527QaPykCiSCHozv0Aul6nFUu9eaj/BbxMG3/QgyvrKAl85MuIGrKA10W42MOM
sL/EH5VBUicbAYQtO7bmZ1xKwfCk9AEXiQl4KDel2dTbWy28twfowZplkB3RIYpI
i7Y42r8NqOGsYcQf12OIyZnRMUTXIS7RFWPlwlAmVsAGMLm6LuzlIaoY0b/7LWYA
oNuydOPDdtBp4eBusaBeYaerZlS2EXD2xo++9fS+c9LcJ1mNuNYHFGbxeYJGugKE
gKeuMXd62ISb1FwrfMEBc8iQhaVhtBWYOplIS493UwBoZvleHAlTA6S3I7n6dpsU
X/YhCTMU9271JHov71DWBDxaNEISHlv5yi2Fu2cuAN6pEyelAx7Z39wxLBJyr1p1
l9Z70IBhS0Cy/AEOVUTxvnGH7WZC/G2GlX8/5cZ2AVIROulU58Lk8iSDMak88i8D
xEMdLmh1u8+zxFTH3Df2DKdYsQhLgptnghRX8HpuWFgDt5QdLb2XQVMqHgOws45f
N+Tf31X64vMTlgx/0MjGzt/vBzcIX97OGnVDSlLYWZ4CZWNvp9ku697iEIsxGyUr
jjXDrpJp2d0fB7CeNX1r5oCSXJRRsEWwYDIujF27et7tVXzkkcCPr9shznf9LzZH
4QutVNDFe1NnTacAVvkq3w//MJ1C98JkVEk37Ejq/yDfMbyUTA0J9Xi/r1fl69VY
WMRMPqJj2S3mnaONUxANy2DoS+OSUQMd0ohpIeOh0inZ8uWztQ6qZStMUxYKOhNS
SY5wpp8IaAP/3OmmVQf6HWYGsKaq3ouZc6wJeFdABCISJ1jQ7qY2fWwIeR2uz16p
YneW2us7rpbivsW0xcAbfvTaGd79Y46pJrN0Fx7bPWAZ7bINW+9QCbAS1CQ8Ue1Z
hH+HxW+9kJkdKRY6ro7fJHRT8H8t0H7cBgwnAEASuOV7xzypSczDWwuI6cuFo+Eh
JoxVt8o7smvtFxF+yHF3zpmXMvMej7rc/fA5wvt/GOkp1Ks+3BVfSDThApKltOTE
vFCnzQcKcX/p5pSpoacfl8oI/Imp7OsUd8HFQXSv6SnrRdhsmBVFIN0ommmNiOfy
BfsFVHKVcezQ89TsXkfd9Hi8eu3rZu2WhBlwE9dVgUZSoj43Mv0AUfG86rqUBoc1
3G7tcTNZdT0xAhOugC1t3DQYZ7QGF8O5jazPFVTMfbs59dwcr9l1Fa6VpAPOkQik
MEnOs8c/JugDO0aJvmUSNLd0sQ+fSnkgk/jJDPCOaQ46zeggyEoZl1BOZkUoXQvg
Z2VcAcz+7BSFDVah6r+9rJfDsLNAz+RKB8FulIzfMIY50tr6Nszs/9go4EPIBZ3r
SDykGxhP2ZeFmabi+sTjrqlme9yZ9XiiKxsbZyc/+SedOsUUBQLOK9wUfM2SgR+7
gkybRoFG82Jg2Ca3zmPpnajMoLo5LaIyFf7JcOOKNGDQ6YSXnjYvsK8yTyKrHsy1
T4xG9S0S1CZyZx7vk0vCtUB8RdldIb5Gx4M2DWV6dMo7nSXS/ZBlsIZTWE/RKClP
AR8KbwaAR6oJBROK8MjRefhI9hcTrkJMepLs94tYSgKdwB4388qyJuDleG1a7zwT
cIPPyX2UYiokMbeazV/zJxtiMXEVn4OrVQuFNFpa1oYPo99Sa4YsZ81U92dWbgt2
WY1Tf+ghZ47etZfcBe4phRrP507cz7rWhh47H6woGA9f+5qyCb2QVNd7xW110U6E
pLPp5LpiqH13MBMsw1FogLqWTZE2FRuBR0IUgRrnH1JiPTMk5a5EbCpPp9hvrlYH
vpxNZEt5bIxnBtQc/nYEpyy6NIJLnisPnc4ad+uGrZy59zekslWC0DV0eAI+YgIp
kgTkZr9CBjCpmvjUKGqbyJvKGkcYUuAZMoLqK0QmWTUdmS1QOZoeQSz5NVhkEPhG
8dgs3Qjbxyouy83y80n3O3D7/Nj1rM3sjJ39PU/aB/pvRPatnJictgh1sXYXms68
KLoCIES4CHBgb3nU55ikbL6r3WLESoL5rcyEZtlPKHYbGQ3NaxpNMl76DnhGbbcl
wYDS94dVQo1LordGaNMVHs9jndHBUeqWkQQRk8lcmyB2T2jT+wKm1+eEcZ8j5zc6
V+MWfVAXaGk+SL/Kzg6S4eWrhK4+PFqcbSJ0fRoDPYklR/qQkFO7n8F1J5hWB6J4
FU7v0ukDgPRTaOC7tjBm8TiCeUv5LhAgI8PXdJUXFBf7KiB+Bk/WTFYgwK+E7itC
6XQDblqdsuchh6hmRI29yrqH5aydZFXQOLLzhB5jU1AHGkA8l0xpR9bJkOxq8nms
sbvLwTWX5lqkYRVGXsrVMZF5w+M9nP3gxy0qX8a8eAHhkser5Tj2BAK/6ui0wimm
Yr/1HjB0kBeCCk+QyhEvEKZ9FUsx9JBVf8X1QXuN61MDVP+vvj0GwpUAgKv7u/k3
uLyLkDYinYP5F6GOOs/fQKcXa26fymTJ8+y+lEeBWjDmaslBdT3wkKlPxzFqD+/T
k0QarztNVPXzUQrSJbz7NdXGZ/KtbzVxjIA3jq90e2EdeQrud/kLr2NXSolp5umB
IucqzkUAx6mCsxx9drFBBh69Yd0/mxBFY+hCPQeW5E/6umtfszKa9q6sApYqB6KA
Z4wsjBkRTDRwDTlvpBBPv3HKPmbCsJeObnIeFAXb7yWVM4WNL4o03krDuHFkpfox
qhxrc9gJHA04dGnwTpfVXN9/CHLWtwVdSFH6nqU09AXYCoxQnctGoym2gpeUMdNA
pG2mldXKyz5UyBD+zmURi3652RNRYjmSTCe0Bbhyl6DGbs79GhaOL8l3y4jjQWdy
ObXfadIScm3G2Y5Dw8zcMHnns4palH7p80XDj5R6fIR1l+rzDMlEsvSnW39uksDq
HrA/DkjvgBwIJ4043BNcH1BRpkCU1gbhEr2dRkikPu5m4OFclml+FsTllHVpVSgh
bfQ+35gVlQSqRAymGUlUHPvUopsw/3SX9APA4VAjZOe/T7fLekisKnFVe3w7oIE4
1q6rhbuUpZ9Mj+a8v0iT7VlHFpNbbqCbeUy24KVa7fBOgKK2C2BCRjXtqhCyOC+c
/ffc53mkIN5kRY1f7chLdZixPh0Dgo3DY0M5l+0A7Zhdxao7I07UF+H6ecyA332n
Ur6Xm3s4bs2k4abUykna8KWV7EIBG3WMkuPFtp5Wg1vy9g7Okwjxp+VLK8qUVFyy
ETE2OWI44MAf6ylsjhc7rBWmlEjxAOYrnN79G7ZdcjMsDKEcMBuk9vnS3Wv7Pj28
vAafnyZCnHbWr5USwAx7nDrUeuyTo0VaayhhBBUse5qNkf65QUTpuYsu034luABW
AcU9Du9bm4R5W9ZvsK1wFd+evoCilg6Z4qfAhLBRuVwsqTI0utNWVpYcHN9OBTp1
Pj31R+yVp2ormq/H7yNqjO0V+WAldg58B2xLKAfaJgEXYPtSqYuz/rLdyVCtfl7H
Q7W7EhuyItmn2VW3EnFECSkCRTQKSDZCViMosQur/lo8bS51WS/24OwPQdQmkgo4
HOOWIvBzX7eFf1bn2FhlALdypcKMqMd9ElljnMzgI0BFZCJ3cW7c8arHTvME7kCi
U95QF8pg+gy/kH4Uca1c/VgW0QIUD0VZr/uAxLZULWwq2eTpTcLSfdyhiywFm01s
QMeaVQASLsdIDt6L64LG4C5UEzsOH09P1tsKuLVYJNUw2XMS7suaP99cVvwZ+Os7
rMw1WO++1V84JQf/lXvWAWndudSiRYlwM/wdpx6JjPDQ2nuVdld9X0JpUj7x8tCw
XAEnv2f5+hwjzaEraYa4OOtbowcAayosAAvMp+MQcg5vK1MUC7zq0a+dt3FaVV/N
TZK6dxxpFkg+HmWEDKK+cjquhxPQIAE1jOl1tfu77Z9HPjrPHW173Dqy4yNxnoJf
heRXvhNcHfxskO/PhiC9RGKH0VBWZtb7tBP3YL57QgtZYupM3oM9y1dJolP0DdNE
DUo2TWowapK//Jpi4bJQc10eOAyRbddqdU51b3BAQURzUUNxZsfJ6YxZ0blQlKAG
Lsufo8ek2HKrgnRccMuoy8aES/2iUAGYOxCHmVfCDZr9dmcma+puuUdjIGYIACOc
CLkHNwWXI3jIV3rqWaKEY9QUNUYE/pFfSUJQnpHIJdDVT062+zLTLY/KxCQwMoBA
orA2PXHYX0IVyXyVU1hCYI5HcjXUZE9yHx0dGr6pZ9brvvD+BGGvw+HHCzavH5Oi
BZJF1Ybf4c7VUtbm/hURJKl8W3g6ESZqf48GrncFBH1fn7IHXuIXemxU/IwtuVNI
r6O6oGC7cJNLo4H6250UPTjBVN3XAGBffzhX9BBpMDBK5nJkr9ZV08R4TkCK3z5U
1zveEPedjRj7C/GzVkM2Rnkj80pXL2WV1WEXdNBQWSVNgWNLvFXGHaX8vrpRsIXf
ZnyJ4NLTNlsOOyWkrdOmYCrx2hlUY1OWHJyfqb1XMQcBW+WmLTFXZ+Kl58JVOA61
kzJMOJ1PTD7HLmp/k4sqgpIE7kWYZOFJRObu67G31KF4wlF+/OIEl3iRPWJMDxZu
U02pcmUbo43JcSXsKXsnYq1OiYHluK1f59QCefzbyQ6Qg8hS8fz6Afsqm7pgtUHZ
dYR6dTLecAbvEgyxdccCGrmcXDq22QRTQW3mVOy7ajtBb+Em/eiYi6bNEFgFqXVH
U4NbFThJuv7KoUbTbiVpyyk+Dck7Wka/viLTRHRpfI9/mqC4xvoP4+JzGCDSgPVm
x2F6PQf+3vEJCdZjEe1Ka96A1JpLbSQnZ0Z0s3S6nQn/2F6wNRnikDpAtVYPSrsY
d5JeDnWUA6kg9ZXlJl9tSbxH2mnjJgpxF4EA3Bo+rRwcAE5eax7LkNuzAuJNjm8T
1r/yYsd8lsd4Wl7urHgBkQZgW+y4da8+K1M9re/7GQCTZ9JCMI46PHAC6xQED0Yi
3yrB1droyCkNsSJ5YPq5YoOpCrkJjBm0RfQ8cAf1ob5YZolDJ+973y1ZGBY1YL6J
UTyktr3HYUq8sUQewz+U3qWsbxDHHGlBiujjA/ERTvTv/wMZnEgEQn6UUiHqZDMt
SKjX4U406RgMsHofgswMySovSmSVsl7GzqrfKLlWNA6WpfR/FCLFcwdJhKDP6Jld
bZZJUTRiG1Ob97u2Xv0eLZTyu/s/C5aEbq1Buuf9QqbKYN4PmB9raaqRN1fnspg3
DXjlnkiZo+W68xqP5Jl9nH4Dc7XKJHv+se8EcIAfEZUfgPCDOAowPLRBBlKj9xGo
Plrfe7s/GF3sNURWDsnoJiBJbIDilKrAWLKaBkr44b2YFsgYJiMx3iY+UDwsxMj8
mAmG2yVpWbqMq9pXlH/e4O5H8lQALkTqZpEld977BAyADsd1UQ4388Ptl1j8d+mf
/mIYaVALC2UDYr7/VewbRzzUDej366kiZXAodP8FITQPqp974oqVahr5IvpQ5va7
XqG9v+8Tu5iOvNIi65/v4+0QyKDVV8YQAUvy/+zjs3z2735+Sq2xiK9dIDHIaAvU
f2pLAtHyZznUtssxZoQa/mfWZzzop/yN3xHGt6OBYe8l6LXqfL3XmLOV7wTr1Zv0
dnK/U2NiefQfrDH+kFm6JEsAM4s6nw5R+uXkBcgXxzmlTLIRQ+IuAzyK8/D4qTqX
iLmSJ8P2/I7FlULE7rTpIye4htPHfllCuLSI6FBFJPM7ooJI4+BHKeKB1Ir06KqE
Envn9oWGHKjXsTGMUJ66KplFpFPaL+Nv2GFP2AZqi3KS/4imVZba2ISELZahJLl9
NbeKbuSXudONjM5r+88oJajYolLdyktnFQqrizfhrakVMNXG9wCnclI0t3lNiK5A
taahMz2YynyjtsszAHv49fZIGp6fQw3XSGysiNQzc3qm43VFr/9HrLEVmc+spCm8
NWrE9tIDnvHdN5eesRoWt22SzidpDev8biDfr6EbixESnRRx84FwyE723gyLHOuP
jQtbRqwe5xA+rgjXp2vxIMID1AJ1UTfTXmSigPkZoxrFJ3DZGwLLlRdpl4lN95FV
K+01YJtOuiiPpfVGhaqHKWpRUq6JyTytAgaEE+HUlow6tYel34JRdb3IGLtZy+T+
6rQfi5YI0vq04ppXkt7t6Egt+grbdons9HmwRzVnfhdhYonSCNrZFBfIUV9h9pi5
yBUoAoBVDU3U9P4qvyXEda3F4FRgGs8RWFefOBYNPSfC2OIWzmN1XNEbEAq6Z/EA
vdcgIX5Hzfr1UAGqQB7hTP6aDz4rfkffOKxFIQQKv03i7vOrHG6M9zQhdGDOUCNP
Gw12bchxhRPvBin8mROOobCKTz4uWKC/SrmOdXTePuUvy5QGb1IjhVvg5220YgIk
gx5k9nW3Z2eZ7MtBpf0XSpdDS/2721rmP623+yo+rxSKgLHTvzFj5TfmSTaa0OGG
HRReiIixcQX2AjgXJO4lLjODxlQsyeg0VLrmAfD59k+zmqRtnIdi/xeKmvf2aDEz
gnS7NbutZjPXgO2wcHGfFo9xGD1pXf0FP0txbLOV+45+ISvKv8bmWRXbDL6TXiGu
vtC6VjBfMf6ygLbNkkhQLcgxNVaD60QaHFjmreakbymVsZo/M67RrsBMIYjGkOI2
q61qVhqtSObKjP2fVh/bXoxmOENoG+fRPbQsLHXC7dlOGrxoCwrkek//KaLMFynx
eI6ovEdm5ZSyVR1p+L9l2UHbEolBXwT2mYo2D0AE8blMEKHvF8Nfny0AFAqtTni6
HUulmhAxoBcNpNN4C41M+XOYpnTKr9Y/G85ZF4DVN19PoQlqklD97SsnRakclJgz
K7G+GjuAMxMJSXF8M8pcCrR98+GuXrP8sG3KyNFnkmIrWxFxB5QDCAnemFHzUWqV
87rLSKeU34UiAmMHAYjyJgFRfiWgVYJVOSkc9o0HMIq7IOoolSU0LSSGDZws1eDZ
jW/QD22F7RSjGFhXpLjtkT+sitb4dpNNYIUBEONqH2QrEq/iutJrHkUUJCbe2ztz
5V8qCvOOAovcJh71GqoX/GRgqaq3p7iKt88XLBBRu/k8ym1B3vxw2r98J70F97fn
MhjsKXvwjHAgBBRSfvES5QcyaFlDoPQQrKTZl3jNtVrzeoFSHjBvBN+yQ7RgKfTs
qnvyZPXAXAr5CZDLNEPC7j9ru6vwKxtVPm79zbgdsW7hVckNQRkeCxmDghJ7Th2B
zROA/5UBATkgDxiEZH1N+x2+x6N/zEsuSjpDzVQuEQMyzKxeV2IwRLGjv3dltRQG
jDfQ5upCSKVH4XVKAP5/qUmSbWHyt4h5OsfaJ4zJ6DGL3Y4YB2U85ksZMba1hb+O
tourusCRsN5mdZ/fBdFEzDhKJZv0hbu1mxmA35XtrV0VKOP65g6B7CLL3bmjmHFt
76tociWBIqRAgtbpFdt5sJIP4iEWWaEQyjJXdL5M/P10hDXNjFhePjIblgWs54NT
mXoFCvZDYBYBbULNkUq/3Qy1jQ+OnIOfFh5fUGMvTe791Co7wBK1YfbU60qOou5v
ydicJ5nqu3zUOuf6kNI1anHVC1K0Av5KIrDPicjDqtp1JuWPOW1pmFJCxkx/DF45
xZ0+ipaAjdppYTKoKNAINrXeLKa0FIq9hXYSx6sCpxPtLR8SMyRa6AzS7BcI/Vvy
aBN4zVS1oOuCfNTVlRWEvaF+eIV1KH6pcX+K2Xg3jqKzjlwcVecDLBy4M5Cvp9iZ
32nshHI9oomuuzfDy/y8toskYDjzLNqoFifS2Z/FxXT1ahbcERj7Sge6k4ejdCzL
JlleVZ9M7zOtqD5ja+2hHiXuS0R3WjoXyRoY8KdbICK+AJXmepV+7gdGaHfyuGxe
Kcx5MwS/HKm7Flmurz0kgIlTgPE5J44nBoMqdK+KlTQkfV+3CTYYJxiy8qjUpVKS
2qmfGwYMxucExCyPAORVPqeHF6a8GX2DNsXbNBQssA2jr36M1vZjE3y8aBFiARty
2x7v8w0wRISySvNANh+MVE2yuTDeEtctI1SNw+4AnmPmBgQ2YtrCZ4N0rAwEi546
Qs6ymbbBH+j54KOuljikJc5tePPFpoTWdZzc9CU/PdifpZXxxqBO9iMXmGTsUzCf
I4C6t26MVXyQ542CUP8fxokkSU9a4nMq2nmzNf0UIBAHtKbf+M+ayX/YRqGZnqX+
ct39SuERyzxQjMMwkswfNhAz7Q856s88wlT1FaUCF8irWK8aj1swF+0jAfIVn/Zk
++8bu54Mz6MkZe/hBBkrZFr1uTBwKhFIqvCr6wQSMXOt0ahqq/nQ6jcPtDHjywGV
zEznnZqLJDeF1dkdS+v5loNIYlZfDe0FfGB0PxtvyA4xBcOsJ5Dsbea+ozvzqlGV
f9iORr7cFioI2e9k1Mun+9jYacma45Xv55qac/H/0YNVzoGjhmT87ku3H2elp1L0
S0vk7zL1pCBqSN7Kh+lt2lU2EkBchYG29tn86qAFZ35g4FQrHp6FhU/jS/ZupXXf
ZyQuyzShFvIkVC3NFiRnRSNNJt2BG8fa5co0LQIKsQ8q2d2ljFlfU00LaJD9STwf
/2n5losc9kpwuTF4jX402ivflj8AuiikYLgMJ7an5cjtWsPYEEG2HCi59M8an5UU
DRsWb+TtscxAHvcK7kIvrabowexo1MnJA8sJ9IykMEkNwWZFvnucKLpOI5zOVojb
0gV8bFjQFrjDA2KsrpYKqnSRWaauhSJwYsOLFcXKDfKaFfb7JAVidPQSY2N4P0av
hv992lVQqj1+Fauw6d1pqHr6/vimaO9+ezyHj9zVWfe64/65bsTXi5BxxoNDNvlx
YiUWlQVZonzHjIYWMYC58/jTqq2r0iQHKgrCY9IInr8V+Tro6asOlcmMRvX99rG9
0uSQVPj3Bjqgm9NeeFM01rx5jjiPs0BFGAeDjUw7AzeOnNd+wlg+0sZSfNKHZNJS
OJj3QODLLpD0rNwP3yqfndhlTQ0fiVIUbf//LVI/qclYkddPKYdz1wTiD2fP4KP+
Eu8fFwRby0xZLIg8HcByWii4IdI1CJT3eTn6eycwk6TWD4MJIk02fOJa83sZo1w6
h2J3QnutLI5AAkeEyqpGEjGtfGyZDZ8Fm7jDtcOCuw/9lEgKqjzF864nE2XsfVcf
BngCGYcqDrEmMb3RNyuhhV0DAr3dyyBvVXitMl9XknNqr5vBQvXObjtHejMmQJny
BSvERCMyTvWddqaLp1a/F3HKFRWsLXBZV/vuY8vCIbxV9MPa6q43kbd0llsYbf4t
Zr3Ok9fKxEXvuB6qIc+ma6RjLrKb/hFWnMXt77zVAQMqSg+Jw8viuD5pF2R6K+zE
VNmH3Jv85UyGShYeFcJenz7zg58DtcsKUfrpGc4gy5FxzMQKx2J1va+5v3Gkl3Cu
6VMP3ASooH9wdqeA875b36mAgCp1hAlUb/IP2XglnC76CphAbnwPggJL5eZ+wVeu
WgrpBCr4c9uNKj5UYQ9pdB1sCvs1W9434QzMbX+sTzjyyfJqOx2C/I0ddm1ucvAB
lBn2uU/GZHZWeHwPaAPZrNE3zfs6zeCbTH8dhCNoFU/5jUoG2Fp6uZuWcdV7j8G4
B/YE9mAn0cUnE7JJ3/6UmEfZtYjYHSX92En16g7j+DkciuD37xulxxs93DLo+b5E
UaBoAvUrjJNHW/XbsN/BoJ4Nu7exAt1LJKnAxb2bzuxXuznWcIgtYFW6UH/Vr8AZ
K9ysCXL9EaEXYVaZ2Nm38oCWgsz5T3wEWcHNW5Wvntx0SMgPQCHVwQ7clYcHUAF9
Ey7ZRUMRsCc/wdmqDcgsV51bt703OgguTTEYIdIshyTZa67uXtw6W5jfsha/RK5+
dSB0mVQEpMnILk1nr91P4z6HLSMZuIw09sMbA25bRrnOhHWZvcLsp/6yoAthACsr
u78FqZeRML4YoMUVavjdBMd1XijMInrBgWmjfyIOrl+ec8see7uxIksdmEhoU7sb
o+WbQ6kipRZqjXOF6vOXjvlLZBMsQ9LQDI8/W9cSGDm4hQc9FLKRDAr7pk2g8iui
26Y6c8/Qp9MLF713LZZ7leLet2GAEPKSDafnC+k6G8iSeJqKOlsd8Q8f7GbiXNsq
Eg19dkFoza334xL9Os10uJm3WE6292tDCHCZ8iP2ku3RIEaaU2HbEL8Su7k6XTGV
KVNnM3XIp1FtujZXhaMOgqufaMFUluxulXKIJgOGJegLbx7gy5Dh1O9C5VPk06MV
L+dAy3XCIYFsEVh4niBYgpREdGACmJot3OKDcCmAIbRT5SMaXeXlLdOCQcEiiC5s
SZgv2odHEud2PremvxRQkOral+h+WeFWtUtJTnkMHfV8X693+rk9m8q2HMtAwoVB
DBvJ+9yE7Yh0/QJ1rIR4ON/knO89K6aZ9YKt+REb79YN2fMw+4yLUWwpEFNG2S1F
MeMZiWjuTWM/L/Zc9XLucvOu+b9B4gcHGmzq4y7GPeW+iOA8UijD3B9fjwffZ3Rl
gI6XTsMRjy10IBjHTTGfO3EyIY6TFM5bkFIDwWCFF09eraLGBlsMEU7AEToJvMIb
GcF4NX7aALgCLOCAILiac4RLg4WsfOBMEGMVw5/4gkbH9hek0jbmmeAS/NNEBLCi
NepWuU01uyA9rBhfXVAtJPNlVGcdJLn7srzvHS3CUie1+m8uLLaJK3KNNRFEiA/7
R4oa+5/YRqnFQQEL7ixm/gJXjs/qULGC9QhpdiTT4rsUCoB9+VHz+nhubUaf2hfs
o+hv3T9lKSfmSfb2jCEkw0BJWXvQVtzJYqu95WBB94BGSRWqiVdvF1yuco4PNB0v
azBV2W/jYSvIIIudXPwizQVCOw+iYhOP9pGlgPgJmBMMRgkyzvESiUDi0xCnjBTC
JbvQISqXi7BF1dKxJ6aL1P8Xqb2GpCEFQwYAwkwTBM+mDIzzsH8Y+qUKluhEfgMp
TNGBhGI3SMVr+a+XuvI98WgI2moQs7p0ZXKtLVKbKNZS98ZZRwcfTE55GrPXThR/
XF6Ewinp22vJsmtgbuFUXABET2r6AhlytUEoOS2UKy0B38BOSVGzOmjM8CfL7Wcg
DiuxVMOfvGHZsMGBMLuKAfcmrk3jUjy4r8WCZ4RWFABkL+2JfKTC+ubhXVGwjbiS
USLK3T03zg4lORJsKB6/YYypNf01qHISzuWGCuux1jM6DHiVYWEcAPH0QtF0AnWB
NWIrGNl/5OjhEEml9NaK3zZsmzuAQ8QGB4X+3OlFeoSKpKwFzLhMsIpePgvnHrGJ
TZ/6eX5xANwkEA9ASlKdW8XJM9sW41MvOFcclMGc46Eb9FR7fOUke7w21LuRqiqy
YoZuNm7E5BAj0tTw5xcqSrvN4xWueTUeHA5HvwoK0tck51CEHhj41uTre46bDVyP
3dOhSEzC96s7Zlyd6uXowGP8Z5Nn4yWHN5zPKny8UDqp/auzf2wZukqSsmtgRqPF
JU2Wv33H5NFAbtTRe2axaa6YjpnB8eDnmXfZXE3E6qnyI4ptIAYEH7pPds2j9YZ8
nW+5LmdwB2XtNF1PXRydhUkqWFuMxvIwKMNj+FEmMZBg/jeZJS5Fo+5lHis3f0Wk
EEvhlStLLsdxcBQDWsozPX1Azd+YhemIYj2KD/2dZFo=
`pragma protect end_protected
