// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:00 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
M6C8yFEF/of0MWfQ89uWguYqM8Uh6jFgaLZl6vuwu7xp0LZlj0bPNtlOwjSkpC3p
SgtbfBDBezVTTVmj8pXb0wqIenAPRSemM09h7SHwUnCoeEkSwEoi8WZbxqG8K5b+
6JD+vajDQrl4j3MYWaA/Mj7tm3Tcx5mAj1xM39Bfuv8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13344)
U9KPzn3gASow4Uu/qs1Ba2jZHHbwGNr+uMcSMXqYLZrV6So00oiT7wAqz/Mk0TIL
sUiGtGPlc+AoCeCEHngqkmSRK1oPIWA7L/vM36+yu4IRiP/y1TYBgpQy42rBWhBm
+pH4wifW25N4D/QQlnaDqa7QH3OOSQORg6CYrrnvA17QwXpDSXDQt1CdoEimMmil
biHPvH+zUDnmAEjH5fESt2Dyzc4mpsINWZDVRUnhKHDTiKMFlzNSFv5QmUNl8xvA
xhAcEnlp28nlu40jyW2TvTFzLlP0HY/jjc91OcG4/2W9h/4KkRDZiBRC7W64fHar
1SJ/hURA7473YW/QHgmDB5uO6EFatzL8tS2x7Vk0sOGCVDRax3UZeo5jedHvmENB
pkfmadjYKFqmhCr/+TzUw0nd/BfZXYZ0adpaLzzN2KKfom5Z6qVqvFPwcNNIx4K7
uXzBDi+k8Zjx/HKTdZiq3EEAM3f7xGhdtqNaLLBWBI5HUQeFHA/0ppN2V+7LU7EK
nThIzNaNJd0Bgnbr2TxcyViubIcbTBpopJbE4w399FzBNMuY2mgnU7xw+wMO+aGP
RaiQELzV3XfCJ8vYaFAlVXQDGrYiwt97l+13On32FGaw31KKA6/yCr/tSL5hZV1z
T4sbeLKcg/831PT+F8Vu8Yku4RxTous9IxT+uecRaMZEQbi4pad3xpBH3CVy/XKc
2R3cOBA1PBb+pYRGF+P9iWwZnnOJoYe9yEBVwYTyeLHt4lHf9+KGA3BYCwoSTrAh
yAVChKjLNKnA0KiuItOutpL+JUtkDfK+AaENWl6Isa5fmYcLHxVo0C4XsRhF4/Cp
HzUYbx0JnDmBeFI9ZCUBf2rBt/b9KGQx2Btd/6mJfTqq2U9upQxTDVMkCuGLgQV0
1rGA0sTNucGD/1cg7gEXJsrBUlpIifyYi0+iog6hU+qSSKTAGlhp9GhEZ2752rEl
Vu0WrrpVvXtrxkPdA1HmXMl7fk72HIK/o+oyGVdCTBM+3HI3VGV4Vwzv6/zrk+f2
+O1f/dgn3QN/nSBVYTRkPANKmjWmvtLu+LCyP/i1GcFxjUYFrZt0zCa57VKt/Tv1
teZCTeD78ib9PQJXLikkMwtloV+p+O+LQ8Yiov3wY0b1q9WEQvaTNFrGjX0lXf8r
VbEWwbM0+PK+u6AwclYJCB3OXSvnBdqvZiPNIt5uNB83UiujURrKNWgZc0G5igsw
fOMN37aJZMOX9SNsSsTmoMokjLdw5Ya+8tGh8fJbXt2xtn71Opm9Mef6cA1p0d9E
Gk5KYedgCMxO7Om20MlebeXjhg2J5GNdL8KSXRJ58lTLRlD6p0BmRt/FF3xJ9hBo
pWx/IYJ3M8IutFZ8yyc0sgxySyKx8Tk4ADJogoJfb+kz4pWBPWwR144EwMUlGwZA
PyDpOaulfxQNP+7SFPS4+IGQHVs/7D6YyJWofgCOug82tBEDJ0RAnnL1X3kRXQY7
/h7FKL1vR6ybRSI+LSgEg4/vn6J62n7RhVw7e56d5mF4KUbX/9kK1D4Jm4+v6p2x
hbv6iPxXIPYLSLz7Y8dhU9JnL4rbsroHhoIkwa+CLj8vFmrj6OXv/t10ObSfQsBr
/u8ogDCasDSRz/IWXnmkQ73ftSHy+anWhT9xvnrWeFJYG8WiFYdNvHVXmn3/GxT0
miCUEYSUDp7JZ8+hH/cbTzreoAJP9qeZNsNg7C9xnmEnOqqNEAkM26SDF9ERm5Lm
n8jmvc1NF0difVYz+2dWtFjjXaF4zUPDnSsyFRSfehM3uFpPZgZ8Gw4ngfvUUx4O
wZBWz/Pj7y2ZecqIVCHqJb3fNfEElC86+mTNilMmUkN7VI3XQ7YSnu/dAv0QvddK
WeR521jWQ//B0A3dpafTmCLdSzvK75I3PNqKT9vT4VrH04SJ0Z4TlDgtaY6IossM
y4xd4orUuDCg0rMn/iz1kBaYaRKajpy8jEQZiO82a0tEoHrmG9jxp33bhp71HsRC
Z13uV26pBjxLev2CKcxaq1PRRrV9gJzZwAf5tm6MfMjLt3FbMyk7xMld4S8CKEDW
Fwa/cLfVijgXtTzIY+JYRSgUyWwc+hp8LmT4+JkJS2YuSv0kOzgOFAjl3AGwFHsV
T7Q+co5sR71zmtzP6y0QPVdFEyUBqcsnxPlBZgVTmVbzbxfjgMZp9gvnP1e7h19x
yHneY2HTYoEOIkumqOCETV7OS1rkPxcxhhYAGGWXsS3WmFMarYrwZ4AvyLsyjNox
PzvmIsyP/JQWI9wOkP6kRHuYsIshUhHhSIOq5p20Xhj/+l2jerxbaw8qyzBEUi45
TX0AmRUZ3L8f18uO/3Oz9cd1ihMGy/A1fVRGphv0tcuB3QuLR0m7naXKfVcsUrIX
6tRLZzek1v+jiORBNRHt1T+en/OWEuNOq+19DeV7D5qOM0WJ0w36nmNPlfTuZ/JN
/+gth6rxa66r+jAODh1NcT9TNqKJ8WIGNHntwsQRWWaWMKXGV0K2BcWiZU1Bz9Rq
Sxb7rx4GmxI1VEQ6DiCI9lTUUIBIxVU+gzeiClpSGrQGfNd5Gi6rP0BfLXuuh6hA
dP9yKWG8r+vBgvHBX5KyZVufFUhTTd/SqQJ4tvlc0RcW5zfXm4YYLzK0hPHrZN6B
ZTJOdFRVFfNG5LfZMo42Tgxoz9tStbvbhutQePMcLlx9pms/NtJ/kK70aO/1SeI4
NYmdDBxNH0T3TGEWet8d9jL2lEUyQRdAUn1ZoFgRonY9+aqdikRJvwaOle3Qcdyy
Bzsq1Ta+RPZpAfCaO+2SrkIXLupQBMJMR83GTLsHeihRbV1g3ynyxmggFZgs9PSF
mDYe6Xnp+Io+T03HxrnQrZXo+kBhNmq8gPMHZTfHcAbKj+CjZs+Qi7ZDINxq4aaX
g9SoC1H+AF+GxgESG9+0wEf4p9LxMPS4untluBAVAL6j3lI3hZ5iABRxcWft+9J2
Ifx/pHALmnaKHjRBql+rtAshxikZPsZ+Ez2h4bA4U1ZeiMYy966ocDRQqFjDVUnY
vYTAM8e7EwQsukVHew+H0ctvmbQwN0DEs16s5n8GIQFriUoRx88GfupPYTVY6vBy
BQmbElILuWpxn+FuW/iNlaKaEaeDByu9SYtT+OrQcUqAvlAiTPQhhCpY6iHtQhvk
8a0TsChxLGx/+ep54zZ3N6b2Ln2oij/9zUZNeK4N9QvYKdIpO39/mIuPN/G5NVkD
VOvMG6agqG++/hYQDbeK7u2aKnUuLHlVT7UN0bq9LqJBFGYo7FIYCODjJDcnIqnY
NjOYKuOKgz8XGAnfYv8SSNH5wPjUbBY3XZtwSKUefAGNS7XvFhCO+98yJihIsL04
i0F0v3R5Dg8OpOso3M9bOxTAFs9F2v0LXByUdJAxni7G9s3PlEagbvx0JQzL//ZO
rf7nW3JEiBFtH47wFN1Kn271RqoiSOcMkR7fMpU5kXukNPT9Ke1pa7NarhE6xImT
47SHwcfz+NXoThnJxww/WWvNfMS6PuPsja/47/xQ31oZimWGcoiJDrA5r9l/o2eD
r23FqU4OhsGAhhcW9OBIUfZmD7ZpS5tRB14DprkDRw8omZIkARVl+51y2Smk83Wn
OkE7grysHBxU0DZEj2mwhX9GdFHhlAEBOTRymZJsEJbmBoxC4D/QLvW6B8rQVkww
3lqM/GwQ3uuOYnDj41q0JOrkyRkQ0DVelaPMYi29ceZD8DzvMmwUFnkWaOfzwQfA
j8I6mD1w3nYpgyUkQt6tNMcaB4/eVpkdR8AtJGNCldUUBkQ/S74s4VLfWNu1gh35
FO5onjL+4AP9oQ7VXMngwRMyCFvW4fKNehuIIho8LfnTIVwa+ThiNKrA4owWbvyZ
hOaUaZCuoHb9ZwtT/D1jHuvS+g0hY+dXvpXM02Pj/DfLm+6mFcPDJqzHWBlvwQVe
vGV+jhw79zjqvSBQ0MECrQbORt/5z43km2MegfV33dZiFiQcBvvRnT0drSkQVdYh
wkAEsGrt3t8UM8uFQgUyO0/Vz6zNTQfUZZkFvBcyO14Jc59LrJX5JnxT66ydwYMJ
3HJy+bq0dBQ138vJfClzxOSi+q7WXo6p8Badf/nsJxTOBQtb+KvEXPOZXCWUBRI0
RNHwkNWf3GGPidc84aEJF3E+cMeTu4o0OwZv8lthfpPS38wcNpvCmck1O2kpjeu9
hMxsf9xuuTB91AWEDoekbUuL8KnTjWmnsQBL2FMC6rgYNQUNfyqG+sYKNPcx6Kzs
3YpjCMGQv1SGoo2mc7vfT4m3IOF9Y/BLqKENVDcrUbJgyFEEmhDa/ypJ86a3t+gN
WlAEpTBynJzkew7iidatkZH+zMD4KDLYj0n+kkUmk6/Lr2Vbl2oH/Kn4dLTuCMPu
lp7RTFXUcdyrV+LF8kZeuVy6SgE1TO8GvK57KA2muhu+x18EagizAkySZDPb+JKw
m90zxFv5Q7nSsnjjwqKtgJsI1cFYnJXUA2YH95CP53Ayd4oMz2diSSh1jBYkMKiH
r1E6YCLDky7eD0k3kJk3oQD2NpTnHMN1N7eLGy/rsizKOXNJcJsG5CTd/Y+XDCSF
F4U+uGr3NIi6mNDfOcLrMAAUihRPXqVKeTvMm9vRU6Ooseg9ITr8pX3S+EdgKo++
lZlbGqUZmnQp84290H8cuKKBEV6q6ietcVm0bnAvpXZ9h4CEMIBNWGflCTcpSpk0
nCtotMNQdWee8rY2UNVAcSCsoBQIVW2IM3lci8ryLh5NTI6aEm41oOEPdfx/wEur
R4782Zx9jxuB2kPyabr7pUIcTLFVn6R5vnAbIT8ftzL9kTgcpGk3MF74GQytil/G
tmiKREwpi+/5ozKaxOqS0OBgfGiBCdsgMnra3lc0qpSm1dNOd6hXEUq9jyYZRtEu
M16haCjgvi7OmWVDzSVHMc2PZyUCFyEcDzdx35F+mdwK+critfVs5ietzxbV5pkS
l2WI3ymDI2arJKQVz6wYodaWJxO2uJmEMVIRkKPtcJuSSIcc6HkHbB6DBCU1VN/Z
Blhqak+h90+InWKK/HJJNnzVRq8YwWD3UtUJApD59lI8YM08Hn8R12NgnETQHYg1
Fc4W3+E9M9/3GALoTlcN1SKFwgVh5FczpBummrSLOYhHqOTAuNeCPPr0DtPl/2xo
vhHkQm81AEhw1ff5gFcBt5v0uKO5WqqfKHcbjHO+XmM2Qq9BwBhyu+jYdaIrx2JR
WsfbhOxXa6uAbgWMXlxBUF76jTlRCREm0BQeXcSFpfLUA5i+5lIEqA4rpXRokox1
JABhjVu5h4p/wwQRLcXLHt2lSbMz1e4HoT63KTGGp+ItMo0+DlVdiIgY0EmHxvs4
TQE15tFcCob1FvGl36ma1qwO3LODje2xw41Uz/YvqiBKhCdjys0DYoaVmlwz/nv/
R0tK4aVfih9ggUH3METnALmpmLPhA0eDrtMXiTqT1/ClSRoD0aAceJn4FGm1mVmL
P4UFKiTNvd/UgFCnWUXyLpX3OfHBpD7oLbrHAchwTnMfdV4UL4TgllbsWiztjyQW
AU5RfoQJ4X016BLEO93AlZZSJ/3hpi9ALDruSG8CJuZqlaQ131ulERvQPDbRciyz
zsBDNLHVNhVyTqP2sJq2BirEfqfdmG0s2fdo5LuBqAfSVesfNAb0o6TLStzWr3KK
SZgKqm0JZy7A7/cXiJeYNxjl0mO80pg6MXIAufGr8VUdPGqAkoVg1aHTRj1yVOEG
qH0DsqszAZmXjQ/iBgIXxN6ijUPLBLjczzJ8dLaX5KT9zF2qz2OUAurU/pCKUB2Q
kO4flEa1dGu4lyI0zsCp4roO2JHRcpPKAsYo/jWxf1f4hCvkCXx1Zv3zBT4oXbUs
xBUM974thaXxAOt+EfkhSA5d5L8zb98YS8azKaUoC8F6ce0MV6UmIf+2QwK2mQb+
+gb/SUjohYCPkJFJSdHnYcZEXpXiYsMq4K64jdWtozsHodrKEJixoSx1ZR/3SHsY
XMvorwJxhl+fOnxvXDajOO5z7sLJuj8qcBwRESThGQRGeS1mBtzC6v2JsxW3GHCP
VDnKCEX6j5BGOp+T5M0IM05KSv5raa5fdBNKdM0QI/g01BxqmFLBk5RKindrnA62
uZ798qrh7+BlcmlotLaBsmVq06sIa4TzstmrWqfjFigT8y4lHEJcFN1EwSXIN2I3
YmcWEXY5rF4nqmSm1xezRgoEJv262XVjsbRltO4X4ieHc1fWitie3kwbgJMveDYS
R5iMwDG5izvKvhpAyrZ2wEK35rpk7pn5Z8DmTtVRSKe863bYMise56sf6SrcA6+q
tWIb+vnpY3UbLab4RuEWBsnk20HREM5FX9UAxutXGwCRUPwqjirb8k1Qc7P39xmZ
Gcco38/eAOk7ZJpDCj9nh/P10y4YakbgaKOG8MNAEP3U7cTOUYjcB4G7bfryltUY
JvG4s4UK9YOe7i+Ey54Lt+d8Ps4JkwNVDOIHQapOukdReNp5amJw61e+0KzQAisy
lS2ZmM+/b4U/Y+ytxMJH5ifTWCRkktltHq+KI4v+66T7OCcqVe1MtWnKcDNg2fpM
uE0FmRFFJh8PZgBl+ijpRtGDen93PUpeRV7xdIW/+pNZWPGywYgyH8WM7CYCLzGW
PKCp/SheN6XpNEqpmQ+oxX2ejcyt9uXHTnzMzRSzMSYwUDs+MmPgUNQrFCNhICq+
ztiwpqfmqUUDuhrKlVyfJSAiMBuKSLM8tDu6bQj/Tk4Ki3AIuONQwLt+knxUR02E
vSg0EHvomg3gTtO6zKPki+kYv9i1xYXmgQhRuJ9jz1htu/Yj9P2uh3f0Tsc3juHs
KN8l6At8gbEPV08hFTrlIcj/qaDOJODKc0sbYVL/HC7ENE6PoFj7FPF+G3qhM3tJ
E8KeCnLq/G8UgSqJRwzM9d0CMwUhK6dG60PqzBEOiaDQ1ziRX/7+JSJmg6lXTlW1
q7QrgVLS9BrZZKJzIh6aO/JXnSA0Labkrst6Bgyy9y8gBYd6kiK2YMIHCwyqhUBy
jVhZSxyUXnXJPIQl10Co5//Tgp1gl6uNkA9Uffz1G/IDYiLyVUkMgsipr6nuZh3N
K84R6CLWGc1Z+YJHzKjqOBJqhtLUD7ue7fFxToc7wkQcUSmbtixJ0mnJ7VjmqOx1
mlgeI60TfPdUc8lgQHWPszwp8sQJSnKpPalCZET24nfpl9yFVPngsdPy+ohJpvAg
Kevt8zk/Nr7857Z5qGhcvX3YHEc4Q8Hxtl+NYTfzAZuHLC+iOxAh0o5m4bik2Whf
kgUJqZMdujELejusPM1MQoREsCInRnRdievuvd3c6Yu8iRdhI77tFHWXYYM65Tiv
R3KcRrR3gMuln6gy1AdfUBGwVFP21C3CymKRKzfsLf5u13Pl7WdUIKM0kazTP1fc
9weg8saMrQ84uRCTtW5qhEpHggj70+AO0ns/D1xtuNngvgTNC/BT/bcdDeM5KMbA
bmD3i2VcbWKx1Lyxo7UV8Wqx0jNX8h/dnXV/WeQwlwref4ad+sxXaPu7jIhfDXU/
U4GDWvZObj8C9foMO702/x4I7X01XhiWYmSNF+PXKnXwIB7g2RQ6lrpwU8SG4cTD
DVvT8K0bEV1mgAbqIJevCraavRiRjV45Dmyr3sacYOm+4kGRs0ltLY0tKDI4bxv5
iHIsCXHppvMLx028wzsbfbKDndCHsXJr29++0j0azxF7au8uvdL3ZZTFUfLm6VMF
F/stIF9shK4v5PJBMZxmUhZrNK9M6ulO7txnlmE5wuPyZVTcn7YtcY8KJTaRM2i5
5SXHICg4fDidBbyrkm5Ybx6gtL2tZNwu+6o6+5DxPxDXrqxAAZ1pYoPJ9h3yHu0o
Wy/ZwYx7uRenCIejMQ3dLVwuP+aLg28q6r6gHuZVWS2gcEqu+l5m5+avL/Ogz1yA
GOcp0L4xBtVoGd+4dylt7J5mEP50DAjpTiOBvKT3palv73i0uLJrMuSlO+eThRB+
6cpbH30Rod4NUJxgepsaYsNb5w+YSUliptqdCSYWIlNqeWaO7jGgepKyNAIA3ioj
Agl+NeYJIESxrEFm5TvOLigcN1SzP4++p+LYh/AUbQPeSPm3ty37aHObkt0/1eNz
qLet57nOMvZkVPamP27/XvKbjQfyMFPCv5UY39K18/zFakQ6SgdrQLMgbBgmG/iq
I38l2xzLzf5IXkNTxpaTnonnr7OcUvHG12YmVa+H9mtNz+vyJeJCzAqY8SoLH4hU
w+T5YZTEhK3dc9D+xkEMoWebqnaLxkSgKTYumlcNWldQxd3qWXJYH7VrE6prmu40
vQxDPVmtbYBt8NW55r+MRIXjQdkXbi9q7cTps5DXBaBxKTuQRgGakiD0mI4gzuPJ
VNVb1RPOgg/99CgQWOMkn4eH02NoTv7bqMzH+XpTNDQk5R8Ver4P/WETa1xuOnSL
k4rmpEvJhP3Lb8MExGzelP/xYIrmUGSzuzFZA6FVoPfnMcLuaAqn6gwJIKs2tr9Y
XLiayWLHErqwKWDzpXbxlTmvXPa40qsrdw8nK0PY2N9dOjDK0tMACNiBUHZ1LWmk
vDG/H58cbpYbnJiu+djev3D5pX/HbMnur6rGNRIfiS1N44zg0e5fJSlhVUbPAUGB
kD7UhwdNQTT4e/YEt9pZ6UIQKJhlqgPGKz/F/XtKxrsUTIh14OQ1xiiIxnO/S/fY
gWTRVrU8e6FcdYytxuyyU+CYtKcjizZC5Ph2QK02Fewgu3DTWhqZrPr7IwoWtpxJ
h3QcP/FagxyKFIquYxq0EDn+m+vY7McYKsdpdEjTmjMQV0A2SmSJeYPyGv8NMV5M
xmZhbL2fN3wTYP24w5Xp0GNwUcS3hLei8KzoL2LakOcF3/RFkeccfasKLwDLaubM
638lDGUDp1gsBn7wIJQSGzAl6d3mFHklRHhj0QO4iaFaFINWsdzOvJFTaJ1hKocD
qqIYF62e08dfduRHzlz+zDVWpTO2J1SyLArRT6JK+ghrSzvDxwABto2JDPAZugUv
pJh0h+vETnVrlK7WBL7VrPab0WPl835193oqdjsDEJpKoSz8sbzhcnFl3PP9Hx+D
paVDIUy2izjVK/GPdFrJoqVio7HkdBDFZqo1c6i2pOiFANxAiabRzRjLm2doQslI
QXwxX0pLToh/fReSIVmUDgBA5FTZbl8iN9Wec0HadHR4yf/08Tf/c8slISXSJv41
rrbRaAA+51B+7jQMGEym0J6Z/MF/EbDQr6Et2aC5zDzlY9mrKRlFHAoLh399gNgm
lvz4YVQIWm7LPeyitU2PwLYr3SaodfmwWIQYv7Q3ci7n6WChU3kGDpagrOxUeph0
nMB6q6zgWoIcewI9Q1cbYF64Qh71bqSyAThSsOob7CVdeZILD0X8z9tS2ApNoOBT
CBDjALcafL1/nccZNean3pP1kUzaQux0lJjdfrqOfrJRomJ/WON6Z/KDjQkfQRp4
7tZuTnWJZCq4uRNM2lGmAF6LmeeKAEXZpPQd08p4484f0xGp3l5VRIwmJueGG61W
XUwOxMx1ecm07ZpN831b5HOe+yyKKhY53j7cnIwSfM/vC+kgJa4iT8+RRuCX28GH
8wfxoFWwdsQYkEUm33ec7WADKWH3NCfqB3Vye0G6P3rshf3oDYXo3f++6dN/NdnU
2PdzvwSpsp0RET4uuz5ZXQT8IOhwbGCiXkApOFYqYfJ4c3Qq8rWnRb37jtqrruLS
oJRWArTGgPMnQYMvbhLbQLDZZs9yUbkwn0HemqwfZ8IqRiPL/n7PNck6pf7zw118
EmsWpC1NO0fq1PDA531GOkcl/MXlaraksfTF4LLBowASy+5Zqn+5S0etLgViOqHJ
xdM9+cYAp8DK8vyJVcCEJLEvUmvyYVc/Hqiume7Yj7YxdOa1re4wmD39ee82HN+V
guRz/hlgqJIpcz72qBCVss9qS6l10Pa9lehWKaNAeswuOZcUkVLYrtygc9zCjPNJ
dzJR9XVNn6YPML1OhTJVpQ0KRFrXuYpApTxBukb8JJmsQX8esK+Y4Aw/txExpyos
XuhwSa5BQDF3ZN2HI9GB6NaEgEwpQ5/qB8KDjEEIDg4lESS0ITNTkPhmYWHn/NDz
73oSq2SDnqIvczkDEUTSsuNTTxNs+oWRtzzsrjNVDBad8FX1T9YOqiemQGbOl0EC
689dv27NAK/ZJkY2ibBTbIs4e7US6UkkbNMgEUPSJA+QUazDF6d55J3ztDTj2P0f
y8N4aV293KyNPJpAmoAb4jukWDijo1Y7Br4QZT7AqhlBoL3LSnmOkEmddmJ40j8j
OAb5bT05IyekXvg6E/fvedfseB7+RtQWp0zoFDBmMM4tYJ0Q5rm4QGt9E6vqN6Tb
kovO77G2JVoIRwv8j3PTQ5WNf82Vu0xS6X/gnaVN+bALpaQe07iFeHewRqzmNAIb
wszT0zp51JoEYlTOVq4tRyfTsrrCy3JXproYsgsxSPGJpOmyJSm9LJVX8mVf+b5t
hhsGcYnxeqhRvx1EoTAl1j5a0wlMypHxyheLWZCqsTmmJucVmXIZMUGXXO7ABSEf
Nfn1GEyYHOlI6sL9LwDcPgtpai3x/kWa2sNTGkb4QbKLzy+52gNSKayx0m7f/dY/
dnR+psKN98pvoDYC+5SJoyH1QiyyDvsk5wKoARL9n7yajW2CMdsMwBf3r9NqzCZi
dJ7/08gSyXv+zob1Bqql0UtZpT8kxgXrV3ZnisrkiP3Ivp0sRkxFiu1lqafcQl18
K01rLVPe0uotMBCdLEaovLWIB7F85DpzVVL29fF0YxrMXxxvklx6YA+b3Wpu4yN7
sWqSvNhcpJGnLcbSQB4316vI7EwYF+fS4ZoI0lFF6B1mdxN1GFSTu9aaCnhWiDIe
zVQFZyj1rpDQs0/rzt4f/ZurYTNPADfd4m5QvobzqXzmlhzCnomj4Aa5Ipq0+5Kt
VWN/WxuNx01tERm8ZWlBq/GNbA1l4fIpBYMoszLUSLJhqxh/C5NEjWA6PFPjpAxT
sMUkqOwSuVbuPsCrE4KrDPKd3zgc2IRLrfuzo/WN+vErNYvyML6Y7SPNbDdIRW3x
x5Mo6KxQulfxFYGKS2Kqh22uuwFnoMHWfppBpg4iDTzQNMN+wLCqpLt8cUSr2jRr
iCLCk3STblllx3D2BSzEWjX/xObEDY2CEBfky5YM2g37VtcINNM5OIxIznogUtiR
edz8afjTir+OVCPkYjjg03dFR+JJxIea1UI0gh974fSUEeU2J2dP5ijyzcu83ShC
1oWAZsecWzaV5C9pEGjCf8Q13yg8UtmyvUsgDwvx53Tp6RalGP8rIt9hcidoPpEU
0ka3Tu4YY5vBuiOcbKpZfkEbTbglVSOw/ohJHqErPhqFwcSDO3TlivqOzGlie4f2
WZ1w/chLUG7VsmLtheVBO71W0gz5Sr/7cjp9jPz02qHlhGFRWy+YiDpoL89Afe6F
6GAYIQiWCYnAzZFh0oNRHFoOZw/vcMmYPCk3LCG4jMOyQiUKaZiS2BplcfBHrsmm
l+K4ClnoS1VAiyJZrgxyS1Jhj9UtkNaMPJGmQpQYkKjrYiSon6o7Rvj9OXji1lQd
bnOekZBc/ib8GCBuBChU575SXeuVOGtwCyLdxNP7mgmo++LU5gI8u1E9FO0AREY8
14vGisz37tIWC4SWs4tlrK4YlkoK7NvphUFKoC46Hvak+Hy6sM/Z2Cnk7S253sNz
hYaXmY9sX63zQ2j+yzTHbvA6THK7zCfkkY53qIxs/zPnMaYuBQ1icS+GISn46brj
AYgtXofDgZW1H3cLKYMifDJDsZy1dW2UqXiAu8xqi74Yoy/ceXZ1KTjWL4rtvpy0
1PracLmkFiDjHbVRSgkpxE6R3T3SAu3bk8qBe1m8owYwiWUsfWJyglvWrgv6O8M1
ywzCX652E63CvPJwFXQpiJwtbbo+UpyLBdLdJ4/fPniEnvOOvNBzc5bgRcg7g4d4
xeqA80XdtWkaV7uTcIpjUxmd7oWMM+JyAoJ1srgv72S0WruIGUFj4RoPzDROJvcW
SbDGfnOrnk5mNGl7IVw1QJiEUVtbgfsA/gm8m91rmHmNrP0ba4nW4H66py1/NnA1
pn7LKVTM3xJC+JEOa03u4QeuV5lGlxb0fkyd8ywHCxwQEjr7OyFElnlwSeMdEWt5
C47ybcI7sj0aLytvCTTpzxlqAocFsS5FENxpu7tTrPL3rLKf5Rdw7XsnkP22AgQU
xFg8Hi7vdr76OTxYNy0WcSC70mvn+0VxTdbdLlolMXSmW3ozLkRcOvnF7QwgwI26
Vz2thwtDqZb/ZL4loRzPL3PfoddTA9Mc6oXc5xiEC0mS6L022/h73FM7JeJ+An7/
KfBDyf0qQhDAVzvNjti87uHuauEzhSiBaUiw0dYk3yA5Gz12lMQT2NLaT8GSAUq1
eYeZ7mV3ZAsLxNc34yFeqNYApVd5AKuUpRmS5W5rEhQBHonNNgkuJACNOJZv92JQ
nTQmjdaluefLGjn3+aYXygBUqLQjCDXQoL7Ftu2ujqzytK1Jc5NGPUBAsziF1jnO
0JwnNvUEexG26YXA/HSm5shqVn83nocg6+DRjlredaAEFR4TCXTJyQhCIFC3kp7O
3a6L46lxUn21HeqXJuigjtu1xyyKvoJcy6T0LF3LAcg1NtXOLAMiQYYs6YaebvGt
Xv79m6CNDd2+WG6rmy5DeoUrqCPvZidKvRibyxSwUM0i0k7oSBHM8y7pqNUzZd+C
URWBnWGb+oK0tjU2nHvqg+swQVbrhHti5KGqJbHvGYsxVz0MWZPqF+UoHGilAEg+
BuHT29GJ2X5OE8HBEdG/hJh5LwVIIYB9UFxp/G/Pd/G23lw3TZ88SN4EAg4coWln
SfT/23xsFy+Koaojcika39jpTUdo56qvYrl2Br6QHj4hxZlmh/ml7RQXhv8Fex16
0y6lJiNW7IvCdcM5EaJtmaRhQyKRLHrA1VMohW/qyFlBNx9to8mbgkaP+KTGlldv
jEODfFlU72yAtB3eKQ7aLybrkepmNBGWs3ncKp7+FW58x1gSdCRMCc3+uzlZ7baC
VG0yAN857Z/J62KT0zzBKN0itq9bJUWgq4F/5pbxKWX9gFOykhQkpDGIhC22yZHs
uj0KfipE2yQi6lsK3/PoW22u3mmbXuiQkgRlIWJJK5t/ATqaIcGQim6HwzShLqrQ
sdaE/EXNJgCyjDbaJfgU7qCd9gXVV+K3nE32PQGKqe3g5UFZBstkVFLkwLAg7p/I
oEfpD3E+kMWqU4jb0P23t8Q2VkPHfdnSRNBqkC07ODIKc303FJCs9ZvYxwYAYi8f
Z5vZ346CVwHOdDUmyvvfBzJWbNkBW78p60VNXvTCf9P3rQHzItcho4sTWXCBi2Ta
Ep1y43oiWidvf+5n+565rsxO3OdiZerDAHueK8D9PgamC7qqfsTE1qYpTrkVJOfV
Dr11BfdmgGFwN9WPOWes9zZ5sA/L/u8qlZlZebt3JkA2D9pipyzbQ+E+y251l90H
kh1RrMmtu7w8LmPyruCbBZEYodjGsHlY/eZG5vC6Ft70r6eWwmP2Jp/OZ82lxNPC
97pxPOlR5zFOPtnPQQKLoXocEOzslM3Oja17Umo3DnuhQ2+B/GSuR+D5HGGD8HGe
Y4sgRI9EZAFltDlt76CfTbgYginsnQL2O49UnZWN91YV4gZZFiVabWTonmskLV7p
E5SccMM3RSRkxghp49moiKG1b89ydom6WwhDdQaPHXzauyRII0lJbg7QMEjvySiM
+6i3Ay9f13leHp64HQzTC/e+FYeXPupTeWTtSDH+igVtKvU/EGPxvb6d976M0GLI
3lNwNWW5sAuizwVGQYl/mqYirHrOWznZ649T+ptBug9TO2/kMazImvpVsw8Kjf6B
1+NFyx4fifuZ8xlyc5Ej2+LfIlO57zNomXehH3dCcwwetaM7bW0RmWaT/n0ykrIm
vH/a2A78CSA+w+Z0GOetzPAAKpqLhopOk0ADDX1tp/jg6iMo4JemwWoEknhT+rKc
lYcq0H5bQLE0kY+i85g53ONOZXM+QuDZzo0QSmfooIZnQEyNvmicmXmL5rFYJe19
5GlSuIwjxM/JQQJTLdN5FFrA+gi7StODO7l3qP/EPj7k54Q6OInblpx84GXZ9whj
tiXqt7RStKp/J/OOjsG/vUdIPg56cTnLlpOkx7TGpF+uAm9+vL//Sso0l/VsKxnI
9jK0CHWqwNihAd7tve4f9AxCNK0IpqVDjnA+8IqemeltiSF8Gy//UmUaVxDDMLBQ
XYPxvND8NuWel4tt4q7f24z8v4jCpQSwRbQUEzraapLzMzAeYd7K8xZ17PW5tqx5
ogbjZBSl/IU5t/ZQIehOh28HIcieZtHAVChIoOqqrAzBJ/kwWTO5ksVJEAZOrkj+
DYdaz/VbbiCip3sqTkkBaNeZQl1fLvATtHxXi6VYTAuxSYlD6JElMsMGDEcjkz/P
Q6AA6gBsGCXOLNv09CTsYjl9nici7+rEapZkyAVXWX6V5MiTsSdvHiTUg5L9zH+S
sUaSzSSi3VyA2TNu06440aSqcBVkOO6L6UR3oDyPRBRKadGEyCE3gOfbh/cZOtqp
rWqRHKMf/bAZgl+dBtzE0Uhq2VxrFhueG92B7I76jNnKaGq7dgIomd1J2e20tdiW
0V9wCXb7UQe+Mz7hRo64tSyME7rt+AsI3aMPgQCPzPBQmSKleJe/RTGd1ZtgaHQU
+tY6npNWaJz7F9sp7oAkjcP6z+OXgdlTmW7EIdR/xG+DV302ifjpHS9XcBkLzTrh
AXda6WZ4kaND3KIeYb3cFFTCszrmKpP7tQuJFdZOi3G2u30Xctn37JcGQqvC9zGK
euYy7NwCLLhrDhqh7/UIOM+9fkz7JUYgv7d4bKoDsLsGBg9cFXj2MgXw+0vYwEgD
v2ZExCX9Rk/RZQV9xw7FyGTrZlGdxDNqxiK5+dmPI1eREeRx9anezD30uejpCeZ6
lhBWrWLDy7RGkJhAFA0mPhdftSr+YarphEbinzV81gGXkhT7Z3UtClebPZx3kxEP
HKlvM/RTE3IO8h+0+wQ57Uu7Mq3B+P6ng41ZLshJKzF2kEKk6lE9VHga9ct9DjzT
kl3IhBD3GwmY+xrndXsaHqtAzMVFq1d25xppqKGC/gXMd+RjMmhUPd3GVmTnf4av
qMJ14yVm9vRxT3HgTgsleUb+fpgmlNfucYkHwlxWdv89JAFu0iIsfgOsHy6BclAq
u2lwPeDS+qyJ5r2kGFPqnIycEqxkxrejicNEUfBWbZJ418eLHfXHdArvib5xhN9K
Me7Y6JVS276xsCT2kYhuhzyti9I6A9AuzuHjGzbI/FW5PRJppqJI7wK53bmZDcCJ
T49JxvuRnXGCbM24Zcu93o6YqSvnFP8QVIAjtcu+4nzR5qW+bhsaMqVJtltbUfrY
MD/iWJaQ6ka2quE8pE2D7XsgVpnO2q2dNNAWlOGwBUl3eNNAhNWHKo0NKc7pU0aO
oxu4qDhzlp2va13c8DLzxb7PK/cJtCXQfEao+dS7p6ifLwsZ330Dt6LdZ+WmhHBd
ATfjJQTsV8+tyixiyppOaK+Ha9Kc3UqO42B5onMEpe38W+wFAqDeG/q0SZykl0R5
f3ui5lxbnH5dsfXKzTdAbab0KoMwsrehKBe2b76Zs97ROQrXugFyJZGNcLAlRwmf
kImB8A8nJaGjNRst5RS6HzPrqhWrefeeV4yQqvlWw9bpezgNKzTPgL9tOPSHM6uS
5v985sOUiFYYvPDRNOSM4ulhrNkslXMYjaCUF8D8ClvvokIz6TnTseRude298HvO
avaQRvw25eJW1/0TSde8zLmFyQxyUEIAM4ZcU0V/liZFKo2+VmIBcM1HSTJeb0n6
T0MrQ0WSf/p3pdZkysj7se38pSklUwpxTWUGl7uaDQnIqEAIaHciyyX2GFSC3Fwy
9TwUsnxyAq34oeT/B3JXlqMHf3FGWht4S7VTo/qs4GGx03DHv5gAhc3WcwFtuJk4
0zkXJC/vyqoAMeTxxYljM1rAz68lt2guQiI6Rx2UhmIgzN06at8c3itPUlqCubgj
2fX6KUmu8PYzfbFVycU1a3EMwxaAtPHzgeEFDp7wdC/hprydiz0C4c16yAL/N3YM
o3Wje2yEMbIs2c59n4s9NPWPSFisjAOH+4Hx5rKtI6bH7sD9VyCfYGtgfxGNjVWT
AznoOKX8ujkQdoezXrPOV3FpZcJyKIDP/miMrBIlM2h93On5buRnyV/B2Df/v5Rq
YdFr3sRRHANAKTLM5zhkC0Am9/XXcCnfiN/NFbM0J1CYPK/5hacEPy3WFp6UIT/L
oJjKRkfs6hz9W8IId2/XEKOVPpYfrfiODQsdSco/76JHzG9/q7jaYJLCQ2C/yep6
P6Ovhn7X3RPFhkqld8w4QBqXPvnX02sJhq2GYxY4I1trF9HUvdzPhpdx5vT9pChA
OiNcKTUUMJHzFUG1sNWN36Y0v9lNUPHcpGYdE9WE2/CnsCcTtyNVDyqT2nMlwzWi
aRsohB4+dw3q6pTo9gVuahBMn5T8VFK1XSmNkxfJDPmyUi7OvCnWhZU5N1fFX/5R
77RP7QeLM3LDykDXwhs9UFhQpWgLHl2IdsxuAcuXmsb4RJCtYGU0iR8f06Bmh+Uv
g5puh1KbwX7OWXhRBaGbs5E98RkuaycCNOV2ckwS8ro6OpZ6BXYbJLxlvatL1pqP
QRFuLVxonIDxp8ETN0TDX8eJufhRrKuDs2BERm3935Z8Qz1KrJbk6rc/eZ0QeJOK
Y19hZoT4BOfow/RKcUcDBbsNphfE+y19z3afgPTVa0UR8WV3pmKD4ikWq4dCJ9Lo
nvoe2fcbxY5fe6Vwpcm+rikAGtTV6MPVszXzBglNATax9b34SJaw5YO6d1POUbDC
G8CTTH5wu5JKCmf5VFMXVfjmti5bjgkcLEigo0JAuA+2qkRBfj8DcaEl5V6WmRhE
vG2xMBZFwZi+NmiTr7I8BqPUwwhFmUmxJ1Hyctby53CleMPrFmX74VIcMBvnWH+F
YfMOuuTk7vO0dgcSvnleVt7YsAM2X8ACwFI4lu0VT0bFIxcI0qYOM5ISrf5wqDwG
ZkETXiJsKD/m3vkK7HYr1MoOxdAyZcQVqHwsdJFumoM1jp5jT3tBnruMzpyTvhAk
AH0Zet/p0Rf+R+87cRxTXoRQ3V/0fIKMVuE6AD9Dio/YCy43ywIE8evW7Xea0Ia+
8T3KUGiXCifK/mq6laQd+qXOn8c0GfgfyQZ4y0hTGLcWl8gX2IbUli2hc8In001g
9kI2rOxVtkMloLoh7poWKc6b/Lp8OMk3uamRH+RsC/HgvQKbtxJB9VfV7iQPNjvB
CSmsvqcLsw0owy1+Z6HHBeUhxoHYtIC9/lt1DNi/ai5wR/4QvqRc18h3MO78a5Hv
MBFt4TrzPYb0NVStB4FndQidJr+s8RGPxpHBcWk36gLzcjwZfWgd3BH2BNz5bUUA
oNnt5/M3Q6oimrvsQxD9pGa1iUve9Ea34mF+Fj9eSwVC44OXjxv/T40EHjlq1tGi
qsRDKWUqRpZDcMg9kc+kzS+xpExkx/tRPOOgYc0FlIzHpIZ1fqJKqYLSn9VnE0o6
P9l0YWwcdrFoIpj0cevnFoncrFYl30YPeUjEQX8f6fGtwIQM9rndEqqZXBLMfKxL
lWIiTrprpUQObhLfrmNUBW3HftFi75sbX3+8rNnQ0FpFizyk+HitnMvn9h/CG4eR
hKmmVUsZ3Y4cucvAhHVQPta7I0cOjdCi9G88Cwe0ic1S/g+RHMNBbCql1DbjkJhP
N2IfEQ7RArLgEn3NHMdzcfnjawQKliFYZLSqViFJcooh6B9vi5j/NGfmxOgmdc/Y
`pragma protect end_protected
