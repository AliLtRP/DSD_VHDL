// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:03 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AozHxQEQh1l2tiMawKCPVyOni3aE8trnDbBg5uWaBu9IpoYXh7+5v2FR2bsJ2qJm
9QFg1IGgPgiJ7Wv9eqZYql+iSeOy/pb3DkQYveXcREc740UojvQR5SEzKtW86UPq
hRIE+dsAEaWxPPJL1E2jzByGrHlpR6dmkmSl3TO49oM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6960)
CLU/OXTSCB/vKateL+Pfuiwa3gprIaTUCK5qYVyQMgk8G6YFkOlgQUTtXP1WpelV
1EiY9l8cKuCAuSbPMLDu7DeEc+SM96qUBmPwx9WaKVMnDPQbEadobh5n0E2tFjJR
/DYguNA4LwH97A7QhKlBP5GBjz0nkBA0Q6MHjJxNVbO4wLQ/+AfOu16BK8J4hrF6
Vf/ta1LWao6iWRX4B2CyuQFVy7ne4EhrITkUplw3xy6n6BWeostPV2iAI/VCVK/0
YuMfAkuD1KDXf+FHSspMQaegAhEIw6igDxRo4fRZSrmZlXsShj8VqmWH44fyIcP4
DfX1NAwYXJAoBuRXLtLp0VmiLfr1KLyNwsT8V/2xI9XBe02dkMDyIvc/GUf78BTd
4cwMuPO0vXsTlActVOBL3heaOo4/pLzohsJwH9F1IQAvFnPGjtncQmkyhgk/T9xv
Uf67P0HazjGqLifX68IByzo5oArFHR4dNlSMGbjWYYQ80QVgMp3GlO9ICcD5e/LF
1pxLOmAx5RKNKAoZtiurFlGIE07hxV7skZZRsFxTHp0/eSPJ9b1QmcPQsSH8M4ap
ebz1RTebczmpEEYOvlDxyBNI9mipT6O8PdlRePLq7z7faO2sGiQKj5YH5MrCqgjg
OULlrsEG+1fGckl5lV1rbx6LegHVYb4BijnH9tttU7dK4lH5cPMYEYn6aN2ktTk7
gxt5GyZfmaHqSCC/U4w+oww8+gbaMTmlRMR/spOKcH/7WgyW9gSTLSsXj4lEVe/9
UcnamQOViH1I/ne0depQ/ewatl5+puZoOxqr6hDEeT/aJbSjyhH63NIkJWHvMA75
atRNHwusaZUcOrsRDZg4HV+y64xrdWjE0Lyl1z0hPZTfxMaLoTuNiOk+3QrbqSCA
Zpb7Uzwa0+dFuqRSAM2nEy623ylcJWJORBWXyj2FsnKjS21lbxRHjGPKs0gq6UfS
LqhSc6Eco7BincvWqZoy1AAqvsQ2qiJFrtq2vb1Yym+6NBgOmWiW7q6Td6ruSkIq
fpRqW10WYy9Y7pv+rhv3MJaHfSvIRNgTnEuW4FFgqsiviCIcir6qhgImoiekKqPm
vRodAfG07x361vZJfONAMvu0pm6AUIgIySWgi+yaSbLkdstZ3FMbT/2bMa5Y0eFl
DYEp2erU1CO8g92lknf8OM6Ww1tWSsIfSVcHqi0RjjSDkre1riEsfwH/4++f7jb6
8LHeQSgrLI1OWvmkQLNP3cSltuZ+Of2wZgy5ToFCn2LQNfYBfg+tVWG3bXK+7rYg
FAcnKJ8LnBUvRbkmb1LjSdih1LxfYTl38AWhu38m+ijNpHvLhJtZsnj13VU4Z4eP
spCsVSz3Y/8P10S10krx7PBcFLNU9DzEYLX6wae5rzgN+HUkbuNKCInCoSTKQPMX
DqEsFfh/8LGgim3+hscPBKPmhn2RUZIYtwk5QUc41xFNywbARiRVQRJZ7cUMbQF6
pOpQvrcpXVv4rLbcPc9HyeEXEoMW6HuSbdH6XS8VTPActNU3TeNP/tFzqjKah3R7
B/Bz1yMWVud63SICMAbniEbJIex1G9kjDqjxoNJfCOJASobKciinYsudcmMvgUHM
UiAbvQpYmNA3R8XbK4FPqtFP5ARMgP/YpUV/5SJT/ZuHbmxIWpImVKik6Mpo6CW3
5dE0s9P+ys5NycHm8ikUKm/01joEkMb6u61oVUAhBib6zMDZbDQfLZ+htnuggqZU
z1js1/hp6EPod0p8FnXdmpcJx8jR86CPSxOvfQLZHGt5EoSt1DS1wZUgU4FlLGy7
fDdL0wEmSnJxr3UZnhoGzsFNYGePgrSnzKs9YMifBE/sFM46M2Qi20TxToq7ieaV
WP3FTNe6oTAeMalsIHULPhWW6EKv4mnkg0muV1oVOHP05y89ESi7f4GLpSyCtBuw
DB4Nrs/++HaxzDSvs+4LHjMx1cVYiUSA0whoqRkHtQNQdkXBzBb34GEscGytkxe+
e6PVD/NJbuzYW94v8m1JMb770KxO0pVpgvgQnLuXCpgB/Y9sJTc2YvLWVPDUwEnX
UhBxpELJ5O6uuBJ6/+1x/v2+I3gVk8aXQ0TrcGOcij9XA4CFPH4oXE91BGyuBHAk
w3iR4QddRe5xCgUpKjkV92err/NWumFQ+qwTICLWMOoClcwG63XJC13m/HU2HAuN
wO5IvCPj6Vc14ITe7ASEfsgwPy969pCpl4PyNB6xRLwLBuBmGPTAZeaF2ICpBmMa
lQMv95NSCetBhLUUJST2mo66w9hgWLYpDbFvaZbn7PEMe+yRwtY/iSg0BWsdvzxK
AvlfThouQpr1/0FOCZ0uXT4hbyYkAh/9Qpd073gtFIkbFz4rNhNkKi3aIUrJ9Z50
0MrYnYP6ScVAg18qm3dXXcJVRSwghg/KJCSYWJe6btrSGfS/n4EcBq9m/vuAF4Zn
IpN+Jz3vYflxBrtdqjxEt5OwvTNDda/AUmPzFeR0mW4ggZRLPbFnlUFRTd/gWriz
X0Obov3dNERzU2XBYI7+EXebj0SoJCrDAoizbpIZuaef/YNrPXj5wP1Vavo8jFz/
xHM85HV2U7mkpatOp5jqW1RIoEOJwDoZAz4Xgk/1v5/c5Plr3NFs9MUWcgOuaAhB
lFDYbNCooVfADj1xBaTmp9wONrjVJb9yRvXb05c0ShqjDGCh4Gf+eeTSvz1XwkEF
zb1Z14eOpwKLHlk1X2ImjSNhPqrz8u0jpeo1K7L+Ff7AMDLle5skO1SzdCvGsqeS
xfXA39cL7IvIO+1l9ydMo5EjU/QY3zLnvHA8VmheaudBQ2LatOByuK90CQIHN3qu
G5jkRwQMt6I86RszJkG15IlajPLIgLxb4INBezqy5N1ovh0ubtx3+l7DZ7dydr7g
zS3dmOLZFIcHMjDQu9NMvnTiE7P5jDtmw5lgQTBlQlpgjjz3jhNYEFcEXLospgwr
Dd+mtQBpW6jC5cgRZs3ybKLPxG7Ka23OAdilghWll1NhAp8JPrID7qt2ndNFIJoG
l73fIRK7taeH9KUsrIdGa9ktG9svKTr+Y1+VJ5pk/f4qtmMkPBtHjrIo4ck1ndka
bDxa9RTwGRFcKfZWwYVuETpl4NPoRx4yFUPBi5P+e39c+JvhpoN176yiba9Nldlq
zHfD9elZbdEItVBmd4J1RtDshLxeYM/mT+YCYIQ2eWrhtkfuAiM/Mf3BdfmwBghy
sB8LVJkqZEAyxzB6/70E0Ww/2N0wESE378izBz6nR8BAsW3CmWrBYwNWliVLXRLJ
nuXc5/EGC2L94h2o48q3d6eLF3kkp++6xgFWAta6/0OjzbFF+614CJPscNzI+uzk
xwHflTpOnB/lwsUXRBQblU9YwvbRjF+USpX7W0KEjyF04NHKnp7O+BHZsB6/9Izf
ilDrqgqDxe/jQXViqIIQynmNqgbodS/1FyveOA1m8NwypuNZ5SijBBRQ0/9HrAmd
uF5c3eJrqKd3WemUl2Qpv8Wv0ZXmyKoRZcaai1Zkw1QCg0wbcm24jRLQE9v0/0QQ
JygtyVosVTnL0kWErwFflBDxEAiprrAFbtd9REqk6nCwlHgGmSTXwsBwoLiARttf
dcp7xvvPJGZiimG9C+1doob0Ii5BP3bbNl9o0CoZ1viEM2x3WozmIi9KUeq4r5dY
7320jLKA9qHxJN67KNbXhnv14v9cnl/t/yo6uxYRdgQg3wgfx1T4i/oSW/zbzuOM
4P5aAWoXoS1Gw9UINSN2SU4yLvj+TRYLK5P0xNqW0Qotub1b5eQJS0LoSTHYBO7t
0fqQnwQY4dabJ4YyEU3wVBrDVsnCZcnK8j8Xbc9IdguXiVJZBaMcAG25qUb4VQKC
K7c9D6b3t8LJ+vManxA7tOgFlOisjD2tJTHddXkAbXmu9Z9flQVvzZRr1Y4iN2UC
ilLdfw6EDpBhXB1+2G4AmL16JogWE4o0ShPx/X0aKYioJ/fFiRq/wT1lAKt662Uw
sdpzcF3zH//mjoW3y0b8IvyvY3actHqkZYJaCzAhNUOtM8BAZkeXze18JOHgc01C
y2gWVqO+z6vs+ZI2+ijOrUoasK+5jxKP9lkwfPOuExLp0+FM85IRgmlve0YzNaM6
COxeS/OIA2/lyyjpL2oNYpuNFPSMSJROYrV0ExuEPw+TL1zyUYsTJY6c1kzQdifG
/Wvneo/vTFBMCUchHyy4UC4GzaCOzOwP9Wm8muVfeTswaNYlYXJLAo0B4KIpSeji
uEFWrSWpZOutD5VJx9ZS4hxDccgwv63H+mcfsMC8YiTM3HQJVISNnGUdK2CooaYs
bZAeYcUrHttUyOTfN28zhdZUxTrlzHE7XP5yRs9UmFGImAD38jJ9y0SwMX9UMnu5
mG5pY7oTXQctb3Rgfx6DRhXMcXx3sfhxcJhHhl3VESitJg4O7K6cyQ3ZE09tPUzE
A2nNKUVC2TtzwH2b35+GOwc4kgnCStF9Rud8e55C5N0l3Z6h6tX0RYUyGGdX5v9k
padCpTMCb2S6tj+rI+0GR6G314yYmmqgz+GncxkTJrd2k0FVdHw9J5Sry4W0yz/B
rr0NQbUtk6RW4FIKvwJOMLqeW6FaCeogXxMVkfIzPGBmBMG3Ftp2C/DEGobr3ga8
x5+Im8flappcf8F7cmhuQUiPJauFTHucqVosFmofEOJKWYddvP20FMgXu9lC69QH
XkYK6rrWAtFiCT5zrqrV9GhkKKa6k4YwC+zSSUOQF5aM0n5e1nbTfn+p0uQPUQ9g
G297XTYldgstUMRurm6kX8ncJzUsIuYWOt65ThBRxlFTqtOYMlNy6NcfGiaarKEm
PvwWSDaW8X0+lZvvIXEfMeN7u4HGUqUv0t/0jU2TkjV5zx2F+fthFX806h9CyyBR
sHod+TPZYWNpR3jHOZG5x8CVz7mvmZIMzcz9wTjCejgLzcHuddFy4CwHdyk2eDGF
PRtO3QIjWN3X8eBSSjcsxJfCTr6wIU0nqH8v/AvVanEEt3FFYmm/h1TEnZT6GWyL
h1YfrGh3RsXuojGs5EerkAPIT2x/xNFF0EeAZDkeHA+VMLYlCKIg1HcDsPfJ503V
IP0zFJZJ/YByJPLMBqZ2nVWMNxesl6Phb3U0782F+uf6VRoJfzu4xIGJmPqSWGwX
/oHBt3pCb0bxnRItidiA0IKhFnSHhdQCyuCHzsVbsU+JTcBeCRSpDbIkd8r7tRG9
XF6fEo8YYcfywm+lKuEMIEtnNKfz86UUSQFr500iCloij0WzaP2apmKczEBrkS6L
w+HwcYfZI7BQ4eStGxIuUXIRjuRXGsYlJZqizS7Zm1aF7uYm8wY7iTRD/DHcjQvi
cSxQ07lSN6Ya6nCiVd/BDE1Ovh21a9VwmVOzm/0j39T/GkyEu0ahO+F1nxTclzfG
ouN34JH/ZfTbG9zdCK1yd6JhK9eyluTN/9ppxmxFHgjXaZhKwVVuT7KSCZGY5f9g
qVa22+eW1/zDbhA/R7gE7W1VnCy3aQuYjxtsfMlUczfNUsxEHUfjM9jqsc/zor9g
eCvVpQlSm8C4mK39/NiRtyoTn3xS/6Be4CFijYRy5wjAv0R3LyVfcJE9/Gdy7n75
IwofjNmt6O3HuYXOx6gNfu7LZIFzFX+fN2A+//4MChZz8JyvYxQzkKUh2DRCEfYM
tRx2ZbQDWEeGR8eWhEGvTd6o/nDQLrJn7SioxeJEcFNUNkfyBTKkQsRW/cxUC6tR
gfWuC4iuI79cHgDvc6GW0hV2OgwqyDbcQCTdzidIANt/eTxh9lU9J5728gdRGEdO
hNPTpPbkgyOTBgRlEaIHxoT2h4jzIYoQkeqYLlA40cBg8FR6XNvUeEQv3H90OGuD
cHiGS0apq16Sml+7Kcc+B4Og2uy8ypiCwZFrzicVgw0wJ2U7rSiMnxUn/Byys0iK
Vgyis7B/qUbC9FON0/G8X4WctUpEkeSpOgRwIHGhilTx6YsUj8GpckG+dYjG+3l4
xnZNaWr4IYzxFifH+CCG3fOqmOVALEpbfdvUzYak3wcNkpeXIGE7sx6YT49z9XAe
EhELNj0Ko5EBmHdt6NBv1073cun9D3P67nzNdkjsJ9qkpQpxipWmrLaqIEKjUbGg
89mwDloIJHKOSQTcPTCPOCvQBVVw5V3vQpnPgC62B9NuXAEY4/PYXRyk9YkwRJdt
/7FFgXzWL5hy2pVQ0G0EM+bslFIYHsPcmeB6n/2YMzWfjR56n+yyWlMsL/DfyrsQ
6y636eGbT/att+rua8xXZf5kQ17NLRCyqI+wvZO0GlYer2jJ+EG7cm5ttwQfdWHJ
k3rxf28LdhHUoXQ78TbKiv/yOvec1AxltXmDNm/62KW68fU6sy1QQV8tsaNYWI15
ub5/20Obg0TCl8WUYpgiBQFtUwPP1an3uQZn4jm7z1Ck+CPSJq8hDu1j5h7Jvh3c
r1iE36oSIZ6bcGr7dl6h3SBxUY+pQlWP7MHN9Y0WJwj2jdSVW26psfzolhjfarYx
C4okXyfEqsIZKxCQy0mZRqmuNMvw2xcn0jN1WpW+qGMR0J4HMujA83uTbhVaSJSk
TEn9vQuZpUVbDMntfT+NGl759cQt0tqYSzY4I0a/WCBFFU58j88uTxpAc5TdH++/
t+E9akprpiCvQXBjY7vzMbAY0l1hNDBWsbGSReoLPYfhy5HOgi0q2nd9CFEUAk53
pS0PsRfN4TR7jBGOP2WCcWpTYhyEj+/t36Pg1QPAB1OfZa1yVVGpV+KgB92/Vofi
9ZemYQHYgeimAk7Dj521GnbDdwnoEqVPeiUIbYAcDx5qClNq7HSAwK2QSrWE+RzM
eFC948kEO2WtUfLHmOTvnNweQNzUwtZC2iG9kJqU3JoamdWKLVCXQfdZLge6Xy3Y
MgkI9S9Fspkte0pcqIjpkJph0vFoNA0I3h6LYAPm4ab8jqUHp8Ce59VGfe9yk7hb
qat3y4mkzexKU9Su3kSxIsZk3f8yZjDyvKOkvSRa6jWZIhhfIkqnzNbh3OzfcWNF
3Er4+KUlMg3tgXuHUkEgbIfsOK27bwhoSHspoWY4NqIAmiWS6TfGEGIILDyhxUyi
21H/uGC1Kb8+jWhZ1Ztdbf/+HWk61cz5KL++JcwazC9s8jLveWumXXqLiOHvyif6
JwDfpIn2cjMlFFr+4zxVTECHFUf/hgn1GErtJ+Sc+SaK2ZITxoEldttzy2egscn5
I3E6D9uUjBNev1Hpdaa7T1d9h2TOnQr044s4EteqZDMQ6d9Yjy7rgP5emvYDS2q8
oZgnFdJ3SVIvSUzP1gutVcDxxty+droQwKQUU7y7oid6+Y2GmpdpeEH+fIdSFNMq
1XLV/whkKiepfT+hW2nkfdrSmIHBA7IxyPhQy/bY88rrXQ8NMyaZF5oj3G1xOwY7
yj5KFe/e8PH45jAg1BNueOp4bGWpps3vax93BrrtlNR0GoYJJnA4/kTpbdO0IN6W
JxxCIJF7e2K/lRJA4w915YyKhfpsx8NEkUTDiArF4JBEYFOqDdyMlZr1oP5+05nV
dXnhIDgA3D2UOg6QsJpDAVtO9Wp1WHwcKOH6H2MuXkx0JVhGhcRchSrW4sxlaLf9
+SRGpaZQ3fQLg3AzGWcGrK0AlqL+F+0Bq6w3ixmTit3KBDSgkPUq39p92L7LcPHr
EmwiR5QjrVDpLjdpgOp9LAdGkJFc9mVIcWjNSCWXeEI/R8U9PBz140uUy3CkXKvK
QYrJYy+N6+Eajicchcvsw+LiCdTy6oEo994HRL4MUi3EZdtE2QI1toFT8w01KiaF
QSvB8AX8kOexcR8D8O5wHXnitW3RarMeWPi7BwmZls0nEIoTQ02ZfFJe60BtHoX6
wLpSd7osgFss0Vbptnn+6/g/t1u4RYw84KsDUuSmfmczFZM8p64vyXUu30o7hQeP
fRRZWEO+YQ4NZHlWgBOiC/qyP5e8WC6RPYxI4K2JhWbVuxm2ObiK4VstfjCDghEG
j4EaQTw8a0mGSnWHMjsOZqb6tJkNOtaad8T63tnoYGPJk5FXl72ZMPqo2gzZ73RI
NXsmHvjqu0UO/7MkTG9pwqZN8vNrQkAdstu3c2VR9+KZWQy/pcGIgyD8Q86ky7hn
V3wVN2TI+kAwOzzY4PpczRz5a+SUxQ9DFwDHafC6m4ljnZwCFDBnDLndd38dgoF7
6+kRaxACDOaHwBOoPv+AVeRvOXF4Qk+Tpu3X7gl76jd4dHSnyC9F6l7iAqVv9Bx7
6oq8TuKZloUbegLp34JVOvNlUdhI5wEWtFx4L6Wtd7dUxEtkz6NyGKNJpRVaf96V
8+mQP3GVRIifpu7kM3hUYtEbnhE3+6e1X0tKL3XXpWVx9c5cE3pmgCL+F2fflM/B
nOebsDhqQ3MN9OSK1GVWiJ89HocBS2rH9CPMQLU9JQLUKPdUTZ2LJgWk3/zsaGha
qWE2/bvv+rPzUkCMf3HPS0mjgGB2nWDXEFv1Mix9lToRqbamVuxlBojrS5mPGCou
aF+GkX8Lsabds6Wy7W0P4rIM6AP9YbKybroFrj/xAHpefGmK9p9Fs5ZcqXlMS6+3
IL2A8iW93nYYgNQCa8F2BAOUBD6L74WnwVwQWz/T9JYXbwX/+O3UiIfBhtR8SU48
nz75mtfLyw1qbuqY0R2xLu5vfbg5kRFQIdf6RTr34zLVDBCmlMWczs52Mefl0jLM
30NVoKoab4PwmZ2fBk1B/ONSJOqrHVBk8URUfTU0lBFbb1zZUfnmMHWffqFIqgFX
hJpqQ2QCy/3kIOkQzwVVraIfvF7//Pnr0tQSay5EX/8EOFPKIbUBCIezVJ/X8+82
t4elQwyAaJrPGs1d/wS8ah+UPq/0rMAwECl2t5hC1TjVghyoIpQrJQgoB0teYQgb
/WBOCiqCXz/t+gcFOMT4T2L6dCTYFKuzxjWdMTNbldiHqpbyXZpxd6EscD5XvW4b
63fU+97KMEIW34ONAg9RDy5P7hclQdodB+PCIF7RYkgsNlxu6B8NcJgJ8NzDVaA8
2jAFMNjux9/cBfxAWuNHyhZGm1UzUsKBYFsOKUkG1s6LfN9tbyh7jUcXOfjz90PO
N9vudbuoS0OHNEpgsQdLrmlowQ290FBgw4LrflRsSfdqSvoKvQCPvIPRFNpTCRC/
r77g95B1212ra7tgpohI+v9NN+gDrjjN9sYQ374Q91o4eZFNcQYBMBu7tbGFwbLp
+aJxtWNAZgL1NdzA6mi70GtMF/C2XOrsjufUeK19p7y5eKcN3wBxJRMBV5wilPBE
wZ+z5bfaY5V6B1t0Ut6bLF7fRV91apMmgDfd+DffJaBslA+CRB6T7GqplK+ji/yP
`pragma protect end_protected
