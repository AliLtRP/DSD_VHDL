// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
G5m0BD3g5GXyhqi/JcjuY2njPC439TC0L7qk8wBrsFsGB7RVD1xz8YlVQCMsT3RK
FHIaErrDu3LmJixfbdudrhHY9nknwllF1uVyUPFmzksN/YtPZq+o/Ml72kCLPeXv
D4GSr3cZ4XEbZ7EGbnqyRFzebv4nN6fr/yDymZvTkJ8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5808)
wS6fJo2kaF2yQJRdSiMi8GlowpBCeSVB2YAwcPqUkbYqyMFrGt7oiBXH6+gkgn3E
qi1/EOyjCPNcAiFI1O3uqP+ffh980piVijQvrmTTZbeHM1Wf+bCjPpprJlazP9kE
ep1SaVL+OUIroDFKHsp4SxQm5nPRtx2LdNGGchLZyAPEBw4+rvk0U1XEjUxyG5sV
Dvnlbp1XmFigtTsf1xFw9QupEwDUUheCsKV56BUaRi2JmUvd2gGbVBQ2AlHTDHMT
wgz6sz1ypkEmXnohH4zxauAMppP7sGvFb6A89VwG0ZRNKGVgxseXq+3QJC2y/5Mb
jheGiOJsuG47AzuRL8quVj0hXZUgNgm/GnR/h/6KU3Y7c+t1e00p1Z0B6T6YXOeq
wPPfj3eL08qQWxiCsEqph9CqQ+/XrPqd9BmSVG5muxppwm+yarGbd9snRi8H8iDA
HQm7VvNnwwdY7Ls5nFzKELu1WOKwXLTdB6IVu48+V6vu+xEY7WWMUfYXpmSvFcVv
h2wzRX3GKO62mEBZcRnqXZU3n12x+6ViVTMJ/ara8uUZbX7mcNnsQYHuVBRKEtHr
9dJZeXz8hoqdwMmkdvnpE/r70eXnCtxJ5Nr7kxOUA5tb/6ESWBYahZAbUY3qOY0W
/MxvCiTMG/ri4VKUcCYgYlVO4hYYeO5GXRaCMM/HPFUKFpuf1kKPstmDiS1wm+zd
WOODUjkWBPKPpMtRrTHLEq2aeSqGuiIEFtjjYUm1JrHDj+ymEVVf3AXpFU4EHe2t
mD8nXpEQpx6W67lKvh40Akffx+DgOKVr+1mCEbyV+KCeg2tA2tzjlIdnYVVdDJKx
U38n/uN9L/NpC3zth3Um7LHspgFpzkgxgKhdzpAqFmZBF8JZQNrqEwhJ/0VMAPF6
DcZ9LAPWDACUOs2wuazci6Doz5b8vzHAa7PotxD1ZgpBTYPLoohUT9d5ZAw7uile
TUGS4mulTIbMViojg0pZK3dN2sk4q94RY+qCfAjQlWfRXeampr0RPs1b3Wb8lvca
ZZbbz/ZWU6H/jdV+S3IStaVtqx+QrvT/n3eDnju6d9YbUcfxcwSpILoKGJMxuwgH
hGg6U0agEM/bQgfrGhA9OqBBCmUbvrFhkGvvdAwZ8UYl9f9/F0RNo3aWzNCLUY9O
Mu9u0sJa13sI92u1E0MPcGlrJCFQ9rZ4xbbCNsyTZRKzgr4bPY4aTdH1jWjf8wGH
ceP6CK2v00zocX70klMDnS8wGqutrsUBT+6u8pqhg1KWHC5NGTKdtoPC3hAkv0rZ
nQoQMFWHq3ATejF2PwxCBbU7w+jtOe7OgGEoV+ODkeGyqmwpPk6SmcNcZp4pCZR/
SSseOSRtVOeOz+Fg/rBzsZCcUmFtnA5pYDbx+jbOsQlflZK4yG1y4ZCdzT/0Y9KC
Miy+janBu1sDw93zYgxT2nr+5WhugMw3Fn5NICpyhx07yWrl6Nuy/VoUTguv0h1q
03CjtJo/XrWWBkfowYWZkk/LeApQ03ZNzsVftmwR2G/fwOhZZQwAaW+bvUlr9X5Y
HrV3CKhe2yTAGiUU9sdKprsPqKt7TUrFN+nCP4cDcCqGFd1EBCZ5HSMDt/rgU1BI
n6dJfyulBsObT6Xz+DgafR5f7Nc7o7S7E5RSxvCHnf5LXluDftaOoYzuGphXWiKQ
q0G4cjxj7u1/l8JLAOvtT9w/RxzXgjo8ObPuxo85qSSklk6e4YhXYNIAnJ09dLFj
qcHKo7QyQVC27b8bY4U8UD5lYervx+McNWJA82twLDInj50XZlec9RuI9I3d0v0u
nps17IrlF1q0qKP0HSTPmC4pY5mB8VHtqNgGif5sOW0EmtAC74HnVoVxJchjMBFK
vxQHxla5HQjJKQ3+jHVZOtvPzDY6RCIPU1K/If3LC8lH0mZg6K+h6/U0Vm7eXqr+
5ix6A+kLWBSKfbwtEFnggJXcbOaOC1tGTSwoQPbfu+SxCBUC0hpkFPq9d6Z5kP9w
ZwAGx+I55w2z4mn816LXUi1ZQwmI8LL7u8wwhnLkf74Gu9VW75fn6wFPNid5EvkB
gYkqX11UDFuNj/2InOP4MkwECB70Lpxsf42sw8Jqa/GqtpSm6RWWJ161H9G4rAFi
bLk0zNdPZQ34NNssRxhZaA2Qs7QNNq9yjTBLjQDphFPb6GFGetXiJA99WynJiz9Z
jm3DsGrNL9wMO2MAkJnOn37yGPF7Eo7f5Zp0aWT81UitxaHkkTFqaNumsQ3iTTMx
95qAm8pkaHBJwA/nPcPhn0+6C8k5Gn2dIv4x5Np1yNL/iQXdPhj/MRnpYAHa2eMC
w7WXsqQfUq8rsr/8byvbFvt844ql1rqqidYKCWr42O5FeOp8ewgqBojzq4hwL7H4
ZKJNhjGwqGyixNUAJINvS299TwSTJlJTe6iNBz5D9tGecsUIIyBbT88A2dve/xiH
Rv+09s2fkPvlRrVRk5S8JPuyUPseXiZS2tnc1T7au+KMMQQWdYT+cAU/RUNWDCZl
R/bdWkjTxjBwa3AQ99uZkY5wKMXhX/i5xJw4E4f6UikCrIvCP9c3RlSg6F5T7Z0v
5Ds72gK9RkmIre6nt+X4ohYEk4tRK5FuYDL1CIVJDjfQLV6pwvG121Seh8A007+X
wx3MI9whddQFXkOxeR7nUJpYOS+izni/08hnkSnvQBkk9io1/ObqVLZS5WmmVksx
mrM8vvVQkhiWue9xUE7IbtizEYYByHhAQzO6Wo/mWCAPpTgvZUR45T3oWo2Xroc9
uLpVg9FAHqSjFClwEu153KAVAGv3xkG21NqJPitfwHkp0IWh0Hymnoqp4QZlTvpC
oKix1ZuDfXW9glSLkdth3WYsCNGqVDHQQ6xr1IaRAXTyFQwwv43G1W2Ew1Qu2Q6U
drMvLPtxZ7bcU26B0Vtjy/HP5VXMQUb88IgnT+H553RFs5yXY7+h1lrpQalAw45Y
tacXZuYm0Sl62AIRnt6jhYfdm8T5sVqxQ7jT7TXLijcblLLWWZXJ747j5SKyOdaW
ApEw9BYzE/idY+n+TLLe/L3pvL9cTpA6UH5DkYNbwlpzAGtVuHiuDEpPRTyZUQVl
4aKr0/u/511UoW+fzc83z5S7bbeP/UGE1VgAKmsBlPl/wk04Z59HSBHnptXv9LCA
w2oq4CWd4ME2YQgCeBP5HyGYfQLzFn5RUKvbfkuNA8jTAjwpEeAOUgoGfIZ5u0DW
L17MtsVjhcYtV6fd1muLqPJNGKPOySuCJlnJfyc36L9nzDIHs7C3SEhrDGiv5nsW
3GYWBK37bVzaXi19kh3jY+4Js9Niav2fY/lIyHlaYa4plooGvPhYyOqPVmk2PhuO
siIXxrqbqoaIenj9WUm+AMHdmT/NC8HErgaUOTCZx8F+BXaZ2mXAX8ldH122uRVJ
2qVhQSBF6CqxZwph6yFUUBLOkuVmvfSG7+DUYIPrUmjt955URS0jw5u0OBzOMfPH
bbYvdozjF21WbPccs4RmUlQqZhYP9omvnSYH/nIC0CKim1e9zAFIG0I2uv5K+m5o
dt3ecFtgzxCp91Yo1WWIMeVvIIWuIXmtEg0FzxnqwexAIACMION4nOQ8d2fWlBAJ
41WE6TPZFK6xSqR8IWDOTp/ycxzvNdAvBx6FRYhWC5qs+ApsykHLHa1WYFuuHPZT
XFnhTkwuBCA55B9XY6/PRoa+QkiwqBdM2kAOTwYsjVGfRbr0pZv7Yc4hGCsFVkqW
lrxsu2mqIvbHddKVw9Jn4M8igbLnmnjHpgMCfnndNJI900EE3suBXuarwIBQMiO3
LlMwFW4MDnYSiN91acph15dzID29efq1owG/4xOrMucmsz8TQ1QbZOyhfYd0RSY7
0T0V1nvwmuXEZ9jbbxv0lUnHtpyLZSiuUD5CK/SjofBydu5mVAUkOBB7ySZ0cyAa
XplzcMVgcyUDhw8ydWC+0Lnq/W09/c2mCU6gu/olFUcUlQO4+Fqo2IQbkX2gqkns
i3hK52V1Up2RoTNZhZpYanQD5FAxO40T22ldDbF6u9lZED8mv46lGvKKffP2RxUB
e7+3vLgn4XUh+MO7qlf2kExwXuNi1//alM+ju4uuf7AAUaAWXF49YPNzYd8Aa4Os
+Zb+t4m/ZwzO2QxjzbS729VxWFjEvkYJdOL7jsj3J88rU/MBukGArtgISpNlYSM0
MyjtaorIt+0U3Il7ZQvFoZYVwKYJ07ahmHI6WPI4Bpto9qTyHWyymBSPiTAlYeRs
qcipVatRj2RahevzC7a1u7sd4yBDO/H4d9X2dvmHre3fWiKpP0l4C3hGfS+5faJh
vW07FyUGiEXIlDe4ulOMjzaAglBntL/OCx5TFsv2u5UubKO//i+j4LTDDdZO9ImW
IKBhtlXOr6pHOEd4d69PTvkVf5/tj2NSZx5KiU1+2JiTUt9taIUpFfJOpmmykSzU
ICbaKkWLQGJ8ECyafSWxJtXEoywDw3k5IZl2IvObfB0+S7aA2Wh80+v5jbU1qAoJ
Odu3QaA54JM+c4tNnNU7CIXHsXMo6CFZjsLl5DXNMwpc2yZTwKYnrcZx0hArljUL
LscT7MPx3Ej9Ab6NaMHovcQyzh1km//zUwhG35PoPCLoXZshtboO7tlxWIC61qfY
5aclg0Tv/8DPWZXQNcD0nnd3oarln2olcKXLzwFlIo0ofjNOLLxNih/GyDAuK6Tn
uu3TptSum8hTeiT/VUSXnh8oHwcj0jdqCh21lSp0c41hWTywwODk9X0NJpXSOt65
mt5Cqn+VkR3e4gHeSh4zvk7QTeftwRWJHkzGRSOIP8Fg7EXCEk2TA8bxy5g90OFw
pB5cLv5SyMuLfk+QEKaxdz66Frqtp62HonJbIydPp85/C5WC/rlFEjFusJA8s1Hz
OSHtmfmhLrhURH6rCgcGW/evUV11/0mMEuxH6mNsAKPnnqqsQ9mcX6Xdwci1d7vi
0D4cqEKfSMzS739GgoURvbn0g0vS8OXg7w5ajnxdQxYQZtw+rgn4HnH11EyK0EDa
FPzrbVla1YGd6d587L1RHjxefkd0lYZk984Um6SXSNEo4jvuTxKp0/e1vgJx61md
DOxzrmJocvE5CIyzPHxY8M91HXnKr5/+9tEau+ZPirX4zo6wTtBSKZXNfCZVuQ0e
onIIstYpDdryfAFrphfju0ssjjRbUYDXQtwVcDdsNBJtv9D4XkYYFtaTWQf+Q+gI
QibP9ThxWW28XnzDvLaaxnH6qU9IhCLnq4O3HjFfCosYZDwyeN5CZgjIPGaZKBtZ
lp6j4cPUi9ib8hhbPEDh8sDUd6jxn7SWzyIrsHHrV8xzQ6kB+ZJNlvNsNizR1CnR
0/l/k/+Ize3U7/kjogDMRaWB7EwdH91Gy1o84Ss1Xbp43/f6PyI2OC19VBMcsJ+7
f6Ro+lR+V5iVjiGn3BpzUjj5xTz199gLipApqyYAcdLxV3bSKydcn9nawe3xK6qU
CIltMPr4Ulnerqp9Vx2voLRwyMvF4+ZYKUPitvKdd305kCuhLseytFxz2X1ka5Wx
p+YzNh1Vqn9/EvEZHi/AkfEl1e6iCO0mr5qt7xSPHqpkssN2umwEYYwZPEe5Ylr8
pdyHe91pC+Y1HU4bQYxkQBrhy4MBEwYefbVKdqD5vwkFfA8HhpxAqMuWwOVs74JF
BKc2Jz2pfs+grSLdT3my+5Fdt5IZZ7zQ17jhDNAGl2Zru+lPXRfMG+BS7j0sJ59Y
37de65G03LDiPwMzk/ucldbIbCdeFlFtwvZ7YWwVay3t2/az6FozSFBWZW8UzXBF
EObW9blcZCapLm7b7No7MdLm3evu2/OoxDMrzmQD4GZAajNDMH5pWZ53DyToJKGj
tSJU8C3/mWEuriMj7MWyhF16WU5WUcvotiQ2JFlWbl8K3nW+Ep5qtIMr73k6VOYr
Cr62WsF7BIZ4wGmHJvYh1Qd8KLDswFzNVAt9uQD9EdNmkR1QGWkyz+Jl/9kpvGS4
WCzivKfSzDSz0pxb/KC2SgE9ersps8tyltYhoiluzWPgRdvtmdHbpXoRYkacNSZO
WoyX7Snr6bb8gf9AS9DvthDlncYUkL/k/8O4QTT1aYlz7xPrivSLiV7mQ6S8CCa3
LJQHhXQhgdrPQadAjZIPRuz/aJnnKj1Dzj48yb4cP/vJyrs7jORby/Dk5IRoZHIU
2rtLDswEwTuRz8Hz2zgIfF5h0Zy31DkRpmZWscSlayI6wdGCPSjKn2J45CHgCUku
wzpkJJ4qo/q180jmiIwdGzMFA5QeDRunVs9H+w2VHIkX9sDCbr2L1fSFdOkFCXvu
9g9mMpvywuI7Rh+PTiBQifIjN/rL/MR+wjoEYdFQZ3YM4vF2KX/PAmw6osd3DTgm
Slk0Zx2Zm+5viTnE4ly1dxqGUjzlArB0j38V8T3FxA3wnmqsBmUh55J4huSw5+EC
ZhdqH0NL0iNntkwoOthe6XXvl9JnbaJhZUKZe0NeNaXiMpmUTRX+UFvaPxOuWTm9
gRqDSISerF56dU+cDVG8iOScNAQrXsdnWCnXzfw9HiAb1x00dKBk8z0lmwRBFSo4
iKBp2aee8o8xgpQXyoPILFn6muPHZOoVgIzOeUxm+E/f6wp8q86ThQwOg2p9YcLe
FVptIp4gIPDb08s47YZfVYlCliGoifDJ+/wqmUC1nP/5e93bPTwZOWiBEZyonOVj
59eOgNTV4n6z4xxNaVjokPCQy5v72y18ICQafBak25Sge7BNqOnnCvcFndXsgaxD
Q2i5Pe9aqKYLEs2WUSiblwCf53ut1DEu+EgDMQvg7aTTenZYzOHMmscayvchQRGY
JCJvzgwrByrEOOF534QXBHzu2crCXxhMC3HcDeMt5KgAtcbhq59ZgHUjStuPvq34
4jX9jnAYgRbJmwEn7X45Iijiiy7DnyDX32JgKbJbsHoLjRNgFPxSrzfTgzex1PJC
emm6UJnldIFVjBj0qca/pVx/2lq2LHa6PY87iVZx5I+XpzkynlMmDfGxLJnXB9xu
bBoPemOH6JxgpUwo0FHcvgZoeg9qqne872rmiFZQRLlld8sQztWpApavnbO5nUzR
keHDFaxtn6Xx1HOF7/sByc/hFLM4YTswDqRxHFs6hgyzSZOfK1ZUabLTULUA8fkO
jHCqNBBJRdww9sHo0SIv/J7UAB8iXcR+0xtWnBgvF+6uCY1urVMc9XYDW+5SpFy1
V0cOdzG9x+FIt2ITKnyAtxJe8bRzW0uYRg1DciWvpIis8IgRNhRf2RBSB9yZIjw7
1VMOalh1OIBeXHY909OeT0upG9t6saO9HDOs2otKakfF2cTEJUjh6jaib2csAZkp
5xXjBIiC0aqGRzUNUzcNELJIei/c5bGZy1X3JkFyDJf6Mrtr62nE2alKLiTGSczj
RrNX+UKF568ih71pnKrXCu5FIUBKDgv3xEYjoVVAI7jqK3XWreNZDH/Ei6use/q0
UcFxRXzHPgFfPSz15izcZFhMD/BI01+CgnhEQOfhnUYXsOwbQhZTvgdHxez8IOoK
ydJre895X2kUS9bNBoBJWaiXSA1St1wH+5Xw2Os3jbNp9oPMqXUGjumgSTD/cdaD
2dC7fDcZQg6wY1j/gr3+s+JsCODitSA5c5ypDH2Xgwx9P9rSe3yW/6CvVj2MJ2dP
ezoAdAhOW61dZ8lHc32B75/+af4ygOwU/40RkN14jfcMM9ml0jjj4CvNUg51J0FA
esR/9bfsdKajitBBVNnyPXipy9kD9mQdolQ/cmqcfPp2AU7e+m5eT5orsMaBfzCi
`pragma protect end_protected
