// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:12 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OhKor3AdoZkmttwjP2j8sB6uSDxbb+terhVv9emPAHdyL+WKVObJnzy3DujIKz4U
FMxEyZA6rvMT+y+BAXPlXyqSnjNWcvyJlAw33++5MkZPTsPsL3OvlEZTnYokKhJW
ZQTWYFvqdF4kXqrIeVyokwC7eolQ2KtLgMU4KbHKx1o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16288)
GYvcBZTCEyMbWuOYlEyPeJ8ya33WCqsOoMZ6Tw+IhD9XDFy25G0no4oTFZqnYVrJ
cxBiDNobSnv9h7fcjqyJM6oBGzd3AaRuMCwlJAV5fcJ5OvhCE8900gp8FdBJrZyg
23uEDJjeNgIdgu4rW2K9VsyWl/BCOACm7a0ZQIYAr0bWFM04RSsojWNkFSENnX9k
m/q4Vohmz8pv2HlvcmjFQZMrteBZpX0lmjy7eNTitVjOytYhYtcRbHOE8qljM6km
EoM6BX3JeOgWdAVgwnWc2c8SW8wR+9gLafROfdth6Ug7s1ScVfgv+KxsYUS5MmYK
OpT0AhdSGNL2rFufP5XjjfzimepWz0290BJMeX2d6p9icNMkWanirl4bdb6yRsiR
eJgWY0tizgodijmB5dI3/3IiU1H7zByw8MbXamNQE7b+K4sNEzK+CuxfS5gylbBh
uon07L75hk2cEkgznPaNAezp48ayjQia8O7xZnWcgIzy3Kyia0wK55dOwBiDjhg/
78hwma3rk3Vg/9OHs1NJDX2Onz8939YP5C9VgTPfcL3ayMu2OO+LcZgNKv8JXjbX
h4ZRt7dkOM5gjv6cSsozxHhgbs54zdKuf8o/Mvypi7/JtpNwiydJQhFiyoh2qvrb
WLx9dFSwCBNQ1Qhi2praj2mZs8Fna6bd+ca8h8KbWBriYSYwcoj9IfA/FiWyoTJ4
Oaex0BV6pG2juwqpgxl+AJ4y9HVMOzxDNtUPNsnJnZo6IrthHLQTbCw2ZDiN86Si
Pviw+XE1xhCzo3aAWBRj2SQmCQSbwrlZkcVm3sZnsPWJ4Be0N3nB/Y/4j3i2auBO
Qm18YeHnvOJO3tYX0CBcTE8neJmASWaRlbp1t+VGEuhmaBpOIyexdpU0/Rbs9CPM
1GwPXzM2huLIEIy/REhVPcSBhZ3G82cuRYRKtSPGqvgQE+OIJpyBCzOG9Pv/tt7j
Wa4RLgbFXJE1+LRVwKHEQcp6vM/itgR00BdiVVS0kxWIT12tyrFA15vIzpE+6AjW
AMtTMp6En2DdGQf0D8cpJFdH4W13mm0/l7gTb4sLL/PJp+Gw3llz52YOZH3ugKHK
kzQ/ueHlW0dbtPrRLLnydcWEWpFyrpPNHauiSUyPh1RbWJ0xJoLc0cJBQnY3MMqJ
Xydx1kOoxzdJhy8uSgeAEDKQ9KslxdaYhiZvU5/NAyf0n3pU/Xfiww4e4RLmLLx/
tb/m0m5wkG0MiENHg2jgtjLeGihSwN5Xg1kZg2s0oyEBY8Nsak/n4ooaqYiE4hE9
f4kXrLIvpwIH9Txf/tw6TfDa4WBXuAXOaXMZemLzuBsdiSFOQL9pNXT0icu7DY3J
zVpmrec9l830GSOJHCKx4ZqK3XLmYOdWps6LvdAnP1Q9CncElVJGiAS8gVfGW50Q
ojcmdeo1wVzAG+aSAegOHOK7YLAm92XmpS8V+RkOvYoF04enueF5j7DQPvIvkWua
DLALkYE5lZD1XSy7NhRPxokk2SMAZemFchYxvNUpVzQme6wBlG2PGbA5YyzLmWxK
qbgioAg1NQ8LoZOBpyUagOOZsoPi6Fqg0rh/NIwI43MKMQkInc8qWkX3tTvitUfR
PJv3Uakkrv1dzOKZkypZoYHiZuonFO3pXpP8Noq68vvVHwumOJTwTf47L8lC98Y2
mvL+wuuYYY2JHPWLcX2hq8ynw8rPPyVbUtahrJPQT6+EKptqWEqoIFnhIRWjcOYq
O1+iGK90CNBPGccvdPUZ8EMzN36cE7U5Dcvf/PgM1BNrSOTiR6p24QQc3x84XrBZ
0P245WtXBn9WzW8rijmhDebtrxbYXCqujGFQkB8K4BakCpxcGRuTv2PGE3mp/qog
5qLn/zim08amrhzaRb2God8b5XPQtQQsYv+MBrO0+QlUrTEYtY/bddxISjRZh+SY
NqLjSXOAO2kNzPFcQuaHizbKRdp+rxoG7jd6HfETpHHzI8jCwMXXTlkIbW0JoTpS
mm5sXupulN418ROQWS3/EqfKg/Y3dgVHnQPqeQYcLc+Bnh8apTick51GpgCLhXa+
QO8/yWEDypc0tCDEnGcFZV0k6/+USuFebgf2V97BSAMohbkoZae7GuI+f/1sr0re
I1BZxaWy00DGc6yRpae5pKcHky94Aa4u9e0ZyY7GtAwiEbThbb7DaBbbP4e45St9
a8pF+JfpxE2TapnrAIcDvhVz+oagi0sJ5GhSfNPRBrY8vyimw+aIVG6tG1dTd6oR
EDLqOpdDqHe3aeA1Kiq4wNO+deiR3TlQK5ZQODni7J5v2G6w2DhkTMwaKLVj2cZI
PKob+GwMKO1iIEYT3WqIbaCqQEw8aQ01Ad6UFUec6SepAa4xFQMUA/Ay8xXjGF4Q
1IQGJ4FRfOF/CqlOgn6Uq2dZL8wwZqhU7F079Zai50YIu3MNHLLN0Qx3OrKxLsds
l/s7gx47oU9aR4f4VfgU+xZSar8KMLjqg9r6qbW3SzgDblhTUIB+gAnO6Rcvv5pT
PfV87h39tWidpV8Aa2wOuzo5FLtUeCHAs97XotouYmykuexTzQWXJUYAAmudJjUx
xKYZaeE9dWzhINiouuCQP+S6SifP//udbRV/eoD5C89iUlbl4WLaAg9+Aec4UkuN
cXaYUh3DxEn83y/qmW3P4Lag4xsPH/E5GCB9562A+Gth1t4u2TpeCT+d+rSV+uZ1
S2dC9MufH9zJ+IxLww3nlJJYWLLUKRnJgo7ydvz4h9wWr4t7zgWk3oZ0jvY7iQaC
ljfYp2Q22t+7XPJeo3HGqd/GHmYC6utTQk1hR3hai3CJt9wCMGyQI0ojn9giCZL2
nOJSkIRzd5pHTfppBuumbMqb7zRWwQ7uTHqiHN7YT4JQId3Tjpb4RnT1quhMa/cf
ms8WU9GOptDwSTD8xJyzIGwx7oPtn2QGPD4CLxXdhcUrGDjbOBzuW8H7qyP+3dAm
36PjtHaDP/TzOPQOyuqZJRBmsuYH/eoa+XGbuxAp86HeWf7w6CqK/ft/hDFEz1gi
tBkT6pXaP+HeL20fSQgVMC02j6LCCTawV59ocmUHKceP5SvlnYrJ0DPH/K3flqub
/q0qKtLtScrucszqnsPhif0E9r2Xc07uX4+KW0U4mXyGWhsCRzt/oDmWoXG/Riwj
K5zPyMZtHHUQZXZFhxv95ZLIAWz6+LFt8aV34VL+gNqh6IxVX6nrKSYoA90ta1UV
vi/vTsmcZXCm+47OgHkjQ7Mt+YRNx57vIiJACZo9+l988tiP48JfMNT8ILmuKXRH
IZMZJKfZZxZ4Aqt4Lq/vHiPvsmERBxGAQRIGbnzg3RN84fslVETJROD2xNodduyn
S4WHGK4+u3yDbrfhRQTZLN3vuqh73RAf8Sbt84gk348Fan4zAkPjY8G537zetyvb
i02GYJORTTFywXP76LjSu7zGa17wURjBkvvLWc4vNrQJVZ0V+3RjWSd94/DMJiht
CenQ3wZpOxUxIDHyMIWh1ZK/Ds03DLVQ6mYjgZ7CxvMZpnf+OQnMAVoZc8sJIr6v
ZhaVLa9oYht3BCOCDnTWLDP2VlyUn3B3Y5FdtHE0+FK8FCuATBRnLE+SqsKp0+HB
7NMmzgIqiwYpHMiEbrpqKLvhirg2v9gW7JyFF14UWcZOmqR44EAcY3WOCb6RtDYO
AEeIqrLQ2wLtncMcxmSR7My/MJyyQf2ZGWs8Ky8j5ZMqtwJIqq8kdxyXqqRCP7zB
/xZ4nPYzc/X4fYVQyVdgVv1Neco6Bck/ti/MWCxN1EvJ6Cgk0y9hDRnua/xc7ay/
qsA/MCPwHjR6Zf4ZS4bnEyVdl0bBzy08uLqAessocyEFWGX/HnqCuWTL632TDown
JqVYB94NSCjklqQ72Itb154O5vNngPA+K4Ee8cOk5xnPlW3aimpvM5gOZglq1cka
MxgFXWFCtlgW7jrfg+4VtN/dVLPfdc3xcZWJfC7KoXWt/uIBg3IJPcfN5q5ygnJH
BO6A/LudCmvGmB4/mb1YWgDAY7Y3Hqj7tKZG7p2sY8BVC0my9XCuTBcW3xmxKSU9
pIZE6p7UfeXEtIEEMtJ3IRPodxKgKSRH32ahoEQxUuePKwnn4gyE/fxecFaobhv3
LSJtZO+4F/r0aE2PI1sut7TlT5CHi+fQRlv08qKDM8ahw6ui8EXKTt+fyykS/V+b
J7j2p8sTrg5o0joZsXB4NKXd7KXPAAcSBfvv6wB1hnwXjnrRLi75qovgx+PWBiYc
7hyXLe9cuZmlLnAN+ile9GOytz94siEGPlmjzarATV6KrPoCi570A7zypV+bHwwn
XpzH7DJGHboH7VmG0uDJ0JFFUFEwah6S6JO4hEkNIgmxpKLmVJYOgvYDwohwS0Rt
SXJVxdIeyqCqCtPtKt0Ex8aYNz5v6MvtFL7uzu0ZFD7W36IRvY4v6fTBqvC6LgqY
MP5rKrk7V9rgro0yZBKd2XESd20mn9QcHu/Xcy+Jo3qkmpmSAj+g2m5SIiLkCiyF
h10JTo/m7ZjaKnv4W2S+fW5BtjT7tUHIQJxUVA3l+xcvYWwvGKzv+pGWV1v9CJ1k
0Ep1IhCYtQPdYhplPCPtQ10QTiFD8Pgb/YKOQD0RSoZH/WL0jL6a+0cbvUySimRp
SxC1adgq10zP6nqTnZxSFQIuKejvvpPlFZDT4QGzqXeUlrBl/CLz1LEY5etO/x5C
/ceOPuVh0cM/s4J7jYgFwL3k1s5irWRbBzjj+9XZ47usWbb2mzM3830mwabLTf2E
/g5D0nS0IxUiSXe36impN1M349YQWxesFYtGfGE8apNgvBecqrXFVH0koQX2ATAU
fCFsMvx4K/xokYBVWlWfZyChPw6LIMPxi1+XUrxSpxeTZ/Bcg3tupzd2sRm0/VHN
s+OK/owzeFpSVFKparW4EVfFRcH9+Ywh1crjtuP2JhYqwKoZFrCvXd4HnWdTVKZ6
4GqFmXcAAGf2FVYnPm1rgaMcd5GrrXRD1rakkd7J/qd+jnZIT5O5ByIEjIXAy7yg
5cIjUq4AICbKvYs97kIbAM3JlrDrcy2nhIZ1HDWT0VtQveR7fd12hxOA8uAZenJ2
0FIze8e6WO6Z603O3izu0dE2WXLnvoXU0o5nC1uEhbBEhYeIR5SRLrs4BeP/P+Ml
004x/W+yoYZc6GPj0T8koBOxX44rpytLZexyxphgvQBczZk4E6iDnrMp2DcHmhIc
OcP8znE6/6FSscrtwyRil5s5mofJLv/rYSIAS7vXs4gmFKLFkZ1JO9R/etCiGvQf
p52/dUgpJJ/xFFitvMQ8AiiaOJ7DoEY3VtTkPQhZthbMH7bTGzaTiwcWKFZ2rB2W
WGf4obg0A8C05lJ8MrtzjoKe+iR1bUli+Ad/mE2Vo71n3fb9yeWzD57jjJzkLlQp
WqULF6aSUR2oLzuHaQOmcKkww90FM9xBgfYrxGXTYmNDIOW4Ih92cWurNqZA1iPr
m5UMFrfb3hzDpX3l76+IvGRrdDbEkzuvh0DHqIWhkNwypCOiW/wA5Jj5H4GVpG6T
0Sa/ql++FYoVvJJ5b0BY+IKYU+rZedvwd56HgZWV0CB1P9GHzYMhrBCw5M8Zp5rK
z/S89IkYSXF2CDyQ5p8SspHwo9zam5+EnnFVs1mZLcSCcCm2Lc5COEKMy/+wvxlC
2/JIuKM7x20nd75Hnp+0EUXbsXENBeSvXoBdwXLXQ9S7ivC1YMVr3NFaAXFTemIW
6qzHovV1xK8hr4f464dTEHzJB2970/fQh/EUP7z4vEYDd6TbETWULV16W6Vlq3pT
tIHjQ/ywiBxAEXozWLUO9KG/o9G+dCshfa9gjXoHWvZ3Fhxkm+gBKSmYwNJ2U3y0
dhdERr6CTXnFmvLOJAk5Q2CTufXbkHYO+NX4aECgXYoq9Pqu0ugPbKo/7qE4Z4Rq
4gnFW0/kCMKHepL88DgjUGkW9CnyW/ZRCG/tC89MfOMNOLoH1TKx/HkN8c0E7B3Z
CFGqVoo4qiVclzgzgW9bz34GPkilLAc7Nd+qcARjQ8cji2bpWBQklqZzE4wf30hb
OKNxk+YmOy2u3EQiDLmZPXMIl1tWBZlShD+eFmwu/C8O2/OgGa5jt9Zlo+CfMRoY
jh2G52JgUG/VD4Rt+2tmPWnrt9EEMnXURmL+xf/voBSIe5jzP3UqMAItuA7f4Npv
wDk5kwvRbXB4OYbyafITe9OXul9da98kjk06dNDG7ywFKEy6jwxcmyckmpOnDxvi
acFY+2lxeglkROCIW6XUh+9qz6LQgIBQXZcx+5GAXhR+IzFfVo+IM89iVzY1lqtj
JN2UK0V7d8Xorx0Iji4c8dk3r2IXwJwnYVjeLtUuXg+Drj9Bo02hjkXDTekWgrl/
DHAoildtt3mPG/XQJR+51O3gHg4RyofqHfhI5g59c0jjPS/NxJ/Px4bs4diTusxd
mtNnyA6KhcLmUv5qpLlR2L0zO6I0Q4/W+5yefQrTa2IeopnB4Xd4bjQiNHFmkUa5
G+WjGoT7LEjgXXgBswPpO3AN9gIMqITgXdlEQfbbrxBsQPvYRc2ukilQIL51RF1U
B3SDi+hNfyfsyooWly1DhM+DtIjvFp6SeBPrQFMQYBzo6ki8QzZsxxA5K26d7Obr
Ry/AFn+Er8el3GNn0WFmj/D6rfzmfJ6W9iLiyWTEXXQgZFU+a1zOjG3mGoUdA4R5
ApbgJT3k9HBsCRWUNA6FB4INLmIsYW23aubkSCL1dQiK8r0VH59uXZZxSfVYT36g
8ODCXdALexpatihlckI+0ZS4NmLLJQzHbGhL5PAwSkqhEtK8UIsj6VWjPu3Mxebu
ZgTS7v/GIL2bfwwHX2P5GrSfXlAq/dPfdZWYZDXmxfLHCyzVY/aWOCNQwKVjGUX2
yJKEVtbEgR0FLdq88XrHXCE3ydsIauTjrwDTSGsSHxTHjVSZ2OhGLvr7+MMcH1Ev
5Rbib5rQvo75sG62rsboK93ju+2G752lO3mWJiSW1UvkFxukhK+I+zEt2H2dfWBW
Mgrm/ivRtgNhtT0t61iLpC5gLS6WcerhpFfAVh980YzFzS7O8cOIoAPhuY3cB7Ri
I5XhSGHuXGcbZ8U8rWNXwyyWIohCXoxaGx3/EtCba7CfwnGWC5CMnRCLgtVToQ0D
EO70nwSuFTuOr//YXT4RUK0Zpl20Pz3GYdW/iXJGdAcZJILLIhEa3qOt8lY+qzZq
RBhXs7draWLqC6LdbBniBstbdi9AnGpCZ7AWKKB9mZFmG6PWLx+G++cyU8ef5fhq
UwlBJ+PI3GkoP3nyYu/s9A4RYIjvGUoLXWCnj8gs+tvqZZfyhpljKMLUXPTOsetk
rTmc1wRciBtjVOPzMfXiDplsQOMD5ySWMT9AovKVjnrdo+526drX58Lt1FmT/O6W
UVsefaKudm5erDF+hFqcseB2+4Xc40agyvWiPE15hAli7vhHx1Zf1iHwPpGk7waq
DL211voeyx9XAhXGPc2c6f0RRfhkYLRGGe4sEiBXQHUDMIUgMQQ8Y17MyXfHb9uO
Ggyxxx+i0JZRs5NLpoctwqEV0iHWmBFlGmwrhOyz2vOyRTS5soqwZqE+Amiyknp+
o+24QCK42xP55rHPqAOOgFks69432JLMVCCJxHr2NC0avqmrhMnb9kp1VhfNAykC
qKYd3Qpre4orDDU/6uOcCMxuUdWuUJX19QR4T7VTsyEp0GRQB/JiDsa3QXIchEa6
tChXYtpW1tLVpwtPmV1uVZBJH7iQOsXKXr1N1q+JBb42BD4SYO31nTNpJffEF/tW
vUmh6DWtbc62NsaLmTr0OKH6pYnWpbc/etsJT/KqT/1wav9WIRexRfB+VAALYVRb
92QN9D0v1yNB9onnlMolGooJ1THsqISy3W3z7Oi9dQeG7/jRvrqQ3Rtd0D3srm8G
EFVsM2tGbaRhY4HngyfYQsRFSXQsFM6uSEvRMGui+UNOXaDWM7RxKGJC75qSAKQ3
1eff7Wyl0hMurtr4U1+QRwhPJej/95qEWLdeN6jaO8bmPBkVs/cI0RzPpJIxXUNE
uP3PUcrtLOtrweL3bSu1eQSmAC4GAb7qD3pqpolj2onns0jgXpidLSwRcHmU+7ni
uLDxUrklY4yX8tJNvexnm9sQijLxSmMJQ5R+tGu4I48u8NwXlmP2QZb1StZXUNei
3alSTL25VJxlRoulX6D6uBJoUz1vmpAaAJj2Qmo6XG0tiXVaXsHWzpA4g68D+Gg3
+kW+SznxA0yl622ehfTQdL5CPUKGprfHBajy+vUWCj7YP8guMoTR8TQx0WFdIBXl
Qiuc/AE56L44UtVnUVPoQMJgsIBfY/A5+vHotPPzeR1gpo4EoCdqahOzEDFgGSub
cynisq70kctrOKPlGIO2nNYDGMbbuqfvT51k+arNr23wdH0tzENDBdVP+YQozxB1
RMnQ3tjKyyHcA70ixM9mlr6cH3Vdo5w7k8pWsj/LJMUJAQGzY1v5EL7f1SOrynAD
YCwDaTpRF0g+F0Ltdfqshsy6vo83kQf/fftre4b4ZOGH+e5LwPpnDnr8ZPH7yGIT
LbiksW7ZVVJlKsgoGTVP0Pvpbg3dFSTKFwhTG6B2VF3hVrY980MCSqihK2jo14yh
foqHTPCdbbTJbr91QTJncS5NezwENUHrO/rprU3mWXd8RsiSxAoCM0tOJPcoE2cd
JWMIQpAjsGIEWtjWhXbGSd9h0oqcYPau8o7HQyHAp929ZIkg7EEAj71VEYI8cr6q
Py8HzZVSyyDq+8mep7tOCj+rE+WllYTjMjn/cl0fpL1cSuw4n64f2k+ABGoV6lXe
lzbLp69CbINECX7lPiqMn0/4mDXJ+oavY5c6R8ZGlOShITl21wZC/w2xs2IMI0Ik
NSjT/k6Z/u2QIavoLvwyi5YQG2ZxT+6NPYz8ItRka9Z8f/3FHkk2hDpeWj2VZCJC
8UAWFUCjYQLmWWvcloMJjGptW8LnLSOH0/0TrASXKCJrpRCo22zari+sfxqBluN7
v0MYYN84KBV3wtVpxw0/gsxWl77qE98rWPNV9+9mUe3c2SD4zAc/KzFo4p2zYxG6
FNUv6N7V1Hx6H1qp0giKBh4vTzfK/byW9x9p38K4eVl+OdGr8J2hsSns6oKZ3FjM
g9cMCo2r/9Fh0IRjvWwmpSoNv7Mz8pkh4O6nAQ5lhrf0iy5t8M9McJefWTanFGdu
PMMjvL2oZdgE8bkiP2Y+Yg2d6RRphKaWXcsyRGVvkdLdUIyv9ByrfZnf2Kh0bZFr
ZQSxzRuhW3COavHKRVfYd9c8usHKfe3oeDHhgVY9YFpOqRK3U8qt6I8phJsoek8Y
17UMz/9HpX84WXgNWNrwdL2xoy2war/riiCjeKnuB0RCDStGz62KwDCleunyXbls
UxOJ/ubcjv8mDFSJct2tHfffrmAO2yUS6nKTPcXSB7a8HnsdbnqpoO+N63mZUJkV
yuSb7tXsqTCSX6AIWvLkQ7sDtS9xah/yJiNZA2k7tHHcBHT/48zdcZiw35ZW1v4i
vD7vQLWzsMHa1A/X3nLj3ADc8j7m2oE5BoqoUAhx1PqjCLUglRcnI1EIOjaRww88
1nTwUPaLyMLQC/O6OIz27yjOb1mqgrZIDZaRLA3oviXFVWQJnDwyXjHVzjS4btH9
SZfdTHu3DY4uKtaCH05ry2d3koPRuu7sQrbW4jKlAS30BU30EvfwtXrj2KnWtMlM
ZpA8vsl83kwSmcDyKJmOeOncctw595YQ1Mtvv7K61WFts5WOUTz2jNO9Yp8c9+8l
aomsH1n4EqNIYrHj77ripnep4JPctX+WRiqE73r/nniABY7GMSM+/ovzWGuWVSkW
F3q2QhRltULPBL1NygVH8Uk8HIMrUvm3bd+k7o3BaX6i0Gt7emsAjRaqBRT1hLsw
1ZNI7I6iyq5wlfC3qZgWfdHbKyjlUlY+FWSOLkW1v4FjrdjtC3LsoQ86HI3QWA2A
M3cYgfHBzNdyFG7xhse6J8W+Idn1b3cAD0yYnX8ej3QhkKlX7fsUuzosCwGcLZmr
a8PCSbLpFsNze9wp7Ruiao8h/cWebSpxiaN0qWTeyz815nHyQSSWFLVK5shGChUQ
e1c0qRUYxMy3UM3VornD3itYFhKdaCtsgFOUi/lamcobXdKGHbEB8ZaY36ySSkAE
U+v8RyvNiEJ2CLyHcxPZ6bII6P5a/R8Q6/KQTQMt6/U/aRMsLJJuKu8HiqjJEY1O
VF99Cc3FjveN8qNvAZnl4cw5sHSk+2zuCrOwsOnsDo03hEtpFsF+CUzcQVtsHhZP
E0KMH/C3ddHb8RZTmn2KuTH4A7ID43EgqR0v3GWdbXNfWQBTsfC521Y2VZ+85oJq
93ZvXP9oHH+GYyOWbcxHRM0W/qhLbx2FpNUfsuofMKNcPGXdIWPOM90+CcTysWoj
URpN6YD2FBR3rfltVR7LOODmD/BouvAYfahkPVXuI9pzHQtZqgj68dFOoqrsNHqI
Ttv5ziZ8I99T3HBvtqQYw0byh31Up5jNKCfajd6JIu5DA+TXVPBA1Tat7H0+gNEk
PDS8zMDdoO1BnlKYiT5hqvCVhAk2jBbyBxkwwTRLsKZKnfZ/XZtODYtyzMIJHJXp
0OdC90WANZjsDt2RqNUsfsYhlFs2PUFtjA6ff33ETlhatYC3H6O3/Um9ABEnfrhs
BNX9DFxDmcsFPBc4r0wBDb+bXtiTIi/ogbb/3kkS/ADFzrWUttA1T/U5JtfiPyq6
deFSyJte6HGGdsEZUSWFZKqhX3PTx8/f3nG1r7bmqQlQK78PRGNArxzuvVksLbdZ
YZxZUrMVFAzW7DlqQBto0lYUlYLCXEfNm6UICEoAqjbPMCd3a2OMpBiSNmB7tipb
or6idkgEBBkqInJmc8rk/p52bBVT8SXsJfu4KdLGHOJ/P3dgltsrBDF13tZxjZNi
VXvev0iJSd4jPEThYAT6nd38d2lV+ZPk3zZASlzWiG46huwGzhB+nDJh8y4rGY3O
Is5pv4JdhPcRXaZKe5DNs84DZft+MvsuwhuwuvVtQkDfQm4Ne9peOGxHQdr6yhkR
tNAueuIDb7zr9SVvxIsj8cVnXOdJJCsZATsWJudqqCvTdee9N5QPC2Z7scPpF4l6
7vTY1/p7BMhONavf3RS+wZk8winAEAq/wsZECzPmhEsXqgJKvLCH7Ela3XUkGYFQ
te9dutH4338PHlbFFPm3X5QhBnYBewlHkvT9OWPBTu9AsBqeF65bkW+rsFTZq6Ng
sHSldgOMqOY3m1ZsUMokAsEGvs7+2qcds7kBi4z52fqETsnW5vBmgT2DjKzdn5n6
sx/EukwfOySLStU4ta9bPjC8eu7NqurLYgdz7r+IHQEwZOkqObOKLMjzhqISSYFQ
jfsrO/E65EN8uMD9NAA1t7/eWWDnRtjKILtlnlSK++vay6EPp1GH+vE+UOAFjBh4
Ke5cJ12OfbsQFFj+eAx1o5QndECCU0g71MoFT26RF4jQAAw3YZOko4mo0S96ysYB
UgKQ1bx2+N+wcFP64Cp+/HdRwrkY+Rie/+pbdLDlrX9mTMLV8Mx9hxAuceOUV2Ho
7u0FV6tHx8CPok8oNmw13dbofbUMQekDzF7EsfMxE27Zuk/pVbi8f/nvf7WlBGZa
bH10U5Y5942/fn49RS468nM1TWkx6YX2tAU/KGdglAljwD8VZFszOwr5EaTbrbkB
0qYb3FOXCPPUdJYZomLEGwEBjVmF0E+mKsiAcz7l7+jwtGATkkS/z4v77PNFq/2q
komTVSUq7y5F7DBOroDh4BykP+Jkb0BmsgaBDY+YArMPYI39hc8gq1XCo5hblZr7
2Olc3yJdVjYvNhQRx3l2hEo/bmG2N1o5YjGd/exy3+2bU4NzbOBt/Hfu8AfXfX5U
pj7AirbStZr7Gyo30Hd6Jc4ZLYu7Chm2BKxgGQDaHZd4vg8+PLglGlvTIva1zOza
+03HIdlpacNJhsWuom9rI/RuJMgnKbkUE0M5i4FlEuw+Vc4AA4nNu9CgHyNBNVat
EulGf2XipAGc/gsnyUbn8/7VZU9fHarPyV2BmijWDWBuZ8QgOM2XWd8ESfTlfMoo
m8iGTc/QzXGugK4FozVT3E6By1JZvL0Kx8/jEQnIu04G1p5QpEjckZ1cCxErhP+j
dUQEZ+ofi35QxphuUoVtD+bFSX90g9Wpo/PziKzvTXnexnOecKvbqk2tl0P9YauK
6x3fYrA0OgiDhTrLCrWSmIZNoOQUurmwx9MX0TfwTD4UohPv56vgFSLFgjM5z8/O
YYrJHP0HL73fdLFOcuB5g0KG+q4jIjWDckbG8bvVTy6pfQbQKrQPzoeUgjFm6ehP
XV+0yaXT9/nbewoprYb5fahmOGQ95azP/KVUnOhCG/22NWWDdWk9CtY3/oYsX8/5
ak2tj+115ZalFF/8VWWgHCXrMUy+6NTCS6QJsU2MFah5ZZ5gDQ7Z4t+M3bclMzvX
oZ1ZChcCn69kCZbVMd8isVAoR0RlT9iUSefeb/HnWg8LqbuHAEH4k3Q4Bb2us1/b
PkGHKuW79a/W+OZv8rCnFo8Zf2fzobV7NEpj0A4DyWwHWRKR9U/uHyJcGSvYLM/z
GIxXjZDqJLPYjFgzmBZOjh9tQUr2UYtUSGImzzbpiNyxLI4FVW/d+GvdZriSvHTs
m6TmxeGMrK+MMlG8muV3/gZPAU2apeactS1rofbLorGp/Qw3+ViIaAWSSV8VcP3p
yKtsqPDQo2jAAHjjgy1HcAjzkfVXkBvm7sdX3rUgkUjoysA1nc0x+Kb42H1hiYYv
4Iw4ekk2NGavWdWGZcM/FzL5+mh0liP7Q62txaVIbzmR49GjGC0pkDgizy+yJOQN
akjJRIJp9JOr5d3GCAgSisq+pu59uyzUmqiTCbKxk6CVEw8DkOzVlIjvnTbreM2D
qajQoT4eJKq6vTmBgvap6/BJyYbfGkLTyto9ySK6uwjWjOcYVepkx+R3vE+r0ozP
nAjh5IRMJVPARGmaCFQRXh/lzxz245VoLBnWswjHYPA4hLiHs7MNmLz9SeMTslDz
b6z8VzGK909dn6MaCdeE1svAeRKyk01vBh/OjbATjhDvIioh3tIFfPAsUc6rOCN1
IoJWimi/jQLYplgPvsLb7n2XeSAxTOkUDupj6W4V6vXQLojK4Th/V9hExKYA2EQX
9zcX/FeYsny2oSEPAZRMt6U1jfrDuQ/77Or+GRneiPlvHk3sEtPpUAj7CUQ90Kbn
QLDOtVxHw6qTbqo/wIBU/3gvYvhKPPuxXDWDKYN2Kc29kW/MIZQkWy98M1P/fswo
kAAOsonmYI/CDsSU4QCoki7sBH8t4SYiozwhHkYzxTKqSIPPOQWhYaM9ib88Qo7J
lVuBDtE0utsQgc6kV+l/EMyTWeay06/03KEBaXhQ9DuPS/Os+2QrKGjZ3LFX9KF6
Kbcjb0GmVnO9wg3NyoDnNtipM5dv9JbI077cwKVR3YDpvBcjkG+Ap6YI2qwjU1K3
cLQE7HXVEW3/+46nG0rWvcgwn8hQ/8fnlJmAG7Dqh4JizTavOdKUTIV1xDMSkawQ
yQftJrzUUIK8oobPPNq5+7JCTJikspChgEYRDCrQeth9/MkAnz9eT1yp+xuYCn27
ifoV4CZUuALkj8krxqqJz3xR8v8D7ZXePRBi7cVY8u8TDjTMFI4dfrhnNXgmkPAv
+GOEpQNHJHRJGC8bRjPdvZlF05zRVkhuhXPjjTJoCkPKoSzo86CjkWp2bqnLYG5m
1rkUyj3CjlPccZpcWJ3S4GthomqH4b2tVK9Rfgydp8cEXPxeI5GI3bYaoj/l6JQR
hLGk53t6nbpMOG+6KULmmUhTULplMLkq9pZtS7lOJKFURUovt6dYd7GAORA564EO
A1go0kH6qPw99ClxRiUyo7qCIEMhB9YTrAFTh7D8ASCk5N0uG9+4F7YggPmnZ/OH
Hpn0ibONC0sMcwbaKP+aAhwGEWqLlg+YpB2thr+HNtNLQ8JXjIf6aZy+fKZ3nnNX
YxWmLzIa2Q9aa7XywghOy67aNZpjJ/tSv9wfPrGIUU6Kw51uQ/hAMc5vnqxDqApS
wPP2XT/BmYOU/AbxFeZCTqQn4C19I7sfMp3H3zj7w7bmUmKNY+C0VOt77G1FyGCL
c02d2WPyblbazIFdQz7bAuyKukwL+LmkKS0t89AvqZYQEOg59H0PWQ7uo87B6uMc
H0eEQte2IQiA4k6v0YA2CNyc2+QrNvw08rhnUkavTya1IXDX3Zz7V15zyup2SjRr
wKFCPfqjLBN4wMbzqytPctYYRBSnan9cLe/80vz9axfUtfAw1ETybmvS2GsC7cDf
X8pqwJUEA7SntRdMmMairUQNBxOsmCcK70RRuW05XPYRVFEF7fx6/VEwBZq8WrR8
zI3ViMpNSYwcBvqfMf6YH6gVXv1cyxUtUwgxyKaAdPn0xTmtQy6/9fjcEseD1keH
38+bXQEwoHE5fFj0AAysJk7IkYgQcJV8IcQ7likYxE1LOvs6UWSV9Q5NQSNAxzra
bwuoOAnkX0vAzJ2r9CgDVKRnaj6r9uK3BqVqa3RPkfu1bv6S/BIuzCmScBMDpxco
MoN08JTff9bAqJsVMaWfhQdxJ3L66+3CrWkcjWE/EE+utCvv/LHPp1co1tRmZWa1
ciL5wqlwAinbKDZHCuBMu10tHWr77EteltaGddy64gzwzKFnh2iof3f9xoOd5A0B
+hp0mZ+6GCPzgVncr+JQbOZbLvPR5vSucr2JGSr+ZSYlH/qweHj37Ay1kxvHBGvA
9H7aGcWcRwQrK9GLKCljEhL/yGL42/QWVPrh5pEWra4XJXT7xdLqj4vmg/vnlWQ3
KMbo6RiR3oJYeWoHc34KPDOiIQdBtCIzCfmAEzwn6C1Jy86apeS9vVK57MJLeZbm
CZEkKl7WFvytIlbOiHusnuPTzKNoQmOi8NXVRQXMsxEPsjRVL1mk4zVYa9ZTz6jL
08mAb5Y49vjXk4gCB6qGf9/f/upSFx+l9M2+gDmMJ20GLcXy8XcXOEDZhh9u4MjA
A6rHmhjRNJ+9ET1aps6gDc841xVSbTam1NgeUdRR78HpB0tTN0Zo3MQFDYeu6luV
L3uFpIFB1c7Xz0WjvJD7iTK2SaSPTbKuICxBpEsYYklry3O81RgHOXsRpA4MDE9s
apcknFt4J2m+VvbqbjJ3icQ8OGTRaiU6KqXKFJUErPq+DkJCcK13Hi99nGxFo+Ne
8GkN0aICut0Sdx0sFXQxnAdeWWJOxRkTWhGiGTYj+lajbaEeLzZy0VemWZGNE45N
+xNbyXRmTDDAenl3qIi/anHHIpi1WLMrTl/xoKXaM+XjeYIbUW5Kbtg2JHcM6YPz
NeAGC4gpeoU3S5jr32h2Q22xPHO6aJA5SHDOFkFUegvDVz4cS3fXcK38SGZtJXw9
O5/xaCd+6RiDOhMPPDvBp6vX8e+SpAzn6AczA3266644p4k9s31et+wGPN/W09on
v9LPclVTULCSIqJerpjTKX7xebTtUdtjznrofANUtNn4ATFiV0JEMMEGslu4lHH9
SjsYzPa8vjDcnT5kYzjsjW4cbtih94wrEM1qYDJg2KTagMWeS+n+bXefn/9zf65H
gD9LIU167hlcJqqKVNU+3DLoCwHiiEn4NO33iZmZHYKhcN9xE9/wvQdVd0Degmav
pKzZ52DP5XYEyAi9rqORUf4pTEOoToaYN/rWdZ+v19YWLiR8IMNhdN+68VPmrjWn
Sii3FZnMCzH4TE5g14wMYT0d8KqWxzGL7tkhSgY7gyXZrNMv3jMXTKoBOOangkqP
HorK3bfxZ1llOMHEb3MvL3XPwdB0zDSM7szEA6shQK552JcSYkK129xZyKlUyePe
dsjlGFN3Se15yzgfAEGJYel0UHcL6QjSkypU1qs8HRs1Ivy1h+ZU8zfoVU7gOf8T
BCl0in6DkLdFHIy2xPY7eO4Ntb3vdeo022UBN66qlvYIBLkq+cqrcOVAY3z9vJO8
6o7HwXX/x41H4iSLyrCLGse2DeSueK9HTYQjTqjz1T7E8Q4z3j3YASG2VaZDDwSa
aggYzYwAN/Oy8qCRIMJBw3uMeSZGe/PKqmvf8h03sWPuV9ie7pamK/mrjqfp9bB5
UeOFowug9yLpyYty88LnXU0X1ZlFw4gndv4lodFkge434WSWi/syd8Z2i1B7voyx
+HEEE9hsaFZLxBsTtLPpZ64n8Sf00OenYfZgPh5oQ96r2y0kPma1SYBJhg/0W7Ol
AGRcvejlVvqYK7uIgtR2j9k7JfjcoOtxobe7oFeW1LbwAtqSqqy28fdlLK70jQQu
eU/vlpj8wy7IK/DCXd2b29qci12Yyn/3XTvEZgekvx2skSaIkKhTdG+1IljoGlRe
k4RMLw2QLCHuEimJAgkOlN8739atKRyL3fZa3TGl1wm3HOF3WBvOfVB+WQ2te0RB
8Phs2gZSWN1+Ttop5OJ7FIgbEZuWOjvkIULvmTTRwNy0Gj46tQLimfPxpHlNYmuF
nx+TTTzLif7XyIq5DRSWmQ5dOMK9b0ReVhWIunPImYOsZ8qCzNr8zkEYKD04jql3
ZckNaJsgSVM/FnVFCmbw7baYQRLod7i6wmEkJ+K4w5UCkS28ms+CDeTOGFU2+027
HhhRDpksh6BjwJ6L0HrAsFQeUYMXuIKOkQn2nLY6rOxsk2F8hiEHrrF+BywAEIge
7ljpX0aqoCw6UigL/YHpUzwGZ/JI1Uw89WRf149wThtlAN1z9VPEGVpCCO+uvxeH
ARZKyuLIbeW+0AVE4+27pS+xWTGY5wOc5WJCEltawXoNoQInSjtzsEWnJF9kNHm4
ldoTRsZEnyk/pHjNPTmym7Sdl+hwCYi0qhmadhVJpyMI+tcdayJ470134prV/xmk
hlwLOcgPIN2yllcsf20sCbi0joEe3yRE4oiOwTT2pWX1qcMGQyNKcVKB/0XTeZ9H
Un9jJLEccap4AStDeO8FR6+bTToQ5AkY6S6/TICQCBjQ+JAanO1bV6Wap7b0/nHq
gZU40WzY1YQUK8Zzlse3hImx0cFUzKxC4jD8Ucd4AfPacDSFhvXQpLTXeM474f0+
3Ue+nxlDRtCZUbDUNVdTcq5GTR+OVFN+YUAmfMZBpIznep/mCxrcqL4+t/dsNM63
hhB7yfrtgGlMvRHSG4s3YI6hiMrmhL4vdBWyLo1Vqrm6dLY+3NnQhgaKAYfRPsIp
bFaZ8btQb8ZHluxI3XNX2HqqcXaT9x9ZWOECFRajLMjmETDeS6ECjK6xVgEAVNIf
vD4OCAC6PbOQrnmHMpblykcQAMgJXYttN+B9xE690xJ4Zkot7BU8uBEbfN8JekGC
N4Wx9vrUlmKiUbjkqJMlq+zh7gzLugoN/wsKy0sVbzUTvgxYI5/eIvP0JR5u2fiX
S0oVVZeFgrTZoz2j1AgXAekirs77A5UjCdY+HfkRKaqusYIVS6NtlVzcqGnhdO6E
0H3KcG8gDEGftQiyDv79+Dj7EcjzM9nRLRAI8ekU/wnZitFAnNM+bXWG9eBIDPnc
X1OAgttUo+9/prSgBVShOprexDVQ9T1/5hjEJ7Q5nEMAP68oltb1CEDvL2FEciKe
krf037uo7nvv3QVlykD6+jziQwxG+G8UXit0L3EQY9qp06sUHHu31b9UlREfLWEw
vdFeAXAm1JbvuI6Fbo/fzv0nFqBi+/3NC3+nkAwXBR+AhoaWjINECJ94MwdV0mRj
zuPkq5IEL6phc7Uy9sXeAipCx3SQA+EvK7m3jCQFyW8JxZF8p9HTES38yXf1Ua2q
2ivYtpTEcGAIQ3NdOn3M7zUX5fe31lkS2U/DfhesBGZSHxKlAm/HTRuCpJLkoXTz
FtZj0RiOF6keg1ZBU/LYOXDNwLF/5oLrzQuWDgyju6NuiogMnExdS0MwBFZaWK/i
QSjIIX6oeZvE3t7AhA9cQTUW8L+5grh2SWbmHEwjzRnB7dlB4oBnMSfUt5o8wQZx
nDfiCD0cXsWPxm4CsNP3OJ5/BfvsM/M2jPGYPNnkvsPC7gOXTFtdYjLxLZ1MB62y
9fZcNsHkJtRjvDW4ykArgOK6bdZjUebRXofpGlYj8WfiJVRCQhB/gJE5KlzfCd7c
oep9AokW0eSSrakZ+a14nY7oQxlTx32yV1qZuL0DQwtDkjd1eTrQ1mSq7uXvlUpD
HOuWJTE2eIKLIkQ6SA8EiZ5bMVYLYgpmAyVPmglKdmTcRJ4IWYfzL6VsorrdNTGn
WZr2EXpUlISTU5wJmPy3C7DxWLPVpUvVfEadhAvphFVqmRsmJk1A9W+qLzF8tAZ1
ccbsoYOzjYksTyH5Z8ZgCrqLh20dMW8wBCv0WZzwwAZOVl2k3UUQclze6PZyMDTj
Diz7p2w9tugwxHL59a24E4XodfHHJf8VRE5WGw/C8m24wKAr/k+WPJKd7kkixm/A
nHomArpHqpLps0PUkEs9iYOtytrfCsWpQ5Hn/8tjpF4zLZkcWsiprEgcdGpPRCKp
XQkGSE53isADI2aXFRQAHXx8qU52BTAzeUd1KzMgqgYqxoUqFtNXAltvdjgg3can
jELN3uwwzcF2u8jGEEXjbrG8iEj2Ggz0pdDszM6b2qdo+KNnVIfGbYrL38m1t2Xl
O8UcwjbfGu6/pQK18K5zjTLcM2uRhH/a++um6amhTGntFw2JB5xgVFBi399SOavB
JXdKKVI2LIUKlX+ALjOaMkcPgKxo091UGD9nw9SdRqOw/hJa+PD42jzMOzHB6XUN
D9oCXhOpyPYw0JSlF21osp8PhBSEqDFYRP5BlfuHqF7wxYDfYKjd0yCXHiWbeVXD
qUtidlWv6tiEKICqNuyrfynoJQ3Ouakt0aYTkCaxqLbh3tTvPhCBHQB7Q4B+leQK
HfYvSirKfytRkxU2vuwau3tenBYvHYRUqPksf5xtKNpKA+QuLAqX4miPVA67T7UU
aZL6OcG0uLexpt3Z/2S3uCPtXalE/cccU3Bs0AQUBs6vr+cjbcmcCnZxZ8eNGuX0
31344LQulg/QZGB1gX4hJj8wKGd3tTZiu/Xqx3xVt8vNDA8Ce88Z2UL44kSJbuWu
1bLFNUEcRDdOG3D402eJ5RGeENV+nUSaj+5h704fSyp7m4wAvIsXatMvWd+DvFzZ
fQh5rgLVMO/9+AxD2DRvp/r8Vl+90gPUdjQsb+dlbdj+PZ6KtmOHdsZMATwXHg4U
RaVe1JvypHpK5YG2Hi8UPNV51h9qRfuuZvyeY3U1SQ9EZAV0nq1ytnXR2+c3h2Fw
j5v6B4qr1szOMdtLBC0IKf4nMjbrXL/J2ucFwoDaPWP0Tqyba8Emq+Bct51cw/1a
21DYUUqGz28arszvzqIue4etxN1l2ghzr8XRN8bh1ukyagZZNozhxV6OurMzlSX1
NjXitMRABIS2uWZCE+AgCyQZLb3S7LsN5FSuE+UMrk8IeHC2q5hZQYdJ4uPOEwT2
5HNgbQnUMsUQWn1PIDOCm8XNHp1SDP5XOXGai9DdzvxdvzojEW1v/OY9ytzfefzG
C8cAhYBsGSHj8XebUdtfHOyAhO1q3gOaWCuokpgxnweKx2ZYFWbZm8/LLTeYYugR
ZLVbFUhD+XE2EoheKoXEJzGqSSfcpBsC43F/A5EUT+j5tDeIera9YcnxYCH8HfN3
tLMFaVWCciCeZtgx7IvOsT5zweuKi8Dvrw1KXBAneiZVKUu9cro7FoIVW3uWHRiy
t9gVSe7Syb/iQHItB6oqiJWxZpTTWQXzxwKTn/CVJAATmR7E2Bguu9jfCL3xizbU
pnvf8Gi+DAMgT4J35tHrT/L9tIn6LmCf92XFI4XRy1SEQXIXvxPfNWaWlubOOusf
scBKrsNfOg3Mr47x+zxUcYucI/v5/OG2TSv/JYOjlfPrpmVdqHuLbvlEA/WeSRSA
k0juIy2oc+DA/ClY7XlV16DLd3abzg+BmJnIvYPTrk0qIDDTbWJNdkZ0jNBS8Kzt
LA9Vh2VodpTV04uRz+WYv9UQIqT4Hjqy8bZoiwxPrAkGg3qxMXRGILBwD/im6+md
L3lrVmVqFx4sq1//JD5v1xsyr38uGszSfCuzzdIy22630NRkLpUGpLUdGxhJwgFU
fgYh9dY1Q4/N5KdpbvgHs4CxqH0gUtZD8yrj9mdq1d1YOHBSzmDGzkoZqIv4BopH
NCI6AVcWZVkypNq1yTdHhHM5nbd487xq3fEINSB3y/RjK+tCuo8kBjmEN1KBJRo9
o4M/pjomblfXt3z/ZGRG3b34DOdNEL1XjSjwye8g/+VD/MEduW7X2TCNZFCJXF+e
1S7FOYXCubkTz/hZfA/ppHfA2EI0azw0hOUmzU6pk2z221h6gGHnAwWBWNkGEz83
lWOreLtn4UhcTEVx2xk3mH/+EPnMoJpxcbO16N/MlyPxOQWPzchDVaSmW6v9RyJa
qbii6YdmB39F52apQak4dgG3wekyoXgbtjgE9c4HNfRM7lnaRjLTxmJeIQ8nO8/R
2fuPWF/NdXjqMeChQAD2PhPKN4VtvdgMp9y831XFcaMcL2HUrAzz3HY7D6n4eOS0
oQldXN01tjpD81TkijQxMpYtcyWGdDAIsjS+NbP3j3Ct6EO2sEKLJridWs9oW9jY
vtB3DnrYTUSKmOvTISMZK4QiSnMm3bEVbbTz71VSoTMCo6l9zmTPeHYWsxZZZdSm
nLwumGG7pjs/cunQNTaG/LHoeKDp7zJ4shiXTb7kaDIy+COthkqVWNew8MciRF8h
v5n41Xl94CWVn4+nttCktxlRG23utCKqEYr+pjAuY4xBv1wfcMcbAQiVHKKLUIQs
M1ho1Cj2c5hOSKYfiwjiErd/IQs5+AtBX6ftp5t63Qcp36K2LzRtiCaB3lITi9sk
fMPaTFnIpxUCtXETO+fw8dchDE/us8mbsOSdM0GVO2A0Z+H5OVLNZbOkbcNhr9jd
3PLV7nUu09CMJ+2g3Q4bBblnpf8NsD0TgQhYvALSmM963I25zPzr8ZpOe3EMNRXe
k1eTvJBrPDRznW82fxSR+q+MuRm1fXfnoDRXJVgs8HvPHl6XUbW3a+1uZHhP4LKY
62/wHURmoRvqAC2FyDlY0UQAQgKQW6c57KULe/a6EF80JIjCkb7+q3DAbiNhs7UB
orYjZhyZA0RkRCLc9nZe0JeC2D8HOj02C6Wi9g614aLm+l/Re1myp1Ff0CRpEQWX
7cUUgpgLQwit7/q41eU5ViVu7dcnSO8myBOWF+CC+HxquuYzUDB2lHkPK6ZzaJr0
Uf6r0DkC7wA9FxKgquFfWM5bHlEZeQP33XxFc9iFyeSc74nq3Yf+VTPJulEIBZtE
15h+galmApPol+R+xq2N66MgtCPxoK564AQPSxuETxnHl2Z1BOWGOiL64zEoXXgM
zoSyrgJiLnPGea+cC2FK5XcXl4QI0ddcFP1jf33pkbLOKqPgD+WGGfGb5wJd3v2y
DrAdN4ma5haDSpjuRjCIqDeAIliEbeVY5q20whUwRjY6ypD6D6A7LdGIC7KnD2sK
49ZgrL1ijED5uY8IwdPRqmlmEt0w04dsWIb6eeuaa0Qfhzg52P49iUy7cAe8CNeV
TX6vQ48Jq5qmondw9T4/DQ4CXRevaB6TNy5WRAgCgUo6jrbo+KHL+tGup4qUQ724
jZtqHqaJPoGgL+qEYSGid4bxdl4+SZBnF3NQzv34JE4UKgnTuMDy/zrEjNUJ2LtW
0LzLOhiU0IVXPoak2hoC00zM5OdhYyJfF0fVbdilzVE1yp2Q+An758ilKVQFy9xz
pe4Et6hTyj8oeasZRvvQUA==
`pragma protect end_protected
