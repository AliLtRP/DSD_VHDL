// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:42 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JyjqDoRWNkNrqEHnpLPPPq7CvYvVPJNvIykK3jkllBrVAyNSVJfIugue3EvMO8h6
Xi3HImaTpvcc657czTp0HnH21aBFZk6HB+v7JVXaBLkvigfNlA2z0P8QSoWsVASa
zCGhNYaczZMsu6luW9rLOQHRM7Qqbjh0yRJ7MM3KCN0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25216)
RJ/wYowZuKs5K8IaNLGV6KuUAfwK3RPZbkRAQdzvvicg5F7CvC2FoxcStT9hE1vv
0Ooehq+D0pD9/0oWN3LQV6zloXuFCs0ffEwunK9I8AXVam8CSbsqXws4+46KKQWB
8k+kqhI1rIULiGJRy0ps+uz6lvLZRxF7upr+AmDAueqWpsGGiQMyKBghQVw2WcKI
GllSOi60ymvcAZo4yPrXGp2Q+t02IXZ0iL08kg4zP5pG+2MuOPAaXEJISAH+su44
evBmbFckea0wfl2tOiz8NXP9CbJRyEKIbjDFvfLbeIqY54SVN3N+Ro9DuxslA1HF
eoR4m/1cxrzh38BanK10QBaf2uIR1/xG8w21kh2TSrpUcylZLE+kAmUXw6DER64t
7u7KVC4Qk3JspEqFyNUOrrRHMDbXzrsMEjaEW6DHBUCu9DwGaj7BMHWo9bDhgliX
I02KC3WQ/VaXcxJruxsdfzTwMA6JV7T6GsHH9dYxsczHatxUcu8ILBqi6DMC5TJL
rRyc3jbtr+Bs8hDrLZOszJjnSNvnzdcrDRQKSJr1cXMYNp4LQMcB7dInmXO4ZdjL
ndNcKSp2StazkRNyu771rAXtun38RQd5lBgWiQDdMswfzARYlBhm7ZtPmTaoeSed
aZVGJQdMU166kqkPeIunRolsfGnIcoBIjy2jypacaZgdCNAI4NSxagDioKsCjVey
7l0+Y7TdjW97HOkiobjms/nwNJHFbikjLA6dPaeiIg8EXECrpNZTQ0kHYIuMGcU1
l4ZHvp0FrqtD4mAmRK/4mAgdihMvzEXtJyrbagHBe967350c1yTboi0BRu03pMh3
9dlzJFHpfjjc6eWScA69DKsY7gm12UoTfCfQkPLaT3GN3/u+txB9WTgqZJeT8SJe
dCng/bBLyN8NB52TQ3x5txMHiLMz861iRLbXJ+fvQPGn9RDKnkrty3hpMVN6FwZO
1FqqhPq1U+5jPhRsZUnSB8AnJSysIXLJ5Vw5fE9lgCLYWdytEa378Ehm/V+pzn26
zrZIFrrzngxijt3rrzcOgKgOJ4JGFreKxjTLgXWIKxnPIt9YYAzv2/f4Qv0imEF/
HZjwtVd9qo+BeB5338HXySxWz7vriHzmiCih6VY9VUH98hvws+jostKta5Z6YYVH
d729Rxxx62+JkFXWBSC1btGx2hQP43vnAwiYR7wyfD10c3gfTXZpN9eBgXkpo06z
9sjNiRceh3C7pVJNmFKgoQBVWqJEoPIdimllAYtg71UPArDd/i/NvLddE2OPKdli
ZmdkR7nQcH/cOeYkWkJB4LT5AFt6mrK6Afc0sL6c0F2PclXRa2lQO8u2Md2vONWk
FNAwbleZavLO/NVoytW9d46c9TuNsQ7NsxfZgFI97QI0foeyQR+7YfrkF0kFZOcU
9s9PDlTeYJo5ybppJ1NLuk4Ar0aengaxkm1WCGfw4FRiFsCyQmEeuc0kDMgbwI9A
1VYB3CvFU5MC50anOjVVue8Fy5la1M9Hh2wPLGRttLal9739HMJTl1IvCyMNxpjn
mqgnt4tMpIYumMOVQRBTtgkO8QP/hMmrnUfpazPdE4nPu1mMFSGuhXdtvrzQyZnF
dEQvY8TAS+3tAWvGyPW0re1c1NUsgJ9PfK3yVJOLcHrhleczwWOtIP90x7ZE47Ft
R+L8p9oRrvBzYcMKG/gEeyFuSuE/CdyTAMmS/R0wb/hyfDWl9Trq6TITqvi2TmsY
JHIABphtAlYbPCkkRVicSKqT0D9JrMHOWSXopa/Tz3tSqKMCjulGuRkkm/PDI10l
T/8VgmlOyI1ez6D+XNTdz3Q9OnKupYc/e09h2YqpvO6WjGzcFP2mFLQ6zZseawgg
pCYkDYEmc8jckjNnxNZyWjrkU4LE7IKPrgRwOXO+Spc3LnOtwmYmhBjq6emG6XM+
bjAkxuN/DpcWpsZnGjmz9kUumo1fkBmN4m2/tsfyHu+wErTScvF1pXWfXkeyaUpu
ekDH4mW9REKFd6aNGT872qTngDPrAddLvIcIPCb5Q3BXz8laO/qnJ0nebG9A3OfJ
lA6y5lCyiWsyfZVziFUSZtlnUmGwTCRHHmCumwygDpY15nmGcfAvx3vd6bmB+tcA
goV64l8mDKa7PsJRtAQ3UYsw0bm0KiasVCASZrMB5P27B+pcQDjxHmuIBamckXPt
q8I3Wej9P38DwW7gbXnv2ene1IShyZCx0Is9a04gxdvCg7yR1g3jn/surDzOBiUZ
55PROUyCwtSEKQ53tXJTDNsNUuv6HvQ9PSVPaknY2Itn4F/sZxUes346MvMEvnWH
CXGa/+NcQqcx/KKYMeera6+moLQBTjup/t67dgaV5EGLwMe4qhq4z92MqWD7y1E6
VLTsA4SpNT8xsTUEsmuRk//9YAcFHDi0t23voO2afHYlQF3Fe0UrG08ZprCex+w5
wuhB4KRqn5M9xUXaPkr1F+Iv0j3q+ZanK+Sb2copgxVeJSPe9F6jXEsKJiOWAJcj
IwZO8qXsKPOs39l5wjH1kjeb0myfFblogd+7I/l/xEEOYXzYMkNhYL//XHcpqyXO
bCTVyFQ69w8omSSbbfWyhQvukQeQjX+pOeWn/IGOExa5nl1vvqRlakfjVX81Un7O
sIvbvC31M7ivvAtFKMpsaW1KXh/Yk3yhWe/to4oD/tHNM8piYpfKv6RZlsZuUSxT
xj7+B5HyuzeIQKTbc7d33oDzfCY1ye/szlV0k1NqNicMDnSNJ43c9GYGvnGkezTI
BN3LTvtlTOl5PPZ2zmZvIpsesxdOaIOmMwd8GLMJ2XtNQHwRwAVJiFPfcUsxDUEI
P3KOsmpO1iU+m52/jVwJqOg8JiXRn4JTnAqWGqEPdbHhh+cerUDhBSEik5uTki1T
wPd8sar5qOR10tRv4EG6T0QRFLlDUJzLZ+fN0pQ+1VpcC+EPJCzEkk6xyfRf9EYf
DPxi+oT9vXiSidFCuG/A2Etkcrmiz2czg+DbaoaCuE7ue3AeGBtQvnDVyWS9mLLu
tfEKo4F5aq89Q56Cq/sZw2rWTvE5se8tJpVqQqSD7u3D0ikJYDj0As0mRHeQVBDi
2wTwnJQyAH9VkFTyhMaCo7dLQcNTtGE2MipPwQKwbtM2c1vfTRiA3cFCvCc10fzC
ARXSWqf/H7ak/PqLy2pnJ2NEd0HdfygwbYVcd8F/gtwd4cu7expZbHGtSQq3JeVT
ksZhcrNZgGcN7evEELbiOX5FGoP4z3zIIQqGi4zpqmvO3ymNUKpWYNhVqQF3ZWpc
oXbWKLE1/FjX11c4vyi0ntaQExFDgS8vP4FJRKnCyyvV2Cb5mbTBsWqyXvx0XzP0
7DoO6BIKjC0aCT2pMpuTP4uwxSQ+LXxOfSAhHS1xbPWKwyuMKj2D0HVg0TSclGzs
yTIL1WNQR+0meMesHHjl9haoZwKzVR8iKnE3mtrTkZKQukkLWTAmXdQfXMiLFBju
tZaVxUgrpx3wWqc92jLMr+ov8lni3aWdZMq6VSZEJ9DXQKba7ko25gg4yA06iyoq
UbK0/iRBdLg4vPtkZaT067qs4EsoXgoIrAwmRNypW4e4OLGUIodkaM+DDEbk6ibS
w9AKG73KSZpuiF7wrVo9asIW0rVzr0Kj3PyNgOP9rAxgE8A+qxr5b3+RgcD1+yNF
OeU0Kk11tKPoOULn/8M7quG0qO57Ob/ZyjUR35J+Hn/i/ZLpac4CeqsvBkoccv84
t6eA2klm5aFga+d4fCfHuO40+sy+ypkzl38zkUVj1a+mAuLw7nnnbPXb6+5vRtoC
ml5NyGjKd0XY8CoU+ekT57w89DiVK8eaHAqv5Ln5m65D2AS0UTJvf4zFZ+nF9chN
OVZFMZR2WZJzB23rXTyWT3hNKA1PoYD+nR2D3XkMmmpL4zrVbmwULSmxqrvjQANS
apxE5l+35P7nunIy5vAYwpOlGrpvNb8FOTxRIjw6yhMw5lgAh95rYenXZPhY3Mec
0YScodn9nLKLVd8y9/W/ZzUkA6f5NrT30h2HNFPS0cIhQMj92CHJ53tHNPGX9d37
WktR/bd16mh3BgfCcR7dRDLs/kE8Pkd5OkeVoa8TKVImfR8qTSDSu2JIznK6FjvN
Z85koNSuWhFv1DIDAt7qgA/RM6GS81bc0KkrvFJv8BA30T7R5CPoOBNJT9qA6S6t
LL87y1W/NSlisoBaHIEIndupEOjRPmIkvSzpxAup5oa8yyj/B88W3r0U35O5lSTq
uZPJWrusetKvl2D+D0JlcXT6NVfCBe7iZ2u/bNUedFHhDYN/Tf3x0sI1+U4cvgb6
6k1L5yExweLiKOWEa1crdLMZEuOvazE2x+R2VEhh25qyK3yK3JR9XsSWok20nsMe
KbqFLzD46Mgp5vH65yfLMWbs0+wIpUxzFf8wWV/0j09SUvHQdbZMd0VDtxoKoWEN
S8TwXj4G58UaNcAwvjFkjUV0Pj90mClM96ir3n2ToXETFhbBS4ti+DAcshgc1VCn
AGiOnn5ZpchBpIcjFjaLfmm4FrkIfdEkcaSvQdqh0+K2creayD5FrjaOzTdhjvuA
r71V4TZhbLRGLHwem/tnr5b8r1gIStxIzf4qYGznqZ+YDTXjPEtS7nIHG7guJw2C
xqJp0ktDlWTBBfeCGaQQnXGzjC1LCIwHclSVuoKvZHiTrT62WuI5nSR2jNot8iUP
lHei4Y4GPcKdz6jSNGSrKLwZp4FYa71hADyzCpDpwmvuQCCz9JNqL9dnLJRXjhBg
360MSWqS8fbe5XUirPVc2F4VpkZ7OWKddiDGasJUWnjBEMYBp0B5RRW/j01cH8xk
dIjfurg4iIT6fUGY4qyEr7r9lBJUtyNEpmkT5FcPDq/SxR+mFcDGP29jjPx2K8sG
CFpTu6RJTcSDV6qui5PZTJWsjqUZxYiOLAtpJpuByC+VYrmBZ+iE3Mhka64ZCXdO
z86yWzZ9SsH13i0ymhNYJPmCJmRBaDK6kwjZPW4/nQluaMmXGm3zrhAzaeeGf2H0
UdyIpLaOO1Ow6hfrxKCKZXOU6ZAzrt1JgG9WWTDuCc9bhz36E29gPv3YdPT6tYNw
D+mSOnDjuOommv85OvFHvLr7UO2fv+YdAxcAO0hs6pfBGAl7EaCgV8seB+V/sTbB
NCKexbfjJd9mDNkM2tM6uBbifGTYy9dVh/tQfGYs0JbIDqXP9Dq7V7IfTHkGqo3W
uTjgReS6gCz7aewtm6loHntWOiauXAi+nMylLoApADHRKG+h92q2H+eXHukRKC7t
taA/6lB1rEFUjLFc3vAsPmfWF9QfRzBVU850YVszAQGeHfbzanIaqk8ErvGX8Cfb
mtVnz2VRX3cG2vejqQ5cH/MbJE/kV98QmcxkD/4vcwAftZR7Ymn+gvQbvoobGSc5
78FBmg3ckhWvKMG+Ply8M9YypBiCeNlNWTqB/5mDwbqTpC9LNouA5KKLqW+J1wS4
q4bamocFJnOhez5IwzPmxk0EPwwoGvHvNG6qj96tbKWm4M6kfQnf3Z+w9h+Ox+DX
NoWm3DWAOYr0OkP9vVPrRxGRwIIKhwj0xt/o4FB9mADWR3flmcSLerkOnEut3EtG
5MHfGAgwHB7kicrSkvoBQvhYvOIBkX/8TfqLYoO4ybpD71i+LhkcZrD9CEj2ouvZ
RAiU8v18kVXy/TXndG22N1smkd8TaXLMIg1NzdOn5NBFpxSEiusN2z0r0AhK3v3B
Hyrs1E0rFWlrPHLSDD9Qgto3lr8kxVLw87cPXa/XAP2NeTv8TgIpepr4eAjPcXPD
HMUEUfalHeN5C+VwKo6r7z350odAxD6tH8D3GKvydQ/n/8m2bChuMq//HvZS100k
LnSsoiQG8isVcgsRfDXM2McdJA6qTatDgpsDMMiLAcIiVBX44iGxVbZ0zSQEku9w
DxsR+SVzI8l/BwKASHbLQKH9kjsXGZwPViI7n6i4r+2/0C8iPTCEJby5lUwHCo1s
wuvZflCkNAbvJDNe6jP+RsYZU1lzWOykZJ40IkhABrWU7zODos1p4cWo5DQYgSdt
5sW3I+/lnYv+5nAQu1P7WHHznwncXqavNwQEaesDUfYq8sWGLtvZITD7VnZUN1br
SwfG7qWJSGXlDJ34odvmQYNT32WItfeMwe3S8WEoYLadSNf3nzHXaMZYwFctRGcu
KnKO14K3ouITJXbcBM04mj2S+deDoMi1fYve/vKMdbC8tJM992HOZ1rXmUN2HW7W
hTglKmSOx5Hf/wL/nq+G3V6nst1p1ijCJBddQFhaxZ7pzRqgZIGqsJKBDYvm9n6F
VLhQXvo9V2SmbmDuW2HWE7wgptdAr5I4skdOsJqVNdW7d4SSncuZwhUqgfqsRmY3
nUQJudorF5GxJeQxrY/aYkaJeqTkmjWAF9EsItWoAr5buZPRfcCvfabHdBibhFpZ
I7DqRyqAbQJ0hnsF1z/2W8KMJOo+5tnG5cRt0zwNJ4lrOgkqTZu0Y6DoFrAFByt7
HJD5Uwwu8JBY/UP9YXGFTcQr5OEiuo9z8n/SvCLN/9VQgSksI/zhYzGaz2porBUk
rBxyqwUh+V/8DgE7AzorDDKHnl2W5t7Xs26a21JpDqDJSzn0lhmXUC82p/JFPwJp
BwcHZbrU68Hh26WStNGt+U13/HW/OrWL1qGiOdVjVQ7i/Sx+XEEbv/7AhL3AahPF
W28eFtnBfN5/dZyNYEvtlUO716EzHIybAE/NbZIAG/WgEAdnN+C04Di+N+ZCACXQ
iBejhLHzB7D+0fCboPOSRXGcJbr306nQSDzx/WzDxPJYYQtIhCnHk1zb3Wx2RU1K
5Bh/tzs11kd77C+EBDsb0gnK9QpOBvKeI/D6sPzPWpSbiUrKSeeVidEXgdwRqtzc
nAgjxUnOGG43M/56uOFrmxglzpBUI7FhJwNqZDQEVqQMt1RKJgrP8tAHssYX7A6Q
xxIO+zxWd2GUcU7rUruTECX23Jp3Rp0kXRFPDM4syw5AODhBTNzZUAmQ/PYxA6Ig
Tc3qKtx2msQxR9GF71rrCgEjZqxeWQnzK2ApKfAd4Nv5WnnN6L9ngCCANp/A8l60
cn9wDcD1d4uPo6T0EFUgKdJQP8Eg+W0Z10lOpaCC+nna+0QI3DnlsQkEV+aRy87o
1i9URbC2AOKQUzKt2NH+8mC44uoesSC6t6SDLqzFuOGSuv9ZaY8amw3mj8L7UG77
aECbmeNT3lRmDPuMp05NfOqjpnmAVDXc80nSizf+bB3tkBB5Vw7snKAYNzcvk/tH
HxhJCUFj/vMFNcq+okAqonalAP4++7PkOjhBJfkkpQ7E5VASgdkCPb9569bDKerB
mcChqgGPDNaJSQJuJBtMcp6q5IVhNwdxhaKItWu9g1IkfZXF2Fbqrznck8QlBJhD
g7pKoz44hwXuNuUAuCVlIe7TlR07B1/0vhiV9rs0h+lt7EEa3LOOC2vdXuNBRK4O
Hakfbg+2uCA15h2MMGM9COhY+jX3qZjg4pEHsehrTaYlhKMVsU7WT5UfQwJRio9G
G7bQNbWM4oV2gyR3NZyJxope2uaPvBgvY0D9NJSRMHcDzuXRtEVQ0HN6n+sS0rab
xFxEzHiHwJ9vjKSj6tEq1PFiJBgmPs+ooUwhWkBIgPzZF4j8hL1WjyduX+7cw7DM
pkqRDRP0khY4bkphwWyNaAGJnnBhqxxVtsxLNDpP4b5CcnDtB2bn6Ij5VDkrqA0g
spIQ6qTRZ/aDFhxTzKYYWng95Yf0yW57UsdW1H3pHdO4/CsTxX4jZ3fz0zo1kn2w
LiqRYwt8IRUzHZwB4Jb7UylyyMyk61Kkk2ren5mJiWGLEGV6+It8ga8oWnbcsaA1
kxPYpkp4BywJCMYTZKBrnIopDkhmSHSwJbS0zqdD1rH0Weg93DyASX/i6/1vHSuG
BG2BQfLYAr3I3BehiFqUAB3bvRC7nPQHIlthnMSvDGdioGAfzsWlyX0FhwPnQk5N
yaXkU9cMoSD2Jx4NYBYxQi7qL8EdnPXkhiq/JVz/61PEwZTocB4ZBIE8BRYBUsRB
0d8WxmaW/CDOEFsIhgWSdhL9KYzTyaXKapZp1Lhbkzdc5+Pc3qyk08JS+TlpAnKH
LNdq0eoX29CTBB1JLtobIqVM0/T96BG9qlkvn5N0EebLJL+HADD/p1bpoVgCp2PX
4w/SMCwlBXVjkj7kmGNtZL9SvdSPpdB0RIFTq1C5oaMuKDCE5mxenYwWPlQ52jLM
gxSFcrNPnzKwvuwuu2/DpO/Gi50IFYbs3yv8MsJbhO80ZJdhNwa8J9Jep5KxXjtr
D4QvRjzhltmB/v1asQQRPl0J9Pn5Ki8zKyYkWOj/idml99z+Nw8eJOqwsTu0af53
uvFN4yYzBbsHABpNTMUZP8PtYgk/3rkc6weG9vGaFVYKfinc6llfprHCGjqzEAwV
9yRDvtqRD6gb0fcPf+KAPdbCRyWqX2myLOZacBH3iiJi77X88jJTV56oX7gdRp5P
uPJMinD769gldla9tXIMFZVjZUGSj2a43iPoetZQl+6wyqdUaX8Rrk7gFJv3X1I4
xjQq1IjXUkuT1UX3wiiRTgiwEPhNwAvOB94LctvwNcgZ2qKf/K0mbUaNfHtsGvri
Jp+nkiEWnRTjKBjtec8x5d5dEEwgmbGX8ih97uM7mQZ7FIUgdeA4yt8Y7XxQthAr
3gojDkx+A0Jw8z2m4+Dfm7mQyx+eu3QAaT/06tC1gPxJhrFjUd9qxxj3plD9mFzj
bQQNh7UWB56/Im8eKhv06YX1eqOCNPZOOTp30m9DksYSp4yiConklFGEWVOYlqMg
z4WHCal41U0/B7ynhZJ54Vb2yI2KFj7HU+/45FLzFpCT0DBLhefF+9bquPfqgSlB
VM79XtgaBZ00HDusy6XHeQmTjuI3U7a1HCVffGg1y0l2BECnivlOG/WLplj9ovrr
259/4S07rI7PswKpXQnUO/MxSpUyioxH+n47JwBXERmv8KHCIe6PnlHmngqtEsib
VQelqVKvkxQ08XYnZp8tBJ0Q8JbyCUClutmKsUGb886ucUTkYqYAO4eQ2lwUBkEy
NIxrZBzYmL7LZFfdeDGg//1ZI5K4h4UhwU2xkZyajvc/dX0rqlqfmqQmyyAELn5H
QwosW04Bg4JvkXOxmoc/anMdXtruOgiQW5TnBpPlJRoE/C90bjBkwJpDGCjET1Tw
4ZzyPKuclbJQvIOZAeN0UuOSLlEmVRsplyPxKbN2vSyAYT3l30IDap7o6v67HKpB
LBusw/uRabmQJWp65+I0V+bNjoLcPY+at59lTWlfvAygZ/1b51bTzDin1EiG4Br9
N/rpOSrFxYqJdzQl2M1PCtN3Tibju27VLq0nAU2z1IqcACdZUxTjXp4xUlETCZ3D
HXhCHQ+vjeYvlY9N3rRFZOOQivFngccS/8SvCMbT40otSskzp5cGhrfy3GFGAsYU
p9jBAdoH/gqqGmRJpmGzF5ZKxpBKkD4jDGSkcdgiLHruu7hYGSjBf72FInhZrxWX
ikz8Qib8xdLpfHzx1Dkj8eX3yEpB38nqIzHMqX+99xPAGXzQVEAuHr8q2JnOP5+n
7HdbP5bMW39VNsdjkzcS1eqjoQuf8OftoXoPV7ss2YS2uYBGGZeAJO6apws+s4Ot
QGJGfFWiuFJkmXgqgLQbYEHD7gMUdWON2ai7wr17czT5q4tGZEzXowwo8+ayMmhq
adqPr8KCFg1GcUAKV2qEe7Ry9asHkWH1zGk6UTBlvDJehxpWSN+wsuZ5dTtxPhIu
goNfJnQ5eeOjoDegXtBbSIYJx0Qm0FN2w/OMXcHUZsQqOh4PBCtqgAWXeUHRmWUT
WD3OtanMqJwaO1lh5qjMEYLA3Oj9PeYyyZvX2MnDtimDw+VOkLmiT4Q0GdwJvYO9
BNRmFHmqBu5P+h7JY1xF5rrjtEbwckJ7OvrP6QiPG+WnW98e9kijgay2jsI19fi8
U8f+xA5fLCPSm7euT2uivbTaER1jVIC/UEd0+tcQoi9RS4cBxSX6GPm4gG5pUHB7
9rrMLbeerg7krnvIWFeiFd0o0PP/GZq/Dv5qVxcKiJk3TteobzNXbuzRfO9R8ymU
tnDR2owahMxeflVnsUpKJuDs5Cyu81iyMu2S+ki2qwgMPpXBIN27+JLq1+Gbo05e
rJlcLDYi5TM5w04PiJxV6Bzg7pn+Z+ewUkOvA3TYnK/chmGzKvp/Pa1hFH/KQPex
tgtPLQOPSPaC4rUJQRjiKBfmhpJhMouItQZ9eqG/U6uJqEXABwsvl0BFI1ypFaoe
CChEvjm2qKcjnhziBGRea0jJblsuamFJmsEeEtZAn4HwP/esRgfmfzjWt2isjZoP
r5fDHBMTWm/InsG/0pWzUI9fd1U6q4hX8PyFpAHe4+ikmMSNXIl5uv9iFLwSgH/f
h07oq/WnqB09A/Ve/DwKclxjhF0EmrLb7Ca6jBipZphlV/ZjSiwkf8iDRxE9ZatU
rNi7NqnInWu9YNI8AeOQhFHuVJb3IBczWOYJL7WG9txIreGaWcFNUslO4Ra7qyQS
2Z0NofhB7bgNx1aXUgfoLZnabDlVnX0llXAGb7e6KqTgNMucQK4lwhfAPd/t6J/p
r2FDLqGAXOd3nld+Yw7XRPNXihCfS5d4jYNKRkcndiVteyWlxmTuy+P5ILxGwf+h
PZIKKzlYjCbJYde/EpUKxcvWKG9OjdBJjIHdzEVB8KCfke9gQM4gWUXBEr2qBUIb
A2DIL396jftHNJS/Yut4Rv80slopZMXbLU4ugq+P+wVQaiRk25kh5kZDBjzLy1wi
lqn1lzqmcObSR4Vg+LW4wXqv5waAqJtVlAlx0KKC6dSqcEscREg//10Fzs+/7nP6
KOjWw9d2Uitj1WGjnVAVGBRcLCYID2GWRZh978EwfzG1fD6Pja6S60XAMciFhnoM
+fRMrG5aKhCRXA4xs8imeOwajWszf2jISyQXqGKRd9MB6IjedO5OkRB/sRsJnr7b
sPG84c8FqQkp7FB2hcVPCwtGFnvd1Pbnug5JAeRuUFvi7GWeKG185Grs6vIc0bNn
3Mor3AkD+/Iv5zorXLe1uhF72rFZsiHFWQYr4kr8LS6teM1gF97sHbP8DnWQlrpE
W74uXWrSPJ7ShAYm6LzXwjeVA7m7VW5dcyMXTmAg0n6pNJSu55y5g1XbiiSBCL32
9e/T82LpX7nP9fcVY0wklOGiBZDhc0wj/KMi6RBmAnWnG2+SvXjrHVOmdqDYVIPx
vIF0s5FTY0Tr1doXt4LYJbXGZt/6XCc8fpg3jcmidMyXan5EkGBaCAFlDqy/PlVR
plSuQsvdB62cemudYUDW04WfKb7g02MvZ5mqlAoxJBty04i0CRws1nal9G74SpUX
7bq9KdHWHDpCqjejOvMyENBqR8p5ORufubk/s6xYG23YeTrkmnbZ4xIEndbHVz00
5iW7Ki/P2cba1av8/QsgllilEGmkyLIU2adrgxbyLZ00TtP6AeJM1tsVIE2Bl94n
rdUKj0itUEy1KCbSba7en8SPb3y7aHjvBzmmlESC/7nBZmW/IQ5Wa3Pp/6G2NB/+
++hBfWM8poutZMQ2nm/6pQu1gp4cUGoCgfCihxB66odx317kY4e3dwBhzYaxWP8W
M3sXFY9AXAcwBYi+JepqesSVh/WSAL6+BB7TacuAIl4dB8mDROeR17pQgGIT3R6r
BKlFQBgntKgz9p70g63xjhXC+4NpmmiWDpVrGYAJkaGfftLmvLU3HX/DuDMNTTgV
Nofx8FHUEjnqVCP5IcvwhzzTYcfa9STJbvxO0Y6ZNPnCe61Og+SPvFXD2sGdxxjB
+6fy1JP83Zza05ZdEA3i6Kn5GHmsX+bcaevp+OjqbqkDn7GMwe/Hnt+5CrBjR5IN
8PqBJ9K2YhBBm9zy8irfYGYbusj2D+W9NqBNaPWiCfbTzW0ca1TPQAdiiHACJqrD
FSThpkFGh/JYjQi89F6bodqZ3EvMv7r0ikOLnRSjOuWrrUlLWnDmYJ7f5QIKSe6Q
7/Zm+N+rEwCP7NwRHOBJV929brfmj1SfWsMbayU1wlz6Eozn3djgbEnvaH9GOWag
fLcNO99FPvmGXYOcXxxm3J1m3JFxFDCdC8ASEh9w83LS2ffN2+AvRjT62QrTwVDh
Bf5/s9dRar5OmnN+FpvdGMVT5P9Ok80r715dA51VFh+mMQIfTiXAtaBIdenOIQsa
dnWAoez3lgTsW8368PBxCTaoBw8IkXSZvn3Uo9Ftq6FXEGtdP+HDROOVcKkDupWL
j7iaU6+SVx4xe2hxs0zWaRqhQm0ON8vTZ3wNNwCWpNdENGuAPM+sQI2VGEko2vPx
zPPnNs7rr0uaFWm7I3GZBaKL7/eo9ZIHYi6y65Onr0Jub4vjgwbHnJ8kq9F6e12W
sLOQKj1kH3aN1xiBjzTF8PxJosNrHdy0RsilM8B9JFzxx/Y1H7q+S0B2QLObtDYJ
37+mri0lxtOdp02IB1QkZNzU/puUhvDpTut81WaTNnBeNn/RZF46jsXwhnDufSGC
oTN/wca9bT0qLZ6qFWhwZpT+7E2qRPFdrMYYJ/YA6ARavxMmg5fPQAORxE24XJMv
P1Ljlu+AwnK/07Gr+Sdu57wOFeQu2hFJ8s+0EzjbB+GIVO3WbJHBjIeHvbQXHT9F
xuxT6yi1QckgZL/spwKxdiNnbtNrpQ8VVSteB1+gcdxSyorLqtDmxpNTRxmi3BRu
PvdIL5Jn0IHqOZ9dJWkEDfQdqIegk86CP0yG1GDURv26QRwHhjSv10IdzhIqu6os
uMW9IziA6D5veZ4o1kdYs0LIOhMKFtdcYq3CR2IvW7Unwj4QY0asY8E6S+yvQFYp
RVyrEeb+7Vr335+ypdgsoO0hRVF3tRJaPh5NRGQ7EN5/kNKxpc2N3wNW02Gbbpwh
pECFmmwAV/u6FczaJ+2yjkdBzsYEcpig/dLIEBsZkpocLw4AC5oWFRhOxScGdY4P
cAHHagRU11CDgy6L5YNR2LNZDRXJv8YIBSzUViHcNtIbo4zt84uuLq+7Xnynvypf
gxVZ9+SZbpLF8nVUOTA9yGbOE3ZIErOQMOnpBNOZiTEb7BMJR1f5f4wu0BkVtsL9
mCyLjyYJ64sNLvfcMOnl8gSMWCLPla8jK7L/WX8Sisu/5hQRhs7Cft4JafF95Mnd
iJakckPf4N/d3hoDVKnZFypqTOD0M49+Xjp+3FZ5CqnlLqn5rIWu8uNf/7szDFn4
p7WlTjweS0wuB97HVROeC+15IeH4Dnxw6HVNRdug4qznzpDs1SsDuRVb7ge4DBEn
uWofzbxCtZaGSjaaYl9hfL4iu5YXUFrmqdpA8HCIEhHxc6e91iSe5krUQiKekmJO
uhhQSIjm5Hu6/lsU6KFbtsEEbLp83Fjw/utfKstW9PhETrCbWq04UKgFzuDGUCxX
HtvKYPtP8BxTxQyCuibdNwZ5HpN+Sd7pyE6TdebboeLGMpOytv83fg0s2/Mkc6Xv
bM9OmSE0h5oJ9e+QHNiC1HrjrekuLjlXeKfWpdyJvMhCIyT7Ru6FA9zvUALpTJXp
J02YqVdVDBYKHYxfz58HD/qUk4mC+qL9sIaiq5m41kcEO+yAL/ZuKax+EFViqARA
5P3zWY5Spf6dMop5EB6+XB+PBbmvZZjPx/aLoze43d2Qh+U1yfgK4qCf1EC3fTeT
9EQqZAeDBvy0rE+MaXEQu8NR6MXMgRe/CUJ+rVBGQNQvjasUiWxvsPFzFFZtOnM8
8hfD4/KWfRl9uXBwiCdX0pgXrbDCxMsCyfZzYyEO3Z4TouoBAtLipYg87Ob1uqAy
0OI45YfAnz2BniMrPZ0bEyslgm3hhZsIpOFEu8xrCcBP8r5gBUKA+claUaYBu0qe
Q/Y24MaEg9u73+XEgZMXypQSlXH2m/CfMAosAmqATyC2Uihnh5EOhh9RXyH+xt0E
26zTG3jjHDmx22NSBTCQ3wn1JarH9rmHfhO73dBngCGpN2A3AW7SwenXXvx8bloM
VVYOPk+8grqlkN44QPNWbWY8DV/XqEElVDC25cUKFp4/mIl8aZKKeq6vL4rVVfDv
mojrztdL6pw2Y65NQQOduaH9j/8gvkgMO5ExvIo8cRijUIaZIdfrkB4CuZZ8DJtY
ZsydK6V/F2vX69GW/IxBPTTPmS3jjxuRDLS6uIeBfjYAccBLzmhLd9h9C7O7lcaw
7AT6Bow4rTTv77fclQGcTmO55j62VJaOoIx4aRJ60C5XKZNrAOyWFeWRB4+uA/K7
sWJtgsOGuqSLWdHZqEL6ClIyCm3UsGlR6ca+zF3m9cUBkYtdeLubYj2BEfM5stbn
OSVG7CFQVcp/oPML7u/tp+MsWPwGjO5RBSV8Xi8xWWLgdm5MUgp7lSZlXHxnS4PD
e2Ch6jcBVj2RaxV3mGopUEac7z3dRkKkpGU9teLXIPyXBc7lgaebvp9tfmxlLmsl
HmVmewUrXVGkmavx/OBcoPZsrDf0orczrSXvk0sJSrb5O4RKCbg2+ym4xppdKSG7
C8dLuIO3nJdSC64D+r97I58GRJSCf0uom6apzr/UP6a5FkucD+3cPfKbu156hAXU
tW8PWi8IuKCr6WQnXu8pzsaFeG6+V+FtSS9UH7+R6zgleDhUQd1BYvOzaJNcCbmj
S/4PaULKMR1VDGYPmZbsXsFtsb2oMDtHYkIs5xc/f5TBCN83M0sc3mhaU7ELlA6h
EEmQJesFM+0a79jFIX1rcfRO3sKGHRzZTkHX4iKa+fwWvqwnoY1CMAemV+OqhU39
3NTQYLu2p9gX9lxkXZHfpQkyW15980Qqzlnk1heJb4MnFK7o7rbTfZrdCBGphPvL
BnyBBq8dFAqO9XUCnYP9bHPowk1CU31ifx0h1ScDiITxMilIwUx0+tDcJOYvfWFX
QNwU3SibFzRqa95iostzm4vi8fy3tFEiqLcNTiMvIvz4tUZwyB1DxjdOJNrBBHE1
3f/9+wqZbvt7c4oww8dF19qKLoUPxzRQBgeWDeoUTNoE8QW2hwEiOv3eyX9XPoph
/4mqbWnnGh+zzbA3UTEco3Myb8e46f6cS6fRVKKYXaB+L/wpGExQnDOV+O4tvVfk
D3x6nXMYiZT2n5aB27GvCb6UAGldgtAvenBTcZOxiSw7ijTLZRjrXgsuhrP3+J/2
2BuMpVx1OUhDNrbs+ZK4L/yfcnP2M/9dUwXVaay7IcDqZWiVIxd02g6F5VV7G3kb
FgPPGEGf7bm+lHGyKqsDEI17MUzxRqVArykhpenvDN0I/ioXNz7tl3S0WVPKlKV7
+RxqS/5+L19pSTjr9/eS+muh/QmSnHuGmv/km2qJ2UdXIvFh3KxawVcBUW3ybWBY
7RTbGiCu7bSfiru/vhHvvDuRDestnN98jhWRakS8F93/hzRrQS7wDShdzw0u3K/U
+bChPfzI7V6KA3M9qRjmNHlMMx8WhVosTpQP7Zhby3JBk9RSCRkm2oo3TYM79kHH
iLFLTiqV2QPiVv3mF0m0SoeGxEfON/J7JTc42A6+VkF92LDRybPpdVljuHsOtsAV
M7+lTU5q/+Czrh8as68n/PwrZz07+rUPLUJJKYyl2sR9Trstne9Z+iUl/xPY9U4M
gj5brKX7Q5WIIiPsQBwLZdsiPxFjKpvTXtWdiNT+GseuUyl2JTG5TsXYhAjlbmZZ
kyARsEzpyXQhdzN53XmqvAwwerHi8e/v4nRIgTmEEyhhotEN0xmpzhIx0fZi9gCg
67OGvV4+Iko4NDQSuuGmyP/FLDBK+0weLnK+reWmmN1inbOhbUMFVCnFO9j3svFZ
TfSGUt6uxN4FpAZywvwi5YKyMpWQEZ5NlnJ0qQh1q+C0Ul6SL/TVzaMO1VXFu9yV
LRt4zSTeGu9o8b1JGOFNBGGckXtVTJ9PCA5vXuQIc7bjxGQb4WOLg3KFOzVGch+F
8lwtf5XFTLD8Yhv4nQNq1Mv2c+QFLbo60k0HKjJr2aksi7rnV8rJvHhdj2LhklxR
djX+OtINuXl1KVYfXDmvhxG5i0GSOCXy3wQ4eM0Q23FSi/4/EUeIUXOx8xb3BmYz
SCQPXanOhYt5eKfwcI7+O2ubLJI+55hkVkn2lKPIIAeyEq843EMSY+b+ldd1ccDL
/UqmFruHFDKUdwUQrdMjfOVOwrso4mEdIgagHcaodhiJ8b4bTmDEhNfN0z60+slp
lfbXChTlXyQB7/p2vC3pkbEg1wl4W42IElUqzTKI+UOMtfHlo0chwvRish0hN1BK
nTaX09NlKupUAR57xXqlIufhzuoTA1qRW6HAOVM9EE2aem9ebJz+RE8qIau+xcjB
b9+HAOwovhrkC41dCRjQ9pZzseAXT6nAQoV++C+pt6n4tLqhQU0UoF5SM2Q+v5d5
7S6ap1hZ4chie3gX+DqMnNxyy6gQNTqXTOL2TYKLcvdZUrh0vJ/g19/ZDIX/wvKa
OpQf51Eu/MElVRrVF84ijEi79QCoLwqod1+vCJ5OaylWCjBL7SwsfGVL2hQVQ5SL
rlVvg+I1HIyBB2dSpFQwhy1iHNdv0kmcULCLWMkcDohpNPfXXs3uqFkTBoiZzFm4
8U3ko4HxW/PuNOf/+ZJXA2d9J0NvCehmMExUmFpVpTakF8b4Oy9BZH1reotee2kc
nBU7qlxAPef0qwKfNe6xcj7hfuwy5DP8P4GeKsM5NSkO9H4uJvCeA4TLPixpFbeS
boOHsB/WuCDY2vcreOpp2LP1TUXJbiLy+fb4ng0QlmEdkMihyxygMUUsnUnjHZou
kAViY0DuifRh0iQygTYs8bgWrfgseZiY2sX7TX1jPsnJmvOZA4+rSCVCjOxWX7Tp
hq+R0feXHcBxcwh3GFL1fPCB9+dzS2rIe0AV6EH5U4gRG9xgrPGVOAWEfvPrVsft
1OG+sVKu/NvtPPQgqqX5YBd0fmwXXvk/1dOwfAjBWaJGpbCuLEIv+WhQT+apACCi
aaxb3PV/58EKYMvVG370aQEQp9whP4/AAuF+QI2+wJWFqQWzQnlgv8a89SL2Of/M
ZsL9RaCOzFwWP46sj3ZrwWe0AefWEUmxRKHVZ0VaBpaohgEa8dDBRap4e58t+DW5
uk8AvxkZU+aFuFvZv+Trw40zNZ3dL4Wpnq4lFTS0EhKdJOWJ9P/qagZv9UzQuA/8
11zF+CSYTSqt7tRlrTPpd3+oZK510I/PIT6+0B8zrctawOIlFC1Lo9HFgh6Jsx2u
L9tUWcJOI9Oubc34dAzn4O7GxWhwKljZxGeBfaaTcItv3xcx4l4GxnEvIQXQXTcf
CwDnwKtHm9VfmqPwPaGtYihxoswUuDROUIxZhK6qyjDttVcY2U6EsbfDp+a/jFF7
sayy9cegDLeI/fa0hrODT7CWkZZOE9mBMhzGg3/W8PP0IdaiLUuTwVPCO9kcT1M/
uIMvdYEOrRVKIjQW2FbAwHiMYcSjaXpO8uZf+OPBRd6YjKFH/Y138ZZj9RiD6B4D
aIpz7KDZ97ZZZsQiHirLA7zEs5ehzXyhq3G9FGTIYAT9nsalbS2VWXHmlcEVdfpG
dGqTnQyK4X4g9SaxA4AAUQ0HzgqEEZ++i89+r9SHcwoNSLV5MnUNcxapmYdHr7Jq
WLzOhWDdyditKbe7eiRMtG7GhnV3xUZLkhjMFpcq44IJIxykr4EPOQ1yJ60vby/F
PEsQnRtMQ+nqsWa3dkm12NyxMwmNkW4oosel0WIQORpUnoE6etHySSm3UnQ1YdTs
sccr/lcuC0w2ZB3rv2qDrWM+ofhs5UrnaQwwDkauTh87b3OIg5Im4tPqTqUU8LvF
tow5VPC/SYtIGErePwzMcC2M6eQrfPKGPng2EUCyMzTdhUVEGUYiEIbpSWZo1k1y
LtGTKUICtUqyKTLUZDftWDNf7GzUuTPUhaBKrvaS7vW+EvtKtzXd4ExslWGjyLFG
6+Nb0giUXsKy+nQnkY5G9+TZO1HdPYCe034pxOB9Pq4b3x/FtPzTBKcQAQm24OyX
9lwc/lWax4Y44J+/Ko3NMsv9KxJtR1eIncZBDlQLYrzqeJ8GwJ0qkVVin4dj18KA
emy4tjLT2u5y39iNM1fT1gOOlCtAVTvOPbV3+l2XPcKiFKxhMNpMyEI5vCaxex0u
OCCH89yBwzUcWITpRaQuy5FJRW/1khrI+cL/XCVaWmkHNjn4UiysC/SGsCkzl7GP
dMo2qDK1NwTgvZx9tS1WCGmYbl6ppyx6qraBRcra5ISfXsw3lIIBYEEnDvlP/u4k
CkjgiNbL4Hj8FcVzoGxX5FLdO2H1oZ1kBidMyK39vHO36EFSxpTSH2G/WOnqZUvx
ryjcGCVZR5WbjY1qECiBQaMmVfT5Lc7onG8ZAjhyRR4xdsrZxsf7YkdJIO/ffSfL
OnAsIA3uflkqwBq02GPOpyFFcaggWR2VkgpkXqrsH6Sb7o23w14/549+dpO5oPz4
KgkZwUrOK8SUXjhhtb2rpwbahTL1YGNpg+CSi+mp1n1+NhR3nn67OW7Qcz+vxNcd
1nvjMpcw8CbkhNwM6nueL0S1w+2fQ1JbQ4jFgeS/+FA2FBKzAW768T5gyoEoQXtw
gbX3BtEI0hVmuDSKCIqMQNNqhcHki1f96vOW89ogvSgoO2LZ5Q4cPbj1SDOl2A6i
a7XiXkGC5CR9QUfcCnUsQVOcpyCiXnVEdR03qgL9fD/R4C1sM/9Bo3pE2oodi0o3
xFoc3bqsmCuyuM15HdwCBfqTFGHC2UiFER1w5H14m8fhpfLT0Mogc82B70eIOtiK
8nDYtbn1odWRgVLaohgbRKCdGva0QzKYa8sEAAtYFoDaB4uVUSyQcPgmSLbwN620
fQBC3W4s3Q581fROmVNysL9JGe9+P+I52IqJvwz8VkHDXUKFFdNwGf4gEK2ZcLZH
a1Y6D7KqXUHj0gVMQDjFtykVxgu8FcDi2ZRtSKYAdn4izZWfrmdQN3vidVlxTFmW
HO8CFbzZsi5d6Kj/aqbeVj4H6aSnT5BVaP2DJoQI6pCcvbSc2aKr6rG1583BXg6q
sg0/GWRwhkBTeK4VUYQmS6dRRC6URmo7xgTbM4+FGEOb2OSUfx3kC6Etx84B94CR
vvN4l8EvkMtvww6MFpVlVHoylAZ912ebmKvk4uh596rvrELa3tQKfrmdxC36AWil
3cqNjy9FJU1kkrVbQDleKF9n1abE5CbiQGNjZeG5iG7XUWAV3FLmYEicAUajq5YW
nsH+KSoUrs2NnxfK51pFfI20gbTsPiSe8mfspRPhQVRaoa9NEwlacPvpQ8Oc9rYA
Pt0U8lOHyIQMVcAltN0WPFEFB6/6ywZNsKLz8KE5RWCifkXins6qcK24kd/twjHD
8XKx1Y6sP4thw86NjXzF5N6AhQWsRlsmxTJW4UN93SyxuCuSDpwrZChrCX/hKvnC
Lpk7/9PZimqdyItHuCPsp6Mlb4fvGgF/FqLi+D4xprYkmeRbXbMEShig86+6I0z7
96F1SxTG/cdFPC4hq1dJ1Mfmd/CCQffPuoidFcpiufk+AU7xbcZwEDJPKS7uUVkw
6oSvLL2OR3Tx7QKwLL/DYWK6JyvXc8+cgQgyIWYc+HlyRE/38/uEiVVrJlrCezgA
Qb1ka0tkuZzxXR9KiMdqBxfRtixwHWuPT0p7q59hTJFsYhgLEewEdZshBsb4xbQa
3HBvllZjDe/NNQTfncfoMcrEjl3U1KcRRmRy1p38GSyCcRAzuDH9Q8N+gBfCY++k
MpIoMtwu9VDAduEFnWsQDd74jfT/oZOJER62v0HV7eLScKEnlA2vYvlaJY6Xizuw
OUIhyORX7/LehChgFb7hkBM/Yf6Ln2SPgMw0ebhvYESjo5m7tr65igEo0qvjXG9t
LiPVd8rIMPmoVjQLA9onhYzdsY0LFkz+sP6W3qFS1UmYOe5vskCp15nL/sVpYa7n
C9rysTk/x66I88RrJ02NVF6txj1O+aVMJIOmiStU3z78+ZKbTGYi7XmLM8VkbUBF
TfPfZWZXYw4W13KYav7SgU0AB8GaOSCSXN1LIX/SF8tcTe65lklhL9P8kYwvHC4V
jhnDApu8S6dU9crK4uQn7hm2QhPvzWVhsUW8iQMBoxuiBPlfoNpmcu9Gy6jfr5QA
miPSgPGE1Cd8jNjvBS8sqB63f9Ls/LCOQqK2cN9Wu1v82QY6TgIKOEi0wqbfh7Ci
+TJd6/KbvllsLjyeiR96PxusMdScB8ZenuYZsaQBFg37JmnCmzJth4eEXTnapH8W
/uxO90c4ZdGKFdtsmGGGOFqdCaf3DOZpV4EEuWDlLrRNIyv58ZgE3VZ+DGRbEHjd
YJ12LfojoqUWaLUsNGX91KYiI49nV4ubJjy1N5jDH3TwOURlHu/D1j4g8D9ii2fv
7gbZILg37B7HfDKRla8hE0TMaSWgrhBeM89fxc+e919iUFCS5ohD6fy83dmKynvU
58lkTBiOT8EzvquN3BdsdWuJlVo3TiA6u65DlTZroZyw2zI8c+1rTGFfE53Y4TZ5
NrxzsIo5HgljJGRvPw55RQdpfYSwvMro7kfrXF30nKRgpTiMMum8tcr4BUaJ5JLp
lf2nj8PwBnTS0hhlYDpFCXiYE8v8v2Ex+WcAD8ztRqlmBJv5kqTl1JHBjuspalog
sJsL1ioyoJv64lEXqkyhuwjqVaQViwcwSOjfwkBQdjaR1FRKOX4vHmnUYo+bBy6I
M+8qel6pLkEIyJ/Si5Hbj/Zv61pcRlO6/Gv/+/q+AfD1SFGn90878SzwJz0p56ZC
ncWvrDYPbm395N0r14vS9ksaWzOX8WitBhDHbOpF2KrPRIo1ewNVN78cq/ehDfE0
Wq06y7Ptgb3kARaKVYb72ozXEpDsuXF21OetbjhhdxUeWNTy/vhVGt8R8vUqgLHD
orW7EWrBEOA8UXP6uijse1QJk3/ngFqBgLO9VJoXxTzA+c+IYN12hrtGxHRSy+zj
SCY6hx/eKtGv8fjAGr7qZDKLhGlMgfEfdrjq1sIT4IZ/vLtCweXyvNWhlzh+Tk5M
eC47l/wfVYvMVSLygj1Tt1Zj0FwQNWls9qSR6js/DLO8cTTxDzoP8t9ySbsKfNSN
LRSUoH3ugVDguihJ261FSVTI/xHlvQFnhLf3I+fgEZZ3ImzfGL3Lw42kW2bSqlR9
3Og2fDk0YQX9WmiGOq/fSUf3+StB7pJhKpBXDh4JULZUb+ePFCsHkXAdLFNCO7HV
FndcPqLbF39bOgry40KI6d5Vel1E/hOthG8DY773wNDoQB5E5u5ktejHDpZG3S3h
VX7Rihc3zB1K9nW/62O+zFj3cvx6fzOBDegVkpcKXuGW8DzivR/1OmIvVP26aax3
X8C4GRRQX5xw4Fewu0cUqUr4GH10Lg2zXSfFodDieGuX6/iSgaU/63srozskZ8YK
CHnlM//I4lJVDTb4Fdmomp2Mk+gpnKeVll1/GfSY/m9jGuqffCidLScKyyJbfTr/
1fyz4604Oou+VoCyyJQVEWw6B7p9fCJCMDQiSaeAB7XdefhFXlDnPgpGxO2jdiUo
naTVEcbqHplMu1NoXcv0UKXC+B7wO3s90VtcBWxs/Yz7VdfOinPV6FSwwdukR5un
Umd38pp0LM+mIbK+ir1emOrLYRXxsMchW6YS/lFJOOZXgk6i0+e/kl8NMVj9Uir9
u8WgmtZsoEOJqYqZ7nPaQ/aeXmpF/ydjn0P1LwfnV291ynUN6P1Ort+pIqdGVbWB
HRZrec5dyYyj+0NLAKrIfgBWC9ZHsTwX3y711SIkwRDCXB0wCqycCx3lzccApbkN
hws5gmvOSa1bJqjOERhHUhf5oRoyGkGGjquFzHR8oRW/eegg1ojcNbJrdi3mzVNo
9/Uu56IaBmG1Grh/pGFqrz8FHhfTNyd8HY0oGpHj4gRpdiCrNh/qwTUU6/KbJm8w
ywIm6VBFv1uSq3SITA8VoaTlRlHrSnb8OyULdOQuqw4JiKQLMZAOXsa4OgmvWp68
qtFZaERijF/UGcpvmwrylQZxoEnctGJe1gC4Aqy2n4UVb+G3+kTlB/6Ot/c3R6Tp
5vU1HTx51sSr54XioOtk5cYHii/1RuM+KQlCAFs7vuRtDXS3ixfIS6C0he5f8n1Q
n01iNWjwu/Y0giurjKciEAhSxTIPSCpipuLqAyViJnWVo+SMPfreUasBrki22lDP
QxQ2G/eRRyq/rMHKQhKoGWKUiviwp56Sp0PWnkzU2zrUpUetqrO8aUZrHhHOdaLG
aAdEEMTAwBNG9eEDlm2dFMhcEC7uMNcWVCu2rhJurkQwCpfYLdKbSpRhCKtUuDGF
IgenEQ2Vcrs3u8wez9vv/nTtocvy6pKdy1inePERks4pmU019Ra2k/uOhTfw/LGZ
Wu446xFJToB9tlALCuvKjA+lxte9X09iqwDljCmtF/TOHZQeP+RxCVrPK31kG1C2
jVdoAmrOJw6JFH475UAnZ8ncC3w8AZi+SSwtgQTH9Bt25Qpky5y8KsMJZF7x2aNv
ETnqD1gVUHg6ZwRHJlaPuq9xh0Srim0x459YMho/FoEuepdtXBf+WUB5Ff/VnXjb
spNXSFpnXefQ9D85TBmGYVogd3qXZFxxU8zg8G3JPZ5HeFqCgBFk8ip3a+fII1lb
LjB1p8OMOsUaRBUFVxWGWVdfmNi6SxppeL9RTMEF6w7ENMAealcUureIRGoLQC7l
djL0zb+uYCJ3/G62LFkkTP/viN+fNjgEmC/5xr8H5Dc3broviFsUCgW3yjjZ+J48
+lrRJ8uA6RfG170vCVxgbIG210qSAlcGoLdee79S8xAyKYRaSRz3aj3iqvYT3NxZ
xaIi9L6TdkJdwNPYvUYhNLV2OlOpEfCIGVmKvA/QteECH+n09N+AA7JA6POcoSKm
JjXoYLkwUwRLx39WtG3/5UaSL4LlsT+Je3VkeRyFz9we1KyHCAxibJexLH2FUGWP
t8to8WoX4q6pw/jFhpLx7IsQT0qIvt6mx+4OT/QXOiP1wQqimjPRQ1QQTHVoxET5
QzxkGoZ4TG8uMNBqdO93ERIuZaeUu48vwo92kPuF5sg8VYW0qgIsNZ6FnRPeNLrF
P8wHEZWRGd0ObfVGXvsah+xvUy4p+f+F5kWOvNq5mYjVhF54eur0ZRPxX+nBHoJU
7dLS7+5fw7nowhC5DrNpg1qSlLmhynIkc1rdr4ucQmQ7cf5JJ0QLUwEmUI7BACAr
xFcKHrwQf7Ftjg8y8DMbRcwheBKkFxKN1WsnL3hbsMLQ+ePtJ9mPJZr9b71S2Pto
Hazcr+nms8STQ8Y1SKGoNCH/seAf2hO53zxa1AaFJ4YP0HIBRa9Y0AX4j3hOmn/d
RnMkzPWS/2//XBM05OB/XHAuZcnHaXw8bSXn4hImjmWLuVz6TMcnR1jbiamZmrw9
WJO5dK5PzwhXruw0PnfUiIzynltZUYmOOrkrXPCOYDoC7bUCfuGyIRhZSVguJMn0
QETElxjEuFTLTOM9k9v18EEMUXlfoDTl/2qCAvg8k0WpVP40ya+8yuq2rzpTelD0
/ukVx4SWaYHlqITHC6AAAB5K0GULhMweAVzynfmbNqGz2V/EHRymphlNlrfgHNBx
My77mi2JfvAsfRYYumS1CevEjUj1kPqIWt2OuXzp0gRLkNGhnO05IlyeBMA8SS4O
Zybln4ceQH09/KkeUtaBA79OdNTDnrt3nEQ1rdRZ1t1Ou6GuRqjJQDyjbYu9SnQ9
duDQQQ4cCmM6mDWEa+gu2wxI9iyZl416LW8fi4dVRwOp4yZ/aOMVjAMXIsti04w9
SmrC/PfhvmMBqsa5LtdJvUVljp7BUGOapkvhukWNaeF19XB2dpX18c5infM1I4Mp
AtmFCmed9r33ZZ/EH6sEbMbumw43Pom7mLXHJ8ptLRo/5m5HL7Mjea++5mgRA2Ut
zjSqFe/+lxFceahfaEqfVw7OtUOhL/On1zZ2wLR3l24GDafk49FSr6XcVOci0eVk
LFcBfdV3FiLLdy5SbbVJeUvvXa2haQuXnqWg0WDv8hq2yrZJmK2Py/5abe4s4GCn
chmogPy5Vu/M1+39x3TBFYXClVhmbSWw5fs0G9H4W2YTXdjlNOmaNVlss4OfZwnZ
sv/wXSBiDZqvRG6YxMCJNu0BCnfy7vqugf0M5oYJXAt2LwT4OQnsoXHdxCzPi2/a
p/YOK4yFpxbjHhFESvR8OCFR6j2EK0lHiy0/SP96k54+1RvelTtCpfvU4IGN0ZO8
9iBaM5ZrvP1D3kTwuarCJ0xCXdvMpNkq0+8U1S4pAdVnsF9DUK8TfDFaOL2F7iZx
jYx97SDlgdqaMK8e21MVXoo1Hd+Mi6GO+qJgvrXSQvzRxI8+Po0QuvRq2+wIwweq
txQ7CLdQBzLsogiTfE43VQcvphlbWRYCbcor/rv34JRfp9HIqypsYmtwSTgGZKKI
IkEiDhvshvHS5T7SMCgKfu94wT1lOoUm/qkfLyjLub4c8QuRsnXe345CM7BNjm6V
4mEJ4Z0+XJ/YJ2XMOA/7ihGOiChBu7gmKbJlHW1vEGI3YBPSSOyadxKAjPaPIoKr
Qv94XdgDYfKlbJIQWWHKoGynk5xec4v49GceX6WRj4bAFyiw/l0i0YcbFC2FQFU7
BDhm/VXYFsvAId7oAg5fTrLJisnbZRSfKkkfp/H9elzptixOGIEp/SPnDYhE5Ono
bPUmOxIwxqYivqY41HE7bSMWde89eWUzqZ5ZKdAGppsoEodMPsjFEyPK1R0bPR4f
ArN61ZLOqRyEw9tDXeu5Sxf8ymurykBelGZA0qeRPAS9gN6D6xGSp6oArFvIKBWI
1esIwDUK63JBfV/Guy2CDxr979W5kEVChoSsgMPB7VgrP+8+61E478DKGfwugRs+
F909517SPff0yX4uLct2/kCupTkj+wawr7Er0kim/v+63oFyF9lB948uE8j9cc6O
PjE1dAm71FM2/MGXifQsAe/Gl4Poy+HL+xoZpfxSTuwA83HxH4WVbLgcKQMDGzfq
tYpSiMfbthAJUhGVRJ1mnzo/73kkVP02xwIgM+Z/QPPY39iijbqDvo5s6jg2EMcI
2Wxlwr9izAND0Nkm8ZD1ywcGtz/1b3nPpr9RpIZ2wezfHy4Jlc8EfcZHNgPWTZXI
ml7NPXj9CP2yUji4/r5VHJnMMWjdQTZ9CW5jpkzDQcH10wxymn6l1AMofKPrpgzR
fju3DieeuoH2MtAbpxrS8XAKBNe2p6u56zqLtmztiHW7CCdrkSv9Wf5M6JBZRRUy
tkN1fcnyvr/9RL8iJZKvRGTBkOHWI1tf7ff9IrY7ICnK7tnVFh6CmdmTnQreNbwD
u8MhFQpd9aoTxgnH6z1tXXg6oXFVCj51oYVGmPEq3aEEZI0yMWVpBim3YaHaRIHM
Kv+zdNodpHyoZ4MQOJboe+hYj4GhlC3Pgz7e79H7ygkbze2qTYlUge3ddKxzf7AL
/jabRl3dYWZNCQpAnBa2sEuqMCV0xStANsodH2j/e0Fzvzm/7WhhEYiOGIMDUwkQ
IKHO/ECOm4K1iE2F0aRWokZJLgIJD5kAsWeDbQsRk5fHxXxw1bPb8UgGA+uXqEIP
CBeyLqRdKCKOWUwIdRRNEmmQT3IGgUpKWqqpquTOKWl7Fm2AGFSTrG6Xq+BVOQLP
d231H0uxMAYesOQ+iyUuPVGYsknewnu86MFMKUUO4GgeTA9PpwSOmcfLn6cJW+7b
c7aQslFRtK5LOoiFfMrKbfoDxq4cTyyERJiqvvk8R2QmMbP6Y3uXjhACAb5AvWix
LYC9jNiu+SbR8BFbD0xCg5Pe96fVngKDC5Q9TrUb4V28q/qCS8moyRlWvbKfXP/A
+97aOvICbsWl02ufAnshsKdOiuP7ZeRsrxudiczFSzjyqkBnmYG+ZjJ6L+ScIS/L
nRh7bq8ba/yAcNHDe1jdmsWtaCpRHT0/Yr6t6cF2abgUTvUz6pdJdhvT9gsXiKCK
y5152NKIBs8XwsURn9sBXddb16BKMzLTJTnjGQKy9pxnGM1u6fDh5+cqRRhnydq/
tJne+Ala/PXp7vf+dzOKqaMcZSCe1bAvsR7o7dgjrEQJWmkJcYTVgAfYeOQYNAzD
t2kANiSY03TVSRXI9GnxNfyVKPG5nAzz3uOYStS7YoY8hUDCt8LhXUcJS95tDY1P
NLN0pFV9e33do8O1Rmh9DjYcin9UujyMTv8yis8n0Ha8kWIyjAg0elJjIl7XMzvQ
xq5M3rxwbYD6avStBScpqKHmEAkwRAZUTCW17cU6Iupw2nvhSjTlgZQy8Z1LkdkO
F5PrKit1dt+ozM2C1FanHb2qwV4/tjZ+DngXFUeKElrswd2hKlZUTbaqBTP98J7M
1qeAYPU4YMIsr62k4r64rt7TcuB1sPvBddRz7By2/Nqc69cbOM2ubwhmJ1Msu0iS
nMRJO6nWUC5xeWOGteW89Exs3IckXCb4Cqhsn0/JKJmAiIKWaDUpdPLrQn0/PgqD
l1Xa2Tjsry4ZDomfsC6STz60PeQ9f3btW6WhzBo/ZxSOOgUKZFrAEPkgGUY+w7Jn
8vE6bu1LB4gotwSTazb9OfFPuCd/juCOZLiBBSoTsi2PI8MzxLdopjW06qlgWjV3
BJXJWs0BAX7DtnWRLQeipDtICKpMxNfBUZhdHPrZldthtHihJIrNiYP1+wedaudS
5JNWVb73OjVhLH2IAwSREyYUlerJXExCMI4FRDHo2CzaP7bes/JMvaa7tz5FSlwc
FWCsZwqIiFsPco3MTjTYWVwQegOSwWU2BY+9RyyHhjSS0b89aGOKh4pydPymoSII
PvIJL6AAcYFxc247arSiVR8UsT5NMNtc7SikDMP89Hq51KOvbNiBHC/nw2AUjzEs
CpacKFTokMOi7dlt+Bng227KP3zDK5JHtP6Zf/0pqj89baMW3ysJ9nhXbGxd1GOA
SIkOCJoEsG+YPOqdDtIrtCSjqKAws+iGQ/qrZWsBJJw2syU/O+nTIa/mnlzboU6g
zV55p4mAKaIwxub1R/3ndz8JZ1xxkK8Bx7+eFJEzKwnz1ZkU9CmdzT9MU6YpZVJk
nlcI4WIHlS+fw4QhpxAgisdUvoMwp79itw5B0I+JdgCxjf1MucoV1QdAcnEt5hRE
1liRE/q1SBSDYWGq9l2/gIVqyeTRCTvhI6D24QmE7ySU+I8HWjT0DmvPieL6j8aR
yXjKqVcYACbZfC9ZIrIiHVrvZXAMTuQgJynuAinHG6iqnO8z4xXqI4BirzxbAVZq
jgb23nzlhN9sbqntIOJ0Xly5ZaXt0WfSY8kntKTNMxQ/vs+U5bIZGilIgjdHFL5+
E5tXwlfbKeQ6L32lxsCW0VnunShD/TpTaeiHB4aKErVUSTrZGXqQf5WMV6X6Nar2
0KOJ5IKR7wHNljoBguVkczjSI26bHRpkm4n9kDE4lbkuFf315v43SxcYq+ZsJ/es
nvmj+hXk7bQj0Hi1VWcF7o6Rd8Vg6gWz3V5kPsPGo7/rimcOKjs/pE9GuU6JjY7V
wTQUKHExQxzvxqieWR0M7t1+J9spIdQWPe07zulUMm4r//DBhcrfAo+YEK18xU9b
LYWS671ZPzezq/fUIsfcvatDbIfEuI97kdeklwo2JacVXD4YOckMwDz8XJV6oFeR
G1QO7b3MBnW7dn1zrZe06Z3HZrqPWinECy2fQAcZYtrDAIl0pGHxNSzRQd+KDiZY
9ymWHEy+c59oD/vt+0sIvb4yz7qf/ChHuLvyYf4RwuG9NDjluxRw1GA+KpBKwrWg
uizRkqw+N6D/tIQUn8W17vsctb8qyvJni2zZIMnA9eZKdM9suHeZAIoU7Y6DGCuV
7QnPdfLTlI1XxsVGdUinq2xKM2r92HQbsGgXsBO+jsYYiIfP5R5ICS96vO2eX1qO
UhwwEjzGlM57pzMI6Dk8L6VFL96MiRLXK06FOvkhzFaxdwFy+J7RKOFc9m7KmUTT
irlXNtDRc4E6YYTTyi83x5TKK6kgSmgLJXT2cTdyldyJ14vHWZljiPpTT1ieiRCs
lVuDhHLjJvrD/wLWYhcJNeBZvIdzF8sgH6k3QqYCObIxZWfqz8fPjEdkb4abt7qs
d+KvzQDLX9uIU555bZ5z/wUp+flwDeP8YeNYqqI8GK/tM2PMcraIiDCHBVEbfW1r
joaw3Sq06glKB1838+8SMxpxjLlb7cYxYD+6+eOSTzqn3myQY2W6UgR4Fx7woAWP
Nba1mAIIxSZ0NQKc5AAku6RjAs7E4RWa7fCDg2xcBwKAdOqB97safv6cZxL7ax87
FnAMUHTH/zmjpfSNp3Jkfidz8FoblQnFBNcYDGpReQcJyHQY0A/FLBfGAnKZFFXd
GDBx1XSakO0T2c5q90VKJq5iH/vai46FxepK71PYujYHjyqMy2e8mbn3SyM5THUE
CN6Nf+U0UhcGc58uQt7ONzu81ygPvdiaZY4Nv0jP8hC9YuydWi4S+GwBSIlQHXDC
8AtG4ccYmNfME6vrKGnsbjHcP+zumSYlONQP679njS/4+HiDW+KlBED3HzeBfsQB
qQM/CLKL7hd5vOx/U5hstcAjRJahJ5HkyG2zbMCaNagTanUhVD5Oy8NJ29YUOSlh
UDm+1NR6V+PkH2Ow+0YuBWHfxskTkUz4naaiPEWjH94EK1bcZIE2wiAA2zTJqmO/
zSGKdUp6P7tSIHMOuRGbyj70wJosBshM7BGJpPbwOUdMQvKJJOTAp/TING8pmkf+
Y8MVxA9KH1xmyfj34SRb0ZjBit0gwhNB1BEsN2RZLgtSZQDrZcXzpcEX2TzETyPm
h1Wz8M3kqAQqoPs37Qb1rI4Zs1jEkiNdbwoyJOwPAn31Y6jy8laws9LuOpU9R6wO
fzQhlehyfqJijfgHk9aGIc8A6H8rIZiZ80/5XvLGR1koKwXeWjwS71wAQzvL7OE/
RGSaA/KvmG9lqpuIUuHq5Bbu5dFepeYRIneUzsCUuBgtTsCSMbd5CF7Rwc9s+JDc
k1N/lVEatFtNnkenk8tUwBDVAySg/0fN58qT3CXeMCCMPrnWND5mKpdgobdM66b4
p1IN6RPLQPjikU45Ek6LZZY4YIxxWEeITM6iZI9EvlmKJdyp0/hmc5ptXzlH24b7
gyVBBVqD9KI7XVlqkpt6dvo1NVkfVk2C3RgD4mvks4mlunVBC6m2eq5fC+y79wAT
VdEzgPacxRzuQRU0xXqLZ9ORROMnt08bM/ybTLJkLkEo3X0fqFBnH5dixBEloce/
chHE4o+hshUGNUiJghB85cgid4/9nuHrMDTRRtud9mhue/fztK91E1tOhrlXVZFe
VpCRB966YdVAJi/y/ki0uLTHpzbB7aRC7IfBpjQ9ZgPkCFDs6HD3Dd43WNxAkF/7
/9gNgZ7c2n7Ip7871fw0Qdj7ki2nvOmWx+/4E1QzBSMx3vmPg+qOduWEYapJeUcd
r1cDUbOTepkJFz1c0gwib8ykqIaGpckZFzjPnD/wZdEeatHJFX6p5CNNOhWmGsn6
QnZlffBo/idyyfGwDbjEf1a8LgNat3e1IKwZH6sy9eS1xeRLwi27n7zY5huVzrjd
tL0ZIIPuJQFEU8erAnjoMPX7NTOehzklIxGDWopoEZOsEJBN8TcsrJYV/sXZAXD1
2wOrGJ6Tvf4whMfvsbK6U4cODLeYA2wmokQW9pLMFbiYGW6qjrw4IrWFsyn8b2wd
lMm0oXg8gOpJvUif5lThTMGpgnh5lVs70kc3sl6KtEqDKxNgD6yYh9sn7ECqIx9i
uB0kSQllUtMAterM3beAK5n7iJcLNAPG/+2QNGtPVqYgREBFE23pQ5v+a6tydxDK
IDkQmSKNrul5/yclerQbTVEpcnXGpLaDmHrnNEAWf8WjVdIW2Dv+OgAoGThrKcYB
GmrCW7yo/1XoRhYhnfz6Vok6OKcVLCdU+nZ5hTwaWkP2y5xLdBAtBu6V2nsX+4yQ
WxA6DQ2EegbAdf/vAs75p5yAxXOKGLlKM2XM9EpX5tjvAjBkP1ptiZ7cxnrNAAiu
es+qzMiq1/Fyz4vf9hJc6RHvg45Bf12n6Tl4dKu8IRI2XvtMRnZwC7q1+RNoC0hR
4jO1bkTBEaIBYEm9K7RbHypVe0tpoz20BkYL6b2lAOqK2GWQhGWcZNl5fV/WuIk1
Kj0cMi9bJ8fY9OlSGmGV+bYGpJA8mmTaJUbu5V5VOzD2KVnvafdJjazi9iceJWzc
KOt8QPfH702Vgt37dj8EwgG33/7XpfZv+WzX9pMxRh6dQKrC33ve70VB23+C7yzQ
8hZzKwpEmmU9VFuwfnn/byvC7RSOkPyUZWuUQka0J8CId7ZvutUNvwuYW/qy3Kxc
/KheJM+Bt8CYLK3fqy8eazpcY0ZlEn+/U4SuqbhKkeJgs5NoADxCw6tQtV2esAd7
uHxYrNb/mpdc+xiQjfxg4uTkPo8fJ2gl3EJJLHdipNUrlDU8FZVePFWhTWVpDGjA
M1/I1+77yvnqrpUvg3hnTFx90jO9WglK8KulSARa2/D0kqbyDrWbNFAhi/0tJXKZ
2QrkV/SBEwdH6sxFowJpMfJDB98GaiyQqA0sQ6+gJNnSl81IWgq3SrgWPAE/Ffk6
+QL8mLJfkcfGGuQug1KLBmUIe4Jdzxoz+8UlE+EWuPg/7/okrEXl3U7TNhEqPWVY
ijNHpV1Izc1RaliN7jrwIuPmKqnK0MSdXTD/mI3JFtqqvW+PmmIApxy4csmBdjR4
ZakMrvsIDc1AYl9HpxNyRDyS8nBqwIlB62a5k0YtgeA13/CqcuaxAWdfuWjNKHH1
V62a02Kim2/2M/halkYYEOdENBRAJDXN/ux730BEzAPWOnn3qeWXxHyh6IGuAWnZ
1oD7ia/LlEhdxxYz58KhS1s8Dq6bblHpLY36j+ZESGWgj3sOpBczud4xmA9A3h4m
DYWmWKUChHHfIZM59nM8Pryx994ClA8/LHfUhGcWB9vrZK/U5ExsPRxbBRPxeJyI
dJXTcE0AnIqgMJ573uRAUUCnLbkF2tSEO/Wj2FXxlWa3RhC0PGffowvDAuBOJI5m
1ZaFyW4AfnVnd3sTNNZfgM+D+y6CoWx4+LcV6+YuOq0PCv5dKqL2dIbPRdUv/wSE
yQ5H+uq3Xc5I1s8ZUpcUi6gfiVElTAfQN/Xmsv5i6Ypw+S7aK2edITVcNYx+h+lE
mfwlXr4eQ6SzS08EbtLYYUMhUCnliOnXj9dgJsSw/OtBglqFVxFcD5nnGFriEEyu
0tUBkDnl+npQbxDLLgyFydXZwhflCFxI7LlPExlPH7FlvumRA+RDkM8PnkA2OkKl
gyLiogwiBKe8oA3AnF6to/d6YFW6R1xmeRveL4FGUKIMuRCtXh/ZmNdFPqMdy1Mj
BV0J0Nk+yupoIznLKMbyE76gLwVMl0Rqjg13uPW3FzR5CgHvXCOFGwmyoj+z0skR
c82uDBQnh5t14Ro0Q+vICorSh0I0s62SbethcAIm4+1skHzM0TBAxf36Xyd5B/wa
/FUqT8vGruNdhSoWdUvfjBS62pgVltoItgo8ySZEfv7Ru+Kzlfln5lvGvDhB60Cu
turYrx+lauclbGbiIT3TrSZKxMgVEYxq0hTMd74wyn6yUrVomcMdUSkImnrfNhCN
Zv3e7nk+DVVSeb718JsZt+jFoQeZvzAwY2ynUzt/wVdFHuEK8KWNJUGDmq6Wo4ZR
YT7ieX5gA+MmgOfZSjj8Y9icKIECZWSCEPgOdRlKPGN4O4ufKjIPFs7zoqmxSxB3
ASsg6jM2mrdC7LuPwxXTqONmiADKSsEz6HFLMINNsSujfUFnQoR/q8JGbfvbblMk
AEECxIq5YTBP63nJmbY1U+/vALkineYehBC1yijFYcNuYM0+tCxbP2006y1t0iLr
iKQjbdxvRMNdFidCZ6AgX3Xtd3xYZXZ7zeU33HHrf0iA5p1+lspkkvkUI+hgb4yo
sDiLLtnRfkrBAQa07HDxJ9AiRorZaY7uFSjxFbbPrh+RUDEIWaXr3xxI8wScunEP
kNZRuQ2gRLlmdEB5lT4YLPCb9vHvGn50/e4JfHOFfF3vlqViQ6Bb9qmcCwJg0w4E
g4zCIEmD4lwDM6yN38dRybzMIwPWBZaNMi7Qlk/Tuecdx3hVx8OWZQ6/bzq7G4Pg
gD6gjuUHmXRo9BIIVCFByBFjBPi6bv0uR3dXopBy8v1XafjW5ILerWM2JBWwX3lD
BZFswXrOBTaKBZlOZT+klBreqYKpz0AfhRlYJrs6g40dfM+7d82XWKjxReIfOOJh
pIIbRmezozB+tYLOtQxAkqpR2TLa+8WlYZho3ANbONKrIhZDy9sOnjErLJpZkEwn
fdBPaGJAJjDEz4Fme7p8ekZZRSnaBKt/NHtwGPBcdLFVr+I/u5WFiJc05OfVtHKF
orrQ+4fZ3osmJjGreC8FvIG+j8H3gE+5EoRzvyXkPIUbKxY8LC0/1BhNf9C7rb2C
9bW/380j170YaMETbam6jkMDcgjhw3QKJOAEW43Zt8q2HZreww0LQp30PaIJBId6
et6h7YS/5dP89fVufFxU9rQ/h2SFV8UscbG/q7c6TVrtaHyTtu/Icnyoe1Emom27
4pCBAmdaxOEMabOgyVfsvH9xTnb74w8Nx8JbXRDAaDtohGiCwXjkJOjAa4DBJzYt
rgILrsEvFfRG+Bi8HxNOuA05zR6mVKFaHht7HR2ZgUJX+OPOsAuZXHGTKt/Veyp8
slIQHH7hRmxMxwKKcV3ImB6daWKjYlWgt0mxvYLUaLLy2EUAsSSKj1whoRa7yG7v
Tx+shdQPg1n/Kp4ZIcG/WIQa4MGicWjqhSkJ8bNt6dFKwoNkzXFAW+97yCx6yU4x
IOvocaw0v1dRjjsaDDWEfLLoR3INANaeAwopEvgdVMUDM7RSSRatP99E9zFhOVcy
Zl9SPfq2QTXiuOcFUthX7PsT3RqYrH0nLNV3o0f8UB+Kk8iXwg1dLJM0y+rsTBd3
Lpt2QvVGAMt1ziT76aolXJWUSnUTIP3FAPWaDNsr6EqmsUz9l5fSp7h9tNEpXC21
fmylVolScffjG3zVxj16UMnnPVbkuD9IYfERTKwQUGs/96Cdl4ivG2w7coUcw0G9
tcWVtUdVvR7Fq6NHAXccVuA8oQcEu8yRPnaE9/AJF0dWqMPSuOoh2AUzhCbLQrOI
ST/yqNoyKrhBbdV8oXm+wKcObOdHtYUzljaeCRTXvCBcgQrlYcnGw0w4eBRiPd6Y
51fD5KU9SfcE2JQM+4kXZJg1DfWM0chCloFA7ZGq5d8Op+0KEs5POKNeIghtXeBE
HNBQL9HK+3grdyBiBEfhM1MjlrzXqETCbetp0H61hoa4+KWER5ynFYxEqOkciekC
9E6SG65MG7OYeReBQiWussw8JmgpTLGiv1PfmPLqEQAyiAvt4irboWsIYwNRhZq+
3BVKAHneOgiv0fnHhqecuBz8HU350sngztBz+d79xMgjCUKJ1rNPQoEtqiIuftVE
8SnNxNAvbp6oQs40o+HrJUCT2K+I6Cju6bSGqIATaNPyVyEOTRfYf7pRYZx5ZjPv
NxvfwTDTfcHx20V9SarEeoSFE7CQEPbN/JgCLHzArVgH2jYZiOr3iMOsma0HcQh2
edI7qj2ha+J0RqJP9+8J4dOaI5+YvHOT8MlA4m7COXebHldU7ChZ2dnVxlZaR+yd
LQJDApdMqEIET+7bFRT3pxdJII7dFL/7D1IpNM0vDa6pi0dlNtxMovRuJvb5vJnl
zOfowwMbyvo8E2+T4EGqYQ==
`pragma protect end_protected
