// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:46 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
V59alWLrYU6RfSTvQPRTFCfdZmaanFrGj6GQp7xpp4j5yFY1W8iMbeiX0IvqmyzU
W1ZwSTYMb/Xo20PpQca8HT9x1S1UEh9XnQYDWe2uAAb+x5Rf047KXxtp2Aa5uRfL
gsGG/0mLWMADjLLhfxx6/K5TLA6N3/EpJ523MbtACUo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 42896)
+//Zh4/XMr6/nSjddjiQWuaL+LUn1GDdQrTmfKfiICFlcz21i9MBrHogQVJ1gN6N
+TDuvau7wJ2a0fmomxTlwwvDTgMbdeqTTEmi7lF56QW6xbZCTNW8dpEYZMlY06KU
iFJyCzr3nhuVKtUJnRmhG4Mg83dp4FTWLuowSI1J2TGXmNRwRGrpS+VDjb3IhWTR
VB9jRaG/IqoFzA/2vcdUTbXTeZ0c1Bl/Qg0KeEWI5oCUDAZuYlZzcKpnwh/zTd9t
YPbjRQN5/p6XVv518/XYnSySfyFxa48NG7I0Sa7HOPtPuUktRHnu6Z6vSrYff4G9
BR2/o1wDoemb6kGkhtpgrFhXVW35d+VwRxGbXejyY10QmB+i6FsDvSEILLkSH6Jm
ZcWbVDYDica7hoJ8lY+eciYOkNOsqx0kugpEIZ0pof6hUPHZv6g0McdAHtYXln6c
EE1xC9hhz4B0qtoDE/wTtC5fdnQXJAJuDAToct7SkU7iSBvpH6Ap8jBhHZkK44q2
JPgqvRoE4lTfNJpB4iJ7aXkTyEFA67d1qFghaXX7UdEey5vBa1xNh/scFoNQpjpN
6xR4EyMnpOpqnRJzLYVGkgvoWjoBkHguWwxO/lj382GNq9JDuXd16BcT6U6iaTRW
VIiwTMLEEKtTvNRbAXKoSioSrwKbMJRJYCAyrQP8sOvlCnroWIV/jsh9lq9wcHZg
UBtAdp0Lbb9vjU0NagEEfIk2AFpd2Z5ZYENRNAbxeQdZLwdoXWeM9h1uhDpVWsJ3
Yitq9mKGbX/Bjd7lYRoSDkD/qpc1P0+4osgfQyY70r+SXAHXMCB/vcoDxW8WrCgZ
Jf0euDRpSptO8Q9xmcnZwCWEo1gsMsY3ls+1pIMCj8A5iNqOlq20wb78ehNSz/mH
lu6emOpHJBUb4Wn8j1KrOHODKID960dX++d+L/ki/9vrSS6KjXFlqKFJ/5y8XbcD
kxPrq9uE4CVecPaPrwcswZb3MYOt1UsCWUEvB2a131hWIW5UAorNTOeCt6ik6acB
wQmdn9PxFRKya798GoB6PQqkBCtXWtv+RsnoN+MPVWO+twUjiG98gty3pmg4E2TR
FvGwEHBGLAP/DetNfY+Bi+Uh21V0Og4kIk7MoKWWo0xvuA13451LNBq4PPXDIJ1N
IxvNTSKXnjqno4OOhy++lgFcaHiR1VWWvB4r/inoFNU37TGfy0lB2UhJ4aNWPABC
PEb4Exdo5Iz16/YuBMooUAYM1g4ssTyhoa1Dzax4kRNPWpov+CdkekePvX3ICaP6
EDqxbihQw4N3LkPLMHquDUqImcCCGdU3K5xhbxbuc+ygAeEUH01YnRCsw7XtVgf+
rcqWAfbH2OQcCxirGVKOH8j3MlekY1yzR+BFxAy2jYPGNGPeAVv5CJ946LMmSlqr
XzoODKH4xBVVC9QAg2ZzG45FmqCQQZDqrOvheqLw4mikyI2qk7w8KXIIQwJ5OxZi
L1O2509WjcY8lJpPgxjh3XNQ/AzkwlDVG0GNIl2dKRKYClPax7cn2bzL8xFW3iEg
prBpFqsj/ugdPPR5sDRnQe+cGbbpWU4It6vrnBktOsqZeuOCNRdpYFImRUfy6wfs
FzzPRtSDwCpqQux0bOsBQrVfd3r6KxSgkSlp4L0rNR6Dq0xX1bj1WHq+3URZ3yWc
tGlt6tww7VCHGcq80iiBNV97VqOQhEhlgUlpbyUKF2qbRHpqR8U1477zZTenOSru
MizIp9Babx63kcTPzir1Fy5MrJL4ps2ETkV4uySZZwBATLkhJBiE0YAYS42U5IQ0
D5eOCZDMCavZ5b5/qLY4B1gTiuai0lyVuiULz6jXxFxHZlD+kcrxu/u2sMA1cQ53
qsrPLCjcX6gLwCumcpSjlh4C51E3I3hWO2GwIb86h71kmDBPHmvAeitllG3DCVTF
ENOUhTh55wQp5HNiDZH/a2SCDQEgZf9WXRLV00gbv01rrEQaYEy77pvG15D4leyZ
Wj2xe6jBvvmWxhz8XJ4tT1dJ+qz0KslrSNoHy3wQOSwX5nUj1DeWYKPBRvMYLaw3
OGuP6B60sohclbNWBBOzV0XZNCdw5Iyj3fwfh9bKWReped2ILtIjzz4qu3apIS42
q3rh7bEFp2y1kH9OkXG/VQuBdU4OdPUYf+HnAOfFe9CzIq3kRcPjqbFcUFd5GFWU
dT5f7oCDUbXmoml/dzaEzcHEMmNYmDK6YytFoEyXNwtQ0oDXS8f/e3uR+5U2vLha
RSljHB/7DQrShUm6bHIiiHyEkz64IGpAmfODqXD15+h6VZJeQSMNAqOFaJcLMOkm
xxJf+YnQfOWVBwFdd9qUuGs5uFMfMqh90XWJqnsSd1bPWCNgcJXVLDeMb+QebQWQ
/vViWb51tjMWzb5d5gE0oR7ggPwNOk1+srfC83HsyVEZl2FVltg0DJmCIGu4tMVW
x7G/j9Cbpm1DnUdMD2/dai2xacZUp8atKyZHEHsT5ciIvNVLoDxOuW2b4PHo+USL
d1g0ce0b1klsHmNvR+SU4AHr3p6P+5hwFRGQ8gYUdyh6qfbxcvBvNJXe3ugusgyN
ZGFAaRjxfBg18grWG1qPqalG1w7LsSAjgbL3TAOIbhjlEL2DiJS58Bj5n3/nqVg8
SxA62TgQhKoaQBvCTUAol8P1daXko9fEwb0EgCh5PuwiWqiHZLqKdkIYzgaNY232
6tfXBgKJNIEFcRVpkGMAdZz6COCMulvaRZtoEUqifxI+Qrglhc/elb7jPZ4t4FZo
7KqoaC2LcdFVRj5skf9lYwu9kTSGjhDPDtsdlfqu3aZ72fUctZm40cQxp01UlWiF
h+KDAmYNJqh912X+PZjrANuS84ZROEvzxmdUmcchGz+fOZrseUdGua3tAcDSbqgL
+GwFyM9bZqkocDuhSusPbt4AEwGdi8crLkjYGlVNRhV15PqYT/a4VhMZaT2gpjDB
ylBpxhzghU09Vv5yjHMzzh98ZWDdHxsyNfjuBTP0KHDSmbYoY10yWcEuoo3oN8uu
xBbFb+YQtDVMLa8xTF14UPbXhkeJWZqpyLImoZbjqCEFUadj7zyakmf+rKEStKbL
PP5stj8RDQ7s+YDC1OSYygIhfvOiKC2Vt1y91gXK/9eWBy8UTD38cC/qWX0sqMgE
inFxhVCyes9T8REXISFT5RN2Q1LO6h4ZUthFcqVsXQpmgQJds0LN5Pog129blUOI
qp2J77XaFO+V/oTKrEY5/8RQDw260RN+Tgb85MHBYKSYL0F2fQNTSRIFHBc8ntxZ
Xaz4q/01cJJYDL1kOEW50HWhwWYDN/lQEBD+tWLDjlGWnSwq18kGGF0VzHm7daaL
1ViBi9Dqw4/VEb73RyGLlUWswH58Cy2z1Cvg2PCYMBc32wZQePfYnX/H/kugmTIn
A6MIyWyp96K7K8RW9C5dYkplt4+RCbwinlPRiggeFytCTXsJ7q5ugyP8W7wn6HdE
7mAmJCTLRrVpuytGh8A7lIN2/xklIe4D9zzjTAI3ECXrgRv3VCWwBe52IXoyuOUO
uxWXRtaFVyJryhyih6Av6LcQazOUYXPHDzgaNvhuskHbaIlhoLLEBab3Krj45eys
oSzdvP5VkitIYSchLiVPC2Tk6wy8bPXmMmuz4dKMcUJnbKeBUV2UyUkaBD+fACvC
LpJNACZ6CqVd7gOjt+rYa/Jl1i+9MfsR2b7t1TT4K0vQJE9G2p9MQPbp2hNDtF3q
Shvqpgv8C60AjXg+85JBAYARz1nAsQGGb35mXmuOtQhyZZDtlLUWgMCm4+gAsBxt
2RNdkR2bw68HpfM4Yq51QQaLjLN5tmh+FXaJ1+REbZ6+E/BZNV1RFrrxDnGb9lbY
PE5IM1OlNM8d1rINIHoa0bYj0Jl1UNzI7mh6lCIJWPOStwyVmDCphsdGV47707fC
tJo154zJ7wRuyBl0KRmgD1OJHlqJPXfiezYua69qSn2rK9PVLC2kLHhK6P0XLr7g
nXScF01qpWAL1m92ByckFXztPs4u0E17e1e9UDHiL3gDxExrofM1CeF5yO0fEJga
CrZXjJ+wu6OhHsR2CWaGGlywixky62TQ4p2L07T+ABP3+R+iQejSHQxk+OvicOS3
k5XY/A/xfFBhsRlAmvEmg/B2stR6cvgt2cWUBRStrjQ/Nzv8gSXEwlI4/UTUkx0U
eoBj7rkc914q+G4PextRIiZXvkGHItuqtpL+eDOIrayXXz54xtg6NfOnDe1Bv9Cu
kS56GFViE13tP3P0+anXNPdXQQSeJtPotp/n3eUW7zTy/Y1Nk97lDib0ztyFLovR
uxdA8rBW8DkBhNIbZltWh6/C5sIqeybZiXaHZaUBtTQf5+Q61RoKODpt+2A47TDs
up0tA/z7k/a0NtavG7T68xNUTJnjjfe9CeDK9Vt1gqCP10rR4HZRET1lRJB/86fu
rQMGo3tYdKmNWxHEYMbx1DxMYiasSJAy3s/Y2HkZBnZm3578Mms8mH6O1S5JVIwN
0Z6DwpcMbmnhHjdR8wGN6xh/7kPriaz7qiP5Nni7Ds3VyI/1TrhEdsnea+5Vk8xy
bbUVWCrKH6oCx0r0WIANQkCG8rmORpKM+j9uVXIlRxm+KkdTK9/3vvnLJc+Mfx67
BIF2jNTGMUZpavjZMfCA/UcqhAOQn226H/Bke4eXJ2yOBS8lc5jZk9xxyA++G2Tf
aCunMdtVbICbQl4DPTeTVJljbnt8nTH8vq021/ASV4K8Dhn5fMRmyAzAPaFPOEap
TPD6lwmbz076ocHXLvufFVDt3/+qBMWhC/chUk24SvWxf18TIr/3YieWfRTTHEve
YWkeaxiBkijPO3a5l27RTaiZ9VVIeFCkYL6DYXGMZywsoA98XSSO8Z2vbVS3vqD4
b2Z+Zxb3oVUKP2skuCbg64whfgTysMme7ocKLTohj2VDrtvS+wHH7tOb+QNuZONg
EiOeW1/y7wY+BPC1KOtZicPcd8gVaS+OUg0hIHPEuPj1rgH1EqwPNITjgReSLT/1
mI2N6u0o7MZKspBQZuFM+FX0j/a5eQxfYjTie/TQmcENHXNcaUAhRlHZPfd8XcFv
dyzwaKs3ETB/111jgoWWqIk5gux2bLLn9xMuOcvbLSxbXZgwJMqK4v75brW0Ed3v
nzCEEinFmwxbE1fPDd3b5hvGijAV8BYtvs1EtC25DtZfPcimWYbT1m/GiQJGbdi3
NtRCszJdPWxaLhLE+zC9+fCAzfeKeAIcfhXTkNsh899RsysYWHCTJGKZFGKeXu5n
xaamYYm57NH1qBiWMwAmyd2rKUZL7S5sCR9iEwmOX+flLZHfSVJeqmYiUBe6+hGT
3Wh+Xh1GupukxYnHZzki2nvEorOyIVSDRbmv7j7DK0gMWAQrCA87ikHsCWmZXmfE
FRipx4oiC7n7GMneuD1yRCQ/EUumVRyjvBJxK2Fox9uP4rCz5S/XS5tQ1s92qoaB
XximA+KZdJeuscQ+NfyxJhGNd003gmBQRaExCjI8vItQMMN1pqp2cp7pELppST3d
1g7aJC1r0//CmnInXkiRNDrtK6V/uMlOWtyPRK+s1dcXdokpU3fm3PrkXJtGsZwK
zMCDngTKTw7NRX5K77U3TBirfjMyccWkdDPHTBsUfahHRDsglCOK3ibl9tH5tEo9
OlW6GfzEO/k5SVPk693RTwm26PJtTOki6JtEQ4eoZ2h1Zy/NvajJY7gcjeDlfoqd
/YCZh0xOpnyuy74uQ1qAByH+ArmzYGNcuwPTrrn3/hA7n7ZCDXnVHyESbvOTp9gK
a4+yhAyL+QCN/yfH094gE57tD7vbzywI09x0GKtoG3KuDJVh+HdztBtkUQp/kc+o
sitOm4udUZnFEbONPgmFLGCf9TfzGo9IWUM0wk2/kx3nUe3KONo4q9CA5wU4wVOD
yN0UjdLszEkC0zZiBSqnZW/aVIGb2DZEDYZvxDnP1NyYWnHmL6g8DRH81yurYpiE
oRiJ2IsK0grNoplcjhs6zFYu7abA7bXPPhKeBqY/4/6xzU1GXA5NrRQ3YG2wJ+1w
c5c/fkmJdMCX5W6BWNBWhaI1GeH0JJo8JRg4D9YSbRIWsEnyLTfdpmX5FT9burBL
DXWmY8Wt5NYY32tsuGrb3949mfxKwnjwEqchYgpFwIIe4g3dVue4svVYWnS8VLrt
qW/7rWFhmmT+lk82HRaXZF518HkRqnP6cG7kTt+D6jikanABGqKOOH+NAV28QN6r
Lrq1upooipDBEbpj9MHQZ5oFkoKIIdeegBU4d5Hw88IZpN+gh3nPsv+HeW5NBBeg
q3rmN2HPqNHqCjudLfKdK/gvugHoSPa27qdpbtq/kVhjeRzx6X1IwWuwSRy9ycXe
QFsL8Ht2kwftIPrMKn0lIikwo7pf16MtQ+Q8FmM65JqA17I+nAKk9JsgLemdDnjE
N1WvrHIiuIaK4uQTg7Jo6Xrcyos/D7yFKC++7eZ8PnUDB56WxN+8i25IpSzbCNZL
LctQsVEQkkT6YDZtL9qaoWBnAU2w9B7cqQO3UieWXWyJpnrwpCBzTlA1T1HBL34t
KP/bYlfXnZWiOxyNyNkfQLzJX7ZH4+xv48WuH1aPkRLTMD3fkycR2LEAiPQe/wCZ
c4sX3KNQNXNmsCe26NXj1Dy/dpwhOKmY/emVG9rL+vON7wjFEALhG9/kUmmFi0lh
FLuALf3MqFYwdGcRX6bFckllb6gw69veNdMCe0zWQZ42XBgyicPuxnNkuOWshYkG
ESCRSgL5KX9UWIkYnzWT5KN0foVMQy19d0KSqIoMmYk6GTPFgQjwd1iijJvTvC6X
pCISm7Cheo/dm1yQOOrNaZ6mcRD+7nOJvgg38VmBvRdpOXHDEbCslOKExAABNY/Y
fGewXJptoIQhJ52W1jH8U5yAxnZEkzp7nl28Qh5+U1r8EU8P+UHw8vPLtELLeN4z
sr7OQndU5hd41hlr8j9vMY/JbBcff3g0uWZ21pA2famlhlE88WBXgTUTtu6J5dBc
DzrRDOw/jb7tAbGl6fK2iw4rWBij1i5PxlUWpLxvVsqE2aR3vO182EGmoQIGbN0d
AyAw8I1q4eb3F/4z9GmrhQfh1mW6dJMwr1W9qd0P67BbuwmLZlSlnw5JPo3v6f0c
fr+ZHitXilNqgLkzi0h7HW5Jdnl9ddUB8k2dL6nFtaCd4DN4hebwSJI8Bz4doZ3E
ZswwHakEcrM2Kg35wvu8SN1scwD2r9PiQOWgl6ByVs5OvCVOxruEHD4k6ehoUDAh
+FYd8+pjhycPe8pFKjd+j3Y7R6UNpWA9ojocj1sI8GokHGHlyNrUO8E1t6L853gb
OiONRLbhka/qu0nB+ZLqxe5nTv0RYabiF3TBkSwTCmdV/K5GGTUpKsQhPFf8jcaI
OmKOuSvtKops8p5PXyhl00+0/y+OtEUJZa/aqv5BCuA1GHBdW52heRZMcAY2AoKB
vgSG4EGPh0VHtLDvzpuKrjJXwUsuk8pEh8gLdlXegwWQHq47PTg7j7WtcdV8RByM
74BWFwylrDyMC9OIxrue6R0ZFW3zcOTlH9nhc8m8/qu9KVA0g/Rnk9HLm5Eg9Yps
vkf2tlrfk06IASBZvKkBNd4VcRhQpx/BwA9lVLdx98/ItcBh+wlfR2OBo+adgJFT
fpjBzKw6eV3pD9HUqYUU4M/4b4gSsIr7FZYnNRCvVQGD2rZ/AVssZidm39NszXGV
uxrEed/PPNDuCwlgShALNfbuqGP0396/nTavFKl8IrYe5Xo0jR/kI//q18WU+pen
ggJouvOvUbWOe3DjWwl0wGjWKw10uPmMKMmPUqVNBQAtZV8cya26sW1C3Ik3NoUF
bY9fUIHGg3O8X54mDW9t7fymL/sdMrPWN0/2BCt6VI0+8avTJ7Ta0OeLOfX8JzW8
cyGyZdtr9kBWSQ2Qof4uZn3swTYw0eyo8MxuJLek1cQnEvi1OIThP2lfJh4SHLm7
4JRzmvGHXANtQaIfH4h3qLWnyjUkW+WYDOA9njF09FdOnPXlRBf6k2xyGDu7z/kQ
vIxw/GosnuUkBPHL5/ZQRtXQMswpfSlBkqNmP0UkTBLRpHnZcPD/H3Xi5kza6vgw
w/iNKuFrAFeub6cMnv9bQtTNwJjBLecGIYnydzRYjciuy51HJQQg9BDc/YJsnNED
/pvCjfoWFkKnSmAdnHuS07zweltg76JyQSCaeLZXZhBARcXBmdGbF92Pp7XpPG3d
S/gSUCqGi3wIqRyxHqdaLQOfKNfX/VtZv7K0bWfzvPwY8hkc4TdlLqssOuT0rt1j
6hK+9K06aVeDw3ctNFqD2tKYzNDSwUiL6WuWtbDTW3dG3iKnS/vJ2pGATUrhavHd
enbhAQrb3aSHc6NjRT1I0isNBVV+lmE9308xnf4Ta9cpdNl7lLxe/1uxQrGK9J+9
ESlILNmd30YB4IKgRoEPl69LXDZhnN72TdWsGVliWMz7sOAwUjUGU/bxySVcSLrG
gsiCCAZJZHt5ws9MbBapsI2iA28v8EPbt++3rSPKVEN9DMIo1JxAE4KM6DOeXVX5
5oCtSsLMDqO5qQpW0MNabef0/0MX21uLX4O7cx2R6I/djPwBoBesI3A60EtQlZ1j
okFFEipKAWw+LP+IvGyxfP7vTRn1+9uJW8IX4+nHDCjKrO8gEk8A7Hj+nZc+LLfE
iGjdVd7v7HMr16VxUKi+4e+bEpPQEDSh2j+7bhHzC1ignxKpL2FQyE7iSBaIA0MF
6rTCANXOC4t/Ay6WGSzQ8T3PHihKiiP+mJoYhVC6le001tdH2ZfykpH8ThUB3DhC
/bI9yhl2/IIhg05rmgcTaK+Kbcdc12n0xNYMu3JYIAdy+mibuFa5Wz/qkOwrdnmm
Yr2flz/ymPm6HksmbbGwDKr4SA9CrCbXEPVblTDrM77jHr4D7pDYx3ZmTfor/qwL
GN9ogJAKsPulmtk4LmJqA375w+UkXEufcrE33/SCDpKn0XDXtaVpA4hBOnPhFfdL
L5in5jxSgTe4hrXpm3yKdhqfR19QYDA8dkz7xymFkahpvUwtNt0VE5d2LoxRekO6
FdxIS2f3UaNZEfMA+xlOOaH7xBVvlhBV1nayPKUgG77T9cfJLfzwY+6JECHlYq7M
kjo0TShWb84sYe0wL0S1Ph34cmNmKSpx2SahubFyeLljPs70K4ntW/7XzIn3Uk/i
QlInUBe5omEWnogZxHmYFS07qOVo0Oiry78QGho+iLSuXxXFH7e/3VkHvg9cJn0i
oFUDpbu7YTRFzBFfmgY4sfVTpIQB/zrMcrI7fX+cIu9tHKJC/y3klihctu2X06oh
hVnWOYqsaeODjUgaRXhA2Xv6qfyFngn3vmJKiZuBOgbZBrgf40JgfxEwOoaP6t1j
MOjmrwCUndvsso2CEBRLDVfirkqPtI4dgzYUoMnvZ27LRemr+7nenXaFvm/VKgz9
MNyGjcbIJHMwsryDaNb4T1K1J4zYf6XwDPC5BYVyhq2sMGCNCUVj5gRo/sN/qK4j
lBKlKOYIWJVb1+RO47K4wVtLUvY5aIkIFKN6EIBEBkOGCo1hST71c+sKopR164Gh
O4SEKa/8mWwXWBIAiov/ZH+V+p8l0LBlp3ndCIkIfjaNxrlaj/lWG2yFVhiG6msR
LtluYCo9ksntZrQ+lArMZTEZJY+nnAmCOiNudD16aNtdQEamlCtUszLtr4gWL00/
HHq4Ht0HOU3+4JpcoFakzfygLlOftSbqfNISoZJSwwa7LNh8vUNf/7LHIUL9cZKq
U46Wny0Xs5OY6a5cGFLrMgYgc3x0sPGV/uB+4PZ5Ymm+kdJ1xaFn8VNxoWLkedoQ
MdiWp5FKpOMagMQXBOmryhkyN0iV/csr22isyJFgtnHXLFI0fhPGT/WGexKkn4Ey
KyVVOKkhvnnYwC0ffsIvfVBF01worshWC/PIBmB8AbxD5ZgkmXZPf87l9XPguy8p
3kHvUNMbv8F2FBqDI7am055QADlw+d8u7EfWaQn5k6FUes8IG16k8xcl0nGQy4zA
wqPNDbjmEO4UjlXwT6QR0LPK7XxZs+RpKFcjDOpTQzCji3A/Gk+18u3UZSKas7c5
uURhrVYqeioHEsHGMaRhvwrMDOsh5nx448xfTqrD4sb/ChbkMweWNUPqI9N/2hIQ
F2kMF1l3xN9ACWTTfp72EP+ZtxjE4S9wmHXuJHC5//i4BnEAglzBHDPjrBa9eZPE
QixEtFMFnUaZYcYllRjYEUvwn0AMIT41IT9VER/1V1gSu0bURCRF81Jny3l9Rknv
pjeAg72ODP7KltCplCneZZZU9vQ2UqXKHWhcsRkr9HLxMHmcpVsuFUpizjClkEd/
3bt2M8lwZ37cMYnZpO7lNRVRfi61USWWJfmfumxtvMsqa3YzkNPTbUv0nHDnuL44
GrLqNxi2INq+k9eikQMCxpXq1HB7Y6CXaK7Uq+Apyy/xSgsvW0hcDZOoaFI5LHB3
1OYFHSLk5vKSyLaMdzBKHGy19z38ob2EnZu/8y4LVQd+Pt+2F/jrC5Q7L75lc7nB
9w8e1GEqQi5suVlPv8yeEp0v/n6xsSrO7/dfcPeuDwLzcXyrtvto5J3kBtpV9ocF
NV9VlPni6Wd2X8skU0EzGy33UDukYvzrT2vMqkY12FUa0Ch+420eqsm93Nt3EkWv
LAAz0ug5U8jYUa/chBSbJ6anwaGWiWOsi5GRdHwgbEq5IH5Kc5t/15qlRqyRFMy8
68H5+ilfujpIHCKcblujabBFm95pm1kVnY/CLUCURy7FueljaDk39d+U8lQxcVAu
40ubArIuISjWzNWbju9Vji92peILC1ILaXv45WaDSfs1cINclbehCiTlsWa8jCkf
n/ul0d3b1Ti5RJ6sPCwT1nftrxBJEqjFtub1gVXXAUmhpGHuckDYjn0TkZhLJt2Z
dMuUtflYeHyVH2bpMXhHEcZQ5AyrxXdsBPS6zxWMRJ3kB2oz90p1ztEcdQxGKnFX
i6aFm3hRCmREn/TAV6aJfrHbJDUA12W2dXujU48v7wvnRogd+VVbmneq0G1yEOp1
CIzH8ifx7iiRQZ8TEBAyRTh3dv5+HXRjRC5Ze8Wp2bUD6UaIA3qZFntiNoQhbE0d
7jgHQinhBcuAgZ+uur5WsDXr9aCOuDS3PH5O1FBAxhbywmsC/UC+SBC+Oiuf20sD
JbgJfjOzr2T7esk4nZcG8AqbIvm183PcXdZDNVNwgnKoP5TubaA+dZP24HFhpBeC
AulSn4bctg25Nnrttos7/gZtxtmZoFiDnuB6Kg3LfX55ZgnA5maM16OLlMkqfiZc
9Hg91BptiiFXMZy+lPOfenjT8H+WQTVZLy+DiOgw+z1eUOJsO99NNnQyK2nC6eBY
YRJlPXuXkrYPQE1UUSdHuqhQCBrlVdizTvpevL2PHQNtNtHZzYonc1IVOMZc0vEL
C9ZtPj44Zk90JdMxirbihRlVdj31RWcXla553y7o2XJ/AZ61bPEQCbfWLoLoUnsj
Z4ulRiB+Ld8VkGbqvBoeoq6Oi2j2EjjHrU26XYBwp+METz1DUZ+wOMs/TmuPZkaa
8QUSJrzePgOBcfDQE1KEmtYi8xkFtt0q1yNndYevFiQ9/QqaOn1csrcCeUwhLiCL
QUBKKYsSc3d8OW0VNJMHREGnkw/dSevq33hUfGeaWP6qDinMfg6Pxy0FPwZSRqVF
SQYeHr9N0PTWryb/bzinAZDCk42hYk9SoycRos5wfTx03gNPRJxPrp6JucQMZ0jT
WcRrugEguXk6BI+C0ZQcSPDsm2YdtHZuu/TaIi5QLje6bqFaguFg52PmDcw9H4Dh
O4Z2iAi3eric0Oksm59kpOMS2XhiIs2mNxJG8Nrhrxusg7AaAvCd4PwjVhKWlTK1
jaT08tF4rOjGnLO41mFpyVqLMMf2EZPkY6Ud82upHU6F2WWAypKxFYgVpy7IWrVV
rCviPUeMEdYAn00imRvVAWbt2KNU1ZYwN2YB4s03FKyBpQnoL2xkFt7A7ZJLXgKy
O3zHUIbdroxp+UgbIPmuNKH9rEeVfnSSPTOOhi6Ja1jvRq6BvKEkMJWxwHqlPrJ8
9Ztyr3mal977KUeulujBXpUqrUfyr2Szkq20JZQ4A6TYjKT9TTsr+ZV9w8DAtQnU
uCfdZ6KMxlOJrwkxAuf7dRsFDaaiJ/7Q7s7kyTMV+vJX3kGcT0LCFPC0Lkz0x3wV
3/OuuXik/YAv1lfFupUgFnQKO6/XbwjAcZwsBHao5yIADpbm6wvj4xWElqS/8LxN
QMpkxWaLVZBsn8LDOsTbCyblS4ViPzL+H/IcdbXv24wWw8NGRLEKyNLU2pjEShvz
AhY5vOeloPW/UvMnh3tblRnjJggrLKmdKQSwGb4/WcmvW7yG2ZqxRjSXvqrbhfD2
PQA+VPpGtxSWaRjGuN6hzdUVH1xEA3yr2EgahhUCKb/WoMgTxifow7Py8FvCx0ac
H52i+ip0u+56Rwx3+MjXXqqtUi6T9swlDSZPSCtut5NLHfJteQHZK3eXtrMWlmEz
+71E7vuyiLz3mHdwpEZQAN1PnTz/hXUYUoMaGLmICxB3KfMI8GbV9xaFZie7wsIJ
KfG9a4vTfyOaIMUKi7but4h6n1XYOreeytnoJn3bsfLyyYAO7uI1RIbm4LDNycFs
UCP//+RHEZgSOIPAun9N5D0C4r+TFweTeouSlkpLdgiZ2HhNbeaKmsTfaEDTjvZT
8jgqItAijmGL0Ka0UIvTw4u6WA7x1Iqz32Nr+//8D6XoRdtgya8NUJEzj5r3MX9P
6Umv4eXUFPZb4AfwLutW60kneiek9ty3P+3sLkEsvEwjn/pwWizexbKeTh6/P+WK
TmfrKPvhMh5fFZ0f380HT2Ceas+QGAv3Uip+ba0Ih1NQRqzVs1PxL77rRUEWxmD9
tjt9oNTmtfGq05CdM+43kpIdiR5i6AIkcdusiI1mlEt2HOU2w+P3/82jyNKx9ZBS
GhWscKlDe3AQEBCRQ0Eb7pUlIyvojaUN7BXgwuMorH5zIvfZLehqwPwODEa/UnSy
0SIyNpq+ti3mWl2jfjlMDfdKpi5zyKNNb05bjND6SZcVzBUnCzZUfd4HNF6pSIzN
Zj8oDrnXNZw+oZpWdkIAXAolzzIjw9C/zP3+7BNCzBJbNxGcU9kGUqafP2uLiYjZ
6wQlXcVKr9gQ5axAbc80NCeEK/Lhy6bywdmxoxlPxVO1bxdfqDHUnhJqZHEHQ+Mx
oPXA9VK/W27SPTKJzu26V0hrfVYo3MAzXJo6k6tK8ACBQLCbOQbSsYYnisfrR+wo
vJaUcMdMfFr8li1/LHbzDUB6HQ0/K7CDQdivfG2YtojLDI6PkpkiYfrKaX/nSVm+
16jpEqI/azQM+osHtJxVZqaBlt23SyNQXKrbOiXB7akyhIFU8fl9+NkC16Cdsegd
hCBc8v3UpBtzK+VvaeIgPgiuqrFOVstXdqUeYRULqYRu+drxCIP3fQ0q1A5+whYx
TmULkxfseSHJr25EB0x5QWHf/l6UQywxNg44oLfgOY8A9W3vo8czHoKPtVXMn46u
qgsAsrbkt+XvedIBJv/kbOY5akugDmnUXeOjN1w4mDe/0NGHsJY57ScWFQPGI5v7
gvGEcBeZ2ecGC3ZZi+rDR6aOFEmI7uQKBc4VK/u+UqVSNk9V8KETUJAKw6vQY+tj
0puXlAbxOTpFwOLMROpS5wl+wMQz7T0R44KstQLGUHGoQzf0zci4/0BQnnBvkbjJ
5IGSbz3tAAdguFpvgD5dBxDDjsyB1AHYfCQOo66pDJl9yFUz8mO9kJbKfARbJ2Ly
zdpOhctpIfFb2C4e9n55OOYrDHfUEj+mUu7NQDGJxqjocxXtai5lQppSUfMD5Ph3
zvYh+w/mQ+mkSiyou05ZLx7Dh4QUA1chnkdesCH263myg/k3BEjs1Mr0xxdt9mPX
D2+0JiSaClVE/oONwbPxhdg/uKPNotHoqbfFBYOUywK5z7Sn45iqaRHTcOh6MwEY
jq7tAAYirQuvJfIoKZAVxVVZTCH5qk3lltQP9YPZ+XwUdgkcXRDwSj/fQwfihaAe
Fmkb75zYrNf52CkD5mRmZ/EL9o1e4FVTM5hnOZiQ3N7ax6LxevBKpxlij8/oVD+5
P7CNIJN8fHvzXK/1shcJJcWyMsMFzOhrefTa5sa3ApNLqtzbUOE7A7+Gp6oGNwD2
D0YHsquDalN4sKTrIBQ8D0JHgwYQuhHOVSTIvkoUlHybCwkqk8pQD+TSk4iVlsn5
pbNlQ0o7nlY7Hx35j3Bu5GpAQorarBCErr4tkroRTNd8LvPOxVf+gOo8TuzgAZSi
vA56OuL8ogLCC3CaN37YJ19oLKlsu1VnZftSnFSjvZbw5tuxJDtlWblKTnk1bHVd
cwSJ0FrayqldJ6ZSbAxBA8qilRvolXaCU0xoS5Ka4WjZO0T021QWD3IilVNOQPAS
6TnuQXa7nx7k+d9+C3gSxvPiGpj369gra1nvTqIRSYGBM6zQRKIv5DM3w8npdivN
6V75DleDPX6Bo1mkDhz2dMfq6Qp2THuXs7yWe7/+moOZHOvQcj7lfwjOeWhJOqSi
AIW6Ifs8VLtIdqS1S8SAZI43fjsg6YQe0OfWAooaHqrkyT3HHX+rhcLaFGvBAEnm
KZxljvixkRNJ9V+YhFQkgEOgzlXvCGnvVISpiV69/H4dDXO6wiIVK5yaMpnsj+oF
4zpJuBBaxmIgx/lkdTghCyuy8bW/0IeYcplBStIKM4eQfnCPQtzhbdS46kRI2xWf
T4oorzY2JYBjd4zlaa5Z5gYLtiP9kxiI3WoWYqjUnxVDFTANWMD7hQJOERpTPtQe
dbQbhbUxvI6cE78huidGlN16PSQID52mL85yZuGxL+3iUyWazqEYfRUmHEb1MMLV
1VlreqK94U9hUtDfmfyiLRz0PLiZbbccWaX3O5mJOus7PkCd//If9/yo0q2tPKcf
lSFqA2tuLK87R8SjlahNEtu/lKsFPacvV5XHh5fh6r5Jx6oZBh17ml5EZjLGxjac
szwHOYPSxHbryLRF8czh/H1K8vgudHolgrxXEMhx/aorOgQe6PMDiwHVfFCu18WC
Z+z03KwFeQ5HaMHA+v9Jvjfwsz1a52EukUfNKMhVdKotfO7B7WNbUWNAgLKnvcEQ
yZDREcBn+gHkgai1syuFORhgmvvaRjpi5Pl0hGFuhZg65MXNo8ymW0f+q9WmTpdI
eDQ2ZDmwuxCPiP616UTOsIOgYQoH3yKkpmeOdiOhVBwXXxbxuNhk0x2mBcCm5FKW
YqsxrRF8ZHyKs6KmMaKrPq6cdNk1WWIAZ7On/nIOmUefR+OLoJ2W0e2NTbkI/j/+
UQohAGBTIO2QmseRKhzd+qpQtpP84Dtlf3nVXvHJ8mhULhXGE1KsZEC2l7tLoAEu
AmH8zlA+wGgC2Kn9YEsT+K/q3DADYyfn23KANoXpDDlUVUtdMB/YiqES+nMpWISv
qoaVFOIpwiBW4bZ7tSS+AR5suepw082pTZFVNVlMa0MvNW7XWETF72puWGHWWbof
11ltWXcb9nO9DF9e493GCsKSH2ieoMpWsWc5GpDZCDk5MmrbpWWe3v2hVy3CslVN
K6KZMa3yZ6X3/oqdSkLIIXF9xvTcqmHjxbm05bantr3QBjcdwF/Hn2PUaRz+J6Fr
WY976LCAKCy/xwPIIWZ5STkWfCjJKgjwr1Ix+A1JgaW1AvGIV+rBnANfKmPIIX1y
SI0R8+D4zQkYVlGFamu7tk4ESUL2x4yroC1wzIWdncuxxqsJ70cXeYsEGPVy9oT9
/wwBdcIW2tBurZADKgcqHawnPjc1PzeAFIV2ZDRIjKuwK2f/pZcOQvrTGT3DpN9D
48ivN7h736ME7/JtmC2xfLXWGpQYhcOkRMHLfuN2yFiHzQXLvyUuL2TCIcXoQZzX
exqtw3swnEDeuxRm5UOxVC9G5plCN4P89GyWau3h/k9dh/HZHKoM7GDK9p2LgYy3
CdAapjtz8dqUozmHlYFQ5wFuhDLE6N51dzVfPTlKZhXmcSpJM+9n2utWTu93kmZX
necrPfRuXwFCrmFZQ48hUI++ZivNLnRe235vjyEaxCKu0Cofqznxz8fgydseAjQB
Ts1W0kV+GqTHVWysGStJnxZEbipQew+gYJEXHY0wz3Kmrnf8RoD9E1OjRLhZVml8
WvcsD5GRn0KtFPRpl3cg+tT573ka2VO2fR8PYKIrcFfgDA3/p0np8GM0luOazE1p
f1jidp39x+HB4gQblKAU5oElUFdVenecOkEer60L2TcfsYLnxu8X6Yf9wEgBd3/X
JXAv25IJupoZ0HvqG2bHu38Iwo7PkWkXh6GYpXym0HwD6XLXx8zkOMHCkq+oqJsu
7JIPowDoDJBUgDdQaYlZRdT/gbb0gumoO4dY9EpnT2AwZhK3tNmsSfzEBD5sN+ns
yspRJ1tC6N44zLDmJQmUFC62Kmf1dArFXckh0tp3rp9mkyDLS/10S9V3/DAnn6Qt
+73aRcOXN38K/bV5YkMVKPxmOvw7o8CiA5dUPC1sUQCYS4KSKEC//QIX5CTbFzsk
ygfw1m41tC8zpu6Pn+HrsqgKekzKHQ65So8w472wIk36C5qpNWVTSE7c8pw8uL4e
74gFdR1kBYC3M+olt60G7FlVE9eFF29Dxebgkb8AWZxZ9faWao66mm0pCsvaGHce
2w805vHIrXjZWsK8wEBQCvNNr48BCIqjYOG1QJnB9BHsiDSkvsmfD+aAzKkGbGoT
soBfPzy6hkUKxzmgPIh5r3yAwS3LaMbWM+nji5pCMuG43/1y/34UsX/pWBovit7K
+jLIMgy4JtS3ikYPLhgtCUk2YG+B+RdxeCLZ5sWst5j9V5uehCeaKW9P1f7MFW6Z
LDdN1+zWI5S/s7lXh8/a4P1sufFU2shVq6K9S78Vfw4cDu7fpAKCDIALTqE69xMe
ocLN45nu+W4IXuqw4ohgBjtp7Eajvgnfh0rBqUqzQLOULWuINS6nS2JiQfR0HXd8
XN/P/muZT0hVyaYzSJq8XK98Mkk5D0PE+bXtxDc/IpaNdH6kjjCYJP+qjY5Q1QU3
xjJkc3atW/dGKlXQW7GC7BZluzlKRgCYRGTrBarA+xYG11mwPNA5enhLzzAyJoxF
ZJjDHuxSSeYCF1CPVaS8pbp6Ex+lA/UdZiAHsIDjlKn+zNwULJtRYa3Fui6NPdYB
iFieMaOENfmXQBmCU0rq1G6AIP/AmzHF+cwKn+0bn27KRk+RqwPcE4kveWS6w+oP
6PG3k15UBt/y4MGobwCaVUsn34dV3gyw71nGJnAuznJcO8zEahNFAv3gY69hKEDd
8ROWfaZd6ufxxwGYog5e4TAkqG6JJNNi09RJCGpAB/m4yGNRvsZbqUNMFA/Skb2K
tHAoi14RFnUh0CAqDn3lsD+aXUOySNC3NFlpRlLNTc0/eDhYD0k1YROYYK9G4IBu
noRHQCGf1MA0u01auk299HpfkTCIKW48AAr7RJvctSUtctu9CaxIzugQ5DC6ZVUZ
YTBOhkr8ED5x0NQYb3yHGjMZgrXjOgn9Tsm2f+OhzLwvxz5nJ3nIMlJ1Is6RrzJt
u2YFlXTPg2VEqfXx1ObxzQRY8oAbQDeKpV1AR7de2Qkei9096qWLUEJEYIV1SyJo
6U/9CIO+R1SrBdYSDL5PklW8Tx4beU7li8AlUfSokhBn91Gas3xMjK6E6CRaJVic
aH9m20wGA8YkisJ4M5jRS12HW91wQpyurjSWe2/SED0Qp8ygVIkupBOCEEcMeOVo
2CalrCEkXOSo8w0bzK1tTDLzR9GOFtw15qnewZCtDwHe99UoW+x7zIiEWK1gr26S
uHnjH+5xfPjPqV2FbzjkGTnTIcODc7Syan4KJRlFNzpe09fdIl2iJ8iqTtj3Mnxb
l0upK+SlbPSU+vMghOFbPmTeMVB6FdtmFqBeYTM1Q++3742RgJl4UQi/hhmPKQgB
BSBNDx73tOE3rOeRINEQoVlzgeAvhnl77puAZMeQlWUEU8cXnhmgsruGLqTutGX8
tTBPuEqaQzM8qKYhWo8VLiCq9uL1MwVxDN8hcL3ytWGaBETQYLbQV1u0yy4cwH8C
f1JNQ9n05cTbwVwMzbI90iy7exqEop2olyH9B8z5QUTWJdnW8PibKVg3vB7awbnZ
DASmuQ++cJLHVKKmdefBFmAqm+A2yPU36q4RWWb6BWprTGTlgaPgZndXFrsJJfZh
jOLe8360Pmpe2y/Uk219uL4bqN+NbTOlvjiSH6Q0Ssvp/AJzne0BBomcrjHWMK8p
XROYIvzfX35la2jFkW1h3obFQcpG+pXrQ9KjKfUdLFKTfxSvkC00jOFKEDAXgxp5
d0Dx1qATgpsg383zAnOVr+JN0UQIvr36JggXmWkVY9TIoKCXsv2ZimpJEE89Oh71
CdnHa2fY+J0nd6/8sdebqwKBEEYwbchEeubkBVS/JRFqY5wM3P7HS0qxRjw5Y1lf
7ueZAap4LD5eFhgpGE8wuee3JoaIaBuLkvD1SOIGo1xp/Hm88kd50MFJsdv5Ge6l
pJ+14/DbuaKYNPDOVOHcCRbO0saObHnV7IKT2Pd3qxO7gD1set+HyC+KOv0yjEn+
c8u7A+Csh7cYExreRxfV8R2TA0IF2SGoQJWDDtMel571BWwi7PTGI4aVN44qkuYz
3I+zNrHY2gHPdmFcSGYOFzKiTghrUkeoFiSjhBmhm7jAUQv+3zDFgkw0WLz1+XY7
ed7Cxr0gJlnPVpqqnJHN538uPu8Cmpae8c0NaG9jMsBVmcSRoI+MsQuGz9pnVy+d
T6HkSiHm6Q430tJ2bBOJJuA/Uv7wuE6uZAEte2NHzu1gOldGHOmLomNN8jEPm9+n
59yj2RVMrUVI06njCVEDdZRwTakqr2CH6GfW5o3L6RfVE2hMKHR/oUjttsir5Kfd
w89EEM2gpm3/fRisLcvZRqFwcLcgInZx+xFqverZpHd/uGoi4T1NxaB4q3RWweYv
4CW1P+57e8+D4rPH7Zne75IS3JderQh67AWUFI8paCx5AbR3YQ2le01eV/+UXtcr
uQSqkmfPCxRyMWwyDYMiaKmB8uheV54ySbphQEb3AuYDWeycP8vuFbjO0vToRroC
IPPZFgnBPmcF4N+Ko4CoJ4AvCy32H6wn6i7joChvgFWaBKqePDPIIRujM5wiRHIh
1lIBNqrma1MhuiIlQFZrqgpAll3CmNojpJTgbg6OAc078l7dTiyH/xSrUqQLU2X1
RCSs/qO8iR0bO4Nqu8S8wBeznTktcqCfR7JJQBkInUMftZjJvKwjPxqMH0eX8oXD
cLwjacT9fn15oblqtpJEIPe8MVFCe6K9tDhkuQmX2e6pAEWey6YYEiZm6q9zCn47
u8wkpTTXMQ4Utq8TKBzU621WkE5uMI7zhU0W+7zLqRKKDD+KXYLT7gtrPDmfmWOp
FP7yqC7hB0xZxa0UZct3dV7cjP33txa80iBwp3abSHrd7arh2445J61B8JjwrX5t
//fv9atw7Y/BmaShmksMGur9ZOXCDNdOH8crVl6hD/gNlOzzMGjI1E8G4F439UrU
Yk3dTQNV+toJELhNOUvmXfs0jTyaM4GZQya6IJihDEklDLIWrL6OxfRUPcuOVCBA
aG+Wz0SH4RzuP9Wo5yxQpa7WZzcGKPIsy78oywGchlrya3fLX8f5y1W3SU/Z1SX/
l39jsWE6EpCkDnq1Wtb2POl8lKDxhJ9IZ+4etQpmJ5Y1Zqokg98rvcGQrW53FUVP
Lm7fcxAVTT22ag8QexP+7WqxSXCGhg4bmhzb9+4msDktx0DaN96wMAQ7n/n9+iw2
zrZ/JLkHUYRJe75I+uUgrHAHCTBVWc+ArohKjaewbYbCer/zvgYrBfGaw0TTieTv
S0CUlOfACpzb5Rri8Zd33tsqJ3sKgaVWR5hNuUIgwXpbscnbFyjdnlwufZ+ddqLQ
Hg0hgFx5tUL6TH+3MeYHSMGz3BtybWlacUBmwIgSXEpmVIf4VXRaf47f31/7tavo
72nMwaOQo8hawcJ2z2ib62FwUYmveg0gKB6083orFkIbvp87+c5x7AgphajuRuT4
VZICH8PQgijHUZX4cbHS7t7YN393Fdf1eCKGcH4K35TDhcBSA9idprl6FETsJM3p
wHVNCNON1Ng1tDAsQXWmvtFyDMcQXysXWdMoYkQSeD5FjW36tAh0iedf69mYouF0
/DC7dD1j5mj0hBOFiMV2x3yGVyoLTWiTSAWD5FzbyR2+mckHmcCl8N+HdHcETS/1
CinydQkcnIyVtLphDLj3B2Uidpu2CCeVYMJ63GhzrJ5QQkklp2GRSjvlPR4mMP6C
140LvBMHKjn3TT26QeZ5B5Gkh0gXYrKdylwBZgBWw6MLpNdFUzJuZvuj0gCeAv65
CiAwszkiz2Jmxbw4aDKZO5YgpAWr2jwzcJmeC6/9BWUOYdk2xFd0dIlw8uMwo+Wd
nSe2nxWeChONOvV5F8RLnp+RTs0GNCZrwoHdu12ncXJax9aORLnZzKfdz4tDg/5W
+JKvhGTpcEsqXXlY88gFO2nYX0T99nXyU4/saOEw2/YZJnZuu51sz85IRFgxbdUm
wKXWFUa1uZwyhU7dWACLwftxHMIpu0etlfMAc+yjHjGuPUedOQ8I4A905HBNDYd9
6WeBLSdfghnXBbk8A0t6RwDYY6478pGHn3s6f8Z0FJBHXYrjDN7ffK/S2YlW5W0s
TiDddhmQkilnmkl/7J7d20GNPoFmvkPBWN0v0Bnyg6AN6J16uQwaNft/wSZm1yKc
4IeZ+eY0LffSqGDMxt5gYhb0OhvFKqd3ybNDc5z1XDfCl3Jcj8AZzzhaOWAHUx+a
vNZ7AKYwS9Wb282BC6x2W+0G8MQogNGmOYFcvcYl75FoeoroQcOezQqTP76j10PN
Vy+wXBYPrVGua5sw1SfR+t8VCaMoEDov+gZeGK7flloP4kQixsrJ4uWi8Vl8pJy5
TYUOQSrEiaTrk8vIowOLoZT91mkr4LK2zPGPH5TPhs3DlIxlx6KGThqVniaBGplR
27XS7EkNoPZ0m+bcl2E1vPX7kyaoubkb/kPjILNEeOHomukyufxGWjygj2zPSaD3
HV3DR9ZBFm1nMbW3VXi/pe60MkCxy0dBGdpCux+nmHCvLhs1Hi3mqPmFk4YLJUg0
cwYVYmQ4ksrv7OMr4lORV/R20+hwKGvX9RWeL+ypZUMQkWfXtT3Ahj3qOhzzYlGg
8aq/tyzCNaT1Z6CB7PeNYzavqnCCK5BI3Toxzo1EK3eCh5bRpi9b/7fVbw7xkk/J
GWjH5gYQ2CYlgg7VAy96XfCfh7D+FKBXUwVZxTM8wz9jxvZtj7UVHWm4vqv87LMl
p99zf6ababbOX8xYkSDjR7paPPXI6ha5MJeyctKZq0v1RUPVzpv+TOnU88XJ+ls6
o2bAyoV3/s2yGV7IHAfUA+w5QcdtohkCMLFqc7ESL4hwU3jiq6+IpPZSD7pw07tk
MPMfXaJTiHcaRi92HwK+HtUYI1zcjLoWMXXGLCD/y24rKll3/8aO6fQd6jHLWI/T
VNKq4axOtJvr6xdgC2I3eBcrWTgnKrchgCx0PEP8NGc5U10zY1sIWgX8exKdY3kF
pRUBjXfvqr/+O4odnVWalukv5dQcbjKr2CtGLQ8wOfcnoVOSilg9Y4B/F/1Ims12
T5uArs5oARVNzbL7Dba/APU90F/XW4BwlRLL9u2u3kqXkpmTCMEjJNU8yOlI30sF
0/T9SY0DjrLu+qcbbcBRoDEdM3LDm51j5qP8iCKzOZ0IJzSFuKnFSv5k9ysBbQyU
6twDYoibAjnXk3V8z5Swis8+P0KxAIFD6KwruSYmGo8hX/d7gl46Dt38jizW2MO3
islA0NFqyt5LsWnRCfpUnhWhjPW7ec2hpHv/yJTN+6jAGn5J4+57Gpm8ed0cedUU
3pH9h/OW7w6q8GlrXc5JSMNyiDxorNPn6/b4DyQP+hi5v3ndGTBrc19FG1Ekk2Ue
azbIKjdWZAbSjLxEViedqTqp/TbP7fJC/V4vxubhom3jVTGdkun6rutCpFalCw1b
Eo7hm7sUIvoaUWTGlu0H5SKlXiZ6PsgFh8hIDzdTyOcOiOSgx2Y20fFwYvX4ocyS
ad7pwI0aQOY9CqtE6oAnXMojL5Rtfa+z/3jVvsz0A0EIWI84744cfTfM0VUJjGPu
PHdqy2OcO/VuEyjzNFL1ePJOgesH18JDQPb1wScVazMYeWbxCevvczyAr/u1HtOu
CWVb3cTP8uMOF5FqQv3bvyxCyjUvYskaASlcpnA7lQhzwWi0OsPClGifWeq3fLHN
fbmi+wKGdxsqf7epNCWemWenYf2PxHG969U2ZbLyBwU3Na+Nn06iys0RIVWIOgpa
PMZJXpAkP/b/zUqlZ1G9LCm9DUZOxQv5emYDV2IqV9a3XlvlJ9s/o5v0TnAwgpbf
5U8Dhy+juDHUtPPGN0gPX5g8Gog/3C7LATXO7LHnmup3spjxx4ApBsqNhMwlHHPF
ZMU31YGVXQWkrzsb5RCQeJDlWh+dhMvr2W9v3jQNsQ6fjqJ0TvtL70pofRdqN8Q/
TUuXeRgodxh+XL5z7yn7gF4U0izeN8VxUhk8Xn31l/I9j5OTMHXwRkwLgi66ap+A
YBQdCc5V+UANwPxK6qUBvCdTLimK+kSsAbXDawwjLpXYyzoHl3zrgf21htuEPTlO
ZhooTKvCISdXOnKaTj3FCrYsAsS547fFvVOpQmkzCkEkaaLgp2Lz/uX9+78m/k41
Ob8cvtTPeGehxWqXcWNgZsAWjzmhSb4MJM/0nqrpKNDydcjcKuhvCNczLPXd3/kR
2J8YTKRQA5Vm6Cb0WkrPnulXIh42CQIh57wmZXaZ35HjYRVy7Xy9o0WL/W2pBque
u7TUhjFMcSZ1JrToNnYvCl+UEYolRLal8XyITsV83KxqPP9PipLLIoI40FVF++xR
2uakYOav3ljTac4JnK3hnWUsjfwv2srstTKEHgZsSHlmQb0aN4y3yUSN8+5+Ioio
mM0h8hLrtTzaTFlT1ngpaldGfvUmu3wMV7vy1rj9mDkM3qg2WYHB6DKTixGgkIUl
s7IEXg4XRlR6IDLJTqWhuY+RLxslofqMhy4hGlsnSus0eIiXApiNPZAMGTCYw17q
OalpAozSjTBYeKGplKkHc397OTcfUu8FExkF+Rfb3ATiT6gO8lBEZgtqRUGLsonZ
vJGkcN4S6DqBW1U3HbqXp4nzeO0/XElRjIrWhJYPFXtxUH6VW6QF/TVdD010+9y7
qjgqrxN0FowmQLPG6R4+hy3RBCeLqNTwdrFd++fssHtPHBOvP9L8UkzyYgbPquF6
HZKW5uEFDXw+xyIKD3oEg8xBBgxOQs3Lbp6y08YSaG29GV6Gt19i3949c/Me8hDZ
si9rP9OEpB83XjkhL9Gqc+shWBjY5+HVRLINmdzAStgOXQ+VOlSwLdxOJt86z+XY
u6cUdul5uQeNSTMSt+SG7fA3lbnB5VmwXN2egHPdMbuZEAuTgsJRNHJrkTejTJDM
LLPWyIGya/trXt9VhbBwl4bjUwZQEKv918F2zGud4zOgAKGuXaAjwWNXp1F0k1R5
6y9pWYdkED2cIGEKkjZ34azYjd1srkFFn6RB+8+JyNaJJ5RV5rLSSSwMGxFvXqSh
4uiN6UiC3RI6Q8DntmNvMd4m+HQqWEZHzDrjEzRcDd3vdUE/MzD490tpwiFS4MzF
NlVYuPc9Li8zINx0pThLe4J0wx7NC+ugPQEppMomcEJxfamKa62P2Ndh+irSZIpM
aROh/y4PLGUH18L4EETgUo1smcyltOR3A8r0CK7Blip7gckj6bA5rwRIQ/XXR5Yv
+/0iJNWqgBS55V8b4pF3/QTSOyzz9sq7Aq8cTXcp0+SfB2v+06w5z1BOmUfIK3Ah
58lSblFB+Nmh48LZW99OfnY0Y65PFsZMbIdJPh5KO2e+kckZtm6BUMIasVi5NmbO
jGaKGCVQ1mOcXzMC/9O+AWeB83p03siJSPvXpUh2dWYkrZZ6Fs+XT6Ke0d6+FWrI
dSi8a5I77YXr6hs/WnQsZNQTl3zwgTpVylTqqsZ6tK+zk6y/OOfbnteEFoHfc4Xn
Mo8gTfZYpPeBTnFpex14HWY89iT7mKQf5J0IKkCmpEsEqSyq/ZnSKuD9XOK6I/Os
sNvTOiehisdjdmzhI8WuOHJ0LGkZJV+9hzCwyT5tZA9UHWpfAjDK78rVvQyi+U84
QEpukFVIi5JHzyrjJZHfTokYFcU4eztiAVeGuw6Zr8WgUsBho7mk6PcJPDlqzrnH
Pf0glcUPMkmo7CTuwdHMIuZNB6/2JRJOx7G+0kndHQBuw7gCCZwkM/1zXoX2sPKT
xEMKmlS3+p+LExOkoIVeBscQwwqvd8TWl/Ff7qQe2oLgj9lpEzGbWFB7DjxIaxe3
PeNWkQ0m6dd5yUvVgbih+EopQYlYMqf3X7FD5lVKH9YFf92CwI+eyL4SFS3ig7aY
LLfXw1GBmsIQuzyyj8wbNqObxgEWJKtlU5TIZ9a28b9+spsrHkx90tie31kgW8v0
uCYkjJREKWs4GoGboQQn9QHZH7TdH3GnnNCS+O/EhyT8ZK9WXu1I6ZGBmFE9z7H2
MvlosUuq3ve7Zkm3hJVPxcyuoHOt7RYbJ4MNwFLGJhj0kodDnR4CLhjOvODSNl5s
WvCpzbE+RSFSZ6dyD9ni11I0R42hnbv7lU0e0flA1wF3rBmHn//BBHVfH1O7ZF5p
1ke32W52vW6NF6R+63UcEf0EtgJMHKb4Sbr+Q7CdaBOTbU8Hc3SRMBAPa6cqJEmv
UjR02LfGjPJgZxFzEAjl/kJLtftzC5AewKy7WkzLz2bpIkGDzpr5NjLWOO9YT4q0
8I5ILo1d8hL9nkSpb5//SPXJDFCa0OMSAR5PPPyGJ6SPgm5FjNg2oBQn0OEylqyx
e1tS/ZHJsylYO9S70elBqwsVBWmZJm38incO4kK+oZO4XxxV8NGCxw9EX3LKo6Xh
kyCQu7Kh5qWVyPsHOV6A/qZ/jE3OsCPxN7WpEbx2l5ObaDIGt9jVZMsCbq3maACf
RRDhkMIiYOFaRLZ+A4ea72Wb4bUpnSFxooAPfSGkwdLo8NjvN67y7vrw/kE8CKUR
RP9+sx29FjDKOMrecJU44WVqu8E/Di1ioQ4GluJPS75SIqH79H1s4CWWvgxiNT3M
X104B73WgBicMEDXutCmJWImhZzRfNtoTeEg+i4aCrQqvvwodpWAUz0Mvb4Acetr
fkcAzYMQATLvqDGxX9/wLKcXG22eQ4yHOo7150dkpaD9ogCIovmWCUkqwFPQC4gq
h80dKtEJYsjoW17kDcYp+aaJWjeTp6AhNWB4bP7FsfndRBup8MhG07sDlfaw4dX6
cmXhyJNVWZ9Zu6MhBEBFbI9l6h6dvSe+KGLjP96TCHOmWtp3leiLieK9iyH+elQT
TrbqURl2Ib8ZySaoV6quUu3foWdF3/GKai9L1rcFH020APqh+c+dg9gGuJazhJlp
byn67tYJpQbDdz2/ibBpLHVGBrVzAppZDFDVHa3z5HbCwtG37ztyu/281ru5ErdK
NBHPyKRDP/vHT7tSTzKK5LvIwE13XCZTwTXO7OYPjCYya4hJrdUtWVmIy0dXYJ3t
MImT9m7vzuI3jVpGPZ2OFvGK3tzPJ6AdtgHKqXxkL0++MmZuPdF6hOC+ZwmU0PlS
oSOjvpflqonaC34c2Oy9okSp+gzh4ELOmQp0Jf9Zlo8Ak0sRohiDIyADwR7jVmEy
QFlSkxpg7DPNldwgL29wgWT1L1LHDOaMwts0c0GoTXRcL3w9jzlPIYzGFVVx/NI0
H4Obz9N1w2yuGqHHjT3lw/IMJMCVkymieu7P6/cDtg1ZyuV3Envw7bL+kmrDqZ0G
I0Tm79UAlNu1oYIzohqRW9paU8p4qnKenHHFY+wcQZNbHtV9KBKNC1CbgntZZRgh
Jo/xoRrF+MlxOf1e7ZzLgjvMdxTo7VYw5MGIMJ8akvGJft5Z+Krc2r2B44i0rdln
pFzBWZ1V1kzY2SsC2R1wARnqQIhP6uEVI39+EWXctwiYoncud6uShx6b+hN1XmuK
fB+aPRsKQtx0BQzbZwLlsdvy42PaeBxJSvSdgp2+u3Ubjol7OFsA+LmnOvnB6Y4I
ILjIWGlgpGTKV76ZGygdLg/rEb5D3BF5NFYAWGWiYuRXaiob7rYy+cMvJ9frXPVR
CuGK73o6SxML+iyqJLs78p3iq1+mQjEuJlbDusCAm5O2SzYKCKpxcWn6FRIHH+vS
rV4zSC1j0j9P3LT1Vp2iJSmTrx7WRgrCkrgRGoVQSnLLpiHpAGDUjIybMzkj6BK4
1vz1KOD58Vcwn9l6r+iuc4y9BJtb0RniV+nu2Vji6KrbbB8uW9eE59AMcgCnnrsZ
csWdwiONnWcwzIhyvnHE3mifOSkru5wlcXhSUnUaXxYwLxYO9Xo0nhbn7CcjD/Cu
Nn7idS/f6EH6yksEC4pNxc5bBjVKzuaMmhZX8oOE+/K5iJHloERrxHJRQ2hmy1iY
P3jddeiXdszAdDLVrLDWsNSodInC3hzwfoqkS+skz5k5IpktHY8e5qnGM9naPQnP
BqJfIiRu4cmch48WL3ztwUXNxsjFhbTSLu7CLTJTP0m5LNuf1jS15RtBSZoMVOu7
ZVL71c4ZdJrJdwOy5lKBYefAoe4pJq3Y0tTXON5RqF9HZBPIa33LOy+PziXFZkUx
MreqTfPGEA/Mj+VIZTo6RpC82nggfR4lj72iO4l/g5+qezCmINrlR+JG40k2Fe5a
rHeUTN91iVJRo+IqrgIdO4HkjtiDxl/TnLVkDQ3B7rZnFkppUrk+iSB0N9BUqbSd
ocKXQ4fnEKa/qLbUD64UUFfJakup9YB6c+jR/+6yKieMDzrARSW359gsoYX1DRtK
22RQQ+97JntMIgpnGaBUec4tHXjcdD2N5JYVpW2jchVNzavi16po3+zivpyRfI9K
kygaPLeQ7jLLzPuoP/xEnPR9UkHsbBrUKgtx1jysgwPqI2RXdmNnGI6dX/GTTMfj
gweJVAP1yURN9zVr5INI+Pbx7sMO2OjDz+8FCWtS8k8g+VcYQ5V017KYzC4KVbiO
3GSMQafkLdJ/TIhdJh+hIHjprKdcQawNtI81hXDxh/I87bHBcWDKl3Gkfn1bRAd5
JJ1mnrgAKo5xtoT2AdGxS7SeqYDhGcHiDKN2Hgz/fd/eVvvSil/mHNqCX/js+OxF
p4h0JQTOvLIu8t/zWojfA1FcySCufRx7vZfjVqEyEL0WcjvpSII9ZR7cPj+PwgBX
gDfTdcqVcDto5JaOrouabe00fYq1T4yKRE7A2qg3f27FFDyjJO5g9wVAxV0h6zZ0
iWPboEquUGWCi6VKsmtv0IEm/TzRSbLdGofs29trFdN0TXopB+5UMlrgmm+bj1QL
q9JS0IGw7IB1v2Spupaa0gCmtdbjrGyPtgoW6QIkhbOguy1auhYwjOCYdEtVemcW
4Hf+Laf42xT2Zk8gTtaTFA1K/dtUTg2Kxyzv4hLSHlMPLYezu6BSyCMsgl22W6Is
9eNA7a5OL7ER9vtpmdzVfTgXKYN2bjHcTRErC50dNWCTUVHhiFcUcFycPanyu9UF
RCtEFMeWVX2W1fEbt+R5OPnKIWxYzLvs1Ssefd0SYm8T1fXLekcrwnnF64XTmqDd
NMqAPi8NaguQGuLeeC9SAzpjdonu8mBw68lzullBp8K6N4OfzhoL4tgEFzWqYer3
eNMAlwjQZJqvidIB++zv8v8vQeS/mziy/M1ji54hf7ZiVHSPppUd8pye16CyZOr7
uzNgKB0gBePUM7EpD54iQ7LM+d1pQ9IgD1l+mZzVwDy0/AmomHJc8pRsk0KS024g
NeOtl0IPPtDUN5sM1sz+tWWmFGAeDTWuq77flTUAmM6PhRgOqIcE86o0JgZeZvco
kc2UkADHBObMZbf8KfcmpR8wggUBoSOMD6lmnITUmApJd58TEfccM9evpMLE+bU+
gZXPx+GYh8aONuz08cBt5mWd3FYfTKXrqOYU/mcGeVd+OoYQyCPpX6Up/mKvpFE9
N326j6V8vSE1HQrDF8W4kMcgBwWNz2Cosa7hgHxx6OOVMApirUUMGzlNR7CuURK2
NiXcHadufiBA5PtkZmcRyDxOEMZvV9dXWweniBCg6NrZj6qAQrhCsl9g68H6Uh8T
qZjCNhT598scCgoNDj0/1C2kV9+sGyLfuIJH6W4a5Ac8fBAZijp7zjwdwXHiznjm
lGVKbPWacmJOrm1gtCDigvMoc5+n1fsQLoF0rclx5FoEJQUqD1U+5lxmNUlftugh
ZkEnSuPMmtqUjROBzdZgvQac5e0qdYqW7KDVkrkHXujgky8Yqc9KXmxrJLt1ElGH
u5FGTNpV49x0cdJIYwOn4s5FfE0lWfEtuQojf6lPd66YlwOBfZs2rmgRBOR6POf5
ojeLlTCXtx8nIp8M5PYSZK4ajItXrNwDY8wbGeRJhs4YpBlZ9OiJZcKe+Rs1YVJ5
6jyyigcdLtlPN+z5K+KBzfXhdfh/18IEkFswPcLWoNs0d6bW7WrhhzA2v/gAc82M
G6qP8NgUDVUsmofG6matcifC5YtVEjnOdc4N0QM9Y9Qe0qNjqo0zMWhso6HXMJwj
TaOeYMA1MeGZlxzJDTTrWTdU0+K2CT8K7Np4d7+9GFHEDlmUq4K1ux3dAo6XjoHE
GFFYOY8KStwBOevHU4yvqn7QvwPFLTFI+F0scmNWN1rgwVzKVYf8t/xnYXnDaJZ1
KTB24YLNCnYYwQ2hY99sQP0VYB+EhfGg8fono3yqR8n5XCMXdfAqhPvCCPDw+nx8
8iN/DccA50ruHykqIIQlvKIsxoAn9bQEknHlF4+2K6TJmOYWQIfpFOHUck9GYbOE
k52Z3xDfv0ralWtp71Zy2AfNBjSf1MwGudfdOITWTc/cDMiQf0/sVad+JYoPBHEv
t7WeZJMzJAcqmtz5SRVbKSEg5wGy7kwPq15hj/3BXmGK4zerXZxhPuFHWHfZUyVV
4jgOIkmQxyhpDnMpYBpGShl+vqenffs1xf++Xkp+vOcaQappyAOSFnd/8VrIwqjO
pYZuN7CPinjs0MFpQgP7TCwdedgbXOKbgGdOCBpeuJbyr1FtFsKbVueqkLkvPpHM
YMyF87BU8IUW1UR/F3cPgs0rH3TwXmIispU43CypufKOd04nlbgGmoNMWQBbcscy
IkgT6vD6ru6x7Tkjx2f1vWik6gpwmDXnaevW2iSo8M23DLorZFjOGZVVEAqcPC6l
dFgxmJyIWIMH5P2GdY8S2C2hdj6DxG/cbL4mIoXKkpFmZa31omtmmvfFEu96lchI
GZkTjmoE6MEwYBUk7l4TGG2aHoFYJuWeagPkL9elZveZV2tZwSz+15G4rCbrdFl4
1VD06Haj6IQ8rJwWknGlVItxtLA1yMH3QsXrhxrF/+Q4mL7WzE6J6W8RHjTTsKHd
oGDZPgRiQp8g3YW6X8fJnNjMgj5Az8mV2/zljaKIL8yLx+ywPngAWgEvGjd2SFx1
6RndoQUjrkmFyhIcoiR1aJb+W85Hgsu3my90qTAdkJG8sjRarLeim3ijvd/ftgbW
RbTehCokZDgxWXUVNKBXeLDda5WDDb4mhnRD4u0jBd0EwJUNbQRA3GDqzcggCpbd
Woc0lXzl5B0lI6FGcpGjG4zOcuyDCqOpQM/oTAzMAj3IU+mgILJkEHlNExygY2Hs
kZUEFH/9nsSuh6d9Y3PY4Mpivykt4ztzqp15q/CssMttaTvC/07qIS6p1+hlHMRc
MZSgjfJz0Nw15xboWg1QkTB/2jl83I9O+lnGDrv+1pKxyoo/U7VOd3Yr48Td3KFo
cVnzxjiQ7bEJ+vxG1xYtLDVKHhlRzmosJD0hDQ3Kh8OdR72YSWdvffuy2noQyxKY
ksxR5S/1okUe0NHEiN/4vM0bz7diq6ule2c6//a9sSr3ZSyvCkfe0/RTZ16hcmoM
Rrm+F6ua+Es+uiYEYtJLIift5sdzn2b0zZWO+iltKoBvOiQngbnwAegYvVB2W7GL
Ti7sUKdYJusBVtm8EvE085qwhbWRQmd1A2ZGHgeq3/dLwQn/xx+cZCMnlFZS8azR
cLnmEJWDUZ3w8569GBp1NLt7mi9r8zPNi296MNDPaGWSW0fzL4NmaEIo3RdD09ed
MZ2/oL8vHFbwjSQa0sQu/OKVAavVzJM7RKFiar8o9fyKRdd1tQ3quU9b+2NjHL0s
TU+CyYUlDRGJJ4P9xpqJb4q3il3ip9oFV8saH16qAzehh/2IizgauqJvitdhFQNt
jvnzQXE/AfiMt2cHRXuPj8wAPSYkKI+FiW1vlOxPR4emHXEz2/7s6jj/ib/bceST
pkleh3wdxE+zGnaCfud266oFBbIssll8HP7VkIDTP+A7phuoU4pgnPCYMS2KHa6p
oUillgdADIP3YrAwAXAcml94EUegz5f5s1RsBEZ3HmZWFShAnW7iC+pIryH5hoZd
aVVBPt5G/mNNOC+QFXYGPf7Jae58IsSoaTjFQbCdfw+KeVy/Rd7GZFVH5h9wye5e
1DtKUMJIBKazHTezNIu+7yWpXkZ7zF3ewak90XUuEEGxtcD/kQwHhQtQul128zjg
qPKS5TLD/BqEnRS2Ms+kvS7D5LMhilqTR3vauVJSz1LSgmKoP3RZZNswZLfzLXfW
1Yg9K8kAQYUaTg0YBMHhDLfjrI/X2QPLbrCJEzFi9ySJ+wP+eJHyu9Z35BgSx+kF
fGi0LIJ14VinB65Nnp2SljR97TDW32tg0vGb59cGV5LE/or6x1/7gGLCi6mnBEM3
BsHdX+4xkqzqTn+HV7bZJxIfqXK5lByI7V908/IXuems8vQIR0ORx0lTo5uz3/fU
sILDqbbnUD7CbKs5v24hS9gurVDGKKKfjeYMs8srrHYG7pO1olrLZUKVY+Y0WdKv
h3XmraLv2bVFGgu9yaVAf96c2w7NVF7u+dL5sLnLQ6/h7tsLkbKwjTAA+W3yKiln
+Hlr5HxibDlYyWiF1RQbcHh2+09f8SZt5qse0yf6Rz3TYy9DSw6R62/RlGV7k86Q
e5OYdEvGwScTftTvN7/xUsc9FH/7dR2Urcq+7bJp5c3L3/HNIGcbCdvLYLBavmHe
ZG2OSX4fgvrAX2uN7FnvXDClirjnKoPhm6TyCSGBXjkUICWqRuAmHs7xsS5pz9a1
9LypfeP8U5IK2JiMhOdXujz/B/22WM5cXp7wnpDL0YP5ps3bQLTbk/vIoz4qJd52
wOn3OzQUIa/512pQDj9FVKyJxonTlO8qP1hC3a2pM/k0wdi++HFmUQeWgWSSFCan
uRaCMvv+ukVjOBndau5ban66uNaOCwSxg9QS6i69AX3V+dG66Lj6It4opBogAeuf
TiMQW5DyOCnnWYXrSVsIEy7775y4+byl7ZIj9W0pOZJ+B3K8gxVHW2vGZULnVsK6
pxsyqdseTQQYffW6qLG0TIsey/axpUR9TOi+pbKrqV0n1fJa2zMlFbGMLsSTPGOu
k1ZWQiCGbbBhZFoksaaJQtVEOtx+pILC43qnbO5bKcj7S1t3pSJTS48oAYr8Q0Bx
G5JaddYPy/UyUE1V/KSLiewGmWFtzbv3TnySIXwin2BhpojmXOXTLRDJsbJ/rWbM
cQMr8RKosPTD9/2YwB0KeQyPqTDof3ya+q+g7iFMNrS9U3u8LAae7MfcxtG/0u3Y
itkveVOzgisoe/Kb2EXzV4XHEyKWCfNruMuLaaEV2+8XI/jERXhmzdqdhSrIANQ3
sQLGL9uivGTMUV0mnhxdFm12dL4yz2AZ2jEbVGeX1mlBY2r603rnRv+VyHjCfkJz
aISB8t5tc8EdKQmhj8fQK6IZCHvXfnkVBm/yb8QXIwAB4ctJ/r96oJnsV+0I7ozE
CbUH+LSwMrx+9Kp5KEzwSqqzMz8EXk+NsrxY2e+5fLTjvsiW7Q5aKPHo1P6iESbF
JkAD7/tDoEt3EpmTHy/g+HsYGp9tAb/yDS1zQGF4LOpTCnHzEUiSMV5Y4fCedWNw
ZxqsocA+HcmjT05/Qrsi41QO0y5LFIqmhrTJt0RR6mXPkD11oqgQraw+TYdP6sqC
SIPgUd9Q0KwLQSCjdMrHDywHWvF+w++aD6r4fH0c/xVFPmtzQqYHi0XjUi9q2VJe
uL3+MZoVQ8fgIh8jfXWNhNFnXEESdUE7ydNKJX80WzVzybnHVTisTkkn6VbFjuvy
zcHuSXpXiUQAxBbpMpxJivJLptiw7v1Lny/KcuJo0Xa4pk8HlKSPi02S6jKCh1St
d4RmG9ODdD0iVIdvqBUrvaeBauGnfXkjj10FM+LLYphNyhFWbaxhMNuCbOD6T6t8
yEtozTksrE2yhr6yPQ121UyYXA41TjTsHka2iASAKquUQtxjqffq97u8HBKhTcBb
8Mmk3hQOZuhXKxiMq/Sg19EyeQBAnMLTpxXkicDZo5yKMv/RJDD6S4pcCtgatxBv
/hng4gNH1OPX+JMxWZNQEj9VV2xZ3B6gnNSEUykFh5VShaxKRc9p4SGuMuNREDkj
YSx1E6C/5uKgPsX+1yjUNIR3R5wWZQVoRubt7G45FRpGQ3NNEmwfEuO1itNUNz3R
URThFcEpyV5o6IVKRBxyEhE90MuctC9UUOt2g7VAq5JuUTHR5selB1ftkAoRwT/g
KwbP46X57yudKW8ZXSMaRwRTBIHNMmZuX0bdLCqoZGno9Jk/9uIYmWS6LAJPX9GP
qeeWZ3cj9doQ20ISXexES6hhE3M7gnzlVlsXIidqYV1SspZerKMjA1j7OrABsmOo
ASr7R9SPCCDTDAZFAalNJ4+wElLuytqSbM3N8i4xSPJomuIS1lF6VTc+LbA0nhKW
1rC6wr/m2JGx0WcpVW9iKYHxFvVCp9ulG2sDAJGncvoASWxA1/Q1pL9+tu93JytB
I99rCND0d1E5FXjvl2IE7/gNU6SL8O/Er7Wed23hDVYsIknHjQzW28N/F0xKGjY1
q+URS/ZIklXTlbDrtK3Zy/Ol2jwBqpcwKNjTOa8d9EE7+sIHbecQxGOnRo7x4ayX
t6P3ZomaiWmtNfYjTD2h4/7TUlf9fQvuQzem/maVl3nTpxz/IwFuJ7+iVrFzB0Nh
dTQooK0x7tyCOgqiFbTIi2Sk6GLXvbix4yaeIpSxdfhR5HrnMVUv8YAQVMLgFE1c
9NUc45GZeNCjRVJf7fN5ZrQr85ku0HcbE656LgT2CeKGVviZgYW6IBofn3r9oDHA
XNZHLhZIj/yhAAA6R8shCPKKtf79n8kuxVQ5POjvKgdYszUEMt9MmZuG3KI4Mu0h
tJXfHbo1a6LYBVhXJqqlbgB5miZ+0HjltD5OqpEt0BQJ8cs2L+T2+8MKgZDfuKY4
X9Nji53SGH3AwFknrIex0a3qTJEScf9l0GZEbktateFhKF7g5wKPCQa/K9FPQBkU
ywQ0H6YDOvxXNVqj/9IknUxF5dbtU5FAyWBWXB7yyutED428xfotV9zwHQs978ML
51BI6jetSMZbaNkSqb5hwMd/aG7fIJL3///6Jpf1LKKBuZxumbGy7smxgRTSPxfo
kLE495POUsLUnqX66/tnK/S0yOOCyMSeBTLotDq1f17kmRloqVDDCrA/q1SSRy12
z5JXZ5MPpS/37RZMYJmxQMNUaIoFWyzVBbinA5rC7wJIgkUcnpaaJlGILEgabNuH
Wggl6lTGI14pYNX+O0iEi4Qwalc9xr8e1BlM/w3r/fmIwCr83ZE9tkeM6tQxtv+P
R/NkKTt1jZcuSbijvkR6WyW5gPpTMhqGfbfMvkUi5Bp9YaFczhOQq9w7rXJKFD/S
ewiV0F32gK97Sv6UORFNHSO1lJmg8yTckWRwXxIGEy8TNHwL2WU03WE68jrJg559
dyyJz2nBfQlaCIcS4T4ekDCEBM071HeeLCzn4N5asq87JMAXt6pYFj2cFe8A5Ur8
smumeakidWgvt9bV2UtKyPVPGIjSrE1AivfC/l74yFa9QzOUufMFpYThXy+atyHo
seULpQ5oJmiX5dErHG+XMEGbF4Yv7BkvMhXRW7co7Qxok7Ra1AOx4ucQ39/HkrOO
gKU3VFn+n3rPcfLIZKBGdCo0e9l8HxNs8qvOGwxAlSJQr6Pxm2pLBGOzCJrzKCHF
fcTeOw4kdREO3Pef5BjUrVZ7cw6ndgd0T1DrXlYA28vYIBUddUffPuA9cTvMT3le
6Y7g6JIjnSj/F/rg9Y2PVfys+zmj325RA6ivW8vZHkyi9jiAE5YIiKFPyWjJM/hb
PY3KNNG2HoQ8assdrJtXrtTUSdx1jHqBxQZARtNlZlUlyr1WKRhbw/UK9JfzKgJw
8ZK21jaIKzusHwEk4Qb9qECkWmP8OgPoTesTR01gzhFaglNbdROmd/OEjkqVfE+G
vwCktTysoK3jEfC0by9lg52Fy4WBnJoGGczSOQayw5Z4hNFlG1urLesqBJ0z1X6l
g+aE6/SFqq2YX9O20AN3XjwTJrzV5EgVDcc3ScKH13j9BkLzAUByW9rwi1QfjsQk
VeJM6w3KSehJZZt1H2QGzGY7dln4lYfuszW9oUA38XTzm0fYrx2Z/QGkiwHh+uyE
wbn9/jbewZhKfD6OVSVl214A9in0Yc6docjAV9vjbMFIUy8ZZq9QODBcWzwGOneL
/G23/rJLpnHaQzYzuf2m45ym7//+MsPl3BV4qkaf9FJDZcIJo4AwPRI63y9JdFkQ
LtMVZpl8909pi9elE8PevfJAhGEygyZWD3AD/a6qqNcxfLc+adyBtSPk2xRl8CAk
znUoeSH0rO+DjMVHwGR2TC/t+rftRiZxBCIpkoL+q8UlXhXI7VZ62hGqZQfzXUOZ
+JErvehO2cr72skJbJdYMPwcnh1L20jan3p81o0jzwI4+zbFoYdQk1paBPo+uZ2S
9bHjKinDK/0cEkRVS7Scj2T7RVi9zQ9YdKSctvvSCfzEvLQwIS3oAA/bHpSK4br8
grIZJuegK0pniXiR08/GiSvrc/eqqLfU74hDoJ6KFnMJAkggBJZR+0JAafnXTV/E
g0/ZrxpjO3TteetIIEhaL/nT7BsTi00gvZfSDivkNqGN8pl188F/lPS3GLwOKrko
Au6pP+mb4HMchq8+ItJVUYlR3Ni29wD6Qjr1zoLTlhSxEPPauWuCPNPrGasVK0OA
L1y96EQWo3JvLcDgDUrBc/nshOiK3CBWZZlz3w5JYGCXxGQG7sa1b9woJ7z/I5P4
v1YX032XKAacdpvtUn0j8jDZEiktAciZrqU7/g6ZTQEEXm5pR2tshYLB+E1+hVGp
su3mIZsrYQpLVoNKlVuoD6k3w4Siu5QEaPMYt0zLwVCXP2mvRCSRPMRagZHMqdKd
7DizyLVtuc/hEEi+EWz3sicMSx87kDMb08TfhPHsTxEvdRGt7EmmoqblvXlM/oZx
XpZuSJ+xxg9D+nKVRiv/x6/Bmyd3OIlkjG2/HbkbeJ5QpobZua9V1jssqz+SXbVN
HYfMiyBZD05Xb4HzL05/8/aEeCAI1Ie6T9JjggAcefGqRoeUYictw6gXRmX8g387
fBKebK9W3TcnA1r128Al03kITecOgW35Z72jgs5jUD3HHsr6NWQgyFqqt1iaebuT
1RUQFMHd2a+4hbmr3queJdWEuVkWNlrbEO2uiu83EacTf0dyswmbghBIwav7YgCd
eslSyU8n4uInTfWa6TnXBKnn2Rm/TnVdlASjkH9PgdS7Bg+axmP0EeVlYuAe7FSm
jbIL7cEiPeqXW/wT20LqVTSV4i5cp5Xq1h8z5QDemoXA9M+cioEGcwzx49+rGYBU
mHdB6O1VJ9lN6WY8HKxmAmyF+3DdWQQEu1YwhSxpA4Ml+b6aIf37ztKZWI7zmghp
GP8VlsVU9ACcg1WYqrXh817ZIUaNSKNkVvRCx4fINGpyoSZ8nTcOViK9ApWEAS2q
UPHDG4t5OqBQ+IQw38hOb8YsPjO6vs/JvMWVmW/62bg8nhzDK6Cvdw4pv/nhfo0h
qCNYhp1dRe+pTVMq/dffE90Z65hRtFvdoZQ32sj/8IeikqsGg0q4BYLaia1yRq0R
Q/8FsAo/KBepeZyeMDfFpRopBom7ZJZMJ+Lfrp6YA7l+TrR+S2IT9/Rjb/h8FLmX
TfQrenqv5O9k/1N23r/JMMUbIlW3ugQoHjuMiXDY2ter1ix3O42Ne2DRev7K0zTq
6cPoIy3JeiGU7wHWNai8nK3dqZzvEu0V2ZuvcAWSIKdLKsCWLbILYQ6fPXhtkmXv
W0QKvAZgOQsZSF3o/g09mAX5zW2jEGjwrZmEVmNFt/ExKum39pYn6fuH4BSk+nbe
3C9bOXZASG2M8YAcs1DjIZ5Gs8FAQIvstzFy6jrPdmzIuvYG67hda6/VJkrYmCXc
T2GYWRmemaqAf5OpKwIOSq+Ow84Wrri3RWlDCJliNNQzUVZ+DhFsJlHqwPVfZ23F
TdY6707hwNQSOw2HBl/L5dlmH/UOWozV0ttg6k8y0sW8Vl2l2D2IFAbr0Uuxo1ni
uJewAGhsQPuVTKvIEcmtJl4/54/a5evGarCnZa8zPwod3EnDbkRp1XkRFN3QFGhe
FH/ei8hX/X/I/LQ9xv7mm712IGbGzsP6UX2unvZK1XdciZFzDeRP5T1Wx000fQfz
cgXWTt5P3Ysfz5T+uLRcqZDhPzwQyinJybFkVvesSG924y3z9ByUlYC1ih5JZkS3
3VVBYY3BlSx3qrUduwuFTzyJ5dQ/SQwep2QGqR+4YowS8bC0oJUiCFE9wg4FH1PS
6gv9T9tiaIpkiarQVele5QRAndwXH8PSuxUbOHvnOfEUSGG3EAEtd6wywLcO9IL1
xQ0Xn9AuSHh485B0GT1OkOr/FeFplMcTJyEvD1kIU+j9HTo8zAAbt24RNGO1iINy
vryjGbQlBNNjj3pFhhRnA+q9mzR76IGlC0b3l95tFji0iOtoYXTY85E1z3V1+Q1w
0P4pQ6AEbUTu2/EHo10ynD1HoG6rISnmGZCldTSqpBBZfYHgbei2nyTJhWjuKJkc
SW6W5qPMiJ6+pjFSAmWNWYePAuoRMbAQZ2ifhj598EsZDYI/U7bdekRjohslauKT
Lo4oxA1v+WAmwP3cQKadVUs8vNN9GNDPHyOae6qHfCdk/HFfGAcvhpy14+ykQdAX
kpr4vdbjfvbMpbDhsQPnjCp4LYwP7/CY2KMamReQiubCol/vkRS4Q+r6fiHqupuN
9S2oLYOH8yTYegnbAZ6yOLbIkKs9lNZCBMLv9ijkhXdGHe3u/ewkCA85djwuMbpD
fQiN4OuNiYJy7Pjx5DiTmlYWVSymDfjB1t1jQdERwiHZuELHcznPNYtb0xRygPVS
ehytkPLwu5h+qmi/LoSnr0skfC2m8G4dx3hr2E8TJJq8QNyhrOC8DVTYc+jhzgTH
5o17Kjfwh7P4AL2mXutNPgQ47GU+6Wh9mrlDxPRK1w9cjYVJeTnhBdQcfanmbMHa
q0C35+Prpxtf7ACV4ELdbPREbOa4HKXCIGodp/ZIRagdaQFmX2Xsn5ZJ4rDy4oBV
KZGBQyC1HxVgTXZxdpet4H/PztT+sEESC2FSjQn3pODUfmb50EOOYU3kWx+YsuOW
AaNk3DsJtnJrB0VSoem86kLvUUWpOBisNtHlN3tpomwLXM/4iXeyf6tf3R1ZPOyV
8sHOeg854bliSFkDuE1TX41dJMsil+/rECUcqnp82bZhs5O3ADlKAKl2WfOKWK5/
peUm1/t8JB3/Hn9FyxoW/ogHeEzAuZHwwqLyohiD76l1BVEExo8yMvXJ8OC/exWF
JQY0QjhaXFQutt++U2h1H9h9MHWVEhSKOMa6jHgtxxAYXPpUpBtcwPa3PtDwbN/t
eYmtADEFnmH8gBNzdZrd/er/fLab8uq1lpdJxNufijb7hBR0ekWau0NKQBnvbEPs
+k/G7Ih/JP8XC/tfoGrCs9V5SWEEU+SFQwRW3gBCgn7oNYIqwNieTOEjh+PRtDN2
qC93dJmuo22HkqCWbtp+7Wbx/o6sgpD0R5KQOlEePe8yx3O91XIAuJchd/FL3Mt0
kzOZzXTa35IB8iVLdVwUiTNyj1441hQ/RwmeQnMVKWVYyrifMNzZEwkdD7ikITVC
we5cBDa8xuP/V6KvYthiRrXdTaZDzotNFnfjaoVTjwPAd99rOSp0GPyY9i/5mG4p
6nWXVgNqDpYMAq2BFMLWKuupF2mxHcBT6nSZDjCUWhyf37zDEHnuokmULoSE7rbk
g+OXY4Mgu3Eq2UezeYw/tSrW/aR3l8br666qKwJ94AsK37jSoFM58kSeczSNrRFZ
XbEwHp4TYs0ECsW5UwdgPcuim3YnMW79bs2np/m5iLBxZZCECgq3es8nlH7n8OBS
/j1IE3/IJPZDoj7l57wwbCOozW1HqnbluWyEPoxGXahkjRIxq4A3qoURro7MM3zB
IH10vJ/VZrFUmdZzwUDi3jzaNb8CTq+Nia4F1hHFdVmz32I/XIhaN6/9ts0uXYq0
wMdiZzYyDnO/QjWDiaYDLbR16bky5JiLDX43ThiYrd6c0RFk9Ki5m+M/+woBkGT+
3hUOyh65xNqkrMmJWPdEHiZa7ksX5OrSwm+pe9zWZsGLEoAhLTSzGi2kRH/qr8qQ
41+BOwuFC13jV7fAeoAZwj78tzq0iUfkvLthwhpu28zJDskVC/RH6WScC32tzSMe
zgrXicoTzXL4rfPfZNQ624Jko6l54x/5ydQ/ZV89nSG1G/Faf9LbVtZjHS5KtkyO
wocbtFSbC/rGIpQvNqkXObUg+eWyWUGKToMODsETrz37w7813x4BD1qVIhYPVx3J
8TVqOzp98GWEa0nGSHNxC0YYWSOscWtryuVadvFN8YeqeWSs14pJ6E06e9WhINkS
6PFW6HWKde+l8zs72JKQDt0KUXoo+PoxJgnMomBs1G3oXbaH2rBxib3ZeH/ZB9r9
99/6ln2cFOYGqLvcWi9RxF99l7NH0WcyaTtOQIP3nereYamtEBvtIkQT+GdDXDO5
TIchg4xG9Ohs93Y8ej8LIkmIDrZ679Eo/7esqIR+X8fU121sdh80/W1s8HvqodEr
YPLdvcAPUCoUTku2m31sDKfzOcJspqh2AKT/TxsjNiD7NJ0+qTJ0CzBK+CadDgtt
1YYJ9B92zTio5B2aBcCWLZLd664cVSDlRRBgnnKgzHy3cj0pgWu2TYSbOk9LKLFs
BJdrZrgJKAoJjpxH6Ek5f9QAZSTnzKctrq6JF9Ys54VknN6octAjR5A4qeH2kAaf
eQI25fsKpSH0xAb57dcoC2dS1wXscaqhAYp7GtCviYccl/Rz09qbQKzsg3Vqm/05
IZ0jTM9P94BBK2ieCQjq4K+umEkB0b6GZoTwvM5R3DbsakqD8R+g/p/QWblMBxq1
VDCnUhtOUzTAV54JLCMU9sRsTxHBdtCuzEQ/LfQZqcV8M61D0h+U5O7TKDQTLTST
etPRkhJ1VbokKR6jvn6DSC0rBhGLCVJUF651mfeGxD9kpxvSMuhQlUE/RrUoQ9fI
yRbudRxRjDDYDN8N7XgjFgK/nmAb7j9UVK2X39z4IyrThpTyARSf6BRrX6Q28t56
UnPk4hwimqxY5iIW2HGBZLahH0j0brzGcE6o5mwBZM0Konf1JPsNcyVbV0hd0F/A
K3gKH5++wK3g8U3NgOZ0y2qzuvYbULAZN/5yL3wqGe9KNpC06yYoOAhdmoipmvCJ
6s3sP3k2ih00TTx1XaZFpCj1usvqGIyAeMqODME0omS6oLMotNDzA2EtoJwQ1lg8
xMl6AMhDPY+SdFYbjNkkR4ajaGnEnADSziGfQpWOSqMGrAfk4Pn9eyyaVAhV94zL
VX9BIRLYxjUyqYs/2JnhrT9DAp/zOZn/dnXb/FfMC9/6DH/j1CMMYDKg1JVGqEqR
KTnYLm+DyIsNbO5zk5FivJqmLyx4L8/9no/p7qEv6F92JsvVlvWZt/d1J4g5xCa+
iIsnQySOw39H0iLZYmymBvKXLfwPVJdZqbtv42JoWC2CmbvH3uW87DQVuS9XZiVL
zQTH+s55P6VBVPdWTjtNMoUTXkKBeIOY0W5r3CBtu1utkPMHFCwvDEYM3iHtfE+0
NTGZIKjhc79SZhGUhLllnxsWPq6l/6QR63XPnT/0+UbnakdQ0oqotMLrzwImDcTI
7HSXX86533XNp//VjzX1sr4O1dKRh3fU83Z0+g8lmSDl14BomHv5cBtoLULiIdpA
9Xd5OFwZqqsCGGl82pwvQRl0p7+aNelS7fsceTFWMmpXwNjlPXI/nuqs3zDN8dxc
gcU7KbYV8ELDvs7tX1K/Q+FdWfvo/NVX84YqKOJuLFqTjiKoxH8/L/LKBFokuhpw
6g4D7d1fCip3YDdAx+zahxmWpPV3MI/BlpwriyEhjvLNu2a444Ub+rLuTMp1LHwP
QwAw1cLxX3NDtyAkifJ5PKY9tHE+X115vfmO7yUAoOQTjHkhxXyfx25GhoUIKxhX
r6L5DzE6XDS1yh3+fHTj81KQYT2L7QYwiJC79Y3l7kJzSEap5aUDg/ASMtpENboF
6glgkGyUFWBXYaDz+pZry9S8Jj/Svsk7bBhNnW/k2ik5puEU7FSe9OB3d87IabDu
Hcmp+Eh/foW2YckBe8BL42jr0qZ+XH/7gleArGLMSEKRYwxpmkBbCsLUIxCs9ykA
B+0v3eLm6kfeyE0gTfI2DMihpPoMtmIg1O8R0QHVkgMQG85PSNMrtSaPUOq08Ni8
81FDn6CPItjqaVkyaAZxdOzRrQb58cJ+YnzOJqW9d6PTlD4dj1MnNG2vcJ08dINg
zV1qyMaF1m86JCxIrYTGbJiyrgX8TMM4u4oT/4exxdg+cnH8HOmNjx+DuQTi3CGR
+5ETZBbXhb8kX/VrrB3lJfDpf1ma4J/V9ECcHZPE/zGrcmCA0wbwzqs+tHybKnOG
ESbyEY3nrm0e/afmIvw46P05zFwg8zZAyLshxhMaR/tg3kTu4ItCm60341zQfVB9
z3yBAda3HUPKK+DO1jSgxHiye79Bn0uUb7gQFGmuoBxK715YNTiNK0NSgqgbN7Sf
Sz08fifOlm9/uPIdc7LsbBrZ4RKU7D3ynyBc8RMzgh8VcTcKeggQS7DOViwtXvzW
LsxuP4CBMwGah99oeu6pLJ6AxgfAcAhFlqX5cqoaHTzRBfRk8WQ71kDwfpeYX6kI
yjDDCZrVDe2PLR0lhP6kuZylzma0hz32Qzz7yNuXJS+7WC3nnwMEU46ykqlEehoK
RUl1USCkbqLDBsV3me+oN1axybkt+I4CGHx9PACkjBB+6llEMSwIAI5crKAleuTH
+UALUajzizh//LZ4foOsbmG+NozGZEUCROU6KLc04MoPYyekIjA8LtsGv/oT8z/M
Ry8WFcG7t+91u7MFtVhkJ+272e+/Jo8fR8O7WeAZh70V23Qyheoz54hnpRif0pK2
0rrQM4ZItl/jD1C3295navITKItcUtIh30nkzT7xH3V6tKx3tCnMKJKakgXD6LlS
LecwE8x7R4dm8/XI6eNnfHYIfml4LwgxQW5HEVngyKg/5YzxF/eHHImjfiatW+xl
QtvOAlRtD/X6Aw3t12hiRnkelR/u7n77+FDdF16umvUYfntrjO/+GDgtTrqoVlaV
2mAbXW7aZNgVzLlgwoQ4aqhfTxPzv44xzpsALmj5l8mf6s0ePPJgmlV3KnpH/ehH
fyl+XFVMXWmQAMhc74E9GRD+pIwY/aS3yMcvgKFoRM4ofsYDgODu+pPDUXguPX8i
r8ynHez3eGW/VrKxKDopNoWlj3XlTwrLoh9BptvX4dBdL+Ke5GTeqYPmYchNklJF
Ajr3qkdIoXqjyCrvWenZAa6/fsiWLa56VzjQaSTPUDLTvENA7tM2UIUWnWzhHVB0
hkScD2U26W4veE4fRdPRrvHo2H8IP9tk4Sl5/K1XUI471Gst2axixZUADwxFobUV
ZiXVeurVoALZ8m+mghTUMtG383+D0dU0MOkvG5tfo7QRJVgWRbqRUbr/0kUHjogz
abiihiJdopiz/uomLxo6P0TIYM2IfRWXaOtyG2rIZpU/MGu0ua41sbBVbLZBmZFA
tZmqt4JeQW8/VCS+Wlm7SOFy0MBNeaLFDVXU0EdoIV6JFmiVePklwRi3dpSZfIlA
4nvCfDBNfYhZoNGvpmSLapdi95d/P9qXhZfFbYYILoXfJm2RKRoDQR2ZpVL/F54n
kesUiprU30HzWjxzMmWYY2v6esu8eOOZ8RB+3JXKPZO/hl42bf0oF1uMe86rRtBd
s/Sqhv4kZHcAzKuHcHpSAsVifniw6WfVeGP/yT26j+G2r/02CFHh5EyGacDbjJp9
M9YIcPNv9aQyHbh5paVvHOCXBSNPsHHquuOXYiEyebI3f6vqtzDhaR6tZK1hd+km
8rIPrmgtRDaBPzMpTpiHbJxKHvX51jtECBUaCMSpAb83WCRdwc+PDa8UYlWkib9i
cHLuJjWWsSIMmqzXje6y9VXGYoYWz3MgFP+GSYLdtfwQlUcVOYKzgTeWKqVRT59s
S+RAco98hUcBG2NjzSPuVEGkD4EKjhPybn+2jYxKw1EHAZ7oek6O3Dg6dorIM1Z5
YLYJJ5qfWQwtQPgmsiUR1yZVxREdHn9MkWCNQ9x+MVgmQee5fp7XvV/L1SuxhJ7m
ZG9vTJO5V5ictS4zeDax7vTdCiKqbIjXq6ChnNu3QvB+Cur87QZ/RV9+HxfkNdYf
wFHwfiDjLaPjEomrrcDiYnkZg8y6WwwSmFLPjUfMGtvLDX3T/HUg433qAV16U5lc
GHKV0mMQ+eoLdVEsJX79Uh63MBo8SyEjuHh+9yXg/conAPFOs7Y3SWrAQjsFyTvC
xDsOfhrrShO9nDzCW0HjhzXOF9fc0RiqwW82Rq28SaVCUhE31NgwqzQ1JAWVyGOx
NerOjOMkSvWkc3Qige309Te6yDXL2QymLThBBInGkyC+4fhBVWhcINBEJubQZWkz
TPZxQOcZX12yPXd+deKAz7oRwQ4IGsLGvvoFTfaUO+r4IBgnihuXgiXKcQwEXbZL
p9pwxC/+fqSEzs+yXujHL5iE6hmHvtHXY8eRjHIEU3GCcg0lG8yD4siQO1mIYy80
+Ou8c2NsAJ5idK6eqdGtr833JWI0ktM7ieGKmFkeqZsOUNIxKrM/+6z0h7CLPCKH
PeLKJkGgrV3y6RGhsTB7Vhx5mfyY1mDbCx1sbHPffaidowk+nn61RxWO763oM1Fi
G5qfl+2IWf0ZcNLQsZ5z4AAzv0YL61EAkRHRdjiSmlfecLPLlSzGNo2EznH2vvSu
lti79bOrszOtEKTi/7UTja/ijiEq9Mxd6H2dAxBYrCoBjH9PJ3Zs2PbvcqnHIFJQ
2YsXpcerHdV72GWh//ulqkM4mWOwuZAlKPKHYpxZqoouLMCdjb/wJsNRPgV130ST
HyrFnW3bD47q+/tzyRVw+fBTDBevazQ12uoLBHN0D6JoLBTJ4yDVsi9hJ9WadGUu
BF8cwx9OFf4oBufJvzBGu6TWwHYYcKsze/nb9WYGrG9AvkoRf246YTRxqL5AhPV8
6A+X1jgejHn1c3KSbwA5LAtzam7GEdk6QUF+DMAqGtNvuwCu0UQnjzCH2nYtggOI
t84b/KNrv/0CUd99YfoeQTq4RJWvMXnOLs1y9Hc7ChwnuyYZpzBBm3h5Wb+DNPRU
xLXrDal7e6Y7dOHTcIWbRvKa9RlFaaevMAjmsV0mQrhQQokqdqi58FORvqvP2dyg
Zky/gVtSI6ljaKASLjbqXCabNidXVYgRpghUsYiLx3vteG1d+PmlpoNhjLG110uU
FKkClidrzB51/qatzDsWVg1Mvt+Nw9IMyE+AeO2r3+I62ox7AItD1hXkPoZWmyXL
ifQdT38/4Cit5ECbw2m2BvnrmDWUUfmO2rP6n7zxKj4Yu1GNr9lVTRmkrP/nNzOD
aqoPgU9QYeZpME4EwGSE1E6kSQZukUw3SINyvDAoM+r5ajrph00NVzHsQPfqMdES
fbTkGqXKw7Ew3YG3EqoI/wRDVWi6PeEXzdIaU7bWtCBEoK/0l4fAZPM0YPzBw6lU
dtmR35E+Xhe3jxkPMPbPvcb7dnt6s09a4GZxYLHy7sRPjRPGOOB+jZO/WmN4xg8L
sS98+Sok+OyTp/kFSXyIP1keIo7Oe1Qn17vWW3+9UMLBPILtjUWaYTT/GQ08Wsqn
Q+4aaJCrqq8Dv+vi0mHPNnBWFs/I5K8AEZNbeP2NFlxjK4riRbyLzF+eJ5xS/WzP
DchUGJX2Yte2k0xYbwtPE8t0qkNti++4432uS2yXaPuY7R0NJBOKztZ+eSK1H62j
A56ftolqlLleJkEGzFEruTkBgWQsqOt6aLadXh1Uf6vlLiTIfLgA2B77eJgxTh3Q
D26gSpCiijvVSq+bsLZVeIBfU8P90HrmMRqBxbDdJJSUtZ9tV7EjsF+47gjkDFjo
gBSox+KoLWqZy4PXEm/W/dl4YggxufJBP8meUY4uu4s1Tqo8d4vpDNzyBNFe4O/C
rghfkQdzURG804pHK2XdluHdPzY/zwg7OkWkIS++XEDuenlnkqvd6iLbLjWLJifC
kz+igvm/bm/x7WCYwF0sByJGp+yqGY4TVtayfxwPOShxh7JhFRSqIB5aeX731qx5
RFCCd1KaxEYITW1QjFnyyyGIVQ0hxZxmOnUvZkD8x9uo9mHk23TnWN7IQmNxLtr3
bzZC5wXjMGZ5XMGJ21kWyY2qmOfMslSxZyGg6ijznSWUCBFVBjyTw4uB1E2fx6VE
PGd4S3LEqC25dOiaOgq2CPGpTLJlZjnQfKwOsK9ExNTxuqcJ8J0Mn6ob/dHagFOA
wg0v8JMCMBOzMcCOsNIG6GU1/8AxGwnxpTN9m5aNMVmH6LIliDOWUPHRGSEG5ess
WzoKcxJs3Gn3MfSfYPIm4uerinIq0n/UJtJulx2Wj+rxKZl+d0SlC5qVCcnCCUvI
ngU/Dx8ukAE+GFVYiJXmWaA1kiE9XsI45auVx6vBqNchD94ZQnDfOvfd5e2e23cD
Pm4dJE9/nWLORD5FLo69GtsVtde1Afj31g4POGSyck8ZsawcEAwuEv/DL6pFAIoI
HaHs2BXWlEr6Eo5zQVYblMWqRh5xhws10vhJ9wWa7P3o0FiqTGq7z4r7bfXSpR2k
6KMYBC2YXBtyHxLmiQm4kOG8+o9qM2suMeqGkjQjXaBezvTWoBIQu8nx3ENv07+F
j9sGcHqRrKaJ7Wk4r42QN4pEm02zvwEQh61xQ6FFY3p3Q4xN/Llzt7+Py0PBND0r
TriSxcu37RKpgbI/oxc1X0adQcRIrtfwSubPTFUpTi3Ngr4ksacG0qIAkOHuOyFK
NPGUfOBfhKKzcWPZr0nHwLdgnWi7o9NnK07g4nZQqQqTvI7Gvr0I77Pil+i98woC
HI4LDCuxiNd6l121JW51KkHiyQp3WW776LBiJZ4mKbvNU9q7ayYGSkFozqfZdzwu
PhZE/lxmM4F9IytU18WtpsaPuy8IlORontxL3gtqUbKmIw+7oxDBDMjoztHjjdkO
lqTh3xJlVPJlS+QtOlP6zb/41knkajARkQoP2maLB1dUdEuLS38BxWKqyk5nLUTI
OzXuQ3Ho/hQ4qkIzR0ym+51WhILwD2avXYQ43m3LdcyDmRFMcBiiLuZ5QyawoYrO
RrSBrpvcrWzZKixB42SSNmhngvOLqRqoqnXszf5S5lB5U9KTm6QjiHQ2gS0TyMeG
iVAoF5lqcQpoLOYOkgtMU4oZvhH7knO3GXXVy3uhfj8yAm2UCucjn9zzRigrFOub
9FjKyzylVrkHb+6sRCRSLvPbU9g9L16/DuRY4OHukzebsRGffB9FNHNOByePElIu
BW4SRINtH3vfy9vvF96+u4Uv5CtLPjUesS5olXI/eWi6aaIyiZBGr8jgjoC/MvFW
ePGw4PS+swfibK4vWJnQlqrW4mA8tUaoIicaHQK/8fNNCOIVP5pr9AS4/j8LQqUk
leVHq45fd70et3CKOv/AMA3f7dKrpT1ZUU2hkKNHi+WR8A50/xiyJCiPbRvOgJJt
ccVLFBQZVou4Sk8YJujPQ4JPX/PwMByLlY/77xLVvwVt4qPAKOCnQg69yXY7cSzl
XqmwK64UOODPEmSyo0HKs6DdTX8gieIclDo4Gjor/egzh3ox/po9+6+o8ExHYP79
JWJ/guWLIPppn9JCOgIDDw4i1J9CbDeb2x5I6a8o4B58H/GLE2VaobqvfDlT8tkE
UsKEglZmgltE3mshGULE4UH3kQ1h95iKXxutMkOuj2W52Byj2AYOdRoxQEwIFDoC
E0VNLP2xdzJamBBp6DwrPhN4A5T/nRuIymG5/DM+tNvyJF5lOtCAoJ2x2f7gH6be
ns8q9GmmQRolVAHDkyoyTxxQAm3PgkBoWvuXVu0EweOrlP+81tKSVje5Q11A6/ft
XbTeG0A17AypREilmJ5cwwwoAtdK+ne5wZnnIFwHo5zjlrLCPmsVY1KNWG6hdcp4
LLaXnCCf40zzumeKtfJgQg3Ob7BT77GM94YNgKzh5SG3BzQ6H3I8P6Kqq/dYbRbw
v+rcFfruKcgcbOIn3q8ESbm9nEx4sj+/HbqcVYjCGv7B3GcTETjhgxaRI10CUHII
2VGkTWnZGeKmU6gLZx9dr9Y9m1aMev9ur+Zo5jOsajU9+fihcKe7Z/MSOb5uZ+yt
vqMnO8aETyd572br46b/qR5V5jgLw/XgrT1YIzzQ0+83ygsaHXieFlKBqnaUbVTr
fcw35NUFSlvZCvNfsz8+66M/9wkZkgcKonjYyB+9JqLsRQv6xrTfSi+Nhlw7ZtSQ
4X2WCkLkEvEsBJ52RzASN4OevQQdHAod30b1hNEWVNG6nYlDA+EJJRuU4hnRAgGT
xiE71O8tPPF/VV08QQ3Z1xzcZl5rAXG51TkfVZ2BjykbS4nXNjFgZlgLI9nVayj9
dWpPrOcB27U3p1F7/dX52lUJ3POiIEMkiux5iji+CcI9H040LqjG9RJW5xWn/j5z
oltPtB4AeAFbzRBjXfo8/mxePrxN+g/ukFNknOABneSDXXGZ10JgAepb9nJGBB8u
Cl7P9uG8+MI+loVAIJ7E6h0lpoBaBLNrKmNlNfmnZmua+3QGRKpfShPI1DO6U9+c
ipX7oCQIXAir6FFSdebgtBju70DqBQGXm7S/NIWRNWCiFYA0Zh79NY4SUBtltoWB
6H734rSSj51oID7AQypItN5c2WkvigQ74aBOnF6kbc2Yq0WOoS0LU+vrEUgX0t5k
ntIBUx4KFS0gKt7KBlyinFCL3krWR6vxsWfdtJ0HPgmIlEdwi/PLDqbHTNEogIaA
CnsMqox8B13YU4Fo0w6eDpxYNJZN8ht/08OGUHEo/XGkkuD1GCctCY9Zmo3KxAKp
M3Fge+PyNZvaBOfofobqnGnxaZFu3toZVBcZH+B73U3wceQ+bzt4Y/Rqz0eWvml/
EUOA7/7I5DDfBgHoTLXCi0V14sKjAA88f/wDHaI7pVwNKhY+DDu0J61r02Dw50HB
CVztO7Ohl1IQAF1JtltcqUNYTiO3R5vAJ97RVuyObG1s91X/JuCrmMugKBDAeWd/
CvTU9KMUL7pE0Ie+9zmO2i62qZMO+5FTe+g2Y6EJos3pKNyZaSfDpVGnMNmfdgMU
BYux72G5eSq6T4dlt9nv5mMH/3U797Qc7G1z3eUY3pzdYAzg4JtabFbys9j+l80x
cHZprhsbk5p0S5UGCGyABg77Xfrr4vipYFPvH3KOBYna9ytLZiuPWSDku6t7lGuK
yNVe5LDEHv6Sd1nppoS/1FXv+8eMCYs+pEI2RbHe1Y5zw0qc5R/g++mzigaWrW/f
E3/5aN7nP6JqFTsJnrQh3PrmPWx+789d8lQYrBJlurmYIdllRVXFI8jY0tB7fmMp
2CKp2iZ3JME1zMkp3xy9RrJKtyG+PsNb9slnKCim9RM4x2Ljf6Cpl1+c6gWPtkjh
eajduEzxjbU9WAw7VyS78KBcfo0fIQ0cCSOuNb2gOXDkXOuuFi7J3Ef86NYWbxQF
UpmTCkkrMX3VRs5BAkQbZXebeWP7xKwuvOHJ30QybNlVq134NiWri7R6hjvgG30C
5lj4H36XY0vk7CZwpoqejOPlNzqCE1P05lBQQR/xGYtibVhuHGSAK9BMxSuFBJ7x
2ehJKD6F0lJxryuBS8pcGoWlu2pqkK4YNluCULPSNg7tLSW2gSAN4GsOt9ojjk06
6KN9CRZPlV7thUaBt89xhbV8mxvTjeveQx49DXrCqOyF0mlBNZIeXKk8fuNRvNc2
s5IFyunDksBZ9aasZbiPcn7PZQbnnYXeZ4YWYAfn/zz0GDFGrOJ4IAuBEyjSSrSZ
Eshxj3jkrm/SlSH9y68tXSc6SwsIqsqGU8TVW2wReE0QQmyYGrRfordV+PkUPKdG
1v+WmZwgG/sSEjc1qUNPNt+gwFxQsWKdZQKTYYf0c5XvMdc+GShVSSBxCVXm7GtZ
hwwmhKcsBGToHVCGIGTD9XXwih/A0SarphSwJrUDc7h6c1GRZ5z0YWH45zbn3LM2
qY4nUPvfdyghqwqhjxa6jxpzVHdB9VnNdGZyz3Y7GMhUHc7ZB0j/y3pLHdWUFzbY
F7Zb9dio2bSsBBwRHrV0niHlxxg+FQt8LlgeiRTFh2EYvRocUqiBx1JHvibxzUt9
hpOLS5osmnfkROJWxWcRBnP3/GPxZp92LziWG9jEtTPhfEXn1A5yc02CjhDAiwmg
1nEf6P37fDhE5qQMws0f7wazYFVFOWkow/55tzw9Hv6saE8ld7Au/6A5hcDjmuVu
x22QG/8dakgbXXadZpeA17Zw8J3qcc3kVHZaT5A14cUHiKZZq4Vx8pz6VvPME0qg
TbwIxOwDMlYaIESpOC/MsMYBJlCAcxiIgkQIdLKtEfXfRhW7QgLvLkxND27O6Ed4
ziQzK06zEvR2t81GyIr3tldXVU1eG8u1IY36s4egwOtjLk8xbSz+Ttzx7KeGv/oO
bdsxGuF/AYZ7lMB0t3+r2O8HVYtI1khkSyfV8KAuf6oaE/6Xp1mAQSbqcSkJS6kr
iOB0uSStc0nc4vSjsR+Vi+i5qXEB5wi6Bt/nvjAM8KcBPilC5VVHt8ztX1TIIkeb
NfTk5n47TZ83czkHaMeXO7wWS4s5WMnkgsaipDk/UEoQz8N3P5lUaFEez2NRN00n
LqzmMGmcIEh0FmPJszxo19e/JgW1LG69Xpc3871UyR1vh7aMFia+3ZgfTuCo6S6F
zNSFO3QThFMo89FJYHeHy2M04dk8sX1lwmig4HFwGItW+MFS1fLg1grs02KoLEZS
0egeXOseN6gIx8RW2yN2BeQW4HIMDlXZ5PcdRe5w1R5gFo6TGeMCpFi8veaxi6ip
tGOTwD3lpEMgOiinbXjXIfOg3NttxXPGYY36yZOZyoORcu/Q1uwqChzJa6ZEyNPg
oXAsDx7aM0iK4/L9ppbQdUfvr9iiO2szdcicffO0bi14V3j8+IEr8oBR2oS0YUe3
+ftDou/DwdBRP9pkgrBNF0CT7uTdyp7zGDormPRHhF5di9QdV6W3U5RBl0rw+DBg
XA6+7ZYXkQCAHjDi6K4vNZDujCtCx2cavGKwTktwbVmAAz+qMFgkpYiwrX5slNKz
uSDadCEmdtOniash/LSLfYrH/gSrbhPRgLjYCrN2LuTs1r1TBTgko+l7kWl7vgPO
3YPPGpPzxVq1ICU5+XL4U7Y4+c667llNE9jv2hNBfZ7ZP2cLbQUcZcX71vjYrUpt
D7Q0RV3aW/cihWaWmOpxN9ZWns56P6dgxKkVf7/hggZ1xLO74IAGKIb2hSqnfaYl
C75TLeA9DEvWrFARPCSKJ309oPUW4h3O+0CJg2E01HD7BL7mxcpR7PSPwCMaN04p
gWxwc5KuPrkd4hg8CAVare11FAXPjc5Ws/4fx2i4VvzBolg0BKQIhB4bHF5fxpJ0
mIi1QZWupTLCfrlM7RW1k4n49xy21vIUttO7WaW268gfuDPJbtJF4tlY8HZQKlQc
fegyldXA5M1GTSwHs/0vGzsuRjMsAM16DK5yDPahlwNMWyg/yR6We2whPam8eWJG
XDk9NDPASzFAc/+140Xsm8mpMOaygtuDVbrAb/DZmD4RgVJ2C7fHAXdcBarXrbGH
32O37h3dGPCziS00kOsZLAKbi8vCnYz58W2GrdlzVSJW3lK/oMskkZ11BGklcBiW
fQsIKmp7N7nhsPuUOX15hSVQeq3el87Z5ARC55dYY6j09lL2FSVSoWWDig7CSOV8
k16ykeLTXuHT9jZiQ/7F7eYJREVaqttVlHzRS63YIk/WGFRsg2bhpvtm4jAihrZg
umvju9wOc6lvqR5GbRFSkmGsRuiHIfZTmr/UB/zawLKOvItUQvL7yoZsVEDMjj31
8+BODTVIOEiGZ0CmEMELp+wGNopEh+u8y2XPf8hmHk14eeNrgzxvVCQ4mIfy3Rxt
f+nuP2YpMZuz9BE1i4id0jhHyc0vpteQ4b4+ni2tNiGuz8R6oUIIxyLUx8fxg+mu
jpg61SR3iOcgL+LIsR7WdQ/OXKXxNlCVjr/YWfacaTdkMb8wl1cneNM3+BF0UF9v
SqDF4dlRmSCdckoSl56NdK2krVktoDdIWY9QchMZaiqkttlEOWjvvcpiHACiKcUo
GhQjgfxnu8XvV+sNoCupB/ELQQa+xnBeGbwea9TERtGF6vYyQPwQDEnD/XUszLI9
0Oh5lRz5wAsbZSC2JyJvg1b1WG6W9N6xKzdYOV42yEq7WzGkzz6+2gwlL4pbbDEX
r+g0OpRVfX5foRdk3JLeAa5hs4uC6SNuuSzwvZ7rANwsrp1W5Wa47q7SyZu6G6LK
a6hAO8Y9uiCxvrUeFPOKi89IL9InaBO8J/gBhawVymKi6MJL+IEsIGmntqNiTZbb
NE10EbBAu+oqtbjGRAtd/2OoHg3GKwltvZtCX8EJWNoUGwwvK4RkxdIr3SqcYnJt
QkrfYLWbSl4UynGVD69wY6XeFyl1x5XJ8bfKKK5LXc/3THr7nQSfY+dvOz8MD34h
EhVcLJDfOE63FUB60Thi1jnqq+VEFxsE/omIcNNDu7c8v3jnCZ/017wO52xNEk7+
OGLUdxVIaT5t4g4NUJyF1THXEUgeTBgpryYD/TJPaYqJH4AWvB0PD6AfeFbA8PVX
3LrYALWPPuH3lZvh3scRK0M71eDjLww+6tS/VJAogIlQ9krqwYvL128uljjH1hxi
rN/sUhTNhNwnHymqi6/ghJ7rsXfqyCF4tu46D4GiTyqOs8meM6ABaPQNKCjIAjdk
tswgYuNiN3H4KnFGWpuKJ6H8Q2VK7duWNVjbJNHUD4m9PNm6lzhSI2WQS9b3sc0g
elBMgypQWCdZB0deutqwHxQa6tzYXlpaItOOEZ5mtyD7qVpc29FvDGoxhqG3Obzv
gFq4oTeu8l4ok3k14rET/FAqIttqbybgRKDdoOCr/OsFdczeFJsIjXEYZk/6A9QS
K0TTsj2DYZV0eOQyX/MaxXcU0sTI7ZN29jmto5AN5Er06uaSj4xhFT5xLZsDkmBQ
yj4SvNwBcnNcfaSTI93Vs4K71Q0s7Znq7PQcNHCqxWb+Jn0Bc02GE+YjfxOSCTqt
ge+nkOwXRQqnZLf/zWPER45UKcbQtTy07Kd/6bfUbhnwB00uu2LUZx0CBeTLdIsf
zNqosAiBckBQWp1rh+rd/ikj2WjOlBAXEy9R9pbIYwUXQRRgywevwACWTGs1oVmT
GeYav7Gt8x++orNC/0q+0O3DJT+gywC6veNAmShki5S2HPwvZfLqBYczRkIQVkHk
oJDe3rF/ZYS17dwfrJco7Lp4FQ9bnBhg+mmeP4migMi8/XxABRFzMAxl2bB3RlVC
CMYlyGgPzJjgSZsxuoEwAyHlMXI9wAoNgpTcPXC7V93rYTwzlxhN3YGMJskwCBSh
nf+CS50cVSEnx6yVNsGDJMKUhv+5+8GFyV0qtEMjYuF7expsP/SkSKDrdz1DISu0
nc4alLvnjEayFD8wbPlyIDQnuwHCPfWs94Ejvqr4ZAfSmbH6e5mBr+NfURHVhKGs
RPle0BQfgRqxNgjjTXNBFiGgV7z3aQ7eVK9WR+2EbJUwEVhPjmGT5RVB4+Q4rttf
qw3Z3H0cJ3bKHovNoBhqHUVfGzNvRKm4U50wKH+0xLTNAoY7BFlFBIk7SEmyyPiJ
M3FFtflV1eCwfjAwD8r3KFdKmQ+S3SoRm1TvSRLwjF2V0yznj9p6fvysaouw+rkQ
D9AYmBnQPcwqraLeDAGU8RKpi2zNSvhafzi1l2l+1ZMQliO0NruPsGv2I/jWyBHL
H3MJt2kKVToncXEavYBWOlhPqAofdm80fwzjN9CjJjrS6aYlA4FPF29c6A4ioJgC
WjHALsynYYVGPfYr3OH792BJlIJPmmdJVVtsf3DSaaZuuxGRTgIB9acwBUHIsiWZ
ShgffzvlC2ApIHR3T/p7jUiKYffCpc3GawzhFT4gQR+fzGO/MZJJRpjccuE4sB4O
9NgZ+R8goeUgjE67fb9U/o+hdwPkXBcJ8fKnG8ThZiuxedVrsmnT5N104JgzgV4F
05wqNvsZltKVE/djO/muGmo0WuUYTyA2u1fS/lc7a7YSUe/sSpo1Wkdx/Pmy5r2C
roqQN2IMahh432ASZWcSdtVQi2b+gbZN5sDVfd9LFRnlNJIKg3SWQBjooZ1UCRr2
ov+BZXa1O9iQ7gSrrBQ1QjuCUMssVHtfpcR6sf511Qd33G8nTlT/Nrkg0VWZMNFo
9Wajh0zQabW3zG2U4DrWoaJlDmoYPlKa7qseqKooWjYQBmz97lbc5CPteTET3BOZ
alLEDDvj1xNiVvN1Zkzk0SXTne4qFhm+FxxmrQSBnyCeGKyXDmqlBYsTwy8gbi32
hdX+ItlA3lonO5FJ/6FMbS6+JYCy9dsrIcxyS8VMhRo7JOQae0HhwF0aHpc/ZujG
Wo4+e66Q4i6Gm9eKYt+klQxHsnWfIoArXRC74ObxWMn58YDU4/U5IZV5BrdEGUgB
ZQVBTkVxScN0Xy9MtrEOUrOYdsZvD0FKhzAUYLKNXQIwTMoIJ5cpvuIhk7i9yD5F
JaZG1WulPcrNCPBv68Srvi6NafmGcx1pipmi/9DMMvYWX8rxw2X9SJ+xI4vBXn8q
lPXDrxNNAa1hdyoAqBLT+7sc3hh6uLttWfPNpXk/OYjLI5es0qbva1j2I2FwkLSe
D8IKjD3sQd6wXmswsxc6kn+48CXpiSeW8KrPB3lFTmGSoJ7sEii+8+KquX8lIkzl
bJBUJQB1V6E6bWvSLIw/g0eiqnxHDXwwN9gIvB0/BxYg35AhmIRJD4VRssMmuQOx
8n/3gm6gIzRegxhrfxINNIv8dJUqAyqRdWzw7c2jaKm7gpqYxW/lR/+5Udd+/zQ4
CYQRYm1zXFCQ1Z5rkGE3WmZTrm3fSjsPN6CnvtDFh+lymurwgfzc2HVSnLtMwLmv
YXSnfj5dQUtKWEAGEybPHZ9nXujrxpz9HFAnRUX2u5JyljEm9bAbt0HxP9jGEV35
Aj/rEqIJHw0RWbAZmzOgZpJCWrIbM5vzMQJO5M8L1dkJamLqKBS0NA1a0iG9u9b5
E1HGiwko6xw/I+bUfLDUWznu7Rp8Mdpwyl3RqSk/74mdqk7mJBipL/XwdeQets3H
mZMvwYYoWsLR7DFOEItX6p/NYoEsSU/KXhbn0Chtkb1zS2bVDPNp03MsCtS947Mr
syDwSqnRzoXbmNcNOtqTPqTwUCyycmhNlK+9EbCaZTHPbPDu6sRe63q5l5DHlmxH
96HuUIY6usX5b6Hiikvqc3SlveWcRITXxkCidWAT8fqtFIcy82hjuAXQAlg1cZAi
n8XPyK9NgIo+luheVRxOhbTbr/HIob+FiXVxjWxiDFxyMoA7C5hl6etvYvCS/dWp
UGt4ohrxFHIi5EmA7y2cE9II9NDbDDEtEXQg9esdUkn9dUtNjYGJ8lj7TO6oz/uF
4BhyGoblds9+UneF7Zg79I/cjSFn6fIkL5HxIwna5SjKYttRdojmj1Atg+1lJ9C+
N+oRPvPa0hLY2rJw8MshlR13+RUeMdDXVwyUj7C+aFWACka49/C1rV2UX89G+Jqq
8lEnp16DR7ZzeB/o+5vcIQ4Z9W6bEkKTmZ7uvfZGrWMtJ9sPFlVj/FlZwl7/xkR2
ENGnCg1MKxXAo+tD/IqRFxoG8BbXMPmGLN4H5d4Rwib/ueryXcLXzmTIeobOqr/P
fpTYavjuZ6M0aIbh9lG0T6apeubF4eKmqkwRujbRBMiuxR8/vfpnpPg7f4n26a6L
yp2NfO2CxLYPwkZDrcoqgSa9KzkKugQHSRiY2xGr6tgbc7L/naSg5O82nHkAhgVx
nAtxLwnT6pZFozvBHrG78rtDNrqCSMP3hKXF0NTbmkcJup/XDbFD3q9JU3jnXQBU
V2yVWbVeMo3AOBAHQ8OGV2Iiq6o56qivasFMainy7kQ9KN36MetIMYkDAn4mUnpz
Tyx4sUKQnYsMkxpH0vjH622e2nXUXW7pRiPRar4CLYLpTSg5K1mAOEVAwQ4MIJjp
peX8xmIODwPrYh6PnujJFmwsNFAitoNIekDQ9PePhHDwHL0I5t6NFQYJgiXqJrhA
GM/+p2rpIuuUcXiWj5tzqUReaj2TWTOFMjtSJBEtvilLS8JBlhP1/bgeRzI9fPu3
1YxIsuaaJO/BVOX5FR7CiBUkSZtM0njqkVIFjDAcAaeNq2n+YFyMRpnSjALljSkc
GdOY8T58LQVPvg/Non30hCR1ZbqW6ueW4gLHQUnAozTzvh3C1FfsH73LLdHTCVTV
/YDizd5MnpxjT4FRw+r1WiXnLcNZA2c89uT7FMdQRUzfbYz7cBNhiIPR0bw1+MP8
fMGQl7eNh2qFk4gbzo36IiVeVIrUggTJ5yD1GMBtXFR06dyeth2d+vsYpQbmJ377
j6/apFruqj2e5KHbycBmFYUXYBoRgmdGS3J4mk4CA0mB+AjY6K0CxEyZMFJ4oLGW
CXzRrZ/lFm7/qkstkixZO9E8q1DMgh5U0XY0gIsA/rgMS4TMNAkYkh2+4Lu1bpH8
GiJ5X2ElylqAMezm7v+tSRsdUKUwn5f4nPnGZtOx2zFFGmZRUMXmrasR+Y33+j0I
frhzvYFI3aI4DEUuJj88FXwvHKmTqy3CgRhJubMhURoXN8D/t17yr6vlUAcVCyhT
mTTD+BVKV0Rwe5oKe7yYc31HK1q5oD3v1BbyIPtwHj7ohbXIuaArcXybWsLXoo3f
5j+PhBzMg8SzKidfjG3pWZOOh3wBRHXDnTEAZ/Dr7iSzfptPYRHUpfdsmlaFAMaS
LJX4hHjTOUt4C40wNN4NHIsw5tjQiJhuMwDxhPSwEaO9SBhGuTaiVtpGM+XmdVAK
y7wStYpcE5egQzhkYD87VCtIIYwz4FGWNYLKft2o0kR2/G0ppXlkTqb2ndW8mrbO
eEHcmgdIqyeDnVzMPt6eozYl/Afx9Zst3RpacZctqCdix/5jjvknpdNIvfJbt/E+
k9UWGVuK0mxmmau3n1TUK2/A4WN67CSVKQk78fBHayVhuMEK/yD+yMSOPqbYqczw
A3sxrut6dBEdjzqV5DopPLRcOMfKW4UuSbnKYFwdrQPPp4Khu30CqDNf1B2LSPoH
Kg4pKc255jWfAummfCrmtT7OSXmHtWxykTxfmbcUJoDkt9PSNkZ4rZ562edR5pSn
PAkEql1UrR5I78ehF8H9+PLftzVzWZ4BRg97xkLOU5ce+2R2yNVKf0GzCKy/CI2Y
YZflGfWWRoyGEVrvYBziUYCuZNAhfMfSk02UfQoh+B/4YjHdY4OqISOraGKPIR8d
4bAxYlJ+bvolsHhaGpX+46Nhl9dHtFyG7hUjNHDDGEkRiCjR/KBJ1IBdNfLNqFcH
jtSoBzRhQuQnCScRcJCL1F6JzS5N76XY9fdsbiy8gzpL4TbI/GpzSy7/9Q4RRAF/
H9Dfdc2HjxD+EJKczi9s214r3WOJFBQoXc4rhAKVe9j0/Tr/00eOSwofzNeJxLGx
dnBZbbTX9YOMxsmmMsS9Dq3sMDFwrLwry/OUA7kggoaf1pLjgQCXaAp7d/uWaNhj
/7EGfskjYr+A4+N6oOjzvERp8Zbgm4ktqifBE2+SPMM9KKy/ezbTNnCn2QEKsiid
C+uVApAbKBLaWx3TUXO6XzpI/9jQ3Gadk76h0J5B6UxlPqJuAhodaI7OsUB6ko6I
NkfT/iYXcIPsns7UGAJv3U33dDugYPNcHxTWBy5/iypZugKs1WvC49EwpQHiwuel
01BzSrik0KgfBEhXSLSgHt0kIbMyPH72VHdpHVXAvC4sQgR6j7TxLRd0C2p0wPRR
Yro2HBYw2igMg2eZbiVf2A2b5s4+bo8IdPXbZEJBAVUnhjqTDw1MJqvCFlRYE7h9
P5HwOJHmJWq/FzfK3KsE+8izaRz3EgVINJoTv4w+R7LbG7/b0LLcwNuO7X/O15m7
t2M3F9vaAhkKoyc1xY5cxukaNUl1wvNowtY15ohBte4Cbzu3PQiycpiNkoaGF3Xy
wjZC+iQZqNtctL8mMqjl6ihlxLEcxxqs3LauR8ssYzlnjyknrDvmNhkeL1ikU7bB
kH4+jG2KWfU3axYXW4pVvdRwVOWVv2IK3VjW8DF1UBgqyQKRB7qnMpi10/h8AiBN
poNmM0O1bajv5oqxdlW1wMq9fi8cKhmjDBJKrsSbFh9sakT29x4YY/MK/P0tryjR
5ngMLpFsd4jTSv/npeYMrI1ezj5ZyzQVDiThZFnjbC5CeRXPWFZUt8+GTZa2BwK5
S/Y919qw1lbaYe3KgVcWKNVvl3b7qUzz3H1RHudElWcYCNJQmkd+KM9UMyPKlyer
T76a/zIGlsKCFPbzgZBTL2Q0XwjOi9BZYtm43S4ypzZhnBstYQkpEccKlp8wWps0
ZO9zQwAw+oLV41tSZVCCamf4b9qyeCvKkOXHuGTShxQiDIf7AegL2ZTz/6KPDN58
qmWOsmfE6Mei3dl3jAHA1jHE8tgh2d4f8KnUYceQ6SfaiRVASrX0aYnHUE+ysMBQ
1YCZdegxR4iM1S0oOKxsOT+TtEqufaOusCkA7g+H7VaYTSj71enzVR0mz0h07K/s
IrkmlN2gk3bU/TgvXQC4osH0eaaC5TXW9OObMOl7TBp73f1DCOQOA9rM4777z0ad
UgX2pRhzh97vfxhU5p9rDQzMFqn1wD7I/qMmSOCn2tc=
`pragma protect end_protected
