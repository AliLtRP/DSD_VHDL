// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:52 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QXBCQjHkh6NGrKSBIVh6UqFRqRkUBu5/pYgsjfRZKppnd4izuSJAkoG6c3gliHtp
aQTNmb8Fx3L/kAP9SugnoaiGKfmKEDach5ZSIQp7r2fuj5+PLG5kmzpNB97BYgDa
MTCnF2kbNSbhD/GJYSLM2Y6R8MIe87tiwZ5Im48XgNg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29024)
e8an2bb8i7V1WdD1SXV+NDkniq66DHukIaT4ILb+Xp1Nogijc6S1CH5BGSQ9ak+Y
3t8EyaSqQFf6OayXtihUjR7bDJAt686odBq57RsDOrlwg7BiyZW/uhrUB8SmVZhj
I+ul8qhVUsJR6yVjuX5CdMnpZIB+rROxP4FJT/C83bM2Qu4DgfPWlNHrrcbRvAKE
EtKjX8srIPVcEABYn0HXnrtvjCUOAg6ZZNKRPN6mzs+Uo33CP+ZVSlGeUdsQPCQT
/2LXA4wASy2CNiT2s9lKr+QZu2zZrxHt3lSx0iMFzSXmspOhgua9ZmAp2MD8M9JF
TXiqIazpd9epKbNx9Nv3xsa+sGdzUDhM2qSm2xu3ISIKnPbcbuNYvqFd3Z/uA8TX
sCnsJNjRLULy/u3MlthkelxdU58lwlrA99xWaSuXWi+xwYgbT1o0aTjyvzOQzXqW
HzuYuW3duBmfwji45jpxTijyiTet+2CwAFkHeiodF/wLehBhSRzagiB1TnSuBXGp
iA/NHJvRY4aPZTy9ksXIg0aYm56NZaGBy8TUAPhIJTzXj42xBWBVB+4+Hxkn7vo+
k/aaAYrV+ixow7EBBOPgSbapWMXcKX5KXoFCmMvXqWKLjwtpMVWeo/wFxaAPxbeu
Ds7UPCx2AkUTlhSlYC/mJHwoIjn7bfyaWakkP5r1Gf6ALCLZKSenu7hdj26CBglV
2wpB4d7rcN0vQM6Qb1cy4Z6z4wkFyiXkG5/x6tN6indcw550GRjAaSou8TeAkRH3
VgpYSU1efVbVoSpqdFNRFvr1mWXLFHlK19SfxyrLb5SJSHdysPqqzyG6iZLqQ5SG
nkjS1AGZRwBwGumq3v1seo+e9ltKtEJwjRYVeaQl/P9GvJpr/o5hA5lna5pvsowB
S9hpUsEG6x9k2/HIDyJ8Y/plipksTnUSzNRUs2oyGttLLOLhcYTT1UY6Mc63vmHO
ikbQzmmR94Bhs4EIxzVHd6ZQCJzGjWnPQoikL897J7PpJVDzsf97RsJZrDoA8bqP
JTOTJ83T2/D0BXeT0ZRKiVgI1WICvP6HR1Yw1ENFSDqHx0horg+8Z7RUoU8OPZOk
MO5LzxmBS0N0CszPyJvy0LGKkrEuNLqzxd3mQjoqCMRe700V8AlG6AEhajusLPkh
Pt3ziaoNT0yiVY1l6luQBisagp0hMTmGgeXkzp1HyJ9aA9DUS1Ecdcc83HOZV3tw
kFpsPw8KTzc1+98BHVpKZcsNqn9U45FwXaM/yYC79C6+JHIwKxxx8A8zL7xU/nAE
qyBG+kbvdGgJEWZY5YCK4szElVIrw36f0HMrs2moBJHTQLnL+tcByU5WbvoFt9Jf
qxOTz6JU/gvay8q4QsbCR9/P7eA+2sxw6sgPuGXIoSn3q5ohMxv1YQFDEjXFHzHB
vHaWeijys/aLBQ0mTbG4xhJoa+Wotu6cs02f2d6v8JW4hyJf5HHe5/yT+NQDbTMp
NeyKk9gQa95M1jfgTxRn0ccwndyCqADavbf73rhov4LxwZtRUwoy4y4xsF2hLNL5
ZosJFrXvxqpd5oBvfK+DOSMC6Km9awLWFRMj19IYj0yowPbk3jJkkFlvwhhTtlIO
XsIx2zmiLM5i7rtELmJCx7uptjX9BknYTpWd0O9E3TeIEuY+f3LN0Nl8AaUq9ZzO
FSXWlIp7+ebJS7uS/TPYz8DfeDHsjluKUgOi2ANyfYeG7y3iKYu+UUX4AXflryCX
IpJuRR7qMhlVhz04MkpG0MJdh4Mu9OFMHN9bbuSFEvi4VXNY5ru2d51XN0ttVsJM
hYv1BAn5Ab8uPTvVmSxREn3ZRp2+HSc4YCwNTV0GW9AjXJU4yfMpik/MBejGCX2Z
7HTIQ8dezoYxcIbf5DDtcDq3bXk7T0KLKak7fmHPXvGuTBdGnyrv5IZcK3SkRRY/
Raomi68InJIZo29V1cbTiMizu852ylfDDDb68qNloJLGpS/WGhprfzam1yhPftOF
sJ7H2qeG4V1kR19nvvQ+AAqiY8KoccBp9ZIYneOu4MTN35w2VnbffVEBp+9CJCtM
+3n7OTQ9ii9EKor120GWK50jMOF8KcZEBYlre9D9tA1Kox0F1K6WKv8qzACXbVPj
ARzsxRnDIy71vLi+5DUQK2zQtzBd+VLt/9vh3USCzzg7zGsVpJ0AD3jq+PfYXiqH
FXFfVZz0WXAl3UW4RDM/c6UylodEZ5kXEPyc/6+/NLfHslMEDBrFOz16B7mWBTf1
+pNd+1cQjpNmPOTlQwA6+DzZC5tBFjyVNPy3alj8JOzVKosoNWDox5fLmCVJzwBC
yxfBOiBNKhEX1vBe3nQN3FBCm4lTlSVW+qlX/eVaNj6XjUFwfEaoo9CZUMiuFuV5
dGPA+OGCxqUxbSOkA4cgMhBJKhb0XYHFW1t7lkstQRS5ZycumWTzbhIc1Pc654TT
9+6mpwpoqHafILNqnq8MXZGZKAfoNN6NShHedR8LK/D8g4lUHKR9jTL5p6kr9te8
goV1jp8en4mFk6IskMIgMrTwBPzPu9ZUH1zp74+bzHxOHcJSCY8xAi10TD/nmQrM
6MqA3jbdJDqKJ3wf4wZhobUQEaN8KDlfHjKKWRUDYuuaAmabFZ/hdTBkin7HxQnM
tnQVrxdQSuEXAlhmAgr3fFqofBM0lDehuq0T+CoYr/wNlh48IA5qg0XQ8/qTcwTY
7blbIsfwKDcKnP5cKnyF22PiMn3GpsqySrK2/Pi4VeEbM8G4NRSLinNfVnYX7oXc
FCz+ICLIP3AV/mwZXj4B+KWEtetf5AxihqiPP/Mv+w9odUCbYozvVCzMFTBQCpBO
cetNjDfNxEt6mNK0pzWD0AEgUX9EFZ/cEmfA9AgW9DqOW3eAg03nqyT3LoQMssV+
8cVW4ZZhoExezKrMZGOA08uc5fhQuzLgzkP3Dzha6EPlb0oWDX0rxG3CsUtHOyfn
o8wPhgT8Q5m0T5lWc7UtsmO5J5BntvQGgR3Gh3f+EH19xJyVVJy010HxftpDxXGl
bmjdkphKrJcmzemd+eMDeQksVRhFhJP7fq6NmN7klVxygYBvf2Bk9RaySlhMQH2p
+HfYBdB1xltu91/VZBn0a4tuZDJ8ay8G7gCGlPpqn66cbSLh7beFvRyRBuPRNH3d
SHXqCcpvIQ+koozqV09MB8/H0igzMHyqef0EOgTViN8W43aO5BQW0jyebAYX3jcP
CYAJ8HMviWsbzGPGCh7mdow6+DAj0Y4R5bUW0ZZL77YKA1ie+vOV5r8d0V47SFNX
4xV89kYsY3AVZe9pgk5ajbOJB8mTjbbRPdNQWvAtOdkAR/sqUgCf59LgNkjTg50u
HgUXqy/oMm5QmGUbFsoo1r1CjbmMJHWltnacWKv11XIPm2N/3dKqurRCbDT1DyjG
RbdN2KDjQ7jAC09SPsbokQMpWy+gXDFI7YJfoOSRXlYJRtLoyzjnDRy9Pc1hEJa3
UuGgVb5bTmcZCKFE+CA5SHISkzyoCKkq5npE3e7UUZq/bwQqAHBYavDHjXy/WvW2
7d7Yu9nBZhrl/u+lkLnUIZFjjTfp/8XihBLsI1h7RQnyTqIAClRa+Ig1pDU219Jw
qE32nbrMpYZlJARfgGo3T2JjXsu+0djh8+FpqXZGjQR7CzI3LAUq5vJIYi8Ul6u7
xf0DDjWx7pzCQnoNBAtUAXbskw4DHH0SRCughpksTl2S77y083umTU5poRS9TKaP
UXuhqOfeBHLjaeLIekAX4+U03hk0Qj5vjg92MZBaPQKc/WhNruia3XxeJS1fsd1a
+DoJKnRV/ik49mAAmK07wL0eRqtJHGYJIY2osK+sJI5KwiErof91WfQi0iSdriYa
XAX3SO8SEfNViouVqu01ySespYlL1dzc92YLjYr5PGjBfurOSf2QMoPbpTD02vR6
GSJFbcfAUe0qDOrcA2jjqF7lOJHrzNuF7ek9Te5lv4ADRUBgooBOKlZXdUdKl5Ab
ouwRsl28cvQTE1okneZCs217GJlx4TYy88KekZkvQeqUmmiE3ssCoT1Jv1wSsmes
IMVA4gjTmPnAebwln3tq5vtoUMDFhuQNVjDSZWNZ0UDhtdqVMVmwKxOyw8zYwlLH
G7fAU53h7XQ1YRKtZ/eoM8lJ9gWieLiaH5UoyDUt6SsFYHnjBKQljzFM4Nhpf7kG
qUxXpZYtFesnBNvc/6m+bpEka+hgOJ9X7uNIF1o2fnPUbJOfUX+kZdWbVtjIdd03
s+/2FfDM+3ilD2OBQEJn1kUHKxp9vGQAKONpeVOEXELxVET+QoOYOMABZSE1lGOF
gndy7e3bTn9BfRh7Wr+beyn3ZKpXnkyB47VMwcTL8gUHPxtMUaT7ZE/amqHnm6PD
E2zuoASuFCebdl4N+EIa2/JMjeJyShjaoTBLpnPFtstHVlSDjB2OVUCjPT6OaGdw
g7V/yvDfD8zHQN6GdaRRbsUysYSXvCIwpcpwa1IlE3NO1wQJcBa2NhQzdgMUlX9K
0iZY+zc+/yqYa6G1KBjh/f0wEdJyzODM+D42HIZ+/mNUsEplFtHwQwEYGogzdS5E
zfaKgnFTeRyuL/RE39aIIPjppyFjJJLEMRsccyxHakpHogNFsyfd6z5aEfGglRcE
he8laVVZHW/veMh1cYqC7AlyfbtHDKZH5fuCxuuvKfY7hILBOJf/G8Zt190mXXhi
pIdEGfyt4E2s1oHKC80cXiWheOuukRF5SfqFLoj1UepwwUARMMeeHBwf0MO4mdoq
hN4MtX6jQk8R8IyDy7F9mfHuqmC7dyxqbCqJ4z2MxvPIezrrjDKDylgWvnnI5vlv
Ojislfy1KE5TcIjmopw1aKiUWcmBB2+vmCKPisXYP1xishMK5nrLzynXAqQEOylG
6Ebcz3rwnOyKpsEOYCXRf5ncoCUBaeay+C1BC2K0x2hjndzodbVe5WZZ3CAlScsY
SGeM2lViChT5AdR+ayFjYvJ9gbxVYs+FZ2oH6BD3Qirva7xdQ7ALXW6tHvYPl/AC
Mto81ODkvE62IyWHZZGtPK2DgmPZNGnpcxKx3aLxkiP85wBOaOCTewCKfwzEJOg2
OWyh4vcYpjAAy5C7I8mZc2mSPkhfXOgG+vtft6u6A24JzidglMTs7j3deDunOr/p
LEYHnzmcH0/leLhfYOkkQW+fK9U8L/LeZv6Kf2MU61vRX4dpilgJz6KpSWFazT7q
AGjvrRd8IQQB9gYT+QU1uwcFwgXr+u6uxrxqlXbs9eJy/QydCPGN9kFmgw6ooC/s
vka+BAX1gplYcH0OK+e1AoORoXvd2R/2XU0xcZKTEc4Mxf/4Ni0rJf9QMHxPWqNz
dIIv+6ycmn1xjIOVyJti7jlu//O2AdR+ruSkQ6htVRk4BbJW9mfBvMcAvIcZDd5Z
EZ405VhoCWtEpq4jCZh0GtjHbB4fl6/W2U+vORC3399GJj5hpPmqHtjT8/AhPc+f
zb2EldG0m5RTt99by5+Rzmt++du8eROy5Sa4BB/SBF+2Ret1a9I4ZcX1+Pnc3A6j
d9NY4Kp8LyejpH8GlnRxGgw6GEzig1Vga2mXt9XG+d2Dxd/+c4XcHlQasjKpDww1
mKf8eN1z9Kxyo8mY/cL2VVwv92q+y0bsRfo3QTe6ZEtD53qnzK+/McA7eBfgPwrP
VRZkPgaZ0w4YkSgv5kxHmr72xhTJKr4RpcQHS1clbT4Q4EE5d382iFj2ovgCbbMs
Z1zJx3q6ZyaSIavCtIUSyhYJorXaL7TUO6EQ9lmk90KO8PiUX6vml3lgZIN8v7aH
yMXzD3pHB/mTeexL/mGHqrgylV97oTnX6H47dsb7WlPVc3r6byKSA/3KBDj8RdAf
w3RRRjUU1QdWwFQoj2GFrAW3LQUDtozjzVHdNvHd7I6/mJn74oDJRMYbq0x5NCKg
lKmsYjihICj4K/fwxIdTsVsr6KdpWmz8HtrHzqJQxFWZnt+ZEkgjpIrwyTm9HX8j
76VlSBSpqzz0vS2yVcmsDz5AWshX9k7MAwbLOVfjKViyIJ9fM/QGE6DKTl3s2diI
i3nEcCL0onivd8FUyamVfrXlI423by+XSSFge1xwxcFp8xuTpOKmDguFHCZy5bUV
fo7bPWcMiWzO2v9Nj9ibzJXM8saXFfIDQ/GqqgfHxLTh1glG7Nm5aCWipInJamPQ
725LKkHaMYiKdI4n1dlalBemqBm1YCXZje9J7IM3zu5tEHiXBYzGCbvINfHCuQ1x
w8JtBOzKn87fmTjoxAhdI38x/GdUWvhrk8f5kPYfIj5cUDTWSVlLijAAgF7jmJ79
iCYfVioGeZkTIOpC4YYpGXGQ5XYN4nKyqt8b4S0ZZn0rPgeOQ4zqSjZw9QIe0M2y
zm0lJl/May3CZoriP4XRDSwmArDY/AjMm8oZ35QkLy7zhdMFvmRYybOdQd+1arPG
a/s2M21N0MmmszNMNYuP2f+3wnImTHT4hmCb2C/wmZkYBPbr/HUBaWuRDGVZQKwP
eGWhlh2XqFE2FPbJUlfGxZ8Odla+1t7K/VtCD4JaPRVg3fTnyFjfkMP0mDr61otC
3aiVTSyCnt2xNZWcqP8byLS4oJpNzqQba+fteDf1MON1DPfqfZ0OhOZIfZIKqjOy
DMj1UU9DIutmWCuVpzmAVq7P9zi3VJuZULrh+QESGXxWh8wTn99mwGPysi/qACbc
VgwvmTgJyo1ecgqjmhBFvPyDtZFBl5VYXIz8k+2Q6RhWj9zRgfVROwYSOWPsBjvV
Ur5PcxF//1BzFwX6pBI867FV570uo66W0MbNjxrCeDJ9oj34YiYWCSk3MK7TjIGS
FGn3fyaoFzyR2UquhpZ36VsuFn+SmVVI54/CBBgGFk0vFS2y1/tzbcfi21NYvMaV
YH8S7gvUgPsiOT6BV50oQBucptwnAiQIIIOfLUvexGAIiGFgKYkJs0i9i2ntzmDF
QRgiKDt9FtGOJ7LQB1+pS0VfINeNFT6VA5+Gk9zinInq0kHnbeg5x6OCFlpzAbTm
JfBYRTwNL3ulx2jFFd/RY5KlqaGGSETf80rmu7Ge8KrVaY5TxHCd1mXBiGezXHrk
FoK24Mu3Ds/8em6qv5FW2rJ5HTtVvzsHfAxFfJ0jSEdKRvbcZt95YQ3UheQ3lYY+
K1IopHYOYdxRoZPqwbm97pwdQHhGCx7LnbtqflvYXb2fd7BvT6qV9Zm0xvTAczHK
C8/K9fmZgANS03l6I7BisDbp3tgRxgMUsHw1/0XddIEkamGXV9RJLwmR+RUj3Z7q
KOmBsi5MQ4v0Gxvmddaebexi5NYLEIMQaVVEInYy2Of4ncePXzHo+t7zb/XWbClH
VQ9bwFp8jD7RcK+TRuj+QOGbAGVcRCLKkJ5FiQjZpw4zAXiY4tunvYCIB0unuYDt
wn85c1TNBrIQqUXBVzggfMqPY7CXtNYRyjkATC8aZ8f82bhIe7hUHzmGsCuur24d
wO616rNOuWk8CwrplK3yFq16wbuu/6HFali39N8oVjpYH2/6AewuPxfocQqj1wPx
sHLTx/AfVnOTxEfUR4QlEECpvjAuH4rNPNlWJaV6ITbEyQ00pOFgL7SFxD8op90Y
4t2J2mr/lsH/kVqrwdr9iEbz1D/dOVrVJe/XOztBPg1+2sRtkBfDMP7QMI3CIB2C
5W2XilC4zzeXGHPs8U4sD9DcRPeQoIApff0Rh8N/V2xA93t5MGOBX0gI3WhB9PUC
PCJCVm7yjIdYW0S5zhX40URyUQ8tv1k0dYGIN3BZUFq1n8eFAFbuUioVMEn39gIT
kGAAhGrI0xO7RQWkAyuiCBgFPROsgPbyGwHcorDgmuTcKYmWqpuXnUTiqTL5ssBL
IMlK22ss7wuEEBgz5KQwU6+LrwBUjTEXJzR33RwgJq+ZGS/UI8FZz7cSJpHiNyOj
PBvfQWgDPEu6Qd3B6kiHq0onWtDQWeXS53Z5xesjTUX0L2W4eaAUvyjcXPSYpJCo
OPHr4/Ptu+UND27yHVGx8fL4dOt4FHo6WiyclCxisotI+W8syfny4SSRHkQmiHZw
N/jUOthnYpVaItUlIv1DzMT29Qo5UoLWfqzlEQ0qLN8PQNBdJZitQ0e+1qMwf6sl
HNEBydGBIehSSeRhYNzzUUhHNFHS/T+Kt59JpcHeFgPmvGjB9WOXfhNtAsxi6sVH
rC/1qAyofjgE43jIuR4DhqIJMEfarnZIaYFbl/MAm89nlrGqnfle3o7YYfPFRqoJ
bK9oLugsLrkfWTt4G4i27ZBfEgJ7hqvMm0FNBa+lkCy62ISEZGdvhC2Cw2Q+8kH9
JHZ2ZW/3ZS9LDrZjiEwXz8fOw1M84WE8hDpuTjrHPsnQVUdY8EWxW+hlbIuFYYYg
wzXtPsNxc8ts4aoeA86wCAs0IVPSYj8P7O1FW8pibAQS1qRm4xurZEMD6QJIPiMU
RyC7mIEk5RYnSt2VuBbvJv/ohpIa2exHCJblN40XEsNgs1kgaSJWyT16u4PE5XUY
uB7iYO9+KzwPy0IwSBQtiQK4AgKKu0q2B4xB36zcRQ2Xxdpd+6qeyQitornHRzar
sQNIt4A7C4ZXhy2J/BV0HnGo0WBSJ0528BTURoY8YH2vSoMGgoZSX3RM2gzGNTAg
7EscfR0OC+Tr+8v+GRrrBKIV2RaVUTZBHlZ2JDdfZIS5WcwHeZVEgzza3/HI2Pv5
N3pSdU0M6QT+5aXrV90wWu94cBozigLPFSvGQ2a9+8YLfkmrBKOAQxY15IHnCSuf
lSCkVym3P88/TDXJ813zqSLyrJNP3sH4ER9kexm5vQ5V2qMmX+8v/E1PJieVnIqE
1cxXJnwWoYO/JyhIHxIh8IMUxK0YupGQjIb46ApyPfolluL2KKqW1XYr9xK4GmiK
5fusfg78jwhKZnQFhY8cOYSsopmPdhh2qiJARvvhbGmMiQn+mE7nMrRm9RRrPKhk
YzwcpwKn6dgEO8Q3sNJ/IhUMI9W/Q/m5Capu+Mm+7/rDV7KvDCnkRQEcR4A3uRtO
2o1RWutqgwkIMCEILtAa2n5128LjfTZSFyi3gG8K+EdjWp+yndSd/qj4mnJEsH4C
YRpRcRompc+hQ1Px8XqpTNNiBuUZbneu7RHrF0KngJRwHyySmBpk9aHSbj6Cklsl
SvpI7IsM6D34xgy/hBgg/rOoV7fsZcpoHxcGpCPrePxHdjNCvhWbkjPTcJE3kgWt
cwaoymqeG/l8kqy3t6AcDy52++N0JaoPCK+N3IoBYQ95xCu/VhYmEjiEurZQFxeM
u408lGHJVef+dq0ueeM5fEGhV6/8MJIO7tAWBKB014VfLAUnWXZfMkWwZ/I4SXHR
FWdjxuzQ82sAk44brvLbjoH+GFfEwMbAreURVLZRLnGeQKSMFWB4ApxdDjZlbVVp
jOjOHQHvlZRuezqmAyd/AIW5Rd28cMUR5PKAqs9S6b+Gw8Su2gZ6J8GBpPRiPTxz
9S8I49QAXCwe75WaNlBjZt9FZ5YsloL0bzImPN+Wat7nu21sqOelrjX3bjS51Kuw
Mnu3MLorXEg+qphQ/QNZBBq36FR88h4oq4ZixWzMf1faq0aE9gyiH5Xh7BXLFSlQ
Rj+ITDj+vd7ILwgKoC/uJGC8GXuF5sOWr6Ux+VIII6wD9rUNEwTK65wI5lZBIyMZ
muL5iX8s+nTcFkwcNzPeWlLtryvprQxdpiY45xfygYIOdgHWx54g0ITB7Z7m/lxF
V3V/a2WGtw1Sst3Xr29R2g3c8Lvx9e/KFySUxbbAZ66rhjlcVARp39upSt5lnr+x
WgCyd9gQoMixKVletDI8aR0VMzmECan1alfbg3tC17Lhx75jv3eUfbW00ezSPmZZ
aRQBR6QmiVuaKSQpHbqvR5ODsWGCAjDANnIw9AYBNM8YOYgvRbWbMaKSHSmuEjt7
AXHTpDwg1LrkGsPYSx1hYTbKr2A0jgvciAD1FN5hkNE/UThnHyLxZGaTH+q5YXST
+YZy+SdAu5Ln5YyF/rOoXBDfvVDMAjRR0EnX9ygV1W/ERmreMrwAZuOLDTu/04BS
lv8qQOUlXDHhlu12DOrTKVntOJnpHkv+PskeVFzSEDeDEq4RcdKtc8W3ZjOxgmi4
nHbxqtORY/c/iUEx0zOwg2UZ7KUDF0Wq+3LqfQX2DQaD/K5X8JzsqdcEBvvuBnMh
RbcdbC1ktDKz5w33JONbmiYEDJnoTnYnLN1UdRWgoVkGG/sOzwRpujWj4rWN12+B
GZnASNhdeP/wyFkMmGd+eniFDCSoOj6YNDbNDmkR46VjWElBGYReCnqwdN5v74Gu
Osgz/RXoLuBQlzGYGdd1pcY3kIbxOGV5ZaZ1fttI7b3NewVZiWFqqjsI5ha0bMol
EDs+XLnRFC911TbJZN5l5Nyv2O46/imYuYqBcEVOS26Uk/H9Ne0IpfP2wr5sae/y
u13Zcmlj0oO7MROjXnNXjQ4d74PEPnCA58Vb7rwz2+lJoJszp9IwflL4kGhLrQ//
dsAkeCtuh0BZ5wf5nDL/v9vdl6tlXz3m9sdYNDby0+wmni8yUymsMBH/G+PIZVzL
byRExvWle8L0n/FcZezmGkLVIJqKa4uLg6QTjkSjoh4JMGpqaIWj5FPIiKogGcMK
5K66Tarcq+TgdPdnLCV4DCwn+CwCLZ+galLUJiHBGDTGwk3B6GQ1hph7WixqZTb0
WWG+tCZSxpLSPLHQjNGOaaBwRT5Nv5nFCxSeE+bdB4EucumDQn87kVR+E5KEVnR/
2ZNsPyuSRLAj21jmn2d0tXYeVShgT213BN5WUf0CWX90Gjh+dsJGXovGDfnv8jiN
AES5QYoLIQ3Bwag/C+nPfm2UNOnfrcSVr9jStVkRcd3DhtqfdbOCzCR3vpT35dEX
Gfr93NsVwyvuahkL+srcyaMY/wIMwR7G8ibqUvN+JJ8SZl06AUIGOT3m+1u5Viy5
PvxYHMnYqkw/7NJiCSzknszWWZwwXDl7njXsK6li4FJl5178h5gNORgvGxXDU18V
mFTrKCrsQFsSvuCY/Dnav9aPO0B8xr/IEwGF6s19LhqwYmAHjaAvQMH+RTPmEYhh
NdqHLSq4+0xJ2mJ8N4AgDI2Z2mV3umUth9D3J14WIbdb9G9ZPp8x3/IH5Bp7KcL0
q8PBV+9seZpNBvKb0IuofhiKkChoKd0LtB5uRf7tMTwCEtZeX0R835yWzOiCOU3p
SwQETB4NhslkmY4fnfHYCFkDEhgYrYDC2DQLdb2qA5ypBO129Hi2Tm++sEoD7EcI
katA89wduC5ik24xEfhG9OAXW3pqXiYs7A47qkH56oAJD8fqTRuQls+AQdBHdjih
sMmdx9C7v7o1Kn59TqXNeicuTCFf7JpDrepuVHOCWx+o9Mma4Pr9IcXydDB2UBZ4
CZ0ei7XnSI83JhUTCYrLcQJe3NpVBiVvNnPi9tATwe9FQj2NB11jx028PlycAP5U
TWN/0fJu7UvrRk4Iqp7WB9Lp/3GXZHAaHc/P2jmYT9MXuemtsdwIybpcWNfM5Eo6
PjhFXg0o7UvKV/066mw8MItn//2EfX/i98XaxRi7GCNeZwTZpmOzqdQTRkYZJw/m
Y2hxHWPUf35ZPMsm7XW/3S9X26NgbfVNPf8ErNGHw6TYL7e0lpkgzIshCOHrON/y
rcuDEQmte+S5EdLXr/rWLpVCXPnBmwGm+4ULy8ujKqquW/ukB8aFmc5ZZ5xgsGln
IRdewiyMsW/lTX76AswwwkyMs/viLpbi3gw3JtfArDoDgVxnewjd2n0FQT32Zd+H
MX30v/4ZbmDnHOj8v0rvxdCf2yJDAJXhERipA8GhVCyFe2LkVMJjYxrhD0+BzK8c
MhjUfPUd88Jq7Cesxpoci6qb6tZUIyKhNENhpuzb95LS9xXBVM+EWlAsd8ZXp/vq
hp1M0iYLUXHcpcoToPq+NkbUAE09TdWo7wSYxqSwnc2ew76ZsYnJLHGsSxTGLBG5
+rPBg156pHIDNHs0SAZSy7ZCMRh+qc976nbQT1o/nT+QG5JX2ll9DnjNjvOmEb4A
ji2GKT5J4M4v9Ft+fnz3t8w8+reTYLwlPDClIwLmS2Lc77z1nDc/YN6mCLQawWkc
vhL72RiVSGQ7WnHtxaOGCtNdCddkUI4H45RX6hxUpIPCDu8RQiXgvv8VzXsQnPOT
Vp+5jwGcNQpeaO9Wgp0kTsZ/7QPGejtu/tS9tW8E0J0U+BD2kkohjFpwjUf3o8J1
z3CJMOr24jI76HAydvl+Rz82/n1fdLvMQlgFHzhgA423Ya6CzPHeMc+IDlSNz5sw
PukaS29QbCXxfrOws0BkqHyINa1Ho+7J2Sw3DZcx4zFsH5NBp4jVUj0v15a0sD8Y
yyC1M1IZqhmwb5YTY9Xm05whgLHfGFKIIY3CG3USK+mITsyhTff9LclTqHfruGD+
Q6uRpIv0F7XNUM1Thzj7stCg0DAHpeXWeGUFFdZgB1XnHerunLRBcbKwvp78ze9F
dUgzpr0ogzYEjEqH6ZL5q64LC6x+YPmk0Z6bB7xYu6k2BsFH65X7pjgO2Mhd0TuV
3WsJMBs3lwBtm9spotOAG+bhxAbWAlvyh2Oetpmp6eZuXMlaqE1xoy9ojpCCAwTz
8GlfoTwvPGi0opruP86DcuG36xkW/EZKKJilOEcXb6sOwaAd0RSlR4jB1SZiOBft
WzxKIXgbSqoFg1LefIJIsKdtgGh7cyxhZK0A99pFRpYnOp0f2si7k43N/X653+fR
h1B9WBDVZxD4fb2Od59NmZMR38FWuAVw4XB2f6LqEMYikGxtalpaIJJm6LvuBZRR
6AZLJ0eWgjxqI0YqAngFr/po1rDBGhKF3dL+d8O5vYDs2DaIPOzrAs7Zu3jwLrz1
pk/tbfDXZ+zgv+NHzsrTWaSM+Q+TsYUlF8oBPDiChIy9JY+UFyRQDE81qPDuL/ye
E/wPayyrzO2xE31BEfp4lhBKCocbudC2nIAiTeJZPL2GrKfE65FArcxv2FjP/j96
fYAjJyTbdVcMCu5dKr4etehwk1wTzS3BwQb1dq/LU7p+aiUE5TqIVyqVJSNRy+Ms
A/27XeW/ecMfUhE41+N1AkIlskJuVMI/LkniqN1iKBZDzMLMjIt4jTcjhrNTI3Fy
uqXV9RIrqQ4ekLPee3L7WmKUysOrEwa1xCHOk1bD+BAi4baLz6dKYbGkp6C7QeKs
mQpC5hrno0m7DRMUSyUp/I3gGPT6Ju2L6PqepMfhQpvjLzekitN4b9ALqhymuJfE
JcXUMBxb8AHcs7Jro7orh95ZfqePuSNhxrVlH0oMG7Q2ajxieNBqQD1JHxYeNuve
Juy+Jyqo5pKnbnkZEwJN10NZuSPXwdVpOfNwh9jNj/Ase/4b2LjAMLRjl3Pj53yD
pVovFhb/+IG8BCOXFrGB1KG3Z3//cqbxGer26hmOpq6UMpOVDHjo+H9/SgVdHOrf
Z5C9AeC35f5nfupn1e4VTHYWIFt7dntjPdbK4GCZijIJPL00PNZuOHtVgBbGVp6q
3at8ETT1przLjqamHKSDeE2GMrXz5iyMSq3X2N1/lLCzefPd8EvPYgMREnFpZ37M
QQKejpePF641bu2dnEvBXDaUFf6dznXSaBFRN3+u2aZpJZF3vssQKcbzoKwqM2Tz
yWFviIVXW32VWclMXR2amgAQwR+0kGSI9T4Yfg9/Hm9atFJOJA4AhXZD2seiVsnW
Vl8xv5mK+25NZvJUZr9HOrqTUExYBc0AOvZYfWbZQAD0hbAMquM8faEJluFsYody
cfyrqcw9dL5Yy6I0nSjYQp4jsfNOmq3Lpe9sbvrizQHe7H6kcSld6EihznBSzAEe
sy0AsVfTagKhIFd+HcPcZxOO0ZJSzq8oHibx+pHTnfZ/Cq5rcNQY6pITBmGBPpdG
3moqhtsxX6yer94orKyn8CLxIs8WGzNxQErq4x2nkRBdGpDzav8Q4WnaxgIqQJIt
15cB6mKpdvRhzCeEPdcFS6vcbpMSyvVbG1KGfGAuxDsIex+rcIZDKB6QGNil3NXw
lQgPO+7ezG3BonkvehPvSaUuWzX0uThP/1qWEmw6VYH3eRlwmEDnfnLZfXDbUN2D
C1+0qwcDskCh5G0BT9VCM8DQk1HkCVYa+r8EtF/CiA2tNeZOtok5188txRE7mA9h
hFiJoJyuT2lG3jdr6adwkhhFMoATmakKxS08DmtFhUR9fJ22mNy5ym15ZTQjoo6I
6gUSqbOa7LoNNrNh+QfJEpdpuP3qGBcBf4eq4G/hfmv7pC9XAgRhWkyfzsbmTz7d
1tSRuzy/hJ6m69I2d3xCcnUcCQAoZlvKA3m1GeR3PfOPYoVDQOlKAp5RXZ+u2Rf7
7KBh92J5VYkBkX2zm9FlksgmMKwZNmuk/LC0cKJYk5q5b8LM3RR9iygLonDC00ML
hmeKaBm1Fc3TlbfIV6vDx8qJ2zFk3QsN+sQ0+DWM/Ec7CP1CF1aLPIuBwBQBUqiz
NlzNUqaqB0qi/IcST4HihTfBasJej61xEh/34ULFys32R0heWQyk5BITs5V4H1n5
f55e3cEiARej0RItqTL+n1sW4/RXm4vgrEZ5DDFGQOy0imTYRZx5UjjYUeJricH4
R+6i0tCg0hUhMlkfy/WGA8CxqJYV2iEwqw3pXCQKLMh4Ku0bIdveoaIlWT6qKT7J
fNVT2p9CBsjN4OGZZd274IdvM7hkhh2mxrfWZZ8llyqt8ofJobmPsMIYa0ycxgi0
uNm4jztH/s97thuQLVuGrreaHA461qFTbABWBRDBsE1hvowk54uzwuMS7oi0VFsy
otVLDGY/At39iBqjw6euCnjGAx18p2RBec3I6A9VFOB0lGc7WTjRtuezACrjNAIC
+OtaZfFCd6YNy+FGHXyMYEG1ITie71kypaswt6fjg7dprP3brP+5eUzqWxrVmFBS
6E81oS4P9j506F937nuXlBQTgtXvrLOkE+ac6zPyhh6l+qBD/gqH0M9qYqPwl146
LdnF9XO65lP/qqLg00atjz6PGW4SvAX4RHSHmQsT8dKobad92yKH0gnGC0zRhAc1
LZoYDGwtmSHlNgjnJQALMyA3MU3ucH1w6kAbosIduKFLNbzFi5CjmhSihIF2zLeS
UcL7d4xlnVNqegBWD8bIMRzNFYg9IokQy1V+Va/JVkzyMc7A5Km0+r+2TeBWS42v
goCgdgdAtN68srivBxpSHSdj137VIPfrCgdZQuXtwKgJ010sL+sEtR71nSoSrGht
OFycNOpyoqCSyB2KDmrPhr0yN4tCY4tyCLDHiFmhIHbM/cC4a1nsK14Eq9cIXx2j
dXharbfH8KyLej0lNhgbR7hnk4Mb1jTSb0jYNVLoo1MS0zrCKfkuvCS2UBEUIQaN
O4SbMgymH113aNSxYQVQxb49ex6KsZaOl+5kKeemHaSDmkXQpdXS0qNPcG7vFAN+
Na+wiTGU/3ueFfJWtG78Qf76ZNnWAzpYIHhTN/Bxl1SA5dy47razgc/UWZXMpEvB
P8MgaWf41r394C58W+jjGU6n96d5dw3sBHBNz3tqpdbHe06dFwQZQtGN/KHsSuTZ
Cyy0vkydhJJDd4n/gBx9nc1mhUhycnjBuD5m5OcTkVBrGaU43ujNKcxzU9OMXz/N
60juIpFY8nLyvZcCqrMEt7j2Svm+M2e6qxAQe4T7utWbMi2kDEkmGXvFG10g/uEF
Fu+8U7eCowSUzynuEoDiVYmcN83sCHka0dnxTNnTYnImUT6u+Vp38K2rLlF71Cvd
Pxje8KZBIVSwk7HwWmTBVT3NnD1GmcbwAAM8KSG8Cmvo656Q2G3bkOhVaAZGlCQH
64R8Remk0zutvMVi5j/5MwtiHzBfWROnmWhCD/jomQLhCNz/jPsY/qDbqJLCrn7q
S7VO/kwZRp4XyFv9zLymRVgxKGQdQ7dMYSJ8MxTsk/+mlkZusf0QO8dASt6xU8CP
kFgwQvJFcvxow129u/olJyj7gx9yHYM3D0ERphWAROy0rFM+4E6OVK7IPkxGOUtZ
j02TZfwPhsocj3PfdPllog8ZcT+km6/byXwSxEWvHcOkRJs1zh8alukABJ71P2Pu
U6ximtcGLdBBmrVXgWizQHqYrM5ZeIxpxTzjsIL6VtQXsTMZmPxDpM0HSEsjMms2
i+z+5XBorAnAtcnM+jY3qwVG+PrVffHpNjAX1fUm1nqwqvbyAtVBzuBZvOLRkMor
2yf373VrS3pE+wDYWAfHnN1FJao1B5LkhWGsemRyNwoXeo7GsAN2IESscIJFwL7u
cter7/cvDFZyX32UuOhdGmGzcu2EADCX6Z9JQf4aVQNBqV6EwYMKwl7Y/97w/zU2
6Xfv1GWn+FvClG58tCKSoK6ErAvICstdTzdhjrsIdxU0UfKCqJ8/+4Mf+juhPeZ4
Zqsi6PQJ7kbz1A/H/WlxygSufbh48fWTzzrqWOpIms7RvMQOc50OjVWtRj/1A9uK
DyTOnxDELofcNlQdUVdorc75k7NddKAXzCxPOgbOYkjuEkNnC0efHgNhAjwob2Lz
7GsPNik/+BcCzzc2fTLW5vTone6N3SFeQap9YUD34fQx98ASN5qEyqfTtB7b/hI4
xWDHXe3xF0Gj+/DYa4Y2zByoz8yVVNWJ3khQHtPrinBlB67LDkCQkCj0RllQIjNl
VtPBwQtVhm1aCP0PyqhD5lIPmBM2CBrMeWTdUpWgBLCV43dpm3ji1eKP1gs5j6Vn
jkNik78TbB/dAxYL6S3O50iNOg/PhYv72cgm18G4PURkDmW5F/7rR6ye3EJRwwqu
KK3TcudJxdzsYRkcxWhP0MyviMxEP1rwKuRtcfTHd9D7wH3Dkm1FOZ7tCtFesFuJ
CDUFeXy+pOcgnK8BrHu5Kqf7lB42llpZYagx8qin8GfptFmMjxZd3nJfd+NLXM2O
aPeUxw47fCy1mbe4aJQZ00tMfC1VTMYEMWStcAyAixBqZkTERw+xV3nxmFAN4b7F
u3h8kGBsjyGPUa8At4fMag1mrtQulqoCpU0EEJzGKVvnRgBMaV4zPru4oqPrg2bB
ZA6ItV2dbeyrpJkNGwr2qUAamEa1tf8PS/NYCYbERPe6itYt4dqYdRBPBAZs/Qf5
Uc55IJw4waRE8Iif8pAPvxu6API2kmUmym5Bay12MOwKpVmRAaD8QhhMMNjc3FwL
biYYsA4hfQLwD7dJcQUVRtWv4vkyY35f6J9MP7hqoUf3Uckx6oBIw8XjYHwadgxp
VWedduhKMl3dlB+edrYcxCt8VFGlFuzt8js6VfxmVODvxg2k9JfFT0vNac2GzOdw
XawHFIvSnpYZ8g0A5Gv3abBaH8Hmqk0LRGFPCIv4WoYJYGSc6K29EClrjC3wYf73
Sc8ovWOe9/wiZeOb1YeD8p5xxm15rM8wKaZfH9LGs8j+damMsuOyR3ny36yCgOWn
sYs5wgtNN1bpLQF09PVBhZqeppfIAykNmDKPZkOPkHyeEuN1jR+p4VRQJe1VEngy
Dn18/OpA4/Rmllrd4w65KgyZKtWxzSRDYd7dRxfNOwXNvpzYzamPvMxnYnrsIO+s
zX74LMSLKjKC5JgwCkfyfh2hjI9mpQ4X5YGQj+kyDhok7F9MlUBGBql7pvYW/nCH
tVy6q0NY9O5yo/RHRpPKoVj4rPvBTFek+iDBkKeN8R1Vxbsos+xNcpxLin9pozx3
b/lfion/CIv88qs66dTFAIpEXu6JNd8AlFiZoENB/hmexHxgE/D4Oxgm7JvcJ8y1
w6LREp4W7hYFlb+PTDrGV1N0aU4pO+QU3FErcvOkcReEj1U/hqLf8appfz/zheG4
S2tuy98KTyRNWOBWEdwwjlTqeBievPdloqczmojOAoWBPeZ8f5Jai7gl4ZvqoRnO
6sT3SltyJnjUh0KmPCacg2QWHpUM0rIYmzPyS612NbNPHuB5HrBGjWCnztWq2TYk
HkTJkSiZEf7WIwxDj+Jlex9t3/YBcfqMhIPkwX22Kn0MvcmpmQemh5Z+QAKtS6Bl
ue2vHa39WXvKzWspxnjAAwndL0VGX5fHX5jzn8DfpsOYZ2M3raKqs8xIvxVPmVgw
4Hz8X1kJLqs06rKns7qPTsd+hqH+ISQ8PG3Me3raQhslctQgvyix0lwv9Kf9Q3TK
drUmqX1/Yh4SvcUoo1rcOdjJ8kuklNpP2+GDFhkxlr/UvVcN4Kq7mLE62qLwXRbJ
nFNFzsu87FE/O0ON1nPNk2eMyvy246LYfUTpl3FlTT4G069jRiA1+sGLB7o8EW5i
WUgUipZ6i+Jl4cPEZkz0REkODIwjIIAw9Eosz35e7Se17TLEU4cZWWJeYiSGfuTW
9pIxUs7aZh8f/ZLaObGVO4l8rR6rS9QZXUc6LruXw6KZW9tYojgPlpWYnkEybiLM
nQd1AR2MoKEKnU4WMHtX4RWYLfXcK2mAzh0+Ubn62S/FEAf3Vee3Jz5EMiCkjG6I
ob9k+MAB0EhbzcU0Ixg2ZmIDp6BPo0YYN96Wn6CJ5Y4lq9w/9a04QONdd9Y6XAXl
cnAFO7Xyx2QQTyngZyffk6ooqX6omr8bXzsLCS2aru//lXq/nWXY0aXdvExIe/jK
FBi0FHheV2U+2cBla88lUCAzQIaBZbdZRELKyBR3iADrIFaRYrp07f7bbQp/qllo
FTKzjwBfvogzveQfygem8Q7+QvkQV0jyxNMvkpWSqsGoSV8hwLnusiIVmnqHGTin
TiIcOu0UhIpayVD2hfVS9Osf+/Vjs3Lz3fWmE6hEeZiseh9o4kJlxK4h8QdZP2LX
Tj2DE293XcBCyLwcaWIXhYDMzkhfr8I1cZJ1WQ4yVk7td7i5cvOFeOVJOmeCJP9x
RbyGWduhbduDQ8mMCOuLI4+F9WYEAzze+kDgi7wvaT3ClF85YKHI3OIiTSc8WFDS
fpJf9QmaXmQB+CCD7uhmRf4B+breh77wzXgC3eT2f3u1ouwrBA2JXqjbivYOq4L7
ksWwRKQZKItuvrVZVl04eWF23u/g5kr7WSEShp6jPgJfQr7dCf2GTHvxdptbnFLE
d10JYBZ/Ifv07U5TTGBMm1yjcHgqu0wO8/1kRVX0k2lwmC//WPgw8+vWHju3YNeF
vc7+EoYtFhus5KSHc5WYJFej9mFtRSSGJRr1+c+Jc+Asow+ABqRk523EAxMCV0EV
KtL7K75zoK1fSsGpqajsFLsa42dHBLSFZT2ZoTGpiDLcyt0QoiyDiY6glkxEruRY
nyExoHDnKsK3OxidmTzalxrv/dB/j5CImUYpMhS/JmpsjHZPl6SZSnBWwstsl0E9
e7dhkZnoxMxNYhs/4Eh1/m7xH+cXfkZ8dxhqjVkC11w9ia5OG3Bk1/GgqJ7v+HIs
9f/FN9QtqgAapo3noJQkH5bfLFVDRTGmZjHvzuo8eKZrDeBoh6UbRjKwStVMEbIw
h9MW6LvZSijmCkQdpEaQdXNaeTUK6ZZHcYl9rO51NtykEh4se9cDDsUs9Ja2Vbje
H5eRkIcxRiO/WAGeSilwzKdNd7VwjHcO2qlh8PDcQCdaVr7gRyfpMYylK4LZMjJL
tCsK9t20KpavlHR/rZYvVBvOzf5fFZXwSh6njCIDw9bCrftCIcJ33OFgp5XOvsaW
xexb6HuaGPYPTMRFOjRD438JbhAvlsA16froAjapxVAYrPtU7767fE21TpPK/REU
pXBr8ExZmaJmobKgKPKO0Z6ft1TSzHegB4lz6FKdFfAn9bTj7pVwFxft6H86lVBA
77c4SiPgx2m7m9r557Yf28wKu9G+CpttKjpYaVM07jm2yaB48bil96TIkowDKAP0
6sfndAiM7S4C9Jf+9oAJQsCWuyCeyFQ1o8untsEhQP4oYiY4yE4pPD61xDcir/7r
aJ6svv3/mtqVRW0xthF7Tdp1ixa6gSv1CjKtp9CIwJrY+3zTVUaxbbTH3y1zq0UJ
HK2PaO432QMKTAmYTLgFD489BJFH6/oE8o6Lvf3+4b/uF3TQ3/SYVFu1WMTYJAsh
Kr/muSAKxQoeeokE4emQQLSpwXiW47RkAPrhwEB+iT4KlxvGkEFkgB8TwhW1pGtI
BOx3ye9E1lmFnA/uD3zSRfnRd8ON/+KwaMIgEJ2AR/elqR7jwDXhQV3X6dUqgGVv
5JVPtg9zyamlLe3YX32PYKioaKPGkhmUMFXdY8FhYtB7N7KYc7Wmttdc/8gZR4Oe
G/7nH1glMvEtbZ8VSqkzT+Rz32IpRE7fCKJezzeaeRcNz/BiYf12otx8u99B+X6R
ynYxFKIFaiM/GkNKav1vwfFoh0IcLrdGd+cI/thREqXpm63jGZupUgO4SuJyVhPi
BT+v8y2p63iKsAQCn1D2mLba0kFH9tvebknuoPLJ0dk6Ea0lKJIfgbDzDfM4Nodn
277DkLHGoiwEd1f2wQmGoCKYR+SsMriY/tV9V3jc74fNLX+snolwS92/IcOweR62
G8ugehGAex5AGNBlWZ9Onsbv9vRn7gMgtDWhEdrxavotdI41fYisQi+jX0lhTLcQ
nxxy6afAJSvihmf/I6uLDGp3+c7J9HrKg3ZVnA5vNL1tpthRFwFDZ08Nr8mosPmx
iZXNLn1/eafjps9PKvF2Mvb4KKyG6c+MAfH06wkapho5kL32JFl6GZ6nPoxHQ/8v
N+XCLAKh7A1KnzoRSg6M8aQtsEosEEm/6tW3B1gywv5hjweqQ+i2zfZ96OehTL/l
D8l5voIZ1Nv+LZp0+4byuj3kKs5oMtyqJS6Q1msk66m4w1om4ztBC3al7gYxhCDI
SzDqkM8OpeUsvp5H8SI1zMKsYeN+/mNy5FX2QMYis21DjegrVLqM/W8EHRoQ134H
OoqaL/a0gcq6ZEdrCj5zLc4h7oJ4mw19Y/7nhQHS4T60vrEOc4GgEmzc33kk7Pyg
Fpe5wgRvIDHRRyl6JcDKfJ6vBTzCdP8y9UXMUL3+nVr7YI05kSvmtHFeenBoCssU
gyK8ix471vpT2fD95h8YB/fU9zp1H15g4noodfDVWNrLydXHRvojiUJExST2Dpg9
TNpn/EPJBAdXkpvpYI8tgX/XVD1dme+s4xAYeDnJydL0Xj/SuQ/IEkp+vpZa5Ogx
n/XjL5hXBVkEkKNJiqJmMRAc3fluUiX2q6gOP8p33+9zeGgC+n9mlrElliO0iO0D
G4QjSal8MUq/M45m5L3MP8gNfAbsXuaIeH/KkSmpQ8OkO3ACuUCnEf3/WbCaZ3+u
TRJRrsq2sx3WcAy0PebvDJlVBZ0EshBVIfrlz+T7hbK+FOre5CPzN6avbVVDzCak
iqZgx+dC8UseKDGYiHiSOfgHzVbwnzXi9XNcGYgeNqF1KGwL5gqs2sAf/O0t0tPM
VzWNClKaE30wy3+l5D/xhzOdUx95xan1luHlltC2V0O+38kK9gUX8j3oks5tR4Tq
ZotzkHSAuwlAXh6FrOzho4LpW1Lbqsh1NuzvwfeeaU3Lv+F0sualIxvfsuQR1siX
JXn7Kc5lEIGlfqCsF4ItgyNX6psxi76Ow2FfnNS4epWDet6NRXcnSsGQO+l8DTW2
wsfG1rPXhlucinzvTbPHnD+cwYDzptiEIRJImIWwKaTD+8Eh6/yKFDIlnYKB8Peg
klhlmemH0vQakcaUasOSaixmQC2dXBq/xOR6NR+IZ1gonEFqhPC1vjYoOi69ci4j
PZMCcOw/ZBKhXYg920OJZL+qLiV/wWXw3OrvZhk1v94BrFnkwWvKTcIRUbwY8QT6
Pr9tlvzjnlIS4Vkps7Jr0NMBnb8XgbVqCN8frvOpx1llHZsCuGaSpgUKIUdaEqmZ
i+exMNrkR4I1OOJ7vv1aHSBaMTOTrBSagWfJadNYuaelkN/6YgLTUOMtfcUy6vLj
rSBI44QuUc2nncltOzvQTHRVhOYRXwaB1BKpTpEYMx6HxaPYJplFGr0/7oCqYuol
A33cUcKN0Bb2RaoEhIuQlSgaNIbkId2oRreZ6Qns8ewVFPP2AtSxF4Uu56ePfyGv
L9Z12WXVKRDMKi+vl0EpQnm8TkZqXvi5JRmjIurpD8Z8X4qP2i/+nx7k1jJfRnd1
h5lhbjr/3PcE+BGGyKn52Z05kp2SvIK1HIGt5PuufmEwCkSVCJcIoRgKNrv+LdGU
mm3niymJXF2WTuFQ0GF6n+kQwq66zam6UkSM7YNpRhHGj0aObMQ8vLGkxkxh+o2k
2uE0C0G8L90ryVK2yl2OHMFvA+7Z7fHxMKipCgTsFSxYrhyxdMNy8rA/ZKYiPoRb
Bs+HKfj579AL5ItcC+DQsCSW7bDqxDTTguSeX8AiJ9VmF0D6HG5BCUH7kNwiLV+i
ti7DNTw1ZiPBjQd3npMxNCJNZqK6fGpbIwguBTurAmZmgkO714an1pAHR/41/1hL
ovy1Y5PKzQQUKSHArCrYYei40fMxf8nsaU0mvS6SUetFAc+mSsJoAy+AMPfv9nHf
/+6AOiuNkrqaYMkd+UGfv/CHdFam1ZkEpulxs6Ja/T80YfCOnICKQhlX+QpN+TCR
W0nJdlMMv+tTKAKcXKOHcHB6aV0xI8eJzNN+Gd6ljonvh7xxGJV6770pCS1DjRXX
fzFwB04ZcyPzNtj6FDxSm3zH2DsPhBtEaGnWpB7MvU0IvD6k1Va2NpV4EBM8CQD3
Phez6h/sgBA4gUO/zyE+QmkEzskaAEfvaKZH8VUy7sBZxNv4IoIyuB5ZPcI6Rbi0
Bo4phzDzBnwy4keItuQyGY2LRMz1nxsKePcxzhZG31sruMhGVjwXg4mPpVoehsjf
JMhqtz+mtL9xg8o2hjcx3AkSfrAsREs+UbPmxnIy4LIxewX7Ye2DtlbYolyk7tb7
lsQoY5J8JfKDAlenzaZmZDizAQfi7JMOH9mKTG9zYTFsmKECiM0ch5x3LkRXh3l+
HEtH06U8A4LKu7n4GMSr1vMJkF5uFEG7WNQTOi3DcWBG0noRFcUP42OcpVQHUkub
9540O0JxtDs8X/pQkYuqizQ8ipDJ1EzsI1eGrY1Hrzf0XJ6XgnH9bLchLg5vuAPM
g6NRAvgZLw5Qoi2MB6l2rzUNVAfTsT+iSc24zZ0Vo8/WwTw+aTFwXE1WTn/Qyo7W
7SO/tConN3+/rDCGmbP8lTNYo6b73pU5n1XNJBQhuwws3inKQ44Q1iOV1XcXdlFS
42MKTQfgrPOdDRKAD15/pAheLdj9EDQ/JgWXghV1breHmvPhvwExjnr6jhh3OITo
6dNFCEkdO2P24S9FU1/8EDBy9ibequyC9Oy065KxXHXsUS60+sOFB6VjqV85Cwxg
zsoQt+PwV5CuOWLi/+3xqeTOcemBtljcyIDMGBw+uZOoYje+jBkDj1ZjQE9dv8Bc
ssJ4VeyixpSFiGtJeWb9sKSNzRT+rvcx6vMDnhGU7ITWTE/tfIUfLooSM3SDt0zO
y2exmkQmiMQg4U6Pey4dylDVcu2gEiXwlP/InZvAf0YyjuVhgpiVVxqD7DVdMyNh
smw3S1K8rHQu0Vu6gBKVHOHaRFDevEOTPD04WhviDKlaMueli9L96d062RwABOyi
t0HYCdzCgOYPJa/gH4PZBOoikM7GxbPcchCTsxrDqaIHmcq13CGlpBbjQNN6L/XY
ehrCxGmGdEbHP+Vr/Xcp+KagoVxeZL1EB/NcyQh1TSxi0VCY1SHPbgGXIKExVqk0
Gn1fDk+IbLABg1shQ4LZmkKRuOAXuaKBaWV8tRL6EQjHbgsfQPC+EAldRnopsuX4
8QYQgZEOciF3uwbkLAyCCRl84VHxS7/XresoiX2+dzudFKq7TEgqZNpi/UoxzDt4
vVeis2WkXB2cHEVV8Z8O2MwwtgVjaCLWfK2XoyqcQBaE7hLVu8ZxlgV6g5cFo104
3yt2hAgWLQXnDNMkAvu4t3DAuk2Xdiu6JrrIMweS3Yo8nfzfQkctgNPQLy7KswqC
D8jO4JpA6vBvSKzOR6OPStaZRLxQoIDzm3GBlQqC/rIzBFYqy+tvuy8wFX0VjukW
N2+sMemveeJEnRis/L3EfaZWewdkTzKLFbofhYniY+F5L74mNzklbpygk/SEEsWA
GuMZF1k+yYp1FgJqMdv/a0a/dJ6TlN4zMXm/EuRtd9Q9rsfiTHKgKUEpJuJW652N
O9BEIQ23i9sLRTaggeoLEN/0Shl8LxAr2DcCJ+8xd1BArgl/p5YESr6ng/cLZIFl
vuBatRN7fk+7RhTr1KZbuotR9Rycs+U2eqHBzCOp98kt74Q1hhn4KkRHhW45tAHQ
hq1PD1HfFScbHet7Y9TEG9oh75L6lsLMrGKwi3wbeOlPc6K7WNOTY764SdFGTent
wFnAgT7r0rt08KToX5Kk0B+qBwN+dDCuIhJqVlRrUZzdKX9Zejjidg6jiaILXQO2
obr4yWpQtIlAjaSwxoN3uAFRJw1FGgVJZ8ZHyegf/H6mSAEe4OrPnS2z5KGFPm9W
Ddjc8CBammG0XGuwKEx2gA+igofmAMd4XW83AxVLmMWUKI4f5Ra745hqmBZ6P9V2
WDWeogwtg9gjd0twgPZMEZTt69fjLTEGvDEeQAd8PEFVUssh1qYNuj/wIvCY4FGI
zK0Kp0LghEutQpFsj7Axp9fBJHAUfPUi9bFeRkHzaRggbKqAV6rr0BKqp7dQq4Ht
gu8VJtIiWE0fKTSt9VWmNJdu1hP8TsB+41xHTF/L3TWq3qSH/jTHScC1FZffESOj
+CrqZpdTIG2tcM2GrtpWXOPnlurcPkB6WC8CcURI1aUWBe5779N/q/010eU8XCpx
gLdHsLW8tf7y/qb+Vgc82fJkB5ZwaGDTOsiwaNtoW69jjd1s4dLxHrb8tckeYCTZ
AU5HqBatPVmYKuZfqtD7vBZ5k+f09Pb3iGa7r6tUdAta7cqXIMYZKvLZyDnAFdDF
zkMBP0oY+epBOd3Z9NoHgC89ZUfMXZ+F4CdSPBT7UERYNCE7SJ7M2ACpVIyScKIw
0ezFJUZcmFX+uI5FyB9akj7H4hSyKhJR582RNUSjfDqSyLKHvLlxV9S7HJmKPvS+
PYzMGwD0BguvmDnmQ4dWvMsrt51n/91AeyPRpiY7NHnFoV1EqXWiMOLwF3fNB0AP
/sj9POcQP+YJRBAWk6jn8kBKhr5esfj7noc6U1TQa2eOr3gyUG2u/McALayoOD0L
ZSMSl1Jetm1mvrXsTCOTWtQnNSOsDHiAFbnG2iu5s/n0JFZFoYrwJmUSYcpK09kD
fVCpJ1t77J3Ygucka0uPeMpBYeam2NdnK9Z5TDDs0B2PfN6lW+V/+7fqYZW7J8+K
13Oe/Ymfw4DenTZ5G2VJ7BRaN/upt5XefWtDC67PME1jjshm+jfIJ5j4Q9BKuX6d
edZ8Kr3ePgr0q47JwySxh3B1WT+buDMwRpX1SB5pNbDhhzGNH3nDIciXxhbSiBRx
KhJOH0PJNjl3yBDbSkAqQQDTrp/wKBz04U/kWH2YHcADETi3XwnuCJVvpM1C6svu
dhyLeFccIf7nXPAmdfV2eJN6gw32iYBf09yqSLoAduwbF/nnr1TLrND8YxkNvSs5
GfbB28F3Uxa8OT+fAHtbYK2FQBbwTllkXkn/9kLhcaMY4mbXtS07U0eYer8RCR6V
v9KMfyIcGAEaxHf1XzlBdH20Pifbwb+LNPfTZlzLP/BhFUtgGdLIyIMfyeknkJV3
DOqi6XbwaU1UPW0lZsQD7UVb9BhUQ3m4eEmDdv28QdYjgVvm0hRnZ+LGTY+OcMiZ
NEzdUzzXI+vVk1SEu+1+jsZZDO1fYEdwqiU2Lk6O39Mj1QPHoFB/8xJjABtnSa1W
Zy85mINGWpbJ42QPGAROPGVVjDoVwfkX39/Q+qeDzm3KK60KfinxLlEbEj0QSZkH
MsgsXI+QthM+WMg9cMGMyVsb5hEAoAf6vysj1XjQW08QFRhF5rLFb29m6vV6adAn
Z9XZAcAOmk7af5hYY/e1QFsw77B9jheeqS5TmKh8eNFKh6ii9/9DDudz7kN6Xgyq
g38/wW9htmooer4bxm96vAtAMlKl05fJIc58CAmUQTbnP1XDFQo9LhMQ2wyQ7+4Y
Xom6SPQkWxvK/w3dh3uU6Tp4Iu3e4c72nbX8yeW9b9TJVP7Vpy2f+rwo4zVD08Gs
AZgBC85g8qXpkbAwV0V5t3sLl6bj+6FCD7a91HpXyeU3zWIgaeFI2kZHuiTGd1P/
qjCZehMuDAKAWDvxA1IachH7UK3fGj5pM1rnbrGnc+4argmnvU3tESu+sUbUnPCf
vS0etchvOI9G6+Et8jtyoBqKAbJ46u8uCqr3p6EzPm/Bdgpk++KBExVVgBcWr3JC
V04g4FlkahAdA8bX2wsoZ2fRsLcSRbjz51feg2/5Khl1mGtm+fxQ1CeyQG4xS33z
CIxN5PGdB/d1bphR31EJ1M7GNnBQ+88TkisJu4E8l7cd0c9PK5ERpWLWXEuQ5FzB
nfGbSnVjm6NiodgfycmJamMUcYFtncRqpLPgW52I+Jfmzuz02Fj4TMhQSmrUQXpF
pNxvRgLZNooV7CRHY6se+l7OWtev7Ky1WMv8NqN9uSXvzwtrCZZPai1U0E5qfYlA
ZmbUzz39Er5MKEaT9CgjFGCJziZbeeSqz5XpR/e4brsrNxyKeot07QSW7sbAbnIf
DdnO8mhltGS1zMTzojFhdXF09IKGaQrBGYxG0YJrK71xG7KeKpySdjaX1Fmew4GF
Y2KXzQNesGR0x5kMcMX0YNFb1KbbH6VtXIsVkRBSovP3RPw+28uNsq0SVP9rDm+j
Go98SLQSSlfzr4Qp7quRNiZ/dkXIQr0YgwPUiA2yNjK+SKv2o3LkgCk04efyuUYy
fT2O+Ew/3ozPeLJW7+3TZ3VM60FjKR05xP/rJeQXlwK/gURXhzleiPIfzxXs2wAj
U+0Y3RmIhEhIriaTgXfbHs+pHCVjJ24kgDEAK2T+GKAZR88gN8rQmEykT9IFlixu
5Zg3/Re+okefWTodBAzcbSkR171xlmR8+mXr/e47DOIe8cAhLE74IN5wJ8sMbyi/
YwlJnCEl/41WxdwrWGtD/8/kOo6muPyuup/oc7WAANrfZDaWf/pSJ7PNRwsTg0A9
rbysvo1n6XSGZ/CtyY26XBDs6F9USwD6ipy0plFGNSDJBEg9V+OInQEGpl7Q9xdR
GhYQFC4OyJcSqkUPGdjkhlBOysroXrWuM7SWLzfG85oJHKz8J8zgf7MPMydwsCD0
eDEORToYSzvUF9uODyof9sYPzzz0F3aWJHZI63VrrFx74vmkMKUsN6ATIF2BXrUF
SgZQqIUhrlF7HW2xAP1mB16VJBz0WA0NaiEAbQUonPDRo5+xAqU0tZoyLOM3iDeR
lFPpAlI/HA9s8gESpJ6HnDj5A9HtI5/0Rco6tSaNdDP9v+sV2HXWE9P44dgv/2aL
nSKSlSId1M8syCiSjCUMhevJlCKaxSaa1YjWdmHUVj6mr/iDgCXVH329jP5jiN8/
OWCtotJVUV3rvNIzb2nVw3OKgTV2qkedgTTx+pBlBk63U2ti4jakOG7b3F9SiltY
/cQ0XG7bucPskzjDPuyv2vhHgCSROo9eaUAOV6e4Ec+w1iv8Bhu1jNn9MSwsUWm7
+xQj1rfOGTUVpr2s8hNHyNUk0/cvgcZnI+2IMZiiieU42cpCUrneQ2/fQBJvp1bP
onMfkU2k9DBr3iM9oeA7DdwR2bgsdDXnBryeR2pzQum374LlM0ATnQBgOHLEELcA
k43e31co1zuvmgZWlZLDnrozO7GqAKpuLnSJAY+MhVTXQ99kDrlABKM8RFaI4G2m
gTLxiSdgtLi4Tb8JX6XH6O7WLVSJy+OKkniUmDGAhsiX+qP4MqzjKqvW1S7s54Qx
L27ui9xSdKypTS9EO8ZoYyVXbi/swUZMkpKi/77DUGS919a28z/pUp4Pl7tGCf6s
Ieq73K1u3HRb8WXNznjNVAFvsDlaQYVBMlXQYeD01MZuLEmnQqnDTWrFhg6EHF3r
CuQ4hvOPV1al46LEy06iyazvDPs7++G9cuZTStRFgiQA0KA6vYdrgjBIDfFS00hj
KMVvKuc+o4g7vm+r2lvK2oLgqLT/SEpjGDCKTA3mzF0mb5yjbz8CEu5dQm7sT+iv
2BMz0KhztP/WjAROc4y68N/89C7zldLuZjnwsMZax3mqg36SqWAdgKPIeDBhw4m5
UT94wzMA4shshU9t67shZp5w9wckYNMEVfaGy+86FrC5LE1it9u8cOR3XXYWcK/j
Fkqavxc9KbfHjRQnaTFfSMLKuu4/n6mZtKkVl4nQ1wQytq7GkIcQ6diY7P5GMZSE
4fs2g+6LYi0MldaZl8L5XcLDpq5CYSSJkSoW+VeHOpkVa8JG76F5YL+G8u2sN35H
YdLmvqo4zXe8DkwhB6ZE+iISX7SnCzKkvi1EWS+zT0TPxT3TsPomNQRLrSS0pyO9
DdEOc3j4CJaiG8ex33IrTOEwW7+n2tUvHryqZnCqXA+EjfLmzu7nMVDWDQ0Iy+A5
3oMiMKFUIm7qHeRlUkUj9JPTJfi7kj9R/XufmsWry7VDYU9u44wwAVME1ybH/6Cr
sqNU5niiVEKhZAEqDv1wAwjmLCuoqgQpkOZgbAVDGKtCnz75cWFtecT42CP3FdVo
jA1s1ZVUR+RAY+9wkKhhAcohMDOGv71SB/CqkNztnyKqx4xwnU87T4zGTHli7zvs
Q1LdON5GZ46jwTNX4j/PxfxIqb3fgYe7RlcfyWFx6J29qLceILHJTbCBjjHX4JUx
aiY1drT1Gz6v8HPA/mcch62TCRqZGfqEEHJ07dxlzzwh8ITiO9VqddDKo8a4L4qf
V9RzvvcDw9PPSi17GEuRHSZg0vg+2ZvgnJL22iuLnvBlm5GnTVp5IncS/J/UGJPQ
wDtw8NsxSzdHTKWYeoxV2sHH+g++mA8BDoPwE5i+7WmdjWRk44ll2rflb4mBkgl8
AFNkSbV6m8S8sT/Wn4KrKOtL4oULv8w8yu5I2GGcdZnZ94b4jVFQNFRBPs+EadFV
/KBIlID6KWb5xS1i8mAU6LIA8Hq7c9Mfpd9rvWO+CDigisVVuUh0hB1cZ8fCkY2B
DWQKEGIf1wqqBakO5hqc+HkELhcY09payYXE/vl/pd9EE/+b8ImzPavTmrRcJ3VY
3IQ7FP36JqUHIboVFsUc9EnCJNusTnLkcHM1rEGIijbyeSrHhPhZlOeL34bu9Yt9
DKEBOIdBX/G/M5dOjUKGme7VIIo9xeIZc7cW0ESB4jYdZf/nQRB2RCXqUxdpqyX2
xtei96JkDhUg3W5fWoICnKI9V5V80yZOhRkvBT0zKHUYDMXEqv1WisJCWr/Rmsxw
PPE4dx21Ri6O55TokWtar1iQUD/6DSnCUpQth4X2EG3mw2AEBQ53TurNOPEMXuqO
cZ+bP2hiD2FeqQ18n6gVeSAnuKubCXa37ueeeZeW9LTmA5Ggp2rkc9UzErrbSgEt
Q5NY4gk1VhVpBXHVt554bvbg2f/QLRPUsSqGnAw7RuJvDyaNtJHZkpSvXdxTQQe7
2ddBHLNNZX7deMJOmYxKih90Rm5aWc1FKYvtJh7ZxdSAkbk35y9xlW7/G70Xgra/
BftFM2HuOwbMHe8CVfLbdmEXJTYUiOr28DLdcESWVXou3xwwADPHR9x5pJuV0e/M
FvibipjDks6ewSNzLk3lUWVPLnlDj8/W2zv08VKpP8bEgN9zRijVXIpdbj9IvYAR
dUDMHnOWlTSj5pLbLxHYokPknOAgmF8xbFYYNrxsPRtgro97N2B0u95LQhcB0cAn
XyyyT/QyMa6eyabdTPk5dJlqFnnPOJqdHbkj5tjUib72Xugq26mOOE3U7v7o7TGp
slRZVejr+wZ8BjU5QFpdBQsXAL9OYKnqnA3GhQV9JfB9Pc05BaNagElvHeNzwOIP
7vRJXLL1u8p+sggBnysyfeCEe4s73MCKkfokp05zTmrteqE5M8pWgWKmxVqLylmx
ipZOn/eOFVHRYm2LmT9wynjSGI8f5vkc2U75+rp9T/nWfO97jzf9a12ICQp0tfg8
WinPYjzRNpHOqEgTR80Y8VfZVWxgKtQlV3WOY79oIKBkr9GSJ8helUBVvjpQw5bS
imNctP7meS2CXh77Rxy/Li789KvB2A/IiUue7saCMSQjNg8jvXpiwLutV7hB6kZi
YWQhhEEtL8v7eQk6ye51vsm8e8z92EkkzuWLSL2p0Lq9LxJxqC/6b4FcihxWE4IT
hOMAiKwU/e7qGagtqbnLtEfAaMnuYIkFbq+yjHwRu6wsFAw06UzOimbgU5VykVwN
ti1A4n9TMq+H1eqPfUnWSS496jRjxwqS9RdTGkFs09LEOzHFrAXUlIBZl8gdHEId
10C3u40m54Z+evErICKXCEOHMxmaNgeKjsCea8cZ0bu0tbUv39+Z42GE2xZNMaof
Vsd8Z4lULRNZ1alnBLCaV8Ybscf5sjk3Th/zm5u5pDNAmIoYSk1vl+vZ/SttSCqG
co++a02+9NOgAR5VRHydJ0Aknr+FklXuNKIACp1/KhoDghgVy/j2BIp5Q6TX9yOk
SIbtdI12FCSpJqLSpc40zozje2vWtD+hwB//Wce0eKEpKGMOfsVFrT2/CyjKVPsA
Yx3KtU+4K1qTE44XFrbvVLi+1CE9RDcA/x+mmCHFfSBln3iumgGqdRNieLWuQkmC
eQeu4AEI+hcTLk+135fV2l46YCb6OPMYPQvZ3uCwyaBV6lubnS08BpFC1FazMaJb
qRRYoAZI7yLz0n2GRf7L2ebrpNrRrzrInAPNfMlpzFrAoN0jj3MB/8IheAkZ7IQ6
P4O8YVxMRtFuhzynEzfYisgotfdcKSckDyeT16qyFewQYBYTRF0X2Lq5wxgRfOHa
hAlrSflsQvlaAACW6c/7NISmUn+eiODNbPx7r0BJeLP+yFNuVWSYa+D1AHdgnNhd
QehPHi49YD0wwSPM39/e2CIw/yliJht2mYWhBv7pGhZLwCjZ7QWoGs22eNzsLluW
pSd1dOvDjHsuyxE6/GOf44M0U6aheAKH9LcGjBW5b/wOKC/0i8xzCuajG3gnATkW
4F+5i1Gp53/y51mQOEbuFakK7hau1b02anG4UeRLCKXq62axHrjeSUDNblbMWyF0
Zvu1rK5/hLm1ETzRWQNrkhip9y+TpFtgYolZ2J6XUnMfNWdEZCCJ7a7zubHLQ2Pq
00ZOuJZck/EMKh/ASlWQVLF645C0KCZRVHHolfYO4peP9DY9JzFjSB9pc0CjRkZ9
4hUcwknsvohRIlPa7aW+Bp6mm7BKgOFrksEb4X/7QBw/xeKAvW6GX5ZNHpNeu8XZ
xfX4vhE1sEl6v+0kcgHwB8qm9zbcZNal/kcPC48JShuNtmRECctsr1r2bfVJrsRv
bnJqTEr1CleVHPby/7JTBXBsaeUXhwwY9E5YOHnEWEsYcZedKpbVwqoA2+Idnr/r
gWmrnVpTizoS6+uqjhyOW8m2MRWNjCDNHg2mYSS7dciZC/H5mE62HuMqjssavz9c
wxF2Wp6TGtSx+CGw6+wIHPKs3wZqVV8ZOwe8am0Mmm2qGUTFgcQqIitpcU+ICrAU
CkvFn1jDHIutLFna93ehKaMCaImoHMUjdoHAirfkaM+dvevSCyYofM1vIuKCAQp/
e8HHJYRp19ZMWsXfFUOiqOG09pCYwRl2AJG3Rt2l1W3oj4DStk5RZ/DMPNednhjL
VNVPZzyeXBTDoVaxaK2nz+n993DcdDwjd9Qy3vRBHZ5rlQNWdsxe/bsf6it+mkWT
eDunWcffUa/8aGYJewtyC1I6m/POrN7p2PnjmN7wbcK+7GYULnzvWBNWFRKmgcGq
/R0bzNmCvFON9qN89jnjyEEeFGU437+pjqMmsgHzGX96on1khVd2Jf9/p7YFbyE1
ZQYtkCD/0dGXOfOiG9ovm8UOaPM8v+lD8fmZWj7SXVOj5Y8Pf+4wrRe0aqSGM4RC
zjF0/c4p4+VAnnBv8u/l7rCl2xLSa16GrnuLzlYcEuA/KBHm/a0LCqnRtUKPMBHh
d0MFU1FcOl3vGTLSIqhlm/BA0y+xnq0fHjoE0u5A9wyb0pgWVzU8zOiJ6sip75yl
OHvZ5Xg9JVsu2x2yDi8NvPFfX6briSzevCKBwQZAaU6Xo71uNlYKcTr3w4fDWUqA
9ri2TGFePBNP226ble0UffVzVWR9u8xgUpjmO83mWVwI8v2X212SeV90BowMgcJd
Dxplsr3jNm1TQdrE3jTwvR3CZSC/Dk6OV9hvYFJXIjw83NtRy9PiDiGbdCR54pfk
pfrjIZBNZZA/YqgwSCSwfrznnS5yKDtsxj1EeJZSBihmYMTbo3Mt8XIfzblHFF6L
bahWjiq4z9kcTwhxzNwlprGgSv5majKx1488+UjqBYJVRTDkhLiGu4H0A5s3t2pt
9ir/awPPhNFAvuAmNyVC9p4JzSmPXaOzW3N1S002+w3DmCQgYNDYMCXHnAS0bNcL
eLNW8yilTME4/meQvlSPXIWv1uKPDKzOpLtR9my+nsjKy/OjMnIY4YKYWLJQZCR1
KnuTkfsT/uBsFt5yZ8wE0+Xu9BVwHcWLLju7EZoOpQqm/kTdHAQy+3nqJ83y3NEb
QUfuJG8Z1Hmw/XbP5yxAu1ASrdn2DHoYuoEpSXaz3InOFBFcT7f5shhstDy4i+Xv
GLNMCpzCb2ETMU5Q3YqHWRMwWo2jnBP1KYB0dvFy299wpwL+Hg4q+zLBaAzA8H6J
NmGOjFdQHVrPZWPuFq8zPs/64sakjRdfQHSObVgUtFtDKOkNUleiR+stwyy5H8C9
OVtnkm6olH/kvB1r+uBJfr7dj+WkLo9NFHKABeHQewSML+dSi8IEFF2SZMAWI8mL
4gAS6GA66NjzBRjJH/u8hsONnDuDb0rDvFViifS71MUI0v3VrcBSLBY+4iXE3C6Z
W21JGjvd8N1G05N914+47IjxCUFO5ovVXFjHzrlKsUKiAK5H9lfpvrd/Qp7Rsz1Y
1rd2b7COahiM8nPn14K1CfAw8+UdxiwZtObyjn2t0Adw7uYlDJ6KT/kFmgek4VS2
oD7eTT8N8UzUSSZlH2xNKno9UUtUBrlSs4gwBKVAVWb2CY98xr6FSc0YtL2ncTl4
PjsQm1FFsNpAUkAYVmKWrCkHkXKzQfmREy/MGSZwY7Sf5o01IBkDK2d7CMcvohKL
G1/OyLiQAp3HnMuQBZWJqpKK/4XjO4Kr3IElIBRclUjO1JqONi6neTy0Sf7tWj57
2iIA7dsLe2noQZdqy2b7URx2DP4zVVBQ5+UPS1rDlQ+xVAOnZB7rkWHHNyWeN32E
HgFWtSc/ZYjoXtqi9+MbfRDLO2S+wXvn7YIAVxx/jPzUSmJ8oMPsTXVDNKo8DSze
fBZN+JuOovYjrDG4M7hRK1JuO8HsJ6lb8+ZzEi5NVpl6jE3ejEfY8IgcighuqH+R
gArtrSScNqpHZhCMSE4eQDxNMqbe/env3p1Fhwvq1b520d5mbgz5s6LUwZYywIFo
NJUQkPvItgiwiD1WPil/tVNWt7wTWMq1cqf6kejxHU1LpTQQ2Z7bXd23ORW9B5Hx
LRvSJgGnPS10w4H3C+on+hiTxjlSmetvGXfbdbPzVuCef+P+PEnsvmNZUEIBqFk8
2Z9YMH+SNHpQsqIcXn73sRU7fleRqvje+dAcULc1wyxqeW4k1j2/0FLjUPDtnifz
O8XGIu4/YzJM/aLg5/IauoA3e1Bae+/4AP9/tDzm0bVTmzUOO0H+3BUzdH8lte8v
8BHKzhWPOYtbwrNmHxVXVmAYGttGPyAVnUcRDJmgMoD86Gzot3DxS1YboCatP1N2
gHNme8lD9kQhbvuF5p5PSfodWYlAGHz84NKyE4BV7mYY4rNU6Kjt7aPmEpVchS7T
jqF7mtKrKtjMyImyLohFz6u0VcqoHS/ar+SnZA2xpluSDrebg6TS4y6hJWcJ2LPB
LzlIaYPh5R/3IBXMuwlEag/AwA3QTWTNqsh/NfEnf7m4XYTfknhX3tbv6S53XOvo
nMVumrP4s81xsZb7JHHP0YqlkOxtwzCGRTNNsSqnIxduQEs+dC0lP2YKkBCemfi3
GsgNHaPAWuBVpyLBtIWTO9tbaDIpkSuUbx2kdfnDPruVt/Eog1trgQtObz+NFuYx
wpfv7Np8cpm1kSW5avhEh+5zvyEYYpIvyE14pklccqZvlEidwbGcKSnux8G/pcb5
fOdcRSe1nEMgQnmK8q+/81Qes6+3gAN90G0b+Cei+ZthQqSYzERiEPH29KAQE5Lv
BCgFAwKhaCyVQFe2TsulkNyHhFy3lJkz9xp5f23+8nr8Ti1uiZLzgt2GvJ5xGBWO
6tQgJsI1PvOTOo9yA/lk8hst7JUNxMXKSFurPweange+3rubefhizjAnj9Lh3mBq
1+V5HRXabuhqDRw9lVCh3sqDxHnZyM8sgquAQY5HiGkq6XhL0CaI1h+Nr+F9f2C2
0bDxrbxo1NKMHZ0UrCWpOPOJ9EaPgBGRZDUjs9EsXts8fTK6FEuWnhGjf5Q1cZT6
5+MfTIl/TiD0ml9Iq0apjTGWdraCyKGM93xEuMsuwYJ8LoMLTC9zK05LJdZwDsLq
MJ2DsnK7fTpRPuF9C/Fxd+LPJAtIq3+RijDWMqZUqu1E+Xe7IyA5vVNn0+68oerj
KQuEtwSyKjatkDESVzyNiXm2qxXxyWV1H5hXvxrYHLSGd44/P9NEj3oqBKa9Ijkb
83C7jAITdzAQnPv8FbSrlloTNW/E7S5L3ahukHDy3kTCfwn7zcQaLka5hVbzleXM
zVxBT3npCC6gMSNWvW937ZGHPeGbYT+NL9xjpLc3FPFYJDRSMzRkFnmLjy9F0VEG
g1cnruLSB8wwWxbdq3935kxoc5DCet7dRymDGxItI/R0SQmgprwk3biS4zPqOVXG
adFm7JAgTTU8dLJh1YxLEL98UJ7oqMRKNaQawlEOVoUdi00TZ6T0nufo5dZEBX8a
y4UVjAKdAGC5ZEFAsf8j/J6w2VLBMpD4KCfpwuiKhAz22AeP6RSBI+5d5HblSeSS
fZtYw2HU4otpzT2BHed+ePhIUJ3QbqZfONvJ3+EhD86oWQon1YMASz1MIMZTyR+G
ucCjJGhW4alkJ3MRihVYoxrAsqd9OShUKsYpW9WjyQVJL6YN6sjvFXeW424wc1fX
yYOJkRjkxnCpcDJftKpm3qdcSy0zU++xAEdFxO09lOC68ym1OrDKoWYv2W6Tka4y
qBNvayl+MqFvOptQ9kiTIkahWYTRbcW7u9zHY4Up78XmUUCvs3lkwMUGN8GCNVoo
Ocd3qijLrvdU+7Va/Jhx211un7pDNzjfoYsAkdjOH45nbTKxcrSDRjTFh5R1kcr/
UYMfKbBDbdioXiR0ZIINTxCQ1TB1V4/OuTY4AInVysK3JCw6Jlyz6gCcZbHjQSlr
zFHGbcv22hHXVgPExeTWdrtuM9lVetXy/SlYEcTdnO8cF3JDEZ+AsAfcRjD218PS
wVdiYTPJagIBHF6amrbY4j8r2h6LatZ/WKsknc0XZrdE6t/0vf0uKFqftEA3Cij/
TmvYV0VD/QFDjZuOSs9nGUAziTjaE+qY3y3ZZsrwDhQRFKPg3n7CJIIaaHshkINU
3DnEo80lhKC6YhmUpOV+46ulpjFpI/uMdz2kTvkE764xypFBukqz3ti29KoGUOQ6
4uTbp+eMC4p+UmozfIwjgxJJfOsX7QZUFO1icdsKnoLIWk+D+V2b3De0sVMn8oFw
Z9x7knQbx605kM+3MCrQSjU0M5assYcjX6PRGUsi5F+dV8OtVWjcpC0UwNtsWPvw
CePCIWyUZpEAPTOfXR71IaDOcGdkPvJuNLMb5TE24sjwPUBRB/ddlFAd2ipRV0+g
izebpp8BZO4pIU3XC5681282I605S6waIHFAo5w3Hjy5ewkEwacdvAqnqnS1Nmqk
ProjFz8BO+Ic+/grDaZNeXGZ5/ZPZ+LoZeJBw03pbUcxfiuPjMZ+IA5IGHmoNtCg
B6EXV/Sgo+qmIIor0LQ6pThUDzKjd2+6pg/phPVnQM9hGioJFrXcPKa5GdSJ8lqb
7Ks6sTvUVHalTFIrWQb+YITNMwOtoQ/lSGLb3NfNaIpk/cCIdYqOCuwdJr2wWf5t
CMJh/FIQ4qxwJPvHk824yi4JZEIi1L+9BvovBIl3+FILUNRoFHXbDeDKCpBa8V9m
2Kd0xKk2bN3tzNXuTkbpHNtIaBfGrBHyE972K2r2eEYGEYPC7UlnQADTTVZwXvz3
KZPIkXptGEM1DRu/BLwluQtU4U6jZ081yGPyx3zesff+FvLViZZcHER/V/mNj7Z7
1fH21k31Yj4DH0Lj8uvZ7wJ6cBYhuq2Xoja4CPnAXcj0DumuKrw1HohjrXfEGA++
mMm1+Jmz/XLFTLUExbQKKXs4xLEFY9hM2OugGEoYMvS2adIRJ6qh1bAU20CyJszB
7Y7cTCG6vnp5rZDbtX26p7pmpD7eww88paJ0gK/D6uH4KBDV4hJsQGMBHQbEdo/+
eWL/7w5ie1c1Ir45OBS3ARJ8KnBcNMZR8bsJYvspuv3EXviK6IdJlImi0+i3nUWp
mwrT1ggcgD9fiVoFsaCQdaI1GIf3mAtPQlJudpkG/R3jCH0OHS2mqqpR/zaQiy2L
EL2ouyBhSa8gB5AKn8bH8+fuaCyv/ikavH67SaVMUmm+XG8Vo9nBzUtnQxQLYs1S
OoU70NLrSAy0mY1pfdGkJ+xhAhBPPBiZzZ9Htb52ZiXeWHs7tEc4q/U96rlqZlFo
2mKIO09ykuoiQF49CLzdKNLiNku5aWJLiBeaCCPvBT7CFs5p39cU+M2RjFL0ZiKi
BRJXxHnmXVTb4KjYacpus4g7txgVyfR+vo8EYfm/UsBjtGCBHnNZoShvyYRxflYj
QjXOvb/Iu7lbYMw7tYs7eOoywj47WcFj+QIT/HHOwe6aY3zc2y32y/smf3pljuY8
gAujpFCtkHKYp2evfIV2tRc8J1xuFDk+FtNfIea/+RtkymaYgk2GnO1rDGDMqyhG
qvoWc9uSNvGibinUavo28swMMtwVQMJgsN3r4HUiQFLdQXN+3+ARFPqZvBOAJAQU
ow/pfTXwvBFK38ME8w9BsPqHVDcXSkJnYjqiCx7JGm11YH4m4ZT+mtXs5lmUNoCi
DFMwhMKzuwyWJwLHKSQjF6ih8qYyKmFV8fp+gsQ4i/eslTnZPvcVX8AnI+vxsWsV
lLAj8q26pF30IcjMbusEaAt9fL841XBE6SYtRLF7MZN7eOqsKvI3b7TirP0ZAObK
lUvCHxUNa8pZhIX5z4TmB+0F73B6k5c06NGd7DqIdC253SCKuAevZOF9Lmpr3DpH
sLTi2him2ZjsfN8s6eT2JJcHC1HTph4pj0U6xPN8hK3vgBrQxjjWcAvivCbub2Lv
OtO0S2V0Pd6tb6FV6bjd44plDyTZSSR5USDsqpgUXfvDl8KaPOf4YIj0BsWw9AD9
CL6XpohyUyKg/OPs1HQTpsggQRVySdHRkO7n2Pag8UacbLI67xKCqq9HEJV1CC9c
AIssnnj3up3jxKjdGAIH3ympuJE9SO79UMEuxltDgWtLSsvMchS3v8MzIwmACVVU
Csr5AcI5ZibQ/K3wNPrEtFvwTx2x60Zpr16MTi52KdcEArLOAUsi4z2UB+wh/1xD
HrvJZLAsm32+PM+ZtJZkvgVpRcIu0b4Koh0Ajc3nd4EL9p7D66v5hy940MD4/fEj
sG3Yv01Tuival1oTvnCUzmdMZ8RZu/2yE/8gO3A7TlprK/hcVCl5SFTnUyagT8iA
VguWym2ts8t+0bvt+73LbNodp7i9EOYCJb+BiiEIEGFK1r/IlFMSmJLaDMKIA6hs
f2qT3G5B7NPhOaMGtV+/ii8zdQxNCGQjdWsfRzfJZI8XKH5t3UoH2I0VbQdoSiJC
2H9KMQlyyVr7+cd21SVkBHUntbgd5iyJf2rkdsMOgbLqJsv8padKlZlcyctG97pq
Il/1vNjq5xurUsUewl9DEFbyrntr6yn9htSstW9hYPaQH2FcGrb7W5ZHuAlL3igk
84RveAINtu0m4FV/wwrf8SqVWJ9irLlNftTr0VS9xVC0u88QevooeN9RPid0bE/3
jV1r62k2flwfHYbIe4JIzx+EHM6jK3mBzMymHl/W8RC6rNuU9u+d1PKakpD/xYxe
WAJWURTwZCypmQ+uSv1fR8PSfmGlUJDMEDtdOYqAKoh6wD781OLOtKq3n0MfSPQN
e6kgWIEg4FBEUc+H0ELQeCYVjTmI1Mb9m1B71tNfso/9cAc/io44aPucrdAikTNK
fkZ7XVZMy8apQId+QDdCmF3qAddVx0E4dnrPCGPvdk2qYuHpl4zcIsR2XqBV4gCo
5Xb8KbpiM+5qpaMJLId/LNXv/igz2uklqybEzbWl7YEX0/yj6WP+Xffmoc5rSGLk
9DvqBKouLnx+5IwtTCL6EQh3R0U2KGMk+P+nrWY6JJz6aTUppn25vnMlh0y5lrxe
rMW7BhJbD9my8kOEFzMQo7vHriGM3WtKw8Is6W8EL1F7sY4VVG0Pfrcm2BkCnZr+
X4/DgFkzcUd2Dz3nVip8HeCdEwDK+Y6Dka743QfkTRcBF10Eza7a6jKPfkoXL0Ji
8yVSeJ5DaYw4Y+6V50W5+3IOqtgQhDdxWZyP/vKjB98+P+J4YCa1l2whe8Y424CU
DUWFXiTypX3MpA3KRv4Cw/JQ3I38VkdJfz7y2aVP4CIkor8GSBUzds/xv/lwX3Vx
FFWBQUeQI6XudQqPSF23+sC+GhNfLZ5rbx3eLyUL0Ww5OGVMKCJx/wCk8IUbhEA3
fYt7kQFXDFJYKWS+FLH2bU6bOfxEq/+WPXTe9qBnIJ4=
`pragma protect end_protected
