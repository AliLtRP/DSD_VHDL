// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
FSl+Wf1RYDHdP7+5z8GQvoSgVpc66h08lH+Rkb68eA9HtDAunE0wg/n8mYqoptJHfCmJpYSp2QR4
a4LVuDao6ih+f03YwW88F8dcGTY5/VNaK/AFaWYkDnHzSOWNyXQlftJ0foIK86bWw0MdnN/q9/co
tY7xefQDNBkd96pkq3m0hZtvFdUL0nVNNcly9gxA1tNBNls7+tw9sXdFiQ49/hiofRXpgV6NrT7w
ofKjr5xE00jKva4+GUDM+pJCmALLcHr7o7gtwzZqF21Y5gCl7qCWVzUzKsp3aVqv7o2tK1jhgjd9
J9YDBLS6rbS+yWZVIE5D9aI5Z+LRA6rq6Nf0aA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
xmn+KDUu3qPS0cQ9aL+Wg/MlKGgiJ6yDgVQT7BibX2+x2pkmGqyTkeL80KvQP6jdSpiBcWIIEPhi
4oMQjMNNOTXYSnY71kJqxwBUL6+G44JrFzdJuVJnqkFYoGzF8zcJh1it0LMRpQsUGDcUCwojeXxt
uI429FAokGMiJPnoxJI96Y6OMALZmM/5V1OVToL+aa5b8NMbBIX9V8mlOxIFYCvoRbxeA0Zqax0/
LVJURzYqrWQJ4YKp9lrnqtLaIZaqw4RztYK2VccIejIVGWXON9zT8xtT7oQyYvwwZYSBKpqxXA0m
HejtUeSdA1Iu/japLMEAmlN+KWmYAHVsedkurvg+BOjd7azAE3KUs/BaOoYrFyA5LnlPxHTw0ef+
Ao2Uh+2DSntdsYyJDEZ15KuzcTRrjQM45A/1LB2Qj+nkmnvVsX+5j8QM117pADEyYhwwthvIZuSo
WReglv04TbY8MpYjB7PE/c7OGDZ6FCNrPZvLlUiKrSzyMfmK5scR1ShqOC07anikJWQVltIT2kXb
qotGItVQ6uEqPkxbP4cq+hhVwTjfBdHXNPbZJ4E5b3F3T3YMhMAp2OQ98v1WAaxKMv4FKyRGiQpx
yAQ+WT5+5gIQmTFKJmGjwwsCtncvqTbgR8969OnbwGDe5P7BsLrn4PGLYBJ27fnz56+WCvSOYyh0
KwhWN5OjV5ZXZBanuxI8BU1IVOBtG4/bDwKGqLoJqO3jSI7voHxOHMuLV45Fl+S8tWyrwVhxo1ac
VwDdt1/DIrg26AbzpINZdPTs+dhAs+L0BJyrVT7O8WS0CZ7S7+aYS7R0KQrFLCFHTd5HF8rzvDLr
0b9gpTRlqzSGoT8KzKIoBMCIOi2HIJUnHg2MNiO1I4fI5ASnzPOV9ERtsAB4fnfSeSrkr0RlhGgt
Y3abm9uPp3w5IUJoS1A8mFsG8fstzcVtVysMYmJgQbX21idmCF68R4GTEww1jeukSv5RDBCyxG2t
0pbgO+2nugHyLzXovoLykJJ28IDNMNpG59SLVUS3HIlpEFoiQofq2K21JnoZ1AZx5hseRfrX9zzw
bPRuuIWO4xMEc3o3VoB6Ut5hJtBFVzTuBpBBwJHPg+Ioms5X00sQRdIPQog/LKxuyo883bGdGlwZ
Gnu6EiOw3Jggc24OvxYlcLfNW86CNxsadkcQegh6SuFnAxJozUcJJun0tsJft6opB5HrOYx3MSo9
ZKfMlKJTRerLAr+7MqQO94e8VI6E3+IqS3DK+i4cFszRugMIeljM3V0D9I02MqRLvRlgWj32ynWR
+Ic2Wy3XJxYYFdkNLChIDUnqeK8gkNKNed6FmAK4I/tlGur/bxiADaKW/MVPlnt3NXolcnBBi1pG
gOxT+w0K3gvRlV/lutWPrXh1w4s1U48tCnQLojATox2PR8LpvqJzDG5eT4JfzYqQdoVdIp5Kjapp
gDwLYDvBSeDkuvbWePknxzh3e+SXhNHJaDJxdWRJVhBnG6olqBXlEoZ4MlQRjRbF2U49vIVtLl8n
ZrRgl5DDnmvyRKqTsvHhFjA9ASz+3eZyrpN1E6LgmykWVepYAtv+Zy32EpkmexP7rkenqGLsEv9W
2XtbuPdR00juiNy11Hk54TGkzDcfagTIv+6R8sm6b0tuRTqo8bpfUKCO2b397ip3jG4QcwaLNMHh
YiGLd/oHoyZqqiPYhy8Vh5VIIgX7MNzPQo1MIAV4o6Tt+4d4Qa2ndZ1+04lEMmtWgYmlL/04zKAP
xrFx0c2+scN2SHGbYVkCFKyK2jtk//yyT6/363CfoHcf3kBg2EI2DgAJV8Np/prI78SlqCoPZSAy
tmLBd4EOCBstMlTJVg0pcamXk9EVPjNe5ztoPHYZgpXZowpevDpSIq1/Wjayft6vHSMFEiTrut6U
bvcVEh7soxmFfEwWPsMB9+N/wnxVAqKMjwFq2/I9e1WpjuNlLuZvLOxKSpiORtAHh85ffAr2Fkzt
ttLbYRqppBZUinUAfTmH4DqlzOrQM6bG30nW7VjqWq6wtpXSQeNW9R0f+WoTlMquEpMb3R2tzeox
QvTlrhqLj3AGrA03z5uB8yaVufgao8qHEotrfIBAPP4W1whpIjgRMlHmYBiepuSv3fwc2VWtkKMB
HOM0kvQuHsa5yFoUNx1Rbfj3OxsPD+nnC9M/v/+S0oOqm4zvEPA0xEBc+qwz0PGn+0XEqvby4OEL
+kSHSC5t8Kt8BIa6jsC8hZtTP7j0Nky6gyuz5HYRcH8kvj0d8ciXJpMX6fnOmXvqVDJLY0yxyZ11
05t7oYYUZqoAExO42Ln+FFNeKfCZfzTBJEQ5rFUfCyUqwHV1+MXDL+z/yYBdIGXhsHN49mhO0xja
Olo3KnhXZl6A1hFiFtfd63UoLqKrNaRWtGEFB+p+37LoFFsYDVY5q0xs3uRzCK+wY4oItLaD0qJL
gd/q9kTmAPdnwKTTL24fDQ9iMhxhd3njy7R4oLX58C4AxNDaZB25d7XKt8BXbqjMooVleub3U1GW
WI78L8rOrBVzaMmGZ2SXMchzuuhbc0ogG3C4RnnVmo6RExW6f8KoIPEjrPwJz2QB58Vvluf38nyO
g21POP2G8C7L18ILLGfBIqabVd+RQxMnZKsUHxwkEPfQVL3jTRX2fTfopndhCN5OxRNpO7OsYAcD
IgBRfbSFPsQ7g6FiuhdM/0ddShWOxwQ+F0+kTzKhIzX9gfGFsz0zMyO8vaiDN9b1lcaCdmmObnaL
y2hVuoasmxe++HFo963jAt/KFMGHnVwsIVkf9+PLuZAWY+msmho1gZn6+TKS2rFqvPY1ONaqbhDP
HT4QBDLj1dB8gPsbqh2Lk0ahV479izwVh1iF71gcJN2OZspokt0X0YPlvIaSuVTRAy97SFKDycAm
PJcKDThTe/CnJvO/EjoL2gr0aN+c+US/40PeO/8uz5ZFiTp9mX3+OCEuDQYy47rfoBexEI4BylUX
BT7smDuh+CkoWwRz6/I9Plmg1kZpCjkqEDZkbGRMJCBjVdIm2h1I/4rJf28ZX/vEfv/Bzk4HnXjK
yV8KfjL/jDp4OrNsk7zK/clp8Hd598grkccyhdL0nUsZ74tncSzLEXerJmA2o9lDnhvoMrPQFUC+
ek4ihOpY12p4w6XUIaKLkUqgnWLSTjRyYXqNBcqNksAqGuHw3VaEPEJtaxZprZG6ak4qHxSWsFm1
4TS/hQqdsxozw+82J9HL9umRCTmT5Pq+vYIvi3UYka/PGqe/UaYWjHwPs757zw8Aa6oh3uG9of0W
472V/3wWfwQBunAz5BWrzkaVrObEtMkJirQXMEeX1ZnCNrAsnrUsblWXNvjADfoNVGgUex3YAdS7
QaPp3oVNnT7dp9qBNtjBj60ZQTn/bo/tb1qpU/TCHLsaRKb+bVNuBTbaGgGIFWscwvyOUmjjVP8Z
R//XXdmL2bCayEbfMSN9f5NZbG7EERith2pQRLzvUmHPuGa4Me3VdZFMESE/P1GeZ1pSSAA0wpz5
wY2+OHlSYBrypgL/dlkJ3dvbsQK1WJIcCEE7SMYGBQq9cLRLAnbx/tYYJkE+UcMoPsjOinXze785
LAeQr+prouJ392ocwYCLRmzWk6XYUU0kCQ8ct93+zbII/vYH4ZFaKMG2zp73JL6HRPwNA/0DRtQu
8uk67ut5pydLgITbbnekzh3Fooci7q7lu2n6abH16ft0aGfKRZnCf3+VZ91IJUajVES1hujiFwMz
y8rMofl3b1iQZrB8kFD/5MqYM51xBcAr1sS4F9V8MLYbmvUFUq6Xu0tn/7WVCwysxIKsIjnKzDdj
T2RVk7/7yoICTSYCjUrAsMBXHHVUx6hS5TcXd+gJn2PKA0dkx4GrHGSsauS5aWmyf6JPm/IdOPhH
uwQBYRZubXQUoOXNOaGNO3ajC2yeClXJrbOSOLTooWKPpXliZ6JzcpZ9y1B3C2Z20mYQc5+Yf7wZ
HL1RBt495A/AfwQdDV7autdFyBzOHsmCCV4AgGYknwWAg5uO14Xu4AzV6mWd5y6PZH48fRw6Kk3Y
Mu7OmVuc9FEq/AN33TQzGZlvrWLolYa2IObjcgnxvhMUJq3k4qnw9G/Fbj3Lv3ls/OoineHkxEsY
abuwG2BN7g4UyQ36kuTwvzJqQopSvc2cnRI83hgcWgNHZl5cgNwu/e8wClcQU449aIpAAke0t8uX
7I7kQ78RxT+cmmGBKEI0OmKd4z8R0zmjScqpiHkks3DxPQ6hPft8FtXrpE46F+s9q4oQeyRQGQkv
wxlTKfFzoKH8btGrT68paOt8JyNK0Li5CKOBB2WgijyGz3uTlqxS7zioeFlq8LUlGVgHhmqYHSYZ
+9EhfjjvZbYTOevHfvO7QARCSlvMlntM7qTyLqMP62avJEHxrF8LszbNRnqZrJEJKn1wVy4/e7VY
Qox5WfSeeXY/JHJqgO58uOY/kIFIt3Ha+haFTbuUZQTAq3b9zBIlrnKikIZEEQRT11WHn9FrRtwL
epotaFXbxkkLoE8JEgQa3HMPH04FgSW19UiPAeWFoWPSRSUFzRJloG8yCDA3xbQtVc0rsEA8jLOt
4YLOCG2/mcpByU5UZYNmBeI7LD7HVRRovkoPYea54JoyYtKTPaM7Ta04Ng7rpPj0zEuDJ7gestGW
tbHYp210IuO/DUz7M0tQ3VcZK3kXs3QLlbblVnTCBmL/ZgwRGCpsOVbPkkjAyOXmgen53vcwcoBJ
KZmzonNoUfJSgeEt3ayay7dV81QuM6ePjwTulFFpn5RVoGwh0IOMUIDWhwp5KjbYagNKRFgCrCPD
uh/figNC07KeB8NSmzI5SxxJbMD/+274QtD3OBomCdoD/11oXok9m+qRLD0W/fpbRZD7z5sWQaQF
+ZP9xQND2jS+srYHholr9SrgfPTv7XOUnvqCKT25D0DdM6g9ElnhwlkZ34m3sMZSuna6dui4ygV4
HfY5Wiqno6I34kDVaeWdLQeQFU6o7lbLRVCBacssyrLJroXcl9MI8E9Q7OMsVLFWUUbjEh1d5Hhv
SyYspCx+5xnwBhCF0FoFnDX5EcvDlK6UKcBwD4RAXOl6f6toHYHL8dh+2loPb0KhiS+pZIDS8Ldk
nGMUMHWwMSVxbGsgQ2eAnpITKlFFKJXoHLTLuLC2CHbIW5ka6bVzxNkUc/vjHm0Cxi0DMZ7P53SZ
W1pmFPOVKgqB+zk99WgQFJNJeqOlIG/lf8NBlsDY3HYf1uNVNxu6IZFk2mlZaYMVCQPCBN6+e9E7
zCsXvt4Ujyiy2Av/uB4vOt7CJ8QRSFyO4047xXlQ3s/HsVI+MXU44o1abzZhGCoqrw2/NWo7CWNd
bNI6VLGujNiA/j7HuLtaJlSiTQL8GpXZ6ez38yQRsHzctYoy446x20mGhOMQLmJeb9aJb4kW2NJL
qMeC7N3KXtFIL0YACkw2bNJLzg4WykQADMqG05GRAIV7t89d64ESz+nQiLDQaDXoWAovemBHDWT0
GJgJ2ZaYFEJX8elNOUzigE+TKFI/TVB5maYqCYCBU4Ni6yVsqb3GAD1j2fR2q5sM+BMmc/8GPtwe
bf4Z7dfS4aGgw2XOmzN6E6mYElR9NqGreGXeG4EgaCzPy34EbVAD6ehj/Zl/YD29KEtDZeDkgJak
yVsmf72+cYxvbfpvuABcjbXhBfxKsCKga1mvRQFC3361fMz46gA18X/lJVXnssur7Zzu8mlCcZwp
W/wbz1znr0IyhQOcaJHz422bVVu13NFjHlZFNO+E3Mn5rDXHY8nxOxCA5mK+hiZQjxJcmbP0i/wK
anENZUqK9OFn2heDExQ4bXE+VcpgvaqT/BB4tO0fHbdDe3Tniylxrb+IvIkmpg8X3MZ67+gxayoy
MQYfBE4HFgR5hbXAuKaRVH+EOVHWEc59YMY8Mz2yjxyYVnmMnM3qlAqCgzaYsFNU6voP927YYlS8
/EFyr0qqG5a8lG8F2TjKQl/I/py7LR2rmByw9trO3a7+S/1Xfh7VCDpSpJ7lcpnkj5oPt7DFglC3
E4UueizFyVmFwijZe/xrpENM36YZ6K8qMQLXIjVwlNQpKXUVUhxTBcATZ7sgOAWs1KETB4WX9KaO
4K5EihPlP0bWPlJCK6C2ZcTNBYo09hbWRi6Lx6j/LfFxxmqrnID6N++BEt+mu0xcHP1J3JZTAZGu
HR3ZDQVY61OutOYTN1Ozxa3hemJvL+7GxkHp7Wpolc7mYEabTwndGjnuqA81gxObyTvldfDPVtkO
paAu8KaRQFB9qRBja/CHriflF0K67b8kd1UC+MmeZXnAtTmJx1R0g4ppYZXTbwDcfliGsF3oBK7D
hFgQHLrQAuVWqdYMPvxQRBUnWXekzhztIuobRqCZm3LeZB7fbbQlvSBfUDEUgl0K/CSJZO1fFgZb
6UUv4JGnwrq1darJw0DXKbWytTA1/FQxd41GXGL4WBzgX/UOk3s/nGepydbB2bDrGCtE0yYE2D9X
4t3g06Hk7WsMxeePzBaDIrDBGU+XZ/ZcdWTa4x3fAbU9w5wWkeRSqwTqJ7+ZiLuuaRcloNSeoTBY
EX3qm3Pp5ybMLNlF2X2TMOCHufOn4rJ4hU5JFTo4uV6oXRWoOQShvM4UCRUYHqHBOkTb7VN1aSDi
nrFK0MD3ROesTfPfpsz92tbkxlhf+ySlIkrTfzl+PgGmFdPOl8S6b1aJ6sK5QSKaOSKs9JuSne+K
9YRIKJtxHKU4ZucAtxMFHfoUZnNG3mfVopUxmjGMKU5s6UrYsDFjYmwSZZbRgezvMtqbq1zOUaAv
9JZP5P+1lRBUJLkdeNF4hpId7uCrKiQkfEd9ej90L7FFmpoRGS8NoKxtKAk2kWwGfqy0T9kdDcSk
CD7uIDR/Ev9RQPsoc/EDrkr67OF5eF/YIFJLgelCLYFEnnWZJTWLfyG7b09rxDViBlbLWB59rPr+
vZshlZf78HiU3WuEHxXqIpd1jKv0NmWqT+IkcMIHO70sdDhTNNu5YTNNx3yJd0KnyRON2J5gqtSP
nSheyWKwzl5SqjmoE2BOb1bswPt8hirlsDCrvRwWDL1ds8CIkOZ+4ysFH7k2P8TsC/mu584kZPsS
F5XQvyvRfvrGyVp9gNEaY5qXjbcm/ry7JA2NPaUGVnwPNPhNJ/ktv7Vx+V7uqWz0Do6icv7EB0rQ
csAoP3uYloz3sBWF68dd2/CWAn5dXQPhDUkU0nskYBxK6WxHHx5uIXIHIfN1Yd3q+9ZX4fTYN2l3
bmSKUhCknIm1EYDF8gFJc3obdbMIS2DgOP4Yp8CkDDEC2BBlyp67rbExHgEpyGbVDbTfmtKi8gou
9NoLXtNSYW/7DmDwNTwjMSCEWH8QP3QUk/lV4SnBJ0WUmm5hVf2LRfnahfQHDQeZtlbvy+iV83+A
vdght8HjcT6iy/MQRsP5o3kSwVvW9Pst4ANIJA+aD/wT019Gqs0rbDVEHKcjvctubosKaT0t1TC9
EC2IhUuQkYRUrEGvI7qlqghVG+phBHloq8dWx2cK2s4woM1HA3v8kKEID7qsgA0SflKScTti4+8u
oIi9Y6sJ3WA2YVuHjmoyvpeRYiX8VX2iqP7GPKfc01BkH+VxzAeCGerSJYDep8WgRwt+bOVEli4L
JbLHczcJY1rXWOtTQyQsLVZL1CEuZBLMJW2Awfmd7lC9bYNyA4q/FU+OJS39J57A02jOdgGofNaw
3uGb74jrZHLRnLWvbck8ifyJlIKHuTCi7wWeS1L2EhgDu3f7CrEvRf4X4ykyIKyO5cfra7lDCj5E
au6ZZGqmrrLVQWIm+eDrqS8/qh/9V4AzluT0ITqUOkkTkPWH5nZ+oHFpi9uek3tKtRntinKAvTa3
Z+sDd/ad/zmYyPn67Ap4LF67vVcn/O0dI5tudslUfVp7hW6CwAv/hGZzhtTQOUYq97VQZKM1Fmi3
92WWtcEOZaXnz1KU6NaJ6ES+Tx+/Y5ZC62p+0IDbLhVOJaQKVAGv+KhnY/N0mMu4aw2Z2PN5bmCa
x2R6Jn3caHxpi/7zaglsrw7rnVNnUpXKqth0pHwFoLLZy/fJJ2VqnvomgD0RPzJ2sXtI9qxo9u3f
1Ihrpiw98+ZwNyng3Beh9oKU3wLHkf7OXCYs2lXLXNr5QnlfpgRRqaqGtW6OKnjGAxUgI8g2yXv0
jyy/F0BnR3Xp9/+VqSiaao+JFEHyTFuhyKIFjQ6ETrQguRJTxK+NWoA9ZvRWM3fuhZtqT3vpuzb5
NxecuobTMF2PpzbkqE9t+Equd2bNcYFXEMpt7sgdMr8GPDUPg7SAmtVjWceJk83E/tU4aJz+/mZ7
Z2ASR9P+JMDQRUY1WNGzEomnplx8mHjmrIYm+RLUw6U0eyA/WBMgHxHJpU1MMPyuKLF5WoiUeyPJ
2N83ciqkU71shqEH6LPhABs4z7SyVkBBoYH2l2KTER18yhuul+N9PFnmKDdF0JHUeWjFvCZQgjEt
RTIZ9seaXasjfLaLdSV0KaaGEOwefTMw7ZZW25CR9y0s8wunu4/idDZCZXOqJoVUpmZM2runH3jh
TPzwpPvo5a70uCHGPJLKgXXOCrvJhVtEOwSxOvs9i2NBDLSENfXKdIDSallsks6czyGQoZVJtVHS
1wCbpGymXhpeyaC1tCw82D+yszpeIuLLek9KjovMMA/HibCgkWl/FLlYq79NQ1doAxG0MONQgV2q
PP6GWh+es5m1C2tWvqWFuRYmYEGSx0YLDiwQs+DtckZOpGqeyat+h3Q/fW+s4XlzDLUhgazbrLS5
gHpp12I8yLQvEciEXSrvh2nZD5qbQWpI/qNU5PuRJZOYSKt4HbrFuEMB8b34eR336u9shlc5lrsO
ts+I0ALqr6IaGHA2a20bNkflqqogb8D8C2rel3CwQSGqj5G1eZop7TITSIceAd148TZBK9jbSpsB
0YzmFWTt5YgGQBhHC9kF5wuFINlxm7E2zcMdTufWFFV/B0vV4oQa96Dzl6f6dtJ29L44WMlqxjgp
kia3QEbtN6BEs6HCwxcVkQEckB0C1doTcpOGhZLxzL1OOTlUCVJQAi1afGAMjAcq8MCuvTC/LA9a
1F4/h7nw5cDIwCVfmxmU1HyfDVJSoumXVH/BbvNSi20x/0BGBPu54PzG0J1WK88uA0UeX88UwRzx
kPciIqpVv6uD6iZGyD6nvO0EC9DzyOqgrSQyjh12yo3XwNfLbAJ9Qg2WE5kceWU/AsaeEvwXXPaC
KaSohcJrQF/SqoSWPJM5MY4H4PgdIEFu7CzTQJKh65HxZm166HK5muiA05nKJC5A8F4djxQT98IA
u6aCsfisud3Cr3su/f2ndofdtJckScZ1VeJmClKUHc1NGZNoFLx9uRJ8Iq9XoVYYQioBGQJMPyjD
JEBwIy7pTaopFDw1nIpfItDKj2vI6gk2N8ZHMyfpCVMwV+T8vSZXl/Tglnmt4OxLJ24v2zxTMhDv
EPVu7UqT2XJivK88PHi5LLvcTgsmOAnSChJAah55t3Cy9PhSfllmI1aZ0uJt9XNZ/elHUPchycTQ
nMGc4nW4EUY6OOa9bQIuMqDVp048gLMfQI5jdBwIkruf8FXCwp6NntndYIZ2bq0+5EWoyjTq7eZl
4k8Eoaaeior8KKnZ4qfogbnnxFBVxjfNK7m2QBKty/vytm4vAfVDcrct1yzxvGjhYZN0oI4er1zp
+qiqCjGYYPto0TdAQ5pf6BZNgUzNWBNCqPj3DMkSE7bK05xnWLqjmdez2CpWlkjTs1rZBXlQYvik
fPjjD9ktMuUStVY4zJfxliy7PzGKzu2BYMuVX+Nk+BBum93JsbkTd1wcsbIRb1WD6DWZfx8I82EY
VHvrasGpaE39ujkjEDrc9deCuZFp46mun0rXX7E2WsxFUFVJ/RaZrt2JmHcpZYe/BsjaqhNM+G6U
tumdhCYNgbOYtAN18uhsOremulQ3q8ZJUbmFkQ5cSfeRvCQu3E954qy25oWsy9cyNo0EdzMZcH6n
qO77MAFYMrdzXBKEsq7SWrkwrewjJYNxh6Rn/NZ2Qh9BUwoI0e6vATAuS5UWKKaFiaHworR0jpc/
Qu3ZhVKFZ+vAYepctNfF3NII64YwI5/nLZL0Hu8vAHm6aFEEglRJCJ9jecxbf9d3XAe7RX0VyN9f
YtlVdZO7EWpB7H0XA75PmyyA5+7BZUZCAeNtdZa+TZVl/EbVsl3h7/Rb6GOCJsx1Vyfd0sVQZBzA
eREmKWeNa5sIEkOasSkkPAJmiSfGd28OUBF7pveWzgqefGMogwDmTAe4dFkcJtCRvTn3OUOqSWET
b0tTAeosZLXwPozqE6UQFzio8NuhDouRRp9JZCusMOtww0NrddzeKryxE99V2dAcWjeohFY3w56z
aDsOiYRPZpzhT+ba6ZAxgWXLA3kHXuS97tG+9qjn3zh1b8js5kJ72uiNXE7FgGvtPNcnygqJJKrd
BYlfl6smCFoa5bqNxN0xw/Jq9X5c6atMqz79aNk9EqglH+8q3ba/K4UvFrSU8+mS6/C3tPhmUV5x
WshJsDOw5Pv+s2bakPMm3BYAXietFF6zSPgc/8DBJFne+/Ebq/w0BBCfbE7mtomlXBHqr8na8/5h
+TtE0mi2TnTn3rxtOfPbCfDZveZeaxwJj7EQWzWs+BD1hlbWVswfRNKC+DdxWP+MTQ62OF6G2bpw
/rHiSTDzXDFFTq7DY6uWPrsJNWIMDNdzbMDFWJQXQ7Tn5jKFCVmdRjx6a+CSC2o0lMF+l0XOdljJ
ArKcbbbG8w5DHLBjpDMXl7ce5HiABqJqMKjNmNQ2LZ/fMgLE/ppfBF6EiqPSZc6acRHEcyaHKg/s
13VxPhPmbivnmOsR13yiHZzo/USlPcy/kx/osGDRRqnVHefd12qad7b6cQfbIiW+LZ5kPLix52IG
Q3ZXJSBHJMrSOQoILKFce1mXGCBHdkOKWrrCzpklFzcfZjo6Ymuh83IkIvfBtv8jaXswOqeu0YEy
+0AAyWcXDpDFftLbQJAstlog4Ov/0hW06OmpQPHap79CPlGJQ1jYh0PDR/+UZk+XFLyEVyGhtDgm
b0wYBz6o1vOEL4yvPnHRIVu37G2J3C2WDLYnPqM2olafnAJhgtCDa/9ytJvrB4Gu1KiijioiZnKX
2XfkN2uox41Oi+Ms1h+bp27kYfPDVBnjwkWtulQWaDxph92RG7/encff2oK/E/0WhCRJVILzouxJ
/byI5qRPktJMGbluqTtYronng94TWnNG08fWmk2P/EERa+vU1LSiO4Whif1jA7D93ScDKOoGsOW7
dtBpwrNUeHJo/CgRCArGqKsNQbUmx8ljljyCuaLEr+9Kyrg4H26GUUDqtdSZNOjZiUIvX/nu/0G2
5RpoN/F4wgmdnPulj2k0jv3Gz4eLts6JlQrt49VIuivFEDN1p91FRhiQQ8OeLJZh1z85AQFzD/81
Sb1BQfok2fDxl5JTm1wNJ8icneBLkCzVuP6S+psuPdT95YnO2nniOS39uqMNmQdmTQkOqA0CMTvf
m7DnudxhOe9qCI2cRhwwKdczaSSdgCjCMV0wbUBJmB4do0CNpN071a3++bMH6jc3F1omHRCWjwie
WflwKKHBs4ejTMTptZuZCuU3XUpzAhdi3KqA4xgc7G4U661qoOcyO7AzmY6KtD/3j3WBDjSWJOL2
GjhNORiyUjgGm5OsKi7DDzIfSeB7rBkVLBrZ/Ys3Z7/chC/A5KD5EQ0wN1o0He5lmWcwJ7TyK6l5
XH0kgQ0s8ijL+AqCdnP41WccM+zLx9Km0MVO6EvZ17tHaC4ANMvVgT9rPjrhb+8mZqPcVAQdNp4f
V/KFd4ZWkL5naLWzb91y6mwerLcAkDT/L6GzPz8yUnj+e72GLQDEe21Y70LB/kSuA2fuA30Wa64m
9S8JFxJbt0j2f8ZzZAbUU3zunSJokqogk8UtX0x2M5m+2CJb9dPE3EHtQF1b+ZcIO6+V/ZWFkwBa
Na8pjEpdezhwsEwweABZPThGRSS9APAW4PCDNH2vl2LkqpMeWDfpnzZqTGorsKkhclW966wNywHs
w0zzEQYj+tFeUr1s1g595cjQuD881Yvh6L2PcuJLHqWWqyj19UQK22cSg7HSzxpOKikBw1MTJ1CW
ifGWcJFKlvowbOfd/luMv/YdyolB15A8x3HPs0aukkxx1hujAR5608wy/OV93DYoYALaYP7Me2zt
iIjcWB0XPSiP18AtFx3WoXstAo7+ag2BSme9D6wGlxh5nRHfnXysXqp5mhtYNX72NkZjvRSJWsz6
smWMUfCtANikvxrUljs+xEVHBkWEXepp9VV8tJlAXEzqSlcTQ0seFWTnCI+dubbpWEZazNVktuV/
jJqETcEvvdbXotpEm7f24guKvbaDsLeFQC2UtLSBxdgA4fRVkSZq7do4WYJgGHFCEg7UOnXd0A3W
X0JFUsRjd/1YUiRqgIz3UoIVqJI1Xwq6oJIStaTonYI+R/C6RBr7dZBBSdb6f4jcZtjoRTg8WIuC
KXKTnYrfw6+UAcgEIkW/+gGl7P4630VqP2TLYV1IEZlU9xZ6kgVv+qByygSym5Q2cf3UJ+tZnEQK
jkQqh0ByyuUg68oTB778HDm5ICsD4sQ8thYE/KIO56dAs5FL/wmpE83d2DSgJkbG7nCCpXTw6/5O
GwmUnqCtfSUEgE6OnD9uBzokrgGr6bufMrJlc17Io5Z/rW3MxWfx6aryJIHYcZMo/0x7WcPq9ViB
+eJObERloDPc5z30zZ06i5oSbpx9TffrLlvoqOgOvPt87rcP/6QL0d7HSzAHSnAUFpWIHebjt8iq
+UH3W1RGUAIlL32D0RCVbrS1l0Rk7g5qTBdwXya7tM71TWuNiCvnJdUWohOkK+CgwcItPrSbYrEL
1vwTmfzN/hXb8COu5zyJjydXxcFijJYDJnDHfQXQxxiKfjmW6D5gcA9W94NhSz/+pxWnDl7QvWhk
9YFucitHLcgh7YRgfCSlHVTYa1+XW0oUXf7Yofk4l7a4PUon1mtmtjvUrTzzw2Z56FFfxg9KI8CN
xvfCBHdJBLUfPSAfcUF+isi5QbiHwVxEgyibE/ekrVOJ+3b57BkJspaFuvoCaGhyo9m9ixESFDNx
b0MttmEl1ecNpqHs6AxUDgiWC7RaBn6Vyqy8JADria/BeMTHEZz8O/G8Ma8blmMt52nfKuAkl8VG
u/a+phE5V4b+2hrEhPVGAMM7Bt+A1tVAb9+7U4prziPfFMGigZGIHwBXN4UaFGHgGRX29A7Dy2kw
6c9WWAJnQMU0ib7YN/3R5U4tydG+cvdYE2u8y9bx+eqDbxARxg38pG5FD6WLzP/NPSqaGsQ9Gela
6NJNGYXZrg0kB4QK+c+xgrIs6npO85QhF0BHwNILXQyYKPbCT7zFhZJ9ogIQn01oG2ZPGRNsyLGX
yu/fPsYXxv2VktTx0b/46b8cJzaHx7Q35jw9+OuOemTEtgF1AadER0vRPHqDzf7ie7n8oshF/z3q
tjeofga7HlUybA6TLypsJfUF4oqS7H6a7cALG/GJCFNHNUolbqDKfDvlEYGF/UxJg7OC3gL6l50H
/VB/iSWvzXrnYTuxaOp8192SojwV+LwUkUicLD6KioJM/pcYyLasYhymnCK6o4lsON/UCOW2mJJu
Qbrbr+/Cxv9emM6jIoC7mCvpKX+uGgZORUAIUk+l+omYg09p8EZ6oQnEJQmNCor2mXuxU1zHAD+D
Jc55sbWe4ssM4/7iPvE6ftiMI/7QxpD+HsYIHHYJZJv8YWEji9q2G757tjFM5Evdhcp7HnVb5uyK
nQIf11ujseZVABD8c+HN5bmPxnlrKRh0CzVFhnjYgC1h1m0gCNLNZQYSLLP8ic+eBMgNd1Z5zi6H
nTM8i/r8+ozpEhTRZakWeizoY5iY3phvsptAjt82h9PU24c7hB+0IwOhz2d3santxf8MK9pFSn3W
G3JLTqqR+Ia19/bb3APJmC9uEB7FhSBgrR0QseSyhZG8tWcWmbMlf/sSOoN59/oQCLv3misVkrF9
ZJFugZi/w3P4COUKLF1WSBydoIKbLBWV226PKkeDSJMfd5PaVV8UJ5SJcGopTGmfZX4iF1/kbVme
V2UCJLWpz3UWK4/SWuJ0qfT3Eij2sDyJnKxpK+C75QTR1e4psq3wNeHmZPNks1IU2L44KeZqRLM3
XBqmZWXHm4ddgO6aH4/byDsZdx9ZR1Vyuv0CAAKPt2oiaNwosHLTnZGaI+48n2RM7mD9fMOZAbb3
Uu1sxYv05Q/HAotbwFXyKNwyvqmZbSCiKUgJWJfeZuTjZ5CqkpNCDXBadc8Y+AGJZidMTWWyAZuQ
8dcyL3Iy5lHgCiZ6GnshwViygLHTOcknQizkBsWVzuHLedmckWTK4rLznlHArmVe8I2pyOQbrHX4
ZtbaMQOpt9uHXYoDBGcU4Ol8r2dKwhkz5fxeWBKVluYlN80och8svHRqA2mCBJou2VeKW04ak2TL
yTIAYPyYRlR3nzHL5MjkVu/gpTK8LMlSF2a7HCDTrGpO96hEyvibvd5rGB7Zdm+YZzkYQU4VGCRh
o4gnKsyn39sScLio/zUVNaFKXGnCFe5gNvN7zFARJmhZPSklh4WnWpbcAsoky/VQBWoqn7xGyNSj
a31FM9rfJzntMBIomGX4S7UFfBgXeJFp1FzBaZGniEnveqI7h+RiBThx3pE/FQ1QNO9o4KQy3dmH
HwNNaKgwy0J5tc92+fH6je0TKfbi0EEVphfGGtL45AIDTb8XIIBnJIqLpw9URKcMvUrcVUEP5QFz
DVDSk9DYy1VdR+82Qko/jrIWaUtXlt9jgyUFjIVi4TKxEsD25hamIoxCOMD8L0aLaOUifCQEVbSA
xrspkVyc+DJAxEQ9+8iIStotSSP3cEawmdJiKcYMcmsUA+3jQvH202KjVLKmNe2GFZMyvtb6ryou
DBrg26cP5ge5MCeVzgaxjxYhUMuUUIjYHFe3b4K2Eec2Gj8GVbH7myFR+enARoRQIcqQIX7HceCa
hki96vkKDOLLeRmCYn1CPDMEWQG6R1RxySoDMwd1pGV3bPi1nq8dD3cAZIk+wgsm+bkiRsitXYyH
Y6zb2o6sdoRvmmlmIELT51x1xu3SGj9xHEwCSFRsROCLwNJMfZUeLoMGleueJbivkvYQTPtxIgvD
/XxESXqmMh5bFY1fptgMpQU8AF2w561Fmjp11sQkM73xuVdkisfGDGxsO3IE3JK+zEvDuBYaoZCL
xfuI5zeXzvI/8rcJm3YsZ2tFCUpwJz5CV2jgardh6Vn6rqDUMG5RDMe8sD3MhSGQAxnf0CsivwNB
Z7tcvwK/h8l2qyARV/e3vBdjtkJH7B1wTUTxKhFmxOpli+qS8wA/lAyoeMIJPTLhcR6Pi4lFE02l
jP+HIEMzQrz1D0fDCDqBDaUhSBjTcExGVHV7RponE8P2XtB83BBWfb6mv5rAkIGe7y05qHdAn2QA
P2QKb6mr/09sTexs4pbrxAmCnFbsjjfutuK+QSbdmzNhJiaa4wXYSIs4h+qsjb1JIzM+jDeqp9D+
foGG/VOOLZsYV3TZ1idWW27ATTeTE7bgkwzvTj3/JgA1dkk7m05N03gvIIfMng5VHr3WBJ4l8aTf
/h7NdUmbyLSI/yOE2Q1Flq7MxLeJzM+4+1Wf+hMYu/CdwO7XiLe0qXv/vbFH/GQ//GRjkb2lBF2i
QF1JDUoZ/jPj1hzeLU3KmtHOV4lBtdwCORhLR0qAyYtdvTIzuT6Dp6i7L1LmMenZWhjqw4mj7NYI
34Z395WaJmYm0xZJemuhbVHLoTO64QIMoD8bYFxlh0XDchzDtnFqpZU4f8OkcTAfm7yTaKarYkap
sNd+65RnwM2vGw/ock3W5KiNmDVEEZm00dDEYQhND4G/m2dTCoLckg9NuhyyLluovQwLMFy4PGyY
vSOHpVvSUMvkZ3OExqm77vlJXn/4Cjf0LAD1jvjnx3edtTHuMtmT3DKF1nJRmDW8hLVzm91/ut+5
+8KipqE8lkUMqfDseoKY5Bfu9DHsx9ROC8kGgAXDSMzlYh19qij/I+YwOGyLJJYzknX5WVl/lqbY
Ht8dw0XZe2R4scOA1g2IDVAVQyYI35XZcPCu+U8ziuGiKoKcNNZVzzY0xM9f7uhHvv3d0S1l2NQn
09ddGo7FH6trjUZoiCM3jOAeN0nc4dC5GRp7igELWOGb1l/oWjNeTU6AT1HwEfeE1huBMWJitpfz
om74dY1VQgLpY7O31lwHj8QVBjLZqsIe7Kgb1EENSw0BcvENFXtgFhcmp3QCNbFVgi865bL/vTOJ
MQVLSfX2u8usntSdTwoL614fJGuBhz2ljSQhpOY4JZ5MRqavM+1DTtreKZmZDTvXqv8rYmnBzmHR
+Q3is3qcMs3zontacLUrwud8//RoOyPNe8PNB9vg1d6BMbSq/KcRJn9ilWJs8YXykhGJK0mBBgZl
IqFP8ynSvrm8GAN+3yCbplrMfmGDbzzlfJxfb6L9xslvOYNtibWrVEpO5A5Yi4LvgZ67jLGg8u10
YGhGUQnPpxANgaRFxyBpXgZCzeorMyvJZhPO6dcdPA8qT5Nm/5NPF6LnXuNXL+usQvhipHC4nkwn
R9WSNrRbg85X7LsT4+pICyITPaxNLcfvh8VAp31EYKJk1V9XwyaeLcsEWgkfBQcusnx/HJAIRDRP
6yjPB9aoeKAJ34T7u330iexo49L/3vtrR6Ev124mGlWsfaxOPxIO852ukoDEj4P9TraeHp8au4qI
rv1UwuM8aAa9I/ip3SWQIiuwBXNt5shk6DF9pI44cCUOR/rDDo8m3fL4xbfVAva3LeYlp5blcc8b
oxMq7sYjA8Lm/8gcT/5dzMDoaYivZteE+xSz1YGUpLBsBmO6JfWHyVK/yZIZ/ewEoLxN+w52LI1s
FRSSH/IHOrluiTGCAdNbVrFlXi7mnCIh0bxIM7P7J0QupxfxbidkDQRUYetToI2qTMEZiUqosFEf
mKTu50HmrEZoaxpb376Rb4qF93nTigMYO2Z3XpPh6ZuHmQxugXDKUsUM7Nr89fxVm8Wdmc3t+7EM
LpGVvb8XDEvAN0tVH5dwvuTZwBMW7E1v/mmtaIuvZzDO96L2ROEwAshQZ/YysIxHNtppDNupIniX
lNsWjOWhZ/z+k3etDqSanzOrjSJET3yZ5pk82HVTZucNa1ZcqBRiXGULeTjwIpfr1SSmT0VaRygD
/S1XZtXVt43amLUawFzEGv/6VslEd8Jdi3353hNDfaQAjC/a4SwUpk5/Sl42CXyzAcUH0sLrZxI4
qtogbtEQBJ4Hl7/1zoga1ehN6Ghv7DB6ovSi4WcrAwPwHjojVPef77NH0DRFf2BBkychmv3+Gw22
Z7hsvnjfMR/7gr1Ef3n7eBXcCFEWtVvxQQ0hz6NOcivC5d4Ba4PBiiFydcHkgZTyVOoRiQKrtDpc
hbEUyNPe7jEQtx3OX3qafsiObAT2vswOp3rXVmNIP99Vs+Rxg/cxYcuwjNcw8lMiY7JCd5KDMAUH
pyUrVXCT1CMD836HuVfy4ELhDKUI2u1JnVrX4Cj3T7pah5cI+WnCfGFIVM6zFgf/JS7c9g8g/2QG
t95unAj1M8Ah/S5N+8wN217fa76023kfDur0jmAfWYkfBaSUv9bIfJczKpCetG7IM5Oz255EPdOT
VvMm4I+o1VdiCul4hI6VZ4xb/3IfGufPTgepJr06SnooaD3OrqK2MsH8wyIfiXypWqRId/Nop33t
0wrF5YnADNFTk128kjvtZ5NcnqZA371Ny1y9Qe2MkSQZUslDLB9AZnD9ptxUsQBNS4CB8C/kGYNA
E2e0qTuSA/TB8gTt1xElvXc/7tb/hrixQyUB5NuyKBTaUI75ELyBAD0Tt1cHs5iZpXP4fc84R0Ou
q9LfTsIDaE2HW10b+UoHW5Cy2NZlweu9Y4iGLMNyltMyJAu7yx98+xji1S76UladcWo/rRgNldUV
K5qM76y/GDf/FUr8sBOzLdGFTt3dQWCrQz1yFARBbI+6vMlLRG8KgFPyRDqGMgTOBNwtoO5YS/qO
1JPAYBspy/+zUgZjPjBfYZEb4GTIT304nTSuNr77QpbAgo26fi/b0/lSPe2RswoXIWizg878PJdM
piMb2Iac6H00GRsxx70pyudC2MavX10Oq7zxLfzYwDxZEzpqkRZA4nTWJXiiyLGE2+OKnzOJ2vVA
KawsBd2rAKZy1x+y/8DX2pz0Wls9t86/fGviOoXAR2bwGbKsOm8U6I2AvzGV6HCO1uEZIASfNkj2
9ovzXMJD+7WJziGtYiJCIQUK7c5GduVW9wuql1nou06bKno77gzFD8tYUY+ZrytDA6cctL0cbWyU
dq+dQNPH8Y1LXJw9SqK/cJoztpNg5aBYW3DkLYtso9a/njKHi+0uuai4msLl5j7u5C55HZ7YrMQ7
2FnrrLQnXRjxHNPM1wsVxVRfS3n2FyujPRud9E2ykUinAKAmXy0lBtnqX5mVSkCDHCBWXEMOHmaM
rikYf/vdms5HWh5w6qcaQIiOce1HSfRjtUvlGzKRqbIXNohdjCxvy/MkHOoQVmFCr2UIiAjow39g
k/uUtQrXaMxWdGsFy8xmo35bnf7Kqf+ipKE0QPiHCj+9SyC1vOyZNmXkx2RgMgOGK507xwB3r4Be
/SCCmurIwl8nN+1xn/27XQDW64UCL3kOcHg6ATW2cM/p5Sn+eDiFBXAFYAkbJNc8H8/8SH16AyqS
8uWjxVbPrrZI+s2upQKwWn82KlHDsVe+pAPSnT0PpP5pi3PYc7y3vfQ8waCz0YcEfWHo+bDRI0J8
SHPiDz6lC46udMsfdxiI9yvsPLhtuNRK+vwiZif23L+Ntmv0dDB4o/dWd1T3hLrw6ZQgqruSyTlt
ly+ovzNXATGZrs0Ztp83MNYzRPKNYbxdyGUXOaP9x+FL1qFp4V2/wPSE5lS71p9ix9uHHFtomY5w
FV2foTd2p65+8Px1/tXINdzk2wLVliDHqHSWeMJ9hhjRRwpHCk6f+6KJF53NfrpFmdaKHbV9NXEw
CWgwlCWM642w9gucbKc7uj2p1/cIBnSMwyrN3Zz2SYIpM9gsKzSbJbCgEDmRfWu8lPCiWNb3uAKl
+rmYzlOHAhdeZEYbHCp6t7gaDx/IxrQgSXY5SW1H020Z3/8JDTzrrd1DNMHVHr5n2SrP+1MQXCpq
38imbCyNK2uiooeCok7J+WWWcgnIpvRqJ7lHpzV6toMEvUtL+AFRKHIuXtzd2CEUhoJWDkcPK8t1
iLGFHWmkMpVr5CsN4gde+GjQ0gHAw7PJoHAqMXeVYE5vIV24XHiNq+BLjP5k1qXiZ7iryzyBLbgi
CpmiwAZVhdYyNnJRinrSRt/DTbvOyNinSYBAPbkCnTMGElcyy1DM6J0mJwVxcnBsEkTihRtXa6pc
n+KnoF1h9NTAXvCzLhJIZt/4nt7uBr1CfTnuLAhEhjcMuQQXpF+nxz2VXdYIygq8azhYdvVI+KyK
n9YutM81AJ2pPDU+A9jXNUQYGMBl21vXc1mQKt7UcKo0ee5QLeoi2xro0X950K9Hh6Dm816vdGEj
t71RKoPYRS0FAc9HtRagiBgKT4T7emqLARHGRaxif5AoVKQB03pDCcGB7Hsz1LrI+XUU+kGXI3eK
rHoAEjOnqaJjbebEGh14Rk7kdKZI3lepf2S9SadS0V0LMHQFB2LEbfaXenXl9CbvDblExYr03VWS
ahnG+TM0qEugAXZqq1P0FAKR2PHoA5MPcHdnpQh/kuG1EKGY4QLatGYyVXdVqAVYH7wMAH/P1BR3
gELExdsKh4g1zQe4lQPotth/qekqrfzrIkPNsZOBmAsFCLT/Kyaa4BIAWjMyQlRFg9/77NUnlVcI
sR4wFo40KWFPclwKZ1/gUQU0Mcud3rFSqyX43TBMeyVDgQpj/ZK/YTYZi6+k1wiek9yyEUGDFpOl
MGOa2R9H131Ylsl+EiYBMfTR4CIDjR4br1EnlJTr+5yR4iizRZ0O1c68l1azf6uppFoSKS9ToEiU
zvKkR81cduQ5hdrCf+O9q47tmOpY9tVKc2GVPGEZYStnGgsiD6bn6D9qMJN7LpOd3/v3dUngTqhw
DtHSSMus30EnqGFUQFORZqOVXVhNO0LtWwJPPrHJgFdaUAarVQWogIHAP/8z1YNjKZSIaQhk7tBU
ISzXoJJ4HrJLrJrWAOAopTOViLUb7SvB5bGugOK5EF+AJsTHlwyp8F3IX3lsJliUp1eRROmSBMWb
4rc0zV1+tIZ5z7vfz6ukQdz2aamy87BEh574Pa26WBxRVYc6KDR1LFRXZbbUGgtMN3ERp++fdPWO
O03KEJVxf+CblleionHje+6Wvtqx+atYQNcFHDmhjhpu2O3fjj2qkHEhvmO/paNENE6OKuvWWh7G
+ojQQ0R4JeFjMOKPevljrvYA8yBQ88w+gqpzghcFOSdmgvFI+4e/Wqd+Opw9xXQ+4ACcY6vFoaMB
2eSKv9/Le3Fow9oBZPLJ+vqk92OZsbHToWSjlRrBo2xCGLOIwVhpfjDvfPL8eKzx9Fnkg788aehn
GXmzphSaRuVHreuQKNEtfXDlZ/FuL5lGgxo6y8/aFLVyr7j7ku+X76xF2Ybz7FT8v5JahwErMEV2
UVxE6zzHFE5dg8ANZjLVJlbexpk109UJs1GiAGINbmDS77ILIB7DdYgaWB+oZoveCZ0bIjBkC1v4
S1KX56RDNm/DyUZ5vqiezQpqOr6KBlVZ2uwtDgnwp1nDkt0Jfvgv7c5+EXEkDNsDyQU5WvjgCR6I
WW/7py29uh+JglNgvYU5AcxBaBbiEt/eMbqpFEwu4zgcH6oES8UmeGhcqNc2nwRekRI8HYzUT0ET
xly9bC7//QFvfXl8wHwwCWuO6fIOdhS2T52EuhmeXYP5wrIhlYzZJNdRVgQvQpVwbHpPw8pq6FfV
VTkFAT8PSNNFkmp9Cx7mhP7LtN+L3J+MtXi1JnYDt/FhiGq5Fk2A/HqXwBE9XR38Q+ZfdWH15BDO
L/yVmBbuGkAs6fZkNWzIlChxnw2mHMzDfzEja14wV9p57yRnKbUWh2AkQjQ3RO6IQbJotaWOfEO7
lNY8dr5jvKi2VfyTCwiL3MPcklgCM4TuWZYWqIDgrdXdRZgKeUXdDHSOFNSjXj46ejnT4KcfqTu+
H4aSzRqn2ImJGVTnYuBJ6iCsj0xgsYcGjkeAU8SnNTX2fLZ+51lakOV75KPsxV9VvuRt9z2VusS5
Af1LGc43dnu8GQXRnksV52f67snIN19jGOkDOU0cJ6p+3lhzA+VKeyByTa24lqQRjAIK8rbSnp1S
x7wvardr0mIKSeNunjCm2WcNxYyyFn46B1sGpCQxl8rcvtSMn/thT6dyta1K/zb7JWkNEK9OYxxs
z125TeWmoeYJN7uJCEdqH5mCnqpSPTKPFchWBTSqcjz1C/3VMgzuA651Yc4t+GS4leg4FutSPFpy
TAVADQHEJLTNkDenPB8qaYgtebr53ET0sSSvyRSpw8BJ1mhh8+gtxdIE1Jb3V8SYF7NQ8ayN5kT1
ESrXWSxzpR6uoDlyElsaPKblxz1MFAVTGm3BpbGzckxdOm21EUkIUBPPP6yBKNVzLW7zMjg+oYfA
vvQuy/9yJ3foj2zB0KqRLTlAqCVMfk7jknQ9V1HtvTt+qGM0fKYJu0+hcj89KJcD6tdmO3dmtiBJ
DJG7bjIh5EgBDyJcDu70FzrAVZieJpQECYY+k9FJ99YmcDyNrmK5M4wFwbQPnniX8bF5hoW549vL
FdeLiW1XqrjqFGj/1NFa08qxHnsmcIIqefi1iKx9z+itnYv4BvOHAQWG6mPCi8ySf6ffq+Q5m11O
CD5HGc68d2f20aGe+1OGfOJt43QM2jHeze7E6g3bHtnz6cLm+Xdxecez3tVwic2in8A3Prwx2KEk
X/zLxXLUgo9Ivf8MLdAycbcb3Nnv/8c+PNhk+Abuy3lbxlH51eZwdkSNAQLnxs1devXoFBpmrcdA
K3uUS0RFtfcA9XRpCyn23Xt7q0Ec4k4lq9b7hH/MXDmvxjuN9L4t0ig3C5rTwk3BUGzrGza6uwY0
r4m9Qmhh3PQYmL01LJbIK2GmBUW25nPERftltvwRCJW2TT2FHmXatmTXffnoCcmE6ecHSfghCv1x
ch7ZVbuuOUgFl/JmHcXywqhbHvhhuXVnBM1zj2H2rNc3MInmMW+SgqM5m45YsSm31+lFPEsr4b7c
q4oLxeg1LVZAfVX/1nDP9WEkluKcK1VDwUghOHo/manf6HxLQxbYPoog1Y8k6C4iT6YmYIluMF7M
4ehRikgTVICiwEzaZlV6wg1YQbn8oJ3tYa3fQzek6oRkgS86UIV24wrd+CAF92h3dC3TMlpWWLw1
ig0guVZmtwYnLcFYIDdy+c1YXfnVDqQjc0xbgJut/W9pjPI+Imv62lv3p640Gz3OrxlCPGpSpkmk
LhdKG5uLGV5aSkSurZS9k3tBjqw82/PaMgli0Nle2qbJZ7sFqlNianALFlNBgmsutEeNggkr86ts
4uuTk4GTd2kpIvCoCjWrTwOlaWWC6U1m9wQ9luZ0Ps9bfTQ0Tp8xhNLp+A106cjXFcA5+nkO4RdO
EzoshhDGyOmvfh1iCG5FazOXykJDMSh1sF1dxdk7+XeRVQwQDw3/MplFyJMFrXz3JzTpGLvD1a1G
nTfnlyvBcjCCkrvr6biujrcDt+ZnMY795RC6Fk4aHmqRyF7RFzMB8j05t7V/OeyeQjWxu4g1+qbo
T8SeSmgCx9UnECqIh2SQSWiJ6Zcgda79u+djfBVK9DrTe9hY9N1TNmoYuaQwvY+8uiS+kuv7NMAK
jwLhtdf6jTqUsv9r0aDeucbJrps1P03s13w6XGJ+K0akpra0Np6pOA/Evt0oZVafgLSuK0I8Ukfb
gKud32/wlOMOsu0vhmqijs0O5YMHBmvbfs8MOIvi+mMgp1UoxVfRy4Kz8bnciWbh4KtKZ2Pm0bAu
NAT7TEGD1VPkjhrAQhQOnNwWZzjxzQzdhSPnfqbpM2A9E+wTzJZOIXVMmiELYOrU6/nwYwAZ1eDc
f3dPxpYfWzw7ljfpSFg/sbzAOIXhvERbC7liVfbk6xkM/u2UECSt2ogf3osKeY3dw2/F5Z06jALe
tjznbfvpBGULmokgMeNBHyRYDGBPtlBSDNVczPHnSkbe7h/dyqmFojahGO1vJqLg/+lCLBx03new
+RXuJtffilzoduWOcOYVy7Aju2rtDINam379WvdQobUb5IIBmT8+wpK1UMrUPqnHdkKwk8T5Db9D
8jnFT6AU+g9CjB0H2E5z6GY81h+N8wEy3q2dbmIckC/+pgtv32XKlCEraFBJWVDHR6RCzkXoRw3R
p+yuwF2OPHNOiXjm4G8xEzduDOlwkp8qMncMyo/jKggdcaSArac6WmLgVPH8d7CleEYoXocT2ZZI
XFpQJsTBtoFvSTxp20W9vc5hD2BbALV7KWZ5L4eZGv2OKdUL95Em0AxRucHaskmb+LWaL2KAZew2
PUciB+oXfItqCoEHjS3+x8IfeViM0/NLpxC0tPYlr8M7sDm7j50EosDkStg3fUfNHCQWXvf2Ahex
qc/DTJYncSl+TguDeaP+QHgvqd3uH2Vr+HBs97PMySA/Af+Ep1d1rCj5hVY7WA6+VQrz6G8bZjkR
3UgJX5lrcfIIncoD8bLF20rjWvNZx3ac0rU4fXBjCVOplVynXVsM/KMMul++90P6AX/4Gwrj2IGy
pat7TavNIdPLfpn9YjgwRgAWCCeh86kk57B/PWgqTHPOBkdRXM7KAdNwQjhpWm1J0l/phrsKD28k
aJdUhY/D3sWPWQzARdavTEbLwt9K4VcfoNME9vDm3ZKLJdYzU2hQa8zkvjWj93JhOAIFctoEuCN3
qcYvoVQHaN1SBBKnYA2g7h03k0CRw7QYCbIW/nxbaoMHQ0Fa6EOjxxIA9ZWJNgF7g7Hykq/Qvmay
lOGT3+L49CMCiwcLpsWmyiWdfht8AI7UC5kjtboIzuYPXIYQQyoZER+qAKsJuY6wrww9AU/ShoZN
XKM6NevZkr94EtlfR3tkjIt8V9TPTHhms6Q9OhUSTb4bG8OIPE5YxGxdxtPJxlMHY9HjhLuLIeL1
q7YKm/FPvTzfEd0ro/RaWWjX4iBPA0GFPWzqBk3cjOmfonrhMrPxjEh9WuViSeafFVE1/5LCvzF8
rvzJziv/XwHghD8OVuXuotQ5KJyyJmsWYIC009wu8VzHfnfm4oy/+vZ+JSjw3WXFf6ZgUv2ZNAIB
kbIXvmBtvgkE2YrMKKp9BYSYgGqP+cdX6d4uFhKt6biz5hoCe0PwN6Y/HaYZEYiSuQwRiksvGWmI
Kssa9E1pZe6Iz0LyZUugQlA02prxeJILNEpRc7v47ARQi1VjpPFT9REEe5EbZQUadS41w9NKgBFD
NVmj0HGkM4CbCAkqNJnTBT5wmubHCo6E5cO9CMQJQ6aCProJxFYDKMkVCbmOXapEIc7adzsHijMk
YVCv3/ry2ZTS73zkg1HZWm0VJDqzDjDoSfYemuMWkDq6pUGmYWeqR1kJkIFIAhccxrXQQ/NzNd8J
zAwecQULhPVj9nPj881sgyRbFa21Nqr/QDTyO3nAU657dR7ci3Ovwv1Pyn84XIyZ0RwxBSd5h/xC
zL3x3Gzezrr9WlyLxuwWtb4wVZXjICwHg8m1B/7pUUGh0JxkP2QrWupmi4wgmv3xKBmgUJXt3wXx
IXmrUCZ8vjkrwLBT+T0QPoJzpwNGID0ognKXxgiFTu4Rr7QOO91Whjck+KiBlqhO6FB4lsEBEueJ
PTknosF78AiN9X7ioXUfTx5vdFCBfwEmbaxOc8xkEOL2MPFq1vXJhGKVSHdg2f8jiP5ZzryIezGo
EBNgqBXOnqadRrNKBivdkqmx+jvvXA7Q3ztR9tbKAMXAnmqBdamitcA0CdfOvoUh458N8KFWGr4D
nQaiaLZtht2KyE1xaGynkgC15vOBoVL44YE7ckpyiRtm5E/VMXj2xaG8YOC2+pnwQGPt9TH/jPmD
k9npCMS4MP5Q+QTLGXf9fNB2b5OEo++FOhgAucZOvW9zt9cEIvzSfNSFeg1YLYg5+9YTtAjdcIU0
Z52v2J26SBwG7XuFtiTpB0eeJSSTNSnFKhKPDQKI396/ldfs4w2qknf5PSDHgjS0/iGP4ufLgvVc
3Qa6wrxT34pR/owpHcIzbIzT3kjbp810509+mWskT6cZpkI0i+byFeca0iyHVsYtBcNhNiKgASRI
s7yOGmM/fhAPI+2Kqcl/Kq7vi3m4LOxfk/7F2MuKfq9rRaTaQioDZ/ZKF8Zp4Zb9Hxh94N+UteJ1
Wa5ueCr5kUltNl3+eS8ChtmibOKnC8hb6jDwHNImzLZVu9AFdUEQiw0F7CbWhET3VIAkroJz026J
trfLYDwnPkIXpK8qwfC/wbtUxUk++rz6UTBpDIbz+eb2Zt86+Jg7JnF6G0wUmHNSbXeZ1l14YlnX
vSskQjQBqk74IFEkSCIS3mAoJKVtYb9zoJiUjAqtkYh5pbQx2CeZVUezOha6X3+3AwbL2qAy1HJu
ELE1Bed0qHwzK53nxQ7koRTzzQ8Umt1qOuD8KABoeYlWSO/WXoAk5yovAk0t3muhp0OYW5y4C0jH
IUfyR9o6l3GIbUW4ACMUcjPLSPs247cbaFRdFeVA/HMiiumYHjFjwYIa8V1uSdgS3lOSWCa/gd/m
rDqYH4IisLRfdWu8Entaiu2Y/oX46C0TA//5dYV03oINJreHnsrdPmrPV2PrhvsbkJY0WEWpYHtV
luXmZPFU2pT2C3nL/jyu49P0r9AghFPByGdee/EqyKd4dFnLN15LbZkmXs9BKNg7SlkuatyOXvaY
R0D8dUMnaUr6TYOoIktQNmR7BO9wDBwseM3TuH/p6zT4umLfQQT0BoAp4KbFbC1lyNFqJ96HN+dA
LwEhWa/shS2P/zjv2YokaMVTF0aZIwUel1FgHZRyTP365f0XnkEU0CTSh0jSq0KpWHJYCEl4xl6s
mXHagePeq8Dvu5kmGtXI9kBGeiEGetTx1T77t3OIrTRlsUyqdfSfsI1p3EqKC7vZYoFiOXrUvsqv
Xl6WMDSc76+BKxZXqOf/U+HSYtejJJnZJxSc5f1GMT/bhYlSZI5ibnE8A7FIfQF72BFv9A0fhngc
6Yw742izmepx8l3OOCfdQSA0au6W3rccZwO8bScFa8GKvMpBbZAU+O7zf4mzWEQBfD0+N7/gJyDv
hQCGI8uX+IpnSEVA8RdiRM0756B4crNmj1T9xoDHvcekVWERP6CigLC8OePxKyiO+s4o/RRuSsC0
X3ekRsoj/boGE/ZSg7/SoqvkHd4hlX/U4dvAr419HkP5vDnJ2TLp/HBC08PI4XBE6SzwhpIucVCg
AnaDwP74sJjaa3BiiWOMdkDaE0kjNqgAVtz09jGOyxEfqJa+1C9fgJxLPwMeSK4kCOyPr/qRQlii
tVsrig+LHoOB/RRwqLG0lj1/nipMKycyGCdQwLnGKsFequzgpyUba8OGSxA1bE4RQGRKr8HN750O
gyCfGrs7oZzVFX5PW5HaxxIE5In34x96V9kyC5w60i3hkjou0FKBUS5/JAzNhUhbzg38eKwYBGPZ
X1aTa/6eGpvcxuxHK73hHOyy0UquQLkVDFxZefdU48p+TvUEn9SXcA3FzoigvpO/ApkGprsxtrhn
oPg1JezEjvJkncvr6BWm9TtiEkuvs2sbH+rFWyM2p3Blw59UraDexZfgkHl01pMJb2PeZEAMGbmg
Qo/hphcl3mLUHQuqdMXfY4rx6veTLauq1HyoUEoZgL2v8I6WrE5LaCf1htPdJL/cALSIp9R2Bab7
6B9OQhteoSk9sy3Bos/1ry2FlpmoAZ5uX4r8KYyEuIBIPGS2d9/a6ipYaMrXmPsNhVfP6m3nz5OZ
2pqSlXuxLMxpdeNLYENkU8Cw2fjEBt3dgRWU0Q4hw04IsYmorkK1TBj1jZWwA4OOa9OEL+rrmeEP
WSOBpeY2S2USsoqSwsRuNo98g9J/q3CacwNfZPJcRl7TtBfpS6GmFqNcV0bvmelgWMe9r2Y1iGtl
k3+OnM151iV4PwYwg1xb/fDEg+7PU5h9rABKHcPZj7zjGIDZqwSyPGV6M/O0i6ZpjnenYlygW4t9
DD0A35JtCDV6fWPha3z37vqkV01/kFHhabzOghYnlImtYMpmoyljJN9l/P2JHDOODYX9j9gKXFkc
Nr9f340eIQd4bQJMceuU5CVbpv4C+f1VDyZXEkoWT8AXDDTqXGqfthwg8MjN1meJ3QvkSO/ks7yG
Rc1XDYpyDqefs2JplrkvuAiLKQOS7Thh3aXdyXAHxFdwcTVeZtQYHHslGSF3ZKdw52Cfio3JJLT1
212IuL8dqqEPFxcaB51TMYo6asg+V6PyHszcxhuoNNTLd6Kr6fx7WCp8WHI02PHUoqXbiLlCybt8
KI4GZmFVXp5r4eC6TKvRUA4Y1xlucLVXOLuVDFeaEdllFRqMbC0BYi9Zyyem1/TR+kJkRhytNqYr
yx5HWvC9rJWUsVHCmuItoHPezPQ4Iw/9mc/vGV2I/5YuZY54sx76zogFGwnlILAyW+jQN2l+nolh
dlsKhC1Z4WQiKTgGOq9Y75m7P6Fav7YpQrMkElhiIgYp8oRA37JzL6Ysd73TwL3Y4zPwhyZ/qznZ
mz5p5iXu3hD9S6Ib/nWiloS7BI7sAml2DuH5NcR1ZWXJtXdY/YTuY2wQRSf7bueaiRd6RsH55UIV
PDRxKJXMmrOvLa4F3+mT5OJTliKygekUhKGPEo3juiPt1ezUTLHSJs6scOh1isFZvUMeKFSNJQSR
HcWdwJM2o2BroMsr0BpepU2cNj35ZShqWozxNHsFxvVCsWivjDjPZ0wthSjtNiY2WNc/Hk2L98x8
ncKdBWP4MyrrKjmBDjpIaE8B2rlrkotply4RjHAchKTO286IZzEfM0kcpHtjUcJW/Qcy7rfdo2Pg
0H+ySieFuPzKAO0iHyNyqrg05UoLWzm5kZXco4I8zJGSDbE25mHTByOFgynBlTgrtwwKjUhh7G+b
/8K056gHV6JMKTM8ttKgDuzEw5onKvzh89IZx7O3EQpv+t2/L8UlGrGUi5YDFjvOxsTN7bgWka6I
8jbugfgScRLXGKozgcBGgXdMB21nMn0xr4QOfRr/0iebdeTtIVX0zMqSNC4rCYKYnwau1jpVBxsW
IXhtZPmCGGT/zYNW3kS7wmgtQHZQ1aZpfWyNzjCaQbDA5Y6xsO7IGXGdXHpftet3cKXz9i6PNTYc
A5S/eXInPpn0tUOJB3+kVOHK6zYlJ7el2Y91E82idHpT8Ld6MJ9VvNCNRG6oshhAvDP2gwSIbFVo
hDUq48SyW/NfDlgpM7n58q/r90W3ByPk7/jt81sHLNzAmJ2YUF3qHyw+1LQ9SXiJKC4TE2+KNWMZ
QHVSN68UjAZ0teUsdl5ssK9af3j4Alm2pmsxNBKCk2L/YO7tuCFI2iHmoY98Ca3YsghFIJZGHXpj
YMF+3dHD8J7iKtpxBPPAHfzRJAYLHFpGsj5tWwvin8vcY8s/FI+Xjvgv3erpsp6+DbplJXsP4xXw
Jvu/7nz6jLiGe9vIBxTLvvo6L7++envuhlXpABQYPYjUDVSB07f2QjFSvAZCOcFJTkhE3uoGbydM
JmrfmgmVDSlYkwfJQt2R3IkIIkEvHnzqOEfrL03o4GpC5NXkZYjC3WQ97nYyVSrrtVu7rX8ZJr48
X3jwQF/gf75Cgutvh6kIolt1QO/AF0fofsRNh1Zl6zyxkEs2Es/gLrxFjbvz/7hs1SnFeS1+t51g
EVTskYsq7Tj5yFwZop1uSd9Xk/pHffaXJ+6LiDnzh5ltopHFF1++Zi9d6iYU6dV40YC0O5Ls3O1X
LicRME9eCxm9wnnA55W3D9HWfcvP5JYSuOiNbl+/xjlP/d8bo9BLxcw3VD7bQ9HvcpxoUY00NJRa
ECXbR9FD0zH39Fqxo9V/V8y3vckaJ2Q2sJfi/YuLebEEszkAXAUQCUlSWtOYmOhgLHwmow4P/rKZ
xsMoM67JUO8uj5GNknfkqJQg13yW4PDcNZW1JZJ07z62/JzuV+MyGVz0TNnQqigHqprkHlJV24wy
cM4DbnwO2aNkuqscCq2XWK3ldgcm8S4F0xDlfta8s57nh03xJUoKNCBxiFwbV/S+BCVoeTgoe75r
kA1KmAdZHDkT2T/mUYxfaSFes5/wyBMNsvJcG1TEjd0zVMUA9YWTDglSp6y10QJyM3i5I4q+mkSl
/UMqvJcqfyldFT2GOGxNjidoRgwb1gzEDhYtlUebwmpsjMBz/AwM6csN6fbt+9VQJQmmwMbHVwRy
OA2gTrAzBtT+1Cxrmbyn4nhCVSe4BdtdLfA8mMRA13iMR/yt7n4EvR0vKlqo9kHNZdvdTMmTCiGD
ykMJO825Rrxy/5YWQL11RK0ejlD4ywy2IZ4KsZSvpmjGTWhECCQnGJNFQeoeYInC8jUtAT97zHQK
+aiM1qrxe57mjfvVWnbRy9Hpc8K6GJ1IjOdQv2LhTVLVeS70sJgntuMiVWbDEdDce7suXpohMHYZ
sW0Y9uHYALAjuk6Ca7p57RlRkuil7QdDJRHHav/gS50212vAs5rxxV0yFk/vFbz/yCugIBIFBTOK
6xlD4Dm4Q3gI2lRlPnCpgljn2LiBS1cCg1XSxPgBEubmOrwHaTHsbImMbzKNsyaZc5r9sgkTJQPT
XTm0C7RAghlrjtcQQJkHm41pf2pQY+rb3J3unrfC4fi/LjbJZ1HdFm9MbyESxDQlXsQ6h+X7irE3
KfDCZKuNkNJN+vQeVZBnxgNWmB9CnKBPTik9pzkOxDdA5LP3h1UB/yhxnkYStVwlIvKIfHa/Laov
W/rXypduMxB7xbBBeY1HmICPVDUllU8VA7rGsbmKYRgN2Lqa1yRlH7tl+UDQdZnbh87VdKOP4JW3
2Ct8GWVRfk9fOurUyfaQ35vP9hquV3RkWnH1pGqoinLUMowCIOMMyFekxBltbSjcOnL+wMCZsP+j
Sl+e82wklUvFa2h5o5UNXbDSOl0QWRE6V9JEiFRtpAfKAwQUG05O54vI0u2pGtSbJEyYLZNDQGEv
k4Gupsgw6cTmykUsLruor91lNdvjoGJG9xvc1vxNsjwomUhXq+CW6gGnF3yZujUnE4YDwIkfPlbQ
fkcfuzE148JLJo7ZNOUIGnwVXMUWtWBgGvSI5ELTC5yoTZeRpPHQkkfndtaMSxdzF//kgMiWHD7F
BG55qpVbjivhfrczli6kndR5n4OZU8ypyLwlu7SYt8tqwBefmA0LyIHH14IlKID3qUuXzIOsC4YX
lzr1oEkWZfdK88ev968lzjzPb3yiGj4G0woTYlsurjHge0el9tm6uImrs8Ttqa7fSGqVMHGeRC+4
tpIw7kTjBCHKigrKMPHjedSxVyuh1XCQz89gNqwQEyO2ldY+KON8F0aPWko82MyMPY5WUGaxny/i
GaQcW2ebFLkfzpSkvrdlDiKHxLiSi7DZ19jhunJVFM9CBKMe1RAIdDvapz8U8d2JdJsdXG5f+wjd
DJcXLDyr6cDjDuRkVhD8IHevTMH6JUj4wfhr7mu0K5eS/LhvWd2Ef8fA3oQd3uxuofdAgE/mrcHW
PRswo94atdOCLUR65o95iNwDbUUvz+4842N+Gvs17ao86ExFt30BdRfNxv4f9Nv+iExSt75aKSLK
YqrKCdjeKV9VLGNVzXJ36Nn7es6IbJkZIX7UCsmwe9e72vhwVGbsqUxFT48RQpkHG7xVZhMErbwK
1LUerbmXJ8jKevHiiAuh/OGar+5dAS++p50+xZm4hGUR7SQ4TuADfvQyv+9efGig6Iixg3A0psH6
1SqfUzGAJuAdhYqmgtdt4YyoORU4VPGCJe8rWcpm5L04uIjjnTBsKkBpqJ2G1W9+Rme/sSug32HI
856RiBAp1/PSxh9M7FqFgnOS+rrZh96JdT2Ipm6by3wi6pgLGInLVDGVVP4CLgDkiFvcp/RfBMcW
Ko6ZuZ94t9SetFL7k1irEHTThVt6xh5ESE0cGzI3phPrm4Rs/h2FkdMIyWAH4veIEIEl+BssGrmt
EUp0ZAvFxeBEpcrPO/9/qbwEkpckURj1lkxNuQ8pwkqhS0y7j4PYP6gRl+dja4C+UBIP2inn8XfO
YCV5K5eLEOmR2w5Qpifar5EpnbJ/KD0qfcCcErMZXS/SFg1vuL4OS7IMGjWQQqeHETX5bGD1Wot7
9123jM9nfN8kGw/VrQiMhVmuRXvConaXsR63rOKTIAni58Bp7/UkVYS1IomS1zioP41ImD0aR0iJ
uDVMHP9HXkIJ4urAX9ixGIv/pW21I1ckCo8rIW+zMeUk1Ayf/jkLeRTEyvMC9M67qaNRnLHkoOC9
UXVOxHXUkYZS4cGRsR8h2LxCe/0ACESp3Wfcy29fJwPBXl4jps4e4w5tX8PBwfnDWAHcs2IResIS
cIMkp9TBG8Iy7/GdmXA48JgTzfXsIo5mRvlP283AoX7GyTVzWgnyFHO1Pesc6X+/1sy0IYYPRias
evrLjV6n5g9LbN/kUAwSOfimF96d91vfqHpswvJtdcihgL+aCj4qzUfwYHQLlMuKEKPSh8N/1eiV
0hGtjyoVDb+J7VzL4U6E0t+Hh/j8/GEshZ7wEQbL6ERxhkeVyKLTBZF+E83oy6RX3VYHlLdX+vdy
kp78DSF6DME6MWyYNchxsqL/knr68+B2tflvlVkTieldkYrEhSvTTQV2rY5BpLxDWNS3GNV0MiOq
mAYDLACgQ7F8cFvsD0q/yYbJCyCWrjDMzToMV1Ux6jOgSC/g9JF2CIxHB2OxndjHK+G8w4UWmqWk
3u+vHx4CmigDk4GYDBtp44oaMDhSFdGGNk1jVGZ6bVoslNVkz2RMyCbn6oTurQkv+LdufXe0tbJH
aHNOEXtFDxOzOGmw1FHaAm16LrlntxUshnisG+sMkJL8o8UQ0+rFLlijqq2n9nM4CavzY0LcaWAy
HBCbAxApOwmJF9m/y2ZIHu6N7fedVSQTCS9iG14Cc+NuVdW3U4pGfK1DiNeSvYMS5KzGXqAHH0WE
qKGggThjsRACLk2lrj4UYcUAqYk012GmqXvEEsT0DmRxfJFqYt+NTVG2VRL8m2e6QjtB4Emb+R7/
XkGhks3jv2a3YvSTgm2VldXhXyO7TbsKRvMGWcpJmE2WouuNppVEjjKokQ3Rpx61klhxTwdnZQOz
q828oOxC47Rq4JCJYiiQf6d7CYdcv5vN9p3SQsz2K38vRtew9ekikGDFNrRbULd9NT2c/sjl1LaU
q5m8Mfmywp5MpGN8vgUnIimn4StA9fY5tCiwRu3DlG8u8YRuxaTDOtOUjd3/I3u5amcJxn81/dJy
KT3TD5gx2NedeUqtwgVateMEGbKO+CppGnCGBGy3eUa62e1I4Yz7w1WwUVQQ+aDFM9qkbJw2kTK9
B/2+6g4YBcicAtYJH03gtJOgnCAKkbRUGbkOcLHFDAAOZRumhzlJuMVfLCU/wu0KUE7nmKB1O0CO
9RDkMqR9SbANUw4mBF+BPj1P5oMXAYA8VIX4etEfSsxC1Zl5Ow3NJVWG+lX38VFoML8VvrMW8bpk
adWj0E/v2JjRayUI+ZFvxdiNMW5OzKz9txmiowxehR4P9ERajmh+wxBAJStNs75gc1ZHK6gqEkwY
1G9O7Wc3PYnJPFnVPajMc81yFxwr8CF4J0KrnsghKAt7kyvKD4WnOHLV/dziMo4klCak8tGT0J7O
sMqNVfZHMqAa3AhklQT/gxnEOR74apxGHQ5jEVoxo75OJJP/KvN8Rru1jzQ4EXUqMtUgzu3Drx9j
1zSkuG4snZuKy/TuDLW+8N8lQxPrc/ck0+fNiaUqaPs9GvjanxZVj4nmWP/IjhzR7GEEnYxN1Gnc
4jYlu8Tb1LD3zqzbXH8FDEYC8pMWinmHJFJ51heqGOQ71n0F1wnt+U0fc9uf5rVauUYJFxkXjk2v
1wxWyrvYnx/YdhfWL/JvF83klDpnrZvuVr68/9i5959fGA9Oc24jP2lCdwhm+wBkbvPN3qHRjfYe
l0lhSjRMLWH/7wbS4wLV2EMwIEjh1nTG58QF9rav1bLd3Kk3bF5MGpNSq4IiO+qh7ldnfDmZ3uVB
ttj3ZwnBrjxo2+7+WKYxmxrFRqrb2RFRHkwymmMi/E9PuYUhYiHMzlE+a9kF5xavGp+32HKTajrQ
zmMSdbpmryd+Tk2g2JaRoXiZtCgnqh6899M/oaiAzNylKJsvBydarGp5zPK0J8FPKjnsPJ+jsepn
z865SrwPkeW8u+x8AcWxbVoBm2zhKg220zvcocJI4DJbu13bBnFixqiamMV7fVnN1tfkAg9CyJHe
nrR7G1Td0MV90Di1VKbY+ndaqYvTQiOYuMW2ce0QaG/cDTdngU2zPlfPU0baBViVUr4opB9JEiqf
lv5McWImmPOlbjDoSXIeqmlUdBunjXS7vtTsYNGso9VwBQNGtez18qTnNXY8yoz4RBmV3P6pSeL2
t8++bqPf5VZnBYUup00V9ZpNDrUwLYnT6fMlPWPvKHHxpUHvG90+JCv31LLw1E1tAfvxukS0wO1f
iLiVI2typuH/gVvqPMP2dawkaRHwvaumMz6Or3bzkd7bQD+d/YSoruOYnFfOSua/5wkD2yZp/Wnx
YLn8ANmZBFmuodDhXr7uHe24FavXzRt27heBUDbZKAmokACipuBpwEDAKYCWzBrsdlacMN2+n31+
78IxsUbsSnqNVuerdX4TbzOf4B9ui1oUIjyo3RTiEJUvxMeWWxghQRy5gL21vS9+NSsTea9ksMGm
9/mJ3alk1QdK+KVHcCdv4p6bf5SuqD9jlsAEXHX/DJq+M65soq0ov7kHpycgN8q+z+QcqJipYVIq
2VRuEPNz5ZfRAANb1VEWv9OOPhj02oszd3yC5AFMhFw0dIVo+wQ6pstK5Dw+PVwUBi2coJ0HYsu4
Cu1WyCd8jmKsjsqDTUd8itmygcV4Rxizz/O/aeOhgGYyMFtjBQaQDROXX/MxMPJHOAvURhuwY9cT
vEjSYj4aT5QjX3/KT+dR4QSSNQin6+jCVc8crtPdhEnpS48IHC++RyfJPhojgmM5ne9RHtVc7TIx
z6WMonw4Qxm5hRbw5EwSeXizAS0xZtrP53PBO/6GQbwYbYwFE2P4GHIOJM+vCKobhO5aJ3VXtIWT
FszvDBBlFdWKqHMPxFxlybBXyVqm3C+CH245kbaAwzAuJUtMkLevtc5KWfzzk9nhvADWdUpIxizY
x9l/CyvEKbtkirxvoI1OY1I5nEupDCUVcfhdIV3vZzJrX+BXSVKu2devKJwKi9pK3U7/MGYwuDs5
1kZN1e9M2O9nm5Zt5REla3S8OJJP04SXTfybQcgg4ZucBK4RaR4E/kAN2AvjOcNIjcMBSmpc0dwJ
a8nJQdXJCOakOmrUASVwa3yii6hArAOq5LcY9cxjJnBg0QY+gXIhWv7sZj1eFgbs+ROlfYYjW51n
nFRjXJO7nDSKoV1FMNC9GBI2L4Kt7fEqERoPNXbJ6ZMP4+pPpw7Z+iBTN+mV+Z/v6toWdbBhYK5T
miCQ0vw21HepCzE+6zC/6wlko/TnNwK95tiOwjiDr7+q4xw9EfBOPwOBunqVHdbReOrS+6eg6DtZ
8Pp5Vd/y6fMUk3Ry2XtmAggBaNx9R41w3THylho1+XFCZa3iV7V2w47eqWM5V8bk4wbFNclXspSq
5QTKdd87GIXHs5r338FUpoZscAFTYz1Ua0v+8TLxd2x/lya4/kMhCs2C9GqGVwVrDoy4GjAQcdxx
tI28lqqs1X5AE0Izbnyy+I2tuOyP34CCKcrA2zupgA4D9DTwx2g9LVC8SchiORfFWs0qTU2pdljU
9rxu28wkoglnL2cHjL8d6SBf0B9XCP3KuWa0pH+Ok585AitDCpPFyySzAXuciijGr7DdU13k3CYh
oVOwrzyukORe05W9y9Yuf7pwoPJtJ8ZKqNtKEu3NUIiua/e9uTeL+7p/f/wnAVRMaOKfmBmsXczN
NFONoBclyAC/LtAEpYPqwruPkoGkgw77FQoSxbVOYZaBDhxfrOoqeQv6UVcUjgG0OAsnDTGIjZzc
atYSh2Jpi50I4gpOPa4rqgxgzItC3kFoUbIZfhCibp0OBa5pp+lJ9SgdkWJbcbzFBe/pKbVDjzhw
PNDQsTgZKte/hqY7Du7wiosjauk38WLF+YM3YnkPalEWMdf9sb8CMXpSNDa6KSavMIrmlEtIRkxN
3oXfgQ+XKEpkrx6gxos9ciTS9b/pL/SeAVaj1jcSKiH2yofXPJo6r2McSOoqe+5y4U4ZyY/6QbVr
uvXx4PKOCOJ90C2lVECNWFnJQJzhiu51wg53t8hhAhkPBy5GOfauzSEwW9ISVznAeq4urTFbGuEY
KpE23AKRQI0EtErPtldpR8SNAqnSy980VXu08UD9NrpnZCtM2FYcoxutpIgQ6PaFZL8c6IwE7CEm
iDv5lH7XL89OSyYlHtnDGOtAgHCxK0K8clWXF1SfXZur+VXo4W35rvSm+rhgMdYLBtE/doYMNoqz
KuLdx/+6ACshHp+tT261i8vVl4EfsEab6MW9lDMhds+SjuBZCHxAsNJTCG3C41U96+gxWwKfsEHH
7opcFiAeGue75OHN0LPgDXq1OrqzTjuXATD6ObKIe8cCuQ3jHiiraio+qzIP4u5G4BtAvvuk6MHB
icuR2dRAOg6AgYUkFQUvk0Nz7J060q1nmi+/rWOoqCkpWpuDnEw8YRhhiMm6ub2Z7fm8rDZi89xM
3CK7iLxuv43AkqyWtsUvsz79piQKTt+mYul2olUXARmnLX4ATfgeybeCeoN/qEgdMpeLq9tuWjZm
0U5orZTR26WYtlofiyfdFl+4lvChzfUz6CfccaUM6IXqp+2jta8H+mCfaZdkI6UjxjUPTR0OQxlf
mdziLe6sKKIajjwfAIAkwcCzyJJFS/oDcixRwf4j3/OW5VGd6MFZibTeKxgLCYJfD8K8vxQ5Tj6o
Q3MoEUX3vy4XH/WFGZTHxpg/zWAFakJr2O9Su9RYl45XvPxEdLifnh1+OBnEwzudpwfqSe/sxNki
vleZjhJSE2ZJ2h0Z7N4EvdaeBCQBK5AN5DUlAupL/cfYnRvrbcO2CZ4xyH7lBOgdIT25cVfjgACQ
maAlt6Ncr+Fcey2i9e4b+FYJmKSou0V1/syykA76tUwQv/ZciocYiEK5SHbD/+QVZIipOY2UHkje
1mECyIyO8GkdoHU150FfsBXYrmmIjhjYXL93AOUaiz4RlqvF5g7EI9OJUH35F4U3/7Fj9LcetJEN
BFgvY5A0MQQHduiRm6Ba/HByA8WuhODzH/g63wEhS6YNfaFGjV2KUqtYy52pSP1sfdpL9h7nmHVZ
PlJwq4J+5rfsXeuGMTG9mD1sIardtirN7simehJcZDruZCE09EZPLimOL33H2Dbwan48ygOt8DSU
hHl8YTwfd4RSVi1oE30I126wMb8JOyMLi+bLbN9IUNtDaLMw7fxIbXNuuJu2lqNzoKz/3WnRlZe2
ZmzEsOlYgIkp789HqwQ2u+EAnJx+uZ2LqjkzKD50UBAtLXze/KFzZxOeu5IxQvU910YtPXAMSxGg
St6JUQfULQEgYhSo6wNOmzAD2huHqUHTP4M3aRyCkP335dTbBzJePo05DNNhz8xcr4Z4Z8aXgS3t
4umfJ9kmrv08wXx52k+TUFAoIDlCqUZPVH/Yfj9wS2/YpSeT6X/KzrCqfMG6bW38Xc5QtynVI5/C
cBChbDfCoiF1XotsO6Gc5Ay2p+U7IGrNiUQWZLJ1ST5lJrdZWFGaLJ0VRpBHH+qHkuBgGYjWDhfN
mE+iVY8Ga3Iyo9K3mZ+z2yyvdsAfkpPjwcrv0gCihHXYVbMfWR0TBlnoCPGiA2hqwi4K6BvZGPbE
z1wNBmj7acv2r5JXc480qpYaaoQLtJDIG8WO01PKydI1ACNCZDVRLoNyZbjaWh+Jv6rf4zvmFTdy
BxDOi9oJXfv1kL5uZu6jrk6MFd8acFdXZJZkuogZMkslL9ul0SmhPVCAPeSc6okzmoYzmmyGPr2F
znWYYubckA5dzZf7hPw9wgZV1uwcU8Nr0oXJFy+nsociPPyU4+FWGpLLqmbbOUwLLgyY+wP08837
l5XUA2GtBopgABgxSfnL/WoYPKR88vnmr+gLKBK4qtZ/yGjia293KXe7JcxnvHDZEKegpg08+yKD
ucs8PhGftUt3PCV2Xv5zWY3RqnOpSo0v6nQI8EhpRciL9rgkySHFoMI2bKswHiibwcbsJvyBua4Q
6E2VT+RgkWSZDlsaktKXU+eWbbLIdt4AO3Mk3nm4+YfofDQC99VD4Hhk6rcWy0kxJj4qYtdceaoq
bm6Y0b2E+cSKEHl84I3UXMclGhOZ8tbwqWWPDm2jw6kmLx3J2I0ZeQB2Q+Z0XKXnYgEzSMHBd4sV
srlnDxbW4KlTYVhd73VCY0d9wdVH5R8yd4Y0ZScgV4i23c7fuiXfvSd2q+6IdC6KgqaMjyD1TRbu
WYmpZ16GhUvIfIuldMNTVM/g3/RnZ8453RxRin0cRYKEzmBj3tTT7TN3PeXiZrOQYsR6M4c2EOWi
EMnxnRWYRdOuFQMgYy1CKWNJJbRmaJ3F96LmCx+kaRyjr/LB/m2vplHu4Ob08t+ELiXr37YY0B/N
N4rLTew31S2P0vBY5x70sauZayj/J5Gmbct9lNWJHEmHi3a8E004YCjmFOkWUmGqNLZXBu/N+a7V
iq0iwJ/p8FemvqgGIWFgc+o1Or5I/+yzhauvlrSkbYU0UWMQhkBU5snfT0kghOkcHoN+L5ZjO5ip
LfocSZY0OcYJstTCNi9ml0y4DXudTkbm+oHCBXzF17I/enXPVMKROWycRf5EtAF5oZnF/ANnn6eH
htnaFaErNFieWG16hd/79c4bHFAbKzOdaHlkwXPR6tOs9WhxIVs6u8LrFK6UgF9aV55RK26s2jXS
aajO4bLVxQYcDUqkaOslf9y7HMInsmdZlpObqEYmfdFxurEYBuVvB/AU/lF4kzXokJp/Cwi2dEV1
Z0G+/iTYAUnEIYOE/o8E7RC95bO74pgmsWeXUe1X1Oe/FFoEpoVIhu6oiIdWJEnn0dsCcFdktb4t
8gMqCGbuSZDbuTRlK+3ikKPiageJnmA83/Nic3WWGMZC4kEc6hxlKumQ7eK9wZUDh9vQJUegQDQT
cbZyFbvGZplHFO8Tr29+x7sZhkosErC0touOSnqbXCauhLQsJOSGpnr1U8caSvUQL0I+FM0zmxyF
Pfy/4W0M1cxzhshsTK5A1gZQ6OcuX3WJikNRkwcTqYAuJh1wVHn519n6YxCr3CLk0ME/BRZAawhh
EImfjjLmRbX5gXbnNGuv2LL0+KQdb09IW1DasCkxv7zn7Z/dQGyddmLS91xuBmEcEaUgfAordKc9
C9+yXYcjmwqRQtgJmTCEaubN4Yu+kC+Kcs25bIsUmu6omfdrr9UtUWXScqcqBFEJ1YIg220K/WZa
OHaRw0Kin30bjyJr+Zi53ess/yPWTzSjvPf2THDeMOSobWtAhJS6CmYowmbZRxMclKhPdSAq+y2L
+BydvHA7JYvfjS2zJkkVz7SfbfeYw92VgQozUpqEe/kMF7oCZQONovOtD5PUiWx+QuhVKdd2bLS3
z/8qc5CWeaIsScD++EparTBC30Dvs6HTBa4Hy72GeQDcgNj8XSdBJKqZ7iAfL18Cym9Tu5zWQCyg
aXKDuqeD/vrOqA4ksgzT68ZBQENVamOYV4BCRQ8PRz5wXHwIRM8q0cq7gbv5es8Nm6KSbcrnZjau
3gbEDuP/zg69yvPhf1jlvk0esTjxCxmkFTbDbEBlvvE4WSy0i/uwrH5/WGPmWMxFGc/0ik9Q0CRh
Xs1qYmGxBnm72PQMeyEYR6qnTTKwebt4HAJOhty1uiAfL46z1rO2B2RbvOPvvaBVMAG50GhGFLWj
slkwRLCIO37rwIy3RD2K05QgOzuWHYRUZOSjX+2MOvV+N49VuMPe9osj11gWTcYbWTsPqPVw8LcT
yRfP8NuD6rubA+hzr07GVs7Ur2BRwWmBvFOq/aunHQNPDAgHdDJg6eWaiYIRuF/amCupTd6eFIVL
0Z8P+5Xm41NkZXM0r6y7BPhooQ0j8u1UlXrNfsPPTbBrDGaDaePuOYKPm6MFStWniyeqhBBA2KDW
+rccAtoRBEvrPcl4HpIci+lAOJ387Jb4w504n8I5cjTAwl999xHkK/VyxsjtUzmOmRnbjNlv6BiG
De79qMSp43VeH5iYtQRlcCbU7Zfmxjpa+8oa77H4Bkj7bxcXl66uJroRqskFyjrocLdO+sJQPCzV
aDCe3o8xN9QlLZIEHlyDQxpEoGy9DLXj62+TizL7OWaa5D1LCzIaw+MsKGMVX84XbFzbkZCn7tPh
luEKv+m+ca6Z5JWJxNT9PbzwvwGRjv/n8R8kS/2z6AOwqfHdVAus24lCtoh3Zl0S1uBISi8PIkOi
PIb1tBVSTiZKDB/uTZedYZqdfl/KazZRhJdC5R3A6owHVNhNKrkdWNS1FlYb1RNEJUNKXQxr4g7G
70Yl8k5GjVM5FDeZL+G777XeylP5SqvLqfQ1np50G9jGOG1W8vcaBYmtj53u/kIGCUOqQrxIzg2T
V5fWaFBXqFL7tnpaq3X3yFuDmEmsF34y66yml2vYRCQWxha2c8vIutE4GX887cn0aANStkSftpyA
5nfRYHYvteol2tmWWeAg86ePP7PnIMTbXTLo95AOJUw3C622SVEuDLRMNw46G7/rmQm8WcYL0QmI
HUvJJj4b/xYO8MjsUgaNdgLx1Ht9I4pSXmZCoX7Obwcgudr8lszK8sS/COQQlmlvzGJ7N4+9aq0g
75E9bkvUBIitBfIe35tk7PaR4K8eU432sJg6DMWccgaSnrI7d1qdSETOxzARZQZS2VwsR/7mYi+X
BYj17mOYGRfMWybjR9EI1X30YUOkf/Pj9nzF07qKTxx/61/x+dsnemYkuP+KQNUq2iLGd7fYBfvK
QDsElZT599AVpNXJ8d9A2b5Rg2CVvi+Csb1DmtT/UzPEoyEX99kYxIgvxRR9GpworILD8A0j9FJO
bC2o7VJC4KAyNoWOUA5tIKbqUe5df0o2BYmonn2gyHkHa4weEVVxLgKkZ6+8MUIDTm50lNpV3g7R
hmiEoIYyqQ5IJbZuGTUaW2B/ksjFs8GH6PZFaD+FAB/5qiKzttp4IMI8UrUeERRR6mb6e5wKtx1Q
YIlXlFAL4NgxMXTdhgKB9wd+vSL1i1yy/+uVqLDyxP8uqv8aXD1vX6G+JJ/Jdtk14akOGqhTvLS+
EGvfRuXj3npxXurSyvhqq107pVNVf5piWM2yb000C9x1hP/aq9uelAiH56vfLknJ7V8+eKf7mxvA
DgxjecWhh7ZJB9QOGQiXEZ5MG//XRgDT6ZWxIVtxOuW/hm+9DAeZS8s42n6VtDzsp9UDYiRymUUA
5IT+BwikOTFB9BjqjYLIKxtBB1kH5sKA4RtdcNP5Ekjxs/TA4JAgSbKoN4ybeb1OYAzgy5L/0SEc
j1VDxvy3mhSDRW9KRNcj8CMn7AAu64vmw1lPM19Pu8d5Hl4wS0s0nQLuAQV9DwcuCTvk25lEwhfm
xiuH+WqPzb0eB++Q70Q9MG1FNm/AA4Bknx3RazOTR73TMiLb+sTjSSrZGRNGttNIWy+9ieVu7L+6
ploVoqx+MCs4BZsFJeOvRJXOGGJb7GB7fE1/SjAsGEKAoFUlhW/2xdF2j1YRjFVLAYFuSObFbHDZ
3hc+Ttpoaq/nDLMNpNiPwiINzf+QZDnza+HcCCZwNI9tjcu4N94H7J2f5ew/avuLSuT/yt80pi/A
DZ8ssn/LpLklctW8mJEh113KhGP+gvvUhftht7wBr5nI4EeOrzq6ESvq/d6X4BGn0AWmgesGBsSf
wjDXQwj5acJP7ZUqjVE64lEQ4f5GowW/Ol9yq7Ojz3uKfonmIgG29AAeiWmbdJ4KQwufcAUny4+w
M0ENpFwiOQseoFgi1Iqznw/QcMI9zp+uP3tQ/Ul8SUJY6PJ/FRCWCSyN0dq/PgNIQaMBkG+JoRMW
bkM+et28n5J+gMJMevkHF6vfIDnOEHdFzqJL2NcoNA3K1tMloThobDF95g9pgA0comN+uFoAo6Nw
j7fp/+M7tLa3z3ihAK+h3EiwKAEYEJfTTiwx29AFrePKuF6Tj478OkWUguAzX1/KRTdFEHbo93Y2
SELYqr+uRAYtJ4VKqEb3yCC8WgtU0qd8OhlYSiILH+bCBGrCumfn5r2YvgDLL+KWvBZWYUAQKh7e
mDOT01dhKy8gFBrCxbhb5GdZBx2beQwkUsBJoxRJMfUG9mEko50QjoSJdmNeF23W7ehQkFCaFB9o
0jYiWy91pxgiJLO0XyHmHpCDo7iME07Pq5f0jYHoRQWfURwi16X/PK5AFb56u4esJMeUgQSV5jJY
ALY8zmRtkEbNlnsYyHbEm2TdsZZxHPeLqqkA7A+n6D9m6yQTh7NNNCEJqckFVzMdcph22lBb6PaZ
MogqTXkcAdDuwZ9hhUdVRs7S/IxGIEtSWGClYe8QFn6mJKlNgbWy2cmmsI9qQdT9WnOP0L2iFSwF
HY8y90XYlpfsCPgR9BmcAlqen0PscEWVMUCkZTSiRxi3aiscN+NikCw9hsPeDE1Aj87czH+8ZmXs
jTfBIGKdq6nIrEELbfY7qzxNBxAgJVxZwa74HyicUC1YWL1lrTADhQfqnQK5G6nsR5pVrrGt6fjF
GfR0cy8Z1PzJwQaQwqmHMrgq8HwLzo7TjqFhGVjqfYaafU4fqhKqJ23rpYFdcmbXrdmEcM1v2oap
zk5D0wP++yRPiR6tX48Wl+kGzMOzIlkkNyO3cyIk1XIEGX8QvhWhrt+0IgScKM+OD3GbCWdYHB/R
Z73qs9uXwvEwBG3HH9ZKEk8iDb3KrYeyIeMaFj3IKbV8xT3qlxhstOHuKuYiR/6TqV03XSCeMPbB
RP4DGuCv4QrRUrbkEd16eZVf/fZB+ZSw9IM4qPXmW7LRP0U5D4ozMxGAlr82Dzo1dXNPcdbquyny
rT3bXLstC5N1KMYpaLjHfYmb4v2BzZfiPGF29bP+Gufg4bdBmu6emlhbuPGD6Nmr6Jw+d2SBwA1t
DvXsK236kmmc5oSBS/uKTn9aBcGBD/k0WG8B2Jzte2Y0PBOZUiM9P3cHNqtjvzyYTbCWoV+iSGoB
z5ZN+sEz82Y9Cr1BvF4ugcY+JbqTYiicUKJy/AmODtdeqiflz2lfUxPzN3ybhnUZcIzxPSrbqle9
a71DrQrCBSVI/O1yuTLBsJlZYCG5+USLXYPhzoGg/AbFY96F0gq0A7xYzhmu3S5j1JKRHNZUYvEp
jaEYcsCYHVDJAg+TeHBSAqu0Ad2tihvGDlGfH4M5qaHoAJjm1XXmKtftEq/pgAHKhbtSpQATY3Y8
K/4BwYIGp3Cga8fQG1/EWW8JphWIikxvD+ovbGYVO0UsB5/8cWSbnTdXemv3U6gOVr6NVYtxNJbR
U37/lrUt6cqKHAkjQYHDxMb1g7xIY7EcKoPC14uhFzO1YRpCzFpkgrb416Jcu7yTaTnuaDP3oNZa
aHoD3X3oLih2/zwChoDlchiJnGvDg/6PZH/Z3jvLfthjMAJ/9oFeL14pq8zx2bJdt0uzTOajCCx/
LpIVKteE9T6XGxVZXg3MR8n7V+GgObyAdGeef0e9e32cnExM1ZfvEcwlDIrrthujwD1XU3GkyvoO
4q6+U1m3m0H/3foP9qf0K6AikxvrV/uSNKUir2VlrjaapwepZXS0v4nGzbw0vzgtQ/U75/C+xRql
/kzad8dfeWc6mX7nwaNUgFx4GxhdGFQWBMestzoXedQ15sh8Y8msDo7e0JC34F4ccSvp5pPGmSMZ
a97Qd+tyUjx/g9bJDhcsO9CmCvwqydfMEZwKdyGtl4VkytTGVymO6Yr4nQ8SLhmu4AS1CAgylwpZ
w+6Yua5VzDYKiozewbN+qI7iNPj2Yus/6X2/U2HuEZFQZYcH+U8hpxuzStmZuqj1ONJaMFm+pNbN
nZ9gmL8iSkPZlTUdxJZAVJjx8rp6Piwv2s0FOQGryujVR8JkUfP1bvlj+hPfCxbeb3PydbvJ2IDo
QElWm7KXKBEfehsQL5c6GiI5WFKIV7wUrR8X6kIYRmwfLQHnHzLbsubW1i/Nh5qTFK3SmxTdIZL8
fS4Q8ZAl0mUAu+StAOqeiNx71B+gk27f7uT6iyzYhjHiISJgUbYdIM/Nminyl/m7+5ujqGtMoKdR
17k4amSrHyJW1xCUtrZFapWrWHyn5u/r4wXCgwa2I2PbpJ1nZZoSMZ31r8a0YgUcxE6m4sOyed1u
/udpkfWXerleiQmaXXSYLWMF2P/mr/V/Xomx1+cx6J+b7rFJLXuP8bwGqnVQjfsQJ2CIut4TGW2h
C5rgKzxkjGc38LPg1TZ0z++MD4WcVSiTTGljGqkktldp4SemMX40P9QqrH+DjdjHMzHIVCkzF4Uh
GNwGwQxIWL/d/92IU7lC/Z+QmWeYcKQRf2srWE9QKMhALfEEARi9Hvr7FAVEi2Aq61Sl2igXqTUF
QOu/QClRSiZCS8bfGUJ6STnRdI7MUSxI+b+vzrfNOIRUeft7OBP/vS+6pzMI+tWJX86KIi0m3dcc
quIPwdoDOu3DsSy4Pm0f8Y4rUgB7z3ikPBCp1U+k8X2Y0aYaVogX8Lp5bp+sB6/kn0JU7VXzUbHk
PuBzM1tgpkrWFVWzsl8bW6f0vyzRMNdNCAUbD2CR/PgmT0y8kExqQCIYrVYpW/pmqL3C+vyF74xl
dv2h1w/52Tb1kTC0nDfwm6tlT5rlKF9SNqJ4rCaKgXt8HhmePvKNrLLRbdWoW9vVennIxkPdu8qS
VwTKC6eDGAcB3Djlc/kKvptrFZWqQhq5IXR0orhDHlTTtIaR9h1QJk6IvjXHj75Q+JqvSSfUpJ7N
3HTAUxIzFJbt/BNpqxDP0PFOcB3x0CvFK2zJGYX1C7kYKBUs2s0W7dgxTSgS1AfD9GhOYxBvn+4l
RBgo+FkZXdZKQF3fznukJ9RJke/p7VPvmoojKI1KDtmL8GlknleveDufl4Io3rj+das+6nPJhkW2
tsBdkmTAmfbXFzz4UVvcjmB1FpAMpwnscB2FKfhWdhvnAmSdleQLq7rt6yI/ApHnO8oPIpPhins9
PW2enBlCC/6DHkaU1KbmzU96qz0myBTa3d5rsc7mJ5nsdFWOQaQShLqX4BbNOxw0CQwHc3SDpbOa
ytrXDVUIKx+CUSOEtPbTgdrEYe5ViSDudPv1hMtt3pLq+XpNvxTFOqZWLbQulZ+jZoGdjKjizXVN
yIO7WfQnseFIIGiC9PEjmpjVuGWNQeoXF/+LfVJnNfO9fDFgv0yZdgn/iMrjFAefVphTziF78Jb/
l1l7k3Ahh/QhE3gzO35qO3gGvwhBMfdAdOuxEpFPeCWaKytFFK6YufGWVtQ9lbN3LAg1aVllf0U9
eFGaBcn8nb1bqqJ634flNbLUEnX8oaKC36wfENw5YuYoT7KoB4fIBODFDTK9hOaoJH+wdpRIZfec
Xt2ZK7lYK0qIl//lU62ZCGaWoQ1ps3GyZbx4CPA8SnjP1I4137P34WqQUD7JD2szz44ilcyeAo6F
XT2QRORriJmYyQ9Zkatm6p5IZxq59OFJuQ0SpR/BY6TEOwgOJpIkvtWGiOw0Lgslwoh+Gya+hAx2
lQ5syBdspgEuTX0yUYLdaAqFU2CrDSL0H8nmB8oh1B44l13V6c1sTvBr3UX5zTR5MCUwEJrkMydj
27ZJSOKao2/G0RW1jcRjwhcAqzfcN+Vgm9GGQu94PGGzISd40+68a2lSzyY8V2I8TB0r2qk1pEM2
PZP0x9shsa+qtteq/bFmEusBXNjg2019SmxbPXgmwJSnDJJk9p1+0OFz+0rJGPjfJE2Fi6Lxwt3f
3QPg6zlG6FUWuPzsQYcZcblyPpwX2Dq2vnsipYwSM115K2EAJriHS2Y4BoHMBMWrLhjsZr3eVrPP
ql9VVBFnUvG6oLKeN97abJUOFyvy2QhwmZGRIe2143yfQzMXCH7JUzhq/fshL89YoE7GZjDiG4wx
CtNeKAEIPr4fPsVUzXgbYfay/16ybE/l0L7gIlMTDKlgeiUBO4luCbzig+QYKgZ6hDGU+jWF739k
pCSbcjAR67IxlyRbM5LsqvUZbRSehwsQBGPsWAa3yvSRXEuM1LSPvN87Cfhf3kttMdsoMKR1GiaV
7pMrsiQpdhHuLcOv0ifqJO2oqafMg+sKI8cy4KWk7rwYnI2EVXgBjo8ivrSjOxSkb+hw2I53rhXC
x6vRJtDABDYv1SCap74n0g9EYIssoCVh7/zBL7QNf8cXZckDvgbDjbwcrEKZe/RX12J9RJdho0nB
5T5i6pO/DHY3JhEa1uSWMn/fKEzvTIAZW1YFiFOZ3UeG2Bt6OLy7/RuM9wKrzk9rqEjQf6fTnCae
o3F7mRWOGwN7lNXfAHyRxASFQCicFHItOJi5mIaEFqRaWM2nBsxi5d3yMx1iw75ho4VAkjdAJhlj
pItbwweoZ8q+gqBYzObcXc00GehE42leUegXFsQ7rxuLfxlTNiVENSGV3aCl1IudZuPOZba3F5zu
pZ37ylXI9fTDqffz/BK4HzaIQqrM+4jgw3DnxTmUgghk+pFgXBwZe1LmqQAxvDgslBQYwzeNHb0k
eDx2DYDkgUapEQj3V5e6iB/wHsw9g+w8dOO3J5/iMuqiqvzLpn3VS5dUp+BhPWwS3t4PZjc6wblI
BffDyKLQCxeqIPwIrDvAghPTx0uRP0ekWFnXdNvZAYx4cKLTS3/IFmv6EQJiJ/Wy2OJXta/+G7pY
yilV6Hf6L+WDSU+1KrFp06lVttgghA2b/TCQKhLAGWRO22TzakOexP7vIhCHs3S1v7LETDrMIcot
g7B/g7xLSn1EIB7YwibWN0dvVfqHBzg9n/AxVa+QgN29eBpmNbKsn9lIJ6rzPts4Nyp7km9mkeq9
/vqJOZqstE2TYqfi5LQHAA3QEnycjWQzuRNpZgj+cFsZqg4/VH195htdWM2a12EU7PDa4mtt0AuQ
fJhyoQVAbNOXysovNWbe8y7aRSGihlAAUSa3LW4tS26VAVX64tNyZUH8MvNEY49W95jp752KiuD7
GIt+wNS8NKHYJDmQDbqF/2Sd81IZAS7DecntvcR7mQjazw7ji0uMXD6iASccO1kQf2sWkvz7Iv3H
2Qx3HPGO3jcu+p6kStdFmd8aFW85jZMyNasr/wvIsxXRkmLMdb5S2nmGTPN4Y+OunazbfOrXRSce
Cx+OfXdVbOeXqY4HECLgySTSIp3/SxSryEXHae8xYKxYpgLXvpR1OBeYYTWbGpTUPZzbCXErKbUa
dfJIN3l1XfM0qjL+QzX+DQcZAUBwhq7T7wX61TdiAsh/ub/zWyr0/3MzhztTaiPvMIO+s8V3n58t
9ZTsXolBxUs2UDE1vFbmj4Z5CB6302blYi6E6gOz4HQDGdAVt8RN3HWRX9yOsqp/8JoDTcvH0q1l
I+W9i7LN1P75yDCLmP87o5wNoVn/wUXk/2sYKzPgZCaWm3pZPCyjS7bakDS48UWNlzKGCLZdF63l
Wg+zl0Sx9krBeyiBm+PNXoMSoAfWjN2w/WI1rBmgvAX4dBGt8c4iIxWCNOuB8pNn0kXKWRO1peTK
lJ4N11rOyyhYZA7AuaR9mca7mRofQ2tvozkmjcj3jucPY5JZdL4UtNkSoU2ttsoa1Ceo1AcBb+1I
aMHyyHh/eberOyBvyPxk/nL6NZeFvZ3KzHwJr8lfDsPLXombs8SG+rzniMAy9Uy63OCe9pbzrMad
0a9//gjQUIXoIy6GiX5xtgV4IUlduGYzmuQZjuykZdGzyj6JE8BOkQUgS8vBctYH7s0vJHE2bQn9
3GcNsqE+2UILy4drVlRX3ru7qeKtXVJIPcfppzimSpKxW5KZkjBopVjm7rle0i0Pxz/02/eYuPnQ
NuH/LCedyFmXekUzGPpmexzmqABPxMbW0zH0n/c2FRYjDHf16coHVPORtMo0WO8xAypzgBAllDXA
rvV65stZiivRBew7/uCt6DjxJsx56VXihqAJ/ffhMEy/79/QLmlxQ3WG1MSJvKxhaELnJGNwQRmY
USn2OGCnAuv447bpToon37j8akGjBYgWcvoWON7LeKW0VyqJM4gdRTQ2uaLCBX7WuU97xHrujvHc
1aqwglPzDqTB9tBYSBaa1cBd+asX7GORl4OgcJ/X5yTlPTalRwn1kBwhoL6ailpc+7xi6XZLQb2j
Ujw3TlILatIkSpiS8yPtjnmUwWeJ6hDxqtUwsGdHOyvHO50zwP8/Kc7wftSYB24GQvj9bu2qdbPP
M6VXPBs9Engv12ylopiY/nuLgCQYMd4SQ1/HQhiQVDytRp0h3OEyaeCpHNHYQ1sPLP5yd6vn4d41
KdgJByMVkKPaNfZuIX+xAWmJmxwsLaOBddIZxgwck0nMIVDRaEzu36psEVN7CPKPplwO7eBj8DrM
I8CBBFGTQ+kn/ciKXLV1N0hK7RjmMXpndwsskIxPWE7Wm6oYNzfXvApdEMQjnExfdPhg0T6LuaYP
Flm+9pdZye4UDauCjIFUkuV7z44AmJFAztc/Was5CZKqRpEKC+G28s0RsPUefzCas/Q/PCvCtYMB
NC50n+L5N5kut2i/5IOYdw0Bhrsb5YpNe7+JwJQfExV3Vuwrvi2Mvu1Vt7IJ9QLdMj74QxfaNJQo
Gkn0m5YV53qp25G650kKjyfXr1D3lN5DFiDt2lTSdFhvTTn8H1alM0C9uVe6iS4Ho6GfyONMQ7F6
NnRDvKaGXg0kuOkJooQJHSwXbOFW5s7vlwq3LU8Bjq8HJHWMA8qTO5yomUw7Exkr5oGg62WjmpOS
p7f3YAiBzdwBnnQhm04aDieFXM1oD8ZCDHLE2iM2UuOIanrHyu/9PCBTq7W1XjIClxe2QAXJJ1nH
U1AB/WOxhLGXQGoSPJiA/bLPuekQO38g0w72WKsowUZ90mBl1ImIjci584GArGS0NzcCfjkgLFXq
OPLqzN9MN24/RHMQMwsjoPVWADBUHaRh8b6ryRb/qgkf1qyUpit45CwvXmLgPGQLoNUKS7Uq4CxJ
jJ3cPRwrve0MHkLEy02JkqKMWAElYUjF/mUfWvxNUXma6hdYRE30dsdG+UZ/BhsLeCaLgyjI5N8B
oZVF7q1ux5QabRkSjotmXrUNr7uwoVx4UtgdlCjiKBvuKFf+a6W7P4GnPJADR4B5GN3bT+wLgKwL
sUrtBd1+RtnFPqmAtaiog/1aifM3+hiMY/9FzUQSPOPeT9WkpC7FFvB0cUppbXS+1KoxfuWRXwN7
AYMCkLfy0eIkWtBOHriUWW8sEvLJFlwvrsBNr0oTZdxUDaYajPa+USVqOpX4cc855rATUWnw1YCc
COi+uVN2drOlfN5gNlxh82TnRNKCikyMGrWS8uDxvbt8P8SV5QBlEdysdGqvdR4qIhHN5EB+R/a5
j7YxugbCLOf55T5wIoGpv5jbb3gmVfDAWwj5V/OhgjczL0isorkSRY9x/WxHeFhXT3spdfbts7Co
NPQjaw5Vn1kN8cM0Yf4ByagRYd3y/gLodnxewpZVS8xZ88kRYxCF2+wen62pO6aexFlmRoKw12GY
jTmlRKWYhlDqKfUCFtI4XYGGIuFRKXlEBqpRkOcGa2r9wddB2wbgAog2KY50VDL3Yotej+nEdC2+
Zjqr1yiXTTd+OL26LOZqQ/52ze3s7L5mMwm1ZgpypC/7wP+mQX8gNKiIbJEv1jGdr+lZaueTbTU+
UQAfbJnxgL/v9ZW16EcZLRKq2/hnjKno9Xu2p0xKkjEaDm9QVYk8JpSJv9JcrogEiy4iRBvVpgRK
o1k5DfjeDZDC0qdr0oXzVrXOw62SCHQIrGMe+2wXbud9yzkNY8DSSLVazNdxH/s7R/0b6749cADq
QXIis+Lf3vyTkxhPWOvdNYmOk+9xD/fOAvQg4JHaVy1gNUWqHm/nUnE74Wj8cV+s9dsId/8d0h4E
l/JShBzU6AatWLzQpEVOehm2tOHFv6w1gjJLQyx+BfU6t2BFjBfqnMv3BJvdIUErc80erwLSkHTt
aC10FCm5OuzDfUazA3M0QpNQUmC85sMe5Hw5NxwsmURZQwLuikko+xbiNJO/HZTBEIpWGo5ySnfI
ewKzAzAh9Rw9i6ENaeenR1daYpH2i0jk4R5+iLkQ8/U0/2wZMJs4kDBnZccxOaEs++rhBBO8OKo9
qCUiJNYdVOuqs4UeGVK1C8wFhMxzXVii41rEg+ThL75tXDlp+OyP423dcIqWBM+VOig7eDhl8yAw
v+TVssWbJwlP8n8FFuO+gY38EqQy31fPML4X+VnvwG/tfEv4IJ73CfIiRcgaDrNDOhznPDCAeLZ4
tJiKa6AwvShDgThlFXzvmz2/ineWNwWtRoe7FQhS/Pkn20TQYU/Q2s9XbXqe5GgE9DPSpJCfOis7
TXoyk/2kPSMHSq2OkyXDq/zaSJFH30Ut200t/zQVUZRc7nrcUo5xu+9s/Z6FJl89GXgTpc00e48P
ydnSbDH5XUIFCdCP1Q9YLnPwPpskEayIUtXeNPOTy2UqgTIF9dJMnQy6dcswJRHBR5mTHNVOmg7p
B4gem1ZdSgQVbBW0HIqXtUolWjtVJOoJKXYsR8O52dKMCOWYnhCG6ANu8KDqGcEP2to/QMKSAOGM
bH52I8eKJUDKAtw91jtDuLkNAnw/Qedo/JuWYlgPk0zp96Ijzj1sSYZxZUitY7dKhs3jNyYzKSUU
J+PLDgIyXsTEPlZevJsqK0butuiXFGmS8qP87+mKJJfLJ1zywVBjgDmO/nWWrGsR+dDtyX8p/po4
SCPr7wT5ouS/KK5QLF747/FG7iUlWhS5ERMU8eSHpudfoI6Wk28npXbILhIb6qjluDfkkwUTQqGK
N/pZmfPLsqx1qly1oNqxAZGjUBMv+Ts2tfWDVWWweYPcIIzIrTy3Gnfy3lBJ3tcfsmmvc3b1z51S
6il5kbxvRrhV3YCxoJBOpX2QrExGiLFiGibHKW5hVSr6L3aHHvr/ev66y5ONXYbP2zPU7TmGoMhB
TdYDXDHSbF5/xr6grO1E/oal+92EAtYILgJESwMZ/8j11xG7ePNK8iQTbbiR8Gie6jGL7/OuXQHT
skvulkg4xSyCQmZ6OIilN7qKa/fIev0CH4XBrJe9aaTYZVntEeGSEPGZDMzaqvGdbQXpg/e4FVth
ZsCqjC+3P4G7Vt+45hkG1UDNmg/+85X5p/YcvT1QZryV01rLL/eH1Dl7cj9iPz7jnZdnLTRh9u3P
VtfQ4GZHqKBJPm03rBDHQNfLOWfmwEKpOcE0MvcH6IsQGIN7XOBCE1o5gZ5jF7bBTR5p4SNcZQtC
TYSltqHWy+LrTMEgPG7eAlK3sS6M2rHOn7IKNMnS869PG3KWeY0H2pabNbMObNYxnUm3jvIHeOrx
HdmYvxLVfzBle0C8bPQzvkhsHmPJpjJA1CCUQWK6UICEuDi9DjuNQnVGcnU6AIV3iduqm3/dVvuD
hCMETeXoln1js5AbHeyTDFf84xDNKGeAHCfYLCvs86p3vA12Usk+rb+ZdXlYNRis9Eowhyj6cmAm
NUPiQJ6PwveV2E96y0zg5z1YIZG/PuH2rJjm6PPCg1oyogiaUJpPhetBdCBVGwbvOLAagBTqtBdJ
idTRLHOMQLd2njAxDKHRzdwQG1KUr+Rj0X+j55WZKa6bpQM5v5GFlJnNXAzPEmoDoZsI3VhMqKXv
UIPhbCIgBFKEhPg5cke8mwhsuVpYn6rC9BocIjVeekJSA39JpQ3rFZfvOkLgohQBgik+KOYogjHB
lrfIT6YzWOLRtLplKJhXaZvV/Zx2EagF2WecZwnnrePCeVYD8+u413FN3w5wMaIALvtmoobpj2rW
yoWkuMbIH+0E/V4rRYQy7V9ZguTEQ19RGuKvHsX0COaDmxwoviKsaFA8oqyTlOmLoeBwPvo4BAaP
/CLtFe+30aSCFbxvuPMva9yverGrI1I4aCMmGiws48Q9g3bOsUZd4y/t7OOx7g9YVM3d2THFGH4s
KR/Zzgh8Q2swbOzvBcV5mB5aZf8ehZUbY7DULq1Vilh3ltHi/Ijre/Alzn/FSScIdD9kNnu7e2Yp
Z25A+DcQvdkZnRwVqAWlXlptQQcu0JOy9C6mpHvrwzA+4wg4HJ5GcbdwlmJ+D3IhgBUrjKvuX+s2
lOrCvmo2M9APvgjizAQakws0Mdf3njZ319mytrTMQQx8MpbaS8Aw4jemnkiKyj2YPdGHzzLx9sn3
5A9hb4dJbJISYdZt6L7301rkrcDaIE63u0/J5sxnlGqR8HHtqgn6mLy+HOE2LyswlDQJ+CyN5x6+
G4KRAF85/DjPr6Y1rwp63HY70JntSK0rdYeN5s7iW3+MsIKF2Is00oBtVtokMMoKNBaqJdh3Kaiq
BvxxyPHMElsYgPyXJgQp+V967NoofeHs6EEZWDVsl9kc7+FpteDFFuLs6dUKC6hb79ZDVp0ZqzD6
gns2tqbAczP/w7HBANswVCLRGdngzRBeZRXmuOE9edz5XR0Fg4deTCO+gtxmOmNYbtAuRiCjPdZu
XgQuMsJ+FAMBCbkoTzDhnFDAxHLjyZ5KNyLdMbADi0bh9HFwPHzQhLU3NKI0GLazv75quTtkSBD0
DyLvoFBeDTkZeCKKtabNC+EPlqnzzXajt6XQSpmHRxL7PEHUpUQo5t/0i26W0oed8BB0uQ3eOQRR
yVWK8zhuXfIxrMbeZryPEROzVu/2T9y8xTOAHcdst+WBLUDmNJrsQA1XF8iB2QKM3iDTHNvAJ1+j
fAiltPAmNOdLnOZ8fYtQq0n7hXn7YABYZ2uL07sd5cawMDAbMVOURoXbQ8p7D2YaGBTOu+3ADXzz
S8j8bqZJpIGiizRWl0NxmIwhKO/K2qTBvb5btGytNVyP/ZgHQ1KnsutVIgoAomWSkuLyJyUz4PcN
R66tJXVtPlWvXzXSUjLGtjtxiFvpHh0HBNoqiFEWFIM+RmuPoqwNWMiktyZCyVX9XxKHthV6aEEQ
HpG7VvDwDquoud5KqWBlBheZHcLcogtcVXGBfxNYeU15DFV2DbNFFjNQnayRoPqKnaJjaB+hYUjj
r0JMTMpyjOHnmiqBytHVbPnLKgMi8DQ+kUtjQd4warAuFDQpmfIqzWb7YftAhEWobS0q6JiSTnRC
tzHl4H1lcMLN+h/Vnb+QlZ/zvvoTukCAw6LonqHcZukY/lApDJwSYJSl9qU19jPZFH63e03me2zj
wGAnoynnOejOur+REycEYbPOdCVbQT5oPjUoc7etv1hE3cJ9vxDBs9PpkTWLtUlQb48/EmcUlOn7
GvDuoSKlUHe54plVDzqcA8kvM197Jl/3mUKDQACPgfvcvXEuq9k/LrSYKyqiBD8KrO6D04xZTzQg
ECHAUm29Ta2hDoQUmS9+zuO7v0azBTwP391ON7J42AD5VRmT39gyWRgNvgI2uYT1+Sdcw+6Mx6U4
0yGxH3j3x3yM7uD/XgFzkq5rilEPDMMH2Cu/wlmWgTlFjROXwZWaxCSN2r71VI7ujp8ZshBPuflu
1j6x0dfUFCYOE/D2vvtOFhQb3hwtsy9Y/A+9ZW7QmdAyABvHml/HFfEdj4gmcQRjyrHimx13sH8t
o2ikoiJPiR47zne6n4rXlQH0ljVoVacgo1acOqvclP17hNVzkDnJ+trzFPxNFTzGiuMUSceIWIdf
P88odL3IQ7kcgzPvguSw9ROCOVuJt0qyiHyfQSfu5PxjNU+yjB11kj1R81cB1hB/y65sXYf4ersk
Zwm06lzBX5FzVsjOH2AbYTEAowpXCFVCuWJPV8ypVdJwxMGeR1zQHABOp5Htv35l8LuwcIceHI0q
CxMh3RfSiReiQBWSVATQMKwvk7RCEUkxrAfSZOShNC6MFGIbrUMiM3H0KWk3oqS5DLKjW+5zUf6B
Ji5F24vk5pg4LxOvsIxTH96gUhroTJxcRQxAjyuofLyHmt8LRT+gtdM7Rwx/khoFerf6jVXGpS7+
njvYNcQLFwnkm96qtpxc5briWI9PYjPYP9CnutbmyQ7svR7E6Z5F9BWv4RYRcru7CIgZ0+L0UpKD
K16MapyUTyUZQiSTaPRUOkFr5+bJXi0/OKf/83jEI+kRRBB/F0hJVNDQLdq7V/uWu6cbD1yJBVq4
GRD3dspCUCMVR5UsLz2v9ULnWFlgO9eu/Z5AZ+DJF+1sLuJW4K9JDMYtX9ocJpQeFEpwHmTTEibI
XBQOqm1ygRUP9pU0RrM/4WoWg3f4tGAAfs3WT0iOARD9rshMaRDDjdeYlRMcXBC40LoEFIg2EV5p
C0J6ZH1BM4Og3Vd53xMe3wC0eURFvyCcodOdX7TVfDgdC6wT1fMRLoz29UA7nikoRBJFyBcKDWr9
g08ksZdNGClEhuBynqZ9LoZS4OrVO6cnA8iRbJCehDGv9S3jAsVuJnvoRNbW3mP54hkB6LJghavY
4BND5/2072MusN48MNfH8YycCCClaEuCr1uIKCZQ2w5eUdwvagn5CvE7YR70dzf8418dAGqqfVa/
IG9lcvneQH6lprxBC1AkvpaciAQfs4+7WMFdBEmQBv9NRUCUHb9+jD+Xcwh8uLGqFmepWRF7fMvN
AjtF/IT67flk9CgLgFoKPNg7LtTxhD309qqnacr4GazKI8eAS+vVHrY8EEeo6SShq6x4CgUieoSq
tT76CtMG4XJqkfbF8FKYajMqsPzVBOrfwquvsqtt3fQL2N6Dzb2+RUKlDDPxwaEHFWjMrxdUF/u2
/bBAim+eY2J1rB3meZElrh7z+UkPmEyC0qzUKAKIPe2Vr6+2RlYwqiJJtYbFJAc7mVsr6ZAFvIoG
pvxvAw2azbZGc/2Y1ELLx2eFhtG6EA57IRpFQ8CtXKfHwcSNYXVt9gkHyT0RtwQPGfWR9QsToDf2
EpBXh4YhgWEND/ZgWGxg5RpnPCpJ69v0yrLVS3GlT0A4MqXG3Jp7KjN2Xknza5YYUEBk/eekJWy6
zO9xhsp/4t3M7kSKzllFeB4Oab3iaSRyarcdlPiCIfeLOXImxzRHlmEwpnzxNmbRgwLB7HfxuBLA
EdJZyEQE6fLDSfhlxl2vQk8gLj8cOHL0q1bYaBmpbZUBp+PKX1hqFaWcuW0OUHs6UbjMIVGKFWho
iLKlCca5KopkAke/Gx39tcfDvrls8MQlEgijGmwk4fuYCJ2D3ssh6+DwFfZEw/PaYGbJwUoYMugE
nRHDS2Gy64WbqoGAJ7ykdpALcywWVWkaR3YxfnJog5WewNeIRxE/rUkhpNor/xlEze9XaVYGzonb
f6k4we7D6XA5bkyuD393MO+QV80FhaQqd+ij5V+nRJOtPqqzhEMmOzKfWa9ClTGbxKwkdS/4+Zer
y7TCQXDpL1k7ogq5P1IjjzCgHJFCY5PMyE9b7D1IMhELQv9OQXjESOypriEkAa5mOsqrPQg5PQqk
RWyUmgSS7/8aqDV2X04m6SFBfRDw4GiYspOCMC/pWQMGN+ZwamGe3XdYbHY0wgJ5oT32cJI8OSWQ
wGxv0HNGR7REgONml2XW5CTffJLWLO9Si87TwkQSFMXBcGcZNTmKELLJr2K9kbUatFeX5bY2nzQI
AFVR8krNkGGaCdMnZO3wGa6+3msz9QYYCwRdJBlXwqXMIcSScp8yA+EAv1EIrPTJvde/Do+ox9gw
Xd/QB+i9S89r4TKv5Gsp6KiAN3av6HGzuHzSPUn66yo3qbU1NneBXHQ7b60Xics8EnT00MeSdowC
7LMpjyQ3OPr+IKleWfnLzdVQc2quV4cT10y/NwUinJwKZVX2j01XISCWu1Kz/mgSVJExdf/yZj2s
jSD1FpIdrJbzBEOpNdzEymIIAIA2yixZRcMdDaHlJfx/kIbjJ0fii/xmOjnmbySNXAyMfLiLudog
QMg9gTkNqhKVnoZD10J93kFvIKUDEnkUURpRgsTuwIlmG4VUH2C1YpdH/DzWm5D27QjugCg7A0+j
CL4Zy9/uon8ICNL8/83/9yA+MZdlKKK5Lzd6trGJVg+17ElYSDbY+wUzdS46WEsXdeUmD6fubPco
Ap+1NT5pW8cX5PIytAbrM8OxN56HsK0N22VegRWbCusLd5KXrFcmSi/9KA2xWaXoiiHgbqBN3gtF
Bo9Y9T6CvV9UCms1378NFOeKi6HEgNj9DiVvT3+kA7b6i5mpm8GP6QCAzyWp2Vj6aBqPYV1HBVQT
FDvGPDkL8HcTK68nAipEcbTmRoQh88jpGDHdqTyLOsMvBrF/5Paa1pYhPt5RlV9ec6ejAsxufkQK
uNNiekpzLBqwNEvakAvEdNyoYLv2Y0xX39wjyKn7D2NK43+yy8vkPyMlJIePswhdtiELNdHOuJ4s
8PJgUtvCmrX595mXYwDC1D0gPnvWlbg0ttJqEZhe96VOV4r6HH3FEGEBPOeu+EoZVyxHT06IkKnN
qcjy9zVUNjGii5d/xIQn0RT3xpZmooJXsTQvUvbu3viwx+HNDWkNPzRXfLMZ/yWaN7XI+Gslruyz
anKYp3EXi3wn/9bO/nFYbheornZ5ulLQsUFe7uMqORNjdKzmTaqv64jbZwaBLc37i/H8NQpc3rqo
WwVlsgLcbuDw6YsZqX11IiP741/GqAG9ri7PxQN+waDhzSF7/prEfq2kXolpOEjbleS0TwAHWMFq
x2QE7/pwz2WTeh3vXOar41jm8l92DHFw4FRr4tov5IjmEDLqZ85sTwNeYAUXy6Mgr7KoiGbnF3kx
khYQSKuCwIrvspmwR2l5mGxHJdOZkUbpwfkoei+UnurONR7M8NOVKywsyS+uHAJRBsThgyAd/FEK
J4upmomU2uRSCKVKHRvTCEYSoQwr56kRiMPMtL189n4HjfcOUoOUSpqwBvKWBG9JkN0+FlU3lA45
UuQZtvA22ztC1mQ/Km7Ia3P8ht8nyB/bjgH3yK3YqcyG4GlQFxIsskaJOee1jm2gULpH0vBCGe6z
hswUFHojgknmrBKnbLQKQ1DVjOn7BH1Bma/nrwCGyFctaDL6yP09CZQzKxRvb5pcV0dLVYs40qRf
lMDrRMu4jhX9b2ZIb4mPW+nEbUrwtqErNKqZm5oss8+0PxGfKF3k09rFESVOlwm3jekkWZ839agA
Bvm8CHlw4fGQYeBhtrp80xWLPxuE39Y9DnRZTltYu41d/VNmsliWQ8nVbc2B7cxQ5nhpx1AD1fKG
VEkgScpySiZMBBBVNejlzhIwF7Zculz6Bkb/FOHu8v2YK3J1YqwOO/uSp+69zTFkaFWCI6xsaYGd
+HWq9ZARx0anwni4/72KeOw0ZXxoI5J30qGzGpUVKZrXj1fY1Uippl9I/7DEiulOtQWnAkfPO5jA
jzvSPRxzMabQUR7RbClaKHuMdYAgcTgMiwhYaAtdYKT5Cuf+olm4CQBbXF8w3HoikadEbVMR54f5
OMlFD07FOmbn30xAKdybOKDxEuodn4+SRMRoSRnBPtB5XE//gXi9GlbxL+biPd3hJ1hIgKB/QJcL
qEDk2hlBTpdS/U8WOn4+s1rV5Rz1mO/5mVkgVTQhHNDbes8AYAXhWo106I+5VqkhH0WS2ip4e+dd
pCutPd8EukEozVKXSWLGf0pWtkgH/pfLNmywLW6a+VYd7PHPQbG4y6mAjUrJ+fOjmXmXZGHk/9LW
ReX84oGqKP2gDaUY3evb7grOKJTp5zwXi0+Y76ElcjIz13Z/LSxCZtsVy8X9B6wK5VwXwdvSEKlN
ipdaZIg8pzfp85RQf/m3marny7r18RCphI9cCuTo7DrnKwjv5ZkSF3I1dHTQqsN/26AjRcSKKLKF
04z0f+71VME0KZMeyWCAOqA5idycuzM+Ril068bt4ths/H9YxI4ZDbh8Fp6oEHBbHVIuTDHGz0AG
LS4Ws6lu31fHmks9LCHDLdSgTjNxH66HAyGweLznTZV7Rjdh32mWqQLiganm9dUPS6+vUji4Tfld
MXMecUJhAK+D9KaJpNyshMkqa1DnV64LfH0zogPF/4GgjuC7oiQ9pl/9/yerHfC0oqcoajC57zMS
1UXb1GME0lXQ4lKra9feYiWcqrEMTxhkEBOKk2edYVKwJpZQ/AGRIlvtxxQXG21v8vj7fuJExSWt
5vMtzLS0Pl5tIw69O6Dp/1wtH7k8l7QDNUAuI+X44hROmfJNdTmYAvAROwgjgyD8Iy1shSUfsXgi
5pBSBLyZ6WskJFXaKHgDN+CmWnv9tfXTF56flGSGJTy6oNW9kftb2OfAMVTgFHZPGUQizv3aA2Ug
zSf7FPpvMoenYbF8X+Ql9HdF1AmCDu694+j0m2VdZZby6uVsNkVecPy36NSNOt0H/96djCSr4e58
a2dAPSb/jjXDNqwLcu8FHQcWenX2k8Lp4ZmNMGNlVPqlYqV/hdJ1Q3cgzhnYDG3S364XajS+/MlH
QYpBuBAP2Zq4cudtS9hBlkLAknU0aVZuJuuCaoq5VXufrCdN70+v9sS+AZWgZayz/LTMVKOqYaJs
aajZfyfK3SmVvpuwuFDN0AC9wW2Ydu2Zr8DWWXKqub0dXEQBTLwPF0wY6n8tiAS7gDwEmwlqyBf0
dTPDYsDVz0bZgBmfmrHCMKxiGHwo1OzUGtNqla65TkJPc3+sw54QahmZ/GZFeBBQgoUu5/5867qd
ovNbS29agnFCSW3dhbt70wnctDZSyqTVhOmgEqinop3NjV0Lq3a8RMV+MFEd1E6/sGaoQO4rwmDO
ZtajvwhNIx9GyKpQILug9eePB6cWkq297hPPbiCn4SYXwSgL43/4r6U6/61ZUmlPTz8LXFE2/aky
jO1txoYJT3AIOuFtLCfIAHFB8jF/tkjGy0mfdb5kD6Gf+K+Qifz+Xrl7QNuKIz04cnU5VIs+8vCj
uQdapUnz6yTMU3nrNlpXdHR903rrAnbO/bgCtwbuLHEWHdcvmsu3b2rk99q6oUx7SOtuyHCH6HZZ
MggXGvXhWZFtQbRtI/8QZ989u8YQyMpsJXz6v7wfLMP+3gpcdTNe9BBOetGNwHFnZaeFsAX7rMJ/
d2fYP6MizHNgpZ0voxzilcsUoVmfA8ad5k9BmpaKCCnFOiSsO6LU+A+pGqt0K9AXwJVd700AoQ9Z
G2NVZwcQA1UydPC9c/Y/HZKRziA8sMGgN0rjEMgchIqlzK4kZUjvk+ZYhB5NV2cIHhb/mILI4gNm
ClWRWJpWtcD+STQC7lDtP70Y+AiEOm2KRTqZa5Oc/AE53s2oQHHhsH0+N9wMhYP9EsM5v4PEdMCM
pdlHrH6nipA9WOeQ3LO2DCopn2Ict6bAqRPBwUfQuiPqjls4OlJ/+/BNZQc8FdbAAp57ydTn3FJk
ZQfO2eyWf/4J0D0GESy5Nw217dZz2Sav9sJIjJexBOzvIm4zdRHcDS2H1alFmU/Z9m8lbtHvLPpa
RU/rHEui5F5cZHiDVUGrK8A9leXZiNHNqA/iymniX/6AiKM1FnrsqTxTdYp+HKMx4U48JHerBP+R
hdeaNVvhW3yPehDHjdwRqH1bXOBAlskTz290mBRQ03tjesZCiXoh3fnAIfrRoYTKx2sntcIPcqVu
HpuPcGqT6sBRm4v3RfnL+E7V02mDdu2NdF0YtGDqYJrcLoYUKFEVfTzImhKjeHI+b8r3RyYZUaiO
FKaC3O+0EGvdwHdiss7qDUkFLSeQZsatMiiBDoKg5+AcWY/RcsTYxUG1hKSRMTXspP+1BhmEhbEA
ntn7/McqEmzvTfY3CCQcMVs1rjjXQeUuyayDEasfsZouxO5M5e092W99y9VuSK+swL0Puu6mqMh5
6ANn/Z5ybzm1txyAV5M6/Ai/BAkAVS2HKidUQ+GMz6unAUStCA69U7d7sg60Wpq0IUIJZyP090ow
PIQtASf4Vt8k9TG5rvQ7YzHF9El4yZRZXAnThyUxLlehT+RASFa/KiAPyNy5W8mN2ZL2RxuEIXcp
iGF0ucvqbwD0yaxTgXjTA/SsN8ThYTcgGhzirYQjJxZxgVTumfrrHgj7GN9mpP0hbsI7+LZFtLoK
Ypej/gn6t147jDrSadqTfkFhv2JxaVoPXTKfGrcexzDQp7vha8b4jggYyM+N7bZJnhybqwqRFEON
aPI21Su8nPZHKSlNuXBG+0p7vRb2u0Ry2PpVKjop1kywwHQ1L+kjU/8O0PVsewGxnQTUdZy+Jl7Y
vD72FfZu6rB/UVSIHeqrAWbAAGIIp0xo4BqMqnR1YswhPDrEWlbB4mK83X3cNcL8e5zDNkeNnjIH
SV8mAB89j4XnzcwkrUFk52Wx32J9chSgSX8ev+NwTAUjDGdQkWhbNofZ8c+FzNHqS5D4DcPRPkDv
PTZKRlj6Q5O9IOO/Iu61qy3YwjNez9tuJcqGFdCBGt73z4wdlnwHjrFzjm2lCHPQIid6tYDcNwUl
PrE8IMVhYiDVoOwjf9Y4c3hkHUP0xR+0ipNmPeRN2ifI8wldxc/JNpCSEYdmy4l3vF2C47IcWT3o
WyhuuF3Vxe3ECu793rKs7e2IwMZ9/aGcom2dxH5cOPg3wE1ZXWifo05IizCJloamPJpKFEn7M48g
P7ofb5jsrvtjCxZrUbT4X2j3h3pFInhUL2Oo49E9mvNdDgM/qZRspEr/+w+kXxKjOICoc5NvQbh5
HLwktwBToa0GJUGF0xWuIs/upC1OJyU6geU4SqJCTt0kMBn0vn8Rhj7dm6n2gR8PYvMb4cXDOyL8
wuxM1j0yKDJQjdNpeuxBHMKu5jTYEJ0eCno3O30Y5vbwEBFQACTrbzMOd0LTophk1YV8KwhfVTk7
fHcVosvRJSaiOhw1hVhetOO1RD5lPMnG2X4KiS/JPVMnPVwnNMOgypUTM/3vg4z1LD+1qgnk3W0O
YlE2MZDKBZvh/QzW3571vMjKDS046zWaMjufCjyfCASNwqRtOgdwfXIXQSxbzaVGgO9sDjtPfO+Z
slY2dVkv5L8JGKdtLl5RUorzs6xvgxMTMf+FZmGtNn+9DVJI55r6p4RBaYxN8wRa68J3c+wDu1TC
JQEh/ORgfoMl3yOTn5UsgPR65GAzLaMN57icENk5AbsNr5lvaXd1w/QOwiYpa5Kp76hXgwwOuY83
kup4rGiVrTnDZWcqJh0GhDTF4xMNHTkDayT4ZUelno6e4ryINvRmEy3pKmBAGZmmEezyDO1GKgmH
BWMY4bGfhmcM4HC5lD0YF9TWpOHqLV3UbtoUJclX/Xm2wpua4ziemYP0TFHYR2WDR4ZfvUBwqPWw
GMUVgdCz9XElw2CEqmgVSNAZOuwyL/g4eBAILY9TUOf8W1NqsYff6JTAzvQy1Y6H4FGo5ARPKSaK
F0VkgaAiBobANyxFsVKxMOrHGXgF5ZYL7a5Jj9nNLlAvGX8iSLAFLf2eh/wnBXXE9Q3Z2ph0l7W1
k7eJ0ws1iYfssEdCFthoZ2QrBwPzrkg8SIr8tL3/Vj4Vff10+m+jzvnMQq4k6caTYAcdhUiQjxC7
Zxn7z3tsZOFRbWcxt+ydmvvQui/6RvQpFVhHCz/GnjYwZCesz/xf0X9SLOp8iL0N1x6Tiyz5m67g
uL4rjNkp8RUYAF41S2MjDNMUWn6f2VhEka8z4qr6yf0Rb9xekU5ezL3kULblluNuCsb2bx6dQXhE
4GAv5RFyhv+/8UaLsj8Ht5idZrHYWTlf+9956KNdjASa3K4ne+q9u/7wINN2bFT5Hi39N5TOOwdH
cPQCknIM62hyQWwgC8ovZ2kFMCcl1S+AfFtgalDx15Xu/FLU+jMRLqk7JES2Y/+D2J/B9pcwNTMk
gHqfG2Ecwi/m73M53QMYDcnSOqbscLV/mScWYFAHRdlGCGxRNafiW4YqkFi0EUAfJBLgLj21nI5W
w1GuMiM1Y/xXcobfzOyx2hMyOp2zN4vkEN7pmoNZuT6RNG4v5Diveyz4WLZf+1Q4KvbeB4GETtHW
Zji3vjQajJ/V8sVSaXWcgoPMBlVt/8AKA57MuxiP1rlJbDl2MK3c9wPG8928vfuIxU3WBLGKeTSM
Pn79VJ4WgHDrX0NrPXNQm4qa4E+pDdSlDPDr3dGAV6iazriF9793a4FksTCnwIRN/5M5Ko1fzMxM
e4/xpoJPMDJFDsSmbNuNAjcsHrdoOaoEpS/pcRnIPiibEYd4cseU1oPR0OiH0X5YLKXf04L1CDV2
nm81QdRb6Lri0cWWUAjInZuzVeWj6LsgeK5ALY/dIFJQFsxff61eFtBlLhNt8rbPrsRMlS1yCNNX
AS7Y+3qR4W6dCto2SM/8qNozhedRY42dDr8fkeldXDabrG4VAoCSBvhGApa7iuWYa5AvnL95Eka+
z32wwkQ29Aqd00twl+cYeKfbXAuE09ewGqUbOZoyEXTf2kQgwcg+PalKo5pyDeDS2OXluMM60A9y
RBOdyTAgmPoxlLbWHOrcZsCGhgRW14XJxbfEm6+T0JcXZYU3EFURQb8EnxxcBkVd2taEg2XUIVSt
5vLvoE8H1vWwqJYZbHQ36hxCwYHvRWRiRW24zHXfbNJz6l4urcrjlpOySAHjV5GYd/jPTqAJJwwS
s4ZKE6D4qHQOHAL6UGGG+3P8pZWYcIT2LHaXB24i6WXwBwiw6GvsRHUBMJf9SaKT7gBSd5VrK8m8
/pA6tUayrnDKSzVfhRh9WViqSQ8nmfWgyOptk9oaRWJbarSKxXTC6xZfykaVqmUbu5+wr1DzDR1Z
V8NhfleXdquDoWwhYU+kb32NAkDcyLvwXs1nY+wTstAxFf7jtlTkKM9CHGaCNQrfOy6QrIUbjuLY
IANMI6qLGtVFZhn4cHAYILGI9X1zeXoWGWJmEOmRqJakj4ri87OGW5l59c0eAr7ajoiR89WPKb1G
DOqOEu8nbKCzXjlmP0ZV6l5yGYjDffczU6HP6yjAAh3JA0RQ1V4IFz7KmgmlVfno8T/HUdi9/7he
SCR1x4fxFmUOZGoDM4PlxBcuAPNPO0IqsDOj0A8aEyLIQbO38hZe7aRZkJ5GO2XQLdLO0o2OyXXm
ie2srnBJqLm6k3WY+GQrfdbAfC14CXaAYtAk3pI/grZkQDckMY28WTvCCF5MhI3fDvJDXD/xUCgU
ePclkC/IWSGjJi9CaTA79HxSWhNCFKU5xcB6EL2IHDecFJgzNslLKZl2oWp4/SUfg0Q4hY5rUNbO
0/hZzhnlMtluYUdG8etyhzCS/d0c2WhnmHNbAv7Y2G+5odEJUBziRX1lQ0F7hWOa4tMKDJgQ/Rwm
FRAh/dJ9mjzU48S6mlct8MqCEu/Qyu9o7cKUd6dL0PzAvqHClKjDyeyszIhyxRi71OfThCo+0VdB
+qrRzYDSK29zZau5/Ev8e+sN+Vy01CmEbPnV8heWYrCPG5SP/3z8VKAc8510cR98b7hw2buxPrS1
nkcz2YeXdBLGQ0/o23J9oH3jNMiA6RhoKEHy6wqq3Rr/5+f+6VE9L8brkowzyhl6pMXmme7yhsye
IROujhanrjcF0P0hL6Jv9y2k7TvDu99iPKh8e7ylZdrOsM6dABwTRtIGwrMpQd7omX3HbzZCsbrd
k/yYmpk3kYjO38XaKYjVlj0uQOFN+/pRq7Gy75MTkK3wv8MphbFnb+imx8Ykic8qcWaFET8HqSz7
CTRYpGqMD3VeIggIhERQkmIkjBemOyouCwOofAJpLpj5VxfCUtGVX1n8Q+xqbS2xZJwHZSXcKI6v
S9ObGAxtfLvKqzBcb4gupctS8Bhj2oPaDKGSMPZ+X6IAwcKfWBbC+7LgK3qYMLa9gUigeN5mTM+6
xEuTbHreXVLgwnzlKy+fRajWQAd8FXJ+8BmL58m8by1Ixvd7lyA7HO5PaJ4+AABsd5UCI9ZqcFb1
wLPkukWI5sopWXxJGrZv79VMssPONaokEXTfxeCjokY12RbVdXBmO0x2hF/ZwdwaKwRMf2q+W6LB
cCk2/IWBfbSfq0XUzyrFexS2pl+Ar7wb1mQb3tz+GjxTkwquVRPfrNbSzqTpM9WANreV67yP46sJ
UiWO7hkJ6hI/OUIsv5IwMcC58zzto+oJJ7Gm5lJemwyXy2z7/kqh/JYI14O0jvQjDsIS+jmUh3nk
phrf+2zW92ciwqYr1vxiANKTkdTc87Igo4lJtsKXAg5sqwz4IH2BGdKPuoeDzT8hn9enQtC52CrN
BfCuj9SvOK72AeRW/Y379SbvKftfidOZ+xcBdz5tLk/ela0OvQt/0AmRzI0f/iUGDxG1PugYX421
dA6R8+tI8nWyhQ/uo3ig4/5nd8AD8d9/NLOIiDixpcBJvmt0jA9R/IqrHAcN5QnFhn5i8xCAnv3k
t14jIOLificTugLDc90WnBb8gja3JHO/lXQviHAXDU26f+e5FlbY1KbTtV4YALYuDSBcmUstUX2n
i6haI+uQlFVudwtbIreS0dPSbiEiWf/LWdveHfEdJ8FBHw2mpAuHh51c6BJO2YKeFkXkAlGAqPcd
ccG4JT/sU1M/Ybn9kylyCoKs0oBTL+InN/ji1ts8bHe5+Xwjj0+niJvgPkdCJ5CbmvXjzh2MT1nf
h+tPZx5f0A1k9z5CoD1oelN64bjZ59pHzy7yYom60egD7KgU0e4ClywU9xcKh+APBJ4r2fwTfrMB
TidBYcG1TrxOUykLgCI6fGAtE//Yy9IRBjm0Go7Rmq4+V4ydPikPC0tvEpZ0Fws7iVd25qj8ENQA
U7GHCjLyWv9m8XoTHHAseOdJqkJwbbp7Gcg2Ox7ys6PfIUJKRl5CxSYMPktC30p7PpSFFihN2USo
5EAJHL97Fo6cWwfK+UMNxxg0Iw+BfN8pgX8B1FHQyXAqAi+uVXPZBhWsjj59NEtXjuQesRU8rDCa
RvgUZ1868ugEL/CPhOa6s41lk+vG8T9RLWXbr9KEcrWEdVVg/yY79hWam/jCaXvaNlkkogeI6goV
7+hEbeIJcDvZ8Dgn3X8Ltsum3JE+0juQPOz7pkhnJPoa8aM5rpKAnPEGYc7cF0IH09Pwsk1R3xQY
H7DKU+/QB4ZzgIxCzuJ2vS/egjDx3tMdaaaQnXLPDYz2imtCd/9/Bz7ZB2gIj8OfiA/mZnAFn4yZ
p9dt0YpgMdA4zIZl9BZUbXhsAyuqgR426QepldPPTYaJ6sRsuMznHe0Cspu0khTAhIzgPQ4z58N+
W38oy3f0DppLKO/kufS1Qnzwt5kBkM3IOmOtnTzw1xkBOi+Tlja59VBfSLsFmBBU8XiCIp+O2tYt
zn5sazHBpPxRoxF0q+7YRlZfdDX8P7Fe+IBz8/o7wR4XWeCDIWli6PRKV+wOb1JI37rAFYpNtp5t
6v5LToySj+lwUGjIg3FF+E0H/kPM1EAB/nj1msrdN2xAEKYa9p38caCM7VfI7aEV7W4/J1+P2Isj
y2kiNg64/1uhN/SA0HV6DPVeUB0w6hgR50G9M+wSDBJQYMExpMdBLbMyToUM1NcLs3zTImeCJ8hd
CbNK8yJolEQFKzPbwOVJ5x7bh7Q4c8UGNVYY7iFBdhgQPH84oBHNjP7u/eQVnZLPeBuFQdoFms3n
gGAl3vLTsgqkc1ckyKxvsPEVRhrbYzXqwCBTestfOtobHCotmKw5bFKxOYsa+sQ7ew+6RHL7SMGj
f1T+lMThT9TOGBFDnAxcx7leMtcHQL8vD4U82ADi4Cd6OeEEwqsz423dCRvp2Ro6TG5t+93G9ib4
xeipb2B15hbSUWoDHMWiP4sa9XFzOa92a500axmGSBYiNJjM1yjA2egGg33blp3yzKqOJj1145ZT
L4ROMuX4S1ieY6+CxMza9s9aOTcAkogPJhmN63ZhJT1xbOFSQI3k7yBX1y10DFOEnTlsDP2EO3nu
sy1njAH36+yGshROlk2/CN+uZtqjOhLdK7zPCpEBFPWMFg0dXd6BlfkGTUoWI2nCZKHlvOvOJZeu
RuTPN+YoPyIi8V/ccspz+3TfmiLUmzYgDNpS3OTRxdMysipHdua1hHJ9aBq5Wez0GM+gbAnfz1Ok
Ej1/gr7hNFFl2QySbCTYaiNqlp2S0XDcX3L1eN56W6URHbLdFnGTYHdbLpdidTe5ia4kIsmiVHWl
bfDKmbBCwMKtKdSIlKgX2qTYuHNGEimZj0Pf3Yo0/qnrmwYwXY33h6pUXQjdwAGCoKSlEXXTMjJj
ytkvdCL5ZbvbGfnnYSd9R82Wog5CD/IMTH0tDbyCeV7BbzNTNfp0qNMr1amse9lbeWk8V5O4qVRG
5feF0/O8KqDRArI479zncwvIF9srQ4KRd+85udmfMuwNLEDpA4v9OCOn3iv0vHo9zdB1SUIq2Xii
sEne8IgiEk/korEk3zIlJBtRCXcX+hgla5Pf3wCpyk76rdJsSxiLgVRpRZDyQVy+gi438x5AIpB7
u/8iUwONl3uPsAYg6pHslTU4oW6z3aRHPewZnktan27bT3mihQv8zA1fCyw1aTyYH4O+SFWWOVgU
TFERl9Ph5uXelIcMdCd/eR/2FnwyGZYS+qz9k4baLwaXk231Wxvp/e28K1qa0XMkFIw2cNNsNDLO
rTSKQS3z0eFWVQkYm85NA22WP9o8H4Vrdke1OKiiTZ3vCTy48UApvrg7XFVvHkX6AAy5MEeQ0hoU
2KGkYCGXM8QNffI8ST9jSg77wHS/1oQy+nkrUMMgnjYrPXKFoySbh00Kv1THYYJhqKFwDxMKXyro
7ikYP7+4O5pB5ur6lI1rFZpaU8UTIbDBFI0PfXI4fFxt/5us3l1Btqaa1bs0CbdCfJgbVdDhFuj0
MkDfExqO3Tbm9KsxUauciVEj2a6yL4xNJ/58EA+026n9ylnDy/K+DWcZviET4L08U18eQhUJ+1FV
t4mP2APN1pILlbeQkCIt6T8ntK3oeshytqNg/N0DxLB+wdVCaN/mP5TeiaOyVeBgjmONgd6KQfSo
pW4Yto/7UypGDoLIXXEpGB56yHMr2kNdTeALove4hLQAMKHX8wv00sAj9Xsej5TngLdxm2GXRiSb
/NMVkHa6hW+a43SqT2fxbMqNFGAQnpIsrOpubMPatwqYPHsawYVsV1tLK7WgQ8iEehocWnxpzNNs
drur36k/yG/8A1UxbWeOT/fQrlwltboRGd3aO+XUOttbp+RzRxVm7smFkx6ImS5YEufPFgs4gAdh
VA/UoVi49rMGrOhL3b8UuR+5sZn7Gfg8Y7kqu7aUhVQHm3IGJAqo3fI3FhKRDlmVPVVsJHGO8h8K
lYwNGg1J5qSPt6MIa7YM+JqvqPv3eA5MYvvm7juUsHdDrGG8YIpx4x2cvsG+sDIKz1ZLgKUKbpUv
zKDLNmJr41lxwQf0cq2vUJbyqPGhLrlkxJ9gWN3krB3hNfo6p6BZj9VTFAaoR/uHEXgnLfDo4AEz
UnLUlHXQ4XDYYBfcGbtP5IGNgxPDRQXIwfctPblCFgoNRYYULyEa/tqNHH4KlPyAfBtVynUmAWiM
xSVwDW4uHOr7+343YXy+KTefYPccHXrk9YnJGR92qMb6Hwxy3X2ECp6gUYMpF0agCdAh7LFCydnK
m6Eunh4Rdq+TZkWMPXcNKr2svaYrmWLDy0FicMrUJt8HqGEHbMAXkGsklztQSaH+PkR/N72NIdr5
RP2MqQm/vmiMaCgyBdfrJmBHdGJwyuQqc9ijMqqcx/KvCGWwCywM5oQYzGl0JWwZHedoJduwMbua
Fd5J5yThNK/YHzfcMM5BGyHSTOe0xJ6wSUS0h95g/rH22nrU2D6DFNV6rD9ua71eU7oWMngwq6nc
djBvCmJr8FUoAG2Z4EJ0K0XYzRUMCKSb+5TxRgvAi6aX8xmtwwWqkBSmi4pMvoNrQLa3BcJuSuoi
h82RhT2JldkBNkfErKgLZBjHxVGiKy4YXe346CkRgYyDgo7LHmxKrkloD3Odl2Q9ByB5U3RiC40h
/eKG1XfbPfPwgC/hHcq0IqUgTuAZlqCAdNMxnZdxMB1TNIuKYbOqg48ZdU2bc/zXwhOrTw544UeX
+csKThpIIbxobw0lMrzl/HHn0N07D8TY8QoJZvMKc0nk4rZo1ZjAo54rxHBaBKBsMa17dIWDCkP4
VwVi8lMIRjyGDfCGJwJKvs/Wdb8HeuV/rxZdbMa/aRdD90TteLfW7NFaptkxd3pKa3WN1d6fPw4Q
mxxlmaa+t/YKvEAP69lfx04JCKjjAhXzaKbhJTeTM96MFIeKrCN9eOWlmzUh7L4gb4wwJ4ZPeMDU
tm1ypTtC0z7FL+xN/A/stKVE9MSWiwcla3nnhMEaSU3XAWpv13myGF3xGCdrghL7KWNXREJ68oRV
XzR/wlor3wW6Iz+awUdY2xHWJTXPnE98Zti9gBIy/pfGKai4dcafo5mdgrz2JjfC2h8VViCB3MdM
WXplN+yRj8lxrUsm7ynFz4+MDiGt74k3P/fQx0ZnRyTqufPY/0FgvG78S2iyi7IkuPIEaVo7Qe05
xRPFI4uSWEzt2sDkop1HmdA+u3yPZdDqpcDrCcbm4GOY7cOcx7+lDm6no1g+YVTRQjLxAeYTjQUJ
rXdVy3B4pADqbExA1TySGYUpWwjVmPAKCAmPOXi9qOfNiuz9NBiUXAdBeA8GqZ0AMTw/JdD4UrAS
VF+/2GRE0uvr6D8c7TXLd4ewyxyOF9pqg+VbrJm68xdel/PJg3rL8FQ6LebfNJ8qDvE1fxnzcWfo
e+LqylNoUV2ELEPWKfnZOkeX/QB+1r1Wtz4rubOyJkOdODKEAUpvwgTvL3n+tSdLcCoegOYs8k2+
ORQfBmOjSzhi16Ta6dKGPy4rDzu75sBtMHIQPml8Xw6rpb+s+O6lNqqzT8DlN3hPBPe2n5TvG0Q3
wlJCkZvP3NfqqF2K10GE3ZkcpCikPdKf0nahBb9x4B7TtD6OpYGbwqBYhOEA4bhXsh4s9u4d0x/7
YR9WSp6fUWYf6jpZxec0m6Af/VhJR9rg2Wxhj3lDvdT3GskwDtVPKtIbQ2HVePk4dQwFrqMFpKQT
K+UXTr8drejjTCOYe3CM0HSjO3fa+imRrk7UigvhFfO3F6js+XpNmXuPfihwrxpaKTaeYxyGMcY3
yJSXoeOjvo48xzY7ySFHd+JgFZSc9JChuNZXwCCqvkMQK9FXxBngJuk7y9Emheg4Ahrh5QZHjfsj
xLjnlQtpcLaBpW7cy0mhRSHbMrUhdOsFc+UimjzLSHMdTcHgxd17mAfcYtW/g0eU1BoJbJudy1aC
7JXfOy0sFD8gpr/GFqXDzp/o18WeYQmfPt94E7sAhJdiztGNogC1WO7Tu22vOyQNaRZ54rUIih+l
p8KQ37ecQ07ReurzRJQfuXbNbDTyzszx1MyKFQkD6YBaB3LukmAHQuR8KL/8VncjUmIK2yj6mYBl
2zYeoOpKF/YtGRMX8XJi1W9ZIdE0y+hku/vPw8WXTpcd9iJNLkl/Odm5s191BL5Of9xEoVie1gvC
lCBZ5CvKnBp6F1L8poxP4k1hqish+EmUj4gDY4ZIospG6zf4mgozHGw1gW+mQseosbFyWbNfWDUi
Ls6skTVmWT+R3wo4N0cWGSHbXVsKQIfh2NZtAf+x1SyaW3bHSMHUTDPgsENzEAWfMSj3bxPC9NDW
PP64jBQISROO2iu5vhSZDtJDeeSPVMjNqnVEjqeOtEL+wENAXSBSgV9I4Uafwqp2ouE5W8Jizbkm
zjlViv+U91ILzdSVT9lsjKRnTVK0RBOsX0hZk3T+Dt3GDEmJ3HSzWYDTXvlGqXIRkNnRObY0jbXb
UBqN4Qm/9R3qTjJAfTmklHScJNaSn4ekGXr4OR7VDjkM7nO/LaHps1AiBOarmUj8P5zo1KqqF57l
OCqJLxe2+hp8ko1YnDThl81TGZEJp95lwl8lTBCpZRQgCRnmDcDoyhkEsDiQJbB/JHWTj7auosug
BQxMnr6XnxMM7PY+8+lTRYrkwLmazKKL/F9+FvmTXfkh3At3MfqCEX4DYh1NuynZZjhGeivjYpEC
CxhIMiRr8QuZROVKuvPawXWgOLr2feYC1JJxmPZjmxO2YFfnGOSI1qVY9NoBvHzHx0od0Hy0cji3
YcSJJZyPb3bTROIESHOSQ13y7l6UVp+aAiEtQ/wQMxbBFWSmCUHPCYsJxcIoOpSTuKBaUi8yj9Ag
hi+adUvZrJXBfRWxA6MV0KDQZzojKo2Ot08vp0pckpj39BzHCvjFSyZr7x7ZSSM6rvOlPyvjnFkR
tYjoWSLHC6DXC7dIfwxk5ntL7mgqTWgYJvd1WbXFdJpRBTkSqeOT5ZKv6amhAcukHLjzrSxo3t/r
XQuOswfD6lmnQ1XCiL6wG9yELWnUV+JVQyD4b1XoaUxEiWFwZ9hgq0jQ7JeSgZB6LyK9JbXfDbJj
2hKyWZN2li9LvmhGlWQvYx2Q/LhoOcnx2f38H+Te+V2MUFKd8EoOWkdyy7KPIHgV4SWEgGxJMOn8
bKozI+c9O0kA7KFUCm5KHWLT/jKvyX+v6B2tiJRPM3aAKPZCV8+rKH5c2GuriIQ2+insH87rVy65
FvI1CrLIAzoyygkxqb0/1LzSK/ty9IJcDz0ifoamuMtpLkwrELEgC88qZJ7WmqsbYNtfR1EIdlfn
gb5t3Hn+4IuUL1bS7tD+AX5haVL4c7upWAIx68ZnSt7IXbONovWLymbfZ2Qbzru/QRG0GR4A96He
/pXsKtaiGQJ9Zgnd1aZMOtk7AVJ5wIGZMZREgKSRpPLe5sBJ54aAus3fCDByAYwZWICC6jMR5AGk
h8Rnq4Se73xGCs4c/u2pzgc1lLkeGE5STCJfmB9kQzCzWkMH8OrVJOQnCIMDsQc+Djpn5WYNxS6Y
BfixxMwkSWjqq9vR8M3gZmhzkzdwIkYKVgPKoHWIBszkYuxY8fttoGjR/AiOReKJOdR0D+ijWnbm
syZTdjtSkT4CtwGAPx2mYL5PowqyG5egE43lvru0UdarXQxWdP1NfYv4dgZToafnAu4sp4s1btlq
GkKiSDyQ4az0L5thW4vCZWqwSt817UPxnJ6n/gjoj11Chc4T0jtpjEC9zSyPyjnwwM2RXTadaHpU
wofkvaJwq9CBgB6UPwXTQPHkMxIJzYlSvWcmri/4MiiN7dcoM17fMGX1RPSqjozZo+ulLMX8tAm6
tv1H7FRoiEovVENEj6XGrKqx6xXk2qafqcAZ1DQuo4aNLr0bMTYJzIRSE1HiAh+BBhl1yTpa8V8t
IqIuiRFl0v7ZfOKrjY1/8LCD+ouo+HkcIZSA9YFrwcBgcR8w5LOkjNV+SPnwTFU+PAletFMtez6J
7+s4bEQIXKo+gR3Q1pAR+N9C4cZ4zfNHEJOncl5T9WO9tUwLIAWOILgH8C2oJAEwWS7uun8s9Xjq
cPowp53S7kRQfjA/SvegUAGs4lp6j9OFxVkxoHmBRRIeXhvJVHI9JKUjpkXDgzAtqwEH5iDOxOZn
eQAqXnEuQ3dj1yTVLkN/labLKaz3bR25E8zK2pW6SSwrtOE00kl3kdy3GLa+VPJQIACrs059yAnX
WQBNEUgpLmB7u/9kXjK1rCYSSoNRM7lEkVzsLgNlVTc2w7J65JDgzlesHNBXVgmQEwBREgvbEyoM
AMVZo3j5osMrJIHfM2LsbirgX/d5tMka8Kng2YkIWDoP1CNk2Eeo/mebP2Te2ILzTjvQ1sIw1XJj
wihDMeogd1E0U8kEij+vl13u6T4rr+gfiOx9pUsir4DYyTQP91tJxvWHDyaDtN4Cp0yTBEiYF3GJ
VG7e8EELb94P/LgbN/hc9bVAkcAdGREx95s2EoLB3bxWA62MNLG2HEfyVRAuz4weA6UnPcKOqKkx
Oq60N54vaenZajbnQZQwEo4uly2oMglvzzNKetVE0ZNsJjyMOyPM3kffhUqhOAxQhS5vwvIQiY7P
45V9/4fFU6AlvyrE2MyoxnOau1BK/5ZI2ll0oAfwAdP2I9oNNL3PblB1+DoFhCduqv608O4bT+yH
nHw+Dkxls3s+CQ08yTiaWpJQqW5+GYTISWpzXCUFHy7z/1gXomwNgAvgh9Mq5To0eRoI6fZO3kH7
ktLpDdGbzLh2scvNd6/ZqNp4dXDOzNuxniYPxKU9+dmGHGDvyknilJ98OyzdPswADjsiVx2Ht30z
j2mtlHKDp/ERck9pAeicXmFNVWjag1vjBJ2NgpKGYv3uO3AkOGTJEk3nELC2Jr3ilWx1ojxQuUCc
lwjs5DHMPA5DgjMawbxfFNeoFbjTVARqkg3fxVU31csVOKT/3ewyJe1OCPzdm9hQYVFip02fp7dz
IMp4nVz1fRSiIn4LwbbM5oLMkxvexeSiQGIQbOb+Pu0cLH4+S2V3eHGprIWqy56+rPjCJS29to0P
TAZVSvxa4ccLzpxSkDPZRYmYJNl3KihEWXYDuqhbfXaKPHjAv8vVX5gQ5evyRI2qsqpd9V3VeYrj
j8Drp/a9mitc6YzMUJjQ39QC3v89NL2N1Yx8yZpmTHF8jdW6JBbwK3YYGqsMibUFsDO+JQfffRo+
HWVj6nOH7VFSmtZpOnbSs5qnDm3soxN9QwGBhz4eqw2xUOcy+6Qj+ZyMp3YT7NXrGYtz/hpYPVjp
x2WLK4gl88a+BvZciLSQWZyA09bxIYXvEDfB80NV0AuLMVQQ/cNxvc2+fohJy5v/ZUGJNhFDwRm8
/nBI79J9yyyJZzzDnS0GJGzI/dYdL9LF9wJTUed8oqGh8H1KxkTCrZB3P9yD19i65pIPi+buddBK
s/PeHW6BRpUt1yE/YxpsNdyaCrdPszsLmOm2G/6PHyLOn/SDO31R2zuGxiCDaxUewJxNgVJVjLZS
VQZ+1WiKQCLjKLdwR2xLeoeNLqizaYs+brWJTKY8PqUl8HDWfweGxYKbku74qiv5PqI0EoUVMjaz
Jg0txNK/kjQnMufWfJUXoOA2Eon+qS1fb+uz2RZy8pSSgYMdE0fucGD9qBRp7hnA3Ve7sipBHggb
YHxbqROFBDiikoXX/8VvvMZEVCqcC+Kj6UYC8KDm3ET/xNAHrk9+FMGdAdU7uTIrFGdPXfM9DX+k
d9aYwIcvmqv5T+n36N/Zo8FmSLHlPzHzXrgkCofTyRON+DFTuoaDwq3aV3p7oqTFd7lGi4ikeNO5
M0Zdm6V2bezmPQHADUFg+UDiS21o1SquvooEb9/oxiNH2pmYcFlrkGD1ss88FPqcxpPNvmx2GNZA
1ti29tpWgWkv6eXaGS691pry+W10XRL6Stj1RtBAb8dwb86cwIuW8an+fcRXwQMS7eKJrPi/+14o
GsvTKm0Q9cK/gxs6hIOtPDwkVvviVkEfHRoq4ipkTCSBurlTbpmn++ZzjbSBYQJq7QVL2fstCbd2
6iCbnY5uonGUG+rYpDZCNVPv0QXSfaS0J9lBSRMriYw5ywJ7ayxOUGksJ3Gi6f9Qb2pW5j4A4MpF
GKJRKUrQ8K9654+zClfK2DreO8OuKNT6Gew8mYk90OEippfSYRaG0t5oRCQKpZS3kYfSzMOFvHJL
b1jxX7P5QpLf1elOHL6fg1LZouegHdiAcx9ILR+umZVT1hoPrQLw7by+goJsMu0WJwl0VyXonjBd
Hlr9FXTjZ3Jq9w3jHNTa8fKC/BE5syw/u0tNUrzBzFxvDri0IprH85aMiji6/YhiaUm7esXLM6Z2
DaNPUQrT4U91fCNroaMJd3WW/BsgBdb1rXRxQjSNFiHWAl2k/j8ufGIg003c2pvYJ7QHKdPwKZCi
hXawv22LSKIP5lI50WaQmwMT9ShiPmmMGpMNRmUa9z2t2XbrzhGPEN8yBg5anKSyFW7znrFL7JIW
r2HBvX3DcaiO4zYu6uBtyYqcbBN8bN88is/NxD3tEiHwgJrGW592XeXpXWhGqXoHehfyCw08xpiv
bakKkZ/zBCacbN753t4M8xOPcXLYCwfJv4pQ7mkrnppg8gjbMW4xES5fUv3QB5bCqghh1m028gwl
zmWWdtWhVjv/gKhJga5M/Cn+XcXp7muJ36LtUn8he5jypBK3fgM9zCL+O/tIP5n8Odne4ZRGVAAh
OnkpEi9n4h/W5LmLqPpfmHMeWxUcE5HukjJyuxPfmC+gw8CVVDxbspgNYs2Z9tJLM+JeqJ65g+8x
nTa2+GaJW9aH0WYQi3iDOh30unNdKDlAnYqx3q3UpR5k/g58IOH0VifxBqqlwR47wy5Q7DVgnPzL
+UkKjDZevu25OO+PtndJetTcDe6+gyoHMcpE5gh0mbyGkRiRCvGh+7KRdeXd3aH5S3uSZEAeXkM9
fgkYf6vmSO1Vz/vqfria051sREQpmcmJ6VIX4OhLCZq00ITVPhPATFu/BApge3y2TaAK+RMEMErP
B+3uSXsnLy1Jj4f7EJQN1ateiIUXlWP+XEmHkjrc9L37xFYPCaSlXuJKU8yW0lkrtdzxLig1VJ3y
hRzbMvCT5rhMPbyxhfxkiJJe7N6gPiKANarLL0MwnWWpk/IIN2XQbx693kyQMo26P5seuyzD4zQG
FBUF4hzrCkV/SbYnpNdd5rYZk4u6FmUx+UBmEp8qI9NgC1GLFBaMQTe+Y/RhaCwnnOo1qOZGlayz
y+IYZ6PB8vclfpCPibaCli4J7K+FBDZAewLzYOxUeAPMqM0KOANXNdWMM+L2Iym9VinqPRuTDaiN
jkzSu1E4LItLwRoPhHTwMn8atQeA5aMw31pyGyAI87U7PmxcNI1DyJfCpJWlgyBHN2RkEtPOHgWB
eT4Btaggh7TaDjar0hjxDabeVh4LNWA6vjtTeWgHwvu7GnfxbR6eO+YodAJUV0a1Uh/X6NRFGcVI
gJ9aKmGYxoOIIxNDcnhRZ23oOywGUUgpA5i00Ed2cqh6AaEw087dwpagy0Gv7IvL+uwloHLVVxxW
JrjahveyzOK1fDlrB1L0eA2KS7no/PJlzSk1IsEUerExgRk6mqN7U6bzEDHI9ByH5mjvOk/PUmXx
MqqZxwU7ZkqWSPDGupUSV/GXvP8njd+qWcJD9yvunM1Bzclkn8Dh2LZJNiig1yN8l4ESeOG2gw8X
H4dFlT1xoLyRYAKprmVYssAc3Pn9cR9lDczpMIVerqZzE8Urn7YEQFRIg82S5y4OkLPTwMw5wtP1
gTKlxUQJ/lmcJuWAPzIm0W+Dgjifh+St9SuBcL08T4MzgP/pZ972+WvkbH2T26U+u5aMvOGddS7e
ESssKU8bQBl8qcFDxITNVZTHUAcVqTt25awL0gH69IKr7MUU/QWLj9fAPHuh6DSdsD1tyM3sb13C
uatujH4ZLBDR5whbaz7CF+hK0Ts1qlz9s67J3yx3c22N3gWCh5ggEfwhX4wEGYFKEw4AuZh/3v9c
wDVeF7nLc46ZYM5eRmndpBGkZk2aJMOr1Y8wEdVJZ4MxmyCUxZ88wLgi+SzZrvuuG3Bv98MglEX3
oklXzOzXlvmiFEMKkZ5UStRAvqgMYWB5aE4SsUTWKEfupbn9GSHsfHT+TXkmAVrlMozLxLQfLtcA
bDRGTffCe2qFxTIbjoLC1POJfw2FXcxhLyDiJCpYbLnbLQxUe6Z6k+EiUOAx4Y8wcrC8FI4HVk9i
BlWBH/dCw7PMEj6K1H0xYMOLpn3+JBap7+epRE1bNC1vF4fgZJIOVeckZ42wqpwhq6wt6xfjibU/
aWfXssPa/3smGYVCh0PEnGPbpysskTzWnHXm67WbSata1bNBibopjvKjJtZDcB4WRFxs0ie4fRXC
WHX4xijj3C3pYg9a1sylJCACMX5zamjHEbMQ+esbV2sXTfpG07rRcPq8WIl0e8jefjvL9mBZAB31
wYqkZJyTwqKGbJR2SKkgd65ZjS1qY7/pzbO8CTum+j62EELhLLkorj2C4Xxh+EUn5Bi0IsBMkRLT
M83jLfTM5xl6Orc/PPO/F5ZoMfHshTxemm33mPgOAA81Xni2jZvxl4bScadZaT5kernHUNfPSTPp
pJRCQpp2nMf1yS3/tXdhJkPRlxKZLfgkr8rWevM9ZwBk4u00mGAqgaOP2KD8d72ePFQePmfJUNa1
zsZ0m7lpU7V9Sl1xWEjBCsx1PfX+VnC36PBUFnoZsuO35PVrbCvrwzwilDg7t9TE5fz2faIBT0xa
1VPu85DgH/pp5raA+B7zUzYQLlHIFv9upFfeH8gfnNZtV2cPhGcPvIqnETcfIgGCPDgXQJgM/69b
GxJOBqhpro6uEAeXlCvE13MbLWAUuhqJJTi3yn28ZJ2Xf4ejXd+2E+/w9KySxICktZglFDL7QmEd
qi9SG8Ya0OEpqrxTyTXY4iweNAVo8IuUCNM4052ZAt5QNghHcODue6jgYhiwEl5NxxNzq8Vy3L6l
MtYTseg0nzTvNKiYfUK5J1VXWQ1wUkFizzhISuGNP39PUa19xsHWKaCltTRdL13kYK98wrxS8WHY
qGq0U1llAg3amqXtlm9+rWMcUdSVJRxe9gboHvnde6yLlVphLvw5HWw4DFBALxel1inXTWIXxtjv
oJ/HobIm0B9/S2iEEyHMotUmHKnNG5LJGElq2WHeClil8321RgIp0SsLdSn1mfPyw/0PBDKcWbSx
zP2honDsUk+B2Q8AuCs90HVINHPLlAPAcOkWQLO7JMv0Y+3WwfvWZ81YSYMA2AveTayellcqvTb7
1J9ZyU3hjfFRn30VC55B3GkxI0wzXT9BcJYGbqYltMKLsYqcxSkgC0FtAHMFpG9VOFFoIfHYJ2RQ
QQVBC4G/aOjPYNLqhpbM7ic1ieSeM8Lsy+n/n0/hpuOaFS4zwRgaWDtE8PJ2gWQlUPrFncsstPpH
KOdsZ/w0k+uzEuoWtXFUHtP1/aPAzkLBr5FdiCeDDYgTD6rPBDxd/dYKSCm4JER9ZnSpdFIDuqZS
cEXjH+ZUA+VLBt6L+o0UusT1rASDnF6DNypBxgocNqKGOE8uPd/vUGU3S6Z4WzSP19yiAMfVAPo8
HYRcoJFeBMRdjYGjAW1mWHAQXuaK7E4oVjSsvO68A02PEL4TOFi3j+iKSUVxnt9EiDqfxkuYrWA8
lxbwr4OjfVLFQE4o588ie7TTCeeS3qLMpyfoXL9tMT66ZE/hFfAjH6dxBOUolzT0snI1Flr0VtXD
TPl+4NA2JpHgJ7+GdH7Dhy5bllzmC0tO3dEgnQebFvzIUOd737HC6YUQpotJGfBprDyKX3gmXQ0Z
ixY4KOHnKuR/8eyLetMz5hkYxPON3BPntz5gM70wO+EMKC3eYiJIK7bT2hMAeK40z6FROKiMPXwz
wQvtcfeFwoRHCVtvrNkak3lDqCob8VxkbEQ0wkPDrFpJ0UR3pb6+GLu3RcfXxlKX1Umjc5uWLZVN
gE/kF7EdSDFqOxBztmfxTlL+S6PYxDuRKXCkxkr0e1U1YCFUhnE8/pxAHaXR1w65z0ehtBUuN6hQ
d6xY2rSZgiMabsRO7RY2Q5P80qWqDVRSATUW
`pragma protect end_protected
