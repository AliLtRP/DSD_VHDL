// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
l/lCpj9w0sIVy6ezN6aqAKZcagufYJsJ2G3Rut0cTENNLyZo+xJpLXlNLQtO309M
gP8ptOQlJyr6sGU+RSYk/eiN1DS6MrTM4aEQNP3c9NTxa2hWARQjtDma6CJbkkNo
aVkJTP8IqrEUWXjr3qItOvfVNoRaHNJcc8fR4fTcJrw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13248)
KKWuSyt2mz0/2UoyefgXaVvS05u9Ijx0s1wl7nq3oe4PRX9fjvBhZOie+ltW+lnh
pqodrLC0sI7NJ41mvOp+rjT5NVQl/Mn34whIAY8+vImrul4FLfL9gCOA+XnrRuBl
SQiryMT0ueKXJJhRa+UENqHFu+C3gvbYQ7GjC6kxexWNZtIM4J782yXN6Fx/ci7U
4Q2ITmTrvZNNhoi+vbc/CIsAoPLVpw+9m+IOpipMDliaCKBaIjfnmksdtokfG163
w5CCuGbERIBu3VLn34BI4hnG0OO+l3xjsCms8lUfT3bCkFYue0jhAfXxY+YjlC+w
CIijtnCZHxajpeo2G2pCMsWVaiseoIvTVktUFl3pZ+ktx8p1Ew7XY+YAxxZTyK5l
W97YeMEUIwNXsjIRYsRLlX3oWuoaUu/lgi1YwvfqccT7DIjMfZqwkci06X7FKcr6
Q7NZh03bPIYq6/rbxao36WMycSTMuEjIm7rhhhTl4qta8Pm/zGaGTFzStPwP7WyV
AlCjy0hgpJtvwDGB5jLCsm26riU1cg3LBEppKHKnY4NYSG8H5tL9ahvYgmS97Uj6
dw1Or6M0hPIi8gynAVAKMb/0B/OJeRB4JU8uDKqykn2Ec0WyOrQZjfoLk/FQ3pEb
FtR0iK0CJrPcw9taEQcXLs0LOHzzswvrxQFJPFjy6BkDK32NQLqxonfmVcHBjeVI
f4nbYHSgvtC/VA5iTSVCqohCvpQxBSLsTKjXcdfVBojWIwQxjP3tuEXQ/YefYxWs
5Zxy4sTNSygNTWs1Ba31Q89AyHRxI3n26NLdqgBTAYuh8907zHiCAfne9Fy/0SFs
N7E5D8HR81Z/Vpbh4QcD5XPZhP/RStxlHmf63iBrCXWmKzzsO/mm28bQxxzk6/bN
uRN6NbG+WLRrC1n7JaGvMU+thzyBenHhareWAKX5Z2n5fToi9EmfHTZWz1nheMK+
ISIU4KxisHh187urbQqq6/xFuP8wXa068kVZxX8yCzEs0WiwdjvcMRem6BGVtd7j
yDAkSp/AihopT1wv8Li0mH7oz43nKHBFD3/lUnBbw0kcdYi5MslfgYq+96m1wZdC
s88uRRAUdzawcJFFP3oA/uZIdnHDi+dhAitWuIbEBqMl53Axmx0fnGM6Y1MYsHPD
SqA9/1YqS+BTK/VTf5xLdk96TUN5G9XJMQ6gX+WdYVICaJtQK4/7STEtWFXg1SWV
y+oKaBo/IdKXbXPXqcsoCo3x1H0dD3n6jbRJyzlcd7VMP6nxIjTmQAthd2KLWLqN
V3frMMhYbnrEwgOkW2v5Kb25iPtuNylQo/nf5aZgUUIRzLrhH6gJttcT1hwSZ3cy
GRaFsqhqZGA4CYyVD6hwbeqsHCa6blWTb1+zO2bOCmf9g8CXhXiEYRcvIFrNESZ7
8H6eURZgAk93rZi8M+j20xOwcfkFjjnYq9F39aWr82XexoynMGmlBfijo17alylz
KDI7rVJ7q8TwGWmCe6up+24nVnnVdNH12lKFzCMJv1l5/J5UO0wWSKyDG6hp+Qd1
c/DHdj/LOsTmFEB7nJcdYJg6AdSI3n3J1bWKu+4Le2RvzAzxn47nNvePd9l0OOd6
OginiMvHKsnwq5+teE9f/FwHvMhwURgl35h8yxFr4/yfnn6eg6ObJE4LtOZLXNZ6
kSwg9hmmw0bWtMFuAfcn9EpJ2CUx4aokLuy7PxuoGvr+R8itrfilD8uqciRyPLP+
24osl6s6wwVRxT4FINVLBuFMr0hLUmEBaXDHqM8bWYiQnh78aFjJsGEieNzwTgxa
tJpUXUG65qMf5y4pQAIvMbdi7FE3Qc1tGBaHhI/fOXZHrraP7tlSTixxcGphBx9c
sDbHSyCn1OhVa4NrXL4GXpY11aPRvLFMkx9SeDwYuPVirCwo1kq9uRH/NBo8Y3SM
pSEjSusFmzqCW/f54HwUW6AvzzrMgcidZhxaw65Flmj6C8GhaU1PoRwhbPly9zh3
TkFbp9Ofh0LpgbYmKiAXWo15zJDy6JXqn1yhTwwp52BdvA5EIh/I9oJEi3H1k4yO
N7W60tJOHUTJeI5DVUH6LJyMuDpvvQrEfSHPitBMTc5ZmoiKOrkzOoO7T9cOmp0w
vYTmRe57AsELp+LI/L0hLGWYfNrv+JVmTX8QRr7Yn05/ayzqpOlFaS+X7EuT2j28
t7Ljy8gP5UzxLhT5YE8ZI0V02rXEOxCcopWCoFxtZmNLClmft61Pg+DtckH/rX9E
nZTL5HsEm75EETem2ugT21m0GeFNudFQftSXWoLQvGv48sYK0Cs/vIZyYsgxQ31L
f3e6CN6BphSOcvKckmE2QjvXk4j1HPFPd09+sdRJjnPQOOl9AvQTaY1bPhh82sti
XRzjhSZncOKRkggI2x3soDSAwdBV1FTn+9e57GgzLqlKv7TQ60otO9S5YGCWllg9
6eqtHlsmBuhuoR5d4mZJ3DjlLSuqrkUXaTTpZaBdUcUA1X3JPJyBLLN0YRMI/M6y
fvtidrEOobONjTeo34exoTbBwdlmtH537aOz+vz83I8i2PxBmx7knWb6u1xCwiz/
BAlNJ/tOn1gbX6hcaJ/ZaY0rSRpryyMQZbUBRbujzKs609b0Zr90x04kNycUpS5O
rQYeoTjVyHeE7nMQVwcuN/mAd7MN2sUc0IYXGd6nPVpqrnM/5wtnKUA81/oag/5X
JvTpGbtURGD8eyMBiPxtGIGJVz4+FjP9/wVregZvWEEWhyvFmTgC6nkiPaPVE1+B
dMf63lO8ps1NBSwtSjYBAlVDHDtTSSJ2TaXBqloiuROAKpqtv9tye6JRh8nRn/M9
YkbQ4IX6j8njQM+jOZjTLQNzo1kdJ37CLYQrJUS1xvjXtksBiz11V++vGeG02Dx1
eFpNDM6ZzfoVSi0aT6MctTmuUkyYey8rx3Hvq84kyY5ql83JVcEoUwPP8S+LVKCt
Iiidn+2KZycuNIgMQIV2H4pUThNnd2v27pLAg3oEwpfvr9LIq+30dvBG0qm//rBH
68nsCyPobpUwvN0lFdN6v0zL811XuDwCKxBv4jiITaBChfaJsqQijHa7imscSDu/
5JiNPmcKS7STLeNMc2kK8xAcj12QeaHPJd0zpCTP0LZAe+rX3R5KSVmA8VWIbV2T
2qqIdR8FMwmzm2LmxzP3/HgYyUetOB/eRUWodnIrW72FJWT4lYZfCSGOXHfEHdBl
RiedceZLlqs/UN01Tm5Zralw76HdhFfTayU+6vNUNMT4VeVlWuRYDVsQRoj8y0ZO
XzI28UvKEguTcdB8pC+nhsNLoSTLRMstNvrB+q84Y+FdjRSurITlrktu5YTV1Zk1
3Khvv7Wxdha2nsRfLFD1Ru+Qv3xB78yGaFxehEyAjBm+eYcHmZW3JKnVa6zHzXG8
IMm5gumNhbscDAPMdRtcfzyhGiUzU2fJkNvFGpUtfZ0OpLZDG1y3V+j+GIXYIse1
ULFKTc37u1IFiWEnGOQdtvSxtW7DCAeB3MpW7glfIqErLqg1XU87BXp1p5+rsNsD
Pl476nHufxF4mCeq6+UkET/Vt4cIWwH5vsKQyxR9GT7L5mwK5QZLxs/wTnJGwHwl
sCixaPpGn71kLa4gZgUYmBelqFtQYe9dVO9Ge2An58vPNNd3PDHee/wigoVgVO1y
10MauxPqZBV3AoTkytxNyPu1NtMKEyEalv8rFUK50gOoBDNWTkV89kHYHl2Rr6se
1dvtsiPE0tAaMEx+ZC6l0f3hxoYf7TNOK3FwLlJeKvZpfpCvVbnrJURvw+1iTZRx
Lp0PpGIbAKAakAuYZucdTZTwP5mqGdYQflvotF8hsCwoeLJC9XfS2U7C5nsw1tsm
9v3VXyh/IW3jGHj+Dz7Ga5vnkaHiHe6KunYjeKWVXGp8uPyk1+uw1WkN1tPUbz4l
mSxMIIKoAknNVdlsw9y1Xz9hvjf6ovb6Y2HcrtVlLkQGtwQLfkjfWXIED5q476nb
ASKfWgoYU2qCKySxJFZ1T8qS+5Fs+XYegejE9LvsjvgydqATYvwMswNb2HbJO+27
luJNY2sSlvWjQKM7xe0uKXt3Z5fkcjOkUZWHb+AMcusZBm0e/KtMRqikMpkCYN4d
8e13X+ak8HzHFR5q+w/aiphZbE7AuClWoQRUK0qIJ9cXvtrMvm/A95bDe8ZyvFPj
8jLW1p7EU2HsywjKX4rNJov+x494KgiTjQ9S1m5a9T68JvbBrpgSEvgI0J/DHW3s
EMIA7Xy7BHaDRtPYeFc1hipuy7u+ylgjUGz8E0jlMJ4U0ufuO5ocicD5PmLRUQPa
w2IKuoYyFKAoaA1Hj1POfwVBMxYk8W88H3tpmJBhfvfUx5b9+UJUBdqfsYahnQft
ir1jKgL37CwAGkvA9AA0d5/PJgqpHTFziPJgPZqiW/XgIrywTJsOHjGJcc1jgAdm
ETt0PXxOmaqP6RBjHZ/YF8IZwz0a3wQMEEWmRccd98vT4YjYKgpdnRyCt/H1R1tq
MJeSBe7VcgYrawinmbITnWrQlyCyYD0PNWqMs/4k1PCjjel3AYccRaHBUvZGttPg
Z3TAXIl1eEwmVAAFsIVxp5E+vfD7NoYnWhNJ9BSPCVHVRSYg7opqWQchqdW96j8j
5CX3ZZHcg1ZG/l0+hlfDx2eHHVc2FA65qeS1OWgMxDNfEkKpuO4bNcOtHil56u0Y
iNgNkqSHjCvvvMhiSo9mC7x/nRLoteeuS34jU5FSnyGW41EnlTrwc2elK6q1EVEk
xGRXdWfC+febFzE2tnmqwmiUxVa3zma/DOmfeyXwjUcweIjLC/sE4e8goVhTTsHM
s4/mqGJpVcdv+2Q1pGfLp436iGBktCp0KPw4z9EY6EYW6jbtsbjQir8B//i6w2xE
fQ8/f+RRdWQNerPZ9nvnzq8og0uPU0u32h07MN/aJ3si/NJE4umT0wGuaden9uGL
p/w8/meDdEadX++GYuoESBh+i13VA558jCRBwBdeyh7BH4RdSM5vXnJPY0NHg6or
Uxcsl0b1RtHRc/tQSUzIKZ3yp+0me5km8WNrtajn+yvUn6OX9oHIZD3hOCuLva2Q
KHGEgvmY+r++x+ZXlI3A5CbjK/YhvCoSZfPZxBQNnQlMLlMcAUxNuxZUXZ7+anIJ
YNhYfGwzu+Y/u1e44kLSd4KxHJNDIzijVBofI34K4ZOrSpG/SkPRCFgR1IYCIU2Y
1jW80e8mmxsBiB5571RE5N+EgQDTVj/T+bYMsS/Nb4DPt8XpUVSvzAIcSnw3VWfV
6mFKjxyKAaGwuai6bwAitvpR+jcDbAQnR/H1DZjrzhqQ6fSU4AS8QHawBsYOXOgQ
VIGo0SY/36DGe5wODQ5nuxmLFtRgbAtyIXsLZPVTWTZda4bdrG6WBPwFEIhmb5UN
hK8p6Nrf0oQ0Wz7Er7DIOVDxpCW6q1gdVeii1y0GeW8EOu1C8O4TM88dEx1zlcaH
WzMB8K+UD70v5RPv7plCRyIXUxIgtjtLvLp6i8rCCHdA3nLl5ibqibyZ2oiq6MNK
P/uHKxVv8JFqjCh/eXDLIrNcHguGIxYbHvm71hrB8Dut+inGmgXnIOeSHni8FN4o
QiIJDzWJKSbH6T0E2w3RTsvJsWcX+koCXAC/GrRFAdIHc0pM2ZNQb2sl6MFn85HM
Tl66Kc2WA5KyNyPhzqAi2C13bUATzKrjOLdXz7vSdSlodLRBv1XnWcozfjDJKAdX
hUUVDIBA9IfHTiqBMyi1bL6gln/hVldEw8vn0gsKeNpAHdBWO5miZzuJhyNZO56+
yBnqirHbzJVne1j1e8Hnw9patXNSKNVs4Hm0c+RqqN6TB9NU2oKjp0g68/u4UPe1
b8FaQzNJSCsd7WPZH4ntseZkcxMswrobq2rsFN+yayDnYzCaYR7RH+mEgxSnwIjl
20t6PeFvAeKP+vuo8hcoFddNRBY7A90uhp1PySe7MlHM1DvCQsL0iusWjytu/Iek
i7w1nsoT6iVwWs99QeN8NX1RHOJZmFoRXIlNJTBpGRoRRHCiJ/XEQuny9pDVgOfw
YEz4SzuI6BFA9iEIj2OmPL1KEKkx1AqEHFnL8XNpHVBkFF4+jauh83VAnlEbqu/Q
Wj4xJDmVfpM6lWeUNfwLAuvQ9yFRHnHgStL1EWA6VHZR5FPDxWj0avbF5jFasLTa
zAE585CMuo1ok8azsObzsDE+KLc2ZXOKxlYjJBIAwUriuYW76Oo8hU0lgtnW0ut/
qNrzJIh0jlFMrbGeePGLXNAFrMR69ZlKrkHTlS0uvNE9/cs1wk5lAa93NO+arDVA
OJEm4vAl1TFgyy6f+CvOO5nWQ/V54xk+9HZgts8F7WEeCcDWsd/r8QyN63g3Xz/P
An9WoZ1RdbHLgA9X67/rwI+kRDtMTpyyXGL0hDgvfR95taRe3iEIIosSn2oDlwnJ
hR0G7pqC6+tMhJXf+/5fgoJ9TC1UqYK7fK+yrzQmTCkKj8hlEfg/Dy8j0GNZiRS5
M6sIARf20ef9Jcg3zOaAfXjhHjGFln6NPMTDxNtgy471dPoGL5NEsN941dsxBfIn
Sl3sSfvT2p3ObHRi/4Cw+Eu4uMyUbUByYoyjyWrlao9kvWsQEdfqrFjSTxCw1BHA
tSa+kv033N4rFmRpJMNKiL9iS3rJvxwyrIvQfh59FK8mnkDJ3hhWIsM1eN24tuxK
sS+162jUnwGtldLfFqUk2YIncWRWsBy+sIFVGOrnZybMbt4QPOlkWpgWq/UShGBM
HGSo5qIebvHVLcSaGh1cKrkb3ZzN86ay93UljjyeIsuBLkLom15B6z9vuJPGcfOl
ryrEHz/ABC71QucxtvtnuJLd6fiy60AlKizHHLZ26XdjQDUkZoQl6BvMpR+3J6VG
qi34f18PTsg8wRHVfmFzyybetsAd/RWgDMtkYXD3pazSbcU/4W6bVcHu2CLTVmVm
FcMP2rbyJBHECuoOqBHHNUm4gU1XMRyyLeai2JBWY3oBG99VzrZeTP4fsGHSVia6
mv6lec0Pmt+pNWLRqOOopSv8Dt0d6xu6EnwJA79sMvb9jgQWJWw6KAfJJdH53CUV
JeMQeNIcUou1Tls4xCIF3hpgVYWt0E9EoaH9GIsHks0akFX2GBYWTL8KtpvSg4eo
7YTU16Iv+onqvCZ8UstO8KX5J9IgOvAGpyEBxAQ1P68YKKrVEvzG3IX1Y7HW4XEg
/yqDrVxDy91O0YUEBIeGFS2ai3L9D/Mn0MjayscflILh40yRZ9dOt7kYBfqrNXU1
YTgLYnVpOAZTKPJVrCzswPO6FRhCZ+D2L8cbyxys4LUg2NDFl2p8VQYPYeQjesi5
TqVwgwUS9ErtZANT40WXly0KLByoANcjZ6AtDaX+Vlq0sxDTf+V8dC7HFvtQEUoD
6xILwOsldqbM9USYz7+nvdrCl65zA3j166I2xOgDcn9sDoRoIp39LHM/2JdKx9cm
pEfSdNbE+8Ea0Tx0CuqUI+v3bC8wBMzP/GQU8afVF2kSEcCj5lfBSSSZeiznv1Ph
tg5vG5v744gUEsg3UDhRI3UZEiAMYcOTwdkUPrmOWJah/8WxI0Ncw9UuSuVfny6P
3tIt6y14brde/juXcRtXV4Q13u50FtVQ8y1tJhlq2pis7gVHSHl+TN6LMCqBGY3g
ZZeFU+Z5zbBp7XaWmQA+IYqimGZa2OjXDQwmmPAPYBs2XLN0mjlSu/NzoLrDZwXo
cxuoBFLWBz51wu1+yUIUPeJkbYyhEoHcSQWrfjo8nNuNu9FL8SFCSH8N8WTL18DP
8c752B5CulHtBfX41wgSBoRJRmOpnmmeA9HSQ28jBB550UMDPCwr++sKShqkY9ba
2SMpvFkgZ/mGI+XnVqWDoR9A0oTYClsjDASnNZkWwpoDRERHtgogIccW/+bI0hVd
w+/TOWAS6v7DPwntaQkSX47ntkudheAK3olvrGUScwqFPQJ5N0Q4+DW8SA6bKOft
Jqtm5fLD6qpB8nT0vdW6kn1lJPujC1IOBIdzu3qOxe99q/P19Uq6H9b7EyLYDNTm
2X7XmHlmEvuElCx4pBQCNA0b+w8HcnuAzMmcLzJRzdjds4mtxXqWb7h49qYNi5V3
L9nUaGrZGx4YO+PWivFlLuLPrTNk+f4M0gPVplcN5K5kVPjBJORg0+bI8S1wUC0Z
gRpKniPXyi/Vocn7VXol6/Rq/p65E+G4NfprgHKW39jMdCZ+VIjjmDS23tPefZZf
jXD3Ak1QMAaWcJAxAywJ1SCnTT/iJ9LbJJAAxQwWWfyFpLyn7dN5I85IiwnVDpVa
Lu/pHLrmoq+jotm3J1dqhvdeuKqOvwX0KMVekCIEezsi98gbR/+alo3yh3rD6S+x
qfRjl0IITJrU3vyyvScXjd5onKwmwQLFjjcZBI64QlgibU7tC/e5ClwFQ4G0EeTa
Nsk/0Bd2I5Dav0YUE+cV4OHWj5ekwNmJPqPIzKYQzjg/u1aeOVNXN49oDJ+Gw1sw
7Y8ieBNvYoH2eHN5iSKUpwYJOHbDbuLZFTR7bT/duVWSSSqA2XdnsPDTmZwag7wk
QFCCN+uW6fSQOVGocIwC8/IPFi46FIG4slmKWt/QBHQCZbK1Ras8psqlNw3z52+j
k893qLCBe//08D3SOVUqyWP95LH6vF6Ysrs9zidJTg8hTYCV8yQ/vhxGmL/OeM2s
W/Udb/w+/nxMXLyx17SpMzG5xO9TkLkspvICZTU1TYTlspD0fEHpsTiV4t8GZ+Tg
lKQKedfZOHZM2bbhdkXkhAdxGfD9QcDWALxwaIDmu/GHXqB6V9mOQJgxZ1LI+uUw
4guYlAALAnN3JRSr6Nm8M7yqhbxEZxZH9f6BQS/baJMoaJ2ch48lI9VrWFKNkSrA
FLztrEvxzxZdJ3EPmrd8RthHkFLfeH6oHWKQ0QNKvaXjzTAVVPEOwPMJNCd0uxCb
cS+iz6krkxoxipixgF/9VCH1nBtixpsDi+SSJ2sTtQSf4ai+7A+4uAOhCKP0z2yK
K/TaqoQ5RsZtDQgnlvIw6CN6TGwFYmMVNe4AeVno9McCdsVfQvKhEsc29tSjb9eR
21lA31vQFP+9CG113vKl4PxfuYUikhiJpHsruJy+OwEYnaNQUSrbapJUyzOTrSuH
YMzOqRGjefQiGG1bEWtfyruNG9Y6dAtB8mHKJN2ewrNNwXyQ49AEGOq6j2oSRtCs
3yAhNlGKlL5Uj7yp87zvBZPMtfbDTqis8Z8RJu09NbPXo1/JR+Kvos81lVSmK42X
ifKMJSBAXdB635uDtgziARgvi6ppO0AeD1WyF1418rID7W3HxVtVfwmojNDZ4xxV
C6r0L0Dfsx9AJbh2m6lK4lwu2VoVLk4lFk9b91+72znfCxm/xoDqdB8SO5EKVTYz
lCMcplTtoQl9TOb1klJedgaCYRbjSovuRauvnan3KWAg/XN/GOfYTek34El2+YQe
UUEXa7celhRov6KI99YGKZWUOBuAb34YjfoVFMbjcZrf9Sq5hP49nO9M1PxF0ZzI
OiwhZHEXrfGj+JHIVNVOGH72/+yT6wSJ0eMvD195Gwn64il/9gfoLHZsbBAHnhBy
1FP18qs6sJniXx3cYmGqhbogRg6hvxYno8l0sXTwvZiY5REtsMwS+lxIf3Aq+OuC
7Sqx7Tmk5WJcLC61ETH/6bSwDab8/yGUyXI+lzZuqwveHelMZW/KqrtI/t+Usj+B
7LlcCKd6HbCCb/aXw8Wn2jVx9iVRe9TRCURWc4ILFHk+76fDCTrvc2HgX6+r35y4
RM2tPvI/H17ng1JCyUwGwjAL1xU2kNY+qoLRwnOr22+axaBVBS4BFALl0VItsUnM
w34MNEYvgr5zgwMKUuMEsBb1WxbyKb9R5x+iA2cLzc+xyvzHxDQxetCXYrivoqYi
JujQ8V6UNUHT4DanItyhxUBqoMnTppESQjdFm8+9Mb6lyKefSCKZoUal3asL4IxZ
lOVuVH4Cf6AS6/LVPjQUrfd50jyJL2UnaRR2aY563iakAfvxfQxPQSpzke/f86EP
yIkSOucqD/VbJDWm/jQeRaEY6wnDrQiMV4kf0EWuyo4AdKssyohsWlSyNwL6+TUs
1iUBqg1PEcq2NJzdqYjnZFH5lStpsKrq2YDvFDwPr7mGMzu+Z90c8YiL1joL6X/O
oEwxJQbBMl4kjw7adX6FZnppJzFPm6LxAXRzYbBxfrOhu45XRENNoLzXiQjf1XA5
1tsvuFXXr2sfELubaWmlKStU7Ugc+TFT6+uRAzYVnGOAFswKaYe3Y045fjAZ80N0
gFj5aMWgwiymkCcwX6sdbQWuEm88RcFOWSfSfXlagX/LcXnylNXrT05ojbESvmNl
bltL8kbGf+7PCdHH7a1Dv+3nSptbNgcNiqtcBTQv8MVlAp0HWzAh3pNeLXxk69n+
2fE1UdgGWIU1lOJeS4ImNg64yzOejvWsB2yLaaVNUYZJWbtVvHaT8nlNk/UprOmp
LGH2HRl6EQnLIcA5KKg/J2oi6kY/TCHsP2YdKbinpP20j+lfVcauOBa/XVgT098R
D3BlUKysBpNfGq+7JMIM2yX5td48m96yZRWbWZ5gTcu5PYr8ingtDHm/C5/kuCcq
mfvSnzcO/z9GzjEiXosb3uoonpL8myGfYARD5JO64i6jBASkpF9zxy/GyUukPr2v
TvIu6zdRuUwZivvmqZ8EcT4l3+1DLE+QnKvIKl8z5O84G1CH7mMjYoJEgp++orxm
6QypgO6FnweyM9bXT2wlfTjTCL11vH4/VfJBXy8ZGQCaVz+Ka88YJC+yK8Pbehsp
4pPKnYD+U6AzQfqP40C5c5mo4TcS+/5KQTw3LSJVlmGLmQw2ZdnBubcdsLfTzcU0
O0kbHCKeW5Psf9qsmJDaXBfwXxAxdFyQPcQh3Ocl20TP8ufGwJp3zJJiVtfaJr99
JGkii/NY+RelIZFnKBiiqwOlcfI+ezOHIoiJUoj/pwhu5gWv0lMZaCUOXw+yOh6W
pMEXn5hJ35jqxpjDAKasZMO6l9txMnEy6ivsM2FfJ6eg4u6ngxcNElm/RVfPwteM
Q8BaeQ3yklcnsz+LsBsnbD4Jv0bDm5gbKht5H2UkLhwJkHE1hOo6up4gLRQSnGFb
UYnXEc34uJrM5baAKkqoC8NINqCw9T2frehtDt4yjlRk9qPhvHqIZfVoZLdsKyKV
iI2u+oaGQbiYJbKCDttamWRrSvjIrY4XLubgefpktGRfXBrKU3MhDe0f60ghC23k
eiFcDuQ72v7e/osEFWdW0CuCCVLxIZsbbcfuN42MwOaJG2NKjtGzHBu6c9uIfWVj
g0i3/S1VKTTartiO2MFPbZCbdOZI479FN+JEF3PvsRjpNJxxVDjhwEQeaYlgNwjs
XDpLgFPFGk1y0QS4MgRgfQdY9X14zNDAqmoNSaaeywJ0zMJ9MQflWv+3sDXqXwVI
i4/exU+vpDYPojIjZNqQpwIsPjqVX+f9Klwgj5E7N3KBNPfeBvgHE8Op6PFOkDWX
SUDgvHqKXpqpw5g9GntICoajKDiK+oIDV4qlxJ8m+AN079wmKykaTm/W3omZsfaF
4GpS4tngLGzeUBgti8ZRTTls3UDZi8rzXCni3Db30QusL6YdrjWa+7l/gVP2h6Oa
SSdgozjO5N2IpNG3UHHx5VPmLMDIB416tyNzWKDE6SOWOVEAsARo9xXexi/0adhn
8tPoMX5R2IK1kiUuXdnDWjhgB1PfGzWeQBq900wZP8IspvMVt8sgsjNK+BWL0xqt
ZMgbb5OqTbPIiiG5zwBFjoraNZyK5XHP3QZHICig2aKE8teR/Y2VGErGP4dia1x3
UrJovYaHOHBpuhkZc520l4uC6RL1VuBuerKl0Yl0GL8qgKrtOH5jHlK0tyecaaHC
7GybOdEpiHhYnSDU/Depy6mJrU9bYkerBKPL0DMSgQkefUymbfc+Go2da180llX+
98BQoSpJswcd3R96BfKsPzL5a+4YmNPYXGZiiLJRMv6e7XyF3nxJEqt2UTFp4Oz1
0whANUw4gASeSiIjZaC7YTGfxcsLYDoDdQrbW6gcvYZ/k8h1jl/GuFXcE+hli/qG
QsVudc7FJvC2oZ7eo4rupo160lK6FFtLPfCZEMKnSNg3N3yvUtxm1uZlPSgIsa4x
6jsZGI9hmFOrJqLL7HRKssEhCmubW9ZaT6W+SgT2XoLvTo6x4nYzA1/vfgl0I8xc
TxEce5d4P6gFAvuIRZmU9A08kagP5Mk2J4eXv47cDHXzX6XGaUceW1oZPMsEauLh
9GzD1zwOoFGyizPNn2pdg3rTUfV/z6s33xKdFZBX3Syvq8Ml/OlzxUgCDMjClj7V
jHWOrSYU2fZCpuhNkn1+W4BF8+UGdVPr8ibBauumf5d0Y0rnwhgP1oajJQQ877yA
big4uHQGf0y1LvLklCK8keYDfXdBSQNjXp8wiXfz+EXeO8INDnC7p7VmnVu13oi2
G3N8Dmp2LMiY+OkWZIR7XnDAWq8KcQabf5lrViRDY0AbMC3n6XXfg+JxHEE0kJu1
8v+7TYh8MxSC4LX+vPLshXVfo+p3PCIX/HlxIJO2/M96g6EUNyMiiwS/Ut/VdAk1
ZMmh8lKqO4bBuyPD1c2HaKuDjKIU7gv+S4rErzmp5b9PJoF4pc31CVgNpUj/JdMT
GfZLvccaPdC/hxaXHk2Fld+jbqhfRoVq+8JLlpqd1o7tHDrH62PxLc9ZqFOHluR3
kYSeWEFruSdQMZ5xtk9OtoI26aBCQcm+1C0jTCJ9xo+OwHVuhPG4VNLLmu/2ttDy
9JKCElIoyrfhO0z0x/DphzbxjNCZbB4VfMH2MdlUxBGs3sIp3mbneZK5QY4bQc90
d6IIP6FWHoCLQ7T3Xn9Mw+BiPBCUsdfw8XOQUl7YN27h/g7jpV69JOKOt9hP26c4
PY1QEMhj7mK4uQ3+AVsV6Nu86q1qkZ4elcb4110zpCcj7+avD5Z78rtLYmqJbUME
zmdmqgqqeCVMI4YX54tajzn+n1X7YPobKtJNFZoLiN8p0mPvA/NZS3roep0538rP
h6BwQbdTsWKoAqr9UpW5hshf9vyjNBFkDWALdBRmI1S1JXp0FzZiXgPR+L80+mdB
XlIjfbw5tOEog6hnfKTFY5ry5gdX2CtITkT6DAl7HH0imCZLco9hPmm3VzMy9lD3
kRZOdCo4FmxQsERehIdvmTH0ZGh0HgsQAB8/MNV+O73CejHYmPvceNo6THmfbbDH
kmuADTPg3LZpyznTypDeL+9OYThq5JOPGy5wft75BC0SHxpO6Oq8OIVfDme+ft+S
cFwy7+zRSI/ZQslAQ5eGXH/qzL9L2eSb3FnpVy6JTcmoZTG6yaORdVhPRBjimw0s
JdplvWtlL4GEh45VpqL0EIeKTk2nCPBSjgZaVW+imdjIVnigkVCoJU2l0PmlQdeV
BzYLdglzfv3c25EcuQZfQMRdojDaV/nR9ZACJScIkfe85jK90rwmi5dn7veCpnPj
8lyxQQaNoKjJ25gVQFlGtTw91fYAIH/shhjB6j5brqNaUTy5fJQEw3VJrFS15AuT
n9P2sQvFoAdhp0bMbLfxVFPI38/lVFHKGh3lkhhE15HxAFbWyq4QmgMwe0LX9M47
37ay+smOENt3QJ1xdkFXWcqGJur9eYUrtH8LcZfpd115vLR/8kZqWGtewnTNzj00
0kyvF8rjFslwwk/gOA1CzD87Gu00BEm4Uu1uzUOtSf1dcvpRz1gFtO+yahox5oLo
o7aP1eQZribBm/lDYhMQEaf5rnzc0FWfJnDZmVii1bjcnvOgz2EL0ozd1qkbJl5P
yEgpQ5+EzvOW2XHZZcr/6+bcAT/WNy0mL8vQPJF7SDIOzKgZNtPaZ+qcZViQP8sm
L+WuW/SJWErFyv02bbsUnxG9f92R//FeTIE1/wRHJCcEPzVMalQbLs/ZKmfsI8hW
HSCuqpmdEfgCM0ELq+qamlVhJIdlVtejjCNRtBm5bRKJ4AXn/1qS3vKbZEU979df
ai8u4vYvkYEyE9qa8Ie/XUzLEU7e59zCIxGJJPekmCw7v9naWjJ7cMpmFZRne7I+
uQqh3KkGSK2ctCUpkT+FRgYG1ll4BP2VsN0YDFU81qDBNfzsDFWKJhnFb4rX6bPj
si9iKY2+9pzE333dNMog5v19XAf3hIA7Ta2l1cOHYUffoQHkIDLg8LV7Aindf/BN
2n6HB6O3pfkYCFVZwaz+yY66sSBKY4hAEdV0FOoUec2MmMB0XkywC9UQivF7fDzF
9h9D3CiRtMQF2tpzBzQZB8z96JRlakcxliDOVU6IGxvwSYHKo1voje264k2S9hL1
tkjxJ0aNj9zsYVFj2fk0SYY7XH54SVSdUTBHIDd2Z7OwqHnwgc1FY4AbEuMlzM9w
2DT60F/4+NFQmB3U7VW+ZDRj+UP5wf17x2p34RLkajDhdxsnxiwP9/rttTE4CKV8
xIwjU1YKeq69jdM0q5yUFqabIrmzTLRbkvSiFFeI9bjweyN7VW8kavk4laVf97g0
jW9ig1nwBJJX2Q0xFvU5Zp5RZ82/aaj83xanJZuj/kxme4hdMkdOGarhloHqdvB9
3GwpZNlUT7mJk6stffBEstOsa3ZHh7kPmVFhqZAl3LfookK4yvJY7pRRlP9X65Yk
2I6s2RvwWBvcYn+WDih+uCPzec+ioDt1WdNP54C351Dv2Zw+fo6jP0ufk213x42j
2KyI/fZgUGcR1OipgrLbBqFTCLWmJc/p1geRvtdK0AtSA6QLheteZh7luDfzjHEO
da87qC/j8h8+LirbOPuzXj2J9XIiSLEe+jK63rRULzhIFlWmjfPS2IkQWXz6rP8A
3+aXtxdozW9D6UU4xKkmpQBfG23PJz7m1oRCWPnZCQ9Ga2fRqAoo1EjriUGVqaNE
k84tDnzZmwZzCvpttbVq6+wWI/5stBANG0zgL7dQRtZVLaFY4J0tOusgGP/vyUNL
5azkGIHEUvN9KQ0PgrGfBu34SfY+/nZLL0sNf6oHqcO0QI8UlDgyQU4wZVamLrjy
aRxTSwn5NzX4PAmuZgA3csh1CH3y6F6v7hIxnUl8DYaTtdB9VnD9BRJQtX0dEi88
qm+b0atPggMfqtSg5SPN8YXJVgMIrFQfpf35gDMZNerJFs+gekkcZBmoc6vxr5Ju
Oi/433CcBUk2xTIOTUpEDbiqj0cHpkLgJlKDzcANfjxycFZSSchx+veoOUmEnlta
O9i2f6/sK4UJF/z98tRZKhFQnL6nigI1pbbrjFK/0xmoYDES6sN15DR2Cx6vgS9a
Ti8++DNwsfhRpoPDr6mDbYCMvvcbCU3ohgC8pHYPBlvYPdJKNEZTEAjpQcOuEIkP
2RoBPBY+BAQC3CB3cwd57ffhKmbtdYch+8VuFCPyCg+fI4H6zRbCnuUHPPidQPQK
wh3vJhFs2zkOR4M2dkRH7Q0AlcbtUSnm4jwZLx3nuLztvpQJyrsHTLkESh//4vjF
wOttXTN7LZh7m2aLrXxfGkG2LnpGEBp1QfrxpQbmnB+LubcQhb7lNeSg1YswFQ32
9tHnTb24RWd5xGSsinlnSbci1lVHnGxj33hk84N2C4ckbqcvcri2z/7Y5Y8FFj3W
XgFq8i4jgL8U5B2gwVqZPHnp31aNfBknyPMx8arADdYyhm69OWkwIG9EOtIoiCSb
e/oXxHKulVJVYlwWkNeUv6ykJbrXNzdTJF/Hx5xyeY9wkTq5FkjUmwwAoWr/mDdt
5GqnzBT/+4RpHOHRlsfGJspapcnngcpc3dgymbMotGCvzB9rUY0hiQGfPbp2JVIE
vlUxpZrqAf53LBXXQQKmQaNoOe+9b8/Wp6gLiP+ZgYa7dGMZZkyj4JQXjPk0AX8y
ZK9NwgVhQtiNKVunqBBWU3r4cQwNfIEFRmYyoYCLwQHyX8/cZVFA9/VTgxuTi99j
5snFRNJ/Anu6Pr0K24l8Djv92XUW2jsiB5QC8DVOTVHUQtrTtQZfno0Wx52GjjIK
+0l4L+yrUMYnfAZUBnX93cbxwO3wCewlgwX4pxK8yXQ7N1s5+xPa2koJ658Qk1rp
hUiRVCqOVNhi5tojdHH0pVhLvFFhPTp7LBmSEG5BTYKuPkSBXkXjEiHKpFmFK+aj
gjX7gQm3hLP9J/C7CFNnisWuleuM9+LTeDBPBiG4qJ3G5Jx/ythBGE8a7mF8hRcu
4wW4JKXXEVp40dRalh8S0aCVH/3Nav/MBUJN2PHixqwTkE/0ycsQkf5I4A39WNon
q6RowWmqEjp0c0WQNpM/kPOiTECyd23aXkXrQxtip7GZN5J+aT9CRxm1jueeqZeT
df3WmONwh72y1f/3Wt5Liusl4IjbP++XE2qk0r79ckdFSbUKF/cO1kvTksY1Eq0I
qwkSKpg6HH6FTUHcIk1EnMeoXKKGzJqmGv8HANS3g4mJdnYg/MzJA7v1qLiBKFVl
TjpC25tJO7FPAJz0gKBXLDkGIb78EatFe8+mOgt8l8jbUo7F7Jwr8wXFQvtAlCx9
xZMKUbtDb/0JlCNOZdKkA9s+HGVld+vXK4q9nswFQSAUodO8kyeBM5oqpRVIr9Nx
qdn9MFimYMtTO93DBmR72mX5k3sXFXKCuNBJ32yth5vVae9UA/vKF2hhcC+RIiyC
Ap7R28kr3r39wOxJ98IPPsVHbSZWdBF6fnO3RMt0NrFTWsora4bQH+MvZPGq7xUZ
2cYbXSXskWd9cMqm7VvqFy94RHwBbsjTsluFU+Ci/FBrTMW8vLbMftHik6fQ0vVl
wpxrFPteihYWdcwojryT3F+dTlZGmksJluLXkt+SbkV1dPK9sd4J+4Q5PNZbk/hW
PrhaU7IHgw8Uf6Mck59yiOd5gAgMbVQKsFH9xwXzxzJw5rcC9n05+hdHwg7K7fma
k8dxw9x0h1+RXd9aWVzNRGiLJ31BbNFT+g7d2/OrRJvgVS0kTE9Og+85OJQVnJUR
YWl7enRVASZSS7ltCE360eB7vvxrrdxGp6XM+EvxWJZ3j5sf2pbekLyeBNYD/96U
wxry1MFn1yxzkDKlO48UySH/IUAUeMG1LI7S2zU/CH5qB3W/QrnYbTYuJBgbUhI+
u9So4kslUlXC+Fg4o0TUS4lTNSTWbaDGpBBsVFlAgPyzKIg/UPvoN3UZ+FAgLVmr
AB7XX36bqH7WHlNYlqna27J+9Gmf8WsyGDuThpFdwi3WPU9bYbm+EV6nEb4HI3t/
sql0x4Q/BCIiij9aiFSq2Afc8iH6sP6J5ZlO1Z3payA5bBnogevt/EU4u1HzQOWH
Mji2yVLR1p46HyOqSDtXPy/6FXyV96a6It6iqGB4blIr6BeEv35Wkv+S+LQIAstv
wcl5oMbj4dncEyX0VrA0LEozS6ggGXd3UZacLN8LJXbVENLIQTnO8aNDo6Yk5py8
ouA+3d6BZAKg5tTqU/AmkGuZC0XHBlSUw/V5gKVcvu+BwfVkHkwuCnrwP7gsehcg
YbGmJDVu8L6jImw7Vfiyhu4OA/rahni0SUjlXQfDnSzhJ/KzSLBX98FCCP1rsPo2
htJjLAvZbrBXfD/mq9EQiwIsyRRhU1wlJwAtg0Qooto+RlwoFUgdSzIv+7VRRpUS
6JBPrJBKBTVTqpPY6W28yttAaFNZZmJHG+WVWU31fGlTmG1hQM+K5XgkAGyX65ri
RJ5wPpdaHbs5xmKUiiQgv7pfVuYsxcdhC5QzIngxAj8paYc+KYFNHbpV9fpmxS+b
`pragma protect end_protected
