// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ock2ofoUqsNYzv+verfrxm8G+QKnab6tjSacoJVHwTwksy6tx3cduF1v/BYsYSQz
p/leRmk5UmU0xL9VuovcU3Sx/X+GH67fX3lPkWAgvrTc8MIjcVLZGawDurz4pCTK
X+rs0lezVV9w3tQYY/o1731PI0SoaUqC+tUb/d/G64E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11984)
ITBUc1mBKGjFpj2FrebRZv31rLO2GwjfUrzJ9W1Th7b23JpJIqOzyxBpLFyB1Jm4
J/BuT/5x8jcPj5xvKdatvWZdA0Fs/D618T7+3trdWwSPoeO3KpO5Y5IaiUEtL0+8
KPGSCABYDo5IW5C/BNq0yDaKvwm5OtTrU8fYqw/2t0okr/HVtHbeMBLr5mqQkt1I
3fn+Sbhxk6GP1Z8c8Omq+rjN0qHUyyLgqLdAK67jkE75sOHNb9P1awkmLCqyJspK
jcH2EiTzPyLuZBfpB4dihmGmd8GgB07D+GTuaC+4T/Aq1TddgIBV3zna6+qJSWyi
D9aO4/HgRLAZpt9H6wzY+ukCsl7JIB6fY6ocN+baBT/StBw+ivuMpFDhUMRcltow
T8Ruj1LHuJLq6Gy/wUv5o6bTxN0al7d7qNp5olcvumkFqbVYWVyTOGb+lqXX/smn
3k4JILEBRxkxdU5NhrrBFY57yC1hwzxnVgjOWQ2/j0sT7K1/gY+YXmkKKHyBD8JV
BGsQCrjrdo/bU7RwZtR0iJ6mmxKJ99JjbVA9Wl9DbtECKXtQgJ+KMruGLKMdrRwp
sSYQ/pGg/hmE1og64qMb9jDM2DCune5pY3NBCnsjoQ7OcwMqx1VEpBTALu7/RTE/
nVkZChqc170CohROm/bmj0SIpf6PjjQeDf2/nE2BvPiGSSTVvcopba1tNy+ysJZN
1Rg93DikNXiZ4BAkTCwbRg4/D7BuePH3pxuSrM+cfqbcSmUDeUlGVPeqbTc0gq+4
hV+6vYdhTKRV5D9NVu+S4Fw+fjCEJlR9hiQRrjKaozQe3DG+/Hu3kkWPQcDJRgXn
zoFgZJLyaKpWStrnBKfQrTzXywhJeTg8+YvhuJummblRq7B1xHRx+hHGVxAzaxX1
E8R1YDGm0dBo8tFgKMhjx1QepM8WgV2X0kGiIFKA8HB9G1hrduwLnXcEi7q7GJ2b
lWiKdR5XZg2Gw7rXVkNFR2xWrZfCw9CAQNKqeqCpt0fEYb4gF1yWh6Mq9ZMR5D4K
tgfj4PQXund5JlTC7+EGGpRGk54/WfTmGYOWDipAwXik/N2ptB3sO/uWVbMnt8Pe
ehiObX5/JGqeZJR/0ZvmqmrVUwTjI1jfEunu96Rg4T3BSf4nAAwrOnXLe6dmaQyN
f6h86HUOArIjStnNCKhNUrVaFzEUqG0PBaAtbUkf+6xV0IdY/DRiMmot6OZlYGFJ
/DAFmJ3VtSC5eZZDZfcyaTDu0X3c/UOsw3NjyPVdqZ2JadQG2mH0mENMxLjiF1YQ
TDV1I2zlmfbxs6WgFUpLA68iNeaOPiclKWwKJAnTwfDJoapYUBHSgDfjaTGirhY9
SeFTRphp60EwCTCtik04s966kzKt6+1clJ76nLwYJVv55ebtI7srjYdskiYuS4pm
XX0cm+WPdxHNZmADzKvj2bXAM3R/UKEpdlScVJSMXyoyc2z7R9wKwz7sFgrogdad
WflwQF3/b+z9kaLCO60cKc4HZSUEFyg2AvRhUtlMfRVOWnjom8HwSgelv1kLHKYg
GKxw7uvS43LEANB9FvK2IT0qshQ3vQ+N9B3fNBpKqUoQfNcuu8XZ+VBCWlzCl1hr
VSctL2nt0W+Yz2RhW2gL/pPn3bbgrvayu62kMdKW9z6Tm3mGXhE58TAeaxnQ7SSL
9yQZx5YQ5/6p3kgQ8Gp136KfmF6CEHBgmWRHljO8dE1JAKm/DJxGQdeVz0Vl/p1b
Ioco/Ka6/LzVNIU+IOnEh2VDfcFMItQ2d+mO0Mw9pKth92P2v3bQFhsAuP6Yb+Kc
he254lD3NcXwuanhjREIMGod4hCHqMtWOqkMQ8FN4jwTt4GCylT6rfjiyIh+SxMz
V7ievlwlRNE3TTQbCO3KAhYl4AHww2Z5jO9lj0E1FZ2XD6wuMH3uAZXydTOPmxmb
RQkFI0whUWi5Ppt0zUKotgYbsXpnuQRcBH3mi9p4/3i797EEzxTg2JCfFoHfv96u
hmU8fwTX3nXI/TV2tXhX9Bre1CLycU6W2EEMexnbhuNHiw8oA+UCv+KaNRiGpWIE
5z2dYY2FMgtcGWetuuGm2ZnTMAPLXn+9lipsVzN4S2TZEA62HZJ+Ia2CyPS58ViN
dih4ZVkOvnTv9o1FVGlRWpTewc8O+zqJEL2Xu6hxKBLA4fHprkWQbyPvTcZz5Sn+
KERO4l8VNaRqc/P5aEJHa01WgU9xnBVPci9MqzYe39jtNcmWAVxWKIKtao619brm
Q+ZJjs9xDSyB5QqcH+2evNTA2AbgCwpQliRrmHuKoAOjBSM/G/kDBpxWjvUM3T36
0GSX+9ftjmsgPCods/shjftRQBDDPAqyh2qpBC3yiHAm6ztHvc0tTS9j2vi6z6n9
WXRXM3pa4aQkUsFoLBqHw3atTp2Ol5eUrxnCm9o+1oxl5eKkHVG/0MUoDu1CHpPs
GkoCqZSIJyOzRzfprouDBVu4w0Ff62QBrjHRJuz2UqXwp66h5O4yn7OGqmg+77U8
JDeym+fuKRP845Je0wbKbAy2A0mq/Jftd1n8ASkpdvKLhAxpgmAFFaRipIxdgwhN
ub25IX6pkfFNiQEgWHdh7E3l9aKcEgKovCWNxZeZTd/z5j1oe8937Ri3QdT4ljj+
0FpDB3gOlamWhRmxTzC2n45gioV6OKCP03naj0E3xIRSZ3COpITUpE9mlBd6M0Hf
TfNsPGNXHHUjdf065PfgtiFynEe/Z6f/sn94FJU3Xbf/P3sgu0cholyIA+mFz6ez
9YjtPByU3KCv09poZneSf3oBIt/ygVBWsojRdb6zLroIHbDOvwnYfTd/2fwTp9vC
vLHF9VKIalzUT8o/EeFoHWS/bh296PY7kLmI4jdVvy3FLgSTIZ4+ic8nlAHglBvM
OrCwi65Fcu2fjl5EXsoRxsAydvTHcwKRLp5tRJCacQK02BG4J63qkbo1lGsvBmhk
ogU9hi/HESUv8+5hcoc4iW4YVvhMolrKSCj5wulQ+gAVHYaMduW98wOfFXXZ60Vg
PCnxtwIVny8mdkyZVK1CQ6WRhU0qTdIGW+Lv5fifXE/SAi0Jql6I+Kk+2m9MSZdX
XujYleMrvlPaAAM8y/NlVD4N9BzBYnLJ/dJBrg8X0RviA5YXZSsLXIKltjNkm9/S
hRyetRQXMkAjuyMWqnrFIZDtnWC13ooLzVIaa2yIeUWFkinSbcrjSbpq3hBAZq1u
ESHQbBv3uxbAVQEHbvs+aJWrj7/g8DbCoL+ddBZ3yqowzvHl6xYvzaRs8IUfkCbG
aO9n0CuqHW3Y0vK1hZypqMTGFZPbgte2dDJXrvLpDWf+uXZMNVxRMOvlfuTvD9h7
wriDbqulO8EpQrSwT7AmD8Hj/AhqpDbnsZXM6Apb/O1hL3A1PzQvnDyC8tHl26nn
YW/ymkcCIoMYLsXG83lkU+Jj5d4s/YBgqPPPs/340vLji74Why4tPOYZMFr/yzZS
Jmp9VfQnHdjafRCgcixW9yt0DYZaVVB67R8txJ5RTpKx1stim7iUbtx7lxr1CwNn
YPpTxmo6KBrdHEcbuVxCXGVT2tvw+iE7dvCNeKvOLuT8/OqmRM8Vj7h+aZJhXuAM
A95+CW3lnAdMgLRDGSJnzMc7l4509jjDP22bisU5LOb4yJva4WmBSwW/ldJjVevf
zfxWemjnhxWncFEPL7/Zs/uNXNFhK+QR/qZY6nAemz1D7eV6DESeUAOVrcSNRRBi
YJpR/y0uHlpDNDci+gcy/fsXUdVWiPZb4uPuXkDOUX371AiwXAXDT/jBRnVXDdBK
ltXdcmor8OfacDt+cLtyxMHS8OP45RkL+2J1kQmj1kQF1llckn7K3G2hRapmNd/K
UPZvonhf4SxEWmYmJVn0lWI9iCWawKTJQD4Ej/yvDRw8piLSD86q+hiiKYHggxUM
tpN7T6uTOSgYqbLiQ4X3MrC6C1SuJkeLFLhFQ5Yw7ohsypEEekqePTM4JBx4hOfi
vDSjaVxyuHxMEVm7g/DYNzsA8UEFAZNVXDqwfFV3ysLiz+opUDNUYbJKlqis3rRh
E4QCYy8v40OKXDSQZcGHEEa9G5g45TEeUR2fQWF1sVRGB/c+2KBbcJImflOXME4d
5rsFblK8Z7MxocdgIpnzoJcZ+WEZfvt8AuXv8QG6UQmqWBaegTx5RofqFRhsWNQt
NL/Zp8nvlKA8JhJXxtBeHmY74xIpnpHU7mWspwKaO/bMk4+sG5FoyhBmeakPqKBR
molkiWp7FKM5G+ojwdLKXMDgbGldmOeYs9APG52p8pPasw2eLtud9jYaJfrQchKq
b8/u67NPpEfMJjevC+sOjL+/16w0VJsWpdnSmY6GKvTMZzrnwWMPTvfk1Flb/2b9
7h6HBw++GwV82O0xKXMymq+xVMX6HYGHIdsItSUM6D8pOxnKVxfH4c8FHnlt35WH
+u1P64cacc62WYmvgHsSGAbAcS4/5pP9qH9c3znLopWzSzuX/plY5g4HhJqK2pqQ
R6EbEANLH8zjgUrqZD9u2NLRZBzCoJdrpL0+8DPMbqQ6+oILu18NsBZ6huEG598E
RxYPJwd4P1o6wt/pR5SKqfuL9HtiJMK4hgcitAPwhGjyXlGesaAnFxZEKwNmxhj0
5E+98tFcBOzY1DiOZFE9+jWKEDah8j4shw5XdhKuYDZ96jN+BG0yDz6DHUwFFf3W
2vQod3ys+m+7RwqfHa3UQmAezxzRVSCknl6mRBR3TngzGWW3gvvxD9m9rhLaFM7r
KsNy1Ss/TiHQxzxQFAnqJcmGLHUuEeUWr7SYIeo64zgElW/9crp/NpaursmqyLpJ
JSvaFZdOnYohX9XNv+T45/n8qtciGBSVPW/+ntkvcX/vFgFieineDffbqVYV8lV2
opYJto8ndocLtmgQfVv3kkbGAPZUpdS1v3wlH0gIscmISDXRPOhcjwuNC1c3urbv
NuszsATZ1CJUa9x+Mqbx5F1JmJXp4uBuS3XB+dXkN4QWxg9UjR1sX/p/JbbgqKyi
zSime5TVzVs7/ikbwCz+VJ0ehRXvWn/I/7QWBd84W9tVMLCP3u8la7cZ2Uk6JZku
JZlD6gJ/oM5OHpPBfU1QjzKTAoMpVT/ymHV+tOlsL2DOswAG0gT8he/5VESZZecO
3una1oqX2tZAbK1ilp4CW473Q9pAp6tCOV0rQclU3oXnyL5gsaHHCWs+vUxFArnM
emPAorETevQsW4xMRtC/As+BXIKnHA5eAH1SnDpcbpADsTINDbvFyzCAJBqzV4mm
oT1RvtVbbSTECNgCkWuLCVoT8/1nL4GyHmiw06z4nrj0L7K9LamMwTy9pNxVQ/lr
87c6TCYppg9EvrVrVyTkP6eU6hXoB6aXscAfRmV13bFgqftXX++70mrS1DbR4mmG
5foZ2MCVVZeWAdv/qbAFv9FRjzRUFhj3QFk7qJDoVnuXjd+LpRBNSkfTKBbWbPbQ
85LoEiqxpNTSHh4+OhnAWmvH7OyTiMCTaFNhg1aljhHFjIfUTpPx+h8MqMjGFbve
xB/yoiZQN0jZdVcKJPkedMMgZx7k5X8cRknvs+CcW4Rgey4/sZurxIZC6U9e9Y55
ofzWsPsqPJP1AJYNuQvoXKNYqg+W2DIWy2ivJioIXVDH8tSkF8uJtAmmkx6tekf9
9gVb0lzBPaxn8p01encFMqm8axb90J6i9qPaHDqxpxsCIyD++fzpL9Afg5pbbjKO
q2Y6fIzpVLX8Gw5fMY3uisA55CpkAX0bd0GfHaY9RpQreofjOH1b2G7pboPdIRoD
v0z9Uw0rPY9N31kW64UcG72hoyRMTGIbvLYvqhZiue2YSCWo1U8owj8+RzfROuDm
QSkY9kBnsZADDii0S6Eks2efDtEMYuibQ3pcdPXWWlKg36w8ZxxA+eAxzXNFEiHc
Z+KYRy4PLus1LmBihPhlhBO++0/ej7DHQ1ZWeWz1FJBTRIvq4j1oTqTgq0PbGJtx
quewAWX0/OJACrgirOh571v90QWWrlcBEJM8ZIeIPbPrORppgA3HiH0BTnZb5HpM
/oSC0MI00JVn3TVcRhVQc3za3Lbrr15xt4oF693LbkfDztj3px0a/Vsm37Cwnugt
GbTdxvrdpRRFjdJ38eXwFpIekdHZyEUl3gLiNbF+U4ORmWIEmk3WqIahYzhajb7q
ZuiP/QVrjRJXe9FZpCkAHfhKUQSrM52xBh5Xa8bIFM4pfXFCzfGnMxQZ/1WKneht
xZnmIch50M8th1OG3YhmvSnarlhf5LPjVHKAXaTd1PhsX71pG4FlgYyEF2RGdV1U
WjCbv46It0X7pbx+u20AQRTkF20UM9bqPN+9UBmqcdSPX27w29DGVJOMRNRhN5Kv
h6hBu8d4n4I8hAIMsohm8g4+xvDvDtAeefOv5/nzDQngYo4Zlryttjua9EgUMyYl
PKw5Yk4HRfA/xwH2uKUte1zQ22cUTL+UQCSfkEtyP4WKPw2tGw6Cf2AmEq+UV8Yj
Rrro0jq8FE5Ah6FcO3Hf13T6DilWFjrp8iYd6qtyok5K5t40FYj2Ak83neMkOyVd
RlZgiBZByC6nRek19LNtQyoO4PWudgYLMzDzbzGHaP4Iovlf6o/7GLy7RXliQXXC
dbQjW8u21LIWyY4P8rpdTxyQNcsxRKdX39uOYFeys87wMhNqQ0PYxTWtT0YhNElf
nsWTnS6lL7izcfQRT//xw5UM8DCKRh7KwAece1Xho5ZfWGjHMq3ulam28x6oJLtN
W5RvMBOvzPPsmdlJvJ5adAweNcElGCz0jY5FrFcXO52CQaHCV9DrfnHXFo0J9W0T
ctEIoJwWK4dGW3QzUmkT38m1YvYZlPld8QQA+l7O0XBSUv5AEQhHShpGqegMB6e5
+zIQc6UBq+Tx/LnOeiIcJaf7skRwf2OVugeoj2qV/3lHE6UTRC4Kzlt/yyjPJGoB
IRRUaLrokkU1gY82+JCGBSpOsftrl9f/bVs0tnhXWrMSFtZbN172QLlGoTglceAJ
kbJ295ZylLIxd9SUCe4wBejkkYfqQHt5lCCBR8LVvS7VU/WqJh8RQojWEUrcJ0Ni
83mApJYrwRNHGT2QMFtwzYWB8wr0/4qBg3HgKwisvDX+/9kqA1EhYpIdMtLswpKw
Cqfl16t3msRRAHsnHsimLYe8L/UoAyLXbGCvax0nGsG/PggmnjlzykFu2CdLo3ZW
OP7Tq7yASVdrdTv1298djcr/4q2ZwLe8kv/Ixjmj9sc9rjPNrexJETpgsn0geASv
93EN3CphYfecsvg3Aj/38AB2IVBJZe78VDYKs9uOLeBdwSlmQlNQj5WIrGs9iGP/
JoUNUg2N+r2oHfpc7wOck6p0itvWMeZT2taDDnFWFshEoFVrtQRHHWr7KTvkcf+7
TVc0aSKrPU6s0PuNg9bCZv77l3xmQHL1qr2OOboHrReJa+Fs79VBbUxWzf+ScKn3
xDun9d0I6vmpqwV8tyzTFcuRUl9shXNb+WXSvKMmMVYMXxKkVJ/UXYS1ZI965NUX
EbCAwya8comffK49bCkIEr2t3dkuyElAUEOvaZxRgKSKpsv/1zaDpcZOrwnkt5Rv
VNKYvc1BmvpCXDkPzakulMvdrWZp1B6e9H62PwueTwD9jcozvJzHaeZX4T/wcdY3
R3sxa9kprrT+GMJJTQrpoWIeiE+YG/MNvt7AqeL40BDY7vqnU6ifwG4GLqWfKYUC
D2mID5Lk97uh7VtLY0+o1UGHmc28ic/9JYzlZIjVkMZWa1cRCl3h0LqGzTq0c6JV
1ASueAUOjtRssyQ/5ifP/U2pcAAqZ+XmzM/PE8ElU1f5ZvVGdSf4h+Uv23WqhJeN
JsUZ2te87c+/IgsH/aRNIWjbRBnbTMlWIpd4t0KINlud9CMOha1ajlGN8RT50Ciz
bZD3zWDac9ESmdowUN2l/N+SFiPBuyDFqcV3Tw7JcJqnVEswiSNN+fmqLdIhxz1W
qLTtxRpFDOmf3Sxef2jvkTZhOi3olvCexaqPfbK+6NFI3lE5eEo4b+Di+sb0k8os
0JjveFcF90FMB0qBkaHre2g8N1tabfmRud18Dhw4/gM1t4loTsBaxje+UdRI/qYJ
0q9nnM65pKRiyFOcimFaX0W4wgZ8q+1RuQJqOUmjE4Ssnk/gFIgNQjReWPi5lBE4
BEJToVhNZCoe6bGQMZCpkksUiKxcV+XSHW05XK3OIjPi3qjP8hJXizv4xdwKfqls
hAzyCcLNADI6QYmyEFoR4a7H8yaHSF7Kk7EnGFbdDlhaGKrRg4XMtoT5dAmfeczL
xCtC0ozAaxMq2jMZrh+GiuAsuWlY8ZNxs1brvKQpUFSbitbBovTmwjVvnzjKX9Xe
qcGBR4dSPj8IcPhHd4+kFKbNhtoDzQVnDoehNLUsF/b5J/sZVfJXcLKt0UWd06RA
we3NvlowSI8n7/D+iDq8u7nCelb7gnfJeGASc3MTPkWuvNMSktGZN/yxKZC7g+zn
yCXSxRfK+3OdA2AqQClsk44gm1O0IC9RhJkzM72K1qWVGgT/sMavKfihaLQ+VRCr
AZvzvlKTKBRN+uo7BvPFJhCny4q6xy0q15BGLdyvhRNt+EJfLYweUb+0dYeLpwbh
QzRKG3Aie1RrCS85PRjTY4MggtYPsShZw3r3Go2BCITtTPXOdQMmXQ4WT5Ynll8G
8VGPey225oGE4EfKYZn9MdRdzZs1UgG5L+hy80Y6DC9m8GssEQnY1wk0uKMDM8gQ
wty5mQRpZjJp0NgxgfTlSTJjfgzAKwAc+PMWvhwmbXVn9F0bHUbXLMglHyqQBG+I
Ucgz+FBY41f9iZSu61b8JJihuxOJozn3t0e5UUYx9f3F5fyHjWBeHma522a+gOu3
6HU/3N75HQIZyqmutwH3J3KvIBmshXdevVsPEB1R6vPh8XkUazYn5UbAMOV2/q6x
7oJ+OpI/4Csq1TT4KFA1f1MTX8Mg8wtcIT1aOLTt3j+KkgzQedKuHArYvEi+49H6
wC6w4f3au7ZC/WrwayWr27ETQnQ9AKU1u/9B5X39lRlIMZwVb1oytuCf4H+VFddJ
lI0140YsRTFBnCHV3RYb27WgYvyGYriIdf01kGbKN1hR7uPvxa6vkHUQEdJ4//yB
rWKF+rd39Oe9KBxh5ab8SWL3tYx86Ucn4aLBIZPxVSWJlS6vxPvfDxg45TufZOSg
l06hHJmHOppTquk+lIckwjiv2ylkVsf0uSZsfZ+W79VL13GKQmtSRBM+9yK/QV6B
4/QFqU1A7F3Yhh+Kurpxl2+BEmKy75IkaHxm0SkfJZxMoDVmEUo6N6S2JQLlxGPh
LgLge0yPQCeoRlR/G4gH8qaWNJ9Eob+bHkfkGw7Z6kIcMHG5LlcmhYl/jX3j4NbY
lpoOiL28P0Dtn8h55cOybjLO59ohK63zOV7TUuco78S3icvmNBlGhF8HHiGISC6N
NsYhxsvMu7VfN4utkCugdoE0G7Qcjb7YMtIuPAO2YQKwgacQOwbQ1KzVcIWKFOiu
+ndb+Yy0fbySRz/jh3cMx9b8X+w6Uh35B8vGDcF7mZ/8cLdAhBqUSlmt/CymBRgI
Gy1pkBxXXTk6loOi/YhDb7MCUvKIQLu4o3eP4ws0lVX687cDt4g3F0pTqKi7fKzp
f5fSa+xYd53ChBiuwN6y1O5JJVd+J4WT+jR6HI9pTYox06JVVB83BLVBW6GGM5Nu
/RdXErvT39reKA1imj4u1PytenAiyNQuVw4tdPUfOsjFxA1u7PoXTm1SI3b80Jjr
JPBwtB/YH/+HhzPLEkWpoYHaaIClwWjNKOhHLvGUaPyoNQgLY2mW9GQyw63oCkrB
zcUNOWEVMGFUK/W7qYFigoy1Awr9EuZfqcv5l8Tq2DssIhyynbqv91P5Wp6xQzlC
8SuvBImcB9CD0J/m8ryZlHk7uJukd1m4Cz9Pitb6608STFS//ZdZz+u4qj+WA4vY
jFMULb1rE45ZjgkQN8kLZcjsfZ4n4B94JonIP11CawiRyHFLUp6c+ZMRZQm3IdVz
r01UowMkcH2txt8SH0Ss7WMo4MSxIZjZ9TpzfylGhnwmoHxLwiA9zrRhqi5BxRQF
rsvykacJkSrNFGA9zULGVOuk8TzQN15wfe+HpnH3ngygcii1Fm6Eu9tMreghVfRr
U6fqNAYMD40AmEhE+GEbXK9l8DNvzFfVvZ0np4sb3JAW63nVVawnC2z+ap14Go+N
wCBxcv2rusW1sEARLTo2+GMwZtV5reP2JBdMWL8oDLBpOE+2DXfbS8sE1j7k3gqQ
CQWKWnwZrXQXmamGtPGcOqXhH5V+1m2zmpgH7jjACcIhZ4ROOvqVuOt+ocGSxxvn
DJBsgiVSNRxIJ6LV/5T03e1mEWhLcRYBFa5gW7GF1IZb9+F+wU22zHmvNrCg4pqq
eXzOzSKNoR1AabXjeJpyVdC9H71IvO7LP6v9lM1DxqsH4shTdAVO6hWm7TxGM2Gf
znKgmr1wcHOuLQMlAyGom9cGEmRMbsjechbIzw5bQPkA4FVE2jxlse3OomVJzzk0
gVuAABm+/GnsFjgBcEYhcG45DvPcyTDpN75xJL7L+QFMwfzUDp3sWK7tfNsDNPtC
NV92qF1+Xz18jG/2HmxiliQpB36qliS1zEG2wDACu+hOU2I3X1gPF22UILvvOjpi
nZwGByA6+XN3AjPtaGMrfPcosbQe46WiSxi33v+gktpiFhDpi0hHuaeUQSxDF7oo
z4QhqvBzz+CggdtVxLyqPvSKmQyJ2hHwT647jUSArOISV/uitLZDEUnQg6C3F2wx
LHC5SlCVb5sjzoKCLRKlhgsQEfJCrBU/lg8+TdI2MFGzrRL/fVRFscx8azNxWR+F
k4SRkqNfXtYZHH3fmHBLz1cArTr1LDHHOxNaRpmAdqVAasGD902KYn9zGxkEbOU0
tPQjPg9sVILqd1zaLOkKP3hChNV1TPlbUZCRBwDnShPuC1pVGI0kjVx1bIULodQD
NPDzHkkHVW1wcrbU/0OtPbbhbonhtWDHgg4oaJL8pPqd97RC30OqG8RWQV+p9W+e
sgRw/9lwoV3dKbb4z/7EDGkuush6mdEQJU2rELQuEQjVl5Kfx/OeHSF6dbppUznj
tARbkSMpUBkIVfDq0wyCV3VNuQuxyaydzdwudviQxJfH+rXKILB/uzGH+z4B828H
00tWHzz8PqlMRwPKuongr7/d4acA8Gh3X3Ue15ri3XYmAw/2VSYRGoX/s2C4uc+i
bj8qRHY7DIX22atXrgM97QBaEsW63Mu7ciKZocemW/Ej4xLnAiVMGZ2MfJ1zhsQ3
8O/dynhVkKGrzQ+UzHmjPcIObtDcaRH43mYfphqNed9uLrGemLhVCiX3g3X5AWW3
HntbB6MHDsIl7iPMT5op02ZPI6JQYmTfOpkBIA2a3NgEjns/OPwbgiPwXfBuyOHY
8pD7LwpDAZ4VLk9Yep/+/970XFQpKHdFub9gTPkyHvk+/LIaadTC/34nOLp+S5SW
FmsXFk1CkK+j5oJVUoTMvunUq4Up4KxCFwLfe+kRnWxBQKlzNUFRhFrp1M5aV+jR
cQ/TbBTIS7r98WFqZBx4NQgQ1drGzEx4WaxS6rQyRil1fDBRX5FOtk5osKTEmqqV
K5hUG5LDjuGOMTnjexoNOE3I1v4xpIVOiM9i+t6BNrwXOJUuvFm9IMMd7H+Bd4hK
EELAaKGZEAt1ZREpwQOsRUrBit/zPvaCKyhZaj7bkTjBZyX4ujE90F04Rrp7Vovd
uGA0dispcLjK9K3LLJPVb0/aSLclwOWncH/GmIzRe6zwycgU/AnTrQA+h9ikChsI
tbajJ0Gz1PdA8yNAFzQK71qUNw5no8s5ASBpHK4VOTNQtIWKUW7q9hfj+eOHIxLk
trgUg8SkbXX0c7GyZ530pj/76LSHPCyU+laQHoS6l+Zo/Br/kfKEfe1kVeaKmbDE
sgcVTAVULPuUNxC99OdalqYnidH/wMdk9qmq22D7o18ky0i9bNi4h5j2H8ehjg7k
kDcymtZVVJx8mDbs0SH0QVqPdq+dfci7WuVZEl7G15hoE4vzmA1nCGWVLBHipSTB
3X9KgMQoL4XlTs0fBvk54kN+ZVpXpAm4HruV9m2YYdxP7FPNnTGkGElLA8eEe6GS
SCXzIW+plLz6GR0MrXcHN7KC9AEk3qih6zStyQRzmbAxmJMLnuZwYmJq04o481ao
7rWiEQRZnerRv4S5XdGfDodCBaa1Vf0A7+4Y7J6swUBwNzGy07OP+oA1iGu8/jVv
yiWYbXf8EkWwtkD+Z18+awPbEIpNk/9S4iccMJe6OETXxUtcBYmy5HcIUPWvv1SS
7HblLn6EaN1Wzu9Q0jSnexVEZPjQ4fliisLWnlVV4+i01wHAdgGQxBTpmIVXxzCt
G6TXKjXXG1CU+d5n5wgN4Q7+V7Qmgt2BQHxDpv4Wg8Hgsot862Sh0pyGNeOWSZYy
MPSFGeZ7UVpgWylU8E0GCX18/FApTJX8brCb6pzMBz7tloBpqNNtpb8XNB54kBHk
XC6HGFRdQ2FXu7fm/D5D0s4XaYrl5u1plJYXplh/nfnKnS621nnUedSQ4aE8+qZI
yBUup2L/aQb8JnO0xcQFGRrM6hO/ic0s5taTw/S4XCTRRPCwmjEvtSaLcFDzdXee
XPMgOYTb57xHNyfufpgu92LD9ceAZPSEQSvS4piFUFJmHLhv103jrWEncaBtwW9B
cUTGBRSjtEW4vdzxHGxWiAwfqEyvDCGXOdeX96zzlkm2hAd1nQTFJ7EWHuMu83x1
+HdGxLWaImgtyoxcanEFhrSguYGsp82j6/4fvuDYw521SOg8TPzKJrHUwNRgv5dU
d0HTBPBPb20nXBQULrId/GheHT2alk43NEpuvr31OhLPHsOz9UxxR1/Q/mmHjb3m
jBNLtHYev79V1ujVAThnN/ay41/Ps7J5dcasH4cICyCMsU7nEnsz0OWxlnMZtO8L
ZILInNBObgJdZR/CKPaXI6obV80rQWg/Bcj2H0fqXKdRy1rsIUPbL/3s4byGF2ol
Y0/x8V8kQp+p6468oMNfZdo7VAELSx8z067jfKpnpnykku80u8U9GMt9xsLW4eg4
95L1utWZikDg/1HCpvjcAQdq0jOv0hXb4Ez/9H+5LPxETlH9S/toictazbyWqYi6
+LaosK6NsHkF0BDqONhMdfKSdABNYQW1Roa5PM9Vk4f18GD7I+XPjqpfE9Wih6U+
Xyh7acSxsMqP+kjdryWf+iyrqU67JDEWgyWcTv05bWM2G65GZ97RHAVN+7pawI4c
0bl7NiIc19dkaah1qNQipw25R9CtwLeAkYNzdOjP1Jl+BBdEm7x/jJi7IXVDpLW2
CTlRYuAnZM/HpXr/H5g7daKFLKsENf2pEWEBP0qLfLlraFsPtqVC/GIfhAUiPMw4
Z71la1ZpXBH6RUkxTYYZvY2e1SvtZE+jbbnshlq1rv8PtlcTJ58KZHfFPzECJYYr
lzDkko0plRzC5lbeRi12+gUhhEsC9Wya6FChY5qthY+AY1tixqB4UcHOyfQIAN+d
hKuOi/L6TdVdYyFpl4KoGxMmyy5oRpPRzUpddRrwMdvvJCyfEZFWcu/e61Tsm3qv
SHDBi/ffYP89GZdHeKb6j8CU6qZMQbGQGYVVPvRRB2tGLgxs4rRyWbfnKBP/ook+
1Ki6eKpn8ViSDPr6IIdLkWVS8Fj/jmJY+OIZy2ULkSmx7+kyLa6cxJPpnIGwjMZT
z4xdolWbQEBeqnKadVD+SsQ6eCrJIEgHSIf+KR6VKmJvMfwC//QYq723K3f3XHb3
1zfHolWzII/thE1MLODemUfT/KU9Xa20p/4v7VaYqK1ZfhEW+p742JsbrKFHglMD
BC6d8r6Nx87gt5HhyrbBev9n6mZD3g83o/YMzyUCimH8HfnYyIU0qfiUZ4VBnMSB
IagrWQZikzOgLqethqD4MDfzGuUTDNEHt4enWkAnPxJfhIykj6S1sEHK11Ev+MWT
N8RwNnbP1/tjHt2SwmAJyrdNkri6v1KVxZh0ssykTnom1+cgxqMUlzOLYeXlkh1/
mTPriPq69kBSWvGGFfZAiJsUoKI3gO0dJ2iRzbBcQgs2qd7Jgl4dU1Pg5bbbwqDt
Nqu3Nnx6nsZFF58CvNFj4hv4UVe5BmTN5FNd8ilY6XP7WYnQlBXxjcQK1bdjjrm+
9kWdCl2EneBAAaulcW/z1kIANooVgZZshJb8+01yQ7Y2FGUpokONBIJCg6PaIspT
konwXaKGCF4tKSMkYbnbH/bfsS4+dnMn8lBEBkLU5Pgh3xEo9AlQPwmLckwsohu0
3g+w/ArvIHh2y8tZ8Q+rZOkGmZPEi7206udkuR85gSR6GBg4C011xkfu5DgnCYge
mpZnWn4EoyGKS9kLGtVte37e2pwibhu0NQOFpNZrfpcxjCAv0+Fs8v1YmBG6xJVg
crGe0sPg3JjwaZRmQmbFLiyb2V4vvk2GVwi8ajSqbZhOjrjIuBvyvssvjQWtAFrk
6CM+CAoR5MuQFjB+4H4cWQmxuM6GlAi2TA9E5MKO9SjIWHEpq6WHOC0uEI9Bnoas
/lzetoY3PkKVGNRuvU3RwnLcYMTOWh3KRtRnDZbIRjBbe9IY7N9vk02z46T+0MyB
mW4cStxOxbnAaflPX18+RjyeEVplTFZztqfNN35gC3jpY30kd1usxuzRYd3syOpw
+mIj4dVdzwW3Zj1fBhW60kGm9MwoT3eocJ1+FSuTJkX47MFaYCdmwNH0d1STMtH0
qFJ8v8zOhC+otr09lj9UHWPMRzWhw26oUoR76fHVdUMsJNoENSy3xnS43vu2I4wm
tfHauP8g1YzPtfxkRXEao0IWqI4OqZD97wiHxqsf5gaiuhUTeWitlG+Pjh0SIe3S
3iA3iY0OZVQv/WEbHGxX70FRcFZ/SV3SZU5C+PSR8wstcu/niyqCDp8tcefCBKJ+
c9Yj4x98C9f+Ic0sOREf1VHmKTP+a3BA7U4/LbpO0XxE+k4Ikb4+S97ocZU6qNcx
MCbcy8s4sQgzbOj8lv8BQzs+/jBRyVkFaUV8WbzeMZYRew2/aD7vGzADtiaNKv+f
8h3I6m+wr85JsdC4V/zhOGV/oAqGDcOrLM22TBOo4n8yr/cDQZUqMEJiKuEM3Dej
LIDPow6sQ+m8rTSQkQRnrX6wO/AqMbvsAAjDN7wrpbDEkg0UTWSkaWl97pj++5qD
afXdmj/ENsrB8gCF5D0VFL6j/aS4DrawdlMOrqDX2K1ql3ZNfCEYU0RVsmrm22Iy
8xozQLWqYwXjfLjsimvO3a3jkqYyRAid6NDZWsHeLJMDFheKCAIJUi3S1+T8hSwJ
zYbaJjbhYx70900sVJAMoLjQ58H7a1hGYFcyhSMl6+dWmj2CMMVz2MAPfNikGUGu
ez/fX+Mk7yrFr8CrH4PZIrbgAKj7Kqed+ZjmKGehWZiC6X2JKdePUkxa4Fk3BE1B
lhKAyUln2R0C69cz+m+pWMokBPLgLiFoBQKyDv7VuLK6uRQS1im0sAHeN5g3KCjL
ZjURaInEOwxRm+fg3ABRW5MYinS7cX/WMvl8/oVwne6s9jdGEsxvbLCyivXNxs+B
yu8W5CtE1oRbn81J09a+T5kZMZDN2zOshmX2qh/cg03wJwUUjuB8KaeQCWsDGZYi
eou+5aBtVhNv5xzzFeDysykoYLc220kc9SabaIg2Aqwp9sgwudw67+b2hkycFJAA
Xju/6jSWWGt8/Rkr1va8CUSeC8CYyRZZjexWJOg3MGt3VZNBkKcdfpqMqevdhhAG
9lHjSvhwXn1WJO/+rxHF3Hm+AFhoQ7Zm5GyQSn4MggD7RHfJjXWpnd6gRU2WjDid
gZicNETzWj7W0xNpHVyEOTnd3RbOxsRFb7b4g5Pqs6jl2aYIh7Gdh3li4BQ8Mo1s
yGlKMlnGsOkDaIa76QHtTw9fZD9QT47iFkjE+Ndd5+fwZNJIvWwcIlTaiteaeWI/
ecQa27D73/MxDx/vNCZn22eCclTmbFOipzQDJQlAOQc=
`pragma protect end_protected
