// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:03 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YELHIT4j2Q1IgRCL8GP6OGv+KGWWqh50i8YPm+pLgyJaEM/x+eB7C82UcAgGG3IW
syurnP/oyxVzeFk4xRm1T68HtpxPQLnLJopwlPZalasBxMzTFy/INVUmwKlA8t2J
f8sQS7LnFY/ZSLtBuJ+HxiBMUAwNgxqRd5nPoVYZFes=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 184592)
wr8SwwWMNAJfga6QWF64CstZ6Bg1o4V88SgJfHrRu2X7pzMOqTAm5ybhtWjw6HwW
oKeASkmFi43SDQgGRM4NoxdHNfYaChagqQxrHcmIbREln6cC4v9ELteNY6BiSMw4
jLIJtljhnBf4k8iUTfrGfdoE66a+yordoxckpdBUd1RWue/naxsUjOV3hoKrU/Wb
nMpPH5rfgape42I4+SM8MRs2BF/47bMxY9/WtIxcq0kLzCIkb+s0hXXCi0Ykm7d5
xbwVx5MDKX+TW1qwqhMlmsCIUUfwjv6DZ7iHQm9EYkBGyBYS7ki5t4995IChmpWt
xx+31mMbIZiPMAXOpWA4i+Z5BEUEacCRWPUhP2eqsdjzntZczIqLDcJ+iC+2cODU
Uu6QPDRqjoKpZM5BOdKrX8crTH6Km/Dv7EYt56BIDsSw4Kq2tX8zMRdGJYE/8bYZ
uyOOJjjrZy5ilH8RGnhpJRfVeQ8lEwsXqJATktoJRxUfnNdS3IZ1MONPAKVIMAxN
gnweuD8ict+SUlykuqjGl3BkhJh3PDfqNe5MNQdiozFZ6LvuvAXBUefMpUf4vbR5
QMxI7fMy+QLVGs3FfORw9QmJzukNGduI9iLDoO+JWchsrsMYFEoKxbdOjTZcWUSZ
eQQawshYXlF3ONRsbd36R+Q88ugMbLohTwmVOCm9Dy/znq35ImMNOYX59taFGpl5
HWd1H0MduYGwjRRsuP4F5CeCM48nHDhkWVwd0I/Sj2UutmLIPyOS6KjZJpGFqVCA
HRghc+J/qgWpfoZX1daDk4AYHSTucWBSz8l/Y1y/ETTw80RZilTENE72BA4qO2z1
yBOvV7bwXOGz/+tGawyQm7fTGGjZUmbDoIzx70UD5V5XJxO7PolrCrkQjxC0Cvfs
BbLMUwQW1GKdyMSxJyHQoJ9IaSMqGyW3OX+hBQ+deV9gpPPnQnV+3Dab12MhBXIz
anEAPS3R6TBabfPVr5q32QxVLTdc9YLz+5VR2xloh2nwbe6ULPAtMdWx27kpuiki
O9jd+k9FRYOvSd/viLlsICk6T/BK3zPjxl9eXss3sN75AqhOWkKDkYOmgRqq/kYw
PHvYK4iH9docjzuAeRPnO9A1XvrEHpFKE4a8rt8z5Cm6Sco+CrclNhAZGnw92n6l
6JXC21VuRs/E/L/+jfLi9cqjCLT32+tQxu5l7c0blhhsOSM3zKxpsdLhwW0t/2RD
ClbdvghM/eA/0jkJzo/mz/5WCU1bYGsVNMuwp4USCSXAahMCrXg6kwQnddWK8sGT
bnozJCKHMjVuh5d8nPCf8lIQ6ItDmuCx8a2nnYNELKNpzIVVe24ki+c8+U+0xJDX
6aimWM5g9OH1Lg+hvwBDoC/uaSHQCvOph5rxn9xzTa9abD3iiltAFxs715lgk4cM
Spv/L5PY+CnHLcloVsVl/Y25ifC/vyfBW65JZMZAEbdhGQtVY/MwF0MhiF+iUB+i
BhSoit7/lpYxVswOL5JuVuQaKcJgHFoaJXESxbDza036A5aE8RwG6OETuF/GqYPr
mDlqdtPmfNUYZeheZLoM6ZeWj4O48zRJsleATqK3JOCUm/2BpolpYPh0PeC6OeDw
/qbgvnjVfOn2mWHt0SzxuDKoVc2R9I0fEMAACwwGoY3L0IQHTEZ9hRDs8wTAEfrx
brX2P9Bgmr8lyqT0+ZBc5Wk3Zo+9vgm7yGKgrelDnIksjibo8rniWX81fUDobugF
np+fBigO3nFCx/2pdQd7XJ3p4oL0PU8A4iaAx5tUmJUd8isWTH3WxGyXZGj8ZExv
ZE901wNKp2n0RpDLKVfWnXcVO/r8m7Xi3nwFAOr5M40IWiRGqUIY+J/BOk58VuxB
Qn87GAO0NeWH4JoFzPsDzjzTNtTIRzwMzAqN0ew1jabympGUTRVCcuAkIBSx8XyN
kkxZ36n299NQrdewYsRvccBsFZhKHr2Lo3fJLinBmZesAbL0j1fqAsd2z+s7qyh+
xD4Z+xz6WUCqJ1ofLGydqBqFyNGMjuB72u7sRMXUg7TOQqLR38X0SR4qQEyvUWDt
CSLH0S5qTvL07O5STxfILrKeDpsLjeNntHwC5HksTAnZmNA9cKAjksfRZUG95HQe
9oKZAUSEJ4kvbx9u206i7eXzNhvNEtGSx+EKe9+L6mTTsImWxbHErJpdeGG4uMn/
zamPcPoI7bWgMZcjYfQuVZJrRP8hwy1aEzCOdQjzAszyRNBhwM3pieWXfMuXIL68
sncRKHPzkvIPbfj6JEaxa+Xkj3B+V03/6eaXv3vC0Y1YmUOtH7HNS8VuXPVJZh9/
av67k5rwqZ8ff0xG8Dxd57yfTRkgKt+cvNsBsOIybxusdimxKQR5JF6fc2EBiCe1
JcKQFrXAlY+LmTgp08wyudzdWYgYywJ3sBHgVDAsuyPSJ/NP4/x9xlyLrqib8ffn
OU9OKhJ7+YI0+cDbYLSvrxwRIfx2clA207/ES0gPdqnQfdF65b99tfgkTuLCNFB1
sz9G5A2Q79HzMLZIWl6jlgjdviKo3Qabj9zYEKSRihwXJmDFxeAh6FlBucmOoFDI
k2SJUDcoiEK92Q1BBdcYvimB4v7GC7sdC4yD2z54lITptboz/MByUJ043fmcz7g6
Ve+g8S/QfSRvNAQXnaRGWoFtMzqX94E1PuzHjxb6ALso8rKecW6QnBOK0sXwAvgJ
B68M9deRxb2ydw5L8xR9sGc3LIMvsYznVSihLBP3Jc21CJKRcJdLDynWPb9/TQ4W
UUQUbuTQ+tHDxAIU01QPJEx6WXA0cINr/bPyMN58WeaD+EAzbhJ/OHhoggQbCIc8
Z9TKXJ78dX/JmHYNDwb6CCOmftWHMUW4Fg78S4GEatftmvKNYT/O311zXSPnxYUt
MuZvB9JVLJnJcB2aKC+XxqHIRrbUrumDiLru6lcj0YAaVPdMMfHfQZTiK9Q7QYj+
fXKHgyomySxeQ9KD9+E94N8IrrDTU9U7IOsvn32QP8DwmtCcKxR3gzXTCWR5t1f5
usXbarHRGUHby05cbfaXLmurgSF3oOJdaNivDaEXoxHKoZMUFfN2GecStuxo/s9k
O13eQ/6t9+jKoEotOGsXfu+8jtAtLxwe14jcPY2tnyVujKWHYmp3TXRmExou00Mm
BlodTirt4CNLwmHF80OEtugwBr0TzPTqNAFOGjpzR6eHXP7pKWP3yIhB0/+Waj79
b2gAkjXO3QOU2KrtI3vflh5hJINXhrymAu+TEywcPNhtyDE/RPuGozL77L0ozn95
XhdqZvJok4FEusvQg35di80zwo91BvXJCcBTdhcMYa8nUs7u6ZCT47R146jnjjEW
gO9eyjAZC8oq4gFIKymQHU5y7XS2eud6TDxZ6HvS3qA2eEraImfkZLT95iPCMXJS
v/0XL7r4npLDe8ry5Gpu8mUdoqr+/U9GoCUYPjNXXBg+r4zD9qdFr+XjugL6CZBG
Q3L2VyKZiBPYx/BJUQWb3YPPSrsEtyToKWgDvgtxy5GfY6tlkaeVWENhb/+MA8gW
H/DLRRI5iveR7iplF8+NdwseRXVukumCFggTa87i+meVb+m8xCgpX0dapMI9ZFb3
J5HznST30oEHgf87a73hk8A9VCFvxnMnn8VFy+uXh3qi/2lnA2X8vfvxfX0qTqIq
r2eGg+x2uRJG1hpDgdE2eOqTkPyRXRoNBEJIVfqETVzVux7sJhJrZln9b06K4EDJ
tkxFrG/3690fPUNhD6d7c5kq6OpS8NjFD4aO4p2GzghTw7eIe2FzY6IoL7BOxtc4
tiRxe1l7H9bMbbH7xLslFQdH9M+2E3WlTPKCAIzGAs1kyfDDWk2M6oys+yX9FEsK
IM21M4UBCr57rqB36zjsYTFfZt3v7Zd3a8FVFtDWPIiqJ+4dKkxgGvZHzpbkpNU5
YRdlWiiEJXYEJ0jDEjt9xH7KG8UEIneljtNV/yfDZiMKmAlGzVnuOxmBUudniXDk
Ull2jgPt+fQtkmobd9vhNlMRu2tZPYWE9sOW6xXXSMsgcwEq1JH+FeinTHhkk1/j
6se3+awt4w5L+wyMpHr0yZdlxlRtcBogdxzE/Js2T+Bxbo6JM7T8/jK1KUOXGkGB
pjH+wJo1XWDp0ZGkpZKghmlBXeOM0xMP4ZBfmmICJEqxVjPHjdOU0xKVeNmVwvi4
SJwRwU7/+4iEHuC19NUpPD6xdGsvP0HzSaqoBnLENbtrvnmh0UShX2Tv0DO7IfCR
bYfTsm0I/84iE3PvN5J2OqySxAVjAnEYeUTIhr937v0usLxayS+et38V4jDGbniv
v91qVUV2Fuo6tdC0qzUWn6phkHaURC8KT3YSYJHp1Ec93qoyKYQQRDkfc1Amru1D
uEhjE1jU5++PraILotHs18hnk+kU/qEJlC+MfakJsK/JTjRvMsfXHND0Z4bhAcJ0
4n4epxU866d+H6sAh9+yBGtWndcY61DbHBIGVdg47YhbwOiFc5OUdWmrJ02d7VOT
a6PbaLeoFLwusahtaMKnrSpRdB0M113OplnFku+pwICEfn+EEuA6woAzVO0Xv5OP
ud0ORrvOvBWD9UOTTmERrWNIsc9reYS7zc/AMzHLPBlTavpc5ck7CCopiA4N5Rp4
bgGbzK7b9FI7Xb3J97/elCMiyfY7MBWJFNKoV2EbLuRdiAqfsmnQLgUTIGBlXLaw
vHlncRhyCANfqDOXpgHul9jWv7Fsr+MhNj7hm8Kg7UYEswVAIzZ9nKeRQxH3NS6r
BsnMIknYRYYB/Rn/wS1gfeGt0pLL1LmxbDbBo1Szp+vKcN1pfwGQzIGn8CH56CPl
HUtmmfnOeAIeUmIKdumfji2JGfVb3GwQbSQoBkCPJRQENyhb+L5JzdTVXEBPeqWC
nA9Hsl+OaarBlaQOb/OFXMPqNZSGsAOMIy1ic92u1zj7Samfyi3F2ToJ5hdKllp8
EmzVJuuO1vXEGzggPXoKZe1K3vjvrZGeBTCXXPD+GJ11GI3k5gzJsag8HIzuXLRG
S/o1Ew3PH6mG6gV7RteQ/qcQ1v21w5iveVC+cUWCUOGjVjefaW1oG8izc/EXKywd
GN/LLtkE3iyY61QYmX7tb9/1GD2IHQ9Br5qbNMUjCGetoFKrbQeUOF9fWzbslfYU
lIgyFCmE4ykbpt8OyhJj8nPf0OawEmBUR0ftmX1QXA/LmKrQDpTr/3QDs+ooEw6A
Eq2dT3GDr1wEmak8OPUq2j0f5JYeS5nk1Q8C+voY8aa71Iukvr7HByiz0n7KFBh/
vYbqI43gIkjgOIxLC1c5yRuBSe90z5ZA/GLiNo7xntMIOZLZAWFPJhrHph6JMkQp
/j+erOUeCfQjXRRm/BmqL3KICV1EnXhIjZ8YYgUoqUJKS8DeQ4DVDSRJJWbiNzDc
EYUgY2rWkdxl11x3YzikDUudy3WE3/7J8L0gZKLwFS4CzCf9TaUM+lcy2kXDYZLh
P11LBHaQBV8xvUPG2dYDUd42SrGx1PNMOimz2ud+pEPJx3wLMqFcHvTL7lph5f1x
Jxx6bTFEUSNi76XAPA0kWipxRyNgs0+UZKSN2q6L6vQKM3eussDELMjOnNdevV2f
21s7Y8QSWOuYSv1cYQA+oIuJjdnMXqh/moDgf3f54dyvrkz4nhFcl7CziIOSkKi2
EnXiW15MNBc0OFvJ080URRlYXnXMaf3mSUA+5N+7QmKFop7DkXuMf52WXFYzSHSh
csznD8fABd0wEwjcm2zCXcYl9qnz5gn4ykf+WZw0I0+AKkG8xokx5dqkMv77oq31
Nk1HA0nYXUIWSOwLqVlwYtRY9kAjmwS4H/uP3XiwWUk1rXlL2KDV7w+/qMdzhaeu
FV92FdH7gvzt1G71ZJtzrM/wEauCzgXlZsz9JBjSBSAwzyq7NvZ0lst31JVFudwF
ClVLD3pYpZtbf6GTqaIZVrcucL9JRNKKmTNinIFp+hmCfiYconbPVtVemdwaZbZP
3YdImNZnlRBqADCzYEbRedb12IT2mp9OwG2kBq3O6NBuap4QRa4ibITRVYFZWNML
rNqH1g9eieSSpxMmOrWp55gZE4Ewz50IhezQavBGAH4ER+VYtNBS4NjbP2InAsdg
ttSzhsJIErQ/4ITWBMJhqJyMgDZ6+pIs3idTue9oYyuc+3TKCRpEH7Y8IR8hVetY
hITXPDsCmJlcEJ16aATU9Bl0o3m8PToHhGRYmZA9PqSXGC0buZsjqeKTtlr9Fm5w
KRqrnf8SfugV3FT12betedY6UJUxeN9Aeh9yg/HP5lMpKTPEtvI9CTCVlUd8haZq
1MofsE3m+9xVisxMj+UFcJx0KkGFq7+E0LdpFyTUPsDFV6wZHxvwMmd6V9TFtvvo
pEZ2NpVs0FpW6kZAGkQCoVGcmhpikNoyrTdZTW3KNiLx8L8ffSt0QMnOGdj3/YHv
zQzPUEZ+9r2gemcCSRCAqKVMgAro13USbm3910Jz6XsUKlH4Z1/RvH0Oye3FEU4w
XZINAwTMZrsz9CLYF5PZOkPWqYiWEj4AQiStL3YOI6MdP3CmXyEHyL80OgtI5VRp
ewRhYKgLHBMzDD+l4ZMVsa1KS+MhNQg0YfolJfSMz2q0r7ulJe4VffzIWkanIyFq
6hCeOymYHh9e0vD6g/cTACRnfTyoSuucRvOPkSEEzkGEOEjMsWs3ubppnthdxyiC
VBpHJJWqIPaXTqXBvJVDUARxBvGq/PO1cXssrOgAqNuD/ZjUYBkbKPs77WNYhH6R
AD/QvJegokdGxEmXy4i+3VSPFupzwypraqyAlvQH8W42Gc1BU05qaDav3BFpnfIz
NXV0j6/3+89IpmXafNyF8K/JMKH36nYyx4K9E6/p2AJCsCZJ4EHrf3+n/FKKdZQE
4QvS5n/ifW35zHXYHFJpOJYu8yVNLEBuoLBf7neeSZuB5qN0d6iIY+CYDXbZkt4u
dqZwwGDzmhgflykuATlkrjbL9hveeQo9NKq4qwK6NaZUh5gggABoZedekV6Qf8HS
I7ml85KA/0g/7ziO2lwkRmRfKJrNu8lZH7yTzEYRlp2ZpcdlVzeF0x/J9dKBAT/3
6NJD8dp1fbvhLWhJ5RWPz6mGGxBxZ+qesK/+rWOUO/mldfDTCaGNziF0V6PJPSko
Aa9kmTO1W/2CXs3eXHMt20Kpu/qox64OwVMQhiAoBgjbBxfzxY3iQ8o2Jd7xjH6V
9hByUHQWMJFCKG8J7pYWN1CybcWyvW2l8HymTKErnSFoUKbAMXxNw9OxJc/tegSj
5PCr2L6ZXKkRO04ZZeDsByGTWNGMa3zwVkHKIBCpuLIdJe5s3UluqGTnLM96h69k
QlENngLt5Z2y7FSnB0p1FPldYY+sacTIkGJufs49EJrAAfd7cO3vI7u8UwQ3gwpD
6QeP8tyUx79IhuFKokRJDKpN91eF4fzgm7IUAS0zghJnrOXZ0jHTl0XlCagdbVUa
ct7uovrz5NaHfjMS1EhrUDHkUYEu6WYfkz5CjHgwKSBy6INt2NwSTTcFUSGA5T9d
x09/6N/B3XDSOy/dm6WgzWRUEK3Q0oCbi1yf5W/m+ChB/opj7ri3Uw28eXl2yI1h
fCHpYcTGgxIo/S3BKJcMow1HtpRH7AkL/2tg15Np/NhHGW4vTCuzz3Zvm1AipiJn
+gxSu9bUapLaB4sbLxhEDAFDChIYyjWF2rInzHyYH0FVi55D0k1G4yF43dFvIW60
6mF0ul24UfYJf+oS9gKhxoMaVBqV+V8ThcdEz+LUTkspTFim6N5LYuJCXHfecZ2d
lXM29BI5usAZC5SuUN1aAkOTruvTfUd1BQQLCQINFzNAFyxleHPUAGBFa+/GHOOS
7b4I0cknLWkfDQfnZSaPk6DrNrPZr21WwIMmFpj2VW2BjsyXGhbx2lKVLhJY4IIX
aCOqMAoeTYkcf1GKfUdBpfboKu7FFyuTOnFH5CdU8fRwwzli8LkKnDHadxpy65wA
Qe8d4H3gvjvqCBxr5VXP56ZhS/4iCjBFy5Tlw/LN8JuvBTP+j22/VjNufFp2JqGC
HIaDhdZvUUVD2y4UwYLGObXyOAFCIUZ91J36LOWouYKf7AUty12zS61gBujnSzOL
2GP4fk/EChA0WkfTwadt/Io3L76iib6SmGfCHiVNSyUBDHcoZRgvFg2WoDZE9dO+
6wOJSGsfTYqXs1kWXbNaF36keN4mtb7aUtdoSiOf2hIOCoikmyu2bz999YI4xVBJ
flwYlqG84rA43GjJX4nRGI7fcu/x9OR65H/pTxr3oszH1ycAYqeg4ECtlKDsUTQE
iy/vH3ZgzknSWV5VUuuz0W8qFjTP0InWiwVTb0zzF2rMWAs9JK9VEE5WSHWtKJCB
AeH0YiVa/6Ql7l50k/OKfQQZPCFogQ61d/Vj2fVT/xLUqDop4rxpRBJNTqPGkQYs
aUBu5759PQ5mfFvuAzpqjyx6W1wZXNQicZzOFeQm5/0E3/2wPC8rKJX97FxFnOTz
uUfm2ivfQwkvQYqIvPpfYMvcnOFuLtEQFFoNszwloUg/vGphByECANqB2rhXGQoA
BSI6fMcu6qoyHIqUH/aJLo8oeLdG6+1Q+i4luZLjHnUGgmyptfgIXlD0eVmZAd3B
TD6RejDECw8nUmCdYj0TCsCpRcyVsXAJaRD5nvCv8hz+GOkm8t+lkZ0ZcRnIX/Pk
SzRE9i/Rf1UfyCK7cCBrU2DGhJV0VCW8lfNxIztHN46xaIVwUAQgfxZ2O9as0yD3
DdPpL85gsEzROJj9dvC6IZbw1TJdaSPR7DQj8in2HW8w4RsdMvePJZbKDEoRoQhj
2KBz8Yw3ljtscV8udwXErdq7g4HX8Raw/KMmVWAaEmi6hMuM6NOX+72ACd9/sQX/
BrR/yABRn6Olur9Dl7mDldi4akFiIepkpALhgfrVTTeNfV7i2sYUWUx3TV7KgLVJ
CIJWUBX5p7zYVRc171LzBJgHxcWR4tbWTsLaTRko7Tobh9wG6JcIDp/ptTG+0u3z
G8W2rB2ZluShS3+LZBAvOz7VUqwwUMoaK2khed2TJuOc3ShOWn4tyy3gN9DEi4dN
LBMW4QpsG6zqxxMdUyd/WOy9Sfq1u9KnS2UvF+jE8rn4M7Z8tvVN9ueDh+Tth+6f
hiCO+7K5/MB6UqUNiXHOMrG/M3fJInOBEkKa5PSu+Aplm6DyzO/LEJfeEniixX6D
CxOQdCaVZxi0mqz0KGC8je+MPAnHTWDLRyYNBx0Dl+wAAk+Me1z7GFQR56EGLEbe
tYDB6FkqXG8g83v90Cq5q7T7pKQ1tdNKQe53ahMJeGtaBi3uVibhieT51Czt4ZsY
7pyT83/Jfqq9aRQ4xVlVqfBwemEvJZGM92Ftv7wp2GP7zvk3Shl0b5XfxdFCfh11
9VM//E3NWpHsMTVJKJ7BBe8FuAfpZ5Ek2i/+SrzGMPhN57YiFnp9N8MifxuKW2T0
NI+k22hFPNW0HsEyl/31XDLIJEdhZ8lZu/FvZxMQKSqsi5h83mZfFGSM8yqxYxLR
xUfQNw+ZJVwocYYvuzgs8bmSWJqyfABJBKKDSUgYnLJqovgXE8e+YpSCU/5aCy/T
CNZQEAQGPqeGpvW0WFluRCBB7e4GCASDO8pd4gRlXm9KO6S+hRTSDiIBaEDUQUuH
Tkv5woEJu2ztL20asmk7oFzYTWexKa2sfGtEWsjSbPViose25TtCgpPhDqJsXEKl
7NHNV9+nZySQSLhJV3tIad/SEcpQ3x3yDXfw6Yimuf8DKVQUZ+XsA5O57G1hGTOX
ajH0fxcJUEowClM4aC8Yhl4Q1MTfaWsf6EDxwnYB7QuVViiWqOtgBgiXl0auAbSD
Hxqwm1l7jv4lHJ+ZR42gEW9NQ9lBbl/aKFcqmzqSrBip3sspDTjxdcSMu+PgDT7j
WIQeLLFRsFJMQkI2htskjGf2c1S8BCzMgJDMMhztDtXN8pt3xTWGqKpGzXoTyKof
pLTOsXB1YEQm2vFCA2RfMvYIn2bdeNFayFSqWg+AEVhIjey6K5vSD3L6K1pfAjfe
T1j8vvh0dmh0dhzi7tDVOXU+64mbxCeFGkOuB89YGsREgimhotV99LSPDIS1cqft
82S88W3md6IPEJ4wqrwCm2+abQgzjJAQbve837ggfM8kkqIz5apG2vWQtlpU+8A+
aIL54qU6DgCdLbOSmkKFZQfAcVozBGxBVCGbWDjb7de6+QWWQtdtjozqF7AH2MAI
OiCp0bXoAVpNLVclu3jRHT5/y6YjscXOJ9DLYWEfKYLQ6NHAYj+ZPD8wrSq9Mg/k
nFqI3aDo8/doUF8WxB7AUPfMRZvscSFbjSlc7pXArf6O3EmRhzz9KQkdKAE9eMMz
jm1fSWhpO/Jwbvl4ewWn5vTVrp8UG3SCcXKJcgmXdbbHtqG6ZLN6RgtmxqtS2FE+
PZ+EpejjsGwYWdrW3bQnqqdFsW1/k4jL5H+uAFK3YUgQdA9XOTII5nKXPaKLVk28
Zfnuz9yU6cjMcPt+039JQ02ylz4uInXW4yXDuWJVDmOXQ2tNvcENLOGE0ggJGVZ0
zW4rs/CfUVqEYOGgvCcJjzTECij6GIqyAXtWA3bCWSSbkWRvG4eh6f4OOJ1XGBZ0
2oP6iwKNO2u65bcjkaLr/BfhDuzdbgohrexHweUatiT0n1OzYEVOGrlF46CW0a+f
QwFnsZSDE/aS7/GljLuA6LjApicMQZu/TjGk5Lx95tK70/qL6upddsfVYENBRc8d
ar1vnBix/3pOePpci5GNW8F9ttESn6cFdRFcs2EIZYdFUv2I1PaXrQ1C4x8wS+7L
g7SGArcMLG40yzV6vRVCt0HEBwKntzn4/Za3dNPRR+YMotOa7OAhK/V5e4j/czNx
9q1/R4Ph9/x+xy9kje8NeDLl+s+lqxP9IIhqD9UIJOWeAJG+KFxrvPys+MCqj8mq
u6oK450CZDDXn4hWM3fylQfKMQGwB7nkaaHzQ0nJ/PG/LphhrrZ8BQvnV53ja1uV
rGRrz3Qn2UzMeQkDyLojkkWQYZ4+WJYm2NN6kh4s9YX6V0pwNswNOEOVrfEjTMKW
+i671dweSeCSunV/A6J0IsLUEqu8QXsUXx9qUvfZijLLQdxXnIHaiXPIkidkY//b
uD8+JUtIQPksYAW3lfdIVCSac/UurMarEkxruXNYJ+WlNPW7bu4Wk/zQU9WcrKLb
Mf0ua//h9fASQhoI97tLUvTUU8rHBfAZ7+3smgI1THYxnKAaLy47FZ8anyw7UqxG
inG7E37E+u4p5O16zZR+cEms8ViBgRDGUK5/5909pY9rgPWgdBBGZa8/Wx2EYZTn
iGNV3Ih6et+NwM4zjzgaRbAVdfaOHw4wFcH/Z61nffg37fXRFV1eHwo3226QH8Po
ki6qfYEQxO/GuqIfASO9hADxm+Yss3GUt2Gdao2NWJzFfFwsQZRDjGrTiH4U/Z6S
jB9Ra7+TwzzrecFcn7m0iR2DI7gp7rUqhoRz+Umu/FtD1T2tMVviW0KZG4FASwyJ
lx4rw5Gs5oN0sFwumP8UP93isvurJQvK/w//tnGFpXTv/8IMWWy7XXyJcLGV+Ff0
ipegqka3AwTwAgxS0fjhb0Fele1ZDj2bfRwRvGk79FQskm3903LGU46BDJrdilA1
+rqRdWf+MN7lI/dRR9ie1G0rFpqfvFdaSTpkWdpQjQE4DuCySLwefReBR/VYUYgu
d7WgJeoPWbGmE4E54hAMLPG5hjhxfBABZFaKFvLD32pMbZr5TNs8I/V75rCQZUWf
sJL/4y+a/ukh2bydfWypyqQZpuQGMCpt+blglqfBnJHPi43T9TTgrXVU3GntoO84
BxIxf5YBJokJ2T9nYGWbIC/Ou9Ncp1p4X6kYfmGTjFDNq2iNIx0Pvpjc2EmURHky
72r3wjpiiLr7Lhgpwv9pCt3Z50TwX42fjc1A/qto69fEm/F7crzvZHJNt7a9AxNQ
MbDrYYgQiFXLbOZI1ERQat2/qITtlkv5anozoWyDmdQRBUNCxIwITaxfbmeOhEkk
KHrL1/j7ufJm9iszjsWA4XB7xOI8zqQid/ShEa4Pto+72/c8zmJL7j94150xc50t
JbmwQQjRSdfB2S11XAAsajRNW4CpC3QjdH6Xv8kh6O55q4q252Iwhx+bQJgDW59p
9DbRpURQ81sUwkiBE9MH6OTVzzD3ym3vdWr33PTvkudVPyVETkZWjljljWBC6Uuv
zMaqSINoj8TyPoHP5pqKhyGE4LLfAoAiSuELcqgI9yD99MaH/KCYsXT6UJ1HUeI2
3VEwx7qPrbHxaSWeBk57Rd3K6u1OziHbI/q6Ci31Ri3mjAfhmfWuK79sVnLDPGIk
UuZ37WSufwSv0L+rtx0Pf8xj6AlfER8OHU7Q4csac9UJr/T4rt4TZ3SzN2UoTnfE
aPwLoKqzKu1qAZL0OeFDFVqwDAy27YXneu8IYc2RurePJWts26CqWCOegCZzSQSL
/tazrsbe2/CL6CjGT9FMgCkd3z6J8nx5Tx9e4xSLQ99nP+pqRGHEdaDK8i1QOts0
fv5/I+fHQ7/YurYvZu1T+Lhs1BrddxHM85MCN+7NSX5rFciRKclv+ej8soou9dTW
fUnF5V0X4ac421E0owncvqW1guJFigUZRZwuvPIoCWBKXPl2aApLxv5Dn1c7tEeN
57tvq+9owhFAyE1pwmXYUc5hxWMQhZzRODBmZF2Pkq10gAY9bUrILG7gStTDWWMW
Nqq3HJC/65wZcdkdMYAAsDcQ0OFTxXC1fOK8r6twA0Bm6Rgowj2ihQxjfDGr7pZE
IALYBeW1TF5ocr/X6juFrSXHK2SSvmMycUgyq21/BxmhizxELxeqwckmPIzFiLXc
02Pv8uTxskUy0qlWVuXjIVHKMeTv2pjkYVOswNNMUGVbtwzd+PHF5VV1t3wg26Xj
Hk4zAK1HGIpQ4rKC7g8AB/6u966zAB3nWgxQPK6YSAkBmH+SJe79WebEAQRhLcLa
tVoSoOZ7aRlfFYUmx0Xq+F6K584kvmP9uabVqKkqo84/9unahh2tvgop6xIuXL44
4yzgFtmCxqRuc/3mkvgjDgHA+LvtUB/ikxl4mKxicnW27Rka8IGYWWW6SnvWn6po
y6LceL1DMmplOBvFM4UFEjYdHVmkoo+JJek4HXKqyIoNbndWJ3wPl4mmRgwG/QEO
pATutlllHoYBRlS/2HRLbpX5USDW702jquSX9tPGaI3rrSsjBcw1XcjhvfYy1G4Z
kLdjJfx2Imt6JCFk9l0h+C7ZQmffTuQzNSO01PFi6JnlKpdqi6+4i8lubnx9/JDM
jprYG+cPax4VOxZYpCr7ICk6gymKGuxyISSRoXE1iYT3tweCxhiCtKawF27rAdsV
f9BuF+T1OQopCeZ+tBridUELu34Gt+U1HqSsDxncopDVRhIHzmKRFBPcfMWEDR5U
J3Q+x5TR/WA9yQfj6uADH68UiQCfU6YYjAQPcLPvytwu41+XVYI9zn1rJFa3AKEL
v9J2iUIehtDyTw4HW45pkyHwBLL81dEnVtMpadpZLt4Wd3o2NkfzXdISvZP06I85
NVRqtR+Xt6HAvXZBPusmK6keTW0BgCg9mN7eWu3M9LHUeLwSTCqPXrRt2UrxoGN5
ka+BPGdtqLaYa+eSBOCEEPRin45PpEOSNXQ1LAvdDbk4ybL8Or9z61aKepeUVc0Y
doYMPbmoG5Jquvvl8YUByUYEJTMkcsqbOzV4NilZsxWACxJd57eSKV8a1zabuU3f
HLgrv8yq7ixEeBYjS8bIL2HQVd1yGmJix1wlyEazlWfjJjBvF+PbFbzTsQlZqHwe
qzv+wN+2Xc4Fo2M+t0mnUZp9XaoxPe9Ns2hHNLShv95icwI/6h3Ml2PXFtW2tRsV
Aj78ywmy+PpD0/l5n85RKpmYDrQLM4GSToN1qA2QyuD/G6pDnC6HNtzQr3ptgTm8
NORE6/KRdGrv+ocNYKAZW6w61yVXyn2AE/aNGwsm5W5SVvJYvPiOoZiIEwxaLvEh
I3SFJCDNKzhHtiYnzxexJ+nxGAn4IhvJXdOfLpmCwlrdN37wF+DWruOtREujIWAU
onCnwtSGCnNRSxbcX7dTfnsyZ+wIsFZLhsy86f3WNRieZQho92TLPDCJw4A/KVs3
kL+HNshfIbt84yYLZnBUIIPP5wb0t0ieZTLPwlb/utZwDB8FtelqTze8RXDSfSZj
ELW8D8NMw7K8KE5t3Jo99zPsNJ+FQyL2bpR9t+PfJ9t7Pz1USfFrhg+oFtJj3o3X
WBqxi+cm01x/XQuoQLBLGzxQKO/UuUBlhnCHzRJCcs/l46wZfk/kAF9foobZsMpI
FWDQY3y51B8muh1YlEJpEuK7ll0b796C95hq+uegdYMU3OcKz3impS2mgEfY4+L/
tGiGxbt/JXs9eyugrVR3EgY0VIJ3YEUWXVFvk7fv7zl9Q4Wiysko1SNJ8Uwmr1Zc
CcfWBEdEsapEO5yiEafBlmYFlunxK9i75zaeoDWbrj4SeWg4Zgh79QEbKOAQe6vN
jwdNFgGvpCYuBLVTh54lCwN7RvFJpc1tPu446O+ffps4P8F0Ibzdmf35DN7rgPGm
rJ7KHKk618pCz5H/WYw2Xzdema/TTJ81NpjZERAfN4dIU8K2gss20kZbwAt+CZ4r
hJ92Zgy3Q9VLb+Gxlaq9y+bEVsS1+G7py9aFkjCfCtl2BTSJbkeBHWA5VqFbx2TJ
GFHgyA4t/Wmwdke20TLtImNZZ2vRKpQZP+6ubNqep/Gfgq9Z9HjyVqm3oA8k9FvZ
n7Jk3CIpNPMydiTveBXI9Wv4HcQTPU8mlnI1bMtgV5so41cfha5gzraOcEhlnwqt
YJKUrsgA2KvRvaA1avpJOwhBV0yiXLz2/n0nZaLq+8HUBvV8CL8TDBdGB8ZbLX18
6PRDDMpIj5OubVbYpvhNxW/CI2MdXSo1FEb9b09OYhOul+LgW62owfpN8+3gOqXo
WtzwO8ZtDKop43LgLV5tEGRK0xTwQBkLXg4YXKOOSvj3b7UlT7sAGOBohQNajsGq
uQjCDU4fZ6n86lHNpPhcmNVssSama+i66wfSbnQMYSKRLswejinl3NFsj4QsE/6p
Len6mBBqceUw+ysqPNmOrRFOibemaCbSQ4hYT7BYQ3IJRXho42A74idHOnP4d2Fm
Gd6KTGck+NNS/5g73HPlTdMDs4cwRjbt4rQLJZzZO7pUn2LyWQ11KguEN4YxL4Dn
iKa0B6FwSADzYPuo3IP15y+3QtSTigzKNspqW3FKDCXyVzeogknZ5y9vs3bFIYmq
E1mcT2idIRumBc96uIUXCtiv4PcEqgu4mTpjNhbAvMan96wcvyj/90K8WtEV/5Te
uZfLmKhJ3LB8YOhuJUKwMcyz9iFVt1TRTDfP3V3QSjAPUWQXd92H1vzRMR9J+Utu
hQxjU2xorMqC4ZJEq7FituYJ4zyUdYkzgJfRm8ZECtONOYzrPGwzm9Y0pcugWYap
o6882bjjUqWd7M2FlkhNbqPX56yEEzGTnFcWxtPZ5pu66YYK5wTG9FLOU5qS1Xn6
faWj8bjtdyqbnhwPcn7X7WdcZl5n9nmIvCDcsHDIKn7PSmWA0l8WF2Bb5Jg9+0uv
OFribQizqVhEmBupsIVxpT2p4Jh4eBraFVOjGORx0HLZAKUqI55dzCay78MT1dOe
By1+CrpNKaLd6ebpGicqCPLS8hH745C+DnnzcGJ9e5LI/6lSItdKUjTW9VGA4U6j
+goag3J2CEzIZtp8K5c07KyelzbUqbFhSfWLC81bML9EjoKdCQ/rOZde0vCEho+O
aDoKA0ljhl6Pg6hYJOi4KhRwKH9GeTeK0D+3CTVnA6eozxrWs0rbNhgXapvhlumB
FjSGdBtrucmOLnvxZnShMvw4xMYWXWhYb3WT3OATGaZzNZ1enz0/3mpktokOgIRu
WN9sZBU8yI0XHUoQpZyWz0KSTOr7+/FG7ryDdVsDupkw3dfvuQq3ZlneWgiwbOvX
ggjr+DNdA6r4PMQl3kqTKOT38VoeIC4kHPpDInWJN3DBjaL3yoPYq4Gnm9UxoRz1
mX/SEcYwNJ5jbt/CyRXAVery9ZRGgkuAuiubskZci3W49jTy3GxK/XElwzuPlIbZ
HwXb0wdWU1aQM+D0jQKhDYMSfF9NqYuVwnz+QsH7KX63kinTAOh6QMiGSJLZEa5s
rE8Q2mRNECMyjuU6rxRTTMHDLfJ5e4J/xmOnKL6cd+q0ZMJepcdu3sCD6Dkx4nvN
VUBcOb7pwRRfU4ewnl+XH4FOwJ5mm1DItmUl58re2j4NLAmaUESsJYt57rbqQ4Tz
kvqtb4Jso4ai1psc1v9Uz594TIF93AcT0UODewZjsTkh+OTYY9nL2qrK3rsMMtNq
AOvaTWJRR/Oy65tGukcKRfKGOpwX7osagTak2x+f3RfmkpLoZTGsK6tipRcgTlfS
r0E1hVoPrkbhr6zNRVkPHTurf9aj5+5ROQtPjKKSMIX4b/cpZJ9qVts2SMWDYjax
nIvr5pf4TmUzU56C8LbsywsQ1rYybNnpN+fRFslgvSyy01qPGmjByw6mUEklCu1B
jNU7+YW+wbRlOk6om4FDqjbUWmimlkZ60rJr1gzEXZTeKMnNnPPEOsMFVJxIP9JG
RTvAyar7kCRZNXoWr9+g+eDN3jHeeNLmdIfV4zjYbmBxNnSWRPGvbl7oZ7Rb5vOI
VQt66virq0m/BGAqE2W7jmyfBlwQY/0IfreEWlQjWW+cpeDQ8FzURClqMJnov4KK
TBpmDrVxkd0dQBiM3xjbtu3fvsdhkS5f5tfRUD4A+FMmXqYKjLQNN8ig2QaQNW8K
be7lvg4juw8rQdj2fS7NeoDtvDQ9cipk0FueB/sVoyI43P3YYNLdzKV8oxdvn7dE
spEtewwYWCGq+QU6k70X/X7cK0zi9Mm+15KLnPwQ8HATuwRDJfTbqW0NRQxqrUfY
iivd/opULgn8Adcin8FQ+3MgfGbhovV9oTqoWSV5OlWxtNlpmeAP+FjklaAt55Ao
fUMiWFuPK9H/naLsF9avgQXg9wPyOoP5JyUTgcl8JXD0LEso2BstEKAJp7ikJbeQ
BKwoGgdK8cwIMyzaRuk2eyeoz9Z0JnNp6yVCkLG5CTKohtkSvgudDcshdwnbDwdu
XonOBvJsPjF/kMlQWjIzN8FRRZePXV2VqP1vjKFmD+0NtnCzfSBgs1XhneoCs1Dv
XvnX3SmTBhwXdNzLaY3WGM7GM/aeykPz9Zo1N0w7ZjIj/4917C+yM7GQKxFONjJ1
YD3pb0W9Z7J26JM1Lwcd5ld9Qg6zf/rIzCQnLF46RfupbAXlN08PwJZ1nT0FILtm
E3+l8V7A7i5EynmK8gY6ZkrmCPxHl6ivLvlhPW+YTzkJ9Sv0NX/7GN7h+K8Oh4a8
e4taZpiNXoht63pphmO5iG9rZq2SQHO2c+76HSohUNOr9FTXAkSWxaOwpA7RNBfn
uQ/CTCJTzCxyGEEJzA2WsP4OsmiFt1MYV3jygAq6n0NitDTWatuhgw6259TEjLX8
63fasP4HGWwhOoOUiD6C/aETVyYAuxms31TiOPI3WxlPAc3Cx2pwaG0iltwcvtWs
ZVX5hF6RDLwQtESXccK0nNRfjezUPdymbJLLL0V6HdWsWX9ZU3XyuQBq8/bYccTm
ubcrAJ2EJA8mbvyLuk9kjRT3avsdXIbwVUAq73tZ+IAp4aQvG+ZiEINffjd2y3xJ
GJWm8BUtkNU6NDaeraJQDI34sKShW7FY96YMhno7mfUceBWeyqUTpYwhZPCLD0vB
QOdytVdb0RhM8rva+0jrhtht1iZrqd09MFDRcnvNrwYvBoSKGJsKHCOJqUUgY2ld
OxwaRNNPz13DKWRkx7vAlATFlO64UfZhFIywwLbN8mcDAMdghwjncrWXsgMFZxrd
sjnDM7WJK7QRz0faPr+mw2f5Veoy/7Bp1LztFl1RCxM6DppyLxN2EtI8NZ7wG5Ri
CAwf+1U2CI+e3ux4ehyfGGxeuXOZky450ORBUzeflr6XtH8a9avtxNZPLrC3f6ev
bCkKVWoppxoh/o6lYk71qoRecm0M1mGtfvN2irWbNPQVcvTxLdRLRkWEhUnVtWHE
q1DNncMihu4rnx7mS/lNxYTovCdmLEgU2GlvHK7V8VhJVMA/iS+oNT75ffxlwxlG
U0erzkUpMOh5EvfrELBrSmiJN23HPLyDms/xe5O7N78xz1PeSzvwVsKrTmS5QZZ6
9nB7II5wNUybZ4d70tgJhx0fd79xSw5DDGh2RBq45nNIFiwnly8wYQgGxHZiDybZ
nGyocpsa9g63zCNwn0EdDeurgU85Ef3QDhPbGiGSQp6OWKUzkrdkRWWQHuOmY+wU
QVh+j5ijj+Wfo3ARD1ARECAwcrSNriQmd+KoVfaPS1y9uo3Tvf4dHR1wYq17BdNW
kQ7TJsh8r1EJ0JZaDdVTzcAWaLBlSXlDsezHcsEf0maJkDc92w4/OLsLDvq3Lgzh
DPB5bdUnQ3p4JO4KZfoQhwuqQu30XgYzbvahzSizQSMLSyCxFwxFfxDAvdl/V7l4
K7Dx3hgv8a92oNQIumCBp8mYK+cR5DUnlYMpu+FLt1Tdz/Gy7M2QEgtV5MLHijtr
oYUJVmcJsk67FiYMPbFDa+g3T1uRzIN+OElCG/2VxQkA2XsXXf1F3IkOMcEIJi/q
XYcu/xTNFqAIsQb6laBFh/2mplmFjV2oxzQaITw8oOGiSJ9gi8o+AcVNpCCUaZp5
baGcqWeJ1v/rxOv8V1m7ionYhuJs7tXoQfz4OImK0SQ50WXNXYsycqPTrxWuiMoP
3VMrI6O9+t7M/kQTKqjFlHn+IcBRELLR2dFzsUWAanisDYns1s8SlGAWA1aMCrru
NMGb07upulcvwvHjU/ZCjG6iv2cWV14jG/6twfMlcVb5Zyr8paXl2RfU+6RwRSaA
Hcu0cRQtPkvvcWrwMm8sCXSMlV3LxAznOjioBtpisbFVdMHOOAFDXWGF9RgRVFhq
Paw/BVibPy08oetuda9lwIL/CKansTryGVkzKY6274UHl7RaJv3WXDNeizhAIhnZ
JseWHFNxQ1Sjad0A6fZls4+sQsw836qntyMKYl9uboK5u1ez7+7X+qkOnPqsrPeF
avNpEmbGIENy/EuCNww+rl6+v/sS6hHPfOhjqc5sQFJnoTkXtF+yrGpd9aTJvT0r
fqNhztcST8VSudP4trIawtUCzx88/u9i9oiwRw8/hTfjJvSkUFr+lsU2Qr6KcH0s
1TC+fMEfjmonZ1Tf9jLrA+fdYKcQdvF0WDZB9WKHxYg3xXOKKH4mFQEHd0dNYC36
ti8+t8l5ejYhnLJGZPpmkwGOlxGV5CPUDIuHPSiN/UJBqmVTGLtQIp0Ovii9MLqq
ZrSS5oWeoHrwRxVv/c1K3DznvEk2dO5HepLYkFtWi1zk2oE53nQ1bZ2+3kmWuvYg
Q1WDNoxU/EXx/yrlM5FJC/zwRZfXw4M8vN6PLPZiU6/plNk20lZ01eGzNMQfbE8p
Yt8lsaI/cWAv9n0w2IX0jDz7Yluf3lWySevE0SJPRLWcaKZOSsxtQkcvlDxd6MS8
oURgNSgQFhC3NxDGkLT7Ja37Rhjf3RyoHHmTYR1RwFrnBwmB+06VYgiMsT6bJ4pW
cWBh5/Gaq1PPdEcqzivBMYzkG6uS5c2QXcL1xESza57pCJFrk2YgYOeCp/1lHPp5
EDcgy9UQ5SHmtPoMDQNRFNQWvLC0xQ1TPoswe9M/jRu0+p5v4t93A6q9zrrm6V/f
d7waXGvA2VPfeZgNpRbPilh04wXmh5QthW8CDFxXI8WVQGwiJd0K1+Kpzremo93K
3SGiH2+kf8rOxUkoXPyxIOJIPrs6cv/tlRpzP/qh7W+hoV6ML9IXuw8KdpBBNrA/
wg3LncTahL1IUklhshCIB5FXTF84WsM6LFBr42dJM2odrVzZJX38UmHm8M0Sp1jy
iv9xQ6P36JnzaKVR9NHRpMlSffz/3PNgapqZnhXL6R1um1/QYPqlySMBEEclzCeT
4VMSC7Pt8kG3YPoGnID0W44WRVVy6Jc6ZsAEoSuDclHl0PSGh+mYcXIf2fmK8sCi
NHvTEEuJCQGSES6Hw5QziNFiiDsy10zVLB5M4wRZf1QM07LGBF7lhjdLDwAkzKsq
FVmWGUcdybAY9E4A8VlpAzFZWQ1dFbPN++JD3HiejowLYpaWMdSRE5BkGEJzzTjz
F+W/s7PGz1PiXVaWtKa8ZfQqcF0DsBoyKcOn1y/YcEeo9Aqt4dguNtVGdOtkQeJs
dHJ2+rJg3yibbL6hr+NdEwaEb2FDgKpMPdvh14f2jzJPm/AaklVViiPqZAbcOwGn
sQrT29AbR/P/C9zyirAI1XubrxsgkAcvOFrh0OOwd5K03bFlxVHZ6fDNp9lW7MB2
qkd17lgsmkGI9j/9QsdwxxIRZAPWw8gaoE8W9wMlnc2rYBNOksNpoqUnrgmCOBB5
4xEcR89cQRR6t88/WpPsyDKdlQ/HvvAjPkz8MipKR0ZU61UQghOTjJnf4Hu9V7yH
Z3sEFdq7/fzbLcXaGlUPcqgE6pN/pOuf4dsHvWoHirk83iNyvbenhc6b5F9BS9HK
ERRor74WF9dPmKUTMAW/CEPEqlAaakr/LyaGVVDTjZY3dNFevgNgawt1YPvdDxG5
EeYcCEW1dwb0tZdMfvWvdz/ApnjcxmBp2pzGSQw5nWILXOAhaz/A+wLLuWnvvplq
rOpdRg2Yry2tqxs8iNNefs9zHHeE6BZsbCkKdmJ6lgNGMAwa3sfmFsIsUIU41Glm
yaOGBm2wRTZ2BssRQUs08xvtB5JQSsh6ulI+g5I7JniB+CM2AOup5dlC60b3n25I
BwT5M6W4kMz2ml028m6eG6AuzYig7Wt7IIBWRp2dVTMVtogXpPXlkCtIm5WRIYf6
Fx7FRaa+8KEsRYxaPHCWccpi8Hi6hmGKX/PxQT3o6rhXq3ubs+nTUHHpA1NRDlcP
Umu9hAJ9pzhMbtupvt8cYvW4mCbxfS3iezkuFEp1lu+2GiS/Dtei0OBlIw0JY/1g
F2npGEfG9KI9Gu1d9WCot49Nwbh+GQMS5BqOUXw+tMuCrxHXW+P+TlmuUTaKxIZ7
i+fL+NXxCQVog8TGZSx0G4RF1bppGPqf/NaDDg1X/EBbr1LczGxeq/yGdqCSg5Xx
x6RauD17tFHjQMPi1I3i/0ZM5+a6GdsG6vTFxZETC3QeYnOw8EdD6ks5vqLckKQD
k+9JSCrG+F+cGNB9RwIQ+0k+PeupIYM63Hy+I5i3PCTME6J44ZmZASLfyaVlNwLB
zk/YbRgmdtnga5quCtqxUjPqZxxt+prx4cRUCGuzyn/20cfDbnqMbTkQzM7DbVL6
6JmF5syfo3vPYvBC9UFg07Y98JUbhEk2TT5h6UAimreNBFCrQPY5Khjk8vKlvYeR
DNmKSkiRQZ5PwG3KYqsdJQmNvD9V/MCX11xgLFKf1zi0TU9NqCsFKzEyqFpR6E/z
Xw2EVhjHwANTNkUEqigXJ/NcviHMrc9rPLD9FombqZ0LgPf6chQaM9BQUud3D7A8
FpxAeQLgT+foMqCVEMBMLREp1cX+QGAx7wVp8ORAtuHroFe8JHO624e45FZnV7IO
DhAAzdhso0ABTyyzl6jb31ydeq3rHUhHSx4ai1ezJ/PkTd4q/1+jwTZpSMBXrRlb
/YcIra5khPN8NTp3GU6yZOIuAyHWKaNAKAR+kAInw+mv3h2CVSDl/jnEtef4orHc
8PDweAcBj8zWvKGISyrx7qOqmgeIT+xaZGi97/z95P56vFO8Qq4NawtU5xD20Iz0
ssme/kjnG0vPfo0rpqJQZ+F9B/SzdJB5eMtpMLt2XlnVT5CZ1sE/Wh9EDJwJF/9k
VKfqRyS8ZAvHQqyu3gncolQLNsbqWAKj4jaTktz/liDTkAiPfpyUBTW20WS1mUTz
MTMLlGkCJkxC8nDydv9qCDcq2VVU00G/vve72kXXNjuTdaS5V/gfpmkic1/JaPPU
gPCqrqp28fjP4ntVRgWj2likEt/nW13rZ/TNymwcRJRUMd34wSw67U7vtVes/bSD
IaxGdfljN4gGjzzT+vAV/hS/3qc8pVsWdsUxUNl8na8it14ozvhYMKttvKAz7BeT
iyW1B7NGrPD8dGNHxwlbIXeOZJVmPwp0vQAb5oZiC2qt4PcfUJ2u+cklCfQUXXW6
7DYT/nzTwQHCqCSrHACyBiZjT/Chhc9ScHAXWmWPdAnbwE8NVqo9FzqYjKUiiwDs
ddGoRPvqdMfgPdN8WqluMF5P9gAooMbyJF5NDkEWNget60kpgVaOqoeguOfVsHpE
XivdKHHiy/l9WZqvzvf8D45aj95bJ70R6VG+u8bPCKTFCaDgrzq08IzPxaqq01Dp
14+/xYrVy6rWTw870vAffucaySlRbs9h5wHpZUD2OF8eMjDgUiaJPZTuvhB5chSU
FEB5cyP2aIR092L+92+6DGddIOJ7Q+S9L+dONGE6oLgy76ki+HKsBiPUZqFuKv2X
fhIFdllIpF1JKmgKlU0+ZzxPIvcvZO9Jia53wp2BvUlahFAf2eBHPfhDOr8hMos0
RNm3qMYMuwuCKS/9ljQhYuKfCLdKTRQ+Z5Wn2No857jO0RzXWvz4am/+KA46Fvdo
4GGanOzaEy0EHLWMTyaQTpggTIBxWxLqJ5HCHn9ZC7GQi6AimiBt3unUGvxv950i
7bX7ELNEwqDi+Xhax/VbEjm1a75L/UyWS7cqdekCmamP9FV+zlJggvcsXnruBHDR
qMbK20U7PpXC/Yh994/vYh1nolvom5R6vB4rT3R9EN9zC5rkYTiABa2Q3ArDe+fQ
y0h6S5JqphEB4XRUP2I/H/7n2IfAtpivAtZMqavJ1NRFQ390KfCWAelrXoDf49md
idr1YbCW/bjHs/mgz6fB3crKnkl7F8JJ2NzIB0scaIyRjUxjpnHOuIv/M6kKF+YX
BJBGQ9tE3gbrAuw0GMrheyCl5xarSUt3OM5caJuG+tNKCvnGq82qHOZktvfdx+hw
rneI/JyjgD66V7UxsYsNBaNERHb8hS8xJdESctKt6YY9V5/dUkPT1QOeC5QvgmFv
sWXS4G6X3YLuDZNzzppL0aZKY+si9IjygVRqcXtWLI6F3fvvVStYrn9y9P9YAmld
xmVV1Asecw5sck45gwunUe0t9LS7MQonjsnpTWp2wRaEMsrIybEI8c8yLqVIZ3Jx
4dJ7/5V3xlsbp5Ju6vvW8tAPpzm0UbhDE5GeZ/k2V3YkN2H0gB36cWv5tucPq5UQ
ru3ZjeCvKqwQvnIGBXHysM0Gbjm69LALo0V4uW7M1024VhFlGmnNMZ0w9d/M+g4b
2MiomVQCKvQkEtCHDFJ9I9/+BqwbpxbDatjp3bNq9mQ5MFZbMfAq84kglxkv7FX7
mkS08ePtIKR8UX9UbR+yJq2cvwODqbLdcSpFLrgzNjCYW1YHJ1G1b2t/rzovVcMs
HJuPkDG+T/BnFyG6e83Lyu1gdJCl9v59pvLwh9v03ODCSNrvXP7aXygJzzV1Lruq
Cx5hkTp+NJ7GyFET6o96qyGFfoWuzcKPLxTqT5slsrbgNrbIqlmuTh60aB7TEOmZ
mZIiK8OXNFfRc6nQNcZndNmTcIY2odEercgCVjkqvdYI2FTgwB4b2yQP9Z5Nmwc3
TJy9IwsLTKRHKM43Q8mOeH5AmPAdF3E2VYydy/kAIng9I9lDHAUSadUCX17ydsvO
JKxjf3sbnpj6UfuvKxkONoXk3n/64av3EhXcViIHFUa5n2ODPyWagUujOUzxhR+S
kcBvbHlWPLitoHFb/ZY6yQTm50UvFtsTLMRwdjPfYM/alZFisSbDF2E22gOwFkfT
S7YiOe6XFPrxpqJ41rPTKDZncHBW8sw0NXD0T/3lk7KYrdyMMog00Y8MNvZxxm9G
W21Gh4dQXM/poBCy49kxVvkJjrMf5z7QSwKlIi706krCawNU1L2dvwoT34FaTEBJ
cRWZFfHirK6AqGjCIKu7Xoe4HjTaXZv2+JwfOZtQilbawaVmSWJmLhNJxrOl/oX3
dI0s54U8e0VUSAEqzhGXZ70gcyHfl4j/GDsoneWTxARtgxhQ0rwf5fGw57CNvRlo
xG8GkBKxHqhT0+0deRw6q0i+i9I90+zP29tt+vs2uBQSwgyXqjsi2/kxxB5N9FhP
/ujHAUsCcRNQHO9BWZ4PtmgxUOeaMxw9+XWIs5srkrNVmMUbOB/lpZ3mSzt1tkFZ
P2ewscMmRa6gUI06XVItUcpwfSDF/VhOTAnvrbOP+U7TQBm9aUnKN4FOrGriuOHS
wyf2k0pNXUIdHy4QfULkuiZZeJLC+DworhdQJwbcYMLrptitJnR1u29S9YMXQihK
IEnDHUOTsvHcgx1jAaYYBGx8jtgMEM7uXqznTJ4DedVBbg/660TAB48xQ1/DZ+72
8GptJkssRKJjiTQVjg1RqpMwbK/Uhs3HjKsSUwtgRchm+9xN58dphbgEoDfg6dS0
tAdtSx0/m+TXUrXUwBJ82yv75ZUUhcDkAZZD2WdJEEKJKKtzxaZKd7Q/ihqakyyZ
7fcfj6yvNdRe05z05vn3zckB6M8m8kLIsgd9ZGeXxnK0ATKSRxVjTgKczvMdiVK8
XwmCUDsLou8SryEbpQm4fPOV1h+4GWPKp+fNAHgiapuQJWO645LZxA3+jZQkOEpA
hAQ6ma9HQFHORTDIqAY4QYbW1t3qjfLPEANMh8OhPBiT7/RZwuoWhAO1lugXVLAy
Y6RFGY7T3uUd5GxlVfCF+Hd1/NKWIMZIuS2VgJKsUtW4R2kIfkcehqH1prFrJgAH
NtFvPLRgTeIkHbd+ari9LQRaU9i8tafr1uEXJbFyc/D/vmQCyIgh4qdoqw6BRdoI
jqohE924AMvMfZLxR+xQrEoNnDLGajmsApi2luBOjQ/4ZjY3/69w06QKu5g3o41q
KaihQ3fxPx4c5Lmx5LIU/qeel9E0njYkxiiBNEIR10F7wp1QGX0t/p5p3Fymr4Wx
eiV0ejAtUqEbeHKUi6nn2rNODnn5+Ai1BglOBRnCvd/5mn5xo21X2ZFcHnJ3Ykes
xSma1lKumUvNoB6Haz5igkiwyK/MZ3XbwpW6QUICiEOwhe1p2TYjkLYhpCdK8eDQ
G06B5Rr+znl18PYMTxMmgDaeoHkNGgvsrNDb+m58pbFwuwOpNI1OJ/NSGNUoR2iD
ISRDEgXID0pdCo0Yl3ZyqmEF5X6EXsNkcBUji6acUvUUqNRvqzGQrPGlG1cbF4h9
F8bxQmM4EEipKm0S3SAY6lAZ5q+iqy048C5sMGWFJapxus7BJ7tyMRWYDygI4Fxc
Mll75WjKwdcON+84QPYO/646Ig7UKGXV5KOxUEpbhkYPFovRDuxUheqcFJADWrcQ
MM+nLc78AAsvJe81s0c8pAvUyOQ1YiGIdNbeRm2UOoh1mUw7+nbR+gJmAVu+2lt0
GMeihXo7/xyEVYyODvUkz6YJ2mxRc3CyY6rk1bJFD/b2yaqhjoJwGuQdTPL11uOF
K1FzXm8AQo5YXVGU9JjmK7VbZnAWuq/Ytm5PbHwtGMyK40LLaYhGcfx2engQFERY
XnaqS8cwiIbofEN+OUuGiEUaE6Iolihg7erA/9mUrj0yhJdQ8GEWOzO/SEi0hsQY
Y0p6xz1OulaV37sBkHmCvaKprAHSZaBBdCHxzd4kn4Uy2yIHwnLssWCMzPD/XGLT
tSMcIHEQXK2KOn/O5yf72a/YZ+wS67pjYodzGLxnjzqjOrhGf0Mkehm4bQv7cwZ+
WnDlz+Xqwnw1XFkZh3X1X6Rb/pHk44mtqX5SngLNsl43B//oaBvVfImjagLiBk/2
e4rC5vUhKCPPEcH0+Cuc35vuIzAl9OJWUTth/WOfmZPHdXgvBdyTsliOCZU74nEP
oV7L9YI7qWhOChkoCzCQENpoFkeLwySHnyGkvJqH50f32jpBuRQxHfYi56IaAp8w
vJ69/QWmEZR1yjByqll2xBJN0GqcF8Dr1cx5Pdy1uEtRbqJ2kkhMfF4lUpR09OSc
ya+O9wARGOyKbCbT8e8M4w7Rt21viU9NLDT49r0MdjphJLPe4q+SdcuL358jGX98
asXizO+k9AvEbs6DWQr5P2a/D34CNDD8N2bisiGDTOCu7wCafEOqjyA/fj9D3z+U
WJeiPjwtT12hDCeGeT1h4Fw8sQH7s35m6hS2ElbdAISx25+waOwbkGpb/MfCGLJe
REMWmeOMWImTM0YO8sRoHmDg8riMXCUVEY1pOOC06KbmG3RLRENiAhzABqQPsH/a
qXQlP74GcDHr1eNkoqY6JJuYF2PjCvZfxSwdMsHnlR9JkK8i8Yzjv26ygBnJatHM
M7GjyzAyQPuZjdlMcmZl+tYKdCQHvxjqDFkAup1ZUBN7o747F4e5DJDDV0DK1D9Y
mUCuwoA/C41uN53LTqb9Lur5EO1W3Utw8rkWQ1Ib9VRU5y3JTwzNuGuUHAS1A6lj
sb9jzLxk/sYmvdjjDKBZYZU+nDiNRUYb1/CtNFOHbGNTbb1qmx8AuveGu6zihPhA
tQxmFrrfYO3YPj0afVRxQYElOrRPV9vbjwYPYzJtgRQbekUZIz0yewJscTP1uK7V
glLZ8TwWhF+cENoSa9lajHrZCfkC5sHyZquJKa3kHSUDakKiVzVj8+Z/NLs1Ask5
wdYlji/Nbkwm5GjYAZLl6/Yry1w3jE67Qnpf3T5SgrYSl8PrH7YK9y2yyxhgV9OJ
qxKbeQDSo0OjWBe79ZLv1SMmu7D3e0IbMjwFpq9VtQPnzscunvVyjYrYrhRet0Mt
t42/BJgO4DY+95VWGMDw/T+OQjwkBiUlm+ur5oZuijpqWneiY8yz5Bfoy4uiFBnu
2udZiLFMoRKKoQTzxqmNJt9u8moMqtwjfudnDkviW7op0A4KhzY6X9MokPGdnGK2
OEmxOYB7/oOm558dI2pgrJ2lHCny+5FVfjE4nEqpWMdnQ1VmnmnphAhQzsjDZQl+
PH0EBtbJAW2hbWUOoeiBSrJ/0F20lrxsvflZiuwbrZbTN+pQDsZ9Xot7Zq2sEGic
oA7K1KnXMTavHrWP6CF5N/PQg+S4x0+0khnNwd9tVH0XqfxCSmCHrb3pJXr5xjae
FrLmWc8PUjoXljzSZiWpQR3PLxCenDpygwz4iwGy231G8CYRdi43xJ7wbZ6roGwF
DmHgmRSZWig48VHJONuWl3Gj/eXNVcU4rel/9p/1+KmpwnLNj8zC9/m2RfEl1uWj
f2scb3xe3pKIcObWzDDxNOYfjoIXQlPmIg6ca32LBuBrR1IN8oRx8+dH7KODAc4W
J1JuviGkmL99Z2UX9eoGWFBVHPoAxF4PbPwAsiRAKxvBk1XEtRKOrizrYQsMha8C
4yzt2fXKMDwgHCquG6Kpl21bZDa8DdNGPtjyy0JmVVGPPOuOj0u6jRl+A2wTgva+
AvtrkQCBNbAAM3xHN/+ZYFCWU+DbQXPET3w5DdEZqN8jcdVKmDyve1tdBtgtr04p
mAE2Qw2Aufhip5JaLaGuOutxDm11ErRCLF5j7ysobyfEh1wPc8lCkvEae6Lc++yD
xaeO5l1Zm1H3Xa4E5o4HZiFjLNQ3QJHMfCRV1Tn6HgQi7rlRvMoCPUK6rgOtGkGf
Rnm461Fo2N71lHBB6WYJ7rZAcbP9LFp4wncEabLotxzPOJrhnGFnMekH68/jP3nl
cOGBrBNd0IfABZP/PR/SULHn0Itn1V5QsWQjVrlekCDMrgPenLXHZrIxTEoT09cW
WpgcenjWw0pP8Z/kABrukmt9t+EWSpxDWOkt7nlFbY/pTQZxEVn6qR+KO6TNVO3y
eyRIvqz2smzRsdgkQEG4GCSTD8RWnGeIsUMqbXsRY9E5sgP1TLlAjnNBYCE9kwYl
jxzKTBOIWx+RqyJWtzbLIFOTjgNaaloUoTuXEGY05n6oxrIlBnS8lX9/rIk7bMCH
GME0YyiP2yXuxy2G+7WuBScmNS0ojWfv6MU/fv6NfJUS+RNL3gPq/GHzTcGOxXD+
58IjnKy4d5ZZlktqb3EcO2z4h4jKpKhKQ1KdJRNL46YuhWgmJPPyiMBijbfjaAWj
jB/j42koqlWNLkc1mKJ/3Uj4JZrTNQdfEJJiZ0fuBV1/QvfaOVEDMbqGPdYteO3r
7NNO0E8mAYqfTvMInpTEdCUUVgllhFBfP5HlwgXs7SJj03Pxd73leslpaBs+xS1A
+B28vl9SNEtIihXGJZM3pnmXOpMcL49FwYAQmzkPJ49Hm60RJRYeve0NCcC+wNJU
STCKZpoz34ZGilpZ2MErP11Nz6FHQY6UCVao6o2Y6vL2rLJGMbalqZy4gEX2JmSu
81ViwIEOlU2ZhH5wMNEqd6orPa9sR0aPjrlegiQ6Zhkr+NAElW+btQ6oXoFEGsYS
SH2nwJ37KJT590nL9aA3MbIqHj0wUVFn0NE+NOVB7V9KYYY5EIAACPCEqbfVbvgR
XAQovcc9c/FmvJbv97N5N4yz8BrKvObfTmKzVTWeiUqHUD1ISxCYlqjuviMsKEP0
9gU27urmwQ380VcA+uclbUJeyU9b9VXaxesGWbhw1qc1nXeg/Fgq4NKA6NYrkSQj
YsAzetFPi9mMD+xol2+RHPJrRgLMXbPn7QadXarweNk6bajpehjiQYqDt1li57uk
xFYTfHDmhamjYwfUwHHxrS2od8Zj0vAV0juRagDMwG/XuYxhPgRSHwlCd2bSPnqj
Eb2QdUxjHpv6VgUqA0+nE/oSNj9CXVIcNKpPSF62YXujkepqFJYB2X9oow/MDF/1
L3d47khtxqIbGNIv6gxpkDoWtcglkZ6r3x6aAqTsXGBgDcnsCTn+DZJZvVnp26Yf
EgGE3VbAOCrY8pZxQGwaHPcDvOSDKpbZHILrtpS0SD3UVKMzCjHCo4LbqtK4dowh
CSCe5IkKVEIg+yYDwOd1YB9820miJ7OB60RCLd3dZozubwlcNKKwwAZ0KDbv4Xcp
DdE8cBycsx+qTgamajMWLMdE1SmPOhYI+K+JvnqIs/zn1iJFt8lLM5ZDhT3J2VJR
hBLh+io8fPIdz5sTVEc93DE5crxhdux2rPeW7g3j4jJuRYVnM0m9qZaYwaqhSQN/
5ikaxAEOQvty+u5Ty87jIh7BJtqlu/IFX7flR0cIIWIYohV/sX60Y40gJk4ffmpw
X/wiAsKgtgkGa9Ujmb0/EpnC7gyjQLXenIz4mwkAvpurYbOzi5Tq0s9fnt9Ho6hg
y7ex+9iwxMVSUkFcMHi4orcqPhjNqMuWbCAffgG3/KIhPXMeKBhHCUMEyOv8uDTT
7ROFELHNgw2wA5+CQKYkJTevxgMfMqLsS8aQhr6L0ZOAOLVNiJXm+BFTG3L4d/41
qzsLlLNpQ1LNl3J2B10UAcl0t2m1vTHh4Yt2bHc9QKeN3wbkzax+8JPBE1r1gohN
EVsyMtwxoH56AY0jhSNvZEikKh5mbj8/zzwI/nQeqtYLb9ObSLyC126bFKdI/GHl
1CbWJ5RqxQnXHJ6mlFQSHKHYx99T0+uefHJc5zAb6BSRR4BtZcvIPtuFKvwE88hx
MgAN2LDDgq3YpzzBMpBlnSbQdydTAIFnMdVBUtADgNugC/mzyvnabHH78JQo6NJ+
EoCgrnrNgSbi5Uz0iGsf7Oo7Fu0vw9T2G0UngHfIgdqpnSrHoDRFoS6Kf2L0eRrz
mJIhzjEd2hW6B4IqdPdYi/JDxBx0V3nRmfGdBbGQvAQJ2iOc8vU3fK6CHihIrkfa
JIAOhAlvfWF1LVhNeSIqlC/RuQhIW+kLIKC0Zgh4n3dkb4IkpITnS4auN0qDdXxN
oBuIdPEbqST+zzzZie8suwDLzYflxiPVNT1sl0rtrJNqV4Z/ZPkSQa8bQVMnTDYE
jmWzWytlBxg3dgljXoZr54NM3vMoPNG0PSftoSZvrbI1f133EgXiFOup0uAGmfSs
PMDa5xed2pgbeLodXylHrQArBK29/gUm35DTATMP00O48AAWnKa+L1kSBCSTV/Vr
3bPnxBVz9w2kvAS2/Di4odbdByO9zY5sJWUhrmMqQPfjjmYmoYX2PYYQyHtDVCry
yI9CuKqLUoz0AWZiAPUrRWoHBd9vwgu9036MqiARGiu9yambpjhtNvxdbb3nw5ii
Q/GFt42VwaNf0WaDhLDz8A4pl4MWv4TLy0gzqE0oolh+1CAZAtF5OSAHEuKLwUXw
incyTCSkG1Mtf9qxNN5LvKLbiv0UTxyF2B8j8ODiADcW2igwppalR0B4hYEKSfu5
vgfCgLvj1O3J0TLibjKFfRgDV/7bXv9lZFxV/eXcjBUtLRJ0Tp5wNc00srEngkxD
p7iyWHWS4ECATpgw6+5h5+hsqMTZe+bVAucGWVa2AdfnPEoXM5Am0yf2FeSZ3iAx
BXajEc8ug4GOMhN4ksIjRPmB7S8oM1PvO45Az5ScpqcnLh4CIJHVAM6Xmm0FnaFu
v7CNg3bqWVYnvNceqdaQ44iDpzlHhwJVQxzzxJxY2ZKQqc+uNVI6RCydDzQ3bgwG
J5DnpcRK4U+QxmsSgfUD57Zf6VFWXbDioe5qTyfyCSq6UC11oPqxyotJgLh20Mbd
Zu0BrEpJ9PrhMm5yI5LV+SutQbJVThELU4K/SY0DJrtHuZSwu58xfxyc79zpg/77
qwTvA2wieof1iu7axoQKo/XMgYRe2BXiR6lOdP2Y3FFxB1eHF7oNdmMwYmFVuopi
PKeo1cM82cffRfIH2KM/QXZTnKXnD6qvzTNo9ax9E9KbuhnBSUbJ2g2mjVwDL5fR
MhOzU7IndAv567tsIiXOHF7GmAtzCYDNAUxz8uwLdi1ps1MsNkULIK0NomfniR3Z
0aGROw3faZ05xKrcWW+0wdf4cOCeKob+8FLjDEdvIfxP9QxUnQ9Yz/FUkD/pdYeX
TZpa/WRH38mQUtm+6b8L9QuCLlt00Plsp/4m2siS5poDvF+xbXBviJ6grSZ59Rd7
MdqJhPirVJY7KQZOZyiXgOoXQjh+ZH5cNq3zkZuqcNiDy7SNnV2I3L6bk85fIAIB
K68HbSYXi7Y6x9wlfZq4EGMHC5HvUi7DQ0hxUUVGAfFBmDmdM1bWGAR8ZPFVcR5V
Z4VWUtJLbjZ04YedyLvyZVnCNArZede28Q3VW2Lhp5M60Zshl8lg2HKBAtntxMTV
kRXusJPeoLTai0aWyl1mvhhvKkisCg4SQL6xwM5Q5pPSLa5ky7clK6UReozILXV0
xVJPhKAu1b+Tu4rr8JyJZbjPcylMJz9IvN4ROdJ2Un6boPhyJIKK/DUYO0AisGvP
DOYRCE3jJ0reKL14TVoriKSBVQSMQDR3SwcBn0Ky5VXUtWmsgZoBwVe9PLPr7KwT
52Cff3milncwLoiwLxx8yfUmSez8APQUn3kkBM+XkGMaAbWyToEMLTj9AC7msKqK
rYsp5dZLAS47BIQQQi/9/vzHuam3KcpSrNYplD4uKHiytgDi4QW1pIyT3q/B92Jd
0iQG/E6eKiNpUCKjuQdP4RXlgHxh5ASo5cH3JtXpcQzPnJqIkoPgUCeeEWn0JAgj
L2iKlcc8Ekiw5avec9/p4JsCykoAwvE0vA5o2re6IJxGH2TfPhYaIm5RDIlkpNd6
K9vOnVzibOXdDvMlK7H+o+aHDiCUm+yrVqix88CEHS2//o+08ewN1rAVsFTfHa18
KqlGTPhRDrElDiFXMWJMzqPZBU/hIZZ+cTui/D4CIkA2crICa/sWUH93fL/qdVQ6
t1ObNISvqUGs52NOANIgB9ZQLqj0RJUAz+8XSPo9bWOB4DJ8oYIDjnDy8dP8lZjK
ob9OmRsTWpwmIF/ozTGSOPYFVFlixNaXZzNwpuAhO0Qs4uQWg+22+qs+Enzos9tX
b+D+UpRDWgFxfVHUoIuSVcN33S4u+vBGy9ph7es5VaLRHfY4RoxaoHf9d/bqgW/P
fX+3m/JGNv/fAUabTnddVDp0Zx00KQ8gmHVsoFlzNDA/u2JzBg0Rrm9fnJzuyo6X
+4+k0/BJc/x4aQXgxlmhIXhKjotZePSoeU5MxNlgpSC8vOYtkJaksHXo+BtghTvl
+DOOe7ucl94kZ/+zfdAeYWbDzbcMcVfm6+vyYSuEU9CL7gbxec+HQ7d2yb23PzS6
y6oOVnTZxDW+2lUOLCKtl8gT2FFDqQ7oLTGlmmu7XQqLtEtEGXwWf12y/d62por6
GW/qqtRsU70lJ+kngcx9aSdBIxW+b6pQRuus4A0NJi7waAKB2o7C0Q6mcUs3yjbV
0RYEKuHTTOSPn6wmUrH21538RLmaiX6+9rQ3EzDx7sRr0UL4rJK8L916aVABlvO0
Aam0Cz6QXvkSlkPxRhsVsmJ7GRaP5BL4c02bXUGhTKycQE2x5OLYAtslexH4/p1O
WYA5SXThqTxdQI/NlE+ONm8hsxPHkLvi7BR6/T31JRN4EZpgq36h5ker19lvrfeS
xsl6RDMSLOB2Hu3md2CfGatFCs5Gnp6vruNZHZN6RMi/X4XvYHGpokr7MHDOU/nD
lCi7yM34loXzepv3m/snRj5t/A995U69f9dkdI5Hgb7eqLAAALKJ1Vl5o/OhhFIS
htS5raHTTe5CHuXUVCSMZ5zLxSqpLNJuYJBTY2/PSeZEpV4Q3GR6GJwxExHz0SVR
GeZIgrb2cirp8iuDoSDvuFIvZYV4gmwyOMcMBgr900h65mS5+BlfUZKNVfDhNTiI
RN2FUpxsiwZxmP5zFgbkQUO1UHjFVFKcBYwNnjxUeDr1BYdWvTxAK3Bia/xiQHcn
Ya4Qp+/sye+INCl8zKmpboxjXbK6vLuQWXnf1xYzfUnjNh6Azh4M3Ey9IQ8+OEXO
1VP2rIqjfna65UhTiqQQglQ6TyqY7FGnSQVuNBTh5QkhdH+6N6PtsdW1kYALAbXx
jogTPrO97LqIff5+IhxjABX3qwRkcPchOmCq0X5RT93PH8NpgmfudyO63j+Y08Mz
QwxWXTgRGHXoO+pawtxo08qFITC4Iiaobbp5JAke+HoX5AFp89du8lPQy4rnYlCp
G+L7AkAyIGno98yd1BOPI7tX8Uw31Ts+KaMq67zTcEwRM4Pes+/sNAblD23wpfEI
BqXiB2wPTIj4pcV8zwPvovN9xcmJ1ElqAGGwu1D3W9H2hRO/rxSJZACxBQOUKZR2
U6GYWLQVd0pxmOfgrgvrTvZO/OZBLD5+P7gGMrUd9UZVN/JlRdoOiiaUNBata5nN
9K/KLscL/HnBlkGtbP3TEDheB8v1Qp54TZ93ib2t1spaZndM2ub9UQhbjJNohifa
cJlDfcLa7pw6cR5hSBa2vW6EI2hvhnL8ZN/EphcpMQsMLjIRom2NejC5cOzzvIFD
4wJWageiCypgc0PPJKQYSPLpxdbBoFomaRwHcjibIybmTJGOXccG12mVuNgmsEx0
3Ss4+FPT2LFsZ5seSXuKhrCy+U8ySqod514+CCem8+ZD4o6CMWn4LCUDWstiBmb7
UvoPe6ydHSm3t/Kb12b61bfeWiu2KmwMuxt7qcQaH456MeWYUpvnMYSKo+/rfQNm
AIsRIHyMEb7ksS3jJETNS59+lw1AYf9r+NzzKTVrFRrGuecGgqKlsfJ5OXX1Sm3p
PrRA5HFOe17KD8khKZPr8AMaiotLLD+AmGuqJwgIj4Lha6qraiZSW2+t1omgI7S4
72XlWyLL0N/A1qv3T7Dm6+oXG0Y7JXhh9uFaiGyDHlyBDgFwyzdYieKnUvXAt2x/
ihGjlIEIRXGSeTvYHi4cOuDLioWy+KpoD8cQjVyY4vywETcrxw8sybpdaJmoIgOp
kc7+4Zlwi0izZVoy/qJYA3/LI3Aa81TJ/RZ4UG8M3NQ6DUVeswvcbyoSyGWQmKbg
sCjnijrC1+iF6cG03nMUzCbThfxcg6vu1V2oqCWk8EtksHWZtaawsOZuq7dZti9z
BynMmZeAlCA/MUqc4ek6cXsD8WXHSGenloa6LrjGAZDNaKEGxwNUNG/n2viPn+v5
l7OuhHGCYuR38DhmDW5YF6Mi4el1YoUNRsoUzn0RGLtCmLU/l75GuZbZCSghj+oE
2Ip0LcYLoRryRV3dU3N1M5muux1DTeS2Wf7wNv7pIkhCTfgilRF7cAUHwJfggpv8
uDujhZZ0C4RDW0SkaduGuwa+T3D99Kp5iyUpGOgdbdT1nrdN3LCUEf7RsgEQIjQZ
7REJKfplPnKEYV1EuzsQw4eV6BV2fCBGyOFo902kiwLh9M/JNzJnNvuccvTRpzGk
V8QbV5S092WA3bTrDBSfANyGapP1+/hHc0s73jZ+ELOhIqzWLAgJGQvAQDD+v9Xy
+uO3H402mmprr3Qvfn7ODbFnjFGNVAAH8w/DXowB+C89mAW89I7DVaiSeJhM9eV7
HEokPCZpPsz3MJ3NEBnjfvXykIzb+NNA0dS6ZPwhRiOX9fxl6BQ9JZ9qQvCiDDZt
liAI0HXTfJvxJ6d1gZQ1u3zvpaicdbnhzIrk2ir4nLuJJvRVUDuz30RL7NJwa3yt
pT3GWx+6wIkRVKh1nK4x6VSoeeMwQaYHnpej89l5bKhqKBGXEED7ubq41cefxONX
EiWVyIFvRTDYYuq7foah5tOL5AlDorfH6j2ettgv+vLkyWpZLkRae7JIXvmYHJwu
6sD1yY3FOxxEg6Hk9qGSVlqd4T9HCh1WgCywkIDFeAj/QrkV5cuIE1Uhddw0YcOM
pzZHuv91ct06XYr/8oFbfGixpvOOeNZiZhwz471icoGH99c0c/rpYpig3BJ39DwM
ZEYW8pq3I8nLzlugLl2yCrmbQ3+xpgDIiFPLjCunmKfD/RRWykUb6f22HAsLolOw
IjxvUON1ALkRmWCPV9rsRYWwq6jO4m8XJ3u9JnNhHQCHdhW0NjlHySK2sfcRHZh+
xREgsRjYq+4wOLVYmJOWKktVh0aTFcQSI2KTAfKP74siAs2KBv4f3DStI7ZfWpGc
q1uogaSAtQy4jeeA9QB1nGt0IGCt2fntSiOVlbxaTKVchvps7sgMjtroTFI2Iixu
LAG5fEgBeayZ7UAyStIK/8ybMdnh/nPHxTodagoodX96B/ZBJBCK9ULrHi2WRoAz
ypHHKqPjmGV6vVk1X0fOvVvSBv34Oed79PzHqgeiUpwV1q0wG5gvayvgCS3xS2hp
5fh0xcqxx7LLOtYNrzfjt0czzBrzr1sZNwrDgu/mru2TA/Om9cSA6I00MMLBCrfT
MA82iD+7v26XyYG3DG94RVByk/i+u4BfXou8O6czfwkmWkvbH+fKYW0Rd2w2FFal
/dACfjS/NcR1/zhUX4G1knCnAC1YjbK6FZXMFef19eoarSqZJaF6cqAnEtTnOdGM
ABvjry9LcIG6ELlfPC6ZSNrGN1w6hBeaQOGGqjzBiBCP+2nOwH4QTzx+g21lXjwJ
wRZBrmXx/Rew89+TBexpn9ijtdNZic+srKlH7nghYyztLcf5IfdAfJXy8Rz+MFBU
uit0Args3Ne6VNPR6nqDWgjOBuDB165hesU8HuWrMVHZtHIOF0sQlxupf2hlmOgb
2zS9YrlngSmqkg/cFLdeW8v/X8Ual/KqKh01VP2ux6jBJjXzP097Vo6RjNMj4q/V
HwGYp+evbOZXTjlDZCfGXUeIOE5ZDKIrocb9xMcIYN8nwRpN6Cm3xkXqJyEksLwl
DbOydgr6i+iLVTjulABmuwj8TCmKWaXAi037Bzj0dykDb+69DAeR8jEjxB2PzxCW
oSpuaB+GUBY2PrLgjgU8qQT4hcFE2zxdOSQ54TsE471C/9YCFD0qL38W3hyGFsqm
pnairAcHupDMqR9ULk103c1uzdWqZD/OWDPmgk1SiXiOVnf/Cu43NtEDsvL5zfHq
vP77wvLmb/JLiRGCNyQZztUZfIiNWSHFZgThq7ud1hNG/iMKbQ5t++ASVwdh+UOs
rNuRA7/33591oY3RMNh4/dMMG6jn6af2NkuzoLdPbNhgoK5g8e+oxrdGJhTfUPXq
F+e44P+1UPS//L/oxNNoz9KRE/HAvL9b7Y5nWcyMWP6/9fO8RmE4NQzoo06z3uHy
B+kWagKkFSVJujbL75p+HpC04s9ntt2a/3gIiyy3/3SKoMlFEknk8UDfwBBn6zAy
tiKqtJyfxgfvh1SDN3CQ5jVICmnFT/zomv+C+pZBZ83N4bSpGepmgMhufjan0zFr
0Ybs6U0QulcVedbRxHKwFIc0UqDUtqVl32XfARdqwGPhTRf9m9yo8/cU7hdUgIhD
mVe40nFEYXQX0NEODqhsckDsRrxXyHotsrvvTNTraz9X/2m1h+leHDTg0RpT/sUo
NbPc4SjsSrrXkvuy5pfj8iygpDJkpLyLumZltDP2t08JaMi8EFPnd7mdAG7Nbdo8
kM1lQHBkuHAZk0t2XDxqHJFbXy9dyvHxnZErbvVnkDuSgcwYivYPjXIFZUi7XTFf
CEkm8GMPycFKqFbY1WwSpZiA3MX/NkPAqD7bs4LxXPGrKmWnME9JYjmPmB3c11QY
epc0z7CapZQ3bWXQVYARdXWJnBZSJ6hFCd7MNDhHgEWvU2LMOwhnA91xKu//FeS5
tbCbRBlZ4oAD5ytjFxj5ZpX/MvXQabG5bIx/ug4fja4g1qbAveMnWtI2MxBkrzn3
tbHucTInEyeSi1y9y8eKsh2QamkUbS4Ja4PWT28Koq9B+Btlpr9+o6pfEUr0cetU
ox3A+D6hYsIEGUCKPpAHxS7G+4rwQCxUT9ziaQfcSLUw86/yx9y67CO45gDJsDUb
neyAYUzTcW57Vc6nsc3Sf2VIMwm6C80C+4ViugmYNsd2mWKMxw7Jx6EkR0sONAM0
Yxg1soxLHVH5SCH8PmqHhuJTq1Bd9ZMJZVSOieIeKcCh9e6iwOawkYLLHEzBgyoT
XR6IksUuRelSCYLznP7+ZqDAyZxB3iiuHEaLUtHUNV4rG6I18tdeXT8/QCI6iTj/
trfZBBo9lWA1QTWxfVHzjxQ75rMX1TXPXUaAFEVRQ0jdELJ4TBK8hNxDc9odUDck
zhc7//5lNeCNrEVYzIbqzjW/muCiI6utEjzrGaW3B83jzCKlAwukJo5Qo7HvlO57
wp6AAfDtgTyLEQS4qISV9+/Oba9JUcp1Y3r5TW+hl2r/X/SyK6dq4rOMwGyQcVwB
UNSvFtvobZKz0NNwkCG8azCbtP8vMDucFYm75fJY6k/bi2hA3U7YJF7ACrWMaocH
Vqe6SOGrvI94/Q8i3qTDRWk2tACbdgHNSEuh2gnh8Hnpfa7vGs17bYGeYXqJRW0Q
FD17nMz5oJJzMUrVng7G9FLBleDsjhbfqRU4TYdMKgJA1lITDw8kDvtLiz3C1sUD
TFwyaaiT2xzKCP8w5cDar4urc0mVbKklQtZRFRzbpNVwnmE8slIUod7CgtDUpFVX
IjRrDtuBDC/NF4BVBRfmSwYzHcNv+rnWaj0qC+197XgsxE2jnErL94KFBThxg84R
Vy25zz97ro3XZVwKyNJ3m2twK8GHEHjQznY2QtOh/g/6ujJCQVXzuZ6220oLZhc0
SDgZZk3xjFXmawFgma+AvZPJCKEguDk3ch2EVXMQUD2y9Oc4z71jElPz8dN7jfjp
kG1JZJTCyjSHIGksZ5zN3EsXwvWV9e8gRCKCZSI3kh9EsV6NaCe4UYSbbs/mKplP
wkvb20CNklps4sDknV7m4tEDsTVaX8s4i20dUehAPY1QrImkbUy+z8yIL+OYF2k8
FvnHYa7xtk3VJ+yTyFo7qTT1ipZSiMXGfwn94sBt5KfNdajYDIIaNm/VT4hJa7Cw
M8/hqZg6ZHST6OCAbcT8LKdBJDGkCqzfBXet1yG+LiYNOmmC0TQR6pyyylfsPDAW
x8wNYQ/uQ7URqRDsB7yAqnMM/jkhAC4c34bFOuNFBwVnorfnR1QfjguK9qj2JgFM
Daqkt65XdcdwM39JM0tE355bIJbipCkypUDQOncEIsQcZvu9zb0v9f3Nl62I7qzb
xjZ6D21xnEXKTahkA4C0DFPFafPAFJcYR9cjWOsWBYcwiNGfPsqBWWc1hT2Pq4Pl
+3WbPfV0wp7E8OnCHv7KyAqQUIe9MYxkmL2/OqIOOxvYdAr+BPqWy9Zi2XyskQ5r
PwwY+w2m0bCMMIfqH6Uti5atgpORcWGMft9iDQ5YLLX0L5T3st2qRXLiHAZZHiCr
awI4j7FrHJms87lYNggY+tJvM2x+E4NSaVzKhuWlkVGPldO7X35PURIypTJ0QfDb
Fkhnnr1ierhuoZKNp4/NvO1ym85x3uuHKn7rMhjkUq95Ej9QQ9K7fyngYUNvLw9y
AjYhaRlWmT8S9YlSPiKECLPw2zDs6x1MQFKFqkMdPGrtEl6AS2euYL+fsXofwYNB
QgQINU+2bhWia9b5lywe3Iw7ikVDJBq0u5A9AnQKszUHDssaOEVt62aM6NSEjQio
eJFu9a/5sMsb9+igg8c86SuNYvNqw/O6gl21v2QNd2mZbWkMyqefeObytH6NAHX4
WINK7ZUzfaFCLDzwnyPCl89VTqLeZV2yTOVEGkpXoKgDro+lBgkgaYwBU9McNRhl
sD6Yc0fJTM5zAsUVUkqNvQOS7Cd7Uw2gG0GXDdGC13FNbKEiBpDBIXFOns8fxLK1
w2+rsoLQ/nrk4bvBhvpWYXeSTViM+1Kyc4UD/zAOuf6OA4+D1L4cykx7Tczh8ruQ
OwUIyMRvCvJaYEDULo9DW2rjMa6nsIPGoON1/9TCusokUNaAOH1Ska+x0Eex1sPs
u0SsLaNOArc0xiLEaxpafluke3xRxygE19ATZj5QrIT4kKNsGU9BScB2eiAVqm6c
mSqGCRZ6dvmKHdxHbvvVO7PtUlal7YieG/IPZ0h3h0zOAjmA+Lr7JWqVhDnMLcQZ
zVNSnS9BFX1Wya63p9vihRMo8pIrOANgCXe0eb3UjJgqglVxOlcko3SH0VC/z6PS
/E1uNJpn2JfNtff/uFs/HLsk0Yzikki89GspqFi9JFQSBnVsfNYFvCBdKGFo6ORl
7uHEgzAQb11HoEg0KDLLDS9tPdGJ+rAGqZyQMOnjoYqaru/XkOkV3zN+g9++wQzc
vDcveg42mKJz9Zhy1jXUj/F+BilkDc6ZTFecVgxZUIov4PCVrjoTceqPb9U9jFMz
c99H5pZyP58sBxJsVIYUrZab2PxucB3e+gWlRz5Tauqimy/L0AdGuwoJk7TwnTvY
D7/Roqf9scEMC3jfuYPrZFAdVXcCUfXadCBdlRkAQetv1124UHhuSpiamXy/xx0X
kvOQ2AALSc/ld1nKEAyzgPti41tKGkqXqLqC05ucStsQ/EqIi1ybjRLi/d6LGyq+
+S+8PAhbposkzRJ4B0Kd8+DKP7Wg0+td8Y0FfHDVgIew7Qh0nD0OOy3vw83Zeqfg
Odek6spJpCbnpb6QkWFDn13x95xeOmoMLBlAFI7A0JWiWt9UU+2Pxoo9roe6H+rD
tt6c2no6v320cUI3IkK3OJAppQmrVRCCD66UXSn/xcEnoXhocDqAoKJ7JdnNvYoy
mStXzVoBqcwctLR0fN1de+y5KSSO+4XSF7xlLFWYA2Nnolejmo+uTNhqbJF+dNXc
2R0bsIHvR59u3zSzIcAV82MLTy/IO4iVqW38kPqqCxb0cPUveEUGRURKs0khA5qi
FFbsVpWtl0JR23yHGG5jX6CDrc+5YRM3/+KN+JW0qjcj8nE6vsyx1zpSOQ/eXwX/
qpPnXWRofhQDH51vDIm+JTqxjqcLFJomfCKONT1jIffloQjq6R0VoDD1TuM+n77a
A/xlXcl4PR5yOry6YD6ls0OUT5BHHmXH7HtJVkiPXOLA5ui1pCJQBTqL3cb9eH8L
or/BKoJCsxJdXqdPqpJ2VAtHXrkPlqxvR2l4DfnQIKfOTobgk4uvLPWn7vhnSSMz
5qzskE3vHM73LMKC/KhkmzOpeOnEQGCamd20POVlpPqD7LFr+QKaMnrVcPlhn9kT
YEKS7wRHrGU4gWdl2Rk8t2KAf7yCMDGdPCHqQKW2nshZj1SEe98c/DUfeZIjzPHJ
H3g3QQF9SwwlDm1FIPdAc9skRxa6FPNvqrWEZqaCutle5W5kr8pa1Zpf78SqTqb2
C6TFhb2Rvi4FufOjJ7sJuFYJNq4u27j07BBtscK5c58lkKU8Hz0Zqp8rDm5EB8iA
hiQvTk34DDrIGbBP70rlJ+mN6O1njfZR31x9G8H6HMGquz8VknIBKfuUQXKzs17G
mNOh/xDFwzEfMygtWYfAwGvFrBbcOSqcHqRHn66bGdMv8WG4tA6kWvyDwwmPc9ZG
U0WVf8VH7ZdgDvsxfiiN8+vfe52gqX5+8dEuRZ2MI8RJ5yo/gSG0TyNTTaFgBts9
dTqlm5uBSbZRBiqIGjnpdO+net/0EPz+A3J3WAmPRm0H2QTvlVZuzck+MDIGN2bG
lwDsTfda+vKa+cfv7ZE/zz4EHFEcErKMKtZa8c/O2i4e8IBpnmnFhCBX2R1WyzZj
U5ZNSbuG8ScC3h8UF4LNW0Xa8BfuYtCg3dcP1+pGk5Dtk7MBoTmMKkeau1aC++Do
HbjE6ZLl0YC05+inaSkyq4LIDDv/I1tGOt2NUUt/Jm3kekJxj2vZ0HV27hY5ovhq
w1xeMx4drgL0FqOb0H2SdsJMMDWy511iQnCBP7Aouyr8hpDCvRGxOVcwO1EPySUK
klxn789n4fCa6LXk9mRKgmpJZSMuPDtZpapctp3Xl/KCTNb5+TI1XXl5w7KVD9Gw
Isa7BXNX8SOjif0AOFfE3sWggkHbsC9Z1B8oUcXcv/V9zs/knlDrf8ZypwX7ZzhU
ZfYfQXpXhg2xsvHfw7mXK0Fwdu3N4qyZyRbGCUsHzjMfI0+2UIr5DVLSL9jePIQP
5obyBlxsUvWY5A+GB2hcH0Pabv8rtbJ0HY8Z/qmX2Ar2z9kBFMWGnhg+dzn7+zyM
OLHkjFFie5SCi+gYiw1XMooIlKVWJ4w9E/pPDyP35Sf3kKA8qE9Qlf9hbtJoyutO
hZLKLeookUtQ8g2i5YOVfFl18GadslqzGV+U2qzg0BE4Fld+6Z3TUswJfuAwUsQ1
hlvQZ9VCQGf+APcgxKlvOmUcvsc0DYyZZ8uheDBJmQCQUBujI56w5szrf3NPcwU4
EUFCaLWYIWbS4tnWIhd8OXmaZBS8CuI9cDm5ylp6Zv9W1JaYqbsGW1HSgI1Xd8d6
qNwaGP7gobWHzEsb0hRpzun/4WEDjby+nN/YMBlD5kCj7hlZxYMIAU2bm+GANGat
cJW2GknaXYl9QbFNbh2fL1h71QI1XC9UNiWD+AGuCvc5faseNQq/MduozsWuH0q3
ObqrZMEpyp8wa4clZcgVtuj3ma/MxRyXEVkRZh9f2lIDwKdQfJ5hNNRG9huhm1K1
KHrQ4O2lWREV14PLWVjGN31KsP1mTc8/qiOPgGt2YLfwv/RRRuPpkMsqmpClB1hH
Pz+r5AL3pR0WTwB+xytb6XI8Fu+04/9mwwJ0gF0o3VaGSTPgSAVg9TLmOv830u54
e5MyH5VDxt3chj7Xq5EOTlg/PrjaHMLXrQ3O5P8HDhUOyg1ghdDgj+qf3U/p7tXP
Xqz5QRPAbl0GVB7s7nXsZK5FUddGc7ANPERNoYoqXRC/OLlbzO6IcAoUEGGY4XMh
IQQc4LEj5TEtbw8Jxz+eiaHG/K60YF/GMV8NIECBHjLOgzauM2qxXX3mU3m9RTCY
E+RNMtsr9SMd9hUz5kLJTskSoICQFA+0OiHMEDJ7aka75yJdLZcleqjZGbqvq0Eg
ZliNe+QQ5lBVlJbohE94teSKzzhrbtg0PX0mDEnVCT4lgpd6p71hWuI6kmFo+IyK
N9zZOnwOF0Of/xWzhZljtt9BSnM0FWnxIGYFRW5MHsTUPKVr8t1DtvanSxXXf+zx
bN6yfYMdulywnvDSdzlOW9ZWW8ofw05M2K4apZ59d7Xlc0lv+2pR7hcNmCnmVzwx
cQ8GMLSsUKBbQDIlMeE7CJKu40pCZBxfqbqLGhUKZFYzArUERTYRc6paPy0FuzQU
eL/LOBhB8yQSK4y5Ho+DDO2iFjfGyYwYf/AbShh5wNcYxg/YDOORDWcpqj61IgER
3Gz4V86zNRrmy+psQFLEQqHz2sF9rsF8W2JAMNqU3p6Wg0ZKbeMn7berpqMlDpVw
271NX1+l1qTGB3uBYI5/Ig71K2xZzzYASXTCHKfxMRrBoCt/YupQUTOok+0pRxXs
x0zZoXK8uv5+UXuCfqnvos4y7xKpuN5q50mu+weLNTZzzwqI/zwDmqQDZkne7jcU
++rjzOsfe0mHd5vhoSUIBUOvYoEXOsIijEa56iwrjCCrU6wPZFIjc1SeeslEP+i5
P1he4AcfPJAntSKqEQN+5jzr/m7uMRV1M0/maR6E/cQvGY2WURyjqSXuKltdw2Li
Wfi7JfrqGKQXCqgpctr0B+keWVhi9gFEzkUo/Nqe6zWE4KQlUUm2RL+P1HfGhK8g
G1NtkhvbC/MfwR/x/HQo09QglWm6YB3qbXioobQ0lPDq//3W2hh8uQLCTJv59WJJ
VnJ7PLIWGQLdpxOsD5aWY2UeOlPWLb+VIsvMVkQvqdEyE6JvLJhsv3EpSOnFDkId
/3tuHGgw44f2opnK1WWm7p+tzoUAOtZFnTbjSKZusYG/iIppEQW8KDvcPpjDbMIu
Y8gvSQX+yyV78IAWxLMV/5Lg6PHYywDVgvTUJakUb3ZJbwUc1RgftxzP3uByTIQI
dqYsbtkllv2tD/Zx/WzJ4s79poNc+BCVpwGWJ7bG5VO75GtS6+n7fREvYKqDCrNe
wh+ZhS8RbvgI/T01z0gimRp75XWQ1uzrmxRqbIXeq95tyCRgNmRMEKwbIr8mqzw5
wQYsqy/UdfRmGFArfWo6A3wijmKr4R70OKAzeqWqr0qhRZCaRzX5cgTwQEpv+HBs
j8DgxjjdgwxjVahd+y0uU05NZ+0v+Njj/rE/Qrizmp0jRejeHiaBQn8n2WhtJEmQ
d1FMtCDzT5oc27IxDDfhhXPnixss/uSirsRbpZN4xlTvd+/+4vSYC/h8wSwpcVZj
DC3sCU6jgtZ3ejHx2DgQGWdj3gcNB/d6fa5JsBhFitCLO5PKP1btOSP9sYDur/s7
xk3F/a3ByJ4YvQ1wdFRFnq4YLzUw5S3dI75FNYCdPe7EB0BbSKOprm7KCtv0xjeX
lBFUig5QSSA2OWuHPKzn0uszjxCEQy4WMwVRdm2q/9JBItKDLQ4boTwHr0Q6A95p
CBS5QAn9Lh3arX7GGfaSs8JbgzlyRL1fgtd/6QfPvmdUxERcmFb6Emgf62/TXV6K
6xev+lr9l5nqK2Y0Fb7Fl7lM0vXJGRnlcs+uhgu7wq9+v7ZMApINSLtD6dJvpn6Y
vy2kuX6mmlgbyOuz3SGYoXDb76AluE3fBbuyoxGTqttYqS2UuOXpaXmQ/JSV7PEq
9+nNOwGDCblKPKtOhLRv7dFHFO9MOQ9JL2J6i5YncM8I8TZIkPLEKJFvL1VpayzD
rUNf9IEQbmgGdpWHHwLv9q+r83hR8YdnBkXdur0MswqFgrcg1smSdraKWCjcCBbG
sOp0rI5Nf6oDYHpP93NjxTGFxWIZAeYyxQDAV2W1KmqW+5dXb+GkcBRA0Gqj1j/K
5HMeBr+ywgbz4iW1O9qqVdF0dtMxrVk+sdQkjj0msIo9U9lfvCJf6gLj1YGNXywt
H8VefumB+g6XUw7PeT39XQr8FUE6z+C41fCaD2N38g1yam5PwK4lIytd2jgqhZAu
8Vod+me+XPMoU6o1YJRdIEVbFFWEYoqMkhsOvvT5YghCYaCpqbhmULsW5/gUQLu3
FoDHka99RT1SpGHRO76TCBIJhshLQTZaHUA4ZNLHQx8K4MUREiNXARRQaaXSMOT7
JO5I7qb8qH5XL1TfI2HDbRZmsSkTMqiy7P6CsN3j/d6XeKqtGumTdmO3BxvPvN/q
iD44IeArPtfHoEM0jJ5oSregUVj946KSZoVO1iem1H664ALux9IAbMpMIe4l9AcF
URVQT0z81lqcU/H1sZEb9t6DJj2rhae3YBNsC/SHS1hGama2DT6PkBmZKEhZTNrv
unZeXu46dF8W5pdX/zuNAGmT/EmkY5swLXY2EeAkQUpU1zc7qWQW8DW1QUyVHjoD
13EnNIjto21E5ij6cqnEDOdRUkzcdUR8WW+kkI1EkJdfqECHWrdp0cwThVI0Vhu1
o4EhE9coUvdjhlP1oGRwLjkICuH/P0WWt2lK6SCdwoJq1AFf4hdK1RWLmXZCCQa1
22FKp+pbm4ZwtSKXim9I+gjxJ7TX7AfEJHMaT6HYOrY3lc5rVz1WAimR1VP6+Jc8
b2lqFNi9tE5StqTP2UhvfMeWy5AVwT50asTe2S4xc67UUJ57yka67Gbrwiu+3GJb
39MHncoRvLRBGQfYXAJAamdhHdFtA4y81mxb2x3KmVCkooirqd6Q1LGCx1eLvZ7T
bC1HZOXRyDILk9iO7AYK2FjrtWxz0VISJyx7gzrsTav9vS5NqRtxDRSfPqFVWJLO
B4LvX6eBv0SkQR+c1mz4vCd8WAoNvACZNEdQk7OD8hqXK5cyLe8QZUEyyAcfrg0r
j8FgZeMU06KeululA1h1XjR2ugicoLv/t/ne9VfO4Jm9XnpEMWsPGU5+Go6TpjeD
2uqmVWGeuCf6vvTgFfGNoftCbvEpNH5RGefnrZc6VXw0ShDoM+4tPu5xdiCNXnXE
IBrdgXk3lXo50/gHPNJgBAa2bP/AkGD/avksdorMehHCgNK7R92sLq59Cq6f8eCE
5XkikQUlKdzQ88d06PoUgVwm2Z80laELmy4hdNkv1R15q9qlaU0C9CNIKN/GwYNF
hIWT87rw+oN7Usk0l0pU/N9q3NnKssSWHSLXRDbwN2ss2vk8nef66AFlUHv3Bwe8
MeMXlKk/1ivWJrCmUpRIBw666XKpvrI2+O/7W+xScNXgJAVAXP72PWnCIV1fdDpf
0KTIoL6/myF3FEwYT/D1idvx4H1ueSx2KyQQccPyezH56tqSwrSgTV0ezisK1Czv
2J1sx3+zoVWPa2uXldHxEXSrp85rcVZvdKQriVwxm1FpsjUxJduFpfmh+Nr7++IB
PHlejIP8ENAE4PwontMz2Pjv/7TV2a/pSHJG4c2e/4WWZz9OTaYwWnubHlBxyTeT
CkzZ4de5QQzTTYloJGdK15bHhWzoaM6VU3R0Trtn3AWNZQE8dLkDyXhHxvWJ7kxB
gM0OMorJpwwmW6DCxsNAcD2y/mXASPsFVABZUXR91rQGFwzIa6F85dhnbmM31qqG
PW1wEziSPjlTRLNQPrJTZ4QpizmtMSJJnABlGd3qMYgP31sTdhdxoEs9e7bOcVK7
TI99iZTd/h6vJW77fg3XtrThfdgK58tgy1m92zVCHg57f7zAYnuKDk74c4IFnQTV
xE17xUGsn/reOJziV441gOHWJOsVsGhkTtuvUtS217XxCXkYFw1NVBVJGIT3dG0O
rjJUuV/wk9q/O6eDweoxgoK2fLXPNSj5POMyQFjIB7pB/zxKByUBy9sLEXEcYneQ
GHonz4jqDlk5ZtnSpOKCPngXZ12i9mqTExYEeWeOFDc94eOhF3qJ14/upDQa1uPo
cXpKO4OE4oKC777w90G9ubY0B4+JGncWKROiCgL5GFDtgAiuc2u7xOqBtxhRS6oP
g4ePyj6gg1iLwSPsQS4RydIkEr25f+NUBfAyCIc9PlPq2NKr7ca2S+3/A9cU/o65
GXUgIWokfSmnR63jlsEoEQLuaxcWVeAHl1qHYsTyifgWrEJ5K514hlfTDj1V6JnI
uF5GugK4KeGY0pe/5hVMJuTL5f9kZDVDjq6m4E4DqQgdhWwDk6f93VrnDhV/Ol44
VD4430NCPA+7Ko6SD9lDpNkM40t8rot20NDnrNVCRfrLpsKqX6BE/5cv4zuZyxek
0kjwzNQbANHTD54cOeoGI0siHSyBXlSVXOILI4t5A2gEgYO+wsFofMn4yC3CYxKO
lzKcTTb5V0Rl5xmd6q8fZvPdWaVDlIc+hCuUcMnJRJBbjrgFQHhFQoEgz0k4sIg7
vKicKuymz2n4BQ69tFVsR+b5IRzRvEhWx4lUeQMtaPfU1iipulXDdxj0ZX4DGe69
j4h1w19/XX/9FTEMDXzb/hNA3Fbqn6VoXYkNw/ZwbPvS55egCPOaoq9wBCTRmKeW
EaXgUlBP3Qj5m5zjLaFNCUlGN9so269l2bnAeZZ2+N+I5db1ZV4HGEll3Ogenpjv
Wwf3KXDTEJkOZ7JYPwU7+5E7NS0R+Gwz3n0a6G7M+1/decVzGgD7H8VSI422SQ46
Wempx1Xfxnv/yPZajJj5SJyWINr1Hwfgt2DvJ/ooO5XoKF25J8OAPj31342gJVvL
udHsQlY4q7WxeZI/HDO0F71ADID9Y8kv7OWO43ZpqgLUeZS0o2Hyccx7Cedj/riS
dvrfMPZAEIxe/FYo69eYibACOU55SmtC2sHtFyo0U5YGSkDlx2+taEEUEjBjg0gs
XKyL/vBOQXqdK7LvLAtvOR5YiXO1dBj9kQILCvtuhI2nyOIW94D5z8maDTp28Qsa
Tm1Gytrn/YWND5C7zLrMkEIGsM21rNpUukRsmhqhv8WhsI9wrF2fNcBZcV8SCyDp
gLicrAlqUdD7o0h7Esi9ZxRM96zAdWBVVnEzOQMjOHtdcqhnct6PA0LtBufpMXCo
ZsP9AiR/NbjQ0dQCFXMUj/RB2tO/0Pnmc/LW4MW4QusH2B8tCkVMoXjeJhirpGY1
IX0TYn3CY0wU/BBasLhdoJaUpvmP529ztyhozncJFjFwVUnMx1dMXdpEXtUubuWr
oRXsQvhJB3GrGvtvs2yOM+WB3wdlky/roezwV0+5Hrg2yXFy6c6IVyrN1G8zThHc
Lq7C5ElqrHtvZpoXeEmMVA9HcOdZVaOlLmblER+8Lj+m9kvq4Py4ruuJyQ9AdntH
A2+v6kf3/k7UBBn1DPe2DIUeXTmWkn8SXG5f0yra88a6JCZ8CtQftrqNMfO52QPG
GSHLurn91Rho0XH500niU8V3yNI5X6bWhyK++M11KzjM6C4QIYx/ilXNIPrpt+BE
W6NDNPfGaHqbpsj+iNYXNFTkulOaCAkcom0Q+5WqKB/w48Xg6UWBptQJd93R8WDH
blSVKQU/RKni/j9KmO1VdFiTdhY530eBVmxN1X9BFyuuHlUnKlXYbMAAs0TybUi6
alqxc/pZhg40esm5FOInXNRsowGD4zphqHkK3tZHSeoGBHjfNfVT/+LU/toBxatw
P7GR51CLwRCL9+5o4lL/hlfDB3wCULB04lAsqnm7hWNL/jubJ8fn6dmMM/KCf6L1
58h5rZxp3nxh4URVcpyBZXnQ/fyYwW2qY0JVtJF5fzu0V1Lf2xLslISvd9VmbPMf
w4t1attPIoeaKTN8hU6rIpiFPIdR1OqDpFP20TmfA+Dqazz0kWMjCPCm8FztOB5r
1O1UPkYK6sgNqSHYF2cfqJnRQBE8uB4s0WFcOqUtB9FDpiT4dpKJ/JTj5E+JKYQl
6xcnaI0ujpu7ZahaKQvyBQANfhStfbygNnoeNgXLEt3UQ7Ig1Q+7X9q6Ixd5HrXe
r4C8/B5vQ3r6AHUUEWvd8MPuWEHQ9FmWNNEQKWY6TU+PApA2LvZy/2M892xsAGT1
iz7bnX4GCk0tbVz1R/7P6Q91kcjydP0rcWXjjCeRWUf3c2aqgsQKJZFP3rbSKcW2
OK05bBL1q5JlEYRarOHq85fPLsI4Q5d+uRyxIV43iY7pKzff5SD8paXjSXeEQQIU
LhUuDqnF30ykge75U9dfxQ7XmG3oB3Pb0P8s8pmelHotx7pxpNzK3SJaX3DlMiMn
qPlpAq74JBaUQWGGjj7i2cV3bwnx/q8Jz4BN4vR3x5f+Hx0fNLKpIKK2lBex3EKD
Uz702AZ1KrFEfkAuxcs/dqRj/A94LhLACzmACJcVxKmNnHOCM31anIXpWgmEecET
WIsTGdv4kfzMIYOyWRzNzzm10IpN27F7PbIz8Nm2q3q/d88td5n1B+PlJO6/cG5p
JQxBBkWXM170E16B1h97jDDSjOrY3hrZdifRCYhD9EGcWf8h+VmyZ6c9le4Vpq7U
NkjG0CtBlLrmYPkYUR94WdsS+QX94d268UJRJeLDTtnTQXz3ecwjjHnlQLz//3pZ
WLfKuxPt6OMq93Xue6670PLVcTW5MW7mBQD3/ndR4l3KoAGNFabcmm76sJZVvyqN
7wjoYYKN1mxtx27xu5sMA90x6S9ZnjMWxfW4NkpbpC72HPTaiu/AkrpcmPPpXNXa
V8qjU9ui7Q1jkLAOj4vvLQ3mEElMlcFt1zX6IhZOOf7kJJ2WTWRyWW8mceBwuIic
YEJIvPrCVnf392BKt0j5oP9Ez0X5/RGBVHY5G3NAwSFgMIk/yrgpTSQ5UO+zN86W
EtWuyP9wfX0gRGjfo8BCT4ccl0mIGnBWGqZk+oJ9/+IN8WE9+g2N/FrDdRK2frm3
4SKCQkODASH1arHVPKZl1ncjqhCj+X7wyuwjT8LWbAnPUS/0zL7U14z+UUrHlSJN
2QU/0vQX/w2kklF2hwbWtKDc93WKAOWrPpDeYhwsGdgRlk/DU12kJHX9HzH4CJjU
rHieNCX7UQyKHxBXYQHtiHm1Z2WCvbjLoXbDRbyCjI/+a8/gglsJ763NJ066ldyi
dMa4U1BRLH8u6+60zST1Rb8N4Jw59+TiinSw+hpVKp6PCPABjeI/Dyv4jBMIkeHk
9YB+oFaooutwecUM2XMEyBBTi++OAbO9AWpYl+EfmhuUCHS6p9PHmrahQd7tBVmy
pYrHjtQ/T18Qtj1xmGz89ZCJfp/PZ4G8B5yv9SFURUoHRpxLrVWMCDuraHXVPFVJ
nnPYo2My1AImaMqKxPuftTgtSQhMGd188cVkDzmmOTmXJb1pF8+FKbzIGVaYX07e
k5YZ6dIIRdFOiuHQzuUkZTxkIC8rPhV/085FOoYRTaNf27HcLBDx8zpMhvum8VCI
htrSUnJy0Rxk07wMCzu3bpLC3MrUN99Meo5kwErYXRT+RqVBty7CkL/cPlkNeONs
UprxCxqM85AkUOfOofrHsNFRpnWPMsUU8fB7gyBscZZnrtzvEUjND0ETUIx2AlCz
HDFCRx8nd3EBLXbe7iAp0THKcfjW2WLl5fp/d86XwgSSxi6X4ZXdyk8stjDVbZsn
Dgk+K+Tt0rQmz24sR3Eo0vVEJR5paJsn9qdnhYadw+/7+DNpXtJU1jxO0CuvOQZa
Z07VvLF6SWxcjfUbLVxWw79pXMCSSWm8HQXxDq2lQLLn0cwDBX01CoOvwAOU9dLE
rq7UuxWwYqLN3zx48vGLFygnsrxlqsWLlosXrXWDLNqwxIBHcU4Sk0ZHAMYa2N1V
BeESU+brp5c4xVdsUW1urYLkCCCkAXNwP2issY+/rz04GoZcPRTesRM1Cj2KgIod
5QYVBQjKJWZ9HSJhGUFIPXJkSj8Uo2R0TdtSAgBzTcKK67w0xGk9XTXsw77qChfJ
Uqw+Dc11qVtNHEoLvl5oN5+VDHVa6mLv7d6yChfRxNzmDypD7dyfVKNx009VIO0H
JfFnzj3ZLuoOuQaEU0qquxplylZcj6xTVDdyqgVVj7fZGXWyPa20msNEIu0XJ7/F
5zfdUJASnzLlTLHUiekY0IJhyOfz5BppInnjdCbk6NG7KLIwUstvHwx1DGx/FYNS
LfQRj4MvHkh0uhFrU2iGydxTirBoEgNUL41z8LFcheIu9v1GMAGmJcVRk972NbtJ
LryT/Ipnn2Jslmkx/rxn7lLx9/XvSK0WANxRwPlZzq7xv1ZrB+tqbOS4nJsYdaVN
Fbv56CPXkRke0KSuoYEAFDUavfUpc+6wC4Snsy5S48tFIYxG1RsHhH0apB11PJsa
Dc8yIHTXp0aMCwAhgPfEA/9LhMVRqiVZm7uaIS9KnaUF8fiDzEPTip5aOQJsMTpX
ehRxKFbPv/1XDn31BJ0vYNYH3Ei72Tr009Wy1rUOfc8TxJfnEUiuYFVonPgs+rtA
JxBxSy9gIq2fJMNbOMgA+8/JgIlqUARgdEmWPNFLXqB1jvrJKZJe48XKz8QvS62q
k67AS3CA1ac4wcvCCSd3m4kk83AW6viIsvWqTC2K9AYVFBDwXXjtEz3EQj8k1zxd
TGFYhzQmWZYm8eV/yjoigEYSKCIdtHr2TSg4WFOlyXTyc7BOY/d71py77wjJmDdE
rYLAR4ZWA3ftKYF2Uy39579NXjE1lZyJanqjuH8S/zk3lXTNJGpBLn9Ow7V1jIRA
RFDepuOZz2nR/+Y36n6GzxhQCt1bycaQagghxaknAc29dNZ/yO3PnJGIjoXEadIK
9gNrqg8vWPJv2hbfU53LiQt99b1cOmwK168oC0sbpW/+00lZ3Xm70jsbz93sGOrh
zOUkwujpCCv3MU4PbiPZ2h70K6PMOrrRxdDB2VGM0q3fw/ebcfIsyfsuOxb45nWi
OVTszDwvn+E/id2YEHrPfWmMhfnNLAdaDOjrpQk43m2TQgbSjdjc6pooTFAeFhvC
1YuiVBOcuXYCWGu8sV9Vwr53X/HZShpT648sRtuHcEujj+TH2Kr2AeTVXZ1QlAUC
E8Omb+DKIgjLrk9gRQHKhVQzj7P394okpMlpaq1ZfhLC8P1NkK0M+KZSvMSmk487
ooZUMElEjDTeeHPQmuJHotTNEVBbz29lW8qfjAX0UrqVaRYj1fy9F0UF8alvOwiD
HQC/aHe2R3ZZj30q7N4elayNRPEV2qwzeKjTFJCf6bGupuM+8c426K/iw5dD1w0j
hn1UxIveLoA7MrWoHh9VrI3XQ+oRP1/nAsCI1TCIx28Ndv8WH60dI1DACia7zgy5
q31/OQE2CUmwkvDXSeqw+cSmZjUiUtQZC+1SvU3w4fZh/lUFBC3ba8qg6DT0W8Z/
l22cQe6/zS+idrcjqPWRt2gPBmGSnoETYE8HXPzfWofvn+199TEWJAF0UWSYqesz
RpTYd5ym3XXi+b/W5khSrC1eg3DT38zxAPAofHjqNB7SxF2stqR6bfHlU63GC1+l
coD0ZNm35dnAEiINdUG1R7XnUKDkDx3SatZb4JshNIQTya8BUQomkD9Zkuj49iNG
q9CvG5vwqQUbxTzPY6ebigUTAX//uiqR1gMAY7aS9lchmFLXYef6oYMGit5YqVy0
D513NlPEWF6fGrNiwpJpPXKwMXO5EfSrUnHM6sLaGv+EO2njqADYckIp5LQLCVtu
MhchmQPw1xicgLyg67kJ3OTECOKAEXV/xj0DIzRSKEsCGp3du8FfeDYbow6Gdr96
4hiIgkMfzJXQImm43rZYhJNQrzX/LP35qYUdF0kgxZs6Ww1T13az+cwmfZjd2MgX
ixRCG+w7BaBsZ7Uk/4PlLGMaEwi5hqlKYbrtIlfBh7AJoF1d5WeWy+0+GjmLI/GW
nm73QLpY0P7ezywv2jSNzpw667wQkv+R6NEfcG40ygMGYnLy4xk9LgrFtdKJbGBv
U/TGIxV5S0q8noy/X6MAPxEWdsV4WPLpn/axUjnUfwYv6i3wTpXGjrVhmZOa8BQ2
FVkuMnsuzyLCughoaWlq4ovgv8SZahu7CyF06ld9+1dO1SIRv4VuiQJsx7hF70Z6
yNDryd5F4KZtAZHjBx3iSE+BWVSnirlVWrGI2M5YI38HuNRaGouzztT+qMbyyycl
JW3oyOttwg1+FeSfRNOEJH8lynwoN6T9PGdkQqUF8Wv/KmboS1fPhrTD+YeLR8+X
HPASAwr3lq7oa/4OemJYYu/RZWNSRnsYCkZIjiDHsLtWFGBVRr4LswsKr8521Dwg
wzePWQDaSFKrauSW1YgQb8nB4Gg8iLz/JQw00xl6qceHKO7F8tjNTIMCuZS2NfM/
vtG/VnactpdsauaceQJLZpLDqj5hOk5iQZseEgnsWqAkMnHXALG45QR2fQ9FDArE
re1nPS/YvgDzYvuCS1l6aU/e0hSrLRNUhJOzzLfVgUU1Ye25r4iuOgnG16NNwUCP
mf2MbkAjt5qXC8vezJzhfwRZcQ666qbvHOpYzOMkw0SvQzqceqjPnRGhLCkvXZHh
I0sNvbIPxd/nBgPjc6vSxZsE3SoWkLqqJZcnyO+fN9kC0Q/NOTBSP+9UuxzVmWX/
x9Al8HiaNrcuYKKkIz5s1tSf052v15h6J7wT13r5jutb1yutK08j++svaIWrQLjW
qJhFWdA0sLT87fkgLxhGjJTh1G8+S+DBgYFqm6yhpdhIRXmc2Qn7F3N5zxlTe66Z
0eGpuOvOzmoWcjVpo1ywdYs/Yl7ZcvM8yAeSbqKkM1oRFr5lSnlMbOwSHQJa6Z0C
501M7boBsnPZYeETFpdWYVEo28LFkKuyNtJcfGqBQfTduVnBbckNhqXsu/gQU3gj
py38xMR5g+uMRxwSI3rAUozkIis9dBwEs2EMm9ym7ozwdsmoaSkU6l+f6SrR6q8W
6o495mNreTT9hzrUCjnx/JWl/IW/K3WifVtXo6imu8MDT5CRu1DaDKcvbxpx67j7
FQzCMhohFsPY3CnB2OvEjdMz2xyEJwaeh5fGfo2LALUSHfpE/1b+tkm1v9/6U6St
IkFEItJj+ov+N+D3gzMwY5qEkwMafITSAn0qb3klmK3ioIVNZvYKkzXZkP1zEGAH
SyPeAwWa3cNBKMkyx8f3CK2kpEENiDmoWMc9n9jBSZGsUhVsIiEcgpexTb9XxBZi
AAe677mtOdExiCVM71mRYE/M9P7KwCikHwqxE30B9vCldRzy9NGZrJzLGSjDGukZ
6mGhTtbyGYAa4QAU591jnKuIfbVhLD/orwtjH4JRJMJ/xYwSTR9MT5dLizHKUxkB
XMpfpl+NFE+m4qtVE04wZPvSOxS09cFpGKUO9aZwU/FuzLM2NvnSFin4rumQG96F
CSEqU46rn2BIQ9N2SAxR2L3H2K0V/LS1sXCqWFUCckDrY9+5/JjqBAIeHo0hSMpY
WOt8Gb4WlA5EwHJmlF5VbGg1mcOFaCU7QQdT6luSDV3niw1FRwGWVQZOO9Ilzwmi
QsdTnqZfbXlYFh0vvLsUDf3tSQs1h6YpZlupNoWe+WCWIIZW8gdnJt07/i3MM9RX
VGXdBvV0w9w/uRFN2QhJkqXo5o5aSiqEYu9pefSAxtTjUq2OGEWy7vQ4HD0rxeoU
kA9QFWgdlXDK0BZ+cueoWMr+RPvd8qq/L4/pP3KLtZyCW0/NTAs5n0DjOASg6UPK
fJJrcB+VXiXUXz6BEqc44jXsPi4DZ7OxKCB9TFa9xxN6oVDynDRWYDIudoeIiVr5
A13XQlFKAl/eP6SQ9XsOLNl92ZWbrDQdf+P1/gdbrak710kj83HDZ9vAZ3UNexrt
SKJ4wRj3ucyirRDKyQH68d3GkoVSBrj70kfw5xEeez1SzsEROBwZFAdfEj40aig6
7PB+tzd8XsRUkHjqkPgGJLtFj1qz/XwLmEKj06raazLWTo7kpqu8fxvKHB2RGK+z
HcO5oojrhOYuX+ZMj8ykNjmHjDHHzr3p0sfhMUcemKTDvGAXwEz+DkeIUnWkrgAP
3pFB0qgspBVaRTcQH4IMIkZmSEAKtKJ6CLuN9UVffLuF3UmC6r1VG08cAqCl5NoX
82wJWUWu5SSODrfgGs5ZCTfROvrOoLNjfBnfgE8k3YrvuVPbdVmflCjxlVJHiYsM
03nPeZuc9v8bNdYJQp29bhjU6Ih0uBfP2vs3RWzEv9ZyDYnRU2LXnUXhFUXMpYxp
wCZ+8eTcnLxpfyN/D80vWeyrYWBHvKrdrVJv6wgp7CX7fIJH6grIHytgqz0pKtXv
QXWh1UW7LvlszvrBv0qoyqRrMlt+qxbaznD7LjiGBkdSWmI0JRTld91KOPU6b+sf
G6i5CG8GP7qsaJn8Ae1z5GreBv4L0mfs+8blWwaVXHeKTjNI2gZhBONwTXD+OPsH
50NSH5AKAgfXsISJ/igPh0XlgC0jbbxj0bhJ2BWVAu8+4yKfwGsmqL8YnKFWK5lG
7kS9mjLU1zO82EQH8n5di+bm0s+Rpx7yOxR6l4OEb8LmJxorUNiTBzCsAB2jtO22
d+khyP/EJd19fjbh/U0rPv1p4k7xQHxAjuzwJ/eziw3UtiKd0D2FLX2vrmHqRRLu
e8ksaIR/I2nO3V2DC9TWgVetnWPz4swKUQ1W2xN//G1Us+OV7O2QkY+gTQ5kn6Is
AG14uwL3Az/t9ZTiVT20Ph2CHl6xfJBcsGSpSBm3gR8aanYNJGMZXlaENZU3pQ/e
XW9xvB6xtO6Y4rIH5kkFJAQtoaUbLxrUjxVU343ptH9AZlgVf2Cv8oGHBxSmam4q
Fv+a++OAl5IlH8Gz9ewY+UyJTLHC4W1vFCFHZ3XEQK1B9D6kVUpKJqpn7d6HMv3p
qdHcxpquMxx+IJ8jzq89DlbifCsq61Drm+PuQcw4Q6uLxwCrINQnW+ABhgJotPqE
qQJk6IwD6olQwsgR3CKi/u5Ki+spz9QF6qzOW6FazrXVHeNucTqQPFTzyL0nTuEZ
QH//nwSXZSdiLDzGPfOExs6Bdu08BrAV/yDUdZwu7b4Jc1EKmw5CxIiEIIbEaAGb
5Vx2xNVg6/hcjeKo/kk0pLbWF/RL+Qh2XygY669AKaH5Fo2rPeBOqEES0EIG4Rai
09DZZwDk4aEHaS2H6P5168oQrzz1eNeoRx66Qqjr28MftIcbzyG+CvGTwLr+l8fm
MOsReH5gzcnBM1jTIiZ8SaiYUty24fb+s+hae8T++FWA6l7rNB7e0wmH+E+AgkAK
PSMVbdPgria9SwLuFwaVSSqX3eVNYnkhOPVdbPs+4FHkzeoPKw6KBHyG/rGcO/wh
oLUjt4xq5x0bolqOCwmnVupxhkKP0o5ya7JN/9h/wvytbiG07ahaGCrsFI+bP0U2
j+tgnqTQKHp0G559dWvuxFB4InafIZINbb3d/7hDLeRr1LSqiOWO+WGo0vKR486A
nk9Dr9TapKOaLfIYv81enBC0iZ9vv47dtiCA+FwNYZU9XbP2EcENfJFy55VwQcEg
ARpLThApClcyUCXbXJrcxzFQe2Z0YTcmNvea3OKS+Q4Lh25z8C1DiPKhewylv0HQ
GpmAp2yicBXWS1612OMm/1heNSM1PN6uKo0WrTFMj/dwdAU6S+7+UJc9IF0njSU7
a6aGMuzl71s2DJ53zoM3wq+jQPLNZnXhRujL+2J6U1LlHoOlcKMNbJJpAQICQPR+
soXi7jLDbRL8m50ny55dOIxdzKUV2AlasACF4oY0IGeKVHum1M2z6Zcv6yv2LdNJ
ej5iuVMrvnv3WNeedpMP0npCraOJSv8xUKEqhtAy815Dchgm22iKgCm7CaUgK2iS
P7DOMKYrvcD+dKU3TcyRUpsL2jRXA+wgcKx1payysWFULQpeFVoCr5y14GKk1e85
S1plv5EjC4Nk2Y0dW312qTR5qb0EfuZTXqPSAmw1p3DtrZAaZR8v4vVFm27ZNmly
PbuTgUptgFIhmv84VQhLPjuqnnmPV2YoHiIO2x+yv+UowAZuexMiBJZ7vO9Gtwy8
DbmzMKmm88AacSqZTPSRHnDr6uXd29tsSDBvQEsee7404gnQYPHSVJFFY/zh77kh
JIYPtk5929ypsYguxMh7++9byCT3KmPsKPI32GpsU1lTnZ/c/hVSUz2l9IJ826Ef
pHFAVQppa5AnU/1BSiesh85+Cc2cwfKHsRKfwObwubgbwzEe2xLv5e1a+HRPNCYn
Xkq/6oEJjEq4Wt5z5qmeVRFjSboi5re1qx49wPuIHp5c0HgrT+9sphsf36jYgxdU
Jr8wgK9oK3Xl+oGYmEFpygDUHb01FytYO1uP5PBBtn20RN3ZoUyFY6IE/Rhbc8fG
4/UVJcdkl5Je+JESLQlEoIXtXqIPKoiBDUKGnvDIouiF37cgqXjeNuRBHdV0fIu5
Cd8eqjLte3udd26UZlWtVg75GG/emkhI1zlnC8Ndlf0QYqJr8RcMmGFnbndCMR+1
m/4lzTy2d3gLJ3bASiD4SJrMGjip83Pkeh8PFQ+o2rStXBAkPgLp+rH2+86csKvo
DDf9cFPPcu2arldpdMcEFt4d/S2jzgoPJAI1T+tQVMZ81IlwG4yN/6skYBzRkQPu
04C3Y+b7fC9AmCwBYgO+Nqde7ul946hSS50hoVveRdzdxwW34FHKJ2ZMa3ZRf9Rd
QYEajNQniAPwCOzF+EKWQiAVUg3r1uDX4hhiTRuw/cf9wdTVhRu8AGU/JpWGoLLj
OvxuFbdQl63s1sTVYEKCsTQ4AaiEGeQMINwaWXmMfn0npSrL/lVS5tlmt2x2dLyk
ZnCUn7H0F0eYdN1T3SdrN8E21uQz/mXItJ5ByrLqjAxoNef6EYlUDNH4a0skyqbb
uVek4C9nNtygNErNHLczLtmQppvVvfn8oC+JAoi2YnNV4nClqF3S8D3uDiiI9v3y
FVAe0EFevwHdWdWpuhcC7ZAAbxNEvRum6wQsmOmvaJXhEqAzSpl6M2UAuHEcFVAe
JsacQK+R4SdhFkrKlkt7IV+gkC0kmEn9+RIBR6MqZWifnOIIo5jKYpp1Rq6AsEdG
G2Euw9utmNDUgLUnjeCtr6/zs3cTN6QTA3fJ3VdMFWqSp1zIzFWyRvTf7+LZx4qb
KS5lho0kHa25BENvypOLwZUaTK0IEYwXzzk22QPdXNT+byahc+HUo2Lvf10w7wvk
cs/TPfVeMM7mmIfDbaF7H7mw5ur2SNsoTKAdF8HENottoq06CfaZ7FQjDASpOtyU
HfUmetv0LCycTt4aij6hm20Sge2VfdET2oWtFACkhml6L9AM0+2GGGHneQxF7MY4
tfwah9YYytyM2sCehs+PElh6Hp0a1KR4sBiehyfdjApGxRrnK38wsfr/2i3Kfmn5
kny3ZznUzowIDjHhnYnXfUgy+ivqeysYyo+NGrNNP5qEIBWExuSq0KHlgguRdtfN
LKDNGbcYFTVC5Co/w2S3MCkPm1v5OXL7ro4vrvdaR75fKcpCgJGpTgkaXkjuIeZ1
MUR5B3QcqNzlR9SKcZTMAmLbF4F+RXUgOzLvmsarrZBR8TAnV/su3FklxHP/v79W
veWW3LAp2hajV2zcG5wqGti7H4qYAqWrW3L3S0VDfxX3p6VH08vEMgfXC8n8PM7U
413nLlQ46Nz8hnMuItGuKGYS07rGzFV5ZjrfXOZS//OXXq3dYyaVF2G43eB3YFPa
jd7UBs1CqikVZcmhTKTPDFMXyNvNliBtfFZCLrEH9XZNs4n1pGJ1Uloi43nIzT8H
06+MGemDOuFnLFKVHt0AaGXwx2YnBeTobumJV+CEFPx+JJ5AQ/+yAHFs7j4wU1a3
pnEmIhuPB17XhClyApgQVkJ+WIXpN8S1dpIfbqhNGalmTWV7/iOILHPsf5u8B1qX
+lfFD0fZF+YQkfm4hA89ayZ1gmEqMwLQjWkAMxUoO4g8cAbgM0fKDvq6ZLZuZf6s
kBHusBkFqqi+Nz1BSnKkAcJ17HMBcY4xfPhmLw5FHaNPuTi+UVTUfHsVOv76Gxsz
utV0Y+FU826JOoN2VThsug8fcLOVrwJmG4wlO66a0H7ao7qUazkQXcmOCeQb9Rkc
P+6N6Ie3lS7eC3Drz1ge3ysmwCbapCJx3tnVM8telGBBuZt8aoXjxGipIW6hwxZw
rTb9IaVBuHfww4OPOq+GjdZGk9Qv0audysGt5wEn4qhn3s1MqNOX0hcwcOqflV4A
KZeaGvJh+kmG7D4mAz4AcaeHUPaiihZI/lTha3tmMnVfhcK71YHvNT9AmLgUBF9G
Xl/kxPvhSEx1lsT2XcHVgFSCOMQXtg6kJXC+B3Z1rvmul7oOS5Z4+dWeloey2LVa
nPkuSDj+Y+KStOBPcWjYxekt4SbEK00IVlqaZirbb+n59Mz536/bDcoUa2krwh2w
9kHCD5NxaJBEojcjKVTsqzYdHLlL37NEk0IXz39Qo36w6LniSA8hGYnAQpUKubIm
mrvpfBi8SDAXBvihsQ9mU9d6t45WxnUnQMo28SQfHR7CE90KY0R0QdOcPQunea+O
AM/aPHJav0Yt10r83hC1DYwAIqXWt6Uhx7DzGsd6IQa42pP0MTdgYqSEYeymTxTX
l5luM0B6yeL1CN97Yn582T14DKSaRNOn7U7LMv1YVVP8/pE6gn6DfzlDULD2vo7T
K4cpzGa1+F7KCKT9z9aZazttOVzlpYXs2v/qAgeMFLTJty0CljovQBLR4aPuIceR
5JcGKha3eA97abDC0PHKLpOuv+8oJHsTmSTi4fBg3Ft3cXkJ30P4M3pn0/XuvaY9
aSl6Da7XyVMisrQOHVBXCariZwWxWOCLjliC6scqYIZ4rOnNte1mpAxHb11PJ0JE
QYWGEBOrN9uCNUKisjUxyvsmseDfWMZBcjW1cGWQHmtQlhg46yAhMko0AfbUPykp
niqf6gIoPbNqQig5388GSZqQig5/Hs68LEBjqE0wqp5eqZvfxdpJW5MfGuJBTSbx
rs5Mnl/egX6ig7MLIi7PzvxKvLbM78BNF7c5FgOtgGjRTwVPXS5nVh6wzqoqts/K
WbSK75X2CGVyamNR4GC9ToQR8NpqEFQDtT/dcSbzAB14wO0gRrSwTVXxmx3054sa
9ME7EmP5i9dYFYhNWmSRuStKgdoAQ3E2akzZqEAdG0G7C2CUUPTvK80EOqAtdS3n
Ho1Ts/9mW/6h2JodNupmFQWEd3UcTKpxfgK+XgjfqK65Or/CiqxfvPEGaam56PPR
v9E8wjFBfVsGPzFU5nycIeYHCZbFpCufg9lX4638Ca/wH1eYV9nxr1cHKSIUF4WW
n4oWOtZD6qbRm1OD2NQvau0NpuhNFbKShHnhxCbo5qalfRbNftLueNpQyeVvMXQc
cVCdGasWpl94lPsQpbbChHekCjyeY+6fDQMw8u9yF4ZPQKt64mXJYIOrJEgb2rwz
hLvhMhiFXNK9s2RCGc2TGaR05V8Vs8Mc26tgvuEba8Lxk0ENR/toDkN4QeYsvGMh
ZbTEj3XAVshq102XGij5UGnNgM0sieY4epFwnfaAiOeqiy/7wztFL75AJVRHTCSm
LZA8D1xj4RwAtUPFsrxbnAiMIqKv7FBrSLoAW4SCHf+TVrydaDfwE1aSblkLzKfK
OylcQoM3DrwTWyWYGHeOHbr8qVrBs8l569xrII47kiDYCLgpv6lpeZIJjlzGcxc1
FJG8Vt8GZUSFAtYXFsv5jscJG0bfw1qw7tqb5RUc8h0p1oKF4m1DVIZZ48czZIYM
TV5Gd1n70vk4NXxRp79SZXy2iTqT+oOC8+PFTVF/j8EQtGVMaL1BMH+7ZgSe6iCP
1uRlX+MdOaYGwWEFQp6nrr1eEWosvNsycUszxLKieV0s/jDv9e8pECHIRXy3Vs3P
OIxyXn41NBR2hBeikt/ye6w6GBnnZ/EPSV0UeEJdjclgTuCMRHLpYlwarfXz8pQH
jCtbSXy0my0VGCm9mbA39MHLm667aPj3Sgbcu2nudK3UNPLHnt36eJX51nLgB8JL
w5xSW1i03CKy2a1sIGHm7cO5y/U1gkVoS52ruxOlggVHdbr/9AFiZQ9hc0SX27uq
dthYu3YEW8yu8IS/z4tqNCUPho14ycfyKnqe5lWE/2jHBt+OD7AMdRw3+A85fHHZ
CdDKE78THJs5tfsamBwCwbBq+kUK9Mqa+1Hlh1+K+wIOUvYJhe9MjHjz2I49+Oil
geO3WCvlF7FQBwxRWD/2MW5af8D0utFqDEgZeFNb9ykvryffInsYU9/u2Ieq+/CS
D+OEPS/RslLb6tNsEotXDwAznYgiqfuCd6SaMsku5TNp3LNJG9Zne3BG9mPSwk3j
joJbiE861N6o40KnaMq1vRqtt1dBQ3qAjNpsTp3XwhO6gKg1bcffQZKfWpgzCkRp
kuZoNQbaPEMwe/ueD3EFTTAJ5kabkCsKPjOghg/ujLGaSkqEBoExFyutAeUGR8xv
wl8rU7boStVN3PAK8m75p9zOD5+B8O2Gv2RQ4foYiHCUc+Fe3XucJkfo0ZaFlIkJ
cicscqxIamHk/NGaakKlO7H7XJyQObZcPS9JRjKfe+ug853mvx8QCeyLg6lVCYjB
iyVsVBuDDX5McVwW7vv93r+c8lnMpr4VICVSvNja0YUXWF2NSqo8zLs5j/a6+FLb
WQtWXkjURiRFen5Fccm8zy1REezZLmKh7T5gisRCnpO41VB4kQiQ+yhXJdiDSK41
x64m8Py3SwB+luPA0pMqGK9cUDlaDPCep/Ybwj0mAYri/wd7yjpkc1E+WmfeXKhk
y45zFfVgf9uZFQkYDBvVVdmGp7DM03QAXGeSpLUkAu/+Uu2jmCpyKAB0ioUR5Uw4
ulu3sx/dDoI5AI4oC+Yt5XKfkcIWVFtBOoXNZ02okv+vZ8o8/4IFPsccfxbak1Rx
oCngOu/9/U2PCaeil73BM6wE/w8llktE0f8RShAsbqF52Aw+m2tmO6n1jvj0fxrg
nYpAKdtIEevdn7dtVCEwnk4ZWpo0fv2FhIEXcKZcKAnVbng16Oad4EC8bsy0fNxR
zEuPY/TveNwvAc3VKM8ZVFJXWGqlbNiJi1Ps4O4AtznNcvePOgX6rpTRiIpeVxF9
2pf7dNZENVg5wZufVEqnIieeFEMApOdEERSNCiueHqvz7PJAeODcF3CyFIWaQSbY
idjLGIun66luvrUG85EpTPhr5oZBTdp6hIQ+JKvZ4bIa/tGm3EGbbCxQvekZiWDb
320A79pXu2hC0gVobvM/1B5vHbL0NnF5heaxwVb6EmBXPjkyO1fAz5qf0sh6ojfd
1KqslGax+9ACyATPMHNM3gawbgxyd+BdC0w5s1MvHb0827RT5SCNAfSGhG46mTlx
m/gF+Gq++U+xaDIfmY1s5LorD4oAyWxIzJ9rJXxhe/HKYIUJvBTVnGWsgg6FOutz
MoD8wU29ARDrfnrUOmYw5cLd5nLn7ts7G407SGMTAlTRFONHnIiR1zvPKjhV59wx
86w35xKxE0hhad0OmIeb5KemQsV+z5zRtH1ewO5lxmyIXXLYDnlVfrW1MOnor0da
nEYgRpb1BnImwtQt7U7veCl0LeYVfdlOsTFKimRvhmZRKf4mOd+KYTw5PxROOjxO
n+zYGIZVq4eqWLKdZrqU2CdEiSXoVzuHv0Zgo+rorJUyRxEBaN7SSQIynp9UZbu6
cA2qcvO+ISz56uJw+UNlWJYRpeDv3YGL3vURUSSPeaktSiX9EsQlnejL9G8oQaOl
5tIMz+eP3oHgtV8mpj9YVnmNFi1t3FjEnNS7Q4kpyf7fsElVN19YO6X5KjRXY3Wx
hJbGiGBZHUZDmvNHnTI+zXQjKYjMiPJtHo0kuL8gTR+1+S7MkcmakMHWymRGlB25
yDdyFRwyZXMgzUD9CjJX5n8Xo5jPDdZSP2uVLGdLiX4VVt7cMXEbv0QJPrRHpPWy
A/A6HfGvvt7DuetbUQwxDbMjjGciK/KkKbTwmB4/k7qdi39o0X6P4lRyEko9h9d4
NUsdDnrewXTIp7ijrprFowPlx+PP9YEcoybOb0ULXK//QejEKpErQt3Dj5Yxs5gH
PnOgGwK1fLaGe7EsqxM63jiQ0BW46gho4wadYWXw5pwoT8WK5vK6Uxt/Pw5PEHWa
7n7SevZw6CJPDUZ4FrGO/g9Z78kxLxDVi9WBiBZY5EGk8gSOa/zsPSIy4iPDZED3
KscaV2/c6ZQwwnOXmbqxcKvTDhFryrSuBj03oQ4Kt6nxwkdbFuNQaERGnvB+9eXt
4b3HuxrAPe1MAxwRkhyAYPxSJ6OLNr8z4hDtJ4CTFNIdIdptCPdto8lyE25MEIiv
sP/T6VWmgWMaPXyU7IQdYXT4GWMH1bGXE896kJFa/wFxuES/PyM9FLT+SvweN26k
0/n30siGbfhzNo/jXyH+oMKMVzvsiGSz4b6ZSmGTbI9Fn1snY2MegyWQWJFTgxgc
4fI9s/8I4H2XMPipuQ4QLF8UqUTRJZIFq5a+T/yCgpnfdXV3fXPyuJ2Vsn+3Tp9r
W/hrLkxFYLZ/FJ5dUlRckn6L3cfOWe/TCVYwnofSLqEazQ+z6+MG583HmFcTc3Ku
pfshOOtZelv1fWPrEa0VCqkMXKgKaEViWcU1KNLIJE7RuyX0zYPuCz5yneKgWPTJ
NuHHfkPBLQhKz6Ulvnp51I9XeCSSf0PVf2EhJOHN1kdEnsGmEFYsVbRmO7PgpwyZ
Yvg3RJmzSgM5wPgMLzOQ2FIMSMiX2myxtDBA0VB8HpFpUxNwVNQksiE7F0+/iUrF
FyrkRnlg7yNYVBfqFEajqnw4zrShS4bfYEOeclPCcBR+D658E6gnZNE6CGCxGfBX
PS3iUGIuWYTFK9bQHXVOhMnO6MhNrH/Pb8lccEhldmBc9YctCveI+ni1M7kcrrS3
6D6rLyNiKoztlMn4JLMxd9pwdnNd0AmgOSKb2uvmI8z5U+LhWWN2iwSKVxu0IPvk
gACgvo0TYedIDkhxglaBINqo+s8wEua0u2u1lNeaAkyuI0BA2pUN5QlIY6Ec3VLc
wXkE6E4Lo5ZtvMOkRBL67U1oD4Fu5A0Ne+1K0m1GqZ4e7zV8HEcWtNE9WL9OVjgw
QXpw5GV7kO5kvKMFrRuFwMwvKnu4IPEWB7z0xiAxS7GMOiWOaLkUYyYwpCWlo3xX
dKj0cxwwhfjKKKbzxKhy0JHTdx47EOElph7nSonKOhai6A0L7da9PKgZgrechhP8
8Uck+9hLWgE7KemNU+6eAtqBQUETwnNTjUkOtRyE8yZPlujWIOKkYDndUXMESbuE
zfnk2JJQHPqJCju2yUa1KXNPQjUb/R3xeOUi0UkAH50h8BgRUOnyWyydtmN4HJ3w
1HkcQlkduud27iulr+f1OHh5UZBrQUAgJiW/LXT/Fe7tuBNavaKqwGz3DlmPkYfw
hhFxHKjpmq1EAFD1fJEIVjZfSFwjqB6BZnnZN7R8nQEvaVDb7QP+m5zb6SA8TuS8
R2QTa3zDjNGVxxe86x1ISpvRg0qyk5pItgiRnx8g6YimGPhhK9ECST0aB1JDHBB/
g1EuoKLsS6Nfd1zWzoAMGp1y2zuOwdFcPkyRmcAKDbGqydXIvSj2sMc5koOV4PVw
Isj/f1b0XdNPVOkRlocsMVXDkDqUmZOgCXY3/ftoF2XyavBLxfLQtQB8KHKrdlxW
a4aFC+GjCZZh0dS5ycxYt+y+Cknf0m0SzVYRQEXft67uB71VokktSvpnWro35XuJ
ga0JrQaTkQrdbOD+wcNw+rNEE3YSSrnXvNLkQ4BN85fXnyXwwzJt8KprqKoNStYV
z+EeMT7eWOdVYS4OtiHV2ZhA5It+irUFehVuI5O5h9Mqh2lcVlIKM3Xic7A5M0m+
6tRcm/lUqvEk7eEpefdZoKdrs5CWVvgZONUH6EulOyJYQVs3D5vTLFOrR8Bi5opV
4HkGfrdsdpzXQBOfWziNgZdim2ntRvFUeKA2ghFqUeuukMA8RhijOucO/KfD+JiB
wgQi1XYpwWI7CpFTGcpzOmLrr66Ph730++/AWrqk4k+I8jJ9uJG9y2VpcYTAifpM
97YE4NPYPuauc3Et1/cBC0AZ9IFQ9si80qWoYNiDiz68l5uicUZrMlQV0G5J/9vY
BQ2piv5YSxDSoyXir0TmaYJeOAwWujAo7jC9OrhtT+tNLO3chwZMRWFR5P6O6l1F
6RWmXVKpZ61KvdGFhJ1SMrv0IEHWnCyX54OqFPeyobwfhYjYA7dB20ERlQosfUrc
tD07/UgN0eKpDQE/2iCQmUOVTcq4qd4pNhPo9JLqxieCmjENYRQZCrKPte6gC0AN
LMaMYXtKsv6i0KVioQdoOJcAcEoRviAQ3ARMbgLU9QSLpRRxq80yhl+JhSw7+Ro8
qyAI7c7i1B0YlQIMrp6Lalw4ClNG3UDsXOJo4ZaQHPJRKeJQ/EilkxO7tlKnKKdS
EM5hmw5jMRgy2rFrlpizXuEvCra0/A/1uaQr8cmp+mP1jNNvzKTf9be+kuo//YM2
JM2MqMPQuaJOQ4g3MQtDtBQvjaP9fcWs+i9KygtHQSxIUWCbROrmc4mqufNF53FG
6uyp5AfrzCdgcpt3EfVfiSYCBv0SujrGEUQG96EhtwNdbX2KKQtJx0uv/pnV/M51
KFHon5FJo4SdrXuaB+6EmmVBypaV5btHLrHZEyhXE+ie/wTaP08FO7xJcT+3ZF20
rwbX0CzKOLzf6IyxgNtVJ5fakTUC3t4ve2EhKCOketcRpE666Zxy4yXJvFekiKrk
YuC54PCdXGaZG287Si5vleePYS4UkYSqEfKeuJFn7fifjbRLnfq4ROlC5b4VxBpN
UIqP6tT82icgE5D7ducFqyhFmjYUOiTIZaFc9vYgR6aAYU0HbL0KUEYyC6A5PhFg
Ccl9rr0MgGjnSpM7QSawzsVEK7wjVNvgAhPDzdm1ECdeXkkIVvdIkwiwRNCmGg5b
vz1M4V2eHlpkE389QcdJIg9h+bAsqdEpgsjsES/QlWl/a6g7vHzBPKW5LrL1xvv0
wHF2+tEb/1y4cG71iL634qgs4cdbja2h8ZXPm1/NinMPnrH9H30d6aK2Ak80RKeA
2n495QACLqwN+ClvielaiXLHYZfcpetZ7tcDgGLOjF+X2liHP+8l+6rtXkKtca9l
TQ4Vc57WIVrq58xOxWLgDDsMt7GxJzofq03GPgobNiN/UPayUiIv8TxjdrgyReIa
K0qDBOHJRKJN4xaJnZvEqTVZIxbGRytRAy2s1ak5KH2MS/3v3NVwbXPmvZ94fVXt
Z4Ws/1fyLpAvhHkdw3eyUNrThMXld8/5bdrFxC+SHEnCYXr7eRlVJujtCFEoyKlx
I8D8ZTM2ZeTVwkJmNdKvJceeiSXY9+0d0BupLqRk35cRSp5bH5dF7THBVPrcdzio
63KTrJpgryfXbylyW34XjsNgb/yYFTAwj2Ht75Au+kK26l3hcbXb6AfD3isAZhOg
q4uYRPKJ65bWwZUss0N4AyVM3KFILijTA9qOxzYiNqFnksT6bipiKQltr+k0abd1
uv6+wo1hLet5e5O/GfeJmi4ngMPv0RD5cdTHWNcrsFxORiQSISMiyOyLmhuNu+zW
qJ7Hv/r+qFLvijnZPXusNN+KtPvpka1OHa2GLYT5RZoXiaEI3rebdtqPsW4wICOd
hdF08vd9tS6lOpk+K6X4ynbYoVh6izQPp0dta0WiRg4dIpz6ma7Qe72ZfeQkrspr
Xxg6O9yR1PKgivLNW5GJWbXEAUkYxopYYqzKc4XxFqKy8GQN+nD3bXexkJ5Dt9M9
kH25frHeBgwGX725N4daYW9giIfIGYJESPmm7GzoACYF+VegNOSkrjk9nHc8CxSn
bH4+n//MuTw0xKYH0LQSZOg6YQhNinfOi8jjT8r31It9JRxmjHYuNgqnqHGMwC4+
NKzXRqXze/1Ucm+t+VVt0r9VNjq/IsqM32aAVZINXiiqF1R7AZYkMEYzCvHxnWBq
G0fCDzJUwW7cr26dx3k8PYn1RhHZ67jbygB04i/LZRzvaJmwu6wuupKfCOk+cR1f
LFu0UG0ietH/MbtJnd/rqmQEFWZbZV1figHlh7y5GmYvYgB/fx2Q6QMQjlzAw/Wp
Q3iq8LcowvUxnaeyiYzsOg25BugWRWwXZMy9y2jU1/DTzCHT0YCENhn8RP2GEqXC
eNNdQfjoWZHOMyaoicSsaLPWtNuow/UtbpOighAldSVJgqKWYWlsQJekj1nB/aHZ
4llNepMAhaoIOTduJ7pOrwHZr1VLRGfW5kvUuTaiOjV9EVq5wbthUnYjstZ/o9Rl
em9XD0jmMYll4wYx2sKxWd1rV5H5srxsFqLusopcVCHemJw5h9T9qlG3QDr+r0Eq
d3PRp8UvGGRSFBjMJD0D9AsDeEfldFyB2Rze4dIjxNsp55+izGwSxDuyohWwKJG2
4zVRYM2nhvn3vTn6LC1QIVZ35HA9GDTWezp5Dvs2WvPEKJFKZQ2ncKuXW4hg4ozW
Ec9CEJIJg/5DtTmBf785UQMv/vfJK/GpysPwHfv1jltZyE5USQCl72egG839ia+6
Jcd0RD/EaVMAqH5+MCdgFpFvk2C2quNl8lNo9ugv7vvyBY3k6oMtilVF1JTeqCwq
cgiJr495hhRhXgySSXPenHvN17poX2/Z/3PtBzqI2VHIlunycktyrNd5/Tpg251p
umZJH8sV0Csc/vbKNQ8L75QBhaV1UAjsYsXPBmYDm8n6LSngI/ZCi8+Ev/H9E1uI
6mjUju5J5oOqZEOYTYedM2SVmFUNIq+uyjpf6c85Ug+SCIvxacsL9QDD2XcEMsyU
MEpwk47C2vdVaNbtbMYPQf5nDztbs2XaCUzZ+SmOs5iYkOxDrYCaHVPbUGdic4XD
Y+Elp02P9ggJI2JWtzONoHjXZdg/082btzRkwD3B8QLKvhGUEgXpMBUu30I2++ys
32Me4Qen5sEDE8vZ9ljXiinDt+abneSiYwAtxlZea5WMNAP0lWXrDkLCedSCs1EI
neg42GDUyI3aWB25FTDwBsvVdNiKhyPv7WBBgv1a7HC/MOAe2zsidN3l8vSCftBP
Bz+vBgi2lrp33SyYjcrKW2L3xTy4ddM0wCnh4ijSZLz2icSQDHlIcnCEYMwR9pzM
Y4TBIxXnTeq8glSQQhVs+JDmGDYbyv/mnOeikBU0k5yuoAl50WbqIiVbdKH2iGnc
iNw2PnxA3xVHZFGmlsH2sabPfqQS7Kc5ZdJe+tyvNFYp31Y7mC9ng89zcFkEVr3+
BgWsqjo7V5H19nHA6o8aMMobTUxcTQrT285y/VQn7JVTN4UUFlw9mYmxoJ8HTL6b
Ijrm891KDwvuYqeIK9G3RUXmId4HuIDSZBah6tCaK3HcIyIYRcsfpCUt1pkuTnn/
N02KchMos+KXI9w2GhfOQnDmBi17/R0QR4cgfXUx9mH7MOOV9jI6o95V6RF1RfQT
rCUlNjsALKXveHLaNJ8zOtkA/19HTy/Rg2OfogkxJ/lLeWcXzXLBdCMW27YyCvWw
f9+h+NZ9GUmW8CIiCB2mKIyHSiyohLSkh+2yC0Geq5SrsKrCz+Up5k5cNf/BAw8i
QYhAICaen2aDFb9O0PonE1syRq+Dfaz8wroxJ/1cPJqbszs8y64TXPo1qL2BZMDZ
MSrh7EDGPNXMBvMINfEyG922Cb6O+nAScr9T7d0WvQQQQ7s/C2YHKsQj/o2tNnAi
VFcOe4WawJuVostvI7AtVRRsRX0stMnR2ElSoMJv+ygWug8RCP4fCbF2eM+O9L4x
T1BE9b3pEeyyXri1zixa13DVbRF56dAg7ptw7fvbKiAlHwzCJcRp1n0iZZY/siM7
dbnS/bokCJnsjjm/MTAAYMUkWvHLog2ARDqJiv6dm2BJuN8foVtjiuTka2KGNnXa
D6Nr+7LKlbdYeaj2s4cUnaJ1p6Q2/eYOg2+ylbMFEBAm5sru/EgmpMuWJ01fDhm6
jfJAaKyssb7jJLs13B219UDyCwYlFDsRAbwd/8+PJEQaNBIErxEmkDOYFrdNibNq
STCzErrxd9MofdfPeT1DyQkgpPnuE7SGkQnxFrgoMmetVqBIBcXdYsIPZJDpgS1i
kwEAjh29uLTBwNgQREUqWyKqk+J6KYn15y+Z4gpjArh5K6/V9ZYrS25Wpo4W4Zfw
FD1yTkJTR/0ZJ1yYjO/tvSys7a6kIXKdbv0mAbQ8dVoYhQ+Iio8piK9nwJpbEckN
Z/SLT4e4c6Xf4vecYdRx1nv4FRksbPg4aK0bkwAbalDGJxEifs714j6cxV683lHU
g6fYkmYEivd/Sa69D6+prgf1s0FCTxPYPWf/KzSvO8LcKYzZwKVw8fV4mOkV0Cvf
MZtak4omaZRkRfYJjujcta5CoitCXNet6NB+24Lj1gxDtoQk6PIU4f5yWsfDPJ2W
8InO7fZDBZApSuKiXo4735xq1+UbMT14dR+sDDL/FOdZoGH69mrrf00nvDyA5kPx
LQzaU6d3tQUaqiBjlPwzsHOdO26K+/zs11M/ZiSCjDoWpj9jZlLroP6cNNEVkQon
jtg6ee6Gcubtl01A6MrAvTxyTuMM998jr5RRCLIPf071BD+dwtEzotR2kiqcdssa
C8BLtyNVTbNJW9Dco2A2BdkSV9rt3oFle8KtmALGQ4fLKZ3Ozyd0vP22RlGDRZwL
DtwigdYN+lkJE7mjOJrdO/kHUdxdHRRN8m2I1rUthwIYYJa0+ZMNaIvEjKAi1BDe
8NNrtn1JYP1pteVfasUfARIGyjXXgTA9nFOaVROer58uV9F+krRnJB/fkiysBaWN
srTw1dEdANgRnpo8TWaxWGlyYWR111dpoAELPUhfUH7grdn/svH6YWywSd+OoRfS
gOKaUqpruXYavAOGhtXT/CfvK+qrnjjjc2A57xI6odDu32sCgN1sk52yI5rJg1l5
3bdZqmAW7/RDD7i+6TzLoneumZkDLNfB2/h8Wmvebd7If6+boUQqVEE7lRg1kiHW
q+0TVCnpI59tQqTBL4lDR9K/kAB0hahl9bFfjz4ET8Yx7tkAfJraXKFShKiUWz53
z2YY9KDRdgKChX9mlqv6/yQEDwBHjNAEpDCb3KoRFLF4lUYQ5uvV1B5z35zvdoeu
9wvdhoE2XAeTQ8u7iPw6DI8VQC2PwDOvhjTHWwQF4A6rYWxt7lGccNcrST72ZX4C
HZ9VONgS3CllioEVV9MS71YiOqw6P5PUg01m/QJihyd40/ENVModDUWtALaTa4lE
A8FIsfX3eJ5L4N6w1PU0zgjtio8AwLoRz/DsBEkQl8Cbadfd4265DGyOoObks4VW
7NPlILFVbJe9P2tmx35TAUGP1M/7ZSOTjNp4SfUFjgNeBRxRBGvZWGDBxUNOf1Da
Yjt+TaJOSv4FnUNqn9GapO9K1B65epfnw1/ekYyuKccChLB5fUwDz3T9Lkta+uMR
sqGlvNQSfN73QIWihXQLIl0+821h3cW8kf4ToWkKNbNiS9IFn0z/+iHUaWMy1Iab
DLKDoZ2/De4sfD93vvJs3ahJYEdMSOx12TFR2fGqUOIjodS0Q37FKMup7ZRQEcvU
9Itb0PiA7PWHOjDo6lTjU6udpZ9C8H3SdPjOV9gk3Ln73IwyXu7yr1EftAdjcDkJ
45LKD/tVPWw1XpiYr7aooayIm6ri13XN84eD88uOOwBmUHvVA3bfZTvWEAaX5nai
zFdSp3wVEHQWejA8Osq7CQFTY6Ad14viOcS5FuZeLvjPHFfDAj7hjOIuFGwJxIwx
p97Px4qmu/B4BfEuIwdubKsWK4HRSYM3IKBVpFmumL6+zK1CsXT+m2q+vAM47x5R
o82EcniuVCodFNjJdV58TVy6YsE2CjULk0J41PltpZAWDMQiDlxthfQPqMc3INHl
2Oja46a4KIrvqkE9R83z+DooB8icvnQdR8GV1iP/9DaJyUIb8iKllzAl5JjjP6HV
EKjUWnku4ZHt8tKhBRLiK4L5Glw5oKiK5ssk6ojw3kef4RP1NHeA3oaHV7X2cwt+
pPoMNeAd8M2dPDaUcRsQCXXuFWpp5lKhF0Bbsl1U4Bwb1Wnp65uN5b4rLCpqNY1g
Z17SKHenLNsOlckOUeWKUi97Tzor2BcJ6flG5lP9Ey5Kf6ONrECeCeWEJ6SUsNWb
cUOIa4zZFWO2sE9IfW3DT8VG6tvYK3FDUkr2DgXgZ+ElWBSl4sFbKkrSMtUYjhZO
6R++qk0/PIrBevsX7BDyh162zG6yQuLd6KZ7POtgIGjeAwIK/XTBwDJQ0PlyJ7w9
drN/Q1xxaGZ2sC07X2o+upUfh4K4L//0qHScMrCHDBFvXmiHcYClWuXYYUbE3mM2
1jJyLG3Fcg5wuKsqyU9QmyHoCPqhk6xU6qNZfCuFTymIY76ZNbAPjFkIyVYWWACi
Cd+8KBzIErhyMFhw2VeklgEM2CJ5QfbYyKmRJSQXvHxPPO8g8qstptgZ1ZiV240M
EicElwQHGHe6dD6lJW5kotLIoEgV6xe6B7L/xTmYuQ2Q5hDUsKfvojlvNQ7GRZFp
kgVD8bTFvvkw5UZYeZ4ECg2dF/tRvKoicK8Z+9Fv+i/fPoRha3YA1sTf15Z32BRl
gOK1C1gGwSmaLWeUed7FmhLnAV/3xWDntVk0rAr+3UqjlPZMI4t95AC2qUBX9KKF
f5LjIe7lThAMidGWDFafH1nZrvgvz8BqVjlrn5bX/SK0hUZ6UPVinzf/Z4g65JV6
AiTYp8I+bRd5BxoSuai7ZUII1FaMf/bozJ3UOKN+LTmqrjO6eX7f92LVyB+cAchX
n+793p5ETlKWoBYyxVz+W6NrYnmV57QKxr5+PvhnjHemq2q757s4N4QzXQkLVSy3
SS1Jxcd6NrAxEi9ggNipYWRC+HEhZv4KSQHiOdMdJ5CFTvWHVCCTHDs0yUxYC6js
S1VRlDMrhi1z5cNnH9I2Xxxo8vljgJVflDt9+rSVl0edlQun1O8iRiUysZP45dCm
Cpjguru2bbo80f9ofjJ/nSw16/P7zK5EMTp2OC2gBoXAcbM0g/SU7fpFJotjo8sd
6oxnm5FX5pqTmZQYc56pdE62Fz2O5fHYvrocEnRYr5a9L25JinBnYVdCsWBpLIU6
4iadqoIRt2rCNa8a3ZSR+QZG/wqz/mpL/7JHpCXkCDFo9LkZ73WcjOAbjJmNuWTb
zQJnz74BL+2MLLYi1DYwy4n4tZ0fdmJZDpL7AyQ5ywPAtuUBntx63sRXsWPBkvUc
PIsxu4Yo3dvGxQ8dEq6Xfae4JzP50/4FFQQBNa//ikNtDMv8JAZQdCOiS5JwPi1l
AgqnUxqxrdKg9SRLHdxBtlF1c8w/UeFQwrHC9LsvNdeJVA6VVdHLUchjjIwnvGgN
3I9M5sEQf03/wI0BcC6/pEUIuM2EgHULj2wG9smWBRDGLRxahcpuQoubgOeW6lUh
sufXh2Z5T3AzZPJn70BukMQvkQzl1LI9jLTiQBr+UYpeWfZk83m8Xbpe17CC1rUf
gm9QoKnDZxaAo0W26sMNBH/oT4ckxQkznBTrep8SBY8C1GjcTR6jYOYGMgbBYXFE
8l/lgDQXWqH5CtJ+G2PxxiSN+r94wp9aGTdmf5smjJJhNye4QUhSspCsbwIfHbLo
x3Tmd9qy3NHKfvnkJEjH8XQ1Diz3SuscmuNyvGWVB0sP7DfV0TAX4eYblgg+Vx/P
GE4h/5KLMoGjuZ8MA4RHAQLqxZepUhLA8x87qxkhsEodF7tcQhO7iiCoCFNUWHHH
QxdpzHnyAKIqVdffm8xHRpW8U2E4SoB//OtkCvyAF4PWzrsixJkWo8MtHCAUHJcx
uda4OQfDApSbtALtXPIYokxjT79OmYB2/m15xlQq867Qb6xPDU2u6/03ArFfr5Wa
LJIjxjXn4hUHVQHDwSIjAm8EuuGZQ0U+cwqsG5PZh6z/EQKVwyVYZcBp58hVnEv9
ES1rcn+2Q6qYPOPLRFKzKmnz0dPG8Ryl3AI01NZhyABJy2ilRCUwZGCUf06NGEIt
Jkp3jnjqNbTbLxLKcenjNJiWsDVG2qF0+U02Mi1PS3pPdHJhL5vqRnnkITKIqBEI
u34BPz2Rfl/srWEFOhX5GHPXKtOo59bx9gj88eqmxpWlZ8JpR8Z6EtPgDPY8VGdX
GjqsBHRJF8Fw6Keu6VxWZ7cg6+QzOraCop4qxCcvimKNTl75zUYWkZTc0bwXvYDX
PDO5EGyqku2YsJ1qERDghO0myuZugnigJp7qwN/w5xJomzIeKXsnl2txJYeAnjaJ
sGc7+5BbQi6jwVuVEELgxGyMNbbnBqS1TBJRJOU4h0G6V+UViarJY8Y4VdU62mbX
bfecwxl+/BdwH0GrLaGJUB9AVbnXyGGlab/lLV+N7vRNHauMaGpuGl1seEzeQq9i
717W5PAZvYSwPo4VbsVXAVJL17Trj0LBmb8TEGonWaZQ4iG4mOLQF8WowtKa1P1O
6AsEU5gq2bq/2RVbDs8D/QjnWKZUzinIOrp6LTb9g3rV0EuaAFfwlpAO3AopAN+9
cb39D7PI8lOcq2ZCynE9Eo1V3A6vfBOwCfLGUnFXZwJyHwCPLrIHcg6abuRXry2a
f+j/h2Gpb/pXg61KXFrIRezjNjxv8gNpCdKwx/qhzEWWpXHYRmNB6Rqa1cerLMdg
G6IyQFlb6tFCgyi/fLWVmATJHB4dq3qF6PHFag3Iub9WDx1ktWI4IN1CfVUTzlv2
ygwWL7BDWQHuo50nxejZ3aj3tO/jrL2WoX2lkOGfsGZ4e0xWEsA2vQwJ9+74/51s
sqsqas/gZxtGn+uQCLy4sdltAb+t8ipKrdKZjR8BSP++evDXWJqETSZ+mb4cPfGP
mVnkgFyfEZtpwsc6+6ypdRr4Q+uGJFnApvn/WitRUvUuxHlc4AgsGtuYKdwGFe52
gfrbZfYW4dnO2I2xeiGS8JKcn2e9fYgYPapQO9814qCnnlVZ+p3qx4SXLr/2tqS7
spzvB8LNidlj4tXpkNMgTNCZGN7raptaXxb1ACJgKGr1+1VpopLWNfrAeT0ZX/uf
SNZwSnpiOdIqCgOBTMsFTVuOlp13h40JqeuDs9WkUp/h/x/7Dpa4EzcdhWntc++t
ddeG0rmsGpRg4EkHSXGg1ynLeOfhSH1RP6vYevuHFq8YeUBt+C/QeWvDMdBlAPx6
YrddEVQI6qG00W7xqsFDphWunX+CX/d3J994AnuLaKE0+dhYSSXbOunCILnpjwbB
kmNTubO/Pq6qpEV/xTGR+pMFK09HUFByVZ0xLl6J3TCSPw9NgFfLxm+GJxWABveH
4ucVEGiuGxC5duFBufN5gImkECTppOsra0F4tQzbKaHM9pW8Pt9NnwwALByJBpTH
YrDaAKF6sRuBrn6KqxPaT96jR6mHDD5zhnk+mg8CCBwAFLMY5W2LYht5ntSaAG1+
YrQebMY2TgV/QWhtfIjSw26iWLTSz2smT788DJnWmrzUebJRIXleJ5lmbN5kLilN
p2v03wdtq9ARQiaiAQFAvZ4CHeTDDz/lKOw2JqTt/fd5qabBSSBHBBC5z/YQwTkm
W1O61zyWEbC3E1huOgsQkfn/kEC3m5dWjvkqawawTqFWJfxADaRVIGfye5I/QyU7
b9gAPh1C9dx8xZikhb6E+OvoKUwt76RMKOGsHSOJ4Hu/DHFJdhUweuw0vIvLJQXW
pd3TQdDfIhIAS7OOCcrclFPUSsyYezMHSz7YX1FmNlTvp7yerIOLr2tshh5itppY
oejqvawH3nTRmqcF3KHEKNFedW5/ddYDry6zWXjLdmZWueuIDRG4DQ+STYmTZWj0
CeK4TTp4r4/SEXaCruLyCHfrpEhmi/IAMePf7nI0lpO30Pqa0dmMsXn6eOJeEPh0
R0eNUGgMDV6Ouv/7/Sw5ZjfTKpHRQSOhAVtkXqnacllxbPFJgAzclCcpzqIPC6dY
VQikc6cKz/beJN/UUMfd6Ot0P0Vshc2mzHDxAdmyJDZurcCgS6sbn9Xuy6JX0U2j
RIRToqTt7OGwHO1p7nurDnESkJJhzXnIJJE0x61ivrzsDG4g2n6XP/yjK06zeBuE
quu7huiLNGRGS9+ZKymOYwUQPKsCvhzHibyFrYK8eCg+dICi2QXVQqYrIzHleiIR
VByZT+3ylz4PH0lMWxcp3PKLlFZNmQzPIpBeMfaFlF+Pu0cW6R3YZYmKcYReIppi
0iL4OGhSLotYN2aiqYlqsEt9Oq9A3vycUO+bGHNJmsA6ThVYOqGSjpj4MsBrGCNZ
juaAg8DJnf56K6Tpv6mE1UanMk3KMVztiCHcPZgtoln10FOazVQESqcSrM9LgUbi
09mxVCdEfHA81QHYwtTC2vio1WEIePDKlEPwmuO9uxgJqexVCbsVbkhuuS9I336e
fqyDcCuELigm97+ZtE07F9wEqYoZNsex+eryh6XkcZdjysAf4C5VFi6Sh0323mHe
SWGgHo+h1Su6ds5HnYtCHRWKuR/kX8xS48LD8iuGZGEWQW1+POr/aCFSJHEqeBbf
jBbHdgVO2pQo1Ub+ib31PXMhmd8zU0i9LK7GodKAGbhshc1EmgQMnbNHGl65+s7O
hLzCsl4ufPTBFsEIuFsWMW/yvpA420ZCEVOv8fVWlpdT82CDOr7R13md5XBt19Uj
ZN2Q7Rd7n50Dw9hb+MweIL8jQyo1/n305gdob7ASHlIBThRjvvEKPH7s8DASOYyx
uUg1mzzo7/qJ18qD2mNLHk4rew8/9P0kIAhPquYBShaYpfQls4uUTwIrxt9HL5GC
S/+/D9+EvNG192SqsvvhcQBpGUw79Ni7JVoPijKIueh+b//xts6Ap5yzkJo/fbTi
fxOrgSbt4eQ4giETHnS2zYF6GijGZSgFzkiAoy6kbHTtwB66WxaYyYFrQaX0+dXN
tPqjGJcoKJCAnomDVPcaygDr/LsHWn1w3n1qS8pzw5OpzUbpGbh+LKCsK0vVBfWv
pl5Y2/gvCBYQEDRenOXpJ6i+8dzmwHY4sqMNWcGx1R3TtdNlLp/CGEylb4adljEN
Uc+qpkDBYpMawF800+OjLPA0SEFOgN5hPibbKaQH8fnhPaIYIwf0NCxBBerfa0AK
fEQpTVPjDh4YcCfDFwWlFOwwcjN5S0skmkkL11odZPNcSJgxUztd67C4XrriQk4V
8MK5NPzJAf1qGw6Qlqp84cVdzV10Jhj5hc1cBceMtpLp0+wB9tE+RjBhgEAHQTC8
KSaXUnIyprRTJ7YFf8hX8MvoXcBcLEgSLoRiYvme/mLigPBvDhvucvc647Kuv695
6hPQW4S6NgeDlfLfPhFab0PxVNJusvI7GmUaiZeb/vMZ7o0YMaJUlszIuYeEJg0z
Kx5kpqyOu0ExTvdh0iVHSR3qPWcR2LsY/TZkUMBinN50pd6TXTtzGWofkn/F4q5u
y9L3zCIKvCialqhwFxhx3fpCWo3c3bHvgA3KQwqo4H9df12qItr2Yb5qCX4eMrV9
nAqI0CLAe0Ncg7SX6uYQRyUql5seVj49JegKJoS4/dVLHh6Y815Nyj1BE1nfEb5c
96jDXhNeRqdE0YqNVCqD3Ha3XbArXwqeelp6RZ+/TSoKS17y3VKr1FFQXIM/XxTs
/vpQ55rclbqeVgnAgISoC3R2aohoAzpc2MLMharnOIGforzIMUEA3CssSysg3pMz
lNwwbBEkImp8BZrMhhmPD56IfscvIF8qkS2DWMVENBCH7K/BLEulz9jl9Z4soh2h
kpPW2c259l4ZhKUwTolen1Ddkh1/6BY6V6d+l08kUJKk5UYkFxm5noKUPETNNcVv
eMuLEYDSVeBvSqpZlQcOvD2VENUjhtn93n2AvFPqg6+H9LJ/mvw7bauZNyjdiuZa
DzD3c9pK+6lLidGdt9R00Gup/vsx7Akirat/ldSzyefOuN3BwUX3hG/jw5iNbW4e
7eP4JL9YY8LfQiriomw7vRNJtGZEFuEVOv2zyLSGnATeL9OwaArfSQRQxB9lNXNd
Ln8waVDrAGELfeykXc9n/439zV86fhsYPTl+cjMNPpKhx+dc0qQbcVphhsxNmPpr
SqxHHQ3mbXdReDwL+fRzm6mOqQDQZutVIpKj4A3o3qdz9ZeyPe4lMQNAvsa23ZhR
hhJ/f1laLLZFIZQhqIJgfskkvPkDVJ+GOTNS2asNu62NIAjiG2hwjk9m0S7Po9s8
XdwEkLSAfErXYgvQAiBwuUdEtC10U3922flcetKa7oND6TPBcwwOx4M14T5+uTQv
CIxc7pFuVLLWrpcksPjWPsLEfAwKyx+YcYJWjB8CrO9BQyd37x5nq2W4P11FbxMX
rnRXroZc4eHLHYUqgi56MBeXLDHtpx/j2GR7G8HTqlRTEAJRatENNqNzXF4bLPCJ
JAm7bKxR+yXr5xZ+lKi/eZ9QOH4xoeoNCAF/v2h1esgZVdt1rnLX7S9WleWCry2P
/NlLqdgr8CslE8nHEzoRlOMw96ScKmj9nMyk//tHhjuGLIGz6Z/3FSmSgeKlOgcZ
IM54B/1b6BeAhl4YTDZYEkQ4PY5W4R0mfZENnrA2orSTRKTG1NFOohfP9SLQAEWB
X8FktBBDh1AQcz8P9zfQBfe9mHlPQZXpgLkfC4dlDEIKM9wz0AgWXfhyYbA8DmM1
3SNSpL6aHbJFmMwqpN64P+NHF4JLwR5rmEwnK1isQA0zQDAfD2TmvvfW73ynGqbm
I+eIK+O24FIUa5lyPgDJcSe1avUJuxfIR5s4UlmWuDQr24cU3BJnU/UgRB1nXq4f
mVVP2DKmUrt7LKqGsUYSa0PZ4xJ2CZ/QMDYKwfp/vlaRGWR4Z151fhrjiuYEBZGR
Xh9RiH/2KM+z4Pi92j04OkUTiFHvarozIo8jRwZVKQbaUhkkW4ASw//Ol6z/ZBNL
bz8vi+ifnYKddADLhy7x8hWT2HpoGKQXA+HAHHlxVcC+LTEelTsL8cLYkqOTjDuS
rodIO0mrUaecA9ytmR0B8nrzKultwnLUNROHoQaWYUO5XDYHGVxyqkvhnSe3m3wU
bM2QJrfTxnXU380mbFBCfTNgrmSXE0iqkYnlGGHI5h4DrlgyIzcjUZIGVwxgAKj2
sO/BiMVOZHpw6UJ+AtVqaZSvjKDGIX+obFuxQrL7C8VC9C8o54Osr8a3ik7G8HVw
wOatX3U9B9Jktw4S45yMcWQmKvuO/JE33xBg9zdct4ZQMpbGY0nHtD/MeBBbCc9c
fzo2ezZEtqGS4pDkcpbL978JkAcBwU5eqeb7+Ss7quz99DZVLWFg7mMaY242EqkB
L8Zboy/WOBdsVj5NZjVFW5Z9HRkk1omp2RRMO5oc+ptw1uPobB5iX589hfw32oay
DsWaVRIpNaBuEo4QtsQhAZjtI/+v38PZgCIrPj4APV4RuQYsD6t+tbeXhpa/Lg2C
UHxda3StQeir8mKEpQASj4BsV2bcdLdrxp3DBCX4282UT62+YpFc4loOliVay4k9
qcEMEkkhlpoTNrKHv8BjeyO23zP1uCMcnA8wkhH8nli7ItcGxIUViy3A0P/KG3fe
wYZpPWbs4okF1i2iSwL6N0zlLb9PHKFyD25ufcWjoTguqbC8Wh44iOIRuzKE2HI3
PAj3AkTZgo3M9fxcbPWhPtXS9LO2Xzhogd9WpXGTZSyXyZreJ55FzdUtZqahdEim
Sv2+XdwZOZncSDN+9Jj3wrECc/4dzF2/mUJV1qiIm1X5/xx3PZhsvahc5Ezqe5Li
S6Hqda8ajH8UR9pRq+YxcSWBASBYT7TixWGmX1abD/MZ7q2MqDOhHQ+qPD3/3xdc
aPfmgQJ/TnTUvra2dPkhAbnE9gMDUeNbxs5EJ3dC8YUnIzkW6Jj1lwVokc5EyZM/
dGfSubn55KQH20dmyLu5iypq0NrWSEiS/MHjgaVL5qoJd+IZIWy8+0tT8RdjWLuh
ClQwT/bXSE2LeA1RRv2usfWe4cCIVuEaHrEBMKp0YjEOVNYN25TkURfBcTUDG/15
LfvI/Ce5Kn9n8WZQFA6P7tqzJfuEoszefvKs1kTGNjY2u0kRneGzk8kowdOKOkdG
2kBrRYr8rXyMwKeBbXPR4lZlpzp9Ee81nRtW1Kkn/CK4fgssVXsUrpzreziiFdNt
oyyHnsR3uoO5Youy4ZqOBilZf/TgyE3w2WNNs31CsZH/fngwTAaZQVzzuspwvzQp
0FhozlgQRkrUlZxnyq7bdAHOKwejBqJ1WRFqKGVDI5NXBZpla4hBqmkzFKWQjnVM
yFM8gGtNFxRmZ2IIHqmQZkN2H3zz1J0nhDscAuGJWKqx5qUCeb6zooq39RIVter+
9VHXSEpyEu6seCMZhR/DQPH95DfEqHjTJPcXt8ppo2Ot573vnCzYsnIf7vMzaZwJ
EZQqlId1SYDwTVyHzD/a70edZMnKsrqTxjQF1YFisIMrEKuKMLkZp9qGNqgpK76f
EslU7LIyG9pGyK/3QnMd57Gvhh542AZLLz42eVokcl0eZj4uKjUP4yqWyoFaAMDv
llo0CljYOlZ2J2j83to/9c9JuQfoWtDBBmRwpRSo2wED8uKef6hLDrKJcnSa/Zmj
6sZgRVdvZzupX4T0XV12ix2pt6USbZbewx8II+Dzd8v9Dx9xpRXc6teQipzQPPgt
0q9rtVJyJ7v6+aBM7345S7Giy4eONVRsilm1tGZYZ1qMQlDEpzLN+LSs8rfdz5eT
qHwP+1vuk7i7LiZIjYSY/Nwdki0UBG3NkYr6ZfvIgleZ5TsVC5OenOAn4tVlJHL2
tD9tkL4uGA6Wc8K2bLYxfl/Z4NMzY1oAuPL1UKYm1fbFISXPwp/u2YUQkjhKjf53
nz9T7nWe8Fjv1Uyky6XOn2rchBlRIEOg5RGwPU+LuW2qs2+y1rasMPPIp/zkmuyQ
o9BU1VeeW5aE/Y7qPDg2rimXjYAx549w99uCKsCyGDXBxkw2pBH6cROctbdPKaQF
D4C6JGuphG+ZffjfVeeDfJcLcyU4DLwrZRrvoddUcBrCFGGfx71KBbGIoKxFz+Z2
GaEI33mrXD967UQcP8vwCWXGGiJrZu5GiJ8oE9GhVuOKj9kCv9SIg9gPKeojVcYz
0YUgn8qmcx1amYu1t/Zu1zNXUj4jr9LN/0obk7A5Eryu9XIzNw5NLXt9nUW5SFsE
2vnPj51bs2HDDUckqvuiJEfYp27Yg4pncYgYs8625CfN760tcslntRXf+mh04PUt
9ViZUgUjwaWlVd7ZSB4xuhYi6qjt6A/tHx+408x7ZhcUirynd+zMZ1ch6jML4FD+
7NDCoxDvvZ4XmSLl8+ALbZdhnZyu2n+EOQPfigRDnPSawLmcBXne6mBMyXI+5HVW
Il3vQcF9CRb10X6iwKsTkV48uQJ3h7o9jguUAdwLsJKGUnY3H3rMdD3Ef5VXPCTD
/2oK7GtIK61xToqpz57hzhk5BIjWIloGAW4MzFGb9f/2jXAr5Tjxp6bjiYHbGjFI
rDYRPDe0HhuhnniavijhqgCQj/dLfVNxWTMmLe9ZK46i5WJ5cZ2uT79htkefJqHt
iqJgAkxyJ7EwIAKYiTU7jKJ9KzqCbIJF3YO5GhQOOP99pQZc22mQgFhv/HpuRdRZ
kMloWdq+4G4MSqKqs7fxz9e8yNv82BCQVj0ejiFOip7rn2XB4GBeCnbu+LuYJOfm
dOQw7s1E6xFhgEV3Tc0vi9pvSnJXI+XLMkabh8E7M2E//O8CDk2NIwVPhOGWUnIB
q3RRvFqjp/3wwWRNRchvk2LeR71zTU4iMgIFF5JuOJ7LT0K2Uj5aEX92I03UR7RD
+PsCRds9ZJ/JU0eEQDGEuwIRMc/MGPT3dZn10gNOufM0wcauSzXsBVTDRSY0sACh
HzdKJZ5RnswN8lT/sS0SvbfWFodKr34F0WKTMcmR87/wNEw+Ogz6MS20KLmDMJ/K
o3QYYBqOaFWAZ9PtnM3GfcKNg05YaXcjZbTb5ZSc2c7fLpfyZifg03cKJ8ojduDa
4GheHrvCgR5KN7ReFZ7qZ+kP/nsguXogmJOTb8LsGjrLWZEjwQkm/NjlV+ngAXIb
ly1dy2doYGVcHwaGIJr6Uv9vAMKlKlopLaIWb76IwaxBWxENJDvurvGW7WyxaVSn
RhqYpgOwdoMwb3kmBHngPlHCM2446uxIqNgl5c9w6llGTfjcXXw0s1+B/9rm8ZLt
x8hYskYgKwXfEAUr/Yuf5O7qJYYX5QPHM3TmEXCe6sFpnttrV04GRtV7HXR22sdr
5wTCkRuqkwiQOqWR2CxZJ46hCJS/LXZD8jDR1hPVLTyIOmAWdZIxUbfIAwSoLHZw
YdTsSVVqyWCuiTfBou8hLFeXWLV9Mt8UWpOGZjXA0fMJZAQD55x2nJtMsIALEXjq
jzzSj9RUqWHWoLTPfWP7l3GOL8FyQ07wPrACBCmpN/c8DsfIaHoEvfz7fOWd6Bpe
B1eL0wUOo6o/jr+AW8woBBaJW9RsZeelk3tHl5M2f85G1cCrj0JzcjjjCU6CFwPT
kWvmxM2X9sFVwWRaeMiRwY6Gx2ckceROUEakxzz9C+8p+X+uX+tYZSzJEw2lR1VK
m9EUlppPwnjHstvbZqdOGRbQNJlOlpbsAiRjxow+hbvcDw16b+lcN2uuSkJO8136
Y/kdLmcCJg1OUGrHwL/3rAHtjBDnCL3of2z7N4wDJjEnmTTJ+YR4obQa8M+mZ+mm
HAVtp/Akmc7WDtg+OK1VIpHtFWNdwMcNmQBkMZ/yAIfho77WvXBUu/O5lKEbK6Jg
1sOdVlJJ8BzvIJRD6CQ2NBUrWsdkKugG0BFnepl543YWGiZcOTneYTjyTOF6C8dK
+zSPn5SUyH5m0H9ax4lwngSdoe6zJgO9bXMqzcRX0fuNkV/yy/9RQCS31ETBqLqF
XxXbqzP9W8cZUfqTEXDf+QunIoj+7eVMTrN+nE3VlAQDf/o2pBP9u5SgZ/wlOpld
Js79DArmqpbbCdqAR1kFpr3e5C35RAiTjOxxfz7WXNMPaTbHQ+///E4rRCNPCTEw
HEaOajh4Nf0gOF+dYrrnjQBzcpyeGWpPHTEBthmsFLJdxxLyWClvsEzjaRE4nHCP
PCqHxkrVHMV3PrQ0DcgqHZYNGiaRVgoq1yJVFlpRxPkXHDCZZ3j+Q44HPNICcZhz
RKYhflQD5qUWhu5JjTWX5yQKsafikEVgosYxlK97PcP1FOdyT2RM5ocC/dagziul
nbBkCG/0xaAaukbsyKvRs8zpP30NEYj7yG0dC4ccvYWKBh7Bo2MWoJQtPKB3wlTH
YARk8DhaLsi3LXQUOR6h1aLgP/pEmpPrCOgNRI0sFPUr0mux1iOunSkpp75gz1lv
XSiPz5lPQZSKIRFRsgO7gGr2dMrkFWyKBJfzGR6I5JRGtRcLqlDoiaYTHr1gN/DF
4rzPaVGPHqy2xrcFTNvRAn7qN+if33s1pWU2ITVHw5JTKolKmrCE9jaB1XA6KGUp
6+pdKUWMRoq8BznwrU85PLnGS7y01Da+MDHwnN4kTi6NNXe8qwUSzJeVlR0yF0Rj
DAHASSE76uUYGqfDMmJttbwW54HTyFD2mv6XFK6SCLDyqQra7+x86beoyU7cTWnM
nTuSUWLVVi626ubX6jIgvZnXE7lRG/8roeyptWAsfAAH1on5YLyFQXBtG9PanHpn
fmy4nc+XWLSiSgvrBA4+cacTNbkhEZazqlUUicc2t3zS52MUKbAkyBbtrbGYxL5A
JMnQfAt7IUoX4EAk3byMArktJUvdRfOiWKyVka/Di00t9tN28ZQSSLYO8/FlnbZU
zjXfVxlh9dHlseKX6b+bLQhQXw6LTb6+DfsYTa7djMll0J6gUbqSgdNCwLD8hjXA
UcwcN72WP/NEFdetKLxmSH2DGEjjIMuzWzrFcVhd6KjZ21TKBN1Sx/DoQzhvus3X
ppd7GNyh1nP3lb7TVIVuV/iRx0dmwdZR7N0C6kMQWjckyG4xl/UAeuuo3IfQ+RhU
e/zzJq7vX0VXhuhtg63S49OpdEj+VTcBtrWF0i/IDlYtcLQYL3g3QdAnUl0cjfcO
ifCx2wDM5ft65Os9LDRISrcHkbADf3THsyKkvyrrCDOZY/mU4/fJMHhxsX0r+rC7
FNkaanAeLiZ/i0PYO3tV1zsQJ1zRmafVid/+PlfZ0VdfsFyhfk2YjyW3mpiAnEed
pgEKnWIiZJ4vT/ZouQCvmHM1DPPZmLcFZekVo+pPFHQ3BFo126Ds1wbYEn9+zSCj
WFA+VB/WwEEkcBzzagbfbjHvK2WrN+SPok+GfmPCfjlV2c8GOs1vcFQgJPq9fT2f
qqE8Hq4hW/NWEtHWqzZ04fXkjTne1W6wwNZZLaNKovS/BgrHTamudRpN0rQMi/Q2
1gkwJ0KyjIDc8a4joBK0EpZab4O4QtAY+pZnV+y/nf49J/s6wj9+JXKeutnjEaNx
/21xmdEupPmVH8u7t71onwWQyw1OTGeI1b9P1ZqLt6RdycjxfmY9hlc4uNwFnq98
W/QrvIcvFICwH/c7vPuwyhglxED63ijbujtcd5XNpo8rmXKmck76wgkqNaYUPvbl
L3RzltIwqfPxDz/dRUd6l34kqC4ke5sRqpKqwW1j/N0abSBZvJtaKwTyytsepSDV
7M+qngAHbbWkEs783dE1IITemHYVJz7i0WNPsSKCyo7wvk8LsDZa2QXCDD2wqJ+l
fkbuNREkM8DXZMyBIM4wf4u0XLlh7UizWDwgyxWkpIh0ncg3RC10qw65XDxzwCqJ
bHYCzv9ZLd3AwIWZ4un9hCzRKGLbZxD1sptpQK2742QlReHHIJVhdh6zm+E5mkdK
TbNSJAyJnxsqrLRGrfEEavRgDhl9rDgIQdZX5ZZGH6NBrrZjFQQGBmRBVykMWNwE
vpaMfseEeJ7SSVd43DlggesU7X2suX8Y+xVM6ZIiXB65PxiSlgo5BTaJHinJyuUH
CpBeYrV2zF//NNl5E7WzeUiU9cZX+0NbqPJxrxgMqX93caead97/xWzUc5L+uWQO
Sd7AI0NY4ZG2L73PwUemuiG6eWkQ4jjMkP7tmlDn4WFUQwXyeWqTcx9ZHtQpuIg7
7/pqIfvr0OYPwFKS0st97oY9+EBcgs/UyDePy6/NHbdJIvmkLn+ZlIsAInXhrVOA
qBvvyKbyn9TaQFUpfitseFC+fLShQ5vohRmaJnirK+4rQpDTJhSMf1LY7f0BEX2V
DLc72099YQs0+aTE7cuQs5cee6Ji0+TjYf9MSxP9srHOtiEs54jrn9Ue58cTNdzm
NC719tVvI92cZXA6sswPdpI6uTBCA7A92eSgt526mLsGW5a8UDpnGevlnpPBq7LE
1ZChtHtv8LcBldazIIxfSDZ/Vo10SLiAMMTeTAJuHCq8SD5ITyP/v3Aj6CcGa4y6
mBCxwDpY0R5ExQki0DKbyBAYUGigo/cfHwkBPQbja0GTI+/qNpJmtc1tDBYiyJFm
DBiZcwtU0fkC03nx9hvtcen0WBLgv/6yuEqgAOOJ7QNroRSlMz13JbaONleIGsJy
j8zZEWAwV5ato4xGuWegOS125uSaynhwtspHPKLmLzRmHg4Cgm0ot42znKXKEgvE
Z4ykuvQAluAeiNKd6lKQNKw0ot4bilOFYQNas0p0c0+1SVQpE2T24jbYuhcvrl1o
74ev8Hfp+/6tmH1dRKCeeOfsR4i8/eQnVVCOI6WSyBFQk7Hmi1kpXfiBatcFCGEZ
3oprnpp3vDWjYSXDd/JgiE7ZtFyyrxJzNDVYzHzJ55+S9dpbQ2sjj6/KodVmNnkx
ZeqCwclD2i1kKA+KG2iS9IC1st3yVwrr5KZ+OKtYKln1pd+aySHyD/OY55ufsmml
GqJMISaFct+7KSIO45lLnLNM28Nbjf1mNg5aGKjudkm8/qVDZMBUF/iN1w91gCtQ
6U+oe1mnjMRNz1ws28t1d9c6FiXMi9vYyN9a4tvLWYFrHlh/SSf9msDMSX3cVn/F
RwgysbOzViTegMGst/iJOCBe5iJSbsjwwlN4vDkeMXe2BbbQxgy9E7MwzQzfxZzu
o1YA93jPJ+iYNSmVd+RluDv8hA/U+aS55Cx3LZfbX0Bu/W2a/Uv39Zv2wlmceZkk
9SnjzOKJsEnt4QhRUFc4CxQnrJZwv2hURAAx0RjHOt9PlhxKWDpUL56MKMdvRdMo
1K4o6si5tT/onKV+34R8vEn4W8EhDuUnrvV7gDGaCrLo/VTfd4imN0fbGVOp2YQi
xYKstTB6DQRSwHVlc25XYqOIvm6s0bdkM/cY5+jtcDnSfkn6EhiGKAvfUs1+DNdh
5uZtET6Skgxbgy4HsfwuJ1bo7PYxZR5jhfJJLYrhr5TvX3jp1NI0tdPMHqcoMHAX
AVYctvpY7Ge8+a2wU8C9HGneFOMWGKTO4Ck2KOQgxw4GLBxqj4GO3QHZdJK87STN
tumfzIDv59jG0mpx+tfmJr2xSXLbN2OzN570Ogb0BpyZxiv+Xn//2ysufwSt3ZT9
QEheh0ujCHeKdHXWGwGgWbV6BMCWLakAdr1Vg9WD5uvHsRinw6mucPrw1fliwL/l
SZzQiakZ5kV19nhlwl97XluDxK9Ipl9fOxSUJuYgUQox0KQuiVJ71nCN03s88D7F
5VNqEk0gG2X918iIRZn5cbzEDbgEl16EKtQ5NvKxlbsgz3jnMNzKUCwWrfgthceD
6r85Lb4JqIuTEGtPMNFa/imye0xOWyVUictZU/bmBYxuTz45wpJljNH5je90g4Mo
RvjQG1IgSLUF9CaOVGk3fB7pfzSL7M2o/WmN8RkKpFc3JS2vxgaKPe1nvwc/PpI2
o8hDOT0NjMQgQB0OdS+8PmjxYwYFyRH9cpVFXggt/OUoz1ZbcSgdkwCZxX7y36QN
DuK1l4DKad5Xr2nc+NxIvfhK7MqisbOaUFY95JHFuutb7iXX5S9A1j4mJYzAiLA+
by9MQozCq914UekGOJlRnhOrFWUsBwgujTAMYKidHZ1Ib0AiLljUBduxeeezOTi7
jsdBACChWNloVSlLqWvlvSlDFbzL5GPmGPDtTvA+ltQmiYdqbhWe1VvkLEt3dYkQ
I/tOPfWHHZmCngHPfEZU82hB8EXW+6kW9i9bKXVLonCQW9QyN0rl1le9zdUVeV/r
xia+6qW0BKEHJHW6qPYQHkrsE2+QGNSndJA/pR9WPOHOuP8uGSUWZsyaUm0mxut5
Iz5ZAXd2u8AM+eR/nJvdm5aAu/pN0OvPOnAYeqePIdqcVmMiE45Da9s+WlcMZLVE
bF2RPoFrmzGbo60KTdb5jqnatsgIqUV3agocjm2vNQPEAUPljcM2eQE9Y7Iu7RFb
onLCh0q7Z28DG/wfTGlTmD+m+fsuo4JWv/1RdKxBa0TY86jHV7DddGimgfuF07tI
7RunzbFLCYbeS/ysNThTAABKMMegoUFPZnFx6ok+f8JJX9RmAtIZiIDYPm4SVcWG
a0EAuiUlI2lNkw0/EyIEcwpqmDHYmEL2OMVr8YmSSKbqIcPVldfj34pLJZwnIwFg
NOIy4Z7PmlZhWMA/V018XuhJ7DE+/bysJkWDzmpswqDcx8okMQszaO/s93MkYXmR
Id1wfg05e0Qbf5sp8NjuCoYyPLg69dAaQYQUmw+nRMcoLx6u+eSuMVkTRy8MHjWO
eMq4ojxnVzmuIq91vLCbZC+Uqu5hcRgIr+04YOu3Z7zmbgFq+Iu9z7ChEJBEBQY5
u/D8yaQ1QiEKFEqroixVGPbVZkSBALQsoTOf7e+VcgaAPbzXvcTO6se/hAAeNxDv
syiUDZdhbxs+trBqqyiVEtR0d6YjM92urLXAhOWGPt2htle+JtUMYjhOMXcJlwRX
oP1cq6LXYBbZFtYMEU60GsmBXGegjBvQC3zBMiAIFjHc+Zi/x+I3mx5GzUbMNuzN
H4rLCqG2HYvTyfS8kvKRfs2qwh1sjP6l38bsnNQnLD7nWjrC4O76nl8FMyhv3MRP
0+8J/6qPIK3QcacVZgu7S1p3IzMCQ9DuElM31IGJRdHvrNnFhHE9FuM1T1bQ7z2r
FfpOdXSmjjvQVGDOkQ4rfSDjOwyIBem2wpnchK0XozGJdS5weabYpi7lOdEWr6vM
2E8qPeUt4z9G+FKb9OwM3+1xW7rdaLzaYqnOiDp3KwllovB1IM+YP+0GyN0A5IAI
EIb78KZ3CZZTh1iwUY/lVOCd9ZFb6UI0Dla5NmA+hlyCvgJ/Ni9EaqzGPPx6T9XK
G+guaFTTfoZlJDH7MlqL1c6ALt/sVrvsN5PMGKn3jZx9YZAQphppbWdbUWarr0wG
xssXgT64Y66MA1i1nYIHn4AaPEWv92wompzVTa/nTQRUnxMZmA6woJrKq1iqbGnu
7sQQuIGCDTC1j0+J6chAGk7NJibtZWl0OiAuFW7j7ZYGTug+MUIWKI5ZF1cLGqiT
0dK1D9VY6agIwm9pQ7MFJXTsB99+NvhCttzoTuNSI7ADQD6S5/x4k4klSOSqOQgF
eE0GLPNEo9n3WdVQAwppkfOinKY74/dADRkhsbKI+h+MsXItsH5TodYWTJDL5DSp
qX5zCly/d6qpPv230tEkxAwTCkbF2zNzpiRY7hZAzA4C3p40XagtyDLjfSzToZi+
KiVNoX6wrzBW+HWr4fKBebhDQmlxeGrl0S5f27Xh78Wj5dLMbpA9voT9YMtuyNHN
xa2Ojb21wi4C0gRnHj86c8gg/+BlKz+nh/jAarXcIQ4kyxD3WEivYuOqdJjfxMfI
ahAcfWoEGuQxIAg91ODZICKxsvdI60h3mb6h4Owh7SQPIIiSP6QoDgq4tJG6Cgg4
BqeRFjHiiwJ2edKOYkiMNSwIYzc+NfA8mVjlqj43U/gqhJ72TGRsGYqHUAXUxwCd
e/HjZIUnROfBF9+1BR19FJLO5/qPx1e49/SAmZOc8eDPmy46Y2AAcbyajmg9fFkc
ypmS2+/5+/XbTuMjNp5onbl9P5HkeOjlWZc73M4Z6Z0cqRxvJmm/zN9su/vU6IPh
u6XcJa/D3kjetRGdPldwlyIBCGqbW4fIGpWFLzKnFFVJo1LEqQw5JX17jlJ6AnD5
xaCMOxbZZUOCX7m2sYkfSs6RwEWlPDa4uaT73tqc7cl4f/USoT7HAl94Ib5AsSDa
o/oNhTw1wAlO98wFqY1Y2AWSMsq3ugGBXugkLa3uvgLnbiUXqnrh5qlZUlh2oQ1Q
GJXLovsPFk0fw+YKJkk78LGS6RvilU2FWCJjf3QMfFH/r4xZRDgnvnTpsxoEoAQs
ePdj7RsWiOKHo99y/SqkqLJprl5EEtwdf6FQJfqu7ly/ITF5L+Ardf6wtYf4N+O4
u0ae23CMBN8ZuCQc2AIGmQOg8bw8pW2U6ZaqOSY0mdZxtNOT88cMI7DXRCCcCOGd
o/8enafcZFdyB3rOcuEzzRhkTpuTLhFTogPfxObvv0Kbdv9Vkqo3RC5lJordLAvo
lM8uZxWdh7Lh1RAtYO7OnwAP28wcuOPv6WdUSLdwxIuWSjh8r+0nL9F4WXZa5xxS
3s5Ul+o9NgdXl0n/MSuJjwP1MvhDDn27PeAV6DuxftoSyYL4VDDpEwky5B70lRN6
RQUdx/ao4LvwGvzRqi/adHf70a/aZr2kWDPvRJPvooe8DqCA0qkXhlJ/nrCuqPKO
IQo/9gtcGeNJTYfgBgdciDx/CYuGeBzLwQJueB4Xx4KcB64lA0OKwj/peTBbKugN
ww2KAmthN/i2y9n0p3TQ3T8dbxfpDiUPxSjg1qVeUIDhSSvLTkII3xTLlRYTOhSX
02Jp++q9gqz0KnD0fBM8KMMipHN9pZf8jV9YPeV/jwa3VHo7kWwG3o7L8mPY4uQx
PdIzP3ttmBgahcH2dUyzDDP69AvQxF4a/9j093wF49EF1ik2E+IjnCEB256ZSFw/
HhMmDJ8Irn7N7wchFOZn+AvXPtqto0d6w8j+VgTVK/fBFZRUuvrUSQuFd6k8fyAx
CEx/+i8usof0Uys4j74XkLRPAJy1BIQK2uRfWUgfyr4by5C2oyHxNNgezczsN70c
52v38E6dmrIg6pjySA1LoPtZNPCzth1F2gQF9TfFxL7vGMToVY/JiasCN43cRlQb
eWZSOwmYGYHcLnUkQO6OkU8mBZnGIiPs4Kkhq+R7yQaTmyyrf9qGhyzfzyHDPfJc
O0I2o08xBXRqpt7W+Kr4JePe9Yb4k0WXvl8jK2MCdclgQQx6vkrT6heJVPjke5Q3
KZhtXazhhFmuciDC5SzAXBdGjX6PwEs/E/DmCGbJ04kxgwQEfGPvWHYnHpjm2cw0
n29FnrPUCkIo+N5y1je61Uy5DVYZg+TfW9mK+mXNB/mOgj73yb9lBxyGNAfAvSn+
gs02l3vVtSqWYiLzzF579JhjBqwj4sQirDFxsCHMJMnvDlcFAIpOP6iUGoXfbust
qBfBGhBrrszHG0ncejnQHAQIgMCwKBy24UAofcHpkLFMyh54QSUQyqhJsSGhbtCp
Lble1KqRpKMinkRlL45jIy9r0yqTA3/GJ4A8i+lMEP+7HQVu96fljZEgduCECCzt
Z2EMTbf46nBenQ2TEloDHTavJtyxv6YCiQhjjtAcWwpKicLIg1LMr8l360Uenktb
Z7EAnuzltZDbBJgjbbVmedtdnz545EYl/R7VivgSrGlTZq+AiC3eKTDyTaFvg1Tx
lBwTQk3ID/zsTsOP5eX+bp44C5Jxqqxih0m8Rkf+o9P5n0PGpt4mnbFrn9P/qW5+
AFM9VRvYJmxm9bFkvHIjFGpdtjfAiWsqsxiMCFsyx2MEQtzaeq39oXVO+LClMtOD
dh7uuAqkJeJBVIVO78j44cHqI46j7FdPS68TeBe2FbMpNlmcrK32xoH752sDK1jB
WO03r0qyu8y2s21APpKizB7eSImokLKzGvJL7Vrie97YCzbl2UXT9lADfgxeQMAz
ySHKZ5RGbaQUh5t6Q7nrhTuvoIm57JUFx9SaJHmcnzjP91LmU4PD4gOyosVmHfwJ
oyyNWMM9PwRS8ZEzUXTpnBngcuGR5WmNfiLxk7vNTRUO205H5yOrA86lnCQQ64+W
iKqsdissPB1fkPM2Mk1+kvZ3stPVbrSJs8SfItiVr8Q2I08a9xAb7fm3EOqkSns3
U6ZTdm05DHGAdvYCd/ypDDVmNSmtrE+j/OtUCsCBvX/mBkWpifqto6B1361glUuL
xMCx/7s5wsPawg0da19fpknihNMOhIwE9rujR5RxnucuVU+Jn4RQEr7fD5M7Dkdb
MbNzrB2wY4BqCMR2pZXS+3WQ/I8jenSnsnj+JLsYF1hyUAXeLzhdIzUIn0gQv1Kr
rWd/iDSAouK3+QfX2SkkKW4Hyv6cJ3Na6www6pvkMkh/4kIdjUNZ0d1VU89anX3z
z0v2rGJsEw0+NP1iWsReGnnoy2Zh3kHytpuJFjEHLpBOOFCSZ+NUtgtsRrtJ/Ih6
QsWful0W8GOQ7g7jZECzmwS25Vw/YmdGO25PdZ6w2jVdRFUFa52FXron2NnymByP
UijXmZ7yKbLWPAMswxUDKtV840Zwi0ZaWyVBG6KpRwQw/oMBBfXWQzYEX9lHFJlq
AF/7Qtdo7h2/Sej4VL8dk7jKAmhArGD0dZGAcxZiLz01p+o0VIWR5VFO9hNueO+/
9WBifI9c4giIGfaEPWCFdZWNflIYdR7c6M9Jtsw3kDngVXBWy8C6tv7UuvVe29O3
InpnC23NBC15uoc+TP9QEOQfVwG+u+aGyT7M0HCPsQutSTHFDt6NcET7CW79n25E
Jwqmb/8nYH0hlOnFfouG3wUHLwr0ZqBv9tIt6ESUICO7xT0fEYPmt7iinX9bYlZ2
5l/7qFV0z7x7F29VFLTz5RBumGtBD6YCN33ggurwGHz1uzRZ0hc57fs7i+Qipquj
OyZbazqHsTzSB15dyfpiK40F7G20mttf/hvCw9H/JykGuTNVdX0ZSOb1En7QGR4h
v3bWv1+vYZ8H4ChafqOvflL9c7PQ9VzXkK0Yx/d7g6OLG/yfyzEF7+MHKZ8ZXSW5
lPpmZsXMStSnga8+MqpKNmnsHl14m/E6nhF2xzpIKn9CypiIHzUB6NRvBGMGadqD
Gl8PQr5OU0o1KcIGWxAdHjQJGTaFAr4ce5vSK6i39ToZ9eJrQQJmULMfP5YEHS2h
YZLcAVCtZQNgoTrbNGhR8Fw3dI/hh60Posotjts4etfpFdhXmIX+Gh/o7QoaeeT3
TAKIWR8kdoRGoVgEcIU0xQLNK9AJ8ly5Z4WAZmF/QuKou5KZ0t36ifidB8vq5Aiu
mkgfe6lA94NwD9CmjyvRRi4cBdAeNkMa1AMR1ErtNWogVMvmwa343Tiy5ViQsByo
oXCf86cQX3JVclktCQk09p85fISrnok9kLV4e3FPsYID/lbJXwx4MTa8o1dKiyNo
oFYxqQHmj3uar6QM+wrOzw4pJOfInPYQj8JscgQdYFDfpX878APyu688PQHOj+6r
ow8atGwxRfb3mzn1ARXSVSXiJQ1DtetUp5RIloPaIpiOY/tmlhh1g/oRAx0loWCd
MMcMTBBfCiErqx4yYFhxQ7uTxR/t5dpTfeKpIMHLsRNlz7/lYpNZZS/YQQ1Qx4ln
xo63rTwHN/NsNOSw8uXp27JRcKV88jqnlQuimPttDRDq33Yhisw1qam2jZWNuDJo
jWAaZMvx1JiUZhVFrfuI06hAQCNDLnb9TtkRMda/PEdro9IwHe0TBCKuKhy6FxVv
f3az9ZvpO6M1MIzu7mUViH0EQLWju3qiP1jYEmmPEkc4j9HNQPqVzfXQcnc4P5KJ
8zjZh2T9XF7yhEOIZfYzJqhD/EidS8l/17i8cOQLzEJo6DRlBv67dZG5qqdgFYNt
s3bvrcpQVh9GGw8H05CU7Oj/QMRcE6Q3UmeL0S4mXl0r+SrZSJl2iiCtJn7B5QWf
KXhz2lSv3fJRTBze4ByKu4+H9oqGfCi2FRFgc0AnA0UpcgOEbdEC8wOuYMIXMYX5
9YhznIBJr3kBzCI9mrmYDO9g1O8fIwaG617SCvKYq6ltKpVz0YcQGoxuJ1+bqSPC
u1op0rZo5dXzEaMyfKYgOc2eE+QhvXUgrJsKzNQFFLGI5q+BZhvnl/V3qqHXNlKV
SMPPj48tA4lP6Cm6qC25r2+Tjx1dpJGgf317kKqnUPq4o7FtWg0XQrRYxyy//BCX
R8WAGEOvrrfEpPf6FjnYc3IyPgvg4PcMIUglvEFRE2/MZTWNr0CRAqNAAsPYymmk
68Wnk1htLf2ZZ5er63K2srGjJshs8A2iXchuJxCR2DLYI/+T7OTeTnLQ6bhSqt+i
bgJCekVhawuWagcshFZIRGS2SNYf9C0JNOU9UDN4cqGLfSE1NHMuha8BKXkhQVWJ
5bbcF+RTO01q/Odl5SRblXZ5NPw88g3Fcr18wup7F0/6rBmgQj1772k0ndV2FV+E
GegHXIYNvf4NlC7u+KAWMUbRtp0h2qsgIcntn8p0erzftjWjiO3/C+LQb95LcGU9
94sDcQ47JB81Zqx6hiQ0VVL3H7GpCa5LViXQZ9wtraDL3xU1T2j0zJ8MnDBfOI2w
bZVn/lCQOXm4fWfwzHV/qdVn3EK6lX0c7+eZvGsXx0c18Fa1YCop7bhoUaTsgRJz
gcgxwk7j8QM7r5VJfgsF6mwhncglJVHLOdzr7ZUPtPMINdP6wN1UVq0APNEEexGk
CRs92ZWNDT7cjC0ovNX+rux0j9dHD92l2ViqMnDxIz306FzoJSSq9/OnHw4XKwbM
ELPIT6JMvm38VAfIbYilUmygmqPxGovXVTHmuVprWFG1NlFn1Ar3e2NpO19iuuZO
dBYydIAjwzijkV+XiIuNMYtydZrjFrtBQVBj4D7iBCPq1so5zaNyrZv5fytlOPUc
uVP4BJn69OWXoApkDg2oTcqNkYM4gkyG3bCD6hIqRykKug+3qVETIc8N7aAMrnbr
racwS5jdYgHnJgieMuk6cb98AhhDSL7wKfMdkU7CG+nwxCHAMTnIPKCjc87u6Gh2
GQpEk6y9hbDYtCJgFa/k89Rmml2kMR24kR5b1EcO0cBial8MdZMk//BVyEwXvGOI
4wSdNZ9wOoR25g647IXGozrcnI5qZxgbBJwJpVlG1pWMRUnZHSrxTzpBcoSZNRZN
QKse/SHTxCuoPDGbmYv+aqG7ejr/ixoxK+aG3zYPAaaQ1XjUeYApINC0tjjyfE28
zbOdlVOtR5xoHCJj4iOhq9paQtprh0Np8PSr8XOvvCIdAsJPSeCmOZvlXKDwAZ3R
zEzxI/sBsba7wR2n8EetCn7bBM84QIv8WXa+i8ktdj9WkenUTbKSIHcGCznEo44x
TzjHOaOTvwiRdspBkPPAD7C1hNlf273Ns4/E7+fvmKQU+YH4p8+kosEco+w2QlDW
XzPqgGCLI6fhC5xpwjaxMH3M+iKwJXysSVFqgUVFVLwAnmoR3G2YJIBCPVXfLI2H
yU62e3wR7PucEHt63F6DJ8OtvH4zZVYJQIcBo/AECGo+KeltHtf0yQWM6AFr4zVv
eKfUdTgomWHrbf6MxAurRWWX8tGfYu1xGDHBsT8D5+/p1mQnhBBo2tv5F0fW95QA
+WqziBNmbjKgXEOK0r5bJdxXfYvmWuJCGmwE+TzDppesiUg3oaJvfRw1cwJ3GTsL
ko89qy8mTWwxHGG4ipfuVLU5rvmpxO+pvKkKhiGtmF8fcRXU5bqz2JCIcegqdaqQ
mJmh8rICNT9mtiQseSmFiJsIriVjYKdB2n6u0ryD4PS8LAjk/68V7C+Qhfm4lNrK
311WYHUJ+jhGK7RlffcnLh6SwuWG0zSFuKerlLhR+8zH+U0AsB0xsvK6Kwxq0Xxe
a2EJ4TKvnfSFXcQTK0LVlW0NpwdG0CZD0IQH71H9p6eElQqKO/LMLyoMgcw1K9Wm
X60c1/GgD/UvTRaMqZ4Muq0QK8mGfwTA5zOKDNflBAlG0mc1FEc2UWpAbYfpwfSg
y5QwVbgvTTeJ/evWNULLN/YRfb2720+D/tXyQgN8CkpBEjwQLX7WXErkHCev4XOo
LTXXQIhvpKDJ4NaSG/7J4CfhA3qvfCir5xSBn6LQBYjaql5VYtApOcMdk4bL1RQm
SCsx11ALtgpve2T0wux0iHFoq2Xgqljg9TtqfRRu8e8Lga97thAvIQKXSVAvYpbB
ojkkDtghoT0UrXdOvprgt9gnbRY6zvVdTxaqFZZYkK6SGnD2hujsoIV5MsA4QBcI
tCgjiHupVI9CP5qsCVNVZ45oDhQqkyZxZ3fn82oo3UkCI0sQkh/FNtjvkg9NC/lp
H3fZ7YVBwndoRQnFEkk0pTDfiBVDTev2gVtwuSPN+Gvblf9pUu9fWnBjc0KQiYS4
H3di4br8gPdpaZN5P7EtZSy9dUt51EoxxEA34DYUMv/JaFvbQCm3dirTlhsWrPXT
f6rk8f2EJv79Cyta3+/kiy6cI9BS85NCM3M+gySYuYod1Own7GQqpor3PS5LnjWr
aux6/2vSVKg6hNKMGXGuCKXXxuC5gKaaH7hduwnTe0+h8rVZ08rKcheTdRKVi8hR
Bv2MQUz66O2F0HsFsPPasH1PLrbA7XlIpyLajpBxZVSJbws8Olp9NCYfDqgRAaUb
rQVjNcgYxKgzr+PvNRAgUPi5v2Fwxz5iUpdniQaT/6Cw0+pqi/+pAiE8oDNEcj7c
Yg3Klwr1UDWVz5VHzxF98XmLzp4VEhZj0TU04LcR30y8b8RK8/Rwgl3UJT5gluKq
gU6TXeCt26ha3WrTQIcx5xksvxBMwBu9pwARG1iZwHpfNEUFMWm8ocCZXZcVeguj
iKy5KoWGI6xdlTSTUGN3iU8PIIhOB+eUDdGV4tzmgC6mcqD1qW1xOgGPm6ZrwCyX
YwWTI4HHaMcFmbH1UcHDoSRTNPlSxuJpls77p3CkC1Bhg9a7cd/ZXBEOfR6IC/dt
zcDcciBFPqaRZKg47nsaAh4OjSiMNTNDw/J6u6gSGLEFjoVTABrYKsR5bsksf1nT
Ooz0WS78mPR8dVXHRjANzsJfX2r3REGXej0E/2iF9EW+uvouAgQFUvteONzUfP2i
VoZd3NS/2dHtDVvHeOqedG/aV6olzArvqJgNt8j6QSWCfF23z1X/1SMJeg9sOyt3
xIywnBUHghg+H+4sFGIIm2bQziRbeJIcTL1C8jSA1PAGctQnk4v+srnJGmsdCTfA
TntJQeelFdi+DMtiuwWOABQZk3vNyNKg5x8BgbRJuxkCNTv5q9CnSqWtdq+IDW40
s1PCPGzlqmS5TbltVZ/QfDi/Y3JJMZaCZrniRvKR0E9bTQszbmfRy41DzjnMuZJM
KJkYVzkx670hs4kpbNwfgjxV/yoXWnFgq5XPvn9sGq/RcqJ0OP/jFQG3c/W8VjHk
v8Za3loQledI7NpYnUr5PY2RZkQb0cqStp98ATeYNnb3ia8hxVBobkQaXH3FF1gZ
mYXpJlahJqsKm8PyRPze8Tz2entjgMBwYRl0dmSxMay3KJkbx9n3QlOwdwRypRkO
NYrpbzSHlLhXnyZH/iiHcKhVEHynItrNG+LlF/aiK6EzNTdYPsRNP3U4iTDL6XvA
GnC+Svjza552vbAs6Km3c1oVY0VRG/GhGpMNbq5urKQbp/7uOR4T+qgckGb177Z+
wWGfsmukffeWvlkxDvyoSJMnDPdhg9pPXN4az0gl7gqWDSexSKcyiUs5S8VLvRfy
Ibuy1Z9qF/0zj+9KK5it6j7fcUba34M4YATxtPuLwJFKY1J2TsTz9g3H0zP/NCFB
tx4RBfktzYyoSC8PmVDQ0mUSwYEBrz2Hz8c5KO6Zgb+NRTYjgRWbnmNhUJNm5CM0
wlBilACMotAT9SlKsLvOTAM2aD4E0wFBz0Z0vINmrSG3jSD2JIe1jHpZTkn+A7Mt
VJXJQZywnxu+iS+BJ5t8qmhQbeqbYg10izJX9NSibEo7Ohf09L373Zl4kiPo94Pf
QOPFTTG0rqCf7Bewgwwy2NLAlPtKO9Qp+qX2Munpfi+oBgVrZZqb7Ewy1VmdSj8J
38uYoQ9RAIiKTRSGHtWcrLVs6q5e5FJLGoRbxMkB74B7Bn4zlIiZc3dJGzcYcdDF
AIF49KdSk9pE3KtI0xVWEI/uCXs7wTZWSKOd1CNq/5wHAG6Hiq9ooo3J/6Q5aA/f
0hFqdWTjhrXdiaeZguxBMFIjYIiH+345WIZdEFbpfJ5EweDgKxf9Q9t6kI2lM6M4
xHi2dTw4CnHnsjXLwQmi6bitbh6hC7KDciiWvdsYPYQ9Bb+QgdZrHOqyiwSYruqW
Bj7E4fY190cxasIdvwx6cKN8Y8e9eHVEy7BTTMbX/wbo5fm99GMyaK1T7px2Z9KL
INjy+M00ViNQ1SeCJPBidCflxIdfBEBqE1rGNR32kSlTlcNbyBGvYmx3C6YEqCu7
ooxha6ypB+oIc5A3uNqn8KzB179IKWz3aa9mW9dtKL+6x178L1jH4RVGuuB1ewGY
U8CKlnu614UffQE7l44LXFmcAKtvjErKZ4Gf23H5RQWf5gTJNtCujdksz5BK0Oi+
jPBzLwwVhLe1rlxXv2B+b1yjtpUle1jkWT/HQC6TqlwM7c50qqrsSSo2ijwzhRfu
Ny4a6m0/tRWeyI8FFDXBYPQOT+v1Q+BBonnFy7rFLk0Cv+a7RfZ55VwdqL+qId+V
ze9MxL02vLcJUFBISU+zSO3TsILD2WVrDpl0dcr3bO2T0ABRhgwX17maz8CGX5Mp
bd0yX6dEbcYIljBXhg4Au29fG2pQudmN3AgHPopenRIAXalxZkDIQ9OVvDvuO1SU
GDzMjcinPyyJjsDRH22jPKCt1v3IyUp5EimjNLZ/2Q0npVaM0lC1AYBzp0OTuwnz
qlILbGbzwn587nYN6rouqfwZNq544NqMRbHt+rkbs7fuzC4cL+c0AAWhxFqH/0ir
S+/1R72/CVqw9opLkS0DGWuLjXsa098fUG0n1fPitYoB2t0Lg7jiOYPEfzOy188q
0CstyIC4U2jyLy/ZA+mhH2yg9nZoIIEITiBi1PG0QiX6H9b7wiUDmhUf4cvRLgyN
ehMqPlAXt5pifXRIxqbWrfMbhudOhIW4VoW/khpFg4bwW20u/rDJ1B/dcHrPQQJf
i/dieDntxu02IxbxUmOLkf0qL7arW7AkQJNcdprztoXV+MRfTQ8usPfdRkgohqfk
ZrxgMXUFa5tQgeV21Hp9xrw+gMtSliYiFyMYeqJ0n6ekE3V+FlE16zH0pGYrAV4j
7pgyiQ18b3EAAvha6ziZmEh31omtL9FcysIUu6X61ijQe67vWjy1/GQPQ5j/1bJW
PBQEKDHy7K4ieldV9tgBw2Wvf3PBPEOjLVbscDBYwBtLoKHr9ZXUXdRWQemHNmlt
688V+S1ZP129/pQg73rkumMKPOmSsulA+zICTo7QZ95eUGV2zgyaMzeU3OEhqKn9
cDm41yS8shtUn0Igit7ampz+u2TESy8UQJtvioKhsAQhVtrS0ukRaBaReTc77uzs
Yk3ka5Y1NYjWDJuw5x5GoJF2mRIFm87RwnEDsaXlNoJJ867s1FBs11zVnL8wzKXu
MZZ01bSnv4A76QbB1jwJOzRW4bPoHkQLx9tHYjnBbykgTJMAK6akVePUs3kPYvLe
fTOUE01Pe1lnlkShjnt3+KHk9VUBobDZ4bmcRswA5Wwsn7Ws+ExBD5nDooZ7nLMJ
vNqq1wZvHM/Q7j4+hoLCb6UXhjJbFm9Mf2WfgVchOqTQabhPnnw3seBFSbfmqC+T
XiyKA5Kkfwwqi7BniOoaEBMUxAm1aeuYeqwga2TRIv0auGj5vW7hPY59lKSNC/Xo
jlgBVYmrpQ7FsKCtgksPUMDtYotfZQh5pArT66/p5acmHL1ChEevBFZ8aKYwuNcf
Aq4W47eZ+VJp5nFIXGkM68w3ccvB5z34r8YUuZB1U1yig1w/Ka+7PMSR96nHDpko
3QnvhA3izN08XqVZiFrZsYcULZRfyUgaGkoH+hHLY1g2S0h4TaaBBygl2BItciCD
rX+UeTNy3g/MZtlpiYPpHPxo06stX95+KkMKan5PA349S7brwH9A8c0WigMazJTt
ezhvp9lpP4DhgLeplVfz/M0Ev1tspdH1pLH675y7XArbqZIaon1Qw8FBNfUb9A12
Kg9w7zubTK/PfIHg1nscIIfxl+lk+/DVL74WOgOHl9MTKOZ1l1RBIs30tvPzLlH4
hCZ6NdzNdEY7Vk9RxTNIFVOAFpZ4KyLo2sKSU+5m6VJBpMbCMVnsO/onGtx2Nsrj
bv/xYDYCGdovXXFjHtiBpvwGzRzKZ4T0N8fCLLdh1xDRRlg2z0jx1N0gNfDKRXag
501tV/Jb+l6n2IhctCcTPxhs9PCdQEJIoxumUj5KUwlptKLVvncA0oLOefa7OcHl
coqGCZRwmTYMdpsZmLq8ik4k/nvzb8JOuwJhNQFdgkyCZ33VLolwD7Jd10jQ+toZ
mln5fBIrGALU8fp9eZP5UX8aaMlaqXr2CAFYjPA+2g9lZfYNiQgvfrcg3whA8K9e
jDPBkfk1BV8nu7ykbr9UXcZd51+2uSu6bEGYUvIrqX873Cc9lINy+CSMxHgeiIgT
KxS43QtiHVLbnMTeqq9+I6cK76+dQufvLPSyvI1Z5myw8NsIWziIzWnFPqYiYYLM
eavYvrG/1qDMCpfNKQciU1l6trLpVFaazqmusLQBKzax2GHSvZuX5YBEqVDJSTIE
bJxYpjwBaUjh0JqgzTP6Dfkg0pPT+Lk+eB8Do5rgMgRsDjMyfuFoBsVtLZeWvNHU
Y7MlfWG2uw14dGTnBz932APfekrEZ/7Y3YZ9XvPa1nwUX7y3fFLTCpqs085+sQxm
QkJOPxcvBXF2YjK/0CElP8lQQJOuJEUaS7a/YIfZBzWtj5rQHMNnN87pOko+cw3N
EFe24GSfYmSROKEE6xGelO7LybE6mVrA2cJnu5IDFsAhNeE/79fvAqAidGx/q6yI
eD1r8Cz9fTZC4uJfhL80tdLuOJWYK61rnj7OMQYAbPbzkVkprkoIORuSy37Yliw6
mWproVkoYacisjiLuSokABohuj/lDiHc3wthaE3H3VCSxXRYkYajHiuErpVREY7O
2fQjiLM22jP80lK2ScKkbWxbrJVGZoPOwyC97Tnommw32dB4D710pIBV/KScQ7Kt
Qv5rlDhhgqrjRLbuXshL6rGipwsvB6mBZ9Ru9lyzhWLNB48lUmNz/MfkZaKQVRFe
NK5KZOmlgcOWibU2lc65xAYYYedqJ4QgFWxj9UdJ6VNDxHrentTCi7sbTeYKAkPF
8asxdqhjfr1V4N3LU6A+5N5unjU1NT31dJq1mk1MzyLwyuq+qfK3yS5wlVLYDTAE
OeSKqPqz9YEflmGQbE+lggga3n+uDIU/CR2RJzo1kbS+7nqbihX+GH9iC5Mx7ZTU
sLCtQaoSM2XW3dc7aBkUf1PrBZuC7tmP/WiB/cQbG44o3JSJ15g7eXPLW/sSBAxn
ufm0t/C3s64Qy3ODhShocCvQuzW47LPkG7o7J0Cm2lJMsInn3h+FR9xaPBsOeXEG
EdOEx4tmfhHVpJjGwtvlgtvS73wmq+KEgwPtTJXuFV2yXpzY4/9r2kBdxBgkzmUU
TRsQY8HMDOaHZFtRIUUMlUCO/2cPWCASHSbn6X5ZV3ntG4KxWnc6VRK7WPPAInyu
H7+Opn2GMvKv/c2eOk/yjw47NZ0UIuYAdXvLDf/IzfBZynVN2tIAy1U1B4Tgk8Mx
3jT/b0HJSn0Vdk8wY+qoJDZSSGzqAAUb/HflQAQaC2kc/r7r/tCuETpD2QBGCBb4
AVMGO/ANY3PhLdHkopON4tQLJGMS0kKvgKMvLO9mF6OuMMXYbZVHJYAo0/s6K1pW
78MalZv9MK12RiHawsgglfOJ/OhLlFIIhsDstWkM5sJETfz4jEEYpJPXsQI3CqON
5R/ordoJtN3S5lx5jE68FPZLKOlrD9l8lgqGshvgLSjpgsaYihFPSSGyw6/ICmXE
zl0vtr71seLyzW91IcsAfCmpveU/FLdnMjuqRk1lyLqQN3SAmBxxn76YfBbWnBH0
2WvTGsv9ad1NQgrbP1wdVj7MEkxv92FYYMA/WmXmPE+Qg8tIxJE4fGfjstxqWLLp
BYU+GbYflUJfgBzgjfivQ9WuIy562JjJqCWBcz+9lJ0DP8ETUtsmfK4tv0TJU2cq
VJJaCemIAPOPhmK9QUYUiFWgkhs/lSCN+1jBI4OGVTtVBLmqq2QkC+euIqLM6MKm
QNyKsaGAkTw220e8uQRNpOey+HrSkUxP1IgyLGWQ5zaXi+jWeK3bbD2UYy1BaZtO
78BXkrLHtgOGdk5Tdqvv6buV9tXi5spRje1vnw7HGpNZ7JVcOjg2fnw3ELo5kT0M
4bW95/G3JYOJljKDy2z+5RSQVfGmpzq3hxy5/AtGYPb5p9yb7xxs4XfcMT/3Jfd/
GMk6bclPHmZrUgzvoZi15aq13ubYEUJ0VpcTBVk3YaUbJCxHTPo6b8y/w2Kp0SmH
D1MDl2TsX2E5CzEGjyV4XMNehyHHkDthP5hZueCV86sqLIBA1l5xOxPgUV2fQ3l+
HEOyMKHqSpeAiy15D3if2Ts+WXgEXHb4YT2+Sl6hWRD+RJLn0FLckCxVElD7ab/2
GdyoEYq416qLzg2ET0vkMbQ9VSVXW9gM0VxkXnYG2pKqJQXRyfEi3Ha7T9WgslP1
WiqFATXW1e9HOu8ncSXCEyFE/88/i4TlUY6hAXMg+JSRi+FQp/88RjWMY2hEcOkd
8c5MW2/Nn905QdBAg8ZC/y6/x58GsoUmQuV/Gfjin/SNsj1NdMigpDriPZVtXx8r
YBVjxCiBSsgrviwgsEzoxBSxil2OiOMqPs+vYJ8g2r5xhieVly7V14XEE3lpcsdm
rQ4FG09l+c5uov47XwN18Qceu+nGbapJWZ1XhjM/vQlqJ2W/uScOK+IuCPRrkaJq
QI2fgHFk7j9gSfEOb4pmGGcjC1NI9olyZr64HayWWFGFZKgDrH1iAUAS/qqVye9j
JYLgRh7fsxL7rnDISjj1Km6LZWwPzTuy8L2ykwlWXAIkyN645PXxF3x6xminSgop
8FFAAb7wadFdjCJXJ/v7mZPr51Y0j6viNjCe1JBIaqY8lzjEgXyH9xN0p45mNlwK
eTiTR5LEcqwFLAGZHuNTIwFFMBn2DhinNYzIeFA42TT4Mn1pEFnIElRijnC+DOPx
429fYx7psrnbUSo51UjgX4U5AXGj1S8/h9tcp9fqq7YPBQN8cLqfMveXrmAZ3lzp
KwUFNfer3CTrim77gbXJ7TBC/x6VzbBEONfTaJk94YiRKRzEz+caun+0Nnur2a/J
ACNnMw3Iyz3xEKzH40uaLFt5QH/yb9tXkeOG2vhTF4lYq3dZeeYOZ0nHggy6ld8V
z27GGaojGQ1MkLiJpHyqQT3aGEmEg6neUqy3twuGf2LUc8V5Uc+TRBN/b5fQWBvt
Bz5TwqCtJdz+KNwxAkGZa/50+HjU09GwWeUqKIQX2vEzdISS4a6fGOPUFS7y4ukl
XJfIkdXavXQUdNlH1a8xKLJ7P0nZdqKQtoEU9VMfofK4L/RD8NBZxCXnZEE49eHA
NdspC+lQN1zcO9qpzsLZ8MitpMNlEimOjg564941sPUiABtdJAYRPTSe01iRdhT3
ReGG1Qb3HTMbNGzvhAMrmZzakOCEkBFi7E72uUKxICWSj7HMnCDZTzLRoUm3G3yM
kqWbD0up/PLZJ3PF0G5Gze762s8SP2aVs1mtiDCDXLtasjzfa/84nCQuhylFqfxE
u+hf7RegaitMvpllpX8EpqiK/ruMc5hoY/xZHaCabUSMvxpnBepKQWm2HG0IASx+
9b54WB5d5bSzKI2CfIcczl75vvq5HIxmuoX9hioxgbpLxnsyczjMhUfiXdigCb7c
Jekp8UfuJN0R6mUiciJdMSCNQBxid/UIdPleN3cvRnlW/KXXrqv1R+ZjADOppZoS
aSADHJR+dA9eyxjDqDpZ3SpWYUatCP5IAek5i6pVMQs2QalBl5gpLrMutxEz3F7p
Y1JO3HJx8WsNLjIIJVIRqBWZRF6kF7WXPVP027ZAmWK+YwOzu36niykbhdXkqSyE
O72+SqLEUyk015EK+5RKRRqr+58HDXu0Cl4vBMH0qRbtteItMYTeDKP4m5MkMs8a
9pBdKBgE1MFspY5jpGYSEqurRv3FDzKluQsnCTBUOaK9CCcmFyRfY0OgDWBeHUjN
0C7w7d3jrvXcpxdqeR2ie7Dj2IxywAM9PM2yEZ/WvBSxQT8v1iNmn6QJb1b2SytO
NAXqDQ+/DZ6sMzkub75PA7HMibbkGKujtB1quc/QZ3yIyMrFHvtQ9o9F0hSxm93c
gL1ctZZQNRib6Zqv/oW2nybdd8HfHBon46ZiqI0PYlKnqz0lTsRlYRQjagdX0n4J
Mk3it4NaeSc4s6FQz3JgDl/q+7CswLGURz/t0Ex4y3hqvHulCBNnd9Qr3nm/umIG
YBYvMjI3F4MU3SygjhxM5KbSmAKMi+UdC6RMfjCoDW1ClAJTJb3VtTYkLeYJIeTx
Y1FAiqBBSS3D6k5UYa5uQBATSeI7Ae4gYttS0FkEXFRyuWbf/Ha1qi9WkkQfG5RV
ikBfS6+WvYkaF2NGDz+AkcXb5FUqVM4R0o9VIG+F463UEGjLK0KNeyVpi0v3pOrZ
bI3eU123hU+1aSpSrK9OfgrnenCf0ZeZ7NOk7hJ95gDOXsaWRJlQOl++SJXpMPKM
1w+Wzk4VL7osHujT9MHx8F56wHy7zS8R/+Sd/9SA5MDFoH50osVJembTQIp6h/7T
tTG4iQJkSvt+hTmGl1XT9+Gx62poIPaQ5K7pQ5J7XhfFSKwGNMEUlqgB11TXjfZK
OggnKN/pppBRtruFcWW3SZTxjIKGSj4j/kn+ZKc4Fg73YV7h2xRaQ+FoqU8VwnRh
KpSWkmeASM1Hd1sQVbbSA7TU9CbktgmR/DG8pU9e0VO2SY+hLS13I7GunAvy/Bv4
lm4Vlbx98c/Ix7CbmnO0cCGfr9TRLfC1iCcC6KGj8bmUSKwz6518r6mDtG/J7bk1
C0cCI+9EyDuhV6/dSDSaz2H2I3oovO5qK3LgNtjOc063iCtL/i/vQpTSJ6Y8RoS8
IxReKGC+SIoD/ioNXRRAskKjSFReXrp0INVwBiZud+1K1F8jRJH8ZDJ91Ep3ztUr
9lSF1fSG2tZj7qhztrgu4CbPVs1stZJfBFe72SriNowL9k7cGOaveuE9EM4kiJqQ
u71J/jDBm5nV+uqAUMCqikXmDfYL2yx+3PWOhPVbPrpm/LOPmMFtp6SGZ6x+je72
+O1zOP2o34N6OoFXmz5kLEZPhP68Ra/3ZM6r73sKxM2Ub78bM55CABHlpYf2kCTm
TdLAWqGv4VrA36X4hSpiNS4Lt9AWJwlvXVFNurBOhwi2NdZ3RxLMTNmOXoicbSLW
T+CHEO2kQAZ4DYNJXKdGsWvQlstrXagq7fQXF7teocg/bX5mjeV+ARhsdsa0BwbF
gGqj3P7Sh3Gd66LAjPPQz0KNu1O+cg3c7p94ubnPdHhxm0WO2r1QC0FTKiEA50L7
cLUf+9M8WoXGT9w+XLDWSSqM3zeGhlQP+Cgt9F/xhYYG67E5MiKNO+8EYpGxZBcO
voH8CwRbeaSTeFX/QS9O+qqzJ19QsAzwR2ElKRvomhyRYxJwUvfUXGlMp+IN6dDw
7S7AuREe1oE1poNF/zoTmvuVmvEs1KJcuLVKBkXIldkg4WSL1LjoU5d8832ix59K
NVLlcwfLdoIfqtC+iN2jd1Dd2803E5AeHz2uOiZRduv0oWDkjpyWeystEuUo8/Vu
efC7+betK6003/1NhNYyOIl8APpjRjjOhGmIF2YM9vTduq3syipb0jGxMgMjiEwr
YZOwamdoQKbpEumy3v/JcAIj7kah2MLuBHAxQ1Kb165SO2ivB6lgdLD/VJkllcSL
UYMIGMcT1PJN+NIfzVVxyV1bnd/qeAW/1Ue/F9TsgTzTVRu2C6+6K16egQHU9w0I
bacaLbjiEvd8pviYrobkfUSl2pX4GYadaaS2OovVkxtZmtxQZN7U9rhD1kqweWIw
5J5/YWD6GXrJuWlsuH77yKx8mnZXAKOGu2oTN8hfdeKoado1baVBrllS8fmAaT4X
XG7G66PfGIP9K0Ig8N2U0zKwul7f82ocBWR8xHXlTcW8WgdDlfkdVBJKanjp7SU1
qVtsFsBbeyz9FI4QIDKgU9zBPAUX0fThKHUysxVeBd2txr9MO99wq05eWqHgxm/X
pVw0OjFfQw77HRHDkjxe41TQberBnHCFUaOuF72lUmL8Ea4/REBhwXSyxgheOGSu
lPsB7Y4QCaZqK+/du9KNm2KBwqzwoPAebwf2uDKNJWx6jSUbcCEJGLouuz6wqoEF
X3V+g+cOOsiCtwUmPcDsy+u/zovsyv7ULhmfroa2BiPqXwCwapumBvWDDIdjsVtZ
ziLn5pZwpAYky6yzFigfSWW97U4SoQEuYgwLVHaRQ4oxsgMRhb4J5eAyDMQNqWEH
QaVArlrFDqlgmVkQUITH7oK2cyFESB3U5YNKIc+Ha4v9mki4S1FsZIPZs0hQK496
YwHC8JDLGlIoTU8a+9AQ0Neg0AX0/iQ6bexA1KjaqVsQoQRGQe4GPx4M9NiTdUfp
5qVCvSHPJiDWq4Viw4NQ4a2n8ygOtvkITah8VrmCNuhuXPSegiccGPRxCQESo5i6
cBXI/QKX2iHBPZc5RpkZ4yOURalxA5t7Ymvcf0JcCwQyqu6hWcfOoir+C0FsTlfQ
UhUG/vsdUVSaMwxVUFgY1if+2YK+flEU0mWZZSHi2pqcPuZDkuX5qG0T4n///y7w
nrb33ce/YTS2wzBiuUfI4orEnUEtAb1me7O+M1NtAdEnUucd9RaO4Pm0eZEpgyCp
GXfRbhy7BuuisIc0diq7Q4Hd8/FVMk3Xp1X+YB1i6mpmkwYSHzb5kaAjm96i9yqR
6x0kwl6/tDfkAlo/uKLb9Jbi1Y3G8CYodAiwOrDcQ9e4FEt5nXzpSL9KhreHWrDb
lo0NQzmesFJiBIgArywR0FYbUY1DuBRwhgsZpT37CoOaUPbJTtqA4KKJK/czkJ6d
C86FxykAdddLLRNUqi7/kjeboSRFWf0ybO3HnajVx4WlLiOyMR26TDDWMBs2ZTGO
xXl+Kg3lyYDVSlK2Fc6lUqOQztfeuEzdC2CBVDn+K7543HoEq6Zv0Iq4Bda9v7aC
ImDiezgI5wNLyvEgCOOJhm1mWsUYqX1DaWgxS3H3NeQHfbj29uXXNUrJsDcE9nDb
JKat2TJr5PPrEAguAY5ag7/maeUy83sICRls/zd+vbnk314pXwSGruCEuNp4s9de
ckyIBkAyGh8OHxI+i1sNi2B2GvZH2SQ0G4CtYP0mY1e0QKLhV3tbx73KrXtoMVZ4
MicniBmY1vg2Tu4spDhHyKzb+vL5SmYpizIi3UiVyVkXnknDG3s5BrOY8zGzzVQs
Cex4YyZ+5CCauUEybOyRuoTMV3Zeo94ZAjjDjSnZeAgv5T3wba9WCTJmQ3Uqfdcg
d1sWGg+QL4eF53/N5Hl9UYXjEcj+7r0CMUqdsuIC4qyyscnP6BqGsDH3EGY6DPgZ
MmTK3Yycnkg0RcVtHQd6KSxYUtmoDrn4sh5zyZbYz8pgmLIxYT8usy+sCOx6c5hS
Smpgo8ulN7h1moLWSk3Pz8Zh8+nWoC+SCnPyymABGvEJgMLvNeWU9QE6+OZRzQBW
ZLuRCGFsowDxfvfCK88c+8U9kaYjpBZHF+CHg6FuQG6TbxxONegnohcheV2X4NNo
gvYitYFYQ5AGbgItUUDm+ZA2zg0bUJGjj9khInNtKyIJjhG9Yq9rNzX2n4N2Rr0w
/xo6hPGKRcp6pKyfUQQlBOOCV2ogWLfMTQYHadzNos5rlNizsyJ7HGxk7seygVwh
DO4FITIKsEZZmw+XmlVRej8z7WBTtkSEmPodD0yGzQR9oDMjAUFo8Ie1xZeYyUnI
YRRaoRh4z/+EHtu071B1W6Q7yIIoobORgPEC3sWLjHquQYQMc8u06p70rvK/IbHu
gxpJoU7K9y2mvW4XZ3ijUPg6qjj18RLVc3r9wLErzWzn+ciKdlsmTZWQUdMp0cZ9
YbQi4pTiVfEJdVvOxbUq6NA9Wiw38Xq/KZB6Ht3QJkvxT4A5QJRiTje0Mtp1OvMY
O2cEbL0IkTYGr/rLbqz1sVFKDxfjvDb1/+K5FKOkjsJ3r9QyGVQps3RzzUiLoMlS
0wLF7NgDxIslumf/uQL5Q/b/9OMmSTzG88Gss7CH3GB/SQGolNkEZZCAmkDhw2x4
/+oD7DoTVA3FOruX8KOxDAZn4hY9X3/hywLdemMow1AfqPWTCElzge+iU7DHE9i0
fU6Tplg7ZuEvdXptNXRir0th4YwoYgjImlk9a6kj9NESmIwl7EF09iabhgCwjtzn
lvNXnoPANdn4C7v/JL9Sx7fOBFkDSGrEiet+bal5QO1qAcpTR0vUdP0xR7xqS3pm
dzCj/YKaVjrDVQqcTOwKlKyN2dZxriQZPeF+Iw+wXLvRy28vZY4YYVWgi6jiDLUF
bjwfftw4va6BTUAXMBTdFpJYuKqPpABh3gpi2kOb643DAc7UNiSSgfMAHPv1CbMR
MOSkdC2fm2pIuEsG8oLdQMvIz9uhVIwgPSP1XSfWbERb60mMow6MQH+f7peCwN+G
XbCWvJK+ckMH+1Yx9UMY0WXESptPNUA2B0d6/jBtSCasIFOubhUUjFF2RYZoPLR8
69Llo6NCT45dorirt/ZVJp+3vYM/dOyhvIDczG5Pi6qxWJEPJo6BC1nLJ8GYnFhu
Zi9n1lf/c9/SckwMtUjZn2LJbAY+TZa1Q6RQEaWXI3vri8PDFkMJ3p7Ff5b3wkaM
edVMfi3O+uWxPJ+/tDq4cKjRVL/iHopNq45ejFggKu3Civ8+AcOJgEp7hHn1a5re
kFz5Fhd9rzxelB9UjSnUqqhY9dtXGg2GcpDFG0e0ZvWGoYx/6uFmq6U2hmbQ5at0
sfLnkc81kcZ0u9NfnSxnj8v1Dmye8j9kn23lyrv6aA3R5UYjgf+HqywRwTcABdkF
LtNEYpKBIWo21kH47HzfLpXEQwDQDQ/jTsdF392tXWNhMUCUOV5pjIDusADz4B9n
6uC+Lf/q1P7kixOdIbK6/sQ7/Fo5Fk3ajzGFACgZNNRM3vFdwgyqacMD/WgXANfy
idwTjcBKK6MUtN+MLk5I87aonmHxEpCTH0ftpRKvvWXH4WIdF3R7en7wSkOMQVEX
rwRvcoKsvQXvsJOoxHERVnZU+nvHwiqtAM2zAwbTHn41ojAz6bq8FbN2MElXDd00
oAYfUqMgCXIKQeqhSit/oSwp2+25KoalDJFI5TnKY5rObaf4ExSSvLD6T61lyD2Y
bye3UZI6oecTtKb6FqJmfqoxTK9JzADILW9R3OAFG0dRDXEOKh4W/eht4VB2XDaJ
LHsmLLBacI4iRMg101R6aNqsXVcdIcZxxPRmVuFjTZyZewIpj/6k0vXgUaUb4h39
P30uR1HMsNAxFGj85CnMa4I0JzKXBh7jHLZ7dp/ciVkkY5w8zUHms7ppBuQKMPtE
RPl6+1/ILSqrXyPZeIPOfKccONqBh08IHmW+y3lSEFsRAAbOp8VaT+J/lIKI7CSZ
SvIElzWOfuiSpew+Knk8MfgnIUW3G/9QwDgPg4wXWzBiW8/3kNZubIag+2FEY6KC
65dcL3jbjxodEUYqEm0fdp6PDvKGMoRr0NC7ZXm0BRuOs4kuJcaW6BDbRjgmAaFo
Hjo2p5uZeaiOshWVThCQ1DlcWKx2PGLbvR4S/d4vfty0ZxP8F+4XEkht8uwc7GHo
GEIIajOWymU8FZmhQfbI2y77KAGkKSEDt1C4CRa4pwqXnY/SuKXv7LNWVouvNq7l
vL4ksODEe2XVf8W1+6CPbWAYtlrkDQn8UkeS/1xx65WnPc+4vMzQ0EpXoI/6+6Z3
QIMkyUW0Cg/i76Yw/lyORT5htAHcgt7ob56u3dzgNOfgBKeKUFNbur8Jg6oEdVNZ
mpY5uWrZMDqT0DwYdB1qJp+St9jiz7daHfhCbYdXDjJlTIcsqVmKTXLWCdg5cJY2
eExZm5IHMK2bPu5lQh91ySxYNWWHObgIgosOglPvYRtsAtrb9oMGiYFpv7tzat/5
G3tdcC/E8JkILbGY/6DDFtSMChVWSRO5Yb8qDbGbWucZdO0OA2BGFVsbqQND8jjO
/WPxedIzNSJVzs5+eucPlRq8TBMVXdkxeFJoqbCyDEhld/OckWvwG1KyLMX5QPnr
MTkQQupWWdS3Aed5CE4o014cRfS32Rt787cc6OAVLkkwj/uGf9OKRkm+daF8n1PO
mFneWoF4btPTPcXqEM8JQvOQ70O1ycXZ37B9sTc1QZvDUPx1uSMeQZG3j5ouf72C
R2v8w8WcGBfXKMaG0Fq3V9dcOmT0PwV0s5NArsk3qggWdo80G3uGRVhfRBaMrv7X
dfurFkMvbR6Y9Bsrqw7SNRfDq1U+a2Md4nkYoJOR0y2+1r75HQY7Bm1DJ3zYrSg7
fnGw3vlVrP1d9e2/yrieSKyT8QUKrfBuYREJD6yppNkikUOuM+U7m8SAqaoGBz7v
karLFw0gmRXzw1mYBc/agduHjzWd83OzdeKvEJAaddvEIb2GcxeAYM/Rcxm4jbXK
CJj8fs8zbwCh83rNQA4LTOA1F7w5R1hEgOri4ObjdRc5ZF7nfuJo737uWjlyF7eC
TOWYbZWt1zO/gJym5A0hM/vTre0KiKDm490eQWVVtssVJz00567waVG97A+DrgNu
Vv7jjBzGOxf7wOWaWhiGv7UlcYgIyeeP7nXvLDYxDXMTfZj6zHLiDWHdJrOTPqCD
RJcH4al5mz9DWzF1AKPP/jIiAYLK/Zl917MwNeM0cTJcjyqKNCqUColc13CkU2uQ
V8FBiAdsBxxqkcrbzbO566kqtlxw+t0xPtcBiyH/h5gaPu9NwT6ixDzrAVRjbFyN
rsP7S6NtcijWE/BIiL4LojtuzlWXsoSVvEri6zlscwrfALOZk9sA0Ur5s3QLWxTU
Q6fAuKoczsATKAaYZ62MxUXKSge3Qz6ART2fuQA2CozqfCypgvg902dZXK9jEjQl
F0z1Dcy7iizjgKs0D9RSXeo9dsYc+uHHt8GYKACsiJc+thpUJ/6WHlNHnFCRTju6
Pm/M4gIrgkbEMSUu50J1ArkSLk2xCYZJiglUlC2LK0X3EWHX9YFIL9XV3BkE2YJi
nIpg7cRsolTSiomOq3PK/2e+OV9mDl+e98DbDCglFfiUS2SWgcDgybR21cZrYO2C
kSX5hgsPvwwpW/CyawlYHMuLloYFDUsOgAtRl3a1jLhIq4Yeh7qw9fUnO+pjUpB/
SoBZ+2zFi/Lxxa9IzcipvCOWvGT540IU79uAlvcrDHejyusVERDzNiy8XY4HDlMi
eUpUZ9tfqInZKoFgB+MVS5C+siKR7h3wUimKihCm2fMswwu6CB+Z5S9T5GIYAaw4
yYjLaMtlP4DrmYnNCTySfRHePoniigho4mAC4etUnU7MmlU9K/8kIBx0Gb6TnqP9
O4hxcSUck9pzgQWQ/DaPthcRY5IxyBWwPy0KUE+HnHOA7V3FiRZKEnrNyXEgy05s
zro7IYFHZ2IRoCnuW10J23IYXtFbbip/ZrPzDTvyauj0N0t5dN1N6oOyD2h+cBaC
4RPTUnzyPa11iZnr+Eyc/8V3aZWgQ48zEQ0iw1oqYFg95d6PPcpNBz5+WtSXE2Ou
kNxA9VLYWR7uTYkiaDBL4QIx82L/cP5t++MdyyVEWrYKThnG0ddJjazLrFFJt3Mn
Lqz7HeXTwK7BcX6wqLXgX6xn4emjvkqAS+RdFSqNrMkx3zFGZQwkV4+dep+izJiF
5mCgSl/z8e/oflDPrUtP3nIuh8n4i7MM1qSl0FC8hH+41Sy0Npc6U8omg1WVAUEf
OfmL0xhh9mfrwsTzZWEJ5C+nd2PUvYT2qnnduhGugUxVc4rzTlz2lpaGW3lu2yOE
uoKc4G1CheQFszO4bf/IVEC258tw2X4BOJ15jwoBjnFdQm5nmXxksnOh+/ztTfqT
kpCdWAUcEH+PbIjj4ctK1zYdqPS5+MhVeHTXmjivUA6t1CyL3RcltxqoGIw2/gY7
hS+7gl1gq740WaTRSOGqRExrrUZy/7cuZSDVYjpOS1BNIUhTJAUtRLH8sGV/ZQxh
wxydJHsQWeF3ZQlq9/IPEZCpPDUbTFSHEw6o/vkVPuJPRzgsimrEvfElasvRBs8a
Vtm+wOoP8LIhbF2GX/C6hipgD1oIXUXmgl4keqStmmLohslUHn0VNDn9ov/p3DCN
TchiAHDkBTxUjZ1QRboEtHstY0uPOz/zov0D7VFYqRL18EXxpwk6gDO3IwL9dZgi
gI73X0kcZII8e8pQdHu+EvWW8yXoTtXdTaeNSwPk0aLLq19FQTArkwgt73jxZHiS
2DWVPkdnki7ugHkgS+JExdUo+ix4TSOgqVVX1Mymyp+Fesc/Bmjei2kGlgk/ioNB
KwikPB4MOXFwAreH2vFszizJf9TdlI74OUVisFCxqYP5hcEqLhReRWqNYzJb6NiG
x/vmk+FcVjdlBPV16aj+uiDrHrwzU9adjzr7NBlKb2qrMRPaaFtw/K+1smU+ax2q
TdzAU2hCAARckqlbfEpgEOOi1FDMm5OYWBUFRRa9LV/LjPoib/B2rQMmuG2cmgw5
RPNbplaGym8/LU+W4AZixr7kZulIn9Wt3+yB/U+cpVhRp0YMdY7TqAqJj+aHPg6M
3A5FW2kMyEnV7iERTubLd73C4nCSnpjlD5Sq6Z6/MFbH+vShegR7tV3cGCD+ddS9
GKP7jpBAAhAoaknyuai8hTpB2ImTT9jR/i3GVRF6bv0sSn3PntMugITWAyYb3kFa
OKLtkf2P1c7EuRSpnJ+kf4YS+C8sGRrl9WrUYo9jhjICOiDAyBl0lUm0A1eVurKs
OkeY3Th1ml0rdVa8Fnqnn7yUeCRGsed2W3MAFre6NpoeSsOLK4NUPc+3pKiScnGQ
iP/gHbrOaJuTsyMO11DcwurFXTspi6LJHIFPDnip/2RLQroWRisJ+8EoZTDXjajn
4cTXcYRsR5U9KgD+vlxaz0ziUhf0rSnX02M2pnhbw0WyF4iJDRk+ggRkGiX8VFOK
M5tNw4rLdfvaRyeajureH00dgpVhzwHGZkkj5Bzs9m7zDrDWWtKLMhA2MfoKMSZN
9W7ebsPCTPgg1VeFWnc3NCVe+6sSixQd7Zm9yNPFt5fMUQ7rgN0lJhw3alIGr66i
ZEkCy3PV79JU0jAcDl1ucttzWV1pMb2N4K7JdLHptKd4sl8QeJBhqi18HB6Pj1Cs
6mY1EuZJbY2xsPHzgN1Atfocn5mh5YpuzFmoVt7RpexI8UjzKDpWaCZiJ0yV9+nZ
yY28DegfhKtkMCxkTiuV1MPHWqKSmtmKmCUvRqBgV+qBOsy+2jKC8EQvUE+LbHCe
asQIN5Lui4pXFSumwT4aElFsAM0I1WpQkTWkIHU5wZDzr0b1qpHOt/MD2aUOQ1m0
EzI8i7MxUPEd1IwUn/OG1U03q3DU1hNpw64FYiH+JA9hMb0rnToFxa8zF/LxIhir
dqiVvgufEhQW2ilDyfDxwJRfAYGGgq0m7KFBN3OLoo1IFttq/tGt63TazagtA7Sy
IjCiKfzw3OPY8Wyq+yj22z1voZqmZFEK0tgLrVXtgz9iI9D7+0fc3v6GC3+lsUiL
Ofe3jUawZ6yQGnaat3nhia6PKM60yFk36tWaYOej3fidBAmxpkeer1fjQWOVjieg
lhfR7e3ufO0JWq/YSRHiLpiUOafhmix91Jqz3QrBuXT7orU3S4BEMGRPtDqkyGEM
PW+sLrJwlChs9r/+JCWOejczr+aY5nxI9hwfY/jSgSVhtqFkLoYze4T1EbPyhlh4
2NfnPa4Rl1DDfzWA97fXGqPaP8kik78YOA5desP3qxIZHUmVC8XLpjNZ6px3Pqm1
kbSP5mUD0MSorvQ2vbWSxsjGq9M+ADgsWFmKGehhw+0904IkHo8sXE9ePOW7WDyr
7mckniDN0qraCyAyAV/vmHnqHoZU4a2qm3DTCQz3VZNBiPB8gwebEx4H5myjTB4K
ObO28CKywiulnUCH8RPHTZVSY/HDk3v8/YljTAwUN3nvNJdKhq9yZRqHYMMp24+A
WxYJ99c43j9yCW4pw97Fqek+GbGIkYuESnrw5l5n06C1PZ9QnaU+wU9HsyMg5pSG
DZ9Q04WvkJki1bglIC2QbUCcZcUzAx1hN2OfK0SpOzBkk7P7nKHXv1/F5Jbg0jaJ
XDI4oilQN4M4vgFgw7u1LGARJeZOK7qus52yN2+TcCxEKL3L/PPI2otPY5pSDg8r
b+iiY7Gg+fWbeNR8deN2jFzQqkDjBMFw9WCiCvgvXjDEIQ/qLMihz5PLrYb+BbA0
6j9P0GHL3+j95f/ENNeC4uca81cAzaX7BS+1r1wWltWd1YZ4rOGTyPIkCINOB8gS
nmPd2dWlLcEuFvFILWYH2sqg4EFkbU/oqo06U4Bf+cY+FQLZ7GkWkW5Roo6Lfe5d
Pt6NlQbEM3N6NxwsbDzgHjQ2taq1MpS91B3HEkLVLtdQhuMvvFf9emonMzPD12tz
3XPuJ8PqAYOUzi5bMXBqobKIhvjmCdJ6riXSKo/PVvOTvy2FYr6l5ndPMubU5n0k
NaXVXxtLunyxMscdNw7v6m1Hig+nJMxrCdmkeyTd93B1KjWTH3KHLsGIBpO7cnLH
0axXMqzNCbqIjfxcVRtbFFKarGvvhoBx5X9fY/ZjBwpPLkuGNEYaTxXruqKi+fkF
62JaBAQvtsm9wPaM2+lx1NmXMIeN1JsIsldm4R5wSgwG94FdLEDJIWnBCtIv/3sV
0sPKAzdSKICI7CuJwxhf0DhYmf+mZvna2+wZ32bnGqaHpljInhnGvt0Fgs4Hj0JJ
ht/V/QAYvsvdA1I3aIIRUCULoa/3cTpSDkdus0scErEJsJt8PXai2gNS9QDFoM0K
E8YDNKd9guEFhifDpGS87B5xvI80ULcc0DOzXSGuicjnFt/jV1WxUDy0Uhcew/sQ
+2Yv2EglN22ikC6x9hmJ9kEEqUO1o7ejZ+QJ1vnIgEFz7O6OJf9vi35mstIw9Cs8
+jZOqboRtFPCg99ZZoYX3cNygWXi3NU8HuUs9L5knYwm9tWrbIcN1p0zZp1dvZ+d
w3bxeE2k2GmXNu4ZhhOT4rSC0NFsk+Pi4Om71TFJ6R7knlnlZxt5vA+VRmpGfVyc
V3rMW376bP/v6kuOC77Fl4ty1GVHjcPZDPXLGlep+d3EGf+lT6LiKEnI6RZx2cQQ
gDm7iEVZXdHiRQEnsfsw8CkkhNd4VE9d61Cbeq5/xMpLmYGZ0LD6Zqsw2V2santj
2+brvxjqd65miPL8PbCUI9PvMeLkRqu5vrMGnR6LAUiQSNdEltsllcgyMtqcuTmx
bG1x60faOQDJnLVBRpreD2HAvnnY+97vGTTjd6srNf03XFEo+1bY5V4HD7WUtPyO
uvcvTMIng0yhA0D8FAbnhCF0ed+tPsyAKH0H8ou8dyUds7GfuyiiKReb35ESxPTh
+yqsVATxnYDKMdJOA6KxdA91L1qWf2mhhlgi3VM4yvNxsgFQmjQ0UG0GIQkkhyHZ
UZFBiIDT4cxa1EWaOukdl/1Gro5nDNfkH7iwKxveDVfUV27fr4Z/SbcdCXdWlzbf
h4hyJzqKBu13TOGsfjQhybmXq+dmVmJvNP8zafyHNh++2ETUO6xJr3YCQJ7yLP1G
tj8AJJSRgHq8EeFhGq9dlEO4vLGtnmHjlWlTgZe/rJnlflx0ADJ5z3y+g5hofbxZ
Yeu7/nJ1qqSl47HPRF5tjRuIBN1DDbbgGjW8CJvfswwHaRU0pLsnShIlT/x0koyI
uQuWRU87xbAo1/8L2xN6GmnRCz2FJ10YJiGyQMJSxaxZ5Fu7IiOOKLKdcO3ureBB
8nU9Nu7dZXwe0V+5tIwApKcgESBPV4BL3edYIslpTqJc3YQtPeBAKlC6p8DL7dUB
AFcKVkaPs/dSKwGzizHf3E48PKKVQqc6gUWj8RB/FZ7/+ngibBmNsIVCoiDk11hs
rorR1/ZVIWl6Wv3PqATlPDwGaIHPxYXuQRD0+z3fMrqGXVQzYlaoPR7r5iObnsBT
1NMa3WNbOXiGPFnURfvvwW1F+Lz6C7mh0JKdD8XHRoMF6MEtEVtGlxvDGl/QJvM2
i2d5dZg/O5HQyGAeOKDIfy38gbKEq6+ERAXM7W0iQqqjiRdgrfFk58ICYMjgvNxZ
cLdgPwofXJl/NBg3FVVprraETk+r6PeBp8d+oBIAIhHW3F9UATSwwUbAr4X/PVSn
X6zRTM7x+aqVN7FYj9CB4sqNiuwH1/qvKeehJ7gCbMSrUcrRVMT80YlxPOtRSFY8
hG16gctiCK9TvedFjVCP+NVRdRYqXymX2IWZkCvztgQylFP/ltX6+AbzPIHLPBh7
xPjFB94NXFFJuz1oUVgTRYgrzPea6940XOIqnouaL0hL/a+Dfd65MuD5diufpgOC
PFb78M/+RqiT7P7oSpG1Z1SKQkRj9FTAx7y1x8SVEYsdYXbpiic0qyUUJ7K3wMT1
A926oLW+r4/wRROv6QHfpOnDO49RalbX9yulVeRrGNq7DChrdZ2inaVYJeUr8vY3
bkXPIMpFQ9vmGWK3EElnkN+hDReUEJ89tdExulxL1DRPov3WnWBPK4gVXqi2SmgS
QdakHZWudxCECCSfQbGfvN58is4JALGauTxoJZRpbUFD19B7WQ5uvqAqqozMHk9W
TLownNsYdAYO8f08lObE/tKEGC2oPb7dprkx1/fYpP8Ts3QfODQJiBvFp/YV+EzL
MQln+31lchkOxm7oUKO2d64xQvqKi1gIunvTKOluIUk3xLRjjm7qi7h616lr4fc3
U2HFin5P6ubzKXRdHaT5dNw3Bwzs2nyLqvhpLC2fb4RVSFKCLyG4Lp8Cyd74yNpN
UDZfFcExrCJ21pkWGYcYZVGFayU7VcyEa0WD5unonyHmRmCnf70pm6l0DlloUuHM
Wgh77G+0tPMTDAnBdZrMnoHxghbihd+yosNTXZpvW6SEzy4lUCJaDZFhNgxrEOox
8KroA/aB8+LZ7U07cmvXfRmdX59NEg1Wq0I5LFdomqfdOnRpxlvTUOoUs3q2uLUp
Df/4B5Ejk9EdmSdjg9y72V0vaDADw/fn1tAvT+PITnymWvfQcxv4h8wFwsYLZ0Yp
Tga+wqj+wbSNfs2PtQelNFRpoY29beSqWyV7n+40xgJspml9xzJ5RpbdQjZIaCkK
XLY54d4tbvUOf4OaYUQKgdQnftPntp7sm11T7CWQH0ZjdKbv9fLdhrhojKY80poT
TvBAhy7PegwLohiMdZRptPcM9JCkfFtN1bCfbdfLPwyps03SblBNRrnMl+VPJQyQ
nTnQaiIlkSlr36yjxUtfuIuCOQUm++0mFfoKhTAzmI457nWgDK1jSAmeI7fkO8nY
xRJd+ixcqYZKbF6u0qS5QpnWUQminvVurGj4yE6ECppFsw2jckrEapLJpFlUXjIx
Uw5WNFHiQHoOXFIJeHPLB/xhQ+9I/5eX0et5ykPI8tPFGunGrx7721INVG3kPnHV
YITPTKC9/XmInBrlAQXmRet+ryiaTE1K+RkaRJrF1/rwoChhOncaKcjHXAtE42rM
FxQdb0Wb/Mo787OvRAwHBn9zYc5xE3ZxX5sFAiISw0RecrKFuMz+RA8Z+k9KY1Ph
0hFI5TACWNKlDGCzrL31H6aiMAII6MZV6jvKlrmSNjbzJhxwVj7VZY7breCtTNt2
8WxbAnlFsXaC484ZHXi+ssVPd4RFA4Wvucfmva8QkJWkQQ2oISBhBMezcB8JadyL
iLzNmc3j5bikVSejJvpmtNmQXRls5rWLqUxPMATuRYozPL/cbVoA0TlhdhZsoYDy
mBFDoy/jzIDkjc+2ez2pINMTn4VMFSSYrAfIxsggUQVDMYIIyUTorjeVeCAXchuD
8VSA17l3VJszENUIJgemakelRe+QcYi9+MkXKcqyIqgx9nKP0H2w5fieQsGDI+yK
aonbVd9dmtg7ovlnQvsiDVj74q+vCDCTsZQo8x1UokvoimOJZGZq+/M0UY0DBlXB
WJzOTpnpo8ATpZ/8TpyItJC2LJtcGww7k95RUOC3W5dbRY7yHmXJb9w7eQtRw7GF
M+/iXKiGeyod4MLvZfe2/HHdOoN0i8EEhsN1r1HPdcMlF+xi9Cb1B5shZ5ORbYxo
TS48LIiU1XVeE2XVLC9Q9M6fsYbzR7w4+W+2pUqgicx7JP4ngfPfO9Ej9kHNGRx2
muCutIRVUmp+301OUB1ImuWe2xsOMW+HfsmfucwEelwFW670mAJURap7Lsm69vOu
VG5PXTOOt2lHAAq+S0z81+CoHMGdfJXIq4Lw+Zv6HgtNRSi1lqIa85/YOkIfBoVu
5QBd7DmWbjRsjfhfvZXkmqXjrkIb+6rFMI+kuV2luAtZfmd0eP2WNqZ5Kehm4Cfv
ftjQAiaxpHA/4pcEPHCo39KhAvyCoZaXD2U3wPGudFrwPJxLlRXHZx5+o535PRS3
n4TVDcXSSZpgEne0qmUkGktcy6Z7nJGXbha0n1+Cq6A2h0MjRUmOlPxgBspAkwuo
FmTl/RcmF0DFBoZCZKyb4sTF2WX9yF0eDaMkezQp6zx3gc1y30C41yu8itytlA+h
0KzQgwR2ndL/m/LmOj1TpPzpAGxP7xAJV9S3iAp68zJbcSF+lX90skD/T7FjPNwC
GRZh3Ne9QW3nulLO6shpMo2fHUpllXng/oyMYeRVmRgaG62vi0Hr8HyowYC2eq6p
t8U0r5FXH8Xv/GYmUBqZzy7yC11go4u06TeQu7eXDU9LfugE8iI84w/djm4Rpxjx
gJnQpfwYLG7OlWWElMNT7hehMxx2q/HaLU4F+npNlGZDLgvNwkAsPrnFaWGZ8+cx
C1nva/I3P3Cc8moWGfpjOlzy6SYCANNbunq9HYXGYjxqMcgQFSgCJSLEPbRc69DL
Lv57ejHEMGCcu7vtqCQHp8Cq1FwICow+DNsPINUJVBrlHIA6B0RDmRkufuMmzjI3
dmXIyFkiqaDmfgqJFCLb1p+3xavqZ1uDZeVUgnqRcYebU1t1YOEDu7XYAkvoDLZ2
xa9AbJbTnLDty/oU7Y3AoT+VWxrc92VrT5UEWBcqSH0j7TAwkCySg74Ncn1TP1lz
32LFyORnXz2q03I1NvP6XSCRT8z+f2Lqt7R1zXxqij7ZByaN9XH0IwIExc6woEC/
AtFU/GbTAy9+uR9MY2w8iCnJuD9x92UXQcKCJr3Xj0d5uSxEjzuoNDc8nT+ZpY9n
RjQ94K+b3KsdS8HdsNSacgDU9Mp6FEspTfcxdfG9k/aetCPpJjiVxOyyvqEUZ2/q
XdjMfT3bvXxBkZ5vmJcou55tFP1ZMuWnqut3en3xs0SVpsrZXijJqemlqwT6ivuH
fn/N6gQbnkwnLAbm1lS0XQEayinv4Ethk9HQb9I4u/X9k+C2HuTi4xZ3qj1BhJG8
5pV1XFHIZZYC9vqwSaCWlKq2PQlWFRZhZx5xkQWjD2VnWbioeDRR1VOBo9iTwYEU
bOKBaUKRAY8u0QGyctVGYHjweaBYj4dM1a39mlvfjSQonblQH065A6xNGgPpx8hQ
VbSxp3TH2u0RPf9gcd1QM2uDZpUIULtkzaXDWjxBoUAmOEXp1cdfa3JlFJZQdfDw
Y9i7xygfbM71KQhMRqJifIIm4O2SxO1yGdpGNwpTDtPWxWLBiyP0jtYAdZC77a3l
wbmaEmWMGOoQh/W6NOpXdkUZJ73JFxeFzj+Etc5Es2IhuLX2KYhV+MtIb/e0aGtI
iMR1DNsXj2MN20apkYwWLFGqwSdS8dmQMKIEN7GEQRjgIFoTIziegXc6S4HBUmyQ
6QS/UVdxcHDE+l+FQsKwBXxvpD3dKBChJOcFxEeCxIz8bT/XZdQ1jPnpnCaQrHOX
ubyLUQYyWrKQlHu5phsZ3F/msEkjqoIpLYgGObYgc7vBM1j2h7ocvuoTo1+KPWQd
FG9Esdz6ppGjphxF0esUUlt0ZSEIa3yo/96dORx5w063rXorQARBUyVrclHQaeD1
oknzfAInrolxfuQmKu7LVdFGjflpz2O0m1oEcKjUda1ArEhkxixACS3kpYphl+Ow
Q+ch1n0zNky2S5D30yexjnL6gGHX4xM9HRi6t0lfWrM4Z07ot+vbMVoNWgsWGTTz
6GfSMRhS1xJnph+c4qDCAQwMkAbpWuDExBlS7G0Q7rzfjWM5oSR4mnxrPk5qE/kj
0qONOo40DDIUP3tLXGUywkem0S3ZQ1J5z1vOi4p0YmGCs++x7TfwtI07352xDl8k
fw0647j9FS1kkvVwLq2qMG5F4HK2lT9cEiFXnztTlVitrNuI/btOLVzPVEl1qPu3
Kl/0J/S7f13bCXb+UcJhWonpsbMmk0wuBTLdULOslDwpPfcvKf5kJ7XThILkyYKY
3QxkjKc9E79tKf4AFKdLXtEoyfvrbmr5t01T0JM43SZ2IM7upf//Sq8xC+bNmOK3
s0aVB4HYKkImdtaNyPuKemXOnHb0QZJbhw931WHX+qaRjImzHyOxz0QrLs9Fikcu
1VdOyFJj9PDNRRQvDL1tI4OovHetuh7ytiodnpj4tU0el4LzRwDlrcbomjmUVuE5
bilpVPJ96v0Cs2Dsbkj78fNxNWtfOx7T3I3aUF2VFMOZt2K60+snk2z20BnRUegQ
/drpJlIdKm2A3jy51bAy6KdJf4hl8SM3qQDkNG+qHPzoLX2IFFYMYTXNC9Ps58LF
ug0OUfsDbc/oVmm25lCr7hZGP0Mrz7WEsjoEBAO+Wum/hV8M6WR0Nc3u6pM038AV
kPPJs9bh3PXW6J7GXPkBIQu0O4oJllpPR5iD0jML3HEy8dbC6zpX2X4GLgVxb4ws
GcCVFY3zQgoPxfOcukeLchEJjCxAgdb3o6Lfaq9LX9vJCfl1sS42ojtZQcp6KgHh
oT3RcE6UM800FdjDdjDSe5MdwHf0K1/ah2IrZZtFc6ifTTWvcf99bLT168PKaSit
9R1+Z4DKSwbV1r8KhQzmoAKOM9uC2tww48cl2ilE41Dmw7lm7QKPTA/JdcX1XohZ
+iacz1Qj7YbUzphN4ueOzA1CF6A4gUDfaO0dcnmjwoTi3YAcmn/tTtHuQe1XSsMj
3OHxtOHmXHrb2ewW/JsOYZsQANmZQbrJC6ZZJ8dkRZ+4ttI7nwM9b7CawMCGnjgu
+2liKzOsWWHDi9M+j1NPIMpRHLUuGjcBSnZv3YIwGmXcGZoOOdzlZKorExjWJUU5
8e33wDpG9RufRRHSfGZDnwetH83emncU9SGixKkGjvru16URu2vdz9k/HjqZ3EO9
m290q0mzgJFHSRm7b5HJWL8d6C98l4JgbpJ8n5JcGl0bB0hs7S1JT2BAiKhJIJhX
Np0IX/l7lDC5vf8zhOdqzZm9lnr08UAHTwcqsPsXuAmxNcbx421Rg6dhTQ23NZAz
gzjqCvCfJpr+DGqhD5xsjghN/SxRnREAK2+jYfYmG4domHIBY6u8TMQvu6jkHGQ9
oLlFG9cDudvimzGg0IwXMQf8IpVbAg9iAQq+uwEzIbodV4AXUC8dK3CLQvbj7q8I
XcQ/pGTfIIsEPtFQUyzOnoXjklxWe4wIc6u3yiSplXwTFaJZjtV1bitXyezBsJwA
9g2CvUXVx/FDJ2p9sRiRxfbaJYgpVj7POlu2xWXYJvBGmp+jvtBxer9gY/ZOd8gR
LaBAQdKFlOmQ9uYMc4T+wU3BPQv/CU9T14ZzRqrMeeVjrty5i2Osb338FiG4gnQ+
K4eUEKyWqX5FnOcG7xNtwK4+nC5xvyHdNx9ZlTy8r65Ise16E6lufYSl8EEUdJ68
Z0pRqFDpZVVQnTkjy8uDQGqSG/CpzQV8pyp1aN5zu6vaPywioqD35MFW9RBCPQ5X
7Qo2urGWMU3IUwfkh96ItNiz4jsvFGjasqBqz6EeODH7YWftcM6dJOJWDTsVDiwK
+MMXYOM6qYnvDBIZc24O7etFR9y+pFo5eA3NCrNQnG4B017VyzjySgdEHq7Vyyk2
vjNPe0oXfAg9TXjH824CTxC2eZbONsBsc9WCPSGbXB03j6a1AZSrTABL10fUF4ah
eAYp1LMwfiKm8KC+bxAd/R/QxprzAE9YwesATFNZr5IlGDbEDXusVtZWqtOJ9uvH
DnihT10uATlbIGm7P13hzTnUEu3JUOcP9ex48BlZJWFB7Y7+0HfiVJ+CwACQhopk
A3g9KnaeMyA7uyPSDpWNoFDaO6tbDduVSs2vitd59fi9U3f2EYQC8VKJO+QTOkhp
vN7vN4N4ZqyTgu9brKML6jGfh4q8VkG1EtOGasqnsQfRgAi1TzZgMJwkuzqSP3H5
FTdzdw7yCqrrDMJHVMBdXp6QPIxpS+04d8baeApwSEvKXfIMDabsEOgcin6tp54W
o2tnwZE4k0N9HiSLCy8GD7Pd/n5QfylXjpUzn0suzNCmUm7kLaSPq8WpdXGZgaN/
NC/MpOKD4q46pM5GhU+CIl5pppZAwNR0dlwgFjrqGw1TkxC7l6t4XYwCfMq8TIeW
Yq6wEenACR+rp9E/2zE9F7DCbJY7sZcDfjy8fytgXm7V5lM8mm9d0KMyFuLyukqB
063TkFLkNaoGdoo32bwmcOUH4a5HdSek/dwE4gRj888SILVvmwMrUeoie7DmGWGz
tseXcW4Br9smFibmYBbhdflXGEcGEWXqBY1Tdfca2T16gMDtBmXiTocNfievRLxs
syvgwTqlWTWeWl2t1jXP9jvZEmFa7iZdD7SDsZswatN1PCiMdSz8wklcUrukPybD
2wjq+9BCLdmDqLL3IpZUfj3e82MT/VzG3RqKyrij5DCgfeWje9fSFdIB/JMst3GX
tHgl80azJ+gyifYMPytSGSpB1tzTLYy+kVWL8wzmXP13eQsoIu3HNSmjf6HazQ3d
YeXvUkwqbUSKDihkewv/N5gxnRMk4vUU7Q55cOJ3m0JM7v9L2qnpdYtyRMS30Hlf
kY0ZQJ8tRCBbppXIrx2oi29lv+yZki3y1v6wTXzY1cN/fCgQeSy4Afw7TzphO9nC
tFiBQ4DUGFcWBwvPUlK2TArxvMODuPcy5HTPQi8AMLWDexDLu38rP7oY5+b6iVGc
e2+icqZFjIQnAy7IXmA33ON47wh8KNRDd6fQ87FBPaQvAQNHCYqtkTGKROeZwkFK
gBWOJwg15IEX4vSj7657GuV+wQk2n8gDBd6a1rFGDzwEP1SJi/ineXN5aX3sMwhn
yccoQdkTjbAIHmFLaYzogMizWz7XHLCRt9zegiTiiMl4lSUBS1YaezBVZWscqInV
UJAmxA4QkvxP6B0uAHCMrxuVvAZCwzJtgokm7cpZYxb6tqEb00SjPQusSWcdHT8Q
nAixsaOf4R+uajV9sk/2hSN+idjitDH89+Saxl9j1ZqGB4tsF2u4qGjFoPnEiUjC
vJrqsP7IuvBsKudfjYODSJq8mbvrgRGq6jkgmsXQkOD8wIT5/cadLFuKb8jexx/O
WLgOhNgrtCYB3Nd7dq727uJLivzSMHBfqha2c+MF2NTcwBLUEWJ3xUiEtx5QwysS
E6PZs87zhMKZ7k1TfdF2PC/fXRdCUl7BhGr8GC3ON7j1QLqDj0I8hnMcNHjEnOai
6oZY6zdYk6m1z4jHIWAgHmiDAWRpJdiPGYzgqp/LeYg9veidCp6RxyY5MI6yBaWe
lj+TFjef+xAPtNAQsKc/YQYd8Nn5RE9tSwyr10QculEpP/csFBOP3sE1mUWyzh9f
0QaWlT61RR8V+vY1s8N/50/Dt+e/IFS5tXARG03qi6bKxq9YFP6uSnGC2ETqcTUz
pHpOe+CYoFgPFm2r7jp0GpmbwQtSi1VuwcF1t5oZQpH9ZdFdW11FF7HAMIPyB0y2
pDcrQHp7cqIyOjJ4rcs1Si7iUedBVYUs9/mIBoBu4gW7UFCLU8l3nqaGl/tJXk7p
grIk2dDLWRSXVykycu1RRQLEvaHlI5KXjqtdT2b0V+kz0TJq0ivhgp9d00zfJnx2
EGSl7xB9F10ySyQfIspnsnGSn7ZC+WA44httdUsdRZAyIDUT/PrUBH8KNM729iu5
F6HVI8Fh0GVaGqU7WIb7jr08ugSdtvjVoiL/qc34qrWiceQM5G+25bKRpdwcQwgz
htsff+AJ6/gQ08RjWQQZEScSXVlY/RS3v/i6Rd3ffTzeoFiQLIOcnQwWwPMdh+fY
Pqzxs6c3lx9T4xkaeIw7r7/H62DqfD3sSOXmQinfGOEFcYpYC/l1pNFYRRWeZoTy
H/S4JYkU/we3TYEcCd3IkISQmjY+CUSPTHbZZnHpa7xKEZnDvdXokYw8PBNe9Oa2
h/ll3Gq/b+vpGUqc5FAnASYv1TnDLhv0gBEyC0Q0hJ9PHjYmSezU8pGOvcM4PB6W
izdObckeX0epyMjSpzPVGIUk1Fx5qgQdl7rjcE9vs/lv5nXfTytQEsD80CkcXp+9
48FZ1aqdQsE8UFfHhAUf7d7FIpG1eYQbeH+qdBZoBJPLO38nsVO4/P+uS5lCsBOY
qhl4gT/fE48cTM1CHbUESJ7CxmmSgeB4AwuNNptJdbUKjUt7kvW/p5kr3fjhbyP4
HIWLaJHnQLixvHHhxuzC00FNtX3WqeFJXkz3xMawyGrM2miGHExDJ20uBrOQ7Bev
Zy2R291rO2PSoRHcFG48bVSEdYi8Cqaq+SxhGwDw1DfLlk9oJzPwJQvHW8mYtT+g
8bXNTEA9JD4/tNQa+tDpDzbXWeMBaO0EoCwEkhCiYPSsucR+3QpIYkoY5nVjkGYT
VGGA+VerkmnNpjCVZl3DlAZi+pbiCDZYmlTsm9PWxFJOBUplSywXs7uyeidGa1GH
sfYAGsnfOF1bZ7BfPgg/xkTUaU5eSJMlVMD2fchzxydMFHHXi1Brj9/TX20daxI8
nBmLy737aBg+n5CHWxfVsZLQtX3A4t9UGaNfz6Kuhbqia87dc6+opGw/6AgAXiK4
i2L1UwyHMSdhOtOK3mLuoQJzXLnKLBskgCX+7VKpYgzKyGHtROnOOym+zK7oyfMH
3ZsiKWGIUzpY/s6H114Y99HDhKLbIhpMLe4Y7mfm7W/VwdrgQU5UU/QcReOv5ogL
3RW2JKU95+EyGGz+HWpHTd3hvSFd0xNUTm9byL+wVuffGNbx94Uhw+EDZnqeK0fj
zAbtfVZvygWEGhqNjVd0wmqVwdt20jDN4R+K5b7ku/kowJoRW0d2KH0ou3HqbokV
o9semCLP5+2AFHLDO4ZRPMR8X9eI/NoM62zGoXhQjNUmAszUpdY3DodmmF/xCpYc
f/4uS0pWQy4P2A+klapuQa4mTgDOYo0gDBeRKA7UxhLCU4EE01Wth48jUaI/PR3R
i26IPlSgptVzhhThSX9ZEk8u/B72T7jU9JDh4JRipT/gD2ot+Kunl83Xp5iioLzO
6h4A4QfaP2N9E7rLYGeSNQOq5VV1YXX46+w/VdnqBZDrExS/HqQXBgUwJpzIpwAE
Ooq77Ll0AbkVNLwO45J/yGV+XHoJ3cG7vi8twe35TBYrrHs3I98aIMaNPZc2eBNc
CYu4npeUO2wVrWW0NY8Zqgy5H8huvxy4OUptq/uuMl6uKhvMiPhhlxloIx44tkn3
L4IWBxGIkSMDxGS1uxFR6yyyv5XM+qeGmoL3WXtrWz7nK70VtLBtH2rt08bVaCRd
RGuekZR2K67u+NFne+ctx44w/9i+B6woAi4tGrnL8jA5GJNCmCzaQrTIqvsCbNJw
LX2wN0I/a6V5Jk7q8RKv0f0H8cVX0pz2JYDasLunrdnzOPdSqD6Br67+pMfvhi07
wZZ6klFl2TL4UKP3UHR4cUuzfhsTta+AqTxHQf14ZQ8aQl1PD0ZPfHVG3P6QzN2f
xG/5imoWjcUI4badFiUMqivxyLm0vdSLAid4C5qWcwRJuOx8Y8+90UAoJud0bvbG
G3+nzUd7Ami8WzTC0BNRz9Gkmssxe6KgpSg0tuwIXG3UPQYQSyTgJISccLzBJFp1
6MyBrXnkSyy3ZgAXKFg0DXlvB4lKjvdDE22/L6LtjOJ557w/W4IL1CBkaFq/eh0P
/n/fpOmAx3mJRARurfQkzjqOZTnpgap8dGTlA2NXiVOkRK2WCvt40lZ65QG/wE7E
3d+OaWQ4Rqb5oA1zZgGxNPDEx4NS+pFrPXWOevhW3l+hp/rKyxoP5/gEKipctleP
EP5umXtK+Sq/RG918u0fq8kopzAhUyRFtsxh1LBERhNSRHHnnUZ4a8giz6hPIHwF
57th6sBcBUd9UHZ9JEtwmuCo64HFxje3Fq4PFZFpAnVZU+DAMlY+1XLSEcUURQl7
KXT9gH5SD50qHPDfSRUIaBU76LxgNmIFc3k11uzQ1DB5VY+3U3lojM1mnGhCkbJ+
u+1nI8aGXcfLwiktZHFA1TCRc2xbX8KLit6HBZYc6O//XFe0gh17ySyLMRIa1bQR
tZik3fj7spwEEPeyLzC8N8AzkEh4hwWVqbM1hE7O7dfL4m4CciKqvWgBv245tPS0
vkp2I4zVLAjne9pMd0mPUBejD/z+EqOL6/BT85UfcDNWGCtM85Rcdv31ABC/C3Zu
2DlJ5JDx6cCjLDg61CtFKo+fIk9JoRIIgPebi1AV3DSjRUoAnISefL/e+GpC2GUF
RrIU0pg1Wb2PHs9f0zT/ej44zAruIfALGcs9tdFZex4S2ntyE3/PHd8fUQIXlQzN
8o560qHolJkNfAkQn2+oBD0x17dCxwT5xGjq7WqBj57BtqFBA1fAzfH10wJKw+kX
Iz8OKV7YfwLMkTsTa2fF1adPH2cRUqyucjgpF9eYD2NngUWGB4eArz7gglabc12X
1KxlGvi47h7rZF8Ju2pVez68j/MAdlQG5lHYZEu8Qr4rr63rXczCuApfs4ZiLPXc
sFYIOrAp8ZLTdz+B5nwlQKGKxLhZQbTPVDYaDvm0Qm6dD77cDeV8rgVW1wd1JU4g
OcfadRnmPGUGoQ+xc0R069bj89O7rjftlx1WSuZPxccrQSTt9MlNCjNzxjtvSmAQ
CN/GM8O5nv41Y9+K/qEKua3Qb55IqRbzQjWPsZBXvEs3/IwGU+D8ShYrxTthvvK7
bsRLkoymt4hz40TEU29E3rHoSMQNoAVbndtJIhb2hZEFBmAuOHh/xrJhWbwhcfLT
4v3jGakgnBjlHEU9nu5HrB+2WwCBYoDXFRBeEmi8iBZDRlz9Z7GDj0+0DOXwDqYy
Frv0ehltsWjbRDwWeJI911YRw34wZuipCOMtZ+z5kKojbcqnc+CaJNlTmnV2cXgx
xH9RE/l9C7qDzj4bqX8P1r+RTlBXoHhKOB8Rw07M+/3wS1jk9ASpaGFSnjlHm47M
g8xvuKyzMnBUy5roK3Q68+riBoQRnR1MFDLeqBG6fq3Iq/u8irYEHVb+B9AsXjn0
1jhKnHSDtlbEJm555+nKF9Fros7me/SkVImsyim1XWDrFfiwvk7LvA0Q4q+2hl06
GhE8XTiwbmsmRT4xFone01v3W/sPX4DAKsoWYVNV4ZBBpwAm1l2KnMdWVqdJ6STM
MXZ4K2UOXSqo/49OOfpb1OVrn7yThgJLwh8qlT+3TKbd+YkTOrQPEjCclZMQZCGc
booUIOLy2BpAKIJONhDYJ6V6V7A2gFP87e9RFSzvYROfov9Mx+DnIx74sgHEy+JS
YtCYydLJiB16/bi4FCRQNcOUHOXO3osPstRoSaAmmfVafjaN++wiLt5FSMrJgPFf
5qIjkJmMNvtRVSOXdaIpXnemr2QrvDrYOWzsudDYSSjXccUV6ur7gtn8W+a1Iz/z
0FkolwCieETL/WHzQmdQMbVnkRyY2rlkszTfjRUAqQFLLaM647S0za3VgnFv+Q00
RZlU5U6H5wagyKGfS3FZupLcOY+4t58Sq+mVzuCvdSW7g1nD8NXJH1a9quWO2HRZ
G+kyxe1R5IkOhOXkf4YdyoEGCzqX6jmk3AaU/7o8x1uz498CCFhg4fLMmjsyJoJo
ZdaRHfgFbiuRNHtU3LR4HNAggSBHE4LSCqoF4UZ1i7ENR82Z3utSTmUkdTiSdUw5
9tePI7Q1A/tPG6qlugXk6OaevEObS4S5qJHHLnLYO8jA51DjGc3IIGqsOXe25Z9e
Hnlmmsr4Pmb6SbXJyCiplVLZiKjgfS6F59Kfq3RmXW6qqYjtngeYn01d8kv+Jti5
+zgZHNSXKccaWIBYkeEJcEe5mH7HALwpNrIn7sl/KxZg7sP6vSwl5wuTF8NQ915g
9jp4th3sigHvRRJddYnc/HD1+ptolZPI9JDrGYUawr86SMlREcyWXJJV2/d4rFUs
H8LhKzOLI2YtzG6qHAJZ6UjTSpcJZtsrx/AhqcsGBhM92xCmYPQoEIlJjiowKS3T
pNFQK8KLxHjsYl+7cp0G+DIkgygV4HvyCvyDlh2UKNnPuy4Q6k/E/NDeKDT+dSKT
jLkr0qL5j7/64WjxhRHrB/EnwlVOsKsDl3QvjP6noOcvD1XcPp1d4APXaKsSaMSK
eLzW1VYcGVloQTx/fPx6wsoccgGx/r21qqQCJX8kq+25wgdlWjrLaqjOlb1zosih
xeMsOEC5Q91i7tJj56wKfkXzgw82D1aQgl5uTiTjdcTjBHuHfQNSxz1DLQkFESPr
JF5jhIdFT6rqT/TNH8by/blNf6it2DsA0DtOrDYWsbIg33RsFVqjbao9Q01sZfIK
wyaJbQj+tE8qOy9FX/JUrURYH+kEINznN75HCPY6jBHHAUIwt/CqvWO3To2qPyUU
7h8HzC/yxAmIHH4B5PKh+emrj4eqY/oVDl+bpl1FiOxUGj9nBbww2MHNOxBq9v1Y
jeL1Q87SK/s27gi7cVT1Oz0O+tCgfKk6TY/gBEpeWaUBq46VNC0ek0Qy0DFJSBIr
vb2FcISG+jA4qUQpOVZY4Ip0hKwCCXWwOl7SkbZhbUUZbrrd4wj/H8hfK2AO9Iai
Mzn7PJumOA8XGeJnYGE07DoXOOc72VKAy1Dv9Zi2lfxuP4LlfiBkEr3/Djnf0HWy
1lgMM/CuXrEf7Xicuq/XKnWT0WC7KIWdCignkuMP4I4j6mc6RkqCoXi7GrckVAem
WIrnz8F0eLiQsahn+EjH3wveogXDqZtOjHbT2hlzCL1/P8R3QlSy5Op21AzaO0dX
lZnWGZ4g6jGF2YVy5/XGTnqf/AodfJFomGxNr3mlFTrC0HnQ+Z2b6Th0zsYgNr0o
IZNLhZ7pyKVIsiKC18uKZrkzupE6/D2Emvc6nbz6LnwjSA7q7OS9EfRSe4Ocwhik
A4rQve7EOl631TU4/QVRGM6jUJGZ70+SDD77BEaRokIVCU4e3csl365Kit97lEOt
Rjv1zhZ/xEtH/pmEsBgCSSekoWHsoNeHHrzvuLdWgPu2JAcv6C+Z1V3sCTRmg1GD
WG0Zj1/DVPxJMD1jAbRCRVOWjcMtCVbvGO3lCQXCI5IOkoYaIaCohI/+85nP0CGz
8cEGJTqgMlO1wU9HPdmIUMz7nnCQFtU/PaRFF1wCpYNr3cNzV9rJ9ySSMJIBieJ5
7N1NXuGd5JM6SKyARfYQQ6uYjo6AAyx1m1/ma4VKdSN4QiIal0Q8driTYJ0Bp2Bk
c6/zV+YSHsbzHIzTYs2ubMZEtjY6i/iVKGSkYQC3JwokYhSlK9icDFqoof1lIzqT
JzPCtLfEnI3MY9pSk6Dos98XHhcj9eeL87b9x6V92oSxSpoeyqLUuVh28hOLpsIc
U9qKN4WGi0H/DdFw8grrbESuCV+ALEi7u51oMTohPRVMX22ygNql+B9JOsXs/GbH
r/n/1/DwiJ1L0gcREEkZH9McDPbxkkXvZ0LSlcU6VhgMjKwAK1y0cCF3DDRcZwGd
VyLz2vCUnr9+TaZW/tX7YBJbGvDbmvkDuCAaYUPWt9tsq2iCTrQfi//mx7KDXXF3
MmwSlraLRCQ3cvfKdunuCMg/I0a0oubFPIdluF5oo5TyVxR3yh6uPDcuTPTacvc7
wpIiAN9tGikCdnXzeozyB/gxwjnXwSMdMwI1U0uiX0RjSvcW/nOXoxnU+4+FdfSM
MM9a5N7o0PT+EJzZtxSmq4Pm9Hsi2WwxmpYkmcT+oYP0PizZnHqJsYEbZYFvsofk
X/g4l+vbnkDrKcW1E/Vmsao30aqQPe0n9PjRCckYwXvGZbiDuPWPs33K4NlWSUYW
mur1fSUpgqeIpu2OtDTq7QunzdnjnWOa9bs+PMFpGGqck0WNLRCPBa7NPPXMwM8P
5HVI8+ViL5CcGib7nmkFGiKz0JoKrPPigC/kUJN9S3LYTr6AHXLKi7m7dQjlx0Og
vlCOBamd2BaFC9AA6oLLqcipSICKxQFAY57TAROVi/4zXCa88dUgZ5VQuQrsa7a4
KqVQhNPr8mKvvYoSYx+ae6+rvnrDqsL2tDgJYU9H5iYHjU/mzEjUWyHbC4Bk0rHc
Ok00Nq6MOHdJL7ixAMdS330uuB6E5LaNeOA8ONGnPrvUyL2LbKi9ciYGyUD4+pC3
Pc3Ul9E6CLHseX8L/EWML2bqdQ2cAD2Qn/sb5w1Szd7VF1AJJJZwwZyDNpJpTzKs
IyczomQrjZL9ERY/FGqxzOdrt54bqc9iUplXhFSLa3VxX3avIVfVICtQdWTMiOab
hf4AIeyGJ5Wdw8XWLtaeB/z6JhX1FslGGyQ1fw6u3O16YW0R+ZC9Mjg6IdU0UGtO
cVthjgf5fB8jc3xAlyjYw2rrq//LKMrf69j6j03xXYK+pUkLTMZlbcanOWlTa+Qu
/67pPmmfDUsSEjG9kHdHacPU7HVKdamKsgKoyLvzkKXXjY6d8OVM3IqKposshSGZ
IuLkhRBNHNOi8QeI+q1UFKgLBxGKfoq0mCVU3SF5f2EhBHGkiZppLnEfESBb40x2
Fa76EphtA8bC1ro6cvOu9YBUsFKGcsTXDLlGkMFLvWIFQrOfXW/AgC48XEX02Qsk
2MF+09KS4CeeE2HSXFJFN1QLWkggupZCgP2g5qPLV7oQdWAcL3mBLXLcchlXsOdo
UwjRmGMd2HVnFN0PQRg2wVlGYR/+w8O9d9zaW9CbuMl9GUbHzxZNLmHBNycjpmWT
6V/jbYNeXhOt+eUg+UR/h2kA7jao/ib/wOED6GbNhdIOahXFbFrXsWuE5AiVsPBU
6v3utv+GMYFvEeUsmjdpMOUtOuqdcd7OVfTgvBepl0iIB42vofm+A2qTi2rJg2qm
jYqh8ZgGsmx5HjdFndmfl2zi2XE7QiWlKGgNY4rqRaZXm9etizVZ/fmPHbEnIXdS
UuW+KMzy0B4fgjLOfR9v5kZC9XReiWfgVDw1fUlA2VW9TR5ROVFldNF6tiNpave7
lnkmGSyzfeTvLjFrg/tVPALT5/9yXgW2cYGWtB0LPgL6ULJoMwPauGySb5zrmj2H
aXaLm+ZX70ua4Fupq87tl+c4LtOYv11WgNUxy5Kr6SvwDrd9gpnzl+rADCwW1xpR
Bujd2HOJfVjMKNHXeu4Qik3G+NAETNpB+PYMCmH7QGyQtYUUuM36zrMZytQN5KwY
Lc1NrURb8o41ORQdPpmPQlJ8dWLhBxqxN/NEEN4UwF2VU52KaErFBVqMgwx1wtmb
dBlBNpXHJX9k8Qq1oHia8X6p5CX5YMWHSGijggV0/HlLNClIvh+RwghjUkoQMn1w
tCYf2S4Ty75V5GYcQasd5mHYMjj925WcOcZHmgW0vHje2lMXpvGdem9YIZo7+7Bn
UpJDAXvlzL8BlAXQJyS11jWpYHD524GSH3zbf4uEkAhqTKhXpsXP7wozILfPDAF2
a7Q0bgJUzvPl9vrObf04gSihrn6HvI0NNcyvL4p1uS0+2WRqTCImhyKMUVgYkmgZ
pgp1BFQ8ZeFCbKOeAPP+fTRykpW+CF7y+xpFQdFLacjQYNugAah2J9uLw2EZo7pO
q8vPyTvDujqR9nO+Ngmx4jRKoa1mIuoq4uRG5Ff3t/Yg3R2c6wbObFyc7Xk8liA8
c6E/5HxWOdxZ8wEc0Ge8t/Xpb/RNO5FOXVqNOi/KGZb7PYljBF7JmOFUCmiIKejC
nEjC3YefLyi3FzrURORYAX06TY+MiobIlv1lTYIbu3e7i2NCKnlhTk7b5Kk9dLrZ
d2TgLt9e4fuuP6JFF0TdjaPKLMGEReAa6YZJ1ZOGw4TvGxqPV9LT94EqNRbOvqK2
7L21j/80/g+5ubJ38lxl9ZbYnNfLwHfn7gnY1UqJChnEYwcAdM8KL8ZRqzqajS1v
1ISuv4eT56j0cMkcWDPIREzwsMhFVw9updYCkgIzKb+pqM3xcwqkid0UoSZOpbzn
2P67y/EH3vqXFAmIAn4cc+iZ2U98/UOmexKXONfwtp/O16zTbdCKKQbetsneMDXQ
YylXh1AtxbH5/Ge8o9yxyXuOl2CjzU5X41gzyAWfPEjH8hserEz6KKv/calnUjJR
KGiHIAj/EB38Xc98+6UZYZGFdQMOeDmbQHIuQ3WrbfvmcwUfqSbsBlv/Z1LTZel6
jZAjeDNFQC1lUTe1iCU9r30InZglO7okFWXybysGoJKzElkXSTUaf10yNDEbXcd4
trv0btfPvGdHIBbIM23c0KFBnH0tw6Ghww/jnUXF/1/C3fZZMZHTjMKTdyQh0lnY
7NlIufACKlA2ZhEpyP8BIurmeY91n0sy/fX6KcO2nKfK4/N49K9idS7ibh4f9dCZ
onjRodJR6/HAka0puIK8itMP+LoEdBO5mCCAWAa0dgWhguIzu33Oot/bYZPot6AR
MAWEGUDSmhfrs4HtOvQFTqchoMIPZfYM0UFkcz0lTr2yqSEgvbV7t7/2pw9ejzli
wc7RtXriWwCUlvTBV4+4Sr/Ud6JXeH91t1f1Stelquc/37quxXTZ1rAc8hNks5V1
TnOMXIFJ9aMjqSAP+ujO3A9KY/SaZjEcU0F+i/NNoNa4ElhYVAiCHplbvhRbbVJK
HNUy8of+lV9XozDJpRau3taRRP8gjfedyo73uJRon8CqS/roy2gOGFev0QGT0pR2
3FgUOtVAaQDRBCGfhRcCCGhVwrM5CBllobTOiX12EvSSe0Xjxc0haqajq42Nwekr
sYluhPYXCmCC15Gsd25K478FcJDDk7AT8HB6+OzBDFvBfwi3nf7CT8rV7C/pbCL1
6fVmhGIFUfEgwO+pjY3FgmvTk9vrlT8xwUlaXyBdqZ53H6aSlHn47EYVPMF+YmmS
Tt+jrU7l1Y9VD2jPgHhtu5JFO/Ub9X8Oew5GpvGlPfid3edky0bqyrdGRAFYsf44
n3H9sA4tOcfOpCAeTwoC3dKn6vLmmC2uDCGL4bDGaMTmah3TBNCpaeOOSx8IyEd+
CWvE0zpU8hGtX8UXn9eBkN0+EjPuVwe0zQzFk15hU28aXozt773OHa/Ulz4uxfrs
Z1dzweyrK3uwmO1/GA8gFzxS3uzQ2Jd7tjtuxd0dCbSQ3AVJNPvEGq6LsyTrc2uk
wu9ryj1FCTJFSueY7i5D6zweuMiCEnwyoD7bXFk3I6gPEh3ct7+rVH3UwiErqA4V
1zYN3WhvdA0M4x7sPCZt74IbPp19/aOSWo2cI+ctmZbn9/+WoMMeLSRf11PVrJq+
khlTJJphJYGFZZ7qYnBkAy+0pqmyoO1JiX+EJRGwcK7WUzlKn7V/z38o2/axUSca
aOuaPeM9/P+u1L7aKep+8cyVCe+kh6EWsyOW+og8rQLrLlQ9CTgf0hgQWrFWITpr
1OoRG14JtSaWS86oHtZIs15mLgYlNZydOipCfNUzW+gjfP0VE2tPvp6DyBfBcNVE
wio/Pu+nJhJ5/CgOFYzbhyGa0fJX1xTHPDp/Vy8LtCnVWsPXTnZAqXjx1+9vEQkY
gtDvlYEBzR90Eov1Qk9Se8VqzPGh0eVOxJweZYz5wNDva9qWfQ0cHsu1YJGMvi1D
v9NSbze/CBLlG7sX/xm8SmG5/8zVVTeZXVf265jw+YbeiulYgxyBgZEULqtKrTDG
M8au8hBc7lYgK5Bu04OZoe0UdQ+8P5FMBBujL3iPho7sGE4vtmJnt71Lq2hz9beT
lSvaYjPpKNafPrO+9E1cERrcs9yoT0xGWGWF6Mxy5D0pppU7ZVe+8mpoIvbXHH9R
XJVJBj4sdErTbyMrI4JRVesGDopBS2sZhkXMaoK2JkZb2s/7jnS7iokDNVz7vjfs
KUjPyJKHx28igFC6/hPB7irir8YVtFlpMC+mPP3oDnNBTWfyA1JzJL2uuF0UUGe+
YxuvAsEM/Si+dydGSQBT6OE40Jf+k2t0oDd9oKVEhr4+fA6Z8bxOTJS4Ti0RZwvK
0x1CpTISvxcDrIdPWhqrwoyNjJCJIzKRv3olYriL2MdUjRXHPqpsovBMQAgRTvdl
X7ciWnh61Natflng5usUtGhS7SwLlXXIVk8V8B4x8Vb6McZ3OHF1d0wSWc/LDuY8
q3DvBnUKqpOXIxXI6UjgdERj7RhmbkkAoP/nU7YqidobsB2pe3dq8mrFlpCtTqla
Y0f0+r0de2iqS4pL+tk0cbbPCR5hg3ly1mBa/4x+dyta8Dm18yoxsFfXj88NucUK
k0A+1ipZwXi61mWE6NmYpQeD59cg6C0/FoQl8pxqVnBcrGcIhT1PYCoVueKUNBMp
vvb9nYQcGHI/KdfkrvKghLOMVCndR35SJuglvdmjlEuFb64AkkPCQGahrKj9I6mg
NWM4WctkeR6xpE5BOe113IVJJk8Bk8YoD1dmLwEnT+t61gP+QzQFG1M+hqcTZp6f
mMqPjeHq0abm3kIXxgsY30EfZTuE6LvFt3FwUBrkK10N3oV4bk/ZqcDzW2wiGeB/
a85M4iqoLcD2g3Rg38HvL0C+ELxdaMhL1+OsS8RrKCf/6A7Gy/++xT35JksmABP1
kubo/OrooejKMvE+lOIC1ZbVEGMx4VLbQNNWSGwpVeTOl2vYLBOWV/lcbuYjDym/
BpGOmlf11U3MjrxTBr9rIn1GPmcxjqQnWMuxOPf6wwr9nSeHN3ks9algYGS3eXeC
Lq6PR5K0mof9JNLP5iQYGZ2/vqp51Z1yIgbUcpVtLroP/YzjQyULxGJMSBEuKaqV
fVrTbFAkRUGrybCjZUSfzRN2vwmxEZ4RAxk3Ne8JDD3qPoPOcpw7/57dfUA+enGm
PfYQe1N5TPTpYMLAysZhjmgWCOmKC9RC+/+DG93YcHtxC92EhOcWbI4IDKojCgb8
Dwzuz6Sz1/7Drx37lOdvD19jj22piDKt6+QcckD8PljghhAr//06cDEaP0jrAOAE
HGivyXeO3A79NIJMTN42haJbblbHfCQspMuU9tvPcTFOMXA+FYBeAk69J3muzzmY
sZ8L5RAN1s/ohybs/cgya1gdH8FXNexuUxgzsksh/6QOoTNUQegYFiN/qqCb1wDK
Vx6G1yZ8oWL8lLjWHg5kFLYclc2svqD6L0iy3dgb6o1/+TKgCj98DODDjzsyJua/
+ieUkLGwDrmIoBrNPE1cEzsgl+ZYYFE4ZO4VYxWVH4kq7qX90CzqJZZDDDc5pLUK
S0QoK5h1AA3a2GQee82eBfua6vQ9Ld3UiGjT7jQ3EBMHxquL95glippCFjbNN/g/
aNLA3P3OjHZlaIQncpbN9g2FOZTt6OsIoqTFc024fOWacDPJq/xiIrivCLXuUcem
zAbY4cVbuW+ZFS5bE+eDzT08N08y2we+vQA1VXZREs/+oAO/3uiTpLz5oHgEs+gb
StJc85j/4wGafjJJ4NgXBZj1kxCTiI3szkhxEBGlSaY8q5YbwDc0TnJMZQfh0G1q
48li6+ZI4kCkHTRkXTU3lar1acxrTVjGLbyzcxgEo12LV1rPF4jsFXX1RhtDZ28r
gN98uMmsgxzan5eID0ZGHBbBuSa4vg48nK1QbwwPLQEtbMps7q+a+IIYoABT1U91
UDRnsfGx8sWbAbCJBR55ZJyPoeI4PG7oNM9tfD8zqTZm7Fai0Kuvj5XdZlkzn1Sp
ehlW+lnoZxjP3PvNUC5BJmpH/jWJO3taav42CsusYrcgEXbJQp7WpViUTTQ2XcaJ
zhFLeyQvU99kc0QLgpLlpcC7TukzorqyyoUumh9ZX6NPx0Yl6pMlujcomkOoRUSh
2KvVgdwgA99Xyffj0iMPXki/wAMsElKIwm2c2KMVEn23AqSIhHevweh3d2OtqpFU
ikZuai6k8nAsQY4DS/9f5TAtSoliRTy6G5z2gtjxiIoZgPqyQVAzFuq2RiPw0Fxe
37U7cWvPp+1CsdRQqMgoZcyQHUCur54EmzRHrt1A2nHC90kDcsm3hxK4K8uVdA9x
DyGBt5VOGfWAYqMk9rD0A2I4fQDX7FrIZeLDjW2gHDleIMvUGkWZIJnMajXzaRi9
tEcS01Ypks34zwNtvDOOrxiKOnhMeGBH21ORHIhd9kiD5bPGHeWbBWp2RdnD8jwQ
ueoe8a1AiAbL1v3cJlhr2yvXYFmc/dYeiyQRBTE62hEW8/d2PNWzEdQZVNk8+zH7
rtljFgr23r5YhP68hyc60o0o4z6xIl1zz7sfnZLbzivFjNzfaqX69u3hrhM6yOm2
MCB5imcaertGAjTmRjkdyMKskr9DDJ0Fhh+CHj1LSrym7o14licUXStTPZB+5pIA
tHAGrujhxD3vCOcWJX36wMYFWxyXnWQwUMMzWguDCeo/wvNvJvLGlpQ9K4LopLDA
MywqFFnVXRnI/XYnGYBX70U2D5v7ya+xChmX4z3kMNQr43uB0p9W04txLMdr8dBN
Q7a6gT6BQfXqADZGuTVl3ewyZ2pxCsAIHDLW1Az5n+jMehaKExJ7xcUBSr2Oe7B9
jyZSUUnZUeVPRCp6qSTOobyt5c3SNzhSdJrLPQCoIKSegzDaSkwZoDjDzHTphzBm
d648USjwYMcwDmZ3kZRQP+Yq43wIpuILIJbftsqnEoPIE6+EocpMp4QUgWoi1jSJ
bHKdA2jngrN8e5pUOuDiQ484YRkzVLMw5M0TAyWKNwD4/mAoOyp6gLkYC2W4Gjxy
C82OTivuibIByZbNgcf7JBF/yr1aE+2TaEFvwkJu+ueFpC3LDNPO5CfqsOBFyfBK
ofl4YfP7trbhXbx4SaegJ2+23AmwO8IoxZDtOvlwDL56pI+VQHyo+x/3hTX09CNu
4LA0GoFliQ+SqxTElndCX0Ij7h52wf26DUfD2gf7BM7MwXs6gMjYzy+VfI1pVp5K
wTu5Wk/cBx961RUlbqNETdG7lDbrLhE+cb0UfmJZ0in/RiQlMCe+k5lbvznoLjkt
mRiSEmd5LvmoqohuHMbwUvgKHiLSLlWbqSNsOBVXQ8u/QKTM0Z4i6MfcJLIKj+Cq
NbCn9Wyda/zVufBSRWSoqOfZ7PaRG+hzRa8xjxFpJzjpbJSpHn3dbOr3REQPLDLi
ONnbOvRdKOJL+HzbdDM1pAsQwE9D98dCBFYtD/R98YdfiwV9Ydg+p0rk/v+93Hex
nvDiyDdmKNEJAInkjYg8FvA+Fat5N2YoVR+7Gi/6qM6j4J1T8N7bEhXadjCUR5+R
AjhDydaL4CZqtFolNyBaP8gqlWHgMNwjN1IQAZgJZRXmI9bXGdLgwwUiA4AxpBpX
iGj+oaFq5ID1S5EhQ+Cmue9HQeqHZTPLnB8e9jSdBYJtKtMNxi4QS/qIFCme6W0W
gEu52AaktliHDO3KDvAheRjxlGqj/2Ek/PwqwTNfMwGrI9BwKp8JVSG1YCOVcUob
JXfWDJJwkFjryLd3d8qIt8A6HCigOq3QNY6HXtKFauX99TUDvAlFoHsXf/1DJUJE
OXVkZFPLjIOco4CV53hVdWMr0vTl/WbB67ZOFXIPdpP61fBF9dSrrxH0acbOlOjq
qyX+H2cy8m/XNNkfdIpuh5HTm982N4R1c/jI0pyDxz6Y8fLLkuHKIsAA7pJYNOHA
tgSLuhfhbXYKi6Y8QeCu6pMvMcGLedh3v2pw4aPlShws1vKyBOILOGvGc0CZpyou
lq97wxmGd4Pmuuk/z27fM0E3A92PNeFwgcCGzCI0h6XIihOp1c85OHPGSWtl/vRl
f8F8W8Vw635Kf+xSO8Frz9DqPVkwfQCPRz6duJTD0I8Mnb+f9KGMuuSX27PPir+5
0ho99ImXFZKzRVOzUkykOG4pGuHeJv1rlOv0P1EKXOKgOxtxPxYyJRJ/yyS9jf/1
zYm/ZkJK2PTTP/Ik4CeHcz4LZYSrlcYwDKFOceGYB/wgThtZBfS6EgcSa64Lpy/x
v9B0bwsL2kvuzk8MEAh9YjaxwQnJ7RBtrRrxn2WlhhbRm0ukFQcRgFqn1E+pVPRh
MoIkcZvuvqBoVYCNLeGrjw1HjFFsTAetDLfw+49aUVfHoVFLFYmPX/pjqsTCX2Ui
fpA2scR597tQnjFBggDG2BXm3u+C4r5oCW9lIE0DdLnCaI1ZZ4fUEAlT7hdD1uKh
salv4N4gmDyfoDLBwyf/HFt5YfVCgsNMUSXdXGehKatcHwZWED88MAlAmFK4JpxP
1kqY5M8v2K7ABE6thFSiwO1ZQ/p8SMMssGvW0dIKATivi4kq5G52qq657Szc72VO
Jt4zXVXEgL7bkNPddm7PEYRS00WDrXlIVm7PEoDzhwkG8D3SIAAHTwErzAlcxs/o
Er1hwOjzGh7MTL73D/X49mU0YW3EPsNuKUVBIZwNARp7A5RBXd7Na4NlG21MKmgP
JPha0VBSlc8JPlF0VL0iLeMXE84yb1uWdOX8vfe+OwZlkzUn35fFwZ+/52keXIfe
XE6wUpNRpp1LVy7MrKO7+zvR5e6W69R3tFzcgMZTIZd49i+naLXBoVCUOuqpnoJD
KCEYC1eI7QDx66l/O0BdkDc/wsJMoppR4APflqjqlVp0gdtmXlAX6YnwMpLh1uEM
eKMlXchQcCzmYn7jZbF6zQRsPXOXUodIsHX7UapaDKPLwdjpkNwmUUhDC+ZXAEuV
yZoWSgePMrhyl8ozINICtA92QVOljGRUn/UUpXMOL5LTaVRb3kbUtVAnCEivR3Yl
HAGDIBTRC4uevxJeQx5RxJ0+9tapKD0PJNplBj9x+g/ObHHdHyB47BynnjGgV7tB
EkQCiAb5nnFS590E9Hk/gxewiXAmhZzqAAeBDg37iWXlRCwVB7EnIhN756iij5iQ
APKJZlv9lGUxV8CTdMuA9EPCWWfaN2vaftjda/euonMUHXyvdzqwrTfPa39jug8K
37/GZ6CnrkT4ldxzgBXwrnNpKivFrB95Nfp7fNF46wzWuNvfoJntiR09fyGcxH8d
AyWDcSpXfuojw/k2YaLsE/EffiWzIFVVu/GQoZTDhwX/6Qn3Sm5LtDm67d+YJ7Hs
Qrw4FHfm129D62WDxX+8v+FbUyUj+hPvXKCWz+BhXybdpesGYFqxPBZdBTFIlr8z
LLfjAXv5zfznoJGShVlTyoWh90iaYr6mhQkcTFtv1oDIaMT9Iv//g/FHU6O+xIxL
+2oeV9rMYPDXY2JefhspmC2q4uu+o+xk9/4ABPFQuCRCug1MS3A1fai9LnTpNMxz
5oBFRIC1/rqSxMgBr58GGgWg86/31Ed0gWd4tvAaradyydPJ2AHbGTXLjWkqse3V
CeXgsoCAibE0ACnGxceraFwGcV5z/J3mtLjqRlBuPAKKcInymnmPT/oe1BQtn6Yd
oucsp/4m49Lxo1CCzTPTF7oEHdkZ2AKeiT0tTkQzpnJ7JR+PuA1IANwTHUKVjvf6
vJ3TzmRirah0rFynvCax4769Rhv68KcRrRzztEIPbndpu8f+tNZbaPZCUqswCJPd
PyMZGKkd/oPub6Lu0RWuseWSc+i9A441S5GTJQOKppxwHZPeB0xbgzubDEsuHJmy
BvMudI15oyOJpy8ARS+5jWdDdBzUDUgoR4uyu5vY0fSTofWPP8fAcUfT1Gvnn8qP
Yib6LTdVsGC4UqiCmal5MggU0vVVEk9ksZKl7KR76V/dM1T/A4qa9W1qdyuZdnZf
SeTV8eUE1cjgyYW1j3v2KwNFFEgcDDRzng94HIBgJO2w8YBRXR9rDg2hEqNzQNio
ekPoGpPSD2EKoznBTOCaHoRCuXCzFKXcrmFSXJ2f+y30KyYgThjHdZMw/q9C61tO
VzPMtdKBoiqWLDDLYAOq+9oLdlxcOFhd5eKcxEOdSQ5j2CEm1cvE7sPH3+zsOPFn
f3db0JU/fXHhFcdhHdsD4J5GEDNJhvo99VoWLV4sdo+IWy2FBTps051lj49cpaV1
4C+XgoPKwFCcgMIyB4zqAoGu91Kh30WJH178tMty0h4dqspiSLI0pwVCQENmXM5F
e+UC33sG+nzxxRgbiPLcCjqWzOQ84zxgeP6F7K0YIMRnPgG7rZha/2P6C4tHHvip
/R+PJ/f6Qd1sK2QANXz8yI/GXGTW3KS0cQrk4Hkipz+ZPRzI+OYtiMudv+LuloA4
EsXc6EgWA0L3uiVBem+OP/ylj/Pk3fXzfXnwxxdXQ/i1V00dtFbbNuCFCF0BhDoS
U6SbWbeukI3uo+8RHuX7le1Ix27oaPmufTDZXubfKSbUGCsqd8N82HgV5j02bcN9
zHSohdSbdaYxvazQoD3w86rVytjZ5EXerTBg0piqoX632nR428WhgaB6dcJFuv+g
BrzuvCe9+XhSw7vlx0U5jY7Uf2gZWV6Eg7Ognbwl/+nINgQgJCHGne2LArK9rifm
3PLaacnDeJw+t+B6BMJLqb8diUM/Sp5nBKwmu6lM40rqMpf9xqUIkAuN+S/Gix0N
JnexIf95yS+kMkp1i9+mUqnnpGx7bYxPgwQ8+95aqswq6rX3Tm/jSMhV8mwko8hq
5EDSDCPDNynsQT9OutrG4evgYj5SBl5gbiio6ztslnVVrazDZ26r8u7JqVD0ppNv
Opsnf4YRWDJSZPcuC1rtLqtToohB6VU3u8JiG+YGGSU6UyEU2AMIEzZiBR085Glg
kOpydPkjBmmO0P1n8fJxdhCTZha0S/uv6SnN8nsrTTuk+xFRGgIjkI2D3Rdd3ty0
bYaqu+sOKJBT1lkaBK0hVwtUIHYDx11wtbActSV1CZisYa57NuTGtddnM/UtDyUY
AtzQyTqKoswUpc5KDGFecMeu+2aEl8TTyVMErloDThvi2pxL6MsiQC4RomEtFe2t
YLCG8CY9+rRKCfctQeBBnxpWIVJzwbBx/HvPyRqahMDFg5Bn5rgWRLIFAjcaObrN
C9faHGuXfHufFtvcvrJYqEZ9u+VspmJPqpp0LpDsHNvdnCgCY9JyRIZMrFUfSZLl
QmyQRwhlQA5x4p9m3cFdbvj3eyBGI4PEtz0SWy0JacpH1Gh4w3jELE6lH+/beg5o
/nYpbYI2/WYKnJiOh/EM9nBqbM4/IQht04cjLxXMhecfK6aFY/PTBDq9UmDh/S0/
IO2VT2vJ5/eXbZ4/yDMnhCS1Z9+GSJUsYArBnvcBWqir1nfaX6GWn5AcyDglp3z+
pALD2NBmV6KxcYmai1eIrAzteb5YPd4OpXoRTwYaJ/nGrEvcfHxgZPO77S7XAP0m
21bO1LBQiBBpoi1+BkRNygLXUxgbzMKjpvTKEFMit8SPZfswacDUyltcN/5SwZIZ
3d3X9S8OUbRXbfTr3MfokulorQm8NrJhhENnf32/CP38O7uuuJtuHHyYHV0VZ4Kj
IXseegd+KWqfnHUPkAFsIgISprSv4MTy0COTvbbskr0qko5XFMTGeoOhtZyrrqMj
HlIvM/bhgyE4/Vv0qvJU79QW0viLlusG++7vCI062k7HpoH8mPGXvmqU587R/PmA
99d+hRRiojcCzyGd3a7PJmub54k/u5CZxWgNESvXxB3p55GfWAK22kQ/8dsHT1kv
3KNJ1LVwz72LH26hTjmp+bLRFuP0CJCEe3uL8/IwNUe20a/fFvTZrwGIQFGR+gcT
frJDFk79ZD0KHRU8GmHA+2tMdOBjlEnh1FZ2DQ4x1djY/Ws/OIvaFV/25p1MQJtD
EUQq1UF1T71bPqtdXSgu4gMuDAUWaweEU5IG+uPvH3X6JJZ82qAhJNTdmWHrjqS5
5GOSX7UGbAzeBIDw5t0Hpi0K+KaYcMlFJXWyYeIeDvrzeKXQv47vQ56Cz3ZNi/ep
duhs2lkCEd+6ioM5Uu5o7AtPkoMs1jWqJG7O3RA1Dwh2Bxb4Rs5WHBsUXuEZjMAC
eZhn48e6iYGESZExJhiGoWLY3hgAlzTkLe7lNbG8+KLvv7bE4X/RBAHp8CD28kBl
HqOSbKiRyQlq00yMHCHT2B0s2MlLx1GYdsE0cmYa9ayNk1XEB3ClOYFy14hsFChr
r6XhJx0OBdvoX1Mg6rEADDdy9tJ1ENyCNsVNJ/Wh0SCy108sv7kmmTVwDaf4gMcy
iGtqgqhYV9UKlwKehVJPRsy8Z5p+h6HYIEcIvFSNGC89oHw6iPeJg/H5+iliL4Ux
ZtLlpVVJi6q0mhr3rJwG5tcux0S0LMjWgfKaZdAleXDKLYCCZqdNuJVUmb+Ay1M9
30IhOJDhZPqHlPRvqhWSXXc+gej3oL13H1oFjOeGreIQVTAW1dH/3nXBYuzLzT4U
ZglDx8SwMBu18q9b6TbHnCiGGmHe9fAFfzxK2TH5S8Iiae1a9Ym9pzcQMMP+Q1LV
jqcGpt8fHoI9cDTBYehsedrnua4oZ67Me7LX3WGMR17do4OTlYkf+21KQ/16tQPC
skpOc0KUuMTAaqgFSdr1FUzbv5XcqVwt0nMTvtSTpbuqq5k0BjvcIu0nrs1c+Rif
qO147RbFDW43jU93q8FlYucZT67qo2ioBlkX/HDW3NEjvxwP9Pyz1y2LgqNvdJYA
BSwLModZ9+EeKQPXaN58IH08Dkg17Smrx6OlzHsA5UReSetdejXx3upNpyVGu+Ct
6gPSWhwJ1RXlYHkXXHq+vaCD/aj2HlRWWcqT4y26K5oHLGNVnPN+Ngow+uZVJrDs
vXZ79nVaOdB8lvjwCYHimREnsyTg8UFsK6qLNx6+OT4gnauAer8DrifKcqLmEU4f
z4UwabYYrPiDlXx76dVRsBwk70ffJrZCTwgIYbnWBwSW65QCA6oA5VSt8d2a5cTU
/iLx7p+c2B791KoKKcBveiLuoYLjJwA0wR7esnoYrpXCm11i8vNo3uyFX1sgivSF
pRleAEwCJO9AoDLiB+wemonLpgeA1FHrUJjDbzGbg8k4fJxhk45iclt1lsHVdjbh
7Fuc4gFZpIJfx8YxYh2NvuKMcrqv1DFStqnBmsNWalX/sRtyys5OeKWCd6dmIKlH
sjuCVYEkNeOT4nXEqyyoQEl7qz1/p+p4wq35w5Ht4Q2HtoBinZ7yVjCFyWMcJxI+
Ci1gRZq+/A142zq89TFQg1t6UvFMrERyiW/aVBupCs96w+klqjfVYK6lB5Zg3fCN
m7ayWllejIP/EifSCnIM2RHWtb75P8Pqyi9Rig+Z1cemDtbhngf//TgnPnOXZlTK
GCXKO7pj6GuM5J0BUTRhXQUA2I3Oe3KvoQnuebxkSJZcLUzKim+hajE93vKMVHEk
l9UTxNU8lWipJHUYXX+5485Dj6IKjPG5vdqmacMq9kbMBHnbOnmD2t585aCy5fjx
RuiuB1AL24UKHh1qQdWTBMDamlWC4Uimdp2vmYOAxnwFVZ2QSZx1WbxsWWA4aPvW
I/RuMY9hh8WVul5XcH+D/VwrfEg/ii+VpY3he2VnoHedDnIBJ0b/ShwDcQF2Houv
vN1r1LdBfN4HEFkAIAAbH8LCoE7YCuRHQiRMMPRhXySzb7ePL4seyOgiwKjzNKxK
+wlqglYM8LMeHgs3VMlZl5lPWt72daZcUkEdzhBmvZkbFley4QPFRt7frVSA+aCF
900zugIJgewPoJvoJZJxsFHIZVYSUGf8edptBT7+8EG+PCP8rVCKi1V7XylRdK8E
BV7Fmk6Q35TunWCmemapDen4J8eMw6oXLixJsWZHZydTqmXYVdEjDJd/c5sd2RuG
pJzeCbrHh6gJUXYG+EjM+iQgcvVa2t7rCMlKLYOn/rTYn4OcsePa/4BJRZ1d7XwG
eaumGQW5qJikAWnhounBjNQeDou0fKSwjFUoNU3/5WgdHPEB+HIP4jE6R0LTV5ZF
kNdcOSxqKvlIt+2iuWFi6/dWX2K8pyeg7MOyU6HFoSA+Z8d/5zpf1klI3O+s6uaY
Xnheb86u5et/UrK16HNrHvLFCeQA9EFtKeyL/KFJsxRxUoBF3z2bHP1QyZV0OZ1D
G5ikvaOhVFafGYYJmjCtiwKRSE/u125tGf1K+0XKRcwv7pFGieDAnnXEqA97+YVO
DX4qYa5fzDN+aQDA7hAoild8hWlqbiNPTOenGTo+teZ1xJCDM+RNXfuj3xj1tR+F
WSNsI705d+oWuPrT209pGAu75dA29sFpbuDDzuYw5b98oWOTdDVVRnjJWpd5d967
Qg9oKYs4LsIuSOPe200yRiSuJ2xJ4Hmu0ZgP2lGfJy7wRsW8Lerni/sm6our/yf4
nQPZs6AbbaLFeC1MjMXnhK5jJpiOkq4qMZ0ctbA3HM9+KQrQUjHyKPQFviwxeuzd
vmYHX8qmMszIAZSiDM2gF5Xrf+CPQofbDVkWV7YRSUyCkVD8Q+jTt3J6WUd/Fdcv
v4O3HYPB81P5yaF9/LSm1miDDroGDKeuIufgBAO5jiFnyo+xtgSbJbnw/nj5FSSq
Y0ZfK7HDvziOy0YyLvwd6uSiVGQkz6oY9YvMqETbrBBGg8q6A5bxinqJiOr9V0Dn
phXMOEh3jmOwAeodDSN8nVaGmy4OJmYADX89h8PGyMpA3MLNKCg4TspQwxgRzyED
N0kwBem41L1/A44wwOZw1Igv/jM7wzRFNGYdTDCYwpQi/FaFCwILFFjzOJjtCbfK
JLNQqv3n2V6PU9B84k/kuzqBMnqmL7bqBZTjvbp14FtwIj9zFgq5Aq9Gk9iyOvCG
sC9UfXmQg3DN/rn5rE1a2BC4i6pZZ3opyx+qTo4IGRBhP/6ftBpzyO7br8DTxb5a
U0cTQXJKRKMBp7XLgFJ355EH9YUELVoKpuNAIytYC8T8A6F/Q/SG6OmDk+F4jm0z
1ZL7jMnq2LQ/AJlIpI73LXAtHwP07HGxTHIsobrs57U2pwpmGa8J4S2bi5ok0TqJ
lc92b5v92vtubmnj/gf3xUpqVBMPQ2z+KsZWskHNk7cL6IAW64Rsy6Bg4iDxEkBn
u9aLzvlYBMEiW+JTktNsenzDIkywRMFxwvhAMfk0S/kKsCUCV3yYOzJqKTbVrPrW
nojGo8qehRbYxy7ACC4XPhp8wqiNamNl/euqeq9bJvOpGpFjlyhGXmeNzJm37tQI
8FrwKSG0zZBpXeHIzsseKd4Oe+U96XlXF+jXuEf/S8hc2kAeU7YCi8G5rep1+hqA
giTR9wWnsVvNxZpQm1wWORRIeAKn+4ExYXQKBorSjLMuCwvGsD6JYI7ZleDU3c46
ZXPuYmzD6Hs+Ct2zSItQJf9A6TGhQ3BWXgMC8BiiXDYE0WqigWAdP8fdTxSNMq3C
j8Pltbe8Csv/XmOlahfaUG1pdUYJnojHtKyJI6I4z7ItMV/kZxCZeXi7fZszcSk7
0MLYM8DBxpi+a9elwbC5guMgGdVyytM8gsV6pSCoBDzhIY+GWkLhb0JUBYkruNcx
TP3g8r6P5kj99l3ed3CsdLk9MpfZAgtLUxRGS1FOIzRKjOiWke+4tdTZUvBQjOeD
jPNFcikcxQ6WzoVPLB2MB6OFI+RgxXt50Lt0jg4X2RWXkf3COUUWcDHQWIQRl+iD
OJ9VjdPj1COWADGrjxjBTDB2h83ZW5sAdXiuDF47ILkz8xiMqvDmf0clzHMhMzqr
qPuYYsCPfjWI+JCD7tVWc5gmC+nCJrfwNKt+eaHliDPajanDfSQ8wSw1nkBExVxh
qoz6pP7XqVQHohktZq3VWMj45wn0Ad4fzasf4Op71stugXWw4jSvC5TrZMVEBDei
f39UOsv7n/429d8BX/cT3zH4BPrSBzR6OSHSZu/K7QLBGfkcjWOJwH+JGFpEwFwZ
H0+TZMtEc+jMbja8zCTTBvLLqKx9Vr+BUiQnz9M5pmCfiyyp7PCv6kOQGRCu6+Vc
VKS84vwiaJf0fY8lunJIdy1x+pJFdCWh6y/0vHhg10TCPYyBbf4/5y8mgnI1EhGI
YtEmZpjsQNkH77LiQLNTTe2tCc5Qq7FG/3kCs36oDHB77AxfrpYlnHV6/9xY95db
sDl9pWxrXnLjDQjaqkzBzTTM/8Yeg3b/Zh1E02x3c/4YP+EuW7QiOfl2ecS9TEjF
/nJWAolY2/TX8Qo1M8fjtNnIuD7kFndITkXaZBzNfeiq8OWakZ+R5NFBooEP6hIh
SrATLtJVBVuZtNDqRkqzwuunR1TdRvxw4iMzuqyDT7bbHx/8qOenCTZFJsijONHT
FLJnQnAtn1iBnX3VbCGULvKoQ14lNLvKbKha/rk4cRLXbREHy51eM/I9mcW1cko5
XP49VvfkU5+dkj5y0Y1t7zWMomp5EqAsCzpiD+avdglGEqXElRMqgZWmo+USGgCq
1tBzEJwgo1P5IAoVneYUqZbc0mnvjoaTmltUxKYQdL3tYvxXcMaCI2OPB0a8MjWj
akM5XPF6N5eYe7CSVZNHl8bjJmbsv6JNHnQtSAtdmOCWxPZUvv6jMqyZuNNt5KDX
0TXeM4IrSlVjeihOuohlU0xN0GY1QRANH+K+NbdZBQ66ioM7UmXs2R61eE9tJ7U5
SFBHblzEgkiX6ubYDpAoEDTe41MQJb4YRndTnFDhhD2arXKjADQ22bmnt+Sc7pKK
n6TGif0XW63ki+DxvcmDfamqI0n2/zY67gq+FOA9LqFhgCR7K+WRGJfxjuXdG+RA
50F3n1KZnkTcyEuxN/vyAvtiFvoetRUQomLZipPRt2Q4enRZwbQcG8XzmLV8TkGO
nIlwuyCRo4yT2fkM/haTk/SknbYgqmeG6GM1f3e+xQxbkskUVmOwnifHThIyD09Q
WNfEj0XcJ8yQD5Sb78gbxL3kcsU2HjL3jbfRKKpvRemeXhBJ5SoheDGwTZN/hULU
peENCX3iy8LQR3+dc4Q9hVZtOVJinlxBPO8uXoo0Hbb9LkbTvKvvRswAk2iHFo1A
mJAlvnQiVpMymaArwyoZvK+TvcYYohgu1KldCGnRBC+2Xpbz7FrifnSWg/O0zRx+
eiE2tM4DIqa1alkykW5/hjtJpmEkpyT8nn60JGaDgds9Yj5V+JOY4MmmWs3CoCVh
d51tn4WbS34wqfeskKuwU/qPEjv/rE/4iDsNmP9d11IRbS5NXw4fA/EexapISsax
LrIo/4AEH5XbiQc9pgfblGMVgKeklQ1tGBNDw1pFfPbCZeN1b+ZGiPcZ4AtTQ2MN
k1GNkRngD2aaYvLLJxV2pDD1RBpjHwDr+COeojxnbMyCxjPOOxe4Rzu04DRo2S8b
d6BsSvR55FrfJoA/y1XeEq18WlW2SKwci6KxKRfgdPECLH2JrtApj7lsAPWws62D
70KywbAzcu9xqyfgXBj6U6DCKSGUCV2hNWSArCjib0Rsc9cWb0a2bsQ+qSsW6kIk
1Q8r5cAbZ7lCW4D/mgeusW17OkQHgWQdJ6WWdCrrBC6ZzNZ9xJbKUWVghZkFym+o
eNusi1b19fDTBufPljUFFkZjBAKW4XhFkBadaJ8BQ5qIKfEu5U87sIB3v2ok9UsZ
EWNugibyIeglDK/KT5mwS09nKHEff0QiYf7mARAalnjhgiZFW/CCOJYzjCcecitT
h3Trw9V6CNddMmOhpEjZ/6yhfElu6Lc90RM5gYzMBkteiR7l77caF8/MAgILre7C
T9Mk/NFN5cKjbGuDb6IfvQcBfaZi+0sCicHsznqnu+t+yATBQJj1TpIH0/tyRMrr
aVrCHfPghUPVx3mUlib42jFm80V8KlZTLuLllazWZ1PkeFkztcRJmUoqFL1T7/ss
GxyAcoUW8AmVeQ5N0/wCO2SqLW4yCGQGVrH7DbfhCTfUFOPuEtCNfVYcQCu2EgdS
RMlK82UNdpXydTQEcJPZit+ITqe8SgVJLw43SM8lPFxmAvLh2vKMfc7nnZ7Ihcbd
2xWTJRgNl74amPDNgske1kHZIPtfIuEBz6DRg72+3uaEDd26qkFHPju2OXyqHWDR
dumMTMbuZbMWEW0C/WSx0fBCu4CZ9lwEAAWXmNBB1SnRCGwuz2sc3BhK7MQ9iOde
tx9v21NXYSd7AVXlAlzmXme3uVPRh0dyculfc6D4MHaVrz6/DM6Kd257EnHBBDBY
jjZTE1KWkJsCLa03PwClxAqFLKY0fVfzVU50eKyV2bCcFT7GkvHOGdfu4XkL4/eE
7BUjkoJS/CzE19q7WUoCmddd3w1TwXzdoht6/WavzwIOyyEDj4cD66I33kYFvZ9d
x52LLdOozsEU1JBZTHTKNQ9TilOvtEAOCMPq8GpfXub2coP2OKhq8pFDJbqEebn/
8UXvko0QrhsByxXb3goI7P80T/x4Uuww+NC18MmlAFOYKP0phScSvYiO1dV1b7w2
wKZ4KLZkojk1jEusovTGFAT3IDcanS/bnPFr9HWg9cMSsEO1JlhGQYjOzjH/BUcN
jJZY3ZznqLLnxrB9UQGMRvCT+iyo3BHNGPKZaAPWX77m/7kCv6SPDaiYS0fwIwQp
Ds1qM3L1qgWsAw0w9Bz3rpTLMWhLZNAm8m4DI7cQRhdHKyUuplzkpZjJVQFxK8ES
NLAFtb+7lTfRrMKnWlx14pqmtNsMIt7sKvwRYFpiqWXZor4zEg1N2cRMjr9r0F2c
gMZYA9ezB3/0asNEk3zXeRQAZR5yUYMWzdjO+HAZxL/ntRxC/JrKp7kv7t6ysqPm
BKTdkNmO/1YnutswxJTqUvtg9OWpVHE4W8cfmPGRldlI3T4k+mF4KOj0TPi6leiU
FhKrqqlrJeDY+nQZoe6utXYWRsg5Xa6B55oGLE5O4JE76jDPHhfhLW0ekLFtebB+
3LuYu9d+NdlBbA/KkYosJ6+uAOGwRYImQrhpqUFHAOJD2b9+/jmieOFM6suh0gz0
gZrNRTB0v/znpVpamBeuKSij0YR/GuGZcxOkuIk7E8fqrS2pdjFVg6zMqFUEvowu
78mqjx+4RmBuehA8qNrnFI79B6yNckW6k3CDuCfy12ALtYjRKfTafteU1SnEdG2p
5+F8kSoa3jldTDQcn1r+/cEUEGBie63bbLxb/XkfKUOu8HIBo26rafjxhm7CcSs0
KiW3p3RyP9diMJMDk0M1KTodSmC76UPa3YOK7JQrHxxeCFqQESqVlB/HekyPy8nl
zFp90ea8FQVUBzV3Vov7bBE8sY/L1yOGfDxOoyFHV7ERnc/JiWKPDppWZXIhQAhM
0zU2NZem0bcanesJ0SeiheulnVoBys3ojsrZut4IyXsEB5fU8yBLV7naf42ij4xZ
Yew6OejuxSRckP6MNhcufsE9mIK1zw1G8+HQL2Bomh6Gz0R2TTFm82eGelTOVyJR
ZzPTL0c9/qp087CoK4aj9/Wr5pFHKDoNRa43KEL3RZKQogsf95EPb4ftHmfZxNuk
WGA+A/SsS2WHDTKr/03YrV2dYEt6YxtGmsVp/WS5j8cr+5hTOjkcm0ravXa/b1th
8DLp7EE/bV277z8aeZSM2TOL+5QbSiywF6VbPwZpFyMsiuDWBjD6oYRsXwVpabQW
uFhAPEzEL81w2TZFvFPc1+gBy15d96ilIjiu3LzUSEouE8F72dGqvWyFzeJDJAow
1XYI7Db7QlIs7j2cpRqUttOI2zipzl+HRXSaxsQFoVDIwohDOCrxfcb3F5JdxSbX
o0w5Tm38Nk16BWqVS3p5Fvfst48WLD4uyOXif1AoUuLyZytI9VII8u35ZEJNpJzq
b4YkKZbfOKgFxgliinuN3KfZi8xZEXZsbkR18VnLVqGZ2XLgU8+u6WzS2m7tK64i
ZViBT3JOEgNlqslm/5IBfy4zfktfXDwYvBEwnLX3kZ7CgYxrBTu8cBsTLzeqGvn0
AZVnu3MPJXVQwyeJjNhXs/dYewMurv6rWpNzi3Lo7cSaHBp9hL45WgeJAwGi3maW
RmbpP/FDwcuW4s5LvgLoVZzJjlWcNKGAiK0RFFv2HAQO53Wo967Lj86PWbsloUQs
Ey3wB4Bsaqb3Oh9dR9B38bR3VcXzPxvyskB76et0ZHtZ/e4le63iQbSh5L7GDJit
ndPaQRzKvBZiujQ8Oe5GeRcIH2SL43dWGlTDOgLYfgBHV3U04UJprAAbrmJeZWZ6
TYO2qlwN0jSww4ZEYfmyaTZSck6zIv6yxB/DF6VVxpivCeOKKMz1hFEHlLLWaF5R
CpzQ/ROAsnPIMhr0AXzHv2/1Tee9y2jFqGUgPiaoFILvsVAJxjXBH0qoSuwH1854
9+Tg9Ols4foK1DoIipmGdejvKKvw1CT2DsDSGnbSDG58CbQcg7CsfvBO13xuUelL
zLl4UV8nzQuG9H9MB4J9g5jCmHffmWl9M0d5qZU3ZjZNGGUqbJ39Mv5wmoE9Wfgv
cKgXtikqsffUVakXaYwC6nXaeVkzF4QG8hKZGlOrnzUI5/OcE2opHYLs98Pj26Ik
EovPw39fsNBCviPRrW06NJkHd0pvQeu9Le2+PigZhjD0mepj2X6rgLfuADg2aKxS
k8SoeT0U3Vfmp381YJfH5fnjMFWcitACTEPSDGzFPJ8ZPt0ar+oH//1Wwf01J4+V
fVPYPH+ngq/U4Duc6kCLNoL34cd6u2ZFYfrKJPMLyYsGKgK8uXDpbF/7gJqx1Cof
1o2MRN1JCb701ZqYqcr5LiOcS/tc/7wIKwV0uvO/nJXe7iz1wba/uE/tdtlkHkmO
A5TsD0R0UQeA4UrEFGA16WCC0cGBPn5b4HZw/VtMy47BWc6UvAD8gPhwe4Xi0+5r
qebol7/f68NlAbcVNwqQiASx7n6xa6LU0UxgG0Z9Cs02nn8YL8fRbCEelRPTUA8L
BK0FXDjyxHQiLH0aZxw4XjZOolYcK7hQ2HrA3lvy5XYiMSEhzzaW3pudppblVjGt
7/zAao8T8ZsjTlE87IJKJLFDXrxPnSDaysoS82nC+WFSAO171Kc/VKeOGDaQTzJ3
mqGQ9hYXHk9GjUP0OlwFpAkdjHSL8u83luLdsb+MRPMy5ruGEOUaARpLsTYNfHnB
EiwWgJ015kDR42+A+uTJWrb4sTmViygsMoH75FPnXdQVFfKsCc4yMuqkyP6toUzM
7ye1bWfC580EzhGC5Y0eqPaHXPWV0NIyVc1utFUW2/piAJ8wPDKUUvzjYwpH3FtX
RW7J5aYqux3aIoxECyTp6KdU+Z/jGlxFGwwkPgyh/YTaz3u4O3Gkjr2BNqijxbfs
vrY7u1cHFHMINGbSBqcbA9nb7CRP/ZWwkXkAWQqJlMvJLOzqgw5CoMBpexs8X91C
Ti6C0jjMtNbvfTwfl53/BfKNCkepxiOUBDzvBY8hjFrvD1od58JPZUfm9oj2t+Eu
5oZVgNQ4VW7FmRZpwglJ3ZFs7gwO3DUCm5D8CFBUdUf9Y6/aFVhk47IlIbZEzJ8x
QSRdwT0vDMELFUGRkavSkTBQge+2JU4I35s49BL53bETuMoYPvcRAiuruz3M+TEg
r2d5Cpjf1eqH8sgRonIzsYA7tx4AToC01ZiPlkfRb2j0gemKxh52S8uSulldwUuq
cc6yR+7V/yRueXTuUeax2i/X+ZdCAYn4grcmwXBxSIioPWaeX4K2JsPi4FoNRiLV
+6gJgTARNDArAutSDDUwYDTY3Yw8P2lFyv9JNkL3WmTTc2LbsPLR2wV4AyQOXVXJ
+x3lBRsnBiXLv/oozdrhb9RbsfZoJ9QtfyG1Hsh3HbEnkC9Y8oGHSn1Ere18LHFb
dGmEZoyzWS7Afv7ZJJYpL/1etDAe6rWsNnr6PG33MSEdIxHVVx26n8NOyAE+uMMj
bezBRG7X1L7i1kGcML8vy6/BfmtXApoKVNCnqPvG+bHkBwtObf+SpMpp49asiaf3
XpljPElst+RG74ssBriAemE4XGUdq/ft3YAd0UbyUvJ8ITD7SVdIeTW+op+3qOyP
9prOKOobgQxN3UJS3D/eLmpBf4I0oaVFns8eP2MTiwXQoan/kLkF3OfD4lTwuhGC
DHEWlrp/wN7RHaHpKkcJVNDY7Vr8udkYnKEI+Pcyu2dkCoPkuQx75zhyH61EIiS+
/J8rk3Ddcmd+E2fOOQX8TRKbxlRvVl60LMTv2YbfxJ27DiNxblaH40mXjTuX2WBz
E2LHV5pn1K9BbfJDQy7pkIIrGM8kC9Fj3l5KgBKo2v6V4XpzcQ0bz0J4GFXRytzE
1Vz3u+nMECSKTcqrGyyvRfppL+lqpuxh5009FQCq66qHquTwr3jpZpj1j0OATcfO
aEPSDBEzilCTbSZCnqLFgP3W3lBcjAQIDwCxVM6S5+7bJjLwXQbIWRmMTtgudhno
dRr+/408UN9XGgiP20MNq3dmAalSVKUywXYv4db1gIf3soTfiP0HNB5MN+N0l7Di
RHrElcFe2GNLviRbw/nqLyQc84dyHWYbiTUzf02mkrXxH3UkTLNvSHCjlPn6BLeP
VqhkNI42cmF9hvirsi/kBmUFXWmPP03f6jarVmbBf9nimV1nsIkQroP2mK3kXFGb
hbNAqb1dWip54CNda2dcNe3l+y6V99zOn7dJEkp+SLx7h6GGd4CvUFf/WlSRTW9T
Rc0PRD4n0h86DV/J1xMx00yFlbpshgEEP9XOEJ5oy3qcZ/wrfisNWvVFz6Qbzj1I
8Wge2/ARvCvNF8BoO/gm5z1FEJx0a4qa7kOMkIgcV9Qfd1kKe+p1ZV3KNQtxQD+F
7MunSbFUPO5goMvPQwrzupgXXLJ219Hov2arc3X7o91URTmFOHzX4cwI3/I71mI7
FnDvzf/Rx0eniHxV2G6sfLZ5k9Sd8KAg0hs/zppI/O3kGAlrKqy/drLKs2qgpTMW
QZqB8XYdIGb3Bg1ENWUlSfRHYRltCSBQTXwyrmJjh67Cm/gYLKGfw9RkqZQmhUqI
7v15EA4vERliee4CrhwQOs147NMlSPBnqn8uJS37iMvoPE0ltK+//bziA0fiK4y7
mHHh3pEjqraV3w4xsRpt9sBGrZaLgMd8MLq5nT8BkKug97TpowxmHnblR/rlgOto
iz9BUc3pHJjAIFvzUiObUSInKz/sditWRRdtUNWNNjZMQk+Wjhg/ze/QT8vAk8ie
qKHiMLrsr6HLr+7wWXehw4Yb5nm5m6ytBTAB05zVgy9FyDyGmqmS9S0hs0UCasL5
FFe4MDyJ2KePM4XK7V9HgpTwX6vvylfohBI5URYxRzohLPQZ4e6gsQVQz9QQfdrU
77ZfHaXwbFWOvnbZvz9J9wWgoXnEr27PG3gHdVA0ShNdw7Yah4ICGsq/AqxGidWl
9AK9qoagU81j13+wFaGYov7KdGQmosN6QVnOox+KXCqHOL5I2vHBwrHSjfF8K0fJ
HLH0069MFSDcQxXMsmRhyKTtrQkDNBcJhcjZWsima8mKon7NkjiPuLwfCvdSRt70
DW0LqhPkPenWzQLpDN/hesoEcILrPuXdkQKOK+jUlgOHP8qf/pWIc2tmnLnA+kUU
Rb/THXYvHxKXxOR55F+2u9V16wu1y74aXw9yjSI/skLF53Kywit0r8SNUx8PKthb
YlaFwP1N1y+2YeXTqnhoiu5SSDdqRQKuZf/xdzSTk3qWxNHr1lrpyI88MrHHRJBB
HVTYtCniKKck7AFaoF9udYEtLd/59BV4SXi04RXrCTi6Qu88Nv9PafzfYvhKG00C
KYiVv0HS8aftN3gDy5oJUS0QAVGMgdDZPTF9Bw7skZaMZDwUrKHjf6tro9sHRl+l
SCVpUa5EBrFwH8JG09X4LEgqtbIYh6yAj38lsOQpl7gyQdLYc42k7eWr12+ocGyf
QdPQhSpRfROVtt/SN0u4BIOV2gSxaeCsUhV1ppLL68hjX2KDRzP9yod8Br1KArUZ
ZC4JlTiixbWaoPw2mQOBgrHOL2y0UzKF1lC9VS25xH4i8rC8DKn/PkSw4oyjP1JW
fRMx96BS7gYUx2d+OfaG1l8TukQSxEuC5wgLwxVkYbcdovXKXRLLLRkFDDTzKK4s
YLe12P8AVZXq4UiV60bWvrl3WUgG6MwpuIO4eQtexlUIXVlu2r4fkh7XlWUZNJNO
GSNUDo8bic/M3ENXO6cUBPlBK2tKGvmnmvKPuqqiqIkZY0W9aoNmbFcd94g3yTfv
QrVSJ+JkvkRhXme++a6HZ4m+3tSSATOmXehZ21hCcTK5PmXd3uNByXCpuM5bk+bl
MnjbasWUFrgKHZMf3iL8yhN/n/+lAXC6XcN0e9IiYI9mh1qzCgs/argAlDQD6rXn
4nVVVGIZ+h1sAae6oB4SaamfU2sGB/iJDup9r8oAz01o4bUUJtW1BRZqs7VpkDF1
rRazRlxZNAdpUjqt5DlIwmomJmm6nyvCiiCNGU8+0HYKRIDNtlAXhI5X7BkfCh1B
CdH+puU2u6/p+berGuk93v1GWEXp+Vbp+Xi5OdY4aBsXE/UfSwxzKoA+O1/CcFSu
G7MlFC3oJv5sPIAKdKtHg63pg8Dbshg/Xo2h9T0NgaSsHQb0W5jTYAGSbkb/tXVn
IohdLw7GAk82C7X2p5CmArwr0UEPFpm6wPopw5JiQOmo9c6AgZIsC2v1wBLMYoCE
fOTj8/1QdSCkTAEh5Yf/G2wua14+87RU04Lxrq30IWJKOCfRP7+sB+PxZIIYBZjv
PcEE7p1O3WhP2n+yo2RoJIaJZj4ld0qC1opO2nahxEo9wIOFdLUsQkUrQ24NVUac
QOkOEExA5wwJnyLm59O5SaTRonQOUOeAKTX7Vydwu3V9Syu+lssjTM2HCeaod5L0
RAK1hOyCqvfGarB3z8Ktwpe8jE/Ubvah1Cqen0Qg8YXeh3PwoTixZleQ3OKozZvD
TJSBqRAQpngXHBxZGQ/zWmI+7+kpmnmm2iT3cL6Bb+Y43EQY1XfWdB+XgeZlCslt
2kirXG/E2loJ8nXyOmTC+pNrr/57a63LerQdTh0lKY0J92K+0gW/lHeDcwdmW9Ji
zEquwrAJCFd0Jgk/waEOuQ5MiAeiZNE7Hy07pQ9Nf+M4Lgipe11zVdxRz8CoZ/1v
JSqnR5N3JMlOmoV2Dk6k8FcrYlgvfc3noTv5fqJzNrM+ZOjd7JN1kB7toXzT41wI
chiAgO/QeE1OR0UW2YNt1YqHDNMG+K5vzDZ10rxaYFh9Q92OkFkSyurNnzeSE4Ru
rhQAWA/QgSstCowrEmtCAqHAW9o6dZeHkuH6IYjuHzq8SaR6kJEhZv0B597VrTxL
0OXIbk0LVuC4E3DUH89jUA6Bwy/krUMCv9u+pgYJSaJdjk7wvrm9dj2GA4v0ALrA
01OggaM4PBFt/gJWxMtH600EktdBJARRscKS+ICeZBy/bUvApuMOOakCKr/Onh28
asRRFFKs1d/Wfh8GjSuucxDgBW7So4DVB9izEfT2R3gbb8f6wlvbY6RXNTNuOMuT
HiKXCm3mitk7RuUHMrCEkSsIsB2IjFlOkSiL66dV1dxXkwWKoeAMMH1YxAZuqMGA
TRsfE4Cu9GjqaD42OXlf/pXQLv0kOPZ8eXNSztri4dVBkM4Rb1JWME47GyK4vKC+
EQHvO6bFYjq7ItsFmUCnH74jj6r4+nemlTHRgJEuLKYZsbu/PsWErGlBrske0Za9
8m3pK067WSr/kFnZiExjsquAT6fsZKt32oyD6X9aQHi40EvLF9CHVlkgiAcrIHdt
xVujqMuXGX4OpcYF7MZxat4AB1TIngO95mDT6lHCjufpYs3NJSsPBGnKoc6aoSSb
+M+UUg6ui9Z07A+29PtNZT9WCMghJEFV9UnfTcLzBJBlrszADx6/sIW70R7wP80S
2HqKpISPBlVU0kTmnv3YtgF1P3+DJRQI/VDvwgKaYq/RBPq9lBFpv9g1QlghSKrR
7dPIgw1ABT6H0mYLDQdOEUzAYL/RRzHNLlxE0h8wF9fohsskHkElAqAMXz4QMgOq
08R9TjGTwVF/F8Tlk/7sQ8ZwT/3xwqXgWcIge3BNAPCoc7mq57Z2WSuX+0hp3l8W
J/ZTbrxN+5m9CNEXl72swIk+2XsV55naSqv3pWI7clZRZMTJvR640yhyOKYuZMGT
fdo0Czd9kppWTMrtYbxiqJH5SchStIXnJ0fLJpfxGJcRlQFjAUHjYCtoGVg8jdcF
2c30gF4VCcfpLOSAtNNouaq3NSBVnr2dzrVu5rfawyM+cw4hsSvVJ5GxKCL9sI9r
BcteXeeaGbUyKdtdxTdmBD3MtS83UbZOYHeX7YfLaYDZoIpYPU9+OerUCdXyN6Rh
BQearKYVG8W5Oq8bK5qNpskjzBsMnnoFe98VM3f/hAGv7HIGwD5V4rZDuO+SNVkS
cUsBo8JdchZku3wla/Jw2DhXYHn7/pIRNuceF2RJbfNWdKmJFrM50WeRhP9SYT5L
4x14dUXkBofVBiO1LwJ0EedLLSXOC2+ZTtAKkwPqJ2TNVDNcJmb+p9qh1C+gpdLA
O37pfNPRUOf2paRHBYnGj4EXK72PkC6UScKKaRcg4SykAsdZeOgzWb02b2afH6vf
TSuEm9ekJ8uPvHY/0n05qVkzp9ypInu1gBWl11Lb6mr+11n8hQjWDDNQMFlBq+Et
dVSpMk4UP2MjK/G2pERxuPasIp3yY0BZuhLJ51K67ycvEx5+K7ZNYMG7VGRQKliO
kEZOwQVW/os8W0R3nyDJHJbaZRE3goMIBKuLstnH2My8IwbLrb8fap7KGyXdL+U0
4bUDEHMk1NXJt2P3j/vF05gf4ILDqHOxxJ2h8xvm7tK7SZiFios9d789jx6gAp2y
/1ESsV2vQN3LP37DloMJ5IX5pQGqVEZMOz35PlBBKoWZarq0SgMj3CoKZM/g2LEO
EABWIVhWM55pGzx/IU73k5iHDUdbNClqaNcOH5f3JfIhjrD0tfdS/q4fQpC5SLzM
ahDpPlxTGJYvAnGhhLm46RKuvjutd5H1D8J1zUW/kLOwgDN8twp7DYGg0fm1Y5Pe
L85nQV9G2bLo5CX/Ywx8VTsPi1vIrC60B573Clbe2cZ8VfDuvxvkkYfqsRv8xlro
TbEZSe1eBJHudRcVhqobw1e/BDySlTBIUfdRmKsUfayJNRsIEUiHhCe0StXBtz2D
ZgNnNoLDG5mNjxLqmlKjIZB0KMNAWCIg5DzNVCHMK4qLjGFS8W3BzmvyJ+ydAfA5
jsrJ595nGioMx4mNLM1Uv9HyBo3nhlqSa3Ri1cSdaVma2Q8azfpMKTrEoO/t9TbO
lNGZRRAUWLI5MaFO7QxQcrAwuY/014iATIDZEMbt5qadfwP8QTZb+Hq3RDdENf7V
FRAAXU7Mnvub/5CeGc2ZqVbI9Rak0GT5L3NnOKauBADoA39GjQoWPgMUHyOp7fwt
ydPQyxokxgw0KwCxuLhclg8v8g9obAGrcxvzBY8dpelK3+7dAL15k77OcPvQoC7o
pOHRhkGeUh+j5AwNTbbhtBHZTAGfr9RHJ0b18PZN0cOVWNQf0StmziQI0wrpF2jW
+dOJ2FEOeSwu85/O1jhWSBTwbiNAfWndzMRsm3gWdtGBcCkbYs3fE0IWfBkMoLjg
VRMVpcMR7JriaBqqFl9YOV9KyPZBqSA6YXtkGvWHmOsWN3rc/RImfOA3fdeAf1Kv
R2SCq1Ugr2OWjkNxUrHZBqOp9U/bI4sEc34cXE9VJ8+W9pVEoMd0MHKYpcafQ9eQ
iZ7LGkUnnQG/kt4pRzQI3EX3j0sl8DznxgzFs8czRbvMiWq8OA7Q6Mfq8iXofXt/
W/FvicAKT6RVfpSPJO487C4GZd2aBAuB4ltgN8af87mlhvPEOnumXji3mY42nlg8
UhFiasr28f00J6aqm/uPhKMDbmRwwW3XNcKzKq7J8j46gAcF8YwkhXf7P/me7IGm
oeosGskv7lFy/zHe13b1fFYZG5EdU2xgg7b5dOlupWLC3/Nt0055SsQVmBdXrxIf
qa4I8d9VPvVcpwyyOILAu0JgNth++C7Yjp2pjH2H8+mOQ4lmDFSIH/ZkiTDSHNJp
1w1GF5JEr6+3E5z832ZMltHmvevBS1j9AbmvVE5moE1yWbztDVc4rDtMpPFz/ns+
ab/b4Bw+AbesJ8cigp5XxoK9SK1aZPhaD+jZ2CwwaQXUun4nrTq++0VfyNFouoj2
i7ebTUu0WH/vfCRfu5bb7tplXENTRca8TTFXR9HY6HZ5aarb5Xo+9QVtix091qJg
g6pWJ9dGuR6PkrxtT2x9/67peHDoD4GfbWH1cNhrpPNUlrxqXYF6ozQwjUx/eVaZ
rioYOJechG1/Bnpk9pNIHFTRLGsFPXnibWamBOrmK016VfANu1eRg/+8aS3ymiKf
vjNgTd1q+QbReS8+3KRPCCIUkw0+SUZzDdn+IRF1X1U5plHAHAiHkQSIqUrnA2pb
9UYwrgHoYj+ul329n66ZMjzWi5pjjjLiJnSWcS8QKTov55J5VIjDu9cKDc4PmpQ6
hOTSf5Ej7SnpzYCB4W8gmjMY6xRMp1e+J+Mt/MGvOvogyqYEwF0YQ12bNTKXfTUE
NnbjIz493whdPLLv1+jLp3UqEuWBbqpZ/sCearHaQx9dpHsmfvMRgymF6tt3jBsr
MoV/f27VunkTW7831TbFE8MShBlxfFUXITUY7hiGJtmOOWkWPSbAVDV3a8cH+YG9
yJbfJ5Lp+z7/Dl66VGgp891Cktx8JEkjQVqtxX4dacKF+vFpmfePMaiCpoIsr8gn
Iggc0j6jttH/uUbsaOobaqGqwlkJaqjAomOwXqf2ba/3y4Cg9lILzm3P0nQ3WjRm
ak5eip96BniJd3VJuu1X6iD4k59ZrRcqn0Ygrbr3hWaWN1swxrWR9a8/YdxCpUc9
MQLfzhTFQ8U9eOKEUYBRTQFPZNkwanLtNyl90M/jdri1MnOM4SGQXkpki9s3K2oc
4TbS2Z+4QKxE37Vjnhz8Ot8ZvdGnmmsu00tueyRifGbhtZ6ha4DSE6E4oN5LBcR7
F2+3AVJLBpZFIj6WNno6O+d4qN9rfF29gtjv1jz3oxlhR3D/47eLbBs3Jrq0+2VF
NlGLgHDcn46GQGOcs/mVaKBURS5MRRg/kpAB8fCDlEYBxo8lNFd3T8c+wyyjCmPi
1ZlQUZ+BAiAEIlFRL7sAgZKj+jBq3UmpnpQmmEzrOQEfKWag3ORVCkUGMskYXinT
bBXjuRaaB60a9maUbxTFUxKQ16D3xFS8NyYbN8j99bxnHUQxSKIlTV/LRVw98p6z
uPvWI5p9oRVwwNusZEhHp1JrYQhSeB6sBgzlYIVdQtbflEoIQTixXOqkVgE3yP9m
8Az1KxpaTBqqNxaVN0HIrKS7+ksxFGE6SZRhweYIfo2X1OkijBB7YljtG98ll5nb
kVCuh3ud5E1ggqmpeUC73cZB1k/gFznODBa5UX3TOlOD776naEsbo3PfqUedFheR
tAqJSogSazABjn72OIwKzaMbZ+c+XwGyrkg0A3i6fyPB6CVhubVr2ASSFwukd5tB
5cuhu9R/htyMW7bhlG/izrbkhwFH97W2iJe8JehyKHr4cLWp9WK/zmGMp264ffNH
BL4vx1BvT9US/Dv1RKV8136+bsBFbiFIlLBP44H1yVO9U4gabA31Z4OTjSN1d4iA
6368Spe4o47ZitUEX3knSN/KkCU+CSZPLRhpjx12/oC6IZ0TpjUw+xZcPDwdJBmr
gxci8HKQtaoULf+cqz5PfdvUkkqUtgyrMaAZyYcUHY40dt0KtjDJzGVlfhO8TQw1
Nq0ysbqqCselIjzwpvBna18aYwEtut3eTd6Mci7tOg1nzcFzUZ8Fweuf+BJQL3pZ
MuDRi6YUWjNQd4zVQcqnCZjN9Qz48Wt13y/jfGocquNTeMbJHIxI26b9K05nsz9j
GehmSpkq0Lcz5Mw4jgSEPKyng7wqJmeh5W3yOcSy/cAPl76Z/xOT8QzXgBbU8kKg
nGEklUoHD+FXI2xradJSpyRckmruePr1pt2PwGp0a4+JhNVjkNB3jlxNQMYLm2KN
We8WGaEpxFTB9oCfHEPfO9Gm3DqBtkVgeuJebbJcw0FK/9rODtMGUKsA4PXLbl0O
C+CWpMJZFHwxw9YMUQ3V4bcCo6foNAm8b39CU2CZ7RGctEhsTKuMcfM0saIz+K/T
9qOrRga9+JnJDgx5gvgic7OsbND5Im0w/yzigNF3GJ5337koXij3BeKDOYP99nd1
1mzfl0SmDAr1ETjVosfYLAVOZ3MFtKhHezaQevucALREkJBnUI5kmwaHL6FEjLLM
Mlkwq0pYgYBS0fKDfPS2SRAw4PXBOugsT99nowqLHgVCBFTXgFzbiiY0fP4S1Ena
9PJM3HLY8P8L+PxXB61ATzUZj2QQnNnyidRvi3IGLLnXc1CHmlFs/I/mvvCMgQsV
GqDCOXGEpPec6RdJsv5eazkgxMTEEZIUcB7w9EmG/oEX72O8mdDoJzCrlLDVCpMU
u+5K6DyGy1RIT0vgZsmipnUOA89ZPC1r3ok79atzPhgTmDym/Li+UeWNiP7VEN9c
9LJxmibwXx/zX7kD3yb3LApLZgzneGfxGRM5bo/jJC/NiBBWMPeKklwn+jV/PioN
t1ItPmcKUsupdSdnx5k7phDLKb0GvrA72/Zhz2v3m3JNise7LPgR1m2M+rD+w3QJ
JjYcGnuOXQ9RPeKUsVtHx15qhXbSDss+Sf3p2i8OHFsly82s7HQRrbehNXXVbhSY
2FsshMppl8vvmvNQnF9yR7DAgGOX5kSV5gD+2GhqB++84X+4w0ydQK8s7DxD/cCi
zdYaawsh3XHc7AhkEdU+YDsjZI3d6j/1VzgD2lm7QV6WwrGgkBAT5jQZ/KAT/kdx
6bsQy6JKWl3iRIwhxDGEdWyNcuGrnP+3UL+jeWVLkQ2tNL+iRm4GKK0DTSK8m5Io
Q9Uz75SlcbZzgag3Jyb1C81ZXEDRYtTPJ7SOd3a8TPMjvS34MXcEg5MVu7Lu7+sg
L7r4fRROGeBTJ+g085NLURfL70XX0guhCX6ZOPYmaZ9JbcUVN+njK3+AVykyFkGi
MZfJKxp4R+5p6S6yO7uBin05vcnO5v3zBR7NUFZ8ryc7QV+EmHFuIWC8i6LosBpg
aeH4tFUO7gS3fJzNsYDr0YwP3VDwFFVg4PdmV6zGXtXYd8dDcv7xDF8DLxrNd36S
eDREP+dn6nebbJXB5DJihuKYCHz6IiQ2YL+j9PweP7enEbxiwrfyw0k4JIjFkdib
2oDl4RtzFDZNW28+Nw883HRaJTUcpNmYDSms7D9ATJTA4qIvUhk8O+9wIWPNDNpj
4rjQwVr3vFVLYWRMUXB+3auQUpmlmeDcuNBJ3DxLi4JZihfRZZD+d4fMBklAM1j0
yI5ev4QD+NgB6vQ/CxumobL5ZQLyGAOC5fQSAFHvdYEHz2BhlQLGEvuyGKfBecoT
fpMCFh6HdgKxfc4WlfY8IGRnRUgvEynTXMI+SAGE6abVuYwE2HkNjNF+wzL0DtY/
Vx7l3dtI5Dl0ZxUlpu8m9ZeyVw/NBVKuz62BA3H0xKI18hVSu877Fss5DWsKKiaY
iYwFSM1UQWhe5p9oZtBPdosKy/hIcLkzBWCtjUR81rv0UsDv0ASvgTHxF35qH0A/
nxINRnZa+GBu+9yYitYqp6nSGUi/47byGjhb6VD1PlATH/OuX/QubiZ6/wv2FxN7
fUDJ+8l1nHcbpvCjBEN9lPQhh0/NU0WKFuKz9toU+1GMu790EOpifxxQr4d4hQCu
QA00wfIuzdrLAyWHHlLpCUKWNyXpkx0vfs2rKQnj+M/ztjKXnfEAmQhn5/oHA7V+
BsNRliZwQKs0pJItsYKTEykY7hWhQyovHM0qcLAzmyUoaTn7v8Gn0mxW5MRLsKeW
WkHys4eqEPHb96NCuJpZ8IXeSl3jv/T4RGxkftnZzbf2au89wFMaLf7aG73DQZz4
joACxMEP3Z9YYuMCxfiGSxkcbKCldw6i+tEKnE6R3zyyBiUr3+d1qXd2Ikp2hhmh
ZrvHyK/AVvWUl9SBIztu+eJ2d9YzKHHO/4R2F85O0mwvOJq7f+nQPh9N37GGkb6D
I56LqV0H6J8t8nYgg9D2ZBXp9fepGbYYvdDy3mnplRE5G4ZqvmLLyaahj9rpNOw3
dWDT+gOSw3jMFviq0EmKZri8uaE4MwB6WqWJG1UJfmS8WwZ/JImWQo9QxXpNubT4
T0cfBUJjFe0NXGXp4ypzMmBIrRKXU84A7BNRJi8jDriJPE2JD1ePe0ZQe7top0Tv
Co6Rf0EnB1gUx1gSWMT5xH84JMw++pvUEWuLeafgK5qRCi9+cTsoZKGXUHOrVsuW
GNCIVq3BNLSq4++Eelg0UmCufqbdVVxJ4jB0LkvvCVE+TikciPnur3ThjbsdZZ+I
YvzP2LBdsf4Z4yRgRq6RZ9C+hmBzOXfnx/l8c8q+n/IclAaHQoBX+Kyei/LWiUOK
8dETxV2k88q3lTViWPFGiBAVmSMFsBb0uVy0KIExGHvKbIgoyQ35L1n7UbNbhpFS
Z32HqFjBQxU5kECDOoGpYGb5cdYkGQH3TVSWDUGUiEx332rlGANMHhaPtkp2Srg4
WHyL6Wuc4LCTEqxXSgpWFdWTQgmqh+SP/ZTbIs+XDI5Bt1j6ZraVmG2/hTdxONsr
WEqoGJbQHhwWzPVKbqpFk+n6uYUgUgykR5UUZibGXhutjW1A+qhbPwMqbyodUnph
HRhYfnZ68rEkz0vTbJPwNmbVaNsB2x42OV4L3LqgDAQqYhX9sGRofSNR5mYfeux4
dPLdjxBjNQszvI89OFvzFORCJWiUnXbJF5t9NcLwVCqkJm1O6gPgUdMEmk3MLV/m
L3ZjAYBU2g091hQVeS12yjuIeXEvahuykpLL2TRaBYV6zRkeh0ymqfjaYvluw0Qm
dXN5UIn15hg4hd2NIB/jD2nKqR5d+qOQkTsWLRJ7DajpKKVugi0/MC4PcH5qSnBE
au/g1Wm/SDI5Xoy28YjZ8JY7B4N2oMsghEjto57UPJ99aPK95CeiJbe2nE98kFnd
TV6WdkFfw67n6DxhIsXlaE1/FdKsm5E1bWijdHsXI6ADIJ8fQLF/rtXDfKNg79pF
EaQCYF6/pV/6Ip3ZaiDNYgt0I7hLpGhWqDZoOOHvaOxDk8k+5xskkelpQbgX5bE2
ViFhe4dHYEaz1SSUmYwoxDI0skzAFuk4jVzRU6riiNrKqdSiphHwxImnW1fsQAi0
KOGiZasKQM+qEl+8VWCbpuyF7Xu04V9UAU4rurEfvp+clCJPT/yG5hAXNWXA3HO7
cWS5AJ8E3IV2XgHMlAQY0H/8f5GV5cHvxVO+S57lL4dqKtNxz4Kh/7CskLDLrY8O
P4lIp6RBp9JQ2r5xHC3MXhxnaR+5Z068YTAcNmRd7puMkt60p+5yNp3xodG44sl0
RoaVu2AR9lvaVGKORX8rHEOyv+6zoeskLZhLRWIutXrco13XrM1PxA/MFiGGurEw
dE1cKdVueWvVcYfxE0/LNQp7YrJ32DoqqC7ssUWlB6VluwAhnDwkpJKLe2/1FF4T
xHmfuEIxaL/4Go5i8ccZL4EKcahYFtxvWIhBiEpxOWZ58Ux40fXzhykyvD+oJe3C
ulcmzpvb8nbKVcB2ppsZTZh8eSY4LaB7G7V5sBVUv+84bvJZxjU++ne2q47tIzeV
P6aJXPkMWDOX3SL1fSG1u+CT3eQEK8IHoFdy6vp5HgE3DpWT3e47Djx7S1qtBfFh
PoQ+AyoPBT23bdmkH2Lyo+5bhoikujxP7WlzeSHw+ttrigWZ5Ls2E+EQ1cNAAAgW
JqJkeszopoX3SL+0qACGANUaIhVC4jc+i2X+lylRGU1h66CYOL6T1KvUtmQQzr/O
Ys8CO6SIEURABaa35wPJ7WciDGQEbvm+QxjUrjuOXr7YhB6jXQ4caYBgOIqAxf2l
vatymqvaBgWMsANyfABHmicfi5ccixJoHDcaDlhgVGZ3Kw8/kn/2si+upL92kVtR
G+hbCPxAoJ8rvw/15f6ofs38lzkywhZ5RmhgwjKTdiEYA8zChw3UVqBCzSDUXtsC
y1MA+OlLwBMXpfrUAGnATRmVoNbQiA2tVbuU+93S089Nw9ObnfT/6saCihivnBlG
W3a4NmPdG9JwTPspsfnLz9sOp4EPYQ0LEiY73VCB/kLhH04lEpfg8+yWIvspLvyc
fRiSaaa41ZrYzDLng2oDhDAo/TdB/y/RuSsmJggGhI2nYD6CfjMaTkN+Gkf74nJ+
l+x4ogHWrzo44wMTpHnVRfBV66o7qHOxJBdFfGiw5Kbu2yKLps3k5Pwq8CUl89Rt
BJtvFcOgPwNiOhg7a6YoZepa2HrJPmmh2HkWeXItMEKBPSJ2ZxsV52+CIE++kPqK
rsgEI4kzdu0AwYMd8q0wMmgnV7zcZGZbWF7vs5kvYR5w7wF6XYwVSq9vX8ggHa9t
ZC5nfG9Udhvo5gPgMpgHi9BdunJsgAvfTl8q256YSVZhOsa3X2Rg7ls6vHrngYs2
B0y6oxdhWJp9TX0IuHbZdoUhFilysfC06MzPFEi9vznNN6R8Ab4QSOl4HE2SXTsh
jBizYU+nIEqVkyCMh5uu8KIjvMAOY9qn4ofM88lTGkmThQu07Dfz1A1V+4v0txT5
t6OfO3D8oGNtN+tp2HWrdM2JdPtvx7bxCrnI28xdeBHfwoR0giwUJGe240JPXqBR
ihLzYshgzuCeeUj2WLyhw31ERm15hAXRfVGuutdgEBxgGb/EgJ1sRKKZcoQbN9mK
SkwaFREq+bE1oZIh3uh4OBUJFwEppfaOgjfwet+FZJgV/Ydn+iEjHG/SYrxORm7b
6UMt/tJjgcX+NKDEgahRyRCgOu3uM3qguglv4hhXGxs29s5r2r0p+/gSpw3SrUl8
uh7I71yHqpsjLgw9/Zs85VBkNRHCBeQ8eFkTQzAMp0wJoGYqsRZIduJ5nYivuW4V
zxqgYMS8UXJRvNeepFoJysWt7bDiaHTF59372lUiADaLAAnzvsgKdynulaNkADGy
ASTyXfPAbUGTrin+P1pUKsFmjuNS41lviT95V4qu1RBpWWMFO1hVC8cifm0oTmKm
4pQobd7ici92zHvgfr4ADcVB1V/TI7kxCnnZ8R1KfleKiZEDNlO1cKUiRMuKOrLQ
Xv00d55kwXrw23eSanAhcsuGolqbyUf0WSLpRv8HgUQkFZ/QpiDFbMcEGW4oy47G
8YN0GqrphnbX3VfaQvjYUeQGgPV2pPVUPYSRTNNGBuMALxGYHr1dg34vlTpU8vWP
wmCt02+MRKpSGvnDFaA3u1cFUmjRjO1baxs/tUl8JpIS7LBCD5GQa96emMgYK7Ey
VNAZQ01I5AQPwqABUY/ov+fBxN2C0liwfImU56ofVq/K7EY+7cXyLtu6KT5Bu80o
w56KLhzxf9g8Jab+0viCpHpfESfuXzqvFvsywGYOBI8KzH4QtHCHI0KMx6puPV27
pri9wXHrUB8J3noIXpg4LaN75Gfo64hCzRH+usJj8WpIEkXztfZNtMCj5AyxQtdy
tWsmfqr+QgHhhzcOHO2FyBg9qPrfkq0uFpxveMFG/faEcbPKhzRqOj7QtvfmA0c5
s60JPeIG3OauZjaydEywg6fa4UOE/wThryi340WP8ghFh+5QuL4GF+5hroYwz/Nc
RlGs5FCIKOhwp3N97IVY11bExwJGXOcvUG8XYSqqfL8vt4FhBqB1Pg3AaTC6g64B
TfZMulfvIa/If+kKpPew3HM0Pz7M4xk71vT4aqowlP28Y+88XhnntSiGOSCxEZ4d
dZI00ZFGCUjiiLVYTflnWOkbwM3TA/2JBvojgUGrVm8F1GmqVGwpLhxUs3vmEKlZ
jJmrAECMKR1jgkNub6UMrUBFr4C7ZgAdbTwZUAeYoH2/Ujfff4AKacf3D8InE3Q3
uqEmIUSrcj4Fg0p7FL8eDszfDhRAq1SeVz/fVNHnNFmkVrpOJEttPJ+tVq4Q8ycG
woKqmejumkXjGDkx1GyV8NMyWn2ZeS23fg/FDWGPunyqHkNG5E7XLWrDeTVLydq/
woj+Ohw7oicLu4+1Atg3x4a0PJLG1Da73pUfWB+uMsfVK+JSczCQqf6LWbThbSA9
v1paKzhRPpz21oACyr48Z3Fh6XSdIDP0lEQxepegGNWkLF0VkkjwX64PDJSMjAAJ
Yjjht4NXyOCYoYGJHC5CEjmKoCKgixu2eyR5joPYAmY4Gr8HZawEjp6EQblEOjLO
gWBRTGYfUM6lmBf/SpznyjxKtrB6ePV53fLMqfA3al/9iVhkO6St2TFvkmkr7M05
lveMalrIoQ1gGTAgos8c06O6di2OUpcuWZT++ah7xUH0ERQ3c+GSUvPCwnyhINBJ
SOMtt4arkzxkK93NYMpYu8Vaj4SA/r9bl6jXZUdgNRvzgjV02znx9CHiu8umy8Ng
uRr4dRy/TgCYt2PSvw+Wq81k/TQuvYbOsPR8C1RJLX6IGFMxZNOTMS0cYmx9TW1/
wJGEn3sHGYwiNvwG51y8PZkE+/bV1z4SkE9gzrxb0zOmkkAEfYh473L0JmzTMXOs
WY6JjUoBi338nR2m+U7GYguCkWBNTcLA8P4HdH0pxeeaq/R1CpH2jywvTxDl1sz8
jL1l64KlqzIuI7C1V/+gAVzBs2eXB0sjNpct+Qb5xQgLE1LYd8BJcCuiIwjbXDhP
8SXgLMCPt7r7AosvnSu+0mP/gZIqHReoO8LMiVGV43TTEelCpZvoNuJRXyC0xlX7
UPbgJlxODoQqqU8D91SfFC7iJkKo8pKkLzJ2RsQVTh+kDTse4b+usIziqXJy+5wa
Z12NsDWiVUsePUgn/Q+JZTORxIGmVq6iVGKtbHxeU4Stm1994p1xN3rGK88YCWRj
ZmS5XLYKEH434AbyjSz+/sDhBWyUUwX9lZK0PI/7XGqJh0KRM939/7Mi92/04Ody
FTr/l+IiIxHXd8k6BeQq1uSqkZdVnuLylx2bvLt3yJYMStl3WHaszOn1gInz0T/f
IjKBKxx/Wde7p5wfoNm1lIHhrhDiYSmSo3ApLr/aSzhzIfMaBp59PTagkmiM10Mp
5mDQv2wdiz+/U1+OPOpRTyvUcs2DNqRgVYk00rf5qc8ZqM+TMAjdk21HYrf0Y0Ks
GKi+ZkxrFS8qVXJNfQ+wTgGBuUtcK20LdllqcPAbzR6Q/8/oUrw2mW+/hhTR7AGZ
xPFOVV3OpXNnAH18ZFh08GYroy+wQDamatvrjiA0iwRD0DW9acE/mKsHd4ITGQip
kzpZIvRTr6eiq/EO91QxNyIriR9f25jGpamd8MEJOBhg69Orl1yuYYwSwVLC+dMh
yv1exrItznHax8G34KomexM8K7TvNs31IOVE5E2XmHUUiqceq5PLipSpundPMMQo
MFxD0s9On27XgJy+XgX0fuhZwrg2eODX8bjJxojYqmobiBfqlTFx/GWAxKccAgyr
sRQP11NzCs6vhPnsZVAc0NGRSGnQSKuQvww4iDPGS5Uf+TPol/2XOmrBanwh0f2f
oRe6F5RigWUITY/zBhefriBWhw49aOsU1pZUKhY5wPdc9mfJDEdoMX7jzXskVF9k
py/vpwuXTWQBbjGDWMEgZf60kRgQFLFtwxWxoPN6kVSlQItJuMmJ6Gq+WSwBZXYa
zYNzw+WSuFPUTdPiXV5wypdU1LLDaKyvc/qOKTqRgWI7khQbH3hFvtMylY5oRsEz
c42RvKClfR7G83Cd+WGsQsaMP3QYwE6LUCBWkmmfxnZc4TkxFgFFYtLCjb7SoRfA
Hp8qy6qv2JyeFNrwdwB+yBrOF/1OmSKdIqU8O+L0SJ4C69+75yX5o7BwMBsIro0g
ieXMpORKfcUEic2BmgloaShiQuU9YQ4iPYOHFbJQyNUlOgzrqmD7H6R681kBVqGh
Pz/nbDC74s8fX6KwncCIvYmH6UDN0GqXMCMjj/EbDqN40+5+oXxF8dKiptoxOTgM
g772TcJbaF6F7AAgEotKp1qnHPCrytQjNn3CNKM0it4CTTB3HWLtHzZfmrTjKy/5
egOIN5l6AhR9o74QNbrlm9zQQooKdMwjoIEv6TXOu86rgQBZtisf+LbgekKuf/bl
JE20DjA0+L1VKX/Dj9vpGvKPZRQCpzLFD5I9WK3LEICOO7ggiSX05h3GDuHyikbi
sn0myAjwhdpVvgpBGzG1qTLKbw5bajg5AKlmNpX/AVyykRHeNwRRPJBcpTA3t6WC
Ue951iCSnW8vTnpWUvhRPTwNEnb5+GXgNTV0Zk1b+7LWQPFNZyx3BIbIjeF0WRRg
s5g0FoFuDLoulFVPXV8NH3LGOr/VnUGVWIDd/ZXe8VaVE/0bWqYQx43rD2kZB7GW
NC+Ys8jyBm7lQlyeBQAaJSLzKB0rRV6uwTkRs7zFYsxI97QYPTekYz2wxMNRNjcB
gAxO1WVJS4QWUa79AVJA8ddvu8mbabPOLr7LetA0ge8AQt4bx9w0iHzVm271y3WO
xGhY7gAyBz19/OUAN4aLzmg78wRrDgEQiOgioGv7i0cDmz37UBdLa6Pg0RgH0du5
0gIiraz7qbA+gglCerYYsO+1GnbTxTytxxJmljS7gjUh6E5z/MEJQAVXxR465+W3
jqR6tGVJY+FcxFRVd3Qb+/gT1pTSK39xVLy0z00+LP2Hquwm6gmlO4R6F+AO584O
x3LNvE2I7xka4/LndGIoq7OGfrrmsgaDLaSDln/F7/DeP1aL6VieE9ogBTKnldj4
DsOLSU7nPGMmEcHOW4vvqybl4Xc48nfEuZJksSwyz5p9UKVHWzPDFjWFoqdafPtp
7Lf6dJdt0LFa9FllZaSmpnM3gTvUTQzUy8n7DSAsnnN+Sqxu0v6bZ1VB7AqWuTPK
kIolyqBtztZYkEg4hwTdUxmlAcgZfKMtBiaUW94L/jNdN6YFFqTweT8xnO2zvN7h
NaNF8bt0qIq9RHKZQmgItBwV9QrXuYrFz5fchHdAdEjK/8MTIqRXb+H4NSqEsJVj
jRC8u22OfIUnQygVdvUdyZ0fXaXPsCZiNeyZb1xKaSSRCCeOPruueRX/IvD7pG/9
jLdXAXpu2Cl3vTn3sxQBtrbGYS/cWMVZRhaxsmKygrfWxmSjmOZg3IfZN44QGR1I
meSRfWGvsEvEIqA9wPpNocmAwhre9CcZUJAW5OTF59IIk+r+U89gbelt2zSCi00H
Ijf5Ze5z5Fr/+dtYWNnuCYvD+16kkJUaETL48vee60pi0cfi6DxO6w0z1NIQj1Ci
6Xt/N++hviNdLshb0STqy2NQ6cGhEO/9iyrYTtceWD+cLh2AipfrKaI3amqs5NPO
nEVBcTjbSZrOosNH2G0t5YyzSmxxshLATPIPIrgvgtzH2wr8VOvlqsOUNAMx31cy
Uv60yFxraGzRkH0iI58ikQVyOVQc5eA9ZUX0QHKnt4C6qgP4yCCgHBmT2+nGucjG
R93sXYKNIyckt1iIx8EV4LenqosPUzR0fP6toAlwx4cUjw6nvT+R/s0QCR+ONVud
OcgcTTS6/uQ79NKb3df/Ej2tc4oi1SH8ULv0I6BPvRMUM22K+pTS9DwZL1eKWp68
OIn5veP5yqBEKDZRgQyjdn8tSNCH5plBb4YXu6hfS51RptiYY6I0HbIg1kFC70U0
+KcenbXJi+Y0GXD8eLs/XkaTlmLVYLdflGRdCrEkVQR730JXzYpxxiJWC3wzf/T+
lUEsufTRsSt1RH89FjBbh/9cAvL+h84fVpBfFlBOv8iI/Jsh44V1N7tUX4xb2nCB
XkQn7xnKM9vSTVR26Mo3oXqexXwlxMf3LL6W2r9bKQkwSg0ikcOHApm/XpNGeYzC
S8BlO8w4k+mQPDcQE0j3uRneLRx1u0iASFkBEPnROBzTxZ7JZxiyR1Ycy0S7sDrc
dWe2cuJ2WOaeEWDuh+UfD+fpPsGc2Wiv3W7wIyv8aEnYc6KMZYfkUBOjByXzr628
GwNwKZNuurTYUbPFFzVm0oz+/UaM9aieIhYH8iPIfhuN1wPrBVzQgydXYzVnmUTK
TN1s4/lWETzQZl8xL7J41tumDXutVuGMuXhgWiI1gVmr9z235wNQvnCTVsaa/1rG
3N/iZ9MKyX/zIcFmFOKVGheURm82kQCgY15PN1II5K0EL8SEBTsDLjrkOGe1Rvas
qh8XcYpfGN4m5xAoRyKmpYqnwsFepkZOa0uCboV6pus1qsvLNoP3hV35FA+lq5lY
40c0kj59yKCjfjURd5WvHO8kCU2l22Ki/ghRzajWZDtLM/E7XNPegtfzqduh2gP0
AGLXjD0GhXY+CZAwK55MdblcMm4YZ1OpXwH/LXW2tqEt8sfgbh9MIrsebAnkIdiy
occeqPy/McMj6ruhsuL00RNUk616BsdTZiHnGVJsOeHxoZqxBjADsP9XXsXoM6fN
P0kYwKP5MKxP+wEm4LVzvB6xQ1GJlYwI9aKQy9IRblmVU2FHjOA9g00Aio/2tYR9
PyBnp2SGeHgP4sNnC4terdDut8j+bJJweZHGc7q/BT0iKenqJHQeLkmAF768sSP6
xgb2U77okJJRpILwehSlJTYHToqgStL6kW6RlO21NJSVRgUS2Rkeda/46Y8PIHSy
/uL3z/Pw46lQ9S3/kgLCa348YVDCAgnwLC7SZGaRUIm7wFKYUgOGQDK2oPyvXz2x
gjMI/8+w/O6g1BnMDGmd5cjaMmFhJ02/qF42dZGlhGLlSzmFUvH5kASO9h38xSvH
ASvwW7uKkCEmoFhSnoo6a75j+29i3GO0wFJUKsu7ozGT4r1mfKeD5M+NvECLufYI
NsFULIG3jXkkRFbWY9OZ/D/KJLI50k9khO59UDiV6xYR75kxTl+TW2XqYEVzGWMr
wwYxvkNvAt85ACQfQzxU7fvwWp4rnmtmPlY4emSBhamTifJzDdUPLTuBMLyRzhGp
ovvpvJNZ+6jlk/DkyN3CSP3mwboLP/wl0DoGa8kA5RCbBDQnrOU31ORZn3Qtq7No
hZwTfwxCNoIranZfsGtdVf4ulA7Z0YamNwqQouSgifGVnBpuGLcpivNe6iUINQbB
xCIvHimun/BgrxWvLCM1Ma4yI+HvZ6E2j8G0yr6oSg1e2VnT0/XODs36HVD0s/qx
BurWKhhH5gy+A4fPFcUPVS9BKxSlwhMbirMaoXrhkWaNZNkxk+izxwaV3r2gV0Th
95ZEUeJKCpscbjcS1nFY2MyUar7xQp/39anrzvsP2ZRrXwpEfTarK9qVog/BSRjL
9C/JnMT3DaGmNr8UlYlvLXUaoRKxvnZSXrYyfssyiSf+iei02kqJR3wTCtnX8rlo
sIF0u4o5nwvjliEbXMW5/HKdsUegrCwbj0D246sUHnKWFqdOtJFPCMPg4uVkbE88
D2pRIm0M6jrhpPYxqzuhpT1eYlvrRFuYcDprRzPmkYALW2SnouY9/HqWJrVYaNoN
ZnrKzBPtOjEHIyZWr5KP9h3q3RCFp6mxLTj1hYyzadB+kLXPYDynCIoR+ENta8Xd
iqN9CV18+dz4SQNT5vL2pCszNOG0UI35dCSXN/iHe8uNppi+G/j3WMjwOHLwvrOq
0FZeHbZVPqpTK9OH2dEpxGMm/vwr3/WnvIiDiVcCEvhFcwRPgGjsyhU9C+s89fVE
azGUxML0dXFIwIlb8rByCaJhCiux5z1mukCcWFqLL/0fmaKCICtrYRxhnZyuFsne
OcL/sJxfWdz0bLJwBaSAPbWLYy8Am9NCYcBz5indLVtV8LunnhdGVt8gcawQFpqC
GY3i/SC0pjKgM70oIOLfDTvyT/+6vU4jv2hA7ms5oIugNtoOQaHyJzGv1USVquo0
q2U2upEhkKgjED3Q9nbgkvREIHYVIAn+X91vuBbrLWWQGThcaCLrj81rCziplW2u
Tj4XFPeR8/FDy2i+YegkpGCC5fHGJCb8/uP+RsNZHDPkkRQEypTaPpAXefRSkcGn
2cWqP+yq9Dd0gsCpWtsNnGYH8zXosto5IONmIrxHIlHgWVHIPiniE4lIUpGYMZec
fUsR0zlS+QBvB4jwy9EVEq4hpU2P2G+HyGsUU3/VUNGYtbCvfF2M0uyyEQQwfPP7
4sQuyU/YKjYBW+kTgKzcmVrQNtsFs4aJZDG8I/OfPgajALJbWBBXsAuMs0coeolb
LaDd6FHiII88X8qHvtLnEZHqj3nvjCx52ZT70KIlgSW7R3BRXQaZ0cA7LO/H2Rwt
xn68A0H6K7uTc8iggsYQafDUb7/9BoN1ty5Khp5ic/AHjLtr2TcXoCfHbxL2+vJA
pRRX6Xy6wnGn16kTIH29LLgFN2BNJqU/TnZA5UlH6zlpxR267lvYloKQ2/RxPKPA
AbqFETgW6UsbqbZ6OGYALDYBUzM9+P1dms0tkre39bqprJnwd+pGNdZEOALkaZnT
XQXELrbjWvPHsRFeT2d59mhLslKf6x6gk5u4ws42CdqckRWX9d8vQYJjoBCcv98V
tG1ZT0ayKhXPGzos/DKXaXkgzJhInpPhBWLlKNer87hCTdHMcUPtsPP6FyiJE3c1
wzf7/hJjqyubM+NHpNWoZcBPf8hj8s+o9BzL7M9bmQ/ks64ODgWrtBhfMwauUUw8
2E1RdVNJTdU33iwb4jojQE41qwYPyPFh9V8IlSPz9UF8a+hF8FMdUs4t0HW+lOUv
4/GcPzqunpazOEJOCeBuq9WFqu7DE6GcpWzLusbke9aIYq2MXeTZsObWYXtupJvy
xaX+s4nOOTiKDfIqH7w7lVS8Shwbez7JVLZkI7bYGFwWXgQyat7ia/md2bOCLV6y
uRZvOvEXLQFjCkWF5ezNeSX2/lDTcFob9TaeHVu8svHwx6Hy/vcQ2q8BK/YlcrMx
+7pG+kPOFUcl0sLS1yY3kwENka6j/Y3hAZuZztZ2mDg/AYhTKEtALEZi68jIVSu9
Dzey/lcZU54sBDVhWFsZU+ymn8tx2GoRMzIwZj8NF5w7+TYxaEVSqJCQ+e96O1qd
lSlIIvMwY8QY3gBfXcsbsB7U+aOpKy3/elaxtRlWhdoo1VYvxMzKdrdA7FeUUTb5
MOvjY6DrxfvjTFKMVDIAVS5U5HZl4m3jOhSvtkz0xIzMPYwPFiS+P49jtJpPRa9M
E8bTnedFWmu7Ve16ldjdeK3vBrzNXCMBuT/BBiohEyYniYPIBhe02RBYdTY7e15V
NudtTm3e+q8k3uCJWNeKInyN1QAFdKcZUufmH44Hahn+LtfHHmmmKn4gM6LABsA4
INEHl4kKvgglDVVZaiQzFkBDebz+llQTOI+RWWMWWXfUUe2zrKqXL6rRHpQNmuPE
PQzd/AcR0mPCvB/CjN0Uib7LQjlGUszBDRgGEczzwSmX5TtSqxFGKFnP3e9/UVOu
8Ceto+gfxj9wAwmyFzwfYcrZIZEp8OJfjAPyN1UhCt4m9WerKuMo6IeautAUYLFt
TigK1YQ4alFODBOYOMUyEc17PQg2Dwm55Td08BfIKaSMfDV91nDQc9ca+ifZlO/y
HrXFnaSGQHlR9YA+lK2C20aLhY+896me/NQ/Ybmb3XuxuSFTbLQugIRfEvhPwI82
5WyTYJvkiyPXKuuISGXlgN84uJQdA11eLz1SXw7uGiBVQLwx3D/Sv6OUFG6w06oP
5MeDMr3hfoFkGgHukRvUbTw/19+gPHDnTFuqZy99AvB7CNqBM4Fys5OnRldC9HX3
y+dlcw+CWXTFZ8ah2WGzY84FZrbzDgSOISYszbNTGtMIitpcJTrnfrPU3aB9TKGh
sDQVJb2QdnvYU53FZcYQ41J4ZX5PiNQPadSGfHE4Q1z00EEtKAYGWeJUp1Hk87DT
sxaTynu4sa8vlGGlfjoxaxiwa5WXfXyaoHBdpqdz//oAus9UsgteZnwe70CK9Scr
9LhpurjK8xBpWn8PPWVnBsVsz1iu4tTJSshV2v/AnIhWdFVDtZULyhvumzW0ruZo
HDGexKWnQ9iwZn6EF3+4scTt8KIn3VfdFIveyoH8pPjkasPqhOkGodxP0CfX0PBW
uVYCz8RmjJNfCWzFxZ1yW5PNV+H/xMqMs/njiBLpgbg7B5ncF/Heg+2HnoAinjHk
wIE4XsM2Nb092iDhSKXkflUdeSVpesJ1vGPM4BniAaKAVWt0stc/kW/zL3Uei/PE
mdSo8AQ3hpuLDiyVMgHGFGFRx0gS+A/DiqpcZEuMOrYq5q3m7ojRgyjQhEyqSHP5
LhIpqFBYKTFegKo1kyZPr23L8nNVsum4LFhnB3JTfgDqASn+nQeylgRx82qFf3Mg
2OqlVCM0xTuasFf6EJ66DSnKmlvalOxcueVHuAJJ/jDZocqtYDk7NdRjGAXEVJQC
eE40N1MF2drSfAncENjlYk1w39cC78yqV6XzjNOmGEo5h92+NC4EZL4BPSCuz4sc
rYyalRUSavMskOra60ScWagsadjAusdFpLZ+en4T2jmbtSdPscGgwoMtY/ro6LMz
hr4MYVKZOqXviDmSY7kDeN2xK+BEMusr3N7w9Lk0tkaIBw/lcjbIFDp6xU3oC+8V
UMI/18BoXg5osRSXRxvzgIBQV1jPacgAThyUIrg381Wh5GHS2OPjv1ktoXofaxS+
CscCM1v+hePhhCDsSofPkVc95eY7LErribUifEanVnn4t1npkcUfmyh+fyyf3Byv
ri+iI3yr6htw0D9ZlmD81cr3f7woC7gVdj+dWvdmIA/Mv5zgTnqDb7EK6/erd17W
lDKWyoHmo7C7OilGFqtpL1iDv4sTLDRx4v8Fzl3k+mtT9jOkQLIY4exXn1NSsJb1
ka7oiN/yWY6qGf6XlCDM4kPLx4cuq0ifFQsfWaTyyFhNlBFDUSr8f4aJm+9NlfdF
w6oZYuhCWYhMg0GLwBL1cRft9HLzBis3v1W+odYQXeuUt8FNxIEE27H5PvU1QB6W
zSF+xCSEF2GlXMxRm1EKIlf3hECyqyWkiuOZ2XRvcGZw6BPlYk06u788FFIo/Pei
PYZMs+a8suSaRIgK8v90aac/IwBLtb0mf48WRzAa4Hvhv3L6dAZwYY2EVtoeHSo0
AETle1riceHgnM3UxuD3QUqMZtBFsrJquL1sescc9NprLX7YEqo4H8kTHR8mLSum
wnwlYr0Y17bWqiPn/zNj6dhXljs9t+0wRXIlUwogSU+8L0Ffk/3Z+b9nHSPQEjWX
8T5YwrFQaQw+g+fZKK3Oj6nczXxk4dS/NGShMeg2N9cxbktWHTMRFitRCbPfskXP
GBMervCNPuhyW67rh3JQz7CEq6Z2gLudbBrybYL0Im+x8/8IdVsqT/3vK2eQi/7+
xC+cFegkQuUV45L+rr0Iag0+4ZGRNNDLJ50WwvOvxdeZYQnvpem/I0OxI6ibxWbe
jrcr0s4SSm0qGKpRx0EM5fkLcAS7W84nQp8WUd7wFD8zOqrs5EST6zBUkx59eBc1
mCSURKVZFeMHvDFzNKhY7hvfZTMQL4zjtnQJF3TYw2rhQyq8Sas/JYt9L3bW0QAu
1yJQcKRng6IGDoXE4js+1nKyQpQfL0VaL4YYThblfHl/uRVEuMzLS3/0IbTZ1Lsc
3Q/OOV18T2pwMFsVl/F6lDmfOKD9EIpOHnv5qdcXyebKhO9xM6lCqaG+CELLsHuS
UY9qrxv1m8iuxnVpPyOBjCwLC0GCpRCkcm8QMUdVOXiJlFNtK28KZoTHo3EVXZLZ
3xq/Hns6QLMRo2xYPY6MSbqbKxr/UIvhY1yGggWsPPSf5KokymAg1lI7Au0oqalO
74Y3y1EP16PPpRL6m/y5eQK0+F2zewza2GlAcKAo/vJd1D1eHEIEewB382zEDCyz
Dh5FmGOqQTNC0vw0f67Z1BkVJ50Il2VJVV8fNnSPGmS71Tow6hqx6rQbfux4volU
XMQE4c2YylNn5LapSNWQ3NhDjlp6NlQZGFofQtbV/jLiDYeK01odnSNdvyBxCKIw
wFg4jgR0Io94LxBk6agwNOpNqa4F1Ykz1AM2O4mbu64l4grzLAkqpdcqIQ3p7QIC
980BPGRYzU/RYRMdsL+mTxy3s12YygNTrUc711CRoc4iapuhupylxxUNGMfbIR7+
xwnbNi6LBzIAXeKq/oju7YTGnJwZsTtAlSeTz5yK9tI2SY6+3eC84sjknrIJDQ+E
AB0cOmSsJvyqbQhz9vpod4mM7K0cwCrDLqpKYGZ0vNzGkAd0UbnnnTPhCXmF4PwX
qLee9T0m2JHO3fbn5+ByqwB+FccqFIlxljBB9vCQaXQkTJwbcHc/zaooEpN7ngG/
WkcVF12Jwgqsd5uFAlLeWEJXWBhDZV/N4tflKMdOD/3o3rnA6rSxEUk46/5rz1Zp
G+QtDNNQKkBT/qdMIsiQFrUe/qJ1Pl1Sc6yCRusBpM4jOkY8GcMzAa7r9kXIKBr3
BaSo4I0kChlIQS/PXs02fbGLSiVAHxyOWAR+MK5+nyKMr4bAcxYC0yABYWllHcn0
5tAsD0481F6gI/R46KtdQWXkSXGtk7LKe79ASGotpCXL9Yk9o4OXFjCVd9GTIOFn
O2p0iOWWjCwRsEdIm6vkM80/f8yqyrlrK+VfgpSnvDhSipAmyqwSYuy544ApxWmU
5DWU7e8yHy6A5noCnxCvI/sRN5fkyuuj1j/IClwq3dNqiDXIZpYe+UYYTNk0Qear
SwH6k2btNy0qQVDgIfLA2xwPFO92eXp10HkLvUOzolnHQhjarFBcSFj7b1K/p8TG
PiijsxJ7/lW3Bay/GL2IpC+IDL28oqmT/I8fZ6UkjalOSwwjkEuQvY5ZxIm7znJK
L3UH7omdRb8GwN2+wOs1sZrieJGVS8aqiZU9nFAmeXG20cGTfHiNuUA5wRrkNP4J
IXuyulBKKxvHGTGXoCuN6TC2n4Y9mye+OHzObuUFunFp0BHrzYLpQ0sUT/FePAr3
uOcE6tE2tEe3THwTeKo6woq6L42+PCspdnO7u6Hf/kJNWUTvbTLBCt4COgYZVHhp
N4Ap7ZlvOtzRDQ6X1TmK0FTmRrFqn0rX3E/dbTOIUy86gKY8sZRhTYVir/GFRGqc
bQhxjcGUfgqUAuMMrX/9RnXihRVkCKVE8uW9zSf1ILKtFMSehhIXnNzGI3j/ocVd
JtH789HqlhS7H9FoCRup/gywA6joPqLAHmVADubvvpra8bvUK3sSEXiFxXJT7Azo
54t39HBvwArY2onbvqQEoQfJf9TaUu8kdP60hgW5a9jBMuo4Gze/cOisFgMp5JTe
Jodv+wkC5U0jPFcyAhOel3gfRTEegUK7qdyJYm/UHVFgoPztHo3LQkkmVnuT6y9m
xcpgtCot+/9TeIF6QDOci1bkoFGJylb+4oz0viLHYWmVxBFqp84XPR0xuwWqOAY4
abjBkBRaZt8lLkNNgT7CKpoB2KZn2VyIM3ME76lZdvQR294PSW9WLeDA8o6hm6Da
eQZoeiucprtqnfI/98WFgOZYHmKGM+pRSrPreaiR3VmUPN+xG28Dl6z/88tuh9ec
y4zRqre2JGFN3vQIwQ4js319PwvKzeqxYK3uyT5DfQETmLj9qgIgIKEdyqA4FMz2
KFABSHxxr/PKW0H7c5/XKAsM9/wHee9WbvfMDRx+6PNKNRv0OBfnCdxRwR7G2yro
Wj4inD/OVlE4hdjUtNLO4qlcYQzlyqI2yKbTulQq1iXXBdk2Iu/Z3+RvngShYEvD
4mSEWUtXsUTfHTOVjkRWoeE0Gm9qv3rZMbKNYuV+XPcF4HbZh83RQT+NP7ZmfuZ0
sLFMiGx5NmbNHY/Ciw1YPJCcGdEm2aJd1QMkKnOgCC78D7h5uMvA1rFUj/7APTXc
Dd3KRoHDZoNPc8JwJVZRknhxJfnrLvJnfqDXfuTUPM8aKFtxHJiXov/mJKXn35J5
jiLKn3iVihEfqbufLkkkin2LPjlbCj3OUCOBLfGfBvNT3ij3Jx4/rikbAg/IQgpr
8pHFSMC8Tqk6JFjPrYO0/QnUF7ZM6ZiBvbwKTqtt42zwVbJwNGgQDBpdov3TUCpw
8DuTTemOYZEm0SzMj0tKf5FzQY3dCw76cX6NBfp4w57lvi7MVpJW/pHQ7+jGnPpN
PtkSHC2zQbEoklVDdt23RqWrw1xYn1/Ci6H+tdvPSMAJKc/vsK8Bz7s01bBnEcX3
Zhm7R4rYx5NnNLoJnto3ML17MWf1nw+8FVFnb3RXpArzJt7sNOnBAQVv9M77GC/w
yws7LsjVCC8ib50Ei+v9p3YDczYcQgFgjjaUE3qFvAIcbOPgNYFyuMvJBJqm1SX9
mYZi7qkx2ooxzpSNOG6prxY9UrubSZHUinjuEmzctY5hlxt4uiwcPu2Sv20XOSiU
rKwA0VeZ9O8DoWkAto31NP0hVwtuCAj056yD3YzbjUIMQwu86jOlJ3o/baTUYChG
vBIQgJh6FGBOK2mGet0uFEkr5AZYBdaU/zzAn8udxLNByUSqMQW/hHMFJqwHyUz0
N9YhgWN3yd9GxoYwOIL6oljqTKh7k9fz80duYdFQpX8f+gXUfc2+nTbw8YACog40
5yIT59SQilYUT2bcu3oc++8ci/0j2ReMC64fuekPq0EW00YVjEUlJWMUimdThmWH
h4zR9YOhH3fJUA2kzPclDAVT/pg5ReL+C7YhpmaFnxIoiq5jDOIF3SmpAhbkm2Qy
DarqGJDs2FEnIBB0053St5rP+DTIU/aJsmU5TLY2H1nejE6I2Wc2aKGSs07LeuAT
59ekuoltXS4FtIR8qk0gfcCORy5GybuaeYx292pF1KUDtqDovpJr/Kp+EZT7asSx
TPLdQ2Ofe/lxl/wTxV6G/2IcHS95r5JpgMnZHYjjROD2NdQktMDxOuxInHjUgD63
g90HhtYVok25goR9T6E8i1vu/k3DHoRJPFIqgVTnl4SLfVmGtpCEGGsFvVH+QUpB
5IRGnipIweQO1wzPiBcZamePKKnqD2q9M5O212FhTDU8jA+BOeYn61UhIElM9uYj
l5H/Aus/iy4CjHH/YwWi1VV6/H8Sj2Y+2LTpSpHyNif5d9wdPqFObrrjk6UvASIH
yg/fLtzG3GfOZ3WQzvDmIEsvX4GG2temOUerjRv/ORn5tVfcQgIr+gi5wc3WqtUV
Gt9Qzkl2ZkKsJR/iKSP8d1O9Q4Q5BXLOI7sXa4lo5I8NbvIyMDzWLPZVWmEB2MWU
Pdr33/Mq/7I7AoU80p/kRcnp+52g+warKQzbws4Xnt9+V0zCgWyuO08xWtUnu7a3
qLFuVASZqI9kzDoHBosX934DoJP9O9qOSrqCTs7bn1dtUAugnUw2ObjBRig0bFf3
QktoheJ+SLH/igOcQF9/J+jOi+1gllKd6KkSPO4JG6MqZgCwHzFyggHGNAUXE4oO
0e9Zyl7PCLk3+sBe8d3rdXPg/IfrX0bnUwmSeVz2Mdi3OtyLddIgF1L8r6QsQgpO
gniLtZyznjA0+UdQvyn4mCh2cpm9dV+M3gt5m3uNhIgxpLowPcpSvSBBuHmYi1mq
xxhQf9l5Ul4XaV4nWhW0EjgxypowYirn/THiVrTs3f7x5Dre9hH877tQ5+Ybrxno
D3X+m/dJYshJsGcTYIgP0U02WlChSFhaNQbIDKjO+4Zrb5JBmTESu8y9Jns5bxJD
gOMI7yzNrtgmHQ0C3R1Zlj4TP4DyFi6kHBay3mfFSEW0x0BqPUSgTxOgzD4nhpo0
nBdUAdLPD1cowvsFyOigr+1pYu5J3/aRXO7L0pQJ52BZ5wQZBxnee9HdT2gM/veQ
Adw5ZCdrDSe5Xakf7Yug1YPRjKYZEi2Db5WwIa4i8tzgD+vMokKvRfQYpK1+i+un
kjdYPt+qu0H9vsHB8PRyuXEhyPYQJYbDxTdMha0oZILn+17I04ui0OBfy5SxJh9j
pa5N30c4CGBrcsEitqIkRwhF15kNx8BXLWD5kPMFelQH36TVN22SwG/p6vAAyQqv
TM5Q1dHW8TDy6hcovRN1XhZdW8qRPDNAyWa/2gOA864ns65tytoHw+zdU1wcEB2Z
bt08wwlrubWWUkQNxfA/ZrlxjtPJNJniJz9ixJ0rJC4VLSBPnvKJUraaiwDEGmd/
cBzf824/0HWsovVOyHYmT3ehfP7D7EXyXqmXX3Bqkj6kWDXgBhdSrkmzSgSKMy1d
StHAjubW96SP62OWYPFylxiLItdDfkRYqb5Nfn8AaLgYrICwRZv3UxhMWznKuAKt
lLAA/3Iac5Z2RId3bHOXtKis7TAQ4taz3w4Q41WGWw3tICYGHYzbreH+LkdRu20n
VvHL8IjCzkIIxlZdT1D3/lam+mY/OgHf4sLnD9cn1OawUcQBj0FH83bO4pUMBTNv
LeqGH6FdWTMGxhcD+Js6GiJndv/gDr/jgYwm7bwq7s424jHSOmthudXc2BUdsciU
bVt6rWnQS+5wIWZZ/8dlRI1MDDyfx/SlOUpW3Oa1Mhmz8yyxVkt6cSds3xuNZipn
VvQsd3yavY1jud+pcG03cVKRcYJZ9ojadBynLZqpqXkOr756hiuOxdWNzUtfKjxC
YNgG0QHbftRYJUXc749/4TBaNtdrTWOZdM0K881hz9OZYXfwlDM/7cN4fpFioWTS
d4BlBYE6ar7xwcBwU+H9se7rEatuRXKhGXoTi0akwsk/v6CJO0AAbDJTaW0ZP2sW
+jkJVMAgkM3txScc5c7Ihk3vLwQgAREjsKlkXSCsKlBUa548CXXdTqKCpDRsQUll
OnPysZelA5L6CCHRc4OdBBJDzNeRtFFlV7STP1sQ6TFuIMZyIrkFXMKqh//aqmgN
LGkgS2Gi9eNHx1JQPCbi/UNAeqrCwt8Y9XVwXZ9UCzwqxShjOgwupj6C5TfCdZqh
eN5yNsGa07+tddg6TAk+r8/fu/lEJ/QZ8TmlnWjQs+wj0l2jxbyPxJS4BojZ6ikA
jaaL8vbrzm8KhXqOUukM9cqqTgKUaBTLAyq5uoYosZkOfRr9pVUpioqFRKiAdDPt
s6y8W1x6qZ3G4Q+jhKsd729wel+ZC5L1j/fWwBIV9SiRUsPolkWteB7o7zLPvYj5
W/3OG/caZ3PKuDyIs3Eq+ujZ+8fF/gRWEfcmOiEdkfa4oqFL4TzQMbwklX9DNzEf
ZqbDeQ/c0MiLYd3GN2/jvV63XgjOPyvS9icSsjq6Ul7YmQS7S4HqF95cewz6CT9p
E4j4ecSV6GXkHU5S7N9pDDW3Vubc0cwPF0QxxyEUYDSwC6Vz2vEHUTUzMJ5ugDps
iRmJU1weKkEip0fL4dVQkreG/p5/4XZKaup1yjEqME8ySwuhctQlgku37D56womS
IkrlpC6WAV9znjweSnv9Eg62xNTs4iEHX5TGTBo9JmAx8j9mwpdhVtU+6Iiw+hyk
RpCzseK87aErWEh6tB6dqhF5kkXchqhXAFzLZpLNmLlsocptTOIosYUWEdhvn5xb
2GtaPH4LIUjuk01wXOsjuwKAvQdddv61Z5/Rsv6ivvvOQmOkp/rtwnXQg9gLv376
D8N6qqyvwlxaTTWlgSitK5z/yIDdefZehhMVQ0pn6S++Ap6nbRqtBVOsQ715qehM
oDUW+u3Vm4kcZd79ThNitGho8lvght8Gd1/oKI8pNXIl5a3YWU7szMywGOxRJM6W
yrnpBHUj6H0KGHUVmWWN7YFhyVChKdT+f3XRsVYgf+8o7MnQKaOa32z59+TBc/wA
OmuhLv7e2ibmmJhUAi7xoDd7ktZ31WXnBZ7iGRoVy5rzKU4wl4BFKtzj/CXpUp/w
oq/8yAx7CU1El1P01IHm3Mcrv4Y+LqKmfparOprMRIPJaJNWs3BOv2S5LDG7XQ4V
fAlJFP9XotuIYXshTQcQWDS6/EchsiYP3guClER64I4zFplkd9gsZSEDifMrNEwI
vGDLr64MJ2oLm6CBxFzOpkkjIu2+SsajXtjhjbwDwWoeYr2R4cObAJj9yKwxn4e4
w5ZNmsv5eo5jeHcGhXM2WXbUZJD0pp3VkaT6u1wJBfj5bBDCGUkWkaniP/TQMgBt
taTSghucnxL0RCKvGXQO1ZRUU4rXzzPQpdmgj01xENcMMXOzSnGEvEWE8jeVKeEf
DTEJOjI+I0gY+moncBi0vCNWy6TFya27/s0T6gxhxZedaXXhcefMK7qwfsSptyke
c6gDHIuSVLsq2jTT+CkvisfXzMIJF+SNaQPq9lWvOjN/wDcF8d/D5Z3gmRzgzOE5
Fdr8nCynCxhTBfAp1yQ3oTPOVK/McNo0Q5JSDC+nb2EZPateItO7P5SLm0YZKnHs
ADfYSLmYR0f2VXM+C3tWQ4G3h655QTZTwt3ZTsWhmQyiejTe6WpgatLfpMwuDzQA
IQotMVJ+yakWlw0MsLvvIlOwFffxfB/OaWx5CBOlxEdsdWC63gMX33yT71jSIjpG
4nt/iqzZy1kcyFNGcERH4IT8YIKKJXjIbwgeVnoBoqSHlnH6QcmYJU8wxuXlEWjg
MJcGpSgHuMPRfHUq74Sm1n6auTlEOSkSRx725X48Xmr+jmMhtcjPmEnV26+6lnpU
VM9X4MCUnUaz73ku6yBJkDJqisfBYGEWJlv0cgjUNDe5hAAmv1x//GE8Rgzgpx6a
HgboWlPH7/gcar/4En8gx5kUdjMHCKEmtBA19lz5VjruUZuGWYbdNeU7YdZ/BMOD
Pf1+WJ7qLzRbBNYvN1OizW/l67lKwOrndMmqo9Rc4ri+w41erNU6i01VS/3HiqYg
rEBfJbFgWdu7pK1F2yzxWaRtKJIaIoMIpd0kbAgZyGq5El7gDVX8X2IKIExxZ7VL
qB0HW6ceiEiBpQ2BjLcDVqWNNfCf9YsNC1Nhay3eiFyhH2aMUdzRrMhSN/NXriBv
roUu8wDG8gyv1A5z6yaU11eeORwFNtaFRD0FgjD+MNmdA3rraPhHkXDBBEuOsgsN
OM9/AfPlmt87JWCoxRY7mcaiCfxDN/H5uRX1kn0hXhdQEEqnikDmEZwQqI68EpgU
7k0BenKReVCcjdRWtIrArbPtKe/MGbMsDXc4pQTO5zZbxyWK5wxEnP5gIKT5e5G+
Ih5CuXbFqzkCfYIr8T+DK2P55iSrZLcWvls9y4jWgi6iKcTrnwZKP60uHU1k1XCY
qo7UpIoDsK55yV6fJg188SluAigx1suxRIzYCpLeBE3QHF8asRwhQCCuNVXgw57r
M9+sazxyUKCpOXSb2KmUlI/Q2593mD1E2UTCWRydkd/h2JycqAL4s62ywIRJ0PIG
zTUq4a1ubvXsbxo7MCzf1FHwiXk9YqhkCt8bnNi5CBpua3wF4AvX6DoqoPYxSun6
FwCpO6wNGcVdpMSq3aOKM7lbUIV+ytKibayxSZcHsxw60my3j2S0Ku8LsZNH1XyO
ErOft7HdHz7q7BLhEVGNOE92eQXlPc5iJnqPiAp16SkN753E49Rhyy60kISRCaOY
R00IedwOInn2Iwg4tZ0WARiby7p0W2GJ+4nCz7s7nakk3ar7nnR6utqqG0EdSdF+
b+7GSPuB26H0kOsgnd+gxjxj0P6s3Fsh/cXRa+U8NFGA6JnCucx4CxcuCvVLpLlD
dXmhvxLJWEUKo+/pgDQ186SggW2BR9uTebpssHMBG8UygUHkjrF/AUEr0TQ9JCU2
cKyLUGeEsKbaxlYJ2eOV1MVd1sdSl6lm8HI21wl64OFtYH2CIQyemXJGb808fxG6
SxNoIvDPPtrTXUL30X7f3kqKOFKOSk9jmjzFjCjqHg+Z8iyAWsF8MZdNcUQ3zRr0
QCg9j9PR4OgvnVO17Om6K/to1kdYcqY7L6XrovxFoxiwTwLRiJZZVuALtQH3je+4
N6XJAMRb/z+g7PNtVUjJACEUj8N6+DzRDOWEkKY86RZinmjtQ+UjMWTDHUq8hgnO
2CBD7zkr3DJPlbuANHvrcKEM9T7gs6SK8L35jESDQplFD9/xGXtQiJUI94BWbfyu
LjSrjSdCM1DQxXV9cOUdMR0WJWVHRoczwMLx+r3MtnE1Vtzug11B5HMsXp6kLuZ4
iXfn9J0FrSyPPaAO7Nh5833xiq7bV9MQ8Fa5RoNOk23h0RHllMekap8COBiceo2D
08sVWUK8djvwfMUD9ZTkrGoL0zk5RJBin0p8ihPyIaILFJyXYM2g+pu+kQdFLbMU
kGnxXhxBscm62E5/vyheG9cBc2L9Q/qjSVO5vgy6NfHRM7yALH7Bz7T8KG+0yjQm
6ylY7A4+Y06PwpCjcWdhCzunv+2GaKtH6Rjeoi+87WZVg/+3C9ZPr7yXHndnW8YB
Kjfi+L+2fXYjs3qaiTrVljdhtO7YTp6yU8Mg/Rufa1rByNbgEKtDYC/T5VKHv6MX
6j23cASx+ctRkDfqO2it5O8Yx1KLvc5/DxS9+Iyp8jE+SK81XugTKGJ/r2ztTIAF
6Rm3l18hIXWjNsK4+yc4p8xjPmwjVwPs+RMM+ovFWFOOklpFVb/CGyyd56jY9Z79
FuMEz4tDs2N8U3eYdW6S0Yym28xrVPAKp8qXb5HCLF/wrxkgAE9f4hZDVOR1NtEt
7p8u/3JcxzCRTS5rmTUm6dbXl9CUqZWFTNSNc8s8kn2KMiQbt/MQoy8dwxUBuiBW
E5Qqka8oASy1ciNxzhzUFbRFmKmGdNRqNshqZLtYhOYV2Z6l3NuEpswozQWeac6L
WMGQBnxa1FCSKKPWBfupl0jCtFq8iq7DGk1OaFgzm4FdFTfy/Acp+OjUm8F+Qu6I
Sc5oEBuN26cTht0Dt0fSx2qL/zZEHaNyBDkh/ILP1yaevM71dWKOKGdmy5Qq508S
5U4XWkrCZ3nFN3i01RvhadJVsnWd5tLKgpAQDWh92gt7V/2nzDZzt4T6dtHVlBlm
w59Hl6VVULxrwuAa7OShEw0+ThFPxQheYXhP4s9w6ycmCbqPa1Dmfeg7HHB6HvP5
5E1bKwyw30UVqSJVnxrPlFxNwbyRfaowhdnJtj2Ro/p+YjeG+Zx8JAuk+NOLzPUa
2Eh/f1w4Unz2+q/AxIhMZrlOIalGKtiuoLhCjc4EU5toxtQWnBh+NXJ+cY6PGYL4
WLHVuLFbYWeR0sBOcUfl22z35UheZh8eBbG995Ekaz5XY9RL6DWndBr89STmknX7
tGnQxu2OUs5TNSPCLYDW8f5finB+nIGlgYXXZehUEU/R84n0lxQ3YOAJ3F9bsaE5
mePbGDe7PkmJ79vG+LHWCRQ7woXbU2RSS13fMrmUru4qYpOh8Ye2vwjDf9nSTERS
vHhIkYOTEGvgF+RkfFRGsm/fc3rCvg9QU3jsvTGGQjuRQ8x2+C9iZF+/bgkK0ZiC
QGweKxpI0teMuTch8BSVZDzGAZZoTu7HDVRT8jZB3l7i29yDYZEMJRwmIqtrQgir
RtplHTBQUHiZHPOlEuO+wmDKLsdCeNK3rctrtJdrYYIe6+mOylwKmQaptfwa0Cul
tys3igt7K/1wsjHG2A/DGMPdAF0gtNusf7WbBE/zNWa7JqDZ+KXrJev7O3/EcuYK
bYqjz39sRl8w6Www1+S3B0M2lcJkUbyx3uHczLNXeDQDKX1pYErKjgyOtD7q6s78
Lv6bX71UxqBnpbob1iuGc/o+Woz2hWDamyNZAWzxAvpXMr8ORzmbU+VGdfPvPqFr
n7uADNkRadJr8UCqI6iWcRjgFx8gpUHlc2UVE0iwNyu44DMx8htto5rh9K0rA+EK
+gV9dzkgcXsty83R0Mmf883GD0BcK3nfTwptzCZZe3w8tXAtAUfcd8mXipWqubAw
XTnJNewpz7XEG1TxtFWPxC0sc/vtLyyHIWsfPbserrKAg0fW/0+5Rf/Nc5+Q7DmJ
azKIiy5jlI0rxfUL2CaNzija5ZTg7RnK6Z3ysav+WMvPUScb7zrSzzaTsA/hsdK9
2VkjXod50cbpi4JsWSEKH0IunzRpxgr9aYekf2vEGeZaPAqNZHpqhid4S8IN4jZI
zelXldkAm3XCJoRFVIIESZv69iLSRGJQEqV1ZFQXqzY0zIQUH7EnJMH9f5IeMjIi
fVytWvHnZ/QU2wtr8VShTVdRBCGrA8xA6hTC/tI2LSEGoNDcgVwkNG3QGVHaObek
DGZ904jwoRZ/UNHXSYpSkGdDv4Frq9PYga74u8val4plbhhYSthmy+HUYKTtwEcr
vyQm6gJLRMKHY3tI8gLdp/rbgs4WjmJCfUmAuaAFbyaw0hXcFrDUIbZLSPUQCGMD
mTTqiB0llhXLOt5gmopg5TI1ZbqDeGyQHOLv4O8oJEdquN/lgn4TM8H8W+Ow/y+d
A34wl8/KRMcfYt6DsuWvlMpuzIC4OXNdASeHayahgZWVYDZDcB5KZe2Ksb3XwVKh
evMvq6LVWH2F6HmiDv40njt9LJV50Y9VfCv+cRBLzQOWGrqemKXLIU/pgP6NOig2
wg98s68/U+dqQjap0NoAnrcFuWUDP88n6g6LzlTWys2vsPyblUQs2RattThQDX2Q
MgA1JsgHRk4T22ppD2QYwm3RX4EvgOGqV6RfkZ1fK7FuPiF2IHialTsG3ATzBFcu
qifX46l7J4MS0QPsxKlyGam40Zn48ONDrxkpGKG+3ZnUDGk/4NSQWc4MODkkOBvF
ZxbQJ65jMG+680/tzcsGkAHhwAgTrTmhoGc0VUq+k7RRs1fgu6lJfSuXeT0bFyni
3u28xvcr9RnHUbcNlUNHk/L1w+h3fprz1YrszNd7GPbwTDa4Qeh4tiOOAabCN+PV
SAFfmI0YozT+k8BFpf4vGiXdWOCb638mfNqUlovaPVyuRBzkqX/A9i45X91Y6nkN
hc2KHfq81UmLhIrRITmS5Ul6KSBoC29zd4h+ySe7T5mnLyRnqKm5vDOiLTLr84C9
R6GF/hj4Te4561TsJq3PbIwNpnfE1oQKu1N8a5Swy8jdlxYKB94U7SV0pr6BPi4m
f2t07Z6UYq3g+s+hYMKZKvohyYmtHKEVtJEVg9z8hzp9Wg2jzisrUMjz9UMpnsdS
C4Qhvs2HDXFuU42CFuXRuzeHz8mPDg4KV6Jvihx+p0jcoAx3y/Gznb2x2dBTNig4
QquYhGWOyx04zeeSECXI7D51rNFvenOSucepsJQARZIvjrAPMguyhMJO4J2SclO4
J1mZiWDWblr+m5PkOECGcOKUP+6UoPPWjdbG9S2JP5K24+bs1/xroidNEcaY/hPG
6fcjNHlnbvT5qqC7unwogFLUYMGoFJWoyyaXOF9XCqaEYjv5igpXqKzwhnggr0fY
oAXyqGhuF/vkpe7Sle0A5cjFtpFHEKLa8ZQrJEWcFnt/DIBsGIcBzbjUZR1kzPmh
bKMuKPolNpLuKnRUTANjjdgDWG9w6fH+NVS+Oh22YPl+xYVcnaXIxfoL11GZ+vjX
COljA69L4ID0rL4MwWsapZP7bR9UTOD/oa2nI+u9TAD2TX+hQsJ36/HY+wC8hR16
Dy5zzOOH9QF4aRIvj2LnrFjt7fVgKrdGrhHehm8fW7WAYx4qn3+I7A2vAcWjuBvS
iG3fI30yRaLz0PVLqRVbTLgeheYcwvfw8U9m0Kg9VLUUSQZOf7K15DZJCkv8upxb
LwsrLqQLw/NeQJgtWlbLQ+u/+70vZUSPo1zwAzfWHCc1eg6KfAXgdk1X0sGo4TLe
hq78ymJgBPLGZinL0TVEAihvITLRtYl/yDCeK8f7vHS+F3cql13gyVxgCuxtLudX
EaMz3vLFNaYbc2uFF+nVf+98ulu61epyxLQG2vBeLv5rNNV2nxHSpzfXrVy2PWev
eSmtKnAz1GfRIS785evC7I0YxiRPW/MUqjXSqLnIX0Ekj53pvAqyNANnCpzqgR21
ip/ACvqGTRjix4GAzRQ6Cr90mbqmvENi5tqqArre95jbpnTKui48f1vMXJ8BqYok
smz73u9XXrVPTU/Y0spvnR9dB50e0loVDtpXSK+Tb19Uyc7NYc5EKTB2KcOvXPLw
qsPyWAAPJH9SlbfoerJ17fFcVxnlRZGkXure8xbVhdN/+LXEhQEnTt2A3vAs0GC9
B8bnhXQbiV4vGGkL39EkhW0MQKIzBKhgPpJCiafQ+lzDBaPRryqX4bVsV27VVlfM
ukPN4IjldNfQcf1HjGy0Eq8YbKmU14UGf5cL6+18eQjG/CXR7BD3VY0SgOut1k5F
6qR8vCinfqRAxP5br9nLYxWhvbRLmmtQNPAViKe4Ujd/VR5NFXUcUd8Vq1KGzHLJ
E9gQ5ArOZnGlmGpVcl2sOx6ldQX5ciWvq/2M4dBqw3p1PXEDyPRIW8QNkH0w6D+u
kAKhyz0YJOA/n0J/X/82XlEvwG/+g9XyhudD1avS97mQ9YwNaOtRy/9PW65/66+s
2P2wvLyOyFJfHIhw7QYoPsq9JYNCBgd0ykHl0mlGgF0JditGIWTh9L3HHG9Xb9u2
rb6SeGl18hkm3nYy173w/pYPpNFfPqAf8fTc03jNeqeXGauacRhmYZ2ddPILl0LY
e0bzceGqkQGoUk1wWIr66u2LderqBNiYC2GovB0Em8AJpZQ+Q5lTUmhxjVJEbSS1
Su1F5Qoi6nW/gUpCORH1m84ajw838BLV1xB916MIKarW61bdhNLJ7fFfXB/0h3d7
rOSRv43uokAanReCapzTbT9wiVAC8/2/OfwXetG3+9XP4G0vpOTyojZsRomHStTB
R5gqkxmcR10pZlpE6gIWZtL8+4vAPR/ObnN9V0xDtm9iUkPf/NhqSFi0GYZ/gjpN
L1xwh0D3FzgKjCHfXd2jpylWh2aWvE/z5sSQyZCdok1nE8nUI6uQs5HV9CvwEoD0
PeDGUv3Rxdev+6QucOBViwZFBczGLPPDoDQvR8//3kuYzCxfiy+RI327EW4vLEiC
zGUe9xWXl8Q1pJ4US97wElLPKBWyLg6NuOiviE+LRsPsKCrC5+k0pZOlHOzu+ouW
CNSFLHmuZiNB9L6w5snfMRhHf6KPG20qq7tlRaYDd6m7lflXa6G3OhpKf/vMywXJ
cLlscaIVOIWdO2RembXLlc5ltt201Q/QXh93cfsYYHHTayApSt64RcZa9DS3inJe
CS4qswV6AhV2mt1/OL1qjoRUsUiJkhLxoVgfES3GMHhRoWH+21JLt2F4WDa4BAf1
N4uT7xwiRqONalME67iun3E7MBRtGAavekiGfNVFr39/6/kdGn9S1OSqmY7GMp41
G3HFS4cEwz+1DE0pCN4rK8xkM3DMRh9F3dvEVGOQ9mVMJhJKk4z5O8Qe4RTbohPg
gjzX/GTtL36vd3jH65ep6NxKwD3nisBSs04iU4/MTSSCCbluT+g4lXak0/Excqyr
ccvQ9fmP2AJbul55QIkW1gHubmkmFzzI5hVoKSBJdzk9f36nICp9UAxr/0TQgFVo
UqerRoHahMVjhCDa0VkkNhV+Yyf5juUFlSGzEVWlyQ96grbSGPipidOJKfg/fWXo
VQmHxsCosdcmvsK3WL9nMoAm3uD72Oj3vm0DM+gXV7gNRGnnegS5IXji4Hxx+70T
w1QBFIhm9v+QWyZSq0wDx/kLMlZn5HLoyHhZMp981/V+qXoeYLUYukawBoJOZ/VS
mrGH0dIyfctxxGECD1/8cBp0UWH5DSkWS+to5Z+2A2UwhKqeffDO0DcnGB+rnOQk
+qb0oLsM6KlPdA6mDg7ayRgVc6znduJAr+eJM1o7fbOgMxVgMDarLhzIi0R9DDP2
2L2VjHt3l+OH4MZ4UuMEwG+e+ow7Z2lu6f9KpN61E3ZvxIGScye9dtleav4Kg2B8
qQGtfhsgnDtfDogR5bv8mHFS0JdTdVa5tEXowaWVS66rtGA6AWA8ZmCP8/I/YZwS
diZWu6ODj6EjPX/1Fw9PLGbJhbcSmKQ3d08Y9/u91clPhZ3hlvLT9sAtJsKAeQpp
QRo9lZyXsecE9cF7YxecNTjXK1+ErlJ0MSVP8RNbAeSftwbBM/tx97BS38SKUlha
kNObZyAjvcaMm8QGLFGSrIlVSpNe2Nf3seJU6WdDUHPHHsH5oY/By/aCjpDrRx4X
oWNwB32FQ1Dy5NCoGmabwP+8NVjIeyKhbbBfl4BZu96WnkAr0VhNYZWhbjcLBNfE
QhPg4CYnTyjso3qSoZLX7BiBbxARb8iIkmLhfs+cy1UHy88Y8LxatDKOYzA3GaJr
V+qBAJ44F0FIoegSNGV4MxQ31mrsLU/OfsgpUgTqFCjnunTIoqjTB7m93tAXF6jX
R6PfT+zQ+c3Z6/2iBmnOP9R4REmuSHBhys4SUO9MNpgH17M2q0QIElzqRA+2C330
F1lwUq8mhoFAaB4vq7fXCeMB88eE837LqZjnNnaOrShkcSml0ByOwKOTo0js8qvT
v/UGQpEMqQQHQc4ULCXPx1mz9O3OS0ZyG++YYOPjpf01sS/ESkNw8nw3d3M/EW+D
mVqGzNc0KcAYaLpPWS0iXFP4Xcr1aJ/jLBuoCwfKrslQ4aDTjW6pgAAGl0hUsVDI
3BiM8NEryRuxC9m/v1QoB2CLdJZ4iybLD/59uZe8q4RAhet72kbpXngOcZPqPmFR
n8nvIbO3rkxylCUWDpnU0WyKPkWWfPqMZAvdgd7rN65wGgIm/elr7/y4EfaVNPo2
XJfr+EG3I1tcAV0jlg5wQaRHAHZ/HWKxzRTneve7ewe1S9fTGOApmAIbJEUz3Igz
3J7vwOWwZ2L60d0ZC1V21cnAlc35ODSzOygqwFJdf7dozAt+8hN1mRoImgFx7Yce
2APqP0Lme5hd4pC6G+/SboNLJAUqrisUWVOLG+pb5joOCaCFjdblFDp6MFVK41mm
6X8Lnc31y/+KLnawWSR7xneJCjDoOwxmC5BkS/aS/jM13eR+uITKwPTbADwsgWvR
OhnOrqQJ4/dG32uQgG7IaiB56JeyrDsMXzlMF21UplvVLe8wYNLJxKSCfVPoExRz
khA5fyFwCZoxJ8JdW4tgiWeGUne16YVSswtcGnLV1HRSMvjv+vAjlKtLS0gVy6TN
ud57XgEpVByqCiQX9s4qM9d6WHtFNDKLiRUbJQ01OhhZM7Z9+nDUXfeFlqzyX3lN
CqhHxAS8z3C2iRVq7DhPTLcfBFbyVZHNqvxB/4miHcxVIq82+QY4zEmaO980vm+h
IWuRgekDI8N4Z5LQ3CQHIs6fPJUl9lQ+1sJWwtNofi75sWkNXtlH3reObHEmUYbD
PeqScWo/o4LW3Xxnuc6kfU98I9s6S8nkVFvK+ESHFgBSe9+F9589ttDonyi8+DPA
9a31NGixYLwFkENGhygdREAdMvb6SxSAutfQHUxs92AUHuiFOqCqKVWujPz6qiyU
ptQF+S31ZDkbfQ8a93U20gjiJr83qpt7Cznk+D+4NuaUa1aOUPuMqONOobzpoyNy
aGYXGqkcMGpM9SBwvMUYcTjg8mwbCIrh5cQYpCxtar3a8xJ/SSOznc65IzdpaZQ9
uYCJsYaPMfJttw3i7+c0eUP4CjB3x88fc7slXzkEDgAhPGicse8zDq/Qx6u/z8gw
dAtuOIuf298DVBfDnaa+ds8zfZOMrpUiby7vhcPD5VYVmORHSF9B8wx1Nf+bebUp
XXyy8uUhNT7awCzWSTEgljvEks+zB25A/FcNkdBSJlVgd3vhIcoa2ggplZpQIWmv
gUG/jkEbnEAY8T+pjLY53M1VNonEGLIZpKs/xHtANmFsiKw8/MYrSJeODd/TUE8k
GcQY4t0hSuquLtlHItMKA5RqaElNyDy1GArtLIBLk7utDzWe4lDBB57FBg4X0RdQ
581pdYnv4l9mlfw8MiFUZEcOVUyHbRcFH82an3femnvECopNM0OtnxWkfGWYU0FH
TF1imBHiCZzKcYKsYl/Lf668KG1JdtkHQ3xBgTCDziu/fkq5jAITzKxC/CbJJE9E
WxPgDPuG+pEi+i6SDxR9H+kjgPkeROJbcV1vTO0uZEwqBDpgJfPadsOWhkY3Rztl
uzwaAs/4dIGUfyE6xXw/+OytwWQbIEvMDJToC751qGB77SEhFfPTArXQJMGwnE4p
qbTvU0V01KBBHAw/AG7ZF1d3DNKAbWR3A4nBJdzjlALYUcwhMePl1tpI59syNqtZ
DMORMG/f/SVmNSZ94t/WTcmiC5Wo9XEcBOzRq6e1Heqc33haMESClbNEmCEl7aCg
mOIcGsuAfYmbwQRF61AAWAGWIL34WZ4QZvSQb/TBjbfJ91t0Qi8sLNEriHLTGW5k
fSiY0zL3EvInxu1kj4tykAxSGpR0OQ0hi1p6eE+Ti5eblb4jayKMSjVivmGG37b0
0rNwR4k5O1G31GNWRV9uBRqfTnHwxWWx3dcGHGHinZ8dJj/JPeXQICNLZ9CZbv9Y
XJoz2Ty8ZX8mta4xbOtzVbgU5Q9tXjtumLr0DT4M7MMlZSyA9CfWr3b+wcMCNY5O
Lbtp6bMEKhuRDeVN3+8NkvnCVLqBDJArgKuUbJGB80FA1+Rr0/Cj9M3/oHXtIqGQ
NPOM5G86XiFRaJnNrVes20dcZw3K9rAuVacHiuVvwUR3hv6zy+Az/sKVYFVD7629
VHbNuviDnV9zjMeCVyBP7l2SALPuRxTQTCbiCD5+BKuC+OyWrqqAtZp+IhXnAIO4
6EeTEV7loXxpRc4eg7ZWxqf77nZ6tVD+SxDA8mZ8BzGIWNfYpkqrthqrxQ67FWfV
+FJVpbGCCXnbIs1InCfmOc2+BsG0QJsrIcTuCtLpkf0xtJ/OqwH/DH0d05au5sIP
jdZY9U8u2NCqLjflEqcPsRt2mhPdQbV+OnKCJCRGKvpAOPjH9wtbSVYpaxkAg2kn
xaNTgmzpY8QqvBbbnw1YJsSvKQVdx2MIpynv6vLQA238SGspUJ+HabSR/KPxGY8/
01/imUPTKgFUomhzDvG5lPM9yaAsnlkEu6/XWPi32ll4baFqOEhLE8EDBzrz1UiO
9S7kBXdWQT57ws17jDIvpW0C6gbWwXLu9PQAt+zDoyuLzQ7lyKctyxU92vlvT50N
8j5qHMMxxtDTv9rnOLSoiDiYBaIVKb/TMIE6QRCAwN14v7S4wcuG2KtQBFgpiNOG
Bxxo/u34DPVRQCp0XYpjusrSWXUQTHk0xjzohSEpOEZ6cnFKjFyEwHnlZTplLOtZ
vZcWG9xOb/BY2ryuivHzOItY75toG4MBIGLGJ7wwtTvSI/+vGrRDJRtVR/nTrbpD
pDY68eeVPCnSpY5i8SOqFwFr9NvJVHV98+uBPpiQnjAQjBtTK9iBQEM+1nvZ1KvA
tQDd2zljNaMwp9yzJ5sty1mglVcZi8UnhA/l5TFbeFrw3yRpst11x60Dkkf+6jD7
hpmgQ0ZuHDqkqgGygQMgyuKoymuOpVZbByHTUEEWJA7/3c+vxTiw+r2OAyYMXal9
v2S+/n4kmVwlE88Qc4C5+6ShbnYJ3B1qgr9J39aTSq8MtKnBpHyfRIj2daLRvLiH
s6lRD7Jnp+uzDQWngxOw0MHq1v/hjvz3EOOjDFaG3KTHA+ANoNZjAqog809bclkr
mNTZhZqYeA1M53an3YMVZ4vPKpRyByZk3ViFtruvVPiPl3Q7AbSpUNAVRnwuj4p+
9TddA3DEk+jeasHXPDWGh4y+vOw+SKBqW6FzD16+WeLTJ019VAX+IT/RA8v8IU49
0iKII5Dm5R2RCBD/ZhpRKcL3pXS9u9gLxRO7F9gz9AhfvJM4biLvFdb1UPdeFq4P
iVh2hoKLtOctLXm9mENF4z83EARCzKaZGOhXVSsQQh4KLVOm2NXgQuTc4LI/4aV1
pBDwMZNsfvEypPJ1N1XEJ72XkHu/G2i3JW9ihVLFd/uWU8RGv9DEihKGbQ6JL8ZQ
wrPToXCFwrqRiDTEGpHNpPeQ4nKkXxTxwaiqBO+q6DHgg4rrl5JrvCyQ9A1uxT0/
NArYE+VKMMwk2UJ+dPsXfV6OWTTQmdflzEbXvs7tipTIPZjYyNYD72mNUu4BVq64
H3C5AYTi6wbcLBcw3BEuuEknQTpWBnJQmZZa6ufOT4iqXoSyekQEveQbOHHILPmy
i2GJfYKm2NHXo7aNuxeFSuee1577+GsatR9ECUtVeulRLbtkhrGNeqdZQjcap8df
t6ZkPC11DiCbXfiSb6Fv58m3MiAsdkrPyltcFfJoMG+y8gV+7+bLuhmAqEG2myKM
2YNtSBkJk5EuqkbmSaabLs38yHRaxQCLtIdWpFrskLoJGcHJQjTTteeawG3WTi1d
AABJ2LNqiCyQGU12cjnuNFg6pFKyHXk0kym2KYw9XDVz2oo3RtQFSdqoIrEfHe4S
EFVUwNDeSIK1ffviXlBIY7jNhGmsSWO1PEcoJjI2Bse2205iyURNto2jpX2ejaBJ
vyC+OQ/SpgSHzFqmxUcTJHrf/xresQclby0gM1jH/Lr6TALWrS9unwCzgGDL2WXL
NkTo6UKHau24mfSGesdiKP7laJ0Is0zr1w3//NcuRsZDiOAF4M/w0hso4ts0tzN+
TDOYcpsugVyOAKU5WqTEOrFnIxSP0w2jkvY8m7OQS+VXdbcBdnIttoL3Cu3GsDh4
Zj2kvdBcnULcIK6dZzZU7H6BVhGTRco+Z3Zy96Wme6dlQ4C4kyWlXcIB2Qiqeq6Z
h3gMPFzCp4303plqnPam+NY9Q2hDEyGdMa3pECWdHK1k8yylefqPksxsvOrtRVP0
0b8iVUYR1obnu0Q2MVLImyAoC++bTrXHcGpx4uNPAyfmYwkwnaTFOAHmUmP01N11
P/+0Z5GENWeVT4z89qWmrUCJ1hmZe6giNK/v9JzbemUDRQWQU0FcdBjz2duuYe8G
ZASJmGo84XROkH97LwVJowQRLGmUXlxSOCvWG8cc7QYOD4I80OvD6Q/p5OyJO3nB
1Wsdyt2p4vsIAzBmABilDoF3//muXUlkiMYpQptEZirYyMCa5gKgwTT7YPcyCN6N
Fjfj6AfpwdM2wayF8jlXcgkQkxvLOefJwipeT1uLqbhol302SvOcmqncqe6ZrCgi
7w/d5qFSHheXbBbbn56PdjGtyy+bRkAEfwmaNN8T5G/tQts0PT73ReLL9dBuq9cx
998L8C9MmHbGjBCE+AvqaHsp+fH9rOiDg8v8V52Bap9CgV5Le2G6Rv9Qi0in9jkh
CrWvBsLHjqHx5l28O6T0g6Rd5x9Bzon3MdC3pWHsG7F7P5AXYKgVJmP6uxoyI9ws
sU66SV5z0j5ty5niXkAlQjdPdjLjvdfl8TcRYYtQMdaBPlm7gEc31MqB+TCZ9wvU
FhPNdG+FNDkHdo6htAIP4Ztitb3AaX1KdlOrG7vWpjdgVbnwwkKyc1plKLOqXRfX
kptvaIRuCF/nJCfvaiClzIHgWZ9exUC53YUXUAgiLTzBIhItQ9MTava098EZYGPw
kXDmDgzft3XYSrXUj5uBIXcYlOGHb24BSoioRhAl3+LkNo8C/eGko3eYQK9fmxpf
bCpjyCcYHS9EzYkN7aUqDJ7c5je5GsYxR3uppqZlQNTD0rRBHJ7YFxjLathUaiyC
L+WNCJE/KjCHN0UZqjmHQMD0Xak2UooEN5eX7p+MITt2kWbo602loJXkRUXW2/da
2lpomdZOMvcn2m2tsUuyCam/FG8an0IkeCNRolgegx8I9ABdHHjC9/L2yKCofSte
Svs7rAguylRjaCB7g/S1DuVF83BeDIjmSBxfc5U1lJao2DvBhP78Wfs88zPDBWWt
TTEOIxHZ64iR0QKH7GTIe57AzOvu8ibHLBKJ/bIuQA7Cmi4rgF8Ucj59wW3FN9fr
RImRaaeybOwg/8XZbeIBIkAo0eqCn3mukcF3eUdkT39MadhVbfMaUSeArP0tzNWw
gPJbAO/JsJMuKb7eyoz5NTQKb7efKBqPEF+HmdvzQw6OgCjtVkRJKZ0cMvwMX6bh
hfudO/60+G3JZZGYiBVZ2g5BdZvIx/oAN6zlnRwkY0Bk6i8Hs8tix0mNIEg/VoD9
TQMb1t/90ibi/Ql1zoAGhWar06Vw3vBg2w9+wpRYCqD9IT+RNAV0j18Qi84TbLxh
6bZUekQnOQqci1atcsJJgMCi9lpQ8jCsiTqhTeSIGyNgFYxcXybhpnP5q3Ck/K4D
Swaxk+hRgIZBenuNDFAEn0R0Ao0s4LG0coB20jvojX7wSssTAxLKVwe6YY0wbcaG
iM94H23eBm9sB+YbxYsdyS9gIGpD41IXM3ShdKQ/95BIhs4aKOsVHrrksLjlE4Nl
njVM+5fNQ3EkPRPmc/MUvAvs4ePHsvIgkK/CphzMbpitJXpqe0gfWgVYsONPqNp8
HbVTVWlBeYQ4hioR319AruIDKhUETAlRjZLnjJhecuXMiRcPRmrUI8odfQffi/V7
iQIvdzX3NdVrmvVKanEtyJFdgLvz8xuBly9a17yTrHH/QTrIafnF++YHDvpsTW3O
1D1PExRfFDXi7tU5NjllFQjCzeqEv6BsURsCw+Wgx1oVfwx9Ov/E9OX7J5u4rthO
9W46MUds3qL+T8w7ud8gSKuuu5t6/aHmn/0foHJI5rlXZS5+20HAZg3dBJ9EnTYE
ij0CmIuKnAO5PkA5tRNamDIK6i53xUkw1jsw5Rea2/P1KqrcdhOUsKRzL2LAOX65
cTlABECMLhZx4LiblIj9fW2QpvkK1r+8SXrCLd7jqB5IfCUedjbvaueqtjtUbC3L
ls/S44OxBD+jaYsvl78opPHcDyUOsy9nx54mQFf1Pvan4Kxb5QYr47MxHsWCxiRU
wyxoMHiBEjoE7xGxKTE00nYT8Im8s98JNnMH33FYmA1GX1W6c8KADu7NsSzVXHwG
996cQizz9WIR5lsUFBwpR9cvDIUJVZs5AFIJTVJGnU8MDoJStxRlvN69LvqOWOGd
M6g0eXWXRpGHvFLM7AYGSB9VDA2zHZUyklJh3NB3/HPIsBELEBiPxi9qlVt7IXhc
GolBPEr1mcT+vkjGsGxD5LMvKorOUBGtT+Pvevz0Pdpqa7jsFjd3uO3dx4DEOSZO
O1ctDwPVuZ51StPfJeTDFxAC3PS4oNpbjo0ezLhmY6G2/d9QQJn95YHUeiN9gVaF
GUwNDrkaSaQW6qs5MpEpAK0fmFySx/ngJ3VS1zpI2FLhL2nO/NsW+sCCTQXrO/1F
qO5I0QVVpns+0ztLs4B11qqqymJkh9+FwkUwOLMs+v3FVlujPiphMRGbbOuCQcFU
uFg5JiN0prU4UOGGlk9FpzQFYfzX9JkxRIRhtXQGYbY8+NK740CW6FaMbDXZsjRK
jlVx+SydQwoHRNN6XX/wdg4njHcUu7UOlwjuAuhnfh9F9/I04PNBNKET3+9ieNo9
MiQL4C5lgXso3h+V+ICqsl8lw7qhLLLnm3Z9WWpnBwTHw6H0HOYw2ind8yDHEd2S
c/9JVZaKb44AaIg0re+B4uGPQ00OpqBhWACiRoRyQOMo/8kLtmsbA7i5gj9IZFxh
QpIESIBwzd0mIV9/MkeV66ToiDbTYomlcUiqwDq42tr8gGj/EmwWolzjduJkmQ6y
aPhlDPlOlt/XTdUIknbtZh/wkKVAsbRdGI/id7o0Jus4YWK7eopVAI8gTDGdcivJ
4aK7+k3VrhDG4+Zj80S1vOZ+QigLxgbNWbqUnMRpCdey7chQu485DZAJa8eGj8jU
YW645IblkqhpiioqdSCgfpSaGE9KXDK0bNnWqUeZAgCnJyJnPPeexsxo7mMPUuaU
FJsfw6gct/t/xIHDPtroUCDz4l7Birac3HELDUcfO0/gLF+nms8lGMe77MTrUZ7+
/8fpvnsFidJBa96/9WvHTWm/omsmGcmlfpoxUTwA4DzzcbEwwGQyxRlLOXJDDZ7x
ED+DKt7C7YIv+eSJY6aNc7nli0H2Yr58S8yu2caSyYdrvekwjRNi5Sn82vaFjIrA
DCFUUIw0qsL6aU48hWfZVTdgzgSxFUi6isUuQg5d1rxaUhPstyFk24nUE0WR5hFu
PKOnAY0BhXsK1ZHHjLmZ213+T09xPxvkcRpgerEzzfTdUi53sW8vXe8GiR6cf5OB
sQZOJtxwYZaOM+BN3J6jElGXGxGhf0ROUMkopYLcsbMZaeWjrXgiQNasVc+rSTg0
jKEQtGy6/Xe8etQ3YvqdWxE65dhXcYwZm9l+I3zXwPnvssOdk+OSuVHQB1QSS/Ql
auv7ql11cHnaTTfsWbjKHpKqVycczyuZXd/C8j3QoiThdYhL4yzftdqw7fT44vrY
Jg+K40R/5FFH0mldPmrNjxxOIwTDncpV1ijWNdcG47oxkVexeAduj8RrYbcg3mbH
tJrGr9GDA9GeknuGAHceTyuFmbhv6d0ML0Vj/9T9VA6epbIgRqc9IKKViRxzr0Z1
Zttdt0ExOUpna6/WxsOoSxApfXrwKRy82URMg3Ig0T/q2JTIfxYII+nuK1dxCvzK
NFlAw096uCUIdGFZQm/sZpnNGWs//x1h5qZo3yUipETcMPk5yJawGC/6QDZfWJwB
IclYJLCB+GkiArFSY8e21D6g8ka2STW6Ebpdu7f7BjLs8QsVi1IYhxN0kLtWHM0G
T5b9PoNShKexsl1aXxlo7oedDQLH5M6t5qjO/Jz4f+XKgfa26IkFVwCDN1k5aPrZ
XlK4GuZI+JZ2j/HozUPdqihFoWtVzND1xdeHADMjGyguJuAPu672uvjiePAaAAC2
1mzrNZIxTGVgx7V1xvvrQcQKuPc2eWs1f/7LlZQzC5vP8ebt7mLbZUCVXxABCBBw
qIxGEUt1ugVq8doqpfQhE/fJ+KGuvukg1Pp3fvo4t6rkz+FkTBt8GHVY+0lQQSCv
t4xxA2Vgd+EWz/A83iwZZeN/0M4CGB09CEpMzlk1O/kwhLgTcBPK1DQwP9GLmwln
bMq3bO2thWBL11rAlXiCE2D3btTVhCxxt/n7M1hHOw/+jrzTOMBMlZ5dd2ABTb2x
Z0sWc2wUKswtwQSI66A0Zi+zYpS+qdbPjhoFoJQDGw3SK3eZPVC3rNleq0t8jm5S
F1pWP5EwbjRfuBIXjArFjxk5AdY9XXArEDr1W+4swMg9ZqaWjBlqRf+QKSSTc/Ix
47EZy6/mcDapc/CVeMYawIReF8E+12G0RJrlW8GNT1aT81+XFv+typ8W1M4f5Qj7
FfUU7l6omwBIHFa9cGH/OMVO7s/ikugaFlxn8hUe7SCI9vTi1Hlm3xQfYVbPdKEJ
CQUEHbGKT8ssF5H/t/Ug96RkevRtCpcWzBaSIqnIly4fNboLfExScxulokvsQ3vc
NrXO3VDXZOxU21ofGkqfqQbG/Vm7JwOZSQmJJ/IopQnXTY+japmuB94hWo6aDk2k
AGZwL51QzkGFy/15eKeXsPoTTSu8H8CEsewyhBmtDsCIA5KpNAYSiVCCdxtlVpU6
gyNsKWcbk2I/016qzmMueB+OAWUSi7R/QuKQUk0u3APVnJy1pWNiwMTirWTHOORC
GOJxVxANUKMJEgk2ZW1nXrcWf7hgjPmui7ksOj+q8yUZJ4+jLoSz2LJafll1ZNCs
HJDWOHzYtGcC5IrqliOSALeMw2l/fcN2dFA7vlslMf/erqq2XQ3kHAGC57uC4u8Q
EDyM6CnykWrxsN/gmp1pBtZWL2s6m+1PSvguy4SCLKQD3iANfnvU9YYPCiVN3JiR
kZffyxG5SoqD169TGyxvTzL6Hs/dF40pq9X2CynFz+UINTLV7BHuKre1nMM0K/so
dr5DLvZ1jH+F50lajl57vsv0XHqluo+H3/IzIeZF33oju+UoEG7oIftdRdy37A9T
avUA4kv853JOiC5AGVWbbiPHZnPstlf++nQ9m6mY7+c0in6ggHtA8RQC+U5rCrFh
cxb+gKR+ggttdOT/mlL8XIsX+BKausK3z9gYt2r44GMZz4G8VAJ+IyKzkn0f67u0
Ws6MkFeC7RwMDZ//+BqmKrR6vXCrlKEslPb8fpVz/55TbKQM9EL9/NgAHi1YsAsk
4TMJkp/YZi7SU723Awx18ON3pK9cJ+QcZC/+EB14mI5L0bcrDSav4liNUHvxhAHR
uGe+BJFpi3jd0pom4GVPQ4kBCGabFZ6DmLx8IPGF/vQ+CUqsq4oBOtx+lHh/E51O
RnHzKbasnI3I16U9aGzrqG6i4IMEtse5FVlMiyCm2BqmCsIY5LkcCOKuKfXTekkj
9Iu+Ahjcq5QlPOSOz5XvyKE/7r4Sl4G2X460W0gJqTjuDKInlFpWToCADkzvnVl4
FugERREFy9NM8FOm6lPmRydLtlSNJaWoPDznliKuaMBNS+Xq3ABItPzBem1zbS6q
A7Ia6Y1hCmvJ1ma7aYGjzFyU8vv1yN4yjODJ0USNw6smPsVfNPBs5OVAXROE+0nW
9nusJDEEx31aKJ8RLNgk29b1/Mdk2mjnyTw61R0lak4g8hKVq8H90hrYQUGOvo9o
eA9HXp8NFQCzhY/5B2BQ3UMInmPM1/Z8/WlSfa8ZpLP4lxMGLeN0LP4WIRtPbFsy
9Sr9HGifI2jk14uspRuo0yF0AYPa/cubwXJ1AszyyjwUHied+kXyiw4/e8h/bdAs
w7bjQ0qZkPDlOSIrphzJPJWFJJtCntoGYArG7K388RRQI3WQOT7Ic00O4DBFbubR
kDUnqigBAGrDeGdOx7FPMNt8IYK+HJ7q9VI46JCSpbHXy5rhNR51pWMQFuP7h2nm
fgMDoLYYiu0y8YAm47JHGWy+QYERUqzHzZpATZ2bOkYbYyrSLJI9exMGbhkcEIy5
LeXtuTFuZ3rZgHDdWJrd3VJC2II5p+7ViRP1giUZH/FvQTMTdIo9br/QKjrCqVyy
3rgPsjOzl5TEKLR6zHlrdSFsD3S2iObIXMC3g8qqxn00Rx+g7HUEGIOakwo92pHd
6phPu1laSJYjHu09mTWHIJJmbNn6BUb5OaanlfQ1RQc7Uz/oXKze/IkxX4qj3skL
J/QRBJfO4mYidZJnTr6AGtNaVEeL+HrzslDquJ8QA60DIDQ+Miv7ahUwnOfDNPWp
/EMshxYR3Iu7Ul9jTS4qEDDh+2HHNYUJxUU9VDmiPMr8EP+X589iLQe2zNaU61cn
RDF67QwdfD5YUUiMCfx3TjzaeIHyek2aMSa9hRQB3AIDqh5KydpLYoz3hne7+Gxi
NBHPquTrZ3NaApuA8knTIfjI2ScIipVCal01kO2WLeaX+adFzMJdhlk82wIPaSCp
kfckOQJ4jx5sMB/WfugucE0Hp4uibBLoaSDpyZ2m6h4YuXjKyQr63TaChte3AD4K
94sPNZrDrrOPpGkWJOMBdgWgYZqb7n4ryL+GCAqO+pcWyXhzRqwF9ljw4mqyG73j
WPGY8eHV6cR7y6+mnr8kT+Jb7DbUeF5nvsOV+3/ouPH5sh7JXtfk8XFklPE6RFFd
nM3UAHUFAzYj+rdZCxTW8OZgRs5IAy2/TO8N1dSSo3l2erMTywxx/BwH6KpL5bB8
HdThZn2FZVVTm+fFnH4owqM+cJj+/xvz1I3oDJcdvsCvhRBAKTGc1gA90KDpw1TM
PVX2pGRnBZiEBuvJc/tFXEkqkAyuWN/qYhIjjQb9QaWmPf65KbtrC7e4zp/rNJAE
qJ59oAn/dMyTJ58bPFtzeU2Box8j3LkusomT6qIBX08YbWJ4kRaLNWrkHWioVXtA
insocaD0CPbrSRrnGZH+m84S0XhY1JhfhNp4A2nPs4bMfI4ZLj6cIlclNuD4+KL/
J1SFoYDhDq3ZlaEObaUwIww9o5zEoT/dZMnd1Z1QZEgWUh4jS8z67XdA/MsY98T2
6Rxohid0SmflQmCEO7yeOsrJm4xeG9jan3ItB2RVppIJOz8nas/TOhyXQabZkaHC
IYUkSdr1C+A4upVeRDBa4dpEyuTN1HymiDpJrjdwXf6VIaAVtkX6OrCMQbm4p8+r
fr8gD/c4f0wVOURHfNvnT3azFxLjEa6v+Q8wlOPLSFska8BiH3pqc3M0eXqOUxdK
+bqQF+4udSoPQcHM9n2KQs5oO9lDM+LwFQDE+/9P4ZJkSTVGVvTagGSovBJG1fDg
RFWb9U5pJV/qWvNbTJ9cmPGgBMWsvtEzCCMwz0L8q5Lw+bERqkQbehCcp7YPLjxV
dOffotfNIuttcsCQ0JsebdqGhH3hFeKIki3tE4IB1JlN1vnziAfbMm71kwdStaWI
C4JVHZKWnhffFuNc2ddSNflTuJLvyoPikXelntfyZj93/t9zgkSTtFM/li7HNsap
Krkxdq/6fdm9B9LmSoD5yfNb4s60MHsDJID/9wqz55g2RQDyrvjTMQDaXPcy4Exm
vKDytazpP0gGeXp+nggyrlg2AJfuWxb4Yq55UiVNx/gVbUifHzx/5w1BIKScPQCI
86JBPLMZgZ2lQfHi1vdSAiLrs16WQ4Ce5cHwN/S6Tp60qLDoqPoZTXTk6VbgfVYe
EOz5gP4puyTrLrKfG3fhm6TazyVkr2Z7ZvcUUy+gEezjBKxqphngntC/IHfNYz12
1am8ZrcbncFCZw6WaNkASftZhZg5ZewTQAFvi8duH5YrRA2gqPrcItIlz1TgbJk5
SxO1nffULWOCHmXwKgSOHnAcTCJnMYeN3+MJmGB3EYTvcPi5IcCXcdetVDD0I1DS
u9KZrdO+IoKZlpNsRcTEh9RE1EsJ2u1A11gCPoFpHhdokQrOiigkpYbe9jpeWMOS
vtJT534d4qhU/Nfd7LMrXzEsBw4PZI6KblE/85xhAnGKtvBvJ84ysYfuH8jpc0mH
Z12Johgi6tso7KAd5PFEw73wZ5ZpH6A1Su2n21AZtlqzN2mzw8iKEmySIR6eDnoD
+pk6FoSPbYqTD8aB0T0D/8Ra8bd2zTH8Jlei06t3FAi6D7qu4D1XtMc/9kgiEJr4
M4V2JjkZHyoSA3kuaQ/GQ3PVoCmN0uh1Ph7fLI5afAZKkqfvhi/tn5NledY16RcB
TIeCyiX/lL+/blXKZVt0cImSv0UPgTqdfFdEwKW/sw/Di2k+D0ZY/ye3AFmjN/ya
A86UcFrI6q9EXVA9feHhkJSzodFKvjmNir5FdTvselGCFAUUcF11Tc1QXPl+3RaH
shYr2FVwdMJlWTGiiRShZ74yAbO2Jczmfx4E4oSQHpzWd8yiN/5z98ZkFX8xB2pS
XQy9W80V+RaWvhYlvfkiqmFHmFTE7YvJFiHQq1kdMrIY7sYhP7iJ8o/BMAh1Rbnf
/rdtYqZYyTViTevFBE9Takw4XA8eYGnVJonM/mGkJNVW7K2mW8jn3pzWpOsgBjT3
khPp5rdJcrCWhWEbnPYUDzPlddBB3N4m+Lvm+yGNPz5N3aCy8hnSajYHW4iVPNBl
bSsq/5BG/nQFBV09RknfDL1KYM+zBG+fa+/NsGFCH+jIoP1Ouu79JZ4xYutiM5Jv
Of88Vkg3dquLJOwWXwuDdFUgHDJs192SfGPWGRXhsN4jLKClNE7o8qn4r11xS4a1
jdhO9a7Yv07yiMzvE9OU8LAUh+DuOn9n4+N8dWZbyB3JEgmka+1zZz9hnm1FO2P8
X9R4Gp8s17HebTS24VQxDuS0OrXWf0X9D68FFOs6cf2RZ0SHFWyW3yN2YV2TNsTF
muie0lc1O6xTjCI/IC2N9rBjNgPUjfnv5589zRHWVkVFMxC6bZ50zS+x1Bhqxudc
UKKOu9BfuDKdfMpLIyhEhbS3solTEPdm6c8iWOSHt+1XjKpCb7cdFOMKH/31h621
10Bd+Fni+FW5bbVS23prYgTwh3BhZIFnoXfMGY1Obg3Vi3nczoHCDqQpnqCTpN8l
SLhiBG7rMlCqku4/UdKoQBiz/SxDCyhhTJpSpb5+kXpUINLwCiXYGungK43hwuU2
HuVf0d84d8C3LoXhagfMKvbJanEj7bXzOGBLME6z2xIf90U2G72Dy+lPMaQJjCeh
oRO2aOhZLt11oUmsJLELXAnSPM2gi6KUlkSX71BbBRSpAC0b8nhgqCR0ixfTAUWO
DfMfErKD6X0SIlu2gOgVAY8ko+JK+GYctpX226gwN1LvmlPbfUy02c+mxwNK0iTp
5dTPrscUHOYJDlQ3oBAXqswDBXAQFLld0ueAY/EeYp9CTTapuuoBhurwRQ5vmbDY
QSz8YPzGzWIb4zcq+aeJY20y5QU6n1foLgogTNmWAsZnYhEFF56cPt3/DtvHjNlw
tgfecwbniBKsMBi17ElmgvPqrFilM0KznFRyt5p6Pp+Z6SPg7TlqeUCMcP3Uiot4
8Zast2hXizBMr+2E3Rt5f0TuqRKg/zKr9lJVXmEkMSUk6/FdVOdkgdCGOh9YFJ1f
63mDDdZ42B+LIUL2EIj2e3RpPQWsRvMT4KIvrVOeP0Ro0B5YVqTpffjdHldSpJ4r
STrd3+ds6LfOnJruqoDftI/4JEZfKVrlL2W+QeVS52uoXUAQhiY2fjdCcGkOdyAW
W82seCELwy1kI4xASNF/GZmB5w2JuT5Jfvw5iJuogsgq2trjvtb+3r8nixFGGQ2h
2eqo3FOlEyYGBIUCAY5eBamgNwgkVTxjRTwRzEq0XsTts9CorIuchh2+Rh9KSxnY
mTwg2e/kkr74SBSuDbaycx2v7onrJ9k2OGzLe9WkjmhPL5SGy1wcl1gdm/l0bSG6
KtNaontlr9j2Zq63KapNJU639QNYXgm8n9Dv/QI7AgSkP1z5r4tbM+GoSQ8w8U+o
n0uupjEMUueXBPaPSjGwVuGMcSabF9A+Ranyl04uDz4Y2GmRMCLVQWN4srmRgdcB
NgU5Xbic9K8X9oMB/AaMYkewEzyS2bWsF3UhsZmjxJi4fa8btXv057wUVTlUuyjM
lz+Qz2jFt3ERcOuB3HZQhCA5Vsz9ruAzjgcPadlHy8q6acQCN/B0IwDzAbHy4Kud
Clicuf7w1+5/tFi/fPZKUBOgR6XDaeR7rRLGO3rXDGs+xwbB8uFgo1fRqokU3a8J
a288DJsU7MfWrLOeMeeO6KTQFf0ZXEw326zIf+6e9f56GCQiLm+0MUzqiUisPJvj
TJ5JsIwgmL3HRuLPHgvMajUpgjt9MfPc/g56oRN6AspimeV+i/D1qyBOJGJp0/kN
JY2VMqwTiUkYjBVlHhLp6JONx/aSlRnfMNnD4O8D5JXnVYrOGxSug17wgHqGTYOv
VwXRMJ4BQFGk6sZQuVaDQ2xkZhYG0xNDViaa8h30vTtpVZbcnxGp76smDW9HWkgu
TB1yotAUhZCL171HaM1pleoUKf5X1igWd51bFt+qPieEoVKaifQsNQ2ByoMoK2o/
Cxd5So8Bcfum+eSyY4N4NhBJTWDeyuK2XSeg5ylbB+bSXuEpeSrC2Zys0uAQEsCb
ZE+Vlhd3kA+7l6Hhdr2RDBo1EuItVHLfzDF9/MG8zR5qpuNLpQN2K737arQeLarf
0stm9r+MIVY5gKMxWrwkzxCvQUH7YTK4cKgam9vBTTA2+e981l7guMjFyS7r9/hw
Ozeppd6Gmnaf1pEgZLW/lyy5eL/gbuLlxzdWMN+oqjpHaT5GCFRCkz4uPKl5z+cM
+oNXNFn474P++QDdmUxJE2aonp/OogIDSHgaI/PHSqhoSTGsjuLXmkTzqofXeFwz
efTN8KSkOHo9Y7hqunhmN74RUoy3IGj70i/7fIQSDlw61n6oYVXW1gMVACCU5WpA
Vh2BN0s47Thk8b09mTLH2QqdUk7qIeiKEUVFqp74fsEWbHtn92H42Aw3nmtHsByn
TJKnjfmmC2qgM40DQcDllsGFT+f0pvB6Tbjmlg3P0bvHhS6C2ZVp4LFLXoOqpPRU
pjO67RinbV/X7bFbWuGKuPXv6Mmm0tNFbly9DMPBXeOxVprspF9zpQuLQpnYckuV
Zmh+7DwzFUC2vh82CnH5Auhp1942Moywg8Zh/6ogHiHxsCNTfUJKmdm7xlpqbHiB
390NWUDR79sEy0QLIEKvPTR6VtTYhw/tsqwSg35JIsotZ85aVek+u430KJqrdBur
GrLd5/mmfeIA+Gbj++yVlvDZf5Yi+8hOL+10VlcEvE/2wcjzh7rwbpf0nR7wVbxF
k2HCJyMADPnhQFZ4Btf92qy0Jbcx2PidMRLx11aXryzjar1PnTyAowVpszlRkpKw
Zzbg3A+BOCDsWP+a8WuCo1Urm3uGWqiZToVGIIbAqFHAUbfCmTkSVno4Fs9JHVG3
b5Zew5OlJnyyj0bJP3f5sn3wI+wI2KSs9GMO0gATrErCpiyIRONWnN6revCmNfFI
RhSqlvXXlpVB6kQtoHR1/2kxvCxu1W0/POMAVHR7YcOwthtCG6A7Yb+DIP019rOA
LIaZtKXmIbMgwpEFxH6xlpMj+tHitkJuFWFXSHNZx6Cn1G8OEtnzctt3cZjYiu5J
dJS4wIrzt7loZGuzuTP3lXzbz6sstNhKJR2Fe2pEsYC+JX9HIsTOKwGHgOs/yoEq
0+p3PSgKyxvTP6K8Ez9xzNAQwTa5uyduyEdKLURps+nm1tO8bhxwnftAKG3WnsNR
hmQqlZ0Ndu8VlrKoQWvKUwaP8ijGqWPRgBzEchNVc8E2TfejOnD7+6v13/A7q6ZC
nGn49cuL192xLfXL7JPNHggGzp6BDqfMcEq9YqXKr+u7hISw2BllyDT7f0tksjE3
AZ1w4M9wjUj9g3yCArcYKmPNX9xsqUZIWNjjT69CxUw+TW3qQHiGT9p8Mj02zyc/
xSYY1HTtWKdF3itZKCOVbHG2ZYq8Z5NHxRhb+FDwjmGpaBacX3aGjbgfqbKX2qPV
AtLlApIyR2bycAO5qctRopoYuzURTmcuX3CQNJ2fYkAxr9eE1klzVd+iRdtUfDdH
y1/PQy3Vjsx8T26iq2ch5qpMke2/Bp3QflYRAlCBETuR7HQFFUanO811W4YvpFfT
u+yU6WiFcT3eJciW3jyID3YwTt4RSgWWbalWI9rM0CWWCQnTjrZCYVn3hAXExKyR
8CiEgeBmiha+sUt9VYhYKmi1ucFISx0XPfstXy5avT/HasqbYp5LCPYjCrO3rHRG
TWNFhHt5lFf7Iud16hP1+DBHipF9SbaSONWFpqsU3spaoFcSDZnWJLeB9yxCvcxB
Aje1wLJi3T3MbF+FE4Jj/R2YEalHf70YwexhX4WoVgF+VTtuJ+wGICxGUBzju7bf
Kllb41Lhl5zT/K7jMProwy+lPBac/lnRK6HO8q2YXbDa2QC//MK14brGvWzohnYJ
lUEwMNypQCXuQEc5hVHIlrxNF0aLjJ1jddnkhvlcyKcze822Rbv2gnu2kRPeRlKy
Vjopx+KrZ8kt10jaq1CQIUnHm6m7XNPmwse+2FRgerG2os641Z0t7tYx8yZWM7JR
ZbM+Mbr+uN+hjuhEcxi345fFGeUAKvRVgmI/Fs5aOQSj14HCUkFRAAzOsBxtTJjh
eXjhffP4iEIQ1PJylhKUV70679+n2/PvXAsg9eggHgQz26KTyql5NX3i3fQvI3FC
9JeKYncXAZf3LK/8WUoV3IaRijs9gspVXUmH9usBCcQgBPSLVSGT5afup+vsgOCX
mxjkeNwvhZ4+O8COb6knwKrkwt6jHeMme9F/Ti4LeLt/QQsCHBhMW0ky1j+0ere7
VVFFqTNMDqDwC5T//Q/mWjM6Wti11FXLyztILvFU6scn0KMEgBzy2b3F0J8WLXSr
+qxDPjkEtmh43j69WphX6YU+PGQ4+NBvImr05CY9byA1x489GIO+FaF2GDpcYnmT
ylRg+x/VYGJn8Ou2ri0jMDqEM3uzb1DkWVoagBHzpMu3rriXcLszxn3bKX2sQmAk
LPOl1Ul6fmcct2p1hBsDUrJ8M5YZ/JOzMYFiR5WeiZuWsP4zgLqz8M3ZDTm295P6
9wZqNXCO7qY9UpLxaaKagCGP2sXVYHs4CmXHYz3gjJDr0asHoORHgcZqcHlOsoHu
NWjViKNC/osDlCVDpRMs2AHtvEfAa8gcDt3STJ5B7TgouKi73ESTOeoaDU/KHlsm
FJEAOsYkJZgamAZhuRUOfaEtMYdn6bcGMV5FszoRybHPFaJX5XLm0UraIY4tNwsV
XNx/PRedMHtA3ax6VR8OjtBGo1v+uHZnTreYP2uBMsD+ZAJvus4Rd9NTxurKO8y3
jB9uDlYMwAU+apUubUB5Y6ijdyqG5yvkGI1V0ZToRCOlaTBrnJwp3qL4meNSYWyF
etycSNWEjsZn0tkV7z5foZhZAGIvTOVFHveWK2HmKR4WmwPKC2XVVWP5jDRvW+Iw
VQYJRpgpuBrE2wZg8F/STQPUmj31qMqF/DosX97kdHKQgrBMLhyJCdTp/ig/F8sJ
NPspxz2QXyloMNbfaoXpsRgv9hOWwc0RnAjBkuKa2BHa63w2xFI+4xOwz2y/YZuz
5f4p7vCg4rkyYCU60Or39l2rnu5UbAntZNqnlTc/dzEg64kntngbjDFnUqrU6RJk
Nd4Lnkazwt/KDGJpqngAdXJCrzOIr39h3hg4MbNoJTdTSkLUNVqrK6TGsUPiQtie
dTiF6OeR/TfVz4dNnLtb9m7FlSkTzaotRiBni7BwjE4CztBRtz7Cxnc0U/BGQtiT
s7s9c4dfqH8VFM/RT4y4WpCcYIN9WYqJMZ2usSCtnzITTNnR2THBCFS9GhuCvfzK
LPkdHZtBg8C4ct6f3QWaoAFWM05656F2HHQV+JHGclIVEWZk72QbtBR1hj+sJp0C
fdVU3vrHQ1571/3biWNjL1NEHT7yiMa7+g6mEl0kwU8YCKAAZePSW1pP/ZAe2UFM
YVlYk4gJAaHZ7H90zBCGsRKUL718Re5dDX1wI16SEl7bvr6cgWoXHJmxp74xjFH6
rngT5iX6FbsuXjY5bxcEgy+6MUjH8XpICyl8bU90yTFKtVOxJwYIgMHn7hB6Jf2o
cds3j3SqAIU6l+FSKjhf+3cymE/3K8FBPMdjMxvgjlKup8ADgs+YNCDXIlpQQCyh
AkfhsKPu9gxyyRQR8C2e9jId7r44UqYj1wsyR+LPuSAiv53qfeoioZMeyl7NIpe4
oAJMMI8tCddkT3iNI70z2l5RkvNd2jxGwzkwl1KrN9tEmgMdOmJFHHJZlI+94z+c
+7JtFCfm+gLpMblD8cnFw84Nb4n2wqHGJsJs6IvTVx3VFPsjcgMYF3VoMJ6uBMEg
vpaes/IJm9L+3Ug1sX+Fc3Vh/SFlOoYpqwJim3cC7y8p/UgsDlRE3X3MJjZaDX8q
xfiEaFVKG2qxNGeqs64gP8cynfHta3DbjiTRFnDo9Es7+bqx9BCdHNaMZSSp+bWH
JOfCIDwZWOk2qEOlfuXH9luI1jfW3EXk/wtXtzNTcV9A3FQeCgQvmnRj5TTlvylG
4RJLeQbrpZWXOTuuX7dxoGMHMh2Vn83Oj9vsU/ErD2ncFaTPR+D/djiYHcCEMmd9
vBlbWT0zQ7LSn334cX1j/2jj8Np6At3F2X6317HCqX3HUKoYKhnR5bp6gy0LEvQE
6pOvoSACisDUrWb/PHmGR6Xae7AP4jaXFW3bvTrscWwu2rTOlrm6dpY+kCUUXYs8
uRylT4qqYaXGjc8UYALHv8FcmcB6Wqi3d9+Y3D6lr59r2H6S/vRDEBAzWIKgNETd
MRL5KoJVNo+hsi0TcRI6NdsfaO3ZuKlLUhsWJDumfcrqeIEC1q7Y/ugEiHFM1+10
yviLbop4tUe+IsI6aK+u0mkY2AxbizMB7BTxTBeA+JX36scztf6obJ+KUQNptxIv
/B7/d/DhsZSqXBDzAdL6+BNupI4uZsHPdpSj9c+4kf8n9p626NzzzDn1ck7NuRA9
wCxYIUqUIwSfD6oeHnAsJ0V2NdFHEN7dQIGo4rZC9aNfHBbjC2EMkroq5X3r6UWy
I/xuKv4JWB9U6nsnPSILJhF9FPZ70v845NL3Ir/Se/PHxUajFaizadfripR56e3C
KgjWY5eXzfh8514I0z+dATs4IaH/x3q2BhXysmsgo7BPqkLpaKEzVNlPwRTjOZ6z
M8iRn++nTToyIYwxr7UgJjgZxO47p46cr970a/kASB7MNP4CTRiQPknVu1GYbGEV
sj6vzf7itpvmov9y7+sJQoGGsMdBoNzsSk60A8yq1PL3aeqmgkcueyu6n0Pfxjzy
ZfKILIT43XiUmWkPgBc7+ZZuaTNbV8SNF7zNO+Ny+uPu8GJnRC/HzcFeZwPrZtZW
z7/0x9tks7Fe5BKEZfIdCEf7NXFh1g3ltqsWJZDzsX+NHJujM2WbP0SEUdR8aXMb
/Si4UtsykfEpKSowGXr/6mBxnELv6+TPmCQxTEX0WHYz3i50qtnavtmSxOroFUDu
mtg4H3ZdfT6GoO6X32V3lT62HGGdZsMeKyMf73DfRLA8Idc7w30I5qXNbsTdvsYa
/NzXGrOmvJokNHkz3xWtkYqdtem0fwvyxpt9Y2mCWk2oilPAVvm4xJmNTlIKmnWf
BfH189ZWFoVsYRjkZpQv/swyZJx9t5171w1yVXHWM6k2j70ZqPn59EwBaGMe6uMa
1K3g8fyajEovVEJ6hGK3aX4US6iA252sT0WjWcVZEwTfHeIY1/otPJd63HW0qkeK
ozZeRR5wBaUE7MVrNNFlEjnL6ABUf/t/vLW31srbuMy3BU6zJH0C65buutZF2eKE
T0avMTB2Sx87hi8zmsiQ/MBjMkdcJe+ROJl1qQ/CwICwrNQXnHMMbjU8VeXkpQRV
lwd1tTvIteDzINjCdCtpskVPamGp4atek9GpDfeO4HVqAVOCFBd5dAMmUz4BlBqp
/pF40P8DHA04EqvgGoM+4h9m4haL3aXkupenlJHR9TbIvH6dBGl7EzDRTVMOOg10
piQfj+Vek9E/MoI2rMt/bODizZedvAW+mcfctPNnOxxDDcXfNW45T7tXrRqfUjVR
G4GDA4OV0rOCu+Nq2JZ7afWIBK1JXSpp0EWLTo3LeIytGVSVFN7m7AcWi9Glp2Tj
I+Cv+O3y3uLaJOUp9xum8jpkKH0LfgEqjQ40wSuJfjXSBrj/o66xoSax9t7JSW1n
NvRF1SNxrj/HdNwHw3T4S2+5bi5o1dADVH89c6pEyu01nCMv3tVhGP502rRBkbs9
3lA0U3CIclE7PzPwGPHsChXtHpmCRXAn1tx4obYtIgiiKdFc4lbU0NDVvrHNrwnF
IbqJnSYA5C/D5zzXnLO6Y85QN2w4VGmRrpQ2kwZaMARldM+IiaUpXlGIY4G1kNuR
dqShFIj+bPAcniKFC9W5bhFQEPPUwDOQa46899OzVq9NsK/CuPdW4O/hUGOI1nSX
zepq4ZdnB39yslfX9Z1xqujfXVmA3plVylMjXCCiKAsdu3fLRfhE3EDDF6LqDA8k
dJ1hznQc4BflVJjyjqQ/oual+fODDBkok4L7VdT6EbWbQpiafL9UPrU8lEiQ/j72
RiDzShaCS2YZ19LlZc/ozJ0aiEDwp4Xnq4A58nwj+fluCLbrBn77C/LFu0c2SOZe
+OtuqgD+PaD4HWJ7LjeS25upi8GcOTHjy1baaezgOmTMgeohhcq7gOghYL2xvuvZ
u5+zUHwoOMiH0zM01YLC4938gpl/RJCpQxxCu0Rpk53MMR9Am2LItMLOPY52ceO7
OmyVS/2wX1MhOZKxdqBTVVIVDHpIfrwFFzut6HNoLzjWwbTa+bZl1jEnGMU4PHi0
4Y13Aix/H4YBgcO8X8DWNVZAkN+gQmRUZJlffZyLxoHHoC+OHM6iV53wKoR0t9x8
Chh6Uj5Cc+OYl3Sohy9aRWDWclSljONumbakhJboNYowNKfQAQJIbFjHN9E+zAHG
JYU20v6N5rIV54d3psxqnME0ai+lb9WUky6yYpwMZOwY0otCiiJZFImSA/w6YKN8
Nofa1drzn2yjQD0zkSmHWqhOqPQz8kyXaxzYcTQtcqss3vEwt9pNuwkG/DCJ0Kg6
0JKoZBQxY1NKk6y+4wbDdMuXOwkfycXWSA/5MeSx7tIXIXIORJZmEBH8umRt+PNl
XHwlgvd4+uSTFBvK9KIeJCxj52cyoHB219LUdhZQCfDvkjx/pw4rPOMyQEgiFbbA
XvJLiCmMYfi4nGAuU7K25dofXA0Iv/+jkF7Z3lxecZNuMorE31FHVS5gajkj09lV
D3y1abmi59d5zgaA1bUKqeGq+nxYf6t6SHD1pH4bq7pAL6FsaYtCjbxrOAH/pY48
fIbG8oaDPQz5C7mxqPPCpYGjr7Mb31PNMbARCw+qfOWiilDwJautIyVSXoKwmZsD
jNZIQou7Db+Xnei3b/4j+3uliThK6zSclo13jQCmpdEMffhq80bIqseFNNoMW4Re
dIqgoCujj91eFkdbYfSpHPtjbNagvU8hCjLcweEMKeyZovyGGGzftgRrRFb7kWX+
VBoxMKr/qYtAgBHcQqN9VWkRd5Kcv8pkXSA6JRGYPpDMlfQ+0h1T566slRCpNMDr
2vvbOGu1RQWT6R8CQPXTC73PsfUAuyRN6v2LFKMSyEv8xBWko8+qyUr8hHyF+auR
Rm4dmSv/E2VV8AQdmFdVhUKMSWGC5Zvf2WhaqvUfjv2NSsich+4VksfZdxqsyXaL
AW4I6HlfS6RbgFAbzRU1aMx8mz3ldQz/fGJqq5l/gsK891+AgI0QYxtqlgBLu+yn
tHxvoRBGXZCp9X+r+OG4w9XfhoHI79ujpxHEP1/cK+81AQb65h9d+KW84C6QHmYX
8FTFtjrDUNAEM8TywdjCt36zw9QBT0Uwj+3E3y7BcyXoOJBXCGiHLMQMjSYTtJVX
JawZ3/wy6jqgF/Y4Bdr2USczMlDQoWA6sOiOUR1BgdOmxWVBUdrPBt4pygoFKSHE
by6NBbifkPFBIaxKfeqIQFraPMpVoFLb/YpgdLlGwjQyGoQl/xh9LqcJvefVa2e/
1gcU0TYPeKyDCQcLsgC0bZ6WGlXTGr9H1nbWODYQw0+BVPoLR1bd0dIHbC9HN6BR
374Vbg6aS4DzuL7Z3thEdoqy+9b2Uy08j8yWJ/eLzfOH4Q5uAdxVzHXRO4CzxRpE
WWWBMN+E48VTeB99y5JlBP3RsqY/t98TTg5DEEE4S9Gb3qKFj+vy7KBhxEOfO3R7
G7rWVHMsKyvbMV/RkzKQUvD5sXJ7qmTigbcTZhTqozz6iycFsuaz3Tb/iqlEM/Bo
KbrOoRsazrz+C7qxAcWg4GWlesdr7yZKlbaq4L651QqK9bJOXwwo3fFe/FIXzI1A
Px+C2Q4U5SNZbCm5OXY3vnP+exu44rpiPOIxp5UvfPu9VRcIMDUoofzsY09VyIvv
xYeOq899BaFSD5sPMK3/sbnbdUhlQiH17xxiZuHQzvqh1kebIgviMatrqDni4ikc
/o/mtz+4IjJQTXag3jtfWDE4Eu8KWEcbFqyQgTO1cWHKfxdXxqSIBxGbzBAvG1pU
sWkyRU7zZ16m5EyMbp6lCVbQRyzaVl1kz0Sz6iAoJ2VVnvQFwNrI1sGA2BfUpgS1
3T8co7ASNOsTdIBSYDUHMQkfYNhc87MQmiY1UBnhUYRbnzdGGUANUxysUII4avN4
i5kOiN0QAHrYhzZbIaScROWjoTtk0z9xpdBBM5yYvONCpelKJ/yRI7Cn3RgV1nIh
8EB2tDA/dpXvB/pzTlq/nDZ5Z7wuWq/We2WbA7D3mc6zrZMUeEOGUYy0bnI+NTpF
xSE8X/FRGXj/Mc08gXR7MDwR+z/EvSY/QPBiD4HJpDnSooMZbK3GRWgfPeAM3UzQ
znPxmPoYCYMMI/67Zcxwe8W8v2vUXJwZ55KUB5q7+cPoyk7wvUMzNljNhuYXYIMA
qtwX6m+ihA+hp3TCXpead323TtDUkDZfPdguDAXFydobR3lDPIibGZWb97C1CFnm
Y8o9E7W24/4zkORmQR9PCfTwMpPNMCygwjF3O8zUXaXNGlfYJ/1ZbkXyNLBEvdJu
TiffzUq6I4iFNyd6MYyWc6sgsP053az4hU8UUBacKz22HNeMSurr27gBsi23SQqq
9h+ITm1qYP48ZNGMVoVZbHG87jEeXAzsB0KeC27Tb31wmG7dv1sCR8N4gNgFZYbl
8dNcKRjCG5e966z7QfOsJsx8mKnaBBShde4Bv8PG11+RnkYNgBtUoJHAG45Kh46b
NlHZgFUijUtgZHrXnbyTYlwVOJRgPGDdTspVL97y1CpWNorEFbULRilQCQRIDc2u
2SsMtwWqIyemGJGQ1spQsYLlyzmV0xbU0NgJ+dJw28003JSnQp0ao6Ac61ONGZ5W
W/HrZgre6LhL6zvJkCnuyBHWoz+j02jTLy9p535JQ8K54vgvtfnyQ+fUMifxvZv3
PLPqr8d4szdd0Yd/ucQWeW6LUGmDnjEN21eFAg+4psm7Erx0Je8DdRKjdwxrcOWD
/fPiEkvQRwCFg8IWVioA00dmxD/Yrd3aIoI6D3zzRC2C0TKMlj/R0E62sZ42PeKW
yyce8woNsLyLLA225OTjvQmru+5MdN6yIE2SF46q0PWmWBTgwe4zZdbZC2TEA2rL
/97j4JaEP9cU4g/6CgOTt7yGuYDF16dGq8CSrDZqp65vnYMYquOiBvoo7WrOSlCb
QKmSl9YpFGMq4b8tgH2c/2mSfQkt3hVqo3V1qMkrx9/qdeYUX+6/EbNzWvD8L8c8
tEhBdf5C2mAahCryiG8zvVviJ+0K/KEL8z9ggphLDwrVYLruRtwDYD5E+Rs/Ernt
L9OXiVLXPOQ4DXEHxZeLbY/zGM01LthcgJhAJzaLdxdwtDYDkNYotXmKGo2k9j3a
R7YfP47COrGvXzkjbgihWOgb/V5wElJVPsF886bnnY6yg8oFmOj3WLZcNhCfRU0x
V3lj60y9BDHH91Gj40GAIgnHvF7miBmsJa5E2nZCBxTJ3Fiad9Ko0sot3Cbf+Lct
DDk0aC+ff1h5M7MKEIAE/pdXVnJnmAPcSAwMLzN9fH93RXUzCHkdGQnBUqoV88CG
cU8ki29htR5/FULMeoF3AzfA3ZqWTn5XwMA7Wb0fdZ2cZsYmM7JgxKzn++vLITX+
SNLz/BVnXNEp1ExX5zICb5UPuwH5S5pL26Mbom4uddySG3f3lUAk196TFZBAlykV
VBByWbs/H3GQsKvn01LaQgCqNK8vOwLvWK1PG1INST+rtgvHW6joMh2BSeA3s8ap
BumSGZ4pjfdK7oOWHtBqAgX3MB+p9BlUq0QjKBDvUD7/Lh4SPom8uAm0aL/TFB1m
zJTUcY13ZuXZnqoIWlqaW8oVTerek5FiPIlVMyub1LZIyTi92TRffOnISW5sF4b5
KHXDlsYNJPnM9QoItiwAD+hhv3mqQbZuKLfFOwPN5edM9QJzhToxtTw5WP432sUF
j+Ks8NrmKLLP2wpMni0B/pQ5lqZ/UnCWlOSt6wuS+n91pOoGwMB03us8gRTJi3eu
R/4/8tR10kIFkSmiW73POEKi3UmR/Ecd81EKwftI3rtpuX2RT/9SHVvgq7MeeCzQ
KXzTffJSTY7197RiXlsLH5fKoEZsEEvSbGUoJp/h2OpMH36wXoCROZYqGmQoFF8z
limeMRXOwCuUB1Chte/Hz8G4fTUaKMS+rldPZ1huX+UgvJaXo540LGe9rRaTwUT5
jCqjr1HJNaMVMHbqqgN6eoMquZL/j/RB30sfh9Xe0zqhLBNucvN4Vq4StY38hpg+
mwuvRQrucpy7dAcVTqS1hQsBmNypsinmirH5odXUkh2tf6nizVjZ67xTV+kpihsg
xzlV2HHdyLC5a+ARLZZZuVBpDTc8L6ClREHido6qm1KjK9uqNoITzsmUBP/6+wgE
dBhJCgHdv3AbPl5TpPcmvNHjEiwqTWV6WEEWNjDpRLpIPozlol3R7SONbqAcF208
pjYY0m95GFGaDTIZLQJIBigGhw2wozfYWQLEXdwTHZDhsiIUfjAaokS1Y5cKY993
Bgw/Z9pWTFaPnYHCi4zur2q1WgYQyEWGeyiwiFbTByocos8DcbXmyGvJxRXaUHc8
m3GxfnzTvx53cyWgF9WUd7FbBkkkIe+vk499hjSayHkpK7jZlYiFmziNetFjLe0P
z8gvI7dorLveiuQpgi8/SATEnQnLSTLccRKx/cBskCIVNUqLFLf22Bq+58NPXr+Y
R3tntBMmfo2FQSuT9XNwGhhBqibTUeh9AUe84ABBQRnZBydrJZvmA/hXwCtndDmc
YuYYrHeMBLRZH6OmAQ12SF+lInasxycrVLxQ6pLwY4XbWa3P3JrpOQKvNh6ztRNp
YZYeu4C+NxPss5DQAS0eqIkJx3Jc/gbb0LT1m3nG91KQyah679xp17D5NFFtqonY
FM6ND9iVX/E1nyS8t+bt63i8pxhVf+2j508WW8xOqVQn4ce8i+U6jvtU547BUck8
2hcrPZ8xSjbVR4L1/SYol9/hvtncuEODNOLx7BM87U9TbByCkXxvkpg2IJ5HvCje
zDOGMJXwDewJA1QqYH/kWM3dm8DHlvRZf8Iq3GC3NIAexFS4JuS/9Q12dQ8U8niQ
rG40C+KNDo+9eh3WdrBMEWjaZgQ6SNobAUhJjBAn4o7JzlRm7T7Z7JhKGPXO47lt
ntfshaWmKCOn2W9RF3Bnp4JYsPrSGq0BbexsrK1wXHNt5y9U6gzQLmsHfOnivhrr
rSs9d94wR1HVg7GpTS4LVA1InE6r0ww5C9wBy9DeYRq9UvtR6pnn7yLhrEligkG3
wIh28aG793gDENC5uVIKMtxSqcYgMDYGkWKk9/3uH5CmUHgTe++KJcWJOHGTX8bd
P/mkVdYzpsIXVvBMAlGavzOgaz4COyGpODKe7TvVoNYGUf0TQIvgRRhM4iUOgEYo
TDVDRsZT7VTpkivlcoOEcFf2bOM7Ph0ajOm9Tx2Ag51lOhiD/k5BtT4bode58I4F
oxAQ99tJy1NCRqW1ErqFDMyy1XMAUV4O9PjBYOGD4y7kdFT4HGzD3XOG78+0aBgA
B/1b+2o0jFQLBXQhue+BHQnV+Xhgq5upKGsD9Ul3Rbdu0Yo+sQSh1HhIUiMTQFl0
wJ/R9rfijyH2Fk+p0E4imS8N5W3R1mOUH0sQol+sftxsG5pTSh6+qBJtTY36QQXI
wmPvbLNDT3tyEfQc7Y6C9coh2kKcZIf2SYc3pPnT52FNeOvX1iq68Pl33BDiOYWI
yLXxHQjf4QmEO0UVS+5O3SkXEQGIx74opocUN3SKh0qhJPndYqeH5026jzfRUjm7
M5L5EERweZUXxfigyOm2DH13Y8F+mrLsO8CugJ1R5rZpZap3Looj+PeZ7W38ef9N
YXcOUGLg4+RLIRjcGovocKDIsupu6jotPVH6s9Yd1KnIsyaV1mRbb4MdGcjqc53P
4QMYrLwoUmC7gSar6m1ymUBokwzoL4d7Yp134N7BnJgeC3RurmFT+69RbcxDiK4N
IJ8s6LtPJouahP2zdqxduQQlK7P1bZQzjnshX/nDkHndkXUPaU/IvQoq/hDo4X/x
kggt4Jip5zkXh8uXeC936TWyiJ13wNvNQE0qQeYYlWuCCLBugsgtnCszZs329qVH
Eqw4dxycCe110ziAAFpzzyJbxFU0fMYvTzNZhNnhiqV5seGPw/HiMfIZ8JfiJ4Vz
UOy/uRRfN6vjMFIo3wwD1QtSu/FsTyvQ8ZARqitXLxnvAibZaLl0Hl7qlXviIPCK
ExgPV3WGG9XDS3QV6VXB6rt7C9jxwmO3KCZ+qe6QpZ+fBOZC48FwMQ5B1anhAAzu
9G6kAzVRS2+aYJTQKIZ5OaQ2p+ClvEq5zeJfYtQK9L/mmSmPmKimkmETY8ZdIfQz
j/Z8u3c3Ca8oQOXMk7ZY1JYLjMC1suzMojeB4mRPUPzxhq1guG8/erp3z6RqkCQV
z+rayefW61atE+ZxBFnp7nKirPIFy/JyKoll7xLzPKayt2hj4y9AaNNKai/mhFgz
jw0arjzKTDgxRS23WWaxh63XZWWmaqhxN+rf7M2O4ybd0505ivFH713CV8D3ae3H
5mqxuiu8XK3Vqq0XAoEW05cdj5u83buZQlePdfRuoMNjlG5D41kaG/f1Bchfzyqy
qVdGhyljmFhZmN0gjKF1jZ5dEaZnQ5EEckhRIGypqSjwPX/U7oAGSxD9oWDFCWoO
nfCvLvoVCGYCW0kll7yrwT022cC4ANykKpvcnlkXXUMAC4hjz+LbkNYqi6UjnUke
Gcsloy+roup9Xfn5uyny+91HFzwM+35Q6Ihs4bHlH8hHVI5bDq6Mv2PAmPkUHj86
3cCtewdlpgnLRj6YgIXPCGUaIb+ZEtm1XfLfwDXt2kVISx93by0JjXvcfjvQuKBG
HeW+J54+eMNnm33Ue1S6vS/KVZK6+wpmu5UPgNgr1SmuEuSeBpzFvBQ7OW9oAv7L
JQ5Wm6SgyzgzgMAAaOQtrNAY+Rvyyyi/Ky63vh3xmbi+pFKcuVfDpxB3M4pAhr3+
Nlc+dqjHY5w39jCLUsOPKINWOiQafo2dmKdjw3gPiHn4foRhMM9FarTEL8ZqskaX
00HK3WOfO4rvu7H72fmpijpKWtEuSEWGgPXJKyYPyBOVyrPzFFXNhUkDp4uev0yP
4N38Nppa/LJ5YXouUrl9j4HDh0PnXR+eXYbVtLKoYy8EZZZhbBuLYMCUgd969fQ5
TlB2dz4MxGqouRKl57om5Deh5vwW/69vARdouDgoDQROB8F6EIKQrqbYTmZCIYvF
pZ85ByUPiYAveHCWe8lFNMENrKHBWhwzwJvbpf8QhyKs/MeqZAgfcf76vsOLyR88
xUTDABz6VbmlzpufBTR0F9367qcP1FR4LGgi0KVrm9nNywLa/Vy5QQ1bvqhO3Hc2
+P3epnMJuvsG7HC9hwEdqciDMavFPQppXKW3pSX6oTLRxeJwrrihxAZ9yjC2BzB/
1Mi1PSL5yOnM144NMNTWnmHWtK3hWqpAswYa6u9MCEEjms3zGQ8NY4BfdK+tGlJl
PO8FCV43zt5tjJlHXEoEiatMvZK+aHGNQzyRRuf2vXyi3aVMwauRQNUkQf+oYF/c
ZelFGa2fNkdfk2idShqKq//jjohbLIcnLYAY9KjhFE3Bwf7N5c5K0pp/TlpB0hxA
GUOZRH0VtelZeWAX734C3ZueMDmQ+mbJ6FL6FM3JDp8dXWHk1GL6rj/pMlNNk1dK
WZmpIv4hTT17GwOiXmPG3GFm+Z/aalptPmh3hyA3lFFAUk5TjC+egQWyxC+Yd4V8
egtL2PtjCH2zWD52rhCPfrxyEQdKG0QTji6ElSR3iNiv9a+M2fZHjAwEPrQHRyEI
1MOcY8sULVlFkxrRbL/Y1ZqIOIfPRFnebmRFvbs1PcEFME6oDqpBkv5bjriKbRXy
GvVgyY1N3Th5IUTc4Clv3tLw7I00VHKnqMd4MspLigAu5/ewcj15c+eEEKGqZBI+
Z3RzpNyDuqltfLcUlTSTeBVZUjYHqSQjyvvhbWMx8ljF2Y5N2dFq8eUzFpFJ4e49
LWzzvfESTvTdNWxHvw0jCX594ivtAgvkZbw1Fwz2PF+GsANCsaz2Evk3fjPiOeVD
QFEa5EMzFlEKnXPyVbEzl1ffi68WaIY9+pz4g8o5zLFFXcs96KClAQL8KdDDdYtW
8HmmCbLgzOv6L/j1b/VdJSSLDlgfCwQqPc0d/PUbbvWQ5Gil3f3bKpBHa5jD+sAJ
dg6jiRo/wjGJdZE3tv0f0COT9sYDc7I2VjWEwEsKXglJUP8I0R3/mnqbF6PDYJ3n
7JMEyhcXx7Os2Ag68BKHHkNxq9r+Z2aK5pcnu4AkG8zfSzZTAQ45MexaX2vAS1Gx
QB4OCWZZ4NlKCRuJANj0l4S/NOU1jBg7dkKr80rg2dxGmzif6bMpihFhGPg+RIO9
RclPWB/pMra3A+H4OasnT0h3dr8pJ1ZdQHD93tkkSdNNzl/DDqZQh7BLo+VOAhJV
ozepFfO6LZJwZCNiMOnjEZVdHU4wJiWxEWcQTEMvlgXEboshEex8u/4Map5fMXeU
UJqHQpGcO3Yiu39d60Mw1qtOYM4Vyjd5QRiFDcOtCq44aZ8Re/3iWPlzTkTQPns4
Tbzl9oKdNiUJIcluvHMid5f/6dScz8dg+DCB61OO/7TGwzhhZ351uD8ByOFJLAw6
3id6JHy/6RTX7JGoV9AVml0Ky613090YDyQuUYkPuac8iLHPMr4KYV9GZ8fTXCpM
vuEJKtsZ/udnc7wWoHMhOayzX1DGkJLZneTwwzbGwSbo/ZC3R1uUhpf/Xg1SSknP
plYh7eQFvqA+Kq3M+auYCD25LrFim1Fi4uudZAbMAj4MvYx/hNwJRdnKhdYbyOLi
qBm6mXRCqO+kZfpprxjdUDcbTEJjxj8Q7Rxvjvtve+NxU02mxVYE+UAwz0HP7mhJ
PJtmd1BfebdGmBH2ANo0SYQiNo5MA8pJWXZvoTc5QQhhrPcdWcdtH1aA7lwUELm/
7yrI/5c7mASlv4FB53GuCn3YQhCWEeZ22giot6H7R4ntoxT8DGzkE3vaBYXJdnYh
KFKv/q4mG70o+7UaORzT7N2XeU0QcbTxE2rHRKv/IrC2TyKg7+9XJDhZDvZsEcyn
GfB5uV71f92y04oXwMza07uAWRGgyQgx6nFeCsi0jcFjOr1k6zirjnepM60iDDFT
K3arkQ5Qw+7bbCG6aFxZEGcWyutaIdapdqDbAMdghv2puuN2wz3a0kNd5EI/3E29
p7nS0bzTOvrzQAMrky3r0MxBzM2pl5pPfEKs9KBN0UdXaBkFf6rS84fmbEeMLLjA
cpP6FVJ4FeVr/Gah0EGLnF8h7vsNWUw3sc0P7aljtAGh4wsnP71D3GTncuInR6G4
CJzp8N0H5mYIOvc5IFwdfnEQGwsob/kWrs5AfcfLT2TCjlPZwHZoergIsNtklA3z
R+nboU4tKkWO6BCPeO3bylEvPcmk43oLcT6XdaN63mhlccMXZJFfHEZmtl95WT3q
c/xdb2qvKcDTGe5c2tH9811hhPuwCfF7Fam1fFl7ftzhI7LmWPx77KKXY9y2T/Ss
/F7e7YaSpAYrWZ3xjgNoWffD06vkYwxrLJj9DpprsugP+3Q/U+SUrUBCsJGZqTGS
mHFZWDM8g8+zA8u9lk9ECoFtEzgUV/zXr4hsy4b24YtX3TXLhYsnChQrd/JuFw+5
t882F5twryhixQfJIfMbhzPo2iSoS7pDDZ9K3bN1Y5hpdfI2nqp2ysxN1CwkG8DO
ZG0bAfn3Zd8CMNwXyiz7XwtjaT2J2yJwaNjmuWVzURPsUdlTsMLz0ROmRpQT2p7j
jt/2RGJX9IaFqAbn4ZrNza04fb9pT7Br1bCP+fQoCgfLlYfyi1/J1CwGWpu/BUQ3
MtRIffpT9AepnelwWaphZcHRIeFDiyaLLReBjL6GYy0e2ojRYK4xaMHoj1/TKsKE
mjAP4Z4JTgD58dAvlpXDFUdDmGunYhwBpnWyttdgzs63Q6zXKZxm4P10IYMtZYlD
at78GuGq6v0JMsOVHQ1jDk3YE17U4CM9nYgoC8OopxXX1OMaB3uc2g4Y5Cjlry7w
Qu/zil1hnRqZ8iati0KtXT5vL/DJg3DPqO7t8jjSh5LS5nvB5pmzaAOcLz2+tDZt
xH99/jU45O/vXKHZc/vTCAHdv5idZLkOajtG7ftp+ffC6xiJB8qTVltTDdHI5Knw
97zkuNSNqSsx0zPR3vOvEcURbmdPYb7nZSxJW/nCBsTj4kxSZa1E7WskC83mSY/5
N7gmm4XgrSXUaDzQIc7SOwsE3zjaN8xaeohEIjnJFyMTfYyJelinRm7V0vx8k/iv
oFwRZsh0GavphQpqFX+l1lhdYD/Cz7ukP/dayGrLacz6NU74OJUt0aQwmoY6mQD1
0029bfV9/SooEQl1Nsu+L7xPGbjQ6iF8y5+p1oKj08/8zpkCO7T0KQhWrUMIQ10W
InT1RmYNqClKK5c87ZmCifk7m8UFI4D27mbRrp7bzyIMaPp5bfZwr9qd0B7JPIIh
roDTO+toiWtMOlaYG9xHSPN2FTcCkNMH/EOfpNNk7IoCrSm5+tJ6tJxoWITzj67h
o741wAuBYqtaI5XXcVdEOrsQpe7kWlai7STZ2WSPvroC2zAnsedDE3N4cZ3jKRce
rfxsCqeOmlYjo9trvTWIyIeASVRXPQNslmYyXV3eziGDJ7bViZRnzDNp8xbqjnmy
o6/WbzABRGOf0TSE1g4qHvGvVUM0pS6EcqjfDtBeoIfo82xCkAfH6Eob3dGWyvvh
/y6RP127QqZ2ZfIm2++01a+2OlaxOrEbOmYL9YUPZSA6i3hkDAnfbzuKXUvH0Zt4
/VDomuXlZ1Ze4RT4Hhjif1OgrOjqUWZrrFmb2IWtMPsRa0gYSRTdiJIErYkVFamB
AbNj7qLBKdv+gGJa0+2jU1ceNF72lsr1ryZ+uSyaD0qGaOPBLKMFGoUHZYorkHun
t3aPz/FqfFjC6/KvpVo3JJOTRQQal/2kEIFZswvOM0C8PFMNJlSFAP/2nbwMpnPz
atHhPkVrVJ3i1XriZPNykVMNlYTQka8bnzpd23Zsbvfk8+vN9bPF2sUTS7CphB4e
cL8TyfgZ4GIWb7cXUSOQe5bO6S2dO2m/Eec1kK45jaEFKhiHvNxmgcPQYILWamSo
EpTTtXqcKTjwshkOFf6tXjlUV08eKflZ6OT4SulprKbZlRBqxjrxYJf3TTYCZ9fv
eFjbn6x7Q+bX5vZ6e8zGuShdpJ+tCS4WlB0kixEeYGFE/t1OG3mgJd8CmZldwEK4
e29bEbI5gb7z8JbpGJVCWjRPkhyy6amcnvJGHvrcoLpOi9G7b362wBKdUc0gWEki
weypkWp3Gcdq4yIZ1azGXb9jsmX/sniqvEthcAEg6ZFvmsHzzVHlqU6V0gxdQee4
4W4Lqx6LeM09C6Hom6Pv6fPAvAq9liGV2yjAFOruy8ChZ6dabkIcFYh1zQ9JTBpN
nzQdd41tQlBTl665fGbnfewyezFQNZw7Rk4t1MTuSTLeo72NG2rb1oQ7dEgbP273
x8Eds57aX3Wq4lvLFQUeY30BRHAjXuCYo/dm0Sh2Xh6Eic89ue8qQ9QaIBY5O5c0
vcY/kskYVRiHx1fhAkYrGnEIxImywkyU2Dx02w2hk0SkWl0ktyObiFvkyxcX8LhF
fwAymRVl3w5S463tfALZB2s++Nl/stvG8jnhGAlPfy6eqUlHY5enBP617nRQXzSO
EB210dJbDH7mkMQgH4eb+6DyVFdjqAb71twQalQcsNn85Sd5V5KhodRoy4U0cm9L
18YTLiOFn0FxvGB0QKpRVmGt858lhO/fn6SEZ8+2xdlpKve6ZiJr3nA4pHKVHpcl
92Wred1EEb2W4Hx/jo/TakQWOHpjfBKtgCyYi11ovBasNyEugso/H04GvfccUJGC
HY8eEGdl1ZFf22wsxSv3ABREZvGVK9+cHb9VSVWPTyv0Mcmoujx+UIJiDIpmTgYZ
v4YKKsD2oBPjoT8eiPLpFsEa5EZhah6zjcT2IqvfAZsykbJm7c1Zs9Vfhk9J8jtm
u0Sg4EK/NRxMAAPFxH61jWrU8cEzmb5uj/bbWkLKRLH4zGCpiRmlZwkgy24t03QI
IOSziNL6AnLICaQkekqTWP3x32fNNaYDfCMYR4T9tr8ziukVeOeCFN350o3i1YsZ
4OMIwPIfNsGcjtRjIhCqb/oC56lMLcM5hc4Er52GzV18GAoO7FT0+9vlp8ICRrIr
xIQ8+6nI/+VLAD60oL3nFa7qqXjCGRV3cuEby1dHTKwOFl9tyWbrNfIr85GmsjwU
8PVS5Dn5nEQXrxqzS9zoVSXLAs4ohSLzzKBTuQ+m9tN7sleg+GsxyvdbnUTfgX7C
qNDKsC0esC9KiJCIQyRy5V3GlhA9HNKWZD4Y17ouY1tVcUDYtG62Ym6EgkeYL2Z4
M1T/H2nEWYtOz/SmzAnbi4WXnXfLLXERLPMC8iqamAyLVMe5sRl+ma9+ubk7frMB
XcLlRZxJ4lsSm78psRD9NrSGUmHgiuWnlmazoeJf0VdCxtWu49piJVAPn04AoxJK
EZE6GEYsH+EtiLsc/vu/IneGBoymxViL+dWJ89/onx0H41yJ3mnLnVg974uQ1bFu
Tui2kAAqNzCyt6bbyuDnEq0LYJgAFE0cHNW2iOyHOMyfoCMIVXDVYDs9OKwPCUUy
i9+VUquDoY9Is4Ph38wrUUdf9a/Bpdo5wz2zlSK76GTFbRKVd9XAm4gNLwHt01rt
JInFDGCo2Gqyk7gGS9dIVSKxUX+UM9Gg0hTlcj6C0+csSoJICGG+9Ok4Cvk2dxLm
yvbt2AbQoZvIsGZMjlkMj5gNQE4aDkz5HD6Ldudgzbw/5td62h8YSjiftlZUYx+v
v+xW9FZ5IyQ7k82vnWtfp+771ewvahfx+EC37HHSL0QsKATrV0hFSRQlAQpH0W2h
1ur1HeAfKDzju9CS6zfSjn/exPglxKmvZawXoEfgzMX/t0MubXB/xLsk7JPw6R7d
JOruJFxQ2DYOuJ3AdIrkJRFmn495YZHt1duvkj4d7Z8Vghn8hfgzN0/YjRijPJzU
YtbNTqM3p4H5FzK5hoscdgOr3ZIsWpZY4KPwAPwJ67VnqIeLOUZ6ijOutwlre92W
pIjUjgu96JnKHjs4hd+h8B1DA5jjKc5vZYjpOuk3YqZg8E1yO+ZQ4PPCxVLCyZfv
ZBWVQfltrRh0w9U/FPhL1aRsKlnHFMmsDf3yrp/oQpnZso5qwdG4jiZoCuRPFPUZ
kbzBz0TaJqsx3LfTipU2/PCzjMfvxX9eJpdrGcz8q7lw1uTc3CW+M9l/lNtpTAW0
NxT68NuooegMfiIEM/ixakvfuk8xN3Kppp4HmwD/QDkpXcsfy7JHyUf2rktx/ASR
Rd5KXgJfsgmk4mmt2AHoMnYxeHTHeAgklYH4N4Dait0mJeeQhLR1Rwu1c0M5jLs0
q1FArLJfkZmgglD0ULCc5qz8Z/o/OQVoPBUKaX5ltxNEMffS5Ui3FhvqEI905HqC
GJLM2CB5vAizlWUmB7PmoHxuwU5wi9FD/xw564lfSyE9UoLa0fNkKINS1gbzgzCf
++3ueF4od5AOgcqyVUYs0eLUco/x3+Svar1cTjWeJTCfv3ab86NGey+10PWbkkbP
dO7871peinY4Av+FLpIVGQhsY7POwCr1E8gbOhOCzAPumT3x00FD2VxpRt8Rhgco
gomTnvZ4P3Jt25y3//oYeztJSfabcNnNmp6IO9rf+bMIMx/hnplJlFVO8MGtKION
ARK13WW7PRR0YCuxtD+6i/UPhl6nel9lCffCHyaYEdoKuss/l/Yj7zdlmNOmeinF
g2MOXCe/+7Cg/4PP6s/YAnsqMojjy/A21nfeSiYCBEqswHx3c8Yq/t7Cve9E6iS2
5ko4252N7go++mSwnOVXtSOJOkGVgrFEHBSjCERaWeOhTxTHJJ7pdKC7P6B9fdi6
2Anoq7X+yQxhUeZ5ipce1nShvihvoT1cFKhkSE36X1HpoSVvXGcVi02NH0PXmA2V
usxcZT6UnmNekneR9LLjV13zwc7i0gc6aRxcX7wEO3aE33NSdFPzVu1X38oMfKcI
ZtLfJ6YfX7eTLJ6jCNEyTctfuT1cF7dl2OV8+6UGGdwimhsC1CjLjH5pnV7wXcX8
Y46BMuL++1O+gq6vk9aoq1Uk2g2PTfPARf71CY3/e3pL9WfO/Nb1v3J0O5PiNeXP
39MDOp3IQUkXmvY/XHjvhfOq/tibOlXEYQCpETAHSixA7/Hnb2vk95EcFBnn0ClW
h32EvK4oaTq/EMbMo8LzUPxercnw8ofD1wSfDRiqHm8zlC6ZRVDvBD6OX4476RDz
GxrN+cEvgslZlTt/MkC44W2huL4ZVRwwJDxKrxfUC3hwTMJ/jdEjICMhWdF7/QH4
2kqyd4LeMMHfPdVtOzrnMMPSff3yl8L/9xVopwRYN2H3iuXBG172g1zBXOi1JPHe
G0aC4gLY0k0ktj02cg1PF+dKkH9Za00jmEP49/esz1T9unUyz8Nnf1h0K2rqVOBL
D6DFaBkcAsolOgVwUoj/BJAfhOcXJp11B4SlCERtikibK+XNO97ZS04DxYaad7KK
cK3c2Z25KaNPeKnYQiiPOyPDIq3hlyI+2xqjl3VuuZJOnlwpOrIebkz42H5nkzNT
X33+M2OZ2B+8StDQ4sN7Zdnv0bPZ+UDpBVcWBuVS8arBiHiV1hsE+r8aQksGOnDQ
YivwVOsLDXLMxzcAXa+y4KQNb1iynh0PXUPeu6vlm4g68iMXPwE2uwa6KadtDgFv
9rShMEn1HUId4j+78eAu2x4BekFPLicYkfPJiCDxrKdGd/AWcVurZkUImJ61sSnB
xhSWNTrX/uz2pP1ELncXFpbSJaV9rnYYl40BY4NDyNJsnDwbEK4pWQSZOTikCqoz
qaDcPCtb5OM4AQ8p8IHB3eSeGR5ageJUulsoJEQQr9RTocfmsVlrwkYZHAs5iTOD
NzCd3JoW24pq4IqxogpbhNJxBNkwA8Bs/6OACt7yk+bmiEjJERjfB6SvmQJFXFof
V1Ogw5tyIZ5PH1B6m5npDy3Rvuxetlp+3N0oZ8cf4aBcZm7jo6H7pf0hHFZablXR
13WHABsJpMvH7NY4v8NHaPuvPhCHllG7Ao89dRHmziRAuMsBtabf2zPaDZCPftYt
/Ix8Hl4zu5taZLWnzOTw858mxE0eWkGB3EGXG9jvdVmEBxGRtvOxF2fsnhoICeCC
0pkQGmRHeO0ht/rrG/+CrlfhXHlpPstFqGHAMt3PcXZVFdfCfkA7VQdM85Q5TtF2
HS+HP4jV+Tm9PQUAnkY8+tmMJ5cXKpc1o2NhVIrIKp/5uIHyrh22J0PXcpmtGRcl
QDga5X0KLWRpcFjaKi3pnbTykD+GCWmhTzJpitKbcM7a2F+WSwpOULyVM2WYgbdY
nDH/boDqVmYeN9v8cIw4jPtgZvnPIl97lghO6qWGK79OfpWl7rV4KRwYbT1SQN1V
0JGCa4g6ThBzHTS20j7zlgdqCNtVpKrKgwRUCcA17FFkZlT0leLyea2BOaQ1TJps
L08istZIladaQ67SKKHnojRNfLY+NZw9lksC0KPRIt35S22v9EvwP6cDUFtgYDAd
jKdC+3IdWxyYQcu5GGs2tDrH6C5vf20j5kl/gATo83N6J9xHUq29i0mw573Bq9yd
f5ERVehbDw5HqTaeAQA5lUjOwOIBN0N5x0v075B0D0aRgRITH5vYi3Axy14iFfg8
VVBNJGcQZCm8QIIXfBBOOgzKf1OTHVpGBO3YLf3Pp+yjcNWL8Wt4Gz6ueds2QpuL
Rdacc/uuJY3Jm8WeT5IJBW4ZD4M0+95dNEAdebAkMxtU3oYvcSfxrTBecK+aFSb0
H2zeVPTv9wD4w9cv+lb55SAkEga+enBOyza7yPu3+3Xc9N4dJm5A+YGAFA37Eq+X
xFj6Eb6VQBR+D3D0qgXlwPIvxwcj/hbGpcReJMrRzb288+gpKuUZuEpZta1eFGby
UvCm/n5Yfrjx0UNMaX32QNoVFw7Tl8c4IiaNifm9E9yF8gJlnQEnUW9pRG1WOnzC
qJnxuRDVuB78zE3flDWsWGO/cczvh1U9XblktLsSKUYg/64h+X7eC43qawSPRGzg
86EZhKfqhFtZxDuZJbyyfNC6I1t6ozgTqkKMUjt/+oAX81JPizDsuw7YrGJVJn53
trDp2r23z65JkbOE7fn9ngS30p/VHljpHjFK0EQ/SQ1RA/bfvM2bPrDGShFR5yFS
xehx6hi6LWIhyLAYSudwejwKYBsrNqfUVwYpF/YPgwTs3jxjawHJcK4qZ527MzUh
KcDPdLP4Aydh8/MnDtspBrcwQhP0EkeP61hYE+40SUlXw28dbNwtJJ3PppHqiarz
QZbWXIfjm1LQSfxOP54YnCjx8nExZrT/ghS6SWfaxPUzdeDutWtZG8OFVfVCAgyz
oYfR79lqnQvfe7pnacN/FLJP+pXrdzyFrXIDeQaqQLBfQ76V/fOHv74AflCxXoPw
db6iB91nywT+nmNF1BYbamzIvkhc2v+nXX8dzabOJHLQyGba81NA7R0UVuacpQJw
lT35qYAIehr8+jC9TXrRkMeRhyRTkVq4ufOqyj5AWsRAPaU/oMF7UhAXGQhH2JGS
Vkbgu0wcS1k4Vxvc+8jVJ3ghtxgnCY7EyQd1xr2GUtkGqKlotb1bQN6CDfim8874
9XTWblcLII+CDPULGfDlcqnCsc7GBM0FIRS+z6tVhrcA31d5si1Jqp1SsZTSPAwh
Zr121xet4Gl2ugv9lSWgm9r/GbRfN662hfen8NQSV1DF2osq4Kg+o+IPJc8vhe/C
tIBgOpHLB1zqyD5fiSOvC1PkY+2u90/8t4ag44YPRl5FSuIwyUHXMSQ45O3hcT2x
qmJ1EPHiSXg68j6+47V1VLUtO4wgKAjPcBB6R4tprrTY1t8tvN4JAtINp0nUYdHE
Js0nH1wl/EkYRLBb7mCcXTOY6TV57dfeKfzrC8CTQmFoXgK7LYcMpDTY5T3KIu7T
Sfa0VRd+Wlhah/IlRiTlF6OoEMzZMUNN8ptUDrs+MbLNff7Q8MuxjFFkHZ4dQ/my
HkMV5Jl9Tn8kosIXyw/2Nr+BVUzeHexgZmIHm+e507IpKUlnZBGF+X8dksoKhJIb
ib3HJoqtPx/ZEgyzaY7It5CQY4sK1yIAHapEFVLFN5bXmn6y9nsUkd5FGtjKmsWH
xJquUrWN4qDhZCdBW99dSIU0Rro6qkRwOsobrXG3jMDXaj8+zEZuOg896wFpciaA
u0+8BxpxUnp4Tj9ocFpkYOgrj53iSdA77VNQgyjAmaSGe3GbgcYJtpznl7DsoQqO
m+7FEt8WxT3fE85u+W0HNqOqJa6FwjvDLUaOPP2oiBz7TO1heqGepG/jqu2pzukL
QzbjtPYfV6hwgGHcSaKTrpOm8wTR7dFV98+FK4NtppRpbzfzrOSKaEutWBhkmVXq
TROroP4MRvu3j+6kxF2EbxDGX5Apq49jnjAWB7tuy/0nR337lj54ctx8eLx5JHkW
QTKBX1wKitTtAVYkgagt5NFirQsq/FOuTmjVweddwsS2mgx506CbQ9pWCdhAENhP
w/J2DGTfSXLLP+equPG0Jb1nbzp3K0H7ZKhS8o/NZdAdCQl0qgLRgT6z5JkyKQeP
8ad0R4OHItlwqFVwZ5rkOWlUw+IimFMI3W5MYlqU7DMbGima6h4APEZjk0mukpNT
TILAyzsJqk0H+ehqbFFHb5ajwnNjXNQPq0fZSXKLRUXVNxjOozQps77ixnYfzlwS
2SjwNLYsakAUkF7d+FVjzWsQoEvE4N1Q+7t8Bsg1wfndZRZo28lv8OkwbRbyDwmF
bKW0o0UVgzuHatALefG3DcECQdFKpDR8X8fVymXgwUwDl/zsZaI+aIsm5SMMstYX
eDhGPyBkHNKW6l+WGKA9befAZs7zubDWBi24lL3L32tJP7aIqyF5GafzzEqX6U21
SVbRKtVcwtheVS1mx0rrp+TbpJLvn+7ZmRJ7vz/0JBp35hnIQ3TNf138qI+rZyIP
mfhRW7oJPe8PUFqS9GFrEXHmQDa0lorrpEYdrLQRQfOVC4q5IHbko3GBNXITdaYD
bRObfv6eFLjrZH6sfIFI7nDFapHRrJtQxThQw2fwJGKnE6x1J7OYQyZ8DWbWGy0k
Dqc8X66FuOPQhk08YMNvnKufJq6Lblmv3+tbn0AEnvrZYf0jvii6IOsg3KdwpJVP
1NXXwiKhSRMOM59+qu3avIIOSYNTUnLKm6ia2bdDwjTBbxW8YpnQ122AT5FXAsmB
5E4uPVQ/3EL+hcVsSlrVHA2cWFDcsTUfoDuF4vpmrz25qCEdIqDHE1EUAGHAW3Y0
jC3qayYtyq8WUpVAhoiite1JErYdRBOz19g7jIXnZbQH2ilLy/D5Y2KJ3/7bCiSR
RdPe/YFeRAUaBkVhdO8B6aFu3hE7e1A9ULHVOefIMm+RfVPE29j6C/4zfzxboIBn
vtYaJqyDGzKV1Gv+iHnKKBfp2CjPngAwt3VwUJcXkVSiZtqayC4y8rAGV7pkohxc
Sv4mvz5AIqbPR6b0AnWqm8yIPumVL1NOFkh/1oyED1L2cn9VThqLAkVa0aE3WnmU
ZqhFD7dIKN7tkptxZWPeEBTgHAx24HNPRBAthDPyeCpo5JnJSSGIw4s7GLxIiMnx
7Ml8gFsB9vWTLbKPvrGMcBnBxnaMIsmWiYrkIx0hiX+nQ78YYquPpCnP1E7ZuvIJ
2xCwnsg5rwlq3ni/0u+5ftzPedPoXX4pd5bft9h3/lcYcWR4p6KnHoqF0nY4NZs7
YB5zr42yb6AsBmsQKXYwY5i1BnLSblKyWZVX2kTlZBqz5kTdSryF5a/vgrZpB1o2
lBsiw4tXizsjuJRMDUWldFvFeW3JvwLxEoSysYElTk5sTd1sGdz/T7kGYNkHxj07
KtIWSFDgqC6u1c7CPCmWvJHqkNjhpS2LrZ77EGdlip6v/m+PfRq7AYjH2xAUfQpb
zWtAz3blIPUnusm+wKSoTQiWgZ97EM9bP7LDRrPBWwJJMa6ABTCIUVn7fok4UzhW
2we0ZGHO7lQj+YaZKC/P4AugbtKAkEK6Qbdi3hFoaePKDT9r0CczIaR4A2yUeXCC
MOczdgi8QrfcwgIlg25hANBJMWFKCPGFN0eg1aix9EBlMgypmdhiexT5nM14Rm1p
KKqq+YBzeg3mbfNhsyjPYxErRTHcDsXm4VB8HOi0mmGKjihKbxPtGG3MKBywD8i7
ZGYv7mophUtPrfcAP2tHY5yPjfAo3qulFy7I9jPtS3uK4ItTZb9cTqbX2A5c2ahu
s8u0jC5PIXDqSQFgFZERbyYl4P8gIw/VRpT/DqmtbTkC1YTmVjhkZEdXKvoJ2ohd
TrW7DUVObdUH7CqduR5ewMCXGBMMmgJ4TTp8uo1vFzZSsND8G/QKgh4+ehdeTRtJ
SaCaY9+ntMZhOCaTXMfbS8LFeX4slzQZAFVFynIbzLA4kE+aU2QhchUElpAAKSAg
uZuhsJyLldJ39u+sYm7IjsWkg/5b4LaPMrYc1MDXnzSJ2lcqmhF0FpsfXkmSGjWd
FuBfZQei9lR7fMJDFaq/q0u7L2sbQ/q5Sllob6pVv5Q4B7v3vUCVL5EyuaT9BSba
wjSsg42ideuhlbspnYIAXrJURbK3Ai6sJG0D/xWnqu3ji7LKWKW88fT0gMgqxsgN
QfnlGjyGy03/N979AIyDIfLtNzP0Md29l1nXr2azzs4wTa65jaewdemCJa9nhXeg
8KDdlMBcxMnirZbpLP/6fgIobioK4I2bbWo9GzR4iNmIp1kGDzgVsduiIxFzsFZj
hcwdOEHTbIP4sxFSWrWtSuU/WSvQ5bxtpdDR6a2z49LEnps2WxJ+gqcmuLfnnF91
GdM43AlzzpqKD3I6H9QghOqKnpMheKjp1RA/sAsFQjQZz8OMQ4kXknhgbf4pS0N6
1xoswuU5/q2ouYmDlTNVrYGSDWxJLQgrRXDSlMkfJgkvv6eoceqRTUT7ndTG4kcE
WlBKaEIts94u8bqBKmoXqqD78ryQRk8zGfZ2qzrFXsESv+62FpZ+x72sqRidQT6w
Kmo5PMpcV/V6qap9wFDjxc/TZbYucNxwpP6fjkbkf4owROR5YC4tg2eMMXIHq/g1
olkMnnSKAKbEgniSDAf7srVL/XIqh8wXIeNrSohzQQvEIHNDYcvogN0fdk5RpdIk
LPqUglCBqOiPDhsjb2VNlmC/b+7bgJ4e1R9Wt56BI/RFJ2cbsAUaIV32mVCME0x1
vu31RCw/wpAnlnPA3+E76YcBE5Z/McespL35aMLcPzRqsTiCTegkNUEYumXftAct
cBn5NMtZohhZIBYlDyFMZr8b12mf5jMW+CYqaCig9cqRrl+H6onGZSFdDdfGRX+h
opUzSYZgpE6WCPgW3XEf0aAqV2ncmSd98YEmToTotd0ypovyqXJQJzR4iqBzFrKJ
ctgRCogFRqsHNLd+AYSaZW/DQYGohaX+GxODENQI9XeC0eS5dJUgi5wGuQNdMGQg
6KDHFtS9ffccf8SFudWiqQ5hPeg/ghk/lw6pWWt6T8Ig8QthTWp+2TNQbMv82LpV
Z4QuM9L1Zp2uEXF0hSY4D/fv6+mB8pa6p4T+vOHwzZ96VAtJq1xwhMt6R970lEy9
cJPK5Vc/EWN3K+7ZofYLX3hwHEF5ZL2+u5ONsIPP19T5XeIpE6S6Jz6NaXx11xH1
fI6YbYwqKLPVJ/L7NrxaTXw54o6yax8raS+vChUWb0Lt4juP4BIKOqMsC4+xwYd7
1b+V3yTHZJvxFgC4D7TUTGvwId4AoBv9TdXfHVJgpttkyZ98yK3Ia6jX6AjGJsCO
tjx7ILbWRBsel2LO1skae5EEEutguVlVV8u8Wz9CM58p96CdhywP0/gLAL/4mdA6
btvJa3S5zi5d6JzxjelvkkM7yDlo/IrSk1rSRRCzmtsSRV0bnhEYiel9jimIONdy
DxjXLhbqRQxEmoKy0fHohwL5kPhovgBF93PS53p7uGhxKYeoQCSEzwpyQlb6okSE
MU8wfW9vAGfa3JpkIHzOri0ZRcbezJ41Sc/OExb8jDDHlUGdBDL2mLQbahFqF5to
FCu/Ju+EQCxmPGjWJx6fXiWAf2pFgKWJ/gFhUFNtCXBvELXp86KZge89rD57RhGZ
BEuQbVuC8A4zOkQ0JxLDAHocn9awCtsAB4b03DP6KOgl1rctr/p8NFPuNoKK9UGq
jKudYaoEWZ37HGCrHHhmKn6nu6tWG65hB/91mRN2FCb7qZ34PH4q6nklH2v8jLRB
zY27WoQONzRWg1mjiSa1QvP/ngVDwZ5lIA99PsH5pgZ+uGEJVespeBG8y3DsYGyR
WhxMhvs/CBN+QBC27H9fZTDvdLQigToH4Be7J2oQukV1WTjpMF0ocu8aHr7WvRXT
5Y8lO0xiSHzEgqtn5T+boKC9NEbV43kAlfmwLTwWMMv4irf6Yc0I+Z1TweEU0Xtc
5XgG1cCsx/Uq7YACQpNoVeYFTvE0yQtzeTpvHHxl5xXpVUTySkICzDXSdwKVPRFi
cVvdLU7GxWAA4RJr+8cR1434/Vtb92O4A4P7K+HEqDs60GhGzUnRGpCqDuOzsqQB
UNMw25KnUQq1wwaPOIp8htgnSCIR9Yc4a2FF5SgYvJ2dVTSs0lVLlpCKxunhtc/o
J72UP6hqLngBlDrRlOd/iyInBfmNO91MRc7U3yb/qBN+vhADRNtAh1yKx+DhmM0g
LWRxbg2iiO3DeFUwCWZO7h/6Qsxv732bzonPyEvnPG3HT1QlCG4XzqYw/QaLdG05
/dnuYR3bvf7CNO5tqcJBsArN02QPMIEA8bN5CPZe2jotr71jfLzgs367grNNjLWv
VbqMIFaYIApWC5SB8y/9oFY0/G/eJZon7UyPuPQEnrwXlsSVJuLkEJUY9FX5QDpP
bif4fSX9Pxn1/D4BfIln3Y6mNJID9/YhHw54BO36tEYFIJ/ShqCr1NJiymx1ry35
m3ZyA4KTmyycFYwfHuFLEBCUYycqMUZGsCB2bDDai0XiFzPQs0AWJWtm/4RLZUL0
EAHZqcq79uuSc3jS+V5Va3W9VYVkXowIdgM0gzFq+E+cE9JK0Aw0jtFiH7PnLCZE
U3tLds+vJp0BdNHA+X0Q+NnA9VeTuPJcV8krKLVTI/moMU91jdSPHYHfTX+Eb717
0YPO3ldISnfiOUiEc0ed/rK0NiMI6z+8DZtoa5/JLIVAxypfeOZ/nvsqSZFaZUHL
LMpOGQ0bZnfjsz4t4GBplhnPJO3HSS4NYfUwkHAsTJKRqZMBqoch0aeTBmSFyn3U
1aX9xDpDt7FTmAIwGG4Q2daemozwI6nMDHel+3VqeqdPls2jRw+eDas756QFmnJQ
s2L3HkA8b0omE9T5ilpcukIoMRJ8/7HtiTlrIP3ZsJOHqB3sPysIFMJyCZ0T6fxP
5RGVF5Hm9rlEGfGR/728I+6nW2QJH1sUOYlY5lfJW6DN9EhGlslIsjknaWcdU+tJ
BrNfetpL76wPjMLsMnYe2tHMhksNZSvNJ9jaiL8FP+IVPFuZtoIW5wi7tMr44DBC
AtuaE83w1rFp9P8rvhp+MbsKvGoCftLZN6vRJ0fchS4hlvwxQg9qry2Bxoz6zKii
FkcMOBbVR32s+A3NJ1WhQF2OD+SL3sqVqTIsBB+Hy0OD9K1HKPYuKTDP5xCU9bka
ttjqids/ZbXU40u4Gxt2OrU7MuugHIRtvXypuJrwfd+6Wo9QifIiXGlEW9uzIG0o
WEbnfkZPnO8s4NHd5lrse1X8a1OJ6Q1LAalc+WtgMTcyh82l0aBrcLzeEmLZQ+W4
WlJC9NCN+n8JzOR0wqSdzrLoaA2RdQifz3pkl4wlXfIIksFeEOc2pDuubpyUSr35
YsRD+kJw+9Y29jwsOjQ1BLSibD5T2T/q9TGOFBZ/CJiEtSk74yF7TviMnOK6a5+F
r1x21bv2vFo0CxEiMSLLuygblg/P6syizy8H+X6m6xST7lb5+k5EAaxLhU+7zyRK
zLq/Q452fU5q9IeSgwEWS4DQsD186AncFA5aXYsVCDUumLz66wKIx7pFbT0wInNv
wVh2K1igx11VadX+Lo1ONALp87gah+VMlXpGAXno/wB7Mdn34NSerauUVkA9Wxvo
wS2YNnl5dvq7e4EaxaA/iuSdvn/NaW13tEYiY0VsB2HLXsqSTZF7NyDiCbdqVGqn
5YbFPPJ7BxZmhN1MhgEc/nxQpOseakaEoIIU4E0RsVCw+802Phh4P+/j9YHQTCuf
etfb3glRJDzpZrQrKbs32DZVYKWtuQvEozj/cKLPNvi6Q5IXJa7PHkH2hs9r837i
WM8XGkZOHz1YU8Nw/2D5u41syC6Vav+8JPCzjQ6hzDl5S6VYZGUpXLVwRdFswOks
sREl+gLSDMyRnThtIw/kQWQAe2qPb90xJ2dY6teLV/Q6bgK3Bm3E2yM3U5JdkOJD
8wrXUkK7InmoG3zt32SZ2PwrpuwRM8XiPJdnyrOCJbNkp93EABuUA151K6TtCAqS
yK6ST1GtYb8ru+mgAOeeBvXf0YrhSVyde4nIPqWQgy3TX/3mtD/nRKcodDJhb5tS
0AG20hOMm013MgKmypxsfK/MSmD1VM67xmk+TtdibKJHEuN6GPwX8ZhxN/Mhmb+G
WiVEWGwU7JAZf/JC3JIOWVVFuOdDFOH5kMt/wg2e+pOO7tIYUAu+OwmNuZTr+FX6
7RUjkrKF4zlLX27LECk7FWqd2pNvnzMzxVPVxhboCD5kQOZ98mOeOVowO3ZoyBT7
lra72eGe+v9TKOlR7kteSWFpPUVM+h1JGh87Y448a1WVr9PjNtHLqBLrZTqmZsx1
pe/THynnVFXcEXvm7gyFWfe//jLKN/WIEGLJ76kNGz7QNULTSCOG/zobBaay3/yf
ZK6dqRh2h6dusmShT1mTMDZztqguf5HTmQNJ02JTnay0msazN39/HfJBj+9LNT+o
ZSqb2ECM0woHXSdeB+7zFs9qFzDJ97VnINCp+kY4WAAqm25UDsXG4N0AUOnWKt0O
12OUDQPR46XvkSQVsRz+/pVvvGAF1CNe+yxFySO0GH2OngqJEJ7yNsSviomeArdf
mQVTT4fQ2ak+fikYFd30RWSzamSnR51LdxOwS8Ad8ZnD3HioJgbaMVLIMX6tkMS4
blH0IuVEDetOHtk1++xmmQpuDfSVaXQpQx8NOO4fwNqpRDRK97xAKuCOCVwIcCa9
vqKhdHb5n4N3u31LT8uWQWZ+6mHU3nXHBI7eWP0BGcDDnVM80V8WkT/d+z+zJF5F
qWZZSu6yOTpIRDwfQb977nfkafJ1Bbw0cJmnJPFS35vhbw6rpf+EneVySud8ED3z
R9i2RDsftZRy5+Yj9kVteuJwR63zTkOrhfD9TLiz4JsZLdZQbxE52zVlcp0Q/fGs
frBU48QSo29vLoHW5kHP9no4kZlfri3H/kaSlNCVcrjjBmgvvCQYvCBCBNcxjxF0
kEWXJud7x132zLB9hVVvpT7j3Y7YpbSCqZXhT6OVAv8vfpcrjTZteXe9VFHqNs+I
Ph/JMrmmoj0S5pv1JWJz77ekpluSKfRRrntiaSZulBPSODXra7FONySeYAimhrne
LtRYp8ZLjqGqW7wgxMnJv8W0Yap25rRq9pG/1BT0gMGLBOvpFByEUzGQBsbIXKgd
3iJHsWesTNew/YK3vMxlF0YJYI0iqr6lA+V6kaleKHn1IZtmua064ZPlXw5txxX5
UR4bwZG2lv2P3Gmgtvy1l6d4Rf0vGTCcOPTIKFQtilF2QJXCW1jT6ktMTx0wxhY+
WgLfocvE8SAuyi3VqDPTf5DnjpdK6m1utOqeI1Or1zQRBT02PeizbYp0h4icZMkS
/bZowvJp+o1b2JFeRyzw2GOyTNXv/BeLLJfQndmZO999ZOGP0g5Op7TmeVhsXDjp
ObJ5oZTtpux5E6+JZwjepONL8mJ/M37aBerAqA3GA8T0ixha5GV4aKr7j7ZBsXl5
L6OVXSP1AOFyD0/CwsNZ1cSx2s0lcsR3HEYYl8/pzRpX9KJmGHlvhkpaHyakUD9c
BUmUsn/l+n6ojIovT1bEjxlhhsqpi7R5qROzbQPk4rtOE8Ci16W6cmaVLQdIUEj9
1yDIyRW4bgLZ/qUlUWCelMiSr+onidBq6zPdQWgaWcTvBHfKVNeGEeTmak6JM9oz
Nt+fJhltcj7OMEFkYT7U6nD2RbzF5owRud59ZRO3rJTY7N+wQgMy/37D/TzyFeMn
Uau1VHAE/aGVzFPSXYkcs+PQ0jfBSbjcWQq/nT3iNAoYG81tEt2HEfwpCLrc0ziD
TiY0PhUfAXfAlPg74JlulmXVQnYowrpoBTCeXF1Ne0oQ0ZosoYMs8ctXkmNXtOTN
wDJbGBPBiCUkXkxHZozUeKIy2eLC/2c5JY0Hq7AawK6qAHy5s8SQauBMa9738BHr
fsapY/r48qFc9SZnHdTAbcBC6Sn/j0jL7pIOkOXxoZ4uBJ4/PNrBPQqv1c4ezrC/
WFDxmsHuBgoBz6ni8zyR11urD7IoAxMQLtj/3k3e6el5uFcN1DziqVoz1DvuZMek
kGufjzfZM4xG38bSI/CrWMJFF/hOTqR0DKTOF+0S7mVG74b9H/qO9tSTuoNnp/5l
chvA1/q/8NKe3jUmyeBftgPbI5IhkXmsSZ+LOD1rx65i09Hz9KY0/ThzrVQdLSUd
kkFbP1Lg2iy3+FPMPI5XkXqvJ2vw4RhmCpXycIgU0a72u2lnY9fAuDBPiQIw3ML1
e+qgLtg8Iss4VQlfsqYi5VWkjSmTesLsXmTSV9WRDFfQRLOLc1jSztLk59GKEMam
E0WlUveJyKGycaezqWNt5eRUntpmnQ6drR5MuCvPfvKdRRFiPZqSABmVf7YY1u85
yUCc+pFVk0pq9TGdMoF4l5oRdaDKR4FLtQ6UNo3SVdt6LWMfj7iaxyr4rvkI5v2b
rzmCQiaP3w5B9txBcuFQsTBl/mmlW8zlVbq+BmAsAMJjahvkUDp2dGu76pPSdyOg
0HLNoryzHtgCQD3ykbkDpP2UTp+X7JMC1TbRwA7GvS8EzVPOHXAZpB7ByziN33ls
hAU81udSiwpor7tX2YHm0iA2o4JNzB0CHcFLkpu2t1v6i9jZGiXy1FIESO5aHOtl
YusemvYzG77SkUg3eSxXB02eb9aZjyFLrQQseJRESMNyaxJ2kRBHFAFdg7mF78qn
XkLNF6yMSzqcQzco+VyhXMH0XXqJm0PTwLtXERutZzzATBqWyBYSxSRpMChTLV/W
u285r7V5HNRSFc1Lg7p8vhvp6SFxRJJ0Qb5laRjA9IJps29TOb4FSJKf49+475wX
U+DIuIj71Fr6/8Pqfpon6XdXmFJfbz6GHOvxZKPfo994az2e2ZQ9QGRKg9RD1/B9
sWq9MzSwOXxKHugwCg97e6GL/zg1180hhjErDLNfbkd2JqU5E4dLQr8KG4SoCdtp
SuqIN1T4Y+Rifdj4BNj2lq68MUCwVtCkfNo3VIqteHW8vu2G4gxrLttH90fGUZJD
/F+6gsCWxKmaEut76iYdQWhQzcw635gTspmJM+2ZQcW0jwbQEBlP6DG6l3wT/SWn
ZpJbapobznrvM1haM0/lOaOZGvbadquGbA1qEvLv2zuYHiImgf9Vyd534jOBM6/e
l3zBLJOeoWZfPhIwECtARcTixjz8YHLeNok3SkpgAQ1huhp36+Ci8CV/FaHGNjz6
BWcnPSVSlGYjrOi5AtaTBxfW1+euSLA0B/kuKJPGH9iPlOU4kEAzS1zVugELBc1F
HKUVLkbGtPdq7sQFIemqczJLhBt9iBGJ7JHFnOPWFLCh3IXhlEfMIl5+loLmG+9a
gZbjB/pthC+H44H5oGDS2lmJeUzdiwFYg04aPmaYkSeO8ceCYivopIyK65l7mOA5
Yea9MDhfXyo4T9sv1yEkhgC6PdDbRZOV6xCdw6kspXj4wSV6m7xblMrYAvuoEaFp
AN7OvjAqyOO4Z1Aw4y1xQu3Q5WblQo8KpYMEKpOkzbwn+Xo93VKxJ1D96DZ80KkY
xQYhsxD+yfRy4gIddWqyhsxT4hkZQBWWJN78xmTAh62k+kF9RPGXMQGBHdCmzy0I
PkbgDD/clh6gwoN8QnVytUukIUnxW3RdK31rSutxCN0H7LfzuaibYSGiU+x5H1RH
KK1b2XCGQBjtIPHXbTkEr0uXRy/3D88qsn8RF0IXAAKbvQ6yTFifUjuIZMTjQcgB
nGvG4PNx90TdE9NVMCgDh2ffd3dy1kv6XETTLNYEV/+zUAWTvFn2DPgAcDZpq5PF
xyrIHeZnd68h12YkpWVOcaSuhDj4epVtbBDBDj37y+azYTIfxr8PdNQ35+nxCAtC
NYbpgICGIa7O40HaG70TfjFb0+Ht9Mwsdiz0Zn50pEAjce/OMVJAWH9Fi1yGkdcb
Q+kzXkRZqCmUPd2gDeJklihnvPmPF7WLB6HA3ypV8nVxswbANCY8xmgeGhfkWJwI
bMenLHvKQ0Qek188r7e2+2Vl9ckEnyqZrLU2LbfyDEy5R7HY6vXz9bVvwT2h/avR
njNH+w+BgNetrxbrkw3Fxp5V+U8nSATdkCHklaw9v5rW2/BRY7DpeTDOy7KAIsEX
+257UQfg0c+cto6xn+XIm05HGNGiNPktYxYoGI6yfj2qdg7zUHIkr24l6DFmjbOV
WyE+ywSlv4WsVoZ9GL4hIYybfNC37dLFLec0c8qkKYnhI/+78RM7ZFN/P0sKM54Q
fh4+ciBCsa1mnkiBicOLITlTOvX+z+kcp9hrzCOhmXZYSRNk8Rc9c5uuX1diBM/p
N7q7uShtvAWKLhfKM9HKJ6M2XNmR3fj40tQsBJUHUwNAnv3VOSmYXEHfNcq5LQpK
QPELYdpxWBStbopzStiedMBGyBkx89BsmFJeVbY8fw0o1WrSNsbZNpT+WEnql/qm
CW4sDw5G+lqhPDZgTaqw9Im30oGqbUwfZoCWh5MOPLI09SgrZkRgnsptf7/BqInf
73czVGDmxKN9Rs8UxjQR39kp21J5C2hBTX21lSrgWYp5hXnkaS3Wh4kwwd9t1yAF
RZucuc9N48TooScT+7l2t2RsT/WWYJKtw2TvQXiwernEz/gcxZ+5VkNWkmKt9g49
eosdzQjoBIkZOSeVseekO187RFXi8wtJjgrFiByyHli7Os/8PvdPu5CHTDxq8ByV
GSzuuJtYVKvg65NXCt3VhSbxDpy/6mm8AGFk4SuEQHb6tLZRIvg2JbFwI5S0r0JQ
WEhLviWGjz1iTyOfdnQMFO46YvgHgW2OIyQB1CmZeNVZ6WIA6zjs3VzrS4NbHYN0
7ZYBo8/8WdBs7VjHtPwmkMIYX2clXwYvoUmTFxQ/4NzSetpjX4TYjjtwhOJQBPjv
jBs916gIh3hFu99nG24vv585SrcHDrWMCVvVbhzm2O1ePUZ8rFVtULrmP28Leyjp
54QXsHwDyVGoOgtPusklHvxVkBzTPNcdIKjxjwPtLKx1AuhZhCzKse0Y83ebdxpg
bOLTaKd4bi3yAIzKSlel+dIm2JQAEkiHADOgbMZzrOTprwUx6NhsJi7iiA9pM/a+
8xml/WZhIJ9tpn/sEsFDaJjV7rnyc2xKcfBgBlIBDax4jTz7nchAf65ocfkF8wxK
6JodXXmuV7Wwe33CRUg7hdx/JlciQFyEJt63YpT3MRxTnxuMQVdEeeK4CapRYLIM
rcbtS+yDvbSuv6xuzuk5pyQ6jIDlrvTfRaHnV6K6Y8p8EsbTg06OuFPxYWWFDKVg
5Zsso2abD4eYHr67BebqP2mGCS28t/6lYuVyBJyyyf0liEC/za5ynaxyVdIRbVfx
vd26CInwLlJZCEm2E/ISWT8kpUDY6j/WLr5F1SfINewI3BTN2Tj2Lg0lIdG/1Q1h
/rHtJnSkSghw0arV5FXoT7ktWlO1tYKtNkTKgunu4SElxeSaUGgDwJYNhN6VYUpW
6MtS/mt8DJR9MXLC6O7mMPp/zTo0a5NcJw+9+uPGp02mPN3DmxnKmFYZ7KGdNAgm
j+9XhlqQ2bWX08TBaZHkZYLftJelYArJaTUUKjNfmCEiUoyleE/tEsKXDOmxZCLG
keChY5vtzsvWcZDnsSPGukdRsUHSTTJAZh3T+gKsPNlxH93YiUkCYTUKEy0Rp5bx
hpdeEIyMCCnyyG07fPGP7VsKH8kFdEtFUQDTfNMOlBnF66/flH7461173cycF9AG
pnvnU1zRJyAlBH7i7nYj/kqlWNRHbnBMvLpm7NpJJvqpBpO+dPf9QZwlAfJL7L/6
4uzQoyCr1I5IuGFf8aPQiWeBemCPaQd2qvQ2xqGrpd9KsvcH1MYOROspq26qg+9L
e15t5Ga1sf71mYLeDJHuQxxEo7rg/byWupETZmfK5OXN2KlWNas6o/bg3sO8mThb
v7OlbYG0FiumO47eYpyFseVjCO4l3Rw2XFMSsQkqZ2Oz+LW2mjvjs4KSslfkQ8UH
aZ2Kst7lULAKnoenMO1KQY8GvZRxzIptMIb/81tU8zdgC70eju2E3K9pPKxxHrCL
MY04chk99eWqxA0fNwxdHyxSEEp7gTxTece8h8jr7gjTfCYkrmRgzuXthaqBQhOd
weDcjBGCumdoZTtLuH0egRTKD0gvBgYfnr7fOluCTYQK1JhfwmwMv+fFl5FEIt/T
B7skJM65+B11fxXmuDib7hW7Ssk1AhFRxKG6idvvlpFcYCxgNP7B5F6/t95m8Mgv
NApAlhSuLz3tt6tiCGwVU1xhPvCCsWIUsCyNPhr+UNI5pAk5Mgc5Lfnx0pSTX8Gc
ZRDrRDGHIaA5OuwOgxOOnGCbXSSxpchKMEKIMfH2JwgqhgsaezJ4ZGjIdmzB5ZPs
tqfOZmK8CCqRWXBUVrSMkQea9YDDvixZa5n9Wq/XxbmOPAm9SXnfcTz2fvTqEsXI
SnZc+sZWUrR5ublbORVQwpfK2p6aNb/GnW3h0ivI+nY6FahXu2b+1rKKN5glCweb
43Sag5euzCqsN1jNpI6ZI+bvko6Sr5W9/YlNn3f9cPTw3EacoJhy0QXABFL0jIAe
/0Qm9t6nGuMuJnBO/cqEWmouz+2a564k73HnAPtOBrUTqUpCYkjQ21RSyxYsDsDP
ScVYxc4eXQyoxAWRKwVVjwkFNZBoKDw0fjBzDqLd1Gn7kRFoHNWIiKJddmuFmPV+
LAAPntHN4tZlc7MFuiNaeFUzMaRa6+N/effxifgYk1YhpjJkRv5DU2Fho6fEMAZV
Cc0TmnocrMXlwHO420fdQn2g/RnQftG/G9ZYh/16FDRNlgASAokzW69nNfCWcU/R
VDHfKc02RBJW1As62YPkkJ1HVk6BXpcfjl0kIJNCZ0jR/29bT6CNMlIxauFBItLL
NDTPymIcZPPm3qhlZq8Yrlj+2VrmlVwPZjnWdmEfZqDbzETK+RsDAk94jdo3OFYN
Lz3fy0rwNb2XSLLJVPDidwCJ3LvVgHywdMxMH660CKBe5tcR9uGschJwtSzSo3uw
hPDjC44X81/QnwmnoomS0QZHwIFHfRlzxsBATXLWN2pdSYm36N9WljhaO4NiB6KP
xt1Y/bbacqgs9ulWIu7uusQHdBxKBNW6fbxP/yNnqL5q+a9OtUVG/KS2e00nm5A2
NkAdMuD5eGGQ8Hrck09nbfwEBd47WIvGx4Npo9bvYLQfVIf3jkxpsLX8S7XPqAIC
HOdtoM7jWyx3N4aeRQy0C8PlYpvwwMDzKSB3TUPLtIDK6uf86aDnCepdw1xuq5B+
xhHP3HXiwWoHxO2xRx3Hf4Lmk9/lqo6BSS6skdFJXdrzez15Q8TRadbDtbq5Cdk+
uD7hrk3UGdGvj5j9wTBzvQtpreSgGFzA8niWVlh37EACXxKGhSzM5Xukdf9imR4s
QLXpsNyx0pY+aGC6W76OM2DxwiBnb5IqX+LyPJMeqZ31vE7RKvjl/K6QQ3tZ8GNU
TUJISO39Ym9gug7skMPraXxQAOrmjCecZ/uSELW2YgZTksGkwh4t0Ch0uhdhWCDA
FS9amYy1+gT6ivh/lOs0lEnDQ+PxcA7I7Iz9DCWzUv1/vUlGrycpX56eCqEo9Myh
PdVAjd8JnQ86rj6cJEOLZUqJNgKYOKTsulDGnQ+gWHkXRmyGicgJnlelhxPRxanL
r+NXRrDLmq0PT/epuTgCIa2ML9ZD2djNRzi4c0LK75v8pAPbTCbZ+atsdKdVCrAg
c2Xagp/oO0xa/q9j8tWyXAPA9u76tbUNehD39KzHQHwRZjUPvvUeCmL+shYCiS4V
+21eOfDRQ/jjWMLDEHCGxn0CmkNnZBmByi0udlLrVPgz8tpKqKYnkhtwtRz/oiO8
7PFL4nM4+HUjjpj0ujrHAv8SP4Vo4waVmlFnVfX+ssHHZC91eG/8Yta7PWcMcEes
/tHpesmN4c+u7nk20saRB+HaLule8384VPmdoqXF3rmjaNZhU1K9W2MMi7fG09Ct
U+9wcNabUegX8esLy2+VfcqXq8dV2TiY+6v2Xds1UShSpMPwcHI+fvaH6E9Kjqxs
qqWKWB7nIUhLtZmV71WfnPcc9XvKgVmP/xgy9Ck0jRT1oePgjzdIm+RSFCwdxs/e
yj2BnDa5ILFYsxYwIm1/CmHiL/xfZJzsoJto2xrVPIhRee+pDIwNWjUt7ESuaDHg
7c0rMH+d2PTSZ5tP611bGaKyA4H8ql3zEqDDenZAjvR10Sr4pnhgUwi+8sKBySSX
sTbuCgG4kMnEZFxgBAmSUuzVUlM0JTJ85ROWxH3iMK5BrgQ/uCfWkc2VdECFFElM
EaBP8QETzH21hK9mzUM1+2Hh+apE7M3yHoOcvLhc5NU3ANWnYwsRcXSS7gEPH6f6
8+Gj8D5kJnoZCTMVr8mvRnEkxu+/n5EX6jaD6KMFr2iNs01B26gTAVZPnTemBOMn
aduwFSM41wfGckeOy7zGLef5c+1q+eLsbE4JcIzQp86sBrXZlUHPMOHtK5MTrElp
0rPckaOTei5FUv2Gd5OuxF9/XZY0TaQSJCIqIWoPhSMogsMdzCeEZyifdxhgRBpc
f+I+eivRlWCExBCGe6QWFx+9WTg8o5KIDF2Gig4fSetpSQiPUSZNUL342SQck3jS
b6KeOx64AI8sOI8ZhTUu812cFqMepiBEhyWwAbtJC9lT2njzHSGMku/WMyjT1YJ4
IbJ/8mXLclPfwNu0pW+b8FG6GsEquok4zIo9IVNy04GUe+d19Kj49u/e0fWWu/1/
701LxCd9uRYzu+hP5huGrO78KbuDj1aokF2mm3f+9AJjOxVThoOdX8pSX90Q9WGA
rw98ieCmP9GQ+2px6TXb8d5qgOYxYw9F2EvqwmQiP3CkWv9+Mjio6sKDAbxlRLB9
3vqDU4SECzdpt20HUAzt/Q1hW2ZtFqrZGJr3TgmCrTfSQ7MRcE197zoU/hvagzcW
b2NKigHrT1C25yAbkoT+SHZLsntpA7JPKiEmdbsM0w/UU8hTEEQsl5gZCbhLmAdc
Zw8+BhG6215fwSZ19uqrjQNDJP9wfJZhqkreXL76glHnlkxwOFHRNmyn4uch480F
VRwIwN5H35sCHgwpEequPO9vWL+bFpO0OFdItAs5VIQpP/u2wQhkcrruij0SB7lO
NsIjF2pamMljbADpUoxOyyK1qlUIBV/07qE8YO4VyEuplBqp8Y7W08nBtdzbbYaI
UUY8RKrjwHcnSgbgNaQg+tBDo+ZgOipbWBJAc5dmKWLRdj5Obl7fxsCwL2QCI3MA
VILcFavmi5jUn9ErPHZ+VjH9fUPhVJi017l6BXolLuR0oOU5l0zP2NRvPBKIv5qS
VJBXGguUivu6yCZDdfvZB15YSJPJt5RLxAKFxUiTTOJ/ZFZgUhAmQQ/EN3kXnfiE
DyzYQetUBGLUspq57YR7JPUXDXIPpM7b5cM//NCKOEOGiv6CZrhmLFj0ljDIM6gD
v4swdc+uJRf1DGdv2sOrYZ3fkN0tVO0f0/IOgZdqSFnBNSXzwkcY3/qYyECT/Cny
ORoJ4YTT0LaoRQh5QKkEFJNiJl+72YDtA2pVN5HNjORxEe0OyMRjbwarJbM5ZLHs
QEY0wBgtIvGPPMs/qCLYQy9jaFOi3KFQDOHfnpeLQtWyRVxZybWc2eaZyytvkknH
OghXN2/rUrr8Yu9opEynrLnKAT8b0xyCLGaksEasTyU803Ng1HyULJbusUlVi+yb
zxoHwtatrjg1Y2ddeDFhuPc8H2q2r0NGu/3+VrDTS01/Mklm7TFOnna67qw7kt+L
BXe1TglgXAQCggKITyyXVbQ+YfP/HuSqbRiooSysDiQ0eAYPx1Dp4dmZNHQESQZm
cMXxvNTiX/K80GNO5rPsYq6p1X+nXvU6MP7lWNG6+Ia3CN/azAAOktCxK5gMfmLs
DMgLj6KYdtc99tF07nu/agu8mkio4QaSON2/A5PoClbrQ1FQw/LhhuWJuoRJQRES
9ucr7+mpYb8n3VIYgqJB1B98OrcYeBQhDnOSvCdpOFdL89WoRy42hsCOYhCYIXCb
Xkw0/WSEriarLgP2fz+yC0GYyQue+0xhOX3cfsshB1FQFFEES1E4P2pf9AWMY7OB
DQxgMvkoQs/Nz1Gy+QYqR1VglMNko0zsGQpNpnEzWUGfn1Zfc37UhQ84fJeAb4eG
JI2o9VVq4FKfvcP9BD2xKXfNDJKqlxmlYtwM/ebcf6m74HvSQpDTuxXtt2kPIrBB
35pKshyybAnpKDMPpmssVm91C92KNAh+8beTwlxnFhfn77AVDM0uFuszPJwItUmu
lSjwgXkt+DscSbURdZuJGeQXZb1ffH/xi8tyQCaNkPqQuOU5XhOitjQODt4LV7R5
heCl5z9KmSnzaDJLg3RHbImm/itw13cbGzaTZtJTLOsVvoRcaMequjPhfLvSF/tr
B7zMBgeezdSm0owbAfMctp9NRIgL/THdxUId4nvDl7T6DyNfb3Rcrw/m7/d+DEVe
tukiGcyNSV/RCDrN4mnScQ3H7Nx1Aodbeat87hU4Z1v8t2YnpUNSwoY1X5j4anb0
/acRZHFfWMWLbT6ipPvl82jkJjuL5pJQRWMdZD3wjJtFeCGzHh7lV5ZH0WQK4j95
QG5it4MzT8O8joeS9ZaPoAgCC6yEp8LegKuXxMWjvW1JnoZuo2hTlFZM8dSxzJEX
nShp698Go0VF73X3FAtW41FmbaaOAt1+cqSn2tgIxN9zDpxshya1w2TCOPGkdW8h
7uIKYXSVPIt8K+6ZatIZBeQU4DzSXe6s18ViqdRJbt3ghzI9KB3KGH0bQn5hPCr/
/4GD+fzUKpRXhftQ0xfYuBZ2MADffU/3pCd5uSm3TZSoePfgh3yh5yCmk2Aq1jbY
d9zvL1LR1nLBKbUxvlKYp7bafibHOiuq6upCGt0fkvyxGCy+DgD1L5YZWi37Fs4I
myeUVOQJTX6cHZFaSIJMkkabTlUXK8iFIDVAojVailvng6vH8ABpCX9PDfjiVRtr
iNJznug3PYrMcT17LC69b+JpBpJdowPCo5ctn7RHZ/qH1GAF21e/sqxSE5FHUCjO
BMi0owXHF5BEj5N+Q/dvmDNx+UlvYn73dQOmTfmGm09r3+wX1vWqRxkBu9K2Xg1i
JzpxPiePbUMdqYnsabMymQf3a2PyL8ym1sPnaELYmw37dL6jxlWM3dTyCQyk0tl+
wdWembDMVYz4Qc6e5ZOBFqzG8v5qhzAaTHx6DMDXWG3gfyyuem3lWZvF07eVFisP
UdOj8gixcJlOvJHGTF1FBHRO1ieqwEoSMVG06QupYjdfMIMFLOnGhfU57l49LIKe
JPGUCJHTHtvApj9mktzwnLaOM1d475DeHAUk7sy43OBdeLjpnPNMTDrDcduab+1x
0XfLDi0FXyDTfw7zCGUpi4V9JNq7SVUkZK2EF3+DOwy+20bYhCjsR6fD1rWsp9Os
OhBjbxqPsezdzQLOlMoRz0wxnsxaEMNUxX2/JbuEEEFFWXzUj5fAKvlMBya9R7Lz
NriHOKgneCexDTNZtNwO3bTRDzwLR1t2OTIjP9CKtpSRweMqV3C0i8bOs+fusEg9
n7lbaBRkYKVS0PBSflkPe92WnCuDxAmOID60CZEkMyrR5by8uBfol5jHIREB/1zb
N9Q4O9WVSoaMoXKVS2mLnlj5OZ9h2oqgIgmgrWP77oegA+HTohMImndEn79rr0DB
XYTUqFGoUm7+dwzNs1SPjWqMcEmrVcLDQOYyFnNHhs0h1dlXLLPZ9pVi9lCuarRk
9raC0JAS5gIgs0LpEHbrnO8N0hhyC9LtBlK3qIzU81VGm2UITPfX4RibZfixfpn8
u5kRuSsWc3TkhrtdeAw2p9WTLT7XjI9lO/Vc6CZjq3DyDiwS4YkSLEx4BL10pBfs
dPA4sBmEUQ7egJElriKFiixIZig43xM6R3IgAHY7jZ/fkeDs/YasYRsjpqSQHr8r
JxWUIwd5+MncTZC6Yc7ZjQsCNBXFc7YEonXU8amJxAimktOi4FqeR7AKtKimIm6y
nRV9zBm0Q8IEmEkRtti2pN5wbd+E917s/LNnzqUvcUagY+5hffg1JisuHR3gG3P0
5Kkn9g8lEPGangVHC9EjMUzZgPSRdNVTOAUqB9MdaTZMyzR60jS57Mbb14m3k90K
JNERr1s/hMfz04vPFwmrOMidBCcZySzxxevMEsf5ddgl3nSo8GGoN/8FzErlpxet
VBOI8uC6b7LSCtfR62DBBntlC4rXtLDEgYGjTsfcQJ8+fIlTM0VCYJA+5l7HMfLL
1aUaIlaiSIYxJoOBuoHQ9DHjPehs1V2QUWhXwkvNmFcrz7iXPUp4zeGAx3Kn3Wgj
Sk2WtauTN9SDXfHqUiBwsIO85Qk3t3FCOzBRRtbVZxQxZgq5CkL861nHFwIvp2CB
E0NF/Oltm9rI+O/ZLWn9YvPz+SljXkC1zAn3RRLD0CwRUxHPc8e1HMxPwdnaOa7D
vLkPqOdj+QotgAdzQK/hgjVvtcPCILz5YW0RvwDUkVxST5/qBd+zJX9GYB17EZyL
P1aA1hO/NKZqm75aCqzMatcfvLg0alLCEo5K5Q5vyF3cbqnqFaIoYsxhxSKiDP+M
XH3bU6zmQgo1LEo8i/chpVAUKcT3oyKJZvGf4j7plL+KLLFqJvRcuKXCnahRBEO8
1X/v3QkQrIg2cSkMgHMqobo/IDSt0IuKmWr6DSUQHT23FL0qRR3pWc+eQAHn1zBg
UBHWIjFlKZnYdRHRZw0ozolBKcNq1OClJhkZVYYywwRCaJNkv0GsfedihYHFnOq7
68twKj+XGqH2eNtQXCZRcToA8qkpxO1beh6ptaYVPKS+a0+9ncprGwdtdflL+Fix
GnhsL3eNWTLMSEREWiaJBfKAludp/s2B+WELl5syyKQmgpF/TuDvkRwXPn2X72Nx
Gq421Ey36x5CofKjKOO8OFEEm4Xj9qgEtEDGkDNE4del19GoNt8KducJY+7OA7fv
Mw5fWlS9nuSVjFtHznO4NdnvUM5PjHEjQbf3FQyIFQTl8gUhocKsGO3s3O2uZ+pK
kKnifGHJDFAVfwxzbW85qkH8r7R9PPwwfR5Q3Vzyc1IybzvTHxoCXLvcZIrz2nL8
atSMF2m8DgrTQYJ6UvVzqPFF46A9E6GWrY2NgW4/EFrtaXibXRyWqNvk6kteYyv0
5OlelzaxbtPE1Y1fGm6QDB/JRZdrjIdpxTGK4kvgoWB9sNvM/YCkkJceVlCySq/e
eExjdOc87GZ5IMsAzAfesw7eyshElCleVVQLrmEGdbX7mBkwMqSh2bn+XEhUs/KT
tzt6U1UuJt0YUKysvi/SwTL+N5/+8gjig75moopQSALhJi0WvHrsi2nVZ678UfR/
YW717EmsEyKpX2VYQKHOoBYKOJdB2lJAB488ARP/D4AAvY/wSsmHlyUqqdvgHJ/t
1J9l03ifmWTvuEHjdUFk5nmtd7IPTynet2wLSQpC+JM21soJ3CZaK7KkpSMmwrWN
eVCyroYJAak5EcT0hbSGFq4BoFgtyiU3wTNcyMi5kiCTy9zAS+P3EHs7ZofQLhIH
uv/AcIgOXcrSKYx5RjuA7UFs05JrH8vlQyUAa4jfQm2z+K/29gM7oGkpxMRr2Jv3
vHmD/ibL50UEp0I6jgKEnsPqH4uLoI1Os99L3EvaHSZXOLzL2hDCj37qzsJoyHFz
bLs+WU4M5yd3DZRgTQo+XSXR9OAw2e8Euak8kXihgYkGGwEWb0i4++bQYGj92HoE
RbZBhpItThpVIHdU3YogmSanx3Qh2cz4tOnAuvvS564mP9XgyKZdkn/Q/OcpSlUf
FdzOwSO9UT6KnajGB0jYGtFb0FhpYgpjRVI/oAMGqHnP2oS0qKRpgs/CgQ5MB2/s
hxpXQzgjyXIV+QJVhH00pQnWBQMFNSsFykGm3Yc9dnMjT1xFNKdDdgVXUbIpUokY
qdIxYDOotvna3WRfOIRsf7RHlZ5ogsmudwtDZP7vFU51bM/SaNNuorYRFijf6OAg
UBH7oytf/yvx+l7/mmUyW+Gqq5eD0Nv/z7Myy6AEQ85R36ArQIdti30xWTu8L2hI
Qud3SEERMDqGdvDC08dAMu46jFMeH2cR/tBp2eUL7gu6Ra9UJCXczQiF2bMWuluP
EmcD0Fzhw3JP0JY2Vw3qql0PR/Pl4IfIGYb03ah1sv6ynAs6ULddRtSn5x1li1jP
xwjMfJ584tt4UKkzvHDlONI58KM9E/lgfBs8mdGiJn32KbaH1yNptAiiGATboLk8
i1hc1Gz1LedfXmb0UlDu3iwS12MtMyZnenV4FOxNYktrIV934aCdy/PFKxOvIVUF
sipjAiSUZuJnVpGURoyOO+l7jpZuDv5u/ZhUxbMrFd7nRXjK6h8SA5RWUaFXOaug
CKezuvUgTZ0RofednKjAeAzkj3FC02hdpvqK69KLAy0sbWZtG6LC/gPWTd29MXZs
QaPtZjQyv1HGXrn9qV2LlrohvOf3X+zAzBv9CntPdgkD+hOnlaTuZVhzA7AQdZr4
UAJoy6KeoVv255VmfC7WFyXDrDTFyQp1Or0MpHG/xQcwYvIVGd4Kah4a/vj7jRIz
Jo0qazpLJDYvN5PheFs1+liqFu7C5bjA92KuSN5FUR6EVjfC+jLuDwbktJ25vuTW
1J+gIrygO4/Ofq+Z0vl27Y15r1jQnqShKkjTfqjmYGyKdeGP89LUMAgBx2v0H2X3
ZuDGWu+39Hk8ypXSXcngu2fBKnY7kcQft/MXkyNDRQn7vTlltC9kLGls7rltZBmu
k3AJjI/go9KLeqXpr5OB6UXCokLkg6/LhW7USxCfsIhMhgNlMIskctUuGAiyk7UV
+MRiqCiLQ2+TkDN6kR+ZKHy18SiAlsHszbtN0wfc/o/ZIlhIlyh4dZAYkgRaF9Cf
FRUQaDf/uaOPbosStBfDGYvjxfMfsozy8CsJ9u3Rh3Reg8jzl8eFxl8YVKyxz6/v
hP6oBJrmA3HDr1Ept+bE6IfhJGZw+aroP9pAxwV+XWpBjnZ+S9U7oScA/8JSBqaB
TYy7Do17eWh0EQBCySjbFIFKRCPL1BJAhj4Zyfyi3EX1/e2XWwu4nYIHdlJWJUMX
bz3qOUvNqgd5v2tF3bwPzHJAXa7Dl5vyXXtnH+r3LgXDphnmI7hJ+FYEOmIxzUJw
DYR+wZyV9F6biR96aFOvFI7mvX/FqkJcY7980n2kt/r6DtFHo7HToWOAe6RxbyEM
vqkLIg7r/8kccnxY/u8wtpRTVJawKBHREpCBS21lVvS2yvg2/S9czNXwCgSenkPz
QKU3QnSdWremrO+rG5MJaR1Y1PsXA5iDmXxynoNQ5GY=
`pragma protect end_protected
