// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
g1wIf0f7ovKxs0vkuglKz3HrKQYuIWSqK14VE6U1NneU3/FnnIewswBh4P38XJNKFHXh+HnSwJTt
7V10/+sdrcMuldo69GtsynG76zZMXUP5xtyGrzE60ujq5/QOJgqTx4ZPs+IENRpbPPZCnutOftyZ
OnPuowqdUfPTDwIhgH3pzGoVcSfJlQT1QLuLK3L/tSqmrtn34Ms+DW9Y2A5spsQqRidiH1VpafyG
dUKP9dgScMmO4hQyq45hW1LXDigNVYWi6mRooSQtAFvYEcir0wejOCp/IfiaRGW/X2TlbHI8owIN
Cyhtbbqe67xlwDHmvsgbFGS/tLqxQchVOJcx+w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
vFkFzugH3kS8TlB9gEYg8/8hgpGqKSxrDbaekNdXMhA5RPzwiQKl97fHF0hZRAoJOPTnqx62r/F5
6xaBvhAml83UwSGlnqJYFPCsjaAa8eC7qyBLCHn74BSI1tU/40BEvT7QlTdve1jQgBLy/qvHGKYZ
L+vlH45E6gaO5XSvU13NsLS5EITQ2RfZvP7kjV9zABqFoOJlKJeLXLXg5uTV4kXeB1bE7Ke1qzaN
Ki97kEgeB68y/up9WHOtOjzzWvLwZTW6ZSlA4umSBBcDrsw298SKlwxV9kWF1yboGwCR++niMU+S
8m+Z0lBhpq/myLA7IYvrTKJK2VJCTOgZ3+JnyOCVQewGIJ5ZF52a4oIHL9PimpuQRDGOfI+Tm18I
AHz/C60TQhTNi14J2cn8BFIyr12xltx9yyi7Jj+jZtD9mo8rClGkki/LaJyS4iLfZCkQ+m9UEJeR
8lUs2K1PqGye9stc2i9n75P9SQwQsCJWFOf/nrcOUglGpXABG54EDvJPTzteWUEM1XzjChCVk9GE
Db73SN6P3g1uWo+vKkFryJ3/O0IWHgWUP+0ODq48wvLb5gFqlNcS4onMiyseWyrUaa5Sg/3z9OFT
0Hyka54hPBBA4uRj2jY+2wWbNaMGM09QFgblVX6g2FyKVtWFBpnRqP6RxWsEf9E9fer9b13vw7O6
FC+c1p739NCo5GWmanfknCO7iArQ/KVFnaayeIzYAbQ+VTRjoZ5ZrIPt+8W6LD+L1yTvuP6ky8dv
Xs0asXTEXatkeGD5LkNUWjUmfVfhTfpWCvrExLFa2pd3JrvH/4IATJCJhjTE8sMAGhWivri2PGBr
FMwdk/Jno1J181z6GRgBipdw2gA8eUYuSmv5tNoXvWfG50QJWxhf2QMSnG0mFBQ0KqEGImoK6t0e
5PcApiq7TjvEYAjhiJC0EKAXquvrte+N0Y5tfic4Enud7H5imSMVnBRhgyprWMp9zI5U1p8GxhfE
t00AKfnCdScWp9ccq5fdO73idO5takQ8rbhoJj+DLPSXNHqne/1/3veWslDnMaoyj2ZVBLhQ+M2B
5STd5CVXFi9la4hrFIzSDs8TlwmV43YbFYhvWNmCDxoZ1bzBG+GpK+ExwNdrJ/8kqF8cnQK7iNuN
HYFl0aAl59JgYs29WKpu+1YGhOhySkuRxuNDej7bS3XajQF48c9EJuoPC9LLyypEagEMt+CFjvUn
SRE8LtmkNu+wSeerfEqjZIre6WnNVunCmumUFt70epqq4Q38rTZtMq2NUw8EBRsijq+xIT8jgaX2
SxtHZNmmwvAiIEBjbLefJgHAhmlw94dm4Rc5UejROMEZF4XGa9bp3wflZkc4eHulM1+oJZymqb2T
GVEDTlBOM2r7OMsUAoREIc3JydlG7HhbZr24NsEEiQMfq0MT5QcAi0RKDNqlv8EV1InL/7iFBGQb
ar5mpBSlDH9+fcwvea8k170WnJDeIYl+PgEd+AbhzzZw2L6uriKGaarpM8nVvL9j2I+5O3NkVKHc
L5NgN5b4cP0S2F9bQDQ+eP0IyjnVV41Qv3SuxLUIOqndXOhGlEbU9sxN55BI2p2j0QBKIIYdmWqs
1ZYoX3CzCaNSc2Origo+KOatOgUe1rDhsUdp6h7fr5mA5ISCYVGaW9gdAYGZJzSBub3o085kQBJw
pX2YrWrmBmyNZWZBawNgg0AVnHevyhCzhneBAjZ0eCYDvKuYhbKoi6mbTD5ifE7Esi/Vkj+hBysR
oCPfl514ypvzhTzoemjBlzjA8YX+iRTKpkBuNBL1EEW3IcJlSNMdhpUeR+m4Gosho+IriNqsQEek
BNXUpG3eDl67aHv3DEo9Tv5Mm2r5TpNVjSBhmfnu38b1BdPK3MFeWpCwJxh3EK2XMgoKWFDLMZfJ
RsweMzWLswm67XVO2eQHnc9TXhjs4VhCrDuk/OiI2xZv4M+ru/9SlNUIrnETiOZ5hleK+3BNMwnw
6EOBIIlIlQVDJaLoFoBjvc/TEJvnyNy/5m7Iy5Q7ijKj34DHDlb6bALV7qV9M1fhHvchIsy71wTQ
h/ANIZifrPOzuL4tl4i8ZFH95XJhApcIpqWZBRBw+3/gdQZCK6cPotVNvb2l3JK5WC31VGA4mUHr
nKl5Vj/PqQSRwUkavJjpd25DE2Zh72pWmRkr3t+SnU6N9TZRTvOKVVTeMIS2dCJ8U4yxk++mhFpj
ixTpQf3KKtIXAshOBngBF4SOevwQ7Oiy1i5wTuZlS/6CR5VsiRHJKjWZ5gBa2T4VodiVW6dIdqrk
j/kcRl0cVpIyf7BEMpcYHYiKCIsFIdx9I8Pbi6/0t12CyqlzjdKBdS466BUNXSb0FBy+QoqA5oSX
5/kHChumQNYmPEkyOk9ZorILGvAq23YELOCt9Rs0ZzlQurTYgSRwjs24hI0vdRMFCFhkXsya938b
9KpG2ZLYiVplbeOyheiZfyZpvlmBgdA+TX4I5JCaHVYb2W/U9RUUMF+VfBOnmQSRQs7GPqqpIcS5
dgH9ucHMrsrLxuAwPC2o0x9UoEh11ilwN9FHmJGQQriu1zwZx97Ag584WipPA7vvx/B6wz6j6hf4
dlyxq33nI4AC+a7RKJFbPNSrPVd/mLHGgmXToqPZ60mjf4/WRMLeKb0l+Qdnnns21JtyGpxHUZVw
QdhTI9uS/grin5Iuq9N1rcr7uTdZg4knatduAED5caLSxw7wXDSeS0h/gORloinFONWbS22bp9t4
vpD8VDgKd6P5U0JPTMywlcem2h8qEWHT8QL0FCtG40EM7v4u1v5MbHioKfmX1gin0ravyEoyldhy
tgWKVKwoLqBgV7D699X8UVH2qSJbA3mutogQWrVTlb4kQkRNJLPECbWVVsktGzj+Pg7a6N/zQ0d7
5DfbmOZkVVx9Yy4JKImNognTaNuoFR8lpRvy7ckCSpdoU7ABM8AzClauoH1K5YKAMT41yBGB6QFa
ZBVOpZe+XzxpVUBwoVepqssbo1WxBSeXf5yX6Y0CdjlROyB9DDl973046ZpTwTyMh6C/xhIGm9/1
6pGwPgjwD4qnxY7cfFaHv7vsqMTCpgkgWiJa/7b+jGj6bOSEnL2fid04HYus45c963CHwq8fBdWs
Q6VlxDPG4cNcvJa/Br/O8n0GHGpbcgXm4NpE0zERNl/IaaP5KJYXs2lCKVxFQG6/F5xX3mVA9ovb
8z9Q5pXYWVc9iPAaxM5O9bLI5mWgrrEnEf7n/I7v5uFcL7CMurkUCNGFflyfiALMaHWK3V2b1lAH
/o8sgQ1WBmfVEapffcwl7+x3n24qrw+qMsUd9CK+/xupdKGkZ7GECRl3Xk/u7JvPIoyuMyiL85Cs
3ENBBHUVcjYtC725twH4MS2uCbFZimHaGXghfG38g1TvagT752eu5MC8G1BoT3nYmtx2z7L20HbT
OA5k2MBLvENNuv93Q+c6qHgtFgmCRYotWIRyOqJpZPGq5okckUaOfOX+mQNyGRSZMeUPSk8WWosA
kMau/OFFE9xoxj5txPZHGiH3Npe5TgT87FqftcELjcB4G8OGRzNdLEK3TsWdqsdtgpB0eexFR122
kAgz7nKRd4su99+3wGCVdt3kwWdYsrebQC0gTZJKwUWzDPwUrBOExzJzdv3mFDSbSshD3AmR6LJY
xm6j/dJ2lDxup+l+1SnmdlE/3xAXooqYj7OpceOQlNSmjQ58Sw8W0bv7SGbIyUzrR8xKRfNXhK+W
Q8HKhRY6a3ytTHnbYaBUgEis6vATWyaS2ZvjdlWbDI1k84DUCP+BzvuG3Y0NGgYvEjv7B6/XBieC
b/MQliyinVFb6QUkYno1F9SLGp9blK1jFgeJiqpvj0jUJt80ssDWBvf2/HdbZVklQqYLa2uStFF7
o66TtC05Wg6JlNiDItF8UkD0pnY50vthML/YYkoFX+aKoM+YZeB4eWz6E22uwO24r5N5a5hFFew9
4g3Eg/YFpw/GK7S32TKPx4feyOs+bj95gofNbB12x2sst14qo32ERuj9+x4cnxISV9J2m7DY4ive
sls1KQqD2T5GEZ3MbtzIl1bK7uNqBYJn5j7j1yCMZ2kJngc2EEwEtXXfiCMjV7UC9mag/FJzUDrn
mlVgV2lQIQ4slwRDo4FFIzTCMZ1JfzipDCoqE3qnqLewrjuipBO/tftFvHwKAY4GjKFGxWIRzSRq
8TYJsMWZGWk+PgV2o4Lj9adW3+Oo5ZlG1q6oZuBuN0FgB1Pn251nv4BMGU7tYRRM0jeBrbjZE0fc
Grs9gPTsMOf1BKl3+kuvo15NRN+94omEkDtzVLGgXCKSWsxAzP8xQpqLWNWPurPbH38v+drdgva3
085b15cQDUUJesQab4VpMd1Lb3+kZQXxxj7q7rOR0aRM0bV6F1M41krlvfNesMTqiEQdsKhchPrr
Ggt60jUTUBBlCakO5n4r6Lf9V/1P4lJJYaCFgAgC7nvoIOv/N2bs0DYI4jaVTW07wOLQiWzmxADB
E32EHGvBcKcoTEUPaN/UzBOg6j9GaZtsM1kJvsx2bJGji+H3+QrUnbnCWuyUtTkIcNoBt9VDi7M7
aRie5zW8WLUrahd0E1/3vX8MtIW/5fdhj3j6jvkn2l5VRiMv1dLSuIX+gV8nAA/JvstXMMCVxIae
FlRH3Wv32hDE9S0ojIpqiXtWkDSCb3fs+acajJY2M2g0WaClOJLfOpUTJNDyMbaWgBI9ReixTzGJ
wVcj+4mCb0CpBtAUrK82aI76x2vATc319VVKGwbdOvQ9kJdcVktkKB77P5w8gn5gldf6X8bBHe0d
e0GwdEuyIaQB94B1mkIVb0wJjyRzpD2bN90V5iV6UXV+Vo1mo+MY9IzXews5cpXc6sueALcx86gr
yCT5KbU5foGmEafC279Mth/iJTzNjC/cP+01+ipOp0J1Xn5VQlyTb+/q/fXeOO0JKdWggZLtJ86f
llfy7i6g555ZusXpQbWz204xiCXZMvZleZtiFVHiH/7K/E8MJQdaIMQLqcVQ3ESYE3bFKey4KaUY
wfBRMgEWjKsbgarsr3MGJ92bcXXP67DfZbz9V1L9ff3UilSK/cX8prb1ZDM6HQvfN4i3STtuAzTc
vlgy238awT4srDd947G1fRX8Ou06YrvH/34kCpCB6ZK8GEY3X4kqjUL0u9EgZNEXejlytd4q0Tkv
iWFvPvTn/0RXfSH0KzpXOFCmqQzVFYPvb9Uc/AX+/7fslrWxd+JdBTL3VTFIJlq2qwLJWPGldpUr
JrMSYIB38SwFdT6p/sy1XwLu1e7/i3Bg3Eq09eLJ/rMEL7zGBae83KNeOYAeOoNsiSFT5T8GyjJu
FpLani+JwmN9rTt5L09OFwLVXz9KVYMlvGxx3B6qN+iP1jK9YRIlR9NPzPml8FUQW9jid/fVlBo0
yLK/JFMtH0y802CTm9h+oNV6N1ZiNQjanzVnvL5gil07XPaPmPYoiACVl71NwvV2zM64wpPLOiCy
cagsuNq8siOoGedB5DXGGwC165uBeakBnSxHgCtaEA8wyR5cRtrP098dwmofSWbNbbllCHBX/gkx
9j96P0Xq1tq/QWAgJeG3Ux/kpksHAOfvaPAnUR+C4E8bxnf/fvbFvN5rWkXb4s/FQZTsPbRT7ppE
6bQwDwlCbyArrmKo25CG3sud7nAX5iO0VeaX/9BeXEH950+JU362oTYOeB7oSPwLNoiMZUEfn+NY
hJqDfpwjomAQkllsr9ybGTxJWS5oaIVesnK8IgRZ7c34SiJUEP+c1gZYRptgVASXUJQ89tAhSFWE
FkZSAYiAGH6xeJ2K/80s/ncI0eKxG51OuKNb7WGzI7m60IybOd9FGZGv++Afdj5tiMeDHbPNoQXs
s4BYTgcOheS0j0jY9fh7zoVYCqg0vDR1TgwClvLK6JKK7h+bB1cw5rX866A9dUAyPeWWSAidfm6n
z9yCzsj3rclV/9K+erXkQz0SKAGlNPCAHe2tVXI+aVfXsgzsIDnt3k13j6odFgOuKBReYWuvhR6s
hLTxfNyei8dLht6vtnXFneQ9cQeLOW0FpeiMtJXvmP0NAGO9HupKzaMxthx0E8CMMOApKYKJr+32
6X6PTrYGhOsQOvBOryiaD0F/aTiaVwm+JQoiICZ5sqdGCKTzGLeT3NFL7sFhpl2YXR8cO/pZTBJU
qIs3wWNTFBQeApMq2kPd3fJDMvQqC7vgWb3//durZKBNU4ZlI3P3rhNK8eZPTR+jVf5Gw+/dU6pX
z3uhUINDrdpskAo3PY5gUbMt3eW9soPyNJ+Yf2/w0xFQB5+TeDPJAXSAlJK+Y8bURrmBrfZ5F+lh
gj/9IW5mEHM7YuGDhZa5I8n5uwTaAYRKgzTvoeMzeSvvI4G9LqPxF1iagzTFRru7SItSZH9x2nDl
tq0ULTmEoRGkg+NXLPj0AdVnLQuagm1nGbs+rvXXo3XSQB4b+hoZkycgs29EBn01iCTVq/OCcVSx
dYxUQNyKacobV4Cb1eqljFe+xjdfzeeaQXOxaqkWXGjfCc/xfCufHmSUml8VhOrK4NLtT1y/fIDR
ExoXXH1Ur7uIUSjdS7oEIgEWaDg4ph4+2iWQ8FieRaDDqBhs4UayQdDz1QDYeeFWumELtuxCuMAH
Gs7Si7CxVGDawIBj8Iv0uAktqtvQ4mFoN/a7NGNXy77rLhj+BwaB4VdEoQIdbGSoLB4zNkTO8ko/
zOahxBentHdeYpjf17qOx0BWEw5gG6U6lzGzb3fIEJsdmV9sokOpPUOxFc21+ai5lmZGucEyplnO
gZ8ao+QMvfe7f/VwqJl/oUZUdRx2hkXSkcSW4InWiBO4FrGK6hEyBbjdAZx8k3nT6WEwICDfq/Qs
Jb8rNZTN675Gvvf9wOPW+T4uWjcYyi3fAIt9aqoeFF/EhBodCX1Fo0+70UEMCM4vK91oX16C6nd6
1izJ0Abra/k/XY/9aae0eiUfG7WbdRuS/Q84CMFWTT3pwGmPT/YmkHZuapuGrjS4DaL+qYkzdeG7
PTFzUWba4E86gesq5Rxna5F4wHz+MwfqDE3HJAGYXpKa9GL2UBgZuXs1Z/GINO6xfgXZgZ6kO2qG
f+SgXZYK1JorQ6fO1tAuIst18KUgIgBsSsDnf1v4F59MCARe64YeI5olW5+7qsASyNm9Cks76OdZ
mrpzRNtUBfV2aGjYonIHRabjrBfyRbN9l2KUvefJzSg66H5lHBpcxEI+xuFRoBEzQCiNSiDtI2xH
fooSWo46U9C7cbVFnrQG41gXn+Q933Jq+1Xw3pUB/RPbEpaus3J5FscK+CwR6y2d4zCAOMMVYvr3
uu4m6YA8KPen+OrhfsBNO+2d6+eHYYAyMTdl8gSWlKntwh0wSQSitwOWPpHPt91gw8gz9rKG6qDL
4EBZOrmG05DAElcRFG1w8LsL8p0RGUgVb7Vd2kFKeDueseCun6UbM6oxPM/+eSopCL+u/eTm7GA3
QHdCPWX3/9NxFTMrQ4MQoghHFJvKSJZB+FE1S9hWi88QqU7izUm44pVht7c9e4hsz02jJ4HoQ4lF
aNWG+gbSe6jWbculVR9cm3A0fls4KIutqFT24ZpVvQk60gHv3rBwyNgRg0hjhGnQAgFL/f8MkTbv
qDrGaJRapk1CmuZ+kUHYai7sSv428TmKBkt5DRMIpS5O6O5SOEEdwroTUwP7M9buzmZ7iEXMpMxf
svZTxE6W9lbi5ucSc+lQ0WMeYSLELxduqaUiLqIXgQIqFs5VGWc8PIez5RxgdZBme8zXD2Zh8TfT
yt/DnX64OrVGNt0taT3+qkbjXp93fd2HX1ykex5yxgfM9vBEQ+vsEnfDg56UjzYvObJNm+AJ0vbF
6IhWMIi2ZcQMVBwapFA1AKxXDViQhzizVoOvNEDOTuM8IRDkRVS4G0YqxBAWOThImX2bcOZZhvtN
7VpKmYI2gtbnG6HjSwsgTiTojteDKXoF6Zl64/GupecG6SJdoxSF5VG9BDUBQeViiDeUNjtSJs57
aTKWo9bDdF6xZtIHwJE4IavvgBN+lqv04VjiOPJo6Zt0YOj0AA6r5Rqs/ixDERgYtYw2v1pz9k2W
Di6c0P/3pW7mSK4LhWHFQK0kOyEVVbhH715V1iestZim2nUkBNuWzkknFlw0G6OtewaNn2m6d4Zf
g1FYooC0RjomNpCOw71Az8EOm76u7tXnxsFLRI3B4Frjm+LMwWIpCvOj00h9XCeViOTbei9VyM9x
Z2C0i1VDUKzwcag+Z1K3RdYmVFmson27JmBJMXXmCwRCW34TbWkxswxSHhqt5k8QIbNQs+gfNidM
VHtjR2VwC73d9OAyfkQAbGKX3wHj0iT00x26c2Neb6omR6wLaXilJgvbNx6OPYlTZ4p+n++MnIuJ
bMDg90Hyo9OxHJ1yh0bOJjsNReDpgFABBlWCDpJf4EyD0xaqeKcU0wPwmN2kWKYEpbEF3sFbTWI1
2QiT58FlU26r2DLO241ha8MYfFrIKq9UsNHTkEaTVvMr9io/t9ZleDrLgnw/PFojNS43COICTk4u
8q5BXL0iv2L52pirPs+hiJs+I3WU1goqLhAfNdwYgO6ut2G/gBhwoRPhs/GyEdxtWJc1rSzuOTnR
PUSDY58sWJZmHCQ+FnGh6I7o1CkPOurOKzSfU45yvbQCU2PySfCfSNZPp9QIGEfTqWbyWzbGtawG
zNSi17i8CZ4cC08sR15PgLdIF/uS+ypGU4Tj1o+wxbrIX9laFznRPULZGgFO6k6R/bilTHQ90w3Z
XZKd0uhN3ZCo8XMVzZ26h4UN1Z+qBvwHb7PWXErixxL2IUPtHlO5N56qJcxvMAvO8HMBKlrBDs3q
srBNp44liP0w0qYek3nOvlbBkYju2QRsmuFDK2ko8XGo1pLwZOuTxTJzHaiM50vaZkshSL0oUbS4
XRZ/3DgB6Q67NrZ1wdxQUvNKjeyQQYq3HQl2K8n3WkJvKLT0U5OJAz182jILwiW1tUEElTPmsqDS
33NbuzAzcy5yhkZe/UpmTJs3dS34paCr9463/5QeuJOsz9p8V+sc9LIK0CZZ90CLKmCuW8fnVaSM
kd1mAu/02YdMJKWUPxsTdQILsUNESBZNLBULW8X8gBVDoB0zeMQeUSmE125l4JPVT1Jw1BI6MuTj
BN/ghMS0gHPoVpq/2NwgxlGlo0J3zEWpH4+ntkJZH+xmnBcIrt3eVJmI+/XwJZUbWOa2QBOQEtpG
8J5G8E8r9X6eJ5swM2e9/nmnV7KLxBmqXKGZAKYyIygFXW7shrlEEfS4j8vLM+OvyhOyXgeqzzXe
4DyA+yaHu+mepHVHRvP1ZDzecY2enoV6SYBozAokKra4TW04+Hb+GaUzvLkoccfAZsWstDHx7Gla
GHcb9LJHfVeV6yoSp5pDKUDroL/2hOscdvKAWLix82NZPSoDKgbDKDsisuw3pptI5MkI0ObOiswx
hF7g624i+Kc+KLpjn2D7Bq5EuQ1iAbR5iISdoc4xIkVbkGIXBBlXm8YiC/7EVx1kTvFo8AVwEP5K
/qOxsbhIJnz+8iPjMdx5ugBSPbQ2lpef6Ym62nfqDnHs3HmBnqmVdnABg9L1KZmjhswa1rtyonEs
s0lsnRUIYluT79/ZCl+erzbCVZFj0+gcgx3x/QWeG+KliRWNq4fyq1U3zPqILUOT8WkNtDNq7QxW
AHfr99P72g+13461qx1064/Xxy/am2gYoEghoOq2iBq3Cc6XxZuw63f/eJmsFnm41bFrEpSociH7
WnjgN/+I62uDij6xcGitAleT1brl5hzG+bbPYZ58YKnHq7mnAcTIHwIdrThns10TDfU7ZYeFXf76
MIkPrvY+RWI2Kv/V9WU/0kjEadvFmt7KPEv7tcsv3leuNg76XkkSqoUD8nHOh+96pqUT6seZknwG
3QNLuFegQcV+szPkhrn5xJFKNWTxdA5YkgGyUHkz6AJlfe/ynNpE1XFRyZT/1xw8WS9sw764Kzvr
g5t0EFMHWWKtCmK0G8T5aZs/HsEC/fUTC0PW3y27Zqq3c1qKt+o4+NpYlNfyBCPmxiFLZbJe+XM5
6zMVEGluCufvuG2xlaHnY1RsQXhd3HIBGZh6yuwzL7xQyNLneoeMp7sKiRISWMbOC/GOEyeBg29A
9kHPBh5SCA8DyWJAZTMhlo4kCyTrYUfAAIT5UqHmjxH4w6V4nXAJscdYyIDHe2B6FbuyOyUwsFQj
+cLrFRyAqELm9Ey1ouW2J56/yNhRJU/OCU7bts+6LAn+0sWS3iOLPWA6Uwz44b9iOWQcCpBdlevM
3cNhCmXe1rPfB+qCWOOzQtFG1zAhOhcw7KGuwsMZ9dsWz5BE1z9kEoW6XkhPIodSFPMCabHgx+au
47veS2LRLKr4z2rydB5qf03uH4bXsjYZx2oMu+MLrdXU9+6QUMvMLAC1jHRB4JRLQuZ+BS08i8ma
6QSCQOL5K5VDIwdaCkHYeOppjl0CsFMTEdGWbW1YkiT9VRqqvFms720O2QmHjbLtRTGR7qrciyn2
8RvQGRdBsD23YNnYkTffnECrLC6P171QqMin519C8YGA/dRhP/233sZ4ul/8Iw85uYrMvF41mqnx
x07QxJKtgJw6xuzCVQ==
`pragma protect end_protected
