// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:19 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FgqLwzOINqL59I0i6227/L4hixgzSlSDtqg9b1DSoisJxy5SkxFQ6YJzI+U8EZ0d
/IwrYD9mOaAiMHQLFL+0rVA3hYO1Gw6/qOLjaH6TBU2yvOKGz47w0eWzz4qcRm+r
ZvZJlCbs6E4H8xZ9epQUdBWU6BmfyOJgJCaWIEKZnOk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12128)
5023J1wBGTEzVtDVgLZaaRVqpNc18YVWHaI5EI2j+Y+m2xj+Lr+1SjZeqHzqOKea
d9zrquuBqv0aGIVX3+h8ZP8B+nnCCWE2IZgfNKOAdqZ06U7Ez/Pbdx4MUEIG6UIn
vPndc04/2GqqoKLEdZsT266703bIOGNWxRAklIUxp1ieOL36e1ZG/JD4OvZqUGte
+AXhOPFhV+V5xZy9WksWeyLMBB0HFWDM3pcCg/qRNClrjgqXNXjZWW7JbaplsQO4
3SqYLevVj/uqJuNPIfU4xFq96WI6Fl33mUEg03HsiyTcyxzGFsgfvxlUbIfOsNgb
YeAFjndPnxcajEOG/xFpv6tPcJ7+9i7g23Tq/RFNlXekmULOvCY6eYG944zLRPd+
usJ6VUHrYV7b3l7bXqlknX3Nyt8joMzqt1dLtvQIYYNyqE77SYYIcfzPiYbVayUv
pkdGwiX9aajoHuvrRoFNuG/utn8+xQZengfgWm/DAC9Jj5dooR+/cjoIqCcswYbZ
8FbCnc20GilpeYc3klLiQAh84JcTnGdLg1SYXFDz8fPQoGdiHc4R7lq8pXt0m+Ua
ZMhbBWFX0tFBV3CCZ1VcyHrGaAbaQudHQsOvrgge4uWwLz8I9rTz8fDfB856125U
rvok+TtB4QA8RAm3c0wJnSVnoh7WGxhIoPJOL+J3X3soJs+R7YIHcSnaFATNcxE8
HfpNAPyntIcKWlAw58ZfP0n7QUmjiO4eNXtuAu9vVBI9z98qSPwoFJ+Rr7lb2Azi
Q2cU+BOPEtG1kg9rxIQspFuWptuLHfDbHMljKIzZckLZ9sSRrmbS38PYTvXoUyGw
PfMKMOb/knM65KD9Xe+gPCGi4Pz9LPQ9wQ34knZuqNxkIH8S5WxjGPUqB4XB+b0Y
v2rAVpC3FyuS/lpblF6I6jYwReF4j2HC6KS+M2xg4A/s/IiYmcad5GGeThfTzf+K
WkVNlEPsSj1QG2mjoUK7oIZ2mPLyLytRxs/rR+CrQrQt0wMTL2s1cjQOPU56Mj/z
P9r/wHoyyKjMvsSyEfKAklhgKYQPpsAn6hA9sZgLQGLvjRoixTFvMVUJv+vdFVHt
B9nPsCxHK7VYHfIkWXaqKiZYT2MmZ2RzvcauisATJzy2BDpWOaZXG1xFMAgVDpzG
ltHq7ucAC6uYRFWrdx1XYaFiPLYdfxpZNCciWZSN4CJdAmIV7LLYZX6u4i2oKg6u
C8E34the1VrK0omyr+NDg8n+qkeFpufrVe2f+Av/VR8rJd2Y4c7SNhD5AK/Hddvg
v+CXdg/iV2eA++MUHCHPOWTMdSOJArdvvgEj128h6uN3Eiu6dvgeh49DGHBu8Bq9
VjSkwy5rgPjLg+9NGsIDVFLrRRBPsGNMlrxQ+OOeF6dk1CBPdz+lLngntDMDB8Te
jgk/tDBoPZ5AqD1vDjkFiOBE6m+9Cmn5+Y0FUvFxqXHdl9sfeFWVCqy9NTt9dt8J
5I7OhfKNeAqMxWL4HGENu7UXFjF9Ywg/8SG04VJY73E1faa4dmgj/KaKBVM+NWis
sEKfotlcOtPphaiWkephNPKfwfB5+fz74N/g+w91lOhDYgA749cH/+YAkwd6iPIZ
4U8at8xoPDd7WZm2caBCcbAEkw4nqfajUve79hXs1HyXPWtqj9ghugh9Lau3Lmt/
+vUY8CyI14g8zBBvtYkK/4OL6UB+dfi6GmQVNhr+sFHfadJ8sHza463c67IV+KJy
x3F/Onzm8yDs+BzeFZVUnl6xfQiYQbAv3zhEBwkXNuEDnDqMP762JBJFOs/XXLeV
YmKaUIS5hEaf5FQXWb+J80KfWgTvBd+e0+NzLNAaJrnCzyZa/ymiIR3mFGMYqgiU
eMeQFBRpWahdNi82BxryrmNSL4kPXDdcPBUE7xvM37SUIrDGylevJPhFnZX3ba7j
wOHffUnbT9vd36pI6EvkoIRye9duGSB4MohCwC+9+5nHyErNK2Dhls5iyiDl0b8T
tUoOlqIwIFCZ7El5JOy9ID33G3LpAFZXlPgQnnCzSdXbobZtNHRQDk7RZXyDPyz4
TMU5ZXm9y9xAjj+N30P3jIUFxcdbi9btChzVR1FaMWj7o9ookeRvCbe/NEHW7i10
nJjxCylq2220HrhzmGSQvmxpDeL0D9pFgXoYll/5pcpMbGVew81iKQpTq89j6za4
2UnbHvx5Ok80ISpGPnt72VdEFIIbuQn9nfNcNb5Usk/xhYUdrrqniWMAWBzRQO1a
pSrzaiLqkXSniEFguUd3MHdOuhXfrNYnaMHg6yoruS2Bi3uyjhZFpySQhcbxsZtn
VKTRj5WL2OgbDIbNjb39kNLjMjzyP86o0dxMO3TjT7zMoPbDmT6+7Qutjculz0y/
AjPWW/D/NepR4juxKZZDz2qQf2F0Vgh9scHIzArJsSo6OJz0Y2FLGgNZGfNH9Ldr
zZqgpG/MJBh3FSFG+C84ZD+qpWU0QlrACRl2mg/5k1OaEhgmzm4yGH8oYT1SlRs/
f34myqAjPmZiLABSTbvDZa/k6EtTszgeI/35n0tJw9I1LFQBepi+cL76twL1zzBR
I6/OF0V2jQQ76//FdXntiPttz8R4N8WHcTEQ519PUHtiDNwP3zCy6HeZLvwd/8Py
hboTC3SyKSb2EryVqbqvzlCZYIxjSdCK7iMb1semNNSVJuRlUGRsH160VF51fxS8
+dHRIxDFpziPVgtsxVCVbgoEzxfS8HOHEKNUFXWZH6piHgacdhFRPd6GHYWEv+Sw
0XCOd7fsTA363j/GrXSAngN7BIXxUvQs6mTWZCZpNTLB2WKlKIvAz462b8LmHGBA
eWCs4aTMzX+neqDIYSAxMh81sAWjc1kVQhaZnTMw+hOXMKHZ09ssCWRBwM1dvSiQ
duJSnPdJmRc7jZhsVpcTZmv6Ugtcw047krn5M9vA0XpBi8wBF0jNnSjKaVUbAV16
bFXq/4A5SXNS1mud3Cw3o1XE38XTka+XJvQmO64gXl0xxqJa0eX3B9V5azcD9YTo
5h3C+wejP5Jg7ulK8LswNw5rWuFjo3gCLsasI5ZwfdXUFsIna8JQ1p6UfOTe0N8j
DjBSqt1Ph9lWGwfFMd3xRhH6uqxIaRhR9n+Ar0MXRq3EXGiCO6jOsWX3QvCcs91A
35qJ/shgVjv23wvQUZSewmB1K4MdLe3VuSainT9/YhMs0oAD+Vy0QMqmmfFA9Y4U
LwFPuT9sOIfg89I2+XZCJscvxyYZpO+oBQJwSoU9K9SfsTClN0kzhaKSbNuyYcaZ
UhFUypBX66mL91qiXTwFlvki8jFEWR6i3EF+urzqVsMiqeuOfm1XVFDzaN2XlMhL
a9lWX9/pzAeGeUycNLZbGtmkzLLo+pme2j8Rga0YYvMoEkRkAFegghurxbY4x6xy
cZDKtAES36kPzcQIhWd4NlxWb7SkYIwCS8Ax5GLGE9CsKUmZ0EVEIiBbMavSpSK4
3m9iL8BqyK4/z49Lu11iTWbd/1WPYH+lR9Qo4OLhHJe65fgJKE0XL4bmudT92OjT
mh1G0U9AmjaJzI70v/Sz2BWVtV32mNWYyTTtViQg27pA/kZvgvaC+SHqo3P37K9v
XaE1Wy/iudUjgC9mIcteAWOPsvF4kmE6cSGp3G6ySibE6MZNMlIf/UVy2azxyMZQ
/seUKrT+neZEgA1VMuq7o9oF/hfCoHPeyIyxptPJvMXNlmjy7UFtcFvLhQvIeH9x
Sz2u/p+iKhZdQCGQSIgK9ajdZYNrVtaBy+R2sPvhcvbzB/RdP8H1a5dbM7oZLjWN
4si0dEzDOALf8U/bHSnQM6XGqhFrO60XPFMMuCFJga+013ygA/rYV7g+U+PhvNKU
QUWzKr3HHte1m2wf/oglq7ZvgSl1EGBz8g1dxTJWKpZfdSga1TeBXuTX1FpuO93T
vFQHmQOE3hCu5PYQ3em2yRIy2QuTXAUmENkhqGzLZKu6Ph5l6sA3SXCrMqtNdjgu
vxSdQt8IW0teGEazgfNdCjN+EA6SYrdGgHswa1CuSjgFu6vmqgDioKCRYK6kt5NN
hHudx6r/8jBXIMQDrMe0jwut0iAWfK2SXrNOKbwnq3SrQfoAy3cww8ebgbdeWaoI
avmJyHo/IFaZZGo01UnIzUOcozzMMJfQPEiIbiaUjX28G7b5qa5kkceSEqbeSkLv
1ouE4/YX+fcSdd2fK1/wTHYoKUHqKL7bdNKXTvuTA+SbRb8oLV0Hz3u3AvCN/tbP
Ik7uHTX42Rt7cDhB1+kf9e51Jh7ZGy7A4XfnG4JsCiB2NjdoomXM89PwDo3CrqGh
gDitVXO8uC5tzpxHfNP5jODvt8NZ5BtsVpm4awIgGUJmYWG8QQ3KwthUmzle2U4X
sw5xBUBSDdVhyqNQixVtZSzPeQJRlr1jIdatnAIi7XYebeuLg5FwsXb8ZV6tvWHm
YS0WF3aLNyIuT165GTHsk8N6T95BOo6VKsI6aTcAdxXfth5Zoj2l4SUZrHJYh48h
gFbfg85VCjenWgV8bgqiZa2Yx9H7gU7UcmvZ/EnaR+1p9ImSE7AX27KQdjGH8F+7
bW9yd2wuufZCON8Tmboh0z7OfbLUUzmgcmQn8j+CcqU9sFhfJPuHuUC9C+P1MK57
86tS9iSpwn77aRhwjWGVRsbkqNxVLPtekmuXWvV5/f5SNq8KSBC4tgx/W5BGv/Vs
xfu6qwv7NirE0rGT26cZad/VG7kidAs9XblKeWeAHOSMG+HhD3tc6RdYSVmVSuTF
EqbsD8sjlXo9hfXYkMJyEBvvR0r9FmGdmhXMav/m/1urM3UGz172xh+znQ6uEcs9
3Wu8LmrCZfSn1GuXAc7sRczsq3YpivzGEejlSEr8vmGlJFPcEWHliUYPiaA8tAzm
JrDAOF2sNgAYes6RDJ+U+sb8Pt5GzacJ0FsgUExKMa84mQZLdO273i2RpKr90DU/
wLQN9lJxNH8pp2mzoX6eabwkXriuDnVDLaEEjOz81UYzYKm+R95Tfb2vejiYavTC
RyxmzewZRWx/hG3XwBDDAyt+PCuGN6TY122fASlzmrI648imLTGqsciLdzAsTlU5
nDDjB5lIXBlNb1FxeStgzTLygQQE54TdgbM6QSlYtFgSBqHCiul0LMXiFRDYznGo
GmMUe4LXPKluNl54Ka5GgwOEWzjQCxIVTSiemykaA6cpRKSquhwp5ZIat3VwC102
w4ZXQbxaLcTwNri0mTIlP0eZSRD059sQ5UPH3alELBa2hhdafeMbhK9X2L4DsG/1
1oCYp6fOkNelxTlVD9VfVlfsR5DMqVNHrSXgxmU2bAvvcxSTM46x3sahGpzvFMvM
tNDJhfrmukx57Sqm8nlfJ/Lq+o9dfu2xjTPV0uqSM/Br3uNzYHf/R32svmmNni1q
qLDStoQwkNOWnZMVLJ2zKQVIyqnA858mrxFPwUb5wiPOvYnAK0aBueeN41PpQi33
7pIrRpF40WIVZ5EzKCvb3HxlMcsCiJH30P5MVFSnlLMVrOkVfARmb7HjaEEX2Kf7
Qk+mD5dLN4GGoQPKxL9YA3t1plqFNPrBuhZmrIfyMbBeumJUlW6hdxW+MOys4UZJ
J4ExPo/mv66Pltm0/6Xi1fnT1jKsnrQXH90zCKWU7SSt57B5S6/lBxxt1jvlM4qU
9DBbFqcb6lrGGcV3G90taDERb1AonHPM10aC/OB2Zyb0lFi3FYbyHR3f6bTipt5F
SNglSQYKLnFO/GVHDjjHzqZP12GmW3D7qLgLFQ4URGVS8dsGyKZEnwjrDIFnXD2T
gkPIYjTxB3REXOhKr1IQKAkeBQuHjnsAnBgiCRXeZ8g6Vb7z4xx/v6gYBm/9qjtl
8XoaTzd+u1Uzt0i7vuHmjVuMWTPtz39VMoZCzixMYtR3BbFK1e+OtwypFXsR2L8x
VJgYmxmzjTcNpR1i/7uK0xE9NpBIIuQleeNgeRX9LiWdN21l8NvPjgMNyhiRuN2b
oNjQwgHXlT1AooWERrmtgZeUKfWoKs4vMbJK+796Q8XESHazTqccAhvXbqKcaXxU
666phWwty7hxtoFE61ACwGO7pnnF3kfC5Lz544xZ+yIOT9dF/2Ry69J2nRhwnDGt
AqEp832bUVzGG4pFiL352EEGOCJ7DDCg/OIuWbS0fQsZq9ehJfKFSsrCeB+My8rF
ZYONRe9aESG05awkLQmb1wqGeBPGYPm4pmldadOG256ZoS4LSiuocM1LkVa3gmO/
S6v4tPhCGcX4+O3WFDuRR4E0negLZId8Cy5LmvKp45eYIXyuzWt+yn3smLQ/RteS
IXzoHqA2gVu6G9zffomF+CvqfVPSriIEZQplMnhgPrLn/OlNi+Crp4UUwItrzHQg
3wpVVDB/kKP/e9o87tvH9T+df3qNPnx/fG9LUXZLb/8HKu8yM8JTPWwmTnYwTjBU
QOQMpYwjNI+vhtX24Rwdkmi12KunftCGb7m+dVRQHmt7soF+8vG3vxEV3LIhHwql
UK7kbh+BmQHDa+VdT14Sef9RZsdiPHdn1yTGLwrQtEKiu6PwsPeAA97ZhTe/8TX/
92KJar0uUSBLFM8o3q7W6VXRiH6QtqQahw9x9v/L0/kRgvMGsQ/UkgMtBNvm4Lj1
lh9nI+kt/pMFsYYbzpeuBbbZOTb8otvCeVVz6/14ZyIART396e0gWGroWHdV25NX
GALtE5sy2jU4cQDoaleqTqggi1e1lFmW4D/IMsw9M8NRVsqPvcFLNI+7rqhybchM
IOyae6aQzGyo+2UVu2pmYbWMI6/C7Figmfk3yUsulGyq32Neq+5ZFzyiKBiMTWnt
bBSgl2hSdg687Jk3HaN1itMH0jIMdSD9ZETJoCPFVGLR0QsvZJgdm2G+NxtEEIh/
hb8aBFhV8VpsDIOc+tZWX7EGnn/g5OKFJZbA6dk+sDGG+aofOBHBPOqW9tP/mlst
4elrkSdwCTpD43Oy9jDO/lXEwkXO3/YlHq3Xdg0nIyqcVGgyWU0ZnNFbLajNQ28A
UES62FaeyYydp0oyvp8xkrGu4+rALaUMvxBZz+hrPHzS3oOuICXKGEa8J4b4kE02
ojER5rHUKvKEdM6gbbLAm9w6azSUYZOh48cJe2HyKXh9U3lcqf1dinevAedICzEE
s0akeERLPD1y6yR5DHSdYvhJkdJ06NvU+d3Pr17LI2ygg79oDmXi1LkzaiyEdwtC
dQsN8ZgUxU8vtXdamOSXq2w90DWPDlQizmZu1GheqPDq/ahLGsGctXHPc72fdjBV
hOcG6knN6vpsZxtCqoonmdURJupTmpV7H3cHhhJXG5b8059kwhaUDXiXgzM1nvXi
3cHSZUgHme6GqXPfPmyKR3hDrVw59TUxflpHFli8O/MrPiNuCwEuP0ISPgZkVbS3
32a6gKUsZwJcQEjBfxHcdNw0ut7jgoK8o4F9FG9iTaHHKeIjsjAEPgoZlaq2i4/B
pegQXtwPQRrJE/54KRylMOy8v0AG+KCI4V6UhB5sjTDzomb319thnT07zvAYEHTb
sItI7uEcHdqBtMl4FUkEH6O/dSLO/YoUMPU9BZiBTpA3MXxcZdRFwHYOczhMNIzW
HSGLltTyi9dhW1xRupmwNZ0gFotp6zTpeGppgz1bvI7a4pcsXZTJjWxdnYIahesc
j/IQ0xNkBvB5aQLQq3aCbI2Ebg70isHxBaC4ScoVm7RyTeP1rU5b6P+VmCgV8AWO
4vnvSbNsLwoqi669707m7vKPRKPWXi/lR/QMbBVrbbbhXut1HJqOU6zUOt3eDNFd
vp4Cj9fG1fai8kppw3LGiPdk6QxkgZwn9KcTN6jxOn+fiDeRkuQqXKOYZ4brpOkc
pxs2TjpXOZ+/WFm9ZMbQldtZb51bNBg9TUmd0Cr5URRruilJxuDg62pd9Z+zvMlj
cZ4c6NqRFGy8w2Vgdzg0kVoMlEl0UBeqDOxkPKJ0QZ/fjGvO3AytgVAhL0DJnXKo
uVUKAf9L3f3TzfGt8UUNzyuFXe25gXFi5oHfwAW2Q5yuKiedNKLEmtcE/febgTWd
gIZBht6d2vrwGCNOzAaD94RY5RnsEqxEYCW0Dje/hFzJ0niF3vx3NMKo+y+X1c5y
4RYo/1Fke/D6hxl2ApIKU/3kHPm29On1TUI3vRS3LVfpuFJTXeyBca77S63lUyFZ
8OVmncIyjs2IHBtPAl7rZ7W6TX5rukQwkVsFiC6utITTYBRA/vARyDufL7gos5Ik
JrGJFs6pH5DzVyccw3u4i4pCedciAbQPlYYB6dYNjaQzs+94WqBCNikRsxGLzisa
nhdJguCcUngGE7hqn+uYkj6ZwWeIoPl8Pc2Z1MItFvSSZIsntfHhkJ/amoYsIjkU
Rs4nB/ffXRa+0f866A5llHJn4334tIvWnOeRHsnNBAgKuWdeAZXXM8MByDOO9eOd
Pa8KlXQEF+49IHQiKV50IDA5s32SWC9N55Z0UxXmwbnXANnXBeZ0GjX6u9hIdgaI
QwDNhxTpILqkDxce8tsTA/zcT/xzchNJuwT8e2pUVCaVdQWcWZc7QqbYfBi9v5uN
HZspj9M/IgaNmPoiN2dUVrU7UDQLvtRfUVBZmpAG5pEfxCCCDr4M1gVUSnXl+63S
IBSOrZBCUDQsH679egzb+H3f8zRmZBOQ/A0dqUPqQ6f7sYzQZ80uHQigCFIf7GCo
hJ5oWv7tiZtudpVvDb1dt32ipfa2HxWiCmJc33WHXf4c6HaFmQtstJ2C4WNyO8K8
Hg4MQWVmc2SbE1dUSQMyyCFAGP/yBZ28mPxz9Hwz/3COQQ0W5cNZ9/g3hohvMQoq
XH57Okbsb4GS5KTtJbT1bAx4G5CPAPllKlJOd1qtbowGB8/Af932IeVxIhWAKNMp
TunbBXzr8pi62zM1tVUYiD0GhoGps5xZongqsshXLeAJ2cVTUCOE/nEFqsRqcWzV
uMTuBT8cRSLVSNHuc63+KQSitCnyIsB1FRSSu8TLp1FnG37qR5+Y1xx9ZqxQxj+5
EeyFdMp6gvIzoqKPi0b1E022kKNFvcHlo1m8b7axl+U6tSzNBGVqkM+wCT1FfUgx
h+ynauzzjnlgOpVZ/am5+WdUTFB6ftMw6uAjgr1yfuYKqy8KHeBbIAKepf0VQirW
aPR2I4DiuQSbNqVdhWOV7Wo0I1Dqtm71UTj6/hKMM2/3KMg2DopPaka4Mmy7xaXG
B10pBm+pwGhiKYIP8juZYtIu8RQLyxAmTwr9lWamxDL08ay3hVVjvPg08xCOw69x
gXd4cvRtweZIGr0z0bG67ntMfeYwfmdhFGX3TOcHay+OKKEMjWmPlZ/XF+73htfv
zrXbVZJcpIXHqs0bWfyKhmJcPU80+Zf9EfOgFH7aWbvn/avgWQVB7xlinVZKmPp5
5D5EspXFdhpBfdL5LZkO3s9USjn8tz3Uw4qVf43mXtQs9u9435mUKNe3EoJeDHrL
5Y1GCyQf0l75dpDJhmNLBSMG61onztQMUkv/RC0qOHbpfSXwnlOyDvhtHOZ+fF+Y
g4cp7ARCeBXIahp2vdQKObk5Lfk8EUOOeFYc4Szix0xprQodCwUYMDk3s+sYzcXt
tUttdein0eplWoB/e29suFfwbisUEYfzMzsjEmIycCDHSZQqbj2qAaDq11Es4Mg8
xYbgSJ1rgP+bSmNRJAN1UQk4QrIdY1Svt1oDkYVyU7kaSmUig5ecGriDj2cIHPG3
CxkIVJmpDgK0RDhd7fsvJJy3V6iSddfm9hB/YzC+1GowY2E31H1QHxXFJIKw9XBm
zK0WhJpslCBavmZ9Uv2rx/UO/Sk/ZtpFS4n5LBleJRJFfo5yZLvtKicRUVEKbofX
xK5woxjPyOo4GYKvfp77Q3QdrRWWPdnE177nF8MEft37U9A8XO+Yq4yZeBVVuS/2
WtxosR++7n5tJ0ijSFgi6VU7C4pw6H8oZMSazD7sxKSC8kV+Pzc5yxCd95qkbBKc
QLKQoeht428x6StL/1OErkO4MKLmZN+mYxFJXpkCQ53CJjOr4tIVaRk1a/JLFkLk
nauSAP3ARm1Pf/ut11ITyQXIZkHJRTM0FJUCYGIpiFMWmbFT3JnpeWa1jxH9e8uD
08ZTi73MdTB3f3vzOQhi0zadOIBked+R72nUvLEB/jPP7gPPSkSy/qi4iWJSqyjp
ZOZ4EcJOwpXxLj27tZk5srsuf4xAGzwrVXV9sY0AGo4GC0RasTiK5YJUowp0FNgB
jjuax5CeTbnBw/3f9GXKrWmDy+Rdk4M/b9QAmVtNVHhAkroz3EfMK4HhHNeM/Q0x
/Y3ET6QLoVDVV56kieihWZ8EHsF1WP0I1uMwL5iPSCThTpX4yyPibq9j66yd9aN6
XcBb9Bg6+jpPxonhAXEaagRDYEliEwkIsFPTSqI0wEx44qk203I8Gu+rBZ8GEjC4
HZld9ramxtbRJFB4MlHgxP7/UktE+sgmOadwsqkiKb9oWC72dZ5AOTxtuCBo+M7z
hzBCdy4dr6l8isrHkQZCFkDgYA3dUiVtXcJYbr0rBWJ6tnCDl5xN3qOZ+L2aVTXe
MF66PU3g0338JIhRISzBdSeupQEHsDFFle6BDiNhxm0ogXQL8MINyJi4KCzQhICH
62Q80jBbBfc2weEMwmz2pyoNeCNr8WZcv+ZoShAWDofu1ox1PuN9EM5TRmrUKBFy
qvzb1S5hubBLSxg1zScMymhPs4STe+UjyXLq4foioJGyFu0bADwmI0fjjHXjLAt+
RvteLZXCQWqs/VDJgwkAtJagQ1p37zfhPQd6jrioflrYbi6HOcS8cawjGk2Iwl7V
H3YV2azwOlESEiQulOfYF431U+WbOpU0MDl+zI/UYMzydJNNHrDtnk/LXqcAQMQ6
IXSHtEE1YTFQ7FvaL7I7Cc/ZJDBD2MbaYXXvGJQFfq93UNxsM1sKM7Y56Ic01wyb
J4vNcuhbKxoy2+lNocf6r4d9KHzzCLC4kyM0nGcfSYb6nwpC7LXXbzkmDH4NaZ5O
C6Obw/YELseueytFrAzxzVt8YiPdPceZRNqGZH9867Jl124iYmHLvqKOxR/fPdNi
lnaVsv/Fs5wg+X4WpDfTPOmgwt9j+ABlyP1fItBP3zyufyEh8GHlTmAKr7VscHPQ
n2gffUwalWMApdy5fIEdEWoFILWri1Ui1UKgnGfmo6+RZyehjoqLiR3PmACniBfr
P1sTqABYLKAv+lpVxo2SthtMqYyLGjCF2ZYBmdR3yAMoPHnsTu/3mVDJ5GkZsPR5
mBP3GnJBtAZZwtTxUd6KWaukYS9wBz0cjc43HKfxf5V+vlBF0DLmZ9Eqt06ZUPCl
E987CEg999uS6grzVGM5nui8BLItun17mL7/AJymC7Xr14RqtDZh5mbP4R0kBMiY
YrWMbQ3+RGQC0SG6L6pur2ANa2hItTeaqZCRtfVW4WTniNxx3wDFZ+uPVLAY8wg3
WwA/R1xTVhI2k1b6zq9FwBDrYhNGr04c16xTpsknf8IVB6U0rYlVwsn6nx+EYubA
kkS/tXL3b0R6VsBQUvaDdxkPPmBtXnMVmD7DIxBNOE28LWFCPb4S6cUxCNz24MVs
IGJBdHfGKUIByI5kA64IFI2zOAbNB6IldtxOon7ghwl9V8L+1xxYa0Jqfp51OGJL
VZAn10pSDinfq+JIKOOhfNMhFtgcDqFMGiUVrkLRKNhnZ92gun/rtDhv8wGybKD3
cjKRt0RWomnvu5RbB6SzbevNZAHgB8XTVN4fyQerLE1nSpGzZGNjfHlQz9oF6IiG
QJckZMEXhgEaavhP7Qwyu1JN4p3un+jjbd03QKo9VYuaV3bz9xbcYKBdoGGi1mOU
NDAVKkAa8SQjP4PfhnchFAOpjZ/QsNCiHuK2cMRj+98I3S7bRijiTNYDi4ZXzyEG
3AIrfUjgSF8pRnyGtiBUD1A1kzkvnN7Yp1BXwtUAJsytM620AG+72ui9YgegKt+x
7HI+vJKhc8bHt5jFB8DwCK0EL6ulIp9S3wqd7qhiQMANXrALxlp1hjgp46xoTGs/
ZFgTyGokGWZ1krG925LjJt5U8QHsbNJMI0RcpeuS1YGKLOHbsPw7pgAKrapHngAy
WO4X4dMOFEiwdx0OtbeN4XoRyBK018M69QtPwrZok/t/Flj8dAqPODu6Ox+q+SiM
JZRaX8nCpJhcAF58p7EVm1RI/U/GV/JOAH44UBNOBbPJ5QfCzxTgouQqH6x9K4Sg
2vJRFYqXnphQc6YKUsJgfmUkOp1YvYpO8I9ryDvzZJ1mKPBbHIVyezIy+CxitSvN
vwnpuRQhD1/w9uKzsZwiKgaOF5UerZJHm5hOox7G0LCS9HctlLn9f32fe1M1cO3D
hns8LVSA6XNGzhuNCKx68LBHe+dOsAGcvBNOCJ/fUTEDHJ38cw1IV5od94tcTUTl
nLkYyNC/a0fE9bUSnzgWGiDiwZUZen5baO5uxLeogHDhqhNlJ4G1L9C7hWriU6ba
PPVZG345txmYuRaoySE7C54RAOVW/jM5AXfR0Fk/s7898IlLLG9qX8BD+4jnsomL
1VEG82OhW8hmC2HqlVGIsOoDWVnIyE6dSEZ7cAenDr/ar1R0T4OxdTe70zdaU9nZ
m6qXy3vkcRh5PI1WJZEIQ2xrDs/eZ7dFoZ114Ee44tK22TuDh//MOGAtN34px0lx
AbgJDlT+9QaASYSUz0irVKxilHC1ZcEOsDNKzgIY+R/IR+d0UmvUwGcgZdjTYqS2
cN8q12rgtVhRNckF2ySlM11J3wSNE31wZi9BkNuwSc/tXt3zB9G2lqs7TtELr9KH
paj84E12y0U76YDySoThVlHjCqCArA2SxefQNRJNdmjof2YKycIbwy1whEJRKWc+
lzZRFTAGxj3sVK7jdnqj6wOthApgRDrNd697wJ4d3cBhmEi6DnLCS+W7qdPsIYxc
rx2mN6UvmopFZPTCCT0hKO3X6FMXyGDBNx2V755RJrSK1tHVKaB71uAQCqT9IL0w
psZ9AOJrmOWq2IN5UQ8Fk0KmTh/Vfoe8IW1rk4i5EmcMHNWw6dTryzm0Ti9cTpbO
LxqF9Z3JmZ3LSE0uP8WkMYej9OBXRBrFoYK0QKCHn0IqnqgjoraBYloQm/qey9eG
xuN/5AfkljLu0T4FlJA1cHzk68W1VbLBIKW6EBoFJD6ZjI4Mq4/fM6ciBU1KRvXl
f4qV4cWyXG/nybDOX2U3y90OEbOtmmZ+oL0bJAc8Rpf10U6/fFiL8V2kR5zCJ8Qf
1u6xe1gglNkxS8cLM0q3pEOldqRlYjwB+s9dIhsf9KL2BFK3Pj78L4KnRGQYuIqt
bzQPZuZ5OKGyxZOBBElc/VsCfW24Ut3ZNx3Q27gI6zeIFZVWboGsWpuaSZpIlFGk
BzLfg5aLwZz/K3b+jCDjOY8eW7XzfmH3HKZeyRZWLGM1aDZ0213PXEi5ZW23u3MR
jN5GRsIttv14IiPqmKnUiD7q9lTSQFMLub0v5Y65KRzXg/1d7ygaKGRCFyPtSwAj
qXGQ/xZ5H/6xOMV8m929RpmX4+czo3zXKe9M5zf8S4hnK2fdZhmE281/BJYpcSGI
noyja7qzzLtgtu8Yy7B7M3wRinxBE3mxnsCgYFa9zuJehDItnI1kzut5Q4vSykF8
Ik5nHovdmOdwd+flDQtXlOBcFEqUr0P6J5Y7DD4a/3QGYjpD54h8GU0cYxrKvPf+
c4a/DO3HGnxG/sQ+4LIZFM1jSePk31cSbG01r3V025kehLOgM/sKa9wy5xwYwYxS
mrS2Zn0s170paq/GW7K8e1l3ByoGv+b21tsq8bVr5+gQfZvOOxkHCOeZGGrqXkBK
UHPMr5os6hmbmIqzH3Er+yz2sk4xsWJNGO74TFYp2+AL6sDLi5LebAOHN68X/xc0
Gkn8h7YeUNy5o0gNpRF8bJffkydaJK/8P8W5lGAa6d0JWlzT9z+DjwId9WU8dwQN
Y++j0Exqy5OsiDQkO25MR9neCUgjV44XsfdpwJ+/6T7wjz91kJwri0g/lKtrB4IX
N5G/F9BGniYx/blp+K7yjvWYr6EmvzKOfeKffhBlgF6u20UE+rA9wBvqjvHxWKSH
vCC/L+ZYqJ+dFaF7PVOIOiQxA+po7b6By29ajmIhAlS7vZi2a8AOyFlLpKGY5tIB
3OZv2ycf1b0MXcJiQBJN6U+028EtEzyML+y6qIbxBA3i6UBXBUEhmx23DVRhGYQd
oQFpoYOnRKm2GTlV8ZZnP2KaaWvArBti8cpIDbhPXWUGDsdrJJi27TZUCM4t/CMh
fF29shGHuwsrRzaTAHKlIfbBdLalJJs9mSXG1bobI4jVMBbeTAgkOb7susvWpJ0p
qUAcz8IZVV6unDDQlTd7V/tPbDYvjyu1Vn7eb7I2pwgWZcA83KH5XVaOHsAVLLHW
e7kNH+NEaMJ9yGIoxEL2EhIYkzADUDYkZ2OkixpP1kRzekBFiJQXbhSoPkLI4FER
iy3tQZPhs9YcIpPsnsThQUJqMrCvKLwXWO+i0AY6lbrd92TG0eSD1jaBBnBPcpOQ
10kOmF6lPjXlszU+BxEWLTDVuvWjZG7m18k4Jh9nJ9+WQ/etzvHpIKzhcEngJXa8
NOHz1CDKjdj5zbYBHlvJTq7QZPMeapRbnLRZOQ6wqqwh/z9yW7cUkiSbadnPJR7H
oVEqWP0R6rbDp9UflVmKrWAcNKvYHp/i7hARVjm8zt6U7ADn+G7kichf1VJSmAM6
pXe+W8MpZzxBegvXCikZfody2axhPFgEqj+M2TF+U2XGd5aKhd7spx92xtWdT3OM
+cEA0iWqK9d8Yop3omWKGUSBeDcOQmbSzA4W/vMu9VI8xoT75SR/tx/UTcsfSWdH
msSFXFZ7nBflmwoty54Wr0sqpldUzT1hAZ5NKcq9b2TqVXUHoxxoY+J9DL3EtZ+9
SCg5v8WqDiUlA+sKh/GP8XPFUB5Jm8EOrLd0j/kJHkKVfTlxZwZeiWMb4DSpvlhH
2TmXaCKeiC0wayGE6uTZIuiNtTxMACfPjBOeZWe9fEZS8zyPJGoWy69Hyz93k23H
/8Wgz2pxm9bCAcD8w1LvyLjkKgCFsU+nNXmubEegjOxTiXXFATQghrxT+89Vorpg
Nsl1VCA1TuXEXDrLOdNWkJXTpwDIFUnMAvdwvhVEmhvXk/O+H4OlboxeP9O/3Dcq
VhD8Pr0sOvi/qZeNp32ZDn7Q7Zz9xdl5qguI2SwqOcdxtNVjH1b0HCODaysJA+qV
4loMNCsyzQEyHPpzWZfkbIdgWROJ/Wry1ic9VV0NmInu9Gc4j2yZh+4O6bYlKZYQ
8/HoTCF1s046z7QuAWS4ROS7MZdorxWkrSI/gyK7CWrIvkMnIN0YPxz4xuIP7hP2
BdFcz3W26fyQqlcgdjS65Emw441Sz2HC1yi+Edp9FtgSADYaTH4KRAyC1XrIMKxy
iV0HGSm7rQxEAx7ar8uSfcVvk1vW1ltN/7VJhIKVilbeE9SEYx+pRk4B9tgqO++P
ZUNTTf9N/++ccnwHcg6GxVVJsNrFLsekHaYELyXnMkmAQgPREeWzhU5hzCXfLAgp
RwP1qvOE0oAwFjXLrlQ+E8C/kKSBGV+mcE6+CNCC4uvBSpMOFm+KJ0zWZ0Mjxn6S
ZCnNTGY+jRrt+a0GaAgLkH6muUknlhjLLeFH/0a5K+O6ReNKEqYp4lxwK2LhLYnv
IDuNwB9iylCE6SpYSBMOwbWFZuaQHYvpZE4vwBsEs7SuZmqha9KoSnhIER8SW6mc
ucZNU1VpJAAbpWDaYgRGDtzZmizRZfDqkKYOk4UMDZS6tO2gw3i6RAJUL9gt3arF
BSTpI1mDPtYQ4M8VcTWL7/s7nAmzfHvtiY6f0JRQ+NxuG7Kyp3jYK8yRgcrhKrkE
rc/prUYYw899xLmk5kSz1tUTA0/wlaCCtxPvpS/iskmOsK7aNpv3VrOg3vqXzmDV
XutkD9Dk6o8a97bqDbrJBFcRth7TNmKpS+ef/O5xPR470Hylkb7PVOGpSCCSkoGt
denj8fiF9oYObSuO149mNpSrMvPFMOPaDWs9lpDs9uW1kQdcYR00MJix4Uvajmgl
bRcQLmIwwYcH6lWracX4UebfNd4uFN+gj5wndszLAUXkRw+74biGq+v1PbOtyYMj
PLQ7zAyHIuT/BSGFS9E9lnY37WowkllP3P/CPJkMdkj0wtvrQr48csdperYoLM1F
AbN46fiNC4jKIft1RwapuPamCmDKKIaym8LlG6gDPIc=
`pragma protect end_protected
