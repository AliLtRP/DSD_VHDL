// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Ys+7CgAgzIQ77hcNJecC10SA1caJiUCW9uFQWiVD2zTBn2KXN2F7QWGgM91gHeLcCNCn3Fx4B5Jp
UnPHO2a+SDzljOjImgrixIk94Is9W+DNpSkklrIBf0EuLjiX56F09sokFcJaHBnzVc3HAqHp0YPb
sZZh0TrKuJt2Pu6i0NFwLyhHo92jH3HDRkv31o6dOZka4EC4PcCPhU5E6tQXQNadUume2hGSEeVp
4E97dUAlY361ZtPrMykYiS6R2np44mBFHqlrX1WVzi9jhIL2PBjT0iUj2Fk0uVvpdgmGynCpGlo0
PRRJ/qo2Fdw5/FnzoHtlMMU26IjdCyoYTrwdQw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
aMYspLgHEDNJe+9+1YAS5XuKZRWYRLexynM7A6JZKAu+7d/LzSvdCiYaMnOEyxy/v7hatJOocefg
/sA9582tu+CDbu3Q43X6QPk474IVNRxEGzkRBkDB4m0OWsx/DVkyogVOV966lBbf+WH5SE7IG7zk
Z3khaBiYjFbMbYwUdXO1Z3XOsyOXjTA4Yp0X5foibc3XMBJ8dXQYyZy67zatlinL58jJLdGpjX8b
9pwhWLVwFvOK/7iE6u4SBaBBlZsg0dJVmQrgg81FUzJ80Qwz0Rzizmp3BOsHLgZfjQozzByEZZQD
bVwoutTLGKETbtccHbz2109vGO5scoF3Vk3cx8hfhZDL2tzq6OGIG9MFvT4iPXco/VKiIE0QkeRD
lh7KTrl5d6dep2+w/wraoHlETCQPulm+V4cf/ubuxzccniloZ1KJsMcbwSmvXNH/Ffv8JmSD8YhM
/9bemc5QfbCnineJLM4wkV0UhDA3ANSRO2WxxNrJux1WiaYzVzZZJ2dR+yDUnICdOOVNCkdgFg9P
RQ7gOxDozMLY9PzaXT5dBmHRwg9IwzIa+WRKJebQybKItpmBQ+dxCdOenT9G5p3JW9tTmeodvAFe
CbGw1dsP1DnrdVen1VffcRTqdkf8sI0tVzb2LVmK/hOtIEP+bv3aXKch/S+s44yLWCzUfSJL1STM
eNFt2fR9Vfn7F0yNWrp8CTpcjuqvDoYvfziQrYD1tAaHVdwq8BgzDh1+B8M14YDlkF8pqvAVMXZC
xZ8k6BeVYq57qksUuTx1s+IwPPj+2NIeJqBuf/3aX0Pi2UkJyWBgc5R6LTYAEYRaboyOUPtnO9ql
x96WocIXRwvfFfuq3Hsm8r6bRe8/zNbXLRmRTvE5aaDanoXSCU5Z28M3y7hH3rLqKW7awfijdZNR
KZh0p9D5jI47gGBMZMHm79OVzyPbFJSfq95LkPDlCjH3S+z7Githrs/JNLMlXwfmmfi27Zs13JKN
IaA95mVilbV7AkBSK3hLv/NMgZCC8JgG2w0pTEo9J7AEw0tvvD81yKulN50Jbiclb7yyxnKNt6Ht
Gv+Ufl1CEhY1k2eyb76Fzi2QZwZNdKGu8l0F/TY4Jrjlr1Wc5Xrrm9UdfTbeWBKN1DiO8WvE4uMn
RonbbOSAY0lo5rV3UDuerVxgZkpvWkp1+bDHep1VnFXRn1YzmlKsUBuLTRfnxeCC4l3TNbP4l/gT
tECT5D/4n8EvTwSssmuK3IWkMl9OB5hdlYEecyHsvGX02zJGGo/5jgbyGHojVmOlcsoB2VhLUwG/
ULhzlu09meXlrk9HLuynIfWeOzlF2ZkUlEDzDF7g57WZMsjNznwE5ZdpPyplpddeEZ/ZyInzhjxV
ShGgPpcf4bVfcgjozR6E0vcVtR1Ko79oX37JCAvBESfg1Aib2szaTmw3zLlckdxjzvdroFj1CuxN
to3J89uBMQ5XFfOR8ulciLD2h/0sSyyyq7anR1sD9XATMJEVEWcsWeUQ+oDjBZ6ntHo2FRZPMedF
5M4oGJ7cHOw8shxjPbhV89wCTaUICu+F4SKoVqjPY+niP+XF0XCFkZyHv2625lBr/4DUY+n0FYbm
ZmYDFY+F261eK/rGR1+WwOqITNI3A68K7cZlQ0mU/US7TjAYbZJCrt7LwjWUY45tNFWgGqI/5fQ9
7y52taHpVkDCxd1nQEILBBMpLQRwSfJ7tT1cSOU1+bvgS3iYgUMZBeKFz0CdsTlkUAg5bgNwIara
9RpqU1cESZjilSHSyu8YLZLysbPPHyTvrmcaFACz8VakZCp0O8ACm3x8lonZGZd3RR79irg2i3OI
Za6qYtzFUkcb++ukzAEQyaYocLTroWn3W4PqEGxwjX8KYQIrNwHZHC1NFKXJBdsf1/lfm1/oTZ0/
yGj6s+YABUia/cDfrsZWnBTaMtP6vWtMm1Z+EUWV5N1d/lm5NRzrnSrLSNgqr70e6ltEFBxDS1Cy
ADe2cKFcyT6+7ruCR6lVIst63U7/Qsi/p60fDTlwoqqmIBNljeXsxOWtglMdqTHKrPGvt7+ZT477
EDU6+JyRFuyPgpHKaacGqhWfEJlCmHOOthcjOu2jmJ2pP4HsQRPEY7z+O10TjLywqMOQc64/M7rP
TUpihCc9Z7VCtGz0/F9GFFNhdTadpYvMdqq3a+rGu26NNEGx1euN1whtCPxHvm0zpQppoAhqbelk
DHGsrygckvSWUUz3V7LOAvFlKESxyE8Ww6XscUD5Z6etVXRKi4dsga8NlorrJ4KpawO946EpelZB
YYLBP23HfYiNWLDg4FZgPIVm/8O4U5pXfa2MpML7/0Y70/gcQ4U2gaTuyTZZScKBWgfR/NznWbKb
Js9u+0hjPTlwE23bDFzdSdJDHjTChBwgonLGDqAzyGfQC4cUp3e434Xm3f/yy9KUIJ/2HVD+Agyj
Bwo1IqeUe5ixzXl6Xp/PxGbAFDePZS0ajwXNeJ/n8cHvklU4T8+qfcbhZQ+tYA8YkBe4dTiLNkEb
5UHdfSpBelzx8r4QpcBC+Ljjcu6Z0HMwHlxcR3ajI0SP25bSKd3IdnEyML1i+TxSr1EZJGQ2yYm2
U4cCSS2PN0x40YkKHG1qhnLYQsymUSqe9XaE23PekqcN/fV5XRfp0Xfi+himHdQdud0cyt6Nylgu
baqM4Yd95V0YWtBI9n/zr47NvL0YFy3hmLpjI0sQ1HkvAPgSoFHXlDcy4YhCrgd9+a8SLtyl3+Lm
zZLn8DEHbW5vdc+KcR52UvJd0aC4RKGEl1wz4+Jvnw9i23pAjY58hUU6clg/6TSXkGu4u2MZ2laS
KQjBSF13FaPx9JJItQP+4jqznCrLIMtvPwK2TWhOh2hisroshhYdsavd0yHdLdTyPhIgsGdXRyXO
5gIVcBTIRtjQ+DeYQgxgRcwnGVNmukGzeOIYB7nnyDPg2wibEFHpWodn0Ft6+Idbr8FkUtXfgK+U
wh/Lt4zGqa6hbiWIACIfHNAO+XaS6inKs4zsMZLl7IPuRTauRUAbK5yvoLjDsGy0yMn17BdgGbHg
EKM4iptLLYrBSYZu1wa7/9btVgku/PZVbehURNJkLqJ5UFafG3yFgiij+VOGxKs7R4YoRiqK00T/
KCUiT/NRnpqj3TJ0+IY+hgpCxEf2/y18YywRSeY11cwsvp55I4Yv2oqaR+UU7Nt0KGYIsnDhebsZ
yQo4E/IkKR/zjgpS3lK+2k7BRbVPTTHRHcY+U2ZONFRDYunSQktBWTq5pgF6BUSLcC307ib/NeQa
N0DV71u45gNCu4p8uv+rcZrfxdgh1N/MuRm+lEqzVoA5RGkJdGt7iXHgxJPCuvBKJyjjRKn02PZF
EZGIvWEelUjRfXeAuQ5YVah38gHkWfXLnFmaiZmlvroZtMGUDmPMWuytI1hFG3rfOvttKrYGF8RA
0B6M2CEbhIz9smq3Z2Hnk5+LcHQtxMqNO/9RZy/lkuYhXYB3fbfer2HsaHGKimBiFHWF/hvSexQB
h7zv9PUFKHKEtF+BIu5ljbLCn/MXx1SKeiiNb6Oc4XTo2WinLQY1Z3bXRAV0H/ZC6HBRCv37Lvkm
XwQ/aKLbZVMe4Nd7c2Y0/HPxuPJ1ysI/Rz5NSxWfg/coBrXHWpxgFO+5m/OpLFx67UGW6eTezYyo
dGYb6miUjPXK0UivrhsczpIf5sWjmiZwOmpaGvOwq0lJrkvxglnhghryFUds8ztMg2bJQuBKrZKh
x4zKvDmNv8V5TdD6XQOZcW+z1Ax2bgfH89zkGaVM52uWPEF8zwf88tER8c6NgoT4ra4wsLy7/1hp
VBE/egc6JLpRrF0Q6mNpYBDS6AV1GU8VGpeV60aC6dFDxC6VuoHu58QwdgjEmoSslN1AJLpbDuzo
32WSmB8SnvqGJ/89CijEktgK4m79F93HCf0orAP7jBF7HPCykJbRl+qvsm2MCsPAGolkbtRUTUUw
OBa8kbx2SZF26emOA0CaUvlN2lhAJkmmAKWKxKKZLpQRtgWN3lHz1cmBeGOvJ+fNgzeQfF2RZd4r
ls88BwuSUY995HJqsz31J0jKKxHL+Pjk/OasiGMBCj+SKNkRNw3E3RQuT50FIMsNW6JnF1O4SGbi
kTQ5C6evVIgSvv6lyQvsEsE41yl3ZS0hszlGqhkz4ez1OMJXmgyHjunIzLeuC4GlKyufnRrQDDRQ
ymE9quDV6S++oWMZmHRzqKKlcRHHYmOTIP4luz/cygMUMG0/qbRy+0/KAfxZnKa2uyhQYbn0CC1b
OtXDa8b/2Cu0gX6RVb4MZYKBuZJPiDESSIzTQtI/IpUGdKGM/AKkdlB8or7AY9P1mmJGLp+4QtY4
FAZNXEtBpHWzAYvHG8gscQ7WVOhRCwIHKI6XK+ZaXiM6VPNvFTxiqv64V6ICEoA9Sc1wJQ7Ue+Lm
edf0GgbMSXDRR/VjNLOC0rxEEeMX1Nfi0xMOHTaHUPsAhlPazq19IU9275fJMpeQSKOLWPtPb04G
G1+8v2HtmLoExzPilsbg8DaNWfN2zO/vcW5JHcl1TcBNOWo+aUr199Hy18Tf3bCtreAlpJ3WG5sn
hWl0BSAufX2IBvaRV2Gn3rVQtp3O885YK/vqfEQoI1QUft2rCXOQ7Qvc5mK/wouGcYzVSALdJ4Sd
NfZoS4S9H0GVIe4GXDPoe/7QsI9NHHKHfbgMtt0rMsj7ObJre8KyW//tEw1VYg+BbST6umASRrFW
dhf26H6EQE9Ltw8yVZ//iRGh2oMRn/AJeyRsaKvvcIXgYGe+VtauOn5SQBG0fjfsOqTvalFLrV0C
CjV/MeWSQsMSl21LoN/qDvMBKm7ZV6VgLt1WQDuJDTKnbrGPyT6ZF7cT7ru4iHAWCKE7Jl6yoVKc
lLP2kfJDdD5ulWMZCR228Tu2G0L0oFCR8aOEj34OJaNHlj/G5eQcxBAip0rLKDYIW2IeVBGY4tXc
6ZsfLkRWHRJMgaRuSRcbhUgabHd19ZxfhzPHnqpCdY1wFtAN89cwknKVlgJHbGK8CvaHQtbHWrq+
Ptt5IIHeRHfy1YSU5JcHKmsb7yStWFDaZFkPWOfHuOrbBVwMwflCtEYc1xKRvi4xHjGcBBuRlLJx
FCPYN7GheKfqhIkUc7qXEcVfLvaEw6CUZ2Rzk8eVm97H88C6+Swzid+Exd1YR0AQKnLd16WC0Xik
bLpae7EtDfRGoiTW+yOPJKftf/MS7Xqbb4bLNg5aJbzcz/QR5rEVsH4L+kecGLMy0nZ8IJ1LTdkF
E2ClpYguNYVKXiWkNrzjB1W41tpz18G41ADAiwezme77AeuiPQ2P9QM3NSPqZSSJwdytk/cDqCEK
w5JIbQrWVn9+9fNSjgvyPv+rCMV7kX8xrRv/uuAj9aMueWY+gDm7exC+E8HCDJJz2+CGXz1wxXKk
K8bI5KkrWCdw70jPoEq9/WM2GY4YY5cllISGRMz+9vlEVH0h+1tPsXUSexoHa57r4V5B13Qpfq7C
52EqZcI6J+d7L+M2OIr8F5HndTiNude7w6VsaaxKe4D5BuvXdGoErJIa3WHM5qfKZ/o8eXB5gSSD
HuAkL7x8XuVYgBCasIAetgQKGRKpZLVZSuseGMWzPozWi2tk1I7nDJ+gtskPX/BnbgAaVqakIxPU
bqxekkrrKvKc4LpcJXmqmL3ryuM8oDzH6gSoROY59/KX6KsWAf8PbEoXN6+f2qEg74d5+5dUTwyG
OALgvWnwrUz3PFJL4MkHuQXXP5OoX674FKvz11aQlsOVujAuDHYr/EWRpJosebMMmMvRTq41tbmV
H43MyIpeKwIPzgHg+AOrZPiJ+u1w/MXkPQC1lAr5N2eyCsqg6w3pCp3O2v52ZLgpGkwYXRKaCoRq
RJDvMkJh+ujGPT/KlLo+rOzDr7QSbC1o+Pvbo25C4yI4Z/RRAJIQRiIUf1wP79ZdpQm1+RJXCsQw
iwUc7fS+wR2DwRuYbf72ooniXvV1gnbahPb6q5+OPBamJWKTlpsWC4XMW8qdVG6xj5EHgVrgv63Y
+Pf8T9ukhfrkyTBTprnbd8Rh76d9bMy+9bgWEhKBWwouHjLs7Oh7Yt9v0coffJWJf/hGjq47KGs5
b5BB19Mz/ZIhU2QdpsQopyNcjA6s3FeBeLtI8m3n/DIfxzKoGVrjVhODB4n+R2rPU0DpV5RO4Fjk
RYbjct7H0p1tALDzvOMgN4qf5sfrWQCIrkpED1BKpetFToR++seV11AL33EbJzfkOquHiux5Ndtg
zqFv7qq+onCzbGWQEyz7Ij0WOqJ0MZAnev+tmLzo41tJwG6ox/PkcvEd3h5SdqTazgRsifRZxD8h
6/LBMHvlaZfXx5wTHylF6vqpeOKuFDncvhCQaIOIw2oRbZ8RGHkxW9kSqHu5Rxyf1DYckjVZDX3m
+y2FbKX/Yrr3RGyhJYBDvT5ZuLlUDr4UJcBY27ce4dMwfLJc+U7c2hVy79y1NL6KV60V6gJvzH11
HD0Vf0HRuTtKrpcYl/DIFxCDzJVM7t3tw95tzt4GYWZ7+nxNDWqPDYAPxv+K5UXeCOoDO7yGtfz0
flrN0E994fNlhcy6d1XxWadesSoTgDqGBdV8v/xITPjC4G+jSkXLAXPsj9aBgi6wd4yJw0qoR5r6
MwNE0wP6JTU6l6orsjUXRL6Bf/OXqglVvMrnMIy9IR/8B7+gmi+SSEM1oK+bhAu13WGFZ6Cz0FOV
7J2u8bKMlZLB5Z3vR24g2fP8UFrtAkE47EWREx6vLUTlsSg0FQhgBCfP31KnIokswBTyyv/CMXO0
xz8P4suzk1ldn1VxgCQpNgrR+zrqCC0q2ojP8o9bHnCCi0tgznEW6gQ/FrZTEF8Lu+MM+pY/fr/s
4Ix1o1TqarRuHW/8r6yxXCVfdG8/S5yXxn89C6GhbrCFdCV+hbBsujRHy3WfPz6xjvQus5clq9uC
zHYJSyVRNRJR+y2xSf90AOjdEnMEfEfO32A7ZvACA/+DQkhM+j3YBJcfRVu1/pBaNRcmLeepymPi
pKcv84JYLcRMn2/prcUCnsmLDYyyhyzFiMmDnF9vjPVhzxOZMBddZRsEGLBClkI5OSPV0Zawvt1H
EA+hvCHy7hXov+SPt6KqpNRhBOvyJbc2zu1hQ6dbr7wcUSlGE5MWF/lpL8FxpFDNm6HM74Otfagy
kaUanPRoeyRnmSTOE47LswJykPTD6liUdRWFIZfN9gkBAs7hlVgdXZ+5OTCO5GisKukK3mrcckDb
uGMepETuXqFDRzLSVa2WON0tg64zDXYfqk+wVuqOph4vdnIZ6VbOVBnVftogf76j6aG5a5hzbEn5
NiphcohwznhoVclL1yduHP1b9aBe8ALbJAqfeD6SUCtjDEfcaKucqRjkZUZlLN2JAkttDP+HVAPK
LICAPXNuuJcI5tcOYkJJK52CagnEmjjcF7Pv1/ZVnOowIwPlE7jygWN2a8iqiB6fjrhjI7SJRHeM
cv94AN0pwXwVp3xWx5+BWvQEgp6P3EhOrjPYKG6QPrpGRFJWOadyqs8wD+0iGpYGqxz/zECoYsF5
7eN5ojwoNrhQpRC5oSORQb8uVjc9woIKn9v7gHyOly01ZfaVVBwxsrMsxmBQyIm2FexF9PWkI8Mg
B8weAh4qcdG5wFfA/qllCnKeiCySE88dz8vJJaOsKrz26fofz6IoZZ6V1AozRFFJwYf7pkXA7l6z
8G59CrS1E79/jDJH7HbzoDpYRX4FRHF4y9cX6pnb/+u9ho4wKI8DFkGGU+DiW/uddcVgUQ/0z2sM
5uIWm4eoLpW0yMWmb0YG2ChZ5Kmxyf0XoNHBTEJCzCkYYIaEnOLywz3VvsyskjWRlhcwv0HZDz/7
ccVm0d2vqYkjPTxNwI4dzTbZ68pUY3sT8KcNJBF90irEN+NB6N5E+s7PJ5WWpWBhLvUi9S7/OdgJ
HrE23QJnhsiZ1e6DxB/0zcRU7Jz/9MCf6M44hT53ku1h2Gi/iyKM+KgNATc52qCb+D63lPxqvC+f
gKNUiOZ1ax+PNf8g9lSkUGKP8QnTfFpTgQvTIgq+YTFFhcaoSSGrgO5lNTRj4ey8mfgEC3h7nWeF
FTuBmdJwNsdztz+lVedT4OOHxNS5P0B9xKdNjrpxdZzgp6x/bdoc4EkHBRk960XHLQxuJ1i3Lz4J
1e6Vg8DTbwibshC9vs3yftOSLHsG2gthxiIzfIA49FnifhMQKsr8d9mzEtco/Ay9GFKOQzxLZRJq
VopXvlzTrUi8/ZganTUa75URH4CgUdwMn9UEiCmWfxkEX+m3xKZgSDSNFKTLDmd+RXoc+kOVFk60
DNal/GJVttMuMx6Qo9sn3wBPR54eM/G5+9bnF9GtVlwn6aLRk4Xfb17TKjFYoKO8MGF+AWmu7EA7
HrOddbOMvD2lA8Gzr2Dp73DTeuI8Q5+3tAVxVJI9IYMwIjIIfupIB+/5dT5QdcZcMkMyLwiKyIiN
A4WUXQfFbeATuFDg8UVS2fj5OE2zZnOG48OoNWhE2fPohA4ZkDRdMq+aWWyztXe3S7bSM0TmJCxH
hdFKVTELvTyYkPfpF2xobeibS+2K9shWmoNUov4ZC1VFKAN6ZoryzQMniRwnsU5pNRDS8MNl9ck4
+IIdl3eoXbSwIsWGcH6BMluzcccLswswhrwfzIOz/rft+RcoVyopwQ9MVpx+Gxv7qMBUNcDItq7l
RPjFoTFd3hvzZXHasCG20ozNVsfQ5ixwFrjHbkBzBcrdUcQGrTBLgiKM3ABbKzWcfw2AO5OryGHF
2BYPsbcirRwqgAPurc8A79IIYL5eTaoUCRTSc+jUqqwY/0DpGGZG5rjil/9lTRLrT1jKgRv2shs5
LZpx3NDvfd6R0tyhlDVQsSf6HMCBLm0xtJnyJ78TmFgbFMJUccFNyCXrF4Ut21Qd8D9bkiQNpIZ9
ZLDEpNgpDFBBK+Y11jOYKo2VzjzGlGtkKNr2CkMPHDk5aFRS8EtIfrRBpTYNLkGzqNLVBPrq9KXI
0zEYAHkjjiI5vuWPjkZHiGfNZObJA/X2Dg8n/52cq2ggfZBygfCjp1nDhwMriVXKQaokYoRyckAD
EdfXj9kGdIPiK/jdunL3u1zm45F38KmDHYsitjuLXj0TIuTZqbdgPP0AK66bYlSaN5SYfAlyM2x5
qiQHS49VKsVCDH40wmpG7cJTU1bwDo2AmeaEoPsXjHqZQiBbpO/6deMZD95PS8NiebcOznu8zqGV
s9ZDrqntNh4vpqm84koVtVIjO5LBCX1AVw2aAaW788oIVGuLnIZ1Y6FmoQPxyhigOPN8FhgcRlYe
rTxJzCSi+mCiOfZi+K3e3W8/sKo9tx8gOO1xkO51b+ow2L6PCpcOR0bH5nWNWZ9aNhGJhsFe64xp
JZZJvtl+f64dNI/22s7nVKIwYjGb4GtqO+VaocLAohcswx4quxgYfZwqd9YGrh1qEpNq9lQeYPYJ
RwlDnHupix6C+l+CCkS/RjRqNQo+7gos23HhT1+WPPCdLuG5rm9YiiZdMULnDfTZtKMb9QJO9eKD
yY7PGnSgshJcnJAxauuyeb9vdtDXSkgzWkpOcHIskE1R1WecD0RvMHm2CMjRKTEbLg7wRCZkp7v5
J7BunHnwPJBL+hePWvRsv9waRTnnpp5vo5sjGVgQqsiN+p3zBGV+jz0UoY9fZLjvrt9VrpDyVglm
j+DyHGff4LU96SVCxyhNYaUjZpMNIssMf07zBGfaK6AaXDbHzIrGgjOQt0u47kwNS+MXO81996Lb
petZj74C7DyU6iJ/kPwc00BcE1dodHjyRJaf9yZdfv/MBQOIzM0Qspj1qgvEysA4bZ+LzyqkRVKS
klhBmipS+LhdN3cut/kBA1ysNZ37OeYyQmjfLMnxgJfio4O1TUV3AorVVTdJD4+IV0zixK1e/6Sl
HgXXR5O9oW+GSTiJnCmjiAcWgZcOSPZ5aMLRvUwz1815uxczzfP6gyTfQj21qEfNeCxX+swYaWx+
5oya82h9LcQ9XW1ANGwdinMhYil8DmmUObaJpWY3Kcq9rNCHbg==
`pragma protect end_protected
