// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:18 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oXxHKvHxxb6EotMEORKx1WSp/QBfjHusDR64g13vnEHo6GhvNfkBC9ntFFaR/S6h
qLLGEDNuwFVOP+KKo3bpyTYBxtZHDEpPEns0gG1RHyysh8YPHDF5Op9gHRRoT0QM
moP+IQ50VvfKEnEKBGi9QFeKt/PPSCbLOkv61C1fve8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20768)
Km+lOoniwE+r9ZcmT1IIMWcyLT3jYDrNALjiZLLNz8NPIVGQ+zSSBxiugwoSBaLZ
aapv4Eij7uweTs7pZHmAz+WmoAC1J2F/MgMxiDXoya8KH2tq0+6AWmzbbSGov98c
cfSlLNxMot6+OlXR+aG1SXks1/hlJhxsZJTYo0wN/nLTC08lCO0plS/71n2PtzxF
fro6cLU7E1juJ1QbkrgyUHs8uHAfXOBze+MZS7QYoPWrytlp5aNyAXx6Bi5xbIWx
QB7QsHinn1hUKmpbL00du0/tMXTIuBPWyK/fHzUGWPfxyBHfYCGsk9RCL4PtOMrL
jvmLryZsDTjdE+deZk/L3vwoFEh0GOlcPpNuuIR2JjaIYm8ZWyR0HgsFBAGFOrMW
dhqE7euozrIfSuT8IzUyCji0tDqyamRWztCwV/GZescz0hqnYZ+hx4kh7fa7OgEd
K1sQ5zUyJyeoojdCOubS45hs0KvReoPm/8yIGaFv2L1NApG3op62PuuDN4L+l5VR
VCiwpfnRUSLi5RcblrqTHmcojPIiZuXgA8LFNaF0xlcFZJVbHOkp5UCy98UUxhKA
5ts97/plAieQqDO9pfDbpVNbjIkWI5A16clyihYsJyyMf9gEpBx0j1znOVf6qMbP
bb/VcAJarcCiFsF7R++VWjS4caHELIuXoq9UtfOJ/eX9lNSw5lTAFNNOdnbxuIm2
SGUnYckOkIlL34KxbxKCCCH9BJPMB8F82EC/XagrRyNLjfh9WNyw3y/FVRKg1HB/
bCr6GLBxSv5InpmEaHxo0UvE7vwUoKK/6NJy5w9eZ+/ozVsvhNJduOlI06BpJIro
W01VliKctLyNT84xo8fxbltc3UmxqlZuYQ8FJW29L9h5t4820QmjSIoFUF6cB+7s
iinzgSaOn2Ue671Pn+t2jfg08gXy2fuwzD7r23oacEbZeoRaJz6hLMxJLnH5suf1
fXExzGfE+3QrQPfXTljXRLHc6wIykeCPGnmRtal/ozTRLgNwT01ulLC30IZSBbDg
8dyUAFu3DSVQ+pmervJA8aAD4w8L5n3UFafTCdCvzHkmZfGqbo/bAqaDeV+bzaNY
2wkJto8HqMxS6+YHgPZWe5cAIFMxwrRGuuB/kMd6a5UHszq4R6cREE5w6aZCwFNw
rlivXsB6KJCEJdUIHuj4SyclfDSAgycaF43zwDIMZoyT1YradtV8GZSsGxnSY+c2
Vovg5MJU4BecPIuX6rBILK3zznIm1TQD/vhI3BrbaTVieIkEXDS/7zRtjIRMADl7
7ca0k9Uknnv0uOmDLy1oMYL2Cu7SyhfSFHtJcj57RxRzbo4apBN5aLYxNtGXP4Ki
9db0VJ4hxZyhi072ddEHsMRXOsUol/f9ySce9xe8XSuprBkWc7UzBuGWjbwr696F
WvJIe+UIDJYaPbopKoV0qWkIkgx9pCDh0cCX/eCGbwGK/QP/gnIhreJsWXV0gIct
sNT9QjpY6zIZUspvgDGjtz/C2k38XlQjs64Sx9VvSIpV+GcPbzp+HU7IRg/+9OzZ
jb+itZ0bdp1RvQsesv5RGcrT9SmwN8tULpdD7U5ep/Rr0bNOPw/MwWLJN+2YMZQx
AAs+WgJusSkY6cTOd9Yw5FhtR8rVfgIyIKqN77gAJkCnsV/Ws0gOr+psX3/3cH9Z
6TKNfOkhg7R3e4b3oV//cNRnUet8eWADVmCsue+gXDcuoRehHxGvXflLrbl9uUko
gRyDR/v1ZJCgdxBZD65n3cM8/0FEqz9OlLJOMot2dsndrq4aYp+YBmMc2AF9eGQ6
OHxoDdyn+v0sHhDyMmL2vw/rMtRcSabO+4kxg3h7SdDvi5PUNJRng/KnMBqdNXuH
9c3xrqVGmpGAkD8O8j8btPZyHzp/ja+sH+I41IR+WTlLeWBLKum5soGGQFVmXRPo
7HEfs8pGiaSVEdnqFzAJZSBGPMxqjR9b2DxCSYYAj+wBs5dnzccoBkQP1TWYHA/w
B+fQ/HbbKXdiPVHN9l3HI++X8vUAMTNOfta+EvfGWAz24yd0e0NtuwFTd5V1n83A
8LAAa+tOWnFDBc5CYPTzQwkFDopGYcubAjJn637ZVe68ympPrbKd/S3SuhFUWqKy
P4ej6RQz5B+izX3QrLIzBJssXCnLpzojBpIW9+BgXTUR6hPHv1BF+4jEv0L7iZKz
zzdTHIbcfFcRUhCrP8PMsnfxIkOcrs+1N2uxGIU5JOlU5P38Ss4TIgII5vcFDAJ5
EgIs32GaY9Ji6dI/h5Ftlc3ppk0vljxHlG7VlTgUGyj+efvcIx9CfBJp83+1OZYe
39qLjlI9YZpkqBXrzBVc2Z0gjEXdC3TGUkoDlnDLRD2XuUsCNepuYtCpEpa0+lyV
0arErRZzH2nt4wEtRrJdrlVqcx/ImChPWKGVMK4UTlfI/PfitlFNYh0UpwahL+lm
V0UZPv0rSpDpSQKx30Y1UHINYnlQEpehTrDuhEY69dofsiIldwZ6qhwHnVD79s19
Saoj71fRNQyYjx+Dram9Tb/iqkFt6POt0SFLwjChJOa3gLwcw7ev2Ed+psJ8StaA
18uVqH0jQNOBaCtC6fepReqCZ9yB7qLtwYHtCkXNrSfztsIA6rDxMxASDhq0Sqf+
jLZShbnCwEN5nOvSVY6a+JRNmsjvs9gccdCAwdg94jYqJAyWxLz2p/lZn3YqDaVC
304qRXCPB5hwgC+16NFRDRJVPL+rUtlBuxyZXOwwh9DftfXnS3dgVJgweRSSl14s
UJ5MwfWU2OxQ+aMelgLp37Uf8XkABQpwyvHPPaDmlmKEtxpz83Ooy9H/jNr51teC
XMAyTH32CzkP7KFyrUBvg/vrWPfD82Fo8fvD8ZYcJI/Kb6kH3LW4wjZEfsD6tP3a
HsibuRDQXPvLF9mDpCo22Cl9FI9+jsxyIUeRNGaiTzmfYL0k2CqYzjgX1OsMcOAg
4wI8sVzWC3TqpkyLjHVc/ZyHUe0sIOT70qg9pKFw5RvWoHOaTIdbSi7WBNIqiRGR
GLbfICgZGHj0VM3var1s/NtYkTEUO1OBAOgeSlH6AGscRKF48d+r9H0Iy0pz70RX
28IfaCUlLrK+Oo7Yis3s/6eHWfzPqwximDQxMQVRrliP4DM+yE93C2IIkZ3iWefW
LYpHk3yCyuYmwqKQP3BGGxprjbFTq/pfUJcnGB6VYYZTPUFSypjt1hm7iL95M+kp
A0p8SRZpLLV25CCjsghZ2IZVfhIXo+iLFl81GPoWv9BUMDB1+KUcowP4ooqemXkq
rHeqswZMN6pg7152Ou4Dcg0fHgDxgTsDNC6QCaSIhBKZnsp2OiyUQCwyr5MlfoNk
cUmoC8Ki4OgBK23JXGluGB8lRd+yaXGl/y9ezb4lA7ClO69qT67neiv/yHvR3Yo4
CRv38Uc9m7coohFNDUy0520UXCgfA18j4nQmWKkJaLB4eaGbeq5g9M09F4eD9qhY
NT6xG6sWXkYShQSycK9iRixym6OkpNlwSTnMVpzm/VHKsIYuyafMkv9aUXD2h8pH
Gzlk9lVtZkIBo/guUsca8idfWvVyA3Hlh7SapyurJfPW4jybUr1hNYHIj8DIxsiU
EMVjPECm+zxELJJmRbYAOsFP0PNHuUW6LOMVV/QMBfia3HfA1/aEd9hfjE3F61Lw
1LDqe8IFtid6OfaKeeDj7leGYXOfwuOscNFWlDvm5Bz0EmGbPgM9CHU1wxE9/myD
wqaVSsNqeYG0XzgeTjfPJbc+fdxTpd4SuW4eeTSleNSRknHM7pIix3UmtTnI+A4O
wa4hbfCRk+b/VlYITHmprXdzUMYb8tePLE35+KLoNJ+eFJi/CfJMOboWzFYVbWEK
bKXNeI6GXCCn8CjxDtRLr55bhN4lzhQ7tVzHNS+BuvsIOYvZUQnmvxhZ6Gunl9lJ
iV9kp0tju6J9U6PVyRbTGqk0+i4RepuE+FCwNUABFqR2lw3Lx8M7aCMpxVtkeqZ9
Xlsc++uoXfAhOwpqoA2CRDXRFDbxTMM8rs546Lgq3E1WpQks1lKRmiNpOfwWnmIC
4yB5DMNM0okgNU5n5mpVGkWpDXKCdFfveMQjylgSA9WTF4QE1EYpH8e0ctfCHzIS
5qkUmaZ9fZP2zGbjMq59QoGT7DQ6LQO2l13xpnWyMq1n1ySfrAUe0Z7cMDd7hvCh
SO52DcbuSe5T30QZShPGc2RbvFSgof7d2xQzkcyMpAgqlL3I9tDRIhSW0P9Ttm0P
Khz1Zy0OXOm/hlFP1Y1OCH4JFign+ZIxhlDhlc00W9JPH2yFchGUZzLJDN1ZITZU
mZV6PK8CSdOy448QzV77/ATpyI/kbD2L730T9o4ZEEo5b121Gi0TdsoORgWquMMm
uqOC35wbFKWd09iPuGh6Xe0kQM+WzNkUcItsrigFsMJNQkvv6LWmQoRGSEe0fQkt
LpXx0ln4DC5Uw8stipQXd0rJfL/xDzznkjaM+s2rFUn0ENSulUCAduB579OFJIT7
+qqohAf3oCtkdBEifctwIJ73FkYvwz0YtzPOE3p2AUMAuaZh7xIoPsdkOWZPsfit
PHLH3Ax524/HzegD15DmWWkCC3dSQJwuLpn+KU617w4EdQpnSiMJakpH5Mn61cjy
aakx3VMkUrqvgL2px0Rn+Z9fzXVMQ+ZJhpBzF3N//FTklwLvPDa4E74QbQjcOVpm
kEnaVoIKDWnGINr/U7zZKHSnkET36oUR9Bc4x9X6n7xLP2cpzwks9a2wMqX+CJ0L
5/63iaGR5Vx7NF4Pol5xUbBqvkwA/9LL8/1+sHB/MkZThrl8CtXUQDFMrB4ISVvi
/w3JrQRRDUMeMRZmlO9TUDVdmkAY+wfwtnuDrQ4RYamDQ2XdHj+CILOnpISWvSg8
R4WliTc7SXDYXIN1Xh3Gm6TSFxN3vLbt1tXTJJ9q5HRqXfOEfq7zxYajjjYA0Tkc
qiPFWArG9egqCr9/0O8yq+aWX1SsmdqwzUdwHWmJjXYSiUU1Vj08RimTujZJgX/7
Hen+wYjf+ao4v/6ShXpGp27hcyPVXk7byz8E3jzIhaxk+BQ3Y9A2vbmHdhga8Xuc
qLdsB9ym7OrY/hzOlDzZHQtE/oRUQ1WPAu+7+gcDGNyKAigak93ASBWht7mE7R8V
V13pYRdlelIkwf0WXyWvqThMaZi28zX1qljxbr1BxFo3oY3Y3J6fA7Uu26tZnsBg
ey9nMffuAFSE4aXxJdTUCbM9P+9IqMUtpaMlURgIMgoq94DXd+/GYKmEl9FXh0Rp
7BNl0xx3D5hh9a9n2p4otiqn47E6oHMYpJWe4IbdqhGBXwGpoliqQO/jssKTAHVA
sb6HuaEH1TMzFPpoPaQCzI3n0j/TNZLFZ7tY/qVoWXoX29OurkPBNnLXTjiCDUO4
ro5xF0LQvxXUEwKGcKtaU4ska1DnQN1Sh78t7idcp0Btd9eOiIN+G88ph/YwA18R
nlEGfnkeEgbnKhXwmOktBqwdGSs+wy5ke4Vd9Y7G0UCaDU55MzyIXaRm0z1TKMWt
yYXC0+JzxoIX3mbpLT7N2YbWxn939ta6Q87qCvYew4GhQ9d+Oc6nOfq7BSiiIMdw
QEoTmr3/JmHoc/kRnZ5P+CNd1h/dpBj8Lc8LuoT0/XZNIzlMm7UflEMqDzznA1D9
MYjK7fHMOyVGjSTrNhpvvex8Ndscw4paAFYmnLPHTNv9pKo+80r/9tunSIXplFq+
O+X5+c8CqIffdGfVE3EB5XfiEZCxA83m3yHqigFEAV0CjpMeuME+hdL2DPxbeX0m
GziX/38XR4jcDNqSfODUsq18yM+f4z6336YsYl4g0Kd94G0PzmyqEgJs5klX6UKI
XbEPoQ/XQJTabKtpY0CgkTEbeNNS+6NnjP4yiaU6Q1YehSqM3v1vXDg36pyEqO8U
BglHyJgyqhHgBetDeMsP1wELC848Jml9vf52MWzAP0CHiTT4qmy4L593N0vMgdYV
owbc2rUnPfkKjOcdMCg/83XgNxBHvN0kWVLurFC5ccbh5rVSAzuPBQ0ZujoGk1/e
qS/nfQkGHWRkniczOpvAcuQWIA9gLGFAGkIAYVyfGpPwCvBEDmQj2dSgRPy2wSrg
75j+NVDbTHlYJjCqSvcyYOI/O9M6KZvhtMNNutQZDz/xY49FTaIqUbR1F3s8mTXh
1LQvcN2a1l7zKI/3BGIi/mW74WKgpt1xsWv6u5ywAmlU7HAnlu7g0Y9FCLesSovx
aRv3iEGx+Wx9AeL9loVQvhvUUWAbhpXxOfvyc+BLi5gH4aISUe/cCL4gqlLkJPyv
75Vd3SAyCDsbUF5UF0Wun0aOgrt4TPoPtvN5RGqQgMY52I+MCgoXmQKJ7WsE2l/f
pWlBROe084Uj23dcrpgl8MTMp34ltPGXM16NLelJHg0B8CC2/CKiPuSbCPlqAP9t
x+6YuNDYmACwrAHGCu5nkg7Ortep0KelwTisd86gzqvYtJr72Ty3BKPBYTVB0acN
HEEW/ftPqMqSuByzmbfDorokj6kyg2JZW0xX+wc+9M1BZop7Ir8Oo4E+nAxhdFUq
Qw8RTaa6CQi/vX209OLalkmsCYXwsPuMO16QfLAf7JvDvZyIvEODOSeNcqoD4Phj
OKSXlwA1uHCdPw4cpIK98VQWfkjPrXTE5nsh63V0w2NLfKW+lpAwdIF3DZuomXl3
6wG8KE+6dC93gA5NnbSK0rzBxdy4X8Hevn/pYscNluN3Jn46i7oAEV4tNejhkzkC
lmydEo1mXj4ZjzovvjLvHb7gb2nzU+eKqWfSa37983B7RWL/aHeBxE/lapQ1fTOP
J29ve7MZJFOaw+EVLcPE7K5hsdVHO7Z4ICnEj2KFVKFV6y+0fRq2oz7MZKmhCr1n
WWhwS4zU+k96ZRvp20U6og9QA3NOQSK67qapj/4OToxLTuK4eSV0gX3Zv5iCm8Ye
zVQcj14WcD5IVWSpu4+gXYcurpke9LoMgl0ZECvkmS/VxSzdlQWX+R5M5dGY9W0b
fZPt9OLCjZiSJ0uxPBwIBfc9xd63UaQaA74DyWv4S1M/F1xvoc98op4YoMEaaeE4
Mq+WShF6iRz8sYXqzxudQjWRiO7lyhOZZp32J4k6wiRZcA0sv83ZwQsJfNnQWtwK
kR/drbAFH08fFv8T3pYKXTNz98WF8xs8k2Ah9Bhx6UXSVZVH4Z+rukAzNOTV1+08
SteDnixUXQ0pM/Og0p0BEl5mrTB2IX9Th5xrJ5WBYU/s1wSjxr5p7rt+fs6Th0Au
BghwjQ9fafOh8CQ4id7PJbO0VIugYSNhrG0t4Ay007nY2WY4ReFPM5eD9N7qsPDn
Z6CDo9wahQk8TOIXk1oupyzs5NnFatR0oIzDZEGfk4qqX9mjPsWV/iPa/ABLDazV
jhyOi4ORhyy48dnT4yHzYsEMooSdXKMkmjfitQjsWGK3IYF4KTHBtNhYRdGHehD2
yT+cNZ0SCVEUROuk1kYO8CYQHqXiR0F7JigmHR0DqwkLM/ggUEAnkFoOkM4aVOj7
BboKBvsPVTu1h0Po0TKLHBy8SswpL2ROUHKA7uD3KDNVPbDGIt6NGVvf5kr+rsBb
LnNR+JB5uTlN4ZPV68YWFTSDf+TbKFONxBrhiKRgI5Q3poxm3BfLWoOGHQPK9alb
Z1Yfif8BhH+XwTHj3ee+lRHuz0auWYTEU137Np78BsBLaW//Mq/7nl4A5gnAFcNq
Y76OBeqR/s47BCv5N+5yQJMIOlEF4IMNHeiLlVUtEVpAA3TdJxGQsYyyvq5Ckaiq
LL0t5X67SQF4F50YhheF8HbLOd2/DrYtpJNU4C8w3l7luye+ukxbM9r5q2dFInOl
5WK5VMumcEkhrpoXCAdxnIvk1Cln+0SBE574rfg7E0xf7cJ++DTgiBD0xKdyFymQ
vabIeHvCiaiRx89Jd1H91UqDHtiEiL9YPohpXr2svH85vDnZ/I1l72xOMv5cZnru
ZVvPSri3dBtdSSzL9DmuzbuNYIFqKLESfj1hu/vtl/LsO5vzlZQwELYLdDcwM9l0
xhiqmird1+Ng0jdJCuvLO/fOf2Srz0659gN6dRV+KJ6P2p6rMB2S3S5YkZ09eS0T
ga9xkipc7ND0ro3yhfpEYAjfvM8wG0apdUkIHF4lYm8KqQjnT2tEU0YT9mgF5Tuc
1WnalYiOxYX6E25A810JSG4k+o+3yxC9WmcT3DPh2MkohqLTZCIozINTPrhpLQyA
kpI2THwIH3CuI1FWvJ54NlnrLmzChMG0/Y6rI0jy7yjJCN1vMUBSdngf+EzZ7yX/
ZzyFXvOK2K3qDUeBMrrrfHqECVuDqos6XyLzzrwrJnBk5NhC8V/Ohic/N9DLCRnz
s4hPQZyvNbwU6xVztI0rVIOtu1RNUf1f923uf44zBbz3CN1+qJFYX+VMEf1ldPiW
pa/Il7LR6YZjmvDZJMO2BEmst3x7dOotosnXtpXAK+cZfKo1Il9lM5uTBP4u/xVt
SDkNbe16zSUwE3RlSoDzYQBJRwnIuceKwyWbVlTmtykB8QQCYEodT0r7XShVhu/H
H+UsuvaTBciQSOJhE6LpKyy1yenbsoWPihDO0WaEWFAgp+QiwARXJ/jV5VyCPbRK
L9+M1vVZf7dkjd5apBF+p3kp5Ag2zldzK3XvFugxKzX0GA7+lKTYKhFKJ6iZDzzx
Csy+0p9buNeasfXRi3vHD1XgcV/kU9ZDCYjZWmneGofELwbJPNpyUALoILHH8p4H
F6/35t3l2dCLCobMZ+xOCbekf1qxYeF7QiNQ93dhcxi6kCXCNchZQuv7dhhJUdO6
oZ/alX9uPZVjdZkyx3UjQM9dk4MhC3YlG0QmTC4xjyz/fBM8vmoDHl9y849dvjEJ
HUiEhqYevT2Z1LpUvLT19DC5z/l5T0sVJQXSlF3se6d/cFOk+6i09utxVyugwlFk
DOKRTUHCyMqE/XYc4lI3OsqYOhCA/1X05uWEhHr3jPAIRBqwoXShxFwbqT+vBz0k
Lw+N73nSdyxVHuSou/OT/Czduq4YyBAB+6Ikb5gsa9dDJ04/Z9I9tf29DKbI+BUi
IRbjR660rqQ1yBCu2SFbOXJWqiPP797Pyrie01iA9BvJ8oMvnBWrG/+udAO+RrjU
OLvrfe0VxvwlBCTaTrZ8gew9s4oPlSog42t+Y/ZyX3Q0OkO5TVHesrqqFqujE9XP
6BLKkXj6B753Z3TPzMZnThFOmesQmWKkoD/CgTrLPCHn2rqZ65YXdtbUW39op9Fd
LIY8M8CeLHFSshQHqi73Dbu/xgpRlb46CKyRVNA791AXDkCNj1z7tl42Yq6PqgA2
B12uOSzOvhqeDs6XxZAjtMWSEf4HpxY2seonxGlsBF2je/4AHmDudOcX4XoZxQTS
rp0YxsG6oxHExxllgme7IhRC1XbUyAod/5x2122yvjqheIDfk0fe1qix52sURTxC
pZ3ylTz8Z9QNTRuv83Cc6I/gP/kHhknA7Hian/z/tA5FcZLe43PZ6PRCVrhJolp9
O3m6T+suSUKP5CA+5rwYRvKVeYyOUnLMoC4lnAvWbTwvzKh45bzcVgeFSZ0VvTzW
ubPFGaiGfaujm1h3Jg7ZIpvhYiqhqvxquTbaLJK5rxDUMjeNV9K/tGaC0f5+XdlO
OhcKBQ28zrBiIIndOtuOly7Y43HIYp30ceVEzoxza4aEcLtcMTYErZ2OjtGAH7Ld
i1UCj5l9PVbOaWduYqiDB1KeWu5YiOcEIiSc4sQhSxk/bYnHFt1+Ts4PMzOub9GO
yB8Br3SEd/Vw5UMfuw0hh4oPzfMqqZckLZgBMLbsS7ZYh8XCGm8Lo/YzqwpY2+IT
i9C5eFo/z3zft1CcDrp0OO0Q+A1YyRKx1rzlACdh/JgNA+JCnMa8mePTF0INZETh
4vNuy7ZWiK2OHlO1YUO6E7Lkvdbhkqg1Va6YYkgKkzKU1fAehka+y0BbxnLq5lur
79c5Ux9/MG7f6BSQLzzH9KFPkZYnVn1GWlTRBtE3UESVwT71xyx1z+up77y7f2xo
VYI8lBNg59p7f6TzfJRACk6RDZaxpSGYU/ivkcVbgZAPfUj0mykbpEBDmOXgGLSC
nPXuVX/guMjf45sznA7OAlNzPsulZppVb+GTxMe9r28MfinuGpc5yOWImEZcrN1O
taK7AQJCOy+zbBO6CWcx9eOTF2W0nBNYOKtzrGlgPFFuMzHL4Et8JLnPCdwQzyoW
tVfawFWbN71a7M4Sezf3Dcpd0EuGasubNpVAKxYYOQuDrOjD7JubwdzB81ZxYa9a
5aq2wsqr5m/EK4vAMjJicnQfuP68ljMlIboqrwrvZxN9CXuFTOeBjyZcqycqLzli
LbkLjzbo74bbOBPqxd2YXPuYeo/eXKJoZEciyIvILK0tvonv40AuUxGd1doYNxgm
B6/7UngbJRoErZnG45N5Kpdogx98lGeCrmm80CA5YlcUpsUrYG1te2dhPFdOvyd7
xNV8wiijq80o4nETpPD6YBG6SJ9lS87BmdBdq+UBIROWtLUIrJv4dIM+XxCZcWna
X3RhjIsLtxd1AJK5bZQYW2d2Lp7ZJHFIoh0ZHLLnWkMwbLrKlmm4Ru8x3xELD5x6
O1NDwmng2La1RckrjeTI7/FgyD8P1J0hvZosOoFmT9kI1er7ADrCtt+vUsrCvUZw
5COVjbkNCe32Yb6vfcVNzYMaM8gDwfz7NJySVwF26B1iydA9JLBeVoEmr2tzprcq
RMn+CaXtX1IUP1F60mKUMV+qCLV1czMpjuLhWdXA80Jg1sWqO0cebbt7NtVeqXXQ
d0XtvFobhzdQwRsJuwxhbiU5Ue6gbRjQnAnAHwvskD5nhtG2lFDliU01UD9vYIg3
5ShnniThR0rnvma1TQvdniYUyFuhzpJNXGaVkX2Dn8uDpk/G7add8EgKCQw9VLNJ
l1b0e7J/li1wbr44PMsBbvPa9kJ1t7Pnn6l9jYY1iPO+zmzpTWlwEXbKZc/XMZcv
2+Jl30YlHjNCXnWqrzvD+5jnb5aXOhb6IJhtDc5nEtvf4QYC9bupTCJEhkSVg3VN
oTazDsa94EWSMDpgpzl33SzCePQe6S8eCqhdFYeoKQal7scmYJUhduAYZdxjNJqE
/yMUUglqxkxA8sXx9Bu5kPSacdmniM2tL6hYEyLUtO00tzPPfjz6dltKcOjHXOzc
sMqtCTBfkL+u+u0XYBB0FeXv5m+89Ola0HvqlwpxM16+Gl1h9Pq3Gj4c2RRe2V8K
Xd8yRjQJXMaMtgyJlH+N+jveEYxgVrRkFf/JonFKXEb1YYYi/MIJIUUAN8xldu8c
r6gpMfS76TvxP6lfG6SMBkXVT9/jo7fuS5Zz+95yusOu1RE+UXhs49Qhqu9d5Oxw
3lgBHJCnG2H/383n9xXGyOQyAoAQueJQ3ebpp9aVB2eNgSCLBMlVKOckPYOBHcPx
V0fmTfDShPGUJWLg5RFW9ELpsKhcXeiWT88KWiJKCUULzO80mwgF220SGOGFcZ3P
1wr0SYmlZYecydsySQvVsACdpElJM1S6DcASv9mzlQflrh1nT30C6V5Oo97xZYGu
tGxcL7XxHQM8YXFztXzRof+HaZMmo4ohdw4KQxSPT2ltHKQwyPN/XEzHQq+mR6pp
sDl2y/Zrll2DDmYTjHHQGKID85rPUKz3C0ukjsH7JJeMeaTz0zpGH3jIdkenEPQy
EUn4sUBoxDAjftQrh7VsmTmLCk73O222bfwBQOCWKGzmG+da2ISlppmNN9qOQYrz
ObaYQSSVEGhxPlV51fz4FobzP0ZPKlcAdefDLHg5NWcT8+XnOGNK5DCLTpbw2LHh
bm5jGAP5IOTt/kUDyaMY05aElLK1p1B0/eHeFgq5kixFCXBa31CXrRjHJG/dQLur
rl6JwQnbBsdF75+MiXZ2YHA1C42nuh+HKY/Eg7NSpTQzAlUY7wWm+isdj+IdG3Z8
XjQc4kfvevXZzsPlvd8TXnbpeM5jHaVueWEBQ4gqx9mrRh1eyPenXKAFIxbvOCb2
zE4SuZ0QcDZRPYwk1EOraKcXJAmVFzE3WodihWCC2s9bSEKBfLAQqraaZa7nseJ/
kxKrCBAkwADZyuVw7lApWl4vuOb+1bsFVqmHvZzmQFi/EYgGP+tngK+gFxoPHCsk
YAIh6rdtHA8CPx3H3JnbbXV7wReC9IjVvpTdBSuDl51xGD4RdENi84bDddBISuiA
0cuqmT0yPpMrSAKmGp6pvAlkcYwHXniasBINc776mGS1E5Vv5YPSBQoXxzyb0y6T
zUywGmxjJZMVoTkVwq231NxboIgb8icjg6LYbxriQpkjUSgGJP13gmGhINoDe9Bw
m+SA3Fy73Zg921Ib4CuQz8jpSezdv5KxyMYLiVUsZXRrGLP2MyPGxokBY1pVGziV
TPOaeRfvTnh18xWnzluQMwt0QgSpVPY7Ahgs8wRlVls8lcyJrxbdDXdOzNLSJzUn
gBwcMWHKfFfP5cs9/7ltaB0hgQ4FR4BOF3Hj9EP1CRKv27mguiXPKwv92dnuf5o0
Jum6WVZMETsS2ZvnY16DChHnRNTlWYaq5ShO/9AuPV3scISwgCJxlruMOTe2Iajl
hK8G6AZRpqx+gL3spYxTI5D0Yjto6nCriyZ0D58P1VEtgOsLFWxQnr/wdP8MsKvf
/mVULOK7IBpSs1v/6WbX5TyqUDqg3M9ibQEEY7DdASN0u5DcN/XfHJv5UHK3hsjk
Tq0vf2mzG8qwFrjWVW3TioZoKOpy+C8jAuJ/IZvY0vUBYoDVs/c5E/oak7+4CBwl
Hcf2wFhtJGHYTfjhf3zTsuB4JAjIgMOScHb16gaXfHGgM/XmdOlig4ziFGH9ey7T
PLHsVXD50XO7IaHcNmgdXAFxTmPe3tuZ68s7jjdULiCUMY7Rrgvtpfa5a3R7DO2+
fZCGxdx6cty0H5WVtSU6/Cz8tQ7NCWJia7ETgZM+B446cbE1NtirIFchG+6SR4R8
2vD5YKPzTqlmEmF6yp1rmFEx3xzssbyeKcj5XS5ltNhOA3zlnANTcPy0+MM3A7vB
9/1q+gE3lVgRc+EIhDMl2iu6jQn13yamUL1rdb07s60NZXz7PS2bz0ciKYiYL6fv
zHFCg/i9Jb6S5Ka95h54ebP2jWxeveRIN6FMeTcNf62CkDmSyF65+CLVmu5n/onX
DrvduRKg/MKlEpSXR8kfQrRiV2bud1MCyZu8+lrXk07UzhvMxIi5cdLTzMTvl+Sz
nLIcr9xT2J49RdxtB+ZpgNIQ4TN2huDf8lztEfVXSQ8SDcE/Pgkylcq0p34tgJvD
0RL8t27JSHp7fv10alM90xabeXMRsazyKbGiv/+eD3V9X+U166hsDVnReKGxPHKT
tBvdB6kB5LYOdElbi62vWnHVlFpevqT/XJaRbDDJbcdDCViSiz+aJgkMPbdv3hPM
UxvSHfVOuPKb75FaCJwDA79r4iQVMfL5CEI14E3GydeYwAQ1HFqnKAwzCwAzZIqW
l9x8sKd0iGVZflY8Z6fABsI/S7pOln6ebcOJw32wI/0HbJsZGXnJkKXAYMKiGQH1
eoQ8S7rVbkjSPFxTRnXomrcdMNF8m67SYMIJjkK9l1mwbP0ZMrvwAro3n+R3NxA3
G3/RNjPtZ6eT5F0MyTsDcaI7mI0SEKVgy5YcAjXG/odEPH9/rL9KcRYB+DOPICCY
DMgLy4IV/kYGne55ownVf6Cpdt9HgSWtGcKmxELFPZyTVLujn9lTq2n9TFdcCAnB
jPAoF2iuzBrw4352ypN9pIOY06C1fT2OmsWZY7Wp0EV+NhBLoFtb1EwAIwIrfVdw
ip9QPGSQr5sxZ/VS3zxLosv15OPqxYVh70KOEer/wEqYPSm03CoeBF9ivurOC07j
J/mgEplfZAMtnu+uEVPut4Avc1DzFY7Z+JRy4tq9A1oMK0mGOcfffqKgEXwKtAcB
8J0WVP5Myt62PVMlm4AdAWh/oXJ6PrIPTxkkmy0A6CcEaVJVP+OYm7Tjvan2I0VM
4Zf1tP3XcJtGpnPc1nxuS+gAMxXVi8/C9DxuRVu3HRUA1o8SY71Oohlj7J7plVY7
3pkzAeOdYLsMdsWK8zpfDdDeqVlcUbO+0GgjJTBuTBneW4fmS9rFjdYphyxviRa6
A3D3hbeBnEH87z9iNoEC9l3yZzgfW/7qXgRWnXUQvqwTh8f6gnSyOLNZhAZO8bcF
Z2KM6djTkciP1LZWs9diVgNZHtzPBRtXdF5tXLHN8IjcOezancb9Ldphi738lgry
dVlTkq5xgTCTkqzo6qOx91Zyn5Q2wP9ySEyiAWuJCByBm78Y7vlNNgLeWlFoGXkj
xaSamTdYKXSz8d3vV1XGE7IB5bqRioHuK7P/p5nOl0S6eAWhqPHKFU2bVCV0VQL1
WDW35j+fVtC6D8dZKORxQvN9gTP3BKM7VUH150MoIpq2N1U9IMzL20Kejz2RaMdC
WZEfKhN7uizA7rd4s2/3ep9FRmZ99FGpx6/e7ym/SRRfUkYghWYlwQ5sXJFjuiME
mSYCtfbyguuBizkNuMVHm9ILHS9qCKQ2Pfx+LHFcgHbDR0ipRwQ25rpoOv+jl/Gc
Hfgee7iNuN9PWLB2Ngt3noyv+vFqpo8Z1q6WsG7UwPq0Msogbwyu/DoTh111Agk5
itRqM075KWUv93Xd8Cy3Ff8h6Nz2zlgzhmlKsoZcYccAjenybPsbW6PrCDyh22Fk
kQy/sjHDq/70FP+S+2VxbO3yuKldTUUf2gmySCswS2nBbufsEI8NKf8Xvp0XX0mX
4JVqLKTIr0lwmXr0C88MBFEStrlpbQREcSaiHGCWB9y1HIYOPA9y6yrZb7Utatnh
ix0O6AuJ6n9q3XSBiG6q9JTbsyK9c96/WtbPTaPxPyU0mgCMQGsC6h2tTyyPP2By
/Tt9GgoqAUywt0byfzMW867+ErKzbMsfSc7QPC4bBn/qfnW65bN2CCgUqyhofjo4
6tGPDBqhZ6P63Y2YrfZ6v9LkslftZAFe/0hgIa9NRyBy65IgSjv5vD92eWi0wOkA
O3pdPn3BM1jJz/eBrsWCeuPocY+NlDgXHRm7dW6FKsbQfciaF5EKBpCzxeeuy6wA
PTa6PM5c8+6mvXl6TZ4c6kDUsYyzeRE73yshtbgIwy68jWxXhJ8GpfErsT0TvvC6
NjWjFnQw9bcNgOHEVzXX+w+yXIJ4pEF/J+DJxAlsd0d6dsu7ZbbvKkgZtzVrtorl
ImWje5hk9+etHtlmzRn1LT2o+uOr6hGfWWYIISa/Nsv+e8a8Ixym/ALkZh7+St40
6Qik0DDvqpHg9E99eiAv5cS2WD58FuwApGrA2wTnFvIWeqFxPz1+UUqHAxL/iZ9J
rcbBdn9y3vY1zijpt9IfK/4jq4n7khTevk2cZte82acAv2dJExfFmtxhv2+iXsvA
/tzT2QWkOFyIdlLwSvBCDlblatZpeGK+Gm04Yhf7ITxdI0zLpPKEIRgYaA+pmIHf
XIgSOP/D0RUK/Ra2uLpf3t4zls9vlMPf1TLaWLuQGkflJbPTnCcsgJdKdgcdGfpF
FObfBsPO54FHJc4HO5NuedZvU0yZx0gtE6e2WZPCc0PzVwzVy5Dcc7Sx04CjM5uT
cOeSsLOPGsbjDmlr7QCoXHmkSN3SrRJsdwjKxa/F8jypAm6VJy+mE9HWLBiixNRG
UBGeOoUVZS/h462l4YNt/cnSzU4gYtaFpWSAejUalySunZAgVPh1VLFC23KccNCg
KvUskqbJdtsE8Ucrl+uF1aTw4bOvsmoKEtNlPC536v3Nx/55tvtN2se8F2DEjOCN
8G2ByPHxjwq8hAZrqG0ClrZ20HfGLE0twQzeAOWku1hl8c0U1eLYwE7MYNt14vn3
nErsqvYYYkPq0p9HuvhZd9XFev95S5M8qOmeQC75i+b/3I6T2vH4XEdzSWYp3kHm
Skkt1kZ/0Orjxg69l++0fzPcR1W3IkCBNFjl6kmktuGFKjwyVt3QUl0s2Iu4wbzE
jo9hLKFJCvPEOl6jTAg4RtIfC767phW9oIpMhuAn2jFNPhze1U/+awFxaji84DEd
mLJLWHQRX8rp6CNvATQxI/eQ7QUMFJdV4+VSrQd6TA6x9RtEiezO9ILDOXD5Gj2C
Q88lMSA2ZTEaE0Jc8BhSKir5pu51iCVx/gRsUh1lBc2DwdEuhS3julFNh3JzG3yB
mKlOcsk0sVpCHkeY/WBUzYEWYYI3YtJBX6ZXka875SHa5A9ZePxMShAqkDuPLZBl
RkwZI706qRpUIuRqpgGl1BWvnN/6JAZeOYJcfMD7JWsH/2IO+pMNvz+U9TQY8xC6
MHy1ic1g1kPMksFcYV/UNWkQrn7XMHXUfq0HZDq7l4UDszabmEc7R948wLUge3z2
wnrnoqQ/QSfBu2y67TRU/1zlpsgGZD39Hkjg9Nu8S5pua9JgBdVx4rdMueM+aAem
APzfB+liVqA2ubr0JDhBM7UZfPP7GuLzLQv9K1zVIVxqMX0GN4E/+bqZGukhKSWW
bfHAF2iNRFJusZ1s36cSnni0Jn4p3D3WtI0T2GZd7ORNimhRxkT9eYX2YFviilSn
jcFuEmmd/j2mn2xK0U8g/ecq75wY8zh5ncl926Hq5H9cl3ylIt/1o/s7gexXNfxd
X1UGe8jsQLUzBlArQ8sdLQKoybNc08AkELnv8s6yEAFr1Aa4Z1ZVIOBMOGvwntEb
PbKIcwrP70KTsSMQ00+miKP7DMnKJQwvQlR65KaK9FIw/u2tDTs968wxJqD+JsPd
DEDzpmETmpw3Vj9Q9h4u1JNpldCKDu2ksVwBr8HgIGYy0rz0bUlE0AVov8kqVHeI
HlQzdlQ7HwvbxR+NeZhjsf7TuuaJiPUeaSAouYcDu/wcXxfD4C5GDJ8/1CovEoSW
CZtq5pXtcZeLezR5ATnA5AYRR6teuHsGfF/WvE8aP3/jAoeW2Dw78W5hTzmcWrdg
MnTDeU8GEIf7+q77VgYqZDscnGgy8WcX8MJcOnljz9Ou65Hwn/J92gLt7lf9470M
oBvZB1Rql1c5EF8tPJN8n5OSjwBVqcyYlWkAqoovf5F4RQpAndzHGL4NGVHrnbEU
mhp6zIO449/8SHMrJl3z0VfG3f+BNtUf86VEaiGJ0VIihjASS89YhciSTeel0nqH
o//GTZxozLGx8FFpwc00SYjKRj2m2lWF4PTcitp9vTMtIOymLs02eDGkNt+hA1PG
ItfLxfy8aKHY5cWkOtw/iyEI9+b+k7wZ0Yr+LypR0LnHLTBO0XsqEYF/+Ad6XJaa
4i9llp0iaHB5pSK2xUsO2Iu7CEj+/ABM9WQuGAYQfYu85wY3JSdQk3KyeL03vPsD
3VO7DNMHxWO27QLqga5YRkBbwvPMFllwxDQWqtUJClIWjjq2SgkCWy0FZXg8Wk69
YuevZw4h3I3Th8qN6czuxPVmV4cJurnblUCwYNqx+MdMwvT+vTcnpEP+fQ0titHB
VIcMrziN35QQ2mQkskrVFYSNbMijpKGttLTHulbxEfjbZORDDVAkI+lq1gq7nV0N
ljI9uHYtOTCJ2pKJcEziaG9qBoFBhf0xGCSO7z77MFbRIKB3McqiUik6AnNjKBXJ
cWvzVZouYkX5Dm0Wpd3NiBltcaZenk6fvZd2CMo+szGxFzsNeblkTIFD+JDStCK7
97VWf8fVpDRLBqWGXJ8Z0CcfAxE+vx3GHXotKddG0DSwqh+bT1u+SvRkrZHPzYZU
3QRBmtdtg1Y63sCCirWOB6mJuqpWGM0YeFoEUak8ZoDmBPCpg9Ey7eJiZOMv8hVc
QV//a6uwNyTUiAbLs0L3xGYayhsr5BUAKuMqWtTvfavZdXszju0hLmM2PuBA3fiO
D3y5J6TayLXwM7ZF2nXruaLL/ptojOrtxCwVFcoeqUAtiMoL1n5Gbe0yy3cWGrjl
vBfafQS7R4783TtbVgLoIbA9lxxKSWaasPXFVLnxHAzrEkNG00FsRnyV7EGrgWY4
Q4CmN14bgyULZwDApR7SMyM9kb8t/bFikj3LP+1xDI51Rp7p+SLjNOWioa2xpyZF
7m9Fm5NT5tqNKUjgy2jC5FpsGqYn7R5P9Ff3Tw20DT0SRYlIFMA+Oq/9sAWyname
zAC4xKkhtMpnpSna7AAeAo5D8RVFw+HnYD7Vs5qbFUAZCpSoqD6J5+xr0TLjmsNX
P7xoag9oDaZ0gJ0btl7V2fODNRrot4k7vLM5ooFh+HGahmLq7tC2L+gNl8lXqddc
6RsdplGSxe9jrvKow0a/0PU8PVsy4Q+BS8LY95LAuZ2pSDlDvF2vu9ABLye6vVPR
LV6laaDoHiQDXhsPOu6vjHUSr1peZR0+AjjwJcFFAajrUWJY+4iN0p//pU8IIq0r
PU76QFKShlYID7GfAHDocMAj8YU4Q3MQ0oMheFx4Y3lw+OwYc12s0z/ZZv7nrBCU
SVjESaNT6KfYe2r8UIDERvhWaLXVKMteiTynLIfkIGtcAyfi8zfdH7u1eJB2Qxjw
W4MwnrpDOoQpeSpJGIf5WWqbCpNbVsGVKfSrEsuhdCN/6VlAkGzcUEA85XhCL71K
28HJtnaVVHP8GGat5RXjrxmUk01utN2R8u+XIFwujUuBeQOa1MjSve6xYhb/kSVX
h90GQI73Gid6UnG96vc5VsACJtB0//cjZ5E9VfL04wuqKI85MOxpHzyPQXcXHlUl
YksvQB1ktIMpzGYASHk5GolvsEW5kXVCLFELgmS591Q1qPwnAsuQGQqc0fEj8EYQ
OavpNRm6diLyxM43+misWdtUUP6tc30Tw+WRe8PMAtwuphNs1t/YIXXBPfst18gB
F7TCQ7q4Lo6AcwjWriDFWZKHj+bPuDVR4XNZaxASKdHanH8vTomYLJ5LmZXM9SBs
5DWN4pyW8AB7ktxUVEhjiluJuNrgfscQzcHwHHeoQYWuIMH3pAsf8lE/a73EYWJV
8p3aIaEx2qzPso5o47Jfo6Zi5iGXfkSVNgzM6tUovHb0sVaHbPRFV3mx63/yZ4Ym
xveLfU2DZGdfx2OEhSj10vGFIia74UIFyNA+0QTJ7sjfMVEegBfSCSwuY6FEuswd
sqWnaBcfkosXd/PdOOeJEn/CLvDNWo2ns6DtwtMlmBgNZR6m8N6QVeOqSMXam8fE
61qZ6nPz9mYWp8HPZvu/oRGwfiPnqbqbhjhAUovBd//rvG04JgnPtyrAn7eWAUF0
+dfaJGXhdb+Q1mnp4hmIVMEW0vGIexUxHHurKVxrW9t5sjPDQ5rRxiKkFb+Q7dem
IAcY7m1bhSPUZCjGe+WUQDMmyE5moVj01aBmiYnrwYu8Ee4B77KZpUBkEqFyUe/F
SEj4ceGEyVFHFn8wChoQ/R5g1hy4r8RZbTh+cjV8u8LCi3xvDCjSMbSk4mfTky5y
8yQiXifEHCdCc9bTnJC/Fw2um7lm+BdQ4IxwYKYSKOdoCSfAyd2DdxivCYkmphPo
8vsoAWiXgagbQkdZxurOcRTEEhU8CS5sbTlHBfrKqj/MQZeYbbjDDpmrjEy3C0CB
4FnUNF89XpPMX8HsB/4v7smb3GDYKLf8eD7zee/D67qFMsFL7snEB/T36N1Oq0ym
UVMwOgnjYolYvIcGiIfqHp556Lt8IF67HUEQGQqxBWz8b8zVcfieml/FW4QU41JN
BUJyqTN0tDJpmuNwL8xnBBmdL0nf2xdkBTQIGo1sGVGc7gyq88hQohx6qnftjHZq
/vlhjZ+Xy/+dea6u/PcEnvqoxvO0XzJ3vKYPM9d4EO0DUm1THCT2aKdcEjr4QN0L
XGz6mm5BHeFTnf7kXmLBCi1zW8bwXrVZ1HPvUjyc1CUpY0dKbhG+hGW0c3lF31gW
RXgRN042Z8m223difhJb05XUGbjbs9O3XnbTs+N+956N8W0K4Pd3ucQSLiOnzi7C
yjTFdSUZ+AjKWMCo9LYLroNz+RAr7lyEX46tC+bHVPxkfKWbUjmIOucjKUsu6ehG
k42J6VKjfyOcaWUK/E8M3oVE/8HHEQgBT5TeQ1NXNzGPB0R+d2PewKB50EgTUcQO
wA7Gc5z2ycTj24Rg39SjXyY9mHk+vA2tRudYuoq5mk0EzP4smGododWeyqSaDshs
UYmtENzkFE6Ffhzi/ePewRW0on30nPOiI9SoWsVHKrtuRtzmtG2egJR03W6shCbU
vtlxNRQwoVQV+ItsKFC4V87WilQCKt+9LgyAr2RwAkExrttzWtWL8uBd6QtLAYFj
MbxXFq4jC0x8/lWSB6CD39UuAc9YjeHTCnRHUOeOoh2uygoHVrzI6poKKYowv1lY
evepnMk7cMt/asVJ617TTnSr0BIw4S9ZQGl5ckgOEii61rDhvfOIE+pqC75XJ9Cg
kUVKp985NYVUecm8oD/+cZFSuRqaW481PDIYCRGq7IUMjOW5LyBUhVLdlvS/yfBY
MbYYr19TLfApOA1DrJPSQrL3a0CEErPX4WzFjqGukUgPKXF3EHZ65pfxLeKmhJXQ
IYo5lVWR2+CjfHl5k3RY25n4isuLU2WLONIQUvJxZMu1D/aznykAUxpluJLA1HJI
lwiS7YBS/FZsL4hV0w82q4aXoZb7A7rTCfCy+n4oFGaTV5APpLl5O4c2XyLi8wDN
cx9dgSXLAlO6K10p9tHSv6NLiSpkyQZNHLoy6ZUnldas5O13KQB9xHBpYLloGM9m
2Wr9fmff+2nG9HxBAdBTBmI6Sb2OoBWlhZu/ynWhOaa20/kfmLa5cWufzTh2+nuo
hXiv7ck+CqBSWh/hJuc/BjIiMyjuDgVZgqfk1EqRaEJy0M+LSE3x3e4Xwd3SgaCd
lU1jDHp7Yem2nN5hcfnXgnsQgHZoc59Zz7uUPuO36Yp+Y8kSJh74T75LZsFvVvKy
ESOE7qAV1B+DCz5nEi+Sa1l0uojhDKOwt08pw5ngXJPhjiw4dVcVxd7zSR5BPxet
qseVffKWdfSFqdUnrYCiZdURgrGVgh/vMw2UIQYRcEnyfeqoBdTgwSqJqNZ4DYJT
XSSltmXD13Es/GQT68Lea2oAAD/1rOP8ZW6MF7ajKyBSrjWSWVRMASDkx31HPMf9
QT6CqyWcqxmG43du6d3hizpGiIZEAFW4C6KOyfgIaX4SZEcLdw3fiAb5ttRQxKKH
IzE20dQreKejzAiAIdxdbzx8bYLyUhM/2+StA0OIcB/XUx0vyscjQ/p1pYFn6p5R
5sUnOrmjJK2BelXtZ3S7gMn5GFAHDmPn6IBsU30Rzk9+WrEVvV3iyUvuBTdmH2tD
TG6OKzd3UHAwr+1FSLOdkRcWLmewRImDi9MdNDNDvi4NXgRBErQhHNgYvwL9sWdm
i1uf58gC8XXe+iG3Uz+SokvodBeRDBb7XXyZ6/9lq7kheOjfppQMKC9/jSjGViRz
NDTHJ9UO+xdOUjpxy/02G4erGKqATf+ZbnrS/vNds7hZbZn9ooFgzi8lqCfdAm3w
BXXzVZwM7HHwHdjFtyCMSVDte1ZgDKfg9xSb7dnxS1R+TU3a9W7XJ6Nn/03Gx0ja
3RFUR/CVwNVJrYkRk3qSp2nxt5oOSuo6C6qgN0f1fuXWfezVAKflJQO2G5P3SG2L
9/CitwDGt0L+V/oQoDCdSwdvyY9Op5e4eqnHrgq2hIXK/r5OCJ08YpDWEEdd0eB4
VG3CGdp685qXrtx8XhtbGrJPN18Kmo6EtHZ8QJfMdilF5sT4k2H2YeMRZ9SyffBe
8wFiHftP8ZG0tb/pAh7R6ItENR62qS8d9vGqIvt5w3N9iGIcdJxfX6O/TjLymgIa
0F+Oyx7qlo2gpiUldtds1XNcjfYqQFHM1sGZVOD8iv66Ip6MoWip6Z8zjJlLPg4l
w7twdvZ4medFjZZvZd54fb0dnydaIxC1msdwBGEmNp0nUM9d6P6yYtvlGh9Oa7qb
pAlyGmfNX1ZZqvgb1LijKavm64teBEFD0Wi6ao5knyEktzntnJEaKc2J6MD5Bie9
3AW4AMezI1HFxblbZmvvoub/rtoUu6RwkRkO8dBZ/cQWbsK4TwZgMRXZdIYuMI7A
I0LPXCIM4pZ0Gd3R5kjxodG6u0HCkTipzNEPZmEqjQcztUXrJvCcEvD85Wg8g/xo
UTiFoLZz87XIJ/jwr0+N2Yus3LOCucbbjEjbkhSldQymOHMjfC11ZDjlWVIqw1eW
MQI1F45mVo5s7y2r4KZODGHRFqSah1hWPR9faWkFmIXVqehCH8QgveDz5MOVFSEI
x25OgyC3w5ofdm7Fpx1bfLdLcWGdVrCJjEgTgmzn0g+oLRy6ZLI94MGGYq8EEgMT
kM62EmzcXgILX0YpBPyiM0z3C85nMHnr7TQUyNDBYJCf09QKs4B5R3ZI92fd5RoO
dSio4SS3HIb4UlUXFBbhCrbabjgFKv+P+HxvpG8JHZN9E6gbPMYSMR4lygAYsA4e
zmWDETEVUUkT+kr40CczgEXESNVtBAOkdUYBaQUjOHGWZac8yL3LnxiXHsDKUxbk
kls5iZh1hoeyzyhi0CHLf6xviAo7/FCiU/+ETO3vxQWn4OGqquvG9LyGHRsUChPW
6g/5h1StLcwqjMjjYp1Z/Grl7zH2V+OV8NSPxvv/4EV7VnyDh6t9IHhzbnxCSaeS
0QJ+AQ7RBQOp6yc1uQavDK5NE/BiDHbcWRrp6k77GKKGjOA3Csawb8eRMQmrKzny
xVAeC5AyK5YTJO/sk16lZLtYW0yR6rlsXQzfpiSbp1aeIfB2PMKAlRhToGYhcQ8W
6cZaQqiVgWtwuA8HxgV74YV48xkPG2oUx60q0HNjAXd8asj5jm7atq3oBcbvt0+g
gs1COZIHRum1gVE9copVg8YgJAmgWxTlQlyDaHIjd/nWPO+JyLl6fBTPXqVLNL48
0aNrOKEXB9swepdCR5ouarspA17gcR/Lf0MLUIL9Dstwoka4jrSd9A2u2WpTfZp3
pywzosMQ+yyxamwVMasQa+lQbaa7MvyahRkMOyjMxAEOqUv5ICj/Ellvstj+EAOq
Af7pr+gB1Tup+PNDMZ3odNolswAuXE+oqPlGe0f/BuiQa5lEAkf+vghAFH2bYsqP
0utKzCVsOiN0TUSuksSQLvsMSZtz+5LeH1HdJYQgGIiEOT6+pngr5boElKEyfKJM
ciynWqJqYwqmknYMJG5CAkEB93QRkhUz0auMazKJFKHf0kwhzMnJYnCy7hvFS5ou
iniEwRw3H9M/7afpgpv+wXbF24aruhdWPxOJIwSEvee2b0VPCVIQ6XswBeRQD1Dk
2KKHaG+VdOPwE0hZDhUXye/8ShVuRk+BZTuN5c/q/+vguzaCAauqSaW9l30m+SAy
SNyR1Ovs61fDI1OEEIGeIbinv/+l2A9B0oLgutv9PYXoI3RVSAnS9+VAlmk3ydJH
002UDywuH0/xetv6R1hw6FrKWYezBe8ZJMHS4qUPdlkNL92m3jnp2804abJu+zbD
O0DS1qSiR6072gIfeBt0nze3SZJ8qw1+gNEdBxyVkBxKf5GCmPIVEw7pCD+vL6TJ
eycxd9szxeN+l9al6mVPbs3BIxLqVr19iLR7LySTo+iOws+PHljRNtpQQo0AO91w
bFahz3jsobRMD/wjF3Pr3x5ZmvAu6ufZX+RG0K24ce9aro/SwsiQhJaKAm02p5EJ
m8OiEa2OYvDp8ttwOy56QyhlRSGw2qZ/T2lTmTZTwUFOnIQwPdpIJaBXaCm7TY/B
PBZYjykX2ZSy4HE2EMUBcYI2FmXc+KNMqPZ5Ggs7pLrz/VR+K3jJ7Kikw7ZIT0s1
ziPJSJPAy0kbwTiClyZgGP84zekECQKZDM9KZCChjCOpn99+0/y+5F7PTEGMBNQt
6RXZoqzLOEpJH+wpmgMkqpt3KJ2DvIdSdmkiVpZSbs6bOhsip9oV18fC3l+x0i9e
htEcwzzgzHe8ShTlsyj+A6vChbsAKRQpBLTGN4FkqEjPkmJKBWCy3YUxPLVw9VLg
Is9s0cO7mzD0g3YhG/nCCNGzdM9bDLTyvBbf6QxPgZU52BBhtCO0itTv0/fWfI2d
cCdQuEuXh6Z/Rxjcjj8WlhG7hzyx/MPQL6rgMDEgxKl8Gujdu0L0QFNjB0ysM92I
Pl16Xjly1b6Q8GynWHh4ZpjWPXYVelioum1p2sE98zmZgolakVAR5yfPetp3gEYW
DEA2ica+ltDvJIR0u7LCW9UkalCJdZM/t8N9vbB246L1tfQjYj2AfVlARd1PC+z7
0qOeie9l8TbmwMTb3sltBEni/EYRlMbXzQN7VDI4o7zajgVnxOG7983EVgXh/vEM
GXBwNUJR4RFzYJHgIAICj66lhBiFEV5bAwSSIB+MyxehXj1qhVvZBzfevQMkDmAH
+bIS7oI96MJ+OYJBFy6w2qnvjQJ0tMaiPV3UMQBHPwqVSct1AsvBqCpjB/MzOo2n
T7TWnFujq3q3SLZdtTTbojR3wAUe5mRhGSSHBkBg7vGyMXg0Mi4NjNcTPqFqs4vw
HooIimmSqGMEGJDdOHnHmdmYrAvlosLZX3M9ZQ0F84BrPkCS0hUQVOVGMUvjQz5Z
+ENo2fVaLYx3d6SdBlbpMHUWoV0Y81ScEn77vXJZ2wWA9ckdMKbE4SDR+qCFFrR1
Ami83c+bWXkqxE6IK9oxAyXOgb9W4bYcjE/0CHAqixE4W+Hmc5htHa3AyJJHnzLS
mLF2bGcKK3Fr4DMDUFDD2JMiJCk2X9XN9fR8/1schSPPw7d4rUznRT34oqn/By/A
AhViz05fsfi78+tLwl3qpreTRGeyzK32/HywQR24UeNH1o9mzXdSNE9kYYWg9HXY
AbK827Fi5jVAFdCkCt0S2sCn7dkO05jVAfOjqN1VXXOdXLT6HzVZiuH3U5b/5Y4N
recy5w1eHrJJvor8pNLVfx/CyYjgx5fUHpLNZwJ7BEHJUk9iZ0np0uzEnK1uBkJE
z/KbKMBc9iN+gU5TcqIiHj/Vmi3WFzsNwpf/Djo7zWN/ifBnLqg0AyxJhuIwO5Io
yGh9pq+dEUHWXa20CVoucjX4jzgtPtQ3ULSKD6DvIMxihcSRS05La9WwkCIt192r
oY7siKyyOIl4rVBGvt38ty3KQamdDAEk05Vb0C3dKZR7lgjbqlB8kT494sEe7g7+
xzawsXO8B/5qDb5FDGdbWbmA/8M8qXEd9JNzrSxwXQrWiEYzGvRdQTQYppCNaD43
ykC7nF9X8v/zlS7u8IU+R1//85y1SMUb5TtglJRyEOFnVWQ4fI1dVU/ekUveDKs7
qU4EFg/kgyIBnqdY5qwkiGpJ4wdBhYckJEVrzsoKvI/P87dvqYAg0D0BL3kUAi3X
rzItfU8RUieUAhnYgr8pbj1cZYk7tIdayMl0S4nrT2puFTeSVbRLoEE1hZpZOPa6
6qYlIgf4x6TY0GGB/lY1SAuUn93CKd8EMbnMQ8LdAk6k73Q5x1o8A+oTQ7ik2qhI
hDqe+QXK2vtRZoBI/ua1X4oEf6K/554mt4OMRmbdRy4hJR5HR9D4J829fSo8mxB2
OWc3ltKTLZUlDBip/6Nyf2WK6bIDxOIhDAlDS0DxoQOjzu8FwyYVpNvxORCohkva
H2jWF0yTWGM3uJVkzh5++2B5psuJa3csw4mfoi3zIovRSdW1ezp8LLOugsriinxT
PVKJVWqQElI/ybmVGV8vyO4jr3ThdiKXuwyU93Pw2bK98SbIkOOk9PjMsZcLm+jC
STeTHs0ig3g+m9FQ2fU4solZfieHfOgQQyGgcQifs8ywD0mihPaT0WgGTJzSab2l
vdNQM3cBp0I1EEUREImCt+gIb6wgoAFOuy+RiCK6q/UHycODHXetuyLEz3tLeuh6
c92SJkqV6tcAplSkcfHNGF1EwH3woBOt1J5B90X3FDfDLF/WUKopXLTArl7uG4Ij
Nr43XSOANaIunpy1GCuRXFoMfL8zatb5KOzC7YsN0yN+Hxqbe5Sxm4RIwY40cGaf
TwV5fANZjEzd1qbBYwI7mTD2FHj1UF9co5mm/TViJLZAATDqezIxZ7U1BO6vJ594
0XGXqH/nvILzFKpmrcj1q5intU7qvYd97kQRhtcX19DyNVKAcEK9Z0p+R56IelPV
dTq7HORFXEmBZBTCRMfadCiTRX81uQ29GD+W86KEsI07rb6BYWRpI5xsZN5jz4Yn
0qUA7agB7Ff2w+FD+z7q6NxvIIXg6uKWIHE1F85KX0d/nSc9zjQPeBIhWtAFWCOK
IsESMChkMIWb42cOv60XchrLf5D85dSImoDySAyRFxo/Ye4yogNZwGINyuywcpmB
fT0vvJdmCRey6oEXQIa2F0eQX+SsR/o5byBGYQhO4ms1D4uPrx588Qc9Yx/tSV2l
pMg/I/pGIh9idWh3m3sTdNhr8qoCZ97+mZ2Bp9CV/uyEEw4MU0LOAUD2KGqT5f3+
6R7S4agHz3sH6XX3SrxGvi+Si9pJu3K9G8KE+PixMOW5qjDD5pBd/DQV60xRYTZE
v+BwIXUyBeV1chRQ0p8bhvuKNCgHBnsADgs5I50+Xmqak/3pu3i1+5E5kxdu4e0Y
oQSfJckEU0SZwwEJVlYz9z4ENUO2x12dREccuSIQAhYIug289Og2nd1tma6y4NtW
Kh4DBwvL71zlL9sRnaKn2jVMG03zg9jPJJbjNeirINPU4F1YBGdEUldK5hurMy4x
1Ewwb2Deru2d0EGgqZvrgpU7W7GhojGHeTyEkZpn85oQAYCoCCgcH0W+TproJtie
4FG2JMloYGoaQQUJhfOkHAvd51nwbJfr7fezQJ2XpP2+htV3+1wy9CDB9eIj+p8l
OH0V1ntruJZNnNShqltejSdqzXQtArHempnDrCyLL+NMEIDxQ8QijPC7i8xCjbjJ
gndTq1rodaAitD6dZH9qe/7wnBVPj5mCocwza7dRIvgDWS93YZEbL3+fjvao7AfN
jftAhbxu9peKy8RqwMGwfbFMdN8d94k1oQZx2bRvSKRFAOatJ64C6VgveW18tUwB
HOUPorsN1u1EzBm+a5rp+DhW/xBbnknE/yiA00UJct1sq39EOBjeeMZqXMfMkuHl
TotYB70hpn4H9uFzBVzgXNb0dgfoGQIoNT8EhsNFxjQl3oziF5p2NcE0Tjb3ESn4
aBeNfHAKaKO78HxMgR4VpE5hJHo9AyjUFfAEXeaWazcF4zVqCGUYq88aFhiFKbrm
g16jR8N2uQweQacYFQIUaxCsI4+87Ek1ktD8I4M9mAA9MGsndX3D0PiXnDZqO6AD
B6hpCS6bnKrK7HQr+KA2iwYYCvxUV7O8P/ajaX305nSXVZtVwVzezqyONgs1wIxE
lG0yp8j/LVyE3I2A2Xii8fXtlvibAM8RIG5ThlTex9M7Zhkr/6b8JzTVfh0DAFWH
bO0WcmamzsA8Thgk2VWWADrwxv75ZObOShsde1hYOM8yf72mHkBWHyP4bM3HbFaz
scHFNud5KPBsWgIesh/a+aNrVdD/sR91nLQ1jr56QvAn1nlgV+09Sc8YxTD2CcPZ
lOZ9ynZ1y0q3CHi3uMr7Kqvvaz4RdHP71kn2ai9wP9zVVto+BwPk1LwUdXG+C2C7
GZt38HPPzJZYelAepFopaAt6AvDLTkJ4WQC+iokjt2e7+B+U6Q2grhCIBWr6L2rJ
0FMvq33itC9UXEnXFIqfBQaACOCgJkTxcoOB+Qrew1m2EdF5nzfV9aj8NAoKfOka
1raHuY95+yLjrfHFmL3yNl3Gr5XDlg1UNcpXfWb6nxcIMWOA1iWMihrmGGKwl11o
vtWp3UIb2ysvXSQrQKxPEj12BR2xLCoHTUmRTY1JjJg=
`pragma protect end_protected
