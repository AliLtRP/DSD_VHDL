library verilog;
use verilog.vl_types.all;
entity ab_vlg_vec_tst is
end ab_vlg_vec_tst;
