// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OHF0qRInv+aM6bUDCl4SPMEKE+Ji8XTlrG/M9YObY2NUZbKIsXffKbUxF6ajpOuX
LNCvlRX+0l7tSDbAD17WjNX4YfkzTTnO43ujpM4l75OEdvYbGZ69GgLAs1O/HlXl
IniO1r1HYd3iRUNr0fY1zphy6KBG6ThSxwg7kA8NhbY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24528)
R13Xwgeq9qIh/zaZ1Qw8ZZ1+gc6SWQwtbBS0yLG5gns5T4A6awiJHtlIoN3xDnNk
CUvW/IJBqLTXc8/rATgJcuYXofN+64DTdQszmDgC8dxnW7mpI7inyPnTTIa9UDNM
DqU/RpQR6FyrHvCtC3zopf76Q/wsj2Yt6hKCMPZK2LCKqfdhS7TDQvT+J4dKjE3h
nNcgQR1T4xx2VfADIAdg8mU9dMykOLsZCyLMorMa2cnxg3TmAgM948xR6BIDuh9w
fzU2QyruXeYVWJaTVs02ryvZKgUAPhmA2Di1+Y1otEFKIYgmwcq+I65G3KicIoKV
8AWVuHsolhmXmUFQ6+z9PE2Xl8Yvm8SMYYqjXJSTTbpZKeQVBr6hBOigRX0l/YfX
+k52l0asOJTV/MMq4Pz5UEzYjXiNpLherGeGtd/sMb2urh6sDMGasYGeCmu3a068
eegQ1X6JrdvHJw6i1QY0JGe4U9kj4nmS5ED/Vm3EyYIcZcTHZqrDzez82GpJR9/q
0yXe7NY/bTnbtCOEsZip6zXBrNfSCeQNd/tNKhoDfmaZ2WQB3rj4Zg4w5l7eqvH5
eIIQXQTa60l2hwz0pG9fepAcOiz+FzPUX/YC7/5e6SMbSsYDqJaXm6s1UjWfJ/wx
KjD+h2g4UlNkZUR6ee4hKa8EtSvzcGMC6FKyqGK7cehG+hgOf5Fkd45goZhNqkF9
ibnd6SUAJmnPabWhY7hugkOxZK38VwqAlZkvWWV7/BmRqT6Fo/TTOAjJWhP6s+8e
PlODJJmxdY1yEQ3taDESRNI1Usl2JFhy1PObaYC89k5PzH9QWazHr8vXISWCn3Jh
i3cUwZyrvc6/p71IALwXmAXILS1fXLIor1Q5mXxizl/9XDJNFPT01E60UUrUZiwN
8mwV9v4sh+vYfFEABMFxPp9cd7ARtRQ45hT9Qw3myKtJNkgByaJuPOk25TfN5D9W
cZbPvBK0A9qb+Vw/xbIwN2unFjot5xYm20hS3uvm9mP+HhRUAqeEW8PzwE6HEJbd
KWpRr3fIYQfhOx5rs+MHGLGBS7lq/sMhx8fQ4hTLqD3oWQ/e0g8YLwZu4+am3+Yk
dMubLUU4qmFPexbX0vRgT5FYTpL7OcNUI2YVUJIPeYHq0ZLTs0HGLF8GyWEgS0Xo
LDMWfPEPO4ZI0Aken2XAqEwxDBAegiYEShTtnu4pSussJzVMB6UC7H+sppYjV5xL
9dcBgXq6J74vV+p0wHUamyIhtwmQg5K9quE4RnU6HLxjZVxDqPvimcPca8kN2/y5
L1q5ASYwOY0so68FloJxgrcnZ+BDl/g8RIxfyq2bu/bpEWT/1GphKfkTqi2MbQY+
81gXH47cBD2Dt9CACKMh6Y6LMr1IODs9O5jspPy8GmN8M0hJjAe9KPo3+YXzNRVC
N/1Urte0XFZgPi9j+xccsfTtgA+p9bZH1gZXHXH6XBsZt83rey88LEVoOfzhZ8SK
rGZ8uUo1bfqjZX8XBkqZksCMJ6MObyjNUZ6RafBJsMUp2GnH5cbb7aArsdNcVxK/
qdBj1siAuSL0sbWWPQr2h3ewgThGEmfczT/G7E8NDfQCCfR7WFmz23A0jQ3YUkvr
vj7vjDj/LSYRMEePnkZLz+YeQhqf6QBb8FKBmYA44CmbGMyJTaGiRUdEqVdpeuej
PhGC70+XLUaUK7zwKtSjLCDuVI85ZHMBKcixcfoC70spRC4WlVg/dXceyKF3Zvc8
mb3aKKaAAGU/YqjFE7VOt+BflScg3coyfEsKPIxve/G/WPXDcL6IZyyTm01NDWDL
eei/jeDTD/UdBl6ob5Bn0WUgMPg1XwWg98+0oehtVKbAbn+KUoS7jT5votXswLA+
c9dJ0RHnS0TjROcDtWyFGkUklAAdKiqfTwN+8lIvmzXeqYXdh8H/rVlcyrQS+jSW
JItB0VGYjuQDN4YWOwD26XZiuVmD2YA8cQHBYFQD88v51TZVQxfX9KTrLWbC0dpI
aOGwFGV0rk60os6upVG5Ra7wLJho/73YytXlDZnG7mNWzAtGjgwNpNL1ISUZKnGt
sXCBVO2WXzivXJ3Ut/MlQ2Tk4pUPOVQGNNUNxiHsRrO2zAu3R0I9frjg5/zxk0qn
+z6wQ0KnRByuVg2vOWSeJRFRB3MX5A+Yq4JYB+P2+tsrUaV1eMQ3DikWU+cpAYM5
7a1jvfI1KVCQrvbnsbRUjAwM09YxnwMNuaROO7BPBAOlApjJxUiZMsNW2pksiQrA
NJ7dwyXPwt0J35LKsUseQsY+HPhhCdSOkrGaZ1aYy34x9Zot8lM3L87EvItLxBCx
64/FONnSwV01jdkogmmcyLiWseS9d0l7JQc/qdy5zledwbr6P1eDwMUFUFqg2g3j
9P6FI/rGuisGpng7THYtXPcfmwUoi8S9dAu+dtu1zeObZBeHNfkagSGeAcNxXHIW
0bmUk5lSuxpgGgj547meKPkMUU92+vX4YajUnFgFz/JuDhGbBLN6SBwjWJ+t7wbq
VDWLov6/vUOLjqDH1yqztGLli6YpT3PDcIcgEWy6uAZjqQPcqWZo7p+w3oqvmkYo
W8xtCyefqPBhsotD3i1M6bXlVTuPE8O7p3Pu8fbBlYydShnIqAcGV45NDEEpAHbL
LXBkzQafEeoJ/6TIjoRnlUBHIJMaP5X0XbogxbbdWZ7KYKXJpuBJmW0TSbsA3MD9
CsP71uy6OByFSBIEjwt1sufuZdJa8EiA1Dx9Zr0nZ6hl9P5yQRDcxm4Tj+0m55+B
glYF9+/lwUrCjfBtiU+5jKI+vU5yHXw1TbuuhSWHGAd4ZpE9SEX4RgT55ntp69m3
SEYx4Lb1VfO1+uokrsXTB3yxDfs2SCrRj1tDc0Pg901sK1QR3F/a9fvNyldwKxPr
gtk3OM3Ic7nj48AKsgieg7X6ixQhZLNh7XuxCk3xG0ZgVeSoGTnXY4a19WjubCdb
gI3WlNEAe7txNaLilZqAbDanZhjrB/jw53M4QofEo2tj/pX/TbpvKmuOm7dVdvd/
UNPDnHqNOgIvA2WhcGSbDjEshTzbsXq/B73rRvn9ufV6OeATEmBaqgWq2C1Zfe1Q
pI29D2Tig8o9FQNjuTuUMa1zDa+3h773bV/8E3mKB+Mq1KsjnIHqReutkL9FmJqe
tbnd1o3V/OE4/U0qZOp/OAfYKObYLuVoaaW8uhe+F1pGgb4bGNr8QyvosJsxyrBc
dpd7J3zzW9+mCBXBe/3eef9OYBUiPyQDwxQ5QfjD1N2Z0+0HHFO3D6ZDmg2+yAD/
sqSSaugu49I6JS4RD1CVwMWU2VgIL+bZjZ9QoHkJwdl/iEmGiZkDdICRrXPOIYCC
71HthYnL1AGIpy2pyy6XzwRgXfxrodUAYmYqq+2IFe622sJMindHyCnYJ8ezqkyf
S0oM+yWiAiLNmoSWxlBNIjzjR3nko4DgQfgNB+3giKGaLVnryUdgikenn1RSaJui
vbsDMRYGoQjIE91U+hvcT77JKE6B5WSzq0/mNJabQyth/xA0+2Wrl7UNvso1GOkl
E+PWZxZiFtsfwIPDXgLjY4WOISNArY81HXdRZZMfVGFi3iFFYUIYpMAPFlYMdL/E
p/fWSWms7DgdQhP2c+qg3anQfGas/n7gEGzxKafdeglAfz/01y8X8wnj9GgtvGCU
WVULRXAbpWVy2a9IzLplBfW0Re/GSXR2zhWSA41Bn8gdtztdLs8HEwkfTnUfK1gs
B6M8GakOeuszc1sYU4mMsaYoBeiAzMSHqv1I6GhJorlHhU6bzWlRoe3xAgS+ubuK
AIBOey6SdxAjHhjLWPNcPwfn470LsF7w7kO2wRsrXLF457VipB5bZ62McNPiJMhu
fZiipe3kgBdRiqiaA9lhJmSeu1T1iuBBjieWrDf+mbJAX4SPKTTUrSQ2zx/j4NG9
lOiIrhNYgNg6B91Pe7XwYR9fi10jW5hJU8YKWCxcbvfUri/U8UWhWKVKCe5HDzqk
cEuF7yplDI3mEX5pEZFts7vsozBaBmy7vdIvZ3NhbBl0jMkRaoDsjKsjA7dGIvG+
Wt+fnVZiW7RNgmZ/LHFi4q0IZG+hKO8bj4wgzrEUO7o8GFqfGJU3OmBaVyWVM8rd
+zS6jN3LiSBp5kVdDhoMWS+6fbf3yXG5O0APxAGaiZiiLA7OGSBMJ8v+Dp/DZ0tH
Ne1PBBF6flawkA4k3S2gCvSSLusxmTzMj8VKtnspTgPr2WRR8smcy5Ozdd1qX1nF
N+HQBRZOaPBJT8bl1dv/9/JHiRM0QmfpqhL1U0GK9zCDCESqQjXSRd/8/hKt6ZAt
nVurbMn92kdaZNNHIUdCbCHmbNyLgPNNEk3okMt311TWbYHTuW2zEF5lO8JmyBxt
DAutvML4NGpP0fUCsUZv+VtrcQkYRf0aCr2xnnq3+xBcPDKSLpiCyZJjyNq1D5kl
2dvU52P/OWxwQWmHpvTddLjTKLPLJkmszCQrJC5QcZIHJ+Kp1diHtLtjUHIyPZJp
G6wjd2F0lhVmIyKafeLmAa4slUqQU9PiCbCKeA9R86k8Hc11WltPCAr0h5vaxQ/p
tQsCHHzOWTs1DYx/Th6EGjZs//t3QX/ircHVmqnF+rSCCbOXnSFwNhZYKaBLtyW2
0lXfr+SUYHz6+5RJW1OyHQGYVYE+qKzRgcInMaVr3302N/moIfLkX3+oqumlnYIA
38l5IFOYRMOnRwAngPzJXEHeVEqgGarpeeX3jLg58Wwwk0dTAWO+JhsLQCW0r9L7
t5YZh8/AO43bGWSTFz7v4EY5pnEuxL+cicd2FZMtF+Vp+c4LXZaKPTATFBukS0OH
45Vs1iMDfUp9GornCyNvCoUpkwpxrq0Q7ewW9jMr8CwtunAgs2WLOaWSxMBVO4n3
W6qAOn8yd/iNjB4pFmEDS1037LhZtm2JQiHVojn+CYbJv5nQ958uAOuuPXr6HSTN
romhHf1CVS1no/jFPYsJ5p9ZPSk4vUW+LoSl1tTJv66YCO4SjlIdWOaVHDh6F78H
CPDFvlTqcR3DSMkfwXVftEsc8QFZCu5Y3eCquEnAoCY0LeOlAjhpt3SJLuGx6q3p
WfbMXk0dbqY9aNXpbwN2BMjBSKbifKhQiBqjGz4SHz2LHdSJ3WSzE1394Sgp3RJP
QqkmGxoS2XtxyZgrNywHyTKN//zmj0sTbfQ3cdAI+IQEh9X/mBhgbBAoox2k4B+k
7ev/f0ryi2oitV5whJ6g60zJEE8FmKtzifyzsy48dBIu5wmwBb+uy6s2p8sfGSaN
dNksunUwexc56p/qOyO3/wYw2TpLh+Zq9Mx3AT/NGQIshgnM2RA6DmjNOX/7MLoF
WAESiNOZo+wox8J4MxTD7k9qzjhP/wPDznVKbj0+4fVXGip0enNnDm1XBpmIPQZ4
Kx6NZWVW6H1XQ5Y6J68AWRTzaPozbpoTuU4xJM1YlWo9uZl/yIkIB524Wb2lBp44
muRMfNiGFpwToL7tCTmqGwoUKatUmH3WtoM84lc4YZbwNUAQh4afQxFdii/JpH1L
zD0qhHkOihNXHHdhle8jHaowF5f3/qI1qqc4mVGbj2+zuJHEeqfky4dzTpiorguz
ibvMAtiJmh0KZWOUgbFnwuV4IhRx9LGSnq3GnJtuK/PkYJiWC0EV6/kNUVYHp5NK
8sExfEgzJkjyfKfweq80E0yeuzashGyrGHyA5psgGa6Qgp9xcXWLKuQ+nnNVMrcZ
hY8gSnm9aBeuJRR/xjn6DhKNM7ITy+uOt255MLQyZHwpXPzM/DWZOGeQkx70dd5j
6GQoYLc0lzrTnfAMvrZru5uR/XzxovJVIAfzkhRhyw3TiQ657hbHtKv8B86l3Lm3
5u5becdD3SeMx/HhymKCKI7l8qtrggt66Fo4WI6p+gF74j+wTyeaJvs+gUUGnkPY
8dLQW/njrzw58eVrvOlkq/WnA8cBGg7We/esvjnnB2w3F259u39kWydmgCe9RuEW
/faK50TXy2bhNl5DYC5zOGsyM4u2WAHStKovx1wfLSzHdk5gfm1QsC//5oX+tQzh
jNfqfLNhrlWjU95HGv6JZwgoRZouxrD/afR11o+5eAz0Z3UIwdfNQw84BfMMw4ep
h3q+JY18m2rhvnDzIr4qnnSvkebPFKDckPYHP+PVnh1iAzsusxeLsjp1Qez02B8D
6Wed/i2SudRwbq4YZpto7gYbMoOuHuljnl1udfm1jWl8yyBGyxdqOUjzTn3yav65
iYXn3ySALMQyp70FYOnrIV04dRFLrc9hFkIUqp7FRVHGk8qGmwnKg0HUSVNjBFRN
OfasCCQ4ggRXm+p3teWsAsRzqT2QQxqxnzClP+N2/Lqmkv1Fq/kPyErw6q0BrVZm
cnkZm4kPsyg07vNle7kZRJOI3cjuA3lMEzp9X6op+xi8Yp3XPf9nEMQmsEYaxZKU
sHxaT4b4h/267pG/G57VlUex8xMhzcxT+1/hGbVSZWPAXca5tLXk65EF0iSsA0ix
pv1JkbionNfFaeIjN6pGEmHFjN0OlPNt57ljzcqDWUI+p1g3OTBiChP/R3FBDGYA
1JAq6tZLRZV7tM1mhvEf0cZ6RXfNM24CICqMcfOnE7QR2DYqwzq+E2t18J2PepxP
Ppzi5m4UH5za/uS1c3yqNrbWANZqPpECevj10ET+eQidRR//F0BZ/DpNaCCr3WVH
NAmayBytun1RHixSqITbMY4946ddNFWOqlyZe3JkpQJpdoPxI3GT3W4ldqvX7YsX
8VqoQSrjQGEMh5oeKYK+AqDFgGyoMGRmQQuAfHvZ3pIflSdqUFkk5c2TvnED+0PJ
hJf0BR65B6cZVPWz0I1hJu1s3Z4N+hpI0tUIHa8g2wU97NlRxbZ0DldpoDoTQTaR
uT1cwFikjQBD8vKsCOpW1AbTk9b19rDzbvOF211h39qFDIpBnGU3hkcPZMSX9ufY
PPxm3Row3TB3wpjZDLolCXoi2hgPnEbzCmiBmIffebMFhkpcdLg5xa/HVDiLNwIK
T1OPgE0sxxGaMW9m9NNsgMG34X9eOPWi6etQgNobxajbWRAoTGZ8fxGT85ayebrm
oRVj+YbqGXDY7gBv8uFV8TmrOVnIvT7btSkqYwMJ/vugFJRPORc8Jwf2zQbJ6Y3s
GFPiMrNWmv1fz9V6PFlt2sxBeRcvkjcpYS0pmlbavGLSdkICvYi2dnKamMt71Gx5
03KwEbC5OdK8cd7AZlwAIfytnTSs0KyH4crEqqOO8Nkepzj84o6hCdcy/6RhTKYt
oynNJLwm1+zxBn14FYQoNW0fwfBx81nDGN3Ackb2lAxcMUVOeo+Anzsj+lhUM7fh
NujCos914NK6X127rRZL09wuhdKGH9SIE2/Mng9lv3bENEmp3boulU+4cp1nCJQc
uibVld4WqVcBmosAobGSBJEqQJ3lBcGMsK6Ej0xqCpVLuEucUGsdCExPGfs9JbdG
TAM3AuLQnppRSQC201YpKuMoF/6hW25I10fB/R30uv6O3+Mcwefe5nqmuHjRp41W
Gwzy2lFaMregHab9DEh/ci7gysbrAjLAoNO9Cq3YdR13aLZ8EWNdEMc/uZGCrtKy
X+Lt19ypHy8b2XecBQyEc1WKwhTsWJeMbmODBUwln1B5RGH/52D9D3ZOYIsc1/f1
8PufP5Lytg4wSoFlYIDGttKAG8dBm3G3SRNn7obQshuIY2WbSZTS+UwsPlnKN/Br
Nec3VQW9VZ1NsyTq/FGzKSQbuQe0F77uiVblOzMq2kj8/hb79EBc9DW23RIIBu1S
qm92KOLyuBj/qpGfLckT2XdiEpaeYQ/Hf//oPuEzUStMp9VEWZ7S6ooymKrGIOA9
qox9QSQO3HitXkN4YIZhvHP5fbWev7h2fcYpr1tL8GYAjgdQvsL5XsbQpPZkonm4
jD3c5b7GXlR3jl42EvSi+86gegDADh39pK1eQi6CKQEY+dBfQGB4wI1V+pPinmP9
sTAMj1ApKdfyB1b5iOjs3wYsFEWhVDKvILoEcgKFkYOGeO0x8S5GMFWJLVzLtZYg
1ZQrS0hn/AJdkTG1jp//qQ502ehaS6vQX5JBE6QTTENST/2WffGGKyCdQg+ebWQ4
2ERBdEzbbbgves3V0h2MznNWhVOrrGgU63EMyGx8jKzOdCF+y6GY57/vgp1sitKA
NJchsxx+s6dGSp4RVH50MWkjCYAERT4B9mtN8vA20cyiZJGugoD1SVwtoUvPfl09
KFz/K0gf3S1n3sx5NP72MpmWCG2s4cBCyknMv+04Jx+3zT8dHKEr3fZb5zRkq1lX
ED1WS1Pesi31YvPNuveV/3DydF4lNxzGgFB3vhKCWlcgjVHRI1NBFOrsVWDTH7lz
R10jWKP9p4+9Hewh+JeH8aYoExSOoY0clztItNmldYCklkOVEtq9ISpKBL0HkkqI
FP625O4py81MtSHOYqKPNkgPXrSxH2B1vRuY7NulZAMQBAbSD3jzZwz45CYZzHWc
VTcBWTRmO0vMUNb/M64mXsS2ggLMxtYvv+J2vly4QUMmVg7CijK2BEo0pauTBLgq
NwL7c1HpjVW0WT7yPe+14M8XW4Vonvwl6m6ZNZBAgWs9vMbR0+/2rsl6twxPWSDJ
+bzAK0AgV+majBt027Cs538XL5LY1msW5Pv8mqd9NfVkLWT9SPKo/vUmCtNS5KeA
OtStG8VawRplFXu7dLbf4ZI+g0OlaT6HXalHkUI+EiFnuLgmBUYhdhIAS0cy4Ayr
nSLB03D4P8DsFl6OiMwlE72hL0lFNfM5OxGMxHIgz3TxdUujMjXdMsGgB7NjKzYR
Q2Hi4FuYdX+6lTe4mRWMPwoXDR/+jAKZDPYDxS/A6DwktwAU4wR71+9wKroG6J5p
BfXDNNaeItPkx0/fVTPUfMERnRaQSDWYam3ktKeSdWdsMbUuK1WWLBDKUq9yw8Ap
svH7phQFGR57sdRlGNPMo/yz7l4X6UM1fOUwM0xB2a+GePGecgq49luv/wZESnLG
EgQoAQK974eatt9PRE+CvliBlbP0UtRylhBadk7eIRo4nhkjS13UuGnivpAjkIcs
yQIjktNY7fgzGvi3wDuJGlggo3HyYsQRBDu4BPzrYjELsBTj0fIjqKCjeBlvLO1T
8bI0cCLkxsUTuVhsJ7xG1feqJ8nUci6ujcCJwHF9lXeXmwKr3PP6gvnk3HblCEsY
aht1llEJc2A1M9EJt3BVU2JCldb7QMgiuTsbxH7Mup+EJfX/CZdSua8XD0ZnyLal
VbjU14O86JEa9Qpj6HLqay/1vRKpGWfVjurAm+1QhmELCBFm2J5yDuoOynXKLpia
z+iAeEjEi2aTPIYM9BXwECz0jcVIem4J3o6kKARsSlqe0lU4dGOlj8a7/3dnHP3y
Mhtnmfbz5hHb80O9goEZpS2iHdiWQqUeeYl92YMc+HCbtKuI2P8tK8poA7HGxVif
xCgTqH5C5LWs0HlUHI9sdCC/d65ZgWZmNCYugxnHjCirXoFEvAI6Dvljl6KsZjus
tAvTJKv2uPvSVTknqRk6hy897cSYVEZLxI/oBmoEYGfYHIcIW7ghSGnHOhmztRhm
HLei6T0ztiRqP7n/jpbe1eIB2jHHtRy/wMun4Zg4DGtkYo0JHYkjKRfu2tE0ey5j
tcVfsbaLxIeI2sn8wogXTcnSJMbQy4EedC4+XVSR2qx1PGBBvZnNnx0sIhDx55qj
GaD0GjfuPXmKUfVmNvJQF8xtdzQma3ZYfy9IIAX99FgKKhTL/lROfa3SWGJywt6q
soM8yaJ31Ztlo+qQVUxLHcXnc8Rjsvrg52y9dUNsjloc7I7133vLm1xokVyX4zna
BsVvoYkElYjhjkhgvOtn0MzYR464o7t0p7AE1LATogv4lY519349ot3h0DZCpTcB
nYXRJhPhP+CHLgwFcXQ6X3oKpabRSlkdrtQFSQQFce39vqbQ/XoZTQzzrexsfxxW
t1btDtPStM7Dhh+fYNkmmFOQyPZfW8z8oBSWulpdvoBd2/PoA3MFa2xcnXTy3VhG
XQ5eDRjsNe+E7k+WkHMUnLBjKhPlt6wjJfnpfr7QZCMP0sGYhqMvlZkTynmO+SI6
o9TTM8DaTA9daOUpPmMzgdbVlHWeA2D+b0GK+RBLKXajpSevDKxtX9sOCcxmGmc3
VhTiiPQxnVgO0WGnt/mwKvUS6rqvB5+BY/tAU7Rvec/9sdsQ+PPls+QKsvvpaqv5
/L4FbBtGEVOG93VkciFuRumbasr0axZpoShdROAONPIDQTOR1VAEYRALRT8hyilv
pQ49ZA9sPJpgmFISS/jkOhRZW2xrEW9kK6XuYJS5FkwjBVs+PDN9jDDV8tc99zRf
kds3Mcufzhl+0V+DKmf16mCflR5s0JMAT7xBi17ZprflFW5ONOCVDfEHUR3H/U1H
KNQCxQYSpdoXO8U+lC2RvxNBBEdV+gECPZ4+Oa3oXbIQDWDATFDkZwkTshYLzEQo
XIvfTt6wmFoXQ1ye1PQiVhx8R/wNhaGEl7D/DuwKG2/y4X/4LBufWJbbhfPx2Odq
XrI5pYCHKBTBb7V9M8LE9jokj0D7URC+mcXcHKswmBwuonRuuI+ULrM9zuSG/N5e
1ZS2gJ3GQEiYoXAw42XcVg19MPhxIAVuH5TISYTd47OFv2Ef4jpcYk2e+tU0eUrq
GIOxUcuRGKoySmGHe1eE/sat/hs4VFc1opzqqCf3+xZFklpJv26Skv3mwg4i6Sk9
IW6qsddiNE2aINIKJ7LuYO5mlaXcEJpEJnawI6voUXNyYopzbvN7ftgD5jsrLClf
wxzgkEZrSwnRLK19Lb5KyI06+krkAwtHH7f8gNO5UvWp9/zHqwrjvnse347cj7wh
s4uYjFw6SmBs9KdX61hdbeXY0fuMVIspGurKojG5vcJ4ySazvxwSVO1aax8LnbVW
EwmxXvIjd+XQfYLgVv0ys6GEOv+bNiC9+0ZBN0k6O7vO8FEz0Us5rcWmzd7yhliV
Cx87HJVOytWZN0kw9IIUs7uxoFS70JT8XkfQA48Fwo6lO+zcm6xyeU6h0bCVnKiu
BNzTERsMYiU7vR4eD9qu8pmfQl6eDoQZWh4GX/10WYFMTgzQ4WOcd/1pR55IBL9r
/tZU5vdUraw8pgvUJ82J73unVKrJ/WJctvb5jX8xt0W3oUju03birqEjVupIoRKg
7sLpwQvZBSVXPhs8wWLcbOGsYCCeNQfrhrUp4TghY8MXkZGpTl0+45g3Y7qT1MPO
xyT7XlR+BnNstpnZ/wrxMK67jb3iXXK5p5D/HUw/BoFbu5BzqL5JriNxOw1oCcfU
yXShIsOAzQlWbjb54j65sq2BiPpw1DW4+USiKHgXTZUhZwTxxu83dxV7Xj2uMbZJ
lOeTuvbYDsIFiJPKTFs2l8ooB8FQMNriel78IFWtsKGaoltWSEvSt4+Ot75qd/o5
rz6DTba8q7Txh8POzVfT1DpRcDulxjBo9PVVgpgOHmXK5zcfmQYFu8LJkEL8J8MG
fYz4HZwZQXNvZs2KHsU0LErYKVOjcPfE6pX0CT3b8Gj90XToAa4fIyDFaQU1hE3h
F1brrXdhuo2iI6DHdeRzjMzTXKfoVZi39kRBpETsf5frCRtDWNolqTuFviOPEZhy
Jc0kExs9aCXGVJzrxCh4lAWJunBg7lLuiOQKjURqUvGV+LKPbIOTPoyHEKHswaPe
n/5bS6qMqA6ZjwOgS+LuQY1AGeY9bLX9Y2JFwE0H7syWYq9pSFmS1GSem1eqGANu
SXAEnHuuibrvO+3SYHoh/rSAFqUmMwq84qrv39TItMykgrKi6f0hvQ7jZGMi37Fg
XN36ciPPDnqZNvPBwSFQkSGK0RxoHUWiKuC/eteTNXrfG9WUg//GGJBivuN5AkdY
ShU/vr2M4fwNX9iyb15TZIWg4eevczaC/K6cNG4UkgU8Cxx++DWwj7t6koj/fV/x
vuxfny28lj6MLD3p5/94ggX8snfmMiYU9a4paYARkz8kzOXTdNYHWEeenWZZDnNG
J8c2Q4ndiBGSGVOoY8rzZFSNN0u6DuVY3I16Yd+4CJdl0jmjfhtcHYrQ4UiXfqxM
15ww/ObfPvD306WAXPyGXnVwX2lCzWB18IMDCmpShkEzyvUu1T/+1ZUbMCqmgG3m
U8V+IgaymHWwb1aXZ2/wcwyZ60CCDF7VptbGh3ICL8HvbB1R63mwGrQ+IYyAvbNE
pZPwLXsCqx6ZsxvGEKdGnMqcs7RoeAstpAVvSBNXpLxw4BVJe19sK6SLdtcPdxG7
x70yGgWskUh8WkL+0h7hAnd5zxDnMoqy5c2Nuth8L4OxgNCPlg6vEqmB04nLOzjI
kp7pimKDOxb8q2OIEjQNiKSacFO2GSR9OfH76ZRiGA1l34OVMewUiVpttMcHchZ5
X9YWMDww7dzi3TGf/AmTU/h6d5SA47hrD5wTCgRIHhu8YltKx5niNvuP96tgqDu6
aQH320uY40bsYYTUzY+LQaE+B03ThprzrPuzwXPbhma5Y0uEAZ1k4EjlEbkYmAVx
rad7eK7L9i2C9dAiRHb0hY8u4ikyh4vn7G2/4tFlqiLPYMG7mfcID++/BGdI8Gqb
MJLQWy9Rk+mlB/aVbJNsCVoRh25L7QgGr6seaA467UTE5Q/7/krhMxSIIxI9SUJW
g9oFso+a6M7meTJ8ZA/ynIClxy6zLf5QKquYe0V0/qSS4TXZthxAkAzgVKhfjrHB
XDylegD2Bo14Jw3SdUJNdjGICLAfJLPHPmBU2IBApAAjyNSbGJll1UPvc5F3HzGR
qdQDmIYEgr+32A9XLZE0iRZhSoPfYZUxOybB1jZNl1SDgn2ebJx6u+EPAi3NhGTc
aJBB5GKVs6Eqyf3nMy8UMvj/XfhEFoTfoDtSGVl+j687Lq1vjTXx/EACzUsWIDpf
Y5rybu95BKHkqBJyzpj+bmsmQUxQ03v7Uw8BH555LE1g9EM1X8NPin12YnEc+xzW
FSIhcK/XmOcjXh3poC0PBQpoauAvuomx6E++C8gF2Lig7mAiHnDcmInkAuUoqyr+
vFGr2IwhW8ns0egMGQTByoPVMkF9AY//6qabH2jxxaG9r9c9ghD0LIb+vcEInuj3
LDC3kwsQ8Lds4l0kyhM6qym4fpUaz3joGLPTCdhwseC1DCngmS2EuoLjY2q46o0V
KrVN3JUbt/anARrwUdnmXWVTz2AJmfdrIrdf/vtnPQZ//egOEoVxr0yK4Yeq6ov4
ZjYRtSVg3/XT8IFnvz79ilkKhuIRGCPQg7r74RlGZz9ubHY0lxpSd5fq0/dIZARz
C9/Vyyf9fHjF9VRUtpRAfGQGtkQfS5WQQO2ccHIFdJ19llv0nI/4LjdfG8/ZtHYu
9Kup8lGMPatfeTJYWxeJvAiUc+nYbXAgwlGKXOl5PS1w0WL20IBB//nwJCLaInaY
bWO64lM2k/CxDCb1c6e/ynav73SHECWLOxR+hcpAdI5r/oL7z+gyADc03hta8W3h
ZlhRvpxsTPUCJWA8COGJpiXTYc57eusIjpArNG8b4TJ4pE0LZiP85qqhexrENTOM
GCXNtJErtHc4864EkFdEE5kAsMzM5uSStNTtKCA83BAw9RbvekwGvxaoZvr7Mz2c
VwHFh8SkrKaKSbXow2n2TelKx05IGbnxPAqd10/9or1Px1ibQXKPGA08fh1JlylH
RfQ32egXxclItu+Rcj/yhIyGSGWkM6wCjEzFj/Eb0Br6FWukhTzmsm9FjGpt2Ab3
NkBhIBn1NSxaKnlm2n06fQ3S7Ho6zMonbKdXeOsXtV8t+iFFnc/xmq8LaYkQQncs
YXCwWSYbdjqqsB8hnb3I6w0upIHRRDXoFWJIlT0DfnC8VUpn1i/whrQes60Nn8ud
KumW72jNkQ+CsuhIXHVJiURyqVo8nkEXZ+QbAVz+DQWEzKlcQJmK1LR6heYbQqJP
W1kaE6fd+poyX+YQmVkil3bAhRXpBkJ7kkf67Bm7hhi2UCpu+ngGq3r7CDSh8F/k
1VTRd/wLYPYG2Y8cLoCCtfZQJ6yHQtU32lK4oDE19p5sBP/ZIId2vuvwA02LwUN4
fijK1TME2/LH26KiP6LTB8RO4uWIaJ65FkCyRWETlSRl8wk+R6qKqZqMgifUsbyP
Q0Pia3+G+kruglZQFQ5Eop79fhSfj51Qr9Zz1g9yCv2H9ZW53/cSVagHylFDOqYe
NgmtgCDoqZO4VZnhszqag1NLwwZc0bo3L37l2wpfds9tRCOcOWRI6teF/oIE676Y
kySjL1q5rfRiJ8leorpJo62dL/c585FCndo46WDEd1cP/JHniJ0pH9wvDqHcq+pY
5DfamgU8rL5/COmZVeaMBjzTo048lWoiTeUoxt2y/DCpO++ScPqKLI/R9/3mdnTD
O0hBIt40MHkbB93F4kw7f38CP6aA1b7MLgHF45d7L9g+iA9dib2UxQn6vpS3UB9m
H1Tjfn8ceshwZmcGDc1lnLZZtFcskzki8tdUKCByObY/I0XWf5b0S/PTDVDovIpX
gRX/XFm4lGcYK03AfchoP1i8CCWYefDPwb0gzSBCUPwfEJOKY9eIAUDu7XVbxbGY
DwQe9Wmc4QVJa1SORfwK0I7Wjv8AF/UofV2TBl0B27IDoUztO4EfM9kPRYXKzPS9
jM/TKjdhCx3y1lO3CrWx0oNhKxtYkOXJiE4x104vz9zomoswBPoQs4voXqi49YdR
76MRoXEN0LJ9K3ea3gZkPxUjCWNN1JJDtRWr5yx+1lMLwNgJxK0sCJJqDwsEq1+z
CaO6UGSWNpa7M3wlLmH6wpyL+O3s+e3Nob/Qn9cRtMxu6sDz8xOTdukVxmla/udZ
bGrmVaEtcTkjqqSCvgEq5S3Ru+bBI3JA+YsFYiFaxYrLfi8zYERkoNb079ZpO/VN
4a7+zmTgHQKo81wFayC1Sz77NJLxvssDAiJRz1Ju8SAb2ODINl8hG9uR/ivtbW4i
MocnGMjdL3AeUUNQENkjJmej/XwZGjgXSIOj0idEk2nB6xJlJNVzp9a7z6uST11B
wyXb74ivzuQVK++mIcqqGD+bdS+AsVUWfrws7HeimwQwg96u0aidC6EVTvIuD0Fn
h+exeoXF9iVMHfilS8JJuq2rO9Fj5e5HnID7iQOS4CyIW7jLDY54r0qivmkYt+9Q
1yD5JEkoTfogQ3MPpyH4E1Xo5TfNUQCEtGn1Xo0eNA5l8gVRjxuE969AH9van4AZ
tQuvUn3813epXHCRoTsceuEt5KVbsaboRdEla7p5gXFVbdY43VWtMSfE2X3oT5LX
ErL9H02oTe9CbS7FKT0W/Xxf2tA5Ig8c6OTlw6RhkHlrCueP++FXpVcjPujV5aDF
tD2p6Jf3rZcBarAAJXYpaE+eIrFArkBfVkqyTIfdNtHYz7srG1ehX/2hSlelMOWR
sKzfPzEuLd6yuPKi2+SsGbeDP9nURsDNMbgHW1jovyt20apVNE3ton9pEADPoPT6
DqTllZunJK+O2YXKfDDSwbQz1GFWVqJSAgC4P/PQpMDCJvzcNE6dXJJJE+B15Qkp
7KtmK1jBksejBCWEGdpnT9yfwlNCsxMdxd5HxLzVoOO0SineD/iPm+AHYg01+/8o
oRoJEuDnkRx9X0T8M1iQ1QkeIlu1IwNjsIowxUGK+o15gsrkwa0/Fjzww2Y8frTu
usU3F1PwE5ZGO77l02piO4wynzosDNJCeOe1mKbz1qqOS2w3NMYpLjkf7vx6gjM0
f67ZjQ/88ZcNvkbLNu1Itqxq+EfOAdrR0j4fXDbwLJYzMr9V2hOYFSXRDCEkskiz
eSLtvYRLtgo3eSlBy0GYqano4pzRbkx5NXQTHoqZFtkCZ0P+Yj87Zxm+Z1aU1YFV
2m9K5RJGjNSORk7chnMuwRVyPSHx9HA8SjLR7/jCGDIx8Ux+Xjp+w1dlac8BXXzP
HrOyzFOUAs+a4bhyHaaHlDXG8dda2VMkfPzCbTDC5vb1GLQsIrUKhHqRKtXXo7le
F48Q8vcCcUJp12y+MjQAAifwNDfWKAtKJEdVJWVYRQBe2padfjPrtokmvYe9chnK
3QebIQI7F0dvTwGnzYQIA9fdcJgTAnJ1wrEkTEvm70KjYjqPfaYNwk+6DVKQpMEq
hHKoy78tjNmFE+OvHH+7yjyjjhtaW62iYbrPIrnRZIFNIIu7IgNawgsY6t0S9t5v
nA997oFjqyihmSXKwzfbtW78HnIglmV2+wHPGLDjky5/RByH18+6mePK6VRIVQDJ
njIIwZVrFrpYROh8IwJ7ZDXENeO66Z45GXwUKmr2IPmPKOR8oTzDN+4n34ETOmit
TtegF8V7Y4KP40+4lw+/qgFRHofuuNn3/7Q2pxyotCVpB13G8x0ZyCn8e8c1L/cm
gY5BLNOaoLxqaZb6q5kZsG4Eo2DGAy7VxfcEmpa0+e5X18ZeVjwlPQQk+McJBbmJ
zXDv4U6NqVJtZggf0RmT1AYdD41CuHkcJo3NjScEwvhh3r3c9SRz/puVZAUXs0n9
kImwlWWwnPpWOqLJZIS37Y8yYeB9A3+bSFhruALtHy3o1Im2WorK5lpDZM1eFqTQ
c5WhpLAj7/VH3R3xu9Uaf6dzHp4R8P8I5ShR/vQBoOeTNWsf/Rc6TEifcDHwBeE/
WpIj2nvVEOpcFI03cGyBnR1GXOHdcd62jwOKD4+JJrYfwagl/UErOMNYMOMjLIzj
2e8wSBpRoknicnMJdojUj+q3H55dX/kz1tn+pkLW5UFOooM/QPIalPlOnortOBjy
IxFVmZ3rNSfiWLEsE/PYwYRW88iqtv+ToXD4GewkAmKHBJ2zCknIODs6qF8UqNPC
CxL9pFwzCEA4HxGwOwPt2H2zfWVDQVWuQJKb3y8AWJJsXNrfWBycOy0ylXNKf6Vd
S7FKVsFxE6bCEaVjsQ18O7tXOirTnWxZAMzLeE7fxgv3ZBYM5WBOWGTidWFhVgRS
LaPZ6et+QlO9HUNVdU/ko3PTwbuKb5316w8OscqvoDCuy6WJeljjAyXx2hOiUI/H
29YIGQQ3sF3/VcntQHlgLQZvjAtlYij2iqXLwwlYWHzX9FXiNG9n5HNuWywD0Axo
6itnZpnuDel1IjCW4XANtNhIQ97ePQ9I/3L7yMzRbuVO3zvRGsFfeLA3OqKAp8zt
xpR9NAhT77aHEDAkT1nvfxm8tlkqFlcJUbAsQ9EnxT97zmv2tW96FH7tlbDbwrdA
3EqRN88mMUR02u+ivc2N8p9hz4rauFcrQyDeY+4mZt3ACjpJgtTuENNojCpnXC0O
nhetaDUlVC6Hf9H5/MblGEuyodUZe9xhk8jU9HlFJubY7l+6yA2YjxZpc2mKLW8B
HiQnGG8x/MLU08qcoCFhmDZvjcgUJHxt6Xuw51M35NaddKl4e/DNi1NQ7GoGU/p3
FX3q4ClwEVEMJ99xbFNeuLnOsCrj1bzW5T+1h10nBvsJmpLpzbF6U7Roi8ydFqBc
Frv8WgHz79DaXBX9+WrblG35Pn7Q3IcbNMseRRk/CjEdopEIriW2n61wuromrXrN
baJYQrVGcqTRfIgih3APuRm2eRRUGXrHWvDzU7NW8Iqt3E+o/OT4iSEg+DCWOH00
XIjFJKTrcR4intPfEdTUnxqjmTefGUOpAK+XWoEzyZldEtx63WihCsySXWblnRlK
eBA1yG+IiMPtH4ApevfpjtkY+S8wDdRVA6k0YLHSuqBYZRm2femi7G52tIIA+gpj
3eFEIY8xt1815XueO9iwc7Mhf3I9oqSmwAKphjKDSQlN/e0ZBnp44a6PokHpcysR
+JGpEp0jYFz9VIOlg25x9eZtU77dUDL97fhPzG0NW4kYVVc8lFAmOE7U5/nOKVY/
nBuny5HmIRdH7s/LJnnTVbl9AJUuOJRb767b7KefVz4ezQ1P53Yf7/CoOH9T+U6o
yD5pLL0jKvoYKhOtT0kGTPtSamYvZQbOG3xdL+SM9SOMUmbReImXNZx8fEivClxi
mZ+VW6YwrmQXllVTEZa14KLlJ8Mw4ocf/PBAf5nmpwdtstJSzLt88gSNLOq4Uvx1
0YsVKGIgSqkTXMLxid+hNEVGYEPKN17avkbyMeCMXRsAasqrFUGeL1zo2iEj0aQg
8Pz6R+cr52PHI23Yfl60H8lM94XgtZ4pZnpckohlXDFfcWUkZrO5xsLawztN7SA2
gnnJv45tvd7pJlT/L/a7ZChNvyYRSXOsUtoFNQofeSkNAvxSZWPZSYrnZL8Io/zD
UU/HOOCm0qFzpld5yjSBFuo5u1rG8r/YDsR+ZB2ECoILmfvVyIopDYHR9DHk2Rm2
jh1DN6GkW+TCeWTh7WC4jxbfVZqMU1w2+jy8crkz5Bsk+0pq7OzXvJMd3Bk3VDSR
OHw5IG3zfO9/JpfFrFGbiidesweiwF/kN6nSHLuqNEQixKqXyWrrJemXZzBxKNrY
EuNlSGenx4L90b8BfcIrQZhaYHreQtUdEKxLczcs5cV8D9M+os8+M0NKAXjZy8h9
/rkS/bwrIHpjvBvWgb+WahAa6SIrcBESjHEB7/2te+W4GE892Jf96VJ770FWS2VF
dgiDMt3O6Ge/gcCts3eWUyaPoH4jThELw8J0i3u2nzMwMZ52N1fWTUeHgAZpEFZL
CWvUR72OOZH1x00+jD2F1XCqDw5iiLyznoClTUL+jR0ukr+WbVwun/vqOHMJ0meK
5lbtGvsEsMMT9xv16fKI6FbXsPbDd3dL5INVpYjHwE4xvfW1pUyXmQYUdhsRN3tx
pVUoemaqTkHRDAJCcGBXU7dHytlQelptMSfVoBZrZMQFqjM2TiWcpYLvi6dTg3Hf
0l7Z83zrpq2ZJENJWQAvUX2wTAjXGkw0mqgHsxZ5uao3SP2hVgX68XgGhBHbD3g6
UOKheAiyRxgYcolxQ5f5wWarOsPQhuRk/perE4ZqFtzaXmcKk+pzuS1RKN+/yXk6
X5mMufyRmRYg3w1XJHscqmyLyDXiHXnj2CdBsfSRgysIR6AMEBi79HJINz+aVEBu
hPzfqDXm+A/RsJkDuYGBtm9r2IxYDIDj8ujh8cHKY+HdbTwGvlYtY3lDuY0u8TaT
nRda5Hw9jI880ZJjJgsgWhWGYTf2iwuxqPVeAGdGYLboZKWzYvnqDWno2iIPNort
gTZgA8wnLuYxh5HtTvBcIhIWzi+52tdugPRKt/RsmC3iT5G0ZN/ISF0rCl8yrN7B
TFFWF06ppCXNqqOD1NpPZxeWtfxMsrvO49sM1Leiddj1YfCJyu8fo3im+mjbvdK/
/33X1ZgHaP+7POll87W10h4HNf/CbFx+Jq+QDso3fwCSCi6fCmq+r2EH7XtaWDNh
sJFSkS7xp4q/FtY+ntNCDEtrIUypX9KZdAIr9FsgkGCupCXDZTAwje2JZvZTaf5t
rhZKEdJ1xDfF6zyoL2saUiZCizeSaPfLgLGdjumC67q7nKMCRnACyR84AFRAB4kw
rEJPxdV42fSUsLtXt5nhOm/vyxPB3l0Cx2prmORV/3qkjt7G95AKiIz5w6yOO+qL
vRtmzpwO/xpu3nnydjAptiVqKzo3Oj/liQNjF1GPljrC7EwfPY4Y8VHyCaR45DO7
zQjrWw4CeE0IkX9uHQ3NlYiGPl/8CzCHa0mc88eTOSQ7zxTYUtJdksXBF/X9syAU
KMCR/cw9hymqBqbp/j5ERvtbErKs7ltS284iY9MtQh5A5bjh3yinVtifIHLd07Dk
bMl7lz4bUQcnUA0T1MV7L/tM5+fY/7ZVOaKZ1mkhp8OfcIJ7EBIHgWVVluUWbAtG
FVF5sisyosDFCwKWKQyziJDQYgRazJbFYKS5UEnQiZRy0U9o/5DFpftonvR7PdTw
wj3fz46S9xnwwQNPtvxAvR5SDwDMKcsMDGxgAFi+0ILf/NM/8LZpn16VGozM+2l1
bknMJmpcriOikkTYF0zRkMYWZu+x5s1uadNSpH7yZENpOMYawYt9OBs6r5TaTDx3
gSntehgYFsshzSmZwTz7Rci8nqg2cs5AmqROos74xF6zzJUpsNXiDP34qMufHXsL
4cOBhjQ40AJ+E1XTUP5Q1EbTjLaPdPdpKPtSUQnWfN0a0TO6XwNXdGmwWXb83CGv
AKgmXuupTngnSw8RQoF7XFKn+9e3gf9O5uHsmf0vY4Xg9VSv880rpBIMKYZyFKsb
Vkey1CeXPCBPXWkadahJRmNyE7se9XtnCDaKXhsA8GCXvuqk9TtMF6dWzNtn/NQ6
vogxtIXmdeEJt0jqTxtT36nXUsiti93k8aNHWRPDx0wUbYw/PilNz9WUdHrLisEU
bdr1AX01DBQwDFLvVSvSz5DtdD46oTtPdHelXXlten4iEUQHhtkJg7bh6p3ET7wR
Mxury41flH4OmB1QVFYvQeL69Od4gWdB0jBgMX9ru4+n+Xm5MpXQBeLtUIjGOQ6O
2FLDm7mOQaokndfElU+iKT0/FxCAvQ2A9h7m7qyMaXQqwse7QtqgoVavPJ7u+/AH
b/1jBCvsW+7gVawsbhxITNuT2YziWL/FtfK9Rz/VhUO8k5reV91XW2iVEA/gLbCw
DH1ae9lCGfxs8TvTlqI1PdbXbDm5EArJeaKPXojp9Bq7RXU+HASGbRvMo37HPc4e
OQbdP8Eog3fob5IeZIrV3l2O9Oqg/M0awdEwLwyCF+T7ihhLkKMiFrIiF05hjOrI
N3SmH00z63JhjJR5UXvmmHKvOHvN0CYc9pPeEJ7a7G3idCk2zAoVrWs7s5ZZjzv0
7tzXU6PW9atlWCOLDC7gAF0KyBAAwrYeSYON0eil2iRmi1srIPIye52FQKEQwhHV
nicVFGruefG67iv+m81gfKXsmX64EQz1dJqQkR9b/h6gWOagm3/ZBYUO8F8ktdu0
TfRWxNdyd0XiDxSoLFGtJwgIQmqr7hlmKrhsyHY3tnARvCLdKCbIQmUJT+Pql73z
f1+lsralFufqKdjo0l+Ypr/Pdk0IwNn8hngZ2c6iIwbNqq2MMN7SKhXaUBUc1KeA
EknOGdLXxGP/GJoHeAGsrDIp2/+zc7FI3rxprLIpyoBYyASt6kDzCMjLEg7JDkpy
gYEjvmEOUvYxko0fLKmjKJCfzZp9SEk0hw6CfX4oaGXuryOaB84HjIPbxwhVZJgl
yu978ABzThEznhuzK17QZoO4O2JdpFud9VsGJ2Y58SUQbGl6yRJ/bY18IDjB/cvl
q/VnuMsCX2u52ITZ5spqHsp3TX+I5dOdgJaL6hAal2VcO1RcGJnGMhrdZ21jm81o
4QV4c2+Cf2jGHgmNbHheQiG6odyjSIFvnyRJE9P1b9uhUNuD8y/HZWn/o1ThkUxj
uaO9I+S9rlQkueXbIXmBxp7m7/wKCis8o5fnZGdr9WdN3M/sdnXmQq4t6+nE7aVK
E55jCrdWgMNqVZQ9Pk2oIigxa/GWpOz5ZdcRnMyFA45kBSKCoi32AKaowXlKi2Db
0GvSPrQl9/VOGhMj7K55XSjjDOcVZTfkgnyAH6bpdXmsGUklcLLIVk1gKwv2JpRk
n9v5Gtvge+ZYcp8E9l0UfmLfDNt+Pg3NtzWLWBummQAt4ghVJBiJAVzHvP+7TJDq
LgrD/jAKtucJs+Nu7wUcyeR4KGva8v1bnwL/VcNb281YrBzRuGia6xCgrSSNDvD2
+Bg3uzsmhopqK9mm8QvMH6TFxOp+Vqll4fR3NSuphLuE/Nm2HnT3MTxFq920WXBU
ekpo9JSzRc1EZpEyi0XraCTq7WxgcP2Dp+vjzZBAHLcK8keysqIsEU2YMfcwMtUV
L82l5FcqueQvPLmeo5vEAZHfbva520rH8ncfrjeVyH/RZ4CnWFHgXtOkQ6yCUU1K
NCGJmto4ItFtVbh+7czAV06z1cqcDNZ3PrRCv8iLSGhGOFXK+PFWKJb7RJEMG45q
S4rOMykOAlaXtN4agUQc1Ci+THl8dINnCLKhBabikZzlANpqzX1x+jOVe3ttXRLb
p/hrmFnXHiPPIa53opZDHgvuUSe8dzZg+7N4lqn/5WG3U5Z85gkeAWmcnThqg4lT
lteU6ZpQWoRwkYs57IKfC+BvWZ6LmqASJa3G321c4yzwHt12P6iPEfoGJmKB6U+e
aFcZKy7qo17+KPn8JJz0YKyipJjgWD64pcZaUeAkpV0ki3ZddZ4c3Bnj5lGB9v2y
WT8srS9N1dJWU4PBfRxAHFaZyM30CxWOL6WSoVbz/DXqHzhWb2psBUONhdCYhd9z
BMJxt64cMnjy3Gqh9AmlE397CunFWiEQq/NpEeA1EooFewMzEgP4a4mdk8eqwSqd
d1H4c23Yl4wn5GsKKRMZUdcZW5/EWokZLOm5zd+B3Vl1Thktcmmz1vewtEQdGVvD
tv0CWt/JmxW9Qj3BpHnEaCpJvaWDhVZNn6dgKnROOjMo+NqbPcHQNDvElPgmp3tR
tXLS9axVvNGcrlMfepcbuYBHq2qUYHUKSwOyV12SJr3OytC778Jl3Obx4c4KUS6d
lIOkDasBGS/xfcQ0/K9/uDnluk7c2DI26O5Hor1EpjBlM9UIg/pGIE261u9VEaDR
w4mzbGZBEXngZnd2fbyA0rTFzLzkijC1MUUuhf6ia41SYas5uZNVIA5L7msew6EO
XNE4GJ2O8BGUbIN6CXTwacXjQp5z7EDNRFA9ZI4wrSb9T3ygdO6t5+qO/zzOTj8x
mRWY95KHTzo1YumvcF70KYJWgy5QCX0xvfS3DrH00tz6ztyXmVSwewCgcMwSQJAN
/jU57mbNQV2Eolsqv3raRzLGvGuhh6kXMDB2IDZXL+B6hJEJn+GfDbKe26jzTWcc
GVwtx5B+ZzUfsh8Bdce1ExzoXyMOZsEiVq2V3A6DnWuafNkC+KIihg+0lK1cni0M
iLH9pKxJ0GQSkX89mZOYZz4slV3JVzZP/NuSWz9E1FJPCJUumgvOJb+G/knMI7O1
zIwZ3YgKYa0hNncpmX8JYrIqiEbSOpJ4mok+TLeG6MfPQiMcIfqG59uRq8ZZ6POU
GWbV7WRMlLFBwDisrefaSejFE5vUjt64CdbHFyhOuDECaGyI1S51QrFj9gPZsIq4
lJ2xFcHP7QbGFax/BAYRKlHVyT0I5bbP05I73UUSf334rL+G4ad358aq+/Lt8bxA
WhjWk6bzfX2HlKwjzu11+XGeTTnwtPN/s+wC03rKC2w4J/G6pEBC3dza1/+KuJdw
YZsBcu37NWDRGrWOAlDS8uXVphTo2aMuJ6q6sFmNLA4P4V4ErxTl/4TJXlZKiRz6
LBiYlIu7nJSA0oSL4Kq+My6YvIBmhzs30cW0t1/m6YzE9WNRAHAVXB41u4YgbL1b
nCYmz31nASltv991+rqi/l+vaZqZsrncTOO9mITX0LT278VlzoRNlXgzzIrfdglG
SwaHbarUavQpXu1Kuv3N5oBdC4SQSFaf5ERzhkzplizCH+ou9FWnSAMYs6B1Nc/y
4EF59vKDHQhw+pV6tkKjDqZoVdXbOZYzZ5WSfk2QzYVsqTvK8GN7Td59d5v3JoFu
3UfL1Y2QlN4JOh/yvFbuoPbE+QAV40uX/SiK33aXqcZ2fbM0QM8uDMPyoxIz7f8K
f0RU6wjnFRUICWvHVUl3ZV2PYsqRcqcou9nuTDHoBy9MfPTvrE2UqU1S2DTzGNqd
mzujgC47bduOLLRAJmJOYW+f/iQz/y1lbU5DgcFx1e/Q9OVVgbCwZXMHF9mXp1Z2
zaKYIDNGU9YNZZlPKPVG5YL38QzvPrBenPEbgBA9ZlkAcAUF0/pNWmn3li2kcSRs
NcJEnt84Pdvm7jYabQtrQzJxzW1E+627Lzq6VFlV+7dxNOQ5EtUhrvSBK9Yk9o3t
6IHlokOwd+WKGRq9QFcRyEi4O3955Yo4YGzinUUgMCDeoOx3QS6ZHh+teiZyDGMX
C+mOHl7lDHu7nHtVn77PVVZwisyJ/xTHue/LiehWXjD3mcq/mlXTlE6m3fK1Jd/i
J4tSmjs+tpLFcZvaerZKg+3cfcfkDXHtDT07hvJYL9Hkchzw4EkBK5qNPpV0gcyZ
kFVxdgJJADhP+9lkFTyN7NmA+P047YcEJVhxA5b0XKp1R6al/CdpV7Wq7RZKlFvT
m1aGjuOVdXP2sAyQC9NBg/5BXeJiN7si0URt289vTXTe5RFZn6TnyBEUUL6kjbnB
j63bJpViHgVTIpT7kCa55aimVpMp0/BzDLCMNUyfwFkdtyPORm5BrrL1SodD0BVt
HtwFGh/dBzZKnsWUXQp+wg8ihErizxNsFFM02ZfOWNPGWVQ7jXjGxzRfn/lJIlj1
LmkMB7JXFQASna/RP6qptNZdeb9ECxDs6HCino1wUII8rOBNXCrG3JTKxvSw0icA
1sCZvR8wZQa+CxkpJUR2ivAV9vyCmgu4Bkr0F7NUHi+zr6ZXyvhDZwbP5yaXdxt3
oBr7bgHv3B5b2L6TtwremdXmIBknqrnOyJaxv2Ev8D/yv46HKje2kWA6ymjeTrET
KVDEdOyzFM9dhpakCMJoeRJMqvOrzlpoyZu3n30IxJWLVFfKr0evL3P0elm7uQqF
S7SODMWbvYw9qXFpmpx8DjtceAbnDy+K+Z3rBb/hyN47vb7RoOtdzePjGWTWlDGO
IzyvJ8jbCsOPb4qhfc6v8+GO7Pr0B6det9npTVaUPY7+5MewX8wMtBCRjzmZBYzE
OWAdfIo9JmGfkKgNdF8h82LU4LtpDd3LTv5lpeaTyyDbYGd4ZinRM0/LWO+gPCPh
/pH9zUafUllfw0F/aF3TWeIbKzoub1Ud7fNojp8pEahjtMVSzIJTiZaVwvXflDYC
1huWlaUH/ssxBsVcCgGYiY/Ka6e9nX0znA2KvjGysdnoz/7+VqzNGDwcEpLh97GM
exUHQsuqSqhv3RtzhYMKAFKVDz760uDOsm5G4v7W290FBY5cyJ/Tz5NdFRMkX92Q
PD4TToYQpnNXpbeHFCkRrWAX6HH0vZSOXJHyq3FQzUeCTmIUf0qXBbgQuIdKE9Ri
4bow2eSG0ZxQx726WMzEfSfNNtNsa8LAdDP1Ig/YfZHaPLsO5RK4lGk4cZ1ro/kQ
ENJqWaQZbsFjYY/ITwsXVMJs2XrSPd0R8G9K4eAnq2miWZqOKwZuCurxVTfAzNYH
FFb96jiPxWy7wlGDVqGOz3rMxi4Ty81LkAiyWruw15t2jHaCstyQ+MqXqOhtmxxa
PrURzyHDjbJ5pDcbpKOTKLoNP/Rn234uOo0ocr1a4NWaCdxoZsZ6wBLEeTcBENmN
9vmb9qKGAv4Cu5JPIGtmKaNaYqKcQhyvUTzFitQl7fc5BAFNd84LvWy6qq4jjAh+
stLZ9t780LGsUJI1iDuHz0VA5aLX4YlBhZ4z90ATNAAfr2YqPYLymycVShPYpUx5
4nSmVSaGrXWGea/Ra+0Nzgf07lrO7A6fH0Z+yKvlhOYnZsgcdBEpy1EnNKPhuIVN
LR3OHxgjcaclkLeIolR/YF6BSReFI3uuaz7YlXU2tUKsPm4VF2xN2qMEay8rPsNc
oQewKKtzj47H7CC1ACgyJAAZzkV7K2T4higPvyowFaF3LAQji2bDL8cJ0vRAxpxg
qSYviW4plELSFCel0G05QvCH0jstWVq9qBp8pY0FZULabp5OM1q/tuPqIw2TSbwW
g6cf+wqdTyd+9NeYquFx957S7p9lAmsXj4V1abbf4pt69KSjpYf9JLyntf7RNkVA
+pVx2vdWkVBh/ABOMzqfF47kAwpwzbZ6TWyjOxlktBUT/md6BrzSeuhCbcGsPT0s
h5fexODLgGlXxvJMIwwk48JCWQ9SPYXPhLKfptlS0n3U6EkvY/uEsf5bKa/ittSS
JFcIz5XRZX/Sgw91GdEo5zcHu5K7+3zm5LSIhv8LSgg0WrTOoehVN1AOaWOy6yKV
GI3wPtHY3uh1/du8yfzu5wBlPyXeHHCk+df7CrOHFrzDQiZfIBRZl8TXoL1PmfS8
ketNAHEk2Tc/Yi8Nr5ObASIXIYEEUzlGOH/K/l0soWntvjmhCp2v5Rox8u7JHMsY
YsPvsYhxKtoLU1nIn4NqaGpdhELShioUvqbbT3yQaeig6OwGd0xxWjOiLBLT1DoV
Wk9MlGQoXWNg7yLxN5btD59fnZ6uBseJ9bOm0Eck4ME3EtSRw7cJC9QQncis9LHq
VP2/jxm7CFXx99qTO+nordV/3Eu+q0IVkGNd/XZNIOn9FlhiIZ7yuaUxkix0M60H
bm+yDGYFCCHFJdImdW28uUP7ks2xSBmCsxFIgilS0WLuZjhqrQxwuQ+PhSygvEkZ
I+0zt4a14Nhv7O6qmp09s+NnlU6E1ErillpqoUIrykOmXTvyKldOtuDgDNB74A99
Zbx6LgwgElhH2j4EmovupAzlFZUncMvqUaN957O9H0UyuYtS3q49DG/nwCX07eE3
cuxAt41rNJMBt20mqPiegoEYIBH/KdmjyBeIWguHChTjUvYrOKeoiEesaIbzcBAz
jBLjq/Cs6wtauEUaLjwir31+UHof6dPoq8cS9cH56t0RQzw+o8J3yMarm6icOYXr
9v5BsM5RZARmj+u6sdND/6RnP9l77IxivvQJ28hNVnGOfgtVn4WBrqkQxmxAzbd/
xhXVnzupIHmTOhE7E0Cp9qMkNMHfXvdBlZB/b0e943YOSeztbXM72ySCiuaaJ1Jx
hX4bE7MA28xQ2tNGAbJademx1zItIU3Pntv+xflRm4xWBktebZ+wGPxw7pCH7Pth
Sc8nXNRK17F8US6S4cDCjYe0IwUSHW+6+uUs02lKului9tQsBZVBkmH+3KAWIlkR
kKYGscmrKTjcG9j73de5Pm380SGRuZ4vLNhSt6XG1gRPn/FK6Dcn5e7RzQ280wfQ
RxbkXt5SXi1br4FPvXsMq4UQWsHyVKAthnO45d9zb8kFGTtIxYOcyW0G59SUauOE
+xCogbvPs8XGt4/Lbz+yQYJrVKL9IO8LTac4GKjFumvFJGe6DTBhY9JT5fxTDA2L
RbOdjke5+4hi5PQROnxPovgN4oitwgPVXQ3Kq0xXSMJOS5JxWJAaKJVyi1zmDX+o
/OmrX271vb8twdpZWVBlUj9Xrxl/46spKTrGNkFWdDnLUioSK1ufl39l4WppvBBm
qWdF9PETy4weHRfvtvBR8Rru7KFV29AI0aeQFflyzAdhhRovIwLKB/10u1jsX/6B
S+/lQUHDDRiTDkhkInMZJs9IgrsBtlJ/rY2oKu/E91S48O6hmHcGJznBrUYRSZu+
qlw27w2jsY7N9axEhA1471RuyJRDzMU1QuiZkFfqDS5Q6yLUEbdLZLzuW207ly8X
aYoQkzuQ1hHVvDJlMzu34iEqiOZWH6bWEjPAIEcxjfyUO/Xvyo3LUR6IL5WfU7C9
Gad6hC6Hr8X29zz1c3f2NV1vKUOnu2quxaVeQglwqu4Nlr7M/d2nAz0wlR055MML
9HuONp5mcLp4HO8LjQ/Xj6LrAFgtHT60Uhfr19ShvvSmvXeseX69zC+9hI/+4wE0
FgTotFHdhGhnqQW3jvVPpdU7H3sc0Y35KidT6jeXWuG0E7+RBQha1MSM61v73uSz
cgWEYHfEJ28xXXEfF1hXO2uxe/ec+bph08mugV47qYYmHKcNYL0qX9Uv8D2jTxUF
ubYwjImYzFne0Uy/5U507mGatrmTZocbD8DtgHxIjR1wPf0VvO0Gy/2iVMDYLv47
NKg8qngqhOTYk5e/h2sV8IMVJ654Ifu7j7hnSqGu0U+DNtcu1wcFGy/J+Pdu2VQZ
rhcf49hx4uGJS2WYaSqOagvm7/AerMuW5Ht4wM9a6xSuwbDtk5CvWItLUhXsde1d
8WFy0ytZD0uqtskxCCIFZ1zqR2XlX44umhH+Q1XH+QAgmiGB3ZTPW+xe8HIu7i+n
0et1xyeUzpH0fMcdBDMREeEyke7nc8/9xqOEGS0y2ACenxkFjVvXT5dkY2camtDs
S+fSiDCrJi4SNmyYE5q8RZPz0sQbebNuFAqtUIy4dK6wOl0x9gMVmPCgfEqD6ckj
+F2H8X9zTTJKs3UlmbbfTmekA4tmC3YvMtpI2+2jbA35WH7OQQFri1uLJIcWLCN8
pKQRc8k3K5oJhdj5Zqxe80BwoYSQdtpZ6mZYrmbhrG/H8frfYpH2kcfpIEzb4vPX
mnsRrFeOc0hYyGPhH178yVi8lRDfkwTWI6mPeeshWaxsh24ODaGbPqP7Itb18Hh2
5LHfFv7DdQykl3l+CELyuvyjs0w3dRsYX2U98HfO50V1Sjfo65ddfkT47mH34N8d
B2et38C7zdofR3kas8s1naknIJotLAuMd9lp12vLsIRbGp8fwlxqtH9C1wqW4Qnz
DV0xO1N2+HOiaPn8Qta9b8N9OzorjvY0ViKtPu0HgVV+a1gUOyqG5F0Ind/rrihP
NRpkPFu2CGD6DSeCLu7v6/VjV9RRiuOCxZPHfcV0qzKENMl+joY6mbg0tXEpOoVk
yvvGXM5rgoknc1tG9BL/1TeRHcTcV9piw2J9NLuVoEi08mvRwx9EFuWW2/gDxO60
qdmGhvt04E/3aKxc6poZJqwFNCkzme4hjXcbDtPlWzAXfLrnYH5EXrOeONTbj4ib
y7pB6odYuDHLdEPNkJzk4QE2/r2UVpzF6547YeFGFaonv+gEBxOz7CwiTGaCcg41
0tRtoWWV/nWILgdqeS755YZr0tiERWL3UVuG/ANUz2Syv/evAOtuNTrpU+eRCBSf
ae3Z8WFuLjV0sAgaTTci2GMi0ZAIWdjCbxBfRV8d+IWlwrLXnmxOJD6Tvm3aJWvj
Ww3mzY2fnsRUqfQUAv8+TyLmdK1crIlQmsPIjnzIcqk7B6qCdUUzHQas8f6cLEoT
wMYi7dJRW/yT3birrHhGNq/s3ihoebZ5xEzR+FjKkWHYB5TzEllx+KeSBtinxNm/
PQrEoT5SLFnJeQeR2v2IIM3dXM5paHEFWnJq210qdBmm/gSLSKuHvDtU50K1CXui
el1PUnWVTpr4ObGmzLTpC8oX7MZAdCFw9tc+kDVe4QGyvKOr9nq3OHjAY6wpQm5R
hNfEr5hM0cQKFFFD4XQ1n3K2VgRqg7Vv0v33njrUzhDDv6yqCtpZEiP650MJhuwN
qp2sCBI3AYtezpAJdfZ3djUHzhsBnprvRg3SMQx9gvdd+6IYCue+VO2QZci2CFGy
+pu5oEdsicKO7O8bXDaFjk3zdmt/rxAC+ZNgp8X+tn+cIsr71eqeGdcbcu5rhLZY
r6wEURAk79VEaTU+rls4vd2mAm21zb7PycznZkl/GYkyJ/BqtWrfmphs8zqaFtUo
69wupTTeUBRJFvkfd3W8ULQeW8qA/WuVkWSZta1+UyhIgnhohj1iom0KWQTxofoC
fleWrzhcsA7RCphV/Pu/oU6HK3RNFPwQo+QZiQ7NRmKe5xmH4mvyjsH1myIesua8
LQyFcLpgIzND7CTuHGhfXYQZ5BxcyKx90oN742MRVeUjGpOcGwoxLkiYfcUOaCaP
LOl1ZuN6Bdkxm3nY93+5QJ0H2vrxhKSuFLZEdsP9wjG3hTEMdFlRVfHNBarXli1v
WWPbR7Pa7peW1TEnGFY/DdWMXIg1d0nQSQHFS9f6NczlahbZalb6W8+1Ole++GwH
vCG91b2LZ8IIFsaaq1q3pnPpQxtvuZ17pEtulk2jNsNIcnhKfTqImfy98MNyw6Ez
SdtiiB0I/w6iWIC4DAmQFNgDmMrBYeyYaJFohwugaOLVQAnXuxjqjhNSqnw+Dg14
9EWaZ+VkxaDcMVtdW5DhzSLi+sIqvY+7Bh9Zv0gXgtMaxcyRbsuVI8vQr/8rd2V5
Phn/iQYrOJoFzejCUUDOwTqqdJUTah1wPFH3+LbsR7KSwR653L4xco2Z6cQDTw91
oWeVc10op21aVB7cMSIn4Ypi2StH8zqOtqAjdNC3t0HWxaKaMaQmwYH8+QFIJhA+
KNfigPHTVlXO7aNwnOYgjrHgwmQOgWYovIlzVE5IlzspZrwhRU4A+bG6teXmqBI8
ImGMYrGsBZwjSXIcwjYnOluKOlKdSSK2k65OHN/1F2Eie4xOaPkdn10fpHqnKL40
6UX7DHy/Th8jYYU7lw6qC6BvD72adoXRPRtcs9ayCElJ/vje9A2V9OTvF7DEl2v9
C0XS8rOxojIV3S99nHuYUiuds7v0D4J1Jy+KqW10J25W+0GAqyu6hJysP8RRZB8D
r3dHiAjTTrrxJ2F5dyrZZkB2Oz+DOfOC4HAukkNXmGw9//nKze06clo8+6pqUURy
+l5RtGXClvTrcSLd8Fc8txuFZSv5NJn6Wk/WhNdDIj0yBb9bbqA7yB5F+slP50I9
gxCojoX/j6S+F9R4iN1cFqv7TQ4ZYTJUeaLjDsJbrtFsjnQGofZlrH4Ps/mSBC2k
zf07NqJik3KKR/n61xFQqSNjoTYs0Yq0batybn02UNQZ1VBAAsLyf82CO4odwtfm
7Ojq2GiOogycMbTw/WizyudloFbZ6fTCHBFm5MsazsgWYzrwf0gagxd9FjIuJe6y
EsLtvAq9lWIn+IVJU67YTi2Hi5dlOGcge2ga/pETlMY4rYvYk+frtCQG48ib4lSo
AXaZPrCDRTLCUcDFgiXqzYO1EMwE0et42+Rj9UcUhtWEGvAWgnavpRkmPBvGqyF1
j2S0obyTBxY98UQPwaVXMBSrAJA9nqlw3jvtvk23ft/OD6iaGBi55dhCTjRTEs6y
LLjjDI7kdkMax+b78ehpbR/jmyMaVXIml6r7VexBZ4RmOrimiWZx/q7X6boFjQQz
d4NCzQWfxyjYOHK8T94HWd+5Sf8ChvBU2F8xWZDFYpZE9YTVMsxy5eKhictXyAyU
xEjBkgPH1278aoKARLirp6mQmgT6RnoJDG/Tn18YkMJMN/fBtQq8qA+fHPm8bZ1V
cAsFT6o2wXToub8BNBD8HKrQnuF8ZW/DHQgSqcm3jqMcfzyCucdfaLU2kKW3XDH3
1uTxpxLHcXICnAlJnk6srzGt7KBsr/KUEUf2wKCMi2tyfR2s8saFV8kwna4YQWdR
7tmMoDlAFt4Y7zDFVjcel1+d479UfmTlL4vmzNa8uU5hMvh3yY0RnByEUDCVb3LW
yhm/qcu/pqy00y+MhkKXRuDSln47oCaVYGekQlWR+a+DGTKNOKJtW3rRBw/OY7Ny
dNtBIFaTOSwRz2zrrdHRrGkhWwScG4ERofLo+RKoegX6qV4KbGr344NywIbwhNzm
V1VetlZbgQJfhWa67U908P04b0ACAcjWFhinM3QF511q2q+smdmnng+5aegU7vga
IS/JDY+NtS0Ak2aMwKwnM0AOhpyyccVbJla2aqbWrDlxa/HeeOMoTMdPSQDyxAJ6
gviLKj1m1RdUeWpjkQlcyEKdytycBBa09bXTD7e9UVKyo4QPxM+iFY4+qx+s9tmj
KrPZC9BtBnS3AA+bCRp5kKvaGlE/vjxzTReayF+oERRsNYdWPGRwN6M8W+6K4W9Z
o2Ag9q/KMLINA5FGdYe0rNJuBYzrLDatIznuv7BKie+f82KVb5N+1Dl4Ez25+z+V
Db+48gVANrZHxaVK7UKBCQu7fohijwYyKeGmizDKaNOL6XBNXWPBPavNnrHJlXJM
kItbbZLzs1KSZ/1su4DOoHi8XHtiuf/BKNXsmVpC4QgianpfW6/EiTRhZgbmuv3E
Ajrl/qKw0tr71v4HYTzw8CnUztYKaiFiw//L3t0ea6m1uVcr932ldfwjui3wYYNa
K25MJyCeK76Bv36ZuFIlC2lQCVlv/1jdsamExUAhR/NjuPqzosVXYcfSDyAQ7KQp
xRq8zWhvJgp2kC5rcNu/BTgd31RxBWTD13hUtp+g5TfFH55Pt91+PXFiV2JcgO/s
BeohcFj45k9dEhgspxOOy81+8Ivhrd9HtzvdLzMVzRUqEEGxuAC8CpF//3KDVKLj
7+PjGWe6j52b6376I7jcfGDPym6FvQl1tC5lmMFNSihv59gf00FJ/9XvvsiEqyZL
vMMiGXQPAi95zUc6lB9XyQEw3DAWMYFXUCf1pMaAy2YxzC32nrcT2aLEesCdsiLQ
C2zKgDvcmeJJtrNt1PsImsx0k/7LOw/uufOeRRf9wDCBHVKCIM09G4XEDl71OW5/
8VvMim0/wNNjJ9sVsFA+QJLbVR0KzG2ycx4oQCqDr9YqDhjgDHvLZk5DvDBeoYF3
XgWFcjAKlwOBvDzCRuIfXsxYwR9RepqCYSntsMJ432sIz2BWZ4105pmTNkQBkDtj
On8Sj4/XgYhjTxbB5slvT2SPXOGI+kWyyrQ8jSCtNN52vSp+VwROUdKCUBRL69cC
ci9Qv5pHcswcZI8VqGeM/kxV3drx5vAxOg/NznOQJQayiJZUkGJmkhuVfrMst7Z4
cq1M5SgpVxEZgdShqR317ykxi08Q/CEH6iw1xRYDEjYDPyC1Xk3mpK92SUuQOw4b
laO2eOZ4fC1+ZhsXJEfg32F3ENao3Ghx8Lqk+f4DGLO01U61Vq+UUzKwRRaGEKrM
OqnqUfVnGwjoDKfda3RKUJVsbQpoGzBNa2QGq85YClx90yA8+KW4qkNvrM+9uqXu
N06TAUxbxVPup26moKSUlzXIVz8kwvrY//2xNh5whg0Wl+72bkIKU9WblKipU1Cx
59ndhuu85kJNdTDIUnmAAPyXLx+oxllPX6OR5j96D3xd1kL63kBB73MPjfSZOeD6
GXp/Rk9oM/jRyDgIOdYC1ggRXPhKZK6/YFeBGHlGdwzWCaeKm0Y72IgnBaBe78kY
0+hmxMJQ63UvUaetG89OhzZZRailRApXotKi8oAe1gI790glqOpIRRpfz7iIL/6A
`pragma protect end_protected
