// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LvE37fmgeDc66fgyMam278eUBftxBj1qFQpsjnUT+96kXIvbTAS9EXTYjmAlfCJz
wfuPGKUvaE+w4rbiNaHHRiPbH4U5wUb+76bN5AxylPTwhtm2FC78T0D4blSQtD1Q
zN4HOCwETKtDIJ1qoaqkOpjWwhmoDT4InuKHp3/JXFw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7424)
MkR5Y/maqOWtR1cbALq7Sic9qb7qv+A7P3fntjuTTbnwDTvFeCd2k2plcEOK/QeF
JTi/pQE5EZJdfTg+z/uwKxQVSTmOOeNXy0/2NhBadxOydxbsldR9iPHV2w+P6s7n
QidwzwHyUN5xM/JmJjZaq6yG6e5kHzhaEckcC1/xID4QA3EnwSSY2FZS0UUnfqKz
Ax9nI7ZE4JHFgIdVdTpwsIGQsrbDj0Ec0QdDM2BG8FDvQOMw4+snbrJo2+GRThi/
QNnLgsnEZxb2RKzsitlHGx7erZJ923ssmsgXq5EXUAPPXd26Hwmqi7iZ2198TH6L
2yRcTiQMREsHqBpHpYndZCY81pApxgmxjccHfjBvbk8CDWz+NgmXID8R704x1ids
8IYl/iey+EuoQMl0AhTVj3d5rlnHdMr37CXCff8sVH2/eBxRAjG5JLZZmxwZ5ZSz
Eyfe/v+73FJeiMYEQM/tQ/W+VIsL848UCXe1a45st5J5SeZFTJTpyIDichXQODHA
/by4HrEJCQwlMCzI3N4iGl89UU1BbrXKy2yT3ekjCYALckY0rbhJ0iykW0GYyPD7
H4nCtrWLKFIdsDUjDwz5H7qUmfW6DY0ydOr/Wndu/ia1OZvXGg9pfBBwXvzFpo5O
f4q+Q8eQNvOH0PTbEDwRHyNihmGsR1CMwUHrxog6RSUWb6o+I/UvEZ6WVHzKuGoa
hv/CWAKvwSdsMrbA5Uv891mz1vVbVClqb56pRETWZVP9mf0/YZsmaDttpgaPz7GT
zRb+DLJCkWVchF5J/hXQBiMjxdDiaSTsStIXiB1fuEus0Zb/kgMUN9zw1DXpXozf
IzBwCf8ptBqcWwfvdP7jEbilsfXF4VQRIPKEVR/+Ls9ctAPy4u+vhskTDvssAyxi
Vj9NbMivV+xbFZMJwdQF7BUl4sm0rRouRYAO4HvUSPgxZOTU07bGwCpy+JOZW02z
QpBqywV4UuNdoaeIKvmIdrPvU6u52cqylg8pThORe9X/Id1DjdWHfgvw+cKt1lYp
MuHZRdWzUwuUqWgwuOKcAz4d6IKbe+dkQaIik6BFMx+Guy+cMF/xWwgJOEvbjwuV
CkAZpCmIwHXj9MyeQEwcKL9m8LYSqRBmLwqJeCycwjT5hH8ptYhNBQJT/iSQ3+/9
N6dL9C/uBILZbq+Ob2X+E2x5I2IT988yRCJWt0EF6ZG9piPq7PKaVkr7hXUeXxtm
BLe4+iJKoJ/BrVQ/FdnnqgW6mBlYyVYnrGwg3PL6h43fe6E5Y8+/bUIEpWo/deum
5Vt6aAinkOyNP7fYiTcsTPsdcA9/qqLOb2AuzQ5e+M/Zckm7+xLifJuH14TjIDu7
IYdsaeW5xqXIk+Jlw6Ywf6XjERVAh85JuHeNd2HZ6/9s3ZO4xdPNS270nrSmWEyh
ki5oJ8aU9OLaWOggNszZA0678BmdsIkx13K4hejnhuDtxpHUrXSzmE3AC0FfVkxi
P1RDVETqn0452TV3h7/gfvj59F1a9TQ1NmwCo3MkYRkilLhhHWnOKrWfdiG53gH3
EkuurlrtVY2F9lBHx1rpCGGUz4iwz6Xs2CIovVdtJsP4inwooKag7Z0lOF8r0c2k
xrbLfk0gqfYLuLpSP+fDH03XuBevfJ4Y0cx3QgILQaYL8Nne8wwmwmhFcGPTDuFt
LXo+Nev4Ng+bgKTCheV1M6j8PCsxHvmqteVEDAKU+acK/uk88MFsR0MUPq98p7nP
ZeZZ5IRVhiH9huj6heL+TAtQFWF9iR/BxdLzV+0xkpB52s/46OIxlTXzwPqivHdi
U6OQ3FOiB/vrI7OXP7yxmXr9n3Bw03FW4CKbgxXGnhrU9o8Sipx/C8gpj/AeDVd3
A8oDmwb5JS8BpZk0v0EjC42dyF4GT/pQ6Zd/LZ0O0ZQONPpE1cb6+WAp+lVBBmhd
/VBLhEr0bbsANwmUQf5rG1pKxUvsPLbWjZFpxKAILhEpmgbB/dhWOqFEFwEv2afE
4ejjQmEB9wFJdx2PDH4q0utiL79NLVz8odVqely4+KxJ01cBrmv6Z3DrUsvFgqjE
uazaQhjRn1FH2p6SSQ8aGlC+gM/plRxhucUtyUlOdzLHYNrKQ1OvBUzLAB7z7+SO
GliO0Jk/e2eO/WgQaZ5jUo32c69Hipi5ym/7YZSrn/OcpvOAhJQQnzHon+fBgFc+
ZpzKDPbL9HWS0csFAdfN9O6x5UwWfxMqXrBgO1XHLWJSJ1TEM7Nx3jaF7S2HZcvN
IF+fGXbHdLdXr29Z0yg5Ns3/0p4AcJjXP//qRCzHi7WMGUgUvCl7HfArzdMPOPrQ
kLMG8PLZX/VhQFXtrj/WrR+ZNMip+eA2/YGY1Hv1qVDIZ1lPOeOnOMEaqfnwTHwf
9PYZ32bTn9R7IQHcGsjxrX6sy9sJwc0Qk2HNmlplmZ1K6FI1c/I8D0lZF5OpLPWx
YzVTpvYWEWdAEcIOirSpuR6oCKx+rB6LEBQB985v2OMizZpiAWV7UvTBCOD6t1II
hrIgwxR4GmkxS+cV3UQzqiN/r/1UjRmSA/dElg00SEORQ5FkLMmjEun8DgzS0tHo
CFc3TIWSHf2G/QEaZTXG+g9y+JI8WEXOkb2qgHiVWbeKjhVzt4KFTq3PGmD2FmbB
3ULmEvXy6RUUq2xXhZXprX6hCF53T5eQtZLqUBMEiDMk/AoiHjH4HSv2Wy3K8lW/
6Prhmz3daosmCIbqlbbqZGH4CyvfG+nl5GUALYydDdrwN5EOhJ+F4/PSHSrsH9Nb
IJ7mLdLX+4jTo9M2q+xWXGDHiryslG4Qlcokwne+oRkeW+0SxLBQT/+Xyd0hl8dl
Yf9mnnneL/oQ5QOLBOtyrpiBIY0V7x+fMji3l2NyZ2sqjPCz9CC90HWd9ywUELCg
ZFYPIuw+Il9JOU9WzkZGDW175Qb1lp6BbN7sBubtktlldwVVMlnt1yfRzRwLHXKe
rRoa34q6XhVTVI4oKnIXsLPNZvNNF0t/+qGb/zHyi7SGAzSHm8jfGzr6KCAnnjpn
o0YQRydoT75ZVUjoUeooqBBCvcYn21t7kSPKSyd88FB4VoptGNVQ4iuHyi0ZrmmJ
i8iu7VOPVSgTkJkpZYHjX5s804BvMrP7DfmeJpwEAKNoycD4gR5NjBvD+OkgaClO
/N8Uy17ul8eCaJ/18eDBet8QJe3YYB0mA1TvqJvCxKEINgo8BcF7Ssf1FbAPcvMX
d0XcpbkXiY45mhTz7ldRnmt7LRV52ykeyh3AgCwnytO940fzajbsuO/zzjCL484R
Iau9ZFXL8dduAsgN5PI9P3Qsh9nKgpnAh2xTaIPMPT3bBeXJrdgYvsvE79CAJbF0
nvDboUFao+Tghyj3HjkyaUOT5afxa1LyCI+bH46hJytyren6w/sw4c4N5prDHrr6
TetK7E8XwO1yCSPi+UA50wEmZ8PLZxnJUh0hZVQWKTmZ7nUIj7MPbdsovZz2KVfA
JVVnYOgwGwMFTcIRclRFMXGhHm2lT0ZLI1hwhlJ9MV6GXSRfcff7lcMbvX+s5V3s
7DJM7p6OY54KpqCxTZ9dkc2PCiPWN/MUtvQVscoCYKs7qN/Rn5O+5ar7h4Dcw7Ti
Yg/C28FpoY94WY5mS/76d2mxkIuhr85cWAtk9wlTsZWSpgSkiThEFyldZgIs3JW4
E0uXkhsYfBSJLhlEceSvaSEEUSxC60m+kLsIbZux/NaFYIDQPfSPUCxGU2DVUmv8
uDJLuBf9M6ZPeDnteTvnrX3VHdbfXQCydlZVEYxodLCKq1XBZUhpTXByZB61T0x1
hZndhWmNWTscTJGhk8oN/9Kdz51Vx4O7j50yuJg/Q4dcvJtR5GoOFkbP+XZx6Zsh
ns8XslxOSPftU+QP/+BD+mqsq6hhRmIF63Ooky+gxUNqknxTgjhDBUFP1HcTB+Tm
OMRZ9BC1Cuoyryj9TQEb1UfBDoT7oG8Y+UFo2qZNe2ZOLO5HODb1JFflRt2UvR4R
h0XqmjqEMsSQVBoMZdaL6BBqf1hKscFIjN893kXuOxoh45XWKDjQAil/TykzNnCO
OtZ+IG3oDMHz2FbP0I89fdhVUKsG8Luslqv/M5dNrLfMuj8wZR8Ro+kXFrR/U8We
P3eOUJx44ZGFVwbWKCZNZB0mtv9ekemspZTrNIn+3MkUlXNBp4ftiAmcGomPNrBe
0UhXnuRYM5khAPpdykhCqFmF2RpTcujF2yB8hn3cJjJCwY488e28yEN5JIa/IdKf
9iK6rHsE4Wh8Vc0A2m9ti2lmIjlJI9mpsm2Fw4nw0E7IzhYg22xEUw2emEf8VhN6
a5IzEyRBcbdQkqfuVX6ohafW9L9WoLY56DSMiZy1BJqXEsYWdSQv8ggBGbD4J7ML
Dcw232KbJDNruiUwPiD4fp33UQ+QhqbPYQ/yBw5EPT5xUZwutxO588w1GxyRZceC
0COsj57pmS3hYDzP90yrSBLfhTGfQwnchq3lNpVDDVCYrdmMLdaS339pb8bR19Wq
zEIQpCDHdrP0wpwNzwZRViDAOsOFMoMT84/LSVjLaRRKc7TsQayySLn+kOVI8qdQ
EJQ9l4QaWn8zNtI5dGeUF7i9eBQRWWzZKJap8rOBaVXSfRVCoEwRGYCFe1T1uBmE
7GGYuZwya2Qj2dvVl1uFlhsGIQTypo/F1/NzqutHTr68WR5YIE5NkeI2BRjvVRef
JLfNi85M73/oqDJKZm84n+Tq0VNC2jlP/zmriTDfDP6b+S3761kleiZwBmJM4cC9
WTeE/UvQaHRx2ZqRgon+dKEQh0mijY9fXmbbcx9WAhWqJLLWQPm+5HFE7EkkldbV
sMdRouehQZtWlppv8gbNJrHuU+jrG7Tmh7GTSfBc5zNZdh9/zXdIR/cyZDYzshyy
fxl3EG8jOh7JF0ann3LPzULOq/iPKQISdvDubmJyCmOl8qd2jGKvsrwxGQhCB7i+
IPsqOyzdUNZZyApHoDptPJJs6QLnFYMBjcNl8UTE6BlyeiIeakdJmdJ3AHbY5AAE
k6JAGgTDFMwsWsSFd4GtDddsZtTRuZvjcvYcD84L8tbw9VAua9i26ADncdd/qmAB
oPSOWVIF6/2gIL2CsOF6t8AEvdjeAGycmAjkoC1ilbcT7Fis8eBOzhTVP4EzLyVp
oQGthK/KWUfxn2ZPl/RXpgBS0lfmyNIO1TlGtfNmoy7RG/oYz5acloM5hc2zHjP2
jJYGmPguxL3y+jk0pyOkzDbtLaVXuzS950S+TQ027MHbmGNRFUr14Vnbwr+eDt/d
/RWmXwds5xA9FOdO789cqOGLSL7OPVgpxp2omAHpvHAaalOyDxRyOeAQN26KCcSP
7swITRw7OxXco/7rsZ5kNOAE1yL5S1TwHyoaFjZe2tZhKv7TE/EuVhIhe9igT9Bd
40jujbRybq8BuEnI/hrob7/JWIOfHhCzObpIcJpnGQTXCbJ4m7sD2zlw1HoYu2IO
cZAt2+1A5ELNTExx3c3L0Aqc2kMb0DfGmSjDnzfkDZN8Lfk6HCKjFIirY90P6Eit
E0CqCVRzamYLvsba3Uljb/uaGnuF5Dh2+Udo+h8CpmYX8d9GBnR/BAzvJ/ZCdZwp
jzqBawE8rMuq41rYLOLQn3gvxe6VjthxLLnvZHFRPsyDUIhlhKs/k6CMVgdwAV3u
m5i10vDlonbD+LARIqYJHF8mNG2RPi8a8cm8hQjBBRZkKFkT+tvTZa4EWFiwO72w
+zFZ8twwF6tWYdTfnqpEWXc754hvxgWf81ASA8T+vF23Y6w1N2ouA45p8m/+xbVd
Tk8cFR4MM2+WPvgngN8HicNKems3KTKsG5YN0PX9qTliSwcmToMOouDRfAVikZaA
wDlhgxASVupeXaMUAQqvInQkeFHy/U0o/EEi5J2k903dKfrwnEehjsTWVDm6CiYm
XMqFL/DPhnoI3HCvHeGWscC7tb97Uwx78givGRvgkCBzjvLPPjWLUry/zfeSje3Z
yTFyXeVWikauK3p5jW0AgfQ4RZQvkhqJSNueZEUwz/8gkJka3tccco5f2SfGPo+k
6kbR8IXTpfkOkSylJYLNyi17zx98/P+xSjAnfvTjKG4Fj0Xqtp5eP9O8bZUQt9ez
MxlVJEpTPWfxL0vpSselS2Zh9XLQLwlAReK1ENdY/t9uQOlvj++JY0ihDQV37Dg/
Coishh9s/1jXvpameCZz/fKzpwltAXoTXEdKYvRlnDQuSIoYhXEIpMGA+QaK+p9u
iWMZ81G2XNe7nFHoLcrTzBHNs5aD0OuBr8vwHNhWDTXY5cA48Q4UiL8zEKic7Gw5
umz2/C7GBe7+EpgIapwSlyyuIUSo9S7OwzTdRM3HNVdJwUpNA5ncph6hPhjy8T1C
Y7kg5OgM1aRakjP4kGg7t36GWfWmc9fLYVISp9FaViobwXMpASAWgXR87aCK+t62
roAbjg77uyKyVkPgqw3kiAzx5xQEayf6KMfuCwqAEww8c1llN2rFKkh3fjjDJ+dn
rdj3TLNTW2TdR+7LzbSsZOoODkWZgElHppz60mIiRdl0oJju3/VUwbT7UFng4cdZ
qCMvgQIMlTLCeqM5fieqIL9zrfv0e18+W82g7bcMes+x/NvSD9zMWPSRGCrDVfyf
eme4mwsVemzg0rQ8VKiNSsgLwOd6gEVxSJi2WNKhdj0ScbloTAlfCTQsgHXTawAH
UPVodwptjBDgAHwSyAUpoH/TGh0eMULPqePLGp711qb4itvFtkWFGqDrv8+ukbdJ
QjCb/LH4R6CcrdXm8ieCPryDf06udwvllEUSmiFDcLGdFWuX63a5kjk2jgcHtElC
FucPt/VRBq7SPwUNeXI5eOKeFGmEJ+4Jp9HU7RrT/0hiuFJZZJwsHcVsppWvX/a7
JK+P1mHcNTxlYp1C/YAiPZJDPjiYqecgM7DAz1fl+R137PpwpTLhgOvRKrsC9uRp
7PEI3zQQxLda8dgK9TFXRfQutOAXrDc1S+b6e2iSU2P3BacFoS5o6QbGprXNqfiZ
hoqRr9H9k+zIOr76n/o79iYOtBJ+UBNqNzOCEqBv+iqsWgTwbRZ8S6Cn2SF9vxFo
MWOnwld8qbd2mm1Uzi/358jmidnfFIMzU0WsDwxJ9WZHj7MMlp39rJcwXILD3tHC
kBiHLkzIIikMybIZV9fEKEqEP4EzKY5X8iVqJnfDzJZAM4zNjGT5P5OHfAVqbRcZ
Kw7IMyAR7NHdpBEZ3B5+kJzTeod1r5tg4vAV3whUQu8ShshYADJ0Dv/GCQFKli7C
axVhmudQVlGj2i72csydb3yI/r9M7cEVAk4j0uRH1B0dpE+suhVeR+Yww0jUC4Na
vnCrpUP86wPCNOlp0BLzt4ki6LNnq0J4qHyoOcxBbr41NtKlxdZcOOMQiVQFXn1T
2Q33poxwkJHJ8HAFi8nMh/Rb3dFwii9efLqrvKyQ/nFGSJiz/Z0f6Eh27WuwEJk6
1FR8lHoQUvr4Xr4Jt8hUDebcnIE4qzM6OVDkUU+fQqGLZftUMT5eQE8ECdK+sc2i
bnHvGpSB+PBwfhp0blsVBUIrpjCew6CiD7tu+DRqGY6HA+bjpDCbzXdozXWSzqk9
m4U01RipGXqIkxEeGx2UNpOczldLJTg0/1ebdPFqLuCWbMApIapBirypyXlveCyM
LtPHwgPkDhEkILlBOTAniBWDcy/F014bh+uAbiUIMSCxy6GOgeh5bJ5vAtfUqq2M
QCxeyut0fIVpf4752QsB2hBPxAbBm5kJNl1HFWg1XW/fa4x0PcqSNVonk+uLv/LU
leXFX9tA/pRb9YsJvy2eAzWRkgkjepEl7vPEDxs7uEUrTKELP7rypAub1+rZqUNf
OBIHOp6TftnazYCnWH+LFn3x7Ay8AS2DwZzb4rARm4f9IUXc3hQ9DL5vcyAIKyfB
6zenmYgHOlRWGoEZ8m4N4rheh3nVq3jBcHahisEPtryZhUmceLQUzpWkr7Z74SZe
tGH3067qIE0Dmk0+zl8STtsTesMLq+ANyaYBPjB/XbeZUSvr0Wx2oP2eQ35fUrEF
9aWH2+jfAx8eMC/a4gzv/tWRiCLS1w+AAT+RAUZAlkkiAxpic7vUE/sMkW1QaJlh
YlowIMAe2+1CwjQtwc0IKeUZp/fxHUCLfaqpi0epLicfrHM10M9v3UruE5g6IoGI
G3JgOBz8AxXIJ/9YfTx0PwmtvkO5R+uWxPLq5KekYN5zfb9TVZJIhdMcfgv/uT8F
QUXBJIrIMOG1pSenTuKjj7VoD7RjaqaJV0FgGhJWbwveHO+rCfOfbnmI8L91RpuF
Q/H4rw0MWXqTSAPPixH4lGEIXZtY9j5pMzQohUvI+JvPSK9nzJkK0Pt3Cvvano/D
x2RWAkfd3KzdwOxxF10LemCH1/wmIvRGAmFUMPxsVeVDk64tkm8FSZS/iej5gSqf
S/6vwrdc+f263alpcBbTdidh9Wf7SHoK4ldFdNYfSOlKantu20DB3LBI2WR0Pf/K
O6ejsiClzYlm7V9e46yGr83Wrkp1iSzivN9OsC19nC6jYxNox99PD8d3GH0LP+op
yhoT0H4ROhITHcExg8LtVt86qdFCaaRRpozSe3WIhgnuWRuqoLd0XXYI65QRz8uA
bttI8Je4uIEOEx/AUGXWoZ+mPpZ74sr23HD8UsMeWTnPQrvMyfM3yJ2UPmXr+LMV
B6WS8iY8B9iePDvuJGnRt0FbXirtbX/IFPxQki8/jjxA8d5RtGK1aiLFiH0K4BNj
ER6gL3pjEfNB0aF48OaqfcFbeMgc8veb6pN3DPY7IM/MUobDa3cPrGKN6uCUNUb8
WnwRVIkeqGCeaqvXUCpuPzh5L4ZJfaBi1xqma0opx48nf17hLzfP7/xbqibxOszs
kNQo6Wyosz1lw1c+u5mc7YKyHu0sjuZMJnsjyLKBZPSsivXr/nTNQF/ZG0pkdAmk
AqmAXhowBw79qKEo+Km9opqP9FwqzvaeGDNHVIgzC7X9MrVfgN0+yrRvdGMP+Oh9
posGJzLT36bH+ntRYVAdbMBhuoQhjcdCnCXXwtDq9OH5Ye9UxLPK2l0byeH4bmFn
VitT8I+BNtGcTcvjIqJtOZbM2gwktnrOS2Q/lrsgoPCx7IXHtJEsfX1/SWoaVI15
Who8Wc0OSPSdFwBsxZvTNgynWI3sLRmGikiy2XSe/svkRRmy3qR2rmn2CQx51jiU
Ip0HMlUfUEiKbMAQ88RJMjF2cDroE0be6QZDOCufE8RJVe3j9NzuPdKTfFBppH/+
J9Wq/PpHIuZxpphL37y9MFZmfR+OCpFQbdmZIGqo+s/pvPUohzZK4OW1Ajef2ePf
J0Vj7ui4LqmunJpR39sxUoGbV5rZGatSh/18ENuDssDQS+BKvRtrwUloxr7ksMnK
kPS45CIAvteTWyT+Fm0ZVQwXwf9kEmv4EIYyrMLW3mL0a88CNDr+v87oFQkNVZrz
kC0g87h7Z9uwZsff9iNwrcPknLgIMhA7ZS9FKuldONAHC/ZiPd4YEmqf8TbvNR7j
m6wUKaZp8QEvJ+3XNRpkmhX4I4z+O10nbGoZRI1TJKtQGlflVzjuvCRCY6RtfUTW
p/lUa0hxzoOEMaryYgM+qtAOZpj1BEj9sFVEIU/ByPOZpVXFw1aZ02L6gwbVYab/
jv3gz90TUSMNFwGirIIjaCUwXL7ERXBSMYt6ECFGEDpB+2omDTaEwewW9Gimnf8b
DD2Twk3q3oTK6qw6dzoiYeMX/JJ764e64qa8VtjFMXd517/5g7pkjqauu1IPviSK
+QZ6qdDUQcbNHrHS/lYsUCB7E40d5aO7Git7zcUYhuTcD0SBgti1ko5GD3ep1H0q
Y+LbL4pwkcyihSDMm2CfzelMn1FdLtbfb59FIPt7Cu6uBqRlzm0kZXZmcf1oYCKl
LfAXPLUHACrfCmOWCCmULLM3QFLRLoS5PgQlIPQDQCc=
`pragma protect end_protected
