// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
GZkHK0eDIOWlZQnC5i2u577VL64XMkJdabKT3KHcFxt69MFMxXEFFgpe8eKPswJ978L5LNMDPtoo
+4l8kIfARSNowDfqz2b0Qk3eCJbNrho6o0dlWcbNy1yqa8UZVlpIf3xdEO7YhO3yqUWtD5N21WDi
pUF0LVWvXZ4oWlvedvG62sQAajEH8TTY5N9pXRArpEkooavIkGLHG/HC6hd0YaEjzC1ACq4z/KFW
d5bpmJKv6sc7Itqcxl0/+4caILMURZDz3HFSWoCaFXnfk6HdmcrUk1Ingu+bWtLo78SReiotCHmW
0NgjQuLwL95an9HdIuR/PhaMz7SlEvlcb25mXw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
1RNnDE4dazD5sxRPO1s+S7GFXFGN1/j8mSNeGP0kf9SHZmXOE6vD6z9F3/51SaPJ0OImCztj6MdO
+NiWbJ+wD3+rPz7oExzsAAfv1gX7WQHuCBz4J/C4bjdg39PKSBJQi82+Ci0Dc1TqY1DiOtqprPjE
JazM0AoWwgvqYyfVo3S1fhuqqQq3PBK68/6wareegdzNwUORXoxBK8TLHA3jooSL72qLYp3FdumA
eL1JxabRGd4jYUhoxgInSZfDDkO+VU6hw2IdWhvCiI40Imfc+B5WmzQ7pbVSeEeacWdcGeYJ06R2
ea0UpubgYpSR4Cd2m8iT64xWbkO8rnwcgQ1EORkJy4mgCAkj3f3J+oCzjfb4Q1kWDBpyoA5FSD8Y
VdVzhqnFnXWaz+SK2n9aIwe9tbL/28sfYHGfGLhp1qLgaaYFOWL8uQIZ26g+OSq1Cco4khbCx/Kw
sR9TIO3rHZZZty+nF6ycx3AUZnNoIfaxtgpu/kRbEronffIQdQLEEo/i38cM9kogQsMy1/XQLAYb
1PQ6Lf4T/U2rnRHyBvbGhRA5DVkr1EF+CxAXapDpPutifXFu8WK8VdVM6zqQfK/C4XHgQpuEJQwd
WOfDYHpx9F2FxkUINS2M8wQZJqcg5J+UGx+Txgvs4IFSPK80KKu5vbgLgmppAydRDSlayIdDKJC0
anCAh2iOteMv/gCDflsFz2nSNMHXCWAtenIDHir8egenU4YANbsRp0dMBpD3hW7cNTVWzwCcxiuw
jdi7Qo4lSMHBnI1cXNHnYSc8oAACXey6hyVsTjaPmS8EbxlQbK+1Mu5pPgfTplxxUAfcClYwQX17
NJUKuIkU0CvycLXzTJRnOK/KDXvOaRWQ3Zp1koh6Av52PZ6jTgNYXCyiPEnuiVwjaIfjfdb8WSya
Z0b0v34UegSKozA42A5+jk5qxaeHqEPzPOPbPdn80663UsYDwOODfPnfEur5DbF3SKDp6lMbv99e
aNbtlhkEzJOowgdVS3Rj50nm0ISUEmNjQvjnaeLwI2r5R8uwXxtvPW7qcFQ2iXNZYwUtZcB1hG5k
aHBpuihky6X2XOwt2TypYKPC6iUqff3wvQA7KsekjOexk2wbcIUl96lf5YMQV7AbSx8BoYL3VXfO
aWKFyI7yxEZUfWcMW+TX8ye9ocG5gkB0g5RERmfMzk3iyjjbiX4qAR3+7qUVM4aFZckCK2siIYdi
8QYNbEmK10CMaChSzUZLHVol5tADEJIMi5cZGS5CWcggGKGEdU7RU4a0Vcp2o9Q59sD8CJZ9rP2f
feTohUbY3g1Wi39SWl57T8CvY5Z1drUt3/Aq5PPRdsCmf/VzPbpdgmkVOPVH+wXgCEM9m0FFK7jz
8NSTyVqfMY7r1nYLHsJgbnvXy2OleJcgrkv7oTnhTsKmEdub3M0PtGRqTYOPKqtDEyCv88puKZoP
1FFyly9flc2hWLkRHBERXEfVYWut/5RIyWJMA/w/7E8P7GX1P1uWQeUGix5q3sSzpIEwTHiLQ83/
1ZpDIfWEx1b/GCukBBpNsRFwOIwqubuHSu5ZW6gRjiZkZ2MQFBQOqozv7fLggTvwbeXxVg+R0qlx
EIjdktjpS2WwlQuYO7tsC9oA6pbEit4ywfGKcJDr7uhddHGtdv3ssyz42ghuVXtOTb2LDJ8HEjf2
2Orlsl5LEHCkJ7y1Ios9hqSGddC4kQSmEusSbHs2LWhOxmlbHnlQUklI7+Z/epeHCG+aluAIaMXN
cOGRqsoBWSRXFbZYrbtZXDV8cdgwpKivIEG7xNFk6LNOQh/q5mqk1ZGmh77P/qnobAxG62eLnUV1
tn5/TpQOPo4MiHRxNaoUykQ9ZbEInYHzgupZQPi68OuNR88es6rxUVqG24cJR2TCHrTzE33ife78
vq4HzVGCNYnVo6LlN5uUesd0qPVixZu0+Crwx8ZBGCrJOS/n7dnoIhooDU4jnkqsRBfkW8jQAwdw
Nn6V2kRCoU588P4fQLHZwSfZS5UBiTj+Ipt5aBbbTfpTHJnas9Pa8R053asCGzEnS36Z6q9RCAcK
sUv++E6PfhCh1heXB8QwMxHSwxTLutIPznmeluO7aJzAhotgc6wudjaPVA7gaUzDXTBZNLakAtY9
XhGzS1tQKaX/OJMNri7cUdoS4t/M9wVdv8yYfZZY0xGhMbbf1lqpJnzRyjpU7o40mlhd4G1b9YhA
oEn+JXImUqElkVGS9/1bXrMJKbouJGY+ONNYEjZc14D8+FANZzXdQRfJpVYTVE8qBG1+b+RDmO9v
GEZ+wSTSr5TcSM7Y/HbIRtF2dV/Hl3H6QAJpidW57+/nnO1KailYMK7QTvp037KWD18NbY0IIEmv
9xrbhl6rs4bWVBtLyS1ms3RsZtqROs2KLi198pJGTSRa81d9+gTdiiUF7sCAqyOuOJ4eukcl9JQe
MxrE0xWeSEKA5j67hgzKwHcScsZf57Hcnea9BmD0wboPul9HwqNG7KCMK+AUoxirQ262XlwRlV87
0Sdz1FbSgfRWY9g+8w7xEnLrN6eeBVGiIjP9SBVGfm/Zq2BdAVK1FTszgMQbzjdvn7pzQVgkvIcC
YOJ3UPwEUjPOuevx9G9CsvwpSdb9i5lx+4L9ljfHhtGv1d6LllzRzcMhlmFUPOTYgG4Q5n7oy1QN
NOjaN/TsLt5jqbv86PCzZcM3X8c5qKyiHC/6sfv9yFC9btmoGis3VHkvwvcitoMrKsnqOIck4n9r
nl7tmHJPo+OAzhJ3ZuK92gfIb49rwB02/FuJKOBU6bEJIH6aPDtj549lBE0L9tD5ua/yuBTHMHq+
THpXNpBPQ5mDFsSZLI8PrCfOmGd1Bz9lRnjc0ZV13mEFboSxpYQVzQHiuxaK+usIFaGINF5buWh9
dcCxBXVN+nwe8imsXurws9hs8qIQJEoGIZbFOThxUJy3R4e97V5PCB6l+mQ2C72wE+vhhtNS8EGt
WEHvZY9BxQ+UQ+P2bopE9O4Ae09m6pjzAHaJXUXJ6KKmmAYozcCR3QSDuCSjewcS7BNabOZBmmZ+
42vL1hbf8EaoPH6g4SuPdFqwuEsKCBwavGwf/v0P40dJCGBE7bSGiY/SflVHxEioaODqxZr7sSi4
toAE7S8BSDLNHFansUPCChIsZbVGA8yNoTKo/KiVGqYe0sLlE7mv/yayojccL4qpRO8SEgIpmWtS
PyMzGfQvh5v7L9wGFCiCX5OD8vb3G1Sj8HCEt+GiLwmIHZ4czTr9gFubbGuI+ZgRriUjcaqn625b
z6Sh7qmSugceQIz2lb9Hj4XIYD3/Jy14OpISej4qcK4m9UXenlaCY2MkVb6eg9lvBQfnJDyJNKAk
czDmDJvT8FySZSleWhr6YUVgqqpbv/sTYDfdbQ2iTc9F3wFZPQy3Q5llKWpE46/UQWycFtTRvGcK
FlPGQJFjtGuq/MzuLjdyBXYUsiDQtnsDWuXYsQG5Jf89ZaI7aADDuxwe28oMxJlSw/SzgFQvM5La
8kbYJcvD4VKhEMNwE3n+cFfkytlcsDWO17zWc8hqIytieYX38OvQ3Fcz3hlq4np9/sfpeZQRyzHw
3qA/m/XP3Ncum1+k8D203BdoUI40dNOB2nH/Mp7fE2Lt+KoaBB7SzYT5FqAvq8lzZJ1vLcOD8oBo
C6QFpSe/85tkwie4T4nkQ74Fms0xMxAvYyUBy3LN+zjO0aoXtpDw83RkxUCx5yQSnDF2hGZ6SaEg
ldYnZsayogduMVPZ4tUqr8sfP31ElgezTDuXD9YWfFYgjlQJ9qDpIWirVp8UB70MthuXgF8OWrUI
0ELo9yt2AmSPqLElRRXqSHJ7BLvNwCZYHBdP/NzSdL/e5An4C1rc4rIIWGvx+tRK/odNMHZ6PjpC
jnAH+B8o+BBGzyNpS90/vrzwg2AMaEJ7R60ZHkNKYARFcl6BuURyg+AjhHClGXJmqW4KBy8qiwsM
PLgm43WJB4TfWJ45Ffcsmi2XcfR2TQgJCrFxBaeQMRg/f9CWQEDR/gqbMW1rw8HEKIRAh86ids5E
pfGsTZQr/IEQlduokL/Nuvf0kPY9OphHqa9lg9yaT2+f3Skh/lhfJzOxorYcUA0XS5BTlPS6KNkg
Gyspt4dTtJcogWEG/YslfpZg98Dos/4wVV/NA90WIiz3CKaMm1vJIHpIoGoN+mXghxEJQsluxSJO
RCzI9VM0cbkPX/q5O5v4sxWuDhN2FsrTU1i1K33pZOn2YznpXolmRlsSa8SdJipjYww9v5rIlMob
/kXq1cj3dOKaqDkVLWr8xdWTBYyHtFKFwhZl8MfmlN4a6msXQOHhKdL8ugiTzNrNTTrACGLJx1HT
aYXSnsYTWerRkKgrz4hkPJ41cS9VGmzcerIav/lp3/PgQOc4RSX1H7ZRgd4g2vqDgl6gz2GsPylu
nr6Pacy+DtPa5BaZvqDUdn9QwfpLZnQmA4pIr44xjiwAaHrM49sV11xL0mFx3BjobbjFVxh6PC2t
8m4u6XPcKn0/Y5OZa6aVsQMKwo9+4eNRg1awXr2y6D39quuWlnLHvVQFnNp57e17x4nezel7geDS
Ccwn2RkpJEahQM3Gh8rTkFT3fAuYU5pqGwKtNOG+sF+8VMPgN38Tua1mbBfmr/cHi/cvJoPmglVm
LwVUoSsfD7plYA9NZGK6Twsbj3LrMe2DttLvA3SL9oqgEVHPdb0nXvAjE8HbUehe79gDaT7tDuHV
MNF6WKelspaM5D6m9G5mmujaveuI2JTn44VMHUNY8ITxre6iq3Hm7xZ8jlwJV8+vDJqvdQtOQIwj
2aEo5VIV+7GV2rqgstcmXgIT/geiddlihvr0lTU67oZxTHr4Tamcy3ORfu8ElZNEdNzeN0eyyTY4
3dtkoHVS0il/fRhUMFxmdY1G79rByOb7vP9tpm2y8bDk18flFR4vogmTjgahyoGR6kZncDqRG3Fe
s0NQ8Bv9EYVPl9K5Jn6kyhEnAqrQiklaDXZKmAp1K1PChmRYuTnw2iNsxAi8nhB5jnOnlKgesHLc
XXVEYf3ySHXOzygG9hkhcbJazrEUnHjhB/UYVYwL6GpYQ/oWUwPCrVoLJned8TNR2pXYgW4FiZd1
5Tl8RFX4VSODNC4LZ7DoB56bAAz8X7lzv2OLTrMxspPy6LvI9aPYsQBAzkKuE0eNTVBEgL8i4qaw
GDxAigUDFOxsF1NwDniGv1/hkPXgeNZdT3g/ix7+TH7gYLrsvzOGz9UPNkWNHRHelOu2HwOXjLK5
00vSKLOBr6zDyvge6pf7X3BsyDf+ebvoqEuUx7ZTt89oSyszqRJFYaR1RaCQwO9WLwPG2TyqCfYF
byPH7aurreQMAvcjdFqjjxvdFeiNMIzFJQ4h6rdt7oY1dzscD7fQUKwijBt/3Y73Z3Xni8ER5OnO
ZcIvIr0Zw41n2myG8Dd0nP2JxZk0sqbG93v4czi/e72IRlYPNcUyGwa4dXZE1BF6SNtiWFvTQubS
dqq3ek2xXbzBNcw0veCFjz870dLPZgtqQhrTGK0o+yFFqtVF6NsII7yrY62vsjI+Qlx9jwPQK0BQ
4iV1pzfykY9BRAslidH0PQeh90XxJ7DDn7aow/eXG5//m4Tj9owuHkoHrG034J7rvpz0mOL/5V+g
Bx/YV/dD+1O1WIrtH+CgxH4qKEXfybDAbkGSMfla+R35wEoNr0unfzwM+L8JCFQZtvW+NTZt9Qyq
qOQTF+w+gt5jcXRtODEpUZdOnarConXa6k3Hfek7bb3W7HWyA1J8HZc7y78w0mcl3f/b1C0p6868
vj3QRA6/TYYzrJSzfSOOc4tbT8GYtNacNAo+dVdCtbf4uPmVDXL2LbBwWkh7G0UcYblB23Gm70Y2
o1OgsMrZKBHcgR18y31gQAbZQUdtfBgPjKwB7Xwncz2lgBLGJZY2LKnjENFEkNo7XNalQrhofXV1
NK3onZ+qe5f4VcQzgt8nhW9Cb0ws01XY2F0a0Xrx95NoftDhj8umuhd0U86XeHaxR/ndd64uxIaJ
5rugSrSLtxH09ec8FTxw8jT09T+n1qkvotTB4laSd6V0v1zCenlq+rTBqe8YeS5pfSaudfxjtrwS
B25G/895Qtli/lYiLJmNssGFte86JofbkKOmd2aJ0KtRFKBwpdYzPGEB02ZS0RVpWgiMPuYUVO9a
50kc+Bq3l2IIPe/g4QEfheA+tC3OmRW6oLfb1UFsmsaZOUIBYq3ezoBwBxbqP8mlJRMbAAw7IHGV
+BZhm6wzijlmHTM5NP26zDoaCHeTFhUxeme4VyaBTFiWFBguunG1LK3/wkmmDfoLij34t+rrzKoL
JKtJgKwWODtj+mIDHOlZteItxCQeNnqX/albMEQEnZIt+ZHVuIETzWk23NPVUgIDRQs9vHczoDHV
ZHylgDOn3MSFNuFqiXj1jq2XGGZWT4Q5jOE8mLgWamGxBocWlKMeOVUKpiQOdO0lQak8c9kMb+NL
xud/pfvYOT3UgjVjzzNcgri34yII3LEzWxkqeLRO4uRz3b9Cm2Q9lW39Ef0o7V6RvdWEBKMBXgFN
j/ZEP4HrM9qTSfZdJF7W2gTfr+e4SfRBGVhxyVKswroOpkWX3fVjBHruryYmdYT5yrW08Z0x1Mr+
TA==
`pragma protect end_protected
