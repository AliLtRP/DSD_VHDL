// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:27 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NH77SUTKgE6WjYe2bRdnCuTLiXNV/OpTkybJIy0l/k4UnXNgklZyTqOD1pKrpTYQ
vaX56vlj+t7IM3PGcKEqcXZol1nt78ErwUQ1PvJDRwvAvBMb1wfj+9j7CvfhbWv9
gSrwTDiTuHK9w70VqmNVbb7pnsJUvZTLAtAGPEu3OOQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3504)
j1M62DVQXY4OWTzGvreESv9DVNnQr0peJs4xKlA4+6TCpS2XgOhydAo1NJDvtWeT
8BYqnks8W+jLDJT0Hr0wBq/uFwq87J8Y6t5L9x+ajwsvrhXhq/N7X6dVM4HcsgZ7
OoS3WS62HfjTUQopDarqOMc4ApMmSPMg23XvH0fF0Bcddyauv+ZMa1lHTYY4cqdl
upfFfMAyw+y5kwF8k6xBVqMciO0XnBpwyFiQH6MH5QcD5f4DlhiNXrmhejew1KEX
MHKUQ9n3HfM1pg9uQcpZiw2DDXfx4+JZQ8SHwzrXZvyjdHLdy0tv/3acQIj1pdvo
alDC/0THBwZZZGlZNfIQR2fXk5uAZyPIRjfzTuvYzmfNWhS+kHTH4ILXZy9Utvf+
9hmv/adZGhV2Xvv3Wkxu17Ql7t1WAAHHMuzvwrxiP1WRj9DeZ27Vw8i+8j6BMPfP
C8xulMp6JBW/TnOgtxx3cP7yS2mvkJzt65HiHECk0H2j+HJwOFHOXcAF5VBFqPaI
cOQeIbQPJejMM+ALbyQgOv18dCdBayP0zq7S3Oglhn8GrZl1YLH8nrj5DP5dM6Lk
qJlMMvso2MFAc6ILBWHUKkNk1DWXhf41ZLjeTAkDkComD6d0p/tuFxrXW7+esnjp
N6uHymXGq6lPWMlTlbCiUHYS+3PZ4RizkRIQAp3P0o3C/EmxE8ms4oqSRTZDDFyA
Hiz4xkfgjDqZc5g4sMBQPC1lIFrzpghnC6POsZj+EB9V5xWLZgRK+8FyXMPce4Qs
olectNufcObSabHzWlNDKDDFa2tny7poG+NuVPVUA+anJEvZl8zgajFEXDTXkb/d
7D2ExWZdCACCtp6e0bK2XbDkFM8PW2wer2OF79H36sbBvj8eNSCvXFfQTc4jXxyp
AZk+MUVTda6dvfp1Ho7uj/4PQ6PYD2LbnGvH1CpFZY6H8iHiBEIcBAUGxC1r/ndY
yZABFGTkWiN9LYCxUtQ/F7CmiWlPWOwwakVMIqHIaB2umiRJmfabO5vwaTojwf+F
d3byGy4thxrvBnw40Ofa3oJf1ULsdCqYv9iBJ09DKQfhHRtpv+PMV5Hq6Uk5V0S9
YWT5i5eTysYQ3SkahWr5prar30zWmtGe7YBBCPhdpz02pBlVOSYleyo6IXg7GL3Y
4L3ydDDnJm62rPEyeXtfWU18G9qVRTNbsynuntkIC64lH2Tx97KP3j0YE43Ei42r
Urm5n2i3FOWGvIsthDRRg3G7gsoeFUQyHYRZj/sicJvFtYDx+t9DT4zsiL13RptD
CfEkW1YSVEzoOxXKnkfCYWb94kUTz/0Dt8C024jiljK87AZHbHM4oTfrzYWcPn63
nKPlPRYpmCUnqwX393vSZwr4djNHoBi278OKD/ZyQSnfFEkXnjfSI7aOtNHcQEVd
mqNdgEYKMy65YCEQNNfcVAnY1qM2ZtgcRuT+9Tugo1kozSSyx8a1OAqwIIr+XhsZ
S5inXixU6Rf4KsnAnWL9uSYR00cv/XPX/zhoDnVv4YdodyzfQqLHTUiomiYEPrhL
M5cT+6DMXsLnEABEXsnTEVU2cMs1NIojvvOhgF9pNFq5/NBnm14rfcnFvmZupHzU
jfDwW5Ug5Uyzak2hS9u8DF5en2gyHFJNfWA+SebDOrPm3uksgui5fEqUIOHq5yOL
xRjL97VzyFEEgXyBdskYpd2usiUuy+v+232f5Ts9swYKNaYMl4+XE64UP32QtDpG
bD3wLisI9BDpYLaGKvLjN9ZwMkZKmcWL3z56MsbnSDsrt1Iu4w1+rqTAYrUhXcVX
7uG5961jo0oIU8MD859+ieRHTKUrUdhoflbt9goKo/Kk3ry2fnNddJhbDKoQY0uV
TLcDEdrl3woGSfT1Fp/7OeiYRy7cXCT4cnSgDD3dYuXRUcqELx9uDx5QCOfIT69/
tanvZ23ZqjzXgALxtKxzC5KoX4S/DiwlpBSky3mK1sUtEknKk4fj7f0oKtvr858D
4ABFtzgMII/1nCLZhyLDl37O2gwiZt+BRH6F1jivtgqLV6bX5KBCVhX8f+VcG93G
V3fkO4YRH2UPD/FDrB2fNTqAc8PP536HgUqvVKmGzxfvX6FDiifi1LT3/6yV669W
XCe+dZeLoGB7YwoOLcg7QzHWQT7cueA5wHa7C0ucsAEYWmyGNAZP2oarLDekq77W
tmqhtZ3DxlgEd5X0N7NSK9xg0+6melc9otRusdWtUA5aD6cZH7+FlcqvvbVCOYa5
v+1VhFk5RbI98Z9ibX2oL4AakTivri3G6No7FH1thVtB4DEaU/uaNA3xFsDN0F9n
H/QX+O+AhrQD5b/FuJkabE3J/JyO+YWabDiPwE4+05tJcsLkSnstRGrZvKRj7u2D
yUiRfEEIkxLtebySD9E1iA0gdqW1o/JHbOJa1nj+kdleHkCz6TGOEkXCPnLYRHk8
zQliCg98peCj8IYCcpSJbvSuMnX4KRn3ilFMIDr+272i+5fxC8zrt0+o5pOUfbZv
2ZgRI/RFfufh1HtwtCdWzCFbur6DAgu0Rf6yGq9BYh0ViFGfCjq/Ae2WHAmg+wg/
hFLmoONdwMlY08b7JdlOxE4ofkuvFzV+7Dmj/w8USJ77VIfvNQFXcd/a3HYKlpIP
ABlXaDpFRVRY04QSNGg11fUoSW1TMkKfjYNXDKx50zQ6ksi+rl3p1ffxQvQ6XoNb
RCDzSaYlyEIpqvLsv0M61401J88eJWYqy0T1Vrf+4RJya58XJQMRaCPCCXC+uRnT
tnT8Ny2ADseeURT8eKcdmANqMvL7mCp+zK+ROr1vwZR2IcXtUTufWUcq7AAtVyWS
1nUfA8t6RoUp9RlwxqHBfyUk3Bw4WcEgr5b3IK4+CA2YeEB5Q2NPgU+lIsybqLGK
eJWvVkC0UhZ8ZmO8H6tORsgfW38BlGz55wmqrj2otfa8RS1lc+0Bw7Lfpxkfn/z7
8Q0cBmiGjKGYxW3fLtEim8tnk/xjpcxRB6yGuuPph0nmh8e7heUWTrBDKr4lLua5
4PUr3gc672jaf8tZ+RceYkoo0Yo2vZ7U3wxRB0EsG7k6ndC9d/3B5ImUMjtStlSy
cMR+Ssq2jjyzJ4EFVoGLqLAX1Xwtn1KAx0LtR7797+k2I5kV4s/JdpGQtqdO9zpL
omsOr84zjZifoPMMrAVj7oVGzDF+e1l1iUR9MC8zVw2DA2SKitWcrcpKb2mYZiL+
GBwTsP6ERcouhPBOP+Fu8NxpRQ6nSx0KSlSRkuRNVQlY9dtKFi2Y6t54uWiT2HjF
abTDv7OaUSWxO/uIDY/YM3ELG1COsXtTezgRC5118cFqKy9yoZ0dtSS1FYdOKIgZ
MwaPI3R5MCV8Zow8f3p7IaUcTA1kf6NNOPRAsVcuFuZMD4HjbF+lFpbZXeFYg7TC
W8Yjtt5PFib47T5mjZYzrWZWwgk4WEWJzMXGt1yoA7UBZPUNdO/06CqeJHbrsV7f
EPBf0GIfYcZLBD+0tFCTQhP9uTicheIK5JffnmZp6Jk6a1HxnESrnZrO9XSZk4NR
vfry8J2q1H4O70HWn64lSHdMvEORTF2ysbJ9i3WpnPjrn6ZEunitajokbaM4SW5t
XxqsIClX1lafnQ4HgJq1ZdHBiSEC1GEqxJf39pzSXPCWzAoEveulVJ3n43Mpnzd1
goC41FZV38U2TWLVPsNmaZMf/j9iKLKthBw46NitYkEa7oNGkxQ15tVzSrkGlhrY
Hz470TlAnyZwgFy2FNy7L1IUhxFicZmfuG8Oemo25Ltl4NFN0UV9MvfUTv6ubtZP
OWedqb7yCSFi68eYS8k5yOXUjKzZNvkp51DmSpEaWoj5mqqESB8e5j+KluNPP/Jl
Plyems05T4qBe5zDXPZcsmuutaFqR0b7qDF9Arcl5h68lCo7FgVT0vasNtNWkpKK
Yx3eJeDNY9zrhXvfLJwbs/svTw9uCTX4aW+b5k46ibazKXYLt2ooN24hBskTylRz
FbII9oB7nn2q8kCX6rqESiewcdzUCIU0ipQivRUZ36byATZt9KRh+4eh2dgaux3Z
AeyQRy2kroBeNT2KweC20+K3LW+YlHnP39gSyyXpQmmVF4QumznWsSDs5v+KCGXF
a5Q0GMxpWzM1J3/YB7FqeWXI6SHiD47eJDNYxFvowuxj+m267/JHeLbCDvAvYSXS
LO6Wh5NrD80zeh8Bi0kRZ01Yt4sOHn1iK6nJdqVrw2P78DR1nHz3NSZi6MQPr2Lx
r3DfQRKWT7/xwk0UEQut41HsWWmsdciJysFBvhs9+ckPP7VtewvomM9Ip1M21ltN
pnMWn27HQAC4wYF9LfO1ya8M59a3kRqOQmmyEFzBV85zaGjR07gmS3na+DA2FYtk
z4bHJxIcoKl05cLLtZ3YwZ+Q86jJw89Wx4xvQ0kT59+RhHFe154luM9DmcOe/MIY
F3spS29BVW5vPp560h/TSjv+TUd6c3bfS/CO73LXHsL76m2nCOL5o8DKzIxl7ZWk
gczLGgllFYzTQ3dAfOnxO2mgG9RpLNO1UCxD6ngNxAHHleo/8F+CNmWweS5RWTwO
5ou7TqWYVqz+uSt5AroHNiOzkRnwNvxwr4dFTMlr2eYH+bEm3eUb4FWOrgNAQpTe
owtTYMPnhccg5eSgowxKUh4BXZjQgUuXwRXRqTJXwcACTRifHADV4QghaydhBFaK
`pragma protect end_protected
