// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mn1FsYziLxOSmDvSTlKtgoYHgBgpAoqF/9JmtOedog2Gw7XPPz3i18m/IVt9SgZS
zpdffOL9+gXEoJhdVWzkplfc2BJicL9gmgwRYDZNfp7n6Tpfl2gAPqbD4GICL4od
Wd+flDiISiseatwTiyiN868mzXKETRLUOEBl19bof1U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3360)
T9Oryyvoie+ibjLpoWO67imLxJENmhxS+nJj90Tv0yP17hRPT18Xu4EDgMk9tF83
kWLqDArrJLyk6+84AabkBCwr5ulyH50oF8NweOUb1q//KaBffSoF/ZFIIzimNSI3
tmJnaN9wjNu0HElB5Ct63c+zmI7KcJLtXMDUYD/atn1VpViJZCS/8SrU+RwG3l6/
lPNZivOoYCK0z1fYult8m9FUE0NcnfKtNkcnmjzMQn9ipb/TnnwxC00TDmZ9SmHc
1pQTDA52DW63kI7pEoou8LDLqL+AHVlg9pGzPi9x9JgJFsQASTP6c9FwjcwI/7+u
O85wGyDx0Vlwds/AzdQBIxYzQFEcz1INvIPm9Wg73VH18ow1zPiP/ztQyaLJzUHy
4wg/KFVH8Qf45x1OlMbDlH/+TSoHiGXNLshAw229J9gfV6v3ekHd1sWdwu1x70ZP
2PsSEgSJllOkPMTR1r4ZavzOTKXISFzps3ULinlolWFuOwfpLg4NJuKcCc1XfNqp
pyHLqd+ErCgWL5NlIsNlKLCWkxAFh7MLtJRG27jm2PAb3taPQHuXvOOKC+IOJVKJ
0hfkxGxWy4ZFagn1Kz+VVIz3ESnedKxTMQGZcBhAgulGa1I60YxUQ04NwVSSGpcS
N3pcyEMHcro7e5hwmEUjqiXmNi0TESwtCEFE7+6sCt+1iEqL6I50C4hcSAKYBZ6G
RvHS3KlXwEpFlnZr8BwHgard7VDz+pP+Si1vXNPam8EX0ToCNXeWKkF+tIH5kCly
GBabApelqYZ2coX4EgAe5z7XseS6fzhM8ystx+PVUOeh7zK/gaylTeVIMyQQidnI
/zRDkEEj6fhm0fcfWRNqrSfSOE+47KNSfHzxTs0pU8UGodjuNFo8wfDzAiJvOuMN
TiOlJae+yamR+mmNY5B3oIm6ZpddY1m6q7W9aRk/35lmM5KfQdjYM+hVurXU6VPw
ZjqZUejk4CsadAbslM2HmJlGiSSyH0PzIW5mBup+zSsUTLlCe6W5o/L6tYHtlYAr
Aeu2yTfFf20/+a68vTcG7TA3FbGZ4he/v5/agnSBljCxF1zx8fd7kbfyfLSWDFGI
8PYWMK59MqagG1azId96u0hFmUpC89nCxqqSaQq1JUW9Qc/WiatBEyE6LGNN+/MA
WXTW51tUhXc7cUBNkzR4LFl5mBVlydb7kAjjNLPYM2IiH9nMvs/YgSDlSq6qNt5V
toZNDlv1PlfAKqY9NIYaCdiXdpTTBVZziKE2uPK7dkLqyRJPr8R9xZy8LrtkDX4T
33t7QP5VX5hQAaMi179lrXU14+8b4Lbz6EkYiRzu87ybBqEG3c9gyPuqwArebAeo
6kZt/RS8TiezZyUJ5d3hJDCcJxPZoyjmYJuas7+ehZfVvtjLhIKK4DxxljoGIKmW
n/NVH3JTngoprc11xgTRpplmZbQN8u56+tZVRbgKqRW1wxRmgRDRuyT5aFlRjogV
9/sMSeh0rOYCC2wLB7cp+xBwkLrS9KiDDzt5ScOHsiyWL+qYqu1f0kV6OG6U1I9Q
CXXYFJpQty/ndf/7ezE6Rv1+sSM6vh1Eds7opXq+6Y17PVB6woQp1S3Wl5Jeg920
as2S2zZuKqEZ9Xf46wcmP7Yw7MfUnff44ONrJK7AciT9Dc9ex4u2rQVP20npBOG5
E0nfnR3JH/anu31xVTrH8ZY5oPt5zf78kqlWsLuRWzhV7aOiFPyNwRHRzdhDevIn
cWu5r/tQmXHT7jEw/sC5Q3fz9aKrrTLagVm2KYMNxjVxuz8FFy+sEzAAvdTQjqy8
TKwUCnLEa8HxvTPLcllia28OxDoR+s2Ozm0P7nq8LNO6xfpWnGlcbhQpcuZOPWh+
VmJgsUkrmv6/1k1A9c1rCvqjtlUN9s7FupspAeU0WNWwO8GEacR0bWWcJa70RZip
sgCqtzWB37Zx8sdh19sABen1MTaY96evKadkbABPePeLFi3Ig1/JNUPIdBHAMW1h
6v0By+x2A5yIs5YquuUm5MM4bPTN+RzAmClLh7Z9jMbEzWRAvjZSR59cnQLQa/I2
p0Sx5uXiqLkNdRHd/Ad2BkZnbfGOqxG+yE9AcvRW+FqQEatsJLafp4FGxU1vHqkI
kdHvx9c2G6t0hCQHyFsRpDad+/jw+COqWJG1riMt6xvW6T9LnRpBKXOkdad67Doe
rG9eSMhwqH1QIViJKWBMtIORRRXTAjqU9N8788UQv3qOHkI2BnOiT6p/JKQKuASo
hZCgjIjtgi8OMS+V6TuoQNDSa2it3EA5AUbBCS1zgVJTx0yHcO9Y02FfFblk16HD
NRaqMFF1TY9PLQVOBvdBsQ4NWOPYPGJxOac07jjjAlroNMy/oE7tyKU2NHoB1uBx
WQszcKd2h+Tf8paRaNitbOJ/2VYzIyZnxuZB/KlVRkYFtW4U8cExIPulzFYqxSMp
RyCJWQPMlAwddJ2GbXDzOl9f1Aclwv6soXNVoSDfeQk5ctsFxvNJc5KRxYPis29o
R23RTnd3xVwKVxxP+s2eH6tFiTFx6SUIBB0XG6/TCqH1Yx8csxWxkrjZa76cFWvA
cHVRqIg9ebFpwgTGMQAEUM8qmTkOuabL1VqEvpRUnc+m408MWAa1QEydGJSzEdI/
KTdKBcrhs99asXBmIu2vhTiYpUO2aSDhpGwJElTZBErptNwO3TGpl3AM/0nzIj9S
VcII3w98Fe+ahhyOWxTpzqlZjq45cAUlwzT4jmJNEprG1izCTMqAmpLwO652fqvJ
52YNPIStZtNYO1P2jEWY2Yo51d6qO6bsub0lKxdjtH+whjMAIU4XDszhKIJNhVbS
WqhUTRZ0Ms+aD6b2/HjU5WvizrCXluRRFvLKRPqalFWpxOxUbRB84nJyEctdFw+V
/wrBGc0zNlMo5o4qvM6MMR2jfcP3/nXEmm6D3RFzOl2weZdnocFsTVucEXQ9byki
dWonAM6LjxIlXJmphqRNxY+HUIVdnTcjJCr9a+VssvxzI3JnRR3tWKn5xXc2xR7d
HuqDY39Lmr4DGhdl5ac+Zr5Iz3+UeL3IGdjgvs1pd9Uk99bF2e+aMNG7bndfMe+m
iysjpAKpG4qU6rTF2QaE9Q4QK2L+vmYpROQli0IBy6zGbazTDIoPiGo4V3XkYYAx
l+vbjH3Tmd6MpUf34YNEfwcZkJeB1xQRuH3acX0ExDPOpAGZv1bqaO+6h7FXCaF+
H5LXeQgvjINBryVuKgnQ8E55hmhPLbq4QT0ajWwsRyRkHKDYYKTHJoRajsMtKZlF
s7UCNqQ8kOuAWJL6WJ1RrLsut5u90C4PE9vsDzL91vUSTi31J7K6Z9Jc1jf/v3gA
JHwtP2dtCmm2BR1RoT9IBbZAf1qnRbbUTKS0czGDGRyWQtIl7l0NoITzDSzrSqPO
jqsJqcxE4+mIm0cIUSp0p7rQCCTZW2tJBvX8ydtsY0VHahGyoAZTHzZMVJnMIX3m
442SiT0l1GglYXlFHYzW++1IwdH8ZqipVkbXLbHofhaRNaiPi2JzXkX6975+vJ0f
7BYxiPZBHOwkiuCdfDJRIk/W9kOJhpKMf+G7bp/5VfT9HAiHoBaEiU9Vj2E3awlV
HpFqoj8h+gxLfpjoEK8N6zCd2Bq7Q5E0QkMBRao75O1w07f4hqYHfKigonjsvAxl
s0IyoG4BKxz7YV8HViqMPJYjShB/tgU/tL48Hk9ubXg9QjLkSMYSkvurTQajryWt
8ojTjSMnXUGpy4Ie7Qik4EQ/BI5J44oWfLPWX4RSeMgUQ0U4tRD+BZJX5/rtHyy7
PTTCO0QB8sR7rL7co98tn+5vj+MTaJajWuRrUZnaPs4/OxMtwiU2SVhEbXpRgsp/
8Yg/OERwNPavsBtRbMBlpkN4AsUIBWA1idv6Ge61qgKT/Izb/ClLJ7RS+8X03L49
iJMfHu0b1MDx8wCCrgYgIFwzY+yYexU+AceF+EAJbAjXkhVRI/Fit9qZ8+TBKV/Q
icmxVav8ita8CaRHcb3aiA6+TCvKe2TQzGyJRDh3FbqoVNwJhW+78YXlXOA1OAnQ
wkmaBSIaUEP5Yo1GQuSsbI+is/WjgXU/kHuybhI9jK2ZifRbnsPDcdmAD2FuMvwK
bIpgJpU/7ld9O1VNDJfELEZt8xekpw8Zio98uOhix0TQJ7s3gwmP5Xq1ddmeOshG
LgfjXAC0LwJ+bKDWi+T8uiD3ZeCVlDj1j/FvfOgEJeI3amZfD0SUyEKrGkMO8Hq+
+8FerYY1gHUnC1kf+N1c4iRIWaAdRg3PibMbDyV9tbOrsdOpSfnlCln9l8QsRh7z
X40mXtO8QtzOVESrRQUBNja7qkEdCKlQX013eRt2PvLAD+TNUPiyZMeX0Lu8F2vs
XgYvpElI6lzXRyFp1kyUYJtxEaDg2sPK1DsDxWadGw6AykcnXm9XrYcyza4N3zcL
0HF6CP1CziWIcWDGyUljyaK5z9BPpOTcEFtUILpq13UC5d5EwZKh/bI2wq8QdTRE
`pragma protect end_protected
