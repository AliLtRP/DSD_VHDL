// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cM1T9J3PHi4AV8zBDLSX3wnISgxzNaNO8LpGkUpa6+lM3NLNUArDZufUS+SEavHu
ft61R90hyicr5FzNj4RmaR2i1JRC8SkWiw0YzBHv6SjDni/3yDbIh2jB+x9flyvm
qtF3IvSqo4tr+VgDPOLnecyOjbbvFOFE98DdhFBSONM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5824)
3bdZdg4oNbJGNKyzQs90WV4HyvVUFL1AX06ALg8kSpGArxnR3g2AeDJ7bfsopVjU
i4ybLRVhiZo04rSSaWiXxaWlwjmSRP+PQ7ZzfJ/YbDdgMxzqeb+1er57T0MGPXbw
7PIOcBL5DwUKjeGLjl30mBVF+cs113/ru9f67oup154pU6LyzodNp2lkvL986OZK
He+DPuipqqvcaZf0u6rtI6ZuTvdBse81/HdzCv2uWHAS6RBrpRZ5h8yS4clWZwwx
LgLUZgIM2uJxzgg18E6atRAlIHxR1uTMQPVPCbaHGluGMoLAh2qcC9ttYHbVChEE
WHZMhwP4xO6Pz+J22ERrLPaJHaHW0Vvz1KSgXUDIJLxKLhDuSn7/qudvPrqX3DlK
7/Yul6x4uX98rn+Eyj4cwm4pNY3DzjHm2imfxF3a7hFiU0SE4oLeLSwHu4GjNiDu
j/dTDQIVwHF23iINbW8N6rB4gE66hLyplZwFIqt2lGxumtzhxJRzTs9onnix0IfL
uii7Y1Xp4CvDE1Sy0+SQ4hvkn1lKQUTOk+A6nlSoxAQISBM568L+l+qV/Obo69qp
wFpAIlsj/4vgfb8OORT/zeKSrAReccpKT9sgIaC3BruO0WbQotXZZcgHRQw19Imz
6y0dYA8HzlYWjedhWhZYBzczamWlKTdmvFDNPkSj8rWFdwp8R5ocbyVipKT+S2UU
XTY3cnT6C57JMdHyk01r5sObo97P3jpzUBFLFuR3ESh8J8Uqy3Zl8B2awM3Bq62k
PpY3C9Tr/2s3ykfICCSUjUUDOrZt0IfnUqVGJYWN9tXjpSwOMf9akEcBmBsZKgAj
xaYyuRoqdQEO3GKV0v5y+s2eZbVbuP+KLB4cSNEvU9ZeDly+hAb2j5+Un3lHuA8J
TF6XBFYR7kqOdu4+sbpNXZeVUKVCXqewjiB8UAiq08j7mKxeUYzVpQhtAnnnakh8
lGnkpDwuzKMeJ5DToEyw4Y9ySYDsoz6XlYxOQP8x+25ZJ9b0V/3F1kW4iafwhAZd
eD+b/xehXjPIpynI0Vj1e6pIHv+nuN0dX0qmqQnxiKHxrbl1mn7LTrFt7XaniMj6
B0KOswveiYteFQyRNkCJBIZmj3jpIBdYkA9oF0UaM01IH46PFwPxifVP5KJk5bQ4
oDn1Uk70yLnAHglu9aHGcRiGUxOjZatDcWWXEjBMinhPp2qWqBdBMMpbwMiGijJ/
ouP9/Bi+TUlcDWmUIr7649GEFusR1yMf+5H/Q7GmuR7F6AEV8CnhqiY+wh9vX1TK
wVhG/6yuKM9Tawlx1jdfT4X75+BDe/P+LAhso18/XsKKetdQRgvIiiIK9iUPf4Jv
1eSL3fE5v0jyexJAuEMQl/KCjhffWTFPicQUGKeJbdpFsDEXF9oYIQzRezUJug0h
8VTpYM16M1LfpH+wCa4YjqWyyMneSKC6wHWFdmuRQlTN6louEw6nPe24YSgmXgzx
7LbpgY6saRyWXu+oWLbuicFmk2n7j43mwpO4HYhKh39qY7lEJ3EYQWKm820H8XMb
deeI2KM9Ptpq4orbNbKF4E5Nl5UqLER/nkuky7NIqR8NUlEqzSax1c6o9YGqteUj
CLpT1YhkdTE//SdjmVd2xnW2fk2rEE6tKm67UzlOm9GnL/TG7/VCrxz5eP9PiJ74
abLwepPPn6tzpKjMX793DCefdlg+2vjRwpHGKsm4sS+S0WyJZUoY+Zls8rOYHkUe
iZDFrb+303ArW8KnjfhZbK5pS3k+yyTSz931DmntsgoSYL3ClqccglJRo4nHxiT7
MLmNIgmADR4ZAnonpRbgQ4TyA3g4toR7Qy5lzEVSDk3lx2PnSpCUvBZ6tjuuLxDm
+fyIUAK2PNhUxcrw1N6iFXNLpjylNmYifWplw73VYgpLmXi5Sv5YKiB2pdSc9Kzt
jaGN4+e8M79NeZwYkd1AskUNMy8ltZgxsh0grUTEmRrUdShSwD1kZLVSFjRWm3uf
kRMsCGCaR1up8jghLirS/8odSUPqYeca+EeYXrSkgpTdq0NB+moDt62+3Y8ZCsnb
oPg1MzEG6/f0VgJ8MF5rFIERzJnZnpzo8cLdvzfrfOTFwy8hhFyKAFWCfc+AO5eA
oSXmnVbPKg2yf+w3i7yAA+YRpmFkjdxClfsvrQvXZz8fkLiNo0hh6u57jwMfsNHG
pA9aAUyq4fHOrxTnkMFasd4+517E7+9jP6gIQDVDcg5uM3+5+TYVlQ58rF3tu1Vw
X2VnlFMPMJVUOSDE+cghMH/HkvpKAzzITj3G36U4m9z3TCnffJc2C+yFrKl+o6hi
Exn5KtAZz/02Wxc4YU6NfX5nA/rGfTWmdGSkeJ7nSG3JPE7DuSv8GfL0ntvqB7i3
JAScgLTV4fdl3zerDp9YjHShk2ZqYjPanr7ceL3Wc7W3Vx+sF9ldL//j4V20zLQW
qFQ4ZqoxKfgY5WzK66/phn59aZFvqVc3ou5GsGVJuvlCoMMP1tT2gDBkh+IJK+BW
DnTF3zrNi0MBr4cthpYBkuyAOraRY9KsKI/lEzRsnF0YI8fhyYVq9Yo/jIDW5bbN
Wb6h/020ZYnrTQeuAKJKNBr1XID8aelm3v/C7C5OtY6keoaLhomK8RHTlUWDikC6
YWIMstBpjgmEssQ9WjdvRyuwxhJqcYVEbRQYcowMG4vhkGsZ3HOk0tw0nsr92fhI
GG7MBR/gXHzrmuxwhiQbGgr1AO7J0gxihYlOTRLpjS8ObBbkHDOyw42Z80nFbrCD
8Z7bGhkTnW0FhibY+idQJf7SS7EhcS6WHhov4O5hKcIQXLQXKRW+EYmclOVUylix
C3t+aaMb790g5RsowZTVcm9ucykrSb4azvEfLSUMbGugNZ4NpNkJxCeYm5k+eDhj
S9qQ2JJLAiP8qvm9fSo7cdA0AWlOWXaImVIPt2BI5MSH/Q6LHqJTogUca8Ksoxsl
2lqr/ksvZiNcuYVzpxIBXJLhuawqIKhyOBn0eddjHCIqn7DL2bmUiiWDMT4xfNv8
cg+Y8aiRLsROAgGaPuGFTqcxVXHoS3NRZPJj1e3my7A35K7P53lqn0eTBP+yYV5Y
UMbeDg3wZspKUYU5mZLeiK688nnB9FJjgMVHOUTxRIJVtArXsY8GXPMSquKC95MW
Ia832THQb6Hu2oL8jj6Ch+ffYfGQ/kWpRogA55gtoeC+PgA9vD1FqyTmYkVo8h4V
m2mrpm6GS9uyE0D4cZSOx4oJJVQdwF5IOzWLcx1en/O1XyakVBEuCIrq45ssa2LD
V3uAonQfzVv/F6LHLXmWsXScxJMQFuFSa4H7RVZJhtj/JVBgGMjgjCYACw3GMKsW
lHd4yMt7eB7kKKrIb8qybfS7UjK/1cM9cxuqpj15gVBZ2meHcSSXnvcT1Q7T0yrJ
Dxfk9S/rpEYJ3ZbqNJZA3shfHuMq4qcisfREeaQlGeSf/peM4LdllEiz3huFrLQj
THa+RZ3aGE1CSwT4DFeg1j6x0NhHCqiEnQ1bg1F+UWNcK2hkeVftSiDQxhNvDnui
PtUwWCz+bGpGwUbtFYEEQGNisZhCC1zmR6FaCHisylAD6L0zau1wsdB/qnjSNgs4
5GDegAebnv3wKs8eYvCVTVwgqEvVgCpoOu7vAcVVMYJISCMpYOi3Lj6NKmSsjzcC
uKybJRLF0jUyZo9VbSWg/FADv/ltpjtB6s8BcQpv79YDByxwsPz7oHsEb/GLYK6E
3ZScExUqTwaTcwwDne15GqdFdEPf8ZDPPNmZB4gRErRbfUeL0l0XMrhlhSVWCoy4
UGBYGPRkJ0hfQkO8ln6xAD3LS/V4qWOba/JRxaaM+d0LTwkNYVuPIUItx1U/+KkA
50t+eW0R1izhTtzL5bFCkUJ5xL4OMlEZDqc9TpJtuxpETrr0563CakRLDYrvTz/e
d7MKEuRML+L6XrvGf0UyMdyFV0437JRa+MFltCNdamKn3yr0dB4LnTHOn7LYA4uU
OqRuuzO4/PcQKa8d/rh9iYRYL5lgoz6pbex3xDDQsHPK/L8KoVyqlzAYNKIyMKpm
ZnRRciYQ5+gKTA3Fi/tW5gG6x3OxnPkrHUjw4uBra/Npv1L2jS9flQnfBdHFJGuL
NN3OuhzpiOeDaaqTSO302a0HbeC9G2n69gkeUEMqSSyxC2WSmHX8GCzwZ7yOgiv2
44R9vwV9VX5CFnlPzwdsNDgoxiDiBx8OKnU+Gwf+zzVCoaU9h6fPNuEYxSHoodcU
j6vqB79MX29QcP5Um7lyNvv9y5vCFQo4WU+Lk2jE0D8JlmodGZp4YZsygvHIzxSf
LIPfg1epukg70L2C4HfAk9kdqkPw5c/Nnfbyz31u0WUo4oy58bwETunGYVlulCJr
hsgUiJo+RQpVb2tzcAUXxLjH3o9kI3Be8rSTm/0cWqyHGM+Zz9qmOP0un3uP0rGA
rd4dqvvWIaw+6+YfFA3fXXk5bQtmiLT1/7JGZvHAKbs6v5gLfgGwpR5kaHDeZ71P
5SaiejH5tfYl8lsjwDUBbbos0cnYqxdyB9fpjb/7VpobnSmeQxzB8Y95bSSUEuzQ
UltgoFvQiUUggmg5XTXNlrvesE8an8X/kRIsRX4laSYsKRwvUY4W+Fuf/lsUra6D
JizGeEbVOldTP8k3Y2XAaAg6y7E1WvhtU6BA6o1tbQCAgeqWaqlXei3RoSEulIT3
+Y46/9wAvkd2zN3jfZutaezQfxc49HU9E5MocgJGWyDiubW8PoNzQgJ2K7BEl24x
9FIU0Bkdz0+sIij6N7YoZGdWiSmjO0YxDvkR+3PzAFVWe5GuSXKTzIyMj7SJM2qH
5qBQFS2lEULqU3wG583vJ1yoRX8r1ZEOsUGUjfvtarW6GalRak6decOvA8xdkxdI
c3+lSvC95IJhFWQ2AGgq3lcJQSJ9lYffmJl7T4m5Tp4Mg5ttReRPOFoRUlQC1RYn
iBIVQ66CKXU1fMhIFEcp7LENUVowI1711zMrxNaEUJ9dWsegW0U7/dT26SZ0LiGE
H9IAmSef5eJzfvcB3Fzl7lrO7mgwkT3DbCdAlm41uK8ZB14weB/p5pJK7gf/sOte
tQGtjaxUlFUhOH+0QZB7eUDQAsrY6If5+FoZONzUBM0NX9HknptypsYNLC6juK26
wVmvu2bIr+XPIlSeokqL6nQZs40QnLh8a5lbG6sxqxpdwgj9Z1xBenFsZNcCgwcY
E5Fvopsn/5Dy68vLJo0ooD0+7iyZsPDUP1N/ISMS4/v6OclCQEHi/8t7zdutT0c/
QJq0fL3GSRSC9gHP0eJ5/a5WAcCtRNXZHCbm6vlNN1HPMgHH5esmSw8WV6RaIbpg
1nIG2o5D5Z4ZUgRkuQRycawyBuzp4TRIq2a2zKT6RJPnXavWTV3vp6+pIvssezvD
YzN0CT1FbwA3IfJFLcYxKoRJnrGnvMVy4JqG1byZyAF6VD0CtxQhKfWpQ6nvCrk+
SiupCC6I2+p5xKEMwDb/LnWHJhp4UGyvPWeV/IEZFXdU5qko8WILPsvsGlZzUcbD
s2NvIpNH1H0y2j+HYfaISFM58mU7voG4/S6reBdzW7aJKgA9tDHLUSBTbNh5ez8e
A4Qg++Rqa1rU6j27VFKg+Ub7Pmt4qb/WojS3Y5/vS16bRAI2vSNCKtCnENYsKLdE
wV9ePzKuWAEKLKoRi0JaUpkWvDIR0eyM4FqpfAWi+v5n0pXnLy9FO2iZwj2fhFEM
e8JihwEGrRuhjzeJaTDtwFEEnqDXUjdwCiWrgtY4/WnKK0ieGSfaoDvviXrBIUx8
kHB8EqwIRsT+vBvPY5E9Pw44UpaE1+nS93XUu8iC9hljr2FWpzr+VNxM0Q866iwg
ncPh1bSwXAF4vSCyH0DqPXDBfAJZ3UcBt0zCaLvz8hJKVhmrpFfF/pvw9c514x0P
xJpsK6BrWqtFgrl8lgbTUZovBLVYvp3JpwDQvZn7mC3lyGrNWgeFHFZW6TTx2K0B
GsGGR45y/6fQ3egJTLwZrKqiXxwdnU5ubq6WVuHueiD8VOx0+EpDgZOE4BlRHaAO
irMwIVHaNtVrMDqvFpBaSgkDTnToVWPywu8kMQM/ocJ9cGcljyeRazfLGZOz5D1D
URJydJzWlGnhrk2fT0WF4lm588WCjDzr38c9t/GF7PIVbctFG9Vzo1ZsWfY/GGgZ
slinVzNqHh0GKrZ1Kn9Ff+axxCgjSFK5flxWb7gI4Xrmmj0GzlkzskGBQ73rtdV4
IFo0E3VodZcjqx62lMOk6JIpVEspaor4x2t30DNRFso7zficMn6y1e/AgaPz3gB+
87tVXig+ieWb1efOeWfmtYaJphxG5IbruauaX7nkHrcfdpl23Wc9ZVIctGDe1eUm
gwk3DR+qTp/n+mCd6CJIj7UYg9FL8Y5rIQGGtD5b9LCs0IdfV+SVG8Z6tlauAova
F5FxjOMcvYomaGpvtIuST3nLhO7ejoiwfuLkYz2z8fdeVKxTcpTsGLrBxNmdumu1
gwLEc0ex8QaRzYYhss7QhhlR5NBC4nWD4fRalLYtgeIcH7JgkCgnR2zGJar3y3JF
nFjcvA2KSTSVRzYxF1SVvtVghtNUGVK6ZpYIfQkWpaFo/haGPxl7fkN+69FLoal9
upIZjvy5Qq5n0kFvQMrlC8ZHTn0Z+tnU8I7y/0SryDj8/+9yOAinI+tCjm3+/wva
OWB/CTtusihoPFQi3uhr2zoJGeXy4OCJ8GMumMYbTdTMBf3XMK/dw4CsfW0L8/CM
ezn42tAi5IqllZE7kNk3ViXg8kKdSxu9jljspE4bjjZl55nr9QhTxxeRT6XnkU+x
fQQxuIvLiS0kk9SmMLmka9AsN0kCbwUqVzaS9FAVuXZI0dsoOpP9KJsPYHcs1n2G
CROcONzx/ZFxuWAr6QkuJaSVq0LQUS5dRVoaaaV5j199WNRzMbZLyUdvQ9a7qrKP
CdBNqsKWk/kZlhEuk/3SaxBpl2VuKDxOCD3YuNTq03nhJUZYK8dao/qqmJssJiYI
6P3T2uZWy2JBzaUZP+TbhaxsQneQPnwaPF4lb0mp7LviHSeGpyor6BMg8KTzv8dm
jLTHg+H7Zy/3RTHz7eN4RKkQ+Me61jgyTJzx+IFMkuIBLY8+YI/Tt5zojXTAv9FO
qvWl+lwQq64Bf7FV8jQtQ+yAsXVjI0/aJWxli97TWvhkczc6caNn5JSMxI3x1/mu
z8qYrMSLfy6rdzgZrLtrXQCq2t9vdxZZIndSsbATmQ/hlasUeV0pIM0YvbSybCWq
zrcyy0uhdOsgiUqnnsXxhvkGLzzegnYP6KrN8siLxUJpd8iemOcZpAD5+HYgry1a
5HVGWcXRwjvj0iGhclQFdr3Cx+DG+cK9E4s6De56PWX4MMaWyxAtTJVL+QktYFM3
54iJeDfQHqxV7ikUOVmUJngWeke6s77se5FrH7RoIoqZQCLjKYx9fT2LouNMVSAw
aNHwaudPkblAG6o0Fmf4Te07WWExqXLEHoCizVvuKEz0JIzLRyiVrYUmF5MxkpXQ
YZdavzKhRLx6MjkEiwDlLC9oMdeg0Ek7Vkt5N0hwQBaaTGbESN9oa4LJHHLtsrP3
Bi0jmPtQ5aBTvEszjL+8zcw2wxRQsopESthGjdtpJlGkP2NkOUcnyyNjBIte2jnL
I8bcx9WEk18QVO4KVXHstl3e46SWM648pkAc7DRaI53YnPTye2gPVMXn+ZXHm+xS
QAElMrJJduCZYCrCF7nI/jsNChhe5OHScczBiWtWbALq1kflI3xvFRH6XO8guaha
D2DwRuNt5A9VbAxAF1/uhA==
`pragma protect end_protected
