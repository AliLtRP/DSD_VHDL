// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
mXt1PX2tOGrdmaLQlqYniaLChi5NK/EkombzQhgIf03rgchkCQBcXD+9ZotVNqttx/5ZwwgDdeJM
POfSFL9LnQoF4El3Zu/sIlFs9Loe5mdgntL+ogM2JAzb5rj9sugc4XkciL2L2d2FBBUq7P+Vgbmz
hUXuU0d8NdKKoqPK37iDUZAL1a2aP3ahYsVl4sg6dsCoXzFO87YakIrBEWtHNp6t/oJa9GJkyVmZ
fGbqjovswLKuXB8OiARCm/6FXMpNyMrSzl1SbcctTCB18hePW9zCgcA2q5pvPZvdYsAkZX7/PVLS
PC5dKGY85Ona4jN7TMV+GgOm9XlUZt/jJ9xi4Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
IRH6EC/SswkzWftkQ2cIP7Q0Me10Vu9ch6DE7ZRpT0/kyYLFIlgdbs1tKBMe3HJWCbeULmKTYzWU
LUUa7J/I7C8G9s7Kao2vF9UPIRgNTOBZO3EUW4I6SU3ja7W02cxyjCfta+f7rsqA/hb9idk5pu42
YE9Q+GF13tpT0792jObFTnRfEbNcqDWS2vTyRKX0kwQh+D36vgpurLZhEywmfqDzVEzwgQ/n+yhI
1FLyV9k2xgx6GYazk2KD77Lv2ygxldfUvEWYklp+NbE8Pys2C7H0jnYNljQFRJF+8pTyaNdwIbc4
09s/WkNSJkOyhnajyXNFKaNzAI4Bf9n7MZF8Kth2EG+L5yeQx+lsOAClD5cLm4wmrH5eFUOE3ecy
WS2c3Nzh1Lq/SO0bQxUvUFvIqxPJfCGsvQFKcPna8CDcpPTxzCmXxJSpjKKVUZ/ghxey2a0JMfNq
MP+b3jHUqd22EhR8+hUOw6z2Nb550KJP01sldV1iqSb997RODzYo41RP3EO5eFPp2wZkJtzdnSu/
BC47y/+fCcSO1oCJ4p8E+a/a4B+a48tWU4W9vkQL97aifKOKgduAvk7PXnL4yNZBEINR7/H6EvFj
u0OrOvyObm4lpnytwxfYqMUqR8LKyR82+4rcSywR6bzoyaBt4LeYGcybjoK1rK1wEpGj6BR7+jfw
P7GJyX5ZmSe6XZEREUSjJtde25AWdEgWNdWQWOMzIYQyWXXjhpoTBwe8QF/PKLI6jHBd4ce5usYl
ZYbFHP8y1Mt8I8poMSGYBVxmUi2rlOfKUuHohI8nvmYzR5ifkahL7/8sRaCGj2uNOdmR4Qp6IiTT
JoquAi/G9t7OW9AJUfAcGNI4KtXlKsL2Per1ttb+PEC9aYnuVzUtTTw/cbzFQ+OdLXRPcHTs0Jft
EFhM+M/2wyLff7+bMuZLPGWvTJTKBjQL7sjkUOjBuQ199YCe1AKWYSD5h4ZYzZl6ZVshsOcXpDPu
6MQindcI1w39ZqoE/VtGB73W0a+YS3yPuarS3RpIEs4w8dY5l/Hzi6aOvKWQC99WtfSTgIyGtofm
6DtxOWS8PXMqgtzDE229O53EqQDvSfMr4oecFmMEqdnIGofINcBIRlVQ+QDr4ZaBjHi/M+0LLD63
mbl9kfw0ykBW8izzXxgKhj5br+/o07o3yIAQkqSMpAs1WzForiIlY+f5AcG1X3vkejAR7jOxYP9L
kc2uS0/emeuW5TCjka+c0P+zplRxKKfooQ6AdLAW3oi52mYgMn7elF96CmW1201CZ0ZUJHB2p6fh
EFjOPF7l5P18LUK7hpjJUmXE0Sf2Ezl2GzD44Lvor5hBVq8eX5ZIGRKhgyWGTwp3f7DSZKl42wVl
HToGBVbR6GIn1WJE/Md6SIq0nPfkoQF1o7zcg9+QkS4HQ2s9nsz+3LJ7a96ovkwXELlz5XQ68NwJ
3mxf0TUftodV2wOwaBhwqkklwJxJ8uiXSLuISvKtI8FqU6Odb/DRzZOU1PuDbFgiAPTEAlcIEOkp
XV1VgaZRh/icbgp1pzDAV/EBlvnJoA8HKrwz4f0aV0zvlKvjIdVNnluRmmY+qJd6JQr/IzBNSFuX
nr9702n55nUjJSmShPToQje1+EDCQyaqmHojoaB+tkemSffBaVN+Edpzw+AWlwFVQnJmSW9NLo/9
LKT98pfsAtQ+TBT2gaQOXZ4MT/acWaOriypjHXHHp5rnOunJmzpe1dxe6NvEkeweign2y0dEAbaM
iyd3IjUOYmscW5eML9OYLk7hnsZVNGN0GpJzjN+on0MvHvlfuBCTqhxoL3218SDhXMZ0FwKtpAGg
3Vptu4PbcpUHmq4dyffcNMUNeM/CUvCJqUKD6BzEuWFoH34HTzAGsUcJ6MrJxH8w+Q2ecRUc55TL
ubZgBXyjzTkLkk2rp68vA/WLY8qVc0SvNUmQKlbBuYH+C5HicYT9t+ey3ilFov1bBZqqU6dlVHYA
HxdLxWLEcpQNrRjGhtDGJBTziRo77SOhsrf0Oj4AvffH8udH/KbS+GFsBDfbVIylK1aesgikZ90a
f2QaOagwIWirbudw7rbaUeehMd9oTvZmrOFShsovj2wJ63Qgfadp7KB5SLLyJVkZ4m2evFt8rzOY
+rT+1s+CLoBzzWQEqlLU7kfxmeWtrjnyNEILUCB3IuGuTsfe7iLMDTqtYPqkBL4auU01N12lRp3i
PcQP7pbtJ7fKuLDRBdtQIVpn/TXZtXEU2GZmqOCA6IdbPOIEDJKzL1RaLX40dFUhTbbuE20LeYPB
DYRLbPKUoelgX2ODlZC8s2Qk4706UqBODtZm3rzBRQZPcptIRYxdif87CbzXR1PMGkTPId8dMPAQ
BXH8oosN1Jumyw7lKPsg2NeSz4K7jtvVW4T3s260/e1Dbcv3cFICeprwwRqn7cYX59zi0Z1TvAgn
BEa+MSjQDJCeuZwKH1XDh0lHZyFnw+Hs3aYK7ltTVyJgsD5nYzewvaW+G4vsveGcRL75YbUzRo7O
wYtQ4rPvQFoBzd/L+dYTA1yPK1Ec9hK7j9ADvxWO0+yfxXqDC1L5CdmM7JSH6jmQ7MiU14hBBepH
HTuu85vkVRilo51/T7X6denamjr+/1O4qCVbL7xNa2cWndpKCzEUv+pDBpsoWLVcPYwLEM9TCbP+
J095dgHvDWmmEspU5x4QF6UFeQZo98e84ICD59wQFq2+MosEgjIHnSzlw5v4H7eAfiVNnLAyD68k
jPZIKTU0z/n/2TiH1dvXeA9XhAlgLwnjVnSaa9/PUf/rbjnWAAPBIYNzkbay2kDez5Qp/uiehRro
A0VWAFQqWzJIWS79wI6Ws9QaLhgVc9QO5n3In0b7apdr03zTmuMwnS4XVqMZIe26kRdcULo9lxte
DhhpX5nCd4MNlEhar+yUYyGUSVKyN37L36XRyI8lZka5f3XvV36abYoBYjkkSOsXdhtENUc7Uld9
w7W2NyxSdpCKEJhnkV6JijeWOnBGsJmkGLDiahhwcQANXsp5ZRjotXIHpDR23N7XC7VFGFOO4dW3
0yRlMZu296k66FNVtNcSJxcnm2zff+S3gwRy4pqCXczDIvpmn0d2k0eJIBEXbW0LT/yuHSAM382j
ZN5NqeqjYoDNIXlvsHocUI8RUZB1Zi5XzsY5ZhPTfMC2sXVGJBWvRMjHSW2vQYcoCfjoumVfknoy
pBPUgZ9TTQ2ocXx0Mflqyz6+A602kRnlVaw5Jnnd9vK4OikApcgvExWO+rosVPTRQU79/v29CGxH
qkfbtVo72JXq4r3M8zq4nR+62okvCYvKMJBIBeVge2ViCYPRU4NmNQxtl31FMhf1jc9E/HFl/bRT
0PFROHtAhKK+FViDlri2m+ClSDRQy09sWGT2L/iB11bogCt/s4z4ASKkSOKyP2TeJzeJcmu75/7B
UtWB/h+7RKlEGSvbx59qkX7piDud/CQadMVq0kzO+E5zPNJToI/9ywopUP6pji6W6M3QNXuAuTek
ex6rMEjkj8j7tuf3xVQ+mzJyHRgYfNqhXBsgxoEKK5HMIsFflLxjjzTkzah5HUF8211NZFz6mb3v
RFWAe9fIQpsD6T442gaK8l9cx6num65HNg9NzqHEDqsrHeRYtbma0pJasvlc6ceR9Z1USljea6pB
Rth8/ZzSwSbmex9Nbot1aW/VJ+ZUabcTy4gvAdizx7m373aapj7HE669MV1sjDVi1q9n7qUEl3yR
1a4XYrtuE5jpyj2s1dIBzPU2Eznk5OrJtAVjzd9j/DufHwTQ8IwpQNyVk3imX4zj5rMI+1Zmu+TG
gFwkPsbaEgBO6QREcVGzLy+H6RHlKa8CrB+eKwoOClM39uf/KpVmGhdp6GIu08NhBvG2vyq6W8ZX
ri5XyoZyY7j0JEwbloprNTQpcT3Gp2y5HcPxTu1djVEsREuCSFtfFmTp8JtchGs8WGG5aUWRByJQ
IBJA60p1nQtxlFA9V+v/SFl+ltwmetaFdHTM5TGLUwVSP0cNSc5xrC8+mIKKmQmSmq8z5fbVSENN
yp2awJID7R/tzyeaVLGGdiXdSrLjdG11GMLuf14yp8Igd+ZHLZd1hQnJRCdKHp22vY3DCOG9Lfe6
x3fDjtWDqYrSILQoN7w34aZxFUm4lLSJV66Bs/xannfbgEEhLFJrik/Hd3A+nrVxgWmYvPr0EuhS
UkVI09jcL/VkHAFzwUk7dndCl804+ckbjOAPs3U7pbEqqf2jL+ZOgTHHLzCfCtwLnJCqzjQVJ3p2
GdmAdPFCzIW7qlBoFS5y5JHpoUXDYBn7StY2DwopkNhbiLdZHt0NmVTMQ+89jqF22DWpixIhNJNU
5QWJcCM3oHMcpZ4pQ3PDg6Dly3LLS5my/rn7/IXtknvPVocTBEQHGbtF7MxB0SofVny0aXxuWM65
R4jdk2zckFE/nzz3jB9aUWg4F+SKlXqMdwCDotbAV8x/HHDQC348pwR4liOnGJsT/ZC/tx+b15FB
V08tpk2+LcY2kfAMbWsLLG4w95MzIwguEOdS8XLRIaH/qCjo4RuYmA4VunB89S49yAfq9qbWCHGv
yOqvAQl7L3bvOWj7CeqW3+x9kFYAbcHkPdKIiTIwrhKyHvAld1hwZ7tOF+1uodpcKEVQCKvjvo9+
EdfTLRo2k7cSQZrceCUZ/g8V5pFwoKrOBuDcLDFtQE/CNbxeJdlWG9Xuf4slphGvTp1ZfaDRe1Fx
+A1MuZ8P6ZkOMozKnBPg90WoHbV1q6ctj35oRtKVtD3ClgwbmMWnP9fS6bumsbdlXraxeLGp3lPY
Rwflbr1mvOeysUU35LUeBUDC7nc3MkVxl+5ySyTuZOK7qQQXQsNFz4fXVbsupl9IRhjwtp44wMtt
Si2VWpGX+rGW+FvdKWDgHs+MH5J2Cgx4GiNpliTNDk2SarNZ2yNYGATNPNmX3ycKIKJP+hHF4XoR
isRf2xHlgQrfvU7lxriwlA3hhXQfrKaEl5UO6Q8+ckemR8A2B3pY/1U09AGnQeFllzKecmF7QIwU
59Eqkp5taWYXBZT0TFYO404j7aipuSkxqoY+3ceoYSPCKHP8084tZRsQyDEMpI91sT+suL/NDbeP
kx6BK7XcVFbbWFZkiasWXi/HVCkMUQEa9PO9ucC3BsduZMEIex9cr/c4KXchh3xKLrTUilHLfvGv
euDNmhA84ob18RDbYqJVz4oAZMPWnv56qAmblEtC88cxiYj+wP3EpZ6Dlzqt0pBcs33oK1z7vtST
q9L3PF4uIYrZPWuvODMn8LzIixt37nf+mVkFLVc2Z5hUdOT/NSQYCnLgxdcPvYL1yw0kGxMNi5HW
7USFZOTDcU39OOnZEtZ0GY3UxiK4PNSjzmLdWX7mtSAJoi+4GMHkNiUF8M5EurvJS8x546Xx1sqR
ARTrdAWifqTgpg2UBOqm6QYNAKX0XqrGQVBrsg8K5SEJG5fS8oN+uUzTPOraphd1wrf1jcniSr7y
l/em4ezZXiY/NfdwaRAHmhZP3KbVqADvLFZZVcGmMTz51HeO39ZrD1Z1vR8a/hTx/OIcxneVE/vn
QE5sSV6JHDEp/FbbDQ8NwlS9e8H3+pWFzvW5VM8JqlXZkNHGtRPo83mJUiwbvW/cWnioFQzDmsAt
rh228bsIq6JfzhU8QPhCvcJL07J35bGNAM9PYZ/I/rdjoeBWJCZhY6UCY75Nf36vZDW26H2barNU
SJxDp63jX/3S0Hko4ACZt3mMeG9q+wEG4oYHUcX5OSwkLTwDsVKxayUAtt0AG9ET/zYf5SfeNhMX
wydraNaZ2WkOkof0lDfb0AvKuA92j4Lwgc/mJ0itbNoVUKWpBe6tnN5psqR+JJqSpV5zSaXN/yxt
3T+RBAYORGOUEMSKPvv4DHwNDjmONr4a7komP96JNNstUTT9kUxWG2OlX7t5xE7MrytisZaXUVrc
UtNPtibaMDy3gA11C4JhNY2e2oFyJbF+x29zbUFBcMpqM/5Sel+L09FUdZ0PUa5ouu0hnE2+VfjZ
H4yvY8Q9qy7bHFJxF6Pclm3Qb+TCP4GLoHSWapN5aojc8vaDXHXdi2/HY+hcqPKeFxuwDIlryWDw
15Xd3NK+LvIYOhf0vGFmBs8Dt2w+vxokT9cuZlnOja1MpsnzLFlkra5RnVxGFmyx+9Tcfs35rcx9
tcVYI00HP8+NirTFxQjU1O/kvDb6gUhHA7hlfSK0k8yUM1tb2MLDugv3RTp4mx8cVdWUsGncprNg
dzgY7QLc2/wODBvubFXK3EKETXbzYZuMIqhZWNB8FxGmnrRYKj7eZKi6gErc1d+pyBb5Y8xD0myx
it0eldxnhPy37BWyW/oreRK0IsB6H3HY+r9jcJ/W8CI+xrsciBRdNhWx4i7fpD+5qp/mci/Cs06T
e+YG2sIqCf2+pvS5sjCeCohM9HWhfq2MY7gj0gZmWhjkW5xipetdBGWAM2jjHs6PaNz4LnVGtggA
mif1fQGUmzRyuxuDWYTNnF0iEqRI1Yap0nf/SQIAGRyN/JK+w+/iQ4Vw3InYDkK2r7GOI+uq2MdE
ueSgN5Q3H0cOWYriax1WuRl0zxQR3GkLkMfhdaD+xAD0nZOWUfsRvNmYgBGCOmHJX0KioV3GsttA
9/W85bP8bqpVChLXgFyUVkTbSXYkN9JyNC7n/QwEyer+4zo3YJcwcJkcdYbr5C1ihno3NdDZU7MP
p+7B1x/DLmz8EfmnwOXfcF99VgJNpDT46Wdtlzrq0Y7Gu851wC/O+PpNcm0FTaaiO4hYBEJGhV/c
9yAzARjfYY8MLOHbZIlT0To4QlZknFgYUMWLP58KMXf5lAutP3lSIY5xylKEjysA9HjlvtyAJQP/
Zng6cI32GCrGLaFCTLrSjgZkOyFNY3AHIFTs8jr7DJwLHuWsJJ/9GRJqL1nJURcbHO+BNdfpO/sp
pdBttDNM4kgsuORQBn3qj45R17bjaELg4Gr3+ArrNFJ/uMyfb4DpGgesTqWdcbEHGTzwBEfxsnjg
qJF+mMi/HY6rRYCiOqhrmq0Hf6ualszUyrR1LYEVZCHpdIsz4RzDHmQWgEPdHlRyYfuTC02oS2Y9
Q1IYcsE5yRG6qtb9mZjY3EoKVFSIAnyT7IlPRlBwNHalco5jVJHSjKBWbKucTfxKDvMxFbVAL+rx
NsTMIJtWaFb6eHBnTdl5eFkBW/IQq77pOd99K9jpKmFEMkosCEK87XCM4w9Q8hgUMFwiscMZD6pG
2Mo/yu6Hr+P1OMU9KnXjkngf1/jU+i0OzCcw2jsJXSgxmYiIC5RIzW91eZZRjqb0vS2WDoohS63h
ICEAleZMIFnZ6R4ZmuztQBPljD9dYN1oEA5NlddKXxPhMNuQHFtI/X321IECfZkaO3h5cDK5GpWN
09nLD4omX1V/2t/4ZCr+Tf/brKdEBGT0VlZtVdBTii1k/NtfU/KQYMVEYuiHqcujkWw3nj2q4pHT
QZVUuyMRUifVLo6X14Mu8Gjr5RasgHbdoI0INE+fmlYmHmomsl4Gx3y1tfHhrLlKAABtiixdWker
JBxAXbM0EhdsueJH46XCoggHNtJUSnBk0E+TLujf9x8S0T15FazHL/wLQTOAfyFFTmrj9Pt/hGR0
V0n01MR2vyL2jxo5iXmZ9EHTeJ1cUUusjTQLg+/y3iEYoJlTedAxTDfGT7s9Kt4o6lDeIs+pe3Oh
+dFsltlZd83cciFFr5HK/4bEhdVasm4EEZ5U97u5F4+zNJRGlKvsIrJg6hJacdKtwc09Lr56sJG5
vSTFs1x+15k7sWlDNgxNqHjPbx/c/+poYQTX5TC5ql2W+2izbc7NTRK61eeUaN6PMBZtZ8nH2Fak
ZKtTCKPBK792PEQDIzacre5YYTf0cpyfk/bWR6PvxLLzmZT1tNOunXSmu1pDg4UzgtLsi35duvVJ
LKZt1rz0wMIZ/e9GRdHGLJstp6P3v35T09eqmL/Os5KLeGH5uDRsk8qP7/+Icp2+oIdhQkTtFGgF
VP3UnzvJA7e9n/Q0r5ouzEIMIzK/C+nXd3waFuIKWK/oXoNxAdE1LcIVCG9WNZTgPLKIbbXTOR0s
84nd/sNj3eDb6Lw3PboAP8R+1TRSJSBRKTSxppQlzOa2UcAmgUlLr5RsdAj2xF2hjqjBPCjxLCrD
FEOiGuBjYRr8peqobq3AXplT8VmVk/g5tYV5LAwblujgtMdiHdKdd7A3Jt2Or+cLu8tWxYQyz5Ey
jV6+xHWOiIPavBRjYbd2QrGvxgf8uFQDGEPlAZeMAYusqY3d/Dx7N4M1d5LIEGs7qAaO9F1Lofs8
pXgImiiCQ7ojchCuAzxEhcY8QcULIpzKa8miaC1Wj8qy2gPMg6aEi0ZqJF379mvj5lfLWs6sTZhn
d92hWM2BW+Of8eb/gSKLNxve+LErIAochliJcsHmyFrvRktwJuBRpfAmK5S54WM5ZUBK8hpyj43d
wsn7/TSi9HwhqOEmlygojdeZsY9dh/5jpvhic+atoNpLvtRG8EXYoyvMqeeJeGjmz640ClTUYTcr
Og0Duj6FY9DFcWifk8SVTBmJCoFmBRdSe7c2EWJzFucWCz0Vyo/qsT9x+aHmy3x/8oJ2doLJ9PSa
NoCwHjUUQEfwYhlRdW3+n3eQmV5wIo+oi6NhSbCE0PdZ4hymB1CKimezJWxcr2Mpar8TL6ujFJjP
fF8tc6S/81YwRJUWsEcUehkErBCNnnpw8XKgcfPGKZ3Ya851nrGV0s4JZA7yA/C5Y7cHQujM1asu
fkG6wFJRij+cplpExpyrKlhqX91/7KDMic+vFnhhOupfweSEYq/bMYp+EO8p8YuWnDsMy7fiN7NL
hUSUIHwx+yzgWBqhPgR7UCwOWxIvwEGtrn6YvcCQnq1Pu6RafbigchEH+Te6ep0GYpLgSVTHrI3C
RetLJZJPkg56DqDHhyLzcT9U4oPEYy1k+fmNcSDgTagAtsRbe6DnBGeY6d5jSXSu7nDcW98atuH5
zfAiloZhaUng4b2nyRiEZHonzPfVYiOdxwbXHzZdxZ4PqU7rv3fUqgbHgGRWryyn7EVUOw2yqyh8
9nCBW/LEz+6movSfhXiVEpey5ah04Nm5nsSmMNZMFVaCW287sbTvitwUBvXjP5fqYXRFI/3ri7Zv
SpEDuenD5iPd+Awgo5ZAPl7D2fd8DbGdgXA6QRKgBRRiZgylkvpoLX58nBV2GX2uhUiY5gWxZY2p
4rAlV/PxyID0q2yGXi9wzj/y+XnP/c+WlkCQRtwdY9+17qa85n+o1+YQ28pM7ingSjaLlwg959IW
+ReGKzrauMwrUk80aN5Bh8vNNilVyQ5OPdOAFc6+3ICYdl65KPcmbgE8MvYbXoNjfuapBp3Pm2f6
QR9BJ3BI8f3cZ0/0GSt5hJrTeIWnNSsGvmmA0fv9fxLETo0e0EnoTJu9rCAvdJ/jymH3xdvRGrlH
bSugXu0nzbmjdfhfCSLtZQw4RE7ErKZDdz3MvobmMzGTnfkUuXGGNS4DTC7SKdjOqQziG4pv1Y61
dKOnTw118IMvKUX7jQkusoeVD63Os0MuLccIlim/uO2oOKMhAo5pzA18HpKKd0/aNNBPU9L0ZOFW
tkKfC7BlcRFVdaid6j6I3DBS3JSwh0f+sHEjHk7p9iBG5VkerY3hToOnMfEo+QgX6WzvD3yCi5SI
Px8etLdgAFesmCQgZ0hNFow9JmYKu5+zYm6lJVZ+UwEVi3PzxrQEcwsMkb5AEt4TeIQa9YL4mZs2
4X8hzGSmiHgQcFmgvx73fninfTNpGx4eVERdxUS4hOJlLNYFVSkQHe7Yti1eG0RP
`pragma protect end_protected
