// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hvsZXMpX4bJBg1FYi7ufrTAC9CVoJ+J17sgZJd7hLDvxuva0DEWRg+Cve4bPAjfu
+v1UjMXx96x9QNcH401q2CBvp049gEvbRzNmFUWm4aFqeW7K4G/bR/ZgEEuk3wZ6
8lmfK3Po7KG7ZHJgmtxb1nqAcZpIjeaZtFmb2gpvrOE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9696)
ohyI1LaZCNStjtl2XSSajUQ7ZzjYwm3RcJ62AGb3z4WSK/5GIPyeJ7l+MPOi3+6V
dYHpTZm02S6VJpojipcylaPVXVAmIYH5WkaVKng4c/klf+BgF7GulGEkMx2wjYFk
+n+SLzdnDMr0Dltnp+6qxjykNfaIxL6rrz+le1UpSPViCjVAOI5W0TqHADtZ39gv
qi9kk27siT6Ylm88hQqtq/ZvA63123zAtb8baEY3BodtgE5Zd4J9VFtyXBIs3y8w
6cHgR0scTFrCwd+G9bQaNwhJGnuEEMeGcm9PS8aBo4gnckMdJG9iiGnymgjfMaOf
fN31Cuu8alnLUN0PynL2J50DXuU5lMM1KluZSQMc4aW6wbhskC0e3RpVtiRVoRF/
VglVzTQpr9anVwynTLSTcmy8UygRoHpy6oI4mwq/uTX/s7yOEl0w0p1mzifwxsDk
H2APH7mq6HG3YqJAcvi9e04mpoZzrXevUOxBgGPNA2IpgN/iebQ1gXJQuR/VE2wA
0BPsE2ug9aTDyBWkx7rSoRPSmZUboHKg2av0olOCYSZ9rDeD0i7tXW2Ko52yBy3P
kU3NmCrooXmpc7xJU14YnWgPLrC2vD87bNHNwXJNq2nExY+aX83o/zyihMPvoT9t
nNMO60Mb+1VtITvSuJfDBbCB6Htf0WkAfDLIg11G2c1Zs1mYtYdKtsm6EptfNNI5
XmtuUDXViTH+3ejQi4c0KYUGFydhnfW6gmNdMMYT/snUxVVubp56ZXDQIN5KWv0h
24q8xU6SR/cFX3ML0Jc1IublP5AyI9lcJjpd+6yN0wJ6OxfPqmlCQdCLQD5JFLFu
i2SDZ9ambqiQ4tSXwj9xSUxlQhsgUuIo23Yi1afZ5yV4ooFcwhkFJ6v4n7h64Jrt
lDVCwrus5U6JvQYro16T42Au5P632ez7dGaS6I3NlY/5QXR108wFt/YCv2eBXYh5
wrd2PpV+MqWEEQu5siIQyQwz6LqcvlCkP/Reo5H/pJLXDH60hTnGziRsWFPgCcvH
DINyFVzxTGTdXnnlcauFt4rK6rhQBB7bhqzth9AjkbAnob2dL55E550FLVFFTySz
9iukCAzQqUn1dtemfHly3Mz8CITWNZOAH2rXRnSteKr14V9n7L7CrAN1cBfV2B9Q
1od+JizbTAzv0sa/PEwTDX7V41RG0M9OzKcfP9rKe6eKUNooks7ObftNfxSctut2
vA5JgE91cdQ5byeOiFXv6zJRMaL0sJCvezppq2MX//s+W1iMKoYXXYVM8nStSyED
X2MCN7kxEbuxGI9bHuuRD2qsMxyrSSzLEs5G80miSMY4Ob/Yfc7AR+s9NKYwjAwF
DAYVxIO5xqwdac0S9n/ppwqTy9VmeLM4/kf2teHhMeEsLWvH4W+oqpz4KT5DWFUK
juwcviRlDV90v4Uzq5P005uQV83hBBABsMV2IEyhgHCBmwr3fBzAOgMjJVLLdtIo
mOoI3inJhdFtrpzkw5DuiyTP3YPgGPtqzTdGmzWLzuJBdftCdQbqkhDN8gCZp1Xs
dFNwaI10vN03xFd4IlzuU09WWtRqNthkj1nuElK8b64UCEYVXrOL8rAFLHZlR49T
SFRj1wnvfJ+P7xoin8Hyfty7wjPlRcfoitqtvjhq504zlWarEJdE/lemXyEKMeJ1
NiWEn41Oi9M74wFh7tiK6egB75QmnlXcoC2weGScDQixbi7tmONSTQKDxD+cUDCu
y/a6ryzk33ep8WWPuw9txt7kzVPkH3UxAlrgu+s3X8z9WrugucJhZIso98VSbQpw
IS9k3OiZbwJXuzGyoN68T7TMYzKE+XkzrEe0LkGb5wueJwzNlyRsTdVm7xDYpDyb
sIgXF+VF30OLx9tUDHEBjBfR+/ZTsehAUo+hX0zm7cjyIrd9lhmDJwiFijgAqjDW
P5T4tjLllHsYprcIJAbxB1OPovuBCWjO3ATGMcUGzOEjbBLTlkeyC4gSaaDobjvf
oyCiDWd5kTXEoMxsGCq1OF0CEtgBS5ObKvAyQGJUbU3qLdNE8DJVriDZgKmIT5tk
7HLMo/Od1I8IpgnWHmhVM5QHphTgmvkXtCmFRHTQtHxfhLHE4UPdZLDYpeoMbjzW
m1H4VrwXkrFkbZbEwuK9dWp0iCG61nrsG83jlhQKnq1x9DC3ECGMCpMWrSDEFh/I
qbRVtLw3hg0yxvzNOHJ9spG6F9HeHtIRLMwhSNCi6BeBU6fnGcIAiwR4yN+96yUf
oAhU6ATIlWqwUp8WP9TibAM5j46sU542EaaeaxxeYH9fGHprv9m/4xG7xxbQs0xP
+CctDT3arGQCnBv9GX9cQ9xEFKQWYp/bkYcUw9K6F4CUUVI9CeizhaBwKJMNutnM
yfr7T+VLI3tK0hKrbPIAI28cFPRxna++5pqwNVyDJIQVvAy6xmgAmBrxi34ryXNa
RW9R+gsDQ0oKSpqvwp/2E/3cRK7QWznIAUF9GXXoA1LnUqgoZApz9LgFtTTlhIQu
xYWn2lIZLXBqW2oHBKsw51mtYEsKtstRM0Jm+JsDEp2gy0Tsrq6FDdoDnAXQVTm+
B5BzhYjhs07EKUrelGHWZR8c7kdP9vDHrJMgFYasZwCCbTmcAqKF+SA9m0obrpj8
wb9uHLMDpSgaUHQPOZxZ9rNszOvNtvbS5AjD6AXn74YEmxyAh0b9eafciQNrUCnV
QiLPnYYIqKpCfRpw0mXA6YHIUTtncjqoBtJ8LknturS4YVFf+wCXrOJyL8LYGNxj
8rZwqNnyrb9elA3pWxMVzMSMg6YYTdTaRDMKN+L20p0UKQ8rvlj33nUhjS8+32A1
YNQpdXnSmaUSAjslTJ0vxxFUdT4XaZTjuR+O1uStm7zYphhGi1r/cSYuRRsjuQuL
oiFylVO7SBCoHuGPFUwLHakDl3fCQM5at4nYewv01gvEHWHpD19PasMGippiJ+2i
VMTHAO8te+looTEslJ1KQc+F4gCt3onT7eHagQAMALA3o/urBzfXuEPd9oifXcY5
NwUVWgXLEX+B1M/i/c8CljVf8TptSuuD0an2Ki5eC1FihVPumsf7ORaH7gtBXYmw
GKDBr1co6XH6kh/HUrIPPpZKwSWntBgNcD1Amgv3/NAu6yh4ah9ssxQmDFslkwps
DW8PTCnh/ictJ86lCF81zrdBKgZ/LG+mZET3sVw16SCv0z9kXog+Tnc7yvVrSmAK
z/8K7ttNkJpKUIJXkFuPyMli/qFpWHPkHeswSUaoMZbE1wW+rLUp/ZtG2FRjlfFV
kX2lUyj2FOzNcelbcdL+vRA6W1qswmZgcHb45w4lRUQHhhBUhzZSzNCp4qlt5nWZ
ayRy3FjP+KlVgrkkeu9K6lAZ6wNlGG3qm6SUJ9E2VLpHBm5JjxD8OtjPv0VihRrK
t7NrogsToE8Ms79pjWxfSb8SCx9qmQXfHPx83ps5e+pC2i1SP4YLbQhwnfadk1JB
Y+S9k4VQUAOHawan/jX1RhR4kWEGsvLDjuyrbXPblewSNfXpV5YXIaL84BrT/svL
CaCo70oOO+ZBPxYUtETtr9kZiwk+HWkMiydljoDxONp+NpvahVHb4vCSYCK+Zhk9
E3i4M/D3gHv+6UglqbgIqh+V5H5oNqqilRJmk5wOz09BG/WLQ6qm12zKe9bcRAyu
eZpsKaa1CB+Gpxy+rWG8Ov4jPFHsA3qf3akGZOSkMKONtXXI2tKdd4mGDzyacNco
2iRxQNJ+OossGP20rTspq5gXew128i7DSgUPTVOcKi77ESvVACu6VH4E9GdjxiDz
U8C8WbB+1AKzj5PE5T/OR8gyUhlcNcAccS3iZyxfCdyYWdX7ppTfFzRKUP6Fw/Sv
7PbCfwHZKv15jzjklnYVsxGvZGVoWTLKYtX+ivIDD7s+sS1DuwsEKIetp8bTNGj9
NyLapgssk3Xhuj5Ba5ZJHzhv4OzMipK1VS+pG5KFHgKlIlzIv/5NfkGrZT1xQX7I
qRXFDmWwr04n+/J/jWEgS03Pa11dnDNCbMJ/SBw/DSpO7jBC9ctSasCLryVaodBK
hf2/aXJ44EtYWhsXKlOGiyOuw5S2/exJl6XvqwsYDGtG2AabyuP6jO+uKWxs6vW0
GVmgRDuMuBUf3oXf0QkTutd7CcKGQRNem5hVIsAmChQ4onnP9ZL5JBPDKHDew3Sv
GVZZ67HNwl0kQoWjBNK4tgXP2RSI8184b6G+WZk4meU/d6stGS6nyns7D65iXyCS
73HFT+PH/ndU4tpj9w8WtxUtan/yl/fg3GVjNxjNmuCa3G9LXUdXsIo6Ueg5kyGO
E05A7leoP4ryoWKow6NjvJxUnTUS1I0GuxVM8FXK0LAFKOZe2sfoAzEyAOqRgjPM
jhfCBOBKz9zMBZbUsbph2JM1q6T3bKalAucfhSbq6g1fQeD19ISkeq9CwzYwgak9
Nvpd0jfFDEIFOtPkBEHreHxcZ1otijpMVXhkyTtYuyCNW8+UJyFjPGMcpwDuIW8J
2RmvyhmBzSFZcS/NL9ff3sjisdMvlnJvf1QPkNrAORUtkhzMe3RLeda4nUVDzirX
k9EG7AJ2IYXx3hFm4/G9xAM/k0BtAZmSnh4gyh+F8YuShNXKtoyvW+DnByxYKZxv
5qph6YZXgiA/V0UAwpvwFpZI7jsnMndjOWcDmpzuUO5gZWp1mgmVBnzwB87dncpT
s0xYMEGCIfzHBy+M0VeFxH/AbtlZ/QMAJzP5rLydzaoY8BKiBZvGMu0PUZdmVr5q
/R4Xp14ugJkKI4/UJeQYbc9n5hSwXj30EXhk+a5r+h+H0UImkheA57noOgST5n7E
r2XcNJfXJUfIitO7aCfQCMCdxxJkNmyYlmriXlBxKAyVIwibG+pPMJLmbITlrl0Q
39vflbwcywaRBy9ALcsT+AZW5E9T1g9X7wSljhlkIvQUjI2m3yEYtGOlkwP5pNDC
+HiiefqjHGcDJUQm8+QNu87m0/UQhMc7Mb4xf5wqXjydZH6ghxSbHNZLF2mtOyIj
FU5CskXzkncwv9uTgiimR3eCupbIJv5TvqDoheI1L6vR6GT6IYilvcaQ0QGrFxiN
2hf2iUvGraTxxdpXxS+0uEscBix+/ANq2VOurLKboTfyYXrauRBXAkFsgcnVWAvk
bSdZLb+V/IMBTAqlQRyUUAS1zGj/UuzZk2kKCDgO2JTDybPxqckF90jLg0f2Wv8p
TZJf+thiDAvU4Svpoy79johSmFtOdOvRhSmyMCE1AwOjjftH5uiy/WzFz5OeBZQF
hwbcP1zORXDy0EtXwgTvGyqcJUw+ljsKwrRCtV6nY4Psm0Hm9WKX643xi+bVBzCJ
bvUc+/vtJAIWNE9SjvBCJZlwdMJYrdD801+iouBA4smGHxKVZOdy8wKGKs3Fd8F1
CNLyQJRskBdXMr1HvK6of+dUqjf0FchPkgWVAvNDXD4sPVX8HiyFbtHZPSN56Rlp
sv3Awo0EZ52g6Lzt6/TsSuW+CuoB3cbtT9F1Gjye50g+S1ToZ9LprPQya0ETki+3
BB1o88T6SWBetJQ0xPfSzGGO50NyX2OoHmX238AH2ACJasE2omLY6OJ/5HFgfPNf
o+DXoL0pGzF7FKh4C18eyXAOm+rxCkikFsrblftRdVdtscFsxIFsvTOU8d8QKc9W
+mCPn4yvcbjAIfpd3iXiAFRPVXXrB9QGJ7CTLLoIXa3O5dTgnMqaZOCkExpop4gQ
Rx3hKbNl2jfJM74eFKnQjtWmKwEKlyquoIc/fbx5Ai8/QbYwqx5lZInPCGERrgJI
7bsL58mD5uBTWA/x5TB/Y7hYAr+QOEaqpDZ4vXumT4CK03vxTT8692rivHB80bq3
LOx7ghjlBXQv16KLj4tbVjvKrvf/5yqhGgZYMlpXcA8a37fBD6DJvAJ9t8EReeat
0OjoXZzuTsxT9Y8BaHweqLlJXyGP1x2UpsEOf58R8NRSfLHbLJDQbRZS96Wb8DPD
m8pVKqfR3Yir9SEkylktJ3Jvfv2S7pW0UcsOxu7FRjYma2ZLPu3+H1bgwoMjDNFE
g76KhNog2owPDGSJ4NFc229tPTyWfn4th2dKIqJanAmnpDmUi6Or4bgnJUmzr2BR
b6Arrr/WbXHzrZyHHthmWoxnJOyhV7dRccqhLvVmkWLfjh7/eAvKY4xr1ZTwBXsQ
ryEy87EcNMFKEwp+TmK3QqPM4y0DGGh5RPVpQLIm8HapU1DV4wgbCFj3oQ+1Prsd
nS3rsIRBo/4cLNhP49cPkEXNF4toHN3+JZL9aXKlo1eh0XtLllA3oJUbhq3oUal/
NnoJT3/sXA6Sx5NHcEkcN1Szi1VsnhNJjP2UYrX4/CghYenlWIT76vk9ZPp1cv/B
ZRasITq5MSoLlEA8QVAKjeCxOlFPt0Re0BTv1EdSFaDeBCRGK/tFmROEPBaL0QqQ
+sVAohj6c4BIeITBORYAaSi1XEXFmlWe/xTHWbc8F6JzJdZ7C+YgTBSyJgT7iPQ4
YR4mv51mXpmb4Gvs/1xf1eIwa2p0KjVYMoPi1HIh2sZgS6Pl8Ze3Len6p2GySPWx
etqaCFAIdB7IfQG3NTIrk/jqElOUwzcf8qnd+BFvNKhiqztUDXp8CgmHiRKNLsOZ
v33U9+jkmoKYqbfzT4MKr2f4X/ggnl6euspCwf4lABIQ/k/9yyMYG73iYkUNTkZZ
uaF71lTkBul/+iEViEB+so6OJA0xb2ZKbNnCQaoMc1w36rqprm2RSghWijN7uvWk
KBfkw1caIDJwx+1cd9lz30beX3Icb25vkuIccdV2Bk+JTf6qDxHCMkFPBHkuFe+L
i2A4XOfqII278jilvzrx85j/NDrumBzmmXGVJJfDAi1vytWE6O2pNOXatKRX6TXd
kmrDZuu82OZx/CNQV1ADDO/mEI8E/aaR4gZPBJHMRa7aVFnKSREKvMWv3yv23mow
1E3poiI8wpjvxa3GlHsMlC03VbaNgs+x6tmtdFLbLJKnSu4+5U/5yqg/GGJWUzvd
DV4EaYgAYxJ6dh7zUXFnYaGrK7liOHR0WYGsx3FQMkqztJ4RHPdQ/KTsbwRsL2iX
vTPLsop56W2NsQyV+tGfFd+irV16hN1MOSeUMeofqZAg1vzOdXq86jtZwcE63Wjd
E0KmxKwQnoWc07Ba83WmYwZ7gwQ3oOQayNeJpVtu3cMxEk9N+tRW3n0yqvTn+++L
ZwYY8sqKEp8y8f3WG+f8Tg7wvbnHsnegq1ZAdr85xdnM4uAqiZzZvXyV8R8UodZR
L/QR09gBolRwHTVFU+cDQZkPxkQkBVVKX8rhYtsSOCLgv4R43XlIE6L7/uHF3xPp
wbFhZaZzAVkkW9TdVp8myIHwFlDWrYO6zUAmWiU07guUB9JfYoRzuzpFczV0RYt9
nsGIhG6hcvMMfqi7hDNsHDf6fyFVr71GF9qay9caVaiPYmSz4eiVpRLNVSCx8i0y
T28A/CXLfFwxfPXQuad+diQb2iJwl3uR7hG1lvS78QjtA3YLLQVQz7sZo16qrMlr
BWXp9JB0PYJONRqBCJaGY91B4MivfIjwKPdpPzuWDTlMWO9aivCVMl0NK52I6JOr
f/2qDoYA1m56JOTa58qjRtJHWbLUaHbyAavA6aaph/N3ghOLpx4Kq7VTvpi2DSQq
Erov5lom/bVryrCj1OnHQsbFHjsEcIgjh13v84MDEQgqjZ0wCTC1Mz8iS+O72LNz
wBwcuRyGbLHbnk6WOJqBVEBPnHy+I+Vd9JawDWQVpw7R8y9zNWBlKwV7b3Dlwv5M
C/laIR7AzZpx2DcfKv8BgSJqo0vzlNj9A6t+sKoudDH6zbdNYfpRQpnKK7UjlL+Z
lcUj4LYg7AKpzPItzvY5tLxzRsr/GuK80LZCLJWgki0er3eXg20HF3jnBV2YWixp
YcFpdYz51anBI3fiKp/BXWdjSm48ZDHBx9O1GWhQC6hIndLLm6827pKtLtwZUpnP
GJwv7ILDjYN1AGp2CTvvz+qKF9/bq+wFGi3Z7y2jR0jjucPc/y3uR6NDHCCTip8G
zTmQ49RxFqWuusrjuNe+6znJs3qKH9XTMz0IR6Q3YPeor0E978ktM5M3mu1chdVr
0ISHgCl8ds3e91fD5h+3GQF70J/afIXIqvDRq7n2oSHN9Ub6d6jpTRtV173STinL
PKsl6/YUt/9KqVP41ll8tSMZ06q9fJLtrfe6GJ3c0U9SxAhnff7TmsOuPGaeKGyj
xGcQyZ1JdAkv0700SFV+HdTVyyFYHSHlK+JJLRVlivrSG1qmdw79OLzfjiIV+N/+
ul6WnymClVf3bJbvv2R+7g+pJTrgPevAptNe+wGCU7pIWmn8KRxck4uJAHrjJk3z
cx+QwZ7CCStXlIu2l3qSpxgt3dQ8t5Zju3hEwd8NRMBAICvQ+E8c00k7Vau+sQXU
VYJtxUQnii/+xrzGw9W6Kk8Mjv943qqnVVI3YV4iABD2RQJa0dN3WJV/kXsKvK1M
qO3WkIR+X5ftuMJ0GJxIKK2s6eWqnJfJ7WzyEeD25ji+pe8xt+jCF4jGxYlt/tJ0
qrWKV01DJ4RSIh3VXkbg9ktpe07QLrcVgpIrGLW3gDcXA7AoXfeEsRNG7lPWCyrQ
Gu9a3A8r6KsWLPsuY+CJUdbOXg3wUvv1UcXG1HMqbmCjWySbN+fBApbZ4yIsoHgi
BnGUz/aoq/x0i9FiAQEjUwN7JuyybQ97Vy9sJ6z1X8ycSDIw+steye5b2LNggdTy
TN9OqYd6d/T3fEdpj0AmITm5T+umO6/FC2gn3kLGqsvZfw/Ux5wJjwcqpcv5ZNQB
EXi7GxPlHGmfsvqxyk/Zip+S3a+NNehf+Fe4OxaYsSKUkHKxq+cd6uFDkgUnY5zP
m8zr3txF7FZFe3lI+EHhkQ7q0/lWVtcDPa41NFd00UEH0DIhUw5r12GZvicHKQ0d
WOLeiM83uVMYRBdxrouTpQrLUQl7ciGi41vRyvk7oJ/dFWQpb1T95HYyzBP+Vsuv
1oa+Dxn+6rkAqs9SMtZ6Aep8Lfw/B8uk82PxSFRuZaO9J4oS7oqlZl0MWv+TBapE
G/Tj5Xf0Kxw1nZrcV8pdzC0zsLjO4N8e4ucdV07ttqZCCB5pda+oH9UfjrVATnnT
pBzT1leGOPi/Sm+ws4IOg1Ky7etNZpTA0x27xJtKfMAodVlOjWBBXFueT4edRTPR
tnAO6iae5i2Mzvr91U7gr6yDcwjgCt79CBXgJ2FGLZmgsE1oQkxONB/MZO1N48FY
ZioIK6TPgs+KJKab6ZRFd62O8EHhX1+iix99iAoL7U2Oq8BZkVlsIKHn9EDTkmqg
BOBYq3PBD+mZkFVhRewaZGiM/rqGDaUzgJKSVDIaTf+ZsIEqZfs8NggIdZwUsUz7
wZgX65IAUkTiLLWGJHiI8dxSxNQWM630KdpLFfuIF5vOzO/P1J2xSE0YzNF+evPc
XfuyFnRYlNqT+SbpwQPmcTXK1GNYa/T90OrTkbYql2YSnlWIGHTw0SPH1V3SlWKT
n5as+N67EY98U1yKr6+Mm0gGHzi+bEvYnPZNAcTfQlLIrSMA5Fm9iO4RoHmiiuw2
ZxyTm5FzAJZA+Au3rKkJ8By9tIhEBt3pS6PWpV6Ige/M4EVMqBXKgl6nyqJSWKI8
+OFS3zKr6Fn9z/5hp1NdonpQZK43Hr0WhuHHzl5ZuiEokbO76dkkKpKuiyyaxSAQ
eW1LwWDwq/Z4HrwDduYBvhIcEi/3hCtYfxeU1kVG46gSWRkT9Afq0DJX3/pWduBn
fuxeOgzM4qDJYfwXAI6wqnl69G6M89+/hEcDgWl9nnuWrgnYjMvX1pBtqDhbD/rx
7Crqc3D/hMgWN5yAyejbqU0Z0Sc4YLmNMgJU8zW2RnAl5z3Dds7U3o0yBRWyxBqZ
A/OEtgIDsEU18pf41ZqZoSPPkFLEloB6WZTXQERI8PvDHvOGaw947q01UbOe9bGs
Nf9GUhPk+qZabNW43kpAqSP+YatGrwRsCcQznBRCsLvqb1KXAdwP6pK5LHP3b2PE
763p/HlGqHeMClkJXN0RGRwGBm/WAwRrMKBCl0KTCp3+XmXGDnOKiVwfIiWk9CwM
Uu+4arDHOKbLL6peHUC7nmB8U4iVs10t71ho05jUzyYTM7g7Ox9wXg7mQCg85/CG
YDoh3RtqxkcIk+8GwYSS7X0vEIbcwnV0ARZL/MmPUGTqFk39Qn43VU2iSnTkZXZr
VjjdUrZe/RTTvd3KVpQtTZ/gI0uK2kdVMleF77Spq67WI4vYflHetu8/A7C7zTGi
AjoGrx4DVn9mFgmA9dQSsG9FivCWaCvG3I+ojXemQsRReBU/9nizXrZ8Z8+J3ymn
4Hc1QVNQZF/gLOUmhGnpEEx7U059Ohm8Ps329BRzL2C7fKhPF9GTXyOfkZNVS81i
QRzAlRb/vS7JaEjpY5V9G1pCBjimATRZRDrPMfSSW9PqBkIIUsXeGprSC2SZsoMb
H5Vvj9yEdsQVaeb/a84BKMzjmpf16cTQVhfiCXlx/fmbq27iFVyle4WaXEMPinwO
OGNNCGM7Y9mGiCvKJbLgZp4WHhoS+QqQPukhdonbRXJD4GlT2eTbatJ7XVfFo8jx
RwqdXvoUKdkw+/voeKV9PIxi+iIR4XzbZmOLV4xMlLExoA0j/tbRIcpIwqCz0Loh
bVPF3TUQj29owpZpbkjCZl0qBuGxh6XiPAmJLgzh+s9Y7UnNVIDOE6kUZMrzSBsD
IJVxihOm/ulpsuxrOdkm48UsBHtu+nFbW8Pg0q8UDe0J9P72ZgPrjy/797QwafyU
nVqQWkoz/x6z4kfkUxNXRxdsbaVvFjsywjD0gvaUp41PS6hfOyETnAFoU7a90aZV
egIg0H8G6ZOGDfM4r422foXkSITey6KaXrqQS6P5trDoUZjNgEQWHae7DtYa0YGs
HHK+dfZ4PHoumOqQvIPm6cV7PhOITWZI3nonGwSNagWof89pg0aRXeMSU0YLZ8az
0HAAKS4Jypv3A9c2kHotOrTOmiztLhDu+Sm4KNcHXOCV8FBeYJ/4UW3gQ6L085Yv
PLeBQiSLhX1ykUWOy1SRdUg2s4b5ERvK1j3bjVJr6qx7teNJ0oq9nmupf6VXYecu
urmo6Q4ubaE/4HFuSrQJx1b1ThYC04Zo0VQPpH/V06GyPfi7WmQCydmT1LsYBvM6
7H+EMYhCjTkM7CBt8lyrihtzWkBzO3tDIdpAxgrx2OgDWHLUeHnrvvrygG6uHvle
1wWkmNNGGweFo0bWxdW5ahVtw7j6Es9yUgplpV0u/sHEI0ijMSItcgoLaAx+BXW6
9t1lBFyV8IDOIRKDoFD9DRS+6RLtYtEuPkkjLQ6EfUDej1mLIxGEdqDkNb660KEy
3yfszuxPRHdLm/VWPAR2zo6bL1NyUVpZ7s9vylxoaZK0fYhU/GDCo4zu6Qg4WrNB
ecsmSowZZh8q19qV7NRlvuHBtx3hjP+507AOAf/s5tLHz4VgA3rSFr/WmISj+hJ+
kUgVILLurV7jJxmYAdBjSCnBgXSUa5CoWh5qJRyNx3d9dC2GG2dEXDpMH47tdQ7r
3wbIG9uHiYzFsjDRkuGWHEvw4UPCxJxYiX1WKFD6O2l+txoU7vhrV9yx0Ly/gs8x
D4QOaqCURW23qN0HxDvTi6mLs2gW2Y0xd4OVzl7YtPHKv4S2E6s38ud0IaZqFtWF
ltB4XGaqpU8y4e8WOGjvt8n8AWKlsDCOHKR1XxwI5JuZXF++zSIrfXgnl+jKPSSa
fuPaCOeJqVvZ7t0Xayh5Nyy5h7bqG6nTlVRNFwHa78qw+p70ECvqA+vlxwveO4A/
6lxRKRaVNe75fbPteRS3IsXVM6+iGGHMtcdIGiUM+PDewhA6C/CMnqZOCzZXGAEv
xtQddPVepuy03KTYDH7tgM2LsAg8UmfDPYmKEFMjQHJF9ZlidCMSKEfnO4geL9zP
HLtvkaECSCXHhZRlrkDxN0vbaNngFhD7Vxm7pNxCgVhgSaZtS5HAHyKSHDNjQ9nf
SM0wl3qZa8l5SNZFKe5lnFzpkzsxToWzGqAS/SRTi850MaRis/+Sz8JuEqUjR6tY
x0kpjM2ummSahSLuvkCjUowbu/OrJqMfpQk3ZKjBD3pFhmg8tLh4meMso22jfbz7
enub9dc3eMKW8JDQQCWC8urYtLgKxMZBHiv5z7d3lnampU2v7U7vt72GMGFTCc8/
pnUvCj45HLPpVBAn0EfZWohxWV/qNeiZOV/0SXCUaRxSMqGQ4nrZlPNtDAB11Qwi
cbg2A3unuaso348r6mI/JOAfQHqyXZmH59waRhM4BsyDLz6Hp1rtDACoZr83pbgD
8Hblr8BA+zMnDctzJ6jmVs/H2POaFq54Qp/qEPL2PDnaaNhdpvo0TbqDamrJKePX
5z3IJrhKdtWnEtoozzuhimVuPPQcraaUfw81BQjzdS0uxFiq9rDYDA7tDg1dP1C1
18/Jq2h8LqNV22i59tWxrp6j79LnVZScjzalb8120iWaA6s6log+QIi3WGRJKjck
AMpZTSHzeW8kxif8IkcqHxH479P2pZGHGjfzHZRSVjaZ49QK6NzZqWdpY/rUeJkN
2ZRaiD2g2nz0ZBBI4UYcph+cYgLH0xdSyO0WDIUHepIcJuWjdhwu9/4foqIWbpId
cfkoWMoKn2HxiG/GPsgHUjWsMpgF6fi5qHppaMc4Mz/ZMAFVBMCez5QiSB/xfKZs
+SNuf/zPW4inaYdFx50u8xZR0TOlcGZztDT+lNRKQnRu97mlINd1vAneNoI6yJEv
OSMA8hFo3pudgFTsa5GNxa25g+5i5joeSz8Q2BPb0DmtaF9fUOfy+rU0rS2YJV6c
1GFcHEtBk0T+yv9/At+f+UYdA5sHOr9Hma2mysTjWEbN0j8+Ewj3/NqwQU8ZSovT
Sh/4nFM2YPIa+zN5GaSSBTynCEv1tP+iGSr+cSdtHW5/3WlwPPsWhwihK2+puKg6
`pragma protect end_protected
