// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YE33QnJ23aVbwiM/yTFRc5xWwY114UPQSJAob/Dl1vF4OAbrjLOB9XhO9GQ/oBHN
k5nRovUefTb3wR0IexPiOi0yDNAemO/CHtRg3vA9ptFk2AosHCf49hyM2Gn2NEKz
uMLo5+zzDI6eaVdTD/6ScWajC2RUYvn5ApVG6eJVk00=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19072)
VcM4whP9ZFfrxi/d9UblhEuSDNOu/JG1BN/gm4LNvhlYvehRfLzsj/W1be8RpiJj
CMcKquI2YdYrhUh4WRJvybaHbPXDpnXwGUGEXRpoKC6TSZIKg9FxK099+M0e+JAW
9gN7mInG0Bs/WEEPRfWr06QPsk5jeEwEGg2FuqCCsMO61wCFl6vgkxEImTp6A0qn
XXW4or6Kd1dA7EkuIlPyk8uwLrIIs7j1VhvtXKCP1QrtntaXQy1l10d4I0UQKxH7
1PB/zdAOtIdAG1Chl9c/82s+ekmwcF8XK19+qcRLMinNVFdCBhE3eVO7QbyqcBOe
TYcMVRUl93lpgovceV15aMH6WwIrenY/RMbUw8HWJuXl1lmukNwGbDQepjqn9zQa
vurp8rlGhTAie1rXe0XRbqlTP++UVlYSvarYb3KzmSPGV/OhCHqUYlPLNoNBuYPv
8AmBhofkLGJPizSxjRjg6txAgCBl0VOpMXyzHwaXilXYrrobXuwiXLR5Apila9t+
jCFE0rhZPBciyVIB8X/kP+1ETJnzFj+JMQ9g+kMFxYxY9jAGjX78N/zN+Ixg38HZ
MXRPktsk9NuYjnq0uxRgTohIsymFOmQAml853RNa08PGdTfBP0TjXkGt9M8cmIZt
LOPKFkpJML7kyEtcEbVxC0zKmYOJITg8lHnfF4wjx4iHA1q12BieIc6N9BfAOP2D
i5jMa/FEDWJt2FXpUjUJarkk5qAmGqXpvLcust3GqpU6xld3qXUDWcds/MCbMCbP
ZyaA29WQoZgWUM70m701mz0sH/b7oW1jBDIP2mgKykqkqCdY2rsCNRKdKOWLTV9w
R4fp/Wy83ekjTtBN2QgNKS4ngOQz28IPQlNnbl9goBVhSSbqglIuD7qpUA5wqdk5
al5B21Qtn4URJyNueciFRtGTNJWShE51pekyjCJ88aQNXXDiYZjIfQVLGw0q8zLE
64T8oMh3toCprZu2+3KRG2pXAROzSgp7WBTBDA8xLMpL8L7SqceFKgP0bhEb1E1v
3J/2EHT2ADv1N6BsxxF7+TZyfZHJA3Ats1WxFHw8fu0UhHVik9+AHhhAtmENRAau
U0pVpFPczbfKzrc/sYJKZ1SmKyK0+cuWlSdMfZ7tR554rM1Fhej/6sh0xI5J8iBo
QRADVMWhabn1DH37MUT0lcr+Qb2bQRF2QQbV7si/RfIypwFOPp5JgKSzhhJLPfp1
Jr3CGv0vMW5maj8sHXQV59lZjns8Dc8CFTG3OUY9Fbrn1JhRoOt/7+mtL/NjZ07f
nrVakoLt8fv4c6oCmj3N+B/JFgTTO0JmAbx9BtF396YeQ37ZgTzoltIpfusp4GWg
h2wvJaT96HfXLNWM08W7u6TvtuBPg/1nv3kP7YmP1uUKek+s8hrD9fWlsiDH77uQ
+lld7xbGdNP0ANiL6pjOIEfjNvI/TveD1RRiQ6D/bnSdbx9FGg1NvHKz5QRCMaSA
uscp3+yBi/+xgr327g8yLC2g+6glAwLCyYWiVgkkdbs9MuNYWQFsKfvMLDWQRU+w
qHYTPRKszR/cX+dRmxx7HGgipa01qL9zL2UJHac4eSET59VgzuJJbQrtPxX4t3uT
6T4ZMdm1zVJYyTzdX96zEZxUNILbGScaRdsGgB+xahdiOXkq/K/lIdATcf6PskpL
TGGnnmk3jrC6SKqSlXd7ov3cMeT5KYamvM5ZJLHb5FngRJp3Pcsx4oE7rh7mljzf
vAbre6umgMJdJUvmvhPYgcYBSdtpAnFmdBRv3gC8GFUykL7NTsg2IAh8JPE2hqwd
G+tz7vps/2aNeu/qAn/XB2nhhVrrYi3+V8Tn7KYbjzDbXfVcxW/3Qe/7QwAMExW1
LYHsdw0XBeDBY2OyW9JjAaff86icovthzM+P1+AZunW6yqG32jc8GIm3LlHWzP5Y
LhXXXJ66zooRhPieGXu09b69GLqb2UECBBs0VE76kC/ntFjc3IffH6wAjfpO9ffG
R4yjUdub4tTngafxPe1791LiLl4LH6oBEAYl+UTvmUGKbkO7Iyqi5Z+52E6VYevx
1HKLhY+apmZd7bhpg21xpkOGuMYZrz7PiTKQ2Jy07s2SOevu6ObBkTUP/KRsWiOb
vg0DlyXpqVqOOv5FbDaKirWcYz1Vzp3wB4mr2LVhDh0rnQYr9VIU8nLXonX18RZe
fxpSG1lLksuzkOtzApx3OX2C2s8glk8T+GddO/oduyNTc9de9su3klF1hC2cBAew
/Y+ImaPy/4Aljz7rWeh6Sh1xa5GLtKzqlxT84JRCA1Seycwz6XTM/T2BbSrS4udu
yVhsmW/KjBWeBC3XwQwq4h9sPshCZcr0m/us/tjgUzr6CMlkpb7beevadI4enzCZ
InUoobyrFzKYUmRC5A0qGTDhHQmUS7VsdSdyMEPkSnSmIqKFYs03/QKZPds4Iobu
SDYsLf6kWemyaDzwuwhR3nlw2nq+Gp44juo4X7JU/jI5mfo2+r1jcTeRfvma9/L9
SDbUyJVnOBlnn+VWfkEVpLiCG7d8SX1cHayPCsfuYi/+jV6I7g59XUNg6JIHu8RN
RHCs7RCOcb99jeKmhCbM+kltROqYPPNEnVmo/liT9pL0+pEomOO81kAgQAdFM7Ty
WIYA34B+OaaDbTHHvtlSs7r1StQB/zjoVyhtCKdUkVtCpcjLjbN6sS+4gDexRjQu
LHNS4TR+HFb/dnNcw8XarzU+gYpCCFdj7A5x0VtBHvr2BzQ9Qq4SzzkBEyRZ9jud
lGq8DnqMlox52/yIS8FzW/E4YZ/+JiFijHXYvqg0Y2aJrus5Zz2bYFID7QVY69I3
1ITwVj+N8KBep5ipPWHD5gmimLmaZS1JAj4q7HPhhhDPVf6Cf7WpnLoCBomcWVF6
N43w5vSZzCROvnxNGIyIEAjGkBW8QF5+YVQ2jtaxAZ50BSNrjCPdG+VXAKu8tRxC
IiQU2wMhsQmX0RpfdR/VmYtfLuUVDJWCkFZcxXUF4caxUTX/IBqpg+Jg7Tb49fqs
DGTVRR0r4AKCZ61CjPZ8tz8BUq7I28OM4nCatOiAJOuKEHG7752Z4sW2iG4X9Nx0
hTgvBuHK34lE7FVVZOGR0OLDASM6Od3GhaZPZ/ovqGGQ40U6qLA+MbDVfKdkzF1b
mBpq/emgGaALb0Aa28JDoIO4P7lS7T29n/uVKUR+dLaWvNK3IPR6yMOrr2r4IGBI
TIItoMIl9cR1urbuwVI8AbF9ffMZTuhLBTCMgG3H1T/FKNF2/bLGk7cawDtAALZQ
pLWZBPU8hOWnNIgSU1ZMZLv/fMLliy3FDkcXgo0gY8vd+on8OdnoPtyk21351b3R
w13QQ9zHcPqMIqk+ydP6xllN3YuchTSeOPtpKRLV7uxvi0OJdJnefPYsqVWhgsIg
PTkTMztcQqwWQ9WjqJ48RsLNpbfE2lYWbyRB3uz4NLf0wP62ANgHVe9X64BWAFC2
jyv7VKDVxsL4vLxan3mgGJYTk5HQgHtKvbNWg3/OFUbGai9l9Zas+yPQNV/udbsi
igDxdZMh0M36J06BOJhXDXW5SDxrZiG2NhKfE224xi7xtMQOgngWjaPqNDjzK5M9
FU6nM8adSnSrdmdFlkVo5ZoE/ptu1KXcpl7G1u43RXMq9TBH9QmzY8BjEvXlnxkQ
HgEwm/Ay9lKpZbNiTqcsjsB3Mt9frM9WFWyB+QXsSVTDupJSCCjW0QmZca83pzOn
GR8l7SqFrxSg8cA+JWqiOf+ZsYBsBaDxJVrH3whufAPh62Iy8QulkW03KO1m+rBN
uBjF8Wwty4GBG16fh3xnDMTftT1jr70dVI0xsDs97tRqza4SrvXR1C7aGDdmTaVA
jqeUGvQT6j+p0sTuLJoXnvZZeA4xSEVowKglvwPP23WJgX8phgrd7DX+J7dOuYWL
YIYxfazr0m5lcwQF2k6cYCzLm1SD0PRbHp47zsAoghLjKXVURDy9stiIr1MZZkeC
7KRL1n0tqmTp2dh9GWqJaSA52yjcQcVdXBPQhN28wy7/NdEjCPX6ZBkgUaIlv0nQ
N1GU/FRkS6Vl8uH7xUWjvbvGkIpfka0wICucHRECD/P4mZK2n03OUGqivsNwB/y0
NcU6yxw7bHsXDyv9Omqvsv4kTvApirY9F3zCQ3kvCFk1NxgJAXGtq9PMzvz+oFzO
p9mLQlBh/I00P4Nqh4TN7wRi2fNJ4VNYEOw48pT6GTCQJEJfVv0v1CLwFjjLcQd/
GCZtatBN9qNIRMmJbJxRkkS2rxZsvbIYZPbDzyG7eFE0LTv69l2WDk1eVeQr8D5t
3H6+kzfMQ6fk6OqTNLRMBHgQlcILY9pc6zkJRK7J8HwqcTNvQ0N9pTVanZim6aLe
260XzSJpnGbz0f7VyLA33uCBEpAh6+zYAFrqtZADFGQO/EV6j7qWLpJWGzls2rTa
PCijY8TXCZ1BjrpMxpM5aVbPW/Mz9f+XE2U8eYUh0VFEc+cH2h2Y5OUyOCvqBr8X
X6KcdF1zvGCtGGVoiX0MzV+6f5jaVEJIxhkf5oOz7nzhQf7aFbvPWf7R3Sqyi7UF
XKI99jPdYU/BtjklMLZ/LVUi4RoSwOOzy9J16Y7rMs7KxcYDe82LDIWPZFj0EsfN
+MQwMTjeT9YbhEets32asxNBd2eLylJOvZ342o/5hKTjEu+iJ0fy12pOs0x3yYjP
Wu4Lz6Dxww0Fxy2j3LiKsGIreMJPdvpHSX+4df2d1k7qcoiAOhqS0qFbeSwZG7Ed
iyppWuJ9W827xDxoDAktNtBavxwC8cZE51+mgfU9slzq0SsBCenVKMU0b+TYRSPK
lI/h65+YkKX/bfCJlwOKNOwv0Q2PAC881+alyeLHSgYlyoaHA5kJMgyCbIYkYWlC
QVZqtdi+sN6dBDzy2guluekMN5jB8gIdO7YAxU1J8tyWoecfpkGrI/y/0rnYxsZg
djf+BeTi6vMZ8s7lfYuDttrYWByLO5D6rfR5oqQS4bF5qk16D98GB1I8KmJwbkO1
dbxv91usNb6rA64OydBtRQshjLgu+z3CQMegjbT1nZN2OdXzB0gkdWwfkzhGRV74
ozWSLgxy19Cj2gYQ5W8H1LoMMH6Enb0IO3iJYyK3Gg7RDbu+i5JpreMdmvIGEK0P
wy/S+yfnTzDnGIyrhSwLJj6ippWW1oge9oNDaicsPGp7Sdheqc9bodXrLNZVh+6P
NA3JGMyWM71hIv8MYqes4x+9FCi2XCka498fjltwW0gIxy+5I+Y6dxYpwftIxM73
q1nO06xhEOGuJd1q2+vb/1Kegyd/DpKNi3aCiqWGejCn5hgzbUiFWzkmVoJoBw0v
foVXlz93MAvJproplkZA5u48I1FNBX9bEvs7yGKQWMFnUf1G1dUdspQeH06HKdth
CAlly5kjZHTCyd2cEDNdtttAbegEARKAL13+jHWnhvjnhWBaSG9cNaW5zx4ZpSnk
2LPAOJDyS84RjJAkM6Atehu5YC7ZJO7LjjoZPtSLOqKZImhuCNyINo1tysc9spV/
OlGt8BAkgEFUS9XWW2hsq59XbzQ5u5teVQjs/O+aELaXYrkM66pICAAbi4WiHYw6
OCA+M2Xz2u2pYZ599CotOGiw1vELOE4DfshHqOfhjwzZaSBPY1KiK40BRi/GgwIN
3Pg4v0TeGBr/bjuGKnCiun/htas0ertvmXu+driv6G55/1RFsgGcumB1h0qvlETx
8SrhSgLaSCXijYawyoL0QGO/lgLdeEirH5XWcg/e5ST12H4TWe63rGHZSSmABnUd
ALT5mhhzpzfkyHn8KuIk3NfmuhGdxDwCXejm+LlnbX2NkjPEi+l0AKZOOSy14OBB
p9gEL6PzKKHjCgvaO/awQYV1eIDrZlS25DHxNXlz1bM/Cvdywg7atTWdOZqaJzgw
Gglz6iYlqPRoIw2KZWZbYb9MzBCH9fwqDi8JG12ndQp3P3pVDMSnNejRQDOPiK/f
FZSOi/oi5CqVdZp8AqxS88H3b2QI8DkEUybkJ1MgZzXtclLmGXid07oyK42RUAZ7
1EfFDbyFSANC/DJadV19Q8srdXXHXDUZDp7mJaVNG6UwWGn/MZaSGLgjuQYOr85n
UOB6HgHCEbkd0b/4/FSG/XHdz1JMVZqUT404Zp3CkSJBWScWiGXUk72mAWQvGAEM
pw1tsUVMA9Cx3qExn0J4MkSsW9kMOECU+l1GGf88uuylqCFnpM2RHexNKVDkY7hG
WFEo0qiC/0neH29o3/7gK/ocLoXSqOw79Fkfs2kzdlkAIOMZN/OhZY/wnza6EJaB
J3eSj4yI6BMWu8sPDpMzp30SEDE0NRdckO+laJ81m/PbwYNBC2jPKvqEKINZw2IY
SLF7QPxeTF1oiQC6Y+uiMy09jBh+kLrIqPat+h78uyGUhBYpH98/Qd5LhtLrsM5E
58+cEeVRbp/vcwzZbMpIDKmMc7/Rqfd8Pa722bxgn73ePaCyTMEJ2eEXj7cah8Qt
rwro5lLn7GXtHCzbWaqhnhy+9VnEuH5UJec4b5ZSoJiluslaRurbvo9LKtjDNnN2
J8PFiBnnQXxc4ZoTJ9CsipOdtddJ10mU3KLOeBPwLU/uCqsR2DBV5fpO6K6srr4q
YzpWQKw9ZcCPOi40GWCJ37JQfS1v4wiqN1hRpbzos2iP8ZZ1nzQtY+s1Ikha9m3W
WsUv6f46q4KX09hANzkIwhxNOhaPzRjJ8V9ELNKOSa9h2ssTGcutFy04dyA7KVw2
Hsd5+UjJns/YGh7tk3JTXfbmHpmsR/m8+U4C+NjUwW/NKttLcDiFIbbOeE87qEKV
2E6LiBJEw7ZaxDzmYcW6brQCBp/lzBGUzq+kThYOF7qZjDIlRazCLc4/p1qWlAsD
xFYGKHK1dHFI8wZWzs1TMlid9MoMhjRitupDhBfgcU1B/BSJcALlxBbdetER5WwE
qiRqPZLipV6banII4uBiLYdi8fnpQfigJMRg6jY64R6ASbI9PWgHdTxsmANq8GTh
SscwBsT94id25jbQVRikYFY3MpzTEvPPHSL5bnqMWPccubD/a4h9S/hkKCYpIHiu
uxpmo4tJ81GV8iHt6g3jrlrJ8E3OUKvvb4TfbqruXVK03Pe/wCDpAndqinI/iB8Q
zRtMkWSxV3jYWfFqf3Vto7IVlEcWO0+cYXa3Nkz93/reV+y4cfQI3IeH+iXKda/0
O8aHhmQkmZmGZc1stUYpqCwBXQehgdAqGmRMnvl0REbJ8hzGluktkK7zNQ41HDsh
fBdackSeZJudQc6jov2NEA+0BO370ArgFHBM8ccPkLXOjZG4t0MJnx95H3mfIbXd
SOV26MkcJv5r5dHCsK7Njl3cVVvofLQWAXJAoXV8zxOuWEsYYzAC7LTN8cTe5rfe
QnsXy/6In3zyDjgWwljIuH1ADVwlLoWXZ5eUUreUPJvJL0jvD8CPTdGCLpR1IHIW
gybV1ale9xO9WRRoEekvDuxHuQ8+cnDpfWHpxKzBNndP5n8fjC2sBsD0K2z74PGY
VpNNctdkYpCxbwZD8+NA5FniILpkIrQXOiNRM2d+bzqg94OcBL+FyZwBf4aN1Gf7
TCzNswVJOI2fCPOPtfx4jnIg8j4znvRgd3XKc+LRtPqROpFbFn0neGruOcUbo6UN
u5spYl/HLxK7pMe64NpG+IbiX1MwjPtp42HrFAM9es5szsr4VZDf/DSntgc3d0ax
NqYGBYx0Gl0dlC5lZvH9KDwnDJ4ZLFChNAAeiWeA5HPkXJbVSjQk1j4fC6pomy6f
rQcu56D7mAd96K56r5TFe6yBfDX8IveMzg3Cw/TgXjs9dQam4YzuJUpKF5s3Jazl
5emwCre/OrZN+XKfi52uU4HlQED6rRFRF2F7wTrZ+JLmXXFqQKn/249/W9bEhy1x
xYb1zuI/Xzx1s8puYI2VPvwUg6d4Tpp+IQFr3oF4BtTQq2rFZsfzK8K/zp8UlqTg
sLwrpnhYHUwYCkWW1KIcOaZIYz55ijoJh7gGw8/hTfdSc1H2BgyqWdUD6LdUL0A+
2IKDqrwX8n6h6+cpypIY/Pl0LAoKQsKT3th42wAY98gT2WdX/QgPAA1+BxikLWLy
HhO0KPMoO7tl5Gi10awpSeJRbZXY/38a4q2zlvFfzXBeVTM0TrN2TVar2R1wl1ZR
1p6KuiANSwpxfQ9WgkE/nPAdb2RhxMrHq7mXqAFNq7ZOliHk5L1GXkHz92VHM0Wh
tcuThXRCgyS/oF0QYphTjGxzjutuSF8aL+uu/WJU3JP/2GIRdX9Vk+WT2Q8BPPYO
rmZ7ptP0CpDvCN5WneLAstewARwEHma7fRzlt7UfCEPoQQJ8Z02ZVLQApCJtrHTI
GKnuQzverwh5cdo550nq2axlkcFW6rTQtab3f1291boxzQZd8fG9o1JMvTJDHbkx
DzU1o9i8XmSpBwtxyy8R9I1ZMPLzcPVxFRgWjRpc1HiaOy7xBGR0DmISMfg9VIN+
HAWA20ivofbFWff3VCAgAsOw0eG/SS3RiV7ppMh0y1SnZZWze9rYqaQypqtECv4p
EUch3qL5reLRjR6BaVsJiwGHUhQTYRZDVKnHTKsN+PM6TeFGxFowXM66EWea1hHH
7vwnvMBbf+Wdxdkb949paOKtmauA73Zi/6QHSdLnPPkGvW+6RNvTgKCa/bsfystY
ruEBmPd1UVsrethh7OMHnKp2+Oamnd8jwt0rdFIKriZvO14DAJoSsXoBWDIMhhKY
079RMY6c9Gpw8GxBTVDDLe3Rkah1BUPcZYV59BDlyhfqMj+hTkW2vh4PAhOqklmL
w/DOJLnJHgAJvagK8RGEZw0CM2kjtArhtVV8xJsEwTQ85qQRfvmh4EdBiskkPfUV
zt5kMr3TkUqToEC96pldq5OOR2gcLsYCULmACOwXdDZlRqJUjVfsxyoD2oAnWTNA
yu/qqErzipnMIyDwHGbqsL23F7ESgtW+1jVhixDS/EfL/GxQA/q/bVjH88OQP78c
xQEvdXZwjYii00YyfbGFptr30nINn7UGUbZUddWskCDkw99ooNVdE3OHwS3IICUa
TScA0tLn9jU/0bEmDiqYOkvSFrbmsJa4TZzxdNqbBT38ULkDLWEjt8kXK3angpZ7
vnCqTm9IksCVZ/C31SXc0FLSA7ftn+bco/LRwPkZzxW+n2W72upfiDqwr7fqsfWd
qh9SBKv5Cm+HEt0BEMw29pyHk1hc1T0MEd7WSr3wu4YT+8aEWxnE65cdsUtsSwVi
2Y26ha2BZGRt5yi28iRuC0xfPcKYhf0aKUptXT2QwKpaMW+44YO8iBmokax1KIT8
y2rnI8+BavlnbY3ipaFuMb6swy6zwUDB1fuoqXZLPOqUAszpGoJkKKP21B76WGKM
IaxEXl5IMRuEVzkVj459MNoEr/H109Kz75IBiNrYMArX0IHHRArL+xfpL3Z+pMg/
MDqZs8Abmb/r30zknNLtl6H1LpoY5TLv+QIeiJ4AePPGJH6yMNpEX/YFNj5Tqq93
2mroh4SQwTSo5KAeIoeuNhb/gKP2fc5fiEdeGjcJrvPt6FNcW9R62yXCmEzPQfaR
Pg2EfW8JDbYJCt3AWfzNHRuChTePAFqMcazhtH0VVXEl+6ea1t5Bq68C8IJUMBdu
bSdBxAzgXP7tG2hzbX05HN/CxUQ2KJosu7mOWqLifDjN96bsZ9FWnrR+mknbdHpJ
zv1E3E4zjo9mQOw9XrVCuv3QG3WSmvT/zY2aHzRg78kCJH07/91B34xN4iVKMae3
93g9MAFQEcZx+WzB37Q7MXyuF1gb8G2V52UQckdQinYbvYrqCu0bcS2fzGnX/isR
c7YdTlrOSRrENzwMigM4bnlv3p2z+uxEwnU8WsFfQJrZEHtkc2rOeakebj8xoZE8
ZlYZGQbRK3lfLqE4jralGGFyA5JkgW0vJNPGjMbVMydGKtGQAUHtnUIS/B3YBxJI
equ3ellbLMIJfVVEpPocN/YuFkvBkGwZsH9yjF252lcRN0duGupCwAVbvklFXDd/
so2is9rvVAnZwdAkV+Kgnv2FNbuov17N57o7pbxbs/KRdbEhmitBDszs9uLh2wfJ
zCQX5lfTdbV1t7ldrEOCpVip06yPJJYHZz4/e/Iwh1M5obE5xkUkFTd/trIUimwZ
avB4dZFPZ9HMluQ4pmrP5Wqp4U5d+m4LPgqckBYqdb9YY1YetrDkGLckfEstcxwc
TiihDJQb9Uz1F/FHkLoHZSAarZUC8Cctq2d2pNPo7LQ5mY2+qrgtR+CIvHf9SWMT
ZipPlOibVi32kkVlCet+xAcBaPpB3JLlA9ycAxPmlJyukKKMqh8vSWbxLeapeRZB
JluYdVBR9WbZ/Qjmyj2UkIXDPay0TFl/UPBJ7iyFNk1ogKW6YlQt7IRdAc3tPWzh
2xXccZiaVJPb1OXx4FEdprhZUtyO7yLuLglyz3+ksf0b1HVkb9HFbSElyexA7vEL
Su99d5laQ44+6wR5uwPAW1q2kMJi+ZgjAfbodfi21hkhRSWjw2JCjwAzXs9qxKTx
qsDxPdSrfj8nBtRPku5uPBS++4QGr2NgFtLal2U4ig8tPXLMaUom3vGx//N4Cfve
JZA2i5Q3eL1H+1XaRg/EYZ9erCagdfknL0KuEjjnCv8PcYSgoXMRDKh1yZ41jz6Z
EzHMDn+7TtKewK8kHZYWIjraO0mcAlsbDg+xxywICyL5lOMjpet898vlwRbfgNOn
bTQPgdOsDogRXQkdHoAAixg7YKMkdOGsZinSCn3iH8GLXvno6W9SgQ9HjA13XilT
a4G5zBYAihwDCa4RNR/y/Ygc1Tzvgqd/fUPD2CldqvD+62yAJ4yDsSgCi2vnWk4C
ur7GDDbgKa4hBwO9o3pz5iZpZgCahNMGckhDoSi87vmpF55ZzBjD3t1iT1SwDMzF
BsJa9k/ULpUypc5szlTWRkzHo0sSdckTH35KtksusfwCdSJECib4eBY/3cdptOg5
JoUeGMayBgM6tz8IXt6C6AanCZHdSvDwapjyM6Z8NHrqWzMMg4+cEz71s8L6AdVr
elJcWEpXtTT6fflTdgPdQACj3NqeN0ZUSIHBnkfXuCBtezNIK8bSccsCEtqgIxI2
PdBpe33E04J4NZRnzPr25itX3J6hi2QKDk3cdlnfyH2xs6z306aBQMU2082P0jXA
BORC9rPV8pkmsE38hhyaLhZ4YaGwmYNR5eaJfli/4WhYe5zArjDr0m4NAlSAcdRE
AbQZhQzuEzi5QGQSDigjLXLNiUs6rmUPvh9t9qMm4DPVgqfWk0LdvoCJUePeuRYF
pW2/FpJ2MeJSRkdd3IOznUTXyfz50Fqv0h8URoLukQcaj/koznGfRVXPsKO1NMNd
g7zIgGEXnq2D+6ZagC/esKP1jb4hclE+ng7RDmpBmrV/eacKmJDzZyUmeJsEUPY8
rYsP37/0U0mAofaJ+BpvxRO4q6OuedEJ/v7KAy+qnlvI9kvJl/3cd3MABdRs/VVj
9iklltWCu++uLfheqQ2ayQiMLFsh5y9opiCxm0KDGUKqzDjdvqUcp36kuuAz3FdC
zsENtbzuaKhZXD2DNE6tM2gClIc5quSeilvF9D5pPpQ2av8dbtJ0/wMH6BgBlsFK
P9fGqcs3eANZN95qMWYUDDkbI2uv2c+vrSowqnrWcucTV8lBoZv+lXWNwgFmgfMc
8sdsuu/f+RzyDgUPeszmczstSlCLE1P0KwRERDv9YNDVnjkoNOY62Ejfa840p8uM
O47TrDQkDMDVLrNQjgSeRDfVeAU2GQ9ohL5GUcH/Dgz5OhYmOI/zWPB0NRlCy62m
BcbwXGs5fdqHzODku+AtVl+bvGdVHrgcFz8xdhndEAlKLTN/CT3lq3uxMhOo32cx
4G4ZCEx0m9d/zEPeJyhpAj2+8OPbofvpL41gxTu8wbs0AQgfjexcei0xgj5T7dXS
lwklF0DtDQ1dWPO7zLTqevlFRBHM2I9x8pyejIUNenwSBO8LHLTFq520XPnJtQc6
azvYE0xSash20NbKZxLPE+s1VmdQ549nIp7nelIoGP6I6E0LFMzNJopEuR5DpU4q
T9PBGAw6kKUs6URlx8ynX3+5dJWs3o4+SF14w2FRM0GmDT2cOH3X/ZeRTvBUqW6V
Qs+iW4J9fjsTUdf0/mtBuE/WGT5kdx/Y99CL50P6aOiNocX7+he03qdrLsDjiynT
k7HumVapgMFGFGQVEbG1ivxr4ZO+mZomTYCClUXOZgwpFCMW3hl3hz4YILkfWT1q
DQIJ8frVbzVZyKVisz8CDnu5LDyfPcXQsR8rFvchAoG8XWIkFWppOLhSX3gdiY8+
FPgN05zN1/uxy4zWF0vsG0gSSdbY86kKKcfuMbf33UkYHzYUhDUiQXvzCsNBAKdy
SOcI3npBjoPH1+lqTA7IMNdNjLCDqSCjAu1/R6Dk6E+svRVoLRfRRz2jTDqFwm9+
SzLVD5SrdZ3iZhZJksJD7Dxoep9PGiK+7X6nlGXyqRudKWSp6WmTDIruESsCHCRM
UiaFDHw32YZEeTQmNNiQO6qMOeMz65VTQr7VUfnyY/XJpyhGOo/NQf1KQUZjHHfX
lfQx0WfpPunl4acPjgW3SUJzR9TqPg+B2rXsRpgMcZoZe6nvJNGyn4sXRjbnAZqE
M6JeTuO3ZqUhbab9nzAbsDvVREnVmwmdxdo2za5MCUpLflTnoH3tcOqsa/wpd/fP
R3J03M7blMJAxrhiCpz+LnGOlxrEF8qH4iTdAMe6SSLKLyvO3uIy8qbCNxtyAcPk
cXHnbp1PuBJzbFTATI2gov+jOgTkmmB/8vjQjsG3N9OuEOgQi90sQhs83Iqw6jGf
1MHJ+P1lm5l7WJ3tR54B5Xqvrjx087bIqbEjgtSVgSD98edJw9FzGMgNbRDcdImx
71dCbyI0+KRSShRhM6jvb1mWnob+THBtDcHMgxerc6O7CU9+PO9yAooD7QkPzqGA
EzgmNImRgReN3c1njQzIVjKdTfQ1pvsj3UOV9v1DV+HSqOZ+3z0SdytvEXOqQwMq
ybS3BnhA75y8dInBXACWRCDxCnLuvhee2VJEy062aHrj3rV6QOCG1Vo4of+90r+9
hrXfrbhtJ/voDlhabaVt7A5I80eKhFYFuBscsDQK0Qzhh7c6LgEhcTWgoHhOP8aJ
wEEX7PFA75B+lDdxdPrj6X1xIlodzDTYGT3gZfHv6meo31zYyVqiHIHkdUKodHMa
fcKqCgdiniVz9J2+9BcyC+IPssl9XzSxZsKST3wEH/sgNjNbTlnjSzgreLQGkad7
Jc7bxKV64O0/JGWxXCP/dJTZ3XiI0RKCbXzJyGv1UvLesGIpJXCSjngZBDSJUgtS
7UffRRmHLU/HGCIx6/kP05Hy8PPUMfQBZdvEfOt2m0HD7SQ2GLx5Bap+VbXF9TF8
nZyxK+YhTbAj5EFcP43nOeHXLlO3Fe86qBCV6Q/6K+9YiRaoBlL39IRiBCylgWzf
dwWNb1Wp9ZjftvsSNJwGm7V+ZHBZS6VJVyK4G/0b3IbHOM8CYKdX0zoJQ+c2GmzF
1bNmGGDfDN9k9cpu765as6RzxrvCVbxUe8njWrIqn7O/4rwGdOH08vjQMP2QvQXr
JCMvRVIOIHL8WTbe22Fi6aU7MNRqWbVUa7hSZ74q6cvW+wjBqva1AmAt2xIR+MyJ
zfrPMhdxX9eMaeQEX3/4CEsFmj3KRVP7iNcekcQ7Ss8O8STK2kWDh8/OgVcVqfct
dlY0FghtkthA1SZj5KVyfzXTw7vsP000R0kkC8uFcAjaLkjDg3JoE06JJfmuH6u7
wAMlV5+r0v0N7qpqpi2n/i6tMreu4NB+0U8J64EEKFxafiQN0r7rJnBk6fz9DM6z
YtJ5HHmfe/J+hN9DmSSTSjS/zZXNKWx5miSRAhBLftAdDrVouaj1E3kXdFlb9mMN
ycVPJgqWJGLEwTTovvUFyodBOsjisULYFanayRNtmt3muHPH7BCK53e4qHFii+D2
1AZ7tnQHa1YhNa5+9mTzs+rjZNvI8fMoGbKC6O2iRVvssN6tnR0pTM2hSwf/jj+t
HVcFkziQcVDJXrtExoYwCNmMNYVS+6cNuTNVcLA04eb0Hm45h0x/1ftD3cOu/rRX
kZpRDTns701RlJt3+95+WGw2nSiwEKhh3vT1/S95qWEDTcjAXhdi8ftSg4zVbV2+
0xAp52UVrQ+hKPe9fQlCWn7w9GzwD3kmeA++efzWzzX+onWKXIA+Ov0PYJxXmag1
AqmaEfLgNj+4Y3F+RBTCzI1nyw1JA2OCQYwgkeOnRP+AXE2pekurYdDsZojyPRyk
kyn+P1VHbDUZCopYpmWdxN5lggq0v7hdC4T/WNe++XzQOkQJb3IdX9UObYjh6PkM
5TvGgdlaqbDCDwL20GKq6Hjsnws9ysRyOX6C8b15sLc6x3NsWfTiyVClm8kJW0yE
bQGDoYvlaX8mBC7WEcPO5xaqsrj/Na+9Ti7bVZxT4aFdmpzd25JUpyUtgKPu5IUQ
WkpwHX3VAx6DJC8YLziOTV/dIITBupBX1lzcVIRUcdEOIlKxirJzy3R+zdAh/Lqn
1hgUl8ndEBlo41HgEfnFmaAxaZRohQbpN0eHcIsr8POEh/xzdbbeiUSK9CBE6GGz
mN8lx/C2Ils2byyIEBNa2ILwjgT02gZtP3hZXIpOYrSHFXBHG55XVgbGy0M/6gYA
Cw/xe7Thyk/5Qfgk8MuWpXJnWF8NfVg5HMejX3EE4vulfupUZ6Bw9xVn+cM+d1ox
tnLhNFKfhvca8XTfcnDXzZ/NsTMRPTkS1XPCXLPO1TYITiOVwe7tgo4r5L//oO+x
yqrjTro60I3yUHJsFkOBha5AayGgNk42+pMCuiQFrIV1VYZJONO2LdtGm4e7Ecx3
C2QwB+Tu1DK8c3Kxg8EHZs2xtCxfpI6+pLSWOlR4werroSjrclU0gs3+n+qA1zMb
0LVFYCJTyvDdrhgcFb78gHiee3FoZDhlrF59oecycLhUsKka163QSQNOi68mWI4m
csxafLmyTLjbrDM8wOzxfWOLQ1vXSyNVJRPavk+8re8zLj1zj519m9qdhN1EU0YT
efl2vQ5mrnsE4CXuQrlqWgA+3Om/X+RbN6g+V6uCrHm/wuS2Cf2e63uzZhHgePGb
HbDvwsHO4vE7WP+9nKyLG0SWLsCS0cDsn9ZqKYNmLXNarcPXpOnOulP+HBDWHAno
VGFKEIXELac2ML1lf1LSXaCYo7QTi7a8+ZBZGHwA7FCJmB5FE02+lI3pBQD2IJSO
gUxYrK6lL5aCwJjm5BUb6WDZjWInFaJIldSbLX9YOoOH/MTtaM6ah5LUhUPEQZoD
6pvF8iIHgjgrJ9tqJW3Ig6m44VgHTl6yqMj/RdPCzIvI+/KoUBaN9hRnGDfZm6qi
0Ok+wN+jvngTLRWZJgkOrXOWju3F+3WXS949UJlL7H0NjGjwA7E5wfDv+zVX0eHb
l2/EcH1eM3eKKyuVUKsFkkVlVGqWaXtWDK8MAjD12u+BFifoZTfmfT92V5DSv1hf
7ygNGKvRKOqm7UCKS5eFVF/Vb+4Eo9yaDeSrjFacRV9/4l35r7dq5H5csFf+wapA
Uwh/3dNsgw/0GqFbsVg/JpKjPSHin+tHAzbTSjmhwAovkdTLcaSiFu/pzMpasTWq
WEh/4UngAZMIf5CRSnw7KXfIYYLZ+cBGYSEwKlF7t6aNAYqv9zOClESycy/dys8W
tZDL1fGVEBPxdSHeNbT05yiGTb5cVjoUiSqYEFpQeL/P8psGfL1Ta8TbQ0bwFwYO
4NhS1G5tFSa9GI61HOyQYvE/hflLVURMUQdgnt7zXoWHXWsKoWc2dDXNEtzjk4ZR
fbt8BiJkhuC7ujMwgaqHSv5g3a2CgkVIHzvpAoKx0BUibRiMSP5eKEaxXLCUPljn
aVDXf+T75e2dJz76lQRgCnlxCOQRscdYQYjZoDQ2kXiMkyBXNxIA4p+4Eu3Ffu42
WHa2v5kD9cTtGbIrPAIPnBmNfqXZzrNQQXalGqBVuqwA1p88POAqLxalDXxeJM4W
nmc7LzbnUIEAJnXbH5GHTTLqapYrSCqm61KCViNEgoTsqHFt122vRokS+bQ61ZdW
lkUw5fbSScCeAEOHFRKVWLyCoBvxgibL9Y+PvhUZX01B+KFkyipCiYBriJCA/6mz
N2zAnwjuMy2yBysKCuthUJ/LgceCM3NL2NO5NV2XjVj25AHWf2XcYxsfdaQIrOjd
Y9c+TOYMSQ1sS+JTiP/xgjsHL76f2ULSKK00HobjHtl/PB7Bv5Ojb9MhKJwTnZX4
72L9oWQPKbhp9kxMnkLupE6Uz1EdP+SNZ/zyqqVRD4TzTDVQjT0dEJLnLvzjgTGH
R2LbA5TGEZlWv1XeNAzdxGKDHgojFcMCfSaQSj6+sZ1J7u3hkT0SUL8G5C6xE1mt
TRmL05XOIUsWu0JqQOpoGYpXUZgQ5qWh9B/M/BD6LvmBkUye7a3aGjVJ6QQVHEaq
rnru7NqgNtcWRjNvUV55mqo0IRpa3qkKpmWC4MzTNgpx3x7M6fn38CqrMJf9Wfbm
bvYJEd94MXcJGcs0a+VqYmY3cn1/kfw0AQojLHD3Fa/Poa6un/zmaTedU8BuP1Je
soSPJE/DE7gTI/PXqBdT4Vm34rE3/8M8PBWdQ28cNa/ew5xS8D/uIihXICy4y2wu
37HRbM9hFPbnjDIZ5GeHV+n5rXh44bfDhCAg/fvRwYbyuAEMGuVu9gygt5Z//Ymu
Aw9Al4zuL6w3XrT4zsomAGSFhdJNBG0JW3SxR3YtKsYd491rhe9lGTgOfUoEIFFG
iOhoyViRWWo+zzyBvGDHNjlMzLYHDa9+zvh4GFRovboUML8ABbP/NQejsL4ri7XR
avcVC0FBZPx17RB02LxqdngPtb8Bw5AYiBPbQgwkgWk9kpF2HZ5XwSxFDnBZaUBw
5FyzRizTqDEK2/jPkrMOJL3FIiZzVSrWb2FdMWR7WzlapnLE790GUegpyCKLt9Xp
xQGnPX1XpAjlrLcdgIn5KAiO9BHbHj0hZXQQfbpO264HWnQ7LoVNqwdoJneXEK29
788+nDDpJx4xUq9rrc1EwOa3s74AhAUQTxdXU+H5Yhj8qSRNF0aKb4nsdOEKoiYH
jBD9a2qKqKh9CosYitEJOpHmYGtsFejLb2v6yUT0D+jcGKioVktgASJmKnFyKQFk
YG3GbBRwkZDzhMquvUXtF6eVmNiE+Xu3/oWUmEYO4mnClLQwqkDjc029qErrQrz2
ygwHmyupV+dJ2H49JTPTKjrYhHrWlWt5Iiw5dzZVk/5NkyPwo/N9gF8BTckLvubS
pLuDsZV0kXXz+gAVSTUnvRIwfO6oRn/zsqKEr5DfeM+ce5xU6FOb9LkWmHClI2M+
bEm+aurj2a/l3azBktnoBoOsn5zxBhzrrHUCCvQOurhVEFNmZkaWOEQoEhMB1Aqt
fPa4Gilue7RTfOENmaP8eWLUh/u/LkesII5niBOawavQyu0MbcTiF1rxTV0aycSR
eAny7oWzAmUBNkrb/VpMoFOoKUxyOkb1kPTKnoZhP9P0Kth4gwabaok3yfi4K2B8
SBZF9NqL9PdbyK2r6RPnxuBS0tyRbqaQcIWlqorRolse5N9+cRHUx4JSysGGCoAW
MuG0TiYS+Hw/EHybzn+TUUKizYPsX7UfTU//pr+6NgRQ6r9FcEbqG5NkDvUkiAJE
vpFydGNK7vrVhD7p29zUFq5IbAs3kK++tFQIJIoa3fIXwrFWEx5MoC/aYGXKs9h1
fkE95I4q07nkCnkmfRjjVOkboyMgkLeFMrEZRaENxoNa5QrdGK6bosMdAYbeV2U8
GdxED9ecYNbWk0j7ssn83oFHsAYE4bowGjBq1Z9f2+CJWZQp87z99b0hQJNSE8nx
4KKHc7L7DJwnGsE3GmS/z54fSfxOaOa0j375IQdvovpY8CVITzTSDKD5vnsjvEmO
z9O+7OuF4lrpWA+cF+7OBrp+17pYwl0RnnICayAycFx6f0kPo3Wl0acNj0GEBsKu
p00mWVvoM2lWC5+A4JJqss+IikcRbcBDhwwT66IWmf0keVv6G4TN1aetPt7319+/
w+Aqwrs378aK+jwzpRISeiCNdfSpH8kThEQTusAtA39Mj17eJPpQPEC8FweSIK+t
oW/LlHm6Vc60Xu0rwqsO4I37Y89oFO1qsi+vy0ZaE0ONLeM4fiW4NEvCm6na1YSz
JPkOvJFCG+erGKqPKgl/sJ4u9l1O1AjXdzm1XcxuCeSBZYvP24mkE+fhV3SXeoVw
DywyDxDD50b1aPYgHaM01mUvIKZ5UWb6q0kl+aZ56DOyjjuA88SqrbTBYj+T/srP
HhE/qqyWemBIif3qfSLnTrvwdD5EaLkeocEu5G01mYAp8snyQ/kqiyVMhDBYGyr+
n6AZn9a1OhZLMO96dOx6ZH+cAH9f/ZMKPbQYfXZs/giE/fHPOKmrF2m6ybt423ac
xd7DWWT3jM69gQTw9pIDDMd/+spwiz4h0qGxkQuZ1vW10mggXtEHNb9Ea0o1wPpj
X8dF4lZ1TfsDvCYGb4q8TgnucSSlbK4P6TkPr306QCXmBRXnZymbayjg/5oZx4Is
hq/26QGK/7/GCfr4jeKWsvY4HaT7aI3+XFDkpHgp34vFSb1soUtcc99qG8PrfrQc
ixJqdP2R4J/ZCmRUgrSjIDkCdRWp4es6+Jf2v0iP4i16IgdYgBiyLsKMmb+8HSTd
PXIgTHxP1ZstExml+ns7DdTJ672dk6keU9b430WRXXH8ylPu9cw9cX8U133sNGmE
ZIGGhYRuf0j6xkCyh6x/F9FxtCJLFClHbI3JBqFHSrLm6LGBMSlom24XRi537bQh
eaLs04Kd0F6A4TR8WQT13FpzXzMBhHD8jmy6fx+BohngW2OhG7xVs2+ACsdJ5R/r
hUZzVFYYs0rLZuFN55Zsc6RfpxadaRq2FFrX0dN+VmuoRaYLoFrMvHtjOdSwSJ0I
ssb8WQcWZ+ClnYLAQ3qYZky4BnqL7k0cERgFTRPsm9iKF7/VLmVYQgkM/nC8eS4B
uH4uqTfvTy8bPGz0GmJd4tTuMJyfhNdj4WRykht6QF3etUgmW82sDFcU3fNnHAZN
HKYmdk5YMKjAYFYEtDCOMk/mIMfRJm3tO4zhJ/IXwvja+cv10LEDm/xIUYE3Eyfz
d62+7e13MYL3pwBTv55+6jmwBxuQuNdHxi8gTV+B7PkmI9Iw1WtYPIXRH+mVqZqg
n6mf2OIFSB3KKwTYnMoF1MCBRKDE3Xny2PBOsVlloaHSQ07n4h5gfyXJors69URS
kMqVafr0FEwFTpesksNAK9shuu5/hkTxPy9q3UFx8H1viyS5Ft1b3u/C0zRZ8Cbn
1jKte6pZVX0mlS08vJCDkXfZz7jnnDAbC2SnK/HuMeG8fICv0NNAXIowzi2soinS
495+V/ykhhdSpVWS5kSNTJYpnNXBtp4Zw/DsVILAA9/uV6tErQdGGsBUs2Un8C98
43n111e4mtofi3nwUns7W/bPdgulSaQGmalWHdqHRDxqVeBvGXIEiE1Zj6Oi5/Cc
G/wYEIV/gi2EBCum8lEU3IfBGwu2RUnNmswWoq1KrVY7IBOWbrdKYRbzXxe25DwQ
6VdTacwHEVsk8hGzk0agCdCnss8qI2g4651gbCEy5EZI4MZQpYBuFK6PrCsC97od
nWW2Ro09NuhAakVbeRM3aVurZl7zVYEWJ5YmKAJ4ZY7kwIo97Mto/KBI3BaRPrMC
n98HNbIwhu9ygqpRs7ghXOnBDaAs99D4NIsHh0QP9DOy8vhfHfzqJhoISiF9mYbk
/VsKj7GMD3MsMdzvELnCdX88s27phNEd69SPGu0NJjaznt4/RY+8fhLMAJufDxt3
GnuU42cPktKy2q7mtoa6dv+Td4hFBWncfC5DD/2nur5zKpJ4Fj87924H4Wcyhly9
fcAG8o09Tk0km9/p/V6AqX+LUiFJgDjK/G9jHSSYI6N7av0GSjBPhnhkxakQ1F8J
LXxAJ5IwEOMX/B06e6swcqDBIED18/cLfMPpHzqNht1+wT/f2+tet2YXT4ti8QUW
ahC2VSEL7Hk6QUIauop+km0uKPgWkQyboLWhccThglZoae5kGj1FZlQMArIJuJOs
2Z8D4YG6TgrqTlsby/+u6nqFtyHYBScicUAK21XR7i1lJClCgDgtPF/a6VB6VVlp
Hg0uNhAHJpXEwWU88yFwT89ggiTXqmJz+48TvOepapAlgLtyJAvXArc+wo7apowi
wvNmRmBavkfnFlg+yIOXUda0uOeOwF7++YMpDSk3DrdM2Bg5otZwTnakoOIn8tIg
2iewxxyO01agzI0wdwLOEuF0XkhyxrCtQk8yAeke5zTuv0CVasyqBwWwMed5+uwV
QbIQDeB2NngMyuD8y3uMVApAw2mDESeOH074u//KoUlpDMVYWISBRVHG5Qhtf0Qo
VmmiaFUbeQ7QNnlifs7ObMd+F3otzp8yU5iTCKKWglnpHzb6vYy+uwZ56R3GYNvp
0J1O1boc2z+o/Uc+xcG3mx1HM3kCtLbhBdYFmfQw8SUE8VRkx3uefm68jd1QVh77
+s8t139dUMrF+K7wAopJOExagvKgEWo90Q8N+jCKq4WjJiS8KFWBDyc4Ki+A9fCI
NfxM2GtFPTgRQQ5+JuhK33YPL4YuGo+uIDergCcAnwEuFPFrlZnI3q2McbSK2Fk2
XoSh0J9q/em1QpZopzZZ0YXGpjkMd4rBOCs88kcQTuHXxjQlHiUzqKLZ4QdIDJpJ
IpKmRroc/WO59z9ROEZOVEDtb2c/pSsG4JHoKDgLhaVT2vhhT3ezWzRNV1uRyMG0
i1Q9t6OSCpdeNJhdc/CPzg8JBTcpiyjRzmk0z6pGnpBO1J3rBjMmGUQo5V0CrH1B
mi3yGp/Ww2mTmR3OXZkn8URGWiN4I8Rg3rxEEEtc27L0YGUPGeJr6PI0YAqnx6Br
PUMgk8NxiG3vW3CFAJ0aq4pKN0mRFQS/slxeur9QEXecZCZaHZi/QTB1D5ZmIjF0
otjpcb8Rwv9yIcjl2xl7UFm9XW5+DwtaLzr5R+eKbgomL6VQkjkAI5yaQPPqQvT7
0aJmCQi0P13yshr/oWZQ2C5X4Xy4qpM3apE47lgnkZqxz0fd+XnQIlbrdbx7Vhnn
IXybDLLZ3EWkT5O73W/NAHTcS/1Zm38Bt+NtsBkQsDl/+GyE8DXn47O8Hcg5fnS8
KAS+0FHK2SEJvMjcdAnF/YfUEL0P9m1rVuQVAFruOcj4tFb6z3qaDPoBjkhAeimw
rPQqbgQPWgdP0STZiBoU1pSy7JRxg10Tzs7Er+EI3Z6K7GHmj9N/bxx4JoAYP6qK
RLOmbKCsuvo5w5h4xa4Zr5Y1mrK8m5PsKteEt4sV+8+QnKI4vhLm27Fw5EKdKNt/
YdUBuUHkGeQk/q83TJ4MWRoCzyQMd9QIA3/zAC1PZim0ljjAGGcDmJ/cfSAznUkv
FuI1jtZK/jAGW/HBp5w12fPKdY+b3cfE5fGLdEs+xvWdsvIfPH5MUyeYVW/ZIwig
6CC/YZOjkF2mnL5hwAPL/1tC+HP5Zk7+m4PaajP6SvO29xRfSIvTvEwNqm7BcqGR
VRI8vqi1Nf+rQXheduHvRcgPGrDNInriSlvzZFyeWWiwhCsm/ulLwCQ6G+9nwGlo
VbSdGm5BuittGaeCH5xMNCzHGdT9lDbGGGmUtYklTPNrPd3v0G85cbPRVHQHN8h+
OeuG31khIYhTVlMSt93P66+NTI+J22/jvcBCc9cOtSFXBX1HrtVp8F/s4JnEQjXS
DwPCSNAjjjoDKgGrhmsRPvYTl8NwyjVTwu4FoCN9893pzO425YIeC6nRxF827tKk
yPqZqIYdLzyH7t4VRLRvirW3T07hSclM2JLDodZTlbQAZyKcjXgTIXJ2jYqpMfSM
jhTJJURiSrRLmcLRPkC0JKH8vXBlFeoyTRUhAgUqSfVJcIPMq4VdZ+qtcoCcGOoI
GfBcDuk29xAKbe1vwvP4rbluGP931+580KU6MMRkrZ+T1xW8KY5FR5GmGKImMHOX
0O1OwvDmc1yCL0JHl3EXfw1TAmplmoFpTGEJxUCZHW5LpgtY7ecH5IAGCnCcyQMS
aW7+KikPZaWvg/aDkq+OStg+k4s61KtoKfIHAchUucGuMmWZvNSpNNSeZn5GS0fb
X/5VQZbr6/YCVDfRXJ5mX1xfj3LFFz58wpuUBEqOUBuLVP1Lq6wFwXZoUbG+Y0Ku
uJH1nXFfXFRypiNJzj5lXxcWSFEqpsE/10rEVZ7aix9xj2VGaik9whVGv3Yj8F9M
nMZt4JGYf37rlrjxHb1B0yrsey20oArlTfF2pZspyMqq3ELSuZo2DzV4HZ0uWvTi
6/V0MXZs57NVsdsWRmrRPJl19nqVC8PcfeD+MRxeBQ0cgrr63O3LnppRYK3xteRb
+780ZmowbNQlyCgYhZLFq0itw8TR4fqARNzR/speUWErvNdLT2ujeEw3acBv893h
7pWHv40ytZZBuRwRbWNi+CwtAFvBY4S2WrxgtBRc8ssSGjtK1K0Ic2AzuPQ0kuAo
7SzoCIswlj4Bl8hIXWsyEUo9oRypkmQXFdaLk0dxiO+UStoF1LrUsBiNBq/Ypec5
xefKu39oziqhg3BaSPp8xYFZUBgBrzWtMd+acU50agEwG9fIfUwepyIhBGrw2mVM
s7jIvuwbBipWsUFq+oJNZPWmr9kv2lRxr+99wGYUGBscZWkoIbxhbPeEoGRKOZwL
33o87X6zqjxHpAwNcsRUL1qi+XsZKgwQHfjDFhP2yeSepUKk7UzZf+t/oBwA9bYA
mROn2w+JMBL99Hl/z2sqmmWBckBTnUdiGwzsfpJ6oiSiJTxIzk6iKfnzr3a8y8Tf
/l0Gb9Um9OLitF0OxhV2g4ruTODmAcXP1abdwDHZL4lJRp4d+haso/mCYsGPBLSQ
zz18jhwNLDFrqvqq7O5Y0qxKin1mo4zv4sbe/jD9y2JqyBgRVqnVd3b+yNb/HIef
sixgI0fAeXjc984+tSXNVP7CMq2rurrinu/4c2oMEYVAbVOHZ4LGU/8HIS/tuCfn
ZKcDzs0CCbqbZvKy6ySXCt4mB8MA+MOEcQPlUgYVp3/C4AV3N1Wmwy+dLC3mxso6
30MC8LU32WQ3UD0cRCFyx2T3SIhM8sP3Wh1q5DYo1r6mjDoQRMJr3YhbGpVJerBD
6q8SAoyl52w4MUAuUKciFJJliYjIbSQWrITVfHSLwPkBTrIWiXOmTBsv6NhAwvRO
mmC8SjVIsSndH+Ba0qntKZxNOYWooMcr0YRj0Q2ddQozIsSGM4UHX6OHBQ6Mv2HJ
3rSIQYGsnsla89hQ2AtC4yyYDUXC5NlxjkrpWDdsPmqHAjQyhX4EPcbPUJNfp6nH
EgLJJ0a7NLozYOeF3jSakKk3bEIw7v8XIJ4/uOKtWPgssFcLrhTA4WYX5etCEH+a
KaOBgQozcYkAWeOQJ6kicONH0e3VVTLEwNNaIDyAv8v+n6pTp4VBAhu6CXm1j99l
+wmb7C6JRSoSUjkOifXeY9yQDpQU/ujVPXFM8QALN7nMEyw9K9yKkPnDp4xWv2OH
786c8Wqw+Q2a5QX2ICdF3MuK/KSgWvmNagMd+fWcIh3Ytae2ydAAjnabtV36h2Lx
9yNTpbvSAljoA27sdk9tS0/EjsgLiaju27q3VvjtFj9H5Ns62k1CHBnL0h9KYQgF
Y0dkdNUACfQwzkVPbEI966ACTMj6GkGcnh1XwYYrql5yCE6KOhjsdh8WsauxzohY
dgn3qzffSBHqyI5WOf7aFxNDBl3F3GqwLldPkjdeiQzZgpNy7XV1l1Gkd+yf1uYt
fSUEkQ/N7o8bX8+uw3y7alyFqmfFmvNCMLzXKokcSmPzSY2/bM1LVODHDqcaCUQC
f2/wSDDta5GxU49m8ZVyawi6vLINpbdu/p/95nivft+itGup3i7IFgYJISzToJOI
XXo2fo5vXcfBB6fIV2kl8f+mEE/aOoL202cZ7PB6DtFtTQ8bY4bWj/hiMCkgDeXc
bgpr7idQpA1QOM01C0R6I6OT/5Q/gdV9ou7DI5A7Urda8OBso9FTSTvA/2PLTlMe
QCBrkqdT66qfE5IJzpeBDLgVe8NOCDWYgvXchIEgLYUIBi5qtbOZQqiMdyKeBytv
0er3HQ6LtVYpf8LW+/fplDaEP1kMBLzIsWmvU4P4k/cMQSsNawCAFS/MsgXNjsEM
tEdu+Q+/b+9HUVH+Laxk6LttXOw7bmyVGt32Cao90XcLEOPfL4GXoGGSB2fW/4mr
gUnwjWnA4wuskMr/OBbjCJ4wnbTTs7EBv1DYFid9Oi4Ww3Fs3gG2O969AW6Yr/ZS
0oylWZzHJBE/AQAorVDejTRBbllpijAQk0pvnMUWjbDHJ64R9ovRSmXFHJOmgqcx
AibthakaEl+/d9gdF+VKV1wVEfur0VtyBWk4Bcb1hE5YOsUvVzv4lbBNZ1fHZrcA
NzTbodENffk1CUjd+Vf+XPDvRSfWNLS/nXX9t3HpSTCkKV1fDmCSJ5dCZkGkj3G/
2jOcd91R8ytye+NnFqaixEd7iMKV4Fh+pgo5D5NC1D9+9efaxG3anmSGga72lPgm
yGT6gLN1tLWiH995HYOfhC66pLF8gz0doqK+ekmznqvcBm3CFvy6uJGeqmtX1aBI
aLulTh4T4yCeiSZxbiqkbSehF7jiuEu5vflf0NV4LoCLAM4Q2VSBb0xjI14BBSix
rDBAnetRcA9sNIALKSb4vXGDCWDXgA1yrC9aKSI1XS0gW1v9mDvNlEHyqa9vCULL
gr768HoGNKivROwW0gmHhOcodVBtf49FuwFEG8SdbYMvkg04pdhFbb3R/gwyoxmm
hevC7YKQf+knCbZHnCYcf5LZa6yoOzILefzanZB/GL8+IkDxfLZ2Nc66cgIiqQUI
x8uX5bdIqQlxKnCDPehKVKyzVhfU8yLe9B4ba5oNsI9nXKCqQPhm72MWqDjsHbKC
JlmqvVIRg8FSD/ha4h9q+Mnd0EXV3mJ5aUaKEzVG8VHX/bguiBrpjkxj82u214Xt
bv0eBfOibnrDotJsLfYug+ziz3GIg3ti1OpPrMu8eB62pSMdLMpEe3r+mS1fBQ8r
3G+pic766Crt2TxB7nZ4eAPKEWxwOw0RW8oVZV5mIk9SRIm+cerWlTM9AxPaVREn
ZzXp+O2dEDPTXnsq7hP82L0/koEEzCTSt2PjMDxrqNdk73dUV+6ulNOf4YeuRKou
hcMe8AF8yHvxIKrPU7kECCn5cmTfY0HT6ycRGwXuDSr7xP3Ga3QL0XhlGdFy3jMO
iPioMLO5RFDT4vu4os2dwdgMIpZO8p68KRd2hFa2sxCl828ycZAeCEOKV7Ypg1Pe
c4eP+sjKNU24zXZ94tEQySyfrwAyReZvKp1DNLttHkkksBz6wHH40wzebPrwmrwK
JbE9qXyc9ig6ueA5RKtWHg==
`pragma protect end_protected
