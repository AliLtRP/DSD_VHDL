// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CnSChecVN5ugtkxowC4MwdxqKycmHwTaY5qhXreY+Cevf0/fz/Ms/eBb9xFpc0XK
bq4GSh0irTE/Cp4nuo+8UmfhjRfkCncXqGrf/Xfz7ZgjO+TFHqEkL3FLoB2m79Pu
nSCAeTnJCpGh7TUdgFF9HFvqAakfrVOXIjMZZsBGT2Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 86224)
jx4tFg+IF4ALBwl/KChjhi7Rge5Wu6moYq/NEiB8YijxAvmJ/yBctJgxYNqKSbCV
ZwEjkqpFOhqrHk8JVz7MoRYwSTuq0QSZh5ysWKRXE7WNzf4vq+6pECTPMX1uRZkr
hRK5zss6tTNeU12bTgCw7JyNP00in8ObqcW9rENels8uLNfv22NYBDU6Nu0RNJWZ
Zk8P3TW3l4YXz3P0W30UYmxkrzyszO+nNmOKnQEWFhgXzDpbbMHNcD2JdE2PzV4a
Qx6mM2MPPSnun1ZS9Cfbe40+cgd+h0U4Az9GLSMGDxRUtxuVLljS5CL1OqfGGyMY
kkoaHjjNXUybBEQjW149y/vb67uIKT6cUs+7wNclOoSw2nABD/MAyZCkx5d1FJZG
pZb5dxSu1hFZ8g4WOPdh2lrqnqTIPkza6c/GR8HgOVGYyzJzVxRk3/6VVz1++yrK
mAFZIMrcalrYnVAJDVG+H1yem3RnNYT0CmiC1nBz5bfS8BvtH+PSVyGq8Stci11F
IPwTotodv6QY78pCZ8JFGAYiyClo9r4DqyZXJbMBX5DEQdaImHHHO5eukaZM/KJ6
Bnh8hwzy8KoIa99GwalMVCxYIjwEvVYIvrrxcJvjcg05lQt57ejMVDRiJc+f8BDn
WB96BsKqRkdLE3oU6mD2yY6vLQOjiXOgWnlVcdwHX2EgZz9AJ/zmWYhhe/j7+5XE
iStnhjQ/zim0mzSE/jaPxB5qLxfRH6FWJmryj/oFQhMr9ughd2M6mV64ay0I321y
Rl7gbPSSV8AEMM6NAFCqQWkcf8DbeM0xFdGYeuCGjqiGp2oUvna/DNjStu2wvatB
h3gBcq22S73/syuTKPxR0hK6ZEbgVDAyxRf3cKgXvQ4BKQV2ARFEpB72DoEG6rwL
NmCmPFzk9XosbqQXgFiDak0oUC0r7aBO8gELqBAVOwebJKSC7JcmiL/TTeoRXBrH
8XLhWCtkF7ihzMFHRrLSjRZ8OZYvSAGufp/LMoJ7GkIiWRmob6REYhd4wmVOaE0d
zkfX1TzjRx16VsiGlEGwuQtq5icNVE/fY+ZIEU2u+Vx2uNk+W1JY/UF/pgP79+E0
65OSM21JcV+91qilC6dFS2+/vL9Y950uKelxXLFawcuKvSm0De4FFDJgz3UV+W9N
3LfIxtWHcX5QO8Tr5YYxF1BSj0M+MdR6gSj8h1xg7eNpwcuPz3Ot4nJ6xQPPa0jf
ac2jeoEq0b4DslgRnREgvVTG3FAcMjRkhp5fOdNjYp09Nb7TPqlzI7No5C+ZmCZq
sJwgMhV3obZG17X5EmWV0bgxExZXh5kbb8UkQZL7BTubtC66C0YwAR/GFRrM+hhX
8oi62P/cWkvIndCQAyQRYDsJHbAwrevzNwidSe7SoJHtoF3awxU1rwtp13mmd7cw
CAQj2Q0lfaFU2CEB5PhrgfiyD9/wzMDaKdS5JgfDitpDDfBlA6UD+K1jojMVnlTM
BjPeGhst77fmssG9NeS9NRVyaAlqJz4boO8zx/khHLAw6MJwV941w7Ty7Xop77Yc
OgHNviQDky3bhNkQbmZakAymRN68NW2GKeIyjWQGkCP+sUBADPwFt/sUWLO4AMhe
VlVpuk4rnCH6P3UdL+Z8sjsT+/z6yZVKpr1ecbqKFo7jYipgFDCB2Gk7wpYIcbKx
MqGqUD7BVEKDGZXMNcFp2kawm7dnv18hUiKVatI6OamJwcVQTMWpTnK3J8MeTlty
3h8t1XHVM/NHaaVstWvb/vQ5dB8myFakp3wmRYsKzTrU53mFJuOp+hXvrkGwXKdT
AT4fUONo6HbFw/SksYjga07KSdPIoSBylyE+k+zsswblZk0PfpS7/7CSuTlOStAZ
Jf8R+D31RYDPHpXE007fDFX2wVZi22OZdXwFkvM1/4o+lk5BRRt8G6dSbBaEOFGG
H42rKIC0qLdM+iO6MkbkOGDM2WELnwLj3zKO2aZyAMoSeXXsWBZHBC3hF8r4c7Iq
jrWRMTc2NYo9EAMb6MchI7BpksgH1Xcfkn3Pey7+OF4HtaPQKQI+9yLBPmOt5fS1
Rq8M4k1lD5XdAvT74s66Kgcjr+VnqbuFUAY2PeCTCI24Dvs/NhBKyH57lM7DSe/U
xhDkayyZ9nutfsEhuedyYSmCUSkF8uXFjyrG8XTF4X0FSNfRSNDyiPs0UYjkp/Hd
d01x2OAxXsqnJZgo4kWopYkFZq4QUWNwyCGXE9Guw8ipPuF8PLE3d8supVJZsjnM
JNLGebt6uYbl74/idBU3jkKaFXNHShy2rLiU+KycnFPBkaShRP+L3hF9IU2cs6IZ
VlGdU+92DC9ISC0cIBh7AsynMv3xiIeLkbpBN5urvKIEPlkszmhhs9bhCK0MWGuW
Vn/GqeWTEo4VARWSpMzeaf7Auro9Tt0BXdpkdop4JFjjbXxykVInqRWDHYjdo+jY
x7pNVJ5iEs3hwx5dTih7U49HaCSxzFV4aEDfL3mp3956Qs5JtV+IeGuE7Sg+xXLq
v7fwtAycETLNInukzXEoCBUuz/lLCkr9emZHDVCzyvuwGgk4FXr2+5Vh6XkVbDru
6K7drqr33pSyKpo1NDE0oX/uyASUE2ck7MW2bcF1ygtKzpXUQwdiggCaqWeFg0fO
2LKG+6tGFi/RPtGRI0AKVaGXwpFccuWr7v28mSWweiRtTRQH/cF7Mk0axAKtADE5
j+51R+ZLgQ3Qta7xiXQvcvotg0XSA0QQyH76whstGewA+dNlq8yQgAjVpyffu3Cy
6Z2JQJpOJQH4LlolEuUjxnw86TfB7wN2OsAQBJYHpwDkEaKHGOoJcy8njMYpFWrA
8iVrKOa0Saua03C8ES4Wd8XFYIqH2lBhZPg+n1v10a6rvDphv50+zPBC792GQEhe
Nd3qc0E6fxsfl/k+TDZXGQwiFddxmREpJ+WT1dzj8hJkTCaj8tQ4Jsf0wvjAybah
DWEVMSLFwWtxen0TgHo8fLgykAY5bLgbAQDlEf2o8TC1tmLQXyz+xIXepSXWSI+R
+Qawl63/lcQ9Hq8bV/KU67lE0lfmJwTap9lDq9aQ/BpvrLQ6ws7HTR3+w05cK5iy
lormi6TFij5X74nTSF9vyMlfSD5rR8Z4ZYgAqjzEQ1tH0etO+OUNrvE764vTQhIr
2+FN3F9H3tj7bx5/eCnDNOA87YghapHFOYi23qX0lViOLKt8WC1fR+7VqosO/HHY
V6AJ1Tl6DlW6AataXbPQv+iLKA6E0c7KOwvN96Nacq1YxJ2oAghYTETKsc/7x56X
tqsPDMtQFh0En0EpHXDj9thqp3pjBEQEBbjg4q2rjtf4hW4L8/bJNxQITpw1LmpX
58Rwz5jV8KlxyW6qFkW08pw96wW5onm2PvVYqx+IzGaa2CQ9PfqdaCNHFBDNaRAG
fKSwbHJwMktZLmXkMm8t/28ArC9cQHYB0WULHFdLmuizm5HyEBFKrTmzXvh5UcXB
z1hX5VzLlE0QZqjo+FkwiD0T0zgajbg45kmOjkloojRTVcIMGw9zz7UDgFk+DykL
OAL5zrPlBMeX6RkeCJhh2BQEBh4lBN/+7go/lZ5t5uVUQ7UwuW+kJxJKDaYvv5Gf
321I7mrIHyVgJGjJsPtJ77q0nocKgXc7b5kFgYkzeq+HoqvLnyRg4+vs0+MNPuyK
IgkAwOx7zliytfhVBoezxCdfn506DEJLpyPQ0AtfUWWBp+LfI/vGtUdH6Sg1R9eK
IvOFtX5SbQG17IV5pn30pXnc6sMp5bTiyD01ISWA44JsaoTMdF2v23UCMYeKkJ31
57pIloo4h+HIqAkAOI4NZ5287wWHI9tjyFhgkAo8w+TGCWH4uD1Yf5/96ObZZrOo
hmmopaFzGtER8YnSvmQofFJMymmcIoFUPrZ+A7KXEhD/uJi6nMCTrAg1h+9vjzRx
WnXyDjqNL74XHxK3yd+QHO+6EJ2apJvtv7pRQdhs4MZWy3T2RhxdGTKar61BOkqB
XLW3tYAqmy7yeL87UQLUE5vNRFiw4STws3bTmo8p5379isy8Te9hzN9cMYmhFitu
yBoRxxaBoeOfWYNyB5Y6FpGAxaQVg0wzllQVIQnckkjD1noKL385IEiZTKZNVyw0
7yMVIdpkSomoTP1bl+nn2vl1lBawtBoslkgoMuIaO609DwDoHphRCoB4GUi+dOZl
slzWTK/TLs0IiRA9BnBFUCYfJ35gDxgxj14tup27ec1Gc169tnmrjycl9d7LwdWP
I6ufPWUqaGi+WhFm8Jl4G5D6yU9xCNe9BdyeIOcT8ca6Ub6IkHxwfiD1X6aWoSL0
RK+xguvdgA3pgtBXQRUF5wUZbnSYCxQ7QsztWmSbiT/ooHvuNE+XdswCmncPYdF1
1lwgxn1CnNSn3NKuj7X3wRz/7QH5xB+EtwknSStofVg2jTNrptUMekCed4Q+de6X
SlH1fjXrHpmQk/efMK3MsDe9fhx1EDYw6C6VYYRrk43WtPPFER8lzwzNDReTEr3e
IYCa72oK8kFq7WDvo5+mvBT0SAoJ+ncP7OhhDwsLP/L+whcHuKXyawV70dheVSDS
jRuGYUzdjBjrMjRhig2xRUArFG7v1oM4Ch+BzJS1a7yIxfS7RSfHkOTMaMVUy11f
WYQ1Ps80cc93kSvphshiHt9THNkx+Uv7BRXUMKO5K76gnvQC6a6CalJylz7NSJAP
XUKejqB+vBTqk/9e3Fu4J/SVtgt+UgNWnACVmYDAJrvVQfM3r/dgGzErMtoRr6W3
kVDTOipol8AAIUHJgmtGaggyQXuuXF1xI9Qpjq1QEmnzNZapBGOLGEMaXWqnsXcR
4Lm8i6AXEpVzutRUfl212EfzzjjMYPB5buODbQ99/7MwdO9fKAGYCVHxly58zUjn
ODej07Bi9eKoxlwm4+gUGuB3j1lRdZfAjt02Ft9A4VDvj0HuGssVScHoOuhtnEC7
tsATn2Z00wVf/f2zHLtTJH71+6Gr13np7eK75Dxy2rvgu0yOItlK8+Q6qBUaLmAt
AyY8h4bcQSu2kcAzKSWXhA2lDuBRPH3blKm+87ySb+B13iZdg2Dj3mMYHlDQtJgZ
AU1uizADnfKDLO1Hh7o1GWq96WS5gfauNVgsa9asz/UXcu1/Z+zB65QTTIBLCUyR
QyLmgw4D6Q2/RsgLXFt/sGC5caLLvvVtctdwFoBBNAqbQm0xpFyu2TuqpCZipWof
H3y8I6eGIRLmxcyHi8zgzybTB3I7Q2PC0wrRVy/2LoQbMpDX1Jifa4MpIcVDVEKW
lW+K5MXXdF2gjKHXKQuMh6/+qKAp7TocSn59NUbdnnGDq7SvlfzW7xXLjZQSAr6T
mLyPipgGB8ihJr9JG9LUptoXzTERS2Kf17CDCQnz0Kev00y1OLH75xiIlT9kW+u2
xkX9FFhwe+0lyTQ0AjDwyvW2ETKAWaGdrAaJX8fCKNItdZ341wmuP+tdqZSW1zuF
KdPR1+DClmdTwrx6/41FMu2CAcJkl0escHSjjYdwnht8kvfsAFobuwJI3dSCnvt+
epj8lEFc/+BMTDCb3Tiwmg73+nsT3IRshd/oNyI7/OXDEOu9kc6a9ARcJrr80VlE
6BiysYdFvv/DXoSnmLGWRX+YgZGoUEMXxFeEMMHQy+aBzj4cI6hgv4lnJQ5TqzXQ
1tI4GSzgvvgA+JzqYBEcbWXu/PVC1AHMb2Pm8jqkAHvVyO0x5MkbLJxzpRCN72UV
fUOyZYrL+Wb4qznZvQFarp1AACXp/imnRCTPGfnMSV/jOEpQjRnU5JJ2Ao4gErtN
cv1v6sJI5xU15YFU+jHzQwm3g9RZ+kMAmUpzKdONtYmdY6J8SPnNPGrlwuB4WpJq
WyO3MMEgW2Hvq2wRPysuKpTnxT5qbHr256SEyppw67nhZx3/QbA6Gm2e3Ci4sNG/
ReoJbU/q9K8pGPx9JjROWKyZvaBazRtRoJq3InI6CFKMu9oesgp++8e8Sxwq4w2w
EbQ0TTa5bwGjz97pFBZMtegqO9inq1ZWIZYL+DB6mPus04Vtb6IwWk/OzDypbDEA
wzrogh9WetzaORGmx5aO/UMaUCOXINaRre4gj/nguLP22SQpEnVcd4u8mIeswqcg
rm7SduTX7Axh3k6bGk9k8qLfusfwjTrA4P6q7R6zB7NKa3Jyby4a1RXnx2/rwE+b
QmAV255Op+RNE2/9KRali/IQ+09Gsu81fNXiqPB0r6YMVvx1ypjqf77tLB95UUkn
ZXSRh823KrRrci+VQpeyTfyTin6XM9kiJC0wzbsthhISqbdqiM1oqfSA7SZHP7F/
WDbLUY+0V2InwbOZEC6Pv9IUXOrl+NImmVpTELRLve8H7J8cYHYu7wzFzJb1rvNW
mjOcTgNNDcwZD2zEXU7MW5os1bC1a1IMEjS8cOTt5VlTjY9VxXCaEOMm6PFAf7/S
G1iZga12NLnKQe9kE77JpVTrtnrI8cjGj7tey+szAgmUVIfM232xrHJ2ebtge/6y
YqNLTkWbvp0KESvEIT/K7QxuHcwn+74lIWdEZDA+oPTH1SxKQELDasdMo/bRq6yc
8UgheRu9lBXwNEH454hldd7LcsE9VYnw2lX97AGpoEDmhwAGRuw9r2SR0nLtjEUS
I67e6aKmOO/l+puvYJplGbgWdbZnQZS4bnwwjfzKyNWQRsmFx1XuluEyGLIKfrBP
uenwdjAK9QxV4SQVmy+vb2aX4Odc7cXes51XGeVDW7BEZIq1p+5G2yJN4pDHoeAJ
1iY9G7Lz0/uHIr5YyNR93xDE5asNFm+53HlIzdOSGWTMibOswI2q3p2hgroXHiK1
/LYCVMmaxH6JGjeEnr1or1WrZpQN15DNifp6pFdrF9ZaPBifhq+8bebLanJGsXy2
t871gkJUMMLKH0I/OXM5GbqPhd9nvWYL4tz4XQzC45rTJ6GbFpoGefixg5bsiryk
6iLwagK9W56NhwRGvutsEB4WS/hcq9YH4Zove4WLa/HXuy7gBVkuYCUjM8k7Zq8B
e1Z+Nn+5HvJnTuAAbCJ809Ve+LSjzZvNX1oOL4gBO6SMGW/iscBMjavXc/LDv9nu
ZBkDQrUHuEpSOrykTDd0rCCWp0GSEqFd9DNbP7+uYPa8aUaG37UEo/D0NA8xNBk4
snL5CDiGCJ2/MgjhV3SynGiVC0h1YjomcUGvZ/NJ7bgS2qcaEQQencX9FlvWv79v
DlHsFc0JX3pXCURiVLbjnuoSokiwxfR450ckSTQ3zxgOBeGDA0q+lAsPISlQjQ1S
s1U4E1O/9DTtiYVnDP+nWXQBtopAYuNxY4gQhCgR6gg4l7aL9Q4R1SlMTXhL4bDg
WTkBIBTBj8GYB6eNisJ8q+2a8AmKyu7Bty4kpJb4ZxwnOkSE1N6qiJxqf631pBPn
au5fDZ5OelZwEklmRalv1aNMU/TjubhJd4kAaYQ6j3fimE8uVXbzMTcqwge7Xp9S
OQpgNyQj0JJxtGYSbQzt4296l81x9aZf1oSRFdg8cPKZxZMvW/BkH47NL0wgfBOF
XkfmbgSa5/CE2m1I6GtFMQ83n64XW6fENcm+j7nzoQpexO6MB75Q+xqxAWV14x3Q
M9WPVX1Yx23WS/Skf4h0DFiqgc37YUk5QtaLedCZmGOUK6ZDSZgPVEzeQr6hB3dK
YrFrpz+F7hhdxgn6myJ2cvn4JV46wsF3zp584kkVV4TB1vrnvu+4d/kQKhsviPx+
TrOyJVlEkilfQ06uyYPRdodPByln2dowxA+ClAQ4LNozE8Z8Zye6YDHn4Xy4X6d+
7dwFkGekej5C9ISxBPfsnnpUnY1yRY+GmQEm6qeEQndmLsx8/sdfCujffQiDGzHz
GEDguS+D4Klgbw7pkfWQhweb8HWWqO1lGfTo1+hGzNL9UHke6jl4cmnRRLc6G27x
V0UxHgTUS/SwYUs8yjmm7P8RYBHRIyP7VPjE7sX/lLxgGhLGL9TSjEPOwDT+lTFb
heF3rb5CDiMn1Im8ClBwPvbKMPcdZCT6ptP5sD4d4Ad09cdiZ1VvxElG+PDHGYQL
67ki2J7fSYb2watStkeXd1qKBzX1Ze/i0GPQnlxzbGgn9GkmGYOSOlrzd4SvWANj
wG8sgvKYwFhyjyUFL2oH+rTtln9prqHsXfDd2+1TLsfs6hJWjbls8QXnYRSGsNRp
1RjPf4DejQZnq0CKyV3hkXcVfb47tFt4dmOA709Y1chzxTd7BVUUaSetAtqJKqx1
H5eI8bzdJZ8nqude1DawHg8JJySPnUq69h0I6KASaCLQ8r/min3bqjkOc+PGNpbI
yc3HGWeH5Z2rn47s/DNh5YTbOLysrG+IdKeKx42VRWTWlJlDPwx2Hb631wkBNKZn
ScVjMuJwbFFfk4gm0R+FTILzy7Ido0YjvNRgzsSzJdtQF07dsdNuiYWL5a/hfXuR
yvlENJs9a07aSPthX12z6H/DWW4Ze98V+gdKw0PUzsyG30h4ZR/hp01dAhzgTTwq
vgb6KeAaG/HqksR6k5nUCzpeFMqBaN68UfpbaFj+YXSdmcodhvGV0R7USmdUa9g5
ikH9VlK6DfOGv/wNtxixc71+k+76bySSdQr7Leh0gTM1zToI8mQ3hpKl8wGoqZra
F8RQEhFtKV/mbElLDdgfRXq1V9zN/WWhE8ezB4X22QRHQY2Aq94ciLfWLuXCO4uc
mUFQmRL7aPUhm2h7NY7s/5wU3ewgtn3LFOIkBo13hHd1gu1D9PuzEoLQf69Zvp7E
2SMkCgbK4scV3I5LWT79gZvCVoeLe1HxjtQ1KI6Q43me1QnmwQItMblVWZ+yXg5R
YtrCC2WLZFcrUma28NLIALEZoACqX567Y/eWglRJaWVDm6a+QHcR+rqtYHBCsGah
DGRcTNdnCkrYqGrUpM+yWYUnwZKq9aYsP8LJBXNqOxfENyvpc1gXfS+GqTVhor4a
3Lv2180iXgM7oXdQfj7tnDpcngQh+1bjI6XBRYMK58C5CPijoOhVPaVNytbeHQBE
NvDQdp9C4lByPf/x8ZrhZqCEIM5+2BcgZjTDLjp31sdFf+RFR0kAo1TfkQGtMkLo
faOxNLIbivGz9hAlK8UVUsmZxgBB5J1XCBbBqwTO+0PT5NKGUiUFnHohk99r95c9
m6zf4uuC6Q3QN0cnuC9HQC+2jVrBBTmM8jlBctnheLcKvSv+qFc+WVQnBQpBAsMC
tmd6IW/zy/6JKm8sN5AZUxtScYnkbDLwnqiusYfLQy41kxR+qhIM/ljyx2WHm11e
3xfZirAtWtJ5g9ANnul2ts8LnESZaZX/cSowA9CGhK4RC9zTp16eUA3wpFu3oAaN
f1x8yULZb//fPdIkSn8XOIFfTPhx4h7WFj4c8oU63vbHPEw3ayXL6J37HS4OhnCo
sjrdaJbR/e/JenbrP2dxU7exZWJStlfiLAVRl16LDcYBh7rJsq+oTFgQ+B3RI4Nu
dxkaIk/bDesk0QrgVhLAgDBaFndohsRl1ZJrbLE8YiOOY0PG2A7+yqf4q+MjoU0i
PnWOiu3DPIJEf0MMrc1KarU77iD7Lt3kaPp2WKPs3eydPLSFp4mCT2a93E3NIQkc
YTzNkHmh3YDZmvRZ2WDOTFoATM2OM++YILneYfu1+fLOOERM9WLAX88LqmDqXHsO
nOpIi/tQYmbfmf9/S/4OFBoaJt0yNUMym1S0aamlZ3dh5IyGoiM+f+1F2bfAzgSE
BC8/5SZKIXt3n8kfUUlN8uQJrHg8R9xcOFecyIQG2HqKo+QrEd2S7zhzEjorOwqg
j/scN/3OPgZ+Z8sU/BghuiYGHSpktpfT/2bIY1dGfPKas0l36wSQ2fA2IYljAbv7
esc0uWTIObVf3AbQ15/IUofYV70mxOTcKNds7tfqkzEUQZ7bkiI/JFQ5ZgSUQnt1
1VmFJDwfxutcqYyB9I3WnzGGJ6gt0ZFT4t3uJi02vTAM42ZZXz6BXKtPSgnwRm16
lnZ+ZIIbELx81n4GDr//gc6h8dRt62W3fexS4rOWkTpqT84qyUi3KxyolMAjulZG
u2oB+pmljsdRGj3+ggp9b5pTWJPNRE7mtxvg80k9JZGg7qzH8SAFWcZN5syBrRi+
t1qne0SUlHJm42+6jR6jOu0Z8xxuLzqqLX4ByY5UseoFFeb5Kw+NYNf+qq+6Ig6c
+QcI/zKiglLEuxXVyfN16vhaKVq7wQnUhf4rftWAnVzTfn6r9cLfOWv+C5ysDiu0
Aa3BTq0KbHlFlr3CxodQ2zX26VgXufI9vP7L8XEPkVCN92+dQRtfGsLRzYAL9vIP
pOLcbMaWBQkbbaG5r/UWO1SBKI9xE54QPFzFlaYE6ghvkXm2GGaxnYiUTIY4YIyF
2hLRHgWv64nWldo4GO9qpntm/CQB8txoHb5Rdto6r45fqGOa+2LHP2jY5ySu43BP
fMxxkq6hjpX9jKRgJhFc4Ld60/J0W2T+aIfmyyC97ls8tu+OgQOOzDFkAAr3tnJs
LrD9+Fiqk8qdXNEoB2LjvPDGyP7yuWk47fNGy8FL5PxvdtIR7xUeuR07MpAOf8xV
5BYSrKB7hj1c8v7fTVk7U1n+UZpC5pS5uvuKgLXQwzx5DdK547/z6N1ij8SE2MGp
C1yqTRU+6cNYTb6CFOdMkZjMaznwwQnt1aGA/AbPp1evcUtsxY+B6WbUQUR42NGF
nT8G+EZhfCSiYqjmKl4ouOIkoq0hcAjUFNONMrHUTfJ/j+EgInxwApC3kZYxGjDs
544DXisQjLT/uLnVUaKOMAmo0ADOVCSg/CrznDakCAKQB8rrJ82dMDbZrxCvUd2i
MXcZkip12GUEsVJhLHbRx30UJMNvoWb0LmjTlOGSp9sgrQQzdjI0SrQ94wn8IkYv
I6013Z4GroHdbgfHPYNyv1sJOJk4rC4pFisjppCkurTRuOjBc8x46IgGiiW2lEdE
rJeCrRf+lHsadQr2tuPjau7dL00qHJZLBAA3t1GUYztmNdlEBzu32HEPGZlDn6RF
JMa+3hTmxMticVyfj69T71QUDICoTYSfQYhjeqFsTpuRRTN06jIbYDU4kz4/1wpP
Dkq8k9GQIdVwrSSveDZjJ/HOJHRFTRJI13j83nx22knphnzzXWs3pvxfCANb3Fq1
gKf80bH2/+CoFGSODKISGARVPVHokFxzFnadfOPyuzm0+9XxSiCqXC7EB3oNl1W8
9DB7GZWt8SFfhGpDSr55eQOfLNinvFhz/6CkzISvoJV5c9nqp7SdwLfrIs3jnKGM
t5SW2IYuLLFtsxf3bGTiGuspmiQRGE90kbmKC9/rz5Ady0dT1KqH26gj+TkmlPXp
7ZJaHb+yQ1AhDCCcuTDeVFbNyquaHHZcilQ7/OcnmDUqHb6P5dHJsZnrNE+GZ937
I55/WVSg6o9lr3LUtyfd2Ma7Z9QkXByPvGSEhEocBfUn5VFPUFhCMgq2yapAePw3
0gCXNIktInNRINjplUS6e6yQlJ24B9f6zjzzy1lUIlhumB/5NHwwyWdZ/+t0fI69
Dr33Op2xhIB9C+/TVjv5rOs+n0osBbDAUY0CoaZVBaE/wqP/Jmpnk+r+iUQvMrF1
3k/L9fBDXrxhAZ6cXcT71LEMhjtiXuIgGYn981JnUTzCBysntL2KV+K0qSisMq5j
5FootV0xkzUdcD5YGGoufpNN678BnQQ6cl+o/TYNycUH8RvGj4B3FUdSjOaXT0Ug
CVit0J1ApBNosG+EAQ8AW+13GgmGx1xTjhLKYxa3t/+xIphad/zzSffDztVGKluG
WfaW9QXv+aUTp+cbgkTbphvacMEEMhxe6csgxHRWabc9iVU2Gh3sZ4q5i8Ady1wv
jsWYzp61WhG4WKxZ4SJK6fraF0cA97HHbaPSYTnxsJdWGtLABMEHEjFyeZgt4Te/
WDCsiljrHFiqoSArlZsvtuM63HfPXpCvAmtsS30jm+i7ySMgLMUju07ZU2QFjEuP
tl5tbUUEl8kFAqyngpHN5+3O+eXH18c5sHAv+d39jMQUjkQaAmLZf/sfon/DSg7i
jGFMTGcuPpGlMGiveiYznyRHZnCDe1X/emZKYSj7M9x00M4X8Yd+IRoQJi7EoKG5
uYOHDv8oFbDUfn32dJ1wc0eDRp23hDz5v7APEfGEZJxwNUABi+J1WixRCfbgD7SA
mDo1Y6LnY0obpQoMTJnOESZ07cxKWXCVo68N6Elg+rZzlQJXJ6knC4ghDksEX7zp
xom9u+1Ip7m76M7Z/IHq4KYg+dN6BKN62dtPwdWf43MyJ40l6DON+ZivpKk3xRpM
2Afs+AyIjj+piQZbeAAU3FwA+aMiGL9O5fZQBpS4guvTOiuURCsRWPEKn2SlRMA8
ZNs9d3xo0GpCiQ/FkzWvY25hXeQ3xvMNQl+PxtkfHb47MZQYqXkUN34r48FCsuW3
wCfnRqEJt8UP3U1INKcVU6XhzbHBi3BIS0SkYb4RrYoW3KqDmUOUE9gTIve7PFAq
qus39/qQPsMDwNpIZ3mj/bLLTXOuET5wk8C5YLDkhDxuWvTK3JQV0V9J0q8HP+cS
tC0Cogi4yqhelI1v523HkiGili0QqzQVjoPHGSIMq83rvi7M1lkELrV/T9diYG0l
26rHe4M2rCgip/31VCgcwjVZ400g7jRIPTAO5PjFXtOgTSZBQpiW5vgsmHaQkNTW
BOBwQp2DCEWkz8rXOII1fcJpWrc2yDDv7MlNw1um7Jenj7bVsACVLECoD2+ATmE4
3eY6MFEWJe3eRaRS7mxOnwe5N0E6y46q63SIMBPVu4gUUptsT7UJhodrzRFKM1CV
SM7JfOYrBdHtddlCajUq9qN8q3AFZJySbG9ERuOFkBA0IXTyVsZL9YRb8i0D/h2n
V8eFuXfOv8vbSDkUAImcPlIdQ+RW6+T7jhpVl+WFzszgLSe2UAosHPZ3qOH1eCjW
aaGm0Jek5WuH64pUkCUGFFX5VjfZLPjaz+/39cdVVX2a8x0z9T7WKzyBhjw7Zf0Z
mEwXudsjw9K/uZgRUpFaK102VlwHCtC48ZeEtBOk5KdcEHjmYWT8Pkc9JDAbZs9Q
Se8Yy+4dtwsSOcX7Hn75oGOOlv8zbQ+AbJ5dlNPYq+I+IHL/gitwiJ1hD19fys9s
h0r1uytx51Qz28c3CZaCgzue68C5GUJ8POsMUfNn7RizYlxTDrlASLUWaj/xr6x8
LttxAPV3gOOJj73S+K+gm6OkUmTAB+Ueqac6o00yPINnaVLeb7oaD0x94aw1Gmr2
mmpwj1RJ1CR/Giuxswl4gZvskSEV1MQYjENGWxMUQD8pLN4u9Y5msMAxjRXRgj4E
Ux3HL9j4VodZq8d/eF1O3UbermZK8l/JP5KAQzj4lbnaaM55lQnVxuobI45MVgi+
v5YkpcK2vaqc6f2oxnCo1f3T7LtcctEDdThUxJQwkVKahptKH36wyaD0dCPkIqlH
/mWiUhTyo7yD0mMUEcWaKyveOWQaunJ2V4ryEg/6Hm/9L1Bn9vqGsRmMv4BpF9ZQ
uTFstO4LYaCZeUazJ3M2h1U0eJN71Gq/lc8htq2f+gmsJLgx70X5l18Gy5FySEB8
99rp3b/EBeAu1TzRUddNUIr4s7Bv7jdC17FOTBbquXQjg8iHFVcxOookj7+9nSkh
a6yOZQPykg+e1EBAnH/D9eRT0wFYowfKCOlPi97rDZ/9ccyd0wZelK6lGlyse0gW
fmLGpUILzHFttcNKvqXAdDYk4+nl2jtVITm3kcmi2i5COBAgu+woA49/J/iDTLh0
siNdM0vFpnwGr86RnX5sn+vU4sz723Qr1ppYVgZLmfWWuqymby3Xfyr7p0vpOk3F
03kP++I0ypKM//i1i6UMz+9Og+p3zPGx+NgQtiBosK6wk32ORECOshFRcSuyq/Vv
XElJPMXSqV+tLCIys1qLULn0qNXLmt9E6b/Btj7vpOLLNEVxoAfrCNEz/xMmBmGN
5p7VZlE5bfuJRJqDZQad4M4+H7KBxQThr8pcCUFzN9Oah0bY5MMYIbTOrfY2ChRZ
Lb4qYnIiiIpH5Uetu0csvIFG8w67KKqvGTZ5QfIpCpXkXnrSF1nuNG7D3ZfO71b2
G3LUGugw707LtL7tO9n6JSBZLRbjLozW943sA6ucNAKtJIDW5vWJADYB2+dLelgQ
L3wn0zp65bRLvzl1nF7p5txWRlbIJ+kNTdogDMPjRERaKPZu9QCVCcs+HQK4D2wO
+9h2tN2geEfguQyAf8uh1KfUhLC1XVfYZD1O3blPQ/zEfkmK6P3tQwJrndsk+XJ3
We0XMXYt5brTpLUADXf3Q+fI6FmwMVm5y1DupHBeLDy/GbpuHd6yqjgZy0OOoEic
nq5VpPyXGcM9LgvPvb+TOanYcgO+Dy+gPxnkd9IHGR8yiTZfH263rADxxJkbvIs0
k9u70rChcUBGzPAkDBK3+NTz8lwtJ1kGV5yEj4bmChGIcATfZZSRCAk1FgIIBc9l
DHXBoIj61rCgPQoyUmtTetuDGd+S5BGYYnaktjiiOkCXvIBoErPw/xxht8r9+NVx
kSsahjVx6oSSqEuaKVS3uMy5arqtaijkljW3qHZyFyZ1cHXTAtsaWesc3P47PBPs
I8YeQthofpa3+IQNQKifVXZuxrMTUKuavscd/l3IX6LmxJ9yWLdvrrgYa4cGU8Cp
w1BpvOO3cdFe3ynTWMeW/igRlAmMJoBeMTCsbKYas7i0HfP1gIgAJufFa6NKzFCx
add+GzI9rNvoYvjmF5cqrDXSlv6OD/kXTg2xM723vybOAt8J7z0Np9bQExHXUF9J
MpAIDvnLGdFhlegWTVyDPTz7ZBd1bPyfxsOGvM+xlddytAMGjvLmAROixc3F3AZx
nreDwbTMwDd5HQ1a3tTbvjAuV+55TJo1rdZ2FR++kroukal06gWDK++uAle4/beM
EGJ5IoVn3l8dOWOVtO+SBOi2xgHcPiODTcUx1CppYtwfa26rO3mZQUHy8Fqb1n38
urVLO5XbMUWtlO8tLNTtb27cSJ1tj7MN61x5SPV1pWRiPYz8vW0FxVxOS4gYzwGk
/Wu6sxDMUlUfBLd37Cp20WQlOKCS2nsjMLj9GfwXVHktrgbRbBT2Ix9dfC6hsdKF
81Gr/Trn1IIbDjpMoSPR+T4kaKABz5TKnPVKyr9SdHPysRnZa3EAbxW1G3JJJB1i
j2tp7n7etdGjeoSdJZFbXCbOPhVuj05xPcHxmneTyDOFy2Iy4tIewMkAI4DiigcL
dMSp4yfQ8KOgo97nWxHL0yrELNUWa+eJ1xa+h2SQXJlufq9LddWlu9HByNkysgYH
DoZvDW/HRtmaIgIiBZbDx5j8z8K1DSsOmUjK3R9R+jpY/A8rWBOwVzFM13xW0Jwk
Qdvzl79U5o4+IanjphCOJNqOOVs9eSdQfbO1NPF2iIL0TFaQetxoENWfc0x0FfEz
IF7ahPKLyR2Vym1iQRIkpMqq0Qg9LUC8H7uSwr3lI1v4k1FksbzpK8ebfQWw+ZB8
x6yw8oNR9hSmPMY1BmH8I04cHldpHfLUIMpk2bfsJOgq7OyyymQ//Myb8yT7fRIW
abfUrf8uJ8MCyFgi3s0HIrsDtgKHhke8f6F+cuI1Ei3YXaI2Xhud8HRCaJTR99u4
sy2Z8etkb9qZr4ynr7DD1yiZfzxRfKPOUsX5xc5TsG6oBLBzWc8jbTyo90WF+C4e
WpzCQCzfj4U5shtgsjQZTlyNJjPpbqiBnRFMxPuJ6pPnjFZYAh1rYL8YOe7OgztB
34Yzaiv+R4IN5VjbrvMHu2O13Jxf5q/4h2hf7hydDNfkSQDc+CU1J6Svy4CLG9a6
3ZS1UF5WoP6zEJAargUT77WmOLOPAt3bGlJX1coE5PN5MfHXzRanac/hyX4/f3Z+
1Dol7OUssy8dCp7mUKabAI72MVKfnup0OQF7cB7BXEHPLQqGKNcku5T7+b7Duazv
QuV4hdOowXxWEqSZYyZpz+RD6sLT/BYhN082qpBAIfa1VDZ5wUvm9Vv3UhIPA2y5
au0CA12QK0KetULDbvJWAHilZ7TGtKnMPtxIJAstWtrisqc2UCmxuZLSRTnS4Ell
2w4qr7j33AjJgga/34Jd0E/W0nud3/LJC4wc+cXZwc32AQZgxoTlrOz8kJeRLdf3
O6JARlqIiQxqk7dLieJCA7my+boynS/ND1rgJ/yZD785+UUeVrQQNXvdDiklTf7F
wmZEx0gDstctS9wICs18WSekNZ9isiQbXdjoszvsnQGs1v0Bmo4VY971OHlKkYqj
SAX27WZ6yLfTbh52+nbBCprSQNZ3Wa0YOkQq3qI0X0E0G4Djy/N5qBLjXPG5Trrn
khMttuCPptPGkSXneBrVu6jCDVkzmAd2KL4U3kCToTUckfNfA0/Nn729H8qiALWR
i46SaszQbGJxrgP+92Sq7jxWx2pc7W2MBS75APGai64CKWPNvAXMzkA4mG8ZXZeW
15EEsCY7/p2IupT+pyGj8yTBx5xbip6Pm6Ga7Zqql5aQ1ucDctTHGrUpF2kR3/x+
nYnOJu6Z9Gc4drfENuuPMMqp5dPrvPB4CTymUfJ0IGY53rXYByfXBnK4QpKPuBx3
3jP8Va2Pv2tKCnRnrolUURDFScq0VoQugHHJGC/V63IBGJKK0cRbk4uhbQve636V
M+9+6TfrkAYAbWEHBTfmBBmoRz2f5jB5kdR/tDjtuneZQjevY+MheP7oYm9h+VdO
R84UIiZKlq/HxbK87mdHsoGwMc+l8vLFeKYGhZWhKvUZsOrJKXr71P4iim01OkSr
FVcOPbu7dkrZ3R99Qm20bHN+e9+hvE5h0uKP29EGI1EkNMNVyi8F0BDmu+TkXLPX
k/9eU+oSd/WxH3XZJr0YxNaB7hDHzfOXHnTUyBBPPRoFDPVmBDrzhdygg/3tSW+y
h/lX7kjHl3NHwyii0Tb05hEhtBXfRBJFDSoLnBsGO1Eq14Y+1Y5oI7WndCQtqWKM
eD8Aeiuhjrq7ELJttmVtsQJAPTDpGkGHA4G/TQsOcOU/nxsDstL991BlcwjcRiwT
jjvls0LJvXiJ2vFe12VRop9tPH7xiFvm4yAbBv3anfB0T98h3h24SS60Zvvz66/w
b6NkRElWoVZgVOwKQ8l6xokQYlJ/dEKPGvUrAwSpJZGShLr7pWxUojwMTS11Tz4T
TZr5MwlzDUct0/au3qSkUx/llyoq1mRHujsj36+O2+pcWeyiLA3f5gEhrAYk6HN1
8p6J2OG+PuW6ghLYFuBMpg4534wFswJfdOHGAoHlrxiLzqY1PKxfyXAwWgQxSu6l
LO5REXSdcJO/dvH2xGDsGAn/hWXTAupIFHnBUxkMMT4sB0USpzfyvFJuPksvlA4Y
ELFlGMhmh9RTJZ/Fc5uDsAGhFsJ/bWQVeXDOH0Lm+drJLT6bRdxs7FeWb4XqsXTP
eii+YmwlFW7xEoeRr7LBdVzXRBY0hBXwblFTqV4/hvCQIBlDqCEY02uSLSauMNRu
xj74fkHfafydk1L+Y306vunX/I/LDQ587O3jLouHBUFi7n+GkPG3k4CYTFIz01Xj
08WZC1BBWLoM6SAvRLIhNReGJESxoEFy7WWWEfznqB46gi9TvtkQi0FSTpPP3gGm
P0UBYOTJWVLkg1Uxyu+DGgNLARVeebe5HaSemPRTQIq5n70fudpJYNWz+YRCgoEn
SA72vn5ixfe7CryMMAMD3CsVV21JdneSTUKD0KbPz9mPgc3NVYx2Nt876IWJE/69
jxujk8mr10QCTiaQJjLcARatZiGn+QrWfc118Emz8MHK4X0BAJ6VJhPJb7YAYc7/
zw/dEJg0m4hTgiLo6mwFyZksCWpQpjwt+aypbusGKTcTSBIJkm39I1bM+vNl4x4r
UqDuCQUdSPrwx3GA+gtkCil6OW0T/GoEcfaivjj6SdKoWBe4TuXWHEmzGZW++7jP
gZgTrGPFE/xzK36AG87NAWcubTxAyFYSDHyjK1l3zU145dYARQnhhzq/oP/A8KVd
Viygo/jssLWjoYujHmyfvwTzQKxrWpZR5+KzNkEdIy/GrkVRzzBXWo033v+MbMlG
G6eLUdj40r3lPT+xc5ERNi7+G+20g40Fv7SiAaPZPtxvD6TV0iVzAzBe952mC6hn
hxw6IWZ7QVeFY25uv4aCoYgXe9G/jKbHVXGC7eVLTcvzL/5M9jJyhGnPT3P6z1Za
xldnNqGrgtwBCHnQlnzM9uRH/Q1UmmGuZwhe/cOKOw5rxD1+K5O6T+bc+1/iyZEN
NlG6MzrcDyP+s/SSyKTtm7JOSsuwhAHYIvipmL/TB/iMAxIkCFiPT3k851er5n4B
dtxbbd5LK0z37RbDg1druyQWkqeKpz0qe+/ZW9aXQG2YBvbuZtFOyL1as6AC5Cg0
yq/EZIcIv/p6duOdFyC1EB3+5ZuN71XIeUqbs/NLBEdtvk7KvXpzNOIkK/6kbSE8
qR9KJZ8yZnkZGYJPVmQZU0tHeTYB+HAIopDbMwaLzY6aDO6d5qL+cL6mrV/lUXcn
IUmF6LXOL7RdbqR3gtrU5uxM6y/PGo+53UC7ObLxs22PtTROeNw/rNitpw/iHaYr
LTKfi6s5tGZ0fJtgdQbiW+qSpeYLLts+fGXloyoOdws2QqrSA8D58Um48k40D4SL
+S7URDkzIWiER6bKJJebcytwWCC0teSoR24xgohvoWuVTgJH+WKLV8L/x83qWXxR
ZmBiG5TUltdT2XxuIazZ/BcC/gcSDG0dnJ1RjUAapAZDZMiPJA+AnLpNdxF95qTU
f9W+MNLMHNl7Hk2HJUTmGbxcpqAIFutwTciGSzva2x2Xhnpei0+6Mn3duHUwnKpa
6vLRjHxO8cW0s+t6ztWaf1mVWKEDLOqGt0FfjtVgoVuXeMVnbi9+7/bM4iqIL4W3
8yf7sjgHTGxbc8Q6ysXOCRzdHwDX7UWERnVd7l/AZVPp9AuTFtJUl7sSEhrBM7U0
aE2BHcj0Eo3DGJQCrFy7b5OSs9Mst25VgEKT1r9uueTc3XywT7eFwcTXFmK2bKiZ
Uog/Ic4UPDSnO64mbnpRu4GbuoikkyDrTzQfr6+gsHK8rjSTHqf3ujkC18u7o0mQ
XDKmNbnP1vGyu3SmJdKYXPJ+D2w0Hr+XBN5aJeewt15A9ntZ4hSYEUKWaDZGXCj7
vA94IxVm2pO/R++KyOY6UYSEeprh3Rd+UagXK8vhihZXyC/1fJHBF1EQYat/H5v2
Djyl6IoplJe4vrhCDhJnrlJwblPrs4+4O8sFazy2mPxL54tQ3Cffs2oBCY/zWy1j
zDGrCYczce/RhY+36K4uu2jeJp6L92P3Zu7wTtHw/sSEkx71TQrZD3WnBDwIGt/0
p3FA2HPfNVVPURE4vpJjNIzj6kB4INgCSnYtN3XnSMHgk4bsXCqY55xONntCbVgb
5Uv3cX5SVApSCbtqNssq95euUczq7Bl81ewKsuRo4nsfVQBDW503m+NSvpdyTIU7
KLW8qXkA4e+F0wESXSD6SXffv9Htik9ohjNmJBD+g2yRFoJG0WMAv3NgTq1YiYcA
aSSzGWsEN7g1+nExq6qzMMmvv7plkcvhOuS3EZjwqMCXnOH6MR1BkJGmeFrJxdWi
+JbGTb++FMvvZigAihk++U96vXaxtZxbtoceKcWmvhA9mZPiU46vN7QffGh11krC
3MZdyyTogGxVXEHzfByOcnCmwkOp+IZjxlpnUpcFE1kqZwZ88N6rcESj9xG7FhBy
Pn5kmE3VaE2h6O7y7zMcan4NAuU7oBRNqq8OXXXWeCgTaHJT3TtgCboBNJrEYhUX
mjLJ6RqSYak2RpnHqRJaUPxiu8aM3LbTUieFn+4XmmLMQzoQytsa53dUqRTobaLP
aYLI7p0S3vLmc4WdpZP1w7NQlh+0G0T0cIW9H8h5zI6LQYWO4mi04FnUmJfMVzY9
qWQfVpNhsVl7LImtM+4DppBvcz0npRPebc1pBLWLoyLdklFL0bKnR01f+k3X+A1G
p3bAD3fXr4yzy1HSdcQxFkH5pKWi8QFOhqWup8mt/0d//j0xLCM6dBoKtS8pyeNm
4WWBCsaN/Tqc+4FykgxQmpPn/Fs390xzBt1ocEn/UpMCJ59cQuqRu8bPgLneaz59
VfmAziAynYBhCvPLmcOpb5cJl6wC+oigFqxKp5yGG0FZX0HFfOr4htspNczL50/l
N73V+4FLsXO//oQ/N2/W+pQEVn5m9uuQGQxqEu2CWSzuBHSbZ479cFVK0lkYcA63
zeZdBvnyq2tIuEmM008BRUUQgWM7ZUXWNBpdN9jKVjPzfdfv0N2quA0SRnHAbO5C
HmmpsLk9WH6ZL2TnRyZzuOKR95hciYTbLrwG/U6j9u0i1EJV7LqU+kvpzzKJpVIv
7Qcx/Vktwd+5W1zun9jsfQfgSR2+DrL/9sY9sqEY112QgEqgI4tG1mVxYpp2t+vg
SjujFzMqEY6CMxdI+ZxQ4ff9EN1MkQBfFQ+E2KN7CtQp1Pu61epme3+CAgLJ8+Io
aVLB/aYTWeuX/z9K7n91OXanvhWzS8J4Zm+VBgq77Mo3fMopq360Ye3hPoBbREvT
1gA/FwWyG9112C41tmxGeZnhTjmD1i7NN9GbGx66LdU2baoaKnzDMK8MYkRWUQ2M
R7sjOM+hEVY+Lb2Hs9eWt0wo7yKaZxDlzxRN0lhCL4dRK2eKE0W6jGz9zRwrcePY
m/HUievUE4iOg+6jZ00A2UnjTlNSyVXmI6rx2LOC0gnj6dwLcUHoe9/2Fd54BZ5Z
4+CxYXGmfb8EAsQyLlVhSo+hfYL1zmYSfvrZW/QCte1Vn7omu6Qmz++FOteuAyWK
nvK1mfVKLGmZDqyZjii22DQkUrcrAZb7e3f4NAMdqtPb37InjBOMnZJJfU3JnyQx
558njKrTB6O0wCLx468lpmDkCKsYjpJEo3yzBzRNX4hrQxnCPezy5irwM7Svpqnj
Fy/FHWK8i7Sj5Y9JQy+9g7QAC3lCFG6FkbAAw3uOpZ4khaPGr67uAcG8d+ZjtIHr
Fw2Ow8IPh63NLHXwxgUuLYX+oKSEiRCfd2wrhmbtRkgkt5nL4B5k2RVZRW0dc8YG
574nykvfOyWJoDkZzjCVjlB4LQtyIFWxTrTGUYBHotcAFcAE9RqWzMV/C/XZLsmT
2EqTy6ST6K3CEGjLlr8NTD2ZVz0ikTmoLrhGTCsBX1FUgSWU9t7eeT6KzhmzXdMA
Pf8ZSTu0fDmmuw3Zsz58bZ0pVAzEOO3PutcNvy6aLf9gQNdVYLs7V+3OmMvWEODZ
Om2BwVcGFn5MqBw4gL+f4j6f0TwEHJmi4fyKgFvlYsLH8tvtugBRc32BrUBEtK/U
htT3MCx5/vFdJ9lFdrXXSrfBVJyMz8oXk5g1151geexa/4GLHGnO9p0CT4oiwFag
G5kg++hsCPnDsjhiYc5GXm/IoTRPISfWm5L9+2Rbzdc9e1UqSylDi2qN6OVb3Jnx
Lqq8D70BYUscQ2e9bcNxyV8+ct6BM/upTVTYHD3Ygf++h3gAldTewebWu1gi2zst
HNKCQmuHZYWJsRyiQ+41bjVK38zsuFVKuBXQstl+O97L0gTqpYW+E2CNU28XdWSC
kXL6Ml6Sihd46LhDb1V8Ezzr/9DhjK790LPGMTTqCs7kMWr+F1dWz+ZpxEB0BGLO
lp6UVC089Cfra+Jh5SRmvLR/OV9fiPrlosQV8NccsxP7ue5mpEONqRmWuxK4VHsl
EckDJr4R8IziBM9zPseLsgGu3S8Jv8q9fyHVy8hyWq3WV3fXfirkl2Ky3yjKsvJY
3b360EXkgGUQVii2rbzrVJuMOt2ODSZY8qghPnzS92WItwleJnnvlUg2O26PGzvr
AtqvE+k2R+Aaus6wGLGVn478ilAwbzux58QK4ytvIuvONlZixQbOAlmb0wW0p0mH
Nsc0KM5IMgD5H/aS2f7wOEtTewFtenLdtPCmLb4drM+4k7QSR1f+v3cMVFXl5fZh
hCL59IzKF1R3W/npg64N9caKguaMEhruxKWEPqAiQFoQMq7z2HmxxL8yEo1L4Qky
73+JPGKaTtUePYjQ7sx8cBqMVNx+tbFubx9AdCY4mKzg084BaiwUYb3eTwcDmqk+
H85olgmMHcTUXJ/WcqxDLADTOluzPumFkKUhRyST0oZDQMKMntshH7fZ9uWeMLad
yGfdyrsFeDhPt4KjueoKxSG96mjGKjbmhFt14lMd96BBq7vkpNpsjKE0oqleDddm
/5AvFLyouqJumld8pgcA2yLl6QwwjiPsdNYk4kn4Jz8ptF72A+Fivulmcvw95TDv
5wnr4TcSKj6m03WtMLcSDRY+EJqU/T61TFkZftQPb6edvSVLLUB/sLB+wGEdNqfi
3Nc7Wfb/hMF0+C+GcTbISOYh/DI2mLmCVwrGF0gJ2PIAzpd9Br3lxoBwp4YhC6jL
qlfNoHh2GHC6Axxu/dQoxJPTnuNH3lEVXVcVa4wdYDoD5EwZRad/y7JERb97hiNp
jQOw70qg7PHtms5/Kvj162D4NgaDyolqmDOvssokIQdkeuBBs7FvJ/0FghceeXdq
QPWpFFgQbIk9xwxX8r4Suok5BKEM/xmquqTvxWBV7H53Mxri0sJQALS2LCIBbvtE
YDX9wc6g8KSlwhRzftp016WGlqfw3n9XaqT7RsR9xncQkh6zF/urpFeb6HCdTMz0
z6i3k8GI5oqPU4Nw/x41f4AKQ42uZiHRxx0+4DgZvgI38/VghN8oqyp9TayqIu0V
fclO3Xd5O8/x/Xeg4Z1JVkMAz90uPQfbyaIBdxmCeaznRyX9XSgpAtjrwOmDO8Jv
SLO4jCl8+6kSH/MLWCBYHffiwAJ2cP6FbJ9X0Xcl/PxcDtzwBvQLZK4WrN2Z0UBv
BVKqT5fbZDR34AjyKxdyhlSuZzE517bJsoraUl8a5+UczMIf2njTaxeR0dSWhAO5
P3GNK7k7vz7J9fZo6b2AWIfPWYn0zLojUnUl/nRR8KC6PQAkSYCO3KuuAn2fs5cY
+zclKWAjIZwWwge9jzwmqj2oRNGe4q2ALhy6/DHQSDlRKEUGkz8InRGFZhEyKlAW
D+LZBAeFYZzfjJrca2/J/m2t+1fclr3x8oM13gfes+lIIzr6mhAjBDJavcpske1d
4OtAjFektV4O3wB2TIJYUB75klZxgp7o8Mk4UwHF0U9jLIFvCUi/vqd7+TI8newV
hJZFyLRipQYXyWCenFAADFI6o/l99tBnYeAu166QwUIARypYtPgb6ADrcELWxxqj
FmmewAf/XGfSy66ifS8ZGyVesE8uyuklnvTYszWcY/Yj3Z+DqjGWOWsSdPRqv5K1
Q8NFGBBltA6z5jj9MBYGe4KlDZePkLvuQbJywbmMS69KrtkjftxXUScIyYXP3bVi
mVYzHQY/HxuqZh/hngeXnz0CpdXA0BEZm/uGNtH7o1VSgSOnICAl884vVef2BtdP
qS0BDNTWQoNvceMzwlI0MkliWSshifmWhRBGqMV0GViX7+ijgbJqLp/+eVxhc6vX
ejCyvncIMsgMU0A1+rSF0D1TweBf6WJ0pKssDzSxb4DjGlYVikhTXIzCiozrO2UX
u6tGB4TpRa2igDDlP5rFyNCSD8r2WYRpEEBr/Hu3eB4mv2mK7+HRTo0LBfCOknDm
JNAyZILOtEV/3QWSDWgotWkVWJEXqOavoSarddHoAfrvDuMKVtmL+1LeX7I6NSCn
hax7Fhnbpe2td67g+wIROfY2S2NHqBSgncBFVhegK12oYnAY4c3q12OcaUSod8F8
Jh+mD2mK4q1rxeyrYLHlRRCX2Wgd5dsxSlgQvwhJ6KDFMKYq0OaHaejsJDMpHm8Q
qwUsibj2m9ECbDwVT3HEInTH4kyzPJKuT89iBvLTSw21EUH9qBToV+mOnZLN2Lzy
oqLu2+BFD6UKdWWdV6jA2LgLKsYLU9w6ec8weeKQh96cbSQKLv4/E2VwQpuf94ED
o8wgCyPRfJtkILA0ESGtKl5BFDoWMsWXCaV9IpwrfMSvWXVzNciXqC/VJSXokABS
pDeK7B74Y5TgCYjbJ2x3RljEHR8MStU5UA772VuUgJ5Wwm7Vf2NIveuIxoUqFegQ
e3HtOhRfBForXnJfwc61oseQNbezTYtn8B2Rm7QtJtQK1IToSDJsfYFR1zltkeQ3
biNc5Fs9/1Le39jK6xJm9Ls3Z35GMqedN/hx3EDM/w53aTc0nZx481vc7rJDL6KH
nPJ8utLAApT3P0QLqdxBTqTkOiZDY7P6jlXGaDmgTf7hjbuXaSt/+tt9A0RIGltN
z1I66LDDBBACBY42nJg4Qd/dGJq835FwAt4Ubk47hDpZoLFwT5UaFiPEPr4mODYZ
U1TxqSXL9s4oIdklCY2mk/Eu6utHXtKXP9THNaa97eogTagd9fR7n6f5KIMQ3vQb
Oq1N+zuOP2Bxt1PWxlnHR9YKWCdtyYwxswLW3z8cFtMGJNtM2xwrCdwQNGeYpN+g
HIGnZh/VA58Uek89CWqsJew+Afhnv9+UFyFNuC3DdMEGYPwHLJ6+r7PiL+3u2RdA
ehAWoSyR8NdB0qaO+rgPETwEv3m4XXpHhKAzDigqQJ4XxrlSi+ScaQ5GHIUTq1aA
Y7xs7qiJrWLqr5w9T90oe/c4TamLb+jC2WuW3nWd3zJ1lJkQe8aEn+MmTzq5OT30
oMKLPfCag5nUAClFozzBxmIVjET8LArQV74bXvlT1d+QvE2Jxz1+sU/KBgAeMwYl
WoJX9bXlI8ot1ca3o+72Ka5a+KqchNaUAYX4ctkGoM9ufuzILQ2NXO2wgCHU8fQf
voCVjPfZoU5w/UFoI1rWscbFDrKZNXw6dP2ck764RngXEC7DbtHXOTek0IjJoKOo
CJveg13Fq5Xs2IYh/8VNR9PSD8M4aFLQN9NupGderMZdtDszFSiu0CW2si+/iCsl
jUf4KbKgsZiNfiih6y+VQJfet5m+bL6SF+bZYkOyajFPpSVvG5gv4+ArNKM9sYfM
XmL2r4HFDhvD01IO7fjZNW80HllbscST1ZozFldFuYi3C1+M534DYbAhRhNIiC8U
kjWYeG6C9J2d3YkCb/A67INLhedfEEglYWxiOShrPEhl6luWe6eGyGevrfh5pW9d
26Ta2sOm782Hw38QEr3eBtMRdi0Jchdyck8soGUY9+5aE4TGVy1ZKI/kxbJyi+LN
NOb5lW/BR4vhM3KbUp8Xci5DE3InZhImvLlvmaIm1z4MJoLKFUiOUvmWVjAk9qfT
WxCyiGdDEoNvGfAi/Ftgh5FXbajj+yCqZx1TZdUU2A88iKqsQc43phLPSMo1P1JP
2c/GdbQmbPT3RZO5HFUOvaGvej7R3t3PafjXZQIW/0R2r5yUFKtzPtfo93MC8daB
UVT3sCAas8WgYf5y74xJgja4TyHksDLRb8mM/gQ/G9Wk7RDHQNbLSjYZE/9BFz+W
xWzUvZtBU4gjAuRzuTc2qZPW3PGR5tEQscjOUOuFkOHORn/e1pTjkBfxTqOUlePA
NYn3jfjwdwmzw6Z8GGHuJLEx5JSwIF8REDxgJjx7H/R8VMvHKKRcsmMRjKHo6oo7
66IQTDfFkL3RPA8/SjsEovKcEWaPBY2XnE4oZmuDnyituDB3oihpP4MtnJsVzMkL
2aBiuQZe36qaEhWeFHw3DKLTbhRG5lQ4zoTcB/L8K7NOGuLtc55RI72KLzZnu1ws
KRFW7F61l0EY+8gGfAsCxsKGwJsgMzJD0bJuQQVk6PxHgWsFxuURfmfgOZoVSXKZ
PbJsdNWMTSfiI5oIEMeoJ6uKmkAkTxp1vCyTFhBOfPp9vdVYwaMGWrLTcT34EkOF
4Rnt63+OuSFdGJqr2gVGQEgopYYcGaFiCiHdBcsioaqucj/605FcOLDVOcUfNwyh
rMwUhdkEVUv9IZn17x5WrS9oAQw7WixUTc5lK9kCDiTE2QMPlx0l5g9HVfaIoPM1
iYvummKpPDBzYjGyRsCxovn+vBnHR5p3ooIUuvngZ2DzrFuFawH7dqZ6T7B2sW4V
/7U/IXSslnIWa1NMR6nZr95s1C6ChjA4rrxa50afpsfuoSMueQRosjNDoExD1QjJ
zXnA/CMjPYa/St0WnPK+OWDpS4R7klXWYaALQqIORAhmuu2+VDNzAyZ0wZtOfaD1
Hb3wuZFqwo55VJEa1vf6uxD81olt0+C0aTO+ZNbmrDfo1k/5PDBODVPkmm0Fi7Ec
4U1UuLvhV+VXtUhsCHe90Dq8i2s1hWKqRhQxRyZnlN0/pfVzDsaVz6UlK1YH2jwm
CAjd5vRGu9XcJhafG7nMiZITxTQuHA6WAtaXoPdJ3cvOqbn5ggUithdkxZqH5MsB
7oVCdGnTTnFGRbWoqIxsrjqNWR+VE5KTJEcJSWTVwn9ZfwWrcLjxYcywguQQmU5O
FtXbmvmyoJxIBKcnhadQRr0ETAmGZUl6gteVtmoGTang1XiQzBornTaHXfYfBQEn
F7NDy0ZOO9k/YTjeuDw7NHq6ycvKcPiuWC0dxRIDxELaroKaTdP2B889DWtQtWkW
J2t3WJhMYTuAiI39e3dFlnNfIkrBZmBHIRn0otveaIF5arCzthuH+imLmH8cePoa
YCR0ckeG2Jfddu9jphBh9/+k55eO/v9dndBM7r8wt8yVJDD/G3YX57oHrZSBd3gm
Tz5bWiUuIPTX44qYmamXomBV0R6x95y3Y2IItCsk+AqygrqugcOzSmlJMkebIldB
Ux+cgxEaSaWPKB3P+eLTZ80RpSzVIUf2GFeGsAfezkxScH+qpTeBofqccVyW71wc
Abu5NEbA8nfwPlcvQMpyNaBLUknkS1INlZg62h2ZIt7ncASnMpDXwvr2p2Af5TJP
PhaLrhJhMyVPYg3sUd0O+EnbOGa9QlYY+rDo3IGeHwGihJJrXw4wejMLAC+E6vj8
+U6vXkjcs7Lot+7FZp3YfuNuvB0u1C3Lq8/dpIDjRcwlSPqZFYeDMxMaq5uYvWjX
xWp3gNLVHT0p175po+yFgyIlI9I5vvadrdxqFGdcPe9d6Kjyxh/GkGFbaV6clKF4
pghXk9xrueo5vbAsbrXimo+m4QgRhE82ueJRxvzfMdbIJV6UQCi5Ku8NVRe4jsSt
JPalLb4x8iFht/DSpUTDElKV1BPKsxXiJuslEPVkRRpMmzxhWint1Dh6bNBqIevf
2fBoVBH9gafCkUZY/Vry3aX+qIuWyCuwgpxK7mnRjD982UxeK+4H0nVQVOdDATbA
oyzcqf7EfOcLntWffI2XEXxKhs4FR7xYnhtedPvY9n2yxWMSTJvv6zzBftp8jpVL
9NQeE33c3Wa5LVZp6nK6USEPDcXL73+WtjVIq7lMUz7FcEyxX3qmej3+JbcuJz2T
x10eqZUuDg3TeiJfE94aLeHVozY6fyD6Cl/A6q5h6+EVpZ26SZXEU/3qd1JJqsYt
sKhF5lFfI3nffqD4wEvfV3xCbm1EskLd8Bo7XCap/NGrdUnXBnAHFRXU1MIXGieV
OCsXap9BkwUDQmsn2evUhLOLkEGD8cPo/HKGwSXTcGrhu9n6KYjMgBhZa+QFQckS
Qwrseb8mWvrhtJnwYgE41i0M7p1OckCHTj2NhGhJQBI9coopOWDjXjlbO1N0qweK
BYFwCS7bnEZTkt3ItmgZ3cLhHd5iB8XdCIGzxtHI7lAz6Ibk7D+IK9QtA5tnSrHE
MsC7Fqd1g84EPwvshQehD7u9wmRAFIeQ0EuXvs7eh8rRVROn//mzn3w2/CCeopNH
7bMVMHbGN4SnPeTouVc9/3tH0wQ3cIOOUurE3LG/c7rnog4IpSTh1KmJCcnaCsWM
881N2PmxoYwAYkkqCJI0tlFvkNu7AElw1rumalvoUTx7GQmoZPHlwqxBT3EKAOhX
4BYCjTVcR458NIr7kTv4nMvgx6AR0hLzeabfTY4oSjf2zSkvuKXfzDQRrP6NZaVU
rx+rTDArvTSb48jjlSdhZZ+b8cOhsefXJtRaAZlSRtag5wQEzBFAJWqGO3bmsAWD
c9kbAWLS3HjJqQh+ERbHBIa/A9rG27BDeTvZkg5pfNJHhao2yLtCS4WRBfEkxE8W
EUbq4l2uQbj0T1TliJSrTB+RFqHtYslJu6O9s/R4fsb3IDAk31bjEaHKGTTCBf/A
DJG8ymecOqOnRGhAWq8V7WLMZfcIQNM14iVrNq0GBVqVD0nySzxQj+jpg+sSKfMl
y/031eCQGZ/8VHQnNT9P1WDcmqfBkWVu06Nqju4pE9zB4aRbXa6QzQnPNFnD+sr9
eIYFCnrMAnF3eZ6/Z2zIHVKt48SGLpt9gwlLZk4Ib+dvXPZV3Qx4mQeH5VYwLKdj
8wGnjhtxpTzlALHz2IvXuqFih7z0Aw6kSbsdcFHzR4f3xg0cLlX26qQ492EzWPDs
hr7lYKgB1WhqCz45fwdrWdrUaVkvPj8SupKlwDWvbF4btpj83WMlUC45Imcg776j
Xo6ShRS+OZPygslwq28EgQvHs4+sviA7owrVt5AWK/TQlkcCrcqeokaKOZODS7CY
+3F+9VdJNEIW3L6eE8LjhWXG04nO792IgCR4uJZ+jg5LJr3l3divSjFNTVgx6lpx
bwfyZOrXX5b4oyUQ9ezSD05eRniSkkHV7PO6hVG3ETQ7vdapJViccvrGAOzKbSaT
xFpK/Rl8h3BJ2YGuF2PvVE+1DlpXa599xlrBQPPYdWRY9RNh3bv/G8DjWWP6QGJg
pIQS/qhQmNc3tfisnhvDrpejqDd1ozKKWY7Q0vRGWwC1UrWICmSbMJ1N2SJ3CmNX
jfa8OZJedmYgV+fqvN5n5PYK8el6Aq0UgPcN7Z6rkRY2rRMLCOPXqCaZfop+cKAX
bdWWGSKUjlezNAAPxHlvexzyIPohzC8AL+BcABQizum6kOCaS8i6faHwd9j+M0Sk
ASIGR4r5D3e+hafotIqKq3iyRZQdjdPPL8ouN/CCb7QNh21mNXP/iuFwnlGrH1GL
nFTGVQzfPWf+JO85UyGh2G4ufmvt65UjlotHrueUwTkEHt9cmm4ztyuAC6XtLSPg
vCFNSqU/XZ/bUsxJuXhTdyS36k+xGL/9EREaOZGu6kExPzepi5+Z6OZjYgWVAxOp
TA9CEFTAvWwiCaFLHWAsOiX5PxO7UDB0rqxT/CxRG6bBgz4aOlsyXK6Iuk3YktCm
xq1zIexkWucg3HXk6yFROlhTTJrGYA3XN/zRLOSeOJjPc7vtM7ieljON8wN0o/Yh
GikZckvhDfKAy8wpn2ueqgvFWQBlnvu9cvxj8w+F+l6nTJxMoMwBjw+0UfZZP131
3p6TgMGGr+aBhV+qHiHe/GbFbxL6NKaB74OUy8g2oN2ri5CDV9xWbicLbG2QjiN8
SrBsAGH5YskfG/lChWlVZWLIoCYL1KLjICEXumIlYAIVncyl6Y7HrtS6h8I+lJnV
8brz0Sl/edkS3ECHXVvWvO99eLIcPtHfTEdcNERQca9UmqOZioxeEzaCNCyrh0bd
JvWHJAl5l0nZe8calj13KghB4LzihomzYwjbkPfkuJbEp+ZVU5N7L+Uc6Ai6mRFv
/ZwQLP1NrPkOLh2HrCLshozpBLNCCkM5iLRS5/czfWsLy4uvTUcBPyDywHkyiXSQ
gsGgT+aesqinoVBQ1vx9t5HKOykK4Pw4argOsGuH6HSo6XklLY3muC3eZr25Bkhm
+q7+QRANXImwcIkhC/7RBMeH+LbkLwP9/044Bb2vBdHz+BTLek6jrrakQGjFYLpI
viFHZLzGTDXKsb7LN87lkHAe6X10svz5rsBLZmBLwFVCxyTlFrpGXVHVASXg/iQE
zHQSOpNqR77r4W6efcLBxNqBIY7az9eCtly6FaqLTvVqPA1RyAKQIjbImeWN2Wm9
/+ISgFNg528wv9sLRqYlAwWnmAj7ZPozQp5vhfUm6WdO5PI406V366WvuPDDO0DF
+dbGpOodE3ucAc68ZPL6cHzLCThQoJQxcGiyQCCD8bTtmw5o1wQH4izOWyUp7+Eo
8lr3nmwqtKwLg4wXtd7GkADDEcVSZMLv7GH2nNfpUmB+dCwlxAEg4vGePIXHraQT
Wca/JOr30+eCrUWO3NlqjiXbXTVA88zBpug3mgO23Bw7AGfSasod+eDAkVuBgiIR
dIPCi0dq+k/FoS4TPsU/QjE/cvpurnI35RFKjEmLFhcuaW2EFeYXq8BbSl0xAMTp
K8teHQPP3YZGNKG6ntEZRyeXb8cKRQJKn4gNyJO5jsbXef76YwqYTpkRw4bbtO1J
jPXqfgD42HRtooaGlEBPxnnr1ij8MqAEwJLODjTqB+htoIvo8z6b/+mGd4rjcztD
L/qCWiR6ago7da1xuQ5NtwakgosQl5YneFbYemoy2Im1cGVNNF5gfuxyoLCs4hVk
2Rg9MlkAnl3lIj3FpREYlkTruhMncRsJOnDQpaTgMKuRDQGDhWNg1zkF6MBDnhdd
iVAFc5rXNz2EV1adpN2Ao60NkLA4Mw62NY7GV4++nP5mWa51Um0VAg4Dslx9swta
E+SuPDZIFkz9PINyyFO8iYaMbzEN2wSNsmqNl8BM2GTnyvkIhAourC14nTZYk2x3
6NXAfbB12MmcuZL6Fw554PvqDuNznW6CFaWAikHufWiIXaKfwA77B2y8BBzPvZwF
k/zXNYmSm9bhk7GQ9vlL7Rc9rB/dhHk3+XvBh2hjB9KkrUNWd8rxo36FPZ+XaRUJ
IlgNLF1AfJ/K5F0D/UxJ+4D4fp2XKGVlE0F4ZWSopg9XxMXAGiy+ylahRmitN1os
MT+coctwaW5d0UAGWf9ca5iwMkqsAhjG7Hm32rQ3lTCoKaCFTvP1vNJxdvQmnMhO
J0D7MLTm9WPwTDfY/fieLr8emF76xyEFae+oo3UWjvG3/XBztz8NI5IwQXdtc+86
Xsf5gB1agx0nIUTdquYBWpjx1lJuEsp097Uz3lV1azzJHjtnvTRpynG3e4bOklCV
OW+nfB8r8NOcSFNRKNwK/rpzQdP+urYueeZw8f/yMqjNLScQSVzSaTkGEOfEVbEZ
mxVDlNG8QAugMawgNafvYkR1Njo/8Crl4DKUFiEB6Log+FugX1RzonwSOUtuUWLj
JiHDgAlz2zQBNiy1ZGKUcMJYPqQlwXlQWkRbbCM/ir21TMogpGomCrgkV2JyzDvJ
DdC17QvNl9kZ46NZRF0Mkq4Q1IzZR2qGq7dODs/ziGMk/qRmjm2s2wPOQofg2HSJ
WWRUfYJ2DsvlN6YFdgksa4BlRaoKM8vOi6f6JOcsGGZP4dOCZCFK61Dj+wd57F/z
xVEbWosIZ7fys/eo18rg2dDg0GzNASWo2bt/P7f8bbQQ86DcTLehNmShUxNMaNTP
BWJXJnzp1PMoaiqZoe7yMX97P8wBvM9Jzxby1FKzi8B/eoSod8H3SZfbAbtp1wra
r94DwzzocbGJofpdshXRGCEj2Bzv3gFLWV3kZ99QSUWo4ztGTLddFN7xejl749tY
1u5L9966DvRZ/7swAUxUkerTT5rkeU5Wpqvs5LYZfuWAO62kP4zxds9HFZLxySiW
WWadK2i7FzskIpO41kY8BnI5ZOh0IdsjNz641gWr1bW3YBRk+YDswLKpMGLorPEt
GCL9iEeoAD6euC62VGY340WklGzsF01k07SteYDsIwzNRYT3j+p/D/DUV/5qMYd3
MgCeMsctxtLGMEwieAso8zoWldMCdjEfInN37lszAuj0x/ZxBBwSMyQbQcgnsdxT
m77lmx8TBo2Q2esQ+bIldj2y9lfLgz9RKmWUi+zOZMva264NcLWfYzArSKQkLDD1
Ynz6M4YMEnUD98bwHFtKMRV712Xa/wYb4ZsxL/i0W8J0iFEptwWMDPPgLMU3KZlX
C8hbjTT4F2diGlrcKRBAugaOtkzUyZtdcjfwCYZ9NcemNc5QFJdYORYL53cscBSZ
C5SPAdq4ZrKP6vRlu9xCVzvJnyazQezWYAqit3utxRWIHakpfDUBZQWAsNR7H50X
iNbtgs3BAEqJpng+0nk0YszOnzpIg1NQxj68ChIYVuVw3FolM93Tp2UJr9ffmWII
NR74w+wChs5r7/WdVGrKOWIWbOL8Y42dAYa/5+HCwX9jYSAiItY0fbzuCLj1azmW
rvuJUGOCECFXx+9xJfno+/fNksWaG27OxjkCLREU4OZX7lKzGPWx4El41PP6L+eb
Veh3XEXZufEOlyHGhYsWuac/l1lv9H6eOFh8MkTloEDqF3Dn9YOCABb8HJ7k6Ksj
5CBy5j0W7ANUuUDnZ8B1aQ/hBYnAjd8tMX6NO3MDB8WcTSaBOvB4f8Ma3iZifgU0
7IL0UidzwVEkmxwX3dEmNl8CcohjOriMR3TFr6NJ/xYNGjPXmN5BNc19vJ4Z+82h
r34HVmhb1ayXqQpWx6JfpSYla0A+DAdhstsFl9rBt1khn09krnQMZFC40f4Kj/eC
TDfM0EuCqddQ1/cbZ0j6jI2a0wnF2j5hdkrlfrvpTG/kLjf/0HkyMPan5pkis14t
f/mqmHve61pjYMaF4utMl3zQsw7S0Q7HMvfwppn3Ds5Wk7Pvb6mE2O9K7EN+kbSp
rafhY/E/1y/5ZZrGTV3+fDuX/TfSWhnIdNs50KBw0aG5b2SLe/jXE8Vjx4s8Q3gr
l55Ms1Ygd5mgmPpaz0sLTaiGXH4qaBDsYZ7kZTLpjdWxBOf6ZqMzt/gszl+yar76
lO6SY4W4fOZ8sTc6dFQjkx9bJNN2HDCpOQbnaEVVEWOdnn1WvzQMRHk0ATCVECuu
ljb9O8k9rDf982rDmHmkJyUXzf7+laW/Gi2Xfdjtx8ujEbEjXcbiZ0pVdLn6dq+K
hotDSug/IrjvhTSVVd06ukCaU065vBlq0+BCUXrYe5onPP3BHtifXjaJ0KFnQ8gV
hFI8PkUkW8qfJXvsQ5E46lNDl8SK2ZX+uSpTAyegOjdEVoUx28zq8dCufvbu5ewG
dIe4zeifIoUnjbxNzp9XMP/DZ0XkT7JUzkqHTBEaw5FkfUkiC/oVkzllRWm59hs3
2MdXoykeAZHU0yi01mJNDQb34Se7g/kZ5gPcUABai2DLmN058YsFnEJu+My1bMzU
kv3W9lmHFuaIsUem0VkKLdiRe3872gn56lhmMzM/IKSssJhPdrlU66Te3l78MOlz
ZR/pn5aje5G+YMsg+WDpx5K3XHYjRAtp4b50djbMEpqrJBfOoJA+WhI1ee5d6txr
0+puyEJpbMfeliPWzmd2nRsz0eAOgcJ91LBNDVVW2EtjTXsRiYeC7RbCybXL5UjY
hd/hVSZN4T3negEzTaw7+IaCGiIQB89ZdLBG1odgzYRWjlba7B+IoVnBK7YoDu7y
0BRComNgcXKP5KXhZdKhgOYvqYp9Qv2NORXWgQ8SczWoq/tnIyoVosEP9eeUx9ze
7PcjxyKc2mRmB+vayIQcLOblhpFU4J1B+lGwLEUSmcaXIZgTGkA9xHdkVh0bPAM/
sLrklQOOYU2ld+e0ivlqEccAuywwyb/vvdvSxM0ry5OBMK+KquuHAKZw69QGCNqk
9b4nfvwIZYONGzNz4fj3hd75DH4cMqLOAxu03Ko8Z4xWxYjbBuKrCHm+ZLY40CCW
EpPnjWWPtv88P4GfHPzzhC4vSoO1jwg+V0/WkJq8q5fc+NXkc/FSMfYs3kTSnPvb
wF7ivd32T/Q+su96z7ldFCsoRCxAWY3FKPiUm2BNtCs83Ql2oow4aa3twL/m7c4j
Od/MjdI1n8/Ew4kdVPoYjTKFkQYeW9QwAatoGwBRi9m+6Ar45xBplcF6RslkQmxv
3Kp8e+vq0KWkfn5B7Gvj3r3r3AHq7YpOJ0gAw091njKHOF0NHgLYwmN5c3FisYfb
PW/AmkpDN7iwRynW69vFBuThFg1DLeCx8f53eQc5m1UMbLZue8rZDAkRWFR4DckU
OcwmdbSkf0eRwS3dcASfax5/ZYbQfKaYCsrEXQVdOsKyNkt1lTiQS+sF0HMYMVG1
/MyRWouh2I8PmDrMhl9nrg0lzHjkXJs7mWeQa0D1eZzP3nESmnyEr6Vnfk5oJjWj
qvzxUoJk8sTYAmxz06BtAKUWd9zCeU+RYRnadij3RHao/42K6Eba74Hd1TBj1z8B
Hyk29Kjkwim86lBNQNFLs0MSWsCTpaoQi5QcxbitI1stm91PKw96qyAUryPT1DDI
6hJPD/O418cW18JoGP7WrjaaBUUl715Q+pGAgD4ORmiqtJkzMTz5jdVpWaQQYNMN
ka/AMBC6/VOx87nuxNbK6FgwretWoe5VyoZkSLke1ojZeg5wpgXKAtJJgBa8GQZ2
fiFCCu+lhKuHQfSRtE6+dyU2oweG3q4aGLIQTuW8KQr7G4fR6QGn4acpu51He/5D
idQzFLq6OnXckyDJVEkx57q28esrEeJELTnAPDanrs8qoE8SlKOWVi2UcBMI1W1d
AyhZDWYOLLovCaZHKJ60Q7qXTUxDKn25bqMjqhe6h57rcA2eWfhWqRU0WjDZ0Kgu
gOo+V/HF5QZOLgZDMKOgo9/gq0m5ilQ/yY8yd3/lHFJlFXyDsYI+feY/fSE70lHw
STz7uxunxuiY/nWw01kBiB/omYnk0lHbVTQ+i4ijTDnUH48iDZKc6g4sGinKI3pp
gIBO5GpwA7tsbCMPHJYGVCyPw8kY0puEKwmfmZX2CINaCU8I2fsgqqAnkrLGlHqh
gWszXK8/ixp9o0Y36mkNucjIQRBooAyc4ReYSsWKZU/uuTkPW5R9SY/ecikjCBfZ
2gIXuV9fZZvSUr8LXdhbq61jLwTYL0UCIhVwms5b5Qmu30j8iPCKZklanqgNr4pP
gEcmLAszTf0sa9bB8B0nXIwkWeZLAYRfP+AN1IYmDWgxivBHh9L8aTpuHp0WNvd2
UgTFuOoB6f7nVfjkXywsuccXimaj2Hr0WtETvYdNyUhF/AH7/MBGpIu8ex60Ub5U
Noz4RlboVmK23Xjf1TpzsW2hP6xuyymf8Wy21uFuKLkUqUXICV28ql58rvT2hTti
0a+o+b3FvzrLqcuarKVt6Zc7hXsQisgQw5GFCJ0D2yDWaJur7DovjGr52nJ9aRq1
icbSWOul8yKxMOwGaG98YYI7NZ+syqSTZbzRZNjjIa02GZcvAy0zDh2cVUGoajK+
rZYoJiK4xuyx+k1jPtFuEimnzEhU13+EPydzim18AeqObmvCg2pImyfBOgtyPtAf
wvPhEA5HnRu3xx7AEZdaDPEWOzFLNPJ8wMdStXlQZGy0wQATCFr8jFA/CyDF3Y5U
l4AgG0tk3RqtW/s9mivzRSpAIvKWBj2XJYDBMdBHZBd1/vHRqVjNZ9d51SRy5YB9
cP9P1mSFqnNF87lK1jbrW1yw4FF4CKNwnzb65WNq9PrxpJS+HeSNw7sVgcEHayfF
3p41AjO5uTqtDs9uF6n7bMxdnRlZAOrPM2h/12QVYKREd57eZTVQ0RC6LcJvr0fv
hFLRvYps3EfC1pdhPlAgOYibtXaGnX6bSEH74M/eAQLLhIYkc+jiK0RtxO+77ZaM
zVXaJPnVALNjtb9qi/86TMMWW9jROdHXcj2CK6KuzS5nds/ODAbXV0J4amJQRsQt
RGVs3rHV2fVLLpzd2QAE9ZJjmJk15x2c4sCk4RdTY1mepxbGFjnSi3/7uYTlF2t5
KkmygGPqSkhmSxLUiD/rIH8qVtzec44M2Wks4ouA9zeSfDQ1ouEAXcIxDd5986qY
HPjqb7K/NdDhbnv5xTPXN1Dh24AKsvfk1Z8+6CMzV0uGQ2zd16s5I/tdlfCtsVcW
F4nvoSvO0qSzu0B0fttgrr5MUwPnsZuToRmqygxaLmekYLC1gCSg1qRQ3OVGXPm7
TzGNwpkQrXN8cjScQxrrQ4h2NhHSlwnkV11uwpxLOFkfFIwp0RYNgBt0eS5qBO2a
sKSnIHdPmF+UhmFWjIm6l54VepBIKFcoMxQytCh5wVQJceBM4/fke+Vv4ui5CL5n
0APwVO527MPqTM1tWmni/dExB9Ov3LIVdEdVcw7+YlKMy3Ap65GCSntqeDyqDyqM
y8v3W/KCHtqUtKELIS6aI+lSEKWLazrs86GQ+Vc4tVll/ubH5SLCTTQO0i9f2luq
LDAaGm1XyNwayicaHi1sHM9WIXuyv1q1lbERyGYyvvkuhr122k9haeITa6N4qxSV
bQcAvrtMNevLeaGDI4iO+053iH92S2vnvq3Fd0CSBdfksviXBY8FHC5z40M9I66Q
h8anwbe2zdvoL24U+/TkB8Ud6Nn+kAGJhMxspFacpl5rcGkCI4t13zibhWiVZbbk
dTN46eCqfSlWgAuk4iJJlwLssbEeg2214K7lfDT6jxXyGDRhVyhdGS3+xH8B61YT
1gEz/h6GgQ7hURVkrZ582lp1qZQWtLwoCxVYLqP8Y/VjFgWOeWtB4tzRsI1R2eg4
PO4WFAprRAEYg9jplnUsGL7nj4KANsgbt4+VhO+uw+RXMJyf7X8p1FWLU8wB9jMo
FCFS+RHmg+UbzskT6d3jQqokJvdNLV/rAtcoom+YpCZJScFViTfyfKT/NQEpy17R
WWxwJxXuNMLakoInogefgOW4HeZO4Jxw0gZSRzeciRlOZfhiP0tQVQ95a1nO+IJh
Up76gCs7VycMerodW8nAcYwQImwV4DRZQhaYbr3H5y/64YsQLGmgQwXCm6CDOeP5
cW22w+NOdxTZSyZJsFPy4bVzkiTywe5bId9FYA/QIXG9bfZ8oVaVmkeSejtbigM2
M2zsPiSsq/06njneQzGYMVs2OwYl+kFf+RtMyshRBIYEEgqWAxBAL/SYLAhuUW79
ebpkh8KMmExqMWv5lQ7J2ZD3wCjv7ClttTve+/p4GojNAVss/Gc5q7dy6/L6AsmZ
Ev0VXYljSNXYulBXLf1BXTGCEwXb+/ijkKhLIov6ADTdtUtQvSF2Gr3f4tWm5TK3
IItROq47oqKyk2f5zHAkHUGsFqsNGdnqftb7l36Y39pqBBlzM4Li/GWZhaq4qpX4
rfvrNZLRi7gkwWfzYkTQ0cbOg1cCddd7cw0djMvgUI0kNLTMfQ3bbrghoORevHOB
DSdFwtSZdzfw5vnvrzEXAdoQ0rw/9k1vna6+6R1Gl699hZvnjU3gTnbzkbuOwDqK
d5riJrwWLyd1t0yvZzgZNJBA85Q/BmNE0yUn82Z+9zUqFkj8CqkF907MVQJpTZbr
EwdgKL+p/P3e2gZY42zooRhuv6pkAH4b+LtA2Q0wL8cOqTVjNdoGwZ8F+K8JBYxm
mCR1MT7YCk/m68OjY6NEyqOzRDrg01ygf3DE6t3gv+YoKysGfj6JW8VmmFC4fMKO
S0R/aZ2rck46qFLo1niPSzbuMckF13ynQQD+5GQ/5McMmsD0xhgREnGer38x1kMH
utfqyiL+HWHLlnalwuQ0qqqmBKTsE+IwnUkHmy1pvWbIA1XeDLGUJOusXiY6oBia
ginWME0VUNcXhT2qVIEtpnhhY6x4MYngKmj7eRHKbz7j1QCddp5gJZox3OnqcbrQ
Hq6QndBf0Ag3yYd6E/1MEc1k05AH97bNUe3Wvp8laCq8eccffuVl9kNJBevdfC3c
zXrA4v1Mxf691k69YFr3ky/ADDnTUd532iyuOLgpOng1i5nfASCljam+/Zk1JeCH
b92ENSxPjmZtZOxmBiZHl7qgy0vFwu7mdME4FC+eAL/Lpeng4/isR2XNWZ7K0sbI
sQ0MNlpKJTmD+AhdIv+tGSY7kWogrXPs3WzJcPGrehPTHpHh9gBsqHFk2ShvMyhM
FXOFZSSDKngG61+VKV7DqpuYWJT68P3Zhj6Vh67jaVstcBc+sP03UqKBCMS9EbpD
TCFULASYQYL0T6k9CHBNhSZz57XWSJFdC3gejYiXNv9yOAxSRb0XPjdsebWsVWoU
NkkWFiWkyVDl+E0Xm8tFgkekE0w03zhcitb2/g99wOAThgVfXeMkMGJD2uU56Pep
nuF3tePsjzOIYypObmOlPVhLyx2MIDwzCT6NFHonsxbrNzFrTGeMuydB4YEeIhOl
QIe3zwQfytbetK/gvbinXcS4695jxeIYxL9vfiLqQtJtK+T1XzaC1E2HuH2nyC5S
PzEntg2bfM5dKSb05wdHp/xfnOTOpD/GTqa3s/GOyRFuUCj3ygZ0lG7TaBxZTdL/
O+vCG7t46Ttk9O/KkyY9yZY0n8L7rvrnpwxGxhAcf/H7D6o5lbUKjXR/QV2uxp+w
LwOtvBXpn1juZLkJcJHoCzDoFZcjLLQpaOQ0EB1LQWajypvTFuJeajgl4tEVPjSF
QFp+pdqZIMWj2efWEudZlvbYlUmvtmfiKaUmZxXKui7rXw1Zn/hF9XA4z0ck7HmN
joWhEoDXpPJaGaUEAND9X8HLIA8mkjEAiZhW5sShjUdoRzDxKvDBEYjYrGzoD8OO
dn7JmhHepcImKsAGK/91rQhR04ZMBPeDCWKhNa6wC2AIXi7B2C1XuASrz0QR14R+
feUVCsA+efsfQZNVcrLKxwfZUGvbF0sq+zQtbueJg0UD6c65Aeaan4qVmFJRK2I/
ibgAPo3ZPGDqvrGQk4KQcTgikorMqwdq1xQE3y34ldZcUDR4lWzHp/GeXsUu6CM1
c2cNe18gAyCu4uBIzayYIrDUjMqkYQG30ApjQzi+nNS0P1J1NHgU9yW7mqB4zmaO
xfHtKNMVb4bW8Cgs7ZUf8XPR1p98BmYHOX8RtEwcJPUAvudDsE96zsa5wFJgA+US
FU/0yt2P9/Gt76KBISc2uggs7enKEj4qEaqdAGAX9OVt/c/47ciIzmZzURVO7VJj
fyvUoilzYyvz22plZJpkGfuuaOGHsum6SsDEG9EFiV7DzoDoYmXlznRh0XU+mtUW
ullADjhKrWoLFayRDihiLDe/UfJ3FfyT4kaLOP2BYz9PV7Au1YZCTMbFzRhtNgNN
zikttx691+qdZ5fTPqyeqihNwMuPh5Z4Cl46QMClM1RRg7BmqFNb9uvVHw0vbsV+
0dsN1fk/pQMFbam1AjaJDZGf7EJMad9JbPSVY4FmVe+KS2t6o7QBA1sL+4kTgLkl
nTDEzWfSD9V7RLXtsAULyVC2npV1a1m8yY16Gy5j4oKpAU360WFghFP4aJrRC8FB
v3T7SdLu8FcoEV9DZ/2e3xF+LTFXAwmVQStsEGP2pcm6x0IDAPcnebuqm1pEMPPX
czkyqc6G/Mypx/7nODd1rqPeGei2I1cbf/yq7M4mZi62WtKI2di+UQujGQaxk2S4
R39flLnem1JATQ0N35US0xSUFnWBz81HBhpjY0xwq2e89rE8XPdTn9+BG7gpZ6DW
4s2LZnDzo51aJz8x02LVFoC5IRzW5XydebCxk/isB17vwcf/h+tVFRdY/pK3ieAI
8YD41VGcf9D002ZpCQWoyrjJfaMhuv/89EUNo8CJDpnN6gkoYcvFuQlg0Ds12Wyn
G6jFnQy5TEPrY3svGTfQk0+wO9vIRMMsHu/nser7i7NqMaF08+xIxlUz7JOn+auX
oem8alv/lk20h8O220psQRRnOL1YNmS5b0G92m2gQVregD2UBGJ7OF7F7G9EEVBW
8SX1DOF3fDxjrYVB5ieNHFcv3YTpIhnE5dHyruuXZrXddIl2eKz1vJsaXnme/oU7
Pf8alYfthXQS9yCbgDelfFfzMNZySIVbpTICRsh61NyN4AmEG/VAZX2dc8aUWyTv
fbbhlfl9oubDo/zsVrf3aihutwuF+lhMSi8msLYK8EAiu1tHrk0uqsIhtYXYeMAL
YMON1cQUS4OPjYA+DsdSTGj4GcxiO1TRxloYppGzZ+PJn+m04umFsJO6EHoFHS8V
9Z55Cbgp0NcDeEDLlpbuPuv3JUZdUkj52eTgJF8R7CCyFKD61xw6zTPsgSbjEnKA
Tf4f8jz/LZFF1gh1ZnHOXKdbG4ABHy187Xt+w0oKRU38nEzH2LBZim1EKMD1YOUM
O9yEh9d8WHmPf8WRJO9eEsTG/Kab2Bgj/MM7PQPpwkyQPZ3jNVJlSsw/bRFo1QV1
vmkELDcfMmT6AWFksPHoGJ5Lxrq1J+l6vrlA11w6nTbInqdZ32LonOodKZJqPv3H
mDqPFGZimqt8CcoaIiG6bmLbEv0GGKSUg5guud+hdrLSct1/b4pujSh+/N65dxw+
/80sPXiREYYGOPCvZNxzQh2hiNAodICXm+EcgUWpVpEXx+xmM7g0Cm8ZgRoevqyI
NcF4m8JsMM1dWK1Qq096kwL/aekFS40Y3dSH3l6uykSfdVx3Gkq1etyV+5MTIkB8
7jDaq1G+P/FkENU7i0aPpkyvYpCHmiAOwyz26F5FK/ms/6RBtg21HLApuGHU7Q3q
s63KofzpLPd23nqjtkiPvEf3WRQp/87WO9EFnVMDI83Pt5h9eDrMz5mF2IvPqb8z
jr7C8I7To7z6Z4NCdp0AC/sN/FW/i2QBAbQBZ9xnpYHc9f6qU95bXmSOt8H+JMDo
QtRaggqGCT9L8N+itZSBEGI5ft/ch6NVPt6+vYbRdfk1OnikF6JvzWeNlfqNZCH7
CFEXKUymMHUh/zlnLxPeZAjgvMP3vzFOuM57qnuXGXWdR+/rhQPwKerNI/PtAp61
Vz9Fn3AR8mWhEM/wgirY1KS8kqs35L+lfQxHGelAdHjYR2pzXnLqjYOVMe1/P0SU
u1nN8aiqKtBe7kgUaQbryjiZX9y6Iq/kVphJGbwoUst4zxrYULyL1GRtt/psVjpH
AIb00RMYMxL8hHTLBg+RMJJKFfPDN/fqGS66PgTRBQUklXRG1xcFyjyXVTLARYpu
NAPvfVAOAJ82ef8f+43u0ZJJ2Fu96zmgMm8WPt0Dt1hkcBIORlHCfkud0q52KftU
JbarThBCoTYfxsvLUm4/pqIYV3fjL32tuAAXvjDWY3BnPM5TPD0uxE09OKbX5V8I
X+ce0Ed1KXyCVzaRbnXbMTbqemq/g2w2aXTPn/FjJaCFLktX4aCQq1q/06X3gguJ
mBhpbToxcoV7p24PGdORNltABolzDkuabO6bY7DoQiGSJbEgmg3TbgcTW+fA4ZS1
PGzqgBI6xxfOF1t3cjJ1Esqmwl6DFG7AO1wNDQsLgpQTX6fHqSA6LByx7DsJQrpp
v4tqYduceefnUrehp/cAHep6rdzJSYKoTUdk1Hlu23tLT55RI+cseQTnMKGoILGY
7kSNseFB0IT3k1gDZPKxZNjF4ZyyHRoD3qsqBsm46rbkL+DooXpTU9m4K0Tx8SLe
CLcNLPEtXtc0AxVVp7kT/3BGPG+b/K5z6MXA0enHqZJ8UQWIPZMk3BOHrvA+G0uZ
T0fVRdHlOw+2lbWeCoF3MHw3K4so/S/KVRM/tQV0/zWVrW5yRz5p0uFMC1yWKmZy
SgyEi6sEMvkED5vikk3WVupNayZPZmaEU/N2vZpxIemh+xu4ilFL6jucges/UlEn
EGhmXYigC97XPU0XnCq5QNu9xaWXOodgNqX80DPheNCQy1zFichBoS3LfEeGojIq
n2iIsTz57mSZGa71bfsk5GmCBMzFDY3ipLtvdU9pn9YKr/FCN8XbH5tuX9bpaKbo
iXLT6n2V70Sx3NqmhmC2oIh83cvmUYIFNRpJDBStF1gP0k1bneq7ar3JYKtIgHzu
s8YRfDvAUxTVTIMiOaA6eOGRaUTTt2/g9It9GIngL68zuWZPT/kVo0Ay2AtNbleO
zJrTa6oS+ebbdc1ooqEET2FUQhmkYSkOFAzR74ynjm4d46l+huu9kmu3M73rO2aw
9FCqZRCoSWAOsu9xwgPUqFYFhANnVLu6AnHPdftbfLJ7m9S3msn5MxwROmuhRE/W
wql15KN4RG38WnXH+WnmUSRHxOeIxkEtkhrSTG6M5zXo0OHAO/oCjn4tQiJneTV7
8cI/8Rrb7hiWaWxQkxOdiAYnXCXX9OtU4vD756iHwv0VBwRtprED5npXMIYdThZo
r2r/KkBImaudq7Tx3nN2INASUOIIuoOAcGd6ZRGgj49/I9Z2GMdFZFARyre2I4zl
JE9MFLbypW1yYRhud4tvUhwZ1zFrH5d0VybnBxx5G1xpTEKw9rGdQtaxETRZnFwp
j2NBwBT1Ga682qeWCTOOvL/OPAUO++JwEnX4ASLvDnFX/BPD8RJPfVvj/UtbKd/P
pBmPcVwUW8ti8r7P2i/EvR6NShgUzLBncT3j/dgIBtlvTPK5313Zpr0xUXmfF+IM
leBZiISpwYwD4JX4IyN7v/nbYChM4iFqMj/dSE+KXD9pVDbCOFYDyg5ERxHeoomU
y9T5lYdVyFwGF80K3teD0oTqys4j/1/dxfKn2f/ltPQfaggWJ+RvMgnvGVYrTQ5E
cDO0EnG9Sf9t/YAehaqtP7cvohyaniqdrBqRayBFTrL9GhTAMlOdMT1gIhehpMHx
JYDSe0WiVRUdlN1ROU0WNvFOSyzMP2lLFx+G7dRNXiK7Vu6nJNk3YMjW/C8RghhE
ZB9ivC1SkPdektNee3eqNMIiwXgJMRVweyro18pmPdjZkCduzeoHgfHyNIBsZWR0
4nUzGQoJG8tSRpOmKGnQwt/g8seN80/EHyU6z5V87de5U78ew1TVPAvVj3A49Rq6
iJe1P0xp+J7IQ2hHTopLTyRELvQECx/9LsUqXjM5LmZVbMCxjS9jnb9AMRGz5DlU
ajU1OWDcSi5yBIVS5o15ZHetC4jCkb4iIy7708Df0EQnQ6q8LYxpLwssG1YJjLc/
lVgVDtPH8PFQRZg6hDKTaC49MryFPFrczbK4o9rTQpvNBPEeujT/a6JxZhYi5haA
U3yZHJgu+PS1sIIplPI1DcKhdZiF+qxze0EY7bqRLhpsUfRaxyPKiHZrynd8sqgV
6AGX9ttH+eN5M8yJ53InU0QhgRLD5wwNVVVPxAnP4BMm5QaWApWdo9JjdYtQ2U5L
vklQAjyu58v8i/nhU73Wp8KiYVi0ITPjsPgLrygx/5Wzh8gAn7VYJjS/yV15pOIP
Yst2KQVVStpujhrom288zDtt3WQBAptrg09YNwlDRGAtSvn0n3qPcoQzO5Xz/vC8
nPu0Kr7oPTaDBN7NvA/o0nwD4JH8X3Fp/0Y5sTAdVKeP9elQxmL6mhcnkU78E7gR
hRmFbRmolQgJmh0SqlerU6z7LtJoZF70yvgJJnLhgblT7o0Rff/B7clhP/fqbcNG
F68S9FF8C4ni/zrPaM9LjnEj3AaQbeeicUX84QTP0v0m9Yg47iUfqUx6bfYfQlbt
S11TunyTYakuEqCewxfvZ8rAu0kXd4SVxofBWBcuCvbmm7DUjFssqSyqtHE0hn7l
s+fp/WkLIX2fvWyOomdGH/NozcMVFLViuuaVzUGdapdb0et7EsK+eEPLGn4Q2gE1
5A1Xm3BNl9NcYrXnMUjg68IMN/iztZICRrpzdDeLxt96CItdtMan/9wYe0tasIp4
LtRmsQWcT7U1jJn0VTir3IWyBjd+xv271kAbgng46eLqeKf10xTadEsrP5SSS7oZ
OMzAqOLhcUQ40oym7Is2OSN11BUKv0pgx+9J1H9apnWsiXtRRyD9tNwIfToCwhy+
2X3IDWl9Xh7lsB/mgxOJrYVFO6t4JC0DY30UUb4kv+rYTmmpKqCumez91Y+IKdGb
7SMXCzaNuVN/mCTywsg1o1l3SJQtg4xyZWO3gctky47VuWMjsFsWexHEXCopEmaJ
RkAzeAtMA5thg3HhwiHMUs5Oo26Un7Ezl5hRENlmguWC5fIAld0xYa19NKhRKiMX
brJj6iK5T73G85xQFoibz6PGLh5VgfjXozGP/WzcXbEHO/DtTdcSn/ztjjR2Z28I
ZChVI6wyEtOegtkD/BQhzOp6EgGNpUQ8HPsV9YEwL8MK8QMT08xhbOJUpjFRhGWJ
Vv9LAb7r4E58yrGrs+vre8c4IlYZcu4uOqrFl7yDS4FASSWtzLjX07/JWg43UXDq
DN0Yug/uq/YNcLJy8VxNXj33gIgDwbecfLRzqYAm+8pUtYu0CprgngfcdhXL4RjE
dHWifk/y8o/5MYrdy1M2jFG7JUSkEMR7UBFUyaXgxO24PUSseKZ5qfMX4ZK02sfq
VupIdHm3jGaZzdmkh2XftXoLdJc7PuTb8Xd7/MMj4GxYW5YyVun9k591kbmr8mwY
b6r1Cu6nGEJUEbD9+vGu+hcvAS1kAGe30nxWt99zBzveEIVfV4aLhEG1xzjXNMi9
bCyoEq4Za9/z3mdtPBoqb3zfF8Tc0a848l/5gZ924en0+FcMaNQeG8U8JVnayu8j
l2cfOKB1+XwKd6GIrQNUtLB4qfgutk9l+BnuEIlrVlNf/dHEBxDpBvELDzF/g0da
BcNEA3j5zVcREPL5vWs1dldnpOvtG30ZR6jYOKm6gx6mFihlqHUtnk1g13DfL9oa
MWHa6VH6gi/0dlshszLZhewyVesFvsnVmQZUIsDKy+UQuq19RyZ3Ml+vyXL2PdoP
j+Ae205D9HxH+oNFlV87BcMf2cxEEcz8+RkEd9704tsmhUdveSEGA5YXPhM7mTy3
gaJ4P4svIP4x5aiZK+r5EssmA7FQEdwp4y4D/7uCa1ZPKNJoWJr3vqmEerfOURoS
oQk5mazQuOBWXJJpwneAjHOiIgbi+IEpe15jHH8hYjMJIyTt8IeKJ0bFEiaFgmsv
KmSKZjVFmEWPH7zcqVIivS8HxGdeJGhfHlM4rqJ9XD6wXzpYQjNzTUR+6xRfWpBH
fFgJe+q3/h5tJbxQSUwTNqd4HLZ8F4TkEZIkJF6tzD3Sv4bDFxIgYDXsF98A6cKy
oIejK4ZwlEGSeyL+CHCqMYtVBL3VWwdjvNerP6FNJ3LIZmclbWPvNI9TJM3EVsA0
RCzhrIlp3txIjdYxuUBRTcX8W10QjUdOuL49xHXCYAyEqI7Bf7V5LI+ayZJnlsGz
ltJJ4xKFeyJNtz/6dZDEtGb2llqQNj3d8Wo3QRuqhCSsnsK+xuqDF9KI5BCspFgQ
dzzQCmpWaoipgj1335T4Gts50gB8y/U7u3DNl1iBu1SjntGVuInCEfqJ23AhoRBM
bvEVSlCBGnO7XGUphc9qxjdnbzSrn92e64NS9z1Hgz77qwN+KjYyBjJeBsMpsEVs
xdOLDnSWx3K/aNFFmLzYZpVOIfPvtUCDCGmH5YUKYpIVNPBG71jJ6WmtCvnEPAot
z8RY7DgX4rdTVYQLY6nQMaSFU4E+NjWA0GhJ6tUZ6jbQRLxbTaw3Q8T4nixYODv0
p+ogh2sFvwt/kuDXLzpHTPK4ArmKi0NqSwpGKmr+nODUCJhz8Ewjb8XoLSdnx2sV
YRjVI/+B34cXx0f8OpFrmkRWwE+m2YI2yA7yKPrQY0SSSuO7M8H3bZqqhIr4vC3H
+mQWtWTrdRXbqVEOn0mjNrmWaiNJX01XwsRElAUUvQq37KqP3d89hWtKLJOK41hu
nQDaz7fUhxSZz9/DscXkMKLSTDYKomxDucE+PlC1ULaL0ZTAlbJWlP38Pyls41jN
BpSYmgaVug8n5eEQ8/DiWkRah4XXF0oCKFQgU8BwNnxWrbMXWISIBRkYYX0HUQFu
AEOxo6uxxAOeoN1vTG/Ck/2OByqKnFRdoevniZZcJ13UiEcq2ld24HE4n0EL8rR9
KG4JW4VmelHwYCfl+l/XJNL8BwcHreqpTUg8pdbfDFCP0MlUollDx/zHjku3QMc9
G/QidEZrnIiKEORVqLXFj3Q4JUorQdwwimygAGwFt+K+4wl/iu3rMqxBEtOXHkBV
zcdNdS9bU+yxDwvC1TnHmnnXfxvPnv2sd1nJrlbKqs9LjrN77S0D5tI2/ZDr4qes
+eBpgNw9bJQxrgjJIkQW2yTa9Lu6wSdWwdcGHqVmTzg+22PhIjca43vvssn9m0Bh
WEScoF9wpU5gjyNju+9Ax2p364gqm8KX4n0P3o+0JBWerdfthlBhK+kFVmRQFm/g
bXUJiE2qAptrKqL6mUcMzlWwulZASdTSkQolZPUNsE4+Z+O5Dh0T2Sq5zmXT79Nb
xukspNApBdBHvTxfSYyxpaQc3NSFNHIpretqWqsqeQx4//NBywyoarJULroCtTge
d4ICvd9SbnVE8vFx6iswRwjxMp2UFOqcIN5fkKKZwzjiGQbPIUcZ7qOT49Uj+bWo
/8LFfD4e2P8bqs4Gg/SKnppShZcd66t8jFjLjHMYlCOoI35Q6P7cK5l3SNq9c+E2
kwj6j0E1Kfhnf6I8vPwsoWxj5tuW10oNbMJAy7plOTp8tKdkhaYYsGiyumufXmXM
0WOtHlDB1ozTQmL4Er5IMTVsGD5qHJnw6PkyzHDcBD/6DPPdHnu0uq3Lf4L44nBN
hGVLgt7F4Zyw8fHxQjwelO0QT6qDnoaisQ0CQ+9DW/b8VnDDSaO5ed0/q3V+Y+L0
ihqAfotlWq2ayNCX4EAqgd7fJiOoGjsoGLOsoKrcF3RZEcbPJbID3nLaTgMHjU1y
/mN88lS8UhJ3qik3JNGNITOqKpwkYhyzbq469qnYLtkivGzuqeGzd4mRolnmJEO2
eY+Vsw0uDDVZf9cJiZuV50N9BuGs6V35nj8Ag93iXNk348WhnLyeDXBOb3GMp7HI
DavJSML+npvmlIfsIYC5qE21oQojoJ4fh5laB8hzZ9V2Bsll1+cdIPX1Fs65tz+a
ST1UDa3X0wcl+8uaCLX6nzAL955MWs1TNesdRG7NjgE9DrDcdO8x/sUBEyEaPpjH
U2U7NKh15zEuCzbcdGeWe0086sQc8lPtQBjxP1Vg9CELtapnC2AMWBTci8ECpgik
oRY9jzdheFK4ynwbHIjtSCroJXARGG346bUe+0OwNm4sHGtzq0z6CJ7LliBidBZp
vbe7ltRZfgxmVi/0ja/2NaIf/hS6lSg35pPwzQL+Z7lCvAyegdIP1ob4hZgpswM9
PlGOivphcvWPD0oWV8TCuWhUlnr61sLlTeoDBqqFNngGlvbdlW+IgTMLb2MPC15K
hSaxf92OP3TQYgiWNWFWfVn3pnc7H2zxj4txuq0kzW7azhTWrH/HRDtfKXFRfaDa
oCXSRtqYkCalHw+YqWiDr3GSOme7FMZrfOndveNXS7zcIM0pX3qCSx/RYIcpxFUt
oBFDeBUTWiOweJl5Zzf0MNTNvGROh1qJ3+Cjkzmo5osodW6pPiOs6LldaSRvQkl6
u263lu210hDr5NRFv+c1E4d54JgeR1CWskOqEPzQQOLp2dhJEDAjFeL4mFLUFcq8
IrXFaUxUB8xlshW3Yk1ONqBdNUg2/HYIaxtbuRNl4G7H6hPUl3wPQW+BL3vmvYSY
JHId7KQ9POKS3tsasyQYXQxeAsCS7RkYFxvCP9LfDcKWdcRNEy41S0srUu4SjEUA
r9qzrEqdyKGpGuvF6RRi1kzBGKhN4z1sEwayYJzW+cFx+j7W6PVO+xS/jCGF0VXY
6EEwX+N7YfYgQdg4TgIL3xuUX6ySb6rgZBri0//z6jMLhin/s/3zx31p8uZA8+zs
e9vwPNYsEXpJKVTeF5XbkcsmPpIjnvwzeFwBMEsKsxYayR50SIE3i3v1eKiHPLuC
fz5sD+yLnj91lkGKGWg2StvPfhiNGimU7eTStD1bhqkIdIdixFgF2Ic6u/KAMJpD
fAOt8E63EDXFWrGsUwq0IL24EQ+wfXqmd19IlpEd3zCKcDlAR8QtdsAx5LpMnvO5
TCyXbZ8RCxNB5LlTBTec4hTuZlI5yLnzikO8hB9ZRZtFRo6QiBAyFyCiShnn6oXN
d/a/pUq9e0pLxhY9e6iZNXaCKM3qOJpuZzl6WJOCc6ws8Y8NxWnV/8zdG+cOSc/y
0Q6HygAH+8Fqg4cugiExL8c70E4adv0XrlDWRokyZxa6k1UtT67gnpAoOk6bvJED
6ZAg5bcRlnMGM00AISbZ+O5uKAc9HkfjgE9Cvg3/tdx/TfeyztRawcbIlvRC34Al
OvvpIEX2oI7JGYqQYEdojkMWWq7+AnHptbzy1dgP9PF2+reHUPQ5KKVbfzERdqoy
GXOfQU+V8WeNtcFN470hRppP2Vi9S+Oc/I2rYMdmHaJ401o+o68KS03Io1HXDY45
wyF6SuuyI/hPXuo4y5B5DgojMN3jP3FrTIexxjf81v/cXkKRs9T33H2pWnag/kCT
GWpjU1Z8h7QiiJU6QiP9fuC0bZowyI+cyeHGOw2Cc+Ni2+efSW2/G21mND+FTeOD
HFIEgRhYfb3R4l5WnT5u6wh7H2j+jJeE1cmYxDI6qk5zgN756/90MzdLy4lczPhW
oSuODmfzuOCEaJQrvOZmgwh5KHpM9NRBpXbm1Z247utzYHX075SQqT1DOy2Vi5L1
K390N6BpAHkX7YrNVmt2zd9Xd5NPA4Gx90RJ+Gsln03gGJHEs1TEly5gWkszpjX5
sNMALWj1D/q7+cvzYE2xzFMK1q93g765aEsWAaBEeWLXof2AdeJr2aIjzGQQBg8y
N1EEL5gLxWf7+g2WeOu8FYphZON8JwcdlOaquTznoofao3lwF7VgkiJdxPoIwmDd
V4CEx3rp1AtD8qrBYACJS0h+LoMqr91qvz4jaYxkEKeWuYRBEqPp46lXnj/sxIuN
2d8FAvQeKQJktA9Dy9iQpUjF1cf8WTGXlIhXrCO2AyAM6hxcuBQ4YwLhuFOE+iSx
fn/Jgm+Pd3EsfM/U3K0TiySxqn86JAYMZL7LsBwgWVS9UpUMDT4c37d13lIA5tI3
Ewy5J8e7Wc4BNvq0fRphhxrMaq4OutWhY2m/yOaPM3BC7DEGloM1Mu9TK5IzTkoX
NVwLaxUcQyyLx8Gu1/MAjv/tKKYzTbF52wKmzG9+tklrEh9/3rM5vsDV2c26U0zq
/r0V4RMbWOkpRwJNo/bUkzFEQQaD06f5VGV+kYvb7rVtG7ve+NkcUPmjjs7d6Pk9
tSInScrWgA97//wpAFqPEMy2cNckWee1z09Rff53eP1XW/5eK4mQo55jo8u8y1R0
YmSfu14ifA2MSRssDkIUsejVw/SNnjrs4VF/XRRdfXitOUZaEtdK02r8hEkb6L26
pbq2sFaw7WK3Cz7/VYgjH/zB5t44IIaC2W1Bc7yXVaf9Cout2/kTrTDFUVQoEhFW
Aj1jcEJGfOJyz7ZEDLx4UfrtD2gx+WhTuDLj4vdDxWMiKO78vZGy+Q57SXy5PHie
j7VILADU1ewv9ooMzzW9GvXGc+eUbtRFlNq3zVx6ZYUW9D7NqWtE8NCPprVupQ3k
2ZoJ2kyEvFXMh7F2YHK4yys3gUVva/1E+QcAxwWgf+/wdVm5VtXDMWjCvX0uFxlx
Wxh88laX6TGFeeN2elayZ0H3zDTbUBf4udK9W3CK9Qbn600qig3uh0Pz5iUWYrA/
RSyiSkTH7bRL+vIkU38OVD161sgrjl/Q1gRqtRIJu9SZdWWRSM4D9zECIW+6IzO5
Y4j0frLUtaM4UHWBXErSHd8LtbDxIJeqZYWmIkC/qYlJJvLutxsZfeL99c6LeKXc
5MQFmelL0lxVy1ccnDO2G1rkijoeFqeIynb+QRvc6kWCcFTj/wMRRnwEAqohQy+x
3MBzRN/Qzxf9tH9ukRQB05CvQiyoU/k4zeRvTTNsl5scb1lJkat91xsWJDzVnsvg
+7wMPYvfzqoX8UGfy6xNII9Av/h+l9OIOUN7egkyOnICq/rfEQ0XrnNlZsHD6gCl
qUQ9CA0RpkUxjQdu5xC9c9ciovXFv7I5ppgAy/lI9d9865npDQpMCRMcKR/LYaGs
xvjrWcEy488aAHTY0v8NGVKf2mxidQtnGK7AQ7vm+pZxRFfZWgUPSlDUlXYZzWYb
/Q8DnLaXGNStzR8eua7254hCEVcWESPzhA8gd7Iiw23c2SWr3VS3UgVlDxdWXp1T
rrtDkqkxG9jykrG1lHskcDI/W48HsBgLkhw97VhV1t60/Bv5pilOCRIHvC9qs+wP
7e67c017JbNAXVArY99thIzsx8IWGvDh8caRgP/k286MHYwCNbhgj1ccnJ3k2Aoq
BYTt1t5yiXbDQr9nbQozlMsJGBD/fO6zywVAeIoY9Rt17LeX0FNVksn/EyMGWKQm
VeRXAO7dG1o4335UmWjuypEpVd/aT+zUGyH2kOzqTl+o2DO6cpfeufEaLzH9T2Hp
Ls8x8k5JtKFUHNesnNh8nUS9SMxPovmK6BtjfzmskUX3x+msjzI6/VvGHZpDvAx9
qHAcixZGXV9okkfTXDTxFpczDykdguAktshBmJeziO50y1LAs/FUh4/xomDFvWqC
8U4RincgDD5IieusvyAyw8HHBHIgwz49cNlQjn6bnDA1qaG7iWWUlIQDMGaCnFyS
2a1YL0h9fKnohpIVYBTCmRJh0hMfs+MZzyzH+oFf3jTnYWInVCor5O5gfFrxQhW/
tp7T/gjaAtHViLekPcxfKEk2A9Ny23bWVmV9MbrwT8KfWZi1/bMhyEqtta2A7vAb
GebGziyqzANELTNcBpT+ocXmZWINjVZFw0qyv0RTsvDJF2iobgv/vfHjtO9wuxKw
/uI7C7JvKpUTlTkKpNwijbvRSZRZla5QNtCAx04JkRznlqmhY0d4thrUJeSkvbNy
1bxtiKaje8w2NLkMjo54yO2Rlhiz7IaOeS76P7kTNAFf/YTcGnhnnuxVPq6dc/Bo
8yKWGwicV7KsFnaTawIx8d9csFUfx0ox75KbpzsKEqR90dFK3X3x9n2UryuC3kBo
FGzluHrgMT4FHmS7BPhgQQfs0JwpPbpok90RgwTU3tei/JDbQueidWaNc1Jngi1X
wozApqvi823x8tHuXWS5Heb//JbLvupW1CvXvX6roLyBXv7v2xTXHsnMLPNoxH0/
pqpu/44/R7ERlYCEaFCAfP+D8f+B0tJ/Et2+WtnMlqjt54wJz74xSEUYpVhBlqrP
jOH/7vm+4gqN6fKDF2VO8hvzZXey89NAR7ior8SdxGMAQL2MYobv6JBBbgb8Z1XB
byD0CQ89zeFjtGi7sT9NBaZkDS4vXPqb9fy/GKAp8w3x3qAsJBjPex4M47qASUwI
Xrha4XgPaE1LBbm2HYd7lpZHjEGvoMX6MPNoJBp5RGw9t/42x9Tif89cDyzyY7MU
3LU2uTZWAGMlV4PPJQqmB0tuUBnYm2UH2h/ImlS10AznzFMReKVT7q+ADaS0YZ1s
O9hpr/SkYzoSCeRD7F7uVYu7ZnQDw4ACmGg13tML6emnEPoPEiJiaS6bdcYH9kUD
QEyObtoIxJo+Dn8czmrcH+X7jAnffUWwEyZf3eY6+eGzwabrWjlL8ieIVXRdCp11
J0DRNAVOMX9DO2pY2vglImujuDZ+YbN1U8W/dAoypPUXzv6DezWhkVTXc1yEwtnj
j2d9uS+KaHx6YiZVHYL4/vYecuJ489ahQg8Cqd/Vt6QrOKWS/V7JSNnqn8XEpYjp
vDTh5qffZjLeIRON/BBDar4BtqI06COyyi3ik8jyA70fy774GAPYc99DrTAou07o
p1HOOPPoK06fiXITZVNhbiOIKVwUq4bLo1IZ9oOBUq0C4cqeufNrLi+Qh73TwdOa
oO+5MRB6l3DEoF022zb++QKb2e2g6g5Ey6M6wEsHg2tXpccrT30+0srGQAqKjA+W
chxAKX0L+3ii6jVuR0S/elHPV66wY8MyWul6NAAIdAFXRQdlsta6uLhXAsobbjl3
4LpRcdH4VUI91LuuCEwsfFWNY0lFiX/hI/sH7tJ0Rs1C0m+Csm/yXU5gOPWSClIb
ugm6wYs4s1d/A8d4ltHiObzQgmo5v2J7IekaP+2w3oc/zm8BkU+NQqICxtZ1TMjT
YM8Lbtf8cJ9fQqnhXECmduwYtr7RpBW3YVW3ztNSn6KyqAfvTNIPCmbdDz6m0EEX
CHvzEU4byY8aL3ZsWdDwMHb4jBnxSXeY8Ag6zEjzKsTmifpxqHAHQ9GhOzzySKGg
T/0K2/CUDazuWCF7N90Hnnb1DgicoZDRk1xqAfgnKX6BwoxfMmXzIfx+NXUZxRlG
QCx10t3A63akodknO/kT8cL94/rCU7ZOSUwkIAy2971YZEfmK4QzrWG89PTFlszN
HZUNbUW6WLItUKEK1tZzUYNwbiZ5nU3pzDy/msR5CF0I6rdNqNkQrFCfCoovL3F4
RKgY6i845e6yiHmRB29CvWUncIO6HlBCpICp7FUNESJnJ4f7YfEJS3upvc6RX6cd
MXJS63fxnNUpaYYd8yIVxeWj41CFhFF1Wz9qW52H5eWwXK9R5mJnDZYiLDTCjVJt
+YopwqFBCInWjqFUcClHuuSwzoa6Ws1G1K3FRUq/e+rhGOYESbyzmk0GhFh7zrGI
09gmW98lH9NhwdvulWLr0pfC//gUlY5InOkPuhAMeqQE5UQyPK2D0WgYZ+pcXUdU
RSz8OFTSHAiouERWz1saiA5F6Feou/gyqzt8Fe3vMWNapaajobgVsXXjH/mVUKYO
EaR8G9q04K2Wk4Ghcu5KvClOxsHQ+d6NUPkx6XxhthcJdp6gixzR3nWBU5DzhhhC
qJS59bUusGMPn5bZGJ2Hp+J2Hw6i/igQC+uq4zyU2Xa19Mmf2k5gDYCmRAxSK84u
7WzzqvfjAbT+pZWixxitTyToxppE/3fBCJBeesZhjI7zjEZRM1uU5OISifykUpcw
qvfZdZAdY8HfvzSbvMyweDCT7MqATNh8QqtWvgh7y20hjMa/CaThEpENHmdGAPRc
lgkFVHWRlkMDTnFqPigts6PjdY/3KCnzUq3XT1/ZXuL65h6sF+iCeKjciPx93aS+
0X/UGTT8ehZhFOKtUyEYVw7r0uTZVFCTIsiR6t6PrKVUYaEG6R8AajDohhzc+jph
zf9OWEs+q2jmpVedzpRnPUwsYczgTJhcnxnrB87dXRHCP1bHAFyKNkbD4Hg7ORuQ
MA0GoWHfCRn/opCmf/UzFstZW5aB+eCKkylmfMGQ45tz5U9MU9JXvooRm3UA4/5R
mHl9ZhPiFMCw7hB68brj7Hoa4Ty9JbkjCrLh2Al6DVvsYbjTgOScS2yGGhfIwHVx
3cR+1T71yoKcaqtXMMBcN9L+d+xH/3TuagKMZ1htHPCy1GaRIDnOfR5ggeGeM+cp
BhyGmmD9JGWPZd/ypz2ku07EBI9HD3CKAFp97iFqEuWgCvb6oN8DcJsQe8B1ilFC
5R6jdDZrEkvfAa24gJIdGo6DG25JcvDT5eunh1tBKBVaxrqroC8CHeRX0NLn9Yjc
pvIXZUNbV9k7zvpfPVrdaI2I78lnHT2c59WpqQkHwolhUoIOAhKI91f6/7t5Xe7W
FuEA4PulaJJXkS+1x1f2FxjVVs7m8NsUfQGCwj2a9F8tzFPLYCxP/pSFUZVF8bFf
cms4mUvX7w7VfEeubWFNHyzAmlqq9W0SxGItOMmxLOSlbnjbxpL93/546K7DBZBs
595EOfQI2aLZ74GourIBC/pQRh8R0u1k6EH+iSfuIEWpXhY87qAOAgfuBHAnS5XA
N4HdeYfcIgn1IxlCakmyhwGPoT/my+dh7XDAsU40uyYIWgtNC+y3peIJi6XX0lRs
e3MiKUyfs9WVCjHIgaPBqEMzMxpGRiSbgM6N5WvDF6cnXU0ucD/mNiz7KOJIDXoQ
C2z/8RLlzQCxixMs6c6O8F0T4omCKEXbPDNA/qCohlonaNiNlDdPCH3ALt38v7y5
veOAqy/vE5talDxLsMHsqNN+ueLchOWr10K4FS5WOSASRWM1jArkNxktBXEVBaru
cZRFZPaHFegjks+Moks2zxMDIkWQiFerpjVyHYF/zmRdHP+9z9DkXeq+3NBwkF2V
uNHrPvk57Qsse2I2g2f0U8kYAIRm+XiEWkj6v4qm+GxZ9FYWXy5MbKBfRt+vo+BE
/4XrrURZhPT2pSbkNtaOJzckJZVN/7yMGDNz9MHsL/trkRffnCsIDJRxE+6F4l3d
WsCelrv6CX/I3BJC5K1bR4157sBjEeBa8f4dUYGZ9X/hGvqqG2bbdK+cm0c+ZSa9
RCqopgSSXo0tv3ciyawvS8TpXvb1GcEZOGIRbhZH7zUdnAxiyyJH4zdBb1WvkjTC
NVrUkicFNuiY8V457WJCU7k5eObdsIf8d/fOVQDHmOGQvQbzkfH2+8KiC+tpcfKk
Uk6tGuBDL9huvOlLirlEYJ/eN2lRKfjQsxlgugd3yPOYhli6XzIKh3FuXq9tI0pC
nqS0ML+zXg+qZ9BGUrQsJWsYP90pbpzKeThDVf4ITL8G2EvM7qDN7DUzS+J4mvkY
h51ye+Fjwupd3BiwaA2akIpjwxM3zesJ0VzZH8i38XBZIMPthG39DC3527SNqEJ5
/whTc41l+v/ytJaUoim7QEJtcCnEdz/To4/tnCDMnBK99Zos/SD7EQ+l6GwGrQJ7
mmK61QLv55OygUPQ5HsxjiVrQje1iwviAQjqJmKHBUwohP4DKfT3cXROuuyE4AEL
xyJ6Z8jIa7F/PizjFLLJDSLP9wZLrueG96zlwQP5pFXUufiK20YSHK1swl81LB9h
0xAlHKtHRCDiPRKib7G9t/BNhqQn8A8gZdyza2Qr0ymoLyZ6/BxhwAiwLuPH6qhx
bY/CaqUNW4f4ed/lnle3quqvxDmyskxU8q65lZCVOUQ3GjkJNuuXZAmXDN29DcHN
WSq1wT/R0kmJVebV5uxnFrkWX9eB+Wse5dFT+0cGS2stJrYC0Cd9R7rq1VzD42B3
QDW0hU7ASy+PpZ+P/1fvcN7Bcgr7c4duiByWcg8Te32ULIC5mwGA6ZW8ms2OmNUP
wddnG1k1kWh9ahuh/h6UEVxoqdImDPHfLqmuxA9zApuP058tZqZeJti+j96FFjef
13t0c0qFNkW69oQ6C3VGD54C/n+vE85rQU71mIYnCoDKe4SfjjdlVbp0bA6A2jq5
lmc787qNCKnNsuV4rR/hK0xxoA4En3JUOaNmHDcxzTHMhRVGc+PKtP7Ak0CgTEgw
yXt1ZbBExgrCey+2uhK8+nwpqvyP8lNj+8IBDv4yO7HhR+AnCm9+ttEmkIfPIkF8
EwVZywfCS0k9gbgIkMg/JGW5GcoJokVuydM6Ku6vq1poHSLBsdpbVIz5ZcNbKsSB
EzWM8NjHz+WpphmJLaN7OObdvRs+W61vggF5bny3MUUEAdtmnHlhEpUYtakwwsyw
xgjGdVZ3zB22XOhqOVsm1blipkjJYlpbJj6DgPRoQl0fMY1GCg3rCMsElP/CQq1M
vHTQv24NGZoE5EqamcxQaixpL+94SlQ5Tm09Imat9MpZY8w45kAIMpXj60Ums0QH
GhIreFSsO602bVQjEwo3rFXx1BokBM5Hc5cyQlGXTVuLA+DDKRgBLVtbA0IfEAv5
UlSd35tjI/3Am73XUd94EGQAenrB1G9xP1CIIU6IWyf69UErXaDyIq534KcSo/yq
qVuYpbDTNHR1swfdHOJqaYx95eGVb0+oAaVUqOjsKMKusM7GrTv54bPKCkmjnjFL
w8rtljpOIZEqVUWJx2ZDw1IYBe00LfT84I6DCYYDjjj5Aqf1jSsLL5x1BUlxOLnA
kQQy5Ycpry+sUXryPDL5Q+5Q7nJtPD3sBpp/WSBt8ICbJFi9npoXYtXzryvn28HH
sZSLSgspUaeju81If2Hrk7OdNZv16CAgnXEy1UjkBzGc9JvNxeSBNqKbGrRE7v3w
Rc8N8JNOWx6Aa05J91aA71aR55NayyXvURYP7SX1ryy+m3V6jMKu95F/uo+77wUI
zE3wu+QTflxj3a8oVT5x9uN2rOnVXHmW90ajiBOkuQPp7PEebhEt/Y6kgpLtRVWD
FrcF0DAb82gAc6Mp6A9K6VR0o5R/L2IlVeSjIVuh++I8QO2o+uG5c8Nf6eOVZrnr
rOyf8UmW09eKmxmfhvtMERuvvtOjgCWmZZChZxF8WmBayWaHbM3fFnvbNK0pAXa5
5bNaUJXVSAnokXfliiPMK531Pi/fGhlLMJNhCSsv7whUsd1t56Dvda6yw71rk3Qu
WdqzoUd1PrWh4mHAupSrCnNofqeY48UV4me7Dzz7OskQAVrMpGMw6G1w/fCAnZuM
h6CuojwwStR+TKl9u4flE12jqrA4fwU+L07HdSAHSI2YLqEfQKbLCjKSfq87aokL
IYzvFMkfp2+8g4KjWPFT+sUBJclYq8m2nyFNRL7yMjbjqe0LzcHn0AiG3rWo69Lp
g/YXyCv/toccTqK0clI/gB2NrIrzT8yg4WYy+sDXyS43+dlFW5jyRxyRy2Jkk1ap
bSZ14Bn0uLJr9RG8lrNvzk+93shGpUPE/apO8/ymPhMX+3I+SYxyhRa76HHSUsln
MR+99atHSoVKG3NZ39E3fSc0H6++SGhRFK+oaILtuT1F+mJUmXuvzxO4+xbydm8v
0y+LHk/hNGQ8uHuXfaAygFTNakELmcMiw2RS2MTBjEl9RBA7vzOkMGAy4IdiwuFG
K55toGQBORrsOu9DoxnEr5WhCz9nje3AFHvdOcP23CEx0EaXFEl/bOcR90k057li
8woac9RSjxGmIIgmxUJc5CQHFzQlHQwiBJhnDB2M+Wo8XIAzV/5H44D3hdl4eJyR
eXco3hXvQmPGX7+THrKSoawjBQcnWeb+QUZCSzAWB7oxJyXTmJ7g8BWS+LQVB+6R
sT/WinJq3sY85RqfFdEferGZW43xIM1BZ4buUJmd5LHOYGyjShJsDSlavYxVUoW3
uhx9LbwCIdhVvPJO4QtV3VJ3VMFzgHvXuyjdiFc0TxUhe9l61/tiEfqMkPr0YH+I
okLXwfUaJCvRX+h4IEHwIkgBo+4k6KnlmM8Y/JMhVJ+LIzzSttc40sTdogJJHzz6
QdhTlrboVJ2Nzy3Vd/7OeRNo1NEh8Cpokq/d0ZDrhWuqoAv+I/YbeyGtYZIRLWAT
CKfvrEs8XevrLMd6g18RmGBkGatTlJ+TyGuBlCMaW+s9Bx4dZJULaGySnG2XVEip
hxxZlp4F6POmYM7LJkFXXTj01dQ/r0FEZAc/F9JZlrapSysUPqy6A3216hkxQari
LvDsmBcim0DAL2DNLsUq92VWDXwlTUsGkdUONM6is3lJx03+XA30jH5yGiuqMzyP
IciUEuXs6nSGpTC2BYb7EJAVlyRiIWuzzgInoU0N7xrHYXA91r2G2yZkm/de4MP1
3jfMNHu1npHJd0ORkUB7G0f0aECQYxBiOalEqQigzVe5CaAdyhJ2tSiHMrqTnwq/
pSNLE3PODxdbiDblr8qRyO4xHfZ22CC3HxxBFaJsZT+TTWX6itIrpgen9i6/f3QM
/gST7wGULs2EWgbhzdAWECiY/iBuwUJWa7zymfUymm1pk2OW8gBUr8yTlaxzKzu8
zQ/slBbmD7dYB4/8tMdEuP3XEkICz8rNUoSqCXu47VdcbtLrEIaycxUkK/1qmO++
uC7YvbaBufExO2vtlJsckRxevUEnV/q5EMNte9BeZtobRtMLPabfqGsn9SegFhum
p3JgjV2NqvWJEsv9IQam30v34K51NkKa9Xxk/6GCTfXu3pDuHjitAj3oWbsNGLhE
x2Ey7HGVNGGDSGwF6/temgsijuqTBuJ2uWeycMfEeqdmqLbXJ20+ZcBgM2MK60mG
GiPSeAX+PASCU1ZRTH2ahkhDbVi/9jdIJyIYbv16+S/FRm2HdLGhRt0DGicgOc8Z
vUp0cOYMcqIJiPFwRO/NOL5mnFH+zNsKjqQE0tYBmHwIfdLBboYGvZIzBW4+XHk8
EaP2t5C93SFX0hzoTdZ5dtZ5yXy5rnhBYaenfZu9or5XjBhHbThJhcRuYpx9uZnq
6+sItOesIU5RV3wZy5E7q0aDm3CRUwRfkzYGvwv7zvJFFGOMb3RAhUrG3QP/eQ7g
LGfbAt8uzjLbXR6QIT45FpIMLWMXtWzkiQlGWNph7OEiOu2rFxrcxxRwkCOr27Mp
52f581/t6vxmzT0UblVNdite3LHBu/A9ubRkONKpUzkbVIUlRKnnvhgplbRwGoLY
srQNL7YJVqHgKVBSq0JkTvLcmlklcHL52hHaN/e+zsRFWx3bXCQ8YSEUIT8IyLSH
6j2sYTNthDurf2g9Gfhv1IiiAj8f5jHlQDA2LZ2UuI5pMIDzqbPfCoBjViU8yF8z
lwU1azL/QQHoBsofOP1y8b2IVHsiqbKCc3p1BEJiFY7E2SDJH1XBLDXDhNf3+4hP
sQyDFlZytKq9LV4b5QxeHzdonqZMwVjre/l6WJdrt7yeQDTVhOdcdJtTaBfYNUNm
Jbh+B5U+njlp/MNf+7lH5JCqBpNMfZgV+BhZAa+2IzBetUMp6JtlnnfxH0kCmWZi
P2NE1PUy7ngOyXl5CNELI/b8v+x9lLylh13D4x6GGQ24jqrRWCqazfSGfUDG3KWa
V8Kp+WJJd9Ze//Bo2RD5wh/AyvDmV3xhUBGZEeeMGwfH4D5ItC/OqbXsaNSSWgJf
FWorNfcivVONYbBpHDwQZe5rhqunStReYAplyx1DZOpmzl0Nrg1rBO7FxrCM8vy6
scnqFG2981xT38a+vXDq1wHq5YN7fY/Sy0TB0JyfONFOdgxYIeMTvKQLFsEyA73Z
XZ0vHwaf9Eei+0kYdF27fk3ckLeH8pq08e4XZ6fau3bOiJEQT858jeowMKJGhuqa
YmHDNZV+HP+4x3uQbvFGdtI8fc+XRJfQYD1KAhhK9NvBqA8mDAnfGMlEhMKpLgca
QS6G1jOcphqcm5CSD+pD6s4vrsvH4nF9NWILQiZcaza+loua1PkcGB1CnWBzzA4A
e6yrI2TIdF2kIqC1pJNPossoywuuVyIVByBOUb6sHmihNAqjpDDz72hh1mDwFP/B
4VmSgrPcZ+aEaOoZyFyBHdf1qIV7aAtn2+09C91dB2kJy9XbY3Uj8xYXkR/w9D3m
Dr+Sv7nVt7UU1zjaGOsRUOEvkPNAw40JTJmqNs/1jLZgkH09OfoA8U5dbVSirjpt
V8almKqtnfDKaQ9qcZ+w10wYHPLAiBRjXa5OeKj2IIGSWBmy//9xEm5S6Xr5++zW
5HH3snHkHf8fjgeAZ4nhEGaONfeQvWm2RmqxCvE3QfgV7o3ZGoTH2UWC3EoYgJpQ
HHkdPJHiAzpzbYOSwbmEYaFp7id56l4crJaogUsg5BxD/ThDsoyBrONaGHdpPYcd
vKjZEKQQEGciDOJ7cK64iiGD9RjIarAurDBWypjRBWBrEfWDE15FSpdYeX32x7wX
XcmksVVZqVkg66k1lgk/xXaFB37yfYxF784wmioSXQBVZDEAB++qdO9q72G82WxY
MPc/3RXc4coDbQFwP2i0iiXXe+J/a0r1X0h7O+REc4mV9j6Dgwd7v93NWtY2Crlc
+Fw/6PEKgFUJCwjBTb5fawfgiruUhPFm1jV4XsZXM3o1M9rvOdwsQZiKRT0GNU3Y
xF1ZeO0Uui5Ph4/I4o+75Y+PP7Aks/zT4HdWN63eoRCeUdjk4TM+bGIub2lJCdts
ygC+cOxvVJstPFMXSGOrMRPvYi3OnpXbicTX8uc1TI1Q2TJJMyqLS8lz9fHdmKQR
W6fwBOx74uZs2ox3pLnCPbYzBe7q6k/UgpOvwNrc8+WrEXpONSy60apdkD2fQyOV
a7JHiULBU+bPaFoymseUCTDxV7SrcM38VA5slnCqXQ95FeICD1XV63y5UXFf9EUL
HeXNvfxdWWyrmLRGkAXPqn0xktH9sWE8QgunXjkiiqoJz162PZe43BYwTEkdPoXu
jhvlTz3SAWupGR2XylrM+vDzJ0s1yEALx83/IoYRva2dOHX6dMcDL5tCnFi/vPpS
OCXM32ElKMcl8AsDZyqCdo3i+9rPbs0anM27ed9JhrxKo4yj+PHSbUTvfamHb0T4
tJEWSyCYYBX1n6UX5grSmS64VQIqZlA4sDckA1LIBPD/iZG2UCkWIpWG6aTr2jFl
REPONGpjW469pis9rTL+sh6C1/AspuZfVYwh2QURpUkDJIsKXIexe1b2InzGOtZ9
NmEs+iF7aAb9EbkCpP/xMUYQVObOJGwwDHpX5Ei08KQag2U0JqdNAcdZsanODoRd
A1pAs5LYRy+iW6KQim0JDfFKG8DopDq/17XvG+5sijI0aZlWngu6zjlB5e+U1Y4F
2CAvxPW1wBpnshm5BqL97uAgSwHf03Z4UwpRLD80dEzqBkhUehnMWdYoDQDtOgSF
99hQ9O5ykRxMsLSJXqDWKG7bh/P9PUclcHPpdlfQyUtMss8nQ3Bg/oFjcVxNB3j8
5ToiNYINl8O3VeLbX1q2f1lOTJ5IQ/qgxUq+I+WpzVd2ARmFgvlYX67o13NjYzq7
CD2Dxbl5sXLz9JTY/yKy4uf8yNpQmNAu+kYLViiS6GtcKpDou3rsifZkKDjiVKIH
LQGB6wqkM08NeagzGRQn5q2QhiQPWgp7j5R58mBUfvqO9wZRJ6WcqoPqc2J2hVFw
GhSvjSuwW8VEMWju3uSNOOXdsn64tFX72Zp/YtL51HQtMa0JxovPn1+n5tSf7bRh
TR97VMXcr/LjfZYNinwogoZZBMOFQmXny0MsucZSJct0eDLsszawANQ0thxzmwTB
4J80Tz+slAAZd8zB63uoq8ms1PZKWXraNa10mPsc/3zk0dr5Oio74JFTleM0Myqf
RzOQ5eJsynq9RwMxb8qxn/vXPMNbynlAcURE8vrC/pFx0DflNDqh5Rjw6/CglmUw
QTFR9AA5hmdkp5F9zUL6xrtbwYWf75zdc61II0rRV7pO11gIj997qmpP4dt+RVRC
Qqb+IRHBc50bMDLQvNUDy+Bkxvy8xjq79gqA8Wwezmptr73jaWgVYTNsUmoiGZxL
Kn97fxOmvOwl60o2asyCKBiwzN0LoAhQV7hRLG5AujVK0xDEz4tj0bf6P3bxgdOG
ZQlXCMHnFUWYTg/vi4J72OjBOAp8IiuwIVyuo2hgcDIg5bRqYraxRrqig0Gz92ey
Zuxmtdm5tV7eBwQnqv1emdr333XGn4EpZfsUeNiU6pT0bQNAgeMpihEqn7KZvBQJ
7Qn/0rwh2vpTXOFziq2S9cjDuZ6y0eectp7xLIz7rpQ/He5mw06UR+dirfFqukZ9
ZmrG3QsYVu9vqCKkwg3kBVgkwy796SNS5cbHzdXXj1NFBwv7sd8uUxGDMdHatUM5
/sHEZdWYITFFNrdQJfRxtYcEziHZMQpcn8HC1HbU/bCIRXkLg/tylnbDGgabToo0
twRfsQXRRa8CmSjZrIUnmYiIxgtYukF2d7lfM5ucXdGxGPFn1HBbVhBUeh9rU9lV
PigtryF6bYUVOWG95A775+0bdbf8O8D5m28G7LybLkwZdZoJmUnnwLgywnx0tpwX
Rf+FImsFJ/GOz+LLK7qkg0En41ACyJ4w0vYAbXrzLuWJe+1ZNODcPBg68qzI6rTo
k9HDPsqLouD7+5eSoQDNozPd3gItu89Nu54XMg+6uetPflN6fK3J6IDtTDYvPH9a
IdWrNDjtMC5sWAoDQJuDPs7QMTcC9IvHqVHQPV+lN3/OZ8X7xdWpPfCAXRpDnnPs
zJ8OECAZ2k62P4UlCiNFlHJ6dSw4XXKqxAdCu0pRmWwBJnfHlDWfnbp9wZQ6xFd6
MMrirlVWf4mL/tMYlmwfcH8YByx2DCmcKh1ZSagyLR5M98vU7Pv14sgpED9Ss/sY
nQ0MkF8S4uaMbJ6JV3uLCrIzW3LVvb2FF6hYdT1GotyF+bS7n5zMAkxfYoN/08/2
uxsm1V65Sw2OvyXBJ3fQ3LUJC96UplxE6Xf4bjBVgoRuX4GkWezOhm7kgCUB42ac
9ytf5D3tosaavZFGNPWVq2Aep3wvOcHcNwcGmCBKPsztMNADgs8lmFn8OjcIMtA0
q5KcIijoWb+/4FAeo6gIRKSIAsbfiBDHlb6r26gUz7LaKY163yEbwaefJ4bZD9Nn
AzblXfAh7JXc7OYCZ/FJC65k2FYfAyEDGBGX8u/sScVhUiv2CA7fM3+LeOJyxSIH
x6fL+T4ZlUl1HRoECAHum45qYRahMmQSZsTqf+p8t53eo5h1FHupSvZZJBEOQ9zm
/Wkz7hNV+JGjbZfmTcos52oGLHbdyhSnnQdfzb6a7fbCh98pkxy0Ny/N9urmwHG/
tRRPM77NrOcYmZW2y3skIo75V3sRKM7F0pEXOFF8CUnRDJN80d5hzQYezWKiQ6gW
iZ4zESoU8p5OX7MgynFhMbHQO7YERSoypVd3pzeAEgYbuwo0aj63rpcCEGxTCuCo
U9QnltIvo4gZb367d13cG/XD2tuI+gFE2CBOOAM3bYUlT+1y5jUNRWMGeXA9cc8c
kpOq3vD3HXresuDRyf946hDZNkdDLTxQmpjOHyE8gP/ttq64W6CHQJLpJLDF/VSA
0xjINXyywdtbL5cYceyKOBAXzw3b//vRs4aJNDJiZ0p2KuWrToWjKS3evNgeBfR4
mT6ksoPriJC6QeMtrBZHgLpiEEQRbYuPC3TPd9aHMLQnqGPdzZE7k2M2hzmmzHrg
6lCspR7LauolgpwpQUWlTchgyWZ9o0A5BaYnW0fZBbzE9tukfLj5cX3p1Osz3gQj
VfQyVdoxih3WA0ClmIB+sVlWDjap/x65qTV5e/QEZbKizAk+9RdIu23d+eEUQQIC
Exk/Bl37tbW0FxOfYWOU5eNDOqosVkFFTvcm1P4p+DqNdy6Y93bP6/9DKqRAKSAa
Ud6IsNYZqZVscmB/RseHAAR/lub1Q7/k+0nAJC4i1ZX4l7y4pMiHnFO0s1NNvhRI
urSrGtyZNtgtmpDHKmfluLx8zE2dvqnPuBpJYTUeH9SK1C81MJsViBq2NXV/FuGm
vKuAr0Tgd01aapg6dPjEsxdVvjJBSw5lP5A+DCvpj8JgOqf0ivR1jflXhRuOUP/X
Dw0BoOHo5Q/8/rUCp8egzA9yiZ0fZayd0DYInJGgY67CeJxWb4ejKm1sqmNdqOY3
ywwsZbGFayrsailhhQxIR+TILVoGKDW08MeByYmFlarLG72l83UK485jFkVP2TFU
XAQZLF2DpQreVQoTn8G02F3eU4cQp3CNOjdCszVl9IrEh9S4p8WvD1JbybrYXAdP
0Glys7evng7UkW6RnPxMGeSpHHYsKdg909Fx0wSo3ncgHF8NluwRSniJsiKkd1xT
hOHvGvbT/EgBPKEHIRQApepfO0WSFKKS/z3BzVQicgp5bMpJdwMafddwZ1hSokcS
RD6cEjh2FmdvJsGGSZWGw6JTeEnW/lFSMVkX7ORVCK/Qu4ECjvGUkKddPSDoBDZX
01BayiALn3PlmwhqnUSGbUwAr35xhrDNsfnXCQKtvUf3G9VFZ+XR3kO79tKKF9As
3Mg513eSWAgx9vLe0+rE6qwkaTWL3vR+oe4/C+cRKlvTUIhdgd621lno13FVjaD9
gX+javNrT6znvOrhpjvt5grfYteojg2AGOuGyVc2IdcQ4rxg5+pJYROmqW2Gi6X4
sY69IPk5uL43ccPJYx7F4r4AvbGXcbB4eeCoReBecToAfPx5ENR73QpFymjf2vBi
zlCihZ7y49aUscqMs4CaL8ns6yMDqbPhFAEdzjI5F6yIrJADzsB+0xUM1KpswvU0
MQbZ3FtjYqIvGjSYSzlJ528bs+Zt7oNkCLz7olZ+q3A9C+7wooUt6so7Kf58LhRB
KnbRcrmS2HpfuU56UMKYDY0ikrH3ZcF1yg57oIAu7VUG/dNtsaygGyWpboJfxkcU
ANnUwBM9G1waIPlFcTBbk5GnDQSZm9AZ4O7ChpeNaLEoKENyDb0hcM/oDd+7P6qL
2HTNbCV7XpF+gDnsjeOlgntXem4Aob/v6PyGRcCjM3LfyFbhZz8GUEVZ07z8Ydli
0rdGHav3PNrwi+L/Ft8QnnovByAppdhQkTKwBxP65/fZUOwnfMQWDw9MB1/w4Mkl
tMuBuPTVzbib/92YoZ9pPSqhH1W3pRhx6DHv94KsAyoYY0XjV9D0SC6KOoHLe7tp
NV3W29bdtF/GYACUQQArbNsHlaSJIe7rEzkSn/0HX2SrOECBVjdzGeDvw4JuYbCi
lETu1Hz/0DdrXeMLHX1LT2X2HOUH3ee6P5jVCVjKXkC8WJDUd9iohb24lweGwZNi
pzNxhNyxeTPk2Lu2dAb6eBlaxOe1lDz9VYzsEsa3bevDke1f81ZPq+LsugjGSwNW
5D6E8027QCxpgFb/v8JbZbk+nYVbXN8fhRVi37rrIwnKDBd+J3wC9UhplkCf+A74
nPn7j98w/oQUJHT7hqjo7g674U6cz1AFBZKbPvfvmvdV1v/iNM2W8VI1uVePEFPl
88ZJ52VvPomstSawH1UFb4BkQGSSB4TxfIBzTMMX3cOiNYKe69RX3pkJcQL1bblm
5+QS+asqllSnJtUs2wZLXaPQpNE4X4TUSUXzcF68wCVkN6toStDkbEjiieAuAhHz
qv6upE0bt1e3xFv83vFKFUOTRtkvqH1SGMBkuC45HW4KheUYbT2KqqXe7CUpmjPL
NObwc6ao7/5dqMxmItJNBvqRiH6H7/ADF60kPNkgs+XH9BAiDV2R4Ih8kvfRYf/O
kSp15YNDImbU5RUZgAn0EoWSHWAnt/4wwzyHBRFnZQ4DdEFh8SvsHElv9wdCmeGD
UfroU9udJ7tcdRLXYD3twYQFlmWRjXElryrl+MbWrh8+SqEACgbL0ph22BG1g7C8
gtGDRWvhU4hX9pVcYUEsVVQv89DuyKzjIz/ahcFJ704F1dgS7INob8w09o4tmbBw
Y3UgJLGH6V/bSqARval29TK/GZ8pXG1GUzeDBpP1q9UQsWtjHDu+x29OuWB91lL4
zJXtYxsDbR5qlJ1OtpvZjuRrhFJn61fZa6mMy4qUn+qtxL6O7UBG8IUZxTBwORVX
GiuJloeX+7ONYACMJeYitNkK61d0yaOilxNHy9ygAE1OtmkXYjxlUzz6grZd0ZQG
y/cAuzgy969vXvmzsCIYamcdANqAmOIs4yNQtn6lcUEsLzTk9iY/FpLWpH/PIF88
hjS7J8qjVAiwT9g1FRf4WXRFGTrKO3oXilBe4iXYwKEQy/u//TFIgcyDHyzvr2dy
G6ENFd8C88+JBkTgYTbU4QybhvkN/YTYzmsa9rJ8eReSus10OaEEptuqhQKYcc0+
qgbNWAmrgQqG2rCEv9RF8j6YrP8O38cne6vNOfUSmMScbuM6MU56r4Wr2B/GG1Gw
Q9xIfoVIK0LZAw/Bu8cyuxXd46m0FrLgvxsnzec0kqdGBwkQPNEUZ9Wqwphv+QS+
2yOtz3EDDoFpXHPDMPbTHYkylzdqnFSe8vw3180hj6BxtNIEyyTP3E0vIWijoMr7
nijv1zVxdwg/pJqeCT6e+guyuQuKlrOiF5eTCeKGIsdEzzNO3mew10M+cDUVyIWT
wR7PqIzhQhJi+c6QYOxZn7SteGjMqT047ThbCUtXZLABBq///Z9P6PAqMuf/BHXo
xsyfcXuqwSxRtFzG5IaXfHujVwj5Kul1MTAIziaNi1DbdKcdF3/9miXeE1NWi2vx
QMgqQlWZQN/7lvPzH5Be0DQbJDgnQZxxaFl1H0n3tzOazzTbICS0+VqsN/8g1q4v
bKF6Iv8Q+ZAATozvUC24qxpXEUyHmdHpfaw6nZCT3RWRrwrGWHMMFv/5lIS5NzST
vF4CPSJ5j3qMz4SiR+UIrmAwGor67xocFltTAYlVM6oix6dqR6f3YeYU3G5vRDCX
1+dWxXYNTmvJFQ/UPzC9N/Hmoe2N4m6Y5bdLv9pEGGk8zuLrPXhHuy9VNeDCYo31
EoEUfAM3qaSc8hrILDKx+b2EdYPb22z9lqDkCRLnifGME1yGJpYQF3WOO9kxmRVK
tuSKevtGXtI0i1dpXrFqMagBllkKfldMqmbkjyZBkq48csSeMqhAFp0wHwt87mnk
OdvLWg6RBnoKBfv/T0h4RLtcV4h8LxDVGVOv5HlgPxqTrgaEifNmurB/k6BSuspN
P3GIb3EwEFPfOP/0EWAjEaLzfLjXo73P6408cCJ/nQcL0pjHQ7n554+9o3JeHH8x
dYynnZNbXerC8RNaH8O4ICC98NhPDD9Vjz8j8EAtMq3e+oET2ID7lQJgcP3+BMu1
N2lynQE6oKuOGdcHbBKuTcqXkfd7POWLrpsRCPuY8IzRUy/wosqpAzxdqnrS4d8l
p8okPcueiJrCq9xGpXoSolODDT1biMy18dCgIOM+RYxjfcz4w/ma0LrEh4YeAl1n
RkwWzbDrJGZi9gzxrRAhoyCiXE/jc7fS687jJ4ckV67ssiXaGLYGLtmkXlAPujoB
J+1Wfk6kocZhlHN7tLoQNlgPi6KARLM4h6xUpi3YidMb2U3I/35diapnk3b4MN4A
1QTcLnyd7bRRPx+PuiAH+ZdERRn7LTIrlNxixX8i6DWZL5IdxAHwcKzxvymEvbgm
bAgJZaiEhosZffc+NR5Hc6GqQCzhGxI1TI2BI1FPWMMXDsGshtHhvukyLCHY9ibu
b1EeJU5s829Qd2kNin8Y3mm9Qxo6Nhg+9Hce1MKa4J1g/Ana9UxV3ofL6ds9reXm
zaA46Gy5/4lR3ptvSqr9sxf2wqLRxnX3/s9K+82D52I2XTVUa/OYuABpx0rUt4vU
FfXPOL2AL7RLaooU/poMCEGu+EoR6rPn+IImu3hgb6DPBUofAa3Cy1Eo4UUiGwsb
wgrm8YpyEB6DWWOhD3NILyjwaV0h38ncum3vLK6F96NsCW0eB4uvERBHplwa9V5J
J+V8fSXN5w7YEhU5sdC3SHUBx/uiEMP4tGdowaef+Upo7QItDpbEF61Mz215oFZe
hWf7ejNUP2EqorYvPVsOqTm7hU9X/Xi0b5ohv4t9UHmCMqVVTnDcNKslvZHy+78g
R5ZQz7kp7UXUtVAGbzFYMciE3MU5bGTvvq8SvRiDFqwv1ZAkGpRMZ27mHGQqGMMq
AF84raQRpBwqDkDe4xvuKcMVwLDPV5T1bkBIlpLMmLuoUxm7edo4xWwSVosJhJXW
h/UT4ANf6jUH4wxKsc+oSEuIIo2qvq9UiUOAXrgpW3hoN4M5LbzMihF/4TXNdh9N
CdcaIC+fOWgKN+FvX3ILgo2n2+KwM/H9Go2sLMjZrJpOzhrIiXGd4hSc3hqH5gqH
JrMpBk3Bg0SI5T9Uj5JQA1Zn2/EeKX7uv9dsDRVbTf/LfjqqcE1mOpfiL3Wtlw/g
RyhW/8VhVB/IfMKblgYDTiFdH6BpLNvNCJV5Zu9ZKcHNbUU0MOTv2maB1/C6yAh9
2G1qOpZlKg4mOjWV1EKJGGOaTV63M99c2xlgn9jPvOXeni+z7R4UieNC0KuatIYx
Zg6HvsljWHD60LX8uJHNXBZ7R6c4CZ5gqjBdPFCUZAJbXoiZvWopGmYYQcJxT/77
aY9aB2t8y/Sq7pF4OSPAWWmlGgo8U0oMu0SHDTzq7FoxYM+BGAat9J0laiEQCquF
ff6Ut3e33zeZSCCaLdJz/2k2JuGc22rqTrJcQltZenVHOcTCPX9SWMIc/LECLIlx
hujXL5g7rrHbV/l/OF43kCfkVqUxu8PiDBQvYPq/borm74hsXysSoGykuNL5/EE2
vMEonHvjkl/nKBlO6Nb5NG0sFsdartH3bEwLEgF9e60IKTZGxXHcACABtLx9+h45
Sg2Jbcvi28LzMqVSi59Xy1VoYEFpexKLeF2h1ClQpHMMOK+AvOrWhlULbCv1mgkR
hEPwUPCBiDXM212vaM+x3G0p6eYx+IWToyfJ4R5p7OH2wxk0nSdQdYJ9d9JE5UTH
EuuC/0utbrci0ItCa4BV345o+VoMVSylyRaSgi1v5Dikuc0WVmHu854NFH2bs7Fo
yhyrFV94nXrDlaDk6M6/omY4F2nTJjnO4lSsWS79MQjSowv1FPUPLPmkQ0HeHWoE
beef55GSSP32PmjLVN/JuPqh43sm/HcglcckghX8YFEwUfWaTeW2hIQ5szKCWhfo
vMM4Sw0MoKkWCHJpw9TmdvxjKfF67Bv3Vij6sbLdj/E/xJR4HvfKEkMtHrHil4ic
jHlFObXh/aHU0CED4uB7noIQjvEbEr1fIkvtWfOSKBgeBGiuARTHE3BxXe3t71Fo
4Wk7/op3s2X7JlhuB7Db5dvzFQaSytFKzftz4PIu0I44xJLcujaPVlJ0stbw6voj
BAARQhqT+q9cjxeMG/pVIAXZnYYHrKyg/qQbZH5TVEgojeJ8+C/CZkW2gBvsCLVr
6/bknxleYjtEqr1N5RXBp6/aPoGeOu1y7sLI8nh7q4S0VpwJI3msWW299efdzhSX
dNvxVobmr2mGwiCq+zeJlfZpCxwO7w5ExnJi6jHFrvTu/4YDblDpRyltaJgQ3j8U
3i7Q5hLZyxt57XoY8YBoXM8Ffq065CJiQqXpODIExd/RphdFWvI42EtEaeEXKgEU
cwO0CMWtOfEt5BQSIJvY04IUmNfLQWaMQMukzjM+KQsA4HMOmRs9eA0yVIxF9E89
8hOaWMG7cL4h21GogSN1pH8k/dPxZlLWzvblSoyVuD89x7VBARg9G4TmYhp2TRZH
q6WF261fZBysbK77FfzXg/BGlnH87dIl18jOj2WcWoTLT+k8cUNgv+xBw8meviEN
zHtR2xv84++MBtKOzvIa2APT3pitml2XA1NH6bQ3znylkqN8T856epBBQwWpus7f
NqwseTQCbJv5UHQVH0gW+UYBYRgxe/4VO7v74O1956sl2o7aJP3QXEM7XgHrCElf
gisF8iuuODp4eyy9gsCSlgBB8kIqHrITf4IxfYIVeIBpNL+M/NKhkeQAbTYCnGUp
kl9zpIf9mYZDM3eGcVbNn6dntBQ6nq734NobMTC6tp3sdKl30+fuhlwkM9YegECu
Pm4ljcHUflxkCcUBO7ikvqvasWckvtFJR/YLu1glUIRUSL8O73delOhfU+IIdo6H
ERAXNGy44Gc0fr2jjAoQxbLLF6HhtcOh0L3BC2NrmraPuhARoB5FiieDULjIoLNp
cnOa3blMGYgErCuMU1dX1UvDIt71PwK40DLstC349qVDSTiH/9sDK8ibv/HhtGZi
+vvvBZARPIdJEMlivgvCT8XNq6kANYvJAAoJGUbfbCFQ6bdltkjeDyTPMrXIR06Z
HlGwFTldQQ5f2gTUM9W2jrh6dk6Nz/NwFsQF6uGkiao64IsqAbJ7Jdcar/lhoYVe
I88MHrC+/0uPpYGXOZkudDmPHziGClGW5MAcxvb+2AAD+PuWSdmYRzFX8o3usPVj
NWn+Yv3vxo07TxyX5cVuzzbWLapS6iKVN9l5xtLtvNFoZrhjJoJ4R4ZYd8BDXr7W
KtZiLmZWdtiiFJmqiMgemueteT+JatIi/D6Rsg+4rk9slsde4zMtVMZQfCw+3t6e
DX4d29tZSRJV0cOpvznfDIZ4fhMXVca3G+0gJtq/Jl2Pqd47nMetmTYO91tViA5Q
E4ARITDHa+LvEtqgwTWh2RzoLGuRnZUKBKeMMLmtXqby+3BcuJ5H/nHnx0IxYnab
/wYqLF5U8ZjwxbWYpPIVvBsfxd3owJ579UY8dZZQ1+TkRhT03lZbbhO2AOhlAhWV
ACtFbloZv3FzmpH1Wr3naeNwsFo/xD7/WUL8wdM0tpalOhuV7drCdzlLRp9QsYLf
Jx9pVw7jeB9SHwY37qZPx7q8d/DGL0Thvb380GBWnu5rkV5bHpT0Eapf6oeH7VbK
uVWDfrMWucpiPwsQWIbHTD3TGjf5kiWexIGrlfdjwjEuDMZL+NJ7R+mxkCQ74iqk
d2C0T9Ge2gdreVmYINjG7bPywdzsRiO/cSRCDSFDzXZ5P4NYVpAI4bPC8slR5euh
/ie5NiRxaywf/VoyGnAJ9NRxa54C4smFBxsfqrFkAJLMM3zwGG89dTUWjiqh6lpb
W+qa4C9Ed1hME5kRrSb/C52rG5eOanmKUfdPvN470T0tomK9UdN7Z0Q7IFer6VK5
tmW3aziyGtDpyMJ1aZrlVkE+rOH/tOteHo/3nfV2dCv4BmydktHOXQ9qqb7rxltf
Ul7Da55nOLBPOqQcA1kCMOwlowj1q/y1WdQpHSU2XAbr+QLLdOnhTw4AY/+YO3l9
tk2zE9gq9Hvzc3IQ4hQrlFbLz2oMTDYig71q1GttFFonBXwCzR+VArAdchN6sN1y
4zXwqhmUyNdZHcqI+92roFhbRmwLS09hNsLUu1owcfQngNzu6HzbMWW+tYeoPsXF
AImpaBOngpQbgTPhumKwNXzJMgRVaDAUAJjbwhmtrJGBF3eOPwqZXLaEC92xkENC
/CJlbanOve8wUUOaxR1/U3qJCwDSAuGBNDeTqzqOEmu6GCiR8P2BQpLZBAoEcZ6Q
+pMdw9VyHKzjlZ1FtKCtDgN2JTOeHcHIyoBWRwGZXlVcdL1b7LDnHwbmMKENeln6
EVxV8d0ZajstYo7kZRjNBLXH95QWcTp5i4TeO3rmSc+Cdd8pbfJDiNBmwlbQpS+a
o3lrdYxbRi1I0YwOUW5cRU0L4PmTSW1mYMaCndGRqHKoxi8jsQqVdqEVShIG43dm
13E+c+85lSfvQhU5MdYO78nMXFigR5oubDj8jWnxl0qA87Z6WgG6i5Zh4I63yMN9
caBx3fTJyJtZ6LJ8quRPASOQPbVFVukbNzUA4llaz3b9Q3cyr/+oXF1a7pe75LAX
GppZGO5dDGf/SqJV0CtpicTjK0AyGjYuuDJkxEEqkenRwfBftfbxPXwSy9WZa1Vr
xmcznBiyt34KYm7syHQY+TUOZ17gpE/la2UPwhsPz/KsXe3X636DTyOOydv0VC53
ElOeiVom+agz1nnQCqVeXjG5nl39Wioq0IoQBv/rrgNRFmZYQ37xos24dNhHJ3zy
TvL2Xq7dNIdsBphVE6qphtVBDcwit6VjurUO12oO9DwGT+JJEnNhlUYpeKf+Z20X
5HColvK+yKmB5FUxKgOD8PrFr9vaKlLvqvgexHHTraYvy/QNCsFzgvF4zBLFUMAo
L7L1fwWzPiFBUzT8dn11b5PhVlTTrnHJvw4mcc+J4nqwo3sTZ/gvPww3dSzxgqXl
SiPYaYoAG/ct9s2xMGlHe8PJUn988tX6kChuJiv8Vbt1tKJ48a9A397KM5hyc2zf
8AMp5U724yVivOf5TNOTkSyuqkLcgJBTHyx33NSHhS6JMLrJD9DxNhAtF0vH+5L+
G8cZ61+robfScCIyVsmCwwZwMV4R86Qt6/tOKgXopROzpqIeyMMYLmvN1vYDIxiG
xDwOJ31fb8+ba+mnK/IpQmacFFnP81fmEeP1kUfvMAe+nC7dM25DC+Ey1rKjJ/Fj
pQ15hioGux77dlZGlSyG298eTomIr6MnVOLxwBsHBM65RJgDBOM+W/1c7NcnlQfG
3vz43vqjIAxd7f1f4vG9r4H8GgB+e5Q7cakDsph2CVhvvh6b7VSu1MdsiInDZDPD
VA7wKecgD2ztrmguBAcz3hUxIjo+TebhHBeLxxHewDsT9B2wzEhBWJBmfYEXmq6B
E7UCqY5vVC3Uv4aEtf6WEX2DLITmPo9ZWsSoPvhSqq7UBfc0S66uFKPXG5quv5I8
NZ+r/be2301a/PC5Xtm1Hq7WctD6DaeC69bgldxWpeInhGh96DxIPOkaJSzvE/Ry
vWzZK5kx5vSp+qpUfER6TUgiTkBFQwfU2VxanZy0t1kP+kN3mXFMnsvEn6rtIHDa
tiyd2bfQflIv5y7YxOAKB09A2AHHwO9yHBD4+6pai0qMVieZEZ565VIVQEpGyOAF
PMi5SHYYspgUr0zwiY4hmFT0B8SrBPpFTGTGGlUpIv3ccOP8P43ndqp4m0IPoGrO
XbwBa23Iqfsug4sTpitEKB+DtgeYe/kzjyME1/OhH49Hwdlewox0bPTp8RH1AaRI
V8mGsC1wFgtb7KD50uYBvFuo7FJpJhONqtx6spYLU3C6dkTYOZrs7YMBViGj9sWM
IDjp4HuQpj+Bh6x6ClZfzr0xoeRzXNIUG3MC78GyWqBzHGcqIxgY4weQmbEc/81H
qMlY1/i8WqK+ihD5X9+yzbu9x5urTTK9RH3Q4nzZ9kIVMOAkKAOC2dYwkx3ewIl4
ve3GQKQh4Jexcc/zK8nZtyvlYkAya2SUCNUegryE5fMeo6UCrQyy2SUIdRl/w0Uu
BWMPfszOUP+zofEenDDNSsJKlaJ3lUiPfaUJn4ShvYGExVQr1UFLfelMfxrv3WHg
pgPBjXvjWwjtrnEmf0t71K1/XUJlhsvfwFcsk0d7kHFD2QWxsGSx16qOPM+0QTVM
7YgOsyR6dTyGHkM39UPbe8CBMQrwanWrid+JDTL/7PlZAwENrmP7jIlzQlpx4NRn
iOuERQgjqQ8gWXG/qXv5QmV4Xz/tlDYcdkf2XDqy29tGm49jNRBgDtZ2DFOnJ/PD
O2cw2dmze8oO/C1M4T0TzME6NEh4xkEuwwWp5rWGVXETY2b8psvqG4njJcKcX63T
0C5Sfpdlf/y9ALie0vQbMnUbd/YGXj7taYO/BXPV8XDG8GJ9uDwcz2Y9+y3dhTDd
kQxaRmvj1uUTFA6SWTisu9YzYJHJ5q5hHU1OSd/FC7k8rjGO2KUW62Op4IzivaHm
NbCXnfXE677Co8DZeIbo5eHnZ7/pICdgEetvf0I0kQh0+nWA1Ycw7zb/qWiU/Iu2
GbyupY+bLgvMkH6q+bWI17QxtAI/pLWCUY1oic2fMlFE0frETo3KgzfxJHbeXUXD
TOc3jdYIIJXqs3eJmh+lx1TiKTynO8ykVQtZYRMfIxZGYqhZhCUXNlikPmdvHTuK
eAbCcu0cE9PG4EPCGS/6KZtPA8/Z+qTwt4MHd/DkJyLf9USv8sphhciWSQaSEs3K
P7DEnNAfus4faI9VIMCLMLMz2UsFTU7vSp+QJlVym6OXBzejX0Ux2mu5iKLVozzJ
Fbm701tp8zOAuVus+xUzJ1M1WFRk2iNQ8XrcvW0ZRcFHMmD30E8/V3JyPvXGqsJK
ILFn6VQyzPtoDDM4l9hJHlQw62NivnKE2+3Ia4axQ55vZ222h4mMwml6hvmw4ruW
oCykYMt48sQADS0gBvWyTsyoFDnrO2JXKcf2EBHowEqJXnfEsR2s017cEZ4MdU3R
iKqBHzLHCSLJrya5B6vdyNFhnTDQ7jZ93TfJLGVkC/GZyZyqWepXS3612ItAuZz2
SYbghFcDgd0QjxKIpOToE18POMJebeX3kVycKo7ssU5T96nQjvSgYXbpcYxBYM4o
RPTw9EBY7PyUKqkqBivWZNIdrFFelIwgClzYj5qeDlqyNVcYQjJdqxF89yg9YLkG
8ODDLvXv+aME5pgmU59oVE5QhGYnQqwHpkxSxwPQIY1NCp7MVphuE+GRlfSKjyY8
a/mxcGtgzP/UpeCs5Pe3y5DQDSeXrg+uLmtEGQUGYfQasdPXbTlXv/eVxy8hHcQj
hOuq4lGSQZJWxpmUQwK1JI1pMpptZVOm/nd+2qIMCUTGb/xJbyHkT+p9jKMZA42q
6YkzlIFwvODC3PLGcBBLG5i7N/5ZFspU1DC3TA4cI//OJuaDj6X/AGUiT8XzKk4T
iQ6xBizPoAb4G0jn8K7JxP8cQT+1G7r8+wLjWd0PgE8CKUXnQxTjvQ8PQM8/b0uT
urHHQI2/j19jWP8gj9LkspyO2q9nNrf073IUh8chbIwUJaKvjd2xZ5RhIfI4SaUv
bHO7okxvbs5M+MC5gel99NOlrmfgMzKUAAn9WMMrermZUg/lSb8NYb0vTDqbBqyo
0gTCdERD8R+P9iE9Puk5jhd4Wp1fWWUJS17kgofTTbZlJPY/Zaf7hR4a+p/TrDr+
PYup6iUr4vqSzEW18hGVo7KAYNDGJxbbPlTqZIhtXBg/mdlCZnb9T+q9rCwqW+FT
jnKKxAB7oqro7yPq0Q3ni9cYZgm3ovrZ1yhEJPuE4tK2jaw7JHPcYzLuR8iFTtIn
pCt2Kc0ddeZEyg/F4UKjjJ6eq8go/4LanC+XN6BmkE+eGX/LgMgfQEe6utl6+OpA
jPtTQxY4EAfwBAvGztGKmOCFtE7hQ5ES5Vm4TFlabOpXlgH0qYISZxNRloHV0K8T
LFCTtc1VXH5Imt2O7CtmUi6WR4GGgFOI0p/EI29Jvx/72vzmj1pLo7QtTseqCP/M
zCP5dAddBDv5dHPnXrCg0cm2N73n/PRTRuzKm9Ql7IemJLqIy1l2x8Kkagd3sHm1
GFoRN+bCmBjMjaIvJkkIowTo3NNBBDMm1XJOC7EMtrCtFMQ3/IAm9wUaly3fgDUj
/lhJ3yFhzp4a5xLG1GyI2AvfG4CoLG8JdO8Wk6FGWrrxpLkxPcR3aczFIWjyp2f4
ReIJwftiRV5ctcb92mXDSw1pDwFICl32+xLdE8Bmhi5FW4GnTRBVG0kK3baK1Ctd
u6JRoMuX5hDHdxsQwsTkn5sAZ6Q9UEeqfiV7tR77miyb98Ko+FaJNcItkUvS2aOY
uGDcFFRrTI931hZXrWk8tLniQn4tBimQtR1LuIRS8Ms3qZoIXDZuuuXbBgSBqy/2
3HFkphUDvreJnOsqCKPnjQV3ZvU4auDrPeRGUR3Hs4KUonEfoXon3LzNcXXRtmNX
0of+jJFMZUlBEHamI5pF155bJuLx6J7NCveeOQsa8kwAV7Tsogqr6GW1Nw89i61A
QscUZ+SSa6KtrPMFO0PZ3LDvByDG7dcIjC+idkGuMnQnuD1E7yV8DjdW/bZzULjh
j1VeRp7Xjgxkzutl1IfqiAZdTV21xdVf4zLEHGAT/vUYmU7BlYkIixA5wCvpaWwh
GuWV/jRpBciDQ///T7oyx6n5sjHYwwIupkfivRCsiTtMqq7WsWU4/bIr0dJgZhI9
EhnIRwgBPWHK8Bjlx4Y4xhxFYSxkECEOJIirCCOkRTGXXqgkGQNIubXWc4WWbwhK
mdtkMTn9qmPUErbtlu0qqvlkn5CdOR7hMhIkMfsTks3p2vhJgQUoOkM4EFhzXRR+
9HiylQYlmBXqxR0eOBw+iEZp8NJZno8MK6fKlcLWS5Xj3lgRF1o8fbggETEZJj9s
0NZB21Y/GPnTuXAd6HZs7RYQ/IUeuFyf14nQbY9uSEUIf2rjPvwWdEL9ujq86hKr
hEYRRgU1jIqNvcENJ5e2eGB1OpE341J3yolgIa2Fc47pvM6cQggBDy5Ydjckfja+
XNvg35+VWyxOFe1bjPed0vyrlpZxXzloKkdetss0N1awCnLT3YhEZxjo3ocwwovs
05qRZoiu9otsgXcjvCBAKhG3Kgbl/tL93Q5+XsU30Rz7Bbmomy0Yxf9xqc5tSN8s
mB3vEVGb5nHOB+nRxCbAzF7xbZaTTqjD5Z7UX1Uvp+pgbuorkUyiWGoQ2rG9YgaX
ulyD7aDZ9vkst5TkTsNqO2Pyb2wUkK0+WRpV08CxNpqCtzNZPxhiPKw423j7k+yl
zzQfX3hec6fAgQiDls/oqzdsFZObF6/jUmqKqsYDno0yiatpPwMk9ZTkoUnVjtgU
iVBMYdqhu5SwpZuIMvxL8e+qRs/vAj+oWSrYzM4SnirWCNNy713rZVHEQH+jNdAZ
FAlteHBXMft/F2aTh5lLtt/3f7UR50dHm1UdlgP5SfaXPvygjAbcFPBN+1Wz6/rx
tXIWNFns9w4iXmXHaaP6DFbG4tOWZkD2r9ylvmYmqV83he3xdb/UHCdyBsMnSM+K
DZJZc/8asNHQtliIgsW6tKBFg02+iR7LAd1kT6OVVAj+DRomrEOB3XsC1LEzWgkt
w7vhjJZihaZYMVMpH6kvvfjSz/8SdT7szR/f1JLQiz4aTlY7qmVmsjoJDt5b/rCG
mCSXWXNbFCLU6qC//NmiMv4XDzxU1tOunKO+ZI4qXrcSHu/BtQyQHVha+eOVRSub
OO62gKDISKJ4/HmJWU28s2xtGCJa6iQcSJaVEh29qI1xL54WAqXgGkEk2T2UMpmW
PmouJsRlUExfcXcwYPp6LI/DIqvgFUFqFshhDouS9mqQleKp8nJnLuYuN/Isqn/B
k0D/oenAFQkoyyt5fO8FkSMt/kxZGbMiwSyHmn3dKOfGBpXrVdG6VlLp7w4Dlq+g
CGyoUjsr39aEEETJXdNLgnaOWqCdThw/zg7BpX/iGdrIiWOicw4IuTDSQnHsKx+h
6mqVMH62kgClPobNP36c/WpZ1tjTeSWtDAXToXG9PyWIaIgyih8EpWLIWb04PsBh
Xp22eVLJsvbHGSKWj5AGZjFI087FkWRNzbxk5wc4XmGWJXOI8E4klgHif9zobKBe
513D95ySgGKp66xz/8HZCJmMYi9yZEa1Kzja9dWBCisJI3BNzn032PzJ1H7FFe3z
pfeQy+MpYNR/VWSwQvxG06ePVG8aBh54doxMqZKw5wHOv2z6bCpe4Z9uXrKUDp5m
vuZmURKob1YMI0ZA2rO2OJGR++kkA2Gt3DIqjZxNy8iiPXIXRQSBTd8jSnwrYTJc
GPLHVu7POTNdGuIdzqeFn7QsgA0UTrYU2ImI+xSu6eSo3VLyYZuys6z2ZLFmNm1z
38x4rpwGdeHOLATO5MyHY5jY+6oiO47Dw8OCFpEX33NAli2xAyyIO8D58fLSsRfO
NoX+QJjluJTvLBIwENv/f6ZXU/Nx1of/As+LXzpZZxOcfMxNyhWgZrdu5VMs4hmj
cPJpboOcGbiifPPlcElih+sYwS3nGD9OaygylfvFOQizCq9kOJVb9N1Uo1p4sqK3
a/ZNWk3xnvuIKoMaV7NQ0bxKfrCnFTZxDUkLbOgq9XweqAnrvAtwfAQ+75M+m0R3
Q/8IVd/I8bxFMm3DcwBxirtqK9MCeXDDeveTk8vIaiCXqJANYKM8jblR74uxiW6a
hE/RHI6434e3VbnZuMngV+H+ycMjUQngRpr4Zl5K7VadcRtKgr4wqYbG3vvwlIUM
iMCe5pxnbWWYSD+wUWt+x6Hh+wDsjysb2xAR/Ot4EJdjVWt+xLcg5nbq+H2di8su
3RGcGurjX4O76iCC6DhQ92Mp50As6nx8/r0t5Vm01ptIengdr4FotatuoL7aHStR
pqIlV+i9Dd0VaYn4Ay+ctTIlEPMdpmvYmE+l7O9LHfSYi2/EVpvFRzIzf4bS4sCJ
nPkMoHrkflgVmRMAnTdv542H9ZgoOVCZT8kr2On2Bl0PCtINxl7X44HX7ubZH6v7
jhU7QhBczFEYJHdMIf8/q9vSxS5sAozFbQ4Nj+MJdD3w7D3hT/qSkPxlYrHCXWY5
4uy4LuX5E85jpaeluBahGPrMcv+E36NreSohu9uZt1nH3RuCK4biXs69uPM+swM1
3Lnyp2ypf7oINMTYTCkEyih/CmZwwioywQqhYJzOMX4JPa/pKUpRcbt7LN0kjFEB
Lu9s7PmpavF1MYb+aoDLSjUEvlNaGBwJL7x/BMc2Rx2lBEKIzpOqMgWf2pDsauzC
4nlVb05fg/7h9ssIunpY1ycikrNUBaxB2SCYoQKbINLKDCIvURmutUmgkjgUwhEm
Xl1SRHl4HRIB+uTnoeNom3UyqEYlS5kb5zstPOp1r103w5KJjISXLo4M/vjzKL2Y
rIWvFGU3WnSDskKxbNdljNV2nLzYz0/E8HsR8aLSapJYJyORxpVwDx2g7N2kzs8i
qdaYxba+YUyljHF7uSELLQotWMTYGKt4ggZUBgqhZiWliDjyMdlktYtrMv7wrvm+
ABk/fvDIz1/k058F0jPvCZeE+pY6sycMWnSr5PtrxU7OB2v11vvemF+jSMD5ZUZ+
JwEv6vxQSD7YNLFK0ZnSMpMwRqi62hpjokWApc6SzVqvV6U5dkt8QnTY0bPVH/ca
VV0RfQD+7cPV5w6OkyrBKgKs9oIXyBHEuclhO/l8+CHZQq3qNtOtnAirEH7ElI2m
WiQ6GO9tnWICFJagAfuNVTdn00fnueV2MUwoLuIle79QgI5Vh2dMtEvlVLZ8+TfK
pGgbliVa0eoD1gDDvhp9aB/if4yr7bINeO9eXzZP+YVVJkIMmygDDIOHkIzUOPSK
2CDzaG+ufdsXVf9AMnUA7i+FdNA4YjJQO089BZ2cvTUL5nmhES46Ner6xa1BfAus
eqNYP5LLXvV8QUNU7yhTwYiDyKLfboG4z6+dKHrwQlomhrBxCy2kMnngV7c6D/OR
LBOX58Jxhs0g7vg+qX0oIysnCjhk6aSSmZ8P0YjCwBUzt//2zVmPojymlyYllVFI
awyvHYoLznEteYOyWXtmuXIS8SXX1xg4E7aMFdBMT/jQLOsF7FO2oqiOsJbR64Ej
jPJtUnVLehYzaNDEQn6ZHlwctKHn4m18IfTItG1bgK9Yg+Umve0iP0A+orrhqf0k
Pm6U+kbJvTd2Y3Pwlo29v3Fe5WCI+TEgYbp/NQtt0zGUDdRVwi3+uOFQCd/nKSfy
CNBidPa8onRCcQTSHGhVu6KFFbY7qAA12c0W09nZiMsA2maWIg7MdPNwzlm2hG8D
T+GP8RHSKvUSyxOIdHtfS8eqBmZo46z60cuhs3QU5B5G9NtzsSa+Bw6TH3Pd4OiO
/cFHu8O1/prK8ldxwrNVc7HumcfR3+LLDFJGmkKGbAsMstaRnmfJXoLLW8dLyFrV
GDS3zwRZw+3bTs0d9ueTOzRr8YR5pg4VSFwMeYbOZLT9JHrbets7UjNm9lLopZI5
JtUmTVsWvrVvxD/mPJmeCpUIm6cQbT/rKBsVfW8tI8p4/gwatnbQNqLiNDIAI/GA
BNVC3XuJ24DIxv0odYyjCjrg2Vvt/JsSkKcAXL7RYcyfx3s2OuKl9bY9UUh+ImGC
dE8AsiY9LW/h2+m/AJYNYVkx8Cqn72DVJPdFfYgG1r0tgIkzg9PhtctBdhrlU6/E
/AK/aza0MbxPykxYaEauDEgtUZQBoK5DuL8efhaVgSeUMTKce9CYFPMJLh6JH2l3
wT85sNDdnmrtpPdR9BPzmvLiEnftcIMVW9w67DLeMexPJb6N/rpSvvVxuc6drbCb
nTtNrrcz79YAkv/xKJA8wvCVZoDKnX7mBO5jO4//ZvuabsOo84LJBc41juOiKIbP
ZFtRZ5W2MJd/TBvQPBVi75h+95v8pkcRhD7q9enH40jVdPTagpFyzlagScOAHNjs
82YwdqywjhHs9KzbAOPh1mJcdYOmAKTzsGQF/hZ8pJHxxAr2eq8E5AnJJHfeiLXu
5WstkioP4u9UIChicQxRstCSisGUSNRQKwm2mvONyOqKMoSWpLiVjMYRals/u1ZV
oAiuboGIWOdN5d0uR9XpxanCA3mJlIx1LEDzY+zP1C5lNrIHxrAWzSqtDQQt3+em
olabDlXbOP1K6NA9jWVQu/RIIZOx6a7ofC5BIbQknT43cPiW191htIk9OxeRgVjO
lWG5fjT6Z8DlWzGQaB5maM6ny2EoAideEPyOHguFgEIujStuGSlzaUfLUOrJsDgR
3+FjrhjL1WyMn4rr8/0KKjalrVM8IIshfTjvkEruaRD0J7mitTJtOO6cBMOZFIph
rvo/TLozgxILMAkVT6G6LY6sk6y1qtL5L592G5RmuZTSzJXSKWkuGBKsZ7o4bgFf
GcaGaTz3ih5n8eaTXCSLW1LteWGxi6g8P+ugAl7DFnhz2IaparZS+vKxWUzXxuO7
h5lLfSvgYQKguvqA96Q6zkIh33oBi+5TQx2xdXRMQmN4Xg6fFzSws/ByzDHZCudY
pP8Ig9/aCcU3a1bJsxAJz5mc1C39YbXdRNbUG8oOW0DrmzGP/v2ezw5SxCFLnE1Y
QhO4YTYS3CnksjPB1A4SaZW1RlBf3fGl702LUCud6wC0x+f6kyk5eBAVk+RyHbfP
B1xeosIKa3pmZIvjW+KE9CyuCtE+9iLJHy5d5zA/hiVuSLI7FLKdwJzF5Ec3bPmu
k6QrDAwSX0nKuGEx0IqPAjNK+4Y+gDYt96WRegYGp9kwwFdJkqDuTuQoy2HxVEJM
3tt0an247wrDwDSdJdfSqMxRhyIS78oz2AJH9rHOmXd3hi64wMep7SMVDJSY/LJ0
xBPRTOrBlYBQyu0iPzdZHtFY5TxTv65rqysgx0qoTef8hm/2d9/gv/8gbkQWQP0Q
5qM8sV5LUq+67PfiBnBsqDW/jz7gw3ZRe+kOCm79hQ3H3PYd2ywU9jZElzN/4iHj
PdMLX+CBa7unp/3Wyg/EPfPTlduXGQpaS17qV2iCiIZ1N76/k+zWsy76NziRibo6
74zdGZI8qPbF21Kwn5NGEyUCQ3R6blLMj79md1hcA+8F6F1+3P35UXkx7JY+UbA8
F4XP8BwItTC7xxlPPj4d60b68Td51plFhbWqtivNDtaZsd2q2EVprHWyj7KE60nm
15Hiym5eleYYH7Vjw2hKqKhHxjTVex7a5d3Qilzp7sSNqMGp5XMd8x9LNVp+wmhk
L9XaOHKH3Wr4ts+8EBYcYhW2MwxSa6r8UJ0puqD53GVLaUMhcwbeTT/PE+Verln7
MafBMnTUjisrUnwQHqIbJy97hxCHdeG+8bDvsJf0jtcP4ZQ7UbrCvlF1/D7fh6Li
P3jAW9isM4KRzLJIjK2lWiRvBp3jYO3zPkjq9lVnQ4f4t96CZqQmrzIIPZGwT7qm
D9vxGiKvs5Uomht6m04ghpHbfbKz3VIegmv8qO5R6tgTbpONidBJfjm3eJazOgc0
cWwnAFrFHZQQS1ahTCRFEgQyk8ng1Yzwc6RH+UgZPKX3tURZJRG55AM4E0cOHF6Q
E3v1AYg1ECoPbIWzngQFjtd9JRaGEQuI2og8Fexgtihq+4ZZIGYImjtoM0UcmFlj
Rku3Y2R5SXdyZQCrBTUaQyhFECRmuFM3vKl4yNFMYYlGRY3QdI0Bq3SB1sFE1LFP
2IbtgRvqx+qgCIM+h5lR/2Px2r7paUkMMhhzshHgyJPnbC6MwGMamzgAzaBCalyx
iyDMl5OgJcogRRQXmxD1z0BbWaPf1qN9sn2aIgHq4XfKY3XgJ0+x6ZIgchFpPjOU
7Bcy5qi2zERjbW3zE8z6AhXM/peDCn+D4TNUx+JFiUydQTZBMkCEFWT3wfXlo1HX
HW2f7WvQ0qhm/MeTwiiDwZuicWYmc5ABiEQUbpo9mvYZE20KZQYXN+slWk+VjAz9
N2aoboYspfUcd30fMJLBBVXhX2i0k34g3LWUtjDG21AYecDEYwZouCAWxE1cOWB3
+BeK4O8k/sL8acVnfd5YLiqx1/W7Pe67ctoUkuJIv9UtIN6On7I1OiRaWSYtvy0R
tyqHIwg1FkJpZcqNSFbvpyQrg1JZ29ZsaGuAh/ojF0h2y73VgFD1hiIIqP5yIHD+
6kd8G4MdkfLMLZ50z8554ayRiUqWj5keo5PNM6B0e8XhmVRtL7BQK0KPjSymUJdm
BBue8MrZ7FldV0xKhzgHMHkF2zCWrt3yJlcnT5Y9xWOZ2T9JKtcZotYCivLzCCBK
1+GuyPvNAYXv/d5Uj2iClMElXvo3IIL82/dBZKHvwhR6y7zx1x1eBJqQWE2KtWtN
uGUy02qjODtG9pFdEaK0XfmlNwhN/nck1dqlu9sZ1TG0ngCWExQ9gc+hFspMlNUq
0mug7hBRc4a5RGWBktVkqzsIfOZSBwQY8d0YK+KW9tGhk7OhZb3Ip7OcxwWdsz6Q
UgyjgeQuvWtDzr48UogSQMLlB3Ng9mGA27t2HxRAVyOQz4CXHly8bOPm1ET5SQc4
cVDTJrFDShR9QbgtaPSezK7VKfsGxdb4ZdakiXEtQVyIUgaa9PSEBkBF10AMo11y
HxxdLpFfOSlpM4zZ7yYopmYuBgg7FmyNvn2+nlSef6Cz27Pdv4UcF9k72VHLhq95
7gigxCm0xDJSPi2i8g5hh0B7mbucE5E4buKXE0FKOmNCrWMV7dUL3do3+lzA6t5i
mfbosZbahvaGnSrR6Jj2ziD2dbWLK9IDto+YBw6dV9Inlc29oAbwve8cj2hKm8pS
MnrkfvNJrrQflWQxq1emGkhWYZHFIZlFDLhqNt/+d0YZbTpytAarmfuwO1yt6PuB
ec5hrEnDhoKu+DmhMr5yX9wgSxJ+EBIH9x/M+W3OE6AwAn6qs8qgdDqWarVeTGeN
0S5LsT6tqF5bNC6lkdyiOv9iJVGP9XKUrjafF0ALGWVhmT14GUuiNqkhTo0h10Fr
/rXBcdgE97CkfYE8bt3YPexxwSDQyxg9i2W5mzvWaFMEmBbCtk8IoCP4og8sw2Aj
V1KsyKh6qP9A3ODOIGmTvPI/7anfWtyonnqwrUhOWcHwi88mNB5i8cbZeSHP/V+J
I71wu2sKgC+7wlGjGyaP9q2DncxOodwgaXqhSBmeW5YOkd64qUC0QpLvBXeNFQ+o
hIN+vSvUMRoHLGVpOIrXU+jtrIBhWkvVpZ5R5S9eQsVeEbhLbFfVjC9XtQarxz8Z
x5ofL5DLQ4e7TiUydCWM52ARLWzkWzZL2WU2evBE8KNFEHTv8UI9JcJN5h5gxixu
V8FfbfDd6VtchFBicN6Y6ISCe6UcTjXrkLeyuBmdNmG4TJmSv1OGB/t89Uf7OQiQ
oR1TWpuzH2TGp3/HS62h6pZxzEUSMd3t9Yph538rDkY6H+K2gARUk/XkllFimEDa
LL0TXcKo2KiKBGDsbidjV1J4dBT7Sm5m95wCFxsphVzGI7a9I6MSTuDBqH+qVgXK
8pQBx43ee9IB4SBGeV6zOfog/qY5JXcLmT3D0gn06dmFLSA8loETPRI0nrO99+FF
5xNV671Dbh/ZQAHd3VZKjXnw/Uutpm+BvV/PQ9Cj7wEe+zfnocEUfDPenxTUieyf
fSISjIZ4xJPB+fGzFK++pTg6OGP9fUCZKD8syo2SRGBSH4BeX4ks2zfz+UI20aSc
vhKOYfpa5YtWec1CFcKkdvooCUQn6HG8G+lWu2N8NaD7cM8ZClwWEwoOh6IRXx72
/KNFurJtjpomQuzDDp+F6DxK4kEkxVpaXFJiBtudOWA0eyBbB15jlSoCWastxS0W
aF3Tw5XJQ6/uzpwfYJ3Gt1hamo0uu9+is4ByAys80XlwympYyxLphuVy/nFHgCo2
ZIsa5H52ryZhUjYrcsmWDOeuBfjwF+6Ivcxi2PEeUMTYFVeT6j+StNGpGMDOR/Q+
FogUBGgRQfKR9n0ZnbOyoCc1L4czVxJgdE3yp8cZNpplnmR8VNPaADqdHvopAuz/
JySunHXASI9oZ9A3yS5maUsBB7i4QnYbpipcmW1YA5TK3ccJ8yqMvS0lZ4B2kAS6
/l/QiWfH5/tlfYENCWixAxIziNuCIS/D6SOJyhggPXIeNEWDbri+YDeCFIl9/w65
p4UkQE4TLQE3SxdMgNHCTkRxdI1Y0FyXmspyhJ++8n20LiqUKX9CBaYwQvj19SBb
6fiHlPCyM7V+YEZMWfNesjIzghZfiWZbS/s9gtyQA8bb9YS55eoJqdDYrDUQAvux
bvKedOOFwcvMbv80AFo7jN2+jN+nMQwhn5wqtzIz9Nq4FPtIkSZ9tuirT/Mtu2Q+
wIUs1wwJQ050gkjHCuJgUmk3lLzs4vsLOfcQX5OtFuMezN17TyXy9jwjGHzFwdZr
LnWpm7o+HT2D+Yj86RXjv9kevTaSRhXFJFBxuMESWyexwx/fdLOtLpPCfid6aNp8
BmimTViyWMVTxmozDCgJbJXrBCmNSwbrQvNnthZxEBwUYR8uB66ueEufD+VrCh6v
/KZmTLWRNcil8nqj+faZ1BBCc6duJHiqhRqpLIxilJfOkYJ39gZZbO3UIeabsm+V
D2hQPnyxjidNOd+Qt9Y57S5+3DNukIlFON+PCTeUicodIOl9zRXVJYxLNMxe2beK
UbmugqG8pDCktfAxCirwSuvHuW7PjpvLLBzyFz6JqboIwtYJThhNJbzZFq4taYBg
78o4FezibKVsdYA8G1BJsjZVu4hx/f/K4DCSJFnZBluL71u3p1i/cKtg0vb85E1D
l9n6skkUWqc6MCvf7L5gKgxN6wG1++xcBuVSOTY9iOk0cwNlZvTHlGsLNlhY6qA3
MwZihH8OE2CiDQmelJZMDq2GiSdJK6Xx2v8i8e3bUBu9T3PsmdyyEqvIkuYzm6oN
K+wHMgvtr6sXBBf9G/y/PL1ue93XeHPeSC4BUcsbv6Bi88k0NgaxkcqNuDIQmJYJ
fPDa4xtIa00QlfhFguOAyVs/U2szCvWIiv+tFjbIQYGMF9tJjiPsGG9mD/+zvO/K
E2kSratTlR34lByixTvAv2s8GnbkOmjlb24GVOGRAnIC6wA8Z5VpZ2s/Yc+TgUmz
csG7/jvNV7dArCoSeaPqsAmbf3jO6fftnnCrpprdaj826wgoF/7KEHSUnR6Nvl0r
1KJLHtVkHLqN5dKdJfx50EZkuhju7HOmZD1EHLXeU6yqRAuMRpJiPiAmK+BxiFI6
a6XZwmcOGyrOmgEAsSFxABTrqBYT5qwT7WtPz2duHcE3lt5oBxpiz7+x6r05Xl/G
YiyHzp2VGj36IDR/830ufKTc2Hasmtb71eb6RBlVdiIvnLclbZpsEhZGE04vr4Uu
+j0gwLR7wwkzcuaNO5iI+lqk3el4jMHqbzj2EiLzfDIUcT78hJ099iQFSOtVMifJ
wAESyfXzKKYMmmMDN1pcC375lYJJAyTrpRY/OoWNcR1NDtdsDkVKybbGqiKPd7ba
d8cJUZigBxft3y9MbyVAQ9+x5LdTcdAAc3hkpag2L7BH+yqyCxPW1VR6hprsxRJM
15PxN45b2DO6ZS4vJliFFfWvs/Pyg5bE2+tAQ3YkgVV9nXXfBF0NS1rze3d4ydxZ
f8VFlzuc1WEfsmz7rOhaJnXsr+w/lCp8RL05V6WPV+VJLxcPVODN3GPnP2nVIsTf
MS8hvsFU6rfz4fd1Oxiidc26ydO0AO+juKDfGjin1zwhaj0uyC2OSsf3xJFH2HHR
0AYM8Aze03EkJqhWsw+KoQYP/Z1Bljk1Li8J1nHNCiX5QuS9sgmNbdtjv1iglrri
0XHaQBmN+3ArJULl0YMNONGJ+mCS9weIVRRosuf+j3JDaL7B8VXBQq+KOmv8wnyX
tEUCNlWcxNCiW5qPzZ3ZtH+yk/DG52rjWmsJDOg5MMQbxyjd20Uhv+fAN8BEyv7H
zQCR8B/U3WQy+aSBF6J2TBUfzOC63bHmLUA0PL6xuNiunn2YyFo6u71SANsAwQjF
kNPMHtIS2wm90OMEanScxxQz62GXZJoaKEudueTI66wPvt4SHBaAXM6O/OFbsYK2
7wxRXDksoC2j2EI92Roj+xtMPpIKOgFmCx1cch5OhQXBNDIDEqkx7CUOd9ydhEu1
bphFXybIm5DcWsS55kAxXaXeQ8d8Hmezz2vbi+aiRXf0DYFMQKcHUWNqJOFxhVE/
h6soLeVPxrwY1aWcyAOF5Rj4yMMuc02nZSy0KKBTKA9s5JNf7ywPok+lcRKObRk1
uaW0xhxCnwIZhJEbLkAILKpn1EnJdP+YPro6qbIP6sJ1VX1YC5/RIIK7R+VLWTZv
mM1c4d8rAnIz7dxFXjCmkIm3lZhpstMI00aiVP+sClURYYxBVBBvqrvRiaUyznvF
7oU+C28WrjaETicqJCto6/RES7VKL0dG7VnFxtiJDXOd3ljqQheMG6QR5ivsdY05
lWaVXxQ1bd09Sl8qJ3kMJ2UdQ1W9oSM0T29SeGF6hvduPiIN7uXzvTqeMnxzDq4g
qu+1EHcfVimQOqaNt47+3j8Q029ewLrM8SvyDmvBzUMQvioAdtQQn3ad2FfD+fNL
yxWmkQj5IHTuUpPLTc0MbgD/o2etEChomIk2iXaFIHah00rLwVBi5WDfmMryhrQo
FyyItFzQRfhyhEP28NCQcrVfowEch8KIyNpIv6/8JsIawdnlHC0BdL71mYcdPpyn
HEETSC0TA+wdaK5JaY6QedQ1ooDGh7jUJHu1f3kxMv7WAlRDsZMEDyPxome0Ayyy
6OFyWgfeNAAA71wozdof/OaRtpnqEWJOoucLnEVmdbLS8/WrpxDZlVvcXaJ0Ehhw
AKSfJ+3MNnc5C00aOC6SKYFTAzgy343REGiJ23qaZpnfHcspUN/NLbTR0gSk2/AX
eA4Jg6DNNRfJmbEHApkIYYr+7mT2rqqTytj1wWTDwk+M7P6VI/WUvVsqSw1aoDHQ
PhCD2YZ68a+0/HCxyQYLfCh6Tstaiyd/+txdviRYGzWZ2aLJ8o92OF4kmLqxC38G
36lYQxngRRFsmEKqUo4x8jIHPtsFc/b3Rg0KB0dxx6ngl1n0YaY7qxv0fZGqIXoR
j+F+zlVFPNzjsH7KtMvDD8QsZjcRzGMdpxzeyjaOHxokN7qnTL/GDAKRZzg/xJsi
Ag0iRlf7zWB73jKruejBhHQJSqC3e8xF2WVQKRyQZqbGpwUiVgoV/A1OFafBPRwJ
sz76u9hr915K5VGwvzXp1CQtq/Fd1Uya0LoWfS+TSpf+GQUO3izjSvFNwkVtev0g
RHkfuwBy1d+s0Z+QRGS1XLCl8FfK2dgPfizUpIaGvgPU3ypRkvnSPFKFmDHCEDL2
BA4mmcPYyVuYSji7zx8JBuBXoT3zDgbg5RwMj0iyLV+ZV5L1EjfweXXGrAeKZDGO
3P9Rc7f55A//tnFziqE8f6ToeNDNa9VYvqY3U81IT8c1tzLQD64HfWPLpksGY2YF
qkKzGk0XzwHUtZHgEvTQfqRq933rOZJcGibv9+ID97EU1P8A9SjjRhCPpcErhrYW
lh0dlUT9jpPoUX3WopPB+SWlDs2BTAoEa7MYq7AmukwRmfa6PSdUW8ht53s0C15w
B6rvFyTQi3Cb8LRFGpHtn5HWIA9CTLo2R45gmnbWd3ei6MjBQkoR/1P7d3m4k9X5
97snZdgAA3Uvpapmy8VKo/bkKPZOsGjktwqVtV0OyTol562SYi3MitMqhzDr411f
wkQ7f/uwiGx0PillN+7JLd4wJ4JAk77dn1afj9bO0hWa0uotVDmp58auMoCtyq/G
fW4YzFo0L36TswAINgBnaHMz2YkXf2/i5NUUaMbvfkk3PWLXOg8jt9XqxKbDAVhX
cfTOMV69rvuFQKVaMNz/8tb+JdHQixEhzOAIxBixDfDELonOLnvlt8LVUgTtq/gr
6ROteum5ocODkZeWwGBdJTh82sFTMI1vN9/IZNkAY+FO8Wc4vRYF7P5+CDL7xo8i
86fX0RufjkPD0c62Bzlk5aB1RsC/qSya4DIOYCyZlln1J5yRL6DR82JSeeXaclgq
Cu3VmBlv6wZ7vhKZwCppg4+Mde0PmI1ZXtLMPa0BpyzMwT361UllSloAyRYo7HIC
ro1Th3h34IGG+F87orpW4PZZk04aEghJBlvYou/vTMqUF0TtjOW92huoxT72B6wG
Hp9My3PLwY8wums+E5uHnQT5sw9NmhQ1yR+eYvVCN6u6lUTNGgn1vQywwmqpac0f
howQgNxxbiUeO4SPpRH3zxuLVI7MV4AjzT7d1LqzzsLIGL+0eZOiTw23LD/H+A6n
yXOHibcvdBFaransmpITKovty6RNv7RUaskjLMy+rgVwVIJO/7lxwJPxnJ23RRBv
5DYq7x0A8GjLk4gvp6KI+axWIjSIakdj5rfuCmKw3JSJBG6uH8UCEfBaFDBRDU32
9UnmN+zRlyXgMol3nwscX/aSF7FcTl8//6+jznSugAjCjOyQgT73dkq93Bk6hF23
fR9jo+/mEe7t+6iArbW+paEMVBooyt+8nDzpTi6WduS7RHML8vbfG3m5eBGJrPO0
A1xPAvZEsWE3klkSAy5foBTB0X1zLTDsnMfSAVZXuL5XRLXGdhZbiyYRxZsonGXa
vsu1hFj2iMPVHxJjSfSgxssoidEW1WcsICkJxbgrcnCZlG1cvTGLs/E6TUE6DHry
qTKUAcv217TAQ9jadjGyuf4BPSy2Jo3+S5kYRQEnIA188f5UagDgncHo1P1H6pEE
h2jOR3G0TLhQnK/9ImiIBcnL9HpJu5ZADH2o8c2dwy7A4fJZVH4S7uZ9VLalN9gx
DSNU7NNxmqb/KxZ17l+Q+SO2t5Q9gSk4GZKOuqb9fWlFt+VfKtRBET3B20tTdLbC
w7kgt6PVcwBoiGacFuMM75TnyMg9B1tGB6rvgwPV1JWcCndr1eBKOYGULqqzMUa5
MF8BB5Qlc+DzMMb+RZi9RhqBKbj3hzJMlM6pseLik5LitAgu4Y7nQ0XM3qFa2CIJ
sgOzPecGSf+JQTueRqZTVtwaTQbyz8qgW9I+U6xx+diPePyW3EzOPEtPJjrn5qSw
SbV1F/E7MCotOY6AOcUFlT/ucCxvwdSbOeSM39ZsmCcRmsCusOTaPao0EYJua0Jz
T7r/uxbFhv70XBK4xMeM17kdsDucHvzZqIldiU5b7f3jAG6I6KzEClRYzD7q2sUW
Lx6hVOJWOA3aulLgd4qOJFS33SIBo4tw3AgMxg2/iAy8RIy8bxCbAo1ssjbBR0er
OzXxdnXTr+vwE8LlfnMe0I/qAwVMP+D6n4KnbXcS42EtJgj7+xDw8PIw+ULxHkMo
3kcC6D7KXfTUBBWenqH2toXi49o/fdHtmNDPcZo6Qabl2UFkfr5CNKhuBtkT+T1A
Zs8M/gJUauWYiocLeooULJdJoMCo9jxl61UTcjq0yduQdLXaogRjfPk2W2a54NeE
PiihTUm1rWlDdRiA1KKe/Rn3EFSvA/8ou2jGKisEY5UliksabE19igai2ufd/yXb
EBT6OEaZF0OA3Oq+K8aJ/gmP/b1XXRv9FpDUbXxPUq+1Xk790QVHAvxsD5Q3BTYX
kXiylv7lh2xV87UGghmcvwPqtgxt3SqgEuiFqBeDM+ng5Ru1qcxzYQ9VFEnjgSSj
QhXDHTLqJpreQ1jyMrLUVyaWvPekAR1tWpKKj5IT1aLYgzPZsZsGwby2Jum9qRsS
V0EgJcEwnt90GTW79UTY5CTpm95YudkLkpu8Ha/fHQHzMmuKLY8LNvIiQf4KvNmH
C7clGSFMab+7lU8XPJqukXJtbPzLP1yrnUQNgeR60EWMIqwAznp/FW6DEZzpaZsD
4QBzyfpCm7wRQBDVmeYTztZX1YQORwXGNj69r4WYRmzR52g9wtC4CnUl8DqqjYEp
gXbYcepsfrwOJQlIY/44u7uAyryG8WM+lCC6kl2fzTMDINtXfQ5u9rrwuTy94GNX
GVgWN9GwQp8Q1y8LIU/+Hq/qeAckC758dRgnUy95a5w6hOvApyJpb3IJbzR6WAd8
12vbACJK0+YEG4YpKVwm/Mdg0kqD0PHqzyRGfp+X1SQcGKqlarjeWaYBuY4AW+JU
e0KxRl0GjDFF8b7LzOwBsan+QUdwgZSK8ZD/HSZlN6ds51Ao6pCQrJONbpOslJDu
pFVgky5V5UyNWVQA5112juDdrKjCgurgzYzBiSESBBwl9UlAyeLHe3fUVs0LTqeD
AbK3TJEZzKQbn/BW4xA1cNYcgTEmmmEJcw0PY2p0xIUe6S4+7UHHmwHYW8M+beAn
+D0lbABO+6RzmMVIqfjdgAuSpod5En+hpRQsVpTzlRd6tGf2jyegnQ1T95t42bmf
RGQ765KaVQPM5OhK/YybWsT5uCkxdVIMpZJYlXF/ijCzwdSLTFbEkf+L0TBWauOY
roYyImvdvTGP9VOfUvskWc202Jt/IGziyD79AVVSUuiErS2mb/qRyKpg9IxwPayd
Euv6JA6VQYlBff5eSGR1ufwMLmRAhUMaee8nKjkby7n7oyVRJpoH5twQiKISNAS2
Qs/S4wBp+RoJrHMnStrVQYDEznO375NV2MUO1W/QyfyIsE7xD7q7UZz5skYuDpyV
8abINiv1WF4Mf3JOVg/JqXmHv5mnbq9YdrHyL6R426UpbYwsW9+WQJE3eTNp1Q9G
Dt1WOMC0mhGIHP7gcwgWp2LYUA+b1ZbJc0GVsHwdaKn2xda1bwwyBhfhIbVBdaYf
/dXd7gDNclOyITWQY3HM/3iRqeFyVAKnsF0+9NJfVvojQfoMyakQeIWVzc6NRYA4
kaV5twBJaaZlwU37MytHTuLpyMEMo/gz8wE5yYrtSY7nC4ZRwIbm4EIQ961FLtq5
q+4ZzvEXSINGTL6jwmv0eJmraQdCfkO7BmyafOPg5tWPaIMLNnDkZuMM6rG45QyP
MUhyzL5Es7NW6Wx7Nyse2zbjAc7GUTRe3IeRrjrCKCFmhteOmnAJmQNLKfeE9XUI
RJktKxVIZNeECmvZvnXwZ316gilSlBSAnVUyxIcHV7mif41xbkq1C/Hlcziubc5n
9rADXwtHv4GHgBZrIp0By6S8BUfc/Js7oLzMUDTTZgpWaFldzyjuo+ZGwnOVdCRz
OyeiA9ZGfFAIp2YjFS6cm/UCcMvgmsp2q59YI5ZZaZd2jjQ48kOej8uF+kHLXiS5
Nb0o3OMC77HfdQyiwsL5gSLysEAGBtehOg7A/M7oBR1aOE1HTCXqgdjwVi4QtF9Z
HGqYdBhDj7VjI+KhfWhSrRwon+qpoyP2nhp9ZFiIfTXW9ma5rQlFRPTQJeD/d8fi
V07ch0nDilzvUD1VWUPk+XtxaHj9oRAKqVdV9oNV+viwYhf2NuG8YQQdu62lg36a
172dBXsnvwgUkGhidzGSO35Vl80JjuasRKbVetw5vbu01P4/Rr3CjKs3tVFBsBJo
LGXPhPN/sxt4n1SKAtqLbb8F0EmnElXxQ74DQrkCU9OBjENBatbOv2r1/Zuct5pW
Fp50CThY8iK8bVuHEkQ6spDBhEZohvKj8OeW+PREuLSWsxnE9qQgimL1XL0+mLM5
/OY63trcvbOR0+QtGAFBGswx3cchrjHZ/2IVQx1d0Cijz/qxnZVdOJCbkaKCntPt
J5M3lPcaUue37RTkv0fGYNzQKJc+alC85QzLwancDYXwJ3mcDFRKed9neN2640xY
eSw35jekU1G1mwrBQk7BSaUOYEyQn2QGINg0xtWtp1FDfnfNnGnOZ6SYobhr9xvp
20gaRSMESMF7bGa0nVjr6Dukpjx1/z8fTOcoHiA6Cl1B7fZb0tLoepL2e8icE9DW
rG101+hXWbqanztOBZ0a1mW46duXMBYznIk5aiOQYnjqHw+PlV9bq6+9d5ltcU+R
qQuKXLxmU6MA0cVkKtFhW3GkCdPJvCqCBqWp+6oHIJ/SHq3/5kVep7RKZ38t/XwH
G3t4UAQh7cFq1y+cfoIzLIr/iN67PMqr/WqqsN0qF8bYel0wNnlJw1l6rrNFIVW9
mOO94gpJAxYJ+gnsIMWOmoiHJYMYHaH7z2Y8LmtUtqEpDLNav5lDkW6qxJrwo+NJ
lPECtznR/nPCIBFASrE/PIXYej2ZG34NpQzx9COFjOeBzPC3ZdiKXPMdMINHrD09
XZjb/aujTE8tXKtGfFccy2CO7jiEv1Wz0T7BH572wq0MGRIdCl+CIxFeatAN5Ad3
aQdDHnpkSBz0S9WneFVVWEr1jdlPZpjxugBBfMXprf5ijVX5+r2gZssGOx30lqjV
d+i0KgSIDpOIDRhuxUlF7sXU/rJAOeZN0cVtSyubCBamlZvixUo7apF2SJTuzoZ4
Pl+WlfbCd6yWyRrxxFLc/M9z1hOqnVTBb0hCELXMrmapsgdllm34IHHGS+3HK5Dl
FwKzzCKVUTdwX3n0RcRirsvAOSN7vrZ/7MiAUS+MvpnwA7f+VOwb3GiDQrAKXIN+
mCrfYx55r9gDkpwZgNJDSH7nKLcwQL1ShQsmpYzlU7WY4JBveC9mG3W7+zPfAhz3
25ia/CUM9tP/MN+lxKPdfqc48oiZjr0pMYepLTa3CvoZ14dA5jTh0yRM1KOa1b9k
bXANmOLMi3cfkqfsc90IDAmWr8t3RbEQccvAins2kDjNysZY7sDeqdH2iTwG+CrN
pnf8K3Fel9+qpla+tUZ17MgYBmujNSZhP5Fs1JFrxl4xKm14rFPsjtQO1dlksi6q
vPYGHdl0OCk/4VUVPJJ6p2Xe67WHi1g4QFfEuU9raZPJ6VenasALldxGB1iEyJex
MGO9gBz08MpERDzc0uHqV0U/ndqNE7OPr3ZZeGiZnewDqD8CGCQUsKJqaO8f3yjA
dEKNnsKYxasyeKVTtqNeoYRAkUSZEnv2mCvEcURcGdisaTrCGX5SlQvStgiKvWtS
b6WbykI/v12BnPrMRF//4phnE199gjxvhpmax2PdOD+MK6j/8RdJ+1uJRnkf/u3o
ybaZZvoz/FWt0qA94wTKsckzN7eG92BDa9MHIA8kT2p+1Eof2mEzxwqs60RJ34Gx
9C6EMxmywz/8WpboQxwhjf6dP86fgxiGjAOzFwRVcr5LD4TX5x1tRgRFtGYf17ij
kYWEgUJVQ3Q+iKez27CUsWzh/c/JHHulBmKDKw6WVsrF29LSw7yFYi/Qh7PFFWUu
QXGv5ipqkcRsAYlv/TuORQqgLGtKvAYKdoWFe9LDDZuXqZgubSfL49/zvsvOxWfO
OuTn+w8lTOYAHw3khgs/U12wCEdSB2Vml/+gpfCrlc2pvIofQZpH2V9kJtB8zqAz
C7UCETY3QjB/w9D3aDiHh1/IC17866aToo/juUjw/mg9EQENh57VMWGsSinW5uEz
VQEaC8tW9/vtgMFCw8oMfGJGBevFNDfJzJ0pprvv1tVd1U5b8xj3B8B4ctJlOBUr
La0d7tL/W1rlwvmL9ivpk+7HkvP7IYT1v/I+cgdabLNuvog83MjXa9fbnBuUShSg
jwObc4RhFK4GcZLLJ/CQT12VVmUb5D3Ft2/OUbWV0MP4lodEPJTl1qBoDQxks5Hk
p5Lr7h1mtwLDSh2UoGdxCWcJjfqE/ePROcHYCfDVgZUrAdAGIYmcuti4mHhTS5TB
qfhK9zOP7UCX9hoos1AvJvXKfKN2v2z3Aj5dygIKE3699oqKQCqUkzvSqT9IV0uX
V/kCnm3qYMBDhhlEevboSuaetorXxNsch0LTQjzDPgFG0t4z7/youAX6hWSQ5ckF
cdHRIakPPvj0g24w95BmYk4oMEPg3Yi0ADbn+XF4BTeV05S5RaQ88MCHIR3yd8gG
dHt9E+1EdNwhE3jQELmXye+098mq6DMVq/hsbr46Tnt71GX5yqHL45L+zbnR5NWb
0hXSH9EP2qgvkhwkK2Q50nPoS3/px/arQ7NhpzFgPP27YCPEea/23sFb9AdO0KS6
Kw4lUzXfnYMKP54Xi6yWKb1Uw7ADyJOvWHYE/8rCufILIUrXs32+tPg7TRoTCiLK
mVdwiJcoLbyCjkcX4GbffGPMGh9H0guGgoAV7HkRaf3zaVYf1jf1ycMH0UF/sjsW
qwwi3knETKFquJ4me8R5pKvDmuEyAVrt+9zOnHaIPxSXVcw/iivb7q4MbBPUgFhg
zZqvIn3O9S3TLSpPPRA3RP5noPclopTGhqlhVfu7YTFBSKLDM2nOZNXLmL4Ukaf1
rtYgpmHVCVdiiYXY8SS9uG1b2mWxOcG/NQEepdgMEEFcVoo34mf1ZLSnHdh3hu/w
H844xBlNTY43vCUj1Huulz38t1U/UZR7Kn+v/VvHC9fF1fzgxW22QPEBfXa3H7gQ
VCFNRgXRR507h600kDKEgELo7dUPUiQwwWPZk8t9wE5XDrlLs2uZ6cfCZK3sW/Oj
pPpKdPYk3aZtsA7qYOsIlyVa0A6dAAxmMJ7MJaJcoNziCt+oci2OMhaPYivMXtWA
0Vw7zjl+dkcSjq1q1tprfzRUhPjzuj1Cet3q8XLRRHsY4P+CIHfuSBYUQMNPcsUO
OdtpFJE8x0UAMUySDUg+XdFUaAxU+IW+IXxytLokKfLunQybe7yGjD8BeRTUgZvz
VNe2lq/P4vVq2wcLcgYvrHvIZpXu3N2W1ahJLQ0c531zQ8a/p8rxwhI7qt8v3mfG
JQ/w3Gb/E2LIAuQCHVM3DZmflZq7Zup749MQ+dg1XZkCKZz+QUlgT1+ELhYpMMvf
Btx1aucbLTC5r8KX9Gy1FhesPm5JJ0iTVQn4xsYZxWl+ZNE+bBfnDJ0DqAQeRWdB
mOGZFuwBi1tcEUFeuhiar7JTjyV0vhBGXmxTy2nYq3fNOzAwMWeg+Wp6J6zjYcJe
LWXtdgpzPfWC9hKjRgxA318+aIw1kR+xKpPQHvXV3g+6ISOJZ++D2Q0LWRkmfwjM
OsRcjPIDI/eY2LwMOUnBMs4p2Q52B+7q4OO9PuoyU7ehRp3tvi3WSVhTd3Kgwugd
F+rZvqvBTTJ7PBxPzw2WiD9JeqzVn/YaMAcf9Phyw41A8yc56zuFUf6cOZmlkETR
8NiJhqm7rXKFzxYdLmS6FHvYEo94zuG47BL4BGycHPa/NgOp14LV0mAW/GlHYFlL
eCkFkzWzY5BfB3NHcPgmwXPldbtGQofJr5Q0vXvxraHwnm8VXpYup94xwYDLWgV8
Tt3nQDJCVx17hCLbK9d6lKYJ9LJYd8fmAKWcHw7GCbItWEg+FO1ptxl/RFmrrwuY
nccLoMa/e+3zV8parKVmdSV/drEAg5gOwcmL7/ZHBavLz2U9gFL5ElnzhrZB5j/a
9H8w2hijLfYd5Jlqkbun6DIHnT796ohcYz7VLRjw0UcZhr/A+B6zgEegtM6miEZm
n3BW+fK07e1gEmLjsePzGCz+bM+UP1mfKqxED2uvXFCg2Qf1C9eS2mPHWea53v00
qcNj2UT7c1ptMA8tlDJv4IFykbSgKUELROJxkFPDlCGocJPq0s0FnPQ+k0NnOLI0
KSqUFuptdAcfA2qmsSU7Z5v6QEKalTHydPVzXF1rV/zGeABKpb0+gHwnV8AXxURc
lXBklDd+9x/oPOzmda2rYOoXDyb/5yfaUPNz/quoi4Yv2zAZqO+EVVparP3XiXCI
bMZHN8aqyDhZwH3/5IchmAa/Xgsw11UTQ1N2RSVkZAPdH9knkswTK/KhhhhEZdfN
nvlQUVLQfjAEYRdeILCpXnS1tMqchD+ZAnKqxpLIwMiPI4A43DXrw6lyRbg4/Jac
xThNeTVqP2JgfEU0CCaTUv7siC2IIBbOSEv5TWiqlpqpVFu7EyXd2Eumz2LUKYvr
JKheObIDOwayZgtA4W0mLAydaX+/melC/fmRLno1SFi7UWhd/rLPSAysuGLoAOl/
TR5d0LowPdAr9E9D4OwfVSwDxPSkUDs8G3fcKhkgEtwom81ulVPrVLEVBmia3YH7
n2qstFJMWLEPhDqW128h/ZKWTy7RmvsUKr+I2cXg8Xlg+BKEZn1/xnIqortxNUUO
paxVyI5nHAyczGUs3wCQJuLHphYAVXnmCj9S9pQFEFvu7NzUlvylnoWkFBGBVA2J
PDtVHPOeS1L1xpQMtM2caX/VMMf9tp8WOfsEq7TPfypm03+reT87nxPH36np6kz+
lm1DYnke29ufRPVOHcDJq0wbFBfr0eIlfd8fyOwspI6Jl4PWhhBJU98nduOunVPy
F+sCYIUW1yrE5vvyOGIxkGT/pnZ3uiFYE6mYY/MXYlUgMePUz9J1ar+be/kvnLF3
D6nB6Mb9Z+9lroe7XpsnJimIoynDmmeON+bZN+edqe6+7zA/C9a3O0E0w3Rcd42a
EynYGCGvxun2l/bu0bj+qtZgSX9X/yxtS5h3QE/OoReCV1+HT9EZRKhsv5KVwN48
DAUUzW61bfbwfr1hG9DBkKXGdVmxQOC+2bx//rTRGQUcmy/NHe04K5VmOdKuOR88
LQvf6ipirYuqcwhbUYwlgXFmidsiuz+t3f4Z3mqClGvTy55KDGw/cf7h2Qw5gCq2
nLEzkUNEevswjXMIxlBWbSkSp2EiDStwubEt48F3k2uq9vts2Yq2loAlVkfusPIQ
qldcORtijlHz2v3QUNiAIFrpMaKiTNBhRnM4wSlJvqJDAef2IvZSAkog4kjuRKi4
tEQz7ACJhebZcouxsM4x7zYwO8BGgg2Lm/Lx4Jd9DOijAivvhh1JEXyTRFYpafmf
PRURdDJDdKWcNV4OOcvR6aaeNxkej3sVfBJXvxzY02E+erzq7qD6lyqt1rx41Mp0
8IAzW9aN+2odIX5GMvETxx6JB43+tAJM21HGrT/GDggJA18FxRZTL4Gsq0cdWGmx
olS10F4b5vYdHKM49uJZl9uqFBEhifxg3uRd4f3rMtqbHv+oBsKir5UTg8P5pyX5
I844bvzYTovnnfYyJPinHTmfQqiU/eqIwUIcC5NMODICohTYgbPWcrq/L4xjE1A/
JKebcV2M7uq1jC1cyNPdhobkUiEelBtxXiTfsj0oeE5kqtK09L8YnAarlm4OKLlz
xgES8P867ArkpTapB4IcTkQ0tji+9kU4rv6hsvwnmevT8zGbV/cHjHcxhKZtYHuU
ZgOmQVCkEo0mC376WkjtYw9BQAgSDThfriVxzIQ8b1YIJraQ2ySZId9oiUdMd66n
qzrf6zb+cv2PthyojUDyn7dP7l8GUXwSg7z7P/W17USxz0z1V90E5Lk9W8WdzqVs
BIDtLxxXFTwS52uV6lBxKAnQYmET174JdH2miBGCdAxBl6fsPORhLWZRXgeTz1ut
G2PD2Z90N0ZfEN8WqdfUvC0tSdXVhda+pqn3wnzNAVtIENyBMkmToF4D/bkfE5SG
ooyGnyrItHvA//BY5Y9G7zd+niBjU+5S+AAMeEP/bJBtgvOurbLe1KYOcUYpPAKR
/X/R5RauOMIjomxJ2FE9mhCueZZCLcxkIXcsUrgR8UhzejczLL0G0JyRxaWhE7YZ
2IUguozAUm282+PTJHPxX8ZNcHAmkAv2ikBUh4MwoPCoiLQ1+5m0WHottAv8djdU
6tsKnTGNAzW0DNKt/Kh6Ndzh5HapeFAzLogSJCfBI0uzvmzZT3IgzDApNfX+jrVi
f10ujZ7Lib2FDenOVR6+z7tUBeOk461FwvhYpvDm61Jb9jIKq2VjBoMkPuxkpoOd
ILDUlhQvxxt1Fr2Ti6WS14R+Fzix2C2Ld2eAqQp1DZzYDNIGQU44LOb1el3qFksa
SiRahr70RFguikkNNiF/MWoE5dhNyCddMQ2TMx7MUBDEzw8lQtQ7+HwQ0+lMnihU
dZSE0Y6hUqFAa1b/50zb2tYHU92ZEv2SFjxEZ3GmQtA5CHW1Bx745dGcg/WM4CDK
4l7wA7ajO57AdUx/MnFOc0D5IMtMkYlfTIO9YCD7jg2hYM0nGFujOhcNeitLQ0/a
6BoyLXAWDcCi+Dl0fddpQcmaXzfusdsEdr80JsS9QMztwxDcM386NBrlfBiMXgnh
zkIqV0l8/Clb2WSsJu2eAxi7AUQOAFESjR4jZl0NIVV4vKJ6Hg6LbGUJPnl++ltO
bLd2F3JtKFUIoK8WKC4C3SuPLltLriRA3QF5xNNy/Ok8CXlOgPT/OUbZU0SMU9ar
s0QQWEjKOGKxl7ODbSbqcR3I8cO2sP2L6dQLSYiLVNKv650X5yUxx/EH1BcRczRS
8vijYOqLpXXlQdvNMAF+9Ua9MI56P7iqJIU1KHBwZqCPDHr63tCC05G2XHEptfXp
+l8eSGHgWuiKpkJbvMD+zaJ+KJV+0WNottHb69l+pBUnTL/6Yj/9yh9U58WxZFYu
mB8ZZR3dXA9PrCRDOjiAVjyL4nM49zVKvJgrBKm1QYuQVV+zIYJnjDokWD/e3LcM
fUMyej3Dj9w4FcmZpspABaspbakvWOZO91h3b7icVPImSqm5ZkV7lgslsql4aABY
i8ZixY2/IgTYzlNjHUzp+XlI6CJo/7MzVsB6BDkPJbKvSnWjlf+9snxS7TylDchl
CmSemGAjabGznJVs8tcMCagWqLvUPmyvgPx3JnAsLRycYr5qyxm1YQNB3la5cyUr
+23dc47kHH/fXQo9E4n08UpU+uECVCAuCbXcniWrvuDQMqoJrrL9YKOYrNvLnc8V
SFazdUnhq8kPC0KbiNf2nlxBe/7CCyzhPbFHat1GMqbF9g+pS3TCD5j97rIlaGbP
3+NL6gq7JVIh2Uou7pm/pK/LIHrbD67mmcvaaYbkbhwQqL9PVJgw5RPz9W19uyh1
phiWeRhath/mD91p80OtntfDP17136z1bOaJbWH2KidobpHwP6AyV3X5yTW4YMQO
A2YLEj674ctHil55ul75YbMAKja7idFkE/GkVqjvvfgbKowAHQsysHs79M471i3T
erOIo/88AhwISUVrAPkdeYsnVBXiuUGlWzdomdNsNnVrZieqeQXBKbHJDOup0L/T
Z/OTLLXm4QKhQRY+InJcy8ycrvU/vv6/rkd/OSPqlP6SgckOwOGpj9HXgfofOk7t
gacDgcznd8fpWWmXIJJ3dHBbjfSUYd1sG58VwfukvWAQPFyt9YpTtT7oshth4LAw
8AS7wgjxEFCvAzfRiKUs1tbkWMNkSBTUjEi8ULGNja5yrb7UrzrMqJAEm+pDkQ7S
tNF8D2deBrNkDK5SVyPhCl62VyECULlfP2cXq742A7R4TnSmqPrUn52kFr2K7YfK
vKfUMirnwpfQStPrrmXDwDfl59yZLnyakv03XlpV8OoXiAD9TEMDKZoSlSn1zovc
g6vc8qudu0WBOmNcvOJhtmqYHvdiCf9zYdJTsEenCt8hoG6ivo5iPzrVuoXSMVsP
ABediGk/OjAreErRZSrUKLFA0hZ6SLj2yO2mOHi5r8Xe3VTNq1jN2G3ZvIf0v3zl
g/Zo+l1SLf/6ngS62Sd48uDaUUz4zSVR6bwu1Y3Ai2yl8He/rkP8BRpzj41l24H/
niiFPz06AhonEN+KCquSv9K6HCvWqj72gpqcy7QFDdWsfIIfztiQQNdi3rpKXjw3
1ctPBKA0UxD5Y/vs1xbocL5C9FZKJ6MNT75zvv21fGexgzSagQB5vG9I7sVMFUJM
s7FSZwFmg07hdMoLxanw+MSNnu/zUWH8R0HXvlZeF9U371Bv1WELmyq1RCTp+uGG
pXPpehWZUJA1uQV1J6Q1jAV+mKiJE1IammC/Rc5a3SKPyS8Cg7DEDU9dp3wsfjUi
/9URa5OxGJyn7YZPZV+t3CHpJYukGkUGDECgXUrcux+89WYKOLuuEyTo7gzkxtrh
gQdYoRvlP3OmGOSrZ5FFpp8fWs73a81GlfBwsxo8BeJtK7bHpcDEjFqmeK6KzLlb
eMrrOThYGmBIYPu3qoeXnjI/qGA79pUdKZEmUaq2ygBzJCnSUeDn27xYG9k18m7j
2N3DWR2Ja06esoeEMjilY5lJ8gbe6rExc2/4iNogfITt6d9zFdVF7gBYNgHUK+5Q
B76RhEJzmu0EJHVEmli/CEiDPw6exf/8IAsjQP5fsOqOl8YlGNXLneJxOSxSyRmT
eAOF94jinYKMDwA7zEx6JW1xotRD8R9tzJkn0fu6085l216TsZ76X42GtdCaNL5y
Zmc395fnqDpz4WxBp0I82c+brKMusTKiJzdel5WoAQ2hxGNAriqJtQZ/FHXQO6tR
mWxxZQISeHkcdCATdm7K7EU/N09GTwm8LF4Mtp5N+H/TtauRYYoM94njAQv3lUko
PyDlgakbk59rseWPneWNAoywfbkW7Oebj1Wm4icn/Yg1jfaNa1G5NwjC97ZBsYZd
/ifC/8uzAdAHLFLDrT7wbtT/UgSxDcp9TV3lZ5triOrLJYbriJw3wptkZka1PlUr
nUYk3DuZXl/5q9IqTkcjadmTAuCRSGXVkp1RJ0MZy2zgp3rX9DEfr8ATAX1sofcv
owygrOSn3PCKiJES7M1l3oxUL3WZ14XJpRcQamd9OLINYvdVTLX5WtaDhEdGnI/O
rHp5PCpdOIResfITCX8SUkCUQR4MWwJn/tnm0nBZYCgQOfJ07PyFvLCKHaTTEIZb
vbHNonhenFqXLe7EWnwTqWwQfl/paRy2XC/CpTt441P4dEhJ175Hc970uyvzBwlh
XiXYhVK+6OWBtT2RDLq1jlJAui3YAeW8dQJoQhtXkDrNfbLFFbgwYo/HQV7VptMP
jckw9aX74JHX7lRiV2uL5p1QEDUgouICQ2ueV11XCUIfyXdpZPxFvPUtqCsE8I3y
jkMA6bjRGA60+p3kJLhJk3yIkCwZ/jxRIOGsl0dnmQ7ioRVRxmh4zzOevoSy+1cU
FFfhuP85LsKjER2WDfOlJMpUPaHWMt19EBiJfTCmnlIIDURdHqdZuAq5jY3w+ZF7
YRVvbrsgTFMI+CfQtuxQm5D4t9C4ucMAiUcf5iN491kwfNrVBSLW3oHxxdoDgI3h
JJBXr8i6uO6EV1dduA4vxn0pjGKG5fGrIKli7aEzEVrh39/VD76BtT1Rj0yfpiwz
LeQ6ne9aazwBwTwgFA8UfTGJmUxZefRRiDG2jbMi+yFPG/iXPMFg9JGc8B2fxyWH
GHi9vSO3ZIetArgS4mrrF/HQvSKTgixQ95vlCec4wZqVZ9+TrQZYKJhV3wiNE2Xt
6eKLTGgE5E/GlWlPC3yqqnBY0rE41owh4I1TT1i0JgiKKLJhA34mBW+T2MztK1Uw
FNTrFp1tQap9QdijirXK3GZ24IwxYMsVq6sZX9EpmXMLuTHpz6NmdJPn7EGRfoe0
6GXnsOPUF3kSwr7GerBJWk5GXuaLmGWonXBxlQ36wS9M1fqkdXee3Rjaz+/QaksO
aC82L4/Hl9tW55OesrenYml6ZIKu/IcnALct8cnr6NmBwTnbinBWIjN6QR2bqZHX
TFT6VFOcj+J6ZAC2cmCCu+erROFmVAIRQEdR0yuyujS2LZAroSbIWZI2XJDRUIxd
RWSPlLxGjOhgembh3Gr0riAgyDQChocXOdo1BIqF3ew/R4gn7EZ9HfRCXQGo+1+u
RncRur01sAiDtU8O4hRJrQ8x7aaVJGqv/9IFu1U8aeODEpt+fEwgLgVp8Euzipo7
SuawdbLiz8DtCyO7y3lAf5U3Ig/EhaSJfwO366+ihEklz3ccZd7Q2PCHIBortub/
9NXBmIcc1BTRx4mCEU8Roa9Xcv9EhQUhSUJZh/DvOt/qDk0AVErh4oEqaftUCBwQ
W19s8CJlrm89pn2ZbuziivJfhebbP7LwSvMHPoEiHh/YxybQdC3p5Pv7Yc7iK9Q/
sL5CZ2VYAQe+mgeOZ8Ivjq3VRQCnK9Ii/1vlZnp/YRHf1bsl1+tEgNgnnGJ2LnpD
6UFUaPbZfhI+E9VOwWpFyq6Ug5wnzkniHv0Cr7SJDCY3R83CUlhOZsoHk9aDoQBW
8zn3UvqRqpqL2VtCq3NIAuQvS7CJGhyV2MtuQMZBdM7WPe++5U9T6KN99eiS5Xaw
b25FwohiKrgbBWARmTVR41asr2NA8eHDh0F33+W/TWbVKQ4bLFvbktZDi1C8i7gp
NSzDdfhYOqoRPtjz9j+J2krt8tmHhsxl9WV/lp9vjptPYNUVnVwvoun7xCCAdAxE
KiYBNOCueGxC8RDa5O9Y/LTG/duQbbOVosZqHll3f8LESlQ6IGKls12UEbfttrho
iYP462rNFG3c3CAlzvAFPNGn9Z3sjRbxdPIat3CVyLS5zNDKDNwGFkldnGLqNocs
1yce1Jyyl3zvON5NqoUt7dc5BUQCm3A5sNV7rcqiaX/gcXQpQ6FKzZND9BUepE+E
VNflhgR67Iw3l53oPo1L0cCkjP3S9oYejK+PwEMtkGOoYLKX7o14fxsNQFUFU3Kp
v3ieTYwPw3ovSyaeBH81ISPD1UqXCzJBGgpwrz6RC1O8uRSVmeLYYdgj1Y2Iicc/
5duVHQDiESBhxsLxhJvED8nbzFAL7zR14y4sapndgYn9EH2d+lk33grA1pd8am+q
rRIZp+da+VO+p2HWWmvUx9xSI4QUOA64AU/HqQRKqxB+bUt4n6YO7fTexB38dein
G3kcBAWAKCVGQVIaMp1AQL+lDSJEtivtoQbYn14OTrQ2cqFgsjoJh1JXdLKUVkCD
cGyoyyEUrvO4MdXRao6lUmRwrDrdBkuRlIvvqIt4FfU3TuM7sNySOOvkwLrLdyVE
8t/MXzz48gSY3veY8fn32TCsOSYpNphrIaj8MvYBJUbUH3fq/Q99smuny7PCa6J6
jjwaZEG35fWdsI8iaSCHVW5l7l0m970AER9q9K4JleeG+MYQKpVhCenwntmd82L4
EY8BPi03D35zfxoFovVeA0JfYldy3muyE/gD0uY8Xgj6IPHyE0DgqQhXpkv44VTv
iT6VSG1wyH+H+zDgsG4G3YaWXR5snPm4+nbgDnFXh4VP8gCzypvf78VDX8A47fUa
pkJDU0F39qRDHUqjYC6a3G6AT+vpEgl+TTqDfCZtwmTPlrPZ1ZLPeoJFJ0OmQxo8
uKkhsl0sd5WfIx76C2Qzf75S4HzA/9nH88tA6/7d6mYRXEv9+ASY1o/fxuryjyDJ
bXNMPwVw1/rC7x5PbFWXDEtzi0HvSaV9dObuJsYEGeacmKqtBZ+YiEqaYXBDCP6i
l5ksIJH3osBGrVhm8k2G6x3+8hLkagsHeqcqLEKfTQ9K4+UOhgxOnvhaGIQnngas
GNJofrXSTUc44uGwHSsKwVYUqmLOWMkBx62T/OY4bypjzDXZ9djDof4i4QmcQs+d
zwljfb3WfdJpJMbOlvUUPpKX0NJxKaZ7orhi/E5lPVFfi81gMZ7GvbMyE5YalN9h
1a00lu9H2hpnxcUIBdNxDCr8PSAI7590J2GLWJx48PhVPQjIE2ctCizwc+3iqypf
i0ElY07QUuippG0lbpHJdD3JIsImMfb3h/mTtxarKcPR9DBYl6LRJmGRPUxj4nXo
3B3bv7mbbi9yIeCnjzcQiwukC9fi5/rejIGYCFEATtihDthfjKXMqOKurVfcS3yi
Gyh1tA5oIq+19MoEn3qRGCSPVhREUptstTfQFWMP52J9TySZeCdkqOx7+lZ8Mcuk
Zowgrgb8Lw0wK+kA12emF57jcTdO1TfNFXlcsFq9KDEcY9335hSctC5n6te/WYpD
cJ7tPJ04hU3BTt6I0ty/dMPFYQaMHpPW9o+RRBY8ta0LUh8Xa50ktAEaVmHOhZiy
FS/ZA1vYYKt5xpj3ZgraN8IweoHymWjPeIQx6H5gX0o9FgFfRjCxiSTW1wD34Knd
oiy/NgTBSz9gbo0Icy3tYqEaXYYrnEKramA6etQVCYKifQlUB4mTiQ05dNiGD4fO
vh9fE2qzMQ4cYhdr0ShcerM+QwFs8qsTYzoVZyKbJJ6DuYrQqIX19QGFqSYjSMxZ
/whfFJ8Eghkw+EZQ1ecTd5cg0TcVNIjeOHHba72tAfVpOQEhYpEhVFxNgUpbjfOf
/F3jS4vyt7TZCsGClUR4cUcn7oXhKI0wpxQ/H0L9NPAOoc/l1PpLvhne2Ket5iG/
0lnF5fT6fXJiV1WgYbZnwUE6dqQEDz1qiQ4tHH8KueZV176RsBHjEXqPZPkc4HCA
0R6ZyREDKHq75C+4UZ/7yE66zc0wY86cRNAqFbVMzVu0Ksg059rgfCxDvXkbUWCf
skSo5HJodW96sZFcSTzrV+e4cZcmDlyRSrSJPQovn7XT+2GnW9pszwhbysgGxU82
jcwdsQpn1PChXPeLS/6wu6hPXuIFRDYE3WrRtvMqGwH1x7bt0XOOf3wnlHDw3B+t
Xy/9OPbRr4v/kEPy4xxWhcR6X41xKIuhgfq009IgaaZFql8P5f3HNWrIpK0WoGr3
5N73O2MBCTE3H6ONRf5M2meUh9LScX8EY+F/tJQIB1ZL1Q3YhFWtlrQQXFdm58gY
RLxxUPU7EfFlCqqyt9TzWBNU/LS6p0YVFmjvft80usp8p3hu5wI8ysHyfdZsWTKU
h0NiidpDpcZhXCsh+ZH/pFN0sMpcQ2xnNTumUoTRuovWn/Mba0sG+8bkdYFC3GG4
11upJxUTQh9CMq6Q1/1iDoxTJWRrhP0lbEy80/7Zz0fZPgVmmzrwHFhlXdR0deLb
VTVWjd60eseaAluS9Qr4xmS8VTjlBGV30CQtNQQm3EbLXijCMK/f3rELT9K1osmO
AE7yjGWiSUSIrdapJSer66CFPUdKyFjZBPjCTxji7/dWwca5VL29Vm5DJnR/yi2M
TZzEr4C6AeMYgfaJPu0rrMMS+JF0emWzNgjm04gIegGpQwaBWMV+At+cM2sv/do5
g2jzBPQtW3Lcc2Gl7p6D4yBM21nIW6FjRfUsIMbXNXwQTvp/6udgwYNse1FiLuIA
Kcd/aGGxpVT0C0bPsl5UK7oZJNavo57RCI4/X9WiHHBEKXSscGhgDffZWKvyje5C
+bhyP4H7YdL2BNKeer2BPjb+5f9/6pOBi30KB7S46wL0V5xWeQUmmElO7JCT26Qx
qFfVzR4kxuP+aRkpM+TmYLyhfHtBUyF9Nh4vWblI0Bfdc9ZCC52hmsZwcmWOYslb
EhQ+gGeNmNnGImAvsgzchMRnfZlhJGUEc7F72Wvjr6JBDKiqUWrms3jLQfgFV7zs
i5efY0XWpTp8/Ora8MjJYokLxop8XMBaLzdhJDgeyejkNV44k1j07aZFu27yf2KC
bvGJiBk7dVBlNYzKO5pXdoNpi+q58NrQFDcIiStzLbXtukq0BJx/Cpr2OQ89BoaY
Jheqi7fkKxlNwa3e58WBHJmllF8qLbXc8NGrUQuVGdDiKTotLmN4r75x8N01pWZt
rICeXhpOLg3kMgBA8VLeaV5jWvBvQmXZcIg9KW4I2Aabpg2LsuW40unsQ8O4vOIK
3vi+chDx2/sEfr2iDQZHLChCmv0pwbgTbsKukU/aiaqXKyIbuEodKx+1GVbT+dhk
+ox3VGK26pM3L5+YGcGu3JNUKUYyFc8btD5J0qIlj3VPLzXR3oc6IEJyKuD+VG/u
gbNz5xer/DTGX9RBBJBwgXRVPFrvLD2YvaQ19kPnzJLmB6QY/G5xDWfMuzF0Z5Wg
q3ns/wWdjACO5hzxUjudUbTqIi5e4rOMQMeTl+HtZENWt/mM4OSbkZuU/h+lOEWA
5iuxq6n2Yii4+8c7Bfe0zNv/y7I5/+EKeaRIuuEEyN84HD8ievGLgQ5sVwzl5gvB
p1T6c2wCJZJa+95ngZEmSNIJVR5JrnQA6pkcFHaYzzdeQKKyPCIF+2WrIXgL9N9m
vBjzsltQbfgUX0VXvXK9G+PBP2oEfzX0yKoSLvGB8g3V1QYnsTrRfscW8r3Yn0Gz
9Q5+alnuI0H9rb/iTWsZkItr4kbdOFU/6hO5D/9AYw18AEvheKA8ADq8L5JDcY04
Oy4q3TqazGbUk2ZAIaVo4PXJI4dRQvnDqyp7DAs2U8llI8Lo6eKVJAxjuP+pklgJ
Y6WncP8dwaWFN+HfhM93eRDMNP5E4nAKkk5Z+vJwUUngJJ4LJ2qHUkxvt5eWYeqx
WsE8csgLPkfRei/bzlcxcKl69BP7hNwMVDOIpSAPzfko270Fqlu7MVoAZxQG4IFX
VaqloGjzgxEvkOO6WGgl556OqV3wZu1W/om28c7K9J8hgwoEXVVEy6QSOdFpWWck
8Q2WFdU8A36b1x/cYhVncfZ87Khbso+r2CvkTPWJl8DER5B/EB24CX4GDtczIDyf
eiLYm9Gs1MRQytZdQ7/Epziztk9lWkupdsZCsAXi3wpN9MisfiXh1r7CMzD9OGya
TCyJj+p6ZqNTsEz29z6SmSmsdtMo8KUuJsMVcEm5TgRaKrWkEDM2yj/rTLviOcn+
6B8ANV+FKNrXmeGV8BzVVXQVoMxY12LJmc5UXeLuso17GKHZ4KcrQvongmnHYxBR
YzSnwG0kPs2eb10EEpxCt/gVuvq/ENoWnVonqFfkFzAv5fBDu/NWmxE/LCQ8sAVs
Tu2uRhLAkvCkKOQJv3sBUv+r2lxlxMlxV119Ewm7uwlFhRRjKkDIOUTn3RHi8lG6
1WP9guvxxwxudX/fJcMpgNvgY3Eh59wvbmD4W2dvPabF2eURmlc2+FujcqCQE/C9
WUlM4Qad/Ur7K/VHqOZS6rMmL08KnX/M8Lf2PeSbO62IuHs4FrnF+M+JfaaBpdbT
r1hUvJkR/T/xjZSNpK5gox72oBYMMOtQEiVE7M1+6a4qJcbUwMq66bszWHmJCp2z
7AztJ1Gb6POgOE+UiVsmMJKkjk4zHybAto2IA8hC8WUa6d2tK4BoaKOirj86Emss
rPSZwTDfzQ/Xr3Sjr56HehgijwXbriJYWLqNJkSSITDZU7pVWj10dfXIHDG7LngD
grSL02a0LuFx2t60+XaavnI8y4pFjdDwWcL4ejj10GltuFP/dmHC8HtaxF6+9FLT
vzikG1APTNogBOSEDw7OpOEBFPyPsqtWUs8TN3lYazyOmMR1Kf4fJMpOi8SzU7oU
MZAD1cAopptu/D/Oqz6+BZC3iCiwgOqwwDfoCDC5k6DtbgcXYkyO1C8hW629x5mY
GssMNxngpQsrxkmYHQszatEEkZUGUTksXRSKnc217GDYh33+bwwDjYWcVVe1TWyf
KCb8h4Oivzsb9yzW6ZK7J79cOXQEdt0PfdGo7xjpR937dXsfYKrQIXuD2O92PJFT
blqHyHy7DkabnImRMS963NPuI317lYcDPEJTu6Hi8Zr5ZYg69eMfue1in16KOtEs
ilRKhia7T+MpcSA3BPYLihLw/s4XwILLLmHhGjQ7fb19b36brREjR+IBhamyYRXG
SrlhWI6Gqe+2//Wd7JiTT0QAQz8C36mhUSGZmAxGfo9KOvsMqLYM9wWLvpUq3o5I
qNMzDhetLtNs/5Zdrepo4h2VXp/Br/vYc4c7HRythXDBdsVFGfsq9UivY155ODiC
5SaNfsg/hIux0QMZcC7UF/nc3ixRlEgJYeUVNMJ0G7jfWWkOZw8rSBWIxGYfgPEy
YWwTbnipuK8pcRsnSRm5tCaXCqQ/pVAMtzS6WmAVw80FmNsdvVVMSVV08hge+vW7
lX9IypNqSHflbSfSPx0cY0s3q+TLUMCcB561oTq+8GqNeOyD0y+wFNaTt0yF16GY
3rmO4+OKWj7+f/78fBVFmU7Ihoc8BrjzqLYVgyCILX/dX94SVlzlFPycJAokoZOS
bGZLWumPtkfDZyNqOrkCBhKBzBh/ZRJBEahaMtihB9AbuTMEB3rcIPi4N0b+Ltv+
tlDKosFaourps0DiaYj+2jwww2T3BqbDWeRZ8hm02m8vqOKX0Z4Xv4XdaN256Ife
B05UznmHmUbHSXEWvg4brwO5o4mO4gkFTR9EHo1EeMHkvDKRUoMrGPz4OEBkGymL
hga2AMEMnq01HAsVJG5MUU97lrAmnwl36hfWcegsx4sM+N6OWZfsl3whzd2JYoY8
BazuPNY6VSknUuDB2JD6t/w9s8hG4T4i6Xo3t0KqRuflZbK3/54DMlUQ8poWyKQf
siBo/mCvwgaCNW1cHPMbSxoAsQqtxL/TOmSVUIecewOuIgXat2II8BRDQrHmPbj2
hnKMrS6aCXWKG3hEcK36X8KaBhTFAPajWaHpriN6HYq0Kb92pgCerRLlvle5j143
cQ5QoBed460QUBjoN8Le/YsI91/795w7/UFTOf20nrMgbSYqX9ITbM/LXEnM2wHb
HozCrXoFmysRDJaUKZgIMrSjPiUTIPhNQcd3lCriP2rSq8CGaMZIUM1ZGDdci+kp
be5HGZ69TkIoellwRmzZii9ZzgzWZckz3RD6tRv3s08bfUjUeJxEorNsUBMv7fpN
r7eppWlMGa6505t+9XeRg2lGFKjbtxPE5vebiOw/OnSgPikdGHubMstGuZ8WGt42
R5pcFMULNf0r6K0RTPfwkePUwTKHFtEqxtPc0HJfbdkIjDOLbrHUQIzYeO9HXP+I
g03Egeo1lQQXxdjTFHSl65/ohYB/C6T8eoURtAy+mpZOJOZSS7Sn9S2ha1UvOmsk
v4eaNPoWuD7AXjJDlp3xJFPAPmzaQwcXBxFBY5lJ4trigWQyv3CUxZF1VpdXmORm
ei/HH1q6ugeBZAMllHmLRt2FP5jpK2TnpvmED3aoHKOO9QoWvAghpSnNg6IFJ2y0
Nq0qz9TkRw0FrQ/QbWx+HxQ/VXaulvpK4ZK9VjZmRP3ZIH9B+saCKq4gCu1B50x3
bdfVjdZr2+WL+hcqlYysMS3Sa2qOYBGhpRKrebeK/9aUHKdu7Uq7f/qxIUa2Dx0L
u2AOLeAWtcO/nDhkkJol7zirTPLwOL8pZmjIFvlmv/O0wRD27R2Vk8lyudxUBz40
wtCaEUKr5sycBQRJXkEh0nBEAYfwcoKmvKDO3/7CYog9iuq/kApZBfAGXM0Vc3KC
1QTj0nkf2lcLxaqJU4j6Qo/3J0XOAAyQnKQkv+6VwxWNnMLFG1KFg9Kmp9oEDQwU
w6q9RmR7p7GAqhkGnYb6YcfFCNlBrylTyXvLqla1m5JRXvMAnfsa212dwvLSw1ZI
ivXJz5lwBca80luufYnftxvkJpqOTfWpqjdz8tBRvVYu6M7+uq0RHcfIrJnQmNKB
99Nf60w+4Ec/PxAhV5FWJbB4FS/L2uatTEALKVmwAcb042J+r/Rb+fQDbob9QEsc
loAYhZLqY7t5+N0K2AxI7P2tYDvyRHhf/KUrONoxYwFimWJ7WdAfi3lDABEj8u57
+Flt/2rXQFzzxfL3jPp+vPqT/8hqtW20bZg8CjZdwUDZb9eAIeyK031HIg0s+Y++
+80JneeHfAmbJSZjkVdFqs0+NeIVSlTzEGKGraaOAXfck+aHHyNrLCdQ3VacU+rb
LcXZJbSf05eWzJQxzv/Wb5Q+Gc495bMMBvrETDGzXViwLkL2inZ7C/oO3W7/NJTV
jPWOxq4cGKG/YXPLv2Wy8zUjUdc2vO7bi9giTaGV9CCsXAe0mhsS9rDF4Fw1OcrX
Q6joL2GRPo6PeX2AnoFv5l0wNkKPfJUg1Imo0L2e2tu/NTdJprYhMc391VfWllW/
Qs+Wv1IRCCergbgIgDUieSCMv23A73WWC7rAGdL27bXYn8aMjdy/wNcPgcbUFvxD
glOQjbTTCfGaXOUbdrJ83km8iGMdBEVyY6cg/rfTvudEn7SOWPDgLn9tUri3sgTL
+DiKyin+Lr9SqY+GIJ2YZPPceVHtbweGcP/76DkUfHkEyPXQqdXenjqiFgzQkxEU
x4BZL/pWdQyKVstVHsKUocPyvhmr+O9C4VkB2/uBPxj9+weM8bRFsHR3+A9iHL64
uFnycfAQSCbwGaIXxfFSW1ofCbaxzOi/yB/RwHZPHsjXMNrEVo6Eoth22J5bJQ9h
MKcGB6Lh+gWlMr4ObpTd+5ekCVXypg4PZ2kqwHC4h/P2A6oAp7jwE57K3MyOpTx9
y60dNpyqojQu0zPSHA2BxOE+7KmETqxWlrNwu5A0hXQQiZlxu1D4I5exO0/b+pOn
MCMp3vG0vpRIFilXNgeoCxPpXHetFw11rNotxCXdJtUAZaodecTBY6FVnXTy6eKY
+AbBcYvALvOaQDbC/IdAEac2MBfRWHQy96WCs9SeKe2Ta8ebvrBkaY/xKDf/aklp
2IWBupZPL6zQ92KXUpE6zV7fu6p6FMYycmsGFE/l3a2sZwgVb8M05szK2lYJ58BU
hR/D01KJPz9r0o4w8Tkm7diFC+bpA7OBWzQctptJli3OWl5Imvb9R7jJevsjBHx9
SKRcobi/kToy4VWfmeB+jBuwT4Wgyj73uWHs/g+KNbAlbA46WyfXNuUGZW5p0svz
l+r267KtatvcN7WjuwMfhCUFvty26RXelcHjNx+uCMLhX4xdZgOHnea4p1UPOMH+
68yvVm47+y/e+d7tV4wfzPXJjmi6dzwUrMD+O9jfXR2N4Pb1EPTyQET9QpP9nfpR
LuCaNEfwEqvbnexAfPaMSC7VubSywUSxF6eoQTnD7GCqgSvqZZfGmUfMJkpnlZdx
MGH/DgHBxgE0f/AufXrzf7eA2Tj3Y8Z6hsTntOB1HPJ/Y7nwzLxnhkEJmoIu3V8f
WjzxsS2rwMMywB9eCU9uk1NuDTLH2Q5UKnAHrzhtMNy06g6NQmCpvUFI8a1HTodr
6rqHk/lj7nRGNGwN5BT9gE3y9TJyRtlL1KUwBUcG10YJ1XwH4pJq3+45OPYh7PbZ
f2m6CTkD79DKy5Y3ou9K5RFili4WMfuwEz4uMvR0h/RPs6QgyJyhQSSF3sF9MWdD
NnMtE6oA9cg6CsM2/Z/MqvmQ0QRhkzrAncwMVf5I+ne60BECasMsbrsAHeA3eDjr
ekQxo43eoChVVlVvZLn47LjXxAnDw7GNvqXoDS4RCmxETLLKmZDNjiBWHEAtOqOo
482c7JV4TLkn783CxhEmelEJcBfGgrlFy8hoAH4Gmb2AKnXx9rRMoV/z26gpngVq
Hx2arNb58n1or7xMkvAqSkCrHFsy8DMbmRqMlLIeRLje62QEFQeLzbMCRud37LTx
azeGCwHjD+dpNNEJo9v4P9nxgeyYNkf4SyTnkcqSEp+Bsxg62ZsqMPCY7OxTzNP7
IluADzriaIzGcALm0nkNHvbELtb5F4D7bxpSpXNvVYWRX6GACDxBoGyOklWXoUE7
Zx+24W51mdanaynbmKs816x+T+s1GD6Yum06xVgkd9l8MZdxErtHOAZKlwX0dhn3
Nvbc+BmpI2DOQ0f91EO2EeyjQNe1SkiZ2esZmO6x0B4IyKsRgT/PLya2Qn64f5xK
oAyvg+OmnOFnCyvezBcWm7dY9/Tf8fY2fOIqITbJwv2oXOWF0ticAWBINBf6Awkq
kbVVBHAzy0ASacw/i/6Ury7cISmf1kP6tnqsllQF/jQC78/xcBspNnuyiDFNm2F8
MPUGi7KekEdCmif/F0tU3/UVkrNuOs3fNODiTvPauO1t3IX7ObLGefBEuugWmLgs
oVymkYsNT4TItkRapeuverPt4C3IfW5AFEz1L+nUuFarNVDuSEN59wnEg8TBjiga
OEysztFuV0NLMJAPAR1aPMRQYkVnxA8OPTf23flzmPFk+KSA7fI5c4FS+JpzfZRb
ubFO/MouZ8KeXrJKboYaerAH/txyOCDK0KfxQ8HOauRGoXqbeHJx7PFQHOQWXJ1X
zqh25GHI3mPrKqZ9ohbIL36hSdg2d498mtznaRqIdDKwVhUIch1KnQm97YN768Hl
ifFLLznxCoJbLV608CRz9e8z1gfnldnEaDlvsIPSt0YUW9xiLI7BCCn6U2wqvJFb
ekxNwJGYPgQmWRKIF4Vj45k+boLJN/R+nRD5pCJ8a2w8FIMtn+aiH0TQfk9BVcvm
W9ilG6hnrsK3h58ivGjxs9EOHFPBRRgmm+h9XoqPVS220BVcDkgAyNZXN7eBin97
O2sAUZz9aGU+MrsmpGOX9pcpu0Wv+ytM76rn/qxu5OcZqxs1wDGI57MtEO/gcpvM
s3bEcF71Fh6v4k7fnrtCoem+k3WVWVnET04ZKlKNxcPyPrCg7ss5N/ZHdDZuxMjM
PENqLR94as9GY6QPartbKvdcySdfsrZMrpvUl65Whw7DkFPLILt2YmYQZE5R8bpE
BENeKxnr34FsuqQ3I08Mp4ijRs7XvkO4kJVN8JPa7d3NwgowmQ0RkhwjvbkYiNcG
J0KiypFXVIB/9lUkOQy0lQuJdEoIgqBWwdFdeFrkCWbOnzE6MxhFA9y3cUJf200f
J+jj1APLej6tSDxPTtrJVi48gGXL9sfOCzDUkSmANTZwotNDaffdPwgYriHtZI1E
K7T5ilqf2m43+wLkXbn3KYm32SVBkf+1mgPuuITsafNmiUgnP7DDkuAj5Kd9X+qp
uhYKuywwy9pOe9gr4cVgGp6FV0XYNRzc3LcwfM2TyG0fxJ4mo6Za6AXbEno8szvq
c4ADmB3NL/4uHjnR+dXyXVc/dTpMe1SQTd2MO6n9vHgd6RBvKh8xMuk219/y4XxQ
ZvUEXWf9GS6CgV9i0PT5lNc1Z6lWQSA5qWK+/NQAKYo7nOyFWjdq2WShp5yYbhau
ivJFtBuswfV52SpAaJXyfEdp6NYlharnZALd+t+RWtAzcaJSz9PTekIoFo4BClGH
nm/pYd7/+/wL8q392ILbStJqvK24ovNkFvz7RPacK43MXtruB+GCGuqho41jPbSN
uBWPHJRDqpDQDWsjdMhmcYo7nmvI6pGGjbBySro5IG4R80/8NlzTx5cyp0ASueMY
4viO/cOd3dzn0zFY5/RUxF1o+1Rq74Tb71YTiBtiJUmxDf/sUXuP9V/1b7T9C4Ta
O2pK4iLu9O8ruhXTps8E0hmzSzcFyfcIh1hkoEe4a77+3zCfi0PH//G+yXAMYtBm
VVEt1JO6TnmoqisdIuI1EFkR0tzyfGzNOylyE1nY+YD10hD5TSQLrLWvBVfSxitB
c9NskPpYKbqdR2epWCEV0KgKeR4gGT9fdouatW9uYQyfMkrlOs7oUoE1xw8ev6GC
KV6YAZh2jcl0U9+DAlzYw7cpvAFsrMYVt8E/+6gt7Gzd0vVde5RLdfDYKZTQkIyr
r2eVTURYOCmkGxUXIEiFhraCti5O20oJKKo/M+4pob8SOOXh9WjmsiAv9TMguIaz
I7wAaspUEid3jQRith5WpqURYuR5LlLEYIukB9IxOeSTRP7rxEzO/UqDSaGa0QBM
b97EoeQyfXFLJKuXrfYciIubvpxrXViHaiCM0T1zUoHyNi7wr+gBLXP14/g4VdhC
duWfPC2dA6mQwl8f154qSfNXboK09HbfjAMum/yDWInAZ4HNcRNGREBFaZfWFjKW
GEcCuhhVZn71l4o2yTHQtC0SZ5ckBPx8Hre2Bkaa8WfjEOMQSXoMcskvyiAWMqla
yAppK16UiSKqM6bsTvwEaJz5l0EFZlJjbHx38tjCBjoWpc7yGxUjqLlE+ddyBk24
jWMNonrSgdTuURE8pJTCt2l+OL4Xqh8bkpZ+loKJA4HP6GM9PomTp7gu1Eyq94AV
y5b2DuLMlWaZkyqq6Z9wPX9oAFJSAXFaAbAm1cP6G0ULaj5GgqyYGbpIEkzf+bOO
X02MQNyH6eJiV7ENcDSeKqOwHe9hWkbgO9P7+9iaz9vxMsXBEcBqn0iJg9HFqjWL
ihMZxxSQ9otLdOdjDF5FCIi413EjqPhOvNHr7zYtOo4RpD5Qv/cJfCW5GGGdUp4y
V1hSMvTeFRLrPko1RMb2zZWTOJ9XkIJUaWkkxo35ruJ8hX75qMJ03MMIS/+l4eXZ
hH5TJk3/XjiFhW2OXJIlHr5sExhMULxVOM+f9YZLN+K7N6gy20R7uyhdrKE6E302
8dVv75VsP5ro+qZ/bTINw9F9/drKhChyJRnurWNyZB4gctfKlFAKCudBkYb7h7Ao
dhhJHVcIl4Qh9SqBw0fmwPh2nqiXOztAA4huJyCYB0Hj7dPkU0mr3sypUMdjd30w
hkZCS/qdw6CEnEUwfrulZP2Y5Yx9N4GpGCQcmU8GGSbX54j+lUpmb+VyIOKSc56A
Sv7W1BZ9epx3z6WJkTBq0EkqWTe8W//GROMT4gQ3wViMxFrGzk7CabX975fXGGhV
HdtYrKNXjLwPblc9zjFRDoKigJ85fjep/kpP2HXBvSOLYZ+GvBD6uQ5zP6s8Excs
/7jdHOTBEa0VMVAo9brHyZ9UQ8xlA/wvy6hNmYEUFCEaDzIs03fy4s8d19NU3cis
YeSvCB53A3fLJd/lTA8jVmlZZ4uiJUK6dyIpokxjJobnh0E5H3b06nj4NZ2Miqs/
jBULxcl2j8i+eysZaS1IBkM1msWwk1vJN3h1AavFm8qS0wdY8wAHoL/hxJw7jVfY
5A9k7kC5syolJiIWe9ooGJWctezBJOFf/0Gyz+bb533LMtYkEhKS+Kpk1UpXU5e7
JUFZVLkCIlN0iLpISJjizI94j0SrTEhwuqsGg2gqZ8TKMnxwQrBxIbZv30p7geB/
QjKLkQVdwCm+2feAj8PQ7Tu72LGuMqZ1VN10+MHKPcxwep6G6x0ps9ccs8fujRwM
qmNdNrgfwHMLIYI8khvgY6B/v2f1k4zeCfzzRgZ6B6g7f6yx5JDFEOJn8/VupGFd
5y1rqizj3zaLNUQHFJrmlj/WoF8xObT0r6yib0DxOa0xTkBWXbKoFyi31CpbYQ+/
x/jl6WUa8dum6TZrpAvTalI8eMlObwWoHHHkZ3aqfucdeOf2WweW+gAjPwoXi+4e
UgL1Ook47Ol09iDiFUHaZw7NqExZintGD4KLqD4cXWeldZQwCqQsVjZtPu9yxXqy
woKEFKc3LORwuAcFe76KXS/Nz/2JClNMqQXopH1rz3baRte7MddyOGgu4oh8QuOz
kInSdi+LjNJgwTK7FGDXT92PuXKY9F8s2o/Hika1Pqt5LwGWv+KJDt5KwEGC0InZ
ClLrOs5TDVkzDpWx6uCiU81b5+v1bOCd4gdZiLpUZTAPr/bO/aZpOtA2THS3VOl/
ZGZhWXCIJtiRfZgAw4wXnSn178aTNLdR2BHYWILhKPAvvVuCqbZhdFL/1xjKlobt
PS4bNZVigfg39DaeYFCMOdIDBRe54aWDbtqYBwDavo07HLRX6ycSAEY927Iakjfe
RWisx2a7bg0omBEJ1APtPJUiIC9RNJDVGJBki9oMDJG0r53I5SMUPhhGhCL6zVs1
VteRzKIr9eSMotP7DcwEehLr+LJplvLdaU+F3u9sMBYd3sWT1SrWImizJj8kLfKX
amZ0hPd5oSPYe0dlhjAn9KLZw8fHRWNbd0WsLSUrkqYstE+cI8OaliQ94ddxtz9j
IatgPJDD1P9AGpIZUwN5hldmLEZrMOfmBou8R3+cPgo+yTxC8SBBsqih9HD3eG6X
x/T8aZIU9vd3Ytz3udUmF3MWKs10cp5PRowxvpySSFMuAdvUW0LY37PTRcHfS1L0
/QwmQKj4siZS0NCbeC3dY4FlxZt9unZ/ql/R2ajbpjbpT0vejXK8I7232znhVe5e
U+5ZvD+rA8cxiC8TEUGlNZyiSEYgB8YMFnULaS2dDc5FmiyNzP4b0K9qWUZSMHHJ
K1CyVnIjMM8aSDyeWF4Eu6Fa9IZpziP56azB/pkr7dWQ94Owf2xTeVMwwe5fmiY7
K/eODjFfeb4PgKaEPYqrXS1RS9BXvtkT9hMr9fB4dIIKVH6FBoPI/NjhsJ3XNdvo
Yql53czf/4Zx6aZzhsISalfb4OP8YRM6iK27Z1DNr+0BX+44orI0s0AQDX+/tmQG
0p9XT/oWE/yaMu7h0+4Vl4VmHZLWfRYCLAN60fo2zescHTOSDwhzaIkACOI6Yxyy
ZXf80L4fuE4n6d9BLLdz7NCveYdB+Z+yGF+UruhEiGE9VwWI7CWmo4C38GmXShzX
kZK2Vl8AQ2Q0huiSposwP4rLK7rxg9LfGnCIw+qbIR1tSHMzePeWKmTaNaR7XWCj
wqmEiX1VQN5Yx4Vl2DNKhg47V7vqhco4FTY6R3Lcfr1B0j+vAqEjGk4aKlRI6bMb
PsUB3BaWldOwyYF+k40WpWZ8xFyeLjQI3A9v3r24Ayp7IRu7mISXijOMVBDbDK8t
rhE8k5YO7ugCtbcQFhRMh6IHsdPgXq3ckjpqHAs15586oHDTueCpLt3QK1mLY/mS
r0hpZs+RQrZd9Rn5WQtzogEU0lbXHgCaL4ljyiCaS32Pns2k/1mbPG5I5vFYJr6P
x1ETyEUOudxyWSJ6Kz1mpE91tnGj7Gnt5zLs8AIQSzXwLsIpZZgiUr4Mqeh+tUpK
E1KlAzl+oigqlAzbTxcp0w==
`pragma protect end_protected
