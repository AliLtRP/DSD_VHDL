// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:25 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Y5Xh0rnOxPy71WjAhcAVGJf0k6DOBL6EgKZ7q1f0ilT28SM+ATPeRILV+31yLbtt
5EBT99QIGmM32UUwwlVrPB6b8I+UmBPew2pv9SSk0ns/byYzcpccLeaq05ILDaZ5
24laqTpmgv+Y8b3rEiZyaRiSnXaRnPW6BttAolNul9A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9776)
YiuLiiNy+MNvB/QHEAf7wqFwvmL47DPi7c1QXYJiIvuvtB5AEEp+zM5/G6osOjYu
Ic+Oh8Z9COwJAtmgDS7vs0EaEqJPK+nCo9woIsD0G2b7Xaz9X1fHs6bNkGNfGsNM
D4gvlTYoMuTGHY1PiRqiiCTxeIubYEf+7102DH2m2voDqD8tPq7BhmlIFkOfFar/
GbmzWfHj9HyKe3iCYILYESSkDV/nmCHGYrL1tqYqWS49Y64Dt/mcyJdBIbMlo4zC
vtr53eW7huWUgbhfri3IYsVWO8NDfSvjxxDkRU00T8tFvm8+f+7WeTSc9maZILSf
GrHIk/3Q287iA66oMhYGR8KAe3hB9WUpiTp3fITqT6Vm6MXTgMeBl0p6tCXx/Tfu
kSvITv8tGVFHSJN4lF3jExHt2h023O9CW/4ukWYJEL50/t3+YtSZi1T/BgS0hx/V
B4Dhx7JeP+IS6rGAYuPcWrlF/Qsn7sszsNAm0HJ5eU/VRxruuu7psK8zjByVzTZK
TW9ecib1iwPeaTO6UWv19tBO+Xv3QkqoGkEuKMyFJ5mgi/aAdePdSoLj1Xn5Pqtx
+YlCYiFNQ6uW0yWG2D+tFS8dhktKe0LC3XABuAo+g28Iu6gouAMRYqm1JYeyWpKP
tFCx3CRJvic95dutCDmV5xJniieo7SmYloivr6lfKbPh25p+ttOQkoV9KE//U5O9
8ymU1skzmikDMdk4uMNYLVvWIwHdMCuif/oPAE2kgiCnFj7S+v7H5yv4tDJFh+vy
BTeG19IKFaadkL0nK3MKxtTQ+qHvLJpyGP+P/yZNGQBFUN8pqf/VYUkH7VAGv85D
lxmupzTRdFPTaRLxboZGN3sNkqulGENKJWHfEfSLa/ahbtaCxBE4sZNUyMWOrt9G
ztq/K3Xi++141RnJcvHyY7B4lag+JZMxiHFiHcShmeKsmw8rAsEpne1JwRAlIp/r
uZzsXQrFDrVJGMHT0wqFklm96CaKsMm3yq8vm0L49NrI9ihMghXKgGxnCTrGhm4d
N5a2KjqpX+E7Oenw0VkoNbru78235yxMA3ensEUtJQ6xSSGLCAPHCIeMoursJdQ4
5XTTdPc3xF7iQfT/8N+bap1rgqSGasGzb/l3ImIRxBhYaJ4S7K2ALdiX+FWMLnci
Si+4775aqfxjgYLYFFhhJgmHJgTJx6K6iqc4KdRdwgjU3zceDqclKmOCvq+CBRGk
lx3QuIPILiC0EBkXgCAOd/lccap1VHwmDOkFWKJJJAZdfDuLwj0/MM113gp/PWtU
H0fyxlUSoOfwxvBV3grexFDTK113uuQdShcl7d3C93CpweF/LVJFodJedVkCpVs8
ozWTtbq7VszIYrth1qMGGr4LS93mlb7oKsHaqGuHHfZFWCYe2J0ZU1L7AVwqvG44
UQF0mBSf2E+UBBOtGXklg1Kw5XnHpiAOJ+kFR8QuUsBHM9Uo2t2nWOyQcXlt76FT
t5NtvyVqFUoy01DzDB3cBMHpPpey6l/zDJGGL2NOWEYG/tfTci+UFhYY17hWZqg0
kiAhU03OX/rNIvXAqZncIb6afCxlsdedaaHFzH6Mx96sLkLHwEBogta1HpqwAUhL
rG2vPHBuM0zxgo7CHQaB9mspkbJXRrmkdL5XfZ82YJv1hVmiRzeMIBknsJgyzZS+
Gq4RpeinDbACMXCXsbZaxX5sODTey3Efwr4BU/K4AONVCHv4g4cWQ78QrWlvK7su
IjPQLivRHigmY7MtkAQj2KiNesBB5CivCh1j/SsE6QTXJUiM9eQtvQAknrhLVvSb
oOojtJrsf86MPKf6QKMCRKPITEMoNbTUYWtkBJo+HT1CLqELUgOTPH7kov0a+hHp
j0+mjLQp9ZY9dN3royllb15EeYz1evFf+CNaJelp8dGvkCNBlKUhdyp6HaUDn2k+
jW71MmynNOnb22xlmjzg9NOFNPcWaq6NghgptEWRdOXsHY7TDJWcz1U3JQMK9M6P
XY61cGFOoTxxgsFXe73YEG4K2saYCz1r4w8pcIkLfbe39kTD4I3GEnjBTBvZbBbd
hOq0v2TsRXRPL+rk9m4Qc0+EuoOsP0zImOaQHC83kxtFbTaoxLTZ/FWTMZa/gAKS
uJiBXbytjHHYtclY9ggJ9W5fzsMWJ80dz+BHZZVQwTa+tXzu3X/2bvFyOZ3kyrEG
2Zp3WtYaUcUTLPl2ErqNRk/gzWc6xfmW/kLss1bSA86e/OE5YS+WxNr/hV3ZThoU
QZsMfw22SRnZsuXkZnEgf1Y8s5QNvBGMbPg+/FTvJEl2cJqyfM48fwOPi8sR1GwO
MLoir3hA1tFEQZg+73Rf/xSWeb540ibWpyOC3a+CnIx4wyC6cZG+LPjc8HZWDbMr
5F57jjc3kISONCHbzTWW41sCLpjiYHr1MpnVcSCQoAkRPJflfFy+4DZeymzM5fqv
YoYLaFKOdbgi1FH8NFToJ/sM51WwlxGbe15XGcPxYBEFcDYi1mu61v2464GK6xrX
kSM0BeW+Fi/w67Gmz7Z++KGSHQHDSX7vwsK1oQM6i3R7+QfRPlm+VYHOVkuTRDac
w3z64V08NiAGii/i/6TPMZ8Hma2KVwF8Vu/nV8U10aZkb4+NYbnodP/WBtYEjbPc
PpjF2CwWgq77p1LTkZcRyxUURZmWb5oFD/GsqkCawAz+2UiSzdI38FnDYO+ob70t
O5lEvsbcLZCHIeMeQSDty/T9d7pGdc+YgLNJLVuvVBTC0sVoFrYScZI/9j/RFX8W
cS++hTbfCZFcw+M+i0uVo77xtHhFeFnuYr9kK9+ff3Pz7Qx961xB5nNQt+BqFpgV
Tel1cvExxOsjaxn9B+MADtb9cyoXO7BEe8mEGzSWRZ1d8voBnzY7klJMmW2zdnpR
CaXVOZ5YwAABZP50WQIDxNCrAuJgxRyJyf9cQXlcW6+xumDnbbjTFZ04+gkgu61b
3Fli+sW2Dj5ecR67RpACwsSwESsjGUcp1W2k5XyMJh02sqSsxvd7BQ63+HHhTpYA
EkdEMvFA0NTysH7RY4uzsEiD4iFErUptcYDkxrYN4wbP9txK8MwFhfwwS4tbH7LA
9BadJou4CWm9b8Ahrx8DzKfzK70RCeI1TOBtwkn3Pp6KeeEVj6SONwVI2OkB7BEr
6W1AHTGIca2qTYXw3bhtU0y/nWZY59uBnJs+ui6nVO83ZSvSozox0GCX38+nqdpL
u7xtCYMAwBFp5evFTMqoNR7hSfr0TA+cDD8yUqiSHVp45oXSbskgh6A7amB7M6Z1
Hpxt8rnRN3/rdM/eZnBTr4QVWWIvoBJvJqivZ2A+JuSryalpHxetsO4xPpbj1iPA
xlpq0H5iKXMMs04DHkDgLFfQuqNyA9odr+RbCq0Gq3s7f1AtQvt7C3WhwZVf2HlG
RI4TM71enjYM1rzYg8R/U8UW3SdTQwW4kg59IQwcwvMVpZ0p9lveX3I5GuRnrooh
04Zhvm+Pjy65QaXwEtovY9o8KzNRvqcg+RI4rR3fSGEGqw5Tzn0tCzFrkHcZGJk8
ZG45fx6DGpEQmrMuxumGjYZM3EGsM+NHeQ29DR2mBypRo8rebzo15IIHu6h2ziX0
YY0CPRLt+gqWghiGpxZQKrIV52RJEetJNRC4CykMKflcEoKlpDdXtCdUZLuodCDE
T09DhbJEAsSCeC1jTfFPKbmqghm7n1yC/W3UKgaSne2WDT+b95VY1VT+J3GHecju
HZ6EgcmdgafDUQqcghoaStCmhfgCd2g2oIfWkJeNJ9Gv+NJ/Cz+ew5zmp6qKvu2k
vdCIUMtmZWmHbJW33vq24gS9BQP/XJVjmvJHBYBCK5Qurkam4LDmQUGLX+V2LdbK
/mf8qhv29rWPmfcydDzcdvhKR9CV+L/pxPwOT5ekzq/Uood54FR3Q4XJ4x2FPLm8
m7Wrk8DRqx0UaATpq9l8xsr6FPLuVWCtXGqCgghfChRcWAwYtpjKW91TCDR65CFi
RHGsr4T4TNuEQi7LUEqqGu2gmEVzP2D/YHyrLQ54htUb6t8yXzTPpdAra/UE2DWf
PRhrNvNr/uHxHaokmhz8jkQeF6yU1Y+D1t0Dh9nWlidO6qhw0uJQhAomDMWE4xmV
rt6Kt1zbIRLgdCNyMFWeoOB2QpAAUDQuICs4O+pNGTVJKP49aIqIw4BXQR/ndriG
wU+LjbYb4rBEJBD9BZuKlCtJc1nqJ1nkJo0LURdc8afsdBJ7orzIJ56MNoNxnTRs
94je+/Sqc/JYElUE9HIfhD9x0B78oXeCeUEdIk+rddHvgjn2HjVksA+JxJlB/JW7
juOOkkTDLi8ppBQl8EuhovOBRr6NbA8px8MhnO/K0Ljo4OF7u2gBzuutKL1+OrSQ
8t33FTebWgnFsi5csQMn6SaEQkm5wnQpzve7dsZtAuveV9+usom6I5j9AHYNLeQ0
d030ZaptTuULRELT87gndlbcm34c4SwqFlLxIs1q3IQWF4bm/AbBxyR3CMTu/RHp
n8hz2KcTWmMAOG24nbecMNEskPEpLO7LXWERZpxPGZdmHG87+zqhWSIUuzCi1La/
yRsrV2XTH4eqcYt/sY8EKXCvOptWVD+A3xKB1KiBlBjdu5CoMjC4wgYItrmVfM/l
8zChuhVArpu3o5JKrktRxYKP7NlWmVd4CG97xBHIIDN2Sr6nXBxwRoSTC43uFG6y
cuzm9nGw7t5kekN2GMcTbmxSbBDJ/pAv8YZfkjehRSzDYYasORaduTabqZ3UexeC
c1Pv4aAp21hhEd7lFJvFk8tEaf0TyjJDYx0NCmBASRolF/Jdr1BqwQy4nk+A8ts0
vSYrQmElAjRQACS3P2NwKSV0/qqt07VtuvsIhmWVKjAg6JqhSCvNay2I+X2BI5no
3ndaoMY75tyOBiLiRdSFNq8Cf/ccF4uuUM76piP+AJC6zzmB/+y8W8gQzTQcAuiB
NNwbg51rz4DUz9KlP6xZMMRV+alEswH9rDJLPEpgogZdfKmZOKu1rJdQuT4fQz/+
Lr9cR36EVKYX1xQY4fE/z+K7pTopv3pqT268FTcvmUoxRNfVLWnvukbB6ZNn0e+q
e1ZYyiC4K2Agw3myYyofBTSdjvBygBMVTM5Fz5/67LY7lWDskHeq5SuJoxs8wkI7
eAYPgydPKWXM2+3QH92BUqe7qjhxRXRi9oEYSb3Fl4eLx5OS0pbaJI+qxM4ym/rS
swm0FF4i2d3xB2VQs3nOYR+KdHOjLeQGwpy/Q5MRNaed2RhUFBxtjjCJr4jw3hot
ePL4xBE3n0qa4AgkKWzOJ0XkqenzSLFebj9+9MLF9joB36rLNLANWZkZgpvtOy1h
jrO/3RIgoNQku8TZDFFL95dKz1sN8AkShv0ym1qDyPWegjY6LCdzWfTC0VAuw4cJ
eIySuHMzhgvJL7Z9JEoMDqy5SSgco+/A3XIdBOeSLNAORzY/l2wCCWYTuPqwjEji
Hu8F1GmAmVBpbaTG8ljNJL//fkrwH83fMrExA98RESPfs99FrfMGJwxNlG9iBynS
IUhdccbPhpUlUdh3n4EP8L26skLe9jJS58rLn9b8np2MKXXfYaOWkQZYqmi4Vnad
snpNB0B7XVUnjaZPkKpwNjjIlOsQXl0uaCPNfZjCRg05GoXVy+gJLQiY0+j70/wv
6zgdjuhC2oFzG/Ljygj99oIpRwrZY0tDewpcN/nmF9jAEO8Yhqp6tylnPM9gmSa+
zOzGqtOCl+z7j3oKLbMEYzyR6GWOEiPfNCKNflAT9+BBxaAgBLyT4nxItsXPfpX5
LDJTNvy6WYJ8RuJRphnI86VozZnngB0JcTKR4GYkHfnSeSPNFyFw9lDuJYhsDGrj
YuB01W55Ti2/3yHm2kCAFBy0tHYQwut1y4eiJNseGB/dJJ/AM6UCquvJkt6qiN/x
byvx72qzfomfEZbAHlSFnYtF30S/7VBJzYsOlNT6j3nIdlvOPtMhMfG2Z0h317BX
KP5mRzRr3B6TAYWhHE8phwaBxJSQgKUCc0X+VYYAaJLDPNzYamGVhkbeP3D3kDMA
CWGBF19e0ZCRhFQo3kAbZvpW6wktozDuOPn/p+B0YxS2VYZgOzQE5VtexxZkg25G
3/igJalVlsnHsN1Rb8rP0lQw2i92/9PKciD1rkNgz716M2cpMYSikLDbR9cdAREJ
d1Qjv9/JEK62IcxXxkaF3bp7pwx3gYuL/uZ20J4eOPpfr//Sxd976hzlIK9j1eqa
eRpCgh0JDfTFfbkQQS3RBnJnl2cw3VinflCPnSPJCgUxhBSFx+hAkGihKgTfU5WB
IN0HPvZVqJo576VrhoYyIfFGOZanbKmpfpxsiP0ul7B4c9bYu5SYDlfwgphGPE36
EUCak0Dmu3OPWv+4isahibjBl7mZKS6Kn7PohrC2K0kmvAIftO6MANCDfvGdICzb
MTYUEeSyCjooRXK1/xsj+PpcvtIE4RWComd6vcmP74cp7dT2NC3mK46oKMKPM8Bs
IlD6TlpaX8POGVbdXLKSsTbNB3li3v+ehRis/xl9hw20RB35ZRZ4Q60HBFobka3y
32/VbePu54LPH+VznETEbPmL6dW5lqAPpv4qx+c07W5d7/YF1Ywyyr4kWTACqS2d
ZmMAwAbvOuB17t4YbhTBrw6yL0FRIHvfMZFznk2hNRjjAA7X7b0nwa8W0vJ+dO1g
K6Iedl8rJ226nP6Sp7Sg+zw4WFT3G9IzHva6Mu26iunIYFrHegPL5oz79Z8Sd/OP
RDWjT/gv0karqgWtg8aZTi3u9WwjsPqK5GClO9EbfFBLumKaF2FVSH299lrITrsT
1uiAQwDic0VYqumM3Xlv3xjIYN2HVgDYX2TO97kCNJcsDuouy+oP46fGkhDPo37m
f4IOzMKsj3wRh2nJ3cyHo1I15xLNM3WVD6W7unTzsTgqiEA2U7gxJnuTwSMzY321
cmTnoT73SvCEIKPIALT9/rdViYP6azigHwgfQHGz/fKdxgyS2uw8L6cGLK+jTo39
3UM/4NBug4rMrIY2z3wdsvAHcWzBRMTWfI3nFR3+So4vSj0Vi6UBW70PW9FN8+PB
hBfekGSyPkBvnOD7v4AqUzWl6xbfvqHKD6dYq5tqt4a2hHU7lb5zfUvR/Z74uVZP
EG66LR+IA3aj6A4VFstdKgbtFkH/GbUBxYJkVD+vjfHywoFtvRtns/4O0t2G3P4H
2OAq48OoGgz/sXEMu9TQii7aTu8J2ke8qAj8m4/i+s8D92aod7olQIMqliv/CLl4
w7GAPzUq2/S86KUOYHeFbVlsjFLID69Kr85fmh4TRn+Phss4NL2Q1D2NGcaH6zV/
kZ+3/QyC0L1g3pwMvX4SbslmcocbQo6uWmoEvhi/sEshX5xORya7TPPOQXexwB8V
w3wdbx3h3oWD03ENIVQsckvjeP3NqqwGb6gLa52eTG3i8zlcKNo1DsylMapiacC6
VxTx3mV6zlJiKzjh7Vh96B1qVyrrqr06XootJuoKC3JTsUxcvoWxhj4RqRYJX7Xe
UZwumoXntLiER/35bH6h3LXp3pKuve+prWDgNCX+sZ75ZkDOTFT5Cn7gmEpK9TFb
Rd6/8Rq3cRYTmNPaafd3uMOrofdSlEFLS0XH3B1V4C9W8+hLEkXlBFhTIB2lpHUF
gS6rfOkCw5vifGuxqQCGlmJEEH2iUGf5UTIiS37lXb/ISeYcvJ96bx7mfjg1Bd7n
NG+lRyzfNjJldWuMCTH6+x0B3pCEf79zoXSVNuEacdTackTHBSJxplD7EbIkjNDy
oNIkJKOQI/+Y/WvyFFQkcPQmnPdg1gOyjGa9olmOrf9MZZijsCNpEqvE3GLSMRNK
yD1wnt+oJASyV7nZPGzqsmbiXcPfefJcV2pnIIEwAh2F6qPkkGzv9+lHIkS4cbG7
gg9Y9hjNu3fAhDny38POnh/l1f/Ovzs9bVBT+SMc63WB9dupz3FYMS6jTXVqdb6r
gd+TT+nBIWWR8hJ/amO/3v5lM8B3cZA8aXd6tKXalUt2CEbEJZ3LxBtVVuGFnHD1
ZdrD1gwV5keQLPHMmvkqT6ILFTvwH9S6I/6RYHZF8gn9GQdaCsq1XXSlhf+EIqRg
6nxkNfF7R8jEMUy8Bxz4xNjoyDao649z0sl6lPOSnihj0QJSxAJ6oOrcyTko5sdO
kb5Kar5UstWTaygGN5cXC3JQJzXOnjBCyosCqtE5lucU45FRuZsqvthpw0HqfY7d
CaRrX1+GM0Dwq49ADf/jkmSkT9eX76VPvakFj6Y0MFlZ+nFTgWrT3XHCOF4f1pru
7s5nk4n/q0BTNKAH4WyVsON7jNGQqHLzc7e7QnS8Nop/CzWNi+HCr4HzXBemu0Et
LGZQ81XmKUsS/r4+Q3Z6Jwf/gippna+rsrbR9fxen/zbwANLmp21gy4nEF2z6+qH
KGR+R9a5j3oe1Cvqto+RXH2hJcPnKZdZ7F+BxX4wXj4RocfKWllzZ9j5Ddy9uba4
R9812ziRDCWEu+mI0gm+3mv4Cho2J/9R6AmGY4KRCNTSqiaEONYSBcWULt6xVMRV
U8x4VFIYkS/V3DYzPyq7RJKkAYFuma8AApMQd4v6M8+ZINkoF1+mFur1RJlLu3Jx
Nv54SL+5OcOeIAl0HOZ7lVY49zW6TEMPE0OzSjPk9yYWTsLjaSEN9tDMwDBDQscF
eBqt8VvRzkEiVQj1geacVxbErscNRxFzC1rr/jr6dPbU0MQi63CsmjjEzJU//aEf
kUtVeTJsly8WfDU58ez94y6Sp7ROQWTlw2m6keibrby54ARnbZK3Jovm+SlQli7J
WvA/9MF3eIU9wMduXKnQsCKl3cjPhOz6Cu0u/Baihr+9dJS/QRW7m9HmJKnUL8D2
xuergI24VNjxqy+zm6U1Ima/pcE1gPZZgq7Hpc3JHoIpyArIvFmGolfvxwXX58QS
N7yWWR7sytRvgDtghylWMUAC59O8UXm22KjcKbUwXCkgkKTg4IqYdC249G+tokN3
PXfKyaxTxNBLcPA8Fx+0NCiBSagtiyMScSmS3lzSXPk6jzpg1R2OuPwAPti3XIzl
HPsI0mpr/WaF29A56ycTv6KTZZnzgD0IJY51LYgdvogOf2mHpXDUzABrAlRbcXK+
L1XefQTV6Mglnm0jY4YBboig6HCCK8g+WZ4mMil96LuLEZqlDJPRjJW/vWYQ0nX1
GuN3twr4ZKCAmA3oAj5raApCkgmsPjgX/XzGk31ZJc5giYcxKIO4WSnWDmBleLfG
WC70IUjXSju1WUOPXWZ1CcLZd4WQMrasuR90FA+/BZGqkveR+mcu637MGQizO2nb
19WmQ5o02wZCuoqMVFxgs4dO9X+4AEBTJnZqucvlMH66aYrk+k6TNd0zPsYPjMFX
PaOltY3fWp7KclY0Qkk3WRKdeJU1+0c7HSLL+u4Ro+DdrjYSRnbGot3mUlmwjQLy
EHL7ipMa1lDPFTL84bcNQ6Ceha3Sn6tYVS8v41bU0hfL+B+nF74KRZgBfPMrd6Nz
ZVlCoSTiZRptcgejhuZ/f706lqtuLmAlsEV5kLVuFD6SeN23oWlKzkctmJG7KYaT
mJS0e5ZCF6hfugSaTq8J/SEn5pfAz8pfsmSsobY9PIf9iTULJ+IVyJ+KesKmT6Yo
wH0jzH6v+9YAI6X0NQcwfAvR/CIaAmvAuIrtW/i4PLwXCX4ctbaXROLZ9ueDAuar
QiwzUtNUUTznTTOdND9J1A4yftsvXyBxIF0kJRBJ0obPjmgTEJ9MgcECgUi0d/GD
RcJapZiwJB1xLHTtNjpj6W0qKHGfMNv6U0edYvQO4h9r+OnOu5s8minAsUIgHK7y
z7puDjzLrr2zb4ca5oJIgxaCz66K7Ayw3AJ038YFbevKVrxBbAivZdkaQblJ5Pi3
hF+ePoCPIEEdM8tT4gWSSLBalSopGfloe0fiQfKJ7jZv3Fe/QBUa/xuAemvxKFL8
bVvXZ1Ir9MvTqP1G/nDWJBZhXLMUPn1QNoEcWt1MM9+EGoZEa8faBWUq+klSavDb
lPX3L0r21G8qFfhxLWToc0rDwy5WvdCH4z5angeLlXmTkOzKl1L4xgdfkEHFPTf8
V0ndShxclr2KyGcMdErGPlwIkq77ZReIwmwRo4TaQdFbEr1rGcflFJBIhBUNk3JE
ionkBMKCWCvsKjwW/FZAJSWfyQF8sxetMfFZXxz4S+s+LF0Cg9ukSou2246KZP/R
srTbPq5M01QQqUZu929RcPIYF+kqG/LSMRQ5vbchdca7bp32F6+pT7PLqAnSbGpR
l8jBv4mna10JK+Ei10R0rjCm1M7XzT0Ub0V90yYmzetBW2d50DkVieMqWWl898kR
GVeQuhdob+gFilpd9d/959dDvLd0jTZCttnyu6SsI4WZhbwSJLvIcVsmiJ39HqLE
BRqabpuPAqYx+W4SLmlhAZ9SdhU0j1yW4BqF/6MNGLMlGtU6zwrUN0+d8e6AaYDl
XvIYfJ90p57Dy2IIKGI8DKWYhaXu+aE9+dILcY9UQG16IfIoE00yY5ypRmYt86r+
T4ND1au5X9ftn2RC8CfQJZ5tz4cHEVx244CInifGh7tAwoYlUGISemexYBxN5Efm
m4tebkgSsqm8T/5weHzfCZd8JpOQjbZNljcMWGYbn5wluTjaDsm+4hKlLlHE3jQc
JG8xsbmEzdY8mu+8M4EJeBDhzTKpLhiglyt37X/H+f1oirQnEesP/SNid7FkWL2q
UzIE/3drusFkxacB5F8E1znLtTNTFwbwF6n5NsvL1WvuEbIOhS+gTLr0o1nPw0Pm
FkNEgzwwYh4lX45UA9+8QNRa4P77UajIuqLdxSLts4pVGuJrC0f0rhs6UIGSNEfK
pDxyZe7xIaaoMpDtEelJnmzjHJXpoHRp6nNWQEnqNt7djHcslUDt9cMrq2FDf1Iu
I+DqfitQNn96cFiL2EtEiiMeak/E9E1JoIgjYshjxecb31t7cqbT+LHsx29yuTRx
Woyfj0mR91EhWWKHf9tnSXKjAss667Wv2LIveUx2cFvVLK0M8u1Jx3GfenvQwM/a
IhXN5bCH8r0YU1Xe0sR+8UxFuZq0mS4Pk9gtfVmlHUNBnhzns3ifFYpwBMldwR/w
GSgJAY4J4Ob/dxfps0up8/fAoZCqcgPQR4ewy8TGjxjVqi3QxoSUxUVcpQNELQ3a
u3bdnCShdGB/WtD68CmpZjFi983PQzrQXZNDlTtpE5vpri/xei4x1hM1lMk071qb
F4iP+rsYKHIq3NXMpWDkvwsCJfnDZX/1JcGZDT8Aqg/QYcbqOgMshmqa7T+eF9LY
A4zLSMi51u4Ucs+ixvbLHDNlld4Ln3GBkbj1ii5iqdUGSn7hej5K721yRBOPe85h
itri7CnlVVbRbqGSfCEmNknZ1v/jq81i3hWyMjoQKeHv5Z58mY9RDNdCfNER9mKh
kFrpT8rL3jbhH6sc64jo3wMLGBsRx5PKryQ0KePytEz8gK+szSqIBmmJV53FbLvG
79O0PTL1M8mpitJvquJQlie5aXGtJgspYsCYJUPK0kbkJ6b364gYDBYwQxNcW2i1
F3FqwvnNn7cReX7W/4T6sLJ1hTZubDMrEB9mZzkj/N3HqU2cJ5Wefevav/CDy3br
LB6u/GGJ0EPwgP2nt1+PCdUzSf6B6CSLZ2bCckiA3JYl6Znz+BWE7p82LuoD+OzA
9iw+joK+LeTO+7b4f5Dl3Gfu5gIFyJUL6v2ReSNgqjrJr/Cbi4VcNu0hNU1q79vT
WuMrZCTIT+RZc7na3C/aC1rxVM+0pm5yIWPXzAXWdBBE9lxetUPVRM8fRdl7dq27
em4nHPy7nKkT1BUaGWOGEp0zMh1MXcqs8ZScEH/1OtXziZQ2wLT26ob4d6ntB/KE
B3TFQZp9eWH01wEUjDUntSil5NX8KrHd5vSTLjMO3WBXICFJyaGoHU5XoImUBogj
ucAkM7FREFJwwt8W3iLOu8I1Mpbdy64xzjdlqzSRQLikCJEa6KmPgj43TJg/uk/R
V/vu+fcEVEmMrWhLkO0AnQWTkHHmCfq1XERqyY0MGWUdWdlJbgvtyl7oLKTl5eyQ
F4TjfMvDzrCBjaZAeTZPM9KyANM8A5nLXzm+GxTlyKo8+ymHuATGlJbXhN3cI9A3
WnPGu44m8XwMXxB7W0fguDjKL0+lG29diGDSerYTD83FbQPw1lDKTup1xOozghB4
TcKRmtQ7vlImHb7+R3nMJwxwTs56iQrrJzwO7Gajh4FomE3txddvIxqluwlO05qu
wZ3Q1OOHtI/LVHUbWQr7HuTWSf2dUVTnhxQKF/0WA1m4ny1c+7L2dMdRENM+atHY
mcLjR8GlL4WQEMGoRByzJ4SVu2RraCKaCUNQcqa3ruafxV3zJJ++XA2rq1D0bN66
fkBpD8d3EFr1LVixkjB7GsW3ArsxmU9/2M1Avh6v+ytMbJsw90K+6gQW0OQvFh2a
WYqoWnK7eoao24sai+ogRrHlyW95D7cX5H5JFbGLwoJcJp8nzAhCQUbMl4ix4GBP
GFFmAe5Q7SxkttIIYE9zKDYz6ILQT0GHCFNYRcBt69VWv7P99MBu5ulzIWb1rLbk
ejONVeEMiHsiPKdiMevFv/abmp4hebr0QjA7J+AahCSTWjz7gnxvsUdCP2IyFgNo
KpFacwtqiPMqYAeWd6eP8v8c8Krndo5Yi8WF4/5AD7XidXyEiKDIevbHKwAYQt5e
EJARvYywWzKshsN3O5L4aEY922apA+UVZCAvBRA/cAPFanZGdhmPuGWRTWuRaqkK
vbtHtAY43/Wev0j89MdNGBwSwxOsujfSJi2A4mjjtA8FKG/eUVyg6HUZu+s4o6nU
un6WZgG/KfG6cUL0kfJTj8tMXhC3Xu0GoLWKHWnm2pDMDUuIKT0be8d7nBKHXsAt
24VIvlonqn9frFxHjJEOk9W77W+0M9t23FI9fofhBQ9/kowpXPaNecif3B1c0qci
YYiuy1fsq48aWbh4tu0Pdf7kVkdVNrETi0sMJeFUAC7jTWPJV3lgs2nt+bD01Vw7
3ggLwbrY4ADWOve03Z9NLRlJcHYA0oYqUPrtQMsqjJw=
`pragma protect end_protected
