// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FxdMPPpO58wzoetQoPZlekBHvxDB5E+k5URiAoSx9mv1M6QyqAXS1dj4drSwnJQG
ZhUwv8dzg4tAG9DAa4eXdTLbnV2i0iQsnic0jy/L332SABHI66zC46tAzJ4G7vig
gxwAFG1Qh7AFdC4USgfQQReYQUuBOfD9DtWFbfFHTKI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 23088)
Hy4E3B2EG6zE8H9vRlPyQsraFmHlM1AzftQAFgJIKZtHwndltW16oy1Y8FpcCZBY
TpRJxkVxCNSgUONcZdSB+v5+4zR8evCexWEoj98wfzwfiBH72Er8V2GOWmfQzl6Y
oAdnk/cQRQEUaysu7SJqC5SVL0C7H0aRT4FuujCvcmIHLqoP3xNm5x8485qmqTgU
TmwZ0itlHIDafRmXmG/1Ze42W0hv3I99sVI0isVwZOG7YWFmnMIkfsUBeLTT2Fj5
FEsA3234snDppWFrny8AkWJ4S1kHB1FtgTUoWb23e94G/cqoQyQerWkv8Vvx5mvG
rG9S5l9X7tjtbVzrbmIeU1dP0pohoe/mdKM55G+qObNlp3q42e586up2G/R690YT
OXnDypryailtlgxLYyQ/8NfQPtFt2yDCraZAMQDrpOstbZbgqWTK0jQD2/kVir8d
Onqg7UcYDmJnEOVxnfTMgnLHlwShUi4I0DN469TDVnitdRtqVD5e5ZWRKqgpwvu2
d4QyXu3HsDrd6SkS38LGstku7akaFevEWTrZArOzA9Zda++9XfV8x+tca6YGP/SL
8awJnv1a+kaYGSSX+rUUElBxqYxiOZ04FbM+CzEX7M4icuxUELgyRTZyE3N5egU+
tZDgTJD4wiKbMOeJmqelxyQlSVQfbKD5hFYZfLrao6Xnycsxuf4SyhF+Vf7wRUQz
QzqZotZcBYpPPmsDmhFz76fvM2cVdTPtxqR3dyCKkrOC9lSW40u6MTsgRS6l1W2s
UqzM17nvUA2+JF3S9dA5OStpU5uneHOO2/nIdrU8WNuG2zTsaW5vVjr+A1x6KiI4
hZMqRByPgxbCqeSOntldA1+LIizZCdmNYy2DBvnYA4b8i70dHHq+uiiMbyOtEk+8
VmgAz13Zk3p05Uffh8Ljs2uw3qh/huDmjwGgh8JEzFOtM6P5go9/PdkzJBrweNKi
PyK1IAUAymlgQ6vWBeaZqPgCxebf5qayXrxckGx8fFrd1gpOYg20DBLLyMOkBVR7
w5xBXowDeFJWgXbQzP0PSLssw55XO66jAduuHUvux60xETU014vOjOj6Zx/8e3X4
A4STSq26gywLcx+AUqxZj/IEd2aL0Qv3s8CYVq1yIrVrE2aB7u4Gsdc/DFSGCno2
lHbeitCtlt4ze5+2MAyTI9Pjt6Q6K4jpHPQw1U8rD9jdFhH/M4uO8GSbUc4xVgIG
lVxLrigURbMOTQC2EVNKtLZIYc2FPDGG2Rc/EV3NE70Yj5mZI0DRiu+4s7GHpXCG
GPOd6ew5JToz97nKZvBmjaB/yJ2ozCWqnBbwtSVSdEw8rer3Qe45GiKhpaoyk4/o
J3+YhNYDoDKwrIh3h2uwAoR/D3UNAV9L1SdYrOCXpOGdA2nW0Z3lDjpGrcOwciQH
bI7qXO6epPxToXHjCOPdpQO4co6U9rpYvumygBwTU8GiMmzmx5w7buVcQg3ez3YS
cZ5kq6vuD/f8EsXcRywWuSQkim1nwe+JfrQeZKH7f2WNpuxtkxRS09ouGVr/wqVY
sRCSyhrrDjD37fojlgGV0V+Bsb0flYECyI/G2GVIiBExNme/ezZresRXQM8Jlv34
sQ8UkeH/jyY9fpJRGgVurlnprrdAemc/swdAIqzM85bJs1sq6VI8zWuJRNdf1fPA
BcN5AzSnRjJUhdwY2CiKVqGqCG0nY1biL0SmY/2PFq3qg8myiKAszobZ0PgdHbcZ
UN+HCsu5IacqNA8YvrpAP46HHywXj7KGKLFu0+lewoR4bJZwyLidxPd5eZgp+/ia
VQ1b3EBePakk738qKsuLbtjDVx21BdYHYEBURYC7R/3ZGa3GrXF/Ps8DWhA8kZcp
Qk4tnIRkwSJxe0Cgi9kxaYT83MNRVYhY1kSM5aYcOLBJpNrTy0ra5pityusO93xh
m9SwdLMKOQE9mZAp09tCU4yOrMwFJKhrsONM949vUwSrjXoehJV0tCfWNYzmTqp9
sBSVt1xSoKZvGwiNas+17MUJrTF2z5Z5aocC001cX45wWvqF92UKTS79o/YvNuqr
fJ+iAQzWW/G56QrKIuyhtx2NcYF+x4TB0prvH/n5KSVD+GZnsACLSdbz51vO9p1F
dlDMb01dQfhU9gEhoyshTUhCLPnDqQfysMVvphJv6DIr9JomNvVUGz7j0CLW/oa/
LWP46fP2jajgivNA0oJpwtdQUy9+9QKD/RnSUt8iQHniuFn75C+fVrTl0Ostu6z9
KgxWfrm326jRAkmlDsU/bVE29dhCruXKl0UmNJle2/W6nT1Qcd47inVeVzUoEiYi
a1Czj5KPoC7/a3etSzFr5wUh6/xI94/EUqPtCI84thyuOxIr+e4cj4RcpNY4/9aF
UoEc+AfNY4l8SS7FxHG+APHVSYaiDY679/ophOhBtXwQLHagksSPdidrFwXIM8AF
mxCWB3HMu9jD4cGUojBWEtzFAmCcxRuo9t8TmY3THCpgg/jl9TXSQR0lFBuCsoID
szh8JugH7aJno6deawDjk6zTf6rTU8lYUyZ352Dh+/tWs1SlxNOypK9VLwrl1ND9
uLMPc03agh3+ylaQiv7ZZO28qImZ2nY3yAATRtxH9fW+5WgR7YHN3SJ9l3BKasRN
cBjeVu5EjyYiEkNt8FERqCtYA00Byru7EGul+tl7saAdBqWMiYGZR0/Ai/D+zI/J
Ojp0SINoFBkA3sy/NACm0Ojoo5zWZIyoUllL7h/ZVa2b1cWNwfYRCHurQqD6pQXA
MYg/BzMiCoL5HMmPogaVrY0IhCdnKTuAUv2ltTN2CooioXFRDj6e/KVm1GHmOZml
X/CdE99B9YH6PaGfVHEJX/HxNINZtue2OSMklepNOtw7MWlGx3w8HGOkwVE+QLA8
9lO29BwbzE5LLV+vJe1LYUo980TIb7y8BRl42jLZGgvy13JCDNFGjO737mqgGBhW
cHDBhfYW0tSLVpniaKe12T+NGjs2TZT+1Qtf+D9NsqDr0YxAsWsRGaXd5nWAkosV
HBTphcZomlYgF4a7w+3Zk3cLI9i+jZifsYNKe7XltUd5JUsYE5KNn7F1KN/jJrbz
B2jM9P2O1Ci8cKKRQKVxAp1hgHDKkC1oFTdLQL7HLdNwPVTJoQO9Ec3qFn4QcQMJ
iAG8lnuwah4rPqVE/Rh5/jlsW7/TTec1WOGbe096wRAA+u4sxnLcnEEWYx0lI12p
grcrfi0eIPONWVoNsmkbj+IithGtCoF54UfThv7Kcb5M4tKSUMdpGQCjYhp2NjJi
kG3jsJgilwYghWyDDBbPFn3NhV0R37SkNypmw113IMaorJRPX5FTxY6HBzAODGgI
iroIkpQEFPUfYuKKa2BAWr/yRDza9PrAMPkzZ6xytXG7jCNWr1yDajc2kTBXhLr4
v0VqCFEdzjBkR1uOzN/SpyiYk/XLDX4ZdGuRRJ/1r6mqaVUxbZUwONH5ijFERU0Y
KJKy4s/6JZmVy0Mid5CsrKdn/P1ioAQf/2TBGXfPdnlOiM7lNneKaqAbAbOaLJPn
NVxPtziLBX4RoiYY4eoR3qLb51x2jo+ylNh4vlbCcYLDXq02FAwRLnGJHBrSMvzg
+KqC9iba2ey3vKlClYiyOhh5Z6BCcFXscTtj2Dnl+pQCZ5veNipxZYZ5wlD41EF6
uIMW3d2BkqwWAlQKDV+ymOLXknMW3tDHgKY+2ryOyGkJdQB+5mXGYczaMngo/7aA
dNr2lbCqCHgX4/VSAPNurEQ9ItkZxmUdh1S3jJG0SMeVgs6zrpstD6K/hR/Vtc4I
gh0TY+MiXY35X6MN2a/vhbK+dK1ggz+1az2pSzj13bga3ygpIQLSrZ8pQxchT4GY
X1sSOXNaQTgdFjKnFiMa3aWiz4WxuSUh5Vc7UfNxs3jlbQ/qh+WtjZBi2v/NXnWG
1/6XQDhx+Vjtw7wTD9ABDor3t5uTisW1ip050frwOuw63hlzl1rROhirAF3cT3zx
RcNzrUEXTGlpLy+I4+YLUurxbH8S8rrHbMCCEPe7VG79KC6IIVMvkSEgUtv3aAHi
IXHgTUIy1E2hO2/9KrFuh/G8RSpP92++CgAT5j39xtDN//0KAjnR3Oi9/KQgEh2R
581i3DQxD9qYh15M0S32q8XR8mg4NohNYjG386aEiynhMjOgQRwnxWHKMzqyPKvz
RWpLEJfSrdR8IXiS0N6qhO+f3t4xnzj/ElryR+Da5rcsdAgLEtXmXem7XYnM8BAz
Ko3psQWwj4dNvOeKuJj1AmwA0CPNx6IjhWaA25TNYePKk7uJvuxZYYHlPDaWa8wy
W5quFfErjZ+GkqQ9IjgzXfT3c22Fd1guqRjWr2+uWdQl1RTrCE/uKdWNS9+zOJLO
C/Nh/r4KSou23i7BcHBPjO1ZhkvrLYYvll/YQn+Kv6NivDx7fN35Pk+PSvdbzjGr
fKyCcR0qzXYr1iz/UQOSDQ/c4voL6UNZA634ySZUq41jnf4xnkaudmsym/SkRhiO
QBVu76rjVbLij62rrPkEa5DVR8mQJxUAY8cfSg3OLZiWVht0eR3lL9tl1ADIDOk9
fHEBl5OiIQMngFDYsyIk1xytmkwbeT1ZfSzn78zGEB0Y8lMpPClThJv/zar3VEyC
5Muy5bS/YjPXRD5wxMD9rn/9os/bQLh33nUgdZfE2fKVabM02DgRtVyIDIPR/6yB
qSlsjwe8riO5kdSr2+JbRj4IircIISYH07gQ9Karag6gaMoe8y08baF8xrp5j2X8
gXU/BxQ6Kb5Av9nRcBdzg1NdYuhyHt2fhXbiuCxe1H7xS55YBMPL7S6oE3YD/Pzw
l8Bmxk6Zmh+6b5rNfVey1m92/G+Kyz8G/fe41Hr/qrvMYQ8OE+9NUv1l/OPCWSKl
FaQxF6u5BrK8Lrk4LnXgJ1EUx6+zuwtZZtdeLjbetakf1aVbgsgoHN2J0eHl/DVY
DXDqQFFJc1x5IL3qmyIiNDvCzZ2ktVtzx6GJcm5RLttzr9F0lwpM1VVmDza45eeB
69j/MA308De1mjRk1rp+x0/VwUQp3UH+qs3StxbHVACYuSPxUgqkHQu+hoNOH/vl
5PubUUKm8WyNCXLG/TUSjoVM79OiNxcwBlldM3zlYIEUsngYJbb100uil7wnzPGm
V12Zqe9k9F7KUGguSa5aW9k0Jx/XeH340AN3oR8hibW0NMt9rt9mL8u4fh0WjMQH
zbeJgxrORwAT+96brf2kCGky+KoxBDHShN7N+z9ReR+JqVcUb50zU6AAJl6Qb0/R
8E0nB4vp9sBWO3kzd3SRzcAEOWMM6eQ58yYDIeAnsszRk4VA1HYq3k27aGZHOJdj
IuGeDqCPWYM2tHHvWW7rRSWXL7sFvlCQHX+xFLPgw1Zc+zVx95Y3ARcRfuVx135E
1cvrJ+8etU/TixySXy5jvMpZmwOSQUBcZIwrqC/SGH06/shTAzLexgLvbxp87QbM
fgKdeJPgYCiZmrEucYAhWs9ca49ijod4CmbsH9yZyZF+oF6d+ayWj8cggjNqIuuO
BorZkKXAHkKhXuP9RgNFWc95IiDfrHsT6SRBEd7rNr7dB/TMJClBUEvkD/aPkoIq
UJI4xi7ErZkcxzgG2nbcJvrkudBHW1NEpPwpuaAYDjt/OboaPRBYG949codfVuHM
TfLYGNDmGWgTJQH/dXSQXjmw+XH3aATrwvvYEMHfLXIJAiU98qTEUoH8ZqfoT41l
VZQ7RKobcRiYH1T+9YTOG3/5C1Bk57+7uNVCpJQYfwApBdRKObndVdS1/jfMHFFD
YvUPle5MrCDbv/3/qGJCKMkjmb3YMJTsAIyM+nGUrCRlSW3tv54iq+21mm4vERxY
TBbnKe02jJAOnfEi+zTzIsRUqJ6afgUyZwMLOoe874aQj1yTw2hf1vU2Ohnwfu/I
3zn40ak2Pes/OdQhhMAP5S5eiT/fnqNVpXmb8bJ89JHrgorBgVpsmy/Ax20letc5
TiF6IsHLE2wIctHXValxFBczVSehk7B4QQKYBNMnFXmiF/y3AbM4cs1UCFrUH8dg
vw2YL6M8TOOWmgODGQ31WynmY16mDbchEL+HsSmgh/E6S2EDqTCckxK60Eu39vDn
P5vKgQoHDkaoF09DOlspccaW+nmgemVxMpwya38mGbVrEo2Cq4oKR9zN27e5zxP7
YQU1dPWSUwVsODNy6jBONS18s8AYGBHCgMBH5lpP1F3PHrjGmV1Zd2eS1GfO0Aob
lEgHPg8bJ2/GN3BwTjxx7hW3kkdcRzfmdnKejujhv6CfafOU6msCpAU8RKFd7t42
B0L256gpyl3vzbLUNtq6A1AQPt7Faz89LAHcztTRPnIBU3P1nKDV2kfXtlNS8gRy
xTGg2SIMXbtBuriuZ8A9/qnQ2H/9clmeznBTkIxzsHAVty8h5Ml2DLXIC419AryP
5cZHvdnF2aqUDOsxgYo4Sj7by5ITogQGaMH1xdN6q6nE84CbZ6uWFaaZrf78+BE7
CS+XnBcy4WOx+QTDD4BdOLx8TK0tdRukZlv0z3uBzsOeAC5+X8t3Mx7mTgt3IQhI
3k7Qnm/mJMHnexbktv7zOI04m0Y3l3wRsEdoEj3u9kIDU97H5VVr23HeNy9QJkM9
erdYvmgPCqaCfC0h58cNJC5DCuSVzOAwOF9RJDA7hwSoXN57cipbXKKvRwMUfnrB
R1TAPetr0TwtDan6rNiRRci5QP0meFeP5MTUd3DxQBxFgFbiGf+8eE9xkG6GVdwC
7EAWXwVztjvLekvZ+FJnEgvOA5PLMPcSmW8eAlclteHf6n9PIxGkMOK8Z6gV0KHc
01UPFwCyk79P+g2cCJQkw9czEuezJJGV3bnTsnJek2OSbqlkpwohEQ3Zws6OXCxW
ihnGfB/7WxfeERpqn3Y0sNccA8CcmSd0B/Up9N2ZP5hNv0yQz598Cq2Vfgogzwd7
1b6TkXgRzeSFGK/UB4TlRCaEKGxAn3kudXk5P2XUTsP+kPS6uYH1gi0MHXK4bfb4
SeMZol75X185x33eHn5MVgQjc6GJonDHyI+DwG33u0DImSe6vYnZ5peqHEpofvA1
nHeV5laO1gRasw7ULx5g07JXQlJdyq3OIoxMIzEPwZRzosc+VJ2pb+ZW8VgyAzCz
NwIaAKEvurNo6NjJUSQSSHz+e9n4ARUrCNvFdIQgQ+Mpx8XcUpVrhHps/Qim3xe+
8QPM9osY49JHGZ+hR45mu1GKCOiogcWPlZwlDK0cF3hO84n9KikfNHr5maZ06aJ0
6XUlv8+VxveZ1oVLRNMIfqXsfsnEbAo4Jfz+RlAUf7Km25sVuM1Kx2+CZymylkya
iqZJaPBLPXhI0D3RM8kQ8ar8QjPLiyKjGW2X7gDQhk4zA+uYjRiKWYgayCBYNaol
whU8QVY26qukxz8F+t58XiHTfD6Ya/wYMhCV4LNtB39g1Pu5eCANDoXTr8cMh+zn
wtjOV2bVSD4Rv1IExqdwzWzyzIXgPz+cMDrYk2QBXOec2mY3BaTK24dhsZ9XrVnP
kObPhUod8e/DZNyLz8IhoAUQ0ZBrfgAto+3D4LL9t2DazGFQgQpQstsivD1olDpP
4cWLilVgF/5Y6dx4FK6HULyaFL/ytF1t1EgsLfzLlZ6zb3IoXrtnNurYAx6xXJuA
j0RNA2H0rOyt+ZQlEtEy4PdNcVF51MpS6WFO3yGpPGDOO3Qht24echw7RPa4tEEf
QLCRlp20SYSim2BexkDAkgeJnSM5eHRiUdnbuFo2Kepjz+q2kBLFgwHcgytTjfxb
mc7JaIFgLei0uQvRpQ2RmIooD3D6ZJ0apAN9J94RvhOsbN/nbbvMlXEWMAv1WXc/
d7k8WmIFkqVR2SRiT25T8vfCZvDWzJvqJwS4Cr0chdFuCIvXFSQD6Zwq9a5qztv4
e84rB/VKXe6iQCBMHCaiLHdhwzF8T3roBs0araEw6PeavO0nQcbFm+3WetS1YRMq
Uw0bnosXKokeKLu6d3wPYG24A02jZFNjTTydVU6M/T2qylSTGAtOxc4dStzCFDf6
cBUwSYNE8OnHva+AH3LVM+YTj6t059WFE3WyxRI+anpeWORrtGYvnTc3B05JQ7bM
q6fNKToqSCH/e8PK5IOgQWOM56jHvBwzZ6mFVPAWuNSuZFmFEYm0LRdGxn8v5Abz
jPAY2f0VxruYNJnjw6UBOD3RFSnDa2FaSuUe+ph6ZZl6facw0c8lePLjULuUj+HZ
Fm13T+UJs/MNeFli51HaMws+u92IKxuVdi0CIhEoT4S8r+ulMF0WX+xPThJ/yV9R
Mm6sLfvtcQCyi9NQhFuNIUjLJEhYJ9MOk9Z+S6Ph4cuSBU/X9Egv00ZXpsXiSbyC
4JwkSM0L6PZ1seO9kLHmK9zE8bD8t+BdIFG8kDFxeTQcQeeBYOV8rdk6NJ2Etr/E
qnN7eM4dlvjx3rUydAuGxK61SbibolHOFx2JEqcJBHRquN7X+x7EDqy4HzqhdvNP
Or7TIZkRTbGOvG1ZlhErhpJhx3+FBuwdqSNeZR6u0OXK08goB4T2fXF+FQnfboGX
A+fGjorLoC/aGbMb8Y4Ytv6GcLQMJsdpyjpRzd9ZAKpBbz2Xj7C/IhtgZkf+7PSO
/8SpAN3brR1WBzWudl7Q8otMDjvIuFk7wUB70DwSuDXUYbHJcPvKIQmwIzUcsGd6
A4m4ztj8RdbBCmdabNiw/49ORZqCNbSLQq6xoGLKftpJlPqyTkU4AT4Iv3Zxv9d3
hQfNpewC6JIhS4i2WF88R48SJfwsL+PAOsZS7KbgkaikYXga4XQO2hdUWbJR32er
lVGGdNhgFFoaTSRD8pV+SgaqYaQf2nZHkW9fYjaprnEPrynDICUZx6L4GRrQxMbY
GCaNzSleQ9SH1OOqaz9BxjY9ry3RxcCIRVEqX+CWIGLyK2Gb+mubWFbcmMXkDAad
17XI5skPutGZChrIok7+gWxRBQIU8oebdZkWY6Oz2qqfOM0KQEN/5x3AmCkf03xf
FLkydgP8Sg21ibBSh8mOw/v5lotgnWXRnGcDxQl8O/jIFGs9nIP7ofLO1MW8hB1L
8u8sIwd1SpMNYavOrORwjSHwOTKUwYBVqiky1V4BOGe4vd+l637xKiXvaQsI6mxU
L8KLqXQ6LDp+YrfKuTSFBGzHQgNlDtu8cisptvIz8b4PXtldKhDPNXqghkGnhahk
fkYt5p3nCNDcwX2GkHZlMEpKh/B9IfUTt1DeiZhNDKe+1ZH6UbnrgXg9qp9rl/jr
wZSzZyKiW2wINMpL5Q6ZRTFDbY0NEuDJQciRKKyTxh9uT5aCmuWlufkrOOPJg80z
5XX02EYYHu/PkKo6BeMY2aWabhKIbYj/JSFjcwgGM7KUxO75yll9pwPRi2G2xxHW
e8XympfU5IIG67cRFKWbZQqdA3lyP7yKTYwhvQv+3cj/Tt6H2cRgcftDUxVH9xmT
6mltr2H52PUowaYBMGINilSHXj7w/cVo7JtlpEzJ+mZKQ7QyKoER4B7C2/cnBDKE
469Olbn6sswO+FaiDvQ/bln/XpgyTMpJpNL7xp+nh16OBcQHZ2SqcnNPb/fcfhyB
CLM1vZM2tKoQdl1fieZiJPgSqDYS3w8pi26zOwlnYKYO1L5HatLQrTrAbDOqk4yC
usFJGEUsskapmPeeE1PFIMoPHi1P7d2GXXuiJk5eih5DXiW1yncDS+seBjUuyzO2
sNJcLOnp9M6su45dbssRzxFKH4rCbpCSNy9gj0zGj/tZ9NrRUw54yOhppH8TY9Nz
qJtC+s4wndCfbU59Qgw3QIZBVSzkFAve35VLg9spJ1XwFMHH3EOfQFPRrarxPbyn
TbU5bnEvtF1hTVuS3LQirLGFU60D0jw37F5G44SAAj+IAd5By29VQxKVbfCszdMo
vG7XA/0zZSRyG76FeRiGlea4HcFwiTrlUJhJun2WrpFGp0mZ9x+ikpNROKx44/y+
UdWV00WGuLqF2oy4SyEYmH2zB781zTC6Xn1XzwzLOYAKsTrii7n/lAybdluj8WYG
pCAT6tXrcLiRHDfxXJf4ADE864d0nReyzJYG6qi/b1DWwHsHywNZlC11UFiswWSt
VGuluAMZv43TsLy+kW0rYl0bfE/BM9ACYLt5EimMtWsJqivcI+OayjWfxmkURo3p
cOwwpbMfjQzdWf5xQkGPW0BYHmiK8vqN6reoDt7LmrMgeB9bM4l43FAv3QXU2RhH
xAmwYr9aglBxGldIPkWECGBT3JLd6K9JogQ0Dp+p0mD7/gL2a9C3vtyvZc65dhxX
TGW3BgVLoDQqLMxSxGw6Ta1eJsYL7v20z0O33cBFv2wJsnPFe40zB1vuxXWvzcoy
tFB7hb2cC4Aroe7FCPOLi6sXfzvbI/JIcY0xTARie2TJZumVTW9t7fWyHq/DJbwX
8cOBL+gktbupaFAeYWKFmZ7ZJFkl9H3Gr6zEfRXIv37K3/5waHa3x4YMq3VvXa9p
whKY0WHVc2KIxKpC0tCJr/aQHZ9RZ/xSzmhunaF+/n36Nz9JRncd2dqRlTsiW2Ve
TK9gWVJnObKvDYAOCmGblKa5F+S4h0BFzVbgU7xrgd3juiQWA9R6jq+0O1R2synD
zQzD+a6b6BsZFpB4YZcb3hm1dGRQlpiFTvsHTpJwO0LPi146Mr4AAb/sdwlu7oJf
Y4MYP7AgMaTxQjBmQ/BhhW6+jSTytzKuANfESiSAF/xB0bQKH/reEqBc7D+hN2A0
0q9AbfMOZRHM4RD/RyvWoAiIja9Ku4M9S0/doUH7NGjgiA2LB5HbZrBO9kvZ1uf3
oHifHUiMVoc8n85mo3UK+W+vWvuPcqXMwe8sFzuALKSJ5ysVKWA/yMXVN1541M8U
ZD+ckYQpo6DfrTgzE45iGFAtg+FN2LVu/tZ+rsMHEG7mKdP2CqCnVyB2awIuI8XC
dbmr9FK1mw4CZfNhFcqLLW4bmNkTbwgy5PiEkvng8D25UFk/6DAmBLRl6VNo11tJ
eq3A+bvhFynG2yjQvBByNML7mfs5YVf5dpuqoCkVWnD14vbOay2g9aMwl+6byGIK
OVK+pR3ujuuoTxoPWRSPJPYK2CO5WkT6d9OBehvXd+m6kY2Z8C3EX8oM0tH/o6oL
9dNyJloQX07AUbDyJwAj9D3x5Q6E1vMWgxGlWhBwrgmQsfBlPP2XTnl5tklxDSHO
EQdxLpI23t23RjsKtbZOrAItszZabfMFZOWL+wV/1gTAX54WI8mUjnqv1DbcjGCP
Q71gVSnvtkPHT+t7RPe7FWj/iaguB3txhGKz4MwktRl/lQJIqVoP3yeiq9qKK4uY
ZTtn8ZI4d/JWhIAVkFhlNkJL+yvCoyCZnksSwMrw1WLvgyue5RGBxsNETkoZPI4k
mY7nVgL6X3C59AmolVkNgsBTFbC4iHM9AI0TqSQHxW2J5uE2un3GXJ+GSb6mea+a
2KiPagI6vTsyjdCuKFAxuadntZv2OMOldJf5grQe0B3gWPQGjCVBznn4VbgudKmv
hdsJD6xUTiN7dcFibq/vcffY0wa0EQnhxUlprrq6um/QPMiXQhwB93PQnN/9mV4P
lNLpWuoA6IxoorI2jLTHbUcixm6huehP1ByoD9lUfZtn9QaK3uX+cJ9y1dm5y0Ml
9Hj0koLMRjaldKQSXzTZgtANjEuQE4TyWrlSivFZ3b/MjNfDgMTJfsmT9tpMLkx1
ZocOxSk4BiSa0qkwpEx//VpLcnr0qr7oOYr2b3nn6cpp1DOIN3RT3l8/BrrWzV0T
m4WRkOW/byz68b0GtW5AU4M4v68saZUNyRcLVSBCP1gHZD7YM8/x3d5f/MFBUmDd
bA5pouURhLtud0YisOnqI/FG1AzkHYLjE9z7hA/sY8vfRuQCTDSR44Yg7DEFRB2e
7cvV4I28yamxl/dMNQjfkKsuaoIMSA6EiqrTAreSgLDI/7E91z7i5f21Bs8AiwxW
QCJ4Rey1XM/xsRyJIXOS9sOuJpsp4DS7p0RVxAt2Y/TaS37lW9t+dJQSxOz2+rF9
tIwbDhj4sn1SKTZ4AxpNzyUbXiWLLfdHP6P/cLwKwVvZuxlY1tkUI8zczh0i/7cL
ETKFU6047tjYhRLXb1KtAVN7kRlL88HnCxtjeNKm5vAKi3MsSAF7G7wTcyP7N3ha
NT2HaxEXR7l40BHxVJ1eIUkvUBvbrAfgw4qY7sMz82e20YBBMdA5Ky4C70UXbJuz
UbsCFIaiNWfx0BBjEi/oKUQu8r+PMtW0irHwwAGPLYmqYFapUkmxmfpue91YUfup
9hCOZmcsTAbEIOoQC4UmBFt1bGxHIh41+LRNUS8WGjRCHIEVImrbYxTzCp7+wYai
10G8vMrg+31cw7kKTOkvh47BdeHqsZHBnveFvm+3eg9rZDsf7G9F9BGlRW2/lYIx
pBY7uS5+m1Hfot1vIsr5fp2qHHdpaZ7efz/Txg+qa8TFHzPG0RHi+JHVxmLpazgb
xTCmrsU85PmBkKSKuTErWRK2Cj3nXAbgbwGwBqck6X/Q5FW5SIEmDppsfjI+/hJP
zTxmZ7nVf+sjnbZWiGu8MbNaOYlv+taR4un5q4rNQ96An/xQeba1GxfyLG7hOlUT
9AKtQR4nGKg2VJE577bZKPFnphhUCkCMAHyqx6o/MERLHB1wRdjTFApMHtg0IrUV
bIACEtWGCCOfyuy91KLctgt/bT5nbAAHRBhYWSBA8oweTELBQGEZzXj5iGtvb328
QRm5yx+5l+0dPsOPhOqGpPmT/EjoW8R0dNvQp8yIDQe4JUiMqx+7L79ZnZGyX9z8
kWNyRQYiMD5xGPHpaWglk39bgqsAqcq2iSxe7t0IdfKw+vECgZ013XegeD4dF3TF
RY0PtJT2t38lUtJZ9Ii8E0k+HYvXFXNmFrmyRX17hZfajrfOFElygb2rVdOtEmoj
CgGdkFDvr7a5Fw4C3MA19HV+UsTaDIgg0Ux2PRXYefpqj9LQo8b3UZCnZHReT9Ic
K1/eQMFFMrfnU20NhjNsh/DkGTIw/BgS7ZGnFVlcgQHmvq/uTi//I7GZdYdGDVxO
fsqU97mEXcP5TZlf9H0ts/pqPbqRNUseElw1CFMqAdYEyFQBOD+UFkd57ThBPosD
/fh59as7jICDmjjlZymqpyELOjc382P0pXCZRyk5BDEqnzpYyIcYVeLMyMq5xq/L
7cPkYekVdnurlRSPzOLjARbesM1pO0UrXSKuqadgsx3eoNKeRuyfMxl6kO/JBqbT
hKOXIicgiidvEoy2WpMVg5T64yFyiUsztPaB62Ga/AzQN/3sZQSlvHvBzQSrQ2QB
K94PAheha6t/DVF92ZKlX6WxLjfA3ZOj83nMd+9smKeXEjsreA2o9dOqaVYmWIgy
ju6zgy6s2Xq1o8Jydyo19M+VF0dRY0fRG9rY8oPl4s1MbiLX4umL3RmxG5TP8a1a
O+O5uXKQsHrIpyZ+KKn7dk2pFn3bIBqyAhPeqZ9sHwzhaj0nA8lfAbSnp6e0U2Zs
TAVrtAZy+bxTtbJl25dCuEavK8EU8s1CSeaXeTWKqXlkM2XZWLtZo3J7tN/xgMNW
jngtBEPTC4SSJVdm7oJeaVPONOrlBZsfSBl0f8muV7tJDlpyDZodWBemWN+cGsnV
YweAVlkJk1gk5KghQVV6EBh8f8gntPblNkfcrisGoJ9OMtP/rz1bptl5NOIX2SUi
Gj8m54mrfOP3rc7NrIQs2omEzI5IP7TvAf/4NrKlgy5qyQD0SIzaIBcm17YZMNtL
HSG50PzR6lILS+T8ozJp3b95nW791+KBlP/6L56/S76WIJKFVGtbJ1UFJbVd3xdZ
wGsG+J0WeyCTpZJGLqM3z+RoqKZhWE1N5ZO9gCS2oFjNMNB1la7Fco71O3bljv0O
WY85It4rGZ9VqWj/ABrXZkJOxl3JMg9bs17SK10lX7UTqFXIgSbrD5y7a5PT/9c5
UYHjx5CLil01H5rYpJN3tsRLAXWglQzQZsHYbaTGOCl8ExHKQ/FbhknBs35zUhST
/SfKkuTYtTtVOAPBWkVADpJgxqf/8YWcWDJtDWc8oljr00KPIinaM5MJsTNDNROa
E+d/7B/KEs9KS2E/nOIiU6EiyuPh/aDRyJBYLOZ7rsycq6qTHYxtVy8YS89D8MmM
HD9UC/GO0ql7svobeNmHm72id+rpwTkCHVWLNo1etFywX9y4GQpc7AXWkCUJLEEk
WbN9E42G2nLnXrupR+H196OD5btpIz0+b6IuSg4nNNhhIum0A2uiREpOExPepuxi
OYuROx1PpLJpHwehF6dydThezkVnzoBq9nT552mHLxEFu4QoqqC+e6NhF4/wiGLN
Ostq/EbDyKlKpPG5UWhXvGzlg8UJ5C6MFXrGzaKr0tgEejDN2zkgSOnkLhfC1L49
qU5uvchHwBOM+8ltF41G9DrjCrTJnH9s1eyKDJjXn5yDUEC6mBjRBBLXub0PSNQ4
E7KNm4l2XZVmF9Ey0OmW3ElcJqq4NDSyJB3qIjvCoqYIp2rJgUnfwa/Rzu1tQb8o
uFEXYk7OdHTYFwppV7HBCS4VmwCOWbmOM0FabbXus8m/fzkGhhaOdRen94LTeyPn
CYfwSwcvQtUqn8PbCTh77dCuY5CXatCUD7zZF5jnfOvjwsGpWgQwl6ydrFY/AzKK
1W3s7jw3cQ6+tgdPgH16vcXoC10A5mMVAJO0SdOVVBWmttKkvePcH3JhwFzgN8kC
pVxmf1NbqLHY5zpIAnFlo3kQrm2LS1k1igss7ZHDlcMWnmMl+F97/6Y53qyMkmeq
OCsHFzcHREDpp5s9bV7r0yES+7MJpd/M6TEBxoyFqblPS8BNBQeaLcFnQTTHpu8f
7yenfL99de6ZHAvzgkMzEpHxevI9VqKTWo2RK8OSEjzZFfAg70zKm1BQ8+vFzmW4
nN4q0xexd7q7G6Cy02OSZ6jaS0w05QRnG5cgn30f9UrDpFfLtm9FxOzzWzkRbPi9
fCbO6K5YeuczNBAnPQtXvE/yHgkbAdBuoPnzaoa3K8y6EMAIyXQ5nVR9biSlJrju
MnnFQbolVmVLlK5+jRoE63OgzFZxnQr59OJi8axQ8GscbwJCvuJnYI5E1EZ3wUyS
YMP32YXg+tvoLAu8S4bT78puCP78/T/kzBKKiGkasAGHcIqnduYcZJBlS6oYUJ+e
NBoOmlG2tmoAJZmKZlItMnmsflgsqPI4yyDqVL0u+XogQ9B3ZDHZskMDitB3Urle
grc1zB61FqIjOSODMB0FQNCXfEmTC2rG5OvdN5iN9FpBDcjRMf3hbxytHKAGf/Oq
jSeEafzXGzVulTU+waRtjY/TrxiwHd2qYbG4wVUO1c0lNGOjnNVpZorWWMS3CchA
Lehwmi9S8eDVIbQklBwA3nKNpmyBpLFqKSbShSzAtJXMj4jWlbwlzWY8kYs83NDy
/6bi6KO9rjPBFE1azsoXYbSNwh5+D0liw8XF2TcGHR2Pf//Ntb3LEGppOrNfSEuS
sVO8inwiLHxTZd8c8h832Z5cbPTiDTeJqFRU8j26mBwdZhTOZPCvN4yf9AS2F16z
zQKet1gDbgqY/joZ9YKCo1vtjwxbcvprn70JthqXDxdOxB5Tc8p0nB/L5OAEPjWZ
M4cviMwRSEoPSanC+G3lcHO0N/7fGVyDyeJ2eSseRNfJt7bD8KODOHDPeFbUeA2g
i7THM9mg9iXUvdr2WfEz1qLVTITyf2szGhCmZuJL4BUrjvQyBPUusD5lXBxYaTYt
Nlp2AksrEuwDvhmA9MZR1owO5pdlGGMIXi00mHcDH/LV7ZGQ8lBwSPfyUApAnOvV
gQSTD7ttOMg+dzBOPGUkqw0rtCRhCqV89NTmAIwYUnZY64/4nf5jwDWK2CHB5I0N
YBvdphp5oSlYzmXEjU1MUaws+JUKm2b6w0s/OuoZ2sHQw7xJsXUJ2WAH82pw2pO8
Rozzf6alp9+0VY0DbYSImPvIjPEQK4nnd3T3njG6cvsrm6PYNiTTrDhnS2vKXbt6
+5fHFLzcP/JgHk9Gld210OZ23N7Eb0q0+3wLwUWbNzwFpbLFZFUYY9mBBbPUh5jM
9Ant8uDAlKdMXh67kEa9mea9jsZFSMOJ1YDGI907X44l4J/DHX8ViCHUoEX0yBi0
K6IDnL/Kf++EGtUuWI/jdf2yLIbZu7i07c6uRfyrwVcHi5+8Pl7VoOvOHFW/+4km
6i1k7K+LetZb5XgL+VZ8m0o2riajkf2Hd0XP7UmrLzpkAzWndpkJxVCFiHTYDgW/
EamkbDEB8F45vdomNtNz9rDoaykr+31EEre6QWBDhVRJsF1R+qcgQjIL2alTs4Fm
hlfXGllXIJcGblhH5OcT42CMh1+wpEneP5vgFJ1c4PA6UY8qg4BAlmj1nGgOKL6H
C8/L8/6RESZXRzbdgkDagfYme2ilowGQYqqKqsOpHnKsuY0obHmqGjB7WKIzNpf2
TjNVGmTWtZQkRUW4KJsdBS+09EeEre3oiKu1tM4/qlMq/BgZECkLCq4x+uYrSUDL
Yx4/7b7y0x1LHfxN2hfAxO8+ek9z76SlT7yHFt2N6GTch1ESSjY6lFcRCwyqmMAV
/C+TY4hxQI2rfy7W4aLlAdcyr5jQ1VrSC1iqwd2B1ZUdsYK0/a8ve3n1gxtfpNip
fGvw2CRbUfWInfs+f3293Pdvh22lq0kg1FDnhlRgFsvkFIJ+07J5FALf0BYRTgzy
QAZ6I9ZOVUP7DKSlvM4tJXgSNHtx6GAq6nsMz15cWV0adC15K+kC0hDFri3f1jbZ
y9h0UWOmtHBrB7V3TmadeJu6+ux6YKv8ZMlv2ch/xJ/HeXs1GjOFwvLnLjPKjEuM
3QNTPU4kSg8u3WtO6ivd5O898T0ZeWslGWlVH1SxugLktPZhd1wkRU+uVkRR4DHd
7D4zQISSCSmEV3ivD2ubwBQgvbPEsw7lGrcu1EhMLOI0A+R7aZLC1X+yDQjr87E7
1hzgP2R6y3JOgatG5PHgBPHSShO132K61dimI0f4hXUoNIFjYSW2Prt/bT/wG2vO
a7kgxZyQ0atdUHaxTg3zJhsIB5x+TdUuIimENPLD+gn1JkBSbTBFOJt+KQk889xq
Gpf0YcezCKTNOLp3RwYmOGa9iCtcGkePB7+UguZZW2rfJGCFjmZm6w2AVqQK+iIn
yP2m1HgCvQJ7Mpt0+tneT4EEIjCaCzkcm+el8a3IWQ5kz2t56ENigXWYJZQM1FgA
6NdbNsNbg/GFaPSACxO9fKf1mu8Qm/YNCG59CMKdGkGoH2k/c7TQwLxaoG3fp/HH
z0DR1jHBfP0p0DPWrZiuHohhdMgqVx8JEKvNy2nqXJ0NQl8wYf9m/uz/os1Owsi5
CuG9L/2cBWHgt+EkXeQMQst8+BWrdF05iiZv7LH4IK81cLy97V7eEuKM2SaDSibT
MRTKHV908GD1ycT3lq54ulrR8PS5LkqOsdlgl4o29bO3E4pqwLFMSxpFN5tpvRbM
I3f3rTkN/2KIWKpv6U/7foSirniAuZG3/48QHwjwywK9Wvmb7szdjYrGkT/I8BBz
tS60uRCEUqQc8kyBI4jwOvhXXfx3tzAAA2xUUlk1wahKpTsSFQ/vFt0026L09ZSP
gnUG/VrMf1+nLOBntVBWhc8mzLvIJAzj/dl+BGvxIQaPzAX51HdI/dKFfSuruixK
lUo3lfG8uW59MXmgJjm/NZrLoEXUel9N1wpmcSUxzidSwa/GWP+GjcySPAexmV4y
DNDAL8Gz5XsUWlGQOMCRTItr1HAZsX0jWKUg2TsaS0Kso1zJ3NQjJ2qVVtO7tWKs
SBMLls3MiZUQPGQy2AnhVwY0BFNx6Ba1508OjA2SKeg7JPsFnsdmLbrKTv6vAFYO
Dbcfx0kTbb2O2yp3Y/yJLcy4ku/Yub3ofIjoS2f2FLCCjJUxBwqxERaKEm+zGqbT
eTArvq7rfeG87UWDw6Ok+kaKWWrUijGKqM1DmvHa35IfPelR2hNnKQ45iVVaMITB
wPrk5jBJ9VSzBy3LospvY6FToO9HL7XgqqCe1aPDSVW/j0fvA55J9GD6K1OkeY2a
MpAQJoKLsrQcL1IuyuuOSnGbVjK0rRGM/urH9VaQCC5zvca2FW8inx5PXBr3clm4
5d8FuJNQwOF12wwSWTQS3fStO+8jFKEk84z+GgGE72fq/YBfJkQBK+JIsLDKVL/l
Dzsgpk45aHjDfL31XFO6r3tRKAidFTwPOhT1VFuU2H5WL+LO9Th2oFZmA/aFpfiS
PYyi9r9Wjn+xnMZZeqJJ0yszoS6asTCd+vCE3ute+ho1xtmuPluW+10CNAV1Ongt
0o/+xn7TTtd2AoD9ETM1CjbDeldf5/ID7FBK+1gtNrfGF8IWmMg0fTf+9qppcjcZ
z3QVjAzLxiIUdmaGmhZiyQ8gpO6IX6z8sw62bkyZvquzCmRb9uLbncybER/xC8WF
Db9ePPnEfijTHo6BT+KvlzrMjSEw9dqAOI5NnDM4mC5kgq1iylVWidlWG8gMjxRG
4UQadyucCq2/ATgRpyrkOSdwBIRTEbykgjodBsG1bOZT6eanN505Gk/OvbcDIf4h
cvOe05W6qOAs2/2ZQ7mB+5iq7WBEVAhB6w9+mAEu313MA5UcliNLfmxHr0QVrnNW
Yft3FXav+W6s4MneLJpthZdcRRFTybPwwTYN7/mXE/KUs52ujcu5NTcXPgHXMxUv
LBTMoA0TCjbervf/XYpJDlJB2oOplOry1QJhxEhcLvfEdCgci0tjMLhkxO4mpijr
Y3sh6my12fRIoUOvs4XyRDZfWSZz1jvu224NrYLBjLjNnWI6M1emgnqrYt0oG/Zu
vGazPCp4xMynZV8GjqqyAWE/StptBZKw52Cx77+ReX17oYkpn0zIBtOv/3cuRHUX
GQ3nReLaY8JD4TUlrzgSTJH3zY+qrlh6Ex2pCBG7GbR8yyZajU5qkwc41S0Y+Y++
+fQ9NRd938h3bKMDHAo4fPMy6GI9NPwB9/Jn9Kerw9K1w3ZZ9WiyJsR5az7NUh83
qDEPhBI55VJ4T09BY63bezR8hlvOs/UlkDpB1upTKLexOLZG+krYzK5rjr64G76S
zX59q2Kao+PYCC2IeGTiHJLKHtDjNEvuW18bRg72Q59RE7RVLH3DVHRO9AhA5HFJ
lM+piRPCVYqfdGUqX1VnEsTH3ma8SIUq43qPhW8XkvjBmT1UoHgx3slKaOHL2iKU
dE6qxosWOVdny4K3rPTxY18GVPI3+9wyJIrMxnvUpSQWV0BBszFnZtihWVGkKHS/
d+NdsnZVJJmtbyCm0X3vNVdEfB1Be9+LHJjEyNGAYB1/KE3950r7Km8B0HvJMdlW
Ihy5Z9uf81m8YHXTn3yEwYy0/gJEo3FV99oXv1xLaK0p6f3AUt1ZFGbTdsJOX4KP
5/HbFmJxhPvlvcDKByoI3j7WZZQE6bgBnM7RFnRX0Wr78sM4rKAyq3ap4L5bRfB3
DDl6FW+zq45mRsiMm48QscrJylbyY4Sb4dYLXvsbhy3cOk/r+dyvHnjbFiwwo+DJ
63pyrgxqrtxvKcakOyQ5l7XhFU4QlVojHQOPqCQfZ5lOiQBMPiKjfjG5SQvKPifn
NR4MBxnL1QaP9LYw+EBa9YVBShBru3fc5yldQLyso5numD4IeHZpYCzhrbTmd5cr
nh7Jx6bIgUiAl0NuqWQgNGo5xGt3BzoL+PTpx82P8zQBRaI9sOyWhnHEXLMSThMT
tZsGna3a4kMxZoVyffvkBD8ylRyTxjos3F+K9w6odqOO9dAdmbOMm+rgoaKHm5kQ
2xfAM/FYEV63NoUjVE4u8RALCJMqmnR6kx+WzMdt/btPOf+fDXn3ek2J4wxIOtdv
XSvbv63Qw00+p3Juyig5x2m6ML1XKN6FmDnwUQQS7o3zdbmxXIzLOjVE2+Hb72N+
Q+quAJqYpqYFf2COFCWK0M1LiGBEOWlxPPJWH2qAjUe1gU4r7+nTsWN1PNXT12Pk
SM+k/k1rjBvtQbU92tpRyi4uSRYI8y+IqpRqHh70NGz1JvqUqJlpRguGZ2Iw96Ig
WFhPnhkvR/Y9ppr5hf79fdjhaHRMnpkdKAUyIVTHD/DiruCNhyuzcXVQ+MzOkt7W
jqSfUHAzxelfQofnNyGMH9FuwyeaazMC372jhVBC6h1AHedXHcTrC5e0PvpEfkb3
tgsWamWBScKdS2LTEZLTwenHLMkh5oVZbFa9b9mI18MMOpUHcvtlwxSa4KOdfWTo
zsv3PTInBc6fwZcVlro0VrVl+iYSoGF04qsxRXuNu/3VuQrR7cDw3JqOU4QHwSk5
ycdImGL45IImXQ+PUcdAsKDuXa/TG6Vi0KohGn2s1xCDojN3YR2sdIDPv09QiuLy
F/UkPoLLTQEJCWFxL3PSnQHOQRsU99UOvCcRnnJGA+rXprVoeRKMPRJzvG+gJj/l
1XBmAg3OedpcLGRtidNh6Q9yg+tXY4BNQRkyKfEXMK6jWNrz+2EzSFhVA39sJ+5W
ptFgxm3JFeDxLuKgRTIwRe1vVieOPmm9RA9d1ZXb1o0HF0OA2GdwHldyZW/b9SBo
q/Rp34A62GOmyO9dI5gmm1pEiEC5Qq7KMwb0vE7wLRTFqch/sogvOV01Z3wdddA5
DE/yTCJOCR374GGGa3WBxm/7B+In220sny1FC4gxIWZglsPwiJ6M67PRJCBUAUjh
6MTY86Z14hb7BQqKsZla5YUj8INAs8W7DsnAVucs9pS+jWJqPz8dwqI8RE2mMS4N
4Zg5qUSZFPftPAt8nYU6xwD9+CXg9ETwJxOo+MDqcpyOorPZoy7l+ukQgBUaXrus
t+Tg7i7eNloj6KLxsuWHs7xkIcNT8bqO/xU8HAmYffnTHeI4SfQytPwtZbDBSQxs
XAFaMyE4uQarPMb89dAoAjzwgWTUHOzFk7n53iqW5/cmnwMPhiQKu8oUCCOoHrs6
EaSDNPhcQse0Il6f4enQgezVwoAoDAnpj1g7SGMgKK68dOtY4DyPgv7VwyhPfyc7
Sny4HzFHebqOhsjpfYxcSUrCFqhVY5hDtjT2v4UYXHruV3/wbcmXSETXHBbpnIzJ
aRUlvDoioDzrfADFstDY536511SQnoIKF+p/hpcCVpobFv25Swp9NIuT9zJBH2pX
Dcu8XA944TVK72bJ5EObFYEwKXUdWVEQBejHnelXwTkS+Ghk68FUTKjcpu2ngFzX
RpKL+x4pCwhBRMZZi3qdqdQ7Z5O14e53MDSKU6XstMvckaIQBqA4rOvcsmdtQY7D
g1ZxH5HuUNMtt0yoOHblMdKVWe8jqr1c8GZEPRu7kRRsll16dIE+QI4yaEyD5wbp
im2XjceLu/4j9bO7NMDWeCkldKuvvKGxdJmu7nZM3ivf/H0s7GerTub67ZNeCYFV
RG04x4YWDKHX7/cBr3gjNLrzZ6y+JRwSDTQFircoguPXp7A84S1eDjRShk5PPttv
wrXh0vGZNklkb6bRFMDC4OE24rLPK4hqUqv2PNceMx7YXti+bWCIV5aN8V9KF7YI
raKOa4q1sNkgdTrdQ5KNNRLeBkK9liNF5MeGyYvveaxF3m65QQJjWK/CfuoC0l8E
3fdxuX4a4IpwLMZ8ljzChxB0WCGux/oCI7nkvmiz2IQh2RaZridV7+HcwVwgxJJG
h+wdxli0ltYP72kdxXu7fVDhegZ6OvmjGTdeKsaeIw8KubQJzGVY6twyH2z4flwK
Zlj+37q/zdWP4DNAC2Wu5yuBpUnLLbDma7fIRplrzALnyCLMcNiWg4cJmQTapAqC
Nk3GwGf8YWpf9CI3Q6XAzoRaAMFSYnA4kboW16J2++28cSUfAmTbFE5OMSTkOuqV
CMblZ8HHZGRXtxzf0Cwqr87p/E1Qt2RwJFmcLnhssU+PWjSvD1h4LYKTpiVoKETp
jxuyhtcWCwP1RRSXKV9nve5QhrhL51kVEZLzKA/zv1zy3V0p2Hh1cTtb+MIx8mfm
L/8v1zRae2RWiOTUHa5yGWC6rGGWoIndYIyx6IXeaogC/2gaziqNxrJzDfXAYfwU
xM+C+cs0kRFdJEfwPKqfiYnk6BcmUhRNLGjqrV8lXdx9DtpxkP0C4T+XsGuPa4bl
+U9vlMHCttHlbIGq6eMSbyYuJUnTLJ0q137L/sqbMmMp5DSwgtTd+eLZuBFSmA0i
i3/PdgeGLETPJnAakITPFdbcmjzkmf8rdq5QtlOv2P1XD8CQEhJq2nqmVbWaxnpo
PKa+dMB2xfMtUS7Ac/jsuihWwAgmiaa5Wj/yRBbPMqI5/wzeqBkk+2UTRawX9rpw
6T93P7VCevx5yI2Iu+PF4CEyNQZ5vCbOiwq9YN0Kw62k6UHDwgiy/2UqXz2YFFku
YIA8fr3tsx4/Jsjh+zyzTBz1cLNqtMrdOoPs2UWHiCeJ732jrLsl4ZB2FF1aalXv
tfa9YFzzFQB+mAC6q6yRU54GbX04iikI1CPUJPZiFp4e35LhU7g1TEABVmbqJMDb
aN+9UgH+UN0qofON97bpcg7mm4NaAa8NlulGNP2fyd9gJQ0Igp34wM93UkjQ5hxz
LnXQTHyYUEPynz/L0t3f3GU0A54EB6nVUO5MitDJG4W/f6DDrvYGBpfFCZk0dyti
bTt0eJBh8axkfHTJzqKDMM8Vrn230dgp3k92xa9ysB94LvkRZqbJtLmHkYdmVOt1
teAJdmvP0y2OBwqypg448ABWwOv3IkD+prqYqlkR1ZrWQLLTxtwGZeGR17SgQiFN
i2E6TWcOAcqFkk2LIE7VQ1Hvb4tNHTFt7hG0gzvtbFf/l2evE6Apb/xY9E1qZ0UR
RjV4zjt15jAndeqZDNpmOSkrktN7258oZCoFnI3y01Aj6Un2ghDjOSYVl3Ur8cCG
jKYKPChFomfsLJqiGoRQHNdpSQhIS4xU7yGU5WcFRnuIao/63RKwRNLajYIXIyIJ
3OJI+j+we0grJh0cnB9fofww7O3NDs+T7ijU1ZOdLU4MDJkSxSxb9VQCddr8vMUG
56BlD9oqvSSMdVSABE3QXKOI4yfGPru+G1SE2w67trfruKGUJfJN22gFjAiJ3Emk
uX0lensqJMrAluPF5SM7Ql25sNX1TsBblrG6bFnKWKLVWjE6KcpHC1BPGlCy2kze
n74FCU5lRuAnRYTKxVthAip9x28zeyERfkIRkQDsNoNSwbWhW/OlMMH5SVNSvZo4
1KIf1ZCaIxpWxw2IagI+X35VT2kCY2WWLKXGBKQnlNv69mK2gWBIXyZtVZtonn1S
owKhIpYhyCmSBX2To/IELUvWXs7uWH0+K/2ZIx74m8OZyv08nanI1f/dyhltVrwJ
SnC2RWXJ9Sda5rbcCU3L0gqPdNJCi6PibQlIpaDUMXydZ5N6Myfh9nnc3kAZtRfE
Wf35gP1tgrYjrpX/NGADqJBXmgfzupKRYgR7B3gHOlz3mdpfiq/PBgncZR6VUPAJ
sZAjHr4sxjXYi2318J/eVxRd7I/lfgFXdApCJeDN+6tWeBwdnpdfUiLQ9/Z5JSbx
ROFkuDCscwmqygdITa8LgEmbWBKU92iZ11yupmNXIDVKJmrYo3Yo+r8o2sAVa5sO
rG/C/37BdO88OP1ZC7CSRbA0QtHAg8A1jzCQbxlaTKT2ITMN+Lxf8AXZHVhJ1RpY
lor9pFFR38CRe9Hzd4dyrP7qTbcUD0hXm7E5UFhvl7azq18CIqwjy5UMPuwHPP22
c2grTdEc2pwZAQF7RarmcyWdHf2OTdXwoulkEEcm4qloOi3hVrs+sA0YxsKKQcqh
jiyLeJ1o0U7i8SVQQMw9ERG3I9TyoFU4FeudD1e7Edkf3ICmY4T8NZ17jFgqgNOH
OUZacDv9R7gbw5WpOuNUFw5vECyRIXZSP5H+82AaRVfy8eXu8Cp7s7u7moK+miG2
YWLYezPp3u7edmsoLttVJejeN+HX80npSW0mP5eQE0I57L3w3dN0il2Hfav2FmDJ
5Ej45NyNNm6sCg2iQie75p2DPlb5qQc1sVzAOOz/eWtP/GjFfHn1d1kTIcdHHJ8E
Wz+3rKa7ZcHgzRr41lc5MwfrOkfRYuk7vXQnWT7KhR9GAtcFvj+MT/0KJTfpm+es
fx40NOzI+TZl0kxusY7U5dIw0BEKLb0sIJS4nfIQqo/qbdCeVNwLj7apozIECgjS
F8yDOINzu6Xs5kFaEZKYJiYO94YpNBMccqfo4qIXrp2f9iJHkxGfBfnT+vyTxcOs
BDxJtzd1PPQOaMy6PDEc5vayXmhp6uRWDj2M3hzjFfDUhkFcHFMqmQihXTOgqL66
mLHJncXw6I3Q8G9N6ln4EbRui/2SzNW2uaS9XGsaO1Eb3J9ykZ+JIsaRK3yclbtS
QkE+Pee3Oo5TloNB/K52eACm6zbfBeqg3xXCzwPwZkI+4FuBEpK4qlQT7XahDARq
UqshHizqkRT6TqmO6hd4RZPE7jVYbHyP4DuOsZ5/C0fkbr83aag7FdJPCczfEsEg
hrewwJMvy8PdGc0ucQP8gHW8iSqz4NXqGMwgY5MSkQwMXWp4Ftji9KkNLhEuZsnQ
btCwL/OVpS5oFijz93zM/d2ydtCSQS8g7Rq9l3tHZPrpJ+/XbXC62ob6omdy1gfk
fuNQpWjCgUdunKLk//Mp/CPN3sWRUKSZFHOi24WQLwGbrYFh9vh+iC0SMrM9wfKg
vFiYy8GoBA3Yh3c0X4u4/iZffpsALcGEgKurmDZKZsiHafJyXDsYQ80uLoU1ZdrG
fej0dFFnA/ll9+fZbemJqZDImwUVhtTcTo26Ug0YqZdqigjqClnISUn2hb0loh2K
QMNjhc34tUAj1f6w0dZyvxVtZOZ7IHbbIYMBro8c7oo3pffrvpAR9bVkvCY6jiYO
gEnV7JlZUxkHjRpAJLCxSl1FW2j6JqH4H4wLFjA5qkps8BZpJyCvvqARcsHfLhtP
Ec0RDBNtc2hvlTA+DD7iXNn/Eosuarh59GfdgP7Uwl6fmt9JtayL9RHIxioBTOQL
Qkd7HcwpNCZOWjY5kIrFpT0R0brs0ocCRk/+Dbv7b9nOCJQfBotSLNxROGIA0vYu
1LSKYnCpC0oZAsKfVpSJ93Jcr/zH6t1z+riA/0nExNn0nuTXXCui9Jry3hnZHRBm
GAWBjLz1CkIS5UcmkGOs0HMp+8pgQBSgcTRxLNIe/LoN8ZcYkc1oSUU61UDdFzCo
8ZKZOwzrgqOBGaW2EK3og1Z6YQlribp8u3JjtbNZ+/sVoqif69nwqN0pJRSToCMJ
XPqyP7IguT+dYr6ifp0uYKQq+BSzBOzk+F0dZG1Gi1dezWF7K3GoiED414e07EJf
LzJwy58Y9BBzV5mnb7SSraMsZsk8L4pB8U3NNEmVicLJotpB7xW57sPga5x81QH3
z8HJuonJ0AcD7Niak/y6vAf6zvo7A1EAYHdSnRDwE+g7BD9RCeDQlKl3NB2y32Mk
z2CJOFhL9f/qE2d8nWZR+BHeNc+pzV9kSMxlk2rIoEdNET9GTS+Gqk9P7FlGZcvw
oUZRSTVKHAfUYRK2J4Wos7QS3YD8QBLqSHqCi+Qbl4llWZfyGlc7XRaajUtktV3w
QbNfIi9Zq5+YLaBIJ5teMLqVOWR99Zc9QaXkL4RRbyxdggbDh+lE0UIMgQntlZIH
1obqZwsDwRDas0ztk2aKChLeJZkIyOS833PPBXmModXxL7WDmMGKYcXbgCZ3wlWk
CtEWCT+ART5Ii3rc1PGB66VZYJXE76RtaR0hRRS/4yCklAk+6c6z9o0GVSHI5kSY
HXSs2f4L6fiikaNV/bd+GjsO0iw7yC2YbdBYNHKfJZb+ADClescuneUuIf3AGVkA
N2gmHTukT3Wio4RzSi1mxZwfwdE/0pFHNQzobRjfK7g9qsbNEM+tJIon4frmtmyI
MqUTeC15rQiNHksB92tLoVRsx14S+7SPvjXPyplak00uK+PytEwZCpPcUS/OHSHG
33Q+Tvsek64Wujxn79kkW6APhDBFW+5XzOIpOsB1QWmIgfs5XrgelAkuVu1HCPC7
DX7qUMylQRvRuc20WvkcqQiXCSWY+DSa0Is5aRzWn3/510CdbvitYz3BwyCyhNhl
xjQbn/XoeEiUHFnSMGny6BmZHuFUAZVBDDNRIz/0oI0kQPi+qC8Hjiyf6jPDPuL1
WUf4+yLwMLVrIQWjC/yiPqS97FH+8gVcGxlUcW8fYoGS1z8eZ2lPPwps5HyGCl62
QNmGt4P8yiBRN4e7f3FRtdHi/FxOE7sLVSf15kflYlXyqcyXvr3oYkASr8YdjLn5
WI6sQ4QD7Q7zi2rnkrxOv+t9tzzhMYEDgKJeahCGG2dnrScWi9ls4Qr55Vw53E5v
JPGvCBw7wBOfkJQg1nagcoaHeApCFVpsfRnVROrNAUVptXVK4O7Y+1g0FbSBshld
+qO3DsyLFHR/CFQtjaJxX10O6O/B2vUSZJekaCAUAVypTMen5r4AI926dpnleQDM
NL5+gOQLrOwMg4+zDyLiEwtxd7bIGEgE5E8a0XnjmD5RKYj6q55qK/bQs+iZoxpD
zUhS8KIzfLSiEul9Nh4ZwS05/jBkXeke9J7j7SEFPNAmLEpuarnm2t0VgkN0xGhm
WvP8R/kvhavHOx1XudrfvZCz0jzl692UXlVxfPVYpaofN9lDOOQwa9X1oAUapRCi
5Y1OQhhJ/s2HkB7KlvmKdLRmE1Tp2m82ckloYhNT4fOfClQAZatCToLkhQrPDxy5
AP8V/w7cZsKdYFzNKTD4m9aaqJYolhCo8Cm9taoPFZA/cIASQNJ2TDN5jS3+MXhI
C2/sUarwHlowdESTU0mKA0LCe8cRYZWRLgcJERRyYxvgAbM8wyKYmMJItx26t8Bn
LE/VNVNhBK8TIYTJA1wcYml8tjTu+4Yajg0k7SY5iMmdvMe6s9SAZogaPmf6Ssk8
+2yRpRDeBjVr/QqW6CRmNgVJcEWUKePpYvZW6gIM2MGn/k+yhoYYs72xeNDJBNOW
VSQaQe/GiqypChty87dJQ5oXMQshkV3Jj0BGKQoJEytUw5k+r5+1HkAqORvHm3rN
PysQ9bs0xlITuiqwzJtm82FuHR2Jme6nVYBKCJh6RS5iCXSdKaIOlgBt/T9EBo46
NWIzKryI040RK0Wc8xWP8q3iSxH1p3zJU8sLpG/Ok6xVFxnx55Xl3hmppxCdGLyV
x3AxtGIW381kns4/UDqZgeF2Qb632j4H2UjoYl7YtTGWRtyqIFKoJQX2g15vBw76
5F1zZ02HcL+XUed4toF42B/8Y9RWz7QW+C3GePJaj9sUgteNeTgX7Qpxse4SALQG
7deLvjPSOhZYxurh+ESdS0Wa3kbXUyuYxIw2xrvJmJAD65pkjn7bsNgagpmOKENi
95J6ruaMnhhqjwt/IbQ9JxD03AKJ1tXJdBD8nfXZsLabU2VVBSIvafZ93RqsM3Ep
CWe8J53Gi2bspHSzi550zdaZGdVkR+2azLNIV2imXqEASk3WMend/RcDZ4CP3LwK
SJs2wk54uUb6hhcjfThwLa0VuRDHnSAnlEJ4akYG9ECoCxtKvI2qaj2vdEcWSXkx
0HCKg++XfzpfuxPWvByvQ37IvAE6G0iLJS3/eZCHNn6FoBvwwZi0aF2oWyWOaV5n
clThgC/KOROd8eNnxzTS60X59/Y1M23aXOYdAzMutDGRlndhkjl+HfsYvEKkVikf
fvVVf4aGO2v85P8kSLKylnf6+4Lzb4GRVVBaJIhGS70md297K4xtjisicfZV9GFA
kT4je1eFuFJP1MEsu2jK85C0ysW0OWWcISvZbzemB/+oxCWbjsZB3PKd2qxzfNzb
Q3faIAmUilQLhHmZph3XqA/tHB7gAYyIueX2QrfUUAdNlAImSrDETvQaPMSq+uSy
WlcVPFZY65A+kAPNErrxG285mi+IOx692vckPN8aev+paEfsdzzEVw69lYeH2m7p
YJw7oEv/1+/z92dOIfncp3FCalrAuIVzhd3YX3PRH6YAtUC13a8SLUaDqVmfzYZi
SBXyMwXHwKVyO55GjQEPj0pM3rhXJaoititnYRRKhDeZnUAFtW8fqueIZMULXl6k
xpaZO4halw68Uhr9JSo3RpbsQGRq/9bJELtwJ4wgSL0WzMLu5wLkm8olQt1EA5bz
0D2e6vwprvqtJ/ayO+22rBsdKkn/tikysA0SsNrKIbYo2G+AX/nRWlgJnqYdBNqe
VmxyoAi9iBOcXeatOJFmX07Xi7+YcZXhzcEFSWwOBRGUJQvmd+apqIpqTqeLqd0y
f2YSAQqVnOXa4Bc0s9aRN8WeYjNF0ZBD+yBH3lImka+zM5J6senyBU6TZxeBB5NH
18UhAjrhEiK7oI05+a/apBrw2+adJoBlRnACe5AeFYcTLxGfkjZCCjKCLyazu5Cy
GubjL8eiiZyzrVW/gd1zxYpiYeJ7j+QYAJWhOC/0OBDqDZqIiibuH1abl69juNKk
SNsg1njQ4rMmT0tyOBYifYTlkHL+sVOs/0ThIOPl3aO/lfhn0prEM+3pP3vgQvty
CTGEDnlcucsdxMMiCfbPmwkyZnfbqx+zuERZgOgD3TPmgieaK+V0fweY3VJErGPU
nsAQxsSdVkbugOHQJRWNrF+wnmVFjEcAiJpfswEyJN5/RCkuQyWSbJgO59hJUn/0
wZVnwYJTSOiWJfTrmHR813MvBrIRP1muNISlaG88O03h4YT8yxAZqEHoXe+Tqo6d
tMbCVL3VzDJ8gOU7fyQWw+Ue/e/XJAyraXFfFPwshM9x/tUkeEo3ecv/Zhqdc6AB
p8COcSq7sD5v05fMkFDdP3gv6EDqqZAAGUq+DxAu0I1+/g3Yepu2mdSnUtxN1Pip
l+k3KQLZg2+kjlayJaJr04wQcw5mCK+H4ZDtwgLgANLaUaE6YyQwSECBmCYjcoav
b3RK4usHYuSHzq9PYFcUu4/026hu+g2QQd1fP6sQcX4J8IYW3lHOA+YOy37Ezo2N
rVz+8s+ojY2LuVAPnPk/p/7GElz+1DDdrz9uZ3f9u3ztajNpEDCNne87M9GF7SFt
yGumo7rqCH60treLT+annjpvCNj1XFnmexxJDZuQvfYpJhWNCbrheAy0Qa2lpa0V
jx4rt+lSYDLm32OfBxT5LtQnv3Wl+Hsre66vGgxRYyY0ddLLvmadzPIG5fcrNf60
O0TF4iM0jITsABNkoN9gmc4DvXYVCVCVYUGipE7DK43zld00Zq1u65utguORkZFS
m6GvYGEM26Yjyl6tbsUH/LGSO6xoxpb71KLR6yKYV3liOWlbhBG8vE9DjIVhpNIc
BOGnUDKPUCS53LpfmqvZ4vRqkpYZ2g5/jvqkDJdx3ZMJX1AbgZSZ08Ib1Fy7JhT8
hlF24Ry4b3GZ3n2lfgmjzpnoFp/uAywTvLoanHcgH7cOTxwYfTnPZ1OZm8wURp3Q
4kcCCOVN9/+MH93MWvqkxfQ8yTJab5ubObSxrHyhg1m5mii1l6+Zo9Lg7O2uVXjC
UyjXLbRehUsQOxmtsO9ManMUM65o9JHGk694XCaB8kNi0dBYwCQRfPN+JTGL5kRP
X1jz4YhbtKZbH3sDBb77lNQdFWxRfC6oKfM4Va37TC5P7IkmHsMiBV2icO6DwOPP
ETriM0Tuw5S3srHeqiHq6gJd8Q2cOOqhglmEPPhlZ6hFaEtiBuYF9tnbiXANzd0o
stzcDYiw+nQ0NP9lnmhUtCz+5ynJltQFUet6aFdRMCTU6weDyTRDtt2+pWoGfNb8
GYeeV7l6GeAKuvwKTd3S3OL9PWn7UQzkwBz/xM9Tm7QjOPzD5b5AWfkMTKZdeCzV
mxmoGZiFWJFnL9/WkekvW3ebY5gMbCEhLacf/PY1DjdEjF4k7AEARlJ2NFR2TpZu
wYRdc6pVjNW4YDyfK1e6uYs8GF1V+iVzO8Vkz+sKboFzmQre0YsDBnsRyeVQBwQ3
Uog92DCYI2PE5GpxTaKjsmiZkKy4KX0wI9Hxlzxv/VgG9LEc7XJ90MFnhn6xl0BP
eJNKJ6XOOFMhagaPyT4MqIEvavNTBURK3I/+Ls38GS308FooEbuS4FFDFS2OCJ6O
334rz8ezvDWfnokm0WeLYv4sA3KqFU6ATMgj+NQHdSWFIsTTeRFO92v7Xt64Na4H
7eJ5r3MHlUtlFX/dWGR+i3huwtPQjMhGHKQSeOClMT+E/PWD61KWoiJkhPFW3fTA
oxDlb5A1DebmBrnGjNqA/pIkXpB06ZYsECFNn9QtrEZvzXP0YAhhzN2cQihLuFbO
AX1TO0dwACfAGW8JiWAIM/Pv7xUWt9a17gN1CIDN99IjW55+oMAMm+MkKIInomY7
C0ZypZ1AfPP8y2Ra7KgCCGZHAnZNONRaf9scWxkbkqNMpJdjJz9C2ZkylDMWJufP
ftPE5749h+UZQJqVySAlpO+vMXkeqSAALOn4hyX5WYz5daxBgSeep+zE2ynC7USV
haMr+GZkYc2VLN89B4mEMcnKD2gDujPmPAYfcoGPpoJWUbOrVgYi4rKnDK2gK8i2
UE98Ky42vxUTX4guoB8sjOloXw1bpo99HpewggOF0YRDbzoKsVI3SRa1OtZxQIoi
sai6xDoPFnrYMXh/ZuvpK0yJbQHv0exLeE8ARypkHLcYbho92mRQHrGCX5YiEvR+
cM3xsP2F3i9gk0n8c5VVeElWL++ohQZl/rljN0u4ABr4NaBQYjWuwQnWB0He7SdK
c7KZ0rHHXoTVl6LNX09aSKc2o3/JhomrN0Q/jhbFwto2OFljPCUs6j68sLoG91aO
VseCej8bJzcKS58kXPgutJ/z/TIdiXoT7C0KpDazI5oVr9fEj9RC5NvQSmpAz0CU
w+WoX5YapPzpqV7dd5Q0D64426dC5BqPGaGgha1M9fxDK5h84XNEwvs/988pvUsM
`pragma protect end_protected
