// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
b2dKqLJDFBn3Isda5ZjBsUiS3iWsevkfin+F0Ldq/7CPlijYeeFef0LKFoVOyjOQ
Vv4cEjECVCPQVnR6gDl70fOIDpMjl3DNQtV6VDcHEcm8mRjS3RbvWg7Qr5Hw4Bq1
ppVFG2gbGYw4MaJh/bNDqAWXtlscY96DEJjyYm9ITIc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14864)
Yw4FVhllgX+yAsg5OMxouVFpgf/V1FLyJ1ocLXyrHBI0gNmXqvs5rD4u/pfqoXZO
qAQjmBgOTPb9PxGf+jdad30y7NqhA75xuB+z3QDUKXzmglcmukB0PdGq4nMchdSB
CwiUueytOTSC9KnmnEzMAkAASg6gEyx9RUPuU6tc9SevaFqyTjQnIS9JJjfq27wV
6WKjWGZpYBPx5IbEPHUnf+L1Df7CQazCaZshFcg1l0STSI95ZMfIaGMfhit4Harg
z5EO5DjL70QIsXeqIKrZmqwd+pO0THickiS7HQIm186pdN5qL01TMQh8cZVbmmNv
jBoAvn6sJwJvmkYatMxX4WtI9FNo4MJSMeXbsUb39+ABQmHvfgX6oBvKDmXgkF/G
Kwls3SVH9MUUplnNSMcNaP8LIryIC7Ze3HciFSp8/gkO32rKdPABgoEUqG1zMMiN
dAdUQMNrMI51u0C9XgD3aZGx7uk7W+yMu/jRHGyPkXUkdU5zcOghHR43/UfVoouA
5Rkc/1q/8UlmFmbOrjVUW0kpmLvaYhvcBDmNWnXAjIsDYhQIW+/xKTthL/eI8wYw
S7piESw/P0t/TuNJ/Q83uY0hB0a+ECJK/4YbeXsGlSQv+q02LV12ekl9IQDcPnnQ
x8a/xcPr6hyzy99gJAMWpiFm9mvKJdb40iUZklrMavgDqxGepcS1pC0NSbxsNNw4
sc+5hFlCEgXCyiGocp+sFvlWyWUdBGfl4gRRHFH5Pi/ohO1tjkHuwr6ynoko09Tz
QgyGtQLXTD4gStZ0KOQDcHLcjnKlpupomes0THYLYUWhNrjrIYnKQ0zabWZEcgca
tWlyjb+t0MRf1RXA/T5h7U7xuR7/V69WKTXfDH7Zkr6BILM7mHcJi93+XZpGDuAz
VIgVUd6owRVy7XTf2V2ACjsA9c2n99aeRckoHFaxCc6GUUYgDVzQejGsdvYmHIZL
u7HE2STnhFVLRppw/E9bDQ8XPbcZHxCLvyCQHapQ51GrCbqX16wH/vFhOMlztLbI
2htMrVi+QwX1n09MCJhfUk26JpkNTTFQ/ybhT+l/RP90QHfYM6D9y4nxK4koxI3e
8psr4IhSkijAR3ImOtzw8srcocmTAqXQnbHN4aijFsZNag3o58CBI/DtbK9R3D4h
sFZiCrQFivaQBKVlgtCZaV4vsVWezcNgXNvty2pH5mImjH6j+FKFKCL1HTLv2g/U
O2tETcAfLIVU3irAf+3ET5t+yW4lWJvfrEbUcRbvqiVuo8bvkp1WENxhbRbXuThY
02Vaav9ced7rnFO0Vg/luikcx6zKsDxiFGvG5iMgu1biWgbJUAT3sEWo8jwIOc/F
lh1hWzOnY3/kN5wBL8PX4u/WcDInp+OPxHqrAnRzQ265lDOb2e8myte/IQ8VwGB8
jH1mqcS1JNTgwT0o5fQqACfirZ5a4soDE63zknGp0vkPl/1vY3AJlKhPIzCp21z8
NLMVpc29BKFVU2xWBBKSNLLostN6+HZuAdlqWdOH4R77gZfoAfMD+gThOlCADUzD
RB5+tIdGqZh714rn8hyKwc8DKGmdedyxavTE7kFi+9bc3zqyAvQcPRL9FmoPeC3/
WR7rutALlPJtiwX0mMB6gpOTID4ImyNP5HqyVkEB3ln4nJE9bL0irW7DS96FM4XJ
WMwmljcPMMuVEvbDOVKvcrQ+cfXO+j7lsCoNtS8NO9/1vvg9PW6fRzXqifUTG23T
dU1nQoxyEPFFeY0434NaCAQY6s73LPKXaig5vgZCr9KuwD3Nu19rynDQ6JA7N9vY
24qYhJUWIl1Kz3iJZCchdPrzPXiQUQn2PLVjdUOab4qH+i2Acx/uOTPm+i/J1f2v
nSXDiKDQQb/jFWUGugjw1PdNJ8LYO0bsRVbzQ/ftiG60WDh+sc+l0M/9Qd+LTTj5
fArn0TbF/mfns3Eskh5o71cp19iEm/CDGAxEsRufOx8iV+TmX8fUj0UNZrhtiIU/
brx8o5KnUd6YXCM9Ddc4qjRuk47L8ihJFtUZEdVFPc1rCklBJ12clpmbmOA7qswg
N+bB6xT1HNu2eKCt9sjw1Z26z4hv2nBubdN3JjJ5hwpj+zixg6lsIJTsa40dLrE7
y3pK7/r5soSAhgJpGE7ILhKIk0GjvxcPQlYFoZDLwNP1iHGsrZR3zR3EYy1Gzise
OSF2pu6CG3IAU5R544elIqtY81EJIeryrebFGIakXobexmHUlIaAWeEuOLOh0B5y
ZZ/k2FVnSiaZLS4QRzQja/NkcaEVvJ+3pV/fTtJtdsnkkamqh9KvQbmyiB+VKLP1
18VlY9+tgJFjD7pgNcZiBblrScYb6DM9W8o3CLBI/uVLKZgA3Ttr3LADi6xQ+dwP
zErQ8nRBiE9F7LglCevC/EZIWMoV7NOBCOUpvFlrqPdJrJsxINADu13bWD0Ia8RM
0Honf0UKCa1oOEpWE6UheWo5kMiUqXqUK9qRLCOJmu5NL6W15OA0qBGLV7c6X/Vy
4VNOvyyNaEmvNsoM7erALzaWT2t5nzyIgnSdSLpMGh5LNHscR9uQ10WTKFX5xL9z
6vtwQZnzZQTzzc2Q8EFVQm+KhZdEXiVxG57kqHNRg/e/lL3bqQ9iqnMfyTE52tlC
ap+xQ2npwogXnfV7Ci80UZjP7+6XwimSW55+39OewhiWQlZsGBdIfwtq38oBYXZM
YLMr+4VykC1oHTt1RUR0c6Ygh0kMzE+0M3h3uSOS5klpowAa+MwoRChOK+Z0JGyG
qZrjIAIlmTjz5xbdmSawMF9vlQb4j+oGH0YdtlXV6pLhjw5o45JaIsmCbeTK8Aax
gwOrJY25t7RZHIg198P3Yf4i3nsOARxYpT0L+c620VMUF4mA1LwKAe2WtoTSifrh
kUtB7igHjm7iLTkKUrFTU8Foal8NmWvUw0otr6E8cKrati7aDQ/M6PRPKdeLqLCy
5KrYfxVaSrhA/ZiKZda9Iaoz+eBfS+JaeOSYGIlFJndBYx2w77+rqjYSS9c15h/L
C7CCW4lj4SeYN6NB7DnEpDq1fx3+N0Orek53iIyIRIMbNaQjTMBKiWkUZJhRwVIG
d3UrcT+Vg5jRZz64U6x+h8m2xKadts6xIzVTnNKqDYKYfIFI/tjkSUV9lX1zc4HF
yfoIJQMKNH9vDidtXx0Dvq8GFemub/FLREDfafutkXDUoi03dJOjtoGjvfpDmkVv
Twq8RItddl4RSGFsNu2OwXKlp0t/9m/q/DJ7jQboexfuYILcX46w0X1f/CRcuA3X
QTsGa9sjoUk2K7OKFvmHbPBBQN8M1nMzINK9dnxscRfSKTCIoAMxqyzR8L37aelF
EsWBA1oNsF+19ThvyhjFeGErn9zEBWWwieVgksCji743GXFm4xCJs1EE6z2E5byt
7hzBkGD5+Pha8QKoLtxT7Ih6tzh+TggDoKglkxYbKzFj4TReBgObHJ8eBoazDFpz
GsieY1KAtOp82ErQaLsf/Nz4XVjwhDnF4/JVjmDmZM3x9BbdzFQ75fkmEavh03F/
UsSyNBLhIOBD9hJdsYPJMKCsPx6A0RSArUV41usTqWaNocrVxKLHXj6DgvDFX1Qt
ITXBdeLrTEieHVuM62cX6ZI7T2O4FQFCuK/74yun86HL7xQ1ns+5PIx220+CPfGe
LOVY2lbIyqHC4+J4hRhlbMaHs6IuCPxEyPiutlQncI4o9RuAqHlLQ7jHyMWe5cd0
FvYtMAW21GufQHUOk0+by4H4c05Rin2cT5tHTmsUm8DbVjFK2CFYYDIgbwt35v1Y
0Edwmwjpt6LQfGn2fvOlmpi1zAK9p2u2rI3hVCICxnv5MiHiTmCuC7V4hfRwHYAk
Eg9yqxEHJvVGLlYFo3fH72EN32YQrrrEVImneogzGsjkAlJoHtpiMv1y1AnyY1Vg
8b5LOGrSXHdsVfn8xZpk9MIepGX+8AmsC0hUqYTiUFvY6zA8gjZ0ylxNmgoHmIFh
BlDv7i+uwuipk5A0F6OncDtcq1Yi/tipAdeX97jyZNCnKv7gp8p13GNFnhrTneOL
ysHuyhZdMf29scpR64sxJT1e1fj9CYt7euu4NoQi/fHYyMHYbjVU6oAl8emH2ayv
Cr1EGQeyn+/EmXHzx/79n60fCt09t2WdoJiJIdjrq5flBhMni3EXxffVh+S7CGqj
VJHR+cCWAfF9XggZFsGQ9EOjJPlLn5wlDQ+ik20admnwzEphPrNZweFq0p9xzbOC
yMl9Dk1FxugrKCv/mm+cC1wGvRCe0Fewt9ux85iZsuJRBBlpbomA3zYL03WtCXYT
Ii8fE1pPySTe2bPqvdK4qxpG4Taw2A9qDUx9enk6ydM3ULTiuhqPSZ56eRqXknKR
Ve+V1Rzn/ASpbpQwkAngp3mZLGfBHGV/TYxQuu5OWYroVOnjzVZ/Y6UdCMQjYKd1
8G+6gM3057jL/OQT0x2nRxS/tdfsr6mArGNtwh1ZogN6oMFXSwj3ouIWl3XAoo5C
QiZ0ksyHoPTFP5sVcx62GUKi1NWk3Vi9D5Gnxp7tVg43+u0877kFDI0idsU/Bx9c
5DsXY8nq1eOof6NUL7C0olAVmScs8XsN2r2/Cy2Xw+Hnj44QQb1GasVV87zgLKYJ
bHCW+KwxpIn7whK8w6NWREh9buteigNpfrGRNCoG/GYQwfzHMWQGYeeIBtXchEBe
Q/INA+Q92nqjDT82hb6gWbVetHwYpGNBZhxpuotTKDto8yybYZ8TwXKFoXgvWGtb
D5dm589GOycJ8U83U27dsEwub3Ho2QlVrjYUIzWU0oLMOsddhFH7Fm8+guISesUq
qST8b7nubgwladPLrUPDQvvdWQcRsaTQoiAT1xfyr772lJXpOCvwWGi8pqw13wdc
6LGOxcIWFF828WEKFu5NOu55iKHJXjeOG+hjCEgKjQdT6S+nh5oYofWIqUE7+qvF
KVyLg/xoQ3TGfVQLHbs+9VWuiU43O8vcGqzi3MYe96OKa/0+v0aeYNgk/O2yYZTK
X5BbF8BdY7GNGhLcZe6qp1Ka3sPl3SNCLo0T+ztdtYK0Ofkwlv+nrxT2Ej0dd2U0
9pxdLwa6R+Re7IUJd+NrhbnjB7PoOYRGl4zRkgVFwv9Sbl1ECVzqTo42WlD1SIp5
J2XyAeY2/x9xgnR0llEt4k1qnyeMdcD8o2ztcgk0Bx3ihKDxcvaYnf6p4JJZUOJZ
YYlTfRvovxzR5uTmn+pM6we5f12B7pvLkQo0rSkMTxjk0kaO2+FsyJhKe4JCYsAZ
iPZq0j6WGoS7S34joaYpk9fu1wwlpuR7dH/i9TW1gMA5cdUN9xG/0Z/8hGUyODsV
hcMSZhFmF7WRx3IziIl1n7KH/nGN8jECu2fzcQP+YqGytK+Z8hSC84SgASbIkI4c
69h9DUzPxSbPrlWdM/K4bKu1cj+EcHT2zjqXzdhPOMp7erFgSYLi92CfZjeQay7k
0CsG0gkn+kpGywFeco9/Xcdn0OSJhJ8idcRiMDsEZ8Sxaw3RPBo8nGkpvrxIRjL/
7EpuLvNdFzJaYc4u0+O0XY8tNClQo+r2tYAFZiHZHLq205tKuyReflm58+m9LLNX
I+UIXHCOEz+nT3Ya2pN0Ep6W1xCE5aIokGHWzpFnloreLlNREN3QFvfooKb0O50U
ewo47O9BkgdCNifFrUL6OnodMyALihIUYaF+Ly0PKE+dJjOvhvx5iCqengtzJZt/
LkHz+z4ydYetWyuKaV0M55OR+pufZrJazMcB4liCcZhI/ZHP075UzTAKvzkonXf4
D4o8aN2JKTN6PWWKL2y/NMSo/h7lumUGqjGYHRnrmT8uUsnEd1kuKL0xvyPIEPG5
8bh57jRWAqrMXICsFOMlUtYrWpEJjhouI0XRBvUK4qYZXzi/coomF7cKf3eSOWUe
76Q3jIQqsQ+9KIGVwtYmpvE6pY+kj1L2MyfKcacoZoBmA4b0odpYRHNxv/RgMzho
FSD9Or0uI79WfohaoLnO10QbA65ux+cItzuBQnoJB2CKaqbZd0q7SQxIqyGHK6um
sjE8eCOkM0QGcbR2q7S90wLZOet60iBYp/hgvrjLg+wvMYA53rlkob6P1oUmhA3X
GuAMYoGfGrFGSOBWvuDIhwPdunRaKV1E0dCGdPrALnvEfW6NJgzKs1/vOKEChdrZ
0v9IqQj75+ZAWdjCfZHpkQpEDwVMod4NbCJ3sMQbVKhCoHmltTwGDexGhl8GnDL4
bB1mUD4lcbao3jcb8rymZ/kB9J9xZ+hPBjQ7n63XhnLHZlFDr4jmH8Scx2If5/Ms
E+3JDbRPpoqpD+E0DHoQvTCR18ajljnaiDqibcnJVuciDoWwfQHtRbeolk7EgwLd
HWnHHJ5aak2zXC+ecpbGs7I3CNw5RqaZoFfeVmv/3RTK44H39CEtXgIgvs5rjkIm
hOWS3wwI1sIfTs1UweDuJXoz5vq0ffrhR7v9khRxWEmcYAXDul7Odf9jOAhjZHZD
mrWL/BL+STx7PLjk1jXHfHFaQfq2FZnyhYDMCdQ8Ve5lBR7FKGo6fgYSfd1RO29Z
IJLv5DW7aEHjagRxZDULbPyExIy8PP5ISXMb6aK1BbwpaDvDscv0I2B9az1Y+Cr4
DxUQIdURtFeuB1g23jC+J/5zT6O61p/D76EdDbfre2KDNSZK0PEDEN3YBvUq5rPJ
mLSZ5HazAQhzpCPlHvSBmJfeGkwhVZlH9pGvoPtl058rxGQXt4t4G7sF234mV7g+
Lt0//r6IONyAtY927b2G6q9EACfW0qOlwOiaiHi+d2NVmq7tINcEgXvIfQOBR9M2
N4y8wm2L0dPt4ouEIbwIqz2Fpi2qZmvQbG5oTNdktFz1ProJR6yN6LOeMZJHP+AO
DMH3h7GLx1KwvLbFukfkWHxhiqlTdxlopD4Ol6sPF/luvOOEkt9T/G9xNN3plprd
nhXUn0fQNQ1+kjSrspsqPPvzGyOvYp9180IlDiJVZsj8r+DRxzGQslKG/t1GnXRE
JmDZnHgzWaq9Brf8XtVKEf0dnq0tDRQvw9FTn0W9dPo3jiqoYcnGXkf5b1sRnRcl
MpMwKC4Pe+5OJDt4DCMyBncipB1FZKbaP4E7UnkXnFbuUytysFLXUwTuPpRCsno2
pnBHGHVswY8lhfzDzHzW5jDM/YEbv+g/ErH3gOaU0Mwn9K87s5t7X93OCYmBOKPk
+JLFwFJuaqHQ9b7Da4i5yIQcYSWYp/HkaEnZ5F3Qzm/wwQwpaqE6T2X55YL5AJf7
FOBOby8Oe7535aUMj7JbROlGyJAQwLNBphf4tIz/RTDIRAdiJMYLjjIXTSNvLF6E
8kNgYCM0Ar+jKW8y3JI9WkPOmhhFyEuw23XXdJwTEtsB+/dcAL0YM6qgZA1+ghIZ
36sndk7Ds4OVuwzRhHu7k7J3vDr3R8EdXhI9tPqQTuQI7I/wGY42S+x2iFNg3eIR
8tT5GBzCwd4TgYQhToM2KYvaoffOsoWFmxvFsYgNqFJe6GXiJM4YBTcTAiHIOK6i
fpWnNFXEW2o2mADctoMknhew8Dr8X/LY2pcN2r2+H1UnyKUX8nqyLt1mcfxVFW7s
ZIMe63Yq+1IZUndhy3j+ktCqIUuUWRbooUh8cLzz/ns7eAMJ0JC9WFxiOih/8vH2
yRk6btUboRKvu1gb637DJ62tWwGh+QOJK1igZGnKAT1TLt6fBRaC8rhL9lEXPvHr
NES6JXKSd704FuLnSR7xR13iFUD38A7DGCDNfELgUPdE0LeQ/3uZe5jiJ1UmogzH
EoKSf8nUh5AKELwKERZYCv8UPx4ury4L/v7coYWcq8bVXtNJpnq4XDi3V9PkkzL4
ONw47KFN6U7I/C33auPllzmGZ3gjXlGrppVPRhaXM96+Ys+0fzWSJn5oPu/QxPW+
qHFXoaFa81Q8g07oolJDtUufatCmTyp7DIcNYMYzY/CT7JeLNnww0WE9U9YlxtSc
1uZLHpMMBfrmwAuHX/Cz4jOdeFBQSCd0MpkO92h8uFFBucC+JALM+wkssmbYw6fi
qVbZWAPAoQuiRhiX90Vuqejhq/szDLX2l7x4wFahff1JWSa03GRPEiNlIHxZ31Tv
vGs3rknbRJcF/YPVw7hVJm7vTaejiWxJZtVo9mJoua37vcI2ntSBJ4G3s+m3AXRK
O7QAlo70uGOw9KSn+WZMnPQ4ywjh9xBVac59Sgi/cYo6JbbDH4twGs5tEd49PAgj
e7GhLlaAp0M1n6682LIAF7x1MuGej1/xQLjdOJn3fGVajY8xdez3C3hgKfKPMQAc
caiweObAA0RnMDh+MRgKWqsW+UY2uY4G2SyZWWvEbCcWKxiSp1JFv+vPspVMNrjz
Oc2bPHtg9PMQDQUEJ1CoPTxcaW47ldhixqdHe6idtlsN1NgBeZcLsUOJYQyMWpDF
WNoGFF9ams3KwROzkz6RCwAmaI7l7DggwFFr6gwnqYCVuBFQuQcLtnsHJJXqOoP/
g1+j8ayVTvK4lQjNkPexPrXEb0ODtiffBH+GOCICfXl5Edvnc6igTl9Z5IzAXm+i
d+j35+p8C9zZjt7NF4eQNDW4bilKCHu15wTv4VukAULDRUfrhgy5Dk7Gva8RJfhg
XiH2zDbTD7FBaULK+prQircMMHbXXozsX4gguNll9jjU2a3hdCzjGUtrKTXJ9nP0
BrCKraE2i4RBFnpx/VM6Rd0QkmLIoUFGlXe1j/8iAqkGvpjuHGvSelCW76Nxwf7a
PO3Nr2dBwohn2ULR4ya/GCbACMWA9Y6DbUCZh9EyVJHdk/7j05/IAJhAv1h8qrkO
UTLY2xj4LQuYgLji3D5tRP3EYvVuOu6JfpX4NR/NUMnybgIbD2FDotawNfo3aB4x
O4ZQgQkNy3VBHJbB3dwEpHuqbaU4G46UnzOKNcY0oJH93me+3XWBzMPbFYstMsMa
bdJKsTgQuL/V83HEJkGQD4C9x/Wi0pjLy7Vo+S1GLBAemEk873cfLiSEnGBGkuVC
4xrFJjIP3cVONwv0Oved1uBzWpfSOnoYuANMUBWQkNPhv5feGOw0hRm3zYIwX5jR
3BQMHk7GDUYJFkzsyi3B3xASssx9w1wbT55PQF3RmnpRMFvhxn0UYjfUjoXtgOsN
P/wCpOwYB697QOQfSWg70iXoPJbuQf5l5015OBFyrlKHznO8BoxEJ8r0Wk1dHxkB
sBis4dB9zcfrr/V2Tagaq8QFxwmG47k1Y51YPDpplC+MEDLsY0f6tULcMYYih572
I4j/7XujM612uM+Ig4IJok0j4FvUuvBVj068Vci754waKpjYZoevx1Pg5Xa1xp99
6nC/eQtUD5nW1whr5V2IniTrUIAiSO9KSNVmHISa5yNRbtjxUKOlgEgyf4F/s73I
c9W7pHtuc2ryv7tNcjIYlrZY8JuhqTxobyB1atIBNCwdAhoNsfipZTxejlDc45Vc
0xC0HI+QmW+Hnr1KJNoZbzbe+vCHD8chWdwBA8T5px0dpb2v1xXVb/UJhBJYd/i8
JXeP5eyANJzDp6bfYxQHj1QIzz9X3Kw86phHdSlbiT/fg86woBPMcc8ixzX3D+QA
t22E5+5vdvpdJdM0SRYXEuafD2OaShLHD9b2PXuyw23rONI70BTUfzhGfgdayZoa
AzBi35zvvWX3WEPt2PETOjB7wzIoOrWXshmN0OKQ8LPqq2STbOdeS4iwXd6sAJ0d
Cn/0PF+BGiNlXeXp0y4tV6FQB76Spr7Td+Ht558aifnkGm/QVf3MtqLybumsmqZH
+IYkzyvciuJ2627lXQSxdyDErsXV1ymM70hPtvE2IstDrltDmaJZqpEvWiFdBG8F
hxxXsRcRjwDz4p6DmO0IRDT0pzVjqe3fO9NxLnPfEwmhoJgc5YPDDkUoGO8RNGuw
ohyYHvUI8t7EC6U7IELMCnEw/DVLQvCeGjCiQleYFTnmIZA18GD8WSaYG018JSjE
tfJQXC4bAUz3Z6Yn5eP2YMlVboRWic1jptA2IQ94h1plL28YJFOp4hOJIi19Cv9X
36LURUPK1PqnY0CvQC1zl0CUi8u+xd8gw4rBv6fjG7zFMvkiGmKbK0ZgTjvTD57F
/VNG3xHhxh4W9nRbd200/CMEoGtseWgG5UPnTan6InhfgJn8SO0mINfUVvtEOEvQ
e9RuG4CsYL0mnf3mNBuxjPMAnJSNE9MHwjEl781TPKnmpqjOb03oqmwMuHNBPnfH
sz0xlFZwBbxHXtT3zq1J2qhF3jUpjnKrdz0/WKLsjPqE5a3cIkoNFYFORt+tpM10
cLaVTiWMA0rWV/LrD7TZR2cpaQdbN3NKP70sgtURl9zWnAX0CsK3ZrVHA7heuXHP
wI5qDZfNxRUVDqT9BHtdEda8PKGjRqsyUwHn0Ojz/NLMETZxKZw2VW6NFi3jyafd
rLXikLm7VplkWp5lQgoRj2C5FqHagwEPOifID0iMAXIRtDyNSrpAygCqnu8e18Uu
8HG/PhlD26gA6H2rBjVQ6ynxWwtp1T/S6CJvyXHEFpzJ0kWotfImPmk7/5sdUP9C
ntbk+k6h6pey7LWrlkJcOROFT7AJ/HQD+pnPa1P4Nk88ZV7QzJHvNksYGxj2n5lT
B5116ELl0XSEKfKa5tqLEw49fHBNMpCXM0I43OYHHWNgJfGpD8WdwDPm+m3yi5Cy
ET5cgqrb0scxxFMzUKv3YNRiHYXeUo5yzZRY/wL4TzhyuqG3qcr3U/R2IenuI4Zb
hP5ET8Pgfvif2TKuv7jcdwFPZVnh64QXhBld+7O7nzAZUJ/BI8tKgSsou8msrqHa
u+ugUv01bDt4aH4uPgIuo1jImalnNA9UEJbxQRXXDvOhsvmIHEpviiBRx4ijVu6A
IRy1OZz4r5jRgaO2Tx6/HlUrsZ3xHZljkP9tWl4P+iie5+OW365ynDJp6Fk+UJTD
gph+K1EWNSwrey5UcRRzqNX49Y3iAtD/3YFQ5ojlsYlGjNMIJEU+yYZamBQSoGxj
5q2Lxq28bJIpAdNy0wz2l/bjPtSpDr+2U/0c72fQzfSqock2QqGoUj1cVtELlXuG
8zMe89kofNCgkiTQzcWmaOvRfpqV31rBz/7F2f3pLYney3O3ZIvykxlNlXXG4Obk
3zDFkDnav/UpI3lZVs3CVe7KoBa9TrIR1BohmmrR9UA9d4A8y6N1Il1bSp9wM6nS
IW2mJpk2kq4EYpcL0vgupmqjysWbZLyK3Nxmy4QrpGpaz+9hzFwRCtPEJofIZ4mk
xQOj29BsEE5On3c9dGOJ8dLr3ozcSHkW4TC92STPktCYGY/A+K1zR+e5dzY0PX02
/0Lu0c3XOlhoR4WQxjadJIH2KxZR5sOgq7Fa5PZlndYuG5S5AcugwuspbRCd7mVA
0OnI33p49KYrDk+MIGm5rzC76s0XzFHI+ILNst7megAa8ywqqRgqzOn5MlSuB/q7
jue8VcGfj8dVRZswA9dUhc49sHu6PNo28ez0e2fg4VBhPsXwHPw2MXGzMQU/7guI
MzAu0CdyMD7DQDjHq6WQzrCnDTZd9BPS+v0j4vSj/e/UkO7p2EQPKbAklb22dhPh
AdUYutaYyJrDkPXyOhDqXThsIN/SdDCDFexqApeCe7Z2bz20rkDcZkr+sHzS8UAe
A7sOMUxAGtJoh2pc7gN1uN6lvugLeyO7Ooo+XxWa30vayLsfH1UKXD2HmqafptRb
/qgKmdUBxcwLTVHd3XLGaqcKKbkJj7sdDDXShoD2jmqdQq57ORH5u5vJHtG5KBZy
l9O/gcme3jSiNOGMepN5EFu8CxlqKa8AEhIZDx+5xck+/5MgSNwm0QeQQXcIHlrT
beINsj0kY84Qj/1o0lFVpKljBTM4SKL4efSYrdYQXe5HwnzYYEZcIUqN4+HGHytn
S2l8I+psSwiwn0o8/4Y+biXfZBtsHTq9x0TwNv0HC9mmpqVHMoN0KPaKed5K2fym
5DjL2zmzB4b2QtzjID0g8Sf7ZZdke5cYQE9E3IFsxSDezfDywX/JVB8bq31hs441
+wEZllcMstwItnmzB7rXAlhfE9SrNkDGcVHHPaJD5+kmyMq3vZI4Ob5xeAHjvzKy
SP6vcbHqfOhyGblZj6NC2pIGjfNIuL/UtJeYgVaz0960MAtrHPhmK6NYv6iqDtvR
A7rImo3pheHnpKiZUI0AiC0pjHlPkkU2y8N8ht8+dDwRxZ3Za9rfW5tk747K5Pjl
CMCQN7NfyzWy0RZlr+77pwBWTUJFOyjquhqL03nSNuYa6OCHP/cwJr0pmNrkNeO+
+2aZDmWsDTUOp0UK04uqpVHdZSdoiBIIewKpyNgI7Q0me5UTmke9Y8k+PfoSuMuX
pft7tvE3mxNBFu2qQgXdoelSM8nzu2sbDV7U+6W5WV5k64Z5lSK2pZRYua77/q3c
t/EWM1qdnLcHrp5isNFAJvTh+hTq/04u4FxdZTikPzRKiH5sheQnw6/6Ib8i5UB7
iYdc7o7rwpGUtB3A/aAxbJ3FcChR+S16ofTraBMa3Z3I53tG5x4pc0ZVoOrzl+D0
muJzMFfZV85wbJzzJuX6ICYjFj2/wSOisDcfAGLTUeK2jdCKKgRVSp7Bhx+579hC
S3Cl2HYY9k680g2BDKunDY/6parM3y4KuqsxsJgfgRm4Z99z8pGk5WTfJojkNqi4
2qKO3krTfCpifFaCuu8Czfkt7H6UUY89RAvBYSVUMaOW0q3AUaZ75MN2pV5ugzPL
696y10n78bYLeqGqZsbIFcfGED0mQQ8qGlnjMF1rtwf0kahnRB5pJk5aV0tDzqD2
xoIS0sVPtVF5lnG9/mYWNwAOBAVSobNSfH35XOUN1uABTQLn8BQ4rRTaQ16FLzKF
uMKJFSuA8lTNaVu4thyKPj+5QFk+RVxi+fhQfdYe5nAnrygLsRAd7yz5zIYfSRuj
eMTSlyO1Ac20gGrNXzte/qYqzGdq2UzvsCFNbrTZgDbDQVpTWdNvF4aUGDT14GsS
N9/VSmfhNt4HMZmz0JM+8lUpcXpWVtNy9g+oIxijtccp6lAEp95UnGlzfOIQxbHV
LMurnlYPD7N3YTOz5Z8ld/tKtGqrdmc81a456B8OancDm9zf5crhkwfdxKrwsE32
kxsAet80YgQdRWyQy6pfu9X47P4aZIjIvqj+PfgG8vn7UL8Gb+n1MZ1gPhmC4t6L
uzeS4m2zsbi2Dgryx3FTCL/8oY97fyztQ7k1kPE8TCfxqpKWOF0n9uU8UgIW6LiU
vFDbzdf6W63Hyq4x1F5EEoNeyCH4MMyf2jJnDbwjzk+gIEFSQCLDhccyFsnU1m0p
V8ZkKrmxR8vzV0vEISt1ccbi018TMcuoyJDKjwsY3m0RWENsDfcUEGZIZxVIUlsV
AWAv18vF2DIaR5KOXYS7/o3cf0lwjB2LPSeLeFskERa1WIf90vLeB8Mgqm0wTh6X
ENJDRUqGY9zOTrn7HaTJdO5OD7aI9O+tPFa0jHlmcClDlVvyf/OkrMlFPuxQBSz8
AfxmXlCxnksCGxEIYD4unB8aYas0mUJVwVeCUc5++sH4YlIZRithpUY92QQvfmNE
uR2rw4Tahx2sf/AhMwLoI8Ov7s3NWXMk5LUSaMgSXX3EwMmXU7XvBFVzhAvAJagx
lULswrKImO0oIPqJY7LkqKHsAuEvsEbq9h+r9sumJG2LSHFaNTyY4HNgHKxzgajU
cqD+1cRdoyFHJQf1z6zZx8ksRUuscDTkgb1Z+k7WsdmwdnptQlIZqPAxs30yB0K/
Wt+Ex2xAn8bqunE4XeWLxoziAPb4w80tkGLZz4iZ9ndbJPPL/Y67on/s7ZVVy+8o
q1bV6HIbWx5GQveYcoXTTdEeEVbO3zhU+hcRGh5hOEXr3E7K0DemwFh4GKI5jVoR
QH+6lKmSthv4I+lChwXwHWOrWORz0kH8aQDN11/n+yJMbFtX03dgfg8Drcmpp6h6
fFsUpZKz2JcmONogZRKk0Btv6L/Dv6I/24ETtkpx2QPij6xusjpntjFdKhKWagP0
nXYTkkYT3Gz9Wgnkn3+RicUdByvWTViL0kt7086j434W+XzsZXQJRgqITAWSpF9r
AhVk93KYqgYe7l8Ke1tIZSYt/9CL/8Sswvtquj9Addtfd8J/owtQu+FbWTlmG8DO
8vVoVuyh/OcnJaeWmbqRkxZRR7Pt4MDPfTNpE0iQw5MMnR7zgZvDSYNW1k2jEzR9
Wtn/uKjBfjURn0agHD/7z0QKf0qCSeCiznZ/b7GlfuWWraRqu2QsShiJVdVnJson
9U53f0UpTP3wN2nK3O6EeQclAGq/dBluapk/xlq/dA8YWwkxoEmi81KfNEH2LNYv
XcgEJnNwWjR67Qkjt5unBqL2atrJkocImoxcxqNGOJ/6Z4trCFhgVUEB/ae5NHm8
BmEZpx2kMAlNRRFBhr79ZUt70PeVQ2sbi2vplB/wIJl1RfsavuoZAN2fTczgqNxh
mgc+4UkZxvkbXGfUq9sGcX4ewCHsmvVF93cSGKPF0jQ3OHM75vgamycg7AiRvu1e
7GuMA8WmTc9fsr0x4tgb4NxHmgl9MCBo5DVE1YtGIywECtvQieUqJpdoBWPTwplC
nbSq+yc7xw/ljAeD+9QqzsSPi5HsZMMwMXuONGirDLe361ue19gOZnCkcjY9sizY
y8DzYzxp9jJHFj6qNuwwOfthmXRCe1EK5VNCqpCwKy4QVgHNuDqQ9W14oJA8J+6e
wX6k6B5eRiTviLlaADsDjXhGoNxDXtinBvU5Yf9iBRjZcVMoYhYddQJ8m1Un7uU6
hWIMaEWPiJh2puZN3pSICZsZfS3Y1CYGsP+E1jKDO2i3TX8tsiSpOti8INqXwUfI
hZ8+9fCMWT5Y/0YxACdNfxMaxxS4QkxCGDXkzR/uE75pz6HS0/kGhTmH4dZcZaCf
NJb5o6SaK/tTYwEZG2q3IIQa5q1ScxAzHtHuENvsoPnZRL4MenjkMHYcg+wkg1+k
NpQa+7EshFzk14+gzHlVcNvfZtjeAM/fBKm/OacC+W4SRM8QKxisCbi+aqZCtLti
etcpWAetWpLgevhWUNE9r6rlOSTCriomhiLtoDTTCHEd7WIZNX68zcpXspb6d4RI
xzacsV1JGpYP9ZmvXrsZ8SezWG2NwDwOzBiN1924WHIPTvFsOityWYgE5vbBDjdC
zdgCZXS02PTphgqglzGyTlQ+gMICiBZFwTT6HDHr2mlTwrwWRx81S6Zv7KdUeXOD
VuadBuO1mW4PXGszIkz/D05mk2UQvor4JAXM3nFroTWBkG9qgMMQziq+N0qe9iPM
ZrBbUn2sczDPGoL1qtgtO0Yd4Vx3Ex+9To4r6hDBQNLk5pZvCKfwIKkJ6TwaiVVK
WfQL3BR1Ll3P1PANxeRqt/EPX07ZnE8Ko8O2r6Fiq+XFKFX1dtbOWIFS+PkyiM/i
byW5JRd6f43YW/kh0BfyHXILc0BuBEY8PAlsrifiESKgCH04T3I9aNmiNrZGJRf/
q8j/mD8R7LFsrDSmJHoUyWk/4kJV21AltSPuNcwJBciZXTZpROe2DXFA43ucS2AK
AOF9gYVsknbzISQTv1APxwMypzzhLaD2FccsKHSrZ0yfVpI27Il7RcJwsUS0DLPb
Hs6mJdQqOFtpBPnGwCNNnl0ogXjyeZIgKVOGC0US07INgKeKQLn4qetVvSDj5N8J
1Js4BgKjwOSYdvMv+tejFo4W1vojcN7CRFaktMdSP6qlABwcC2YDRaGytHoz0GNX
Q1Dr5o4iWGz1MMFCUki35Qw663AT3KdqeCEhKlIHhcqxhXzYS0OQBxGqJJsUS79c
G9LRnwTBBgkkN1P4HfjxAlgcMCofG37nKP7nAKuix4qHuvDt/PkYXoio3zvtgnTU
W2ssnSROGQOpXFgB7WKLFAffxKZ3bH+hrZj8qgUGXTMWrQpc6x1KpBi8ISypFFB4
QQNXLt0VCg3z7Tlogmv9K7Q704f+xQMKDgt5WGp+pgjjhzbYsq0oWjFS7sHVJEFq
+6tYDDM+6HrLd5CeDkblBQcJBO5B5YuL4J6a0d7UTyazdYkULzYiDjLj2qsxBDvx
JUVvM7dHdy/smoOZDEBFh7UuhlIz+ok0gRHHQ+RbVXcGXsP9BW4QRLFmHyuguvK4
+TY4x2rOpzr/pIFMtUCbE6QGtj0UkByMmVU4366GIFd94m5qpVC6oP4FjumZCI6k
88PWMZghwkNyJqpBl0JtbmZCmoOxwQ4jxeZF0E2NVcLBpF1nATYaJi5D9KW1W2pJ
pHGX5N5EHnOfMOenJo25MyDFsqgvpmHb9WwWoNoQ0smeanIIzMMQVGW/dnpXEE/M
oT/uTsEHDy4JaI1w0f2hNoTPp9LqhsLx4S51aopchQKBYyKlk7G+UUuN6A04/kyb
ggYrwieIGvnfRqto7/bV9cmdAttqinyXxI2OjJ6KFjp3351y0IKzEm7sjENDjv7e
FBZOJS+x4177Szs0OQTgB8+UiQCSNXylKbHSZAxmSmQMS8YYyuc7rE74e+NA0SpT
z7quTXxAmQcZ7MDym+G8aEBbbQZTYPhi5PWxEs8IgBZadDHtj6mnI1k9xtpwwpVS
flQRzKUdtLe5DtmIn834As7LPFHYPjB/KoTBHdp1u8pmhXr2UV+1+x230kamRAgy
UcTlQlipZxDwXag4anMVKDFh9pCyRWR6StnlIIcTmhA86U2/HK09S9r59t46GLSE
QVoZp0m2FeOMFKhLHn9Ufrhcsexpmae9IaC5YtShxpF7Md7QE3YT61mAhytIEB5s
lMR/ar93JXwHU4+V0NBdjjUnOj0vG0KZk6swVmP+UoZpQoKXhp/2MpJLby7C4hW9
kL7+JRgvztkToRAq+9hK1RRmxv0x25yPV7Zvr+mz7iaZZdo3a5RKHhosaAgO7oHO
xfB5AMUejwK9dlsH9+U9Smsi1TxBrJGtEIryxDrdCdc9SS3VTgv0Y1wc10R2G59t
3LtQwZzqVCDQ0SxXJherCT3MFdl1k6FJOpwuYjSgPRuTgYVDYRZUf08DKlNAocOj
E22VtL37Mi6kIlAt/F1185yDYAD+6yLxzVC/fr9TeV0boi2YaXrCfjA34AsjCLEY
bWQJXGUoDx5KOeGZQPFShtjh/4knKl22GCo8NKsh2EBilEDmQAn3ANDy/aLH9WfQ
+Jl9M1PaaxTRvjps8xnK5ZXPxYOnmrvAGUct/v7Wyy/Ri8l+EJ7Gdy0RoVq3Iotn
6cdVZXg4vdRE4Ldu2eErWfuwCSqyU/X8FdLsDURs8J/hlfD+VbCXnEWLT87cX4L8
6abb4fpT8FhCV2eef5cTZWz5T3GtnYpLTvNhCuW1ODwnVyhxTk17IQ0aD4DPPE5k
yQaPLJGgf6UGrqRF44pJbeoZevXcbAe7BDHlSxS0V3wTktADYWibrK2TyggFE62a
lo94jWaiOxPTAMg/9uCbjCA1jJEmcdomQaq36VlCpWWU9cBkLS/OvAnwN07l3Fzf
VZx9/ehxzG1YKWvDohfRJ4bYcx3TtxtCnt4WeVjkS7CQpmRiXCArbGRwFtu8uhtM
XXzKf4NRU6oBBcQ0P8QeiBjaYnvEtKtE9QSU9+gQdMeC3N+aI1CnyKsSM4HOh0Mn
U7YKWk+gOxE2mjwYD8w7Q+KP5A0shzjqdOkdVDoWwzpMfyUfnHk/+lKw+9C6/0Zz
SlRVg9moA603UxlzXX6Va1bs695puUJLY3Eb0jRjAtQ0KFOwIdY9+5wmkSPgUWnf
GN+YgQgBRWjtMCGjaxb1vFXtcxpDtSGrvg2NMIgezu+V3cgfwMApplA/tkwCW0Zm
1UG+594KlpeuSykINu8vjn5HI4ghMHXIK/ZWZ2ks4ap2YVC9bXQnouhNmMjtnJps
XgitekHD9mv7Q23JLJBxRLukm5aRMdzBQl3dsK7XVjwmJ1u37IeGWVTrTX//ZJkC
KpYGrpJpJJtyNR7/8tQlqZwf7GqqwLqIbjPsJWlwYNyDElzuDin5/yG4rN7nAwQp
PRR03QH5CRGVwmdbW/1QVhxnEe9UX+QW4RHnP+qB28350kmok3QTo4YdguCxvulw
i2il2AMJTU3wJgPtVACjVRVoDVMEg/Fb+rPW4bFw701bEGtYsFmxZt1P/bCJRKrR
HtyJ6VglJHPHc4cmx8u/j2IU8R+6i50K4rry+ni2TgkIbwTCIT9uAM2RZWMCpgUY
u2skpbFxQaN4GWhKKyH58SpEjYzsCGPQgV2pAG1MzMaZc8PO/3SU0GGNRwLD7OaN
DmLwiXIogKOZVW7WcddJAWVkt8jNN5ussqvKaG0A5z6dDLi482E7R9uTYgPqN4dE
gsZXbtR2eJGvjoiPuNghX9yNx3vQIZcfDVGSYzn9kP8FfxjwUmdStI+LUzs3ow98
6tl+M7lY3kkvKuKgAxTxJ2o5kUdqF69LveDUt3W3p8VThXS7imbL+8G3PXXz1tay
4Xf9aLVbnuIWb757/69FoUz4Y+Uyq/pK/3g40cV2LYu9aIzLA2YexzN3MjR5uoc1
keAeUJaOsy14UHOYjXkkLjOBv10x+sR62swNsVJVbJyVBslHOG6hvEoiG2fTHbjc
YigElUht+lZWBsWisi2z+M4nZAVEGpYWtXn153fFSSVZQWewwfkfxP/tjjVCyvbM
epRD7VS8iAurxPYzmJB4sPFas7tWxxXebqFvIDOEckqtIHASo0jgkGc7Fmg7I7jW
ed8/SKVZca0LrlzFW2Jg0K2fdyiCfhfVLEc17Go5lMCWzgN5xuTcq/+l52VslbIJ
hkT+1HdKqk/cE14F9e15gkZZDsgKdcLRjE+uch70NT3PMO1qs9UoYCTRtIFEq5Tk
dDBYE5ozQ10ZGKdZcw6GPCYjpgZ6J75H49bk3ktSH35F4wEjyOxgCRFfNCmJqJGX
tFDMvtRxUona4ZWZladRM3H4B3obN1zi8qZDqBQyBMzBJ2oxoFz42KelYNu7rTwD
MXxv6pzL/MbFXNUoM/SW/0dwu48Fdsmzs16Hja/OEwDO16mMtiZdrVSZm5KYTtFn
YKHcxWSg3N6ik6Hf7NaqBW38j5wPthPSLVOBfpiDhhMA+MrEE3EUlUHfwNRqweEi
eyC9MVkOEz1F1qTI+jnD9VBVyIQhy6DeDNdC7mNavo/OHSQxT3+0k4R3g6GvWuMM
E30D1bX0lEt87Q2HuJLDEQ90i4sZ67D1+e4v78exsNfG5+p/Lub1V1idBnq0kWeO
pzMC9GVD85lgDYpxpZo43m9ycZkO0lX276rX9r7gXSLBs2dsZ80HG+yCzBx8bbu7
yzl7/CNSLaaOgF/3ZHCoejfdETxRe1MFaaQ6+RnPEAYa8GSe3TXRvKI/3W6U6ye2
caOTnkaEWlJTy1xaGVcaBKyziLCwk0W2cWyEn8ri24d1OUlI0c0XlPYd0rb3bXKL
Uk4OaZe5stuxh9DcCsO9KHpxL7R24vuJJ+Y3jzBNk7XIKX5Tlm56R1LXaaLBUDV1
sIXR6bOrNoaY2CJb9Q2xn5NH4E27Oecko9F2wJVekRHiQFUu6V53JlnQS0t/3NWj
26TINiXC9I6f4sqQicOgH6fDkH9s/0wrqWa4fEXSFSGmZGtGcuC22o2bdcR2vV/c
pFO1I94ynArlFS8OuUPDJGh57SA5fJuVTeh6ZA/5quXrbUH7N2rZU99lL0FktHFq
S7ou0kBx7CO2CFf6tDJHgwivvjcIZuTmmplKarIZ+p6pjTN5Q0ceLC8spvW5AsKy
5MD0DJjPOiG/5y66WUNam07/0bUYSdpSZYsivtpXhtM19GJhCfey69cEEOJvnya4
4q7Jbf5NxqjSjTPoEa0gYJ7tip7I6cq5m9VPh2Ok+qlFrVqjBMxzUg715c0BJ9xQ
tb5uozkIHsU4o9TS2rAXfHeVR85GxL1fzWBEHQ5NGU4=
`pragma protect end_protected
