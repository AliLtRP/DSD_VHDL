// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EwGb0IKs3P4y65F9ihLCHefjLhpprY0anREtUJ+lp7meEuvVy08LU/UhsMSr3+tt
vTJIQR24lnKLdqq5iWH8uarFQOcs6N9un7wudeKkJ9Np4f0e/XYD4qOHfotT9hO9
wd4DB5QvuBjPetYA1pVEtZNmjGIAb+Dbt+x3vThd2W8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5424)
p2oaKxhAKSEWQqMfhnpP+45uO2Lx2LnclthikGsIbkwE6zuhUisj1QdjCJzsrQp3
yLt64ul6OyNzPpUOMe/T7hLNoTvEoemQUm/vtB2yNC09VdD9e3vAnv9HU2TldtEI
IBDYHQJNXgfoKMrvoKrJQaThFgFSVIyDYDzm8zOYMVHvZKLRSJwKM0IaRy7kkPGP
BNzG2tu8Sn7f/7tRIJQjSKyEQJxaKolxdm4LkM4LJ1ufuG3YBxFocJe3eKVeq4oU
4NoAKrGtmP2VyZxsc+EUcLcahNeIcJk4MN6vEeheTeNl0iNPZ4DKTbAwIxUQpSOr
4gyPwCU0PBymMLAjcWrBTnq0nkajWLD44QYBHlfWA3lGt34fygS1Ra+BUHtqsDEJ
0HWdfyBCvtMlJjWb+rrkbiWWL3xehDB5ajVzYVfIK21LWWY4NH1FMm/RFJ7vjF74
jAMn/fQeItbUDZ3j4ji7xCVwmSowCBba+ye11ef5Py9rLufPqH3hJX7Qtdwv4JvO
Of/zTxusxuxosPRyRmMXQJZX8CfgwRSl9uvCLTJzpd0ZLwoZfQZd4MI3Y1cdtEMU
IXkfDB58B+XY3QpXmd7CTwK7LD/NFrVHoPqabym21LksAHP7WSUGOWGQdH6Ok57N
75MCf/PTJjC51RbZhlDfydI4OMVy9moJOukNB1wJFsLZ0JaGK8f5XEjEEiJhK84X
BLf/RUjRr+kdElRTkj0sKDFEyYysa/FhH3r4yFULhi6XADIhhygplZEmfqJM1RRJ
PbU7e10Tq5KbTrDz341m5zbOUPhdcHswLrjbFLZbf4bq/7JvobkfHo1kSSWn2aip
GiY/ev4Lbl8mTfavgW+oOi3Z6MXe5weOduexT5udflkwh3+ukha/nBDgg0WypEVK
zWcTnSDnHO+FuUS5zx/wzBJGx0QqODOY1WSCil/7CIFepcmf1c3zmtZDCWPvdPER
dPV5zhhEcnl7xkXc0nIJE8qKMqnbmy2qZ810NSfL6CxN9DIMYzlb0SBGTuovziSy
DVh0xaldRPllGVYgdjLmxKBDI300zZla0R9rZjDfYbSHbQVj+Vo+UZclGI0D0AHC
8sFKtjuH6xwm2l/9Y9ajU8fF9hHbf7Xd98KVagJr3VNEGoBW0KvEijP2ZMordZf5
1S6kQK6QT1qp1vvNJxstJPtyiY4vhi6fU8i4mv1k1k3JFAQxl8m+JjlsaWt0sPas
GV3+WQcI3I6/8UEKFt0bDFxI+Y0/YXWtJuqgPnWODyrJcylhG+XkiVd4UX7Vbs2E
YYRRJB8t4C0AtXWf7g7IA0ySa60JeUfM3KiCVgNANety/qaDbhlo7tWJsRgFgw2y
6IwQvykD6aRe8JjGNKZqTfo4ucj1hzAWrunYDI69pXDmAoZ/Wxmgs8eXkN6ftZHc
lup68FGOJYiI8o803OUPPEGx1HCp4IvmtC5t/G6XpTgbx0Dxc+BuD4YFv1S8hSn1
s+UcdYUz73fZileoYSwhSPZlhFpVBP/bK8n1CmbW1JaDu2S8KNRI7hs0tryfy9HZ
8m2aAVliIpCHBOLOya2pHFHLCy6zVogviWZ5ctL8VfIPWKjDFWMDqtUHmsWqC0wW
DaW1GRvJJex+H/tzzbAswj4p3TEkDzJjJL/63HeOnIr1OKj8+FN6uilr15trEmRc
jsIyWrMyc9RC3t/YqG5qM1Cn0MNN8PjLTBUfQwr1PEW/5ZaLytTtYr6eMkU5tWoP
k5ZhpX8Llb28aPHdPKmZkR90h8zUruUyNRudKKvLAt1rlFawZlHqES3klgYZFXHP
zhErrcpUWxz8SnC/Nyn3Lj4nZLXbkCpkFymCqfkX4kY6GtMbkJKYAyZYK+JJPc9U
dEr8DiAhdPBVC195yF9onNwCDt5cVstPX1Mi5Dcw1AxOD8ZthyH7krwEkF/nLol2
rI8QUDc46/jgSyN6haL643yBKkJiexSezRdlj6PvOT5CRVFvVFM2L1jATN3GG5Po
5QG4QrsltYkML98k6pgtEzoAWI5dF0Ur4R8uN3vV7R/p13mHc0CpNYm7TX3gwW6N
DwiDuPYktq5H8peTV3Mz0sqhPuX/+XJ6krc0V/NT43vL1QCRpIdwVzOOWsbnIReb
9fpaDKa5Q+6yy+1kCvPqG8AdcJOISp27QQCLSJ3Slb0j0L9EzcUWc3J0N4QNhtEf
Ul62zoZ3y9jrPoa1ZBIe7ExHa7V5ndiJVCxOnFNmAt1o5I0aOVWs0y463FSZQ4te
WuDAPcn9ulYbvvUh3FYZrw2paFZgcDuswv3RzDzVSXjcpaFBnZEeV2oXuzqWUPo8
xSZtWK+2wsJlVN4tXtJ3MfWCVImSJys1MbCU5sW2mJv1EQm7t/zvr2gty+VBvDeL
KHFQJSDteHj2l1Dyuso9PrvDQH+vk/g2+MnsfkMRyurkJoNmcolOzKYHzVc2L3Bo
ajPdyXSJ/oS44rRt1gs8cZWBCnVr/aiM8Z9DM8aKiZGHPvCPA+AjBk3YlPtwvTVN
f5W4Y3rWGSTzawZFmXLHBheqPt8dpC3Y0mnz/7tuc0W9yxL6gsTfyj0/0MDKRwY+
QFSOCdtbN5MkRP9y+36R95vK3pLEXd4Mtsu7OmT4JjLc+0HuZ93VP6zX0jVfDKVk
DGj2UYXbFcyp2SwtmuqevvZ/QaisveSMdmP24m5tpu4xq3Z9Lzxkgi7N56as8Ax7
+vRG1hl05sM6WQq1qLPk4JLsyPVOTWSfoiypfKI+nVKA0tmyUpF8rQ8Wkvh8hZ1O
ctObSVAsoZruYaX6gJZGhxd4Yi39mKQ1HKO/0rSv6bYVHFtw1kcuJa9HBZSU6lVH
xNe1u2NKsyQwGgRgU9W3NdZ/QVFHQofvOgdvQ1iYRrGdUqZNju70tUdmCkLUNmmF
mS4+g/sLv9mNcQ/rplyrnqg4ekSyyCvtZ8EtvGTRZJ848WDxQaTzNAx5eZiaYqSD
z+BSpdC5KI9WP+JeVaR3lg4xmQZ+grbPEiGtaYa2e5oJS18dRmDU3bB83+7E4MuF
Zkw7TjevLJJNXTYyB/nADnKEm14TK7xACu1Uv9XkBRhzGI7tBuzoCnKC43eOhmlI
hd68nnvLxJHMczsWpAPUHqCQ1qcYK7fTjn/jNRzGE5kF/YeGlxWDj8hdIwG41Rv9
QpG597WEhKWakmjLA0ubtbs6EOpLfznaICxWpmmgU1gVU/0GrkjpiMqklCyvdQP2
5DvqMKlYtptQgJIUWAZ3uVut2NOTR+eQYC/seAqojkKV+KoidRbJEL+1ARCyxJQ6
oAxvN3pTNXnn/onR7Zp8tRd1YNKJIWx6d7BrPARWXs2WSOm6fC6jsk+tslUhG5U9
YPNAHX/0bDJnEkp/7mg8aUKMuhHHJ2APQ9NMu37aWNkMbpzzwiaOFK1cgp0cEnDE
1UpVSdd7JGy5IKz2xsjUuU9dH3/hx7W0A4KYsjH5TsbfAJ29tTOzP1g2XcvMjZ+C
OKgdaTWf8wKIrY91CQkIs6Do/I9eit/KSsCmVjAZS1MT9vhAK3U+r43i7CsU1Mv7
ikeoqc2SsogmOLYHib6CQYC+lNOIVWX/WLeTOa9D82POAuu4zsjn2uEjiLuJL2+Y
1huuJ7CtbcYpNNGB/6SmhzzGGDwTVLgV/tnH09G/ZmcZt4ncQrLfHNjxVNSQgI+N
54yGtaXTmOVPFg1rwJLXt9H6fr9MtrxWMrcz0lxVuBU1HbndNHib+NYAwvbyxH6G
BhlEGKjg0R7rLZcQJnJXk1zBUWOgmoC+RtcQE7A/QJAmmMz+44+WTrrNmcUG+SRs
o1UkBGd5N/HQN/fz6m4B2iAmXROgR2sFQfD/J9cuPz8b2QOlSnYrRrb3QM5cA5Cg
4snjz+pcXkXbmmRe70IJq0U3QuEgUqz30jAxYoRu5hXT0IW4AtQ8zAtl3M7mE6YV
yE7CrxEe3X732RZDsxDke2jpxua7hhvyqO1g+9qSl+dVKBBUYi6Rth1m54U/sPCc
hunj/wCZF0bHS2iUMnJ1NwYFQZ4ZAtCvauYHXicf93HeaaxabIyMyeK/KsoooPVX
rrO/cezLIRoHBiixI8MqWmYxTj4cQ3HztntFhOI9jHDqT4KqIsbJGg8CtdA4Q9R2
uYMiSpzBPXzdhY8t4FE6qcU+81JatR3THhSFoqA3N0MD6FRU9QSe8U/ih802jx2i
LCXf1z7/M2sDhA0LO+0iBEPZMjlwf5sMRkckNccGgCZEikMHh0kZYC2Gq9w+fBuj
mPERSW+9gGYPCePP1qF1WB3vpl34GK9S2npoO+Ld/DHGYYvbu0aOIF+ppijnVybZ
dGwC7DLwrnZKnQ04b6PqUL+YrA1QDVHVcdNZgr9XP5dXqJ0UQoAnrmLsZRt7J9ha
4mQdgd5zwS/AgG3HhXIG8tvqFSPOOcb9dcs0RhkjDXApzivYyHzIc1KedQToBsZa
rL211afnUoujcDtSqgAROWMDmoUVeJZZPthKGaVKyomzbk/QIrZHKolPK7aLcKKL
/Wa4YvxJ/jWXIevDqi/y9fjiNAcogxHkZXBnd6Vn+RkdqB3/2XCNUoPpngxMOe6j
PTyZJi3RuCj7a0w2JN9u2iM/M4qBg4IGb7AVaj9LLRxrvD4aKq8dykEfiCehSP05
9ylGI+E2M1lgODit5f/la5c0FnITl+ZKcq+b75IoC8hdvWXMwr8vWBR5qTuvV/ZI
m8aFNF1O6+J2fmLsZlY19hYHWB/7uU7yAPbw8B8QVu3otkSIAYnrKjccFFLhTTaP
CUXtxZubAwUrN+bz/jOBnEOz+9Zk7gGE7KsJZVWF2Y+E/nBRz4uTDz49EUkPW0Uq
y7eIqeqyddIj/Fk6qKh1XUibFH95ndjxJfAAi5+qLOklOx2WtkgZBXf833pkLEUk
LC7AJKC/TyYoVtfB8MgpjGRGAPMxOHbH2gIlgr7ERH1BFIbutYdRqQMdpbZXtQlD
M+BrXv/6WHZUSiD7QsomhCf0clgwNAZTAk8R3mH29IAgC+1yDL+RUQxNCAaeyARG
gexi1+QWlkVVrobZVvRMe465z4aWKgttbCX4U0KMkfXVo9/mzXgtNpYTSAiyRAZd
j2tCJvWJnJ6+9NVWLdsSfK6Ljidm5oHFx9w3NVf8JQtQQsWEUmJiSav0M4adKWcE
OgeV8zQVcMG2WqbLkIEnF+KVW8S18euxsByJ73dCO5ioUEFnvLQAsaTR2qma6E/t
DyFWbrjH7FHuwZhhR2W0fKDIWLyYAZyaH7hKK+xNCTmYsTfOowC53JGtB7/M3WC3
0GMRstgdcqASCf2FDwxrJQ1hdxkDADrUEhBV5auDssomEMSeDs0K1T+fWZaRleQz
SC9yhzj9XrP5j4LRSTDVYJGqLleom8gk0a2N4ISjxu8k4r2+nyztGUEHxa8RFvZs
uw2w1Jvn/ixnJDmdCORnQG2h5S4F8sefyrnxslPYL0WQIWjUu8GYzBPKeB5wcdVW
00fLYBTrrnukcenyR10aOrrs2tKyZSSIA/zn95Jq6xfRHLBzLMf6iNaX/bODVuv6
e9WR9g7CDmYgLQ13f/Om/UlSiEmzqIoPr4+FOQc1zqHxQhVGlYB2wTfLc6bH7Csg
UEqqpuHmy3Qa52rLWLMM2y1OdAnrfmriLAkHW7bglSBgYugNDdxASpsKB0tyQ8+D
qAMPt3f098qxkugukRlJlievIqri6Rqz9HVAqrbNlLkR4A9U0xi/s9ZXdDWxWF19
KRkxXMnyqIdk+LUFrQPxTORwTE7dCVzFO9lGaAntVPqRzlb9ZkB234YXMuC0TzXk
Vxlp/7F6jKUjGYwEosOnriK8COqsXDG0SL29Kb4UYZPvM5iv/feMycKHX2ZpdH9D
D2qhnXNW6fAw8Szy0aEpaDpmwmSohU151LGom19SIRabo4Tp7Q4qGVP0+gMMuPA3
WJ8lahn6xAAkQ10KAN8YZvlqRijvaCtNc4gwKJGRm9bahFNG5auTEXqhLV1nJXUE
rP9j3R3upcldNwvc1VPfB+kaTf/N25gNPbcGCnTJefNU/+NYmjip35y52gtS0TsQ
0Qc/h5JRlRhwbdz9EcRuTaMvIAt523PSVVYCWHWPEPWSjvU1Hu4Q3yJOQGf3Qrop
eiAianDVrDZnUtdWGPJfZDywZmKVpsCs37+z9YqpcUM0SJHaq/uycCCEDmF+yIIO
aTXpHogV78VOeXnu9Zdf2Fdyib/CSg/X4LvqPAXgZjqe8ddEF9/For/FzR6bPFlo
0zkfuHxjFODz4QrRDNVrDUMC0sxOEUEtAyXnACk9MD5IQFYEr20bX7v86vXBapY7
a5PnKF9TloTXBzEbRM9QeJ5Z4spzt02XFwbHjACYBaunm36sszOB15z73Wxz3qhw
dZgJrxe1550USZkt+XHOO0wgojJ9YMezvwXGAtMxyf8S+3HO1RLah4EBIpxBLnhs
b7bcFWHvJorP5hzeFOZ9ZOUwTIyFEKlnxbFVhB0Y4/3yc0sEyH2k6ENWK03G2uj1
Es/U+UdWd4ksxcwQFz1yN07UVCBSCTVG8EORYjrZyeVe/N3h6j0rz1dqv4ZBgj6E
n9X6AZAI9lYGVXoItrbb7poVYQz2WAr7f2MeupV2VlM4DoHHvDyklH8iCJSr6Pvu
szs2p46Lo7JkoxkTPt/WjhmgQsK6RMvy6EApuCOWqfLMpCidLqL3Z1hAqT17fPJZ
qfM+9Z+qg/hFET81E2lVIs482R6QxPsXoHGn/oA7m6pThJAhOMQaav3WkLyfae00
ENzmLwePDyVXDBKIzYm9IMBwraoMDkmxAC3ht83G7DupZbbpPRhGxwVMMLz2JPol
GndmgXwTet3Z9z0SAWnWgzJwZ/CjBU5Ojujpu1jfcS1YkQYH0ntsNRkITF+MGU6/
ZDJpHEVuT27t0yQFlvYnxt6siRPJr2hU5Mj8fJfcyJOfy5+IwTSRSdzXoIKRIPMs
B+tWUpGwAVEsQx5lDoTXpzFGPoI7jbkU/LiF5OQp0KVaCc2yxvf1ZApSzDyD9pwN
06mlUt8iO+qylInJZKEBuwxBZsluiolBcGNj90MwvptTU/d4hxEF1/jEVgSDrD41
wC0XjhOZ5tOaN/9m5GFrwLeM7jAepVbZoVIeX0MO+zvAlcBtcPy9Vj0xwuI/eYhu
wzobeV2fKgTOKRS0dJoQJvMaM0wPbsa9didGX5nyh0dhy4ign6ETmAIHdufhq14x
JU+TENYAR6A5ur+O7n8vEeHGHAf5U/Mv6SPPNK83ozOtgXdJdK/Gto+5FzLO6rXG
`pragma protect end_protected
