// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
DKsXqRBAu4QDhgs5UPFb6hpT5MgNgSTjxwkigTWXWyEjudEFcETTAiouN+hboLT7n4PIpiXdtF3W
93nL1rskGZ66AuV5csCklxR11kTBOaP58oENbqsFXS4viBQ1Nr5aQszSw3TgRsPUcdupCD/K9s5U
TTJOhNsC6k/v/8K8hw0ENGGU2gEWn2EsVOCL72rLNVsTT2Z+sBfi+GNm05oGu30ePHkWnCZhJ4Hh
2m0DSn3DpjZ4mvUMcPyUduQNZ1xrualUpwImKpP+5dCQZFot16Q7zwTyGdMOUGimRB3HavlSsfkb
MD4LWeRYtOOgUisAcrNq8lF7WoQzLtl4y3DnUQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
ujP9Zrcktp9v2p+pESEeNflDUS+if/0VO5KCGp5qCoG9yW6wYJOj4xiJjLuv72edwz3UGJR8cR0H
NgSzS+EmbDaIJU5UwNbcjH3eYgw1/MQk42CYunTIQJW320A7ZkKevd/ZTg0wGMd82HkAESbOHnGp
ltxsqRBEMqTJ9J8Zh1AekonO7YgvAfpoNjoKfPkIxh5wV43nFMDVF7Sz3dULYSXyjKpRH6B0gCG0
/KFwElZmLuhB7ltY1MpmxVyWWxQtBgN6OD2d7v35FtXUrwPEJQlGibUuEbeYWbYN5tMaTqAjGLW/
l1mZkLCI/VKMZVtytjdutH28z5+jzYLJN3lM30+iusHaml/rKwP4EVc+dbDsOxatotjIyu1DihvM
luhyS0syWgilVnN/372ttOA0of6PQWH5j9+kMDasRoLQfPs2bC50jUO4OELJuQeKHQsqJ1pLMMmQ
pzkcWwQFXXLxTpAdoAfV8OZB8dCqJAfNXXPyDh7/h/Sg6CWPxfb/jQG1u0nWIPpjMYR6S6RyGsGn
X9uhwdz/pUpY4ixi30i9j6/V/tDypK6/V0x96gM+MWZA4qgASZ6HS0zXTVjNuBv1NJbobLObhLFl
kyJKnvec2449Y8v0pXNdt89KKs/vawbu+/vl4B+0FBjxbMNDY6y/Qjm0X3pRa8STLeqUsGNE/kpt
xnPwNDbaVbZRuY/eQEevrvQy/5UHM87VhfzorsQWeAYCmhJAbQXQf4x9oW7JUTNu8OFdwHxLDHQ2
fdAAxkARysZj6igQ2j43yOKSluY77EhGWYulp8+0jcvhTGBAWEnEYzp3kwTSg51sKRO/tLjTUk3B
eNy5yXwr7+eyNMuCPKJVivXYYe/zfO5rpN9kZIrsCZA8gXJO5IeQqZaiFXLZZQJQzdMOS5n4CDak
3Ovqo2YRVsnOmehImZty0D4KSOkiUiAIoyueIvEtiAPKUVqqKVBPYWkTgHGI41lgo0iO6Yyw13v8
SLEKL4max3uXmpQDxOiwjVMhMYLLkK1dca6HZp/IFZS4T6PLXYYlR4VPgEWcZSSquoFdvFC6ziUz
2s8v8OFOiqiC+C4g0oA34fEQRf2gnvaVq0CXLdG8fNs0hMTm+3hRf5lGqSsv3rmq3iOJbnOoUNpH
HpDYRW9MSsG9aFCSUv9xt7ydiNSbpMtshTCgobaNg91otW9KPWFqS6VO6BR1w2kNwcPHzj21+8SH
Lz5uiAx4KUFg7ZqT06n1LwLvm1PB5YivTqb57/dya2boYg5iGdQzrGjlrqKEVy7yyCd2sWmJpCvs
/ocKx1ickMgekahQV8UlrnWNCEelHxG9xicOT7JuDggwK0NgRp7RPJb/abhbBGWFuQklBomjUrvK
j5UZTPS05QIOYhj/TqY6o95VV2ErUjrztr6boFa9NEZYsHhfoZ0v3nN46hgrnLp0yl3cybZDmq9o
LVrtmsFe6NstgVAMjWqpqc683k72aht1q1TDqoYmAk1oqbJys/Tr+qXtuDWI2acmwE5CdPcWA3sz
1a3oRjUXOplrmk6D1LBLU6quK7D3CqLR/u0+g8+FPiKmu652lPKkb+5irdf4sHjLB29Z/ec7lXq6
KOqUDI95Ts4oVKGHvpuvwB68HeLqOLae4/fK4FR5efYiROQDtWwlG0GDt4bEStR0WIMUovWGYlh7
oZVdnc53eWspAsuL3thEZIeYtthAMm3OOaECGfHgHUrJsxX+pW7OOPHL39Zxpxe/eHJP+mmkIXw8
NqxuVnGARb7un7wT5eMmD3/ClTE438Dd0wL7Hu6gv0iI26piUihBNxn/iOqMtBsXVtqTglIH+RX1
mVUD/IHrVBebjWz0zQgf7y1tic/ZUdOU9hQXH2lKZaiP1SE5JWBz4PZFxQxwAk6nQX0buXltkdDO
3cL2g+OKJJCLFnjv+wu5NQAYhSrxi1yFgo/YA1IlP3lHg+D3b0PzaR0c/Clwjv163vkrOaMDoR61
XuQXYVl8dsMHEqLCbG0GtbvPlck12mtBd7IToF7OZjEvN6A2M39zQjQO5K5Yi0v37w3q8Mywx77I
Az3KtVPQeRluAu5dcgsuww7rq0NmTcoTmKsF819gr6NnitCVpakvbwB9h832JQ1AOzE+VlEgVgTK
PTYf2RsCDwP7ETfoTmZJCbrrpFAzTi0j1v8paYIl8KnkzrNG6E9SwtzcnML0VjeyxMn0OBt+z4iR
2GH9D996G5oTVC7Ru1SdhvB0e4QEOkgEuoXF65DDc19IG8307mivgfIRoCEO+6HdisEudVanKtGi
saioill2V8TrYXy4L0lDhLNbXKGOBoTGGOKDzoVZkLKk3ddT6oJNecrXbAcEbO76fjzuVqXlScFS
hb4Zflqhz00vaAG3pbljWh5ZSQPRvVUCnxyZpT/KduJp2QKaJ71+VS8/yjHR4coOu9jTGz1jAHZ6
W8xc/+K3TMYMGnvwzXPSZwCe4qCUjaeDNh1EM9R5Pq49BtNc9Jqj+pIHkYPUn1hTgFJRH7PYE3Sw
y9W0DfAgfWEJX6V7rKG7lm48t3cbDUnfv0QKqWdsYverMvUQJdks32TCqNXlqF/S5COwoPW+7tOI
ztwvQ9Dl/OZtINhIanjskbyCAislLa98bagwhXWpY4wz1o3B+Of9ZYZlFxVRBzssXQ7aNDe2WxWr
1YFXYikbusHqkbFMRN/d8QFoKWFFdOwea6XTlvGbVMdI7X3UjxUaDmCPQ5NiWxEBX0gQcjgXt653
waN0FFB3qwGs635WbSa6c8mNG9Fu324uR0TX4GW2z2Hk1BfKeTpOOoL5hOKj02gG6YUsfgG6KXgn
kDWbgAL8T1NqLSbUsq2D1Fz8JvLH9XDmLwA715c+VRzZwurf8ACC2DDfQoqk0rylv8+4qkpet9bC
Vy8YimVzuA8exD2KH9NTDhSSfhQGSDlFhRpcOVzr0xPhxv/buaMUheqLMVebTH4s0osuckEeJvD7
NfEtW3k7xTfM4dIniNeDe+jBeyIVYM0Ip4ROzC+y6IjwOcopTqnRi66vA2XvBLkxMeG4XazsQGCb
5Zdfz1bSNyuvbqgkatzb94OaKRFp8UMx/k0sUFISaRS1z4/apuAmQ6IxSBi4QBtcAlAOejc4GORE
jzW+RPWpATkqdbZAxFUSojnr3nN6BeETVzKAbXEVvKg9hwFu+SVf8mPO+h59KbXmDg+lfCE1qy/0
LwKNGr1o6DFqtlRJeQ4ZH0gTIZZxsLR6D0nAbsk21hkI1htd2DHEQbmGpHlTHzIGlwntpdfZDTE0
dkW+FX+kI39LH1yWjJWqYYijHAwqzpvj6HlgvrjaIXT2tc5bs7erLvO8HFesopQrVbAIUY2/vy31
QqOSSzJH0L46MzOO83pU3C+xzdkr9G44gCEndsyH5bAVyIlFxQlEMMrNpFJY4uEzv1LComUokX6Q
1sbq/HtjxaGvORGXtL+Knjve6ERhSxr2p0+gzeQofS8fvoOiF4yRn0YlRZdD5paZQkMKZ/+OU674
W4AzYrNL49Nf7+QqRwTkqddM5dJefMNw2h/wgW3Lh+AOMaCvCoq/fjxObvh0HHvP4hKApVE1Ci8C
xhUB9jv/FqwTmwYqf5ndavksBJgcCtnSKZvPSKfCWEZ/O1MMwlMi8b4bFy+kPHPbeN2AMCW50XPF
I6Yx+Fg0dlrk5kYDiSjdKQAxmdWYhB6Qold14ecT1rtDh2aK8B9rp3cFBIjON/d/hfDhSJ/wUOJV
Mnwu8hQEdq2NIJwOLtfd00kYj8ntmvGa0VowF3U/GNOGKvTsIfaubF9s9+kVoVcfU6EfoAIaGQcA
efURXzAxMT3ME28+sL4MvN7vnXtsL2Li2V20nNFoEl1kE3zNDPXPM418suNigPc9Xr3BKv/SdEwH
wbpt7CvST0+n1f31K66e/c3kEsxELXr6xD/YS4UUaad8cRN5qe9JAOobnL2j7609vCV7y8ab7Z1O
GP4321JP9AqihC58pwk70jG5t7Vt1KvPBNRmC3AAxYqP8ZTr+Z71uUVxkBbUAXg/2/uleLMYVwn6
5CUPhpT4kOehpop9WTU9a6kLrLa5IWE782pdz0wcflXtPPbE6Fzd76SxVga5kW/pfC2lNHE1Ax8B
jYOelzksuYXBqawFXf6OZhWJsXOhty7Ru/vNhzw4+CjYhx6lYg770ncFW58WTDJ3FPm2CL3K2YPA
3dHwHQ/betipTKqfNYqMbss5Gatk2cuE9urrn2swiJZL2xyQTIEO6l6A6c1UrzOFhrK0gi7z+Vj7
oOCZGoJXwFMfdU0CLyf22ARImOD2T0sHp1IgN5/pTSE/y0/5ZC33JOWGHP1q23xRAEkIGsCjIA1L
coTcZBqgtEMouxSCKKEQJiP6H0rqpCnt0IlusPv5eqGnV5HKyPFsyT3oId+RRN54/PxZ9Lc5uSmk
fmLsqIQV2bmXVCmiskTqEUpCjxR6Ca3mDouWRtAT+o0qfh99VViRmslAxa+LvLvUNFDp/yMduBHf
qUCAFA+LnjHfYmURt8mF/f8PlsHu3TzDXPDkQZXhp3885mjCBB9VVJ+EX4255vjIVO6oVEcfRGx3
T2H3oOWEASabHUJAkrYPn2zEr5uN9GtcA7ki1kE5+sImZlMXMwUsy9boBWLrE+DNP7FNI9Lkg6FT
Cg+bzPBK6Nv6ICrD0UGKACN+0o7iyUDyT+2hIv9v/4SHZU54v40QQgDpwLFCt9z+TuIqXzh5W88P
X3iZui4iUZF436cJguJYPB9u+3MT1C7MBkzaPnBNTQ/Ouk5AH4oaeTqHHLVW3K+Cpf2FxIjqmMDC
fnbiFcmP3IFmfyMXYHILRTmSGaux3NKKJk0EWpS0HU3A0luDyvN3CchT3NzbHjIghlOZDsIbBWuO
NQYNtmgCSxhwr1ywXu8OfV+Wa5Wai0AmFVq0+kN1Zc4tusDQlc89ucMz1rNKWTk/sx0ZyRZwbyyG
AJbp55d1NOn1SIGvX67cQ+yiVSzmEFxxJ61XL8aXq5hF10DrRDRU5KYaav9ZwRFNrnbkw2x7+U85
hQbZbjhOFkZt+yVaw1AQZVgtvpx247sy8cSasNSGa1ngUqQRcN+XQjjJadZiJxN5K8H8Nau77tZU
DDQkyXXc8LiolP0CrKDjA5zVcaHtbGNZz4+GSDC68s4XNA6cednN80SwgHVV3BFLa4/ONb5o4mNq
oVK+nRV4yKSR9IWcM0Mt2ni0mBPCpVVA+7lR16U6Jkg6aMPXg2Tjvn3jn3Z02tvlxoHo0RM5DRoB
Kll6yceTNPi5M53rXA6yTaecbwJHxHGUfNYy1XyYyobHs670JtTd6IsqEVosiW41PQAcBOIKfv9+
BD9CYw8rGNeoDUsaivWLo0DKJo8nk81qLpqTsEXCgNlzsXnxWooQF5L3WdOHugMlwVFM9Y6TC9QE
3+yAehpFd2vJKw0KK95kAPgi4Yj8n8ysl/tVFCWXPcvmAzEjeztBWVq0KkIavXxJO8qKo/ssxpFz
AZNuPTOpr/8q/+1EZBsy+7A1LZm0+Z3ZjYWMy/UEstQEhGL43jfKCzOcPis0TbuPYqKAABXPtYLu
9Dx9ft9cqJ++evpj3yOWvmrwKxneJk0lKWLEcbb4tZPGKol2MV0ma7U0Wto8Txhfc07oPEmUkMk1
Gi+R9Ty+wXXyFwReFWgTPYK0AEjM30a3CfyelbFArEQXIrml4/GS5NF8NJSYwJ1qccv60HNattX2
uWbj5UJH6Nv8XU9O1FIqrqTCv44dTlujQkI9EYyQsHrkDQFD7a2M6k0JeMRmSuWzGwv4lgYS940M
AftvXw3Hduxk9w4kfuloOVZf4I0hdMs7IlFM/IhS6364cfTkUSHxuAGcs7JDxwX4j/a0fPdBtJE1
2X3TUDjeVo24VAG4kuvkAevYY+5UFmIe4PacKQdoQK2RCFfyf8VxnBw9SOv2ktvJ+uD1VyRIfum4
zpIBymGAdSSVf61yU4AJPEaiZccCuDcvYOoOqbdWeM71wZ0TCxBK2fWDHg4HrDdNvoHp2jpgbRVR
mlL8HrcmdtviKob/Jz7anu5sfWlcgTtgwo3gyy4Hr2nYFMBmf7ZMN3hl4IBJsw90Ru7bMfWABlkF
vPw5XJGtYwXIuLHE1qwokEs46Iw5X1FoxawxBg3gSaTNL+sR5jCTz4dPX3UY0iuPhZw5KRVasGm1
O5jwVpleDVLXuzMxrKzy8/FIJxZ7H0IBEZy7I/2Tr4bv0cR2WlfoMdtOB8eLW4HW976unDg/73IP
c6Tbm4jhtKG07hKmyvUiayYmbv1rF0Ne4hB+CRH1Pzpj2/ARj2WujTS8ozPUd+DL5PyPmJ1T8tZ2
OvFzx7gCF9XoegO+nAqBB8jIpi5A8J7EJjbsDnS8XVB6HmCVZu/z3ge8nLGJaFrNzVvIU1b6N/pY
Bq2rMlOi4FnK8p1l9kI5iy1KWBnhnLStm/FdFSLvHnRcT1e4+D0ttuq8KvgKD4Zms55cP13G4qVw
C4thmlcgQRwnmT788J9J00ai8SHqUJ8fJbRbP+hT+1hyN0fQoIKYnBB9enFVknprZINRo/AI4r0S
5tMmguC7ff5PgNFFZdsPIvO3DEK24qdBIw6che2foqGP4sFkn1ND+Rm8S6pk9sJKmvF8wROhAnVf
oWK6tDZ6EDyoJqUgbADXm9C6RO05PYWwomZHzpN+mrrZSeAR2hpf3O7EK3gUZ41+N5BRMWu8KpJu
0K7yZXdRNmVh7gbhLDZyztr8blBGLkp2JoOPCsk7jVX28G7yLoucC8AYQtZSTh1cpAhyCxvug01W
8jXMgMQ6f1plkDTrrEZp8nNfNDZYLpQJ+hJ5fokLGaoN2pCI8Ye4QRZxZXoYRfQCI+K1ubnbMdad
6yH3vf9BckvD3MLyfXdDkAWdAT6OhBVHxvV/X4MlsusU2sQdxM4w0jxG8yGPkU9aXQaP9w3RTB0Q
yM0F3Mmk9dEM9ewJYg1JfC26EYPXOmBH7y8CoGg6IgOEXtb24hZZTNdmDdaSAD5fy1Uwg95EWHkK
NFIMrHXUkTea9qKNuafCW2Iu00akZS/C0JLd3O1JEvCOkp1b+DvaPKu0CLi7IRWWegXTPvxZilRH
V3aysTeZiw0yia6pKKaQLAkJenyLZAJpxxE1Ui46Pj81V0f1LuVHak5Lzn22S6gW6PSZSMlghC5A
2Fk1g0bfJopKMtgS4BvhscHWAWczqjvSTzntD8KcswlUlNxFXIXtfbMdNN7lufe8/8bp6zy8oz6v
2hXl8jvjm+Zfev2CWk4KIa9pSAoRdEqAbbBp/X1zTI5kOTsqk0p5rmrbIq5G/sCB5VigCa2apnJc
ECjY44jhSgswYrm6QiIVnjo+UV0HhdHUAAa5PLgafq9ZB3EPJuWMBr5JvAizPrnQ/ZvVTL/fsaFJ
xzFKgDLurPAHpGth5R0chopKVo/Th/IRab7YmlfcjrZlKXyIvkeRdbfysVjq31mcVHNBtq2JL7lj
OA0DCFun+aFLEQTvd52MU+8BxN9hbWV7Y9nXIwY4FLw+1fRPlioARsOLVxXnQJ2iaSS7pmuY1GJU
Wn0zVE+DEXhYl/quRzMG60V2DNTKxbNVB6ubPl5rfo23Ur6muLo7h4hsTDhF0JXssrgo0wUtyQon
mndzucPc7OCmrXTplYZs6x+PI9TgNKvkXDqZHhw5uzZlLr1BcahbaC8Wgyw/+n5OoJvh/bH4Wg0h
BclyVLWZi6AjJDdnwz9AYqWvMJQif+KuRHT93WwmC/InpETMhQB97CmjI77jMq/0ssl7d45oNBz7
c0ZmFtSUmXLGbtcVnAzwsX07pzVsdXfoy9pmYXkTDZYMPVqEKvtdv7Jot0o/L4wv53enKDErrs8m
9anw7/h46ORy0J4OicD4CfFE6rbvCzKdV9SEdaSh6SqTtC4LtJfuRrIA0gpWadQjPQVVI8RN8b9x
Z383RVyzuZfpt/jpILbkqz1p73ag4MnWg6Q/b7yrd0fSoDG7utN/WXx2zdM/i5HOmiVHheQluYUB
mRgWG35LkRzxWsfJgJsXM9Bmgo+PlP4GQ/VghDnXg8+adV1fL7UHMq1bwfEASjrTq8dY0RvMXF70
VavYwstNDGZ10mb821F+zY+2OTSJhlU7A63aS8Wi/753Dnbu6VpLnLkueXS4Imifydw+Ss81I5EN
AxHZT66mqVSIcM3UdSkXUV3YpV04M/x6rcZ56TgVBhG6YG/bW96FiSRc/1Qt0zW6U9Egpzx03MnK
ApmCw5Rnvg9n0ZbrPvs2aMvqvCTGDIVA+Vgj6jE2xj3Jc7oiB2JIPT/Zrv4Tx3tnqpFDdh6I/Pcd
jTlB496ZVn6TWb2hLYWs9wmI890Ix5cx09ejXg7eC6+VTw5qcnQp6wVAbO90th139IS+R9Z0id65
FYbtFcTeKeSSTh5hYBB9OglmRwvMwLV/PLXErX9Ttmx4c3eFhNdUnnWkD4IVzVY8BLLDMqEFQnZf
kpkxLVko7qEteTm/QMJrZvLIoLiTzPa3QLoSHqksl523WI4CmR/Ko5J7HHqSS0Rxk8TQED+VxZMF
UoETq/FJ0xvh5UCvGQJ0S9AIkZZsyl0bFGHoiXUqIueQ4FRv+YDFgiTksQLFsbiPcYspeZl0Uf6n
j1nm0lmCZkBSd+LkloyUfMjYnHfE7bAEo05SRU0uREv8rnkprip4EANDIAYAK8NSW2xHQ68Cl6hE
tngg1KCjy8ynunnCeRYduP4XbcWEiAVrFPZ59cVJyOTfOSMxUvJ51i7lGYcb+AVhkt/kyWjgZTGv
+7AKBgtwLHfL0aUyYbB6HLVO5EzfsVW8ufGrCy2IDN1NAopYmI14v0Cxys3pi+83EGeEol1Py1EE
gU0YMMVcVg/XyWmWYHk7fqRa2WdVQwsOdVIjRdDyXbuWDma7WygQsXatA4BSjTSfnhWN+icKwlmw
Asc4RdjPieHjaMZ3JjAKMosgssHFWMUdsY9x72TcjStlTbaQA4QXRFmitAEbekpa1Uktemf2FqbB
3wl7OEtzwdsacsYbVOK5nmdYfD+LcpiihdE1gultdowC/SuPAuEgIRmnVfZUOoI68728jPd8twp9
0s/7IzFlIXVXiifdDZVDnrmh9MbhhjNQUvY+J/oXcKQhGxld+WuYHkhrOlmzJAQtWxvA2TExXYzG
tGNBh6gTwAQkRQIreltRkXYAJ7UdrqQuNO9eIZXSmB4n0Azo6qG0lapKRndtAFhE5P8SPCgYTzv1
Fvp7HUVDSIgIM9umyikHbTtwO48PwLBlN2GhCcNfJw8f9i13MNgxsSqSOvmwgXxEvw+7ug2Wvbgm
DP3uFhT54OjeX7p386mmAQ0AIerFRS29wLxeKbmv91kPb45yTEcVLkTExKvJd3Kp9DcevTYJI81t
TR9ahZE6DJQkG5Ow2TD3Qf5MfXan710cMzsJ4fIyckwhUWbd7v+kbuS3Dirgw6cvX5IJeS7wIwGR
cQjgNVJwK+fiQI9+jFED2yVW4mhD/gOpZCCkN8h8o1YuOOjLtcrmtrNSLmffN/WqzSXeHqbNR76B
C1wrj0g/ZqSL/+BRxoDoWlUPefRErAWYClwT74s5cx0ij4N1JU0vIWiJbIyt4En2g0MoortmBSWJ
LwO9fgU/kN0J2kw26LLh1Hq6sV5CYF/EnI9EaXYq4LytVjquTI26SiA/esMe937Z4KPVj5xcS3pa
Eha5+aUqOQqJqY2J1pu5HPdaIJCiEwwEihZTDdt7U+R/syb2YeHniKCscrUQbQpN6nbi/XXTUCwG
pnkMwmnTlYCH8E+K63OHK9rFP1jFtXGO4/bBPzogCyfKUrwWz9zezdUsq7S5BzrgdTfS2slZSeAV
ZbOtHUVj1jCYrgSNBElRC7XAgZmV4U3/yJSaOScZ2I9OCB9AAx0JhjC9UXOaxM8/d3DCXdbnqB61
kCLxKi0P20qQ0VN/DRQ0zy+b6XCvlkfzUV0qaMIbIo9hCIX7VjBhGYDnX2FQN32flY1Rpk19WY7W
c7kQ6I+edtVvtFQ9mFap4NqmyQFiQ1xAJ/QhibK00J55bnFA/dmc08U2Cit1uqtUYeC8QKpYXeen
7RKMcn6O0rb27PNZme55MI7mZsOm9sDp8zeJiwv0hV9mCjPrq4fIN9tMilqKmohaTYcqygJCu1IZ
QqNoUbyoW+2wLQsU9s5y+4fazs9PqZwvOHzSIF9JtvflcD0dP3QcdqXICp0bydfqyEshcEqqy3iK
cwJJAN327R0Yurp6k9k1or1aaQSNpIeugRauIzBVAa1mb5TN9nSoeuO+BDaYo1qfBhmZ80Znwyew
hWetuGLkNoguUULnv0GtO+ByYBfkcxVBBUIAF5KV/TkN60f8bIR0ielv4Ekj4gomOmRVOucMqxjX
WvBCoBHekSAmdRIxviRJup/LPkEJRRVNVoE2Y6jYIGD15dAdHZdjY407SE6cxcplVQYaNoOP4dX2
DiKpwFsqPzrnDeOUlllMN02R/vSCiAmSThlgOz7KLF/0k6n11ZDxlrHs8s7gbeIv269bxE5cAYEi
W5lpE/kQzZXryse5Vxv8odxnX+pF2Ma+30wsrvmVkVs6sDSvpjRj0tIxex31eaQ4wQNwfi3wZgxo
0MphIB1GOM7X6gcOqeGVLbRtRyN4gnN5S+3AqAMcw8DQNVrBbPUenPQuyStq3Pud9ebsQ2Vs6f41
6i7pJbfw3evk49AFB4XPSkNOFfErhAzCiIn47yfBtCpPCzCnftfFHpuW2m6iuiuy7I8gChMFWJbY
VUxoSORI5X3siYThnuo4KJFZOTeCIgwZsisByVgdLnVplmiYA5pfD+CTwDEfojw9zQ1Nrv7WiXja
0TMdUaeIyQakxMqeJNUrewbkYw4KsFHuN/saA2X5mrQrhyJoQsS2gbtnqfxDGLrvMnhxn7tJaGWh
9lq7k7cQFCJehUnupp9AWly81hnilhAzjQLTo+VrhQnHQWAoRDkHfqc9T8xwtqC13GyccRPf0h7F
Y1xPzSxS3FhdJacPIS+fMJdk6Jo0RCsmBJedE5c5i+SDmrqKltO4tp73XVCDpZdxX6FxlLDHwUki
S9j4cthriiLRVwe4ueDaZy4DUrYoXFNrCIxdYDkje//ZaljryR3BAY4Yh9kNa1UtYXwr8Boj/L1H
sgIdgGGZLCxSPRmDuRQjYqTB+/F6Z8tKBR8uanyH+wcuu4LEM4Uzry1TtgLoCUoMuLAHOTCwo01u
Nmc8O/NEjxFAXOkzzXYsocWrpE9sIgUcAjwLEKQT+5YrYxLRRgu9+Zf7n34zGoVgJtLiNOp3ut7a
JleFS0gfq/6YtPd6WluDXLYZ+sM1HnvWivt67P7nhFcjZO8fyNN65N/8YF5eYQ6ivSxM9yIZmmTE
lbaQhogDsPFQWlQd5ldLr8KRNGF1CtqjrwPtJM0hToI5/IbFzoQiJXFwLP1ffSUwlJer0h40Dn0s
bLAjNsWktZwDScxiB2tTwhnkFpbGyj4WjrpbhcRXBz9jBuQEHmiogx6CYXj/K7ZvokYPYcPegyJ2
SDkjv0uflCrNrr8TFCNKYqUxwnAPuAt7pO/NwELM0Zt0zynT+uYzD615DoyF2xtvZt0IYrGXkOKB
jgXGKxcCTcyGSNVG8MGqptIp2DOkYP6FTTmD7GiUKRrSZ7ljAnSVR7wAnhLWB1HrBNTtOGReb4+w
BKNQMYGorxdn8XwW1Pmx99RTWP9cAbeeB9DAVKK5Y5i15gWfkLEmMtPohSnkpeXvtv9LtVL68aRQ
qkNDgpEAtjnIiNilul/1RkCqPJ244bS9D25upS/6ClKtbwQTj4Uy82bVbWA4zjhf5/uHYZl+b0wS
hb+8E1UuvXL9Wu+26Ev0pX1H/U6P0RjTSjTdihcLymZnqWCOMM09eTqdAvxpdZ2UMYjUbjI3DYjd
GfCGSoFzQYP00TOs7ecEkW2Yaw0l1R3EyJmukuYGaLFWtXGX4pRv3MZ9h6dvsAksgV+xkaH5M9pw
WPv2vio7yOQd6zFL5BRxoLPWGbISMLPZfKN4rGdqCUkTuvmGjAqlERF8WbeDeOrGTSxxfbgahApT
zJ9rrucHtgj8Y9j2n3Kx9NCuPDlgLXoL6WfglcePVOzCJGnGat2Ky8/k3Giv9Nn203RkubVquVQp
IUrhs4E3tycB91c+VSO4oIrGg4cwAzONXWdkIZAYqeh49w9bfs0E2BdqwlVOJIy+oHSi+eucfWSu
LS2dozfH0V5ZnwvpEYnhqVJLiJHuZ/MT2y0hugO/LwgYWXCmJWj+cKXWifmz120loqS+Ftgzyn9M
diJHf1hnQi07e/BzwIFj7S1iddXQovp453Zko6gHim6QofdmUxsfT3hc9Qo0vGtuQsBuj8wQ+8ul
wbwWJ4sjJ1yKoDSJoP1k+xjOKNZwXlG5oL93GMJtUP+n/FoyqP4E6ZZDxSjXHvp4XYvZ3R/jLWNw
34Jri1UH+S6ub4DTvxEUylQL3mAHdduyhfHpvvcuzHOcED2xKXCDdPkdWu7KDN0jtR2T0waDrzBr
Lm54FrJYN71rK94RtEjT0mZ7UlCxdNbNMULXsJGvwrprsEhsk33ZOikGFubGZhCb+vl2x69bWuia
Yfv8TmbEVsS0lPhuHxSBpFuz+3mXkzEpM2G9DCnIbr+JAlm3LOj3FcqphuKTSxv5eawJbAWqBWmW
riTImrMcshurec2l1GQNSiF/19AjiKBws6koQozzL2UabCsIPc0BRRLDXnsJXSURJCCeWvbSoHeJ
o/PbUfbdkpWYWU9owqbl2HKocAmonqxSBEvEsfwm7x8tH5ia8Ns82sxQONKhZ9vRKugPyqX6bLbA
6PkXCoTYlD/EkF3ZWDAj4j4ttYuTqYBQ7hvtcbdsY1AdqdRcvjmmt8n79BUHc1uaw5YjkfgnVW9Q
+amm+aNZ6QE/bZKgKuiyl41Te9ClFSrqQr6kMI8EqD+p2BKEeXkFQCfTfzKEREddE815MICY0NcL
qKaw+DKoqkTDvFLWz/s6sUTJ3B+vhfrcE/9Z6Xp0fAOLvtAkAUM3NJay7ZbTTkiBoYioJNxYbSS7
qTDu8DYG9RaQkKamYDcKi78ZCBr9Ua/TqY0rZIIvawKU6BHdt4TY9IL0IDT5GMHhA2YtY+nCoJ8u
HzG0Mod+C5+FwLcyzkiL6aMNj0lF2TSc7fLmaUDKW4UZQsdnBydXw/Vw6rS5p1WGVlEpo3R/QAgu
LYEZHvF8XT/E32Tw1InlX7k31J2ZazJTghdOx7G10trCAnOS88B85DFdmb3m7wG2nVLtKxCFwQz3
gHAcEAS9cvOgzjoTDWj3rutuFGlO/3mRPVuxqshRInVIHMFAnOcjrm5bqnsUqK0SgnruLyvXmyl3
zCkwMXEZiTWtEgDaqSxk7A2bfQEV/2Mqr2PRxlOC+HJWngbvU63fMWEv7eKJ2KexgwHP91Jm4G2w
gYMEUL46llpNtBpYjE9ETupxRgfqkDjqOSbv0QKn+96d/wenwLbMn7lBbV+UZE/JCLYe8xbv34up
1RitdtQgzhw42pblcMDyxkvRm44TcAvrU4j8H/Owj7deWVUUqlj4lApc3PlW5umSsIG654HiKAYl
jl5357sUpRwgzXCyqgjSNf9HDoXiD8q6fTV98uCYW+t7uhL9NQNHL+AuH8Fgq3xUHWQdcjMbFKf3
hFn4YQ6Lp2d16abJ9mqq+pt07JuQZ4X9nvVQSIz5X3pwgnA2jC9BPYSSdHC0H6vL42yM7rs4Dc8q
TDeDGzrf4iL2dB3vAkh6R32bmnfqf18wuYUJkYp44jv8VVBCXGEHggHaWtvsroutmiXl0XQLp54F
f0+X5o614lOJh21MQxOf2JoXe5Wm+QN7BdXshgjSJIQ5khyWXGM0/WxahetVHng/MDI9nq0gxTL+
3Ee/mUgJN2qTN4e1QeIaO0o6q9D+txifa6oJiGtpRY+LpqKk6D8yYLEpeyDbRKNucvRkhJ1t+BvV
WFmgj2kFODHxO9BFUTVNL4jnpno2/L69Jz5YgTaNWlYdg3OdxlZXChsGUZcbOiwovFDX2L1IMvSh
/c9dQRm5P9FYEGCiV6NfW0QDfFwvEY3aRioIFBqUXjXWOTMrWDyxFsxDFhm1TeqyOZ/CIUQtNCBR
M9hmYGA+J6JW0/fEt7/xgqElP4GM/VUGhy7vyVPkkHRPWjx8yGimEgsf/gcsYELYCWeyFisuk3Eq
+EiLueEj/i/HJ3GnmZ1hS4ot2zzJAW4/BqMMNKONMLtuK6mfUXmJ2+2uhSZtbyWgUlDaL7S4l07i
WUZ4e9QGL6M97koJ3BooMmxXZTsYNsPdq/GAQJPaGVOd19U+FKnAVtnsgYLweoQH2tFeA1nqJ6XN
kKiRG/nGJXhruvvoat6GGqgEUevCnYOwDFpLxGILVsj4sXS5Njmpc6/AENRp79QWoT/iL5q3RX0r
mQvsWx6Xc5gV9wc5MrSCFi6apPnjDC4Tt8/z//yxaNxCKsD4m8VCvd0yt/RWN2q4JQ4bBXIzy9Pd
HJ942uxZEUKA8LqcAzLIWzkWI+0txG5onS9+uyZJ9LBiAjMRayZy9ENpOSDv6wabOE3jNBWwqnJP
Mc6u6rZQLt9VO4zjw7ElVqKkf3cUvzgFqJORm4Cc2pno80DxlkD6fblUKUzgPFmpT0BLjVDgxnu3
G7PRJVfb39JQKhWFPvAZ3UvT6MYUbgFDKAmMLYcWaUm/7us8CLqnMLIuhsERy34OodoGIri8Ctr8
mk3/P/7btYcxliCRgPazQhsrrJhDZbL34PxYKKyLZooTzLjVjg36jqflCofmkQHmDCuo9Z3TMxHE
Wgrl5TomZD38ADoeFP1x4/rO0vX57mhUBWY2B9/aJ8W09c8r8YOM7bZK89Om+duk+cX1E+FWitJf
qFVWHxOAnGN9jfZ74pkpM9oOaoHz9Zs96KkTUSC+lgXZ+Afg6FWrKsMU4chhzvbUd0g2qDxaX3o+
iYo81OEqv8/A0T+MWOFqnh2XLbgEpO0V/5LBLgh15d8GCDVVXIYv127xEFWFMHJoLsCTBHJPajJH
hbZgADojMjJccdpUypfPgh+CrCCNzu+Ug7dGlPaKZO1U6ZpyzIpzIMFpDuT0cEnpwjznBrwjGIGF
UPtq2bvKuHut0xrS+WDyJpcMLblGkb5uzjIbiVs5ghCzyZ443iptfiBo/dw38WbiYZfKzRXWDZae
ywL48mEOZh3iAA5BaVFy4jFIyv4XxMzskJcGH6eTEBaWqq2ZjD56i/rvpyTXKgh+mIeI72kqG2k7
TNMGUS7lz1clt11xUlYTB2ATKvlUgbVXJRnYAsuxFx+G6FEw3T76eo/xzei8QuI3HL3MXJhug82h
8Ej50/3fDFHxNjQ1QR8cJIFvWWslNd/uKqloUEuvOlTEwN3dfEuhocmAJ3U6mf8yk8VXoE9kFejd
MnJyzKuFVq3ZvSdcpQMgXKOELnhnnNWNEyBYVoQaljyYmhAPu67vRE2IX8IBBw2iOn6b7Xk+sN7y
SmpoZS9Sw16n487G6hVlcRhNDZdtD9GeU3sqPbwsPQnLOxjrY52OIYLKDUfZcWZLdfflERcY/fOA
nzdQAT4GH5VRlsklHtjjb9AdOu6XCl4y6Fj/ZySk611+dg0c4UL6GHNooaBrNU58FDcyqa/2/X1y
CUvVRaDHPFs61QnCnU8qfx/XXmHpB0vHcHzIpiqRhj4Qpczljkrdwm2hLLmh0XFJyhzRWEWOrVLT
1cbnpqdOkXM4eHH64izWc5zlAIQHv71AONA3VONbqwS23BqgbbmrnP0LdzoaqIFY6vDtyWrxKLgZ
QhVnTYurEsNE/fd66DSHu8IAbOgtpAE/TWpBYb6exU1zjwyHPhPgfdxnixRGSVfgQwwIaNNx5LI6
uSuJrUdor/EHWJXpOHgY2Vv9fHnaBZXFm0Kc4yXpw9Xdw2iXDKniqpmRERkSXHwoHhqZrBQyVCXb
aOIkuiYvjCJsManjrX2XbTI3VYBul928na4ZcQa9LuwrE8J9BJ3x8/SvXVVW/fFhF7XeXvPUAEYn
bROpvbwELlcf91z7qSA5AXvCt+B6+IK+I5QJlTqRP4I3tQUkWWw1gNvk24O+5pHjayBwPdveRWZI
OSU6Uv5EyK4tlMKrauHHIQ6ssmhUu6nQ4M0z023F8fWRPEf+aJRpABzcwcnwdTQwtNyiXgILDYVq
+HgUo/DWmU2QhSdEiay3UkjIXMib8DDWlytFhlRthsjrzykoWTh7fH5+XgI/z5i6E8EQtWldxCuK
0Bvxcu615DKMR8Xrpn48tCGY1j2jO0b9yYzXi0k6WmbGjr8Sox7FgPL/76jxZSQHyrHZGgbIymMY
tSEE6zULgEBB5/y+mZdvXdnmzXplTAQEtyNQlZXoFP7F7YnPbY+If2rZgBtHH6C3LSVUqf2isgd7
AahpMnbNUQ2Dza5+ccfZmP/Yqqv1Uw5got0YDHZXb+q4D57SpGfOmF3nNEoK3hJDzWaUeDqHCD1a
fiCJCNCfZ8ZgEIq1woIgUZcrKK14asN5sLAy5r28wO7RKFte5UjWOh3RQK+mtOVlnsWASF4GXOFi
mM69qywNcH8iA9eNx9j60Lr51lKImB5kNbqUS2wRAifmxd2OFgTLOFtz3zr69UwYi9q161NMaGjb
2SlQLi+MAmfJMIodcIl/XOylUtWyg4zDPAVVClnBw/J1l34QsavOv2vCDQExdNpjxGxDosvMlsC2
cSZ+lJ0+ShYEqAGmSNa57Xsk69k+eKQharZTs2i0G7exi9ILtooFqkU3kwiFxMSBHij4b+UTiefo
t7Pq6e+pAp6+jVBWWZAQHaqk1FMjcFEjEgDQlU59tjrom65LfdCub2+C3nwTY9KCKnWa9o5MQ1qQ
c8CR9nCwnPKhFG05mvI96IguHF+3nDPrweuWvOAKS8MeVInnFiLISWASACE2lOM82jm/NEnXC1YH
IT53nuyR+YUZefmDqDYm4tPt78yGLuxToEZpT42X9wDTRjRSbAOqDC/KCCRxM+VRhocBzRlIeFvR
dDeW0pP+5Jpb2u5shwutfY+frFAusdKsq5Lrv5/ooqG/TrSfSudplP6uRApGM3uXiWMm3wH/dAvk
LwDi7CxoMui3rt3BmzgnyGG6oZRxRdgmz/RfWM62OwvrLYodA9zV3dkAW3p04ITQnlOYHPKwPNyL
Ra+kBNcHyqog47KEgDNdeFvRWI+SIzFAI34FONh7CXmZsRcZ8VVeXDwP8Tn0TiC9GzGbS5a8e/Pt
eyx8GWWI3FtYJ+hhTM0arSq3kDr7nXMFppC0LGaVt0HFsURLLFRxcmrGyqQdrTsZ5tB3pPnaXPIo
l5Hk823OybzDP+6DtSkID4kauWvQa/PJ08lf2mHK+V8TuuZ8bwug+3HoUhoRGxoxrkS1A+LEzBA3
jEt/BUraAt/6K8Ay5FKD5UKFE+PLc2r7dLb5VrLR8N6wHgSksJahtdLI6Vh92epgg6y4ILMBF+m6
sdB4/juA/fCte6k0wKo0eIrXeZl+/UlaAjJHI8q379BJN0NfbVdx1crIqzvj3nRs567Jg0PxkXJ5
j15YDBi+TIaHLslCoU8JUkOjv2gGLgNBktih1vTkLoLP4UEf18A0R+Lk4kDqdBi18rA3EkOJ+5Bx
OtrsDcgRknG2WrCP3qzplF27myojOuvBnmF2sfqirAJznbjma2Q5PeQ59AtyHfkBS9T65goTkIUk
H1/7ItKkWqA25lm8EmY07N1SJYxjUTRARlNkGuo37NWTQQVbZ9327TY68MhAwh+M3rRt94ndiCA9
g0V/2oYn8DgiSKfovjdncKyR9XRACE8KyEG6wcr/LUCTbROaa3AUBnnIe42HG5Gd8Anb3A/Kdryo
bkcPDbeSSUOOeppZ1n5vLy/CUVqHQgZhJv7pluQURxOZ6qkQuVSSD+/N4Fq8tSF5VIz1F6RIihxj
XkH9JUlGAnpO3z5SiySqiw1M5yNfYx/Yjc3DYPZPxB8nHagV4tuIbscRofwVPZKmpPwDMRAEx2lA
MBbXio2w/7wBoW5aRti6gNpwC+0f/E4reH6E8d2MzcPT9HldUysgCtuoxKOipB5WC9J5/47BAEHl
Y922nOe1hVti0k/dQkfJQraAPin5nj2A49uZ0Wj5uVFBy7Is8dIfvJh01x6v4hApw2EL9kSIEsjo
j2oT24kBwF1Q3kBcyhhFQoPSDpX+5koamH9Imwm/MARg0Kis9iGjBrrMsJNuKCERcy4NE8UJgGiy
feCsfRmxDbHeZjtzwpsojs5Fjl7rsgSTtJwZXgIz1RRFrePviiiB5pWAqteTGWvKWogk2XVAvId6
vUrx+Z/C/fA/ksTt30IxfXuPkuwnoKPj+Ej/K7wdTmZ4OoRaPGycodTYz0cnwh7D2YyG7DOAtMaq
7dJKi9TVjglE7aXdJ4gIcz+iovzrGQyp4C9Zy/mtmo2HhYDfjLMpM9Fb6QorngzVSSbAGYX4FjCN
IdJbaIsrtPW2D7gdd8dpBoS3P6aO+QI8+3lpV6x3BaX36LIjoBcauHUxF4jzllyETc0yGxkfpX/6
XU6P0Jhj61sC7/wTUhwd39HG6ZIAjzO3/bMC7ELfL9z1yxIlFai1z0xgKwcXghWaSfLpGNk2CVAF
Xm489+gZTxMCqrkJPrKm0+OKtFYyWPrg9pUzphBN3wqwP7YjrqZDe3SyGUT1iTekVhSYUyy8pTYu
OsvLaG628tBawONIzAd/8ZRajaJUyYpOm9GNT9Wm6Dg6Ql5OwX50owT7fb+TnJyGHaYethIcVWQV
hX2aSUakAu2H1tJIGpMKkGKi7KasPEPV+YAFOg0CJcJc0bNIwdxJB6mK8k0mRCGTufR37sxJVCRC
S5Rd8uqGIyKEcYt8c1uDlqU6RpagIKuaxD/7XfbPFD33ygBkjHgMUCMy5Np0ALtMCZpNOUcVLVW1
fgPYcE7HhqVDw2mVftPelBHbmsvXw0yC1pwDFfLtHvI178wwCFYkTwD5b9AKPEbbVkGdathZPdim
/73FPFFOBZbjvjAKo4uyZFOK8dOCW1w07/pLlQew8LkwyzpVNyziPX9dsWEBI7McXODLGs824DKv
aR0Uo/H/5b/JxNeLVGVQyQ4DMrwacB3zN3i3OqIp+XR+BJq3uRC5kcgTUSGn6FHx3nUk3NBjDNHY
eNVZtR5aNB70dVY4kSIWhOz4IZdojh9wpPrHLhyhRRMSX0zMbLugbPKFJh+sMUfqhp0iU1zTqsV3
QIhaJOIFhJeQ2XkIVVG/r8B1vZcA96QNXzkq1nUvtjC+3xglvOESEf0DzalCzKO35oC9mO1AWpAn
48LxOtjZimHJzUEAR2v68DzRGgfG/FSmli8Du8t5bptgsKiBhmiWm5Meof+VYCKhpLOjQ5oJfejs
t0SfK1Ll3TEu5A+e8cqFjhjaTBFIJG5sdMfytLW7O3cfIELXjH792tpLQJloq16pu0XIDYMVUcLP
zJjXrAbgk0BUtt8FGqrlAi2X1puVcT9Cx2QG/fYl+f1+YnLfFmq1brbjc4vP9m6tcr8oMVNBg5wz
vevFAD7b6Tts5I7SUKtA7Ujq1utaqpVQ5NJt8xnkYa0N6z1kmWvB0wT/FyzzvXiK3AQnBcTvO1W/
neyONCv5e26iNfuPWlE0LA7Q7KuPdHyLnAemftCIDkUulTPQ2135BeFDboJWO+KOUdC0K6Cd+FFr
2Ex0VxKGv51UxYjK0vFd1bPQcQF2O/KQ7HnVq00ZN4S0GL8P5uJmVdACHejf2xchuzMTTSMo2CPU
bMw1pqicvp25ObjbZUvq0zEmEy6vsxUEJL4RpXzNol759VP+18dwr23Ef6V2PYeJ2XlMYRq3FhdF
8Y34GzdDigjxD7lRNHj1DBsjDFn7etf8jheNi2ArKF8b0bHyhEGzDG9elyQ/m4FQOz3xdedVN6jF
3ApbhQ6dQAng2bTpN9Z4InB0JzvoEjjhSuhl/cIu2QU1hYEorLq1mAiZGqVFIsD5rsddqfS2Qmin
1dzX+SKaESsASNHFwER7KNtura9Z/nV+qdEjGxElVwCdc2hnGzSFkkgG5314z5WvK7HcaFp/offd
fUIaD8PQM3+mpyXOEAWR72lJXe7RIcmnoRhivwVMPHyt53s/mUmyIgz4CLTLvWhPrdA/ZdVgDkxc
iL98rPpzgJ24iEFagXwy7NK/+flVJ+tejwXxpRtvTTZ1dclJPw6RfsnYB256KghXhQdLOqGe+5yN
Gh4WrwrjaoILk3oBPfu2J1fh3cF4iDKhmv4v3ob8+ebYB3gxYfwTHDiz2zw883hs2BNwlzS9k6p+
wxjJwGGhscrA2FUtiE8zaLJwdjFhjF541Xx0Q7dnbdIQW6hR+txReX1FcNxbYwsS+uldF/QL6bLr
vxda/aMo5GjXAkWZyFrYVaONACiVinhPkGbhQ5wMZ18ED7mA5LKenPRFD6aYQRPdLMzKquNEZzD8
26D74AmGbiHVEOOx3GVynP5ph9UkCoXfBGTmE9IRHGtpwHOkaj9XxK3geXoEMzOPYdFzJDe3OcPm
kUF74iIn1ViSFE42C+NHZPjxlnPQEsXO3pXVKc7f55B1spOvyWxlMzROWbcIVcBMrRxIStVRfioi
tVuF9pDOJ5eZ/31KRDjGRd345i9dmTIxvPBvMJzDm/LMKOVMwzQvydFPnD7SMH54L8SdRVP2MEjC
TySuFPfoBGkfO80YRdv02gAA7FaN8VlF93+ghfV8Q9lv8hdNiACeFn6TKvTzVs9qLUzyc0btPtex
3HBOzuZZsLWn+vxs9BzTHI1NbRghZQw3qdFa/X5NaA/CPGVcCS9LMcbjLd1eCtaw2AuiYidtxL6c
epKHXFbDRcPLrnLKyoN38mYNyLL82Y+wDlnKLrwrte5hMrmrlC+2saWbliPJLvwz0zBvZGKX4Wj6
/tf2N/M3k7E05dW94gXm4bgUmI2/g9vx3gyRAMZZUTb0kxnBffAUhKob3uCnBzzhkQBblsaPo8zc
31BQB+z1Ldov+fpQyldibpSec7YB9XiLUTkQpkpVT56GxfL5iq90XOXMmHZc8LSkyxrSuta+5GL1
wQL8g3mU+JIZPWkmAbZpcrwzZIRoZd8SbE0lcLgPFsZZEGGmzt9AUZn0OGo4Bbyo77/JEtMhUD+5
2tU+IYr/EOZCiWuDwreVyTGKn2nzTEo9O688wPwJiVb7wnTJ908TlsHatnd0vlQtMC/Av01s4Uqg
aoecjKFmkbLQtgo4lwM2GW+tTO06m/KbL6PHFa0jccmdWPaQNA71Zjfp4mmIZERIDg8KgtgLsUPN
5JZSEW9L1lAiYuX2ffarMJba2GzykGPV43XkOOxl9BSb8dFLpN0v7AF+dhBHUEeNn8jHGBT3CY+a
l9Uvts1mZNSDA3GW8Z6IUfbHM16dqOjqKbMvo1rZ+fkZZig0b8eZdj2+wp27o79XMPffkTQZFwIg
cGL12K710/VKqQHd1zJRWvYb8yTkc8gb9UNOZpTgKAo/bdooPJbsJImV6zZ5ji3mIPmcXQRmKqmV
ruji7AFWJKlfUcnSnKoYiKGUQtmVopImtdkEjzRJMdcsJaAEqS5H07y9HkTpaplUHNK+gJV5FP0o
lzTSG5eAECWbf0aRdxbWOhuoSELkOn4k1AM9vuqT5DW6yEzu5dN476xOil8bKlER663RdKIUfUmF
zIvQCGC8UE/t9P6Pa7RD1WewuRXfdfLqERG12uRTHqDfLexf6Tjc/3Bu2h4t5gTROKdK+6fhzI+h
sW/HwIz+AtsnSyGzalTxB2OSGjj/RjBmSg2kCIYqm/li0APRxsBilqeNhFa0ME3HVAaJ0wfRN026
bak3/dISb2wEYdtnhd3BDj3teRVsloHhF8JT6RTQmau5iO4PQ73WzEu82EQkJ1KgUbepK+F34cEc
4TTILRe4rx9sUPRl2+PkenPPeZPOlPdFoP+kcMhWtV5W25odU3MgcrbB3fIuHkixFgZ8aWPI0x5H
7fbtM3b9BHzl58MTMVglqiUWx8hiuLQQmSDy1/E9CFIv2dTOIhxc6eDZYSOZsnMvNp5kTd8Ktl41
S2AQPfCkCCwn9l1WRs42ZHq8S6k91/SabE415hh+WOsInSJNWtcBIbk2/0AFVhj09hMnRueaoTuQ
H3bzAfVwY/0+BxrXBMQKS0fQl7xxujvnweShonh9Rq0xlEgzNaii4KmRsVYSjqjzXrxJrvAxAJsJ
97omogXP0du3aLDY8jjMRWym1cnhqqcsJZWBi6jBXfMr9d7/lVAZ3rMtUolr0zi0JNbPsCogTKwN
Q1NunmGbcpi4YB82HgmIOyBQjRdBR16RPl5apjhVwpQxdUHcOttsN/YUDbeF5WLnOEMNigDQRIcQ
5aFxWEREu9gbmz15UYB4WURvVXUTYXJShlcWDqtT9Vtu+Dtx8XDTE2bZwSNi0BybRb7K3RUsBl/e
eYqH+0uhprCUYvH4B+xLCgi2/sPjZN6R3BXDvUSnCmNFDY+ACDU05WfEiK2rdLQEDm6RQJUBekaJ
C+/Qlf7fFtBj0qhkFqgGbnqLMMynFZyhKwc80LF5hlTg00Zl2/p8Lk8zIsqsDoQbVDjTeTqtn9Il
go1s9Cn5KssTComy1y9ZpMpCXzM8UCYCNXXKP5LdihxTUs0UlSX4PhTI92ew7dufczIJuQxRZ/We
84jN5t61dXHV2YD/RiSsw9QbA3S+19FIiFz/djjcngGBstPGYoeFfgk1iGjTa9P7+TEL5NNdZIgr
YYOvHg2c0r4L/cItM08DX+M1AaM1Ja7gFPJmTcuSwbztuc6MTSKCXuzqE4Omvf9OHmQve8TK/j1v
FN2SEc5E6LgbOyHwIEmgNtW/IY5OhPAjgHAzw3cgxn0W0RRJgn2eFjqGqxWeFgYDXBWaRhUJLhdj
pD77I3CG2cd+3Ii8o9VTotJUNVVfPdKV2ruIIOGRIGAVtYcTGW1evrd1ZuYJ9b/UlQUVk4yGpo6t
ePJ5LY7CLqUP73P6dPgtCntlCFO81qO0yKEpkjS+yRw4YLqKUd5qoab+Ee/0sP0H2cuoYMXJ+8f4
/tUSHHXtOQbUtUf6Lp+pr6Nonhkj6ZQ/4IEdBy3gFhQI+GmpSRCYLOUThDab6Rar3EjIXYzmOx7c
Ed7LF2kfnZCFbBMvys3Mzby01SBZuZ1DqVmcEBfsXgKj2+r1/+K38kDfHJS4kx1R9GbOK431r5Df
TO4fBNi0+lmIuaVYuuKsKDpR7uzv5+36BBcEJ36mvEK33qXHjzilze27spPSZm1v4reepTrE1c7a
FGYxuwsjCqrwOWkaKmRcSh1GvedWR6iRQ/wUDfNvfVYuq8vePN+ymr/oiQjA5ApELDXTeIkdXNKG
TWZlJBBdHsh0uoR84amNSiXNKkFIWzQ2DcA/vs4srRd88BIr/5eUUWQ859NlBoH0BNBff3u0yuHF
rX31cTASdiZuyyBh8Vkqg5fiakNvRlRNJK91GjTwh5bhiCpNwK9yTpedputES/V74FNuwd/OfWxn
NkaIziPkUQf0IAbIwXp8yGdI95SOM4IHj5RlpnEzpCIKRS5EobZinIrl3k1xADWGhc/oJ0YsbQMk
5VncJ+YooqFokOYB2rSw6lhWvSMfTVGSmX35/FLQDaXVKiS6MjVOE/ljbXfTOm67H311fc2bRuB7
FjBzVUYzT05/voXzDi+x+MdAFaTIYY5PKGWlEMZ5huFaZmkYzQx+kbMA0kKuPxejYWjsdPkd/OIE
0+eVS2qI3hUVNRY7zJLasILMHGjmyvT9lnP5I8RdeNwGvw/CnFrX2NU7uErqYfh6XIrrCdlblDXn
azYQvEvXIYQ9TQYIlz9f2NCmF7x2dGQdsh0zGNPmKIpQQrC6aS4IFzyIe4XVKCv50qOubxH2NPw6
PddaKXUVvDSjbzYOcrjh600o8PY6OO6orBf9C4YLsFA15unz0lfEFQZ4OgHdCfzfrN2E8DYnbFhN
tFWd9d0pVVvUks3J0iA/BvfCRACpQx3lJ4NMlFTvhTGi9qa0MRr7eYl20rp83f0pqaq01trrlr15
vfDrQOgJbc/Rw1rwOiThHDp38/CuXDhiZ+P4Pbz/NLjMdeDwVk+rSuqucIZEtex2cxUortKqSsfE
U16FV2w0SZ3n9Yzoe/SLv/iWFbuiFZYbZgoSGnap8EV2J15iptaoQnNjjlVzQDOrc/5ktsKfrzpQ
gne0gdTC8OiFfbJm4imQ5/w/daGw3Trcy8OU9tqYXk3OWBP85C8Yu+x3J2Uoq7QVLAPMAb1gO9Fo
/7sHB6iVeG+T8TSChFxpOuN5Pp+UjsQQhISgyz1SDJOzod90UWm1u32c+kt/mXPYMLjnkLg9Gbvt
LXhqYxiA48jItY7UsDoFkrh4aqcmehxBQBs8shwQo/eG3QVuS9SctH9WoN7XwlvD8QM0Jt2YK514
DojsnPqPYw5xNh2qqrBv3jANJxqg6conGsxBeF7lcu70g0tHkdvbmndVx8rGvbyy9hoXjzfGWf0O
szpF1K/Ph6mWLCc5OoLnm4EH0b+j1S6+f9K4ZazFSCCK0upk7UX7S9kVx73RVeZtKcGebBRllaFw
c3XeWkORGFyFwoxPlWjLfqdmJ3Ufo2mWYAn+IvhT6qN6/MiLIX8cxciU9WSjJH3lyzfH8AlDa4+d
6S80ZyZooLiuzlMTGhUqxk0tmmtfA5j+V6TSJwbqUChy4c7LXKqEO4aqvaxL/QWTQiUW4K0DLGxa
7RQxrFcjQQr7LG4Woj9fxS6UJignOjQGb2f4QBomNgH1mVVqMxzgtgJG/E7bh9VRZfAINfgDWD2G
zHiyzwhtmXjDkFIZjYpEZWBp+VvtDe+KDNFJTltJT1bSCj9azx5isHjhyF0upk4on1LGRDWi+HOl
4+MJhjpP9ZsvWyrLcuxIBjcFDybqfT08eB/i8vDprW+0JfoqTGcpsxdfYvVfbxPPODjSiDeCrzvW
TsmSNyvY/c1HVOcMTQGcYoz2LF2zG8WADzzGeRh7KZHLYH24AGaWKOZCn6gxPy7wOj1E40UjdBca
jmZX5nsvKRDZfj9qLeUHRfCNDLcLuo8uCP76VGBu6dz1EUfqIZjt/bW0UkBlZepp422uzJ255eda
Mt0an6OOdFux5RUJQdpIuLYrrEQKOhMocQrkjlX/SApbca/UZZqpNOJZSJ5+m7JU01p4iq9HjAd+
qJX+I7jatmhZ6hpOd1VInXNKhMMEl+jDUd1ZxBOUEb4V5o7P068XlsGGweuvIuM0sRGXOdc3wdH/
0FwMWJVs31W1Bz8pmh+8fgRvagvrTuAL1v2+IWgAtF/NJ+R2+iLnP0CLlS6OJkhVrgjbqYlZsSOd
vrvWcd4P6OYIe0RF3EMaHBj34psUdUtYJZ/7RPE9G7U9I6FCN8QVwi3nUILRi8NUVA5JSW53dOxH
36SWMnfAu3a1YtTBL75vwzRkIGLKeD43GkuPKhwfjlxiK6EM1l+WaSXtKk0TOtRetKVMB0Eo0Kxh
kkf899YG1F3GXtckKwUinIK04KbML/B6H0kUzhqsL2rQt283rWobGCEB7SBR4ZZffZK01hDOF88i
JxGJ7UWQ0ZBz8tOn5yEjRo70yf6SF9yxW2NdmHRx+XvsM5njRSnfTO1lOn1anJRB8Ft0JDPMLL4+
CEziqf47L4jRo9K24do9ewIShoy8l168hu14rVuteUGbtsWJowcaz/37J7tlNRykwVZnCOoejW/W
kk5vPxFI2UZW0VpJPvi/7UkBL3Jq+ViyVqjWrchW1Yh7MMBN/bk3pd3+R21U6i3qhc0f3I5QS87+
cCJQYowd46i5wau1OnaCrroKLxHDgeUzp9ntiZeDWrwfd7lG4GDpSY1vtr0d3mNNGcGh7434AzcJ
k8hLzh4iKJWfKIaNhzoC7VSWlVvKYzXvcsEMewrgDems8QpvEfyULYPxRzhQ+JieiNelODYeCpjp
9M8FbImbNic7a5LgfC+aeL5nBZwMSGx1M4zeTkJlb/sIkgOLsi5VlBZ/YhVitsSBrYRKpOu4V49T
qYUyxSwkk6/+B2L+T6Si2Kfz1jMQLXPxlPxxrri3hoiOsVOeZSEehSjxFWKhCJKL76zU9o/nU3gL
PHwRR4h0Xd3otAN41WXjpUzczlyV9eU7WIGqyrWlhWPsTWHGfbDuQQpVdsDFDej0TpeSvcJ8IuzS
YElgl2BXzUlosMJCbL8feBsy15Y4Ln/0tgzfx3xDeeTEGDpzBvVYGMZARnWfB5rAqrCiL4fTxRI7
fkjxtT/shGTelGxf93tGhVdLm1JwZI7H9b7II7H4BJk8gESeWP7zMtQN4JcFGN6HnL/aMJ8z7EWR
Gamrjkp9h3iCbM94yZs9ApI32aULR+p3FZLaDOPvLXr9g1JpPKBWXgkA96RaXtnS9Lc/b6BHx0do
P4nypHNTxaOdUcck/VX357gp9LKpo1+/M8nd1/2JGKra/q/NYfTtV5YqIxACMHjOh5gUoCQBxjG1
VBYQ235Sr8osP38bydMG+fMTNjWlJs3uj7I1O1a6zSqhrtLAq+9HdYk6pHV17JUtSgY4poecS3TK
xPzJZLMY7STV4y9a5ckYwKDpn5GQyeFAw8Y0hllEZygEl8mF6m6S7Zf91ajEcCJ0FJZyeNJPcvYD
bqIXjmg2CDmZuyuTgAg/JQZUNfHjAa6tsSjFcelEMWb2gXhxQrRpFZoaPVj86tA9UsmHmSlBiCBW
v0NAT4yMgC5uO+F24QvMqeB75JozI53kedsanGNzOPmaYUGm4bvC7PQqh8y8qIwGZn/MmIGn0pwL
SHnW+T/a5o7WfYt859K5XdCJxcZSKwcr+ZtCk1fNKiFc0vTMSVpLZ12pyKAlw9Y8b+dC7bQz23kK
hA6O2gDUByWDw3Nr+p8FBE8X0DZUtG4BfTvianJOn1hEAVVFF8CX4r6yk90oroEjp3qFXzMSuTbs
vJrL/dvxJjnZ33qT5GK0vKjwETmsKnsAC4ocI1Wd2SiCp+9zwEctShy19ZSt15CWK5fadlLevJer
vNQJH7/OKLR2s4qXpXaVyD2zKBC7KzywUfB2aLFh0gzH1oFevpEf+0Qzo/LTaD96K09nHH4Rfr+4
8Ki/OV4AYD2dWkISKV0jfND8P9q+A4O+5YC3mmMSS8Q9A/qOlgTPtCY7mXm3rP4GRik/eEfEgAFz
Axeo9UZ7rAWa4bx9Po7Pl3XL4mSuNNgqR3tzCAZg++DL4Az70rkhmoqtcQbZFZf5tUJk35dd1ofM
b5Bt7CLgEbtaYZAqYWg1kJ3bozjLofdB4oPeUNLPWc0iiBSszlbiooO4R3x7iOup0ojSp87URaZ0
Ysmm/3N9Px6m+Mib+If8rQsrUMhKXExK94/kabMtjUwozf2UbphJWy4DkyAq748gnWZriO1BSoGS
aegjzYwIrf8J4RcWOOOrj9Jgw+DVdmdjOx3XAZz7/mnpMdEnM8Hz+aNJ1ARzuevtBNv+1p/D/nF5
U8uoahIqYU1pMQGkpGRdAJuSZMp1HYfATP3QPVM3wAnr6NqCIM0rjLqpGz/RRC8YJKTJZp1JuLQA
IBgui6tYDdXhqq/I3Zyp196HzORcIKwMXei03xtzMaERbvWKIXSFdGpN4N2fpZSYn8u6rzzPBuVQ
wI+G0Pl0OnqiuMUQcSHo96gOtpDQLlk/CsZ+4Um20uA405KaWG87wN5b5gllgrU8m8ALqFMk7Sz/
2OOTIhxEViDKwP8BlvCefE1sqyHwAIQ225lAT7Ec9f93HJNUl2uDLMESZXtDD2GBs5b1HCRbT3E6
IcwbZCZlvpxV8/9ktfuZjBcyWnlOOpdwT733PAyHvi3azJIcwDCe5xoh5ICN36LZN1y2VBx4Ak2V
Szk0sAdiMoxGmm4UwCSiFsyDlOWKu/BG0p5z+xuJ/aL7CwPPLVO6c0rayaYiHAFVc5crtDnsd3ZR
sQUQE9afHyt0ZH+//kguecIOzfCDdaHBYN9FmQkaFNvrJMZH3vjTGMoW4dkS8cGZ+vdPITjJNskJ
xZVw6LNB66Yacv9lSWi9tzqJZX4opk7oyq5nnxyZfkiCX+PagjxQSzR1JJ2Reon6KfiMV1m85dUV
GY70xO9sUgQvEwx5fvHyWHpCKj7ZBhV6+UniVnAxiH4/I9sLSb/I6U0+de8wd6R2vDwUyCLmxbN6
q69/+LQ4Gp7kxLVfa01gtVEhcTPn+viyIoSeqUyN4ns2lRa15AEjRTYND48xAId1EUef5x7wL60H
BocDXsmObWLBHSou9vb0QWOT8ALUxkV5DtbzJ+XOlKh0kwneWou0vib3uRqMPTSj3aDnELW2TE2v
A5N29mwoi6xPsi7SZkn2F/lmUBjq6yR1OcP9e5Ln/wZSlayxCcgUbm5ShcvsNNrdAic3Xzra0Z3U
fLJs1oojWZcsVRG3Yf2WVbI8SaCCuknhZM9wtBOCTVb+QYO0ZKnpsCFKogdSWrQQ1gyJ1G3us6Kc
pdhdzSMbob/6HfVzuKGF1F7Xk7E1WcctQn9G+IBvfnJeTUNbTVci6ceoPw47GPSB8OUySpO/mI9I
2pvmdtWAqLkxxS3l06UqX0TkLel0yRey2NQ1lWGEah1ulw8+QJ3heQ8cAVna24fOVgBcT6tS5YEH
cLktP0RlFeaIlZIm6/T3vv9Ww0qpnLPZ5hCCJM1OEsp5tfsFMKzsU41aLxHGfy91a0z4mWzF8Mc4
Qezv4X0bcIAaJyF/UsHdaVXO09YtJSrXVVbeWVyHADVQkrNgsQYYB2kZOvJmUTYRehwwAoA+qHeo
0SvLsxBsAzNAlEvSz8/4FyFTNx1eviskvlUiV77YCWFPlJjbQDrVT8U19IujrW2C1hUk1mkDE3xE
0ESu6itbBl1CXtChNxDnP6Nrt/ZfSgjrGKc0oAcnAXvKPGM14ZI9sU561GJAKRIma3BYQSJqfboP
Rka+dc/KHIb6aE8Dpbq3P7Xmvmo6d/6cYkobB4TyNZCT0Da+R1iVLCwSbrXiyHIH99y/DJ9WwAyn
u9L95jpaJEZZFnUYNIfVkYjVuMNN7CfZrHfu8/zjEfEXee/S+NmHAlO2XOm9jZ7q2O9Ctpc7RAy7
lWOX0J+ucmRLZKcVfIsRIztePPhQevtYQefE0X+FI/TpilIyR8xZHqOWagGyZHJYNhXshM+JFlJk
V3BGxjBzht5ymfRrvRaW5f8v71S9dJGc/vHQ+n8gmcl/0Tm5yRdOfnztXZyZU2s2IuwgZfDTzPqA
Bwbu5wFgXZTF/+HswNeCLOKbqcZeSaB9GYElDfG2diY0cWUaxzqENeBw60ws+hUd7w1fnNQJAT6B
ri5StFj4CYj3Egdh9/HTGn6Eys50QEoeS8rACh6oFLrGaLn8B6pnS4Mm+UG5HLgv0rZtt9LPNM7T
uh+BGh+bXdC+5xfHKpxvTcVtVufGf0sc/WcD2AL7kPJdGDe7ac2wKBZ1zUxwzT8uVdinZMLZuTBT
2qga82D4hv636XCr9jEbHmnooopSecSVRiIV1ZQa+YhOoMomFeLv2eWl5xby8NE/rKLuXKdThnFZ
jZWfKhCjHpcZ6uFF2rVJx6Eh+MXbB72yGFF2TXRxPKmBQ0JAmAecuWr5c/DU3evD8VK/jbP42hJ/
Z6p+IA/XfkBs/t8lVY4ErwZcTm9FbEEmsDgw4H/Ta/4FxfX9pUXNaH/7oMgLmzJfLzpn6281+pcM
tk0MBWRBIy1FpO6FUhFajJu1+YTCVHlTpxv2XlsxIjjorawX5fcWkPRdHZg0rVt8qVcui0+UKSIH
bu/MIdVR/ZaZrMWGyo2Tm9wdGwHhUocmEQ1akVmfMz4sVjxAcvGLAJDErU/jhcYUQjqP5p7tZqfN
SCbTC30Sz8omMB8ZueL6s2UktMfVs6Vly6USF9kVBv+zICxBFz+UtK46ImkiMNxcepPfT0kk0zc8
7CHM1tBhh9KObA7y2865saYdUc7HZmKEf4/ajmsxrSZkvpBmJZ7Fh5YXvo/A/2DoG7PSXUQ8/JZZ
ycRkscztIFUMKzQifxeHlvagoINlU6EUIoN/0l+ntg6/+0Pkwn9yvZMDhc8kns1uzXG4nNLh7QQu
zrDlvcmQtOBUyK5ssHdFHNnD3ExCr2wFgEkXirFhjg/HPN9gUUAkO8ye6IdgB89pnwz+XAlyfRHk
a4x1YwWr1pdmR443mjAFWyzC3KCNq651Rp75PmpkQs3LZKVjEkFwxLBod0sQiEUIbRTV4AQ5zEsw
aY7GgiCb8eqOoLVKNyjkV0bWz9qtJ16Vo4IDsgyIQbQUrOCVdQ7SNPQflS06yj9LmkyAgJVb7shG
BLIDaNqthl46mrvGR02BQJMCfxrB0tGM9Qplbfpm7PJzsZERZcHydyAon7rtq1n60gP1fxvJwQOm
5r9icZkFfydpA7NfIuI/du9aLvMz0gNypgy3ruLIiQFaHsOKilAd3KE8m+uzgTckBZyxN3MVwb6t
ipxmgQQWqEWKrTBx96lOFD1YvD5w7ysKC8foaR98mNs6JsXgp+rch9PjTONME97ut3joDn0sX0FJ
7UY3R8bLsgmD8CHYE2vh+gardmFdCom6V25rOzVdSF0Gxk39QxKvcFYe9F0x0icRlJW7h+CGxrOV
N2wapXSgPqrpLpULDD0fTuUGibHDY5WEDDJJwJks3FxfpSMh2CrIjoDgg0rf61JU8EdqnLDKt5Mp
VkeTPRTl3cIGKI0ErCNEs6qyP51NkVAteVaVkbV2Fy2S715UdqIhjK9HTqrpO2Ek4w/YUMFmLtyV
HWhtFKVRFQMOt/ZfeGgbmreSPGb2LuvYpHU7i4SyfwI8C/5yFAtDR8A0FRsHxChSHxHTjgsWTrwn
szAdcTX2EU3Sl4RGzDJ9aTW72B0YYDRm74NrU92M6xPQWAszW7NO3Nkaa3RUKtzdhVimIvbsjnnb
lTcV1vVa8dflyksgO2Mzno+Ucg/QhEz79YIqqlTXKa696PPdR428cTjWKEEHmCf+nKNHKpSGxSJJ
pzQglKY2z7eb+PuV5Mf/wrMKiAGiAjvnuhCJ9ySPKLbNlrOe8rqE0OGBNhgbK4nCNtS/01/MKQSR
YG3lsdOJwRf51vl9pmPKKj+H0cX5KTdqrVCmIRK0LkXf3ptt6G5piGhqFdZK6H1d2WXysmkrP0Kn
D5mCqoF6CAEH/+yjYNE2zJmJ7pvl6l0RBURT4ewxdHyE5BJMVcHzBRd18AjIMAlBCV2leMP2LJl0
sGfjiyFrAXuvuux7+W4d5bFGaPv1B88FPu12JalpxV9f3Gfeaie+QlAIwsqksV4eVL0THlzFoysL
0HkuqUcStKlsJkOET2POyydMNctt6gMddcu7vjy2tLC86/MwYdoyYhat0JbjEXspvxlw2S2vciZq
UpYGnZrgO/fXJuOisRTvOGqWvTM+AuX4V29huXobxWXK4Dv6T6+TbFEbPq7+zcAHmBSy9xbWcqoB
P3ajxMmwEiN8QCpYF2N4fzx9T5QRx5vJUY3SqYrlYycX8KuIP/xVacpLWfPPyl/UQgc7NyslSJrj
7X78KXKRKu8k8hD85WGoy41sTyr/UdooO3D4si2Zr01Dutprs+D43TSi2zp8UCevUJOfaa/Q6tY+
LupSQxjUAQe9xjfLi8lXwl3IBX9lFLOQnEVYkbxkuGSyMvkaCdvKAEkyu1tQeKYMRzczpIQ0Anui
pB7C13f4j8sgQLaf5bDOs7kCC46W9bTmKwFIipVqjM1IwpqEoco3NYPdsJGUC1DJaT2RXtkRLhLE
9c9JnBw3q7AQBUDVkqIxSYC+zo6AgOYIfpHYCj4ATBmp4l6F/W2TC08zisnVcILm7v9Tqfwkd2X9
UovBkP5LZOUQxPYUgsvjeiH4AYMpR9IdsrszKcnEhgw4wWym6kTe1czfemYeWOJure8BaCc2H5sN
kbGYWYO8GGks6n7EYitmk5sMelRNuajK2b8pgi+mJF3WjwYUyqR5l29RXPiFDNEdov0Oa2/Ywb/N
PqchrGcpQb0GWCxcfTJYDqzzBRJzAR+HX9ReEnXNaYWN6KQjjc9lDJL+PGa4T6BIBeiz2uf0PuoT
OjUVwNRIl/rbGiROwNlOjHFAbqJr3agkvKYqSBFW51bnwv/GTY18ZWgOsNPMPixgJo+g23UtgHkL
uD3uHPBPKZ9o9odUNAKXIo6pf7cJ+jGVKDFbEOW4duOIEq6B6NHXlZmxm8EE2uiRYfZSy12fQJs1
LNuQfUxmvO+JP7ZCPwsRuL7yiwtE72qVMBaPBusoutwY4p3GPxHvVr7nXAuG2d2stNjI3kDXtKAg
XgeH2H3HvF07fRod26255rfD8aq0lChQaiXk1anyb1F3We4peHlBPBYm62VTcwPsGhKRdySNJDvf
An/OZ3hlwY10uxE5+uyaMjaHhPWIi88R5FaxwSs3OBok6c4pdLeDUn3g0bbdYt3ZtR/SAraKKC1j
gRLYophZWkT2zCKA+/G+ihMatY6spG/LkwUxOLKvgwrQnS5A0sSp/EzE3y9c5+s1gvpUoKFAY7pZ
CPJsljFfi7WuZ5AOWtqUESRkTBfYUTQ0lUKpFg2EQNwUEn5BrLcOi2eEDukuJMFr2PQMpTVKEEBL
o9L+14c6fFOh3jHtDmsH09gL9Pa3P0jT28J0395GhrezApAvLWRF6xTi2mUR+y9i4GU2UGv216fq
PmLLr6YUUa/P1C1STrgva92iRKe5IFmkjwh8VPrS+EuxAfcOOgoWjgfev1tREJH977W396iUHg+b
U8hGXOChvzzybHsPJchYLrKItmnghZgQV+3PVt7e+aX/Dt8FP8tBbfokiOEyTImOl0WpaxR4sa8O
wPgAnGmbyHXqYjXIrTtxyGBHpFKFculAbFKnr/zc9smKZbXsyjhWFWD39wWBEn43j5rHJnnOm8Vw
Rn+aq+gtRBx6WwlodsQTrpCTS/GgRA+uSP0WDz1be0Oyz74Rv83fm4JuMxr0WKoCUH25HYtLPN6V
6GenNxbdDN/h54WuoRKNrVXy1oYhnM64HkBeXErVN8A1N1kgG5po0GI3fEtcycvZDwoUxdYlZ1Ei
kyzKAwOA7XUOmlt5EOGrgHAfI1JOS/ehtikeQTJY4y+hLLrfvCyCVSqxtNZ5y9uT9hjIf98EzwU4
kDqGiE9P1FuQl6h7p2jvidwdeGHe+GT5OonnpBqpkaQRuzngPFEGy+aErLaR5ZC19iGy89rlMpqj
WxskfO3I6pggM24cTxcT8rzsTwKauBagu4uf79TfQuOHtHkOe/ZfYfiN1wmXHoiD3+ShAyoRy2ed
BE1wXLXC/1VgGAM4GRTmPIrKwNdqFLTdJZxR2ad5hOfBx39ZBscrkhVx/1smfDduWNcB+LZhcvoo
9ohzdR20RLkK/7Ju/SNOnR1k0DSgZaVsPD7A2xdzTApvGxw2BCUFbwxSc73iYSf6pmkII+rjY71C
6LJFhvF4BsdnNHBIhUUjnn5GjFtbkmgpzmR2IyqmxruC6SdKAn/kOw2FCwg7upVy9305Y4/PsujL
FeY+XoxAOBqYh0w7rEiWrwB79STf+BH/uIwBFliPH/GTji1+mmSJUOaf8Ql2HgjixxPiO8wLT8a8
Lmd+uF4nzHJiUGYoVQLDXF1++mh9p2k+Dg8MnJhWLn9+8MADGRgAQ0B148SV0TmXlg4e/HArRANT
B2Wh62PKzI5Vbczv/NnXhQjrFQwF2PX9x3gkkjYWiKSTsMlQkN//py02HlGfIzTOHx4EPz5McLYR
D52Zs4G5qGbJOs8CBskK+M6u9wIH0elQ4Y5ikt/cGgDHcnZjlV6Mprri9eovYrK08Irn9xiWX0qT
9RvQSEz0NQdL6DEvaTDe0vKBHIbEB+0VRo3aS03MC6bRad8kKIoQzzILlsQjIci7t4HzidEGhfnk
6QMGGCbhlIsgLqEwSpwUxB0LbF3xGGG/jGOGNFBPcf1ah1i3ImDqmdimgFmbdwQIdYVjJDuTLR6O
CF4nBPqM2zyUzoG/F1S8jV3OaFoNTbicGJuCrTJuV1GTi9qve44fNtnqyx7VEpB3nHKNwTynOaYb
Wq5VGO4urT7rzbMGyMx6jlnpLnsP9u6Bcg/UEFkJNiuA29ITVxsWZgY/uefENNJS23bp3u89n95s
KFtowtFWI+7OeV+U2sTHzYPy5Pq39D4sePSfqf+ktX/KsaJNG6nicfR3mdzwNyaQ3DHRIsCXC6n6
YDhGrv3PKiiPZzKW2+CDO0ulDxPxjxkDPfNlJn4AA6MKtil4CIS3llWZGNNviKRJxHlRHbLwxO+R
aJ/gOysyL+uCEKx7xu4RG2+yrO/EmsdMYgMU4HLGpfDMpnk9gkqbk6zJ0xHtA7asNBWvGdLyQ2E9
50PvFbCeSUS4xl6mUYCmcjMbPjsvKrXxuBeUFc1f2ulVFUu+zpyg4cXHrj519HKFkd6ORTqY5dkm
IFp1dyVnzxH3glbkO88PpHo33Ov0MOXKybAFDXF+UIkMH4f8zsYii4YPQ5P87J3h8TR3+VGH4yAL
A+VcZz4nrMTOuCUSrdxs86zm5KROokb9+gzB6wmflTUW2wBO1+YZO6ZtL9Z9CmfG6x+h21aZWU0e
g43Y6Kqi/86ff8e1JxkAT9c56HxRw8o0ezjmKmgKfeoPlZ28Hy6OriecknUhaMAgSJp9XLgk+V1H
UdJ1d4GEr/n/zGSGqsluxqbt6fJ/qhS0rYks616uTCG3vbXF085Ky8DK2KgJaWtmau89HRq1KBq8
U53Oro1R+zJ+Bj6rxqB2dsbVo7wzMJq2ZiUvAgLcTs5Fiprg29Hfxn5Sqa3cf7W3k2AhjhtiZedN
VI6UAIflKuNXyU4REch9hs0sFFeHtoop8h9V+TyDVyRMDU2uTh+wz5c806GkLcjTaDUuaLKIsSbL
099zE/CG1nEEnvulmurP1HTuQgAe3jXjgPcCP6370/lRH8ASvon4YD/ttNBaH9SCIrv8yDrXPnrB
CU1sxH5TeAhQSBCYYyuJM7qmEforvu17ammB+gxcDA1UTvhT0Orjt1AUbxK5u8fkanAdGfMCs4fi
b52ecM//NcGqp3PEww6LNadrT0ult6jaCBUr5ih4roPW6l3q0zEDrFwp4ymZ8mHr4owwZUOkwYOF
LtQPyRcNkTONEMlMwn0trS2KszKU18crWTgLwCrWJfUdKx5tiWSAhnHAHcsbz5Qfw0zxUrp/iQtZ
e5tPHva9VSYaxPU9hWzaTrvpNCqyDHSoA97aJdooedxmewgohLfcPNmZ1+uc5+C+WTSuSA4+733b
/b7tpR0/nm7eaY3NbWA/qcCGtkLnoPkbXb8VH7tvmydEHekypw4hQH+urpE6CMFwc3Nhb4Lmi5mY
lKg4tRraeMXC6bvtGMB29vatHoxcacIV/Lzjk0Qeej+eBa5YwzlHdKY6s8hYBa5kxqieJ1e0nOon
jA/WTAIW3Ageid+qrtbfonQj7grqhIHFMZBZs+C3eSkHbSdDvTjfgdY56uksR8ZDgZBNt4yMgozZ
ra2QH7hK2LPeB/MBEQvfmA8oWJfDdYt5zCzgMKkVQbHkXpmd45iAOsV9/HixuCof7BvcodnYCb8j
knU+XX6nDoebRpNdYid6iw0t24mxjZgkQzPtRKZDHkyC4xLURb+y5U672p5T7/t8Pr1WQqP5l5Ri
FRSXGnqH3e9W1tkQDFo0DIvVPL1vVib6Ibj98NmMOS8N78Wod9pen2hiVFeoW0M2cYZN5KvZkZFW
hLVsN4a3NoCpHK8dcbtU+mG4g9pBcnPBe8zBgdbcfkQzgur8/aBdylvIdFTuCk6pKHKWL6wg48oP
t/+Ijv6X52PiIWH5IUVI8G56RZeEW9ADhlKn7v1Ax15dt0/RGa11jAzPMc2uqm8ZPQNe9fp5Owvu
7y9JNTKmi+AlQeXZtR7zqMKVL19qmpq4X9glwejPKgXd/+tRPG7fYUc8p3uW0mWmhlpbG7Eosc3X
9BYXzComrHVYtLvM57io339WDmwvClJOZG/B86SeY4NHaAdwkwfM5T8gtjq2uy9blcpAsEEHGT0l
QHM1Tq16iYMf1PSJYsrsXOK8AlD0kmxIFTJTmi+DIQUe3J5i7fzT46IcOcL3Jsm7sl1gBZ+rNGFF
e+GN3JUrDm7c/XU7aLyE3LVCLBIHwrQRoM3fwjnh0iTE0or+hS4elIMWymrCPu314wTiauvmJ0n8
3FzhjhwEGwCD0briwC6Hldy6HITlJnC7AijRnLZ3pQT+Su1SUHo+syaZDqz1EMLE17LGEZgxhiVn
cLHaXIgkYpeQJnOGK5zfOrq9sL5efW0WpWR6mfox+HybfoGQxo3GaRnhfwnfTguDHRZr431mlC73
UsMYtKGxqlm6/IixviPVPqcbaDxQCU/BdiYHw/JojIaghzF/7SdOV0Z0a9TwpbHQ43Jcevhd/Z/9
WdTXZgZvOn0fuuQ+WQS4F7ZtxWIzPIqWQY0XH42eyisvhcQGqHKFYSZd3VaSA+X+TnYWS2X6eU6p
63XUMmfxtgsZIy2qammqMtrMHXA/TMkf9hbCCa3KSFaY/qx9xzvtIS2h8n+C24uLkV9tAmOjlbrk
X3Hsm4rbmrYCuAp3NBynfuzE6B6koSeDfuut6+KvSBX/YGB28E/ObjPbiIq1TmOb9/pBmxjnPKlw
DwIoWq+xAfFfMUoiN1U36dAdel8d8u2rFiWSkMmb8O/4fy9rahi68vQBGiKq9ymBPH7+s4TxRjcw
vlY+JGtlrbqtQoqJHUp4ESv0i7nyoosxIlfppfZRho2oxtMtnKr6vHAWAOHpKlhs7oFVaNp9Cs1u
2ase/Hu/fvx3zq3tkhIL5XoqFojk1iVz1jVZeC1yPLFbkM6jUJKn+fIFgTyMwl68ehmdpAcY1/4S
JAjQOMuBP9AKify1RSJSH9aPcgWpj/47kYzp2aU51vSHrMD219wEaK9G5X0iCDJeQjrAn7c82cst
F3//MJK4NRbmRqJCrSeKZGseWcmiSp+9EpgaMlFLyGX/8Se0GX6/lDm3Yuw67xczHKAAqwnUcm9n
/rPmrACAlWF/sYuBEoYvr/6MiI9BTfj7jkx68XMDnEObgimQbP4OLWgIK5IiV01lqeFCPk8OyYSm
IyCiRehp7JOvZjijdocldIgbcLnMxcqdRk0jg3ZU+yGmd26D+RTKE2qFgUM8DBLx1RnLvb4bgrHt
qiMaQ2kc3Q2gsbJSyYnvuL0v2w1hBZZDE3UFQj9n5Qbq1eLdGa6i7tJKzbWL79KZwaBNDbdnNDj6
xmZ+xV2loK8Ye65g6DSwZnu3naQkWW5jqOwy+x9RqRQaiMCeGhmMdWE9/NagkDsHGHL1/VCXHk/2
MCg3XUaouystM5ZHp95DdUnPvLld0DTsCwx9wyNbsuOx7UDb8MdVbFtOD9OJpXGR6LIQwHN4tsAc
qTC5SQQtVultu1exyBdZ+VH/iTAI0H2l5Cpl7GVTkDUEc5MPnxUZXISR3ZiS+FnHhgtvupply6bq
p9pG9ox9ekNo6yPk685flc4pAuexOXy7GPvt+0t6RqoR8FVnGYJ8Oej7tow/3cnPUlTI1AWE2n7X
yfGt5GfIYrmxiJmPyENIRcJIMJ4TypM5W9SYU4XzyRCglySmPjky1+j4oJ42kmTJmdjBV1bFNEeE
7BMuV5rnOesmo0yK9EIRLG1lcHZymbTHgmPAtzgjqHkRjfmKhhQzGyikhCkvqSj5WaeA9h7jPHni
plvfSxujSv9M4hM2bI/pni0X5p+FrO1v5JOX+MrCB8WDRnZvGK7lV2tqQYOeTlO17Edk9GCB+ZJm
XELcy4KNL0sujBs8ZF47LaeSz4zhpoOfYb2EeNxNJfKZYL/7BBtDlj1hU1iD4gANnpvJmSlX6RJ4
lhPfTBhFyvgvuXjZ9pcz5zHcvPvV4Ccs/TqmSlB3U/zQsxeTF0KCqhqLO7/oQrRpHbdFtOwBUXLW
SRLkJHKKWppYyJkh6CTwp5AXqBf2AratSCyH+a/4zCxmSjB531zErWdztdwrvQTS8k7jTHEk3RJ8
mm3B5Dzdo3nHII/Bu8auqvjaYSvnGq31bsU9G8upDbCan7VYC50ZMx+B2+OkP8YHglHjDqyaRGsK
S/A2ZiaRWf1UPq1Bg4oWoESWKYwvfyjxzcLM8ut64IM1Y4Pe8NilSPgGav7hYoetgfm5zEjHu0yc
Fj/tMoTklvE2jCmOKkwmyR1H4tNNKQP5G4CdUF933Mq6fRDuKtKsLpX+Ou4OLqRcJbYpepZEkLS9
8son49S341T4nxidVP6ui8WQqfpCeSu4OBrR8E23gXuGU4TqhAtvGDZ6DLKmmSaD1aDRlo7vqf/k
SmPIs/2NIZn/OF62KGJSCqpniiiB3S/R0eorBeGPVCgTQyrzl1k8yRI45poil4TVsm9BkaHITIFi
5SlmSlQMq5crZLOAlpST9YV5cQn6vfQllO/jFQD7s1pj8HUfbzWQEaag2rlcLK1ulL6rrY3pigER
4ofYAGGDNw90QALGPkp3txlRJp9tsLVVyrEcnuSh7dFZ3bDTk8+dpANkzDwqjw2DH5iWFFTvhcm0
HO9i1TIddKl5ooi5vQIC4FLbGsYSAtMx6Ak+Q5uLVarp2D6Z7nB+V1uq4hFWvY6jdPgmVvrNPg/2
jqap/Iig1jWWi7lcMwvBdNqdaYaZozkZa+aGZpfefz0oowhG8u9EW5sPjxKAyFR/xWKxK1UMz1ih
HHRx+MRuBbAzyCL6uXSVZU7bDzMDBAnTWCm3kw0b0q5ejS3aeQr5f2+AxzsTurxlu94QkVDVmKxI
qK49nZUZQa1LuNmp7wA0ApwSnMtSJlc0wOQOQep6Xt4xWyFnn5bRBQO5HsSA/5iK9zJjPAQu+i92
Rol3W5FhPb4gCI52/I7CN/s5hBA+CvAJqIua/vYpiSo3PviiYeMdMy/ddnFolK2MD8Vz5vA4ekBq
yHYLWDOHwKsDHR+bj+th/ePnqjhcycIJXTo+8meP8CLkQItQp+PTWLWRKINHL/OlL83B7cFaFqv4
6a2OZG24ZrvVzmLjXmNep47SzPaSJIUryAoVLynNpkKDdpsbX5DF9BsW6WYFRqbqmqADbZmj6pKn
BEgyWkFlbA4QiGv3s0lgSlyURPITC/bztL/y63vC2Wlxe2KvQLlmm7I9Q+KWDw7tSkLZUX4PC3o8
+bz4pyhMGgiVfuh1Yz56qPTEZn+fJWqj7MsUdphsxep4wW0TNAY7yHDFYFUm3wBVCMCfMp6M7Vco
URD/1hj1/FcgPLqEL0JM9na1bzhd/dw6Kc7bkR3Dmxj963pdFsDMCd/1BrmoqFeJxm4PZQmC6K9O
G0vUiNLiNA96t4jI6qNBzTKTeZ6xcsha5I6YXnhvdHOQQSqCgK5q9uYapVUIG4szwfR/haO3L+3l
bCEvDxCFvq5Gu3q7D1nRLZgK9tO//7B3dU44L0lExWa0ylJVyQVV8xbfGV23C5i6uDJjBIvkDe7Z
S3lyuJt635KDrYRcEk7wixiwcZe2KawO5edxrXfTwHqyEjxcbADYQ1k2kCQyGfZOn+X5y1nfVMHh
sq9xrYbJtgqsHym1Srg7222/4aIrapj76oLvwYslEFQOvBuSRqglE2oSpskS3HX+aqG+NgH/flRB
AFymQY1btEzD/nfkbRd7KTNhnCzRG8F2zg2RCTiby3CslL3DGRESokqYfEdiaJ9WqhK5N5EfkfE9
nHOu9ntUfV5TGx1a0vKz67DdugC8IlM2dLYlWDxuh/daJtxQ+TkEbj4rcAguJpOtL0mqWvY5vTO4
n8XCQG8Nc1J6KLwdqWFX3VnxcMMQeb+exKru9aE4Ba/EDXmF1+/9CvI0vVLEhg9/9W3lrzNgWLqH
3sctB11omkiiYE5h96gGXYgRwvu1x3H039Lc/tXNK3KWJX8YpKdHeBWsvjL/i6ZFUzQ5pkb3Rb0p
8d3WsvShCz05yyP3oVDXMlDTMeWAQesdakPyfyCDJI+jnLRYvmAwIXWX02SFugC0r1ioKSv9KVO3
gJAIhofN6ydK2NGFgF0mK8JgN0WzvCRy0RS/G01yOZ0XDTZ6Za6XNhVeh0DT9jBKD3muFLv/kusr
DiG8cNFihcj8DaieE86tAsCBr7d9HEHO4BAku2fSCLeonI+XObhAmjrOH0FfzCfV2go2CyOIdekm
NGYDKWmGdu7wIKVfjtdnc0lYAOMFDR0eLRPPG85ztgWmvH0zbWPZOD31Ia5Du3mRlRLXmwajzTSi
FzOIS1qDJUkH41WibQZ0TBzVTEleegKMkqw8f4i+I8kTCcGMNigw00sH0APtbN0YaDeAtP7wu2dp
TWDSjPy28ZzQ9ow4Vwvje0RsUcRFVx6jmFAzBZau+jy0pti0kQC5x2Zfp/0mgfEbaqkhieEiQYkz
UJgYS3RusVGVAgUT3FzMR6eUwgEwkPrdSC6z25nmOEKEFVXq19DZqB6YuBlT+wDsD+7N3wMPXmSr
FZ/ZlTV3aTfQ5Qk6oMya9VIGhNURG6p/PAC9+U6DdHnA3HEsY/x93Mnlgw5e8uLky5Mdu5aFk1H+
w1GmuJ1jmKDFMfZDukkr0kcx4+abOP7eQ67r0Ve2PtEi7LNVjRNOowhaodwnzcoAQ+U1qRp7RZHx
A8op0ML04gj8XRr7a5eX9AuvK0CrRxzTGG3aIG+6OWYwnJIQtnxg4mxosCuWxz0pfJwRk+Xa/NGo
JqLpvgAnsxLX7oJx4Ih+OBBgjBws73AIcSYwEc2bUGmNbfDe1oJOf+pSfMSKSP+FwNCaTLFTA2nl
tQOhfMXrZaZc2+s6Evl7zjmHv83cwP4bnIuCIttrDndkLysSNPAwPyZmvosA7nzOkW252Jfs+Kex
c4KIC0WSQ/3c8mcr9oi8h1zJFmJMG+uj5N4YjEFWiRsj9MoQk9AkQY7+hHMhf/Z+D0mgKbrvetpj
3SvmyYkkmow6BHDpNBevho4y+Ud97+Xfs3tUcdd50ryCIXYE3J7G63A2vjkSjw8/b3wjnTWySSqD
BhTFpxFyUobS3RCnDmlr7YN3B822KcpOFEtHqsspZ+0GJ0M96prR4PJOLtAGA+Jh1iMKlJ3pZwmi
mmErFUgMMBTXHJ3mEQiAzer8V9WlkZIVTw7acfsIzy8xHtMqep9J0tvRtJ60RyQ0rFbxDm2vDHZk
SJfvBwfiyldBEN/JuUEKnCS0qDFX37lhDUk9gwdHg6wDFSOTDSR9mawRtWABK0A6wN1UkhoL/mtK
OI3Sl8hJAUBKLDBa8p1ES/ia+tRbdFvl9H4Gm3NYZVrsXBIY0qrOsbBELxpFxoMpq2bnFJVuS7fi
AbML60s6WIJD4x8GWV7QENj2VvGYxNNnuJqfZ1/cfsAQb0+XU7PaF1kgCvk0OKEcI8YWL6lEYl3U
9ZxTjCBtSPI9abKy7xUw6cqvJEaLYM7uf0Fnw/6ED4HpVlMGmKzehC4zI0R76zcH/RtwnUIj3Kyh
4dn4sQcPY+KWuG4tceN+bz368h7UBCKfXXgiwwzyc80MA6Bs5GtNBtmBXiGMSmuXovsFYJGaIeDm
H264Sed08SZoqZyrtvV92/ht7lzUkmVqMO0wxMy60u8NAx9STsxuqrzpZBNRFJi1kO3YtDhMK/au
Vs22m8If/wJKOw8NSU5rluX0JAdA7o8XTog2NPVdjiLE0bsgz/azlREViM4puJCL5GFCTT4gzHoE
s65GQfn09w+SoPkVP6/qBNadV13LJt6wNj9kOJkxizL9/BzGwfA+CwdeQCTidECPEgbIsNeeZ7yW
iMcll+59uYO3hKiUXUfCmOx5QcTV3jhAGu3bGY63JR2l+2qJRFNEp6l3VkTSRjvOA5oB4BXPQEbE
mXgE3BGo5tCr/GzYr08eeoNEA3d1X5x9XPUa5vNSFbfdrxUdM8nxiNPm6Doskt+Y5KoAa9qn1tGz
EAiq7GfnjD/Zp2hs3vkmhFyjCVKoB3ZsWvphOlwz8V1Tus4huN+VTctBWHPFUw5IWUmWvvCh9fRa
sRKW9ISFBYOO6lLqUASOREhhd7KC1Y2DvkU4fvzDa8lIQef5Qxnse+GcOT9t3ssfGn6LC3LVqK+y
uGvbfRGSi5UGiGBjJbV6xyORmXafTUrQtsO3+UnhtKtTiT2hUiPbl5EUbLx5LRtmpjfg0NFUvc4l
SF0kJ7wd4kxaunMxcmb8h2/RJQxrtltb0eJ5GvGgL35BlOwpHw7rtvs3xgKIKDnvQ+pfaW1fioMI
vDxXYxHgS3lPkHvO8nDbPeDP/nFVwsSawLhdcrPGdkUonEEZKyVs+1bIoWxfaRU2SRJHMNN+UNn4
eg4b9G0ms7lZI4kQ9LTtbpWXG1yNep03uo5gjwqTgFWSanJNFFSH5iOnZgH2pKhpCuasWmdSllth
MYbmznZHHyJiXKGNinwf/WZW+ssdCxb1iJDcImwH31AMax6skpSOUblA7VjifQ+Mb23I3ndWYL9s
6lSpDbjuBHTWRFoPJ/0nOmP70UyoWeGMgnz5uyGb6H7dC8vFeMAX4T3D4Bve1tDgRqgNhOlYVPPG
99le2fRIrqcgXXhcvnGiH4Z5CY9OkfOZ7YVTQREGBzpwiRD/wArMKB651Mfg4JUm6f/SORdfmpCL
QXhnXr9DJADyUhiv7fj5jBJ+Q/zfIv0SrTMtw1pfWNMSXe0O+q/+1OMt/Q5qN3+xEwM8adm9CKXQ
jYDx34PFfj742uyOlg98XUKo9JUJBobbZeJGpA+B2NqrntZ9NeYEp99OjFTJDuwNTlVARctgiURb
RNfWzYFQ4xDExz22rlXETwzTRtBvyhO/W57KxRO1K/9NfUCC6ZP4rFMrq2BXkGlj2aeh0LFjb9yK
i302FKObSpDJbHgrSXqJbiQlJUL9ZgVI6s3qs1PobUF6AY1NflXuuZJ1fr8f5vVS7CeZpnGN6C5O
L1kYjm/VpKVVUPXmT0pEjw6cg7TX0DOqldhJJJksA9AgXEVa6b7VSICVbyW2mZDGEPaNGZRPXjd/
E+FAr5ATj3n5SXLsQfBchfVB9fOYaZ53eMPGs50lBLEh+RPOvtOUSVoQPUHlDDyTlJp94IPKEA87
YqoHqBa/DfJxGcx8aIizX4vKYClON93AX6JaWIWU6AwnNY45nHIM79ftc3SZpZR+wPth1+SCso5H
P5uNsArdM+NqjB3ebV3vIj4j50gmranCdQfewyO2U/v57+bkaetF/17JPU79/w5dtrt8Yctl/peC
LozKl9CPRA4gsTzwlden+kVIpIVJ8rXyhrn/89RbYLIlU90g72OQ+rQd1NgXoekLzuDQ1wHaN+2E
NnX9z1Vcc06bvnkCYs9hXzBdzssFL053TKgjwHnQ7ZPD9RmqYer4UB21aaxsX/Bw5hmsEV2RrXv9
+IPz1ycD+1kkJZ98ko73eNUEcc+Vs7RB5hayKHYpztrHf7MwuI8lpJ56ltt4PDtZBKQQRAQDsrVe
4PqQruk/bv8AcB8g5psrhuZyaw467LcoYAT270A0A2GJESgzrDT4h6smYPF5i2FyOxEaW4arIFXD
OaIXzQTKA+5HVgXPZymhygWz2YFR09oHTWOHOLk5RaZ0eoKG6BYvSDZkFVFHWNNlQz1sJ6q5SQA4
fULgVmJhXbMY2GkQdAIKS7HvtHQGNtOL7RcNXzUrcEjRhC+DIxsutwJ5Vf4afGmy51AzdMoMUDE3
CUjh/imoKm/Fs36uCwh8dS1Wuaqnk/TG06r/e38JJaIMFvmBpcavcm6L+RUc+cYDHsFaeu5dzIRP
Xn3TKvgdTShEYVEN9Ud6TPqHLmIb7vYfz6eK4w+SHgPNBNsoVNwxIvXnw+qGw9252ZJk4X05oUvN
oJGMcM/fGP9OCp1XUWG81ntYzI4ulgVECYopGpnplW6Dqjr8nIF1cJYyLcGKdoILKONMz0h2vQRC
AucUpStMSIgaqZ9Y7gQuwdG356UlL3QuahMRDWGw9bShn/2g54v/6NfRhjCRfoOJjKBb/CcZvTsm
QeD5Q4hM/PH2GkhVIUfgN9yGFF34KxAhGNbnNg8poXFFC2MO1i4mERIXNYiAGAWnfbS1q22tKRPV
P3kJ3vBW5uKK+JntKwqlHu/unk7hfEEFzTAiCm/vC8KUj4obcaJ9v6DRRMN7/PJmE6ZQh6TCYwMa
/IuExs0aq5cbzPfgS3QKvzSCTB2uXW5STeco3het5q0PvkcBX73xgJzp0WcvgoHaTJYvtFgjpyOD
8XXXO91bX9mld+0MdyW1gHCp0SZ8qwYiXZgcw4CcZc02laX5V1kYDAIsna3JTzPYaG8leDKxto46
E9ikEGwgRbI2/BGy3pfAmKvjimLLly0YjcEsZeXHiyX6DKMtW/QNi5JhyxLDIE+BTt/8pg1NCsRY
zx8tS8SB4TAWayk9w/Y2uPCZJK8WeYjqrfFjruf1AAjejwKTfe+TUfyAbj25/nTlwwITtuFsC6+j
1gwGsK5oOXIYBRZ7RSc2BAZjD17hoNz4uHfsFrWYA9mlKQCsUlIBH7sE7kuNOimWUOG69Qp0ZaEA
fJHIaaYfvAjFiQqkhWe0DjNjefwBGlzokAbtxXHBUPXSlboBJhu3+H2Wtt9RCXx+nNtbwUqOK0FY
HqjbDNYUq6i7aNWIcIG8030hMg2OpP6ehjsYodOHFR0RUunxU4KLC3lBERb1EXjuDPtLbYVJfrfh
ffhnAw4vdDhnztGtncdfWhNfyuOHUR0FHBTLnmHqVq96BgxGaWSc9cNPedwek8Uru9Sls/GaexMc
rOft1muCXWdp7CevUb86WJ8BoEk+hB/IvYfpACoy9h8B6/r+irgu5k+JxBFVItghPQMWJGITazo2
w9Wt95o6Kc+1Lt6zc7TxrTBL6iXvHqg8GvGZ1Wc+ubk+HKzVhNd6Kbmz/k51IJ2LnSlQXzZtG3vA
5Mb4LvxbHvVh+siExhSvIBZ+KYccOAXLEfpPVH6MqoHJQmCdFE1ihamHMhm+lYvZJF3XowuKZyLp
lYwG5nyUhR1+EVqKNJEfRNGv/8XoC+un0rFpuXU//Ao2V0dBT0XU866JfM6MI46uY4W3mgfJDKhQ
7Db7scYujmQcvkxhU/WYPRBaX/oo1g1CvxbjOUsD5acP/lMXfW0XLITQ7tU7y7BbiDx8wc5855xC
YybgAXyvQnssvBWn4FwY+bkoe8ATKyTE6JhqlpOJwPz6jNYTwHtkCFcNYbGsZ6Mf1HkoCjVn7ohO
87+P/3PoAO/uEV01vGgw13MbFKimr+Xy2En0neV57uWntat6n01bP7dWPyFQYBCuKzzQtgOE1tOl
x8mDzooU/Li+ZrclBm0oxUs9SCGmU3pbDz+f+yaC21RWHif7C4AXMj4cHkfNBRvsIh5jak1b8TLM
KE9643mixL0NNyUB+5SOdqwKUhtxn1zkpDs1+gE00VMNg0aB+VGM3+g4HUb9LvX0cO0ppGXUDyI9
n58CNrcAkcEkIKN9cZxBH1RgQcDaYJQpQJMQInnWMamr8JlkIJ/5BmYx19YQgQk3m46rySUXtIjI
8Lewfpx6OLHyDCrrJv8wBD8mcQ4N8FHhbOWdDR2U41wI4Cee3N3MisErQH9BNFrf1ulJWqso6t0A
NFnVMU9vm5mGJWrR1WlHhTsxJm4k8zFZJcnXpSaUKGtFQQSG+NOcw/klSBwhWjNfVQEqUDz+7Pi6
Ok6PrNrCePLI67Mq+jE+/ceN8xDH7pZ7PRJlv5OctZPvrZmrOJ3wpVN9/6U1WVgE6u7sBKbWBJGW
rPvjlNHkZfmZsa0M9eY56Z+cuZYlbv3f3X0HINWTFhUjwxFGjhgH+sXkfTTjt0ZojC9JfthlM4qY
sCw1ZkuuF5qpzGw0w2wW29L9iEYU5pTsloiqgX2ajDEj+VUCLLWjkf4N9HXsJZ9DfYIGTzXPXg3E
alK3f7Kn86g2tyTEQPrbg9X0qvdti9MZjHbKRWlkI6bKIU6jWmrPjDiW50MuGTiur8904e35+cJ1
qpCjK+u3HIcDJ/SfMx+jLj/oyhgd77/i3cBU1qb6MIRXTm7UJtQhFKJ13zAOsDgFX9shjtOqfaxF
UEdPFO3UFryig+LzkUXUfAlXyUdCT6xjjyH+Tg9KfNseml3Jku2zCdZjE6Sf8sGmQZunMYIUkf4R
5N0rPwOPBbvMqcTCn7da5IX54IA5jktI43QPaZ4JR5s2NnYHPK0CSV+UJBb7ViaiDh0usbjHE2Yc
xGls/opQLeWmyQYXWglELw4vq/i/B+xc7kYIet8KZV6EVOSO5tYzhQayNi+E6i4kNteULgkSjs1v
MdJ00aK3delsdXvxP1F8gR2aId1MOJTOxzNWSi6DMJAUgLZG8u/JkKj0CsETrrWpKhplGsz+/KF7
wsC9Xpp+x+//syWbLTNtC0d8bUARIuV5J4iZW7kvy4RUzjBEtx8Kh8gOC9XIoFbgyGxPBFXxpf4e
v7xfDeDN62oobekD9cO9SWWvT+MzkGg6+t4rcsv9Dc6J2Fco7usrGWVAyElF2md0HiFZPCX4In7W
DSzGru6GSUWlKEPT5O6p4nED+EQlj3gbPVIpoeSphFABRRkojCiOMKh3q9kgSGYLELyvvWmS+5hI
+4K5jVU/Y71Vfq2i4RK7pVmJ1VeC6y00pBfmLmNBeWv3hK7Crb5OZoyHhtVHlXQqkEqS+jBAMKxH
4ePwjOZykzDWCSy347PelH2A4CGemUCdzeTp6tdccP9qdjlz16qMzCwcDRT5v5wbE4DikUbRslbl
R735VwZpkBv127rQKWQNi8Ke7BxRtBqFcmdilXJFekpTm0kb0/zzsCc/lKrE+Il+qTDiMtklFGoh
FWwPTyZaJ0GlnOh6YASoZ5zGHWIUBAq6LStbZbQvL8zheFPLMHWpdhDEhtK0vq8op6WC5UjDrtj8
OtXPRBL42qJDYQq8heUx3stWP3Xl1jn90TtV7HiecZo2R5RW2XNiqmeh9YQyl46Q8D83nQljDiWE
e4Js/Fwc4VtEjXa/g7eNgIE2m+LqtoEwbRpmlXVPPCL0rjqTYTSNRw8/Eq5dWUUmOSVr2PSPIAqp
9WT9gnU0NfQCo3FSijLI6T3Q7LPxrbGfjWOXR4hy9591s0goRi782S8adyRddkq3scs2E2VJqUmG
GnMvr7i+mMFeR/fRTDetiJkZWm1EMpB5YbPbrRGMPluTjqOSRWiq8WfcxIFSkobRC2RO4Y4HQbND
mF5CBVqRDfYjdg2HXESKmWYpI0ischfEl6ikHwfQghstUbwTfdKwPb9yPCIpgc3CHDQ+0kuGjcv3
UERppFg/RjdLY3kGCOWJ29RgzRF0muDdZsh8lYBJWlD6XgcTeRAYb0Nzpa4g+GIaP05qX8O+SwN+
S98M4k5Qqi5sW6hy+g+ofwEeAvv8JroraNsdUzXXUAsugrGx1qiMbUczOMqeYbauCPt9BeTN/TGq
ty859o9kKeVvn1irrhEzYeds1Ug8noB9sBtEGevBdrX8VS62Z8Xqre4CWBgC6CY5OH6HgZUh2jkn
hZNU+8Z8emcUlmknQstKKetwNbIUf0Ob/TMqU7Sbn4GMBhcojcfc0RxoWnn3f8TW82QZuCA7dmCW
nk7pBR5hQWtyuOhapvI/osAG9/FLiPeRSXfBM8IC5VuAw/swny1qKu9QUWuUXGxiLqsEI2mP031H
bYXUurnlzSFWIRPXYA7LVVmV3UVOW30+qusUNzh6NO9qJDzHS3Q7CNIecsJrOh/MvO9CkjThQkCT
ZJf3itVYbbxlfdeWKlzyjpLKiN0+pTUXJ5VobA5beBNiWpOuBodbBxdSr2nStkN8jN7Jr4nZQEi1
fN7YRrw1wRayYa/Wjl9sxfWdKDLIYyz5/l8cat4IFHbnM+FzL/VHPqEBeoxWYzbAkC2ll1xZEm4N
3QUHi4r5/rUIOZGOoa2iwvYfoHFEfBiAia4efCUGJtZZO5VKSIjv1IDXogWM3AR94YjC5uwacy7U
pgE8LMBaxTL3yhFd6uDJPOLE1MI0H0U3QXJUK7UJqGAuwXmhvwC08aUsso+bXoH/KU+nw5ku3UAL
BCNccfHHTPrEFvO336mRrz+6fJnFLhgbHlghe5koFxMbiIkZQhNP9qWGlPM4pJGrXuVwBbF2ioA3
2l2pC64kogpJmYmH6iyberh8S/PcYnavsvNkc8T82LL4K4bCP0QrpQKxzrwC3y8Wefd0RZRoe53a
AGNRp6tRLEgMRJc4L0BmzxKA4gfGSCN+43NGFzV6+inB57nzCpwKIXTCWMNWKYNd5dc7WkX19jxo
2Z9tLALqzYTDFo1QICuT7U/rWRh00UP0jBgdBFu1dY53RBNWiVIVLlj9pwvor1XWYD+/ejVyjz/D
lkgfTxFlEaQuAMHNyIgGEC8EcbIYF5Ctx6jhTQ/YNSYnwQdv/7wMbzn4WxUk9vYtRMnioJTY5k06
SgB22Z4eWKX3lcG7XffehjvV/3g2tHucVzcN5cGL4VEPDGinTzj9hLUM0Tv7sw5I20XMQDgdVHu+
QwF6iN/99CiO3ft4nsl6bPugBkSbTFI+80lWNraLwtyYfsS87wvXxTno7hSJ8f3ePJqigkEnw15b
X7jiZ6yj2CV90iv6eXfFtLwcT37NOHo91yKhW2jx3hB1IXVZOI2SRBACK7X640wOyl7/1BwJh6nn
1e8mWIm6KDdXSfSFOfiUT8OHsXc/bN2ZV+l+M3i9EPJNul3N2lvh9NgvFZ4+ozRqjy7vKqjjFar6
GFsk+v4cvb7NgKjJ4oqjy21pfpg5H7lx+OSyBwgs02+HfV38TUEyjWkOfoScbPky67R01vQGoj80
u9uiFGWUy79xltUqaOuVE2iAaMYcg5KdVZjYBLC3WVZCa8aUaGfVnjoiWAUSvWFPuFCUCZ/n5aIL
COn+Z96AxXVtMI3Gn/KfDVeLTr0oiHHbQ+pthuIzMVlgrCcsviJL8R/4jRLW19hgh7bRLXT+Wp5e
8Mh33vcB9U27iyjiFfmDDCgc3D8jt9g16UhHPdC43PFBCnu0/SaHL0xVPihRM3aeGLj6HxAm8DzY
ubxem3kjmF/O8T+UbGXaFgdecbMRJ+KFfNvH/f+AnEDzNBL/V0LZxVPXGRxIylTshEZEsa6RiJlo
ZlaFFAebL7swCzlINB/0mMxgZheb4Kmcq+RqbJyjQAHn+B0yaVmMdUxYrkTPxL1Sks+9KJ9cRI+x
7bDJa2wlBgZjesSS5WncdjicWai0dQ2PyI8bETR1jHuvcGbJpmaPl2lVM0oz4r3wMoadmd9UyEm4
6XEReoXnkW7XU347u7nW+Wkg4mjnwmnAaFfk9+NJKi0g2OY2AZV8l0vyPR9kMOQJyZBf6HJn7ohe
1iarjtrFTxd3KZlkhXtZVtziE1wKxIgwbDBosrwVf8nZ94ZIzNyPn+8TRWyNNeCF6ZMU9w23FYVZ
UvoZSmMu3jcewpSJox7D3zr4VvRGXzfqaoo8Bv7nwwfku7xgM8r2pOfuUzfzldldn20vdIdkiUna
ONA78k1I8I9pNdrl1Ik3qoJ0+m4iXprSwEnblk05nOSWBzayNsaKt2hIyIa7D9Vod/lNOyblGqvo
FEeRUDobTOEAs3sdb+APF+pBrXWragGoqhhevqabsm7Cjy1tRwUOtZ12en+l0CprHm8mnOT4W7Zb
9V197zwr+52G8gGiUBFp/6DVQDTFd6GSj6vZ3q8Dag7abOyRS1QsF46WMWqV71VMHM7GAuzvZDHc
IJA732O2dec5G5QBOT+dEg48K5DSIyMtxQrROvz3gjMyrQLjsXvXHTYcRBDZuDz03GCtasKeEFDf
aSb0XqUVaNSH9K/h9HHNETfaMLE4la80Fdy34ia27pBWHWgwNAJkcMCYLfCaEMkEOqzUnCqS3+uB
u9CnN88sT8rasfoHwAgkg09VGlwljz6Sb8i6SF4O9/nCp9MWs0gOae1FzMgLog4pRSfBHZZgSFr8
rnZ0PRwc3NsuUF9aEgTYXRy2Xl+bE+2mZCqecqACzfOD7iaRyyeMbqYaV/xEYETNHV+uTOUPqOzt
VEXgyLMW1O4NRw8AhoCdwZYZFr1M5aqKs64nI1oqVHV9pLZljColTEU0xOmYVa6dC9XDchMFGOei
Y4z3FC7usBeHT/2A+SGroo3aHc+qPp8Axgii9yElHoKpmMJ9t94Zv88o9wigkBi8PwX2QmAFsTDZ
Am+nFLT0n2z/hs5KOnRqJR8qXDzoxfsD3K+u8iLCszZxU8Ic2/A4HbiXJmbqbE0LDLjR45BFldoX
br5KwnvzbcrUmTREd8cA6KzB9CC3HEM/ceNnWNyFk+QLBZyvjtixvQc9VoGeOoF12YqFCrrbgqGZ
4ZmnJg3OMbDlq9DK3I9siIxHsAa/3qcpc/02NGNin45VpNDlpZ2sy2kh80aFA5KKKSaI944fWRNA
bwHDAN91KuhdR5LtWwVIRHp0pz3ZhzR05OshoWtMEfQihQvIiqbkJZAN2ksOzb9Iz6Lkrt4aMAqG
616GDdD+gNO7yTgXv0ZADs+7eDAKH6ZuIBgdl88NdC85TAuxuE/ClURqG5QLcF7Ylm9/CXgTBmBs
rHhfPp8iw3xSXpckSFonXmeiJVAqh+XXcFZVpbw34b5521xRydSeiSqitmZT9lYsgV+ho46qf5kh
O2Vx8CaRFEFvN6sIjaT4Y3uqxt7kqVxPa5ac+YFz20TIrbfnayvx1fai+1lFvlwIito/dwb0IG8U
5jOlkwRyag6FtmSW7W80Wf/YEcpjWJc+mVZwnqDb5F3T5teHlEaPnstiyTyUvMx3v2AoO35EQEKp
TWMcq92Y9q7WIZx6qzKiy/1tHAn9Ci6kJILdm0H/vwBcpqUX436MybRg0ALMXKeWU7eLdVbDCtzD
PIcvZxJ6COYN7Pt/+nEtbbtO7yFPIqC9/9Ccjo5euxUI6W/fwl9nGs16p1JccxtCVsuANpuE34J/
vpFZlbmdPcdMpN2WBL0azLQnG4Iaz+fE4PAInyUBRp5ZFj24SKW7ojBWZ1um3wovbLDL8W33VNly
C5DU/eqJz6S3q8PUJv1w6BCFv/08ZPiY2DSE9MvR9NxbI4GSjkwEMMXUfIS1FRHkktdP7zzxl1o9
+/SUjF7vd8PzM86p9Zyx4SoulsQDd+Y9HPkOaXIUBillHZZnm0P3Yx76BNNmnSDNiCMMaRSqUJXJ
o/59oFahdEc74Z7ou9fTtLJPlmtMuGJRF9rOi14OWnP3mZCv/pnEetPz9yWj4Z7G2aD2wcyekOQ0
PVFFwCipt5RCZC12bSKHOD03aHU0ju2nedRi1bPFqgGE+DwSRCB4qsHMUu2CduDQPeWuiEV8RW9R
MxE1ZUyAbliX6UZfnCW6AFJdJ+JWnaYhsnjaGDd+WvfXoU6nxyqVFbnQQhBOLJvUf9kI/eb2/I6D
jrxjNszeWycdqw0HmJqV0ijNnfYpxyEC6BVCJ9Yz12wS2nra+hm1ItE/t/HwzwHQaMeP8FcIRf73
KzO41/IDY/cDyDfzys0eXjq2vZp2vPF2oDkcvWy4ynPsCHzm7uWh/HIRNywNHRApXo+AzGrsCwcG
N3YJLFb/kK87xkzAdYyeLuh2pB7z1eD2H+2qPK5TAmsbv3S5HS0kHZep6CbpLLBr+OfGI7LnvnmQ
+SP/JLjPHhj0QShFRAUnZUEHOtffnJUOuKKndXThUvbgQXtdaO+pNp9n3VAZpCxuVQTXpvDh0ATR
Zgaf0gecxHGU3MjfADxz+D/vBB4mlkm8d5SemXieKdZzBGn/9+rYS5n3Fi/LNMp02SGn/Iu2GsLw
GfKH0JONLNKNw1L3XACpFxgMgR6nqi1d7LRoPoRQH4JtKv1OU/xZzWRommwmM9WhjSPqANF33F09
RbUrdaiI5E0s8kVhxYZxTh7PvyHSryrSZag81KXAdr7xJ3GowVpxGturMIamQnn4LNqhqrxxD4Am
6gKDUeOgZZuUCQA8XBzQt6wuKnEZQ04RiR+/+EpI+FZ/rVyHoTymZYYBM/49tqEYqu0E3qXbd5oF
Od6uBDgnmUFH2HMnt6pCjUJ6qSAEEwsagZkkvRCMKHylWnldlf+VCdL1NiRyAOhWmXkJzWvCocwj
O/onDIP7K7/SpEPO6uPHR1EH+RS7XPBZpvAJ2P0NyJ4Hn549MmkyTojngPY7isxyal0uGMAFJsZv
U1QWqGZcxXXA3JZhRo91clXieQrMKE+Or4XrBsKkp5L24OOSy0tmqPYn3M/vAXu4JfI2P2MGEkXC
o0+sPiBPzTfE6HVM249WVLsW+hXXQgxGLTsIrS5mAKA8/KNkCxm65jsAB7do+VE/dWFUtjq8pkUL
3gyVP59T+BPDVSOA/J5BaQX5KAz7NLqrOCHMYqizxNZeA4QOJ/J57V86AKDEio+McvkV+TgdNVX7
ZvMYI2NbMDrdFoAnP1WFlFtEUV5vqQnsedeFh3s5GaqK/efcwrDkb1nU7NKiR583hDkTyOWtphTj
7YHGjwT03VVb5AMapovDd8N/c2CV6UpXr12mC3GrcP/WdYtNO9e5kutPYfv9x4hkWk4ZKLHR3f4T
Ph1l4eAez0jhBQVgEKejjLPoVA/y1Kzo9RYL5ijcziDWc8wwhGNaIZNN1eKqhwRlSxWrhKNVem+C
oE6cLoTTr1rikA32GUYGdX+aPIaBmT/VD0Ni2mbc0AWcAq6MqmQZ+jOfqbMGkNh2IwDcslN9ypYh
SHuAdFVfyg7vDUCWoEZWctCSNZHfWKEhTw/U8+mkOF9ohfOowWIWr/kzS5Lz0EBUsU74KJVhAiaf
5K1QZC9Ne5o8hB1jDHB3z7ac1z9REn+LDpVS7K0yWlDk7DMRCMpsceRTVS+z3CQtPyToswF4Zg3l
CgDWZBUpCclMmf7q5eZEHVz005ZvmEnY2p4y1BqRtGKLhPn9wsN23NgR0GFInLpH+gcEVt9uG94m
ioQ9uOi2mxszCEEARPk8E4+oiGeGENjm+2AgUTxDWkP71jODYYR6PZtDeXwZdifoghVyIgKo5T+7
B/kkMv2JjQpxbeu5Q3YZvjuSsF6JLn2syLN8qxCTQsUkeXTAwU20n6PfQDqUjhzmtnFgzW4Uvbyr
/yDCh5vV7+Ft2DidRdJTynI3QFRQ2TbZTS1T1lk5PfDN2vEysYQLjFIfgkQoDnB6jXVMUQubufm0
Ov4xhoPCNg3TRSTCGoXwp7aTPiUGU+jM1S1ahdfdwaUM83Fkcg8lEroedZO6w0qZz0CVIzfbVX7M
K3QVE7NmFUf/xaD9hRGqEPjS0KCtHK2V6VMsUqsWrYHSi9lZdNM+EfBbDOjNR1EooAYRCdNZlgs4
rmjxWn+XJhCRPv8ZWjMai4U7pKh4A2adDqaljHDOXEXpCQ9hf7QNAqoAqJFNvgwb0vQlOevyzkQj
W6ljNnnM872vL0wUQqM6Rk23seHMbuHZk1DniTRjs88Fgx1XfSIO9Szx/2V6PTWUvzIds1XGRrh9
/+gMSYhnLgjR4THd1rt7hOX5AWIHISdxanJIBvpozxr4W9qL/ScnxxA1k1mhSYT02AES3KBtIHJC
RWROQrDZrg20jq7PWfIIv019i7XOqtThTfhxqQMujq06S+0udoNNz6lhJfgDa4OZJjbUzhTavVLb
IoipXlIzsujKl6xEyB45IVa+8VsvhEp3QBQ9QBilL7fDTlNwsWKO0CstDObnopNXZB5rHH6GzJtE
KZgMFdwZmde9IJYAF5jNAggQYp50N+kpKonjBWKQ2S2UtTihcCS6DpjQ13SlKenHR1+zaiIYlr1y
a0tPH7Ag5Efg9lHwtBq3xWbySPWXKN42Rx+hLWk4qzUA8RfIasfybmx6o3LeOs146WWF2xGWYqYy
W8kZQvYkwPg2FNeODtySIzg1cQ3BGZ6wJ1lUQfKGZkKMmanwNDgz1/ymLRSeOWgt/2ym8L05cHrZ
3zOZBUfBmB8BbXYNS2NPQU4IttWH6vg0Z/UheRzsjl+mBVzG2W/YoV/VE9x+tpkYd7PO45lQkOnI
vB2tysvs9Kcq7dbGQaczKVH8mb9dnUx694TGqHCGE/kythzXdskGpc1CuHJYftQR/I2BKjZ4T2oz
xR6pn7jVx9syQVoq+h+D1R3AyNBgJbDIkMWGOd7nsG0MOuNcL3v0jxh3PruDy04qkUHGSAgXP0It
d5s8lqyTb0vHiBwfPWQv16JY/U+R/osN5mH6cnUpiDCPLo7/uG1K6A7QiKp6qnqoh+A88aCCNJFC
YW+TUqSWk7FbkEGOMPTsaM5c898sZ5/v+N65h4I9a39BVIaT2IKCwWQoNmilKWWHuPHYXumFheiu
8I++tZH5FjewsY0zdJ+OuPvPyn+/AhqQZKqkiYvUKrsdUpad+Go0wl3nUUG1Ftoz0SpgyMidtqBE
Tp8b1N29/AFGW50Cp7CYHu/Vr0aSUsFPvPRUkD4cgI5AlyQaPvz+OOvKSIMKqWTuh7C7+LOa/fx8
NTDN3kFbObxxutLgdnALCWLzJLxShnRHeX6liavpL+86RGLKyQwf5oc/j3r/X5RjPy4Y+G1ZxSit
CzTgAq79G873Wv3/YnVh5wPuB2OkSym0mwNC3d9zvYU1HtyZQkhtm+6RTKXpFuZmtWwBUv25wvEd
b7SP1FMsStLsBze577jkB57VwHy0yrhe4jdrWzlUEBvqokJU2F1QrZMhVnJqmTbDp4+rfkJ4CGK6
xQWxQOqGO+8YhsPdND3kzVDiXQtKhtRsvYNWNjjqvHTlsss1t7rs1Tt4O3mzH2Xlo0a3bHNsmLGP
09Dp/m+o8oLgIaJmpZJ3PQwjUBMPIFwRBgrs1EBqRuVs4mVmuntt2EPH2OiRzDhctq3KkjGekSBj
YVGyqgMTPXcH+ZHmjsMikgxn8ya1hLhmD+dhZvm7Iqsh9hcrxOWpQzlFfDegREC5i0bB7j4yLmWv
y8tbq5vbEy90mtsd9grfvW8z9AJ0wlTb1+CUH8fD/Baf3RRvJw3mOiW5RUq8CwhdUBoLSPoT8sTw
llL5XFv7GFp+jVE+ZHCbkKLUuYDrbP9F7xtaVQnhQ6+UWE1Z3Yab/XC0tXyJfkZnypV5TDiRXku6
9YlVqjNklQTmfnRp+b83Wv1n6TPf6Mzt5bCGZf1brFWH6L0u1rH0fPrl1UxwEVf6zf+FcrU1rvmT
eV/2VBCno5AcJRogHb4LOR8eU9ldamJnewjHpg0aK7dPpTwx/DDDbq/v7HQA5RN/xwYD5K1Elh7m
BeNPUtxHSyAed+e/QmrJTyx8uuIecsRJZk5y6frhdsTiO8y4/PJU2GPb9IPLit8zeCp8DvbFVLWP
IHoqCBsIJwYNLdweonx30xxlzRBaZUndtf919qR646qCKoOHMGxqpOww8hR8ABKRn754SRTq/Sw1
hheLa7wy4PWRP57RhI4l1RpYALFcle6ySFFw97oE3H+nC6uxwjh/c0tS2QmaAjKbprXmAV2zC0Bg
XN8MfaYfwaX0VeAZD1cdfnlE7xDypo7rZv//HjLV1YRsZGSdojmyQk28I8FFg3yRT40C68+KTQlb
HixhqYNQy2hTpIAoRGGASIoXgNaKDc9KJ08HcWJryyWSWi7Q3mq62YXB6LZr8+N8wY580CSPsOyF
39LBBtJ2wL4up3hUDvuO/PRL8a8CXmM1Sxpo8e1hfgBfgxCd40fD9NdkQzZPPa2oVowo+o+I3yYu
VKYSsl0Hk1cKPKUuTkTmPi+vfsIjMNTa2vX81jgwUN2GUnI+O3D9ay6XJ81yLjo2N72uZZymE7LD
otn8DLm3+/zQRZ20l2OQGOvNmOIn3NjA7oLWba1wEs8APa8t91gRoozXfbc62mOwB2k7KTpJ1kL7
j6fRS+Z+h42/1K7duUp8OFsv9DtJ+uMuQ5srfn6gJqqMv8Yu+20LkApilFzDVkRCFIiqIzIy64SS
eNLGTw1ZUUXP4Gfw94D/FQwd0+CVCf7bzLuQiOl15VO67qKSa7prMLCibTGtder4mo7ag3tn9N3c
/tcd+UBZkptUMoqDLJlLbEpjeIMFdcLwdeFNeavGrWEsp49ZX6SBonG89NhmeDmnRA87ukR/upW0
nqerBhLV3yUfiq3hhQPPVNkLsENom9OwjndtEpnLeGYAmPY3XlWJp1MuLfGizBcHjMu7HPD3Xiep
LgYj/E3Q0kYXocmjqtEfm8cejmR5LNIQ5toh25qV3rqtIXPyEZFIoi7+grLmYxgW6/BfQ6gKxwL2
K84dGeVI+rTX7aHMQCj52XrlkdIZrwG3gUvRc7a81R8xhrZpQ/IhfVvuCwxxL9tPd3evE9UkXa9j
yn5ww44PUB6NvfoPae77z2Cer90hUzH1+yidMABC05BR4Gl1FyNpnQa0sQzgCHXy/6LM12asELn8
Kla6nol2K290haILsmPUEhzOzw9lUcN9pBg5CHictxQg9+SQ89xUgD96x4iCuKLNzYZX+DBpKfKR
NziT2g/LP6W31ei/FjEXFwXahhsnim5FSd2xXqCvlY68sMQVHqwo718FgAL3nFA7tP2Jw97dpOMp
LXFCmDWREUuuji7uxtJiOm7OJ9DH+XpdP+jbmeUfy3fwrSX3J5RHt4G7DfJ6nb/sHirwd9TNf70Z
OUU4cDNCpsBj2nxB+4MEpNhRhRGhEJdToQLPh3In8rgbjxc+nD9rhr4mykhUU07uGqgOZqGM8Sl/
/Oz4dGh1GV8Bbo6R358vz4OkdssUaisXfglRlgGYKlDGAGekYgMks8T6YYyX0DOB/PLJV4G0WxQ4
Ip0FDPKTV+dBopIxLnpev+boiZKIaX0ICBC0UlzrHKqXuJ0mbUc/3YguIy8kGNZ2iQ83dfy7nJuB
o3qLJXG1Vri97tB+NDb7/Hfsg+1KQnwn0PL4UDbFI+C6ibBOF7GeQAccATlUspPBSlE9h2VRmoRU
HkTpZawMUEW9N2/ukntj0NRIcwNVYfm9EWVQIii6NUK3SriLQBl4wGwdxDhHnNDHZfsFRG0qPPAW
KxIUO3b4ohEyFmd8u9T/QiaP71dCf8Z9uvNgrOLg+xyvxX2Pa9Ko6QF31EHaebkaiP9VJyK2YdYO
zMENCc0KR4tPr9R5rjAxZeaQNYz4IUtoq4jV5NHyERMQCxSqnIkboutm5Qk/ZNpuObhXQdSEXKto
bFEeYXqWRQovZyMsCXtz2oLSdo6QPpF0UGkIYnOgaRU/VZH5qUo876vDgXoeBBHeYaslRKcM2dUA
Ya2n1U0IH8wRC88ITKWE+0XDhsMaVwVQ8nbmbNjYWqgDEG9UY9wOHskrHqd3ZjefP03eSJ0HkzmS
5mz3Vv81Gcg7C4GI2YLH2r3CUeD5S3EYPI9OOoEyufv5xjisKYxdn6AiNoMTEVRNNSWVEQzVQjBG
I+JFMoPwfA7yxGcOmbw0oSN4BoPt3k8KIAhnrDynevvxwTLp/EBqgvQsmQbBwAroWzhx9IC4WoSY
actg2g6559a++phZSYZWt7tq0bAqZjXO0dmBBohR0Kgje8LaJKQTcdL7VBvZ9bQJyvsGK1P8FUML
fSngTMnNVKSPqlGFfXz/ktUmpNQhmkSoHvpUJSrqdIv2yADuxHtKSaSZA1CiHrpiT7/6UcMjxCxq
2rClgGTkwMSi/7UAK5UNPRxLoQ+QPlPfO/RraF+FIyE6rLqX0OqCqW5GECe82n0B8WnGfrvkXbaF
X+MXa30MUSFf3AB+ftPIE2ne+Y7f0LO0eMKxSKx6gdpGihxN4I2hr++npD3Sq/xpOkivMrY6W55O
DBdsltNnM68nfZbd+AQupccvodGyhoAeY9+Ax6q+AUG+TvPaa5bsBPLMov2gBGycKl1vziEwwi2k
smlzOGVr58huwltZi39jp8prRdwu7Y12sJVR/tXjgLg44goX1IwLa5ypeH13rdTOZx4O2/eJzMMD
Sel/bW9NwoLKSWh/KdpB1w5HYaYOlVY8+Uoqisfc6/Afz/Q9/ae22k2Mku+tifuvnJ0ckaIxV07e
nxsDN0oW0c9FWMwx7w//jnxqz6m71P6H1icbJ9NV6rsZj5KN2+rtt9tzWjS/PWic82YvBcGJxMPZ
OUulVBCeThFkU4CPtuW4Jb3djWxBmB6GhspeJvGJygLlRvQe6+HPDyGfwysHbJoVak66rYa7RSAD
ifWzlFDd/7u8G2ANUT/Dg52YR9Z8XUf38RGCzQvCCPF/8odlMLZPlbUONQd1J9KNa4UAMM9IWv+g
miw8d2Wr+5Q0VHlvOxfssO/xssH5kI/E+vCIBjpaZ+CLYEbPQIUIzoJbkthBUpkUIuXqYNEb/fv6
d5/SUo+OMKZDyd0iSQ1YrbCJXlLKjouuoRQoGFs/B7xWXMm+wEUZafYVYFhaGyMyAFKh5JRIRkJi
/ttAxRIYdRspvstIVKIBBHM4ZfKHk4JOtXADQ3nr1EGdjDxnqH5Qac73JdZrvCKve/TiKkwMKHLh
sXbIn5kHrFPVnyM+tNL1Cqy7Irmy31WE4G5alnRaRYj1ch+KQDLnG41pSGHTLQloSDUd23Pz3LwU
7p7LDrSf0YAlU9oTbhdQT/dhEGQkaWweSqyFkRte0H68t5UMAcBjQtTgQpaqQvwYNEWnqA7GX+1v
gI24TSf4y7Or0zPKFZD3wPWfe3K15qyVD+gj4Jd2z1AWbyDDtuG9ttNx8JmMfQxTnLebLpEom7p8
+BMjl+iMt/4/DPEFya7a93hfRqzdR7DuHnEsyALbkMA9Cz+1Z6kJ+kboHhQkyu+UDLMv4BCf1Zwl
fTzSdHcYZ+idnaGvk9SLzuOsURpNrW4cJyR79CUTRzoSfbMZftaQ1DgZ667MitJq3ynmVgRh6fuB
MqqQ1R2Y7n42xSGVQoaxhTYDVVtyN2Ho+OQWXZ2qdIZf8eaCw3XTQvJix2HSrQSIc7ajirkCal3R
/WgtNwDGLv+/DBCIriGfrpLkLwPfebMwsxAhuqh0yrwBSgukxM14kM791bSZr3c0L9DSkzShBFEs
DeDG5kaXP8Ygp2r37kNAjmoECxStTLLCdR4PK4w4EbhUDXKdAz7sTUguLtnuWBbX+mC6Bxv3kNle
VWDuSSm/DW/DAJ6deUlQVXjAIdF4HEtmMqMK6PO7SO4XbsOz6DWi2pH8c/9dIuMC0Aj3lZLJHKtX
a0S/Kr962V9Mrm1h0tgJi2qNejahTOdJKdAoz8qjXCrt6nVFI5qV01vbTWw47JcemGGrJXBd5y9/
gQuVffX037llQw1wJxkOExOCIjjXLq/sgRJfbCAnw9B7Vn5rrUE+UKJlJuFQejeSTZ36zeEWQ//N
nagE2ZSbKk7ES1tO+/aKgY+0EiecaWlUexpov5gzE59yfoVjDXfAjDYupnfX7suXcKH2rZFIXEAc
6W23Wdez0+oLO0Mk9RwK1JG6/FdcocaalaeM9h2Jj/25OAP5M6t2UYFOQLPKiRyvhXRLXdny8569
3Ud+DC2cEM2alYzASgYRRFA47ifkSjyM2ugamPXvXZb7LyL8UX4syJBMySYzN7fg35g8FyGn0pB/
9+OPmWvXEkO6Dx829Kna+2wBI1XpN0Vefw+AydVu1m8EGe1Lv8f3W2vrQkP1HrCxwsqKcd8UuyY6
F3RF5I/F4iPoP6CgDDmUAiMwdlxBmT/SYoIsBXNZpKzwSbXTzvbayE/d+YizcAMt7giivJr9VlXm
O0JfsIin2LEcL3izKub5N6HYeETzFDcqMcQq0DWh6DDJdaLHczsyla7Y2YfyhKUkrdh+362Mws9I
mUz114HdAoCMm/1yX9iH9bnwrYChzHTln/35IYoUhwAe7ZfE4YPvBlENTGFbsAHwgJeDlzD4AiYu
FsuYchaqKwZ15nSeZkkGMnI8aP2pP5A2lEdZkiqJ4GRgNw5sg6px7yaLpk5xI277JOG8TFyfq0y2
TTcFa8lHvmS+abVU/6iXMq6/IkNY6Nxuh/W7U/qWab1aRLmUDBHVf+D3IP4MIq2aVFE9RZScXz39
JOonm2MfmtaFUzxA1KwMlEofK+v2vyVBWU8Lsws0RMnbsRVXzDhbfL+khcUPH52N6YsEdwEwKn6m
UY+dhaIHlopzZw+nS6PTHYvIrJq5UX/TDl5qNHrFxD5u/FOuF4mumb7IWAESogoWA1ci8R1Vgz5j
EpkT3jMrwVRpRTeiRgo9zfqf0miPv4sN//5Qz9xNMVOZNjoBVVHpYpPVLFi7oI5pFsF9s/WCrN7L
apfTb8IcK8D376iDHprVv8jGGtfpm9j9e/0Hdk30CZxsDh1ZY3R7WfmZnvjVj1eBMmD7H6eXCjJC
LIv6HHakc3ywSml0zmoA3hDt92xCzOHhDSQCKuelSQKkoQ9nd9A6+IVwzcC1A2DiaE+pUa3kkBjb
Z4C28//aFS6dEO8z/3P73qm+bN6ydQKek6rs5uwgVKYWSbwsxwK4dDCkXLNpzT5JorXw2+TmiJ2m
3pFjLMb5Muc0NVQ+xo/A+eLMPcv11WXAgesMChAagmeql0+t0nBqhRE1tCalWfDPXo1YrSzMGWyO
JhBvmHAXRfTtn+WZMDzIZO22YI3X25wn2K4KQwShXg4rcQnzxDXI2NUr/atA39HsbWUDn+f9qbfX
1z8UrZLN1MO5fsRBj215tVgjZDMvWB/WvhXuZ1cdf85E3GTzVGA1xMaEgz/Gsih4g4NhP33+FRmF
RVDFza4jqSPlEHI8wZ+nSx6m1GMi4+BjyVLVHIgzOFSOkZU6mYGFB9fWs0YTc478I+XWp0vKQUrK
RZ5ZWTJH9g6mIFnZACN6WS6oPWaNi01c80oO0hlZOa//rEyHFiHmVxYaPSoI9QW8KdcITot67TJg
77wgc1oiQiUbW+k+5+4zE86nGBfR/TXP//9wYTS3VNvMUyF71nwd4P5/aD3JZ30cKZvVGvx8t/ZF
TITSJcPvFo+ln6rG0JxHvUuAesrcXy6e8LHsaITJTuqByOIlxukb4KT6VLUbOlZpEPZ9a+Xu4hkS
YZ1AVTXNlOCcgDIRppJ3+/cROXqM64LvFSRStuEzJTYdpQeq8ukVrE5RzFBod/YqzzGz/QcukTug
Jw9QrGZTM3U03vBy9BGU4gyuNdGuufSunNoVo947lKTF9sQdg4RQ91qkeqaMOIJdKjfY28Q0PjIg
0xoaKRX75RV4942c1yqgUw1CwbezjKcg47jDN7xQ+afVNQSX8YAb1u4icB4x6cAHgUcWAYFqjper
bFCdg/q3LfUmclFY64jtgPhHV6/YZvFv9q+9OzEs4JH6VPGIii2JCtZBV6jSodjEnBzk+nW1u38c
XzOPgrUp54B7DLOlcPIQO37kMOKBcN4Xwb062w09iNjX/fnAcuc46tNJGkEC7uVFpOgDXlKqG1iQ
Xs+eenJLd5ufVggGsE8KRNBsrtWEcco6MCrAVvf997fctp8Ip+pKtMyeVNtR+W6VJ3Xyy36o8lOx
EZ2JRoROadxrco/V11MqDe1MN+RRITTdOS+3IBpPKoHvrHmwsWME6yeEg/hv8GVMQIto80dPyZXc
wwaQvBrynDzhkhB9B+pfhzAWBZVQpCxVPkO18cxy9e+VfyAFs8d7loXxZxhNlcxIxuhSteSmH2Il
fag474Xp4oRqGlJww5+D/OaFhI7k6SFxrYnGFCRUotrk7aHeK1cLx2CE6IHOdx7iDkfRs9DbVEWI
C2lD/rjXkW5Go1IvKZmXFS3IUyv/2l+WlTepMV0neWbnGdqrdQRW9MzmRf2XDL9QnYiZVM5I/W25
W011jcjSLMFHLpKQqPNLnr9iStT2uZlsVhk4sgTSth/PIN15dmAPfMKpNkIMbDaO511GykPUFQwr
5eMm8sWh1vhIPDGkqgK7q3k47MYRjAvQ3lfDjdHCNj42PgpL/mND2YRQqz9Zt7OH6kJEKuvIou+S
xExwrp/yUxg+1QyDVRr0hXDAvYAuYPpFKVcpzOfU7nvj03hBHkS/zgPWypXn3KGraTJ2CkmKKOOc
AOIg9ZJaabxmAA/9Ez46nuQ+3H6Y0rtEt30tDIPqjw1ZZ24XAwCk3UTbwPbWg8qv2gR9VhHHLYik
TfSb/DsbUKdHLuqZXUAfGDBIYvzq7jb5lj6zx3rI3Rz5X1r/BgeInlQx2qk2lbHFg6/SNH0CaJrb
CiupPNJnHXb8pfzwobS4YjC0q5Y6+nt9p87JoosBxbojfbM4OVD6kFEh2I5JscCY5SGl3HRvvwXN
kXZ8yApCftBHjN93WNFzQa5dq4vzYPF80b/eUFhRVZavAH6bZmGxDNMfYVDC+8ccxzo7Rw1ssEbF
XT481Bft/XiDEqaNKZCP6YumTigvZm8Yx6kOAhBt3SqlO8eW52JgCsi95mhw1ytKJLOADeklrLjd
sIJVHMtbNXDC02GmWNf/GTKyDdf7sDHVzs6BYCDKwKRS1od8kLIpf95daIsu+axv55rSsdZ66bYV
jfKTLGjgkCIGaiBnJC6idAKQHRlAUiqK8VetFIWtZuNbV4J78vEf2nQ1No9AvEsdmgncm6L5Q5xg
xMH9IGthNGDgWYjLfm4f4AHZGbMFB4rmv9VKdKCEBXLSB0gBvxUUaRT/uRinfp+seqOU53Gr/x3k
QV4f/QZxUMZiL25vO1EHt1JnBaeRdqx7IrlXdvgVZsKLcYlePsoPLeKBzKgKe5gGKtPzQosl8il/
z2Dm3RoTHlHGB+cbz8E8w5l/4O2UAYM7w1NmZyVtib/6KUtUQsbANBBcRfnpgqTHSiSFfkkyk2UZ
pYClmaccBH73amDfSJQ4Wk7frz4P4R/ZucQD1z/sFJdYhCAHcpwD0DgDJUXcxWIQsKTQVIQcfjWy
MqANeY2+VnD2s2QmxS2bjhQeEAifjDq/H2WwqvqHPkUMJHK3XGnIwAD2PHNl3Njxtq0bgXhLH6wW
rLPye8BrtbwLe3o7zcYuXbtbruaQToFsXFxKTOKfLnPyEJNYaraJaGrONjFVHfOKQx37EvrXBCPj
YzJPrZZ8NCwpcj2KR4SVruvN11XwfVaQ/NWo8wPsoKU9uiMiQjKM0ZjevoK0fZsfr3xqzQRHomSe
0P5qS9sYcDaWDNjHif61FMk9k8pfw0ORBG1cM92HEn64GzVXhOCAbl5fuqC0Xfot9VfuSrLPjjk3
5nIvdGrY5pUE3Aoj5yG41c1uyMM5g01mY195nHIan9js77AluMhqWI9n0RJ7alNfLVVgh8jb7wa5
YN2sw9gukDrxxxDGvoBnq5HPeJP3jQgEfXoFyoitKsFaPR7Mj2xhHO6lvUtFeOsk74eTDWDTRFzq
Bggh4z1EnpDmrFWOSgTLGEcfV6v7B/2ZXTt+bi7ddu/QEJApC9uG3PwvSh4EJqduzRQZ8ycsaxx9
RIzNYsDC8eRMIaVonmvaZxhCVdt4ja+fmfiu/eZ1Y2k/2Wa4IfHEJn0NVUB3hPm28kysLla+bUwt
gJmoT66iHiDp8HTa/zkO9Yl3/jzJ1KyothycEftRnjgJwUyeO3IArsIsizOBHeS/x+Kk/rxxEUSq
gct2RxQLJ3HG1xjIvETmXTtgENqZmHJIuxjc0DpEGfnc+rjgY+0BmraRQHFBALnsgQ1zkU76o5Ei
au1K/DwfJHGbi+YnJjKQ8W+ALhNl/gql/Zn2ipUWhunpoZ47XPg/ZFTHKZNMlNxC+nb5bQTLgfGJ
Z01FDm+tW1XnATvJIL+Og33iuxzcT9kYojGfjfAxrdkHXkxZzaHgOXLLLeBuQwCNzCZPy7HeiTXi
6tXUQIMoGWBFw1F5oHEkYEYNVKy8y4PCdT17H/Q09rkzybPf0BGioj5KqLSqCRsog996h5eGsZS8
jYxq6ked+Z2msJ3VmCOG8TO5vWFPiYwWH9JS9ANW7bPMxDUXLYDGHdMODoFRzINFNTFDolRfNWU7
5T/09fA3geZUNIqqbCAfjXNYihW6BBuybTu+uajazb7QlIJYP+LGFKau+5vaG4IY9Btxs7oOKthr
jUl4NpGLzvFmnL35TgON5eTZp5K3lgUC4iHR57k2l46zTDInEpqIklcxRYMrtmZNPe07HipRX3rz
Fydmg6ko7IUqoH7pEKuCXe8P3DBRyg5psrGC4uilLUFm7GNccDmPeQFbjcEsoCUf1lfRTduIJrEj
3JHGo6U32gHTPY2jxJH+l+/jhysCdeRP97NKCSxT1SnPfCCHUQHAu71G/gSk3n5Zdd+V52ZacF9B
c50p+k5euvQ/keEvQoE1l4979ExZHIuzGVRV9DWYoCvMcS90Zht1PWzYYcLiqBbcjoLiJhOKerQ+
wZB0QmivjJNltoRhe3Wx9PiJl14sz6Rp50EfT8O+kounRwza+XjkEYYT+E+S2sp6GcKFqI9t3haa
FmwlrSo/m5eVnqrhPlQOYNc7aYDNCIhc47/KcO7/6tqnPxbObTqh7SBpKzpuV5o4t66zNry+mURl
o85WkRbtuym+P/ry1eDUN2U0+h/zkGsvgTV/fUAZReqO/Eo3ItwBqalhjDnJXfkygP+TL+c1wRcw
ZiBJz1TaOfZ99JKMeu8MBiBB2DJmWpO7/wruAnTLDrR5aAvqgioYSYFm4VHSrQsFl2SIN0JPQ+7x
5qSpU+SVm5Nz3+aiiF49teJxZSZPUTgMihcKrvHkmUE0XqH6Yt4YLlNfeFUHO12vyg5EX8DHIHNk
8Cp91ErqGZ7UJv1c4+3DwLr+Y/QScVUKXHkHsn2dFV0ow3Ee/rm9ZcqKFK8yckzEizfNhilDor6J
X4RooOEaUKIEfoYU5loCkaCC8pIOT487rNq1BhCNNxDk6cOnvojXk4CHPORCWwQ0f3xm1OVWLMyQ
dwuICSve4852bd/ARIw/Ypul11pDinD1c+OLquDaIpWcUXYBNk26cQlfxLFQdkq3yVdqBbPyINnk
W2EjOnezEVPd34PqAcTDUmaetxGqP+14c4k/+AXspIMzlnyl4jGmvmvPk3/hIboRuFMJ22aqbbRN
pbt8SUEPZt2tORTSDqwNxWMKb7NwBxnwUBVSK5G0TlKicB50nWCknefZtyBTuuvyCQDh62I3Qn6U
VkVk9LfjzrtZgVpQ/4VYIocyvNvThATemHSKxqfgWWL1tKlM27fZ62BIrELbDrf7c5yzfoOrV31S
ywHNAe4fxxsWprHE0Mb6vVL+2LEZE+O/DoAuiBQkUh6yaTpGQL9JLcQMM1U7TpKgX/s5uZmpvX+K
Zgd0R6jtTogh+gl4X/pox6wvGePE4NBerx2DocTsy+3HSdiYSPUzNmLueWM34jCT7POVy1jEhv8B
8KJtmStpov7u6RwRuuYRye5h/ZujrClPYzwgBf6yr+voEGe4q03+QzvjpCPSsIbTS+wYrQPuBVkQ
kVq6VV2B0dE6WtLiaEE6+NxPO5xtQqGL8TrbqVLxQSBQZHsEsKGahAs1KL88JA61OaPt+1OooRz7
Own5ygwqKpLsw6kHz8K0TRkiMvRAxefAEySvyfgdhHHSoIp5axIEAuonMNeaCFaHqNdo155uHPRG
AsEo8Lbdtm9TFyYCbtCe+nt6eLPD7WnTW6idRYwIfEIHxUvc0TzcUAEeiml0i77NYCH4VBzqg5Mg
D5215eS4f7FtkroMwd3yZ5FdcjW6iSWKxXNFOCfPOOT4Pi0dmX9GnlaXbJaZC/7MIG7oI53xINfq
fIEFMd14kD3zldAnFug4wgjgjGqG9SjlvfFaYk8b/VJf69noSSPgv3QSqrC8vp57jIl0HataqXV0
nw8JU0In7TnZs3vW3ive7w7rz31wv3R+eoAWfFSfIuPgxWy2b5wbvIg4oOsf4kKd7U/c5MLYsUzF
ldGH+i29NCt5fxTYB5mAnXqkrXeeaK95jpsLxERE48VgTVHjkCwAD+gS5QjyCfurhSW0Q3KNBtUK
w3cU7cwTCsxR+QnHOmKZpwpSsnQsCatQxoJHwMYWd20OxOUaSa63ypvtD4m11YHbmIedzff38iJ4
NGvlo2iLtqO4WXseKfDtSW5CSq18U5eDX+SbPriAocI/66z9i6UauU2EDTkiEKWCGKyxOySum0Yy
OzeUat3heOg9051zT4Ef085IvXf1ZqaXANEVGpoqiMXB7dv4hXYhA8N92WbHKXxaqMNtk8FRq43H
6hjvTl9LiIa/fm6zugm3SiM4+r2N5iHOVN/QLx3dG3MD4b/LOhOOS8Y9aFKYvirT2CZx8f0mKAZs
0DNhjirV37oCQ0EEXne61kQ+byyTjqPqJ6DnJAR1sU4e8cJaPDJFAKKfy3m/UkC0ZpLesAo1esSm
nmSX+SZVL0Nx+nS1fOsgcuz+Vjfg768fhqE9Ac5Pt5ctw7cAgqwWkVKquIlGTHr5+ZBj1nHGM/FU
K0AGWjqGxoMYS3XvpiJ+uotIUGc7QhMA3FHMjKhKn0po+a0+XPLnyKTkqROVEQiHM2umPsGO/3ow
LRvT6kn+h0Bq1Uo4cCZzsVhy8nNLjAur11bL7iLlS0MJggmUXkNO+LDoIoT63hzWLfC/hBgXnqYg
7E4NsExxa2fpt+v/jSLWTCJKTUpiPHmQWDeP1BvBKYcDNGH4MwUhAkOCp7l0Ta7ZOOvCBfG+IuLQ
cGrKyv3nxL5A5Bdd8N4WR5M73lymFqBAjSe38fn2CtP/DRb8qQb3d4iss5O+LsZC+Yd6dI2Xxr22
2QD1yXwIYTt46WADJQrONFnQrGIGJAUQebNJjF32JVzNtCE3QUY6y2FEAcsQOuNRuYUW1/Eh0rno
CtmRdCYI7fEQAkUrbuvSsz0O0DYML6ODLK3shCmUhKt8jAqPAuBCmoypLRTO0egSAxVLbtHyuvMH
7ZTc+rWMcu4UMysEYuYM07XrS4PDMxrVEthfmcbE0I5FKBNVD2Uy2XubITvR/ma2gMxQut9j1W13
d19hTeungbja+i5D/1XFNaCLDyb4EJ02yKPHTRAyYgwPBiizrltNhKbL8aK4DXSW1iB5A12ZB2qh
nz0S3RvxI3IXVaHTv1tOxY8SwKbxUB2oCyI0rlmvXOQzK9wXMQkyUjvWyYcQy2/NS2KQwK1gTY2F
Tlz7sWu9bch5z07oqPAcYSOehCkZVJqFMpmq34KItrlFwTD2optJAmURKwYSPAlpTrXI94im5Xar
wwwtf7h8YI3uT6Ow1wxGE5KFMQwcIBoRUGZ/ZQm+YGa06hc4PYJAjs8e/NBVZIUZJWx3V9/kexmG
CTVonlIxJVnYlQ4l9KBZUuQ0V/zpOQW7Fc/bgrFiVPoRVdp2R1Cmu3CZk3t0S40zfEKVs4rYDpv4
8O5UcVSC+f8/LOF3kp4eyTsoeKAKrTdcYHy+CQYBCpZ0JlUJFPVVbau2BqAPJ2M13lRz5/rqoYBA
l3yDUEywquX4m7ywNluLZG17ybUqV0o5/4E+8fHdXipycYGYluRlKAtSRRYu6xCm3eM6KHBDySfs
CCIfgZfTUe+QV0pHA4UBNiJMMdtzH92pXxyYfYja7UVEr4nda+XjFe5cx0jgvh0aAmcCuJMpr9Rr
f1aGt5sKTQAhlV/iMExDTFD3P5McqQuObwnnsfd6YlLyNUxG8Um0zMRIZuYI7mWO+yxvpS7zPbkh
iQWdlMJpOfLmi0Hw4fglU6v0Q52tZKW86Ilq12tVzJkL3sANyPGLmXuOcnJuC+0nR/8/LOP+7QDJ
cmOxwOcdLDkFWABeCnB7/bfnm39PFlfjT+YmPnyagPKBX6b+SzXRYxHl5nGfZsLbnYgA5KpdoJnV
ma4Q9BsIzIkWd3zJcuu+QbpPQGPDjjbROJ3G0NhLyFy/Za/HdVBhSspOf18DRohX/ZxCQatup0mm
MIeabE9Akt/yFr+IRWq5B0BvMQXlslMQs4IBIgEDEx6zUFoKGHxJy186b1g1vnELAb7uriNC7pE5
Y0fTkxYhJQxzdK2E8CrFUdzByNcSkAwEx99eTJoZcfQFXFR1ML/9TfHchh1UDKX+DmScWSJIY7sm
wXgesY+buWS6y7uCjM4BTJQOoAhHJWZMNeiGufJ/yxiEzPXj6CO/pCsaWuG3ZHXLAwjakjb53vDs
O880qw2QgAO2fQQbhuD6SiHmmGUvl2ZFNHO93n1u4fEzUdLIfNa90mmL4m57Y5n6trniArZsprbi
Cmo/ie4nawOsp43+iVcrkWXBas0kLv40XCEqZBfXlc7Mv702A+DnanUlYqF6jQ+I+RrgbpOVMyr6
N19d7woZm2pdLWS05e1WEY/catIIDnXuUeP5f22IBb/PBpd2AKZj0hfhXTevGw+EXLxvJfCjwf6F
1oEZuVvkyC9NMsvwpEai9eFc94XqDBIENGAV4RyArhZCu42KRGagpmu/wYz9vtI/gEK9ISrTf/kX
OABOI2yZN7xUgjibFhuJbCCtOHj46T7/V3ZVCrd6M2zSBOvzJ2zolsvPDcNMShUuxmvVvSHHhFJq
BcCCgLsjhSLsSnWLRB0uLutXiLayb2z7iwKg7+uX6Npd0P2pxddnk8zAGGqeC+QMfycG54lAs7XV
Cu33OrvT9OWwkn8/sKW/T2M6VyfQrn8kHto9zuZafhE9aroIILOYp35FqQuWulbORI2bdME7L+so
MXHNzwQgP2PUcIMg9Iw5W6R6aOhlNvOkJx3ReB7TjWBJoSf5IYrmKEY5e/JXaBKxykNQC2IXa1UZ
UmBVsQT7+j4/hD05s2P2pl/3fBdTCPKSC4gIZ3SZeZNquUngpPW9Dcy/Zhws5ZXxOKGTU+vr0Yv+
0UHc8+u/uQYImuABZKXDtj/kOWcy7FubMP6NyPMqF+u7BqB/UqDWQ9HdRZ1YQfY16cVQDqbKXkPx
LXGvpTzBRPIINISGhZeUWzVj+F6aceH08hL+fFKnPzQTB9fjFWxjJjoG8cdFJ9F4AO5aurDcP3Dz
Qa4a8L6oZfvHW7sr8b1dE4io8w9BF32NWODLfa7MZGQadhi66ixN6DV9BGrNn83L6GB3m0AsnFSb
Zhs6Cedsyl1oLaskLDhi7vj4/5K/ur3ygpOgJV42pYs//kaY41+njYTVDg6qOlwE/Ffu19lI9oRt
ulxRmzolBxa9wGVhhriThvv0lxjA1PLagc1T6xUoaXATCuK23MuELX0Y7qoNSia/LxdI1+6QxwWX
pA4QZ+D1g4ECTb99Mb2xQe3qu5Ww39mHgxUJobtJK7sVPFbh3lxQ+6YBnn/ziazE8UN72DzQjld6
e3fy00CwBzpWVJFP5pre/ul/P5dq9yKxb/lmBEzpG1ZWrVrz25zMVv0B7t+pASr7yvpUtYNk0oyp
OQaYguBvjg7JYUtNPDife7ErD1GtUUhOtlvgGGr2zUlkr9YRt/lyjUFm2ztUJgdYUEWuTsbfxKRn
uv3Fb0rmfx5vUJL+3/b35pmjqSqyycRH39PARNtqQ2s7FiM3JRbCNHOFN5oIA25Vshyx9jVymofP
iKZ5KAboCiIMomuffHqc9SvsUYgOZLX8pybXCPYQ0WTnPeLv/h6fkXmG7bkolTaFysqQQZAUv+0H
ji2pkwzTIkoKzxsLMrdlr9w9OOLsqfeBbbs44ulOPEirDUyRo7Lj0X6oytrGQMEV4rUkytM3ND8x
F/2uOqhJ0j83CGHOCYUaDtqKtyURlDkqkte+TCfv2gpsOlr6YEgAlJuvB4p5SGTMvh3uWiXgOB/S
qBExka+USn/QcqWtNeB/h7L47eIgMEMwARfbP02SZR4v0sTaHiwm7dHjsloWwMc9zx415B9CC2kS
tL+JrIQocXQTRXbCrjSCchU6gUAu2ohlmLyoxpJmhLLUjd7AFpMeZh4zgdn5L5h0QVvGV1nQnhG7
0aN3B3Hh40MyKkNXGBMDOcZB1K+vifL6xC4JXB53GXeJcMWF3yggRoCuHPF5LGA+xzay4zT4Xf8Y
Ai5yfFkpEu7G9/Ip3+k79UGsuYqrgfhjAq3sWnfsgW1dElMltOrWoosjfrj546vNdgTTeSNz5422
dptRgNmriPjrvAFNJ/jBAjqP2XmLUS8O8depzQv1woCCt28vYs36Xcj+Y26AL3plcPtYqPWzcz91
YzlzOVgRVNTwz1/0GsQNudzsFjP28dx4Tl08BRe+fwT/5GlP18Pj/ZWleiK7Ct3+nb/uQQk+76t3
HLhqX3v3rIqP3IuZUl770Avaz5p/x7umZOLY8RmjdHPrYaueNky7hRnOXxIkdvNmq7IZuBUGFuO0
y90Lo4nayMhm/ZH/STuiqWV/WTcBAAeocZsjp1Nn7FixISHkgTmmcIRKdGz38m4nwQRbdSyxh5AD
fDtXwEziPRl49YieBpoNszdwBzVAHe+EYl7DOzLlqShl0DHkAxuO18EAOwI2dp/qNDGUp98pfEsK
WloRzo2WHNtuQa1RJiMQwFvU4At+CHPU0Eb9FWkoIrO0QzRqE8UApUL2jJNaLJegJe9HFoJATYOB
YSCJAeDOowmMbtYsO5y+hOuh4hNdA/5R9pFwLiGWajxoxrGMmzHgDhRXS1QNIwFYjAAJX9KblDLS
Moqf/2J1moL9vmymqRC7jTRkM+lTYzgfvshslJN06HnNpFS6zzOGu5qGCyGRjoIiRIBWMQRCpvQ+
WvXV0yrAipcoFrMPUmSPoX5AyiqG62t5QJ5/fZ374TgjX/lwV+av44zHop+kQAK+Igu82BTcJe0i
/+fpzOlbNhwIMg2LAkDUy4syuH0NxqHIvvlBpzpG/PzY9jwOB2aOguB1YSu+STQs2HntuZ0GtcMO
8JiTtR21EigQfwqsAsPvzajSRAn2i9jLUlPRzN8hD66AU4kJdDDHlFUgoQYLG1wkTGSwp2Bb/LuH
gbyQgIq2ANARDbbwcTGOCthw9fWw3KbRxSNXQ9J2PKpNBO50QodYI2Q9jU3ROC7dFibhr6qVPU2c
d+eaLdcGLmeBGahnT27+CRFOdisvANnxqKVP9Q44hWcu0xsEIEqKut8ltwIz0o6uq1zm+6MnTP4q
TFHPUkXzPECGsEAHpbl3ScQb4CB4Frn4FF/m4kQGUmIc3w3zFUuH2TeDURVr0DU42ifsQp7ciXYX
fgNyZ5ovIotuPCzu83E6COYzgkN8X+ibLAZ2IzaAxls9Ph4ohJxWLLXhdzdECkmQXhO+lxVLPOdb
x7KQ/zeI8a76pcpwG9OXxgThnTmNZQrGODeATjlvMoRhaVBRs257nTEXw1vuZaNay5TnOlM6kCbu
xmnnVHAUs1LzZ6hBoO3pvoCS+KDH9yOxe/jtrD690jCJgIayj8fBsOe8cWntR7D1IL25sjI/fGit
MAClFNaTyw9iWm+xEwzlp4hFGauNTtUYLYqwrae6Cp9BuWiEpCWsewGdTPDiUJa7aSHEm+BNN16U
OAHJipPWnBtybySYyBnEZryr8Vd4AS2eNFaJcybfAXgToEAxlXSLPBonyX0xHrjIUHicTASvxGAt
/Iq5IMtDeNsXHNwjq3iLYzUIkAwTsbc8ULGTVMLMpsJcDano7WSz2bacq1BGR3lII2vvWUC86hkg
bSAPCh+4zCTobdwOCUH/Tbf6HjseO7v6lvPdk9/7tPyGvj1mUMrlelTXi4JluCFV/rBSvU19PK5A
RzgguCXiEZLmoyM5hli10pK26LzPSFtSRZInx/WlkFKmPWLUkinFihcpbLuUj7JZxZj7h9SS/mWb
/HO0HHz+cL03eZEKrF/5AiX3BhCR4cCkeVRBVh51lvjoqe1eqOEMU7DoAlAtC3+HECQm5gTXBy/7
JCqXf2utlBVCeeFs5C4jzrwctAf9SRvCZVW1ld/gPCnXm6RL+/CTxkx+IdXMJLSfWf1HHP1ttVe+
hWfd5edetLfv6B2F8R1gDakgGtkvkji8QBjC8ACS4k4zGGNVH25jhrs06kLTXhHM2oCgEES6HILu
DbhnUbvWWlQC8pzRpNUTRUeHstoEB0rkf+xLTlTdielaVly9cLWrE5ufhuQVNjGt6XVhOe/bjw9T
YlLnUEVQtJHsF5aXN0u6wnyy+W3oY9+7DqBcScTth9+88BQigNysGgAS+COHjB4Np0isc1tBl8TX
ae7JT09me3wxBFQCq7zE9T4iz1dLbhTxtQxi/mGuqmQmpC0NOow+DV93S3d+LpR5ErwggeLlBEpZ
CX0PSle0E0MmYWHUTUm+Wd758fWBynHlHK90b/nJNJcIJ+xhT8AW1yAsHl4maAMsP91M902+Skp6
GPjxIaHzl3F0baqFKyHCbrznZHoYWLmC1tuLvTRMg3hXpnplQ63BGUX6RSZeBOx0vHH4ygtjZMOP
hJTGOuSDsnOpiRq3ROSE4gyQJihmCIwRhxIyarjJP1uv1pbQuwGRV8t+t9Du5+XzfDdRuG+TKS8X
1xGTA66R86qlZs6QqZDdwXj19hhlx4VVnbmorJttK5cx2cxXqQnN8oIPV9cCH3gl/GWHkOfBox7Z
z8g/vFV3IFeL4MmicpuNuiEoQ5w9QyDmZdy0oFk9sJlKgr9KgxD1hUKrZJy+wIjAM7JGNW48zhBK
VC/AAmOOnYe03qvt7xuvhBdaSYHke9N1UMC9JTFURy4ZI1MFIhct7syCkfzN5uSWFomsOpZpTOFo
4iElTLuA852w1I4A5P//e79b5fVlCuHe1WD1Vm8S46BbztwpJOU8+ynnLEcQB+qD+hBeL2OFFdT9
VFKa/0RGejwYXzkf1bkPwyo9Vsl45RS2UeXq6GnXTx+qIcXr4SF2GksC5u+uszFac9nDUTpqJLok
KCI+Pk7pMXCV/H2rxNxIktGSLMy+9kRJ0WUNJJqMsqV+T89FgnCqk/gMW5HoBSbbFBlDpF7o8ONd
CWVURQrG2urLOD4090VZdl601jH7wlKAvNWSZVeuyX2JFpDXpieilwdSDdkhaKbXebsUKtRZ5stJ
aF7t+VpVS4J+uox6KjCiP2WHCWGHAA1gZsH5eBAXV9AvjNOq7v1nxc1KtgVCVJfvogf8VsLOmpSM
Nb2tork53TeC6V+a+JhzcqckdqL9Y4TLd+Bbt3HdoiBMBJZnSuiA2bH4V4u9BLXS85EMh4Cr+d98
MLUAiTahInOeJozMe4NnOGcjJb1rWnPcJMeKIXdjWUJ/tm4pofjD3aXRuxVRTkHn5G2DLlogDVe7
rm0q/5IToC2iD39y/jW4KQJ6mqB61h0lX7LvfNL+hpmJoPy6uP7miNtjWpCwjyIDwTSVK3jMfRXE
0z5dXF60ZVd3Zv0dv9FXiurKmGO6SA9gZ8Dx8Bnrc4ll5APr0XF5Mxb2g7F+K9x8SKroglgXsshW
rSzI22x2kxIOA6olbb8Zc/2CAVpMiNbDe/oq+HNuZmpL+K2/VXsh8j7PvWF2aXFpo/Za9kqq1Aup
noq2kIHP08qOBzvPJdVFmdS7tfv/kGWEVXdhQwCvoaVtmqr5VOOOfFga4QGhnE3C7bVLwVI1jcV9
RKQmLuaI/+1Vc3bTuqnDZviOY7Rf5vmudHkxtWo2K1tRa7ohwzH5WVoSyMnRyRyy5Wy9iwPz8nAn
j/m7AY08cDUQQaHU+lCEzxiGfYS9N+NOnPpolrbvwkpiMlYNAv7t4IPMK/Zc363X/noW8+zzEyRA
HXRjCJkjvBL0RZegKNRsWgLUrcFEQF80tPa07P1aeWAXM8WII7vUa2cJtaC9uBIc6XpyYGzEQhbk
KAfPdNWDj5TEOHYQkx+ip55cRViyRwhpRpc8Lb5+xyEvkT7MD2Eajf1U8TMpmu9tk2QzHqClZSMA
5RToev/89j+cWaoAdMpWo84iTGTcO05h0SWrkSTzIp4faFZlmwOgYU2CFNlwJhROoktpuwADBjd1
0JWxoxpD/uxYx8Kc8QfIf1n4AIV1irHAgv08J2DiqGKGX3cgkxz0nAfP5aqSYMkq/lfqz3JI8f9u
ThldeBWMd/bjM4H2xLN654cKEkeyYK0ZiLABP6y25RbmIqLtYfKFIyTPBpQVIAbQPzt/OPFgmtOU
C7ue+Az3wE9yppHG59e8aaMkWa+AamVsDdE6oHcLyywb4/Vel5xp8FbLzu2hQQDUWc3OmocWIi3u
QehZbB5A0LmnAhrtQtLwg0v/TCWXJ1SS8fEESN4LuKMc3NF/DIIqafVnVYw1zN089TQTrxyn+hLD
S9A0Yac9wBBfdYOwnWZxiRny2lfbmd/Lpe1GM+1R23xE9taeeqIcMtxY/YZty0df1Wcy/K7kekxr
D0gnUlkHW2N5dIqW5AoRe+Hk9PFmWZD1JClu5iDQoxw77sJ5tn3HpDOrfUFFSNpUQkqKurb4n/83
OicIosaBKflXE5SxG7TtJYg0ObExToYJ/hEwAC8nucCQJqT70ZtsDNH4UQYzO/LJweQQfpWi7YqZ
27AYfbyH/4hhJPPHvo5/A9BcN4tEVlCgi3RM+6Yc+jWLz4Fgas3foL7Dny9s0rsDkoZwCS/pFp1u
K9r+lQQ/X0nAVKDdXhefc3+TE1Bpnd33BaKZCcfWywdomkae20nTR/TbMMnq+A7kLNsdwBdUgXzZ
inVEWnT8NGq23RbbTwyJ2c2XbsdTDB6hEYFgYoNwNQBiKbGTAqY3mr9zZ/8bzw7RTGDp5195pLyZ
KjmlrhosaGsGoE/+2yPlCIB/XLqw9vXcSvICqoGXUh/og4DQV5XSKoIuitMuKC3fpL4UcCLtlXZO
6vQR8fqxLj3Fn1K2CxyrOXcjXKu70R2qCxfSltNq+T+3KKaVrTOzND4itQJxH7W48nK/4wa0EpmG
Mn/nn3MqzQCn+D+bhGT4qfgK4GXcOL4OZ9QSQJ7EXeD3yAbj8cZv9Qf7CzbRcTWEE9IL4BSe26VB
tqM28G+QNvCdOW+aRbO2tfDaoxs3IZ+aDUxz6zEbkS04Dcw8eWh+ohifUZh+ijE1rDX0vFZRpF4R
V5JsVcJuytk+TN0vXwHMxCJhHZD2n6weAwU8SWCEOSyjw80kKW/x41KLIPvAUWEz/U/lSy5dMy38
vZ+POj3v2iEilr/4yQ2wCowUgv2N39hCC9uNql6XUjr6HrLGOMISvHEM+ZVJd98V+TiG/0dBMJa3
7PypHWDWEjsa8d2Fg3M4vkMN4WfYYIfNici1s+kTEvUzLA56PiZ2/+CDIXwHQFmYJvlQDra+JPHB
SCy6pmwWWnDDd4gzzVJdkABQI+aj/DI5MJHSiHeLuhbrkE7R2+3nJwgw1vf593AKL5uVzKvbhskc
GhqhwAgKgy9xRrppHyUFUxbZaEURNshT20PYHaHcCpGVSHPGkfJgGo1b2lv9jzZ+GY0cZOhyQN3M
Rbbdjx+Ph25vM+/jvtNcRMd1sDQD2uNIrJcecMoy3d8RLKknvm+i3ngjej71lfplfm+Am1ILEU6k
NBFVV3WZcS+GrB5mz/mS0e9AoIjbwKVObWjV2uyWeNWKPe27fXJphyQUWWs6+UqzVU74FBuSUHya
t91WMS4XeKWKAE4dRf/1rzh4if8hceqXxgC9CQ8dZ6M7qsspFCPkeay8QKGeruWyn1Ve5SGEiS2g
Ox1ZstBL7qZCfUBqqRgVlt0JrdNyJAsU7X6vKGyvFhREhoyt0dFk7fqyCOcLUJvdx3cu6NswNN6T
5Chw4CIQoAVydUgkYVHlZwvDAb/BLT7X0KWO5KuzPlJT2kvO3TrT4GRLV1zeG+eiBonfvcTl0gr6
DVvMF6kMVSGsUTY2GicnEOkwYUjFiKjU38OkUtgfrqeOOxDrNYAa/yqJRC9mrVHlrEUCbyyTB6Aw
8n9NFLzZd5MWz4OzI1BoaaidYZgWxeIsm59WygvTsuZQE1ofXROR01OOhAnQZas094/U2eQyVETj
OawDpwoqU5XoEuLpUMOvWVm37+oflFoA9fdRlRvOHO7JaoTC/nwa9sfucZbs94CyJ3hlBuKrSAG9
li/mDxE5Spy+W7oM4GL7TxwKkb6XO8wBj3gbLzL8lY6G/MwP5W2u3KkGSmNtjQu2gyoSzBNnQRQ+
nXn+hIgkP2OeFo5HbNr8xzq1DL1YBmM0lmAHN8cNT/Sqhx1hj/Rp50wf3FU1KQwcICNgNawNjwwK
i9Z+BuwWajtBAKXWvQsw4pmGYw9Y273jAXhMOU4j2fig9CVtOKcy2On3dJNfETd1O51oVFiQbJcu
IDSTxJ8wFKe52dE4iLQ+Bnwh1FPMcqydfHbiuXNX654HtxpqNq5yWQd9F0nM+rPE967fE+YI6+2e
In1ISACk9lo1q/Y8OTmIppFMrHQzmX5OdqwFaytl/+mSMoLzoILmIM0hwWkLBdoNGh0MsYS2TePx
H2mL9E38o9SMmdrOQFS63LfABf6a6U1xkmH2IrNjfYe8SW8uYXJdcfY0L9yScrdXwtlooUBsdSL/
lGMp2NvPKd5aW4S14Py1s1AyRCp9uGuPTO6GW59SW0IerIfheJsQ2hul1H62PZX1khZg429koGNj
RO+a96s/vH1gLR+2YHcsWwrq8K45FQsRVpIyQKoEF82ItNyE9KP+QEIZvOJVGKD1+6exYMtcEiFY
qA7op1qWB03gUTY76chaKcCDn9nCU3bm9UFsKjo2hxmQx11C1Zn9l0Xe64t4d/Oq9rGcNbao+nOB
oNOWpL8XDTITBQWYf+5avqsfB9NchyJO2rub3KB/Z5YJTOBw/xpJjApQoqWDFym442ne+1FtOZS4
x3nR2LSVwBm0YaHJefdvNP32/7o1kx3yLiUuylaQcOz5j4ugzAidMvVMFEmNsR0BGqgqNeTPVBCf
yZIvi5G9epqzgokQ0py1BegTqitkFoGW2DTbcGQM/hPdSeOgctdtrEsTQaTq/EQi8f0wGROBBC6f
4O/ElZZtoYyHYs14jfUf4Wrk6/LH4hbSze4mem832t8u44ZK9XhslCOmGCIFmT9n/hn4XZPg4L5Y
7287jqNSP08g0KrmcasQ0SJkS0yzd4dydTn1uh8WhKRkztPR34aw65Tsirg66iDM/DlLi5o2qH33
szbbTqI/e/xGXJCXdpDHZUkOdQ/ApU3YYMniH6Rqb4DHSs5aWna/Zmu4mlGFo8L4IQm5eFAxMtXL
Eh/6hkc7xRM8Se0/VVhOamF58rlIbc6lewZHvPG3JdQzgLEmUSlfjpUf8rYQ4JG/yJ/Oj8F91HzH
tr6KaD9rR1lVfivpCW9bvRWEmtxDxTIr50BWwyPdYfpjLY1p2i+qw5tZktan7se+xErtWCHoropd
cwAIoaBbawSQoqcEuVeRAzcTXVE9OAjNFnTb16GxRAvugfBUglIL/N5ObK3IotIE9ha8JnNFh0P8
9d+DoOtLNK7/2rTnZqIO1Trk1BuywXXp0yewDs6q4HvPLh68OwpJy7jqD8tMNFfLia7XgpfctxmK
DKhCrv3HEHUHsUPlB4wob9BHS+MgS/mZStdbiJHSx3HFimTSYT+tDHj+ugfFx7F2WFjhzD4mGoxL
O+oDXDWIG99WwRqKYK2ClqVRxoWuPRP2rlyzMia4BiRy6HEgH5KyZNTxm1TNbFQJOoUdFuxisV1I
cSL+pQXledEoE6qx/h6g64SHkujoz/fHuQroq6w1moOgtnWYmN5rnrkH9q5VEO1ZgCzZzYPbgg6J
CEEoOrNlZXxXI0o3XzVMOqGGs+ZJKNmSeYhN4arayMQfYs9iQVrbaBWd/Qr5UrZ8mN0y0qWjhf2I
FK7ncB+0NoRkmGsVZWn+YOsfPhPGUWwBUYl63dZBh54MvKzXAjr39+zH/epZqbjBRAC0APvqALZs
73gSP5B4mHTPOhyuozOSZ2o3yLDnUPOUOczmbJR8BPW07Pzqh2PfkqyBSn3JHMYxX2fM3VboFXwo
sqoNyiAN07oyg+vNmYZs7w3aCeI/R3gzZ+M3CH3ULWX52P2UP/JvrNjm145E1Hs+55wByQj0ETdQ
CUN+r/jVEDG9QqmoKRVieTp2BupdiSXe1cuAQh8OnvtE6Pji52+VI4W1Tj2L4pDnvWNgjHg+oTZV
TEXXr1qcViNquQNy3UWR6Cka6bIMaf/woCON5Boo8JJs6x/IQ3ZQ7ES7iGzyMGus0ne6GWH7s+uQ
iBnBn4r2w2nqs2yagb4re65novgW4BwPhHnK+lWBVm+GshmUoh9Osk5KVNc5MVPYOBERj98pPvRD
mqvWf6jDdeSG/9NAZqAXM3R+C0w1EH4gPDl7SAWQaQhZuPEaXweHFIE1W8F/j7DJwJlFTVT3LnPh
RuESwBGJSPPMD8PsXT75wOjPimkihvFhA4beGvd0WLQN7NRNSN6cMJhFkDMm1gEesY219Uzq5TZz
wuGTDTqdI0VE6M6+tBVidVO/2eP3Meb5N+ZeZNdcJqLsRoSn9md5W54hrUY3nXdWwCciCmEtDRjI
Ex7NyULsM4trhW6vwhyJbeL4nwoMTAvOFKr4W6pytXAr2ZGN+ZFY8szsKXZXxWjIMw4x58pt4pLe
27V8vtpPRGITYcZAMVdVsLVi4bTXVbrh8+mrpuRT/Imomsd+54A4Rccg8/p+NwSqQIlhStvo9A1J
LE5AXwD3Wx9a2xjoQofD3RCNx7SAWjQQ0TAUyA0z58ydLKwoYTy4XcxLyMkN0eoa7w1lc6aXrkxr
ahPVU0LT9FdMQkFJe7YMl/yVw7eXO7YuNa7btWCWK1H+ZyGCkmkgE97jbwwmOxJxdUrhfTy0zlrh
QcdYrdczj7L8w8BotmQAopPE5AzR7qwkuHBbzuap9ZMuyMX4ATrJqrM4xQBJwzqbzdFKCfFAO6IY
nx55hsl3YE0vsD7dKKSVjuEtROfptnLde2bvKeCqTtn3jkMYbNhlfB5zonsDj4gJim6VPMNpg883
LXHH8b/Vdls+Y6eHql3/JZd8V3IUTMsQenLcp6eRcJB1sDcRyosWF+XP/zq9bFcAT2GRDHpcUr7m
hB+iYT+RsoBj+LpV0u6tnhCGwt8/syoEy1GkIXELaE1eIlA84fX/O3PLFMecgTSRBjtvwLq68VPJ
uIA+2E7C9ECRK0sJLQ0+5wnRd5mb8ks0VwBreFGDUhusQHv3cVbMP3SSl9kOl6vhV3K2pRS2GyBy
A2SJl5p9XquADyH+n4DF+qEE+H5oKs+MYZ3NLomvlzDgsjQQnWD14vB+L5oCQf0C1xm8Ffpjy9j+
G1edeoqy8+PCk5LldDpwW3YRx5RJXbJwoKVHFE+1exN4R1Msp6lHFZF9VMLzwclhdZEkOmiiZPdw
448tNXahPsOVwvR+qDPxGYLXkS6I3d0LxGCkr6/Iy+9T7dpAinx2q8fB3rcDuEQajekQyhVEj9tY
D1mJqyH8e4wNKlPru68RrT+Jiqb9+zfsF2Nkr8JM5MS89H6fALiRemV+92snsY/ocCzkmPWj/9mP
3QT33Qb/zuVnsjAc5tmPqWMo1zn7wnzNGUISnLwDSSOpllU2GivsXsCDDcnPipVLRQ4ZNkhcBN6F
VNf+f4JbMhx50anPWIq2Fe8UcwUFSPYv+FwiWvT8vFJIY3/XZGkAaKwLzZvVHwfnWzp4CM1c/2WO
hGXbmIQDyQggyJVzSAe7ctJsOCt9QfphTSf7BzewYFTASUEH+tLK/qS18JRgzI4xesc2Ew94Ht5D
m/2yC/YV3G0MBPscafuHOXh/Su20DyiuaQx3AIFtJBC1NEa7qoH/3ZS5fbmvpBGrX63A5DO/xjXm
WAxOz+tJFOOFIZne5r6O8lr45hILV9mQ9wf4m9S7p/5cqiG6aRbfMnJBW/wCcdKwJatxK1iudxQ8
R57qidK3JgD1+L79Ynq4FQe7F7LLN7JfGSEXE3m7abbXDMvXI/3bvkxGDEf8FxJmj2mmtX7Qz3vi
p4PxWAug0xBfjXi5HobL+UZwx8f4xYHhOd/jj1fZDX9o7s9axZVZ1xRSGMFwEotK2XH7sPnKfdzf
5Zu2TBQIJGw0FFMw+2iyPn/2tOFS/NBvvy1u7I56BlafqAPUkNC2PmjHHz57ID6yWa0O9yvQzT9n
zcaQb4WOTD+Ad/XZaQd1mVtZCr6tOHdYBsJle/7JqRDTADNpy8YRaOt6aOMXbEdEwVLJ9FjWDCKP
9lnZuck3IIm8hfgT31uTTsNPMbmUq2jJxHk1eOGCOdoxG0A4vOpEJxfn9b5aZUL0Qw20shFsb7VQ
e4UIPF0+3vRprXRaUXjKYuh211lxDRDuneV2afD34eTUTEA60oqD+lfvtEXWOBoE17L0vkttCIQY
UtaWp6gfHzbNm/b40eu2mw2GBxuZn6ubpOioDHSYu9X0hDq8rjdqcXxU79Pi3H7CZCug9/aHDi+m
WqYMq960o4VghVEFZAxFYIVCJZ49BaXfxDCkXMZRbu+/ouow7qkp2hovbUhNHeaK5YiLDzvAQIDp
R50Oqb6YxnM9FG49NdXDc2jych5MCT+wJ2xl+7juSj21hLsX8gE1ukV7WIPtABNea/6sif2EnqG4
azONmcBFKzsQyPuYwBoSyViRE/akeV+Wbwrr4n5UUp74zb25G2+9KiBNwoodCLESIgtTVQLfMaQV
gIdWv8uFve+L6SHVxkF1NqdsPSjEGtH4Z9e6j/WAvGa2r6qgnkZeT5rsk8b6Ui8TMKXNM5Boy3T2
gKBYy+euF6QVGfOP1YGMV6lJAxC5cNiIkvmaxYXFblAZdjETxYJbFJJPpLTh8Gb6c/WPQu+7XlTJ
Jkf4/IvFylH3CIPS5Q5qwwr0MdN6pYZ7gknaAwKg/tFDFsgcIZcK2wSKGdHq1NCBPzi0BYH8hbw6
qce6ZxJHFiyFXuNmEq+IiY93jdRH61W61ZTwxvJOTHwc0w4ZED88Ej1TIFDJE3dESbZEX348rg9+
1FNTRcZaDvHkHPn4uBCiITg0OtrAbqVFeMXDnUUlub2izDm+YYkwAnk5c7MYfzAdHEGGch6FZiwc
0TRYmRQqiT1UoR7gn+emnP5ZN8oup5zHDjmCaMkL6hAKFImIM4Qzl0Xwg7xh7lv0XY7Kz+UNj7Zq
u742LAOWNlI4KGYWz06XRSEuT609U4O+D/c+VUXo06rcvkC1EQb1/WGW6aYKzAta3fCDpTa+olHj
Ri76NOfjkEKOlReLtmx4B0pQTOvov6AY/eoIGNPsK5ALCopPmn+knSLED92iK1sLuO8bRGYvZMe9
fJguo88HSwh49evvJ9GLSge8tNHh3CNaF+i26Ig0XDsqTwgO/0afZc1wDFJtWT0qcpPn5qKm9XS9
KW/67aArxyjjZRS35QsfORLEALDZhdWs6z/79YZ2Vynu5N4VMrwzyLJWNc90WJbb2QH9akB5eGmx
y2k2t4Qxi4lyNEB2wtPgEy2Rw/X6gSVhW5BSonNw1LodR1LsREGvyXP+e4io31HCxOiWdXjnENnZ
YCNPkQ2CMmpds3TEHZXQ25n4ZBFdR0MyvFIA27PJTTQXIiTZkO6vHyYd7pVLTeL6pn3YFEw5LJ9J
dbupNCch8W9V+Yd0GozvYjoM0MeBUPNzeVsbgpphTSyOapY+hsDKpKlAd5isbZlaZsxjOPu5Lykw
R8nOuSQ/Ujljq/2H7ePiuCYRdJhXnIVmw9IRAsQKC4kAt2tfuOdlNY6DXBmxLhLMxVTYjQ7t8xyh
KBwalfrLzizf3VsUJ8+z1fb1RnmXkIys0cfeK+Ob6KMF7PTaR4hdNa/PLg4FKrmNt+uAl6or+eGI
MkTZW+2gLRoc+wthPtfHotvHEom830l4xNzX7uvKHyFukCeRNSJMnEo8ZJ+yStbd6e8Yxh6JVJ4H
qlSuWWt1pdrGZGQF0R8P7j3dNHv318kO5PdrJZhWBDLTL3ZDoP4e3PhNfDKHwncTmiERLCPN2ScA
evCwDCmOd6yf+hQcbnAxCVb0kZZfWtCcgXFv9g3+YX6mObrZi+9Fm+CA3zupmuFp3RTEjkXwHNRv
6dROVNSr4zpD3jy/cKMVidZabTFj5U7ZCOXgvCVfmwaKG9HSnbBH5UYutCAONk45coPNcPPMKG5m
YEF2BeYZTew7XTpEX/lzg+SpyLL3z+WX5DuCUNbRGtD+14TEVymkm6aI9XZeITkHB67LvqgsiZH0
+puAy3QNE5Eye5jyHzIC3IkLzyDb95MtBgnV7pCQzC6RuDwT6W7/UgXKKGku8xmy3CW2BjYHxxgC
IbLubNHJsuHPUFzsaTgpkKYOd4ffHF+wPtwbEDVzVBf9yGFYeyrv+0e5eFIAAwwzp3L8pzr+0eSX
aWaC4uJHJHxIJ3NPauCHO5RlSGFMXVkIuuT/BG+hNQ6XIND4dh52bhn3vkKT/AutgV/wrFXjF7R5
IBkTAS94DUS2eWN78KE5prAb9uQZ8g16nzlodCqwQR3pj/FpiPH7IFu5LCX/UE5mgl59w+Ws1l4I
p/lZZoq+Y3qN6bjmvfyBiT+EoqtviQ1ikQE7+1TAP28Yb4KQTQ0BL5QLmtTNVK5/XOHknrUb4Ub1
JOKyNNJhzIt3LLK4wZj9UGR4xr+XOjf2BAw5dSLTa2vawSqZN6DjScIh91MHekomrGaK98sNmta1
zn73p1d0Hlvd7W+0j7FJPN3N4wX3IAzkIpvWJskoTa9AtLUD/MBc5czpQs8owQ/NI8X9bqAkYnWh
s8IWCOIcY9b+jUcd7brMOPT4Vhdm+/4jlKmHBa4oi8a/SD8fSiUd8hUjziUjQYXtBP4fGCvQlnXT
JX/ZmSPqXyyHjE3+lnicC2ZY/dOzQ/oorwNnbRlPjiljdTlsVV3RjJoJvmBXr2wyaCGps3DVnhx1
loR1zVQhptW8Si0FsUSjLm9WDAWqfyw53Wl5qKJfd6pGmnJ3oMZmuNU/iKrwnHmE9f0eVWQBMoAU
kgVkyeSLLhGlZeZ5QzXwvuG0bjPdbsCgEWdfaC8sXRIzK+/6vIn2+RJmy2fu8Z1y2pM4q3wcGoLd
NSgfx9K2Ts66g0xJTDsKxK1xIOhiJjGYKo86rfGQDTrO/0tmTGC669m0OwctF+h32+9GuhPFsyG1
CXyP7HEflhc74UpADjG9wQOSbqr6VUEBrTYS2RHYLiibibGvDfroHWtPvIGtnc/lut289lXjAFsu
tdS8eeP2wxF2Fekxm2qGLBhROnMH7JFOe6kpigEF8kAtPCtx1aAXXJQ5KU7KI/+EM6K5SsdaSgUG
BGRXzF53tS3nYXAjIVq7/ARNL3YMDv57mMcfh84zKDrxRJlMII2usAsuLopfFc9UWvE6lyDlikWw
lxJ5iQTETRZCuvUpggxjE5N838PtIcZWqMBHAFzEt9m8wVRtoE8UFv0ouB2oia98I5xjmNh9LDMz
kFamavRnat3AF6inrhDRAb79QTjYRYjPGF+zLIFICRCtBHULHE/PO8PycMmn7FRW6fMCMuRsuFRz
3K6giIvEScQok/xB/25jl72plc62L0wzPPaOSfPT8YF2WAlg7dELQ/Z8Cxxq4zzLZjgEpF1Z/Hgc
lJxZ6VAhnrPZVJGM82G5MyGRnQGhRiFmM15SGxCc6JVPewil6DDcTBf38w0QEl2P5TJCByozrPJB
g+NG1+8ep2Xsm/pEVjV6fxzjTY1BfJgTmEbnrGLQ8jfW1HY0XM8uo36OP5OKy/IUNruG/QXeaMgn
Q/7RKXWIzZEkht2lTGNPGeQsDAzV97mmYOX6QcuSgTPccK6IBU5rVKMxhpRZLT16biQdKZhwb1XF
vqR2e6WNk2E+gaNcCJxvIru/JVIirR9b0tfqTzFcZ//qgpaZeagt5pWeQ/cDzM/2BJ7FBj584q92
WtNOurqIt5yi+jDWC9zqMghWoMMEnL+fDXl6NRpTSlvf/xebmT2Q9joy0mE8KCYIDG/aBbwqcpnr
qcy8tJKRfUUMlGR93Ef8BAlyHskmQERqoX/t9uYUaAjORZtkvwVz1B9ox0J2D8DItjxffN8Na6um
wCzDGgozvEHDoj6A7vp/CblNZYw4mKjGlZVQd57XA/4E/GId16SoEJlxb0gDcudt4/rg2oVWlhU3
gUgetPqe05MVus1Y7HBsWO27BCX9gRWWrQf+tv9P+3wZRn7Ej43h9XOZltQ+KSv6aBwOIitkFCXo
BXmjiycF1aC6wDjfHDz6CG/F6/+GE0QiMsgzw04Djoz6PQKnukfUy+Rnoa/aIigf67j6fm3TrG6v
comUrDRS9mx8o3zXQ0OWsvC0ghfXonTvAafeDJ4BG9F1bLsc3KL3pobkVmhMRIN4eMvf8TAI3xmy
MiQM8XtpCzTOAFnBzxb/8BwIoH6Wo4cJIkFt0ZXd60iFjNNELQwzIRRjs1j4v3BVJJRUbRTmhcFR
922pzRse70O7DtZTXKFEYAm32TXorDjHyH3xiblToojQQ2mN/XixAdsViV0oSAOr2y/Vhbrl3hH2
ujGM/3lphWdr15xlJd8uUixZSnKG3UxCDWdaf9nGq1HTi30FWtp+EIzh+7lD8/WIc0t5AMBMWtyU
a4B1lu7aUYWLWDW/acacHPUAPZYq2i27qlxHSbhuZ4pNUjAYp6HZcxzH+h0zho8WKq4V8hucNndW
LyoWX8CBS9kWE+DLGxxP9fbnwAOaexq/doeGLQfAyhS3Vfc0XmZmIVHf7AWyniU7nJJDXScDsfRB
ZWRR90UqIsoYvH4Bru8uL6K2Su1N+JGW9wqYhW+ft1GNudZ4HaZCHH3CHU20tr6VeVdKPuz7xACu
NOiwGssvNXsXPpuEtjzNgf9kz2cuF/31EBNgDkF9ihHYsIxAnSvA0AePEs1CquiVvS/G7r3ZICEt
iIc7ypVAKk24UoCgsZKDz3JLMQjFTobYQ/Idt/hDz/xRxfflR35q8LHjuNuTzOzs2kizRSCvx5Lq
50Pqowe6+tBGoUSSXEvqD9h+aNRU1gts692HwnyUAM7wndmlohkcGYzrh7L9w1z0JRrqv8K5ACkm
oIOHwC09saLYhH8V6J8yxda5zbyDFejhKkSGAu/3SR3xUe9AFEGGrlMqitvudtdfj56dMLRh4H6a
SMIl1wQ8yExjs6CZICuKCeGDJJ4HwN2zHQj299ye6lsgArc8fKSLEtyGEednXSBaO3nXc0Z9kRom
uJohsQjLKmBNIwW3YMs4ExCSwub6pZ/+tFYQDXWfsdlI1eDp2x1r09lq7DwxY5/KNFKOil7eNA/7
BGPcCwkIlX4igEwwhQy0cPZgnm+jv0FJQ65FDeodyWr0CHSRg1RWnA57/bYa+gqZafr36i4INmBT
GWOkyr7pUKy0BFzdBGMSx1jUt1rnQXPaC0L2ZVBjuEPxRYgUHKNVVdFRdrqkfMvL5Gp8rughxANr
NmjHfoIlWLXp3pUnMylJ02792pepeOOuif49rfAJKl328+GTVXkOzrNYppabM6b2enfCvVunMJi9
xETTDzJtg+qEYWXABXd80S7VpmWt4LZ0PMsm1CXblX7nGCETeFcRoLqRk2/ZJkKpOMFQO+kT6Bi4
CVfakK686y3AyOnsm0oYyrIcSnuaAQP5L6mcIZUC6MoP4A6SE3kiCO30NwOudHnijofRxTF7rpdm
lCDvt2msZsnpvhWZz7JymllWqu1cR0VICx1WAPTVAMCJUJlyGtYZePaFq2nj05NilIYXF/VZCy8b
ZpH4/N7dyt/G7EPG2g9vj/McaD6NMyWQQpS2ypUek4ohaVm9yO6IM1wJN9yDESyukeYK6BTPzO1J
CpDLUGimBKiG0IcvPpzbW02sZfSDRXgkpP2JYuCc2wVIFdMv7BhRicW96dyKDBt4cA8pqKEn1PxU
9CAx5nPff52oGhV87WiGK7U6i/P5nAjJNS7t9saekK75yMUKmq07OOPvqrMs5MkIo00s9QOsOCIM
neBp+m0qxqns+pKr/JZdDd+6fktW7gOM275sQbIODScGss58NbCqzVEHhSZaFRwbIP06SwnTH0qt
GtNeqea2BX9UkDhKZZOx8PByOQ7MCFFG62D2/oISKWWN2P0795q/8KHcIy2ZiR0sTQl5uHpVnzzM
VJa1Cw5mOlDiG6SehqU7fVKJaAHJYDRaHQt3krD+9DhrTom4/nm4h3UiAwlsViHmHethySmu6Ugu
NDRlcl8TrVzcZaUGI3lsN7iVV81Y3X1A5Yl7+MU2Y+1QK2QG6xfBLpz+qz46QkkA+INGAAmyGYRi
nEgXCyiXxcl5BR9SF29VLI8xJ/AHxhhG9fZqFuqA4x0w/gnOLgT8SH3RU8wKL7Hp7KM7vi3326Z6
frlPg81t3grueYSZ7fwJBUM7Ezq1DqFYRScm3FxvMmTyU/IQbjkQdS/ajweNvzzkjV43YhC8XaBK
2Pad04rXY+3fillEucaAwoP6Y6RvEbseKW0DhOY0pNNDh8EQIScvY+zBkA/LO9ry3vE/nTDxbRTR
qS7xp+6WblAlmvjbWFeihZ0BsOJb5d6q22PO/lKhJ+eq2OlZwxQvM/k4FnNJfTzcHlurY21rI+CU
lwJxP/tP2PGqzeMjJEJ1rHDMomeVY+/C4JnEFhImel8dD//ynJyMq6oPZ0u5/4u3fgbH0yV5uXfy
RTl+XRnFHfTibbqisX2I7qa8x23k6AeCnzhwdZszTh27OWrAzKeb2HSRDMckmgZthFUYw65UQVcT
oxPUVsO/CPYfl+r8fqBiKFa0qEAOopz5YX+GfZLaq5Bl2otvekm8VJZwnPTNAuTqoBgKY8xxA64r
Cd0uTjcqRttkX7l/2P/mlaGo0oagngQSTge3BCjMHPfczhp4uj6Z2jlEecTwOCcN2gX+SNKwlqws
Ysq8EJa05AAoA9saU24hJe7aW7K+6qGLiKnx+/7V0D2jJD/k/4S0+D633FW3WIGVcv9gQF6OZVVk
gmG2oyf7/kQbR1opBtxq15sDXU4QW/RFKvUaLfvfZEz9i6vGbqPN20+peXBVpKoR8eP7GbL/HHsE
5uYk2Wb5mSYi3a0sdnc/fEMy+Ycbtx+vnw2fisRiiQFPb0ggFE3T8miv321vGPqITy55LZ4SjIFS
4fWGX8ckhP8xVp3+bOyRVoV2V4eXeCL7gUYAX7u5xLhR6V/iHPJBDy/hUa/1ZpqLbs+uyQfR7UuF
wC/UEaXQf4rFvdYB8Ki0m1D11PfLy7npJIAQmNLUI69C17O9dj9QSDfkYDJOU20QKdcjyuQNjD96
nTtNdDzjUnSsV3HcG7RJIZI52e2Q60D0UNaEXSeStpXc8EO2S91Dw13hvJgNONBmYIlvsj2yi7zn
XBMMqRAwMrJZXgPAAfMjA4WM9558XQqQI4KKYie8qkIo8UyW62z8Vy9Gk6Zx3vy2FPqvmB4j7dSn
IrAfMmGEDNeQYpQmljfeaPw7SGyec3TTWlSN6FYnzhuD08e68NVWcbiw/Z5DiR52zUvzAUFpk+TX
EP/Pg6WoJhbhhSIxPkQpS41Vjog2bKk1tEgdXRf/awFA32n0uEO0ZYJYjM/qRJ8gHRCRXheio3fY
DbpO9wEKR7FS3Hm3KVWqgEDwku4JLPOq/WfJ88b+2STloNIoBnPa9+xXLGmI67dvdgt0ppm+yAuv
NE7yKYlI1IAU53pLk9qChpNz51w48ldAvXy93G5dvmu6IQkg9kgDZvtovO/W0U9YII2YGHy92pqh
r1RPFwrYm/0VT1v6Bq6KVsvfLBNVdhCnbuOdNNzZtUe2xy9eIFjgIW0orlJEHcOT3gkF0rk0TVW9
0k5gk0n0ig460LlkXRpOebLCq+HDxyIbZiQYHY5XGxa0CQagAAI7SiPEB156O57uUq4l+FaOAt50
Hh/CptjuDfZz679yhBlPsVliJz1Bhu2rhQeJdosjvXYLsJPpIT+ZklqzxpY8EJNLtKBuRjIbDqwa
+I5mNSUMRujgV1yPANDjTBfygUkF9h3cONnRnU8FyzZRcrly7V7PIjrqRJaqVPCnuwRI/MeRpynl
cnsI4+xVNh7pRf0oIOabWMs/PFpQ94ZGp+byXLsCZ8o4iTPPxaXs0WhGyObQ2oCjc7cOYObXyAss
ABknG1Mijt69/oNiDIgPihcWtIansuIyIYUxEBGjjB6cxuZL97x8ioJVOls0vI/T+RvL+9FjFTp/
Myc7q1EFcR8n4komftO2/5Hd1iF0kgj73gOSCKn0MMWl54+n2QsqwQ7xVwetSZx8WZ1zlN1KbILo
FRQLHmPzXEBI0LEjVDijiWZ2WzC00nbrC223uOLA4Mcy5e2RlCMYilNy7AbS8nKxAmYJwbfV1fCW
TCZIT3sqg1V9Gcxjm5r1vUn6vUaIf6zDqpUJOZodC/AI5G0s8w5ULVxDvd/yQ08rHxDp56rSQphW
IIOWKr1jHjowVVYltSdAc+QJLba1bfwFWhmsiCqSHCySGtxiAPHqMlpBN3gkhGfA7/tRJYi3J7Wl
lj+yhviWsik2u06/c0IlcwCd2Gw7lMuqkcniONNoWu0sgqUEfToWPSjNIALO3g4QQQ9SJMV8UJGY
oAtkI/hSjD9VUmGRtiuDccCCJSpyWbBmIbI0xcHMEoaaemipBZV63zRB5NB/buS6dxMGKgStI2LX
kFofJI9TccAiJe91VP4/FRPoG0n/PuowoaBSU0Noxb8giL9BYOqeMGUBlhI9hTBhLXPYjMfI8u+m
trpRy6XhaDZzRdQgl8Xpkkrvj2y7SIwTDgNr4PDswEyo5ZYagM+0H5sQC/BA9VCqVvwwK1pJaMhA
ZHUXFr7DZOqHtXwzarkEZeWtck1u7RixwLD9MyBgsCopgKx4kvdhIN5bV2v9lIkF4ScfP3fYpTgi
btXZqwtUxZ2F6UxXBA9XDMwmikSZ+cLXN53YITp2pwXUmylPks7v1paLA1hITRJ1OF+8EkHvbzBC
vf9D95P/2AkEUop7nAvpV2eBmtNmnzemzzulN7OTbCWW1CmpSxv3DVHF2llspdGikmrkDRdKlzhO
N0+c5kLk5ylQDfBXwf6XPY+ECgTCrHtDKKpO6ufAtHfgR/IbYRUVwTdoaiwiEcBEo8lYX0KQmrwY
bTq31FRc5d/WxglV9cGXwYqYXAHbEkUZYx1+oD4plChb4BhxdUmtDlwT9BKQoUm/20SAnTdaSPsd
aYIbSYjASjjOfkmhxisoxih2CC6Vi0K+oohFhAevr80dZO94QiK4z6YMEuR7DB3Ho3nDv5T9MhG3
oL06uOityvQhXdreX1Vtc0ik9F0Ci0flzNX81yzlg3QApeycsTkTZKk6urEiq2EpX4nzAIIiXcC3
opKsOrzG7MKOaSYiTo3bUbyqAGBKRYbiij6EemrDXrgQ6q8zh5k1cKQ50hdRecVa7lXyRdlbe6Zt
9q3njKTQodOP2Bmpd6mUnzfvlegiB/LdYfkhn5l7bnlRam5zx47a2+wsxTEyWGuZ6m6Ep4LAMZ+1
8/xNQHjwSdqftsowT7kkC8QQv/JOGNUyflSjgxd1HXUNJM+yvexw2qGJHvvj7ckXRoV58849Dzm1
1i4t8Iqk98yfCeVuN06dn5ulvnF63gZhiNSdO86VyHuHUM4Ep75v76EsU7gb6Ke/BQa+RCiPjfDi
j5P/OnkQxvFFbavQxXi36XJqgaEpJJBi6HdjCwR3Fqk3un6ZA6yYNm2O10N4ZkSF5WXyPgTiTL6C
hzxI94FX88NhjficRczJtD9wgShUpz7U3wJ7K05kaSZqc8ZDvKG8wKnnSJAM9UQIFTVDArvikuJ3
YH11ZXQMNvufKARddNXxCaFtSP5CONTCd8ppiiZczj/bNemXQXj3pZZ5J5AIOoUmgCtqn6KfuYxk
UVp1YEv7sbok91Jq8p7chSHLP8Nmue/ApOgZ0zXyf36MICJ8NBt1ooIAVJs5OZwopmhX/8IixHqI
WXI4T2WodjqZYS5zGB/AsLULUza3tURymQkBpdptVvB9NngcvozQFlnd7hX7mHDmky9hczkF3CnD
Zu22YUVBBGMuRiei17sPJgqww3pbP9v9x1Bdf3v2/QuqQmAWNUL2s+NydTDhR8wHsHAn8x1uhe6r
qT7MOX6G/jqGID4V+6fdQ2raE3uQzi9llppK12FgC7Gv6A3+eQkI75D40L9lbHoIvHhhHLSpewQQ
ZPm3vIcULoz/cAne5ObCkog2XMCHm+LXd7Aoom1gMMfqBI+DFKjFhJQv09zR04a4Fx0n5EL635TH
cHOSlpiwrwsZSlfJ5IWM0EZ7aPlx4x2wfRbBzc4YTzN6QdPvRCbjXvF85xNd4RJlNJYFBO6O8UM5
zgWLT3IWm8ezm4ZavpKJvIRtnE9NccnUEBVs1h3wUwwPZiVUTuIESm543ncaNB29w9W6nFp+sWel
zrf7kEsh8RFN6UWwg1vhpzwNi/OhKIL/dpTDKEg44uDTc5aDYpn//DpPXIuNDL353WjNH8GZ+N7O
ONkLb0HlYoHkqMLc3rMTQUI3lu20i+pikLoXVY2fqJeiG06C7kx88LuiUl09rPVHrLgvodE4ckEG
Zk4UIHPewxw/+RPff/6D5M5oUWJNW72FdVua45mqJFY5R0MI4U5eyruE53epd4oOGflnoYJROWxm
2LipCEUeY2oGT/5706bJYnBz648NQFE6T47lyEWzt0k+0tXQSJWZT/3fcHKl0TvHS2sYr+ru9xED
W5/ntONjGCKmoy9fkeOVBT/tNBX6vK75yzRBqkhnIa5szCMdarolywIwkDGgF4gUQiGIyB4qyaZZ
Uu/8taaw04SQsB5xGBTwoErL+ZF0We3FQrPLKr9pu4ZnDejXew++E2HecqWsMf3iD2z1iT9qqjiv
v0GAfSUmwacfISQvam6hiHVFvEzQ/K7k4meG6YTGlAavrOBO9EidP1F4oHDDgLjintplJE+qxs5+
MTsK1C1x80Ye6ncEdOM=
`pragma protect end_protected
