// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tmLJevIYnLannLMnEydbc32E2erAjNAAG40wJD28es6RiU4SXtYaZwG9iskHabJL
Mxqx2CQlFmqBAaNNtsFJgkQJmEOIpTmzsn1/wg0GD2Tn5RzrtzkRV1lXV5V+XqWm
Zap5UqZWoYO45sCZCrnUKrPrGlAmON7c1DRqbXah3pM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9424)
d6caG50nz6LEpXIKUZlrpMrxslB5xNsFrtcnXMJfj6p59/gL1bV2+MT0YcKJzERL
NTlF2FXFTdeWZS9Vh1XeBmsFleCKpF0wktXrJJQCxUEIUFXzMsgDIiiKegklmbib
idD9iAPrAIv5cdd4kEuFrCGqQo6ZwkQKT/R2DFw34W2nmtbUmAYtQo57jGJ/8vob
0pdLj+D0fONy+PH3LMUI+B4Ix1iYriuiaZqkLrQ+4e7HYTnZYDs4LN4ohgeVq6Vw
CuS0XU56qsEMuwrm8Vi9WaXqjcK5h6/RqbvH9d2ymHcXMn2JWnJQQBLxGq0p6p/r
3yONpTmTPQk+xRTU/A45d/sjt8Fj/Scip90Fg4LLJ2Ng81qQnYNVWQEj8ItgsuqH
4FfjgVLCHg8ydDCVO3RPR2C0a4n5Xu05FRsj2nXLaPe4NcZ860zUJZA3H5fKgdWq
2pZUvohqcnmSd+X6Jq7UZAEz6lj/qde7mD3QC+C9wylsglezZVUy4sJUiiLyuXUB
b+qX2nniTzNa1d9sczdyWroE0lbnnOgyxFxSK57xNVV+aoVsaEPEVq41WXJBcfxn
v+D9WflJj06kHPbrYwVsdvpoa8MLGt5hNfDpNuuY2IN1KR2eaV18vMj7Z2GikfK7
c0YQxkbZ+F9t/NVHHkjxUGiAIiFTAysPM+pW4IgXzmxHDC7n0RzEYBpIW7jAVSye
OsrtORogNDFg65zfcBY+xHMu8qZSUT8WcCJyfuKjr3TF7hCX8Up4Y5XQ7ao5K8ei
DF6jIgGAnDL6EljzPwfauKx2YJ31Y2M3cZplAT95PnQWu3LQ5X98RaZXsDbtifi4
QR9VJ8D6PqDMvT0Pj47qW61zgelJxIfPfZJgHSHPnXrCeR6+CgjXAj/RyL/itKrS
WHf/Tz/gwZub8/O4W6FCJWebJPnPLAtKUcaSdjyxKnzACce6zpcoYr6Bmu+GUu2H
T4Fc9fmOFES5LjTDc2MfKP6o/13H+rLtS07UzPcwmGLUqHfWij94cSJTUlC6yoNY
n8PldvK4Fp+LvGigVKV5+3MSevJHd4Z975aCjKqJ7Vf+gtBicK+p8a4XUK2RGZyT
6zt5XD2ibrTzeTTdqfteDmwiUdE2ob+22MWRLXxos9VPSx6kFmCJ3umuqztLXc8x
EXQ6YPbsHJLeg8JlkJQsyuDvD5KFXlaT6fOayV1ydM1tSZowDJbKTl42mHIZXm8O
P4qC/q8LXJu5+eV9OMRklpnhi+/dP6xw9f2fy8qLUK0WUy97Zpl3CSD4P9ofZskf
YDxCsrSbWxqrgelqtAUNujQuyfErVo3M6t2xwUAlfXldYPZFG6TfEH49K7yyHO/F
8y70vUJmk/1uXEne/YWAGHXMyfwrH5IjUWj64fuXXFSrRxF/79sri2E30wW/1lvl
WOldTjDg65rDuw5YhEDCMbcSMSNeQQIsAW6IdpbTMtibWBdQI5/r3u4W6mULJXhn
ZBGTtsgRbAfrkhCm2F9/79/FXDd3v7uMHjoDGf4u9jtDjBsddxl6rlECANRgO1Hd
Zpblpo9SXRnwRtiyAjYSBCCF9KmMo8d8xb18I67FHTdYyHtPseGV1uUxNBaD9xoF
E1LWVm1rAhJI7VJp2KL3jFjJiauiWtRhNuI1LlTuGRn+nFJTSYS5v6pZ54Rt4bH5
FnPU5kB+DPCXfE8PzORWg2FYd0x6NXM66Gj1bjvlILe4JRk639damD7MqScjx3zc
XegdLSEoHDj45PtqUP6Wzn+tPFH/0pse7iKGK8N20gOhpdRnVIPi1n7eC2krxXRp
wy6uI1Y5IgMnKSlL1WSbqht+IrLvijJaHbge8h5OwXXxeLaz19PY2ruqGLTQiPHv
zf277iTyQbV1mjWV100XIS/eHujf+3MUIxw1tGTIkmLUh6v62pJaYyj9a7Mw1eji
k2uMCXlgtbi3A0RLvIZfmjy45J+g84C163VLqid8HUjARhha4Cd0JVlXx61cuF2o
K03uiZ5a50J28nLXXAVKLYpVV5S1vavvVslCdfC4SmkxC06l3vhMcQMVrFReAKpn
P/Dl8pOMS1IvWfneZBBe9AYAOQVquv2qOYd1yQj7+4NMq+xH7ADcRyp9Nlv4W3E4
2QHvck5+JoDiSb2cz/vcL+iHjsvNwiutsybh3PaViXJNNBlUh9WArFiuzEiIQQBS
uB+wrdpeeM6jnqcJodvdrLYlRh6sT86ZBdnYfMM9naLJ5qhu4jfGJPpJ5QGwlVVN
O1Dg+kz+XsndrV3aCXbGFzDQxle/2xPOU1F9mXOQWJFKJD09CuAtJ8mFqRy7wnq3
Ibd9DwyAHC67R6JZgVPn9SAVJghRIw0nlm1hJ35y+p/+Hgt35aYomgYHvIztrZ5N
SF1yg7Lo97OSl7VEqsEGTwLUMCrsoZBkglyQvkNmKYjiKUNjV7HbhVeGU87zNa22
ZfEg8p9cIEt2ah4APQPtlR/O7pWh0Z6acrgePmWd/ntiamrGfnS3iwf3GRnzsigJ
+nGd3SyflQpr+vTgoRBRZe/5RDhuIGctuZlrRWO4XZ3LARsW/OqLlh/0TzyiS+1t
uhv/VKrgVU3Jg7YnNKv9NGnPjTzJC9yqlHtObD27+UMtjvUUK/qKP1l/d+dZSWgs
y8lmm4X8bUAjYbQ8VeCbk6dN884GQeB0pBQXK+Nh1upHAJ+aOAUwaN0uPbWU9ILE
kYJ3564Fbzk9YZSX6uqt68P6HbbnonG9jXrQdXfVlqxljHgaCEFf4I2mWS/Jz0EK
/5HmO7tRyiUh3h0IC9d4tmOiuYGrvultumWmq8gFfytVFonhJWKMHoDsyPkJIycM
qYLSWGTP951Ceo3VbJTzMJepiu4mmzJsuWUXFWdh7qHoY1NMkQK8Hb9tIQXj+auh
IQuTFsSbCVSfsZx3frzqr/GhbM3NFDLPHoqlpcyBm+mpdbUbrO68t6tKvD0eZL2Q
PWQZ1L4waIIhdQ0SYNyJTJjQ2AcX9IzH2/AUhTsbwBhqmFudL24Zt8VoiY/FTgTs
+LXN5+Qh+pHim0BdRNr1JCcjdcdCB10MmYWlrpnM7XiU4DPf9nwYt/D/9F915Ey2
rV+DXJMuUXB5u19JoewfrlryqiBOSiXNEngquGKLp0pvLeNhnYEvQtgsUiex46Yc
nRWysaGGFUc028WTOthONOVqbYaPlth9EtXE1P0N7RynJoy5Q4xK48bB3LzQ2sjN
NrhjxzZFL8rdP/O7AyRV5Fbh/sIjk+qtaeniwsWFwRDTDyZx41N9t0y0aMY9z+Sa
T3NGkW0BGXiQn6TV4ZDqjrsti7JeuSACD/Gsge38JMZpxdmnXaSxr4HiN7RqyJYJ
ZQlBjlUpCSxVaD/GKt+kgtiO2mIvTtnEl0ZWIj7sKu1EK1gXg/cMhWwgic/SsI7Q
tJFKmnCQQ2VIF0voM2ZHLxH3e4av4+ie0gLfP+qwZUMLatQJ1mT1hywyJVJjyhfD
/m20PouFvAT2Q9Edzc2e8D0WE/n4uprWn4gRQARkoJP/wz+RjSAD34Rcmv4uKYfv
iKAqFOCrqEyEroFAxZTnr3SmfQxr4QV9P35swSq4F+tgAokNwys6ZIWTkl58CowD
JVMRgbAwcHHC6s5bjTeN5IRn5C3znNnxoXlth5mEgn1JEV5r+TOcHF12963xaw6P
c3z5w4Om5PIob/o/M+Zaf6T9QaaN15S37gKOAmCK5b9wcOySHkVsafPik/22VUS6
P4qbgx74aSuqlRyPVEctbQKFitzNAbMyn+Y+9TIv2VPOwjc9iRMpmvBcyg/7PBho
BY1rDpvpaJrF6AR5x1KVreA7JGDOOh/yO9OXmy4SrmJx7NCIkHMV/FHH3g6y+s4j
5XeFQpKTo8bYjh2I+E+HN6lpc7U0+mKDb+IJf3WOzc5EdniXrQfuQDROhA9kOEq9
0lS6ACM/WieMYPk1G/CmTVVuJAXTFEK1dxQr5ZxhwQcF1rlGWi2QZrBrOmcj+WBD
iuOo2iFfkwgXqex6fXL+vgy+MMYvb5jCbAlD+z6v0lUKfZJXeOXCki9KjM7oc4+Q
juHzfxAr2GdTVjbp9mdc6B1JVP4/tqff6Yi/tGjAm6orcDGnKFTOlnenSN2vf6mY
LtcU1rb147s3x0NqcKhXeHD6xjsRNVJAe2q+nXo5kV8EI/9P+6dxxUMfniv38kQR
1sgEurp9KZoUXE/k7iuvIK6jhgn36PsoYip+3d+EC9psLiws617tudk7kcA+30Ws
NBvwMADqgvIQlkKNKEWAuji2M4XAdNEO5e+EnhKyoXiPU2BqpdwVfQqp4kNSYqgN
FFwASSV7cZRJSPXia8yLW24VDAOFqid2mRUUs13ML4uJcvbjjYnc7+6ZULC0fO7n
7GOiwAemx3mb1/1Lxl2S5yLpQ7Gg1Sxg/xNTGk3RRdQd2fit6IOcu5DLomBcm/sU
1j1wVLfnF6EEd8imayex85sGy89idcZZZQhPHCcp/qWmgwiCb8RUbUGOGz+ojYmT
5WpfaQU3U2ZRQLbUnBfveK+e9RgelqUNgkCPJFDObnLzdLfrE3bX0fHxI9b2+VdW
mgi8DXUfpDNJPzMh5RpcwoFVIktg4/kKg/+JvSIBQDvMy3Y6cRJXrNsJGVsqBqqp
GZ/LFSt26jNhxMehLysA5/2z6kNNq+BMBg9mknYo7CIXWyzH7Mhi5WtLipLOeJPq
9e8TGwEdStSzQCNyJE8/77hwbL95fiHUtjf4r+mu2EvYRClYJjuOpwV/dMUx7+wr
j3JJqmU9zresq0uuO72qV+gScmEdtuW7y9jhkgHd4Q9WW1Krea+bzJ8QuA9znE4l
fJlh90tzRPs/VFG7p/8cIFNfhtNpbU1d0jQnQBFTWE9cMvm52LZnx1u4nRfQwJxf
xHQYtDs3tovZfIEKxKmfJwxIv7Q8qvxAXXRKAQgh3oUsENfzfjSHccSnL80jwUbg
npGkHmm/XFe7XX7Vz1J+rXXE5slKb6MeI3D+y0s4a8SA1/S+dd8gdRsydm+SQkOi
8NXL1MSlzv0UXSRRHsefU0a1kCZkpZvSpp6np+RiCY8DMiUnu7THIe1yCyaL1p2W
fAUNHbyJof18Yjv9s8FBR/XiFSlK5O4EDTYCDzAk4TrWPBKLcRhFTfXE8/HZo0Df
c4oMz8zgI650p3nxuZsRWlu4RTwx3zZHqhR9ZAC8k1E55a94W7ob2eEuBe3TVUu3
Yo1kGw3a4OnMzlzvpDB0QpUsM5SxgqxEg753RPXysUgkqjjQ4Ta5+pVup/DGPSBN
xDqc5ffco3+Znwh9FAW6wRU67fzGCj3Cizogl3JmQpYTRweSFoeJP2VFK4LodbEa
6fdkre2/hzi8cEQ1KdUJaReBw1vTD3KvFhKr6Dbs54ZooYikTL7wXHrcIGnK2inP
svH7TGAc4XvVQhwq57rGGJSCM5Jg+2+0tTtPXw3Otq1W5wqKhKql8HZwehEV5HZW
PNLxLsSOIcNZOxOpt0EVN5a42tVenLrDzK4iV49Zp0CtP2XiqY/64yJJZRXF+98j
wiLtVgsc94+JekLfL/3WuTX9o0qLxOtmKUIjIWQ7QUAltdI1DXw1fqfo/zuO3aCR
DLXe3E2ykaLb32AHmAOAuB4Hit28UM1PQsKrdWRd27BbwC1oGTEhnJRX40CJzZ5J
bd5/mpUCKM8H+1iQpVa0OUuLtTDxnr19rrU3BwXqurVyGBjIIBLgqoKC1uThBUXd
fm9tp8ZkTLgz004MpiL2zmFno16bjm0NMI26+r97zJDxYsKJYYHTbEAJWgSgp5Pt
aSWChitSOk1PEvV33PMKTgyTCQtMrLqstQhExYDqn7b/1kIfT0UT/KBAPVpcx+0a
riIDn3/jSWSCpPg9Mbkcz6YLpL8oikxd9Imhz//92bsBp5irV6tG8DIi4fcpoDqD
VJgj84i6rSLiMBe5/4M3a+TmVuGMyLtOEbv0r0sJDuVDZSf2N+pU4YqGJVTBhXwv
r7mhCw6wGSnlDLhBq6RgXmvNfjj3113yUE5qaIovqDq6mnswdx91F9rTyX662oTl
JSI8EFikhYFcqlPTD5O7Bxiis3nf5WxcaWl7CuipBKnHnvtZx63R9T/yZ/U6FJ5n
4lqlLoP3J0Laodo5geWwv6nu9LrG3FM7mVVawk/SwutGaSBbxsXI2HUKwAk4+7rl
/upyA7a06r+DKyvSZ/KjL1FnSg6zX1s6jpV+Uk1Snsvas0qjK6j94u48UARSNowb
5Y/614935BM1w2VgGc7W/S235sN0zdrVD0njlmalNsGaWxoYtMpAzdkajeqOEn/G
rFM21T5pOYcDcS6KJ7es437LQqVyW0ccdmNzaSNPlxY6efcRQOReGQrvsMiFVlv9
3UJrEZ2SVgyh5g2QrXDiskETPDcEVomx5DzUGS8xdmZIrt9MreE3Vi7r93Mm3e3l
zcccC4Jpb2V0Gv01lotNxc2/vA/4/uXGMq7whjv3yCbjdZo+wcnvXMhMY45JOQAA
GR8xqjHelrELUH8gTHUuSYWaxkPK4ZTNYOQLAAF+ktaTymkrWXzmu5t4J6eqpBtq
AgXb3K8TEOE6mt94Tu7USjVvwbNZTUcfzPT7zPlI5lqfuobb/ZOm4bxCzZ6M2MQZ
E40zEHoupbkVqe5AcGRqRSysc5XU7HeCDAXoDOJdC0vJHZVevgHRi1NEa7ooYPuf
LnChksekMMZ3XMpGswmxVWhly5V1r1xpGSL0KksFohNKjP11Wlw5wG+UvaPbvbH7
Xb2FNyzf6s+FHxREK9qvLrIvocdWxBFtMkQh2CBGpjxOnJoCEZ3a9Rhme64m8gE7
pp4OBvV3NY4t6/QZE4zaD19wTII4QMdpsTxYzda7aE7oR/WQq6yCYToa4tqMHW5/
5W9CznS3MIiRgEnksy1bDUCVwV+Jdu5zZfu4e/JdfX2ZVKrh9wpzAChHc05OyH6M
TYDetysNYAGEO3zIE90OEZCHrhoCQkvXgYdRAQzSyZ3671xbnwgIyjAEHXyPhlPP
oWA0I7Z8I51zQ+wSIWVFuKt2JWaswgYdv0uVlOP5WEP0ekUCLA8W8MguP2Z2ad/6
TYdTtnR+vTN1Ycfezu4bY3K+v5HqMiR1cz0cZeoYJwkBms9G7fqKUzaYkHwUxuUb
fZAigBbHFwSy9ozRSlkxGkaSlvWou3ahpQ+Qxab6oU9Lv8FR0RgkJ76TuAfa9Y54
O/D4Sb3IFNKfHi0I68HtNrHD9dot2jiFK96u8C51WwncTZBV3mCkJ4aFx8vJM8YY
jPEj7jV+Gfi7vRr8v/zYjwkunYH/8bscbUw9CfJCW/97awa6SFIfE4BbYwGr4XgU
YO2B5jx7M0dZB1f1Qv2TeDHnhLCcUMcIiZ8pRXJtE1mXYH//FufjbrMHtyjvdNN/
2hB31uq4IaqlTOHjddSCA1GFHfUu4XgR5w4JAQ6Gq2zusSDGJHU0K9TMYRwNbhIR
HYV/aY08v6yFWZWZ+/hhCb/vgidB3Zd1qtk//sHrOoN3xsz3ON66CiOvBJAKlyOS
52Uh+B1xwvQG6/QQUM4gQDKZ4EWlVGxuBey6bndDXkRFvTGi0Dxhk3E5yO1CYdsV
DgglgC+TE+5Tj1VIuiPQmlyHDxTuoXQnVNviWpG67HWR/nkEBQkFGeWKjNfgu9ae
YM3xPSUi23o/r91I/IW924cZyFKWfs1IskNBOzDYNM9+KKKOnO4YbAELw55G6aqh
mTLSFXSGEvcQHfZKm2JY+jmYhqpwc2DL1Qc4Vl2EC8ugYyL8EJxsczAb36lmxFmv
dgzRx4NZcu6mfo3VJcVJOZS0xYaLe75X2MDGBP9w7BAZW+DR5LSEpk91CiSlDpaw
mTUllm7ugoZ/xMkx8Jj1uNgYEefCIUny5l6CYM38mHfogvQNZdKzpoDzgqE9YAQO
PfpHug8N1G7pgCyAoqlOOGZKb4GsfTCT1KsHsn9mpR0GY8OwNXDnmipBY9bNB40g
LtFu9Fy+w+LXRJNk5aER6DbgPn2zdRx7yPjTCT78nBG6Jo3cNUCcBzwRxEjmmpqk
QaD+TVyI7Q6j4mYW52UQbMfeAmjK5SsZLCKpthKGH4NnYecvZ+iitiW9KVdleIJl
82FeyN18cGwXk5pouAXgWNu6l1qdB7rX0rz9uImr3PJNX6pKfCJov0E8agnIIF8F
aHaeq44Hj0DGit3znjGt/PYYJYXyNIAYPbTrB56u3v/gkHsfZkarMZKsrp1vgZ0I
pb6q9atQTup8pa9oEG1kCOoiWYwoHFtKy3+dyRlZBpi6MJ/IVGZ8Oi5VvR9/hoK2
tFV+yanqlA4f2iO/LAMRzBEn+dtj4xlUNkI+IgMDAxNpxovZg03An6eZOjPqzK3M
qSVE6BEX7Ph+y2awpvW9JNBOZcrKD9BTegBhFmiNJM2M0+Q3+jZl+RQsUH926Yz6
kuhJTRE9fbLW2sVQkF+Hd4iRU2zYBP+NL7Nwn+OPbgChxmV0zna8ktjcEpcH9vv0
aMwF64i6cwFQgQgYaIyi6bO/skSZAd/l3RTv4tTcTh9u3e0hCD2q215+vxp7xx7E
A/B8g2vS8vAUhCbfrRBi+38q9unvHDRenwtjCOvahZ7DQfB2Yervq3lN7x9NYsSN
A8CbOHZXkbfEk8MV1Dos9Oa1b78Vb6ql5KAWhXqyRa8IFdWGt0GGp0Cy6piclHCn
2PXCui1nKKa29duf9ddzQfw4uUNanLETpUjpLu3UGvQgcmjCggqdTr3+AnR90kL/
rf8xybYuTccRPE4vce0O6VtycDC6RjvMqTwO222EcrVDk1WQHG94cXzn9SXbFtbN
HoZ1u1m4yA4eFL/ZCO3IvV442c0+PrpGGfkIClfRwK5HrNYYJkK2vtAJDAkIiyLS
fOeYOrJa4eyrHUJ4P3lJp2Q/QvJvKQmwSRxfX2LZvY2psLPH5q8BS0hYZ1lYWQjh
PfLJimUQZvhCTZdkRx8hMDQL+PwEgp3DDjqHp9tc0DO0DSqd93KjCPA0D5GRJDkm
yyfPsY3p9R5yI9LrZnl/E/GnuwMP8VoR1b+WrLWOZQhhuo6PwS24IRbo/yhwxclz
9jGoq8FUS1yvByS43dhOggTcZRIRHBIVk78a4hEefICkNfaDAa6Uqy07mSszMy3I
6PTGiwe70YRIHgxspMXoFeLH5UdoEgSQULYZDu6yTERpl0ORDIfEcyh9PPDCi/Gx
KNtjHuzgln1pwg5BHcwv71DiwvG6ZARg4Z3fAUjq5cJpnNc7SZyM2kLxtxv0YonQ
eWWTI/MT6z4fcgHR4AprA3rQWh67fDAgr+Meo8pL5HAvzwRAnFcL0P8hN9Rz0Ecz
St0OKSEdAcVSxFsmNVMxcoImEwyD0v49R68i7T6BvXbVMJZVgoZG2cEsbSTVpuan
wRYYgJnfrcnIgCXErIaGCDv07+EnnaQflAvjnc7XyT7q14V7NSIZDc31IhD7cT3r
3yijk0SKdjg6rqunPF0lqK7kdaHPc7/22xbfs5DprCJJVckigHbOoaPhL6AjcEY8
eDm2WPt2z730tKA0Z0i9YxC64b/bDWqXb4zDLodW858UYx6BzJYuGnDuB88OHIjm
Ibx5vnF4+FWhntH8sfWVNXDS3v/P70jnH5JBbILB5zSTtZy/V9vxdT+Fn6wBAwrU
6+lYQjhuaoLig6XR0l9JE+2dB7M9XhjKp2GHg+ctKDOWaYiVVLxwryxmrnrRQhq8
Jr/7FqA1biVra/Cg2AZofqEkHqvmIEJmp1LHXwu7WQFwLtZVa2JdhKpFg2AxaNK/
f5mhe3k96sI7MJMwNvIu53y9LlHUl1BHIvH0e5C4PM+V4JyXC2YIfkUvMnHGtGQ0
nzoJaWXJ1ij2mIsdSYNjGCwKNL2YkKfKnMeL+2vf9UwjUnjrlg4htTa4BRHTyMic
JDFDVhXFHJ+AtDJOlifHqW3Su8dhYcFL2RqZ/R3Ebj59MSeQWGgAza1S+/GjhAxP
/qO+GslM/eiDtqnwuj2qRxvxEYdJ3UdFRZDUVA0Ecop1S8ZGP0TGQ9AiRbZRoV5U
1buLo9E6Bkr+yr2KsCniXRLkTSJwuMd1d6HyG4qKMYmXXuPj0IJc+W7fpZIRz/fQ
0hNhlev+NcOsscFJqoaaT2lV9j5UHCFlkyw2cZrVovqAtRyrywfrQrajxY1SyQua
nn0AhVqoxxVVVSAlxw0NJuwJN88wS2SzoqMU8OFvSyJsGyAZ2RaA738cy4vNJYip
1ELGbhkteqXejvV5cYfdzNirSJCbfrSHhA63LivRxlOROJvYclV/mqQDdEKPNIXe
N5hP9GiZ5bOiGl1ehzycZIq9AEHZhlMewI0SvPgLc2Qds4JKb8qMNNPBgnX6vejB
DwU5bsW5DQymKkcFvsSXpFet+wfXwXG1u9rY35pntvVcJlIWWYoefgVMAPrkehNf
I8sKAS2ICU0Cw8ohtdxTmPWPQvJ7sjHw25R/ny1WnIJ/AmDJ6MDGYg2Sk2DHPj6N
SXFlPAeYnocUE2tmX2Wfr/f/zR5m8HrJL1o40cly4RdFa/CWPQEQoC9ZvJ4vKbnr
eezmlvbdQzEEE2u8VjEvHb2XXYnfnu8kl7Of9k8C/gLMky9M7UfHQ5jqtfyKVMUR
2l4DAIZB3mHz4suCM8+jD4HG3t30q7NcxZ8Gn+FSZnhodl1TtDXolRa1kN83G0uV
LR41sLnf1BIEugjYGvzepcKiD3qOXAKHMEojxhv+8nqQumTkhkfINjGS7rSKmsAg
Wp4piOmyFRYv5N/sklQm9NsERapKzKlTJkHIIiu4ZrB/xXhxz1Kk60bRvtzqbSeH
dRPgT1WPXFxg6H7Qdm5aXHcCofteF4RweXtBimKhUsms4udtKRq9X8I5DZIPPIa7
W2b+eFmgw79F/Psy2sJHO+VjzCcwKm/vYuePfoxPHzUjtYS+Nu05vC5R32V7/uYP
qUuzgX6PAPwWEavQd6UB4VDQsiTdWGWgeWB5JIRoJjKYMHklWbLudaK5Sq0AFWUB
QWLSQsE7cG05vlyp7oTDBZWySRpKi480YaDFIXVu64gTp41pKOVu3DhSvdqtkMqE
dyJQlP26z+k1Yf+QCfvk8rf6GQ518/w47+7EO+b5xESgnQK3rdZIfoakAWlJuK9e
3LsZpoTSJfPfY7yrHsPkZWM7BsA0CnDVu1OT4QBqNI0Gq8GqZHe6X5WqlWp24lVT
QsKSjYtGCBUPQ1NokbjVx1emvyDjj3/NW6r1QE6mhzLCtBoBZyilSTrkBTe0OpKx
/BUs8iLH/mGZaogZ78Ne0+eTclLZIeHODDH+NF4PqZlWSlJ8YAsKwEq8uJ2HJMt6
mtYz4boqgDrNSalWpREVadrPjzY+P+TvWQqnsugq79CXfIe+bFHnrBlqpWy2wMse
vGX+UaCP4+vy1IkaQapTgRRmsE2UuRAAQd5M24FADL5U+gi+0N0SJA3vIdd2uxXx
S6F98aYnFg6M7BRu7LOOCF9+JTGvNDF6i/iVl1DxaBwFuIj0k20QvOtmNIhA/crR
/CgTREaQ17ersPJYRHjzeglA4CjXWRecu33lbkinOO1w7ck/BXlnCXuV40r46a2a
V/g3Pr10l/4irGgGrNqng09fVhZ+sziMQCtZgrfpcGWmYzc7vi30iGky9IANFJn7
8TvoWTUQYngtVpRRYefsfdlTmKUkYN651ydd0c4U19uqK88erK4O/9/iA/3qd0Uf
AxL7s/UQsSbVMxpsmSz3jhBdo9ZJMifMG64W4sH9PRCCfOhnEnsjJn+YHT3Moz2F
RYJzt1ONJroBLD/LZtl6tCM4B4fPn0hFUmNT/sujiXW9A7djfCYOfDsFLv6+wpzs
S/Oo/+unz07QayVVPTskmXokqFAn/ufvWUlLOLcajhpPE/6po8JzwWcAn25eMjCO
2q5sBbl5/UQLxFsYRGNOg/imcrznP3G5C7+lXa16E/cpRWKGOqgvV2HnEbOdnzyp
doutW/pqU/w0U8+UJ4tv/otRhEGmqcGcdk0a1tPcgBXq4NFATPuZ/xPK7m1RA4qQ
gANdrQQrrcVd3cAd5StcSDuP7our+HlQDqUU0JC+bpqWIv94Sw3wtic4Dlz6CAFJ
Vykhg+n5T7u1hq/et0KJaAAM6QFPYUzR/N0lO3+jLbc/WZi/Y1Luby/9oTbvxNQ6
UJx8uUsIISJZHH1kQsgEFE3yiUy/AKZm/YvNP329r8fAcSgEMahJwYTZ23G3F+vl
edzISkA5FR5ND95Rik8B8/M48bgDAW9q0SZ1uNYvERS/YsTuMJeSS4msM1DNuzj3
ttyv1olBGyCrcfnfYGPowcauts1GIfPMyXbnFCydQIHiWlKxvFKLakp7M02tSQQI
qmiqEyuOZhGJtVPIWAK3zBKE68NH/DuXHnAd1QgYZBeXaex0dsvCzVlAezPZzK+n
uo4Z/KQiMcAtxPYeXjfO98aSO9wwbiKjF4m7gsHmZfzUC5i1kOR5y9eXophF4NSG
XC3LwvJBlEsvXGWXYHI+6Sj0bIR8S1pX59cRbfg+GaXQc0QmV2GIBQ0pZtIzXgFI
zlfu4/S6XsSIk3rTxyETRs9rtAYcpcSJuBV9A81sIkusJouAOJz2erkie/r8JbN3
2NQT0/ViJLeZtwfQ3a8F+Q==
`pragma protect end_protected
