// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
n3O3qpB0BY0JHQUmmido+IL5MFFkXox7SptPxGelBKptVpa/+xKSvRULPF/pxjMw6dpUfSP55t1J
AAH1TSvu1/V/jBP60JzP7ZSrp7peWsP8ZaJd1rVG4CGYH0lgJ78KaUw0RyHM8Mxj2oGarK5M6uz4
D/ss/utuTh0V/cL1I80p/i9VJcIb7P/y+Bp3YIKsbfn6qipFoeYKKUhYSUkMnAp5bANdMPREC15e
dFbR1tW2iuUlKDal1VAbDXH0GurEkKvwQBnK1l36FBU27snWUKFmXohQmKx1km9s5oUaUHwM/Gue
48c6YAFmdcpTbcW8liyVZYhzYMavgJHhtkdrXQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
igT+9V1sPxZvAEsa6LWr97IT0vSbQE7Pl2e+YqIij5hl/9uPLcAAy1l2MQy65VLdq9kLAtqYZ67Y
/1+Bx+vOCU7oel0Qopmh1Ow6dNM65DkWaZj0P2YP6t4sDhFFJOiaTDJojBtpqVLztJbh5rUjez75
RfTGCZkIOClSV6fRnmbEf4nfAOZzkjUX6sux74CCC+fsg5imTPaI6p87h8FP0Vz+PWVMcG0WxULU
0C7E8mjFBLP+6XKEqD72LQc2d63xa4s7sEiNm+Vtn3rmcJ3UKUM1r9FhV18HpL0HBp0917+5fcp1
Opvqkj8po1t2rLnjBSNBKrAsYtErttkhpfzHJq2FlVXostpMloo6hrJ73oewEtZuRP1gLGhcFRzV
561oQKKDoo57THQh0GpFq1pTNSaRD+v2oZ74e0Ppv6Gev+hxkY40ITnTCjd8t6wlTFoA2AqNn+4n
D1QrvOncpT88gJ6wJvIIwkZVGwXw9bURZY6akpwot06HYtdRtib03DuoIY4smaWYWq/Y/0f0pVV2
yJGGSLpupf9cuM4riJoMrgGrT9xgB6AizEVd8eKKvSC1i0/Z1+WPZOx18oSpKtmaujAvZArcQUIH
HEiCuIkn4bnS7x0PmenLg3PSL5zzJOAZ5PdsNB6/n2MPSwkECKNIsYNzEPlZbJfF3tj6ZVNXUsHK
ChYjAV0F9NXnEqswVE8JVDZJhW8JEJaMlQZBS9aM3OlPWTWQdusXjuW9DxFJZiFesuhiZ40EKFfB
l9nkmKCu/uJE6AJSKpkkV/gXeTbWL6r2lYBwf0G+ZQPReqAkR5odcFMRVARQo3CFY5+/RdvEbWZP
N99qk9cfBHgC/n7cBJsv7RtggaSsoEVYzzc4NgJWCDYygj8f1aLZo8nulDY4uGWQ1Q+nIRzpc4fr
kGeCozZD8fFILrqFvPca/HW966LzOwI/Q0ZCaoLPzjvNt4HdYTWa5D0Wjxa4k8FwoxJFAJJKKRrX
HW3ojEM8Ae/K8jkBxXbHxUeQ5dBp+5soU22CoFEb4+MT2MrnAPEfVuEaI0QAxN588qxGS8cbFlYH
YEfxnNWMc8vB9H+iDO05LljnPyOMuvfwyEKifimaLcpEGzVVtiPvqzSjipQPRgzopjWa0Sxh1I3g
bIWUgp7OYyVzlb8Fot3N7+D2WPRlWxsUDgv0uMXi/WPmuw41//rCaBSM/lhOnCQ/6BH+5z7des+F
xkCF+Rfye3lESt8JMri1xleqcmDODdFP2ZkW7NEOAnHp7Rg/7CtDc2OPJjRxE86m3wOzgRzkMAW8
rxmwQRFay+GQdOXGh3639GAf0p3ZPOdaphc44JEQ0hV6uh3Hg+t1CXoEvwEfwcoBlS4i8V+Q1MFY
qSdf0BvJPIViCX1ke84PbkYvmo1Gym84KH0jkV6Dy74W1vWfhYwFi266qMK5ztx3vDMWfLod3NXZ
2GhinYbhqTT1qT6OlHMMI3gUt2RjvJ2EQIW+3DrVqVtJm0+YKMWWFj9/W7nharbG0qmCWhsoMT/k
HLSA6YPdqYXi0y7vZv6yhY+vk9hJ+3laHA3mHOYfyHm78jRck8UtVmMvrUiPMViWycF49gjLHvs2
2nj526fyf+I+Siw0iloZvq3DSpi+ZEnZk1jn/SWS9hVBVP/sZXBGzYHWeWIkP8hzWWOW+RnTX2bs
zhDsYWECkQsjtHRAc7y67n+wExDeW7DBWSYdOqgPS4vR5Ed+zQ0Wdhvq+ER19kV3HyRCBpbHDYqP
XEvHEmMsfugma+iTf+JubWG3z9SNnf4W7X0oBagplm7j8tasBpC0Uc6QPxJ22a2JtWnkn7kQOxYK
hM65GspBslnDB6UJXdxryHl1MY1c5qJccwc4DKN3Ihp8Y7Epy71LnSBl5Ei9/ptoyS7gtWq5Rlxj
OMHJsaCl1ncmirWhXvr9wKOAzxK82JShrLeM4UL7QrCWnCpy6odafZIQeenA2z3yRM2TQtkOykwb
XCvjXqRHveMWYgsmCsXTqdxmUbJz4mmjfkVfk32ISKV+AKlYU3MoXhn+Km8cb++EpEniUt1ZIGb3
zU0BtwfF5b40QU0jiuZi5Qg2dW75+n7wLtty5Q0NJ1B7i+Veu81arjgZaLNcm4opp6y9e0gpzrPL
k0yNoHIJUJ7FOhGktR3BTIK3lSJ9Ai8UUH3gXxv6KZcBWF5/S1vh53VTX5/AHDk1L9ox/osmEmIN
IgdFX29rlAZGe+7Oiy0NfTOJBkI+i28MNSKJlXCg2/7mA7Hegs34aa3Eq8VEFhAcnSVzxlXObd4S
PWE5odaG5iIH0VNncCmxBK/1nXKhMu3Ig3Zrj4FyqmSm2kYeFKiVLuGi0zSrU+poS0jb+hTjwStj
j63Jv0Y0Vt/0+E1H+1F198Tckmn0ipgmcs++b/Y+W0N9DyTWRcvX8XQbQ5Ps4NDmawL7NrtyEmPS
Pm+oJenOaej4qLcqU1nxE6QSj25jEyOXvgl3cfoEQKSayIeu+eSbPO3437gtE+d19wkJrWVS+cjI
X4rPxTrDQHHmJBmonLh7fBNs2KCXAz2km23II778BfqhgdqHvkVA0POZrMa0aD4s7QgqRNlcnw1y
Eg5EaroMVOEACoqXc5fr1cifVPLcm6eJFUYuiBlOyAlzunZAu5/MWhO+DTZLLQgir1wXYjXEYXMa
t61nbwtFPwuvijGhk9zOACMIvnf21KEWFXFT6kcGQC1fh0nygSvYMrpGOnBCDofQ/v3jlZP5+3gd
0Q9tZHHV8RVyuJO6D3yv7zfPVbpt21yvVkWygJwJoH4lCW3R+3esddkUlCxRvHjBjL5rPknoWINC
K7eNGUJ2Nb8gLT4cHfrW/oTDX29o7Mg+QQhMlmW+oOzknSq4c1sqHbmVY31JGD0bGSIwckB+8O5/
jejCTB1cwy+Caxd2gaqFNPtgDR6Ddbzm7c7d+T6OUq556Zu3cEutPwOUY7YDcCzZ1Nq+pGX+dx7T
6FGq0NSNE3vhDVj5OmuTorROuwUGB/HMQfawclPfvBBaS5d+L4LCIXEVrVEY4DI4/LsmxyoXRjZR
YdD5gc0c/JdkB7mJ8QrFTQCNCfzF8UDn1QXQpSwuhnOm3Ipq4E6j9/805kxIqys7S3r641c0km7r
lGx7kEkdoDxhSMGO8e+83fYTviCk01aj+S2GpiCRUOIa9Zl7q0e9b5R8Y8oj7nPZ/QJeQzeMHBBe
F0k+4qL7gAsdrzwyNjJ5rbaLbATNDuhnO3ijlIYufDX+A7MZ4jal6KU0UhHdWuazkEyiaN2aU8HD
Zd/Yr2tDGgIee3Vgg20vgGHirIZzH9pbabViAHv//aPDVM6ph0QsnIFjKnmO04mRrwHVDdLp2fjT
YoGUDV7HSmHFKXTv5+MZOB45c/ElAiom0JY4TpjAXGqvKixM4tjpv6w6/mrSLXP0lBjnoYrVBQUd
MxWNlAdESBENJmiR5qwleCcWTSu3ysK2n7EbFAhW4CHbkq/LuDjbC0X5utl8MXNvL6ufisDHKI0D
qKKh6MG6EYfeycXHXPcW2xNOiBNo2qb0ZqvAb4qlGsiEo/8HU8wVs0dwSFpUjxbCDvnd1LPEYKRd
1oNrFQuN132Sb9p6lCiqWKLbdXCFIpTIVqBFykskgTYzLi/y0WL/qBT4daCmNDGyVNYF7a42YEa6
taQp1TJui04P0fdjsXWzpnHGAqL3vkhI9uQXi5aZbLbUH8FAxWzb4S8dRChQ5r/n4n0WEgxUzlRF
tSIhBU5oA/VmVX2bCV2XiCR6LbjM8zkVAOZN8IMMzXZzcLZTWR0IC4MG8jC2tQMmAMC+X8nKdc5+
VwmZPzF8xkUff/zwI7T8d3yK5y9U4e1BE8ddA6gKyJWkw7qUDpmyftU3oBOUb0oolm4JnFPStopF
sI1arjufcAn/dv060u77dQDFds30jEAYYs15PnFBo20jmRUg/ZMnOjSbmdYIrd/3xIa1rhH4h4UD
g5ucht+8IRErFGlTa1HpQQivDTFCl2Q+vTUUgA2CTGqoTXiqUp29wXhe/1MeSXL6YBMoaO7WyqEA
9p+r1MFOcXdvwlUHd8ODfPs+9wI389KbDpQNzDbWj2helig/mx8TQETYNzrYG0fEexU0azq31nKs
9rCMoUlgc7kIgWI5j4W6XnPhSkUTmgZuapwC6NaFouhnpfnvfIpiNLo9tGs0J/BQFW2TdHMdZXlv
LqPPr+Z7ynohZ5n7+HD1PwzxRE+AvlkCKv8/CeidwNpK41SU6IuAENGjuEYY3cKBxmPF8MuL5EfV
scLMbP65CSMoDEEmzJJEZZJZfIQrEczoNpuNEdEVbAec5T0KKRvEoTEdnsY0XMCKbk9XJ4IZrRBn
1rUZQtOjuHb7hHzHN5FPcyJ6fwoz+bBTSM9fBHawwCFAz3Rn3OUqKrwt2sDNXMb6GyfiO2nj7jeR
YUKc9YH1ozbVzKek4in4io7cP0bP4WQfO6W+AxmLL+pE1pHf4QOYUIilZWMs+Xn4DHMKDonjZYHF
LY2YmWNsoFePFTxc88C41AKEWB4RWghN4Fqt487DhDwcmI5iXqdrsRs26EfGPFurbExnmtjn0bv5
ACoTlSTK/BO6VcdDX0FgkF/SnHOmQKM0jTesabnnZZDdokDDaihsfstnicQCwLab4Biek3JYgHWt
Qj/ovT5/IDZoQrKRlnDF7NOgc9RxsJ8z+6Cmaikt5en/8r+nFVIXXePWigz/7TOrb/X+hDAxnpej
kn0anIOA0SW3ez/Vweh/hWu17X/hTfMI92h/G2W2qJTN6Hg/YUJsGMjJv7HSlY3/9kGOgVas7W1p
Jdhrx6GOh2wxpogWa14t9W+f9shhREIvhNWtXkH7k149MB75JbrIzy4a/Gt9Uc4/BRBfoxcO+cbY
fYBskdkQlQdGSiyZjvX6rA7te3HZh/3bOrJ6jfYkWEWWu4PogfT+Lxwsxp+7V6xdlEb1M4IMDbZ8
bxgB2xkUPrY16dJ2cimY25EFXZQ5Peduc8VZhdjt8acXcJ2SbUCi16C29MsnMfMs/CqQMYaB0r7Q
yuzxoSuWL8PAtS8uwQpS0Ljn8/z3DwwrSwxaskZM2sPwhbNKJz6ItlMGmo9x/VYqayStl3V9x2/e
XM/jkpkvK7LmhHH6EK6XLV1tmqzrUQpFTFS1Hs989pPqZHf97Va+K+if4bTMcVmGWG0h6pLh9NQE
lBlWyEWEGkNUvf+pp/VM/j1YwYFDViFq/BuOoHP8xbR3Cjj06yE4UGLB1BbQeFp4fugZGm1wDi0T
+s3KO4NSNrgj/BdFiLJd0yesxo30x2AsXyD9WeXsom6Pm80TaAMFiQkm2jIAvkKt9d9JWOg9vGC2
lJr2tgkc9V19psc1yohCDPZjhHj8dD9tCgL5i6ESnVulVNhAuVHH7+XN+ukVfZvfPsmK+WMc+aff
HtxohQX4oPEqQ/yDyaRwKfuWK5AhsUcJMNcLPmEuJvylP964gt56Zg6ka4sfVA89qJPaPlGY4tbO
sZfMZ+9QadTk/uIhtciFOYxVUGdgp1bDmka+7nC9QHpKNYDzg+YFWxaPx4CLGaCKt/1An+DuC/rN
dztQaLf0hZZjsg+0YlCNEozQb/sBhsMZtEGACj9Y8POPgz8u7fZc8HRbw8jW5m3oliuzVrgHOk9y
XfkN1QgVnxj8o+y1f8+D6BK9TGjDyXs2i0o1lb4KjULq5HfGx4c84KZjjgePTtlIDpjCaywFwgFY
OjdD6WcgFfAlCIaXR2gNy+4xBJG+56h1O3bs5uSE2Ynpgyj4qCmIM1l/rxttf4Z9rSEkLK93J0xH
xrkIRIwMvCcnGnjLctnfuj+vO3KKookh2vTtSUd86rw0eAQAm8K+xB6hefmCbIa2S0fl+fGcDwe2
mCv8s43G1kNkuaqeJfQHEWkZ8JX8dN4JiB5baBr2f+pikQQnE+bTWxrEdMDJ3FAizOM2wKI4swks
ZF+oeUMWTD8jwfNfMbKTJDGom1l2aO1oNKBfiMjhlOZEWLTU9+P5CAuiF1R+WidG9CIvxD202uY6
Gi5EMrXrItKV1ZdMUmQ3XlDWtFoSt6bFoP/mwUrsoB59b8NJfKlVQzYs9XvM08x+lwZUHueGeQT1
GIblm8NHkT/tyqFMSfBnF0JQRLeaD76t61YOyB7ICN21hWzpzqd/IGfF73bsZ2xIG3uCMlRceq4+
HdZSnScOnfW8vSBveIHSKAogbXPhDmBaPKqpxLuDJQLPTH3OX12akhedyDDMyo/EgD/E+BZsng2/
GzBk5K5P54uEBsUO/Ft3GcVix8leLFdJ4QYbqNC++ILddbTUpNWG8e+4h1CnmEzuQeZWx+kcxxj1
BNRST5VNBP2cOYAw+IfeJYa6xzaFGaU2tkZS0ZOyOVRi7MsJXivuhx0FKm/wctrSxIogbPga5qea
by3NUUZ4S2M//OjL+Rc2ew3YiL04zEIjfg7aMAqtKgJIK4J38ISa5ir8sWQ0NPAT4q90EnTLn+f1
A4SfhkU1fo4St5xigBtNeNz824cBk3YfrhBJC8xn2cLm0RHfQC5DezvXEgkRuiM2sLF/6tptOTVh
kyu7+OxC3lbqJKztkKEjXTbWmg/nadJbeOT0JjB9eHgqr61/hc81DscX3ZVc0FlxwuYN1138ycPv
k93QVJkfPjVKoGpPLMRVAietXCyf7uXHCR9w4M12INHhmwndDb8oOv3AatUQl5nfGsOtXlOJtyou
KPoE1/deULujurCOKGtNg+1/D9+DYiibwoSufUTvPqeor/JLBQTYp1mSSIwAh7Ot3LID3VxXmLO7
tv2mW+wcH3zkTRmODNOxvLOXwigQSPGpU2Bx6HObdC1WRQMGV+GKnVgMC63QQsBb9VyWgHmL5+R7
ARTQXJSyMjgj3Kw+0cjIZrxIjH9VkXpSSZ+xmTZ1yXTYjbwIOgiU0DYrNIIMVpZvVRCjmvPQbQhj
NFam0QiLooVVL9vWTA/qDj23E5SOikD9XoSSD5fA/1oPLqKEQozvviXOC0tbb+BRAbyaemLtav7V
pu/XPaoRp4lxDb45aZIIVgcIPZA4mrCwv/1KMlVi13+bs0LZj1P2GjnochJnVRJfD9S/PTvzxy25
YiE/5GxFn6894jPZDEuigeAQw02fYC/5rAoT3QLkERVjLcUgJiV1dHU4sNxO2Qe9CQ4YSBjW4frZ
y2NmNHPBtCUWjoa4Cv95ge2q5QMXChVRKXaWRh6VyyKsUPKK8OItAwExKIfvfYpUnKxnRWDPCrrg
c0oKyBB+JjIV15KRkwIhppNMrSAqJShb6Fu7AZtWhkWQKJIwaUjovCLNSvplALsmBOjdjtJfByIo
aKIufzipi09bkk23uEohG0kQGG9zOn3y0sQt1zLCJOBbmMxW2WqxiWYtcFrpa4ci
`pragma protect end_protected
