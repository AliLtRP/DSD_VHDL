// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:05 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LSrQU6vmNNNpZ9HQ30wRdVVEU3xREZRTYRnrNnmZg8Upmh42bP+mLfSvLJg8eQ6U
vW/7BdsjUlZZx6/dutnDpUyTALkAIKSR2F69NtuHyYwgazRzhsnRQ6gww7jVyQ+L
ZEXcStFoZAIUr5rfVFPdwilb1G+F4mRWHJoVno13Rfg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17152)
SZydPLCa6M3CflJMVEcdFgQqssM1aVWsej/iTyvSBMceKxp3yvrXhb35mkwGWX7m
XhbfVXJQhyniLK7cXip/PcX/OFJTAGZ5RIaUVWHLdBIcbDllk31WmPm3EtL27W5q
5M5keL8TrCqSDWwSOMHKPhhIm+vtrStk7QiByQ3XtOGoEYmPUXGzPDc0i2Mq86mo
ONCf/Tgxavt/XkihQdVBr9m8K+vDZO7TkJYLPa6sRWn8eZZtSigy6IcQCjVNMW/V
PiHhe0e6Ej53RQFSfGQ5rSqhRq6GkbdU9Qa57ngUG1ZC2YcJbTi8w8Z6sDJaOz4L
l2dkQz96TDV3y9XS53AxnYc30+lCCKH9UHAhxTDoK2Kyk2y0j8wnHvBj74hnhMb1
OvZVdjbk7I6ujiv9urM0yzLAvESKbVcBTJSsb4u3hhAgMoAXGkIO4RyhxfNviuMz
RTVnmTPjtGxMcdvTmMbVXvk962YGq2bLGoXoPsed0IwwtQx/oG33UptdJ0/EUoSj
PvVZkX4nXbmrnBEliaxmWhtukLWL8BOznLjZ1JIZgD9Gg/ne45MLC5hEsgWssn+4
cGhj0JKIxXRXlhwWrLowhvo80M6Xkr951CaZ96kbh4bwMba0znCIy96uVZUcbax+
NN98pItl5hJ3NrPMs36aziHkOzw/8/mGIAAPepgKHdfee7K/ToR3Xf4hLJm3iIrk
ZG3cHisl+rdNuYG7KPY4KjqFCQ1J8CtlhEdzh//TaxZIYWlj0NDzzgn0dfyHqjRv
TK8xaSGcsrD5Viz7PzK7L2KB4ht0fyhRfmJHXcj11V1sTwWv3t6mT7rsadMSQ0vq
33gmDp/Hn4X+WYbelTG7QZtJcsY8khsVvKArgBjLvdkgC/L+EeTzCXRHutUoNvdx
cBe6Ha4HJnIkc9FuVgyab+jDj9LaqBzj8yf1HIjPr3/KTCBOVqMrqJIOak7pioZ6
vISRj96yneDaPbFVPsubQYnOM7sS2SUwJMWyWGdpOVQnae3j0orcogX2qQkB35ki
mSgok8Vpv75uFaEqHSczCmcIQ1HTOELH7ixdTSBwM87eDs5qwmN+9zTnLnKvnKKl
MlIQcfa+P2rkneSj1M7I8fW/S5uuCOfUVwNhgI69XQVrkTzDA6sHZ5GZZS7V/Qbj
7ngTRld1b0d4aEyg4FKuJHF4PJVQV/d6Gmq7T7OrIAfO+7rl8x9E0VDxzlCx0tj3
DcRfAjp8g6b1FwPl3ZTnEn1FijJS8kKRyZ1aq00hG7+ITZgLSkUcULE5uM0BXtIF
E6/v5TWzf9vwgREkA548miXC643ounoJdQqU3F04sxaA+vrV75AYnWzCwWyux5Ce
GjeuvCuieGVpiCRMINtNd5JfjiBysKtx8dKYm4jJLIleR5Qo8Kk9S5fAA2M1e4cr
X+Q2A9hqSG+dypoBo+CC5LarVS8QaeytDjMGUMgtp+zZChq33xUuJ468vqRtb3sY
R2ZcxcjS8GDPEJu8CylzpCo9KFH3D9ph9hvjZE733vwHoWdcgnmoohTwB1tacBcD
gmPqlX3yq/YwgHy5jG00E3LoIkUrHn+TdNGB0TzTO5V8u4+PX6NcHv0NgXh2REgY
BeH+0wc/8IgNUiOa9t8XfFRQg+uXd4VLppazWvxsd9h212eov+6s29o/kQgYJyBg
/Ganq/R5insrY3hhXWeW5mK5Zb4q449GSeJvixmZCm9w0Ib78ymWkHbGa9BRiJS2
qdkazhw4DzgNNqrhTBPBthKwsaye4q9cmIWk8dOVtuyt2Uu0PanP7xf0WYdlJRaJ
vIhbM7NRMaDEkLP3c1Nz5aLoL1HX45vIUc5fxOcX53gs6tFlASvMjo3zM69/lDym
oD8MlzeksZki9k8XZrn44ISQonuETfL6LyogTl6OPlSbOHBTREp7/xPl8KeIkFcw
cVogIvYsA/vKmJdtYNQ3JwHSgKskjIvlA2x30nIm9O1qacK5q1fMYdcxElbsfnnX
LM3w0i8TDB3uWhDurzC3Kb8wHjuikjAzpz2tJUbfH4mKHESm0dgKHZI0TKxOVuz3
u/VYGmErflo1153Q8qs6lwY7w+oVDlHtHn4++BGDx8L1DqD9oAzE9cnELLUwVdGv
ay7Ry+WgjblYe8wON67+h6S5t4TyDDUiI6jgLPqOVRegZK5Qw7ifh7ayLFrxhXt0
zlDOKzmKdjflsdLnrGV7hUWweJnESgfY0QPEGtoBVtLTTllNAY9TA6JRuyrjAMqb
4YTwVrH92yyNz/RW0DrYgaSu+7+K7ceOyRHuRdBa0kW/zOyxmO5UuFlNVNQkrt8w
zSGX94scovqENPOCyi4O2bX2aZF0JjKu6MBopJJfZnGUvcqiJqWdaBr+Gu2oZfxy
QqPdc/2zT8tVlaUppG89bCsby3CgkvX4dliQwCHb+CZwgnIubsJyaKrcR6Ub8Vz9
8bHlLBeGKCHQQbaMAopb2hBnaztHt7RtYPX3Q4Jxb6r7qu2i8KNa8/zQNms21IYJ
/QLAw5eceFbwFuim857t09To0EYRMVPBuVcyHO991tNZT6CmytNhqXZpUQbpy1DL
9y76cY6feLa19Dox5USCzi9EIYruYjW7LhNp6alItJJhxto2e+u37MXvXQDr6gZA
/zhOUdFfWqjrOva2+SaZPQL3UvN8F0WBwS3MWRtWFRphWqjpqk9r2TFM+Bo5bqgY
djN6SiKJyh3clgTli4nKqdwdRV/7gIGgqyL/FJUseWnOX8WnzMTraDcIsBcUosgv
GTbLOvuOwh1+BeXJbYH3CG7/ys1DIMPKXHGGTS7PQ0x466oo4Ldez9Hpedlhi6zj
I0mhDo7Z2sDOK8D+a1U0pxGrs6dsr0e/C4D6i5qnO8S3nJ7xyIPAxTydLKWMbyqC
05rNBOapYd4uKnQdy3WR8so8Yz0GR89N5oG8XwS5RlN9GQ4xXzZVuyFaRIB6BPjT
cN1Ju8yfCVU4GirHoziv6rW0fVBUE3oncCAOhASqvvLBqriFwjuWnh8fUUWiYjBz
CJL6r4Jiq638pWqAva7XjnNSUcwpywmx70Nkk+260ytk7ggDbHEa3l0dgL/zyPAw
aX2sje++nSrUJzwiXRzUETFyhsor6iobGDPFEZ2aosqRxrVq+aBwNMc6fhOScnQA
f/VbxDS5OnKRQ0Tk3l0J7hPXPCOPVuj/9pYqxGFvmVTYz6ijB1dKm6k0Aaqhy+UF
zxOMCWNeDuWRSeWiFGZQsplV8TNk6CKCGPmtU2oq8B5Y44cIZE3pfeUq2xgKJBlh
sf8DyMCItbbDgTC/wUFAU5B6YPf6hRwqmx/NNTexBbrBEbEDkIPOwWQ0sp1cn1fv
mTpItXaNc0JFgL4z1eEwOUtafrCnkt7tPjFbWRBgFpSktv4esm1huDTowOhxIPNf
VyjwDTXuyvZaGchgyNIwrrbeV4kOoCZUU79wnMfQCgqksoRnyl+wWdhQTp+S5uXU
OBJ3lm5sG+QMCwOKVwXFM57P9jJCOHLzAkd3LZJC4WQbUfYzHNx6+gtUc8JvKs4w
1bKo0A9efk9lFvCkec33mVIUnrD6U2gGn1vjKytpbtSJ1rcNauiifwAEd6mht6PA
Q+wIpTEb1iV0d/y6YiyPC8AFM+eaQTX2Mbn8rrpWNNXvr7/26x9YrfAo1QP3fUSh
hiaGCq4Urqxm+deN9w8IUGHxeoQyGDauPg1BDEPd0NzauUz0yK22I3DcD9W5pu46
90zWrWypM8vazLtfblI3xPZjBiP0K1nPvTpIccEqNzZbpI0tJ4A/ULuMEIQr+Ljn
BOzaSTK5CkZIPIbrvoEd0xryUpc4QlrxlVUlnMXNkVifVbakPfUMqQKnFRoiKB7y
N5IJYYHLbiXzNS/5fJTjJRra3ZFJcRNo1BB+6DAVgwsRmmEsAknSikSsuXtR6L/l
dPwTP9Npfi5cK84oCguBhi2v7STNVOxmTv+rX4ZTt+usKEwGsl7eMf2q06p8CYU5
u8M0jPhe4y6lnUvyRLaLqgVqDaGmZHntS70n7AgMKNv/quH8YL7eegiiaARQObKi
01CUW0biWb9aN2fXZCFrBJZHteAnz2jKc/etqVmAEIOm3fjpd3bS3OY9HqkHyc+5
iyC/VtpAZt1t9nPHgR5X24o67ckV6+RwJIdiAua90Vbul2eI/HvcY/+iJzdrFTte
Orp83RBU1xc62bI8O6zDYRCkOX/MHxe/+tn7rE/rSaSPzkBoAqA2LLh6zIpZLC+q
NorvFKF2mpI+mhe0CTAwoNOqb7f3f6VnEHlxXzXO8CKgbWpcY028E5bVm/L1Peyl
gkS+pWf0g2c9V7bQuHmT1xcX3l/a8YSmytpJUtCRD9ehb4S7XGkcqMO8AmrEtdxy
ZQmDQuYg+SaT4rvrkgQqwh/7RV6bUwp8c4FjTjyK1ygoE94qpFtSDrfjCLcIpg8e
K1/ZDD6cifbyHQWrUZDxeSo80ufcwV66YM35rplYB8nWvfJcFcekeDe1SN/VHNdx
TRoKqJxOl/1N4m6W6QQAgBYaxJELgCmM6Q/Ci3pobOJmfSOSPB5PMuVTi4vuk4Eq
zx8n3MBGEhxCnDjsR7OCh0VWteMhnSImXhoLOZHK9yFUYEAxd6Nm9YA0jzM+NqWB
uDbODQ+MZAXyO4AMV7f323LmI8bVhh+ATpnduN2dH7XjvBj3z61DvUsOTSUG82++
L9BfFJ8cPjZfRFeTYjTyPQdAG143OVxHZ8V8h5t0ox6kgXIPgpWA6XF/Zl9MONkm
S5EwzUEgbZtD5hINXTB0DyKkH7oeINzPj5MkZ/cWhplnoqWQcskkjTKJxxTnAMjy
yi70Ggd+iZdJhtG3sUn4V2rT9vcc07SqXwnkKJ2mSUOVNWDYV9V7U5OSdOgl8woF
PLCGI7Nf+jOpArrVKBg4KFKpIFE5XpL8C2ISGeU/pQ6Js+rKvIkj8CSe2Fz+JmjE
JQ03KIx7YiEjatMMwHSpSgtv5EocSfj2kV7eAB8CE74lH1c9LMn6jFzRs2zeSfCz
IWgcNs91PtZbhBe6qtH6EJRhfJPe0i23odS1naFnA3adZzR/SponHI6Al7S3V30n
160mGVZ44fwjLlytCcPxpjmBI+HBRc+XqdizWSgZth/uzBqs8nSDJSQFh6OwB4+U
cBrH1fxCRUWdOaIEU5O6m8xY8QFWr3JlbOdN95tTAnwy+vJX5VGurNZYkb4rl1dk
QICLJWsTdumBuGrM5byBGej/b4DHtjXCKARWfoy3g8PUKZWlQ5hjSfyCPbPGh4AI
q9d6ixdut1D3AMuVMRcN9HCmE80rtDxZyUzwlyKh3I/L0qc7tR/WQQJTQuCqDd3U
tzMdcMhms30pR6iY5tVM7DmXBmOnpxJeSDsmhbjJRXaD00l87KMKLYLhgPwRqAFM
NqvBe65UQhSNpmz8HLB6U+BHX5su5z2iTNxlriJ4z9/r+q7gISm4jZqVvAi1clZC
AMlSaBtC9Qz1f22K3OCVxygunhYmY8DOlGwKwQ9jzYrZJwM6pwF1nXxN/wkA8pyV
y0SzO7IGdKm+dVYEtfTx7w1rT7kKO3kFdFKF79IjUvGrf0+F1mkVOaRfHyGbWRAq
Wkh26Fy3BQSZXCWn6/wPXBvWsvj4KWMzA4awNH3jMa0XavIqUv++ph1toNShtZuQ
vjK3T9x8b5LAyCa2Ez+B8l7oTQKV2533oW188zIXvEdwVibayaTyO6N/LrBtfU9g
GlIMYh/KEzn4EIN17/A46yIpQjetL5mM31sNbd3yOCxMOR77ZVmRmLKClXnhSNXj
zrtw790Cg40ByiuwfJlyVJ/fYyl9SfohJt8COrG73VdewEEBxcOR9PbUa2bCdNqm
fLre1vWoO3mJvQu0GQCisD2w3n3/KFf+8mPY7MMN+b71cEbdRPBit7qdrRrOPEKt
/ISIHvcF4R8zq6MjALCL8xzJtK8ACOHIexMAGjxR0LopqrxQzSyFhcnjAEiBMN/z
s9mcUmEll2Gl3j6kiKBuI5wjcOCroZzB5lt2EYw7vw8EZHWY4Fh8pJ8MrYvrTIA+
PJpRAWT8QMo6dPgwHbyolFFjr924z6hnDrY1nH777LWOol6kisDRfKdnpcesbuNB
aPc4xaMROmuPGtweiPvCeMb6XucEoQa6wFuP7HUDzWO37bQktdVEdY7rEO18UxkF
Q2dfiqkqbcryuoqrftBqcq487ZBtQ0MoFSr8ymtIGAjiEcLFEKl2QpWJVr4wljpw
GOO2AiZ4uYPCCxLTTOjFzdwMVm2Z+redscxfcmVa/kFwkVH1KXPdKi9HOltMgPnT
8OAh7w0yUM8b8uV+lTL+PuLkv3cwvUljzI7IxpPGi9DpI1G5uX5fvvO1OA5hXNjZ
MvcE4Lm1Um/AhnkHZCyCPPApphLC4wAWuBsOJlt6epiXYlddGjdyTgaR2DXRF7Cw
IomZdBHbCde6QjLNmouuCL8NwBSrWAVxnLfpEJc8qs7riNeccsY9j7OQOso2X0W9
EET1su7jkTDSkPRKqQRB+nv7pBUXDstIP7b7QuoK8xLz5CYfk6d4g7BgSaq91NRR
OzmLs68ZOprK+G/PuOXG3qF32OboBfOwWUaIG0r0zNV7M492pnZ5qOB6nL3Zlgo1
93S77KPYqQBFHjDr84nqIVgrwuspQuDDlYuFhdEoymL0Ic7b0swehA7hlbDtIlDw
sRq4bXFeNk254rxsXsxw1hcoo37k5WTHUBZSmLIJu5bjV4QQuH0qJMJL2HAtINCj
gbetdpovYsc7swQKf77UNmByTHcosao2wrMgG84LH4miqa5C/iXDw7DUir/xFdwM
eaiVh0rI75SywDOhsRBoDoZi/qmyXSMU8VIx/fZ1V4F2Me/v7OXpH5frU4u6Zr6u
BNty2CYD+WOnub906GGj5444leaEvtkmN/GZ0LRMlRLZTp7n4Ws594GiRjeZc+kS
RCd6kWnnpabcg7/4/JA9/wlJq6PYiNkv6HvWA4Jc/L28Bm9qbYogSYSynly3BnDx
wQxLWpnSxJOoTllpCf7/ArZUDm3t6lxyvEBkS+YYgVtlZ7bWNq2Oqd4tuNjzQnfr
9lN5hL/NZ+dfFZYotXta3M/D79jV4v+fK2UrBVFlsqQJddjvlry4Dm3c3nX2n99V
OI8Bsw3dngWr9b3S2+X0mXpxgPqRQC8EJCaVc98yNcyJmJMYEcxa3afnOwASavZd
ArDvqRhnkwaS8SvY7AJHFNtiWuva50cKpRI5Zdb/JwHrmPvfah7j3Qw6AQG1itJK
QdP5/tw2+arOnYXfYalXBC3bakFABYooQILWkvjvELWViwBzbu6jqM0RZaAYpjBt
BBTn2Zt8Ws/JwjeuD9pRHblZ78IwcicBrRhH+oJAiyaIM2je1u0xyDPd9lhx113y
FkSFY0ggmj9QoKhDWstV3cmxgtIXQmv58J8XXJi8c0ijnd3gFpgpPgniNCF/yGse
yitwMKzv4RVvG7OcxPGDyUs+V/sr1bjDENXEwqPOPYdph+TkLWvfz8nrD3ItAC4p
l8jV35xj/RMdncQJx6X7vlpgc1wXTVK1DncUXPj+XaMkt8o20iEmuHglGB7+wsBd
m1ueorSBnLPoQmOLceL9Y4NHF3ljn36IKqp1Ttb98Cxxn+MYytvOK0Gte9tIFEy8
n5MIBWzfEWLwiBNZ52XaNjPZ6LJbplf9Vd9s+D3728oB9yR8PVjRG8rZbn8yrpSJ
1U6OF8w0KoK/biSu6ZXnqDC7pKjVjTftWpBF2ot5XwFmoz3Ib7I7HTzAb80Qz6dv
+sm8v2+okrZ+yd+BONgvT0FLCCWR0P5x2hPzGoiZYvD6ZSGiOUSBEvLkjNF9RM/w
wqyqKmE+n8P8enFCHY6ag2pseGroH9C8+L4FBTYXqg1GBk/V7Xt1Urwi6ZbCiIUn
iBPr9u68DubTosIvFTiY+qmGkP3iTKeQJMhnWyjFw09SfLvOsm4StkfxpXDMEtmx
WQmcAjrqS48nX16trHVq6hrWvQ0gf+8a1Z2c4qL9rQx9UcALX9bqErO8e+cyBaYc
pt6lLVTWEz2ncMfnKTsXL2K3qc0mwhW1UrwxBN4b6eNTkyweYm3/sbQ82qIyF/cq
hucS2ZieVgpQbTX2fXl3sAtogSKe0t3bAyiDzDXXlqle6mjEMLw0Netc3rxPTW0o
Je7leQ7PIneQ8EGuYM3einnLJ52z5VPyzjlxVNq+2ljJmQnNaMH9qkrUKYFb6XxJ
v0G31F3qa4qNZKtwQQvNs8cveDSIaDBJ3PDhnOgOG6DONxzwE1VHE5f9T29T+inM
9Qw9L2hNjYeXjkZZpBMFCQw7qRCJaHOdr2TC6CT9hNO1qC5L3Fj6PrRinNW7jk/d
/6orXtwtDnpZx0EHS5wC8e7g+RkD4Qgj2x8OcbosP6qNeuKkvo7e67jIlHbAfbIo
eSFJDJhtzlGoGaYfOdepY3GVB6OQYcY+bP8jtyhlH9Sg5/lYWyTEn0hw53+LvbRu
AZtyo21yyovR5STDZSU3VUtKELLTDdBMy6b9L4egEX5EWZYwK4ANY01nsG2RxNgC
iTWjZRFEmso+NlrgzpQOwLSw5Vj0zsANgYcWu9SIu7RMlvsFRKN0ko7RrMvEXGZI
P5MwNUfGmNrWOOilkFLn+3YgF1h+TQlZtO0bJcY0iQkSrAHkCKiegmxG7T8Qu8ku
i0aClofI9sCbt1MwbUr8rPehScyraPjnwE6NjpQX2GJ/ps0wtxKzr+ipiwclnf25
MCYm24q/SmUwfpS7iEqlOqRaEGdieCV5zUIbvPRcco3N7GKZIF1SmhEFQfh4NKhl
gbU1e8U+KyxfpkGz+t7veisOJyKush/rODE9PGE7sQPA1I44lpQHrVvUGNDSBplj
DtlgdB2A8SeymWjbtBukhaZRGa9aHEQTvr/xDGgEwqvmxx5epf5gWkCw47XsMjjs
aEVGm9o6dACo0I1w9VmX2mwCgfl/dUdk/EP+3G44rEo1VqSpFpMPpDAh5tE8UiXG
nLetEa99K+DXfCJ1bxJ8aDmLRSmwemQAeDthuFkk63gEnfVWxIRrZTiecGAMR29/
uO2ERDziqxEkCK+PuIPYvXMWdvKyj/aEtQM1wL8hw2sQAYZ9iDy98jq6XaTpAOgs
caBLSZaj010mcmuqf93qjvpiIHpjIN7cxXRiBQTvf3H/Q+c29CSDzIusYpyPTxDy
T0gjfGp+CM6LyAiHJH1v1Yp/frBAU0kgQ6y3zbhxkZqe9eKSoqV2Mn2S7qAKQmpv
fYkR8vbXKIyVuXrryQtu/LU9+DIUuLIdKi6QDdIEyJXxTarM8W3rQpjMsgRT5bw8
OpY/0ya9Cy2SSN8kAWktDiC7A5VWTBAugB8HPZz9S68/xA0kyKhIK/mwy3bLz5Cr
+NprjFbXlIPuSSNZkdMjaE5RxmCC7ciwq4aojBPHxizkdJ96G00tUH/zYSYmg/6w
nAA/m8ZOYpEaaN5kMMU9k/tOgBcrE/f9CMcomZej89EAkqhbN1FWfHWMQXdpdgqN
alqOydVI1f0+GvYXVwFWPA66Ymv9S81MtqwmkM8/Hkyr362bj0FlkevqR9Xd10IS
ikbI18BTJmRGB8pJx+XyPVrnDwQAD+L+i+SVB1h1d0vqAmFQePKFzCGZ8O8F4yJD
+eeQqgdO7tjZSwP29v+tR/7IINGIuP+u//iXE+5VUflcQvia6CLuVqN5hG3LBsis
VlfqJrSuZuxFvcdUtxS7WonsVe7FqYLy/Z3FvIGzlkIl9zBgx5Xq0scgHjPPbbL6
NvNEE97vB1H6dOO5Vu1UBNi319wIcilqdqfsSrQS0Yk43ZFZiTmbtDq9lWxPy54A
qbBdx75te6pH6uxNzOliPUI29clUKQooPoE5aR/XwrBvxc4sIos/sxSUo6omh2YT
8j+Rv8/W+blTeq147VCdw/UwCNTPGrdSo21W8JxtSy0qpxDAuBeKT6r+k1RJrPS6
LSp6mDtOkNL3S4Re30rtRBziWKjUAYttj31MM5CHUyq/PETxCTNtlRZ8659hY6N3
qXoiTAiB57gINCjLYKIdW9newxtegq47o4z+WWNzkCDYZG7JEkMee35aqL5mWfV1
3tjwmdaF4FuD2me2Bdjk14FuoBb/SzwydBBXbC+S1jaxKllvVbAH7DFuKiDdE0gb
LuQ+jPgkf+Qcy65dOg/1bmwcBZJjWM6xWxLqkYB2AoY33yG4OOzrM/HD6bzFkCbL
dM4gFzmwSfKRyb9sBY10xgImQZelAhUdOH67ePubDgNZChD/ALwdjNfPYK/dChZt
jj8JHzszi8iTfcyaYgKFa17o5rkJ8lfBpiPJcr/yMjtPzrbP0/KqSFOHI3qttxb8
/PmLV27r5hSj3IRWKTj3kT92U1jwUKSkyomPhH/mHmDBwk1xU5HJC/ybfsbhpVSR
FIFCo0geSbaRYZu/ZM31L6A7M6CQZQIG56ooJTOOYfe6gMXJr3AjkMaiorqZMvek
8cSD28Ui2XQUb/BsM5qmk5kygPS6rJPeGop/K3TM/qLwLOcNb4Awbn0DNE9o49Lt
6kJWQg+cS/cwJYLQayJqcng/glPlYEQPz+m8JCo849ev73xifBJ4TCckeemAOvSJ
pluOCC2scS/bXuLlNYgS5ixUl2kO0fvgDn9StFjq6AZPODcCpuAM4+f8VURLRq50
Ef3zH1BE/oTkTl1xiNui+S12Ohzim+sF6x11/b1BrEKF1GuyQJS+AGTJZW9KcQm6
ejOQJLkAv8LZUmkJVwIS/2fjc0f8lgG6rSLTKjn0ZJesH8U9YxPACSrIfx2hlAxp
jAl6X1ORfVFgvAUXreUNnl2fIT0uQaWijgtfryKGGSXspZETuMy/6Yasc83clzNa
U29rcv23VTrL5TxSpqTWP1r0WaTyqTzsjXRCo/JZm9E8we7y9CN9dRaCCdcZsmSJ
6mRD3IqWwMnTRUi22/PXCl1S2Uv+oDKLfb4BVLsxqmg+NBhqbK4GB+cikZohHXZT
jCbOI+Cw5wSLIUMfuFDVDDZo9oz5+8RKmjaMDMxeESx47enGntjEv5VP/+FeoYLg
iPaJBBpNqRvr1YTC6WwOXJRqwbyzYTJ4aekSdER4bIP8W/tfFsseZ5BZdQ15EVFh
MXeutQlYYk6WWhR6su2rO3Uvz9ekBxnHcrL6WlmmgNIaw7CXfGJbtqVZn4hnCEoI
Rb1zsWgrcS2e61GjPjSN6+1kxCDvpTlTpZa2qD4xlCuibil2UE7uOppEf1n6n144
eiLvckNEj7YGwYIvr64X61GUy9BvtiJRWhsiDV3i6izX6aJdN7U9uZsGYGkZXcJL
eq+O0dPfGfdgBkNM1FCRhCCD9FWsIlUjW8FTKhuRCtOyWFavyNARhvpSq56BTEdM
k4KIxD7KHva1vyc8wDU9E54tzaqzKerdNAyNoGUKgnTpS48n3DrEAHHmrYpm2a9S
/HMoF0YgiDDP9nqDw1ZUM40AW3YltMbBHromIpXhynBc+n1PYlbL5xLHXW+uDdzo
uAC1FP0X9as8ThQEtxFdFnHNSyskkNbmGUGCkA8EJglz8IJFTPHPcPR/nskZ5NpI
iS7helJQ6hESlVEacJOiV4oS6478LXliOWWkN+M+yPUcnIFYtnmEOmN0PvdidMKe
JTuaxmtQsA4wS3EwMZEkksrmiHPWMzSdX6gmInZBY4s/yhp7jGjpcPmPEyZkdQNB
VDCNV27fLqgYv/V6hEG3CzDBoobC0tKBLLwq2eeZcY6q+iMANFHAC2Bdrs7abWau
tbP9o4OUfOCeyJkXr/3t2147uTsWgK4k6E9P6QvQPE9K5JoPVUqk1MRSoCgY7hhU
++NAAsGbqH+dn+zEDZJK5x0rGKwZHLGSyRLV6m46/Xndn8/IvGPvTeSfpHhKb9nV
Wu62Sw2oYC04lwU0Ywcqi6BKcKvcqxdDM59Pskv49E0WzBatb52E64b9Aqglm/s4
B8ncngx3Yi6isvFTCQ52XXsoxJuNsPEufYzcuCRFXMst3jYFA8w9J2R0sWyaet8C
KVkd2Wvhxt21vOKAFyYfNNCIfFMGWtNvCUBBG+46CwvKZ3saJtO2zZpt5s01x9XC
yG8Vxwor7qY8CHCC5x1h7Hwg3i+nk9XTOGyiU6+x6kNjDSV8CYbNcsgtAlKiMrhX
+n3FHihdhFt383Qdc6d46m3W23c6EiFmmOPTv88PnZGb2NSdZesUm4L3OETKDuwB
zEH7yVyk5HOWkXDsh1S9Hbr79Dxo8+jkM87jNFtHv6tAj4J5UwCNfmI3rXPhcGfo
p43vT7GGW3PM6JDjFJfh8EL0QldXF5qoaWRMNeRdVtlCx4C0elHMX4jCk//+9hIW
ikd8P95BXmB14wxfq7G1tkQehA/Pt/fkRHPiN4PD0NFsy9b3Ap+ZZdeLcBzjR4Fg
pJ/eqbQntHpmZWsshfcPxPD9Z/5CvNoIA9D5K/0Qq6d3HfIrAP2f3twGlC7r3687
ALD942EPxfMB8FVWKcX81CAKvqRCzVTLATOJpXM4HZgodXF+98lV9yRV76cNoNXd
OiZ7oIUfpWapBetoT/o74i3+nq0/C1XaEXmgjQrk7s8LmkJ/K+7umO9Ij7k7vdCV
Inrdrhg4trBDXzlWYiXCJStWF6yMH3Z+/zoVcR4mbolGaonpXg52o7n3Bgcl2hMW
xP/L+zuRNlJJx8HdB2BLZoZ5og9NtX7LfDLv0C3mRKKYoZcaqJ00UOoPvas3RbzO
qpqhHR/vJjaHpmqyB7kl1hoQt6BRMuh3Z1lIOMtSgsCtdGvKO5Jz43QHHIxK9Ips
9dWsNF6O+i5H37v+Eac77e6gHTIa03CXNhbPPjQIRAS45eZfv2zqt7YS/PdOK6yX
ITMwtnN/9IO5DuWR3fOUZb/PNjx1/httJiIDRwP3u3Cbu9IKXyZTuMWAVPmpam1V
A/E8FsPl7A+XoGDfZ6PRinMj+2bWWD0wIAg5UZFXQPQ6RBZdE05RlGlEWpSgs6i4
J/YrqK2ZFpIBIIDKgu2Cjtx6WXLtcwkDluXxEwOT5J7P3vDGGhlVMShNEt+o/I2o
xpWafezSociW6YJDmiHG/LnDaEhfTJq9oF9EVyQCcGSPxlxX+HY+A5VuhocLD7nU
CeKW4v4xjisZU3PKavfBIf21rUXlmSSsyxBSoTqR2on1uIu7Fq4UrAe7bXLvF+Yb
/L1fxSfEcWIeNmIoLfWmQ/LLKicao6qkNoolpHV+yXh8MlVz4aTFL6fZvd41r7jV
5SfVEBgNeS3A+AX+015a/heVYGbaf1eNcv75IR5ilbmiVobhYPiDdZIXUDTxyqzu
EtF2JgnOmQE2EcKWucSYd/ZTzf1ugSAggfP4ocrPtvGJyCCZGZYEdYp+EU5h2sPV
ZOqJmau+6aRz7tJkLNWH5Ba1l/AqMlyszm4f6VSG2dwyGZBpE/xo951bOX5xPMag
1kqSvtnJVNluG2Vh+BUjaFH2lY8SziW+PuKH6SO+IJY9nJuJqaqMnb1OaJu/iZ6N
omuud/d+XwSPyNXXPl0WRWIyVc6Eo5fclV88LEZU8257CVmhczWx/BW+h/miOnSf
rF30LdW38Oa+NoXBGhJv3qXU909koVOsMdFWufI6DOPn+welNJe7/iSkwGiRpv4K
/O4rL81U3yVYSMAxKYZI6bfqlb6kflwH+OV/g2xFvNMc0lmGFzzkrYRqaJDi+Obo
wcBZWYjD/nCBHvuiyQ00rVQz7azR300FzODHISCJcnk1sPiLFMx4QCoCjWKWpP2j
ta9zSqWOV4O9Q24Vtle0GU19aCv3l8s2PwxYVxA+DGMTtaFydDm1fB4SNPfRCywX
5vuCoqTqLIk1w7VWkCEMZNATQ22Ui/yT8y1VY0AoAdsVEJH7K1nPHsuPOnLlhlkf
Jdr3q8ToSBE8LBsPaa8OmXYmHeQLggRbOqQMUTNg4NnIc1AGj0zugSWcH5DrsENr
vTLQWmxKsWhdzSC4c4hXqN8ZKCbTi5kVlzEJ7eAxCIGz4GIOJrleQr/gNb+ZUPHT
wESRtnk2LcANhLk8I0jcnbqjkqsuK4I7yoGBSCAhCHLsfjekIxVVOdsJBTQFzk/9
d+4D9k4hY48mlXxBjA4+gzMwmNXQbDN7u6ZPRirsvH5Me2DUsQyenHf3og5CgKn+
4JHAU+waIj7MvSRAQdQiJmU8j7wZadXRxbspvD5BiKo5VaJyPoei6OCg+UIQN4aK
ArBaN8yKYfRbEbjvYv/b+na2dim/EbAteH/B3s2+NtGhFuDA+dmROCSmSm2rWgIe
n643+qnF4EgBT9d81ejDtG1oNVdoHwJXUq+W2GhigpQyA41IiiYQLBnYJIdeA6dP
Poff0e2/K5TmZcnZj12fF0Co0OeReLyJDEutWdVn7DABiXHKsNFdKQlPTR/d1FjQ
Uw+iIig6F/l/HfFO8041RZF5F5Ibh4eRC7wySM161jKotugED0Ccn/SpmE+9zN7X
5Btw+/RYwawzXcFjxiQNjk566AHAe9QJzupJ0rdUoenXvbCyTFJHjmQ+xNSWpTOp
h5L/qpaJKFR2RbYn3Aaw6et0ZRqMcfJ/fIdz1YqVkjsIi0/b4ISMRBkf6SeDtdv5
J0J5ly6yqSs3KJrKtz1YlT6YspQf02WqEyZg5FizXR3x0w9u5K6UPfRX8dyzk3SA
qerFttnwjRaULkyyjvmwbXky4jCLlZeQLrUh8T7uEUF7sEwXSVX9LYsodrRYZ9yo
NQf6Dm0JP2WmvtasS8BjQ/83DmMfTdM4krnRVsRcUonO1MQuiyacMSLATilkYUdN
SvJn9ewdUr9v8YHXG0HfjW34a0D3USfU/lqYdJNR9DahXt43axDat6hW2pdWYtNq
g42Utv1d/eKjs4kGfEtqJgI7FVkD5LRkl6oTC9sMyOcdpvq9DqRdYKj9KjGPERmR
OmyUY2UV74uF69212IhNWGaA/UMjKpTWm62v+UaEBFzHJbK8dMTQ2A5tRAg6vmfp
GEbW7ht565gtV+ZcFGBYbqbQ+hQR2nYhuYCYExx7xl3BhKEtp53f/bffHrEhdbf/
mU7GE1MaS4FhcjpH6Lw1zliBpGPH7Bcuk8fS8iUv8PQfoTI4iFrpqR5SNDCRbf4m
S/B/86DmAocFOb/9a1hmAU1sFvZ8so7vGuGGaJN1QpFU4cwaJFzXgwiBWa9rjqMb
ndMGv3qW0/V827jSJjbNgRkJUMnDtaxS1HEi8nz6EHuTYQB8XytaDynOsbgMKP8z
AbVGQacalUDZHUuR8Ft7GpQWxuky29VZKvq7r8PYOwgM6DYw/xUG432xP1yi1z1S
vhQ2jxysa3p7FLOGG8lTmXUzIaaefzNKuoCuyewd/HQJ6GJJ+SPZhjT9fiAGp2LP
sLCKFB5bXoxumoYGqJvhgLPNkO2w8mKbI7VnimGS+frIySDnjOVhTpTi9vnY2LZX
puu0wh8fEzGcDIsbCcMKUrJVxnl84nSWIuwHyAU18IeTpItsUIPiR5gxohGI23Dq
N2kx/DsyjMRgwgQXhpfpC8arM2GhciileKASjNJ3RKw/Sh4k7gXuujWHnu15YaY4
Pgp6Kw8feP7bnulJV6xQfC8/dNkq09E5YpkYbtLagWZCh0kpKvuy/1G57UeW/B2V
mjH88UVYJ79HGzpuE0Vub82+GkjTXftGzucym0BfXmcwXuET/UC2xE/fjPAhfs2a
VBSxCdPWutm2fQjFbot933ov4MN18/9F7nzSUE1kDISlCk1Qjk6oJ+BlMMH+wyzq
bRCyg1lOms62mYPoekktP9o0+Y4qB0Yn6niRMnS/7RkcbhDN2a+fEZeyApLpMG7V
2vJkRxHxuvAG/+C3JjljYICR4RdTQ/pMSd9WFNE3f9bR25KvqqFjzOxICPC0q58u
S4wfU8r8RVa1gnhyKXgOam8mcSASUmJNQxg8txZnAiG0iCpV39/GRuPT+UJgq/XH
hReZhroIo2ozXq9nRR6DyR57OFhL93Jz37MrzXbFdNcHx+6IawFClChIdK8MZ9ql
B8ZrKn2XTniJy4KQ1DA5qjFdgKW07r9CkZr9WeFv8dMeVaIPrnKqmZdUjvEikxsk
YL8Vo+2zZD/cYHxAoolJ8gry/QpB9GwY2qQ4o+jfKDs4bu9Tcx1DAuDCdBIeG0rY
+oql6h/aLjfIID4JVAxyV0vFGC94mTgTcyyQeiN7vKMkt5Szm13qQ9WO6IT3uBRK
E7AmbIK4VNRCOJgxAoGAQI6WhtBwRL3MrfCs262kRvl3WMroZK0Q3YjzBbLXiCd4
5ZoeF0qPdeSNbTndinpYH3uaCxlVOGYzYJ9PnH5Hv0i/c0A7AdThFwGD4s6k3Stv
Lm+aaZ/wpiBXX5/DwOjBCSxzmj8USIYA48qMrde/p0rO16pClNb+dScIKphV4V+0
SINsN8Ur+cwQWNtMcZC/aXdWd3St37IsMlhz9QC0mmqjvgBBs6Q855eJOkAT/UMQ
M2YC5Bc2MoFuEr7NjIAXjdiiuB/ViETWViYHXc577TmgQGQN3hkc/cmGfFQbXNOb
EdnGCcI25Pnd/QEK/YAkZWqXRA+gwP8I5YWhqAKcV6lgp61MHlqzy5Hc74+qTUJY
KNvYhMyKBuwmkzpPt6P/akgVqZ/fZNbQz/8EFYn6Y4b+Kv1Bbfi25gE8H7KomCcq
EA0Pep6VccmdPwjoXZ/aabFoD5rky41wnzKeJDxnzerRQuq5qEwemWKsHzDZzove
PiadnmYCS+qw2zyoW59A83ATw+rnZBnsYvz0LoQWnRp9uPy7uHCVEhZVl85BPPGp
vZ/L0/jf9zKF7vHaWm2/NOGCXT9tDHIl2oFtJ+/X/53UeyuxeigcbiRh1Sw/X5zS
2NUFWypEI0MgH00DzLobrdeCHbQ9DaCAzwlF5jXQqCFLzuXJylpwoEEjelvxNlqA
2zEfzZkPzHIn0YcGF6JhzqGESbnE0ky8N2y9fEfDFmaFDak9/9gamX4OQxaWp1CQ
YqKRB7Ut0mI0ZfnfmQfllwO8KAydtlYO39/prZ0UpmyoYpvnkwvFrjpuEDD15mKU
XZ4CduSOrpGNtEMOEAiWwbNg0CNXj8JDJTp0sJz8ft19JzGyua9jeaR66cAOgPH9
eZ7W1O0eI2jLoyLClnWUHK+oa0arOL6HqOSGiWao/E2b0vOVmvALEIWFKgejHICT
Ufo6PK01vM87PQ7Uy7l8w4WBqyY4HE50TlzuBCexulkBKrK7Df9N2vmqmhJQb1eD
qcK8T9CYtsco7Bj5FnrO+53aAB9DAgULSNIyW/i0kyICUgtrtcrkcJ9fQKr3y16G
rgDdhERZGYoaN6hrkmlnlcC47kDvOtXafiwqRmpSYfrbvx3iJn3hz1XTsgO2/rj3
81s3Yf4mpq/NIKNP38MbJbXbswKq3i0bQPK8TjSxfHlSktCcSUKnKQ+zp/pa0VM2
SxIsjTE18ZSoiFJjTZxpAiEjvcEdTsQ0lwZkh0ZxZXcYwklrXuGfrz6ugB2O3tvR
4HaIm1sEnwtkoO5wCufRO9bmOmWlFdAE2Q4ZryxuoqQ8luLtvpi9QXTTJN0Oh/Jc
+d3FV3IlJVioG9Ap9GvTEYlKbiL4bUJTCVqAVjVD3sLwPmrdSQS7TyjIxza7bT/Z
PdddqlLe1QM4igpBsNgx3NbLYPTV2x0hhEIU6jfmnVMzqbFGQUskM6Zk1x0ekZNL
dkKDzThYBMMN1b42fDv5tDTZRSZl6nQA709UAY5I2lltmVj8zKVBjRG1v7e7EMQ7
xrjqZM8GrT9xTczfJN2fT8QevTgZaJtGjd6o5WmiShKsOkb1ZPPy8MCN7OW0FK1M
BL7r9+pDO9FFqAaRwHvLvMvbs/maSwlfneb4Z2Bgf70S+2oFcjEkNcZv6Kvp+BH7
HhQEUsgSxCpNF5MIGTy4dkkwk6X5qeF9aHkopZVHeMd/pkjFzJ/ILymGh5bnXF6V
dIMRPhcr5O+HvoKSCfRGnQ8BDqgPch7wqmbr8VNjVmgbkk2/uvearPZORzTd9ItE
a/phig5kaSupbjEHsB+bjOZmaYfPzBq/a6XAnxCV0mZsdnHslaoVC7nP/x0qMKuS
7pvLV+qXKXW7oTbGmK+HPkttBv8Mh4eP9v15DH0ChjpXwoa83ISDTtJ+oSGqSbgM
wyc1wpB8ApCAZjbIx9EzwQJ1BrbZN8pmSN65QvLyIAUoaK/SfPo8tGKNGeCVIs5Q
Z2S9bFsnw4DUXiHnBYZA1K9U3pkBaRFuicIKNedc2dF1j5/i5+HruWn1agS2CgZZ
2hYHogZaT5+myKEnV1IbH0dVlqjoU9ZDXQT0tvHjZllAU61UKdoIs2uo8pQk39AU
/7OQJDxcHwvnEUNn/WHE71iyLBHSgG8UxeYbkHPYnDARcQEbmVFxVLkD2yfIJCjL
H93X1TOf2vW2fiAlXf6o44fFLnyo0/biXLvqN2eb2hckMYvdh1vhH+htBGEQ6E//
/zG+dm5IAeTI5xX+2FkwPUIon7PL3HToiDa6JJDwcabAXNbZ3aRmnx46vKrDs6rr
ANVI3tiYEXfKFOlKFyQNspFVrq8G3xM1co/dKhbfhe0fzEVRBjj6A9Zi0gFIAQuo
pHigm8e+LksRTZe+dReB8GF6xOY9PzjjpNubtDWwL5dTbKwtQrL3Y9/GOQw71hHU
TzNjgZnKEf72xRZUO2F+xYBDj2F/oqNqSp8rFSrSAR7V9I/JpPwEIYu06Sf/G7P6
Cr5iDXfktfVuOIvKbBPkIf9JQvelWuuQBpOikH6oLX2lVgOiNujXLWPzI9Sv0WMd
mRN94wQ7rQYbHILEkeJl0ZzbMI+3D4eUb1BA4JgUYdPmg5ZM1ABZFiWXl3Kx+Qze
LlVh40yddELj925I5Yl1mRUmbyRi4lTEYACE/puYxjdQ9U9/z/vYns2XNptSOHpR
Jxs3CGlXx0fRpGDDw2P8UL+hn+qM/HOi5M0XlnOD8vjjOO4D5ZcxvqEb89c86LGQ
r4TaCb+sIZZUa7vgXn5LL2sdQp/kuEdX1WdGs7m+5A874dm99Us+69okzI5ndQXZ
yo73RdZDd0hgS/jZm/tmn4geE6Ua008faAWIlC6vFcJbI5N47dScxFMaMTM6EjF9
iBndsdISujSQyR3ZQrj4uT4BdOVgvwbFpvp7unDjFVXECUNHd2JnMe2aH74oXIfA
5dk6+jh56eCNB0Y4zc7RTAvBi/Xar7F8YK50y0yKR/3/5U6lpiBImAikjP4z78D2
glSBIQ4RYvFBn5UWVxzcmtQdtfC2uMaPo+NEfVnuKm4WLu4TdMDH8PblIExeUkZl
vxEk51UcPP86yzKz0dxrOawXoszqzJSUDl5UZmikaYrxyY18PCE4Jamh6uGD8FOC
Tld+t6eqZECWukSqxaFEILB3A9e3cxuiuXxm5kLcSRhhE0dtkcGn7vKfXEiQylgi
rMBrd5pRy1EoXQN+3uOeD3cSOpLpB1Znqc9L1AaK5icUAAcomMJl8FF6gzJZdzGm
kfI32GK2rikd5OC778h1q2t2qrU3LocOrvz0WN1MZP9Vbk8gsJr0Fz+DITUakBjx
9MqXv9WtD5ezyoeIPzVi23vamMhKWsjbX02DOkNnzX0lxJmWWD9dVWsl+W+JEH4+
J/1Hqj3VKj+edZlFwm2vP7xX3PeYKvlRin3IgXQLw/bYH0niseVCR79sZoaISGUU
tM1avTfFogeir8LSVuZfxcqrKCescsW/phtdjS8OuZ+XLhAmpH5oTd/gvh8uL365
gwLEB4WMCOZ8+WxfKAqastsN4x21JSHhvKhbnCiK7NUtmxuvCMpIYLuACxkGQJIg
JoaHxljcsPk9H7soE9iO8hZ4hQgvJDcUmojSmQk8y/PjkYAgjNZd8mRA3TMH5N2T
14+eaLq71jplxMZQHyWPtcSmZ1YJPqi/sQstuH+BKmFQS42gXBFMpYI1cbGnDIEM
GJgfyb2XgoViFks1oVVUBh9ntCkKWLBwtmH89z72fG419NXjaql9enE2srVPOsM1
CSw2zNd9AHVhCEfk8rVP4fA4ogV12TXL4GSNgSsuGc51bjmSQyXyNQ6mbyaNJ+Fj
Tf6l6Gt+lkbY/YWqpCRDXIkZlglQWFDtG5l7CODhgZW0pAbCZGl+r9bPo/ht0FC1
fUecdBNx8AOMmXVhqWssBOaxr2VZcPHr1NOUyHON5HXjXXEU2/Oxbg7otB1XxOYr
lmoZ4z36TQ8te0swPwaYHB7WzeUiAZ4QVyiQpU1zSaIVu1qRNd0X2AaKdnkJn3Zl
pcRjtDB8t5YDBqmDz6TP2XWdrbrDqHH7fbXyEi5l4HYBgIo3RzbWHc7eksZrMcAp
tskim40lLFGWqPO1EZlk2kW4k07wHOK4OpbbW9rDYkkN0TxhiLmuYiX596H+1aJF
IjGN94nV8l3zzMZxHNrnznzqupSo5jXX8f4kLA9cIJ28EPV9MbECXl8I0nHTzgjH
9vx4xS74gGAHxL2YSkg0DBeFogwlTeROeYsVwTQOIh9LGWSzvzNVrWr5ix5ig95w
JUd2cgmLNeUHgNtcKqUMEAvpqs9H7rREaLaxFM39ei9RjNmXp3e+ylfFJNXcnpLq
G6S3qgbcShByeFOCdy1eaYQ45iLHq1RUm/NB8v9AyD0NhFjgGMV8qFfh7/NnmF+S
guGIrJV6TbGSc6dI1woA/uYw+QmQ0pws9y26eaB/0kZc6PUz66KvONgibSMvywXk
bGDbnUOEyK8zA2nJq53h/qSS33c7UWHzb/oLa7e+Yqd3pj1wN0susRpUbD9K7LJV
spq+3cLo+JpxHX8pDVinjTenEQdIFaRaY4HRY4d+vOef8OvuecZiVNNKrAYl3xtI
ifxdcv8ebhFgeuDZ5rhr1nvrzHrQdbp29O1sxzROASxxyVKfSlp4FbdCngIZrJOg
R7ru42KBd5YvDjw0btR/Z/6vDwXJZObjwJ2LhqrNoXtJss5ZMLdeLn8y0Jd7SYt+
LjeCrxTA0TCTDCp+l9Jio+h5oYYz/aBUlB4Qvj+Lcse362D8j4VPwXfljuLvNOnA
+TeCsVzQNqa6nbI9Ck5pFHi7LDCQEe6b46TtnIinuFBmdMeonyPECZskkDtRP2K3
eYGZCRwkIxRT9RPfrm5HdVJdmmzlmFILFnWNnZLKR1u6yMTES48vfuTRBZItpiDn
Np8WjVFQudK59qcJ3wb2xRmeImiqzEP6X6JnNyGi41HtN5rPWOHiLzuFFhhSve8q
NzfzAzlTMvKgW1nfHHbv8JEua9huUpztYnBqRtLPftFwohwguztmSXE6NCWG994H
8HCtzZqEGBzLHy9KfV8PJ2olT6IxAar7qv91PuI7TiyluJ1MI8YPkypftMKVCh9S
7FDV0J9oy0KjcOS7w1IRg8l7g28SpYPThh8ZmQdgzbloYkVnse/kcRe9CDGDdiJ7
P0Jmyiqb5iYRPyUT8omjIKABBkhJhjbjBRVukY8FD/iydiXGw0oz9Nnisu9p3f+y
oUn/BayeL3jFrHORB/Bkv87MjDytElkXx+Uchr0DgpZXIz/RihRWAbFswDSohfOU
0sHKq5Jg8xDNmdL0F/etYJFYksyCPMnOFwuwijdZz7tTleyoFtbum1cen2EwaSJn
kKEbCyW3WeiIFxbSjrJ8CQin8PzBsQJo3ozLuGTfv2rr04Dka0eTj1X6LefElVst
L3Zj18CSeqyD4OgEjEX7RqK26XisC6Kl+TagZ31wWxaN9On7q6Qs1HvELM7ezvfh
Auko53MS/fw4j5EuDFXuC9wNz83KgXtRDjd2WXX4RztvVNdhG0/KdEWyptrVDsqs
E/tCZuWMYi57anK9UzTAf9akxMaNxIXKiqOugyK33aTTXIsovwhVnPMwKwMiwt27
Q9rIl1d0uxP5L1UAB7qh5DhH8LTUXiGy9pcPzScz363mrJeo/ejR69f++gvIK9dg
KZB+3Em+Zz6lUja7kfC8beEqpzDHA0gUwG+S2oQWkzvkAdFRdJbDxi5rMHXGis5R
8rIhQy9lXkSKLzWhEM3eqfFB/1/LlJe59jXQLSfq1GAWPdT6hzRInP22E0AdMB96
oXriWabnl4I/pGgruGwdIYyoIXbayCO4kxUH6N2SV4hpOnd7/265yLpGIn3AkXbH
pbLTKFWWg7HOCVR4SuhgAconKRuWF/YjDORsW4bejIm0Nm20F2WS4XwEpJPfaokg
CotTQyEEiKBTxVaTLr+LPzm36SONw4RU1+9ZJIM1IiIjJRU3yHIjgfyAvO668Iqs
98QpVkSHO3luK9Md37lThgEw1rF0ycuqyhju0RLHX91BHmaWxmCHJfvd7Q+Xt4Yg
10K5fWhJkE83JSmE0X5x4TC+BK1J+SNwP9XuancsmjObnmkWGu7qF0PEReJnbM8D
l5pBMQ1gH1fW2wl25NW9grg1PhopelkzXhco9uUL+NNWbcp1uIntUZnKauaT9Qb1
wnmvBE+tNdqL0Q9up2FkoCXqjj/43wkmJcO78/8VKa+5+yf1f/xB0fZ787KsB4M6
qvYe516mN40BO9SmFhqtgbEpA2Rs6xbJ5gElo8sR48iK43kQGjCxVxQdNs4Gtm53
4Ks2zy5bRwhucJ6AiA3q20OCmD5kCQpDgs10X3T3+vh+cvtFl9jSNh65Tt1MIBgk
EePnjlRB3N32SKWj2q+jnZ7P1SxmPblZTmUNUsR6FCjpYjAjwMXbasSF92dnsL0+
pQCdnM0713rLZzpBAesM5k90zTBkVMWYi44vCRp0qIt3hZnFIOya7KJAKyR/hHWp
GlF7evdQX05WjwtyLrnUx7VrLdd+6dl1qA78SdA+U6fxkfZTi81c4e8+GoJtCfNx
XCm4jEfTptw5dGicAL9F4VHzk/T7S1pZ1eWWTKSnGamJGjO/g+4p7X5sZC+Pa0Qo
Nv6FRtD3HbskiyZKopUM9EcerDpwjXJLUVnOAKl2leKcPXbmj8zvlL0o2vuGlirW
9jVaneAj6WumQR+XSA4Iag==
`pragma protect end_protected
