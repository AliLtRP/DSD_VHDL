// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
suUOsuNW9+4DSWFA+SdbYv75SN2z/lqzFlBCpQ7x60TPjR9DTZ1/Wy3yLC7m1+Ik9df46iQbqNb6
l5g5BW5BINdlYSP7TtoxATykhjK1jGUs29XwoFu1EuPjc8Ictj20nc5uBf2OQ1LrQ5V4+q4wi2xk
yJQbvuRu89iVeO0exHYSGqdC81L5ImmpsDa9UbYFnlbChwm665+eTGxK1j8yDfW+F2sGon6tgw7J
k0skBwr/TnTXlcHhJ2lB0JRQNfCryWiuUCaqwwDjS3psPB1zyRgDsfusdLnnhBY2sXTvCjZjrDp8
hnzf+DY7ksT2iAaGKZeNI/PnoB9dHQM72op4dw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
4VJq8BspKxsS9jtFTHGAu/7UaKggMYpm604+VrFb48SWPXO1r7V3Mcp9T02xgpVhnI9bTG0fo8AS
sWJJxFSoz+AlaCR4kx5DA8lbvIBzI0iaMzMuC0jTlMn8N1biy+t/HAag/7dbGrHj6L3rMaewAdVD
fiWWjaAfXeF5eMG/rbfJGIqLuWsKbYVut2gkQpTY010JV4d1x4Cs57nd8vfRaVHn07zz+Ik9nGjX
66D6qBlqZ7m/z70YhT36Gtt8vodX9/qy8zIbi2FidAaBPA8PiOfRvdVQ0s4zbSwxaZb+ajWZppjy
pXeaEezsJtQgn2Xj0A55G28txPYW80dmVmePPvvzuekZZD4p5Y6pZ3Ejb9dRfernB5T15WAqdo3S
4WFH4hZj1tC/7rQV6rvT1BNiYXMrQ/KpPl6wYybXum87bVrWwUd64Id4Vpdw9lj0pnUCOo7n7rJr
vOVsROStFZ9aRVF7Zs4+Q/jUJaqbQkyCzxz1PVj2bQd3db+typAF5mJw2qnDgx3T5BwKR0Ao2+ml
oJ58SdxEVmvPfP2ogvEjHLIO2FXWuSDqMnmbpugLV99rMod7QSDXOlb5DqUrfAMcA6Jdn903LEsx
VxIyif+UqGmEAlu/cal/t9dTc6RU7my653SHvNIJL7tvcacvFodXAjjAAlJp1cvNCiV2YhNk4dwl
EIGkqxuB3/sqcYG27xljuDkwfaNt/6yFImDf79gcKw8DIKnatmx83g7eqIebQTGYFIEfmz4nBzoz
YuJQXvQBc6XlO1nnS7j4P3g4a/tcRKRCjjVBJQkNA9bgPJSRtEuemoOefZVK3rWD4FJk1028qWo7
BKzTbqo8TtUzGO2OAL78OsX/GR4NLYy8+kJa6ddkhZfTxqgXN3/SgmJaBHQ/om+++lj4r+2r2Kiy
cygRfPLLW2NP1Z2usL6gMRailVR+pihyfj0I7tLruiNROoYMt5CpMkhblqSrAd0oAls/OWbWrshF
Pl06jlIKGAxTkxLYZX0dP4Yde449nE8VD+2uAA4mC/3zwXtBjIuIkVt57865B5nYSqa34mZWlnwk
gO3HqvwTXywgD19Kv3ZOwLA50uvZFtStxGhJzVIhuf5isunNY+YPObQ7hn7IFNCa9FBkreGZfle8
jC9I/55vwTQGVfxu+l8qGNXgRRRN6aGAE29K/E15Q/sxj0boSWqW/E5ENeiM38Q8mNna9t+2rDBn
SW4x5IgJ5ArLhpW+hvZeZE6yLhPzUCjwAxMuYhGTz4tDfs6RwsxJ0/pBzMy8ymOZp7SmIgRfWE3o
4sOzEVGSsMBcyViZ+U02x7dTeyNtkDTHYLtmevfqOmFnqBS1EJJPNfYM3dLhskbi5WkMO5A1+hpe
J41kwkq1XMyuWWjLZbdoUYJTwIl+uW/glGCcSk1UyT3v6/KWIS+z4vl6mb//iG+V3IVjpmzTDlOq
staGwBlAtsJRLVogYOu41LaG6a7fs2ngTwle+bOKHFXrwwpYWOwtykQD9fg2Crgl3uSYCQ5bNDfG
NjctuIGp7ko9hTNB2APakJb1q5EXJygHJGL8wa1H2vsIaJDjNaf5w46QYn23Z5cukA5Q2Nz3cs8w
iTC2kt5CwcuoeO1lX584OjCDCOXUfnM+p+6chUUYSVVNK2QC2hObCNvAdfO+15EzxBI0bhd1a1b9
WCFFKP0FBcYpiJgL79FriqaZdW+bYt8WUkn87Q7QJ5cJ5nF0TtX2xnnGPAOBNxeZ9FmZMUFDbg16
MOL2jVcxpGXduJpUyOuZXXzmnQj7UiVXHriGbkMLA56svsoy323bPkmkkQJaFEL+XU+B7qSNbRUe
EuNYznP3F6hQ1yhELCLKq9F6VKCKbamSUIkLIK6iM90+k05Y/kzWEqoMBpn7Dk61WeqnUXIQLAzU
EP51RD6XMoXKR0mJ5K3X33vaBajcEN1f7qWF2D2EfzrbC57eNJsPJygd9kNU438RK8X6Ptr8H8fA
XrDoV2C11NwZFzFFwik93wQfOzbAFdd3hth8zlFjqBQQ+0R84+st9kVKD+HuIohBSpVF1j/PLgOj
8SmbvIKR0sfe47gLU/yYw8D0eI/eCe+BmeWD4nnNImq24cZqa9iNznF5H+3MtgBUfHQGf8BBQf4i
rLxIaGDxBDmfcmIpeQPjqgu6OT0SfIrgB2t7y1781ESYFVFgRifVtPr8z0A9GfCLzQXyV91Rswh9
wgPRnTkDyPMGzanhHqlm2oXZXMMgvKnE9kplogwMnxQVPHhzlv/KaRbTAeUFBjZC1MiZeAheK5t7
wTAKdSmn/ftNyTTvbBhZcUWtSCwnL5TLfeadUFU9hAPoIaaxUZuilCpf6JpfbwfFI7JzDXDDcfm8
Wr1AbNCjxbn3uVf0xvPO9NaIPCVLHOdX4KCNk/HtlzwiUn4fzhgPiAkEFtBBGY/8p8cVad4LpG+G
xfxp+P/lvbpdOkptaafr3qecCAJ7kr7m8PLn3ohO/rYCDl50Kglt13XWmqxeoCE6thAxTgpFeq9H
ZPhxnoH+IaBRKp2zOhzr3fjSeFsSWwhA9gy1KYQ0T04u3F2/s6L1gg0a9tMC/SjiYN5v6Pk/bWYM
adgwbRyXckKdpnZixzteFuLF/igADLFzJOmOCFGshIJr2fQiop0qmvEhypiNmFimxzkDJMocaznm
8m8acVin41OQU+uhLHKlcKoP7XpmaG/SpDcKxEz3/3mus+IIUVvR2uTKeMLg72cv6oKUWen0p2L4
wkF5hcLCDxyTp29LCd7R1qlOg71Yr1HKAjsoC5RoV0I41uJrDNFbdPQmxoQJKpHhi7Mf4pp3XY8c
2wZVUDt8eGY5qhdSLShlRYE5uSTK0gRRH5GYfi8ErZhmPcQaoDMVT9W9edxiyB4F2uGhX6V9IBH6
/wUGT6etBkfYrahtZQh4dlczpTUCEURJOZAmhYbg0XwvdBxp1V0iZGwbyFyVG1zoc7ofOu35Tvfk
mEi+a4y1mbeG0XgwwKeC9OQEw3Mrv1Rdft8NO+4ygW0NupSwr8stH9nIxAK5K4Xy5GId2Kd+FH6G
yNlOz0f25Rqg5AxzbN8QHeKDuxHZab/kVSEwEXVOOEMXPnstd73uk2T8L9AYI96LxeYb8iPKiyih
5nyvdpZSXuHb31cQ7lt/S8+8kfYMLuPRAX/ifiwwOXmyenRo6SrkImLs4W2HejGiIpwK632DQKV8
42Stnu9k5Z95St91fD2kxAJbeCU8Kf9DlTaiI7byXsw3wV3k9ArzSEUbLqPoLj+WDCFL8Mtk+4zC
kSExiO//+pkgq7ckXPOJgdQSAX/fq7P/ojJFo7OAZ0brpaZgDCJPMelM6LomQJzLi0c0P71p6rLM
DqrqtbWCoh7wrikJLwyjQqycR91c5Co7CPCzl+QvJyW98FkjPliyD4CQrzSCsKOJHO5NMHbb0Lxy
WKaJ0wqv+0mky58iUfvgENoP/m3DUSQ4FZ8vbgD6VjOFxL7Qq48xr4nHh/TlYpVCPU+/QjBZ30cu
fLIBks+0ijaQFX4QXnk9Izh7kbat1GpwRr4q0RnohX9FwpeMbKddcPDNh2zpN+ByQuj6WHmMCmD3
T/ugxu7VzAjTOumZmZvJQBmWJBMNLnMmf3B7zKltXyqjTfnoDtKjygROFcdI0weFpinwM6vfA9f/
exSbkqaSjY/piwelPAbiEY7SMwXjXcuPIGM6JB5FCg+g1qpijTUNzNyTMGON5+tK7fTfT71lp72y
h9dddRd31l4Q1LhSFiHq2e9v1DHqk54B0OmC08Bp1NFjQ0OPs9Nmc42yxlLLT6Ztw7sO5Z1g4PG4
g+vc0OYcWME2V3T+59a2GsFo477vhL/vzcz/MDY9JTqHGv1FaxXMzDU81XJfNhjqjjhgHIkqjy/H
spQYy1bVSm3TyCjRl11WJYu6hY7iLOzgyPPVomWG9r1PnmkAWym5uQQQcZ35Rg2c/VUKz3AtVMcC
LESC1TXMpJPB9pCRTDAh6EWsXSnAl8CbBdepm/hFXSuWphQyu+uKp4aqF5kL+8kLxgmGZByi29kr
Gk52UK566WXLLV6w3ZBfNdHETrleZk47yAKrwgwN1JBIRXdcsyDS+6WlFetgBS7Inc8OZ3+FqSv+
SfhAQzyaJwP+JqLMMLZsl/LJ/+MpEjaqIDXVVuYvwIFVErZV29FC4pZ4a61YPuERobncmjDckWgF
Ji5OmJvhJDuGKtdXCBG7sfNwb1U63P/pmX03IqtWzh0zCOJNZeaL15tgbFNrdU5dM0h77sCEMr5z
d6RZd4B+sQNhF/UCqNBC6O5TjOvEnn8B9TMMGIyuGY0xmgr+RydstVUaJ6XDtcK9chaFfN5tZY9d
uwFT89B0XjPoLagadwL+k3bIJqXd4rjFxVfg2LcYCcVGMvLZtdrk4ZmqbUfE5tNJ8dYweP/3QbqZ
adKqzxlOH1v4vGe4/8myNmVMrHKkT4+VaCrmH2K4T0yXESJQ/K9PZNuplLHpVvIHIvMNOOffQmWv
er67pC6KgD9duku1TCdW/UFdVEolIjxHvnnzW1KdnjJbXvuRde4Mvd+5oJUZeFF+IglPfiu5AAnX
DEkot/eg3KqQajG8rWjz8lcdvhYKaCW9GNXxMyFvLuYiLc/L2+cFdbOigzoTswEGWFrggarLr6Pw
TWJa40ZdNX3sApqGH9IBzwJcjqHCQzvF4BJKBuYVrog3LD/l0NBi9iSZI5CxqJqAUkD/dqseksbl
bWma0gZABewvUoim2Wq95w+out8/Tv+Q3BmG9pCDFeEbYVZ77p2t3hCwJGnhbAI2E2VxwReCdlJm
3+tvzeR0AQDZUifsrTf6imtfuzoqnRRXqqkTkyz/yhp8CBrYCnrk3dg1+eLkpMfsr8zPImcdidrh
LhA4Fzd+A1qVxWvkWzpYqVDv4geIZoQU5hLjJKZpxZGL3mpMyTksU6l/gGJN4t75bLUbQo+Lg9AW
/KOsElsPt1f8+W5/jnq6i7841aV8Ao8ZCfyZbRmaoqN63E86KAiCjN+adRJJnB2SvmhbLBkDZ5KK
P4EC1Cn0uVCDN1lA3OGx/Wb5pD73lIXTXsXpB2dyg8AYFhFxG2kIHqYhfL4w8CmjM8V1INq13CJA
tHCORUnNbN+8fmpIrADdBoM0I/PromAJsgPYqw8nbwwknMsegTZJAs57YwAm6GpycERcgwQQWPt2
BtPaVDOedkkQ7icKJ49Lqo7WgaXVcJg+xXUeUHkxyc1erLtme1RKLbrBDEk3w0W4XR+pPgoA9QBN
KTqnlyERNJ8pVPDAlxqYtT5d90MvTsg8WCPqJKyuQ3BkidO7AKYE2JPT8dgEgivDtmkbQhp4Bof0
vWWyMko6j5q1JZfUdtyCcxCLU976UklkP3FksamOD9hi61jcTqOivKoFrWq62G8X2ui6O64mMhei
kTyTgf+CUqalat/Q/H3EWunllEqXzUlBP8S8LFZkECZqOUA4ouCAWVlXZDx/8+tHmZAj95Y3YVMm
xq7NCq7eQNqkYJSyDoQpNtQgCC/RUYO/PNJolSQtagDJphx84hITqAJXYlNL6yvYLcN2VT/kR6EQ
VpwpxyuppnOlmUSlmC+ytXyOD2UR2xsrLvmdjPT7z6YZ8dh8I3xXACbgo+UUZc6SA3Wu+ryF2SNT
N/8Fo8La4JaGclmapPJHyvzpc7EdinVsoSg68TPDRlISzCq2FOmu32nqNZK/kiRMug9W7U5O7oeJ
1NQ4hIa6IWrLbQUNb441gYZmTh+Z0Ryfw0ydoCiCIepT/o1IbR0/Zej9JWIQkUsZ6F15Sk1ngyql
5UlliaNjDlZpvyFc5ei3QYKv99pjGVTpA2LOZTsPc1sZRoHX8C1vVrl4S4cVrg0io/Wk7Ze5nPp8
vqEyE/BpNG+7eLcEPMpAFbsGLq8M7HY/jluEc9gwWWOms1KI6olHfpu3iKofwyYz58wq2k/wynid
jIr9nrqAmtihxfUZ1Lu/DcoVVXCf5rqJi+b336fYgzr0W93GCcGhRGEiZ2NpUer3f1mJY/CpViQA
Af896F4/1Qx2WGL8wDt8huQ6JSQYWNz3VmhK5jOd5OGS+zmPJLcBdmurIOEtIpOZAJQSyxy4FN0R
H3ucNfUh1GHH82HipfencZxh21sZCkr2qT+fQ3I0qpXe0UkIhAyJ/VC67QZFskcWELOmM0SQPDsG
vNBZvHH65e9JdL3ZZF5xryd+CTEc+L9+30A+AtbgFY2o5UOgZ5h3KS1iHeZ1mn6Wrhln2R3HEO1p
HslDXPSH1Jp5ItGh00s7cttShmUbrDUbXViHysrf08Ih/j+sRwL5YjtBl9Bnc+xT9PX9a6jCUnuI
m/nZHMVVC7/+6eA2u20tZ3Y0luBbOW+4YR4xSYvgNo6rfYws4W4e7E/p9x8L02QNA4/IUHo4zHHs
vm8BNcUnIwQFlDW2e32BfULMemOESgPXYqDnslRgoO0dxfaghpwt4spM8wJsjsmtMZKQ07+SzbD5
5k6TNCOHC9+88nHcsP60V+Gk/OPT4rYnDQa7DJtlozcMIQSfyAkXEEKJ6eYJUHMu1zzx5sRLMUcV
Ao84TIi7AITmVkX7VKiA5hqGLRSkDkVK1aFqD4R1U0WzGy7tisNXTLdhYIkSiSSn2E4djULYFH3o
FUVMbBUdgM1hcZai5lizGvwsfWxr7pXFd+vZb8MnOyoe35QH5B1xkGkGiywm9diHg3VZdr2YYHoP
u4EG8t/zZKYpNw1RQs9a4b5ehUI3VtIWnecbee8Memts6Kzq8wSqmesCkG5UzA6Li5Et/Qpneje9
+lAFx4U5X1w43D5iEds9A3hg7MixX62fJUBYzpKrW84egm4EA9faCclFjbdDpVdalqWgOqeBR2Wj
+pbubQqzFALlblNk/myLZyDuDJOuXQXHsfPcz6o0jOgr6iesuWdafnqFxSuBJAXxAZ7N14HJhtGm
X85EaehgV18RNypiDGKSVyDIK+BnpJuvdrsD8wM9fRlA/NxLGH5m24k+RnXALh2pwPFk5ctzqRee
Dih43hvc+SJqGhRIvOtL/r7UhUNgJgIjef6+ASRBuvZKHnETxbhWG2kttYXbmoy9n0/CRYcvTgeU
pJeOjlw08Pt/lZcs3W5J/9YAxY6NMhiTpXGo1NA4e1OII3/UUixAkop8Iqcx99E7QMjvar/Sn/wr
2uEYq9WKVFfhjcsAHmpMe24xx+McLeEe6i2BAwUDV1aF8Ej9weAOMsUdJkIZGDjYreXkMm7qEI4+
eyFbFmQNzZyi69HoRAVXUEmmHtrY/bpwmLkTQSZtg1HhRoG6Zr1tS+TuuYU+8XrGvbAf5p/7zYBc
w0YbPL5RX96z5wvh7mDVjcTkNAOs+DLYtvf4Zkm8sPiFo3pSH8WyhYNMtPncUBqeNUwuqgVHX4cV
nUf6mLWE/wAOJE9olfjEACZRV5EytiUqcfxeX9jm+1jqVT6g98AKQyHbTBK7Jr7EBxFJ7p64MIhr
SgBJGO4ZT/xj6mF5C5bCvML0iAZNDUFDiQOXawAhoB83mKnNl6aSZVHy5C9X2yunuuGx2Mf3jUir
eRvA7DgBY9apcmT/pgpCfoBMExnRBIqU9HsbBSdt60vUcYOg2LnOWJfef+lChnu/s0O2f3SNfNhR
Ys9driQedlE/dyi6W9O7IbLYLK9CG8MzsqJAUMsDREHR8R+lt1elgDwho+NVzcGZVsIEkZFuXZQI
aa8A1GotaTiW+hh/bQcVeIdaSGFTt2wVCbWLn2c/v6pSu9r+WpIrN7lImMNtR6joKkbgpo+99x1x
qJhcNkxDl2EZ1BCMHuYvp5t0Z48lj3B1iCIDFBHvxyDcqk502KFwFrYoV9oyMRCtdqT68IlI+7jJ
sQ8xuLM5bBTn4oTTmlZ1T9H1Q+E2ahLIpdyIDgIlLyKK8uOoPqJ1y8DLPJpvKu3pMzvZCFO8sDkI
8lAj6JmS7X91U7d5++TDFTdZ/1Hof38PphUxfeON6R00IXn4G/8ONUzZUR0trsRI+HIF7GqJLfcZ
FnCSFxvIXmu6Y/FKTVjbramYt8hd3nklF2jfvCXy744qah+cx0Ygmmn6XTC/a+f3kWxEYnpQZyVr
mHpdarqgvqwAVqhx8JPRc38gXtiVGYLacdfFDJ9+v97/10gQvc9hN5vAeD8OoMqBQ1QFSyc4vdf+
q2h9PU6DVrNf8qzgI7/00VuPlwanT4vMlcpKhho5/IaFpsdiCFeBdCltAWcf1hNWQeiJnPMk0R6B
KL7FWHHCQZW4QncsNm2rwT2uo3ZZmYFeBLwajpmEqxGUKbmrSeYQNuKyK0NXqTjxHg/iqdIDJhBw
cI3BUmmG38LEsnTADtVOTxsYlWtLk01g2y+db6/NwyxHhlCwzN8elqS6uKsuR8kfxfnbt5dnJAy+
myWXOl3dp9m/u680Fk5UrMPNnJJDxeISqpcrVC7n69yrFpCgT8JDQ+cz/zv4drm9iYHgzXtmNg4T
ckhBGYO8exPEOZOgEMv1AC1MmhqtUvPP5XHTpZTxfGVgkKowDQ06hb3sA2Exk2KOpqSrMqGAw09R
lQBwUwP/00FVN+eTlMlmzWIE0oz9xWXV/chp70qLecjG6vOO13CEk41F+Hc0mnJXsCV6dSYY6Ua5
1AuufXiIYp6Auyb3TLJzg4uQRq5k8WeJtBzIws4PiOtG5W+YzE6SFDg+lwmyOIQPX2SvusrmEgR8
YXsIkhIfLPGZSg3/L5snVmd3sudEfhYJpzpHBhHoP+fOQPjcqUVoRPMufasISHfvNjJbh2y964Hz
vOvkhVkvkCh8XR5wgBIgqlZGF4wmx7b91QNLvoaDii/5tiW3UGuy7Sa45BYdqL3lKS/OaTZGIGtI
L8Rsd1tI5wnsJCiz8NUXQTuxkSxATMsiinFpG3ZFOaFENxY+DvQGcedf7YB7vWwM8mX7Pv4cJ8dJ
AWCdcCmjU8nAOdnNR3rfKFuE57TWMV53iZdDVk/tfWhWwX6uAKyw5AxxjlgKGlX4qtubiHUT0Tk/
ruGYhgwNKW80oyCnhdyBunj8ITNC0gvNgbhSnSD3feNlFzrkNauEaEa+Xd56XMg8DYe8qmNYKQNw
G3+mnlU8F3ODClAvVM8pmYjZR7SPSeKZKdenLC7rHXNy9dW7omQI1saLOKOxygJ/n52xwxw832ra
a3P88Ia4uYw5w2JvU3C3Ix78vTDlK12vU6oZqwQSM89b63WYpgPLvOX8SC27050FI0MiI2oRilbV
1zdcrDRCIaUzJZWgX7+QWfGASkCnMAV1hLDxzbi4rnn5LWqCu3gKIcIOlt+5YS7KIbFUf9HrQeEF
yukc/f0nuj3sWilt6ClqKO/839iUImKLyrW+0xtg3/VPklRCgGQhhjWRM95diPzkdpwMlH23TU/k
qbkr9jMVnOq6B/3ezYZ/tJtJiPnFXDuzlJp3neIOgwAtRESBFR3sRIvHBaz7agxSmR/Skz74bdIQ
oQFOHt/ipjJWBMEEmdwaslf7gycxIoEU/s2d/RtR/ICRarE6nJ0yEMl+tqT9mhirDIDDiwL9h1mG
MBfoyfspOBL/6tSjUtkgYWuxNHwxTrx6L6rF0RZ0d1yZsVZfutaFLBUV4F+NpXQi8zwzmamjmUmc
70MGJorNGHUN85BR+HGWaiuh4j8pnfDV3V4dEEgM/klSQLoZOHBsxelpMoZ5ifI/XuBNhLJUtKEN
90+nVH0SxkkiuGzOBxCY02sDt0126e8QmRflURQAQOHqrPPN9u8CDgYlTTKnnIchWszcRWRwE9Xu
Q3rdLw7juxJ8wjEoVBNM/dqLbZM2zoh1sEFzz8hBZBrvSFKM84eaIguvAZ2NRicJhapowUOqhh+G
lo4fwgTf9x6WLdvbIUvFnkqYGMunuaTHml+K5Kfo6YPUygNEKoLQXGfQYd7W+nPFWM7wKIB7xWdj
5qFcUj72A3WYFWXiDQbO41X7NXdDKkDpM6utTpr2bP8msHsLjqeLWLk9iL5DcfgIOCOCs0hkcOtM
DCPTjrQPetqM2rXYNR/K7OxrQqVCfc9aRcddDSNXDJh7Y3EEDwTmTNHhzTid5ESRp7Db3A5w9eA6
qGLMKrNVg5fRXJObLWq4ohaKCqylTVo/De5lgMnFmuW/rEs/4F63/gFrmJxL+jtwWtcs+A+b0cUp
/tuT29Pblqh4g+6yW6UkizEeoResSkwDu2Wx4LNQ0vkBqhgABgU/KIkBZ6vZHxNfBXNItQoWggjq
Cnb7hWlAWSm38CfmlfUVZkGJM3H+lS8gct4C5IbCr6vndk/8mHAXZtItEhApyTPVqEfNMNJ96L0r
MGHvCRhmZEqdmn3rD9BSA9a/XzHLhli3b7+o91wAN+GDTgwH++DX48cxtaII8vDzXb1WcWHYtbI3
gEW5mkV1KemKPy0nECrguZ/im9f66FwhqVH1EQbBc/qA5gNl0pxrykWDsLF4v5KouXu/KngclYph
zPAjV3dOxGb9xAThlcw52L0eaEXoSYEij/jFIDTevlAvZR5kH7GAdRfS7QAke+xBEvWBlL+4M6YE
JHHKqAmVMTE0wHvO9AwM7t5p3LH5uk0BJSIGizfn5wj3+LxpqTXeik3TfEHBLmZNZqvz5IvgnXmL
CIG+3AJJvGQnLOkTiyTL+5YU0kbbuoQv9h95Q+hAn6oU+PrXHgVX6ipYWAlrzRzB46BXeKZK2RlG
dyU9cds/RXYib3B1kKB3+GeYKVNyfeEr5h9iaCAU5mO43jwwO+3PZC9fbqmIoy5YaWNRd9yPGPlb
tI3ROBX6DVTAlWH3dpNex9Cqms9286AmeS75XDUiKY2gLDAUwczzDrx35D/o8KeFdgqhs7F8O0oR
3LZ6fsdu9srtpkK/n/soqWoWM7vrz4LPZYywZaXu3DB1GZWew/gD4Q5e+Zgr2KLRTu5501WIGpy4
uGMH4ZYpX3JkdbuN02rPChkWrikhUgjz3Py2/rmQh+gM+gA8snsKFZh6fB96S06jTY8cvjx+fNia
PREj47EAyzWY8flRAkl+TFdFpCZ9KUan9DJz1yXMFLoN5+FFf3WCy94VrfowLoWmb3IcawfCyjo3
SdLVOJ++8+RsnwROaZuXwO7t6mi3/IFMRxcdx64RJ83UqwEDAjDGkcy5/yTGjJHPGjkpTc2ielPy
B3XtTm9VdF/cZGtPDzWnlpO2HcMz0As/OU4bwlaSbRA06bSSZo/gXbiJiW15jf2uyoGAAO5CXRBr
czb3lUZd5fTNfdfJx0oo+PjGZOJURLG0IFAiXfNXvVQgUaCJsFysyNtNMdEnUlTZ4EdK2FHxY3qv
0PHTFF6sAsrmB8KsIi2RvU5MvrJlPv9g++4dJNit44gkgBLCUFSL2JaFwQmi7J3W26awScJZdxIP
YZJ68MS0Y9ZTWZUSWWji0hhQr3g/QJ4pNWR39lx2dPuQl25ksxTcOgcqPGfYoUr568PBn+CfvcEM
Mzfc0wDpZCrZXRaz1IMySs+9FORGPdSEqX3aCZRrmkAGmsTXWOgmVJ76YEHHsiBm7EECwYMfsfzr
l5myfLfOKc8e5TIvcFJoHxyIC1RVeklcEOvUaQWFK/7ZXRt9tDM2H0984++8WNUdL0H+CPIk8QMN
DGg4gQ1ez9FKJGnvA4UGjhwTXWw0l0G+F2UsD3ae+lI2S1w/t30Y/AUOLpbpZqJPd3elpR0FV+2D
wqVgHBQ46uPrQS4Df9oF1NgI/YC5WuZ+ZdiLw5NSfMZg+emoWPt58UB99+Q29BR97wYsUCK+woJ3
02yXPHbgp6XnsjUMLzVD2FUTNdGN8DzNf3l6L0S2EPIxkzTKIGK5bORC1xTZ2cVTvuC+4LGciyDr
VJEsPNG9H3bPkAhzw0+3eZKbC1EBkdt/8XB0T1bhrq+scWoPvmvy00HjlRWzOZyRKTowd5uiPzxn
PJkk/fbJ78IqVCjCrnHlSaV4dO5ak7RDEAMyReEyuLTgo2uc9LbOB40SlwijczX9wvlPveT9mqf2
WO2ubarl1HFE607bfBNL6i60bEN75k5myzrnYElvTmeCyyoWrEy6cD3MJ1i6wy+2YQ+4QFqLe4ks
ghyrt+TQbvzudC9ytbp0/LflQUilSaqqfw69nPJ76bB1jRYWp9AQrZ13Aqarr3+gMdMqk8xq9CMu
mlAooWWWi2qM38lrSoPLkPj2Pxns7opdyeFtUuG0VKG5QOPwr8im/cnVy2pu8EEJEeakmb2a8MdE
3/UIdo2IUOKc6NTgHyn7ysTG+Ha+0H/RHXhQaQzTF1y1zTRSmLsJfqWwZqOh82inr5S64OShxPXd
X99ukxMApHl8sTY2TohorLtZuyu2JkF+22ZC2UKS+4HJzEutOGSLULB1agBLv+ItL4FFElWq0dPu
3srOfuc2teBivHQZIz6Ov7Cij0c1YoK5/1+xgFY65RYQJCnqGJFjamHOcg/XRwvV89sPfLR44rAX
wulANXuFlChqT7uZKU66JwAH89yegFA1AG4vvvqQYI4Zy37tj1xHlgh7VXv9AvI56IELVG0=
`pragma protect end_protected
