// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
HWZUjVsd4kHYjX3LbBkoZquzE6R1TJoeZF2pV2dRMNSMlL3fBtpBeI3Jasg96yQ5GBrhvV7PB/95
qNvruMRT8pUl/36XXx6Ur61VEMLpaxxRcSnTgcEMLAs1P8zl64yDAdvHozhM1ixSNKBRq+IzvheM
UYI6IbK9zg5Sof89nVWhV9axKHluM4QgnOzQ2snYPr5KNRcRHSBAop366L2863AKU5IyV2AEmKQv
R1OOk4iUZbIMdMvPXLgB2BF8VeZX5cgmlhrFJ10h9/TEL7QLp+xaV0XjRDB7ibtNcls6/bFBASyY
9FfG+qlbsKFgayEoXKw8L4cUnuickwswkR61+Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
hZCt5+5PJsGvhod5MudczMLwmtPCSs+z+MhU45czn/MSmmCMuRvcxOVLTGJSmY7krF/RVN73gCsP
C88AkTi8dPtp1m0TeVuo1SmALJS1UU+BEc26J8IOWtIA+GhqidZh8oTtr7gkWl+KUVZ7lWE8NnRi
KItGNbJIcFBb9dnDSwXZsCu+MMm4uZWFO25cUC7ijHv1f+M5bfvZbzvFYvNR2GaP+NpkVXfT2VSn
mTDlpY/q4+UMYvq8HW6mH9Yn7gpQxwJkdJWD+Z1zCqKvwAPlJlvBc5MxVArXU+l+BpnyepswuTFu
H4VxSJ7cImh3ej3tmEQ2wZTKtPC0LcEampdlrYBrsf8W7Fj3hZqYiJnGiFz8dFI5AKxxsg/nbtzk
abjZwjesiEp3Zpq5AddUlC6S5ENna9wBoWcLCtdP3G07qXZe+UpRKxufFh8oyn4cr6I9Wrg+Jn4v
sRM7VCYTAU4rKBL67KUuin02wOzWZcVXMAXKmGYr7tf6BZ5AZoMdsx9xpKrVnThPoZGWeAJu6n2k
dSylvhV3lzniYtitr4AJ/5Q+zIAxUWvkQ4zsmu5hNlanJxImcYVM2a0s3hZIXoQZPccCZwHgnEp6
n11GUDvaAKKQA6whhF+yExklgs2+Qb9nryHzsDZGA2eZSD0ArRfXkvkNeuMhwKihDbmWi/2p293/
S6Sxcg0EiuiadHHf3rP44qrp/ZTjsWMctY3aAleaWWxZZcrDA+AAzr2y4nsHQNs92DQ60N8uMoTP
GeV6Ttx3NeoX4S4pDAMxuC9a/w+hMuU828sIjtx5rx4DY/sIYBGU7GiE9Ru09+MHNIBzJO/rueaz
MLCNZCjnA26LvYsi7JbLBiEl86kQfxVWNqhukIVNDElKx/SbOd8FTwoJBaw96bp6uB6WGA9V5XLk
JfCAr+jJy01ibSl8vhhVI/HSH0szIxxUqI7mLip8/Mmvcvr93ka7WZWfeZ/dleuQLeyNsH6veBeV
zO7al0lC7hKe0a4czptEaf0GJtGxJ6mMCfZuJLPpr8zwYI5uMYR+o6gwhsGmrhEGFHMqBwJlC54v
VejXm3oi+fwUm9mA1iwK9pomavIYG9vv+Pgnz2RB5G/SpIJ2+yPDLnOanCtA6UqYBZ0MKkenXeA2
StKPftnQeLKPz5wBluJpSqQf7dTM0cXhgPJuiL70N9SGcLL2fMPS4DpXYBb2RFmutdDr4MXYSf6v
6gi+LMVOwWMfisj8IK0Q1jddl2QLAXdyFcwh8rmEnoHFf4vh8RIDrLjsdLdDpXcaMAC32w4518Dj
cEBjwBvo3dIQ2xUBj6/Pi/WzMNI31L8oXABM3M0+tGYgHkcEM4nCVlv8Jy/TeF08wCcQtVH69d1l
Bb/94VH6dF5s8eQRaySrUWYIPFbux0D6lZIKisS6eH76P9FKQebboIGrQLOLsH5IVvO0fPJD6jJR
pkaLT0biUtGyE8NUPqyUL7EpSPN6SpMva1CiSkLC+1xCqTxQsznHKeZTowKXbuBC5xTXikcMec6j
sOZlGIQad08iuQzYAEFe46zf+ShlzEcIH2NO56wzkU/Vy9mpwCLIenSwO+4mhdOyEeSrkq/njwX7
xr0cRr1pTR1RQnQgWbpeceAuBlw+4QpkmlCJSvFun8VsqWENjIOmBqwAJ1KIzx4s4/2pG+aD3BWZ
9AMxDLk4eqkceXZ5atzWzaZNwyFRYv6or+EbjS5/fBREID46SPReSnJdpUQtP6nDwVo095ryeErb
BalWxfvQxD2fViyAV8jAvcrRWLmxJeAvUsrziivck7rO3u/KGK5VoCwp4Hd1G3h22rKfrQUve4y4
r1n2YgocnxzrDMOspWOxbVo5sCvMaYZ3ADtbmJpwwmSvsnFG+tbZmxCmLbUbI1CH5h0nWTU2+BZK
0h6XBnTotR5NtXxg6ofsMJ0ixIMb7O2ER7V3owyw6o1m77Nt5sAF7cdNsgKQW66JbjblQ1HjtzqN
Ow2GEIKHYCmHXGP7jkd4AuU89CgoSBudtzrq5MpXxC6uTY9lI85vUU8CUE1Clm6Ijq3vmQDU2qHM
Ho3TCqEowvpECkLLSXs06IoP3ldHSvZYeBo8AiGRgO1sKsNWwk1TI6Cou2P+fxxjzfrXatvFu7g2
BzvWplLOSz9sn0aXvUx5kC/jHecQs/r4gDvzvSxV82izMwi7BTPQW5s6qnCwRaorYDyGuEbY0lTR
U1+Wsjhb8UJLhBwdnILXEqiIrnivrbgf3Ptpy3DrFkgQmXTMQmOOtncIufQf7IxwXNgWXLfykhj+
ZDWUIPvfLoI4RX7Nzl52c/3plXDXzjgfdZlygE2Z6k6kG3YwAvPBNiCVvWCpAtgQ1dKEQP6K7FBL
Ttzm6tYz7dRqzpdRgIcqETxW3u5uxZFQHUi4Q8m2ExiLgpycdSr97YnYOI/+VLmBw4nQ5Ki8a3PZ
GHk0oA1FwZ7/S7ZS/KV3dCFUJuFyKEPMoSmo6xXIdFwm5kbw5AQMuNED4YeWsJMemBDkEkmIKRVf
4XXX6imH/K6JLz2SrmsOV6bpjOD1Umx1jUG0Ay5gVPkWQT5k6E3lI4RGcmzyfa6jGqwyScxZ60Yu
CjpBKmPrkeycIwaAaf5kGkF7Aez2HXPisdCofcpN16h1otijy4jP/sC5tb2/mNPaOevrCeq2HSIl
nBpRRMOYO7E+uwc9PX5UasU8An7m1meZ57iPJA+tX1IYK1YSxIaozwYdv7oDKcj2/6QYUix+KLfb
VNbmRsmrSXVBYIaOp6LzXpKdZgSkbbsABEJue6PHMzc6W+lpUtngCeP7HuRPy8z8RWsPWjr7XD/s
BFCyY48OrITWMGTR3FinNRWTUCzp61ZjBQkEPaJ+vSC03zZ0EjEKLa9iLeuFmoiMSJcPsU0LXsD8
SCiNeynM8dMoJI60gWpBT8HTmGMxu1/CXjcUdYXPzjq4tz8EzoC8xyqG7I3walWPjYBF2/+nd52A
LG3tHB+/apDpaodF5Y1w0X/TZ4ETQPLlRuhZ8zZNUdEwSfo1ylHVHOGae1jOw48u7zC2HperRJY8
towf4bi+KVdaAi6gNNOIddyEHPhMaWEGsMh/eu4u0rxKLcnHsjKULIJ7ACB2YMYgHlsR4JBHBm2D
lLLn6nipna7rxCQA6DiIeb6IO8pPhSiZAJB/jxtLleQgnGDiiAkTfTB3jGlZy9uyRvfAu7EvdJFv
IHrgnR6pb6kf8AMXvBFp+lS+e1g9NkCgviMt3hoWyxtNE83eDV6S/OB/oOr8rckxMcPwOqtzAXp6
iZ/j9rJBZRW/6QoFWGmxibaOilvOQX1vVaXgbqdIBxm1UxoVS2ePYQhGoaBjLtCy/a/fNCRN/3vx
1XD6e6nK6Cy5DME46P2DVx92mpCoWqPduausjWFXLS+UIxvlqQooj6LL6DfRHFRP4ALEIfa8qSdP
MPNOngTVpmBvwwGmTBXXKebvwTbFIb3jDzCjAE/ZHoHHppZA/3Zk4vap0XZpQIEL+SpWWYIhzDuS
2kphuX18EQqWx2u33LG8t3ufJpOa4G0FxG5BaOOYaPAwZDp8xkx5WlNEV23alIicTTdIvFtEsKGy
pSQ88Uyw4Xav5V5UUVYIHWqVoTOS4OWlgRiq9osOejg+c6bnZi77WK7Ng/EDvd8EbQi86lUv5Idz
4y19Hc/GQTETwlCbjD08ThvqOtZ8Y9/wvjZSHBxqRWOdPubwhtaLbjadqhUHXL24Or0sKXs19QoC
4CHafda/a9ElGWtuTPPP8pFv8GCaD3D2B6cEw+C1A8xyEvvWmmNZS4an9nTz3UHD+vEm7TT66Ut8
xXljCSXY5X12Mv5PlEqHBTZmFBFACxXSPTeiJBfTodtXEyl/9dbD32CGgDm8umR0V4HWhLyDCOAx
iUMJWG9AzmMEHKCTZ+6mLZXmBuKSoe4OaqwGa1cCLCNkEn3PLo4J+rQE0G+C3nwKqXp6lpZ18ryh
O6Im4UoAyeWaQ07JeLThQMkd9SJvw2eGI1PxLZcfsq/eZRv5s3TVu5oU0cPB/NrYfeGLGlyZwXL7
oN7zI50vB51D/62uDl75xhZc+1wDcKSMIv1F+Yv/AhWoTMhFv3X8/KCjX6iThdsizXe/RAkKePlX
U8M+zcNw64RaxtuRZQBy1rm+PRQU5X0EyxJK+AJ4SUeky36GTHkv6lrI7c4bngMeD7sfSv0itrD4
MIJfJ4S41hI8+YXFmZ58pYBR01w9gIc1alNj7BlQ5zO19AJUWgvXlyqLTvAQOJbpOo+UtX0e37ln
TulHwPe9uetBs/iMaVEgfEXLNMs+1282W1yeUeE8crMA8iJagDSj2mEJhJTShm9M3h/i6pLbnek5
csczV7DvLScyzBDmw606l2Z5GwBmDyqzMINSwMJo5CMBx6WMh0B76yvjDciSyVclbWu52jAY//zE
8V/lH6ZLdcY6bkO+pEfd9ALJSyfePhjouEj8lD3A5jXtrszRUhah1dsO0rfB/x4dPn4ppSnAGfPS
PEZ/hOROmODQj76w4RfgxgxrphUqMNiZ1TGUjw8JEtC6Em3l17KBRgEY+T6tWZuJITqYJ7IrJ2s6
LrEIAac8BCniEcdcp9Tz1FsF52oN9BeQVQcmpgQFFFHPQMjPdv7JCUXubobUM/0svJWyfJ5jDCUd
3YRNqlHwBzOSEUOydfglopWxkl+yP434pSPp08/1Mj9Ed2pnVxvqwWBxPnehXejgcCr4+BrnuWRm
MMK20pxUN722eDClw9OydZ4KS4hov+GusOiA8GKUA23K26OKX1AuLF48d7q7wJKlWOJ6HLdHjRZr
w+tBclGmIDoIdHIVtkEF9gtfx1ggwoKZM8YsMA6szJ9N1z4htpn97NXDzBBHXsWUhEfZFXmLNqCO
ME3JDXMqNWJoL7jeMKCjCYpBE7cE0HvVyx86ydngO/BCbsqxIoX7KCIb6fux7bPE6xDVEwg6b5Mh
DgXugbzVNSJwY8NIksf9LA5XoKgKOv4wNuyaexPS5oehLahc51cMckcSM0LLstauI0jSisfm1m6i
55m/x3odNE/517QPB8L77d00/pZBvR9cVc7FM4PagiY5jsoU8FUtFn3CzP5eRnwtdT5gLMIoCkN7
lgXeO30/g0u6QwBvted7QsfYfdQTvtUHww8i95xRLpntdYiw7j1AKeLVTtLKBIDYc+KQveUbvhl2
fQHmZItWMNhA0Y+37HaeeZCA9GKyGUTlAUqNYu4ZgPYTWciF95w9CGv7yZyIR4k+VrcRSo6fN15W
Zed2zA4nf3C/a89wXcrF8K1oBX3sBh2au/MV61wCKMJOaEIgmdc2VmsmFKQBiPPCqpCqTs2oX4IN
y3ayIOjfCrsDZ3D+KGqUKyRvJGtPpAnahM3GJK26mPyKujhywaajgFaDeW3IqmR5xacCnVm+9Sel
0212tFKnI0Q7oGvpx9PHG7UrSjOFhktYa/ii1HtORH1n30M791ucduEJk4Z3fBBvFL0XWlpOpjRO
QSptEO1QsngfVqtCV1t/j4B57Vjedt1F4WRRK+vSTWQowVvH94/SFc/H1LEZjHPjKyoamo6SjWNd
l0hUWoh0LMGjvMK0XvWImx0eRisQg6nY/gkgoEDFBidqLqTOR7uqZ8z3nT4io6hYnVZvjzvWZGgo
hE4IGF9XdgcfNeGbxTyreTAwtfCbHytBEIVZMK2yWfcweClFgyHX3B7Mrcv/+f8bUVq2pMzgGPTC
7W95ky+ozSKM6zREVzOZ0u6ZCfkDO+PZsY6AWI2ou2pUyst+IF2VYzXpgN0fj6BHrGNWBgtwpccS
ZxEtUCnaym836reWlKnVlCjg/5U8cvFfbnUeXfk6an0siQ/Rb8yQdiydLHYGCGFT9wO3AmMfLa96
LVmSNfPKCoO3ZkHQitwuQcjaVpyui7GIfYWESmxUn+h8bBCDNemjWZs4Hp8HRPdbgcV/He7K7tEe
++vq+l2T4k9e3Pjy+ZwPeWDraHRz/CLMA4OeYs9odL/UniobGlFupfJjHjD9wXXh2V7x6eS6hp4e
DX6T1sT/b9pFxCXvjPrRDbczpB90P8cgyZV6CTrg692gryMhYyGHl/kHeoNpv2fkJ3l3hoZsHAZf
ALDiylsWgAIr/u3g7Bi0mgMWti/nCiiAbeKLwE/el2lvF3PM6TQvUfX1Et5v5PXWzu6PSFoUl/gy
wPFhCa4iKAn+C9KG4+ySIowlQLPnUNhzmJoeuJ8PEh0eCAkAt+az9uGCvTzVF3TDyydIE0hMVrx3
Q2DEe01Cpx8awpCiar17RUO66qp0a/leQv9x+pddJErzeCRACaMJSrcW/STYk0U8zRsNTj0AxVfE
OzmKXjYuwZfTT8ccJUSK7xDwiYipZMtffqzAqmMw46W07y/ns2z4fSO48kZFwbXKquKk5WSIe3SP
QV0XGopY6PsUPmLFYWK8/z7cgsSV7X4kIKFeP2F8/zWJw5PTzl8UMPqGx8GBFhS+I9faVp54v6yS
bMpMu9ZdGO5okgX/4n/2PIHNFkQ7hLKaBxKXz60/Ya4pALNeWBIoCyA8O0ZTeiVgDplth79fJoSm
IcHpFzUYfPDyKtyAWjtYbtsnMpYaKfrKd/7nxuzCMYz7ru26PcEX3uzOoPl+9hPkwXeuyWFOnUQA
vJ7ukH30eLSumzONUd2BA6KdLMUgunyABKXV5wE/4+xf8XfXDoeKTXNpoGbAKimoSQXQSdrMMNRw
Y5aX0d1wGHw6DafB0BxB5x9P4t8XJIha/xfLcB9SojHU/CvHTGRBBUjyo89ihSPflRw/duvHO5vk
gNQYXtKyK42pzOM+4GYO4HXeflqKAmM7zJ616uXIJ4Lx8dkQYcTKDeOZxe6YjwOlXImGRPGJaPgL
D6wwILENGXI4NrPgpMV5chHmz6C3ypECK7mT8VXHd/xCLb7lTSIvuhX2RmUa79GjOQTlUQxx6FnD
Jm00KPjunGgIelM3NKq9+e0peOw7j7Xj1ZXoXYCv7xEsOomVsAMgpujUC8MjpsOM0PfwsP3o1kOn
e7mInrYuyMT3u8TL0EV9hfkn7QkHk3bJwkANppP3cAYlaPjdASAeBl2LzXj1M2VkQMDgt7K+vcMo
ifROAgxTdwa/RjbkqHgaituOe5lf4a2om4j8oqII0jcmw/5uPiDYVbaHCPOmYuclkrPDFpaqGCd1
qFjt/g/uLT0tYEXH9z7PQeyo3KTdMmHT5UotYJMkp/wl/ws/lMuTUBnddh7pzydiu5QyW26Dpi0q
skpHY018A6j084LSPoOihMwo0reiL7yJqcN6b79/HbnJfkBG798D0fd6oZXrlvCDCfXstsXpi5Fk
97ZumcyekmArV6CSmFrtBhY7YgynPDckDzxj8nEllFsB7RLvw7bCn/jvn5/tJ/VTB3L9AnyhAbnw
2fnyO0hkNftckfFvtKahlT9KJSz2XC2j6/cFjxqqBcv8psiwF+uMd5/K79yv1sT+QCk5APxLR95x
scnmHjXffF+pwBQCKuJQHzpaQ75LAdo1Fl9JdFwA7XugpPYtfO2RqIqT3RBjt4CBw4SOyteVNSDa
8Xozw/8nEIWE2rIKmstWNSZhX08mGmTu3oPjJedBzdrK1+kHduO3QlF1KJdpt8PvFBMU4NGF5DmT
/cggEltBHVGb7KkE8NXavKvEEZIj4b6ZaS4ZFeQxdBA/DL0Sn3zk8GZVz36EwWjQThLUmk5yBwVb
PUjvNl+L3tGp7LFUf6qxP8RzcSoxtsXnyIgyji2d5Cx5aF197XkSOEKkpDKWaovO5jmRkOgniVzx
yxk3xoUL+Qf1VwzerHvt29JObvW/w8LtKM220Sldn+NMGHbkcKZ0xYtpl3BmnbVH2L/Cguv0yDKx
/iqgSzqwi7PHMrcTpwbq8LQ8l+n7PUL/keCrhpgkm1ZcV0UC5dfrrxzgDGbMvwCTD94RtKZ/2ju6
plHbYJ/iwfOaGVaaDn2emKT6TGCd5gjoCgn6f42SJIVkh3FYxwJmxtRbo0SHzYwtTwvHX3edOt5E
e5WiwO5Zf2m6Cxiv78QRt4xn+jCXz6UU9pSBpwyQCCJrL5qcdBrThvlmIpoEl//Y3CO24wUL3MAX
sjjOE0vmm3JjG5X3MwPZvb4EchArN5PFy5SlAd9uZ1xc9ZZGEtolPa6DCmk9gqIVa5UPAxKEx4VH
0t/GI3qiOk3tKLL4gFRqHRBZ+NKzP9eLeiGnMxk/i8nITowF17ZXWocv3a2wR8A4mYEVsoyH2J2M
ZqL725KQPa7zhfkqse2sNNNGXCyGGRPu9g2EwvOGRAbk0sW5cvdyw/ueIEYLeGrxI3YqOrbEJqQt
c55oy8K6Fu092EJKEPYs40SD+DKfBN1fdz9j9TvpjloAmeR8P3uZc3t/FWzxpRb6bl+VkA2M6AgM
tPKm9WCOGZ1NC92yumWgcJUY/22RCq3HE9sqmAZOPM089wEL/bnqYSq7nGM3VDFmJ17GnCaFeOBJ
2gt4h7NpVHDmLmMSDICSR3ZtuOlAEtMvy1NVxScmC0/uke3o4Jaq+rHdk1h1Y2uLYtbLA6s7yLKX
T0PT0/oDyGjcCtJyUVQQDqFg+OVebiarJ5qaK0zmgWd9GpH2A2wJqLNOJXWM5NU0kdcH+xTvLjyo
eN1aGsZAatcRdxq46rA34YwFN7/j6lH5Ep9lKv1ChLvPox/2x3FxlJul2//ZtvgbYXHwX6rYkAeH
L7ZsHETMEnFI9vw02lnZzBo3gpu5nM74YfMvnujotacVf8FvJ16QKVmdK5SrhbRxPZau/mAqDqSV
Nz2FSkzi/IGnq9nqm9wMxzA/KS4E+gQrsQEwmeHlNwQgC4gVXlT8f/LnVg+96lhYV4MPbYqsds6i
h7am+hwW6GIKjooEmS+3vkzkjuZ4+fwiJ03EkLDxD8l32cC6UuhUNVY4owARUpyX8XR6T/rnStHE
zsZ2f5bJfC+dB9coQAmKMYkYWhV7khXGPJQQVek30tcdLHTpCNdYjZ+ktGrZWL2x5Kp0Iq2UTXov
vpG3TbpvsKR/7l8pLUorFLWJpjdE9uUCWP/Lrr3SEuBajGnFcFipRnkr2D+O6rSPaML4nkZAtnXG
tMD5dn1xHgiNSNncLAJ0cuCg54nv0KO3hl3NOQRiI6yreukURygbbtZ5z7pMz06BStB21w2lhDtX
yAt/H0JkbFM46eVUjE6RYX+T/ndDNGCHCpNS6F/ar9jDA+csYn2Ry1GruiMBSUl0d0YVPP+dKhLO
xdN4QgTGMu1DbPjFWym0XUvX0KsEy0hrb1P/e9C+JnnA0ZnwMTF3WG4tKGzfWWw0tvn7MdELT6vD
p8k45EPyPXPm/+Zx9Z1+bxLNhYWnuxbOoNOSuJLW4hfhVucmRVO9hXB5LjLz9ZX7YgIU71R4QI4E
nqrmH5qvZFc2ByLUIB2G1aN+zC/XGly90yLfsvjjv7L0DAqGnpyTGEarmgMZN+xpyU33/27/IAFq
CpIR0kiNlNxsR8Ys5cSDT44zebUHZ7hl1HaRKTLAOc0P60dTtrHp+LijRw4ecP+Yq2qrcSkUWMwQ
rud/Qqr10+QxYmtWe+ykHlgC6HoxYrVHJRttfxdqX7avIvnDjQAx2x+ipKm8ymSd6zdRRtF7rbjK
yS+lF1y5vv4FXs+3vIsqcFdVEjStZUmp9scp2l3HcK8+qTVOPcNsJOkw9AyFAYrNwPjiAJIA6POH
xMGKzCH4OI6gwnonXDWKLwQzOk43raIwP0pJydkCWxesK4oTHeghz7N+AMuVcpXx1gblk3TR97GZ
QTjN15yv/LHCA2qF6L7+Ut2SWFgDAovM0WOZy2vZiHx6C3EK/SnLYMCvdbRgXkA7JtQ/gqIprqoK
fBDvV09ezTmWQZL9VKTArl4fs8xslxyLUYzKVUe0LQldv79gKnXo+L+wsFfSFeTcsEaiP/xJS1Ie
cQhNzD3Pqh+daibXdMvDxjBzbpWd292ShEDqCHksDhkmiICVqJOowR5yW+3Yx8d/1G3sonGdQbJb
Wdwv3oUZsNuMSO5zneKvtp7Kw8XdcJgbvLDJ+8E8C1e6L+kZskKXcKRdT5wAhACQJIqAf70K7kCA
F1iAUK5fgqFt0gIVXSNghl0fqqkSDvLmsxmsHSsVNqPq1rz07P+Zj10V0ZII80jPzSeX4ngdADbJ
SkKy/RTcTMAfV3VkGyQ3IxERjW1YpS19kqUW0NShAspBF9L0ZWd0SxAtsPsgcI/+6YQfDnrbPWlx
nHLfzA+HvsxfxAgEFj3B3Wo3bHEqDfGyzMTiK+mlEQd1HF6CFQy/QsyzLyjH4nnFwTjzXZNmaaI4
zBsdGF7RyoSGWmuU5KhQpsOz+vrujwaiox5eZ1iK5yv6xIRd5Goz2MlCIjH/7KCHp7uNyLZztxXS
9kHuMQEMc78QDmMdpj5px+nguI4ihFeHylQ2Oc/q6ieqpKv34cu95a2oyH8cI1DYs4pOPJu/XIgg
4M8oIJpU2IbY3UJfqv4IApndvGq9UnBtxEccEe1J28inyRXiKIgnqqtyBSxlqVw+WKsaYTQh4Q8D
hH8abgXCCFcZzh99eMfjxPJr5l+N4ZcPMWbMl+AjSxOWo/Jnn2pbTG9qEN69rtSosqxMRiXwgNp2
VOGZHPNv7G+VAp0zJhwe4ZYRJKzuuJRZJEy7MBdjZGRV1+oxKPwAkR7cNZs2LjWfxW7o+YPQIhhC
rnEjE2lIAIjOC16emUansU/FVqz4mt3di1umIh5ffE+slRZ7SoSgWi3m0KOC8Lzgw8YNV8QgW4X2
ryO/jYikXNzmb1nD7T9jmP404gVMmhx0OWUgauUEdWdejKC2+2r7wXSx8PCYkzxYoYQyIuVQYx7K
3PFYUBBal4TudjR1IiXAoKADGi+0YAkufxco5oTUZDANnd1sz8DvKPy3jgdZyzrWMLwpH469Nhg6
klutCFpnewTlyrf7ZCjHkxVnj+UwzFyly9WDZWxGB4T8Ptx+Zj7Zko6YffLF/39wL4EZiGFo+k8D
0Uc+dBAcnMDA8kegxoBCWb4CuANiZtkIGHnvByHZqRAhjpfW0A8uNLRKcDwy+aoWQZ+NPEmVLY3d
GlmHWSdG9YrQZ9mFMY1OrqbupgRrN7P/a2kKJ+uP8o8wfWyk9p70c+/iXhQImg1pknOImpSGKIn4
VYaWpj0CC03J+B9uQ7+k7aa4fwMXqpTyS6EpH4sXSvM8TUnEAo5ChsnGT2dQ+gjkS3i5kdf1Isp/
ldEFhFApX4umbe1N1ZZfjLz6+28vav1Jh09U0pwk9eIoC06nEFqJq1eE0sk4Fvi5D2caqvIKUkUe
wiy2GnoKgQY/4t3SXBA8h1QNj0ynupPQZvpKPcYSZ6NenRuvCTZnR2WeQj+SzQJ+ogsGGC5IORqd
x7sB69gUwClaTHe6sCEkUmD3TrcekX5ddDPTyjq0uFP5eFr2qANQ5XHXnh90nxqylDgEIbDPpEUL
xNJQBqGavkSWG6LWyL2sLWNEfGyUTVN+EfXOFfT7EOOJpUWlQujbt6MuQCAmMxlINr6+XnTiHn6F
0wnUUEyBlkumdrkzfe0AL+vObkMuuz/r3cCAyvU3WqafDli3uRnrj2IyXymoaXIuprlMobrWRGBe
NM7XK3Ju2ifvfcxYcZDXjMJtcfjrcaSaSl92SspadT1ozhW0pFkU9SkKzXLVMjgqPwuZo1iCJqCG
z34yrP0GuHDV7lN7XNIkJs33+aC/uUKEDBi94089b0RukR3deb0fTUd59l6ulPm2pg3xT9XzJcX8
Udgchbcxu8pGmZCTQv0mhU2Eq69WB82wGHrrS+GUJ510SZmVKUQ/K2jRKQ6vq+n7hBiTQLNxNkse
bDA/q4JBF+dA+2qZN5vpaU5vFn2IcdgMDvRndHe0KQal3NPPl7iMDgCmtP/vbrIypSSvVg5QMs1s
g+XWEuwZfNqg5gA65t6y8Y9Vc17rN7PWrFm+rUNVpaQ4sOlSlwO7eFr1Byg7oybUlnWiV3eFUHI5
XDZO2P39kjjQU3E18rjnuBW4Gf8tpMM212MwfXFZIDzajExdRg3zA4ttDDaxCma2Mw2Le/LZSgdf
FiFNalgMPQE29OomqmfoD1bvpo1/De0VEcS442f/xGJvV6EMg7NywlEp1By3eDExt1KbvyLaWa3+
9WHA95E5csWK9jj2zPR05w5bcHIsElS2M2GPxkE2q03e4lIkruKce+19mHLyI8eDPhJwQQL0w7aY
4mN/bKBxOcTKMBsr3PKcMj4wcrxI4Kxx9Sd25ZuhMhFhMl2C6pUg8MIlLK9K4+01AOdM+1L5bPCM
QtxW2UXy1UKOcOEAa2NnUO0m9nWKvarYvgdlka/1M3Qo2KOxi/KeeoBmp6vrVEeh8IYOsjfH+zKr
sWAWGzZhW3+LLU97VEilAsuUGZ5vOWLQh0SUR5VBR9lorzuUXwxG/lPCrgohzd+oV59s87pj41Mj
gaTDFKrTAi5waTicaQ7MUGqF/7GvHyR12hJJmwGRYJkTyx25T0uMAqhEMizNxD2FiGuaBK/AxCJ+
Fzs9Amr7JGNivtSLxg9AdfDqfzNkOQoaR+wiT+oB7roEndWNyh+LCAQM0neET1K758gX0yNze78W
oaTpX1iO6zDTHE5v6AbPGAYEaQGdR+74MYTtqxC2D6GmY11TVoJ9lQah40UHZNSlkkuyfnbQhGse
NgW+3Anjpb58+mEBsLIqKg3ZJ7PQRnL20bAGygsrJWlzpU/lS+PufDBKxI6qVvqjHEQXnc1Dm0Mx
1Slfwk3T9bNz6VcbEng2zaMg2+PuYW/IX3IoeYFOaomkrFVxXO9R8wt18JN/gABtdqCA+ioHDD7j
kiwFcO6uxpE435sk6sIcZPs/sMq2Zlsvrldr85Zfik7c1Pc3l4Ajhb1HdbQYJgorvbKQb1qkYtI+
MxaqeYpmxS7l+rH5bAwycSYj9GT4vngvefO6+6cZ+dlCKPxkYnTYYplUBnFeHOF31hgx1QtOg7v1
bLjwt90mJFam7PDyuv2LZy1zj0fUkZSfxhuSEvqmWn5lfJ+5Bb2LoHWbf4GmLDBVfni+LeXRb6h3
SCIDZ+Bq8LUUOY6bVarZosrcRccHy3V1O0xz8yRC5mYaNwm35hQk3ugXyClw5NIxBPuXbqLKiJSj
AeMMfaPw/fAgtW13fYQU2FPtfQABs8RFzzyTzo3qC2yjwUBPp5vPpUKW69pfC0jmjOu7l9yxw0gC
/bwOi1MkJi0t4B0R0HzD5/EfD62XaJwzXjONanrATRP7JFfIVAWr3c+iuTJ/LmeERvRR8MPs14hZ
GEak4KJKPzYnbu1K40P1kiIYjuVGWqSyKPaQlzT1QtIDH8mTMSQOVdDrqMzC+n+ulwyZbvvoNHXL
FWeiNWc4YrjjrdXlkX3gZKZn4qcvW0xD3obuPWUKr9bwwdxYsl16CdWBFexOCRJqTk+DWZpt6XfD
T6Nl7Wgkm4AzsfHO2uwFm+nKzx52cZH38BnWDwGjzYURhvjWHIseKqqcblom1Qxmf7eH6A+UhyB7
bOUvdr9mNPZqZzoVfJPu+wC+R/8nP7zE3lUw7bO1XKjiQ9/cEHn5OcUHBMWVitV6+wTcx1tE3yGI
Ktgs0/wBfxE3HTSVBc5Msrw3B+BJ//3f4fTRcQ3WcqIcmzGnFBRfqZ4MM8ScKcn3r1S7a55nBpCD
O2i2LNmmGgVQQXZjxczvx4nBdwKnrX9j2McKNOZVA7Nn2dkE9sMV4Wk7euqeRJeW84nb26rYsnKN
yRB8LE2rTLXtWc8oNkujUKp4UlXKsTAFPUShXq/LbdRk2aXLu5F2SV1DcyD0lSW1tTQsYBh6KRs7
jdoaYEPSvRTR3a/QeLUcEZwzH077hDN9IyKNmxIyc01uR6yr6kvot4THCPZD0bOrqa8gDlCNCWNi
Qb6oEthj/GpAm9fZynfSKagfCNlIKRRedTyqxVvsKREtlF1AFPPFVYghbH1goT1XyZWybT0hTW0X
8Ww4667iKRelgcG+nEKFdGgCxwPYj8KXnfExq8J44IAp126H3j2FgnrGfNFwgFFhl0y4sEWWE9J5
LFh8ZNUg7Pt3zP6tJP7+Xvp2+JAPddz3gnEALcE2CqjAo6ZlBieyWJKvHVFBhoNbezu0AIrZgXTX
F4lDeIgLzhza135dnhpzN3Ki9SS6JKrx2PUNXe0LQogfO57IGhLvMRu7r/Sq7gYpEC4lNIb7bdmV
9BNkvuygMk6NdEp/KeRtZ3I/7aVp3AruWlL4azp5uucycvmAFf76iztp1rTMvktljm67ovLwOA4C
kzn4esc+o7iJmIOlHmQyUqEFedqemjyhNAenQn3QuTjVkfe0lVv2uH9U56HvbxUjcl9LJKP/HilR
P1wofn+rREjDnvueaO/JhSfgGxFRK60AFosXOUZDa9NZsi1pIUyxxO6VJTWyK4nWalo7cOsYfH3d
tSE6pYs0O9RMpXVTDF7VSNVo6tpzVj4MpNVpLHnzglli7B2MZRsLagkDAqzGiufgD541OjJLTijB
2BiAYDAl3tpRkZ1QQRvHMxpmdG2kDVcGwJ52F+E5aT4yUfzLRSjsbx52EEbMJkDopEYakVJpRbvO
sGepQ3u2/XaUvtsSBATcRfNdtOboKPXo0m4fwid70QhftzESRYWeV/ea7UNS3f9ZSioc3ImZmNwn
r9LySEV5YJnxQ3XR9DY4Ktm8ZjFNJbaKEapQMAQQDJXd/HqSfx972LdO8/G2Ee79pNIeflx89Imx
op86Z90Cygt3C1H9HA6T3FRmT6vjdgOoezgHXSLKLx6JY+1P93TtJJF94IO4LBJkvomtdtmrk30r
jMgE3gWsAeFe9QQuS/fG5oCStc/UhcEVF0ExkloFvb5KcmPF1eRHA6ugKGCcbVP2eyP1VA+y/+xu
IiM3MAsB36xFLrjwAqQT0K6nDJhpWXprUptbVolQrtVFhHbk1Cnkx01Iui4bAeGiyJh8dbCBJTKA
ML/6GTLlsPXUwa2ZS/F+j9LDsOWpPoDLlGCffBIpxYTQwILqJ/oLoascAMvwsY3VNylft1KHYVck
CT5bVMiJQPqAXaaggHhD+bjjLtMcvBwKlmJx0SaBzHRNOGelBb7XDMyhSPAMqOqtXdL1/Hn0TBe7
XQ2DzUSw41mbTHtoPf6K4OBkYkNX60iNu0n4twCH+NDvZb2AFCBw80e9r8WHTJEjf/U/gcKWlsMT
ibg/mw4O2i0PbbFxgPuTR3CGmYv9fPlihoqMC9+ZT4gUHJE2JQgFMVhASUz04LxJ6QpzRxQa+ewS
JjK5b4abPC/TvnOXR+uKhkVKYOyep+0fO0yUF5w11klB4zR4TvxY5JtTuxBSMZHCsbuvfKcK31hg
f3s/vKOwvixKXsjyz2MbUUWwsTHoJRwLDz7dEuDlcEUHUayQAlZ7xHlZwOqrTF+2YGsEKOwehRK0
qW5IG7In+nr0OVMpd+3rs/ftSJc+fcZv2MFqzQL1u3VXijZWvg/tCzOUgSGboNCzkNoF3l/fYa1v
0cMXnPt6oKetDBbBElgMkn0aIk4EiBw1WGfWytODZvJr7m8aMNESCn4iysmST5aiOgSqNMqIfjDU
x+plz3e1sg9L8gnSfgvEo0cZcxn8gYCcYEsnU92CeeLgf5xiqzrF/VsX72H385XaTvO5yfKJVait
XkJlNOc/dc/azguPwkgL4mxiDsAVH4Db8ThReii4Q9XDm2lUDR78yw6m4AXjlY8J3g9dhhkbM1MZ
qQ4ZELT++kQM10qo3ZrdLOv+tGhTyaM+UrLLueIRXOdEfiSOOMvIiwH2nsI18K91+xDQBXo5yZ9S
39MCRHGHZXkNhxUwLJlaNA7IhKhN4O7+UxgECbFw96Ma9iAMLQshutciexmRn2ZRxOct+KfTCkrO
3IMKLWJBa15CEw+UP9jeUBJFCg/ge414mIrZwX61/3QaPuqSyvGPOKI17+KRWDzchihdsVrRFcVf
6cCz//DlwHRq+lve0iXbOge/8lwZHk/tmMzKv8rWSFMJB5pgJV0c/XFJLWTYosEevtOx+PPN+Rv4
zi+Q+RyTTQ/8hRhfu3ReWq7J2fJsP77bMtsYGW82uT3lXlxi07/wtqdR1NTMLLPWYSyRtakGP/Sv
+gSXl7+Xl/tt/S9jb6YSx0poJTBxC6AzfsxkxZPQtzRj4ZBhAgbR6UkU1Rny8Xplt3Zvuexe3uks
BhO7bduFzBfRqGdSOr+zKfuOMsBT08MW9l72fTjxVk0xXoVpdMknj1wVbc37TmnrsLd7abYcteE6
kvJs1XqtGPwOKSceH4NwTWaUdMkDGj63WPEhEwbMocUsA9IPCp7ZaCNcLpyyyjb92ThJPYzwBHdu
6PSFS34fE77cij2GCVU7ooVP3j7UlTRuMSQDLTv/1XAq7esYujEtUJXCnyMWLR7zp10PldSXlSIy
WaKxdOhayROMk/1U75B9sS1osLHhVzZOPGheZxm8hLzIaRPC52bdESn+1+y9J13dbhO6E0t8b8DQ
VNbXNMwbJUwF1uDrN/aakmpJC+tCLdjKhSDAmQ93uBX/6eBANvfKpIERXOVU1VjBuNB5OfAqj6s6
Knk1yCjMgrKXm4wa9ZU5PbSinCwXFubgU26d15v8tze7nHy1dAdD4/FXTsU+qbCIiVb71Ipzm0bo
NvZ9fBxqqFXCB26nXSdsJ6YVmXWF6YDpn55dLIda5hYRm7nVReD392j5HOMBwge3jqryJLAkMN60
PU0ONXtb5jyvQ2r+boZuoo67pxjzs8i35XpqEAr7Ss1zKPBsldNL8rNO+rT3h1Wo+va3ixBVXKNv
cf/O2HyMhY8OHx+8xEzPoapHaNkTAp5HwJkQu/1aXDa6LYHr2oimBkan4glqSKCAjo0ncq/3gyAF
qSbGeT3SbC0LBE/DVMPJUP90t0OK1Bu+6EjXfJGuDg2EaHKoFJO+WXLrTDIGVYx9we0OsuGj7TyX
po1Vo2Ypw5t7e3KSUBMw/Sqqtp+VVt+hTWMEBfx77HCxmvMPmRfZtiDisxcKPbioO4hh51sWb2hq
aTI1UNdsUtXShzL2grWWW7316Qs/1JEvQM/YlQdBI52gP4XJoeZIUMxLoLAZdouxjzgjqIHs/6L6
e35ECoI+ox2g6hR3OdrGoxrO0jkIR2wLCqmx42lwKLJTvIbN5FfSI+oW3L1MaLMgOOvYPOwL6QgX
EX4r17g1UZW05sOUWNO7SK+hDhepKEw2evCD8ydSuTLqykQXet/AsXyxNdNVZN1f57L6nDANq6WS
rwdb/f5sXISUsS8YyLwVL5hOwoQNTH8fpYdZrN4Sh/qmWUBu082BVrqAWZeYlhjxVTZAlkZY7GNd
f1eWJdg40zOPL35XTqrRNuv60DQsjwcQkrQQYu55YJyJhAiZAz1+XjcCMWd279I8evUihoXTv2Yc
jO0djUvBHNdg4om2Y3KJlSW5k0hwLfNc4G7x5UYb0hoaR70VTfWnLDTzQA4uptW4nC4KCb0HWOFj
1olt315B/Gp0gtnt+ssb5xwV9QkKOBQzTiKBqEp5pobF60QjWoRA00qSidD6j/Qk7G1/YA+VjvXA
wHMfwdmAoPQIOr6OyuWxAEIPe/QnAheTEgcb7pMXOqtUx/rcyGc03VZwOKMxr34YzV1YXt5yVBRW
rwhLxCwr1j9k875krqjEf85R2QS0TBsU6RX35vJ+b9wFdBR6YN9EiE67NOUN5YmmtcTWW/eDsMRU
Vq9Tt0fkrzkspz0JlhmlBUKMOdPILnOe7JwNhpnb6N1KTUf7S2BJR6se0aouUvo+Pd54WrCotYr9
CVsU0m2swBWH7asVVCrX6AfMumVscGoB1VqJq245vS8ZPfEcn0gr6P/BwTwcyAaaEBCGAAXnMtyA
eJKK+cKFAYKTuYtxT/AMVA3BBXYMxZU88Urb+y++PTXFvyf64D/nsyDRGDmhgJleQkhEttPNqqRv
OjcCJCgTqTkogNLfqu/1XNf0ftcMZYKUj+FMjVMLPAyaIiotXDniGTMDMac+irFzwNHtr1bm6zIi
0KDftQG1cGIXpfRBh47InrR/4ClnU2ud0S2jc1wHBB445jb00jNEXMfjVonfxw+bLUNNA5sPfQJJ
2CLlUr0rwupPzJVL28SeLdGgXPVWztSW8MmFWvrwnxqse+SH6dhaMf9eH8MWfVEHH23wfq6/Oe8u
XvUj8DkeJo6+EevImu6yC5s/TNW8a4K0ocNnBCCgiPMOuwqML6cHvYTA773Jvrjp5C61BiraaojC
X7B+3O/B9ryv08xKErT+n22Q/3ahNfWpXkUd6PXRCfGmOxCbWIUtCST6fsGIs5k3GpIot3XnOQBh
QkaMHROVMyewDT7HG/v8I0bNIv4It9ljJMnns/WMTjcs52tQe1Nhc0o9qePVJB7H/yxIVXtcQfxu
YAAcXZOFLszg0imY4r2GQp7XUXpVnpXnhBRQZGNHSVWCcqi41X9QpoJzwvA9tosVxW3kiTseFF9G
YjQBIwwi+M8kYO/o0gRvOyQUkY0V+siRqTTGFRmhnAQhqhblr2bMmKsSqJY8345aAZtQ12yMtjCX
oxQ4wXZQr8bCRoqT9BbWUj1lxnKU8XGVfzy+HSwMltb1jOxM9rKhFLoCver5jSgKmU4R2YFpnED/
B9ifNyXGjNbRq3kUSmFeL5Imj/VAs576kc66teFOlyXCMRFfxNYd5+aYKswnxaoC5CDwSlRR+k+D
pw5Rv0tW4nP/Jm8WXmqLbogTpRYpXWFJkPOmnDuewa15j8RMb9zY8M7wiKN2h8jX4wgGKLy1ZEI2
zV+vQXipJRqGICMm/0lQADBLI4EGXani5YCtt/t70dMjqRF1+egw+JDeZDzFP02q7h40URZqDMkg
4J1EoceMYlADOi0IOsZJa/d5S+GSpQ+IWdLow4fRggd3d3UIqQUUDPW7m4F/hQjQnGDRjcWXY1WO
dZU/KbsesKQPNgX5kPGKgLIOFzWHKJSZBnwJlBdQuynFJ6101byabZVwP75eFlX5BWpAiT+SbmOi
5LlWN+TctSEDc0kyOpXsaJnt1zPINNzcndLG8zss1Ma+00ttHLT3c9GejDLqbCfNJlWXA0RcY1cs
+T2MJgPIg/VVjFoxep1GM1SSv6wiowDSP8LV3Y4sBhjv5vzn7/T2Irjv9Y0L0+HbJc0zDkH1iQCh
Z6FHBYiU+X2ZFSIprwbFWaQaELbjo0ylFsp68iCg+1dXEgCVU0hRfsThrN4dk18NBXRYkU5QpuZs
jedPuvyqesKDd18Za8lpqvOaWMv8qIbtJAsgIUTM02RjI6kmjC6cmcjTPfR8eWo8LlUuFN3ue5/u
mXs/ccgsCX8ORJ4KrfmI4x/bcYjnocVAoEP9RSHFVy0Jbux2iPeBwwmdsg4MZStgGNrV0COYLqQH
G/28Tc1HLEq6/tL7oby176LMlV29qtXsuLFsvUjnDX4YiiEdU5Z7pcho2GSOrnggXTpHFEy9OWt+
V+wqdEfLykPVoyQHcEQ0yrDR2KGNYtLhHY2BAMpt3brNjMsi4b8W1qmfRR9+oukeUMn0L4yFYmbi
ieFcA1aF9hSLXzgkaX/IAvLDYsPRpWSiBGkUjf/HujW+3H2JqFYBqWc/IF9qmTotV4VuJnqUP1i6
FeqaEP5Oq415kbAfUOr3IrM+oZNjnz7zTPDf9qfImIAaWK8q0j0l7RWnEExhhE9QXe2wsqudah16
6yW3BfQBNpJ7gLet26ketIIX6I+6zUnOLIsfEFu7G5GwbW9LYJJ/AOE4gKY/8lTDc/bD2PFO7mz7
fER62h4YZFvRT9LB3VVvzKROZ9TcnN7AHu6JLP1HK/p7Ip61hU11j+otsQ4zWXpusOt3yzWpszfe
tNbO0BlFn4Sup+mvXi+fjrWG9fZlrB66s0zm+7OL91GljPkAdNPzZWFj+fmRbV7ZCvgUiH+hcisg
lTiKcn11RopNc3P8dNINHdatI2gRqscR9wDnnvQ36RVfZ35rPlsK6SizJ783GTgV3JMW/WKKf7bs
ApEAA6S6lwZ0U7pkR//bQdOXtADwGlqr9gSq9qUhGnBpIKe6DpjS1Dz2kEFQwvi8AEdHIqb71KNb
epFXezvr6Cxr2w2qsQbaAEK0iu+ZFURj+tCty5wXxYXGWJwcOXvBGvmgj+XltDXKFifxyNFV9U6c
Ggp119COif7+w5i5qDzAMgotlNbyKAipmzI3Qv6SzkkCNL2ljrv4xMcnohxGeE8PTiQrkuZoOb1N
nSdLd7aa3EGPI7BVBkKcIWZRoHacDOKYc/6Y3l045PizyVhjo6CaleLDO1R9AUVolM5JJKTWqBrA
BF6DbymeNn9t2iuEAcLj7eoNZ59TSFm+MgXv2lq+2izI8rRJCq7yWiOxafreV4UzfVx/ANDjKSow
5DNLEuJJhH3EI3x2HHGguqcliyTppoks0LAJRA2YgUjWIQoqYSmW4y4KybrOhyEuDQ/WyXU452e6
kYEugCHnOigN29sau55m5wdF+K9tRCJ4DgOl55ehVRMxk2/bEoCxmHHLlxd6s5FYJufWDsG5RKTd
8WSJO2QeWU4IrGqUKABW1vDizplUaH3L6j70WjScMO3FjuQlJ2hwqrw5jeqBoezWcU7sfv05ijRv
BMHQePmp5sVoWzVLPlaCO+7ritF1iIO9DN8eN254lS50/gH39kYAGDIxTyd2vbUvFoyW0GDEaqKr
dHOYB+DcA/l0lvxR5BY3cChPyFudyDGQNukEZsuV57gD1xpHGpZ13VpbtK7RF3gDm+Pe88cnpKX0
DnMpizfpGYvasOH/fS5AROIQ7zMCkF6XkKLkYBB8yUpyo+8YkgpHJIQtI7THQxd5jYPGuW9aMsBb
qeYlO55UGeBkOPSNnRHQTYGDFGHSbcVHzqg0d+sUXIxy+ZrMu3ojAIvcHl9kDm8mBUKDllEJwkln
wBSdRhYw7xAjUpjNZ1cizXXTnabWIh7gDXcdJp3IkDwHMq95Irtm3mG23pGqPxb1eAWeOL0lDaOa
H1p0NI31gtB9kS5mf6SyJLayxvNilXMnm7w+g6RmaJrznr1okM4OtXxAgGzGKAubYKYuGs4qVo9l
Kep1tgHs9Gc5eNfoh1SU42XQg/jjvw32v8rf5hWM5ClmcR2WLGrPX+DcgJdObSdsMJSnmcEQy7rX
6Ddq3FBqbCjzYu5zO75VCops/m+S3AyuAGG6NI7xEArwbt/xSgxwAur1VBipdvlDZ9hwUK9TDnuO
HNBDKln3nL6KF2GYt9cESGAGYvfCshUb79ACCNczU2G8iqyZAizda+4Kqtm5jTnuxmF/GSIaa1GY
/ZQJE+eifwP9jsrk/GM5v2c6svG2DwjlI5uvUiqRmL3slsKNVb9/U2kod/ISBYF4uIxURfv94Kb5
LDb4NN3j04TqZqE+w5CUMQa7ztUzluDf5TyE8EAv/WwmE7yPI4AKJrWmafT4HYsThUMW+EnQCjNM
8HpCrjHIUYN/E5XIbscOmQfbV2vSEw1xVkxMU39h5XgchPUUJSV5ecGNnT2IO1281Q1iPJy3FQ6e
vyCGE0OaFkBZ+GipkGnVi28wHlT9q1VTG0xw3nDwyCvBz53mnXxy2EsAQhsY6DbNNWdxEcuILP8Z
R3A0dezyVml68PDskl9gxB/+1n7ETw8e95uu43zgRBmY6fXrtQlKDZT/HemefSAHNiwAGCVcaXuf
udl0P4ElSfTjvstk/lwMN1owUCjkzOqOs3z4GlxF8yCn7wSkDP8AViWUtRygZirhcq6+Rhr2ybxY
nf2SVg5pB6YBDupOYOKZNZXewe3Kb92Jg+LGWQRrFLS1RCBoGmapUw6xr8dNKHmxsshaiV1xdAMV
nmmngAfFngm/eCQP5EpvKdDJOC3tbV77Y5iRMdzhtFST8WhN63HWeMGpBri7RktpiqAvK5aQUJKy
rPc0BiO0ygIgeO6qnU7HcvcV/K4ABRlPVAT9q+h25GrVAS0wmeYcZMezTDMJeoh+LIdDfJ+SvZ63
02s/gRkx4HXWRySJM25hOUFVpgc5F+vTK2EWuGAy73lMnLmWfN+mgaHKwq7QJZ9bS9W4/HcSum0w
OYtZRmsv2yKjkqUzi8auVPk6+AUWpWhOGtZ/Qh7X0QDEJrE3fhMLcM+toMjvCaUC7Uvya42UbSJX
OTgTljidFUNEYsg5I08Wt920agX1w+76SnTZK24+u0IPfc8STWdBlTSypEcZ6e7CfbLduRdR5bQU
Ey1GT8XzEiVX3F0RL6goyuBrZBRB8gZ3HFx5AV0iGVuwMVH38mSbqLcHr3Vo7ZeSwyYpbl8QckB0
8usUxEwLqfLU++q4tDVJ+foPj51IToBXAcr6QLmp53FUc6iIKpiLJXVCtDfD0uQ4s1JyJuyjiXU0
rK+9qEoprb3uUrMNRUojuAM6RpLvgcIIa3/UYSqoh8dfiTlEEm8DBDFRVSVS44zAcb9tJuVaTBH6
uFZmK5F3m0FwFPLrKSOre0j4OHsD/oTqfr7mdKCp3/WX5A6KRIKZnbUAzNlaBJx7gwUJveyyDQXh
3IWiRrE0l1LU+epuq+bp/7awel9HjAs3n+2a1//oJ+zh/3Tu1roSR+DVpbc0PlvR2SBsPumhM1DL
4mkbGWKjM6q6k/mBD4PcZt82qZ8c+1Ur4pJFyvhUYpxRzvJyjGtq2qh5fsWkehR7v0u//5yDE++T
cYtjqEtCzhbR5ddVHB/5g1VpmK0y9DrOOy+xBdYt38nKEoGjceIzLHIdw4X3kMUw7Mh6QeLYmolm
w1dVVOBVQCeGa01H/RX4MgEe3qS0krY/+y0oK6ZJ9aggBxkhHavcV+B/EJtXJgwqc48mpKydODY9
PIUytMo7+sMB1VVa/MVEaP2hEVGRZj9uvr0tbQoJuTsAzXNEcnaLCAnYyIR9KtkyBGPXVXu3ijek
fYcq/CbNcjVaZgL/UQjXyLpvkbh4CCGVbCTsZ1XsdM2ilhgVDi8O7jE6KeibGRZiTj4+arw8qFLM
rnDIPp07++SWZZVk/taijw5x6E7CLP+yi8N1XCQ1vWBhY6sRpszaSRKSqx5SjqoR+oaiK+KVqKEZ
wmZJ6EJtoA9mb+3iCbcdl+uqIZnfwQbcalsnA1UjEd2gTlV6lbRcFUp2Uz9JCjv+oyUC3yXARXvQ
p+zl9WUOulJK73Ep6sv9g3uxK58vXP9s1KAUiSQ3+nqDmIy7p3itbHQ8CSNfLLUQ/uZ93ArKfCl5
PCVMaeDqGJRKnK16NAKVDY0NfGE/qegfXp1xLr+K87mu+BSrf9t91WQYXRhtsJwGjQnn+BMtPHOI
GyzkO9WotrTehLDbJq6ounaPnz+gSAwsI75/nnCmZKREn9uijSYCgU68HJPyAAqMK8EjOXS/tY+K
CgBUZz+wf5GXsQPWhb/Mz8sKbcrXbUR36GhxV19AR9Xs/GGvadjDkpvQYyxZdQc+QEan3dUSxwKl
TENs4fjnBmydvXy83ulgJKHNvraai/mUYe2HPgC+3MR1apwlRVct82HDYmfnwSvxY3I1rPD8koLN
KYGxTIPnfWRquDFVfAiWeVGAYGZ1H2vabLf9GsgtJUHoQ8Afr8V8uEknZR/IfCPSHizX64+aqG8u
tbGRwsc+txeCbme0jOqXX2X8KkPT5hig9ijjPMXyZNMHoPFukSnvcXn6rxMK0l2EZNDhFTDTI62+
h6QiG/WEq70jeJldeBoxTq/lJZH/riIX8Wwv/bLAi1uNzF/u2d7+c0vR9WoRHXwdYCVNfc6mBvPN
C1oCQbAkcZ8w+7vjwMyj4cxtTckXG5OU1XZQGzawR5vEjS4FNQAq6l2cY0Ju8jcc+UQGjDrmblhK
dhSfmBe8Bb0jkL9ywVwYAwPo/LiYJueEvmTEMSPUSTdwywQYga3nkwRLwMDVrDWQMt4knusU+won
tAzW9phio/JQRJdK0opKlJlc4iz7rU3BfP5lU30LC5x2WCopSf6YtJy3UcJ4NgQxW+PiqcTZMJvE
EAIeDax0N/y1+G33+l5Hrr3FPGLp3BHa76I1lGhTDYQNTBINi0/LCz7qOLRFha4eC/FL8F6onKoj
tPmBO3dNnPXxTEJA7i1jYogwdhxW1PmDe3TPY7zacpaD31gnZ8NmJG71DD3h6ewIcgZezoE2Bmzm
urcs5Z6IAYDb8SnrArAkueEzsfawheFWufvYzca/hbM8++J2eJlEvf16sJkGMDWA1z6nnJ00M9tZ
nnAi5/MXFjlNT2w2UcBD6sdYkJ0+hJaIfxuropCbSDjeFLeZnTF0ZUICSZCEGg7o5coVZQsPaAdF
NhhJ9oXzPqVgwphBnu0ntHM/2Vhz1wYCBz7eZ7IoxqYOyLoFP8cbD/KJjckBRnplf3JeRV/bRrgA
CZ+i9E5NrD4bcatZgQTwnHibRrZ3LM2cgh2WDyK6z0lDA3/4qhuEhzeVqV3dBoDRFj7C6galYxSy
k8uI7S3c6d9RGP2X51tMw48GW/lB//+JD/7nzEouBzdnwkC0cOH6DRYhP0typaFU/61n2d3nQUL8
KZBEEd81ZOnx3husxI5zHW8Dw77BX00QRIL6AmXegrW+vMx/huRef0Be2XZMFiubqHGW+SKXgwlP
sz2Ssrb1ZWkETpSE2EMoB/IuthqG8V6rS0F6skGspiQFTLxveYs8jYASpsIYjQIeOaZ6NqIrQt1G
ZgcbvZ6vnxGJbbLvdnkZjekU98kQz2jsJycmnGdIy+DFC1z3MtBin6XEMc18M5BIfE3iN8ja8VRh
IqftjWxbQS8PVOC3Fx0zSTZIxQBfuzEEaiWRLIl/BYcHTL+nxrhwc03vnaO/e7s90S4IVibFF4Ya
JIsGqmysaMlfFw+hS9KvSPEHbRIpKB6z/3KjXxXPpBuowMG/jK2ligRtbuFsgYWGTnPwAXIo9+UY
ovtQybt8jSUnjBIao0jkYnQv707uyb8RPn/0mmxtjF4jOJUhQ8lZ77ko4ITHDBk9lgBjzEu8h9qo
4gcR5/Ou6uJSYQ9Oi556tPbVGWsO7Or7vzMcNt57vexmKPKn/HhPPEnbs2c+Jp4+QVu4PsIyQ1mt
xDAeacD+hXgyus3xYpLAKBqhBkBQw4GMiSxaShVZcd5hDEUeAbFJbFRccKm6/66GFLbr2WB5RKsC
r+Oba1is8G7Oz97BJIw2HneALyLk4raRFkTzk+6f3e3s+QBX0rk9TE9yeqXBQviV096OphHchKfU
K71HkuzC+/Y0n7vnjp1aV0LhAZmUslZG7ggDtZqQaB2Y4ZG1le/ilCyEKp5k0T3yIUf0w+PitYIp
zsaKKAFB4hYe34UZgjMLM3FptiGSB75G+OPf8s/WXd6z3TVSoZwAsJPfX7zDdGm6IlO7csMDeuOa
FFeGjKKBY+f0Iji/tAS1bBNcG6oau1lzIo6Ua2oL+AyFtEQHiGjp92zr8JqWmYqEtmzj2I3GG4FG
VkAXR5+y4f32YlAsKrlWL+jI0AvFfNplkKQC30fOtKbDvZJXbMhAVmRw09sV61pbKehoy5veQM9v
Nk3IkzNJYqgrIdmI1OPalYOPUQiVOaFhqhqrWDk+H+O+vy6GkkaOwvCzKV50CZuJBJ6R7N1fzXsC
2DXvU2gfPKSpwoie7HgrdRqmKHvJtP80W2Iv7YyiD0Zt3RGkSEGdKUlJIM8QurMzXPuGyIGN7ghJ
t9qpYn+7xUeH7UolSE9Tgs9I616M+cs9GUNNV+is/hPpdDucW9isLyEe2WGs0z631wEW7iWlzhTX
BiMPn8cGXVZSx6v3vFMzcHVkwPjrj8qn0cMicCuyXsTG0vqHCE/mNXr9PXH54D7S/S2+vF0Qe8JI
WqI4R6FuUcYC6gvu5uesa4P2EAwLa3eivBazSMS8NB7Wj//K6v+bpvGOlrm0OTOGJwDsKPVEblmj
i5wGu0sBinRXpM2/5g4DVh9+EK3TTLZq1wHff7mdTHHN/gAwHekQyOLuL5K+AaiqPpGafR+GljK1
eK5Ra9sOPaljCqwAEp8nasX/kRoLmC/bSTktYZXb82UO+EHD5wOktTKR4naRHB0MdmH8ZFeYXNA2
80Y1hCo2u2YlfdVeK/0Ku0wOFHbS2FDy7WqWHTloJsGOKFBcgF/cmyNMIIP4mcc10PPyxHXpWIV8
LnsiHqNkM5F4veZWgX3uwvDe9PF0I6ARxSORPcwkeCSgFFE1DXdUqJM2uHoCqVYj/yv6FF4p3L0v
LCJU/J35SvHLyGT1PGAjPjBgFf60X6rDq8oyslD+0bhuD0x6/O9On/gSSmMpcSfEv1ZP3bONlape
N1U+IF4YeKOBR5SJwxJrCOQ0dpd7vAlao0BOr5N4tb7Lz+RQxEkYSaV6lH1g7OHX5BeFaWDxo5JY
Q9XgvzwR6KBlTBB2SN/fw4os+j8A+Buj7xVM8TTA0HVKAz5X4YWaE6GiFVNRTg3nQ7bPoi+c7tM3
ZZUazaNHdbcH7+c1yWoqmFbg0/2PFhDK0TyXItmIAfaYHWhtE/CNE323xVKtsKh4MDkf0j5ZD5fR
d9um1oeo12jqSTJZbCVJx3ixmv/6EMtsK3sDz6L1qN3LG0McXuGqA19qIBiY0OeH/dJJKKbVgjns
jrA13wCvwIHHSGv54Dwcutr/0sz4McZfdK6mj/+5GY9vxpQn+7uOO/YWDrNLKVrRDMrK60Ir25bX
4TQL/SdbeqzdMbWE6eIKn1G+zAc3NNbHyiP2ER+q859dTSTvnbSh6Wlm4xLt+ekpH0LUDMfmt/ze
092lBVP4juJGtLj+APpMOwMQodFdlv/bLG1oIkCHvJL2VWHgv+5Cq4V93nVfhHv+XiuxKucL3tAL
sFY1jKeH1fNE1Ryd7hPTN0M9xet+GKRQ4KcPGQplGVQokmIky64EtS75B1ZouDwS6yK6Cowqz4kw
HBAIQcfJbE9knLQ4m/4WVnsPJzeNglTcsGbPyPgjxbZJjzmg2Z5iTDOCybOl+WdGvvFMQNUCaGsR
m+aD2QKdagmE1MiIRWYZMdemD8zR5fvUiDhCGrC/1egsL+BODXH1xBj13i2L2J5hMQRfzRvy36XG
dLP1ayvQX4o5+86ILW1v8KDAL7uSjCXTO8hj7uO5HgdVVlBJIBOvO1eo8Zgdl65hMbUXZvbIUArq
/baYD75o/7Ir8EkxOxFQSrJ5Iie9TURR95pnCTk+npAguNTG41V0Fn4KYp4oUjyaIKTIoFgnNLQH
1PXjJ/j4rqxWlFTCsODeJ0whB6u3od9W9W0rPntnboWnrn9a4LYUQ2Er9+tXic7wDoivC4NEqYWo
Vy3km3lzJ5sdUYtVjTIVa1J5bjintErd3woCmg+hCV9gFMWzKNQyTt82tDowpUJPCNmOWwNsBTMC
SCfIZAu4ny8RJXBP/CTJr1/XHjeJiDlIHGd6MhaG97RosQPOb75ATGrholpPf3O7Da7vLYnM7bov
jlz1HYkdgJuQK4k+Qn4zXxWjTMUv0wlfZwRtrviCyRbgBv991XeVdWhIOIGu3ltpaXHlipdST931
wr6AuH1B1Hz5QnqUoQVD68mHTKBCBKdJYIT0bZmsQgC7pXfE5j/r4jLTVhXsBZHsDvHmNPGlLJ9W
cF76RPcs/5In6wLAIq3ksvXJayCR2f6r0e9PUzqeffoZ1ALEp39OQ2cgwG9bRK2QnmUCEBk+7CjX
ZSmt1uUq9JbFYpt7le4IlGmPh0rG61hkRfxpmdPxEUXkGTgO5iX/bwPfH1ZwbHK5+uDCISPAEL5R
EVUsO1NjPifv7tCKD7Ma2UOMEK3slRPtFs/l3gPoVmi1gIZchwUJiE/R4iA3wKQfsf5RY7/B6jx+
heWn2Smi5+0Z9zvYLgiB1dW080rGfPZ0+FW4OTJxx+9v5FoX/vyCtprVZJD0yPfhPbYSlRnDSqFO
jHItC0TvTuzo1BTah4OFCwAfjzIWI/BbwYxMDaw+CapTMa06lx8+Nkadb3xa6T/pIgeAiH1v8DNV
EgsKkJ/myTXLZ3voHxa69TpMRREIw1eeW06626L/H6n0c9pwSbTfhSn/wMABELPxaY1UwQX9QJf5
HTSM8Aw9FunxxgKq9LPU62qKq24K9kSFBv2PYqFXoo/J0KveyOM1yhYAXNAHDCRsCfk1K3WbBh+j
Ch8Hq+VtJdcn0Nok62odjTWhrPDXm4lG2BRsr5s0OymD550mz/u8mljJUUstCGxjiTYVfKHmCmTs
PSH6n6GFbH7Uw3rD9dV4D/bLiUxLUgRF4wtx3vJiC9ZKgn5bifEo2pmL+eys8rHzeA2m+wwlWiIP
MD/HdveTIHEXu4pZ4Wylab7ftxqtndzkozoyFWWHWj9xVhmt/ZLcCuiDjIYCO5ch/TVsdQK/jMR6
N4usCdihAKndGKLSTRdaj7IeZ0B4NRUxww4HZnhlQ6UZSXzTIFL8TOPgF9Kc7QAC0HCLki8ql5Tg
oSHTSMHohFJj8j1ZSDYmxG8acd4shHFL755ixarMpvG3qI4AasnNahVKDCCASvTeN4PaP03AavGQ
przHO+yfkfEMvSvxu2WDFhG/u/pbQ6txLkMuXgIFgdmSRxMZS6/1iKTqMGgWrNAsS479PYtRvBB3
edR/Cj+0ek03CNmQHQZZDBdzGj3Dvk+kGnbPNfsGDNZH7DPAWVCkEaQKd3GrfmBznx3eCGizviKu
QWwpXXr/4doSZJFHNyGjgcYKy3sFo8fLtFnqNi/uUVsDUhXboqn2n888dOM3lNC0treIVg52fRl6
R9ZH9vuiFcqqOwXCQNnUiPae4BtChZFHX9u6Qdo8hmZD6+sp0FqVxA8WPjyzusiwDul/PE2Q9rta
cFSVGBCx4KPiCge34P3ivFZWzcwVsM6c7ddVyT4//2RLsZWL/79RJcH9uUa95sq1NQAZZutLWvMe
L0y/hCu5+NINRXju/UEATcEvJW2I66MS4B97pDxKpXwO0/GWzczvEjs72sSuVaotjEXhPRTKMMBo
SqKOQQW8dmkaaEHZAaMqVKNG5xIPQ+qcoo+tIiFSiigrobY7PWpCDVPRCRxAyemDygzXrag9Sm+y
leh6eGdmZFOjhiLX/zPdv5FUSvuJQUaiDHXTGdJ6FkWOdn7Y3xmHOwtmmnbSi9yplbaZiNZRVYcN
CVcL5ZtZRLITrfBk6g6nnTv1cZDlVVoiuKb0sdgdtUk8LVWKQ/3bgw0yM5zzvYVQu+uYnZ4QGtQo
kz52KqYpZwNRC0ExP7zsdC1rnEASbFr2miLqZMtVmFRTrE4eWTsG3pLXJg+zadFktHW3rMMq9SkA
WdJycauZ2m9h3s76xTKrmNX1eWpxa09LoB34SAvUQvL465eJJ7xXlpBrwH4VJqInD7tZN5/L8Gp8
lEELhnMdUMtBGrHn7GG4tg/sU1NEkzxje+csq4V7Qc8apNP6uVsiUNYYHYcVSH5XwDgkYNWkv2kS
Vo4rWfXmrw7wG/6Ix5Zgi39KJvm2bPUH/RHIoNiSIY9LOkMWuIgnIC1XQx8Ty0u931O4/lBkJlw5
1pOPmDqRVPpzaBD6tuI0Rn9zbClw6dwojjh7IIuyPWNWTpvimzBtKUSl0NDSZDOp3JyiX4wpVReD
8UfQYqpY7GYIqjKEuB0S64p50y9TxOmIBheu4udrlcaBOzqG9BtroNC4Fbwv69xDRMuZjulpk6TS
Yu2h/8xtZ3LzyFlbBkG9De156Mc/Gkrc5OIgyIK7W1UgDkbVlzGcMuSeKSphWaoj7oJpgpvfVAVQ
6dKsfg4+/Rl3OeIaKJYUVZ+ePODS+k188E9gJkwAKLkK5+x8Y3vRiWk8btxmW5+TU2rev5DzZHCG
YSapEUadLL3GMHkMpa13U2CW07zCrWunCDh7F4VRdF8IQlF118OBCTylGGhKPvmoEf8rR3ZfJyee
y/HhHk5J3Nfi6lhN89Spdqq8g9pc50tnWGOw3wkvgUxk0U2HibBefkIk7NM99l7uKHSoUPex8rDj
lZTIaXAEpy11ah94kjC96K+cO9Kv2FlLssvpumfVqXOTAJfypU2ERlPr3pb9TqVEuhL0xMAFFviW
zuEZi5+8dovi0bypz3j2m93GjdT4J6ON4mr88oPZ1EzVepgYOAF69yRsS7P5TgjgWt89zmqK0kVv
3sSk1q0gmsqt2aluI5wH0C3jYwwuYTLZ5dUaIgXuYPQnYat8qKU7gBnwE5lchJfjXkG7K1cOhVkv
4ak28OPSLAalF/D4poU8p5cxPajzwjOKPrC/zVa0k11DRnTa9Hbi4zy7i2DLG42FKoyfojnkU2RO
wmrUDmUYXvzpdGVwWA6Kf2aXLdtSzmBqD4+dh1XzYETwtTmMJ8b12UESkSukNLWAMzPh29A0IVi/
0qD2DHcQDzI7puRaYGoCqVZwboGyQuC8+smEx4l30odzkG1jKPsNEtx07bx1DjpDfwZy+t4untll
UJXhpwI09nZthbN7IMXqg6+5hs+KBvsa/NGO+wzm938+iT4Xy7An3uDVHc3Nee0EGcXEgVGYYKcV
KVLslwKnecZkn+hUsWNBhkEXGeC48MZyMnBaWNdonMd/E/GhnA2X3ds0XgVZcwuYB+/XJjp2Em+e
KDH+3eymluPMBGKhYOvabywXJLNv+7imDRvNTK2yzc+eCPuSYsw+GcPiatnIBcIa54mPOfAgMsWQ
cd3jS1vkAZjVZYAxS4lP45InZrjd7UIwTN3eiy9ZOqH6sPzBAjYNms9ae3m+n5aiqJyqSRqurVQD
IEVzy/6GsvTPGetvPFiotmRdLISHKdc/W9jL9UNOSU6soHt3SUg+3RKvDyThtKBpq+cEQPb/YGQa
JmAb6BHmbcBNyHvaEvYLbDv3/hi7G7YIOMnOb4cUCxCCbr77KYzHoLT/Q65hWMSIfk4QKqtrAaNi
xavucreIvEZOJ7dhlo5AbvyAO7JIFl1f0k/mnMTq2xCBSnH7wbrawNdM5Vuj6UPmwnSUwEj8+wN0
sYLuFDQ6E+BAg8FuAsfKf0jbEckP70du+6HEXI7m3yXzwKB4KP85YauCxMl7Iq2VO3TdUrVFGsqB
nLWjPfFuWWMrTvirTLLO3xQ2jndsRPbw+OUrBgfwgttlP5flGxilbMfY/5VRBAhJZ73J+T+aXYG6
kzpN9FNjp3edYXNBODs5omkkmIt5HaDeY30EGIi9O1IWzueN12e2ZDhpCnMmJ0BvyzjSs61xIdyv
wsh9a1NqzfsnMVrdaw+EJYcHDOR23q6ES909Wiat1krDpKMYIg36/AIKDCWNblNIqIEAcJuj5t4k
PsB7g9tkVcmhdkqretjFVxNcMkkZHyh8gLIf/BMPeTyCCSufDERT66Epu6o1PmazuNjyZAMtzZri
UKpaoSQPJBWjKYRZffCWl/ygA9Lw9HmQytxWB5LrwkCihDI5VemMVxtDMqzofncrYxzJ7lS2TMYF
IYIg+gTP/OidRKEvGYoX/DWVciTmNC1W1ogEkFq57w9CkBhz9jkrs5yNd/BcNF1ZKWPoy7wmTGkD
gR9HQ28FXtvlU+WzE74j+YeL7W/gfR956Fn4f6/5yfB6xTH0L50tzTuHiyVB2/Ufqvb97smJZXU8
/xnbH4JVQ9leset40ODpqf0Hn9JYl8xli22FRUJbZfxBU0XKDrMZC8hKxVgaMHMDSW7vuu4BOZ5/
p4VRJrzNMyGOzDcrCEblMQmBoKr5kcLJEowJAX/ovMPStucW7cYPi5pj3weWqVd+BOn0xnqfwSbm
B74gWsfofZExle15WbrAh0PIR+VHegHun3R1stXM2mEiOiH51reG1vUhfeD0riKgdyuoCd+360j1
KnBUVVL6OtWG/P6vMIYdiKJ5S/ZLobHfR7/qDRz6RIagPT2M14sIGoyHFdNWnjeRdM1SyUOUUJCT
URnTtt4XaVbZgpmhQnhfqL2M64EHcSTLqMGpBygGqw+PSLgXwbOHfdmYNkx6DNNIE0K28hZ8DcVQ
foBd0sMDG8erSwUft0MW7ve5Cjyn40YM+114AmqS34OaaQj7EaZ9gahCbIoA8uemAOr6UFiSKgf9
We0oexcXvn5yajYzmZUH2mavcjR0nCUesAYZeHv7sphwd+e57x+W5o+KJ7sQlPGGQQPhRFb1CvmS
5WIfeaTK8/P+noYW19Ks6PwyyYWWS67Mhb16xpTICABN7IvNNL/wOOHPikmJlrlurJOmUbJdITMv
EDV65sgwGLIBA6ArVA16KUP1EjMm/11GeG1VWZMAW3uqtm+6i0cP0LCp5OigG3UWGsM0IDnZa8My
oJATDn8AQ1aHyvLqQFu21ZsKMl45Sfq18sw0e4Vq26xIiUkp1x8wB8fDahyzktCar75QjL5979Vw
Ca+P2OMowsib+1cN4J+eOs15NWa+DYtjNZ85ysMBXZhP3D5UMUJ8f6QaM8gxZjQHNeODBIehht9P
XAVfj/AlocwGK2AXr72pW/+4Nd0EYOFIGkfIzGIy5dmNzBaEUe1isNxZ0+7A5h2hIA6RS1c8G8CB
YBOGaisc6b8WInyLvzVOsiUB+YhjLPUWvod4Axs/QpSWot1t3WiB2iCJ63vhMF6v3gl/BwrSlYoo
LgsNEuqAaO8PnfETxzZ0CSSzDIwzxtnioWKoUABblYXHAtCg1N8Kx4IQTS159k8/TURDCK08YJwx
/KFu+pP9wmI52woP8uTA9t3Cj4PfV6znZSTWu5YHl5WQ4woTEDQ2d0yim/4nAWxxNkAh5Gptf9pk
MxBc/S0z2g+/Firx1+EkZqV9z6FWlY0CJ2ZtqitumiLY1ugyoLMcyXG46xcq/hYO077MF49sUrA9
JloULoXsN3xdVg7bfttM/68bac8EGh9dcX/MISMZDuLYOlU+BUoCqftGwlTjPofNPJ3bRFOuRbPj
NNfUA9AyNcWI4JqUZ3eSaeefgsqlAdPRLilsLOCnnr8kvFuNYG4Bzg4+Xye8tvsFQrERPC+kDDgK
Sn8wKE9Hpyo1PamV+jv5/XuJ8BISml8IDBAYmjJ0xSpQG/eV113cze1RKsuTmbtPNLceOcFVfrY9
1u7bHcGNQHW6XpbQYgYwixSdJSKv0toIGo+4h/wXWDUUPI4joVeKDiTcIc1/Fr5C6V8+LYiiqBne
SRq+eeeQzElNd0eV4qCWfXWK6CZDqQBcxqi2QSG8/kll/Q/IAj9lagPD9wSo3K18lv+Ze2gj9MAL
mkK0sJOT1/PDl9XLqzJOG4mtBzSMbXhMTqoBA3EKX0aiNMyW0xX+AKkIOQOIP80EXP/MGhgGveOF
y7Zt5Mgu/49BfWBj+mhS/lYgBFFpdV5k2u/+u+DycDioPIQ3f6iNdW5QFy/aUkxEUEY/FLrFb3Bz
f93IW+W1Ft4WHve/TdVnzCFhPsp42LR4vN++HHNS6oPD3pQ2+3aeQ5BanoaQROE3/+uVsOb9uOm7
KtSQ1mDJn/0ae01S+btyIhDnxEOLWqa+NE2eOwVE/xHGGWYtHOJGqjhCHeSlS2njdFOO/4uR2i1G
bPHMbphuT1LsvQYAiFwfP6f2rCzNyaLX2nzWF16EDsPJ4hG8mBzEymUftnLmDrb7hD8gZWY6yxfM
pAojlPugnD+jN9+enYHX9jjnQR77avut8Ur8Ko2wCT8QXswxFQk2uuxtMFFoyLaL/fdaO4pyRqiR
l9LYpA22mbPq/hMN4giIKcJYY4FOT+t+vy6abNqkwPsVero1RIVQX5c6dBUIxSe/ZBfdjRIswvjR
+w1q9sh9V46H3Y6hZRLQCTpbrI/DIQN5dHa5QBH0GD8YJ93ZUv6iY/EcEpfhhrZaZNOyGwnW3wrl
Rk3cgGJv7XwwbwpPDmEKg7Kzb2lasjCIqoNIYBREpmVMtUTwp3CPX6I7eSlin9VBBTz0knmXN6w2
6ya5ltVN1xaBIxBSQG6RMMQMg3MTvo1+jD3FGTAUwm0AScjmVg9yAdZJEtxKPeW3C3tqjhQmClh9
+GXj2J1gNZlqTmSUOsqz+/o2XXhikjOxVFWZ4QdjsNw2fUTt+WAA3iPbcpxiqmVlQ9wCDv1Vr17y
28eVxEQu1qg6mas0Mxt3JxMqmwmo5OXOptEvrX4UTf/9NeQO2e8J8SBPPfkqmvywZTFHFe6jARbM
Q3prYdfPG5nVhOrEVNPBP8/DuQI5UsQjtO5PvmvCwLQa2/H93s8bKmj0GOW71q56WsJsXxo3179p
Sd13hyOFQo1apWzYjr7NTKvg8nIpsUv369WOn2OyOlXFffnVSR+QVdT9+hnxiWczs9Yqmj+JlljQ
FBlmuLKKcnS4miLrE2KrqQj2AzsJ7nsNJ2MFxNBLMasOHdgFqOC6NqJqqYXLoJQe0Tq/QqTu6Otf
ZnlKQ8ZbZsJJTLx32eYud9Y0lvHdESkra1JQkCCEdoQSE4VAtZ42kn4/JflveDK2Mu1jIWdAKvQ3
mdzBeCW5J9qqd1Y12smP5aRMrLDlZxbtrnqhI07wHpn0Y8ZrAkSf6AsjYIy8u4Afr7waQ9/wnWeu
y9E/eD+kG805o7781DlGpa0HjMf1AMZDCvxVytNpz1fDoiJKUrQ7oven/puk0eOxKZtEMVLdhMAR
c7WXVq99Vr6BQTcByh5Q4iQ4M/tTmuRNNqAm/LMUGb8zScmF8s39MuIkHmUMEAr96B33z6+E/gXr
4bNRacTpEj3dvzyXS0Du1Yx+qRxc3f5EAK0F49V78FFqAerr63/h3Ycro2WGT881MxVZWzBP93kY
SXeD7Mdvi+fRxEOdPD+DtExb3ZR9hIyl4rPzxqLjT6yIHLK1HghZJG7yMO8PCDp/frmsKmPwqy8d
WxeLriDGF+fKaHnqUDiYbEop9LQ/L67IPOAwcx76gTa6W1ywnfDbzNuhHVhW/lHb39BYJbE6vBo9
xYQOZ0A3NxWyc/JQ12501xt/PbTNcFQptb/XXx5cJXPiOEor77NLfn0OIk42nWMEdgpG2+gvRCG6
aRfM+izcNejjUD6zlNT7IhCXTzA64X2kiULXKpnIQjpzBUsoCSvjU1a0ZvnsdFjRzYizgJXhH/ML
JfnE5ngM5FZ/x2cY1THFlbk18ukzYBEcJCILt1+4znjvZqHqJMc1+T9iqXreUq468tACpl4JHh/g
wITtfyZ/5mgcyPkTgcSPrx6nH5/hu31VRKB0RlV4w6JRXQOGE8wf3NMVG+zpa/iTsEf9kVwdgdfa
ojTNWMshyj2C0u1foq/UAjKcRb0VT11mHNBvV2jx5H0lZBdMCze/ofPHW9ywSI31ItMwiB8XWl3u
H4HxbILlTzRBBBbd71sZiGclrCf5bYSe364brx9VG+P2A1jvnuEbT/09wILqCHaNQ4bBUKWZ615F
/cpaXpTQrwYKq5NzHC+5IrHRXcUMxlKKEdAsYFfQVhkyrFyXOF4ZPKcrhyzLZMaId1t2MFkLXpHg
8yBv7+56TYPLyo4Zq7O+Vz5hiyiEthPPrb4dEXxkVfgj+U6wdPufdTc/XFfhlNhOZaHhNEac7zD7
2LF9qpymtd1oFG4mPLcRst4PQZpFpiLa3dAXWTNU0DIX9TKJ2y0zg1DihKgOhxp+QLCZ/RPS5vSY
mhHLsQ04fc2/Vt16adLNw+fTisdWDDOHi72O3nM+di2dhl0Dr/lW6b939OeG1bq35DFhr5KLEHXH
LA7CvjJhMvLMD7Y1VbNQIC20Mbctw5pT+6TCfjKU/WactYcwu9HfVkHSwNL3A71NGdiPmLqz+UXJ
MSjprbrwNDBplDIwFIZeMl2yNNn/EYv+WO0eAOHar3GqbkGwVBZlNjP0x8oGmLXp8Tbg0ZO4KcCl
uMFTQKVvnMhhhDznKqHrl1NEsfNB9Tzcn/BGo8uQX80PuCz3FkhZ/xk88JZvrCqOIpD5158veWLk
gl5MRxZjtIEkh/+I6TKkaCtW6N3Lgbly9DWBlwvqrhXIVsnuxAlCTToham17iJmdpCfS3yBQY37/
Nc1dA/ybHvnlxCBnXHgiZCGb/64nAJVcgFna+XQk2IveDrOyzXiIDDGxxKdbiGXzB3cExMV4wOSm
1LoQtRBrFvcc0P84G3F71M18tjoc4j1VVLbrTwFO7lTzCRT/4HA/Aji9lWWL5+9kqPB+1BXPrPg7
tx+0xOeUoNIoF4i5BCIiT6ogiLLdTM1O8t5uP6Xgai+3FCU2Ei9FinQg/491yCDMt3q6o8I2/dA1
z7aoS8sJR/tKr3V8EsUx2ZF3D5tKikNec54o9zkhmuexrkN4hcmT0JZLXuGPNG7IEX1SeBiFYGHe
mwdSB/AzNLmQHqFj2XCahyRSUCEpb7Gee3mWHa43HQ1pcoDVh3vAm38tldzPBsfHX6eiqjJJm1OY
K52rDC97eZs8rrLMHt8oTH/JLvcsbtk6WLp9segvgduJIXufUVwOXSDQIsopKi0oSkMEhDCuoL3b
vBNhyaHi64IoueWoLBNWZEL1qWl7xc9coYHtzL2f1kk9JkYrnsV4g2AMkI427OloiYZi0a8qqDRA
rGpJdCMNaccjdKNyTp0BKLsBkTnKTxRP0uB1ba/fTs5Y4Gd9Slf//8dZBwVedPsUp2tm0F4Dy1tO
CiNDVM9KtYQVDEC8mhRJOwYYDW/TIz5b/E8C1mIerLuQVU84bScilDhjgC+DMxgiOJA+iV469qQe
mQMZJga0hBjcYtQ53qOGgcScIazNhHraOAr91rGGD6kYL62OMTGfEF3MBGfehf7zCjHkmcrG+Nlf
lwYWanrm8ovT4WJnISdSbAs9j8Vkzj3IH7xuaOWTita2yNmjcsKuIf76nwPFh4sKncGjqQmF76qx
VuBNv4PkhBjdvNWzg0zloxlKrZof0ToxTex/oQ/QmBFetjSHiwncbwbSZAx1hqV7FHkEvUDqFwsJ
5mrHJlGL+l3k7HbdD2xGv8J9hKG8Ga0YYz36NDk4K5twTs6s8nwKJDw6/ww8LkwalVuXltIY+iG1
O8JveSPZazhPT/cxqdZT0ka6G/xJ+xeDn43WHYAKSCDyjZ3dnK2rpHhFZQESY0PtkwYnUJWSN8JC
IOcIeU0JbFtbNk7uhDiMQxdC8byAspYulRXqETsXSk3rhV7lQWYDLrFgxbrhNs4ok2WWFk1O3cT3
fyybBfsaIPnYL7lMUQAkVaEYATOtWLPhCp8GQiNnxt2pAk3IuRSpJGyikw6PtFlirNdYBYCL4iHy
N7TfEgsZ58hLsK4FQHEubzI12VKR4Npe+1Bwejo16v1vLO8YoTOC8KB9K/JgTWCJ5+eWI5mCk0yO
mcCY3X3MELTNuHsKVPcNs1cBZlid5GZU9v77LLqXEEflq6Pg38Q3G+x2xabLv8gBRBEzZJjy43A8
lWOb/OHLFPG16RtBL6bs40sgqAzdVfzIMd6YJKaojTW9nA+9G57GFmxWKsrm1nPgXVEPCIBvw7iu
kVPqoOnQorOfxV854H2jP07UHKuYMLc5CWDRxFvAwfZm96drBZE3sU8cbkSoV2pGNXtfHokvqzaz
XSQz/2PfOIlM5KKQKVZUZy2Z1ZuMl/kyLdqd+HddKAvNybiVIm0mxFJGUuID9GCYh+tqGNX87N9s
2LfbmwpglQB+Gm5YSY+E7PMbn5+h/h+9P1m3V/piiUoctW1OpNXTua8dA21OvqTiRXI4qFNKkCWF
0VJPOwSQqnn+1YnT4Z7twU0UZow7612F3chBQLGW54s2i1wyguudzvotb5CLOPOVaWssZF+FvSjX
V2v38oQyOGWs/3LRxfb3xyEOTDUaMeIsTgYKR2R2ViED84JwtrdrT/nRnHvCv2oEsHSrdcdKvOV+
y1HxKvvlab1lRXEJ+cOrob2YP0/uMDPAvhrrMUaS21b5fZHb/FlEFqwRSnzYwRZjSk/ux6yNgWw4
ocdbCbXWJwSfBpjah+v2ko7LS+/gb++VayrEw7SbKiJCdRSy1d/QWY1LZauK1IEJSIS8k72aUW/J
usppUFmO85ZxxtFxvCR8r4m0xBwcECNFKgFvEPu++wr+4n+IdNtdy7llqZPdbQodgEDHY6SMxFiK
5Qj6XYVLrEU7fAZFLaSiWCU87LNAc17peB5pPtUEAe6UAe9PrvraT1aNdxP/XZft6kR+WOpuRnkx
6mF5zHpTg2kpy8Ii6zYydqG+xpdxkWe6pYRl4hprRKZQILJsrPURn7ihj6ZaVK+i+jIPbUF8pBY6
2A+8+HW50NdQTeuK1Fkyc/ChymWtIkCSKdKsAjxogq1sXUgBzjEdafrazKUFaAloSj8LYpFqXb+L
an6tMAr7lnyB3T110CyzrIFLgDojm+mZCIrGKK7e+FQx8ZMFUIO02xDeUyQLbTfiDYYSKenGlJlP
8LaNQSBEsXdWZD8mwHF9I1Ylqx86eZes1KJ/RbPnQSSs+iyl2jDTcKBsthgUCy9o2zjQkkRSYrbl
kGBKuBw4lMSKaDcf2sJdIrv4K4IG0I9vRHLW4F4KDH48K7Dq0a9hzRcm4uDpewd7Rpj2OxTBZ/gT
9ONWcs4ivsBbnUMfzD6mbE/Ifs3Ezy0GMWtBw3T/kmygNCQl1cFZo3dC3Kbyffiad+GdLkcXWxn9
lok4AXzoEneXsHFj6c9xMosknCTd88hXxgMkCbe7cbrTFmLWugTb451DSHNO/k66LrvDh+BEBNSU
MRofJOpL/d633dH9ms2hyWDpukTH5Q+EyiRWTQ0IX7F5HHPz5mxvJH1JaJ3FVDxJT266/8ouO85d
Wzag5EDGzwa6Osnpr89BuMumIMYpYBPb1aNFuWf3vtXVL8Twa9XTLmrh75q5j6668TjbW+VamNVX
rscRpcjNn1JHjJDIL4hfvzoYuc+57lBXEC2g0aadELMDkaWC1c+KE6h4CBe4QmEgqdbT33ZWXYQA
CBo8mdxuZcGzqNZMdldq8VrAUPRY3WZNYjd9trzVkxk9aPDnV2Z7+ly9/N/PWxUgWwPvj1sCHSUL
0NlG7+1Yr5n8bfq1HhIiTFFPt9WwstpgnZ4jrLdj8WxHY6XTF6n0zYEe4SIxmlojBPitOfVc9XP9
vIL/nNYRG3v00Iz77vEYBwbyp+MTtgUNSZgBh7dQQWHe7mq7oKkQw8lpA6XtpJvFpuGnOFP+tCE6
W404P8v/35wRYNB8PGjqGZut+hu3v0LEhdxst0QBLClFLEcXT1P2C56TU8wyN4qBU5t/geL6wMKA
WQOSw66TGtRqAJtVhLAOFOHLuHYrk00TXzQc9jK1x+K1cJwqBcBvOlQVdwElAtp0ewED9ZwjCCeV
3Dpp1fjVkdCIejfw30M+tX5qx8bkssQhi3MUQMvAFlz3K8ol/baJDDxwJtd/QL76MOo6wi68xKf1
6/UHn6l2Fv/d/3Na+la2BhUD0w32sA3wUZYl2ocJUTqwZ2VDzUhy8f/YtEHsyooNqe85oJc98CY2
KvrzbH9FSmid11E7s7l/Gp0xL0/lhOMhtnbF5hW/wn5T1MR78e2Gib5IzkPO85tSb716KA0PIlRR
1xvmOMvanAw278sNhNR8WYpxJ7zZQWEEwzKdAg3k9O91zHoO9YVwEOGB2ZWaIldnxilZRmesx3MQ
z0nn1LDrsRFBzfMxWvnK+flPb2lXzITvUu5/7IlRvGQb2M7lu6gLeiUNX2YHr0pHBpC2DE1alxjB
W0I2Hr1kq+hCTRGpXiprcnV8y8jxbBK055+TT7v3J1MFMAFVyeQ4q5BiQwSHVl+08guvINNq4U/p
pK080dnBzlUYDf6fvwQT0VOZyCjY4zsUXA0ijhycMY8FE8di8CaBIGQ9GGoKxcSvvmcQQxi1l33u
dN6LWTKMSYC9hBPMdQdqlN7mdpjUKtpayLEou52zvJJ73UHwCE/Ddwwo6PJV373gyTn5yhXHMfff
v11WkUrSchVc6BLLGK/6kJGSgexxD3nNgqBsZ77BZGG6MP6dtdYmKdfI91NzzAXnPdo5D72WYUwa
wmydjM1OZRLhJl0WdWPO9gwkWTl1ztWbzngRNBCuN/3EG+DeFWeAgL/6XslO6hWE99nDmbABUtXb
S9GFNjN9NLD1soC/3vbW2VHWN1FMjjgW0BYdPjAilYrdsTg1IOSUGblin+va1zhTHcJ5zx6Sim7Y
naP2L5y9oOELtqqsmjxZS9AE7ExGxSN9AxPEdqulWHGQN2WMCiqQsyCNxHEAIHcYANpxTlpwFFAJ
0BbGYQuSxVBGg1pXegfDbOx9xtoHuEf5rBKrc2yqxyxij1hAfI1o27IhBHKU18A9gSRfvipPQEhD
shHZXb3o0gIn8eQuaLdargX9jN25RJjtuETp2Sgp+lfvYdNvZjUecQJNVCyNwp0afYmRZOqQX4+8
UbHsTXAJbxNVjvsl2u9B9Ujm71ApxTSHshyK/NUVUfxT19EgjZxfK7yS75/sY8mekxm3srMV52wf
Rtzj5k8H2jCk9q1S59erRSoLmxRz51IhVsrVtK/HCKj1KDm9HhHszVhwYnu81ruRVq/8Um6C+KCT
8PxapNNW5+JezqQQzEaQFCbbbRcWRxbWaWjj1KGmCTpX4UfjnsxnvYBq2JIP4YUFp2vrI3W75D1+
QBYkfDGkTHiTWU7VyxAK+9LCVA1L45OQzZdxEH3pkJmnJKVItuCGRiSZ5tf5WhsNvBHWiSBJ+wsB
uG/hBZYclKJWnaTEKhiGx8AqwYmyC47X7pWv5XUgnRH+swdshxHkfX7pK+E6jG+RORo53zGFO+Tu
19HToo/cRGFk9tem5C3FGNXmckHLilF2NtLj9pgofltIDoL8r5L8MwX+jtRF8ulOmInlyyqljWL4
tv5Ks1wtM8B5LOdGTLKfrAKcJhSRNiH3j26itr6zxsaaC/WI6vScyU4yIvkiLwjT7IBcWhSvhgHK
8whWoQVBLiIekBSY9Enk+Tx0epAEtk34Zc0GAOxo9bmv6Lo3fOo6df1X+XKC+NTQABvZeoWQCX/J
PP27EHpSoMAjm3VFxT6OYsPg/4vEoFc1IkkRjOO/IkUHvEmXGR+n5hEZ7Ix03AVQbcP+N7dKLlri
cVwI70bz1UNR4KrWWBWQjprKQSdZ+7fDWhnqebuxRJ14gge1ox8PsoM7jR9Ji3ayIRpEVmkZmXZB
db7qVtD3UVPQrIC2CPkOMyTMee7a+RLZevmn/fwWVYiUioUTsHsvXU03QzeMWjK68wyX+PKgLcRx
T8kDzrZyV/FVBNhd3ruV7/s7/ekR+WAarO7oWAlGC48r78sMLhsg6WYfiTYagiO2wt4C6K+DUeQ2
0oKqJ/8OZ/SZQbpCyFV+rh+DpXREMG2mEjQ9s3BC+xCKjoNHjaaErpvWBL/HmfCrMzhS+EDS5s8K
yrDOCfh6siZgYv4U7F5pkhy/wjAo3z/Avfy3mpS76POue/JD2onfD+0MZEaE5vl2nkfpEugpPDvB
5+hf40E+lKXo6FDywQnjfMlCPgZRaiG9rkAQY6ATrzYpBjCOVdGcF1mqSG/LVTXQPs1ss8DqOy6G
UhYZiYZdjVfBpc4oOEqrFB3oVxz3OzSMSC3ZrCDugmzxy7+Xt9Z7mn/DjTQ8SELKMWy7kr9npyzA
gr1UO3h01hxfCRvDhmOSC48U7/VdMHQomSslGcqx6QL20MfTmAcG9K2jBF6pUxzPLG8D+o1uhc1S
mSB1GGzxzJ3/h6UY/4YDol58zMFHY5rpGlI7LzFlKyx5cih6tuIF13v93h0gJmQpiSqYHEoc9n1T
7yG5TsNlhmmdekhITvlWQgWq8CpDp6+HD2phlvB4nV2W0eSIS6g1nIgCxa0vWAwDZPjUj6k/GS4+
JRmjuxLN7794MYuAte1wHdOLsmjmVELdvYxSTuHu0A7goMQ9o09lv9tEbW/Dt8DyRgIXs8l9lL5g
DVudl/Y/KedZmuRUw+2ZtvW1EH4ZPununnnj1p0SB6/OZcDLeepE0EwbdG5tEUQYPt2nQHhp+991
nVsuhay0WzsGLV0Jz3qTuqoFmRK6mTFPAnkYtHJBYXs+sqGzUh9EKip7Xhq8LX0CeUYN9R+2z9s1
cyshZfS+grZVgIWcbUbn0fHYlj/Nb7k4ErfoXmA0CODKwwJ5eK8ue0oDrSDPIJLdQlV3N417VsOd
accpdZgsg1LLq3gy7KtNOtuQjGMKt1vdeR49GHxyO4Y5JxXnHPSEv6tqgTTin3WdCxjIOAIWNSWI
Z+/JoErwsQGYX8633mMxh25yh7QFpawGpA+A1pXRhe5f8gvqTwx9gQcWJSPt4mRcyNalXuyRmSDx
tM8bVWuwF9q0AxfVDIUUl2RqAc1mQHNiUXP/PtFaWsvidsNht50jK5Axf06lm/7mOTqGJyGilBxX
GuuKeMrlM4anidWv9Puyv2dLD8ExmXeg92uK247LAk0YbvAcsHe7+9IKHGo3MNrg3TRJgr79umPl
EjmgzYeb9Mjf8EOx0bp1D26vEjsIL64FM5TeKQr9ErJjxYsh9H7ZnnIJVHvcGYA3zCGieieplMm2
GuPT9Yhs5Z93cwZ1CWT/7tGbvtd52I9dtq9EXY2MepQ74wmbABm1U2lM5SJpaj3JOq9UI9D+UPju
NRyqlN1ZF+vVs2F+a2OUkF6WSjfq+T0fcfVe9JbctCWHvQqzVlhbL3+heBnwdM2ajF7VNT0erVfJ
GSrrrP4LsAXa9dve1Wj41x/DUTqP04km5q4EHd0pVXFUqPbzEpfRL4JA4nA+O2NVEr1wThrZmQaW
+4ZuAeMp22oxCuD45BwlkTYgNMbUO+OF5InMmqkqCX9j/Rt3iAslHv5+jcH4jOawaJZlV7yBL0LD
Y1FLx8ms80InoSi3fWrlwrxF3rieMx6GmczcHKUIpXWk69hvNl7obxalWZKvckm4S/drABYhKZ7P
60kp8kq0SUI7pij5oxDakX96y2y+8pIRDfbgQkvXlVQIrDuuMOkbZVGcaYyR6kbZfUywYyvRz3qB
vXCwQu0RmcSdzvKZqk3M1oYrzNQC2YHi9H0Sw1tMNehlJbMTwB3K1rlCMYmYsSP4AFSLiuNTJqK2
kvES/GFu63G95wrZWZAAS+GostJS6HxR+I0OS8IimLvWuN2TtVmwFvcLwDHA/HDAxGl2LmHYMOOP
N3Se5lMVwXgDlqLAUPWuIuOFQwcJgHL6x86RLCVSt/13N7tcObSG7ZdnaBGqFsGMectYMQkh2Udn
iE7M9M+QKJQ+08MnHKWHqN6EvzHfWEVTbOVW2By1cHEsRQ+8Pme/HjmBv7WOXhyYxPf4HAIGKwry
ycFA024iz7bHipPQ8ToPcWNYhbQyAjqAckykbSS2xPKUrNJROu1/7MLXKLQJI2QkviLlL1vB0IEi
KpiQnjQ9VYS8cvWm7RIk4vluRZsNInvVh8tD44iw5h94v6WFMsmckkeZqlUH8DAEpXEN7rnpoXmK
h9zmcZ4R4M/Md37T1WfXVk+JobQ9WVTUWMiJ/RWfd9+WkI8nFUYgCG6MUdaREOtbHogGOzjdamsO
JDwvTfWCq87exs8k/IUfbnfGWHy5zIbzKl4ofv4w69qJKjWT681RicYlBukaQg0DahJJ8W2b+HV6
r11GNsgxSUwwf+JT5RmV3ewV7kTRWfbTsTYu3NJMiux1DO3CyfW68oyKSboxsplgo0xNX1rjwZNV
g5a0lJutASMnVcZKEXkpygm2xBjcGoR2TuMFTCpLXQ99whEmCi/cSbDSH6lSKlg/EyMHBl7M9HMw
TR2cPGvwjl0HCPcWBiiZfArPqH1Idsn+xh3FSNlP08D4mQPGlc2SMk4LA+Ag/St0DO/MbOpFNLtK
7LTxMoorOTJZBhYLa/oKoU3cTs4voFzTGiNipvXurPJeeNjJhcF5PWAE8itAUXfmNGg/VMJT2Xky
icTMsULysgiB2qSOkH/dJ+na8/W+LzoUzxgKpsDkZHLQie2L8yqJShLTV04wX8KKNNk5oRoIGJrB
yOI+zjO0k9xjMqRTC5MFdnngfmf6fzRD9AWA5biWkYGw+9bHd0SiSvfCIElAtqW0QFfZvXUWAohF
sAHvHvjrmXm7GTsRk228CyQjmeOusAFlQ/JJEI+7hpxp8+18qFXSUyKvDh2wwlhPcxYL9ouNGRBm
yoQ6AZFB7Js+SiClYFlT9thpGpWTfzsOtgLJjzfIfEs22Egx5fO3EfxBYs51B1I2JYLCVCcf0tGT
t3dLCARndwYp08tf9t4j0c9t+nwh/AgLjkexILEXW2g6eTIez2AR9TrMnUEc3rhmwLgx6bLJr0yA
mcCEPwAd8dDZeuaFR2iP2+QcVbxFbrSf7DseKq9P8GDdoZGrnW36aOHfw4y8YTuz9pZNUGLV68RR
1XyUKRx9ZnxbfJX0h/8tp9Z7ICZKlW9iXOasXN1PkJHbNowHc8mzndNaGLAIDqkNZGquB5+2oLYT
p+Vgx2UTHRZD0ZsUU2qaJ3dnqIc9qo8Rl96P4J/mVbjS3+v38IHJ7gJGp7hNHbPTiNrd/ru8I4kF
bODWKXox8WtIIGzXgWlCbj/UrIAhRusOzWM97axlva/E1uaV9HsmjtB5jW8PVp28/soSXOGC1i9r
ogfFt5Q2nzhGC10ZhBUyd7pF47BX2CgCMa4g+VZ9knzPBOc9U0K9gb83K3ntEIWUFvmiQC2hN8AW
zo0EgDX173NpwXiw4uLyJUTypxT47fYu7tO4XZDRmvCWkHmnMqVC6dYnkKrNDB0daGt88mTqVZql
lpfrQlOdAql6uKlpgvyxySX9JOTPrFWIU2O/qCVUN/wiQw8SNXfe6Lyc8FA/a3u6gLW4kgdLUKr6
jdbEdzjVFORzTK6yWJBUXrZl90SkDTIpqUHqdy1HRNCcOLue8BpWeCGbk2MEtLFAFbbPF7Jb6/01
yr+19bLoWmkMaCFLu/K0NDBT1AH72Bmv63daxjfbCV2GxPByW4H8j8fYfYKsj2nQZCK7UdXfhet+
DKfz93efRbgKcTw/gigMazEzH72m4Ru5xzFT/N1AEjbDW6ev6PA9mcAMiA1mSZHEfd4JfbB5Lah5
I3PWeCR7/h7X6rnY0jrfbs/H3bGp7DsOjrI39ci/TIMnqBnyKhyH+8aNRpucA+guAHwVoVviRBzS
C2NXQv8YuuBvGfgr5ZyIP8yeqk9f7Np8Z5z0jJVSExfNLWH+xPcXHmF5mUag+1I4LRjTMeXXQKQQ
EoouRT8Z+4VR6h7NRkL1Hyt8mjykFStK//1qkn+lUMBqkOnqMwC7CYMpzj4fXjvwSZCJDKKbsGEM
wuKbmOnh5w9bMWaIhzdCg3b/RyK9frteG0gTzHWmmY8NpEuP1XrhCG82x4kq9pHHDJcsolyf7uH6
FLb2YxQGATxSkvh4mpBG8zr3heZB45GgeTOW4WI/y22v0QvXaPzuf6QX1u+2TntHnjyi1n47yfeV
SYy0RbqNwoe4ZSla9HLrYh4tCE4pUw3WzDg+KI2EjTUIVmKgbJbZWm38BdeantZjrh04g04Iv01+
d0hpITFUiXOb2bx43vu0L92VQ2g6EznMGQPdjIGCuhdGfay6Lv84cvbXckrtooZsR5wNwbe4GxWI
bnC2gB7n2vJ/3KkyCUtk2bVahWmciTsXKpV1ONRUZ0ot03eq4vejnGiQTytVOhK8KH2ympeby+9O
ISHof6zZ8WQwjSfsLhhg7ck6c9seRIhbSGN+xYi2DHA/ZmWX+MBBH4scZeosFtcUCazbKY+rKWGJ
307K5sbqzlc5ZggEKA1QolEY0JSCE8AKQlMtBvEwUzpxfhqXOTTC3PF8OpG/KEzuq3u9xAABENUf
cqwxLY6tnfWFIDLKNELX4hmkdfmt7IoANWd5oImZar+Isuxzo2PbdTgiHujK4QFZZlXsixBiyy2d
dlKqohoYxwScd2Q0qI609l5sogMmEZ5WtNzRWNEAb2A9nmoFPQL82m8Rge6Dz3fr7eewk7wSxUHm
UGTV7BUuMvl14IgdsxhqlsJnf7x3uJ89M05/K49VgIJ2kCshjDOEFZJKxPC0uUpDgvhZ1DpIvFSi
8ThTNkDfjv3P2OLXX/qFJn4OwjFMfVUVb0jGABINikU1UBkPxNR6ifqJNq+sJg8XPKHQAjQah9lx
0nQ48T9+GE0M3JPPsiGJZxgAmZrHSKf1qz83VRH0/a+5tKTtzUe/EIndeu2S/RAuw9msL+AzCc1U
mlo3WZtS7zwo1GzQhi4Rfr1S5x2SuV+S/G5C5guMH4XhHHDg22TKMgXhkPqW3Pa3yCS0wi7yJXtT
bMlBHLDp0Cr9pW1A1yjkeosZe/wS/ky3Fic0sFWLBvqXpRfR7/6ba5unuUo5+9ZfD9R0j9uE3M8o
S2GI/L8sDz9+RaW/GuWHKci/hnadiguLltDg8srYE58F55gJftliqzKIq/t3HXM5nGmi8Vrh2d2z
o2TPuqE1rvrMdLS9J8HJJZZ46JqIUsKiGafQw08oDJH9x7u+WFZVbamCT6KxR9eohiP+fP50lS1e
H+vO1mvza0AzhBM6XuNzasGQfdhHwe1Gyk7vF218zpJoqgIzNBgbE0URXCRve9GlGIkEIfPB2T5l
KJniLc4ldANck/LOhCDeYFWvqvdbB6fmjYfl3OS6UM8HIQDHd0kUmg8E6qiGBAmrzDL/Mo8ynCv5
noLO2FHPkfHZE0r4oQnqC2p8o5a4CXfIDAzc2UHpTmytMDKwWE1RokXu+PBgaG893GrwHiaEZgHj
mOOlGOh9j4opI7t0vPby9FUHEjDo9z+5O77c0q4ExYXold4Cff++QmAgXhcUE8yRY8swgY9WRZAL
gV7L7V2VB/H/Vyg1IvAcfRavws/lJWsc/IMDB5jykdOXMe+jQKahc2WT/wEcKpzVjA3Kmhvu4QMg
wHyM8XWan46FmO6cWIbFxixzkNn1/huU4hzGCmjfZTwq6oBCopeIRyPAZ/yz836U5q8qMad22yTr
idgAx6uD/xdHXdwR3Q53s/AO/7weulqCwdjyehhNsZYNtKpVCK/tOMc3Kp8z34P9Bvrcm39neRlF
A3wd1yWrTwZxNfR/hDJdMd+ixuy54R7WV39Dne5bXFu+yF2jEwGDcdyRNQ1jsxbFx59HQG3L0JW5
yj7tr8xAyBEuMqiUdfp/GwMobXQtp9gvicNei+0zpbscrUrI9x19Carly6EGPIilxLcZ4EPBJyH5
jIKbSmWVqx0PwPzcrwOYnZQ9Re5cw/Oa17Mw2FMw3S1H06IqLtT1HepmcSMlIqNQARo/wjsLcuda
IGvSydhwHv9rIx0GieFoaBf6SGMDqzlmA2t+vUgpchl1D5XbEMI6h1AokyX9uEwVfL2Lz3HyiF+M
/Ungd7CxnEOPKdxQmvOrMRA0TdCwq1u1dJW6/C/oiaulbB4zftHBcF0BVVzo4vsuVZIGsCIIWOsF
gg8V3yQLvwOhgFuv0nm8yidUnGvGt6jSxY6TCyzzB4vE7FjUok5h3lL9PzRrr4yGCFXb/kIUapCo
T/jcg6lbEm60Uwv5h/zbJLc97iF0f+0D1+2nL6K/goq4KoA+VQhkRRB2HBSdKtcQwgNrtS79LIMJ
HpKgrncyUISvX+Imjl7ILSvx0gqqP82YfZjYK7yWhsROLOv4AIIuNhlFTiIOyDJLdQbLGn6MTVcN
hO0kQPdMH7hF9V/8a/BHWVexInwXan0pqCr85Sj3GgLswrdYkNm4t2SY3PgRcRdPLsQsdUEy9Zip
Do+7CWFRpYROVyGL8mMm7XaT/pUgxw9m81NJD0aINOvr8+W1ufLhTmp/ngHDjkqR4TICcNeEHSLq
3FKOfagaj+Gl0iRFfh3SqEGwKwDKD4NTnbbp7SkFygdjzIR4y0PIvGkafPUAQzpJS+oAcJ2zNT03
aC48Yz9HyWlANf6JUtLSyVIJ6oieiHJ/oPGozFSCbO7qlKvSutZi3BoPFeNbR8TdWcK+DKxrn9LH
6PyFmp/zRufeaUSImcykJQma8z9uukEyEgBJREK7FxHDHAMKQXG+st7r0PQ9LtJMbEocxG6v6XKy
gIQuMS8W0ota15Cc4o3cuvi61ILZpwVw1u6DcUV8kpdhjXgSf/GdkW9hPXeNArcsV21eXGijk6ZW
gTPCkselgXm4Tpa9B4Xpy3YgxWSPfCKgJadQu2Wjic/7Plceq+BHp+PB8amabsLtBELcYuoRos/I
zhidCCzSoc4rw1xZ65WRH9RskJNlMj1BTRUf7DlJZ+4WxmaMMVANCb/FmB7sobraXNNzpk4KpKK0
9coY93XnvwaHXbXIpFLWGC+Zt3USfNIWZZaifiyDJPQAYNJ2Vbo2Lr1go+d9mDX9kAcMgim3X1Ie
geAHMwdaFuO2P47qVCg+JPipaDeG4w79jlvXPbSNaZjyWk8uEcugLlaMFVwh9z+PZ/vQfaY8qAxU
C/i4pZ862gWxUvMxvQhim58a2imALrGiT3bcZx4/QNAQw9IoObJitvCUE3VQhx+YTqQL9VtJLeU0
PzfkmUQ4vH3jDo9XdzeGj1YYR6b/It7QBhqrnbsi/tXgYNiWh1rcmviPTULrAir48CnCzXMdJ729
lMbDq4PkEkUZeFSadwWW8/ENKfEQRd4OW1wPwqINat07vv9echaV3J0nNmMMOrmsyhTfJ2AdS32A
xlmuzYlk97siulu174T+I1ZUvvXS419VUy8B/uXt3qLPXa8+aPE9huEjlFVNJ4heUERwPyMhxTen
g9HxIknl2G63qt7Cw/oTbgDdwE9/q/zSS2jvzeCqXKPRbykC71Q2WvGpKIegWhuZiDZ4m8TDPOdA
uy3HLbaRBiX38dFV29SZKqiBiEm36pWWjRbJij2mB7CCeC+IroocNnk9ayULIhi9efs+h66eA0Ml
+DlD6aCRHKU0e/WGcRvzM+mi9RfBZrSDeNBQCMZKa4kw8XqawDOiW9/xnIbfwgZZyXY2Ft6Fhnax
qNcQgnuFjQoBm2s4jwX+Gnf/bfULzTkfuJehnpYok1wF7pKXjQqsQgAvttDCagCCtavStpcUjdo4
HQJn18DMYYBSY9tM0sBrpidKTQk1K9iSPKBtOxAWi+REPS0/gAilNarBYUgn+9IjnQQliNhYFxkr
TIVNym9Xed1n8hAYV6mfLdaOpp9F1XX2bSzSASkrc5fh0ERlph+3JD4ef07Nndm714AMGobTM+mc
EcOSm+3Hnzdb75PrfR364Q2iyxdOiWkdGZQ9fW8bpLtsjJ+AlQ+li6LtHRRO6doL0AfFPzkQ9hhG
EDPev+zcAdmioNg6G0WBivZjD+4kOZGtV06Tq9XWxgyQMoOr2U7UCobsO8zDSXjrTYmCz7MrmI8Z
Eh2aKZerheEnR/znz2kxowe/mMPd5OkS3Z0MHDNLTXTKMVgOri0XB2NUkZDqxgU/2pSgvLbt2FIg
R4UuIvMZ42QogiMZYq5lrqclDo94tyg+wvGeAJDRSfrAOXxm2qKgD/4QyvWOdiuf7TVCC/MogHdm
lJmlNnJUkk1Jk0kUdnwJAbePfbVjrYBPJWUfHTD4thZYF1F+p1myEzaop2Ha0EiplnkiNgKpb0cf
81qntQVH5RIHX9hcXbe4DN7rkeSmQQowTbGWy5TitfbFjuU0y5it2M2PXI1j9IQfNZIo247Zrgla
M02PB9s+3JFZD6SrkNEuPXNVYz89kDWHo6APlJK3Cn1Higy4u16Y4iTE8uvSPu16U2sFWUh3Cczt
Kx3iCqebnxb+ZOp0k3EsjeZgcG1jAdOH2U+aAXRVgTkSbtyQZYCJgd0GQuDFv8EOFqbT5GqdrE81
+38cYKRHbId8tLTmHt7yvn2LUhX0Djh6w5KymRMlW2k0mzyYMMtAUvXwak3EZ3nGDG6EwayVod0B
iYDVumPwStvU/bXNlEbP1tIcT5VQDt/UV4gtupd5VIpH3gif78qM7DACs4a9ycEWWZ3yWwvz0JGk
gNSBjcZ67MUcMy5haryK++aHEWvO283u3NMN4xRbFrrPSfqJRfY3VIHyJ/ftABvzcFJB0u67wHRA
7bVIxRwQ85+xg5zOOcwVvoZeco+6w4/9ljDeqGNYLz3JTJj8A9ukpsygB5F+0KPmTkOdvXejFKlV
Wp2f5GqAAatx90y12DzKQCv4PY17rnz0UuUvn7mWd6epeuc1pLEQUyIZzZHzmmDnfgH4WM5x/BhK
BA0JR6d3nt+2Ck13lAzb6lH8+STQizv9IGGin9q/SA59QxrHj+oG4zez0xk26Beo8ZTwCh1iWXXD
CVFf+7HLIoSG54V4MhoH1MshB/T5YXD7l3irlw/guoGAr5hS8f/ZbWlGkcMXohaZ8Vjyuj5D61Ta
BeO2smKp9Z/Mvw5fjQDNTqSkTrnq08YsfP0YV5xY/B5whjpkB8ingKjVVAhu1X0A6nsax6UCekrn
bhVk1zyZgM0jrQ6MaW6avYQm6KstMv5Yng+1OVpHDFZX9UwuqbalB8Xll5RFeyVR5Un9cwY/iu1G
72LNMpfCvHQk/cvi0voGfLbdZOxicQUp2Dei1oZP9VEjjtMD38xgQwdAWc2qNyUgoBOjhYSM4xfB
SVpYrXGfT/O3QI9DvDTopLnmqrlNWLcHTI0yPEp8zYhaGxpgnH/hdkBXmYdiNOZEFr20MwPb8FT8
GXguOeqPiR7h3I9BICqHCKAA0Rhk2mKBWzn4/4hVvsBIoJsujVhnkM+vN83fCoOKmWVVfMwLBEkA
oc9Rn5sjt4ZCDOHwEKU2SU50nkFaJ0uAJbTy7vy+nxpuC4+n1FI/Jt6AC8ni3wqrbFJqwHOnUY+i
j7RYkp3Vp4MdOjKq9//EHJZRxEAs3z9pZ89DbUJ1vnUgQ0jraFcz0EI/WdpY1GdxLPunh8l79hbo
2yXkRa6HqX8zhmgUkQ8yFT+HsL1J+l2GTzl40Bq+ZFHoExvGrm1JxTRfJxT9/OQqpBBTsGu9ls3c
Tw6pUyADEiMw66Itg0mxta9J35Tcm9m7Atwvdw5HOOR93IpPg2iOqOI+y1IOUmqH+iUv/4am3TKG
vzZob/i58CNpDOdsoSTohVzfkV64nyVRV739MuEAWd/oaXXg64U9rFoF2VqfAr6x24mHplz84O4S
NFl8xisj9upTrNQtL3FBPGPplpzDB/5ShO1pQ60WcZg7OpiheM5Vw2cp6FxiMyc3Rt4uRUKnpEtn
+MDEqtfug4Duh2VnezQSst5bJ138eE3KItipyEJP0EYzZYBD2w2h03e58y8NoVbbW6WhHL24xtTo
W4AOan5XaDekdTeAo+H3YomICIxAZeEIJ4nA8Gh9kjtaQCIRPF2eGjQCxPzFrgS8YmgKYvSWrCwr
Mt6a//ZS3gj+P/cygBP5DuTgJb3CEnO3P4BVgMLW/SiAthyFrxeHooLoh/az3nX1VY61f4b3EEYl
1P2oNThzd027qPj4SaefSuly4gvRqFhq/jc9cKZhHXpb212AHPCQadGTDexQOVg5PZUHVaXsrGkc
IGABRiNNqCkAko8ULNJpmV+umyAIAtwF3f3rX14iAW0AcgOnRbB3m7oj6fTiJiI6SNtdvt3JuQTU
duN1CiMHIj7O65mpjR+klBYFW/pJWoBnRzG6/Dt2Q4oPyjmICURBt3ac5PlC028iTGXhtX7VC43z
OjDdlId0nTECjMMEveDXR/ce1mkcq/fTeuIh+ATI6+lMKKxsenLDE/uB9g7k2VtPTwwSWjEe9LDQ
hQYy0Ux+n+3Ti7DGHXBdPu0lZ8OFY0M3vfBUTp+v8d3fxan1ZNXcpecr/hcAXLMAAWTbzneNmx3M
la9m9YdhInjORcVzzbtChdeL+QlEZ5+XH92qSmpgBR74NQ9xM2+XrxkOA89aEUYUsrmiz7hMKt+X
O3PwFGXBgPiqTUIvyFWkZZXxKvU3f3hT+LVeUV0CtBOEk88jrE/FVhVr/JbjKxE3i1I1wdCxyVgq
Bf1nz003u7l9nWvFD8kKkL+1zIH2FE1vFUoLqKFRZF4SeZ/D3KTbVvD9BhyJR8Dn+i9XZScMC7HS
m/Xpqu1A0ltKS9FHK8l8M8tYAbXUye83NCloPLEvbrjlfRUsCNIfVq78M9EiDd0LNaRBqzNovTLm
IRPmRZ2Qxc2A/4uC+EMQps04ST4xAjPn3QXG8/kSL/4WDQyzBpOIypXRhPbqHwPkuCsstbqyucxV
DXJI6aKF0ZmzM/MdZWxBmvCFxKmF5ecFB2a/rBywI4XiNP+WEFTKVjpDpu8dyLTs3FXvH5nDmxca
8fKmw99VNofpjH72qK/FM7qiBvM+fSijKFQ6QflOl4he2oOn2uxFc2NmMK56IsFjhH15bbBHiMD3
a+tJ2pUHIkKo6x5hJaqlC9uv3rDwBJOO+BDO7ZDW0JRafcXILI5zpWJbz5SrEUjXQa1lCoU5e0Us
oQn4VBjIR86wz4DB74ZgAeo40Xx9O1GZCNT92hx6qlgCtZt+qWewV+Ccoi4PhQ3ZkCpLQk1enkSQ
LtkhbCJsk/312qGvxD1VPvHj34Hpg0cASGjSJnwE6p1nLOiFShqDfVzXOiDm5109zObNyfMCz8qw
2zm9ePCbzaXj2RSufLK3Pqz7KwJdVCt0nOyCtkJtiC7HOyMmMe3w2FUhFf9XLXkPAQVewnxyMKsV
VzBRj1D/v3NvlkzMfXQwmBgOGawxGcm+dw4fXxqgJhCYPNp3UHa+551N02zh7dHIYZ4FoTXT5tpx
MrxiDpFrf21beh+6igDLw5meWd+EOkEqB8cWz8UDM/RRFZJVVt7lIAnHCKPn4F+tuHLF2iXqdPCS
Mco5C7HA5+9VgRcOx7yLfSpS/0FNTQ/lSDzHl3yxdQXTe7LwHAnAf+VTpaQ2/de3XscSmyRjhLKG
tIpCO9mxwqfA/VloPSRxUtTyrlDZ86N1fRNPUmdcVHE+N3HKDPZYUpdiM6CnpEK1u5n7q+eR05kK
4vFulvMsA4bG/xGDyf/2sGCwPsFrUAvFInjLzcAKALxTY/bDjnMOGwLMZhcCzS9tIu43gID6QGhw
1BfyXTkqlnG8NAcjFOEoMIthoz+gJaMKA9pBnpl4x78Wc2R0yDqINQwQV/VR4wVu426NSWJEpm14
xHxGkfdT1yqPH2jsGwsLj4oh27T616DeupFy4um2oE23HpHdhdzomaiG8VvpPhZsC7gmdUwVx/QE
ggwxelt1riQ4qmgbZNTjVZpvnFa1/6YHi8XHu3F1dtMQGprZ1BtWkyHKzU+5ojMTtwEUYyZXo+WL
ewQAGcuOxtyg2ijxFl30TwttgYwxuUpAKSjpw6Qjwa7424VmpUqcqGO0g0rYQrBWHD4FJxIivM3l
OSvUcBNABWnsiZXlJWGj0D1J3WQ23r5otLcVmnWpNA9lDiIeK0XBtAJjvNi6KBu3xK7zAMhyhDUr
5rdQM3rX7FBBXflHDWuJ3JD644JmQaykth+7FDnIGfr9S1klWAn5o/yduh1SN3KKXelzg0eAPicS
ZUWVN9vcwsNXjaouzYktxDIyQ+0505K1MHG26KySk5rFazh/+qz9HVR0RX7F9m7ztThBJV2MKbS6
CVapW6huOu0UvGZNU3YPoS5kkzIEFWWnsqEdT+rMe6/0LP6rRiAIAR1+qxiE7MSWld/kM4R5salT
OUhwYfl8e0P39pSKbptmCJHoh7DM0VyP9ymK+5RWvH79tbJYuysuetZM72PxYwrrsH85vHNdJSQF
qU+938Q72d8Rz88=
`pragma protect end_protected
