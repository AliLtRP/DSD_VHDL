// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
eI6pTk/e1/niD+qEcZIlgIVkMeAvOt45zta/0JzChwHWiAZ8H2yIskkXYz3dpKkBt5RoK49fykTP
/13we+mHqIkqK19StbXsDvHHWbErMnECPpszoTRRmYGQZiZY/G3CUp3tQuwmnFPaPsSnuNLuGFKz
FMUcE07obgbI3AW8eXEhRRC/gJCiCFCiQdLpX8NmjNxItY5WVFFOs32rtU9OcHxVtAIfUbVekHPA
r1N8vvr5qe5Gc+breI4BO5e0Rsm5gkErxwtdqVD2n+ciC+OecPeJS/f3MKdAIxWt0yaeKGSK/ISX
CgscJA5NhWYq1HsOHh+YvktRy6TPPspX8JmU3g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
1vgf+79FpT9KLaewjpN8sAnPEVUiQVJ6lkiqWNgpBLWmseObs4OEtrWID+BcvjdrgXL7UUutO+sg
6pKZGa71LzzQ0UH04e/4QD4hKZBByss7TpgXi/jYojcDiGCjDlFKapgosGWifSLeUSyhpt2zW6GU
UUkyMBk8omCDyjM5jKyrdriiOzuSjvP6avY5LMTypl+g/84SmlOEAkOAlZjKZgJtZvY+I2jQG6/B
DURbYSTwY62RtpPo50i8H++Qcb8O48Bp19aDz5n4btnfs71B6coJuksEYCQ6A38s9NGfqod7OI76
N/p2DCpx6d0F8S+STMrABayQDTTONOVSSpuwLFw4sh4P4IF6WCKiwHknslpRe70kBmzydCCsfOfC
CdgTQwi3d+rchQrJEo/fXNdqB/ny+3XcYWBIg1S3PKiICCXYCoEnkZyNrMC8wJxqqUBhqI4Z225K
41b9/8lO8KC2unEUrJoOldp4fzhWPf1+vbn97N3msN5QAn+7fUUUsdG+vOUfMsZRU4sH1oDlyDk0
TKy9vEUj4nOogg9ab7uzISUV/3rIMNtqEj0Q39kCCSduoZYszRM29VDn4f67fPiuonvEWHWGZcgx
ZHCO96qKCF7qa2grfSLqfo6ZHeTOgoaQ8A07tEbsK+2z1SXPo29SXZRevvPr+cO+QCUUwHQYSbnl
vP+dfWc684PUl1vMQXCDTU6BBPSdZz4vKu2sgN4SiPcGf+pagdTH9l+qbwK+C5vNeIAbUT3d68xC
maEDfyu1C/xjJq5ES4m1IRffOOoU5O1csNXG861phwPZbaub3yCxKuhXb54eSVOREC7npgZlfMFA
0cmmk/RA2gdhmFMySyfEjluyDs6BEcV7q1NRuzeXXqYIsNJQVKhtwhOWjvJbB/KA6Kj0glPBX2tT
zVHTdidpbzNC3Iy3smgC0Zu1qJcVBAivCiaySTB9ejxM5Cg27/lwadD0mV/xFNMfSngAqOT1TFCb
f8uOHwbCG2R8Fdz9JEdBQpMyBhlLfaOMAdXvuVYqr1/IiPowlcTh2uhc/qKeHlVjBJK9Om93Jv7+
F/yiQ9XEyZn3bEJWDNqkDis84LmssTU3H7JjNVoV7NfDRxencKuL8tSq2h8hRUAh+rQvtPmJiWFu
u1vjSsuD+5/oo529WWo6F027wby7/UPr/a20ZBP/LvtsO3ACh0ATrbqB7yA69KXASvQBaMq7sEO0
M/3Y18igQsRdRjKTv2eCeomCgRPkvCBXuQbi5rIcYRuyycHltYD/bP4LDEwqwi0iGtOVosbi5GTg
xadWQuW31Twv77lxz/iXWGjojdMKvqbj1GuNGAonmMKV7dlj4EZ5kgrLzqKd0DotO6G0HKrf8XUN
vdbWVawQMhp4c4cD7o8+uFxZqWiV/dOysdD7pEm7yEWmKnO85AmfebpApDvvKnilIJ2G4RvZAsu/
aRxgF6k0CMZPVrSVetEi1stQ2/rbluC5+4qnMuPNKI70sEQXFx3fgHK28qfRscqw9u509cZLCUKn
9VsUSObPiZQuXMQRvCg8eRXoFBsKY/CuWsufVtOltl/PAmFc1tgS9eNjARubM2M10MNVw4VQizye
BMGzV5IQljUGprZaYCoXvUM16iyp8fHpe61Hx+mqYRVwJKq71zBJB3NfggOQ0BQYTtj8Rv2Qq732
AUqQAngM1oKNZhODoqBXcqjTKIQ2Vbwkt0LsCek+59hBGiupqBQ7IO5jFUTCFmBFB3eTUyf78YWp
He84nphHZFJzDp9k0dHA8mE+z4LXf8lGwRVHfwxPbnuQH1QnuA0njnrEvhjvSs4TCZoRIjKK3anr
4VElrb+rClCPKYJFZriHg4bdjiknDkpTdC6SVoFTUqPUH4MNjokKz1FhL3DzFcpnC3QgMHSODViJ
qIUa6C88QQeMxOJDOGMVo0D75JhOUdaRd9bs/uBWBTKcrT76OM+Xzd16D6n4YL4rh9F7QXAIAvTk
s32ce+sCVNKsCHRyPMFWRaaweesVwoMSlFfX75AlpglmU+xt9b8qQrs3SRZx4iEWgETL7wopJTZU
6FSffgJRmgKkrgwMqOF/Xu3e9JJuX9oOn8Nri1P/GylzL8aegqcfzKgT2yhhobKmIdwzPNnuaUd2
lmPLy0v6f08iqz/ezY61HAkZHR4aHQ7C1UCosUIr2jgrxWgVv7P9AhnCbUoe8YBf0IyilUDNzEaM
5bbX+z7mUXHwoz1r/xYD7CHDXKl8KXQX53A7rTW+q7zvDmJp7azSKQBlJc8V2cG2SIqX24R9NWDl
GuSXk742ZoXQ1ZPJOE4HnS5/2RFEaBvWKYoKPhL7lh0eLY0s7h5KZPn0xUz9wNpnWrQafFFOmg+Y
WksmAz7934TGyn+/yccmQYkqUzRyXx/BOkCVSN89d4hcK8fWM53/r8sdwopplrE+c6+9HHvNrUlK
yRPp8F4NBiY+2Y0YlY7ncn+jBv3TAPJW9theujl5PLV/6ZJuL5dWy+pGW3n4wgubxBr4P+CQ+fIl
yy5wCGdf124ppK/arZBmlXyNA9bY7A7ITiKRhLv0/MXsXQLu5DYpMHQmhpHcFsb9WelFi3QDVpG3
2aMFS6dg4s35+ALxchYSwEU1u6YSNZxHfTyArwam0mCsVYTrk1kDlpik64o5B1oy5cctMoFq4mVU
hfASHg6IM4Bupw/8lJmcjlyXtj5yD2kCthG7pisUFp9haEEx9UN8GOq9KAZikvaeZT5FDPnk1Cif
DrIPVt9Ea15NlMRoZH8sOG7PxvWsCRCU+vF/ovSX0lUQeph8oJ9zz3YXE2qp7tZIqteB2N4HOJXg
NB7yjFzefR1Qs48tFLIKk11QKvteOVjLc98Xlt4soaJ+e7I8+WjUew1bOc5K6WVhxjBRQHdH5AZ9
mOCDUkXO89g/wA+L03tHZkIKgI375lCxaM6lEN2LvSofEGnLg50lffvkla9iMQP4aOHoLscc+0Dd
A/5NLbsnJOHW2VUDG1Zj/s+Kyle6fvOFXpTXA7BhPBHN94sMvxGRkNHaBU9guXoMzDnzvFYPm/CJ
uX+VuCtuOlzGm8Yuj/FdmE4hSVA33KlQWQ0Tg739LJKr49E7yfV0F/ZsXdqzafuQUIcVreXLDv0J
qrvRRLxo8fH28K8WWtbbPVzbq5gxTPMj4G+pNjGKIh4mpKfzcf/+qJGFI2X1ef+btR0bL6tTAxIq
/Lxzjz5kP0muF5NFlqDMHoHM7BK4kEKLpv2Ek2sWVhW2u0vcJCqKBWTmewRlkXk76u/sPKI9MnAo
cWn/RykP7/TyMWC1AajQP5IS1DLa8hyUvdGmaMtOq4yR30xYXU5ZKYw0BH6r3pKHaUJiT6rZ3sQC
zNT4DhmWigVrcQs9GTiWRP/P9uMpyGpi63cekLvqM9CKZ1j0G8G712jqJa9fo1LsRoeKV7xE0HWE
Vwn1ESzOkGrPz/uGAk+QM3KuXNaWb6y+vO9VVmehUYLzpz61X1bUe2rrJlC0oBq29heDE+LvZH2Y
L+Up6de1405uj6xecPMCyCUC1zfawHTp1vfFNb/5vAS1BWgPm87Ydj486bro0ULc9C7dwrCI2B/m
Z4zDircyXE9ft1YJeTJp9+dPkJK8CT/5jSbNjaekP4kyD1Sf0okxcAl/OeUyMZf3sPwkwn3By/KT
S/egUbgYjP2Tu09RVqZNQUYOC6AQKcg9baPrOMTf2UDNXzkxZaKTYhD21ghp8xY2GGcLv/SX0HEh
D4TCtZ0jrHEnFte/OetJ60AVZSdm78juCusFpr/bq6VWn2qANH8pV8QQ6SoEx5YLN/3ExFf/5QZ2
9IelmaNWqiNvgHe4yfGXb/+Y9zWGE+GzbUO2BP1pmlAG8BmVZ/N1x9WsmoG8fpvxThRafZRIqn0x
rN9v597XEPU/V3McsxNcZtKis4OBsKxw8Tz1/lg+SBMQ40LOxJNv7gjc8y9gco3gAJXRwoHdx5VD
dsEBIkr9qLVaX+lL1g2Tb/DOzKjDxrnm61IunVWBjLSsYUSHbdC4S+CHXkvDSBPwbpqS2pUI+MQI
xTpvdnd+OMETFd5SgltqKtBJv8cV7paS9/7kzkPCvXDzq9fNt+hNaXTV0yATsuTcjm+F7jEMk/Q5
vqjoLj3KYX35wYkIx71xH18oxGjj+hYYObi+w180UXsoYi/kK+fT39byGXNMIWVOmgeiDwazAcqP
HkNzgKzxnd+6ahw7P6/YyKxIUmfOk9xNNhB5M1ixN6yi2OWYbA6lhm5I4S2W0gHcJgyup2G9HZ2p
3r0+s2MwORxHUPqQ4U3Fl0Ut40hODNRhF/ByIu+j9WSl/xkBYe0rJy8WVrjV8FpcUjm2Znz98tJj
3LJWQuW0XaUq0JrUNzMsPRViXrcfUNxMTNXy7gA1dx/GpWcNnEpKveIIr8rL3fww0yFRUoeuBBio
ak5Dv1U6CELhRqPNlePVGmsfVZzSRWuVtOlvfSELneo/8RiCBl9h4cEtIwdRUwFI4tlrVkbVu+7R
+IXaL/twKbcqJuwaDBjfsB8JEY4kS9HpV8UYCoUQO55HWNtm5O9mJwj8HbfDNM8E9bhUJB9EPMri
2S5nyO1jG8Ogl8ICo+k5uIHoXkYbM7V5yulA5EDjn+GrkpmJSNuqSOJmz5wYjuPKMC/LeuNSSjSO
IUSxI7Fgue26t4/RraYBfmw0MpjP5okiqgYQONfBGxMCAitf3ke+3rsAzO+f6BsRARHc+Shx8ok+
TdF3LytV0Nn35gZ0PzFa6txB0GUXcABvmah7fyXyBT44in4ilhlaKAxE9vdh25BJ9ZYVjK2HVMM0
d+//t0u3yk9m7XPI1byPvhUXJ87Cezmsv/0NfNzQFd7+Kt2KsrpXQTadJKaifM34TjnwLkg0cVpy
XB/Y2PlvrIeLyzAkUuUrfn7tkotElVCelCoDqwGrBA9yLVHWNozC1Knusetmbr0/jwnjOJtNEpuA
gGIB0vkyug0PpEWpL+fCm26kOMjvslDBRTJUHHzy4y+/ijjFyc+TItfafWYlvZZOQgx/bvLHOCj3
eJEBNv1AdxxxuX+wx0UZs0cb6cNiE/KVSnL1jBimpwU+6/l9tZZWsQa5fr6i2f+2Jvd4Dde3nzID
0ZjKyz4osF0NUnLdGzxuXI1WvonPR5T9QH7OGF9QjMygKiMp7UAPfKiaaT4wc91I213i+oS3+2Pv
6pSStps+LmYW7mzk2YoXKUNyj5l6yWhP4UPkcBObJbvpoU1bwqLCIQqWmuXsZocRLoOd3dMK7h2z
nN2ZXWXgKqYQV0HDL3x4gIypslMnL8MdObYxOu6PWYT+COeRo6vSmaBl8eaowD/j6zPui2jEShLq
8Wyo7BChbrbtyKSq1tWOEti0+8fbIWuPYlmO3CH4/KVcDpVfIk+n2eblLiuHlF/U/eWuhSL7FY+m
mOpWKlr4rnkopbXguu4pPEoATEdjvc2Gy2yZgwHzfzb6OIztsqT41jgUXgqzk99PE1G+jc8C9j8u
JNcwkBrmkvJSP0ub4p63SKrSWim4AXdlXSHC+qgMrgIOyHBp5kt+dCiLmUfZKaz+NmmyocWcUoI9
I1WX8wXFbe1PC7isCLLF+nMJluujUPpFAowPg1UcfGpq+qex6moTfDM+tPWc3Q8cR6o6lxUTX5WL
4oRtg3T7V0qIXekyB0VXx8luWKgfo5LyE7dFi4l8zZpDU3Z39NnHZlosEGcCrRnzWYq8eD2pmCrI
U5ePp0cQgcu57l1diFQwEsd1pTul7OD922M6zppXFbu/FEAeyLZuLfnKKnG/AgYCVr47bBAHG2Pw
Fdlzk9Fr+6FLt3sQI0v2oQFNd92w35kwJXrk09fCRp/A94o9WHzPveNbaslXoPAALcSna8YD73n7
GBPw5tOA43rAvXhzPe96J7DxK1uBE2/iCgL329CfLJEl3fY7Sc9hRnHM9904GBco5Iz4hMqEJSn9
IL5tq8AEVj4HIPXlHwniKGwl8Yug/LGO0TUoIMoLH56fgoVwkhme+FrMKRAwrh/p7UaARNy5oMWD
tK/Epi3ZBKNBcT6h4p2IK0mqT24iEbaOo+6h7ymxfH1EFm9jdb1gy1pqkX31owFzsTHiKdN7dkVS
tKcqyeTC66I5i/5yxCVKlqmvSl0v9jmHvxdNAAexu2kY0jV91RFOWuhYBQKdhoCWrNIm776jV5Nd
9U4pPyy4rhLenL2rqaLxroSxf4NkNfyerJTwVuRY7jggXewj+PY3m6roJvAudpPVS4jGhtFqCWzL
mH3uo+yyrStcbUrs72nRpHFEQglIanrXJYmnCyyyAih4kTKyA+AySUZE7o+FDuxR5cFeQfBGhlZj
PlM3Dlod49cEWsuk7tjqCplT3zmMq57zKTObvlUK6e6rQyTPg9Dyy0sDthl2Qemr97ghjSLwGk7M
DJV4pNsTiLeAu+ut6fekXbue7NSUrB4McjV2pYYnwwnHLEUdDp4W9dfretKizIBKhdiyyusOzPHw
uOOdol/nH0z/WKdFBw36HbLcfHw+uebjgPBzL28YFcOYsK++4KOFlgL+w2dh4AAjdv/SS8iZNdKz
ZZieIwZvWI1aNvzGpvYQEKPoQk0blfxxbxENMrs4cjVcNcMlRNPGsaFoSGrwgEQmEc3nv/7yritJ
+ERNvY3jIIYVnjC8z/zhXoJexaUwQG1yaIjYSxpKuysSl3/PNy1SUMKnTcIm6DaXZaZhSug2obWz
+STJv8MFTm0kboc06XNMzXI5YXEqjNql5mlDnn7xpxLahJTdJ2w5DCJzRAK0vOXocO59uW83gDcF
SjWM76HKENatOmm0/UhRMmSQbmk5DcwVCwiC5097XMpabdNd8aua7+ZCACLAA5aV+mFO0DkgeYXA
B3d+lgo+5FKKlPIK7gbI0Qr+kSTtXmUDvcuoUm3v+fpfPbv/MyTlyiafn7tRCMRot9hbrH7IXF7C
iHrejZ77VTWRO0dsfot0y+6I1HdwHdZF3bp/1GRheJQam0zJIhbGrnEyZJWEwXePGRgvRwJlOmbX
8rjMz5+rcZVbTQrfBLhbSCPmpCRjbiSDjXUVGYyRy9ulEg9qr+MwBJiSBUg64G9MswpLs4DU4vwm
CNgTwRrxA0xEoFsLaXkNhgQnQsyyppBA2UtIbnz5LV1JKOiL5vBQ31r+nCYlOdeWQUKfVsiVqD6C
31Mja3aUGv1BY/64CJ494AUPQ6mrBO9O3sCTAKNTFL29MjYsdIiaeJpbDdYwayPMV9I71ChDTudD
IvQPzXwItC69CP0O5qHyZZNY8KHqdGWIi5XGve0I2iD6CfZmqi/rBZ3rAOnSw9N6Eh6qUt5MTz3t
B++SSczod8yPbnc228mtPgzHaGeVyDdn8N4jzGjm+tAoqdhkiymA4W9daB6vSSQeuB4mWPuRAXZA
vcRKA6Jl+EK+NuWrkXnVWSAK616acaG1X5uXjEsr0vspGI9672U4hT25rCOtZmDSuCPjOTkXI245
lLr08bk1QB/NjbJ643N1nvQZFuJ+zhMXB3ks0k0RvfVyLGc57aQlJdEeT0s2tC9aNHoJnmFHvmC6
nXnjmi5LuCRxGKW30MGVMWmTiSOlceX28bmLHzvbRzieDaBmH49BnypeP03KGcz6vx3l6xX1rMQk
dP/1rjY2A67XxDSOwiouDCG5TkCo0YV/t2lCn+Pi8JF84CKB4AWhV9CI2XrMt3HbCexDblCI4PXn
CpEmpw5Sth3DSJna6q6KFhm9zXQeOdYpye1g+edL1GdscNE5uv29EO4JsE8JHkcHIZcUJInSaYgo
oxzdkG8U/3MtdOx5+4KlEVjgxEIo+deGnGrwP5RzakLafd+l68Nn1G/sk5cgjMerPwvdTucMCM+O
jX0NDpqJFdCRmfDkwHJq9/QyO/hCmyzK4wylMtmlsVZ7BRmwNYhRCZZA+yKOsA2y58xbQ8phXA7m
GGhqOKuoIoXozaw3j0qNc3bxHaxGOFc9Tl22qBpEnysbRvfn9pAJ7eqTDgwZqcdy3PV080Wr7gER
8l7nGq2KhRSgzgtCYmz+RV8d0UspsqUbAbzwiBM931s+flHsM+OIUgrZJm4wBUW8rRjFK/UycsdO
QSAvpFKcFb5XvzPd2M1I6ab5nfasDopQS+5kZgrT1J9Wpgd0q86wNrjLeK/x3IflZDNCGiNg2VZ7
92Km1kW4T/4xVb0JTrRtOcJrpJW8SPasPPHzKdcjQy3i1a7bfif+Z3Fyu7hCXsuKbs68dgj7D2C6
mZ42McGIrzdYZAu8uRvn2jgBtjXGuiCnKPONBH2Fvf5pEM0iY93rwkO+twMOOvsujMbkAvB+xFq1
n800800HxGPEdLC3HrrxO0nxBzgXzj+/0EK8g9Hk9LATzQ2jn2mMk6gQJN4qXHe+WT36Drq44YO2
cPgXB+307PWSXNR3RuWM/0Rdmtg8QzKLAAwftfZumG6X1RlM/dNdcRG0zZCCx6J6On4+8JiUkwdX
55Fc3L31KQFW5T7JmeuHJW1BwjpAUNGRAeWQhSgviRbFDbiq5Y4/2OJ4PdkOHOY3AX1DjrzBlpBk
WXlWRoeaYYVqXRsxf5Jt4s15/+cqemfXeOp5059B4tAHgpGguB69D2YhXsE0lmfJqZH6kpFrm++n
hGkPJV3yPHYdzyr1buNzihvN0VRtBf/Iwi3SnOAUh8zqjy17SZTohGK5zXpZIHJ+h36PDIPLsGEe
5/xxFf1s1FdijB3YGoHb0gaGAwCc6CKEh2lC3nBGPYkUdjPau0vG/kJBk9dd2biJx8XEIuWScV/c
Hy7RiAXVadQ+TkkqR0oVXrtWga61JxzlnucykDGYOojuHRVGWkcwaStYLwWRWcdSJUrzs8RnzuBt
/oxQLbSIkSY8cTmpzD1RRI5WFKsw0397kjDtwQ2T38PlGBAcJtyM5hxoeUDXZrVQkvkfWr6T+z4s
u3uIlVGKRQbYpewFMSV/TUOf0LQFgGOSI1HmPzzvuq7ejlelL88sNbFy/I3PCFiGEzTtlpE3OcOn
Ct72hF9Huu0s37+67Ps3cDZ1EAwlWUoDDcS42A7sO05G+HiREqFDCIfUtnk1wvRD1UAKiOtwFkPw
6fPmB5wrFZGgdXo+1RGK9LbEnNG2ABYgFxikg/G0VMDdv1Tw7xbTdmjvU/v3KbGZqj/2fFVQ8CN1
5c2bw0g9LXco1NxKXcMOfQZbhJHMXQrDB+OrXREwWbbYBn92iwWgc5n0R9b76iwpRLnIQVSFtFsi
n2xqgmwTgZZMTEp8Wr/1hdaGxiOhlAoKEoAHu3bzNABsmKe+n8k2iNX9oERkXWljo+RNk7MYxDAo
xIa/oSojvs0WCeT7LtrJnTuf0cTXPeUlIKAVZGy2NibHXGGK0xuJlT5EnohAikE3N4us+t3p8Am1
ZT8CgC8CxpX13+bt4JsKgm9AEk4eRffqGs+s7XdEUF7SS0RRe7ZRVj4lTWCPFrY0vlslPjqPD/12
nV2rGWFrGNjl8fyETtogXP8ACRs8nZdzFzWsNCpXLrM2lrMjWY9KjrmVrrZ7CuF8tQu7xlAKerso
JlT25jkNEUtzbICMuwUkQtMsZkOuLhYUms9ICC1pG/CNgDCvixMx6tnKDNBJOpY+3Sco13U/nypb
YIsnnmvf2bhx9BRjvXAVYiGZHquPOPrQxqHtJshfUmxiVKpqk8qbLupxlQ8a3+piXDLFUoWfwFv/
Xkw433NoieX4gSZe+9ZHn0tP38BGxwKEMDMQFb6kr5jjEVXWf/NATjq2Xw1vmfKuhpYTTeTQVjKK
IUOdOikjGNfZaOG3Ya136KqNGn8KhpEozfREBhBjrpHvzUaKISrDnKsZCIp258tVZmLcjL6wpoxa
61ip6Xj5aTOeONtiG24jgH+UORsI04y08orI8vYkFW14Yz8VMER1xa/uQYoGzuHNQnafQhL8vAdU
pZ6eqTO5XTtavHpmlmhl2rDcVjbR2SsCX4P+uDLSpwTzgAO1BL+nNCSKCfsnOm581bchP32pjCYJ
MAz0rV+3Lzai/8/sPd30F6Prxr4Hw8l05ZzKPvNfZTR02eOJF0aoHte+gIGbcYVHD/xHvl+QIshE
m9Z9XqMXQiOiPYzjpNbte/J8zyjCVA/q2tx1xT7SkCmRSq8tWvcVkbN+xd8H/fofp/E7d0kkqtU7
4EIO0E9rBVy2uVNiE2tJXr/If7E+Mh6NE68CLdMtO3H/4ueSii3lF+XKMl6LUtFuTa1qiIvzeI4Z
5u9o96VxtL2OA3MYjuBMz5WdCA9i15FK1VctVITfiotoYbkmpOIEjw9OqTM26VFpD/Y100OMFEqa
qf3DZR9zJFg1lyEL/Xciwwr+3Vi1YA3Blcr2PdgQqmT6SztUpfWwSUVD3JqT4kNy1mDjBKWIkf+2
02eInmpRkX1fq/ypMHESlza4ovIB94F02szubWMugnAMC46Qn2DslPEwcGIBZzYM0/Q9ObTiHeDd
3YsJyc19wk+jvayKUPTSglUO3vQNYoaCmiRcFG8kMbzlVm1/lqytC1MrDOOWvbmMTRADMAAK5zqB
ZPPwDBfFHCc99jPiGNj+QA7Qbc+KGb7tC+JZk3NWRRsnR9tZ8xtpxtpsJ5HtjnJf+GY/O5pBxqsH
aCXCPwrto/t4vLeSZ1z3f9F4QtNLkX9O00pbKfzSbAIIC/J6FHnd5l4vJXmET2zgFGdtB6BM0pbk
nMkJoVAPottro83upppg0heq/s7oOZPzptnEwYO3wQ2h6SZ00/VpYK41DOYOzrZqL/LTRWLv/oGh
8EYxKjWgM6J00xMvAWV5Gl307kBffje3fz8dubqH0y1tj9s5q9GS/7dROkprJqYwrz9qn91wcVXX
9+0d6TC5dL0eqOikyQ2qM0Yuhm2UCEvLiSt6NN5xefy1pk9R60xeQ5oZkOXvnG4ypvSbZBdhegMl
tJajabWxKz0ykt/cf0CS2Itw0ETgxe0eXExYaTn+MTY4Tl8u+Q87BNIVWo0wHt4dXMsQ1bueDpmy
9IICMUlZqWvdQhh112j1W3SmP0tS8v9krAdWjCmM/0OGqGnYWb1sRZ+MFOHNV8Z4pN4hPxakXYga
ka5po2VzrwZH3wlX95ZxzVuQvH6qOK34KJo2NE/Rz/tO8IhWpxtvEmc27BG961Y9JVJOWLVys7mD
zzLd1fxKQJB1XlaYOtxEg+/BaYzbGWLs0naxs9orbvdhnxFnivyZqVuONzOA69PveHW4gbua2TL1
n/iMuJiAwPF62Xwl4TD/F0W8BiAqMgZszEMXNWPb+XsixZQr85LTrfeSs6VLonVYhIZOlNs5B6gK
VhIVoNdW/WKOVACfxdd71XrQIVo2M1Q9PP3ZiX2Ezg85OvNED0RxxnYhpgFG6xhI6HhGp+JdWEmQ
SRlQyX37Q1bdjlqnpu/puQdIc1xz8Jo4OgEZ46Fzhn9RJK4wun9mqYlsVkiwFct0W042F/NyXMJn
OiRIg527Oe9GoWZHtVRXPMvRysyN/6Aw177Gf3wtK1+SyEA2RFP3UPvTTe0TN5ERK32+4TO7K57o
OnxFzYJgX6QadWPknClD6bkD3PY6geLZmCwjjYxMoZFf1t8KluQC88rPqyCYKl+lBbj0dQR4RVx9
4jzN1oci3Yl1VFV+y8+1iSi0g5mZU2AwLk7Ur/KVIsxqrDdVbR7IB4lE7AfAuQVr8J1e8pZqWmNK
gxwcOXPLzDMk/PY45AlPy/7j6o3iy59T0rVjfCB7afupk3d3sU99tSlbXt2s6ljq70tqnUp7L/fP
jV0QPNGs5MdQFj3vW1Wo6NvrZRxmJtRNRH5WL2NqtFA3LnPX1iRZDv8b6Zo51jEiTZ/c9neCmOTV
G1qdMcEgktrGzHGCMMphiLLd9jq+sTFnEUvKUlZwZE2AyV9cB5EPMsV9PIcmLL+dE2MDhMESBXoQ
x2RMDcbVWJOgQmNxF73QJRgr3CCV7btjuNrW7aqfsGmfzMKtqSJmTfCC5Tb+j4W6DMmoCPXEyzNt
OtwCdIgGd1bQbKPbPnSxIPlFP1L2j2NS6pLDCnH4SnCnD4zhK2Ycw7Qf1yfLvO7KVA8nbncpNxmC
lwvXWhZtki2gTo4zZ0c0oNsMSBfq5kzZts9hur5puLUnHq2AYEsFhH/bkTlH1Xqu+yEVVAFgfQTS
IEzxUwSX122IbeCAIc3FZ7u6XiN7wmhsrG1tQqutUp0t4yJPf8K+us/2O+qFlvEeu57Clj4wjEo2
j/Og5bjbsVA118530idBKThH0EFH6Y1rNakdcM/EmvXKXTNbl1J1Tlgwu3WfPItB89e0xZt2pAAl
KoxdvyvDWsMyJTZjYPq8gplbFDpJVUHSPvkXFmeGtpeNdWjIu0FdfkfzApaQM2d/+5iyzUw7nihf
VkenATDWmxWmJjJK9mpj/vH/v1OlhX6UkR6jTOa+EuSS+XnZOeSNCIeN/vL53KCjlOsBI2PLKa7X
4weaUmvft5WZNqxlAyd60WgZxJaWNHapGeqBVr3BoUHTIJLyKR8GXAOnt+YNpAUQQX3CTb1vmTCx
gOJSPozyPdk2iAcgdDvzeCB3M5lvp9JjCvhBhQR2DUx6tO8f/F/W4O/FSp9gQPpYy8K7h8QiW7Kp
7W9IKs5DFCtPzOWdEF5Up7y41UMH3112cgYG1Ca7yMiq8vg5A41tXcP6bgDmKVwpNA/6
`pragma protect end_protected
