// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bedmziJ1WqU273dwMUr2/kAGFEAcbLR3Xm4k9NZqkbJJrUIZcsp5CLpnhduyYDXg
5N7ccZENDENlhh9jUPdOk8obsFcrZ8rYAPcoOg9hOATfzM68YkYuwLwbHjhWuygF
BG57qeB3/+bq9Dx8yzJtUe5c67HxPqhju2kzYODuBVA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9040)
RXqZhWEYzWj7xjXbNNlZqoEjfPlzfpoJvgWFghUxtXIIjktjhA/WGvTuUOgKah8o
UJt8nehBs7bXiqODZ1OrievHTf7Ryctlqe8HiAvC9S49GopTyx8idMMTTUtPXzdE
EQa0/sXBSL3Upim8taCdNh+PEmmsHDvkvumAE0AW9SgLcOoW9QwO3VN4q/+r42a2
o3z7NqlUeMKP/pMp7x4lTOBKnYE+VamMByhBXAo8UmXyp8sLHFGW2Xfvls3JCLmu
0Ii4OZpWTfgxrfNDkojVzuWlsVRFbQGpLjevvLZ6gy6g73vogYke1pyCRupTxz1c
BKM8xD1jsULVK1E4XjqIXspALQP7gpuYdWoozOLNmKASXB3mf2GUgA3Y8MiTfPZo
CRUA8RDx7ejcanwlYr6znVYPK84lSrBG0/gdOnzX8Ge65OH+jBqS7gOokWYBR5BN
beY3kkRr8g6XePdyDPfYO7CrFOm5eZkpZBP+wctzlCarF4jgYYP3dY82uNJC4glr
CwlZJYVXpyk+lvqRg52ZpeIIWUGw5HWz3Qb1wUEVv2i8G2BAzdIimXsgzz1I+6ah
5P5JjPjFMtYQXciLuedE0MMgLHsTvJecDlEoDQwLEzMZYlaz/g4pt5FEAZAtKuC5
Vd2Q95U98dFAoCWYSd+qPvb243mjTze8rmTT8gxPjWwGgTl8uThPkqcqf7jrQjLH
vjdZIZOszHEFMRF+Ri9t5Oz7VCCMT5fmmXYLX0Y97nma7sdMJKkiK/y832WQhZY7
1rz7CemvDD/0aMtczO6XQwttjrpH6tCYUeHfnMVKhhb5zOUtUK9IMh7+Os0EJO6+
BHLiTdKWwWso+RftxoKdTRUpTT4XWoRvT5H+4vI8xfn2xVBaZ7SyM9WZ72TwwviI
zl2IUZkAtY3gUOH+qVDmw/jfS0yhbFFUckCim5dopwUW7AhewQXgxQ0dOQUQpOdj
MmQ33ZApN2DmFW8PyIL8LqgO7DmrIiuUik/pZ5I/DhZz70HCJ92uLi7oAckO5OoL
s4JrfevtnLlhbK3KUtNlRcGMPsCtV8VvnrW3x/HTwWgADX4NDcYFbuymk7DwCjCG
wrwtvkxgHz+d8vYr8f4hz8oGivF5wlKBi/u6GS3RxY1OHtFrzhCI40Kyek0W69qJ
pDiNjesm2fRVXp6/ImtgelfRwxv91rvJWIB3Nm+pnjZp5RSh2vJuPKm2av5SJsw7
9AQZUbinvV0JrkrMvy5HuW7NfxEN5OBmbKpKeZzokfvxjHBUQBUJ820j9LNnZHEM
1gxbTwHrO/9pptZ92hPmPDVG5LodlPxgwkoY2tphIvjfYDnNe1yUa2EbeBWjjnr6
aLgbQUR3okHjp3uk6U9aNXbaRNvQ0K9tuCZEKAC55sni7mFVGDuizfFOYZA/qItS
QiFGQt+Ur+piN36g9lM2gRHKtn98WVsrSvBd4Pp2jOZX6kKlwMkuNZTZXr1j/bv8
CRkWRSz5rAVFgUizV8fApj90XwX7azkQpTMtUlaIWoCQdUqrxmymsP6KPHqofcD9
Y5YLAWBddT5XRPMOc191v6fJbB2UdeT0STVHDC7CZINZaqVjZb581bzG/tCWoHBD
AUvrUm+zyBBkTiUGGCCZfqPrDL3NVAWlqUilwGGDQ4MrWpbHxWi7E2SoROTGyHD1
SSfkeMvtkCzujfeg7YLn7+YxkMGVrs44PxRCxB6sAcgspNM5QA14SnDV8p+gL+q0
a5bThuZnCZq5jWE5XszinoJnnRJS9dvALF8bz7ltNYMPmCCWaDCnuUkpNcFJaeNH
5qg3GpP8Y4CjZDC4d71/KU0otqOSW5a0PnKZEZfq7AEitXhr/QV2unEt0wQV7fRN
TOIxov80+PWGw2UsLb8/gevzopBSBEKV0seQ5aKRQ6kHDkhXZ4OdPjozDVUzYKFy
QOu7n5qvihMWwC/6SS0YP8ZW5YJQA7clkwGEYOKbazEcnw8kVBqvUfuUwPMlR9Yf
dgaKCDw/35mKlLkRrjc9K9djtoEIq4c02NDq04pca133DwasvYt4mMxRqFym5hJo
vuJVC9cAFtP9MSpTEal5a/Eful9iMhHHavddyqVKqK9s/xhbVn2NzdusPia/QUly
FcDdnhuuvtz+no/pBEPTbVpeO/feIeUqr/U1AoKLl0TuyIm5HiugCypHTTp3+BwO
v2Pz7pGdZgofu3mgE685ZQ17+u7pdJFfpfhzL2oSDrt1Zche/xI1GOwBTuAT+SSZ
t3+Nu/VDWuMcfjuceS3vS03rXGGwvxlorTnOWHoiyYe++qeEVpNeoeOYXyJtnI42
efq5gp/t/B3eD9KwUrIySTr9TxDWTsrUmHFdvJJWJLB1YtxoEa9ohMGJgNMkNgte
tSUds7SrXvOoZfJjrQEOIt8yihIEzKwpXRMeZarIUYO4WMWOb+jNMOri4rCZVG3C
MxR9FKt/6VrljSzMgkTwWbyukEMLWCsaUvfEfHfDpFLkv6Q1aol4c86V8ldDBNZs
nWdU3rAIt0aISxF3rZ1Uqc5Ikda9P/zsks9kA1cvxKbwEiBju9Qx0Vd2RDqRtD3M
nrFY9qClPdrVSwkljI2HER4ZUeFWBgloFO0K9B+VpuCnBrYrcUlUx3EMOAbGchB1
fPmWuLd53l5edCG+9wmlKSzqJDGgNO16uaahlsO/5rFnJq1eH2y/vLjOvVnsmfsh
Dcd7ufS4eYhC2tA15Ya59L/mMS5bF9Wu1BII33LexOEvuFZoyL3JnjRPsVlO1/Hr
blZGqTkdNNOPk1L2Y8ZVlcgty9BGkWhPln985CqAm/De/N9POE/s9LEqFzahp0Fv
Db7b98MKHU+C976LkwF+q/e21OOdlgMVKmptt7VSwg9ZjF5VQllhOoJVFaZe0/k3
BoaKYO+jjh5WJrAhvuNcheVm/nRU0X0OBV3/QQVDgkNcHWFeKtgDL0LOjJm9JbNv
psmnc8tR8224ieVY8t2CGexzAmtkA6ILptetszDxwGkNGaJP0pwkQtuc3Vf5O3/C
KWIneCKFpM5zkOn5CuxEhMPXDdI9SCrki6a7OPfuDcqcBwo4of40LaPfRqe2j6bf
V7y+Tyb9PwvqwEwdRzEHxT4abGr8Gsz2jhO/cZSU08vADCpkYp4zpodjViGLiTvd
q8NyisPMc7qJiKqATUN6O2wd7uBC2mLJPfe5It4Y6GsYrvZfPJW3DCGs+8hBip6h
Or5jqJDN0MILmstrSuKNODjAowirbDXu4cDez7yIB5JlHwkONmyABKky5LuJHqJO
jbzh/2lNG64a4OYfmQlW1FjxjJJDDAlGnw+j8hCeP6pbxstCuc92oWiR18cP++hM
ivuyPPrUKVBwEtkgIqIKP94jwWbjwZLJoJha9gFpyQoHy+7WyxG+kAv67GXM9E1V
Fu/gRYs3WKCBYwslgEmPmodQiy21tpvPLwG58bOT4VzkmVLMXL00OVqMlNAo0ni4
HrKFwWBVp63R66x/4QmQcb4QT1EMd3mqC+3Qlay++y8AU5VBmeJHey3AEOtQsIA+
2D/wJP/hzVQO2fvkqWwH5FJ6Csv87K/ECrdeaCpBoJiXmUJF7VvpUm9o25TSGR3y
uOAUZcSczjLLHuab2XWMfmE/dEVMcKztZrVoe1sEso1gNdYDTxGprpha/D1MDLTW
+u1ta8/BNdpxmGr7NRSYHejbxDX0nD1HeWaxPMXemdmmSduZsASAcQlYmaTnMDZ9
HfbMYARBxbNE9h1GNO0uMP2DgJOIUQIK9eO0cEQSyuTEGlSaVCKlb7Szg5jeKndR
cuGTuF+XJ6410oAMejt7X1c5rlf29qIZNS2hUcw3Fxg/E1c2rXoyfu0oyQLHnrH1
yjc7yq/5a8yb33nZhJi0xsCG7/jJlVilgSSinZGJyY5mIF90GGy6/zytz+iy4gBy
Vqw78YhoXtAiWWMzWx+eOW+5UhLRIGLfZENHvQnPeZrA89QVxf2js6pMZIT11oNM
JNoGbkAq7OvL6T/bUuBaCCaCuE7JJc/RDx+HWVocObYMECqNAscDSYQZF+ZnVBpC
SW+LGVaviy1HsrkpZDtxRi0BftIX7SeScZpwqvLqJ/C76jbs6K2RBNpzGdZT5XjM
0wK0FHA1zr6PiY9e8RouSYqBCZ9jbVYF2mcqSMXNxDN+jZSBNmLpSKpg9OUoDAdi
k63ayV3aWU1ZFsAMxy8qRF7UzUjRbMeWoQiYga5mDQQPUugOTnfZKlLxnDuTqtfn
J8z+f6SLnoXZng334oYnSw0Y3UT+Mfuz6rakaX0+f7wAdZdCZ1XgrhqQieKZwno3
nqN9YST7/m/vtyLcCEZEoSFbNxu7slYGlEhZDm4MSwVfVEUM9zyjTn2FxHyNJUkr
aFlqiyC6GsWZ0FPnf66zY6HQ0wLf8MT6N9VdMaIN3LGSkhEs2FkJP0U33K+04ZXp
cKbm1uDBlT3zM216GfwvY9m9fsCCKaryD7QbF9iRHksuiSnKkvNKpnMoMrdgnNzA
hDjT6+l7O/iCRt9WqEjtxCPn1nxcFa6KLND8FEyV9e8lkK9Ibs5J13Lbr6nlZwFh
Tl4LsxSHZW6YIFr5KLM0jbsRpVlzpD74wp/jZoypcnzh4VD8ZQdyiQwHxlkhUf8O
iuFrZ9JQTZNrc7Qllnju2UNxQltx6by8yymOS4szCQMGpTiUpHXZN97JeVZW1XZ5
RDL2+SyD4AfJHY/mVnYe11B/MXe82WUDnFQSFJzXn6I8NOloQjvvQSEjldBVmNVW
zJFp3o36y47GGaBcrZdbSVtYoKXlTdUShoNtznzaEPQ0c2iPDbrHnco23sBTJE95
7kjrbujUvJTt1tO44z58VEf8nuYN0GpWHvWCA7jKGb8lJHHETMbEA0gCjH5fCwcG
cfDS634bg8jAH7wyUknCp7VQ0SGkCym3R2SbJ1rk3nNZzQ72tktVaUcGBvGLQsk4
XkFWHfaLwzExtfNkl4x605v0J98t8BhCEdos+vFVguZinI+YVCG8CVLtbNJ500wB
YqL8NMB+5NGHM4jdR+wAHiQ1dBB9keRUrHc3OSv0nmzv5qhK3OeOmRe/nHVZyllQ
y6wy5oJvFtN/6crCGBHE8xj69MlXkvnrjMJnxEkJmMqAKAjLveVAYQ8DsnWezLPD
PntEpzg7E5M6otyMVmLhr/xH3lz5KKK33r7Vm3ssQvRMDclwSmV6hLWvvbN4Jjgg
hrzOBiHBQe859O32ypUESFIW4EsfyEDsROC2sEwUZRCpoGMh/z0jOsaq0Yh0yuP/
AHW7W3docUd0O/jjdaQofsgk02RTlWoQoTDGe5OJToawRB5SuUemdq2L7zyQ2/MD
gxdc0Fckja2mtXrO//xNm0XZIh4HpKqCGTtIFma/xPrlCTciG0hSf2mr87lnOJ1s
gE44zQ56a+2waLRALfiY9iM9XHiN98NOs5cRQwWWGvWVYtKuEy/HnQZXwx5Eci3W
EKLej0SJpO6hCC8xntwSZSFCr64Wa4PzAjM1fv6gDwvUKpa7Q/vhiFtE8LrtOmjd
gNL1903RsMAb2x8uB/2+nuFLMCiduTGexK1g67pbq5R5K4TGQ/koKQhLxV5B244F
+wpukPVEZSShvXDqW+iktgTjbpBAgEiimXDq0gTRWCGkOkqzl9dmhyANvVOWB0Qx
AyJtlDX07pk/zETT2xTAnik9oLe0JWX9DPM5F6KFydyo1PRcauMNt3e3L3iMZjn/
JYLhtrN+hmZy7Uq0AInY3GBeVS3SKEP9pDyiQK1ID/D/+8a7BXF+GPj6M6oVaOL7
eUml6soVEnxVt4Si6Z6LzIZS/ddFfqnTXHmO9RERigv+a+IhWcdPxULqs5X0iF4S
RSgp2Tw7tdlGzvKz4Takpni13kqHlnE8vWXEJaOCpwjPvHMbysJnPJ7+QK6tEW9C
rofIYyEOqJghfYe6ScvReQEryBPntzoamA2ah9jKuuK+0+s8YVQLxkitWTd2oqxT
oDYy9kRyzzxVFXZ1M4O4U0NjCRqjRKulZw3XB/9In3N9Ae9NtGosqXiBboZxO6Mj
W7TB3lf/btX49IRWdiEJiKv/RsTkNV0o7mdqK8+0haX1xEJKYx0MFhTzK/K+03kx
/YJRQV3YK8iRh2h6+KenLi7r7+OAEIkPXPHo/3xZty/Y9WidNzykcpA7W0IijubX
59Hn/VKmnuHd9ifsVmwnxKeB0ofsDzjWXDBiyLCiI8MaWyIfdWtAbgE0Vtq4+32/
vIl/9bjdIyyScZ96/h06Yf3zdfRtrSUoqGPtbnSC+x0QvvUUwpFmg4wJDNpgavJI
nI443oJX8yCwc2LQj4tLqyhaKm3vX2xAI+kL/5LP4px6S94C4vnTSTyhkH4uvZek
wRAI0zO0YIvK4f+q2YyfynlAPJKqqhqjjVbpl9YZdgMGv+RGKtd3OSD0G0SrY5fA
z9dRWtXXszNjqlwXIX23qeMM6Rj+w3hGPfYAOc4YCnAN6hXbJpdqXh712mKsp6Nr
n2ProUxkJAFYYqMAiyDfKTFYH5lLv+XddA7HFunk5EAImtFBuJJ453lOqSe7J8yu
Wb4N8mjHkAj8ySlDQIe9QvFB3591KyX0+tGkq0ykyz2Xd32xjBvqJx949gsiSWd2
XlIyq5JYlyIrk3bGE8nsccUBedlSV/yShVx61W/wGaMwj1coUV7lDsI6QDInXbzq
dIsT80iQb2Qi6GvshMTjPDCGNsKLhYaGbB9iPaXaQrUn7bbF145rnp5PvPydNQz2
iKJBw0tPIOz8P5Yh6sda8kjM7M08ajXr7QPN90e0amd6/ii1FxVEc/PUHWwJmht9
hr8RgQlzjlKpsV8qUM0uSd9gYB3HhPVE5bZjZ3NPoKOSE7fk5VFpYogeQb+BlQTr
SD6nQ0iVGK64GFWpM6MfIk0soQBEgu8uDsWT7GoU6bpHBsP7BIq/an1SETBsJ/ow
NtyadSou0CuHYmeENWWnTNwwk+UxoDOZhRqwAuVuZI6mkJXzsq5eb0yBbFHmTfYn
fsHHVhI8YZFCIcoxm8dxSH5GAWMLS9datY+Tqz0X5tPvWC+KcYF9noh3YHYpENWZ
4N/ow72gXNp6b9IoG47QFFF15t39piTpMvA7+B/tvjNks0YcviNERKdDOPQerQ2G
MPtIx16GTyBocvj6ILreUh22WHZf7XWSU7XZxX7im3aDTJrQFoV/OXCWMwJ8wHGv
jzMujo/eymC1N27QYkXCsdSr3JL/e4W7Ic00pEZurw4vQm1c1hRAudHjmVGh1nwB
gP+TsbFpX7UKwYSBl8uYvxceQ7uhTV9EJvywPsbmOKNEWZDsi878Rq54yXkG57Bi
50qNvcJ4MBFcyV6A+ZG3Z0KgbaA/0GUE+Kniq8Mp0KNS2tOJhx96XIy3pHaILVvU
B7S/ItgIuoiDqz6LMCu+RdygoGp9KHyc3nIWPDxqRTGJqkQM0cB+9+JF3ItXEocN
EEbHkjoOidqeM22Xh8JU/1ZOogUQLwUiqS+ZY3k0K7hM5wzubftv2sIWB7KtJRaM
HG/spoge5VJ06CNRs5sZPnBUHZz+aghWyRe08z9ZbQjEUuIb6m9lRZH0RUuitWEx
UvzEczdZ22CzU1a4JlPQhVZX12XHQ0gIbhiUC39BFbDhX+xyH+nqONyNwrJry8iJ
V7nbBl3Pv3lWTg3QxcbPDYYIxic7yB5bhp0TBIgkhYC248AMj/CT1qdtPbBSXSOr
a5Ab8Tc7JV7nPpTh0DKIMKVDJPzp/4LIVJFYTw5nRY/NkfhTO+nprKlvVGMFNabS
mSMCZ7cqKmkxffbwYVIE0fZoy85C+dn41m6Yyrmrz5kOL/Z8R1N52CoFbUef5QK7
XN/k/I2gP5DUyNQRK+/nnv4i3808Rbwnqg2m5+WGejsBN4Km7NqhFvbcAuH5ukeN
Yq01+jERVQEaiww5jmfGmYD3+kx6n8uyYhobl4pAhuXHEKSP/RDN91nYORRnfPSc
FFTJ1LQrJpne89cDFjS/kNN0OXoErC9oRcOUK/nOvk2eF7/VNBcycqBli4U+gatT
PuFjdh+wft/9q20kGeFXHFzM9StME2fZ4GDm1PmEUs01sSRgN0FmjlrdQ/ZP9E1Q
Pf98qyBx98RX4d0cg/igWIAleljGqQ2lJDQFWKTIvbYMOhbgfwwFEQtw9yGfjwOL
ERz8ufaiaL7v6VltNWBDUXBF9lZHWJ/wsj2DOvCNK1tf/ozsgYZIPWaPcihczNj4
c0Nq3QizFz7E34J9hUO66TZ4NfFXjkHu0JhBHNqVoan49NsOI/h2dtvTvAhYvQ2K
KONP9bRtia5HGkNNMR7jaNibrwQqh9Uq+ageiCtw2O7Y0Y+7F4pNWy5gBX/Kww2s
VIqdiMaEfHIzN98VzuSMvG2fcnOcDq6Ev/siSleSF1mSICidHGTP8OhgHRoWcFCd
1XtrSfaNQV6xkVEu6hfUlL5DyurDiYRsw78EZ8xqLeYecpArOckIzFu8YwzQEdfE
zqkZh5FpiOoos4+IwSNE/qEnFwek0AR2dEN6PKM0P+JFAlpGaka4Qe+2hGYsMS5N
CRLiOuLuKDYNzzbrPML4rO3W/4Dv+kfLPPmGkGZeT6Ih/c9DiIPSR5iRf2who3Xe
AqpgTGABRwM+otiTSCpTATNqJaNpTLt1WZm7jNKVfMKIIacQKBqZNkqAkVrfw5hK
5oGmbd4Bfb3BdvTpgWsmJd5+ogZ0qxe2SCFSFDiR0D0Yjwe8uhOPneS4vMh0FFgP
7tCc0sGZxRsM8vIzuNlM25CysU4S0P0IJ8zIGQ3zfcWQHDH457wYFVzdkj/3BqgZ
LTBAR97typ7RlA+Y5wtinFSBzLwSW5rvOoSvkbc3GXgh8fHa3npJGWxKsLJmVxci
pIkLFpEhOlEYTnfCJaCbDYbZhp+XiH/LK1aVXd2q84AoSb2Z9Rw38g9eyYWph4GI
7wpf6k/D/ErROHbfuC3werxxb32h1NNLq28nwtkgweLLnCss/Ij0KEXwDNoZQCGs
3rBDo+XUUul4W1iDeViVtfdbIY1TVrIZmMo4WtOtFB6RiPL3jpyTauMTQ0gAIeQ4
qpfKlftR7UTvOJzGxK8Wx1ufSMe4Qm1XLKL8ez4yB88eTNhBCrXwQzalDUFHJ/w2
TS8ZkGkU9YL9/csMYo5LBeBF8gnCVZ2tG5z5zSPiusnArzAV/WRqwxpe2TH7L4dS
o/KIM4wI3e9oztvKqghxllSJ2Nr+dNkAkIjJLvK2c77I9kQGyZ7SRLELhaOL9qJz
Stkks5ASv6KhNWrvQo5ZgFDif71BnS/zUgPqqizIO4RjRqWODl556mgIgzNTa8r4
LqaLIdJZJW4qt+bHrBpFwtqEFzR6jS1Dr8u6mUiPPIFl5wsZfAXbg2FDTlK9Gscr
sTyvWNvbxge7OTLxHrNYVmGHa4W0yw/EbZdbU/BOhKMe30aeUlcKUCNElftfHpz5
y+Rmr4bQQ2kCdB6W5k4R59wkAWPd5hYzy6k+C4sBL1HtSafyo97p6V5tgmcYkngD
jaighUM0x6i7qerd/6fRtmNLdYGpw+qTRT979gLaS3Ok37AJA5mHXd1gUmfkdQ+5
0XbaYyUKZhSi1ENxq0yJ56heo9/NvInNwJZlZQgb4x+y0URo2kEwRwsXLoFITR0i
Ieb+FgxXCS2cIPGPMLRKT0ofroNoK9AtsmElyG1aXbgSjDrMA1TQa35WcX7uzDFC
3nWvBVYksLRg5kZR9moy8ZbqbhBclQHpPk/Jys+8Y6LPBMa82qhSV6TGqk3YvO4E
WUdm2Pu+yt5kU3RNbBUV/iu+fOENz5deGue4VfbjMpLa2eQUIXtUXLsHZwhmcVtP
vArLSZ937085KgjlIadRqyA7tXKl3WhCGtNkCEHAb/flNGKPKdI0wSP5OyeEQd+o
V0OWOb7CbYiJD+e96NvqYKKhlx4hCBW8zmTRqmeuLo30dv0/FCujMYtgK/jHStYD
Qkuv+JSvj04mCCiuW2D6wDbaT7LeITdVw3XCaGVYhFflnc0L059E/sE+yHnbWwaY
jjw+ALIiD7zpSfVe4aCDXqvyavsk7vqdy0+vVD/8T8RfPconeTpfqKdtTL7Wplnp
efSu0riY6yOPwMdTwrV8gJkgWkDaqGSCqzLWpfnX90H7TY5p3ZMKXAMxqBU+2rSl
fXssFa+8jlPsB8+Ra+usXZYZ5bzHtrlpwq4kg7rj4jMQ7rAUp7RqhqJBroij4DEI
DvkpQJ5d/pDPy+gNV+iWHsysuD1+PaXCg/1HyxOTB5ZVKry+Enc8vSTja/QAIn0O
QOnpZ7qmrg/2/yaMRSdcZX9KMp3M6hDDKv9Fq8uR34miftaXkI1QUYLomketkOnP
/UMHU4daXb1zGckVbVZGq3K7n2z0BZi41epad8oFX6SQwszXu63IqEQjXyo/HxPM
6yOq5TOTY/g7jV4JdgKsxqBzmgSRoQUaFiuD7hN62Wh20OO9efCeXuZKT75kBkwf
r+CnkgMyceHp1CJyGf9ozpego9IHkF+H7UQSZ83uxwKUqxRbK6+lzhhCdqFwAcek
AgbU2xIBHC5UsSEHhIygkF8Yd9/nj/uvs3zKiL3IPvuiE6sNlOtcH5SUQr68sOoH
//oeoogRj27KkcsOgKtO1Ayxwc5VjdgLZrPLqwuBSO/BOHoCRqHy+62i7RFZpB49
P9TNkmUv/sI0OrzHqdLXKXGzUknmsom5ch9Iz4XyafBmsJlC+byYFMJ2aU1RQ+K+
mpgaYAQssOSUbXdp5MWEmXqmCeQ6/adw0cb4wfuUO0Px8Qp9dTENC5eEw8Yem+kF
iSMCGdHr32Hd4bAVJXN3iYvW2I8S8gCKcbQ2/+zM3ypn2yfXgVOycqO/NEo7oh5S
leszAbGgDzTuD7HVIEVNpQ6vW3qwoFinb5K+RUcWGpMbbSW/wCgA6/0UjOg+FCQQ
g617JsZkY/Xt3Hf+61uJXMyPtKTIj0rT1/BbJ5zYM/7nH/DJFflkXcWx31d/1vay
pmRi0kztKk6VgtZMcBHWrUnsq16oT5ot/0309mAreh0SAEIf9bQ13VA813ymmVLt
CA5p+w4TSSFtdH8fIqSCzG65SIWy0HnH5Ry9G93vJuQlHV2s/iHMDETXeM6Cc6kT
0FxBCcAE7uSOwrOIjCQwpzcLzFuHTEzx1tttLbvsJ5MOwDXXINQlLEzof5uRIxK3
10/ygYEHaY/b/8zTYThyUw8lyNqBPlMt2nWTGsDWNoqkVXH3xp55JS9E5h3ZWeoW
JFWDxjmqzVNZKAOYVF5wCVth29VWk9TgI8PX0On3vgEqYPWIDVhisVcYX5J6KU9N
PaLIHasSmHSF742wlYo89nnkovVpEZGwSBYdv89erMxHp1WgYz8Xf2wu8GIOPh8Y
eesoUxyrG5EQYEGJBQoHBiCVk4P0dZF8w/sIQaqakgaTrGaqJV59uvf4o5yaqBAG
z2gWp6HBp3uVll8ykiTKBUZIZH0UWUNpfKvii+AQ1EmLeEQOJ65XRrUj52Kq3HKP
J4kG4DrarZXDuCghsSaB9JvwYqzFEsEAASYKiB1cp8I5pBLjZLoLwiFAlUZkQOU/
iDA+eZzItV0U/ShEeeV5VwAYLwgEPdbB3ckgUW97f1D/cK0zVF1kwLyBHzlUbRN5
6fJJrNr/GnXEl74QZYSduxjYt47kQ289QyUkG0vRNGTzwU/SQBvWQWxXoZmbO7la
1TA7aGd9S99c1VMuCh3SsNBwE9jebU6oQfDoguaHwwMMk9RgcjsCbytUY2xg4fPR
1vfmGu5LNMuvbiLoFDhu06L6bttvqaNw7OQCBQcOvZqyMQ1Ugjkp0AgQcVMZGHPt
lmn4uFtJW71ifLKTmrCPARRoJHNCAnVzuvYsAw4tp90+Fi8PDgLM4ew3X6UXNOQR
XZqDORz86bpuTx9rJUbumWsHIGKgjcASKq96It4gxAWhyba40bO4n3Nf57KYjf0/
zNOhjCYsVbwHjeyy2PCrw/t4jYg8sqbGUjmeDIz7058EpNgXXLpwl4HgFm+7v1pj
rfRhlFlA1+ECmuocFyacVXoA2lbZe7ucwvsLOEWlroXQCMDPCNNcEpdjQLhTFxYw
UZOm8DbiujzuHBo/9e4CFw==
`pragma protect end_protected
