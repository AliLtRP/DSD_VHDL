// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:34:00 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FRRRXXV4rw60yyJPHE6TaTBWbN27nByw7nxptYro0KD3ukFy4AHr8h52UAGgn5bo
YMsnpHpswwaq6jCRaf0D3l5VuGiL8L/cWlvW+3dzVEVNwNt988bMnHF5rC6uBEt5
nVqhwW57Hz3r0/dCbR3EqhY2ykiLDGbtvp6lMjHxpN8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6272)
NewLYRyCFofb8XT+TdF2rcHGVdRaU3h1W1/1WbcQ+MuZwXmG8Lz0v6N7/NmcDUgl
tuP9GiBwWchNwfNTBKKS9nygeRT2X1sdQ0HaiUT14D2I77Zb5iwSFjGmEcMUJk5n
0nf7olu/RGmENHqyXVrfrQmJeoZQ7Y6EepbiQZ5JltIVNaEjGLER/horVzqN0VDx
SCPsQyoA0+op/m1+v/z3HIQhzHYPumfM5wFQEZmGOcoefl7NxfqAuoqguEV5J5o0
i81+iZ/H7yYP28N2FTzwvq0DIMBmLB+CJ9xEPeN+2NwPydYwbGrV78i1Dy2KDXKD
NkkY6kQeJnkAMwU3nVULm/tDuL/4kdyb5+UAc7Y5WWfXeVfbOlrrR0oQxXHztqoy
kZoS7cxHe57fMwhEIUqezDuTMtAoec7dVPpkqJ3k+0+PRKbkf3PrZRraNUHtzK3i
5F91QUNi6mszoNZlEie8ECNRZ8lXK59Qdr7Ojiv/TIZTepTUqmYNKtdegza5nf3e
kh+SRHjwYoT0qHuBd68gp9p7gsfpfTgNchD5y6Nq58nJ5gG4LpRulcGWyiFc/M+g
HO+iyNrTY2c6Cq+4PGVLO5kqcwz+OuT7PC59/a9FiTxpvYlcvvZ1x7nRGGc6cJ2J
0b94FzEIImSSoGhZ8hkUVk/eAedulxOcNyKnqJ6m+Iw4rbGOXGPipDmGn9MfLmOF
6j8Rlm/j+lXz4fZ9hOthdMjovX8IUUPQXkT/9uLRvjehToeKLcJwaCefRwBoqUck
5ffqTPDMEtJmfSVq6dre2aM27+PvwTfo3mL4klgREKQlVNuUkZmPSaBg+DTSAheF
36tWnK6Q/TMLthU6LxvEc9r2+AwBuMvmyBOimNitp8T/pvXySeJZGaVPfjdJNKH9
PJHeH8x3FIPhunrBvkaKt6rmhvk+qpkT/SefHQSLmSMv5EB40EqIFwDzE/EeIPvq
1EOk0sDzMtHTU3N2FnwKFfdwlZOxXtNeNQulC3XpDc/bY90HY/iNlzO0yiGTNjN9
EgmSN0MrxcZMWiBKveYXfxfNHjAPpIF0pZfiEmo4GGcof7sjD7sI3uSkkYEQXqIT
XfkrZFiGQDM3i0/pzjEdTWaltVO5Nz2UzLQDZGxgwWHpIAXcl5DcWXPkeMI+zaHj
+fxAZ+rTscjK1dgBUY0Q19n0lzaX3zVGDBJM/SA0UoJxqONdjnhi/MLso6yo7nm+
0c/yNcsxf/bzuUQ5g1AtRhe4ziCLGfkh/UrIOuMR1brid/pHc7qTGbgAolBkwCrr
Ym3WGtJraEp7uULxHLWvarCyLgF2uKAV2NdYpF7bXpSnZIpy6PY1/7KXgYjdJwHf
unHUABQTaoucCHXpiO5kv6UMwEG6cj23udPij4YTD2RW7iG8IcH4TH32wht06NFD
NT0XRQwr+blWZh9M7ek3v1hy+gV2kkSkvuWTH8pIDE1Da0ILnOujK5ZFcN+9Stdl
2xmhPELqQW5z6NPSE7FcUAIaWnS2K8nOz9GjhLq2S+LjeJlzmsxv5M97FWd6bVE1
dwKMZPRpmA9N7WZCN+fy4qW4fNAXMdexq2RqDhEnB1glC3kLnHdZxnVKM34fMKtD
JBq8+pI5v5iii5RetUaqloPiiIt8zI1hvkCLoKpfzCfQhByN0/ERwtAwfLIUYTug
gcQ4MN2Yn+fZal4UjgU0MA6EQkvZKtjFq/zL6J4l8E0RZy/NUl/Zxqdh+OztDTe8
mIvET4cCK4F94dRuYhd52mN7SKXcuTAMfH3hE7ik2OudxVZcM42/9+57RLzv/OK+
92/2AaS5dDChtTGjEnIgOKm0qTWgYHadfAmSrAietFqWxizvqqPn7U3nD1KPMj/z
2o7Dr8BLStmUSELdlrVMpvudtVqTZl4Jp9dAsL8KP8IRMkZ27DtHJxqFTUGnLBUt
hhPwOlVaDv9ydfDzm/7pue3XNJu4PeyEP1iXhMvyFskHGCv2NIDuIxd4MvJd30II
2Z3pOWGv/Bpaa5+JIax2AmoIAn1Pjz1fyLHqkx3Rla9WXN9xTt+BZ0SyolZRnK5N
ewzieCgNQTruO+is20lwxrmultcrtnMx4C5SYBt3K1CHqRpMCVbW/3LsVDD7Tkh1
jHA4xbFCXKjEmhyOOEnmAFQTyQRM62H21O9KE79GjP1XO8YhMAb0yCKhDeHlVkSr
NBdNZgiMBbllOZs8dCKvQCGCO/uCmDKxSoOhiqzlPvQN9aEGKjQ0iK0AvHYO5FbR
WaLWA+VuC14/iFwnOBMPg1ybP1nxVnq68sZMyLpJBiMTFc97u2M1YMu4eeCn8UF9
ItXpb7aU+S/VPalr+na1jLo239L4Rikte/Vgd+5+SG8hEvfX0ILuEi5xxqTdF23K
YSbFqsroQvie8nEhIGW5CQcCcTtiU42Mw2JoY40MG9MlGJ5ovim9VviMVXelwmyI
FJMjFg6/QnA84TVfwWKmgUl9qFP4ALLdxyASshHmHySE8u9wxQI46gXS56xHJnEl
oxqjZOz8eUOKvNkay0nR6xyHXSJ/RbRQF7uOAT2irzU2q4CyotvHjpPvxfiWy+PC
G2EkkvL7gEfR3bzw5yT2FVxMkVGtrnTZ8VGBvLOktn0CnPvS5zcVY5mGWvukidpE
lhh2N/esqFQy85z+Lb2mc8AOXEJTiPTxF2LPUgsP6uFILwZB3edKHTBAga1y4ANf
BgqeJ79CiS1bYlsQwkI4jMK2GXzhHk+iHYBUwJZu1LeP2Ic76orNxoCRUj1l3KO/
kS0aZYk4KSBcSzo2Tj/RwPOp8RC2lSd09H83n7Mmpgr5ecge412hlYI0TOJUVg4v
btMrSIs+0uKJVfXnZkLHfKzhdy1LUFdgoN5N7YOAvbuc7SW61kJkwNLMTONt4A9w
iJbcpuFO35x5GLxv7bfwLEjy9d1Zp8sGabDlD2lL8ysyyMII8+ufvsvwxIY2Tp9/
OLToYVFnf+rVgW83ZssvrLq504eGRNvtL5D4PoEUZ8kVENrkkpLn9fFDksjqtUfY
wYP8QHZ1+Se4SvOUT0cUyrA0ThCTXktW720jURV9v9uRbSDLIoeeB+WdnwqTE2o2
9L09fGY2mVrp4Ve7kjtp3ScUsgNGauoDtzWjS4TOtJFblP2nRyk1bZ5C5U4wicOc
eD7/X4o2HuZ8ij4ZAKuWVGpYFzB/+0In7NfK9+9NiJM1gAh+z4nM1fn94JMP4GnN
sbqL6sEY9HOVrAuYrYiiU79Xm1AOB+6+Kply7RqWOKHELw/hKH116P2xOneuAdYN
bv3RRBY3B3PpiOI7xbB5zqdWl3gZc7UVymKFJ1ziF68VIvyRYu1IOPOwjaTz/4dz
mj+59mfQ98vAZ0Gz9yCJI8Ge7+RXPcO7zxyGYP1u3R0YzVPQMg6bXk4SUAw+LihA
5ViGSKUARQWuiRk6KhoqlSI/SK/bgTTG28vjS59EF+HGBqhgAYRQ4YhfZawwQItM
LDBZf8LRfgqQieyDnVH2fzzTvbecJnNKMB2hUlMX10FhOSNPpUCREt+hN0YP1xYT
x8Ceavh+rdAFfm3Nf1wpkGwrais7S081Jvo6F17Gg5NXreaaUa9VcE197SvVMF3W
AKlQEGMu6RGXSRMbPgBaJ3HPg1v4r9Po/V8eBp05xexVGV8cR1t4q27FVJfaW7LX
NS9bJT2vZgH0lw46WyRnYTcstW5pVWRXGdzoetIsYV2ADgZaUqMuOcXocvlCB83Z
syb4XDusPqrwsyUA4eUKPp0jg942zt+5bIDd5Acuo689GaFKJBRDywPsxNDLL55N
/Kd6MZj3pwdGq3edf+gjfFw5Y2WJSIxgRp4TcJ74TLezRDIW/apMjEacoFuQ8OWQ
2nYVQ3a9z/T8rBsy3O1kXiivZAEb/zPhoQk9DYokyjq8lAmYLmvfs7jWzMb2bKSr
tzxqV4Ai7g0WMAYnUdjT+eP3keCK0TexA5KgTf97b+gHv8SSFOb43L7TCfsdKVdI
JpgHKwM61yE7EbwTKDSe1C+jze4/R5Y/vViI2wABy9/jbPrC1sef/wHFYqyz2Cr/
jOXbuKlA21theehp/Kevkd7DzLcEgiBQX7OozO6kK3tbJzeNUziIfPAh9XGTpDLw
8TAxrzjdvQhzSqNh11gHhrqMjIpoZ4NNv1SR7tkPr+Llnoyq/Bz89YmlIRWPb+4T
rzBrIaR1KEqSoEp3yp75pXGKECOR9QqafhwEM63X8pHMW7lIhakdb1NlRfetS10T
rATjMxrA3NjqDKWTVrl70b+OBDBuYj342Dx6HTQj2w5H1r2R2q5SLyI0k4Ud8NtR
PaXdkcfz0V2vNJ7auV+xPS53jJEeK+ItqQ/QrL97W5+SgZde3LH1u22GVrFD25rN
X4dU1owOdlvADKkWKFT2wFYHf3aEq4H1UBhO4unQgFYtbj2kzt4t/AftCVPX6SuN
A9bqef7Dqpmvq39h79mK2ZNTPGFAkOxMmz18vF0zv1oQRMsPar7gMgAb+TemrYEm
ClTBzw/tDpeeI3qMX2Z+mycC7UKpA0dOo5jZIr5/SBMy8kD30cgDU8FoICm3r+kX
6eFY1PWiqVomUV7ZwQz0lZnRMZFRx74pBv/hTmNv2KuwKJWkWH40j2+AULQFmDLg
rnX1ZUh6VhqRcFz5Dh6MRnUV+AyIeilaVYlnOfbMyboFXJmRB3xVjQXtgW2MbZO0
Y5R9xBvJitKffAuaeUs/odNDDxPsigr2OvGD3j1HM/cg9oU2HAOgQ0BDfEmT5Txg
gAT93tQvAGc5QoAr0u9EmWjzHfzzJRVUH/XMMwoj2zZZC/kCQjs1kaxomo8HTB+r
4O2zohf0kvzsKQQfLIY9GMVaLrTlvnRAX1c7sQb2Bi52PvH4bNo8934OUkbYSi41
9LGP8V8LEymHmFzj4Q1WPgjOilVaL82BdtdVBd1hXYLpJPqyebXxI+l68mamXXKI
HJSPFY9kWls9pFeN+VqFExS4YG988SxDzMj4pOvI37xKwMS3H2eZxX1kNX4LT14r
A2nbZQwz1eE3oHYV8i8P4Dzgm2SwXWMWqW7zh7tjYi4p4nXGs3MEgo8TsdgwCY0G
/iKSOAVhOSjcmAaCU0yAa7rzACps7v49LP45iEUFANVomVfy4xo0xzPbIuRbO/Sz
eozhaVbIEbR1dPVVikBOUXdx0Q0YnG5nKRYQScErSNKdOoWFP8C1qq3X7+AI7/lj
yu/MSlhOeFWktnziBy/i9tbZIE3U/l1jFtb+MpCOLPcAzhQj2zMQoxvO5EdL60eW
UKwz7EnHVyuIc8vriPM9NzXneZGh6aFqQ7VmWxHmtriEt0DOHyQQYq19ZXmFFVBK
yMZiIydzT39sxaKtsMqhoc7JThfEH67+xUzK84hlmFIw8p466ON5UlfqY+XWHJkJ
BOPVS2LgLse+AnAhpZ90/TkvP3N/ACGj5NCwq/1CfRV768q5OYnXPOB+XmbUnFv4
yCzfg1aWbJMeE8Xdv8T4khtfB53e6JEPaZ/ZXluQyBkxwOxoLPy2PGdao+s2Tu6w
HEy3ae8PgBQAUS+SY64SRB18gS7fB8wDE03RNjIL2ZeCAtCQ6EgEmKiymLWLPkS4
C4Vm8lRsJMKydLUurTsYN35X0Ox+/+/bQ0HvFNpXne3948mt64srvYPLq8lLYuXk
hZS9tE1zkSzTYh2+Vox8GSRGMdiOmLbNWK13gbzDne6cWP0nm++GF/d4bQud5WoD
m8pb5zFUgq8wV/071+2Az/onrwd35X2ZEhAySjLFowIEysgQV1a+ZJMjvFclZs+r
7MDOuvjve69NPpogQ11zRj8321z2jqdwmOS6pyGriFBRKxsrq0XHndZ3Q5Yteei7
lhINGODRAQ43XE/x8+M3wDK1VwnaVJlmv4AgfU4wE34xw0IDiisZ4501FTKhvzIw
RgOvBmbtl3lOyWv/x+lKKZm8Ir3DOXkSh6Lq+c2qCccTBzproliAn0hROluMo+KL
4b3gTYOSf/p0VTIdiQT4LxTGhwrQdq0kDdu6LpcJFQO7zzjAdoSwlTSsLQUnT5Yq
tPORLEVu1zEGkbP05Q23t6XKOcgHwNA6Zf/3YoAJDcq9WdUvdku2+MdOt01/elqf
CJX8JNyLcUboOSmnVA2TuF0jXTqB4qPcpAgmd3262LzicPhfduLh9S0nkU3ErqXX
rulFo1BDgkpWo27Z7KYwacQeCgrMx3nV5Wxl1JDtaT245kuiX0R1imAE+RwDaugE
HGxjJM43wR3pcODRY4v9IRTt+nBpsT65AD0Hj9l1Qo38Srz5NfONeC87JknyBYPg
5eKRZq8rqioEcCq/kvDH3V0fAfVodMzaz0FJzFgydQw7LNbjTv8Elh6DN6O03TF7
hGAJK6yBHEj8f2x8xyfR/EGYSPUrbfg+Q8GSc01MqEDmRIo4jLAd0p+yv9o89M0P
1Kkwhu4vpKq4Vj2gunNJmEQGHtn5sem3mQKZaYvO5eVmJ77Sc4vAG6cxg/t/bUsp
0X5Q9jrjd3T5TtlwGSlxg4Xti9G2+CNgV5KyIPsSkdwteI7amUnYxtdEo7HV0jQm
78QGNzP7pM9ZCtXheHD6tU2y99jBQZemv76ZnrCawdp3wXecqHunT9kAQImSaPot
BtqRyNGc4LzAgP/1BllKsrZ7GOrdJY9ubHSueFUQrEauEOQgZy3wGvClw8AfEhQV
J7jPddBdgZJYT8+rMUDTVlUVOj17iRyjefU1FoB/e0s7Bg/LYhlNK1OcBIR3xuXl
9ORyDI44sZ+6rExB7KmaX3gHAqQgST8sJkOqnS8fe+xp/YbqU3nO413Y2mRzn44I
e8Hdz2KNQA7ccMyTKSxGLHSDdN6IuYif/ksoL0T0LcrOJkQoLnB82rHmVxGcRqG6
kg6s+xrgNyqoNYc479HdDL35FxuX0eLlzAHLdBBQ7k6I+zhIokSXb5rIglZtHbAG
Tf1aa7vAJl/JjFcRYQrBkI1eK/xrdnceLcdnQ2DjGb1njbUvgibrpBFMHH1K1XMT
TGWintBAWA/SDlMOyS+Rmfh9Xe+1Q6jsxIDqhrDrGa94dH/i2WzXtMeA4RsVqV0l
oNJWgrMrTnq7AXQDPf+KcRdDSbjfO5+s6XTYnaXYkzBzM66xuTAxIvht4aA6eb+n
XpT6Zm8HoCZpXek+nPgXPdOi9dfZdAbFUFdhudK8cReHeu/56oMWxLGVcSrkRFZi
A/BWSZRkkJcsIYwxFXW/qmt7fXI7ybnJqAP7s/1fsVyyygIlRVpWv3fxCAckbozt
q6VVPj8YVjclELQwcEA1dZ7SC3PgnNYLjxtjtCsO4u7rKxNFvteR2R5J+kpbV9AQ
dRtavmANfcqZJfrviti2HiR1IaP9H0oPr9eNNAfWz8/RWkyheMTAU0Fw9rCdFOSi
UmrPDkuNTxH1tLxSjgor8Oozx5ytuIlDmPfo9LFWbjTOagRU4A5T6jh6ebCZisMY
dC/qAkpHqEiTZxHHEQZ7Gjod8bOU92PKXJ8uJxQqFW08hH7f1tBeNXlVdJyjrQ6f
mqGiYM9F0m/1ujpGF6VzYB+eN4mEHpmylEA05W3aR31qBu/Jfwkjh0QmUsTOH/Se
Ym4mNTuNbfItzl4qq25R+JTdMfoH8zoJui08Kuv7CfSQRELAFxhDG2DWRoOTQbQQ
2O05I6e4RSdYWZUB71PR7wStTMtnVtpmSpWpxZCQ/LXHg7Dh3aA51t+6sjMLU5vj
amnEanzI8WowWOjwnJdHyokKNaBrjY2zSvjhrAOdG8myhDngPZskWN9dle3weWl5
JHm/RUQ1xQ47XCAJ+2gpos74CyUYyd1Wg2/wg34HjoYwcJZwtrG8sc7fIOQ2C2kx
F5ieC/dKW4JOi5VnhoKBXFyJ7PbGEB2/c1AFhKCNofWxJQvk8vh7OzPqOrqQRJfp
U0xvSf/L8KVCl8Crb3hXOSnCLPf0cDsTy1jRpYDKYrlAOtCRGTvk4e8dPdLtKRDl
GJpmEzcsB82y2471+KqZJuUT0/eV6oI9W4zTdoBzK6e4LLOrwD7OiFsKQQmlk+t8
IYqKgCkFyPaw+zUTC3cma3xnnIAszS60a3kwXLRomokzsN9pohCJL1chDy820mUs
nhJGZufCCrY6szWMuRTl4cjP0nI+6r/TVFLi55sDYlPBVntPElSRN76Jt5cNWDRJ
Gk1wKSlk3/0MDk/FtSuuoJe7VQI/u9/XT388K0WD0ao2o0nOyl5pPPrziXcmR5Gu
hjNM6dFaby62/LuCzfsCsk7yF8iX4MENrYzeW86XX3HXUCWJpNlEvqJ7Ypj4p1re
f7+vLfJ89e4hqdQoAey/sieurtvBI+hxhvaQECyP/6f0WjRgwHrqAVgCdhaDtyJr
7+KRc5YTBoxG3U63hnrZMG/MAmaqsRGNuxzYxIpbROU=
`pragma protect end_protected
