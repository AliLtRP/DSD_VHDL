// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
a3OxrtZK40bgunPi6MXDWxfRzCX39SmHrYMEtfSIwxXI86AG5tVIpSNSHDDzGbX9
cfZZw2ksVJyyI76scBPfooBMZ84LVSVqxh9ie+JKZrsGIY0p0WQrrfhbwgAjx9D8
pzEesihnyFOkVhy2k3o8gQ4sDgo9gy0IN8EE12VLEp0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26960)
aNMDniL8y7rOiRbmtU6kIqjuvmOk7iBdWawv14iQfvA5rEczw3RlpeVlubTJVWIp
5VIL1ysKNPLFGORR8TDcWzoHWJT1RQotjz2qqJ31DcVps7NTq8wVvMy0AzdNdr+4
SU0gh6DzeSglsrZJ0ttAwAbq4VX8vxtTk6S/3l7o2uK/jaymRuclaSKg5pIlEWI0
ypBVuRFCaN9ei8i4x0LNGGY9/L1wWXG7upgT6GcI+lc9mdISdSdsz5BgEnQWt3a0
48b3pHZ9eQAm8jibAierNubTKwYUlV4pI7Enql9kMP8jzWI+fKsK7X7TiE+zi3Jw
4KHnEeo86tS66TiW0TTWBN1tjH3xy5IeJPtccl1x4FAAFjGl9der3bn1+AYZpTtW
v8mzlIKLqR+Pxhf2fIqFBNNEcxuRnE2+SzD+j0ASgz7XSkNdjc019lquHbJYX+ih
gWYoByNHud5NC4llryVbBGhuGUebnhNl0H5gGRHCwd7t/lweHHL4hIXGIYsYx6p2
2Rqmkc3PUVWhj04YOBgsWMGWBkUWy6yQzA1giAwKS6x7SM6yAz520CBCBuzjd3JV
9ZTnNy4qJ5qu13lXcZWIhfjpjdYC1bNv9a/VEnXzueyq1BRXggBHUbWijv6FFFLr
BvuUXxHhbCL9Pfic4AeCFdvnLtfPgElLni9NxS9Gmw4gMYiftrc3YmnQK2TcBlq3
NBllLQL5Q70BABau6P+I41Xz8/15PaaspbZrdmg7tJntOzdCQRPhqp5PuBgoC4IL
eGpaITgYHqBfuInWDIGnO7qwj4UnBxe7BGDhcsuUCqXOvhc3Poeco1eWXtcsZ1Ue
TFjsfJqB3xNiP/OjMnvehsFj3ZDDIapu+7wvIUrsb014phXQuapNCjlIXrHvqKJl
64huBUBjqbWxbgNxAp7b6o7Typ4acDza2K3AM3JQahfqG4WRYug9l4N6K4ayhMhx
HXXqkoOs4+nN9uTE1pdZ35XyD6WFnEaEuvN3H4tV5TW7xlNredJqgDTArtBqgqGe
eBvwRt11inhDwUuv5M2KEYPmXSTHYK04E1RaIt64NSZ+IO9VqpbPISQyi94GkKVE
FKJDj99WJbAMjPKqZnSG+PF+MfNXTLHBaXMxSs8iyDRIIwUq6dZuGlvuvuF6+aPk
DzN/4fRpqLprUiI1yu1/gr6gP0w28PdI48PUIeSA7azwy9lniOCBclbZyZ0Q3SVs
un/fWR3MW8k+cT/2o9vkjQ0IfXFU4K6d9TPTDBNJkJy6jfIQr1GQJF/VPL5FW7n/
svAnVWeHn2YCcOzdSLFg/8KuxQs+bYsNEgfZXoJxb75hWBYCpsHEk9lUX57KfyQ0
MfnWKzhEUy0l5i+iA//LBNYn0HjWorIu31EuNDKee7oCkmUYrwSkIqddqdrjEx7F
HJWpLY/vD5AM/VsJhY9HnCcMIF6mg10XB/tEcXtGm9pT3nqN5DcP56bvZfx9NyTW
BCRo0n93uVegbC/CDiXvgG07utCWZC3zCaOZVbp3DT8kap4R3l2OSS7/XApIH49e
VHg6caCjdQwU1GuKry1O1gmDbM7/xqQggvPY4JGLUN28z1ObzMqmEsHs992kj/kV
wyoLtZOS5e4+nluBZaZgNDSHP4HeGISqbVfpVy+Ijna7zy9nhdN2H3Lor3r7ZtQb
8z8yZs8UAlVZgS1cWstAtdy6LE0LUXbyH5/u2UpwjBqFo0Wpz9r9qd54CYkqV4xv
Z0Xo2/QOCuDW7GsPPmipJW2DjGx/kZ4SzvzIcJetzjk+Av7Gw6C8Bk+luIW1DADP
74AjplZF3As79FErnRDJU289SzVIbxzJBG/Gey2RHdVkZVgSmZUgDBQMKnv+6kjO
w6i9eIzLdn+Ji9XhMaq2oLG+6U0cNNCPq4ZxXFD2D6jhOlmRnpEgcyAWojZzuIMa
mFn3psnqJIiKasT5YrL14aA9Lf03n3QeykhPDYkkIu+zuv2JLaTlcfzraBfLPs6o
Sv9MPC36VOMo9xLORRrQCwqYbqudRXkZ8VhlKCQVvHjNgjWSlCmG4LDHMNAdPJ83
JFhpqweB0gyWy0eoZslN+qMNOcUPHEEtmhHnP0k/KAXms6K3VEl5Cd45nP5xI3WE
qt8z4uCi79d44KlWLzIlbD+w62xabjcmP6wzrODr+ad8JHa0nk9vaeMGsFaH9ANZ
coK/UNBlamrtvNWmg75fVRpgzZnNqfV3KCGZSeG947WgFUCBjZ++wKkCWHwinAYO
qhl9jS1oD4hFECL8RAtdcy8yEMz89N6ypJFbFklkq06DiulOAcxbFWoqBf36L25U
ad01MrWz1zsJXYik0MX6qFVspRQonjd8YV6Mt4U3+k9X8kC7ZTsWmfKpTjnNZLEf
KQ9bFVH0nOIDcs5jfwhWKYwyfIO+3E9Hq6dcfpPLII9EsOCS2i5SQHQI/Fg0NZM2
voHhBHkXKEkL8ZSGhn0IbUyaN+oGYlb3RQX3Ipaxj+2GP80dLsAYR2FwE0NTPlnI
4ltiBjYxo3FvuJc8YFgOc/RxgJ505V7MF9ng+gwumyl6FXLwbq5Ntb6+eyj1QioR
q4I5omZ/0i8qP3qGKQ7rSfH7zlD7c+mA53uJiM7XA2g7bQVPdm2mNpvgkU4KLpA8
58Pfar4T+8t3yBObMowWJZsNxH6caAFtxN1PNcchT3gscd7YYlkJ36YPlwM2BS72
PXkqs9MIM+1jE/m1NDjPBRCwzJlMQ00vBT7aPBUKwBx5e/v/tbihUR5ibXJma2rx
KX0eLK1pYmtl6V1ZOb4Z1OXGuiUQYeirQQVLaZS2/GdOIdTNyt3Hw6jiiMcMu+lj
jgBVwiLgukOtJ4rLR7emDLJss/kBzQjTQJuvgALDLTxZiKcUm0Z707foN0jTvV+e
ZTqwIes55h0ht3pDkMtuGFw9aoJpRbvJ3puirQLkCw5OFV45T7GFK+Q7b1lN4HDL
XR+GpDKIQApP/xmCA9pWHz5gvPOcHWUwRkbFXmsTP5NOO4LJyhpuqvHpsRv/3pFE
AoKMTTT+4AIgGj4YTSK919DoW5+XMF3BNaj0DbcgqQyoncC3KnHI6GJA7M9/yhZM
74/67C24IXhIjTk6PY279cOUhOKzuj5yI59q0KtElPX/b8R4vzOTCZF8DQPfy3WJ
eRdk25BIhNJU2YE7D7+CVnlan2N9cDOOSwEnQHeFfdb+4wjkUeUzHBf9TX5oTRQ4
xBczzc4fjrWIJG+OkMjag1v+wMhAtZ34yuwZQh/tWDsZoCx/t3sOBtwoWhh/qwRH
4buvzM3Sywch8n5g+QBoUizCBMsBBoKalLJPBhGgN50fE+O5ueBhcMqu5GTHXl/q
+YyKQFDZDymSgmru7e8bDP9Z5UjGeenUQBCKOoLUmp0/aI+h1svcc5Z1lLB4f+6/
XE5iwxtbSulSyIkmqX7vIO080Hm6higu2oIATyyDuE2pPbi8E0bz2pDl9BRk1G3i
9hQhxALXXkGJQA9aYl/q+czQoXVnvacVNUkEGXPZhDBCWvWFnaxj93saTvyBk3lg
w1uVwPwo/cBEu4XJxnvb/zwyht/lbkElxqwYvZ1UVqXNN1XjVKOaDfmdm7mnkNyG
22y/5IKDuwspIcfKtE39DGAsF8D0PxkUEDPay+734rmN48qDL52ebQUp8Zkfl8js
87LhfpRVW6wMCb0/aIi7vpfGBYvoGBZXzEEj64HqpSyCQOWT323LN5S1QSq8D1PT
T+QyJ4y7ks15hAGMx2cpLwkU5amFTpzsEaLX0+phvth2WD+WumbkVaoJdOxyPqMS
bXbraTGV6+XnDChH5hPt8YXBLBLrrUn02HSMXQYL2PT1L4h3QEV1RNU63BVF1lXM
mcmyYERWIdSoYphxU0cksy9W+IkImA7HGK8Hh5Hvx3Sk41n/WCjug01MTcYgsizF
YuxCHpbKs7jkVscv/zBpY7VzzjjxHrKZQrcA+nUgJ/LU3BjqXOUghF2OsTg+PMG5
y+GKx3qcfEqnRxv2N7UVCeh3uxIqZQytKS7BJ7fOdc1G79jJfVLeD0Sunom0E28M
sYZzRzkRRAYaJ3XNoiG8AHyYbO5r2cMDNRXVF9XqhdEgoWVCIybrxao9pOf6Nem5
tnow2JNjyBvYgP0hbh0pDcybtlxqKWhDhokEuGuMMOrPvdrDRzGQFhFmO2Kj7csD
Qv8ZxxeOdM2Q8YpblITD0OLos4UtUt3oaHxIwFshgKB7+qZmTBW/nWnmYDcFITsc
5eun94bIvH4NpJwWdV6Wh7ywWJDJEZEWUicn38GF75rsM0vt5fPpMH7F15MbLFai
xc19T/vRCjqRehnTtWtziHW5Am14LhrvLjZmZAxZYXSfyhDI4NxYp7PggxlRvJr5
mBXXYlMTdrjkl9tAayUNJqenExD8ktyNUFdpgVsmQPCJIFo4jqAcW0FHQKiTAOP0
akA2ABsjyrnhiBP13X6UvP8gOe8KwNNPdjwo1wcD/alwEFnPvCNOcFpjYc1SbwTc
LwFZ37spomKxme22fTRVf77GyOWT4at5ROMk0CFpK1JzUQaWukmURRIbmc+odoZg
yqX+4zdnXrvIxkgGAhuCRklRixbtb2T40X9GGIPLfyhE5FrJ3quuLo2+jAORGIma
23mCH85OL8jDh9jpvx5LOayDFqbwRMKIEJRnWBXNCuwI0St2AEAz/CeRDbEFwjen
SIc32wV1wvtfwoB+j5GaLqzfLNr8Q6btO7jWDr+/qg6qIT1WgzaRpNQeDlsxSNQ5
b2JEaFHBRiRdNBUwYccp0LhQM6CnoowcjqenoSqSsl9UNKz1e5wmk1vIKQjG7pzO
I+UgAiHXd2Xf/yPCONaqe6dxdw5jGxAOQUiitxAN7QsKT9rka5tjNf2GTZVvFARm
ab+oe77MOwHuc+E1PTU7oK0UIIvJ1c84TdwlU9riRW4E5Ri40M2JQ6KZsOqd9KwG
kZWn6OWPuZaIY8FH2x/iVGFVHRpTB3654nVECuD6dUTtMJO6T+RJndFp0cNp2H5R
Gj8rbEL1OoxSV+XgOZJ+yEu3bO5UAzTIw9D8sYXFi0Vh/FQB5GpajG09oibVOLXQ
eJcS4dC5BLp3ZCU+0VVgyE6g6arKEGu1TVKEFAKpGnizrVDMdZTPICDm/iDhRr6d
6jL2XAym+L6pEVSzUChXPRpN4W29JEwtZo5kMTWzPoHgXcVjakfjptvRwWmIixYL
4mVG9jLKYvVMNwciV6ZqsIDzu+dnc4F0v6VABGe2yyrFR3AM+Na9nn5a//C2KAsC
mOD85q41Hd6qk5GEcSfViOwzR+cAhbr49cKRJyTe1bGa6dBwjN/FSmwQec2/e5yQ
qYSfkil9Gp4HGLNIeRCFsAkykIs62LG644U17DdkfSLJ9MWGNFBQXljnPtqsXMKV
lrea2oWtD/LZuZzdldFK8eaL2RUtm9XFUjcVVjBJqqZa5+JiiGeuHWxtfF+4qp60
4l+irtLIZ1mEcOeR3s2ODMauoI3JpsYAW7YybPiolIrOMEgwh49ZnT4Kgt8/dufW
lf39BJ8c43zrWgkXWZRbHMGg+gtU6r4/0MRVmemiigLM4/GBkIrrIWfFoTE0qy3K
3QIFFFNaUlpn47Z95gGrObgZ/IZgOFvU9s50J1wLq/2URXAgjMxsatW06fBePgJ5
Cr1Ci8yygf0wXCnbLnu75zIXaZXp0xej9mR1rkoCr87o3RDHto8XpqhVqG6PDWXV
emA3prHVw1DvJ7y7HSFl3IKLNW9xI5uhxZrXC1lSV7uv7Wb9N4JWCDPfGNMoA2Iw
qGLT1L2zGSEmaWsB+TkJIw445DmjwcbC7VNVuI8DL9NjLv3vSDy1Zx+IF+N31GMe
Eix9jNe19X5Ey+9wRYM6gvpxMeEX+vYNaRu4nP7tC+1joQAe8+BUiMjop20aIX8K
7ESnU1TAZGtTThU5nP6t8FK69c+pKoO1LqlkEWPySDbVgjpebwNzFMvR5R7HZlAc
qZ5Ap46G4DWKlBKlsMKfJVs03FHE4r7WRz5DAYcrXIUhcBG+E5Guy/VptTwlaBBJ
sfVC4YfBa3sUO4oYYn/wWv/K2e92rU89X3kAzyBEFFQ0T41c9J8p8ebP5z0xomIg
ay2HUBA2+Nwwg9BAlKQdoJwPC4nQSg2n9PcOrp1qHboPLD4KM3bX4N6AjYFVKZP4
RUxmYRpWZTfMQlMYRaRuAo2W/kM7f0cFNZrC1+0fxd25YlYumROR36ZUu6Khc7wT
zn+amPXvULJZF44d95fYOjl+s6Z+XDmcxA+g5nYOVvlfs30OnmpklOSLiinmpTde
VNBUvTrFnaoFe0y554TQ8WxHWTX6Up6Po+m0D4Wdar5XVj2dRD2YDaFBzJ9rJIuS
KEBQnYQktXV+bsESCLdZ1Vg0cWtpwijP5u+4DPbbTcnnLLYhDjIZbZDl5PbfU3Cz
I1CkZa6XeUL0yMne6HT4IPyk4G1+6Cq6VJShog9YJHdOOSWBuYe/wxnVv7xu8Jq8
XxIP3bCQAvedQVClBG3gyFoudY830ilzqefg4UCA1jo8XB/FQqszL2ZxvWieITDm
BdXrSx2x+rxjiTtTEPbL1PvpHMYF6QXFmK0B/3qe7gsLaeo2gq53RUfvw/A6H3Ct
QV8OHahJ8gTEf0A9IbbxzcG33YS++Xt0j4+/sjV30HlJaKETA9BQS++iHxBf28Po
cZG3mHMImxTbBHRwkJjqR4WT23UEfn9NEZu/K0J7e/xvtENgPSu/KuAof3ioeopb
NDbHCpKQ1vK/8EQR36soadfNwkx0xA+6ezub7LxpWBzfeHuaLoEIQSznajLbx8Gp
A+l7jx6c8osITEu0SAwjevihkm6Mp2tLy6HNJfkVnoNXN/U+5+CJnAffeVdnsAmb
arEGp4cePggllMTPz76sMP1oXfceZuZV0x4JzK+JWmA0+S/9NeV9Ddm9IytZNH3+
pK/bRQeoqTNMKYcoezZu9iBXRX+rXU5W/0bJXX7ghG8xEQr5YEd6IaeJNHi7MD2t
0BH7g6viRWi2k9JQCuir8TmUQEf2nbkeZUSrHofRcpUqRejvEW0MbksQPvq39YNh
h05LZ6LjZ1BlSY8QE55EsI7kOjs4fBxO4z3+4DJ3aKt+5z8TLWakOrPo9cHpC+G/
9oh9qzb5ufzem9lqnIFV5aXqAGOHXyyPjgf+DpkOIpk1FMk8cxJ2DJG+mx5YrIe/
RipN9ETLr4MMxr7CHeJPIdjOtBFx8CBlB7YrQovNeEQOlEJFyNREvw6zAC9JOeNp
Ti6F9kz56nmSOe6s8C/Dfm4YZmVkkFNoNFZ1A8y+9JIaWMT/OWeftNX5gebVa7zp
a4iPdtFHCuj97oqW9cmoc7s82HriKyvypSKQqFlU07HA/yYxxJvIfwSX8rFQPDAx
zc874UZuynDTKIhxEGApReSmCOJv4BQvj//oOL6ITX/1GJ2RdE+l+OtfcNdjgFw/
Ct7pF4arMmXH4r/6mLCepCvL3i1+JJ+EgzG94IwYKdNR5hCoZS11h2S485mXtU4/
DyiiimycOxOiTuJlc0KrSs+4Dl7yddw2+7nuAHnok+LqxdmyIkuMzIMks3W5tvf1
9jvkyzX9MgKBbSbcJqdYCBzidv67Luv/z7AFCh7HhoPG8pp39wW5iUjMwBrJyllP
KUvTSDtRz8FWy11avV0vCmIjSmqmQAG2/IZ7jXXgQB+TKlMXTADo5kDVfOaN/Lpl
cnqWSwz2yog1w5tLL7GH0Bk8+UXPatmV/gFNuMExpziolXRPpyZvomGyjoBQR73A
MmpkQ/3vIW1CTfsNXtUJdImjmttixZYFvHdrxb7ZS8HyMt7VRbfJ8Fca3jl6i+pf
x9UunTpG28VLbzk82lboUA0uYFebpflYh61QLp6pniyVGBlS6f0Ug+hvSCTbhcxj
S4q6V6c4cN/f8HRPK3cF++5PAJzQKrd6ts4c+YeKPZq8KnTmJikJ8ODVnl2tUgwX
nWsInEglUzpLLBmq9A8QsxJedlubBJZi05sA3I6H949JZnp80/w68zEjd/c4zcW2
pGOtJ88CRhmzW8EV/pn7trdpknI7JdmT25iGYIY1bV8VP33RW63qa4GydEzKIhDe
jJKbwR2N9oDxF7HPEmLVOVDGUrSTNdlravYF+Zu/Y8Ij9vt//+neSRGHKr2pGNDG
Uz0dON+QAwKqBmfgMiGKdmCST13OtICLlvXXPpq0bdh3Qj89p65Szef+ntc5OMbH
kf2lXnyE6tPIduQTzCUZnULYkEqCupE121NIfwUOrPqHFUia+2p102CiIWG0PLCM
02x8Ctx/+18SnldXvsTnM1imkr+l+gIrZUPTFDCvC4kHoZZLJhgfcrpCPEqvjfQd
+2wc2nTw5qy5UZOjnc1CVHwZ31hALpv1aw1TDVWJ0Hfm16ewHb9de5wMqQ18WM6t
Low1kGp6MJklsir6MR9bymjOhgHWjuz3fySurvvQRJVTAnYs7lPFM6AljdrRT9Vq
8Y1jtG/ZYQErXi4EYsm2HRRRwpr8ruziYGLZyv55+xfV+zrNJLixYKyMChbI0fLe
PGWJJ8EVEy3Ai9UzcRDTB/hCpBVMjOjqGPD/ZYEr9RevaKxaBUGpd2XV5uahRRtJ
iYK2sFfPqfOdtadMhIaYJEX1uMFuTgo9rGSYi2V2XIABUcpFIvyvghDE3sGt6drW
tU5jX+Ivpp1YApmA4A3r4vyY/3aXc5+PDMS31gogZo0sPOrpay7LHzc4Kg/5nQZH
u5N4GLTg/o9+O70Ye2GQh3+oLwOR1qBWLEk/HTr+QgdI7Djp06sGJ9W/HoPSpCh6
/lHXSmjzhAjSDPcL1IW4TDUBmBdm/aleyt+7CdzKzrq/aWsJgnMP5cYnx9ATbYRQ
3txVvjxq4XeoewPshREVYSwJUjzpC2IoptRFNGjYPuO7ojGTn4FPYe7IK+kfEFkz
+G56xPgPb1uIOpzKRbgTY0D8hP+8yBqbYPo25KyfWKsl+8R5YzfHjduJT4ziJDBg
aPcH9gVWUhRzDqBYu28FhSWxvu2WdQ850txAGaWSNIHk35tdDtGZrHFEq6llKEsF
rOiqyRyYWsBhBl5o/uAQoht/swxu08OSYDPA5dTD9oTShUDCIj4rnO9JaecnNCd+
/uJjNtxu/54EVxQgqs9ysnzj6O3g6QVE6q1HLU4Lx2EGIhcqD1DK6QOX7Yaq/e6z
+Ij6Jysi/MvTpi4Yw+IuVpiy6w5qMiVPfO0aatIjCJTJEWstsNm8/MaaatqEO9/p
963ZaU95J/YI67MrdbHAfhLywGeOyfsdwBUW8svXmRiDlMqArVvfvXuEdHxXh3jB
j9K8V5HF+8h8kxyK/h6TCLZhKvrSIUabqU+pp03P8FK/Zl+4zgwmNuW47GovaKQg
JKigR5ByhntmkrJsOpuNPJ5W93w+/zvGSYBTskI4KvxNPyeBqDY4b3uAzTiGBplC
aezAq9sUXtKAvVOwhHl2T8wDREUpHGRhvzYuq6H/GTJ5SwIw7vYOzxLbXoRNIQ/I
BTj+415cXvAjiLe2NLIB7gq0Zk4yfTs07a6LXfCvfwtoKmXSmzThIl+xdo70yRW/
OOy1Aeg8O2eVS817X4cVNTjcp93k62B/qMJcwUezWIvN3D9MEr+hmyQhRKkZIihs
2Zy7FZ8xwEWDw8pBsJ4ayL50m1CNwfcxilvACWMX4qRoSMyThn2NHQiyTjAYzvxQ
VwS+C1e1sb7+u9qrCHJtW+6tEOsD9UgX305wLjxYTRpJa5gLM/f0sL8LS1CToWw1
xUHiINHPq0366Qq7fuT9bBxS/zhoDEWVgga4nn7VoyVi+RdPXMI1fyFSs1lWc96q
179SW+4bIrkx6DyYhx0f+cuS82MrpsF4MgGJzBXcoNU9JZbKhMwVLywpz7SWAcaf
xIEGB28bhEhNGC0VZrVGYrvzMloOm5ksCuUiRGpjOM7gMtKkVvVDIvHN2sMf5xqb
kjXRY0jiDgLuli05IxeaQ76MGQYM6wqMaQWN8xhexbV1ptyi03zjtg4YAb1vIDO/
k/tetsuVuJpOvmcmaY/nDStqsopmmN0lLdr+nAeOae+nIjamceX/xUrheptnL+pz
gDRsXseuEn1zdDLV4K1UDfVnhxHWIRv4An9hzZNMOkkui8qmpn7NUFqLfzCSRsK4
Eevp4PXIpOK/v0bMrwB+W1uwVjv8lR+GjSmeZI3sfOhbD8IW7f/bfVheP++62yKm
KOXhAEbuJb0lVr0MvJecOznYnO3PLo5dRm+BZ8Qt5yqMrcyH7AuLkubCnX3A8oqq
lqnO3Q7fEUsi8fCe3UZbnijdjAzbmcXSAJ4ievHseMoCrdbCIn+c7lvY+5YfmRRc
96S4wlyQDvs++I9QwtMZ6HpwfPdaTlNGsqP+5BiLVoWzziDoSTlc2hZxl/s9g2qE
rqt9AifrVPn8v7AEzH9VmuqBAFKhBqSd+WtLCl6hM/TZla91zVV/3fDjtliBP+hk
jjQQm8TK4soTOMwiVwHZGe8sr9cbFYqsCAb9edj+kp/pftzXRNS5621/M86wSlmq
wZoGthJ5tDYBEvSiJMctbkgk43Hx/pUiRauWqI4TTaxZ88rL20xDa/7Rbn/pRNSZ
9nu86RcYJY6S9DErnq/6xpx9pLQfEMbp3hR16514/I/R0tV9cbq1hQasXmxYB0xl
if8M7rsrg/YIymENJlQUKqSeUaF5Obs16AgPHZPXrGTZ/23WiK3Pd3kP2xBd23T7
Z+f5OVRiSPpKMjeIPfbiqsmWAicKaDaXUOrC9VRTQyXJhVXlqPN59DBPcPG8K7jc
VwVWkfv9j9BdMokEBkgTTQLFR+/F66z7NH1D4uVzMWdQ+CzWrBUbaZ6NbAXdic/a
YbnTYLDdaxdfqRjA8j0aAPnZexLwM+i1Q95oSEHW3Ua6xd0zB71SCkrcQK96Oy11
eLYlTi+JlUehmB0ihmFHRGba6T+89fEjAfDAmZKE9R1TnutxylGD4JDgXeE0/ZKT
/Tut66yWGAnhBi26gnCDZYt+EOh9aINN1/cDynSx7LaH+m1+Gq36QW/GnNDIvUM4
YJht2TCa/LLzfF/5gDPAJk7U+02Rws+8nFB8f1kTvCwh9vqpFVMqOKyRC5IROP8F
ytTB3c7ZOByAsDPyhaRJh+fwIzt9+NKap09qjDz98It/p4lHVHCcM1Xp249LCR3J
J75l5Btma1qisahdbHbN5nu1ytibyut1bHdVRv7hkR9jGhL7qCS9XAldy+cppuw4
OTdO8y5epoi+hNlBrIco/zof0xv+VkR6tGGpCJC4AxehtCximorxr85A20J0FYI2
1EqwZ2+P3hdC6OY8hZZ9vPNrER5iitxsMi3uLK//B8aJgZnk25KyDEh1Dnk7pyUj
3thpp2SjsmJrLV2T8NQ8vqRPzYJzB2O6YC0ffCLqSM7QIGip5O/xnGYxaYVHpzDY
LbUzT8qV0ap3/sRG0NRlcKc/Pdc5a5Dq9nY9Px2iCs6NkO8AulwwnwCJ5Dj4knOn
f0pmPUEFefS0vs2LdL68Y5jGQb6TXxCK2O6I8KhifVR1760e9iEm/u8ciJut4mLC
GKHVF+ll+CSoisxRHHmDmF5tzY2qQqIn21yNqx3jAsxERG0wmfRuY2i7mN/rwwwU
vwIQu2QDXw2Q5nb1dD6NOAcSKdVYJppJrq88oX9SADxQheTzqNokgLHzPcxeB5hv
mgABK/yD+5d+Lw/S1m4mRLD+0M/CI4u5Kf84CUGoe1gAt1BoVKotBcXA62G4zdtV
mZSxGnYzKmNVMEyTPhJzTRUml9iVA1ldZxEPPtc5IpeAM63Q13i4rMQeL45EOdDx
4m5EpWTAUnWKUcX49mpuqdZVntq++gryGDXL8vTlUZWeyNRIIGsfoHKkCK/h1dJ6
WPPqxbBXRs1n91y5vHIfEuN6Y8Dvl7Ho58OMkgY2ifMz4QtCmzgkKUT6I4Li2wpJ
HtSqOHIvrWJhkakLaoITGgUPkifb9I1LFDpp377NzWZtJigUuP5hVRsaIi5M77va
RqMHhtc6Ezi9L+yjhfhVgwqCJnF08H+mfcoJRVrFaVsB+e7D2Qk25VRdwjas1VK+
1X5zsfMleHVPvEy6cYxqwDVOKIz7unTwiLA04jt5o8sAc0N3cmi2NGSPe8bmvyQD
EVxJBLKc0LRZSbihsVU1cyPb3pYgbfGndnXidOPxgYqtmcDC5TpjY0APCqrYFIVK
+jNzH2Rwkq9V2W/Pe8ry3DRFYRpVNtUEX66/lCOFsbVrAiS115a5PSsVsRpKdQJt
+R97pKOY6wm1/k0BydnT7v4K4yLoctkcFqQNI3dWAAO6p2bIrNnIzmc1v5NJZI5G
9VtuOy8ANVKSfHzN+QOS8iQQfxWKAFLhHkb88Iml+JGLRIhkZk0U2+gB3SsClIUt
fDFtVZYJ34ORL1W9rbX0Qw9qhxL89V/Z8opF2uE2WWPVLI1wuIqd+R9n/rCmIWAw
xbHGBNLajwspW7TRsr+Z1MWDzaIxJ4YneIOBo6+l99Ju2NURsvkxUKtbZK6EC+6Z
PEqMuBQLK+VovU9e88YHtOOPo4JhFPp87aAdWQkWkkogws98KKoF85YGuHejWmCR
CrAM5axLyaerS2JYUENAmcwNoKGC/L2d9iEkRYcTnGnsVHFP6aOLH6ejoIGMJEM+
f9Qlkqj+Qh6/o5B9BgR2pt3Ncuq2QDCRKC0887wOhmYfOOL3/PdcBfopsbFI95E4
gCh6t/lLomZvDZ4EchxC2iGblOuyshg9vfVdrK4zx+xLSOyj8Z+JLPkhna8+5i7u
PTRyYuS5XJHpWh8gRHK1SZCdhk1oy8jeJF+Tvwae1qkjO3nWOMiqNxjkfRunwbv2
DogcMIJqUodVz2toExvIEDX+O2t6MS05LMurQPuWjRqYpsalmDhryBW9z4wA26Jg
oJcR5BryPxZrZSrRruCjmZba0Vgd2sGeVckJlYRQjHeDDVuWQ+ALM/S6q2vmXDs3
QHOYouDoSSsojSzgm/IzriEBKmF/cA/jGzdDzoACreYWDh+s1L18CvNOE11j1Nn8
4j4+fiVekyeBNc4XYAB+ObPaldPU2Sg/O/n8h/V8+CypbmIM5BgrgS5GRmvVPL7M
RFtcvWNxfx8hHNCmPhGEiJkehk0pj1j1eiEg0estvb5G8khzUN1qLMUKNL8Ha8dh
FZTqePlsQd8tkFRryjK4tXX+9+Ygi0/LPsactdkHZUD2ZI5HZrT3Lobf7Kzgx5jH
YGmJGDaIuRzzB4vGpBeNQaltO5LW3ILPO3kqcNebBJPAhINlw8ZAzzfU4qSi3A65
tb8CK8QN1mfbXqQsnGBEFHZyhfhkKWLKRnkzUM0nZ3geLpwntgaQthjVQ+Erh+Rb
eJcSErQ48DkftSBKYM1VpDdZ5QXv2usKikQ50191abXIb2S8td5dzyeABeyx1rIV
AsyQRYYSdTFLKRyjJ2rjEwgeDbGJNqec5zjHN5uRXdJ5sh3mCLNZ64kkmEtv8yjY
oJeoV0L9U2YJNV0SnLB48rdCq5AqEEh5RuS7ZGIubVWm9bHu/+ISpVtdNIxLYUxQ
LohLcxCm02wMCZ/Z3Nk/XC3VLhZenBnSFDH0I6yehloiJcIk5NErRYGlL+KI/Z3S
HXJy8WpUjunO8QPoPv155NV+eklNRXuKMi1SY9MzmG2Rcpt5ewjXTDOvwmOn7ip7
htqhOYFSKY5VK902Y3wGjTVGqD9+iJvv06XpWPwl11ebeOnDd7kgUfd1PIY1FZK/
5qGohsZSqLfaK1mvG8cDa6Mfjlg/xdv36ebWCHicBoGH7Oz0VGQAxJivqAOFNOGt
zX/SA9cVVy07i62nHVO4ESm0gnLfsq2v8GdrPg9ngT+8RpaY6oSjYVqj+AUhO1p/
TLMQ6XpFeom20iCKWAXhPbjlqOIGab4BtCWYocVM5Vi9znMDSUgDaN8jdrWu4l13
Y09nVHqV5sBX9bi69sCyivujvxvaC5w7MadPBUQfOBYQnByZ1xM6B/AnDQJMMmHl
Nkprbuu5sgNuTY9z5HCFm6rIa+hyhjL40iRAEyxKsQuvtRWFy3rcHhP2S4FTHEdW
9KUREmVhFQTtALx2j1SzCOybC47+L+uJEAzkeWjwqiHeGURgJqCLLadKuocwxngN
Jj5+7WCGBeLeuUDcDBeuV6w2vaqCCAvGDIjAG/49KhDXLL5iJ6TTDjU2QCfByp2X
yPVZB6w3Mr6Tc5E8+gXxzBe16oX4o2kPZ1i/xVqUV1IXOkMzOgZpILu30nIx8F/5
jGq+pHe/72jr5sJHv6/OSymsYBjB4S2DDod0aTbBlsk6I6BQqtmvdOLx/1BLccuM
SlOL1ic5zZl6jhE6MXsIqOOQ1EqI13y7NozlHJE4oywtAlXfaVwOcHPOa2flDAEp
Swv37QsWU0yj0+JJqqA95oPDFCu/t95Urv+HtQs6BCjLCRijATDEjOiBfTC/7EG/
9wDSMJmsQqoU7uf6X9NlI7wLrqpP5pW2IBTKuL5Jb7F1fi1VAh8bVFtPz4wuftU1
5odG9KmC9my/epR536bfUbFoVterPpysMIYOxPMt8C4QwvxnQpzl+BI5mapnX2XD
1NAJPkNhsK5cjn3Yq3XRoXQl25PbpUqLeKPpZV9eRofRE8NsZGukdxgU6Xp1DaPH
5Z4t4T53GBrk11EIFb1Z/JnKR2WmceytusbHh0aaxODs929d0nL9cWrkQz0Cjb6w
pvjv1tMm3e/ncWQtaxF/H4m1rBv5hHqX4cb1wZ3T8dDa/ukep1Kvp9Y8Z5r96WUa
U6rJ0/2/9dNzy0Mcbccs+i/N+9WXC2eARZWm0CbgLUTguXOMMKQGoT2SqTuizH7c
2ukfM6Zq6u43XMvcSLX9WyBjf8m1tT/YqfW+Mk8p1gqrUV7j/v18SLr6T1psFkIQ
KSLEPzU8krp6AXXy8BfApk7f0GsGFL/W+A/ZmWviu5mh5Rmmb0V9oOuSZz+k6GDw
6zrTdUiztqVb30uRU2lJHy84Blu3DRAVbQGs/xbwVy0XL4dhKBGDbHNJMVi+hG/V
si+/PSxXftu0PHM/mqoxbX7kzBMwezxQ0BDb2LkxfHK4OfD+lgmkqjV9569PJ620
BhAJ3+5PyaggLo46P24kTchnnvQYKuLk9LZ5NVgi2p7uUX7D8vfBgZWuoaJ7UsDI
CME6i+Gc4pPnWRfTfp+ptSxjm0PHyYlPLIwof2New4wIoIeHSxLgL1jhQSaKawAN
Hw2r9PKW+qGkqC5hVCMAEXpyoikHjt6+SDe9WS9kABVoOXTZ/HEjit8w0VsZyU+2
NjQpeBg3QfBRjAORGG0sU7XFWRhPH2DAoOAQzcdMiVoyX9iGgom06ia2yzfmL1BF
QxXe8yhvVXGBv7egLlHYjAUSHyity0KB1xhiu+Lxfu2rJVcJPjbY8YxnAV+2qU5z
qMTHuQr6WJXZZxWVLTmM9woWTfTuDqfd6yBAxfRMxSSV4gzLBV+d8LDMYKFMDzRm
K0NOE/ymHMNcyir5BIIxfHY8Uz3rSHCRx7Xrj9yAueDEfrDc7PkycLq5/F/LePeX
LHu/+hP78UihSNyl81IUYJAezIizwv+oWk30RmOWJp8URKWzuFIkhJlJqzGUjyEt
CE2ZumZHKHoqUnGTFA2tgYrJJ+Mhjo6DboG3lkXUvqk/hNAwV36qPgyDtrjQ4DhN
DNmfJRgSL4KBJUNO9DuXvMQFr2fyvd3Xft7Duy5iAN2eI6ZYMu7I/tJ/o1jXFmli
wEiz0+JO931NN6z4+T9fbpTgFpJwVlr8HG46XsOjA3BHFs5YvG2fRjHOudUdQ4U+
9MX5HIUoUey9LEIyN3Ill0lnqHV0gsRStuNl5DGC8nNVO/B/KCR86+GpdwfIpiOV
NWQVnA0fl3S9gLfg89XloiclfkJNPybCf1ZdVlfeb6SXxX7YGdQ2n3mh0745x9Px
VVDv4rQM0nrwcpurG7wV4+X9U3Cq8US7LbMhc5wIQLyqtFeU7M7ronp2kdotbcmW
r0C/TRBfg84A2wt+UK8BozMjT5oOyLeaZgUCHa/TJyXNE8FMbHDlY2hnxJHzcTma
X+gR+gM1yK5hOeihLjo0JdKHF0AnGjLpLlyCsC+ZUl4YLaX3Mz4u1m1BnOHCqMK3
K1EJCrLm6Px4jj6SBzfNv30BBmFJtZtt71wspGZJO3MbpMidC4iWtbmzA4JNy39L
PAT6T27Dfl4xncdpL6nEOv6dmytjJGc8mhZUSko8G/x2U/aNl5oAqCD8ZXyAoVsU
QRCtWLZDqumbqYMSHzy/LcQsbEGXCrmm6+hnwbpe3Q+95z0yweKz7LRRVlmtwqYl
XCvV+2xBl/ndZ9hrFt5j7QW8XybhRm1gmKiY/jdsxHRGlCJT73nwAde9hksmcbvC
QW77D1zh545QRMib7MPZ+U5rnPrQv0ZxHa0K5iO+jImnMxxOV7vnchuGSaCNP9bE
YHi8pFR7YLrFmqtmFMuLNMrK38uNyF3bzruu6ZP14HZgnywnuht1VyCAoUh5tDf2
mlRNwQ5J5Q6lRr/cv1TghUZ1pmU91nlRVonuYcr8MljJjyDdQVktza9s2fPef/up
xjCJ8FPU+rmOBYXh66yqV5eNQCS1gHd/rUHl4kaqfMb8bWDX50RRiqKbiSwE9w6n
9fJ2Sr687ySzgbU+tacMnq4eVJ9fI7BBbdsoVxdEMp6eERIga4CzI63wfzMmzSI+
vUQU0FBb2QTY7/+FYcmc6f3NOMZuPZYw8keAm8b8QMa8WKp9dxC/DCPsX8El1rwl
I1tuW+I6olCGigpoNGM+LtC5RSMmRfyrqhAHNv2u9MmHHeAJmLMtT23pKGBP9K6V
eSiII0YVg4DbrRatz5V2ji5mLC6ZL2idn2xJBCDIR7bitkO0zXZsOGRHAbiF29Q6
29mO8JxPQb8KAJ/knnOCiEfuWxzsIPZEgQB6aUqPJPCa80G7TIrNjM556K/peKQf
u7FZEL/ZpV7dufUTkN0h1cRKjoLR4SgWmw3NSrUmEhITIsegE1tnT6NgW7Kahent
BNNkQqyF+QxxEGENqBCLdibp2e1JzWT08G9b1DltSNsjKtOo+/5GcU20F3jvM8xi
aXVq0gFPYHkSrICWJi82J+Iq5Fe7lx7qqzMq503DWFE365Rv4hkcOnP5Mg6gnIwc
QoKXKlkV3lpNXPvAvTnyZ9ZtSMJpRHuJh9bFtEK1VqJ86o8K7SppyLE4fKu1NliQ
Vc1mc1sVDN8ckrc4iN5v753IUk5fvx5/ElQJmvZ3U9yIxwYCxJsod2Ld3p7PvKeh
/+yEGVAdkFcK49EBF1jhHiMDgHk8+08ckhdbBaRdW43f4USidzyfU49jO9LkkfBC
ieqamLdZn3MWjb6yngeFQ/V85Uj4EvmX0aUCk1ABrVB+3U1LocikUnzZuUZh/pVC
g1yIAwX3lnD4BeJ91kK/KNCe6ncGN1FtalFpbJ6xZBbJGwMzf4xBlXrE9713kRdP
03pXxlY2LBXEjjUTMIwv2Ve1gsQC3K2wZM+5rbEp5GuZ+J+OR55w0ULsEhAJZotx
RXXSx+c/Scc8kNq80D9IY5Y9tCp9/obflBrbfJ22U1Z4BWCr4OYgXEkTlBXxXjT9
KucJbCZ13t+eVs9yx6LRz3+Xil4Az1O0Ss1aoFd+2m8WNClrjVMCjcmudtLKO/QB
cCMsLR8DHP17NehUSsC7jt3giqLVzGJ3gF4t27+PvPRFV5v4LlBJr/mmqI7or/RZ
ATfwna3GYg1dn+uNvCz/6u2W36liToApVEmhZY+S0tmCkYMjWWXjYT1zgN4IA4UN
d53b9g3L97aORVnL5YFQEfC1OX4xh53yv4FHVn/JUv+JyrIqMFnCcvMWaTNbLgqT
hU2Wmenx9lzg0Xmpd+gwFAaBlHirmzUQC8biVPSLd+TUOzgjo66b5MQn/jv+/LDu
J1Vx9ZgR0P1K0ulT8IRX6Cmncvnux7lHlqyFaky1vjU580r3OG1PhFutpyw5JkQa
tmou8OWd1AoXfJswWoz4mMdisEmPqIAu8ZnmWRi7INYPB0128C7YF0uATXpp6jIk
g60bRlZgTlVETRf9tDZn9R/75IwLSX/kz9eHjumpPCnEEMZbk/MLKXmrmV3seqrH
5HswkFjLXczZuBHWz7gtl/HtPh7SGhA+Gg7AJQNNvFw8aOYZmAhDI9/DgkB5oEVU
WV6xd8bka88EQQfmd/pB2aMnnERrMCXrGS8OILuXs2n9lHpaB5ZoXLuJ6Gm2m5Dy
H0huiNJRoZzvSBgPhBhJ56ZaiDf3UqV2gYRcH4+3onKURxCWK5Xxy5JID59NZ4bq
s/2PvTinPpIRzx5taJBEeh+4VE26Y9y+oRDcQ7kPyDBCC0q10TEV8PANjpdPJvrR
MGIIer3+0ryp6z08lFotccFIiY2sKoxJJP7Iajsm3bnqOIuMP6JpHx0qs7bLjyN5
WMFwbxl1PpZ+aTq0o5+n18ENN9mlNQFjuqDBdwVPRlKHplS5VV6mhGgOm/y/nHMp
doFvqW+02Y0lmfQFN44FGLFduZFQk7Qwr59QBtqtUodX4Cbkw4N9X2YXDKwodeFr
PePOkQ3pWmMfNbE5Dxqs7LmBtXxPe8JCoQz0kN2PuMO5EA21HWK2T6g/8SnyYo/M
upwQqeHXG87yEnL9/HzlyKCRkdTlkfatHaPpkCLCLbj9AjLsonTpJ2E1VaTl2lwd
fTkAUn9YHF7LdHn4X9vbg3XmrFv/ZlOaz30RCQSyRmactPpBb+a4HyNQsFZc2qrc
IIEVwAKcP2xjcAfff+QVy7zrh08m/etbbnaz5TOz9tl9Nx5nSfT6lh9pBKDLz7b/
SM/QxAai1hPOh4u2Ylr4sCxCcsgLe1HWT7zlp01RzM2+2Jw3GyXsrJmID6yXALga
NICLUcCZqINEX9cttjAQW94D7WSyjBWQwJz2WjZXfBUgBpxHj2ppVlJDsRWZ16GG
TM7+LpZFAd8q1GSFeQ6syhsaeBkgXHsqiJiYaFpg9JmtFu3H0dHuX2oibCZSV3Zt
pdLBng1W9nReJh4G2rtMrBmc+cZG8cOkE1tf9b1w5XyNnNK/96OKOzorqIhdhHE/
QsubiQ6EURjs9X98RFRSDlLxe/2qtM1wKlPR9BWa/joM/Eb0Sz7gg9pU4NlRi/Hg
lWvNtTBjJf4MSy17AIcTh4f3cB2nATYBYL8K7rdSTso5d1TSlsxDMasltHBgkOyw
EUof7L7b7J9FrOfNHLWr/xY+hdce+SJHO6bmNw1WvVkI3Z/UDQpfF2UHOTogGPpP
2ivfYPagO566uA4EZTopxgANDGP/bRltSstBzVyWaXU1A4n7rbKhvuzJzL6xmsgN
u9yaPuYHeTckIFRLs5RzQ4hIeF7drJ2t/ZaHJKVdgUvs2QuxBMHfE8SmcUwsnZ8v
jN1mmYivPWHjU/5Qd0IqXUSe0s2cek+ngMdX7MVr/ebZ40ixCojCNNy7eizQ2kg9
83oRQ6HSgMkgFHfTKdnZobXPFiEUOn1H6ju2o+WQA4a+MBYEqQBFREP2zc/MIOco
3EwSgHZeIcdNWqS9LRqWzlJsx/wsbZHq6rJYzroK6+dL84yHy5TBJ6AiIu2NQ9Kq
4Mcqk/ipSPlaE2/jWOjJpA6VYcmOXK+a/DLwb8UNC2nwT5MR6cPitW3MelFcjmak
QxNh4frjJhQctgOU4asGpDDc0gxZIEykCcClXUjKQxDYqivEc5/BMy0WQ4h164J7
FZT+kNe9h40FW1oMb4fX197I8JyguAwVTWEoZxz//IZ9DyugWIOjsraonKSzCzNF
3TgRCtVbeGP1NXm/KmqwESrZJMzP1pcJESfjWzAv5/bERXgMabMvhAQUjM+fHrKq
NU2yxvX64QNhigLiy+km42Q9OO7cbmWCma/hkONN79p/Lqtm3mmgzWk0JLaOTI1i
M4QHejHivVuWc3Hh83dE8JKE6sTHEjaJLkmkNkuteadgnFS5cldMP/c886nUHzLA
Fxhsw0BrZULFxpL4qz/GtA4nsJ1tgDrzlJS/7fWu5kwOoindVI6dVY9VFQ39h9K8
7g6dv4tT8GXEHsDqJghOgNLj7HHbnfKPUGIqw3NmZmRrwK69MZ9oBDxZxey2XE2+
aBmEgw+hDJUvv235L3WnM5xClB51Tb3d9u8RrB3843o2LrXblCkbn+5PLX/xegv9
snrgJbDUvZBeiXvJmBdUp85u4W93aA5ZnzA2yLMTnHTkQAgmq5V8MxGl0ihj+bnT
5FrsjZDJpcKK6hfnURwezPnqvoR0JFhNge+7mb57+osvohh0Z/R9m7YlTYFTzhiB
bQ8lMYf26MWl2pCdfH7I7T0+sEsxIlHF5Kh1y39iwmdFe5TsFmzn00Hqxluryfsg
wrmm6Y4Zcyjo1crRKRPW9JhVdvmq9vb6QqKp6LhaOCGOG3Mbrnbfi6N09ERKAYFE
H2Z/KH2sK9tYBgzrHV3kXhiOtkN06M5FaHqJ5Fr861b67BZeH1vi12+2+c45u7Eh
gKi5R0JSuFTQQr4tJbJe9lOSB6OAqlwqojCT2nsOEibi/pcl7vEJO2Swv78tr2I5
rwE1IuuB/OxSBQL5YIGeyObKGjkME2O5+sBDIzia+l1C4+xtsBI/JGduAhSXNynx
1Oer5wuBgLFk6K0TRh6k/GbKaibFe49IeBGgp5FYTNUaNiEi+2giMP3mCWsGhNn0
5dU8PwtC8VAcQygmboQMWnRFMEu+kF1XWpWfCSqsDvF9iaAWcWkxJKkiXx39h6+7
NwKgZJWTOnn3ZUcIEjg6NsTA5u7J9jUJkc5hpLm2x2V2b4/dVR+clZitZ2Kf2ylt
9cpqL509zGki9xQT5H8aTEe3xdoOfTvG96F9a6upHbF8BvPicFXdvjosfsKJ5Irp
otgiNbpjYVnacnI9MubruO3PVtry3vqagnZMdtJR8HAUE1fVDatqjspH8AXFoVbc
TANn9po2Zg0H+Pj4c99PQ3WrAXP47zm8Ip2aopB7nu5Mxpd+iMgw3QbkAKkO3GJm
8l7PI5a8C3OM3JO219NC686e0bUyawmmcqWyLANtLBhes77vB5lHxpa9beUhpr3l
8TCeTXzjZfstecBKjw2pO6yAtguoqA8s/c+F1doHxRrMvvL5Bm8yHzvM2b+29Tfl
hALydFUsmo5+tbNWwovNyUhIEDGEQGy6Gvb8jgNLvhWVS/fSykDUQBvMLDh9k6Ie
B2ycu+YbwkMRcosRhHQkUO0w5DHC9wWvs5bt10J2+vkOm/ub7TFds/yx0Cy7AjYt
OIO9uUDPva20zmhsNd8DvalD09pP6A15mvDePLHqRBUd8rZlLZJoLtlRF5WNoDyL
ab2eteMvXhe6kkYgRPr0syoIpr0/LlZdRExI94xgfwTBXgAPx1L/z5wWEsd8B9G2
EZHug4Eb3qDKXmBjctnHfi/Sg7IUqG9SResUrNb7sKCcU20dZ7rs1WLQLDqQDu3a
Yzo4Ii9bV7PmNAatqBHmDfzJIUVjOu7Ymz85ihypIaJwUm7VDRVgELbxyCHebe6k
L0BViJbnWYc7+Vhg5/Mhg4f6kKoIB0hivPsKAzZrTCQYrgDtCW8aaRc0Tl3xICt0
UfGTQhUU7aDNOVERB+3rkPq74wcMxcPipKix8dD+OWo6Ndf/Yeuls4TbGDk3C0Kx
qZsrsV32ZKJfilDRkeTpPD0n/LBTRXINxsgo8DlmqJT71Yz4Qku54sLxRwdtiUGY
VNKXUxK3RWVAMmbdAQttMwRFVKHgDOnoUQouZS6Xl8d7lnkrmor9i6ni/2+t75y6
ATxvJRf0Hho5x7AZAWB4GeiajwsuYwNwDZnmht1VJAop+fM2kvifeFiHdRr3/qcK
Q57wF66C45AtsnQ3JfbW9XlSsj8vbqYwIn3Wpqg18pAQxX7juo1EAwj+MbrI+qzp
Pf6kzh+iTc5lWVTNTX8H2ZlrRyNVchSIqrhXYbSZSn7rpAyTryMVGZy26/EBLQKQ
nqMwou68bOcweHyzybTJEVLXDzxZn9npvcxvnUU8ZXveXyuIVudB33XP2Yw9fglb
nqUCEvHq+S5KAdSTopjy3S0l/Xxdxd2l0XQmiTUsSaU/8HO8q7ymV1Ei66ynJM9Z
AVjiHl0nfAn8v2igWl8iGeN4FLKLpSoYFbfL/OQFlhAdQSrqaSRBXlMsaLjcm9Xv
GKWJoHJEuqSh8fjxPhpSHT2RQJMzN7I/33Fl+PKghAjw5henPe2f/RCysy47gdp8
R3HfawfbjU7wd/CVh2sh9erFQB2TgYyueHgqcipYNTBCaBdtgH9T+b3TOOzt5KXM
Y3kkRZUgkRCfDcasuagKSMWvMytZ8bnWZCDc1Hev1NC1nP62E6PDXp3VAspA/3Ih
WWr55N1is70lkb5T0qO3JBuNXRNBUcIiiySoY55vImUPKf3fM3nkxxXtyqCcQ3zB
gHjdpWkyPQxUUdF/n+gykqoFs1HIt+a9V5EKbC1nh89wQaMC47sPxDZyDrrSDSy3
bdnSOb2LJHM7OZyZ0vV0wKl4h34skWfc2gPJBLC0qvBDbu58vPbVqo6zfE8IVdtB
kwWM18UgZr0igDivAiKrSqDunhKjOXuzXgmJKo6lB979xHhW9GfwPtwRpEvnmhK6
66jR9KbmBCG8Xd/acLU9U39jDaptBswrPcgGAy0xVBw9Ij8GjgEIcPclkbkUkhcO
JVXgMbk8AWFLaZib0K3XrSj7dkui2BKVbGEAjIvARPu5Oy5/MQglKpftO7U643eU
f2pe7gsf3rK/RY7JpuG5OxxCrRpKH0bI2Y7ZJXxEEKx4y9rQMeTcpZS3gzz7zLX+
MAv93GvBVNPaMmmO/WdZs5M0UdDDO6qYyUcPl5bClr/F6Kb/7eN9jc/tmX3hIaiU
ebHiPJbj/IsZksVYikbJ8hw5Yp/CGW2PeidRDSnmWZ1Qqs9HIGQf1RNn0KNiitCu
6S0LTZvFr7XesnSIa2vNzYL7bvediig7SrwUBz7T6O7sSW764xpgq6+zpUYg2teu
bt0yBo3P8zKGi38ZnIVqKk0dYM7k1cfZoUNH/fEAVHoRhEXP/PJqryHArmVlNnIT
rB3ryFVgTYIDgj+P9l5efEm1XY3MX4NiEXO6F52cy0jFRrrUo6CGA4zVFbOsCu8S
8qfAEp0N1zTwzHfflOut9u8g6hLXvkIHlaIed0q6FhPsVTwpEJwjqv9r4LFUJcFJ
da9zLrzsUJEOyfRorFxWAdC+A1pVoNV5ZZ1OjA2QaNRNLNNVUEuYf8U1wj8YbVkN
mQvdAknBu1w79PKHgtIfzJnGr0Kc/aa1uCPASTSbwfyIhX5yBGBWeizXdHzLduvl
VOcuqlKOF2uzPefx9DRxM9IMGY2RX2IrGsJIEgqhPNqpQkRiGOOBrrGSiw9/GftU
J7kxyeBCwAQ5sJu5TJOF2o1ws9ro5XzDC7Oj3XrWw+H3tcJjECVGryc9iiCjyORb
QzYV9pbi3wlic7LDvirvc4CsBDKt/FHajah77RBn2MzIYf40qO/mU7gibKZb+sYX
c5VipFKHgHb60HLwbvqvSxAdlUTzpIKaQ4QSbp5SXyGZ4iJNGWuuWCFLdkxHyfbt
TquBrRJOPIZJl5PLoCpgkgpqV5nMZicq9AiegDG56JhOgBtygy2v3icBhor+c6Rh
lVlrqjYQfgSP6amWf58PhtmwU1pYyk58t5ftShL9Ig18HgSHCYmGLfKsyGB8mkdu
W+YWp+w3Kyv5xhQ6+K+tTBklkBqLtTg1fv9Y2zmzKRQcFue3y7r2DWMs7vvTgOmb
bemtlVm1D1GdYXV8FbfJUDlZBoNNv2Uwu92hiKZQSexlT5xnvyDA+82b4MTVdB3v
DGhcWv91x8KKRTCXPZPOb2cP5yF7ldSfvWvOtehLCXI8hZvY9+NCLJ6sd4DkF4h7
66juCv8HHvqkVgawAlbOrtOd/eTd6HJPBZSHjZLBX81URfTkxvLcHfNXPNYl4nD1
lhgGIBl82JRDXetISO6MZp6uNVuzI5lwtYhHNadptH7MLHvg+urC4Z8P3fTC7fRw
EJ3karNeHN9UK8gx54wivEed5a6pM7o5BQqVkpkPIVqZmxAO8VkfX0BudBr4fkA5
AUbDu5XIlSIwQPFKHbzQiKxrI2a+5m8zj8aVPysEZIjdBWqJ5tPl5OwLAMmUTkNX
MVdyQH4HifPxmZHb3rXgggzv/VpN+4MWQ3RSVjzf0O0txTaC8Db3e7SGJG7Ds9+6
OTX54qApT1mcXUVYv5tcxHWr6x0xNIs1enc0c2PjNAjalOamcDZ/EyVvgtq05Qtn
rmfyVOOFyUjvaUn3w0IDHP1fI/Fs6pp6irdhfUfegasNNlHp/QGmEeQKUu3eWoX1
jRUQsV/FoPb1/HmD3FcGPZ07GfMXpctoSK6aaWU9UypUKPYuwc7Z5UKVFugIYOoS
OQDqnqtX6R+7lf4ibaXwKwNRUHCQoaOxLzY5fqnjry86hrI8X8khXQHynft7nnbh
RisAKS+qEWa/YsApJmMxlZI7YOs1bg7APyVAjlwuJC+BaVVbCNnzcjyYWxpZbgsk
UbaB557iaZCHlwlwlOTGT8yh0mEinrC7EZPtPONhTU6R0D/d4BlnUWn5WdvEdSgW
7X8GnOxQ+fa7N//JD7hUQ3CuV5rZs+GrXEJLK5HNcBSxK9VsjX3XyvU3euA8GGO5
FqFrOwBcxdCEd8B6LT/0lIa9LgGcF4yZq0ZwZAwkDveNe6OGwazHfcF7Kvtkcx5e
ov8Uppf8zgzYr4JyUDyx1o9U0hvObcqVs9hKcFLzqtPxiVNVVGMXCR3Xuo2iOJpc
o6zqRaR4d3IqBp/glnk3ukb7+4RxZl5xpEQn/Y5b1Wv6rw3PLIIuOXA1gxKOuNg7
XJHHEyHxr9A9KP7HSIyx0E+fHJMHG6f6uvlP/cxTSiOY7PKlk4R3ICIo+SeDGayS
zuMEbzGGJIKcIFnh0PsVMaZit0y0MpWfdhpDjDP1x17JzQEigM6Rla5M1Ny47vdn
NKqa/ZYLIkdwSKKEwu+qTLQmp+cmRarzNOa0XGt88QnmpD5DdVHDhKUc54egahO8
1uPLhxWkYgxYYt9JHNqXysi3FS1M40up+XHmnGubg8TQj2T/UmeKJYZo31ckQp5Q
V3EczpjDZXoBEHXzzBxDQV9O7IOKTmLzUWjbNEe1a0LDvCD5XtWAUfOZ84TiEkn0
mU+F477okwh57gQR+nc6+8pt68cs5poqt3rJP+o9wFSF1WNiXK/Xc05LAaM6ADc8
6I/ET0v3pWJH/f7V32AhRF3O6vI0BLjeIgxIWgYFNYW3HYvtFo1pQRPnUPmf+uYz
XwRgIF9h4+jIJ4QXTbqY0l5pRC3V6RWQuhPfRbTbV4YOaxLCaO/SctZGN/9dz+zk
x/49GRLuCVQoGN9M4O4XnY+TKAl/2/2geqdHPX4jLzuhWJTmkENUoO3t19NZ8+BW
/G2NLf4dytp0deyz9Erv/PIpnrwfpHV3mNcb7nDpSZMF6Cb0FrJ9RzcZi5jK9KLR
oR1ymuzFlsvqBcb1RcV5GFA3fMmr3LzCLTiC0PU6JDyyq/gTVmrzNGgqLiqa2bLb
b4BCnEcDJrojuqvI+a+u/4Iycgx4bLafCup2WCVgUqIKVynwXTw32vllHZUSwH7V
DjD4OqaHzSe7Q4H0+ZtdpHspl7rKhKKSDRcjxHem5Kjdi9oTUymLZJ585fE9bHkn
9HINWoUctI7szIDqn9Q69D7qzOQEo5p6eatRQEQyege36AP1uMIWRvemT+SyG3dg
KyAXCckjrm20MVfoLFV4tV8AFryIaOLRPd/P4T2VAvGB6b0WSGoP0dcB74vKh/au
ZzRo4Z2VeeyFjnrm4OzMf3IOlIztNg9YqaynIH/eHxqEPTjwoxcDFkWGRNG8ALLe
NR6QIhD1iOZaNveIVRKOLB4UaCeA8DS+iW7OzPDU62snEoYpmsm/gX8QOYnIMYLr
3ruQU6IvdJKSaOiAfipmtoyvO1xqxTCECQg09WmZ7BvN77jAJLRD5DBH9fUxtOAu
kHhdwTkf6/DkzazZMjfNavYZxcdemOEMs6moqDUXz+ftIIHN0IQRQJbHYV6sHfuu
EB6OHH34Zef4sSn7yS6YY2r5Xe9Gw4e7X6H06jg1mbP5dxi0dYKrTLZLrdTvh+HH
Me2id8hmGwkNYAl4IrZgyP0WeEMBkgGi0PLi8/bkkPF5Uspqq8eKU3QN60CtPoM3
NiAIppNYOUuP3tjtnV1zTlRSJ52Is162xtl9MflmwOw9OudWSk341QJJL72SnMYC
oc2T4Vw8shUE7XcXlv4Cysk48T03QxmA2gwjteb37Slf6IbcdiM2Sla5SAPmwi0c
6IJbmBkBW49A+Uz/s55SRRB1r7nXr7NVCUgkPL61Wwz0oP3cmV9b1jmnwwraneMy
Iy6dwbNKMT0Q7lnhdmHe30sI0pIBVty6yBxHCAdm8kMqYNNTzgt7beNUZ+FLoCX/
3NZFxjQJArK20n3SnvUES1z6/FDgrJ9wm005ORb7wIGkQTZY4kDxIMqf9Mz8FnBd
JLH8EwjYlu/BaYh1Meq8arMQPfOQZdG4WMYj3Bx8I9h8h6T1/35liuP+VwxYJ8B0
dCeSljfPNmlBhbYIxNBXXrftbdl7uogsr8e8XhcX2JWSWoxyD+YJ2VACd0ossh2T
dMwth5QLk4Y+ZrUauqbO2gnQYkG4da0iupvZ7uACa6/m48stl8GIN+Bs9AYf1bf3
zEQZe1PzOMlOXlmRgaPkjoIr+NKvXBeEZ849sckkS4gJEoDMRIlrqg7axq/PfFT7
mKAw1gCbaiEj3hvJHv5Jpq4HdEND5/G9k3Xo7EMYEZbHg6EByInNm92j1aeYGe3v
UR1wtYcosnoupCOobvv5GZpD6/VbZ8go4d0gmzzf/Fk3mY/qssgNujPeUMWqLiys
ZTLalhGcjEKop2Rs8qEVpxIgP+RmFq+33P/4DootOyyvlZa/HnOm8TjUFb2fzqhh
KxI7UhKqO7EUGknV9C/6ZkfvxiQOy2qATnJBYTH37WPnrEAshPo/nqpa2XWkAM1F
tDjN3S6F5RXrA7cPN98EcvRu1sc73vpxs78ZODTzpQqHKEBIyS2CUwDOgFuvVckr
1+fr4xeYx8vIOyEqUCVZgPtej6a9mwh6EGXK0ZVZ1jqkP8AgyBZQCmSIGbq58Wim
iSB24KG6WiJS1acV0b9R1LMBiN0tZ3dyIqgJuI9OFA7O0hcnAXtXrIywx2hn0m4q
IFRa/tIMe7jn0HT+/rA5hZu8/1BbLRmiZ6Y+J+XQZ8q4D+IYINaMnD3nkeQ65b1z
WXZmI+HPZK+4A9l136LUwb8jSQIIoBdDI+oTjNf0873Lzw78GxPoEZN8MaU1Vzop
V0U+honISVCQmK8hE0K701PzaOCQwTRSHkOz8FNz0pJAziEPEQs2oFM/A4ZZ8R54
/bWamgL+PtQWGFnS9RprFKhPUWJTChExEiBBXDost9/a2uRuxAYlIy/zwmLvdBph
7QOlqtK/CTMkmoj7boUYnI1Gh9uBHA2ZNG1K6ap+VGRiIFCtAZ+VADqBvvQJgsB4
Ic38pIpcvKm19ErnDD0sWF5dZBgDUgCkZEsAe1G8Bze2IPXpvBrW7mNFoch1ss2/
fvhPrZjBrurMf4CVJ8xBX2Eg01dQ1QiT4Ii2lc9MDyluJDi+loclzz5Y4kZp5i5F
WYn4NMqUzrTPRrSSTlHtI7nTpm35XMXrDhPzW5oN5jAtNV7baYMHm7qBh/x8j/nV
lv6oLJx8J7xH+Yfe+/nXP7t+Yg20Lu0UkXlXojUAGzjKE1eBUxP6c9PYeHSQQVLx
PNXDHZKiZmr7yIe9drC+gaUs5v5GDTmPrbtFTobVanyVvf8dFFLgwKZkjL1/sFp+
usWqhRgB4udilSWQFOap0cwxTZlJ/MgjuUxSgRIxmin0vorELqFPt9wHfbHyJcY1
45u7HDv/dguUgn/ZF7gXbuQxJW6kTwujYTcvXq1mjmYe1Kml9P6Cx/dll0sd5x5u
vE3WX/ACq3a2Zk6ICbDShDNWnWH+geUFujdRs0PFfneThMWAoLE2jX2jNcEnBorm
X909MPlPcChpnCX6qPqtIvJWCYOrOTANRCgVNi4TIrwmLaNwQ7cZVhZnQNSuW3Vq
4WW5zTOLqIlQwG1tpLjXrAXdn70iXdEpYCdpIoFyo8D/dBtEDtDGlHxZlNGSHavf
Ra8y/kNi/hhXmsA6aUuMnmKzhOCZiJ9o9fxw9Pf3/YaDBDAxReHcCqk/MgUJfk57
jdHq5vHYdJYNDLU+5KBFd6qNg5YVpQq8Sv6S4SqFuDH0lW5HBWaY+nYJZV2IyXfh
eTcfoEDyvPNIvEop7RvbODEdfKHfWy5O8BmBnqZBBMTooo5dTx8UjRTvSf3EGs2a
EU5qLeQYuXIE4YLWkqEbO6Nhd1QsC6VCEq7eK7i9dJFE3XvIBL+YYd29btkMDszf
Z1K7m58jkZBSSHjsMqj2u8UtE0i/Hh8gSRL4juDL4OCw/zNv01SlSFTMlGIEdt++
2lYmQP6W/IU5yuLVPeAznCJErCxlvAhYFgcICYCORw4+YnVAuHpQovPZlLEc+eH9
ayMgSA7vLrdRN/1Y428u3mQDmfL+uSXnN4/QOM/Q69Vimc6J4tZBbHpIHZzJd0Ft
JXsOWF7agQ2eDbq9qPefVYpoZwbBDov5Db/uFiNcUBDRIpKfT1mkeYBt7uMs4XtF
HGJvf0fXp4n5Jlq5qS0MSZdEsZHCB7zH3I9reAhJubV54p4YRvXhnuM20pZ/eVkb
uN3/5GZ+wUAEO6PpBkd8MF6de7QtR65D9Asumcl6pKkqzRDhX0bZfBHGixjbOUj5
Mg7LluzkgBitktjXODXUomELSiNAIkxYB5C9nL86xqIxwHGcoxxzwn8dc8PvDHNF
bOWhyl8M0CpUjKjFTWityj6FNn5QBb+DTmNOTvLfW/r1PvSn+jhOmpRtjiPVLAb8
zmHDDgDYMs6t1hCkZ0E2ngAUSGvkbi3mp7k6w68WKJGflvwXiq5fC8NOidpHXsmi
FksdPMQif65/dEUfylObkiCyE0WuFe0NMIs/yxwFpbbHX5C3K+jS8fTLaR2XGF2E
Wz26irvuGjTJUEIbLrDeA/che+y5MtF/ap9KbHZ4XZSkHgkGHl+oWL3ABNndLM89
mekOHfbmFQ8nuOAYOxoc8Ut//6uyAv8R/VQoYCw6qLq2b3fO+DFHJPMXdehAgkVb
nxHr6dIPZzVuVddgAoNSl0D9MpYjp7a6J+tDk+FoS0HTil+qY7McC6y2+kyqtUrO
8NzCx0TS90EzbkHdXPrstnLCZejZZqj1R7vnWhf3KkIaqHpIHG1Jb1A4lJsHp0fm
1pHzEvcARAOXW0xqdXE2+ykJcA28w8djHo4QLHRSQh/3KkMgXYlSVUyXWlBQN5ba
6JfNaZmOsyyZ2btHCg0tTOxX9YSi+sK2JJkD6//WxigEXvxk2Fvu5fDKxl9/HowR
XR+uFNKxHREohwq4yDK9PM4JtsS46npU58wIZdZE/BwwYvnV9moe589/CyIgVvxh
pyQBs3DYugBSmN+S0F4RQqfFPdbhZSx6X4/S7x5kR7oINr24nokDODbWIxJBf7Rk
SomBn3EHIyTkLR1DQ38GXDpp8G5gYIpL6EUrYHcQMVSoWiBfchM7tu0zkTeFgEuA
WGrhySseZ9U9Q8GAb2vrUwqwMdoMyYFcD2xa3HYShDGuxuBdlDAuZeQs6Sk+v6SW
Ptyqmla63hySBAqOJ80RJsl/sY5StWHWYLlUe7OBbwEJI5F4bzzWoDssI+3JNFVo
KBwZGQsjJj8obJX1jECOBU1ULx+nvx0eq6KKFjk5Kxp9ponLBSkP63VRoa/QR6az
QdrRig0yUcoDINr9h52V2rCCq6SX6X0Y40EAd/qtlgwVNTscoWYTdFqWd6ywfy+c
tQRee0Y53bmRL9XP58AFR0dCx40Fdfih8TbC9B2/fU3MtG97YjZIbGk12IQNNsA5
Q6fYvncfAL1yswlF3O7lSnrh3lHNmMohcbTIaORv4dg+FBqu+xzO6xwrNqw8LmJh
xSHgeCA2GQQebDwbou7kmMjSaFlkogKuAX65B9TCeHE4ijWnkeEuqDchy47YmkLZ
xs9r+YSLe2J8l4CeveTF932rUmQEQ11WUOT4G2w9RDDlTH/zT+lfzuIyz0xaA0bm
QgrDELm2ySuYaKV48p1KhREWDDBdqm11nVY1306Qi2iN2VMQthOHu1kt8AUmlblt
w8wzh0zpqKhYp8uSy46Q34ubLzT7zZJ3R/d15UqXQrpGxFyzgcug4plyGZQN6XlY
/F5/pRg6aNG/o0SO4Omd1OCLSw4xSxGphzm5W1UpodpyxJ7tvdyepHDAG1XfathX
Vo0+gXI+mw9MlcWaKVOFZ1bTOKNQMqhuzuE32OasVdmJAAu1FNBNk78vZTlJp8a+
VVymSitQii3Zs8/I0ae0/MkZcm6q4+7x24lTrMl8J81wLPorH+Pe75wq62R35ing
RYWZbs4pVz06x3okNxwZej2G92AgY41c6OhLZ8tSNsaA+AV6CYdj9P0Lkx1ESaRL
47kG5QWcXSZB0iIgIi0Vfvfw/bWEBHT8GcopHnbIKxTZpvzEiPLH/EVZexUZuxRy
95h+kecBkeY4QbLCVTpA+85VwragJtmobvVj18jYspq+3lwylq6t5It0lx/x7Pl6
5sRexzB/ATi2zJBrjnqMz6sxwoAL+CJ+6y3fGpy73bKoHu/kRkUBmTwBjViqClfY
6xJVC3LxeGoeF+CcZsFa0zE9YUDgI1YQJHG1KS3ZcNLNI7+jzxYMJ04SfKETy4VF
JsbFsRvRhZgk4e4yxpi0ZxKr5JpsX+XEehyyZKQzmObdAF32QpaMJgsyLY2SdZ8t
RW+MVdBB9qO+0Pzivip7lSue9Wi6L95QbBSiT738JZb3dfuIU8NY5yJvELNBqj8g
hsLpeHsuS3pfMZevgglapURULzPrxcdC3Tb8HkoEEYlV8r75Rbn1apM3vL8RZXYc
jNpX8PeF1FUXc9UTBzf6w6DgM9uAPX+N3XDyGZSleyek/gmElvA8OXJ6BawfEJnI
SL2xFzAEd4Q1owJ0gi/5ebXCCq35oOujqzffPez++x/Eu92BJAXWnNIR0q2h0kF5
QRAwMUkaMrqgFGwkB1njzV7nu2e09QY94XjGuUXDuogh5GeBI5VTISqVlzVlMtb+
vNCaTap3YA3aJgfhgNmrHQ87NeN7MxfGI7G7U6+upJ6RqCiC2TIAoIRQGiwR07x+
A/IYXOeWkxO9/0+aFH5slY+6VlzxSMOfGr87Elq9RHW2jviwxK+IUafs+r7jVgDO
2R/5t6BkMMFz27BPGV2MbiUGcyz/gr86kuYb/w1NJkr1XSr1bPzBqjMnx4yfNtjg
zWLmxh6UzTwN3ZkE4XOGVIQvmtnRnk/7AMfld34nVkUEgSp4SvIvA6Nq9kRL5s7c
E1wJnv5Kkeg5Urrhe2FO2x2pnypLDJYVwr4zlhECBXX85dWWyWNhUqkzfvp7lfJ1
aYBVxZmzo7hGWAQAvMyjsXH7mppoTlOHoVY5jUk0oTKbicT/fk+Ar2yMq19h/rg1
Q9rjY1d4P0mb/cOp9/ixPx6mrsRz/PR7UEgMdjfzftdrqbNKLoCFjmPmPsaepLrL
g9riKSLd7GRSSfNwO6oX/PyJ2RR5jjyU2iRRFwLhvcoPUNNn3hstWbyi6SrKXOla
IFPYvrQRNfJMS+1hNNRFUqEGMFtrJOMSf/H1tjLtnOf/g5ojK4t/y6JrhbArdq+l
Ln3VH2y6Ru61rhr6/4Wlvon1SWYVnUADtr0fAs4CXGhwaN1cXtq6bwgWflzVI6cH
63rQzaVfr6X5JvxmfX0xE4OeLpnlFSzkPOi9QUKeoJKTSRKMg5Vapx3HpHgQJYRU
bYDeIhEtlHqHPyMh0ujtuI26KcCbmeo4Kr+tSMK8BL9y1QYyQ8/koPveOqTmRK89
Z2QRy7KO9JpBGwNP6RWbOohDj9Vapqn8w5tPOFq78fpw0OPgQ64egPGaEzwfOjZc
jZqNpRzyCsLEBpQXppe+HsdMkf5RZrYpYkcXO+xbmknzTeIXwh7T1FjMltkI9eOC
KQjFvUOChZ7CM8JnKoI6yMoJy8L7kt7+8GeH18O0PTWmtqcd9ELdo0LPcne0SFUS
NRO+aUadbz5lKW7m2tB0gXA/QY2Isqd/LAyqMDa7pGLbYsW+IE7PW/YJbjjaOCb7
HvK27qpW/t0lUo5FAHvpCuJhlo5FRvcTavhiDlCtfB/4rOjszgygVZblO06iC7QG
TJZonLJKAnR+LPyXwH8jvO9Ne90KYs67ww1HyE72i/algakjy0GT7Ob/htVEe9pl
z4cxvYq7ND/t0Z8+AfJ99cXQGujJj4LKJvUezNPEJo98ZxS2n2J7pjl/RHUnqeos
bqiCa0Ecb2U0RUX84LjNwVHFubdrSj3/tL8+VBWdv3TQjCTahm2yDYWIpALb5tk4
Gh2pHcuWsTCwADGiGo70efNedUB53c0lJ093FLzVni0XiJUfVohjJOJTuHjJToM+
crfB2w9LP+6oOSMUH4jo1KojlrldLnD+rdTUEmdoBlfCPaznKDKvNu/J9DsgBcJE
+3h7BWIwwOvKhQLBehbKpCb55k0K8x6jj6cDwG3NFEPdaHBMlPSc5s7a/EKc4ihv
iUaCRaPeViRUwH5B0v+kvj/3D897Vb/+tZZEzYFfsnyizmQVtYKYboJLXlJ4Y5GB
OB6tLcBsszP594oVbF0urOtaIFB1Fub3TXRIrzK/66yJRvJdYYFC/J5mVHRa3oKR
QTkQb5V/dgWxNiDjcIr/Qnpx4khje/yRmHoKMEf5e2S0ivpXltiA5usDenHlbSsx
klLAvMpN4vXtOydpFkW/Yh4v5zTDCBTps0Mc9M6meCl/cq5BpbMjpNfxR0riToGa
36spROcQXwhioJzDLI1/ymw7QcH+naCdZzVjp7U4TzAUNi5VT8NFDJRtVbirkl3W
U5+AFlaf182J37QrzKVuFy6voRD9VaIlLOzjEZtwBvjt9KlhZxVSf3yp+nBnDQxj
AKAxM+xQiY3q2MBN274kGmgwCYaVQOIj2UR5Jj/u2sL/NRaX2qvgPsOsTZksmQgE
vS8STHOaicNjzzouv+wSyJAw6xKcPLivkhb6qjZZYm9dYpt0n+WGSIhlPbmNmjS3
HPxpwZj5A9RxVKet4euMRWkFG0U3tKmm8JpRsQQMOm5spANOTns4lsh9xsD3DOfs
RNYqLNX3OghQMHzGmoz1jd6GBsq4vovulyd1VcBndIvNpfyQ4Nj3slT57D8hqeTA
KdszkvhbowMhKTw+gXE5/HJQ76acK3EwnZPOQE34DkZgx01n2lt9m1pJKE6sG7i+
47xLtcYHKccDO6aJS4Cn50uRe2fRs6aPyeMcOQu0Ymqz8u90uUd13VKhEzuHUIw6
p57+R6TbqZ5cBsnZyoXyz7PAdpK2hEHqJpSDKaM3HIZhZgiLxjYSzyjTI7WRluRF
k3d3mQjDboQ8QP8ilTZzHAwpZh5GqYj8fI0QEHpCCgxYyRen3jJcZeG7moA2fl9u
DQPe8rBDSDtwjGSs3Puins+VGNk68hwdVqJpx53mJYjz8RQkkD0FNbJ+pXOc+pdx
sgqYOoNMrlv8fOA1wu9hLCYjlLF08gmm5tPW8LqwSAMeVIhl1oVyqqlk7nT8jjDP
ow2mnhss4NWrkClzXimNJSl+bxFP3V+S2VXal3/mNQtl6j5cRjXSOhQLme+4Cvip
sLB0BvGkK6x153kAgegakDyncZxANpjV8ylU2B2wN2aha0K1pXiyw/r2TVS6/zjI
7+oEVDyYUp4PeZ6KaqmN0c03DVOCuStge8aTOkX63xV6Zeiy76u8K0+PFHAbBAer
9Ksv8uH5GRF4N9Ed7Kb0GeFUuVefO7rK1mxV4ma0Fni93Z0+5jCgmEwBDG8EdmsF
ithjSbxtG8vD9hmubYz132xuq4YBfeDkliBuxf98RBS+RQSiPmFS8SHSAPfdrsMR
LF3jtNGLOelXMOabJfORWRCdXUUgu7xaxZ/WATfGM1dSx7dUgGYtSOizGzNGic3h
4TU+6q5549MByNDKrd3QXRVT9/PycYrb1okR8XBmy8I1pQfIEJKjEm9QIZt4nDbR
8dLGGHQat11NrASQ6WElaVnBOQPp8SYntqIj/fk/7MqeynIpb/6Ncm+0cwBJjfTc
bErXwuMVxG775NJ9E3vzkxaw/O2ldSG7meoWoQK/VyikL00Bd4E8WDUJs2om4a5a
3ee4k8Wieae22n9mygaSRgawqVSuen2rHYV+7e1/V0+uSw8BkG+BkfnRrTEx3kmE
W/kBrcylvs7x/2KPOBRpAa18o35/3fbcPJqv094buaRI+D6e5/Mz6Vu9KYbRMVfN
rZx1c7T+64cIH/mO7CNK12IlbDOF5XSdyitnFdspFfxo/cxhFN+3vQM3j1ACG4AJ
vQ/fBAMCBI2i0F7YoL/ZrcwDbs7UwANvqQtSlIvr8wgVglbVbdTp0CGX6czC4Fim
ZYJHq55v+aGWXvBX2OvtvVE8NC0oYi5tYoeBOR28p57C46oLF0Lnp2C5P9MNeKBO
KfisUEkxH4bkBP1MNFqwQ2rWXfzM9MzalYZ+0YL/UjocbVhIOvfzLOg0UklXSbuM
+zBu5nNM/xLMyO5MwmtmCDxd4H0Jr/8IL4F9TSz4uDr6YDS3A9Z0K5XRGOf/Mqwj
HKlr+jNCW0U0jsr7oeHupy/DpNdl4nXJjvxSCofKLnztoDHcTJCM+/jUEFHrDGqq
C8viHI60qsyqeRpYLWN7yYTKHTOxlmsajdb/RckOFsnVVcSuQW/DgvOfORg8AKcK
DaCORmZaxDmgjBTfhBwZ1NfPIkNvVry1dUlTDST368IZCnWmibaejTNMtJXaPpe6
TOnm756WnhGADQavineMTuSpyfG6FKVBdmG7HcD9h3Nj9e3xJgU36c25gD1uOj6A
jTdun1dwQifjgq3TjG8RB0kPhLbw7OO1onQV2S8ZTr0KnV6DB0H6QD8W97iFOHzr
qtCdzOfRXJPokNBeBLYqL5CF/TKuzkc6Vnv+NvSMdmkGljunup5sVPMcZYpddbIj
2OtmI20VrDx0vZ9bdAIM21BLEekHqxaTY81gi8CBRHKcvfGRgPhcldMupRSDJASK
KkKyppIJ0w49I6fPuE6MIpCU9F4bK3DCp7UuW4DbLiNmEV33UACkwOppi5SRK2jx
1P40e3fRWHLE8L4wLab/oVrojZx+c7aW1nprvqccFceDZsUzBqBUaGneuCk/QQ0X
bvA6zRAr+cPaiWYbwPaSHnMJ8FSyySEFJyBKFN9lD2+fJ890og9GLtrFuVE8IEkW
yVIfZMZSji6eCllocbEe3GqBleGr/S/UkQwxOt/P94osIUi+0UY0AJWPAiGJfLNb
3WybJD1ge7au4WRvgpJL7WxTXkfe8qpQH7y8VAX5XqjblU9pbBkP1VDe8hixUmyM
Vz0SBq/cdIey6WajO38QnOtG5TlvEWfailwnVnZOQuJcC7H0dpiELhOU5lq2x4LY
lffybfT6t+z5eSaORxmKbEGZkqS/QpjUeijE09f3JXcB2gRqAw8zEuaOdjPADO4G
QbVi+LbWPYMcVQZ51LkYLlfYkyI6wXaI7IMandao4j8qm5dHjs8wyexOewmfJ1My
o5kjmSewU4Lw8NXDoVZG9fgTItdEKtfxwlmLOhuc6e9A32FDs33EPVeP/CrQkEKE
JeC7ysdoY6EE53EP3uEtLmQUudRqO//cjrEAV8Q/nfzTswMJpZ54EDMBbf5o+6BT
pyvFcNzfAKJJgZMAsT2Ag0kLIPYK4kd1R+Szzmw67+HjjeC49fJFb95O74aMKWWY
AHaq3gZBFeMkaGmZF+yZlXeL+yFh+TuKW5GSHdkTzVQ+10L6GXEeQgj1f+z4F17t
YqCojgx7uzAbGIo5ZfE1aTL7zzn0DeCmlxleh71xsOPv9Bf0HGCmLVniVxtAH1IZ
hJgy+iCm91clBF8Kk+rLsyQJOevmVCLildbHDDybFn4=
`pragma protect end_protected
