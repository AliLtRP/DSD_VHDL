// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WAcuSphOVXFa/0qxpRRsFEkNuqumJb4VfjU4UMVGAhTZS80lBUbH7a/ihmSQfCOx
219MYq2JehoTL9Xmw3vou9iNTckvFlJ5Njzc3Ze51l+ICBQR+223ti9Xb2tZGWdI
tMmY/3+hshb0oigreygkld0UZLYSJoTJREQEcsJN8Dg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57824)
mWLPkfwhXN9FYhEhhGGdFOY7eDI25JOXPLgnalmQr3YPu9PSMzhL3Azf+p5877XC
D1dC9C+zwx3Exx/OHNVGLPe9aQ1sgq2wqZNnLWXdsurbUcolPaGMTWNcNu7BFYPW
tQku2SVhF4TsoAnv70c7yHt5dgh8f9A0LmrD1XTqcvd9Z/Wh4ySjnWfv+Eqrga7O
TueIAUFkDxZw5bEJFbco0aDpTzMzw2g+/BJSc9oL72qw9bSxz9O6BNu+ujvSsuFV
xjhIbrq8rOWF+zlXzwyUokUa6gniwN0U+/kKzS301zBJMQhUpm2XbiXoeQUSK701
d4L2juQ4dBuP0Zg5geWbC0nJ4Y3vaIo/nlsxlj0aPSSqUE6BcYbgeDjTN773mk4y
p/7y2/OCa5AfSVO3Deo7EjjXBC64WThZdQeWYYiqiFI26g4GmXjZjLtxGjHu9ydP
39TjQXPmVUjnTQH7xOGvwLHEn01PzF2//6tVIFrhR+ADkRDCOFMbW2qXUHQrE+E8
GFJo5iyewLWCeuUpHHoV56zCOPzE0b3j2iCsIz9p6bwRekhTe+y5KH8BnuZio7ih
NKcotePs6DcAz5t33AjapAhI3JUYzmcY7s5NMeHW3Zqb9lPUND3g1n/3LD9zjBsk
D9RvmexTK4LlDRGW67/2CEJX1MDUq2B03cFeFJ/cPwCK370vnAHOdMR8B/9C4HeW
gRIwSaYwCXE3WUXKNw84IJftGUqiJ9M0xMtRSf/YLw3cAPt/TthZOYTulzhaUzYA
0YXTOoofiiOMDcrlFz3caW+2gWbnQ1L+iCB5sTzmMkErn8BJnEOwsPgXDDl03lab
2Z+IMQgAxL4HdRwoaDipgw3vPamEPYfZWBJW2cFniJX+g0xiwJJZ1rHTq4rlcbyW
b+rjRrtN+8MepMVd7g7bJmvV0huaRI7pnzz03X3r++Qw1S63LJ7c4Yike2Qnk2qJ
Jg68YNIbrWYBRy0boZTDhKukMZm0mXZiPoaZdLuZjS/OytOkZnrYbG8nCacWVXv3
HdFaSIRKrWyLHGAZtUXC9djcYGfFT40uhK9SeubXJrfYqydpxy778yk0fAx87y+b
3lFhA8WsHTviPS2dPQDq8i8PlnL9syB2jVcTG6V5P2VJiA5FpyRAaJ7Ie/y04aRB
sYIC7so+Lg6ekNd8dX2LU5lGvYYjGXvfG/PHwTrId2zwgKRol9hsL3bKBqcfgY2+
4g2OcWO97sSZkW8l5YWWca3AjM4GN+TpptVdyz9HXTEfgF0aiHpASVy3sYcjZ35a
OonDQqkUjZC/zfL3uEp41HHmNg+05IRuZ6gQ/UX/4Zi5LNQYt3hcfRsP5ZvKsfrz
lnqPDacYph8xtpPnMqABlm4oe0E6NBpXZBvsi3tgIFZA7Gm5eBnRoKLULcljHo6t
5EfkUbVIpKenVdN9OpFk/VuIZ4rADgrKfADTvRyPCAQ690ImAMHvQb63zGKC2UyN
VymhT0OoWV1/9+aiJbX3D2xWRELxy2Hb8Z+0kHDHZVaWi9Zdz49YvuV7tVaDDg6U
u6qOpgZlPz32Cc3ioQ7wuf8y/K2wnYo35YUUOdrokC0NtnbcHOqDp233xwjfcHny
qyqauAaoqcabt8zsBHCqHtKVVftBVdBILIDUYNJ2bppUZqVy8zRq77rtMCXarUPU
2fN9VRvdizLQ88WVwvO4BaO4+TNG6/ktSFVRPWm7QAOYmAEu/9q3K7ECdNAGH3rl
h/phrPVsLQCLQKJq5CJmXOoESynhVvcyifuqz/txi6ebPd+GEYzeW6VXiq009nxA
no+f61OwqoMPAiWEVkUo2GNsFybaj8qemAUvOO00dXhPxyOVh7BT/PsY0AkDkZpf
Av6P1aPu04+ijwTjZtENcTr4pvUaK05xu29081t6z7MXyl2+vqkTqI/9835nm5UZ
17iMx+yEF4WhMdjRGOAcp0pw0AkulLwVh+W3BydrDWTYGSU5KVzMrDCoaXBjSQsg
mPCj8C6w/cX15leFGDMtZKbBIP1WmYIP5kxaH7C2PDsbIAyHV2TOviQ92Waf6Jwx
XyI4NgMXtOfEO7cIKhZ4QCL3LwLKv8wZrj3+OUZMR3LEHzX7aPcXYRWJ3R7tD3oj
RBzQ0UYaQWNQ+78+ihjxhQT564iEBG+pPYhYxedaofH+BEX1LWnLlsYSaAyOFFz3
2OXhcsgGQLNBt18Kf3xrbzev524giu7fXuhaJXhhM5uOSDiA/g8h7BhSeLdCQ4Xg
MJfkcCJiXSkzFXPGclQDoym0k10uZg5sXHFJb35SpPSsFkGY4nM1h4Vh51gOM4jB
gI2PaGsjVx7/YpFjdMsfFKkavbuLGP3mc5fHCd7zgeB+gJMhQ/PqZS8S9+65NXYr
W/a79se8RiH6b04+WnTLVQ4+mlLop8erOCgxmMYY+/+JLieUS9Nv0usvXfBRbYcO
7M0/d8mYiXXc45hqS0mXoAyNCt8tzMwC8NvsO8x6kw/iMK8t9m6KdloAKXQjEUjb
c6ChM90nQwJENbiPpX/O7SacQIG2dHWiyFbTYsSh/PlgckQNn/S8wItsj5lbDbaa
n9lXaJ/UimDmKY9OL41OazKRnD6BEzf/ziTEBS7Di5C4mg4doliYP9I8z1YAYKBM
LrA5ufcZbatmlQFjxCyQ+LioGdULPGj1h6uJ0sJln5ROxkBkrUHJDDLv8URW2X71
47qHpAnUQfNnQJH4VYxGsOTnDMEGY++fo/rPPNbDgevHCKiWIU6Xv+IGJE87RTBS
2DQZBY/1rarV1mMpHNQdPs4TebT9t4P7p/pvc2395P0OyPA/XcFGr75NOKLeP9AZ
9pXi2KAOEpPYMI/quVHJsAXP1YxcDL2U6kk+VsHWsDydzXpF90hYkLNwwWJwRMDv
NHCpXpTb4afpytds2WI6nLprhDC0UC3YRY9YrYriwH8kaUWvyWoAU8Uve95BV3mv
OLdY1WCyKjdeMmTbOf7SiTbk5/ajvs7XI9KksnayhEQG/korZUW0dKuxBOLA2Nde
26iRRAhsvumMMv8c5d9Z2ou+x6Q5q/Zn4ibIsmuDPnzo5XznUpno1tl5mxA0w3yI
T/kJpi7VyryCWuoEG1ny2YyCC+RQp0SzLh21qBiyJ8Kgn9ijU72Xj4agD8SCzHez
Uc1hn/IRxsMyrLHh/Mh7k+4Ssez4LtPXQZsVjrCBeXc6xmFn/gDsK6YmcnfZ/rOe
X9Nh7HsPblcaC/GxnZeSpXLA+8a2FuOcM74PHcNpfjehQ/I8qLatiNTcDWGRgjVM
ZNnLUdqKuYttKSdrU0sR2h74cwftp5DBkPbYgnPAjUdGGCTnQiGnVoJbcLgqT+Xs
X+d0h7t/dAyBzDb0n1gcsu4K2Z5XHV3FnAS8rbDwSJoUjtt1syVldyhVhv+bJP4W
g7DfBIPfsJ+j1PCUoDozwQY+e3RubqoBvo7EpzuTUlo668OwwuRQO3T8CM0HVBqM
4yTVocv4qfJ5MLRNQ0H8C80xRWqSURln0J6EFm5LiM5dbn7Zml8hvJjnM+L37jZu
iKvEI5ckxVYLPsM6DDkWJ5xuclsNNiwetRrUcrEbAC6g1Qm4482jGrFhjxnmP9JH
vlDXCC5ll/NevfCY5gBKAtGXUtBdp5DJnUYnkbOwUUDmxGXBXVOXnn3tPydWq0Sq
vQh3tE3lUEoHAMjqCXs3Uarf9yfsoaZZUhpQwimoA0LJLx5zRP/CdBXjFR2O3a5e
qr+Zz4YwGN5/lq1p1NtHbYGWsbNJDcE7T+9BTtZCvvBHrcpFBSQovj2Ntct09GC2
puImv00rneqkIai3E9Aqll9ghyNw7lQfc84HOLc7gw94TOsT/P9Cl51+t+SVXYzv
DdsCsIFKV2nFiHhnYt97LNpst4NaPOeCNB6hbphfpZxGzmQgLoxNnCtxEU6AmCSi
8jUaXKi/6LTsF5+JOBk+xxS7CSDequ73tn0pPzxdIhNDqIRuyC3k9DiOPUGMTj3F
WBAqH54yWWeXu+iM1Tn4hYAsoNqXU1gh3ALMgQepIa//glMxK5o/aTNHtXOta1cO
R+EU3Nnt5qQSnC4MiSdzrqEIgfNOGKe3nhvmEpkrKrIKo6r18WLUV+EXUQ+yAG5l
0/4CjF7lRYDMa+ZtMAXrevBgONQ8BfydFNfrVtSdU41iW12LkiAb6HsMdlKm3Cdz
SrOqD8KSUElGJ5fJcYJTJC8BHWXy41gYo8dJfyk6r0eIKS5blLHMWXDnam7Jw9E3
WD5A1jOgu3XlNCYGdBrVaaoU2PWWMpVpEGd/Skle0N5voxQt6I21AxYRcHtqP5CW
13A19WmO5kkGOTKDOunoGYWJVruBMeExZmWPCjSAmotHD7u3SPBveV6eKJTIpyLP
KNhCaTXwlRLeGVNSaRE7pKQampu1cu0VGYXO/HV8DNyJCoPr3lw+ne10Hz6hqd1S
stRKtZ2S8hvZHe/V4RF+Pm9DKKzBCEr5s47HbKXgGR/yTgycrJIv3zcbJXiUe1v1
TZqfBghW+TOgx2c0ealofhNdqHpxp762mRISDTATILNGmo3gsCLj5T2nJsr2k3me
6q96ns1UQ655/9BvlFP8zu04h2IAipAahdbdL0Ux3a13u36g7+etDxZU6XnSvMs3
nqx4IaU5sdN6efhTKzQVLtpdpbbNmovFKULo5pm86upQ9mpHGPc2fcXNFXP+Bvz9
mzsj9/gezqeuNs86tQQ/2QYpdhT9OrcA9QXMGs1kAzUnM29F1mWsuHlUAEtikFvP
sL0SbB248XwXYz50CbpuBVWtNoinQEuLOEwbvOjavLlHX/eo4lfl2zXOMNvwrfJ9
tDB5/asc0fTbnPM95sQMAQr+ZngBN7ykPeWPn0SyZU7ZXgreBnS4RhWENXqWmH0h
aMybKWVxHQ+JKxzEoLhww8F1h2Et0L6LVpn9+lWgpx3+BuG2TzgJWMjeFtJ6qrYj
ck3ZJ3Ch09T00AEZxK3I77B97xTkyAnaw7M91yBvKeyilXgTNMxHkLGe80IplTWd
SGWBi1ITHkZwKzJ074tAr+/LvlcagYGk46TbK7Tz5yBGPBF+NpuNWQgRNymA6Ho5
/njAGDQS8w4N7C182phK9nHhCLs87OeEEbQNUhRir29tCSHYOVoT7+LL5wihp04/
aaCnMENIEB0qqQxhfY1UdUHsG1suGt2Y8FQ1ZPZPwK5oROVlrAbuIP9WnMShtcKQ
WgKYG/GDtYQqRmaJ6Czbsmh/1EIF+icbckCocobBt/KI84vltdUKXPZHEb93shPW
zRV3w9o4ZJKyn12Lf+se0ri1KJsp7j2EIiDd/E8y9mjrhZ/awkQ5MKPJwFuk1j+Z
lZxLP/JRGGdRrcx5Z6ZgjW1HantP2X+9nVSh/PS6PAsDfzF1k/U6qx14BYPp/frM
utflXzVpVT3U2e81947sz6zRXr7Sk1DgAPJbkBF/5uIZqxAy2M4AqtCwbeBbclXP
rWJ1KJFTUFDZOY/+k0OB5nxwbuvr65PvEkBEw/sMkp9iSREc0Ur2f5cqTwr+Lqxr
Qni/iSCqRd7zeWm36uif1fB3DBwEMl0M7akw5LNqXBG1yH/zeKfaMq3bzAJnQyt9
8keYYuB/f0GgSG60FJuCIyz7QIeKPKh2CddoMbisk+XQJr63jqCfWlGzfvyxMYKA
80SCAy98gyG/eDBVF+iSFqioqnROlc9qY8dtpiiIbRA8yoaSkcSTeAyFNkyAUfLh
VfsLXNawLT23r5CYF0JP0uU7oNU0aS+dZLUKql4UGzowsWXX2yllWn/UuD3g3XKK
k8EjLwkY93GyjOfXzetA36Der2MmC24IlMAw8U1b6lrOp9/xu/op6nuv3XVEkFqd
y7RP6hoZPTfEQnUIUCLJHhciGLF8Kkwq4ESvIYSwpg49P1dzS2KkmPGCPR8j1Obn
VpLAai8GbyxM52ftYDNGgh4A3JUSQqaxz7XXzvkRxzc9gtptJrHgDgbPsYiriN/Z
P2X07qVCcetCk05OSc4OUl4VEnWcuOYASL6KnxQw9bB+Y4ClPS9PzDK5A4F1xtMX
A28ZQYse2SoF+glgbdxwS01istc0OapwMfN87aZpHNg3kspbvVJ0hHTd9eNqg+/n
qpIYTknIKOhyjIY1KD8lnT0R4f/DNIE9XVJIzS6dNtG7aLiAjqJRO+BOgMf1rFX7
Fv/CEPv/HkE74y8vFRg0wWoG9dj0d0Ennt3N67p/fGFwwmhFjIkQmGy/EuloaYBL
mGwNdgFJeh39nw9cvbGOshsQOisjChl3TXT6wgCM44jmSNGj5cCBw0pJKLfhA/iV
TS5bSXOOaEG66pKXtRzq8+NsJyPwxbVDRHE2z99s+suII+tUOQotAh/iMpLDuKAU
C/s21BQU4/+idTyLRdohq4Oolx68ofohXxhuuGYu2QdQi6JiFL+J70PA0MmfRkOK
rPel+J1C0z0pLBOYI8rfbuVZ2ps8wYV40Icuhgt+QaEVVPrFGh3IaWjGZUnH/HRA
ep3V2lJuvn6sGPDqMFf6C2F+jbwC9or9eI0CsCBmLrjgiNocEnEBqgBunKc1ihL9
jxaitM0Wa74SPnyNMxHurYd5kMLa7Z8fGvIq/ghhdX9jKithbDdLgqijZiQgJZge
GvvieEmnEUqGFgReeXtq7rzPD95Uzbda9m+fEPHNZt1IIvDWF6jpSBa3QrO4JqPB
sFLk6phSzkROnQKv23iUw8ASCv9o11IeoJt3/+qrBlbFU8maM7Bn3KOifMVB+vfJ
uFrRTInP8PaWnstF/DsYZKpMzzKK0oy78y20/Uo9u8o8H9vQr5tbpPfdiWQZN7iL
DwDm7AQDeuMGRUs89hvyl6AfNjeX0bmSopuH2RPkvAkKLXnCGYd4Drtf1Xtbi94w
Ef9y71sfljeL7prdrAMhIWLkFB/JqY5rKBmYWgIfX2qobRlq7bTcQQ5k5NEMjqCw
JqHb7cQ4v1B/wXIuB4sUe19gAGWKBHn/3AsJpGAkKlpMnbM6BhHDZRdi5gCsv8+O
QfpL8yUojhwF4M19AIk79CCaVMVPlLRtsR1rqkNgC0/XF+iu0r8Rusd1jCLpMAtL
F0S7nObMdPUWz0R4Xmhs+JBeicAIY5PxEf6VHGVNSfDgBz/zHtjhT9OQlZgTbA9C
hazRJLyZdn9xs8eTr/50qDpOLJEdZuC+7SNjrNPHqlmcW1QADgBQK5f4SUGbiAQd
/3u6iuSYMCsOTq5x4loAUk+LZl3bHWfBqWLDZJJkcw6pZ8K8HCSJlEzkw8bRMnyX
N6N1T9QvT3j3LRBpbDxVCjxOV9mSHzMFIY5c5txyQUtzFOciUWUcgzRRPkZUrww0
lyCIhwpgJhhcSRO9MsMUnZYF0MPCBdutU3yMZZNtK85zPDh967ym8Wh31urSBlrG
0yGAv9yIuE+cVidi2/a6u8fcKnvFk/c1yKZ6JhHDKfl+8qYXZwax5OwRg1Dn4UIc
JDfmbeegq6kaQIRQaLkXb7d27JlfcdL2/R2aX6jZjVsHJyDY16oJFaJfKb/74MPA
OQVzVeHK5TD0tB2AYg65/ErU4o3owb4J+O8NBhET80dHHK7H4O83xhG3X1j5puBe
rZ8eU5ZD3IUtm3zhQQpyRDqn/8pSXxUnZG7L8WObAV3R8qWuF3u0sCvdljKCuD/Z
fp+SdHMiLvGyV35GjEOhU3axHLLDcViOVH/cI38UgnSn2B1SfGdKy4XpfpbfDHP9
dz3f2HRhq/vBEEDjpcyMlns/bRW3kvnDgxhbIWI1y6hA99PYGfC1/15RzwGXLtle
FLBRGGkHhYpIS+2aMHTVsMEFmmLo8LTSi4AfZG9DlnpSPy3IEWWXUmGu0wvm98D1
4FoZpETEk0q8Dvuat5k7MeIWGWYAfCm61K9Vnik8svMwSfdMUjs63IjDBjcXdxTM
DkycGGcvAJ1E25DWbR5uZzGQpPmP/mhDdt9ManmTYvNNRwXgdVC1ouHMtMm41eav
WQ2sDyz0aHh6qPvX+vebRDEHd7H/VLowtO4Pwv+GxOCtyBZQPjQmhN4d4i4AmkYt
lf4fi20Wch2e6Ie9pPMoSQP7EMQvWrMV5xuV9uCXZjlmweS0kzDgCVOmHy74H9Qx
U2VMzHuNExtSpu31ixyBMAG1+DCjoeXB1fQrm9FL0Ly9YnLTzT2hKntUfoZl7sN0
fN7FNzfudj1PoMdpa8LdYJBVI7IEUTiB0GwrANlTS8hDJMtAQb9upyzLEaq+RaPl
BB54Gz/GMW6Lf5gCT134uuYXNHZSJcWlEHt7m5UERSTnNLhy6gl9pr/YDazWDRln
FNfXxobFoL+qsRSlVOUDYLdtiUHI6K0AmxHoy1nLqRvxeGsn5Z068jqcjcsnWQhz
UBnIGI0vgy90mDnsYK0ofzVNZcCuzOsMdF8DlHh3viwlBkxCdnrdPUX97ASw+VjY
V4UrW8a8YM5/GHigm6Q+D5oCQ27Dyruw4wZUCYp/RkcwTzK0Tq5iVKtKI6B8gaEy
UMQk5wly5q3+bboSqIKm2B5qGeSjQ+bOR4MW/bLuGmex8K3thvFO17T1LTuU12t5
4L4O+wOiI+5vuOkp29GosBZUEYUZngWnAzAGxmScstYIFVcskGhPmpwqlsci7uw6
T7mahuED0QPNwBJU9Qy07lJZjw/E0O2+fiFKXvgqicEdHQIVM21kzdm6D1BTwgfl
M1EPeeAz70z8HKRR2bAtErjxghqLMGEcnFhOMEpknN1+uYBce/VCeOo2BwQfD3EI
S34E+IXWDSJpsRnELsGsQb3A9JjvVOSkK5liwUbAivjvSLD0aqW4jkwPzK/sB01+
E2tUQhPFsRwQZ9Dn4MVOC86ybL+Q34Qq6L6mQlcxuZ6yo7fRgdpVqqsgXsD99Y75
TD5cCsKYPnl5ndusKXhMUOp5xLKaPvUKq1H1dKl0YG1DOZeIzemVD0t6I6OAGBfR
o73jIfOGA57o5lY2VvM4bcjqW4yqJgSVPsCso6rqrI0BnsKNCe4SDm7buV6L0E5N
n3Xpi5Kia7bJsEt/z9GuXHER13lgsTU58TPNnPkiWxKWueNUetE1+LBowqDcw3R/
IlLQ6NTIWZo699CoowdBkok2kTIUd4C/xjDdmvWL6f+WTH6coutoNDtH6azx5gbG
9BOYyMWDdoPTrboLzqa0Sqc9zzYkZEnx/tOPNWlsz1X7Hhf1SK/jypiwZeTR/XV0
osl40actzuzRPDl8th71xtje3j6l+4GP5sUMjA7DoXEmc6gxe4HBj5iuNWd4cHEC
NW7/uB0dNGR4SzfDfretUNHhP6c3boK7xNKsxnA4yFDfRQiOuB30yj5bZy+tKAYU
GQqlIfriOScvXyRSe8vRxdcLTZ0ILq/45lzRotytHRxVj/pT9ySFPj3QUTnxM5VW
ZSSD/rKQwRa1I4kh7Efdwr2ceTWmzvAdvCS9Q6Yjd501xdt6hv8hPeedoElt1430
J4+OS2My4Ve7clSCongktCRecCL8G2LAJwjdZ48oH1hMQ+MXzSsrtluqx5G8Giba
aVSEoXTcOhq/fRlWMTOqoyCFdjNyoS5k8JuvIGnDhx5pk+NKXqTb090/q16nK4U5
b25W4KSPPMZ2WbTOs8hRq32/41Uz7iUGzHCx4KdchjDY4Fajs59exgNhoMjHCQVt
SY90qE2XbhKTYQOa7IMI7rozPYCuM4xFFOWAw+znY8sz7LK1dkwMMZmRlANuw+/K
CEQOrtUbps9rtlrlWJZR3irwk32/tzngNP+p9JGL8Cco4nXnga1E/OnzJNCgt85C
pm8edqljXuDtHz4+g7lI/xVLoxv16gP/PBVZZk1oSJOmfQjJh6LgRi3zy03zbQzW
X0p32a/HY5GvBcDleySxknLtieRk8palCpX2PzYr54riZ2lcmMJ974nH8/edfZyH
stgQ+ISVsMPFE1ylojT1GT8NZCsJa1hLFxYKYaJPNT2b+Mcl5CBhh7A7Ze6wzhcy
0iqvFMOzak9Lta9KH416ZswJ1in2eTxMLmKceienHdfEFaHD6SxLN2FazVCU6xzY
MH978z5qnRJDVczKuegGKqn1CPgUiisLUCwz5SECFZeKj9AYFsSkzgt/YeIWb4bF
WBG1KtLIiPl9YEJ4Q0Zcr3wMn3RGr+XsvrERj6nui2a6MiOR/TZq65up8jfogKZo
sjy483lnK6fIluuOn1G5jPZTPYyexjBfmRomtUXfeVGdO+thvt3Or0pjE+1VRvNP
P2iTE5IEjXnYCj80XQmSl8naJ4K6vN5JcBJT9VWBVnTBVoW976eDoMbQ72nsKiYj
YEAecvrRC2NUS6i/+iAlc//agKzqVfnNkZ1WaGMY4sJafnhB1YyEJgLYq4VtPNqM
DJhcUqYgxx85mX81V5461klfWC0u2rCZP6WlxnkgSAvCYi0+2Wp3pDYzUyn9TaiR
j3dz0JCQH+uw5tUcxKcEL7fJ9I/uSdrBZcusOC3ESnxRWen5rAOSner4t3Sxo33f
aZQ3rmhW5GRNj3eQgyvGHK5ScJv5IChsMq5mLn36Y/ShqUZi/DD55UfY0BdUjNau
cXxpdaXHld7h81DRjcXPuEWoDMDzjHjzld6JqA8Nci7CBHH5wUt/WG3ykqv0knA5
wn+vjd0VYcWgTQkaJXpA2rbkH+arY/nsOgR6fkqNt/50ihrmv3gAmHWp2tCN2baC
j2u8Z1w/jm2pbexAuWClY5ROcerflS9bz9wREaoQd7F+YCcke/keORS6FOOSXWkw
gx4vdSOdzzYYuG2l04P8KHDbxRMh7kXWzfCf9pWXYHuyeB7yskL2T7yg/s06nBXv
03VSEtw5jXGsNAxO58/quMdoLNa3NAvbpjCKt24xnpburadYc5DrU5aoO701dFQp
kNFsK4QSR3BqzmcS+lU8FYzD/bgi1GnOU21xzJpemZVezmR2CqrbLuBypveB/mnf
VPMoJxT3RMCLHXXFmZkiM96asIx2dMstaPxQ74r1x07PPwB9D5waKLOZIIrJRoqZ
sdJpQHYlxzdGFSzbPIpJnCbICggIXgTew9z6TcM8qHGw70DWaHge3vJzc+t7zmWn
WAlY3dM/2uEC3OWF7yD+pbynGNZ2e7w+V7QVn9oWpDE0vTXI8Qq8tB8NDFeBZHZ/
aOt/nAvI9v5wCMNnC5ANtNKfdXeq6ix980p8zFg7IffgdEOotpCIPOLp4DFVc5tX
6+NK4ft+kHPROdkD35g3iO23VsrfVBIgR4+8jq6sHLl+YO8DU1OosyLEYbEniSjj
L7WietkHshopWHiYA1pjVZnOFu/8pFFsj67hLVgtgwFsLrngHQkDYDjrrRiE9qeR
fvUgA1iIvvhuElev8xjlmxqkVPcnHzxsxSASdj/H7dGbKMbeeMztG5+Sf2LWapOp
lHA/dKlxmEljan882eRvplXLNjOSmvqvnpKtvOWISAnFGwAPHpXjtSDxnxm4G5y4
w9+kAMSU5hudet1UwHTQs0ZHwul1x/TFNIbMKFtdCrGvbq9Qq+qbWh6qquHcGktT
0AmAlZ7zqlU18QTQq7qSO1r/lkAdD0MenNqX5CQvoZrYQxpDrabp6YYZkXyVp4QE
us3ZMw2G1JBnqDdFa4VDpTKJqCcmwYTekXd04K5h4u+ifvBd42QxOx5x+YFN97Vm
Maw75xlZQwyKggvy6ZBicpaOmDrdnmN+dbsFIOlWhH6xbyIiF9mminF6e7GZY9mr
5WXeDuCwl8Yccc91lmhmMJROhKaL2vQXgFlC6ONUphfQcdRGI+/SGNRvgAS0hmZn
gs1W1bp0WM1yROTcWdJR/aLP0fQwVpbZuvr4AhsVA5hgYFlQgTBLHVBOChn9A6AJ
pmwzLQqZ/RX/5CJwGlvYRXdC17zGR+653S0zDxEFl5yx5lgO03LJZJglMb9bD2Fl
q6oJN6HNvRLU+b7QY7j40ntLp4VZvV7oYX0kMWciSgmahtvCV7z3UHMDHb/WhfDD
pUaf+mgbJ89Nx2Q2VACUu54uNfXUvMph03U+sRqPQhoF/qKlJKxwnN4fsqmStwBO
lNnq4eGYvJiO80LcyV2+XLnVVmPyxMCPjwamSokGpCOV06cbV7OCrgMYhwEuqefN
+Ls3Ft0nzmpIPqAkmcNuJ9YESwL7rFnNtlgD05vU5Gr2CEWCrCATT55PDZ7emi64
sAn+DqzDUmZ0E9DZij/5gR+P9XhR6D2L3aVDW11thFRhcJFNK6lOGlDaLMHkdWt+
eQosqolvjY8OH7/4DDIywHzvxwtD5DuNDdIa/QAF4uqLe9+fesl6qVOpJza648Ne
o6FoN3piM/zDorYTSrrUAXqz5/eVJC50ecoeXiom+0cdR9A5CUFHJshihMRIrzcy
oH6+QoMCzsknVAXJyb8sDNqsNRDxQR+Mzv8FiHgc2kWxMdNVzKZwIORaE34MlLqV
tar/Gn+BffOAyq619qVgRngV8/fmSnzxM46B7OhkrZLkVXsVttBKjyyNJfeNV7qq
pa1QsoeSeAGzRCRv3QgfHscGvXLtkUIFaOYgWomCa6NTL+9Jzp/xQBcHc8OBMTAa
pYHs68Fn+oKUNBYsl2PyUvPW4zllK6kGU94EMKERK+aeVPPfNAfEkAGTSLygZ1jK
1WibOFODjqXSLNVB9oRcx87wejYBNxXxRXwvlYe78jK8ciJKqickedV5qy0zEMTn
E3nO8pANJGRVakAm5UXvwycOuFIWl3TB6viE2d7SwgRpM4t+FOStZzdeQaBiRbRk
59Ce/2dwyeUE0AOEjClwxo2w/37LKkfSljYUJW2eDQ9vMbD4gQyLpd/BEHZ3RBpM
RBm1SPDrGM4NVQuh7dA7FGbh1cEzldXpD/y53XK8PFgSLfS1yT/C19M1QpWDxDI1
N632V1aS6iNxPQQx5kVlPpg9AHOE6PD97ubE6Wp7mWbz3dAl2o+FgRDdjvIW4u7a
YrEEAHc+4iDYIDDNMZCYyx/Ky4TMcKN/Ao2pcXbiQL3dQl1JFYfjPhMwmIqOMx2V
Rp/o6bDgmaly/E6w+lOs0L2TD7IJ8ApEJajySHjk5QiVGoIjerCm85wTGXcFekD2
eb1Y2eEiqL4qBIgFrfx+BT3iaa2UmucYg/wmWwYjU5CBR9HzQwtSBpbHg4hifdUN
21ooRSk59sxy2fZyt+YRxJQbgrPHBVGlpSwPYjTMDPjndFzt3ueM4MzO7aFwZByL
hgEoT7MPWbtzRutm2mmrKQj4ROpH0YWx0dOi5uaXf/uI8Lt0hIbnruYoN5hO+NEw
UrcWhYGgA78FrRgIs1cwxUhvZixD9xFAKSfP+RLgU523n1cxY+D53OPZXzu+XdH0
kYDMpJoH6LILklJ58PrGDFW+Ucbm9GWOAFxRSqBBg0HVZuFzLCMFImkEyT0yKO0i
6Wjhyl6Y/A9DguQx/XMqR/uXCpNGi5N6h/ATOWqMKnJL5D2Jv0cMgAAoXntsXd3u
WTGW83hTwDTyQ/1my0aeXM3xbXvF+KgS+wpklht7gqQEikfKCXNhSJh3uIzsRDSO
5uAmievIafww+3QvkZXZUhsdK8ox9CgXAsJ9dLMKjbFRlP7gkkVUBd4l1EcqLCZs
qmtJjaD37N6a4fPvDhvQgZC2DKBIftyr/SfUG9aOFsA8/i/SJchpebZ2y1QPAtjs
WdUjW4IBQdbmLJpNXQeXB4855Gc2jMWtGZ8EGiCjQlpofcoI6cBbrVvPwLbP8+Iz
id0jPMtk0eXIpbQFnB+m6jo0034aZQ+o/x+cbquPqMCiS4NEIFVGtjLCwLAL+vIY
6Sv48GrFEjRgIpFI+t87Fve/i56HlJ4VFwiahm9MRVOBartrolGIk/ZoYpAm5kVe
yfPcESZ/L9/W0ky1wHTZb3UKLQGh5+8ySXT56UbpJEUdPiHMCJsgRetcopF1ANRT
gseB9dKIWHy1HihFis+5da6ciHoSTl0hZuKYd+eNPfCvKFa2D73W+QXM+QzJxqFU
xLAyaJvqzMK0RU3Ke1cRhzqp9U/wFmxFJLHAeNHXt+TDvx59iu71TG3LENAQ6EQi
pM0NqHYW0JYtvgfqLbu4I5pctdztehNXJtkzXv4w8oOoWEvKSun0cv+hivaxa0fl
YSLyAFpfPgIiX5oI2LiOvOHBM4GIcBotqmCMnsW8l2hhoMUbzTcjQJbSPNsfuDLK
866Jd+8c6xxTb/RLQ1pha2k2KW3lr5pHMcw3tGIfHHSBpzwuonNmBoEc4caPr+f3
MVc8qL2yAhfb1HPqcSYfewCnWCbePiXW4bVV1rcrhdqxJEsdsGpEUbPf6huRnwnx
qabeOw4zRRmBH7bVcgeUvEA/jJk7bAT+e2VgaGFNfkS+FCdBzAabUEdqE6VNVynW
RYEpV0Ix+a6TLh5SJO/mNCBUT6bDVeWEfNG/VMJpIwuTaZIa8MLe7Ld/K5yih3td
GyxQT5wqb/hLzmZdUyO5dduSAxAFmUC/FmQ5KeKB/Z7MO4OzLGb9p6PDEl+si8TM
XO71rKJ//k/9h1iV0wwtq9SXAXXUj04M0OfryF7tEbdPi5pVtk8DHKJ9ZlmzK7RC
9WyuezjQi4QGc1QqWVEqsLZR9RItsLVD1sZrgH9B7xbGoyg8VEJsmGSJ1dIyReyV
FtWOrwSwHK6kKkc8+ypuQt+Vin4dKmDMHv+rRhGCFMBxT5B0WigrVfEZh2cvLv8L
59abDpnFXJJkqxy8QEZp2mAef4ht8m1tYgUokFJeaFfvQ216O9kmM7+CpZaSFYFO
g+Z25K1zp/ymzlrmgd5thnPBIpgsU94OJl7aBbx8KXw2jMmquO62KzRt2uIFX0Fz
pl+KJsNR9RhinvphhIjTQDnoMTai0qTrICPI1tc2W3yBSfW70AyD05ujqNeVumM/
B20SR5xuVm87EgHvkQPVwwherGm3FZas5RS4XuWLIPXKF9cViRJV1S+sSIzVe4oO
I8lQJVVg8qIlvEoYaX+OrXhHfJm7Zqu3nBuaRYlUZODSejd9hBqltQQBhGJ3xaxE
OhtxsGoz/qxoCxxpG+WrDu94kLIEBF7FbCgy1QbPnPAE5dbQb2E+eeqPLO4Ib64b
4fsDHIeK5S7/dS78Pb44j6IPF5mWh2ubNOh6CcgfuDVJ5SADn5dlArzoBqxPlLRD
06LwqqxhVDcIX5ka3fORStgP1zuFk6Bc3wKfvaGNFVXVWF/x2grer/pMkwTsZsTH
9UMCI4IPbGmif2UHiGqIsVOlClsI1P+G5tcW/WvTOrBpGOkxFRLOy8XwN5IevuWT
r4CN3muEeBSJspdjoXcyXrZzvh/Tj5qg4lyHzHgFPYGN1pnpC4jOddCeDpPJTXCv
zMBBo8JERKVY5KW2s00Gseqy1sjZ7oq07NRYtLGJkBgQ9pQf0np89p730/OdqukD
xJk9XkX6jjceIe2gISim1uEeLG68XljfARJeRRfaxi/JkoWl4yEv/SowYFh4zNAx
D2bSPoDygoa4AS9863N+7KaJgYjdialAog8mkxEyGLYMqGiMSUjUzdNutxD/P4qc
N2JHUuzAjhQRxZPXfp853iDMcdeuxRQxEKrS5Bb06uj7xgV+6qRcGJ0h7+c9DIYV
BW3tPEWq3pZMKgyWd0p0hjKA1Plbg76XMHec0mYpHEOjA70uDHAuGpPHTVR3+n3P
LgVKsKA6Mz/7DzzsX5WfKS4PQYIXju6y+WDj0OXNu85Oldq4NJz+orXylUj5sSUM
naZ2xBgxu4m2ex0+TARH7+I8WchBkEHliR+mPC8SBD3CTOY+fqwadaEOf5pl4RBv
JQ8mQOMLMMRSXkYSBgVvH9ElhLmLw/Mr30mZUtwEhaBTu9b9Xyorh3OpubchZK7V
mLydb4CKXFtsTVDUOFtBhuXnFer+/dW154jeSCwT9cuf4NEWq/ECxLlBQuHB86/R
HBpPt3zLUljmjOVq5HtDs36ligGfWghBrCysLAQFEd31X8G9zXgJGBkWKP8mXwQW
mbGjpAL69JBR9kSioilynqoPW0zt5S+h1Sp+ox3PWGS6VlTYCNvL+LL7JumBEfJU
nYg1DlJj1VyIwuG/oe6d6SNF3fP3wzcj37Qd0UHi1Gm6Ge8tOe3LYlhZeG4su3lB
CvyHIgy53fPuOchccUlOHHFaPJoF9tXq7ePmnapoVRnf7jTBM0W52IIR51DHTzz7
2htvQ24pV7uWcEfR+1FLYD7bNOMvEszDJe7uMkdt6lcbfcAdkJK9KCMyTfYAe8p7
XTTh09RdojyJihJtPRk9ZQFuuaKaP/JJA9lKsx7AbFQXInfhnX0w8RK6EyMZ/X+T
jNoKw7+XAubRpFPK5oDah+cu2G2LR0cXA4Uvsw+EskH+YS3JwCu+uYaoHTQRJnIV
BtGQyQZG27CsuFw9i0jEWJRV6Us/z9i5HdhPo+lQuZpH2XUruGDpXs9da5hfowWY
ocOiyQ5cLqgECaz0BtE61xIdM+fkVdyTRSIUbbsHU7ZKmq8TQqqhncJxTCd4K2Io
0nwgMmVQgvXoGV/cGNg+3Uuq8lDOsUSfyDK15P4Q74+GC/a2lIvWA+reXDsfNo4Y
Rasht/UfF+BdCUHtwYSYkbqBvxI/U+qHKvN/NSAe+vzTlctZBrAtpS4NJYELxR8F
oobTY2sa4lm+pruQaJkOcf74g92OjlXFMBOqTir+KaDOxwsIo33YliF/9C2xXu0B
4GdedZyQT9jO7pMMXOplE8EOzFFfqIapKP10ZktNac0+mMqKmujwqtsiCzMg6CmX
1KcAiOG8BcOfJ/5VX4o6JApgsZl9woazDkDHlLyByf3EozYLRDiCAWOMkt2cotUF
WlQm8x1HVdYK5bmeXfmp99jTJc4kfkinqkX5iE4T+BDv1PHvJgk7jgGHC0CAOPux
OLOZxT3A1wGhlKWnBHqSO2nZVibJP75n5SnoNXd17W+qv+Z/zHbtqQGri6dYekKj
9trnMSt2OmQybz/F2pYUGfgmy6ubjn/dgHyR0hyzvZiTVvjgNqbyzdii39XKoSpt
wjG5upvbf2IJq4W7jEwBHLvxkXJcxTq+UjKB+M1rMzbn9fLZ5ZB5zp2EpPjFmWr0
YQLrbAAqpi5w2sqJcRInquyg1NqCg5TIr3d34c4EZv1WW4h/IYDeFZTR0cy5swhv
jbo39J1TYBVR1x4Czsm/5V5YxoUB60xA39SfxuEMNABsvPgFUn7H7GvtBUttK8Gf
txRHT5FFxAmL9HT02q1QiIzTAPkR56ZUVE83hPFPDvYA8rO+UeF08an2efyKf4Yn
7UQElp8EhUiGNPFUlpUCW6AM5Cl9Y4oqbj1lzf6AFOtAgDiN5GVbfZOXH3k5sqVG
tzEg/MrFW8ezQ7Xe2QQ5vXrTXxJYSFh5tie0TqBuWtk7pt0/28xwmtjvrh2E/duM
APNhFE9EN4u9FOgzGO6U2DmmAIK6rtJdoEoTIPvGf5GdV+66I+cH7A13Ukw3ZMnn
nDr323CJudM8uZCuSB8zqVGGV/K2tRtqMVoQoeYFg5bWL+tS0QqW4ajgxUiSyBaf
+tWvSYJHSl6+0Cx/sNNpiTYEi6+moKlk62hsEBcZWUeuKCQPwAtCjXMImCAdmtWg
gyeiSFMtYsjIr/70Iz3UyEOibrAPtqJHxW7Kno2VKHeK2AsluWhY+wPDL3dvOjh8
k5k6XL2XHLC+ActGB7MJJv8yPjYGsl3WN3FBUPW+Mp+JStYmOMNqE2OLg9EuuIre
hQpctpzybIx4P6HUioY6c3xcbLPWo7o2U9nJKfO5jCLmmKAtaDj+IJ8ztQugVpRk
55p+O8zMJ47LYQLipOfh6naKK8ZJRi+OD15SPGzJL7l5OOV5G7/TC3DJztAInvyl
wJavI7DbOUOWlgJvZyNLotBavkklk4Xom1rkT6eQEy1KqEEvMmuhcU764PuPh31c
Oz2tCT65M2a6godquMdXBqfxST+LvhXcp0TKCPYIeb1lCwjpCHYnjChxZb6IPZ7P
a3oghrVyJFytNZJfUXlXTG/sOtXjBtiitR6XTS52KFRKjq+Bx+MytDmqr4CH8oqg
WyyttCpfjnE28urrjDezoJesB592jN8aZ79WoSl2urIvBcKgdYUcRm/tVWmFOZxR
KED9vvVE5xX8U0qUk0r5Zo83kDp6kYohOcnWhfgAdUFmXHWFjZTliPABxNFktSoE
tCGBOM2IqKkLbjm/sfEDtGWTXQKocxfHmsbQzv5INL2IpBbHz2RV/1sd+w7PUw2V
i2VxVUI/l1pCFgFJIngPTpPCJmwST/+/5Ndna2u+8uzG9ibcILCxzGd4p82ZEcUv
0e82i3ZrrgK1Hvpy4xArE262F5JhO9yzn5lI6/AYwr6miCA0u4qR1aWrQcbRIN/X
3T8cBuo+WypIONX6oHvX5UZ43KNFt9Pg9NvFRyadvorfqcy5WH7nEgihFBop3sMZ
2m3SeDwZujTriqzrZLIuDID5dRgBm05u7HYp4kapp50hYpXYTel3BDA4Gr7gpdlH
HiDrYa+E2siD6CGNmw3+flY+NrtZDoY7XOsCPGrTuJAaTKj710X3PLef64iDO9Zm
auxeN+PXCAgkuAP7oB1iD3U6TptvhalCw6e09jvBt+Vb63Nbc14a+hxNC0LO/F+Z
BDzyG4qOsgq2m6etGQCKCeS5/rgPLXxRyQTBBf0icJzaegM18kyLF/TpkKgyGyA7
vJqujCSHzGKqIm1jf5o0gDaRUN0GsxVvfL8TUXvkxLqYvXqqGOEBbVYtpu8fb2jE
wkBRS0LtHw3BQ2cwTd76NDMjOUAwPS3byj7EFdc5H9XMtv+/F3EKriKIyVyC7LEC
7C6v3jOLpcGjr810BRZY9Ld9xHE/JLBcsIInuBdfiKE7Ujv8Cx74y+KTOFhIrDla
hdAwvtS4B6DxuR9so8L192rg3n3ogrNOFMDo6HnEIBPBvaU11VaKjGXYq0pZWtdm
DrQuhGGKQAX8hI+1g2cwzHp1EmYcry5zTxve4VR2Zz1NQuE4h5V0pQfo5ixP2eYt
qQffBuBLmj6ULRGbJ9aMHpWbX/jP7LWC962nXjjgW7m/Bx3ZVatvsS4SPeURTfPN
3+Orb72a4P3EvG3dspF54kwH+O+UHyR56BM/5jGQw30Jsd5yz+uKJqUJRsIbl3ZP
jsUpalJszshTcy9+p+I/WL9Piis9R01Fy/f4zu45gKEDI7lHRy/y4cYoeqTxR9Ax
nKos+6xWZ1xB8k2DYQ5fK80epGwBuO8lzWZSMOT4h1Z+if+UnxDhazX/IuvhEEt2
YGWZnNHKNSAtzDIdBfMiwJAOIHuSNnVrzzXayndYqkB1oaRp7umyEH/ayzoTZ3FU
38xbZ0yey8gojqQsM9uk3VibnrojbycAJ6RmC99Kk/HmTGT8f21S8JZlwdZic/ac
ix5e+zz3NrSVEbTw4cm2LJo1OHAtGrVwkKxBBR2bjs6V8KHkJgyTCjo7jh6DxeM9
FEm1YhtIrjLNVpcTRC0KDA8PPnQrz8ec/TzdMloqx+AfMBqFn4x3XBUF6qqofg9u
d6jwkAy7fiZW+HhZMhkjDtxMa+xSBUUr0QKs2/vF/yVBkwOpAJKL10i/+chDXvV3
ZlGddBt/Pm3cqZDLXZzwANc/rk3hUa2aVxJTKKmVRdTVCcMVmYSva9foE+u+6hde
3QHJZ3ZvkfejmqUJsln20qYstBEk7sm+EvUPW3y3GpB368M+26eGbalEr2RXss1a
FSUsOD7OBbJFkkQ+uhYFzMlIQWqIw+UT/61+jyRTOLcECt9Own53dH3JoCcDc3ZE
ssb5e3mWptskS2d8YpGCTm/ZJPA/x9eWgRAQI5AV3dl46dRJSF2PaCubbaKiab7N
PW8Bea0qyVZmag4ET/M5nRuFPMnyrUSLl6OG55M0JQwd1XIheg4WUMFTxbbJQdID
KAGwrTg9Jq1pIBWPLN1jjSY2oNepYmyzFlreh1LYtKNgZFZMrdQnwnoW/zHuHcy2
v7awr2TF+bZrPwH59tSQ041JQrGyoAy+ReLySZvbz5L33SiWjv4+Q6MGiGXOJFmL
YCBNpjKAXKGvfiU5ZpgVwIHI83DKDB/quEhNSK7oMb2i1F0MslhIHi7WwpvXsYKL
J6CmMcu2VZzrJDN348Jw5bwrYdP/5BBvhhQwC0Wmz4K+aVhvkF9Tynp1A9IVQpAK
whM0xcrPVl7XMe5t2BPz6A/cqPqMDySFOP91i2GqN08EbJ86t1hieFPdZzN/qlyn
685XhRtjSUw3DjIDfzohDyZuSZLse48X6B5mkfbiM7M5jUh7nZsSxPXjWmLs4Koo
AzvOrLaa7N5jWfUx8G3lQKM9/1+NhfL1bXVl5SCOiQZOz7mQhN7EyupsCejwBmSx
GWKdaIAuvX/dvdMQCC1rHSRtvzu4sMJ7Ar359D3PLBD2DGagqyl20dKYO1yFtj5T
g8TAPKbe4NIq7sGEefo+Oh8DM8//V58sBuiPDX/x1c4bcUW+e+k5Dq0QAMdOyg59
cBtNq8WVGuxgAlzqLf5IRQ4Kqmp01yW4URRbtoQJGEdv8oTFTfZ1OxWQWShGCtGY
65HrA4cgq9Qq+h5jnaoh7LE+g0GEfcJejbURmhVDwPZlLeC1Wzn0a6E9hyq9OqhN
W2h6SvjKwaSkTgxa0SNnMr4FDuxjFEDrSAkHXZV0KeD3DQI/Nyuw0T8FkcGCrBte
b5RPgTROtowiKSPcUA3pwJNSRzQD93cAmuo4DLqQzxMcXYT9BzdzlixFMJyU6aZv
7USZyCDgh0sntt2bbSxc/WW/3FHM5vHmI4sQfeWyuKOFB5sp08tpTyurmKmGZo/d
F2d3zdHBHJI4rbVdpGz+aU2dZt4BgilT8oi5mw1CGd9c5fwXFzzOQ2y6Rlm3auD6
SRs8LEFbVYaBkrySNYhiEmuOiF8+UK8hXyH9JUSiOXxETUzHOKJmcHEl/sYeMRSU
rJmTnvIJ6Vx+e2mBXM3BXV8T03iCkX0HJtovRreEJ8j8Qb3WufrtEf6bbAoQJWU5
lnwyLojoEt5vZMw1wLA4/UCvJiPoHJnxrkj9swX13OZBVXTTUyJs4S1FnnexDaXm
lro9b6dBt87YYHLbxfv+SdLUb5GdkNvxrcT+qv97JNX55wXUGfR1/OejgG9eb6NH
w0ixWWwGpaExCDsaT90EZjLdK8Ps8GtnZF9ZhJORgdinKG4RTuwhvNabQOPZe5uJ
ondhP5GLSWgohNkddcklp5dbZd0Bh5I9PaNTn2c1H2tfvYPNU0UP8NmjXNEbKtTh
A60im49KHrkkG1W4coiTWwJQS04x26lX5c/Inmn+/nYN3g2v9ObSsV+bGxkKtpkl
MChh9FuS6Yg/do1wb8yOnqSXQggbYxNVlhQy+bQ4Ht9kZoKTPEbE19mWEY8EkAsE
VW/UInCgPvuF3ylVlmolFmLC5PVzQi9XKr7zeSPdLmwmSR6xOR4RlsbNnh4Nx/lW
o/dfKRFa0q2EiJR7yRT2lyxnaPmr3etQ8rNenGGWcDK/QwdE3ODvploMtosSpw2H
DTyM9Re6EfFS4VP5uOt3kslWHf8QZY5jeg4DwNKAClVQUxSYc9Of9pIkC+iozu2V
eqhqPrq8p/7oSlkJADo6/jJWR6+t1rCFT/+YqyDfpxeg7ECxrhnmBY0vXOQhz5WL
oD/gXyt7dj4HeKxMJUEN0GGUC8LmjP2uO3K/5bcbaxLD0cV8oGYsQg/bm2M6zBzl
vrePYC0T8+T7/GawYMFGxNB4jQFOpkVUBX8QverB29Ufw7jsimeZesDbVkvHaARw
2X5gNH3Ex0OqrFY+yXKz9WMg2Rz42tm6Ld7rbOa/lS1SxknAVAVCjsftBLJCdC7+
Q7nNiJYyN7ttsA/rIOMg025sou6RoZV0xoygxkr/7fqPirhSN6Y390xJ6otXiK4v
XY4zs0ewAgBXE637A/ywV3KwzRrssmriI36KaxH3+TgG7L/MkjXDW1o3+hVuAqfT
OzSErygSrKVRKUW3Tba/GkxdHOT2vSmjWk3NIwFAObT9ChO7bxB461PQL/UOlsAm
9qGfY4MRLCgQfM3cxDoauwvmi1A4xkG3mk0xUWF0ugsHNakBGsUa713wbAJbcdsm
7Ju433FBjNndWLaUfUU5q7DChYcIXkRtjMvnpv8EAfYSY+psLoQzQD0b2R85qSQQ
X/l357/K+WAdXkl/K7NX1B4WE5Z37rUcSIY3OL8Jpr99sqLBCPsbohtLDqroCTZI
sgREMGXfWn9wP1mEdjqz0CNZRAIhFUfQzkSPsEEI+9p7EdWyWEsTcnGF+FwIE7fu
m8oM7pqRtlm1vsvf91hb33X7W6HHyLceyIb4jxj7BVQ0G4B3w1TD/7h3P3U7THz8
V12ao7OgyngTcgcUUQcGdtyeltZTNPTmAc3S5ZG8WoHlE4Ixc9tSSCIhvdDx4hvk
giG/fnlBIeMWFC5KgkifG00pWqCnu62JBjCSRwOGgRisNUtrJek+ym32IpvzFNjA
/sLwnGrQRN3y/TEwl48ZJrtjTAs+Xptg1qNR5wKdqDIQFcluNl29V7SYx8oTnEN9
brwGRY9SXPM/fYFLCVTtFk2FLBY4nt2mZXyIQjHL0psuXPbf5qKcwVqiHgdChHfI
4yh/4uJ1y3JmKbELmAv0URhdNGdU5GyAwCeyTpCfySi738IHrti4n4aWy0PCIq1g
sAV902r3dqtVxjos2HUnDVBqGMuDcWYb6np+tN+BNctvb6DLjxKVCdZ2npNEuExa
vHBOdLjsggOZLMn5hwodt4ja5rBV4wWonEndDL8stnLZCvvGoYzJ8oKFKLnJWIG7
ExtyQBWEbnulHVhDpzfN0y0pgzyFg1q4VtBjRLHL/L4UKgL/MGVI+kTFZ9PKrBUj
WM5fZNn6HnJ3zOtQzI7SfIYGc9kTKBe5SFC0ZRV09gPCwMbYqb4GGOpmKsTCeJ+B
6PJjdSWa0v9tvDdMEHxBNVKOQPlEZC+PvCJ3Di7aac/hj02N3K1YK9jYP0i7wxnx
S+o6CrkCJfhOlDoIKAvwJYK8EJwajxIJ8TWMPzg056xR73lfhfAabC0W6p+JbVYJ
zrbKjuD+A6R7AU5T72kzUco0yibgu8nWY4k9VbVSxjSgOy+c8M5EgMUE0ckDN3bG
3sJsHW6pJl4xhF2y/6Va3xP1F/Bmk4UQuDNABBObYwvUBQFfsUvMydwJNz3EJGbE
zv1/L5JAWTpZjnEib3k81mXhI1tNc6iTQ0cqgSaHAYPtOpWJQUozJn742oVp8XgP
vuyuA2/EKcJFclIrzIx6yJlqY9E5fEyQR/oyeHv+AW9hDJUEkRHgZdaLPZy4PLDK
toWhMFlcdbAjVt+STkQY2U9hi1nqg4lZns7uIKqBIVcqEXZB8qe18HFxtlO2CfqU
4WmlzGU5cGxBPrJ7N4/BLsj0Seid3r6sc1oxolxb5ruf/+139o0XDhXZmKeBU9fU
kB9HZUZnA+KQD8ySaigaP4Lstj5giLte1oJ54uGuHyUa8bQ6wMDc4NqxwBYszdxt
j0VDxx3IFi5jSOq2uXA6+/Y/8bUh7zx/eZBOUb2+7D/oe0P02NbbTfc8VuAVhue3
iQmaV3lNwvLmGgGjetsrLnNbMaC/Kq5aKGf0J20TPGDQ8CzTrmmwY/zlQA/zqFY8
oRugdUGUSPRYaTNYBHuKjiMmQVmEpclriSZ2hOpx06DsdVslmtARCP5hORr+vwv5
Rwyl1MjDh57xyATv6Ag/0NgjzDTlPhJP7jYiemz6GLGsDI8fM6zgsEd9MSj0PM/C
5meukpefkwmttCdAc6O51cGEJIJPjsdhz1AxLc5vIoq0njw+YWPaIBqTWv5HIl2h
0U/sPQsLD+h4cU6wYBHAZKltg4rmARQyu4rmzgZ8WoPC5FzGzZT+ddH5QmSqs+li
EdtaFiJQiebd9vyobVTiHxpFNuZuNHu/UdZxJCHoYCXbdtTzz9+b3MB4ay7VrbRH
W+LzOnQJfIgDZ1euTLbWYayItXH8gPnBlQ4aYjIqufga0k3VsdxAwaPNJDItvdv/
gLI0f2FxvpjsmN8hz9NOo3jsflCmSxW0T7yFbNPg9vpZGUFUhtehW3Ws4G1IW2+9
t1jovTOxbvAmq7IYyrtzhdo5fofokzlEhDUF7bHKcLvAWbMNf9qZYrhJJ+pU3Huz
gFsFg+I+35N5gLv6CNqtw6brQ7MeCo1MlCa+pK1riSTVQJ2pSRAhDCh8C524qJO6
ifbTpkBDeoRZjjMFVOiuqBspvRVV7c3+HvWPuPuq5bfnF1yUqSS9VaxrYEvAwmNI
q7b/cxS69U/WZN5Ve3raKt0lv+eOG77tOLGSLMS6iGqbWYfF1oFcyojyBlrGkOsg
k493IYno9eXMzUwc3gF09/2ka95cQ05VI0POqnAInLuNleuzvGAnLBh47itbR9dK
3L7YGcEFcTf59zy+/+tLIXJg1Lq2rrCpHVvdElDjd/1vr6bPmXEFNbA1uziNueFx
yGaP1sc+shwZAkmEf/hx6yDMC4kOq4l65lzk6Rh7ql0RfFAiMe5P4KV4SFo2RrbJ
iq7JoEZLz7VQ3sxJM7y41soW5FMLJ0HFIjnvnlfX2SLTaHJrfDP00SAGAc3xQYvk
yaGwQ79+23ME3e8qsm690C/DbCZSunmXZrUPIJzQFn6d/dXf3OU9BD9faRWy5qjH
wK04geRVCSLFuMN4dbIoczlj8tu89Itt1Xlr5LOy8iAIUtZ+OF2YLMkIp0M4d5u7
r4G4d3aNYFf9kjS7Hoodzg9R7mN44RFARdNjFHIzuUB9YpTpPqYTTnAFdSkT3pFB
aTPN2TVrfQBgHL7/ICWvBzTWbJ85n5Zc8lZdIZDocZ8QA2W3JOtt/ZqpQPLicV7X
V0uzqj3zOEC8Sd8twxTtmalnotBOqrSakb96t/U3/A2Vy0FXEzMjoT2KzTfHfcRu
BaN17llgRx7Fh90z7ItEVVM7HLWYFYIlKEibRZz4fZHhG2UZgMi9LJaX34JDoCM8
Vj6T3kgTexsjEJ6wgKWTG56OPZkVPTN4WLt64mSpnmdnBKO2VZCywD9GvVWzTQEF
rkip+dY8MR15oozngue6COJU4U/UPjLX92wO48M6BtR65y/Ldq207mFLdBs0sOPl
IdEzjXJ0dk9mB5nCHjzhssaYf6YWAG2xChyBxHqnk6B+cgakg83IN9Ur3Pj6PXd7
uCi6Qd4hJnnJBGSSz3ThnSvz8SxBU4kjEQ93iq3wD5C3+sem79ETe+zN3IcFNDlC
hO3Q/jNdm35e1bJ23GekKMYAybDAsV1TOVy1qyEQCHLKSQZad6eAK7Z6BI652vtM
mL8OfLu+JTtNNJ8oVx7ddUaoveH5EvDuGZOZzez5E9XIA6YzW/dqwxx0HGNZF/QJ
P65Azw0YdJ4HSCYuxiBXJjGXzE2PnBMuGDZsZ9OflP7yKwajmj8Fw/iP1/nPye4J
UNN0CL3z7EIhB8esA2Smngcd4saE0rLyRscnx2gIKww6YSHDPPbfD98jwhJD02UD
CtHVf4DA+m8VEWBMk2rdXorIwqYxYYj8keXmyNaPZzBX6iZBONBxxU0lO8KrtImw
p/kDsb2vzWK+SrfNeuzCDWDaN1JNadbyP5IVpDZx+YAod8V6yUW7d8n/+hzFHyVp
L/lG4i5Cp2PrUIzH9wqx3dVWGMOmTGDHMvL+u0VfklRci20AYHoALZfDhIipHJLj
wmavm8ClcnCtf2NZjXXmhbhrry9CNPZjT2RJ07TchWs3yIlxots3MI2K97l3g36R
Ut9i93twFbc1FhgT16XX29NmyFjY+054ed2Bf/2vxcOR6CroxxkhZvyTbh5VvzDg
hl26K2sDQe0z6bggvwhK06G2TTqEXvObZsP+VrExCAjGMTtGP8I3EtMuaJJxQagZ
4SMOL1gn/ZQPmJpLH1D5MGOXoV2efW5s9krIubv58a7tGXvq2dFSocnAMWjAyL7s
ve2K8ySFR0kKcyIc0bvDNjW/MRlwGd0KrizzyWUAEPBB1gTzsIrBNn/cFNSUfOY9
92pSa5hWWykVmyIKro4rXpZXXktF58laJDEsToqvAW0Tiz5LMALhrnpFaZiUmMV/
nws8fqFoZprEMH2+3llDFmgLiFOVPmR3kWoxh/NclqwQlxfFD+6+oqHyMh9Ju5jM
mLM7+iwipToEjHu0bSR/QPjuC/P0LpdzE3smVSPNzboy188Nig12CRAeuBoUr7C5
+dq4rJxqYoaWeAKWQJeVdhYbZrxVXKZzfI3f+vZtZdfNI3eqF+rdRNqKXV5WNRk8
ZFAsmmsGZjteac/BqxhkvZFhWG+ZjS2LrZSgsHv/MDiFtHGr/4gf+klTp0igzX2j
0uQQvktw2ytH2LZoQOAKLeJzhwYUbyhqzJVaducjtz7ADB0zFsz2HqwzPeoZ3PgL
s79U+sILxICOnJWsBeM82gtbE+1n/I4zYMAczGQ11z/YhjSRQnSpeGE8MD6/8o+z
SP8gQZQDtfGqRnrzB1Zq21g27eKmswl/aS4QjXDgREzxM36p3wRMIFyKxcnPxsGR
UTwhHqQVigUTjx/Dd2Z36sC5ESgnwpLF/AtmlDYEF7891kj3+ygGbULM2JSh4mC0
y1Pe30QzYejuks0dD1e92lw/z7IJk9P2kwm9iZ/CcNtRihYvbaL7z4KdboMw5QT2
7qk96X+nipUAObHgPOswYWLOxEFD4k7MMhRu2VIFjhJWVXhp9Lu87EGYMpnh2iO8
HL9paWtoP+IkQE1sEnLi5mgq2gxeUSFF6dlkt9tacR3U0qoBjWN2BoTgmTHrA9IU
A5my58t+Ek5c4vFDxImO6iGXlkCGv13ybcjt4RGk/gjRzKmQlqvdFGXxsYPKrENc
EIRmN8ShE/YZVGKFw36FC855CMMtQGfAEbYTMxxfC7Ynmfn65kGfkgaXENCSDtXr
DYb2smvg8FQg2dL/ObOkcNS2OrsHXQk6UhyUg4f1fhZ8SCA0lg99Z9YVwvO+PgzT
hS7XtsSVj+jFh42/+AayNS8mWV51oIo4tHwfwQAx4V4Cf1XWTIooxkssCLcKjyd1
zqPbTMajhri9pwTGlUjWkDZCTnPT/MSnIqHTlEfBICdGn9RMoTS87JKi/DOuLrH3
Xc7OmzMemcjPfLsJRGUPTFEiMuzgD93wO7ICCTMNSdxLTbaf4keYGKlmyCSGKY5h
ZPncyNf7H4B1PWcBkMoV8DKB24R+eo57Dy99J5km9oIfgPiLT22uDLrIDoSElV0z
5I1bloLLpXri19WhjCkZ9mcYDbQ4LZ1wtZkHyakWnV8TFrC1XrVAdzIsdAUow8Fi
1pXbltq3yTyxXEE+xVJpeuNh2Q+essuscVBGH6OLsFmtwIBHHEqS9DVfVBnKaVyh
62Rvhgy/PdAyn8PjFLG8vViwytCKOuYDMySLjRxr5jWB8JbPmqusUGdZe/n9U1zd
qqpgIXXMZiPYJwolLZqYtdWaC5qA/fTd2yKAnVZWMXckVoejZfeyBzTfa/GPO4Cu
f+XIT+nkrtKK7bVBlLwzZ7sHR0/nynfQUl41Co62RWc+IE90TQjG6BozpuZS1hLL
vB7QeJAq2QNSRd2GhGZ7i06OhR5JzM+lIho61XPE/Y4u0TMax4joMlRwbqPPNnnd
1+9RSN/yqgamivC0VBg2+Z6iRpli57LxT/76C2OyeCyZaNJeWmEE0aFBcR4BsnfD
xwAAwTnkwEkyx+5GCV2b6J9IuqgDjug2axgy0z436RZxGSt4xe/ZDRiLzJz5tRXT
9BNFBSNWYJbMUK7ZiGgySlG8AlIS/Bh1rT9GE35WDjIkc1/CVBf+VJJ9igJuKXvR
w+YFdwcxiLMPrmMUpWazjus9me36EPUb6gEvAFkozFVh4LW8q3VMLxNjMXZuSHZF
91p/ZzY1/a/AEjaQKk9t+wMt4jpWE2QXfoUmiJl3cEwiyNZy9C2qVfqv2+VWF/l8
QwNaO7cjhU66PHlfy1ZLzMUZtImSk8clcWlezh4CYX79bkjRw3CrLByB6s8cAiSm
wZ0ezr0D16mc8gzGm5vN1rdFANQ7TQNPfFiJe1zQci3BfFlnursNS4C0BO7rebLF
Y0Nez36jujw53OkG1o+vQhOMkeNMFuFRofg8qVTt6WVjeW1BHlSwQEUOmmtMdips
MKFE8taxmu/WqgvdHH17wtCa7TjM23wUNC635Mu+3OpauAOBqn+ArcICpJEDb5ew
5s4qzBRrcXBryExxZSCYuedHNJUPt4Qy5yLhga5/AdLRlHPDRXXlDnYaKySck9Hb
INoGBC+Y8X/kqMjrlZIu8OvMKzGrYQtlPQ0jQN6C0R1Ey7wDPMBYT+J9sWn7uAUN
CTGykHvdEoOt5K6417yVxcmYvBeLz9G+ogYjHzij66ghlhjR7O0Ou9bEPCTtH0TH
5aCu5tD5urE6lzJEkniZVo1+RRgZ73ZnsRFCQE/ZnYsg2PDsIzi4kqURWpx1B+wU
HkiX1bpvCGODY+JBl0KOidu62a/u3DYFQ2VyTZd5JsUlKRAdQkpPDHhFVTzhpZCQ
ICuKYmiRipS6ipc4hPN4q64NxeyPEocVzkHUdlrQxi800Zy+IhFieuuxzUosvf0Q
mKrP2JHykwNMcFXzqkgIo8JLBD+KN8Rl1wMH6rg8oKOWdvaSoPKZAk12Dt8WwzyL
vN46V6SRZpg3XJK8Fh/H86fQAWA9BRBQbjt8i90jXeNGYt5Svpmz760wScPe/VjA
Sbe+zCjl8CJDt7J27neWggIlt135snjdlIvQ417iak8ZRCymvli9wuiuk9R10oEi
o7P+g46nosricTyP/3b9/AryGnHa2n8v/snVDOC/ukRAehS0YEL1kttLp5F3Pu9X
i3TIpOWz7K4F9k/bre/FQVWt7PI09cbEI+bWQmjJL9fuiANYK5dYAruIaRhXBvbv
DbhvonQa6EHf69PeCbCuUGgVSvP7JOM0F0NCG7n97yaiI6xl7oOeLbPSye1EDjpd
1JZOOGcw2+fmtqAhEtwM/oqZv34xc5pwPlCgwVMuB38PpD4HIhS7XwMJFO5+tIiz
bKu8BD8e+aAnEqwHdCSlEWGt1zMRTItzLCjsgXRyYRV7RwyAhRBEC5596Y5qN6Ar
+AniSx3wwE9dtqWCP9YAEMccB9vWOeny/z6hsXnrwJcI78Qal0jgY1Hxkf25gVV1
miNhrbXIsxmpXafbDFZ6RBq/XMV6afEHq8sGcQJ0M9SIYa0MEVv/QjKr6GYDuak1
lkVzmOPKwuv3gmecb1A2/g6LOibsqB9OeBXZeGEIrWFNOd7XY/9VXvUG6R4Nap63
01sxfjYKy9tlg+SVbShvyVHWF4QraEenPxF7QgdDk08Nmw9Ke0rtlcvUcNzkOwQ9
ZboY0E9ikr/+2cP5JJEVvqIUpFxU0xZG6JvWjCdm/oEpocMS7jTXCfUNsTf9M4Q7
S4mCsUChT/h4bvfgn7VSOvorkSrzihRNBybOLMTJI+N7K1D2IeKt21UPosr5jhq8
2GnseIC+zWzsVQ/k49MlvyJQHmiO5oBQPcAhe1DL8Y0ZdQmIfIf5Uwnfbsi4Pbip
U0d7xZFFdAfszMZEbd8WEb3sQjv+/A9+wMszHbbgcUUDiwH2gN8F1iGEA320uDim
IB6JYiXuY3Z4MV1uwHXAqZ64KZZC9032FguXUv2JYdZqvMqd30bdhkIWI2QqGxXr
Ly+tUVL6ZCxkTWCJ2H9LKtokixWzX4YX1NeGD2OzVy0ybPc2r6z+LOcgvE8IUGFq
V8alW+U7fLGEOSx9jizhUZTuds56NcMaFGZT9+OZfiAq0UjaSTc5tEyy4hin61ax
xdHYLgyEvu7agmchsycfaKUa6yRzjLutsMsGc819VstNZZM8K6gDGL7YoEHh5WdZ
J/a4X27IpmV9AOvpheTempGRDDlaRpTxBgB7Bap3K7CL2poVJrBoX1gGG3IfbUC1
g6F/4YIcmzGloRdamLoMqSOK9ZmRE7LoYsUhrvvBDL5UypYTouxlwBL9+tUKl0L/
I2g+V+V6149xeX1DaaFhEuEtOQRx3RUjh5XWChkb+L6dP+uvZhR/FPV7JO5JRmta
gu/0bHgLnjvazhsn1VBlSkL/mXKdQ8UNy87aepNsYqBlkCZVOn22yOIfw84h8tWI
5NSKYoYXl/6wdxAa0B1ftWvtV7AVEJXGj8lEW8ZTc1KaAKfVPKDweBDPbcVey3dz
iqG98g4m/Uf4NOxm9QtNVXfcenzcFPIkzU3SDcm9/Cftn3rZhwX4AbJdbaSUK3/w
Ywd2PoHVD0eg2Ni8W6EwMAIcjZ0MQcuzb9yhEblxU5M0vMdf/FARpXDGy910YPLS
eQVqxWolFXNhjVtGl7AV0QlSP5balI3udcA/6/PCJGssJDIBZAfIHbv7Dvlh0/gL
8bdISiK5qN7UDVgHAI6UIae50dKG8qNH++v/lF1N+7SRhY41XVe4C9N/DmdtvA2w
VFUiaBDSomBus04CGs4knp3j0MUSUqWqsOxdUM0vXJy5GL6TckTM+K9UGh2AkWvF
MAoCcLxQYcFxXNDfqRi/IhmR52ZyiN/1VIyQ4YL932ihkY33btCzMCt7loG18QFj
/uK/lhtSLi/pH7Qb01L10ibD7obx9UVUEtF07B18CxpMp07nOmpfe/M6LjcDR5yn
4YnyYgxLcf9x7Oof5GA1Mw4lji1maw+kDpbTX/QNUIdn9Vus4BBezUD6WfP48f2B
N4lMMW8wMthDeFysOZEt0031JT9zhA4m1Z+RXkyOSy96eKSQEKtF8dguC6oF8EnJ
aj0naQZ/avs12Nmk4IiYsICLDBnpoKgkpHGXoKDV+Eo88jMlgbVwl7bd9sKhBU9X
uNPjgUkOHdA7oYZdYUkp1yb+cwK2fGly2Q+U7z4EnZnHMuOju14+O3UVDaNNrwif
FrbItF8j81N4+g2tDLuagUeJrVAhHo7ebLFcbpG/BVIpwmqoX5ULWXOzBsrDUWuy
ZLKdrPoW5Xcue4lmlgSP08it4242VJSsGctnc37x6vPCLhgWvonSOZWFWHgJBkh9
wAn+0zqD6PbZPZpMqgqCQS3F7m7mqCF3gftHuwgdDpMYL71VCxgJGyF4JOLI+jom
s+AJBaBuyvOK8rTIKaU/qabD25t4v8SkmvfnliyNNraa/c2HdL3JE5DsLx/XW7hJ
xLe7XGHHuX8TiGI0kMQV57LzE5iJQScQ6fFvpTC3hjaOLK+88CNfDjr4HK0JTWWv
OBcaP0clsFc8a/mrQ70DqrzBNopB5YFAQV2+elkhV7j4ZyAR1xcA4xBJYvk+cpIn
X4zDtKEPJPSmO6oGS1C++l97grt4alVIAqS56CLTLo1NhfloVfnHOD/pZMuAVg1q
+o8c8k7XAGkcV03ujjBifFfNe94jMRMmzpocCBckNSXJ4IC78kfOSLgSUfVm1CuI
B/sj0mpwxE2htKCuJPf4G9DB0OrcpD6ysTr4+s14hXmSbSgh7ycUDymCVUaCaAj8
l9iWmIJsFGVb+S4jyVLfyQRqezorFLJQox8YhZCLMQlgxK+1i69ON/8HOquWy3O6
WEXN0is5p2MKgQftNeroC6OfrQmvcZSm7lkx1cZGWn0GrJF3qR1iH3Qhm/aKePlY
otoHaa20Qba4df0o/da2kZhYzse9cfdOFY6j5JUHjGZSHUmH5RW+Hd7PpIbAdf87
5DYQSfYxry86k0DNCV/B7aKAA60nP8SYaU4IhFW6R1z4dG7EgduDGu7l52g2+R8f
8w3VDDKRc1liQyJl/3z096rrzKaFwG/6U8zU3JrqhbyqfCNjFxkriYJNrBsdyHAc
9r3Ymp09XIr4YCfQjRRHwF3XG2ogya7xuo2Lv6Dd+E1032/R0ZKpvpfWT+ulEjEw
rWSRhFZotJUP/qxsPGWf3mwMVDHEyuOi6ch0JYNrE9Rv6XDB3puSBi1/CESkrMeT
jGaRkGiE+eSMdumSiJrNnXLQz1MTad4miNJcbBIdLaPmlS3bl3fd3Qz1O9Cw8YV3
gk4QXmjsX2lidiCeTSh6h8wqIpcjlFHsTknJ688JHl6YM5LSxMCor3AfcSGTj8yW
whV3mONoosN9DI1iRiuDNfij0vDlcJv6Uh0MqJvEvccZLdilBcuq48vkGznMlHUU
rPIpBgfACouX19dcQ5AIB3odNTdEBcAsJJKZOSiI0LrpeB1vdbBxPYQF8fERl9e+
8h6AX2jukfhTD3eJn9uVV+VLpo28Rykxrxv9D5A7R51Gdp5GjNdh35cIeZ2cckOh
NzsPUQ91zaBDlPZMCI+VJjzJ7JtMPo6gZK7NsRPlZXLpx1MqJy9RsMOFXJb2IRrQ
+YKdleZMZrkewTfM0Z5kQveIl+DitQE6q2ypC8pxlTsQ3ArpoBYJDbNH4Lz8kCB4
eATBg3uNeQrquhX4LWPJ2JEvo4bYiz10R1W5dtGEQbwWCgIHRVwDNffn6OapAOjv
+H7xyHAH9Tfwb6nMmAwV6GB7Nbthoj+3vmw7jRnV+8YkzFnXHfBJ87iFSpsvnFFV
gpCtIsJHwtixZ6FcuKm+ydT/4xFUvIdcvHsZ+Fw6eduIIjAqcWDHI4CRSoGK/yxj
Y3yOrHUF1h/f7numOVEq5PeeCLF97jNQEPLl4ORUlHa7A05v5JPOnUa+CFSGh/YY
x7r+jfYFkljKceu+7/O0Fr5jpqMhfgxDaYePtcm3LM6VwIrl5wrpVQITwxxdBYJJ
XLdF63ed+odSGrUQPYa48Sxi95XhOn0u8HCS7NUYdoUweRTDnNj9MjgidXn1UKh/
dgEEPLJZhd2iV+sVzs+YCqRg6aCS0wxH7RYG95y3bylhFFFLxtVNXex6ntSweJYr
wr/aPHMUH0TuiQ3r3XJ+0vjhFMVuPP76yngSgdgX/aGEyOW7a+apHIk7q7hfYSJo
hYIEhfLj32S25YWliUktOQr2JxRB10kLJoqdxWKqYC8/SpJty9+DqMNSVq4oeJxU
4iDTZDJ0zu12S2aPwIKBowN5i+LhXxInJN185IFCOBzyVqWushXGipAo3SpJm/0w
rBiwRnloa808efm8DRJALDPs+DvueCYMAd9eBBp40EGJhij7+yVHyCs/W8UOHLln
O2WZAyIHAnOp3O+VYoORA/pSfZMGueqzTHV5h9Jo6cgkhg+w3P3BB0NvyxL6lOx/
oMBFA1g6roFOB0UwlhZuam6ZveahjcsQEJKPaGOaOCwSHa7lLIr5ki2ScIh2xvUD
A9fn5BXh3QMUNbyPjVc7J4FNE8n2u4tHtKu0uxXQmrsjyfHQ2lrkfYYYD0/0WSh3
au1TZTaIs0ESfprzkZKj1t6n+rKtLKIWklHGTBoMTrz1WtRj0QtNdWb3GLteluJW
SYndbFfZAtClLdbRKCoIMkQXkI3qFKHqXUgrJUI9f556SzGEFKUlq/aId+NQd9nz
haHzpVd/pYU51i4XlhxoyRKVniphG2ukt9UnJ1KKt+RF5CaalUrqZ9m90H93RXnl
pGvFR8ZWmrANeb5DVIfs/pjoyfAjjGJyO+cTxvh1ZZ3FZeQKy/qE4w1BMEePFYVR
DpufJBigy5SJFNDci4CfYdpBo51MmqwQl0+1D4AAG0GdsQUc3Il9W/l0b4h4MXdl
vTKSUKyiaww0nzu7wPkbYGy1Uvzca/r/2++jv81rljlVC7OURRGJnKDNBMzjlUeH
/UWI344CnMdaw3E/xsheK9k9T0K4nFcJ/J9NVps7OdBWDcltErQclhqun4ZEoURm
iKhaNVECLz2WCrzkpc50UHS6BwkSnw44wFGsAdaojOAxKZ2rm2kREKb6icL8D4iC
/OVAU4S4OT1kAukCppF8aFScitDeEdKUuf1NQgRlVgHO+6f+3SKJ7eh9jcb4mt5i
UB1sDPPr7u2wk/3uWcA42mHOsshpIIVxYq3GU/Bv+/5s+mtnmRQ5nCaoEHdVxSJH
hU4qIE4ajoHgveXXr+7g8YrFz9gE9LY3tn3k8SZK44C0ags994AQbS3igTY2wTpI
Snz7Fwkz839g0nnSfMGc1yZgqlgz6ICO0H4tTJ/zxxJ9Qm45WH2TPqD6Qn3oWQUc
2fE9APlNZm93PK5ks08sb9Wl/Z79ktbPJjD9XfY9jajaWpIF61lbm0LmszlN6Dss
JbcA2kqB8VvMNsJLGaP08ncSCDIKnHD+PwFpKztb3sfeSF5MpyVPPZMQT8k4Bv33
wNX/oGEEICSHSgyeDwytuw2s1CfpTwywoCKjZC6+uNdzvmA/0d133DmcvP1SPU78
dvfDQXYl7c9EAyizJgJMuSGq/fWDH+cOTYS4IzcfRz8EgVpfVXFRNMNAd7ORmjsU
pCL7yq7YOlEdBzmT1qu8qo0qcZ8srj1wK/SxaMpULGQzWbwdYmHus2ecoC9Nz1Nk
X1hWSKq1phiSZd229U4HIQybNKu+q+6Indoub5fnN/BdbEJcoFfJ0M2hQusYYttR
P/v9TlbQZt615W2vBH2CqnDw3mB9EQlDqvhza2Dhyw4Kya8glWefcHhOkr8382rl
90LHfz76BrqsMurAt6sYT3df8nV7bNK0usyqWNL8KwZ+mIKylMzRCk8T4ZZHtj3M
zgADjR11vpdhF9WKSj/mK73RSaZ8gdn4g+3iwz/qEX+BjjWGudWAywdZJX3dUvtm
dN0XzdVCtmQ4ZCyPdhuW9lZFK4ic+YA0oQI3x1UNlM1XBwQGzxJ/VyLjY4s1YEeC
ijwXdtAh34LQMLS7+VhD7mTL9cq4F3vAJSZS9J8YWF6Vhyab+XJjsyMh6g5oJBvx
YM5RuqtB9a1aDXZrt0gxreqJaTpz5An2W9DGsTgIPNvss0QDd0lyrEAuLATQm6LX
Yh2J8NJB9S+z/gRbQSWElxUbFAmR/P5/2wv/zVKf20pZ0VMXdwRcUp8lIWPruDzD
8ACoHtRDmt0maSLlyAsbLmSht7+ggGo2pXwINpj2knH2XMqJUXo2c/hoQ+3T6ViZ
qBm+QTcn/KSjr/bdlu15Ml0VgXVolEb2PEw67tsGrxcoZVkEEZLlKEvTMRbFcD2v
r6mY0VjOBoRfF+3BeRay+DvVkml8P8clliAgTaYehhO8RCHCFDuUnUaHF0S1K4Kp
UKz3QIsQsoZOrwu44+Y2bz/+Mepv4Amdnt+uKIpmKGPxQmDIpGodYlb/8Btha1BW
cmhaXaOcRSVxtxxxmQxxVZSshHC6Mss5RalhBMJF7illUGRELCsu3IVCDszEi3j3
/ObIMR0Q9IFd4R+57gx+TKN9kHrunSDZhH2zkG2zIdX7LYjwQXuX4p6xk2/4iFHG
/c7wOupOoN4XxtsdRSZYTkyPP2Ocg7/N2gDBRBJZuqovc3Qnd2gz35rN25iaSpry
yWerBEiYszGWHg14lqMFXdxqqeEIwP1zW44Y0QtO/OXTrrSNexDAsfamgtmDof3w
mDKkgunHBRv4NpI7SHf/0+g+q/n9WQVGPGIUvSlpZnWv4VvGb6fWYTcw7kNRxLCh
KxAFJX2KbSuB8AhQqJG/w9eeXgNDVDnpN+XXxKPFm4IDEV1StMvHXm7Or+h2kPfa
9d0q4Ej8ydijBk9+Xly1UJfbWJfRmAF/BFAZYe8Pko2jTdfgAI7RFxE0huRecAge
cPTBmjmzaX4joRAHQjKAEtUtnGG5ttWERbyXC9BtS6PY25lqwqETVy76MmsLNTQf
sJ+3l8T7mt/u0RbF+N3kuxO9eRLsE+4BYwEwN9HXAaa4TtUXpw+L3fNhZIkeYy53
SQOKbZQoXYYfkE7UkEoyKLW7PCtZel0sl3shUdTQnvPDWkR6MhTEpqr4pY3LKMC3
kwmsFz9t6WS8VDp6Sd5yapVJua8VneM97Sp8hReWX8lCEjDgk82TwFFBw1jo/nh/
yrTjGRSTgAtCcQLFC5/NanZEJ1SwqJqFvAQGDEtJp6dw4rD6Vi/2oyEo0KhmwOw4
aXEIHZOozrsJWAMXx51giYP40VtLHvqZZfbyetcCO0busleRjw67+9T88/eiX/CZ
v1fJw3Yn1NVkOeCJyf6PUanEyNKtxV91U4Lyy9Tp2STVd//hKha68dxmofG3azz1
pzK4XGvYVrEDOAqp1vfsH/fWnEWk3Gh06mUsZCFONP1sUO1am44SlFQJ2G50BVoF
ZI3E//J7sla325J6TA/S6DRVgWoTk7RDhF1JcoU3jlreMLj5YQMjPAXIOjRlz8KL
/ydCWErZXfgSIIaGfWS33nNH2ctXFkzT7LCGl3KjR/a3dvlrHD0b1V+Q+lzqlbSa
secA8aUK4ageBG0PPMA3J4d8PHpOP0zK796wLLoHqpRt89eDEG34aeTv2FLG9++Q
9FnKKguct4tUhDX8I5ONVyUTp7ncF1pr344E7dl83fBKXhGtIWk8cnbQzWOMM5fp
krHls9pj6wKEZzsGBwlvEX/1jiS7kmsgTw3SiF6pFORi1fE/aAvLf9DPEFDSTMlE
G1QCR+bu/84u858DTOmxg1lshrjzPE0marl+C1W7QcXzDv7OEGlSVKwaf+b/xUld
16c6uURY1we4djEFUKGj3FJ2D0zxH/kAV1x47iRI3J4znvz3UkWAI3wmNVK5cr0Q
5Jmr1YQ3iNeDo/TfoQ2hpRWovfvQCxkS1qsVaq4eOUrKPeI3mJOQ87uLpyPndQhm
z5netYPPPtqKvlBng/m6Xa0bJxgvy+JfXE9WsflWjd1iZjOWK61dHmnEr1i9Dq31
ueNw1hdWK2D3OMUqSlIl8T3CeoKv1U3dxPCnDVO4TvdkTboQp/nrMXYpuM8MId2t
2tSRfteq4kBzA5Rntw3XXuhZju7y27gLDwh81DI3jpdrBOY2RF55gBzmnrN7Yk8K
NPwUbsCIEURiS5ObFPDstTVrPmUPQSFU6qtzFoQdpWEoDmqqWHv+nQjmjWQF9MqB
FRk6Eju239tdPcK9WJKdlXRqG79Q93CRdU3aWMqliDfwZE6GxKxfK86gJ5oMxmbr
7YBVIBbfyZKz95u8//nrO8VT4N9fh7TCDON53PKQHrwbb1i3Wth+C4NpHaMrFXSr
tWusHD8qnNhYKM2tY5svCVA85dGGSwzESAdsLA+K8HMwDljnTkl4xQqzGiy670AM
YrYprc7Lmtk1Q9XEhHcWtZtjuM+HXp4fi7/ko7pxa5edVQm9Ftid8hjh1orfYKyz
3pmEVnRhK/TzObuwmqtjWHU4dFgukzHQsp9teyDEC4+Nl0fewU2JCLhaTQyLiwaD
nt0cg15dSzS9lec1/Pph1cEKaiOzH9D+fxYU+gLLd+vzG+pRyDHeU9hNrpvLZNuI
1KsowzoTqRLMwCi0xHTICLFfbSEKeBKXLQKbVlXB9OYjnBcBTEP4ovX8/5wpdoDX
cDCz1ESeVdApSoP3Gdcv7C6Eoaqvh8v4QPoqb7bjX5VzWuGJ9Zp1nIToRnVEp495
c9RSZQ4Whq3vbfV4MyprWzsmqqn+xHZTbTxl2FvlEpUIu3J7wHZe1Z1mP2KE6FPc
sKiYadSDxmKdslGe2e3cREv0I0fsP5YvaWv2Xvu7ws4zYjJJr3iiY1jqimGoANHC
gUFHHNJU2yINj0OrvX6pfu4wv3UF2o7SrPLtWUHEj7tq7RB31fkT6PN1cUhmJ15L
MaPAyo7rPloXdDntjEUEy/ercnnUHlWFn7VPl6wj2Os2OX8AH1+X3syd7fmvzlDo
/EdnkMSV8y+Fl8N6XV7b4uGvjyPnzkSHnYY0H2YHinqnv6NpU33Wv4clCZuLEGbo
LplxRdAnF3qwXjV9PI3/QGheq9KHD7ajBb968l1QlaM8ZDlQJKvwxbUPEHiGxBLE
HUJihaza86mJR82t9WaKqCV1ZZzHpgCTXi4VJu5lYQGmKcC6Y9d3quYfvdQWFTs8
O4HTurcGWWU4bvpmmFnLCOXyIxJq1ZRd7S8VAoXw7dSd+Qe/PVYkRf/Js0hQJKVd
1et2S0r/vY3yVZ5R8hKkWTq+4lc9QEfYUp+BdtraiHFB4BZQOM8B1d6VlrZuzrho
aEzpw4H3YBJaSapzqLbHXgnVULqGf4qX0GNpx+tL0DEIMACixt1bEeauNDHUWayO
x0serL7cBuArO/wZDHQBXu4pLqqlpZu69bv+EJUGwuLED2vWOPMgoqDakk69UX8/
cJE537S6LHZgdFqR9VwM5oYzbkocU94ycSiKkaftXuEs/HmC28xEsHt699QTDkuW
Uow/fkNpV1bOm73kI0lY4IJrPjujrH55CTG9CDG1ts5sq9zA9GwPiHm/x7JiVuo4
GokjezxQL1xVrvp8NRbJdwYXUUTQ2/BVCiy65+Um0uL5T4nnSRfV7dubutWVEc4Z
O0vpE3r/JLYiBTA67+CnUEUg2pPF9yHP/8z7gOIe4j2tWtKGttl6Re4wft5XnHXF
BLKB6uNS8a/sPjMM3WCEGYBhZoOsfBIbb9uo1ZvqtUJ14ndevCMuSznyS8XyYSal
WCSBpnpZgSvid1hWCO4Rgemn2F705l8DuFdWjKnp+QGMH90Cyy75a5kKz+pa/uaQ
jYmXDnugBTw+FrQYg98kh1+KGgg7iRwr+gAiHCQy6vYSTkpBDjc1QIzkCCKrK2ZV
FoR7Lg7nGbawBkvh6mc6QkAQTdpMKJHLBEIjB1hfsYpsyNR3lldj0GtwTWG0IHsV
So5ICLgpEFRd4Wpt2+yk85bUlEhVvtcEm+ZvajBgHnEI46MWr1kj0X+64zN9Zm5b
Zw/fDFaVC6+tsHCmtMkUNwiJGrcE6dVk1vOuOjYQIJZ6If/HkrnSJs7ppmJdyENV
ivsr1Y2uhKviafVvXhmRAwrjcKHnn60WeEeWsN/8Sp0mSuBygb8wIoZHQpTPxuZP
cd5AdPMxnhydOCfNOO5dlq9SOmGQlWXomTdqdnRqGBKN+Js17yRagw5/yEOpmkyL
QWlg7bM6OHhEkiUPfyKKlYJH8ceWAvcC5V6VKS1EcqqEaUNBIjwmmYEg3j7Te/vv
xqE3JdJgZe58FMUq8e5+BpH3CEiig7aIviMcq+NeXpmSDkOqATJfosEDjjYsU5Xz
Nk6Yhq/s5ahHy6qSfGKc2dqHPO9DwQxnPlmcqIzeLkrI7tlUf4YwKVomqEGoi+Uf
RAP9kKyQyw0asCTZPJlya0wKrJs2iSCFSmq/ErREfacizxKIWVWJMC5MspLLQmMV
JXO39ikZuAsyesXd3r6k54jmX/Tp2Fl44lcvf80U3Q/wu0iFk34broPm5P56kKkr
igQVDEl8sdHAgRxRp3tXE2dj1jNquNuvu8/++6Gf55E59JDgqUJu89zTk4IzQIqK
lYlj7JkIVuua+x4BdtJq2+b7Wh6zgu+vTmsiQk7AO9tNNA66ZEsU7xmqCSgAcYgx
28FydjEKH/iyZckx/eQ3KL5KrvDgqYHHMppW6GAQtg9UWkb7daOCdVrHAJ3D0p0B
x/9nl4T5qf7OnW9gtHOw3ISCcRoSMM0S9dRwMDDMPzftW9oITivcTAzJ4xV8sPSl
Dsm+9MV+itGr5sozIRrp1YSjx+eR4amik0/Zxy7Nap8ol3rAVGhu6xgkEVjJeMFI
A+SmP4GepJLClFo9kOiPBk/tLqDb5ZcbB63nkODfsnCjHJ28/Cfa0SnUNZy/VEkc
pQY1Qp57em2WO3Bd/c93OcRB0UCOTZo37A/iEGv45zYl3YLpqybrpIysuUj6qe3l
Q1eglAoJ5AQBNQNe/k8of/n1k+rXkF6tBQFWFv/r1qooNdsFkS+sxgVJkythMz2L
M8kdqSf+skxINErGhvvsdjA6vVoJh2PGZ8lMrrGgFMW08Zsr+8qNHl1qITHBEf/D
JWAbhBdzvAx31kdTGc5Y2wRGMb8eOObfNyX0uBrpjY+yQNjOcKIpmGZyP8SCG5aM
l2YB45mwMM6PI2mYgJJ9+ssrpbR69Gv1dsjP7PAee1YiTJAC65fysSDfmHh0/5Gw
tlPjhJ/RXW5F8sevmCYQZMkdigURGd0zY6YpUfNW8fnvC1KN24/tGd3EloEXwBa4
uXqDkOyMXQhqbVKkMCNur5L3OsD7BqiOIlcwpgQwd6vFLsSt1qezsaR1uIgOKKbt
Iw7RcBdneSsirj8abUJWeTzyK2AQTIYDRrPv6I0pUJIGP0McYabEb7Cz4DSVrV9z
fbqS5lCTPP1bYPLmfO2DMBvS8hzX+SuifUo5Rl7GE49YJGjeA7q+9KeO3rukrdLG
+BDMe9jav58/PeUkgHTTS+zCqb0Rv/xD0p4PWP612hZA9YLCvgdiZb9WPGYu8Uvq
k/ksa9XNZi8L8bR7+bS623agG2pbZlMOsdbdQ6pkVluTmDHIFQednh1FcTBelCwe
E54j/IiKhO1ifiiDFYrIiT2nQ70X/QSdp1/9PDH4TngvdCGS+5y9zfVVQXRZ6MMf
OGXUXrzPQ09DXVfxJz7U/3qdUe9O/n2OrQ0238doIvMnXaqkTe0AC7a2mrqepFbp
QhBX3Mq+kKb1W/dyBE4NZjDaMK9bTzSEMEBjZqfpfRKe+8vI6nqG6QYnGC6jjAZa
+XqB97BIedXZ3nEnU/b+nwFjXRAtuO8juokXkwmGS5aGvXZhwaw+yUvvC+we5G9x
7vFLUyHc8Bp8U1jNbyS2KBJos6HnsloWct0czrNt1PHG0am4Q2kspsh51e+Q8bLw
KqrTarb84mZGnfZm2wdOBkrRdYwoA6daIT7S6mUdVwoTttmfuS0Or6ZGguGEruHr
mOeajmE2OUzdrjcI6fCPCD930R+6fAFFvSU74u7phuL4J3JA62/Ls2myIPyCLKwL
DTrDMQxqfRa3TuDwzptqaTuHX/cvuSe6G1Nq/VMgXPFS5uc8detDJtFpkuCN2XBF
+ySEiKnHnJ2lRxMKOghHASlJoexk7quNywltQgpR198AHHMEreM6yPsqsWy4Xz/n
e0VEHrFsLVJFW4WSIWwD41ZyNd2GGPRFuJgX9qtv/RWb/ZYLU3aofC3KE6d7x0nT
p57YEZRiWhbTZEph5vId6C4/pt+bdAOln0rmGnX1PbeFJmZ/TOdoIiIyEQLEgkd2
2O6HxNXGuBBnX1bcp40D9cHHKaXlzlUFA0HQ8UIJrW+SCVXtq6i+X4PpwtWk5axM
TdRL2MB6a0cRQ28QTsgIWTTeZ+oENMx74A6flb4DVKDuVGJ/ld3maGZjZKqF0b7p
C/gqAFB73sgsBEYaq9e+IoGXJRGvXZm+Gl9/CjEcP+QNwp37pquZRXTZfpB2Xyhv
7wLwWD2jN4AF/wlseiXUlXbwssiewlnYQapoMFnXfX3cooIx4r4n/L42FRgMz/xR
QAazttJ1VHfotZXwGUe/fCW9qnSWpMJmnxO6lpMDkSkJLqxGf4N+01sEMbn1LMoK
OFI7guY4F/Uz94O5VG5iM0kdotTa9sVDkmODbahotZa2Ob60PWcJKCFGcI+nIzD1
qOUdL7GBPHnRHKCaXDZsgOHg5X33PfEUJ+dCrBRiymEHae95zeDbHV8d/Sj/kqhe
CSxkkBPk2vH39jirTTGNeIENdYqWJT4aXCKL1VWYvcwBUgViJQALX9lHWwzMrUjm
yRXUpnQv4JWv8AmCKyFZXUXz5rXN7gy0yzrg7r57H1nIU5la6refLIS/7VaktLP9
evdWw62qazZyYH+CAkYvF2jjeJAn5T8hnmd1SKL71t9rObGvBVj3mi7aMDThZecx
6/IWMxY9Uchqn6xU8WkWg/zuINfX6yugNj+8K4KUvoezuPyno4dvKoY9DIiEQLBq
I1FRrrJCDBnADRm8a7pnZFvO8q0xXJxGjrRvTO9f9QN09F18M3/pAvpBhsnz7gBs
deTe2A/0YJk2FE8DAikRmzfXkqFTwoKxEBnTmalMQnUt+TtJFn+BCWW7Zl57hDc6
vfA2kLt/WULG3QNW81QhdASzrwYWp4mqktyFGNSktCzSVA/7C1OWn5WFwO9xYMoH
Tb3OreqTRGygal2sOVNOmcXHD0w+iz+eH36YetgVzBVX9PqVXr+hezsvUhmKmTrM
BlC7xfsB6UUT0IbqRqSQp+zEGQ0MXG84gBZ59OGqJ4WJ6horTyNWBCljvajR6Pai
xXIerNsYnUTojpAYguxpi+iqQaHd/2CSoeWTdAFLWPqS+AeyxMoZsOMcOzm1Aild
/VUxut0Qco3OWxR+utc6f9Qkke1wmhSZIR/w1pFjslwmt/lw0xVdYvUWZv8qwb0t
klDD9Pq2ITMIWcaBpCpdFT0aho4lo87YT4ltWwF1MHtnaHzNu+mVChTVqo0HcDTg
5wmJat0H4By3SxwjL5jQSfK6j/epcri05wjObSiyVR3ojY/4x0fbeE5+qiG6cirX
A+ULoM/1B18bX92bL8aXu7CfHj/67m/wad2AGl11UtxXek1j8Dy6Nlc4SuZmXQNs
Y81xutdtG4JZDO84cHw6kiaB2UwWKdRQFhpvHgb8ZI2k0m0z2E8VunKIgsmSTJMn
5kxeNyrfVldxF94DU0km5hK6rjEwvV8eNnEX1qwIqxjAyDyuDbt4lqDEOqzTc4og
orhxpjZa3C+inWwR5tgPTOs2k6s7E6qZBQXff5viRqXcDiwb4Csa92zT108We5KO
qgs5eoOGBAoOHGCkur6Vvn0EOw3fkrvnGme3coDEE6MFJ31gvgNvE4gewDHVBWLt
O4bMS2kkL7sgR/WJlH/4XRdatwG9tDsYeLcv5s7qA5mIY0p08tw+u8bPHPUmRLnT
X5Skd1rP2BoyGo8mf7uxFf1Cy1Js62U6MqiSMm8jGxjAgRqOzZQbiUdRRhUvih1r
5E4XKT+frAzc35QRVtBdBt3cHWt2UUaLp3BrlmWOvldpXxyaC9pF3rdaRVPBXrMv
8MIjHmLeo5o3YZHVPo9Hyphxe/LEeVXoucK3TjbYp0HhVJmU/oN8ldHcJ1hq8nbK
f9Jit+polL8uzFIm3rm9ubIlTAAS5Rqisi8pIcBPX5YZq28JqBttfB3s4ikuyeRW
+Uza/to2AJdGUAMjfXAGJK58qiSp0F2IJ2UcJ9qvQfpr1ebYszePOGD67tcrGXec
Ao9ZOMb2g23049cuYBh1rVyEwGEc23EWtKeNksN1u7/lYiD7zYK137eUadSe5wrZ
b2LGV+pf1EnWj/Yl+Lv9Uqx2/jA5fWIfst2FfvgeR4kFDtVQ03WAZvxKcN2MvT70
RpUgzNlh/VYPzw4CfqEqvR7GIn3xD3G0nfaF8TG0nxrdlFBs6QS8pPQ7BRagJd/2
+b0/t5VQZ2X1DsM/VqHLTqGEIrg1ivV4Ns6u5xMOWHVWiTGVRLeZxPTvIiD9gCaQ
VMD/cXXSqe6e5oB2+nhlJyAYJOSC0UdJtRHHmBsgi1cCK08545BNGSibHs5iZ3LL
jPT5nLOt7Zb+q+m9Uci+FzsuKG1ZGupcK8xFA1gOQO6ObNEHF9pW0zKMqMX28cgu
ZbJlBGoj2/RVEDjp1hhXzjDuOF1F7FK1z+x+CIxIvbTv/X1sKLIptQLO81Q8r5KD
9VPf2rnj8PVDCKmIhbUBb5GZRSf2YBGRK9KbzLrTWHd7WGS5A3eOuivh2ybazi+I
K1krjTTK5Y2oA+kPzHxAYE+nAALomfHtlqEZ4K0LkCt32RDa5nqsJE7Ic4UB435f
U95RIzjDo7xgsrBzoyw7KAnZAjfmyBdkGjeVTt8pjt66c3+2i1njbcxPVe2egdf9
U8Q2KWnfeJX64WuGCgEgSZkDzySFZxFqIdHaLaGsSMHHhyLuXgUTBp3wOLc4/X1/
PFkjxvZABjLer0JMo5602pyxDXdNiMz0c7p8xzmIGtfVD7grJlJHwTC3hJlC+XN3
Mz6qHhi8zT0MAwFUVhtzu2IVz1brU0anIJ1FIcQJ3y8r/eB45LgS9AvPO3mEgT+U
HiQ3+s6Ewgco+Du5hi6D46pDiwg42k9GbeEIn0KTTsa+IrurY3vOU994A3FUqjwv
JW1x8fUH42u9F29l3ycC8Y69utZvPOIyEB8+7ov/dIKYM7FN7Uf7f0dkn5l+1bYB
Rojnf72W4TU6dbcBcpOdbP3ebRdpmjwhbHTB3stHVkI3zhiEWshzNULv9jWd0wrv
RwWNBPhI2x1f+B9otyRtho1zIfFRU73RzUJcURnMGDKNf0lnVi6+F20Kk7YjcYTh
sfya9p8X9/5Ou1fgSW+dBXU4CFBcaRVzVDN988i4NzndbIpY1ggxd7CKafmFS5Lq
6W33U9GVxXdx07ayclzlS0/v1pvaVf3nVkkG8cxw2eClySxC953dx3GNWkIt3m7K
+nMcNeiWsqRdqW7UTtAW3mKEeqk6ifJV6KAA9LFvkdN8MHxy81WUEo1NPJjZ/mdc
JbGOs5AMeSe7w8AXMxbuBD+wxphDQNOIXL0FpIML4MxgkthR4ZiSF5Z/nL9hUUlv
qG6j/L3d00lw91Rrdh2zRGL0rcrqQE75InTBzZkFetaFxv+zZ5qXBb7+qziGVLDw
iniIdoXyS9BnvN05P7Vo9AVLoBUSi+jioMvLWTjYYbmdNx/ktJBP4iL5M/Km89p6
RXVBXXKfpMNsVrZIJc6wj6CztmlSmcLTvSzPie7dgeWjABYeuJPU+jX5D7eZzd61
3T8N6amRVqHY4vu/qPCinq5TmPKu121PWstirhmBRdXMTBMs+AvEIcmpq2SeIwrr
GOnRClEF4UTDpYP6pU5xxoALrloPbL0iHpxsBA6oPUIQ1EY+SVDtX3gh1YFvsB97
8f+EtvCw4eP2LGVmRit3+C66ISkaAL/Fin6KGFCGCaYpPr5/nlG7dherUDdAc29O
pe6cif1PrHQg2QWf5H0sngFui2Ve8gd//okqlObaJluyKfIjBB6dclqD6JtqLWhE
bOZr1HX6T1XXg2lK1LeB7D+Sbfv13ChFNXMYFEYBYSpMY/ECxk4xCNTAF4ZvwzZy
NF12FoHsv0S7tFbej5cADJX6hGbZyKGleO6HP+ufQLTBJCamRbxSOsv3faaZG+vv
v13mhH2LXL5vNboVC5IVsDSGoF2+iFApc3kelUD6SAhmDh5pfm2i9cyS/Xy1OahB
BKr8S+4yx42/sAqnAXY1RTfoAnybPSCKwZKzyQk+v6c+Ij7xZeqmGmt0UZBbXF2o
PSDp5cdp9QL8ogJ5+N9sprcP3rqkVqSXiDtAfEXrWxSQR/YKny+wK9tTT6HCYw/f
b3GgfYt9ubo5/D16aNZGM2B4K4ZgL0pjf4k5BakbTiT/tkSEpRB7WLNc8E0vXDSy
7Spj05zgZPCUPlZL0FDb+ukKxgEXsX2CCQGzsJjRz472RXzlG0VU47sDWBIngIcN
+v0KTbuYZIqe7StWw06BsIv+hKAC76r86+cJF2ixo2pNc6H74bv6ggpq+BGlLo5U
wNL/WthnsGnmw44KCtigvPa2QA+LiHjASY9Ig6ZvhkqnuOj/4RoJkOsf998x63Vf
Y/kscRgjaX67wx4Zk+uyw3ZgMbqhLKhRPfxKCYXCz+6KCIFn9nEIF9YdpCnUcAec
cE4Ip3Sh8N9X+a7rFRxArz0hxQHl7xLn3jxfWskR1fxZLi6TKjTpfp3z/asqFGmz
hmNOjzTfM+uUIdXTkNvQEXYtUr/ti85WJUXqHpOdEjY/Py3wmx5BwNHZiyvGjdeE
r7ajww9gTlkcSFREAkkLN1FsBZxKY8MhBCjapTKN+jCeVKde1rVD9f8Xrpc3sk2a
CQyNGfoZoQ3KNoVBWPp7RTP2Uu2fmMU9XLU7hVk8t7me5JV+6oFTZ+Iod3IwBBg3
Ems4Q4m5Fab+uc0LU/ckmkdUBDZ3kgDt1I0AvB64z43UXlyVRWMr6YP0hNuyNWOs
Abk9+8TujcTHbfguvm7ZB6N9q/L/+sb7OvlvI2oca5DaZ21L8qLgi6fPuqknrMFb
wdt1xPiwDfac+QGjjzBog4yqjUuFBGyUAEtKG6mQChPP5opPndZLytApoZdudGGM
Uv0xpVO0fzclLUXznV5DSc/oGnMk/uZyBiwn06PMhO4FS/1CFe+cSymSAAwGIykC
CCVpU3ZWjjdn7Zpxl36efxXQ86yMBskQDYopvOek0gZjGRJDoKlZ46gTQGwfo9+H
NHRbqgRAbSCWFu2hP4MebG2teqG8h9SusdIsrnz7/v7fGocjICjduOz6gvF0PAgQ
8Cb3iuCdkGVnf4rMSJeLL0UvLSuprPQvyHz5NUjGXiLkunI5GNBSXVkbF9XH/dlH
W4xwjM6FuIRxqkInFAQpYyHfZUoZHtj6r1KwNk0nExmmHlC3bmPf7kNVhiZmxfCR
4fHgHsU6LyXr7pK+lnCKWzqwlsO2bBTe+PvCbaY6URoGR082fwXSkRzYVrh5ImQb
QFd8Txw47dSDXJhSL+XYajbo0PEGg8i9D6N7uTWEOxrX+48F4FwJA25Ug566XPuc
R42qkH/aVNcag5GlMXQO3WZ2M/WMRtfS18AsG2eOxfC8ShE39qOEMBIWH/bW9xx+
jCUNm7NGzQ9UuCeoT2qfsUIVKEzTFIML+A5tXiewL8y7ChEvLPzYaIVI/ns1DGrM
8dSgiImTOdUmgf9omk89NgxgDBRGMO/RCQLeMWatQWZfyinSBDjgkI2VcuZZybD6
eaInX9NU3DBe5eRjx7oVQ0JAdDalhL11UGWaRdDLXySEvD3y+GJcZmVULOg1/Wh5
HYdcOkkjmyK/anJk0k22OWmuf7KyeXx2kyg0HvBC1uhxsJgV+F2Zpy7rGICCBstU
sFEEEmWUiJBuBWRxafOSSNrXucDsrbX9KV1pv/IaRJFhmREO+Fj/Y8CGy5uj/gtZ
+8SiIT4H7tcscenVd4zdIXxhMpMbkoB0V/3beQHOPTY6o5HpKviMwUG/fdlqTz4V
51l3KwvAEXsCUzFcnQByy7Ip3FivbtJNrwDF8SRx80jl+FU2dWuT4xEc8id3FqFQ
aY84/v402v0di+h4YbeOwK0w9IsWICYM+9QyMVa2nctib1r/KC38v9uea3h/ygXK
UgFJZsqRbZrRri2y7hpJwbHUDdT6+PrhbYPtrt/wIWSMBUvFf+LE+H+eFYY1/RFv
hL566/1eKksottWsgCjxcK3ZcvncOCbWQl2VFL453v1S1aewhRjss28chjP6kJnz
NDYqACDtPC1oT4nMbudir20LrIPTRrSxp/9Nrh1tLiQGrMVTghdtNaEys5y4/KX2
p3U5pHqTKiawtNIi7WG37accph34zTZKSNIVOEcZiuaDABJGLn9gMbPeH+k4qc8e
xsiIkRFdbwGygzxZfcR49Q2gwWjjwTCt34dQBDmm37bfvA0XalO9QzVL2iHsWXv+
27GF7xxxRYfBijjcfS7P7OUWvoD+smlDfLYRsJVCghCf15ZD2ApBQkZoc2DRadmr
lOGMP44BKcV8o9Oljl3Va2ubaBjEi3njc1pwczSG32ETEo3n+fp+RG2sYOloDxrv
ZhESxFeDCqVnNyM74b2FfP5MlmR+BmX242tqnT30qGOnhxmf9WmrPXLHnNbBbweK
q/3N54pVCEpiiHMisRkC4+zfPr/TM7atwUoJtLxCr2VkRiunu+qINdCPa4or3Anx
qD7CKCLui57eUl8K2cxwIaRCI+PSHvFgybx8KXf1AlUul9t3Sa+Oz7Uhgbsu5ReE
mfRCpLuSDDCXtTYroSxggqRteURNj35y7tofHcjwKJH+yLDZq/cl2UxjHyTMQuVd
aeHLVLbsN/o0TSFNl766yOstRVZuABbYjSm/vBzTpRGNXcrxeq4uR3ItacucspH3
AgGmx+hx7ztD5TRMGllA4nef2BCjn5banYqx1yZqMn7hVXMRgRmNPiHzuPpSIG+H
NYKdO3fIyu/YSMvUIDZEFdHhEh/eow4iq4mNCgBPO9/mKq7DPsavelJDbYQ3Wn/g
1y5yHgA5vUiIAmyzo6bmZWjMXfuVdhkmMi9FkldkQihOZijCwNwsl61U2i/JEtWl
UiX90y/XAcyXe7K+L5Hq6LOgEWTRoibebj1I7IBXVxhvDCziopqppG9WOqHeatD2
+Yx6MNMhuKbO8NfKJ98IeUJ5/AA2ReZOTviLZxaMwSBJthLedQbuR5OlyHbY33rn
1BJVU7H6axdiWNnUdE1xs1eZgJTXbSlseEeqZkM0/OttJOzL5/H/CdQ75PATEjHo
NxlaYvpLaEyPtF7T5NZMh0xNQ1vU8wZsFH9g6nB6oo2s+CWP36UDib8bZrhyDAtn
IglFv0c909EPITsmBJgqVLxBQ/Yn+C4gwTWbTA4hvLrayd4lM0KK8KUPGKLTWETz
VEPudEG144AiEtEJBd6Rhm06nTtVyhcnVX67nT3vszh7i5cRlVAwn+CoNg2DzKED
lOavo9wgst6NbOrEE61/ONUuHlcEJ2m3sLfaUeolHBj6PYoEZO5acuCttONsVbHZ
SjZO2X3ofAm5PmYU+CiB44oT9WyfQOhChQDGtQnvKxATCL12s3ZOM1d5slAPggPd
bgYMgcTavVDOcTCABFG3hWdFAX4+2zokQ3Wb2XJZbTUfFH78YzdTMYuwyT5jt/0m
Bs0FmAJKer65smcraZ6fapspObBHLT5W3P9Bs+mU30xFeKdIbErwOYT3F5NEAOSm
EXEcd+lFtGoEr+mWt5DXTagG+4EVFY+b+VZuFIzmm7Uqoqx1I9wysGACk3oLXsVg
3ThAMKBepg+e6VitIdzKXn/s0s8ja5TTHAZ8Xw2BM4QUcWRS1g+doJcnXX3b+vHu
jvO9347f3DcIWNb8AZAMxtaFTeCb7nyjWihuc6czfKZyD5gkunqk0D/0/soGLsgi
6nHrR6ojXq27jQm4ARArdnGhO4rwgQwKTHI5C9bgjbhNEUXsKrE6Nf1t0jC7C5iy
ftttOdAvAXnnM6yxrdLl5aM3Vpj0J1y8h8FVRsJvbIwrF62eo2WIcqNadDPO6xtP
Ca++W/1yP+2pcDIxHxQVnluXt1Jq9E/OkxcXBrSTNU+Mvxcw+iG1ucKH4nvCdyEh
JTM6Tc8zD6V09Xaxfg5F6X8WloGBgQG5oQFyc2+zkhCwW2Swa3SNZTjejWmiqDt5
yvpUPzwbo0UrzDxbM5XQr35aszSS/aUFhzdFBE6h1Gaa8Fz4XJF8tlVixD9FLycQ
NoYRCgcxi30242for9rsilUKu+8j2njt9YUAhXFpBcuS18pF/kdV7wKI3ItGxEhF
FUMPgz3VuvtSO+BAxPses/McE5ZB0AZrVeefK9tBFxlnVqXurR/LMT6Zah82wBo6
khvZjk7PdccyLKqwl0XRCZC6ulmT+103tt+eOyQO7n6Ihy8Ky8epbjjzv44yn0wC
qbwG3yrzGLTJyU8G9mH5S8I/yWZYKsr8/2ffrVdYKo5xGNz0Knfx9PXR0JJ0FduG
t7wUxEzter8N5HMNLtbiq4FFpoqtd/fH2e961OgfMrHou39FLCpaEbFO3YZJcBSn
O7r/d4p1QqWFQuWDWJFsn/KDIcRHXP6ZjdbY/Qf8RrdB/WU53pSyTQAo/dEukhJL
6TrkSmFiQnpROuM+3cRPXNsjnqaHJx+XNx6XXw6AzLhdGJiBjsYbfbj9VZKf/yHH
qI8aSZZlq1UvhXz3vlOXGbRLGzMaQjK1Mydw91a59y5lHfNZHg+ZPAq/39wWOZWF
MiZ7u5p4+tjU0+0568ZSp8DUnK0RXOBy83MRvL7NloeXNDiJLiFt6d6UbgSdyNOa
fZcPLdLIx+3sym/8uVdgq0jzEdmH9sTh2x+Fz1ukBiMFS+g2HisVv+huFtzLyKA7
Q8xmNSSH34Id1FsB3rQ08HDRopp+FC7XDDbaetZAgP9gGkVfNJiYNxGY77++LmMb
Pa/2yZ7y5lyxMUQdUcjtrEADLlFsP/yKqH2rgdALcNbGx489782Laazj0VjNqGmE
pQou/fG6/oYbEuL9dRfAfFMcfCcKCIAFyC62z3a6otQkKoWSWYX/Ww3jBgEz20jY
5qUHDD/TP6Lz+Fwx2jbp9/PNH9byFGxdgnirsM//BZhaKDmMF/Z+7mMng7z4Jobv
zPDrpCDgfBJbeJe920I2k2uEfscYevC4dVhStMlf2nRiQdMRq1FdkP6F5v6ayY3M
+GQFeS2i4zTqeRG4b7rf2gFeauHcepgU5q54Ln2TkEF3zMbDkpzf/b9GDO7kyV8n
pgVGXF1TbUZZfzMRPkPzyadOe8OIZnDw83zWEZokCBzbfj0rPB2XIs+TLWJjBoWg
PzGgzVylbEjdOKkaIY/qSEmDmyGKXbY34hnteEp6n7auMRwwt61w6VGk5f7VfMcG
Kn3QPU0hEz1frR8k0K/1Da//gWMy1L8gQ9xH2JXynkrWnUunOlvCrVFQIIdwxgzc
IrYQ3jvSaqejBNcFhKz8iwmrB0DB1mFFp1zpi63v62kHuPjGAiiBJTUnSU93j6vY
ZSD28A9p0dAVVq3ZBZBj1vpYQPrEXAbWn+ICl0DXfH/hfiHzQDqeaPQeS0S3xeGY
saNk9SrF5b9lSVV/2zuwvwJ+J0r0ZB/QonP0MbExfJngiWV0bVMkYAuHco5B3nYM
+GqBHHOiEg6oqjEm/JOBO+P8DmrXyUGQPJibhCfEWPio4ROti9K26r+Zovu51BRs
TtDFyqpvbuVcbgVChFzOmLnFSWznzOslyYOH+Wx7tTKsK1E9SBmMPnUQI/lYgwKh
9E/RLZqBrC+Wl2gILEkELUbEwoFxnOtXgAABWpH7P5LCCH1wdId5Ho61SRAc/5/c
tpwBj1UdmrlAVoMSPQxbcpV2sw/vXpGezdBWaziH7p3e7pUFZcq+mEt9HTcCB2S9
NhT4jUnCs66PqCwvkH+Qd3du33jTvjyDd/JJyO+6HBTinohxQ9xEPzkvj2bzRGEW
e9z2OydLQAWJfcRJjYZNDcCUhArDbNe6CfGUGdMOS4Ul7JH93jmy0XrCKVJ5mPru
/uyPSTPzy8ftxCJhsUH3ewVEoYIYn1R/U0W2P7YZGLuJ7n1nuXhtVgn7UQjL656q
i9WWXnI5ZNkETSFwq72rDSfvemI54hKjXDqF+H3uMYjlKO1+yu4hhTDFz6IhO7Ou
nPr8xvX6wBTTcSgK8l+8nRb59M7wKokWzZq/uz3eD1vbwmfxxnC1BQj+bS0+97tt
d4X8UC2hBOPOewOaMKdXOCB6RC4lAe35UGzYQnCTWOgRFcsu86NlHFkdPpNBGtQD
xcaZpZq/WmlKs6Tgt9Jb3/fjGpR7b7aex0mgvX1bXysmMt5q6TbQdO99qx9DWFNb
0HbTI3RuIXncwzNNdMyMEEm+w7BXYUrgtnfxzM4qH5ZEZpKLTQ14z0RsK+l0i/n6
e/RN1HksKGnmSosfV7zp+3nwIdyReG03DGlI1YOMQOY4NKrkXv+7aX9Z/fiGODw/
r8frz9OmydBU2ZgJDJlPtf37ZWlrlk1djRulWk1hSYlfNWv8Q0xydDulybwBKim6
aSiNe6kBdiET1Kk6izyTPLuzFyvcN33cTa2b2SwOs7XtUvF2AYH+xy2DkmzOhbqw
H89Fy8WGdQ5dOk/Ur+iBIBIqetE83AhUfwAESg5xQ7UG7THd2c57zEqfXbUxEP13
J8azOKgQepZCf9DPtVJEXZ60diHO5uPgPh25O+qies6G8jWD1gO5RuFm6JU7ywIy
dpVPTcJvRKMyBOLO9y9oqigGsfAZogWYsW05sxCXR0H7lLectUW74CEVehzgq5KU
W3fFCWaCC/1fw2M9YLJ/3jDQ+bfQSKVdRQspRwalU34Nky3s7IyQEsiAovWstEFe
kLXqDHQjSLFU1fPH5GxlWgsmOCAPyK7ABUFKqSeIlmBUG7Rsv0nYxLeuBud3nIby
4/eRUTtC6Q9eU7/NONvYmVQxcz/GwcIwNV+P6+AJAqjFitE8Zk8FiloD/xJmLfZj
28D8YV3TQ0+bvWrhfPI53yql+QTcQH5U05KrX1l1JRqXdWbZumHIwixC0rKHv3++
Ncla6VNjxIQPlQDvS1lHK9NPp6S6V+Q/iKEzrpU4okTDuiESmIraHiyzW4Nb5Z4M
9o9bUvtOtbeffxrjgk6QYhEvTfB0Y5ebHU233rWlMsVMmosSLciOLNr7HS9wVHgf
F1Wn3a9c5eWsbQpWntYf7/FEOHfJJip17ersqnPvRjhEzcpMbpFNxXMSDnCQj5Nj
Th6WgSIzdjWc9MRqJZr4k+wKYwevorBq34GlqvXQl1dcpjp1jcrANrt8BsjOBU5O
HKlwIu61yhuQkwKKhW6eqfpWcaosxPvOO3ETmD1ForK3BUVBX11/H/YYY2VFguDz
QIF4qXYN93Ro4gBrT35Jzq0ATs01G3QRD0qzUV1Rl6NyuAHOc8AOSeS31rhhBjmA
3YZlx39lDSo88wNduPu6q2DUbxkfU5gbPEJ2GMQ+kSyI2DziCDPeaA84ayj+pAWG
V3fDBOpxO5hXdq41fDiMhXi1rmso6sDKSgwJMhU3BBG0uinsdeKNrhhHVpBNYg9s
qc8Xz21OcJHvYrfj8VIAdQBlFdNdQcSGBCy0oxTm7ZjUJSoYof5bxFFFi6YPF7Lp
iCe+Yss8pqAMiqtG/FwL0U/ms1LF7r8NoaoORPhgwaTp7GlAK1AkppARpwJEtH5C
LQhhZbgIAVU0HrmD41xDodzrvoPsA69+gev5BX1qUyHe+WE4tgmPEsJgoR94LOR4
KKcd6jWSiGGO0ValmMFAFWK6UZJnfkh6naM29z0JXNDVssbLpclkxEr9ra7vp0/l
HlnvXT9lu67LNjkvnuafKqotZ8BCssinZ36wCM9oE+SbQimI1IXe8WHP9s5Gvt54
0bdgWP6afBOama50iKOaEl2CbIlBCoqekpggrNWEZBE7nGpwlglEMoy76WoP9AE3
1FYrSlni1SQsAwJasf65vDVZvLMCwepWQq2wSBXzki896D3K4U1e1wZKYFnQe0mk
CFbq2kHPAv7MgDAH3B7XoTtMmYXTi76oo9uH8hsUNIKvH61EM330pn4tuIor1vif
EVLmOkFfhFzNfqR+uYQeg+GR33TDs8IiwWAUSicr4wOnqMWqkevIAXpgXJxNcrhl
PDGtulEBLQZOBEtM6tojqx7toBEV38ln6pvEV/NlyHuoOrjZhI+uPqkURU8RDQRJ
1hjyHuC9J9fyZM1ZX+WDikUWF8wmU2GHh/mQpuTH3QlpYGynbZIhctX6FIOxrJwz
QG4zqVdJA7L6wSEmFzqHHXcA3qNcMRJ8o6j9XAN5jwQ0fI+eddDQue+ClzCeH73k
4qKJ/tKvBv5yOxxENUI/zJrfBiJtx0NEr23quW99imrgPyznBnTxTxYMaA1jSjxo
CAD2fYj3stThbbesOcUuluegnttrqGYHY2jdJouhcYerMt9P8GuGsrfbbatUsiMi
eSyRm4EDxdJ9DqYQY18lPSiBInoViPD+aT/63TuYUln4SwkPMXeH5/OWZmwFvSKn
rgDiOsUBB8KuXn2vYNjhkkCY4UcDPoWYOhIbg4jm1qoChIc5JJeqGdWV75vJxxLq
4zyQ3tNoprtKYtwmUOmgzFD+kFb8Ym+jsIFoN6KFMzg5L4Rn3f2zaf8kf1VXUYkp
OKLDbpvY+pHpN5kkjmkpPkhzz/km1weOHvN8aEQOVDTg60ozg4k0IanlTkf1eNba
E8B6SqwfgsQMzjbs59FZ4lNCsDsd7UvgCnIantqjf9lPvgsSyKkQidf1A+vNBw/u
cRqF179ADk0F/s/X99M+3HfOilAx0za/ySO5RmIA+zZxhlJJBIHBVemo+xfhsZUy
b2PnPQTi9ThkCvE6N7kesXC5YmC+R6PN9ni1GzXEVNaXLye/O6gAF8+uqI8Ypg/s
xcst3s14r6ZyqQqP8t7XJuUYby2FV9sF6iaZNye27Z/Eaia9L3E6UUVwB1m99yGy
sK6ocs4OrWiDoeFKfdN+RN22iglq0amqaBNpSNUqKWpkcktzkHGS9zyPvtwAX/A0
2jYco42r6KpSkf1WOenQGCpqVKSs95bLuZ9m8dnq3o8QrwGFJhnO8JySZdgAHNeb
BW6MNyenHGd6czi3aMaW8ZLrVXlbvJYEkadAUcxo96Y8p197IuUTnM0msti1+qcK
aSepJ1fXskwoFX/nRRtYZBVMU3cUVEF6RksupdknV9Vc2XXSZYdU16EFQMN3sKm/
NcmyDmfnsLPkCkaymQABKatC4BZjJ8Gac0TPY9MLfMoToSbQy6591qpnknisHYFo
pD9EcYILxAChkq+2ZZZIEk6IuLZIJ0IpCcI2+c4mdolOAqJ1yWRq9uJJtA8DUXLU
yBCHIeqaxs9tmGwf/COJ6vr1tv5ukynCc+sg5QilqPD8S4sWbt5v4EwlTufV78FG
B2neV2S7gvxQkORkX8J79ukpK7AinvvsBUzjlS6hYIqHPxCyc9ajPj+LGttxeSe4
34ad+S0EE4SkxMZQ1tA7uiinYOYPqnmXnoWJ0Gi6KakANRiYMGxamPfSRuELPcqI
QJmLBch/mCXXxSVnz/4MDHc02AIm44iYmTrXAuUW8DzOF/JVg7Tv3TVxZT1Vwgps
qSkPFwqZ4pZa0tVxsz32COTRd2wIkUvPPTcS233Zbrpl38b4YbIod2kb8hqNfJsK
c2sUQBlLWdyxCqj/xhAmY3hI4yvSbjvVP2KEy2Z8X4+8DfcDltVgfOLIMo3pCkwq
K5VPw/weH6hSyHl8gXVCRr+693nxrPlK4CLFPW8v8psw+zE5v4rln70fGfQ1uZo+
p2hwsToeOOpONj40A+owaG+iHBL8LvC335cAT9M6vH0Q1AzkLBIpkkzNQA56pIac
FSJcLdJHiFNQCR2yes5wDmQYg4N6Wpg2Hm4JNFz1+hQrgRB95FqeCLtu0axVoUoH
8X7EFXExI0PKyfEplJ2oI2k7Zm9ihDqT05qahGWwjJwemcVXsQMdsWketDZX8sJx
FAqnqve1V4D4EZwa1Sm7vJl7HQ3bO/D5eT3vNsdgHB7/6aLLtOeRBOlUzlEtptKS
deWD+1AcqOar+BvpkYgZNi01G6ZvUeOitKjz4ONe8P5Z9bUzhIvP4+Ai0+LYz/ju
5IXWQ9HuEde/JLQ2Sfhx87lW0uXcK8D2KSeGLpf9BgyxkbhIdFaO79glTMIdiREW
VzpqV7ti1LcTyjolywxnpmG0H5TBqk/j6z9l0acr3MdrK1YpDWCwVeNUJR88uqto
slxJnSk0+bJk3ZPEhF27j/pgRdC+AYO42XXKWOe9Bal0CTGxUysT12Kf6NzTGae4
WSN3Xp2YWRV6NK07Iah9OxwocjQw2TtdjQTIasslaLt53ycIYicp9dGPbpghS4lh
7u8MNcQP92Ygaxo0ZkUT7HBRUnJgEAocciwJEcbNj9XGkAFJcQrqviwDVAw2eImE
qni2dXY3gJWKtpZlGsBcTlfWv0o9kZEqUj59DBAEw6ygFrK14J9D+gKKmotsshsC
AEjXx+n2ia1nM5RwDEqd6ef6WPSnPl7UzcT1p3uL84xoplvIJ5ofjlMDvNCGgUPR
UuPql8inCujPn8FAShuAlmeD60vH4bqVL5TX7XYcX/snTtHZHf7pcbjHzTIotby1
2bJa/qY3K+h93OPAfmoSFV670Sut2An1F9FJkEhGaKZ4SeXZgoTY7yLH5Pczt3Ih
1j1enWXO7UbuHn/v2Wkww3lMuBGpYxWPx+ExcayWTzete7+E1OUO9++wYLgXPXuK
fVcGLWT62iCKIBwHFrxlH8Vzugi7b6PbNzUhUMys/DXVp3v1jaiJBDADWi8j3xJQ
2YMNslGvt/qHvhN11TnZEUZaJyRMJUISIF/kBbAJNnTbPI/+oacj+Z0S2PH9rmI3
4LzX0u0Q+3LnYjC2rgh9Ecsesr1LDQzMp5LPtvYsKGMhNaRIaNeTxX7dwDggNGIE
LmJWRqEbWrN/xreANTj1BG1DHGDrxMMpSJ9i+5P6zvr5vfCAbWvXs4n05Gpc3t2W
GwQjqZWXmhoJIT1Le3k4upo/Y2FSH+mG9MaU50ljfqO0yMIb7oagoamuqLKAx8DS
2tfaYGwVsEq5+fzhZRA4fjS6h9yqbGgVdEkMvM2BFt5i3n0W+OfHhSReox4j8lvm
K3mJ8j99Thxo90CbAKICyoB1/AH+yKOEDiSPefTeVOauvKEdU720BUyoE4lPgShZ
iekY33kJozXDpt6Smgew5zTGj0RiAxsmAH/tyKASoC/GeQGVH/m7Ed3ztG0+b1Fb
1YI8L5wXy81g36tJijBnuc8XBLpjYIKukEbGCpJNauJZRBh9QijHGJZl5CeWpr/W
fcRZd3Iun7m9NRpLd+YvwJbdeh3fnjtFQ5vF22aPEWjRDD8lyRghBbgqzbRoypxs
NIL4ChyxYTwc2aQ73nzRk2vueraWQcRjU+Gj7J8OCWPuU+unpPql6HryeU2XaqCk
g7w7YDWzMfgcwuMbslgPbstrg2j1d7V4Izz4OWWtmwBAU4K6CEC0wnwwNewlxVYy
6iYhocEdnJW/U+ma3n92VmoKcs6QLDBV2YOEA8SOGjch3dZw/V/Vh2I0+db7VFCg
c0CLXVt7o3VS8Ig27HRI4ez0e9JO2TU6OQ7IRcNPjPcYg2OalbBk58ty+TsPLWYN
TAREO3TIxYqsmUAqoPlIAVLj2/MG/lhjh9n3O61M5cCJ181yUH0g9XAqHF7/LgU7
dSWqYYCxBar+krVryrAnqOrxW2gbigeJuhefQnJSs1XUj9DSZlwsgZtfAhgh56gh
v01a/mRdIfvCYqi2eqakfCSRxX+JZ5EBenp0WaVATONnhM+pDDNx2+dsG2YITFH4
wk9eLtD8+zx6mNnJ5E9WbSAY+QjXWBEP/Lj5vZ0GUas/b7nb5HvIXakfbDMPUTTB
KYl7MDPj1MmJgsZhurOIRffcBMvJRMdwb/+sALQNJysXvhXtMQuQTgBGfQCMAbxT
ILtfT/xRzk2rtI+ryJJCxLtu2j3hUKyKiD9FXvIJiNhIWw02qPiN5MBAR3cT3oYi
T78sPO1oHSHAEnYMxD82cUpfOfx7NljLSOgdRZxhijhTTMD48LKQN+j7wDotoOmY
oH2sZE/z5kCBwF3kg21m0yYOKWeXVbTvZwz25Tu3WePLCaOLaDz/l+m52eVcE0ly
9BUfq0aTKzD+H/GANPBhOctSvieGbmHck50rzGEKtrFIKEf8yqnW53NxNeED1XSg
fn6DYtPPCGyGNr+1shSH8xFPTzwAubSn5IsBE9G/+T4IxhR61pIa3dZMneXfFB70
Wqs/U2Lwov5HP8T20yOUaln7uX9EJCXejLOTZ+HrEKdFWMbJgQTby5wEHrRtLKUA
6SpGALdsmpoBe0z0ARD8JHKSDKY0cnxyso/ojCBFWK26Ynq6ZKMN8/+GCyQrHnVc
MG+DOXXNKagDxmW59AYYbhQ29u0CMZpnYbiPMjf3jEiiqAVsg4vcZJ3tqjHsR5t7
qClpCDsnDbzzLxqkTUi311S2B5ikfi2UONCzVkIqieXs4oLXEpBaeYBefELD6BcI
/gcCqPniEsWTEn+PiNRRTM7YSM26f9tcyPbXKYhUY1eN5rYUWzvlf2w0f+9Jot+x
XEjTa5bJrJMoGGZhI9S9wJPehPhE+R0Iu58L97xOsx3SIYRKw/+SzOm019EpJ6WE
uV2tKTObObHPLat4ktT6FauGDb7r24d7XhcShcChrML2Hq90muf1hEhkeTBFxHBn
uDYRPR58blCZbR33aAKJRFiV3VtgSsy6gC/wIvOT4f6TtFSpbARDHFm0TC9guj6Y
KXOzTC0kW9igcvwLjqW1tkedoskpV+fQj+sbeuCl45FotLV/18OSF8kfyLQdCITX
7b9vmqjS2T1k6O9LpdR68/n85dvBH2x1va3hFSKOgMrzRsp+cn89oXiZQ/Z0HyhP
uP4sERUW0NVAAiBi37NPDWDzE8B1vwvTAHkpVFeJWFbRGW8oxqN0vBUkGXycjD61
f7dIc1W7BEUWA9GWKSaCnA/8+cZTyyToqc8bYkQIdubKc/O8/ZWJNwrGbE3I+Swy
E9jEtEzRES9SiTQcuEIUODHeDEySyCvgkEmhXU/uwYWcNkeRyPAp4Su+ca8rxJx3
dzcMfwohxQMl4JZYcN3f/LYylUCvwsPCulOqCKxkGe2pEsu4QDyJv14nB4R181cM
6GypATxtWiWmhHQzgwtjJkYko9oC/EQ0eSlryAl2dSz/k4nRR1/ozAuqp+vafmrd
GKfaArGNwripZS5NBrhSZ98RwjkLTFohn5ae1l9JmUd6fR0qWk4WWfl8Wqlsl+NM
oxTT+u8XDQo5KREgULVp/3HTkKn3awCaS5dBF8zYiZnkH1e0x2ES9NDeg4XmpTKS
RIjvE5qDAJFfEe1K/miUZWhdjjgEOptGQZkT147PMMBLPZt635ORqoyd5z21nLQc
8JXPcULOKC1JUO63xm2tigtExFaeHN9cvdFyvXlINhKGV9rHwcjow7lZ7qsNCm2D
yc+qcahcFx0IZ9niibndwGQjbgbPF0vXZ6jhoVVSa9xCdDsHeuOY/Tb6DrfNMwsB
Pvso+bKCzh8lnd6VfjnMq/XoJ92KH+9DSjUHV7KRQ7VCZhYdsQNnFYO5DDq2Ejbl
5uUAY0/pWGo1EVXPfO2lIM1zoatbv0b/YVqVc9dp9CvXRZkUVR+uJkFEMPzwyvYg
C9deWjvGTe2oJApKbJ6a0JAFAMwb1aK386+aW+g3HsyM7JuvU6SCFtaLQYtAd0yk
iv1mq0ZQfIzeoS70+/0IQhym1U3w6Mi/wXTowhEzGKc5KhU7gSicjCt9u3CwIv3d
ec9H6HKW2d14MpWRj1xrUFBSdDWXRER4h1BknBFYaqBcozRyLAxdMjBMEHPTy21/
7LPIiSWOhAvw4GCPFSHYtwKDp9EWsqwjGj8ikmY+KaQ98m20cRuqQHBSb/giT9nO
qA1gvSAEeNZot60a+3lKFy9h3PCzsxH2FGMzNqH+7wxqim4eFs3iRGX3w62oXIzy
aghfOi0Dw7q+IIgQZGkhIFjaWQoLRqb5DJMgco7ljJT+cbySwU2bohQ2enURtPvO
MR3Q6QtRGOPAazq5v3l53no6V1QZiB1Hh/77u+Q6wfPdmco/wBpL4l2nJSkLxFo8
QjSY1pWMj2aa2RV7c2ZJOjexYCZSJFxwgFQJv+RUx49kRwKW0Pat1KBbXnCWVTFr
Zjc31kVtnFv8Gb6b/O9QdWyVaMOyHqifIKqedzuIfxg9L54v3AT3kXbQx95d6rpt
eyQXZkAVoVxomdSKCnhXj1OL2TcoX4l2+ypefDKXxGxgWMKBBRResKYA8Y3FQ2TC
s8ayZFtcaEOHKh0Th8KajTCPXKkqHIHT3RPY0yAyug/k8fsb0xxFMEbIgy9sn+kR
IXu1W4vl2AO1aQeIFxELoqi0FzcdKz4OHkMY7UwbIGEs5LryN/Qe+03zj7Oh1DIJ
uZ4yV4ka32FejS0bVrtV3T0GTHo6GAz50A+uaeKqKIhH6HdBQ9OvkP7cOpkHeZ3r
x5/2E6pKPGPV2OKhww4tHxZ2rnLXvTtfkNhHfJgOc8JNAQHtOoNmMPPvdVJiexzy
QEbKW1rUNcsXhk0tqriBzazDtYqMErTvGt47nC/RxUlP0K/JFFxktiWSKDmJjMvA
9p4PJNkIQ45nL376DfX72ddaFfY0Md/7Z2gmkjJIt+oUX+7L/RjUm9Ffk1/tWhYr
dz8/8BbknlhtrjstmWDv/iidIdWvTzURY4LVQSo2rcJ+TC4/zn3C4+bzSEO4BgJx
GcuuylFzxgNyEqyeOI0XhM+nWsvF79iFSd9UYyubOC14Ym+Emds+GlkdoYjX7eY8
lWxeOtEYyytGash/4Lskx0GcftH0Iru34niMaG66eh3JoesohcTQdGXPzVAef8Kl
GepENd08ff+9INbDHYvedO85RJCXH2Gj75juJIe1wcEyXKJEnScHmuT2Sxu8YvHL
14qSuZc3cnEY6td8C5aWH+6bOJz51S+BPWEsSGWBYGYe2vOuhIiVr6hpReh+HttC
UFOO3WUXaXC7Vsm2pZtvF+WbNoh0IumGhT7zCHMwX3Woak/EbNvgnfY5ouh/fHKq
V8Ua0wmg2hcNOMeI/CF7SyE+SzzuUm3nSpMp6MxR7WiWYWpgXmkYtjBNPggydDTc
PaqRjRPIKVH7guE53bwN+ztKjt5ewx65hoP0409O0jiL8D0Hxr+dVxyjMpJvo3mr
WjMnKa49wMfK1LdJ7OoiZenhzS8BbUeN1gow7+WhogomkkgIPGo/56mmtnSjeVS+
vkfbigRGv8utQC6KNj0HqT+CQojwFbJ+hRJT5ZO0DwckBCTvKRdICn5bFFrk02Fe
HwpBnJg66DuGG/OvTffEkO618fIRXlMNyOTMtYSPa+DLhAA31KzWLnKlReeyYlPG
eb6q5F9dakR3F1zJgAPMVkZTTl9MdzP824F1npzzccUo8EKNksMyt3IK7UIh9qPk
XkLZh74tlCiWT1wsXZIv2SiQWXBMDo86Z7tu+eTzG6rLyKuswkGSbqeUrZneXLWP
vq4OjmxTg00djXhJlMizg+ohlBNrqSyroeXwZ03PKhhr4WCiiyciCRYSlI++i3Gt
kaN6lCIxmJMCBqIUz7DZ40qJbrzb1jOaf+lwyt8iDzVH2+aL/p6n7kN0dK2szjG9
G37n0V3ggdTN+Dyg1rGXtZMe5Tisz6QKCJyvXqlMnPQjivGsNsm5zCNxdcJa3cXI
JDwVdXKyhQ3x1oFSNdfA5pMdYzaP/QCURnNYlOtQ8H549a//Y/mNY7tEbhfeeRIM
EuKBc5QhOCwfb/4FoyIbZCKlFrmcPTd71O0PpsKSBMDw/aXEqHCz+DLNsVryT1/i
ZRIzBF0XpWID7IfEdqQOIPzlQ8+3OZlSksPe9hbK++vy8/JwGXqycNoMX+TBSWja
428TkthMZh6XzDurQwDNukZEiHFRuGuYjN9nSjHcozfdYP5LTyANrTlQMYlhCNpX
wcIr+u+bHRR9tOC/7sMrDW+Sb2R8CqxQnJWQ83LmA/y21GjL8tl+jNfHSWyNTdhQ
0Y1v18BGJAizAN9WJy4EwSBrQMt3v6EMKRrsrHpdbDUjEKoZQAFnv7M/9FgdpzgM
RDFc+pN1/vZljziPliWKPG+ByHMjU9Wrsz+SfkhAHY7RQ/Ds4HrdoKUZUOO/3mD6
rU/YDkbz7xQRGnOE4zzYkJwxoAHfbLdzpxEUT/SM77qdDeRALmplVCCUbi3JJRt5
rnbCJGfTXPN3RNs573XqACD0VVYjHKEBvHYWMl7w9ZCSVyKhK4O3diwFCnVAkb/1
UW967yUGXdYvUiu/whHrhSyPsrkXCubS3SBWtcYKhGOuHobKUwKH1zHh80MLN2o4
3tolFWZ8Q7xPQXZaMk1N75PQFAjTqF6AU6m5aOf9FNAP2najZO/jGDhyDmTrj3uN
03Esx7tplIUIF9hJGsqc59e3IQvSBTjKrUAS5nNgUIYXF6niwgdduKgRnkSHMo0u
shOUcFHMShwqJCtnDEiHy1XVWgxkKSQaA6+LNTiTmQ0IAISxTr9nCxq8MsQl/s8y
v6v01x2ZLt2nicvRGsdu+bXc5DZwqcQjE4u5tIYeHAvyOPYgO4i8fOVVNC50kb62
RhZwQVWS+T1PKihjWQdhcb+Yi7fWzI8Ie6Xrf7H6vfnX9M9E2sOPy2mWSlMalsxZ
pGT+3IMtAcOZj5H2p5Oneqdn/RDH7/F+BfAwagVb6eYVBvjcsQ9MpWlFtnK6ycsT
2N0Ilt+yP9gdb883iXHIwlvnhloVFZ0luENGywtnwspPDUVTdG1VoTr3iJwDeni6
kgQkaddHvtCfQFCWD2nGIekIuzJD88O+K/Q6ULYIj56AcjW+g9FpkC/s5VWJ39PW
siMDyZDDxRHDPzR2DU+L4DEK4vfjSsmgrcvdMsAUyU6jjLeWha2fKH4lY3f4jJx0
mU6eG2cAWkVBhVbUmF4sSKcZmxsW4ytOe2S1N1wVf7iaN6hW8O1Y6ubNukiZkY4N
qQsaM9zILPv58kcehv+ecszUdLIkR4aTdYTkmALva95gJuJI9wHbRcPEoOgDbUyJ
oOFYzgKmS9VIGI3fdcsLbwznvFRiVP1HoDS43ImRG4R+jwo+Lv3y5WMT2V1P79f/
r2sOoEkGO9kbg7p9qZjc0PpjGmW7kVMUVYIj2jmSe3j8aGVm0d6sTNJqtbRJyFOw
r0Qn/pfGjHXwcPRljQ7MzAjLBsJbSeYTD/2C7v+6aTAl+43CSC9A4ps1+KHH16db
JAUOuUFqTRW/sTDFEBRAlu4yYH3IYK9922LFV2RMfXrz3ITutCPwt/AAh822E4eo
xTzWVs6d06qIb4gmgNBcX+3CZ6VkvgKFIOQlQdlGG2eH09/d6pwsKOhqfRrGLf4y
kY/ke4fz3SBV95UlDKRgFQSuDiY1+5I6I2tZvtV1vs0mX3V8GZKhBr+johXCnpmB
XJ7AWvP0auhkWGANjmz0Bey1EBwFQ88lYo7q/YNYiNu0JdeR+kMkaJcpfwNQVQGf
jiMvlYsYqzh9KRbPnlu4fzrIY/px5NEWHNqLzAdHTPI2U5WYX1tgXr11LJEM1Mbl
Lt5carI6qoVYJxA1l/joNJ/w600hq3m9ulC6IyXTfx2Q15ADbUnso6Mw3IgWU93c
tcEZ474TaFoznhcTtbpP8y6gdRLBl/RSplc5wgxIVzeAmins0FMcm0fmQ1KOCm80
p+ncaF6Kcbzz8yVXoWGnQzfVwdKm3z7kOGO/hPQ5zxXTrnj9makpz6a+FvjEw640
fXHk4VpSDiR3MS/iAW1crwPRH9on9lNr8E3ytT9SD1aZFLy/8quZbBSF87wgOoZ6
B/WOyVX3IQI6hJg6aRW0Kl6D08yv2Q4CJtEojRn/gukWr0/QPBayKlph4R3+lsQr
XolitVOqzG45P+cEIfb27FVlxVGpbyjaUugXLFW7DvThgR2vKWcqRJK14X0hjIXS
YBkPsaTeCS/cv1fWlhw1XSETrQf25Vklyy3swVzfsfMJh0tbnyCCSsbmMiSBsM4x
UgVBFMj+0huWfZmt1DPFUTASPdwYI7IzsrYpNWmonuHPQ5iQdIzI5ccLYtkPLwCV
mVVBa2e+PNzjF07Nfq4sY1XJfevxNPr9EkR0B2xuqTg9lUcE1mZxiRxpjLiPfMMw
Fe5lQA0rZHQnNryNlD6QQoeTjN9yxFk/GET9krNffkG+bCXOqYT82IZUK/6zEXNn
Fjw7mOOzhPtqGTpVz/injdXbWSoP1vor4Ck4FAErXJ2szKBiU8SL4fEGwDlKbfHC
3RtlSciLWJsNt+oBHVcGTazFE1UP8oJv5eyFlONCcoURDsh8EE2YCSHMfVQGcEyV
eChe9WARXpkEAFCtMfkJwS6BWAw1M+aDNWXrHSKxTVfWj1XWnNnegFVyLvOW+8sl
6F28QbjG0EyH4+Wyd+1mhojfaoyZlGwofuKdJMSRupZ8knBzJAVA3rEjyY51ah8Z
9x5R+2UM2MFI9rL8qf5GvjY4cX1kQvetJOdr8GmcLDKrdBSjm+jl7Nw4eAzQKYTy
K7tkRS7WBCNaRLyjrQq14KqOc6iDxsPZaNAjOeZNV94F30ti1HLX4BNQrKM7TBWN
mX2K5elLZCauHuChYjPGg3hg5ymxFa6m4zcjX2L8TJWpIHvuWtky9hyCfd56R0rW
J2Ts/waaLd/ZBZenEjzSrDNYymwoi3oSBhSMyyg1G9VfON6d3iLn997ez4Oo0Akk
c3hd+5wdnVWr9qVVQZ8jswjkX5uytG7xhMpOWYMUw+pjVaRA0KFcI3LI2DLZgHc9
3agdDIuA91rLqGQ5e1DL7AS1fW5oL5gyDG4k2UFBERH5smFVdTihgNCCiKUN9Caa
8Q8Q9MoW6+poNThhxsZ8tex4S0F+/DyjVPCKTX7x8v0D5/ROJO948dyGjj8BS9qO
6I/7+o0DaJV7zhDXRuj883k4IBymN0eFHJZSoXhC6qi8ggURFdSxA4Zl1WAt/Pc3
jvHnYgfcPW1GKHEsbEmko90la/y+i+oCL5dgdOPWwBJsrY90X3veBpytYcGTXzW8
DbXlX9yM6XUtbGy8nHvNGD+9ZqnLq4X8nBK99rVGJOMwD8CRC9V+FLZX37fSD9VO
bwprV5Qo8ucBrR97zpfoBVxLQ0Ur8ssxc1zBRUJk+VwHCngzrmPJyPJVhjC9Rl/C
n6UykLsxKkDB9ffw5scRPRxPPGt6qL7fYPXX+u+oer/xkCz3UJtsm0zqJwO+nUpy
69oqNo0MxtLjfnfgBAVB/GDN/ObR4duwUOlafwPbKuEJtJJsvUJc3Qev7IFq96pt
+0tGDc1Xm2vJLy2jT+Y8dbf7ZQRdO3fTToskdr02r+qHxCGj2WLv+1rmWKGld/jx
hXA/kaF3asX7yntLf3wnVbMIlEL4Xp5ykhYGwYABt+ruI+JsRWfz4i+y+YvxH6SQ
/4ezvJJPKD89lgErogjD6DeCwAlv8+cUOe+dWOqy8XTKCUgoTpSWoEdTgnGit/Mw
rqtPamHUpNte2DiYH9msjXbbMnUjWo5+RsAKI2iGmNzB6hmIg3KS4PhHg/GIZp4w
Jo4pSGfnHTD4O9ErRIZeKW4DCfjuGaI+lGsiiMWqR9eOI5fsLPDZS0nGCW9uCkK4
Ppx8Ix+5l+sn+TKSXP7rfc4rxSlfhZ0rMQt/DkdhqcCvrxqJMXFIcgFDfBfg6+Zd
MiwppHMpoZcSSofe9zdzr5gasx03Wf3VXjBMkVv8N8X51+9eWVntjNKpbocgWKuF
f365cuRnVuP1+0YL1oJXWdU70oWqtCQ2aV4tz1mm1QG6GiMPCq5Bf2l0Md/xRW64
T+hZ0Hrh/UzkGbf5hqfli5KYEaGUhS3rBp8e3L9We/Z+L5dQPPG2pxHw1uwFMZDt
Jzm6rFPmwnd7XOrCD5hWb3C2AZWoMiENVxftdEXjFa9t6ekn3S+++U58lHhYwGgG
ytNH9mMWkQMngcmGuF7EkrPE3++YMAHSAoN27f0kLYbN0FhdK55ILYI0NTAJBzy5
taRWC0i53ct2cPJh/T9zb+uUo6l05SGIPs+PvI95X1etuKg0Ok33dD1ShULtz6zo
1IgIgQi7Qe+s/aOqv4fCe+q3VWvsonV8xO2pI8BfZl07ns1L89UrCCGXry5Vp2pT
zJF4wAClWbPFMBVXay1/LCu2OhPiLYiaHprY6gTQZ2TkI97tI4pbi7XjggeeRj1d
ga3ynMlm6sRmreRvbRFrKspS+4zXrUDko3kI7CWjbz4g/4jIJSyNiop56JZw5X32
oBsqPvsk6km/6rvU1zC1zxR1bBfawdpYmT6CC9U1VvW5NKmMI7cY2GQXxBEtyF+/
NDEENH9Qh7EBkBsnPpTGKT1MSXH8dzOyWytzJHVTGTpnmTLuuYKDyqIscMBALFQb
NA1G7YiMhSUCAfQeT0LWLOPKyiTNMnoF62VzTyojaHvYLz9xYnslbLabS8sIpf7f
MvEGmJTsU8DsdA8/WO2v8jCzTm6J1YDiouf8pAbNZhKQDX/Pd7CyYVHxFh2dLW01
vDZ5HZY9rtUxO3xpIWYAHWIyMnf+9odFCFdJtuR7K/AkbE+Z63dLcVaWtLEOTV3p
jM6jm+OOjmlWdUMUTE6HWp++JEOrJV7oatWbrQ+dnQPhYrRTsU3yfWwn9kQwgn/L
L+9cvDRrCW9T+mSbYcRWLIC2SUhLu7szXX4p1GeLbMmNjhV6zRVYzahA82f7od6n
7e+vhrDSWeAc+JyhS25scMe/Lfl3QjrV28wDLHUpPIjKPNEU+J/9O5BOazu3juEz
pfwdf4y2J9xOnNHxVpeAAGccglfPxJOYwt6HRtmJdYQKHXziVvmpdbe8kbWPt4u4
OOR22l93KJun/0E0ZxR+yzIhAxE4sfp4JlgMv67LlunCDFd7oezTfA5XUUK+i1mf
yj+qCPToOwpw8+Rr+IXI0VxbQo3ylEaJwyLtkqx6sAA7/lRJG+zRY+N1IT/5pF0d
SV7erv5FMPWA/38glVQT3dVCyDe9U2N682Z0tZAwW2G6CU5eWn9r9bATDbnJtTKT
qPTs6FpUr91iK6WjFwwX1J3WBt/bJq48oUzEEPbbz0dgiK54SYzteJo3ML/BEiu9
U5DaAApU+Jilsk4QoP9h5UXU7suLvBaF76LpBJl8yqEX0iSL1bDzCoWKeymHA4od
dBe51HX5xYwyneTkEwsr3CJKI36I0rZlNQcZRYJXmaH14Iq+V2NvvkVqjHgEzDsP
JRh9QR+jUNtGTpnGWvTtldlw/AtS10M2HViAp9iFvdOEvT3lUZmJvEfaz2NyJket
IXs4tMGYpb1P8W1ncpA7pr43Z4X94ycXwpxqh2R1R5zoDyYqNzepPdOwB3b4jheR
kWAn+1B2SSaxLSGrM4N73AkwALWdTfFwv+XzkXL0hS5wUZrRJXN81beN+0BWcxYM
EMw8Z96QBLNre2AFAU6srkP9mZmkfRCUNNA9khRYFdRFOOYbCrjp/HfRRkJBTq8m
qD3rSs/PlQ2YBUtdXKyktlSkhRZ+/S2WzrgEhaI/tYu6HTDmIPy/m9WD1wLMUMNn
MTb1dmU85fiplA8BMjCzJ9rTrn0zn4JPvlHbEXzVa13/ct3ZzwUCZYk7eN9BqdVO
S7NgHcoIfpdW/0H1zgtlv3fPbDbSKBgxvwboRVqJsHE0fuHplOlt/g6FofebH/yu
Vzz7TEd3pBlFrfK3WC9T6VN2fKIMSkUQSovlM8bXB2QkQi8rv1K6aQJ4IA+URzGX
dV8rAAOvehFgaYBQw5iTNbTcbvS7+8l089Y17YK7L0ogSzsaBh4RiXTRHM4VK97A
VlGu3Gi2yNzcQZmytw3zJHKXI9wUZmy3Bl4nwEvT17VCEICcCZDkbVsdpYUnyBAV
Gra7NkO0R2nTONMYtoTOpcfi+lYnGUcVwuWzJhqkdzz5Qrgn7UF7pxhxga2NvksX
bsOXqkFv1RoMAu+YYPTLEO7qQU6ZDoLMiUiqaSeiJjqKyOzhHA0VZXzT5y0abwkR
Swe5saokI6a5+hnwTCYWvgCbTsg5d/QcwUgFAPxBf1iEtAyjHYF7u84uH5WG5bqo
kw1OuYfYoAn7TUK9oGysd3g5fkA3ak4rwu+6ZUye/nbKg2TEXxKstl5FFjIcEey5
0ZRlixDc48iUDe3m4t5eKRjFU2Y9zz9GoydeyfxVN3vEToRRNAUat6R/tzCxJYe8
Vp9ZOInl4pGLwBuompB0VmNb+Rfuf3ylEJrvqs1x/pMi/Z1VLCvjPVLPA1+G0dxZ
h2I/jCPJUejIzOdvKYWTtZR+UHii4bBtybWrxy+H7aLmR7WT2g4+imkoSaASCi2h
n9mNA5+gQzZl0pFlvsRRzTki7jR88++dRaJXrja2Ni58qJ0KD+qaDq9PPeizkK8n
t4+wmlI10JmZ5IG7GmesKMMhBMDbGulG/AgDqvj5SCRtu4kkvzPshtcLtLJ/rJ66
IwsUgtJKW/zsiauqlyLTbI2Czt9ubhVjrAY7z0RUxY5AN7U8vzfo3gUuH5dDhxVk
0OXhRFxTcHhXvvL+oHQ9YZcDk+aBaR9gC1lO+2UjxDOFXU7lZ6VNn0QpLkCtUr37
iChqMEf9JAHdGxWzdDtz2Y+DBMxm/tf4QYM90SFjWYJEH3v+Rmq5rd4X6BMhY9f4
UbXZe2xuwVGbWKV9P8C5IpgkUou1nYdi2huSUiBxa8DpmGA1ZAr2yENnQyAWkO/E
OGVXmPnfggLrOwvxGxWQyMyQsGl7mI7vwOor/Z715tqVNbc44hfEfxhh6EP0TMkS
Tx4uFl9LVYCDUi1XALzBuyGl+KNhXLG6C7AOVrQ94/W0pNLsYC89ZfmZPC8vw81Y
Q0ggoSsOr4Edgr0//V4pZKip6EKQEPJfzKZBlNt42UskVbaBuzFLNc6cSz7UIC1H
6Q03CiwNbOQPe8rL32GZBLUCEksCeuwU4UbavBuvdLOArmmExS7ev7LDwz43wP1B
Tu5ASz/Sln5fxbda1K6aYawyGdtZUt8GosO9vJ4iXx+ZVpX21gKsDqGhfE+M+hX8
R6fHlUT2JyYaNeeEVKreBA3n6rBY0dTzN5zKB+yewbWJialG0jOcPVeHaU2Eojc2
Dhn6HMk0c0+OWvKB7FhBHnm18W+TCBbI6rkerM8i3CiQmf+3slhJzgcJUKT31DKy
q4I3dure7lPoCbgOOTw60kFclQ2EsgAtAT7AaVjem7CBAewk0RsudUXAjE+c/x4n
eM4voTzPPU6Xk/rB7WvJZ6IUQJi/mC/n5OwtLXTZ8pCBtHcVILB1pivJB+mg9B1v
riinVhjqS6YjGDjhy0/9X0aJnLol3vrz4dYpX1qJ5GPEaHuJo3Li/AadYICOq3Lv
099rWoa+ncgVUrqYIczEQlFv2j1vOQy9/2jvq+u8LpJ4nsLkf1pwvGcTU8N0Gmz3
8PIrnG1aUOr0YyNevgLavUOAeyBNPrunholpetdALbZdg9HjJB9+FaQhYWLQQcha
ajB62ulB4qUsqi5V3XQwkOTJX5ovoydXO9L3I35KJt9AQsUVUL0cnqHaO13uiZPK
iu6ym0+sMm20neTSVYxRML5lJVkpaYR2kHbi7GBydfwldm1E6ntYrYQygxqNT3uU
Jh08qNcMeMXIPDzL5BlkL1PZ+2OSHFSV7EzKKAqX9lHbHPv9u3Mb9CQTyUq1/mfl
3rWuxwfJxY9xvS87mc9SM9m6zryaq6tPhOkYB12YdoWp4aWZxqOk83UE4kmA8uZB
PDKn0p2eriMMAOt1eI+4dDDH3/jWQCFDD0dZj3FqJqHSkSyVXGBeETRMLA1c4vg+
3Ld7rwp2VtzyFwIwNesiOzzU+sxDXz94GXqTZmnRLlxqZ5YtGlz75mZNEUOai3b4
1HPLiONSsrduQpjRaTjIJhaxcKeX9AIUdnSNYOtxUwOygXYjfZmMUG5KzhHgF6c5
v1upYs2cu/ODOxLXug8OBXeJ60X4xn0Ek0HvFRXoIFSRgkV5esWdd2BnXP73oazi
hlB1Jj2f2ICo0anj3P6+AjzipruGmIVDtsB/nIS7RAILhO2XiVghGqaq7J5ClEIK
oNZt0d2vjITIS+YTjEi3SPczh1ZPUyhXSnLShr/oQJimKrpUFjjnp1ysqB+QRFv+
QOfz3zeRfijGjppeY3cFHiLaBOfsXDZrGbHUT2nwxUdBzBDiZqdIdzKTPHrJJAkD
fDj+ZXpeHZpGNU+Dx8hF957CxlhD5+9JCvWml/5fIm9Jc5JjMcU5tI3/MZ8EXWuq
r53pwK+E5aqmfs1vJTC0op5gsbTWpVss9uVW3ErZg3o4m3raYOGAkVBRCJ1bkNGJ
V4Z+xYoMpz3fHKEW8Da5w5Pjwe1doLpfFCF9CXBjerRpEFRMCAEjL1ND2yQzFgDv
0aD9AHZKeLyp4QKTL7NXB3RVlnYNBzr3oeFEYx3rwmmo4YUVKMRz44vuUrGK64Xk
UnuFkENQ4hdhHZJALGWp2/sEqCW3EBKpsugxos2eOTeHJloWo+TBTTs2VXqTuKuB
Z1B0VNXxyobvTa2ML0h73CDUl72WY8kd+fCkiknNVIo+/fwTksqxDfHXOWmgVgNm
LXSZ8R5+GulcG4Vt69RNyNYM2rTpC6Q7lk+V+5Tt9f4squf1GmGP96O4fH/wTOEQ
h8uDVeOE49I3FQhDupDGgvQW0aRFBdPzhlpzQreSA9Ocn3MMROLYmRqXB1kMaH7W
kqWDYCCXqqCV7PLsuxCp312w2PJI1lgS+WIc2HnmiqoNkavCPlKpKXuUzqydIj5u
XxYddv3XZTohO3gdNbe1Qn2dCxVa7NZRtaHZ0u+uEtMNqcHfwLFG2TD3gZ37AfYv
FmmDbOKYFnNn7O80aIRsymx46+4+6qYEfhWVc374FVqN3gFFZMKXVdvFZCFY171G
rglMDjBE55VKLcGWHfvqRB917VfJzf7cjEAtWei7jIDf7q6RYDC6j09MUJivGG1y
5u0jeIJmU/L8lOlBLourwzkvgWf8hZD57JQ1efJmj7iX7ibnpj8kWqv//UqjU9na
uC8IUovLQaGXixg7eIhKmqmrrR4ZCwHzqI3h9AvAfdI3EQWFS63Or5pnEhk7OHzd
JXGZ/1pC1BJDmG2x949mnIRHtbRxNB7yAU4jOg/OqIn3C7JdhUc3yXAr/RuMOtEm
czX8F8uV3msfGRtLxyioE8a5/J9//Dp5GP5DSRwXrvQE9WtO4LVvsLvTbRmMQFw0
inrrUQA2wrqMA3dKR5k2sww+WIPCJ6vP2upeFKdLBAEBlrWStMf0Gek1sqCk40SG
jITJvp7yd2YkE8lo+NDzrriuPbYCQYIrSvBVYSrYR22fWQCWJMhXKE7fiMoJCUG/
qkYutax+B2FlPx+bqN1W8CcyB4Fzk0nWhF3V+czUKgS9W/vzXJikbIx1kTSbWS2o
mAALjc9A43cd5LPs5ONnOqJKprtQQ5qSvY3JmME8nw082fPb3YkOkOvtF30mK8wl
2UDJm7NPSdZD71u+866OUS5Av5pcexH65L43EtMF519C75R40Ki7xCB4u3IHm4CZ
y0x78HEdXyhmfhCfN2bLfQqIxK6YdPFzt9HYNvgWLQxAMMQTojsPl01+szFNDqOk
TULeONcnzagrshiTsnt9O5OcAY2XiL+8tzcQCZ2GGXYyXLQ/munXtoMB1XVdw1H9
o/0YSR3sL2wzFhQrYHE71XQxAWKpFcKNo0c19dhdRdonToS/Te0vX36ub1rMDRj6
3UCgY+fU7v3oLADKzIStaD13ML5FYXTS8JAs8dAMgFilPuce1vuMC1YQJtxl/BuZ
xd/FvrL070sgzRmOyWf2AkH8iTr3mP4snJWWLCbnhulC1cfASf7H3icnU+iLlmGK
FvbOLYObwFi/6DeQpLwV8j0XsrL7V6SeiOUlKM7qnpi/fGsKwrMRqvgsZ8CPsXdZ
PqhWYO5vYtE1qN8IrmI6GtzdEJ/msZz90umSz+uEXOa/HmX7oiYHa1wUBxGjaaxe
Xp1T/XpGfGb122WkDJ8sa/xFp1+VQWZBzCPrjJpz89nkukbUeqq3eyS1yvKudihQ
jXpIXrQWDPBPOZKqRUXIcwZXF2WhNWjqkyUr6aQt3h2NEbT4mKcFm/PY4ikZq7eD
ALeppKj9hsGa+rtkpWFiCRr5pFfmSol5yyiDrh2h6DTHMGeyZbNEjDzVHro07d0e
JL+I2S/HNAuaLPUGJbt6V2bbYk4qA+/z8V3W7WfZau/cD1ujbfCjlQ3hQ/ArDqJK
S50HirzFiVzWITcpcc1Jk9YlU5rtIRwQWVgIoeBrmvSTMb3WCVZiP6tLIBEzg1FG
1k1nTUGSz4STLuvXDugCxsH3dzHinogfRMY+gbgIKetIm8aB9g9D14/7l0mGxG/5
9FNLpRmMttXvmrXF0QfhoyYLPoiRp8J+6JfI+vyFrDDa2AHtO29BcYjJW8VK8V7+
ldCxVVvlUbOmHw7KsX2txwUrbjfpf8n5lMrNNoqG9CGRLyU7tDxGYkE6oc5jj2cu
y+Rsqz8f4U8ptsfKh2t2Z1aCIR8QwxJ+cnnZ1cM3/WsxdKfhnJobnq8SsFtfYDzN
QnuSXlchXimCIz6r3prSnkySNYTk3w2OKmC+TUuZMp7RRa+1u2/YAeNwI6JOuvBK
wiOGxVhlJAChZuw36fZnPJpwqhjjZm0oGkZEuGhWDCxhAyUepa8LnZJWbURsozz0
hlfK+c23EO1qHQNQCxaRZnZuxfdTMjc54ZtPf2aAT1P/B442zsHuo6WE8DMOSAeY
KAxF2YNl3psLlsMZ3iFtkcJuiXIiEoIuqpeYVAR7Db4ct2HgAGtxw/OmcfABKWdg
TqXa0BVTXc+NgLLmtYs4mN7JVSfXnVJ500CZVtjIhcInCniVUa3cdOxlhtrOEUSe
13krLCPePkMjy3IRkZ38EUPX3RGzsbaBXMPyvnhPhsep7L+GffGP4N0ea0l8KGdV
ogKpqOtg8OP8nRHrBIXLNt46Q5zwmvNo+pD43HaKEAzfoPiC4vF+TZQPejmcJe/9
ypUXlrzT4N8YEbmLWjCY65U+EIUq53k0QVUFvsyccDbK9y95osjE9+G1R4yqO4lG
USsvQpJbqx4BAlepl34214qiJHntbToSi3Oc3IYzFZcJqFa0l+GyRXstP+JKDc8z
IS3hEdmzCd/LM+qE1UtB5KVuDqxx8jIztLIk800U3eZqXT7NUN+kIH8Q0uKeZMcK
RyJ0i5ui8/8uBG3gTMFU0Kn9RJtR1slQZbJGyPR14m/5Q/L0qTeHtu4WoM6HlG7i
sY/072upYESU/eBrdpc7td9o+hItkQsWCimWoC7e3f2M93Up3vP5rwbxpILdX/iX
5J1dODe8EqY+zoAPRtIuASX8j7faQCCcuRZEiBKs4jp6e6l2fVq2THArMWXMBVK8
UlmWP6A1BHv3wAul170n0WUxhl1WuM8hN1Qjqc1kaiI8bhXzZiJzmscNEQIKHPGd
vqjK+S0UrF1Qyr705PAL7lhY+Qa5K1jhpu+hNQThLXGxvi9H6FeVlIYJDRJ9EKbv
tzDKYzlQutTeampRESfSxh4jIPNmhWqVcLoTEEkcsNmGB4RzOkNL78eraEo0HfpB
sXPt4YwTN4wZE1J/8UnAQEM3S1NpKX20JLK1ZXO8S05b6Ju5b7ICdnJ0j0pf4C0E
xgXYAbDIRhl0Cif/ZqQhPQvJarJM/gOzjQnFhqMuD8BC2eE3HT7vAeUjw4jDLeNa
141W6YjOfZIEUwQXMd+Atq/jV9Fb6bRacYLo3FTbGkoUuPSxvOba1NehhPUPJKpA
jn0BLCrycTNXCE7XNIdA9xlXp/XjpEJnFO4yIljx7vVmBLlPRmYYTOFugCqj+nRw
z+4rL8hsPuzcGJlByX1Ht0deT6R1qwuBnLWZNAyDIdz0zEZdn5VUSdTnGgI/8cuC
NKx5PGpDsIb78HyDr4PLS3ZNluK5hLjcqgpsGuCCnihIgvOhOJ3d5wHEb+X9L+xY
skDsrV9kBCyZt0VDX0D+Abu49C5iIqZiVavHiM8bToH7nmxCLesFDTAuUg+/KmT3
AF6lWRalzsg19r/aHKXGLkzJpKW+QAn2z8C0zrLUQr+ndJyqBETV7JIRvM4p7ToA
tSS4nh8OCcw3rpeFEgv8RWDCH3Tt+I8WgZp49ilVM7AddZVCCiyQR3ImTcp8Ta1U
U0sC1hph3g5qOlUFsUQ5QMz0fOhwZjIqm1AmBwbNDqRxg9M8NdtKu1Js7XF27vUW
eD77lfSJhlwRucx5nf3J3trTJXGBl7xUp1hzh7Hh4UT8FZ7mIqqnueYrF0oKKCxM
0CZ9KHcDo0i2QT5pWfL0QQCivDUr5MciQukoeQ7aziUfq02JHY28k6fPFEQ+3Lx1
5BQDhvLwUhBe5qTsPK4SkPnab0gkhZnbZ97YRPBLkPiwuRSUX1BEkEpFkh9quspi
DI64G4YPc3EtUsz8jGyTNDBOq0CtwrE9MgaKSxcpQ5oAwvcTN4xLLbcDFIyoZLtt
gSr7br5vSbKUJJ5WWOpQDVcKNjX+CyfLKz2qb0uCmP4VohgOh+CV12VD2EmzTHql
e0AE+WHziRwo8gdAF6itgaTaFoLuAXY4RLRON53238L/uyjQQLqYJJWkdFrG2C5p
0OZuF/iPUmQm3JYE/WppdO+PLQJyMjAzBTBZOR658RcQ8qVVAHUrojfPp0J3q2Sh
uv/sZ7wxyHS4XT0L0orLfShqnTuJvBlIJRjWoOaX1+UvS5NgpX8ZOQ8EP9O4JbOe
uL0qvfBjNn1PjPTJ75K+c6/RBLslSEXs+HHYDlJr3t31MD1m/ni5fDrA4SiwOfIn
R566Apj53404nmUA7NViHsiF0TmDlnAl2jD8ACaneaWRdFxpzsD58JUbUsIa1W8g
UGulssNGFm+Rc2zdU1/8Hl8+F6pRCVloVPeMbwGwjVwxxu/VQT2V4r5zx4ZDCz3G
7lsACHK1EHFWkcUcfJrA+6ny61Osk3xofKBcgZ62i9YZkyMoDxkc56xfSsinQZmD
/ZbTQ1gKPP4WXrQQK1NxfEZH7yyDLsJEltxSR+drCv8KgFXSLRCeIin+VJ1xs2sh
Nnpg8xuY+NL5e8Hj7APDSnqlPVNnN8M5u5TWX8B20epD7JBCyGtOpKklQZqp0mWO
FccNQwwzU6/gzGcBz2rSdZ0MD3Ck5np8Zq+h+FhdQzsbvDSZwRF4wxFZ7Uo9xEbG
T4gpvfFQn9zLtnjEdwAe9Yu96INKMzvpL8mxWfTOCLHE/hSQyui4GxMoq5WmAyyx
IO6VIUsGr2w9NExr41z6f/OahzwJljbcz/0/9bV1kKHsyfJmlet7d8gaXay3EzAR
3/dYlnxO5Bx4QJlffvh4m5CanG5KsVrVYTx2qmsw5mhIV1Lg7dB3RpKCMy3c8Rqj
XK4hyPcjW0AmT0csY/oYyIM5OIwKQfwzdtosdXG8wBHiA5PTBQF04uYkThl/2dEc
hshUiAuTBdsuMzomIa8U09TobaIPuFnvPkR5WEa+OMhYbkQyOLXsuZghlcUsqqOI
2PA4O0D6n6TFtqnN6TaenOBcM6OTNwNAwKV2ulbhD4cvQT256HrsCYXBeIWaufq/
qZCA4g1ffHj9QbvD2v3UsjZTUUbUVIo5QGG/+lYpxfmrrqfKB34cUxys/tEEUL0R
8I64s0HX0sKxS2AFpMoTQBesm6L5eGThkE1MjjU4zxq6Ce/YgL4xvTbIUa2d6V18
hPxoJ2N+e+aijA4N4uT+z++F7ye16wqirBRtS9zEryUR0kln6IMNRF6RWhEA0ovW
zWmv8nWatqZG/HPFwu6prBIQsVvxSSBu7NSihqM42X4kyousN6Fy5atlsZYV4t68
xakMxmONBRHO/cR+La3EKNhiU3jBMS9ko2GM8B14CAgKj52n5wwQ49ITNMSZJVy6
ujZcK1/smU8eDdFdZ1a2uQFy5UKWNd8hAuiOx6tJ373bJCLG5KaM5GrKumBnMi9h
jvR4b39rFehtuSQ0JpQi01IWAuIdROpVukiZdYJdeowmxUZ0qFu8WEB76lLqm9lP
xrfYShdeDOVRS6NeKxEhkPV+CDZGj4jD5NfoNPeW/9AP0+szY48r24fAYLwMhljP
SwAJV+TLlIxTHpWrrfy0CPef8qKtMgIwUtiZ21hYit0ZRvXXInsmQyRUYndiLUZJ
Ty0V1gFz0ahbJY6BdZaIA8UZl+2turv9+ZOzsFseD18gVuGjJh8izil28eExG57r
R/0+JIrqPQ+OHTXNaXv4fbzWAc1e3gNPGwsUaTYdgDYtDTvUXIrmIF01ArwllBgV
rVLUx8X7QRd8E1/J5X1ITVg0Kx3LkDC4OVgQUkhwKaEVfsrO5HkjmWdU6KOYRsEJ
05464GsXMKnCj1RCz/exgwBIzQbCSo4cL1VfTa6/UOnMd/l60VJpIGObRiM3UPIj
MBGQOFLQedSWPk3RoTyEs8aIPQ6a0z5g6eFstKKVs1hiq7mbFrp1zy7aq1DNfvU6
ubX3eN1OTxxH0kCLKATQtAN32/88y7ms52Np1p+kWEa8ejvM7+4fi4PZARJjxlg5
ekE3qum/23pvbTVwc73W6XaZZOhxV+qJID8kJdiXKUH80glun2K7Lxx+oqELj/4l
/ojrHngSKZQ66lfSL8WioXzjO0U+KkXHUZ8eAR8HX1+83rvxqeEgaiTbT6MZOs0/
EOv6d+HZGO7H8w0rYz5pjglVcSEhd+Yfre/RclwdCcduYik4zjBDJPUhP56CN5mR
VwqG+w8Rvjir+RpsANg/TQwPF21rSmnJYhlu0TcUkAI8nM2IKQSilGnoi04SPEAq
iCVVx+/60XyPdw9d/MGXDG/FQrc1qpCNHcncYmqhyJQm9AKbjPwsiK4dChxvMBUO
mpOtzaIy2Vok76UI282aMVjiaxNJhrFxiW7k/NJnqCpkz3lrmJGdrj7l2gRuY+QS
C2fgnUyCLQSHpdPMC4IdBEkvE6sJdTZ0dW7gFTbtGLXHIYiNUpA3VRWclFyWdP6M
FHmaAiSEv7+naXliBITd4n5mC/UHAKqBPKBkh47QSsx33JyEy/w7UMez5gyEdN+Q
YbM+QIQnuuQWuYm4pyGFS3hXepBpy2bna7Ly70YgvCqPLWSOjvv/DArk5q9tZQ04
joSQ5ZHs16YGpypGTjsOf+0OgJs4klJRTxRDzhqQRSkm4YvGRVQ45G7iqqUkNz+W
sSGNsduFrfOhO5DX4St7mQR+azjpH9xw2cN0ZvnwtCIZm2Rgt/dfztHe8uLxSYdA
hWQrMjRan6iwXwqB/nlZ5myw11XX/WUchTzEI4UaUayYX4BRL+wPqmo7uQPNlOo2
ElRidmHSq75do879pdB4QieqS7EUq4yS5rGrEjv03UIVpuJtx1rWJoJnJ8Vt7Hfg
diaCO8sDdl6Tb3h1a+TM1QUbUgO2oKomGQvQTBU7trXOBvZKdu9irlLAz1FS0zvw
1IZi8VvBOfTRHGwYNJG4gZNd+NBLJacby7L9NUmrqDZ4K16xbcF2Ci+txdgToklm
XD+JQl28SNfOV4ZdtYJtj19TDCpHwdzVretd6tX4wP/Eh2EZdxJGhoXuJOliHubF
AdRfXAI48BPF4yG01KlEykJXFDOKVEY5T1aCKCUkcql0s9JShjj1y4Rf5EWPEiSP
HYAqkCW0hLRYeFyj5Hkg74gjTJw7HTlydYO7BWHgtioIwvDDgf/4ZybUdf94OWR8
9pj8J+E9/DPFpbfGHKI+EfklQmuY/gk7yNq0uF+iJ88UC/WbnvBmoP6GdeSCBQGw
9znB/7ukoJrhMh2gIqPBKPIEx9Uzw1EtznMCVSIEix3QIpRIJmC6vNeBVZbB3wwx
OjBe7PZqcRMqkdTCBqy6oLqrEp+rxflVfW+tkZufhWtCJVbiQKOWDxEDY6ifBklg
BV92N0LTJYmU1qDnZ+CaJKWkRoJjt0rBXjweYyDZGf+3Mr4H2xbUUide/xOFPLjN
s+yMKsJIkhman9VqCE1bdC6PlFlbW1roZbaVoo8HD1balgse5aFjmPKWuhRirqYK
k+IPyWvaSHyBKUlrQgVReYRhWPhY2D3KKSJF9dD5mxl9n+2Cx8kVN5eUn/MQKNBF
aV7syCLM/dfTukfJc6hOmP8vgYnaax5vt2Bj4Hnjdxi6wfMtFBdlUkz7rjpmcgfT
llUSxi2yyUE/lURB0kIQ5bkvy7XheJba48e8ro2a7cMIMLpWVxCi6Dp6yjY56m4S
VdbvIT5OA2QtiK0Il4PnzAZJOxAyYIlD1E3UtTrfr1/ciHoTzaG+T/jjivkqaMxn
+xjg0hqS8H1RpzvNE7m6k0DojDphbO5v+lpRO+7qYfoxa2+ho2kLWw/zIlYxPfUo
W8cyh6MfTlHp3IxIG8dlN0+QnxxXRndoHdXbkGxEwam8IwZOMr27XPiEONd0eVE2
MEPfezGtpVq9HqNH2Ky3b3tgfBHN8EhBikiUzL7CiVUOG5SNQp2fYUROYxD2vfBW
7uVTesjCJ8G0LPEGMieCvRGAt4AIddA13F5g42X8W9kJPruApkcs9Yl29CA0iHE8
f1XZsQdnAGi536Mqmpsixanputwry9wWSxHY5fmisMY=
`pragma protect end_protected
