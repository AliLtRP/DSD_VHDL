// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:25 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UXjsHKgEcP1UkjiYEZ9hOiXqqUN0facxFAVqfudkrELV9DYhHzf7PFobWuW1cnz9
7WOUwiILk3G6AmlL9nKlLNGu41U68+3+M8DbPviPbZ1dEKIrHDPzQUJR7ygPw1Kv
Mxi3h9tmtVh3QW5qSmeAGUuubwlb0RyoodP5CfaUB8Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9840)
hfyDK7wJk63KvSMfNtMwWSLo8f2slGxae/LKzq2+6IxhVFDeiU2TifQx0zWq2jIl
OMGZRTgYNtQJBcuzSnyHGeJlX/OC2ApLGxc5v5gh4xryNCBTRdyccQV6AiJg8jS7
0TK2uJMgGNGV0wPxler6tpQ3f2K771ahczWzym02YlW3UqkvFrTvJcYNy2IOG8zk
UGhdMWwIQKzCEmcIUhSrh4RZDdJ8R7XJpF8nYuYlM1nG/3t9JmcrIOVH6mSzelld
24QPNShe7HePs4JCFXWCSuK1QvPWzxJOhYlw/voyECPjgRatZCUY/EYfLas8yBsf
GnWL1+83Ub/d9CTVRFAY9zIUbWS0R61vKvEEzc5/IPHYarKB1cb1mJAZ+kuNNcIF
eCmmErKmb6KM1T863g+tkzQhSjMzUDuhVl2on81/TAtnvMzKdixw+cwiwY7AAuCM
caBChn+X1qRXk85vQYQmH+uqNTMK9DwUMyzEyL3l1tgLGFvA2B1z/hWbOCH3E+Xh
M839YjRk09MnuDDef0INIfqqrhvZeLGFDNvr+TUhfFneNh91XUCGDfW1NVui6p97
dRcbgQIHxj38CGU5uwn7dU/0q1E0dKVPvE3lwP14TfuupHhEMOQ4ads0Kj/fdCrw
B06WzYLzup6u7I6SQVKGNWvA69XY93xRydqvv8lbQBQ7VqwcRuNrzjnVHGqgopoa
La7USJmBD57i9maHnigrYJz7pxAbRop913E6V96hiiML+amjyx5sJM+n+YpM8SJO
FGbG2Rqvat/NyOmLtbbh4WdauYrTclOio5ioTE3FZphGWiw1cWNfChHPj88FKeLx
Ejf0411pQmdE49kPRYImJhdv7iVYrsm6lnFjplLyLISIf8KKRhffqFvxN9mBRJVn
yKrmNyCU05krlAZRWa5SrleVRqvwDkcelKiSMWlZYpBChFndvPNPlTBmgN9Ces75
f6n3scJDGGqHEo2OY8bVMaO8muHpX2CKNKy04NOxa4bJ5Hl9mKVxVRwSyVJStcxJ
BIZyd5PRKfX3GbDTC5I1Y5AG5CLNJFU4qyGHFHpDJhu9OH8/e6VZrGId4sdRbco9
uoIW0ppDmxH30SkjRuUK8vOCqpr0LRGU815Fcw09AON6DY2wq0aEcRY39cl6OXeh
pfxcTLG2ECGbycK2cQoeYjsuYIdn0Yt7W+JiwQC1igEkF03rdfcOE6yEvifDs3wx
SLmg4jU36+TWjgKkmGQwJA7LnIDrGeR/hBiHcB9DHXWEHaV68xfeeex51WNB20NB
+z1/lcsktVgFmqxWrPHnbukIMDyVovs656LoegEVLghTUQ2aQap/MQ3+iEfFX4iP
5m7xmY5e81MXI+DY/BdrGtLqxtN02qq0la24jqW3TTFvW3vGOP6rlpgrJ51Jqzf+
1IsNedb0Q7ha5leLWTaD4vOUOUAGI/2Mj2qwqud98hta22zn+bUGJlDqqDQsgp9p
UISwKuH/7qtUpZJWwOlnRLv54wd+155yKTIjfqOra2wyIsHX0e7J3Pw4V2G+H6gz
ukageTeZbBAlRWOV95K2PndBy/vmrwaEE9IZXKfDaW/ZEwMD6QvxK82KcRtSSB0E
f44ffDnvGgFqGlDv6K0wHuwGeCDQWvUnc4LWW+sDufErIs8UF0ikhDFo//qvl8T6
MyeZM3uiU6MpI/oSwrRMuzQn64OcNt2hVPU6NpCZmQHiIVIxalGRD9DIyqvlS+C8
rfGsZUSOjjJuOoJzImWTbz46kbowJPvdFshbo69DhkKv8RLK+9O43lJpo02Mld6k
E6LhxFhjelSYTG+E0zsZ3tePRqjIOyv9WGUQwf+ZGjgYWs3gqb1tPgElJAaksWbV
fLwd1v1KVltxxON0XI00XYQ/QDdz4VfbmUCo+Sp9LilhRYAY7zLcZz3Y5L7C1RaI
14LdUvi3k6ogErNYahvhHAKEBc7UJC1MQVWWFplZoFADsk1YzOJy83LEduCwB/LT
AoevdM5m8x1clDJFYlXkdO89T5mFW2PW2/2CRTNDRTfT/Stgbpb3K5nND4ij06H+
bs+M02c3ZxiKI9g8R4rDEZQZ4Ia8iSg+TR8Tv75y1JvVZbrOnN/pTzHvpxQ6Y7sC
w/A3mj/AF6kKpHyQXYjJz+gmjKZQ8SjgCnEnxDNroFBykWyFGKugHHOnrWsmGrqa
uOJS0vDjVK2XfpwJ/4t1iPfvajes8yjrpLClWDoQo5gzxUzwUqjpCexZMZYiPUq9
PeOaJgbZCleqdSMvsjlptinW5KM1vnXTHn+UsQ2nAHfDzyURCSaEW3jYgZHavqP4
0u1VyIYVgqplIeyxFx31Hrv7+qNQNpADqBoyaG46SgV2zkMe55EipZjp1ifTLJNE
Zt4qGl5mRWD/4AM52Ia2xRFPxZ7v9VxXKz+zFaKhFE4Ouq0OzOgtrodSNNGJICzS
KnmZR7WjJacNwIxUNtYg47cXJvI0leaQ/dTkSyjn5dIJxoJfylYwLEVOx0V2Q9Hi
DJ0vxEpMGMmzIQjUJu/DBxCRmhoGnyLGan3HPj/JxbtjxBkUuveHXro3X+p0vuAw
g0d3LdJKy/98SzpRy/8AylsVOX/6mhSQqnJ8NFTZ2lUSKBikpvL2mjhxS0Ho5bIZ
UvpGH4c3OTd8UikSysXyh7anUowPia/NStnPQkV2ZvvFBvNyW1HMjuUBytMlJI1L
xelplUZJY8IvJ7b0+QqDs4RGB6Ic79fhVILduxvfepmqInj1Os4lNzwSenyo+cYM
wI+4GddGc+RAsCxSKwBCYoMRn2pT7/eZ6LGAoc2EDzosGfKBqTLXiAdirGl2m1mF
2BIuU6u63k0XmzoQ5wycR2ob4qXSF2hc51OIuUIfUJfQjEucylyX+2kj1u/7DBUu
k+FZmze94XkxtycWcBU8+nXqDbBWReM3y/WnNoZRNK+GJPBE8ypbe91iRyr4QNYl
1LcJNKVQusg23MhI9qMoY5p01w+gkexrYWqOFfghLYD/fozhbSIx0WUOnD4xhohl
9V2k1foUfFYsFdqh5b+OqLZe56BgmGinEQ/HfARthHre1SF/03W2GGzxRI7ty4EB
ho7Y1x1xfHwgcmMiqP3H5kUJGoXsBVeMpEzXzMiRAkGhzbuSF4SCvKgwRWlZ81qF
ZW6DF7wNhuOYj+aIM3i2jxgu81+i1+mIdaP+doXFOCbII4JfL/1MdyFYvxpAI6bY
ITi3gbu3bujAR6vSx+Ue+WgRhxMvQ0FB6O86WoZyYy9NLjUbBoQ/13COXxAN9S/d
YYUrOqyvPGl+utjhpWxbdWiNAok0HP5m6drZPQ+xrsL92SnvRNlCTSwZBMmCu7ko
qSgAHHPYEpZ9K7TsrFw4GDXeJkdqTm2/PdPjA656SCJVIJ3i7lDA63FM3J+n5lXd
vrP/3lTYq254VeNnmlUFHIHP2dmdhvIVJfos3Bfl8d0qWtEKqTYAG0gcKrOL1m+m
nZzHAFwN1PJ8L6aqnlm5g+um+j+C/g0VXuzPpNB0HrW6NJxqMKlEZnseA5sGdXg0
lgZS8dk6vULt3JmwDRY/tKsRJ2sPC4FEsRVep+Q9OrhPRJHOmkDAIgFS3g1sSVN4
WzlwhILykP62D5As+uENjrUSTZ7oSyOMpBN8YGiPfAIUL5zfivNhM+fJgusNBifD
v4SCAME2B5kYmkUGdSTeOBAeJD1EiVER90YEF46sSJHnSDqKGbZGpGYG9W6/f8TE
YJ2GG6afp5Yj42mSBpuOGI9eCUfAB85zLqcNunFfEY4DLFLopnfyRIqocERknyIV
QvLoWH9HvJqYsQx+kCRxN4IZtRVx4DsA1Z+d9jRMQu0jdyJjcRYIzRzpBHcXKBqm
W1Oft7mYQfFl+qE7/n5G34I+wwFnV13sK7FL+RDnIBF9nFRZVdg3RlIPZVnUUpAX
lIcNZ+HniVja/N4Kd3+F0h4I5jWGNh6JllCNlhaLZ9TxTBCT7JHdCO48qcTn4X7A
x+NcNh6FW0ZEzCoyqEnzurnxPhZ7z3RgSX3PlUOmRayhqAz93xCAwsNK1e9sk+U8
2BEFQuR/B1vKLLg2Lr1zRZgASTP+SbnNgA5oUPg599YVAk5WU8owbrxx91vx//0c
m6BbNQ8+jxEBZQehaigm2FgJtMIIriVVQ2gMiRUEYsX1fdV0+kyAoIy0SSd4rD50
RPOboMJCaDSmwN9HaH3CCins/rSDp0Ph2E9O89o0W630iPst1itIaWkGRkuMyEqR
9JQ+P2+I1TjK0LhftNz06D5rhoh5t4iBA9vI6nYGg7oVXUnnfbjbdP/J86lB5EP6
dOX2iBPZ6lz6x7d6tPKf4zIf7iHGrIJ+Kh0KHEKkJXVjq5+gswnaEVkmh4mc9f26
uBRhAdhL/sq6aGTzaLesqjxnyBeUOyZr+wQT7iB4nrV3V7xQ4vV69QyReKa9E0VQ
haTqikvBhQGueTUoIGRYkNyP53cg9jfuFEAyTSpwSlv/ujxyCHoxqjX1NDUhTsTq
p9HvpHRKcwSW3FpUDkwjA1wFMU47kXEYEyYsD/Zw2pdyjLvuwulTYgBWo4Vr4G58
h/6xafRyijTrfOTUzU3mDBC9k/3gOUIEIbB9pek8mlN0Y3V+mRMgQvWS7uOh4G/X
YxLs3FM+Meb/3aUWnceruqMOqGvhr+KNCDz5RkrJd+m7booTM6S1n407De0IFJ8F
ThFoFBIIUJ4gByUUM+axXtoxoUpWRVELur3HRR9ebASGC5Ly1r3/umwoXWxgMmrK
UJSm2Fvfu9Cb6xnPChI2kxnNoKDD1syq5zZWqVjJ5DYC/4QAvvsDtAUjr6Zq9Msx
VVozn8MavuH+N2uu+a9l8/WKAxNWiYw3MgqpStE711OSiW2OVrzWkeDU3Iv39eOT
za3bFy+8gHA3BODnmyIkhxtJyuFo7lNvov6NCcD+t2wycZeMhD2xuAnnuC9RZX+H
mcA/UT2YxHI7K13MCmbT+k7BrB502ZKQTOD2gpZsY3PcYBuyscaEt4GJaniJHb8y
ZeSiYJHJD389go15uExDaVDLzlQKKziY+4uJVckFEpMrbYWGdAtecZ5DmerNvgQM
5n8KtIbHYTWS8bu1W2jDCPfJ0bBkIRuWE1Y9nLhND58ubWs0jgPpQiKYGnkXrryR
3IW0NN1AEG8341jqmA0/ZvfTvCVSpXTBv62MJrJWad0xqHfF7CK02a0GBbpXj3j6
iZdKy7FOF+OZ3l6ww9K7LDYDOLg/i9ayL710xPxkOfjPfUCYkfXuyxcY2e4iN8IW
kyozjnPrQs9udcEL768sV1a2jbKUx0GtJlo2u2YQmN/Qtbzy1xe1Ee27mixUT6mo
2bC5v6Ap3ZAW9jzovCftfZpcVpxTH5qxSfQdqc45KInIr+ryNGFYfGNleirAmGk8
c3FIEHy7Vg6xyzv9W7i7R5uJRGwBX+gU3g+mRQBvJp7YuZRz91YyhEZsrqv4xYqS
FPiO8V5ORHbiLrFF5Xv7a5TMy2AEEuDnhbjBdjWNijhr8VcalFeMAB9ow6vut3Uv
oeZWVvE7oqdZlN3AH/iyG5PRMuqpCdGuJD4FjV7B3TCHgXL/QB6+hQCgm/BniIBm
gilq9SO/mG8coG/1b1wdOscm+gvMyadV2osIG4ixz5Pvxe3KxTMCRN1sFK5U4ZBI
y4K451/swKyHRVB1B8X/VKDWk9OuX/Ue4CuEXvFMALyw8me+tTb4Q9YPmeP+NXm6
3mXzxHI55mCf+IRnL/Uk+wYb86QuSgWn/uTw5g1NoKbnZTx9vR+edOz9L23HmMLl
k4amdZ/r22rgQFPEmE335Z33wyCWpGlddQajOGQ5LPvT5UYohHN7BexRWCEsRyJt
bCsbnvR3aFVoxOhuTPPR+9i6wLqsFCkU7h9JlPYMHMlw0EZVivROWwQwbBByLOus
WslEIGwegbEBjLHzP1K4jKe1OvwOnOWnd/fVDWv3FnNA+BSRDlN0JKrILpQ/9tjw
2Q+Dn5vWfE4pzcgMT9aW17rSsy7iIjIEbel9BatqJBumRTr5HXB6ACqLpxnEyofT
8TfOYLtEcE7XE2Ivx91Qo/+FgQjkUmdcnjeW9kkFp5rC/v+8hnHPQzryDH9oBPbz
6yTGzfpHwwDWwZKC2rT2Q+pz9cKZc11QG3SBVExoII8yQoZHS/2tVbx41OL4mkx5
TkLWQgRWmtxjPO3hGNsTYVQk4vY7WZdmXsxRGbssbZFJDeRinv0e8dL4ZKKy8ul7
SgmsxUaBYtz5p/ZUl0L/R5hydbcSGgUo4QmZe5fnRZgXuUQ0EjBNB5RfEEUFKsU1
2u6EMJ27PqxWcCNCSYKAMF1h/dSW72SDP3Fvbx7BAQSYAY3DEyHX/C29/GpSkkig
6GFxyqo7rNMHtOt9p02UpB9Qnm3p8KR3p6OabTX/ur/+xXUbcWFtH/TjzfKSHdu0
u8n1frjfCEWdSyn9bqwNY+gjtAvJuubck5mG9VKAkJ9Qn+R4hypbgCWDjqTlMKWY
OwvJYk7xFZZ0tq3kBODqc/98HzvVQpuByY9pkQhKTMWavA7fXNGwRqFWOv1Y5jd1
fu3AQ52Wfsha8EMA+NAV5TsyECYIpzPwfOMBxv0dmS5JHq6XSuA+0GU0xdzvyYhY
//8CzwMMO5X+/dQBHjCDVBp6WImh24HhjTTrSC9fWiCtersNRLfCa/EoEMfOa4rr
sLxjbbN7uNDqEgMcgcVSlqGjrgjEer/QMpQx+b35zALfIKVWz0ijrivSEQuPv7eK
glj0kr31ANEVdmyHXE2gQn9/xPfWGLwnDY5VAOLb5Dm35dArXZDIvHvcpkt6kOSY
NY2UPeCQOd4d7i3nFsE+meS5qRF6WCCphBhJjbMve20P4O3zfXvmTKP0aHUS2UXw
2g9JIc9Aa0nlC+FycXJgNBr8UCp6p7I00UQyV1SUkGnWBapi1RPzQC3lWMcOTq4S
cU69ocB4OmpLsv7WqEciNumlDRTDqSrMg11b1p6YO3m3H2Qlm8E+NWaXy5wroRIw
/+7eTKpqKW+jaEDGZy+wJMRlMdl+FImd9MVVblFAjXXmrgy69NPp3YJKb8H04pp4
I+GGKnjE89Tdmqw7HPTe7/uNIiBMtrIdsT07/Mjf5x+BToz/wUICkeDj2pGNWGpW
hFd5Hsq9SmH51Q1VmgFJBxaeJPrKOrGFZd5bSoNSKZkNHb++RcahQ8b49xlh6JPG
+MnU5eCcS6fQBtky1ekJkpkFviPsUmXGie9Tcmve9IeiqfS3YCzxZp4Qt24R7Nj8
YLNTxZIAU8RIeZqLxI0pSa+VcGmb3y6jUyergo8VqEwxkFHClMtKDpkqPpPPp7KY
4a9CLmf1P0PMm9IERT7UiA6oZ+UFr0d/tPfim//TKNKbOnP5c91jhbQTDIw5Rs9b
Ij9KGJemkZ1L4IYuuVoDaLygmHV7S6rse/utBlPkff9+mNAnADaaN/VNaQKFgN6W
qbMV9onMxjjD7DOv3uZ5iqKXn8S5KsaoPGEdgpROe8LOFpODSUcMpfHxbAGEDXso
X99oWaFmLc+OYgYNPdcrDprJEsulvYEDxlzAyxXYkb9qOXkidGFE54NuxMLzD2g9
RnrJBqfAQjx+WpRt0MJCkgCsCS94PA2rbkUAdNR2EW3g/RIaABbwqceWP7hvtfa3
gTybs9VXYioDGEU/0ZB8oudKAhXBIqka4380Z5bmtUNe/Tdaa5bd7XQqTYBwl/m8
8BcgTZimhzSsbWofkev7vG9sVVvym4AHEHXlSMdSNV6iEfqULerFUniKktYEwSpZ
NK6vKd6Ul0Cw1c25m+FxU8fgWoxayG0dHh6/AXTrG5Ll9bByk0YEKVXezseUQ/Ct
u7zXQXz1sKsPZ+94vHfd9wWd7Ade9Z/OGbfc3hvICfBLGylxMsXDIJ9/X+tkqCyd
7J/vkZcQmjCb5hvT3hFTTkCqPd4QeOBRGPK16RnXOgJzNSrDZQgFy6uWxn50A8PE
9pD9/gPxm//sdTkGGTprA1/6xTqeHSlz0W0gmgBTax2rWVW8V7Av0kYcw6W3vAnB
ER7UFLGBL01aPvrxWO3NyjPan29QMklMmyvZtqC2Jqh/yxCZ2HrV7BfCr2cAFPK5
zZoFs2QwEgOcBXcK4on8bVuLKxdvy/b+qH+GCQvPfmUDLByYHPknAa2Gq7o9diqr
ZDCK5zIr/TRjuarjauXwaBZaArDJZhpbWxyuD/yqb3Ox71HzhS/y9l4Gz3ZD8xgE
1e4qD2cwXusNIMxv7AebIQVobBfJyLEQpJPEAjpdihagsYFseoFyTVdM86EJG3j6
pazMDgdFdq+19GQ0S6OWD5jGuc5rXwjEcNE1ufdjxRGsTT2286fEQJMN+6zgR3QM
dNzVvGneMsBOq8E+cj9y5cb6TZinlcriOP4ItYhjvwZzIqWM4AmJoumtiEKLOYIJ
9mbfeh1qkLqdOyx9jylFJ9AD4RQCnEiMZU84o9Fah7+yHS/Vy2FqWUjeE9PHEDvZ
/JgIkqfJjDiK7bXRXuti0I/kZ/Fp0dI1zUPBTfRxX2c5KOKIQYbZsUTnXnLX29IO
QMrRlTVbXLV0dOa4cEtC4iETDu7t6O5TXkqNFcBgkoMdXniWPw3H2YMZ58q3yr4v
GJhgsQQVgpHus7eMi3mOPgzgZcSpT5hIN52p9iafAKdQfkswIvk2TEmqBtR39kGc
9rGzfyijTOf9U6Q04hFrStCTYyZ5RdL/reGMa+F0l/DPeXnP8AgkgLcbHxoNUhfs
efFxaJO3HbWsBotgz9inJdqM1GRAKrrAcPE5nM1tnqG5eDC/OSYRuGyYmLCykw59
Xh8+rsta2wv3uJtUsM3t2TyIW0x4w5r0HC82olmbl8/qc9fOL5TTXFqargSzpGsI
onxDMId2f2IL2u3lbi5fDjbUt/52cdOyIQGaGBGrupxO1sC1QTIqRiYW64jsatJI
7sb5pZ1et9WsZfE2fVfNEPGS/+uOKEaUto6TFFQ/2kneZF3fLyOtHKj+nn+Gn/Dm
nu1O3QL7WR3vconQYSf3/BW3bkZlijLRD0xoX2CFlqeUsHWbmeyRxufiK165A6KS
9w9KYFPofxDzfT4EQnDqHPjcFbHa05b+VfBI+XwVIwY9L2xywcvDTSNzBAApCsEB
G7qJQpC8pOCdxltJDxakev+02GBpXKSg+pGL8bPyzXNhMPlJIBxIkXPW9p7Kgt5A
b9YJ3FZIGd1YUwV/OJl6+BN+VSgl1AHnQW2W8AYiYMw49LIiJewMX67nhwY4/Wua
kPF94lk/aqOZnsFSnbwZRxG8fXn4psSur9dchzx9YfEfK5unVxASfglfUC7xAnVO
pVtHbcn9a+0g4EM1U4psb4+POz7bV/AiOZpBF6dBSWm71t0KAfWbFHFzDsyiZfnc
GD4gjhew3TCUTCNvudB6P6n7nlHvJX7CCo0PQOD/IO5jyyhbCb1aNsr83MTVkz04
2BE8qhwSGNCJvDL91aHDPNN/fKE4wIFsV3mekYkLEaKur5PgMU73VTdEnQ3WTvgE
3sppw3FwQPBd2C2BCmB1sE9QTOrq0ANB+f1eRx54PU6HWWLtJDTlZqEYMPxFJQWx
cCVul4IpQFuAak7MaHZtY3ig+3hlaEZ6tfRyn+zFGzSvBIHorK3j79ApowNRBB+z
iZj3DyXuLNa6DLJt2OKdA7ZonNuTp0hfHiKJfM7WNYp9/qSsDBLibvYvxoBkPg43
xPaktB4zkBVhcm3gjPSsDIkp6LKjhmb5CEAmRm1ZzoM/e7nP3uht5t871CDq546h
Yq3o1ll326L+gFUcC3/c6UnbwDW5spUaZlgHisv+31t5TYQsJKcosrmy7FQyW1hd
e4qSP1lV9yRjVRszMr6lmsYILlEIZn1s5FfFkVEvK/D0HcCoFg3srf0OoML4zy/y
WnFm5Bb5bF6K3qRclS4C1EjgypfArd0mV6nROnGvqDznV5xmmXk6ermpg6iuPa+p
xPBMbx12lCxWV80JoscN7DJWVYeullverS2zGkWtswl7tfnK4gF7fhr4fyZ6rRPO
lc9jvclSHKVSq/UKo7Z7cE1Ccme5KmXGM3GantSF79B4yd3Om/J1HewKQDE18cky
EZ+B5x4Rg0EFWZmcLd9zcTdiESEbBCvcnc6cQmFnqcrTSO2JyP+lYHO4PKRyN4N1
uo5+Cg9DM+GzJd7aesE8DCXVubMvWcxWZoPH79aq3tIUSjJ0vSLQx6leF/B39PcV
5jwksGrtNODIuN0s7LPJCQbfn51WhbzSyuFIpdvR7U2zVAkmp/wjuVIDRTL7GqX8
BsB4O826exBEB186351VYDRAG50PXh566W6iEHZdV26MXzj320euxfjFDxElGVwQ
2Xk4oOLmMy8SzYRCNQuCVghOvZ9aUozbI16Tmay+LdO4vbG1e2LQRx1+dAgf+aTv
MdR3cv+SOeS0CpdmNBlRRSd9JFSDOJGX/PURS/O2SXkEK6emZFs03+qBYzTgIM7l
tzc6WgKdTRDM/48QI2UbnJT8RTisBEybcC9/+o2rixo9/wrr9HjDYNFZpC9UtXoD
UxwKPIrAr1WEXyIJPT5/4lslakPKdA+0Bm9D7OJdlHpyGASlJrNKk42TCgUQyELY
mXEpmrmn9XwSFV+vuumGUNLII2rj4f02Y+tGu4UrPoZF5Wu2T8sb6axG4RNc+3pg
aIodUD1253c9bjI/cGz2xr/p7urHTRkWbUyvpzTVr6c57hecF87Gf/3AxzPqftny
JmM+rUeqkzOpRy7d2nCes7b7c02hPuEVtZXJLt59lDtOBhVV07jVH/9D1vg+kwA+
5SnmwIlrNMiZS8knw5eFcEKQ0kPbXwURxM45UWyhQSbxl0qQH/tuB2fkey5wp6e0
8ORkZPGRk81N6t3CnNAbqczrlAmLgz56gf0gtZcNMY6BmuEJ4dKYSsGw8n6n/voJ
Gp8xvSZIDmFWcg1m1XKH7kASmDANTlIpanGlJVsu6Pk2fp69VRqbrT5o4dkE82rE
AAMt9KO0nrm331xXhTdF8Hc95o3ICb/kME1KQVXm+Z/PuXI+Tgw9jE+g/8GnthJc
f2Sa+nBJIAAJGLeZqglx4SXqjBKQdjRUlWdG6u+Zw9qAzlGGKoLnXL/vw9SbZrhd
nU3ol91ZxtD82pFI7ZE0onVjB/63FADlmWlMVC4SZ4HD6DaZfVhO4mpKrTI7M0aD
v13KpHMUA5+isZZ9ISXJfR/4BLfXR35u6zEModjWvARGh4F+t7JmE6DgZQ00UGR5
MKH7Ups/SWnbOTforo3av0CDWtZ4sWwywILnZ1yMlhnX1HdJ7ls5lNu1BCA+AXn1
H8+x64QD9L7YF2NSpm65DcSKZiHKoTK4vEkFDVaKR8kAUA8oZrLiVCcrpbWkQfFr
LGu6iERNxuWwkCP3N4yoh2K3v6gPi8rOjazvxwiSLmDpT90V1t+nQsoWDcnyo5I9
8aemTCWt/drnVNnsG8F0PjxhJU3D+ADk7HJB94nt0SdLq4lino+xDPrYtV+9TsJt
uDtOZxmzYostKh2WSQXkf7gb3wXVn+DvJWIkbgMw9taZlkKbLS4yvl4UFqtyU0Gt
r8mqvgDI1OGRls2HCvmCvFzJBBt47OglirZEnBOC7FKhYmX1OhSGYkAWnVmFccIR
sZLF7zBY17hjeDYOgcyIhenyPb9ESnFYXnhhnqKg8XKoRgdz3AzrAz8QgfQzrga1
mQazFfMg0TAiDnBtLOgq4Lbq/VnUowYhQm/09BlyhQhdApW4JNrnPfRKC6cUiGdH
WRTQHZByrb9vEEebwTwsVvznHdYCXy0Wj5HODNN9GPYSXK6cFpbqh3eGWtIKC2po
6dp9zIBkQXWKZSdCqw4tPCLhZoINAfvcw0SKsVjRG8L3TRoe/XxG6wioQKwy+4KX
VP9+fqmEBpym9B+LpI2dXjhNOERsnu2C1NYHuAKd9/BYfWvieto5W2znttfmLB4h
rp2tnrIaHHaq3I/b1bVN/ogSLav4s1vpPnmb6l0VZ6hQ+yb9H+R9rXNMUQMcj7jp
Fef7L5wbZObSjoy+GGPB1yZVC9GRIV1HWraZbzYahY7NdbV0xsAh/73YavQlnOfg
cCk0Kj3MGAD78V9sDeUpzS/KFfRpbCQeEOJzCWaLZC4hR8o1QAZJX5JaqrtIIPJO
UQUGPYanPX9QwoUSt8/gyPRbRx/6gzGk/gQClZUMVgJ4Qv/kgIV4J1c7ac/EF7ut
lONLETvzOErOSNo0ivfZ4l8Gcz1tg4aEA5ykfVfKy6RE+yR240ITwI9myjO4pBj4
CRtEcN7tylyDqACIv3Ti02qtwqC+GniEl4SPsvMFcVn6MyKXRuOYV7bkLHEn1sAD
/1KDDGeJ/16i49YPtj92iEU1QPgyuzzWfiHr/3EVllJJ7ATwBNkz5+JG8lP9pLSZ
j5INn6i7znpfquBb0MpCcs9bKP5MBEuEcBa2UJ46+ieqYkfS1fdWjoiQ9TTXlYfx
Y2eJUhlkdCTDGrX0f+WO0ONkKGkj4poWmyRhYHMasa89cyrumOQaPQHwmrs6zk2S
B3y5w/D1fZFGHheRD+z4lMcVKyMbQMUXRs6xyauNiEmnLgJc5gfwFQVMQVnlXK3n
HFnPf0zd1KjuNSvxpQcvd8H8pwGYggbSuI07nr343+umFZugztU364B6VoayM/ML
koviVwfLoVfHSZq/bsZ+MpLspd8WDEs3HXMX5jWf5Ci90SxZKbgpT2A0dSSMM09L
e6n0CREtD8+LJQpPafCXpXmyGSDRP2Jlb2IgNpYLcoMsS8y8VabdOk4JPfstx8kO
fYe6sDDaQNeJcgTBgvOCy9HsoWJDbbs/vJPmF94xWYT8aOb41AhmIl4nOwDwgrEf
t7CaYqHyULxBeG5OfcUtsCZpVxIxm7wP3W2bXrwVw0sh1B/GmCNMjAfNHkxG3oBC
YHYlalRJ5TWIzAjcoav1cA+/xaHIT9uIPZjDtugahwGpYTnKrczw/jYxwxTb4JSh
4jRp21ui0M628NmfstOHn7zxskz44RDu/lrHJ/bK/3urAtXqYVOiQuHvnYipH2U+
ZmP+4HJggFVOkXeTK6+GBasD3C2gMi884b6X4rm4oUaGzi0FKov0o0UPVCvG5VoZ
AgmWGmDkb08d25F324e19nrK3kzj8IhlPiI5IMLPFsyD7xNxsPragds8O37Gn7kx
`pragma protect end_protected
