// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DOjgkkX/dhj5BqLXcc38eFVL83ZMb1OhOygwb8iLk4OsSlPdZsyuPexefzXRMRfE
PQ5uuG7Cp6dm3qU5KFg4fX2dLMVQbAumXRY5fxeyoXkwSdS4OfkhkgrN+FsDQkZU
RchrGTshPxOm/4AFXxsHNWD+BkGilnSG2FGqkyABFRk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7360)
kurq4MSLX1Ps6yHqVLGB8/7zsY+wr1YqI1i4npZlxjkHpF+TuM/llE5Zq4yoXVNQ
63gK/9ty4ZWAr26MjIbVl4yhOZJhwiJSxx9FDEEh/F1HSMI3h+swkbNXQYAnGyJ9
L+j+pXCNx2wt+4AVlHW1M2O8kX8n0RCaTV4VtNniAA1XNorUUyyoK+wBANm1XkMW
I08w+2Jay4RlZ3chvTf5SDCgUdqrXjwfqFionDzKoTGzyBbOw9H/wcVuVFqaEDWf
AqacBKlEcBZI7Ft7lNfxblt9fTzUFdF+J8hclHqqh7yuKWr1WF7UsKwtGbiozEu/
iel/GdV81K8zC0Gbv2Z600c8h6+PHL5ghbGOMXyGGz7efLQ6jASWIYTlePJauMep
RD/nQD7vJKDtzPyKYFUwTA6L61Onnt79n1145vU1m7HL9tHbK7yj3t3vfQT6KfFt
giwZ/ieC1b8jrkTnneCsNZxouWxH40UE1+ahGj0MAo18G2A+ZMEqlBrZXQ09V784
b13PacYjNymeWeV61/KrBfEpWFa0vkBrhFQi6JZ2SA7A2Js+m6MlNbv0B2JbzfAC
Z+ZGof9KDoosl6+HIDzDjifwRa0UxQyWPQTKqeT/YS6jzp6PzDmAOxeHnHrDFtv5
1TsDl919i8lys7nRrS4VplF4g4AmcEY7ySSObaONbMq0Wrf6ykrPfeFhB7fK8qVW
jlRwaU0WUZzdaczTw97vqPGpI3CKNarivdQBFFpOHX5zQ7SdnXGnmHHk5TO3h/+i
6d+Au7/HNvowEKGNhHZH6OAdsNkFRK0vzTKIvL0ZAilh5kng73JEOp0RFskBHHa0
lGlOQlvzBFGDkHmHPAqkYrX76mscywkQ0d/XCQebH91qkydkucfVXad4T1ywk1DD
Fwb60xfT3Wtddp0WcUYTYC7tiFdF5SNv7Mbo1XW+op5CRdtXz1hUoO4vpZrcfmRK
OlpxEUQZ8yZ6/Cm3LEofFwh+iLtoi/EjP489c80MMRFjNmmS8xbcLIAyuUHYhgkE
jU8SQ9CiVJGcGrsP9mbfje9+ixdxWYah1J6NrGEgdlLK+1VvNeHvWmL1hzKqSUGZ
jNu4U1UZrIZn5lMShoL/7Lw3b/Ofki1obTtcHhhv6nuNVXDELT6UgzcwDooCJ1yL
bD2Hlk9ky8nNnJ6ZntUjYZdbsNOMa/HftIy3Oh8h7oJuB5kjiRNQf90Kzw006DuW
3JqU44tVmUqBzyM5Im8ORu/axBBfva1oBKdbkf2fM5ZQhdcY5ITtuFp8tlEQpvb1
VKvKMcOG3PCVSITslXQQVKDjrknSg4pxv3MlPS5Tp5StpFTUIhFwfkoLkRuLPyjV
puKzlKsdVFVgO7sVgXZ6eIfkiCaQjDBK4knxsWOOb6rKtFncHFV69sotNvzB2bK7
Asqvez/Nk0djLFgu9a0E27Ad9iyZsj8RNjO8GQBNmtLnb0mm1S6VfU3c8hDuGPIF
Zj+A4ime8NnzHQtpWmHVt/WupAcSKFbIrQ2UQzIhLGKqqgKYjPgnGxjTDmmV/eUb
d391RMv3+S/SiipC6De3jdaSAeSdJDbSi2CGLuudPywdBqDKMXRlU71Lyw5LKENA
5M1Ysk92U2G4BTm0dOlEF0kXRhP5eewtG3g9fXyzOll89aSwAQV6rsU/e+eAeuqk
OeBxFQGjSX0x6YFGGa1EKIsY5C87BlA581YJxjhWtHCtiBqTPjYHUUmYcIdXNT2F
TcEc2D5iMS99L8+wo9d1d1pzCCOBwlrFEzttQ3h6aYD8oyftS1Wfd0vqwNWAzcO1
T3vfVmvcUyJKv8KwsBVCsi0/Bmtr5JRIkBm4OGYelbpU7k8lc0r4cQdkjEHvp97L
hnKDEpTrjQFM986tC5uXesn+9c96qR+LfxsMZ3UMXY6vNQ25V1gsORVpW2JHjSKM
1hwgEZx8hI2zhHxGdQHpoKcdrVp8vsUMO5pWjvVZaC07O6TD38D0xh/JNvaWjuaD
d/+RjQELcv+aaSS1qRLns4io6AwEJYWA4H1l8TUC3OsbNYa5+GaJPR9ae+tpsffW
Bf17LKEmcYRo+Ep2H50dBeijWoomvKRhNMq9UtYS162ofKyvqYyDDQ0gYzCXDPoD
m7JnxKxPJVOwS6ZL8o1z2gkCdzs6wRgm0H7gX40dw3kvUOuGyMXC8xI90omGusf+
8AIpI/+JL2tLvFG+i/eS9STGN5INpp7IV87A6afVcdqA741JGKS95ZyocXyO+uew
4Q7XBKzx1o5zdf445rHVEwx3M3ra9cQtR7lqLRs5ndGDK+jcfkcRmmCqZaa2JRIm
mFWRLmF0y7KxdpJ+hTpy+swknmpFwuLJmJEDs7KJt2gBi3UHUswtTgdVqc7sp1Ut
+X4+qoaPj20ET7R/XX4C4Zc4LtCPh/aDHBc7RI+xPnbNbt6kTpC1ZvVlDkQdxypW
2KPV0VAMixIoktD98fltFrW9nvTP2TwqeGvuz5n3W2a+G0GhgMAdOQtUHaII069z
IIQqhBdhc4DMGAAiuvO2SbYmOsAODgjZ8p/CMYoMaBfUEiYNGq/C8N6QGJX63L4a
/rB0NiY/jDgJj8qNqP1DRqhL1R0aMjD9nULU/GSj8VWD8on8itQDGixJZIz/feu5
sXWCAcVsf2Hi4zumDxAJJ+OSOfqJjYDvliiYYf/vvLi3jgczGFAZ2HgUh5juAOKO
cWQUXIhDgaUFRMQw65LOPziCw2MabCjEDfFiI4qu+zrk7xfY395nKafSrz553ZyS
b+NDlpBywYqVCoDb0yzHMh0yKOQnxzy7QHo84qSPxUOlDZEqEwaXjdGKzsQ5/Ffb
aLeikhjKnPcbkeTGzNzIVcqFBP1GWQtVVVAfVi837IQW6cTUKqNUnDPLAB2ANgfW
pWlRwNvsPBEnk7NCpP/6SJDrLriW7PEmD+2CnW3EfOPaJ463LOkP08c8Azcxjcw4
BndfB7WFy5JkErL5TElURNpXC0mPoOx83O/XZYi59apmm22rSTX/FKDhkgOUKszW
0DiHSR2NOLqUD8BbfcvaMIcmlYOhkvRUNYtaRAbaH7YQpQpV7Zvj0CaBVZeFvcpB
3g/cfJZN5P753XHup3AB7ytnDy9bGCHodP7Sihb41wfVyYEeHQWvkv2Y1jETDMh6
IRcXNq19kitjtBQ2ACgUUOgMB3zolruuNp24OV8mmc0IPJw65nCrZeUeqCl31o76
WiLIo43ct+8n60Lb+lsjD/AGEQtI9q2cVyxtTvetO3jWuuFQoIo6tIacJYNFY5VT
wQPtmzpsozYBK5dkySo/9iIpHMpz72j6EIzoydtjRaC4B3H0c+TZp+TkBWKPRNim
PpJgKW0cv/f+OWyhLljQpPcbFNTWLAdTmid3tN8gJF+qMKxcy93LKOiPlN5CGGam
01prLkRwvLMVCHBoJoBLzVFekh9uj+lo7pE4Y4WYUzO1Gl73MTKUk6Zz1tTp6iok
STVJ5v48bV2HD12o1FN+Cm2Hb7+9bwnRiUcPPdgJ9VJiCiVDY8gTHbQo+XNyrBYB
C/LoHtTwbE9rlRt/gLChEm1ylZ8z0odqUer1NSCjVx7NJABZw7uXJbl3coiHophj
B/P5sAt+8Rzgsk0rLmQ890ZKs4NcXKFqIY+a+H59sc4/7CaFlyY1NT7NpWj8ya+l
HGz7xHmEspGjhmG1SuqhP4rNJVYDIwyj5JMe0keAMmnOv7oVZWMxR5YXYCDtdgqH
E+GIDzvdVJhkbhQlljVieKSv3WTLkLyzZLzCNz+68sRVUZKTCBducHKbRlQhEs7L
RYzk3A3Jk51k9QDD2wb63c4tWf65YRjwQ0n0fgLkzcW9E4ZLGGf49SXUHJwwDzP7
93GN8uljNzQp0iFuiMpB9L+AUUvHjl7JOH1QXzxcPr5kRPiEDjdPvo1hWKVpK0tC
koz0uGjQ1njMlbvxwn0NHQP7M6SkpAG8te3XWM5XrpmyRpPMI/AJ2H9h9EpqO8JK
bT0Ig2a1SlimpAU7mR/yR+l87GDM1Y5bmH4Y2XVAOZuy5BiRmPbY0U5EO+5XJ5+M
WcMsc2y++MHtHbgS5tDvYOou0MWn9rN2D3lnd3ZGSK99uyqAHbt1WeQfQaMErzCV
tjRfy302EcogdsUiOLcerKPDfNwtsfb8+RyJnihexF5A4XKOugTAjNrjKrwxeZkr
AtKhMKwaEuxVXY/fvuSlPtIomg+zWlwVQTHqRdm2f6KjjZb+zULJu4fzuFiX77Lv
91wxizETXUQGITguQ0lIioMdCVBkglP9WL1/YuEHG/DFh3H90NWuQ9BSnVrxgOAH
ByTt0rBW6g2nnSEDRs2U7jffXQ0Wd4Zl9qPG2isklq0nXp95ONbkuroAwQBV1CRB
hsDzfxeLgpwghPJLJD4YhxjhHMcNe+mewUHvKB0ohvm3DZIwOUufH3ZohGrdOlPT
HmZFcinrTRzCvxwYCZFSU2oHaZOA9cE43I4shMuzNUCwO7+0ndp850QvT06ZuUAQ
oMglo1U7NUKCum9BZ/n/SmA4qkuG2dYqJKwdMb4U54HGoNxF2yeQfBJiVc6jwMf1
4crGNvLLJI47blaZjebRAWq9InrCBoJUQ7WnF7Fd4DYKnFa8cBI1Ph82wI14S8MP
Rl50v9cKONvh/rYm/0lm87RFu8r7833Qw2cl3ycmGcpSFgW88s4TQ/wRbAHl5JZO
bIEqQuzICN4Q3C2120GIrVmRTaJ4ZJ1RkDPuF2lp8tiumWtWT+EksS1z2AJgzvE5
JtjPxcuZUwi+thUOb4PnoVWpcNSRrLf8jLbA00QUFdzCbw1uqBEuyLAOu9RpMcnG
2u0oeNotB0uJCOfBGBz/xcbxlfvZ4myiH+LCGpx66XZX98Fh7uAYI9rdyt+SnQgd
UFy8IZjlkDNdmJSEhZ0OI7x+A5fE3N7YlDTaxlV79OgKCpi51sffUe5I+ByGAFKM
z7AXi37/sCNKYH4xK3g5TeJSfxzPcfWHR6d0v0X8A1GJ7NvUyU5TFVYPAJHpow7S
bs1oHo4p9FjIicnlXLUdDw97gnhEaI8XBxMS7N0sYFaDJkt1anrK9UTmgUWLsBTX
+51C8ch6SfPbJTYvWCtj15zsELdr1H6nXZIxknW+m5WELh3VzY83uoitkL9mr+Lk
S3zteQWtqwIIOOnm3O72gd7Qj2kDENdebY7tezLeeegirOLcyDN+ZSpuFCnM/Q5w
/d/hn1BrXE86Mxov8evzj2n1iYItvgEaC7Vhjt6XX0AHhYBtJgi8n5Dy15IylVVt
PDKE4LhXySxgjbm95XsOKMvJ/4fsnQbiK5Oul45q1PD5zckW/rulxGfYrEJ97Clf
QcAb0AmeQywSCJxfJ2WPusoXs7NbbxkKaxVLTkM/YxRJbMKhZCe/GCwto4ziI5Kr
haNo+7kRcnTdZUzr+ijPXun6klIp8+1GU3t2ofvMmUCh3/Gg8+Tx0r01Q8Lrcgz2
aWTMBx6zpJbRZHv+TPCUHVYyfHB23FwhmkP3iOSwwFJKZA5nlpLizdEv+M/RM0Zt
yA2R6nyooVRE3Nn+Iq/Cgk/sCq0o+7bjvuFAxldF8QJo5/CvXV5vpC6UPbNjZa9y
X9gEKPPcwQVlPzJb4p2sObOrxl89GC7xy8qCoGOt0B7hK8vVJGON5ncFsJu7HVrt
edCHmI5sC22GwHy+WyuwuRq+fc0H7A98YGgApLxnSaAvn2SoiY+BDBHZfO2cLsDJ
4Tad0D06mFKP0iAzBMkTQaWG+JWtimUKRmGIZ6vduux1xEcAoIis4jTGP85eCYuD
d+vMsTArtezDS41KU+OsPYYrSMd0XAaDtsTsy8eAHUf+4a7e+08mWe5RcVFYeoPp
nufH5V6PPsTU1LToKL9aKmhPh4HqMigmLPmcNatmDlDLj1Cy0eKj9md3JxgYpWXU
iYXcqWmcmgcZFvHyUJAq0AOWpUQBO+05ccWNBUJuvAhGr3nEGngJdePGT0RIoRcI
bNMcpmOdYQvyC2FsC2NZuLeeV+OqkWn+/zTtYzGasfdklnFKg1A83uwu2f4Ypb90
vSHMtRGGm9vnH2VnwQemRJjvROjY8y5Hze4dVw/rI7tqTkhM+Wh3ETFQ2VmgYnXm
D3lVk+CqXFsU7tHksQPcCjiyMx9oYHQalfXaqljfe100mOXagvquw9GKUv07HIPB
5jaEmbqytwOGtukT6hoofCcIPxiFYU94F1gdqwkOR/28mE32QZJd4+sI2cFepv5v
sVnV/kXq1gOqlFiNsZfpJ8jifTnFIJvqBpCsegXspIQ71uLQpGlRo6SYDoFPKBkk
X9e/DpfzNj8gyVdwh9Zqx0YrJBrEFP4ZqxH5zVwcYETFsPpk5oHQ/q7sqbO6S7Rj
ZkVRkyKzaCkAcCw81oB7E2vIk0y8yavpvCvbafHVbU+RlIso/90nN7wIuO42QweE
As5c1GKcdGx6Xm/RYk/9hPNYS3oI4b2hUaU9utgMZnWWZYrIkIc2JhKwJHXR6j4t
Z268WgcIDBZgmsw4FbojzPcMKA5Weh4KYqme3vjpDR11E1MzM+GOCyFyxr4TJUMY
/HS2ILK+jAe1zG8KWRJgQQDhlNQiy3zziB6wKCsZKgPZ8OGpkNHCEmgWMJRLp8cg
n22joTGKYJkXf8lA461M1axkw9amSWAxyO1Zs7sOlxH7OUjEOGQWL+Gkniw/ASpl
OXzGpun0wOqTeOI0KIW58WvGgdlielaqs+78HMCBGJJI2wSZ1spXQdBIRlH3jFCR
4LyVXelVheJ4SlS90+g/VorgJr+NIndOaoqc47Eba9RJ93s6UZShxsLxPBsHkzOa
qLPY1DLXF6MbDirerIEgFYmZnba7m2a3l9xxV5b7wEpzhs90GGy47lprdIOnqtdM
OwsQHrMzw+giUrGljjgBPqTwsDGgbf4omkwEsslsLVR9C1CbDFENlsTVaVMz9r5R
A4RoMMUUfkiII2La40R8dKgb/TyaADG4amFh3smc+p+UMRaLCpe8lxK6KUYofTQc
LpK0cBogJjNr3dW+kMtm9SYKoG1X4TQU+1m8v7NvBe7oAe80ZQDnqaopbcM0EK1d
bGMUrQpIaQTkrhKFaml7TAldU/39Ov1R5eojv5jxILhpFIo3BP58D95/mUcj65Jl
YWljOVDa5xzfi8f4nOMxnaczAZ2iFVLXW6HbkBjz3DnBi9M/JcKiZ6bPyxKh06ny
IPoae9inwYjmsmcrVE9Vm8h0cKY1bbI6FKqV2l6WEivpIA1XIKmPZsttEhytOVEu
lO5Brxh0pu1bBybL20HlgUm5k2LwWv/0YMLMZ+2tyaoi+GyZLQ+si9t0oVQXg2rR
/rH/O98QvHa+b3rn9fXdG+9cHyWl9Dl+pVFfIKbia2P09f3dA0XVhSRx8MzvRex+
D1vvtrsn4LKoo/nVrzIEjMBHOrxar0ft1dJwlFAg5KvJdclKqnhisJdVxfmWye2S
41NVf/zFrj0g0Fp82cpLrW4i+SO+kGIxjr3dEvCRO+nC/oZz3m8z6KIu6VUkgfyY
SMTq54BPtk2CJDnTtdevPVfhsZ1n0ld0LZn6oxbJQM/pdPhNRkyIG4s4MNYQvu1t
L/6Ip3ZF42H2uQRRFsog75yb7yUPlYfITmym7KUiWSp0v7l5Iu95jOAh74e4RbZX
Hh2ekl9CT0FL7+NoBiUvUGCbF8zpVQ1MWse91ENo8R1gZvojH1OqT1DW9WNsgGof
ciECH+mYx9QgeQzZo6f95OFe705JuZI3N2x/IGB+ETHMaLyAgoydoCgxH+Kk01Uh
cz7PjIrsYc/NYZJjLLydl+q7PPzNsKTBPFmwebgNF66uV1TZvffvcgsqdu05w3qL
XbXLvgfsl2BnoydJ16NxyG0t/JYaMPvtjMTyeIkH2118hsgOnC/pXS6XqTyGlffl
FCbi4W7nOA4CH/6j0Umpzk07eD19PoEdccV1NWe6YHaVd6Qri0f+MJdxRWU8vJYg
PX+0bYBxwwXEnVSH1eKN9JjIRIeW4RGgwwTnavTOMDTGQw2+xn0zrXt+JjBat5fw
dLRPMBtNnm1JDw8FWA/icmjdkWrZqVnEY5NLqHOsGTtNXqbTxvs7aL+jM97EK9YE
eATYe/MfW3qP1QBRw1Et5pVX472BFR0VogavSmSKPNXZ32Lp3iMdUTXdKmxe3saF
lA9jMnuWdwghuUgxh7bTRln3f1ccVcGwi9J3NwjwOQqXj/PU+G2XjrEyxdryHUuV
iechiFPOTB6or2goYZ2j2KrTDNAGkI2ZvMHYbfBg4zuTwqI8fAUJsbK8+zlJljso
T7W99sgJLTKhnUH6YxiWRTg3Z1AauwFLd+F8SbZ+NJMa5/859W9/aBbSuLJfgwZo
AHfXikgLNHHpRQpT2Fd+mbfDJELNLeIUCiwglu67GeARWRiWFZvvzCjFDgL7xOLf
JhriPdKOJWwGQu26Ha63cF3BhSpubKW7kvxoSa8wfAzoQbU4CJr87GvcxhU/OWXn
vxQTJdBP9xoKcAZEXFAqV4ObMEUHfrtoUQvSmXC8AXw/pU9M6gezlDxvvTVA3Ttd
QcFjWqTjMSPxnEhpDUFgfR9hKnT2TvLT5EgRDnk7NawymVS69HmciO5c+Srx/uWG
pL5Rlnc5cpCE/k4U+VEamFTcsdu++MoQM0Pr1GDMs6x+qGt/mQqANd6H1jwyTy0W
ila5LlVZL/F8ynfjJUNj8sDYYqHk9NBl3aixrGv6RBdEqbb1VRcFlDxmLvzHnFSO
u+u2TFOA2DwNetezejFMcxNM0NQ7d/58fv4389UTu42uxKLoVrW5Yd+UN7hEJxb7
eaGyQ5+BzZdAbh4HMXfV+YKDZIt7IT2UomHDHQ4DURP6Mh7uzE1+PyJjtXfhL4lB
d4UcmYIQdn3Gttl1sm6u0+6lbgUljdM35cdqolBarHOKBssd6HAvzw44lSYdDCCA
fVuCWWFsy+yCbhrb1E4JhErBU4kUNSio3RWcEE1Od05N/9vgUyF70MUS0zn6OGmM
Ensyn0pMz3efBktyH6p1XwUpHWw0uwx2D509lDlRdovtgkehNfiioyuAeVQYWhAv
eeTl+GervnecNEj0+nTcCpBhXVn6hHCG/TeSrtChYJKqhAGo/4zHxtQ7DnV6cndE
rtF4lTp3HVP+lZsj5aqZZTL8j5WcNPDJrDME57JvCOF0IunEqyRyieYiAEqfBfIh
lC1xuAaOPIr0bKuIFE9TYyQmLfLploI1czq0msijfY+98k/0G0Chj/1zdWOCKfw5
92uSQ9SDhyPN5RZlDYfvxYxvN7XU2zh2z8YxapDdOamB80r28ov6P5SZS0r+tclW
ERmCzzw+QBkfusQtHOaiIeb5S/ua/wuA70GjXrNXcEEe/ZK2w3icOD4Has0loo+O
FeF4yXnZjtLeSqvJQYuOnKEbj2OP/Enme2icOvj9RkpGhpHsIgmxXcpEPek3NZW1
PJgYc/BHAi4KqTpvTI82D3feTX7iTeyExJsYsD++B5Wi7FnrsQg2zJVPIofdAbXP
3eZzQ3XXEjN+LzyLTKnVIrfvHRM91UU5s7kPuU6ABdoR10IzUENFXd71Mu8i7U9G
2QDFrsLyjqv8qkjxEp0piRR1fH3mgl7roIjpjjKx34kfChKO7kcfGJjW/sVp049C
BCLTsfwhM2dgU7DAS4Aytoi+4Ru5b58SZEbD1BMqtxWiGkgtJpVvLOGII0H4FJ6B
WTCbtM5IHC4mmHW8rZPuOpzMhCRZr85fQG7iH1oL4BVN5+zynZZREqpS+6/4rNHZ
FrtlHbZ615x/Dt3Rbk5yKxEeZtg6v40WGlQGDPUVchyx0QA1B5DtL9jVUKNr6+Mf
O0wQ8kCMfAeYe8RW7lRPCw==
`pragma protect end_protected
