// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:16 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JPrMSV+4I1X/b3cyuctE8N5Ug/HKPKeJaL9Qj30YfQJK7TU+WcUS+VAzyqtAvbWv
6Z8/7OzJSy08wuvxQa7Ehx+pJttXMPz4W+wiZWjV4OXi5Ds/HbZT0Ykei14gwb9P
dpR1sGnd4hE9Tf8M8c6hFuEiscXJ7pMoD6RmZ0oZujE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14176)
1q6t2JWK8/9s3whdiLRLPrWdsDxMqj7ftn7166c3v55PnT9XuTIJScO711kC1efA
U4qMpwz/Geul6XWeXGACb4s/7RbfA9/dqRqpe7NPauNWfiMJDitS++UJK0g4cv0Y
/MLDs3ceJnGTGv6tCR5JAF/+6aL3Z8GHM9TrqPrBhpl6fiMNI63Vu3+afrukbyiI
4FhClQWfkejBOBFzguND8knlyiwuOlTLJ3KJxrQ110FHw8z6IXXP1rGZJ3ey9lay
cgd2pp6WIlrfdj73MB1C8idwtyy5AgGVMqZ/yFUpEfhsX0BbqwcMFOlCEQ97qKEI
3zHRe9gqoX+Hg7M6CuRxg0zNXX35aYUZSpnFUQaio/tHF3yZS8yuAQFdlaIvSISC
AxZjf5VzmN99JkyowmcPbqP4WPqjm0fvMJyklWSi27Ecjl/JKP4hCMAGd2wlfg/L
NZ2eA/H0/XJDypKZQ0fdaB42pm+pvQdicJlFogeeXU2DcVuGu5+no2GCAic2SVHp
J0epfBlEkxZR19f8Bv+B7wK4of54+5kE9Qp9IsiuRYNZTONmp9fQuAvpwlVe/2un
8VoNhBLm8HX5zHQbuRIjuucnQNiZV+K0Qz0EbKWUgwZApoqXNCIsZCzTPTlPgaKT
aJXEQ76jBp5YChucg9DBNwqR9mVOzjqOt5zX57nrAPm07tSOVaahS27UkV6aQbuT
iIoXmmOJfX5kzb7Dsxd4FzERe9Yi1x15n2Ps/ybor+93afSXtgI1ovj+6vxg6Ab1
IRNrzVhWztrdUrUEV4JQ6J4xoegcfkvh7ljDRc33rE5jkZeCVPkPQTFk+U95GgtA
D0EbrZIDNfmOESomVd2inW078fNEVBmVMVFZVne4JuUzQa6oGMPit/srVfk1MCYe
kQjLyaiNVdRxzozqBuM1C69PftpHgmyeJvSSNW8jIrQ1tHX8BsJn9yYhyM25EXd7
XLiCG2O6LQmcQjljd236gAw1e3n516D+7IOty+BmPkV/dMb7Oe1m51r5Mr59qlZp
MnNZvZbVXjt1oz0PSKYRoGH4O1p15ujg1ityMDXMdgcVbur5GtQbxWGJvBo5AMIU
AJ5GgnaBT6bCTKYo12VeAuMzUXeZgEN1qwOBnwSoDNX5clP+9b/2Vdhb7qhjMvOC
NIkTPQi4UAxew3N7sNJT/I78Dkj+nhzV7KS8RA5izNFsuQnLrJQIkbXmLogqTw3M
UAstH9gV+6D13Kcde0fKDzoyNb5QXiDr0sY3/tRWWVLr+tUAjq88CQ6H3EjsTmdU
irwkQWo2sdOnlRncjvxI83qKmKBfvp9gJrY39h3y025oQFU/N6x+Vgm7j3ivMOs/
cqmLQJVjHNsTLBuNeEEmOSp1IGBvivwqIYm8jPUBpEnPUhisIYPbPY5rrrnCQ5P2
Rg/AAm1wGxdX57K8JWFOB9vZxyevNFiP4PLgoR9XoOiEsoaeYRCIjdZPSpjwEA2t
JIHsN+Q34p/XsXkVEG0p+daYhFtkmf0qT55F939GMaYfys+fIk8TaHcyTen7u/HC
TmghKCykv15fjLfBMIXIScWfdj3mNfzRGTdwg5grRVVzISRnsRzOFAqZd4LMAK0Y
HSIQKOSNIqVzE/qYMP8J/ZXvaJUeJKpxiHImCyyQEUsJQKQSYvC12uX/ELAPaI1r
efCBbt7FP9kgrJLZNCTwnV15KKwYt4aX8dnYQEtz87dV6vCIduzRcTLMSq920xZF
XMYGX4AohmePNgAUiEan1TNV9jMV64QnDo5xyBPBrQXbuKe9sYBExslcoJ53a0oL
w4AgEGEL/AqrAvq4ILbJt24FmUB0Ujlk0BWp8kLYYqq7STulvpvyzxLT8b0XahYM
dlygODT3euaueMtWVvekJQ0/Gd526vEt8L1Nm0yDFIiKPaoE2fE7JUHCPYxhhUr9
VCQnMEbgGrrhsBJfO53778N+FHTo+dOSbUbLXt3PzcLvriyNu76xhHNdwHZTpom1
5gvd4han6+AtiLT6v1Tsdj9HY3UGl4jykwiDvf/U9xJx4GwHD+TEtbM9xviEU/Qa
lLRzDpKv9ukpfdwDXw49WE10K6mW7Eju/ObNgzSjyWwckhfAs+CQ6TYxeOCVLJNW
JQ9Tdkmdg/geAf/wEW45f+XBCzp0k/wa9j+UBWW4Kpp1M51qRIv1oYf9e1tOA/6p
pwxjXv4hZol9kZr54uyJxlf5ttQACILLVUfKVxFsuFrwNmcL/DgFrm1n3OKeYwS3
WYUJcUtfb3hMnwojpraTe6N5bEmsiO3j31Ye7Megs9WeHcK7pP5cmURVNgrmDMvI
kC8D0uzWT8rdV2Y1uBgQwgeSU4Brl1XlX7Y4L85wPlFUEfPUThFmaOXbxi2j8M/m
7p5MXR3xSBPOsLNUxXNXkMdh7noTfuBSZP8905+7/V+OaliFjeAry8KAjQjDZtBH
+d37WLCJEZgBwyQNMuGRaazqZ2cbg3CjZn5LnlmqEIW6Q9iQb++un4fiF2ONXRTK
yx48wa3/umxiiAX1Gs4EeR2hShbzlgTqt5zTrkuj2ElmX0dwPjiKqDyBPqGjxCJb
PH4vvZv1ypP2jCzo8gcKxo0OML8wz/Ss4z6nWpRSwRbuQW91irddxmBgqbtzcBkh
vP4boV1Ko6s4s7081FzNZiUaPHRxEMYUqb60zHxJey254I9y6KfG9Z8TSAEaFySw
DYRR+Q2TWdpdZRYYy8PADTc2Acn+QFHy/C1mu2n8FXqqT1Pph1iFVHMJ5jOldPw2
U4WA2WOWNECDPBn0eDoHfO4JglPfLULlO7ljqpfmPnRSAaqWHmXO1tDxMCb0PguK
GicINtT7x6a2hBJKaGRvIXosDGwTZ1BrRA+qrCXQekF7VP8myBlDAQiOxNKb21uz
875h/HW+RfWJI3VWOgvVrakGNFhcEQyVAAA9+Xq9eqiLAwdD1HAQqX5HREI0UqKC
8mmAYEX9GDCVo7nMbqUMAO3CD5RPSaPlw+skdezgs6YhFUxnnUKG0rKoE8XSVlOT
jKlVixPCpVPL8EYcfsczuqGUx1sBU/80WRnH1S2T0sPaY8iouV6X5QiPad8RO/su
R6OJVhen/WbK3O4gHOLo3dvr/t374ThyNq84aPEa0fbWOL/lRJrQtX89JgEpbu6G
LsGmh2LYIiPQDkeRR7mOG+L/bSNv+MJinhPP/f2Qjx0Y1GG41YuCndXuXhLD9kme
miwuFmX9VacEHm2gx/LWDpo3WWZRyFbjSskyg2c3+Fjoqwm9oAmBxZ0CqkM68ZER
zytUqbaNXpGDEhHcsNmdMCBjK63Do3aFR3e6ps/lo5MnlZzQgBWJ/+6q+5tKAWXo
fyVA2PavJztIOrZzA5p69WPldWq702fvq6u/JRo7yYwapDP+GzBgvdNbiG/EeFIJ
IGnk5V7AUGMZZOOGOmFk6Pz0SDj+6KIxSn9ewqrtapVpKq2mfCKLzKWJZcxkYKEU
r7DVHn6Fef03LYwc7srEXdaPR1rXYQmNikXeNvKCDyi58pFX7He5QixMwXAnC93T
4P4rKv9+oifkwaFOKHaIlan5vpq8OEajtAVyXO3eabK7/aUQECrzkyPwIqHPDWUj
43/bMCweLCqs9dFOShfgT8s0ZqmR2M0Kfgq55KhykimBpEJRjiUAMV/tuEhnNhSC
A0fKpbTmYHa3eYa/OjZEyvNiu8FwqHE3fWx78dK7QnkiSl5sLHNQUfreDqbA+fdE
wnhx8Pm3gxAKanNMaMhNDLh9P2FYLJKUFFNwxGKytqKNS1FV0YEtQ6r0ewbH/TWL
qEV2h7xeV5rrW/9p4GnlaXhiw5sjkj84z82UBx3kyrWrAfUHOCBoGShV8T77xyY5
yM5NGX1B89yhES73V7udqoqTy0v8/VGBVxn+7QKSc5GAq+HFG4e6mIibM3mJDZa8
zBx36t8DQe0wpjBVOLwE7i8DKdcxV58udvUzS3JPucRQjAONIONLcLolFxip/FhD
prD46Cki2SCeCHYoqgXvHKMODraxvfgw+SkzMKml3RhZhB/WcTmnGSrkpUE8Wa8n
hwi/EN2Zo0g650n19+fdqrtA/bLfOhteStFPWnSiMAvKtXTcwtAE8dYf2eAJQK+w
kkXWbMd0VWLPO3ObLU9i/g9+KsEM4OkzRoLjio3K2X7VuQEc/8lchSRbaDG65Ywb
/m9U475RJ3oLEXHzqKWEcU/04cC9hudArWt8XEl9jzefvjr2awaTFHf5UzSrgMpy
e7OZ6DUHpTAbFZc4KOqaRBwTMcEf5rkKh3z54zSnUd5OsprJETG5acgWKlCE+9K0
2XIeMqhy4XrHS7LWNT6omG6SjN3Ig349R9qkn2BkOglC5443iiw2WHjyf49AkYP6
PiVnlII5FfRiZuOYJRLIFMvEFhmtFQ+fNxY0p6sFVvm5mcK9kdy7g1ZfiBsfviix
umKtPj42+LG6fdgI4hr86KUgZM3cvcOPbskh3ij5hfa7cTvNI3cCqbKVy4ya//EQ
xVZRN/Wg9HurV61wzfeHarA2nhAlVGP9ySzrlesfrQlzTvZS/Apfm7D7iYA7Hlsv
5acmoa+vVjco0z+db5vs21WX4PIRK/DXfYTsKy+0eyl4v5jfc2jncDmjqIP2HGck
z2yt2t3UTdpXPUj1ZS2DlMKonKFuIXsKaAMLTPx26f+L+hy48yewz/qOOgu/biKT
LZXL7rhGFd9M7a9asDeLr4gjJDSHAOzjlo5zwW/711Jg571yywW1Pri4SCe5qUAE
7Bez7UGDf9s6otn88vjYxKRsWM68KPMhDvotT/IdpljCbZtGPevSBekE8Eijve/L
mRk0HqUFf9l9PKHkzbK274mqIoLtRUHKfWRv7GdICFaBL88Gmh8pNNdYIXPlGLjM
yGMI5ignomXXkBARnKI52G7pTOckKr32CnDEl9DLMhNU8Zw0vkZxnGwGwfeDIov7
lLQ/sEBEq4p/oSRBJELSchWvpxuqHi1k/6/wdLCD7NV7N1DwVrBbSNDi1bn+J2Pu
m5lcvL932cxNXz81mZ29B/kqqVHQb0Ycp9kfk9oQP1MyryZVqildZfMfvYKcHUCj
pSIiyvB2myHlly5FOxylXghjQnOMRwpgGWT+CrqHy2B56LX1uCCEW0BIFSfee4ZU
NV2LhK4eEw+3Wn4I3ttHb1SRVyM32kEPAtLSetWeDbzqwGmDrQvcqWBOdyvTZvaf
TLtPpmtenRmMTiLVmZdnGl1S39YyhcGcO1mPmTnFQIf50J+Vf+chSVu2ZTa4OX7v
n97kUVd/Xk3d9IXHSczIhPAUCFQX2s4y87IcUTGmEK4HVjg4aDMfGAA8qU90zhmP
gDG6j3yEARlww8aTVCAdcD8bf+VjkPLMIAvUuwgyfsUb89IE/+R6LFUinry2BGUh
9jjd7YgIMKkOeShcS/V+oPOZOXO80lhVSsYhF6/xKbA6JIrx8qhydkSCiqapCZOM
/NEa93s0wrUz/3i+oIOvjEGOtCc6tF0/JzpkO96j2CKiwSC4LMiO49BsWBUDjdoP
oSU1b9kkf3fUCqpL0yxRLXtVHwoHNAVXpGaxvF1tdxKOZEvxk5oCQQj8mpcVlkzS
6K94sb1TVZejaZ1LgGhBek27dQipUlFc9H1FgAYDe0cGAYg3YNb4/HiYr6JGQTfL
MZmWlB+2A2GBPMkLfGJ6lSXmtgwLwBTCpLPxkSgUO5FtTqwWv/Hkd75VK46qIedO
ZedLK07orQV4JxTaDsvQZOyj6UPax1hIM9Q4h2HTRB6Vno4CffhdxGfr3uTdOqdh
AEOY3NE32N4y3hDsbsDi4cNhytmq7QAfBcpgjr+TKKlHf3V++kZzzCYuO0yAd8M5
R6KLPDwheVF1rtT54USOepwUEN6Ws/IqAwDbp9HizHnIpHy3qkb1TEHweTDnND5U
480fK/bUtXNn6BIBSUdOhGaRrb7kiyiYgorm9qTE5UX/f9BiYac7FDVnZlg7TMQW
83Je9EfwVhaxaWu9K9vbz4Zauy2Sr2M7sCbc7NW+TZ+9hgZSuEDT+0IkoBs87F43
g5kfF2Z+lhM0FWgzYIxRXuorwqSynUUlPqufrVwSmIh1JBOyXtdePdv7Mkd30u/6
WlyqW5+lf0AQ6gQ1zZXit1SthayzYZMv/+ZjdhcAK4WaqgyGPYyrY0mj3fBO4MUu
A96H/I0NM90qakRaT6hjlPKu5RjlZiwHzaqf2V6MjiBds521dLH5dfi2/x5QnysK
6A/SK83s1zgf7lDXBlvp54ow8EGWjFjfBb8/duKeqRoabPj5/kdAICc9PdMZWvhc
dog6zoLKdAmlJnWqrC+wlIQorpXp7/AS0eJY05xA2b9pbbrpDCMZpPOiAfenOifE
p+jvLRbZ83qBI9rG6B57LnKba4hce9iZJEY5REnF+E2+DgPOwEstiY0z0G7ropZA
eGHubpiIfaoU/UjXKa1+Cd16XO9Ks0HIIVAr5uLGHmLh/eB0DZa9sPRKilujYHTM
bbm+tXav49+jC3Kms7G0aYdjnYyxnoCt1ulLEquwEcPRNksvQxXj5db83euV8+mE
b32Xn2Rv4mRqx8q0gZ1pzTUpbJiB1LXSvzM893fqywelQoDYeFuUPGZYj9TCiCkd
boXM2OLeTS/eyM8Zn+z8JYZo5BaJUTxzmDn/qqAoqqTlHbRlUZvDqqjLxh65TIoK
E/mhYKOjMRbkHqo5moh9tQsBCmdwrynX1mnCLESpGFQoO994J3f7cm7JBRwSaBOI
RacSDZLlWrOM/VW9dMgHTo6crI7bvTQo16sP+IVrcsNCmQ/B9wQC1QndZ/BBQFkQ
vlkMXCivXkH3CjpF3Dq986JzBHzGqxrm0VTfE4DqiXMBXmzwwQvoM82Bmuq1gs0V
3m18eOp+cEvH4uZE8+0+rv1h1JJJRj+hZLFue0BJtWGVy6ixA9Dq4ZJ3uz7jSgME
JR+fvCPBgqpT25wfiWN92NQetSaOciMtMdN1yUizFgLA6Pjfmx6EEW2TcqmHgZm2
Tc25OtTCaT+m3+7mlISnB7KmfyftKOyJ80ZFg4Pkp1N5jWXJzcGjU6NEGqd2lx/B
39z6arj+g/joU+KTTM7YBeSQYzfT3/qMMiRfMl51PlwnO5gG3B3rgDg5pfamgZgC
Un77Xv0AwlZ97qBVQtTXp06qH3vrZnHMtv97dKQZTqfwjf6JeSvax4lZsaEm5Y2k
mIsSwr7eRcW16/7m1rI+aIzx0sbtd6HMh1h3GlH1ahEUAKeL+EVAavZ8SAxpNeud
98gi5T6j5IKHXC/gpTIOxTqakSNu5nWGSPls4i3bhNlQ02bxeLF6QI268L25aznK
ve8jmn8MRuNKlj686m390owP4y5j05hPHsNcX+7wcyt2gqpnF+USABK5Yre7N4ug
jdoVhkXbtW+a31t1wUev0TF9UIXeSq2aCAhLcurHkM0gCzYO4rG9SAahgewgFD4Z
+VaO1PWsYmYA6f4ckqj3T6LEFoBSnSZIvuvY2yS9BDkmH0uCBNtlvwvQdw4LBviZ
k8ftlWjo9gHKDNapucamhw0PNMFKcNUgtFIRPtCr4lv9qWtvkr0eZ/rhd7W3UADv
hhxPm7WwJ89zM5oTUTFXRBv0F8MHL4ACDFZBRwvqXMGA/H81gwoBDmMDjZSFxEaB
Ck41BPuC+h11qctnTpEkY8MGeYXbaHJdbiB1ZVi/a6umf5/n4XRQ689gGRs9y/pM
3jp/lP3jk9KH5rFT1LPgDLZ6k/g30mH4K0TWJ4qlmQXuITYCJW/4vWrRhwB6FD1z
wDOrEhxye6gYlUM883liG2uRzgFSxJI8QpPxDxB3JEgZBMhkYncsj6cCkOR1x66X
QH+wFZk0h25898KUPyPUF9GlNLH79wCZb20uOIkgjJ76XA+QOQcJ1AfKaxhMYWC1
8ZZma9slOpAEkLhlfpvObosUB6g5G9a7tXq0V05Al2dFEk27/puQHqjj/ra77bvu
5ZLEiR4MgTXOh4pXVKFBU6Fm9lJl0nL3mxTh+8fr0+Ox+nwCT38+qxbtZo0kPqAT
FfnN56glcHUrSko3BMh7a4VPlKsMRvVBWbZ/sU5FvwQY9JXFb1HBzY8aRL0TmzzA
zGLPh47AfdlAYGaxrZbbyhuSlKCciJ+MspmWev7QlC5iTASHlI5d8SYmtTy57kaG
2PDjMOGzTW+Qowl2Gq9+CspA9i9cDk13bnUJxZXKWsygcQSRvDox+d6JUcK/y6/w
8GmmWXbMi2oxPnBGxtWen9Lv/K71be+5NlX4DqSvww+PeoufGvjnk3RZcVFs8SPZ
x1pKOoidMlXdkYuRGt37imvyVJ9yAjhKnYtDE6XSazti8gkqSjPcKzT5bDLeozvr
Sh1RsRoadiO8kYpg8WvZb6Io1c29jb4Zm8AhLvU7LXDD/NDlnrHzIBse774+Iktu
CbIgkqppdko+/VbkprkUqO25NtdFpGTpln8Fz+iGufEMEPZhO1fWnRCFnUm4N1zP
XF0wkw4ZCUlgLVrhHR2vwZ9nEhVxv5GsLvHpqKTzemRUoqvheAnXOy9/zq1NVdVK
ldzFFAkvx3is07/nQCEG5N2pSQTajUPTG9O5fz9BC09QdGwK50SL2pdp7ul+oCa0
L8h6kRV11mRTOgOJ5qsbqj9fBsvQwCp91DWqegVFk7R47Fx+7L5nSXprEF/vv14h
ltX06jzvPmY6Mj7chrz7C2mGFMdrljaMuoP0a2tpbwZHmzPKm5MLIRRyQwZR3juo
9npujuyjVzOC/fiEP1wyK02wG7DrhGRxFSdY4uPLuw8lfV3g024R5hGaepTgF1aD
3HrxJEyjYBr6Rpw8s258a8X4YmFmgqvx5BeOQZp2HG0frEP7py7hMVxyTGqEJ2zY
QKgQocWeGI31ekbQxzEVMsPXIONl8eoaHzsxXKEfJcYIlA+IWH0zh1SIRsmdYKGI
vTzTpla3HdDc7oE72y/v7s1JBQ/WSiOwA85c9BEuZyhxWS61xmxXEk9oe4rFfTWh
7m61rlDOlgYfiIKseJVQIb3KhxZIDcptREU2Q0tOjHIgO8sxb9cSh9F7XMozAefl
Jm36FtbuDTTr311yAJ/yzdkV2tDMoD428zFscbCSc9IqLl4qAwEEqmoEdwa//X4y
peLNugxmCVIUEnRrQ7xJURUnDEgsYykpNWPX4ne7xd1dXEe/FX9+yhr31+h6bZaA
NLFPa5ygkZ1zACV4Iby7EfCMSC8VZHmoO/CneTLw1KyeI8gIW6rWTedzTEC9WDpG
m56Lr9GWUh5gPyatwWpv5ny87fIXt97EPAbzfXesefTaZtfUuLjtRcBIzcrApl2l
uH4q3I3PoeevdmpILIX/ZsObFDJ0jAI4/bf6iGZmF8kqaBeM2MIS+ZtM+8W9NUXN
WUMaX+AnzMdF7JO/Urn3fbDHPIjVuZlcY21FnM2bCdSt+02FJL5j0wgSh8JQXho1
ZzXXd50Ii6mOODbP5gZ/OqTDXOtg9K9174GD/+wVy9YhugDK3hJ8RIcxwGqMZld6
DGNB1PnbOPncF+qbEo1NpGko7UKYjp+DSbQjB/CoKqGkdI+EJGHoQi12t0Y+u9ws
2xCPTRgF+xVVBvIPMbG6dLtsckQKPwc7zpp9L7YAG5GMoTEXZ+RUkbOK5fnMDfV0
wRCxOdg8Ne4MovLalwfNZj2zam8zWeCimKuoxImGdjKrF09Ln4SnivumNvVCVzbA
tfRU44bBlsNCLONyVzAp0jfXsEiXqhzueOHJUAxThG7EeATwnSHA8B9L2EotD2nZ
uE9JeMu9hLHhumK9ilpHYfyZOBxCr66TL7GN/XTiUkwNCrqtFXPe2M6cMr5NTxu5
tqRvGjp7B9EhmGqkIfPGCKQZrXuKGXZLSU4r6SSmi81XM8AFCCtoOVeXht8NBh9K
2BmQZ2h7wC3UxeFCRU+Yocuf83PX+FOfg6yiVDCv+VmgfdlU3dOLDCW33zuzViI7
o8pTll9ZPp+/zaTlnIfo+i17nAG7AP/+vrWKo8exgDpK/6T0V5RDaGkkNVmqqu4i
9SgEbw9Prdf34kg2du0+4NOAYlnZ5UifrWsxXYzvVlC5JYYvzKTAm+8th9yZhT8r
7fOZdhGBUz3giAe75meN5O4GnXkKxI8VuItBNZC4iCeRrnl85lcY3yqJQPZHOlR/
bBNSdH8BnPdyHen5nIeSBNu4utr2XF9YDWoGVKuu3q7cWMku9XSpjneammWObowL
GcmS+DEustgA3yP7Dms0LwqksourcQ8M5obEyH1VxKsQ7eBtekF+TNhMGz3GIWwN
fNP1wYKYlE2w4ltqd5cZGfkFZtzQyLVoF01y/qdXvHsgbT3a2dEGCK+Sn960lkwB
Sx7w6eKngmGfPggJu4NNf9wpI2VWMvCxVg3URcEOli8HBiSO7VD7Z0HjmIPwB8d8
TQr0UfEuAAdwb5F9EJ65bdz6TfL/W3bydaK3d6+zZztO22HBmATiIrw61SJGbslW
z/9+syUkCNQw9YMIOrBhMAd5HL4FkW2cBBpfhBL2/Ei3iWwi6PDzWxjuiHFCuuKd
H5iiAAiLRqB0Tj58clazWqIkVrppRK96xj6tBCR2/l9/3vSHc5kR9FRyGs5lhJfM
WEViAs57XXSFOfAVjMdGZVgKqmTzvkUTMp8S+xUGKKsK/+ImVjojMf41jov4ALo4
m9KcqmV24sUnnrhQVD6VouND+7oX23OBz5czG5VOhC7v1th1wJ1akzGSpF4KqUM6
WnSEWCAF56l0pkolEe7D15Ug/48xcaLFqbSbsYcAsZobY96z/8YWD+gDj53d5m2T
9tBwBHeyUBs4/4gDQujktP3WlYuGBTH6Kz7nk+LqOCLJMyjB47vTfOj6/3bhQ0vU
LuWyWDbF6yj4fX3F8ncbNtsccwiKHmUmDizDqe+IDeI9derw61r8zu2rnSTxEYxt
1OQwWt+3P/99/BzyEBfTglunJQSXfASjlUnH4eX1EsaCXDFM0w081KX6pIZZp3ZG
khinUNAc9XrVFBpUTLViEh3etedvhEALnwbMhTGa3vmH5KwezCqItonXpr5YA/uk
ahqrkg2EdkQ50lBLs0G/vul88NbyHQ+Y4q/nmQZNPqGbtuRc+V1fwdX1s20EcI6c
yn/+UR9ZxVc/TV3Yx8qiiTFRrJ16eI/HYxw34f5EQgvqqNUakNm6mcRuqmFudPqY
FhTVHWyiXFORMwX4xqih2xp0K58jAd/6iqsef/4nupHjls+A7BBsQgZFX+KJd4Ql
mNyrZJ4pSX7EOKR0MKcMoQz6MJ7vQw7muKD451MRvLtuwOpXo5YriD8DezsdJOHD
LCthu9crXERoKs/GeJ311yNGlLQ/dy7dXF8d6anR34N88bxXljg+kfGZK5OWtoUd
BRvE4CS6jtTsOlD63cNTJpRggZJ816eZhndGBzFhSv9ckPVde4W7YQ6k4t0cZAEo
dklsrHWccUmirUar1rHSOi/jw0IyycHta99A1A/0Vfdp4v+omvhNkW/KAeBt7aVC
0zWWibsAA+Vj32/Ksdh2wMK2UIrOxbr9nETd/FKSJmo97OVXC3fvx30JAY7UarJo
YY0NGCOYfQJ0OaPGh7qWiMtF4wnDwaq43ixzx5i/4D5obxMUYHj40JWO5W6YLsty
DazHHIjNiqm0RzJ4+OQ6xXLMnmW9n5NcCUoq2Z9y5giwl7dZvMOpBSlmAMDzw4Ef
lUlKUSAMmzSeazCDubOFTT0tX7eoviO+8Eh7bo10piAkBaQvt7yM2oqxq+c/GP4O
pTW/vuYsnftw0JKBrqO7iBLFAlnq4fIYv2zlkH0Ef321whIXHcermTwvfd/ot9Ku
FjUt3apbhtUt/ff8Mua4Dqe92GpvVJgqp6U2bS4wRJIyg62KP3xJiqW04HwlX8Kg
9/7qEFEgbmpHQ5vCpcJhP2/vyvTcC15iVOLS8zX1TDGsbs2OHLHJf0imfvHVWpBG
eIQogKUTlXB2uhgKUVp4ISoSX5Z5QxENx1wCkoIe3US2xON0Gxo7IujIscWU9jsK
mAwB46jwCebiykGLbI5ghm2RsMFXPV+YorYRp0d/Ieg2bLWVzkGgkK9Q7NrL99Us
s3RfvVbDW9kkWZayLA87FYWgtbPZ8g+5ka7YXCDXLajTlJWWYEBKaOtAZnVf/bRU
A4+H4oZvXcsXk+CqWkDpW9GMNN217BOR2haMFnwwWuTp2azxMRCNaN8IFy/5d7rW
noErehqJA/PKeiS77GUaqxrf3nE6E0zTpwVgI2cS0V46Tk/sIhW0OMnu8vVf9yR/
mjfuX2dynjl+0SeGzMiSMvnAhMGU5Gm6RuRKMVASKs6l3PwJjEpPGHxTnCK45Tpm
H6bPU043o46NxeIrDAK3wBCw/KFQb8LphA9Nr36Twg9ItZd7T6a+qMRPE1KFkDtI
dNR+eWzyT+PKnIIlqVocGa1CQPM+hbC2GSoeNZeA0sH44IvFJRUaTi5jDFsYynGW
+OpfxXC4zQaJosMxkLFSys7s7BQ4TzpZdEgthSgB1tQ/gXx7/+bimwKxcsecK4MN
S+c5S4XW3L9yGM3w0zcMPIwrNofC8aP1ZVmkAYdUwA9XVledoXsd5PMedjnS/GFC
b7zXE13wkQnRU3JiLCN1PPOQor+eVKTbNQbSAYEBK3nmCVOp8q3pv6pyhOqLDXMS
w3ddsZQ3Sp3f2D9J7wyB4oyCTakSg/O+y6befUUT6xoqa3xYJwJzcLBgpuc9/fEP
Y4nQKKAL6Iws4dlH6cjfV5nht/eT1Ab0NJoH6mNU7ukEvbag30ABi9UU6OdMUZSq
SgN3toLygtbw6dqwsI/1xUTJDSU/KOA6jZdMG8rX8JaNEtUd1vwD2bbJar961I+Y
dKXfXdEEl6epzL2roarQBdR+v+zA6PsND3J7HTTquLADkERHG5A0Pb90ln3lxeGR
PdomdubOsrOyLAE4zH2hC7giMecyzWtbpzbJ381g0c39yA4NSLSJ9JUdmGtmyDE/
15berYTfyeqFGVGfsfo2XJxrtxuYECLyIaZ9N2svNEx0aXLfEqrv4EBi2KMn9jI0
YpLilyHTb18Lyoii/70Ap9bwH9EgL0r0r3+tTJS9RbTlx3O2OCR9qOcndFzc83/9
PwH5zYy2njwSxSueZ9K6MtAb9EsBy5N/Bl6gDwbEtHoNamIpqCDa5uwPH7rzfRG0
oNS0kxTUK19vuDfxC2SPA6cJXBB5xRvUsjVydEJATf3Uy2cDXRi6GBcUhhoPmEbJ
KEpyWrI6oHyqLqB0DFd3fLX3hTgVB/Ua9i0r0NWno7TZwVCANpnxMg/0mzdgv1Mt
ox3d/NN9I1YDR1J/y2lHRl4y5/LBvPJxCmBaFOuhiCRQnfxUPFigoyVXxwbPcUja
4XQZiFkpuS+g1iRZFtVZpUdBVxSe0A1OvB0kZumKgX7jI4ZbLiWeGTVLqxC54iwt
EV4rQKF7KmtnMY5q4uWvsznjGbYjjiDjBJWq1h+zwCxFRln9VTcZVeWCw77UAAE9
Wdau3eZDWhSNBoRRB2Q7q+hcOGLB2g5cHLjLIuRtmc0ZP6uJJyxeFm8MpEmTQDWF
H43/Tgr4Cc9dDHQ7XTzuKsseJaZiaws4OG5eQrhTc4fMX7gzPViaoK5toREWGAGU
Np4BPOjE38392KMbezSo3VyXV64mlVcyMgRVN2+6EwXCjWsplf4DwQEx4/CWn9pl
Cq+zI/q0kzS8cJEwYuilOGgwsEL6GYEH5Su2JipwRgNg9nmDWEkrZJq1Fc8Iy+fa
23FmsQK0aTBMMU3duOK9r5jHvxGgg7SK0CrcvxzYseYAmgvuz/QpZR/H6oB2Igz+
KcjV2LmwG9ONInNLcd4kBhO3Bld/FnBm8ei8Rgv4shT+cROBB8ApRdJXDWsgWuc1
+JY1ZKp0vrOfJ/OR3U84vqq2oWGZUmms0vbbb8OmXwVYxFoLMcelf4lbpYGmupt1
Hh3kfQ8ejw4Cx39IJ6t75Nl19RN9r6kziWtxUbNRbpjN8gg4ag5ULpFX87K6i9Ji
nySQSabt9o6VuXL3AEXDGToOfpHWNNvk1BWsWZh5uRF/lRvl51sMNgdoBkQI8vbq
fN1B4+gdijMlr2qZjKQSaJ2uqzbS/q+2wlq/6Hg1Cd82b7kLtNww0yl2kjbvO04L
qCQZL4wAew4ao4gLS08bJP//Upee5k/C9hkj3R6/1yoZsuKkQ8dVubESGwvQ0g6j
H1EbMDFr5Tz6yC8q5kqXQWSOFa8NIUIwLaS6RiWJwVtEZaAcANb89dJeloKfkRhJ
9vJDWsy3uE7q/pqhlb4WvrygKLe6c5VsBc5ArwmUUmaguUVANCf7u9t/8yPNk/4l
9C2k/nXFZ6R048Luhd5gguQFZMx/WxtNtArrFgPjsUV3Inv2igWxNRrXQrIBkwyN
jEYB6SgYzMd9cDAJKfhF6yGCBH8PuzNGuQ3Mkozuqh3zR1d3vJYiLs3aF8NU4DtY
Ynnc1OaWPHiqdBgxFPq5tNcR6iUi6FtK0vejCDRw/98C6nL5QhCz+Iy/M4F8pZq2
rmUIwfhGaKi1WsY7bouFwF9Yxl1Etxh3kakzC4K6EXGntIbrASqsNwprme1P9Hx2
8jUt8alZYtJ5UkL8K7UP+f2Vr3HxIHM/uYD4DsMuaEQEsYA3lOjq7yL135F36n17
yvSziSH015DVXU1ZaagGnrGtqSrVUm29Q642eVm0ATLN3D0WTY+dyUb34aLAZ6Xv
uy/5NczjWUuP7FZPNy6sL5q+jLquwXa2zGB42F5SQlBaX6xf+TCsTEFU/OU/tFXA
ksiKdtRO3u+/bI0MfkU7mKU8MtxqvvNLrb+pk4wa3nUmfZOvRoOdg+MLf/oi9eye
V+OFSEr6novALKPLDL8XBL/vQ8/l5wfYn94ToCRFL4an7Vf/cO4f5j9gESHolWFw
8yhgbnMLwcwsD1XsXmVn8ai+mRctjZS1DlcHnc7JMYDb2sXckO5HAI9GMeSFSJzQ
ViniVRnQ1fBntzlH3860LgcaPA/AbfMN6Xthhwlx03p+iGpXKXt/l5zdkc4UqvYf
li+7tnVA7oo2qBo7dCxRUeAyK3Xi1232Rgf6Ont4bfUwoYKhQKXRYBqCo+QU18qN
7LseZkh4TFVOpC+FbAI2iXjiMva/12oDQ912uhxEDsmczWCqVgSBb6UzZFe3Fzfu
wIW2GgIK5TwWtYKiDN4ujqKSlC02puVdDPg8qQQnNxCzxbtxNXR0bgAeRILLnQp1
ol5IrHg89isH1QauE4Enz9r7gjfaJvkM3a5FsXQtG2OhvqJeLU6kzQs9u949gvDN
iZiUCU+LNJpquSNN2G60GSlpjq24KwJXzw2WtgxuXOX6QvZkj7hZ0hmcFOlphM3s
eX+Zr/uCq/ZROSLjCTNI7RnsVmCzquZ7tMQqFp6BVFVyPiSmKYpP4Fd6WxEzjlYt
rJEI7SbkdtifEwOyNcG6odSHFDjOWB0f40zaH6bMlW1ZWQO8NbCvOj16qqNp76FE
76skduDL956bmRrVtmrMtNxreAnfelABRqvAxqHjnCinquwSTJ9W6lxPx++PSQgq
4Arn7+OVDiwS3UYisK1T9AWF8JmCmcnffbwL5R43EJc8H+L0TmzG+K1bc8OTY3oA
dU6Qg+4XNTB/QrGNK0Nnc3w2OAnsPT0vIhxuyugBGJYKQtuIwmfHmu0Gy+EqjCx+
9KYU8D5KKsjJKpdDxZTJpJQsHR7Gdulo9camIZQ+io6sh3POmkmNVFVNV9br9ESv
/A5C/iGadzZJQB4Nj8zXMJluVton+1NWgUFkiODX3gO1VJkVWrv6lNRfxK4AONrG
xmASdqC+P0AhjzEsUP/8hr6bOo0BMSFmrSVsClWXjDiA8EoShHQAbjemf+u4+elo
SRNtATLPW+CsuLJZlQ7e8ffXq+eoWywsGYz8lMAmF+vSkbLD5zmq820xTgcgY7q7
zQP/BTDvmykOZiF6ngyW2YPMH0Cf49n5dxzGKqQQ4h2P1IJsri/wy0AUQVhyPlMn
MeOwid1M4C6nWVFNUMIv08HHCNsdyaWDDf4pcs7gTe/Dis3XhMS1FCaTiy/Vmy4b
/AL1/WDgOY9eoHPNYSVOR4TIFE1hMwFlW5beyVgtsJEfpuRKMBvVJ5AOOsO7EesZ
BaQQklEjCaZmKQBID2ylFrqwCygX6V0g3G8BFVtcT/kx4q/3shajs89vThy7hb2B
wkOXVj+J+Wtydb7c53nVpdmFUi66nMWJf86u1qGUdxXp51OrZwrxvw94CwM9g2oZ
b0UZXqed8WfXAX7dZXjw0jzewUHu4pa3pin95cS9WGKWOcYBfRHMltpy7QcdtxQs
AWDOcGcVAV+iPLlqZYvcYNIeEzIMbkp9+B/HScIT0DPpVNDfHcLtykxWikHXHtb8
XfZHhOOvujsp1i61RnTM66vOSZxRP4qlqPNNGsFGSYHQeNgWskdspznm8A3bTrIs
lC+TF0KPxLfO8FX8ggzVOfIx6XZyYaA0NYBTWmnqvgcsIevjPQIedZ3qL1PzCwBO
JF3xs1sdKlgSFv+t4iQ4AL1cZMdSUv7QDLCW/GfmlM8MvEwEICYA6GMutp9cblEa
CgOoNn45dkreMmcA3i7rmecc8SIhWDzl0qYJezFBkz3Ev8QtaMBoH1CQ77WM1tG0
MLsc4ckaM4gsQmBR3ilgJceum6HQ6G2fhqNxfm4p4wa5Z1npVqjWX/let1vWgMPt
+RRpBYx+MDK1/F+/NKjWpB7phmuu0GFS0w0AORUeAhfYgym6Px6zzAtfMH0pSjc+
T/pGJxjF63lk8Ls5IX4Rx2HQV3IytsHIM78s7zsGFA1hRgExJZRKDdhBEvl3b5ta
n90HD3v4B1fxySOBmyoT3dIi0k/G1xAPX/CbTNGF1P8zTRsH59XKzPt0xRPQ5P8Y
VejkF5HOHXlv+Mnv2vLF0lER9TRdDyPKhpSMXQgXck7ngaX3onkAPTdq4F6MKdTD
0W3GotJpvtYI+x502ZzHKY28ajMCvv6C3DNb4ccoVPgCfVzWMobhNErPRS0EjkT+
uy6oUUiBfj0ssKcQ0z7D/OB4qmWAeTUYaglKLe85Kcf2aHVxss+8KgP3wxkxUxZH
FFwLyU2GqqyO6nVAMIIj6YRyCcmDssV1MPHl//U7BuhTCc4qx5YhK+BMMxNiDmry
aES/1IINBGUMQlxwx60z9hCnDtfL2MTy2iT5Ijg/pKit3QhwdBTLjRz7U7jUDXEl
Xu/yFlhR/0NUOCr43XX3sB5gV1kI7LCPuY1SQj7nfna9eiPmeDc8a26Y42Uf4ykT
wQsv0SwLxyRl3nwf2dyqSprcpk5VGsmEkVaOqsBc6TOd4kHI/4Yb8dvorj6MQrOS
Pr3zAPcEqTcJPWjqmMjQ+wZe26l3QeVFJIkGZSHoUCQc7H2BU7gKQMrFEKJ32BV/
2msDbzhjdCKbc1e0TyafajUESgxUtiSeKf/Feu64vxOTLxOtNu+CCKibh3tsFo7T
OUf5L1fcPIo6/9Qnnh2eI6aqc0pIhGqk54FIuIw1HMKMdqvC91uQOFzLYwGlx3S0
efTd6wQww39CajY6n9JN3wjf9IcjpwMHcQ3w2p9CsdpQgngan2ZlYRq4nGzsTGjT
ylBv3mm8ScRF6o78xrnznnqlXBUmGRLk5JMpvV+ROqDxfDdFjE9LSMwszWjIgzIc
Vw/aJpbZMWa+fTf3lov/JCZ0PDVXic8ptMrQhaKZv4bawRsHYvE1SVaGnGyXoK9x
ZGY9gEp7Ll+rVyR+QJGcbwPxeneFGvcAlA5JkFuHVrg9Pdf8tohnhvoCTk205Q4P
/JyHyjK8YNN+sv8nUJUkJ4vHqDxJVJcTuMQjWFF+P3Fkyw3ezz37f6/NNNzJVi2I
b3gMSZh5dOpEm1I8dLOt3FPkDpDM1LaMct5GgfDgbxu+qUkqC05r04Hat746MA+U
x+Pk18HWP3Pd6EiO7vB2q5Mw/lRHbXmQ2gNsujbYHEmilRoPhmf6i+ZJJYL/yEQb
dbpqi9PhSTfqY0o1fEhs0YTsQK1UfsCDrgs4XIZ4nKwNoP7P0JWsSa14ScsnzI4y
v8YN+YJgyyqp8hBvlcvUMIbi6byqVSVRSdtyB8Xnwlg/n1ikz84gcL3mZF6qiiPy
OwzFQn1Ed9picUeD//Gy/33qdZbX0CFCmfn2BMcG3049nZ7h38KMHJKoKWtZMly/
gcZfGT6uc2tppmD3fIiMVhDFu/oB6kic02N6FJ9cwCETGhnEDXaSnpyi60WCdSfW
FGPL/bjWAFQJ6fKtiQqr1aiJ7hOqqQAct6FvZMyJPF61UXWxabVwGgZajt08d5ip
TCp5gdrLcgB93SMENXHMHsgqfJUqC9RXAcSGM51gdEBb1jGGRkUZTpnz0FdND4K9
Oh9GaiNzbBo+b69zJ6J+zY1pdEcxwosaALFzE4UMNOEsKHklmDsO8VMjnq66OKsg
NrH3PNt6B7BaP5RroOsbYuJbJN6r6KhyxFbUumQBwonJK3czwsXRSG9CiOZhSG4y
8Kv/b5+ffCYKYky1YpwSspFCvw9BcoMHRuE3jJYujfHpT35U4fgx35ljx75XNxme
HXJ4dUwViA4aA5XxW2MpB+RhEjMXK39KWD6h+eSTzjEx+RJbMXhigQ8eG0LQaKOO
Mnc798EZzmNBcr+Q1BQ3QT6HPpzdUgB+LzHKOKTzlgUdPPbNAwcV4el9DWZY3dHR
efZ39SRYWFtEN5dFRF2XexsvXNGBHPo6sVk2wZePXCf5NXW4K1uHxcM8H/WIC8z8
Yi443q5xo52VX1i5s8nqAuQbBnxidOinNWowJMffar9GCR7aekIMzzSCWPwoIcGs
1c7NCt4riXbJ9k+0osk4iZ9tXW/93H1tIOySJrGPTp4UiQrvD9Z/Qk8NnuHFcqZf
yOnQs4eBAD9Js12MeQ4pKTN/zj0JayncDiKSM3Pxbaalrn1LeG3TbgIbJLfUJa5p
dob73BnA6dI8pEVjnqsE8Q==
`pragma protect end_protected
