// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
EvcYVD4/vul8+7+RFAIcvSJcb73Z8C/swkv1gEBU4qBgfPHbk17ETCD4nTWEoaxNGNsQ9Z0K42Q4
rWjvDHGHjR7dc7iSXG9eSuISzYeKl5nU3jaJMQDvZBhiJ3QS/d3Xel4mKT9n8anAsm1pYgRoFfaT
aDwXXIsJCGYh6MccLSk2F2sp2wCYuRceUvSTuYMzQ3LwTR8UJAA2FtegRkI+om1xrKcqY72KRAmk
/6HPMUNzm1oR0hXwCrlN76df86ayvi166RMzktuPyMY+hu13FCI5NAAkWhLwnY0OnxwGXkwcp2bE
qH3OAuApt34p09LtTbGDF+HfQr/KfWOcsncwdw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
eYiQLFga7oU8Sx6kmPCabZpc5at6YvIySvHl+NnoXH5FLPh1sJOe8UeGTYFF/9pweKh3v9wAm4Ah
r4tlFB6SdYeKnI56mwSaY3JvDemiU2Qlt5WS0Nt9HizR7T3Phh0SK3ZvOAzO8A978bXnfxzQfC4c
tEwBTqn+Vhq/hv+NYqlOnofxX3tt05prGFCuwWNl7mMkonLmqFApcdHOlPYIMPv0bhyfDxbmnN7x
Va9OIcFDEDpPbhjtwhc4U9I6omSL8JRdBjw18Ka8mMz+a39zZcoWwl0D6HafmpEbocXFkBxUjqqB
mkm6rUdSt/h6xqCLdL/DfYjHSqLCzL8w9RnsI9uyz8WsA4WUk8n0+k87L5ytzGG59l9mbA8XYx7C
vkgK2NQEZo7ekLMSd7FbJErIylfAlgExhTbTzPglV3R6TqqIu0vwxZfDxb0kD2w1ybowQRwGsgE+
sel6QcLdR2WupPGWlihYExW4tc6oTPWb1qgqDSMquoyG6GNUDrY31Y4vpsjZ/Acrc7h4q83XOAos
Q41lLmgyP4FCzYNTNTbH6DlwuyavRIIy+7TtrJ6xrHQLhGcajPUsWFkruZh1nesuuMxb0ax7zEeg
p+hFDg57n+6hxbBc76VNB/31/9Byf1DJmkmWk00VegthkWrGnwsz6UF0odCpB/5jD0DpM6EWKcnA
F4lewrr+SojL5qZtbasdr71NoqxZfWN6z49vvSonAVvsbKdrOQVJwHwsJBcxeItfwUXMF09f7GYH
2C/O4JnTtJ4SgJtAPtdGNmt6R9woERjIlJBJQJjBLp9eSpewC+TaiExyH8G2gWQHwK+RfwNZLsdz
yI5xJxc9hbKBdJLgv1A1Bv/M1MD8hV4AIQ2i/Z+IIYhFUtAZp7vXcNezd7T+2Pkx7GwsO6GnQ+oh
5+zYbs834hJwukppWqcrJq5m4xPpPjtwx2y+ejYu59RMj0719gywvfoKmGTVKWVyTPs3FCZKfB/y
SRg7grEWvuASVjcuAAzMd4Sfc2vIq4IeG8ejdmTUxhgw/Icp1hV2P8POsDETbX07lFCP39v5MAcg
oF8MNk4TXWFB8Vcm41fCBoSFAR/5OjWNK3wt62Vxqop+mLk/HVGfzmsbgVcPG9Rfgv+zFKt9nNxV
xgtbq6FWkSKRMJW8KVlgbXcpbMXPcVcZEX9OPX0SdWRNoaNQDDXs0VtliEEBH6TG4u0m8TYl07a1
UPAn7YxqWpQtpx6f2GLFs6fcPQquf0pgAlCOeuImx7vw7dHn4DOZYYU1WLuyPvaeYsyz8cRRjHa0
8LGpT+Z5XkikhWf5v8rXYdwa4UPczxGeeiZnwwh+jm9+jJy0q0MyjAhbIfsC9seh5bIh7cv/1pfw
CcQ4+smZwwBl1jUb6tISJ5ZwO+Klvh15PQI7ISgaIeVgTecmH+Ns/DoWEunj82CyRsUTl0N5jOTT
09OmISMdoQVFphbjySNztZu/mqrQ3iKuwmcMUzagm0vWmRpP0lpTlMJuL8TkXguI1N3RdSCRUHhE
qx5KmSh3GHbmIrip8sRdTmBqYkcNleY76u/96NtgcRm/lSnGEYEvZA4ZbYp2UEPokrCUGsstR6MT
wFYqj4w5CZyuIUAcssxqnFDTriamrJla3Jw2YuBzTfZqfuq+aQEzjpyi2Bv/+tOyW+UhXZ7uYKro
95r9TwC6x1r48ysdMCcKkfJKcFrXpATxPljpcoh3aVhJ4FJVnbV8eNHNHzCRlc3X4Kguun8x3He5
rwM5iAqfmbEx7ap/fhxMb+JNTYcL/wv25xmwApz4+khz4Xko2l2i4b/wipOgxZMcahULhjhSzRuM
oR1Q+ULUSDiiM24fcsLhbYM+oW6zxSPDDdQMzd2XSgJ8NPCtacRyv6d7lZosHGfntsat2FKFEIhl
2TDIO9S3fLwxeiFbKCSjgBzIPa+2qZ3V6ys8XSTTvQsBwxxA1XcDdBp94N4PKSJ/J10XuXSdFbom
hPUePkGptA54mSTn4CnvlTL4UHGpO0TJa8Bhd2oSvoCupR86un7YPmSr9FSFeaxuxfiw8v4x/cd/
l3c4Z0phjYcOdfZ2lzTx0JMA6ChW5Er6+NeEOAG85J8kCt7kULn0eyxwXS4f1pWcL3Sns/IfcGl6
P7NwiZQU3aqUJaMbFBgBgVfBFQdMpAUTw6dL+AGy+o0sgFvXMqR5vwUxQGOKN9vJlMej+5Er64EJ
Iet9ouHelQyttwVnaO4TuRno9G6Vb6U/z0TsBooIC57zgLLPWv2uLn8nfQwj2juzeZ4lD6ULpT8Q
50TRQNen/OFLcNtyEbpt4ihMlgGy+HSjYkfJyzuLZ9RTjpZ4UMq20/nxOeHQuglECx9JCQHUShyn
Zeg6rUnqWzMzsfJwGO9nZk82PHmBmfhEegO0ZkveBO6vIjWnD3AJNNNhUFiV2wnijXNDih1Z7Jmx
zdeqdBt8pheEHz7YGE0SnYiIbZ7TKX3mCjvjc7K5CzFZGS7SJnSBCqqPdpN1rz7tYEt8LdwVhNBQ
nRcIsUgIPYnGtCgiGwgWMTzxpWGsc8118T6TXSBPtQb8XNXvlf025788CpP+FmwN8NeFrh3x2BDU
ooha6veJAElKcJLD7nfIIb9sEnyiaZKxDiTaCJ7r5lgc2jHKmIQ3gVjZPc5IOY3fZgzYpYOzSdQS
yo4Q+LlP3MrrGTO7oXX4JfEANwvFMCLyh+T5rEQwoCKnDSww5dZTj/FQSV8DZs30IVKR70GeLZTz
lo+c2bLX5qgLjcaB5vosMSkSj4GADjMMAkf5xFSea4I8+bIiFGkDkbM4awQQAXv/49WpERH+JL1K
2HwL7OqP6hdMlKQM/zRe5Q7V13QKhRmeHSXlLeusrTvwXCFp4N0jX9jwD7vnyq+4xb6eQ0Gyg8fT
iAkEmtsNEmBxwsPr0/kNmkHnureh0//S7ykgPXwLIJIZcz/K5McFK8qU1bVDZ2Uara1WzIJgj/bA
JECVVUsJ09GQ7GVWIte39H2sGB4i6mlOlUTSeLE1f+tpOqFFs93+a66HyZj+95AtiKazzDknxlIU
B9DRevPgyVjXRYNo36dCYSRPvVkiYbOzBvbFC8HM/hPmnCl9kKPw0FC1NyysAv/pPUv0iVdnnqle
8nqQMe8+LUAi87Z4kvBHHyG39qOcc3T6coM8NcJktNnakOqLyAoIAlJhXxxKXDdDLPa8rg85GX6I
nwPgkxJHtfFgKF5BxkbsbeIr+PjrH89ZorSuxXSznBaGq/tnt/aj9RDcHhKL8zD4Hj5ryrnxVa3H
rMCVEBrDbNEiJVCzuGqC36RW69z7CdkugdrwWMh3I+LVMjcRGomvBmKtwXQzehW1mZPXpxssRpzz
8/DYsZdfQ6qIaLymvTQrdpL/6B2KPLup586y+4OqnxHclp2jMAHvqAEANIvJQ8cAAQYxJR8Z78cM
sEdRjn76VZVPc9efCqIFRjg9fOA5KKc3cTGfPDJPGnNMrxIQcicGMXgXJyVVS1DzIEqTl67n99Pf
SaUD79q2dd7SJ0IpYp3iqz9sQVtZBVeh156RS+UyxOgivPONjPr+MBgodJI2ujIdzAUjeQnVkWmf
JdImWn8WNlf7+vsW9gXlvHtTkW8zSLEoa6jLfFW8L7wyPhDkFhrA43jgddT/jNVLw+RZWfVC1FUm
vfed0def4Mwq75g4mXCXF2CUmDYfnZR2RJwIUE5+rf/LOes1RnT8mWBddLrS3iWTASL2T0QLbXWh
vdYk1Zor8G3tdmxcYiaQIxr9PqKfAJ28qNeHbBfD+/4XvtHpS5b+goKyJcjJw61TW0uS2M3NpJ6Q
h93h1dtLpz5rGzJKWxrwFETDDcNVCu5WEt7RF43fo+NXi7PwtFoOS9U+Jt16PIGLn2b5mFMBobXQ
gc4/9CPLQfaVm1OHYudHWJ3s9ZepVouFypUTPCsyOlzl3GJAUx3ZyadiiXXF0vBZriyydGmOtzui
iSXqutVFK+bmX16dFkRVDJL+elO/z7zhEpj+y6QFr+JdjtEADeX2XwIXRE/MTjWPwhh13/EW4IcE
rD75nCHLd6BX9xmAjFG4fOiDgW5EH8isuPO3r9EyI/k1mlcGEeLKUo70bpMzMaUIcwVVJDovf/sV
yUGBYU3zBm1NBmlJhuV3Hxz8tp/L1cJiyq1mtlmK3ysfoBk3/i/5cTr96vo6enjRBkTxfSYq3LQi
KAW4/1P2yoOM4kJFFcFuSZsE02d2/3NsHbRPG4zF9TyY8KqIedMH1XlSJzCHEOUwx8U7wC87Fs/E
3Q8FJmwMiWPmh6KZfZZVn+qLdVQKfvKWHx8+lmP0uzUjEdXxIGfQImXL336mHGNmHw+k48G0a5md
O5ZLkwxsCChcqj+aiJFb9UYlGJTMtn6dY4ZXHv77gidndEhGmvdFnDCpYtpa93pc+eSI2YJMxDX/
S61XBVAr5wQB0YkwVHADa6qOyT9zQTqiYPAEidobhF5tYY7TSej2c6rPc9s1jbC38gazqrD8YgoW
ajTDnhzHigdrgKFBPzeI3U98YgwH52QzCTxvoJ65kxHYr9C564RVz6uZDKHea75HJ6jIddx+kvMA
4Rs7KF6v0FQpIdKjV6Y9k1wlwqjx01+JFcP+v8syrCHSifmUu0EbPXx6qGOaUlezIne2chFVCNEX
GihJd3Md8H9cJhk6Iy3FFtpzf0HQUIuvrbC67SzT87GHLJCez61bdM/oflAV1GuezS8UqyRY+VBb
PXtoALdjtTUC+8nSIngIUYqLpiRo7H8iLCnZ9lumBX7c4FpD7juLgkkKohRE9cbMCOEj12SeMaf2
pi58ls3DrlUCs46qPpqhXdiiB1lP2B/P3shA/kYgR76rvbi3e+s3iDRaXmAz1Mm1paoYqB3s7TYo
PYjH3JjA3Le6Ttrne6Wb8WZAnHMxUcKmFoSDFHkNeisI9Y7k5TfCV4Zav5DYW2ZsPpQKYFZrl50l
brvzllhEK2l62wj3xKwoV16R0/0fyvJFwEuvARmKBBhiUx90wxeOD90l2+gf4B0NW8hpxcdmzbFo
RqQ1h4ONbHOz9ao1ieO6WXLJb7/TKBiRAy9EXtS3heRum2nW/B7ZF2+DbV5ZW4tBfGz4FkVxKyCu
0JU0k+KE/MNEma9FoY/WZ7ITNHWyHqN0RLRmeTZXXbilM99I08/7dyOG79wL2hd6I2Ca2K/ALhkj
3m3OhmJ87qlylcc3xEkory7/KvT5zMYOJj+Rmgn7WfgTfucaMwjObmqPAdVTq3mrYdVDS7OeL2fz
u+ReDcezAxig5lFj4Gz8gNoJIRqPKu7Wa7MGP3+Vxj9unQzH7Ge8M4eBDY0+qb8olFhozOStODS5
TbMGgf8cHnOTJle47ZxDEZu9QixWgtNSRzTMj0LoaRP+PkCNYGGKjNOuXRDjy9Ac51p3GAFF+EbY
0A1knDwIT0Nhev90xWtmoQjP037ReOT5nl3TVZvoJifI8UDfpfHcgKcqvWFdwHcGElgoBk1kadTq
2eFHwMTQajsU13WxpY5+s5bww1miSTr47S3/H2N9hdmsYpT8bPIb8iEGkfUhQi5BUrtdfqo+qCNZ
nWHOYzrSAO3giXiJCg7d2rdV3T4yIhCw3P9///NETNU6HrLfSADhPxvgQGU7egOWn0it+PDV0orN
uH3Eul7TKgAGlfwgN1C0ug0L45nyFJNXwzSsTcYND9NkDw2wfZIKldAX+chGJeaEuBVKoTsBoScD
ko47BSDyldDGbNTSi/1r/tpKxJSOKBq5P1uECi/eVfjxz5oxx5ceYxwkmIMA/m6cDGnr5jOZv2mv
P1ZRfXU4ytjJK5BwJHAU6EEd/ICuUaQWFK71pqeH1xGVhjH5Rq3FiDN0L5FFsMtYpN8vVg+pF4tG
vPs1epdbs16eoV//WZYJWUsuh0xBI4ziZHd7DQvxj3/0xz3m6/GNeMf1z+X8ESu8zDFK0eoSLZzD
wUZQ4rVzfAp1sKFpqj8wCnGAbs9SY2sKVTSL8LgFLDD2t/4hZeym73odxXHpFHzphDAm1IraOlxf
MDl/+5sgLoANJWn6OhCzi4oPU3nGqsjZiYoDWdThWOI2TadOE/90ZEFRkrtq38v1pn4SzIl8tXPe
rnAxO1/YghLVoS87BdyQ6R1Kyil/hwCKfUj/vcmbZ6uUENNRwydxzpEzn+qIjiEVH6t6DO3n5Oi+
meQyr5l8KDvU6+i2L1aEve766KI+jBhn1G5w09ZbWHsVhi+ztgPfnIa2mMSVbOwzcBkZYGOzfzMA
+RFkLVw/6n3OpmEhULz0PavDhUP7TpMXn8vgShk7Z7N9vFe921DKW21TQt24OZJaVP7j2dSniZct
6MOWsyUYIKa28alTLxKE0XuVsdKZgJHT82f3c8MJo8AlGWWnZc0I5uA4Xe8OgiNy2HovUlEa/rQ/
S0G+bYEu6No6tmcCE0sJgvsoLKcmbPAWZV1zw0JxkUND+AGmHYH/8uyeKsO++loGsWl70VyC/lM+
b3G4CZxQt8LiOU4MhjzWqL00/Q6IQRsmkmNZZJaiiZDizWtPz5jvrUOV0SHL6glE5lQce4I9z/cK
ygNVQ9LFy1l3W2Gib5iODRSv17gyM/Zzb6uubvI/sFzr2bK06KPbsAn9kfUlP/pjWX0pLo7iuksa
NVwLve1SvnyOSrvp0wq0+C2+fhAvwfqdNT6c6EFAP1WW8yI8JPza7yN9xAp/Ruvo+4TpZPgCz9I9
l/zifP3wkxRHKNZz6WeaWxGjLNayIkn04azmghbAu0/Ctkwn6qL68dJYJCSh6S20OsmYitAmtVTk
Y3HApfY2SCI8akOas2EA4f3z8bCdbbJ/n8us7dETTM0piWz1gWWNS+ZZhgTX9rAaz8XZBEKgzh6S
Nz3wLEhkmL2qNrtjt0E9F8CRyLrSP4L56TBF0UiIxmCDYodZkyZFODesojLbapKzee7BgBylBHtG
hF7Np1Hidx473QsiD4Z0cr0YYyYr7ZC59/N3qvJ+Sx7fNWdmXlzZER12vunHMy/jEagA6unU9dld
pRDIeZ6aSaCAh7un+u8aCEyTr/1sRLefknfGw1wyVXLUg7KLxkNaMfWnIUDiZ9ovjudm0iv7GHtr
IU8vAZmoGWyH4KG6cjmI6YBARBoMjYfQcolzLkocDPAWzNts7VNQSYUvZNSm4NUk63pA0eD34LEw
TolJThidOp12SWbvzV8t4MTtlJ6bMajy+RjVZg2agA0pngcwHScyzBGLf7G2NdRIqvY3pZ8ywUUh
V897f8UdFcaAhdjhGIAVGnxZen2AVc8XNgh3y6dC89YVvm7xzQXdCiVc0LfjCfIvT76txtKcd6zO
RgtgEcDd03aL5e+WsI/3mfrwaz2juIUWuiWpSMsOAdEXIa1FgI+7X6Yc+8Fq/ly4XG6uZ7xByWSV
cSrwcFTJ6K5X0Be91okDl0Ag0Iwaf63o8fqpmbQ4xEfouRKuzss5mXboXtJk/hQjre4uoQfvkdzP
8pRxOr34f+CLctkj7jN7fiVCyLf49OW4hYmxiC2gIhnq1WrWRfj4Wc2w+aHO2xn7EM9Lmc+n8jl6
GqQjzdTSYmiN5rRGvZsrNwwQN+6eFqFaPvB48W7/x/BOTx/MX2hNkVCEfVrLotIlhAuhApC5n3zI
1T5muX5u4D4wusPJLeY27ZmH0rSnTYlHMEatiWrHrRsFtkb56HAs/pWzQ/UBhNxj6czAxmkLh9OQ
yzBxryPb6CoXGXTmH/2eQmJKCRqxQYme/c+bui69r4q7LXneEQIeaTFYthFqVkxtZJsY1/NT7eFc
XYU361xJ31B0FzzUHMHcro+t/FxZir68skwI7dARdOHzh5gPcYbcS6ojXxpa0U9wrZ41sf36f0qt
NOLu7A4PufAXjxojkH9QbYpa6pKeVE9Id/wZr8TUAORLYN7LtWrjm2IMOnQiKr8yHt0gTqIzaOkG
cT2a2p2HT+ho0srBZv6XIQM/qrYhu1sbrQYQGhtKYwV5mv20TCHNZpH1Qz4UJxYeFX+WSY3s5LCz
/mjdQWdxNVZB/wHJl2ahJ9K7QPb6XHg63yBVkgOlrffOqJxwFPt4S/8OtwKua2ld5PRz7pLmp1je
+A2YpyimjZCvXrmIdXjEj9+dEpaxMBiG6kjYvI0oLLopruTDF8zx5+ZPykoDDt/k2yXAvaeD4dDi
QbZeKxNZh6FZzXdXJBVOycMdx6UsgCH7mfv7qyFqrYdyuSeNcr2/goeFbYvvtZZldvyhHmlMYaMi
4OxmlL+SoQqLdQ1WUl+C3m+1oHpTMPUFOocKK/emaRKE+8Bq9m0+oUw2HHpZJ9Fl8pGOzVGxKu3Z
xzgDnjsRoPHNkEd8NDeG6mHIlrsp3g+m8zqDkHXhyAu6tcihVAJ3dbzzOtZSYItKy5rGbiHhFFj6
3p9//Bi+spJLHDRS2M63N63fKTcAnb4bXnv0xWf6crjJNmPw3e8drTIYMf0zbYUt9jnPQK6vv0Q+
PMflzYi3NetnZI0evRs8wTL8Fn0GkdnohXhOS2gTyvuunFV3tOPH5ZHaptQ6qEMsI5Mki1U1lR6s
dMfMOowPFcYPrQqTSd/big3lBpQSAoxtAahR1gBQ+VJm3OEoXqQvFLGDdYgbGJ798CCNCkDxVJ9a
OtjPQbYxMrQOc6/f2LJeUMkQDSXM5R0wmJOBtiZfoFx8XyUSGL2JUtqEgaBCCAE54g9vmQrCIjIM
I9ri0mBGNCLnkhrvuZSH9EH4LVCFCSXrqGMrs1PEb06Dj3bxNH0P79dbayvb6WSskFbCzM3KwlxW
1UpJobJWtEwKDqS7Dln8ev108S+qdnM2c9aEHx+LTTuVVW03dDOwxTolUcRlvTclCA0AhIGm0ufd
AV8SVnnt15UU6PcdnsjNcHvEyJsoSVD4UN7HkwU5Id4HkW96l1GHNZJhneONaAJ3xJChUFSFQiSL
Buf1/1VOWig3zctmGLD5iLAHV0bTwlrDkzyBKwyOt71yX2xx00XXtpdp/2GDhyBsXQSc+IHDN5ob
wu9oDufaBVf7IUgxuPs0aNvksAE+BFlT6aB7N0EdqVGeIJegle/zoYnA1cVefc5EXkup8DFknYqH
qkqemIZ30PmFq+xadNQ35K2Zd7ARuqICmxaMFZj/PkUPAyEpOm+HRm49vxlX2KBBKrdiR3fanb+D
lX22pVsKTMI1LYozTlorgxgb33IKmMMWrHjGWDNSRK3olY2XT2+hb2G3QeIpKoZ1odkX53q4SC2D
oUWlg5RD5020A9V7n3pnTyyl3+Zaj7YeEo/zw7CffsMfaf1Ckd3FnxQ75cM0eXGda3dEb9pRRku7
0WpSvHvI/ixznNSAe8eAuEaC4ZbKSfA21OhZjT1/NPaDbgvlXNIu5e0tahAOWYQQwWsl8K5pd2qG
kQEjH/2O7wQyZ3fHteSoyw2XTL8piTjzmscbJeLZVsibemf17iqf130ug/PNbv/JwMYadPyzxXzg
sK/GpkehO2aGMph+e0Zm+uZPzoeVhE7Y8ApYviNWgstBYXQYvKGpLh3HTUAqfKt6O55msbXP2coc
3cO1g7FDwyv1sCxGhnoB5/uaV8hl1zCOZqx9Nhh7L2s+ORzVGfRDAqfD4HWV2+GLvKUBn0BU4KiG
iSy4iQqqronXDdRGO/V3K7rWjmowf9obrJJUBfHXMx2sWX4oaWuxcjq6W8iTdIOBcJZo9HdRu5Yv
5m8Dp4B/aFiE0sq3sswjuCjkD6IGyMNWFWLkEGYoriiEP/TlYDkuZGaIZJFOW2XWI5GjzT5yHucc
juAeSdXvVrQxi1NEXbKWWQZtqqiNBxjFbMsaQSzex0HOB/XoTBN/4/X5irzpLrI7p/XegcxpWM0h
1aiarFdkg6l61eyiisoFnyBzgK7rdWzBQrHVL0LQwfDRswQ4Iklm293k4qNB7iUXjoCZvT6VQuzH
ePB42HiNLh4/g4QtR1ANKcPjFMJfQobr4yU1I1kKbLT4WDtdryjUc+JxiS1ril6cInHwNanCstWb
OXQM9Tmbo+eHtCJ/74ceE1p9hBm1XZS/DU2EXYTYrZaB9LRjHv2L2/9SZP06ViWUs4TCUaykmNGs
4D5+XOfat8t8igiM/iexV4v0wI9strRoInyil/CczjAFbhOPQR5BseosFZ7OcDlrasQ+T7h6cH0K
oXhfoTGW/tP+L4fxqk+7PTccuXXYkrnmQ9BnfqK5NQ3yEDCYvCHzn2Nri78ivQihO1Mc9EhjVpoJ
DtKM04iXWy9rQVTm3VxInF0nUagvCacUF+yTk5MAz4g9vU9vl4n7ZeXp2Uv1fdJSrMgB8wDWoFZ1
91jvx8Cjuy2hQq/dCskfc/wt41GNGbbIe7ImcPjbPmciMn5W5F5pH2X6MTgcfUas+rixbyVJfGeg
0aMKIIW3AEec2s2OfwxkwF8wi/JQjANyqvQKr29C5lPURNWURAqT4UO2mC3PnKCigJdoDtZfL0dS
lwTIm6kIXmH7hl22Z141rlqVIelCIgpxwbkl5gBd5RpHVVdJzu6uMAHHL7WQErQ5OOrqaUDF9Bsl
YaRIqw3b0bHql6X3AZsx/VQGEcWQsp4cKq0j+tgnm+plXLVbcmgPmvqf4HZVFjbPB+NwYxQU5Nwh
Y4puUJYE3jKar1/T657/omehhcl9bnMI8UYmLLK4OewHp98D0PKZ/LGBx9RCDZ8nnmDJX7kGMZI6
Lr2lcZHjPHhmMxnyhERwOXSurH2AifPc8t6sHAvhlQxLxU2oIyqxV/c9YGL/EDxbuiEzzVKzBPWG
d/genSY1lCUwUNvDBCgzUtYHBmhiHPDRoaeiOoWhJJQ6jezMVA0ER4VP0IQg9Ut4v0Mmmvf/2Oyw
dVTm6LfzhhB+BTIfh3tXqMKbz5hoHv4xk08ZRJD66h5DDEFE1O1m6dNsVRbKvZdRMQHjC7jSCU0c
6uCYDEVUE0NVFYCfSyoyeWvLs7es59P5VESYjCimS+iztCVU1otUdXce31GAksG0/bQ/Q85ZAJtN
nvQ9lnzaLYjUKwDRT9iI3rXsCM/NpdcvxhGSElMKA2K6836hf2RQutGII54MUFsKUqXKZrWJv4+5
L6i0ZIjTs9D/O9BEyDJ+x8pITEmEiOwwmkvxghN6gOTmvkffvN+meYyVkW6D3ZT6u7nsVCr8XBWt
IJpIckTJFnyCaid0W+jmxHlmgXyc/Hcr/3DDDBA+8egry4JGqwTnVbaRuh1o/s7a+BxvaxJgJEUG
BiTRdL4pQZqllRulH7u8rukMW13ht0/J5rHaWT3pEGyTizEvxwFol4YmRTO4y7lJ2od6TD32CDS+
j4YVeqOixsRXENG4HrLYIkHcQFV/Tfh4xnS9YNGnFeHQedsnT8dXDxNrtce90vEykQkIWwHVP9yt
RHyp83FPSYyLGiFw/yzLYW2LLKz44t53XzfwCVdlDVwwMIJ22EOx4qfpWLIUkeOZbQDkpOzmzhsC
kcPULIaq1InuirP7yIp5q0RAnFSAi0PyxEn3EccG/pgoj0JJsBwKX6DgcOFDFP8OhruBnOcUdtMK
Z6rc2XUN9NMaXVbXV+ueBMCq8YLP1XPPripz902HSLEOU3Qcizhu35o3rzST3+Dy8nrlkWJbfr2k
ZIHRCEtuJtqI91TgFFClrlHmGSdMAOfVMYkiD/8ZJfaJUaf7+DFyWcgU/AdgYjG5oxKHLggtxyIu
AXB5Pd7ORpt3tnwP5Hqfgr+2TjRz0Nl95k/avbGToPWsddcAAiD/ofj2qnYkvcQFTbpB9NGXJbPl
w9eZ5S3s5qfcOhgRTPsVgm52TgEYwPASHO27lucFmAsTgcjI1+ah5qWE85iQx9EkXqos8FMUSOpk
tWWRtxuR1jOvkki6mmL5xxHWjKxyertshChPwFVDXvN6Tk0f3rZZlu59JksM3rZijfGc8NPXY7fF
jeok3tLOhgnha9ClcNLansh1cEbxDcsVHbD2Vmb5SG7/s60VfSLe681FvQO+WZIO0aXowHYmq8ai
C4XraM/0zb9uSBa7dVDTi86B7I9Xf5KWVEzQxqWcu2N8oKl6pRbQCWWzCz4BWpqIKUGzxptob8jC
Mc2SlRkegQ87hagsGA+PYNB5kEYL+W0tnZ4mf/OA6CuBKCfjBRpRGewdFoWZse5v/zsr+L5O4agH
INfRMA9zY8HlFex9l9yHhBDxfD9g//TTRmzLOjORkvRpwVmuA9sRkWlg2EuVlvb8q6B5ezJB69pl
3eJbfsDW9nFH8BxxuiNr2BOoxippcd0+WVaqjy2yJfdVC16jqQ0SpUrj4i54wC++hD57jY98gEiB
DEVUpj+dZ3l8C4ETjOOQwLDPK4tNzyoTIVTHQ8KXM/gT4eXwHWi6V+I3h/5d0nJXmtcsNd6dDm7f
vTVytXrv4g4VXEYJkZLUnre+xw8jQmcKNEVMeypqlXqN49Ki3RVJmRTo7dtGikbEhf7YXyXgEOtT
QeBV6PJsk3ZIe8kJ+6MGsBddVpf+rpH6F2VgoWi9qF6Fogt5uvU5dqFu0hJ/CXTrwnoIKSYfBsfF
hi0xPg4MJMh1b4NmbBQshE5Qx/MOLo6aR+mxaEv7jg7DZEw8qw1kS3PZrxggxzmUbAiy4qKkBkmG
9CFURDTFeRbiaMdRsM/YydmZHKiyyM9q5vtcdh5jY7rFzNX4M2R3OVHhpxyQq5EnJZTd4QuXfWmj
lOzKTGxwJ2wYl6VpzkaM0ag8nWx7oTUvR+yp5cSaubeOU2F/+0EUnEbB8cw+EBr83zKWla8hecif
k1Vom/ufOAUYZt/NQoblJr2sms/WUbbo0kPVdB828iZNF/hTZuRc7YOUHDVGsSPfw0qAAbu5ZqEK
jgaA3hy7dYcYaT9UiTh2YltRNu5vIFjyMJWhZOXoJxI9SMfzDgZHaJGsI9eqgHKe3d7B/+gvjFP3
BA/EK+wi0Lxjayrdv3elEEQlV6SdsnKucnio22h6AOWZG6HOEsfspuGzigCFBvUuO7MMs2WnKjYC
ac7LkSh87bnDgmP3nm/PtSQHCjBtciDXKXjiQh1aIZ07y2xyEGi6E5CfBKEcpW9urNg5dcSPGpFx
HmiYqMxCjGjgXkH/HiZN7OvUloiTZh4rLDRx19l6s+prWVy98HVhrq1C+pst7mcm5qsZP1//I+5O
ct92bTzuX1kfrDYW+hsMf6udpCDrUX4HpMPjEbpPmisiyVWr+BvMlzEF7EjFPnurOyEQsEIUBWL6
dt9Ld1B1b4bbXFtwGzwFZ//z95ZOnjPvBrNZwHHFirEkwwZ+R1ejbyNb/X8dTjJqtgAGQUxudxCY
5Ta2sWpJmZatvoh8ilRQ90yBaeK8C6NF6PnPPVNT1j5zstpaNb4qfgdho5DzhJfCJBFH905hpE+U
rqN0tNjXTvNrlJJE4zPFh58aZOXLXcUXWeY48GEK4zmy1V5FEWDgxmVuExVlyN9DWcZsyjoqqH2N
fM32wmTBIMa3TT/SgaXeablkowkQh7q8x98dtRLteybmTySKr4qHBSbShK/mTT0FkSwWwsohUQFe
IOxWvZQeeeIncFH1Pi7mP/cM4UEbWV5v2tTuJhDq169KXTG3rVJXv91yLj5IYGVwGDwiCRcIi+nJ
RgboGgZ5uPm/tdi5c5dn3ZtrpZaRtcFEJ3E/K/mwlASs8D1daFtKkl+D7r6mof5m1+1HttGJYPX5
gOMYjnBCwBonrmXaKzTMtoBr7mVJ19/KdkLtsgkge3UBstf9mprU7/O8ULpW1nbPTbg4QlXLCWYI
qOTC6V8X+ldtvKnIzSYE0kZiJ9l0dvCFo1YiifstSm/rbSwsYEV+qryBUvSp2qknDj0FS8hSWjqi
B3W6kmJh+dPlzsVnZw8eDvYNfa2KR/e7Ud6MoKuTCQ0w5TGlcFQWY4w+/NojUhkVPg9cWHmMFEaU
vNyREH/f57S+9/Bzmvrm+yU6vTBA+fL4x0S8iUgJ/+k/7yb7lQr27wA/+Rz09G/2H12+xAAED5GH
y3f56mS6euaEScZNZXetB4Kb+9RK7vxYsHSZPlHTqZuzWLdrgRO2Z9696KAEMo2NgGKvavM5TFpF
Uw6yTnX9rEqbGcnt8ObryrDcJXXJAyATLUXSuyMMnOiHgQKI/KJ6PeBY4pabN93TP6jQz7kLTCVJ
RfQt7BUbfGUvbzEvm2iXvFkA3PDW5XPDenERXjpoE/xn8Jtz+ChjSd5hzo97hZ+bqfuhlOva8vor
deyMTQcvRN0lK3G3x0sJq9rOss5VTVSZGB9L6saoV+yUuaPwV5Ac39qryx23fzFSqydnX4Rn6dd5
W16QMQucwpo7M5ee0UgJ+nZuaxXr4JlzBFAf7m5nRQGpBwCUJxdKlvn4Z1dbEIon4CC5MRFM6jHi
zCDHx0r9K2QP/JcW2EpxOjcEmm/5LUwVZgGiHT6AYML04nZMSZybNViClkMVn20FFW1e06ZpIdYE
jIIXxQ3O0kFipZTclYAYGd2DulEDzaJ3HJMuu+kMLG6cm8mTwWlJbb4+eE/hKYbIoPT3UZAnmZc4
O1iCwB+4UGwG+EwCFECzlYwLW1mK6Unl+z7DhguYKV2sHfmDL/QMpcmAhHAOwx1qOL3wHPn+Ump1
d1Ukocp8hyoCQigQJo/qAuCs1Ba1KdJgI7e+YXMRTd//fIO+GFrprD3nMCRWzrCYjmEP3CVCU4AA
Pjb9E5oj8Uvi1K1f8+E61pPdLOrnG6RIoSssc7RQlhA4MkTtP4+Ko2Fdcm+4MqZe1inhSQZOcdei
sxl3gaerWfYZRgsVLCr/qJfjQCwC+m/4xP4dtGkp4TR0rFGIx/RK5UoM/83ggT8dnnxMVnYWGe+D
fOQuVqMIwTRCauj7YGzR6uB8JQRUTJ5hI3QHsWuzXQKJOkWmnap4cxl21ITlst+kSg/wWl2ms40o
MWcKD+hs55eCZvwMC1Y5Wgml/hxg/C9/Gmk2lZfvooVsT4uPRvfSwgTeiRDoSAusdP3LEyggem2s
iu8npwM5fRt87WhsNtXbL3W7XzlHegS8q8nCGL6tlMGhqTRXuCZl7reWxLQiFM34bNG7UrxBdglZ
fEvd26tRaDyiVXLBmDMYhVd99SPA7Q3zVUgWAJXGb2RNTAkaJ5hiYUCFpm5/D93d7dB/WXTRji3D
3ljo2dvo3IvADzbv9Uiig/TFnP6iSNK1rsQLGkrnSURwMDAaavBNx91asbxvBt3lI/IprI4XsEhZ
QGe3+Qr8LxtdVXHiXGUjaJhgQuMBc2J74N1bheQTczDDWzG0QlsTo2Euvyg861s7xlMklPR+mL4s
il+5bkoqzxT34+EHiONmBDKFwEIwj7u1xK55+C0EdKe6okh+R80IiWYiB+j233bQsu4Ri2TO6Apl
TnH1qNrY6JleLY+i1as+O9Nckmk6tXhVZWML1fxSKWn3X5JkVAvc07jC5RZv20UAGVhJirlYPM9w
MEXLqnSYuQg/82hgSC1+ykYQcM3U8fHOQuGhFbcFdBtTi5R4UcUmLDxKC/wvkPCklv33NHr0kk+8
nU7W+mFJ9UQ0qlOuipgc5s5SDDyKQgJax6d9L9S6ocgOAcBZ0KnT4/A10oI1/fN53pC0vQbCJTGf
z7U9uJ2vp8puGb3tLwSM743O8YAIGefeezE4sn2hAN8k3StWZyQU+OT4aNHzNHMQb1adWCGeB6hk
l0ClKVH+Q9pigbloVcwmQpP+MP/kkWRZEUj26f7B508+POfPpGKZrh51KRu+PjbJIORVP5MjIi98
AgeoIiUMfXwg9h/5gpTpkJjoRGa5Z2YUAKAyer+fuh8+riT/R7jUobVkagDj7h1mZTytIpiwrUGG
p4JVzasM4ISSFAWVBT1WxNON4mUeuJfdv1QJDRfFKQZs1qIu6L3KbgtE2vrHH/GxjNOmpl/v+JD2
MifN2TfXyITiPLs8WoDjVjEkyInW0BqWn+m3ERqTzKGdR7YKoQPeEDvZNkEwDKj0OhsTwqm2oqAa
m5QMwunCpVo79j2NhgILECdAr2xHstYZlY4pSUSI6LlhF1tcs6aV+CVRZSX49N4PHp13tMWhKMkk
6wCgojLziIVth464bm5AP9pvbiVr5XqVAFftbXUfD/4/O97fj8tmpmXomR1shy2fyo6p9gYG9Qf1
wXqy0aYpLuyVzrbXGEWTlyiHzAz31LwqTimvwqbZPekwTIF7fIxo33xchSBR3LfkpwataUW8egFY
BDVxOeTQLYC1xJU8YHuepWEti1Y3PUWV5PyZiT7ILxN4kipn3VIAjn2asSQPJWJJewV3QfGsGFOj
h6OsNCC+R4DWSK00uGQiu3IEIFvTZvkYmf79FjcyZfiaGlS+VTRzHQumTAuLISAot2HXqdfk2tsr
242ifSQ042yr/jYvEb8Lk0GDl/6sN4ayqp3d9x6Q1Mh/evos0hwsiQU2WGtu2P0XvfqUZ/T57K5i
Z03dyA5ZiafKvRcj2q18CKMZlQf5+paX6i2l4dSwiZvYNfxD09q0BEnempOx4usEFeC1uv/7P+kZ
d+dH2MwbCxON918gJnYyeAc2cwLsv+RZ6YnzrrY36ivNNw+EXUx6YZaEmcv2wv9cEnuRf6VIqLlM
cF0/JrqRRgeV0EwmSj8VHG6RUJFGMfuQQp8/DdJzWFYmQf4SMBK5TmvoxpiVa8P2/OXBhsMIUK+V
MgWiw/LOwkMk9UnIbnEVyGvPCzDBg4GR9rjRxOzWbMsPqP9IYQ+AX00sC/9TiKr2y5ydm0o6b45o
EOHG5ZklAju9UCkvEWAl3EGcYKGyN3QfSIh6DYSWeYhHf4faW75ZZGrDP5CLx+lRGNgm1p1sq4jA
anaijPfH1U+UZm19UbyIiGyCnF9QBJYYAS7ZLVE8zX+n7iZOpgGT609VbVZ4Eqmrtw1ZPBFpvO47
MRpazew/l6JySNmV0dO8PEy2GM3qK7WZpgijJaM+3D95p13NPTclBDtEDheH9N6Powwd4pXPqam4
N5Uju7k1sdZoHkYBzLyyekegV9DSVPPvjN63Pvz8otyri2eTCMUHM8wBBNZWoc7gaTujcWyq2UOA
N55aM6V0c6G7lDme0VK5Ci/ZYlqUx4xtJHSuLbc8zJLsJ7XOS4GmX9fOhggEO/uINmEJW6AOGEIg
RW/z8Zwd3qLD9NeRgFJ21dWDMGVOyqIz/ZeT8ki6wuEHkq7JCMkc+KgZirIbxrXu5AGbx0NTlO8x
P/3AkhswFFqfxZVj6a6rNSAfITTgTOsqHN3HM70syELq4jY5GnFvbtueu1lzCyg9voXyaYEj6ZBo
9Q7vq99SUbrImQC8mpMEz8WnhYl1L/XxnvsBeWLgHGqhUVsyA/af9q0P8w3ponwzQsYOEVMfeBw/
ZY3IupUs1toSWJFX0A41bqCkO78GfnhWl7wGJGdlO29OPCRd+K8/shCiXAQlti9fMz7OCgxmOAcl
Atnpu9ZLKq8bbHLEDoa5hsjYDayDdtzg14AG5agefstcO1rrFdYQ9HqxTSLIVnKENLhHA7HGSiVQ
86UUHZVdnrpSqhGmXZRYPCMZUR1/WP1nFY7ksV6Lunl2ZBaD9RSHKglC0uKSYCfYnIbaAGX/qL5d
7TsLA3iqTpVwWT+BkSnHo06BjAgHw1IdK1nYElTJFk1C1qihP7O03WM48xgv/3E31GKYtvdgkJu6
HkoGPxZNsjIFsV94hKOfp1Pk2J+yVcnvAQDgFVgzsmtSgS7tnCp8hHX9C8klzewZivLuedWu6HJV
XvBJQ+d7hZM3ViZBtkoqfM1hIO3PYUDD5z3y0P/fw8tIa6dRH8WLBXaXiBxZUp9V7N2oL1yKZbFd
O0f4ASmS1ohLMZd0c0ba7DJjfL29U4/xPIhOCtfnK5uCIhHIRhAW2HZ3oeoqtIEMWM6RzQS2mY/6
OJOLKeUXwoqnuLisWNFbXQ45g/om/fng77gv76/rB7edi7LKm7CiR5pb5i0PdZHpjScYUxOW9ISW
h05l7OYq3n1FbCrIVyFa+nnpmiNOiTxssdnIhNlQP+dZM35HwWkCVLrxQDg+QWefFIRoKrAPJGEe
OFo2rv1kTVgnftsfenY4B50PldXeem/j0AA/8ntDU0Odq2KTAbiy61ezcvMKJnreA0Z8yhAZ8ByZ
hg/5oLnGKWBWaeIPIQzMZLl1RW2lkZhTnT0e/3mCYpT1ROYJ9/eyBYGk+kDpVOPBvu9L9gBrrGQg
m4gNZP9dtMrn1LZWirzx1/PVBWGnkWGNp8MN4eixVgmrAT9x1kDp9TFgE/e5EPJbtvlDeRH5ntel
47ZVFwyO5W47tjUmsmiSNGPJyNoM/Aie8nx6oHiZHiEZ8wKt1KMJ8GGccxKt63rRqerUcbnsilXZ
5Nx2ew9yGWfSXb3Xet3PXfDnh9ZTHb+pNILIg4ALsfpRbJ3G9Vj3p4PFoT1DR6U8vxDOB8pBNDJe
4dcPgoPNGsqKY5Yjk0ztsOLejtIUGHTjgTqLumj7AafroQPhKNzQRA0rMuqnTjQnieQOYv+6mwW4
IobbfpbMv3s2gVaVSv6PIdsfRrOOl4qrYCSapSj6Katgm4iBesdyFwVv28XsFJFZTBdRH0y3u32e
TT9uv2Bvb9Fsmi/HDFbQFjhZRbV0Kdk3CCpGLgSRnHkokE24rtbn1i1cZBMwF6aSocux0UQFqJF2
3NfoBWY0ZnHwN+H1DjZezVpLO7bJRqs0iuBYG5OqIRE1NMaZBkO7Jti4kOsoKCDiqyks43o5/ADR
TrvPqgOCv0jkfkM7f2zPVNXqL7e+7B1fkxkXEpAS+92nKzA/7zLWY0dZAdAt1/oGMGjKVGvR7FWX
Wp/gmq4YyYbRnbqNmc9bZpMWsj6FryFQYRlS0XlNvAjf3C3G/UEEu4PnUQyhpzwIkYsceeH1ZQLV
9N//1RWVlKpxLXn1WPc5h+xEa+QWQ6PTsEPY+xymNzxRwBa7cVUbyCVQLzDRfTUGEyEzIpNsjDDV
mrYGOnBqjHscoqlla7xEp8qtS/WLPoa2B2VZ0wB4L3rJjAvQ125m4U9S8vMklrqOSPDPwYtYYodR
daCeKeUxC+NK85C3XuMU6ly+ZMHnYXJdOEL5642Y5vtyPLjOklR6QyBBAJkPJ48VYCbAUseWeEkw
Ju+alWAnh2+N2GagB+oFjQouM5OsMJi07n7CVrzIlkE4M2vspUsguy+1ETB5EgFnBfKibE53m5xz
wEPxzPBhBdsmQlq/BFz2B3/DyQH0MtZmTxgVaSPaDfwjqpBTd6VInAGyazAzGEqe+g/6KIBfNsPJ
/etIaCLjL6ML+4RJEKpPuEGk9eNjcKM4x17+Z3lN48yykhsaUBIV4sglrCLlmPAsCHV3H0r/A/tE
Hz8qCPe2uvYD6kwmZut7j8VBgjPlRMoIG8HzM8MThtWkPOpI3o/MmNJJRut1FcnAerGtpCxT0XBy
Z4BCZmFwXhYZrnC/h8mr9bXVb3STskgVJbRXvAyJ+upubCB9gSkkrOk/Ws4sJ3Tw6yEtgB0qyJNm
1eYhJncNM4N8G7wD6rU6CXIOgkI7/jY1P3K/zAB1Zq3KZBj7uvxKEcEVKz0eQmXxRsjP/1LXdeuC
rIPkfO37J8nOT4WleJ6JR65lTFlU4uNZbQ0D/Ixicy2t8jE5wWLC1BJVclSRYtDra54+Fv8HDiEX
wqX6/9Gwz8N2kgnyXaBO0ujT2V1dNMtj9ComRJoT8KX3b7Tyu5vnAfmhrXqYmBBDn03mRe3HO5dI
UyukYJWXOFWPx/yzQmt96jXvy1b2AeQySlBX3WIG9gHyHDxASz85seAHfO7HD+ImCeClepOWJ+vv
tvUsozWc89Gfv1sFC8fuXFdwov3xrm6upqzoiCKhZbOOG+8laHkukQQ5InPSn2cQqjgjg4zyxJbU
zXMR9sVr6TAH4V9X9kIIVZy1W/IUyAC+/4oIK59tEHMOMf9Py1DaRNPEu2d5v4y3i4MYpux4dDUG
XqXL5EfcanTsCi4bWC2KYcdKIe3RZNtVa8E3f24aXLqaMWnele5JcVsCTYWAlSeYpR7DgOX+Q9rr
s7Rg2N865rNuzNY1xnH7tEHvcScmO6ZR6uiWXIaPvBwr2SZZ59WDj9JLmoZnEdE0chyZ20o+Oifz
dVR8IUKSQ0T2u8Yp1QrPt9vwBtfja7coH1isqD59AXhRADXwP5ikgN3BvFPcGe5yzJkROfK/6s/O
hDeou3w5PFY+NmfinqwHs13SnzEST40dtS3I5SCL/FxYMRhu4qGvaSMzrMq8BzzqJkrwYe91nY7d
kzQ8vxCj/jwd7TO0tisWcmzpxtyzBhSWaEWPfzCq21NG5OE7rkYAancJf/DEMlB4HN68PqPt77ry
InqbRPNRRrWLUsAMtNukZSwcFRj0mPjE9skTTBNeDUeIJHWhr22MWhmdzYPehUCoXQHJmvOz0m+r
2ThR6waTI7qYpXVf0SQNL2zXEW9Afxl8oozno3CuHsE/Tq1bDPKF27ZYDjozquU57uhCMWOI9uPD
YI7DGSvCDfxPaPHKbjXuTVfqx4iO8VtL9doyz+I0v4/g1ziMZjE4ZI7EI0cnw+XLqe3diHVmBd8a
+QFZMSFBMBmZqJe3AMtWsoBcIBH4n3xkakMlbtxUaeo5UEIV5vj4tnnt/j8k6dD2hArUc5LsFmc/
RhUofXWpzzWE+MpG6WxG8RUz4bJVX0tFQYEaTIPAgA8FhQru3DxqQWOwJgt+bhyWbrXrfjIyWa8c
zE5Ss6vU0HHOEv700CrZGGmYQ382zsqb8v1kOsn+ADaELBDUhqlo5HGGNHvsmaKBjL7fKk+BQMDC
bNi1vmsvOtoN+tzo4/O85ba8ktzfCVP9REwBNyft4Gd42L0MRKSdHNFIBMdLetbaBgz6rt5W6TTC
PLKRNRB0lWjc96DT3hB4PT238tepWoY4TxWQRHH6qxYQhqXODAI4VxEUndEArgNdm2vNcEKQ3hTc
xL5qm7UJ3Kuo5oDWD6h8huk+c8uCV/G6tKkmP0+9kxNBcaQau/fPiGFBJSI9XezHbytjgv6ErRSs
uai/tfxvZ4heSI2bnqB8CM0TZqZgh6tvFbe975tWjV01gDqclzCgg5nQ/Hn37VBjOXSmQFoghcr4
o0oafm0qxuMWlS6ePv997GgCKy5/gFPCpSGLlN+n7KkKqSlZYDKV0mrDkNBKXUPnLiry58C2GZx3
XOT7w4QA5FDz+vNax4Ih6ODQoc1CoSXAS9DOxzBKnXfx6qrSZqu9q5DziQCV+FEEpIpA+FfsYrS3
exc1nMybytS5tW63uV1eOBEOr5bZXy+4MEkFO6Jt/CJdJyle56dL7Ett2OHy6USMp36R3KYkCQft
OyECmArNAtHKATEYcCCvdVDbOcC5LLONRw16+ys3MVVhLhqo2hO+/woSQH8nWO69KzrznEhXfS+B
u4GvS6bjtp+7G2cgNlcduQ66HukBfxambCT80xr89VQ8gt6tSY6Y5yb6ji75fCBDnoO+m9jXE8zo
wjf++vxm4fR04I3X21TcoVUteRubVti1Y8osEaUCw6LRoMLPYLOdLkFXKVw132sQ3uFKq5NkSgnH
w8kZapOz6MiUFeU3eEm3XHV4pDaxvhbpLLOlAG0MQhCHQZ/N5Q1YGJJ0ykJZ2oc5tyJE9KUzCERk
EhlvrsNhV1oUK1MqMrgoGr+No4CSBuVVVHaLpJuAb6/Dx2JdXpFEBBqRGrxX3Z5MHGyhQhSvYS5Y
RWm2RgUQoQkBXoXRRYhBKsVJVwwoHXlG+8UUcu5zjO//ZeSHKeSzGjcKndSxmdFzL/Eh4oU8v6U/
o6N/qP/hmH1QQ/Xl4QTQLFECPgsRjsT7K2cJT/5JdCKdIRkzmZdLUgsuCxx9V+jsYoGoXgdSfBq9
7UEOtU839Yf/aw5Q+zYudpzkmQYLndiS1GG4mXUT3u+j5JqxQ3eXlkQge5geldnLLb8DBcgfHAnP
tJmoImAXTl6vHGONetZZZhBmox+3d2rrKETk5ob3ZinRVQ1EwlTqbSopRIQpaNkuXTJYGgzNfgWD
+40qb9LkDLzH5kc/bRaXsT81M+v6bZHI/7UlmXsZ16QWKINa9YEWYxAnr6H/hDYzvco3fA6sdYoV
tkWGQhjSQZNUlDr7xcv4FJZRhDqAAeCaf3aE0dP4+Lj/TfhXWMXnDIXPvP5GlOG3ZNJUYYPtReUo
5PsIrz2SaCzf0WaZWc944dXFvJrzOSM507C/ALm8f85kl3CX1lH3UdQrBrqP077UWga1tzb0C+EH
PncpApXCQBC87H8l8CQAkQFQPftKDbzWDi8cCDwRTwsqeSZA+MYAN2jo/G8bDkmy4r5+3TrVGYx9
kJ12b1nZ0xCd4Ecq6fwNpjhmXOmv8F1Y94aqrdyQWiNtJgui49SQMRrLoxIsgkHeer7juW+Rt0HA
ZwFC7Ni7qeUPulabnjlah2Qq3HrJ4XXFKF5Ih19Td0C5tvXMnMRD5rzcvmfWXwviHQgGlKHbyPSm
8nPIrefFA34z3JMY8/0N8rpQ4Mou7KAbnAu385j3nJ4jWgQ4NRhUtwpRH3CLH0AFzAIae18okL68
8xBI6wzFLBSXY4Z/KPWyyf8WGHfY3e4vK+hqozBpvp8QFMPhHLCgqWkwqY1Pmt70ILG3NdQEkeAN
Yf7UEgRZFysbI30j/BvLNbIHLVpXJu7E/YbsQF+nTxdRT5a4Pwm7gEuWGKUz2XWi05+S8xE3+583
91NiL6VKs0JAU1Zmx5m/yx9fjiFpdWSKo3Lk1YDGTK6LOOuHlL7bW22lWJILIUQTuI8DOg7co8lw
3nUOdjOB1/1tyUh2v3r9YpW6alVBoHIQ374aMVUrBmaAqnorsLUt9f8ox83mCtw9bw32eOV++U+H
M5bPU4wcyZfJB8uGhqd+4x/g2Uhuvah7uBwoJq1jqLqzHUEFL1Sx3HdDpQ71sUiJLp6cOuuAHdYC
0O2i8SbPjCo/tdmSqmLagYYwMFI2EbxAbTshzztUafEIFljUc696nLnX5RCadmWdim7voINqh70T
PmgblpTyP2fWhUh8REUqZiy1ciYPmaXxMzRT/OmYMFu6yaOQuFUsDWt5/DzHgMSl9L4fceiYzHdn
YTkK4aB+lanWiKN+k6oLeeOpWPuUW9VNjTFRzDO6mW9jYlAqqrqxnznCIntKtRQYkIRd9c7siP3n
z+cDEo1ESKCq1gkS70hPVIatzx+k26OXMLQgabpfSR/ieC68Gln24WU9WOTS7DtlgLxxr8PF0LLU
BtqVF4XJMXvTQCZRr/s+EwayuIWGh8DeOqzTMhdXpkqAw3E6IUJYrjsKbDgiHnj5OhRg28AFuHMJ
f80tp+Ut6ykLFUyvapiBTa97qSYXY0CJ/H1vifrzk+Kzbyi3P0tJfceB31v86RnI2xN6QFdYf49Y
kYshty2O3Bv02U85shwaBmwYIyN5b5LpmWM0P5I1SfsjJFoT/B1Jx5/Pg0npWGSN904ma2x3MX9D
nheN9On7vdc2XAPBUbL2rj0O/z9CwIjlU32CixrInicFwiXJ+oJXg36q8jOCvOtzQye0tVp8hh/G
d7JinMW8SQLzO32cpj4bIKwxDbfrKLo/AeDJ3tFz3E5xNORoZ0DindfAZqGWX2myDIiOVSV/5MMu
tAaan9abuBQxGlGCT3oegma+xs7tw6tWvNnZqaR5rJF1MsGe8hYD5l5sVhq5RKF/eQ2veZotvAAg
tzev6FTh08iFUYbgx+dXR6RCEGfao4qQ4wlEDY5OH9TqExM/GBgehJ9FpGDWi89CJw9yLDSgeXHs
CaEjZhskidgGY8b0MTnRoIXuIJiEFZulDnevYIUZMQA3GZNW4pVeyfDFYD2ZRnTWgk4ZaszsGIAi
O4DLguBpEfJL8whdI32ERFBTNGdRwDB/bjDOW35lpT5g45I9peGGfhspqcPQ4AzDxRl//YWLzz5w
jd8Wv4PI7sSMpGO8El7ISeMCAV8dPhrlDgLK2jfTTdzKYAeUJgGC/9AVGWZmEUiWpE2P5N1uEe/5
jwb+YcprOJ/UpmW79K0sQexCyUbU2Sey1J3RbLGPzY9DMMcw1KK5oU9dVDHvuAeZZ5YKGed6DwuN
iusicHriMWYSBugeeaQDziX/Vje0d9hJ2T+eDwI1qwKWOZaFQ7FAcRG+NoLAxw/kDOykjfn44QGt
kseIbd71r+OuhhHPta7TBkqWtnnfq4EhqDK8HtEpMYTfix3LHeywruDHpzuHnl2xSYKrkm2sbbMc
4mNVxjv+QpJ5vwmFpHmisN1cxvf7K7PgmIccvW+Q/ck8d45ybBzE7gPe7F8faB/+XYJqSiyXp+SQ
LCc0A85Y1pUo4eM2x/JE9HmO5EkNTqrL1e+SEjnXE+6FhUBDt7esZBsMXPVgFOJlbkzQ1tGy7ZWx
JvYt2F1IFuqMcTNRXlHOlzuqNJcujwPzCLHfnWma/S04YIeWfXnLPGn1WxdT8MzW7kiPA/wUudya
tZU5M0zaDx62QkMi1yR81h+aoa7R6M4GUKBVBUDp5G5PoCHyt18SLEg0gZvnfTGTCP1WuUseoPEK
cX4BJKCIilSapeXRQx9fJseWyiyvIzRRjVuY3bYP7i5AQwwa1tKXZa+mVWfEkx3PJ2pCC9MVolXI
FUDAMv96PQNvUZh7C74OWZxDemi7/9DLbKdmuE+j9BvQvsA/qL6R9HKckEkR3Ki8YmUdG0mKVUPN
lI4lR5RzSkl5ZVmKA3NKb/qVSjvZDBnq3gCg1dHj42R6RoJvaU+os/CWj3hiRQeur79OQf77MX8u
FNrtDoiGKmLsOd1Sg4WPWfXI8w9djuvwkKZwtgAitk7rZkZkF0vxX1YisXqd8Jk+J5W8tOzxtSxL
1BB0VtujTKYvCaP/p1+Wx6G6GbcoKvUrcFi2SpBd4a1Db6BbR2m+4MzCdpaW35eX5BOL3Q57F4j0
Ld0CuBaYAsw0eBnc69hBtjS95QpNJ4Z2GsbJ5Mw/SnCCgrhKao730qMQ5Jq6d1bipShsATZ1jS2B
q+bdOm1QQAsRaNq5i/zLCodCyLK9IVEwDDdBbWICf+erWRBwLZcF9mQiaojJOO3FKj3dC310yxl2
7zvidMWndpsIqq4Tpc1mDM/hsK7EkyyPMY3De6LnAKPiRQkuJr1NAJXsdwpm6pWyz+4nknJXJepA
VniUpnNqZ3yg0JXa94W1Q4KUnlD4rpn19u0IEQCBkQE4hlXdmvx4m3YRNX61FF+dli22WToH+QtM
5SuYPXSq8FGpm5JsvzAFxMVQ2kBzC+gfRvH1FuBAO73BOJlR8F8h8kC3yABnVPsTzjjShek3x4gF
/zGtKJpAQe6WqcAU/U7FV7naYq7jdMCr3eRsGXtcxPcKHl6zC0SrWRiywMVjqFgDTJVP0FTvxSwI
t2WmL2wY9MRhQzz007VDYpSY2J1ZxhunpJWoRoRJYYLBKe9ErPJnMPqOLZaBDbNacIAVjcimQ7Cr
P5NSsw3bCKbQ00OwrL1fI0B4+6/ERRx/LlW0z1XSJxIaD2Ts+dVmAkH/DArBmCu3oU52KP/xvGTU
622Pbx+yykJ3ROQaPKbGV7ZXKVPfp4Eki15DyZv+SADb9V6leQ80zo4aF7ioNHjhO5IRjllH2ToN
uBWrOQrhmfFYEF2epZwfK5T/K34rQAJpz4NwcPYjDVyXc3rWiWU2o+Hlqwk0m3MIx95KyOR3TlUH
J76f4J0k2X38xJouP8PL10NZm3JRMR28k4rDrSCX149DiPkdIzEObtMYyheFQPCPut7rGqAcycxW
AdCftYZQmr9+3XDyBwiiYT/k5f+WTejZ4GFGpd8HwkwUWxbbliodaV2Gu/Y4hlo6d3udTD+Dt2Qu
bqfBKb4DZsuTkU2n+axNNsf4p6Wy3017VALSuczOqECafdRGYQW12DGNb6TwgRe/BLQRLlCUXj5g
oSxh75EPZP4qMEKrdRavN79cA8NpJqEiyh6sojjalBwJ2dMRvtNx7n309f8aLz/tG6FFxvYvdm6y
6/kuiCvuVbvcc2EdjfuHzD4LIDhI01syhXB3AKNLv0jJrsyLmwK2O3nR3w1tmgC9C4QQ9hNGZxKz
i8dC8K1f9e8oVFWJ/k9FLOOwF3u2jNscMgDFO1YoCPQckurpVE0jD/IpwUcEhn72yecse/pCRw8u
wMN/aRoCHNpFwVxjwtkhfn/f4Vw8y7h+0nfJtXSnK3RpFrh1GioL+s8Qix8fG3QQdJ5kgPhz2uDZ
/4JXPFhmE+1y42fUzzb11HQpJDqu8AoLLdZHEPJV74dnvK+ZmoxrDEc4cBVyCCASH47BvKiD/wTp
F3y/jAsiGI6aemKTbnKXjDKrNvvYwTj9hoKAWWbG2mYNaacrIEnEQsgJRBs15P2646m9r+xq6Kv+
xwSZ2mQQ0s0bG+xur7U7Wf+iqcEhA80CzsFwC2K35qkIhHy0qCI2S8VUddXhQl0C+J4Q3X0ieblS
etbRCtoM37HbiH75dZdf4fmkOx/UA9xMRbElGNIetBqmAw16Kmw/OqRgIRq+OI3j/iClvBzOD+OW
BSA6LgQAt8JvrEaxgsevD6r3MjuMY0e4VsOnjI68CybRonG7n2b8VENaAtfw45VJ9Fc1t53TYGC4
H8iuaCSUjSa5d0KqP6pcVi0hxGZIl1LNed3+VG4UdVleQkLXNohtcsosvg1iXJH0NfJ6CKRA9owr
hLZckjro/6Aacjdwn36rttOdXh3E/ETvGmjkMo+UkPEuQnnmz5+LjqAr/pJ6QtlVGnby9jiEor+L
72SJcVesv99fv7ZJt87X9xXfqT/lboAazGxumlLZHhZ63xRX/V2PQ5JWNEJfl2bKPsZUUOBMyZvx
2qDcDAi4unswq96FQNlfaTBUnOF7m5Xfn0yxP5l07vXGWvonaGNbaXbPu5aK0idK7/35oqhB2QM/
X1Ut6kpqD2DohD+mtWQajDvmXn1oliYYqZRHtEtVboQchj0W1ZfCv90sFLsrUhv1Wat9fsjV2tH8
W/7d+ufW2Q0rDK03nRy1SPioDWQeLdwmnTsYUAA8sDViTQD30bR44xzkSyDbZGzRUP5D6tWg1/hu
pEIf9RkSq1g7oy1u/JUWBfAMK02QZv4YAHNrUzu++vCH3wKG6FPrg71rqgvYoj+x8I3CSl1NTB4N
3nBooeXmaGs69GHd53RsFprVj3n0af7X3zAJN04tf61tOPZTuPizy8P+zceRx3iHwQDVI96dThoD
xUPdv4g7OPvdMe2Gnxc5WRMmrRFhK73HPhgK8BBR6uba9D9/jw2TItWqUeSLmhNSUFz3gFm/IrTZ
XRMxyQIAumabJ60+pi4ofkL9jh5S3n+Iu5TZapE/f1LkXwfgRlmmu4gOHZsfNF1INWn8TzbQigtR
c34GfJnWWQgiZio0YWuQE23Ea7SkEj0kc2/kQ1slaV1JbFXoB1hTL4r3+oE6fC/RSy9eubMGEZBZ
mWiE4CFGNEt95UNTlITCsjU=
`pragma protect end_protected
