// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MSmSYvhgTlKUEcIZmeAU3JEafk8alvxz5gmXvDDRrV3PBSVxgTnbeFg0Yk5uV7rk
qomPs4VYCRQHBa+4fWjTozhOFrBeGi3pe6zpjQNfTPxqTDLE8jWR88GqtGQnO1TC
krkSNOS6m5NhOur4QQGd/QwX01O4nW1ObiOZTRGY9yU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7152)
PKyDAIb571YN+nQhIMggepLki+aXov9sNEeKEXD6D8xC/Bx5WRlMiz8enOcdrI83
ZjMZE+2UM4SgIZVecCNAlkrmdJ9Maw2xSinu3Muw7HK7aVskykGZUxVOHOYGUnzP
nw71wmLohln1c/uDu0css9JjicjKspR81+t0rGDVW9cmxGP6WuAjtAHoKiNwCtfZ
v+YgjoTCjJmj9PvmQD+kHQMMAD/o8af8eQzYlLyOCU78mAcRNE6dnl5/DvV75geB
vLKvn6wY+eksN7D/tnJtDL3mmNRGboaDVptOzlY88W4iu7iLg7FR0my2V38vSvv0
gW61BuM9HDT236Z1DU5ss7U7983Hl5mTMGbOXKGjsX/+QG8SaCq5cDBU8DZrqLlW
rG650eVyRhKDiWWQpU9xN1SdoVhnQMZ3walQD7hgf7u2dW1IRBbL0gWDizmp0fgV
XcpTlI5AwlL3I/tdaAgDC7D9umL+ohcC9CTaTpNLA91k8gP7VLOQPzdlRScSpHYt
jdKw1oM6rIgYwqd+f42woqdjnbHqc3316MhgkTaeu1w475h5yVr/PPS+/C0yAPB6
Sm7n/dV5q5NBWvlxjVvwVGK2go9bf9YCVTyA33CXo4KxIE1eZA+UABexTLkQ/QK7
0XAcsG0ekj/R4MsIiXMFIi6rQdqyhepJ3jFfctzNTl6B+1qSKDOg63euMO/rPNCE
VoX8f7fq+16PE8b5OuHb8pgiG5o3HM9X7osBXogjkreA0GYMt0lDwcd0lpVrtJhT
98EfINieff2eaYtPeeThs8148dKAWwLZFHVad5LbGD2HkbVEnd9kOcXfJO8uvf8G
5Z9Jg+poihCaPjk0Ggk+35u32h9eNySf/wD4auetqEVT/KLTIoo9PSdP6oZkPQ2X
ar2YNYKaQ/4bvrSWU3lW4GOBJBr4ZRu6OIpIpJbXU2CykGOQF4xzRqg0YRKAIX1r
HG7fJnIMk+zxYdZEGxAAzZ4WB6kOTB9C59zIy2eR+VdVDQMr1L6jJPI3xTFEwNuN
ELlszgIq1XrjRQWNuEfOZ9BUbbz2nEqYxEJoxUaO7ZnyLwvA4L61W4VsWZXhphnR
OawtDIJTPh5M8LVvg4+ZPAIayhxariLnwYQseNPUuOTPS+uXxRvmfRhNNK/eW7y5
HhLdW8RbcjExjV72Xw8I0P3Q2jyCCY4+r8ooUchVXy4n6dVAozYqHgeScCYKO6K/
zXzTtMUU/2ViPv9DpOS9vNH2H56oUIEns7TXyScLNzVodJGsEqVFkw5qIRPS9ZXe
poNGIZX+Ahmzr7evHFdO1QTQH2bWsnmcvoqAw/OUGpxAG3CGIgGFqabwFReKfkxK
sYg8pRdJSM2W6XXWVmBipmM9OzSO7rvYqoz85gnGkSv7ToHfBRTi06hSNut70s7l
dfxCA080bKJupPQpJK+almu6M7zJXbhp3sWYHNcweqQ16biz2fOSAM9EEFosPN2+
IS5YibqjSK0A1lBW7rDvWpW3Fh+rxRtVseVsBibpUg81Cj2AScPOgMweNErNc41c
uQOJ8kQ8SroeYTXEP9SUN09PDgqN5tTnOTM4ojsSoGFaznKXovUiLu0r2Y0vNz6k
C3JuFKs5PJNeE2b/d+Vsesz7j75CMyDEmyudFWgn3hT/VismenCFdTNkfA1ggw02
6oQHvQxlSra+1WXSFc6UVYyMf6QAijYla6YF1AEzFIJ3L/qis27iZCLlhYvOsP/5
plr1cLSBtaLLnDjhreMOEzyT+pkYaMs3P3xF8Gb4faZi0X2u9DdZoxRkkoSNsLk3
eATeZ3J1xpBNbrGlFR3btXNKEyI8wSc7dYr0aLGMx5BUslCPdgGA5wHDJ22QMv5n
Is0hyQQeaJa6BBti7nMMOAfCvybicKLxhzD+/XgS9WFAr5HDFse6Lx3zQHVJFpFq
7OGUJKKhTsIealmgx+GvV3K14steJX0hXF1yc6BvPZu2grLHShSkrGDjFasBCLEG
B18omZda1Mhv0xCvs/pYlBerPaamNAXqJKhG8zGkjp7dJ8BcppPJ9TU4VriXGSec
ci59OY7OVYgipRf/qoErCkzFiRhlRknpvMmwYnqF2ZVNzeuX/85zFg5mq3zF+tlA
vVRh0OxSSD/hwEge8NOxSkx/x2p3+jl7egOOBKs3HNUBvTcw8RHFRoB9UZZDD29W
6WaEAF8tQgnmRRcqs/tQ0fsHi1nNFWCM7e6DIZ3JHiypHxcXKw6l/yNIM9SRlu0n
6CB/O5Tt0HxxN6pQMOWx9vDfu+MbQFBGdZ6oqevxEkgYi1BkM6dHeo23H25s1brm
HvFc+P5Tez7P8r99TAkDRUHCfqblHSjrPPIlbnqP0eF1p2Ab/3OmQGm9VEJEP+gB
S6Ur/BV1z9Z4r6PxmHgE3wORlQ36r5Kyv2IaNAA74huIu4lisvxmOOqLZ8L3gsq0
o6SFiGaH7HVONNBCsPPtQDs6pEep1A7lFlG7uvbMzEYM2GbRuHszIvsRfaByajGj
PeQ/ozdj7pG8hm9kdB5w9wjqKELPhUNeSCDx+Z5Qfy5pz2SUUXZSOJVjKUdIZ3OQ
t/mZOlIGYEYzz26ucY0ks1CSprv1qOzuy/bHOpkaUoWxklxOUexY0WD3uT5+XBik
9XO5mWC6zQSYDUv05uUAAofFd+Bf3SdZdHuxbLrF4PnVXUqD/3P51BiyQuPXhjbH
QGDik61Mkhh+a0VrS2gbkuBSJGZd7M6S0OWpN0SEgtDXUpCu3o8dvaT61ej/OCHv
h6xLiHsfUDkw4HXLzEnuj5Z3hEw3YTBAgZFtssJfhVK0VWarIYlEAuT3Q3F+Ta7v
GpGk/D4dyFUMvgedhgAb/8GQHQsZUFlKJ23bL3za0PTwnrKp80wXZbMxsfO6wtPk
XLrHoht7YDc1sH7IzC2g2Si05VcK2tSUOuKAw/WAOkfrGstdSjZNwKsHplj7Cjr3
PlQZKmkAz377qMx/DZqBFvovb80D5US92ReB2d+xx4CVFMe0250VG64pe9lg3sEZ
dKRiTO9MPnwtb6EAkDxMsGKFFZeuyPDiOjdiCOfFO938sZCQvH3bLLr3Ps83Vtkx
A+8H2ztU5BoiSd4VfLAurrYzgjGuVqMHDTRCMgJOIAimlkveswlTMWnftBsX19e5
RhteYJkRTo1ZwRZJEhyS2+XlcxHmA4kA9KNLXm80cR9U5qCx3+EvGJSLp+3k1eVT
SVqTY7Ut0kWQzeWd5S1lOO4aAJ8AsbRXXwy93zZQfC63kc9381mjgoiBNAhxWIGi
jYGU7anoj/sl1krhYIh5GiuAMLtZO54WN/lCw6z/SFL4wyTmoRoms//2YhKo8nAg
mVqS7SjlXoPqfvZgTDUucdeztvWoUl3XIKtNREZ0eP1HN3iD81B3jZ/Liv4rZpEq
aZw5Uc0vnAUAiyxjdrvRBFv/QwLKCaxMcaV5LXKmDassQon90C/0nQxxELzuwVSZ
jbEtABZM4WwUEz0mXI++bR+cBzNPhnzpDy2h2pKaWPi6Nw3O+8oITCl5AXSjFdja
US8TE8TzaECZfXuBLAiMtNZg7/l0soLzRqGFXP+gqZWtzbRRBk9VUk4JuOov3Gp0
4Nnx0jyYZhjEpMQ5ahVVjF92AvTm/7jZ3B8C6jUo1LEJYVhlZsw+VXo6k1vBNuZv
enqdOWPqNupRBp6a1is/1reioe/q0putb6TG9VB4qwtPF8LcKLLOkGXGwL4BLqrG
J2QZu9L8KUc9iYfREnK93lqeSJYKt+aVIJ1r6QIwwmnBuZgLcjTR54QvU8sdlZ+A
WVb5YqCf6WOfV5EV3huLlbfZiKICafF2sQ9lobJkFKluwAxJKTcQHjXbIGNAs7wt
sSEWwNUOmnUt8QQ3JtvIRdhUuoO4rdSBcSzeZc99um24DIlY2xpIZGR6kAn9quC/
K3jZGFeHH1tV9clk5A0mkLS2P7R9H3d9WUaVtrHX4CCbrZ6Bc55vb9wEhPCtGaqm
GaD9l5wrPMG+h+t+XFMZkkG8GBX7a9Hnd8yR/9ncHYTzLQtTLZQfML4IkeGyk3G+
DzqxIs4rNRsKdMMgctgJMCUU77zlFTgZVFFvTnNJR5E0ZzoRhf1RU0k4ssl8LhTq
Qdt64PhgoVPH8VzsjNqyeqoHm8dCtwrp49MXCO9D9RmlYG4rnsPj+MFYta2i9WvY
Y+fo+TgB1vnlYbZuzrMceOew9uXxVM3NVX9Wd0EgzjahtTr7n5f9Xs/ZDf2qIwzu
pGv0dv+ZdnjFJ4GB2xbCo5JPS7wRg798zvYI4nIvWBKcM6+jT58icgY9X9KOFFyu
N0n7GJlEPJYOqDmNIrRSJtPaFV87VxvMRlGa/s5dW37aXjNsQv+ez0o4Iv7cf0o4
H0aofxHmce9ya+5jCLHLod0H/0dCNAdkhzkVK8V1R0jsuWi1Jwe4UX7EMDDMkdCJ
fF7VRRN2ARWMYagrMgrl2AicXE/itpU+4jyJwsIVx0KQarMWoRCySWaKyzJlerBv
rHf8qe0WlmAM/9qJghURF6ZMytyDwgXk8tWUb2R+qU7nautvwejT9Jz8N1o2tgmW
sP/BCNTuOiuXYdCEzpqClocHw7lrfe0Xk68X0gXldB1oMYXTwYwskJKqZz3yNiOm
0w84UpLlAnIcE3w1i35hE6vhk9UikQ6JRsvFSn3uEjm26sgWmej3aYTFPXKZKu5e
4jbJ46SYPiyNkLFHgI2bxvXORq+QdLxDSL1/Z6RsZFcqdKg+XyKXd0/LGFKnrwOp
w9UFAEaMMbxUpONT4ZG6tjRXIPi9OdCdbt2FTbDToAptq7KN492jlpQ670tnxqr4
Fl+tVwQGG8DMi3gu0BFfsd3LYvoM9RQjQ+n/Zx2FYlgfWXBHtYnW3aWMAohSlBEy
FyoTJFNECo6xZetw1QO1prJ957SsMPjXu8yy0UQWFELXM/5G2KXfLppGh83U4AWK
dRlKXgHIP7DqZjAz8dClN0k+309O8+8lnl8dqD/phjy2szaALZf0K0qtyt+BFEYe
CpaBhZgiu88Pw9liA7dkdRPHLttEo8k7eInE9aPwnsLjLhHKiGGplh9Y6xNwAe2W
vkjtcdEqD4hM2mVIdKLKCSmL6/h3qTQl7JlFlEbIAzlDsE0TwM5pmnlNSzg2cXoS
XRq9eP5e6Z+1zFdKCAbuKOcs95WNEpdHJOKBGpckoiRIvneI/0BHIIR/DpxIFHiD
PTrNp0O9Q51Wp/4tiPo6gSEla1bOJSa6jiPauEI6zW6KeUTP/tByFERi8MoWDion
254fmvPfIL3lbdq8oKaRpiZwnV+NK9YHkcRIVFP2zfBhYZ396/6qp0IZ2FPYElPn
xYFgKtQm7PxfCnmMjxRnYU0U43PQGTQ5Aelo81aoz9/d0OaxtRlz0tadeCCDRs2z
uYCGT7r8I1pDA6Qbc6SKkE3OzsNwW2fiAAcZxYlXpqsr8rwA+uxk+6cRG+svhfiY
qqGc9AkwqaskaAmWqH8adu44oJzzzd0wpSfOf+6SwIXND2x2BbyUxhQDFSwLUs2u
+lPmIz6WqbXjChDxKQA7zugHYgGPXQbu79Zgn64y5o8N8z4icAEvRK9azVOM69Gk
IFBaWPWMKz4uW//nv7hSuBhfKNr8PAdYXR9O07RBwu6ueNaSEQ/mOUIH3jOE2q1x
jOHZu3X/1NgpyYHNLqiQWTsNaRiWX0J088JEB030WeRCikGpjlFIaOusovPD1KDJ
ElwF+9Y5i0BDsFuMuuj3qeCkJD4msIEThZdx61Cl5som81FA0q02MexSOQS16d1S
aX9OLpswk/1zPiv/8pAAQBSST9YFG2r/LKUzui71xshluJFoetGLIXS+ofeuMO8A
7juYNQ3O1IK2yfQ4KVGSRf03zITOnv33yO0v1Y6g96/o2N833vcCmX1YpbT31+Po
2bCBFur2zk1NimN0XE+n+ASwZSWoU+CvdVAvUYMeU5TeK0vC2DzT+WEWpOR/D0K2
TVzat/J4n4QfpvvnAWzmNqu2XB7tF/fUTM6gBI3Y5SUztjW2M6sYNJVv4IH5a9Ee
jIrlQrE6KKxoPDD0rgEwQpn5z1XCFdIwQIe/7OxLSGSsYaIvUNjONbxjSRvtb6Xi
GmfHOkiccJDi5nUCXK99WE5OEUK+DsH57nubG4ZlbOAdolzSCMZCdehGcvSGSpT5
Si4h2xWcCtm+k9cSIUkppm3mo9paC6CvM0416pDlBE+q/ZoPPO2fbPXdDBUjwov4
Lf4vpUJFfshWSpBgnn/pxZmiTHTCKEJvrOuAfYU1x46uCw0L34D+ErFeU1nEMtJF
VAxswH0UEzdYFMJu50ygOrUUUAh51bZOB/wwGvyUeNDKyjUBUkGgMY/+W6BV4U0t
pCppTUwS0JAiWiiyMKXUC6XGzzbv8LLCs3g3QTibh8/5PeX98I1SZd+zx9+GhNYl
BvfqGeCItfIcl8bno73GU5/sVqGbMOUoJEMUbk5b1IXVUzCaoO38wIrWvhLOWE5S
og8mHh46j3MIaX5vor2tPNIB2H9TWLWwRnCoI8CGdnIbQ9OQ0PrVr23vQd5BG4Lg
Mj5cXby0G+iSpm5+MdCNGeWywfdz+ZNZ7Js+Nh5STxM97CnxR8xDZmxUuI8A6Vi7
Buf+jtDB5rXzlNpju4mSEq/JQvbIlqBVdtafFzbY7LA8ZpFyReUw3JvJremzi2jr
5Arn+IWL1rJ8aupUZYBQJo45YL9JIQuC5306ftIfm/hmop8zVBdpMJNDHIqAmzj1
6Ha43caAvsNAFq4+eKa1r5lI3WvKBNmnpJsDScPl5s2cY4ztgxvUNju18OQI+v2C
pvfM2ERqVrN6SasRr9TcpjipYeGAhEIc05OubZX07sz1mui2sOtol4oVkz7q//pz
lmBvdYxmL56Wj1+IF3coG3uBAszxMeJaxLGlLdz8PYPUMIJCK547evQMzPEASRYH
NKaSSveBj/OGEqN5Rp+oQom2mD5Mw/chd+K5buGEALC1rBGDcAHBeiaHqIv92P5P
jYKIrfQyPhFoGqu0tgoViRUlzaxatGYz7s6OoOSRraaXn1aADzB4SXHKjbXXbCMI
A3ZDH+qpRlhQKXPwIywprehDuz2THNT2XlVxLdM3fWRSfIjeyVHZtea2S8boy8de
dfkT3s3jnXlHUi59Mdj1lo2SJrrfsmtYQ9xXKpL60KZ7M95bc/z9klMUCc8/HkD1
V4bruMS3qRZcnjlgda51WeaZUo/cvQJD3cPd0OMtKDE4Xk9R8lsQy3IR7FwXjHpX
gl4RXFIa6UtC/16V8mrW+J77+mYO6uebuRn/txZGdjx2Hw0TiM0uqHRnY4FB6KJ3
OHad6P+LGNd9mM4GynF24f686T5n11VZlPzKj+Scrb+rv9mpFDFNplnuhFVHvY5L
smzA+wwk/u4nq7xzUATM/BhfdPBZ6UGwoUVNzuCKVmbrh7vwSGQeFa83BdMrlgqc
XGi2KfJaLMgXD6FQ28GO9Zto3iIspZzkxTUZyv5N7N+Q2Iw2Vufszaql0Ku5rP62
gMV2LHV0FMXjCeLD0797wLXyosRwveYz/dZfXX760xVuPB6S2R3FZUrEV2oeGqRo
YYdY0HKPupUIl/4/UPU25xOlTHY67O8J0M8F+q4uyJcwGqVKgAExQs/6CtDBJX3q
6W5IJExqm8pET8utzdXsMTvDU8T3lbbWa+ONbrbx2QEFXnj467RqydFmHqLfqfza
WlWnlEoGGlf4e5fzUcRxJwdb6IlxpT5urBLSC8cvOP4gt5TrvvtBY02WeSYQLtrX
xVNDeYKRs7fo9XATo65niKO6Ut239ApE04EE9hZ1Q+2/5lbUjl0G1ONwW5raL6Ta
NOeQbAnY0Ab2lNL74jEBn/ysDTxeJdXG5g6F2giyHi+EdM3To8JsVziK2WZijolm
BSUI+Db8twE3/1kerLoro5ve8RQJEYcB8tFLr45k+KaUP+SkpTdWclR0sfbe85I4
ipChVPo3AugyadabDCEsjeMKEppddZ+97Jh2nNOZWwIX+HyocEec4DYmgaufyIPw
vSt1Yv1kGPpCi9ertomCaSuXeH1L/fLIv5eWgkYTBoWpuKMy1BIEX1xONXBjUJgA
tnoBm4UpuqQkXNK8z1/oJJbETWGmiquCVoItFP+/QRd7Z+M2j4jAEmg0JjjwRx8l
hr7ZnONWE+cS7vhKbHPoSgQvDbOuDMK3o1v09qwPzZrIPmnbs6gQak1ug1K7AfNK
CdiiMD8tdkRVilcbxTXrQjlYROGhflPhAXZJsIfXQthLe8euCDdkj3gKqtMvnSgG
dopxkQLYY21a0PCrXJMRHTn5uY8AhxEJt6DQUAPDAcIbKzvLbQ8e3Sm8ot7ykxNT
y9xwJdLMvI+ADNDYJ+sAZmIjE2mmoSrLts124pO9IpqhA116zE1sEx0aGRj+jj67
MDwfGKu+lweOiPG9WoS9a+saTTq21/V73qQjpkbIGZEwd7HdrarxU3dB1Dk40Hc0
NQTtft7VBA9XWSYIYIl0PExU0542HNGi9PMce1guCPecPnvgY9sWodynNUUZZZc4
QOWGnAHbH5n3S20fjZK3uM70MoKjEFUzKIHMotKglq6F9v/nF/N95k5DKChgBPdm
P6DjyBGtvH7d7oc/vKOWKkrBsSnjfc8YFwz7eJerP+bOvFSaMfcSpD5IHWPZ+9SF
r8l8X30TVFWEoJZerGCA8lpC5AZ7hRWBY8UrLpU3iu688q8s7K2gZLDfgfaMJ0Yv
t2snCwDVIPb3M7lK6pwq+fsyzhZRTLKzYoHz5ChRM9+3dISwKaIyNlu0jeeGtg52
q2CI+rBOI6sSfLHXjwm6NERsEkSCEzghq7Wb6a4GG+m76MINThBnHsHa7rfnViX4
azxGjg1J6OHU9hwBRLjpWNUt6zPfqTTPZEJQ7VrMJyFangoxElH1ZClVIB9bqffL
ZkFjARULyW78+HosKtHBxR2MVtnottnuAHecKNVoqViQbeAfEvk4HdpfNcGuI16n
1DP7C2KV4c62ajUAMhs9JiMr8JOQ5FpKkiP43+n3Kxg0AtmsupoJ1NqqUFap1sH0
mFyCgEIF/rjYvR3CNRNi2yz+cTFKuQurtSYpPXC+X4YxQhbxoL/0PH3NiS6davgI
TdWBB6N0Kp/2xSZQnLUzW5lwamVTCVJuy5lhNIchkPzQtndrI3SeVR9ZUP+1sxTA
BuSCktGKnuNGz2gMLNlMA+sEYCih7iWqKdK8wME594enIX60IySMinZHj6AEMPlv
+3glIXmbMK6iPWuPJ0DPcTinfJfYBCKlS3gxmI1m4/dsl0+xuWlHqlZwlGJ+vRYI
gjywZ9Ea+wtDLs6LdDCubChhDenmSdTWyPhOE8ogn6ECDXRUyLBZMpjOi9zm7p1G
86CXlbdhvvF7X62kF5nf5Ie7DkOoLCy6/+n5e7GnmYYElq0yrZE5IUnxvPn1DEDl
09BM0OttlUBU5nKF40p8gE+2wJXtdQ7qWOAnplMkun0MSrkr170taWpgCjnjoH7B
W0ZPqZSKm/l1SkLLtKSzWlKgdOE2AtnodcDp3MAKoVXEBy8DIxYfjGe+JF2zZqmF
`pragma protect end_protected
