// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oZ3hw5b0334Oc9cEvaPLtjFbsMEJqmXHp7kGBztyYnrBtEGSBus9NwSJjXPiLa3A
NTh5026vsWyNUVoZz1juKy8DFtH0KXtEW+S6h9IXzW7N/ltZamHv3YPg8nwdDq/C
qfv9MTZMQqQ3A7PJwo+Nq3Fdx26e+W7FnU6Yt/4Jk1o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10848)
RrY09G8s7Kpl9m3ToMUrK7LNSSxxB8467Z1iQfFpham/WCMQyoq09Xau7kySyiYk
1e3bGG3mvoq6Ik4l8rXoL67YqXCN4PMmtTGAuNOJk/nP3cabG2jzX+ZXZ77IfLJN
jDU+Q2N0lWZGZKAqt9pojew/L8UGend2Geg/TT3FUZY2Y8MsUZxLvOhAmsA3XqEg
/Oym7U/8rTM32aMN4AlQwxS3cJaBbWrLEBVAbjwmhd/vHOpoCpE6DNgIozaysPvS
AlsCNJSkh2iuVkm/ZXMRM+YeVMBfAdqcYOPoy29OhQxBcDzhTFxSrmqvkHmJwwG9
mp4xMYRxrClh2iGF0YeGlWosmeRN56+my7feNMAC7v8B/VA1PLhM+flsnIe/g5l1
PQvaoT+3AjDuX+TslPu8+PWntlbcp0jYeAmc7yiZoGWYVdHppWa9PuxYelxpob3K
0R1ci5JThTV/glQ9N/1q6Zroz0ngh6zuUv+i6QTkHPFn0lld6lln4kjkNziUd9ig
gP/0qaZvOUNVwOu1FKWOUBw9FuWQWPVQDPESynkWdZcyhcD/eORYlurBzYXu6mzc
d394r9P2zm3/GlC3O94o0rr8glrzdS+4VJNXSqScIH3L7SB11FPnVDAtnO9eWxih
69OLbszz+oslNSbqHXGIX2fjqorbwx1Juj1O6gWWqDKoCP5d0KTD0cPCqi87n9FZ
8pR4LHAyrYT0UElSnP/Qb0Rj3V0yzr/4imS3zDD+O5PMHnaBD0tNQt3gL4IhVAuO
veBaLPN4m0NneZicfgeE3wEWDVVy8BY0W9UeqnmscRCmt+ouNYlB1fFAmtXj9cHA
dUHuHW8XfrEvTPk+eEZ4WBQHoLfnZIn8SJWJXQKjAFsepoF/NgE/Y5kpxiYj6C2d
g00+b4CmuF0awIbzZQqWSCvSUSESqA48rhr+ALI3J7OQu+IyJ2nDoUIRWgRZNKLn
aaJcDq+K+D/DUxoqVFP7NhSJuBbt8CwF0vrgcR8oAkuTM6slV7RXd/sRQqwJOOw7
UTbaqRJM2jkYOcAvm1ZabK7g8fc2Z3CLbBU2XTjSB0c3UWytsS+8/Ul0Kz6GKJqT
MJt30ZOVWiZ8hJzPlDgNAmx4E9ngVTcH4mG3IbIz/RNEAETazOSkU/oKOYobcc+M
n6nk22YjWv2D7z9Nqb4v9B2Oe2MkQPOZTvBVYAD32/QNDwhKcN+s6vZ4SnDpc+Fg
FumatkqU2nozK+PV8JaXfHHiK9UargQdVhvm+AWs0IAPeM5+s0RlLCEB1l6Xux4t
quCQXAzz/zoi5F2DbSPBhs/d0FLxqPYuK5GDE3FzFojhen8/X2MLjPcOYH6UwJ9e
4YEhriea8nJzfnNEW4VU8ViniG3g58VBm6B1QmeBm6NqCv0bS2qhHGcSaI32NSpe
zAuDu6H8TmF+y04nTgbVZKdUYLBFCXMYLL6Jsm/5+fnXw16wi08ogJ69JHg6tRGZ
OxKUpbPOgkrb/Bn8IpUEi4xdMT8Vik/31w4h9sG35Ru1NHhu3ujRgrHhaX6fgssv
KqUe61cP/u1F6Bt1RBkt3dgOpa+7qGHn2mS1jc4Xukr+VprGBat0bAyoueYwHdXt
twYeOd+Tb3nY/6LYeY1XJ+PBPovHILkmLnBum209JeuobWfaiUqyKUTRMuiUm0d1
JvoEdnUiWjsQz3kJcEDZvzIDG0w3fXyI4O0FZAkT9RvOh9/lp6eCCu0vbTvs11f0
hMwBuS2fu8aG8gGnDPYEjVvXpYeF+k8gLvbK8XB3Z//9Uw9toTEUGmNc9n2oJTSb
wVK7SdI0jYYVKfmtzeAX/7fEmdV26pq3SRwdMBNxDOhyyjjR/HD3Agu2GwfgEdzR
hYQH8ph3fLKRJWDukumcdCakdUu/lPi7p2xFgr52dziYi7lfd1NbGWItrRxXwUog
sGolWrWgZSvlFiMlgC3L7E6j1cGemhRYXiAlymOR6a/Y+1nAYYB0jiO8ei4FTILd
hfdZLTx1R8VQmiV7nik9mbWQiaH18t6YnMnsAeWH2XxJYQ96nUgZW/ldto6odoc4
vcO/6EHcSNE/q/AdT9FzcHfkWvBy9Byj6gPf90a2SA+1mofT8w9p62ArBCTRXH+5
GfcSs7+8a342EFIu51m1nsv3uMaK6WrnlkJ2jYBYl/cSPsy47165tMZJWeG5LJCL
zn5HWfeCPrSx5FoRBRZGFq0XCMn7dsEzxdGUQofutRQexbCfZ5myNlfdARgjkm6e
yLmzrJYZmfU4n7PG52we1drzv0QqFYZ96JmryWoKnfr65+ZBgNxZ97SiKakuu9Q+
hLK2Fu87bu0JV9Rt5jFQycyJhsNKZKSPG5wJySg1YjtXB6/Ssqj+MdqCUxdVhovQ
alaaxBEMv6uLD3F037pDYoBz5m1lFg6P6hCce6htX8nldUo6X2xzAfQRXGMkJJ5z
hRhoauCpZ/yu91oToXvlyOMXwyiWFqaaf+He2tshuzCUw/BwkrkSpbsIP07QNKih
B6qpIYrvkgVM8S/HlElF9WEftzOh1cENjFI5IYDwLQzuCcFSCCbNiqcLuiqroe+X
RFu1CZSuEaasaua2kgyEZupodKrBEWlXsnvdK3wPwc4AIzHMvq3TBKQmNNNfMtIm
t2yiGdRXBzjMkpVGLp0ZS4udWWv20Tl3l8LqF/G6U6yxP3lrKJvl0lEnapcADEYL
loD85M1ow9r8x63FeI6eZ1YFHF0ApBKHxTXxR4r60Y38X2Z2ovEauunAvUXT6D//
drnLzJY5ncsmqR5pIjPjm33mC5tQQoO46PUO9IKB7ggudsxn5iINQpOs56SgpsTL
6rj02CJjSNgUe+utIDOpJ+iv2t4y93jRUmxyW1iz6yfAvun7uMAELUc/rEICpxE1
4IZqHP6GSPiYUCz0SPZ++kqaylbiGRKlT9e7PdAUWCIlbRPL8Xj7GO33dwEvNZcI
qMSfpDRu2ZyC27YnSGbJo4cXDt0udNynz64KFZGY1sqIMcLUk3r/iKaQZEcy+WxZ
w75tue5zKJGwWSW231o+zU/g2sDiX812fS5paQvz3uZUXx/lT2VTX4xXEiQxFMSg
i8eEU7/3iP7qaQFTCq0yBJj5jnp61nnaM1LKOZjEC3sE2BZ85uiVpLv0cEvMVejG
Yhp0gRg/Gpu4pvl0tf1qJRsEbeO7IqXc+Qu9BPPcmwgUNqXEnQnDvCVvrqUJgTIT
seGQciGyu5c7A1DsqVVlY099+EuvVX66l7Q/TLFvRkPPQgg6slC+z6gAToQL4WSg
lelFUhUG0RGG42kBXvfJbaTknNlagNTQNcLuP6o4584MuyDE8tyOvTq/8Vf1JlVm
5uCKyA7qB67Ri0n0zi5LFatVKcZKDx3B/25JRXeGrb+OGEYcRgSYvHhtij5K9oOQ
+ziu+xujXiWfFvMTF8s/dXBG2QSQXD3Nw5W51YD2V0D0t8lQeYunHdjA3BuVPVsU
Qrw2JiPQO17wOSViHv3Nif5I26HE/nCXwWwspMtsIlK6Hb5fY3N9hvGe9e/BbuK+
oQd5qWpJDNTnswy29CISFPESmGQm8lU4+YY/0xZYCH1M8KEP9TLSmIVOgEqM9ZhC
X/1x8apfVT9DClSTpImePtNW4y6gFIg3YkBS7WWQ7BOjPfqr3wGjpJAXyyCWzIH3
MiuM6ZP3iyS0vDLu6SCEJmJtRQZIavneaATiwNjvGvmvFxSyDYutV3cu8zhjJ0HX
22472dodvmqLbqNK3/cN5P4u3ABamD8hanh6/EQZ2l1OHkLib1SI4VakL+xdNQ8F
76STaM/0bPLTOWDKq3fBNDmtiOfw3Mex9a2FMSXs8IfvYwqE2HPFPoa4PLjDwNuJ
cJeFlf5hqa4e+13mG6Dr1nMzyFKIMSk50PpEuu7qKjTSEm8K2ifDOEsI6IBSCGnt
nHxvgC+LxDGA6SAsmHhKVn6dwsSBqCNKf3CxIpW7qYiola6vhrgqDGTH4HzrFAgg
X/jxpC90ZE8ux82Qk2ETI6gHACc+2hsAtY2YTOWxyahSMO/3QZUwfO7qqNqlTkeO
mUGJ33PtFvqFEFxLP+dewNZFTqrI9lOZ3exsSJYv6YrpRFaKzYnBSifbrzY7nbiQ
h5cBL/4xuFnu1bV13wyeFUVEKlsMep58bF4PtMYrVXYv5fMgZpw6DWcp1GBipOVU
USTJqBQL5lOypKn5b+6zIVM4P62dvDCP5zs89h32x5MjuMCuXPV962VU3Hqp9Yvh
ovKlS8oEhBe6XSN7ks6sJgGf9SomzCrDX+zeJdW6V4LJXJqCVm0zGsGuOORi9Nln
aA4VLt/wcDYItufW8L3S4tO9xOFqbngov8V6Cpq2c5yunKCSFdDDBQo6DgHr3DSi
wtGtgrdHbVZkyjsoq7BWaLZe5Zma+W98UMjCGYiMNrcsXnVVoLLdeZghT5OtC9/R
jQHhyX7g2nJSiWXAXi5VuZZR6n35ARzJkAQa860IrUCNfNXqGzIwk0SeMLkwuRSj
VO8UY+kKKzZS3MbFhOUJDwOcP3HI1s8pVMBXECqOiFq1WpuXqyt1soFN+GHrUXWL
bgsGGSWmaFUG2NRVYaEjmiDyeYqV57SZO3uHpr3c0hdd/Kq73CFGZ7V8QTfoFG8b
1SppmK4gwq1owmQ3kHCNDh3sCqzVBW+0sViHBO+/Hd2gOth7bMRWoWm+L+Jq9Sr9
qTQQdzPKI1GnsK2Pq77uW4kO+NET0Z6rDJz6vgTAATFDF31A2surRSZHBDU/MuyB
DZNWHSTuXzuosJEpOVlA+aTtCoN6+m/SohCyLO/VPvJKha8p7rtN3faPWKzXBImB
Swbo0pUYWji3ZFXhOSU5/UOZvinNf56gKgFjDYnrf8dGJIEHQC3XgiwJqIN7m/z2
BLOcqYRYY0kDrH1/9CUhaNRrY4hDUOzuiRqu4MqN7jDw/J013f3kzmPzbxRcXDin
HNcqJKC4+JtxWcBsgUQKqPJ3yILirafbXbGUhlBGDqqRrqy9tJpLZbAFLTsRtlmU
rFrN8sW3DPX1Z2UfZDQami5Moa2imSjUJ/4YZgGugRDTumaJpvr1dAyuul8hPdq1
l6m91Pg6XEUaxX7hvdWPbXF8HA1wr1SeN4F3qjksxDXsEcPzL5TeObfreeNojS5+
7hSZbcmYKU8uWajYaldMS5sfxvrV6EKZ+oP1FbdKuPDvEJVCxfjFwGy38Jp8hLTv
DSGGrKkP6eM+K4Lztog6hBtXeNktLJJIBddNBeS1q7jK16XbLx3334Q+YDZh82VL
3hnPbgn57AaePqNcpp5Q02pQuno+1k71RyQGHQpJycsaL/qoFkeppWnExQ/W8exZ
cGYv6SoVz0Rt2rjrmogQmuMbZcrxHqjpToT3pbr9nZNIuFfLdwVuUXmvlvbz5gff
7GM9xiKdcEn9bTpp8lQ8hcsSjfmZh89NDXGatUx4Qs2ryktQbGgzueWmEZQ0inE8
0g436b82zkikoboyp71CKJzKj69f/Ay+2JsuXHY714J0lZUehJkx6/dyeWDaZDYj
uUgA4CjiZMZsptNLGz3628ZEpdsLsCT4IEZK4gKRiKHaCT0z7O7UnIQKcudDFCzg
PCrJ5oeWXbm9RAKnUXo5XsmT6K+i3p2TWQRkDsk124VT910zdvQe07anqLhEGBzk
gGVmWgMX/opZ9njyjETVv9nHnrnkMGXz2aC9swcMPEhB9eRyG+BuIutE/Np4PgA2
jpIfyqmyt6CHrcV/C1rXjPKn7bTJeDri+L6Dxv5spTAESfBGOu1rKYny7JWJ4oCy
u3B23X8wPRKDfa1S8ZxOlmuL+ebRyIxrI33rk1TwwSc5zcvWhY+a8k9IV6lUWT6n
UQbVFZEeAbTqbj3Bnjf816gat7T4cOBbLxFJnA5kedGQ7C5Q/IyYazfC4N0LCZ3I
vqWVw+UWjLCMYynu8sd9WXkBpdInrQ98H5TCxThDYetAt3DjBOYpPgpGbArb7LvH
7EinbFxaqoO8u3WYgPNc3PNTDTcfcZycne7KXCqWgFxP609PPcT9kspbbBs65C4P
55IXRFjBib4pQiBsKlY6iBM4rl54fLBgjUKP9mYbRPjIDCWvWV1gi3Rv1IropzmV
lQ9Sl3Ge4Q6qOqz01vF+YX5oa1WzJdTfW4MqvHl3CDb3Le2iFDUg6HJuvwcx7InA
g2pesytIWhEkGa8au1oUBd5Dbyg2ZqiOO5KLEkUfucma6GoD+a5MXiQosb1aEEXo
Os5g3LMOiL2e+19UZNzE+K2BbkVvfAwgog+fKnI7pdESESyCxLf0N8kH+ZAj4Ml0
F1BHziUFgmynglXyhNpo4VCQ0Ay/7R6e9pLdoEsy2+cDfPFIgohlRSnCU4nt/FSH
zpL8tm2Wc6Ob+W/V1VH3RKob3TzgtPtUQ039yMy0ESwzHvQ354N0fQxNX2wvUgTS
QZSdxOLJKO0TGdC7FLWvjPy4hqk4jpk2V/ir6XlP/4T9OpG7fC4dMm3BbrZN6TD3
9C49jd+wcq7R8NKkz8H6/GOQabMY2c2l88N4tOHp0U6r5jENyIVcpFf0p+Myj1lc
E6bL+RR+hhKgaFUqjObi0mivPfSAf1cdUspVezv4nxJZmCmXJsbwgIpgwUl98QbZ
8graGssh3/7IDx3Fl3Cqbc/n8Z2T3cSCG/ppdkU/TB1eK4PIWKatdgLX7hFlKC2G
B67DtEcnzGzbHICZSMa+xELGR0TD2OwHbb0iX+jhxJNlywheqYumBZnCmRT12u9o
MyGaKF9ZVDaXXIUvZr+hcKonREDNw39K9ESOnuUfDYG6Ixigyn8cRv0LgM9dw69n
osFUmUIa0D9jDjnKiniuqTVie+HcE1B4v9Wiy0PHSaZwGDxbbxedxxwDwsSYy3OP
r6csooXqMPJV3KogWhI6zmXmY2B6goISMezTan9WgK0Norvasq7d+qXkWgFu2GWw
ehj+GiqwWj/hv38/mJTCh7jhfpeehhNDYZkGqSnWgFq8XeuS/xYH1n2BOsNnzv1t
znBH3W39bN6yDReEQluqYV4IWy4hPPQPI2LPdZ6T+pImHPSHxKBJ8pNNEClXLPTm
HXcaQrNI/tTc93HiqfW7CKez3lrF1ePpgQtd5OHW64APZ6gS9Hm08yj2mabBdSfx
bD9y/pISmS2pXYK5ltDf3oCgg0KPVCNQxE+poHenxHDcQFa3gYohe5bWl9YyeDri
53DZKojGjQWMOXkBzmj8oJvI8LykJPzZOZEULJz+jz5PlJBYcoBLbqWDUAFKYnIv
8Hklv49dDX2OD3KAaUSrFjaedlwdDwiQSgckXGji7qXFUBff9yQ4kRO9OeM9X3jm
RC9Jh2ZqNRhCf6gQYgS2pQ56FeQ25dE9fLbi5OQ0kBixfMRSO41al+FLlYnfIsDW
S/mijGJS/YLcnBjPr+6j0hay6kMo7pReuI+VUuF1f6d4keFN/E3GB8dj9omhWAEq
qsUJvEDatRCDRuJfTH08Cnp3nsDfKvZMpcTfeNIboeVGawz4vdJLgOG70F2R/Ynq
MvXC/6wcgs44CGDzGCyK0JW+sNb/dYJYVzcpFPMI3yPCiWq1jecmBbEIsOC5I1hs
Sn9pU3wJEdeLkHhTEBBwjnh/sYtM1C2GCDetduCx6q/TpIsxPVrb5TdqIGot7zMF
pVZOtYjE9o7vonvjeuaHzWdyytQCpTBjBP7/6mZ6PxUx+gb6zAvpAlN8JuSeXNRc
nMXLqCzH7l08uf/3hmBtZJmZirOASQhiCoP3dHeeKHF4fZ4aB2Fed+kDqdkSroJ0
0nGU7BtixLHHgXIDhlFU9+QaUCeJwZlx7VKb/Ym/wBClZIXogd0sQSDa3ePxrLWI
v+HpUw8ozP7uBteVWpbCMY8YQIprCnIxIvxAB/G0ascjjrfJyDR99cRkOpQ8CVTd
pOJSrZVIElDtZNN1xJ4LZHQ1UdR41PZEZL7Be8eJfJ/NNo142wPEw3u4JGV01sPc
20Ac53ODLSo7HePur5QE1oeZ7uoALozEbxDVm6HU4ynF2YnjD2qhZd7VRUyGMjp/
oU9uliqdtyvN3EniLHQhEStuOUIOVHbu+oFAZHNSQR6RX1v0cJL0wMp5WGdob7Yf
5K5bUBG9O3Vick6KM+DoKgInfSW03mO8Qg1XpfivA5KCqzyDGCmVjRvJkEtZGOFJ
yH8/CvHRuTzzXfHsXvNAM7PK0ZLwrJH5yf1IwLhFw65X7Y2Amt+5I2glfdxfXrmP
VarCoj2dJF19YMqtlUGBQL3XQpS2OtccbF6lKwcdLFl66JgWTswO9WASphPS6o1N
wBAGOS9dQQn9FxVe/WjSKjkF+OkAIjU13usJZGKoj3MQK29NeuwMV00BcW7JNsok
nK+dSErIWjNGYfCYXzhwW5ZVDvd4CVqXBuCkBE3oaFQV/GVycUXG92pp8rP8ULGS
0axAb0xk2yT61mf/MZRCDJvbuhGLVB7kp1mcxdm9TQZvjAhR1uoiehmNY4FrIm3y
peLcAqgoQ6idkcXUI4wGVJSAYUgRa3ewQA6hcIwLbl9q7wpg4ec4lkqIHLoStx4d
vQHllmQ2zTivSYRaUyT6hCGX8Cmrj7Md8aQuok1hNBU0eDWXXBiE5S1sg9qIPajY
KAGCY9sQPAb1sPfpjNtftQJhYB1BSUi+fEvYUMcgxnxu6xwlNJ7y+s6n6SjIF+5t
yT3Co6K+Ys7DU1waqUPsLPaUfvwDP2WaDwTHzpiiwZz9PVHo0xRVGcAGFWlo+bMv
yKPdb2viPASB/rw36v/wue05v5NASe/pDGdhremZNUwhLTsLfQKY3kroLzLuzBTJ
TCDaHizBo2gPp91rJFdHTND5XHPEJuTJQoYiUM9nLyrWsJ6b/FuEAQ8F6GFC0m45
cDgtYWz3U8aq/jb1iDaSPtyY5+3kgEs/nwXPqxboCjckavaMARlm9fWc+TXUaFu1
jhEMh/sUk9ILdgHC37vy8NoIVCRTShLSkPjk6t/LZl8iuHlQ5gFVM3jKPw+NS/9s
3xYzO5pCK1Tg5D9rZp4+wylj2zxZx7ZgB3nDGP607UJk5UipVVxGu1SyhYe9M3a2
aupRnzKL08xPAjLARBFmCmbApNfFf6+x1jBxDitG2sNyVg5AG/jNF2jX/pLG/woo
dvuaqRcJ7uCL6bDrbqWqr8Qo+95ByBbNHpIoVgA/TML6/Df0euJWMMnLbbBWps1H
PR04ZGn/a6Za1X+dGhEGg9eOZT/HXGQocrUy3e01qdbDKnLMYqczuy8W83G5Zsa6
8qg+avj7ak2xyR4s1hLpAxIwmkISNSZH4D4HHFDpq24+HYasfyFEFPuWfYYYxapc
iTcI5GEDnUdQODRZhZDp88uuFP9qrypk9msT9kaF+5XB/lNJbqyhtVfCZf1ZfL/L
fAhV+UMTWFOuf4HzQA1ffTQR/Nql/aDUswVDlnp6abnTO+8PWmk5ccOF7d+7F2ga
/lrwyApyqiE0g8TTo+Py43ONXNPSXzzR70ZdBQEYOH/Jz08VsJaq8ATt3JniF4Si
CCAf86cnGoOe05Gw3FEBxO4Hbumc92XXzM00TG7bhjJSv80M7Z9rqd/SuyuUuln7
C4qCExhfNmAX/D5lxoi8QRsAS4bzwsT7gUdpLUfSrpYQsUt3d7FeoJ2RKvItGwX+
sCFdcaBpeXMN+bstiRY2IyuEfPSi7BhauUu3HVPZEewaarqKhAXJKd4Nq3NBau2R
RjGRG3QgCitdE7/Ih9s719HLtoAwT2MDnNRR2yjDincZSzS0oJBto+KR8WBYSiyp
jS4H477e7m3aH7Iggudcc5nmifBNWAafBSaydoyAeuYaRYBWhsuQu9ex5SAxOtqE
B0WNBZFZ0pXbkWrTcMYjmbKI9c0CWlcd6/VRpvjcfOxW6NndYGDQgCk/kYUrfRQN
7cwSUNvo6eTEJyEpzQDY9MDc3JC63kmZY3/uBSOCYwrU5d/XGvdCJDIysaF4mxIq
Vf8hBZtIhjjR/xAh+GZXO1UWoJP07u9di163vslj2KEjN2eFqEM8ryeRBOFKw60h
PzbZMJTYJqnKkHF1qNpbn7A+2oiuLdvJFRHHIiQE4DQKeVDP06delbpmDrNijqLs
7dZRMf6HnBCDHrrYmeGmrIhFjIwl96TSZAGhFXwoZHgHe7Pi8cQXnUkrNfM1kaT4
1BVrvsysQyIByTGknV4nUC8kmsEX4Jkgm27Rv94vrjVXQo0/lEFvn2dGafqQoKJv
GxteYtOzIqYEUYgdJ/LyjiILUo/ZLrQrsNBoFNTVnxZt4UNa4J2WibRreoba2tco
T5eKJJxgoYknanuUZQSncdknK1c4Ujlib8VgzRzZlkfo3+YHjAOALw1zP79srPaD
lyFuqkbpFX7uoKsr4EBLCHYZaN4ZRY3iftI1TKn2p5HLdayx9R8wg3mZwszjW0UF
koqjplqkY3mGxObKGkS6CDhH08W/lpDaRD0plOdHdhrIEEVqNGw28tnfbq9ZTQDp
2wEDsiPZ/j4VYyO2doKoqe/bjphYqo56QW+NdzGckqsliF1h3ZQmGA3o7woSbGPF
NKMF7QKlmfTbjxP8jYpGzgwMzvLxjG5RTdWOUg921qdo9vuZNsh8i5oIX16MJBw8
eIvSdkoasCg9NVe42zO2oTsMyvUwhV5OfawOVIHjGzXrqyQcAw4lYzbyNFKwtcMP
x6U4A5jbrDS0O7e+xTU5juUsUWsOO7iDX/m4M8lhmyo6L0AMkyW+PbWQ94zNkQ5P
dnlcqxRiiNiSqVmgYMo9Bhior79QR0Smo6Naov62wzH5o19fO8ZdOb823gWSy3M7
zwrS6P8rKyNpeBbDDXHR2Wkb7nI7qMFspUcJ+740mjXXqTORqH+fWB1VSkJ98SoS
XWH31l8t2Ytt254tGpr+jYnrCSa9OXnp6pizLKw92iOKPWQqOBHhXlpkrFmctcrf
XBt6UwdyjvOUXBvWShQTiL2XpLo+T4LzhSXqTqx7VwF/srk6Rv5QcxmBLPId3XMg
ciHMnvoNJ8GCMa/gndJ3poTIZbYJ81ILjGYtd/TTiv5L4RdEOCFRVSCK5T0iL39Z
g+diYl66+YJBqVpe5vx0YbSYw8SBu+W9zo6B8bz5Kws2RxkxIA3VGqd2d4rEujSo
PzR1Q6MwvkRUZs07c28Eh7YTxvdkncR11Pkx1aPyFSHGPxZFiUXaP/RG+GSgA/Wo
WWF2HE/ZVRyfLKqz6NKzd5RClEO1LIaAoMBMDC9iJNs+VTFrokKTBkCI8XbNwxDy
RaldcRpdY6XNOUBsjYglNSqJgza1oKE7BcC9Fo0l90lVyhbsS7sHZnk/c5Cb1Qjo
Nh22Jki04bin5tLERS5mhmLHDiuq/D1YAnJrC3B+MG4gMox9BX9v2s1HqLYpDi7W
bUiARavnRzWi158ph2mudWp2rBa3bZWNYI/vlBRdk/FZE+bEzF8b0Mlqk/6eBNJJ
EXOpxju8J1qHvXYo5Q56FPoVPvYmaOyPztlraOGwfpx1WYYSrylSKk5ghhcp2cfI
DQYGgZqvS5dPvqCk755tmRMhIRLM/NX7zonywORgR2x4nLjOhHten3Ea2048ttIT
7Ia+Djx2L9i7ydo70/DnHaJ2pP2R9rmWD2ReRMWA5Hh5zXtsldbSIFmLhh5lzbEG
N4Z/HvzG5ivSBAVYrlPdTLXA3C0Iad1ztwX/lhBc3DOpUITRn1hV3vP5n5XKW1co
71UtT+t+TNlVn4WasQFWeZNqNKfljoKZE7gaafSQf0RP5ITEs6FbwM67NpUcKgNI
dcQVnNTp/httqdDXFaNEYqLvs1M95qvjMcPrEGFkJnMIWU8HhP9X4jcphhoFuX2I
4lFvr/04gcgUNaKkHODxEh707kTKSZE0LZwfw3HwYNgeSMu0/G3IZ1wY6r3SQf7B
DlLBf/qKVTGhY1W2S+U1/fKDGPl+F9b9DCXuXO7sVAxk2KOJ5umkP0mYEzMk6NGL
R9A0qcGKYDxwe4XFOpT2S/SokciD2WsFeE0voNoiPswBiAy6e4edGpIYL6BND/QZ
rvezgyma91ZUNsVjsKP1qEdR9nCWnV4Yd3GKrdUTS8THrhKyPAn50Any+kdlMjyx
65BMAFzeECjURR+Nq1TioJYUTkCOti/t8V+0qd83HLjQ6kpR0F5mvXRTKHXe0xvL
Ltmdyr6zFTEq/n1ThpOupszMgP4H0PfoPYOX1zls6S8gxozpgX8K+K6mp1jBtzxn
qCFM/G60Wn/t5xTHpqeySL8FVWa1JrUk67tYTdeNS9KK3R2Zb5dV5SAUo10oeyN8
pbFcQe4HLVw9o9tM5iNzpFi/F2sJsJAVxMhIMEY0fyj7kdLoo9+Iv/mNLMyD+8C0
aCyZhD1nFDjvr3QvtLH1fGZosCpGPucLgZJWCJ9yVUFYZmcJgOKmjsfUhMu7ffnI
HmFQ0bkLUVmk6RWoEvPqaP0Skn72qhyBxXuR1u+slr/bbsZAo2xabC0r+1Tc0jMl
tcxISoj25dPfJn1XjBOzIaQKUjny6ryZ5ezBuQUccvzerkkm058qZKF9wIPHEhAG
ANHJtfbEeqaD4F3bOu5E34wSfls1FTVsagzxMF35h71rxjHYzR+usGYX+MiWKNb0
YpOp0X4O1iFoQqf10L/ItTu5pen2bfHA3i941/oPkCHn2oyS0IvJbSvFVEBmSUnY
KnaQUGiYl48SLPWh31t3yLiiAat0WggKbWIFdfIAuEn0Aj5L620WCOUnoEWWeSpT
T54Qs/r1ulfH/A/inKyxW1OrKOx0Fz9CrV4Q7foxI2mv5iz0+18rrOYqxoMg9nIh
M82ND8/W1k/hVlA+tXFXPDku2+agCtSX/5EjXbB/E8/10qhcPYeV1Y9UFNXVGL3v
wVhx4W7t67j5ST8T2Ck0BLQiRuTbzX27UwdVFddCEtmtKtBF/0u80iHOeZTMkW2P
0nRnUktlHdpyQsvNq4cJORctreEub00EK01n0oD2KTBQVRJQTVAf9IcuRqr4AkYz
dTZM0dXaAsjgpMQEd3Sjpv8N1qqAqGiy5DkD0MUobtG16GYyAUHu+I6n5EhhBhzH
dh7rycyIYlITNyYxCn/v2v77CzLL0dIKBhR0zsR8YcOE+b5OC5Opgfvu/73lzuUn
QFSmfv4d4XjXEor1vAoBbsR5hB/L4Z59PL+iV6xN8WBa+hgolJapgJzE4qlZdBI/
IndrezIrpx3oAn3rKLc9ImRUBNM4nMQ+a+lwbw0jABhc442BhNrfH3WHSMWi3cp6
KT1xK8BMCxshKZlFB9n/uihKLrEwS9OzNtCwuJdPf+IBSyv7q5C1XT8MlP94OEVu
hN9oEGlau2nYGw++wT4TF7ONuaSLr3x1TsADahshEBAo/O7ahb0Dvd7S0c3wzY0P
HBoe4Z+bzOCOnHsFhTVaf792i1ihwJJwbqcDgjiovlNDjW4HwT9sVKwW0/1lL1Ic
e1S1vIQVeZx6pCMF4RJ5SBiEKsL3aPw2F/UJ3YU7swQbaEtHkLxTW+pqVuDjXNj8
8oZaaoxftJTRMGBfooOndkZsq6Yb1aR6oksNtdwJJmlES+XKiTBm8KdVFeFFoinw
hrfCnKEb/v9N6das47SU2mGJDvzd862rBskI6nxx0voEeacR/1xzDJUBRaLvDQTv
3uFXGqC+hlOr05BqXpIbR5tW4y9otkEEeIL1UHLMBGh0/BBaKvYbe7eA6c9gI02i
5hALM+o5KRXlA9ji8HSHlHCujaq4UN/0uXR9TLMN096fyRUe1wRo8fn/h1sy+5mH
JcIXv42hsJPxn3XPtZnBDR7Xdw9zJK9pLO4HbitJmJotVv+PrEbuQoECEOljXU+8
f5F8oZCnoQBU+f+mKH5t/FyhHN/UZyWuQ1VEDvZjvx8r/vxY5XxCJOtW8dP+XS3F
eZexpZftwXSfEI9H5IKLoUAf2wMFd4vsyRQ2X3+xw9No++it4gLNVSgKsH8ibqK1
pHl3m3RQufMq1vvPRhplpJCpSES4/HN9xx4ds5xBiDVh+/05uCtqR7lSy76G26Uh
utkq/Z3U3VBGUZlB8XTuhiFps9W8ZPck/5E9xYihRqqi3fAvGBVAGYfwuljezZaD
/sanZ7twq9YkdofqimLq8EqmHXywAh8flCo1DPVABEA5MJAPrBh9RF/voZecTJ/9
zdjBehPps/5IEc2MvokxJCLhdnWXzyrktBZqDLsYIXljWJ88ucZwPISR6MYVkYj3
iNAW9WWZ9MtrDdSLCS4ALDa7BIZDeSDURjhEVIhXkuxm7raqYHZ5WU/8twYvw43m
Cm5Q5Bp5ykT90KjDJBw/TDPwPQZN8Ci0/HJHUyR8P6+7Ae/+7u0rIS+SplNgBruK
ZCKhdEWCRD5RQPo5Es3DrzAGAeOSULaFpGSzhgoja0vmddPF8vpW6UyBugLoyZGN
QhsDpqQQntW/mO7vB9gemfEmrcSZZAt4opI3vdO7N5DW3sPGG1oA7MTPDGWkXCy+
2EGSTTXza7hPKprxuMRteH1yyYkSQsVr2tFH90AiB8BlCc0XFKRhKNRwbXiwyp97
`pragma protect end_protected
