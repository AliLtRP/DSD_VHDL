// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
OyCXnhsHrTNT2MBqbcYc8JsF9rbMAzdkLuG/Bcq0Gb2uGwZtWObSW7gxUxkxC3ulz+9TSfrkkql+
hQvSR3rn2QeeGb4ytSBkXaTETovtQVgng5LbTff8cPunMAKPdDrhDZiYfGkdIKMSNOuGUz/lKkiQ
kHQscJY9YRtCzkuXA0kM75MkTGdNnesIwiw3xRtMm8xrTtXnsg1isiZbHkSgr7bm4Cm8SEymTboE
KNFrGBIzTOky4kDbVhIgOfkiasNyievMG2V/0kYRXnIDqk/VeUC76eJTAye0HSIKo52y0M+CFsMq
U5Bg7R2mcau88hq9KRVT+nvochM7pcBE1BWCgA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
ZlScGP7XPBDqkrRIw3IXZK0PStlOczGUxxRKEt9gRgwKMgvjWY3DWDg/+XnKHRReqXJwOp7R2cU5
ICa03Bw45esw/TGRtQS4iRieCpNiUeMliSuURS5CSlaxSo+qq0RMSXqy53wGLDKZq/2VUtEJz+Tf
cespWN6tzAeuhKgT0yI7/H41b9pqcGeYgMClLTSa9UFigzrvTeyAKqA2I1oAuEKIZXijbXRrOgsN
FESy/mJ2tbelf1W1fsYEofs/GnLkTVMtSn3GeDyEBH+2qH1mDOko5/tc42YZVqblWE4UDUYDwm77
anEdGk+c/Zat8ZVYTjByRKAYL2TAhRTdHWHb0JooVc2P4r3+68aXspo8gqzwQVeYqc8KkULyZ9gp
5uLQIhrD38tiLOm6U3DSC3NxhjVgC5IJTtYvcZCeuvMt7KQU100QmsEhEihShL6AXqup+JOWB4OY
CefWRGIgwtcbODGK86QFOAVTSGBXK3V0dktplNAKxNiJH79RyVZv4ntmIcEsNsepw+F/N6h3Or+G
auNcA2qkbfvTBxexqeXI+fQ87K+F1Zl8EWBaqQLBhhhOTG3k8/IH66x9ePRT6eWCka7hfere37Z5
sQAxnBLIUFxmEBJEyPdAXZL/n8I8gj+OiqMTJW+AEfGtIlcrinxhC+cHLii/9XWHa2YzaVtJmAnA
Kyv53kc05CksT7g4hjOVAjw3MhhcOj+bNqImvNpaZDqzPkmJ9mnUI0K4X/FiGK/mhH3CBlXhVMp9
2i5d9HbRV/og8TcsBVNtoads9hwt/4c/XXCnPlp8N6IYwStKb2LA5FvmSiItJleANpwD3zZ4+aAs
jw5mHxT5FnnFGgSi894Hs6c5Ou8oxWQP3UVl3SHIwPirXjMNi98na0k9b13wF4DSI8AJD3J47plQ
e9oO6mzWBKERqS93D9tcYNX2i8wmw/fkbIOWtorDZ0ESvwiczXPbeacglShq7j506LyXFsVrJeRN
b03QlR2q68ohltVZGs/RjLr5NlmQurLLWZJ5p3rROve2D+fcoNrDX/C7BRNrVuvFldpEGQBD8bz1
sKG9ms5N3YJWrwVXkgYU+cCyxgorOi9XxP97Wst3MMj0/LmbJUy7TrDxSZg3ubyVyRp7Cxlwm9+n
nBHYcdtFPje551OZLGpkE8B4W/V2Sv8YztoSq+S6A0gsU4toErHUYDfBSfQXaZPQXO2sFixtEkyU
jZa5j9OE1IbAJQ0LdVeOImzUPp4++BUt5mPw6EgRjYRfaJ/NXVSzEgn4zQn0mCotagjS5GlJeQI1
4vMQqNDajc7iwnGtIa2YecP7ILqC5pPO2DYE71nzW7UPKVZuQwVca8aQsAVJDTWt5Ah0mWkxUiwk
TT6Mu6Dlnu3eUMsAkZHaPcyBTfYgSIRFCE7gY62xKPN6hcjTSG7Bg+9kJv/gojEFFlngeN7+aOXf
p66yUv+8KeF6TV0eGNGOq/UWsI1fiCBfth7YkJJ2ICTYo/2nyurw52DQ0ls/qC09O/mGMS45mSGP
KTJd/nRG1ou6KObHUSx5uD3Qe4S+a/iduG2vVUMbWSnAdTAdmByXRoo1YLgqTe/r9uFaKxni468G
4JLzPJtE7FYliGEQamyRzocebTzkTot1R9riXgOYEUukb5CGRavcGujyiyJptAZN2wE7/6U+N3H7
Hb50WrmKuNQbepRuzVi2jOAsl4rcCzy57VIoaWzZBhmhnT+b3jF3Af3oZBtXhuLyYSZbsuCrg6kD
jYbyPLraprxKV01GhBEyPj97twB+njKXhiE3QyVTJ5pfSwQuccGlklwkukTHDAGKZDfdqxwfksrj
XM+LY5QSJPfYFIxTT7DV3odnJyLJjqtiKlxAkx/QC1Kmcx5//Jdiv7AxfIyGC//0Fwz82a1Jr59Q
joeNUDGlbk7FyXgdr7I5XfL7W4/buiWcE6oDS4hH0bQvS9NZqYJAX6FUfSCk+7wry7EjW3gCiar0
+VIc60fEubyS9ZPXkAd8BJkQW78JzfJULhvoaDC14IL/mSvYm156+EV2aZL5TqGSKJYRv1ZOTJR9
+zwYb+GwXO/Tu5SqFqrB7BHdXnG7y8o6m1b67BtnNhEkBkmZw6kmVjOQN3vgnocrM3CCNoaRaixA
XngSQuTESjtPPX9AqIlZSiKaEelRkPVG9kXrmboZMxxuPUu7iiVkXXGxp9PEig07mf58VGyvVw3h
3k9RcT5YjkAbgYdjjUKRy1w5JR0deuzAXZONBU9oZCurpju5PTXg3kYgUgn3YwoyChgumyPLbbtw
vanQHOBQmZAmvQ6AstenREld64aVjSHX5NnDt6Gej2DQobd68jyUmv4dHzw1guYZumO8lIZMRWKp
BG1B1L3fCNQyIVaBbZ7Jf+RwOPN4uy7AA11kghvESiOr/Nbczi0+fhc1cOCZm5WXWhahLMreQvJz
GA9iDlvT6ziKCaeGuZa3Ir9775isK6DlcDr0VlOYWVHJrI42T2KrZN731LPkQqElX0gWFM/6XV3X
J/xdhjqZjW32hMYlILFR8WZc9830qvgMZd254ZKmykISl7QeylaT34KCYLXDRU9VSA3Deal3Lfbo
ULT/nJ5UIaW6mtzyFYH0KWDaGfVKCTsfU2V1ZQji7KYTCMmS9FMr9uaHGVlvu3JsmSgYLp9g5KAm
ldcYFvoJW55UTVdVenxXN/dpMfX/ziFrmfe3SlsPlN/+f04dMHT9XZBSlmxXfCIxbNRpPmd4dnWi
nOhV7ml3ug2PJOwLsQNzguslEqWwcwQr3oWEPjCyMSWVaOZSO++2ggtrcX6HM/f5OdRTbd4hBlLA
sRM64oxsxqmTff6+c+NMf2iKRXSCBqdELrMQpZG54kDmgSaswexv1vLdG/eJrYN8nDuCh8TGU4kc
suhQze6IT5Y4uEz1VSG3tKlKeBG2GDhcF71KBmk+I0fkk0qOynwLbTJBYb3+9RUxZKgEuWfljyo7
fbUyiAbpk9T4eHA6dz0GrzJJjp8g5YXaxnpQwmh5/330oghBuBn2wF48KrWsj1iOzGVZikRzgC7o
uhqqOM8/vzpkWcasKAJGvWtLbi6yTIpO+AJ8gT5RG4vuuqKeDveOU+Iy28TBw/pTyf5iU6Jhy0Az
jxGSf7QPFd0PMdPDshCP8NVC0xNcUng0F57RnXFEIqL/jLy8FGPgLAe8mpPnZj3wENjwgz6xlR03
+ytUicuEawW+upinHRDqZs4T6ZE4A3ytnfNMef428vlj3AbQhCvWsUPf1QrJxGjCfzG/N4oIDL/L
geIofjggkwEbROwJOWBQ6dhNV/NvLrewCZ7/68xaOwvnlPP603mektiZI4LN/JjHvNjrlAkcZMuN
EAw0BNkaYaYaeAo/FWr/+N+PossQUv5/FzEajsYvS4vgruv4OVObK5F3C0zj2wUi+Tm4SVCFrjdL
py9BQsL00Nh4A0Jg7mODCxg//r+B+/56e/QyO3wYQTb7LFO9Lmfja06FK4k46hxifF1N3p1CbIY7
1Cz4VF+wCJEjZVvLlYEsKHpfnT/B0/21Qrb40PYmQjkYurHW2dZDQyLgObXM5dK44mjhL7TiFRgQ
IR45OvorCYTtvY4lnMlh23SYiJmN1jN5B1jeRo+F6Op8QyX0qTJ40ihQEutQGhqz8oWyQOaTPtM3
nuV3dzN3ZxAGqNQjSVQDQlA/SiT2Td2JQv7JpjeW9aAAJ1qYfuMAKq/JRfnung4KbKEId6pMiskC
W5XUu+J+PXwWW0jMnp1HJmovUElrEV8ZLO9liRQ3rm3LBmCxll1nk68SNAQLAvmZ1uvuk9CpnP7p
6DjTsf0z6SPnsPT+2f8DqMEl+veNad8nmFO5hySTeQYicZ592qMrhAMfPQ6YajoL44W2SqNUPXYj
TbePGVncCnb/y9IPszIYJHM5AK6FZQCk+1uRZm/Tyta5EDWEsfiVlJo2I+vjF4C+hichVfcDHKaP
pLNukS9IGq2ZHkHXVMLpKkCFepQLSkhLvxlO9hw0nPtfvwQqI95/XZgdBi1EStv6ZyC2eU4cDbtn
xVYVJsVtgLZOt3I5Gg9PWqkWTX+Rcyd4nuSKghD3tZOJGmsGSCavGkSpmzdrxG6DyV6vBGaW3bVw
DlS/TCDatIAeI/ucpntKyOXXEeUBpZcHcStSpeeaIXEn7t3GBTLt20JitniCHV1ptXyRl1ozUlTs
Y0yTZ5hXV0ENPHAzKMlowYYQ4EpJwyVC1MwSSN8ObDxRb4dihXX+Jj2B4Iwc4r2E5pLxUBqFZ2Nz
JY/uVNhP4laC5MdKK7+2jdHF0RXUOcvfFXHY4+MDs+vQW02taX0A/GsBTC7PjTMhjqheKvXcqPN/
5qnXko0Xl5f+dAgufyhFcrLrdbmgGdPwPJGUXD/9vW/ItyshEG6VdTPaToYCSn1R03JKE2QuB1+N
IN/xUL+o8kba9YWI1nngKy9oSaNtdmlnI1ftzxuTyj1sZ4t4Ve4PJxWvdQtomEuulhzUGnnGP3T/
IgT9pJZEkHf2hotgeZ8Idkvb5Ay3NQ+Kpr3fwh/WDW8XPMrCiPcanysIW/kFUgBWRApcBxSuEH1h
c0xqf4ylzftgu5FEUHdru9+IvG6bSWr5vFrqtPuTM4i4Yeq+Zfx9e72XO3hvwUPqwGHEo8MNVlQh
ZiE+Espj3NWwuGtEAhIjnlcWTEV7BoLjK2vC1RXMES3k84H/cuU6IlwsELd2VYLrax1hJqi4wdl5
Arfs7K1i1rU/FH7ZaiDNoiTqk4IFWsM7QbQ1XgHhTA/+iCk8fy1KSHyXi+F84oSkfkqdP5sl9PvN
wELHDLkDpRadV2PcPOm1Gsy26SgVPVoiDehygAxYH3N7WwZgT2o4q//5ItNo5qfqYw6EJ8otxlrm
zCpVejxBRSfLGJbCQ8o/AieQpoNqLHDfs4uGokdwfWyUSgJPKvmxyaJATS82WdcyKl6C9XM8XOmp
Keg9TygcnxTzAjXBwyfUvsW64w10BDApyiGgjXS10woEy5Lpby68UJuFo/f7AndhhGRg7iHG6BIW
L4yavGY7KZnv3+xwvIg9egI0xDGZSALeLCCriGLXgMHk/ubp2HxTya3bTBYfnUxvfJ43EMxOdutL
1UpsHszQTf3W0AJCxVXzqou0sV2YaPJLjS+Y7E7JqNI9UXPgd6sq2cMdbTIq1xGNETJX6rAmXpXa
akmHnVwtl5KW4yoxSKgbEz6S/bxTjvOhxPKzlgHBqYeOX1tF5Wp2rqDHrx8h/B4JEKKitStLHqRb
3t33bh0pnb5osPIrCLduBF+OMh1RaEUChBHvsnMKFHtgXolfDlkk38CsRz6RhJSn2Pg+HfUlVh9G
DlYJVS5/COB0wDuIjZjFfrH+vWgRA7NBTdTy4BKPAqIp4/ZNgixyefYhArn5nM83ZABPPu69VMQS
WEPBqzPCsvZOGm8WfPAlobuElmXwaWjucnZmEE2TKMwT+0f/H3zl+o9okJ3P0kFDL+kuEqWuiQOC
81Huf4lSSoaLolvxSwKTMjFrI+/FUl95vuxed6AwGh8eEDjDIDG/Ax+UcBVZdoXO7nmt33K3bZcS
wq69EhR7XT7nbLJyuRILmCuSP9biPgEAC2RpzIUlsQFlxILwy/Pgsi1QkXA6fEIU2oj/XVXZBXSL
MwBBjJ8WlG+rdnqJbYb1Mo15YOzJ0RVXrV+10FVWg3iL70RMPa15d9VZYugA7Q4HmAyRwOO7wEnY
zsVhx11BFOhcONHm9EFfFvShdMN0Q3zXQQ/tNYYFB5f5RqeVf6hpkCjXSd+cVBXtR9l6kaUqKahs
MIVHhV3ORTKNQE11DfoK3ZW0TdPnYRt/YWWrSOkBUc60ec4JmiHhgsd9goKU1Dqtx8WDDcpmp/7A
3oayeX/jKb55cpaNCiwN21HVKQf+TEYxTKZFaI5jun7htGec5TDFA7epNKOQBHebsdRPLwuyrauT
lmohTGeuZrM30b36eQzL5X+/4QjWUsGj3nUlpgJAFWaExAaq77CU1AzOsP6ipYxbzqF0A6Hy8lnj
38tmQyvhBwAdRRc/MAF3sgYtLnpKSX8aADqt8mtg/duf5/JKdPH7IVJe6is82M2+RI2COFYTvPto
gGKsTas6jiZjLMPZqLRBlC95n61xocz4OCbDecH+wAAR2Gov93aek+ErHYa40ywT+tFJ/A2Kexmr
PlzNcGMf6S+8+oh6YbWfyJvr428fuh9McVrOE1R/7H2VcJd6SbOeQTDQb7ekWSfXPQ42TveZugdA
NM09iizccWQo/BgHArepZZO17MWfFx47AltJp/wWXADwy3NOqveAuYq1GSO4YgKQU3H9xKhAakH/
rm5LoxNwrRje7ZMQLli3ZFwVAmIZk7o0ff4emCZaW7qm5zHtiP7g8QpA8ekvZrSbvbhLcwFApZYr
t3G7ZnsWA4MnlWaDM0HY8mvXYdKeQuoZ3Xn7CA53E6A4ff1an/MW489r2ZiLWm7Mcu21ccauaaxP
iiahZ3UOfDk4NbM3mHYQXbPXQ5AyB8lXE3etwGws3uyrg4lUMX+cAmAOjOg78Lf0QBnGacxx9NoJ
AGKkH9IUbewsM8s2MoH6kMjaF4TrLWgRE9ifGHPkZiFEJniICY7A9AysWiw17ELoJ8/vkV+r42Pz
XfFDogMvxPsvDhj0oAavp7z9V1EI4GCqhjofIYT5AGD80qXWRRLP7wNkqvNO47I5E/F7e0VEOqs3
CMqqhdxzVQUVaFFKfDegogDXNJ5LASVUQ6SdUY4tegLJ9032APeZcjye5rFZELu5qBWXO+WYlwo+
20jYii0hlFkEWevqFTKfUWHwfcwHTJni7jeEeLNy7SiW5/1LDbCDZI+qkIK0YF4VZ1gwWGg9e3FI
MrJ2/kk3s2NL55o7e00wEprGh4Ls7WU1hfE4Hk9fyjdJYIwT6OPp8q+BnG83JpAPhcufd6zG5tME
h4hy5E0Vch+jlFFJKYX5KetofNr0yuvRXr94DQdMfHbNkJoS4n7DBMdyn3th+tX7T2SIw72xcPnF
/I+rhCaVU18Rr0JrwQcKq6U5zfnSthXNKQSfvjvNO3DEPeR/gbpGAVYD923SmxQ9IzMC5MSGtZLy
wRaBgGHG5wZXkmPL9zLGtVNN29+zHpCQSUIeptJzEW/C8BsMu2bvBZQObIwdk/+SIUZbR3m8iiVe
ll0TuhhV3+CJR1x17IEDvNxEJ2kTwtKzesdDGONN8tOUxpxgmdRZUR58WPmNC1dWKerb4deLZGCG
O51agjrZZEexNMnVQ3YAjlD5NMsPeiD6dU5DwxQxwAtadoygfVsFCWdOPFqDHF/LV911wh6H1XhR
2FIhVLqU1E1f016/chWFhfll5dpdAD0p0YYrAAESPkIepDfohlcYewuGzOxW8Ut6x3OLXGGwGMLl
dt9kUwSG4UwG+/ZY6LgvbDwiezGoi2A1MWwq1wKlLUFc7BKQuQcYqdMm7opH0jxeB/o8OnYzeTfM
m+InPdo2IkMYJ7CZUzPquNmaE2ZqgOPkL/k43hDS5lEndIh5k9bnollPB4+LIKCgrJBXrEVvEAPG
czoKMeupwCBaOuPQKVQ1cZan8BuSW8AQvzR6eTbtcJGLakm5gaeT2HZ3vFIpo1BgJpG6utux+Cbj
OPrwWy5rxGS/6sJUYMqpWWpEIiqX2miD2taz6SjooYwvCPLLKkVgyHEyADOjXOsnHqEpUMXaAW5L
mVPqTTxDFQMNSspKgrRrbsFTr9oXYL6Bx0GLaVc1QC2NsEbZRm86urwJtJD+NSeIWj1ssmqlEFFB
T6CnXHsMZLQx9SDI1IdmO1m/fSveTWn+NFkmSmyYYrxnOrp37230I5NHZH8b2rqaxkE9of8a5uHt
I1q3JflJfftFxlIr6mc8DrFdqwS7Qdai2Ls9aa0Gwkz+WIVA8uWdMYcvAFPRuG+9X0mFMn9Kt3c4
sA/PB0Du2zRgX+Gg7XN/ndvM8+4r/V5rqejtvwifvbVqxoBd7pWMigsKn0iN4J0wYZDVoiqAxNvC
LQai+Zs0qpcSCRfcRb2wray3nSqUFIARZj16sEFvKdYyjbhAQ3wJwKxbcCxSrgM+rALjWAoVmk3w
HUN1bqEJnTZs617fEBlD/agqYUNOM5R9H9zwk6ztm1v3pIydpfSfe/9Gh+BMVFl9Hq9vG7Np4HLG
MHFvmim09FbDgr6T8Od7nVQw5a42bzNjCM4fg/g0D6Sddo4N9wUSufUQ053K6+qgI9/QiL4etPzt
vFOhODkUrnfSXTFbG5SdQ6USqB1UfcvIbzEaxvKO2Q+Hp6z+JsnRS4B4yyNzTIRRmMVSHCw6ANIj
F2MqhGqWdd6KvU4Ldq/zlH7nfP4Ev8EZpBVuAk7oipHvMerNeRtXS35RxofJ4zSPfxOTkpVNWs0l
aqg0D4lieCldsYQJL3780kdhRxdHqLRW3RfNpnRF6mHY3PnSxx4OJe04tMNSVaurxM1SFBLG1Umq
wzCQWk/fWfQUtkRix8wrMDggVxv0rkQ80NSa6RC1Rsd3ZFapdwdUhInd6lyQOq1ZjJpunK9E3TC5
sYf9uiNOYdfc0VWLOHjBAAQlpJ9pQOKlRMwnAaOhjY/79qDkfieDjNhVEBLBMFUArvdkK018oji5
B9omrH+1FBBNFTR2O4EmK4ijqB/hd8yZv0psyAJTRuk8QWvNM88oJW9HTq67czra/92Uo2AFHPnH
r7AJo3wCpreUlMNenV1L9ZgdHDqEMaDm+Ms07vWjOp2pf7dBijFEYPDKOeUhJ5BIFFI1GSiZb/iy
Q4cJCg0ktJenJG+Oriw3vqDj9KYICYdyDuOqLHc5e6P1sB0fH08LOBlxqx0I2NoNoblVn4gPp30b
fpgSthww8qWjgaQ1MyDRMq2CZCOH1yn3uuyMEKaRViOhPMzyQDbD5TKDP7h94wmJ+l2l6rK8Xcto
4pL5ny2w+In5UiujHGhn+AGNeAu6Vm52sY77NTDG7IoiBDG7TDgNulI1XXDY2OOZvAUTWMyRbxru
cImu+OBypP+MnYa5si3V+m5pxBM3/ilrHL1F1aFRtcIkLSjoYTwYlueaoDX6AoO8+tRmALHW7go2
Lzb84LABH/Q+99PTHGFHC1DmeHxJX7MYPwmVSi06VWF+acJLlKKloKu7+Xb/6m3ghR4wrEXSWRhn
unOJH6UZMvhaxoXLOTC5iDLyCcd0x1MZWKSMgqacxAdo4KOcxYlsSNMxV7jqUMMnc9xNxBhS+FQq
Ey5buBeW0YKUFqaxMAn3tV8jBBUnYUqms2TK8BQe8tw2lsEgzEUFWC7DyNrs3nDKg1KO0gR9onj1
5Bm7ZOcxJAnuseoKqYHGWt9kSg9xvE6my800JvwH7hHeP1hUxNR3dOIdTShKdo3GO079/yLyRbaq
37zqF4atyHmwpV5BUyEMC+YXCNmkJruiJSNvAgQ5G01msG03uQOZmV7/1A91SqMPhE4Vya7TOzCZ
Z2xGQAL8kdhoPt2mpc8N69zNZtwC8PzhhsN6FhyCyMBTDpfp8vIgCimTnhH0JtH26QcU32MuwSo8
iUEvmxSCEbTZ5cX5e1Kncn/fgAT7Mok7lPUg2/mLp8G5x2xU9wxmMt9zf9dE30zz2GEZJj0GyxHh
mjnK+54hD5Qq/Ocx6QAnjyKrUbUZK51q7K6GdCaoziocqCBu0yIoG17H5SPToNE9MeDPyyUKrQ6T
40XKZ849+Wy0DmR4Bk7lcctdddoU3LdZ4uygVABwAS6jmaIGYlk26v3jDWVj9++teOFQGr6Cji2H
jsgQKRXr8O+yyleSCP7aRdeLiIyg+4W+IuJtTCQ2/6Qmf6CEkpkqQA+pRt3qtyVVn0xjkht0nO72
+BojoPUTUnPsvk5j63i8kI/TweT0i2dKxA7gYmG2XEA6FOXhsjYTCKawwAEAabrdYRcdXM+WTNfk
URjHKs85Sxddx7z4BKK0mKyJm4Y9Yuz1gdS+ZrbQn26iAypHOrkTGkcUmHEsPLkBIFodS/BYnzUG
W86T8sTiyu9zCYwb5+/LA4G9BXoXY1b4mvBBFX0TGNh6tfCSMlLndqWobRn4wWlWddTaY40QOaqX
qKHFaHY+9Bg26eLmsVs4SL19UzqWbux44F/50XkEy2AupG48xju4pYIzWeOIb9L5NJmIvCzmtxJK
e+XL0C43rWsJ91ZTUVttBGwELupgSVKlBY6qehC1OOLRcSHvl7if5mNtybTkkZDXwN6TrzNWCZ2E
ChfShTeKEECD8/xdlaeUvUKXOcQ+LDcnJVpeUA/qH0Hv7KBeOv5IRVQZF7/AcqQLrMtbfEfp4Jz6
upnvOWBnoIrAQM5Zzf/FUQrTuJsEqb2gIH+os+GrD3VefAz+yW+8tZGO/UNISYd8FZgsSPUsfyPF
AbFVusrFBVLrHgvEQp3G/RTCrz/P8mflszCJkuPirfx25CB0MHJ/zvO+/mzU73wOznvXts0vRKZG
pmkh4LkWiwLUQVpNupVK9sxJWzfAEsx6+1MDPlkdxhSvFQKC1YXpKmwXLyLgjO45xP+z+G9zzV7s
dBfdFwzJzABsGhvqjdVEimT1H3xKFbMKqDXEAkX9T6VC3RRr5Qno2VitsTEaizkvlUmEnUxI7N4N
ZC8xbrQiOM8pam6PmAIwDUbDgGlUV/u8c60ICJo8VuLl0Oe5wwBqBBj9il5SqHBkGx1x+9GcLZVD
1J9WpShOzUeKQ2NTNJSVs4s8DxdNBe4YUMIWnDGT78dkuK+4edpTtjKTKzX/4tbkLCEAwejP4+9O
TOffIV3Y64CQ9y0kkax+i/tKQZKtZ7Qz9IcJkJro2VP0kQlohIovIakoOzXoYNYJfDLRlesTeoE/
QRMMXlYDUH2RN5JV5sqbr8jIKOiq8DbstyE3rmAkzZgIXqD2b2Q3RNeR3L5DdkIKRa+baAEqDGMk
0wQb1eC/dBOvne9sL+LxibGSj1AbIdDzx6el2PsqZOnLvkr1jXk0OzWHvlAxsh77tH+DQeaXvSIO
OXSZ5yJwELK2Ett4nC2ERaWeL9XKF8DeBxPkK7yNMkNVRmRZBA02ATg7PloRi+ZEOcMGnCFveX1i
rBcLilpsL/FL4w7/qWRk1XqYk0sxZ84C0Est1vnCnioMOAjJ0P7PXrZampV/Ojp4SOuo1jYHiaIu
8LFnj+NT6czf8aaLyXMOEoxgpulZg9S1IBGHuhzEyCkp3BYvC9QAqmFr+9DSfj902JYOP3MB1o9I
baGA5AEsso0dfYB2VHSlVDl1gM9ItnIb7XY7pIPmL3E05i7KrUoXpQeWqyHbWTWmjpwKAT1QHGTd
fJjP+IP5oTFK2uP1+rF7YfqiYkgR7a0TpmPJlmu05mpjfC3FlLO2fHSru1mDgsVwOGnrT9OJwdI3
+aadu6XmLN4NNQVz5b2Fr8F2DiARZpIv1+aFYG2o+ty87FFr1fVzBilVxx1pBSG+tqpqpoUPKMtg
onsQiSY92v4rfHC8w4thBzius9BPvfOsZKTT/e8O73huGZ39daevHI4S/tLAgoHRmwqqEgcNsdBB
NPY5dPFR7kWcGlrHARdHORfRX9ViDVdE6e2xMxq1eVkHUSCQgE2lTNBTx1sFWsbh3SHCQjJ+Wu65
yvymbvD2fcF7CskdF/mVagfwRRC0krDHkcQeJhDXQJLxKRsHnAxCdkYXQ8kZd+igLnfR60X6mMeQ
DhkwPSEx05tvVywVhNdYqIwqkk8kXp0UN63YFPrdhnxxHgjLb2rsdvD45iyhcSKzc6GCD67Pmu2u
Ov/BOR1c+bTWYdBJVVXhAUhx3zFXCKvphrW1I7XzbAxvSVFdCfipfBhrpbrbULvn2juibYfChrTo
R4zYgW9jsr0ZjkbYjZb2NRikblZ0Oj8u92smZCdj9uQLpd2ul/tyE88Ild564+7fz2IjZfC0o09f
iaX+wgSnDu/fs9wqALqjW0cpPNNoMU3efkjdRtsF8ThkQ2pAUqgPHDx/QOGPluc1Flh8PdVlJp6I
xGZZ/UC8rxC5+2hNqmiuQuiLds6x2yfCU2alm6lYBXoI7q1IeApsEi4r5lm6oS9gnFnISI4FO5Qi
l2Lw0FHk6Pjct3Q/q7ub8/0/CSn+//TPMl892jem8QDmtt8bUUvRJmEVjPBEZ2sN3O0=
`pragma protect end_protected
