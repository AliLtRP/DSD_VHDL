// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:24 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OtDzOYosPtgT0Z1nSbMs0P/kKB1RdqGcflQmzR9qMwtX+7Pp38BZsvrUmXe7+06A
MnyMB7fqoJhJTztLtmYyGssnfY7lgoE0QL7IKYFTiW877OU9bodgipgrg3LtXQEc
qDVV93flyfAHSTDE6qEVK0yui/0YXcWKTllJbx/oyA8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8128)
+q9XZVMiKzB+peqvOEsgxHC/feKvB/asi9IiY/vqus7VOG5d+jOugEse78T+Ppwo
/ppHZNcIGl0dGDwc2dBt9DujF1FcxaG6SQYLhVb7mt7sxoGLNEw8pStrX5PcVIra
4+c2mJPaV2JFzFTdxoXfidb4mQytOJlwrAmR4V13Ub54M56MYcwxoV/m1dJZjioW
ia0PvEre+KK7TPqF5l4qrvRcI+9J4lLmadjXzGQ+5hf38t9UdR94A+9LVzYWpLcJ
UEF6VC/QU56lfRLFHBRgubHLOZ9eKC89o8k2eHkjqAdIJKlXTzIDmaU0PcHXRBuY
tQe3F7poTamqlORDK8zrKjwqXkx+YZAYpeHDQd2cBadZJItvgX8lSn9LoRlKgQ39
8DJW6hzSDIybkMows5yZ5qHLL2KD32JtkoHcmkCqjEAyx/kSXdbFopM1a3aX2pNp
hOEVj1lrNWTA4OpjvJoe39GjelC0qteBYqwF9jq+Lcnc5eVZu2+Sm3dASiXifNIM
oaJ5ieeA9Pe1eFfTnClaf8eFwltX7w2zqnp9GRRlTZM0DtpEJd4ZKqzBRXuj3KD9
WGgIwUwjSrF6lL8R5bjRhNahWlPywNSktmkryEdy22Q8wWQbBtpcYKElJQJWfbWj
7erz+qCX+kmCl7JlkMAqWgHUSCMW7lkx38Umq/YJmixpyc2FIuCSfOy2SNKDC3Bv
HbrUFd5l0VJuY2XUTx2X7Lws33EuPffDmuUaLPizWBUWuYXIzPVMsqDe6KxFKMJh
hy8Nt7p2jvM/3yyfwef9xRKsg7gkha06Xu6C/kTSVDgVqribJBZcSvBc+r3Wc4mj
keGwKuOtrRyuU3Ekz52aBKOM0F72IqmHtXSuyLNkRxU8ReDqq9BuWulJjkYe8+gz
dPaQuJEZLYEgcSA0V51FkQ4q60o4rJu1jiM+4GdiMdn+pU8yOANtOXs5fLSkE9Cs
LRRtA6aCUlG8FLnTyle09XY0jbIGGPj8db2K3rMIVoswoyhVQ0WJ3mav9ocU8eJq
2ggaSartpDshxl7HncDRAas7mBiNJy23J15v+AmuOKwZUvzcuhhoO7+HOq3g1gak
rIDQAfWgEUbSVSP/OZ1jpKLvqoxDz9oERIDO+TAcHje16zxwAcGFg4LKiQZfWGxo
f0Nk1EoJlp1PP5b4ZuwH5unFHRwXzuis3P8ENL7hzW3ENH9ansRkz/QXlqRG9ycy
pEWUq4fwE8Qe8gQ6LN9Xf0IGAxswZluLLsYu0eiDk07fIOsrTHTMvk+2XVTI6DMv
NHjc6A0/+dZ039WbZaQdS1XaBYH31C4GkIdX6Bij2vqDoiLErvIHaL2bDSxZAWXe
+6UuS+JIWFirKvR7ILxPLco1fBEtaoh9R2vyTIYEsh2YxsHPKpPb+oDR39Ie28gj
/wue1rnridwXPjve/weudX2hYAkWhbx7TQZGilfQFoUMunmQtaJm5tFMxyxgooe1
S9e7Q/qfjHaOccLi+ns+Yy4qXpLf0WQqdcD9Yx3MvrbJLji/UiLT5VCPxgU1RSlu
qmFN/mEPQndKJc7pAR6imehlREMduhLGxdMVpKDA/5kDuqs+/wNwLVeWm0od7LJP
TZkUn8qMacRFDRSYnYXKdRSIpDnq11PDG1kKOHERnGWpnbTEEoiLQjQh2ahMlMtR
HNAznJndJucfCgx4KI6aLOwWZKmX9RNUaqf/rATsCaDD5h5Wztyq0JyNDi5cUH2d
WC37FJ53w2v8l5kiimNINfi+P2QnAxs9g8QIEjqLm3gNTgCxGxc39G30it6IvX26
XdfUegoGZLERyfWGSfKKAELMICyaMoon1iCKKMtDu6xAiP/Kxr9zIQfvuqHxqOmB
LlsiWdM5PFkmW9aSwfjKUve3oC1aXEMFbJKxee+lcdRj9wwSdNdbK4WGDoLyoybF
VIdoHEQRRhQi6v1e1Ku+tt9KPXiLtqDFIgw6N3lilPhzcDzzzgIynmPlyXB4I4Kw
+OEso1aQwEQ8NKwQ7/Rhs5f5017n/DOBZcvTmw8f8BzDyj/vjHG+tE5WB0OPYc8H
uCDwvbmC+LxlIXtk3uEp8EHe6+Pze/4XwzO81mHRR62wV1NhFFlWbnqB/LJWIEHT
+eo6z0Xn/wzg2oKaLjVljoPScz+9YKb8EWK+1Mx4us7bLWvRW9NuTYhbS8fo7FpU
FE2zFxa4PHURA1dLB4U6NNZJGrue7hRSNhkxrBcTW+4QQ6TyBIGGvTna8KtP89+L
6CDO1yA8l/P/yf//Ozg6J70qSQQwI4QtBiWWtE3xJ55IHm3V7phmsHanFNEKNuZu
Opp3TYgVLKQHJoBx+1LiB9opY7yrfXjTKUxOfVTa8YESGQ5Ev8kbdfxaVM2HMILj
VVy4QcaUgWQVfNKPyxQqe0jvJCQus2pkpPOnRy7zhhu66P5v/2kVSBz+Wa0724Sm
dcg2wCK035h4vVZ6tM3vMwzY7shDDfhgbNqt9roYN/Dx3pfRq3C1g3qQ1YxeK3To
jwoaTSU+R9yOp8QJwjasZamG/zVwihkU4PPH1VkoFzW6DFu7TaeI/cv4bnhddmJ8
o16STsyPc763sbbf8AFqe35vfbx8YiacO2UxGuHGt9GTEKGe5ZNayZDskpeuR4Zk
+x9HBCntfz2SzUwt5yEmq9o7OaGkww/NVI8d6bH8Y9EvGII/xGU7tEjRLjBs6nAu
jEgzyZf1yQwJjtU7MT7e4xpNml1SRKXYiKAdySTahBfe5xGnt6d0NL8pLa+Cxq+3
puFK2D/EcNDbPyrnziXjOH1BVOiwCmUankPeY8byYmdTwtYgn080PU6gVE8Qxso5
PWGW9cjiI9NgaowMeuL6/0WN3p9xT6KZwTVgiafIv114qaKZbk2HOnCniKaVJ2eO
YL6fEV2yvx+wTZMk1SVaO7Mz3mum4le+QMkidEJvFehPl0ezvhy0HXRkZ8T1Y8SV
8I3c6YCvV2BuvrXdQLDCr4H8KDZ3Ij2udxlejK3XNccH/mfSdkSCiNzijMAKB8g4
lVfvxvKaZ3s056aw/gnSCvn4z25YDkuElutRMRaExLS5s7h21H1piBlc3f2nHI1F
sxCmYn3M7qEYvSVrKQQuQbp2E7Yls8Wz8IkWCllleaQw8OIiOxt06Gll9VUViwVR
bI8ZlZ1MJCK0fAPRTPFTb9Sl0blrVKaq63maX64O4IS9Z0UsAj5zqATF32eugx1F
vBAhJY0s4isCAgpqvVigxdaHHtGv2xnDghEt+PLP+MN8ZDh2+zZEX/hYoWxjbNl8
htTh0ve4UuG+EDkO1k4ZYWJ12rAov+SrlQ4+6rC/eHaLxidDl+ztydutSB30wLoj
k9QMMv7iLe5bwxEBOSEeWDLpXgR/Y9xJu7cmWJ+ltyY/PmymczKWYgSAvjd1lyCh
E3oTYoMFFqjO7RFCxPUo4HhkPAHHCgHpK5keKLwviYVHioDpynFfHlYbk6i4P1kM
MGxDiRdkLK+i6OpAcsiyOMDibvmeSoqky7w3+YPE3xidNfvX/wrB/BdU6xg3YsqD
tp68DPiZLKQUNITfm3X3DupyDdlqA8rMA7p+t47yMXJLsdwoE7OvGCEt9VL8oMBR
riSlqNLB8tjDO+h8KWlc7sAArd5g7vD3NAiC8BMgWa7Uc40i+Zddg5GvL4UzqA4r
SCT7dG4yk6CLm0WoyIWhRPM5uYzji2zli/41H7Ez6bpie6hGviv7/gUFzuQIRzaE
wGDJkOsMInHpnHuyPALIIVeNRo/w6mkWejUnl+eFZEexe1AyRa+oSDVW3C8/+9iP
IxXy2w5wOJCnTTOYpTpfePobiM+btOyLsFT78qIYs98zH/4Q7TppuK3hh1yE6+fC
xNf7azK92x/xGDEWrajWInDVAUsepU2CHdukELIoZMEuSdW3bqnMowVQRpAIK/8T
RZaTtZvK2SDJyZXyzUQro7eG/giNbbQcF3evXwugk3P1osdlQfPuQ52SFQpO0j9c
Y363hnbfFFlXA2nRvSxeWqCAorexbKq/WqdgDuZN3Hye99616IttobM84ar3Gt5W
abENwSj4MHk6QTvQk5LzaaKKzg7X3KMy0f7Qao9w+vj9eREV7tnfJFwZyGK2bbYR
dgqr337PlrSWAI8rrEDFP5y1efeAgLOSgiRjTlOWnwrzQHqIlwKhQFLPzA8kW+8O
3iuKUakKQ5Ei4GA3Tpk9kZxdSTvZ0kfc7cM+gohTBEtSUm8/NO3kLd2pWC8FsZYt
lNXeVvTgmetQA5Mf4BBKMXWJmqv2hvG329E7PC77eifYJZvr7PI7GRjP/RvjoBmR
88ihPskLPgIfLNNDWVjG0a/Ijxqr9ZMssEqcAcv4sZf+MjLnouQk2zXLFus3IJSU
KxWg3tiCmKDz8muSe7zx6Eb2PzSQa+SFdJcJkStCRCcuGFymeABaYDV4wK7Cm6Dj
5WkyjMY68b/7BbVPfUkkvY81uYeiC6zjnJOOgcbhYX2DbUMBcu9gR4Q3j6rXwGH9
klLFBym+gpd6ZyAiX1SjLY2NeNweHDZUDkSK56uaSAkJAjf9jJVlxLMHOPwPbPld
yeTS4yyy/fud5TvX0GL6Ptf+kK6Aw8wlCvUiays++5CjQdCECigsDlOIJczwuzx+
jl7dfWPWjB9d8Gd/WxFPvZ6xSUhvf+Ji1wwdQYvA8fhziZZADM+NmT5UxOXQgKGZ
CMK64XjXiu5I2lKBZkDZ8eqyd31QufWATWxyNJ2Da0vVZAsYpVIjefkiYBEoEfnU
mxXcnSR8nr2AnHN8g24uSk8ypmM45PrnszHCqcTeuMi4AqfWb8RqiPdSXzYHQjOD
ciOmD6SVhTR7P+chOnPr7PEAxYQ6F76uJTZ4qFpQcKFmNEI+7UKQdDFxfnEmracX
mWvloTMiMvC1clS32EfiXTqo5x0XLgRUnlru/1/8ggois2QFy+3VQcPz25hhomw+
DXi4D0IaVgr8qLs0m5ZySf9ibI8M49KPw/puYTd+T6eNVEDbQ8Ic7O+8eydku14x
NbCndIctqCdGgNM4/iJpOqsvsCiKqOvrK0A7nYhtjmMvPDHeLWLSHh/2MZ5mNO5C
esTHzrw/GJSTiGDXADMtBQOYV33ZFc/cjpxNvqEBEEGqHe5SRvdyo2XKPCylV+Oo
Vik8vc1uriYU34s+eY/QMF1kcQuh531NEqewls5BiNCn60gE4tz+uCFg7oOusFxK
rwUlm7t7DauX6WCkEuqxhsG6ZCQSrXeLYi8VlS9sqt1BuOXmxLQpND6yQIdzqJeR
+SF24LWbXdr2RsDrTP8i1kH/7gHS1BnIg0Hp3FVAy6/tgRMSCzashgAhjBui+sXk
OBuEgpLOBRU6XVflGdhdaoQplqpEcD++Ga0dzK5vkW726lRlMJ6uvtDbm9fUoipP
OonIAvbJTA70D88kaNxTbw/2zzTyM5QC2s9NH9aWWn1eTq+VBK6oPIUxEm1CmkWJ
DdPxjSelxyxzEK+ZDaAA8Th7iPeDOGlfXBAyWSpzvpns6TALQxb0hhJkpT6CRaMA
GALKO+gHnOeg5tZBFzPH3cujKBb3tl2x8sX9llPuL+cvOaj63zRVJrTx80pNkfvd
B6XX9VHvab5EfbM4ZpFdRY9phg0pdd2KJeXI+V2duyo6hDmTjX3BiQNWJcBsG6Zm
7qgcINnCtJSI7DLW10tzyooe1Y8GTXFVZQ+aZlA5TUYuQTBUTfwI70WixkgOd/As
Aa333ZI1aAjNhMtp8Amj2jgaoAtc87Oc5EVtmFJ5gz04L5sSQNgpzjZj/rmHI56o
BMEQ3NSNq7ExXu68T1BWXqX/9hvDOFIjnQXtdneYbD792cIr+e36+2rU4UHx8wll
PwaPllVVNMn4q6PpvN1k283swS5bmBpC6NPII7YzCvO9j1Ft4thZb2TbcnrzU7ut
iLq0kVuBn/Syr3yZlG3iWzwonNx8O5wZkU70etLx++/uRMlyDBz4WRUi27YInBkx
ZWS0djkx3EI/8845Ob5yGiN+UZ982maxMOJR6lqH6Gj2pv0LtqM24TJ/TuzJxH8i
NOXCpDi7vWPWreW34Dh9QOj6ylp1XrraJgDtrEs89wNa48jP4PqgrhlVe9fmcvyw
Zc4Lg3LarkJtRMVZBuxpPFaYajv+J1JAnjClD0FUHSj3ozw0mXo3sUXvSDBsCVqO
0E8C4STFL9ag9VlTB3z8FX5tSmfJ3tQ6OCrdL1Oaqbrz/yCI3UDDaC9ZJ4klTmWI
0+0onwqoKO8rkL4V4KDTA4yd/zoRvLrwRxPneqkn9ycj6unY37n5B7XQqOXm8ewD
A/fHHBfoRzrnCKZKJJHUdZRCTWEZVEnfV5DGj3DhyKWOMEJJ5/pqvwucNctfwcBB
VFg7aJ8mtnjPPXLV10R+7uKj+gDY2AtjTu115P+tWMjzXpJZmWFfoYT80axgT6RZ
l+QpT74dFGSWuygbhMyPA3SzQT1/JjdC9BiloAW+h20OWow0zxe+vIgwyL6KIxpR
Zn2HahqHnmvo5kjo3ibspXk532xH26TKc/lDaFDbT2svO9L5aRGWgb0RA68eeA5d
CS+Oc5MtCMjHJjfIEeVVU7dUhqF10XwR4gtDeeUcpejqYTWIHmdBjn09TbPZ4ebk
ZV9rgWo544JegHdE5mFUvM2UkINkxGIALRttjYzctPPQU4ZjKFhdP6zrQtmxgvKt
uKKy03uLvvEEnFQlIRA4ZGOLbripcHs+1NiTDIxqJjfnGQbLGvKBwjbgDBS+59Ww
jag4b5gndlxP2TJyT+EGLtDFV7rjoDCz8wtf1JncOt9X1HejHJU7EuRn55+OE9Ty
O07MOOTeJj+Sz2NQN+v8BiFgn9Mvv8RerClkf1tPcETvQrtidJUzRO72RG1OMmDq
ubxJ/4uKJ3C/jFG8IHSgQA6+/IpvyWXWqiqgFEls5lZWXJRVY+ceH3Kp8oboaFDQ
hfHqQn2s6ZdQMAusvo8/AjnzQIVqR4KSbsXtnCe7QQzz5BQAo1Vx0him2Rony2Qo
xUCPOnVN1PMP/iKb0TZeiN4j1X7CP6ImVzng6Xr/ZnqTxx1267lzhs5yUrTi5mTN
2w1ld3ViwGVrbmahYpcLqkBSHLSE9vCbXFgKOiQcEMCo2rZmS1KijJYQWypG5nEs
2q27/AsFn2pOmP17BDDln+2/zi8AgE/3IiAT9407p9D+zVhLpO8b4PJv3Ik4pYQu
+HA4tK45K0Oul2y90/+3uAMb8zuhn+Hiv6beBaObsRuzMcGW4+hxijyl1u0mBH0e
axGb83Z5wHIAhu99E55ebt24gIVLg9XJu+xAMNYfM3ODG0yGlMwM7czTTofGJuyg
NBhCJ3ZAAR4Jhp9Y2ICdA2nrJKMt+/UNztwzxUzXLCGt3r4OTrIE6VR9/vvCZkWI
pdDFTgq+CldRY0KgkYlHplxsTfi1UfVs8Ayl9GnTaEct1s+dp3sbPM+l3DSqLDDX
AB9ZdXsJCgRJSD1evhdUHL1I4hsACNbeZPQHLafiez2Vjjd70abEwNw+6Wd05+8h
U4BixX2Zbe7oJvXqZPBSPNvtgUUxanTYSU6mqH4+Rz9VTjTT1PgEgyXc1wszE2wZ
0ABOZW7vnFOPKoObyyoeQDNAkz1TbwxQogD/A9EWlmRSIeXpeVBLWTHoOfsIExJO
0NTbDojZLfWox5xeIBnpQ1qk3X4WVD0kNR9OCfHKuIkPKGmLyPC5/13niC1mLuGG
MbpdJPV8v6BxPrUE3PMpjUON/h3Dr9BFeKwR6v04KCTTnhnBU4g/mutqRK5gM4Ij
0U9na5ly8t6zwI9qIpH1Ie3a86woSicrNe66dUMm+mf5aUjdynG6rJQwj+ez/amK
BP3h78RHs3PZ/T4VXEkaJMpT7LIcMYQBsOPRIhQVqG9XKzS9l5UzOtkSYLzOtGXL
6AKASy2A9x9oqMSRNvXk84sw6d2pNEd891rJozXtaLE1TM6FFyJpmCr+PyHIk4Z3
iqojee8AC9KqkxlimSMwdIpQQZqvWS4vKTvOtdMJRLHQUci3PQjbJcY/wtzTAQ5C
vAjbVatOLP3kT2n62CfVHcNUbJsTR5IqjjhUMncjfx1UZBa9PJCjHtBfvrpcB/1o
VZexkWJ4HHqob+Sgbq+j/E+Jv1vWCZsxpzpfBd3YrxObfUiRDlOXdwz5pBcZyz7c
Lv0q3K4n/+LzRbQzTYbDui3JQG22WDPqGky7CBpNNgnWwlCoKM8KWyteJEsEdvqv
+0Ul/oOWHr0MoX7VTeZTkYzvqNQo7CJCA8g7+UmXJwAL9M+z41Zgva3IsBr3gUZF
n7w+jB377P4sRIKUjDjbzMVTQh5HWTe0dldxtappJ2c0bibPDECkCAnjX2hi3EKF
OvcY023je9s9qFoRrZXfC70Utk1dsQ0ZweRZO7TUqNwu9r2K6mfKLGUgXHT9XyDm
XUUxKXD/0/9yGPZXlPMZPPasdP+NRVpA22a36KDZvq6+d7QfG5jaZiA3x5U+yVJN
An6waTMu29dzoUXnyk3AAgZtJGYaODNGzFnlLaIZ0GuJfuO82+rHQEK7OHSkV6uD
aBx6ks0EtN4+z0WvEiT6NVR7eSbLnA/MWIlibeXfcj8Z1x6AOAx1mVVhXryWKU7m
tUHFjYhrWnCwhThV36qnN/73Zubkyarei04HNYW4qYxtc6d9wrbP60Dwt9r4i8XY
fjrFk26NSdC8tQ62OW945uzx6b+cy8qqNvcAIeXtq4e9CGdxohyTAsbpV1OBCKNg
LXT73CTZ769QLDMz7WPz1pBDn6y6XNXiO62HOl03ae8z5fY0cMIjJHOoFSZvt45c
pFFktIPz9KoRAXnYtr8McFvWI71Tfh1930beKtOokm7GJfCZqIFWekx1jM67Y3Lh
tyJ4DCanCLRSLjI1qN+kctahEXEVabjobB/vZ8bkSnOcOTHQlSJG8DgZZPEKUhu9
V6TwGqtNYma3stv2W1VcmjHIQpGyFL1wZYpPvgrc236b/z9ezyT1RVuElPsMZULs
8n5+ScxJ9CfcWZgW8giH4qIExjJ4OMyxm5AyXn+zO0D/z7BmqqAeyfMkPkNWgjnu
heR1I1VD8h8rwCKgr/wUzHwYmbBnx61kYyEHoSkrIB3nWR1127YIbbg+35qOo4NT
+Ba/GpQEC/WS+gV2BCcXdWqGG5xZvzsYQFgfVMxoj6jeg1+jDi71mjJ+bsJOFz48
yYH2QkMqa+90wEpcPQhkl7mxgn7lXkOFZuHjH7xSpCm+HhhYepJgf7HunU2KnjS4
OJ/WGXyk0pUXSsoyPva2lyF6hKnswLEsHgIAxRirq7Nsz8kKfmIwfasFu/fPXVIS
g8m79PO9ce6dZtK/5+RTQR5qG5NnvIl+FEJzE73BaoVNWUyzmT/W69pjZkjuat1X
7TIGIahZ+OMMFFF5KmOrBZDPcS92kD6Er4ifla6J4kXD8hQExg/n1BWcRXGfl7Xh
zFVkudHID8UY9Mcgqu3IrjZKdIz+JQSd2NcZgEiQdXDh7bjNZTfeEPZdkExWVK8y
3+VXRgLkrrokU/cXRoT52KqGP2rCLj2/svKJIIBzTmLEa8Zlezor4SnBwJsLLCXk
DsQv7S5cgDEHvGJYEDWFD8P18XpQalTrAV5/B/v2LhOBqc1mMJCuNNJf+s85DYTk
BfxsRgLHexPCUYCnGWGE7XwYVqRZKZ9oDALHjDdGWOD1kDNNyBhRdUdNgvzDGZck
/yYAp8JphS0Eb94A+tZmGA6Fu6Ag/DSfvN3PH+XM2gKxRKetSSx7XuqLreORI5N2
TgcbFN7BkOYYcO68srSuJoeACGzr/Iwt2rCF8du9tATwc7AQ2wiaQ2z1xGD/KGlH
ivZdhDfr5V+bunEfLo2lgT0x+siRm8m++ZDHY1jlnwS7L0XFsmZARaxYgNcuC8tg
dA5eqTAurfXX1TGDJ2gDr3JS5pyHN1kHl8jT08HIPdb6KYZVFMnyA1KHhQyM8HfX
vsbql8eerIlc4pOXe54R4icbUE3DE/bNCuXS37/UrUNYv2MZJt0XJYDo36lmnvoW
bgMQrQ6DIYV83JjzWkN8c45cQUPfCcqkNHYxPmYjJbc//PJbEfJAsaZZMJlZUyR2
CZI6HCKp/qrbfBA2YpiD4KfnKDD3i/kDbG9M3pQb67I2CmZsWPVQQNYnpZW3gus+
fuJ6I6RfJXUA7YAMecA0qBAk84R+Jfz6/Z1MpiwwTKhu5kO+2mqFXj++mQbQdrbV
/2aI5Fxrhz/+MX+H6jOjbfwfh/FwMOcGKREXRYZJl5xzrSRwKPPJojFyvbG+j9Ty
m/fWzFGPy9PWmqx6x4W+NhC8UOfm8GCj1yIoOxdKnA6aw6YbP3JYKN+ZzAKTwU2I
D8aVW2IvLr0bZzwek2oVcCOTwi4bHkmN7O7DVu6LLkfQjIZzENBA8R1CgIJj9hBZ
H7JS78dyq9++Yixvs4jNp/OLW7QJBWPDqTBoqR37iAQKKd+AKDZw86XNrBejswrH
eh197RKqvS7n2c0kRUsyifwSA33+q270uwd7qENfXz/vLuSUbX9qNMib+klK0k0R
f57cfEFrfb5k98rFtPYMpFJOsApxRc/1JeUAfK1bYQnvcCDwXYaB9mjoDb1Ud9y2
VntYEMVpyknRUwSCy4pOu6AeA1kw0nRdgeTRC37hTHvNB6PkI/Gg6rlaOwaw7oXM
vOf4SWYNzFeET4mvCCPaLWqpFlIqToYpPqoUtxXsJVTDAGKwm0npI+g7PFUFOUUs
MhIBrgX9xbUrsBfDQRtvfZGplx8O3bG6VFYxotZBc71E+cpzCdZ57dNdAZlEor/z
RPYyalb+Srs/6RQg3yD5SOlUV9fq9tFuxS2smOldrNmfqXyH8Sdc7vOrijfnxtHT
XTFJ4TNKf8CwqKPpISIlyg==
`pragma protect end_protected
