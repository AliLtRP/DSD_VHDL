library verilog;
use verilog.vl_types.all;
entity one_vlg_check_tst is
    port(
        b0              : in     vl_logic;
        b1              : in     vl_logic;
        b2              : in     vl_logic;
        b3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end one_vlg_check_tst;
