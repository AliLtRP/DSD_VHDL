// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:19 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ll3AkO/919pJDZqn6tjq5jBNfQR2N4j+u8Vl0pSwcvluXJdlXXOTZL6aRapditOE
LacMIW/M8wRTZ/ST9d7r36SlsPKvspLUaQwI0BO6DGDdRqW/qAYkyA167i+ynf+h
OCVEGMplwk1dMi7VCMPQ3uNGwppI0lU2UQyj0GNw9G4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 47968)
GYGk4CD3MbjF6qyTz4ClEhObKnvT7559+aIUUF2z7rLFigc0XXFWsdYC5ZxVzCbO
IjMMD+5KUMf1KlygTYnpuQd7NeFXUr7w4ri/3x3GqJsq9anb6ZBPuMT2lft0eEDA
Cji3XMN5Bzb+/C7iDZpK4PEDCrS2Z3p/+OJUbPgg94hmcFbJVaVqmW9yPr1EwvGM
CNe9WZvF6igy3/1Uw9aTOfViQ06iOZyRWnX0r3go7H0R3x0moEP/Ln0DeMx6V1kB
zFsM0CrwlFhx+a78X7hIqhwMr89eulJ/8w4ueN7WVC/frldkL9iRy2fvvRT9ERDd
IcUyM6LK6BzPXyGarmpQbmpTHwOoqHUrR2ILeoDDBtVRvIRCE2zK+5mCqoYRcqw7
EWYLsd2iq6wmQ3yfEbknWnJOnzXH9DU+r4h+XY8MxgMcTBu8nwWuoUdIElm+jn2M
OcIbAxp+d9K/MYrZZFGuKkTxE5e5czkoVtR9xCzAYTs1rA7xP9JWGs8uIa9h9YnJ
bzSxo+s8d1Laz+rNfUkaQdwoSH95Y1uxE+utC03LE18fbpZu/AbB9Gjfe5ui4j9b
AOc4fjHuHHjw66JKbXt0+czhmJ4yZcc/cUims3+7YhibJiER2hw6qJGQCLWorfUq
cb1xi3fJoGlupB5az55fEiR8/fl74mH+6N0fsVgQ2dlltIXPHTWmhzqAPFk5r9pu
Zkz6WhEpJT+jsMwyhGeP6V7JWEHN56pPFxVo8NYrhBjnglPcap8VLkhBfwhvLhsN
yVhCKINIKD/ZFbjsQvVkA2akeKIxIP8tqqOq4R+EHIyovJlotNrrDyuOKI61vORD
vl/w28SGQVPZnOoLQgmswqW38BtFD+WoJ5D+f1Rn3gmxLPGpG2zNMsQmLPxeflti
752dusjepbZrmaS7C2PzYiRNNPbycl6yrL2g0G3xx0+dNhVJ7DO1+5xrMiHKlZ1y
7MY5SIaYTaUyIsUZYME7zvaWzx35b6QYvdreU52GxUD6QwsmhPQKlr7ylkrEnJwC
nWApBWEG19jOTAqlwHeLJcAzYGYGlRJ13gfZR9tdjR6MA+psMMtUA1teVSfzT2Yz
8+HEp1HoROUFrc2eWhWKP3bl4cTCO+Pm75CI/eH5bXOf+p6TR7lhfEL4tdKdTJIL
CGjQ03RawduMRGVdmZ1jIhG7F724qELJgQwcH1RFxBCE1ZPf+HAs1HqGiCJoYMQL
gH9NOtxv4CpHuyg68VIOsypUPHXd5Q5xomZ+go0hr97Bnwxli7wXj7zgAtydTvjf
pMzgjjaOHAKi+4Cxhonqyy+8/O25lgHxL/DEudeC0wETMNXhRbMPcPB4uGQOzOCU
MnQceB0Nao2YyKuJKxbiERABmlgahzhx1XAZQJMlD2GM9U79ZYbFDMixf72H0XWB
A5TAH2j5EHov4FHsloWfKhRFtjyxjzVewlYNeycRjOw2vnUxYrdKa4qT6BSCKwMa
q5lVgE+X+/kID+3uj8dSKlFpO0dRnZL9JlYwhiWZnlHhS4OpiS8ImvSEqiua14zl
kvgd1jJisgO+9Krconu1sGNrlWMUfRebITNx5gx6PJEHu4RPyCWhplsvMvhazi68
DOC93+2BpoJYr6bNqhy2l0Sl9R70C81HvZGsm6RotwYPnTY8ee/fag++7FMq5Il2
DUfMvxcwmVpV4a87Bu26Fc/Ee7ORwyyRTAj97t8sWMxWN+sRRni9yVhtw/yp4g5Q
UO3VdMZo22rV2wP39Ddvi98eqslpF2WGof300G78B5fkj8JGIfW+W1hx47gfjA51
DdDjSDFm+N49a9BRNxo+RGIpZJ8eMJDJM0mb2//6NA8JlGsEk9M3iDHrk5phWaJn
VwVgFx9LZkpwqybUAIx1LSmiezkn8321PXI9I1zIn4fRooen39tJVvqsR7uPcBNO
NCglLKS283Nhz0ZtVQfpPmWHJ5fUwcrONYUHJJrmoH6XsufWdBJI86uAqJczAeLd
UeNVwSmcD7uyUM9x5c8nMN7ymgS4zyw9naGRPEAkSQ01jsX/9SYouOuqW2swBFTR
OfO9SzDOgAA6Zzvi1saOhflW6JXdl8Kp3V1GkwhevQ/L0do5/8Lkjn6lZvGomFbx
Ms5rrI7yHFu8DC5bWZy+G77vk5FBIzu4UGDQUDoqukrQQ4PCqmWfCpb5U65a4Cwc
JN8YCa/8brDcpCEkV7HItWlRWUzhNG0GlY6Ol438WgO0QegO3AqQog1uZ5/J95nG
ws6K5mmVVIFVa4yVys9rG4CW17JzQO+UTlLxxAS35nefYkKNu7JwwxcxzdP0Lr5E
yaf/VeHm1ERD+Izl9dbD8etQBeWKWBCvZpE61cxpFQgSZGgsOsXoWmOIEi5KU6P2
++k4yjDHpEfQHbe8lNG7rfQj5S97Wzj8Jo2Dnu4f/Y3l4QWq60oWfBmJIhc0M4dc
MyjUZl5QbXv1VlGZI05GsL3FkCqXOOL85J9k5yIYHxPcgKZ1TvJyG5mJeETgMbBk
65wswChWK8KCGKQcnGorgZ36HT66ENA55qZD0nyLkY+rNn94YDsQWluZLocI0YeA
icmxJGm+AGyNypPjRi7fPptl9m9Yq40JPbweNJv/86pJ1u2VQR9+8U+BAXv3Sf75
FqxSQJ3RH/eP+YoeJs9yUginFDEnK2ItIkvOiWz/xOt8jP0bhD8dlZWHM0464WIC
HN37PPh0P9hzU88pLGi542TkrPP3FR4qlZNc26to5ea9NPCqCjDG7OVBRBiY8KT9
xlrnAwj3j0rmq+0UpE/8u70KagKH7ZQgdiMjSjVcX7aksUB4SSmna6NL93a3MyLp
5DXKMTVCrH8polBlBn49iDpN59Bv0wSyqh3fe7DA7H5F7Pf4XvtmymY+vmQasKru
uDpuwv/DojyG+aLGef2/FXTkNY/RYRzk3Jdi+K0xGmsxgANtmLu3qwJufh4NNASY
HTWnwIZfBMUJ+kACiy3vRmWRd9gAxbyJKk52nRz+ZIqq9rjCXz+0KWX1SmhBJ4+k
Ek6+OBBBeFDE4D6KdxdnuoX03BP7cjXUTp68nbkbFBiQ7QMVh33K6K2xBl7oZVfy
m1xU9MqbEsugZDguT5dIg4A2A0An9ANy8f3MoeuswVXsxL0tlTMhrIrBLXJ3pXux
DQeI/4WIz95Z2ky07JC4GDUiq2k/rWDpMHVVClpWaavaSCdvMY02VegcmvdSw7YM
kbZE2e0S7LUHH+JXAnkJB8NWKehdupxIfzgq9qGSL+1BsvWGlixycmpwS1eeR0Tr
XLZqbIPb2nQAFAhhcm71e4yv1Z7nb2vnV4Py3AxaJGE6Thp/9Ju9ypdihOkbh1wN
F3BJxaTtfguSSfYYSHB7cm6lTqvTkOx1QQxFw/cnOIqRemBWhzmUplQo3LkBoMcF
u/W74DUdRcVHzFnJ3KCleTjSuBXfLNhgveWgEIPynQX61NpF4c10cWKIgymVKfjK
DYCvkpqBJ04o9zzhxmt9y8bvy4w6TUCNAbZAlx0NcnrvglP06gTQvdhhkCfCjl28
t6t/gQb0+pY04d1mM7RayGbtPxRVnXrfCYxjhqH/9R2E16S7AXD8H5shAFGmRZNj
cZ3jSP2z8OExZPqKZ3IcP4+yAd/Oz+Z7BmvgfCYMqhrgSOvcniI8iJWL3KCyAakS
O0YxwS15a7HuiG8Bsc7qhjOgbrRvFJG5qIF1XXAwnNTr7dWt8kiMRifTPstbnP9a
A403jkNksmKFg+/zp+JDuoe3vtEUSCQ5DC0WN4SCUR9tpVy6YrHbVMx0oOcaCYdy
lA5a7HQrY3V+VJC0zQRDw4GNuSYs640qVkPovkBeOd2PM3GbRlCrNzFGwhiHOWwo
Q/+AeEUfhjeXhWLnef6mCkUjMkm6tnEmYEwFF9nKrG4W/VbYp8C58ER8DP+FknRP
RfsJ64lPv3vKF3hOQMUDgDqaI9VeX+qsXuMI7ZLAQY6Mbtl1cvUiWLfkBS6z7pfK
RLd1M8auOeyHwxvr9l92NU6StmLnR7TVgp330WMJQIeExoRadLOhhIlqgfQDa8ZE
Uf8MY8TqJ03zX+LjaZOOD3rwTsOVJ4YcVdHegJxElqD+aA8XbgifzmkrewiEJORh
hdxcRx+iMhzMe9Qn+qrxtjwW/sTglwo77qlsqAneHaN1QwnKlMzW/LSWCaxzZel4
lJghpzuAoZvwKNAR7LDFcTrNkKwsX5YKZWOQKXUoOM1Cv37ithRo9YjTbLp2JKi+
vmXwzTa86AWdmiqPpFqjb6WbfvjanqIWL08wP6Fc3wUp6m/3kehp+E+ELJFhs2OK
c8tnmMSRQjwivZ0cBDV5lo6DhHU6fNgTCxpAoDdicWyehetBxOAi+W3OzTTvwIIC
zaYVNDEVEUrx0nJ6YTV0ufBa4cg/WDehOGLud9n1APH3QV9iS0SUrUV8E0OlW2aD
s8hVTqHFjWw7n4E1sfaGQbSY7ajlolqRtrr4k7pinzwtPiL7HzZHXM/uPre+8cYr
jztHrufSXP4vSsf8k4Jq/bgHmYK4add8TU49Ux2wK6iC0MTJrul6zozXPt6nXZsY
3nIZ5CONbGPJyoQPu/FYIUPRkYX3O3/KxADbu6xm8rplfLPjzxMnClRpsN7S+9n2
VTZj1YbOHspAx8EuchpaoK2IiqRB2EGbg0NbBYV+cVZ71N0/qgcANqeP2rWnhTZc
6irjAvQm0SjdBKRLKkCPZx7bVg3s87VpxjoDNp+2vFYsKAfzNlIYB88f9XfOiupB
ckfup6bE+tjIBcun8YjVBuRnF/WhZyAMzbj+cWslK7bjfnzH3Kz21X2/xHCXXmn1
Uqh3cLdN01ZwsY4Rhpuw4Uj9iSCfGnczZaYuuWaJ215MKoBLDZR1dxonPLXFkWvI
zc8G/h5AgVNg2dVRU0T1xdo+JZYJsyVxP1Sx6IRqVERArS+HXg7EFtWuZ7yYDuEQ
e7rokT/PNV+mX50wTWDQ8xSNL9VBS2JfN9UImZgcgTMjwS4Dc9ByvVwdUF7tSGvy
PYwk+BMzjQMfFH+Ry+MLQDGu7vA0vuscqfVgt+9jXVN17ohZm4Vz+Kcyf7zKB0yv
fmpn5qZa0WGftkNFLe/ScbAPJ0+htCXSBoH4bndjECpTPGSJJ5UEyOQaJrohnTjT
xCstBWhhG3U6b5ZVx7VW6yacXUrd2CKizOkiGxvochHd0N7T307yAHpTCBrcCl0+
tLNiKhJsQYf0vaH3YDXlxQ++JopICyckh5N56d8yQTTF/P+ABEZyz4J3nIhvz2yL
2zKGVDqpL/V26hsyNXXL8A608HmKGsaGXS8BJWQLuGn+39GKgI/hMO0Qw5jtVmu3
GEojNQX+rt5snTFD5qOvsJedBzWLRgtXLB3tRbIjMRiT+TRMj3WlC56Ylrk4n2Zd
WHgd8MColUzZ+urRYclu6fO/0K2IzkPosXFB9bovk0p8rFNFNvEA4ZQA3/ayKMO1
E2C4E3lG0j6kCKfG/pYWZo49tJpVjolrFOWc3nDnB/mfvLFAPORunhRED1IsP6uG
Op8zBhC9ctYrqRX7oDiY/34pqrLY6ndjYkGS4JLeBOuG289T64oaODaX0O6swUt5
dsYZEQwhEDNhy+mUsNMKYGhVSElszsxF2J98z3JMjyL0dqvcq3+vEvdtRiUKEl1x
iYgGS1pz4+NV2LdhI4H3ITaJfqbg6rsTuM8snjPBIeCjlAQ3nLcvl//5hFbYmbqa
P/qj89fkR8cMdii0WJgyDZ4aTcpx25x7gZ3KiajLATR6rJBcipZYseKEXQoBgNor
OiQHK7OiG+KHQGfJnjmw1y8h5u6nnjjBEf6V+imwqsaHClbC1qZgFqQcT1rD3Ygz
/pubgvFuHSz4XUr8Cmkw68gJAGW/AYmJg8bHUZA7EBrjoZ/E4yg4y4rYf4d41shW
3/S7ZysIh4JNo2gyo74jsJIbKbfGjqkfxb33f2FTEwfv22WmY5OqamTv3/+Hfbq7
p1I3KEnV+E/F3oaUIM20pJiIb/Lg5eqlVWKZKNj/ekDyoWY67f3nyC7qJXMVtjXy
4CxyQjno8Bj+Rq1cNKGCm0mTX3Zyl4XOQi/OPsS0HBaBd+DZQryNanBtm6PhlZsW
MUSFcqK5xut9t+3znwaQIskHV3N2J5SFKH/Gb3nZoG2qWRZ5X6/zswZWSPUj03ER
nJMRdghd46whDHTHbQFXuClmWvh8f9vriaQoDd34toRb9aDbcuqxR62pJktp7V9s
Aat395s7E8wH45nUSKxk1e/ahCmLo3dwru9SONI2XmfNdrBNfD15DPIZ+98L7aRh
EjtfHNLNTwqLH9Tb44sNmS9Id+eSVutee6jInhv5DseUxYRSDJgVsutM54HM0d/4
Qwx38iAcIJJaPel2SVf5oh+cLJccKl61lGv4bX/aW5KyAzJbabysV3swojItJ9dD
3GCS24HPuUQwyP4GSRSJy0Dy1s7M1MwSbCuWa9e0HtLzFYLZHzn0YBrWMIYug8Wi
bYLNv9XGjXZJRApAQvaV52DFexdd7Z2zXWmI56+ezNSC7Bt2CZV8V/A6DRlFpnFH
RFyW1xkQi4ejuI53hpcyPwri8FQMR46WQxi7ufyip61hKh7SKvdiYveAv1n1UQrX
xTC7ays0r9p6ePZEnRZSvhihdKy13ao2J05FxfTSUYLjCYskIfWw3mGZ+je/KYZ8
338Q4obdiuZhZBXGmS89yUH1Y4mNZbo0jPkcCFPbu5J8XyuN3+dc5qy+h+blTY3c
p+y5XCy95Fcr7BDlb4VoRD+/OnJjROnF789dE0hG3lANQv7/xHs1CNFY6Avz5EgN
jq8iXTmQkFmgrond9+2QK7bDzznL1Snzvp5f4QxzSpALocEMuHackl+wKGAyek4I
nQGcIKQvTCG0ICWEg6whY4W68dGk4y6km0Feo1o2/JKqNpfwfeXYV3aN2eGaQ4JD
s7ISq3H9ga+QRGi7JWeJJ/YzkJJD730xvoNF80Bjldw5bdVzI6mjZ0TguUT8tw79
Q5R8s1VapL3ypJeoJs7nLUuD0SNsD2FGs/S8Vc5rGTLANmD/OUR04fEFNQUZq5bd
x/I6tlmYac8Zn4LOv1NdzGstUEQ9GD2Cono1gUUT3P0gIpyQlb3EEE/mBwlp0Fs8
4wyeSpbXsFzg84xVPjrbr8tAQAInF8ZVDPFnN57RZB1VHJ4xi42+EkVubL6yX+vA
k2s1XgIje/ukc4PA23sQ1V4MG0mIySfQMj0wzr1iLBDqTk4AorarrR+Qa/qmg2qJ
NH1vLeLhO07Cc6rl0vnRlla2xrwOryb4bOL8Vh0INd+nQ/r2jS2Ohk3pliJJpihF
jUSRcW5f8UrsamCZ9YOWHN8KChK2KbJFmjDCnxeiP/SDhfe4sefqCIVhu/nLe+lx
Xc18KRm0GWQqbqPMEhYFDTy4DsU3apvF+l3XoJ8LYJFgc7+QY7Zt6e6IiXi0Z64h
YjwZ8Y5UHMTdwbhf/RjH/Q6Eb/a/h1UnbkXKu4sPsbKKja84GiTrCJOccGZA8HnC
IB2Nwjvc/3Wydl72aQH05IPH2KSHonVCsSDpviyKtskhuYvCo6V9/q1fMaBsFUWK
OSwbM7P943KnGK7TyTM5WX7gWqlNPIUDWv0WjgizhQZKl8PIzuY5ccXpW7x4IURZ
dOSrtgkzR93xbsF7OVyWZyYOTCUtXwkYjprx4Yp4Q2/mvdOkg9q6El6/8XE0lwBp
BeO/6U1qqUHuMTrtmGgHv1D6+TQft94XSfz4Bj58RQHIIsOFXoTwmt3+Sh3SAUgH
vNlEcgVby4sQcgx5UGsexc3HGssmRdUdEAvGeTCnNLvDoSml/IWGf/Ck22UbX02B
7i09ysyomq9R6sMf2t4qhUGCyHhscAGYl4NtoNpMPTZkugMHv489M0G0b95GMJNj
cUswiTmzhHxa3mwdW2Y/wQqeaerOOEQZN1y/BSZltNqvk1DGdPcxnyvmkP3kSwWE
SqCtxTLdSe98a8HPwVsOS8QyEZWxcVry/fCXal1alk15uYx646hASO8L73whcucu
Vywf8EhPIrnyligyPhuTMNIv2NShec8sfScydEeMxXVOQJ7rH5MPx3hbiOcinR7U
+4jd0UlxTm5ITvCFTl3kcNv/LXE2SujCZDotWeTu8akcx8159y/q0LZxvGLDFWL+
8pz1S4Qxu+soqrxFwgfCuPpUXb+RWKbuDp6yR2EIK/p/uaR6Lr3cc1QjSv0VEDzK
UJg1Rnc58g4WhppYKltO8UTY9IUPQ7PXONSzzFJX1WTnc9mlvX+X8xI+RMvZ7RmH
lW51PVj9R5zDXtscJ4axEvL1Sz+y8Mho8rXLof90lrWTZRi2Fk51XoahggOiZKBF
LKa3p9vCb8fx9BgsUFkdWKaFs5LoXbMJdxY7SvrmeJ895LNRdKN6X0+n3PFeCDmt
If3q53fa5RLA7gTmGp3KYGmNMzhePXYqhvsYW2mA7EsoqsJB3X6N9S9LSVdRwGoh
drH26iTegQ3a83ymwoUDx6Aiva70vWZyBJEnv07jmCMeekerVPCfEtJTcPeq2nK1
E3AvuLjgcrpobOyRug28HH0pIWq/lG1KyUxf3RSwAMHRVLd/3mDYmcBVsTK4KRJC
vEDqraH4QmnHHewD6L621LEpeRaxQfnpf6X6vZKndbIZZz/OBn+FElguHu/1aRPE
/ngSsyvZnA+eFRGESWVzWezLNY19O4VoHHrLzOgupr/UGKjWRYylJkeJBT9zIHfm
tKV9kB4skcEMH/rEMNhowo0AhvevJA0scmSu9YNB6d5aI5WsT24C5BfYRX+FEp6V
NfHb1/3HWVqHbAEGw5bINlBDilVKupTTfaFTs8JL7v4zvDJwubBoAwvdm63GJBF3
AQeX6pw+Z033Ovvifx/EJsR7ps2mb48DgwYqCMT1Z1p16pcKB6fnD5gqUTTdX3n9
mRI7ddsvefUyr4rujKDbNhR+4U8MBtLNAJalEeAdDGWIHzPX5rJVRM8AQsjZVG3T
rUrxr1yDQ3/wBDS6DXIXQrgHJZSDuVQdrVWN5kfAZqX1FOP0j938JoWAMnIcl94y
ILZY5WHj4mTJikZOagGRxakR21Qp7bFlFc13QyljIsGNp4A1VDrUCILd8bELREKW
uKwSL5zVNf1dutY1fvKIsxvtSaaXl5BKhe21LrdBecsgVHeiaDVJur5AQ5oTccJ4
K2L53MLPGKcV78/BSTntilN3WdWnLvJs1IvADQUW2FK1v51Z6+yi1ftiu173YOZe
OiE3BXNfaGvzWdsTq+olGUTFAyHR93E427IDGbU9V4rHQU0lKQ+G4xO7+78vLShK
2oTVq+/bsHXHn5+Vu8q6iJDq5h5gyj6jFC3R9qHEf88vkx3TcCEm38RH4cpz/ZV/
Tdf1uUKrlcJqQx1Iwg1cXptcp2CmevAHu9+yqSR/QZpy495+SG4JPGX2c8kLC5oR
M9gQRvr7Fn1dXS6pr3rUyrnIE2DpaLp/wQTvoLIrQd/KyDXYlSqqP7yxt5vr19Dl
UIiPVEAgu5/sIp1omVUFZbVA0VKZ2aaxz48PkAL0DGqquTbMqxZGeDjZo2JlvRkv
LFDZBttTfnmRUJjmbdI/TN7FYYrBMB4FL3TAWlqco9uyNsjehynljVB2qDblt2fy
5Bt+Jadgh9AUnoNyYSnmf4lwAwUSYrNltaM3677yUmi3h8GpL7PV82SAgKzEs/5V
H09Upy6xOofHG0Ck0FLTnwhqELIMfTgNGFW8cR2IkBpkbaiMz/MehGfrxv46xD2E
BSRzxCQ82q9C4B2DBxrTtYCk/DiHNqIPAg+dnhOSMkPrL66Hyj7C9uGcFBXNbF9v
MzL7C/YnD4Q8eS3hZq1fEUNZn1FtSNKJm+EuIOv0G7yNXcevXv8anApQs00AVrMe
90kbqBA0G2XxK8tsSfh2YIeVKlCAMbrVbObEtjg8edGyAblomfYqfxnFkbkahvpi
noJUEq6LWio3yubIsuUJYThD6ecwkAafLRMypd4Wh8fdfNDbI6nRJ2X5pfR3HxO4
8qfJNAzyNA8NeIQQ0G+VfxzzdlEzHteVD5JCPs712T3HJNFbaPHQTiHzSPoO0hBR
XdvlkeUllTsx3JwONG7W41lj09H3FYcNnxlqZFm90uv2WYB6D4Jf9vgWNYp3Mi2d
dycnL+hOYTzk7YiWURzsLavg6s8twioeW/GtU7aSOY6mLHPw9/VHAA1vb4ruhSwt
tuUjR0QiMfrjnikNkT+GzIS6VzCPIoQuXoOklXW4lO7vGO/fs4Rp1AjY26PTIKsb
pgeavKs2U2Qt879iib2y40HEnnm01dfLjITGG2f8PRoZK7j5tatvW7H4Bd2t3T+e
Z+Qln4iIv8JFZpR69FbM0edRdWzDbXIU5yd6WiNxn95h6wlyonZ1L7N/SXxzJYH9
WxJmsVpiyIUKaoZsYvmoWTaND50kvyGQhxD5GQPZssFNJ8uSRBFq0zoqg1WpAAKh
htGRQulqZ5E2YrEL0xjM0Ofyyfr3bR8rAERD4eYo9LUaR5SaEFPIOuKgPD2c9VL2
pl/Ti9W5IgDgUTympg7xXavK4S115/hddbDjGdm8D48v2J1i0WZvJobaXy5SxXbD
i5c3l9Ckk/WBgqkjtMPWST249p7u8h9HqeXqfUgwSeMkA/EUeIZdMSDyjAJvCHpG
/r1XFByllObUP3X7kuECkvkrcFvWkNU5IMEAuchFyIVkz1TZFiTkw085gJx/iZL6
/2Hd7Dth367cuundSgfAom48fuajZaZQpP8bF8kHKMNgeSArrj8AbRpnjRg3shGX
fAptN2lYz3e29kh+auVYryxR9zIS0FaH+OzMMQu3x25V/fFFJ51yg1sZJRYezJAs
RDvbRRvAK9LFNVrlDrRwDwJsCqZ6Rw/DWmE2K2EHytkBcNGxVwVzr5H8DZ9q16w4
WeBgGw2mzxhN+LKEPt82dYjUKz3JgiAAnFkjh0wMEOsly6NHZtrTo9VmAp06T2pa
MQ7Uto0OPDf1YwFpoy0s3yE7ANtuw9AD3nEHCYopGY4BOPTBEh3k5laX2TtXI/Bn
KwZcqVDO+qdse/Wi7c2m3+Vqql24i2U2DDi6rIv2FDPu5ZpBvL3QAjmWJI8n4JqH
cS/Qx8PBn6XcTHMiYXeMW+cKFgItj39eZ5A1h8E8ZDGRaoD889XVEFXZjxGc9ctt
Wb/hPeVbkodkDAiPKoJr8RdjMp/80EQNFbeYxS0/FD8iWWkZxXvNP2nO097woiBj
+HHrcf1uAbwvGulqFVsT6MBLt7IyIZGvaVfIaW64oo+M+yfUvsVXAqDatPgIODEs
BIMGQ3FeidB7oncq00ZsMtwuPWTHAm5+t9Hkol+9M4Z2d4r9QgQnN4gsyl/RrxzG
TZOXdZkZM+EW8qVc5ywRunYNPHEfZ9r8DfVOakoW7WZ9Pe3chmQM2+dZsgIIHLAC
2VnBJ+/ubyqQgOEpgLCDjLz4309rgS7P/sui1Hn1Oz6Kqx6zYZNvomznvEkAcx3W
IdPFTztk8E4/BLnxjAebPYJrq9J3M9VQnOU6MmTjchd1xXu+wFYpjvij4SM3EXak
NT+KsuhyyvuFa30qsP2zCxJQ+uUDicdMMAQ1skQGpeyjNPncZ5d1Hw+eF+8kLuR9
BWwWEWmM4txvSawm7unA9sdIpbHXRPtx2ymKKCbnu5fxb4GUUBEnRZeTcav3yrpf
vEbLc1XWw+amVyLjRjnnojTlDJ0qYl/seVvqbHUl+VLZYUx5da78cTCvUGV9hxdV
wO7bHsd7DW/7JbKv/wLwKbuI2WKfwZKs0BD8yLj63IRG9g78VVr9YMBMOW7bkvTp
bpODZKI2tS1EBqkqZczHFdqkdTU5oDmuTRu2Ak6zdRYTNCtFAVLN3Xdq8ti1NmiJ
n5qk7bgfUnoSTTUr5bbADXlPO+ow0v34gWqhuLG2e2DTA1UCYesF8S4mf+knjFXX
AVN9uoPgTfwZRrSNuxrE/PZiYqlfIIAzyi+Rk0sbMJbdzjvkH2bZWlopZZKkCXAP
KO1nlCg0bxzVMm6Ag80ZM0a3ln6VXovDM9eaxOl/ghroFm/j6YSZOp5B5se4zPXL
3+6mM3lnMYt4eT3dkciLtNU+ek6HJBDuekqVYSMNCLRNMQkaD5ZCG/CzFKC3gFZL
AokUMpxxQ8VJJoXaE9/hinkygb4qYHz6MiSR94xHb7dxNhr5MeyKL30XgklRHhX2
mZpFEUz3NlZ1BN/1i9T3DQ/wxzZH3E/zRubzakTuTo3uN2wHsNgRTjd1MWhySo1S
0lRRjNVhROI/C0ST11dAOj/uji+HtdfsTY7sPce4i6uxUsflh/MPcLox11NQk/UD
E9E5kTkWN4+hWJn+JGsbBiNDWR7bhbs4itphILOpMFGYWZQWYeAljwHFLbAR7jgu
W1gv204+yUUZAjGu2H9GAn5bcnKSHDxFn1ABWbj+kzG0dprf0RdalXMh001CCsS3
PqcWU3zcCmu+5rp2bjDayHGeof52q2zjkW59+71qbC4ukibPBAco4oTnkk5YbqBW
kmbYKhcLtsOVrBX5cbdf/KZwhh/UwwPJKQzFzsVxyfekSJVbGSuhOY5IlhzHkKZV
ZoErwtL64Q1yvmyUSMnJ1Twux7QOz2CRGwHA6uzvZA+BGbCEpaLoGYhAO6DXtsQy
EuNH6euwST0Yx1JJF2DKnY0stXpHtFAiR2KRIhwW/+hmsMpY8rYac4hNBy3G2nT9
/aA7O2vqjnAJFpFvNcBuTExm+zCxhR9hkEzJFFikidPWGHe9l/eQB7IcawcV7Rgo
V0jV6xPIGteisKd2YrjE3EGAs4HMsVY8PcLNoKmZPMbpbKTcKICyqfoXh/Yd4P9N
TD6gtyD+QO2NcNEAOrIkx46oVj8RyZcjADB+fAcYV9Q3uadF2SQG5zFdERJxnCgB
KxzsHtPOfsQTb1qgcyxgjSGwV1ecgeKX0+zPraphtdv6k4ctfh7G0C8ugF38JD/+
H2dBnhA8L2s6q8yZL4jspWckYzidOTTaCBaEUtCSrctEJqd6mhcCW0ipjjxlOxck
rn02vzQRD2nYDURo2P4B0NmVuG0FIrWtAWrj3D6i1u8OfPeRhQBb+PaYM9s9b62w
hvIodxWpA6mgT8v3waDk+zPTlh90ye1jF3AAJISrt4SxjPyGrgEFfl2wS4SP8FCR
BIJ2VTBn2TX/7tzmQksjd2pnTgC32vlfyE9bAqgaggbjkO0pW1rzyDIqEZwc1UcD
jYZfQXW/MX3NQN0YShrZRIwFhYdKZyMc6eurSkRTcAyGquVDgZlZYJx2LUoBQm10
RWC0IcX1mGbJ5eVO6T2z6UrDLoopgPtWph+JH3G7ScpFGHULMuKp09zIVi9lJ4vo
N1RxJl9PbhyYf8+qtkUMpAu43Yzivo0/FHi97rYn2fY+QO0TR7I1HH0zysZXzTtz
dXgoA1Crv9GLGOFkLRmOln2lJNWLf068RoPG4sJtaH+AuJWCR3BT8qxG6IPLJQ7B
mUTxKbRIU2YXqnWf+njm7J4rYR6brKrQEZOgjei/Ok1IBbe5voVKZSrg6ukXhWOH
fNUAHKfBW0Xj1P8cQRDP6wL+bS1FSQbEFumIOzUb7dbCf/md1xBHgdaQLPUjWIrM
Wm4j4S0j4n2ksWdJqmHoV7rbyOtLZKCPqaOdy7ddqgPF5cNBbtk2Ygb6g/6LjaBW
ydhky8lOWWTPDWvmqfjVf5Rb7OqBSKP2Cz+iQ3xUCOqMigBuz0lu/8fP9wWXr4Pc
h9lpdVPhcxKp1RSV/ahY4pU0eQgNLW8PV4Zs1qRzuLrTb1YQJxE8mRAyZZmDd5Fv
UiNa8ZZjeRySJubC8I+eOKQiKRS/jLqvZ7Ye6BWKS6sRuXhQg5hGJWdtfVasGFRG
G0ly4awLpSrLozKeyKZ7qfcpBO/ibzreTq/tZOLop+RHGF5IRp5nRRyHCCTOqL/a
uk7EpN7Ujsi3WEsoSMq+aljCXJu00LVtQu4fOxP2OJ2HVV8FfmjlLVNJYwp/wQJE
07Ur6xQmUL3s3vEPYKb1PTJx64tuD273ULGYVx4qPwBy3v6ibuscikEQqAwGq0a4
p/wgIQVlVqZoiEzKfuibYEMT2OzCW+vZOFzPN+hV5jIKvUfrsQJLxNj6rgrykfYb
oujsWR26LWxcwR8z824wzUxWdc8YlLG1u4CYYX7pZB5TwNs6StSP2Nm4LA3Ziq35
/RlOPxJboep++3v9071a1ccDGDJyLkgbJbxHI5gUnPsQkgapXAbpy/hQx25bvjon
CDdBbST/RnT/dffRctEj59ChllJJPXFXp3AtUtF8h8cmm2oNxKi6pLyDQhevwcoO
8wXEiQEgNhoq3VPDmcyhG1HcPXIkSvTOx5BVjm0+tsObzoOuMIZH7AmGShpSQfkV
lWfkIURgZ1xheTz+/M1HlVmMQEU697NX9erQAE02CDvD6dsyug3eBcDQcauiFhLg
Zi/0Dn3Y8jK+cBxoD0dM/0tJ8+lUMe828DTU++EDLqzVQblzeTmGDy3gtn+T6+58
WSnbRBXZ27CJAhwQ1/fVpHgCBUTJVANfQtLl25YtyURr7urjwwxYiLhODamtlW4E
jwrj8Rfrvj6LbAxzQ5RH4WrHG75XgdhS6Q0+7A9DQ93oGWZ4UV5IFb88KGkfW91i
qkwebTMh9JwnZxi8QiZwhm/jEY4wvfktuZuPXbR1rMXsk9hmaxRztnl4R/ClbKyv
S98r/dCNyiseKb+y/RczbXlG7+oMMXIAyKUrWzbjD+vUh4VHqWIPv9lBEvDMn+Rr
35b/so3wGln+px2ohc5/wMb39KcUQVPOkPeIgHbK/F/9w55NVUhQj8W6lLkQmgTX
VPp07BMSGx02c/v4siBDpyNoX4K8h7JGLfaqPZQWRnAnTmIbn0CGA19oT//deN6X
F/hHu6njUPLPbXt7wzP5uzyzCLEEd2uVr1BnuX2U8plnXOoadatsyM0iKsfhOwLU
MVBU8D0JCfns2Qz25lr1otM8mPojt7wpT3J1jFQl5OX+Lb5/oZCpgKnIbHKIINcY
vnILLoFbX0H86HTtZiozB+VLCgjZKTkGP+ijqejxVf52zjPLqe2vQAT8SLQwXNrh
fBm+9kQevsr7oii8Iem+/lE1gcPRQ8+WWuO5U5KrRhJqyKAisCkVRxnqMQBBJg1p
6obkVusCvioBbbpxHufhWtJpnWtcqF5oDPpu/9qx5wZU6/yGG1iyKoedQ182lCnG
4nXjPhwvktwvnt1uZnMfqp/T8sV+KjUUG1rEoA65Jq0+SeX1Ny73dNtbdj3iF0oL
/J6Rk7KtDrjXvE0jAFdHgzjxrhwWDNzSMaE83S4nM2j5AwIdoMWXP7ZT+bhnXb06
D8kMSeimlA/I4etfs30aH1Pjx7pvxSjMPI11o4zji3yxgEI8IpaKcGK8GNaY801Y
1t2qqW2GoQx3UGx8qh4URxoLs4cMicgRvK+S9Yr2eV2IbOeB30B5XrWv4Tn4LxcL
UqP8ojOJbLKlM1SbcNkb/u80L4UbDMekSJ4Td/Oa0KQDBfHPGpWaFgHZWYdYqipN
cTaVE9mPM9W9FqTO83rnQjP2ycXQtLoC6bsVrLQxUtfzOpRhMJemOh4S2juvS3xg
VsQvA1bOmVSlCj9Uv515ehxG+Izl/TwnYQg5hVAnrn2/yfjDG+6rQhC4/aNOM1jL
7wsn5TWAAaNp+TeJ6zXCiH8hZU9yk+BMLrSmy1NKKk66hTEuhciHBLbq93KUpXOU
YTB1ojDxKY1fhIDUDVoKDOZV0j8KNuYKmvxWCMkIaAPElWgsVT4lQkdBt8BflTQ+
uYaNbwpJb+udXBsPCVnOh4u2IloiRcR1+sohbSCjVKxJQDUaetvoAmNuECijv8tH
0NVUGBHh+ZiZFtRqvGbBb2EssJ7GhMC9ExToB9DzqHCqMe1ks/+WqoK6C9ff+kVR
qDFHyUocYY/yxYgfyVRr0yPyxFZu1oprp/1+Y62Wiy0a2p9DbLGpCL9XaDXN6ok5
qgsn3smUk8ZJSkpDBN/LlKWDDCzGAJD7xKgoo4fRyYKoNC3kXdBRLHkr27sgbLwT
nypxuOI+Mw+aQOukgIlDL++J1NOnjMuXQz2+8lIFziVUy9d3fCUoHN1NZu0r+9KB
K78MLRuWXep/eN9dr7Mxg/vEqmaUzupndSqBN+3MGTwZS6R2ZIeOQhTstPAAa8lK
QQyvbat1wZisyDDEezbe8UiaHnWDRK2xh3ASvcUuC24rNbKJ94Qnw0HCAk5WJ0PB
qX6NOJUhLKAA5jnA7j3Xh1YxMeFE0jtPu/7KOM4gP3eKlocKQWaa4nToVkLq575f
rggVK/3KmI46zxFhqv8mjWPFr650sErxCGsGRNRkd0xgEHbGTxq9Z9Rjbu974rXf
vlzM5lN4hmkX/i6gd44Yyx8SLcaRyvoaFAl2oM8WPtlGi+L3yI8Ce460feXzaaox
0Nunrxh0zScfZ5mcnFMhUd0tY0+Bf1O6ZeFvy5wjDjt4Ieqxa7EA/mpKp/w4wRQ3
lHBiEO4HnA+UhMI8RAcQkb45uvskzv9zb0jsEvkBEmlJslUvwbhVUHWnJrCMyGBi
53G/tO9xyVH4DiIAf5pauFaPy8JSIM30b5M95b2kmZBlZqn/Mvjpg9Cb1D9hzPlA
xFeaeLM/qZXOFXlm6KriO1SLdxnyVCp6z0rGBjIKLYdlV1YcVRofnWClrfG4+yL8
IIJIGvVX+SntG087PJdjLA1XuQe6iv2yPFJJtxUFOF2HwNbGB4J5LOgZC01C0zbZ
RnGizAbFUYnw4L7Io3aBEGA2fHY/oYgDOyFuCn0wAW9iETHLFxAHatVID/ETkfdl
O/6qlgvndb6bPnk8a6aSRXA/dc/v91OVfY/UnjcaiB71ERDfLCLpDRnUFeO5MBZF
fbcjf3X0LeL1bGwamlzsgxTQgE6iAWSMGTSHR4uhZpjDL2mUDmxVlDlS5Pict+Dn
4vBZCEj8P8oGJ/JYgNBbN9qWbCmMctx4BFrtKY+7e5+cI3J6ARCH8wAG6VCd9LWR
dmqbfVqz+ISMlsIZT29E14zMxnjR4Jyqo5PYv60rwFvpUZ4rd0YzCDBiuezEeDds
IDoPicjBQqO8DQSouxZN6Fy5WNitvKM9cgiMwW1zanUTT237qrKAIUT5Zu63z9K/
a2ZBjphuAi+Ka6t3JplPKp2e7e7UoLDPt7m2lOSDhuvT7YUikSR/sewOBXNvh6Ln
YGKPkoEV6YpP+0rBmt5yGlJd7RSN/v4tiIAXTgaaF2/3v+ptBxYHBuWjLmRQs0Z/
hF1/HkfslFaGKOt6I+z8JSBN/rV5xXlqF0oi7g7VsWoAluELhnr00dDx2QMkh63C
SrLSjP2TgWICQh+HJ+WwQZcgzh1MyBmccj6oVqDwhr5xB22yzCZOO2tzIO/u7hJ2
sE4wb+7r5iCNCaGu9IqHeOV8ePJq1DujXCZamxsPU7JGSYFg7xcXxKugH3SAIqsh
dnFO0sC1M3e4agdpEJUcGkgEZMWz+CTk6LED4TGuzQCrV5I3lGUEbr4GlXNMc/Tm
TZNeDJhdNc7QuJj32tQ0BA+DjtMBTUaKWlTB/YyfXV8AEp6aXmdlX1hHfCdj8suB
0jyVk6wvJtxWhE1HNndRtQcLgqXZ3FwmAcW9jb1X7bOqH3XPLeP8ygCzZsrsfrkk
VFB43XH9/Km6jUp2+IbZWIPVGlu+Y4kmDO1b1jX1RkbVCNJiU8/ekTxyF/XHzxo0
3uDBLqSZ1R2pyQVbcZ6jl4xkhB16PmspOexFXC487mKIX0/7ZJ7lMW1LgSzs6eud
2i3qABuu9qufb0EEKYNWkq8XqbSip+M0KJ9fARarUBpEMiKT2ElFnFPEptZ7zLK6
7W41jGTLfeXJhH/y1Ri9S29UbYwWZFyyIFYAziqpbafQ8ES/IPDpuKEG4PCFBNpE
bMOaMh8FCvoVzbdaaujn06/Rg8JxTtDCgUrEbogAUH7gWp14cUyeN+FkrmEtEZXS
XU1SUxKQHqwMNaGZmtRyh+i+7EvMAstiwZfATwAJxkdM5Qy+Cv45009ZQPwJEnDV
GRurjjCsqFWKPZduxsSpywSc0VXRzYi99DxKYwzm47qbV2+9Vc4PCePfRvBaCB0i
THSkr/XVU49ybS+FsKVoSe2R1H95cfx2pSV4OPvhis8pwJHL2DV174Qg6wodWyiu
Wue9yF+rdyp0dQlfm1ws6AhiaUbimt7jH8uZ+38cyZFHosy37weg1KFPB9pIe/3x
fGUIuCzcN9ZMc5t5trE2yDHsf5UgqeU5OaTqekMFgrDYolXZ8+8iTmqTfl7JDx4C
bz5uDFmz8c4YyeCXybBxv/Ay2XQYqlT0no+N26mC3dEU88naJZ1S7EFOo4gB7yEf
0j0NqBJZTy0brdwVyUQTrIldScj0mBt5XgRjhinq0WtJWBSbcciHeORjVrXoWwW9
Q9+wKxwQLDeWWxT1RrT2tnYCgY9WA1RgfNOpFAtw1dbIbZyaiKrcsAMei4AEw33R
+Em6wLfIuh+4iI0SekUQbzaWJQckxRnEpG4Bndi9pkeCB/XjVUgJRVz0WaPC7l3s
jxxZLQJ/Hu8FVPM6ZnQduKKu2IwYvvYdV8fy+UrBavuN+o8AZVSjOlH+Aq3YM7be
ElX55w8n4tLHYWjTVqZV+uhVGwEI+XF0pBUdU0itenII714IkTxM5CViMPqlg3SZ
n6eetkUYgF89tq/M0KEOile6saMoTVCJzs9AaCoXZmvSC7xzvnSHkbAOgAWKaW/A
t3PTw45WkRWXcdhbjSZ6gEp+FjvADBDyqLlZqEqZhaFNKMAfnlxQhsmUNI05hXH0
mr8DTQrOmR0mcZBQeFdwX8qbFChErChx/7FiKE/xcTmnuGJfqtzdztOsNj+PMgjd
D/BJsEjrSdEPn2aBaYcshUtSb2urdtnJrzRupHwrbxtCTDEVp9umWhxqtOdY48oD
tHdMx5XzRzxZn5Fdkb/JkTFFAkMLYqXddJm00R6KKK2ib1i+wAhjsj/kH3twE0/j
4hZuGBFpmDp49PPPGmUBpdYlWsClKxvX9AhKfddO9nQk48cyO2OyJ5+CPwa/Fdds
t0nM7xZILpKQUCUXAsDjYT/x/24+trrYSFUkpqLx2bqwb9ZStP4UqZ4SDvuYCkSI
KmvzLzYM3Pg2cMpoIhvp5Oez+A5qC29BntIGSFnX+6zRXA/s3WepsDhm38TkXBwD
SUdtLzW7P2T9y4lNoJIHcVrSyRcF4xgWaincj3zy6blqTaHKD1Irs2OBCzfD01oM
UxgovGJyGZKMP81oydT5CqkknXlG5d3+eq+P5QfTZQvL7QnA84pI8QmlwuQxcRKo
wnXDn7CP45WXs1zmWnNXQieUvwtC4TlKO9E1DN6z/VCCfjYlhTLPZZo9YCLMBEOm
mk/2hwoU+fnRDuQKrvkmEIXM+Wh+T4hHNjkwK1sHF9iaxPDP8iZbI5chtKNPTI06
oM+TdLhyikCArA7NOqJVb8UGw2iaAwiUGi47FMXXoRj08JPDgbuwaDCXK3rMUrqW
wDMziZGhfrev99z97b8M605Wy+sTYdvcfQGAa4OQ6V8rX1RFPNPnFkLMQqga4QVv
gH8tebaD8UC4Y22z/QtdDTajBavzgmNlBoA8xP9MzknhXQk8pnnOV7Wdksq4KsnO
eM1Rsy+POSfbo4lYFm1XRATfLLsAhjK9umCHD58ueeZ9SVtLJ9VjrPMKv4YgdKaM
5SF2ro+d4Byg/MSoPLt3Cq+5SzHHNG9o8uKldxfzBdB4JhJ+t0J7rt8ouk5AvmYP
2l+t+CW7qP45Se2g4zF/Mk4YpbHth3vSZHZYxNpdJk/fDCFx1hc4RNfJCg/w3lhi
jCecknPGOcULrHhZC3g3CfZtIJsjyYsOc9lR4UWpbAhSnNduIHye92iI1Kso5+ZM
jwbhIZaiv2iIcesn5kt2QMa1MY8U/Z5JTZ9rCEdr837yCrx18tyivqKdk3F6wELF
T5xa/496jseuVklIg9vLittPoox4PaqsZsJtygVXKH0ujLO6ilWHJq+uBBxrq/g5
9DNAPI0d6JWDsBRAAp5up6Nm7hCQEL+QZQW01RkUl8NcIj5Qh3ML9OkP3urVw3XL
tSo0dz+rRWJSCUzP3xPAt7D+z2O9Sb8qCejk1f3RCMSwdcGTYROghSoy8owiXCxu
T92WWZAm3DAZGnC8Raiy+m2K31iqqwjsSFtJ4RHq32WGlMXWOUfknkbMhFV7IWrS
iK9AFzKNJ15GtFaoCBfbmKLj6EzjRtJzTorkEXy33IlLQUyeQPyeGcY2u9Nk7ccg
SI3IH3Dky/Dzye8YIyF8jiSTPFeW75pYoJ7vT2W0s1wNA7PN5iYUtekTIw2W6adP
viBFy++l0nfBw481hlKXF3iY4uRsOCnKwjqZcD5Hc91xsb7v35lC8jQzOzaMlhqG
LKiwk5nV/SVitY0YAL6FywC253VziKQQuMjUC5nmyjVCl3jUXObi8CMOUikphAc3
Nq2wc++Pmlw4hxiki4prPvRvcMqQSEMR2JjLL62e0e1Zg+X8so4eOH7oK7mrMo0I
WpQ2jCjBiQ8afFa+Xk42PqskJzT/7a6z8ZUNoefnNMLCYw8QFwIK7IbutobOc3+7
o2aGGyVV5vFGLPI5D9BiNkCpWmCGSvSdHwE6AuR9BOmxWxBWuB6IroNFT3+9Y7Je
C1WZU0PjaYMQ3MUBoLYwMHrwSgU0SC449/S8e6oJ6dTJ7apQkMaJHvAlGZbsUgnJ
rPgLDC00ZwMKUU9oASM1oStJ7x3uxYMG2YUsUnsy3+nYINb+cfSOjQJyeF/PbuJ/
xtfVMUbRoztMJzNF8ZCHp3om+X6wiTh5j8/BxxqCZ6UHhDUaV4DXEFz/r/lIljmv
LoWS3VXdinl4zoKJvPeLRPTo+JE+cs/YvVXscU5D8ZrJxuw+vf4gIvREPWD4Vbbu
gMuVragtBSMcWFULY9xLnK3/z++D0XR+1q0cEvNr2F1SGVIPl+BAkJXHpiBL9M7B
R4YDkyizsci6Q9oWoBx8DExlMrnR4C1piQ9vHzwUqj0Su918gp2OxbHOpjxUoOEH
pxiz5o6OOBVDNVCMn9M8H7756ldQyo2XCjDWye1b4Br4S07HF8LY6WWgGdxZNbkn
1XC1xBKyChlHMgCNj3hDvTCSf9FD+Nmlrk6I/WdwTvNsmuUBKXjd7Qma8ijiIopT
+nZsCwmxzJvt33AG/tzmN7us+Az1Xu5nPfbbxEUQKWtcrDCgsZ/2ER7v+y5m2jHQ
6+ofXz86kqz8RFIOZ+sVwsa43noqequR6i5YpMCN6OmMID6my5qeGunKPasCIV+4
PBTdT1pOboTp5yRYhDUWTBjKLReuusXQpjhELEQQmGE7ScLU6e7AGMElu01S3QzO
iyL2tD5pjxyehrGEVUTZZ21xQ/PwV4tC9P3WCppxQFw2k2bB1dHaS078bRII/7xX
yf75HU6KRT2bD0qyqVC/V0XviAaO9N3aLwEIBZ3kC7vlx5siA7AHPx5yHQ3VhRgm
zsa98Ys97hNeTb4tM6KFPMDbIsL5sThzspWrz03J+HkF/XaYsQ+cyOM8LVr7Jzx9
+v+ucPw2bYXWTKxWUsDKavd/CgV1rAPqow2YwMb0VDbdc1jXa/porT8OydVJstPi
VaHXwXThpbirL+Lbs0HumuZ+7aiUiqlUTjN/TuUS4rorq4lK4U1zWk9xdXTinXO0
ZM9HHylFmSwiLW9SEJs1PYJc+cA0SBTA5cZVcsp8UN7gM+zt75fFrrmEyvmKV2Q3
7l3NkTsZ6tEGvjPTPzJE/VOgTZRqPWz0YdtJeMSWvOaZDe7v88kARHexgGgc0iYw
ZcL1OrIwC6ibj+JOQACaHCqhE7heYOiZ2fLSvc05n090XLQX1SulBCfqo8UJGAvf
CQweHyuwlCC/c07Lv4IHXkaTq0sZWsZd1NsYM/JibMcewYB3NbA73Oj6iaCtRACo
XgpUv59YATvAeY6GbJfo5frPWJCDHTtu13iVBe/anFESwvW6AFYd9kxD83Pch5N1
xlW3ZLPuAiUWi+cg49N97ZuVQv6Rr3byDCJHwDMwxnOj6/qY/9hLsI9hi7qZVm3P
zKym+WtfQfP8c7zsXtL9QzXGG52SWtpp2UChk23q1yQ68lgkqwz4MkdXCNvNRZiT
QCiijI4JI7VVZ+GypdUunLn0gTefa8TCs1PDampKgC8GMQB6y6AwB3Ts9K7flk5c
TfC/eBtTslIIyw3cuvNF7zRxLSNlWAeEmvfrpW38CN+uuqoEUVGsH13MiZF909mj
6BHY3neDx6fY4yGhp2FKzDwtgcvZfbNcp3/vtpb8JJaZkuBGOruLBfaHxGpKt75K
pD0jTLjAuo8V3n9xXNYu2qjHwQXNFuqgKg2Y5RS155QdpXprI/8M2zXZAc9BfKds
rJpSCIKepUkpjyMwI59dtYC4xGaDS9oiNczMjz4vdsgk+9C3ZkKJphun7OVogYrY
lj3kXaMBL+aVHuPLiZsDcjGyrSM3px2jJ9HBBkhfZezWmoZ4R5qgBGUM5OJG+3VA
Buvujp6g9Hgg39cgCalbbgJ2A70IfaqohdqVHpYVVEGmTiQlNCJnFMQiKVDxfA6t
98Gju9VtAuSuOWdCTc76pHKO72WfVarvEYQKfHjuauQhHDLHUd5QgZYi7oF/SOVF
jsDr8pv0PguOQ5zbjRZe06yoE9gFZVtYFkYK8sFhz8i/Vlen1GE3IEcnxFshR1oI
Hjzw8SwSF1hLy9SCkdZLcii8CuGhiHpfHPJfsfjiTdN0DGASnga+q4n1XgRmGv4w
+J1qhS0bHS7ahjkNIM8X6dXNrAGjTAJedtzVPJLvEEbzfiiPJVyOKU8GE8+yU7Ye
zzGNMuzMbrkOqSsjhC4GEKwGW91UKZ1ajowObkCPazr3PMJCw6sIfLy2M+feRTCd
DNOK3RsvmO71qUnth9C/DwNSrec65bBlZApUeYChcwYf0/w/FEqktwbyeFfmQIwq
gV2S6BKJNawckuxluw9t4qew7XCcvUroTAuhZ0EQjjYvMY+zCdNU5Vo/0HmeiRAk
SuaFmwFSZfzUnuaM/XPmkg2/JGSDNkojUT7DQ73HSoUyP+kWlRt0jlj6bemAla2x
f4XuVhHBgpiXm+zOjs0VzoO/We9pASw1ciqmCseogyHOXbdGXSJjGpuu4z491+1q
QoNHh0pkqVynXo+xhrOYAavQMXTiBMZMdSLlsvToGQfbhtxVa1dNE3vUAc38CHjx
cgHiqFEzuQzTTVzjDghOWDLhNp1EKnfOGPpzabT2KVCe9MjvvR/l5i7Xb5pp+PW9
GyRa79sOfZk5yhaJrdp+UG8RGzCs2L4Qpwjg9OahN+UfGBCnNwdj2UQiIdUTXwMf
/KSwLbzvoySdx1gyjb7WrgxQ2QdXnqhwdr8TOoupAzpf0kUt0DRr8mWdlmimP/P2
xrynFnxIoKkRmkAzbsUwQBNRbdmNPTRg9Mf/6FrWtzoiP3BijxjYK2X9MgJbNcaq
GJunKxJsNbtY5IKwGeMCPSETapyqk5/CUhIx5Lc7HhZ0KDna3JtumHARqUMur8lM
aB9RhsPLL9itO0x72s7S0dluc9OptVWVFtKkvmXFWpHKnuuahALBkDJ5Nh0lYHR1
GSrkXbi5e5OWWuMYqwiZC2u0ksSRA6qqJsBxvc0gZYYNo8k2nZO4W5uvmtWpnm9u
wtzX8rEhZu3lqPEE6+B5xJduWcjdKpRKaotOisIXeQQO7W6GqSDxqLnyxTYUXwJC
mL/uyCyL7olwx4cyrvBQtGzYIEUz3a20186K+OcCnSxIqI2c/zz6vN6E17fTMSVP
l/utwDFFe4V9idNZScmq7NHT3emNnqOzC4uMTxmoy+VQK+vzOJ9GuJhbpOfzSZuR
L8fcBeNc/tLYrTPcWwegwsmWh683Q/HDJN2hFKQ3KqbnTE0DGYVNQwr6iB1OgHeR
w3SsM6xRqSklwV+iw8S6Z+JCV7Dktz4/qNeW+PGkVBl9xTA1c1d1tsu+jslPsORX
0U6AMyhoIOqXdPMMjvr5MO/89ER8sXR9z776yb2m7CDxi/CrgI6cjiyJvnrLJg5v
ddzgeP/shcXgGtWRcXxUdlO52xccUbmBSXlYWNa6i8DTbToVFouRFVbGAJUTpxPI
KgAjVJhMqUVelTjsoYeD2Egl3zlPsdW6+fp6P/e26OF2ClUwhQ0NDvqPu/yPl4Iz
GSQVm9ceV3g6d1HWoZkK6lrxjymMsetZVITRtHT26R7aor9c1B+Y6bugWiFIRLaH
67g0oWFQ8iC/s0P5khH7dWJkRx+/okRUUg5kWvdP4uJfioir6Ht+wkS+f6VYa4rP
G4Wq4fabbjK/sWmaBNAmuXa29CP2D6f5pbtRBRMW27WiHzahtsD8DgL3r6fGJWPV
PDHpiSi/9271LiBRGK5CtCD1KBucrkZWcYC7//tjxDF2rCSj9Snu52D83zsSeWMb
vn5JNFFvU9/pVNufdzqcZm8Bb4I14+fckw5YUJ3wr222hF1lU1CypSkjdDtOqE4D
es0lKIAEDbmVqRIaptOvVGWYfXtAiQx4oaHxS3PIa+n9599ANigjpG50oXgeQE/Q
/vP3ZYtxwwWQHN9yfDmVPftWwviY4YPAazBUe2YyaOqcJAhu7Qf1lNYgcWLtczIR
42d2FDCTdJO+PgMvH5CbUuL5TzO9Tp/MIYot4+hmKIB20gRgALRtu/7DIJWP+ttb
1KLeIvWPbf0X4+k/3pevrG84lwyWOSbmg85qI3BI9bIezUgoRZvalcQ5A2tNpnqj
IoLwwE/QCiXqIKg/YDGwUnnx5MZu7/H5YpfPndcQUdNfqhhlR0UTSR5MYmsCVI4J
p2nBxMZZbJ0CcGlu4a5BngfBBdYKc0uSq5X0D2csOPeKhkyZRhe8MMZcEV0yxfGL
kJKSojBVdPv5Y0iVKWaEkMAFw3wk0vgwlGTG2tZa4WCGLfnZposj0F5tO9hsYYqV
sPmPgHzbK1JeX+fW/vps62Osef4SA4HmOo0gRDFLu5w68SEkGSm9CDYExYRWE+v8
fH2uBeWeB/dJyoy+XOyAx213nAV3VTsmF4TBR3T8CU7eVBsZMI1MzknXyDPdIeUe
xv+UvjxiJoKCiVN5ExSUxIVuiFIWProrhPljr3+pykYCI5Hbia06xeED+J3BWA0y
TRbCXTd5mpRl1mXnAtnGC4Ew9JV17VcMoHOUDy97dXwX3gCUxD2jr6Nkheqke9G8
nEalzZ/1zFS0IgHh1iuRyPLrG1EwiML8vcEory1ErHeCBaE9OzySS/pdtO2RU+t1
DZrYs7N1mOx+DuOVZRByE1wbF577kSzYjT+RmgiefvPZv9HR6QsAO9EbNknhJ1aa
A4c2JpMrpu9AqiA8Y8SqTploiNZJZrj9B+6I1RCfq1XFc2cl2gWYQ16A8M8AxkPF
ImsWl745P/qZeaKuJ++Ae0YD0FYMn3P5pLg0krlvHSr08JhMN1SXJR/h956W/7bj
U7KMCizIC4FHM1dOKZBiKZQq0CUMfIvTZaumlpl5IS8ShVdt7nj+wuE9zjv1n1NG
s3V25h25zjRR/vQLEshKYYl+kQC+2IF5/M4YtkkKTZD4uxx41FUIPa5B49u0DQBN
zY4W1ihR1YVLC9QnvyC1Lznxp2eg3dcVtpT+Kz65DZTrN1IiCx2HhcSzTreTNYud
ebkXnZ3SHhfGpPkUDmmVcfip+G4syIVe03d1nflJqfy2kb4FFZ5//J9m8ZnNlGqS
ezM1m7hyYFKlqQfxAmV4hayqcSSo29OLRtWZipy0kPgzF+f2RJPZZpZYebN2C1ta
2wurbJdp9F5B6WU9vIcPF105Z7r5fgSusW3kqgluHfsaz5duOWXJZhiGJF0OEjof
68b9w06hWIrnb/JpQItXPTySJTzytCWuXxF34TNWQE1dCAvfWeGIa4BFA+P1UCdN
mlWtveIzHi+uLy5DpA5bCyhvFihJDz1s+uQcK2cxqPICBVNgodNKGzTFqhHZ+rtY
+0juonZdym3N3U7C7eh4WQKPz26JVuoe81Bt8veld3S4urTjMSmMVWgQKszg+5/n
x/Vw0868I3ujHODLTY8X04HQL1VxiAiWlbZClJzmuU4qm46hUBf9+3kZqUvl9+P1
pxyEAc5sITszVIYGdhO798H4ZF1KTMkSG1SKUL+ckHFXdsPMFqDhmYSVLqcLOtke
S9x9Jhx1nichlLWMENGrMMPj4N+Y/8SyRRKN5jqBHbrWiWlzY7RCD05PDrtqumAL
Df2HYEaRjCzPL3JhcPDmMWWptm0RWv+9dHDVaWZa3BbZNAHPzPn48Uo8DXaBSagK
E4/hGXA2tGLwybh1+edJUBnjEj74QrDQ+0RPKuO1xCArJdMdo8WF+TrbIaOiMjz2
uuWAEuRIOEQkOIUHl5AkCNhVVzBr49ziV2uGqQPdNqPlozw9QU2R8V940Rq8KJcM
MVpfbyBHbSAoMgETDxLdrxi/F6rkFvLagiF9le78pVN3j4CO9SbTe3pHz1RGweqQ
rBECTcG0JVXS229i8ADpYmUCH9w6Mm+rxRbX1Y6JpoZKa5vpicqtsIZA/ep4cGRW
qOVzZKXmQeotolX0T0VnwXSdHejJySGeI3OutZHkbiRrSUwYi4eyth8AHqF+baCy
38YM5zHdfzdwTkXxdktDEdBn3HuecD+gWW5Y9d6dBXsEb/hOnDg99xK29MfTjdJW
kiELGiQc9wZn4Nnh1IHjbrm5ARwwFjp3FQ9+3FhLh8H9zbRinZyYPpnNiifx3MfS
SPdKI43QhaBMT+ch1RTuy2CGiehRgf3QjcCRoH34FgBvXSdQl3v8+4X3aKVkToFQ
CnoYDt06bHPtAe64lL4w0BxjJ+Z6ZMniGK5D2z2JqmuWXec8QWB6qWrQ8ZmOgJD9
8xgcxlvCKLjCkHD6g3ncd9DCkkNuuVwePMVVIeHMn0GGyyE3vEtoHCO9AohtuJks
qtS+EBhSiJbg7G5FsangcEYuRj9zRQDFCddt/UrUlNELD8nVTXbrrw1EbS+0w2LA
YYDzrB21iK6aqKu/CdS+opYRzvvrSgwkUWrsofU8M38ln+UzRH9TqUpJQDhGUZsP
Kq6eZhWdeC/HuauGicVeWK8q25OgQeGK5jlSQ4M2XOfKJkNCYFfTKOLZFaZCp9Cr
cOgucNpdUnOsYUGWMhoBhcu7NqOKHx8UntY/o/b1XGEXshcCKNvIbUgkK4Pu6uR+
sbkIfYao8j2etTqn7cGWrGhAp2vKeAuEpZ2uOCUmFptvqFuFtM2nUlWS3WZnC5Wh
qcbMW6LN713kjznNG3MvkUDIRP4/FGCyFGXcF2LTRlKzOF3tepthbzPo5KvjchXd
6O2qiZU+0bDFrM21BoAz7jqPUBXzD+bW1WVKg6N2eA2rO/kRyC9k5ttj+r9/cB+y
a12XPKS6SUpXgwpQSUsh2LstdgPmWnjj/nUKdOK12Mf4iZOTo7FOCukkFiMdH3Kh
4ICqbS/7e8vTn40sJ+erdhVAE0qXD4GD3DYJLk+f54RJSSt34edvJ7uF0tB7pXEQ
jGIpwmRO133bklSaJQMyIOc+6AW01tvYB/7bmSU2JiN+udopvRD7mHUshzL6GeNk
5W5dvpXwtABH2heOVfdaSy3rVrCu+8cOfoBKGTVgLhUsiopiAuokP9eHxvlwrOH2
oUNYFtwl7F9dnUIErAA3o04CboeR5ZsnYCnKFIRz1xhu7nPpvniZ0lmzWYzWXLeD
LELdBFlJgxDkXsw2Z/Pccw7WEN1tANuGCq+Oy3SwsGq2NDxj1R6HK1I9K/OrfGBM
FNY2uUHwZ/Boc1C2gWg8Xn2K3zPe7lrmGIl2H5hurb45zImE21zbh0wva5Nmeo4T
0S9+wtEQ24OFhVVLGFY4A0fXkFTkqAHgw37nc5YuX9CfZMjT66yyekyzqVbZsczU
A7u3Z0/C4UVVs45M4n9aOmdnU7tN+nVxBLzjfuMTFbQrVt9R+eM1QfGOVxAyrnkF
6FiDXReoL/9xJ7PvKY/cWdYCh/mM34GDOXLRIhn+Sc9PvjjQJvwjVUJJjByrNgNw
+1ODLaLMcNhimJjGM1i6jx7OrpGHkQFGmTu/XBz+25/vEuatXryx8FyBQfkR88ea
NsBruWQ4h/N+a0sdUBRfBmE2HgKfGC99xU7/3eXCmHOlqKR8HZ7y+3GRCqCNEHUb
mk6B8hycB4ulYPd4wGDI+JCM3OEZKAlubyY0a3JaH/iPdSOMLAvD5VkMkPQhsFPL
bJBtgjD8M2ADYmFsUrYFIl+LM6pE2SPCqMuU1xYqZ87i71j+iHtMwYm0pK4UTbtK
SFxBfUHMmbhHe9XCIFvMj2fqQG5xN8OTFwVqEm0AQwXzfp6L0acbnZsBOfdVUqpm
nb61FYSl7Rrn8SN5pxK/XWLN0JiUdl+W1go8eOq9WzSeSPhy2+KZFDdrSKLjZtmz
b0Aanbjg4msjX7T8+JDlbyZAK5PM8+Ya6qrOx+di/3FmuLa+sHzbv/QGmJG/spFq
q99B87GdDrUU3Qhdy0KInJzCg4fZtHz1JNGTot7fTLmDm0cSGez10nNutjWB5BPK
l+UgvjzNk3ZTVQAmM3jQNQauQjtjXjk16yBZT0kXnF5A2sJekfm4rx275D2FS9w3
KdshZTVXddixeaH2clrMCa/YyIBvGzqBMam5tWiF+ZkKlejOl9iMgKcyP2QezkBc
GaUokNhz41N0dxLB3nn5kcbIao25ERrXT2XYA6/jeyTMJAkD3pDCzS3sVc/DLSI+
oAxhFRxv4rRhIugig478rl7XyiSxngYRa9iitxpjuqY2Jt8rxQTR7qNclSedU6rr
Q3sGp6Pzv0KisH5d754vDgU2Q1Sxa/Kd4V5jGdBiSENZxS5xgEKm+tMPKA2KRReW
uTQ/LohbedEZuShqWamgYCAWCc3rJveIDMRBSeTG8YrX50SV+6PuQTgPXKUio5B3
JowC5FPrcRpNaHLBfrSHi8nvtT4naO0z84tEKDD5M8TMtP2OsQLaVi/xSx5fE5tZ
L6IeOtZji6BLszOs0Q7UWwrBmLo1V9efbeJ3tafPHILUXg8fkCMJtLCR6bc2RZQU
agmRtBPBiNT9ATFIbqpe90V13Uov4yElpZPIXUHwC2lN7gcPsMA2hr7C9qHo36HL
L4iCaPaji4/y/3Q53vKOJ5gT4tDrA2B3IwAeyqX0qVvWB3Bvu96LvyM95q2cFdys
qqiagiZFTIRur3RhfZ00VojvVNh8PV14uN2dRW+7tu5lQJvFrbZqsSJWocICBIH3
eBXvQprQx7nAI9snNFUYOoA7xTcaQI6Vs3qa1GHksP9pRMZfq72No0oZzJvTe1jQ
dhTzY+vYKgetmrGodmkUJfr4CdW0RyFaQyn3M7lWRib7cPnNg4D38pf1rEg+pwms
wv9VBFy+YSdkImWBKjtQ6UgBjlWn4LLm7bXkC/JtloHhv9+S+QnoDaeWqe2rzWrX
XXfzxmVgMGJuNEAAn8Kq/37/cb3YFuj/xPoGQzlcOZOVWMGD+iy1urSb810OWkWO
AkQHPJah2D7cdqIPK/tINn38FoJTU/LotHWg2mFds+lc+W/0UpiUDqtSX1umTr50
95YDMaQr2qbnmmSl7Jnqb99t2YfXr/KlOeqj32wrwau16OCcawABkK+4qo2HwI4V
r200wXk6lB5LD/awJhekXmNtdnGsI4FYQTuSYqYXGzEMnAUb3eMXOsobvvN6wzN5
oS3xNY1zAYpfVuUW+wCNiLzYmRItJ9+CkOoCJ7Dk2olVueqMpE5ATg0buYBuJCir
5/ozjnetpw/v9Bg4b9f+li8I49npUeB29nk1zlSxXXWkKJGI5ntBSGuDTu0qMKRR
boZj88qyEVqejidGExN3bhfHl/sJ8OGzHrbN/7SjJbx7XnSOX0uiREkjS91lJz1o
Fp840RkyblSvxIWSEdsFeHMaO4MX/AioL5I0hocJAPIqEKRoUraUX+LaPh/XbLqC
i4Wv+4Bh2rhQGCtB4xSzEsd7zQOFQpt1sDhwMuNjX2uchx0SM/EAskSNiVmD2UdN
xiR0cSPBiWFKwvKfusnaNwlzVndicnwfZBdzhJ366m5UUHY/KxZ2loHllJH2MjC4
25l2t+9+tq9PtjiqmipTPgJOhvhx9U+2FeegJsExVZZthdJ+s5/eLPqjp0wivl+d
m4+B8PNI7xThr49i2b03qdTC0ododf0128vJskLR/t4dP3Pa/LfnoQFcSlo0LtMQ
ldQVjat6EboEsIm4JZ/FxCXJiJzf0cyWxaJTqKjgcs0eSkfg08vkQoWcDd4gaQFx
wiy5d+KY+Rs5KxWH7/Zke4VmH/HpHs1Nrkk8ESetGB78XOuXYOYZp9adYoZbB3uO
JAS5xgEYJsY8XUfvrXGmrydHKtMl07hjrjhLYgkI4RfoaIoQbM7iAaWZVoqhFS4p
l1uyEYvEEACTS+d+ngEOb/f5pTtiUeT/sZw0jIcy+XYiOcpbWxA28uf2DNTfJyrc
a1jBaINKFTwFq/9pP6eZXZXx5MXogy9AsUVe+fEtugy0/uNxZ3A+HMueGvO51c+D
m3ptwp2EUecL+p7RthkCktAnN8taBP5cX9dInZry9zi6QEgtJKJGrxCvooLqsRc9
psK4m9H0x5XifVBICqpvSD3hGMjJ7w+0DhhFLVjtur9wWj0t8gL39KVfQcha2o2W
oFBioM8OfR7us5vp9v4A2IFAA0yTGBjepI8NHcZ+spN6ImQj6FUGesAIwtGyOHu1
FmF8sidxMF5nS1RUNbArkklGCxko0PA6Dg5WCDvkgznJ6ZublVee5YXVvPCRwKpM
eDooSgxfnFNinXigVKgXsgm0R8PrYv5m/7X3Lu8ElagIBZbV316mHU+QoI+Xh8Tv
chBHoEKtb1U6plgmDYQYbx2av+v54xKiFpqd67RX6J1cCp7gPJqfsAwOEryDf/AE
QgeudC+2xiUb15UjGbe+OvFWEdNOgL9J/5wFnMsYTV1bq2BiNy2ihN38jvlQ76lx
1RZ/rjiiqndDsyrikvoKITo4ZswK2oCCmvH0JJqUuOr9CTXDKBdOo4FLQugBxefr
9LmdbZn48xUmw4yPVB2bIIcsDZRXeDlxc/yhTikUq7yU0rAkpVM30yFte8DgK0s1
Iq+tIoBngZfjs7NKE7xsgTwUCAEnlSDhNcjURvF5bbObAcj4cpcgNPfr3lM2n0Ts
QvgT9uCpOwrTveXittsT/hUJ3nvj0LqskWTD4wOsgVRd0xTGKgAMIwePoPhup/R4
7lJHUCA5tIPmTaR7WDDCsiJccFpiCfsNMrYvLGHa78tTsCuDrBLdpPymGVcDl32F
GW7RrcdAA82AbXWtGzK1KRHMA1PMCXxrWvAcLYXWt8cyk6s7aV2TGxYWX9q5hXgi
GwB1ru8cfzKy9fRn3UJgNC9Dl4a9TiwuZzo7Vlt0aWt/D0Ogsz8vmhoTgux9PKMp
PrroqJiUwmfLOFmeqAiP+EJes/4D2zwLK4bMDZMtfZjQ3ce6VBx5Uzt9z5mQff2f
uu942n4Mi9QnaYQPWGf8vC2XdkGNLccNb7jsvKJ3j0qEg76s7tLfKGcH09w434lh
UZVHwcnt8RpuYrlgZaWRBx5yJSoDeQjjKUof+DgCfjDXJEATKt+AaMQBfdZ8RhVI
UYbjg8mKj+9Zu+AdtHKp8S7djVD0f5gdfSkPDiLHXtHUOjpkRBFH1lbty9XssiRw
X+YDahLjCQO8P3btVjwDfEg7Yl03l+V+D6onjVBTzpkab3tTUwwLSm/Slh4dsYhh
vVCqiPSnev9O/SD+w+71S3yNjS05Cfr6MALcOuPCGV4jh+TpNnolRYTYF5P9Q5VN
A/OrA+uKRuFxCYvC9lAoRejP3GCN768Uh7PEGNZUJA3I9YldSUpA+HiJvVjl5oZM
YEW9W9GflSK4vJqqtg3gK6qNJdIhaIN6/QlQ+hvQuWMYdqif0sH8nB8uFUOn74GL
4p3L37nytJWVDI5wKZCpI5s5t4NVDexlwe8axtAtAcPTZKEhwprbWUJWdCbWnRLY
LAN5zkO51oLKwDhpH9VmQb8lb/fE5tDWQTng68Jg0c1JKhg3N9eDHN9SMUzGdXIo
s2m6aPJbXFg5yDFD1SbiBqiUVCiRd+r0hGtCEgvWOpuMj8TCvlVx0kvg3pdzeikc
o/ecwfomfHbF1JhkbxEG0/qV8e6SZj8dnzc/yw46NTsWsAfB3hW5bi466ONayblW
j6OF22HkzUmWPZF1qhSmavysaq3f0RfK2UeUlrYQjhkbbdnpOTXWv1MPWVxOyLHo
zWQ3fP/GxeZhA/xeyyZnyE1rCC+vqxPq79j0vK6/e0TT+dh6RkrKz0n8eQyQODml
hJcM3ud8FGLgA5ZUVlVmG6KBIZ42mdNsj6gtHApoYaXLUJ0FuVimoMJdLZxWNLIQ
CCxATHJNM27dSlT4v45rVBTsbeZOC9aUW0hBIr2GAfrczd+fEjxgWKbGDAX9PVGp
WEcgrK9GCUaZh3+LYtXyf3Z8VXqVELID1xhK0lN3a12cSETPi8YsPHnBljvfkhUW
YqxG0l1BCjNcDlZvgYHRRheVSqzU1nfJogO2xCatjnl04vGNbpOv8IAJlAIwLRkH
ktmR20cHZ+JpVXI7Edfln4DufT2IVYZon7mC32lcnLH+hSf3ONcA1lLe+5cVuind
bHc/WeYHjKZfYU3n00UahH3Xemw4Rjwv0hCDJHqTi18rUK40CirtPVwp3Z+fDZqo
/5OVpAK4jZwJZbNF17Sr+9OKH74OZI3ibwPpCQ0+uAAOLNkGrraQiH8rORGHaPem
DA8qBUNXycDxmQnGQv9YXRfhVaKLxbDANmc01jMjAhOHcSPxVlLdEpthdS4sZGLg
bAD1HrRV57aUZK8VnA3G/T3UKUtMde28gPkF0exQIUmwUosEQ8YO3I3G21jzmaYp
pX3Iyb9qf1p7WhgIT/kHkvGTjp4/U20qpVnvaYcHsGBnTwPqp0hT2jPw5aVWr4iU
kAgwCHtDSGqDqRMv6ygk57OJNMOJIB08/dwTQcigCka6d4Kb3UbFHdUQkZCpf5vZ
dmMsSx2MRteJ2zl02J0xc3md8B2eu/rUvQdS2h/6qso9IAXbF/qTaPR9W7Up1zzq
HxL7xPsvXQYcUBpABwzG3fLQRciQQU8MNlkcFFPAhf930fhSrArRvxAxjrGVbTum
+x8aAVEV1GRCt4nXBvu9TesI7/OfxgL9At6jcT8QnnhP2F/u1hBrPntL8YYltR2T
p8m2+QG+ZUABBwqGJQcz9iiKWJZsko2HZ2/idzt6I7jtPB+t+H1P6Q6Gy6l/L8bM
xIJSCcmLIC1sjivZBDl1dq/PTgn4vHhr3RfwuaSVR5lKdVqiq3bFSxP7FGnDz6/e
o/mleDgDBBMaTIlRESgxJIs9WPPmdluLK50lHqWHywHJtSy9yZxu+Im/il9G95FN
B7NuS7F9RchANQJBouDbecMbKuENqyy+NRpkd38mZOE0Ut5bCxEyvUGTsBBjb9lZ
EAknRLmRxLMLm/fuP2UTA9VhFy1enn1z+TxMNmILa0BE+ENpBAExWOvDp8fBEIA3
J03P2mGJ7RENbGm9VlLrJdsS/hdROBn0ZGYxZMl+CFmfxJFki72Ta8f1b/Xy32cX
rtM3GBtC1m9fIjT78J+q95ekvSLyf2U46hLq10P+TUmqyOxwBCCPknJ29OZDjbC9
sWvhx4300xMqmpc1Hc6GDWHEE7vaHMeGZy70arB2O5CJUCTHbl9jtP8+eCLfiic0
JiiGt6N+rj9A/NN6rV0Of52+KSoQElO9mTKDWKj3WIjoDYRUf/Ay2B/GRDMPwKKl
KBpfcAlniE0Hpm8BLnc+WaGnEkDEqRwnLmcNaRkDMcDJo1fNvGdUXiVaWNfsDxYg
8/fS6IUDBcmNpCjNl47juynfhlePMYZR0beADtfgBp9cFdYQh8mCXdtkXPQgnLuA
uYba2SxvTM80m11Gt3Lyu28VLgwDz+puBiMoV7+aQmZheFj9te5KawwdMjjuLf+j
AU4u7Z3g8ZuLNdLkd3vW1NuJzVQUFnu/wFv2AyCgm0fK1naNCagVzJI154cRKxSZ
fQo3PGi66oceimHWKxGVLPngqtt8kRrRAHSu6p2LTfCann7j82UMzodDfumqGueS
rzeMG2l2nKTfJGDEEztzKLKdttT8vyeUq7v8mIPuoZB4771exd7IDCaGlXMq8isE
oCHJK7LIg680THyqyl25cNZTsC3SEkS5joSxZfpLvsxHz3tx5CGlb3uHUeaiPlzc
beMvRHB8NZkCWSFIsArAK0kRf4DJP94X/gtzWjrig9fH0WsbWtfeeEsMs317W9NC
GM+nV51ycSj1zNacom6nIJV+bJvU8NTSZ1ZYT+8Xv3xXYajac9ORGA1geS8L0b7j
vOjOA8nTSILyWKGg6Ukc95P2pu1Yc9CKraZH9DfJSotHgHvqchAJbapvO9zkb1oo
+2fTXlwkC+xxP4yBxMGW0Z3bFlKCE80b7QZnr9TTmAc9bQCqFI1/rhVdKYFgTvRA
sONXfCAJTlO7ZrhDgPD87eBjy0ZhjP2tqIC9QqfQfV3BTxm8MLm3EMM6QZdJdzjm
eDdewLV1gnLPtdscMKw4hF41bro0kWFbQ1JMg60hOrhM4WylH9CDjQdfC61LSPCx
8Ovu6hUJ3ACAXlOjl9I4i3onL4yR9hMDNWyn3kYT5OcI2zmAQJsR6sIvM+C9bW1C
4PTWiTi7g0lGvLKbiMzvp8tliulsAYbp3eUr0+RcaJ8lJ/gqvsJ2URnxeNs7EF1j
CG56xkCWq7JeCRfXRY5K56vSpwUDHdZdgAfG73Id0b7MPIa/catwNk8Mhe+mNqFb
Exdwq3tfZTaKeqwexysUT807jvry8MLSTm7phI/+Wx45lbI3n//dnwP0aYiPuuKZ
UqBjvA+LEQDPm5I+S0liD6pyL45LjnFl/2wOIg3xN2i6gWyuHujWjdkhZkoPiPMA
d6dKM6E3u/+V3woglwp54StA7t1fVqkapQXNPR5hqIra7xnrwzJLS3u8QRQSQhwc
LqO3oEv2/wnWoeBz4t4vPsR5M6ZZKc6RVMYCgeAxAq+w2cgn2uFvOb57zSPsXtGg
9bKLjJM6Igo5oYKOmLmgwi1pSmySrpJFgbruSghzlcO+DsJx6k+nI6UKdxbCu+zI
ihQaOt1SvXdax1FwiCx0HMKxH1w83HGi/2B3keY/uDVTNhAKZGfTWsV57SBcUWzL
P8zZlxG9hjbylbOxCWeLVZoYRvblxvKEL7cpm5pAxtYxkTU93h8PEULRfiw2+Yjn
Vlhh1J87HCPiOnSIqSOHsP2z+YYdtkEr+zHrSzX5ukL3IpfrUCrqna++IluHyw2m
Xs+HUNfJuZUi0mqKBAUHyL9H7iamyzr6cxbUL6BxXj5ZAPK/mmPCFhYk8/mx+AG2
irexo0K/Zus5/Uo2rz2xUeFtQDiLlXmwNjnUNObJfKpcZ7bDzv3LdisnIrvGWURf
MtUJbMNWYS/sELuxAc1K1jTsErSMOWGaUqnINTQC3DmqRKOutnhUKxJaj12KMqXe
inFKjB/vPUw19D2lIR681NRNGfKCPlrySAXXxmOXKU5TK9FG3t4OkKjoCb4NZFpL
nSesEidPG/VvL+9cqQWU2T9SSt3vOWL2BoLs0HrMytJps1sa/FaE90Mu2/LFT3dK
G+vTLD3dHdSVkDCCKhtoGujZjJMXld0GWeuTYEHlHzosJcvzojIfk5wpQnWFCRAo
uA2JywbiUq1LyxKktvyhLglbgzFrRtCUeNQmEpgZzN7/JTYeKf/HaDf55G9Gyx2z
uUyJdGvKYYx+Ww1MmyMHVf1v9nWCVB52BzOzBLU9MsFZWy4sAFoUxZQAgLOKgjG3
hb+Hmc/10DxptXN9h4UOUZ4ChI5NoDDd52xCZTLOtaBRzF/W83LOp/bxgIhFDepM
NWEBjYtD9/s9hXzRpYFnYhl9UMRSvyjv7c1FLe1NkU/jIkobgZ2QGHoFnSb6ogYw
uAklKCIFKsC+74fyHkt5nGyiv0tpLFeAgX6d4SotVyFcpWFlXTISuVpKMF0jdFW3
f2whGP7ne1HcxnovGp9fYbe3NxW/J7Ur6x5yNFb6PzNrrLOSbt/9ZtNmD670fMqE
uKeoZJb8nX/565sg+JtXgg1kJh0CcPRL9J6tuAdwJOG92E7vpiwbH6czhZ8beXZB
qvUIx6D0VLO7cIpxo6q3g5IgRQoEBLOsKu2tdC6nTqJmL2npD9Qx0IhpWvfxFdRA
THffyD+BpgjMFuZbnSVQFOelcYLbzRTXdu1QxqtMUmSQ0LoqB0pHaWVi8PRU56Hs
HYGxFQeXrHzdomXhvT36CaZ0lYkwSB5NiAjR83Qu/zwAw/4Kor67mHVAI/mhcoeA
C5rOs4kuGo4EOdByf84MgeLUWF9UiFyQrG3qkOGhz37CqGAXbFzUdypSLmPb/vkD
pg5O4gmGRJAkDKVj9x34sZuHf7OTM0r0j2ajjIejarSqAIrc3cLgxNza4B/kNhI9
z2ydjiwwsN//EP6GnOwSrtLXw2V5EfEpFLnPkAdBOhSLba9Rqe3T5Gy3owKGywQP
3Od6yygreu6kfSJ1YOLrrfyhUHVfczAD1c7zHQUCFT+9IeWog1cU0W0JVPX0F0mD
KiWRCTmlwTqj2YLwFIBq/0pjU4V1VLye42COYGoi0kcqczirirtPECGxvnUE/Gsr
pYhfiS3PSfyMdfmJBq1dVfK3qJux4ujXVbqgdrMMmsDfvIATC2ay6Egqc49m32J9
N6bOKH4QzntaF7k00l0bjIpmbqX+nHyWjdwZfpV/9fD1EhsduFcyT+l+80N+xQ8y
729b9fUmXMVnaJsIQXTdSpEuaQtW1FzH5Yc/eLmeKTDaMNB5X97ngFPZWyXayVyt
RBgq7kzsKW3lD55smsRF1fh+SvVyZL6GEQ5VEO7oijwE6xkm1KsGqdxCjQCovU92
eRP1lpUJwHgUaSYp9JlrOH1SBccBJSQ+lZVGeRplxVc9Ai9cYnHVM9rFigc8Kxxz
OVYxm0OIhwRd9OWXMkt/dsbuzxaw/hbiVULzD4oUYIBRhZwNcbgMouG2uShCj6Gt
lJN6hJt8whv8mYE8fWPf0xqa+/vRnjkOMbXvCioEnd6pAOZadW5CJF/yr5hkxBxV
WRIPLlm6OV5Z+czpSDKZAwyHpqLaejTnvy1V4ko2roB+fJDuZiuChDpXU34hGJ+y
2GIig0P3BbsPMhdMaQj4NLGbvE+91L2Aeo54bTrsR3CYwcVawvrbVJB+6Hrz9mkH
nQ/Sy/ED7GjkSB21s8lPdO7KW4L3GdevlRjJqpwsPnnjrw4lZhFICnzwwRD9+rBk
RUj/xg5YA9skxseojR+wGrZteGjDqoIQu8PeFrzxbXZuIkAODjEpJ0X5k0pnsVx/
kW8RkTijqEPTRj2+QnnIo0ix58GJiIdZsWBSksQUrVDeFh4j+xjUXAzRZH77+xVN
iE2gTsNECgkRIK/XW+jrStmlQ4naIC/wx/OnmjBJUJ4EWfF7lqYuW28LDoNEYSdf
+cIV5YQyJI6lzQNmBfuAHBHWzDbG17a6sNCG0HABccPJ3JS3svJ5rUIzgOwr5ww7
HcYhLs4Ge3tnaJEb9hnK7VjWM++JN9R+5KoQ0OSfMd9AgkS95DeIcN/zuXUEIkP6
nExco9nEzzqWxJ42/b6ERshUM11x9C8NxZ4afoiL8u5xbLMPNFuWy1s/uiG0BLF7
a0JbrvZD6xxNv/Tt1K67RWtB8OxMIUsaaNXw3oQhEuThOf/mCQlmxxWUjQj+L8rj
B15n/tRd5n/DlPNHWVaNVoKGRESDCn06MbGYV7vUF3+n6zhQCjEzkfOV5HBzYqVK
cs934qKjKOVa01OS5qIy5JqGs4y4c5YAZCA9wgu0SSuX3fTVdNitfew7KhfL9JNb
IZuoX+mNEZl2FRRnhG/RPIWyyL9MkJh9gK7BZ1gtZWZofnL/yXg1aZ+XtESaHsPK
5RlTEoLTU1G/kQxATrQ/pj7jdsceCKtcdZf/PsotDXzPyzXFPZOZG0OYsXaRkQOg
HwDMcAhDkpDu8Y6nIagOb2YTrJWZn/WAH5ut3Ueh2EfVmJMWrGASoFzlk86W3f8B
sENTbOPGgKuMlVEwxDPt+j/yjwdjjKT8hJHIb7k6lWMqA5VpXYC+Li/B982++QWM
5YeaSMjz5svYKOqCL6wWVot593jiXIFTPmXSWt6y5GIv8wWLTEN1o8pTsTS7FZtP
zZU/KPjZt8FSpVqCJikfAZrfb5DnTkyUwS35/xqHIOdB0yuY75lb1cMqZ0LOyQrt
y/kU1vnNwfn4lIUJ+uZnypKJF5z0W+f+b+LZUpV/+If6RGetcIafuTQ1x+mCATEO
tUD2lbgyI1gwvVZ/2sV9TvLDw/pVcNvLp2DiNY/BRGcxqqjdBDCL27XCSlJgT+F4
HfkEFNd9IOaDOsFjGWYRGidxXjjOHTn5M8qaXXZmPjfv83XMCLRbcIFUrRfTgZqk
bN5z97NBV3yI1kL3//hLCi0EbmKWxH4EWl1QLx+MvoyWGfRJ8F7eU5wGc7wNZ7YM
JtGH/XlpXx5VX/UM8NB+F+012HKeTSvMy6AZpBbRhazXCZjgdLFvVJO5JjgvN9cn
AhW+X3C7RsHimjclPepjOCY177NCuwoWL8RSn1V1hZRGF3juNIPqh1DIw73Nn5UR
nDpUnFo062m7gKpnQ5unsC8KF0MiN55F3B/dDcgfMNuLwzjvNWgT//+2eubux8TC
LVfWEWuE2s5Bje41SnZffYYt+tRkNk6U3wygy0ekE4YQhc1R7X6EdT2TjP0E87bt
Ja9UNyibTUpaARsb+6NGYiPEghDXL0Ra2Iz2Ixu8T38vFJ4qFod7EkN9rQ8hQC0l
qNkbittzjimbyfobZ8QnNbbDjfKFeFxbtaHngTBOnq+JE11hkgWvUQ+3gt6w5Ubb
OyMpDwIMbD7CDFJke/n+YdUg1sk1bxrMNS26culgikZcZCtR5+/aZheVng3SJw7j
IISvULE4HWMl2p58Px29BvyqzNS4/QaiX8mC/u3nvwdA+sj6Z/4rxU6LbW1b06CJ
jl7MxpkwmPQB3d12SV4FgdlRH5Y3ypWI6RVbhHb65/Xq8wtK34MtXIcOJDJomWd/
dHgLj6jldASRuwShpVp586ciGOF59+eo9Q91WhThKo9NOkCMcekO9pec6YvMhrNl
JIiJPip71+qUn6FD6/Gb7RTrie/2OWviV4UNGPzdSzkUOV51OphlUJ1I0vSaY217
trFGZSkkaIBQeQrXnZWjScVgzbMh+irv85r+rsf2Q4JgjVl4ERBZWPLUDl8LJjcZ
H4Feheftk/UVuFjvRDv3YLa+uloblVwca0XLxPXZcnz1pzD6w02DdMg9g15G6P06
6Q4vNK7ithXvgq6xzr186EPRSplo7sHNgQFVkCgBnfJ2EW2aCVHb78o8zuqggd+d
iDW/fs1UIyoXWOFNqRWn5TBm7MO2p8rrog0TRsLYKGak9t/J1J2jHJITo8m9dCUD
J4q2K8YYFREEe/xYd00RdJDjtNM80ESjPoeV2J3FDezJcRr4s+kgjzrv0FJ22umz
ZHV/DRwfcvgP5rP40aj11fK8PO6fT31YzEHaeQwWopW4Rk3xMAfy/c25rn9zpRgR
lbRuvCgRzB+pv0Tm/BKeLa4yd6g1g2/9E1Icv0hoCxJSoFlWvU0FQ3UWc662+sgg
JNYKo+1jQr6p3JttfmkDCawEZalsbH6bdN98tQD0KcaifZZu4z2Xj6a9tbGFK47n
6GGm7Wsbg985WAkwViCTi4HRo/ZaT3s2GhUYGUoXqJnoCpIrMkbIiUTbWEOI6yoE
SFcE4OkkTHA2U56Unen62Ju42IAxMWvoAUUPxW/Vc9+I4p14wYDAPYrMopdL2NRN
IiK0saE5X+llSluSna+3ur7MhJeFbhF1pXUkcy8TXdVfM0eYE6XFI+NL95V5npXp
M+UZWKJ4Mwt1sjW5fgATZYs2+UqfLZNNv5eyjVCfE9QWnX6EmTmfOzoKp/4FJI2F
0f8WLYkeKNivD6PZ5gzNs30Rfx+IQKL8FO7qIKa070K04pjXObNpyz+XLnfefsbN
She1FruJaA6OQOGx3RVCIq+GPJfDj0a7hBglMUVQPCaZB8Qkzmk2eMcL7eada2jg
GU4958arlWEx1a6UEEauDXOJQFzoPtpuAqB570bkOncSnNh6GENtgXTzcSQad6cG
neZBdvf6gfUjV8dOwu3LUcdmFoCdSvejPGfFFLn+x3CzFR1bHnSjTGoX3LaYNdGI
W/2JVfTKRiOcl3UscibhE5HgB/YDpCaJKPHCTz1UrtI4hRghoCWp+mMd38BbEBX7
hRIXnncHOykPz5p7ecUi5kBZ9T0Lf+RC3Nxgt+at5oQndPEaJnCPKNUb4GPl0VGY
pXpIeTPSN2QQySMHYqlmlefDI8voOCFDXCzgST+bt6ccIwSvBV/27adYRfU1pTms
2lpG/iRynHphHec70+ZErfR4a67RTa43vzQYiL5tB2ehjRUOBMf+a6zWrZzdZpbd
lX1qjkwL3ALoHHZ3jkr6IT9UT56eDbY5kpuViWNoJ/nlQRyOSqStwl7Vnjq0UHHA
hHiCVYrdeCI2Lxb1bu7rc+qXKjSmq67IZYLa2wYol/Hf1Bbaa/Zx9P6mUK5lcZea
sk5z+DPaCruOBYScRRRdGA/3KfpquhRxVZXowwlVECsLFKgrCxsU8AzcVCpEwGwq
i761AK6ZxXFOiS3OiVHbE868aJyJH70aCMxzAKC87P72xQUzCVbUB6d/MsraOKIg
nwtb0CytNrNpWu9T0TZCGyge0bh5ahjUGFMKkQci+jMh2klncdsQZL0EoTIRJWpb
4a7E6w393ZsHEWCjVtwoatD+9RHG9bEF8Y/lieUUgGqvHxUcBfEFPKAxj8r6zHit
QILk1Ogp+AWPc5xCGSrpVT6e1ZhzKvwGuJV+e9b7js4m42e3V7fp1zxa7Jh/grGH
NSfVF53l8W6ercJkMkUKL9PLKwrIoYcS/ZhhNqkuEtJK/wGvBhnhiQv3xlVZhFBS
a0MEkHcWpK8rLIbUjM0tzcwqx+AjsjeN1JB4lmc9lLYugF42UTVESsN9gWCWRKz4
3CE2WhKYdvt+nwURiIefN4DxR3crxU+Rzcr6+cDiIipehxBamzm1MF6UnoYltVN3
g8P5EMHYHviYwO6sDkKQSdm0aKoQnpqfuF0FHyp9ZsBDcB9R2pL0I0VsXtXtmuvs
Gsb0zrdUeME1rgSqZRIhH3Sa+zCZTZ75JnYHmzwDwfrxKgJ3FuYZBfQQM3NQppYK
ssplhVN/HxeAClA00UnX6EK/CSnsQLf9KKldKHrPzGIhJsQwFwOTwNpAgKlwOzfR
tRb2Zicy3b5gd+dAyqP9oe2uJqonVn2hMLjEcEXHTf4BRkrvZzC3UQqCTA4fUuyF
3RjFjPPFq7wzo1RuMEreHaE3CeHTaDveMG9QM23Mvnypf1yWzFf09ncHXapWQfni
NfpdFIk85QVXKaV9ReT5raKfhTAsMe0UN0KD4ZwdCfqfyGiGnYUOeYBuEpo7/uwS
2dT1QRYa/5DpaczpIwk/rQdsIQoH72EmyUnoaguzerwEvvMMQ4XiEENYl95cwZ6U
3WTuAoysF+mlXHhIZXhgMM//rTns5f55yazbBwwQ4nOdPo3t205mX7YNJLPLtQKx
1364HQdWGuaE0g1kNXH634lHWimC2U27tIMB6a7Rb/YfjHPoRsxWAF+uSPgZsyWH
Dlhw/rgTFnLlNLfvmDfxoTo4SJK5DDYC9+qjcPYk3OeC/7P4x0L4Rnbv9N7aPQan
L85vV8dSt5Iw21Mtq6QP7yndLflgXorN6+bOtGwYCtygsV6XQSlSZnfBGAklwDUf
Lszlfz3XgLRQeRt9Q7DP0ZPf/aXx9MKvzcDZE7m2ECjQsKTVp9BHVLBpl/lpAsGm
f2HBP1WzEVQBbTl0XNSimVTDWo+8tpzdBKknkxUajH7tvSF8CmBSR0YJ+y35wCQG
pplA8OOAoWmhfRSLtuL/dyyyoVsHG+yxuYlliFwhilgBrAs/I25xq6CxpPOAT+Xt
TinppgUgrMtX2zPUCg5Gcv7UjxuaH1nLLEH0FOQbf94XYTKUXGMMOLLqCq6vzKjH
yxgik/rOqzQown8zpD/FCKFPw3d/Cshi5F3trXPAmYFa0Ng5VjDBbC8PjGsI103/
rYFl0u2HXAobReGiMyN0B02WijOZVSAuOIk/fgSRAr4OgOnep9sECb1YISy+9FwJ
+AniQOvt2ucDf5uj+wa4V2/tzdU4nxHmBzDqXVQeg93oKv1Wn9wcdxaJTVHXUTfM
4VSyr7ksUB+rp409j546Jy3cScVKxV23AztFTtZq1ROV/LC6el4NIDr3mwxjycsc
TWoK4HC2nM/yhZy5Gnkpdtfj+iSAD6Gnr3SszkBfG3Ug92QdF/zSwW/NXLN8dyo9
pM8RixuUt9DZtQv4bVNLSjASAXEuHhl5VTi7rQezgFVI/o2U3xZaN9PENIwVFJox
ZOdUcbdeh+jP6pOd3viWk5GqL1kT7u6lJFrHyTVaDmA5RKotYV+M3d10On4YC7zB
cGFt2Conx+qVN05UAB2lnK/c0c6s9lbahebJnjPciNzsweLnFRg694JqaKw4VqlF
O+oFQ170e764NrGGIG84cwlRAr2bKsPffM1b94m245halNkKbnuKNt9mOvEBDkuk
ec3OvpLGBeJgaoXemo3NxVSEJc1U5I1WnRpcKrrq4O/YWm7X62LOSUcxHeeiFhOE
cg/e06zuO9xehO9RUZH78uS9RFCI/UueVCx5nGwm2PKj1tnoz338L1xIu3f6zQFS
UujZTCbh9eEwaFAcUv9T8RCXitXzXFoPN4ST2v4HDpx6ziUhJ6IgXiSYyvYGAgfW
7ZbexohOoRR0sD5FVOfb/ajN0B7lhbZCZqXAievJh3zKsVwZA/gujSLsstmkcYp+
YKmhLJrUPwm/lTjoi4BYeM/NDNoZHw6Q3x4XEAUdTW8JfClsoFztisxMMObzJj2+
FYrfCdkgHaVSz7/lQtQfmV1fLu3x2YBc4KtP9dz9k3D2+7NKeud5xVxUpjmXD6fL
zXm38/6nI1Wpzvv+KrY5UtADF83/JDoXqHucur1xbnw3iH7Y9u7O5vOIbv7hFtrD
xn3gbirj1g4SAb93n2r7IYE9wRL1EVMCWS3pLgqbzkkdlx/0mq8KGWQ+nJTsiBJv
IA1SCC879NGeO3PvujJYBc0Et/oFtMdOx4b09NH3YI12tIDm9ke0GurtWoLZiNHd
yQ5oCr0rB4rpL7eQul8pSjOqby1U6AapxWtGxWvlfc8Gai1TCSBk0I8xyYPN2fzS
+TpgDg8HM20RlBM3AIa6p9xSkcNsBF8EKbv9Ao4Cc0bzRVpfEeHytL+y1SfCN133
8Jv+Sgh8Pcwacc3X4AEZe6jh1QTu8usylPRkhPNTXGvSXj1JQjaa577FLixlkAO6
IGfwcgZe8ZfXiz6tZ3FDu3yjZeRsD3BM/4zAVS5tAdvQikq48aq97UWA3ZOg14ja
DY5kt/r5sW1+cdvR3JILpCvgVla1/anvZ5Gqy8k55OYHSH+TfyhHfMICwkaTGuiR
0wKnD7iMEU4Drk5BpQzZMgWftSLuRPyn0zwzoLtef8dMhvNPubZihnsoU4rAiobw
kgdCmaEfjvcrkR20ysJ1CTrEcAgS65fYQvojPQlPGFVGTfCaNFxPM5bW6BaqLEuf
Acpq+SpzZdaJ/3qMQ00LkroJR1wGZHH5WGr1yIJLpzEHEadYduk2gR2KGtBnKku5
zd0p9XkT95xhOXQJC0xvIwLv/oSWcXuncTLgl76hGff4jaCvWENhRMEyD3jxMPLj
lRshPeiRcP2L3NfhMs/iSOE9t8nE871jXeuRgl/jfRiwFfZ2vrzN9c1EXPzAysLB
ns0V+URsDfpudhfrfkelg/HgV8AeH60yzIDLDCKcHX71i5CneCC88DDd3KX1dOkD
bAkb+YymWrTjXTCk3nG98EtuiB6ZPWhVx7tBBSeCGf29xNrSfKC5IMo3ub4I8cpa
b7sXfI+amA71wfqsibcMwoOVw14WUxA08ReU9BjZsirRb0FBZGKl2ixRnxLOASKA
+ptgXKBi181lgodM/RyT6vA8mKRBZ6LbqwDDF9i4LGUZEh0Oa0vNNUTGlYRxWy57
Nxhk57WjD6fJbAGMQvCtHC0iCv6OCTfMW9klLKvgfP85Aryq79R8NdlAa4L2vYCB
WzhBRs530ymt/SqDMKVuChsjUNNeinsTOrS/uLjX4LiUwmd+Kt1mdBO6lEJF8FoG
mvPvFP3eNeWy93VK1MY9RCU5RoPHaBfCoPioJmWQcpx2WOOrG7tw06HbpJOMLzAO
5WoE+ecJpr6elvn5Ufno+tU5D8nedfRNS8VRaadELD+2qp6cGB21kwTCkJJ30mnf
AlwCjHhEJGLoNxq1dSejRyesR1QaNgnKk9v02nBxvuSQQOm8d9vUJCEarDU1RIMo
3nEqTVMnFQt2Cn/4UkKaR6nNHqyE+jw3DpJygJZ7ftAWig+A36nh/GK6QWAThM93
BHRfHvx7Yffa5c9KOnxo4sHyNpZIOFJOu9I5gGPztlKjvWchFLv1LP0C3LwHGzwN
0URXQTSFlbj/dO9r9uKOBUDc3oda/5IudsJY/CRtQ+/GKAiOL4CGCpgvhue3q7gn
CPOqNPrsgRVaoMVx96/rSXtb0Wz/IkhIvbNwQiHVD+fUr0sNP5XYm++EoR02Xsho
73vJQYrUbk1g7GvGtWM719nnFzgV2WKwKbwFowMW4B5mEXqcVMiYWiKKkZyyR9Nq
F5O5RLZSVqodb1Wj6UCJAw6Bel5bz3jDfqjhilG4HxLW9JpFy9nwiAjCdL5wKNBn
JJ2IYn/HMcHh3oTHq+BabplQx/fuhu0hH8LqbmZcCoQShvbhxVVo5jOj6mgUdmri
z1s8IlbV9O3+Io3Fg17lMUYuSK/p8UmlT5dhWhOl/L2hD96itB+2AZbKzdDG50yq
KOyJcE2rmkH4eO/64PPAT9Xl3VEfoJxz0Rg1bvFzVhIpKkVcrIKmunexTtw07YbU
Zkj0vezFCSDcpDsFy0V64jO5JzsVlt1HAP+DhC3ARTM0BhC4S8rE6ZD4fPd9KvqH
DwFKw8hY5EgwJMnWxoe76glXcXKgs5XlJ/m6CS4Au7yaCTSStcAN3VuQ65Zr1avb
ElqgU1J+GjDYWcqlbpJZv5ZO84gkS4oMUMY5yvCSmCN7DL6KuJkD8eQHqOK3Ym7X
fRsH9W3F1y/rpPxz2qnYyl60QZaGaHpcUW8vRHFklu8DvVDnV42oAjtHsEtlifQF
Ajp5WQVQqm3P5IMLloaDSXhf1RkCympPAaq22Hw8WFBTW1ux77BVgkBtW498iycr
BdQzGxGznB3uNucvE4WXvdNvXu0VSVdM6hfj+zQRax6hVRdxNITbGIW76MGpUE1K
nl4vNJsGezZa1uyLEDN43gwgThqLAXIDh8uXdseKfP1BgWcOqR2GlYGzyHQc1Fga
oyX7YMn1+dLYlC3RClKhvcdBYc5543zez3NVubyWrz5AqGsJyu8zmqIustZq6yZl
HHHiq8jWvxvGsP4j0z+wTZjArqzTvws4GQ7+u3xblhCn2FpHQz9jULZuy81BTAga
hWITzGhytvKopTOnJSsELOPQChtQileKK6EVIIQ0omp3/Que7n2414s/ZTlPy9Ck
+kHSbQfUGlOEDxU+HtU3f5CziEIqUY1NS8p0XDuL33Bc1FcTNVhmjRaFcNd3FvCP
kQBef1BAVSPOHT4YKA2Bmcxr6vXEO+UzAx2eEYlG5dac6UR13Q6cBxn8Ih/17aXX
9dDcfYWUm3/WGpJTVnrf0lI4y/yvQ1G5i+vEL2/BjR8jYiI81v74y3w/EmCLCtqb
MdBfqgI6fhDQo0fnj445QMNbvdYq6OQppYWAMyyFBDKyPskP3FR5iIHHGUPq9aWt
unj8Ht2BHs+dGcPiApgRlNTJdSymJlnTvRx3FRSiCBKojgRgk5KHCRftHB2+kTPj
IUU4pwZn0yugakF0zWyR3oUOOU5yfq+XEMoAKiJ0fT6h1/eVRd0COwG7Grf3itLs
Lmx2OVDhejJ6ivHtW2rPSMevoFIgSFcwI4U57yxU4YppLlwmy0DwNGu0QA2JCRJG
rg/E9wCBZBKR/LlIcJiTb3s0cF2NC8nUpFB5BniOb/OZqJGzNsF2uKxohiaYrIPQ
TGBHkNF+tSQaSanP0sa+VcM7mtfa/6FhaQgxPzL0PmItY+2RJz2EYPE/Ivj5EE8A
OpsWfAazdCklR9w/CVwzIHk9L8qWPCMTZjKXznk0DXwwYXmtjIHwK9tMUBEP2256
hDJw7uabi/VJCSHgskGZtWh4M8GzOR+LTPL70RKekpwOg1oM2P42OAN/QqIJrHY1
5vN2TdJfKMRpNee3sHzuzgayI/vbSvvf1hkSxpFK+XqBW2D3OMkMFIOQUmfeZpSL
390/U5iCg8wdKa1YWoXOm2uqBaVbzsrWCm7WO6LwRyilc+sBCJ26rJjn4EWqHVSN
HQo4M4ll5Dyr9JxazNN8bSqUckIfbirSOQVWm+jvtksD4s8buueiaOPTb9LCTgUg
tEiJ/8KXaQbDKat1KX43mGb69VWukncT20mawBfU9FZ8+D0Ow/3py4hX8hhb0CRT
zK6GYEGPP68MCpeoEi0twlnP4x34GcrXDZCkjgNdchqTZF8tTNrHsdoPEUo+tUpF
OilgANc0LyvY+JyzuJWnh8ITR/z4dcfMu54xy9bgRuF7I/NiwgLTwie0Qk+6TWUD
OOy5aa6ITuCCsGCNtk/VJAQ9R9BT0bCuYABo6o4tF5I1jIYDd3NloH5C/8hdw5Cn
icPGxOLrWHlZ1AS3+Gvoq2P1rAhBMNEeTYbNxHF+m6vk4C3FX0GrpIZwxFCzIb8K
5TzgUkH9Oos6GsAveAEhC42B7qF8CpkAiwnVtMTDn8SNki3TRqpQitVGNUouvYJl
tm6H3CU1+lPSrhSdJqN1jpieT29FZdBLJftk2Ms1SaLvJZdq9zyEp91/JICYFeA8
FlpdihhLliexdPjPdzktBbmR+qbbWkhFHHraph5F1U4Pwkc0rhdba0HWjZoKiNqQ
4qfNAVFBCmMedp21zm25EAzjdIvjwCPioFbqtGTFNNNIcFh/9Hs8tK0/LcwCFUhh
bIFNhojr2W1T0GlPlew6QIChhUdEqOEh7wkacby1Ozvfd3w0xzs04KxFD9PGCInu
7BOHMXVbfWbqhSyXY9hFleuHnrK2npvjLzxzh0Gp0DPji95TBK0hcg51b+ii7W2r
e8pM/jxRJaCimbv208CZfbR+nvamxKLBCdoEWElDYRgRJSbMw4Yt81FHd3lp76QB
oHlSlku/yWzV+CanJf6nUkJ+TvfPbPFG+OUPZ1YHrMr9HZ3nRxw+2OsLv2byC9M6
Zhczt1L+7U8zTC0TINII/qjB9rK01gApMbZLRpq6LZi4f+HNnqWHGy0OZs0Mb+jM
xsatlSlQo1qe7k892pf6RKZ/Bb3jCDPU6xj9CIE7DwwY2Rq2ot4xcit9uCMjobJb
gvZsjemYFU7naGYWFCtdm5IkG1sKqLT5mWW0aOChEL9PIhRj+wkLDGC76v8xevNg
E8NuQA6rccN5CN9Vjegem0T3oERnBZAXcmrZnsTmdD7BwfPR+9tRBujT9eac8RBr
rIYtZjyAULAXNdQJeqXW/C5Jf2gbyqb78T4xSX1SIGZK4PQK87E/F5VvKW/5uqRN
JV9SQy366wL5QQUvHENmc2243OT0ifksHWgq7GnMWZOJ5GJSayI1YGQ7IeYWBWPL
BQV12V0KIHw7I31EebDphIvuv0hlPDNmvSgAEV91r4GJnkNLoRNslVxpTR3FBtuI
kUlbzc5YGIlazFuahQbWKfhobkLVXc2Y0bqVqmAQ2c2GUjC0IlgGbMnugtp8YRw+
sGXh41hCnP2jKPqmMxMFgzVivbshsGuqenIg+chZVSNFZ2bqqP2z1FSwdyCXzptO
pt4F5clL+Bkbx04vxfD5xDp3lkF8EV64d/kcTk7yL9lFQb2BklreqnkOe7PT4SbV
l2rGrSn94qunuA+M+Z/flsObbn+LHEy3uEm1Fi7ZF4p1KDF+SRbYqhY60peAVsN7
shADUBSqntnrLzGWyHiVjqBvSUIDYFpWEXhMC62FpoGmGYH8051nUAyN9buJUACO
kEM0oS/4eU44NAhHUAU8ZA4bm3KoAFnl6duvzTQXKYMVmEjRK3q8myYoSs3Fy2NQ
ErYaq3siu/b+QIf1tA2dS8YDBhOV2A/jBJ6lQDaT2TneA9rkX5IhrJsIQe3S/xdo
2DGBh7149D6+KSs2IfHs9VLDbbSVBjLxj9vhzhE/GNvq+aCFEICwHebDrE7udugQ
M2LO3nqbhCZglLtxrBs5TjrUwdWMOGP13bsI6znX2+7vu3WWZGPc5UrrOyQJrP9q
TEBBwSJfFDxh/mJQqTBIv+qvekQ6OlNy7+A5fXJKaYASzB5HhrH4mECHdA6Dzk9u
LNHtBB1vqYj+VgDfCiUkXOBvrrhDxjWgyr3+yjgHUSYPNVejum0LCnqiX0n8MJsf
gBG6ZmtNHQPZ/WSsmKxHmUljgy9GBKm4g46ByYdAlWEX4QiZg9O1IJ691BVucF7Z
3y6yv8qdevAEEUNKqgFrDTg3ngPlXhZ6KKrhXm8P61MVnEHs864vcT5SEpFvwjO1
pgRsyBgNzqgfsxM5O4bZvWKqEQLk7uRc6JPtor315rqL+hg70M29NE5V4QbGqky5
1WJ9703NaEw0WVhhLYiR9sR6HOP7fsdW1fRO8JrJzThcCSeWiuCoDUw70m6NNxKO
1ZNpHySpQKXW7cMD+UTwyq1yhAOiaSfPO7AZ5+WUizojYQ5yeEBJXad3Emi/ZPru
dDVPrTqIrOI58kKVLMy5ATkv8s5c6hL+fRITbQqbEGlk1Iz7zTxx+3Q1teuBWEGK
02T9am/gn7PoHGpxwo0I4eTf1bRnIdIE5IDhFCY1K88sQGmCVo6fRrw1YogNu0Ax
boFCE0zLGof7YIlXNX4BQk/kyNZDs24m8telI5+v6z4qs5Oi4TtiUDEP5rVqn9/6
pU9MiBRTi9yMKOXCnDJwILXY/9hbt94cjVKcZSxo9flEL/mQIZk3qRvwmXXqYkfB
GrA5MeUJDZAtYVOJvesKJl3r2PyojIG2qRUd+MnaMuuxy+VY5sUform8mBrZu7hj
v29GJ6/KyyXxDQYn0O/XU3iU0DsIMXL9GSCuqwGK0ZKSLIi32PHLCdywNKZDKEpJ
4AgGOpzF+34kjzzoskVK23CDOuIs5+i3jxQpC8g0lSPtM235eqbAec+cdrvEMEeD
xjATOmAn0/X8Vi52L75PVZAmgwxNmMwNGfJI7pqG0dpAxDE5K5ZS0AuYeB991GWE
XAvAXoVOboNu6yBexA3IPt6vgRKVyiF2M0kLuWi8r0oSQyD/NruDpNEDqo3lAz9F
P71ientp/VE7AXw2uyF7O9iIIKFRweZqddfsZne59xsMD8Elb3Uod9ejAeLPOcN7
jBCqTUPjG41dnbWXqG+CsUp9mavYALQYtQMZhZKFsiPzb+QjfcZ33V4Rsh53la0Z
0o1rlDrd8CVy2HyDa796hYxIEznnnSR/GTD3igAjO3wAaPP7h/AofGADWJ1fqr+w
MD27FIzTz2gwDLpE0rOnrMh3Wgu1JN4NP6kE7+VpVLZIoh2u6WTZfamMPM/p5d1P
kXlsFoMoHX1Sxb7UUWhVxAD3hBMkSp6DxpS/KLITNwUymo8y0Z493zuGgmy3//IW
Yyagx8Q/F580XKrHNUNAOhvrF+vyrs1BGyl7epHQ+8Hu66G9djmtSlqPjXPDugv+
CtG5tEMH8LuHUFYsd3EYbbmG5d7FcR550Jvum7cHWNmDRrmPFNzZG7nZdwN5ddlt
RQeKsvsA+8h+kc+9uRyaCTncP/5G9bdkjHHr33yOuh0UzaAuHpXTJfzZMnc9KSs7
SsgC7SyhANLDT5mnMOfK4JBdvHrdusFLgQmwNIWsNUVKJK+GXGQ0Fe+Xk7aEFj9S
fICwd3kGiNhOADVQKY8+7sarPgOacwb+pbb7DpNLzLEQpckks6YgMbYvsYjJCdwP
Nae8qNuHE6DoCXwl3YO5Be6Wh8BQIAmMieyNTbu0PmfXHHj73mVQ1HQ1yTRFOd0v
5/JAxhA61H3PQZdIcmYUziRZCDKX2fZDoIyJNyUhgkl5VPHo2D1fveMbqae6tDm2
Sq5XyikQCilIhixhxyqNg9/BGF98SLIyJfLh68ngQ+/6EagWn3xMZNoipnZGXu7z
ZFcKTRhahC7zTJFq/r3xhkF3nTZ8FX6drv0IHwa8L5BMVQpvjGugVV3rD/eUGiwP
bQz4xiOq9OFVduWi0W01jok5OtxSesdySwjnsWMgJ7LvpN7u+qFEkTtbQESMHzy5
5H3DEWuFG0xW2zqAvsJOddZNRKlzTMOL9gNg3jiREECvx1j/23+z8J3aIzDUzabP
agdzUhsaoHyDbqpto1okM9quH13/kTfqltIkKlG9/fLQsqCICLNtKyigZN50lDUW
TZp5FMsHqYXZjNquTGPicUpAL4nCED218jbSgSghPDoMojmZVpXKlGi4MoW4eHC8
QWObKTIHVuTTFjteAxnF/B6+lTcU19H6fD29eEGIPW8mtVsiM1exhXoU+AMEqPdN
xMLY/i2ukYnDweEy0gqQSQeiy3aw/hD776hAAvyI3Mu/O98d8mRHt6bUx5jiwyjx
v2HSjCy4Sv5ujrAde3ouhmQ2HoCUD8sEduRmQHdG7KOUOYE28SfEByTWWu/8JnCI
oSwAJIKQoCE28z4FR2iI8d7sQB9uPQCw9SB9Ze4hgTwbCUaGPKsCuIv9joHH/TSI
SBgafXLm9AZkvvV6q6RJVY6k/CkRpX1QK8JGQQU3WzTo2ktz9b09hgw6Fj4V/DTs
PwQncXuCbUkUCFDTNKDYpeZZ+5dhdbZncuQeeo+qk4Bl2hmwUnWg5pDNghlpbBn/
c1+PVIOWQ7p8AryLs5fiHM2bEDx9pxSFOucI675CWl9LjIiDK0QEmpYHMNz20rZD
P3Qhu012Ua24FuE/9eC2C3s/umdQGRrVLBGer7FMdsIE0Bp8Jj5l98Ths9xXcPQy
bd61CV4BB8pXP2SIuX18+Se3wnrYLhN5BBwTlHIAKrVHzJu3SXarrV1ffSGWs+mV
clxKAGHwnTtKRLexwanvmK5r0sEoG1ea8/O0IyHAXiNQeV5mvGWSfXySiLuZmdlF
8QtoxXn7AnAy/fA0O7rhrAYMmKfuZNi2V14TY8LYmCn3pJiRsqLyxorw45rBp2uJ
NC86cJZrCfwfJj1/g3lPt51Q2Fh5dXYshWGBuuDM/MYiYo/yx5jbwKkqY1vtQpCn
5dgYUQz2F25pws7/4rv/u5Uf9o8uXVZTXDOWT5TJbp9D22NCTcX6oMWsmY6f6zXV
Xb04RqnduSzxGl41ScEz8abLkq4WJT/7kj/SlpRJCGJQvW8OMLH89Xui1fGY4IyO
HzOkKHtWJl5pgWwwKky/qJqmdVehaOT1+bQjH2Aty8imcKpgUIz/c58eOFwKnjzd
N+7tLakuV3deFUGyg4BL24UPvpP5YZuBjS4KelcFOW9FUlHkbSZYgDrDXO+S8OxY
o+spC2R/hXEsqeAwt0X3y4CJTMBNo387xxWhvl0MU5LZhRxH/6uKe5eWOunGTtv1
mx+8YfGqgnh8cpOw/LyCzR3gnP7L4a9x0dwfXKBpiX1Zr5oLPvWPJuLE3xfZ1HQb
kzwfjPiSKeJ5KDxJqzh+BMwFFHJLUoTNixnc3hhKHRuvfIgOzyJIZ/g2+j5uP7pV
SWXN5c+etMtQVDxCHT1Rp5Z+T0Xqy+RuUvOJ5Lsdslw/znR+GGKFHaQaRPxFV2A2
fpy2oDlGaXyi+nolm3pIIpeTLqWNwo6loDiC7OLOefm6tgt/b5gknDhgUfqb/CPf
RVBF/PrpWPzH9XCf4plF2GeC1ozjHOxUv4Ra/53nGUrE+ihnHwylQJnCM6QHwPLW
kPwObon9DccEQmklRsMzIHgPJ9S+uQCOQJaeedpOgHpvtYq1NRubcFkq8Bkx+Cf+
l+A6N/IH1fB9KRBcLlhp4E+804HplXwvhXL2XGvt1RasCGxeIz9zEFeq8aF5sCA5
wn1AqOhRcabsB3mofbKmEdCTUvMYtT8wRXzvx44L5jD/SkNjeSxIkGEPCxOgycGq
lHK3mreE+RxHxbnho2SfHvV2M0k550csK1lthLjRfzZq1tObZqm2Pl1T41ZKdvWL
QNt9YXZ+0FCx8sRHwXctkYLClYSbviv/FYwjQSBB4lw6BlTnyp0pWiyb5Hs5ozz3
4N3lVCE0horhUltlG+27uoG01kY97Qb1yiXNouAlTY9T+y5zCZ2DPDh1VX4tgPuy
C0jZUi0LNrX+MviwXwYeJlvKmo91g6aVQrhlxRhNidJgTTunkBvy/exbnIudfQJH
f41z28XsS0SkFpHFsiewb2AHo5Ztceqs20E94CE1QMJafmhDq8x1kgGHcUU8OhOZ
m/L3ExlCx2X6WKYZfDvhQqUqA6+fr1ImvTwOepOnrunpRjL1rQTM2YLq7QJxiFRv
iF//kxn1USDATKrOcDBGuc9PWDIt5pPKLZJoy/HcOcRMELDusrhN7w+XAeYelkdf
HW6XwCcvEHu/8DB1aupHMg6nvnPrOgK9PL2qXJcKOc9DTNJ4xEHP0iW6sxhB1Etv
IC70xnjDK6j08KWNj0Doia+o/9qd4oUJWop+X4lTtx0FT6DQMlj2r0eNO636UF+N
NixukAKwyy1T/nGaFR9JULzYuVWMpjfxmz0/gKhCaDZMoEDKwHqLrN328A94BB2J
PPvuiRLgzwWCzMqoTF1xu+fOtTAupfWvv3Z0caMg6sqVhvPnB1pH7PM/YSwaIxBV
le8guyJYjvPTlkEFYKAxb0nRj2n/YJWr8V6V1EUWQ0IopTIFfQEzIr0osVBtuQB9
uk7co24LE+mSfv4y2TVi8Y6CLkdPDeFPXoJTwORsgI+0xlmfdowMNyUd3V8pqjES
NJrX5IIdhlb2fgiV7R6dDvtGsX05RuXFJZTdjpwn0MXnqnzbn9UNLodhch7BPmS5
TEFEa0fFvkrQLbGzHInUrDnpHO9K8AdqTy29h/RjK6cZtTIiOxZ/PJBFxtvsOsmc
X1itxvX6I5GNk5G8nt37lSeE2ftr0nVMQFY95WX6XPBXgFtdqMxJAHlXc9FRjIJB
NrwvZ/DnVZY69038Il99qj+UVjL0YZ21iXxCefJEzQUxqhJLWQIe49vixCfQEHZc
iFnd+S4CZ2rmxcD6CRPKZd+Vo0XkGj2SIqaNFGW0+3ABqbM5vMRM47l2coU3uxny
7ypxFM0dvC0Ttoupbi9HEAQgt4z8uTEIBKKNysyjaWU+Yloa+mnuGdQ+OVMEfxzb
/DTOB6fLjnX/7yT4la4exSlGXZAa/OhDZV0MpUYZmiVR7q2Q5+mLoKdoBTPUjuFc
eLvJPuViZjxr3BT6ctFFA4UJAPKOsxwCX+fAjWQyd9c3IXgM9y3+2Tic4OFAVNHx
GBcJbuTwUNUTX9ndW9I7nrEbtRJlgCY6HAAkFOUD4yJfWEyhYm1AN/qYAFH8xJJJ
tIA7S+iPABE3CDnQUuQwkeYKLgKsTndPdEPnumzNnKT9RF0JniHfwpElgOmu/PqH
syNYzJ0tUCW94lohOlOHELqvJhYc76CbnkC3t2j3spMB9QuVPuSYlz/gI3JTS3m4
q7qACjpsQJDCbOUwGloRrIrNWzLpKDmWkDtkKeUwXWphth3yLCF78mhUscsNPP0B
9uErepniunBHxG+aSIGMBP5bXzOoSZ3VG0zBevV4tUMALKNmRkUthS5vgWs6fA+Z
M3m88rBrkkNkgUPBdqizIv9fh69fnGYAihyNmoVuTsf3aCqgAsjHXYiXWJwXezQ4
uE0ydcFvKVygk/EN9ule7fHLft3fiVicAIvb4Mq1HL5/lq5HyWFpV76Y/HpIdjBD
ZYva2G4QQ95n1auq5ua4lOFNbMOgvMv/JnF7geYHF3Eo2J0C4vI7YW6Tjrh8Iva7
3O1P0Aoj/LamudQO7uztWV13/vIpo24jum5GYYSslahTloeIqkPNlB+4px/DiYOf
jF8JSeNrWQd5k+i47dzj9kbfgWZZrObm8cia8htNUYMRIEOs+SD90zQDvO3omXIM
yjYX2AZ5/Q2TgQntlW54z2g9cpHerMIrUVV7V+6bqfjoIM6Lv2qH1v1h36qqNtth
QR3OesJ1BIMr2BxKcRgQ3ZoUARHHIuLQy7nmER6IeXGzMJY1AqzH/kMAe9tltQdz
B/fjRGdNDR4qY8wcrcEEvncMFx8mJDsJnd1iLGEpwDQFw1hNHj5OcyT1hpmrCG3Y
bQdvplUOKVxBkSF3LODNi5AOMlXbSZHapElF3Bvh3wJiq5xFHeolU27rIcZ+9/2V
qLR7zNu5PJil5tntECnqrxY3vRe3AyY9SRiN0uTf+RJ5RS9Zi0/WG7QkKU/kHOvh
/jxQYI/ljz7eYBs4/1SYNiiRxXHlL8V3/bdxu1EeYpFEkrBBnl0n+vv1ubMqFWuU
Ak4OD4YPBWrfYv7qGh5A1aEvZRrchOH6NAm/t2vHiRaFtnBVXGqQnmByR6AdwcUO
daXRwIHFqcug4Sm9N297ok8N2wIXdxy901jMvOWFRzorh8VspDSel9RHAMrXlfPT
23kKxts2RRg+am/x9ATkjOhFUQzU2ioRZajzKMGhV6cA52KRO7Os2HnDZeNSbpW6
UZyo/nGaUzS1hyk/hmgnpfKe9JobHr45OirSV5BiVklUVdRNsznINxL5eYxNbnPX
CONRvnX0yLr7ScwaDmaQVAQGf4+1nWSRl+wJea4Gq77sKcNpkpgDaP4iXZ0yMl2Z
Jv8CM/CsnAXv/rnth2xbRn59R3uKW+3R3d5ovDWZfrsdsLqfsRZDVyRTc+Z6QvDK
GFvwvv4vYDtAObbLmkl9RUN8MgNVIlEPJR+x5sLsiZnR96qMy+KisfyPooQBkzlP
hkdRUzEjZhXt22n81ra9dHbe/C/VRC+W7QS8zB4Pzkj4Fumaht4WHF7AoTuy49qY
U6zAtyxn3/piVwqJgfiIY+Ykir29Jw9fNgYKHu6ixpTSRniMM8BFmpv1AyCHNScn
1WmyjjVPgQDc0Ie91RUNSOakm5jeD6k0O+2PbDSWG/bf2qa3RwWVoR8OAJj0IEeV
Yhw3c4RMb29S6Sg3Mu5esDeII04z5EP8QjI+XfsLody6+gnIwM8UvnYDrxk0lPER
gjQLpVODG1sJBkKo5YYA/6oC75eZw3io7h5N5MMqoBlSe38IWDEfyYc9U03uL/kk
GAbTZX+/DESNDFnD25spFbyOQ/WducLrCZBKgrYPsLmwZzaEgOCfG16YEnVFOP1m
14hctTbQ/OmtqInCpZMlb5l+5035fVmq043+U3N0HGWDyl3IBJqUsEXNloj16B6L
uRZyc3xOZEc30gZkO5UE3Zmif/hvbs/+7wsOgZpjHu41aRRh6DLqK3nkRMd7D/Kv
FjaWw/3cOyzA+JOSsg49xUHrtbX0f9yaXLAkxBfH0+tqnmvG0V8gnGsMGV1MswQT
pYj4oT2UPu9Pef5BoeWD0TWb0/hxDZN1F8CCljluViEb/kbcUl15OTQdLHheDaia
hnNfB8W8DTklr7JoHs3PjcescAl8kV67VthA64/Z/I5R6VEPhdJKav2b8PzFFbfn
3/2WhGrgMaZAi2E0pBkO7hQR96iCRQAHiunyWMKU0FKynTntYmvQZyN+kgtmA2mz
9uOuvICy7zMHfHxU3SEMrT2tDqDZihWMHfvkVfm9x/0T1mWcvc04djExMpbhVfMH
oztWaIXc81hR3hPULw9LqBYNom58nOy3O0m9JZgdlqYkcdzhTeA0cT2VYPnQ9B5i
H9iULTtJuubSSALw4zDnV7o9Nw/koqveRyQuvpu29q6LSRKjATPlM+HchU1/O3ub
doBLDGfw5xa+VnBl1m+n+lh0UlfLjJjc/S+HAS6VgecywogGP14iH4yR6pOSWGAA
F4Ju21S2LyB36ddNaa/LXOld3OQTE0P0ylXyZpFlIciY2QA2O6Y91cDIgAdfSHcH
Ct7pw+n/ugKkvYhUvqtPZnZvJOBvOAvBi9wnecy0Ucyby5FYi8UxvL8VQHE/PDM3
JtBG8KMsgABIcRYAaOimmPUMin5k8zwVkdAvByArviSXKuusmPHMJq6WAEMIunKc
NJh3Wm5pa3/uDf1A0Tci13k019SYXimx4eSuPvtH0xuBk3FAD9d+XOuqRm/J91/S
jULDiIoVPL+v8tZN6WMteMbT2gxR39JZs4Mfe3S/sI9h8eDaiXbdQB2XxKhGvR+Q
6BQrHWHSlsdhPtRXnKVnpF+yFvoL4xefZ9y7WY4XZZSlu9nx1Cy9fo04oh8RszhN
xB/Hjud7fhhOSFj5V2aP+mXfdezV6D9Bu/GsmydRJYV4gZ7KewN3MoyRwXJ0kytw
qacGPgEJC/2uEuO9c7F2TihLvT/X4mHi5oVWqzZv2BNVTo7lpSI1Zd0aTDYwK42b
ESU8WL7xn3CxaUDxJ/djgCL4aIcJJGAvJ1AMjUNmDDfg9ApYedcyQLDtejWZQEBT
Ja4jo57mckOttg5PeT855OEb/aGs4uiFk95rO5PFvaEVu1FofIpFqa8g0oak5Iwv
q89TeyTiRGkPEL1BSH+MTGY7r1waHdjP6IS4RUHfL6dfJw/loNguNm/l4Bt+3t88
RTtHhkXy4v0SxF2khndVxedWQA69eybus8UmHc6iN4dTdqbvlvsjIai/IjsoylJi
SIpv10J5kewdMgohpR5WX30q+Pg6XQaQ/W5+tPDCIqqVuUMGCpyvGhpQU2NTVtOp
hfSC02T9PLQ9uZ2vv0sU3vJQ1Z+fBDq2tBB9FAG1lGyo/UN0w81QOMAPXf6oVg6j
49nFdjR/H9PhHIQiISw4WIv/vSL7yiB4Rs21PTBjdNLfeLOQloNjKRD/IMa/D0tU
VgS1fwbw4k1eYZn9omICX7KEqY1a2O8KMapGUd+LZqkKlsDCV/F1sOO8i0NqANee
CvmXs6HdhSeQoc5XAixh+UDAvmiVkYqo8OPB/Q6/TUM5zzCC0IUMjaqMGM7xKq27
nRZiO9NcdR+GrIPkD8BSbIL9dx60pIZh5MP/DBfyflZPWeBuF7YdvRKEP1JJC/I9
pZ8kMLTZMGbz2lg0m0IAgDpGLH1jGgrveGSK78e1jT462ztixCI2sMbvL8lwWBWx
HGPBjt5u6Xc2YY6q0fTz0169ARQqdEmpSUY8pEiFNyNJfoAdmyBH1N4spbXW4IVr
KN8XQO65Phsrjc/9BHjk0fCBEdkgxOagaG8asHeQCACkqwr4FOiMdjXmX8wwdUB2
xMeB5ySBtnyqygmJ2ZiFrp7KvOXXaA14po9Qf1VfxYQ4Pm6xzOxpZ1x1kYfuOI6v
sjDMZuXsLso3txM0p4/9d+jQsD5oCRm8lqUXpIKoSia1whiVCm95aBDTDYTvxIoJ
mQONAOhc7EpahHQ2JQWvf8Of8buMRdFGA0Ql62QduzfRP2PTQa1XXbACQzz92CQe
Hhm/YxADaQo4uvQQaZTPwohPS0Yq4h6HFtFQFXLyZZZgY5KRBWVwQlKOss71U3Dx
3uM0f1WZGxUugEtk+8Pw6qhasf5/a5C3bsRU/rniTDCXAWLzjAnhFa5h45FrL2IE
Wcdmp2UxpU+6evX4+QdtMk43e5Xs4dGv5nYX/cjzr2GieFyTAAkXFh1m1J4/4z3s
wfR2t/iLccpADR0d5rzTYeNIg8MjZYMBdfZiO4ZamW1x+vVfFcuJhnj6kueiOnne
Zl9dY0hh2nr6hIESm1Q3sfHwOdMdbM9zVXejLDXfPKVy4slqEdjeuT9SxV6Sdyxn
JNHtp7xv/K4IbC/LDC40a5Ltc/so5jZZBCsfiPjXp/XgcPb4ZL38QqNX2S9C7kvo
tn5ipD9x33CjjDdjKokR3Jc8TfYq7wt8MD/8VEi51fKkkecdBFbpLHJw5mUNoEg8
5fb0MQR1cFMni18nFsQC4HDJtM5ZO+iMe7gF753YqTvDwCEhRSpAsIiC1aYGPvRY
ofKZ3wY/YL0qwr3gGNfSPT7hfsiHmCeGmcgXAC/OKBpvsnhc22RTNoCe2rNzqYwN
JBuf4LMDMwtkj7kVaBaUEP2kKRTzwEQg54+wNrFvxTtAvhuewTvDbkLenaXckkm+
DykwyNaadj3A5nNoc5SW0Z4HMIbFKlwgIKYbmlmlwpL0g4pgpatZ4klMziZgrAXc
VXpy1AEwLrcwRTBFig9UhEIpmJi2hogekxPZO0P/rImxJLefqfXt9G4d8qupyI6K
bZAN4uy9kOSSXD8BuvxkZSBAJ19U7O5kQ/mKF7BdIHUx3Yar9vLU75KqbXBoWRUq
FHoVD+O0jY/5WmJIX4mZb9th3k/R8L1VU9YyImFykF86mFQQD8jqPabY9kV0M5wJ
Bp0NHxZFmMAJrgR8Qjiogn26bS3vHboM+XzrkaGQumwMex5hI7scv0c43KasIo2m
xMynwTSiT7oVDKQopZ1tu/eVwPap64HxwQRhS1DiTN3MDSMX85dsOYi4d3p8BgOH
ewjUhF574MN31+6uBEqiRaR0SELwm2F38I5Qo6Q2NiPKuJRqhI+GIzF/jRc+Aqfy
hlgIYdcyHvJTmiMrx+uxe5k1SKibV+Yi3gMtp5VgFAaF0Qjm5aTxoVEx42a4Q0tq
pkXBXH2C/x7vLFrArL9uqOwb6/93u5h71zHbA8uQkqqrnudnb2bG83YXmcMDqdbm
+0WX6679ziIONLkZDQCAsE4+nCiMjQcIiBOf2Vl/r9eCTjgwtkR/OlyYlF65pEEv
6Iv8bcwx1sk+Je5fnXc0Rg8D8IIJf5+zMH4vvmmY2HBWvAYskQrwvtRSHMIqHVsR
EL/L2zi/DGz/1ecIVAgDnfuZlfXMb+I/EgYwYNbY1QbeyYlMGgkocMjrCCJ9gKMK
XBVxHtHankbxMzEj94LyqR9uoeTIsp1AYLaLmjRA4Rp5Pe9uP4LZna3guEgSedHq
7zsPI0arQMnZ0bu7OrVVodP9XeEcny0r74XwM00MaIUZG01plZuWaNWDkzVaRsxM
KAhMGNgd8MWbZwP0UqFbqvcHteX7olNqR2hcDIQgtnZsPN3pVzDCy/LfBKmvmm0u
Y+Rgoks8VhLj7VuC7hoyQmZzjnkxQcqSWhq3I/5lpaPO0W9LXsFTky9jcWdjvpCf
bPXJHwhNEz6Mg/kV5tQH/syU5GVr6tbZjhyiC9XKzLma2gDqg6f2Cvnwl70zOz2L
g0HUUwKkbt/iYijv1MdltnC9R+jHf7hBxNjZ5Y8uQ0lECJ8uoyzFzE5WoPmBtJSd
3K7x4iSRk1CDuSdcz/pLX2V+zVrGlHjDENTF2bF/VlBzN0+C+gVdASYwJLXNhC0F
ZGRTYpbkJIG5kmvs4A7Nb2CvJJ8Jbx2NUv9jrOn2xsCbw5ymvAuU8AOnTRePr5CH
QFNuVFr77ecOBnEPBT11BvuSYcVgPaPzQAWmtqgbW3xeAmYsSY7z9n4OSPTXWYmo
dCZzeHpj7zlO2dKl5K2ePewAuyMGxgW3Oev3noY7UYOqEkqgnwFssESqTVNKi8Tt
oYEQ9hmsf4pmKlSBm1w+9iV1YfwJGVFZvbAXlIh0s4keMTq/DvVWrFgA6aP2UEoi
2xCbpoZMYvMYwotUICqUZZnVLLclvXbQFsF9ls79JJbVUIHVFBYV7RvqkDwveuH3
yqjF7PnsFI9hbp6UcemKGJ7s01A+G9cqOB1uperBGImimPEAQ5PMMvCRgl1pkOP5
WQuqCHJ5Wv4GKwMAFNmcVUVHjsRVz146+2yK88xwMtYLitfz8YkpLV6Nsiwt42DX
XTyXu2+6ufx5ljqPZCpGRWTVCDJ7OzF6tyRTl6igPtsPU1iFKytESbk+xn+68qSM
QcBxpkKdP+m5BOFGfFtgZzpCMGAZfGFF3ofe6v1ffyzL5qjqE29xjIPOOmikJ/Jd
HXvZet7nnWrpUSNuueRtEJCkSESJiJAkRiXms4BL18rNAlvHYfaWdHcDGF8l5wp6
ujvy5a7f94wv4hPpNUM/cX85mMbss6diDZfh/7TD/JNwWPJHDddVhwWXuerJAMiH
ck9JCZHPJ/WU/olqHJcJt54IpipzQ9dj1VSQqHY/xgYN9Md3b+xISNmEx+kLynu3
xC8xNg1a51yUSU4B1Mn8XUJiJWAGwmHr2w/FRogXywZGYlgVQOTYameQPM0b4UrJ
giI+tCZ9zj1A7qpFbzY3J4hmee398a/JsZSNTLG0rydW+J9ApxuuwELivG0/TV+b
NBWZ3bDbHRrNZgYfZExfRuQQq7I9PHGZP8W5VQAL0wFcjaiiAkEi+AOv3Tq2SCgQ
ulsjsVYnIpv747cDJMnuH9sNq81F/hfnrx4+ADIbiLxJAgkU1pDbmFylRG4vfIdK
vyY/DlA1d48S46cXS0CvOonCfK0l4nQsRgxoZbzLpJ7DBxsMAXKxpGozyq8zKzEL
huYMp00kK2eXsgRzH+Sm2/uhu2b09wDzRbtuj9LSmGIMd/1WqXRU6ra0DJP6zwnX
NopSCw1HBhv6FtF8OedJHWI7gsdqVkTuDXSU2BCYn0H2j8nuX/mqdcSCp6CzqXuN
yaF+SnAB6fdosDXGZyil84WUvWZE0M9nehFrQQdgFV37efOJlCAyS07qYwMjLo+L
bBL3SUHMb0UzpMv0wbpbWT9H9eM2drtTimxNUVV/5NyHj6Z7fMJrLSdLPyk2RbSX
Pdmb30Pzz06AlPzyilB+q1c+5yDj77ZPUHURTdO7hHmN4n9juf1cE3Oy3MHTnsXE
FmVIpqRsChiDMINs2sUhbYuTdcuWHBPWLEPc9zpSlfQkJck23Jza7QnFxa8gbcQa
3KiFCvseZ4eQ74G3LU4ErhDd4MwDzznYsubFcBYbnMDs1MdpIVg7CgjwiVsz08+5
JgC66zXB3bPC/9MCfcc4GYFMRvla7CzU4hlJBUwdxrUpnUh+SaM29z7ugE8a7j3G
4nf8+tbNcjqz3tU84aTGVb0eYc4BQM43nIRGpbS3uZAMTp9ZHzUQ9Z/snCEBxdH1
UqsY4xRfFcaSIl9vSVLVY2oZ3k7A7jUGa+kgTolajGwSxXq1n1QsUnIb44TjJ/20
f5YdYpauukpdPX2lJjYnm0a92sCZh6lrdqVEw6WV199SfRXo9c0h7Dt+1SoYsREj
5Vus49Wcua9/PqmS3YPGMI5MFGQv2n0k/0+yoFuOcHIQiZeCwQQTujnI7Z/4rkh4
+mIztIZgaSJ6K4J9QrkHe78hMG3+/6nE+nSkRs9qbe/8+u+f60UTkIJqpXxYs22+
+wQq7u7CkO8hjUZoMzxPXrmQ25PMYqZE4Pv2VU/1aX7AHbQ5I3/mG0n5BDTqimJ/
lsoz6ohqm+UL/5yrdE9lMmH5sxM+wDzARcFRul0p3una7UNXpDExYMdPQ+UF4Yuw
VTZKZhln26nGXzbaPtTDD5J6MbcNK7F61q+lrJjZBH+ZQUgiBmRrhZsCSmiHEZdg
6D3VHBsBDaABfccAiAZwfegEFk2opU3sxkcYILPa09J/K07PIzLbKUy4tlxkOAPD
az/4EwemYPKTkTkHCRdiG/PELXRlp5DkoX6uPLmATivwVMGpmXInppnJ0JyExLWH
/VO3L7xgrnS41rbOGe3giOAlYrawJxoAp46umHaeYKgVWkeELZefytLKMIx4fUvv
tIVO+m+Xd8c2WPe2JiNykPF7/vT+yWHldU66okV3v0JcSwP6uqaq1TJ7GOYQRSAF
LtHOjpqzPGYOFKM8fJzMLXUsnd+SVBIDwsfZkQUh6pJ7wvWk9kI+KwEiASQGjH/A
0ri8QR63lG8HpLbs9WFruabfV6VmYkjdwimyDvl1oh925448oyg21i6vDWOzgMoS
14OmsIaxci6921RLdJpXaPI59i6/zjvt4/hCvyJOKZ42DKRl16Ae4p/WGf3RMQZ0
5jVucwyUnd95Sx6sSqW17jATr7s1SNm3iBd8ZK+v2b7k57OENgq3U80WxG4qncmi
D8hk468AoVSNC0BoNWRoLtQy4V/O5pLiQGZVTV8I5O0WSONTpxkNFT8qi5Zmi8cj
m8UFEti8DE61gJy98Sao3nH9NNBMY7XXPGa4ooMqGCMzyNM89tjhW9tvxJwcFQZu
y7vlITf8I+cqibE76t3pz1URt4D4LaDEtIf9lojzznQzQa1u76Eg8FT06ODlzjWA
5Zmuhy6RiGpL0nllv3BoC1QwTOLFxamaV1V7zL2kOTpRvDuDJwkIRU+S0ptOyiRP
LX6/WElz+xr1wLcK8rKo3c3nuqt4lEBCQWuvSbOzz3G4VDGQz6bHxU2XOTxJPAk1
A59/h/UK1UYYr0XnZzXrcecr/hZ5+ziIy7eoITpKF1QIMG7rrVQXB6KdybU8qBOc
pBCDGvegCDb4W7vF8kgbkAoh/hxAUsID5tmYaRYr+4qFMKCT9NNE1Eqi30BL6buU
RS5lqtDGfPeyEAbBWBnme3qm3lX66sjEgUd8l68afESall05gW64biKDmMsv3O5x
KCy1eoykpXmGUlvdJzyIbfXiRw8R+TmtL3haccgyI0hgOO0PRuMHYy+uGsa25zVf
g4Jx6fMJjBAlDBAz+BGRv5R62j2aJelklZ3ajVvfY/UljmUDlgx3Ekmyvb11BEvq
VklpfLw1vxJudcV0V1W7o6h1LHTeiUeUMDjgrjv7g1RoMkDSBY+C/ELXzKx44eOM
f03GHj5t+xlPR3N5U3MvTfOqWyoMlx1LgGIUVBzsEM7vvspFM3SwOT5NCc4oxAy/
q7slUK318M96x8SC5p9qVyqaekRvG3OMwoJu3nId+hkQfaCwcBdpbxyE5XXuMV1G
N+KjtQZh5WHkCr72SKf0UJqXTger6cPn/HkkAPYVjOiJCQtk2g+Z0x4Z+Ad1a76k
kw3+aXHOd3GGTU7WttxRv5RhLxrKkbiMT0rQcchiYseDRidSCbL3khTO6BacnnTr
8LI2xQb9vrh/VcgQl5NS41FeTzeESLwZozPZ5r3W3qht62S1fPtUwJeOaDEn4wDn
7jwEOSHJh5ZqkjtvCHvqmo3SAzP+zeWlJpVSlRRCqVP5cw+4gq4vUX+kjNwGctSo
mQC128tHudIFk+wG/aDsV/cC4R2cl4YCmwPLIrzxa4jaAkBWT39N9+FO/T1Qa5qO
71IaGIA9QOBhqu07a8jLrpKfqy5rR8QUYTBIgEjZs+dQWKCxKL6tY4e8LJXbefrO
SC/LZS7BgDJBkei9/+ELO9LYVhUSvdVwQU177Xyde+GN4Uy8LzqzqA+ddjVxK5wk
NE85hDgw9kK/c3rT9+oxNFHr4kZDY7sNHu9rvT5fNEiUxqCau4zHMZwA/mDZHtS5
OALnUbJ9WVJL6qK9srVCzRWRwNhJlRevhtkC6kfxY493NMJX2j6RQ88ahANlvOCq
rqG//Nu+bnwjrq1+ntw05zn2irrMJtpPN+FIyyq4GRV9J6s2WqNjs15HOjrzZJBu
iVh3Am4n9FZQdLZwC5k9HWb8xys84+uqZXt4orJWs5TF7P1EwN8J0B3i2AnjPhuP
XW76YqpX2qGDAYsZvrcpt6Z+yIy+88+RBDao4zQsvvdKmaNkqKxFDPhJ5pOrX+bD
Fh5daSYOxRN0ucy6CC3xRiazP7v88Uq8Sot9M690eOmSCpdbqBSr7vAXuLsyRNYd
EZOWtp3S6OEYR7YIt9lgxRBM4EWJDEohS9Rk3e7eCSgBf+1ARp9mG2NBQpAG3YSZ
qDVXvJsvRedJ48PW5HtniHkG26yEACrdX0YY4RUPbUgc3CRcRQRzNvk8t9LD7l6j
xn7EcaSSJ348/M1OdbwWMNHTrvUeIBprLdW8Qgrf1FS7UAcjJRN0iAKYz8SEzrMA
tdGs3jJLFgnzG059yPFlEHstw4zKZem8KIFIRZPHauT5pxzV0A+EEQ7Yy6yW10V9
1uP1iCfAbfSLmaIZc+RHkQ==
`pragma protect end_protected
