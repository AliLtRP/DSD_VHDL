// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:18 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HaR8VysU1RcRSZGALuRO663+lRUdKtUWbXzmh+cDpD/PGLhRdACDD8D9vfa6C7yK
d3CxWNpox0geMSr4jWXT7TVAEOXiuGVLqalct6mz091msuRmv8+MCObbXtnR1QAZ
0Rr7MZZ5uSAtBhhMa0d8hwAN9UIr9LrpD0DtNqiKKTs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14288)
E76KdxvzKflr20Mvb9hrJBjbeFTrV6FmamRdLCHH/+/sHtzSgrN5zcaJxwMSjf3j
9VB4Iy0zek1u6udsUB/jjYzKFFmZ8Uyl/OU42pJ2zoK0At5oMZuzjbPLQRFRL3BX
Y5HeKEMzPu4qGngH1IaucN0VM+zQtR/9MsEnXIVy3J068zI/SlmTZ8Z/hjRHhqoP
Ppekbgzg8PtZW2a0kHKk6fqCma0uSocFrl8Igm4P39USJJTOcQEQGVRZHqUeAzgh
EyVmhqR/8Acql84VRApLMSvQaY9NVXORXPJuE8PHatoMyx9t8e8s5xVG32QBB77B
dOfK4l8aflus5ZIMXyPA8ZvS7hmL3TRPRl1/PtFB5L66Ura+HoPudfzftXJrvxXe
1VFZSQNk3scn3bsNd9NgWEpbpFVoFsRnOz/PdI81F2e8evg/iFYbYk2NGEl0bo8f
4Y9dQSwwwHWX7ZU5M/XM2TQBPKniOfbtygifDsiqmvlIk1SgQdGqtjwW6vtVGrgv
wQS9BQTk5Img21o1NYPb2Pq1SE+RnWYYG/4TdtnAwxZ+pqrzAm9J62Le7yfnMoID
AjTR3FSnSRRp8Hl7CdR7VtivurRioJqjoSJvNuJya29897AZ5umlAPFAajq/GMs0
giMc8zf6qKXkrdG2AOqu4iKRGiULGapCU0BcQgYuR3Z3hDdbt5jrRc3SlzA8NgL9
D0vgtZW0xvDUZc56nkrtkfdNiKuMkW43+BGMGXww1rb0XV/kYt8oypTFLzslD2ni
qIGTdWb/daPblq5HKvKpQokng2KsdKnJktuFBevhWAyP7yZfd8lQpEh8vlEGLo4x
7GF+prdVXaUKUWVzL5VcQ1nUyP56CK6/NHgTpoWiXKA0ZJ/kM+x2JyikL2OIDMT+
1vqu7DOHCPXWHWfbC3aOvRTgbLZozJz4mzL5FaWHcJlZXmkMtGaqwXrgghyOt6R5
bqkVn1GAfz+rMoT5OKRe0JK9Bv0ZgSW+Azgc6hk4XDu7wOGzaDLcbrUAvvAnU1hx
u4gi6kyEKD6te7ZjLOuq/AzuAQP9jhAVoSXhrcOxLwIl1lTWyzwyMyDwAFFEWN8i
nHRuFl+FyQI/6gXJg+1hH1ruZE6EsuE3PaxI9I+yC1zU70SOLoT54to5mwv/R86w
dhRUdU0YbIx/BY8pPSLbKXqfgcjIKDerQttTbaGxspdfE4BvYB5t/kIS+VrpnB7k
XzhSIyEfSBxQKIOgfiy/LPPRQHPKuUS/9yZwy+ceSinH92cgyLb7QEk6xNPm42sO
7SsGDO3CysMaTI9o97b73LCnc6EluS391mfJyD98qG6/16h7oq41WO5V+Z5hnMqG
WdpL9GHOh7ri9jY9nOsAuzpYQ6VvxVwK6aM60nDR7TUt17UHZegdhx1KLzl5GE8D
t1eVfdXYDB+nAmFDq+gRTxyObB1PIrkpe/oKNecC6eV1y4IXdFUE5GtJzLdpAXD0
lUjcRCOYO+fbLGrop5MYBojRmGsRg0cByQI1YqriptPHVu55fZQ6S35/nh/mi6ig
zm/YBHaMDN+Pe+ryfLkenWYKvChs70jrNW4vpQVK/gWYWKhJ6VNaRNNah2+NjU89
l8IrNXdzSBzHsa1xJ04AaqXqfQYpaThAMpESpyiDOu6RlHV7RP+jcOjQwePKNW0p
ifoOUJMZZc2SPX/xziEY41eJ1CUY21VUPZrKyuPuBM3DAguSdMzTYFf0IDJPV3X/
S41BzX0m3AQ/mGRkVDS13+g4ApzHHoQddqWtCtI0lPQ8xEi48FYBZFBRoD+7j78g
8tmjIRF2YQHzBmLTUY9/RTXLNjHVQvQf1xXSftz+9Af4ePBTB1pCkarKnye4gdA0
USRpAIp5ejdbjq6+5vfVKW2EECdpnzOqrL6P1lAhxflBeBWnGs9iD143gXBH5pc4
lLh+C2eaWAFR37kYg1CMMjFV4raxwEE4j7BXeVV+3dOXTsuMiy7gtzxmpf9+vwRW
eTaW690RTHErjVy0S0zQ8FW3t7rmn0LATUyQ2rjf4fPsqAflt45cFBe2mrCDvf6G
rUa9XY18kNNZxrtHDS0aBYvqX/1dEdYDZguavLtsljwbTz0w+IRVe0GgF+MnkoEl
FfrrecqJNQWq/88TcUqngnTz0ylqnsGKymd3aKYvQXs4q5MrRJM5AuiV2WlyIWjJ
P2bpacm0Y094RuH2k3X1j95UY3BcNrFUm/qqSCEPqp5tvRXixMZ8HWjsfjamL5oA
yNTkwAuEFF4dDR7ECtDMKRf8rsvhuL1UJJRKRGIEP0MUvFQ/j59bIa47CsC3Ig+s
7eAgVCAmRPIWw0yE8y+nEzvaKwAnxeR7UefSZH0IbRfuGlDJCXr/n920HpoU5Csb
qw3ujZd12EmRMzRM8lloHtLzxn4qZlO8/11+c+0YB1B2ZEo9tqOqtRWxbH53+7T/
EsfJSmIPbHLGhsKYYZm6Ea9gwR/UTrcaIgCWUxGV+JVz1KNXZqih296gEs33oeGW
njwKSpikyqG/tJqq/Vo5aQa6il7SEG0zlga4OEYvbpHa6Sy0ZPtSqBZwKlUVb1ga
U4veCII4f/m/kpdOxuNV5bpjMhbVk0yoJUJgZv4TzHAjdVTp+chZW04nCsV5afa2
ot4HGAXK6gVQ+QDg7oI6KjVRlF1RxDmaSV63aVADqapITypVzU9hnYuZg9eyCPhB
jZVW1I0PVnlePePD1qVnP9539BCMLC6hwneyTg8sxDDaEdmjYy2IaHM2TibATGBK
Qokr1e74SZhXrpE0v/uWhYNC/ETiJRg3SKah20Or2aDde23lRW5kKsW5NJlaICGn
EmmEqKM2I/2kpaNy3nzAHR1ceH3/ts9d5snsqq/4YN2LT3peNTEliMxMeQSa2nNv
IGeoZtJFTfoCks2mlQFZqOMdqn4ERZqWblOSKu4nZin6fFuuMiBNWV/Vh679nUlu
fSAS5Lw6KywBpas/kLoVXpfmWB/kqPzgLBi631Z8r/XCzWufGc8oTst7DQh0s4CI
OzTW0m+FvzslxSaJvxxmXl+o8mQ9X5tzvijOdP0q4pp6TxUCmU7pFTjZbOCerexi
P0KomVCVprgONj/m4ZNDmuU/5DLf8DWgBG7I65wgp+TdufINC3ELnkZEbnXVqMqw
e5BqwKR0bSq+7dAh30B7SC9ERdmmHBEK+64k4uoi47oYc76SeLjUoBvl/N2ZT9Fu
2x1CeKe2ry0zKV6pg6NaWo4EYdKEB4Y0onOS4/wN/Eg02z0Uo3XmXQB/ZCE4vCmv
PpIqGDWaLW7NpM5r76MfR2buik0XrftFLVzTGWZO2gDn0xWCuvaBU9VBMZNfIrRC
bdWDt9d3K8ncu0WQUNvQj/xEb1u9yNrjflVal1cYh5H55VYV13r0xJTAPRBJDHuo
J1o6QlvLCKQKALzLooL1p215p1jouynT7H6IilDAdyyOITu9H/GMA0qUimbFx0xp
2BAuFHOGlOf+68FOhIdJpz04xFjHKq3wR3ZOu8dTRG8lvTCz+qvOtwZBsoKpr8VB
rll+ooMjVPS0bjPxfZf09P9d6Q+9LNfl390HFhhZzjrMcWJ6wuExA8vyZLft33BI
RxZYZ6C+Uiotlo3I9q9vbVKG2XflMXw3kXcqm4eMCtMRZdKHZMgT++5OYMYo+Yfg
Hy8uFJ+2+4zH1qKnSA/PXS+2tmVESAu3lY6UN4NCEq2lsm7yCq43gTPkbDT/nZBN
Jf0nXTl3C7RIV4xyKEEqpayx/MRmfljAeb4iLug3eTvpYz5TXf+cE2ErlahDys3Y
nFYT5Z1L60WR4xfh9zlZ9xwMcLULze5OuFyROv9/uhT67xYZ0FAfbaJi5ZpEbrz7
Yoecnh6/NI4diaTPEk3QRzWNyayGJuK4LhDbWhshvFZIUgKHkRY1wgKvrTSIv2Ve
gsIh84PnBadcIcMtYCyjKeV8YsZ/PNCBPn7/ASdvpuD/2ck0vwk7IZFquGg+8UGs
uSACE9WzrlLjiY1uGmY+yhtiXF15nabtTkIUlwfNXcCjyDDOzlPL8rGy1PoVb/CB
kCxEwWh4KWqEEOA4MLLyD9N2I1Bs/CNa1L59qDvINBwOMgtWg7aVPZ3BAwLaZd+z
SIwbqQLZH2puaKz5QHyyu4UdbUwCRwUpJiSc6TZsh6XDVmZrY/fixbJqSvAlXWE7
AQpg8BjyVuNxalmU8e+wH+5PyLC1bgFvniZxCINrV0TIpQYlh/2dWNO9K6+pquTM
4ExBR9IRDB+VpHd20KZGZarCi+Wf/kcV9jM0KnJ27nTDC2i8bWRq/2xtDDlO10o9
z0Y31E+ajqyoBuhoMQlt3CbgftNTImbGLHVZ4lh9GMFFF/r+vSnaQrcHLt1JeXYG
gm19/us2xpdf81N9XN/hSVeJ6YMetHJpHV8ObCuLADZ8mDNRxTs0s8AjlwJJLLNw
csecaMTaHV94YruqY0DESyQjzbWrgjvC3XBJ6aT319GYYWH6LBL6PJ/uNMDSZZxu
BKEGp7YxAbTcu+Bs/ww/4NVfV8BklwzdOEaOaLuKFqfzeJ6FfpI37r6pyk9TS8hq
mKnOPO6n9PE5hnCBe5yAKVIQW5HizIpfUUkbVyJd/hqsArdVSJHz3xfQN9oRNfnE
7L7AMpLgOSneP9Zagh4vEJpr0BEMJTJB3W535fVd39H7g7RSrXBqAdW6lv7DLFnx
qqt8/Lypb0nzQf5/1V8DLlMXw+FO4UZvejqQ7R7XITURTmGc9FsgsGKYA1iuXqs9
IAFbh0VYzd2nwVeKc58t1zGfeEjm/I1xH/uQgh/o3rEm0Y7n22XTikB/RRQNYAd/
hVLHHxCkSB+4urQwal+7JflcOuNuWboXcoMrKX+RcwubUJ41kD8hOmOn9uHiJpes
bap3pi6TtcZNh4fcvqPLBRESt+WuMqDGLcNxr60i4RqgpyTpuVJH3a3uiY2Ye0lb
CsGyrMGm9CCE7mpCEhEBxtLnNrgs56MfXx6RDT0C/qP2RK0GuPIhB0jjRYwsCg6o
3qURS1XaobLQ9DjHwixPn26GJIg1YVnSSNwnd04Ed+BnSl34TvJ1f9j1doWBqj2O
Bo7sM5caHKnrWBcwpT7BI5BIFicn+9qsdz5rdbn881ei4WhhGhYKTloicHyMsqh+
NPoQDZOdkfIXDJ9e/Cxz2irnx/fFsmCQ3Plmnqc6fyOEXzs5jSeciHuD2FxpEG23
0cu6qJbTMVlVHvwjMLxVvs5+vyjU1zDmbq2tjH+kqipk5Eysd2ed3RJ1E68JcffQ
8GMW+PKSNjJrpke6Xg2XsakpDb+fcjJVmOfvWMVCJU0YOV6uyySAx7btLl3mXaly
E2GN8amc9srVdw92x/5QH86x6TOrlSmjNjEtGjeN5efc0XQXyH+aGeI8/IubOsin
4Yx5Uw1SGn3Kygf2f9Q9vMudGVnJHgLokaLPRa9CcG14+VSGIHRY+d5V+Crac7E8
pDB+GY7ds/AgT/ZCWph1AhJ/j2i5TTbXYOJF0V2R39hrf2synlkzBV3S/KelgWtU
gTi2nuq/GPWRjozeg6a0ll2/ipW/z5HVegLkRsXWMCyOocp9Bv2TF8976Hp+amVX
1rA3egeuU02bYq7GuyeYS+BV04i8CntTQB4v+vfZqSqCo+ulZs9enUiFf8HCSDCt
GSKpowC9jTJDKtTH6VXpux585JMCUFGrdbYsZ1s8usGYZirkdNvQP0QS1SxVsnuk
hJOHimP8aDmSwGOXwfGc1u5nXLA9gKdiw+m8ftbG0D6AX/YFIN+nZJ8GETuiJkNr
3vJjtlKz25E1X73IkybHPZn5w4/x4FMZJ6KVWs4bSn97bcYEeupl4Y2VhRh3him5
vK5t2MwWAqzV+CRJMhf2umtCShU6yuYQl8P6bPzjwfJ4315QTpBAkuiT6Z5T3oTA
EyVya5OskxMPNTVUna9orvSKhMmfr4F5vDXgjK4ChRZysFK9RVtuW8excXGuzLrE
tfTc3HBEi++aCTVH1N0bWcFTKVLVC/BOQw3m7y7PeDL++vSfLW7QIxwOMpxigoXN
KMVqKsFuI3rseDhZiOi/PhmMlxTAWUI8U6C4zGtELrXsQXTsoidKN4CqdAK7k0NH
rTZ1Aexi/3rHgiWKdCwZcMXqnTwjqn0fnVJgJw8VRDarMcH9OiNGpunSXdM99Y1R
BZoPIjV7Kr/DMj0o/moU3xpNNHmeycSOX5Qss19FO073+Z8pIAFrACvf1epVAzaE
JxR+WVQdkRvrc+Mb3yvf5nZHZ1/60SwEERHX5feG1yZbGTJB1l8TS4BYX9RdfSup
6cNkRo2LEPPBGCGx5ywB9ycA+wxAHiEcMVbOH3OdKUj1B0lSasny9RWXIgkodK0z
e7SORSH0E+RdbQ8q550tcVeky7cWnbMwa5/J7GxJfVyf9Zxl1pF6fF1FM1Gos4Ug
VzAC7vsZ5u9BARGBqBZCzlv0Yiyil8ac9E3H2fu1UjedQMcIJuBOsCmFqxKaAG+m
05fVqt2/DYzUw5+PC8khU0C90RYWKCqs/8fmWmkp58BeBVWZ4zwjm2aQnwlmA+gL
So9/8A6MtvE/ZFLhTbsLogFfMLZRRwdGrF7SrFCeN6C3V/AbrRlMepZzMHKMt2Pk
GrLC3qyLgId1XpE7LK0aCwBvM6pgwF7XNUAaWNM1M/CtbTraRLHpGXGaXg0FPu5R
f1XJbrR+kvfXpsX0xTae1VZ37tJ9k8kDuhmldNLbiMFEu+6gxPROb6XVlfETs7sv
BPR55tekxiY5v5l8LC+tP7PXQKyozxWh/7CsHrT0NjXLqdo3ekzTTgf3woWTLmg7
UhaLbcFXsXaTXFbn7EXb581MzRc1nkSELlqkkGh7Z18kXGbOQkff/E4CucurqgK8
MhmIGOPMAaZaFRc0iurpnj++RsJ3a4k35my6IetpnqdKToj4WajFPb+ZSlGpcxwh
+UdE9hBx7LuxK2AdDRzrso0GDFxH7WqD5ecC74FfecKx+wzWsKyrD5+CQrtWXosC
m5VMIc4R4S12Wpy5VXimA4CZ28hE8+INhnEb6giIsyXO9PA6HEbr5+YJ1HUW7YVw
TOOO5W4B/LA7h/+AZmaRk2Jv9ar15f599SsX5rqV/gu5toBaJH4RzscCuFWEmU1Q
ehDWWq2HEGrDwXFTwNFiIzT7BbR0DqM9BR1Ll8lUNYi8vM/wd67ENLBFB1oEy1a7
NE7fJ2MoMAdF4YOXKkIlf9dwdITvXKkJ4VaB6sZRd61iM1x5f8N+CZ9JCtJkl57K
MJCSjBxK44Q2O3D7cXo3tGvBiKmNOMm/SazHNsKjr7aoq/mOh7hp7q1WkChODLsf
S5a/MegP3+YSSm8PVHX9Q/Z5O34apGuOlnZzpsDINa1Iim7zbo8FZfKmSlhFDEZL
qVmN4pikJjfb7CHp95BS1ShLkCwYI/6nOqhkno5q8psGQzd5+kcgpQJKyEmLzweH
CGLKTM0N4vQeRcTr1vRR5ycX22dNOcX0vH7B+uH+RzwaiKj479WJXh3n4YnMBsc/
iZFvvoTo+ixv0krPhxZzhetxh2Rd6wMtfzWAvIzMAHLP7fTfZ2/VQPfWhRpXxtL7
DNCVmzn1KdyBSoxomlXcpYwzegfE1mnPF/sNlkNZklc6fBcQaVvVUTLJDEOBTf6z
zYz5hNMOgVNnCofvU1/D4HkpmGw9waB0zNPIRZ9E45LZgTR8ZzklH15b5l+zw2EP
E0YKbghm76bgHmdbWT5AkHwvdZKjfrn8DepAUI8Ioi8Wrtu8zbIVyb+gMhhOsAnC
tKgNSYVFnJ2gTsJRJOB5P6hiNFR5uXlY1qo43PfcBClHVZn21yM1n+iAnEuZ6sor
i5d8n40I3gLCIuvmCDLdZwcAHkp9ePJs3+xAd3cZCHJBJwiMUwRYIfbXHa6XNSp/
r4ZCIJ9T6AEqxdqCsUKApw5Pvs0Hv3oXq0oRBWGzi/tyaSFBagzlNjw/nl5fm8u8
mbNIn9y2NmkDrcSr4l8eQdAPRnBnzsRY1furrTiVkUF/uVS1jLFY+FN/EiKeklPg
MsANloec2hh+RTwZ1DdAJK5Gcbaf4Tpxi2wrruNUWKAvyIvlIIh4dmFvc4Mlk3H3
00EZA+8q90XtSn8Cy4ENq5QVq5gH+UyvXP2XFvqcSQoySwLaGsa+CsM2B2VrZkxB
qZIKDZ3/Qccvr4IvnpUQPZllM59Go3DjknkBSmwzCgMnP7sjJwOYqScCNlDRYSAM
sGRKJcwZTzmloEdMYzlPBuqwI2qgrK8N8gRS3Rl+xlJPPMzBzPbXhsQ6thOYMOms
p1AVqRGxjCa2vk7lQ1CWbfnHEj6d3IFom9Tgw921qHs4fwGTa7uYFoMsnbusMGem
Y6THGaqhnjFrtd5IJOj0uLDBgviP1/KquQusoFcwNAfXNsn08NBO4954BglX56Bm
py3fBrF44dv0sS8Ljtu+qpQHKbXfUtQDqbGrs/X/nQ35FEpuN1bGHTR9Z9P6Rlut
08mmS6kH23FJaHqPdoZGVDv1ffrQyDA1/ITv1wZaqJZdj2HoSzMTsh5PtvOPGROo
f2CPFWoCpsCigKWJeTfOUZeNEsbGmuha4RDK3bXKqOaOikVkYEqJXbPUfQV1+VZf
8NFh7F2LM/JUg1Smmrlz/e4UUjyKKyJiGNjytJ6mmsWpsA3QXEWs69g/l3O3//MI
1ZIe6/0BHK/pdNjWs156ppJDt5ehFMojsX5mJ5dEj2lQjKGLVGEQVoSx7pDoP9B7
rwhKIspVm4C2rSXKovf33m/7g4cPwgDJ48FmkzewnAOymF21xYqirBxiHz+eUR6C
bp4h4ODrkbMb7Yu9oJRTMyenwmVxDGyd5Hch32xDsgtA2WoqPNxWJF2m1ij0qmkn
8jCVfmq7MFqK5GSBPN7wHV/0FDcaPHZZStLG+OuQLks/vmaI7FFRxhJARGylNYJT
D40JedP8ICEKvkxcZ711MUKRz2VsgxjHw+FzwoWOsNePSx992w07kTbb/VzM/def
wusrSM5ov4B8WIRioMYk1Ztep1QICzUWFohr7lQPPy1xOi73O02TtMY6/mgnhV87
rjmOy0DR9k/dMtHj9Lfqr/jk9NWgUc5MaVxqmMb1q7gDg6ofJYFow6Ytq4DQgKeY
mT4yJ/p3corZ17/5DaPUvfOd/W49O8G4zhFOdz4YcqgxGsmJDxh8l2BldfyVrTsG
6aycNDmT3kQL2QTLK+3UaCN91UGDwIngk/fSFpYFOF3zoPnD+DO9bGBODl7u94xW
QgzvvqldXQCkEXN3FcVa/J7sQ+aIfxO9Zco4+tM4HJXj/UHolliEXf4sHbmTx05Y
hXDsRgbUYtWDlbh3j98XAkY2SZsosVXgg+MP13VwnCYXfO+pIRgDG04XEeLFPLHn
XEPKC2bZfLYFNY0ciRT0FgeW4KUq4OU3WHemyHtHmi0YnSm/ph5hKiwEfvYf+2KE
z9s90ZOrARoxhTqljae8sLIMUjN+xHMIMm+JfP+gxqxiYmmiqFya/wPNo2s0os4S
dZpmhn2E/8nUREecRaGt6vuvxbPNVqvbg8mo9m0fgDwaCjr8F0SAprEKEvRF0gki
RLfYWCWHi9l+0ZdaG3GH3rHTQDUqDJrxlnHSbut0oHCU/K76ARQTxbua2AqEiMXC
oeedufbXOQ+wX+vbhJLlt1qkMTseujOylKDTWpgpmkc3FnkKJm1O5eI6fBe7hKKm
jnvpqIl2QWDc/AeJtHruIb/tki5iQc6LpWYB2A06UfP7VVn+IcIfFmm7JWjBKApq
p2xaW0qfijRVew1A7cEQ8hYGbj5ajSBMbEI03AWG6GMUTNMnpgk30Gy4JYDVEfJy
9NzDZzHsMan0K0AkMIyE2CxOaAJ/vjfkQFKPyk4+oFmWc8m8E6x1HVeNqxGmfcUl
enKkCxxWXWKRBrrLApbj83to8sLLvcd26Th9XyrI5NquQ77gz+nuck5eR7/HUPOv
uz8yvtaGOLrU0lDam6lQHqAmKLYtqiOHs5xq0pRXlzL1Rsk57EWxHuztT+mpP0vU
FDOwpkm8lyuV53TFMnslQB/l/ysauzBgjr7aAXNK6uhBTzsjsKFSaaKBHKZK8+T0
hngOIXi89XFiiaZZZcbZRrSc/unAPP5gG084M3mWZTRY/V4YbZAUVzTjcX86riMi
2v2A+djJ4PPh5qmR9dVj3CzywQA2dAihzFVX/kcgFjvu8/Ijo+2VSibCCvsKpbw4
sHrZ059WesmIekS34OZXO14PziYSKo0MM5zXdsI8U+XusM5EaotgZvixOl+JZqr3
WyGwMXU+keSnEqeAL5wkPDhQtWsN5s7h1TzliFSTMJtKFCsJqyG7CU+SLZeMNrLj
xnj6vwh6cBiRubTsEazwPiTVG8Vtu5XSLqkVqpxz5rDB8y5TcrbqZyjgwYEyCeGk
BMnXIK4qr1ogguiA6VUlPjQaKSEfPcH8Fxul0G05G9LZhuOT0nbvySxMB7jK9Qv6
jgFOBYtyAexu/jFBgotPsWdSkhwQKtLz9R8q9oZ11D0aqxC3Bvm5qFiusYDYsd+e
3RJmmFArUfFz5bHhRfEYkT8x+KaEPU2QhOOTnDDR05ZKns8oGjFoz2DBNQoILGhb
c/5rGXCMT9bIKb3YL9FcWAK8QxsIfnQkgq2nlfciLcsBWVjxQSzSQyFeCru1ZI+j
E7e2rorReBpRAEh1+W6La9GfrTQNCfggluSMPAf5SMwcWq/X6TsRQCwsXL7sb0TF
AkRlG5biFQE2+LZp9F1+kYx85trx7RmBvnrG7t/2doWPM5uGd2zRYjQDJn+VNcSF
Ttjwmh2D9HxhluY6LgGdzkWqsZkslx4kR4kEUVhRkMrp8a8mY5sW7WzPMcyR4WQn
NhSTHg2kILsv1Iq1v9MAAPXzb5qQU/3gJ5IY8VaiAqairUBudGTY2QSbz+6h4OvU
hVurYfuU0fwGTG5KMQNyY/tkZv/BNnah/uo2nxgmxQ5R3jAt347VnamyAGaoFhKk
isUtCJHW0bCka1oshhc/VBi1ap4uY2BMXDYDKd+KzkDJNgrxmc73OdzT5tV084bK
j8yCSygMeA8QpMqUI8w0Eb6EArNgfolXn+5ZHfOfPfDlkW+AQg+pZYLM5/UbJbdF
iGUaMX4JKUsku4TB3z/jgDpMQ3r4nC0emQZGgsShUiVkKYbQ/KZtmZWigoPyc3fQ
CzwUYb8Kpw2trkoFTIGmmgqaDI1guHyXzVpgsZRIoc1yysDUyqUVFxZBsDmE5N0g
VTlfZR/7Lrl2adiNTK6v0Kx/By/NELqupqYL0mxYemznqcUIrQpi1rJHqJSYu3Tq
rXlIV7/BVgQfotvICxg0ixa+40IXmyDjPEK0wDeFr9x6Q0SPqJx4XE9lNxoPjWQA
pPCbf+Lh1MEwhSmFU4Q0x4al4sON4g3qjd+S97UNhkH+fgXvlU5YuiJ84QiiBpFO
xxmdlBQzPNadbux0LTbgFHruYmjKTWyQ4HyCBgjbWzK3MPoBECAkIFATuB72PFCM
GBr3qz7KLh7r2Z40bHoV6teYMiuzBKH9/YdqDOuFno6OCS3LqLBxceMAtryBR0WE
Bh8mflLJroMW4zlcNLrqphfYTP90a/l7Y1INOJCu83Y3O167A44eIl7Je7MrySrj
8TkpMVf/Jea6G1iebcVsKhnGxDtbF9AgkopwNNMQRETHOcalNgzp8XvsvYbZ4ntz
XJaHdN1PQSCHDOv7K31tn3miPFAt1MbgyLhdNg7lwTyAc1Vc+kGwAXva4MONtbjO
6rgpG9/ME0RHq2mvvYUicAWygL0xw304/cFYn5IzFdBZnsJR0WA5WGyMLV6Y5Ym/
JtyWdThW5IA3O9pcu2rEgw71XTXfn+P6iwGVNp0WhufTsN9Afxh3bV09FvDTghcF
pKWtZ4hFNtVZBiRdTsjXhuxooXkgwF6pvQUoGeERGvPrG/UCo97SoMO3s/7iTtU8
uBS01HjfheY/RJRRFn6OjfTzfVI9faKnH/N5yy+2ckWIt/qVKHm44ou0++6XdM1o
ebdj0RGgzewclaph3md6RjzM4A8kiINF/Eui1inBRIyqRE+451JDh6AZDDUfbSwq
5RBhRZQ6VXZPShElQCp8jziPv+fxkKp9eAp+nvWMbMrvbYNipbYbrcKCwcU1DOvF
UcQx2P27ftnGCKf8Wo7lJmeIaRbqSjVkOnUAbJ/hheHsadYyhKUoTlF6qdk9ESs9
eX4ncEz5DFuB9XkkzCJKjseQ3xfwlTwX3lsF3zDR/3Qh1YqRKRmCJVEXzmllbM7S
aeCcw/3Ys4YNlh7atYXQ5YEWVAbu9JU84kdR36yF9aevFpzZM6NG57F817pX4ym5
mtaw2wccOqmCWtiipdNP46E4HG5rRR0e+HsKd0DLWPYGRmkyLWkV3tuWsDRVQvmd
uS8lF5FJrUdE8BWLymW/L8aaVgyJ/VS8Pq8v2wDIaD6nf5fXQIUJ7k5AYw5QYQGZ
LT+sJAAA5G3fijuDkbxWiPJNb++yD3QGBHhEJk60dc1upqgTspIVCLFkT34T7ROY
9O1ba73ohL4C6dFQV4ewH+ygkY9msSTTWh/lxm2wN6nnYOFB8FsSGFQAVVaFtx5u
P5WUJEDFCm+/nVwNZH//1T8jvrPMIf3sn8zmPRFbwUv/tgd6zNBxEqla3xnfX2NG
DZlbRTYBVfWmHBBKh6TwZ3J0uj4B+Lp24uDin6IdBNw4ygZ5LQLl40/nPYUH4AeJ
w0vdjOpMAU5H5pxksGkeJWWsgMSbQLGGkpfTTLmL3ag7bXQPFm6uQlGLKBh47ede
1AxSCVDBl9bWu4O1iui9MjKrY+dr+AZySihh85oFW1TM03qDkxVUXzlsNFiH54P4
4T0kQTF6oV2LUQQqpFN4FTKIM/2rmkOxVwmJnieGDTlumv4D6iSJKh4bAwpyAeN7
ykcF6Okik9g/xK77uT7niZUfx29RSVIZgi4cxvePV9YDTJBZGCh+m8RH+dvSLgkt
HsRy1l8ZsXAvQvVxKs8ym4k8G1NN0ysQO8ka7GgmZ6qqmiEfUzsr1qQc86DuJ0/k
sD2J0oE1wFdtZvsQz2Jon3Aq+VXFMkLhUYtQkfXtg3U043hS1xquj+dnEza3CsOB
EP1J/q6S3OPvFP+vi+FTtG6F3ZI+ofriVE3dWjiiqs2fVEsNzBQLnz+DJFaRTRrW
6u4jkVjVS72miTF6PILouvBalVQ/upV7TjY9VIIvKiUYILEOcOCx/L1pS7b0iVgj
n07vkBbZTXm890VQOp/RGG3yKa0dOjsKmUQRWwhH6DDEztX3DioV4pUPvk+zNqqO
2QkpWmGY3a+yx+3tC9uMZXxWIIKspIMfePxULIA6OhAyVCLQVbDj7x6ORHusCvY1
h4X0jGATs0WsMb0n72og2UTItb7tz86fDfN/HZ3wj1Y99/3OHwD1fTwLBkaDWTM1
gtWtZJSAFuWCU0aa4lFEBXkHl2uizn3R63tu+M5xIdKGEGS1w5yYNKz4nyGgAoi7
h8zZuCUkBKRCnkbFlEB4EtU42oadrejbUbm2soOTWHIEebrFuhWBKdhlPI7tZFNp
zSlC9MC4DaZN/1i8q+1bVfL6MKKtujzE0gUKtvkh9850BWpHpIp91qsMXxmkMeIa
gavJ0DY5ze21oVO/YYU4rsbkILYuMl3lX9oyncnds5W+zmmWg+7lAGhgCnZG/H6g
zungo82UgNlR0vFTwQXmlNMOFCVob52YRusjigTgufZ60dcKUBxZkSUAd8vNdhar
DZeLcLO1b9aheBxaOEUeGaM2JxWVUMXTiQHep3+JK7bi1BSFV+j/r7s/xPFcGI0m
fPE3pk3Kv+yRMRcdWQ3sWuuaH2dIg2fqBzc3gOPoK823yf+2Kut/JvTCLclGAfYX
YIQx+wcndsQS2uFPQE1OGnRQClata+0PJUW448ZwidQm8lfSbYY3uDPT84tHwRNE
qOpfXZN2vxCgBVN/tETCVFaQAbvk5IngEGtUSXOffmj1TA9SHRHvkv+jDqcjSHQR
FVdtIBTmTqN1F6rNey1CbNfkvYZ8Hyr4lj8PrZgQq0uJW1GEg3tLcvFPOq9fgxom
8U+abk6P5/YEVWwjLtIkeTDt5IXpho1iHcZjvbE7NFD7BLzA30Jc1pDVLYhD4438
XxLm9bttVlPXzVMk8rpTtkMAuAFlKTxWEzlCBLblbYiA2kXfyqqnqStknZESEvnq
eHD1OEZYPT3+hnPVuR9QbYeb0S6oJyztbMUenG9Z9iLmq1Xx7k8msi9tK7q709+c
fKcgTjq0OL/h4NDZkGl/Wcx/AeMR/QJWwyR6xrC+ZN2NyR6i2cQpaeD0zqa6f29/
/TlddMFKWWTGMAMnAfK3eYVzk5zkEPQ2NP6GmDS3lQcA0cxdicKpoNZNbEGrPKDE
2EsNfekR2JzgymwoI8nK2T4R+tMDMNyDHwbHeXTJyIlv2aBXnk66Pn5rO1ajCIYd
krPzYMAKOZFivlwPYLUV6obeUF1Z0hxM+NCunNDpTWnZDf9LjkGxQnCg3fCL0Pbg
buhhJE22YXYklqjSwPHNtwOlKHhT5xKIFxs8Ep6J06DqzgwF2hojcIQgNBye0izI
MS/mjJQQiI0ulFpiBknxIsKpXFSHExGtCbgjIAZ5OiSvE6J7xSIyUJPxI+xLNaof
1YkqlQOpeCWZUlinVrE8ivAQDHR5p8AfG1fqB/1YEbWDfKr8eKoc/SumAlB8mL7g
ocSZFyr2DMRBnw8EpuTNnf17/TqbfZcACNjKTKKgzSLvjqvaS/CMPOqQzeSfMAYe
NiGkgcJvXnz8mNkTZP7Jil4rPiT9xmq6rzk/iQHpwAGcj+cLmfkiHZzZA+XHp97b
LYMqZ3RDHcDJ1bTpI5JAAJLMyDK7A6jZ8qeuguvAIBSJs9MBaFP/Mm/MjprrnfGe
3eI/EQWaMilcNy6JtDGeIfaksUsitRMOfR2tv7NWEbWAX1Sk1VU1TAaTDklz/uDb
i25ZSoDBD5H5UummUNeXfOUBv2MpDwRrNFPWNulfB0c3G/ME0yMjX2Txq2LlWE1s
BO7Yqx0tWQjVngooqUCsqefbr9POoDQQWURta9w+qup1Z+nQV0+fRtuv+cYPVTzr
TrA8PPF7f/EFNpAdaMBWK8ypEpZ/KbTxft0D8Fpq7iRZ6Id/PsNMvTje2DdvUGPF
WhGQxvNamWKRcZhFHstGQbrpKJ4TjnsS4SmWHFwZUWwztSlqkjtE4d4V3jtCTbIS
CQrpatZr7scec1sN/CYGgdy6ff3gI++Qv2fBzRNY733RWZNJi//kh9SflxIlUYap
9BP7JL7O0PZUyzzhJA7WvaW0ACCPPXem1jbmaDaa6yqnDFd5lITekgRluBldrPhI
afWlGfrMP/amSIlyJi5e9yo07+PNNdAaaQMIQIXg1rn8/b3w2JzphL+IaUlIhBQk
cGUzFsLdH1lV2UyQQDu0X0bAncMEag/6GPvtWgSv6rl98nKS6ypdaOx40sONaRJ7
5LSH+oGWg5eTBLAFnftgHdLbpas3q2VU/cUvATxAm7jh25zkW5//ejpNVVmcTz19
1fQBsG4TzGAtPQcQLC+FEHz3+N1zopzg38JuvAWDIfJXLF6pTTABw52yNN0mJdoU
Mjftr0BxbpbeY9tIrM3HnKRjVyK1s3/Wlwd3wHJpjq2x/UesaUVgMn+idpdd6Oor
S4DTDiUx7e8GzCxpE/2/QHwHTTHYVThnugfqzn5Wg/RqlXhtz/itgJGKHGI3/ECR
eAvoHXmqNgPUjsuL5pBno9tkBXjxuCXYQwG8lSZrTjGNClR/rmlMqfnnJC8I+bSS
UqdNxHCCOarIJjPXEqeICa6VUTUWSRfjlT8yNiWpggoX9WYFBDRHIrNv1qd+HyYE
7xTF0oCgEfFQU821ivrePcUL160fepFyxm/6SN3rSCp/QTgnXiWqBFXoPRx0vcdj
njZcICVYfs8ERNEMZb8fitXhDmu11iAB50J3gV1q0oWY7EOt1402e4gSbZVFEbU5
SlYpBAm0hW12Sgj0ERQlZsCjeIMuZxkkM26uESjfIRkAyaAqVs4SAxYuQJVWqf9G
DkJeyYVBnqV91QoZkTKVMgQWsKiCrz5A+UXdtLUWi+eEOVb83EJa5JA8OfF8xsML
+T2I55QR8P0L1qeL3fBNRNxVSdMEuPk9LKZfw6cDbIFIIBrEjEZzHH7Zka2RezT0
+WNGPPcmMosvsDIU9G0JHmZfhNlnEfK4LY/Fllm3JTumUXA3YWXMd+dC7ZtiogBu
bKB9E2Gf2OSaVGKSKvT45cJkP0pMLy8wQ6EDe9tyyb9haXHQcgKWuLB32VG0da91
3BiHRai1iYyoXQ77ijA0bNlpJDL8Zgthxxg10C5vj+72b7h0JBCcesce2tV6h7WW
qJrtYz+GAqeNke7960088tbPnSAE5hpFYqM5c9kOGiWcLu5vodR+bNmgkUMBON+3
ICLPl5eiEXGwj1nmehGupW6ZM9bKE+ItHWDApUH9DFPyZ1goh/XClbGePNsPVfj5
aFGKKO3JwgXRcf4wfeA2zEfmmNo+wxdO4W4Jx97cEd6Qm5JOtOuL9CGiATHUldTf
4O81c1yxnCv4Q9VUTRtyVT2gLfRZ8m4QP+/OsXQVmL5Gf0xRuDffu2RzFqG9Tb+8
c2gccYeHf3SO/0JNYpgwibipPhWLLRySo55P6wnp6kAWSjf9tU0pqh4nyrxvFEHG
s0NxborhLD9z9w4OXR0oLhS5AALnCllEDN55tL3xjfNgQ+rfVYoIjYd+WIF/flQL
vA+g7e0dqTDtU2EAI9q5wguwVEF9c93VEKVBot4h+hN2YHlJhSpu2TzHUDvM6C/k
WRkIJxD15NvnyQf4Q9YCypljnAFTADhEFxo8T13l8qZYBFKp9K557meW9QkTTL16
8yh+BFNTjP43NA6cJ8PnTcsZzDZgeVE3IyK0WuyKMKOlBote48nQUEdgLzx4dPpO
1dM69ammldC8gB4IB20WVsw3xKxCua6+YUTmxL+WvVEmYy9ZEXRojFxtCYf9QCyB
9s0LjUsIiFHMfwNqHnonT24I6sh//cTFO04+WcCR6ZpcqZRYFUYnzB6bwVwGZRWq
KETnosxmkfqmIjjPlwQNJUFFoYY5qpekLXsmh4BBWpftcJmteIP9R1yd2nRPLbJx
EB2lMxq27vkUwgg2DYA8ksibBCEK6ONblJxDpUaMV7HTa8PJT9BopqcV92zE1tQG
Klo+JylW+aS/jBBf0d8lKZwMUIpZt2y3RFoPVLu/PwMAUu6npqYx2tOOGngHKCvo
C0QqdlxLGohw116n3BGGojhzgGvVPLtBtCDxwiXMLzTLIY+4PqvCmbLygwPcOUvJ
xSX+HPDobbnkTAnHvEpcpXIpMcR6kRkJQijk8XoIZlcVFwjg9vG4+U+AzXR87yGN
h0JsF6GuU8iZF4xBQ25EX1nzYJGI9xEBVu8+OkTUBaU54Qv3p0imG6eUZBsAPDKU
woLUTgmAW+z8dERKsru+ajL/3vWE63yWaTu5tLTpoR/JamvTz7yipV4KNfwDR9mo
ENR7RvrCONTo5RSiCwf8KaXlM/q3ml90Xb3VtV6jOMaekPdWnhDvFnL7SeYV9E2v
fwJBroCOcS2/L3FKxG6XZUqBWvg6lnP7hUmTphDKRcmgGwW+Tuk5elNsaZvmr96m
HI07QTD4bGgYQe5G6IeK433haLWJljM+aDojilY4qGzThAfvJEf+MV4Ka2YSQU3G
zEawCuXadG2SU2lCrkUYnFICjq8n6JwAoY9A86R6v/9kjPN8c7CGb9wVvUYnvRkx
xEMO72pMF6OTTkSAfjIlqCzne1kKQ/cwL2iUoB+fCIFWK+L2RP31micGAQyva+yq
bAjkNqd4aZQmzrEUIbRzqlRynL/hox6C9rhAA5h1FuPjS2o89Hf95TSo26xlpOZs
0BvnMIDNee9l7mjc0U2R339oB75hqBqFJ4enyRtb7iXHxaaG3+BcTlcmXbbDMLZl
WYKoQ8Zpr5ca7wTKvRlgxF1fG3JVYcZvtoFlJE5oBGOpn2IvKpI100EvGQX5nGUD
nElapkE4wrjDtxvTBtU2OR/I7pfEXVvCLZH76XSSnlvftJbACcAbsh2Skc+nCo3e
cBkwnoO8j8BHx1jitrsx8rAYRZUFbSUqiAyfftoBwHCPGAqXTKsJwbcMJO+21Aky
c6JQtora/GtAH71JKC2hXipwe6CXsne47VY7DBaKxt9xoCxS5sc5dTHl2ODyPskg
sxJwwP0v/Ei0d5SEn7KhGzGGDs+GAerdI2vPKP7NOrnR4IdcSYViUak9+oU0AdOL
5vuleBteVpxOPsIH9t5Yscavt2DU50t+TW0yDpXkcqMadQAz/tKHIusbO90IEfw+
qO2t/v8MdriGI5NsdfbC8iNwatn9QSQoqaBM9F1Ehwcg29ErKEtiVtKBda8oC5CD
weKo3JUUFaVZUGzTY1kXC2m2zo14Rewt9znpMHR8O+s86PfpTMWZetJO3tnYD6Qk
oWpuISLpWu/Ifn5z0aEWOMK4BK0S44eif/f6Uu1pTEsnasSgMkFN+hXZFpXDSE5P
Vaoea0JxqH20cO0XYRBCZOCZRTdZ57KnNUFW2eyW6S5R12XpFYlMtkQ06UjZAYVm
YbQ2BskW2o9ix0/OK52XfcAyiYQBtXQpV/vmGd9c42Jm0+jBnKSO63AUM8N9gv2X
4ok8LgL5vAKB2J5Ux/K8GbBivK6OmlYKhwawl5eqeSo87V0PYbIwLZpX6KrhCRbc
hYTfcTzg/fQO6Y1xiWrUICC89Dv0XcjNL+w31tpQbE8wslwmfo8L+aIEmm9uTVdS
wsCTNqFrIbT2h0oeSlpr4/pweeGkL32xNx9zDBZmfTj5rgcDcOgdlZrS/70RVDsW
GjfS8ymNKpFFJXng2MG00KcgoU+zFOdu+Gph4OjVNKuVeS+9HbsWf5GvV1oVuiOS
w5rk3/c8wvTSfSEBwQUSZ7trgxNaoHXro8jcaTffouM22bIhuXy//YvqaQSs6hjj
aLRNxDtGqpCX+M8eUZ2C54N+N6V4lNS6AvsyNZ05c0HDQLY+19/TZ+XFJeHKkX91
SdPwHqdKebcKO3R65scJLrDzjHSX+WMFmL3Ut4QeYS4=
`pragma protect end_protected
