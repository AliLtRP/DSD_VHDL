// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:02 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lk8FmDG94inTi7V1cp84xPG/+TjUHr5fOVEEKIFy6y73P7H4hutOy+TBI0/DFIW9
HfqGjRylz/blmEgHdXG3Vf/InBeBAf+fOdgOODLQg/N8wxzwtEEfwgqZ6YlI027q
gvIsSGOusJ7+dgZgabBUX+S1Sli7qHK3kj1OGETRYUk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 58432)
LcIkvHrXORM6ZAUecIVubcZMkBueSFbcud58dvQOgAniAqXUTq6Cr4jAs457zgMm
bii6vdNnLd0ZnRahUyAnRUGSMIPUCdt7ULnkyrPBj42XxRquf+gIH9I/MnKASt2U
B9zQp6SBIPPa8waE9E42+ZdSy7RLuQCB8NPIcNQBfRlX2R6mmUsNPVfyhgTXoktM
k2E+XuUHzc8TBnL5u2deqdjZj/Vpj/rgk4iPZ119ETElHnHBfRvtX46BqBu1jVVK
s3aJbypLAra1eEAUs7uhH4798wvb2e+FONHTTkKXtdps1EGCkx21PJ1uWmv0Lj7w
hAjvXexydILYpNeMNtJjt5YHiqEiMm+6qnEeQBD6rU6aQsJkw7+l3u1WHPJ8Ue0O
STTv0OmKLyRscJLC3cqVTVjCDM+QQ0eCb+7DjG4GVJnUZ7+neopJMX7IEWP5oeMi
7paQCvmQ0+GZc87Y3XWh3KVmEQopDILIBWqd+jxt38Z6w5DNXqICrmjMuLC3Z5xB
kU1rZMQ83F38MYzNgiMtVR5zNFT5XhNfCaCfThMLAiy16Qi1/jenIpAFzQUuOiBz
Ga2SVRHIdyWv54gw/XBW9jGWG7BWhkns729Ge1R7fyYLHzYKTjpDKqykUHVGLnDJ
Z8A/Vnem6EnkPb4+JVMjvks7aqB8SX6A6H69botZR6s5vgAAqnMpcJZ+UH3r1qgg
ZsmCPvnpvH1Uz4Pv+4S3pi3jpWI7F0jTcZSzUeotXoxzOj9URseOXZRWgE2bDYIK
pNoxscCpwxaXf6RslyGpPHE7ICFGgZMKjL7pmJSsoOMsQTOaA7BSP7ulxATmiA0j
9LhRM1zxSUMjP6J0nMyAAJuhe7IJsqxF7XdNkwo84+VCpTXC5nlRRhouDtGhtQfo
Sc0YNEyaRHKpP3DvxL/pOSlsZ9rsxddrKrqb8AuB+7L2u2SBIxZ/BIRNlmwALJeO
6LC0yEBjm4t4zdB8DAWNYs5sOay4Dgeu/0KTED5vjuUo/KgwyagI4QPBXp8Y4tOx
SdOppFkie943A6fHt1SyQq9XQArVUK42aek/aZK8NFZRI6w+V392ahUAdmlV8jSe
Vrntqh+txAbz41qNWOwySlnRATwUDCtKG4j98Jv2Kim6AtOKD9L50dAQlN34GtsX
HrysbnOzMQLfHlGZVIiM4rEV8sU2AHlB/o2Fkk85rNTswbTQxyIW8B9pOpCj9c8Z
rafLnUR2jtHCUNmaBY4+VTKLs3wQkyOBQoCvTTBpmpTj/jbjnt600Z52kFKM8dj7
0AxZyDy19VGx1WTf6zxpOtzB0ejwkKfy3JBWRfZY4MagBraD7lr35LAM3D4CLMf4
9KMXewyB1ZJveX66f+XoMsXcovxULVN/872RcZEHd0R0pciGefWqK3ASB39E0VjO
v/LyHKnUdqHP16QoS0DDSEnkU2QrvHd54I7k1WTJTteCu8Mclg1IYlmGmYxv1OZz
ybV+SkPQ4JuMBsjFTJ+xHjtmR0CwJQ3lp1SN2ToXNy1P5S4q/yZ1sUku5LJXRvK2
kxnn+0dY4tCNGumzMpCnI6P3ZlMGp7NjUW2O41V4U0rapL34oWYUH/0btFYJ3Xmh
dclCVwzxgqSjIOybuEnfm9nTNwZ7Zk/PFNjLyP/+2OEPhEtVafmG41MOxNOTXOo/
jfPdgNMjdx6aOB+UqNxlIdgMfpphvLxuBeG7auoP7gY2RZ72ANuUqRiK54EkkvN/
wTmy2zhCIM2Js05MgLWIdFxoiZEibG7ZvY1yOJOQrgk4d0/HlKMpCOL39vW8A3fG
0yIocB+FtzjbPvUWv9PMFs931Mo+gO5r89pEoIrwGt+8ytPO39n2t05F3YvHMvf0
MM+PTGDLMbyioN+ey8lP7/11AcEQ/5pYTdgPKgbXnrMWLS1dvmWl6Hdkzz0tPNUM
bzWkLCVIAkE7Ck2cMDornw3AXRebxgwGG/jDqbzLAyJef4tL//x4ZSSJD2+StoeR
YDsCFrLQwBYFWA+wQzNghXzpzU2RU5hLHuOM1JrZCUvDILT/I52dV7GJ+dW38lS4
YzV+gdEdyQgB66bfbVO1CbPDmmIwFZsjbZgZkW2Soot6piK4tHLCzxoJCT9xXLrc
1kE2mv70XFWFrKxfgm4YrtcBR5N+VsZkY0a4OhRpCC4eDCIaL+9hLI9M48hq4MLj
CZ8TbGmCdRjCf3hB6iDuREwwHdmq38CV7S8iSFrP/zo7brvUxULYi/IsZOVJdMrj
9gPe9JwBkuLKwLa4+sARowzfDt7uLx2WneJDJeHPPL/PHnNu/QntaPIbGHorcVkI
TS/Ze9yc1zy/fcvfOJIJLuwGc/B4i4V1TFn0mNYXUr94YSDLNzTDdMJmVlDFGNey
VKwRb4IIWRN7a016TyW5LS15Cn1t5rWWoDdTqoYudfxy2K3r5m6IA4SaMo0FpN7N
IwSuAzoCdx0y/HVVOsQ3/lG4MKhZQMp7EkDbs/5DjRdYu7/UFNhZNsAPkwmjrMsa
fb/CBtl3m9o9plQzPehFDzWf/DnED0x2jivEx7YQF7V+BdbIqn6vutd7Q7VO19MZ
GFwjqeROYeqw0MoGvcKShVlUYjyiqSmaThO7jgpQWHHuhsV/cVohyX/lE+KQU9Dq
MxSjZW8DaDFnGDj3GmuYi9SripB+kzk81tsqMtbT2mfswhpJP+4F4Ib+l+rNRNcd
lDXl0LvKbuuk0RHj2vpYXfiWL3Av6WeRHO+uJHjc2Wr3PMxyu4M02Iw49/LLUf+v
ZpQQeJCpuo0ZXAZirW1WKbr7mixiDYSSaCv7hK5BD/5M9oSiOPLtICtYgNgv/Ztn
HbqPyRPjnBixIFSW5SAGiF7xs4/JAet3qAJ02w/SUKpYy/kW/W9u8pgwtY3mxIcr
u7XGxpue2EJWdg4+HT4jkDyXif7SRLnnd3iLuOKv5ZV0Nj0qHhExLS+PMPyPopHW
F96Nf+ktnjnCgaZXnSIUxRpH9nkdRrfLerMMZdbjnuvlAoFJfuE9oORGcXU6QW6c
1G5hpR58eScFMpACx5VO/Eh25Ks8N9S6TlWFKWAeulpUyoz+vvNwlgGZH/455sf/
DIFnMAwq5wxUkW3Jlv1SYRLyOGPSrdZ+50ITm2F9NNeuPWgANdhDgf/N3Nv+aMf6
panXS5/MT6LfaLHTNwH1ZEYrxxBJa7YiPSfIAU164p26DbAh7cP1qZANNrPb57K5
A0U9ocuf0K3hjhppqjHiUzmpWzSLgSePz97QgybVr7Rbu3PEIngZ20dCw+aJ4iiY
mkKd9IZtM9WJ49s9TmOxucsHlelRZnt2NFxpTCAJtkc2Il3jQtXkLPxatz/ytrAv
OCS2J4iWihiQEud7BUI9gixgQw0Hnct3VBY8/CmHWv67VKwr5/QY5uS+gyI4bgzJ
Wy+R99OVTnDHJ9Hm1HThRCeUXR7q84hN3gtcCm0ERderzRVbINR61I4esAkpbFOo
b4UttUBBcuC520podWo1E1SzfdzMo6lX8LBshh6KCBr59Ud1esBgaUkfOCLmEcpt
LGbpRH06N9uWDpXRlrJWUINbukxzUaKNe5IeND1uWzoQ6G3u4kmvj2b5Qss5aqGK
51FSfgJKDTSCOiBbFEEwJq6/EWeeg2ePPIBUc3ynLgVprEAMNB78IGZMWUCRiMrG
NqUYhQsk3WP8Ewf8VqYgVk5+jilKWnimhGZrACjWCKBllxTN1Q1UBGOD8aFkjf6C
+e+xTQa4jKQMYhmQOmpOiGjDHaW5b2naSDL/sTcu3Ru1pEej6Q12r/mscgarbzja
s/xwfdBTCidZIScoarmLxo1BWXHxYLs69Ny/vlgLrQ/BXw3YzxfOkb9S0cOazRuy
+xImFvaT3vcbrUh8mhRScpOfaH8+0q5qYLX2Z62M5LDky+hymom9QSfG/LZqExBp
zuDzqDUowcDjlgvEi2WPdbbXNJ7U3L1zqp6Fiuhf8fewmtNDw4DlXjZNG8EI/Xzd
cF7QUQG7HTpdvoGe2YUNGdpYTcLcfKC7i7PZmYg2KaRPidfL3ZCquKdRYtHPyQLq
rdwEVwh9f3ZoCEqJ8jFY5UyboP3TfMPCRX+fPuQfU8b4C4c+r/1pmTv74gZEdgFB
YulBRyNevPDyMUsLOR8VEVnfMOA40j9ab+OKlPLEbpX2vKStZJwdQslA+NUhRWpm
0uuZR93mY4P+m/pCxDgh70hHmBwZFeLr5jTVqCOTDyvzldysuvj+RtQ3vAXTjJ6L
FzPSMTeye9lWRZytQq5dHcdrMd7O0HRAf6NbIspEOffgZ9+2Rchhl5SGNfiiaPje
aWejmzFY60ukY6YsNQoElbGFGtlncFkdECghK7eqBGvh4a6xgb8kOV8JXo38BI98
bbVeykwTVxjD2kvd3Mu2P4Jn+IwwmjklQyHoMGPaz/O1WMO+HlJsWZS5Rx0Qu0Jd
hU06i/6LwRpCTM8WLRX0JzCVyDCCq1KYhXm7S7f17zvcKmuVr0ENyodbFADCEXwQ
ezvSi3TUmPyOovyjAFXL8jp+mojJENzprQK6fQmp0YmrbqmJZREyBtIJ+pr4u3+H
D0Xo2h7EqmFxH1qDeNT584Xou936Pe3uq44atLlezB9UWa87wnKWUPcNtECcUw4S
6biFiW6m+kzOCwloRN4mRkV08uGmJzQUFJ799LdSIiM3EpFrca9utUXU3dCRuCM1
ymfOCSt/HFKnmaIYa0R5I5mTrQaoMMuyUqDTfA3ekj8sg4Tp3Mzqbz7BYMcpUBWA
fRSvUdOWmj3kmna6RkZ9oVGL3ZH6PFJoGeVCYiBYhT4HxHhCaCNjkIxTUdps8ULK
PsD4d5esMWh+K6eyV89eMrfi11xb/xgvBHJIUxaQZQ2eeWNL2cBAo14QuPwYal5I
Ufn7hadwpbJqi5280uUiNXcFt4yq2ADPN3YUsIXvBi0e6HVyBnHCFciOkY8ZWnU+
51vr3tlVyMMzTOALdOWcsaauLYaOd7H3Un6Z/mOkxcqFOs+phjhUfeGEsVpUUW6F
DvwUaZAjNql4ivZaupKTiC4L74JwS73T3whzHxUs/5Ck3r/+C/oWqE+03LxFr245
yfRWEB1SOaIjixPdMqwHQgUtcfw2B8eQSIklaeDsiB0rqCtzIQnS5A/Wc7MVVIHY
Pe7qYtYghKD3ueytWEKe/hlvhBn12u82F3++lrVfbiRg6g6mvNNXKnbEa4OAuz23
N9vK5xCjttk/V/Cylg372t4/lOt0QMtOs+oro3OEN4dhFk39hSQieRFwjqtSLLtd
F7OxDPmI5Lr87wbuS92174zB/7Xc8S8ry0pO6rHg4blGdk5vItegUhzU7ye9aeGd
gWgkRw+vvcYgzcc6W9vPabK8xZAAE+80RpCKEzDUg/jC/c/Lnkst9xtYJZdXtRtw
+QJEtOb7LMBEPUNaLpyQogKYnXjkw6IFV9dnh3kkI90YHZIBef8M0FcIyOlVjS8o
BxCDVm1vM4H0pP5gdTOYFMndsQ2h9Q6FEg5KisG0NnSkgybQqc/MR9P5Rr/TqBRc
F74iXBbjbTt1MEIigqcaz2nDc2iDZsBcH8YyV3T8wcUxJlh+NhJaXjdmFQqtWo10
TknLcme8cOSZ7eLHyhADbBeCWv3lTwMHTMP+1uexQkpuc9KBY7te/xsxYxoLRF5J
IOJG8iCp/nDLcf3nfPH4rB81orFf9dcAZ5+kGxzofRl3R0p3Ay6toK/nI9jvaMqO
B6mHyVO1bc3HFQsb7O2b/5MM0qfw5YB0ihkGRzPSxL6VHVy3PuX6jnKUnz0E5C32
XpzqdQSlVHAjwNzQAfl+/D/Yt1F80UY1JkW+2/gsHM7SaxUqO5NC7Ym7bbmHLVn4
XyAkt3S66YWS3lSALS1D6x/AAfMXrvdsBVlyrXLQDtqUPzKC3v/ZUNyM1k+mguJL
zqKaUJe7hl49zMptiebmht63kG1KuQMtuiFOwcXcnOYd5Ch8rqzDyW9gYqkzLmnX
UzjY9IoEeCf1Z331Zbbbh3NlUZBmNS2TlPijexjpCuWRBgp5XytP01aD8iHgGeja
hSjFAGrpLX1NfTVpPj6EEp5eMXumQvtWeQHjopD/uraessOnb9yZyPi9jG3KBhWR
GQ8s/PpDaT6qkv1LLN9ByXeFPfytFFtrAlChESqhr4Lm/Bd4RxTp05Ds2SQjGkk3
Kr/V3cj8ys+h0Ykmu5+4wr4TI3hi698ZUJlrGRLbCY9siQ6YTS0c2207kG5gAFWT
FqWBnO0IX8RgE5RO1ctQlmAj78iSr/EZkvMNDewRONtYy/i6fZukSAsGPY/LUsWZ
L9lrwlSph/c2IU5IkBnrwo9l1bNgz1Lk96BWmXN3LLFYD3XUXUESxnCOoG3v6gbI
Oc8pp3C3BWrbqz8Zb4V/9RGSYhimJLj6JgUsQSjjBtgG86eyieRFJLBqFNlpvjWh
LZXAkof+z8DW4Wx24p/4sN/hOrf/tZE2D1FF/emec+v4qNXC1JCuFejZZ8BcVAIP
Cx1n4l9TWncMw30CIfkTYoJH3tstg+nGtSZS+eivVOQ3YAnj5SHRPrcQWZyz5pxB
xtQAXf3T5DhbUzvynzXM9ykQYGquZOZmxiEIcbwgj0v7Ql8A+v0xAE+t6Ic+YKaj
S3BX/AvT48X0kQbXepnFLbFTWR8K1QRidlBKlU9M1TWAsXZOu80R7cLUbFQCyUS7
t94AZfb1CbybUYgjKZwX2lBoJLZUhz1kK4MJ/XEH4+vbB4dItMLUd1e5yZgmnKkB
TExljOWcAUkcz0YXWB//nKxIMqOojfxvG/fe2axOmH1ZIcJAzAgF2jCdqDS4aZmv
muQA3WHEBCgGc15v0eshq7bakzpHb39QykhEA6Y4WWU/dv3EQR5a3YBtS8yOmFe1
6a5767iWd1crSqMbGnfA26tg8+bwNTQMTKNsY+Lf5hfcLjo/6dxyUCoBYgY0LusC
0b8frkGfNyWAVIb7jmhSHJYgSrUl9ERWg1Y+BTFjf5OyALUljAOSHmeWjHTD75ji
BtQuC4K/7q4Plgg6CsdI6TqPrDjVzxX2aX2016TPdxymb5viUyclhDlrVkXmUPbH
dA5PTQZCBPP8QK2l7xx3W0dJGkDe30rurris33lhaVY6C1JVu2XQbB9e8v0fKHUQ
BS+p2I7dcG1jbIZSBj+QY61gzh78O+IiwxwZNsdhc7Bw6qGMWS6uDVI8Z1H1Nrup
k8oXm5rAQQuGOJig7+6M4NwYLyPoPmcI9ZHQ/pJjf27dF+q3h+U7/J7/T3+xXiow
L3Jz8bvTklvd/wUot29cpQaRSFRsbxgEa0BRnFEMVjwzBPHnPOUjepIC00oyAG3C
ARQRjiUZL/TWOFK7dc6qnUtHGJm4RvanZZgk/5Vn5x7OzWBan8MTK3HPpjQaAX9b
k8FrlZRkPCIA3yNJntycvna83KFG6UcBhAD0hEd+8WFnuxFZaiFeK101t8sXeo0J
lZ32c8MjHJpddqPPgCYUys9SkY4MEcUR364NXU8VpaEjHHiNN7vaI8hKlqK9pCZo
sm2bNQ8U0CNiXd64nhf7EZFHmKBnKcwwcpCWVoN6rXZEIhXtlcFo2pfqlGHyxuyb
9bPN82Uun6syReMcDcJ/GUtUjfoaXZa1B/1apmJ6s8RtggOPgpyZDM1lOXyeEezN
OMw+g2S+EYFInFlN3J0XTIgn7mtVQ5jDC3SFqjcPqA5kxLSc7YH37JB23IwpAmea
wgGW0N7bq/agx3fHBo7CGSzvwz15nVoGiD1sPlriDrW1WHEgPYNWHJm15NREbtHM
Fv3t855DgSVF3+16TImL790DuETDBg5G1rYfCdZ3bdEb3PDiNO47Rh9MS+EZp3lM
clzhYbLhWHyeDsPmqH/6mCmiMFrrGHqi4WvB9m+AhZzjpqQzhZREn6BaINsmKbab
K/S6r7+JdKlGv5WeD2S/eW0YegpVWiATYP2bJe8PFMDM31uvsWXnzjfWjnBF4x/I
KcZURaaVSs4s5mZK+Lt7PANzL9kGxX/z4Qzad6CcIy3aXxg6EajCzyw37/1dOo+t
ivm8eJfhm+LYOO+D2aMhK44Y0ejkSIimg68PcfEUC8D97NQmFq4/M3fl/V/SgKM/
MA/QU559lGdySYk2D6Mp3xfVwgoKgFDk+ZBpd/WDsBT1svtXPZhlIbfmIms4awmv
UxINI2FLHiJTSBLKEHkZO/N9zY12vyu9QvLN+66S4bVM6B+ObLIDiPqwMVEIjRSL
dg0yc/WJ8GHQMUNi0dEb+rWO4l3qQtKXL5c+PTEzwjX4A/M88dIpPNUYZ+SYAbN9
7iFlncniZH+AY8UBYNl6ZipbvjypY572n3RSK4pc6ImYubx+jjEoq4l8+FiG5DFB
JXXuV8H7HvQXkq6YD4w4Pen4kcxg051PUthAjFAhG2pc7ngHBCmzVG31Fs4Yh3Dn
QY5RzkuuCy8yOERgig21HD0F2Ew4z6DHSMODilSf5wbCnGf/zd+mx8junv/5pyCM
2PYdhp8QeZjrveRQlXD738xbV156q9gItbPxSbqT+gqPpc2ZzxtNHwe/JvgN/S1Z
303OeW/Uqmmg/TNuAg/3lEwOpgsSJB3H+e6mu69givFaab41eL1cX2VYKfArDcge
U9hJvpc/tgb52rY3K8lFCPMWgBQAMsNqgGb9YMduqk+OHDs4ZKOJvUdZ4V0WD88t
VzkwUyFCKOi3ds0e08m7CTNG4hTP/uKWtQ4FXpy0GLOleAYW+fO7b2ltwKQykPds
iOcIdS8pzrhgRLB5CE/BysQ9LjNPt0ZSulcqj23+05Zc3zImHtdO3RfadB5ZOJMD
T484vUY4/eEZhqo6v31/D+52Vs0bqgMfoi8nVsz0RiHufjFq4G/MjX0T1Iv/bhhG
oSDfHvAbZX71Q0Ipl1r6QRf1kLVn8WfpUYQ90Py6eQVyICB+GSt4aQ7ZFJZaXsyO
76ZZdbtkEPkyCj7ljmY8WojymxR/bWAIS6oEfhN0Ib4wiEZAezD5l4rSNaZnK0S1
QJ4R8TTuJFVvFxBMQGAQNH9VMbQ5tVBFUB93RPx3AnqWQE0lGJ5hTS3RDZm8+3DV
07/6l4wSVqvZ+tOHMjDO4F0YHaXyNMBrp90XGwP8wByAJZ/mHIUVZlhHvSbePJt6
rZsPqUhI7JCFEchp+VtfQnmymmXwAwrKFXIqET2HswY184YgM9fE43K7WObMCSp/
PTDXvjkNCFOzFAxCMvi5MsRwBoWMDYA6lhbbxlfqMH7WtgwmSA0Tn4wnl+7GTrgh
TpftcCHZbUJdtJVTuL3WeKcfRGXWGmMdi9TAdVTFUHWn2REcJG+ton0KT/eLsrCi
cpn2WPJ/YVXjk2KnvtQvJjwY6sHlTkB+g9Io0OKNH032iln1WuTYy9i0kTK3jNOy
/VgWYkPJunv21RaTHCUXNKXPe8lDeq+bHPw6x6Ngk6XrScTQG/INZN7BwxZ58DDB
W/bDoHg6R86clM5baH1ZUQdtMY+hTLFhvjpehTyYLyjIcs5+/uZn0EDnobXCMdmD
FGynsddK72/A9n9sVqzs3ucnccSlR8Jw00TDTIJT8beefWQGGVUTc5ofR7eOCDDE
L3Pv4VaTREK1HUzWChY3tu1CHJVoXBdFC55rn5V4NiaX74XhiaZ0LbM0wzOXbTRl
mGLdergSbqyUBEvZe5B/kK0c+5BjbpaidizZJ/Y/RhJDhZynMEcJ+emc/AcH5zwg
flG9YUfS/5VrEYn/0r9l8EcCHMCZU/PCGl4cPwJGIw6nJDDHQLM925QGgNAoDl1F
bNujytk+cKh+9qFel2q6IC9dxZ+lcjcZ/Tco6t8eMtcTV4L3Evb85npPFJR5MEfo
BLh95s05bfCUijsSQlJU68FBwCLibBT6VvAaWWvpiv790gJIHW/9nouma/AdjKyb
DKg222DC1rck+WnhmcG8Jv5pln1lLJynTgfqFQf2In/r0O9vKa2V2vmHn8X7DZlT
dWKRcAwe0ETrJY34b2cZOp3XC7lgtWLxXyPRqcoYQPJZTRZOyWwnCdOu+DETYNEg
7YMmUNK4u9c9ibboce7fUdk0BTA8aMn12vJJdopDzuv3cmXqxKSbj7DlkSUfE6/P
8n5tpZolCmtpsKElag6MqaSxs39+1T8pe+QBvdLhmWr/9TgCM6YbkyK9p8Wb07gi
m+GQ9fApnQrxTuqSTxmmeYV/VfiZ3LRbjz9ZlcMu7fNc1Q2L8mA10z3Ags2vZUzm
uF98I1rrGwcHcMs/1fF0pZXBDxH1RgTJ/NfdxzuzbexPLT+BrM+DS8Soh+/bSjsA
buKuS1pr/gWl5ehxFgJtQbvajB99JJFw1yP6nPJnra7QcPaV+kiElbNw6cxwpH1H
5QAdjN5lNwW2up85yny2Gh7D09vKiL9fNR2B7THgeS6MUbnCfsQH1aRl25Xy8Q3/
FnWfJp+cl+FaRLdo18mekdeUu9Ppi5SQuNMJovA+C4CR/oI4w3c6NlQx+99rg8fe
54VqPylY8ncUxcfKH1J+ev6PDLMo/pByQX7o+CZJLpUXQZH/oAg+tfmp4Ba9YzkM
6xCDYTlkGBCr++0jYx2waaWxff907cR86n83SpUcQzKVJGWIK+x5GlxZ5nQ23QZr
8DnqB6mLRiVquNbH3DKOqiarqkceNZgMw/oTdcAxf+fsBir6IjOxNn/8I7ep3hPI
kVEcKQz9jHRiCfffKG6mJXL9S5wx7dvcE3Zlj3SET1u1Ry5Xm3Vl+945ErQgYDOq
dTKeQmFCaAIGat7vQ4+xrfNYXzSYiVR6WHlpe+0E88t6QGQ5cVYvu9jVrz9n0z9Q
1jPkwvtGx4uVwDEVwru7nYAlTCH29UCHRzER6zV7S7ehyhm2zHg3p06QEjeoIoKb
nHVjlz5WXiVJ3I+94rtZfNPqYHCTizWW9oNxN/Ot47yFS9foYLD4Ngc+twCY05av
PRGC3BSSjqhhC+7wdkdvlN2PqVHX/O1KS1C2Ky4xPkQAcIhKaVogSWgBZOqWRR5w
0aj+yySxO+dBCQLbHLkvgr6eBt3OTaNavb+bWYKViqHGvI/WgtV3AHDiz0OHCojG
ppioFrZTzQaM2lLvUZk02NOlLzLiLk9lXNjh4Raiy1zRrq6ClaE9/TkPnrDGy2uG
YwzGjG69AenbzpLQqay+SRRvkVWsBHXvughztDmvPHSu+XoMD5EONN1rkVE6xi8Z
XxkZ596pWxK2p3xH+sJuZlHqrF61Yq1hK2MVtKJQ7iREj7Dn9KmppIgxU8fPWL6N
EifpqZIXQMO6JMVFsydRudUXcYHZ9dY1GIInlNvJuiSu5ZqbxPc0mMkAwESF9/hN
uDKG+zM91RnYui7XALvXuYRGMOb/0UhiTCj5k/OVl1DNN9B+ZiE+0vDY35EE5rXC
j0iY7dckQIvp6SiYiTF8l8HMEWTamh0Fboo9VjuQUKEXHC7T9y6ZPRXI8mFxEZiX
Lkl26BsRNEJxDt/Hd5iS4gTNtUOcgr5zDAO6aNkinDKysqzamrIrLO85EMWEAfN0
s+bVWLiR3rceIJ1YHHAGi3dCiAKtHy2BcPeybo1gN5/JPnPCK9YRQxWctVEz3qqi
tM96bSE7NtKoxR2ykE542K3VYpc6VaU/+orDT6npzKkwxb0Gdi6n19B0hhLlDhgM
aKiU6Ijse8WuDiI9mJuQY6DXwtr3UKB5rrlMu83gldA3FV4/B/JF8A+p2o2uM7tN
EJEqRn1pIZ1zzyunKgpJT92Ykqob9VY1iZGu+q4bAja5rn1BPnZf1DlbBLbOn7mC
HwYg0WwxL9Fp52OAsnXaTN2AHRXXkcnOxpOK3t1wWmPiaOR/2scZ+1Q/jPesz0l1
gIEjYCRh+qcUO47ZsrmkvLZdyCTBJO7Pp1ZHWNXA/BdGRYX+m7QTowrrdAwVBt9D
kCYZsI7MMUWJArcJT/ANsy3XlkmrNSjSQTRT4XWUueFiVd4pjEjMXZ/7l4A2KF3B
moyBXg2cEjf9zmv8UejY9kDW+HtQJlRiK1g/Uzhr9s+Q9+w9V6k0hdcI1OEdJxf8
czdYLSBjZiRNy7RR/cifycw8pzwRTEQIjnFbZ6CuX3Zw4xN4N2dEUCtnN+oovqFk
QZpnNNL2svSFORyCDWTTvjcKo8ANrrAvgoalQmemgMC2fw3FIEgTupIcGJSD4fJq
qqRYGDLo2bbCW47AN7/4SA7kseEnXegRmZxEPIlysI/PrFybOAtraSefVLYAjQKt
lBdsSLobuezdhU9PaalZIRorBhyV0ovLLnxgF0fKAGUuNTTC/94mQbuGbLjp/rTs
XqkVi5nS23lvIAvM8OkySbqHno0DrfuDlxV9qvYhBDrARX+ahdlE+J1CTeuPvVhY
/qEfmYNzcEapka4Wp7+2Y+El0H+ZVK9IGx15D0MWc4D3gCaHz7aHv2d7iHPfLygY
8NAdI6pMnuXSHG6xhTh+ygR+jjTt56uL8by0Qne6keB8tpQrMfMPc+IBI8YicAnH
MpwNluAEgYQTsEV/rWeDeklhOUcucBMnArmrfhoI1tE2DQQMHL5opwDOYIApAbNa
XgH+/9iVqDKpchk5InV/UjhcW9pblpqAJDrI6F3Z+pp5VKHbgS3Ocnr0lmIbDgpr
JnPrZhPcg+psTB1k0m0YEIbrP6QtNwga/3p4nuT8wh7A+9Y8xOt7ehEeOg97ejWB
wTdoQ6IJNBohWa+mFrgoudEKHy4OsNoP20pUeo8xlgVqsqdUDKRKS7OyfRh50OEQ
kEJwS9r+r6O5jyQMn0ntecXazj5idFKN1nziL3yne3u8NaSr71tJwTlSZmWv6YYr
g3StQRisBseToc84BU60s/E/a/rPgUZbiElF7VsP7416hkpq4tf7Nh9AO1ycPwd7
no3pUvzm5paDNdDyO/qyqsf0eFs/5SXsA8V+VVVco3eJMBadyP9TJfypnVTSqtT4
XDx8qO4mXzTIxUQ2vES4nRXgSfS16ImtmtTgt2EesKmzpV8ciJqLIHLUXQ9GXPGh
kVgG+Aa/uIQpibbKrt8NTycAM27RnaXBbBb1L3sD4fuveR4mYPDLljCyjgQTEflw
FBRfbO5/FLkCnK4+sLrrXx6XveF2zNbIu1HopBolDb73uftNOS5Zdu/zr6PTJ4xi
OpwUUWbcm6v38ieNG3ujGSpCzvKwuDp6am6X4M/0VWriivEF2YhizfieSERss695
B+ppNx535Cp+esSGGzqf2T19QfOGs7DMQheJo1Ew1UGWlbGAsmnfUmXXY1be3bTA
A0PcqpK8YbKL63lyXbkJt+wFEtJvjxKXy2UzLqKMtLFGsltOQLOUnzO2LxnbpLKa
YwOEiaFfT1EDs8/1gA4pfOBVuEoUsaocaeCjfmZlS9ey2a9jOM6hBi2UJ0x0WNVr
UtcMPssYu9oibKbJ0U/eC4HaAVJVQ6sJeR/xZUJBzJ4jwLuXiwS4B66VFQzhF5eh
75++R0cVHB3+E0LPETdRbJrzW17WQw+inbWobszvmoNXBSsbLzm54+ETodDuGkwY
QWLXQK3VoxPqoV7Mwo1Pf3ebIIRfGCLKPeIAIZ2xzmwC3x8/hvRHy/PrcToxjsRz
lwPICNQo7ADIRha/xUsrLL472RlcdUOB2bOnaD5QCP2dtlvS+9DKHS+cpG8/SzMt
ThbEa50NcL03Kh75gotgqQ+SJuLhGzGvwxkEtUQaJcwUuM5g3LqfaTfcxNgmt4l+
37RACo9Rw9+Vk0K08IjVK3NlDG0qvcNjrCE3oIYRh9o0nLRrcgZu2u+LkhuUu2RH
1NkRmRIJLn5Tpasfm3PI1lNdHP5FNLRnWTDICLme2asjZnuV169YecHvY4cqlQvH
wdichyn+rHmxQ9GpOvY3tcKPM1enK2Sa93fl9aiOaiHse2ctVoq+UATHoXeaOA6z
frFPcSI8Nu0KBhiG1FMW9ESOqu8fTllQAExGDwPftU9XLVOi60R1oZS/1Y5ZW2QB
2B4TdOn0JUS7+iPU8/n0iyCDBkADzIl+tqDvg9JRX+h0C61Rx1Snn/eY+An34gEZ
kQEdPYufJ36IIO6G97PuqxAtiTWaRDrzsHrOcz3l0JdGey7pfaCfE+RtVy+Nq1LR
yayvYyMa8k+WkpWjcnf/9ISgXw5fKjHZZdzCFoR7jO1oNJhZA0Z0Wbit9RtkDIxg
e5s8kLHpXfuJC2YdH6VedMSLLY7Je1lYClgunm14k+w4jARNqcRNGq8wfMPa34px
oQ+icoKxQF7y9nzGVcqoqY4zpQOjdAe1riKm5i10pOoH4f4PripJe30Q7ZBSmXq8
M3zDot/pqnQWoqf602whWWj495qHB9h+ROHoYoBg46KNIaneeOpWbxhPYICIniOz
yT4JXPAG0orSRpqswY2VRxVQTGwraUMOG7OLrCvig6XXexF1NbrdYxHneXpjPXYB
xBKX2kZNNb1fVldglTwqmtLBzUbdtDb7Tnlqcng1ymgvxDtKSNDRIhn2e0R0CAjn
YLFs3NlCJLH/EFvcY3bu1Z7xwaWz6Jq9lSeD6oANy7N7SIhAbuHBc8IYlITYKSYl
IhUxlfSDFFcNavMnS78rN4cEul6fXbPMUTzaVqdEttk19mNCfyTawHKQXyo2uHCc
Cj7Maqza6OaQ2jzjunanxE7uKgxiPRAl5V3leEoZzO7B9u9PgLhwnzFG6Ql89RRN
qrb9Up9h/v9uUY+3et2xsoszDgXgzIegLgbTDRUjbRKJNsjmENRrjXBVRSyo2lkU
ZB7y2GIENDDP07osEZyMMU0rk77HsJtUdNDHDGL7jh6EwCWtWhw253eC3g1DaDrj
lzcz9J8c0HsmoZNXA9Vz4D8clR67bwheuHxZU/5n1Q5HTKENC/DJZ8xMaW3ePWpB
0p4qx/g9a5tPFcW0H6BNM6U/3GZjrrSlJ2oZ4O/Ia/LKKxGnonb90AlIJzDSsEG5
YOsXDUrySlhZWOBgbi6LQvQ0c1FIHbT6GvUpzDod23zd8OUl7iuS5kG+l8PVMxBb
GEW4irnVjwQ1qnohrEskoo7zFle1kiu/vBPKugqTbaxYd03DH87QWCfuROBVI9/3
jfThUIZFHSqbiM2hrOwFgxFDQnMbjObrvBDx2DNUiMfuM/FJjiXhwfq3Dz5rANgo
cw5NsPVa88/TbUOtJSddcsMjFh6uxFyXHUCzWYMxq7CuKRgOr/agHrC9WShvp9ae
GBY9IHA9uWk97KJj3K1WXkd2kBOVXT1fY6x8F0HKT8AXleWmuCwHjOLO4RaPhH4y
gzv7aCjJUwXJ03KhYzGWrlZJuYWfuq8acgJgu5vseXgry56OTBx0Ctb3gbdiQJWG
wnPmIAIrApkUGnu4oN+HAWKuF4bWFQTHBa/CpD3ccMcKUkbnHoF0Rm6yEsthmhGg
ayoma16EwrkmMog6CZE0Y0h11SeU6w3oENGhnib8tkzjL7nau3GLYDJF7EsACCHA
XTq0bm35M6NFWAggnaUA3BBl2TAa06pEYqDvLbnXefxk81IZ1tOtKnxd6D4B4oe9
UmXfkaLezJLTQBci0+b1Pdd+eeaa1xX+ip5l6uusDyd2zh1SGlkC6WNJJnm7+7Ce
u6udE7EtjCvQ7JheJqAI1npIPbua5WER8cRMVPJveP/TF7JPlez4jNlhs9Jo0Rk9
pQMv1LJlOdUB/luej1HG5vpPxW+X3O4+LL39pZI2e5uTUTJTCabWjEEuwlpR1KD7
MtZQcSh3MPQBi6yuONSf3D767dZgqvBWe3nw6EH1Fyp1S9dNRd6FsP8P5ZUQmzZ/
lKO6R8t3kzB6aT0ynfdU6+RZatizE0kH3XrX9bcgQghr5ncOh67gTlU6+6J6UmQr
dMyGQcdHuyK2ndhqSrBMxKE1JkyakKN2PRNf/Jk6VOYMpTs9vYR/BU2ByzdnrYDq
H9HUaPvyYSD3b+GMWU9yvbzLKcrNvtbOzi6yJy5v6StIkz4VP+VWQAjxJqce2Hng
6ROM6VvhJJHZ9xKHgV28tT6yTgW9Eq9wsbfreCM6p9yX3nZdclxu1kWdFUq0Fd76
P3mfZAR3zORrcLLOm7jkdGBKxeMWnfdcndq0jD97elGZ6NqwnZK5UK1UNrioEAJz
FoQU1ZcOixUoi0uReum2LNQJmozmet1mWX1Ku57hSSmfbtIKVaN48HsUFZrPcYP7
M2NT1KkGojja7HyFc+pyPGIhvbtxwp66NRZrrQK0S+O2LEnpfxBF0SnkGXGUXNL2
R9WkvhVuYu5xgXqvy9ilAMFVm+I6WXhzASGFCZaftUVpCFNsG2Y4sQePrLWeJnx9
P2iD9yEMNbaank/8A6PHHbXYSmiApDVHqonlHUVztzpOENCEtjZNiXxhkFdbJUWS
aETjvbrre1pVK+/VaEqvglJPnsmGGiUnX3LniL4aj9E+H7gMN224HK0lj4H5PmSd
GvAgq2TcCSod3Hs2WwIRr9tRDr8Duj+7QIb4hDR1cSlhTt/NPZcr4Gh7f+XVYXkD
pVgvVdoMwMLWRq8CY6BYqo7Yl+tYXJOftgYuN8DqWcvzp0aADOSOYKR6q4YnnmKy
VjISfXTUW1Ggb7t4XGEJcuzAJaENMiMVIqUQccqvQIMxT74FqhsnyimVRxcph7aD
G18HGg1Evt1uMQSdpg23jqvDPLfwpVURT6L4Pb+Tc6iRtaLwmR/vHCtNIReulz2+
rSz7P3EWuZmspGf1bF401flK6dvpDxnlH2cAGg9gpjgxtZFwXx0KQGVnhCPGDqR+
MqhBaLClZubX8g5J9DamyJlWF+jY1DYnXl4iScdKFRhopyZTnuKizl0y9AM+T8Gm
qSTVnxh4R1fCvFGhPFdv4L6+ldUQTtilnXUwmUeApuAjN1G0eCAqvLOshAh8wlww
gvWzh7aWd38qtNSsIywIVc/xMyWnuFga14Xm16SaIPVoWKThcX0CUcIWJqYLerzl
S+ivzwOjzBC0waIUDoj7ezY0qeWxHtVKYJKI/puvjtOQw/ahS5Uzag7X8rN3YmyH
Jbs4/Sk300sJ6lGViYjZ09stU1u6HNOGEAKfXKlud6pCfDrCyQFONSA0tpFD3Mco
8t3mNTgUonXyg5YgWn9qNGITyco/juYiANJiwD8i82U1iJ7NrocbmHpVEu9yBg6U
eL6UKdjzL0JeHCG9LCL7jiSBV0sHpu/bGVuzpskyjo0OTzFpiIbkzdk9tds+4TP+
MbD79cdZb7t9hIOm/osajeR3gQR5FPzqoMAOqfK9je5sQHD6L/cB4zAqT8IroA+L
G1GqFC5tIm4slFYiL3FZwfzFfoq4z4Y0vfM0CJP0/W93PQco1Lww2bVZ5qomXtLF
MG5rTvZC/fEP61ZU/pReTfR6DfmJyqexoFymb2Fa8VR+y6k6xhiOkxOYc7f9b74e
tzlPR5Fpdua1PhClDO+WH6olcnzx0V2bQBh3KSNzr1E9UW7KHikCpjAiyOwPC7Rq
ErQORzul/LhpmHqiDUaKIhtE5h3WurFui1GEg+8Xx0g1FjvF98VIJ74WkP+eGzLg
bwBuQcxNOiiIk6SoXb4fT0kGfvRbUdrGkngczkrAHcKqx/tn7JpAC7E39KLGFwg6
30hipIQXv0K7lbdVY0b77vhCw0bVmpVmNGb8jvVeVVsZuirdSxuJ+0e+7Q6+sGHh
FqZ66ACtS0PtwgW+xXpyP6opGxES2/LEWinRMPZFs2+TqHKlOpRsaWUf0d6vz2/L
Cz3MIlfP3mNX35P76e6qTQ+idWLr6BLGegN8bsTGZ6oQp01hrasHWBxaZZUx/8X7
kt/KbrrL+5OnzksBZZ82uIKcSehqwnFMAS0ryhe3AKNKBcl8bmEJiMU4/1l+hwe2
SKFehFdK8JIszWxC/6Fi/TG50WxhvehNzUXeliNTSiPrG50Yj+H+gFMKFBt28UpS
kY8w+0IiQxNeYVJeczBjDU6/9gwYTeDoV4kZmArhUBpfVFnae5FHz+btryd0bS02
D41lO5rbXvcsAxBMGji3Wrm1GIZStQXnbGA7axLpxzj1RncqsH7tBvYARdKm9wpC
n8toKcu5omhnFwh0gFsBeUTl3dtN8h/slzPZM224jdLaJ++4l2ZR0zukWPxUI0ju
VaTPPFsMWJOc5IvvEhKwwV7bIwD8CR5LPUcXXRkxbdu5jWYZlugBY58Y05z+V0+/
76RB5Lq/e72g65KK9PRUtvecfCefRmjYRwJJPHXJ5iBWCfHmo5D+iaEp2p5tZCM6
IhSusYeeeFfIn6/MPyMvrC3cEMTOgU7RAZCW//20TFc4ZhrMldiw4R3zi7LMijSI
iYoHwqom+AxfWuFmDrAhIVxYW3oIq8X6LhyLHIVq63J11EhoyS9VQ3CBxde3RJOp
QrFFjapX5QuOAO1BaRb6SMQrnDBPgXWVxjMZ0bXyujemMTPHdHM4oSBzHAsH9sQv
jSrbIlB7L4Hbc6FwITmcB8K28xUUNY7frxWZEZc90ek0PfMBizfdoGTwpgt3XU8Y
6IzjDFSvbsG5mRxZFV3b7RiN6XO1WIBu3Am0Xfy5S2NlktphKqMZHLTGnD+0a//8
9bRUBT4NEMXFGnc4StAxy1fq3lOrJmjmBUTmSFyqZ516eAATfwCjQxF5zOboVwd/
0YJPzAFGvI8zYYZebRZELyqDwXAJ/cT064nWdR8Fl/v+NX9AKfENDWecTeqn522T
MkH7SUog8RqjMCUlanuXRMpeRsD9id3MI7WIdIivjWK9yErIh3qllOVIatRZRGNs
YW/rMEXkV9cXMlD6Ogj/G6BJLdU9bCCpfiMYlItzXdBc5OCuLMr764OkGt+v/QCZ
CnccEEZ7fp1LVIjSbi0C0bdLWLDmkZliCaXo/YDLfr65SIW9mK3dxagrKwIJLIUd
u7CFQJVJF623EDZ8e5AmzNdmDUmPpFEPiAts11N6tAAkUPugj89I6mKdoIfvKqN+
zEcVOfj0BHTuFAQLo0lTbUbdjSkPHvR/shUfjbVbwxVKQmTt4NE5WpJ1LYS8N5tl
/cfXKD6kPcOh5nLuS64DUnzCReptjtPVhYzdJ46WLpjGfXy7EgaeOuboRQoQqO1/
yrZL6joX7O45fE3aDGRQMvQVvLB2oH7NcYcGXP1xLo0egzGQ5ceSF1hRMccPL5Yr
/KRDTpv/gNmb8B2nNy41K1rfcwEs+NCxswaxYShc3s5SQEVbyWV76Hs7mNSrFKHj
MTQj05np/7fVBlyQK+PjMKTGaKDWUtDofyNKfXXCNabK6T23nI5VXzL6oYEwTFdc
FlQF7LnaKmE0aPHQSmMO64M0xtfOd9fNKyNB1T83sQepYNK3d2HgYFaxPhh3xQIW
Hg8hwjLnEdD8pmmZ3gkA7CMJlftfPCwWVk8Lg/KEzgzlKi7Mw4NPSyKAgt1zQWen
43LC62KA1GkSqBURd21XjSVepE7c74rhVhNBpOZwzkhhiEelcKCXq79NLy3+D6QA
k3SOFFQaL6bh8WezQpEau8NCB3TU+iJffUM0D/a1clmJubOJRV4Y96KqX3eV2SA+
HpLqhRYq356oBaexB26pL5u1nK7iKyZ9TveV7FVHwGmWbkwANWcXVHGMKQAslI61
HsJc9gQikeBJ2s2WcOJBkSJKpv0IUugHEI5l7/57E05xQRyNP6Dx9wlR0PRAoqh1
5TlKkfY0ArHjEh9v7utcbu6T044wIZz3x6exWwjtOjlvSC6gxpfdjMvaqWHjljKc
QzR2rW5ehh189D+YTyYFpQrHJKAC+V0nCykDbyRYNLte9m6tBWozh+LSglV0hp6D
DdeWBnj4X/mC+tLv/HlMwy+DF+15qbjDAoF1sJE5sLviU/uy06027H3aHmti5PqX
q9ywOoDdgTo3ippE8wVQ09K/lRVgt9qiJDpXfymtTmE4G3X7ZTlHaE9bbscItegE
aN2OLbENhAZ6SVvKQN3/Uxns1G9eZXHN82p0sBo7X9+VtNIB9yD0FH+4iJWTK/jV
9SQth4QQ+ZWedQOxTVKqLGD9rUU3U1R4mShW2IKaWQq8XZYrmcs8SJK1NCT9Bw1M
g57AuYVYfEkKOpwRYPXVuJ/cwhej+NCDX2rIK6CLpH0uPaXoW6NV9xCN7C9ylDDp
gzY0yW7SRpJRU+peO5xdJKl6Rxf8K4zKyOh+G1zk8P/9AvJya3bboRDpm19gfmXt
0VEe1psMQcn3t4gjaBAnY++EGbBokTCQRJHKEX9p/JZjGLmZF7NFe2RCeh0T+ncp
W2XOB3TfijfzNWg24lEsJespKF8O6odQBVpZdQkH3EXX+kH2f8tvZQf0YFRIsiOt
J9DDgoYCbg9jNVFNIuWq8iQh328ndOnKDjWdaY3g5I0rvVnlsxB4k2dma537LhyT
i1/3N9TvB96oUwKTX1h0ce93pW6MEGHpudiur8krBG0aKBujosD2NAf3zHJZoX+5
Nszm506bYjOt4orQ7fjUYyAj36/tqaFWKpYJmgqs9uMt7NoGvn+RUD1zy8IqMeXx
BVjiw7vwJ3fZY/BEuM6EGHdLtDu3XAQkGbNP0z6414mDL0LmeOfPUZNZU6pBDSMb
ILdhPWh9JwDui6u+5OprhvHh4m+g9pl8sMlFPpyPWJo8RH+nw2aTEqHRQH4yNIiD
pCfF98yHSKu5rJQqYzUoGuyjHd26S1JrtsWwnFtfLvot0vbOwAxj0j3opsYE0ijE
CZRB7K9G2+vmSGU0z6IEpSqK0NtHBqYI7x+JQAPmN+ZlNhHLnqTeu3nm1AaqQlEe
BxtyJ1vDlGRM8dt9lpyCyIQn16EBCAqpnlT7/ANVeqjkLB/k6n0TrbCHlaj2CtTr
zTPjImoRXfyGsXY/r4waearDAuvFn4gz10vDBi8AJloCDFNsK8YiLuZADhq7+AaR
wvNMtYDGtvS1aq9c0PjMSV+mSDTlJly4FImj1dPlq2sNKINirIyoq/iBl9pTv+JX
eWkDgdYuGrubqN1abBup34oihsL2qdX0qhd7sNlcLHzRnxMU3h4gbTPgnuVLLl5d
VdmCmFY+4/gdNYa4PsMlbdC2hYxbF2GzdIAnHPymrltPgaSM3M5ctsiAOMJtvo5S
XrIwUxXDdLKCEc3Lts3Ef2jNIogcUPlk2I1hd7DIP2n6tUADlwvYPQU28SWuO79/
2wN1z+OSmCYU/Xa8XKQDLtau4V8Rmdgrb/ySud1x+3MLqf/w5XgNHQSYRx8bRpOT
Qr/JJJJtmYON2CArDah/dStb+/0Hb2TYDlSPkUQ+VOHtjtAudb6oTtz5deGEy9TI
hEmeV42DrD/GiA5MI9hRpQ8MqjBtd+3r4QGjyJJvY86h8vUEsp2wV5ReAKYjjPlz
/3o53Hs4AkMOs9K8T9fCuztXj4GlUm54xrVhETxu344jNWdyIh+axTTNY3ZdLrWr
xFLF8tDhu2siXYEji+gqLpqOhSlAd7I+DhRR+jqECm0OQ4ASLBTDA5GmXGt/kc58
MYI0dTh11BVVsNnQfJ72uAkl6b3JSMtlqsNUqqwjc+SBM4qh0n74Q96tpX58zP5w
17b+XypUFOYM1bnENet5nSgPSeI9TOUKDkK3PuLg45tcEM7YjQleok6i39dUSv5k
GGfZSAzB2fC3kxqYZIRwJkJ2FTM8o2ewX5giTV7vW+2OI5Anbt0btmWRR8T/SgHy
k36gnKppM9bHXo6rttQpcl4gI/HiH9C7Iw+4xI7Bg1hGwBEQi3PZdNmwhhbKExEK
ixQWPNiUbFJF6dq0cgFXsi233EnVQCXC+UCi1ZlviGTwDFIBsYWj+PoefUhkNMqn
q9DSS4mz9Z/CSn9kU2YeclYHAV4v5daGhm+89+umLCEgYKYRId7Sur9HedkxGu9U
Jz/qE4Hfjia6eVCeKhxteq+WNEi9skiwcWtUyDOS7t45eqUrpfmVk2iFIyGhnxK3
A9pVl4s+nxYyT9kVffxbpxmJ+czypZz2BeTdEMgq3DanaWWS2t7SBaFyuN3BpfBo
a0aEk7f3pyvyl3S0Bbq4fvq5xhdj7n4HY6tJ8jqphAiyCNb8ATZbVasYvjQU80Op
/QVhTDH72CN0CQmu6UDAznbX7zwpKzEdIILWHTWhs9qkUYVTjw60ClAMQba/mP02
ljVOAnxz2STP66kfAmgJFZhYuYt6rzUyh2Fg6u1eWdBAkppDEEjiX49HL27CX8pV
phQz3jsVdmLE20eVdxoNESwDgqCx5smd65ORG1DYQzPWgUIHt+kKn3z9Jku1wYvT
hzdHGf+l4SsdD0uBsgMJ/o6UQBtp6x3I1FIiJBWAiJVdzwkqtuh5LXzzHaHDJ4LE
S/D9c8hCHA/Tr7RJ/Lk87WERRfaj4j9pj5bzWgDZaq/G6ADK74Y12zwI71T3fzwx
Z+RlmceyzUd11jsPvOYvUBXi5rrKzTrsjN4pG28wbbE+yKQGdZ9JkYKHkIaL9stB
vc9LQ3cZ8iqUi0mwl1vxufAkM3vvH9t6DBKPMFupXM/k0rvoaj871QhLVuKOOW6W
ivR+Z88bvXmuQWQEyyqAGCtE5tUk2ysfeGEYSJm9GOMYtawMYuKXm3JsCG5iLyCJ
MmSK0tgRVz7V7VjkvR8qpn1q5qhGj5VCyVg14oSRTt8duZAL3rJWlF1Qe6FostqR
4BRqlA6ijreBOAaQpRe2D+cyxG5Umvl88bI0+qCJf7FRYeuVLXHc6nFtRkYqszK3
YYHri727kovx1pKRkFvHUmZv7jI6Kw6b0KHxgW1KUjXf3P//yXJ1mNGWoBexVjrV
c1hKc2ZkTAvjtUCnO8KNfJIIjNrBYQXsSSV/qDaU3yhJn9HRlAhsVYD7hDd+SqXt
9Aj8zxMsSfgM/+oqej9IXB+sslqfX0mM+9R8CCK7iH/NevymYgQUnDTpO8TfuHsj
5528nls3rAUXWiyZw/Xz8ATHpbGH7H+02xt6cph3Zv/zjERjKxNo3zNdRLeZEhqH
RLXEKIy9I/iiWIsxcbaQ7hGiK8ZMNGNzeI8TO+nQlD7j8MwCNfXFU6vR69ReqrsM
AXjXUaeXEExSPBGoRWHa1JstXULKFcOcWRk7s1ftU5Icb7k/9g4jwb2E3Wh2PGV4
idq3d2dbGwEYf0YvQlnsx7ZDMhhR0tyU8VF5xDI9snzEf1RlW6v5o0iA3jbQEkLZ
2pPIRhnRhVeS3yzPwX4oKkVaL/u6SiUipWgGrcj0vU15ph1WdmTEV4GMNUdBGZEk
kGh2E2SGhPZcmH1m9wMQ/Wf+/lRJ+U9VXpeP1LEUgMD03yPzzPFCG/vzrzLk0UgU
ZJHFaDz61dJiR9muLRdb2XayH7dEBRazWWs8UdKTamhgYKgGntq9ohdZj9rd9OhB
3uWmnM4qdNYBUg/OgNXFKSFGKk/1bIK1jpN6FSOy2aE8dWHhlj+zv0Mj59qkwG9s
J3eStHuEB9fr6O+9rHZwmOu6LxRislkZ0nMImcaydRsH9mpgRFk838CwEq8iJKzy
kt0WEwpbbNk28TwWF6m9w+4GlykzyiVOqwC5VGe4SHrmQOaLsW7OUYaOoq+x3zyl
ptSM6ozMlunkCBu2sGbEBjOhfkeJhYZsMBs37neZEvl5HNNwoyNdjAy6U8vA1s2A
qDY1Vhn1u5vnefW/agr4Rb5GpXUmNz+m26neTMjS8kAshFSzU2Nvq7thV/57TvZR
ZQ74IOpC5yg9+eNULQBcKtoufR1WREqEnDgBM1O4kfyhmsNXerbwAbxJEz5zjfhV
qkb6IKLKRztceUEqONUZDMOdbyWQ780zLMiPxJvNQuxRoC0lHiSfcgUv/1oDbiaB
Ahz1jFXze9c3Zg17NbCukZznt6lPO//ToeYxRSFnfCZuMSyVNDGboP2dFdtqYIdX
cZWGBZeP9STDU4l4hUHRJDtcd4Py5OJ8xpik38RslkljiV02UDb9E2WGVbiPAfPw
65dlvqIez4/EJLqns5jxko6eI3fNRPR26YD8wb40GCFv+fn+C42XtY2bcGxvSmbN
jSiYXiVtDND6w588qrgeo/J15X9NinJbwq9pMH+Xg695PdZKBFiL6EVfPPJ5mV7/
ShJQoxYRUShQQ7M+10Uvdxkvj+PTDvBX46xtvvMX/GTyxdJnYjIAMWawiYnHqaZt
LWKAldxLpFFJeoySZapQUoqWKuOTG+RrKl80CwgxtpaHwp/MgnhI85GqV1XYwRFF
ndmscqLZ3uY0TFJgR94DPwHfFqS0ajlMytXnwqUmaokjAVI7TPYt/9Nsg6CyH3xd
cZITYXrACvosnoLpdR6Du0TKOCbWnlUTkEajpGX7AgsLZotqzvf6BmqirJ0KwaFa
rjUsIch5wyEXOrpUFARSG5gWvkU4ljHgkbZhTrbiPVbNNg/CZygdLu2CEpSqcoiV
H7/ssLWGYuVfg2nwaldkni931Kb5MG54o0uJeQz9SvFgpEEbWSzikXGgNZdeSpJf
XRx7psgUMGdSucPIESlZe7zi0fJ9zEoRbv41tMDX7ciFZsRbfMpY+cYzo4f5o7QZ
MGZQuQEHm0sUubcrO3icVHyi6pPCAuVaHZmfzC0Gfj/FL0xCePRNeqVyHFRIG7j7
SEwJZdQtdKB9ZSIRvGMgRUT4xTaZt+FEG/EehbplBcLI6x+4AB4WDPvaSg8jZkBZ
hT42Ystyu0nZZRXk3Q0izn24kNIQzt6uIKS6NwryObEFsGs8xSqWf/gw2Wzx/0ud
PtWX5wNCKEu1MMzISWOp6yTpsTXAVWimHmIToqc9yw9xCJhJasM1BaKOpoQfaoaI
dttzJdNHKtBevvbn20VJZnl4ths6LGOgPm7FQbVtSXJQTVx/ZxmctYYOnWDKTbTl
zl06fmDuzI5nleN0KVCUXEL0dPN2zs4/xyJ4kYMjrKevtExcXMYDXUzhfKMrrgRW
VhHRAbzjgfVraWCPLZQb7wdZdqsyw8V1mnc+51L2pR3pAducWhMnOrEpXP+Rzk2C
mVE8wJK32jfeiVF3Kst91jXBk961E4V/ZzlBa+eL36k6v8gQh3a+Tpx23OJV85Ym
JOTqyJfz8zfunI12t/Zq32qMFsUUTLS+hwlQD77UFPcZH/XcwkZBLxIbFLMJtEP9
eHjIE1t+nd7LjzzByWMz9hsKQuj9ILEBPougVd8O1drjKvFGa4v4ldRDj/r5f7iE
2LHJuXJW3Rm9SvoMZ8Aj0g+JMdXbz9YdhrteIYy0m9FlvJfxnUwFiEHIUcqGioQG
cRUg1XuO3s3Faxag0UoGhv/sY+2yEWZVMUegRM9DOX+dIeocvpGRx84a10resUI6
IHaKaGGaG4eZAnPYqpdqkRfrM4p2aI9pLtGRf+lqEFsGU65CdgtfrsGAzaTgCsB3
mgxHVhIkZnCyhZ9oi4UIsnrLPDQzd45xOOzO64vl2sLkqOnf/NwWGYCQr6IGgFNo
YUpbXAQOm9kzeBmppNas1LGTNt9hXoJ299eGlbqYuv+ewuiqfie/fMON+eeZpHF7
TqCSJiUT73C3qyVCQxJSQepIULm9GEdjA9LoqO4jOtu3oTSmgE4vEejtRQwNAdr5
0HeHmo+X8ZHBeROrLZwMRbWdQu+P6OChBnBkHrpR+1GNzIpZVVGOLxiHF87UvCet
YvhXbnUFWcOLcNC3KMkR1luYIjuNv34cxgdl4skjuWQretP7o135CwxKTZQRV8gn
ICehtJPiVljj9N2XpEpE9FmUunBrUg4Loyd+B7R6pl2MzgzmymbWJdt6EnzEalmB
MgLP0+v2aZPuVDpJWWwxRHjMdo+tOLWz/PY0cNTohsPw0RszGH/F4R2rWwccIDWY
QtVn3juhYLXmSI7LAeXLGaQBOfQ1wIvfy/+JOeJmcpm5ZEPbkLXDdnkpEV4U6yMm
B/4DxBDzc8fCWyGzcGqCVyLVYrWWzysCSpLk3H56dfg9AOh0bOVxckFmlepEhRus
16E+GGknGJX0+Lta2rU075umJuJUQZDD4+s/8yw71H7F7yYPwqJkj23+9RMVsuqp
vMoOsi6FUlJBWuKTsEYjHo89cm/eyY3u/xaCF28qor8oJmWkJbMKWRGlJ2kRMAMw
yglAikrDuCo4Sdz0oX8+rCNRJxTYmWM0S20trKhhMJV8grZdL713FymB/Z/bib24
9RAb418EcJd7unwpJtIVS1r7wLcc+JbUgfTtPFhCVZvJbD0mVgS+Olp0iDtCgArB
ZDcETPwLuHOHOc8HMLMstrC+0LkvHR8+puTyYQSrOM71XqG0friq+Brt+F6N6NdH
sRV5x6cyuTVGYyWb3j/fxOVS3Q5TddFP1zVZojF9eMDVFEN/Wqd/0nYG/ihJUuvr
mpcjcWGEBEsQ+4MT027HPzSHO6mFaaviYG5Lw7CtDNrk15emjjCuXQ1d0wU7F8P0
OjBEe85C36pS0OKak9V4RqlsieauXY2NQ76HtcU/Mvkx+I378okfLdMtErJNnj4L
zwSl+ytgpK3Je0Q+MUNqM2KuA/lJIgi9AjbAdtA92ApucQo98JQYCax5c/2MHh00
efuTQIF8sNfUinmD56u3/bp8sv7HK6vh1NsDjy5ihDg8piSVcV2uVgVawtGnQbuB
sAPnztmKjXofNlBuh9YDexfsi+cRDQcsqcSVHBlpiIVEfg7A+pyUesggf3i1ZFWG
Dcw+vtiaOkTqnVAG80Yms2tbG/nspOUnjDCY72on9r19zbXLl2GwEbtKgQahmoN+
EWPG8kflu3mjttS5o9XhlpJgYnQPtjauMO6JTrydqsRoUbT7nuJpHeSbWA/J4HX4
s59QIYdWy1ESWuK3GI0gTnGHVwTE/oSZGeSgpTvee/lJcKeosQOCvBQ+PHF4GUtn
2TNrBZ/7pBZ1A7XwIbXYpcEoGw6gvCO0kOljj6HRVChfPfegZ24ss7hOo2TagWTr
y38Ay649erewq75uFmD9uczw1uW1Osd3jtXTdeziQpfL/dO2xdt2m0SaPxiZpc1y
IT7YQM1j7/NRZJgVue8hpqqtX7UTJvhssxJF8wpxmUax2SwQVkoAqb3IBSiDkYTu
F5MOyt0eNk3JNAPTR8URs/UCRZCyVCijpTFc9uLgO4oVWI5IrWASr8XlzUJN/Ens
IpGa3B1+yVLXQjjdNMMpBkMqvuDDDlLAc9hjHVSqFzmkG1m6I7cOeF/nzNIr5lRx
EvF28Hg7kM/ao6NuJytKVFwLehi4/yoWKbYm2VAfFvK6XmlQ9RL7BmCla7De2vPx
cNiuCKA3gIHgrm0nkv+NkQpy/PuEfl07mo9gpkNz9ZF9XowRgakGMWhYQK5iS0HD
SdkweHuTofNVWs1w+H3DTIxRVWu651K5epqG4vAFb3lwgby+MYmsmo5mCtudrGgb
CS8CuHZfhRSKRZEsqslo0kyIb5fSuaVw5RuXyFjvJdWh7WvBot4UC4z1pSMdybWn
1IfXLExi+quJdtsREMyU0AxMiJuVuP7GZi078Vee0fCTqQ7fSK298R4V4oj+C4wh
cjpCC8vcJGlRCPxlgTiwsYebHSlC42NJErFXiKqnP9idfyFKLcZSZY/4uiQgpQbF
3BDhJXE4kYKB85jTB3c8wRMgKxKRawSJvfc3znUfuJZ4uA8llPyUTvMnzVHAW2Da
DcaON/pTpT9bNkwPX/cGzjcDXFr8/CJv5cVEgY8dfsfNukNB4pq+Rp244zfMGTSS
T2aN6z3WYaPYVRvL5KPyFLvqsFPDSrMWNuyHiO6eWpDDgzZeVYqZqHWVUpGDFFJ6
Tsu2ttwotvDt93lGbgMpCj09wdP4N1JlpVSJX+9oGpAk/8EIZmvu1aszvywq3elS
mBqHmXPIZV51fSKHu6pHaUKN3z5fnyUKGnKqu33Ig3PobuiDy7z3DYW7ttjwWHfO
/H/nZxzG1akQBqytPphlzshmuUUnQCYNiy1saXci2H7zyhwDJx4sCmkiM6Hx9kTf
jomcngH+PO/37W9O8ruJTAgQsF8zkXovP2zSP5roljK0se+KAi8tslmyW6uB0Vp6
Iw6LpfGOsaU+VOT+shqyhlcxFQzeegdAtcybx/UadH+6JtoXROz8YzLHa2/hTTX3
CdUeZMg33Zyun8zH1dQLe9x9rQ1ov6s3zrjYexs3qpS+56NQ/VWmHHzelydQDuvu
aKT5Od5e2k+o54zvjqPNB5aUT4Z4jjxZvo20uUczFXyE9qPMepCXnqj42DpwjbVG
FIjtTWnNyTs2IhubhKKo4OmNDhTnUhIEVDSsV0PzB0+PmLkOrbH8pmZqQQajzFCP
DdlRsAzvBDJYD0VRwl3grLAj278fIF6UzBnpzpXetMo29o6bYQQnGf6NzyYJnwDA
9NsAmcj/KpG6ITLnH5jnWRH1xPFVTx3S83V0LkelrBdySMO3KQaL3uhfLnLjbkFn
IrpfgYyrcOrn7lMpoM9cImojD+Frn41e0qxM1k8zc4SNJQYkrwLUU6IdAy8eysRY
fEMrNEz5Vxx0u3bKxs+5OalItUNGqTDAbXyFNvE2xeTGfJ3El5sufNpJEzReCEOC
ESKIJaZM/XK7UKZv+0O+wmHzPbSRXni4G65G98h2ZO4Aw9LJNrfNI85Ep7Khvhxt
NzaCXVbiXNa3JBdT7VWjGJ391/9e7xYOIUGM+vG1vDN1VVgxBJc3cTbHYXVArTVi
LZjzGgYQD4YDwnXCpvJtxMyBDJoo/KZPXaIz+ZwOEw2Ys3/Jlhh7q2QYUrHGyqQk
fZXnzX+UO1IB4UERbedAhCpSfmNPQR+ct4A1PvE3WKXY4J6Db6zgPXDBvgqyrKO1
tWCsw2c/CW7QdHr/aDNU7LVt8inhnmxuY/fbvwhk9jbvhel2isHt0oZKIhNrMlt0
CLuFiSq4LUCyrBS07z3bBKz4BZqHog9eMx0lNMdNM4v0Nc/kJEunU3rGkRoH3sXP
JS7lbeayXsdglEo19NIxMj05IbflLdgfOT9NWr/db+QeYNykApXkWBYxEkhDOKje
6dy6cSZFhzix2xoMAiRuIxgyYVDJGxYu0BmcduVIC/iIL/huIXu+hLRczHvy+wX+
4EdkYUl8hBNPtIAlmViZdHwTyLYfmIOdUxjpPuFoRWGzay477BoYdT+alo9S5dfx
KG8XIh5g/A/SKoqg3AlZdTmepioPg42lGdkA00iOTcGh2osvQRnjr2r/fNwqQQI1
4iL63eJSVqxFYteZ98Tki1fvLvEb117cJq5XuVS/h2qcTcWLD8yxVC509gNiYTIs
5+oHB4Y0mBohN4U5ybdGTvBc6AE2KUrTqUe4A1WFcZsVWEIVGwRO6mqmI7UBRwNu
6BZKG9anAS2nc1n+K/ogHYrIpVCQcxI334+R0Vv7BRje9eYSsB8iPQREOX/U0mMY
v6jzLNUxhL+qggIVGhIzG7NG+wOCJARj+IhQiJqb+edi7kE6tSWDROhmiE4oK1lQ
jiQIoZg8Y6dyvJmTNYSfIo1CocFprV1svKyehieZ48bwSpg/0BvlB0Yr1Wr0jyO/
iNHZmR1lgDfuk9bSdEW1aCElvK9kNTnsXRiMkXz4AgHQAvE2376+qi0DMMLiTeIP
6s6ZeKYKrPHjNQs84rE53MkXuA2IvR58/1UlJBIubKfJ52veYo1m9fyT9CJseYRW
wg3MJcp7WfLyVnV//d0RlZtamq1PuWdC1OtO4yp0mmY3u4mNauZ66eq8IoEoBrxE
sNkADnLnQeeLo0VsIa1ANXDmgoih0XSsDIky3tkW6qF0vh/h818N1D6AiKgmd6l9
khK1QAIQe5lv6GrMklmMX34kGDSiiAFwjmqvFqbBX+TBDvnDJ33yVOLembrPqQ1v
A6ZCag4WNFgYOob/bs0Nv5s3f+6sK2fN53YzD/7/Uq7y5svyHG/Ixg4jqqK34tn4
OvAH0YbqLOTfqnQhvJ0ZhnrBtQkVeTzTYgAYaDTaPccpESG+rO2NDrt7FbiH/DFU
4VLHM57WY+DlEHzotEtedlbJ4xqgzUNp3uexmRp4kll38adyzMs6xKgT2e4qmOIh
puCxHorHyQ9VvKWuKtEVyinY4qQTi+COqJJpMbIkJfSfxfLyhMK6FrejOPmw4K+O
wz2uCwNKdr0iVqHaJ5k+NWsgvrKdFj/mgi3JTL87tlbNg3KccnYHBukqjGoAmRf6
iGC+sQA/tCXl+6qVhVbTJb0kOhP/4KiBGZnJw3QNANUdP3VXfALnj58HlM/bB1YJ
iok62yRWZcEbVeXrBG40zS53nSz683ne5zw0JxGfiP1533ftZvfBA5pkBJg8A/z0
EC+KEe5cQ94hH8dpESeTuFCLNPidvNafR1oLnR9jyb2fmPpd/sAi5P6f1X3WSqdm
JRibl1+Rw1y6/lEcEmKFoWkSdBtO0z9TNRFzHn7moZlq5dzUY5zgJNtO/ZnuuNo+
sg+KZwoFI/qCsnh4FLrOi3TgKAt6FsaM7gdYClDT3XMqrE0aS5fCSQ/H1h+41Y8U
BxrkUFeqz8dGbzKgB6FoD/mnJ5gT9FzE3e316xSt6OQk+/GTnCnStM3/0pyBqp07
XPgHHfXscXDm0hY8QOgBFJsaun1sGrIkm3Xam+hkE1vKYQMpgpJFyFClYm0KtgWg
gdLagAW94Nbd5Ke6sla1HjXbVDVtM8sH42igyy6r/SVf7GFb/v2436ftf5Js2Quf
AIFfFEHCPb9DCKiJz63+c2uQhXdy/RyJNUnFdOmnWQYEa7HvfJqjbYxsknY1Linf
ETcKDRMJibtnn66qawnzLV2Mz+NmkgmwqHlbH31qDD+4rVcW+mUDHyouTB8Sqqpa
uPTs+/kIgFAh8ovOoh2tNyTtnfkafC6++gkr0mqY34itgi/+DeW1EekjVXl/AGqc
dLutScH6YG7C8jA9qZpF+eTyFaHd5VxPSrtxQhU7KzguDSKkhIokcnISj4HDOr4u
kyLiBGPHU0k30QfCk/hjUXhaYEKYmegxwB7ihn2qX8l9pRYHLiPh30HdWlKRpqX1
9IH9ztdHUcSClbK7B/fQwETPt27uMTGrujFEqW4J3ruzV+ZzsXNv0HLpHDgH4BpO
Ro+yEn8KekGuqED4cemYkYxjsodFwqVES0mCn0p2UAEA4FzGiHGszQasP35/0gX3
iMpoM//oJJLRVoRCtYf0lN5U2LvcCUATfnmWNPkT4Q6wVjF5VThldqhD/p5Jgvas
t30eOxiSRTkYevlyapnczJUgSxHW+MR0ZIJL/ROIQHFyYDv9fEDGxWvgbr3zT/Ex
2m5zEEjkdUUoT2XtBC5FxF+auVPAY3i8dbrmVndNNC3CFh5/AJIJBrKVoEMEog8D
PErA1oSVgGeBT8DnUCTlrBCsmAjDICpD4lJcWpY6HYqB4V9AUhkdSAaNUueE0RIv
c/VgvgargSMeUsZpmUE7drIpr9hSSoVhfT0cw/SuI9XFe2vshDQ6J9XTNdw+coVY
RtPZKPudsTlgbdHZooQeyC4Q9pAs/7XlwUi0K7SpTvEtEhGcRWZ3h4zD7UnHQoI7
CAwOfyUJSZ9oiEZjkgmWgpnEKZfkDLQJr0aWVhSvXKCSpkyYt36gBxfY7GAHEGwn
F7Lt5ZJT3hVomJLFWNidld4kQxf+ijyS0vTjCV7ljb7rEZzjsTYwGRve0hed6CLX
okaou0FcQW7XlXo1FjC/pdveXZt6QtpE2T4bOznj5fNvqHBVpoO6yb/+0fSC8pUk
M/L7MBYSLuYz+vGL4v7H1XUQik+n2wj5fEZnSCkiBJNDjLTNIDhugiaNL6Ft6Kgy
KZAXPMeHTuJgCEZReE5Kdaeo8yB206/G0aphrkL1Ag69mZ6ZL+GYL22HruEJ6DAE
dUHwmyFgZNUUVl7UpBfJUGcgutcazkgiNKt52Q9h5pHYRrJgaWwqAVC5GPMWv+vR
lMKLIk2ctGd9NTUwni6xu9+nZ+T3mdtHNeFOta1Lrj69QNQRHaDFQi56WzgyxwNS
V7MIfFhSso/M0K2WnaBR9exQ+3FbTJ2cj7Ll6gxCyd/wGRw6TQNaoCu80H/0JFG1
Mz0gA4tdwosSYuu39QIZKZdtluUmB+RlYh3iq0Do1rfxu/wJytCYTyYh37b9nys+
6sOpF5C5aj+CGtlqqynAn5IHBl+CyRmuYf7jLW61jehqB3UaIWRxP2lh4K9LcrX0
gJRdzMpLTmKPyVxT+NzU5bxglcZh8lfLZuvUTu7+xPldLlIyjMqhREDFZZ0tXzG9
G6+UlRyHl/J1RHoTHTRfUdB9GblrYhH1y8ES9FWFbArT9XHxPS4tt7bJ2QGd9uyT
fw2MiMivDlSexQRFNnFBSE6PenDjCr/bnmXZO5jd8V5R9fOHBcemNIZhhDJJz+Cf
gkUFL/3sT0w8GC4gChqlcyQRRis5839IKHNxGzDvb/Mj52H5ZPOrrfSXo2EVeSWC
LZbOoiJKrAaz8Grx9Psdz5BnxG/96v7+sgJoK1ephzqZ53DZjZNhBM7fW45HVgp2
9mfwR8Hs7mcjxUNmgmU/+4o2YEqz8pYKRWPQBj1qxby8WNZ0dMkfCojm9xMg8bd9
pbPqBhSHNbZmLdLRHUsLs+ndvAJ+cyKHwo34Edq7I0stFpQZmV4/CdlG3EKGQkRg
1zIY8ezkACUCBvXm5R1wlRMpuUwybQrRGCtWG1uAvAarYVwmBzglTiGIPZU9Mk+R
9a6vaAk/k2rScLDh39E4MA1S+US9oDKesmvFqGhvdPFjeDz2+uHTpWqJs27vJ+Fy
Ljaau193tn5WiPzZ/bYyi3y28M1jHx9Qdj9+XX3MHZm1mXmWihHgzcG88evt+vjV
bPOQA+FzJnh/DgXFpsM4imIhC+hjqaM2OQ8JVgeiAlAB73no3hrYnK+Lvr3uS2OU
2t+8J1XDN4+9i9Hv3M6XPK0D8Plb0dvloZh7ykbjs0ctKEfAUb4q4cyV77pxYuWa
XfkWp3HgGveDerqePEC/RETYneiEm+ag85a2eUVmToF8/4cQzkAkktwzNsZEo2la
8shTJX6x7ul1ZrvXJVsfzliGEI5ePsFdLjkrgSshbXnHRH9dPX2tt2rB5X0FRsVo
YV1+febg2qBVzqpeoaXIpDFIUNthuwMN9EyPC/0S3Z7+bMF/myZxrO3X2B3/dhD0
OlqrYVI9OkEkSLkfvX9MHsQBf/RH8FgF06lVVcRd551ypSGExuOsZ6qhU1UIV2jO
WFTWk6YHBVm0xw/T5Zm+TJZRoNukdIQJe4ewZyhZQUiOeMjWTgW1jZ3eRmdXEYOM
oWF+PJzMYXTfVqd16gnxDnr47YS0B08w/73wz67gCNtsyc1GuqV1JeZDODwD40TB
v3zFh5go/mfz2wgQ5JkF4Roe/Q+Nq94SNXrjImXfrFRlp9mlj6QY3S3IVEnGdcWs
UnKvVIChm4N97qtxZg2ydU79/bw86MGhU5ICLoTnT5BLQ0LC67tgwlwl4LMgvfPt
DuqPTevgCD6jMKKuM0qY+Sx9ztN/Fv4VV3rOS/arq9pOiSeMCmTIkzg5bNPkRsl9
PSlgvl5UWB3fAAwTyRZ/E7aMq9ys5lEJkdcqasyHVS4T1DNabJyoNJv6miLzZEBS
SPmk1sKIPoGR7x/+yGIwaJlCLqTCuubtFn3j/pD21j/On7fhbfLsX2d3NN4W/ZX3
rXmzzdy2g5cDKTVI3itwmQz/g/bVaFyKoERcH9bA0+LGBtIkADvmS8ZLkkVfOh8I
y4I7eD9O0+GPCD3XFjM/GiE7mxNl/wByJ9xPrVJk404v9ndpZyrfXPaj6tNXOGwJ
TY+dY8u3GJRzCAx65OO6NoyriT307qDrepBffkrTZzcRjdCM0cgPEyssrhakKXPF
KfMRwRQ+aHfcQrA9FswfZFMGbEnTtVTeXPy5M28RGG1Kz24+sC2DDrxalutRRwPq
MBUPsvolkeBK7GtC2UVEnaBdwZLaw8gxM8e72KsWSkqS8zdpYhilGEXArZEeOy+/
1Ty6LoeJWtCdTGNOrWYlCUKxK8w8xNPbgzFa/uubZvCMh6L6d2DjAdlEWNe6QLWF
sQt7860aTvwUw0LShu4NfhSIdcy+CKQovhqgHrWgWYD0npL3X32vklE7IIjcKr1X
6pfuK4rR1u13w0xSqiQCiWakWaTiONywgIsEZCVMptGEM3DaMlFcaR+BkUu07nL7
IDD/TbjxitArfWUxlliw1LdLM4whPIEY5jHIuxNXAm0glMbyBDzFpSoQxwoI7qI5
gbzsjDAxtGndcQ26d+Xv572swnwwS2/qjDGmfPvR/OszmOdxBq8R+aJSJqPo9fQY
9Kpl58HsJfm8Gci4R2O52vA4AE50uQhgI5zd+UoqkzXkV/LwXo2vwUqRh94jiu/y
+t482PgZmTR8AWp5KGL0Rdog7FwXxVGtjcv7wQc8u0V7ij1wJ5Ggnp/3RjkCfmoo
N4iAdEGrQe14vtYXCs3y3qXuwR/cGVOfDmHwsa1v00vbQbNb1o6+vV6+u6VQpfqa
AdQ8IpoMRO80rGKjlZY5M2kTCfegqG4IGZs1JFRa2aRMSMB+EBeL9TSo0NfC2LZp
/KxviZDAl69EcG8z80n2IICgCkBpS0Ow9nf2ZuD20MEmx/3Mct6P4mf6VusklRS/
6f3Z/Dnj3akagIkgIldeAFL60r0jLh1dPBSG125emmcTyYEpdjkiUvE4WnjLnpRc
3BLU+/TS8C+yiT7q99/gDICyhOznReZXn2Paz5VGla8ZrK0Ql16y4w/1dzuhGPcM
ApTIKBlTyEALJ2f28aEkL645cV6qVZlALbGEUABgqypRD6MuYAF7pJiCpsB0SO2q
vmXYZnrATO5auF0iKwTks38fArFOTi7yjY/Axc+lvS8tnDjzXHg4bParGHUVojKR
B/DujVj5vvx5IBuKZ8ZDTGF7AhUCdgXRLpm7V3tuUU4kQjJw6ZhCqy+D/ASMogyp
n76BwCI87h/89ySuJ4orZ8Gr04ZedstfnqdfrZi25QAm9Zm14KYeDvqfNMIlCE9N
qsfYP37rX57UWpdKa+Gz5bS0MY4bZKOSg1G5FB1QAmaPkAGC9TU7WPoNYs+mE7ZU
Z52PjNgMR5bdWXHxLQ8CsBIRStlo6cwiCDid7ZMmb33dRnObHQTAxV5cQjqRm7oj
My/aLN83WkqIHr1BFpouiXuJNMDOOq6IHABONg4ndHdwwjUqYuSE7Ql5R5+4u47d
GrkuTPHh49X4hstMapRDKg0wL/qVxua1fg+pnXDlnBKnAdxKkYjlZXgdVt6dfP9g
tFFMNQ5oOmalKu+SwALBx5jqCYME1WhcahU2FAc7RuGuFRgLOclVUCcUjhrlBXDn
BRS48g23fdfou4Gg0WoP1/ICuJDgc8e4UvMvY9+HRIfhDPVJv5Pf82eZqQ0lEgO2
WFQid2VmdIC3m02UZLDVLYv0Y7qOEUouOU99mvV633AQ1U3wgTechkkXPXIRNDPV
Ez8PkkzLOGMDI4086CL5f60+mFct/7soG/TgFLVkilC2un0Ux7RoTogaJR6wS1f+
XKsTu9V84/GmD/KQVDTaG+lE074Spo47WA/AMVgM8+pOqteqpkMWloSuFjWEA3AI
TgEe+zKrB1TH9ObjsHcpLLTF0J+k0o3hJlAg5Ch9CiVvkShe3wI8DhBsZjdIhvf2
mwZ46U4IN+M6CNlwlTnr+FqTmqqYyIHTJNe6BvJCDB6wUvII8thoOPMlKxBeB9zn
6DCeJBZu9aNyhJbRm60YukCidFcYjJOiIa6NMb1geDAp2U/NhIvuo1URqvo8bpfZ
mgJbSRITn/lX/rKIo1HJwh1OQzodFgHJ8ifEUqPtGlsL34KSDBd2BA9434Bt8eLp
jn4ER8z/BbTpiiGzgpvgGtACMuNtzw8Ko1XesFEcnnthw0CBjyupUg3sAcZWaYk8
Wsr7ZJ9m71ORfHhTx6QRcwdlXUtAKJqDNX2QM2SWhdF5KkfMQQOTqLUEs6zGGFMg
KIcAeCbb+D1lp4JOK6qKlyLyFFwgYFsa/6lcUFWrCC/iLlOEc+LGiDUinhoIZaWd
Rw145b+LGhS1vJctx2NYGgP7nLkYl2ixJz/KI5dYQ1K157Lh+/Ad6WlMUnWBpKst
7Q/OvrpBTTAnQKp07qi5PmcrC6CBug5h9lj3QKihKW7e9JzefsM8/ZagCkwFtnib
fTD1XYFHIK4qyMKhj4Nd5Ex0KK8udkCFPPNUo/dUuQ3dzj8sowLYTKerNSj6vD9Z
dH5mnqDZ1WAUHZVZ4YhtnTYZym5la2pzZoJEIsP5/7NI20aToXLkqqKS48h0vcrI
1UlH8rOSOlgT8XSCSVE4227t2zT6Bs8jaDDrUI63hQX45RL1QjgNnYMBuTfy0Txb
A/KDH9z928fYM2erhFeP4QNVcCwKzDFHXLDuxunQgPSnllV3h2pzaJNrKk/oJwgI
qF4kuGHW9dVtiO8me4nI3yrcbX392ZIWoL2PgfT9c9khpTiEu74PiVvxKgaHPv06
OPj+CXVJSIPayqlR9vrhrhk4W8+jWuKMprCEzurpFL6PIokpxtApsBiqgWJFCWMO
q0WvRZ9eK890fmbrnPUj63KbB6q1CModsMw37omElQTug2tGX73lYDXymaf95t/a
2e0L3XfOLhSvZnCTA1/3tdehUgjgOo20vobMTRZWqxuQIklcp0QN/HrbZzXGNhTw
0dXSXTlM557ToHxpkAWabKJacJCE8fxIqsydJo/JrswgTsXCX3OCm5HVySc9bnmx
X5imopQ5RvjCtczeFUt7y28ENq7ZMBTPOjZloR6jLIeIhnx/uJIHqhKWk/E+YF8W
ElHx+JvEITk/wD+F2tib6ayq7wjtWU1xYkJxYmXlVWugZSmMQ/iwj9iZqqWo13Jk
eJWTGV8UetQv0lvjsZpPcpwUmilwSqLYZ8DCWEiZdJk4LIg0qA9ItyyDci1WPHoz
QsHL54Lv17TaDdwpwk43760tN21IJCeXutlXIUiHKPDJib5Q7qnOaSxKcguw3gDR
ocmeW75z3rXCadQeedQNE+ZolJKJK3s3d/MXekxLGtb3Pm5E3yiWaf9ZlGEaarYz
K3lnYLRnnXpa6BlgCApXUv8sgzBWAhbKrDicnGlVZU0mByoAV88BnCYv3/saTuoJ
zLa0hhOESKEIIjnp/FdvYZbJVlHiZYtMdU6lUNYpxB2rncdhlcrVmUHNwhRXlfGb
stBPt9PSxtP6zeM3YZfnqVqRMyjwqfMxd0HphPwAT08QQN+BCy1SV29prkpxof3E
crHDLr647SsUkJr8QzornFOu9Erws/qVnjLHa46Gi1pkNTvsqLaLVFZVBXr4vIVO
xCU5wjC+YRF5+0PheJUciamalVcjWKJG3sftD6tPk3vT8s5wrXjzo78xkIjlsCnr
1DIgArXDMgyHdrbl4qsMeOFB9dUpxsLxtlfFuZGPdqvr7CuGF5Vl6OLLUR7EGCvj
FMqVgYRwDRtkAtDhN+QpT/C4XJIynJ+jQWXueoVDnuGxH7AOyTZmCsgmE5I+bLAm
1h8lulBLXALd5kHoC3wLC4wQ8TnoYSnHf4yd/jBLux+MV9vJcaRLK7Txu+qBVScz
KrVqjCh0Rzjv11TpMVE6xViy+xoJi/6glidaZZWyZwB4EVfQVHypGZw12nObXl7C
bCVq0cmnKD0rF72NJgrqIAWy0cjWeNezJ9m2G/PeIlohj5pCcmu7IKxbQ6tygyCF
vbQq+Yeb3xg96z51Pno7cSw12uMN1/gyWrNQoRKhI81LPH08H1l6FDf0hkjWLOBA
gSSyy8Fu10GYcqZ/gqyPmuusTLCDpBsaqWwj7oiJiTHocLEsoaQ9hCAYdnK63hSd
UMWOGgfQOn9BEEiLnD523lL1X+YT2Wi4eS6uM2as89wHLqGu3Tl70GwXVPgIaRD4
o5BAGWxAmlv0xWW3OntTArBmkw51Y645drF6lUvDgzucXFaepYFRUnFjt7r0ZcT6
ngSGSKvWhcdG3zK+6dLiu7uMGZEiUa9NSXqbjQuw+ICFeChh+nJWEk/rVPUtdqdn
ZQ/7NcBPkSB5JaF6gsO01ncgRa9h0sG5eZfY67jGrlZGqYDAvxlhZsnvilai9l0t
HPKWhIsIt+0uul/tWguVAqTWdhegGCpG4XOzjeN+MBhSGRPadIbnQkiy8bxua/QB
29A1F8vWErZVBrr065e7T3O3DOYmgvfyTS8QAvpysgf+26/x2rd+/ujJhZok34ZP
dQ2378oHyf564Iaa8KFFgSgZk1bZ8Fn54NLQePrhQKmu6v2CJfFqsOZQhFEygBhv
f6zAXsTLbwhUa/M84nmvHUxSQ/RG0GjpwyvzWr3+zyuTGfEdNo1vcFoLeGEFKkcX
weqUkIp3ID7MlCBZbTqoqqJ7yq2ggBfh+A7r+qV20IAakEQB7m0nHbGt8q649IsI
/LbLWDS9D3ku3Iuy1t7K5TuONfRJripboklNGsruRqosGdBS+776WuPpE77P8Y9b
ksGO1ZXDXzNE8LNV0Fys+eDEQDW4EPlVBk+roUzubaSfx4gbk00SVhuufOR23Uht
NF8aTq3KgA3mhfqLX2EITgU08TVdqg1o/Zy3C+8VSOm30QVvsqciIZjpz9+fpuDw
irlYkG7Q3hLbAdiV5/GSLo07JVLQZEtVI4EgxesGBLZ0uRO1siaQJ2STzDq2716R
TCCwvaoycG+ZI+DpnAu6daxvwRI691aTsrdSAnM95I9vZoFNja8YRAIfmx/8wxkN
hsepb9fxyj3x/Djdvz5KiqmzFda1ObciAhDVkTAfz0aSmyXADbwxVqysbk1zhVRg
MfS/+J3FKrVbjjIQBJkDmBifCyuagtdAnbQY2+6+QjTHD3s9GFbk9yxDmPg7/Zu2
UL5iWRlXLapYBY6g/toFUulMqiz1W8LyrZ+uXR4UC3nlp0zlKi0eM3BkvAua03GN
vK89pDAV/b7fv/ZIL/i/M8An7R2OEf9SObZUxhh2siXmCeT3WXaUw10vxSk9qaRH
khZvxgzuRQnGyCWrb2gis/tQ2dpqSKdWi9uXtb/05BjpfdHe+gd1xFHgrvoADKn5
rnnhBG8ayH7v2xfoGsqn3aUDQNn8LFrYPuJazIDbAEByKZ8Ke+drSfPiPHQiV1Jj
cP+7pg3TL0grZS1qHJMwIErxJkRfy8vcGISsfVLwd3o5tGfPp967IdmEXmasUxY4
D2Njvu1vJijSwOgtbGt29lHGP6FW0SYXudFyuEx7qeY12QtvGGZKEYPWQk9ZOZKz
O/aLGIl1iPw5nxXYbFhUYrb5nZt7Dc9gOsiJDoLUCuq0UYkbBBTGf/0iWH/KMnpR
uUPwmjaO0uOjxAtcl0E9FPC6l/BejOFHlnqzHEcY+550VoBzNueXrihGneb5CmaU
HeF5CqqvYVeyTcR2HgdgtSdFRIwHyKLR1RJ8+CV+s4NFUd6J0rBDg9sDMgBshWBt
MtGQX+k9ved9ZRNV9gImpyPVoWgXNQ0nmLWgpFE0NKLpjUX/OBwRkoLeyYY9B6DX
hAuaebasQFEIjxVfOtzVZl6lkmFeIHKCpKER/dSQjEL9PNeO7Z+AfDeUqE1N2ux1
Bqw7rdytSjCzunJOqwl+MxBv5/Ims0VYJ2//CzDYG0hk287Cyo68t3CKoTYrsVTN
v/58i7aJw+WZS1g4D+YOhNVxBjhtbIE73MaYf76baW/eC+Ay0mH6NgnamNakc8jf
8JVpXG+u7YbIUAKzFO2bGyKKf7GC4mHSPm9I4phSZ95cGezEnnyjuBrJikodH5Z3
wLJNEGnlEGk3yS+Z2OgYQQwqDRMSatmGSYNQVFQKDgRcNPpSNi0hwh/SXRSnyLDe
EBbdcAJCxYK8T9DNTbhEAeQMi2ft5b0gvu2URJF2NelqYjHZ/AN9lOe6bpQKMpq1
QY4qB3D1CgKXoVkkH1j90TNFrxfKoE3QJi6tIYwe5R5ueJOIAxlmxSYK8K7G+bxF
iSYyVDLT1eCz4QENxd/qIrtiGCSVuwXrvl2xjAy7wpeg6qwjTeqVkZ1C5WnRGufJ
2+FXPUR/jjowLBE67HOGw0V9TfUIeyEWgaS9QkfRpcm5ZgxRLIQ7micU0otnUYPq
a5US7eEha+WULFFNixHQHdhirMMmkJOygMMZl1U4UJ+vcUPjPIKIZfNMyo2xyLDQ
lIIdEgIkTgB2LqeRTE7hDjnPiGlTIKXqx8BfrDpHSQ7IVFo0zq8i/35euPWoIgs/
g9UinpI5mygsH/7SA0ksFAdgV2o6LWSOx6F/AxLDfzlvOgo2IdGwNTVhcs/R1BW7
HReQLrbTpoKs+zFoMQ3aEtClvUw4eDF2UkP2oZ+GTiPs5YOd/vQ6/iUHyZJhM+K4
kL67qQB4JN19NuhfrisURFwpYB3gqUC/qftWzsERz/i+9q6ZJ3UUcqZ4hkSetV3k
41GkQEBIGIu+IsuTTf7VoW5pHmB/IfrOYCdgDlXdY8IyWIsJCsF9ZCm+5IhZv13F
PDDl5yrxHrrmNbDOXDPRXlUM8befoe+EJI4i7JwMWfIgxrpnB64Q8+F817lXr1M7
GSLqEOAswc+AyHUdLHL50Ekh7df83rSC9UOmFkAPekl70EeyFFgptCfmzO6c+0LW
PtOG9s5sEMd6abZYa7Mgp6cDAhcjkDv8/WAkHSB4Wfgn746jxC5fe0Cubbvm8LDW
jpSC2jml9AuUax7i6otWAE+PwlJbI3I5KX5b6NRS+YkSt+Zq2rH7TEEL3nvibPre
U/M3BfXLEVwyIfqa8BdPa/ZIhYaL7DC2kYLtDdbujSjFOrFjEQDpPleeyKIHgU53
ErE/RLvmPSzaE/CNwbrZxq902Lb9vwVwNjfVxNJYPureHbVX829nyu1/b55jHrkK
vpFhn8Jrophg4qz37CT85U619xxy8TQ3cIkwLsrtqatPFohG5xJpjsZIpv+qOdhp
kJKS5icBtdujnCiw59DbT7eFCAkTf3KtPLjkMFkyE9lO6vvtuyzlLtQPt2n2dWrm
QgdRZZJeDfzj5GnO7FmDJgrPgb2giLtPwMDsL7O0udTWCYBc7cdLprXf1u7X86IM
OeUoLtlo5wPWA8UApyW/sPUxmtoR6VK+B9u7OkuVHJSHp2i2mdEYIg6O9t0jIBFM
l6mpiuAaL/DxGWKCZ9I4RI1VU3+ntckpCMfkk5L86RQPRFsxIYLsxBwxa7XHP3pI
arC9X6u7uuuh5xcelTa1uqKSemr+Mk0RkuZFAEvlpNvPZzIeIRxv+Bfy5/S2OMij
xiwKatAJvYER+DBNc8/+I8cqfP0jmCDwn7Qd5+SzZNVXYGD88lJdy03mvGiIndlK
nZYpX26SBQWajFRQRTPUGFZKPDGMWwjphhskGqBsQh6iVAvCmwbYLQwkuReMQgMk
xoBOf2OhZB3AZhEJ3Ahy4uTb8ejmoQBiYTWw4pmXv6onf4gJElSn9yojW8pqpiNt
DBqJ4nqTyO4XPLgzZwAlrAAfDVV/SG0nasKNVO3eILYii+2Ip2Kgwp5to0xAyo9S
5O6wGU8tS3M21zoB8NplWudLe7W9en3ZzbvSanxEuOIr9YuhbNpdQPVvlIftR4Dm
/7TEnGNWKHG+skBwilx4zaTQBMFSdXR7MEEeVSllEE0jfeo0km4Qf2HLdhLHvIiH
ey0D2rfC4aXrUFgYHTpMILxoQjtR5x0SOuF5z+Kf+EmBcCfnGSzpJsCzSqMVyWWh
tQr2aJlqDprBnBfMYnYzjtuiHJE2xGoMCYDR5P27WxNg1Vwyz2v4uebMGiO0ySOl
b8nTkBfDDHuGBtQ1YairSFdIzTrTKLAN8pLc1aZKap+5ix3+7nqfoYdsk4eWRRh+
mcqwBoooqkFpATSG3rw0njMOXGdwxI+10DxDhl8s/b9E9aQB0d07YBO8Wn/bTiiS
jKi0ALcMk5o3rnMArtjWXCe49pHc8ciLumLCQb0zdXGOU3OY0lCmQMAeyKt48cXZ
7DD8/qkJKKZkHCDCNnqK7J6osV4fYM4cXJUh5Nokd8iFb7WVqRhUig3EVvaTlEm9
mcz1MBqv0XLfYq57Dm4mmucAEbtuatRo2jCT8wR0/VfhgLtn4kXLcoDfopDYRpHk
wXhtO7uT2uvuQ3KPuAZM4HuGmra1FMGwmsiacSojmCPzbA1VKBYt2WgW01114c5b
j3zs/nn+GmnUt5xnSGGdnz5vZOpjREdpx44fs3XwFhYLJxVspM20Yd7YCIX+rw2+
x9C1xGQ+oSeq7FGOG4v1dZt3+2WGaJ+GB+F8t/q+u+gd96Od8T8XboXS77Cmndqr
cSDsgw7yjjgYxBACL/CdN74hzkMmk1WdMZ3zyhgIIWRtBQpVDmPBgBF6nbqKpdQs
jkYeLbYdfCpJq1FgBGjvZaqZAvqpY1V0Y79DgrIZQq5KwW40jxodJk0emnWq0PoN
Mkq9nCDI+OJZ3+AVSyn0CwcuOO6o8+LfBgtJ6ZPD5YAnlXnhCNMv72vnKMy2D48c
ujqRdDMrCyULAa2+NEZLIm/Z3ZSIHV2ysyHv0Ac/yQZipR2eRQmYAfD8LXlXiET/
PHLJO8ffIlWEhm7ouyKkXYvi0zcP388Oi8LhLnYmoJdwi94KQNHuHJ0FCsY/fFZ3
p3ietCSPKfVyJoW2QN6ZRnJ5khwyjpDz1THPni0YQf/b8zF0/jD9VD8PjfhBZ/zh
GHpDlmfebsdpzbVAXY+PkC8e+bBJkuAi5EArVFhnWVV6PQI7sUFXwWYIdsgAxAv8
ZD60heCaHAhrtoZ/mtE3HQByhYx18fgPRcb9UGWXBTxirmEvi14T2lozjF/DdvMv
tKBjwOswlYtDLZ8LMjhGvLr2FEtxGZeJvH9yKobjtarCbGIZmjN9QS/Kp2R0yW6/
TUFWooEB362mKfiKtpub0ptOUFxThj7a0Y3xGfaf+/AZVe3NsNOoqP+ZVfNmbhWI
r/sMZ1KpM4htd3rwilAaRksa9EIZRpsXXAeeMXVWnE3gM31VrXcgFErlNYZEhwIM
tPOAvuakUy2KjFDK7iq4xDnbZqLCSfzAPu7TtWLLNN9EsIl0SdjxiKzCW2L6rMAy
bLgu0dDae+dJsBWcHaICTWn/R7VFbrT6oWFTv6OxOOiyA49QGl10zUZSVgSa6cNV
D0hEHrtkfPLu1cV5J48apy+uH5VL0BU2FPeZIVuMn58kdRnC4lZzVCMwj6z6DRSX
/l/1CCxNSG0iL1LgvALPpR1XtBfpJ2SDapuuAL12uSfxzriYZqwts3wGpbC5GTIy
sKfOmeC5jpDJQgON91xMswASP00WAOGq+j1pPAEEPset5hSJcepI8araWU8jTrME
HAEGZFhdB8jy4dzkRVKHHudTZxTZrO6VIm0ny8tAGaCg015z3BJy16UKE4ph+gvg
q9x3ayQSesYwXHfxVZbmSnmTn1MU32ZWbsnvfCxLEcwQaE6lfTH8JrGVAcsVwdDH
VxOU3+sHI006AXOkDGlmH11LSA+AIP6XbjmP9hHsbR6yVJhtVAz5UT9PPuiZDX/e
3EA5nktR0hw28fBw1XmSIRegPtS56wJyssKHKmiiuonMC9ApZQQhQdH4gEj3c6wt
t0QNuHPLnHoblz47SGGoldswKf2q3uDSlHw1NANharHv8QF+FJKTsC4Jt12lVPx1
VGHcy0Hc4uMyo2Kb7a/sJ0gH1q5TwC/DRkPx0+jiomCWmhWPOLBeCzqbvqo0rMdG
x///7+eesqhJwVAb6hOo8VpEq47g5ZJZZuCt768hyWmybQNh2LrScejV5KVvp2pa
BaDDxZ0JDZnHSCfTCvcYv1/3p8imMxZf1wjgXbhLbfE99XswGHYRR4pqjmAhzto4
p2MseHK7IrcF2Rf6IzuYeVDUcyH2uFuFfvnRU/fma1N1eIUiC15zW8QKdY+5sT7p
xbAcFM4nr9s6JRDkA6rlUOqlsfusu05NJoHyurmanWTuBAQsH3roytarNY00m5Rr
fIJPhG/3/KKA+4IrXVjqg/iHwePeXzTw5WL8WhX4OW+2+pCY713ZHby9baFTZSLM
+5oync3LMePPG8kd+CQ/IQ9Sst6uHrXQwu6+xMcgZTj2h3LA2kHzWQ0Hfz+8tRFL
E+rNJ8vAKEmSjcmC+wRkiwPkzOhHtQy9M2iKTw7+OPp/BuBmaASjp/i1GPijQZS/
4bs/0s+64W1wAmverhTgTi4M5XsaTFHWdQ1ubd6y+MSg08n0UDB/J8Y0f6KxIOfq
VOUzQwU9JdXrprRyi40LeStPdCXY+h+9vbD7PEoB2GpYJeLvNwOObb6lURUdGJ/h
jKUFrf6y9hzRA6WCwimU/x8LYZV857LDbRyUb68soI2gPMiaQOBizA3RolBVL02N
pZ85MrqImeiXTBw0jM7TMMjdF3ED8yys3qvfABanxz3JxZ3e1G0w5s92DjIygt76
LuVBN0LaAnEeTiaz0Kt37VlSerB1MtBttCfwrFWLSdCxNdawetR0/azgrhYjNoN7
pEtbCxj6yprzleCMq8QScJ3MTEZJkEqVyYSCt2CgJK5whsiHpF8s2kHyOSYPu/2Z
uCtzcTFrwEQ/i2zYPJlsHHXUyJ18KwD4N9optHk/ODTd3+PCfCKeAjobjEM8SLRl
C1vcDHnBbU0eq1K0iwJOWOF2dA3hYtAmUKUj2S9/0UkDhJvGAqQwzdRIMovnn1K2
tHHikLP4vU2lbf+gq7uRqCpDEBVnR1ImSD8BuhDinY59FSsuchE6rgN1fKwPDd3P
Mkqq3DIqhkqL93Vqq0CTWILRN+Vzn5PB9ux5Lzzgkpr7ba4gBQ3OJo7rMDUGe46h
XOHzEpB+rvObddE2N6jhwFYvfUg/6fN/xHx+sIJC4fBDErxa1LaGNO8zLi/YjRIo
2qW0QGccaTqdtLwDCOLGEYVh70jhdFeaKqVDbwVRpH4i28+FDWHwBLSlpn+xpkaG
4GhPKkdvFvW+Vs8FTOWf98o1uNb6m+qXXGOTJb/HQtmFJrDX8loe/84wGk3AkaZJ
5W6wxAQewIzN++ZD5Li8d3SBFdermyZfC7We0dV+xYllc3xVy8j4zv4IHW8+w9Uy
ryTCbxXrX9kwxEo8fHdS3B3yjX1FVvX61ugTNsEth9W77MfaE2b0wd7BX8VQkajn
U9W4RASftk/5LNsjFc7u9YJ3faBzAQnqfS03wQv1nECgXEXqf8EfA83AcQnWKw2x
zfCt5FaldO+SRB4U91b+TTis9iSHl3pkfoqshGXUB12bUgWSoApwId4Uxhfgqxk/
oZzFSD1/HXjwvg4Iii2i2ai6VaHk41WEiMNTtqQQhX/Cuz6ob9tquBn52XhQtsVO
VA5Wz4w1qv9G0/rUThAk9rH1wYRpG+umDF58Lcc89xT82bkYkGobyaab54FOvLVu
ePuf8X6RmDDbbN6leDPeqrrkv2RqhHVeJ8ISBCQUD6uvB2VDsWyH6+9I0DbbWTRk
VB/1Fmyqxq8TZMbeFbB07FSy7CshCcBQlTbIHFK6FrjaQY9cCaugiLwKN5mqc2LO
0SayFjEMgHPN6VXi6HIRn99YvpWyzMQo/uyBakCot3MowG9wSUiblmjLlGpok18q
x5h8pPrx5sRB16D9gL4zjPTRt8BJ03n0wZWWFbivqDtdizG4UKWUop6Ln3T53KQw
QiF3OxDJCA28JfBZsfHDv1AwLIBU0lRfnMEOIaRoBB7hBPON/tj4KkZMci7lvJPk
4CBFeoZRF6odC3rGi57O352XmaM5CKulG44JPdTKJzB6/FujbRYmxDXENXHGDIgw
RnY5DLb835POQBF56A2hVIsVNoTl5dCmhmjEGldjZY1SDI1glpR++WpUJhh0Mh9D
GOKs6P2T8Sf0FAgBgfHtZq4VO5iFF6/xp4ZUe/wdrm3H2JjwC1+Sbo8ygmuFMjZ9
TFPE6bbijqX92NLlKrWmZhprlf9KYZ1UQd2tWDC9issH8ZnytQmqn7meVFrZ0ifx
gGVE8dvAYqmVVYriF9IXF2F7Jbnjw42gDZkeU4sN9bl1SBWfvUXu6EZapBSPEAt4
t5A64ZVdVyj3tKEzI6g9oH03nNmf6jrKnARKacpWXpUCytOPBfI2SSVsqOSdnENq
8SP59r6fmM23iHx6lr8okplnICE4FqLhaT0CxDO4ysYMazCEgPpYKKRtLdwxYNTD
D3lgK5XzHBI/EzOUKhm9//QJIVbksOcVYM38Al+2WIkreFObJ0XL6rWBLbOtjO1l
rDUjX/NEBJsilOOPORoMOKmrLIfnt9N+1VFuu0vCfZCXwSazttfOwv6bpYpAGIr+
BMiis2SFR9+6ibp7wZQSr6SUra1KQSVr+MPFzztteDDY6muLIKmkSYiEdX+9o0lA
D2NWypol5WP5G3QyAKsdAhJ20tBjn9IZTojQrshKmbSpNjH/vne0FUA3XG/zfE2Q
sACRt2q3fF9AV/036YmKNgWpWGHBhrz8q/iIbFLWiZUUEg4/iHMBmLcuREwgtUq7
H5nRNtmXGDfzEw2sIzjMGyirMpk5GxVuEamgBfMwvWS0XnCC+/xbCb8r7GDGZxZ6
ozH5/PzvingddIr1iJXZ3Huw+MGjInFowl90cyM2sE6qvVRNwSQUmlii2WAW3zCI
HZsyIN+8gd/54q1Blut8BJzYJQDupAqlYcHY9rq6mUdJIZmL/+l0gfjY9ttwKPlX
0WP6u1A0yzM/NcERXTJ1CHK0BgQ3T3XDri0PJ0yJq6QbuGkf7VI7AF6yNZTt45m3
6j+b1M2XtRiacnTf7NnRfBiGWNyWJiHI6z51+EhvP0YemKgruQBAyZCz89ERBoDi
1yTSJncz1Ee2FyCmKrzNOFxvBQIXT7vUjj3HYySYajiuQ4wMyghWJvJz6t0BsQs+
Tt9C0w2Y2MN/zsOl5J7WIfwi1mM7i3XHRp0nmBfBnyj1SHp1xIaZzIvb7v5FDqgK
VkNAVNA3u3GTY64C1XlFhDoiX8p6UMSou7gELDr9vTfgXryGfcqmFFTPugPAobCf
hPTpaKBQxTxJrSZc2qb3bAWI7Oan3CH0akh/xj38/g/Mhi12GTI/YZYyPFAabVbv
IuKQutUap2rEtmUzGWmCJ8Gy2/WNpiwqv0cDXBzDpxTtQXCckGJz1vuNZdRYoYJt
0wvVm4Gj+6TCgTDrLH0v+PssC5paEL9gORAV3Tilz1BUPfn/BQ/mDhb8SQiLnHGE
SObVFrtZnw9y5JD7G1Pk7cy7khQEwoSfRlxYkCIfIHN99oVjoXWbrysshaZUVGjL
dn6rZrwTPnJWVkT/cSBPoB1pJA66UMYK7hyaoXM0x36YQzlpS0/JiPHid6pmuzem
U14HSGJ6Y4F79K5sTCn2pul4jLeFpQrBMjV51MUyqU+g5l8wmrTbhSn7ZnzBHJOS
lP/43w24BydAK+DtKQa8qTNRYzEa92FlAMs8XyXRryObmrjXkMbD5GdOwl1LTGMm
EILKgYLkKjY3mXXzAflZ3kgb7kgAa5hzjciAstVTn6ne9OwKSxqKMllVYS61lYnI
r+VYvPW5TFHAB2oxHbR1cP16G5VABTBAIICkYLPYpIL5WfFBi6NRUFSwmk1kDbXy
889pE3Q4XO4AlgY/5jJsElWBKAsjeJHZIPYW2VXOUwH0v8MJqhjFYZ7ptICNOAcH
X1y8sxfRu8twWi9J49qFG9f8aZPDQ3MUOwH55LRsD/gVAr0glbTOXFDfM00QP1Ws
F/Y52s7JQ2gG/xW46TRAiNOFR6iEjW6+SgoBsjHNcItcFTgwj7Yru8imFBym6fa8
z1/GlFVLIpvPwKt/dMNw5nGl+22mftiIUE86Eoor5O1aysuA00xI43iyXjhlqnqC
sGDXXg4pm/7eD2259Y+2BQh9NoQwzn1gLBZUAXcQu2oIYSxwV0CeZ+GPeV1CcUrF
qYetiRz4KTK/AscAoyYURtvfEz7zXfEjLf6m1PXGdeZW0FeD3z8GES1uFPg/QA4h
dKJPaY5fWzTt8JGEBwMG8+qWBHVR+7i03CElLqPnLzo0un9AtnUpTrQrJCMD8oU3
/sTXyYE1Noa0raNhy1FRt1vJNNjWx/vKeG8T8cxehqgr4jaoIQ/LK9M+0iOo+MDK
QnCoTdZsewJ9ja/4bc/FurmtvR+EcU4ct3OMkcbpozMNamun549ToPebXhu+R58E
MO+cmXdRVuMIXnKq+ocwJIwtScrJ8b5tJ+iCcFvPGN9vvUu4aBHzbhbJD1uMmCK4
Fh7MxJMLP6o2oY+g5+GzRaXoB9OOCmhakHPL8rx9WHbSUIKkjRcAoGcFmvu3o4iP
aqef+Ph2nm7tRhScONiSId6cT2Ie674N/hbPoEn7HKnvCFw+nqK52kuNyWCk+CN3
FVC78CS8mwy5aKm//452/xPsl8zbNcdbml3ThjjrLmWPz/JeoU0JpB1sS+h+mKnF
SO4uuC5p/TpYziN/490+c2XPjnVVyQ4goebOQnaV3jYhw0XqvAEMhE04h61e3QJf
W9Tf2CcKUO8uP204pVFn9SvUTOfAlOyPCaqJtoLdwIIskWGZfhw0fwU8nsM2pfq0
P+1FgXvvz+1WAH6qs4ITX/F4jSq8Hgr3+DhoKfLOfMZPiUnjCfpPg4fcjkEXHsBO
IqbdiylpbC/rtdVF/XpTI0ZGMOKif6xjUKu/g1rtZlw6qFX8xdUsWgfEhtXQ98dL
Uy0WobjZ8YiyxzGrH4gDkUblR2nlndJq0Cine4dW0GaF7Kn5u6/rS9gI00JffuBY
o+60YaMbQ3ELPc2Tn+ho2JZ7494fac5+6MYr4z6T+ZowhuFB1cnIHFNjBxSOPITr
4xqeg9wbOL7krlW5BLlcuNremoN/oQnmzaJ2/mZIasSzFAE97tzhT+5HS+OzvoMV
qSkz+ZnsThzb1wK/cR8DGoMIC0QXY+aX56eWOhddHSriK8OIBbFjpJ/PYxscOhs6
ZCVrPYiNtYNGt9rFML9aHKKbJA9xmgr5ALRcVW4ndPmfUR7J+eygzwQX1ZVipVtg
2hyJ+X+P6SLLbCKImjh9rXwf2LO+5F3V6Ike1JanPg3mzj/jiBmCBspjotqJaZWd
AucHGAkG5sNSyeYo33Yx2oARPeLDtiNym7WKEXgjnr557CUHS/ynnLayuQ+kXQsi
8UsAwjJymevAK+P20Jp+uq1vuUnECwgl+FLxF2JDHgXLJAkQNLb3LLkaKfpQ3Ynt
XHxmPZyW77Jl3DhPfnyL5o8fHJuq4myziOVtrchyx0G5Sv/x2iFE9w1pUipFfTL0
AFAROaYGLGjLwI8IRQBZeEv4JqqcEHho8vP+xL9SeHu9cf9cBbgwCSyIt0u9bskL
4jb+h0d0kAEVmGR6M20gySbe6BK+9HmQfEfIVXT6piGpaipQVh4B9+9pLe8HYT9V
dM0sFZSSbzffOwHjeB/yLSxTocCP06JGtzu3aXjMtLo9pX78CEZQ7+kbtWy8v86n
vvWxY5sdA5MgTD0iqvH8WJ30t+e4sy9wJT3ulafwiDmZPoq0athQDrncD9v0C3tw
bNvfQFgFCl9A6p17adE+vz7yyrgg4tav0Pp6j6xPiRUx9f84q/4yuh7+V470anQh
v7irLpF7je0ZD0C1etF79s6NZPq8b182o40eb4kGk1h2ZDLUXp8TOx5tUTwKPTYC
q1nQZT4i1NLGDAbzk6fRVpGoMxc37DVyBuvEkgy+LDuspKdq9xPZKrlE4kvNEz77
X5EWOFI3Do15D/fYvgIuKzZV2QkKL9jkk+8If+ez9IxdXMqlPgbP0wZeLTMwjV9/
z5D2lXIPYhBirJvyOAUrFCkqglPxqzW+L5FNz8K5wSvWrkScSPtfa0YH1PDB4hJU
dI1YDk1adCd1fsJEWE4ax0lASENSG4DBhcaVK8wKUecMiuXDXgn/vGSZOWzLBxmA
Yx2w10v32oz/IH14xpvym6ZQw5XYyiaqGrwlVc5xKEVgULSHC6Bs3wOUmEfNcZf+
ae0J8qsrR/a995dXegn+cew735ZllaVJ1dYWjJEFz8SgskI7EMoPy3JDzpl2ZI3G
tjCLMN4iEt6nwKMmQWPhejOfQR98iyTpKaBjps5dHglDpkqwIrp9nASdBnNsbMc1
wOhP/CaHL0KtTyJPfaDYVpvPdTgbDfa9xJGcFmMz3HbvFrnmj2+FvhmW/m9ji8Fq
Ng4asMT5MuCyMxT45HOAaDgQdCBpbXCycaQbR6erwkNsHDN7mctBMs2rXrVoGRHD
FWZOnv78ePWWrI+MDsevkkaBv4ZpcgBZ+r9xJn7XqgjZ1n6f6UvRW6GKWTTQoFjD
FgeWhQCZ9f6+uOyNPEc9lwfOobX3B2eoDJxaDbCf5xMM8jiedaN8k/XEoxVHY5iV
rz97O42heGCEOKN9gbatNbzl+UM6w25n71V7KCFVqg+RzNCZAnGUQJ7ftFxyKvHj
vqGSyV6q6dpXr72amxfclilCnq3Szn5YHttahC/MH9x8YV8MHRX40PvIujA+Fa/z
zkmXf22KqV+h+yLkmP3SSqngyCVB8QU6f2sNa5vkvjr+Qe0F59iRqcm6vCryngFr
zC4XjZkJFC2MCCUgfLIRCbDdxTiZmu4+As+oVfsVZe7NeiZFzGmcsvIumSJ2tdV+
rJ3FZlWRpBwY1mCp+runn9iAzptlBb1IrgsZhwTkpEx/sJ3dXkwbBXQVgqBLVqtn
8fHQ/TTpTl9d5DkqME7xZDXoeZE/7XkPiXkk49xbi0fS79CMLvtWR51AHz216Os1
789FUGJow7qXDadn3PejRbdpO1sdDxPrgqvQOKhPLvoH3ybDTKJQTjUozL+E9uQf
3Y2adFYq9HrXi+uJ9WieADyWXf7OpKdiSg9+/W9aKvVnjAqZH0oIQ6ISNWziBEJn
NBH4LAHVl5H+ypnSAhEWxTUUAMsZGQMUbfzxD4QMUR/C+p7CyaZfXW3Rh+VDHKn5
CbLQd6TtHLUP6r5ww3SoF7jlO34yBlv95qugSIBG1E3DWoTgftzWfSI/j7psGj6S
E6qAaMfQENdbUwS2YEbtT4Q0QAivQFNL92vdv6csrDZ/PishRi2QtKtEIlFCZVhF
ZXYFQiVR6KwkN4kgAVotrTAEc9ATbLZgIzs+TEfNPQSYiQL3rXK4Vj3LgX913yhv
YTAX0mkLwW+v+Ezk9vI25arElYPntKcWKu3gCHtolu9aFCI306CuyPwfd/VUBFsF
t0S1ZanZAzY8FMH1aCGgiGMZ6JayvxZB8jRi8um1uAc6h2s//R3GMCQC3Cp2cDwt
P70JGoHSA/EvkF84fI5sPj+fMGFGoLr/ApE5GUU4wTeTZ8LcwfjRwHRvUuwdXpLl
8HVb1SsB8sBa7rkUDpzPLaLmtRNigCaarYLBLbR8bujGd+kIDd7KJcswWllE0NZB
dzfOOgTqGt+HxHruuDTQg0Bo/RIZNWRuNJhcz3nmkJjDEEVvb7iRQvh+KVp6bl5F
O2D/CysQcagtRPnyCKU6llo0IzCH9bBL6dZGrYIfy2803qv/2frs/OSCyV6bdqGF
1LT7K9051d93rjYg2pKXGCzWHhOT6Zilt/AEtYkmi5pfLItJpqfX79jGZAVX733+
Mbb4IyxIQjQD1bXYLGgYe3SZQkSrUtLfwcBZ9loaG1Spd/BF+PAT7QC7GWGKZt0e
4zHz9iOxS5sUjgFri865ImWHeeFZS8c5WoLIFqRkSRbTl7N1G6Dt+0BSokaPr1Jv
zt4bgLuLW+n98K40cq+gg+tE4Fs7/VbTssg4EMzA/Dc6L4NrxL7TwdsAbDD8GFPi
hKsaHZeAYHsCU2LeGhB0QUIxQE47YLD4dxy/t7T9gZNyTlZ4xKpquMcWNvnJYUw0
BZAKfS6RuYF8LE86XfR4YRVteKAOqIxe6iH2tZKaTpyMBVT1OzMhuqGOy1fyIjH9
D5u5W6QrnuMI/81LNIVninDBOM1X0rVjrS9L+li7y5vBVzhk/IikM2XBRwy8ZufU
EgsYTmLAKiXPsG7ibrn618kSQHSkRA5bUlo133rati13j2IFiGuanE15DfK65RsI
bVUpxY2xu7TP+T5GLaUSxSj/dc/0qPTnb9WXQsgR2E6J78USkxeyMIm8TUqR+AzV
GFOSRTxnSE0oKqqg/ITdhufRQCESVo0vogxKL/Y46Kdfmhb1QtsyrBH1DY14+jp1
bvhoLaMacheetSZt7gb0zmNQbLHo93vNw9ljbEnGp6LUpgMhZ8X3lgHqM8IZUSzK
m8KlfgrFXHGxhtBdauI6GBDNDRTwbHNAZlNAXyUrdx07JEu9n4THx72iWJA9u3ef
tS93o++D6zUEl2Svt1q9ibkwDZlcDszTa7pnf9EYMCIGESU16vrIBPR0Rio+YWsV
9qug5WSHsdljWLWb71EaJfbT3Biy2gcASwg1MYTvCmBJ3wltOlfmG3OKpc1xedHV
S2cxNdrPxkP549vIuLD8VYlVLM5TS0PhyEZxl0vzCuKrIM5I+3d/oJkn8x0i1Q6V
n2FaVAJzsOptpgwBKs65Vj8EXYL3ulYds7L+SsDsSA9XgGTctlnJbmILrZgjvBL/
zj0Dqn/xpQAKhGIoCK5jOGhXFX9Ja94deL7YUedG0XK6ViuyHteR27luS1mPykxv
Mn2u5jvSXtIjNHmwSfRKqpZVZoSxo0CK0AtryPYN0vKjlhygO5KrLW4QDTHmflLV
Ko3h7Ruk/+9NE2NTuh+jAml4G4yU/kM3scGmMLZT+nrLp8l1oT08BC6xn3d7eAxg
WQ5FDTZP7pelujI6D0NBtGikQ0YUnXkxT1eG6s60XfouEUjHdfOFkZ75jtzAamuq
x/gEaXJAedctPwr+vMVtHi/6Cln4qnQExvEEaVGqfVGBnSWwJZw9T4QOTkUTResW
8OklJ5M2wF6/6DS4zEUlYlbMzSVUs/1Wug/opIlwKBU9hTpVZ4QnNZuesdjhdjix
5Umq3got8I2K/wQGQY1vHWooz9vT01dVnYB0DYUQAC0f8A8uCW0PyLT4U/hBuQfz
EHB/77LqRilqZP3uFDJRVcV94fBCrZKGPqZwaJ+xhXgn1qA/3Y2KmbkjO50YMHb2
Er0SX8oPD1gL39TzYLAdbIAfapfBklOr3l8TLRRX8pVWKd9IfH4KUjMmi8eIzJSz
pWNwtNDpdMmX5rc4m9vSsQ9upIiXKkiugXj41+BW5iYOXgGRVv78atIyF/lIcvc6
AnchoVymKjKkiEPpohbXf5WPaOgTYJ/g3FRnNZovJIpHGSd1wQCEycdI85ku2TEg
ROpLeyMiY9lCYR4mnFpDoMyBkFzrlmgXaWlR8n+7EAR4/hiVOVPzvCVvYhAq4/iu
qxdcESjarw/IYNlYE5Omhjqe92MbuujAppX+qlmVqT1bVT9/fCK62/xhDrUhELWJ
w3FstUlPoZKh6nz9dQbEBdophZywsc+GkiLKfBWZcxOom+Z2r/oLOvSVnaHh+mpv
h8/ysQ3u2szLh0T+f9UmWey1Wl88LpHNICazlHvJ3jzNIdK9oeu5i2obbSebNBsM
d0gipVm3jaeB+m9r4WZ3VEePz4foi+MKq3eE4BD0/Kt+ILodnoHTveryaSdrwVXd
1IYaElLrDdZ0f+OlqCj2i5yy9cxz+miNN7NhaETBu9DlW+9w/XVSwC5UHMcBzqkm
9VXHiEtWZk5/Fv/WpNubWBMJtkNVxdlAgkGHtTV+xwLlDITJQBVeZIg2pk1LioRu
hesqUXEg0RkwU5BfXUNiWPOh4aD/8ItRNRqZUainsEZoBbGegQo1vckZFi7nB1uV
bDvcV9WLX4EGPkA0w/d50TuE99VGHNa4DQU9TX0nnH0UGad992GIH02ZM5tYPSkB
v7I0uFYtcewWQAB8Z551O/oTq/JCJVnY9VxJpByo+DpqPCVKNo3Q0KZtEis4Fhxp
JQHz7Jrd0BqU3qRZ1aykSiY6lD7MWBkOsTWmjli8yOYesX8YxEhuLa2nJK9Udyxv
keGCAaAzKfmEr1WpoUqGgBTGIXXoY/wLmXduV4+3dPp68Yr21Cu6f3srz0zQDmq5
SW56Jd4LwHdpOM2P7txsUZ4l7iEeXzCiMSEEC5Iv46HsvRAgvpD39JwonphuP/Q4
sPiZ3XZ+I+YHAmfaqGEAeL3HzeFG6Q5/nHtj58uOj1jWF3uHlFb/xi4ux7Yr1Zas
B/cjOCTUUUdKYC39YXRBYR+XED1y6CgKXoQN7oHu6a+XemAsHwBtbC8BAkC2EPpN
17m1110tIVUwlxQ3Bl0P90nm0nifvip9HXYxpkl0kAt7I45AdZssJtSBwnF0ue4E
h2Jzfw/+WxDcQ8WYRAM1RO+naC8S0iBHqP8Wm5gFIK4FgyOsxLPpZsZZ+ZUvfsex
pYygBOZBdhkpzLxRORV0yPy35y8lQ2saBO/XbqLARcu9QG4qt+TzXWpvnxoq83g/
f/F6e0EoEYnZDx7GfV+Pnp58boQ/fg3Z2RaljzXWp7FyuP+kCHQAfJy7hO4zpY6b
8o3mL1uf7ZYfuTstkKTp4WlMTGVqItPsNboKWBifL+rnnZRwtYkVVMYgKkxzLdse
Tb6k3U4Q2sjlYmt0udhCz1gJQXvHG4baBXAFrz2tK9DCpoz5ShleY8HYcoPIEbOE
AGF/x5AIPyiWG10ffqGR+2B/9zr/JxoGAjNzyI4h7yl/Wc8J43SKu09SrEkbK/8e
YqlN8wqhp2UDyOeSVUK8IkSL2fzyD/94u/RgP69C9dgXd2EzuJQQsEEaa2I6Nfnz
/X82uCda+6+lJ2tVbMd7g932gHyTy3paV+H89+t+Iwa13XKd+WFtaKpuOJCSpjfc
s5xk0QSnoPwaDgUDNQrzBn20kc0mRdLqWlYci0BkJZWScviHjIF7D+dg+0ZhQf4Z
77L/Fb+39DuiYjTxtL0lGtl3vS94xyiO+aSE9QaskEYpOnVQ40SOSFU+rBnZrpje
dnnID32jp/aT5lKbFIrKhgfUKJCIigg8wlNu+VpOZrP4ptlhrSn15QyCQI4DvMv9
YtTe8q+rnFK97d6hg4qZcr64X+R+Fb2cmSdaXuc2YUxl+mDuvKBXCl1SPnWpLtCA
R5lZZJz8EXZHsZCY3QAPhwdc/9y4VPpG0JM170RQzo18gOH18vr1Mi+oiA2OfpJP
mj7EVXnnF0H+5aqkle1eNhf0MIhkFaWw2SyxaMmu9iEwkggLKxYu6gEGjROTrT9R
Gjc0xe7kF8QYhaMa+a9fbCVbwKvbM3Glcz53RYVCWYrqCY4FhdDdYdDxbhGDd331
I9TF91Uj9MPu6FccavfIYMyXlvNw57s+/+8G5hWV+1UbXdfx/TjzQv5RQ6A9iXX4
b5T11ltgr2mkUjsaOpaoju0CfR73BTKFByeQj2ljybsjBIpmcH80Ak7UIZSOsL1K
/NZt/h/GN+fs6SWnU2V4uZAbM92cCPTrOrUPEZYNlqf0zRZ9jzHl8t0GZvsVwFW2
qon4yqOxIxw0a4kqaFtZbyL5I/6WsZuOKzE+XiCtKGWWbz0y0Ml6NQsj03Vc6jRi
MZawm0bkUpFFLq/ghvjTyh5xDS1ZEqVjASKnAWBxAwhR3SwRdN5oASW+bq1pKgOt
uQ/XmtFS79qBboZixdRdj6oZJI00N/2bn6t3YRtMHGgcjV9vcHI86tRfIYmlfV0x
ICNxu0bOvuWBmr9E8gbrecenHnLhroNDiF8yIQhpe3NXTP3N4x6mGAxjDz5cqSJ0
hQARRETsI4JBIy/KL3bkxpa0GmcEAePT1zoHZnrAvZtYqGsoRRdNqCiAFer73THw
rZDvMHgjU+etkSRLQTeY5yU+eiulOLjXIKPBK9iAoVM6rP5iPuXUhDpCxYa4nSi7
CEtdfyUV+ka4qpmoGd83sDXGUXfatH10IJKgdzIHaGZBZqVJv1lX56xMCOX171nx
hqW4zj6WUT1jJIQ/P9ViBDYbputqsVb2iE3kFqA2lBMxv8IHTTgMOTHfkzEcBtyA
QFoZk+PNqn4FjFcmHjMJjpj84E9fBz7Sj64RZsmH616WJBOY9NAh1L+RSbSW7K0T
cmJ4dcWBe0a+GzwSK2dH8t6LOgqFnkxovHCOuijtUvpD558ClYdLRIallk37Twa3
1FVtrHNpJgeUS+WDGe90TBiUnumpxv1mADtyxugZr2GaxBjl8f2T6tGdrF8GQJJ7
M9mmosXez2XHuIoFM7F+wuMB2r/2qhEfHXZAcliAYF+rsVFbRNIsHXanEup68zsn
9lN6WJiH1w4bwQL4KvwBzJo4HWX0bmXScoDpZrbgf+hsX3Cs2KjOIiqnSzccwOty
BySoC2AXsPasA+QjijeqX5Ievp5ZKYErytBoyHgnpb3mhcNogc/mE4JyzGaLlM5u
Q7h6Jk8poQegumUdSKyI1v7zIq4j6ddFS2VYeTspGlHz1Y9DNWQViOfCsOOEapXA
tXs2lEU4TKOTHinXh0C4C5YJcSMMo09EB3FULSc/1R61R7p+6JPjsvcIkZrgdac2
5XPaLd5L0cnMtjNY0ubVwXKmo2BX77Fz5z6wxSBJoUTY2Y8IcKOUh5PdnGgGiJ4C
ZWxFrMHu7S9VHYQqIgNTJTtNfrYTOCLnWGgSoJYNaZ+yUutNTYPKWeCxtTg+ii5U
ZSKTQveDeGvH2YdKUwVXc+H3RG0YRk8acmeura4pe1m8W8hgidzSV39oSYlsi6XV
Y7N1axpJ95ioI/etp0OpnMH2QdC//ino4Nbib814YG/t115IlTGD3nwzxcCWnGn0
iBLBApJc3/AVALdTvQzlpfwJX0tULT3lE0Cz0/tKOzq2xTfpB9WRO8c+Q2EtKMKF
mTqAcs9Wp9SrCQ5kMKTmCo0+VnH8jBf5vfDcJdc4Fy09kMR3riOjEfH/X31tVuCl
HsaP87//Y8rfW2U/7Hws1Tm02zWiFmW5AZ5wFWbxJVpILStfCKQbDRBVVyb5hDhE
cYzH2V0CwhUzVNJEFeQqa2l3cPi+SnS1NE6jjwH9DGNFQm+4ZICAKM+U6ZjL1N5g
LK4ecilMfxLPCCnJdTjF5Dngf1YFPLCpPYHTN3yDPCHYdHa4yA0PbGqVVeYJJsCo
Om2zimSBpBBspExDy3vqlR0dEjTWNsm2ynhNcAWl1DIYt5adfiSKcwLrGS6G1Czx
XDuo2RtI1W8sagTeg96fALKafZDCU/AkKrUQYO8hu1N31UCWiUPijokItkr+gQhW
il7ypXdei/Cw3Sx+/g9fTNU3zdfCf6XFHdqW8lO6gtB1mDL2EJQdlnzr5teSJJRI
HAX7qw4/T+rHo8CTcF4Q+6+93L15kuWV6HhCKlEQNbMo5p2gklEOOc8E4Ex2O2X6
dfL/IjXcllTLVxTJmrMTyORqjSj+3lVfvcAqXvVzpiDkP5b88VW69IoQO0z4a9TC
T7T2Xw/c/dn1kk8YtYp2C6rsVO9VNNVlapOS+/0dOKrWN6VrIUiWLR9168isbcXM
TRpj2ksoJPMPXh8HGkqU0isdpasxccRysrGlfT3VryiZ3tCiZkMAZpYpX3SHXq5d
DHWXxvRax7SUsSfmueWuLt9zCW++syTvvimhNfLFoUdrfIwASLzY7lrRDOIPT6Vo
eCVtoQsnYh6bndVH3bqT6JYbHqmHM79Hh7kxgqiTZSyq1sHOEdRZsIeffn5RiE+/
dU8EPr+kvWTn+YGapRKXpvJ3PnlyUsoiQoKtq59oaVzYHrhkmKQNSHMXUo37XTsy
03k0nBpuN/iRkWW42ZnFz5ej+EIn9YviDN7pL8JvdgpVTZX5Neh7n06JMhE56TWg
Rwg4ninKfuEHqPzsAHl/Iv8ruiQCt8S5qgzQv5Cc0FvfiHaYvbOYhQrTpDh0L6Ld
IyYJ/c9qw1gFDiAIQBB079sgZKDM+Usvwm1nH+0VsS12Vn9uOmLAAfvj1ffo02gS
757Nsezgvx04r09WS4vTwumd7arUfnVkF1Yc/vF5+dSAsAeLZOXPk58lEjk2jqWo
DNgeomdLNILkcK2QWZFwtDjaJM381EwfR6S6iDWOcDc3+0BwOarzOWj+UceuX+7k
CFtcvL+bBvu7uGyOhii8fFuhTbz+qPYHzvv1Lr2BXz5ijsl/+n6dKrelLzHv6jWr
uGk+v/w+wbyAEsClzFbw0FuCXy/uRJ1+mxLvuxtx+0gAYB2P7olLyzWWpncv4BXF
05bRgsrcCs0xQiprleIha8S6ii2sK9wqMGX3xOMTYHuLbK110NwG0QBVNUJ/F1+J
mEwjCMyqn1kk3NhurZF8QBB5ynD6z17EOC5BL9Ll7UHaMwbUSrQUwr4QIhzMcU7A
KgIj/n3BHSSGEgu38rJI0OAgEk6pWXNX+q5w48BGKas4CzRrbxcGpR/yfrQWf78G
pmm89k1AnvbVKK4FG2NlY5W1cSTs/bxEu2S+uqgDhiugXaWlJXBBtX0Jwr0A2qdJ
J1MB6pmXhj+kHKQGe08ix6xCt1s4/9Lb/TcGH6jdMfhVx2+0tXebUUWI/cZMjPXe
vYApTKK6acW3gDH5CE6cnVC51+/WE5YlzcOr09V1gbMdLxf62YTbp3Jab2Enoexz
hpdYgZypxYPEGjX+McWtjhf8kxEbY6Y4x/0CBvpZZTKDKNCy3uhqCdPTkGKN9B6q
S6MUXC6MD09Bcdfo9SQKpr/fxHGI41ZuZYmkR78E30ydgbD7IVIpyuOL1udthECt
vyc2451rQ0REtIPNanLPqwIGa1HkNY127pbGDS7LYDmE8u+2d5XpvGnTj2LBA4yu
EiXGxfaw6ORA/ikePQzVL16k6f6H0W9yMgxZraJAT1rdq5WFSJz49+MYUdh3eK48
tWtloql2zhGiK+NM9ALVaVAvEg2AERlEewSTiJ4oF0cVWn84Fe+AHCMPcYhmP2rG
ckmBVjctHH2fmQC5z53gayKoZ0H2vH9esK7j5wIgFiwSyjDEACTrKKG/WUjwc3GV
rtZhHEWqDBB+6ZsrEs75gTuQ/T8e6b6/JprCqxHIUzZxgQxyOVazM7t6GF1VDYS6
UR4YFVyzLEE3aVPOQZU0mLzycBv+ojfZQ+DR1O2jmgBYdAQqT9Q1pzt/w9BEZIKc
2RazMUpwvoGlRjGvT+hia0gfLcl6pyFjBCubKw2m0CluesIzz0ipo0EgxI5+v7Sl
/ZqNB0Z1PEsHnCdcPCJPf1RMfU2FtaUEHbduh5NJRlcsGdU3EP2MNFHOWV5kxkFW
TND8dOGdsQrc6qmjYcGJYmqo6aU3QPOFoQVLAeh+uMWfw0g7+bXHGua7QxjDdx0E
u4mnBiyHOtkgKoEund6Dt/h/6Bji0uH09puulRpVpFav9CG8+p46Rs+61mBVFm15
hJ0NfGryPbdFz23pWXuSwxPbQhVLy3HkfDcXcpkTbkEwea4PxpsV4OBV/MTTwaB0
2w1oM1Ji1eXhcGKGB6aPV7gPL1IIXOvLdqzwG+rN0rmO1Y3Bn6OJLL0a7tqvr6uc
tB9mv56bmFckS6KU2BbFktxdZ+ID3hMf0EqAswPxUS0+Wtx1QDsrd8o1ntJJwrKL
xGktXieW76yyEnIgmAn62Y1qDZ7PEVjg0c1qRSvXt3DoWcy1GmzbaiuOVqfOUR7z
vhJjtnW9UI3tWgKxWBY9yuMdpTfdz45WCyblWUs0bo8nHfw+qnSvcfLB5EEMp++L
MxO0Gt8vGcBHgVsDNRY7oQzwV9Vgw+cmpz4yGMF9N+L5K8s2qwHOg68kYyq2KRbm
4gqlHuz0YhP05VyKkfwUWjZCopo1J4xbDw2KrRdn6sH1cKQhRDNRVR4G9V+kYJcB
nI9Qzx5CG83VOTG1zKZb6BktgygBjm1/JlV5yrmTl1jqYegU/qodkRSN7UnBcCoh
zgshaaeArxr0nAP7+hq11RH4O/HOcxyYmaP2pB+DhM9aaJB7y/O7Zmkatf5pG0Xa
0rZd1mnCiF6LELX83oZssNpdYzSbjl4+fFKMU8nt1hjWmMt+Y2WXLjCM7m7GymSx
fZtLQR2V7a4APsOUDQeIWOVVStWs5+y1Akmk/w4vjG393yQp3CjjxP3df840mBBP
N9VhKGd2JK8bt3lSPaT2YmKZmWGBwYe1Ycar5dUvx/VNAaV4ok7f2kHHXTQbB+pK
zY8xbE/Ka7av8VmJlOzesRnHOfX8WPusH1n/9G5Kk99d7GE3Q0J9LsQ5wnJlGplD
DiFrgXj2jJe/89x8tT3Qm4Nv24RqJLT5YzQ8Elp8GvF5fk9F9TAW8m2xyTzw5e9/
DNLJDxMgkBDiYwkyQzWtjI2G+TAOwlMlVXqiZCMjELZcZSLTZb34PjshVNYeiyWC
wf1PYfgvGD538DMZ/zKpHrpjQ+78uE73IXBwgur2M9YePZbcMNa3gMfWNbBzkE8U
tYV3FzRaozOUanv6DiR0K9dQax0g+r7B3M6nkIMWWC5+YzUMu5LBDZLP231cv23R
LaICmqImQuTGszJziJyNKPorqaSbgv7fKK+epKSuBpYkzsAinnFbwBIqwxi38DuW
ZM5UC/qtMkfdacHEbPUjGT7VMViFrcODo9M6xI9zD7xszssaAJyRTCpx0ZbyyBCL
eXFEmFzBhbJ0ZV4wul5J0YeW9NGnV2h4f57U39b8eb3wKpcH3NxH+sojuOHkD7L5
kpQ2kCu1XydRTkR4WWnLdaA5v3uPavIzdWTZZnNSQNkX+9MlDBK6N6h0LtQMuow7
ntGNamA80Yg+D7VyHn8Iu4/6tcIGq1/L8ETKwEuZE6yIxRr4JUD7SzMwIZHlZziM
eydzWegcpl0w89RgPnxbvNu+5hdxtuCBpb25C4TgN8RoBUKdlf0esWuj1OebEcpz
TOrZIYdXdHLu1eo2iFo8RfWfV9C/PgKx83YXm2SdQrX8e6qvxlgEnK0DUKqTnXS6
1c9yVWhr4xko0H/2P2ryvhYf20W6JGCW96z+42IEfCwYnx1WkKgkAkn7N8icvXnd
DN3jRUkJqlUNO1U2CIJOIYJdKp8qrGH2N4YZ1b3OVno1OMBUU5FP0eXmPz/VqD2y
E6tj+SJolbDchg+AFq5bRNFmi7YD8pbLm3rSCQKKyyC7xU0avnVOnTbx/xqda848
kTrO+BmGSt8+oPBHbZ7bv5WBp5t+V0H9lj15sqrpoh7CO8pg9oeDDQMaYAcH1Cpk
pKaJJr3MccNq2i9f0wMfXO5E2x5OJu6CfKiS+sMdpzSlSYEayen6eGujmEE75vWT
naiw9WLstrJknEgSos+Uq9Zp0OmUfavZMj5lNgRzQkb6653gg/reKPdz2XfNV7sc
zwDy62TmaveZJxbvapDGnvBqIEqivsOd7ttOb3zjln25J3MFj19YL3tDMtg01Qy7
2pEoOMjGqjnY35vw32d5wP+r7ZizEqQX+tA0VntkkcSAd4V488zY+kjkrdYro01v
OECi0xbqvl+q+rAt5NVP4JIBOSvMOo4j/SRdP0zNqQxcYukVrt7LdQevm0qSuQEU
y98HbvU49Wz6Fz+KET1a1zbEbkQYpQKB2aUthqTv3OPMtVoGgKJvY/foz5kBStaP
UjfRIhP02QE/eqvm+YujFHwN64ecwE26KhufDU2A1qpFqjFFtgp3Yo4JmwW0xFqE
JYjZHFtjPN3tPfXLHs23XrpSXtP4u5die4Pyaj+Z2MPN2ZxOCn6GX3vkFjqhYpRv
7n2RNAhOrCg1o2bXBQYi1PPirKMqH5cVBs37M3tSClhdPzoPPv+36qTAFmbH6qPR
+bnLRilnLMTx0SRJhFaKgM7IucWsM5WQOZDdNTNzODw43SwrXIx31yeKTiXfD8KP
BiCwDcgHYi9inazscpqvenjelcqFs8QlIOgNyPMk66JqJq+SFNph/2XQJjsqFBxC
I33m8UWRMD9Fref++euxpnMPeJ9YLY2S846LBz5msnyN+yDe/hwjXriOgmgCGE/0
7p6iRzNGCG37vwbHNOFN2qWxlevP+MUQh3XI7DZMO8+KHUcaOgFhF+IWCPdiaFen
OdWvHvXk2+cfCN4EdS2fk+ef9Mk9+KTRW4HETk46GKY2vVMZW+Uzgrlir4vpGCow
j0RQ9dQ5q9YxXkBygLA+QPwtcsD86AOaJYjrZlNtBLLkkIpYvRqwxRktJ+y2ofRC
JqerR5rrWFc7byOPCgZioKGO1qjDR2tryutzjngmdL0eI3lOoV25PMEhDJjzzAYt
5rD+4inKu9lUaH4242a49Kl04f//dMdUx5/U57vaGuxb6APbA0wRLhuGQ29Cln58
xV/fMhkxLF0G+M1P9lbEwJnxVwEsbZ36pfqxLfnlWdZE4nWc25c2b/v6zvHsSfgQ
QRtmt7s7h5pFkgvTWPC5Aw5I308QmkM7nkWx9Z/Ko5ctR9kKgm/JjJd+epczlz/L
+a0duDYQB5CM/c2XuLuiZFL1QJ3PilId+RlVPzQl8w4vT4ooGuZJJs2YOyMuKJTV
0Y4Gk2ypr51wyEP4KGZWk8On81nzBf+W8v7JHS1RBcnV+tB66OXVUbq8nWXP8BJA
3TZlBupK4Y7NtL/IPBnPq1iCPdSdt+3urn22Z8Ka1aVHwTGVFtv+mqLhow9WJwOz
yE/I1U4XpChBvGrpLresF6gIyijZPDidRetv43WxxQgKjyPzx8tVTjQWjGvFhN0T
RK2P6PTa3+Wk7fWmHI6sZL6qOEnjU3dq6ZUaeP1elzm0q9dNwLRb11I7dd+bSqHb
NSq55Wm0beB2IMkdD2fZDYqF84KyAro0VQz/K1KgVIMwzSpdhcRidMAF6ucneHSJ
CBhGwOfJTRgTQD4cia1IhlHIifCJM0pm9H+mEuAn6Ri6VAKQ9eudZFSlN0/FpRma
ZzcrEo9mAbNqpag+l/CSgKgIlO3XYcSgKRToQJnFX6xhIH4P3UUOI/5gZbui1HBK
dOwQU5FoRlo9Tcj6Q1mdXQf/FDf8tivvV1dmLGTQ5Ti+wb/RvD2FTrhOdW4zubK6
7Wa062dVyDpuxX10e+nv28UdzV99mVrUivohey3eWebYbo0MEcNo2xl9k7+R0hnJ
EYOGwB+qbvP2uQLWrU8/7W8c0MYhYYUJhjCFd2r7tdHkKsX6kUJ9TNv8oP93fTqa
UpVy2GSDUZwuCRfQYQX66fkg3pf311QVfSh9MX+J5YrbdCmClQS17ufSVmzWuzPB
Giv16UYDOve2mrSVfqg0viyaYx7yFBrs2noko4SnyDb+nvqMm/+LkDtJSTdVMl41
TMfHQcIQBr4SSgfkrOf1UvIPeT78MJLXARosLds8SyT7mAFkb90zXkSVWib0aOAz
aZ91kQBchRQuvr4oLuirsxWEctCixtzKTbF+vce4+KJk3OAtlTqNBSuXrm5VvAgg
HEypqhOVRDd000wMzyogPFD6ZlbLAhQZjMqit9keL1/M9n7ZkNmbMy4h9SErJuWa
pbNHLpKXwzEImYJHheczDw+nIh5gwFGL9aMD046zP6xvZwZ8AhtuYTUM9zH+FiOy
HXNQzZiLqovmKEkLolrXybquW79uXdBCSSJ96E7Y7BOnC6AmB1sm2Tkb2C1xD0Bu
o2UsLMlA57SatV5k9sH/MvBL7pfy0wuhSBjg7Vg/VqeMQPiaJugJHZBAR1w+W93v
NiGE9qaKmWJY/PQf9aAyNspvof6W6hScDltXiCZQ6sbrSemINvbTDGAlfNyL5AAR
hMwULz6jm8HGI43qvGcyESXeXi99wV13f5P25jbJTfhdtvbzti0uzqmu0S5xUpdA
XjP6bq7DzK6mN4gX+w/3ITWXDuLQHmCdnsZLc2FMt5jMg73e9W3TrW3woLRcHjfh
QjjIHR+V+ibl3ygf8C3JpQqDvD94AUn279nn8fBqai7cgxZvi4J7HLjUOx/cfkb6
2Cq9XWZH3Z/GxvvkbiIfIwXpVQ/wuVCvhiyWxCys+jx5j2lRuQE7hLgkNYfBR67S
2XesDOH7fkmOhhofg4TMSER+g3T09dvMBYSS0MzbMO1kVIWQbrVp21yTdeyGSDtI
CANLMUz4nsri/5HnQ7JxdtUa2Rf7k/YRn93JenIP8s0zfB8qSUeeEGWvaz1JZbbC
Dhk7QSNJ4QvVlfBw5Y+rn9kZkLK9yr6TOUCWok7DTLcfHhNAEXE4YmPnSnZIIDLq
D1kbO+l2wwI+CDnHMQXRWj7YUnFdAl90EBbazE/V1V2rAw8NPZ+Oc6/sE7oxTxny
lDxCO55x0SmCngBYCJiONRSM6wgeghHPAvbU2Kuzz3X5O/kVgKilfCtaBAqn6eeU
/9Iiji1NL7B9mXQkKoVAH4sLehndIi7Pbn+bASTels3GgmUF1Sn8aaZQYmy+e5bK
djH9iLPiNKucKwQJxWGPFtEGFi3IcvIjjADjWD5yC+xRKFVbW8G9CpAj1JMmM4bJ
JSbCB+I8lcFwfdNcsR65P5h2UPCe3jNol38gVl5abbQscdL8IvsBCn9XQlU+zVeJ
tRPghJE6XPnhx2kHQkCPyKpMOLg8ZDpUMXGM26N8ktmmFxtKtpNvW3Wy62t9QPUb
ZeZ8l8iz/V1otBdywV/hgZ1sbY6reWTuHWmbybPm4B3xwfs+MCUEoy5ye9LbsgS/
+1OdmVnmb6XTME0uyGnTD9ZIct6ju9vNRVo0ZkzJ5B+Y1MxCXL3/IJmUPFj42QFt
2tew3hCRwau9O2wXm5/hZUuftPfqYh5uobK3goi83D+I6cWas/uiy8vjwhv194O1
WJv4C3a0i1wfqCGLoB7TF5hH5ti+VOT6RmOab1g8QA7YufEgFDPxTnIMwEg1Qu7m
WXxbaPOgJ0d0AockXgsm9GnLoW9BVww9U2Fojhrw4BqyclTZVNty1EKRiPabRNsf
AVm1YbWXqhWSQD4hMPhl5lBTBHnN4ggnoz5Afl9+m0cmqLb2X63K9kh9GSHad2xJ
Dyjn+Du/xfkhynvAnLCIzLMIB1LtCBy/Va4gGXwE6X2tKV5h7DceWIU/tkdbOkzk
K09z+KbMewn6rnji3NYVjgq9AQegOxYR67xbUX23pn+VLekyHLYxTGrKSWvfspcQ
T43eWxRyOhJRMXjB9KqT7qSQiuhDmC5ra3YigktygphW4zo09P4WbPc+D0osaMBJ
QHGok+dpsQqtjAQ4NC6Lzv1OCED7snE0lVvIJyFSJ2tGABd+ESMVXtrV6oIbhsHy
vFWtGbVg5dpNEmUGImj7iCqZzin3jC2g8H0Pcla4FwurQRDkJKHkiZBLzrdwH5G6
g784oa/CWWVvtuYCOrE9YFAxrnvxumwopN+hgWVnHu49DpRYUHpVGcwTxA/p2IC/
TX02IYoSGO0YPqr4OTxYs2mGg5KvniZb6+9Ejl6g6D06UxMFI/tI27PJN4Rj8YVP
/YcNtKKtBfkB3TxOGs4a/fTJRpsI97YYHqPdr1VlMhifuYtJFQhbjapoXfXdM1wS
44nhiEv+/D9r+DgV1wKsygJ8x2YOuq3EAGnNHsfilb+K/g5m/7oGQ21d9Ag+DrnO
2tXwaBSMhQBAj4/ZNB0KuVtFabK3770iPcKZgMUsDeUM8PmRtOhTa4PGnmDjo9z4
s08dmkuVgxhLYDcuIG9UmlraaJ4rTu0Ai3+vAFR82qdoFC04HlkzrCCNdAQBVbrh
L1ksuREjwd7Fop37XnQws3JVjyL4TcwoOi6Tks5g1F3tctIxhzIecY00XuFr5e9r
5C3NBEgXZMf+hb/jOXEodP5yhUCTYICjd8pEHkPDryh2iSnnsOL+oSgxppIrodK3
cwlEo6S4fu4H5JbkgrsE3iRScl30i205Dk+uHvoPXZnNWZCDWSC7ih84TJ4b7cq7
hlnMPDUVrglb/nzL+JOgXWeo4iKSwKVTvIII5itYutTgPrQ3KGgvwnUVonWJeTOs
1LQfWiWpt3dJiqVkXZIy7Lq9nLIyHSO8OurbyLHeIzt1gChmy1DSGDSUxAgJRZu+
snIWnZ2sjBzaasyyL4WYmLJV/ogHMz8ZDWmYMPgTE09bfOisLtX4sk4kF80sUc0H
skr9bTokqxcCXhCyqOVfazDtNTXZA9Go6zZjPj+eh8qhVQdm41i4z9cksCdUX9nb
rU2kUhN+/MdPRCRvkzqEvqcbHIwgWK6fyoz3eskM/r1e67nrOlPxQyLoMt21GqyI
O1SQezRnD0sleUxfs5DDPQEaFHurYoVRgKclGKaSP28T/B5ir+eX8y+L3ynrmepC
XjCmp7znbT9ACEs+VK9rfiA54f2qMhajWingwWaBshz/QgyrlKUy49+P7rRzb3OV
AyAZ0GcIt8WGMQjNE/HfiZCU8GCvG+p4BNkZu6nmat5Hh5YOhVQiWBl4T9hgXOWm
wR5iSxyo3h9UaV/y0ce/wl31/jHzH34JsmzIgKiFD1d//3ljNLs+WENS+EwD9MDR
wsZlKd7g1rb+3Od7EGXlpT0QlYdiGNcT8Ew6MWpkmhYUBkVw2ysjd28O0YhN5erR
YUHFLNoaYjTOnEa+AF9s8SiQ1AbxnNJbHYUcXFn3quGeimkVl0XmS0h/hAL4w9gd
LimWGBXlLnX5uV+lhgCakgGzqPfrxGKJxKcvCeeJy9PHBHUIaHHh20pqeMqswyp6
AyOJ1kT9PSfqg+XWMBddiDB/CxS/yItOrlPvZk2VltQVA9CkNEqy2Ms350wzlAgi
nu5AEPBHCXGJzwBArF8gx+jzINRKfllR/TVy/O7uH40wRlSxyRZ4JP7XWKVRVDvZ
BA40X9YJAXe51WbzrKjd/gveVC3Ywg5vJim08bGqrcpgfMbn4wae3CaQZSiHffWz
VaRYF51rmTrmVOefC2e1bFIYXu0IitTXDCplwcG1VxnPA+7zwbv7H60Ck6560H7z
4zhqLzIHduzk7iVXFSGMATQn33mta0+ZZqDkb1J72fzjAG+/Yp28Hgmwc2VBSpz3
zYKC1iRhcSaTAsj/GFoSBf+p6rvyGG1t6aLL23Y1EB90a/moNnqZVtbs5EYoH4fF
9FtjA2kU7b97YU/7BmNMqmCMeXAsjqqUNqO7r4jfPZrBGRHLwBvATZ8DUHSH0Tae
4J6pJC1UpL2aOonSZqo9U5ZxkD6IykgjrNNI0Cm2/1jBY5/AtC+ec3WcDWwbfDmt
BHvOP3E6MkEaFXbAFms+BGEHjq4gzmC7Yd0YyB5Td79xy8PS1Qwjbn8EEZsW5K/B
3B1+h/bJvLJPFELOExkEs9ig5OymAvXZ58hDxGXLsskOW50Q+MMJfdIJ8ZAkCtDk
Ot4aIqyl7dgdf3kdgx2Q0DYUeqnbZnQ2r7JsRfnpBflMyoGS91NjT2oObYG6y5lE
ywQPLoDYm4IKB41VWfDd2Uht5sJYRmpUt5CgB73234mxv0acn/toukCDb8M76YLs
23fDpka749lPOqmg9y34yEBQ1dzmj2boo5l+zW2FlfydPRN4STRE6OZgdANs0ePV
fXbPH21o8fOyGFkJcmOJqBUqclBnzpv8G7vfLR7oi3flyLEQ4LbjOfy+xPdNlUSw
QE0eXzORPZfxHIUb0fi809dHo6EG/HpRkxhR5Y2304VCUUW62Od9jqh3BTEUVcuP
WciRppeJeSPNma4R+Tqgtp21IzMmtCUN6anauKEykwvNve5qGvz7Cpzl0AYIesLz
zQbOXNjWbnpAM0vI8MsOQGuH5IqeioSW4m3/870OLAVHZ/aTHwv+W5RQO15rlJOh
GWItX7ojlCYwdruD1i3wIayJ7tVK+40RWhYsxQODoVMmjZiXaMwqjDX8+/EmRRuz
BKUr3t1zwlzeKLaAGKVPu8xOh/AGcrsVbI05Ss4Lmis4I50c2cjaBeZ47h9lKVUs
6XzCrnyMzZTY2sFga3K/pOYKUfXMVV2ImUWuJ2xXeejpTXuGyK+bs77DFIba551N
mvzo1czyz+sTX+WQ9qK0wzLtMj8AH9RmArIiPDUR0U/BwH4N5Zs32hnLQodgYF7c
mOvwPnJEpYj9YY3NjzteLj0YWT1vBz+HpPR1cK7BT8io+24ZXpbnlCPUvpgw0dki
JQ0tOQXvkCghwX++heQQK2fNxyZuQFVrWdpDZIPp0uW/MFRZ3nWOdtqAq7JKqi5Z
u2Bf5Nqt/bhc0+iLU2kHUIUxzUhxSNTgG5GElTG9K6QIhRLuXUfIHeHP26AwLXf+
sMNhVjhWDT3KJnUrlNh2kCDF9z7OeTZFCqADmAbVRUMi72V/YKH+yFDZ2NKanMtx
UYeoNbC4zuz6cACCvXiYhq1ws1DHypW89ZaNMN5J291wEPz8cR4eLTIxF97W3J8D
B98QPFMkh3pFFDBpCFeQanI+ilpQ/0m5O/HzF6bu/I1T/vUYc6FeLj6Yk31gqRCe
8LVpiqmw1fotbEJALaXo/cwMYEuTkzprqirwziYv3ZXfUz6w4Uydiok6xLjAnZei
Ol06KCveg1bwTafae4pe+1Uai0wSSUkELgR0w0x6X+XiuCTxW4tb2nY77pwFHtqZ
bWwmOq2Ttbkk5Ys8CkHBXqkjyF5rqIhfkfvHXlGoQDGU9BlWMEUFB0lpMR1xKIkK
q+AHFXy0AfJtZmj8nMqodd2ubs3Mla6WCe42BAOvtHZc+y/KpcQz2rHSPU21vuaS
bESCoRZOfkYef36cgxcvwRXeNxhBxzekntl+4dbJZMmbAtW0gg0yf2HIwlohzfGB
iad7NhxwO3+BdxBhtn7Rd8l6Opg7OUjYf9q2x4DIR4u3xlpvXP9/HoqKxQyndYON
ojIaWrfuAK4xE8pjcMa3nJajULZP2J77C1fq8UttTGkgS3RFWpMJInjk+/BbDpWW
r8c7Rwd6k0NSaPDA0bQzaShCObSDmTHMhHfKfmZXBeITqJYXSE+WcW0OOE73oH7M
wm7jEJKMtby310EL+xx11M3PzARFUDZbQoIw5EJOAWmAkXAzRJWtJpfUmc0KDe1C
7mM4m7ynUPEcrRFpx+nf9LCywaOyh4RZZnaEnnBf/H48/+KO3g3675twd7jtvYtp
l7EHg/WrzgShmPjpeG4ltgdM+jst8az+Egl6rc/jKkxlfvJPul+ImyCAq81Wd4NT
kBvzGXbnl7UH/gMUklGNPOqv/Gx+8b4Sy3anYQ3E0nTw6xHLw2PW30pt+Kz66BKf
ZfNgqnx/yRNB1ZmyuZedhEjIqqtixUjtmJvr/FRgNIPUftl6axmvbhog7RSe8Af1
Gk2Vfe0Rgb4KM/lgq/mmmsR0oAY+KiUYcThUHCGkaVhWaIQnk9y1W3TGAtzJ4ubd
mNptNbUyAuD88shSoRaZNoo/EvT9Fwtu7E57VfRBonoJhtMEY+jPiniAT7/WCjNp
jgnoDy3UqtcIyXha5K2R7rwwvNLBMINTlOiK82SKHIvHe1TI9czcSOrnhEbn2qfQ
xDO3QxcyKhMWAIS21acHKcQ91cN562khdCRiGLbipGGoMA1GNy8HQUkneFRBtGQK
TemOHQgmLh0UlWReI0r+JSb8ABUFZgUWuVVphBMmf3mVlOAyoS4tZFZoXnyixcZQ
H2CYKVvUC3kk684de9yPsFexKz/FQ/V09AaXWgXJoIBbkl4u9QJCtPO2XJqFm2jj
yTZdoJg6DpBwo1+VeGfQL/3p85IS8EkaLeyR3S3C4myz5mSZEFyhORBVon9AJOFg
2+TNXSCXi1A9bhYw2nJfES+4m3kTRTBdFAa/gDxeG28rFX47mId8B4n0b9sxVulv
FNAHD5nLwU+tWOC0GlF/i/FIrsdV8/HM1A2tcvcedY71YI1rEXIzh4tO3MWna2L2
UJpb0HWU5WHdadg932vEyXitYr+xaTluyV+xoy2ZA1nU6v05u4WiXrS6o/L0CXZV
ILRz4oIPrB7iLU+i7V3+ikmcAa+Thp5ulJVe1YqkvKoJ2gd8oJ1EA3acbOPQZ0WD
7b/fEn/WV71aM5RrtXczN83peBxoEDNpdtXN8vYRKCngMQZumlYShIBR9n1x24BV
SMrsmYACSE6G12s7/rh5/aLo6haCOQ4oLhDpJAztsgyfbBDUfve4hpFDNoK+2gcw
OUFk1LnY4dJfHCvCSZswJvcQtHu52pfmxeQDOdwnELY3k7WIYDU/VbWWqHbpVrv/
PnGi2al5A79Pxl7xtPMMZNesbsaDlXXy3yBQWkHGM4B/adN0IICCpL3cpMHbfUxQ
Mo820F6er4d+j9QY0Lvv91v+xDwRqXpC+Vq8F/D8gksWZ0FFRVKEHEcWqSx1lbY5
R9KnxEc/RgsNff+KqCHhjDlPEXjWMNdlMA6FvVCCq8z7erRhAvd5yXnxM2eGsSQu
CI2SDi5QHo3fafA5mCWCJTFqYl8ghUJAT0SKTF5j0uZwIn7t9rX2KzBOI92En/yo
vpBZpoq0lufNXyv8dwnVherLPA1flt6MJzYn0Y+WPeM+9iVCG1t/PjKdNlEnJFh8
azLfQBicb2BJjPB82KGpuHeIXsbeOyqFN9o2HoTZt2kRsxsEqs7h3tndBT045IIP
DNqKiLHN4cMVjGmy7khVXgEVSur1lNq/U1aC+MSHmnZ5WhRm3agJZqtr99oPMwBW
fRurmrSUhDy8EXH6JW8Nw5XyoJV6wmWalNJNVB6q48yxrfux53cyqwuAoyTuKSg6
77roMzKd5ZxNj+jJOoBX1weUyORdyM79pd7aMC/mokia2r+YpsIarUzzSGBBVVeF
phnC6lOGzSqSVKA9Q5Qv0yUdmsrDkZrhCQkvi2gXQOf6fkl0Vub+GuHZIB3YmvzU
giqfqNxuVF/87O6m8jJLCIC/RM7yl2NnhZI2rxap5W5gTIX/aNTfSg5jGK4zcWV9
KdSaeA+SxHVckdO0Gqxl3cNXRJ/7n8asusoVmSWJ7w2J+FVXzTEWQT7N9SHD4acp
2/cM9FlnQUQgYTejAc2kAVjxAY/JS7FeXluqlSLgM/4Io/ab+kbeYX04zphnHwaE
+dRT9bpFZqmnDa7j0O7zyWfzwQSusnfBp5/7Gn/WmtHeqH+ja3WPkaeyp1hA/lND
VOjSwUn1dRPSMMfgZMFTHzquW1VFBXDvpbtCevKpOfMkc0Rp1ahsN7rKsCGpoW31
YaPjOQ6uxNsNFlGjpthpRjohSxiwrDO0CqedUd99rJuBp6YV+J8jgL41YBOCYpH0
iGID5ZBy41EPls1i3rPaeyAU0TYcfWv0ytDjgjxfJI/c1cZSQJfOyviekHV8+iwB
A5Ek+rZVedsPEaDWfUzaNXXAPN+zUkj1qtG/1BrrZwr83zvW1j0q7ZFhI700aWvq
dH0hIpXlP6/KTAldyK32IJTzv39PR2LqtOjdhqtS86reQ462FMiMtdDnwq59sUaU
RT2hzGkMXwbNb+6qCzefNSFs0UOLsuEnc5DlqocSWB+bh6n1JVYrWk56CqqOCKy8
B+tCSy0X/igoC4CX0qXiqH6RrUCo39chlEIQ6bhMY5cElaRcjvd++A5Zf9njSjcm
eJQQVlacjlrCMOObFbr5cuMGoPkBgD9NCpMIdnA/Z8GkP24qBbhMAM3Vt0wSGT60
L9/HR4+dW/DheXEZFTv/MepoqHG8vT0dp02joK76w9GXh5pwoX7M3da1kZSbmam1
JZe2GeP2C5yYQAOc3UXRuB1wt+zeG1bhknSjEadzL7BxqR53mYNruodM2Gueuh1R
ZgAwmvLe9D/x/0znHbZrLKJIz+gQEr4wFXXLWkqNTxSB6ABrqtQaJHM4RqMl0FM1
04+hkOrlxJWbce/jbTR8/atC/Zni8tDIXStT4LbBs0SpJmYDKlmCMkT0ZSnI6oP/
frAv+14XENy6lUdzq+NRJ4wyN3mQky9q87ywl+OIA+ou+FCz186NJe6H9CEaiCw2
rA+ww2TFLlLQ0pMi7x3Qp5AnNVBLMr5e9mqA5R3ZNJRezR/eneBlonjBC6EdmEGF
wfX8pFU7ZD8sGzUG6En42x+jBk/O923TeZWOHqutjB+dtFJNfPLyP/hOlDwzC7Vf
Lt5gkK/t811iriU7p0xaAqZhoHKxRlpJPM5wRFdPRJb3uGjbcm4eBB6A5iHWKlLP
ZZ6WDted4/SaXJYSJaYPRlItAJCHOs3xnksCt/GZWMgueqWTtWxD8/JSNlWcHHSK
Po8AsLiBM6x+utjos3FrfxoSTGwAzBkYhdNdvF+jPxOhllAvbbAXrEmGNWo6Caft
aKi8idy0wH/UEDs9PCVA6dPxAXYX0jDihwzrBfG2/hny57d9ExSYWEoD8CQHLdst
BXxxejTl30LWGx8atCTLfbCo9CdhypAgtUICrvJeRv9IPwkjrHzax6LATWs4F+FI
EvHBCRszd1OvucreDjzp0WLX4fMMRzf8y+cJNb3MHjPHzjDiJh6LnbtpSHU9EPIa
cqw6rm60d9oiI106/p28mm8iiyymhseo8fsVs5InD3Q1vwxT9Kno4R4VKmAJbsZM
xVm6qqncv3yfAkRELUeJnreua5O5wrSeNHbyyc4hDdgk7S7mb5JoJFkM9ua8YWyF
IKuO22k9KYGNRdB7FmJXn3njJvWhwxeYmxPuSHrN+eO4fvlZddK6FPHBWTF+WfdO
EoZTipjvFpgnWm3QELmHZi3mOGldZ2+VJ5R44RJzebZzgLy78NCfIbxTCfMwVRRJ
1AKhSLjEMgkKvub7F/jX9nseugRZXAdgBgFPN8biK3xbUSFWQIS/DuG64jCuHZCz
D4oBtithZEzIWg1wrkHybV8NDAmyZoNvkMEFRp7uYUyciHsBL87QzeRFO8uwdbLe
lG7hNAjYGkdm2n47Au2EleSPcPhlDyiEgt4Rl2oUE2rriwurxl+DOKpBTEEXoR0j
bS5L28yE2fji/6aM76bHdMMmnL3wJu8jV5T1aFley9wr+pD7N5jTHYQdZhj45UBZ
VmV/SUA3BZmHZo58I6jlZr93wSh9UXRZ2ZwjcpUIyFk785787LmmvVMzPcD7IF0q
dkuli99QZTTHchVlEzqvvTiELDybDCfrcZoW4sDUGFZzmjxXuFporJCJ6+7UXHBX
e/cYmOwHngi+sAfKRfMkaY5Oo4AnrwGmVHlE/nQZs3enN+mk4/nLNegvZhIS/I9m
zui7wMC7BinqJ4QDfn4z12dJ64AC9Qdxh1Z5sY4YTAXUgb9A+MiflsGx9vwHblN5
X3tdICOCwCAelRVQtP4PXJjK8s0DhxbFs1MB8WLnif2HxInGY1f8yMJtyYLkP89+
4h6VTN7buz1AI2fqto/lmdvx9ZptaUp14oMWQ9WN5oFRV+E6GP/BszHKQdPRNG3y
yhEi2P1IqrxfjG5yICC7dWU1NLj2E2A14WvJ4gu+kmCfyFnk0jzMjMt8GtL7GNtF
oSF45Su+DrUMLqNPn2ftAtUlBnarYfua58DxhEwd5gQ096dDPSXz4yJUNg4MM8n5
waaN107g5RUG5G5dQRb1bW3gW89QtZXLhcBNiQqbOng8PNDtjLoj+j5PzsNS8sjh
xZhNdJWx/+aFJM2ZaK8uR3P2wKAYHTt3D6fgFkBifY7DsFaUqBmZgBl/Sel1lrjI
yOhc3KdBfPVpjKaiNvB0lZIGzYvZ7d/TdhY1tmVZTPL8GWsoMosBhAIlnxWMINzc
Jwh9Ajw8aXJeomERVcABNzu2ySxs69dHkS+YhkH3rHOTnIB7ehi0bjqDTbCJzEdo
6rD6wHZxLc20qPsja9S44AT2lJIa2XYmQ0jAm/ZxFuGM7Wft0NiCPi58Mq9luVzp
zv/w1JloscCs04Es4Khz5rI38iCuy44T4fY6/fAXv7XDo5+GoDT7VUj/lPFLfA6Y
7gSZoTAd/zM/H8tCzj0/Z+7VLc1J1HGyVf0mauRuqOoWS5tA2J2FToy2q9d7o1lV
FZP6CWiByOV+NMIYLYrhrV8bECCxQuqEAkCRiApqFu6T0fEPxK3L1kNHt4nTSv2r
coZbeKLzrr3vH7GzfO8uIy4oAzkpFZRdRGzdLgyOG7Y/8L3EhytQfqptPIR0Hz1x
LFP2JtrR491S9ZUwmNbx50CmSvQR/AeekXAZE3J3UqQRYohQGOBtfeaGa6rEkHf7
Er4OF1PVjH5c9Dh4sFchqtpNNLpgl74jtkhXMAamhLb5P2HAY2CNUDvnr2lgg9s6
ANkta+sd0hUHUN6sdD2tuAGH8a2GkGOXEcKFQ3t7lzTavs4vImfGJjTKzbB7b8eP
3JNBVE2eLonRCxZ7EUgwCrcCI2ohmrMmsPmmd6StYookOffq0ivaKoCtsoviv2DR
oASfJ6gckjUTrfzg1nTEzZ/nyqUqsH+6hTy8cUSdf2xvDQZlFE+3+ezusq1xi6G0
Mqpoz3+xHgkFc4nKbNDMDnG26jRV1QzXo++LArlQtm50y4ga+/61a0rmtxtfAw6Y
hO/OVrBCONXz16Rhqk00pb6gwhMQ2S/o8G0fFXxvrPwFNGKWjdi4CtTJNdII9ewP
gjgcuQazyXMSws0G2LYbuMgEXy3taNXbKhFXHE4rpoGE3mYmVSQMKtsO0xAJyKkA
EAPF46YRSTpCjSvMQppWE0bFFJMpVWbXDnYb2ajWQuQEOgXfS4TFeZApQ90js1M/
nVPEEg4gsYGmAn6Gv0yA26Hyyj0GdWtRybuTZiDzZ2odro71a6+fgZr/nxx74PA0
AsIivoCuPqxgwbXFho0tnijzRBmihKbaryhbtos7ZV2G0DswPjwVbJoqXCze64r2
eN4Yue0are2aZ+8d7s2PH1W4RK9uCM3PcU11t08j6wChU0q4MLdT3TaOKUkAlw7E
3Nbym5DUPQics9NW5oG3Cp8xDu5GZvQCNL4EAdT/6RX8G2bfHs7ccurypd7ElMQb
QdUrQKuW1C2nlSYLvfO5K53LkyJlY9G0WDnOj+SgQnBEpoDKS9yKXDkQhPIKQ4nN
Am+OyrwR99x5retoomz+rmNyGgn3pUdzAzyz28a38K+QDWnAE9bigILepsg3jNqj
Jc8zBwJITjX92f14r4/VtG8lOhy0M2ltUatUwt6JYsH3I4UQ9t1hl+hsXdgxHXvQ
6IoiGYqrRQJHEwNO5FigK/K8pQTam1sm+qJjzggoOOD2t0bykYcmRun/OW+IjVeE
AiMMGnCAqYCep6N7iQqSu2MkqatD4QdzQJuxGas1puwbRN3Y9d1tW/4BNRDmtxnv
TuFH1cRwjB9Xbqki87PnxZVrDFIUF5GUoOZPdQeK3EvnzdmkAZh13hMGL0m+zExs
e1E1Xfoj1EEIv10o+kdlva3k/Rv4VS6SyDd/1WoUt65/bvXIkW74aZQRjwLkS/Do
qOHMfI0Skz6+WhdlXVWedUxaokptSIPkIe2kkp677wo96fEg6vm3xBVXcKUkKzKT
CDdB5/Tme8TXhNAy//2CiX9MjTIGF52kyQZAKckc/SIOiy+MprtZfDnOVv/XU4tR
M6jIAeUQn3AeanZ6kZWdjaRrcldAOeWXYTVEA9fqK7hroWbRxmwXXhYpseMCFm2A
QEBXJZ1f+14L+90/Bir6kW+cDb81Vgf4Sz+V7uygj3jSrfDloacnCLcDOXYpKT3y
lkpLqxw6/ueSkWLdMbmnXnOLiYpeDYCr7hyc9skVQFZVreBCdVwg53FKEBhTAPrs
V2BKkK3zl1q2RCCxZIkF1+awCkXC5srp97pbaTzhIyZTiPQibAU/0He94MFV6Vx7
Jz7eblfiY4/MdD24hP58rQEIVmaV+Bb1/QfudyMjiAF+5/0fTSbLl2AjW5wQ8dF3
EzVqo55kcLa1nj1c6Jhl0YU8+m+CfaYwojNn0EpuyeZo8Vb7v3KbGGSXmObznm/+
/99HHAyMdufH7Y+PSLsRSHu9xKn5SI4ZkG1GmEoHPfe+bXL9nf9IppHMsfPg1TnL
EoiEg9ssPkq4s0k7Eg3bwpnkUyUdQVcApuZaA911acnrUY+tkPgyX0Lhy6Y6VDch
E2ixkkzZxSwaTAMv3JNhhcl9IOvKDBENNp4U/3pVgiWrMdQhC2N7Dl0rwAmMuFe4
8WPgeUhC3ECaBP2HlTVmhZJUAEKQg9KnUwLnENPLkseE0ORml4vo5eKZiByh8QWY
ghMkh7RXuFk7KCnsOcZCnWLAM4Tb2KzXHBPhcQa3R1x4Mk212F5mJMhuCAg505+y
mG+4YAbItNElmuLYruWrAA3H+RXaOyuGUHh5V3iH/Gv4KhUNPajj/1z/1623lU8y
DcmsLNd0R1+1TpfAZC8np1tuSKyNq0JaelwvLYHrSBDE6CG5WyL2UXhr522nwhWn
QbWGmrvEHMow+R8HBiBhWv7Ju/POCiNrc6ClFHwKJdHL/WjTtFX9H5kPLCcNnwBd
fauRJZrCwUzDTPsA4bHRPjleZg6hesufL7w2gX2PnTcVBdhCrySKo6WaTJCV47BY
E9S/Av/na2cLKd4BA7lfQmy7zha0CzlqluKnu+7Kwd8z3fRPqaWoR+yB+wHg1jep
Tz+j4pzTfKakx+WvSS+RzBh5ADpE7N4hrfmkSnt1yxNUmwB9obxI9ek+9rok1W5s
RcIabl2a84FIxkV/ND88GQujpzTnfBU5FGJmlPmUtWERSt5PVc+SSJKc+jo1SL6K
rh6wY6zsoXkiNxD9e+9dG1NIQvzpcm2eyWBRYYXLeqszC+Pwuo3eMcmcCP1RCUh2
2ZFof2IBxJAxa/DOzwCAEmkWcdYTAhR70Q+sTfE2VQasegYbhOkSwEL9ea2hcnZ4
A5k/3gXzHdA/aXF40f5J2wM04igVPEEwGXI8LgrbKBFVUDj4epoAnwXznvhy/uW7
qtq82dA/M435HkfdObB7n8oEMOqWesOGvmVJnnln2lGGnufAWSpRov0U18SCq0eV
NTZHsPRgyjBtfSQtxGzceWuRpRDie1yK6K3bbe924UiT/9+YwrceTu4PGFN61y/A
11PwX1NLDNAtrOQYX2d6vBXfBR4EeTkyR8yUoSV26Dwbu1oed2ppYRerVL/ar/V3
dWVo2qe5cVxWJSrTJ/ZqP8B291yyUzMfPBMRzi9vxtwv9oBo08nAuKVGVJdn2HcO
0tWEDpZhmFNNQWhSqVlTTzSwyn9an2B5i7EUOaxZxCFflL6oifefUd0JYtkEncJZ
ArAOOJcwdAY9Y6lkwDdqZ+pxggnhBTktkaRYpXuedJedyQseY2EkYC7vwk968SAG
xSO0h38J3je1+LoiHIqy5r1LBwJqmwrQ6EsvC6PqcBEjdwTPjG2HkD1gqDFZppCw
bt1E8m9cq6SEiHOEgwjgpZA3f+PbWa/FcEvH7Or/yfQ0mS7pLBg1647ZQlxl9QqP
gMln4K962xmZaOpRqYgJCH2uZFMkALDESbKSVqbeIriuTAiMnbbBJfsCT6QUK0J3
V9BWFyKUHBgkd46PkNPIPQuZCSgPXIQi8k57afgzzWITwOcuUcbFYvOYZd9/jnHA
zCBcrj31WcIB+Q+GzJJebaRd+QOrkSKzDwwSYeLZnWoYny6fag+rEKrgr2iGpYwY
D4/NSAqRhycUVfPqEQ6AGU+7VUgEceUggH9TPENRzqHRgjRsxPammtNihpr4lYvN
6IGTR8VmzUXCQBN3aPTsOtS320wABm5K6n5tJwmMmWyK88g/RVLiWeFttiN7Wczz
D9MPKp3Q32ki5yXV06rFonSKl/Vv4S+guDVKMLxVKSFpfLPpNdJqun5mfCOPMyC4
woMJdndnQFoqhYdJcd1j4vJVWQPZKu92BSlzAyv+iUdd4IB+PSajdOMq5xIBOAcW
e+WP4KBWZ5/RTF6wMe66yl7h97A9PXoKA1mCp/9qv9kQq8pPj/BbE/h+2hXlIkvP
DXgk58IdjMhsewvpxBYhuVHgxcOMheVVWZHIfuF7mqIGnPxuTHWTWXtsGu6wXNp5
pibYELPfuTuul61w19BJbsVcgDaPLKzuF0v8etcXbcrHbM+hPW70IR7X0GnItscI
za7B0yP/ueledHEYkU5Qsmkt/Hg1X4eYQG9OjpQMakE3J+SJN6zWz/zPMXbfVTFR
p1cRtjh681GWwP9Q1vjvkcU1aOPpj9MQtQL4k1rW7dLjgR7MIkjysayIeync0rKX
jisSEaCnxcSDtLyTUYK+YK3K61pKPUHI5P4QLGAxgVd0YWmJvtomGXy4kHEwT6Wi
B5u/moMSHZjgs7+5PszjxcaybFjL1oI3FyBuvCUqRmgGDIwXWU2wtkDt0XUgfQkp
yAWBGGZgv7DtF1qMBNI3uRW6bz1af7tUK73XucEXM1WKFHCKZMteJpUQhe7zbqe1
u9rsX1G2Xl3hR/JpkdYdXRiq0hXggTDNugbkPmQL+PSOhdpg+roZ3trT6tf9UbOR
IM6JlKSvUT0fS6SqovSPqnj7lL3lnOVGYVWVudMVMUwEPtHUqNQag4JvI3ujobFx
CnuJSqGmhvtM+ia3+TMZJM2efGHlh5c440X3krjOARf9OYn/pmsi/UmxKAyKKTY1
Uufm0DCFH7vdi6Gj337CpUxRQGkQFtIbo3vyeIy/stztIYLVnEsSgjFqn164LQi+
cB/zeSETNeTNBUaE4uU7uyblYwM+dhi9rGK5Ja+Xy4Dg9/L65CMBGvlVC+omi5dl
3blKwS8jY2U48tZl05BqR6LSFKknOHMDOXJ6GDAbF0KfERuXZIcJNj9u6CuNMcn2
8hF0XTYjc+yb3NJ8ERN99A==
`pragma protect end_protected
