// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
WvDtbS4TErX6pPnOr7eC3Wdh2gBKbqxrXauEciHuMjSyWzDRVlBQ4xc0LoeHLqkkvBXs8YghMlZP
1Vz9O+32DXdtQRio+0L6KDeUEuNP9DkyXm0Bb6PsE5wgZZCGo0MeAgiURGV/cMZFAETOcIQB+CgY
G3Q5If3KN+hzHrokxf+8QFiURZmaCelywmBizZwvkBcE1l1taqJ72fCmntylo51vgmtnjT95qLbr
gAYT7YSBLmbkBcBpCnRbRAhUuttYeibOsJyQq+Eoytk781Q74684zlfbxpcuCM1CWaKde7Ye06i9
VYTaKsPBmgPxasnAT7SfIFt2+7cR/sq77JU6Ng==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
kAlC2k6odW1L0/QrwfHqHqPGHj/A9DQFhJfXkZPQkv9AP0UlVetvWIR2WYeWlK1C84Ll+wt3CX68
dv2SBoagOAyGxCuSvUeWqCxQu2BcDxOwH3xDbcOMXWOyOQV9G8gMWw1uFM1qT0CnpNJiD9S9WOlm
T+Q8oE3xqvsVZFlsIr50bVug0VNOYKhYjp504KW7T9e5UBW2NcyBDk7OnUfunadQomf3f3uoUkjL
NcxhJ7pnpAu9SlO/4KgIhB2FPDuqRorPdfWI5jZEeX4fBNBvFIupXTGY/Tkx/Dn8wRsT0cIsNYNE
BQRn07HLR+MvwEEVJGFSKCJg1Zehjp5bdwE378WsN1gkPjyOYWlLMpV+mzvoqi0eGev+/eRgXrvu
1K1c4HGOISibic5Ji95qBSFGgCGs0Q3xeEK5QUI7fJBzZ9vJHQHdIP8ve4DSCX6cNrakTjSVRFl0
d6/7GMIrnu0/4VnzASb2F+rNTXF2oAXa6jOlisxkFdQJHylqf06V7hjh8bQlCdEr+2TWfnEK+4zC
q+sBSfWi2R/SuR4zxnOLgYcfIoIQp6+51ZPFN6wnXBJwo9rN+hFgqf20Z5Ew2Egbwb5Zw4OkWlKW
ZgPNps2eUyvYknJzNgv/pCkXNrtcJxAwSqlassPubThOInIjkSmzdkn0tZmUDavSM5An2y35XBUI
AGIvs9e7SDguZ41AnUepZ2I4qWELSegbrPxJ2nBUlcEiTI9wLFJdzD1NMu3d3TZ3zgQYcklds8dX
/j9Sxu2WtlzTXntPKTVNjqlp99uEfZFiwlpTAXKGdMSX4NBdCSg+Vb4ycG9ymJwwReI5zZYudvkh
WDA4c+UY9MWq+dfn62WMuJMee4SbSjlCLl2Edwkr+QJXakkoZwrJFWjUd9AbT2lKq1M5eLQgogAJ
vr+5zYwr+jDhjxnCOsqm/JFs9OQNp3fXsNoaZBNJ/njbRPxUeuQUO0O5lueN2xwttZEOupuUQmBF
cAo/rAlV1F2SJZ6EGEu6Jh9BSJ04LhXq4l/ZPOEs0NVLGCBM75Sp5sChjTX5UC1Q/Lf7/d9KSIc8
i3H7bvmySV3HZuEAEApIQLS0LYL38Rcv1wpkO2Jknixkn6GKiOXBnW7FckXWqNfGqCyIk00WHFNm
pnvqf+sDFaxn4XmNOdhy19diznxfd4OL+q3SyoK6GVlbDx1x0I9Svwo2YLlReAY7JpUNsv2+k0H0
LY+ky1gF7JX/DcVWQd7hVPLir/Y61Ru1J+0y3iZM5x2fIsGpSG7p6QtJzp3GLJ6RiTDQg0SAmaRh
TmzsUy4vQeq/qYo5QTpheSRYuOc5mh0KiFDYzhL0YNJz3Ia9SZg8B2GJm7e9/oOsONQksf0IhDwG
nNP1pJpiiD/YTcio7FLrY+N8JtNU0CLPejJ66befro0n62MUPD/VIuHTnC8KFzqW8JLPcxf0lcBP
p48C4xzBx+zKP+R1cBItnBTVnogxC7Gj7RxKr/JdG/y/OdjvDT0LylMQEre6raCNVvOlb4PV/P0g
/vYrTL/65VeVC+sHVs7ZTQSelN6uloka2B7px1C7gxchWx+vJYkll0vecPAeMV94mupYLkdu3YEt
fPfd4CQZJHG73A2O0RehRYMtQaWbRLgq4B5euk0ZvW1B+cGvwpX+tTIae8SNwuDsH9IUDnYvqCC4
bp7Vn9HruXTTFTXB+WM/zgnRJdcsirROHxLSrexRlWgaCgdBonIyqwpw5Uo7xLcBg2XknHoRFmvz
77zLdmBQP7ca0Trp5+jjTGx6pXEEOo6OO/BqGgKVCRVcD4NRFegy1652I2PrmggULdTy/Y0zYDew
wBTRrI/dLwlMeUToyYzBD1+498o7wjtoIRfDYzqmaEMjlIs13gesZ6lVqjtnTZSKRV9MxulrpOcL
MoqpjkOYr0i6ckZMxB/V13VTMjOXLFsFKRaBBVwxJ+W0w2XxC2RcpQ/lXnRiIQdJR0R6woFUgERu
TrLIt1BE1YPa10HSJw7+tzfNz+kUm8sKtHU0Z/HFAT25czJjQS+1apRYQtdxVjz+gc6kLkVoLhhV
6XsA/bljcwJgChHfdCBksdrfTaWZkO3ZP3TO/LlPbgTeruVqFwzEt6DKu6b64D2PG+kmyhAAwRt4
Vr3q/+gWoeCOpl77InRv4dL+3J97Shpvkuo/X9tErAfEZo658GfNak7Z34mid3JVs/IM+orTuNTb
onkFzxjycABN38GEIchCXrC6K0I+0yle7zUwMoc27kAPSqn5ytuZ7Q/3s2eVup0MvfwVoVh7tsPU
+xY5sUYhXUzOnWwB1hcFGbuSQ0kLBAIHPEwv/HPoaEW/A1UcLKvSsUGCJXj1PHvp/6pIcgvtnyCT
LhVc2kRRV9SRqfD/JC2GzZ5Wy80my5k3q3ra3hStCKRzNvQ8dHcMPRngb+oaZszKaUmp4vvGhDOJ
N4O0mc3yQAAaJbR1WDIWmXMCCP66sZsT8Vm01EiSqdmEp1Rr0VTZ2LPpnZFxqvoBv6SMU6/UFIna
1RmcA/NhLuWQs29Hlrb9QwBZZqrdAO3W+rVZG2X6apCazWtUQO+HmQTd7SQCa8Q8fqoJ6tudpifG
8zKnJkwggyE/rVvvq4SReZVQLxgQm7ycNIMyRAuVrSyUnKj+QraXal3wO0OJ8pqajk3J9D1/xrcs
cN6+eF1MsESO9XgtM0AtODBa+c1ZqES4rdj6OtCX6cJ6TC430TACcNSFHf9iQbYCTf2YPQMDNMkW
JOTbMdBwl1jhMxkkMRcoRDHyQaIpXcPwpKeRQNueRZdxNfabklFpp/YMsQ/T47Y4bmursefrjzZb
nYoUtTEluzG39EPi8mrTMTCaBLLlmL1RI7Qiu1BoB2ucH2nd8fsh8pDuo4mVktFvL5idZQxg3KIt
cHzWEB7A5QG4i/myct9zY480+p2OEHM5yOCntOFCkb/wCHGjFgg9GgM7smGgOHKwKqQK3y1j2xUJ
yKVdW2vOpYO0kcz9KsoCSNRyy68H16l0/Cp43tba2uqjNuT6PuFSKTOcf3/0r9HRklxDkIEXwDX8
KFHBeQHGH7iDf9TDcVYAQwe5uFU0xat4bN/bTuBQniCm/OXlz37h+w5YC4CdwiBkvT38OCLpFZFa
0LbVhRaAnVTiew4zYNchh1N0pMqoTyZ28f761xKDpzA90mUWf44hKf1Au/1mQ9UY1/JZycg70ecR
KtW9xBwmrCw3+wz9lNUVjLJFaO3V/G/oz8/7Tw6e9GFSupNfcZ2oG/3v2j/wTG7+wO9D9J3+TJmX
DrNi/izweYzv+OCj6MtIQTQEtYsQdCKHopzKEBZr1M2SxEDkEksxw2USRT40oXBkFbPVVqYqvDlP
eRGJe4/5KCk/UwNxcjhaQMhmp1pXvYwwgP9haO6eQaTDUsElIwbwNddvIdHPSICwyJm7lDkMD6z/
8vHTi4rot0F7SopjBYYumQKdL6XRY+PHi1Ua9Q8wiXmjF0zk4oDHc/C6MM68q5z+0jO6/l2hXmag
UXL0X0UQAEtcGTeYafSfbUtMdOkGYZVgUUYpMQeAAwwlrjQ+Loa6CPmd3OA90QqAgmVFz8aiPpBl
c9R9n/l/jcgD0XNcc0rW5B1zSg1B2M6yz37zetQ67N1sHNXvRl+1NsyvgKtT5o7joWIQz3NLFR+0
xSr6+3V4WTOjUU4+2tscudX1J/hJHbWzhYnx3bNOFxuPdmjU497Jim7xHZ3Vy742d1ULyGjie4mL
BHuG5khFS9SzQu5/B8xIeJPBTyJ4U3AsphC859df6lUO/ZIb13Exjku5YkjIvMyfbDpQ2NsvEhzS
acCbp+dQHiVVhUDL6AUSwAyX15AdQGvAXU6rLhXIBId1dOcRE+lutDriD41nZplPD6K8rjEFw2R7
YUJ0/kRlXv9c7IQqw8NXyBTe33mFxvy8I7SF37z5K0ldnrjvQIrpZz4O47OexQms5Exg6evqekoe
DIxBaNZhGiU5QXePFHIzJ+jF2NBaVws7cGoxBmwEeRbAhn339iPPDIHinbeBDpGD1ML3PNdQ+h3e
EC1QUaO1+bSRMBS6J8MYnKm89O+s6iamLeChxZZ13zMgXDOqY3fWaeTyKYsPE04tkezk0ARj6DZo
G+JxUeXFmzfOMdtY3Ii/Dsd+rlnN1EY3OeddlogSO4kN78UH3rruqzybV81oCBKDY96c7B0p23/U
qP7wq0xN/+uhSSGGdase2y3cPO575ar3RBZOOl1NKX7D8caahXpbSmA+TlXreOyap7rbf0DvqLnA
BGkvCl1Cmy6tRIHJnWR0AM4iwg6eznCNFiH2EssDZyOGOp89nRzpZhSvAemcxGP24FIghh9IO/TI
qXaOu4f1kqbzQDXqolTobR1mueNom+DUf8lnN0nMFukQjLAgOeDxG4vkF1nyWBgL3pwt+yKcDFe8
ptywfmVjidDFJIMwox4UP9wlO0GY95nwIcCVG6QdcFLRbGdh4Kw4BhxPNW30QgViRrk+6Dbtn0Rl
AaNBxWSochMLaWpA6jHKI48nn6dPJzD9YfrkQaT6ktvS/h32Gq4hedt56+edTADQGU7Lhn2ZO5jz
dREOZ4VAwaQ6YnSIVW5ZHuheN65CnCLtj2HgnQXJQx2sMzOWlCGqJyL9rl96mpdRINGi8qvJHHh6
+XXp4o03aMA2lJjwwDpWEx7/Mk4C4buXvWZ3morqD6enhT474OqQrs2wmhEBByecTN5LK7YFgCFu
6cw8zS+4cm2m7Bh7tnqJag7vQw/7moSRRAUE+BKl1wC8EL3CU/Yo3L0ewzb8dDzamLtZi0ZsgWi1
dzDo2ak6qRRWj6cozv/K7ZyXNlBWIJec5oNKNuTHhder0Xxyb4glxYsMX3onAv/me5j19+QuVo/G
90juTySC788sacl9PXSSz5785QKmkUXnp3LEJFGe1XKMLay0zDWlOYrYaMahvN0v8ZU65EOVFl/O
UT5rN5jDoTdWoff/aUJVZd/wbXmGRiA7ZQcp43++6qrFaqTPP/bdTYbjmCdWPyVb4kYD1ktrZDaw
bAMw/y+uSKD08T7yVWIWSDb/vImaHad600HsEVMYX5q+9nmlNkK23L0rrQ8Ff04a/wVX79wFFF49
+8xncWn8aziAqbiWjww8tNVsadbKlvHujkpIHQTCUKhzyjLbp0Kr98dGZj6ueefLT2ksnv3rmKrS
MTJNFxqlFewK0iQ6hwUGIqqdflZBlvA7rZr5noOYPWzCFrwhnGelUg92/tBTDEf+gqNnrAFkbvCg
gEIa99pK8okPsc7jcCK0+X5gpapvH712ihJKOPRh/fZdFNVIzKEtqxZKtVMN+BwqZ90vKAiayhZD
fIGYFILyzLIyKnD4FUfiBqFLe9UhQNDXbdB6OsXQ+Pp+ROX5Md08WzMiVtIPOsEmtNKyoqw4RiRx
GzDDuGwQ10Ci1HAkhyi2s4tqmEXXZirC+DX7wiauK9UEa4AlcZYCQlErCXoXo4+T3lyqBNx9fekO
/B8ZyP8yEd/bN680XZP2PUQsFY2Lol08ZsawS8xsaY3VlUiBqlrJmu4xq06Uz6qhjO+yKNUNHe1P
LjBR7KoLdbIhbve8QK46bjGSql8BPH7NsPhBSL2vDjaAQtkSWbpFyiDjntIgjPji8NbZo8wF2vum
2Bz8jhYsHjaZ1wuAHIcTFAtY+uJK2F1bgC5ZPlpVy9O9eef5iQQZ48LlutfrJnJrZPo63CXvWwT6
mkB1zOx3EarPfI9v+QtYGnYX5F6jIJUSHQ1OLztsNaSGyS1vAtZQKWIABEGSfteMDq3g4GP+nAj3
Efwn0xfVDV8rePdNqLkWZUdTr2CnGe3XKyHd4H4hdB7Qh/lMltENtecvm1x1DD7V5z2ChiWcbeIo
SROH9bV2G5Jtm4rcjE5IYAaDsgyt0ymBIL989kb8iE4925o5PDIOHkiSwV9ofbu0/EdCAyPs8pWZ
flDudX24cpRdH70QkD58GiCkNKN8VZxj2gIY/K01bLsklT93NmiU61koDORbBrEAlMZGTNC91AYv
b/t2c0Yvdp5SdukEb+FpZrlKhN21vncuWNoBMgJ5DY6ZgtmmrJKUKnYH09XHW3eA7YfsENu0day/
HdllPkV3y5UBMfZfb3WskmE6QCI1W/oLbgQlseOJo107fbaaOZhpFlJZ/5As6UBoNq3NwyciWtui
r4qiEKQyiatZi62cVApjTdIaJqgl6Von1XOCetghLD2ycNS6tjnokFnroaUbOl1xYVQdHPtZLMVk
xucQmchWoKHhRt1rRcHfiWOfZey/qF3pjNKYt/Hs91v37zRnlj5F7ipms8Je87L19n4+rSLf+Eds
x8k7hFnnpQ8GXPOZCQq3LhhC9Z0axBF/yRaLzBax+iB386t03KtMX/bn6cyXpldaHl4VGZ12pFdT
7x0iyPDrNwW/QLgVveq3n42gJrOQ9Ud31alJkkutZdGbF/TT+FpvQw60nCrzJP3kKT+brFXAaelV
xpoerDhn06Ha0JW6rtrqzSYKg419DZPqWNnEgCfn7Jplpmm2zwfY0NvrpBIdDbUUsU4oqMKCjOX1
yRpyKcpALi2IChCBU7P7pwcWS1McF7qlwpZetZn6iqTO2vztpFs/TdVo5C6GMANvwRn/5WL+mpFD
OIWRPb43gn37tMJCIw8InxlOKD6QIrPNQsL28YJuanFTGyD4AwpT7Szdwx5EGvc1ggk0XAcvnfiT
VpyWlTWSLjbenHMUl7zJXSoHQldVLFVUfxAaIC5l/mzJ31o/nnDwsAGTQzvXSF16e6qHn2EpdWsX
sEVO3zjQQNcj7pmcXyUmDPKtk8iRS6c/O7eR8zDRsHutdoaWdE3H79ISwcGgUozdqSppjF7dAWV/
2WT9zitLykqp4rPewfnVIuKM/HXHgqGyyLD1+72UOZi8revEnOwZb5BNkOM/FxsJgURxXcO+z5TJ
3Y/TclJfxAP2J5jMW65CXVLRG0B9H+SI0JCjmG7u+tTSzKnBpO9MuBRs4pX3iWPc9aFyWg2y+UDk
mLVLnwenwoUOQs4MsBGpymtVwveto2bhO3ict33/f5bah0zNkl6xzuvPCF0c2xBtMMH4z5G3g/SG
sO9pgrLcYXIoU/HzgBtlUCLgC5/VbIg5I6etV31wQ/ln+AlxbwiLmsw/UugjnJdGMv2VWYaKh3PA
XTby18NhvV+PgilOnhbTYQ+JR6JmgfrOV060dA8CIkFNNaE3Wj+lACDPDE1YXE4C0M9xBTTPujSZ
Sro3KRSqONwype3bq5EL6aEkCGKdxIqKfo3v5DYWAJZCzjDabHkEslhGFSjITeW+7a43QJkdI1/g
MEtqWH0CmSWag9SHyxbsyaK0lDRJl97flZwIMHWELBMHOL/QfFbEUJXGzBCFe1izbppPU6gtyiSn
Ej1Q/6FTlBa/rO/+D4Bc7vdlyzZKnzHRR9WKmnx+OlGI6tOD8/beRJbdmhtAPt7x1CtjdwRLby48
qb+7ZPpUidx7kJZKYaHmUZEFX+FgfqIUJWeVluFVti5ylcfWdBsL4CTDIyhuPpzF6X6GqpbnaBmr
DT/Xuqq9XKbiOGcr+IT3jJmhue2A8NkvDSAOFjEi/UlVwbNW/wKn6CBEtRbiHgFucmaOYrGg6stn
CflKdNp1uIyO48DXz1vvnrBTs9pyrmk3Uu2hZ+NHomEBD+O5wgDaRwYbXcT9vRMlmuQstDEg6gP/
ess+XsN/+zZVgrrDbuvelrv+JYog2SjaTs/3URybr7CWettEgZ6Bxm9ziccRQy1O8n5/iStLNT1L
TU4RvqbqVc8PFStzmGPaC3PdvNkGLrOa+Po6CioiNyY01HWKQQj8xM06qH63TVin5eXCp6BTg5Tp
4HHay97nFCaozPUKrjADHf7uIT5hCnbQZ236/ybiAX3qfm8hjPIQ7PKFvpDfrdURdQ2utGgR1e0K
Udc7BCMqvTQy/QVVrL8kAIM8kl0D+ApolGeGvMXq/QzZH+VzQ4Zltkt9LKM4zQFw596Vj1TlBSBL
gEHCv1c1+alGQjfw8Q9Kw047sLgOP6VuXxrJoeZ62OuyXLjCltRDKsHa1IaohVE4dgKPc3bs2fpb
35wxhH+b9glwtGoTXRvHPc1xdbLrh7sWRAXwM63iOIaSZSugpvjbUl7Bp9TgA/Bwds8qida2kQ3y
YHBAck80sHD3HWHnLMtUPKf1bb75tDhu7kLeLeritWeYYYoaJpNIJZnXSO5YdwRFhYWEY93VT8UN
YdmeYirVoksHSa6Ril2eHKXx6lBZpbU+sQnkOC4RZgusDywJ2TdUA3BaaUP5ZROSMcAle48XTlLM
3/LvDzfPXZ1U+I28xnnSCVT6EILFqVa0tQaMvLZ57Bgxptzjgfn9PWBBzzlxv+QAZ8jfbPe/Rsaz
4RPZRL4Gw2RcPTXpUO0OT1O79yf+B7yDK9M8h8Zhhdll4BDjnS7sENbykzpMefKnsAfSqybyakWc
zdG62TbFLJpSyBowZugbNPlwmev+vH1cVTuynjiPVgvIYGkqqfwzpfB66P5TK42AO5RhYAqEO6R1
6JVXRPf0RAKuP3t7CkwwjFlDy4GXM6PfJGSBuwjaYnEVffdkB47pr5cOrKJqm6n/SAP+2Wwhy3+5
U/7NP0YvJW5WYd3sRVr15iu0VqLqMa1o7nkDyDu5QyE6XyymK4OCt0F9DpyXLBIMbd1Q1QsYX4Yb
j5Tph9l8Ux6dSWMCe9LiIWa/y7UpTt4c7l0kgoaAlm15sUfkuVy90goF/pYaqYTDd7jWJIDtpAqh
lNAnJZvitYTY5Hn3rXqkTOo9jkyMgCVT578eCRcZ32Qz5flLd5yzqgaPmFUj4x5A+0U5SjZcHZMd
visA8j8Prj94rB1tutqCBnBMyRikbRZBLAGyUyB3ssbmiAsH+QXf7vshqeuOSoqH/5J/UwEiUmMm
DLvFpZwbeKSh8uJ2ymRCTasKehnOt0V24QCSVC58lWRl2OKObaI2S92cew5+GJ2E/2JqWp205w1B
H6c0WXeXhbMbG2P2sKsCtPdpjnvT1YRH7Keh9d5GH/xdVPw5S5QbUveKWBj8NlRmBeWz/Usy1uo3
RD+Y0wk2aq4owKigEbDGq+A4OwGaN1vaWRWw5ncA8P6ebexBNaBwmzGgCCwM4iyM2fzI6e+IZRV5
IDmJo6BNIqrdx4NelFZMthu5fch4toFQrE2dNujiM0OLzXxSO5c3gkPwZUaRs8mGPbUkZvPESiZ7
2GTF+WwdX7fTdtGt7Y9ViM1ZqsBpopq41j1K06nZl/Zqd6Th3qrsEqZqh3uP3huLt8jLQDqgVeN2
qk9ElovUNWCxyKkwX/AqKt227P3335jE3FK3IOfs+OIH9SMpe+O/Y0fZew/PVCq1i85jZpO2WP2Y
9XVIPCpPREb/41WIn68LsyCj9pY3GZB3+z0EIeL6zgADa+CPrP6mrf/C+dUyUM7k/FSQ4vz1z+a4
pfx+em4DZfKMdQzkA8/+0/pn26A+uDhYnjxis7EBXzUd3VNB1fQAWuaB/MqU7XzWNt6LfRQt5PF/
z/mvY0tE0TSRGh3E33XXJSf1f4lVgYly2O7ozR05nFF85EWH2B4jUmLVT7r44SDKFs6EYPfs0IZZ
SU3fTuIIrb7+cCVgD1zwdAUvcdU//FpJ31mStd2O8BnG3XXxhr29sYRMagFQF+GDVCU6WnrSzqpg
ecLYHcJBKdBZuIDdroZL1y6pIqigNcavbB/7bvPFZhoFaOrQfVMv0qA=
`pragma protect end_protected
