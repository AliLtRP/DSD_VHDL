// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
p5SKX5RuqhwpYIBdsZH3YIoOk/U5NCL1C59uB9Ga/NPsEKLIN7H7JsKvpY04r7fc
VSTIwxHyJkl+JbYwv/yvoNNqCuGobFf6nd3LClIciZxj5oCwBWoKI1kHJnXdEFjO
uppyssRxLI4evqTo7DYLfO4y2kY4+4an0lj4oLidVRo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3904)
+s1iwiyqiM8S1vsnQQhKEK9cm6vDwL0sugVfAPyoFORmwCVqNBSPnE44h6UF2RIb
Tpu4uxhA31Aa0QU5G4yywU6k05gZjJSoSPxnscJ1/0YHIZIx5JSHA+1RsTUHGokW
WYGKyghO7T8OdGGwe9URLdvuHTCDEUt7d2OHRs01n8BMzNGGHkrRTy9YioJ1feEn
87TZrgyytbHURXft816AV0cfxhYVVLmAByBIMp7A2UDq0GK0YK3upRjVt1K0j1tb
WVqiG8vpOo83rybUKlxXrpXSgq8muZ5mwtNZ7jucpqao8Wa6Ww+cbZx8TmljSHjc
c5WdqW9Nn9BdmOgo7wjDCVbBr0B2UM+AfKMBokq8Id2IenxabJlAbvSZ/Jy4cuuA
BQJx4Yo5REDqKFDeam6B//TzjPH5qmTAGmSPEVr5MWpn6hox29MYI7YDzjr+goiK
dB8NLZNcokirNpkuBZlcOA32rae0TuzXE0tNBazXH6oMRG09GOdi6wrLOVj25M/C
5tUNiVBDMtnLuiQWMsKqGnyRz/lZvzovT6fC9aaJIV6x7VpRdi/IxwXYeTb+nwVz
MOXECezxNG1z4VBrtlQgrJzZMNxgnbPKatV4octOCTP1fwvxSS3YaWdd+xOR8WZu
f1vLIPC5fZ8v0W/gBxmTixj6h973QIFJVOwQfUcLcq9pWMplisb0gbcuGpxBSTV/
QmV69ackbKM+gpQnNu+Q8VtN5rgE5aTeLcmciBB6oBCLG41gxYwgmMueToTxsrm+
PJl0BxjLNLpy/epsoojj523HPNu0EUq8gJRQKMNJs2XvAZBOf/V7M9yS1Krii89t
1Zytvr+hNEAUuMoaQPMJ7GvOHY5zmWOHjbzPjDxIGzDVq7yBDz3YUZ1z+PYhVY9M
Hry+ttm9++b1TySrRkPe0ZCGqwBfAZFWvcmVNBFuNOJSu0gVXYZzeISnycjvpCb7
rc2poINW9TzYWaVMvLNhyzjQKgJAWLiHwHZwrmQsmMRpGvJrCRDw77tdW6SyYX2l
6fh3uOT5BpsgIX22GTyRjhVDCdVfypz6m7BtfMW1hsR9cPrAHwJJu1GUyGwOnLWd
c6J7aydODo2HqGrrDTV5YuhM102HHl9TRpoXoHgwKck7uAhIOKyBDyqnytJAJjb/
TOXo4osR4i+uWkkKwt3eo3tRL0KP7hpbFW6MC1etQ3Oi2c+DiVn9CSR5ipC832hm
PE25AR1naZH2kg8Z22aYBB3FjZcVqX5lPk19AeG8m2vSR6k+mlFWOZ+3VsBGaYN3
hjp3+yU6tbC/An7qm/eb0GF32kHiALbUAQXX1t/mzr+p+cxpjHW4cfVAjLst8Q/4
IHu7eatA82gGneHjrbPPH4zp8euACIeZMrf+E1tkQu5T8FkG+qG5W9KmYibCA3YU
Js6j6V7xgyGvvQCUYXYrKUh//yURLYtyTDt919lsPUE3gsYL0POhb2Nm9toChT3Y
bdFjO+DOMgSKUPBDJT8A8Y2q9cFB52+u8JnCg70MXBz5hrAvwT+/Ok4IQkx2qkem
/KeOC8KV2GSYEis/l/lb2jLwIzSdXTeQ36WvXOscGD7+RfOQXrv6e/TmMGqcxilE
fLaVDDqL+6spfwcF0WjTFMdWdD+gWQLswhOKq9MgJmWlrniH8Zzy4Ld6NxyFQ1Nr
gWkNSnOWfolqGL1HJfgSbXHehHO+8eCAutTysymyuxECeozcO7NmQkph5wo227lk
QaXjBOoz3pfEg+6b8fLWVPu1EYhwBtHnJQMACqWjKBYWwf4ozMrRzpB+6JnCLkrv
PX53sVcVRtPVU+/F6lNoEizE7B9JBg35yUHTd4iOqkriiCqGMYYHSWnqbKgf30qg
e6QMOxGchlvE0e2kgTpn/SL6f6X52OS/5wdgS45c87FJaPfk1JvPTrH6TpQB4Pi8
Vdghmx+ctBGL5er8AeLi7uT0bPPBzHqM8ctxedtLdWZ8gh39LBCQHmKbOzRxaNNb
xETrdcS1xrOcXVJ/W+wbb4uGMDf0vjbQHH2hx1FicLhg99swueDdd6ZCERZ6HTSo
jpXjx0bdwCTTdvjzk3s7deqf3xGGDC8swdnUZhSkZpEwfPYrqNJLKgBUqgEuBuUn
Wd3REPWCl2ogkncaiQaFfZTVw36nNFkFsXSnP1W5fQZiqgk93zJGmowKXdz2sOkx
Ye+NmM6EB8rS8y8KpRRDOUYEuONkW4PIeOMH2UWZwBequjRzAbGcyukqe5OB/E4J
KI1ASex1VzWQCVdRtgyb6WjQnJ0qIXpSk51VFL2/GDIt2qE5Sqqlik28o8ISe9or
zWlEKZhyrAM8RndwkrVYNnkA1ZwPVvOrVPKhE078QthB0iZt1ZhIB/FcPTN7Jfnk
NYzLVow+tLJhhuWIWZniFcYX72bQ8gTl2pgILHVuXI02bAjQZ1+IRhtzCyqWV9YH
1VfMPAuJIbl135wIwGEWFpfE+yMLTYC/GH3mykdKtSCMz35+RSQNwSXfBA9s0eD4
Wz2zomKuie0JeXBGdcm78XZxJkEgDw1JRZaKR9OAMl0kebgz94DU8Dgv/aMBjI9O
jFViW8SVPTZGVSvXtyIwWBtsxgREvn7arXFY2tSnf8T9lJE7nxFtz+pgT4C6cCSY
5dpUiclbu0VlWG6LNjRLfhRn59N1rZWQSMARAc9/btt7S2ReRxsJ7Hwt1UkGUdHN
DaRwscrSodgaSVVJFZqwXygJKsmtQU0Aluk9cv+5IX7HzSFnHHzc/1I+xjJcTlrz
JS6rF2uGw2OvhCIZeblmZPRGy3k4xZZF9nBHNh2eHUddR28bwTRhevnWkmjCl73y
4NVndLbuzloyhcxZZCZP3BGGjHMMIyjjpDgxCoXZe8M4dV+zuKSCbWSFYg/I1kJ8
EJ9wO4AlVlffOiWImS8mzOZKytNz726eHIrlvEcow7o3YMxxDkM/QFeiFQDqMbxp
NdsiXaU19RvTHmiIW+Zc8xaDTGI0KKuyiP39kndiHY8hrkhFg2HXVUvgw4NtVVC5
qHwfzUuDsR/v7HUHc57hKk35khs5OwdObD/fkSq4IMudbEm1B+IntsiQWRpR14wn
ZR7WUmE5FOqUrGuon7REB9KqHZhxLGz9km0KexSTbr+prZo9fxYZeSH+rdhqd9jN
s460CppAjcYhrQeW9TotUhfsLWySbdy7PoLVqTD6GdWEJm01wGRz39jF88rbypFN
ApMrKAQ9Fs/du5dsudZMbuMmqgm++OHeIfy/9vEqig6RYAwm4m5X0hC1EaCLgaX+
t1APWzA6e4aDK/nxo6eN/4LWgEgd4PBtzXRIhUDENCk3okbwrV2fSETg04AopOVk
0FQViT4owpqBRaarsvfSl66ylrEEP8sL4NA9onoEtJOf0kWeEOpLmb8W9IU82ksB
tNRyZ05feJgrwyqLLoLAECZJI25P3qMWqFu2yrkPmYROsUncb+MyXuKZK9dQItMK
sc61vbBdTdUVP0SsckvP1Bx3bGdmllCNgrTZB2x7FWxojJKtOENie0WPJkbyqmjp
nekBhQek3NmjJhx0GpeuX++4+IDu/x+K7Ah1s02DBw37qD/EfCGDORoKzoHlJioZ
GlIE+Qql87L6hAIKVTdvT0+20Lv1Bt4jlwHq+A//M2gtw9bNZrrtRXd3kHUgRmrh
dkD7UCqgLNdGrOdFP/UBCnx7C6lAgQZNE3HMNCfv0JfHrDXEmp5BkClo9Gqdigt7
QzfoOUzHeeOPz2DoS6ABeP6mpfWUmjyI2J5dlR9HODpcrCRgmpXZKEhS0l1VpC97
ZP/XQVmwIt2/0uzV5WMRRBakVB4jhIi90iYcqPsuBy8+iq/CQINrA7yw615WGfJf
J2qLxaNJffs/qaC3E90PlumOLBuXMXSN4klwxGUxyQLqW5V69+FOrC7Vh87QJ1vN
Opjmx1QtMkwzmbp/ig/7ygrsb5JCHECOwXHZEGnutHKcoVrV7pJ+JJI9ky1/rB8z
kzvlRZb8FSeq08Xd6XNhXSmnH0LaNMDNjt/j5doO3ERf/J50GecFEBlwstoNgL9t
QP67LLrw15O0ANCFfT+18EQyzdGbmFT0hJOMpUFETqDjTlyB1BT0Jp5Lwag6K0U0
bIejd53X6M9WFdcbvKIGDJSbWVMkVEXzS/9+tq117ceL0AtwDlJnYkz2Xu/0eZpb
H4hTlW6/ezkmHIc0jGfortTYO1rUgpIB70Q9/a0D/UAvbLBkSDYSz+4am3OddpTF
jLUOuYJTX8i1QZO1pRlo+XzZ7cWeU3jKXzxWvthFl7bHc1nCnIhvLVwPVOqzSIVy
wR3M5SqW8FtaFtwNIrVa0Wen50ImHqBtetkfY59ClGRiDYs8FIPG2KuEa+UvhC4a
cisCqr26gSeSI9qH30rQznKDbosw4ExOqWVxiBkkEPk59O216Ub9FsejTwPis1x8
ZmbCsrN94pBTJHp7WbiEqwG8tBplJVAy1PbvLOyIEnqhiA+tMadvUePL9TSI73JI
9BZfavls9xASf4DOCCOMVZM94OWnuspOYmaBzbbs43ZoOx/OYeyWMjY0+bz6J04k
ZeCuJY1fogDMAdka5kMDJuXIKv4bt39eREzAw0OrxfIdTznuDzoBCDqETJns/1B+
WDqjKjAU+ZEKjc0MKkqTP8DGioNJaEOELL3IU9VYa7nsHzaYSjEG8WoH0v30Jsf7
OBRpjnw9xkX34vaOuDWO1VT1wlm/hWqBM223utE3tzJr4LFzNI/8xLYLKlG/tzPX
WujH/xmVai8APsKGLCV/3l4Z9+kYQAVe5EiY1d/iyPLlMgmZgpWFUzBZLX8MCoza
OCcKv8k0cNolvCIfM+I16ig++Mehq5h2eHYRQKJzVyJ3NG3wvlg4PwSLB1eOZCEP
KLKzFjyRqtlP8b7kCq6F0sVKq6godVn+WDbH2gszbYy8JZVGc3ACFxRrqEAIokB7
Nqcdjn2HEs8mgYinK7vbvj03A+X7Qw3yXpOzxg6jSgAKKr70iR4+raYMzGkfD6Zz
EJ7BJ6AnKSpIHRDNKrCQ5AWwT5A+QOwuunoDKp2oiPGe0uD+apG//eRgbcahO/08
29NBJQqakEQq9vdJP99GFC2u/65RfXzsN5YDDhAdFHl55EaAJyKdmByrxE3R7EXw
PkS84iL1NT640XA2DJsgtcYkJdXpUhKHXe9MmlnpxEUkKV2/5y2KB8QdfJmhtpfJ
RaBXt6U18kod+frASdcFXQ==
`pragma protect end_protected
