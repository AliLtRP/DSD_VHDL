// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Xf426+XLGuObwXe6SqMvS6srmqoBc1wfP2G8ONn+8z/UnuFvrbDBSN8544A5sP/B
DNsZedRYKJnBNlAquG0VOoex4FoS1a+aDxZDLfQYFfdJAsyWFysl6YfLGRNNRiFT
8N2Gy1O3GzOZQQ2+fqi56PvZ43hk/rHsFFAqqpXkMO4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7248)
0EExieti7dnzF21GYn3Dm5cWrzDESyAdoNYOSRUz2xAkcoHNlWcC7ZNC0YK+Fh2Z
y9DKN93BdR7a0RyKlxxbemEcvkMTz1Q4njMZ8zNBS69fcJaWhvpaPRCIPvacKK/4
tpUNAD7pkiC+G4D/ASQGGL/rWQW0+HFfejKuT5qvyThCprDCj2H9i+lBOJ1Y50cw
Gcqvs2v9MpyImWzUubKS83JF24zTF+7YVKpKiINvHa0CMfVAgjPytFf/h/AVqLT7
U0ehn5nJoJdiqNSoSt+EBylHXNbVN8TiTnDjjTHfJ5f0slCuWeWiZdaoSzXEFqPN
wUXVFpDTZF0aPbKbY1DmrASk0okl0xDyHe4k298l3HZwbDXzltVFCELT+ouziVTu
9Y3wPlNwst6QMIgoEk/cTi3qWMM7icZmueEATCc/P71gSUtOaTC66tzgu60ctORR
598HeIXxlax07EbJVpcCZB0TsNYpvT9T4Lb7JnUVaLWoYVT482DSzsZn3MEbU0Qc
jWsbC6b3fDeECL9b9h/RWuqLutZ8RQSE5wZJFov+lBx5NicdZ6aqWYnY9W7QFeN+
7VgRXYr2gFX3aqgMwslbPzjwy5EKRxXkB9qKbUeyzNKE+B1D2Xv465LvV8kaZkwy
bTVyhDTcngf+B6kIrrGp6BbmfDDHraenS4i5ZN8GSkzcYdJ5BF7gy+pNecyOQxCK
ckmHqS7R7HaVtWzaJBAQJN20CP6OkksDdF+8p8Vt8/1XDaXs2Y5OB5mUt4OUDuEy
KrzvGfQC24Zcsx2PXJy3X39KERejRDFMItGiSv/9d7iF3IwNrG/NjlagMGtD9v2w
J6KNWr8RvCt5t95q0w3Lb99KUa36Wo/d4b4jaM+R9oKCH7t/ZCNhjNhWeMI29b0I
WNxQiPzg05++BTor7QGlTKnznayJvZYT897KW9BPox130PZNiuz6Anz8vqhw4ICe
qcv/3OzK/bLcglayf67V948SuhW6kDaFRa4xGR5YrEU0s+mv5l7ec2P8QoQIVcVJ
ncsvOFOcheCPd7X3tb3smgJcGu61EZt7zGFlS50TEAXhsZqU91xHWdiQzoK4StHM
IqgQsvHqEqW/Wlq/kfItH2ZEZXX2Bn44mz2z5R6sQRWt0dgEdeqoiClKB+Bz4SAv
KRbT/3lfnE3+wDM99RCO39wcC2cOd6b81vuFL5333CsrLcJ9roQKMiFgGCoslMnH
BCUfFyIBmunXSjzbsJ6qSi2zFDWvNiRSwRq2MvjR6NFTFa7Z0+uyP0WP8lY1OhqM
VUux3xIuOL7NpIasWZ5vB5/TPKPi/BdXDeouERTDW4iH97bOYEpjyBDS6jz1wHdt
mg+pO9ufROE4fS22TWWgWTHXJTFyKzqEywM1bUGQTqwcepWhRyhHigCFrhgpkOuv
lTsMc1sf6zpMe78atBPODTp/2KRR4tuRLUpOEyh27ZckHUc9rLvS3iE6UJdvBJu/
4ZY8t8NroI7GB4kgdBZ72awejn34TcB63As0oCYaq7947BE4gCaIoxh20xqtOSZv
Iu04VKftCCZhj1dB2gD96AUfoEPkGUZfFG/p3LWu/7IfztYt/kMRqrjrCPXLC+dD
Ilb5rJ526cUNY62CLYJ/8y64dRaEIVsCI3VYlets77jvq4jB5TQ1emB2cVaU8wIi
Ogbkfwn+ByTKo1lRoHeDXhDP7HQu8QRInhX+mdGGKj1NVYNtmk/ds394M8UsIDvI
C8NFQb24wirgTOLCelVNvAlc9tZpRPnaLwfsKTT67Rd4axNVZKUMst61oWyprN1M
7mzq9orAxyty3d3z3DWCT38FW57a2h9yjCfECzgCTkEXF49QSLCxPkYYi6g0ywnq
w+/MUOmevH4UvQuWbkvkP6OuZqcEhBx+NkChcGGYLufBylc4G9DcrJSt6T9GHNJt
2uajj6ktKyF49X3Qht+JJ47e9Do5pyC6SIdUBNjwkv0b/WVllP7gJx63Pvow4Hku
ZhMZkwmIziZ7wFwa4hmI12vKNwEx2ImtlHm7unmmjjS3hfsEklSkpjfwq5ZXAefE
52JjLOapF0CfDjT8oLgPQRqzbCOoerfqZ773Nz/PgbWX0rUEiZ1OyfU1g9c8Wc16
atmTCZ3N1KD88bDQqXKQvlNLO/e/j5nN96HMJSz82spscyefCkwWOLfCubXjc3V/
8WYA7Oq2godSKoC2d/6ojSAb3C6y3GCXBk1Djx8oAYsom3ei/VDyo1RgmoSrSAr5
ioEd6X0YM6A0sIdLbvcRPec8QQEZGWtur3OvQ3XdmmJeOsEwegYn/TeBZ0ctvPvT
WKDnjHrifC5yzh0Bfq83uQKrAEVKmhC+CjdexfpqWjEW9ZZWkpvuhbRPSAWkKfBj
OWB4cw/PTbL1j4HqNWfncl904xob+j1B8043ksRo7f8mv0lwVLtWfXQdlvyC6TmU
3KTjqmo4A9eGCbhTyi9G4zoZm3vXGNjCElqJ3H49/r1F0POALWaWP+K/hJttaLCm
8O2oNeldAl4uzTbQLiKRnzw2BjqKNNTiN1g7hgUrL+LWwHsHpA1HW70ig0MYkJ2/
FBBuZ7D925drY49ksWikkxA2LSmB5oC9h++1VmvvTAhYQiAS8ELTuGIsLbnwWGKZ
oekTF7eykiMuw7ViIJcMybhqDDXOGm06ePOHB+kbSBuOnYHR8VijvXnBx30niX91
mhSoAi1ITjcIf77AfPckPlDFCdFBtlumqj3I5jKrfGzA3ML+dW84H4fE3IJSrYnq
p3CXY+ZVHZk2QTt6ObVsXY6nPvlwlNO+ZiXfepE2nigD5J9MN2/pm4iPlnNsci2c
FdmEbNqz1Q5HThvZIXFNbZu71jGdg4tQ/p5HsBuClWBPkl5fIbAlk1dsxPuvtm+K
/WmXTuavkSA2oaRWjPdTijoLA80zULNUTQu3wiKAPR3pp6q6KgoADQ5q6bqICTsE
bGEjVns81TXPwuorNaz9o0GiuTyorTsVllDHAj1K5qIYvX5k1PIWdcPhYupu7Q0y
S9609WW3h59lELu9k04bLjGE6UHLsuiA3ipSI5Ea8IAkllgy59zgyjVlNJBWi/QS
ngsU5vV9WITQkDWU4HNrfOicJJSf/dcZ+5u+adbTMY7t9WMRGiejF5Nb9PJeQzv+
uzZTlleaDfmrBBx7wuTavjjbmrSzR69JSNadfeIKFm1JcGPjGo9AttonJxxz9fGW
CKKGfTarEA6ne1ny8rxUsJWy5OekOSg/HNH1RoBptBS6hrTODWjMnLOsf7fLDnf2
HeYjiintmloyDO4PXFtWkwBEyRI6ot1+UkovCLgsreEeoSOBpqyO9gg72nKn1XYr
z09UoUSbdcYKdxcMyZyKbHh+3CxhDkYMAbU7xoADCLbAHDxfvMwA+0IBl08w+VL/
j373snfFIKdoIaPJIcYmHor9fCY2iP4JE6ifA8L0hvTxBV61rEqN+W4jYlroSz57
8gIN5IoL4GZmL5owtUVLEm+Q3+EWC6jlI7+VyKsnnMLuoqllLUZ8zCmjayq6WE7u
DJuuID6dBs3Jdj/ufGeeJjlaGpfpVbUHEs4KvrGZ/ATddQ74hG354tufsZA1cDIV
f7TZWbRI8kfIO25gLC6zEwkg+P19Iy9AOLXX0Ck1ifthLKHPkiWHwrIe/xJuB5wK
9wZiSqkcEJxSpT695HCTB7cmBZE3PJJPqI+6s3vjOvMA+0hW1duCRCsM88jUDG3d
akiFUN0tnTtLyqePw+YZSRzFK/kFUJHYnegD7+IhKvMfVvO6LqGyI+4nt+lXHxqs
6hgmibEG4dg1kX3nsb/vxb3EJ2Kx3Lw2arOTU7IqnAIhknJI7HzT+wzEcT3E0JHZ
T6MGMu2ZZDX19zgcJ8KB8KQNdqIYux3WpmjV54JKWIcM0A9ObVBQoCBC4ePiWhCB
1wc5NSEMu/CW0zEL8C8qhQtPSYt50REr1gNX61nerWePCrRsRfenkRQqbFaYIaCO
IgqX/m6cXP93TOKahCXt1Zxsknt1wbfGlyC/5rO8u7xKs9x/Wd9aX0li7bX35AVP
7/Do1MHKn9biKEFSdEP0ZGrg4XkzOJxPG3F+Taw8HUSTUPMv0EqktkYz2wxg0j+y
7Y0pUS974WTe7mUNcQu8oRU9VhIgot1f7LzitjLaEqqNjyB/nHn7TzDVtaQMCRqd
GQhYYiK8KzaEn/3GAn9Do+pSfCBT8L9tMPzmUBXd/8eEVFc/xMeDXiSF5ybiuapa
lfG39MsuzoB/rQXEpK2D/8Mr+hQm7htIPUhn4+QX0gpfdkimwLjFGRgjLj19BCxE
9Kv0J/2db3WFZADnF0G2ERmJ1Uj90DAf3aB8Ex94v8OHQc4ZIW/R4xZXTDejoATr
AwM9vmzU6ooRlCOrliPiqHAJXqsPwkzpVS1e1RIaxNvjO9P5IKAUwTgqdg177OAd
bIJyaXAZi+Hc9VV4SiOzClu3t6KkBvw2X2hwbnkG3ahJCzC9Q2idd/VAwMTOjVK0
tVppwcbOp07LuAGwWzbbjE6ZdgOOW6q0ebBZW54hgShf/Kf+V3G/PL36jnpvXTFw
zJrhxroLTz1CGzETMVQ4IgpsvBdatnU6NjZMCvRITXJtbQHi2GN9d6amCtBq4LjJ
DbZmDkXysbDS5OtgqKPpiFUw4Y7xJkQ3L99ZbIAIaNWz8JgMoh1erPnBbVSN1EIS
Wt7JIC7ZKm/etzcEbYupnWW9vaPFhr8p3Ev+qNxlRopx6p0t963IODnBa36DIqCk
pwUAQdYLXIRm9dAU7PRETn6AFy/PrTeL78pSGQWs7IljuOI8XqkUezxo8y0N4prr
O3Z07gN67328iHMW7YfyzHYEEIso1XURdoFSHgg62SClkdO2rQ/HVf8+LCRrvU67
RSnuqlAK9YVqGuF9JviJ68+osKprgIhTm3vg5MC2nusFvhhFm31DuSoN7GCX8mNs
8DuR0SZCs3RH3jLTaRE8swyn1VAliqEvdoE6tmLFORUW00HGzIcqeUytTwjbKmQp
Fi7l/tTJKYsF1SSyzozumcHvyB9r8jex9nni0NMzOfoR9zuvvJYhKV/WNQ6cguAV
yF7Rk5M24Of2sDJDVvX1UCej/ux9nt+56K4KuPN/LSQgqevGzU6MUNU9yAYw05rW
GWbDPt2/sMQY/20wDxk6tzvh7ku3t8o9BbgdB16jkhKzA0ILme9e+Nkqku/o2ILn
q/XSfaMiQcFFEVrj2RvQxlxirdQrJBV4sg73bLdduOI7Qn9JW1HIOj/nfM6srH8H
vmaDlh26ka3Z2/zC5xnplfOfm/QYnIM2EKD+beKB+84Syqcw5PRojLN2JQVM+JRP
c7iUH1dlbGU78CmtKIACsdVe1kmXIraogLZfqe0Exm03nxTVIR6OirS1ceC/h9UN
0Ovu6/6rtRze4SxnUra0/EbpeUHy8lWjKlpVErxgvi9At3I3yP5Nzw/dF6Y23CtC
lH6D7B1Uyk1aCx/Wy/SIa3l34GbTBTlh4fQCwNBUOHTDAGUW/oA0IY4TN8DTuGH8
lh29BF9V0BC3VUG8RPfCHYerpugQtKOiIgqH3+ZhIOSUHhdtEVrOiZUGU+VnAezr
zJhZ9NZ+20Q61NetpxDM+yVhh48TY2CzaOCxiVZ+w/U6ZdIoE6WJARXi/+0U2Y0y
+ZGfkeVaoqWrXzBjg3jJtVTMW3xNuF08ERa88uoSBbUYCkG8iaD9DG2XEIJtF1kz
5PES1s51mFqbMdmBtUck65uJqf25ps+2sQzxLG0Xy26MXqxq3XSaDeKhmOUTaJ6k
0x/shNu/zeFyRVKEV4wxS+hD+JQ8IWGu5FqdLgxfTPnOLJzFeLYiHUQAdYVsycrE
URznJfuzbQ8JSomfE5WG/oFX2oYepJ/AOYVRpD8A8PtgQl5JbR+t7bkoA8ZgHePM
PSC42GbpTs9FR1+gTJHBL5+UxsPHZTa52IAMZs0kCgN08yCfNT6CTdaO7daz84+a
QFR4jeb98RAy4fP0tG6fSQrLm3kcfx+Nd/bVpJdppr4fH6yQ/mI35XJ/CodNe7S+
5VJSmET0dzqf5nCtE4wcLxB7LNa6U1WipnRaq2bzOjjeT52A8+QXnFPsebLISqEz
ks3dRrrsOPItBNkRj8vgjnlhSjZNIj/PYO17GzhNnzclibtLAufSgEc9Z3cqFrDa
KMeKOojh/jvOzWg7vqfTvrWXwSPVVoQgOIyjjaz/8CxBJuUqDTUR0AfOlNKezw4P
ODAlLOYCJ9WmYGCHBIWreWwJXkLqbkv6YLP4WCDMXpRlJv33sYn+WyDdxNjCGqJx
VF1RUuAs9OHeVZFs4se3n6wj2hQPg4iXRQAnRleyLVnQiAqrEkoMPiJTG9/aZsvz
O0cveUgYAqlD0x9L8vSIwONkVliK6TwuALlqy5UwM8JJBsvxV3pusm2JkLPsKg3P
uDCo5H5tlcEBdO6BaquR5u5ZK13txZJB+KRNYwssmKpa7VtQAdKbwtxxM45Qathd
lGz8K9rbuDXCuuNpxuM/pVmWUUZuWXuznlNZi0hSJIHuVnO1x6ftZR+2sWlnhXYW
TLm8ZiB90f2knuDpCItrxMPlproaEAnLz62fgZG4GeXPPagQydHOS+45QTkZxEyt
cwiUJjcjkZUMCun6MujV3ppFoUvPGeiMC6FwPGHrG3X/8+w664Yxv3hzPfwNTCh/
cewSMiLH5NaqJDy6lczMER07olL0eOhTKOUwXqmHj0j4O+5OqEtMPtQtLeNqJ9R2
MeuHC1AWO2C6unitQISYByv4L0FtuE/y/Aaa3Db5J2rHM7BOQ8Mnu9s14sUqP8u3
IGHVOTt5vWMrk7iaH7LABg92GsXqH8zD8nZfK1ZzTVBz4aelZAqjih8AMcSknZG7
2SiwJMcwiw3ZeR0SdJZaJ78S+KeBO4p+P/mrXJkR1zXsGzkUrjYylb/hwGFQOzwx
0eEOZlHLvxJpLRR8KyZpTfJtgMq9RFlkmYoAOrl/uICV9FaOEwbtzNsqlUBnVo4t
N4szILjbKkXuZ2meLR7ZWTdOD2rxYZKjn3EhM9SU56YnUAvaM2GbhVehL/sjmIgs
xw9adc5dWVKIMWt/Evf7sWzmxcJiVH8+s9VTKx4na3P8ma/QX97GPZo3eBJvBdmD
PW4nrUR5CtVQNtFBTIXlUz8w3DIw5UPbKC3uCuzh1tWXOcfLgaClhaCDZ6HwbNxl
wVNyS9QmnSOQIySUs/il21XE4DbPgImDV29jwRKq78sORdfetcP0jeLXOyzNJJRt
+iGJRn1uqh33qTn0VOm1xyqczPjyD5DxcCBngat4lsfxjzny15clqwXAuAOQ1gd6
yWoU0ZKDm5pC5UhfJzM5uhjsZFA/y9nzl1LfPwLq2fY3eIs6/jg+1QIEqXqMKPKZ
WYWBFsSmnbqyzxnEcbdInhKzJHx7Zxo0oYth7T2OwA+IwCNzK94AR51qjUvQT9y/
lSRpqxZpihNEJfbbg4DSfeXEQ1JPmaeYx9ns1J9tTvIqY4Kqd5gBz8k5lB6VRkZ2
vUCSAMn6mKQX6ePtSjjd0Y6IXxd5PiHj6o8JwYhCQ/YRuR62YW79keCYpKY0G8b1
OsK3wMcqHXHRelWB675gzu9bFPeA9JLnZ59V60zrlZBiMMvveipEXAF4iYFr9EmL
KP677QxTg0FdYdh8CR5O6b8c+c3y21IiKcMDxMr7vMRzIkuJ+bGh9HpAAJf5QbUD
DVsDfg562rHLK95EH/XDimRfXklEmPCfXY6VdPmYyBYgyAa8NOR69QlNBEg21LrW
ucltdyAj30iyOYtU8F7GiiAEWGJfoszYtzNnHgNt4BcvVmYUHTFdSxhmx0SfVJod
uGJIQWFgDXUF/ntIxmehtz89NIE7ctGgDH38jmeX2/Lhylb2hn6kRBk1wGgTilFa
MoqkHAzFe8UOfqYjvNszSr9Bb2UPM4+kCCAVNzdpBUKHC56AM6TFMPLHIdZr8o3g
RbqpkpcdKq9MbTadEqjVHCZWLWaQ9aqGJyWMa9PlLVZ+6zH6o1vjap1DXX4058Ee
voNufVYfWJunS/hb7qvNf4wbULq2FEdqzJ45BwVuY1L/yjB9sHjOho53Iz2/zQ3Z
O3XN/BKTzJGxubWU+Udkoex6IAw2cl9QNZ3mgwm4jk4R+PTYDcqIm9+nON85/jWX
AADPHW/8r98/aqP5NJ8oPxOpqvOpYWb9oHRRMZtS8baTvWVLJM77t3c3eCZgSVQ5
+LAis/5eBsnj55Dj3LKGNWkimlYwuFgbOk7ZWMq4/+jUXPEFoqJSdLGJKPFizF7Z
u6eAbiBOmSanHxmDo8Y0xS/hOO3c3zrGWQW0TqAOWXfXK04nBLAItwfzvvyx1h9y
M7piFW5jxZ7lxt7aE5Gm37V109ntV7Eai/NKGR3D3gWfKd8Tpw+nkBw/rd5gFdp1
wMm01C96DqNvpifWXfw1f7iMxTZYpQHsLpCSTCn05SAYyQml1p07rV3/0HQYWF6S
f1uUfh2OFja9NFaf5PWz9/lN6omGYaCDJ7VTmyB2ZY/qZBlann7dEMFGXAjUE6K6
CgIM8ehEbYT9jJH3zS+jV8O2B9Xqbfpl3XzNtaeINxkia5rh122lWRLC3RwBhwJB
ODNgBZF9jZwpRseH0OP7F3R7ERkzPnEFVhsKBd3HLaNz+El93RDhzM5TvHT8yEjW
T7Rpl+dEREcH+x5sTEWkoFegHNHMteMJwFcE3P6kkgAS4BM3bhw10hDDV/XjWB/6
TWJpJ9bqs2TCLGVAMRA2ZHEjPngYtbf6NjGTXyuJK5BhFLU9vHPLUwtS24DfCgGg
zBAU7NUGLwGhxZCicABFD4ZmuCXLKvzGYTvKwO86ohi+4BgQY3/RrEh3IqQMD2zH
2Qh5jDRgyG9dpLxRSiY0tXCJ8pax/cRJgidkyOkidBnSSDFO4VyrecBDoDWFcb5P
LCtfVoDMAn5Rcv0uaO2/Qi0+30YJlaU+MP85kKoY/X3yU7wo/S3Y/J7YjKu63nIu
gDxtQNmnGTY309LAOxXxM+Ixik0B3ov2Dk2BBum0JAPyQJ2gFE89PanNgUrTZujp
v8ru/eB1KsTmdaiiv/z9FdaAhgPnK191JGXvC4bvNKAq2p0AP+2LoKD7bYXYcmx+
5ME7l77S8YC/bDbJeR2wAV4gENKdnsGgqzOQVUg61JGaTTlgeuwsIl/nkjkIaVvY
orEUpolmswGqac89c1H8U2adKxPzuK8WS/uTRhvGV7v85WoQnB0wgFLttHVQ4/4B
ffIQ4pzybT3l+HzCW0r4AKAZMAdbY7ri7TuzlgE097wS7tIA1IZ4Qi57vIBclOrG
7phmomU4lUqnj/PD+ruBaGo86R+NTjthJDn1cnY4j5LM5n+V3tFUIf1Qh4LwkZDi
rY+VAmtS65R+rlev6yptbxnD2omMkb+uQqXBMHBjNt6vtsc4/KEB0CqCeZtAzL7y
5v2kan0Vp9wr0n1uvHKOsA+t0bsDoZ3zDDvTanVNyHDWtyuggedsOloit9yuv6d0
H4Ll40K1jDuE+Nx1WWMezpmQcELXvIS+sjIp7KLWK4PiIt8VgFCvS8QO5HLRwMbP
GTlvm4ZBRTSwHUIH5jckKVCaNvdNTV0r1rlbQgZn14zuh58yuN2bpDHtnwcZo09F
KM9xnCwUeglcG6IuHXmoYowKcY/msuaNauQshN1To72fkDGL7cIsMx75ftREXXYe
`pragma protect end_protected
