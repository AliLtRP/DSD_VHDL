// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:55 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OMZjjoYAQYqNedJUiDXVthH3ZSx2QyENO4Li+cHz1avaxmtPubcmqR7X50Zsnex2
0lu/5y768nDnKeJs3yTzCgfCZWqDN/4natY+6Pp4E2kJBMIzhqMHIhnfxHQNu38B
31aVvaG4VyNA18x2bxMMEmZHao48MQKn934hFYi32pU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11904)
ziHPWcxxqlBDYBDrsoFsoHEzn9nrGY8PbFimE5kxviFpdD7FB+vX2jTnHDP5KW6C
UbAp8lB+fA8NqtjyeO4Y86ua0kyk6N9XtkL5NRzCS1HqN5f+MZBihbKJUKQuYr8j
fO42d9SmNV07ETed0ruxqtnB3q2VR6GVza7ynXK5WFZtzuUjr7Ij2axnzuGGKfhR
kPQYzkaVKwDkzgD/MtKJiCpiy6GdqfA/T3QJJfZAGLj02gM6W3QYGF6jQ0k+bvtW
c6PCPtLaPSz4myvnn7BdkZQ7pdU1VxQ1KIC448G3cX4HHPGj9AVYvSmr/N5VuVRn
cqC1i9Y29SA+fh+retGRacyK3KBX02dEo4Fz2CWC5JPe4qODfNiM07cK6y4Wtpqo
v8BOXWJJH3iPtC0AD2JaNShqVTd0GftZDZn2wFI589TAt+U5wsNDL4lnbS3xYquX
dINN1bP+cfuUZ228mwjm0UQ/4p0+X+V2x5NKMRWCJBT5ORugArPXFHQ1X9AHL2fG
f1OuOTkF3qWCdDva7Kf6N7vmQ4K+621PGndZAIAbgQYM1QUaLVvLFQsLRnvlCu/r
j9p57G1fPfWWgXxW66/YAMvaOs/P245IDQ/jO2uvEH3+XLJS+0rWBZ6gRKdFH1R3
RaQ9yhXqerj8ODivq9Omx+/Q3jVtHxyMPcRQJXK2hgPhKu58cHRq7ZcD3TcnSFB/
azE5mfaM++CblK8bB8kwTotTfxFZMUqXMuRzZQmzo4bGyG3zHAGnaNzRcorRBxQw
Y9noV77Y9FxLtXHDAa5Db7WfRZ3ZmEk/CXqxMtPA2S8P1Yb8vvEjGvAr2EGNi3FX
VCj26HECfJ9aDmBM2md0ZgVIuHxblyJV3KPZUxyK0j9PuGq2Jg5IiWVyHXOhKQ77
IByoDRKSoqY1onLqB/F+Dzb6D8lsROpxBVTdj/Z4++egzi/hOZdFq6m43tKg/bPT
djwQx+ppEPQA26sB4sVVCHt3AUzuLD+hIQ7QDds9dB1jr8Zl8haQld6tFFBzhio1
M7slJFNyEsSdekja9xEIQXYQK7FbXYa4esqT/2ckWL/5Qk2kJl2ny1DiMSG86htp
fZvohowJykYR8hBnwCLC1if10cH9/iSvJsaXgQkwopmFVjkOd1KKdVW+h/375tdX
hsVnDcsRsYDki711MFT2KPn5+ZmoKIGDDoNki8pDJAnhZ+l1Ye/XZclEdK1ima84
IeCWvirzXmKF34+ji1naJEKK7yf4YDTKhQ98Yi3S5z1HNa+FjP8poGfsXIwYhrxP
sP2DJYjGtzr5BUzzP+ggRQZwdnWU39iMkZZJxTZxjseYPVrhNieR+4AKTMnhs4Gj
cplU9Epiucf4T9/fCvYntbrjL0/2wOEsEkyO7pemH5Vl1qYxoZMAWOgKwFX634tf
odZ7lhwI7fpO41jgrUP4Exa+TCdxGiJFC5c2eBkNMELlDWsIZrXpNAvV6y0GsFGF
U0jTaDwwqi1Mb5Txb/Ebw4IfSoRPkioKx4PJc/sijNOaRKQAiKJSHDx7eI3FHjfI
/OLbazl2qjabYNgZMk+ED7KX3ISCUx92KXvdeT4mZ4fRs4sN+BCERmb/qgFF9D27
1FSlURSPZEeUtejoqM7BmWTwpnB7B6xwoggYIhMsioyjGDKSpyNAXuiBscbFul1/
twJ3uwZzdwdXCaI7XgYymfYBcQSVPtCQ0X0G/7A/ZTeu9R1Lwje5L0uWZSjfjDkC
/60g1TyxEozXmr82jQ0EGBasqukOw6gsKQ45nmMQdezI09ni0GVdNp0ze2tuEcSD
9JlyjskujleW7MBcqSPC1rkYrDCW18sS/0DOhjaUBXRCCzLsJImICxavS4DWEyVX
/9RkAU3An+Zlq+JcOm8yTrqDWTPbuOIt8LhdFGbZOLU3M1Xy6KbjneGBoibPtUWt
n/JmMmcZIS1uOCMQ+gI82Rc4b9CJiBFN5zPMKiIPiXqhbu/sxBDznyxmMrzQdC/t
BUmpcB/k+dB+G78e/Zm25azyzD+klLKjcc2kQLsx6N6UW0L5OR5xUUxdLSPWThP+
xDdvu+upxSUk6Hg8xm3kaOI7NgEsYtpdvqrTa/Te0seIFNr3rqtp+u5i28U1pqsZ
6qUl0mg+irwexjfG2xLhLU0SrnPnyy3+vMJdIHiJMvgTfTYnX31vkYQPVOC17oIF
mC1nAoSWj5hpfEFFM4v4Am4cjnpboS8MixuohAUsIMJ3DispM9r47w/Cx+AMmdcV
SjpwLO1eZXGWNflqcTvWl3tFVTYIJOPpwiYFLgFrvBjWq3ufS9wgYX6POeY8RLdf
LhEsYl8JpQg7oFKXYh8ZNMHXbTjip3YUS/k1xgeDZ1Mo+G10fqI9qEU1uyEntBbu
yhv4fs+Wn3t1PZk5NeshRrIfl6XPYgslNEvHXLmNLKbpfTuhJvMu3hBnEblC+iew
Ie5ACgLNE5AdEWKkU9Nl6sLDou0Q7ELj32BpssYHanI/p00ZIa8og+yt/5Gcp20G
rLDg+Of0c9Eae9MjQdWbB9S61Y98ViuqSC77Gi8RB/hanx1n+l+xE9a1f5kQcRVH
6DFvLUUSMFh5w1PjBfysNmsLMORgxyt4jsocnUpomN7JxnCWkMQDdHo8S/2CzNYX
D0JevMbvDeuoZf2w94BMP5DIGA3NVMib6WcikauTfitXh539/uPbGG5l1Zfd/JjP
4m56sXbsO3qgW2M7VhQKBnzgu9Ab70RazBtyMn4QDX278O8wJpRaju5z5VcG32ta
ZKPK3oSCNJUh7Sqw1g1gTaFZ/3mqnfnulada81CDSOGV70brvH7kfgUSe3YAHtVH
0FwHapVSwABfnOiwSAkBXHsZzYC+Affh5GTjgDMoBIYuN8nsQQ6apALQVfJiRjXQ
a6bBW/B4XXpU6ovEXt8EllPTWLWX67XCTgjdpUr1prJiF1ifr1S6INltYn2oJGmS
rbwKeEaL7vfLQVzWPZNhKqDk7oxgsyP9EpDrSZv+eyX2HX0ziD8xAU8NIUWI4o1F
ZuyAC2jeErFl8wibzs80BDtll+8awgo9avKrcwL+jkayIeX61d/x44bCZ5rqgvAU
bnQ2l1U4yXMCvmxxHniiROePgVMN6Jr9RwAo7QKyB6qB48yDmVjpxZBTSazG8S0M
NrmP0HuogRsm/o7C6K8YI9o3QJO2rT3sHRZfpG/j779Mx6jYPMgJdp3FoYAGSVxz
Ot4fx6H4dx5GUn2n7Rq+HUuhDKA1kLgausOHeBPUyAJGZRu1nb/+Fyj7YP17/ViG
mNo6sUWntxdsOtTGxNdqvJip3GD9fzjrGxSisX5I7DDxoFRH18cEAEUct+elygYG
SbaNixw3q1q+xIk+KP/EopQOz8u4MskVxgVElnN1LTZXXp23g9hqkghBYQ0MvXrr
7elHLDwnYf6agCikjqGd2wfwOUaaFnUYM3IkYyUsmAyNm0bzOw9KTGHjswNFs/QP
eZEgYqslZALAa2FvLKw/jnF5iXAZXiH3KABY2cwW/2KMILe8KQkjen61iRwobpwo
OuCFZPBqd8ULSGINEz7op0ffw2N13fnK1WaIgqyXf86u0gnfoy5vv7qS3/TijL0e
1LxMHkpJnRpO83PANx6BJxlt15iAUnX4e0VVurslcsHo5yxBCdnd7bzYybfkcfm3
aQotD9Be/B221ztLIErz1BOTHFxYXTHKWAoaqNT2TJgEO6rz0Vk5+w8P+uUlKZDs
pR0JhzsoBYLPpaIcP7cfDjJA4JEACrUEPwF0Md5EQiWGk9SOylZABAf0eJP3M2nO
vbcdZEeXmPwZxILf6iX3CNCI8UkmVDr5dw81I5zdAxq5fY9l4TUBCHvZxxJmAMzS
U+oVecybU8pkhgcHpg/HwR3qOO85SsMlWv+yY9vuJ+/FWqILAuPkK3Zy3dh3WQqB
INoDGcbH+yagDNqIEFMx7B0vSRvmnTKqRmA2qT5/8LU2o6pR/oHn5X3rF8PR/EZL
k3X+uixPycVBadMix8BrckAu05OXXvS0EjFSBDSK9XNlWiOnX/htjUSzcwgDP6rs
eHQ6MeZ+RMnd3s6Rt/kVYCSDRo+ek22egZz4/9SW5cqF+Qq+s0jmSt5iSX0hG2uK
Fv0Xs1PkUS28HuCEXVGTeI1b/jhnYNK+F91RBpsbN0lR9T/udSipik0IBdluG8c3
TI22qz3H6neZCd8zUS85cFAP73arg4OVQ84eYQ8/6wFRWmxWlTf39Mv3U0heurkn
boSHQmNqkNIlmiwB/N4+UQN9j5//ADaJnSwY0lJmyZDSNFzDn+ZZ1TR34QLqxkfY
+yElaG3GjZuj+VgJoEHLux4OK/tjvjrlwADiS+GkXqcBHw3nFI6twGId5rgxTIm7
+wysGTbq/KwUYEezgBz1HSxxTDWKXYKXKJoycvWYwXVwG444byKlmCKeQNP0IN2V
4c7xiqAu3w8+K+5pNFDuQ3WLk2AeDkMw6fjDsnFe0M65AKmvfFnaOWFNRmLQxe5V
n+HZdd7zI2jMMNjB1E4WhL0aq+vafoNEiGU5nwryD9QwTd02MVC9AOeya6C7YCR8
gtUNPt8ZFNVS05s9NjCYkLHlvCM6IRKoDWc9hDmQ2OoD7E28R0L+scvaC+cIyL4W
NOT9S+4LVVd9F22/CXF53KFXWcVC/kQUzvto2+kaDq9jT+NYqfP2CdxsH5CxhIsX
E+cwDAdLrbuuf/jw1BW0lQcmCycpX9OzcpUGfg0V2OwA/vo1eLL3kQeuxqMOKWCE
Q487vhfGw8gaYAlM0dOX/5lUL+rWTeVpDDGzC5oy9AKy+kBa2LBc3VavwYQz0VoI
UDBazO1FM5pUCdXPOjcnMtvlSVKZLYhcj9bXnXviw7D9u3AlVPASR4DrqXbxaQ2R
/16OMSaytjNiz9bQyJYITtqGZSvgtDGnEGyuNQ+Gxm1Ohdgb8bxNCWtJEpiueyLJ
IL+a6WJ0vWMg0ogbyXMV0FXQbQS5cQhjINZmk1/EQiVBDqxz/xgWClV/+juHIdae
0qs2XyvDxYXh7IKgYP3KMCo7JUYLBJIFhbA3q9Imp1npE+X7e5bkdQ7+fJeo2tR/
qLI1SKGLtklANINsaWdVZa11hZuuSaPAd7xntgA7bqxdawi9uPS/dXvddMMiLFSJ
cg59dLuXZ0qXMCNl7eDut7CfmbFRzuE5Xs1F8cpMMAu43IWrBlPqf69d/SveWGQ7
8cWzqYlS1lnCb1edsoHUu8ZJRPOahHO+9qVWJmxNDDq3aKqq8F2Jq1i5e3yof+MG
jg9wzlFNVxt4OcE+igY4bol0l0R3KxGq4TSIj99q7m9M5I85oxla5uSuG4EllRdI
ohmQdt/RwK/bZv6aPiWN2X4b3dyqNfTEY5J9NcDlyh4dGYHaf8LPEwSBBSP0IAv4
7/UZTMNhdIHjDJh6Dsm+Z1foEVTF0tHOvtZBiz4aFASzwOOXEgrYYwLIBE0LT53j
G7Yrlk2fDNNxI/Tl2WiI1eqeX1zwAf9qlpMU/xbGeDUaSqvlkOfp+EiPNI7j0eh7
ozSnZGMDY72OGkEZgEA+enkm6YeDQr2v4MXY6e+d0QF/unr2dRgZAE/WSEAn5GxG
IGFh9VYP804xKDY0R0jsnbYtki3k+E/EbGNv+yfMLjW2/zLa1utuAV9UMd0a/68f
/XswFMX9c1OmJFCC4uyPSc9sbeU9SmhV9RYlfKB1kB6j/CCc0YPtmq50EX1l+j6v
nlZp88bXPRmT2vg5fmVt7N0cv4wRNRu5M3CkGb00pRDfqEy8Xa0u5/QnRfRT+Oa+
dejC4WwD8J1+HPHNEv5uHSycXFIktFUZAiClNynifR/O+jzuCzpso5+IDE1Bu31L
sBuAM2WhynPca1V663jzg6zUcjBSLTKfGsJczej0jq/XBss0P2mQIntxg+FkOoTo
jUuyl3jMFrfMAn8R2ldQVNGm8oXThejbTlsGgYgOSzqelMoYvy0iUaaViOYar3R5
yqKmSX1dBF1fWkZpqEovU8KpzrRvUmz65ztDJG57Sk3JPDlOdLhYJeWULA5lxFnJ
/jwyDl3iXgBPBJBSkt2+hztD/Pev44L0c/XK2iw85BsAJce1MKSXvQcFp1lep2Eh
bNUz6p9nXFL6b4lLyx7tIWGDsypmNggLw9P/KKDwPevHQWaN2BW7RGe8oxpS7ivY
vMA3HUsxIubXheyMN51qhoV7hCSpmjrORH4s5EJvZhnycOP6XxfIKfwRjdKplaQr
BzMmPuda6MfWhJW8g1qiCmlFaRRS9oPrG5uG54c+xCSrXMjFKRaWFLyzJQ7/m7rZ
9pdfpTHZzw4etx6jbIhxLSSh9rAEFneyo2Z2fh1uTUmI7N1nwyO/vtYFn9dIL5Rl
H/EK+FViyn65kw4OQdJdgvauzWo72wuGffrzGaJHNVvxEPlcuEpRHaHKSqU3HJdo
I2WpKBEehvjgIU2hFutt/a1nKQ88CwaFOfSOi7L4wIZn6ePaG9ZbjnpePOJWpHDi
xDbHarPgBIGfAY+nsDO7Cre5wKnO8riO34g48FB0cprtJj83fPcMZn3Zely7aOG+
VSfa4IHxEX4IgP9AEvfpasS9Qq4sfxi39bamPB70whwBDJCG4XqHn62eGcNAt/rV
X1HOgj2ml1RsNuVOk/NFbv7li2/DxV9HvA+Pb30/Jet9+EmvLeiOHVvv6IFdxykr
yH4lxE/8oEMrR1GiQUqofYDfPtR82CA3wMivKgOtmifS7ocdW9UVlCJhn8oXa2g9
wJ/o1+ffgoH4oe5ehnL7wJUZdYJ2Ux+w4q2ogiNmP3J2Y/mRVAj3B5qLtqxjaUpf
SaIq3/BrJiucGWQlbtucbeewAHWAWbtG620gOYn5PNwW9xUjTvo3ehODvUGidMGD
ZiYYeb8sLIgVppema8JUw25qLWeMCG4ZmeR6nKURpO6kMdW5DOM3zZGfuJOKTa1P
3/UbQ546UOQoR25DX7t/UfoXtL0YsPudYWtqkUWOsKsv2/1lYSzgEHFB9N/4RzAS
vcSoA9fSuiEUkLEyR6CDmepnJYDDTa2ovIXyO4wm7Ivqi0rqDt0YEpU0CE6B6rbk
VqCLHmYJR6tZ35BWQMlpSEu6O3mzwbA6Pvx7590KuUFbZPB+k5oviK55QDw0t+oC
NmSIRkV7eRaM5hMd0v46Igtvl57PUsKSVyWAExnaYGjQ9fhZSQ3V5kUUKC+MwX9N
QChc45diZjIOl6cECB19qQCppPdS1NqzMvFwNaWHV676Dh+p25b+KgrcKRiidPpC
h0ZGfRn2BVxYjXlyFWcVm+uhA/uZu6qUP8/FBz4f8bG+DB/duQQvlgB00Ki8b5rR
+1KD6I16SOiFUIqjR2HqjOgr747V3ecctFj2vLnHlDaMlnSwC+FuTt2ntB9Amnr6
gUlTWNHIjxJtt/1eqY5DJk9nv5UFzN2JQ9ONbQ5HjIxXBvR5o/zzBqVE4IjDAahH
WDEmOAfu7WWbfVwApAML0cqlWR1i8GkTMa6pMMuNGWhWrTuebLcOII51LA1joNBR
WUUIptDzUGhOylmmoCescLt2wXKv7aZejfg3CmI5mEEe9kmZBgT90uqKyxu0kqf4
4vRV6aNuFGSY8bdTY2xvI9QfIiqgZUapYLWrCk0sebS3TAVEZEHTnJumQLF4PHty
/i3e4rC+H80DM+92pr+RlzdxaUBZhQpwzDOA10BzF0nRoNi0N+osoQDlTcDDdXr8
fs/OSqjCgwDEk0fMt3SN8jmUhJinZ3HLwgMNO1YmyRqOgVeMaM44PZtpZamfNxeG
mKkQpw8XvlCmayc+xtt0BHK9v2E60FgL/AqVQrNwaU1ESfV4LDrtxyYUlq/RBMlB
HCeIQIGcu4afnAe21/7QH6aweAl7xLEqNxkcKGX5p7pEyDRIr4MwRdmJARbmGwcA
LoqvdkJpyDeqpIFlkgH8PfGzD6BBR7NUjx0NaHXK5rCS6asqgBeVwCeDwKUojqPe
UI/ZoLOOClwJrfD6BUgvxXktT5NSGr9QZGdVb5mWRh83LO9NEdrwc0Va8e5ta/zK
8fEDzkK2d1vmE4Df7mF54LVzlfIyz46Qr1B5P0ypWQDHPAwMam0iFrCgKbWp8p7n
rTidw9NzJDuAK4m4OK3nBMEBxSlD5TVZsrv/6Mbgn6f1xjzOru6U2VM5h87COKBg
6bJpVXAqCnpm6c3JmcG5Oaj2/ruGwBk8uxddhOYuNO+ApYff+P63oD0KvcxtN4JH
6YMm7U8PMj7ooTTVhLbVxcDWrLl0DQ/eUUrwPyIza2RFtIW0cQKdElo5fXQiNZ3T
o7H7frIdNYd/7kr41DrCHUBDh+7hCIGLhsSCF0p1QKUn7cGGDRnMgFNAziNZlVr/
PeEGwWYvFXmb4XskIKpp1qZKp0AThtZB0bcvntq4EC4x4HShmauQw8jm6plNqXcj
l12Ra4WehXYEpQSEPQ+48PjLyCx0zNUqZIfN1/vVoVxG9rUMJV9ldxEWp1ZMhK+P
hbtKXIpkHIZzOypSBzwYp5G59fQxSTPIZRJPKcxabDbXICqpBwzxvrtbA0FHoxUl
dw4QwNCGDLpWmFzqV8maNr4yXAQA5/lDgCLllRljY5u/UmPy7fg9cbpF2VilTzzQ
A65ubpejPphwWRLVNnY3a6zKMY0rxSfIF/mTEbwsgD1qcMojMlrGtya+iwzRFEd6
5hfss6l8pnyITrnlyHlruC2ChDnvrcNDfrxi5222nTYlCMmPPxAhiVYpgJnfaapq
2ENjmbQ2586yaoOZ0Pmv5mpXq7a2BVyPJuPhisoyQdwcth4OnDCSm9gJ3jgdGKCP
DcjcZX/y8fR1oqg71s0ofyRSYL1+MZnFeZqU/KEIVRd1Luhqo8DiBtogfiHKFnO0
TuU6npj5FJ4GaF6hUe+jYrhnY50fmpoyrNybCXAx0JjAEasOkOYMuIvPZSHTirHX
0MsWHGGIk4JhPknAYjIL/vMTfJS7lJ1E+Ec5Z5EWcVouqgjP8ViFvkDxdrPrTdxb
aLgrxY212hK3NZDpquea0aK6gAyKc7WsYE4fTuB6qIlWfIfSSGbTJ/Kbk1F8TCo3
31MJLauSxEQx4UXn3XhQjCtwpILrp7VG/xtOs1PtajfJ9VMobUt9yftg9VsqvukQ
VXmnbqIBCvaHEWlicvb9iOBUE5YH/f9VgPoMbWTr6I/jC/hn8T+OivAWzHNuOSno
sO63Ux5IECfT3wB7RZNK/0hkY3W2o4UahW+IWHuc8VBgxJotbhDKuLOvx4AzuZj1
NBoBE9KsfEgbAS+07qaa2BGp90A20CWr2S9FZlhSgkH0LHlbUNwQqCbM1MrRJuLv
LZ8kvRu1Iw08wHxCdtv5H9hvWPNHvDrb1Ex08UyMeOcYf5FgZ+3J3Jm/mBZhVsSI
uEXdlKbk1PhVZTNQCDACTqV8b7bt6V5MQNwDE3ZrpJXeiERuejpp4f9AIWDuDXJC
tqK5OQyrr1tjzFHQNTcsGC6PZGvBgt1G7v8bgVugwnRlyTxf22HNqbntQKeQQ34H
n3P2laY8DUeTp3/1zGUIrhhMIfcieHKPp2tl3LaW9PRJTHJ2gueM3RDy0SFJWVOy
WweA5GJuTtHQQ1GWBFTKcWiwe4Q9t0nBZPJSBNVJnmpNSKEgM5IfZ3boH4XxxktQ
kdhHEnI/NhX9pXFYJZzyj+fsa4YYuEku7wc0AlpNJPSG3Zb41Xk3M6XJK+PCU+iY
oII0xilxyH697mFGyfD57137qcgvDuj7ihfdHSj6XUXGIl+bA/0YJUyGcKJTCe/i
kqfvDZrtZKuGwTK3HWX4b2xN0053pRJqQBykj2zqOOwItZr/2cYcUpFQhXyEYQr0
I9LSCvKI8o7twODAQphi+QcKcJbEdZjMlbXl2kqpYa19CTYl0z6Qv5jhaY5epRFp
n9USEpqWrW1dOzzBsIfVtuNw7ZpdNoPdTyriuDSVbg8fwHJ9iKk7ZFDu6VCg90eW
F0t2G6OpIeEouqolM6AMGOrABonZvZSsayBNQPrqAJDFvZr8bVoMBMrWPOhYdQSS
8hrDGZ7wY8/0HFvEB2gyn13NldxHSoSiDBhLtIzT8KCBlk4C9YMqOxZDo4hb9MxQ
wlSANYSGbbHOJPH9vbcAQSKNQiDuUiL7bdiZYOLmUK3xVdHi53/7u03qL69LFm0U
AXB5z60bp66RhJaqh/Yj0AlJt08JXh7hsCHG8eI1k3LOINqMXqBhrz1J11GyAVuk
QxHI9KZAdiJPuqRboY8HXx1sxIhTJhCeTVb4SkHIxzqA8rkjW/oK1Gk83nti+/pr
zQrnZqTNLSYnYTKKcNrboR0CCqJn2JhvTTarO3aBNGwrAs5aHV7WHEq2LBi8H5CY
Be3XYpL45RjjjTHpz1LlJCguR66Rde9x2fR1wM0zAkFMx5P26JlBTykwv7p36WUH
VxOHkb83mBDvppoJJ9KpZGRMYw++mfdVrXW7swc5komAC6NFlJI38xQUH9t5Zp0t
m/kmP8EF6kvbBJiGKfi+56wraCwslU0Az1ZjPSsuBci/o6CpZtK3p6fZaCmPTstG
ZBCILMOCsn103NSyMpx4SCQIIusgd7DHqH4fPjJI98cNOOQLZ8U2uofw1idSVqJx
WBqYqCGUyYRsdHImhsvNBxFarEqldfC4VoSk5KNn/rN5UcFF3Daq+dC0fzCcFobF
rCs8Ta4+7rZWKSpFpMYM2euOsaJpbIckBp+Vyv3imugOBLS2HE+9VKwHtd0e5iyQ
0pSCyEvukrDejg6IEoMJR8Cxf8pkvpCpAt0n9XIsVXZNulHGxuctbhKQxJ/RL5Jb
ffmFl/ebVXyE/CsHr+ebPjnswsaF27FzS1uUX7X6gIfsMcsCg5qFtEYF2j4HVa48
502+EVGN5PZfibyYP9rldy8Q6O/9Wb/GamqtQXz3KRLBCHSkErYzHbsMyDCBNZKJ
xald0f/mLbngA5XQR291LY8g+Z3/dMLaHgR3xe/Ja7GD4SJ0Mmvj1CncvSFlEJXl
+uBn1ZKvXmCpzrkFuAU/9roZJlKGgS3fbeutr2GpK13uLUZDBwdwM3p6IFTMeGj4
YqmbggCYZrcTOZAhEgTS0rgPiVf9ZEhe1peBz3sHjfpbSRl3/7vZLlj2PF0Lx7/F
aKahfKTlBN7GCpLq+UPHv4soGlQRqdyQ5zpk1N6Yph+cdruEhIx+SVW86OH6Rzmx
9rzMtj6hh7xW/ipWITWM6Zkr2Vskmv7I9aaDs5qxTElFpOHk84Kjn76ucLnpDN/E
rBjkGbumO7WRcycmCGfFKqn0YjDPfsZiqXNcOqsDzlG2ZJCtBNvPBeeJnfUYhqem
vD1G9QIyoKj98uaSyICyzR0LAKDR/Jdng2eSJ4EDqoCVMEHErJbYWdOjk7eo8KkF
PV86aiwdwS8UNM2fWYyatoQJvRUqDydcFhfYu33h7EaBQ50feJrai1OuopRkK8Xl
1IvxR1xrEyxMh7mxWF7BVYOEg6TdOj73vsQ+Maxmyi+vFnyqDMnPhYbf+Ngj9zkm
ACSUHG6Gnj3xGnMDMnCFBjv4AsAbIMc8wKciS8bq8SGKxJEbnQvHcJlwJvmtfNHF
NkZthDrgbTk3108oJUIRLqWxUAPEuUW55rBxEIHS6V6hND+Z6tZn+prXilMSh7pq
FFdv4wTcOHARN6G4ElIUT1jyH2nUku5NOzwhVAO2Ljx1uxumFQk6dHOUvVeDO+Uq
IxkWjXLDu8fHZJIzn6Ta86hGgmTes0cRdlsntpTx0+zYWyU9eE6T5EuPgft4/IDU
thwAyaZ2mCAdePkD5Wr8oysPF+Ekf5Yi4JTcHCsG9Dqz5Mk87ZRjWllwRSLUxNrT
0P8AedAa00T8eoXm2RIWIBJ8Ebl6sVrYIWgFmbAOQkU+c+Gr2LDrhXeEvvADsyTz
L/xisNTHZbFdwvpF9e0HCdFkE6ul+Mma+8B3W3VBLItMnggF95HnfJmJmEhgq/ix
8+89yyMiocWrnh/T70RR1QBoKr7UWeJLEpWTlf+9uVc5RsD51wjFis+FeH11k3sN
/TG41yuzzLIBcvAHom0Kb3R6zQqNYHyGnZlSBfdZuRM61hl4yCtJgIOgyyNJ8z22
Gr1iVCYEpM6nEPLG+zPFZnOf/Ap/XoOYuBjiP9hb/xDfrU7zqMCf2vZwucwC0qD+
7O0jM1tKzPppJoIfQeX/9CMXq9DIRsHLfeNjJEeCz9wEmhaKRSay/783ndNynWSR
00xYeRy11JPDRNrPJhSZ4DHSwF34+YbzU51oc6TpcdPONEcwIDKOQPnG0NNLntzF
Z+KzC36rfuc/CYtrZD/KtmMftfScnnlEHCsUP+Lf9tafJMsHL3EuOsRd1FauKJCM
AeO39eUADNeORajipMH/MOO2jF+YwW5n7hQe9LChep6nMNhmLiemlfkc5fMwAFVY
A/zpOwDI8yU8w1/Ot0WScnjZka6CgmIsh8qtXo0Ifp2TNqdXytG5oN3DqsNeH0Ra
USdqlWLWDAGuN+IU9YYwQ2pADwGg7nqvI+5Cwf0ot2gSBAaBUrVo8rKbGzar8a54
RzLqd6vB1ZQQ92t1XsHH/eFnTWHpgqcbG2KEPob21toY8LuRrpsCauG4oICizCza
Vu3GMk7RPMa6flOFoBAiaROAwGxcIr1ea5zllpvXdtp1TTrjVJI38LfyABEAL4kL
b+2yG6X6DHzeJqH5+PhrxO7NCaGZAZn+ZpgJIIiO81tCCPE/pzHzuKdsl0gMp/yZ
qK/jCraukzb8Msgfw35WHpBq6Kv5seNySwsz+vLhOhgK4Cg3qjzdddhnk5RucVlv
F5ZN+5v1StudLxg4tTT2zeBwDS3v19VmDUw0nWTT8Y5TNnhv+53vK1iMjmmstvdp
6tKqAe/TWCFeG/W2MxdiDNTmnOa/H9uxTO1f3wb37zeNcgxPqFPlrp8iX5kSwve+
Y1lDAu+YQid+B+u8aUoHCIcHJ2fNTRh6lWRfqrDKYpRgyW2TNosgJXRvc/BR+JXd
7E/dKUddErr4Ju2/3np9KvKdSueu6/Xu0CIPujoXE8vliVYvc/7LxXXfthgMb8x+
K32Ah2+iuOPrDtQGvpBt5dfasGxBeozKyy7w9rjvna26lapnipURfDs0YYgBIV7s
sfgRg/EF/26g94SBZa1e/rNSD3yCyV2I+4KzVp/jRBM9AGre4DS06vj0PymhYiPA
GP6AcNty2GnQlf2v9ccRYZrpuMd6tSO11zuUf/IBYv6VaWx5nzhPQSTYuos2HIqv
VI/RQrLfsOJF/PHkbFoKIv8KOOXfMyVggrmthtKBknUEFzFWGac+siY4SEZkPVfC
kvjlXDkPzqFOlapKfK00kERvBo0t0SQR4Ri3f2AcRKxOOTTXIkQRPhhNqn6bR73v
tG3XTomFlukp5yZBadYTah4h16nN2MIXnA7GAbjJcEr7FqXmFg2sOk/9O9abZ7fg
xtg3BhmLvnJffKUwBU6+IFwL0aJBfoD6JcJyw26gKkFrf8ed63qKodnXKI1tQwUH
kpcbsD4bcojHg6+zJJ62jl3G6mmWLPV1d1n7AKfPN2eGXnryC7kWYhNmp0QiaFjx
i2YCDI0vZZzwiZz11VftVnRak5wkBs/yug5uAC6I9D4vi3+FdmUncNt6nCztifC7
HJTGwc3c/UO992sMFChi9wsYgOR287CvqxcxVdQC3/S7AtwoNVtuHN9cHfgGz/XI
cCvqfr3bypcyTjpMEvJfmnNZVu8JThfRo8b+QFImFTkIJc1X8NgABpa+tZ+rHaFh
Oxk+eMlUQtIIydlwn0/0uZ6h+iMmI1pGfP8rfsVUHfwlxSbqjoogR0VPpWaTrnlx
kBzCgS3i8qKI7kEr+yvSuQINXd4D79Xeadp6HJuC8HRExEtnyYf/YKGWbxivIF+L
TIsZW6d9vWORwVpJGfTscuhyTCIuMyIOIGZcBcI04x3jbjXM/thIsVrmO0uOg1JI
WoOTXaFn0pOEtG6kxLRd//+qwa7t6Gk0m0IU52CZVezJ4baKtOiy1Cu2CBBhVzLm
JZyd/zjVSxAJFdWLlrdEiv+S/+Hw5DtgSKP6P8+7Hke88bkfZ8YumqF7j9M6Hu0O
dhYj5Tq3+L0M57jIvqG9fuHgjTtXvpmyAkAZ0ALjhehn42Dz8OhAOjmOHDqj9ED9
NKlWOAGhC7Mxi3+P7rpEDR+jN6UKXv41gZnlcWvZAO6qftBADsks6AYqgrzJs6R8
ONZxyyEYXMuFuTbgoWk3V69kTcBM+DYpgwqf2thFecQ0nlDnwsYKD3CGCkX72wDy
Br0d2/r9kZY9ecun9CH9/KhSICK+ZM8dhLWwkJpbIFLb6CairIDD1FXK37ggdhjq
jbURBzH7c4IxqIRm6xOONGBJNyhNIH4M+ECu2OZHRVfObsLktrwDLTTRIOL+evgK
ib+K2Ccyc/HtKV6i8ZwwrCEgJpyBPyE+RX73SQlxRZZJmekabxupoFr0vVnDW9ws
QVZknhlM7pvv21+1qOhtbapkUvlWvgkfB3RnHwJ9joFtU+YRLTV+GoxbU6HyYijY
F/He4I0VqBc36JiFEwSoKvfX9DQcteg3h5LdGXyq+pLA5RJQFgGI/87dsccugiw7
ImSQDm57KBa25rf8PBoQV7MvNumsAOyB5IKA495hZIp1Rww7N9LFLf61SjEQcApG
p7ckIOp9lymY8ekJXKf/GP2ocrUDoZ82mTYwhzMabzpWKRaip6l+M/rQyjmJVNO6
CCA/ofICKm6MZWI/D50SsPmOFZM1ip5nRYkDLyMxGDwIh31UA4tq3cfId71DUwxT
NpZRL1LwRCyFS7XRaixHSmLGZduB6y0b97wfwoKOww/FBAovUqJnO6ohDDu8RcOh
YH9/SVmfChhb/lnUrRCedzJ5OGsSeutC1l8uehX8P+tQoefJTXrGd+5vQsvd5/Kq
aIvIVUtWt+c/wJbtiDjCS/0X2MnIGJ16hjwQHeyd0R9xzriS93vwL0n1dAef9i9q
A6jtsI1ChDwx2JqF4zEETPeLv4mYkafl9n3AbKx5oCnEWJ+oyD10x4qSAmAXpPa0
/Ft5pNI4Ds9t2jWGPKVoZr+vcBj2bL2qzMSbCGcz0SWHgkCABMki5MTAgmMhNoJk
kdEeg30al3I3amRSfiSlcHNSJFdgGKKPwpqrZ6kV/R1wXFcoOROUoN8yiBC4DAMu
BrJMehIR8Ho1PDLnWuMndPugZPq1bxViWCz0boppf6UCW7EiOvHIVOlI6/psAP3R
vo339Br2FYaHpVmeiwdYGKtZrF2qYJifx7dVtek/5MFntBrn/MyCmmeD3OKhvpfG
oU0b8GQaNqfP8wTByrwjaoph6CgeFdNHK4qUyjh1hXjVH+0dYIVfnK4DxYMtEqJD
Fcuox5VeziXoLI5B6SXoeSvp2JUaEKm9TcukWSsEPaitgp81rFfgl+405Vr4lugD
j7rl/O70oejgZHZxQqUQP+uU+RUnuMdS8D9Qih8aDGsn7+LGHXZ+1RTHWHRfgABn
knTdG9hItp3m+YDyb+xfB6wDpcFgeUSsOhdHMEWKHoxqzOdoCuYRQoqj1W/w0SZW
19JnVS3mtdsHeSoxrjAO2/AyP3TuWJdzHwMkL5QeraXaLMFxIWwYPq08E+1OFOyB
CcgXVZlusKQaty+KE9Trx3iCOGPQOOa/cry8PsiDRDmzjnTVX2VkeHPsoGS7qHRP
O8wElW1vZich4eAiB/Z0811xHyoXODiHc+Nt4dhwdHO6qdORYf0+2Gj5z9r1Hu+c
m8OcH6ZQRwngfcKPWLEIe8hDDdGbw0/UMooQnT/36iJ/O6hIBf3pb0Cj0PoAHjYe
juKGDr1VWQFKVyTLAMnIjrB+z8U6Qnr31UGUcJDfZCxwPUGMA+DIcYzks9tRjGzA
f8uc8FT+COfYfMZOkq7EvwPTyo4YmRSRboxrpxhSvZ6dv+xKjwNAkxwsyQmMm5Dn
`pragma protect end_protected
