// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:56 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hX1+n/W/bv7iVi8kYFJoKCjqU6OCaQDgK5Opx+ZZbfQiW/LgaNe2k4VoZnlNrdzk
rM8C3cYOpAMHWX1WIzBzuUFhqj5Sp+yxYEm7IPA146d6kCtP9d48I1vkZiS1Vttm
eqGeVTTPABt53q0Xa+RUmurMbcr6yx2XozGMSFRh1lc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8064)
ixK+2BduitlQlxVgONejv+kbDnx/FWIyNQxRZMeOcQ8BIz6N8khKuxcdpY4ZqlDy
vrPJNLjTUiH2lnWCGpeSuthE0auFm0LbBiBdMktgOKsHNihqKYgPqGzLhR0j2SXO
HpgwYJfE3KsdvUHHMopIAXxzBU+S6M1QHBjz6MHzz+CzGR0ikfSjhrP6l2YjrJlu
+T9paeH8tPGmo3MCzKvyAE05oPkqu8ugIwC1YfjnjMFJKVmUagSqrjQ3Z+eSl+DP
IpQc1o1y+lMC9MRwmapugh73G9ErEps3N0ARd14BgJoSDI2l4RdwXeRrHWotpi89
LKEcPx9KQPFAvAWBiyUWMQKIz6KoPYAnC5/bzy1wZkaXxScEMsLuiknWgiERW3mW
HWDtWs377bDm/hSshuJ5OXECvQdeABE9EKHyc/IJLy+Fm70e8OL2cq2ErKHgbXwq
7bJetKS5lp5Jdyq6M2oezAYHDUaf4tiwSclT2bt/1SSbJjPRxrSjCdOmAE70sQrn
H7BqSeuMjN++drGCTRQnUetLJzTef5RYQD25sgpxYmXHb9t08NhHt/8x1otLsbur
5LhGvM5Te4mnE6rligKeXzbV3ry9DQ3Ou7wnBjvz1bZOCYFPuavGomppH/ESih5/
ugw6mCDUPhl4Dt/LGfxKeW7wZTqXrLHL2QQPh8alQryCnOrwU9UpPyAtjAvRj/CN
zkPlozbFjDczfXW1r+hryD81jDzqMBqHA727oqrxjsWkoh4iHcO49TxvOYEJaSa5
yQXtdvM7Nf/+7rwZtuDKCvZN25EojWSC8SYzKbFNXz69cunNm4cNrrleta9EmLFX
hC8vihIRK5eas3U1ypElRzms6rXMrQkeMsKrtNq3p2ev8W+89tiqZOYJdQcTzdJW
sD/GJc40aW8BeeWWaQPHqjQOqrNbI3AhXpOquv92lN1u1Eq0eT/eX4lmoZKdlzih
2+AxSGNaknTcIDPsC12sH3cDnzOa2Xaw1RHhLLXsxV1Buyt0RGnOO3rkXJK1twBG
EuBrGVlFBNkOTToYT5MEHyvII6UqAzUrrpEIAy2w87ecXVrjpXK8P+0XkTXQ7ofu
g+kIHmmO18++GY2DUE94PVsnrNtfn+No6XWUPV6mlc1FgF3B+BAOfLw+tBv/IH1a
Z4Ul4tpYmDBZ5DIKE7p7nZVRocM+VIk4Mk/+ERcS14nxooWE3dUyvJG7j7sohDcm
tNu+bu/xzYrS0nmBYfPDP13eITvT4IFSLEeTSewYll2WMTAp5x/S8CdZlwZwfBrL
pTxjtT5E+kTnw6xvXhYO/uo58GxARSxz557E5uS9XyXScw045FRiouOEjtLZ7vzV
hDYq7+egd2aXk0rsW7H4dtolPYecqxyuxef5HQWSZdx5eJBOQeJhXPyxL9mHBzCb
oXd95RSLGvuoUXrHKwETZL67Zr4yNCNoeIeDATETKfKEH2EEgepGjsUMU9j47Rbg
0whCU3sgssPZzaVLDYSw8i26TbycxeY3qfcVZK9+BA3naEoKQU7R6AerHD9Y+OG/
EeayDh6+lrPiZrpQdeXY5VW8HbFLNTPIzkTrnKWzMuII0Xw9e3Pj7X61aBmVEeLe
qzAdbf7m26zY6oCMKG9Np7NjEvHDLB5p194jLH9Mp5tqzo5LJcNeL9RKJ7unSAb0
kAE3ZG5drbgMabm3bKa+0omIcFb8v9XZVhAYqYhKUFh9YuuMTDIGerwBJKjwaMDJ
KwHUIUhIeOphnwLTjeSIF9n9i4iO6nK+j2uf5pa7AWSloLlSWabrYcqgqpvBURc8
Dl9UELtVFWxk/FgMEnKgzCX6uRQPpG6+doEROyPCxdY/bNlW4tnorS1Jyn3Nwr23
oVpWIBsBozsOiuob8KlnDrPyA48rnTQz7/wnFwbMcghYDvaN+vqOrp3f9r2jki53
4lz8fG+F8xu4ZXjQguw3d2wld1B5fo6z5yLL9F+X6isSs5wiwc3u/ce0PGlkDQI3
jdxeTUutOZp8kjDbnfQfMserQaC3usSwIFghltXBcwFQjonBTlKKPTqVyTw2pLDu
DcR639GkWSCdh2EqYZRkL3vef6qlWR0DhpAeHLQ1SokVKQiXjSzcC8BHJ5zXw+ED
1uY8EBr4pDeno/VvB/qVNjCIjfM3XfD2HM0up5ITaSL1HhHwGk0ighiLAHX6LJyO
mgfw41e+6u/hShtLD2NIE/kgJNr1GjzPpWuemk2fY4zVbzPgHX5D2BHGw2SlPrDZ
oDXUVxTH/ARc85wIblmCt3YtE/ZDjk+Gt8Xf3/CPRVCKWADf3WZV0Vu1dUnY95za
nC3KPSzhIaR4GRcKYziQMblI5X1XQgFUfbFKrla6J+KujWQAbeCMzBrw0jeeqbF4
qddohNlO7kJUmmofQri7c8/n/FMnYCr6Q7SiGx0NSSTjkvDbKRA5HF1FTMiHhAn9
e2xgUNFe43nz7esRBFO35UqfhuNPJGb+t/OhatOh6J8TrkT9iAeP9LE+4ci2IAmi
uvJB05H8GDrZAp13QPcweMg5iV43z68VPML7BX82xHMhYcKPD4EAPPDtNKtDTWHW
+FFM1oXCIUcY9/50mEVaWB8F5n1PoiIA49G48JI7OB1UMVPfio+HH0QH5VHUXZkK
vrM13BkeS1XBwaw34ve/t1sNAtKBAg0+j9aX75p0Eh1Xl34WIwHSPQMZOhE4g9DV
5qM+4lbu1B2+8oLM2Kp6Yvx8V3IcfTKU2BZGVa5RORVZtz/jZJoMoeYnrdTaAqqY
FuC74JVflASLvitz7SC0wUhhWdtFIn0r9pXWlH/wMZMBmDu4ISESyo/bnZ7M91QK
yQVT+6hEKFRyRNxs1O9zUKyFJSKApt/aRjgS3hLeyFLhPP3UCJznGhXlQTSntpBZ
9TfmQSx8Y+BmaWy/LlGBGOAtstBDP4Vb/XZ6QVjU/GwlmAXcqQM7/e2Sz3jDvm3B
joFdFNdd3c1TY7Hn92NX8kBpuXNcndlJ5Gyqf0c18IByYlaUIueFz+387Xbbe9Pg
3avu+E3tENFcUJe+M0fzp/YudiGI6DFrJ5exw4pu1Pjq/bCHFbGFcAaBsdN/xZ9t
kp6O119EGzuYiLU/4Hk/9nt1o/Jfm0zISXobdIJZT39WqaqXncm9oFger5LTyNzz
/T+LJdBWSUM8BO4WL08DlcQXfVgmE886uNiSdJXSpb8vA1p3KOBios5uC+Z1l5Xl
/NXZxWrU6obAhpXWeEGinnAQxRryqbcU3Nvov5C9kUr+tAOonaGEi6RUwN4kDnU8
yyDVdIpiiGg48an+g/FQtpTaiPEMu6jz2IIZb22jhfaVqBkxv4yW46KiLV5c/eG8
5NQVYtucIxgVM+VHjf2bGTaOr2IBk4Krqrk57MaD9x2jYHoV3lDQ6XgvFlwosNu4
GjcOWPav8QVW1adSuAmiXcJ5e259PE7fCkPcWjE6yOLUmkC6KKr0I7M7TKFx4gXC
CWxma2TDz6b1IDJRa8iMQhduc1mdUsA81pgJ7kME9bhqL9oa4UswYQptwOpUoKo6
sernjrImb+YVUAVUKYaIKh6Rkken40lAzfRu73O/VqM/RmfKDQgLTPU9+lYbJNPV
qZag5srbwgbW1Df/Bc5rqM+O5x585HEEgMtHnBAazZfHsFCznEtagHNtXjZPR16c
tLsqlHaFFwwuVFQEIXkmu2hcUaQ19uKJCL4wZjqAh8NVgvt8qoN5mGUEOseLDjM5
9SFmcPz+CiuIu82qKCgF6trE+37GMA3axgCl/0XRi0lk/YgQduRJC8wjMhcUiCEh
tB/DEW3nsXXIsbPW7m9T162o2yhx+XBQJnPY7Vd69rLspp0VM/lZ1nCgUxuEAoNJ
E0UIOHYeEstRT5Kcs9HPn9M05EUPzT0kCsLHnHJOm2gisaRvDVSSWt1GIvFqyLci
GqafoRfKnJh2773ZUcjBFlzaB3QHrQxK7dEcl4vubVL44My1KhOASpXRVH6OBJhl
RRZvimqOXKNXUvzPOD9kbTtyxc2KY5wnXdJAxZcos/VvY8J/xidi27e9a30CTVyy
TJK1FOV8zKDg4VXkgcYKMN24i/B15D2QvSHfl9SyDC1cYKXjV5Is0bfY+Ei4Xx5M
bym6schRObfIUnK7nzb6UTJwrwQMEuuY04/garSpOCLIxx6zI24N0LzGGzIyB0rZ
A4MgnVxYEZm/t8poKTje49k7DmSFsF52h8Ucl/Ycvlzui63QVOOFnsOgJq3mBfvg
6QNpk3MBw23YOWZwhXkXiJNmGDlrqKb3kCj6yZCtY6RDcnwYTGd645uY3muXdKE8
vk8jsR93NvTmPVnvRo/w5huWUgnJGQxQvsYuCPefcwzBcSkX9rYmtGggUAVrZj5b
ETsZuwOAnXm798QA27ubZVLyMbMQuvq2ddec4AvA4rAMplh4mhfM7nF4vr2oQz25
YztB22ILQD40ZyQ9tfssrMHh+x5tIbbIrxo9Iye9ywWMI1UITfTOxuRQ0O7bC1jy
pPwAndUSWeJy9CR92sv3Obj0UbzJfG12mMbJcF2jaKmulTMjADqv5FdkicVo5G5C
+a7UJIYEU2+Q5FMSrUmnZMPUfXNPmM4fOJOlwwS81yNJ3TuWWqgs9uWL+oxNq/QA
hkkWUasHFXKdZg4uUMbPAjMlT+ZyQjbmA+EmVkTPvuKm128ImSVqafD+VZ2qkR9t
36qDrCBsZkm+bz4C2BZLrWrkkRxM4afD/0rn0yH3lqOq4ORUyWxbUFZvFYAuYgpg
tb6sZMHpZnqBeSVjG9+7TeeyAeSUsGoxAolyPAFaXvFKhsd1dIpYGVn4lnwHguAr
j+w9OfLOzhtaEyzPivgUaF+lwwzjSTS1lL4kA81u94u4vQZ0BbAwo1kvuon/GxaZ
ixay351QYxMoRhB9D+A6SiPpdQIauqy8fZXe3w9fWJcIkAWnXVXtel/EiB827L26
e0BEOg3aj2bsCN+aV8gtcjxWX11oQ9Zi/3Y+KbCUzCDeb8SR0t4YO7GU/IvbcFk3
5arl9QLkpxzdsZFa+k7k0zyhPyJZaXkodgV5XfMcTXeDugwka9lu3M6Nu12cuHpX
V03ygnxwW72FI6sDn/hR7eBeYURxca0j2I14YTXxLx0DHwr0YSj0OydzAHke+FKk
vYvlzfSagmedEDmUb+GZzzf8Fi4XnkuvsTsvRXSoCSg1oJ3/FgPWw5IHi3yodNAQ
8ZK8/8j/C8QkSpWcT/mxrlXT8ZEA0IvFh/hWBu9yvnEFT5fjCsOM9agMo2Hd6hN1
XRYkDjD317TKZr7inUW7wdWgqXm5fnxnYyQcgqYZtln7jcE/JELCN1MmAf5C4nfh
85W4mK45fAuHAiyKjoM7K5PaIRv0bfpm+/ZSDDPW/vnFEuQ0maPvkuIXVtBnMUBl
DLTZ/TXae4T/ZNI3REQmTbRxoo+/GlfGmWqNeL5ZKtynSHHd6FxCLCoR24vjUtX+
8P73XQiaspgxicHv3GVGPsSKcp5NpMhkEUgtjkhn0xzwPvezK9f4wXd3TAfTaK5z
v/4bQR/HE2IOk97f7nDAylBalZ9oYo0JmItsoPaCsE96tCCsr+k65A1lzX5UUdal
VU18zTIVn48rrU8H+gFH/A0NskScH3K1hDK/iIQG0o814gTrLt3NRjla0cVOfit8
8jKJacYMSm8FhNqoX9S+IN+TnnepB9Kz2HFO9KFKwKiyrPgnC6XCcIiUFmU6Xg0x
Zbn7h/Mn59BD16mk5D9ooIbuvUhpKnVtRogc32hGKkEeXo7ZlZ8K0aUCAuWE2Z/E
c3fouY7pHuBZ0PVbjYDpNZzv6qIZm35EzIMCLf9NPXncVkHN62D8Agxa3Zchw4ek
w03xSDaay+VebvVl/qONotwHbx4vtI1YJ+fkqDd3ZgfYyQ6+UhDx8qk6jmmFrSW5
DuBdKCZze5hrTr7fQ3POzBvPipt1ZvpoOesXobUSBp5Ky6m4o3c7jpgIo3gXfEjR
HwWp0jYyN1Q9o0FqIpMC119DEkNHM3VoL4qbMEKKuUrE1UhO2IuRoQLAQPRNcQWQ
812FTZNVhjj7UqnpH+YmORwdpH4sNBveBd7+dupoWJ27F/98UXN4KrK6qpFCFtOn
LmUXu7G9u4xlKNBz3AG/JlM+MMTvY+DlPCBLZnvYEvhogvFIBYU5/KOnr0pIonrD
eK/6GgzlvB3H0yBM2mukh4zs//MSh9+n5xpfKNKJaYIodqzS+2YDcMSE5pOsvi3P
gzQJh+8hbKbomP+gHY26A/xJuRvL+Re2gKxXFTadsVWmczN07UZmybRCdOcqKNY1
MbwIVCGJphYgRF0W//K5HzCIVKu1pYNc/tXXW2QsyMUfrLk7lk3zDWRdz9u5cry1
6tatkDP4ie2qMwRmDimhOG6XMnPTt0Q56CPBgOVT1Opfp2aUSGTqZSVWYJ+GCf1j
IxY9NuE1UjejgGpIISRkDaNhv9u0ixwSJeXvTRqwBRcPcUyjMDuu2qvHNxpKGRjl
MducQF8fXDV4lymV1svFKk378/T5w+7jv/uVBZoTz2tK2HIcGCd/QefyEyT+Mih2
kUrHdAdRHs66uyMVg8uQXA9bymyYc07vtUMAD92qLHn5Y2CAmzPAF3knkHskTmf9
XdeVhb7+rbpTzfQJbJU8AtjZd3S/yDmlrw1sNVyKKYpE6S6ZQaGgW+ORY5NeEBAe
BqjlV7ucmlao4ATxfkbf678j8dvCpEFepSvEzrUvPAdfnTXgCaH4KCFaBjPbeNRU
XWmX8vSVE7RwInyPtoieZNXtezy/lKlXg3DTGe4t10hbYlSAoV4ic46E7fQ08rI/
mLeM0KhkdqahllbQxVZEB2AtizzrkLWiXkkMfXOSIwZwuohagJ1/fs8rvkENd/iX
r4aGg+/rPbaYrJx9uuEEvRc7nwvDowlvcSr45GAdhg17ic6uFuyG1yWqzVpuRNrI
QtZfmEO9m9LYGkUYntWDbbxcJu8v9WjjyUSuY8m2NRGOMJAGsb6dPHoEmUQLlUmk
eOmrQEXY8WNoM5kMSwPltvKySCjYB9oZcPs5+z4ZDKJ3z+gDMrddNRPb7Gof+RvN
Lzqvcp6VWN9vNQHGdzOBelMEWgW+udcF1upEyq/mqvJQazKfGM68yzWEcS0cWqv6
iQysBl8ULZxfArxFBtfHm4EJPbudWZQ0/wdrlUOLd2H8WpEEa2up0ZaHdg2JYzzo
Q8rSIG9lZsjtcLvyGTR9QLRv2NYcc7oHnbst+KBpWXgJ9XJiMwcIgmxlvQs1WRoh
SeTf4/zMilj/IZXjThRIY28mrnGfH4gq3Pa5iCS5tvjdJLNTbJBmEcyYgf2h2iZb
n6eJNtcJTHoV+io31MQccqpvwyJAMpjIq8i3m8tmFtjUijX4j/nt/lgR2ETlVtM5
O4JYZt5D8t6UCAyWZ4cWzzzNw4KsR3dPQi4flp6Eck2wdXr73nNxhlPFYzgbIaPJ
olg0tWGuTUB+h2Oo+Rxkksu3f8ei6Wkmj9bGHwGsGF+is8ktUWbBg2Dr5O1v7Ak2
2hKRCwv1Sl2qlVhw7ociT5+WIkFLpRQWX8vPoPJ2OQoeGkibQ1uEt39EwSHPfGp6
fGadYOZcDF+/ZTR14OlVbPS2MNPjqgBeL+V3cdL3PmbRRe1FUvwCZkmclXH6p/zT
To8luQYFUKUFF0sf/Ot7gHZqqAjBJhF7cdHfnewBCx6Bpbtk1jRAUQi+d0qJe+q6
oMUnEKc0KV8toVYbiJ1spTEzBFlKr/xJVuFYVUC7Qr7qUH5IKMCE9jlCqXBC1PTk
9X+WFBPcqE/cC+RFnyoTyA+KdW3ZJdBzRC8XbFVUfPZ0fDv4SCNzZV0y4a0+DxO2
RHQMVs9v154I7hi9q+IjN906fq7Nkn6oxd/qTrWgOYwPzW5MS3GjmME0ju0ojqyM
OnAfxKeup2YjykHjrTZ052a1L7GfybpknSZZBC5Pq734tu4CgnCTFQd0H/PYFiRg
I2X2yBdwa9uAyQTKt4FXaofKWiqViidt5ARrwMInOvWmcmcnT667qCk9cvHYBlfw
KMHPaKMlNmgudnnivb5h3yzem9wNGrBcbwTQHy9C5tNkjVt0c5IAcPNuQwFimEn5
JJ8WzhmDn7CZ4D8hGIk7StxajBhT/7x7PTCi1A0PSRhsAdrPzo5vQ6rD0stw3rV8
EJ1KFuQMU0J9TbQSaX4CORfEBHqnaCGldizLn6A5xjL5iszEHZyGutl8+Vqjjfvm
6MsmMwFHNgmX3XeDZjG12a4oNDagkaUFxWYeHEqcT1qkSH1UEcczHfecpKBKJbwF
ztmm8Rbdh5MBPqhBBv2VfOh9wbn31lyYt2kyWVYe60mm6pmAhxTlJpdN8v7REVQt
+jOsErZnQTF0OrtFBo7v1+YEyZyTniUtg08C65+YLi6/586uznaUmZWo4kLJFO8J
JzwGbZ/5rPqCCWErkAi2BI9EcTjC84gNnMB3RCWRFZPf1FLhL1/3nfQ7Gd7ZnHB7
Bb/xRZQTpllGsfiUQwNJlfMj/Q2lmzKL1KPZhspgIS6QQ+jSoV6fMGhtnpMUDw8G
YHHxPR5T+zs8EpwBr6N5/3Rh145+mZSwi9tdqEJz8T+sCaSYf3ZqaAek2WOorPmU
/f7eFTlcXPozGIxaQTecG64t/pDlp3SdsVLXUixkggPPdUqCbFBTmR6NdHRlFgfK
ochGWI2+bj9DMuwxzDDjo1Vr1J7MvhIxYEZYcjPH0+eSWjOPAm1500+QDrdnE2Qh
5eTPqYTne7o+pcJLceM31AEwwHqqj6OH0YjnxiXM9/68CS1Dxob2i68LAQW7y+DV
USB3oqy+C6WxU/hibm3TBzuqBVK9PayYkQCNTlVbd+4hgPfKjxF8S6BlshycybPI
VA+JDMlDhocWhefx69ZXO5RYg06HtXBPyJtixaD7KCgwK9DCKv/b6qQdbHXGTE0a
0PhwAv5U7QvQm9AICiYwJwftdx8Zg85Hp9VSye1Pc/7kvEVFgRkifDCeAR8ASD15
KikamHjxCR85D6pcHPbbDyhWXQE4NtmpWDp4cDcysbgVCeMFmrDsw7SYqgykIv4T
OFQH/8sQxHhLGJ5/1EkESXkHsr2vHahx0werqg59JHwmWd1L8wkFZG+yHuKnjGLx
GyHaP2CkZfXTC8a3Av1n5rYIzvt+GqbrDhtE4/Hx7NWlzvj9HsEnVRHdHPcW/XZC
LrKxLb1dJxfXhHsUAGtJAhPhVmitDY4OiyrAkSNADWaLkQP3IPso6di/AHrsoMTH
wA28NjWlyuKG27dWGzjjaoMfFsRJa3b2TR7ADhNwaiZO4yRiP8H7HmdWmnZZfSdr
9KIpIdXg3Fecn/Nwl4ybJm8hDG6PfQSZpZ6WWyyTa1Z9oX/asPGLwC6S1SsH1f4m
+D8xW++VuZJhp/LlSz9wYp7WjfyMyEu+QAaQwt13djswUA2Zg36EPhxl+Vz9wCVU
i4qoFPwcvcqCLgwkQJkgXpS3bjvtvCUJ3S+l/0XprxIfPgY/zWyYe600x3RqgaOg
CHxoqfqeUuUHW721t4i8y6wT8AlV3L5cPOgUO0L6+PkHgFUNUIr+LSZRbfyc1tNo
64RbISjILHg0+5HIXxRFtafUE8rOeFc5r+SEl7lTUdeApxTZc2AsQOehggCXFAHX
Cmo4xRxIZ8VwLrY20NNKLCMgEz9ASajVuhkP7XHjYeDdJbPLwp8Cqg4xb/oqNfkS
lTm519wCfPsRRUknsZUc9okGRQ3bij0oz7izVUVySrLmVX9N2Ma/y78o16qt2fL7
Wpic4dVvYvqIGVBXkz6f5eyLbXwQb4eT7PXBkeVXI+Ss+eg+NlxaurRMlFCH5sVE
6oa11JWZ+IC/ixkRbiRjRmZh0jQhAnx/lzRXIXz9rOZtMqULrXzEB3raoXLcMVGT
AggIK817KuG7uo36DBnYBCFmQBJgHaPtXAIOOMuSoekO3moEy2LnYAbWXIgBU496
Kj5qx6unoMmdYtvc8lbIaG42eVm2pHp4PR8dxUqiwLJhOhoZ0yYZBirWzWk3YYKt
yWha73nJfB5DruORqhjVx/6ZTKqrusMNbzqydA6/hewOEHODfN6O2jeb7BtoJ0+m
O3kRJrlyiIfVhh+wfgvzcoS/WMkyV9s0fecPEegB4IpmUYBB/CyO/1NW8Xh73NS9
AZQFbZV48EQzxQS2lrlL1WepZXPmaAz8aVljhWiFt0qT/8xmeCqsB3HEXMphpkD3
tih8DgkbnHO7ODkXklrHtdtxoIPNr9WWnHN8CF+6Jp+tQLWaiLTJyDBZ0QuQxLPi
JVp7jyn5Jn6HuMdb/Lxd3xjH3PrZBeYRHV5dsbJj8rIGpmnI/YVrLpGVcOWYezNR
lowzKFCmqri+MpKqNszHZ+8p+q8HNRt7OGfqEEctJKjZY4B5mv8bOmja7jUU3QYE
RxGi6jarOty0m0YSBe6abLS+olJSFJ0NsH0h1Rm/5uB/446iSmLtwLaIpyidgQVN
BVhWCi6GAFg7VNl7kJnAJOLBavuYRDVUwfHRrBltGqlHSitofAxnwbq9F7F3j4U3
kXxKdvOEJBEYfm8hyBGZN0V09OMiaOpCsN30EcspfhQdvDYpiz9gu4WTKdnfIE3M
sL7lruk7TXnR1OWEO7Q8+iUkxq7kll4KaczgUPGgT+5VzXld6KZ+dXYI5nwWki4O
g1cbBfOjWeX4eMtGjOI5d93Et6rUduuXueBFz2hKPPT4cMM2m1c8DssaK214C8o3
g0MTQBcVFgl3gXNYsB24OfHCtQEybMCY07Z7DmmAoz3I1NPvRQm/LYjrv14V/Huw
`pragma protect end_protected
