// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bf/jjClmoB6QrrVEPLpNimpI/GCQhVvVxGFUXUd7ILC1leUCzFZgvA2l13tEkIcG
1en33j/H6RQIppxZYTEykPbEpf3PgE0zWJj1CWHj+FPEz9wDJsCDTBFhM6BqaKf0
q5rNJs+fAitNTgIVapBFRWLsmfLwm/F3tqZrmuqpnrQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10992)
MJTtNFUiXwns99TwPLAOse36Z1pzuXRFLlTI5sNumgvQt8KUrWpTDUsHwDF4l8Dj
2dlOxXo+eAnOkgaiL7fOyjuwbmvcG9i9HGcSS+AxOzVxFVHrOU8hOF26fB32ZLCY
RQRsErjACDg2xlB9pC/l4MPO6J1Ij14kuoEH8RRJwOKbqwPp3gY5sBHiVU9P20aF
qGz0h2Ba53WT5Eiys1efvHRVUnI/09txjsFdhuVrlCMd+oRcOJSWrgcfBOF4xR/2
rbAbYQLtFV7fX43AG1HNIVhFVNkbAf/IqLLDlXKQ+IYnJ0eNGIHObQIivLUR2Fgo
42LMBGe+rgUltKwOrlmQjPXanRP139sLqYG4SgKfmA2uz52LNgE85K7YQsrDJ/Jk
lT3HbZYgOlj7s2tE8DXATGw2hH5EfMtWzmFU8u4hTLsyCqHra8UVEFw/cSPzqoVZ
9/KorydmtbXVpL9KSUcGGR2RcgzDV7VuwuM/mGrxXp83p/axnZ2pFDKH5RJAVQgM
WdNG+X3SQ07ROTHnNuCYeLwt38esNc406wrH7CKgS4L7fkVI4MbHcYvliCL6Ob7R
93V2HB5Mfrhq4Jv9pvMBj5bdOv6QFSMXhNb1YemGMYgZVMe6MsXSEUP7lFnOgdq0
Z+Ln4wt9keSXp/aQb3svylsFNaCQYZHRET2r7OBZJVFGPK3sWp9gbqcKWcp1fYqT
es8h+qTaGCI8JdrOnvMv/tKFSG9nv85iynh8dwdL7fcAC1Ul3qjUaz8WxqZxqO/x
15ONhXF+DZTRH5GmJ2G2ZhiKAagkIpZr8wawmfBGeA3v6dI61SYzy8D91vlYduJ2
yw5ynHkXHCMJdnYPp+cwI4MeqETXy2HU44JxhCW9WR/xcwsXCKAOZUKGWLN16pLZ
wOFB3uGnDMLUNtC+/pJnCvzi/aKNt/1FJGjdo4Hz932yC0qnsbA4/MG69bvluAYG
eumUE0ynvF5NQCVJua4dFnrCXHlNXNXtcjaEuRFTgCC9rYU0NtUuCHv04IqO4YqZ
RYqv2u62YKPhFey7Vu7qCXt1CjhzTji11dBPfh6DifcWl8Wopr6TEvuFkK72QAII
9+6E2BaNklWNI895rnrMgQAzmYHEIz9kr7LKUOQvshHylJpxRYBmVCXWq/1uiER0
OI6RT8oLOMW0IywPB2X1kzgjYjHLma4AIdXnvKPtIpLa3tNk5jKAEgATIu/Yv+kJ
6Prkx6YfiM0IqTH4KmdMe5DQdSTGarZp50jxdhs4pfsEsG9AcephSgow+WKPaYM7
vETo93OZRZuuxxKB0gasyxE2Bs2WWer+8KL/lm3+sN63ODcfY/WLixCqi2ynUkAJ
cgyJ/t3hLNRagWjjNfgsDFDkq5D0aKIb/9IO/9tTMidZNXULOteJKFNdIGOkhIW1
nmmH94148/VYvYbv9AFIXL9IvtNsE//EpMm3X8gb/NAWKotAOsHOr4s/0jm9VZFi
r7j80uNhdPi0gRRMRmXpSO0TUG9ESpzIrRb4ecyzZxMNYd0q0I0lu1xLJSpxMd2U
h6GQm0y4khoZ7XHpkU3wo7XMQLqIZQHj+qtVR/9tUep15Q94FYwDLyu+EXVMH63N
Yev54zBzkEBVIzpZurb2M00NZYwNa4Oal1ShMCWuPFKgsho47zQr7GxTdE+bbRRp
HReFg10es46UnyJagkPQCsEmjpzU8+kirUF1ZF/ws1Ent+eM9J+BK9/orBUm77wN
0/skWUUOnkQwejBG0JIyo8RecyIIb+OS6GFuE9OK5AZBKJsZkqjeCTK8bZo/csgl
h5XV9jaidgvqX6Y3hdnV4wUFjKKmiaTTDuitukTwLlFFVSaIcNugTeTd6I2Ef/nB
7uxdzfwQLS/L2NDj7DHk22lC6O73Msh9c9Ae23r6a9usyZPMzg+PtFUqwpIqWYIp
hOaS09U24r200lqaKfzlPvxDmUdbo/SQDeIJ2aSpCw4K6D7NTjkz3zp7vSsPch5N
mR7Ayr9lvwaEWAUqUP7a1PquNHF8h/V5997YEQksf3m8mrx810+fQ3Q+HLzqtq/z
E5rXKKQfBbkK0xDxvMBQSVOGqMqWjhDga+sysmyg5xS4wB7c7Nzg3lB+/4D2fgyp
x5OoM/fw4tIlBZQPHyjJxuEqvdo+HHDie5//NrNJVW80fdyK9afG9a1a+su2JRst
t6El0IOVqGk1S7mHhNo1tE5k3+d15EXb+L/NLAswX50v/QMTmF9QJqfh90UM2A3T
U6gKcFAqJW+a81NVPDOSTknknFta/ZrQxMzdtrGJewhcvPQURXJkEm7LWlq8M4M9
CeMWwrTX8A7CxrwK5r+L4ZY1ep1Jel9V3gI71eJo6S+AFSJNnHo7rQlsIR/AAzA2
xYS6Wo+jMbfrUJtuUWQTz8go1Y+FozkkwYQFz+tIqzIlIGclU3eKa75j8r956sms
KDnWt7cfjPLWvk4tidmSqTTvIKiMHGIT0VPUYKxnO8KWQaBEu2tYcb1vfxQYxqH5
8fbu2N6BpwwkmE+k61L2l+WKbI3X9ruCM8l+1OUQZJwHqKS3va2aCbxyAPkYuUeK
iamF0hq7AyM1uJrwItVR0KxerNiatiYYLjgbjNzEpuQhwStIBRWnDHeN9uYbsp0L
Lfg1gcYJpE6853ZSezexJEE2hketz+MSYhCLafFhRbAQP2yv4GL1zqMWEYipsqxg
ggJHTrKEjut3C3Gh+NucqKk2uW+F9VDmLJQU7Xd3gkVyUtOxkHVAf9HFeqbOCNvn
pqNfIfe8lMlsplYGQEMUpx/61gQdALj32l2Kwy7rFHTiyQN7AE7bcvnHcXM8T6Sr
MXCIo5yhj4NkCWGwg+V5Rf0vDVIxgKsrjLt0Iq3LsKzicj98euqNSRmXA21r2sj0
s69lR0I3SQdZREDKa9AOIYdOsLXjL4eqdveCgBjkbIyUSqxdhvsRQE6YfcOOg0U/
n+IJDsFD/ZMViRRSivcato/8C4yd+z07vj6So2mVjUGQ+hqOCHxDGi2kV0jmIfah
lhy4F0Khvzag3VRPuItfZq5kf+1r7sjWAvncWa7aiHaF6L4BUMFumKsI4Y6GrgH2
ikjQ2pRUaV8TW93Fjz3oJSWS9YBLpitcjg9DVizM1hH9gBM6+1xWmDfT68LOP8HN
j3o1HoHRQfe01k8Q5MslbHxka9ne45AqBFO6/m2zylz8/1h63rYX+zmBDrB+Ombk
0n+tFbz4/CON0JSP5e/0SxFVj1Qxi/ZITWMM0cdm4EXm+UOoYZsQPVt7auZWJzNf
3xzgKt+wgGIR4UK6ENOeRqV3AgSE6iSffHm3SZkNcOvgULMp1fulAnGsu0tJkN06
ZRYtm3mJ0S72mWHMgtVhQ5EERBFCYUjakBWsv6z47lC9Vqo2H3rpEDbHHQJMxfKf
qtxLnpyhjEFAIOZg5fpXlmqsdQhZ9DIQWlLYOeRCpRIzZMNb3DM7hdcCJEKSkXM9
xkXWMUfMxz6tk++wu1tpIi7ZV19Z+OZl70bdQhFQnMtKt3d6ViCBp7ZSDqAi/WQt
4jYD1O+CtnLkBIW1lzGSoGovSbWSavrmQtffYwpZ5Z3JztZreL2g88VAtDT1hxYt
+HD7gl6wNBsorBwNxVjmE8/xEq8KSCj4C8q3Nfb1ZypF6Q7gckcdXDlYi/8gg/Sa
ouXQ+4jhL5H6L7xBXy5siCeKa5ItmwYLs+vfadqtdPXMFHa2BVha5rGbS5MeCVK3
a7+vcV4WRXNST3xQnYsJ000vNYD6hSudS7UTAXbSlJJLiN1iDn7bfJvaYGgsRili
bvTS5QPu1+BL1tIwC2PXX6XR8k0UJFIIBmDbwei1uyzXktvfqPIR/KU+KaxuRiTg
r3i9KpQtEpjOkR5COXvAOMMmvI1mL9f6zTZThf/u1HH6PFUHLtpAP8z1eQxBlnnz
SZ9auAcdEZPLMTDb35rkhGVEbJxQV0ajIPHskAPLyTHjxIkjDrwg9Mgp7CnuECqp
gquIlgi+OzChm0dd7sl1UmzqphsgGRXZZAy5/0CHiEff8n2zN8qF7Q+HuH2WjD7B
opDo8aC08+XLMd48l19HO2/kXVJkUD3VhrEpeX+AYAX2LPaBb9VLJ8zdTkAKeMIB
GtvC7bgQbaB9EwQ8ywK8CWgTowEX7sP6hXjZxqD46XLy89Bsp9Fyu+V8jGC3rzEC
QpGd58JsmWmvXGURbsF9tK6C19p1G86joMzaAIPWUdRiOvdhgRxRHvGV3sz8ATv1
p8MWdPxP3ZbjOmqmUkcGhHvJh0DpMRp81aXb9ZbAktyRE23uurpikP47b5TZVIgg
CcUYUPSQrH2z5UXXvLutCI4zE9XcjRVdAB+p30H82ZlPzYPt+sTQ7+18mUQXUcKL
IsnpoejZVsLA/LgdhqpdJi9XP/5hxJEkEPhzjbXvUdXQs/craeyLsJWbupTRiIAE
io5IqE2hU5X/f7QTzlMf/mOFe/9uWtd4mxtTXs0fmlxDgUSf5V4TawTWx21vLbfo
bOpjbwUsuTtQS2FrHzphsK+P/Hcr2Z63SKtcP4OsVaPvA+98TmgY7+r6NoatGWlF
5N1bPcO62WbGpTBiqiLmj97nPRizObQqIzdOEqPw0IBQbIishtgNvu5SHGdcTV5t
eoFLVHIPnjKPujTwmtbe9XgCSbx88rJfte0QjXDSdUdPMO+RQGpDNctLM8h3mrO1
mlaDE69zmYAMyp6fc7II7x13x8apWGa8hMyThe66XT07HfRghuxlzXMc8NYctpIV
7INLhwmPo2kMdPB1DAdKRR6Lzy1mF1Q1DESMY3pGEGljoVhR+HWBQmjNKUqencr+
xrAF+UZ24jr5g9SmXzdvuJur6RHXmnSdxS8mBbfUAdJSvJyH5tzFbukfGOdqDiFt
eW/vIXOZC2GD+eTWF+foddmd4KvjHezw0A2Y2m5Fl+FgYkEqONj7Xb1qsNHQ1775
0Z3wiY72tMXI0d6kqaOJTAwhlr19yZkWiQiI4BqHB1m3KHkbQgX62zZpSzveVPZc
qYoJzMfS0ohzlg53iKiweqjisJGoTWIX5oOTGO2Gjlb0nIASgmeC07hZ386E8x5w
UBB84ciSBgf5msCbRYz9sox46pyu3P17e+YpHAFZ4hAb31l3afNiLWxAEt2uddBg
DzWVGiL72ZMlg9Cm2ZFhSIF9JVF/dmrJP+hruv7JXM7V8GH+J5YSFoaopDB9FCLq
v4EurYM4luIh5Kx6tZG7sXAXsDdhHnC/Ki8F4VRgCRZHoqO7guXmYDiYYAjwSq/T
cfWgZeu4md4w+RmUBnCnEKLbM8xgmDw7esEM2T5CiZw0lUIN7ueAZX18J79+pw8T
I4s0PHO7LICHDK8yYl0hMliaikYDqlJep9gbCUlcz26T5r+NKXfXEj3cnAvlOt0S
m2FfSaw74jGC/ONl2tpagSDRFym3plHszOmTaPDslkv2pmvGjDPJVonXP9zunXiC
/f4/6RWOCuB2s4Kj+5ke+6L9sHS1DhnpsVMH+AGKcD/HV41xKAc+TqWCtW5Lfr/u
R+DGC4aZ2NDTbFaDeP8C9oP7YdUM+eyOwbF/kJNvG6P+q30zJb2cncMB4Kz+cL/M
OS27lsmkE/du3hNS/9SMsdus1Otvtfn2xkl93qWiKlJiM2ccgVSdVvy35cDeC7yg
cSuKXLfMlcJypUlYCLVTwin/YmTHaNM65TzVXXqEtqlC+B1ZI84sdniqeSuTkvWJ
weqH/hX0O62YRMoJfpIaJOntPhs4xci9YrkAAS2Yw2Zm3Gh+yH1Pbfc23Txenu0H
QPbXSXAqd1t7+vEOkauF/lK2JRSsm7yloXmDRVvFRoTnQL3k5+cYQMttkolZKoJ8
ZqhgZbJxOr4CBNMWto/mWovFIjxu1o7gi8AeeaoTpNr4J+frNjndhyMlNpyoyox1
7gnSzx8EJQPTwnXvK4MDpeVo17U34zTwI28gxbeF4lHH/J27RWdmDHiQuCvYV3ru
okBMgHzRw6EFpdAOAOQgmRZ702NWHEoeQ1Fl7LGWopLMD2E68oZTCDl1rpOo2ALR
lPCaU7SkaK3UDBgIA+KcoAx63pQmAwAqRcWqSVoiBtNKxoi25Wn6vHypbe4d/p/i
OebBMi5UkL/vrf6u6zEHvI6aLRt5EJMiqfJqc+2Y/gIRbQAzDk4f+KMpzVUZaTFo
1M6dHGL6+goAl9hboSrKwDP5WUcWJ6D0ARtndw1hE+4EKp86LhcAYugpa0XkutkO
FdT/XX37jPHEkX6fe+DZfAaIrP5TUruMpJzTaZJAJeNjkw9uTr1JbC5lwcrfVjFP
cqV7lNnrNt5LGwr9kU4S4GBds8xY1Si+wS0Vr9mavMCcnHiuDTKEfH3dM2JmG2Ft
G+x+f0JXqaCTeRbQuLfumueav9wDgxqkpdRojLmWnaKXTbNejYqmZHcaaamA/XQN
TCkeXF5mu9vL0vVQxHM4e3hK4/bV1nPw+G8YtLUZCK6mAvu0wqYNBW2g8rksgMHj
uJQ7j56GHK1wIdEKFg4IfO/4tzCHqkFYy2e+94jtCL8y/EACwUfxzxgjPFUYAHth
cFNKKva+tpqrf2fTJ5lqcS4USxgj35HHKIs2B9IuhlFFwd882R9ynkp85LoyCdAY
+mOO+fFn8g1naWH33dLgxbq0eJVDQgV4TUiD9QrCyHHrX+/IDjLUvMawuz7EEnKc
XiSCdNehqPV0T1QaaGJTq8db+nFesblACa/dtYM6Qwf63Y6iXy8l2nz6rotKgbtD
vHyZkKPn328PHkV6kuUzQ0t3a1FPDwbaezWaON7P3IavsTu3PQDojHXnr2iHlRBh
ID7oHBw5CCOfnzMcZQ0EqpqiZ6jhrGvb4/i39QnXhlsFYy0WZBofbK0EUPxM5b6i
8QmlCynwI7IcbEGNWQHUaykphpaUidIbBZ4RLvihhptCPc4yaXQqWoTgtMzfhOgb
1AXoZcblo/YjUVdqUvw7b6oAb5e8AkmI8B/9c87xhKZk6yFxzuneRSbPISWPzXxO
7stpio6ZuQNawUKGeFmIZ3jrMtcSLF++RI6lw0cNy+Ro1/cxyB2Rzc2c6st/OgEN
wfrMoqBFZJNL4kiiCX13W1KngmqmJv6JZotF3X4JAQXNFPsidAD3Wv+JWrA05T7D
ACeUJWYJ7HMrXXTwOp9di9vzHMtiVJgTGCyudXnHzXOWQmaLIxHJJwC83RGQ4Mbf
4XFPvJUyvjeR6zDoX7AdUt7rfSG5pzat7pv1jAz5GyQfzJOWjo+vz7Db5rgEHGI+
2qeN2XWZI4C69u5U5xTa6CTnedwkgkz4v+VMbigY8ohS01Xj4rDK3Kd3vi2gWhxh
Zj/vPbJjBLsvCVqaDfiOmcbqmH/UgSKspxYmfhBCIYPiQzmdtCACQGVK4+e79S4U
CgLMPN4qRVpisoJTULi2CyMlE6wvwX1oDSQpO6ftJ01x13AiauvJquLz2JZBhxpH
6+oFYc08eZdCIMLxX1rOYjPg9FEvsvmW6XhEBWKnA0TqCkYeqVR0+M+vb2oxJpnV
Scm9xeR0siOgLXnyyHEIUh9tGQKOqWDCxBvF87QSkxHMAca5mOw8Bj1h0yqDxxG1
3jhFSpXDUQjewLTfgF4LFrFuvVbUbUovWcwsxz9bokJa9fY5zSGslyls+NxcwtGt
PGSk6AfJVLF0dPeZ6cokz93SbvyRV49Aa5EGrO9b10eRKNDKErQ+euTUWeMS/z9N
cp1VSWKbsatXacqzjRHYx9HjbexwlOOz0eUgjOtcov292XVPU7dUXsbgS3jkss/6
zqXpq4FI1b8T05Ed2JPvuCLVe3ZLTsT6QxYZkfAdaX8Mbwh4dF8i/pkzXQdvv7pE
Lv8NRwjwPsrz/aPRWn6BWLrs7w3ezVOFDeYKwcPdOXcG7z+A0zrqa5W69qibElIf
RYrZOee4hf+8j8+/fG+Caqt/LplxhGOUeXjuar+ig3JIjGdvdPj/odmmt+WTkoIN
pIjvCKGmFUaOX4+9Iyi7+cAaGmmUwyqW/0TYcVzps60sRCBriVdJVja4TGaWGNkE
osT6t8X6JhU8su2FQ8SoT0JD61Wc/404EYdxpnMbo2fShmeQBPkNqigAev2W6eDG
4Tvo2uulN/EK1/LepFdNNZeZfOwwWEqOBqb2SKvIfQwxckWfSDZEz8IKk+0UI1fk
h9ihmNg4XaXF6BEvZYhsoZFMqaeTkox1yhqhucKjJ+HIxrhN5fQhqFCdYomPsL6Q
Cv8zhqnTxXM8LneQuhCZEKOGH+LWaNg+lgEY3Iye7uaAnnqxvhYPm+ZQiTdbGRjp
cU9cf6gd+yZioOYwr9HZpebxYqh/hbrQgub10gPQYMfX5ROlaaCJoe4ABjY0aHTi
xf8LXvpqC/LQq8TxHdhf304gQ90R3c3yP1IM/Xmw7ylyQtzJCC6Ej8yIZL/b0rTz
T7KH2xZEU2f6S9eTmj2Jt2b/4yYJzxKI9QK/kIMYJjeuXgdHqBPq8N4gb+BreRHR
80r0p36mBRMTFV56TyzEwJiK0Yy5wX1LIFMvLOGVETWGJPvmbNlflBUHk30vmOFG
mA9dY+T4kvLymB7Sf7mBWxA8AJ6jW263WlYOfYyytuDgE7e6Xo6Ok2yja2buA64v
C8NicnI6Rfet07w7zsapFVsLY+BhtiBEEqBl+k+CsCc5K/c8Vs6RMSgrgcJTtccn
KTVpBRzfMzY0W9dVCfwq5QBGhSbNfFBAYJcyGATSzgmZDEgsXUtD1ghm4QOIZIhH
MYeReHRIF9/hR3JoofKE51yUdshoOU9qw6llruLlvwzFgSb4IDaPnE8XQ+3gAFoE
rzIxUEtK/cmFpy1UW1Xam8BcjZDyo9Hlae9jBQiliHKwyyfI4sQyLZ6ynbm+aVKx
RIYq0XXJd0kLNdGBYNFeM4AkKiSffpcknn4WGiRRLvk/BgCVbOLPnhuo801zobB/
mr5zkYR63b80AdV1+QK8+mv7Ch5NeJVgcbYp8Dx+jUgWItcI+e9zmZ4mGEz1aUCT
CgkEj8KU24PBg2K3qi0h3x1PIMml8YZO/jm1UheJu55GGDTpZaeTVY8Q2qQykgcH
O0PqSP3kzH5b4jT53z1tBzwPGGflXbPJCAcSUqlWXtUjLkB95n8MN5ejKVfyf9OW
G4BMMry3dWUs7FcfF2ESDlG6BI8a3DVH7gUhMG/t+W1Sgt7QhIJYwu2pkVOAq2uq
jTAemsHUQRNc3PC8u1EO1jhs5ROTiv7/RUl7RxcVYO7YzI31Lkh2GfdsGtYQ9nhg
23NsRj1xa4hyVRibM1SEisMzlDH6a4cyetCj+yei0pvqsCeL44ncL+CmOwTq15F2
BAnmJt2BcJqPVQQyyrzJGBTAdDZf7PjlXtEaobGqUD8egHNxJksaHZgw4wfitQTy
NXufscZeaPzHn0aYcjuY0HhAWMvxE21YJ2dsdXRc3bmVETD8YDzYANZtImZX45rj
B5ZfVniKr7oJYuCdobUWTciM8WNzRDf0fYDJd22t4xmJaS2sHFQR+EUfuzjDmrsG
CvwpwTbWO1l2w8fZzQXtMm9bcQ3ehFuwBYBPjSLed0TQIqzpFK9UaNfLv3dEkS4R
wkm/N6ZhUJlpE5awDY+MKmCRGQbgmwC7UYbt5ZOdrgaPvxyyDiH/ch8te/CWeJtq
aCTyQdPNut8r46ajtzfc8zx09g+Vw3ccl3gtlddapUa4Sx/omPgWqUkJ0sagg2za
S0dqR5sB546dElXARQ5O7ByVjIFvBn+8w2exC7U3cNo17Hz5efY3lYb9TDfMPtjW
tgFAkdd/GdSvRFnDPWaJWVsdzkaaWA9GML18n2Dhq4XHoYV6aJj0gYWXCs7WwQlz
FlMAmricVrYpfwgJOMl9xv02S6aPV2op7MM0ide/+uadrH2ijKMQK7KeOTYh+FIF
SDXkhJdYwN4uaWzFSdSeb0TPj2m09vFLPO9dbeIAa1tluriG12ypAc8x71GAJ1B4
W20JcQD783CSP1qBrGld/rsv/A0rmClQvo7yn64xFYtx9Izg1hpUTwyaVbPFck+S
zFnptVYaB+Gmm7Ziu3n1XV4k5Qdt/E6x1LRV0G9sGgq15OyeRkurGplZIcOYn96h
IRTmwe5P7sg0+38Rv8qT1+nJ4mFc8idccmJc32hpwWagyS2xYfS6EaFUqR7xcHIP
7WpNth0yQa/w0Be5qkeWDsBGBy51XB3pZTnIeIcZ9x6qm7aLFsdeg7R2cH2xubjb
PNR4kskT+dApLPysqbKWg+ucNcaYvy5pabb+VZ2jzZOiDvDiAEoGQCOfHwfmdh0W
0/+c/gozMmYxGh/uMiIe4nIIX4ml4OB4GrfXMDG/aUWc6MhLTvrK4gSVVWZFRJXs
V4zDrTbe3RArlOnstzR+3KtOmMh/dPPD0Ta0Aorpy8oJBRtvu33Sbr0dLmHWrFTD
0B97Dl50mohaHVnqHVOWehdKyRj8fIQI+wsn5KYUr3pwjCsFU3kD7rk8f7ODDqod
ANG+hvPwwZvTm+C5AlO3jakL/pWMTiqhEc2/WxBSgrUEh2G6cylsAPawJRpEf6UO
rtAgZT4wUAm4pVTy/udkzOEhwx7kBU4enpV4iOuX0YM/XlnvNfNJD86ybZz/rEKO
J+3tXxe82gU/xWH8WUZ+7nLFWLBJ9uCNXH/Z7ZLrP0ndm6TNp1qHQO8qM/+NG9A6
ibyGefW6oK0Lp2mm1TljeFkKOcCR1gwnZE02P2h2eCcWZ4l3CEpBzDejx/x/Vfwz
5cfqAggwb/bsfGN0s1FmZ0CI4ae/oaHLkOUg2K19Pzxa/UFxXMADtZzUzemGsGKs
63fmhBVHqMhMm/G+sFc3qqJjtmMbHZLoNmMqzzT1eQaTsM/6nVs9DlJBtCzBNQe8
bJZlGmVYTC57fXoq0YhUbszlPYT0suA9NjjGB2F3/KiHd8+FZWLZyWvOENaW20qy
JWHrMtuV8HMLPQPShyNVWcWRwP9wU/C9rWAU0BpCMwDOFa1qxgWh6o6awLwR7EAd
cqnB/q1nhoG1Hm8Mu/kc6mRwNI9RY599sSwWRhv3vb01lhFGVydpuupDAL16Qksd
QCKISfWtvQh0Mvg9koOBauz5WtAzlAsDT5CSiSRLsHmJmXut4zZDYLxaRZDl7Kpb
BGfEL+jsfmzuvTyPPPNp2s569LW5SvY3FfeGHL5fEQZ6TBXtNIOQkOm0k5f7ix9k
UdY6S1/PipHT/jEJzt5ASm6hUbIPh+CpLD0bKOKjUKGKYs+x6d95PAB1UpZD9zSR
LOV3nZRZvTWDR9hDrbfrsx3tr3XLct+xNyNtYcOLj1LoUXO8vmDbyUwuFtJV1yYH
SzCXU1nadFXcKlKqdOOpURVfiNoUp6dmvDOyBsJ4u4eLMZYXzs1zqfkBMcF58LuT
Bh9rdxNAoX7SxlqlpfLHdJyAJLRuEhPsgitBmQNOZLkTGCIVFOpolz2Ina8W2XYF
424V2ndQRWYKUKjg8wLxOPQmeuj1bmHh1wscnhwgpazxQr8Cb44ZLuKdZb2KT870
9bBjsCDNM7ilzNPESqaz1TLmmYCi+izJg02ilCH8u8sc/GkFwG8pi5PH82uzUJ+/
kK0y4dYOuDt1oUEAG4dtVrWhED/OKcv3sWFa52/wxsBbJJ2q+4PhGumnM9gQ0Fpe
0uOqEjxYSbB852E84YTlnA2qfP/T6J1mxesh7hQUuSlBuxhZppjRUTlwQEPJIL5v
gbFEL7gnfEdCf+hCOFM42e+QhQkNViZ3eEtUy5IgFotpNqD3pn+4NuD/zg0hPEGv
d/kUy01p4n6RqmK/wxtEvXLBOrA91dYN6gIKtvMqiQmdeBvvFiokV8iEqlI+vPQz
1cg8y8hnziCwkluIHE5Pl2J9niiqddaXdU3n+EMfAHa3gcHJUAMx6IPV5XYQbmPK
b68Myk9PM4785DyH3WyvAdKZH80l4xLoRc9rfw6wJdhvhXGCjmZrsCCLMztEGErF
gTvPDdsi5gujXmkQ6joTy4cRKP8MvXqidgHS9Jk76A8LFHX4WrP96NkR1JNBUR7u
DfwLvXq/4pZAbw3R8rvMqyzqbchsWv+2PQq0hvbdH6Q5K4vNLM2qFqiYC+/sGR4S
Q3X2blN0hOjKgMElmVZWxHlekyS4wqw65NogstmiZ+VQLgWiF+WDDQhPyV+t0C5c
qgwEJSYc2aahXWjDcNZKt9sYef4tqsN6yYbIbdA3Fg6OEgfR7tWlRrTIu9EasfJj
yltbBr72DRqPT7eb6aCrMDg7OcTf1I1Li3tLf0a4YasshKJHyCnVl1j2i0zJfW/b
KH7C3foJyEaKza/WLQF4HEzA4lfEOe2xBWz7nt/Nv1MqWkbj5Ytb9eox4eBsIpld
iPSm4AUsJD7pmBCEza3kEhsB/Aqg6XklbQlsnjPleHfUDqjYLBep9IScek/I/UV2
JK9hHgW+0f5tsGbuNeQwJym6sLHA83xAfkJwWqaSuBgOoLmm4esGqwwo+XmIJIre
bmOginwF9/j/rYZ6gg6Vgw986p+BUVuUs8av+7EYPRrYBPfJCMZU8j1hxIpH1N+3
wHL+hlLztKCwbiMBzcJxfY6PAFyHRxu0untsXPVbjQxuB+2r0L2ZUmHgBMNsdWF3
6v6sT+yfXh1Y94SGcW5Rq2VOFXuXhwFhIRmZAi21ibpPOxFgZQylGKxkvt15zk1W
c+qAFJIoxHvsFiWjQd7TG3SV8806hC2B1V88I2tSjanRAC+KCQsib+jtJ+bhgZmi
T4E1L1SmgO/Yc64f24lfxNmOx4j/xgrew5lXnTqn96jS+kVTUJAb5a1RTGP9xph3
u2CK5hWDWtRdSu/CmWo+tpvDLBTDyt4ZaEiXXg4p5qCaDC+PbPwbeLco6AurVX0n
HJv5zNydhmVBnQRSUGg/GTCPIeTJz6ToVDVEZelGmnvCPJ2Gs/Uxwzc+tt5gsUfJ
e/fsFEhfqyzxlPJ4Gvu39FR/MMx2JljBhKegSxbUq3CHf2csIDohwiXo4q4prEcC
oX7PhTv9t608XFAQO1VXjg5RTtxb2wnqlW5/0bX++PGVFal7vN8sL/vhRxGKpobV
x6aSmZru72NpJy1Ag6P3IXr42BkqsKWJzicQlMz+y0fx/LSac7ab83NBTpVnaFWu
KMSK+iG1jltawGhdbC1QfpEWPrZw96yEhQK1UVZ7ZCbJtaCncrL2tesCOAUrgul5
flNy7Nf4At+et+sBQnrS63eFf6JGdxvXM5tb6P6GEVKZsF48fMWwh4q2BAXVoKEH
hXjmX9PyvjJXF9Tv5AH/hKSzF7B17MsNZydd+Zn+7QKndvl0FYvLOPSyvFEcHVNQ
YF2uTkwWlQTXZ+7WaCp0ZGmJ1H1MA21pt7VlpqShcT2dJvOSkMYFaEbVNbqCKSOM
MBp/bh6nWJFpxY4LRB8jVu9OZKoqYNx2h7/kpKmHF22qxtDUkIEGxJKROZ+lZa6R
g9OLxEZGe6ZZYaON3Fj1EwRJVfvj8GqhS69VyadB8Vc1I/bBnhN+/uPawTUI45Qp
y25+WdoY7oc9hJ31GU+kkkzYp6e8qIq4iFgrZ4tmX06xbTL6Ws0x4WigYTIIwZF/
dx5Lu+bjvC0PvSq93x9fXTIu1wTkOhN5bixlmOtND/H3xnvM9Ql7cQLnTehLb50J
sKRM3EpkhHba+CTkxYr8zAPP3WWk4WWEGH2hfD+QDMz9s2cYzuPMMaTxhVsqwLuQ
gv6zRnNt0x8/dPib3dczKdU0eY8QHa4gDZei6r+B/KSAfzrK/dFwhhhl75tyZ3ip
EwAEJ8AUlAhWFnzIrHESYoIkw/amUjlIxyJM6gpN3TNgbmZktLYHBJVdwxAh4wce
DEY8GuGbdyFqFKU+DE8l+FKbnTuBUuOG4SkQmwIht14JegtVSJCYn2g1C07dk+yg
ul7QQIbAYchU1DP21lSoTGryjneT3SiRnjVDWPULsWOQZNsy4g0psCwI6R8drZe3
fPdYGL8m1DUALtRbORjbau0TKZSu0Sb9xHZG5YP0gE4g/a+/n2aKXYQM1KjpLlgl
Q7b3Y6dku9VE7W4qFF+BEIfLOVSqn2auUhHtJ0ueSIsCE5ncTzT9dgSBaRI+Fud9
/0Bo2Na1fJicBCweIuiudsfO2fkTRiDz80zYHDoBIbhaJw3MYyB8/Hi2cQe0M56x
FqssDn7wljTVu2swBm8mBQ963C6sSliLLQ9cPliEQfwpQolAUnhKeOviVd4wvPAF
6zOd3xWvmvoYebXRvSkEnKgoAwQPcQ1ooVIg3tqpY939is4dhkjotm2t2hotkPj1
Z5rA8DyqGRgzYg7ms+B7D/6+X8s2gDJ7QKeCSciCt635INv/aMC4BJfd7xVQRxiQ
vFYKKFtdDG06HFxWwaRF6rbB5xxfNyeNCBV2GRFL3pCdFv6Kv02LFlHcSNlaBr3s
R2x1ssga8DTquc4LfaxJH5QfAhymqkfqox+x6IdCRPJHOImonJpbqOG7oin3CZYR
tQ27BsRaSoDOw8tMiDuyZB3vWkGuXy++Z/SLFOUsRmYMNBqKKSrYX3H0XkU6Zhai
uDnJy8EnXpFgT4as6vbV5WnG0InMeLCtGgnEUT5qLwJNum5ZxocTOhjeZOX5i3cz
sST8NdLpY5K/CwNAKVWDpLo4ERPeRyd4NfNTLBKn7Q68zxke4iWZ4lJRuwcYdF09
cxRoDrjjxcWPGpJ3EPRf92yVNwKWTDNFTrOUSYuBiU6LsyUFmAO377qfAT1t429Z
`pragma protect end_protected
