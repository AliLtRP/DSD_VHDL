// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:27 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BzznR1SK78SeYFQlxzjFSBb6q1A2iRdeZJ+q6vHoidNjuJc96Zdvl2JBUrBL8Q3r
w4MYyPFdtF+5rjSbLKV7cGmnToVA3tj4PXUppNISyPSnLkB+Hbevp+rowBOPIBfy
FU/hNqDl6UPgFDzdB/OlwlUAVaKSz8wM8YAsZBeXSHg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9296)
4Wcue0Il9Dz5OmBB+dzE2kT99hh/fI24BjdDZz9bkDVUO0HWKOPoZrnjAblqc7Ud
LrkZgMYSRDTVzTipXFevz1M8GO+ltXmI1y6VP3Is7xD56Sr7/bUZTF0MzSwU+1v4
wtGP4XWGqk7voyXLdwnMSZXqvb6YiOqEBufq7SLOizIpvjLreXOeoTZtRvnGV288
EZpcHDupiD4XOYd8cc7XIRNFx/iRgKKcpN2gWqmy6Fi4ed13TuotLnF833oA+q9h
0J8zMFvKsFn1TOR2boj7hOnvVjDbRnbmZDjP29RdpIad+QsMYZYdbZ1rpHE046Xt
fftTSGpraeiVz8g4pbVuxro6XypX2wE6396MUh2TbxB4zAhivDcFvxWZdqXUlG7p
d9xhC/TAezfoy/T0OKsFcbp/KlZdkH6p5ow6z3j83c8sYgXgrHtzVAfEuaJN5FIv
uHw011bwKqvSRRKAD4d55i95CFvVwXokGCgAv+NXzXujnOAtnkizwa6D88boDrty
aHvPi7nn5qJEGRs1mwWELiRCzlFjZlaqMpOlBdJ1+BPazRw9knY859UGBMVhKf/a
9SVOpmNeikdxEY7zo1nDSBw6FFp9zz0bqBTFD6Fh7Eq5NYMUqlTjm/Fm+GkVljlQ
YA9lZmo9q70Wz40TEFPxFoySbxz3/J1kkgl1ql6YgrewH5nBGt9HBVtOu6I69B9G
DkZMLjEBPnMoT1p0x1KZ+DNmpkwlp8wVEqh0lGHtqLLMxN0ASex12EUy2Ofn+oqq
QjEdEPy6CuSJs2dND2kcQf86x4XSB3g9b67MXARxu/u1JJysEpQbpTx+/n2jZ3dP
HdHuprFN8PJpDR/Rhto64t1OIXjw/wXTA7h3qNaH2gStvaB1siNCFmvPYWHIKbD5
E1oghhzOpE/Y7wnkxMI7RkHJZeDI0dkmhD60/ZnCyVR5h0Xd8AEvDVG7bMADFroA
SjzNmnltT/lKn8tPbO0YwcG9kytEsKRshCf+BGoTjH6BYlVenW15KMC8zArrPG1g
O0PnbfQwp+hpDgDxh7T+gOIdwm3uYdaTacT1zHD676IAvugYVZmJoQDHeFo0cbAo
aXZp5MYokdtjNaVU1dFzKYGmVhuA4b7v4ribv4JFAUous25IGUsQYX80Yx7nUrTn
SO38+LBHmAjFlZQcqaOd4WdMnogDNBvFFMl+v99Vro26KCAzXewsmoqMdTDSm45x
xpmseWPJzkXhkc1XlSPh9bBY67QbKpHrn5H7s2MV9TejodHf8GrHH3z++xhLgC6X
IY1+kW2BD81wNGwoxK/U55a9BXS3hHLTmd9MDCg4T0Yc6/E4ILQPAS86HRgqWDcf
jzYhSY+f+IkdWa2vUswR23wH4V7XIB6vZFNVeE6xKCNoHTKajg8ikq6u5dU5VGOD
iNqpdHqUbNp3Eqg0qC8+9E4HykD/mSIwW4P+THEe7MZjvWWLuBoUmFqOD04AoJCa
aFs99/ZuidIGI+dU7oOHFqlUyO0SriDCdp7Pz62ixwuLmwg6viShO+EPC6uKrcUw
VLN0iblmZu8xkYv+qSnqHp9fobkbz+XQRuwU/xOZx5Fp1URwE3U8TufuqRR6Z0RP
r85QjH71edQVGbQSROYStD7YoRTc44CmptMIEX7sURXIEsQESvxRxWhEDCPtVKQ5
or2X3vU8f6teMII97aDa64mFBWdWFO8a20ckA1FT+7p9RFk5irGZpIPxYMGYGhUs
9bzvrnePbpf4diYjPFAZkVbD1ApZE3JiilpTgr6TNSk+vpS3pUWUBNTSLMX7560B
+XXTQTp3SDmROXMDvbw5vF78NfIRB0dfHS+Wk/i99oL0c/RkmXBFrB0SVSP86d4S
gXmVbdAvJwGFKOJROVmuSYXCuJw/h02WQbA9N2FbPIt3MO7RdpRZpPcmtUOgSm5E
FeZaHj/5t9/H0R9JLGk74ta+0Qnrs635HwDIbSpzRuxy3GwYz3zizN+1PPvN9ApF
3+ZHZPCnQYqpbG52I3RZvrmOfVU7scJuNxttmoy9RdLCUDORlzRkYQqNsLZXSegM
RIxnAL3ZJ1JuEahvUTvWxKneghp/bfgNLUYJl4GDAox6P313DbSxQUu6G3ND8+Yf
yncCXWfI9e7IHXiI4krycMCpawixKgEUT/UPCmhn1xsB8q1vleFc+XUaZ6EmeLqX
FenLkcMdoAJ4inp8WJZvZdFlJux+ywO3fY4vtZyUvglaWLu4EkayQCSKqpoRSVdP
2Jhx/RKTrlu8rHjsljPPY22MyLkxoL8n99rjQQUMEpETC8h5oOqi7gO/9DjixWlz
0ogonnvqnCjIj14gp5C7Nz8k549rtPXpaR+fk86Pyqz7/CSvaEIjL4Ds1RYAMCB1
1YNbg4QmvXDxPTjtGmFxYLY62LBKgn/neCoYScjSSiYSHo0FxkMGmRfHrnPvCXG5
/JDA1rnGnKxju2bEDftWHkRgcGx5hgc3qUt7MsIV3GMdShOrhRezuts6U7VVDTsa
w/sdTVBYZA8JPgESOYNplZVMgpFIBR4N3Wgj2EbnQVKB2iaO1ovRD/7mmurvJGGT
j9YaBW9mZVMmPqzDtAnTnzjBPLmk4Ublq5Na+aU3ySPekWEYKdAL8R/+fRR4MDMV
hJye6LKSdUwji4oa2P05+f4N6gXQO69X0Jbf9AaH80nf57U8AVS//uOlbr7HrhGK
xwuGoV8BUjW6GeyRqqIW3KXi9LLsnmkfP90Mb28TplTf4NnGnQnenwPtLBGULhit
MTqxEmOOQEa6kNHy82ZyJV9z1YGPrdIsllNNaAJzHMjJjtQ7cDgIfZWY7jjdR4C3
MQZ1gd4WJL+lwnCBeRyE3dLVJ8ZNaEQJ1Ub6fLBesJTpOpYeJ8iarHjN9Csp1cmt
ys4DkEzp0P7vxM3+l75xsblwNPhj5o7wNVT5JT99Ve0/dOfzcQk73rUZ+wuPJ0HV
riaHiVVAYqmovZcxrR+aRHtkiU3KAC9pPB4Nij2hY0aS2epHKwPKaEUv17qA2SRM
AfaQmSK+Foi2WDfh4K3OK377s+bXAsMFCwFMINc5LVogiAN+TbTBhuJ+xQqQ7SJ2
9UjIljaSqt5ZFT8dft7u2iH8bJfuvTbsmHIxRPvfZ5mnHBu5LFTJynf7uXIu6pTN
MHBJojwE+1eUnXmQNjrqQVZhrw3XfU7Z3Oyltimj26D7O6Fls71piTsNXhLu9ycP
WOIicy+m0WdUAPwBStlyBxZrKijaO2E46koHYSrwo+/Pm2I0lN3nRfStbVzCPs4e
HGR+KP+9dvD/+R0jbVbke0O4pTiyYll0YWQx2k1Vc90ix2yPHOGEUZ1XyHntIO5x
9ze4e+diyjCSseoW1nnTyGKzG81TTf29eDtWZXuqN5hV8qpIitYRRppny19P0VC2
OSxAhK7AhRuXKMFVVoPonk528w2XLWE9APjnAkbEszsa7SooBprlWx3i/Ggf4x54
ENVRVhNol9+N/cGvuptPTGzbV2O3KyqMcfq+YuJs7uFWvARwK0Y6Un+br07ofSJS
6Bb0P0cTUbsjDEo/yyqia9XSt5OPXGDoZxq5uud7ovpm37WoOBIdHAFWDkVtVnz6
EkkPdbzQx2N9K3YNlcXvuZeCdsc2yitW4jVdJOUlRfSj4aZJcj1bZI8yw7b//p0X
pmZ5Iv5uiCkNvoa+CqGKXa+u2+NbTVyu5XehapfFx09PlL2sMnYlEgHFSqS7vdwE
t+IqPzoTXP8DDo9ozoyo/dOEmk1IhgJFf69aQ2e+mp0njxza7BOJsFkkeOMC249O
PsuUxrm7Edcy6N4kKE1iH0g6k4r8AGZ3NAXXGKXZlwWvhgAFEGqLKv3yvTd+Y4Yx
DANc5IFSfHQiBMUS+OmEGQV84TeAr6JZc5l5OHoqzJXKXnOCfB4x8F69lK3RGw8y
kNCjpfnMtMii8/qpvSf8Y+nd+S4jdDLFmK4PxUMWa/aaUprHubmW5kXJrjaggXBU
t2FjIC7MJhrn1UjFv/KUsbiTFk+x9RheXZMaoN1eLjsZQ0usmWku8umpThA+fOZO
ihQYDcdFjPysQbNpyHpgGbdcs/hINBuHHgvyK0Iuczjjsd/VwJ5QmdpHiIV+iWme
pG4QElvJPFYGs4RhGjqt856/3WJ6bmpu6Y9Bx6xHRdg6kNZDTiDkdPkBCzNedlI2
xfkS/8V0gdEit92yjvJz41dBhIzkhp/BKCGRojSBS37OYIE7vAKBfqdLP0bF1X8h
YMHBjIe4H1x1IxZ1YVxJN6nbbrAwFpkmsMkwzxoXhfd5AeRUW9odi3mVK607X0Ff
PCLq7L5yvPtHjZZCPSY1GisKYtRICL8nHbDahsrCr/z1hUFDBiyYji/MI6C5ZaxC
F4B19AUTINu9GZLCE3s/8lHoYxlJVvUZ+Z7WM3+S41ud6v43tVDHnwwzQvcctuo+
VaeibHm6rEkUNggWKcU5ejVCUF6vKDe5KU5Nhz5ZKYhaWuzQ0b9NiQGhl1HV4+Tk
jrV56kAVJ99SMyWhPFK9gqM+XTK6Sv+6U9ei/7tbW5mp2rcswG9Aoj5skwOcI71i
D5sZEpUReetEephCX66DKpdCRS+bnRJ3a+T9bKpkrfxsjCQy4seoIk3Ml6hvne5l
qEhnGNBHqbXsiv2naQL9MMvvQANLVLchTHDlUR77q7Grs7zUrCi3CgaP0QH5L27D
kOVpsps0/2RsmZRbu9w1huERhCAVcCyeYj2LIMI99rK0UjEjJ91mFQ5NcBlxbygG
N3jAPEIV0vU4vGPSwQf5MJSrH2E8/XJFqxhxbltq4ARzFMhc3C5Q9GqcvffmmN+Q
06yYaNn97K5l+aXSHqukPgNYDOvnT/oqe/vEUmPXrnosZdLARoi7fuVhcK8kkkTb
P4aH76f1qWXRDX4iOMlDyCpM0fe+53BIchcuxBaXLpmq/i+FFlT8XJA760cKhzM7
BykScLEOe2QABxYqkU/YmtCnvUp8OY7bnI5aj2M54HmDXIhCPY6YJgp18YVgOVUl
LpHcrEWMDBW+A36pgak/TlMYYSsy6hdFcZ0C/FRAWX/YGCfLwtoYPHIe2eSYdJcT
JQ3rdt9RQ0gws/dZ2DaA0yXlRi5E4VyEXTi6PBJeyH6JM+J020Wcs4nqdgM7mkIH
pYJq0W9wcgCPX20EKSV17Ny1eje2eJW8CQ5YScqJZd9tAqu1N7QeXCU/t0mkwABD
8Z3RpQfWddJxaaKsCeVLnxtn07QDHQzKKhHgQd1jj6alfSnKNPj7a0xYG2V7k37U
Z2ycXXjeIySA+AjlyhV0pdj8E6Sx5Ch3fxeGpAbWHFKo0Ep4Tzjecf6rvkSqu6x5
iF2hxVGEh7vMdIs3GGaiUl4EDqM78dLJlvAK91CpvTrzxG0g06Od0cbOmmWfB6OL
qqaFdqiLpsiT60zaWwbAA9bfnpB3+Qaw2YkpgIl+9ImbHjQk0drg1ecm31wVfN7c
FCM7Oy5iEbNu+LO6HspGRORlT8nCHt4X4oAS4Le0tVGa4Kibx6QleyHB+b2J2QdX
xL84ZVZ5tFXTuDQu2sllVunl74++dRQ9FTucZtfHTMUavpskePFQBLZt4UqfGHpE
lHa/Uhz1HOd1Mzlv7qgFXOkuElTfBxgi/EQJ61/k7uFaFwGmY05XPovNtJaPwrDl
1JqklcWN9sADAt6/0WHlG9NBhMFTSJIuUBf6m5L0w7vZFZ1YhMo7V5rpHU4NhRYX
i5d13LHb0jPA+0VUuSSCFHBd3TrTphfbakdFOuOodJNf308dYxTH0lZiUyrlWMJh
OHD/6SaiBo6bcq8JCeeY9nEhmN7KPXskSt1V7tslzzEV4fyzfBK+szsk7aopmyR6
7q7v5Ea+J7ryBB8CLwZV5UODhfYDgq+ofky+ULKayDYlDgoCoQjsvGh/XxPLdLbH
sg+Xp//6XOhOSNgKK9InnbMw4+I0jxqs5B1z1g1PtDhNEpfoUS/Zw2F7KInuzf6x
jzoWpFORo7mMrSh7hKjUMkKehOkWru2+gUNOvMhtc5n/Uuqz+aOSGvLUhznSAfhD
vxbIRvyTmWDLEqeVebFz4+FCjKpLrGupOlw52UrDtwpT7Msu4gJFyWAQ4WzpaFIu
n+BTQwPkhI/1UniGZbZeUlX0FqvD3LFTrQMS1MC2WahR2SC1b5PkVMtRKucllsCu
yHB3Y0xGvxPeX9KbLgMqiw+fujWhmKqEppqYALVaiEizEY1LCrb5IDbP4RyO4HAg
IVWrDBhs+4Cryuk7Oh27TksA5IHLx8g1APcN42yxA9VjsQCc1tnkRudJClLtnEsM
OqkkfkrcwOPqQlAkb51k5nrQJfG+IuxWldrO6GvHL4VzyVgmfgS/nPayk/xMy/op
5BADk+gxfk9RnTXsh6HpchGpdQv4foHttYaCmYg5zUXS6/HtcVwKocObluhxxaeN
uaICuwEUIgLGp5AYkNfO1TISsFTZJ01+FSp58pFPlkmxCQb3DJLJk8mLl2NVvwmS
ZsSCxF2Mf5Jd7QCAsFNVHq8hJKVVxQcFajeuVB+jx5pEVPgP5xw3rqZpiSNx7edU
iOUKDYudBLn3LRDquO9OzaGFv7UDkFgIxuaT/G1tqqpuANqL0bfFIQ+gNVQCo9Se
qhu4tCi6TmgtMpMPu6Q6cHIfjVHaa+q9UyjtA1UcVCpnJxNF4k2/g0e1pw6l4NCD
0RhxjUjWSWEbVk1+FhBrnKDpcRYrX04B0rcXQvKBhDuC2g8biFl9bbBhcJMKq/pv
AYT5W5rHjaLKwk7c+BeyTEwWtyU7fZI9sHNpEZxX0XWyq/68G2NiKoq9swJq3bA3
IhgUKkK33uVR4VpmgANIHs1SGLOfNhFegN+8fFdE/y9EssQDYFIi3uwTPIvINust
3J60JSI4nAGSljNzopbkkE47Rcor9sRvXATPXodO5ANHkzhzyZcIk9m3m/3PmG0Q
LlERlV/DlHz3uyTt/s83T0+HqAKemVor0+ZAY5oxwPxMvpGv6LMrDmMONp54V77Q
+gUFZafNumiYizDIqXBincagoRjx3BMFHeLx/VgwvANZMTwd+rti3+KH/jrLUScc
rB0fJdoJG8e350lisckJeq5yeXrzfUXxhVBT8VDM0oC9st4CZJKC0DU5nDT1UEI1
TXLZR9LrTQGK9eEoYsnR2WzIfTOGn5qvsbg0H1cG7LGAoutFU0ZpdFqX69eoD4OJ
AedwVfIxtE/U536uRJGfPv1G8NBDJhljBI526ooyvFd+Vy33bnnop2tyc0EVtcwT
f7qcAwzR+2w9Ht+raNBjnLOTIOeyE3f2FQTeDgisDM3fn2Ittsxoh49WS3CYs3Io
ods4jcSlJUSQKE+Xsi1nlpbe0M/F6lB8NHKXcQgk+XQ2GWILTV7hYq6S0pc7RnOK
bGP5NakDq1cQnfQPGo2nTW8mlBaVpuMl+nOoeCaFEsYEjsBJ1q514nZ4C7+ZdIGK
XU1VmaL28h0RNF9iqFvMLtI3My3tibUrmFHfVUpvWuu8MQHu4M0rLKjHWHSj47LU
54hkzqm6TY7zLpvB1gNW3gjdov4FrlUmWQw8VwbjxjMvOdHN6d2SL2/uNaa6P8Ti
6D/Qm2bN3J/reoVDiWhGnXhEn0VeCtFsjN3OFPHfUJgNYhTi/Vp+MToXNn8Yc5xr
q2rc87KNbA5kTKd39VPNcH8amnAoTP1hljTwljIPSC6i4kehBcQedy6vPBUMBDNo
+1ecYMbEIT2t6C9H43oUbXN9dDvud9Fj+CGrBIdznMkWt9SFAcVLBG3aF995XaF4
yXe9ncRNidPXQPdH87Y+Y9Wv2ReDGcGaVW98Mz5KDqThjlVFwH0eLn7DVwP7mDOX
KqMXI4nKhMsSA0JBgxZK/sGNZFc8vtvwvJUFdYKT32IdXqPlBL5oSq8Hd31m7sQV
oQWkOGkpFtYJB2E200W4HVjJYnxA2k407Cqu8pbORKNRWM2Xh9dksIVsrcGV6pfo
YTtBHJ+zOa5q8i3gVjhlDpjCOFxpMbQB7wfEC2WHCf2BZr7W9p0jJ3mkRBIN/maO
EIf7n53h/L2b1EsxSV+SkVRLDM8w+5+OA604RrxqSZih+qcqQkid5s95Lw31/fs7
pxgkzhsyz/+3Bv23HXdkUGul/tJehrnXWq6kkkpm2x8at2oxGZxyZETEwO4o6uTA
T4AnXNOacBy6SMjY5Dxedo9sys0tQH4/V+vLhfj7wVbUaoT/stx7AM+B+ysxNl1g
++yi7qdxlzA+rZQ570LEe346HcUcmi7w17aiJlHV6jpHbWtnDoDrpSGxeypGOAm+
VZfYEw29YfKltVFWWsQEdkWHOL/g44aZJJfGLw/CK6rfSfRoNj+44FTBA7rJogG3
oJVafEPw6Pe4m7NXvJtcxV//xCQnv7SFTdo1K0NsUTsXZScE9JMVHKNDG2uvUI+M
zBkgQoij0Xz15RcQbKRwwHgI03m9jFfQmeVSW6XrYPEVsaRO8dgw4iarBvs1unAP
wzTH2DJdPviL2nzrBRf53RPwuZEQkO6hfBFEZKJVDn7nyviqRIehbGoA/6ytwVw6
QYC0mKxtkkPUHNE32Mzo0/PIshqvjCwf9LxgODJzeeMvMIcGAQ3eJ4xaFqK5cEVH
P4aRnfS1fhs+QbS9zMYUzm7/OEOZuMrTSqTskoYNPJyl9Nllv7BB28tEzs9VWp26
RBYTMpwChm9xH8lvL49Mz2nZid4sbaRKAifK3BFyxH20e492wV52nJxuryaA7Ldy
tn2sY0v4txtkjgF18xsQG2LL4GY028GRsE3zzwJNOdZSoeJDgycjC9dOK2ndYiof
3JvHL1Ub65nc4viPKwLMP2nCw1auoBCTMp3qAM1NktulXrsN29hOJPN7lNZV2oVZ
w0rF6vdl97wt7RCjyNMjX0W1d1ouL1Rx5y1sAuvCMq3BkPMJYCSr/CwS//6JuPK8
ufFJkoyAQeHnajB24McwGXvuA8dk2hLt80C9KQ2WqHzg7Wnxcw/daCaHFkKG1I5g
XWvZVk7Ywwsl0Roj/OMXyVw1RduN5yHjl82wTQNvK67FHaLfpkgfbM4Q04xDOOqt
OO/T2gnSB72PemvN04bcI5wxiZ+EeoNwG7PI7Bag8BHN8ghMpGZvv5SePAQ8Viwp
UjvV3aS5rnMLn0qHkjq3B94a+xPek0XpS3j0Lllf2HUZMxciraxeViIKdNZeaSMU
kfyMly4tu3Vv8Jh43PYPfwKJ6JSAJ2qPm/RksEUkamJESN33hRhKWlf9tFWaa+EY
jkgJR5a0WnOCyVhOhPZ1Gl/YCjJJe3/tG1i+Xt5LrtKPVbXihN3yc2vjR5Pd1/Pc
rr36dE2WdVbnuavXf8/qP+6osIz+fYz6u61oLOPbawtmHF/3cILa+ZiF+IrSH11K
1j/N5uBWrzxmuCK+JsfjR/ogKPndfI0Q/W7LyeYtKY2RbiOnaGMwWyiiEd8z/nlh
WjjN2RL2bpEtzZOrRIsu+ZjbDm3/MVuUqj3qVHaIPol1w+Rg6Tfk8ehwMkzYCRzT
fkjN67FHAR6YO2/Hf1Fhkd+a/r6NFtLDoWHZ+rOhphoQoFWjFyQlKdbYvdFq2wJ+
qncJ8jAtCen6auFA0ls18JRM77rKqL2KMi4/W2+8sfpssK5WEWNTSVR7yDGLdtN4
J81Mv6DAjf9OOxb3xRDqTv1+UMPcT2rmaNFAG+ESHtHPQxkhXyBV+4bnvtEecUDv
ZtG0mqrxH4z+AxAx0mykfO5+ps446HGye4zE1QwjXSbkZc4sOROMkUVokYSnCO6k
eUi4AqLhE/mjsoUloyCov0Hn35B838WokCaGvWd7XL8JiMXRdheQHmveh8cZevc6
KE1YETDA7//fTzI3Qc6qy00iKQbbi5HEVeoPyVa9cKWl8R/E1L9DxVrCBNQ/9fZT
ruDNrrCWNe4V5D6aRNN2IlJtQigAVZdOIRYU+xSdR/8R8PN7fIN1WCH8YU21VD+Z
mkhmiPtqrMQQZQOXvL5j0gir3s0IcXuI8TrfzUR04QU33laTFNWafxsc5pSXNs0S
BSOuIS+uHvNyWOhxH4Ys4wYvWSeYYHj0XNAiiqjvPw6jyPeYRMAg+6+cIeBFQ0FH
mIvjVCQf4Zp4Y8/JEmrkfLuygjvDLrvTmfZ3/eqQIF7ia8kCdLIwa4qYFkSYbDEn
3zkFfVGYpmDxbE5m6ksO1NE6TsSA3F7TT3Lp6uBCwYT/AyktbgC87WheGfRrw0bw
SnyUXRWXt8VsBbErYLFUU7yROXrpc4ElaYaJoPxS4ilEI7hnHLNWNwifjp1EoXQ0
Z4rO42zGiz/CCGNT2Wt0Jr1gqSOvMytyq7ErUw/gZzBgMxFooQAxVA04i689DSnv
NmHW1HQhBiVLyRfUpTIWLMgokPx3Vz/bh4/aViQwE4UZrQinynqn6k6A2jjyQFFS
4qsY11maGcsP1TUz4W5/nzccHDOapcbR6Yd4lpt9HQOjhVTZVCPT9HWhtNhm7alB
D/J4BfgbGRDmVWIAjTZ2PomPf3seWAx+1NrJgbJLtirMj636GUGXVpZDYETbA+ci
qUiKf4plmcmmx39kF5iD4ECEz4CYy5Bu+txuqTQuMvzRxFAMIsQXiDjD8WzldwSt
tYLi6O6Q6VhJXfQqewf/m487XEWo8I5QooHggg/TaUHOettRVKjsAlBlzRFFU1cj
g8qJ7gyK7v8JFERGJs/pkqK1N+9SR9AzYw6jPJ6f+EtMle8om+ZSWCR13fmmCmUR
1pMMrvYtj4GwC/s2aTokFlxhhqYqivXz27mP+42D1y+I0wan5kozSlh5steMglPc
ZlphvH78qRK9C2iKISziLD7gMU68dvLRg/ooGwTIE7jSX971890SjJcC8jW+951b
GlEul+QjvUqcE/5NRx5gcQSoiH119nrgAHLzvgMRGQ1u9naoUjZ4wKpRtIYDM9ud
8fCdiE43inl3IhjbLYUALlO3uA6eRWIs7Cr2+EjckuGMMthh8UP/0v7Vz6vuwj3n
nlN4OPBOOyqWolAZjDM7yypLVupoazYa47MJ8x1GkbXVEbIBPaSF3DaFodkbfXOr
9d2ZmxuQmSi2LIrpcBaGSO/yXF5G7b9C/nDEFJshSD3ciI3us3p+N/taoTNAwcad
wYTTkCwcoEafaCIMSp9574ZI6UaomFiQi5Q7+B9IDB342gscjaiTv4wrPYb49ijC
YBTuq9wGZzOaqnirIwzarkuzsyETFLUa9pidQVt8fq5rmjgCpNvOqacAqLyNcMsU
NZpCpbLtuSLEc75EFB9NYVgQUtTSXitnU+007MrTEAuSoysdUleDSTaO7A0ojpWO
XT9g5LKSReOzapDdrZ6N/P5ISl4GN3jA8WRWXiFQM5zokC77z3m2GaSiJ8JwD5cz
FEMhsjqtp/uyTZm5g90sTBOqKLDpRaIB/KGHy/ACgAWxt0XaxbxPko03fc0KX1/7
y4UENUMhWdHuz8Ur0A26k0dNJCuSiCrXhl/+sYHwiEtKMULXubmbJR1SqS29ta3b
dMsdaiGhTBxL0GrGVcuwUdRH/fkKQyt6nrlUPpRUTU5IBYJENezDb/reLMrN9+QT
1mcreqwifBAajHC/S6h9HI0dxoG0e/BDebaZfTnMPIdJRW1Pe2qKQ1eJcT09U1eh
PVhr7E2jxGnVZp85sIqaEOporJBT6IKna+rVrQ209lvz98XxByhlLw92N1qtLQwB
9w1N2uUBbEhjT4SxOg4IJwlY4XojiSMYUtSLaDrKdyR6+cJG9xbBOSvIxji6S1Ld
Jy92OV4fN51+P+NgnXWjy1lf5mj8fZ9PqkUCnbfAd9gBLR+esaKxC4HwqeDiqa2f
iT+h6W/Il4wNQSbMYPre6WbNja2t+iqPt1jt1jJ84INwlEuTtRvRtuBLFk6ks2xB
ZtP9BP5s/LntBWSCfUcTQLTOT22UQwf/b4zeUaNqfqwJ7ukAhM4JC02ms6wZttMe
v0ElD1btuNKJuZIlxm49nZ6zSZcQNBZizcoR2FaI8ifqhXJSjafN8eX03VokqSbq
/m6/+EfDiOQisBK1jro65245KL53OGFLwSxBF0Pqx1vYKsdq+dmWmP0be4nWEuLg
Wn6ZWVSUr6omL0iw8jR4zi/9JMjIG1xgTvpBLC1lubSXyQ5BKJUhaqKRFcM2+hqT
sGMWjx+ByW62B8xyvF1nZuR+K2MP/sgf62DPulivIyyDbU5HorlswLSj6RFAzvfn
FejGdE99YVaudXsYDh/jjEDk3aJSNJ03lgGPxINFi6khV9MNc3pgh0wReQ3WZLDV
kJicPntsDhFDZLj1fHSduRAGNGQLh5wgdlQY1LNPPMrtwRtlOni7S9WSbmlu9yyp
Ty5GQd+0lKIJcfz2MayVboi4Oue3nsNgIj65XDePAtQgDNQh5iXCG18aVUJvwgbb
II3QgjOkz/VtoHSCeh9QqyzVdYY1cPRS7ILp8+S3czs=
`pragma protect end_protected
