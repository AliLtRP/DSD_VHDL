// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:23 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LSIN5QlG3Tznte3TwRSVHjch90rDfAbv/22SFArc7S2VpB6IdtK+lOtO2jGYgGi3
W1NNdmhD0vcxdADoz6zI5gmDA4Fs7kjEpVcvLzo5dYMcG4ffG2gdUnvsycqRRjdz
VmI5wpVpIFacdnRP5MSOpbVe1q2TIC73S53i+xiKGI8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6768)
DlgGadH8kmK9dD6EyaWV53Zlu1PAu4MG9C5kCZ7BAdjRglA3eh/ZHEZIEPppGKB2
bsI9nOCFucKxBViKttyO+Q2oD+3pByBwvGS8w1gE3FApMRDvwSzCOsdpSr7RIRP+
mO8qguSwzLrKgdO3BxArnb1M2gsuvA50oidU6+bHwdgZrFBKrbAjBHqvTqScwcaB
tpLn6XDtqKGFVMuyh/uCXPrHDtPlw4QhZRdSXZqwO/P+MId4kJbbqSy1oQfjZPGc
aeX5XafLJIY49UoTl5h5sTjilqTDh0sequCD3RSFeDSZ/CJaXpwzjcDwLqs3VIAn
xhY07chIczBe2XyFrYAOzrhYMknNgRgW+mcCX6XF/tRbC9ny0ETzwvBvhb8af1n4
QRmBjhixY4mDj5Kvi/SgXkzs3Rv3ZgLfuKjP7p5AENga+TbomGmkWcAlekxs16vf
vdq5GXpVlVdbj814qdOZqBxnyyli0/xnSk6b+Y8BzEOaUmqymgR5z6E2lbyfPBVv
QRLKdS99QCJhdydDimuwfDZG/Mt4yH9Aa4wss6g6WJhGBwzqU4DJ6S+W0gbusfmq
qQmmu6l2zXJAl0ERsYqo6d5aU9FXVreTIKZqIsiELkYaqv4AxIb8UCVe/bjJBsVL
Seml488a5dtFtkYXPQNWgVZKbrUnEg0amuA0wD4qpcXW8x1Ldzur9HAqm7cSKOz+
/Jr8hgpgpsGjTmC+VeDuc3YqnUkv2lJXd/xPRCaK3nCMRW5l5vqek/bdiIyiNf+m
V2w7JlVjT1yep7OiRzA3Ddgm0tV26pmgxySKbw/FZCF6N8qwsrUM4ZrVE42giNLi
RQ0ALrgvKbfxJsu/Rv0aFTlnmw8Ds3kLkl7KpWJLrY71IY+ZvCEL9h0Naw9fgBDZ
oAJ7fYJMb9ABBkcdmVZG7UGJoy0kqcmcgmpZ1zvxTSr5ab99C52nLcXCA3ijfR2w
/6X2FYdqjC2/QMIWnW9a5TRWSPj+5Isk6fXM8/pmM+AF/elD4AgaQYBCa198zNUk
f4hpt8ifObp66uqwlUUD20UEIF31Y97lDf0ShPPg6aHicnDHqhzV6+Hi01Q3JuHq
f+rilrOjXuNFl99rVVkbgKp/kh4U9IOeYLCcqomDGzqLV/XAB1yPcjI7Cp5CyK5Y
7oiiE3c99iCVNJxP4yIgT/cfHPCp59ZUBE1DxBYy/YYHbRLJGy4JGcbL6syMcAS1
zBem6SeSvmdMv4oeShpc50KSNHBV3JtKDShkzyoOcMtqSBkre2Mrmx3b1bpcsiI6
g2PgbY8ZwkC4TBWFFN9peI3S/apIztkiJoKwrTVY6dsZljWpxvhLocz3eYqxvVoL
eVGqydh2674aPZgwtJVJ4aqMYV3WWsiCiUWmVftkCILldlaODKeYlDxQjPexXBll
aENdXbF8tBf50m0fQkE6EsvZdmPw+1NkVNKHd4561r3TQKenopXs/5rGlHdBBIDG
6oIlzknHNAHRRvm04QKK8+tX0qBwt99KRPMxdSHHAl1fu9WYfU1sHFrPxTILFbPr
fVALnq6hjLfs3H63Pwnpf6PPkSb8BpVpWj12J5y9yj12tt7k23dlBrgzCvHojSlM
QdWYaZ0Ax/M14qEmdnCEac99l5zRlP/mdB1ndgcr5eoD6Ci6gAiFzy9yrj8fNnpK
OlI4H8Wr7+IWFVN/vuMANLKpRql8D2IEK5l23L9SpFyq4bqZ71di5HbTvTpEDhsk
prrUDNtWvnDazI5uSBz2P6giavUb7UuaMyVPdC2Pj4zFP7oKwSsj0l7t09JiKDPv
AxeefWaOyV36Pez5UDbZTD2P9QLqOTVqjzzDad1ql3Jtjww3chWrrvsv14Q78Wqt
89x22FOH0vjW+WKsaQyoj/2L94eIXWDDXLkAf+TBwl1fj3JCzGukhlQeJ4NANwZz
7yNUg6ogSXaWMODMu5gD96hHrSE679eOIec5kMiJZXU4S2FuLM66OY8Ht8iG1AR8
TOIHVUwLvgiXv495I+LlsRgo71Ww5hFzPLa2QAxo0++WjL1qaG50oJQrSe66InEo
P0TmNi+U6Fo2NjJDlN3HGNRVAO7/h8wWTAZLYbu/oiKP29ZinAUmEKNk4jSdZ37o
GY3zy44acCCCSw+XPJiUyqB6TW0uJSN9BVoEX83TV3QeiFs/2FOnnDacfeGUScQQ
YlHZNYP/S9FgmgtshVljLt4ZOYwf4tGSRERWcANWy4qzPjh2Y/+O1yC3lg+/61RB
v/mWxuDEPZL9AQ1BmxzfW1FH9be+K2EiViiAwgCo3QcQFIUxVjWXVoblAWFqZRGH
0JIdM528YB/Er2LtRIdEaSJk1yJsSWpBsn5tOsBU1giGEE0TvDQcAZyTifNZxrzS
g2Z5e146uRBtdntFkDpjjGiUSgYE97jbhANd7yFJVuOwYRZhtQ4VcZ/NW8IYoBsn
GKi69rTc8dctnTamMM+4NG1mVaR3qF6AOzgJ49yy0MzpVPVTVWXW0ECV4vp8TLfV
Qo/2gXAey20wC+HWF7YU3yLADVwXlTCkCvo4BaCKojRGSoEm7ObyngdNkZLouh8s
lB+Ivf8TnqTwKl9mjTbv348fTMOjH755vdTKFSg7vFptVsbS2aTEbMeavPc8pWSl
tMFcw4ywgItZ3uE9zVimZvCMcJhd67dV2kxghKpSp+f3eP2BXZvNn4nExKRn8S/w
+DAPGNIBBPgRRwhrqofd6UP8d13hPM86UCVmYfEtXmGoNNMBJLIdHjh/B+mVrV9l
Rl6fsFfJdfLKKuBFDGy9mqgaKcnf0kRKaZP1wCwytuE7dWZo8lp3Hxk6k/ZDup3a
RLHQUxeD25Zr9syVEzm4ghVkWZno2Cd7Uo07hSzK0Q8whRVUZryP43C1M6oHEUBM
YzqTCy0EnDA8V9To+hIVQSIhdDLDA7tXb+9zk3eh6lIcLtdlwnKLsSOW82af9Mnw
PsE1MmU7/XTYGTf1M4K4Ouo0T8yAqHQp9rsCGAL2CSSqSJecmzGqeeMu3fu18eaz
dHo5JGI/5UF96C5jiSIjcDB6Jp0nK8evHgtkbyHVMtJLhPydFQBwl987Xbg4NDAl
LgTYqQzpMWODbyyt2JM/ZpsXlR4zI3SUdMJ6NZmRAVEns1iiW+zC6gPvruhU6QsO
PfoTXxB1x4upTDUXV3iXkzp2ttzjhpazV04PAgrDCJvRZCMtJwKsNo4EoW1cdR6V
6fxewqrSgKmN/f4oT0CLqsnGoLYxle46YXB5YDLsYU+gnBuGdmSo7WwG7qQbuzNW
NmhcKwe1Ywhs6+9XgAGtjoZJAqPiBJgQ8TdVTogIaloRlIl+k2yo8LRG+j11Pg1v
0kCSLF/sRANTvJ5gI3mvvDCnHVQrTOk0DGulK3DfHQRPzfnunqAOeGHPjVhqnse/
nmCJ4d1juiRhOWUKPjRcJp030b3rEZ896nITu8ZYvqdiIeRc0rTQ2b6H6QuOdQV/
FiD1A5G7+dTYPsK1caKIHwwckhKr7+YInXkHv4i2jyBU6HswSASUHtCDeHLOPbSr
AxP4aJ75FukDWsvTEUBkk11yom4OoPzoU4U8+dHrUbR+hCWjLjmoXoD5L8kq/8uQ
ZUbV2Z1mmYJv2ktpGv18h6CTAo0KV3054te1r/nA49eAHw8DKz/pjqPjg4Qr72+8
NHFxAy8ksZUBCAJtyZqhNc6SYkSdwdHWfPQxUQ5DApyQiCG3ype8vPu0x/+RvYT2
XrQZpl3e025OB8njPHZOOMerHnd8fiG12LHwR9aFH3ZB0biy61EvgbQna+9g8t02
RoOczfDZEF4uU0KYYP4dVgizo5W+mgGTnP6YUh3qoeOLSdtZbks5LPj512tjdLXK
gYOoQzax+esII1BrCQ4jDVLjvL0XqfYRJ/XUuivCZpijgntMKdu5/MCH6rPvoqGU
Tdq7grSd4lTRlKrhoLSU1OzQbMVPrDoHpbsOtDvAYSN9ZXm5V+O18L5epy/UEjKk
3HCTOI/QvxH6IwSaBN2t6tIdEaSBf81TKb1mNCt2y+3dRKTkY0x6CsjW9I7QnLHv
FNjAN2tllI2Usc361HyylmfpkYERGN/KNCvqr9fI05nwfMNwoPWN+TI/jujS4lPa
K2CH570AZscKsZY8xmPDarJjwTkKIxVEqIaXYF1m7YSOCtellyfS9xswBuS+mCQt
A37W6OjgAsObp+awsTZIF91QtFwTI6uBGzt1BysBa4TwfC8+8FgYcAoWWOn9VB1v
BhUYpxI2IcdHGrfvhkHP8LDNVxPVdtaHtmrztPG6CogKI2QhDoiUfvB2r6otAMuI
+zo+czt+jgIdOoLunZ7VaDS0UfzmAYr1VLXzlR6J0W81yIrvvCvCMAvqdJFO8RQP
bQFqxtRdyz1ziBzJg5wxW5+jT1rTsL1wBHgw4R0LgJ2tqkw2XE741OKdWbuXRE6L
R7sr4CSr7WErNWcuYEcXW2Rpskoj7nGY9gqmiFyT2sXsfCzIwYX1UBLXDUn3R0cX
5+8bbrBlm0l3KkJmfvo5aVsG1496wdtT1SmVgSmXAkbgX1dh6QKM1kiWwA1E8r1R
I1RQfAanVgVwcC9kUHJB3ixiXWp7XXqPZceViXgynhJp1unI90sGmxJ0IkYmC+Yr
TuiYF1gPJg8YDvocGG2Et1M5zdVqRi3c3epgfZYlyNSOIzL3iwKApU7W6lNRFdQb
7DI27hc+ohPbYNubhzH0OHqLBSIkXevg678nftBKEBjTYisHpxNeDL4payl20Zrl
STyNwWucTDIXszncwRE3qo60FPNPITCdDQzzBLVsPkglyHUdk3nCI3yPw0Q0m9xF
rY+b/SEWUGcXXVUPkg3ho+Xk/K0LvjhtJpRMuhp+0uSa7kMyFiMg2zNIyr1P51Ln
FxdYgb3RJ2CRFRw3kafaP0J+vX3ORUHUT62QDyiJwc4Hj9Db1aaIa/GQVV5v6B/u
wTKnDMhXiKWAlarAtwSMxp2iB8bpRW55JMdJqlxqDqdMgjtlazAm73Eq4lR/2ovn
YNBV0gt1k2dAqUzfNSfskjovrJSmHt23hQ/pTVlA06a35Qhz/Iv219NHitpHjQWv
IavzzaLKAH3SChBEWdEm/mUJ7qZpk9YKKFWSMYmy+2ViW1o5rvKVUUqIRua+lOTi
J3fmXEk30kO5hI4GBWnx07ZagGWPXl4MdYN2Uvqw93t2PpN49L1D09rkLBj9DJTs
iTHOjeL6XnCoBjzj+XBLgVGDR+FEeC3Qw2/X4X7mUDLB50Eb+m6ctifn0w9Bo6iY
cgYdopoz5XzpqjPlwnHrg8UY0aychR9ONJF2xrD+T4kT8kpzcmg2TFo4Hpp1FGSD
NP+k2Hkg/ZIm9VWlD9Uvt9da5OAznlS4Ci2H+oj6m5XL+YfttRnZ06AFFeHDyzOc
xNoAOCGNIQX7Q3P1dw0qhTr6V/nAQ/5vnOwILN7+hHvXllHwk6i6bcxQyl3GJeyK
YG10rvRm2xzAXcNYDJcYc+tDZoaOyYtAf8wPBfC3vf+fTZFIkjyVy1qm3Nsf7k4d
hUuNvslAyngIiowzwhqgBM5M7tZuQGW8JU/FtVGb5V2b4plXXzPidQZiz+SL7aPX
UASBE59/Su5Mgjg0hRMvGkANXAMGou+CLZd+dUHqMfzsukJ/Y/7rNi0nDWd+f8Q8
YaeL2F+Xdrk2z7B6Iu8c5priC4/wWX/7GW/wd6oqAKkC6pV/kykwF+47o5j9vr/T
055iynARdhZ5cO8dacwbRqZK4U+15zC9FR4CyKrHEM0mzWNq37vuddcB8gykkUhr
Dz1wyqZkvVHUjjqMKi9h14s+mkoBdK72eON6hJq+U5zau4In3u2Lx1GBCzrPkL3M
5lSc7d8Ax+IR+OJMBX7QN5xpkbyM0d4mstXV3ycu1/COLcgau5suQKCp2JD+XQ4V
snLU3iwLCFkOYQR2tQj/r4a60R+EdON7Q8MRnjWAB9a6jTLphqs9P3moujtkFHDY
JIgMxoRMvHNd/+8jYw32qnPPDrKo1lYxASAiXstjwUlzf9SQ4i1/s5iyP5N85A49
oxAYjQtB7W1af3OAiLgzYP1wJlYcq+IQ+FMos7GyMcoiPj4SAYW470qAgncunovH
rx1agHIEfUPYKK5nUXtVw2CSrvDrhAec/IMxtjCgp5INcQRKBnX8pswwaYP62SPh
JPUrW67XLWVLyigz8fB9mwMQSKtb6Gz1r09i2uaP4jPXF1+aDN+PY7ogPuXLg/oj
dVkNZE6NVHSpPYdYaBn/EwE16GeuNkxvv5TxK2kvbMoW5Vq7Z1Q2ztajPfEsJjWR
f5DOsSVOnpJ2zMzH2cPiTBrf1lx6+CDQlLuYcOLfbMVYDHdB9pyxxG2raiA6qpp9
cv7kAcw0Zx3oq6PDealQVPYc19p14DJTDm+5J9e+L0shKvn+cI+IDI3IbqWwy/92
OjZ/wMpMpFKORNznaQrQ7L42h5OR8rrmwhLYjwpzZ5b2RVXtXUqTQV1oLcHz/jlc
7OyU0YzW6Fe5PlXuatD8HOOhzl0LUy47NaPNrt05lHdZ/kGK7/d8jpegRD6yjUAa
SucwK4yyv4TAkgCtf04ePw/XOpxkFHzyQqH9WVD8wKR71Y869bCVYMuXXBt6umMb
Ku3vyOehWGSj9Ys5CKhe6Fj1TBHUpFtKdOKqxLlFZ6VNaD6OwdpQ7Dlo0JsMpNbd
zVF1VBnR9yrPxupVFUxH3I6q7luxY93dwfnDkbIIt4mC9kHrfr74qROsi21SiYHA
Jbtb5jBIQv3X9aBN3cosGtIowwycyrKbvlbbcSiUUxL2t+0c3D1wqLlEpKmZy6US
oYDz8WhIW4TorXJxrvnVDYf0ShiDe8l5D1c7dLfxRT+YPtFyDIhrHQH+5CIAPunD
kQxXJgCsGlMdB7Tu9k40iDE0Z4j6mhQos/hs/P4t5W7POoLq5XDDzJK6hpdlT7TY
Kt8IoLOwGylHL00/fZH7yZgqwjJ7Iim8vIKTJ3597SKJ8foPluGgVoHgnldmeWxx
aNgKkmHsTvtMvxbeSttMkKt2oV2xcnph3gBd8akd+I4ZiCnAQs/3NBTH7FuihfpH
e8fWXXIn5wqNb2gHD5KI/7nU+36rOnp7N/Mr4FQsbx1DHRRMMsYE1lrzHbnG3Z3s
SrDGJEBa7vdd7FPQ1bRaYmEyjXoNREWIrNgaAuVTcCuBlavm53cT1nLRZZbKM2Tc
d6JiGlUGO/zKVmbFuGYJx0RBlzA3ePgxntLHDJlKO7uNYvDMa9ldI9k1xIBMqK0p
LkyR0saBB1cGnl1yQV2VhRP9/k3gD5KtXUciqseE82kHofslYLP0p1v0g5iEuTM/
5ju2jHRhHAgF2yHJuVIWhn4qyEaCnge+GIPwfV6vDnckrnI+rc32FuKQZoURExZn
3jUvujYpLgbah8nv34pdBxP2hVboH8aiaeNzIWOuDnabqmtpndO/n6YPgd8pEqdI
5HhJNlpTmKpIrbYnpKL05edpkZhJEbYRXCaRitpMKJpW6MgKnd6bIXufC0f1NlmW
0gDdKmserhKm18OY5DtZgYsw9nx0c7awlAsItFFK1dwJkrZpFudFiLBp+x5iRmo4
3X5DMLiJto1g60vhusKI2FKrkoV3yGGRiuLPIeSM4z7d4EckyZy2PntRfQqTY0GM
yZ0UYoAJGQjnB6zJFCVB0S6gO22RZqW9oreKkqQBPVuB2WU7L5lCmFjmNGNDx00m
/IhHdgRYJfjLfA/Z5vcf7nRWCwASrZ6zgsHYM1bF1F6Cot2ozvmXCApSTW8hiOk+
YonCHo1iONxnqi1EIsmIf0wAMerFQNe7VxWWM8lXCmg1QPoKEu4sBSHWmgk5EVwc
tEjxaZtSdMBwPBL+KjNkR48o6r1pnwM4qM8KcJRremKTi0irWE4hkf0qIXBnnw9R
3QSLS8JUOhypbCEER8meoEHHzgldv8Cdus0jlKo1tmV4kVTCqC1bgHFdxeOaLHA+
uH8blnssbpQMK+TaMWPCmphVMfbgVKgbjZzCI2CZTh7zoFAAMZ5cuvThDqk9DPJ0
cP6ogaNrTV1tWmyzNurPYoPQiZmqsgm8/1ozdcJBfS6tsh00W/13qsr0wcGjlDeg
EK5tmPNPMv9vjJFD5AWR7sW9ddHc4U+kc0dMK4D7rj5JBfqXhcZSJ/7DJKhwz7KI
HQK3scCOghu9uiss75pkvwvxscEIBUCDcTiifkyoXcRHmjmhBuazCve7moSDMG4F
2NnHqYu1IuW2kgzBHn5hpFpgPx9uZ0aTYhKerMISWOSXgEgSGTY0C+ZFz1UVoqa1
+dZG5VJSR8G3mNJhl8LWTGcLOheNQxCFHDssuuE80ZwuMRYbiSyEYITpVSXeHn5O
gt5IPEZFvtRb3COMsMTDTctMYjT4tup81jnwHMMGjr/1lFFe5Kjs9W8ScQHZSs9p
PSyoSz7cYw5N60h2FSKEp7JmpC8drV4U0FMNQr3mTdJ4NhZPx4r+3i3DEosbW9jV
+HnmhsUQNuXuuSOo7eMWjwCXd7r5oOlwW1h4A0puT1E+H/UAHEHHCv39rZOjiFYW
Ig3j/vxXmbSmH04g8jnTw5UQKyYCIkT18t0MHK7H+OINR/s84JKw9QlHxR6I7S7/
me8yWQwQB4GcR91XaBkx81fEyXeTdFQNGBjKJiWRzUIplRdoVmDDU0cQnsp8HU3m
iuFWiqZeeHRlFn2GuloZ1x6260roXmERgsRBAisZ/YvDzUnIYmwMHOGSv0hoMJit
sQ3OA59ObM8ySTbJzmyoMK5PSQBjrJjUCWCuiU+sKdhQ6WUK25x5d/jNm6R0Kbb7
toSa2Z1TXUZsp/E7Kug+5+S50u90YuTTRSTUJnMPlT2Q6d06RuMkJwveX6iuS9XJ
a/MhFyqb3L9eioLnQafIchAa/woR4qq0yRrgBkUh+n9LtGSigigUYcnVph58efGz
OxOK0ojFegPIi6r8/T/2zASLJkpHy6ArGRDH479fxb/EavcUXX3xib6PwCt/F9n9
CEWjRIn7Iqla8F5xWjnGbktvEx2DgZTpMVRXRgJKoW/NY++V9Cm6u5F1gAyCULFm
`pragma protect end_protected
