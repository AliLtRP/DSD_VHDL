// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
e0frKaLEsAo7jM2fUonYxgz6ofdZxguyq6Nf76GHgcxQ6nDvKeSwwOPkyAaaRxplROGHUZgQCE/r
E2x66IomWa4CmlC7zWxOiF83vP+bhtG46eV8zl12LbSxCdOqPNMl9O+SYQLMR1m0IIxnTUZxE5rO
l8hUDEss1ognF4cFy7RQnWMpr9NjW09gK13ZuvGi7UqCAVCuZ/l5aA2DSnPaUS1xSPfFQpqE8Mnl
EUJROY605yzJR1tbYbI0LnTHlGHL8VD60mYgdoEABJ1QilHrLOTBRoX7A18ar+P0u8+AbT9a0FYA
IFmPOUIRsEsHmKhpHI0oqWxzYqb+U7F5OkxONA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
ehTVaHapHN7YzP2hciEmPwPnVJHYQNo65XVOFAyhDUvNgewaBY6xQ+pF1qhUvjBwHtKvH5QkIbeW
aQHBLVqLg29pR504S1SAUEulnmuVcuhwq5nFNuSb8vfXAz/AW2eUOWYvcDrREK5KdAWcO79wpGI/
yBjtI2Vfcr40p3nY8snY+MMzoeqyvz/LAely4LpH4B49MIS+PWYFrSfwTIOVrYD8Ui39n4Lpf6ei
6NxajbBtE11mu+BXnQnDOfttV3R515kxnyIptckI0WiPCS0MmFz5e/di01FbthLw6rd5t9lH2juU
3v/3TLmrfjNPIWfrRAV2v78BP9SOg+/550DHWhPz2ttwWvqUqu9LTtbjV8zzEsd2WIP50f8KPFC+
iqP/anf0NyYEWLd2T9LcmD/IlGGV8YBr1uWW1kMNAwt7+4OG9K08R+uAVVVSGvPoGQnbCnahPYiB
I9ai2tpk2iBOPN1glK6yz7IPIce/6g3g+OWiAz/6FrnhCIRD96EpZZC1ZN3m9I+ontelYrI5dBXT
03mfgnCilqtMB3MLCG7R0TD5i8lHTI9HiK/KYuXAotc5jloCjOGayOQSnWIo9zAVp4ZGyU4kOdpd
aoDC+T1ZxJ9ikDkPcK0JqJAkMYPuCvF3iDmisQ7ghnnC7mKwup3L+pVbQiwaWtmjiF/zXIB+LXRZ
6/4UVerXqouLeYVTmIJJ66Ec0SYHE+lvfzjjdYeRziFrMt6DiRc5JVnOcpX2Vz8UN79qN+Ru8z/t
x1NpytZE8k/Tgf0jASysyG5/UNo8G5NH3d5w8TOsz7uFPpGBxR6HCCRARWaq6REdsi+FvIfpsjh9
rb3orKys4Mrj6JqnzPAeF4XcMkCd8oadBQm0YI30Ie/BCOUH3Xh6ZkQhlW9gJs4M/Kve9Kr6jTeh
Wms2YH4hSkx0p2adGGjfa9yUMq7pOwwoV7N5NUY8pfFydg76LLYoBWn2TIXSKyccOhIBVr9wrOlc
H3ANn6ce2V3ocogxrgCjTfvoHLmHEnd4QDOCmR66SNkYgb5pfgnMLjp+dpku1+pS6ZdDoyRnsroy
BeGmWTMfWXYutaxTbvKvOqdvAanqpGqw4xyN4Y01Xt6JSpuzlhEhE2QU1m276SV8Q7CBS+gSVUcY
sp9yd1Hk8pyrC9bVOx06EEBF7t1kHZn5R7H48c6qAhFMkFTHtIzBt4gdOe4cAwfJwWMguswab6YS
JfxqMfQAxf/SDVaoNkEED+UFuPMnScToMwlZzofkPnwJPCxyfnvhx/20Kv1jsUXfnueufatnw7zq
c6YhNVoGvV6XUid3TJVHgLL1ZrsIhLGSIsAwwE1bxxAdL/QdKhuiUPtVEIwCceOudO7pK0YQ4R35
/KznxGErYGAlzjueyTvrQ7P57IVDm6Oy2ZmNiPFTK6EjsyUfEJFo+jiQimP3+jCxoLu+c/HEBQlD
gP0EmMJAdoQZOfv5Hst0GI8VueEPqUqXrvQDQcIYNFIzdfND5/GCW5lc8704HrJNolYqi4eeOzAF
ozI1xitGnYxwhujwg/1Qbt17DaP9F+T1oDSCUyma2tegHmoo34nt8qbmxydezNezqj4sIp7I6Lo6
88rekKJpaQlt8MpFOKjnzQvo+1cKvz9CBudT8QaWZ5M5rew8b/2YGZeiAI02dm071GTM+ZvmKM+J
a0sdUwzpUM2PAW6yiv9qCqOJfrQjggMR3y9QxdWcNkFFaH/I8tC3cep0D77JhX6PxVQU3VkC8/Zq
FVO56p7/cYDw7TSCu40OpL02DFz6URf7SrzE/oa/gqvS2Ww4VN5e11g6p1kxGbRFos7NnK4Cy/MK
vjFLwpUmJbKxTGTn4yTbZQZpMIKzYfhbArs5qK5g07wJO56sBPjJxw31/22LS00JD+T2K9vtNAMB
ToLPDkjx9qCSsXXfisQ/PKHAESyvY1x+1Ud6xHWYsgr+a6r5GfhOvesyS0NHzMGhny41HC3JQIB/
vEjFIO04CGhQNz6WCfi4/WeWVI4xVdOtbZmvw8uhdHKPxU2Z4oQpwAlumnoPvlWtXsQo6P5SpswY
Z1tZAingn+p2v1VCo+bERdGUIS3YmyP2fFfEwqNKC2/fdLRAeuIwGEj+H6tn6tuksiP+FdWzIO3B
vXNRLsbuj1ah7PHY3nrzOBZixocq6aLZmNPpkcFFbMw6lAYOP/tCsCzWqvWu+BgMohw0K0/s0AbO
pyy3+WvB3wuwo5e7tc9jvkXec/tYmgSB3cR3F3F7Ol5sahu52n+dWQed2MDE7qxvtiBgQlpHNIxM
0xht6LJ4GlDCtdIlTxzywAKp6bcQ0v+Ewdy+BEdes5Dt6MN/GUM1CtqKZtOObD3wZXJj23D0b4dU
W0nCIbBe9fum1CDbQdZbU218o22qc3ZyajvJkKQW1FHVAebHTY4RfSKkUeNCOk5j4TPxonYYGEPV
ZVoHG+eCW5H1+DWXeW1HHQPpYVL1thplZp+TxiD2neRe98Jzebfa/G9yp450/hIqcmlPd2HQQ51s
ZRDykgs4a67LVnuWHZ1MWb6c6K/fZNsQRN+ZEFxtXcZRhshwR5UZSdh6N2EQRZe3vN9YYVDz1cs1
kJukYZljjFYcJlf+Yc8OnGe9U1LHGyRr1GnHKKIK+gu6LPPUiRGQxvnB0XO4pp5TyqSMgnKeYo7C
hWQEDEE0bYOcPH5yEygSr+ou+Netdwd2TSi3NgkNCXHJHalOuwjnJpzfin3/fHFgpzjASCE4wh1t
9DEmg4RPX9wF7E6gzdg/aANjRcmrrCgXe5PoK5s+1leVRsg6+hA0gzWhIrJeevbmZcNPdyzPIGpJ
WzpYhUlV4rf6LSwwVVFekf1p3nxMiWenfA4bVfm2PKcvXGNpfaRfDyiVBi7hX3iUG28UNfu3Ff57
DJB5sIiJ91SaXYTHrZ/dYlBSycPFuVlDd+lpkdYyLnf9weRiHKWKvlDRlgolaEfbWyyee2GU8g9k
CcnNgVb3OnIB6bCPSBwXejh2jg97nsCfSi3yHoyZ2/aVmLqowI9QNFdUU5mgBQVDDRTQGx4GmQHk
OXdMG4w/IF5aTeQEZMMKHaO7rbvuzXjkSTP+1b8WDELRX0Qqy1arC4aXaBPGllyopNLXJDLS1FHp
vtZYy/C3HfSySJDsd+p+pswgCE3RPDFRw2kBUK3+YW1i7ntuM3AaLiZHAbdMQmX4veYDRXw+2LQq
0jPqOa4qYzrc33Ifl5bJF24cTTKbqo67+Zf/IE3s6QOPCYVlacmkCy+IwlCX/dAKc4OL9pR7KJvO
T086p6DxCoZGDhnUvcz8SzXyXD6N1NzvYUFQDW/t6oB6K2Yyl1JZkPZPOiGOIny+FhR49Lla1hak
IMTbvAPz+LHarZxCkX1PPqCMH86V/A+FH3Dm9NsuXn8LzpDO8hX3oxg/DOj0bQk2oEGyX6/MNBD7
+wh6h+fHgMGrZRwrvR+RVoNlkJQINjIsP0XLZyBuyc8ZEjap/mQ0r08N53KJhCwXHjiM+uNzRbEM
H6zxKPwWxGFeuMi8r9LHPeQYe5bHdx5wPWRiJfNdUM/BDAcZ/gH9XWp3hWeiXkEkngwuOioV4OOV
cyC545AsHRllI0GWq4eJfImjK1JRehncQkelaQFTf8NhMo4jgt52HBc3q+Hu/nfEwfYgwIRdk/7j
nGwPApg9Q+iKSKAopIvrSDHq9LPG5z+fAtMAUBGq1beHobxV8gvkPVeoQlC2qNYy/q11NlpriEs8
LV1BPphbJ8Psen/rFLFZIj9UBkiXuQXdUEySFTpDFftI08exsCerDM8xT14asediZ1VlDCL7g9qQ
Gx2gxVDQt2W1KLwR/Hj/XCC7E7SHnQ/JRMSreWxUGRW24GYjlMsUQO/TcQIYLbd18wM5AXmPvAYL
ZGJ0iSYJZBFZfXvfG34xCQ8QEqy9IZDtVHhya30t26pT2zlKZNu3RYpfC24aNt7Q1rN6YbZgaJze
f1+HkkxRlketIey7Y/c1ek/IC4j0lXsCdAfNkOlQZ1OSrjVrzTSgvfs2jkBlC3IWVG/sUXSnw7xc
3iyvvQYW1ZCLHqG8b89cN49TLESyCWXIE2JYZQIqVs/u5XjmrI7/riBPHsl/J81cLys937zoS2Jh
Suj4WCHqLSb/8N5pJClovgDYI+SRmZZ+BbJaOHYBQnFJpjpBBjyMKx4KaP//zDFPPo/YBKj3k8y3
gadP9qw5lmhizCDlZrXaRCtAnPWU9YJh4T+Mn1dwmezI1NQezFAoBiOlR4RKPBJ3Btv8PKciq01m
NmmGKUxmEb2dvU1flXqqh9yDbqVD0BQoWxzSHI+NSZtq66GxB7nGe0xpgJOgBj+TsuZa2uxTSjGU
71GYU1w6M/Z/Kvq+iwes8vtghVMmUJ/WvnBbxv8mlJHojHkV3OpLzeYZdNUZ+e6o3ogyyueaQDmg
9HmMdRYJnEJ4F6rr0ZIfI7eqSqJBxpcBvVC1v0JgvUDkVxzyqtPpmwcCMGVKBCex5uD+EMXnLhDi
zVhDkVisIUNw8LBvvtJzcSItnr+a6kNNcxXsMRgYVVZe+HpDXsZmd60QzjYIB7OlFQYEaqPp8gFO
effuA7//uNR/6cgSVJb0JtarrTneaVKvcHFtSuxWfqrRPLuaBAMEoAL+GTegOIuv5D0HrndGSQhk
3vyA7A04AxpN6gnA4bAGMBmNlT22GHog008c+GevZkKNSxt9MQ6ljQHJOFZ2kIwT2zElfwUwudAd
466rG8AhKR2D3AlFqFHGI8ohvfEfALtxiT405dqFcfNTOsk8yRXOwCOn7VekMJHrOyzHowqDWAj9
9NjnJ7Z/XJn7kSblhnX6hkIBHxmhHOpYhVIwIUvuZaS8ZN7cO93Gc4Ts1dbk/PG+1OBBAHIhNwgo
aV7n4b7GOBdZwfnbnj+OC3ndNAIxNw69jylPwckzcWE9dyW4fX9gGfreBRignATe6Gjh6jTFvPLx
hVxJSCuaHeiOZlFahtUOA7AFyyOx76vQiRPCLfbTD0aqW0Fro+fT5Kiduzpa57QI8MPvAKEq5hmt
sXxeK2bJSX/bS3jtBHty7a6RGiZInDxN5yoOMPGAiwdpOKO829qkQrAw/yXboznEfrSaG/LxGD3h
6Kw41rJEM0YsXU/3LPE2sTiqa7PxR5ZM1c0tCbvo0mRXHxTGBXFIY0JWR+yIqEean3xOPvYR+0qW
ncosl4su8Q7Enm39BX9uWUajEuCI2hHi+wQFaYi5ArY8+KvzhoDrHkZsP5avpXuhvhUFP7eGbeIb
/DTOJhAj3YGP20GndMCIDNLZ42k5wJN+TrAVueaBX6tgHpgxN8GsGk06h8wnylylSd0BmFO7QC6O
ftNKLZ1Ntb/f5vwm+q9v55fOe5w5sE2UUFkf0DF/Bjfsye+UuPVKd1VJkcns8hki4S2XjFv12dC5
CBPTTNvs5nEnv34yYvuf57XnLoVX9SGaSnqlr103BGaJszSJE2pIIiUXeOBma9Uy53Ua3S4ocITE
2kFlHdsITSRLd9C4/K/9rkRrmZNTCdxcSh2sHCK8YjXdkuFKM6j25HHgnrk0hQlMbSqN27Vu7Sff
z6JyhdU0G8/EosPYVxFHVTfQQWg2ndwzwQZwMD7e0LE0CKRLVbi+Vr2200k4qjVPK+Rsf24B+niR
GyUu5Ba9rmDjC5K+BwhtKkECow8jB/WpquGogqLJvlLfhoqClvT4LRc0BgHQ0gO/mwaGv3Up4l2e
s8nOoSNsbGKYu12KqhJXyXdbDxupdMVf6dITtteWpzs7RFQG324LeLxizE9P4Yu22jw0F5HG7aME
C/k9hjxPAsS05EW31xGsv6Gl8QmtRd2S6YLCLQbgUqHmwycIM/IYgfRkfHMftqzu1ZIIhZml3Iyi
m1f4Gtzid3fXaA1owyi680IyD7XCrngSuhkyC/espjNWhu/MjK1emUnK/1gXSgJ71t293dppGoNP
EXBkWFP2q50+GkhgeV/MJ4iC3Yhyp1uD9sY8OkarGJZrOceRS8WaFvE58PYt48fXQBtv2NyAB5fg
RBKyxvmbkfwz5tluSzfQd33JmfqX9xq/JwKXKCKcCukQlTEq0w2gsczqWRZaGKQWCZPI9tc2A54d
QjoHQhg2PKzPavQ3818LchR2w2F/tJAsVAz53hd84/N91GfxhTU+7CeGgAbyDhnhnNP2GImaF5BO
lMTE09bnXdbeF29srGRdijY8xvzLM11S8LO8H+XHr4S6gPBQmVpMuaKc0nhUG8SsiPtwxaLFfnWS
24jyyonozDEMKoKjzQqjQgk1stQbbd/ASjfzfWjTJHl2x7x/NBG36kH1LUZ575yzGtBfCfRJjE7y
NmbHF4z708EAj35dnKu/tEGLadMB5SUEmzH5w5GK0Ap4ko5jir+aOLUy1r8p3aCMNTj4o4FnmnbS
VxamEGGnWdWb3C9mgnw4qI0sxPvx2rd1QVAy2dVruysXtHAxt8JZ6TDKq7pxJNsuzJPKnfS3ocbw
hC24AED5TD13Duul8m135MF0E0ZyJTltiaaMKGo/EeeekFTUVSO9git0NE5z9hHpegZt/EhCAPWE
cXBzSIBqky2H3eswImfCmjhUl9vrpC5gr5jr9eu+VVfuPu2cRsCsPT/5bcCurf9sA83SHHqgwamD
wqtB5CNGzLs3/G8dNDHiXQ0DO68je1ItC+zS+q2o2RdmEhHqDPvNu4PptD6l3AVdFaQMCHz2zIc/
1Gkez9JlXiZGi5jmd9rgGU+uu3risp/W3LhKvyoAhP/w4FhqDznBkSOOtLTeCxeGKv31c3XoNoSj
OfP9uSxwlowjf2zfdc+lIDpG6udm6VmhCogrLFUZnU4rAj3PhkU81kUuguNe82p5SyoTu2QzBruy
sBOJbIR99pzeeYuaophfUGh4dAbcctNjHO5S4zW4u4Y73e/0OHtvytnu8BVZkUgGgP6yuF/249ts
DiG9dUzTrgA4lg9E07NgNEi6BXmmo5GLT2qYwEXUy0Zk3oN36ObTJw/scxFMhDVNSDenQbKU9+Bk
l9GeB4qu3V7XUYGTqxeWFQ1tuB45lA2I/PYTncNZeIyWFm+yP9NnbrPtk0VCCIhyz/RSaswmC/Tf
/73kL/nWNEL8znk6lRqlbMGFhWdsTTDSvw1q449Zw/VomhWB91+43AQCptI+cEm0tmgUdK0A2W/N
icrQ8bDx+SUbKAtiSfYQD3XtdrA3925pGwE35kHmYGVIRCWseQeCSA6ez4fC5dEaFJN8KuYL2qLR
eoL1YLhpqoxQTJ3/VLCZqi/zvlGoHXAQq4PPlONXxQZ8qk/8S2zmhqS79hN1PMDHZt+s2IfQ4UmM
cnTr2cIOJBbPOc2XiJbYRoLa9EU6xlNAX9xu144NIn5Vifhl8Gs/YJPNcnhxbZcT5L+dUXoOQTq8
ZSHyas6Uyrv5yXEgtaEIlhWa3HBDvdd5FqXddywxN34YbLyfWoCp7meyHYY+lZG5V4QYqvDNI8c1
OYiJbqx/oxpEGQ5/wlFfw+zvOhrSasMNyKoXIwhmk+0ClFastK7cI+5BGZmFO05UezjQNY62qKpy
St/AuQAA+XnHg82QWxIxW2iwOrWP+IJ9NSKDWNCROM7RhrSg56l8QEHIrfYhzzKmuuU6U5zZMIOH
pjP8IASSbZUC7MMe9oJ0F/bPtYCm07vARmYsByA06ndkx3AzHT9D5ZGy01WYpx0EmUyqt8JzRRpH
khS4i654R+NfqTbCWROQzwcc6nwPGOPZeorBW77s/Ikq46g6l/EogEEFQuOmuIp5s3eQ9QOvJa90
PgvIq+ImqOB2kNTMadKvQ/9UecsXz/Daq8pnOrWM9aLon98BopMQIfhoR1iYzD7b13hy1JLZPG1o
mQ445d4QhMgYpQDIUhg9tvniHuNdD10Lkd3oOQ7kQRaqJVcdmRR/RvpVhGembQBatJ0zr/C277i5
Uyym7hhRkkyxDiTkFOrYzehjx56LEAtYd7GHZLO+bvTXbjKZbDJ5C2stI8rSQDwvSbpLwliePPq0
sAp4WqjdvrO4VimkWc0WFX/rrzCywMcSqPBa7H/5K1W5Bi0QOLARyEtTF/eWLGVuGIPJDt7q5Y+V
6fzRfs0CibEoONe1bLNVBEfLFC66EBLUKQi1RcTX3P0/GeCALNeTsGtY96qZsexBxWaVHfpIQxPA
vqFazTEplRo9F9OwsbAaEtWhYh8WFEUG9tCEGhdSungEhRFjOinDqcnAenA+GfyzYGDZUWxhYM+f
J/z3wkSY3GCZ1oovpfl7AiBSvLOG1B+Ha6f9qsrFrUEFAX7d1KKWtTKbyt+MqOXMkm1QMb4o54e8
rtF0of6AXbH090JdrmO2plLq29qqtqD4QoNZR8TIJoScO16wl1wBMwxQOJDiypm4e+K5bC6Iusof
B2boQ6eXyY2quZjToXkh7FJrSX0GuAytbDSebzl6M297w/XS5eExV1Vu2zwTIPt1AaonOUVtKgzO
Ez432as3DoQDY/rWOMbBHYn/inFrqvFNS9TywBmGiYqqPdjFgDrPxYelSF2ewKTOHGJKyOZEFUDa
/WCHnAsySbVPRGPNTdFrfEEbpBJjmq2Bw+45fXWcatbFpKu7SbPXbV86PJ/DV/YGV0s3e5UordmY
3ku014UR+4AsuvDB7bjc0viiiEPG9gd/l5QxLKH3jTWqGFptkwOUFejqcX4L9zYnv0sSNKDhpUV2
4S8C5+Gn4aNUetOAq2tZPQCjruE2HkVf3s+5f6uSP2pAfCqoiobIAlk2ag7KXeri0dLWgLZeNWst
1CrFsgmocU2YIt1duXrMBEYR93CNIdL1Bc64T9Yxb1m65CPSxPu3NFXh+mLDs9pSoGfEGzi4fjGI
69SSL+lLGIZ1sI2IbjReA0qxVdFGKWl75PTVbXtkeyXyjFztSAo+nzd9pbFGkTwMGEzGqZaXWf6M
GAwgngKr3ayOXZZipnnitS4quFrygEwj0aIhd+vCQsjBUJJr0fp5Ya8IayKgjP2ZErcxWkZlQcHP
fVAbTGE5u6u4A1dIn7lngJVKfahaMkiviIgM7bz3r10qnMRbouLVywsra583fo8oCNvQltWoMD85
tbVWSt6gdlhXRetaCgfJM25gWAXKqSLZejfJkqb/huwx/Ko7g+fjFg7jYupFJVhwZkLpgyYIglks
VN0d2kZvSDq9lBDABkdGZr+rhLJXkhUr3IrA0QbTn+O/ndQ34XyJCt3dEOCFhurpQmyD1eWrZjV3
9g+GBuIEluhFGcg7MA+zF1ZGiZUEIsDuTGnVHHGCkXFQD0mU2+yS6XlJ5L9zY55VL9cKtMnPYuj6
HdznfrB4Ep8vz4bZ+BoPTHlBHlQTxNIM46oX6QIFLU0wYXrSJGq4xtDQaY71XlugrvpGoMYE7RZr
gEfHDIvhuLVf4Sa+NNtxFJiD2LOjVcXHNkNv9Bkq7bHBcEiVbvAeKOXqkyY1TEpOd8WeWu5f9vBh
4PdqHHlgSSTK5c64UkpPOu7pdv6VS3Brc3aWWF3ywJTA8EtyKL9WIQp4Qi9E3+1YylZm+ObCtjy4
IIpE8MNm+cHTvSzYwlzxJcQVpqHtfZzhSPpamKG9/rRw3B8aKxivAmTupvBRCATp1rzAxqnq5qFh
dW8LxBCDN6wBaQOmzKvDZHLOUASnqmUYi6x7gp8k7x8SWznZ9d1bsPss/i5ODoLQZT6bMsa5P3Jx
oEMEY64Fzde69cC9a0Umw8w2JmJD3HlauNk7Q3rReBq+u09onLvnm+S2n+v5CqWaBrWptDrwFA1l
+MPbdMdrL1jUttSnjcSxIwpcp9nO9L41VkHx+FVeBUmHWzNEWqyhVLaK0e4C4N4ADRnOJMjVXokC
MvqaLHVEsL2xf9Rk3R7izrsSCB9lO6Xv/ifybHG5JbNYGU+UNiI18j6usmlylNndqzKg0FyQVg28
2I+usc9xWoCsjjqilyd2jNTlq81mlnrWZBIMPKWtrzqmREbtPKuPoZ3jWLJCs0EQGkSvu23gEHvc
F1pGZ53JFrRrHvLL7Yz7iV8C9rSn15yVwgLCM+DiCSxwLpLpiNxHv9MeQwnshar2DLUS7dbeIHhw
I8LlzZ0QZKCgLBFXVtIIJ90bnkngK/r96UIY6VvmzwoyoD1YXnCfL/nv2aW8f7ivBhvA3rq6TbWA
Pwt6y2HkaMfqdC0nBYaF4wQ9PwQOWiZ157gIPCDM/0ItG7lmFIdYcqZ68SDCR2j72sRLwSt9nx+Z
aVeJNyoHKRjKeWFwDl2djJFatPoJQR1q+dh95viwh8d7ZVQZRGcGu1YHl2vOSnziNvTtOTk4DVp8
fiLvcXRtEXzBwV4pL1jU9EvE6JXSFnZqRCGgSGfrSoD/g2HMxNe1qdoXDtJ5mNnsBAtnrjSuZMno
FnK+raNOjKu/9uVs+D2KP1pi/OIYmd41BpkqeI0wJZqypHJ81eqVybn5byvjWiUSnnMV+IwkG+2D
xaMAUKxymw4VPaK55qvQaqjp33c4iaF9LJok7ljUsrkAGAo5W3VWB21EboZniqc+1HZc4NKG0LKt
9R/1B1yMVXTv/Rnhbd1ticLnTKgQDYKNoKWphlNqaM9TgPMrb5Astosme1NffyZ2rH8i09XyUj1i
6GyNHU3H4eLrVNZXKRW5kjf7xYMBbqW5Z5OaZmXLdyZYL/nmw+WKF9oh0ZEokcXsFW/Uq//+QQs6
L+zf8iTcJ33/ZBh+1KDUucYESmnSwXdCZDSNYEO3Q4R+55vAk/WBSWKdVPNnwpcynn3yJtcQ74Xs
5QjJLLgnr7V0CQpTvQJdg/BdWjNsrc/i9wpTa9FCd/M1yiYBxAqWBRSt3iUIsSdAIGgmYLWL8Im5
nhednRreKMMStpdWGeo6tg563dbkAAi25mVmAHQ/KA+hntCi8vcIIMiMMOk5RniJHQbuRw8eYR3w
GOPisOXg99rbb8kc3ggbcdprM2Lw9D+6BAX/iobTQeorXSosg1Jl0yUO1TusphAVq3q1ytHBDyA0
Hg46hqSbQQwoGj7GltNuYF8NRz6vWuqkk56UCJv+6sfEe6ZyqQx3krEq6b/nVxgGqKdAArdQ8DPe
3s0qalE1yFkEMUKyCpY9K/67OxUhxlHi/jOa1TmiPAeg9D0QWSYLnk9r6ZENtPgBVVsjp5MKo75E
owoEnSCaw5Jp8xd5AQxSDv5yjVimd30DYMyraH9f9aap4gAhXFhOqbrkYOc/YovRmhat6YgMxudV
LKWJydbzjGaCK7kcFZFahr3X9vXEc7AtRAHJqyNZpyT54l7XkuVbGn5OOgM25vCK1VrQpUG+/W87
t/tBrJIX8OGRFrpWGjfq0XDjmlfHicl2VokNIkj+D3UKVWuY7ijHgwbXXBQIeoVGQfpP1g5r/0kj
o1q0MAOso/bhDWOTC2x39Ge8IUu2NxpwamqCrLLQWzix8i1B+8L/cmFpwtYEhZuWbpZk+fh0OBi6
A0glpuskoIruAcYiz2H+KE0gX93+g0w9M0VP2JbwcIq1q606w65pQfTRv/XHAyQfC/OOQwwcMDAt
d7cxlvabHwg7UJodiyMWYvMZeTnCmelywxqbx8l29HUysp1+b15rYeYaOPrzjmY/kcY7BJISWooc
NLZCLlHOUjLyRHleGytd/RgfizElsGjbXEtq9BtusWf1WVKbJ74OTq9f6d12by8A6DHefoyjS/ge
acGjknKwkSUhFeodaPx8UB8jPWQkf1Mz00DK2FuoLwxS841GBalW5lUuahihJV9B/yoxHjEAjucc
XECUovAtW6BO6LYNfoHX3z182uK0NQ6Hp1NZjcQwCA3GAtlTSXT+kDni26d0O7LymUBpB/i/kwxF
TePsLqX+vOP5L/BL5/4dJRymMqqUpOyC+uqeHfOEPfA6clXjHDqRV0cmahctIxI/xM5V8JqLcUXA
Ze9/MijqVJeUn8IDU7gsaIwvibm8PuxCbzAm/VAkwCq7M9P3lSutCNOWzJ6NSjoaKtuShZhgnnIx
lWjrovsCwZl1NKieLBHQK4c7n+UBQiLBgnzm2GzABMSt1J2l4weeKpnC01v0KB5HsEvkvl3lXnkN
yZ/oYfVQOuYHOP4OPXJ0So/C2g9wiiRm6TGpf0Pc/7471+2eCW59TY3Z2CvoRehHrAvL8TVwfBRo
Grr0L2lzhYXuiIxEudujOip32KgtnJHzm1suqiOxYEO3q8hGsW3eTeZ7EWW94CzaDaAgodLJKJDP
Y7kPvWPY+8YkQCeJyC4d2L/04q6akRoTo4DgmuOGc1NgXUkXJm/sAvhtaj0JMiMowIoVt8buCy+7
sfF/I85q38SQq2PFetj40BUqh9sPXtInB0eActcA2EmMi9iVSS1OmX2pP3XXylDrIa6KFmIBL+6W
1jG+LmbdfP1fWviw54YqTMWzhGgiVvDrtjBXyTcYEHFcHtM/v9pCC53I1ZU9rl3zyb1WaItcT9NT
nnDfvVzVnhi3ozvS1Rfsui8lhSs6mNDvr55k6kWIqjSBnzdl6VC/I5PoVJlO8czwoahC0/m7Fpxl
g1YEI+TXe36iKe8pFblcCkxkglIe225sJW/qQuPfaevmwrXsc6SkV5gmyfhZ5a9vR4bSyWeorRny
kRCv068ihoOYMILVbZJ4eXF4I2yhBPRv+s6JfPwv4vISY/1+02PNwZOInm7+eBhv3/yvOvH8eUHk
14/pZ60Vbjp+akGSuwoK1/lXa+eDnS0zUFJzrbf7OUaj8nXElxpy9BQ3GnFt9Ep09Q0GPz/so3tg
ynvIpd569UAz0ssZhmGTdVh8RVNI8x5k6ecgJ7YvnYVSsXRxHlQM9Lnki96r2tIgPm7EaZB9hYB+
6QZgY3SZlUC10tfqb9DrxXO+GtwJu2z+87HWbNdPtUYnDMZv/SiepURmb6dNdnlH0gsC9UcUtngo
HnHeLVuUmaqMmq5c5XfJspzFNwistHbRyvdSFVqsD72xnLDQWGVrOFrjQPEfKS2mE7S5XpsM8oTk
nw0/QJAMD7drSgApONvebLBkDCpt1JF4AIsSoNPqwyPmQD6Vb+QXW4sbzDzBOeWwBQw2jIhAmCgv
ojV9hczU7r4LfE7gsC/CMWX9Yv2zgleMrU6Awh4+QppDZNqBubwCCg0c11qe0y5TFmh5K/6O3KcH
STC/fIYxFaSQOuZfRHfbJKunbSJG03CeGmNrXUTuVplLFd5dEPjlyg//7fkkP+TMt+DtJzDlFwM6
18p72PbIklIWE6vAe8kRRoMussxzA00dcReUmtHatzQDvEBMPwTj30GpBmGGtK0xiCnAoNxrf4/Z
4ke38ThTxjuedPxEihkR1N0pjPsfoah+N+Wmyhp7w2wFTGrm/J2XDhuxCzv4M+nLqE6W30eHGrLn
9uNXWOCAveaMzjyGpRFRj+yNoLoVH38Pdy1WvlneqyGQEvn123NXVLkkVOb/wLZHe5HKzyk9+Wtb
TZlHmsBdExdBiPzHB+GIBH4qug6yKj+NtBXKyBCfUSqOmfqHRG8PFQrW91Kw+qfWEFUt0fOKb4VO
DncYfH2X9p52YioynMKFUfs7jfkEM7Z+VHtoVU+lmfo8vodJJz8FGN6dQ3Kn84agtUNkY2djDKt/
9c/HBRCyBz/fo2Xx1ZRpSucNlKwwqV45a+3iKRbYe9s9oMcub9TFngR2uwNU1cjjXLuxYcBC4vAt
S7grn6ZfSvCvY80EoC/q4z6onSrz
`pragma protect end_protected
