// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:15 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HDiVaNkKMrBBzRxze0Sh7zUNn1s1ixGOwLteJX6+NV9wG4p0VwaqfmgEMVh8u1X2
log/at9GIdPan+1bKZRXiEWVc10OOS9l9rEawjGwZRL6RfRQxiK44gVBBEHOnsKE
7oXY1RmgmxCBkAOFwTnRKX4tvNKrCo2zGCA61kckyDg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9664)
jIrgmdHV8ZhnFN2sZDxTry+XnZMfmuayBKXoDg6Zh47C2seCbj3/F5C4IvtA2kkm
oMuv4TInW+2Eb/1QwibkzyndBaZG5HYAh9PsVQfFI3H8mwIkOVOy403c4O0UYilv
cSy1V9hblcWhajUS9yGuGGJT2PzOj8wcwq1W7pc+cK/V3jiQm0eV2l8leUWzWQL4
Hw5/AS1DQlt64JYTe2M7j+rC5ORKtN1Zeze9PDclwCp3nVP7D9e5hqTTp5hsB3z+
xmmI6Gz4AiCbgbRSd1FdqIbDcVwVSrKSJB+sIkFMfAuu8dSNTmrbsyHzxvd8lnVN
pvrakKenaMGepEpb1xM0CWNeaLhq/5NzHMoxXnvs0Ol42brAYDrgsgY1n2VwL8Jt
O/NtLP8HPocp2wIrSoSX96CE0dZhMSFx3fdXKmCXutMZwwdoAegPia37umPtKEqn
mdlntL5YvYRwBBfATXYQ+4e+JasQieVlaX2pbhkfjfS9xjQlY3KLwjRpV7AJhtVl
p6GN2NN78r5UVVE1sCEGbcFN6HEaYQxk4UEdKqNiK0ztSGXXpjqMqVrqgviQUwcc
/1PJfrtmk3JLEaz1znPS9/Pd+EqVS0/lBx3EbZaji7TUeqTLqOuLaQL5fXnSNRsI
hgyucV1Fb75+OCVixaeXD1mTNnAvs/dG3jSiI65GsBbxEdjEYKDU+m6uhD/lWnKV
MESewMnSVRvyJ9N2p7fpsfqDXOnnmWUrK0Mn8YOpmLQ8+h/5vIJwBYvKcaiAOxlc
Mw3V4elWqWP3p/jy96uuFntSH9xgMNIqw0HmjZ7RuLQ9e+YRMUAMjsRUwoMbGNEW
pQYv3Jr8oEogEjwB7lnLexdcdR53aGpB5/i7n0EbSoWDDQVSB/G0KjM7FIGsdYFK
40wU/XCq5pZdsQ+mHGuUx+gsFNlGzqbCrWwIq9irdrfzVQH8TfvQTuwIM+fk5G0d
eJybsgDODJF2UVbKVDskjFWnQW04hZ3A/PUbP41WvezLE8iS+WtVkrhcykoGu6yL
LE9nZDi3FLHRleuElKvoctG67YoqSADHTrTLjaw7d0G6ywRMs5khp7y/T5SOZ8Vj
MitPMveYkkPAuMXhL2gcbQsMiAVzwIZh6EpZ/OqJabQmZ/WplftwpisPYVjtoOW2
pK9Bunx4rajv+2rLTp4H0dbznU5rMZzgdddJDJ9VdpxGK5iuZcNjs25ZjxMFRzxs
MYP8mvgnt486YUkFXBHkNWvqaAPHEgpuCIlNcQX6LksGHa/RH2J/asso0pYCYXbk
vu9SuXCXuEUZQruBgDr7LaBIri1kAoQucSdsEyIAS8bQ1rLOxbUF8GAB8Bu/1W8B
qA6kx8wNzXdo46QA8IfQjRbRyu3UFVQizCi5RfEQKbB+65CZ48+sqoOvIyMDra7M
PXoJx2dO444sKUIhTYnuJwk+LfDNLCj9lhM8AxgcLMfgJyMN2xnSHra5TacjY+Yu
ILPobi4T0nsuEl+AGwUmyneLwp/ZjJsxeRygmzUhHVGSeKLoglXJ3xxtzB8NeCRu
loj7TqtbQF/7VF81Y/Lb5zBpDDELUMjbPiVwHDqEj7RDTsAou9OcBMpBP1cWKiLs
gPKg+fp3Ug8+I5/vh3CpQ+jTB/VJ8xCGVWPTwUM6GxMoXSKL8w9Q9E9EBWVcC43Y
MS4AT3PDxLZ0ojeGSyZ2ohan7h6L7p1OXuDnaFnyBThvLxCLzhPYQaJNMln6PIYS
4jNukG4oyIJCA1J+GXppLGyyZYhVu5oVnX2yvr34bKNW6uws1BOfuJ3C//ucA1bY
5zau0VjwK4vbiEckcX6mM1H5pNIvcEuaRHhx48I/GLTvfWg0VKuHIherepG6k3SW
Gp5fINRbcqVUErQnYvIfb4Xr8jogi0OCZ14TveQGtTVNpwtDMPMapyy6vpurlIL+
8/qQZaPpwtyVcVLstyHmFdY0xK3Lph5cOP6WOUVfubuu7JYp8tJO0Vx5loa/1+db
djk5Ndojw9XEVrSvMToZkbv8VvfmoThtt4+tS2BHhcZdOi/oHJsRZtQ+4zevZwlc
nuEXLrjrE5c6yYZqB6/bPoBngXF/WI9qDiVkKj6VdzSPJ4sPMHZTkJZKqyxMyQlB
cGn82T0T8N9HD3RiAjzaouUXSaltffn/h88kuQnWLEfgUJqG5yNSP7CDp0J0NRsr
rkMbWUkMilhzTFmNxVSoGAGW+UMCrpn8DvrRqdVBFOPa3I210Wcgs4+hxdkO4G86
omNSn47GfIS2B/uA2D8D4YjxwjMLh22zCKxymyNUAWQT1MYU1KbjASlT/4gE+/+x
vmGTTuEiXjHUot+HIGcjHm+PK4eq+B0D0kLT46tWzc6FCkMf1y3ar1FYJ38o66M/
aafPfSQJix0ZasIxoU/PIcrMgsJ2uN0jrnMTwyghLAjTEdwOtmALARIJQkrq/f3T
3qE56CmN+SmPvc+t/Fz5vVfyb74xPTTbbIsf61V2SySeeK+XJP5JZMcGFWIn1Sg6
3rEBl44Znpccg3ZMqz2B0x3WLsFd1cLtgUcyvXxQxF7I4LyInHBslR9s+xDFVWsO
ma/hggulxTfanAg+iLR3uhm65jjfVIZZi78Nuz749mBco3cyn74iZpEjx/IGqxzv
quLCuxuL+cVqlug9TyN42IZMDRC13pNUZWDZsL38v6wTX+jPpgGyey0K/j9+RRi7
OvQf1J0e3999Hg4kQPhVwJEAU/5Hzzivw7Wws8WnYmlaqOcMDEAcBgkGaZZGIM11
iphTafgJRKLU+A7kYmNJ6ysEZhZbtT2ovyUoApxTBr7/8/CmGESxy8fpN2qiiUII
MJ6J0ABr1VX8O2+hQaUB+ND6GTsYJZADY7rIPacKyGOHmy+babiHSDUx0tSmu1+l
ADEW0cj+TzzWYcZGDh3Sn838Yyjk1/SyZX1Hz5ZO3darQV95M7jLZJuKbM2/ZRq/
r4x6WehJGUl1SV0U4WUKiGomIjlLYfaZpSNdbtNOW3f04MWb6jwmJ/kOnIzgk2u2
NjD1u/R3C7W7C6wIiV+ei3NdqhcH8O8rP62foTScvjyaUBq5DApxco8julYpFJS5
MM4u2co6GIxL+UImK8QN1D8nnQhg6X3e2xyMkzwZiXs5xvlNkTsL8AtPY/Ro+Y6f
SQMqBOoBUzL2TyBsmTzd6W7+tVVCic/g3Nkc0cL/JfiMvu99aTzbewk0SC0MhFZj
l9EZeeRONB4NwYOwpqITIeBqgrTBNFR0twQVFKvUh+ahBmKwKFYjucTHy4b0x2Lu
Uq3Ij+VwOfCDCi+YKwEErmtaH9SzB21DGYEFL7N26xEHqmZX5E6JDC3/COQl//0B
jJJA7jhjGxcGwd3GejCbXVOUK96TItJRKJYEy0Egwjhjq/VBxdEsWxX/IOuP+fmY
kChCZazV5A3SoRjarEV6pD0NfKVTgbPwPVMs78iCWDv2SMVVOvtNDspMEpthmB+f
RbrluwAZSYGHjJuoidBgt81Fb0Y9TUGXKPH4WJZHbq1vvkd0sxY1k6znpGWZc8OE
Gl0BXwWEGRvTHEjCkekgzUP5dUazsNSO0P0sCeWcvcN8b0Qm67TUMyBeAiarqPDr
SI0+8hhkyHTGEvym7TCLmo1NztcvhCSJdAOAEVqhXzMhjVkxvgCotlE2ob2JPSbZ
DosGXuYs8vUKB/A562On9mV34H88GyO/jRNcN4YdDacufkhsCFQURjSrsGw9EYVk
IXHFbA4ocPzeuTNKWlY9k7W0WuKNlSg/ZrgGXyjq2/xv8AMQfho4hq8j0LFsMwbZ
jsn5KOJFR3R8YVeaIM7++aOC6XzUbKzZD3/IZiEF3y6591WdGJcF46CXKNjyphSr
sBktrNJtciigxjwwE8Fwj8ykB5Nkh4iUEHZtKXIyoAVXK+Wh0Xf1Bs79vO/qtZll
NtyzzIhN2/kKCipk5qCA8AJMz+qBnMuhojRNQnadb+ZTJ2PRpqs9SeKu+IbAJ8D9
iMSRZ7CBaQxEXDWOeaPW57g5gesfboC8lainXRTeGYqZUUq1QANHl8U2kIceWE3+
sOlnQQu1UELRTrmnpF4h8iLqnq0JwPzbtn4jIjdu5eUjND9ckGTBtBJchqtnwW9x
rS7EKFGbbhftGfvaTiQTf20/tfaHipUO9gP81ZDfwojdpRUn/yvZk3G3igtZnHz9
H4oGYU6/3N6mDchAjr6L/Wt9lTwGwvBBWQKV/L5x5KLC6NokfoeSdP3VoUzumJzT
WIXmyeGs6yPKwixf+wQZRUlBOzNBwbUvNDWTNq06VK4StzDe88ITF1cIHzNgnsmj
rTvbIp+9LPi+XNiHAPryQJ75rkmS6kO7pdwThzHaRCLb9YOgUhjrLS88kk+8Llpu
pgn9dfKNjtOKMZpxYVAd2HMqwksHhVzOfqO2Yc69XZyUpmVREBVJ4cfpo4ByI4cC
6sUBefvibduawF1z/YxQBTQlWCCUc6+4ejlh2fx/jNJBEimyHg2GH1pRwUT7qrUT
BrVYLA8bS6zYMZWcY5x9AYs2rZilYIKI0xEF+7cUcmilk9CBjRYFVWHCuGpsdW65
3Nflve1Kjf8bAPDOPpMxHyTCtFcMXGIyIdNQFagN46VqDA/J5ssBopTOy7w+/Gpz
QisCULAXRlnk+IhHdn57v0lBLuZHgUI6mrBDbSVSo18k9CFc2073Lq65miC5R9SF
Gl5p/crGJbvyL9TkxXMa81h7TBIgjfYS/s+wVATHCRWGnIcWVVzllsiTDQg78QNA
B5VI7lC27AHaVVbA2bpIbhfXdGSdSNCwVyzELlCi58thxDtfkYIgebvwpvxtvXFt
gATs0KvIkSBnCDaf4M/QkFOCTe3pFjQKF3eqVDwVa2RMUf7Jv0mSBxO4sdoZZVTn
yPXauMl9zwXBwI5fLGSlSbiT2Hv4i5rhMG/61tpDPEHlqKw3ItsZaQC0VQ70Emb/
IH4TBj443bqbW5UNouJPaNGWIKF4Spm4Ia5taDuU2pF9miXgUvcKv2blssHCHS5L
CHYA0Mk1Xpmj/K0DI7WRPzY7Nb5wkLXy0gy2MNpvFqxHGY8KtPyosrxQGnW+epxO
PxVtgIeYesSQVduT74H0oo2R6jwqxzBVe5RrFCmsadQojolJXyVWCFYNoA7NsyJ0
8LJljb3kOX3jqaMuxGJRTtIcb924AuYZ0OyC1tvTSyHD/dH5h5k9ykmexcvCaSaG
IVpZd9KmlS22+ijtY/uKRE2znkdKW4/MV96BcMZE0o+m3DIx97MD/C16wcsD4h29
iAdn7dI9NkTUAMdnzxN0ViPBAEaeGMmXKFtc/qAMpzkBsoPIcACu7V08IiOjNGU4
ScDYN5r97Asg6ZtvMx+A7EMCqr8n1aVaZC2h9ysY5oWM0X24OWj9Cbbgi533IwmM
GPNyEBLZYma8jv5JdNOtNyPOtrl6+NydvbnP5tgce/pe/op3Q79lOX4x+RVvFOJD
6VO9n2+f4s/bluYDpgi4jtovHFRp4FNuZSzD1r+cMC/D3Tb1QPYOzb8C1UWmh3tE
CCaEnxkGH/Z3QmCaYFvhn+9eTRLR1UTKFPsGvK07RKwOPA4ILH3PjZRKOiG9wMtL
oIXxLuRa15iHIGAUGK5KGpxtvnVul9AWINpNlGS5WdvHhTYMxV2G0ZdKk6/mZbkW
c/l2h9yUYKRw1OH5X8EugUh23YrqN5/lIAgLaXxahl1UoiBszdp2Qz12sw68xKpR
0ajzD+JtBsflUz0A2RIGSWTvKqxZbxpv182F5T91zyhjb8hi164TJ0WcEDTswfp2
VFnhYcwnGw7PXwmUvbpOsdfFoLu9eC+6lTWquzm9kMaR8o4vZwT8M6f0r00keShw
Y2Tj4V5JitpluDTffLix/IgmfYLCpVz7dBwMTiWK/ozR9ZY8+JcufnIgSAV1XUoB
zdthKF5tlqunj+zCHToX/1WgIyPAIDaixISOyS1fq4joG3r7Wib5oAUhaUVCDTqT
faa0I01WSf8p9jMLo+kmwXl+vdcUaBLg+unjWWmLYCDfEMNL7dp1vD51rhny/LLn
7xvu3TjoJqGqw2KnFOvGpSWsZOgteAHtz5P9fVrtlhuqcGzpQquVgZ0GX9gqdDcA
Y+87x13DJueie/iZpzL91LJtv4L59sgcXAsz5h5GkVwWuu/FOU/JTMzBvXyoloml
DOiaXtVguq+31b4WB8xf0mO21UpLZ5OVfL8fhHxGtRKF3jmIGvO4ZdPf3+9EzwNC
VxwFlsCW5BScqfVrhRZQ1BCzSY9clk4XLXCqcv7AzUSJy4GpkfcPrEgQGPKF01h2
TiJkiFWaEWit+N46GyyxoCIbw9iWPBcCz4+THc33V+1dqmuudo8HnKB7GRaTOW/D
8MqWLk0ajnyh44Y86vwR0s7JhKZAWGnRBlQl+d3wXW80f1NmkM1wyHsqdMtJgXeE
ywfq+WEWYsYD6wTu8i05Bp9naX+fh4PDJ3og4b13NcOMiyFKGquiRKym8/gX34WW
BczZxIGMII/VZTzY4YAO0iArId8mmqtbk3QynngPJXvVIQGC4T503XS0TP9osb4z
BAzXrJiTMOEK23FHsycBY6Fo2Ir8xKsOp9ecWc6uDrFO02qbdNuQhK1zFw+AKyCk
N5RMDoTGLypCDDo30bOKExUmh1RjY7R2a6GyaYWWa3vaNxyTv/aux/G6tl+2naNc
1/YEqrM4DbfoIKJGJ5QA3U8bv/LWa4u0gehp+f6NyrjmDL5s5pPN0w8Sc4r5BKjt
kCu/QnTA9eTsGKtWgS6hU6P6KSPj9UeFIyybgxOJFaHWAJBgF3uvNmXvdufE0/gn
KynzBwnuXhDyemiJ8hXNluHhkNvQD9ksRZgCnJGKy37yF9uSg7PEMkMunrPJhGcu
s3vVhPqYvgIxPxDlyW7sxiGupEXHKfQaN/I+ANBdx/sP9B+TBEHIebstCSFnaIyF
9KZOOTgbRA+7OYibZvj5rgq7Cz0rsdg8vbmDS+SfJM1x1kwvBXm23g355Mwj+dXG
ANznImElYZfg/817Ez5/DyhxU4f32evjdJmHpvgjlthUrJEZD/hihINrXY7BwMKd
x/5+JFaV6vZgjyazRkI9/3+CINV34/U7FC2Hd8x0MamgsjEymssme/0V5Sx0WUdY
CaT6yHMvawkARaEL2YZwFm3+Nq3NOAAZVpdOCtOhd39MQ3D0HEURid4i8aS8W98q
F/LPRHgJOP73kAy7VKFgpagqsOTub/m3VeYWYr/mqqDYvEu1+Sonu8QygyhoK9Mx
WOG2Al6MNtbZr4fX6lr4rnxGoLi1KSV6vUX0vqrI1cLZr517vtSaaAQYJiVKmJw/
16O765WOdrxCy7dWbL4HjJDcjH62cv4czexAVX1N7QkYeRMKp+F0vwaT6+UjJdgv
qrA+xzSjvk9KrwNvVDTF7DFCXNFGlztZQIZquI7OKkpw7YEMNFeTLnSzdjppn/Em
WrFwD80L6LTDAq7dW6Sb7aKol5tIwbWEZLETk6f9v6hUKXr+Lea0B2PLi4Yj0yCw
Wfo0ad0g22BvygEm2YnTd4yZdR3Yk1iDUTLCVjQBiPCwXFDji+TeJ2xkh5AGn8lE
drsg3iu8oXjztVM17BroXEyR2eC6TVuxaZVoLkwe1uepma4XnoGLlxOh4lOLEh0L
8SVaC8+xM1xmnX+f2JdUR3BBOF/TxcuqWMfXCK2GhCYI9XMKzU3hUtBWAiwzEY43
BoGRssFDz6gQCfp3rUoqTuS1qkneS0AbGGYa8veifYp9m3nt9Pxg+YddjW7A4k95
zY2QBgUr4YJBYSKRjvnBR2FFoi/rtb+pUwobfbadi7W2UYMNd/8enetUJufK1iO2
dyCliKqL8eWZFtoSwBSH36/dkUQxyCK3SK7J+EmLAeoFLlHqD3Q8nZiupYrfd7wI
qVE3Ag7aMqw90G0Rsv46IxFFOblxNr0N2fzf3cNPQ8ercV1FiR0qPj+FifmusKAI
Fwkb+lIggVAz0c0IOcMawo87+u1LaGibWNRonc6YMFoDhBmlzy7T2OjY1GsGBrgu
DPZHF8sI4MvgSJlWa7lsVUJ572BcDnS+weHysm49Kp5E4a6IzySfUc1SIAminGdc
Xn+zxqpMzN4MJO7jrI4GrUa40p0eTKHSC/4xIhIRONqqE7OxpnrSSTlRgoGk3w4l
oAva0YAKxwJzVIbRVO6VdjDJrOWPO7GV6kwxufd6kJHKWTDinFIQGx+azG7oJDqO
YW79/L+teM30AJ0daz1qM8TAcAYwOrSP/kVQhA1Umq0bthAamYcLspWdDgs6ZZwL
GEicanyeaHY8R8iShJHYDEawr8ev3ntHBx6XChezdhWrpJHmYQmsFS2IJ5eJwSWm
RQfbgZ19vYbjnAaOhQzz4YMbzVHQCKjdiIF7xcEmidSWdg4CRJDTkQBCEi6Qxj/U
perujXIU4UkKAGn5qT+/EDYmqzzRaqv05bHtoXhKcx08xjphZMljI3lg7WLxSlK5
KaxZBteoZh2mllF6PeTTtrnSWP9WqkM755x56BpW4mlCHbVgrcupdEz0TRbk3QYl
qvjw2rrub6w4EYYKQPWlKhahWg03600SFLWk88UsxRaQ/W9nfY2BZ9XwuT2h8uDZ
JEkL6/IeHmtPMMcN1Bpam9Mzad2BdiFy2Dhbg++kd87XsOo50Z1656pnfz+DXdTf
AK0ksw67pSmgw6qjAWV2jRvSSUUOR0bS2Bb4lHu2k4eEdBCio7OGoLoPiEBCOMNx
jUhVFmTIhvbHsHoq6PQmhHkL6oK5ovAnpfI+EmoNZy8Vc9N1Jlxh9+cE1r+bmj12
knAviE0n3IPDzBauG8vGzWhGux0IO5bGBKzHWDbNcG7yHN2pe13M96nzUcrnTjEu
W0FXfMFDM9iV1vNX3KUmbNbFcX02XcBrYvyfhj3zUPka0M9n6tdzSlEd85LyVMYB
/46fe/h37gcDD05RdbOBfgcv8jYfeX4LQrvpTj13GQUmHKcEIyeNznvoUYWJgTO3
XNRrBQRIwLT4T0HkOkUFQ45Or/X+UuqiuoTfkHlm5P016KJ9EHXS+Z4EmylxKzU8
oW5MIc7WZqsrPGXiw+Hwaj6V8ZxCdNZhcnOcihUS5N9t+DK0xS8QOw0V7mqO5UUa
EKAOD9ypmakk+2Hchjaf+dg8p5FNoiWT6B8plpzZ0Ptqal3/RnsisDuikYZCzLS5
iMUY0tzB3Eo9hX0Uay3l+nBSdS8ikd37KjhFHgK3JmFeZGcDum7/lBSauUUJfV4N
uUGVP+QZBycvjRbxb2Z1SdL4T2kbaG6ZEYf1wwJHtcXlaSuXYfw1EMQ0bna9ziud
BEI6eRb4JpSch37GvkPbKKp8Gh/zc/4ooUarGyp+TaYnxgqxSt7tbljlc1/EOT4y
j1IyZIqoiiPdUj6nxZPfyuiEVEgBoKJkRX+Du/WkWMo13sqgADa6xG64XsmeSBeM
JUB/9ZENOArshsKwMHinyGketqD/qGj/WdnVrIeXEPHGNKNRBRGGm3REPPzgk5+i
VQBiCfvEegmrr0CFLcWHdm7bpD/nvQ7RM2+1TZ4qPiAQZqLgymU5GA6qttNasLn/
XPxJ6eMyxQ9oZVGW8kDNkF3bM1hefJrc2iki/qa72JwTQKG7S5G9OT7y2c9Z9aKG
htiq2pvG3IUB8EUm5FvN5KxGz4UMqZmRWzvmgs7eyhkp10QDjMMEmUhRLU+nArn2
R60g1+QvbVghDajvxOMFBUBjMB5kkHXK2HesYPp2yU5i5EWc1EnF3L4e/WFI23y2
cx3D6AwJVeQR1ZkfRHouHGHfvO6C8iErXKK2ozNmBMN885WHvxx0P+lSmY3FsmtO
DXEZcslhUuvMXCt+WKGciNZRK2SWKEztDrgFyXTQh4/Udk/dqGPbXTI8myI0lCT0
vVHYKzimxiKNpMPpSFT4+SN+EmMACZXKLKoG1Zh16oxjyUq/puGVBVT2HHKBv7KB
gRJ4XVUyPc9IqWUJbODIhEth6QtrrDJvs/iztP3R7SiJOFKhOxBfHVKF8F3bq6my
LS5dq4rhwxq6NZM3wa1FNRb+QJwRDgPR41O7WwyXDdRLjrSo5m8rK4ftDQ1dKu67
d8JzXuwaOy3gZTH4P5gFt5UjpwURkMMAvp+G7FZg0tpC9Cwz3zYi4RCr6uuP3mU/
CebNm1Ba5N3ZRwQM1YadYI9PvLS6ytTRYRI6pShoQaPtxANNbmvhWtPTyzeyBa/s
Ex+mAoj9aRrsjUUm14Vjl+J8jM/V7x+pDbPuoSzIgvGDYNTI56+B5JyS9ynaRJLJ
gRgpfMLFQPkTwlm7c3V4bRUqEdVsLYnA+5u2tYHepPgNYam6GJ0iN7mf07y9UYHh
InFOfRNsa44f+Pn9q2wXlGr21Dp/omMnej/h6LAlK5alSLy9FgegsOFnJAmuNK0U
eP6typPaCn1uz4j1N79YOeLWeK5N3m/Y0U0rkhCna7ZC2DoGvkiLDU8ofm+NgPF4
V3+/bAPpZDuBAvn+Fe2fy9KKcveTIayZQwrSTc6SWElbc+m2KxLL8o03VHouNpEy
pz5Qj7tNo0Ab7tv2CW2N2gGuuVaseiEvYIY/eDePEGXPE/gEfedILSU8ADqU0Owl
kAlBPElbi+Oy/fsLrdqQNwaB3Z7VYwKsUAsRrZsAA9A3i5SSUpYgNbpJ0vy/pfrP
MJgLFSNqVZxQ0FiArb0S08aq6juVEonVkqb0sTbBWzkXuRIcDwDkIdTITEjT9oJx
V61c1Xh6hQjXR7I5ln9jhdTbZIAQGrCbjxqZk8yIHmU/tHJANafjvD/3QS+e9JuZ
Kl24suz4YbSOUvLxSAADIT55RaF0pSsoaUcIASgZrZQUYU3OE/QDDyOnCnW/DJm5
tR1tMyAbT6jD9Z6yfGDiydxB+0JNADWXxbvXCid4LdQe3n/7vrXH3pRCVrEOEUrU
kahlame6ov/uJTRNOJ40g6baatJ5cIz+cJbLIJlSnOFfmaUaMbLIrQpx3WSUa8cx
sPYjhQxe6WlLtD/yxUfYmW9e8z86ksHkhQhiV21SULXHZ+MDIZcCVy7HwHPDshzj
EJN2l61Qcr3FprM01jcrBzD22m6NPRmcJ7r8oCwHY5eZ8PHHBo9LNCnUPPX3d51b
fB44h3Dfv77CpyhE7hIWQa1PBM/Tw+vjkzK8nUG5THTvynD8NrsgE7TcS6T4En+d
YiHLR/JGzpYl+CDxhutpt/buAHEY4ute1KEzRKL1SyIpXlQLKqTE3VLNM1dUrGfB
Q/XegN832f14XtfztoZnYMXzCVf6n47x5Sdqq5i6U+QtdnYdo7aFgAgXXTRzKDR7
fl6tjOzonN15gwBkHw08gNK6pju1HSzbEzFd/5N8Ug0/+F/AC9ZnfbzNGg/M/bO+
0+hwZf2mo/87bVXjWsVESHvmXvZLypjrBRCtLED7NphSSuLslspqD6pX6A6Dsich
GjaGCdaa//SftwLRATucyScsnMN3Mat2lorGTbSuGUNSfKkxf1gN5du8WupPv1vE
bXmY8mMlZFhzqNHvcCpsf3ciI5C43nC87NO40f868uU5zARf6/Yxy5i+nn+iLhbw
lgxNb6E+20VlOfNbnnfpf8RRJ/40R6CQditlmApjGZEDtmNKcsQ1m7qQFR6PsMyu
pG23W8SAFAsmZGUAtswaWyHGodzaitOHBv/zI07Dbe8vqhqnrRLijaduOLrju/8g
4cBX45xLK50/aTQevuLe0clNmTnc+06gI1TALCh0BqJxdd8Hxk3vsBQlqTsittdo
1I+u/zOgDlcX9HwvLbD3w8Fn6p095+2jcf+iTTFzy6RhmFO7tKSj3LEpmv/iAowg
c/vAbJc23V5Oo1wbqpFp3YXtV6J4JmmBpKaGzxuvHkiTJYd2SUivBeG0Pe50usNK
UrpHJoGdrOWHKTa6eI3cpqqnJfCOFo1ZBht69W3CuWyHKnRzDZmN7wFWuEFlYfPK
TOIZjBiuqEBFWioNV4qW3qWtTP9GQrYXjekO87rqLeOrZEVPS96kr7MvLhp5gQ8x
9Np98MdqOEzs6Wvr2uh7cS+0/Qv4K/QQaU17qO5A1l+Z2RN4Sm81kneZYwfxlyv7
rbuepEt4K939Z+P0l2O9fYVdexk8+OlMe6Y5Ahw0DExbarGdS6f6gIKbLgMNXn/g
nlba/yF0jHFjuXjvEbV0CNUyjlSG57KJp0tdZiAU+vyhzi6r/8F6MDyyVhTHWr5s
C86B6T1P5lYUFqQ3DemTQo0iBCfN4/lSsXUFF97hGrISfnhiokJVrquM6uJnJF96
gdjREOf30vWhZ/09A3dWlEZdqVbUoBAxczYkfmVtrlUw7VOMarv0bf2oFOWLaQNM
1hdijc50ufnLph8as2HkteLOBJASYUjoRGwa70gjPfAuPc3v8RWOk5w22SkLDv0n
AETV6N/5jLaVkXOQE7MaD1cSL/r6/zQpoUrIOoPBwx9wvV8DoLa4qALAex84VipA
Jvtz0I/VYBSWhvwHxNInY/FLsqdeMyug2fKpEVOjHZmEKvMR3bdej0TRa7sLAQwN
WXiBk8CTb+oV2hmV1d+7Adxks1P4vP6uJgqCZfpNDj2VjPlJsIiFBgaTgXHSCgo7
R0Olad0UzV2ec6h7EBK0ImZIuO6vWhHgXvtJUFO2eX35tWP+r8HycMlDEQoUC4yc
vvE9K6nnYJikHsj9CGPBJxgS0TAMFDhSMHUS9xMeYGzfIVEhrm2TCjCyoTwFWJ1q
caXbWyvskHNFpkYYsIN/108u7P2eszOg1hUG3nc5vFgMfC/gBXVL3GoAifc68n2F
qOQhXQvaeX6ira17VtIOin+7xJrad0wwUuM70pxnaTqwGneNwvbe+JDz7haZYav/
sDLBAgWKMyCOKGR9lMwg6a31XUbY5gMZTM2wLdt59W+BJI9kf2tU4pJSPLc6o0zk
qdUKVNvOcGXgBkKloFQRSQ==
`pragma protect end_protected
