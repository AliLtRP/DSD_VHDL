// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
nVUjz9sQJv4BAqNqIC+w223ppxM3yK80WDkohvasm+7GGWSHv6TZO73HTNoDUTWbiVodz3kM192E
FQeXcCVYX3rh6EWLpeyWjouM8szsXj/AtKC+f459Xlu3ak+c1RG2wF7LyxejbexcBfJDtqkBe8TQ
1WF1hIDmCekDUEFKlG7RR0jqsoxynDlHzMS8xj+TmL9G3Jlc+9RtKZvCR+DWfDbpvg+BzcNBBcN1
aMyUENxilpSB6nsgi29LYz23F5/C74sLt2I1j/ucy6YZjNZ8qFEAY/EUy6CI9lcglExboO9RXlZf
TE423mKg+rtNLImJDYSIyYw41rSut9OHzBv6yw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
TcnTsxT5u+BWX9/4GiMVGyZvVUXF7uVPY5PyKp+cs8Q4jPAQYP8Wemy4kEBJIyQN4s7n2J89eR8L
dX+pHovUv/UhUWofkFGFipanyxpdwCMtxsxHqYr8yj2pJt6MTAsJoWaS4Ars7zjL8GOKQYXMHoBb
yOjeGRwFEbc59Z4I4ekjgi/dTAEVrHDdYkISQRmLGicKxyRgat9t40abMZsMBsjsael0VzBZnrh7
0oc1xS5tZUKFb4q0DxjRC5IWbluE+BjoVY5j1gCxchaNLC5FKINS6uZBEa9EkLxJSLgfVWi0pXaK
bRpRDuY/qNzlZnrWnfHzO00C/lctgilrFgPgjKnDsjZPGTx6ghJq3cvpAhqjaWvhk+FCEVN9YHJ+
gCl985+rzUN+wIdOGGNKNImFFInmJ/j+8dIg3SGWPhb0CTSAz5ePZnjBmfF5mtJP1scRsTcIALnO
Ukb1MOCVPj+3PcgEqBnyylX90vMI3MYIVtftHWAkotDEoDdxR0485JEP6NDIrH9UfZFG0ag0KzG9
DrYkrQYfdEH1Kz14uq6UJkN+HA9A5T6fpU7jGCCdVLzB4TWCRxQpCdhtLrcgpp9rvKBRtGXcFITU
gkPD2Jlrvr8795WrUXRqHFVCgcFho93PdSdqliOzIVWQc/UdGn2Cw5BxVCZC6TBeC0RxBOwhC2/x
2aRB4ZMDqNUl3pbRFxmgS0NxcOlwwTCLAPfmfTR+JKv8+qZFtqYtO5dCaPMDHI6OuveNDt7lnr6H
bcJxm7/7+JrwQleb8gokEOJO1j5hBSWtxbvH6LW8eyr0KgOb9ZrXkKyowJ3WkrXCMDAHHmhFl7wc
qmstGfaBKqtGQNsCbSnGU8It/cqX/KtI+xRzJxk2lUwedSasrpDam1N6x1QJvJBj+aSQr0Xb0JN1
FnZldtB3mMnVT/Yi9nGe0WcJmG4XwkQ4pu5x6d3iY603MfjaBgKZQetU+wnAlfIVbuczlYRaSkS6
NsPJfj1s2FJDvp4qt5iXF95HKxZnVNo5vKdFvusCAg8BuKDQIOqJIV8VxzEXCu2+ewbJPu81h2Cw
cUzc8iaA2J84R7Rs1OG6BrSbau0YWqqClUv7Qwexjt2E8ctD08nBebnruqoWeY8cSOw/FA9/drD9
h5HMUOYdPnnGfIaGfH6xFerwIeKdD1znYuuvzhxZLMOJGbwcntx0Rm3+r3g5vO9daknjYmWr+3P6
BZna5H7NAwKOT6HhMYlBJOrrLTylyDqs5HHFjA8hVuvoF1TyFW15tm3OqqRA3pr6DIMpQ6A127Il
37fi9cKoKPFDB6Xkf0ubrid1p4vpj1Oj4Jkj36RyLrZya0dOnnbxrEare3njMEdqoOb59W+h754N
aUf5hSH9vJl+axNg2WxBZIsEQ2KQTra+dpAmg4MpcbXJdLL+QzQsL/flRPVK2uPIZk3UzGQtbLeF
PJS/2SErhO0oEXtgUfh2AD231u3Z6mmt0L7Iljn8zE1DLePyok4jAYn4nOwn8PCYXB5KcaARzcv7
+hLqsd/aEYQw4Rde7Z43bWcyRv1PZ5qYcnosAFliQZMSpxCE9tM0TGDGe9VGPqmPg0//OU88MLoq
lM6MfGZiIaumCN6vGJ0Nm+c0SUbYwVqIh6HQpE5hfV8z8Z6pPOHgWE6htya86ICtxsQnEm3hJnzQ
ECZ5bTc3mT+mp7Zi3Rlu2ZlR3Bdb1L5K1ha3KviKmx1T5DiVn/yezIKjEhcEv4JGh6Z2JomYvGlg
+G2YYHxHhRwPpNDqW7/8U/QZ2fqdzdMuO0UlRINqsAJ0syl3RXstNSpQt1J8ZYquHcWNhP/LCRHK
ap7UHlCY9syRTVdxrFF07HUaogipCXda8pGhhIKNYcT8pIdnmD/1hfMyZ4608R9oJFesSqjiS7GW
e6oeaTFYc5eFh/XkfMP2/VZDEDJONeTjykeZYH4fry4F3/SS2HlZNKb1cj5NCmbzJWB7WqQm86y5
0R7XAOF0sK63cHCbjUWvu/0hmklY+WsaKqHL9fZe38MlrYyfgxNDnd8ioSg7YVFunTtaiMMEnmVa
bUdGUo3ysZqj6VSbmeH/3sjSU99o9hHGRsLbfdRq78TKwEwO/CgjoxGB3sAIc9EBFcFXOLh1B2sl
Ib94nSx3ZOJYu3h8i6Ia2qQIj3eO9ba4ZStWu1eRdcyOwDEvLsO/ldFgPAWtWe1ELEe0d5ZPe9ZU
GGM6UISa4Oz4GSjzspQtlh/mxLFRxMOrnbumgUp1JVVvJPpt9fXy1TRbwwUFcXZupWkVJSIBnJZh
pyF6U135MDgRgmG6mrllkWtc3sE7A9yiXIJxPNn7slGsBAsw1nJdhiRc76w2UO91BoDmzik2jgvT
3KcfeokAmydFzXkpfZz+LXXPaaXu4ZWHiVNNvTxstxpDms1+Pi2uNPtlTp1vm2LHQxjERqmsm1q1
FAclePVKSWGpyjGhZ0Hwxc0WRSydBhEgO2E55LJibCqJYtXvaxAvtxjc3ewJYTE0reZrnGhKYAXD
uLByVmsFsRTDSr9BJdIzelsNvvV1lTFHQs5SrAjEIwf/qx+BBqMjd5BnJlAZF/FllGIpXgk3ulJg
An5ceuumMk7CV/sNB/lfqHd7qDUUQjV7AGoyon0hGDUPSxXdNNuo9Oc2cJAHVqIr5a6keNb+d4qu
Xhd7mh01+IQfxqKRy0pgqmHqrU+hW0x7ayfxUsQqjBxuHUetXjOJl3G1JouQl2BZvCyRs7KxFj34
P8sn0aa6gvG0dMaln7nKHK8Jw5U6g3ocab2fLjwsEgry3y0IfRf8D+cq8c+KJDPfGXrCn2hvT3MQ
4wZApD2DdxcnCfscXyGOO5rlkTbc8sS5jVVAFwr0GxUZ5ufVvxXJqGM02Qh4Gq83rc7TvUkGtDw3
VRV3j0oIDH4god3o7vBgYoGSCNCveFf4IzcT9yJuwXDpvSf1k6xhgxIEGM7hIzAK2M9mJ8sOd/06
829AZWjquanG2dvemOQqVhLM629u/cirm1iKL2KEETkpOOCBxGswZO9bKEctvuyvr26LtM66NU//
SQ9Tee/B1Qk9MSibio2H0LN5HwzepJEJRQ6bNXhBHOfU55eAAbNd77TP8gDDf9+3t9ujFnfNRfcN
oCDaGelfnlLosI2LHo3tq9SItl+toXZrz+02WGCgV1EYFjFYkPAhwpLr/TP64807Fgn9VLD09URG
X2+HzFrFvC9cVyhn1jBEHRQRxhqprb6y9DB8vxurVA8lvLM7OLzcgcCWIfir/UIRL0Z92h+X6T5D
DC7ztYvqrJK35xwXa53Yy2DQTexlEfQa3i86L38E3+fS1aEc8rIPt7qyHSlz5gt0ykzLPFmNxutA
xDDu7ZeiyErSLDMIrXgGNdZu2rpe7kEvH7RklLSLEgmggbiwPWA0ujeUNP9zGbtucXrwfkALp1/V
6MSWGvOgzzBqXA1UFrJ2n0uFXzHHF2YliwpgVV87vE0S6m43PEbaMHpoXvNzgQPV7cc7TsTETff/
hNzweZPyarkIB1w+/6qrEGNoFpnWDu6XyuvgMTmQuvpeW7S1sao+BrkjFiH/wSWCbA/UcGB1TEGT
146FhdJTQ5W+BxO9UERvBhgAMDBA+Gnju/xoopWa7nfDx+1Lboja3VfH+lU/XMLEWJ9UPcLssk1C
iWt94wSYCKfBPz/3zjJClPl+AwZtNnqGHuhBozK/Y8n4XlrAulWn+rw5p9kjLs11DuI8d9LkE3UU
NzvC41GVwsNOgP1yHuWy4XSGI3BWs+emE4aYD8LGhX6YFmWTt07fStnOew2wOab3fSF5m53aRrZ9
KtkZGNOHjXY8piFTl/QVA3Etz+TvAyZv+aXZ6E7nw3wiEnnwiAvAN1q6uKW1W0lRPR8AwQ0itFoR
yP5V7GP+2VcqTPbCQivTAYPD79X2Kwgs2ArG/k5FV36KtW0De83TLVhF2r5A9C0urabVyez7lW2l
AB8iqR0eH98DgEZLN6jcBSZ9C8Dwgsy9EneTglheWquiaJATyGlr0eK8ps4/0nw9jrgLJ7Bi3l/Z
hiE0o+jbg1NZ/LkIeFC4ATq6nQkDId98+tGuRHq78idj6kwJKgR3DvAkjY/7IrNg7UsUMFCvEM07
J3OlAS6fmaSYmSYrtaP3nOcYW2N1e17aPQvIl695tTtvFM9ug2YP+EPrpLgRbqdf9GUWgMX9616V
tO7LnQ75luCIz6sFAprOqqWM3DIXUPucpVokJXHDBPQRp/sKpYtjahiMqMfBl0uyEdLpJ6mTS7dE
+dlxf6hXU5UgIaC0Xjpk26HxYeYQlBC/caXDdYvrn1Qkh0Nh4MX+4fuDcUq2J9QPDREUhiFxuOVm
4QKwI788pC1cDZ4GY3BHu/ilkJmNBMTDugskIDLPo7pG41rmJ+G/st+/CUt6KIgdDaC+0Npsq5VE
xZ8XD9ZqeuTQD1AO/yZGqKK52OK7fCsv05C5nj6a4Bk8UCH8vgupAH/M2DTRJFIV7gsAf+LhEDVu
xsdapgx45+Y+wo2pfzlrCJk3/Jpxmug1xYW/BnHeUVuJ5sa/e+d/Df6rz2Tg0mNO4KVnr7JK2ylo
pHaoRxCB3PRav+IBfEosIYy+JBqrACksr6MEf4x1J0S1GN5gSEm+zrxlLHLFpzpJz7j7Sg+JkCjh
Z/cRMXvjuTTzCjNc2oBwoGvh9EZusYuKYRYbYkVhGqViRlQF6m2EYE76Q+GNEyu8bStNkC1NsCs4
PfHD6zILd0pxSPdBAULSvc22qncKnSwvIXRnb1hhdw4zAwg7PS+fRdrvn56MlpYQ7SHC5CoOJfVF
BynEo73FyW4bjeGndpm14gZv5o0i0zxqq7sbVxX6i6Kv8kGxyhRb+Xc7DQrE4V7jFZEav/gpungI
+rMlX2xqGPKPCBsMp60Z/yshAB6ltfA0NCCRkyH6FUe3dl19Um3XehuJvKeUn06rHmLTgw21Flyc
8sk2CgH6+EtSWkucdavfEqIZu/xDINvczmpcfhBnuJ/maCZm/C1XicLqtD5t0QbYbZeITMck/6IE
itp/GC8Ab2DxZ59+GqrOp7PB+2H0E5d9bj/CpzJYEipJ6CwHfxOvVGvbFsSPdkSGt6RhJq6gzO7M
uVJVTuZvoJim4Iz/edbn2N9C35R35bqmSMqoeQyDuGagvwHITD3PKgVxpKT8tFqN4QSAzPVm5+IR
0wX3Hb72IPI4Qc+QMULu8R17XE670Zhnhm6YO0AfHAM8ATv6w2OQYh3AMSvwaWU+zCLuXO1Izglh
zz6veGw6e2FfAZj/CEd/6og09rKAE6/Ok+0msPhSF9l7UmTizLuPelIyhwI2lx9BM8BAKRjFfceK
/BcDAPhmUE5ROt/KW8QR45oJyMmQSQG/0Vvyswu97k792SYf7f53ajOb8fn0R6A7iO8XEAEp0iee
GNnocRk9bFtKQVxtHA8Xjrq/x/g70lqPkqEEI6bmTJ0KxL/nE/bXTk55UJhle0NPkE/rSoL9d7Tp
pOe5frEQ6rKEQT2LnR/ULrT7pSkPJr6gm6molbS2boF+9+5K4tl5AFC8cnrFe8LIhj2IeOtb39Gg
JhCNnSLuefTQleWVfhGd/o/ZD4e1skvZwnmqBa+fkBCHBPorpyQ+0WVSX5OKxm4hYV3fIvauFzyV
VzIZW6y8zsjVFs9Lfnk2CeKvhtEpQOpnHxg8IBQ5Se06hTzgA6vqnCrnC4mhN1XMcnB0CJoxYdYU
yoK0xm60/02gR4qEGZJ6ki5xzPD4p9kyhogC6Nd4Zb83sJAQ/AD2B1a8NAqMQI8luelSDfqPSEsh
nL3jMCUt0RvPj+BQjEkpYB8JI+beu11sj4bVAy5JZRd3icvi0+pGOXkPVMxFzITiGR90srGYUUbc
/MAEUnNtCHF8iikOKFDqUgmsJhVM0x5mDnKoeseAGdP7Pcfrhr5UiUKKQOUNqs+iYRuU22Y/5/5T
pa2SNAlflOWLEq3a3DNkWLH9rEWs8/LBusCr6+aYTSV84FGS8nVYUUfb9MDLvCcUYZm0PxcH84ly
/I6mRsLIH1nzvKRqArWl0jomIotrGELKPAbnhwXTXpU4GNl+4c6CQBYJ6fplQa/GkEuS2uGS8g8U
AGywe5qs+EUlihyB+P2HU1pQV5W/hoFdYlJtUUfVZSCMVyiNsJVBjyz4Q+rcDMhGhdb4AU/SH+B5
xAB/hh1NRnaXeM89lfSN4ErelFvil77foRbRh8dJTOZ+gczLLfWDrZWD52LeCqQRwTJfovyaRosU
bNGfBMVCNK9cKsN6CUVVrGJaYTTTPHrG20WjfJYzyU5SrFuWTQy9GSK3ovB2uFnoCWESxF29vGb4
F4ahrtF2IKVOYtyCsS9Bd2b7hTzKif/NsExtDEdgnbU/HWI3q1V4C2v9e1tnllvMrvQMCtD8IJc5
1YJV+ymhN2yT48lT4qMFvDWnMbz3Ay0P8uHd7HQBIMgGbL2NQH58jG21lCBU+1lSU0j+YzBVvPp8
bYeQSkB3suQSz9tlaunz3RrOJqw5CZev1ojwcpwDkwsgD+Lld9gBDGEfrSHQo1ARx5PD3RdgMVcI
qk5rEqfoR4l9GNDEMSSjHBz2BEa5OxC+Yy81Tc8a0bpESjdvNzm0Rfjud08jCRUDTyeX8+fkAd+n
45E9Jp4G5BHIml6FuJUW/HPTQLUIvT5h/Ap1kPYpuqUjL9WF9bbBLXcelsNZ7nOvE/4/BIGBu2JD
02izkQBX31AYf8Oh5gVseFP/6fZ1NxOJ/FvZ25iEjmTWgmKlXSw1e3YULNu5dok/HNFC1sa3X91N
SCcsmj+/AicW62YziEswwKVw8cR2mkU6s2nXHcFqYOTOSdviURBeZQbzelLLsLV06Fwcr7BopC1W
wr6abydpToDGAy6zmG8yOp3CwLAzcyDWi47RtzC4tZYxhDdjj9EN8thKHQu8x2mUnd3tTBWZ3kb2
8VS/rJ3d8aVJYw+2Yc6uBZAe3fQZGsfzJi6gP1IqHxsX1gyWfpP2Fc+PODJagnwWDzpKyx/CUKEN
KhcY/5pCQx3mSZ97ggcAnAlGopDtDOH+W+R4+eQaIRsnkDGoLr6SFGvArESLxZDdLw7XaPi5QExG
zT1uW5jHDW6i/ShlBJbK3SwJVQR31REVLPF/3KqRXZBizA+h7k/rDJ2i4a4yCkklI40jydkU2I8u
sMABf2Msz1ZGIie9TLdXHdxhBorVUoIOvR9+GjJ3Op1t4su2I8/SByd9AQMCU3Z5GcUBHzkHsbtV
lFXDiM9k7Wq88MmhDKlcCwJE+gB4rabl7CjcOhNFUQrEe47FdGirKjDvnFmMf5c/6F+0FH4MHSaB
cod4gvvjL2IRUyHW9D34WPrDsKxkpuhdNw9LAOWGxKmEY5IdLdKC+8OJASmXVY1EKJDFaG05g8iX
lIo0UP1NgCaFCmAGyDZX48kIiH8PTnjqvgtTop6+IR2jWEnEOoaAMCB+auZy7NRhcLoeD5EmXs4J
ukb2kNazuZXTOVxMDg8gRvZUc3GldVtJMoE4es4S8nVcgm7Xzf9LJ2OYk232RzaKmZyFjcP0R547
ZIHN/BrjAFPmcrPwmGAt60BMPeOnlAorzIIAcxTEjaqVXOZM9+fiBHrFSlkI5QDu3DHmT1r4TNA1
ylzHqAFHL1z0ZSLujaaBL4aRi+71lzouP8Q9UdvJ4sO1WHaWgSJX3eR+4m23AzMK0ZZCf8iNMVI6
EbXavKeh6MT00hi7zHhGW5iXbeyb/XGh2Q7PUFxy/GDpPOJ/A9kiC1LKjsvyDmTIjlEIxDVH41CW
AvnM7TvUO37C3UXSNi9txdYysxD7+fvxEdrdSllgEP085Su2WgFFEaB3BfAbAv+DKBYK81pUeb9x
KgV6q8xNWNDoCqECqF5dHhoiAsmaw7bPliiA/6dsSZJmHu422txWjYsvALShF5mOemdysf+xv/DW
liFKpqKs08CGZ0z77o77vYTh9uAayejXhhiD0PKMHL8i9Y4Edxa8UNbfLCsiPGSz66x31nnpuL+m
noW64oDZZk3yFgJH8jrxxRSRHgTEupgSIADXyS8r+NUOVMuv0rgN30JYmbCNszc9X6SIALj41j8S
+2bWahOHy8x0vlAaV+u+pvghmc9OQdEQQ3DpkjGtkESxqHukoQs74HfygU8I8XJtUdHR9fAk8Vx4
AcDMtpWasStM/UOBRRle7mHEPJZRhGRCHOkBUoCKT3kXotzARwZIzJI15Z/vCGHxeklK90uFjO3G
3LeADepFQ0OyMJ4AInU3L93CmJMHlGhq+kEsKwuoRwfJuH91dlc+k9nLWWQiqsDdkdc0Ow3KWL8I
7+5r4Rn59CU1tBewlHxXdiyU1rvjnQ19TQxxp7uQ3gS7rr02ortYSptNRX2DBzUfkq8/TeBUH1I4
EsOO64JLayKBzcY1FMWr4fCU4QY8S+xUb2uVSJPqhEZWM4EHjI8iEoSx13ENOee3BEHSnBLpCxAl
T7iOmogAjr4EHeEBWmGD86FvTAKFkzdwpUbaYM5i45Bh/7nm4F5h7Nr95Z3Y3DDhnxHRgnJO82oL
WD4L1ekMYBzmtgI1oMvAdpLsLXbs4YeTbKa33nKZb+cSzt5rkpwZJIcHzPLFDIMUih8Jzzi8fZje
uf3GlDx7/tkBRrVyJHQRxcG8K0dqbrVzrW33zfxPtq4olreQjOKesAHATsjpuqiEDx6v8NmvjJRQ
xNZlUiECNmEMigzuGlgUi99ZgSeRtk4FF873ypbKgNS2F9tGXY29U3IDyCEXU0bF88DgoEyl9y+N
tPY7H2w/YigtbgdsPUuqVnzdyRMCy9jO/Iv43zP2VZ0kXvbk9ct2WKNYfA89XCm+Ao3nC2vsBIdZ
5tpZRJQkZZXpO2J+vbDW676HhW/c+XOmPyqkOqJdk2S+OoKK4wntOlbuq88JFwEjKSCbhqfU4wmB
k2XwsdfL5h1VEvLmor/RO1Yp2tAPDjqFMyAkWSo1s+wkwfeWHJmRPJbro1HtgCkwNzqgSImp9MWG
3aAPeOS9FzeOAzjksEnk65Wb2i0mPtQUwDum5SWNnir5nvOvmigLggmd3UhiKYMdOz6q1vwGxac0
p192zbnt2SUJEbC7ARyQQNOvzlr/TqsehKGKrI0O70lUDrSQaVnVyhqTovjzAG/lvCmXm7ZQxALd
AxKhRuOuRn2OLEl++WC+03M7N6NhdBfq5wApvSXgsSd1/2/Eer4KnSO8yE9edc5qlh3iOgRGJUJs
zYlhQDMiH22meXHsrfvaHtHu7MJl4vBM1gbThMk08L8N8ls5j/aLNesQ/MpjItPI5ROnReTn1zJw
Wj7T7o3oTWSJIHx29njS1VtL5T3KFeCIsR5gjd8yin/54E42YE5qmcZcUs96ToUXucGh1ZNppJDF
3KZdKtyPD8TML8oPn2SW5mDVfu6plxKIUbrvyJl1ydVfU+35P1Nr3e++TZVIqujthAE+EMRiL9DP
FCfFcCJxv9392iBwzu6lLTH7kKOP9vZqzeKervPRkFRVjzJNxB9Ohci1yurtSSCjS6DuNxYFNBEf
STESEm0YmaoqKT6KOe1kfzd7Z3DPY9FmsU2DTnAsqhRl5uEsXV08GiU24HY7CMKaKdUJWzPMtka4
oK4r+5uzu4ayc8VlHl8+UfHdt0FvTWgnVML0DhT30JbaiPus4N+OKAKlmZHnxwLknFVwmi3qoVlR
/fSG5ZBwMF7T0z2OH06r6FHRP6UWnmGBVS1xPt17XtI4n8zDUePyPnl1hmxos0jakL9zW8fwDWAS
gJ6CtwFgvzVLb+VkpqvaQR170vydC0pFSpBQcNb2TxgJEjwqSRhIQtu/nNUX7qjhKfmWi5A2Ozc8
S9HwbBSMJjtPbgzk5uagPAXlaNCvpP+cT30O4ap4kQCgWBmbPvt0x+sWGLLcPSwIq+t7zcINOg8H
XujK7gt2+273XsmL/xefaHJ4ILplZmuh4tYUi0C6Nxf2pdWVdQ9NRgzKfRy3tCBHYdqBlvzWVbS5
W70HnPxkwXRiKngQfRKgjGuEZNcUb4KwD6RgwMlEyKtJNwa0AN7UM4Gc2mJI4jVifLETCFW8y3FO
9i5gIfsM1W2Xm5rQAkyYkvggFB+H1GlHrUETYge5VXIzv3gIAaq7NMRbPX7BeNi413gxKkJeRnx8
NDZ9tZc/JPRr3LbD/9efKZYuA4KZsGVXhVi+AtBAIGXh3AOZNOsi4Hd5LvR/qK86iM/MYHgXA8j8
/zMHFmHcdR9YY5BasO/vGcJPKh7xUJ4Uy/M/4zXgWEoMOmZe8l4aa5N2m9bdprkI+U4ULDZx7YFF
usTNP8391TvXwokn75LUUl4D2k3/rE8ek3BqUsaRA4PtK4BSuiV3u6Yju6It156rtwHn3p5Eo79A
Bb1cIj4CJMe3xKXKEz37tSX2JBe2cyW8VwDyojrH3GO72Q94IQyin8Q1n7LoiIQS5RPDEG6FeJq4
7plf9KHCYzEFGyLTTMGfOp94lGRe41g8IcdfKNq+PkCgryIUpntxC+9R03EXby2qaBgeUklU209C
m9ZNKlOGGlXqrjk2mRjplsVsJ+cWwsk03WCCqepiJ41t9n9l+wEMzdVbzVK6nFv9cetQvpHm73OS
ZDUXxtX2jgfiQbOuGE3KZ+pcPjgzYhFSyR+rnXEJgJYaLpdUV+VnVGrUaaUPcFwIWW3SgwNPe4Kc
8KySq0k0hx4pIFRIf4eVSi07vgafZUuI3QpP/V2hqvztCmaCPE+/GNqwd3tZUTfcVZKSb0Tgn0UB
84u7ovTS0IIc3DZYPPKo211ahP1jt6HLhCasPfHz8uY2RSyhWF6MY2A4IhUi6bDXjy40wJf2DySY
oeY=
`pragma protect end_protected
