// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:20 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FxUtGcsaC2Tw7DXobF29Jt9F/NLlsD88xDCn7E1n5/fkqD53Wg12Uxn3qYqTYNZq
yisfGmf2xJAMS5TH7hdwnf96jIfjkfnqgdUnnRTW0MH/0JeoW0/9O5aceyYxace5
ciKjj+dQIYT5JwXKnjb+GCL4AxWg6mP3l4det/XRZh8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3120)
2GTnYjrFXcCZmtLdGnVd2T2QFMltKPMMmPkmvEFriMEfHWQigi25txwWb+VZGenR
dmxgk08eQwfo3Y0WdMfDquUgL2tKDblQlMLxK2QQRrmfd2l3eg2ZoIDjq/2YvNwH
+6v7Eoueuu5Bkpa4W7duwSutm/7NlwdePValHmepQolX49IS7vj70VkTU+WXjsiH
cKIG1dXYru8jFMdn+gon9UrkMp+oGPAUkQKvtzk8Uh/wRTdawS9EhhKIjzuNi+Q5
EOpGcMwmxGuPRGt8rGLUkhufCIk6tMK1GLznmkRu1igiiBoZYXdh89WXp9FkJHhJ
xFS5ZTs+8t/egsTk5umaU/GAjtuOvJ2VFZDV0Tyg3757B/RWIKpQq2HyC4VMUqHZ
Rb5vyUfSWRYJ+2hLotZBhdqRtKQbqQTj1PcaoxTPXfGyhtSjQbaxJZN0VXGsMhpP
ZKzFrWiNxuewUV5b2HiqyLYRPzcUQu0dd/3r4EStnAykI835+9d6HMhEZDfSA0t9
+YDE8aOBv+OqtdYRC3NIp13NRfAyWufuo90VtPvVbXH4wghiEoVe66QH+1aMvt5c
/HUZcOa8qprvkLS7bL4FIS7JV8GfeuQ5YQSxV4fkZIQIafwYgNrIUd6UsH6W0/jI
tnFkCWyMZE9CQF1dD+BGrzms+xIs7Q3kse8gsQXk1KMWBRGZaBJHaWlrq5WNw1kT
t08T0ah6D08j7VFci3kPy0f7OiK/AP025YFB8FYGijNwBvpbwUWV+qjwkG8QZxIt
bMPHI4kmDj5TvVMl09L8lJtkv0C70S4zU2LcNA5fHVEcoWDTjADRjBDvAavKRspa
uWYawVnOe6VR1Xo413Pa8RWPqI3G9E13S9eMrDTmqtxL4h/IyFTdLSCPGDHtW2d6
2mEXu8IWjR8kVCKhMgmvGxuQIdnUrrRo4d4Z5zhmfv0rZZRnHi6h9WlxTtp3ASVs
O3ADFtogHtqJcTqyaAjBYFMuZsv5CkUPoaIFnBl89YZmg0KJoHHM2O73OrayUiik
pu+m2Um88cQhXuvqAlJiJUM+yJlLTcgz+FLv83s42SgkBSuHF9GnhEVfI0Ck91zZ
dQJlm7u85/cgp7IiK7hW8qF+waGnS5Po14RXG6A18pDhN/YMNvDkl3MF3QaQrOdD
cU3yWZ+ap/I+woQyMOGrjmE7hQ/pzlzPj0rGtINpfI3fSZGuT507LKHhQkp7ks0w
1G7Gup2gXMvg0aJPZ2uRSEk5hHPz0b13WAwI8eYM9wtAcBeaLYhniJBUWzV0w8w4
TMLOaQcNbySkwacd+WlkKDVS+PajhEDCJgmofYhSfuIUK7noVQowYqo0oTFZ5+Y/
qFAjvHUXHWwKNSvlPdkQ/GaZNT8WVXpq8TLwszi/Up/X4sE5VcocOWQjTtYOAqJy
hcycgV/rwqNU4MlP5Uh4Ta5uLnUajjSB+MIBC5nZoaaKvQ2cdvEUVebf577o/NS9
Om/Qt80PhqFecwnkAQLb9+KCqPvvHTd8UXUJwpMqiK5YI1BmkOvM86eovVDIxflk
pRfok62QIiDMJTmWmB+RotKw2ZWq8Q0YoJ33NUvKW7bkH1OLoRy5ZA7FailJb+pS
mzIK3aTQ1/dqK+IxqZ2vo4rCvU/H3hFVkxGo6V62u3b5yUwHK04krFRPki3H5wIC
mVRk0nMckT1P20vxjeXZu7beWH/Rf4f/S/IaVG+omotn4fhIDqcV6AUbGdKtFte+
udqdpmtBFNktATYUIOLY9TRG3lghPCtRclzj6lNt77py0S3Oap7wnkVsr2eFxAZM
Hq1xEKC7juPetfPXiljI5uDhIBJ5VjaEAdx39ibWMYYx6Q/8MoWhvm63APahaUqU
HwRpC50c7Ou05250rNuIKZzItWBy4Mj8SA4JbO3jNJHZEWjUgHDLEbm91bpeh+fv
3VtOXUBGjqT/PrenbfMJsdKavqWx190d/Eefkr8KT1Y1/r0Few1T5JKLvd5bE71Z
APmDH7zsSWFg/5E+BOyIwTxUZfgrsZ7w6MXCORaSwmDTYI7YLwJE4mBFFcM4rfH+
1+yNgOJaaircDFb3gjSouBHaxXUZIIyEWu/W72El8819ug/S7gfLIqCXyugeXEed
0CdOEwvP2AItf4C+ys12z/7Sid7J+synDvbC5NrEFGwea0IJBUzb48dvoya4G63P
AJcvYl1DAYlf34OPJqRJVK4jnusxVnzBagRPYvQ1mmreeYAB4CvqCSKsOvG3Cmnf
FuCxtjglHIJts+9jm0CGLhzyf/Fw6mN0eMKf6tRN26PRXeck3RvF8s4Z4IPJFliF
AsxuvP7Ln7RrFsKPtMEMVO4f3XUha/KU1X9EWqBRZ5ILnqPvZSBe63/cDxTsAJr9
XWTFMsh30brQwR1yJnXZME0Ai4wJrKgkeFhOh2HkEaUhk9T9jYdb0xKo40eBq99i
ZAH2gsQ4lYgLsFMY0yTYWx7s3VcJCgwFKukY9/hMXvmln4l/afntVihy502JRs6A
tOSS//TKcObpV3MNYhJFuGYF7FhxKVrapA9zGXDx1mAn6SBIVbNoSW8ETEVa796F
PFTt9eRET5nxmDFmloe3ls6/tnsMvzJo8kempa+/LKW/9sJp5zzmSg0O1RbkUspb
82jsaxpo+RA+jPGUDTeqMUbVGR7tCcRlM8WNkJRFiQWS9LbfrLnT+YVgUESaTF9/
/KQLbxxzQqgbhSoSu9p6QACMzVwLh9eI1EyzspqQki2fTMqG27BSlpsdxu+gU+AP
QjSxd1zynQJ0EukspokhDgmrIjyND7N7DXF/EGMes5T4GSx+HnUCBYjCKc5w+T8+
lAfjwwcPOCC08H2LG8zvseTsgAvei3QH9cSG16OivXbvKSAsVV/yJUwVc7PDtZ2U
qpmsAWOfR639Pk27sGjQjGAvoDza/6YMf61k20L+W8yV4qd8vRWxtZNeGDdFbbgP
nkV6tGuRtJzxvL9V+cSMx9y2x3kAZD2F1LMnLMaF8UgOxX1MLgg791CgvaorKWET
2UfEr96NCU915kmfV1uEegFCyVqva1la+RzakstLsWJP0J9qYVjgu17hfSxV3IsN
OJMs90xmflxL58znQB8OT/4r5nQsYozu6UkYEbHRtoMsyy0a1wzpCkxcDjQ6u+Yy
ae3NZsXub7aOa2hJSAd0fMM7RmH6NfPYULqGbPneMhABXMsIl8LH84zXBcZqCE8Y
VsDrcM6OFnI4iiRIQsxOfeuXggYc2BMMWrlHOtQH/RO6nyu60kAn0PV7yVJXdHs7
eRCbIBB/f38cnAq3uh5/7SHlYB9kzDPiyKFv1NaY0GANs1hWPh3nbxddgr5e8BiI
bWxNmGpsJxwiuLJM0QzlhPW9PV95XJcJA4MKta5XoHUFg+aBR6VYDJytc9ZDxa9C
IWQDr6zabeUT78UkDCaVNr9YJgSV8rsNCWAuwu2pMCCJugQhCpcV6g/FvV/AiMH9
bcgZ+uYnlkUiWJvlz2NBtoBz6elJxhA8XJKjqOpyCZJVqKuHh73w+eeSNg/ocLiH
+E0vitFS5p7SKN7/0iviOz4Px1jOJAzm7lFDwAADRPYjrL7qcHVTuHu2SNzz50xf
u9kvQcktUQVjK7/l64oyiPEPPitFyw5/KBDHheoDRrOlc3yB37rNDPSPSfDKJl5a
3usR6jatP0+uiGujqqhKGsRH2xhbOjXLJ4MIYLh2fE+KABBZjglxzoUHPodLd/ZP
DDikAlQHGTZqhIRrmEoq13/cffzmMn879dLui79f86mYTXIFpN+GxIvbnejHmEIF
mY8nQWU7p4gPzcniUDEWJqpwqcGezXjH9EZVlcVPjuwqcDLzGQAIUirOZg9KHpvm
Ywgb/EDamwLcZ3W1s88dHpooNl6UnnxbmZVP8rRVYBm35eUIw7aqeZvYLRnn5ZZY
t+x4mhcM5xn2qhsfXREzLc9KSN8SmzgvZor3Cen4SAsEzmv1wutrhpkmHrcK3GIl
tdNtmsnX7dI5q/zPLrb73JrzJFcwojLOg6Jf6tQ3rZc3tl4mrAPxHAEhTbZvNOhh
Amg44vEU81w+JLG1Vy9cbT98DFBfwAvJjqaON93m3u156LSvn2ImsSfdmgL1HtbH
3XBKNAuDVLYmD7F/oiQ9yRH+0SFdOctewIPJqQx3w3XhFJwdKbX+8RP5tfE/cwqi
`pragma protect end_protected
