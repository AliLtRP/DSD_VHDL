// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aDPgtJ1UKVE33VlSSpiD+wevquYjm+vV0h6VBijPvau3UBJ7CD4QjgTRJrf3P+Ti
K38y7O/EHRicliR9n0jz0DqJIfH5hGTpfB7oKSNEQ9LOySaYjkNIFdMN5+3tAcTy
2ZYF++wuHzmSJ1SY8j9LDglIGSJON+nSUd2hz1V5kdQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26688)
vmgxoot29/d48Aeqnu8quVN/5qbUf9U51tBCYadE3qs4GUfP/tBMJD30AtrHiKhe
olBVz3jcX3QwfVspmfrts1u2tfKsEBvjYdevD8YG2rN6wUr1WfCVl0Pcf2PSe7vO
0sz7ABzRlc7HPn6ouryJ4nCmgucDCwB6q0/YL2fLc5rvHZ3hvYMhpSyHQoWsKit2
UrYT4UzwHG1EwLZPp1X5zKbvBle0ZV+uGdFgOsYGfvzhledXuemJ20+TUOkBq+Bu
jkMmQywzXbg1D+VERFfb5ETjFuAtb2++p9E51niILYEQ50DSQraocLMukX85D/u8
8XU/ABQaEBUFAB4fWGFfXSd9hdC6/BrW8SShoFNbOcTCxsQq1y2vRrQntlNEA0I8
WCTOH6G1t38dGR0QjkwJOHM41eZaFCZ/UozxqGQeurOK2PH/myaO9ac+cH3y1IiW
wJENUBGkx2atb/iGrY9j791rBqBq78r/V33RB4q3CfOwmr5bmvZI/KBNbvKtHDxj
ihJBn6Tl7Tl74JdPtNZZT2dYKCx4njW7fF4XGCN8ecwD4cCpjymKuUWqhUCg39LX
HV3HWokfiiouVb6gnlIiYdxlAldNPib5iZahhlQzoT5kHOnda5aLPJiKrQXhzr7M
u1ufyUDw6iRa2RHain55Tu2gveNLrTJmtFKKPlTOvZKeJIWOToH9pw3CqIvWejWs
e0WrJt9u8ME/9r3jSnBepUgDTjP2VZRe36lhE/5ILDKO97YHUFXfH+Hx3f/8jSmn
HHBXZjIv8lGuyszQ/udXL0UGUH5J4yPgV6RTIvXmWBnjkUde685/XO5tq6PMW7ex
E6YpaYYEiLVwvX6EUFrvajBhGGs5auH2322xB0eu0HcV1y++0fGiMuNpLR+1ntOO
Lh7BlWXRoDyyY3R2vbgGCwp3kft2a5hf2HlYfwUQKyy1rY8RSwhpIy02P6DIrauI
vsuPMVhQQDClpsygSdKVWKg/3KIQcojs79MQ5C2Z+m+GPO3U8SB2umhzvXNxAAKz
K2q3ILrnG0yTsMq5glvjGgHfUPA/GaNpHihYw1EmTVIN3AMZUUt7OyEuURbJ5FBe
p9xlQC4QoSJzz8oY8hUj8qoVmtLo8zP0jnViS/a0K4S9L0lRQmDJl4T2WuOD0NdO
qNwedXmW1yEebEi0+WsIrY9oC/e+SMX6+bX3cqudluawCcMsmO7r5AArumCrTzV8
WAHx3ITiUysrSU3K1RsKYoqmBkedypfmEeMU+YCZu2isUBIc/mSe0DQqT/MmiEzS
RqjVBcvNMaUy4b/AFo+/I4+l40HZf4126u3LqyCJz9CFHQeRkmxPXh+pW6v26aK1
Ilh4dhOE40duXPcBdkO8kTo7VGuc5anyZgZEg4gJW9exLqsfPWi0aXcV2f6b8CVr
oXc8R/xEsSGFXo20fFU2FTM6OYJFzYK/37BVK3yayUcYvgBWM8o0kopY9zMB0oRy
z4V6I3tCs28N8trNPH6/LM2PuIqTeRpUej7bToEdcJST3QTPHLxqN58z4zI2EhHA
n7vWEJbj/5bFSzNgP/Z2ZX15x5i3vZQ5lRqMpuMaf7tFLIkfG8sR8aCXRwscFene
MPWhlFKJjNv83KClHl4HrKx80lXVvsvXwPkmhjlVm6L/j+pc/DdyJDRldCdtkeVr
qbuw+7t8JIAe+sUyl5QpKew2qGp0jaKDeOMO7klnFj0BpueLoiWisydEDef6KCyF
/GsyzxGzr9Xp0/7kVKc+l9pfO8CPkH525tsmsnhzVbhl2PMzO15zORMQDljT8u0d
GPowZPgPtyYwpTDO01Yh/umZhN5+cPIc5dPQYEYze1p51IucOdv48PJhsvlO+BEZ
QWh99mx8Hr6LayeaPnhP1NlaURIy+NiZk/SetzH5FKXqxE8L7jrhL4aHN8lQLkwl
3No8iNk20g8iMbqeqbLR6TvO6EDlI8GLDQA6OV9DwWIIW4S2tGwOOXOY36DsbOVB
lOKgUVIcMbbACi3Mh5ip3RZ7u1hQO9ywrmGaWkd3pKD+5K9zGrZRQq51iQoFqhVT
NWmKu4oYzIuVNgFyMnRVhTUebd2Aq1dReHKASH+yQcPbFuRqjHBUaJafnABLtYdO
WfKfVsnZf/BtdOGuY7nFE2DeHUQL0KyQ61tHPcmzRK+82vYvQ4Up91CAYHRMaSLD
fQLmKh5SpXWmb2MZQkORLa0yB4F0eHRBZ33eUoYG7hDdEjyRmFdtAVfzYAZE0ahJ
YkVjZtMbD//YrfgnUopRQE1P4f4WYEEwO8dsHfgy1wGvj+kFpHpQj7ttWjyGoKGT
K0VYbbrIDsst8QuGCCp8mhZIVfa40Z0FY4QwF4jmfMhgtz8DdFZwq9HbZ95jsHb8
8Nh/0m9ZE0lIgF1rmT+Mv1htu+QykVIpdCYwaeb/6iBqcx5bZAxNJ6FzO6b8MryP
9GNu0Z76KBROcP0rKX4h1Pb+CS4dowUDMnJeQ3EmOl0iBSBXfQetG9CmswtxxGhU
NMNdcj5DntCOGLtynruRb8lFpfs+9JykJL2MeN34j1RH6m6UBp3c9eUuStOb4I//
fglosJcyQk2dkDRtuu9rdn+ulrALFchREQTw5buzo7K3nH+uK23HFE4rV8KgwrgY
qcio1qOr8DeUQ+kKd97HFiYvWkQOeN9zjqI8UAJYdetpaJF+ssOVsfzRjDF8vDfQ
wstA/Fk7eudWe9NujBIVLA4pMONPjoI2eWmxkfaK70jPw3FXZtBK9L9xkF39xrEC
htdzenbr99bgOso5XBloeSeggX4DUQ86f2wcFSOBCPMj6+dDeBzNVE6iAPMwTmDp
mEU9jnoHpxBMworHvg67Cf40uGjtVksRdw3/wWbZkNcvYfaMaOl3Z7QpmqU4COAk
xs/LPSTljRICDZaHaAdA0axkhJcJZA0Bo+U8SaU48C1Hpb4GTTxJz1Jf8n4nBcW4
ooGGv9Ah1VMxdClwpCrasfTSQOm5Bub2eYgNpd2hVVMz5AWyQDtmdU/BFVB2UBi+
mNnh64pNJBq50ao9Vi7cu7JaVCrpIraZ0pzqOIv4hW8iwVBZEJ1FhVtaoQ25VTKp
ODqXeDAbqQxCmKw5lX6ewyc7P6pNTDf/V2OdsE2T5vx2lAEMWCge9XceBsyhECrT
tg+fGSdJBu4gNrY+pifm8S3L1NSLajGrxS7AkP6u2O8D0xe7htflKUa2SnBzrHpo
lr3LR2F6fBbdNwn6PUJuXSctzJY5Z+ChWg7N6lt5FEk2FtajhqSPfNUAKDxbNZlk
OFV1MDo/xTMQ5zDArrcYZ7MTKNMboP0f0XQbAgDXy8Bz6Wt3KnYot2ctoMExlY1G
NhTxU4BQSUUoIm9vIkQ4NAdF5bftdTOeAxhjbIKH1UjlS0V5QY0zqN73FKqbFueO
p2mPYV35KDsSFOqouNzm1sSoR0sOWd4VLVmBjbbe6pG4itNa3DpXaatIhdqxkEv/
tb26x53B07D+KkAaRT2N5o0xqOCDHtnCahF1wbkDVhOKNPJuBrn1E0RcS9hrRNG9
tv7nqwLltUxjfF00eDrl6LqIPxog0nDW3HerI80kaqJhgUwfpqlFfxknJ1lPx+SV
ajI7sM6eSENT3x9OuwsYnDi6NitBT7QndCPiUfWPYA5f8xdZwHnE4C16t96PAsO8
6yLbqd+b1Fod6vCZ76vz4XGE/sIKmgjyu4dxfrwpq1yY5w3d3EYQ560kmFzXP/yc
FophrVKlIRcuew5wYTfDVUoXShTAEs6AIzROU02kEgECUfNO6LV33Q/uVfP/YZ33
q34GIQjyJOj95gcsoFrB6O3fiV0XTbvueNXQA+b9Nrhxt7VMmrjxSJspWnx57f0s
3uNI8giayCCjfkCaPGMXnz83hbLE0divHvzSco9og9r19URrJdajGTF+c07sJtcU
w/sGirtFv63BvU1VP4RNuSbHAD6YETWbyghWMyOdajcO6EmpfqXUaydWM4DmE8A/
gSYGkhMoNj+CVsHcFXDy1pEWJWpb98tRBmUtY2d+BJrInhZM5cGgHfi96fPt7kNv
PWdVjMIZuSvxHr81kWABq+Afq7Jc7+t4Q0Y60/AyDRRhL4QLz1jDMI5l6R3cv1BN
AzblgAq1FW86RASHH947Iz7+CoSJ+7aVub8ycRXolN7WOZRNkbY9vflR0gatc1hy
1Ck2Zt98/lnOD34OUR4tmDs21G8aJrzQnxzLqxRB63VXt+jPE0iqRqoszaih/G4g
bM2G8DkWAr9HvFTa9dfmLso3VsFUcto1dZnW3dl2Idb6hwvo9jdX16Hlzu8xB3a5
UMEX8EtRPuciCJSe2SlV3LS2qa6+2dEicJLNvi1VGr5eyZPk54DOio/Hf7kCy3tS
FZrFOxMnaHbprWbd4KCiziSu41CPDmRikxy2Q0xOao9xag6IsWqWUgiQMqt4dvgg
LPKsBb4Ph/puYpl7vZG45AVKJPcpEcpbIgyTBZe4+GXPULacwUyYONuNVkrKtKr9
g5kPovSB1ZZP94itTJafJhuNR0vQRdaIeEL9Ab29+WmiwLFUAeo7kMfA/76dbld7
hCfeP/mVIOgnxrbl4V0YbJptHNOQ5qoDuVNS1LYoAl6tfgROQYSoQBuo8URSq3Id
tZRBL4pnlK5URB5kWr48qN4ozz+egNnHzN/vjW/oE2f1tnds5sEv+Gj2XIDULvtW
liL27642stkZm9v6GOS3x2r5X/Mp0RJ+nR6keBB3qWkdC63gCdrtKdDW1SicdlJ/
N/qg0GSpW5LAXeXowj4r5tofS0NZsg20K+WIdy9UEVYKHpN3D8Hkg61UPbKheoSu
PZSiYVnaLaRJUGTOpvQN1forG6+275k8Hnpf2WcZqhvgwN81EESMdIEMotFsS5Nk
0acG6GktpqS0p6EIR5e5W2XJoqvDAo0OI4YhH0LC+YFO5I1ox4PFCue/hhRSkHY8
VPaBEz9bpjoUaiKqJyqrTAN0bSzr0R+IXRYx+Au+WksyekwFfOtTqDJdh86aAXG/
6NKNRCf5dMESFwDeHxYzm1o5agQTH5OnsYCwTTUvtN2p1LH7rEWLT010iKEOAHPZ
5ypLabHz4UylfSLMnBHxjNWjqHY8CYnELuGy/frJtky5QyBbhiwtsf6ipRrb2cwt
cQZ4ZAJNi3/7FiWsrc88rDUKznJs1zmq56HaBzqYyhCalkSiGtfc0TxoU48vHn3o
5wB4QAGHurZUCtqoPHd/b0QUSMxi0/mwz41mZnd8lycs5VCo5HJAzDzHF6LH0V+M
NK5tTEbIQQX2tuEHZfF528a3sOproyC4apmyam9dx7BEgY9skhv8ckq0ATjpPlwS
qKUIIGIXnpOGXbxM98BsIdCn9KMOjhtcSLCBX0GeKXFJSYJsUCpjCQhVoWBlfY4r
UNocXY8UsMO0FaiYG73V4LqdGkCEH1zin7AbEU5zDyictPz5o4qBT06bIUIZIUzh
7ozECL/BnHgpvWYpMrWFu4W9U4TouC37AfVB4BsU6yYX/d7V2yhglDFB6W58CaS6
+rvoTaQV1tnZnSHv6FFAb2N8ZphE+tkYz065CMa3tH4fsCgKwNO5cQjUpOr4gTKD
k2k8fg02azUu2S+QPHl64iI9tBwrCBNX7oE2zAaL4qsUxu2+I/eDnxg8gyr1his3
LfOq2VupmnlN21qe2G7tx/uCmTGWrLfRFBRohxDhYDyPkjWiUdxmdI/JJs0ApS38
NzR5Yp7Nrd/LlHKxpQ4j5xVqEoQ2gbMEqXOuitCPrWa0yosKLnFEKw1C+MLK+KF/
zMh2NEjU1S1pO/gWT6cC4+Y4RJyBjimBnRVRWw5DbvAahNX6EE0mMBLruQye/++x
qq6V43rLCpqyq58lISjcBdubQy7hzzQ+Sn3Ck7LiH43ltjn4M3MKtn8icNtj26WE
wXhPtnpqYWy1Qi3HPDaj8Ke6HZcat1uCwxZ2GnyQ9URKdvNWM8N8MHcBUzhkbWae
cSyTpN1OqmuV18bmFlg3A1CmpR7wOAt2rJJlnJ5z20aFuT3n7RD472USoOPFQ3Tn
aL3r1PoTSlTC/AFlpPIlgg6sA2wMVR+p3bskJzMxaOLi5yzlj5J8ROZWRUrzXq4g
3gtDb4LrWF3RZ3RfRuQBfaQ2vwwA2XMrcOHvuIAhqmfwHJ52bt3A27xyqmbfsFk5
AZilbNvBqmBsqljNJDyVh/Jt/DqEX4pkXvoWW5BBqARtI1cU/6TUFItuL7d+udqj
ljGMDAmVmWlI7NOD+BDeU3QCmWcSzCcG0Of5NCbjwv5FrjgM2x8XqCo9nk8iGgRz
BqSebhIA/re298ex8FQpR1MjIWUSkM+9f7ximpNQ85gxmEPVL2BTa5u3leU3JpqT
AyvvnRFPpeDl9PMn7cLo9WYZD74gaLN+NtaKNJZTOwv8FIX09NzdEta4Z0iC5IRD
mOtV0ahHkyV/J7jdc29ol/kVrm2JcNjn1NL13ejCzmUkNPl6ukvy5PtUwzZqfEEv
7Nhq/UzFD9WfcIrf39IzRqzO9p+7FfJq5YFTkPwLsOZ/qZuTtsxJeEpGLKMqH5YQ
Q82S/wnbB/hxRJKubahBZR1DlAzTypwnVsVAyNvEHBluEq8TWuB3wO13CG0LXvX3
01BLdKnc4cVrS49sRsHUl4VyXYeoJlylqR0Otb+X0nX/0yJ9mLVwq78kQPEcTjQk
mYd0ZF6rkd4MM6mCa6c7CNdy5wlQTFwpW1XvU7KYaY3dUuKuxMDD6jxQ/0TgmfVu
ybmFsGJAazLJddqnGi/Es6vcmcolaKxM2CigO0UwUy5VaTK9YuaIUeVJLro1TaP7
wqKQjyPQyBytJ/JIE2Cc4xlyC9iu/mooaDQ9oL/1G9MHXcQiL0acU20YfQzo1F3w
pKGz4lR1MpV2J/z0e5eccXxVKcfAE9RAt22x/q1+KpHXsKv5REGmXf03k1L8doze
hEQEaJEOsb9jC8CrTZAZn7jYWW3fvDxrIQHFZ0DojT/OxJ8NyYSOE9MunZVLLxPW
bPSk8GzqVFIUaB22NpQ/tUxavLS1NB4mqLsQEj7zIXf7l9lz+ar0ChQXF30Zu+/2
EC6+ACUoyHen1RMzVmyJ9HfM2i2EYajnJPC6PjXU3T8u7EEcZqiQwL9AjLmVIFN7
4rsbou5MnPkXte6C33H2xOAu5m/KSI7PMpVpiFnRJln7xGJIiGgmPx4Qs1tBfwKk
nuMksUhyvos6oEVKkjejydo3ckyT7dabwxUgNhXnVdVFjdHxMrwd7++zzYyJcG6h
YmaUaRDNz5rWNgJWWNzxBWmbYn9c8bwvm5gQeFJlKePMlvk39FSgF0X6sYjGMqp2
uDBxnp373YaIArZZnNlAbMjMCExFthHG2U+N+UySYkhvjnlislP/v8zpl5JTJv9u
aVDl8Yykvk+dbWl035+3P3N+uZmECrtpT3h2rZe4MA/xsxoIuhES/1j/IYvG7UKi
mnPauYrQ3WGFfoyP1lN4rzfLHxUZCKy8OvjiinjJGQLyVyFpdIFIKgMvM5MNccZp
+tmHKWPq/gHW6mLiPpWVqlwt3HfNglY3ATlFP3O6mwmYybpEhRSvBZZ8mzdUsexJ
HTomcWSQ2sz0H2GeGiWPkdJtkIqjIdIbwNv2ES0hmNJnn5cqD25hSTZHsuL42xAS
gXbKTbIfcPjuKFyFGBKm/IkgakkiVrS6gw8Tga3x4S/Y9BRE2SJ1b9eujHGoYDp3
QbWb10fUzT1GwjKFurRiJhQDuUyjOKR6u/JBnwdDYDFEU94aTYu8fuVybSMNDH8o
/5kUyashNFBbjfmEuEjE9wTJtNva65T6pqSU4DObd4lopxroNHyssXH4CILDXaPE
ozT0cXogjev5nTkciJBXJN95ltcfb1I+XjR2SKFclTH2Oq9Z6T2PJ2z7t9gLfaqC
l9yAiLyqHoBv9EPc6u7ae/wcKbNc2ieO5LDb9Y5XnX7VIgjHQ0p2UOerR8xaCTHw
z3GSrjwT0+lvXI8o6cIaxmfrIWmltsKilD17rsH68L5bIcWrbfWhMGX2QgywAo/s
2CFWJ0MemUddM9o0xBwe14Gvc+5pyKdiGHe342CLQd+I9g8pY8IK0WW6TWExxNIn
+hz3LlvgBgEP8MszDmaUTVzFjWZRm/ccZF4hQU6we7RmHcX3xAe9dp6pW2n8uNAL
zBlMVk6r+eRijJ1mEdrsrUzYsa/H+KVpfAV+JVCSts+DiR2hnbFdhIDBoNbssBP/
LsZhu0Tw/TwlGOnO7ToCTIvjSggUtDaCZ+VA2h/FysFieYhaU0MloFJipSEil+O1
JCBZydM7So5QkbGscq4CDutkUIT8fv0dOwrvwrX3jrFC1+1jrxTQbaTOxwfi0Kqe
8wGM7TgQzDPdDPNKXgjXXKKroJi+SAVfrF321n1xcxb+yE7i1gxKPQE/2VQHLTpb
cmgUbQqkDr5NBxziC8Zq83bFHKqE7N3qirflWcOXwTbOD1n4S+A8HaaZRc25hIvn
218ef0CRmmumyhJOB8eMtnykCSAeLvYbo5POa5NPH67v0/PlsC5HFV9tYQEM/kcr
aL7CQ1qjYZS6ij4kx1n/5zRBFEw0SAmUseMApUpJKgAs7tfn7KB85AOX85n3raBF
6zhEFmRtDdyhVkhae9Hb6LlxDUSH5E6OzkI/zKFftNoBll9WqaoD8yS6uKDxUmZy
VcdJjal/S6ScJjKKjzJ1Lnr1aMQ4nLYVCQAz8n8ddGVLAW98Cf9S0qXo7KRuG/fI
LSDCYs4/HSXQDJ/5obsbiLyRTzv9pB1tpTeuElMSU21txClQ3i8m7RXdpMN7NyMT
ZoQzE0/jgvOvBAcQayypIg8j2DYlLaS/qywPTSnhuHodT6V688Dn0zUghdTLVe1a
Vk2ar/NNVbSoI8sjEH15w1StUgoUpQvKIaG5hfhsjlBcY7GKow9l6YfKvqQWWdb3
grUOCb3Ps1jcvyVyJPl0UETmt+G329K/61B/fG8ebq8vN+CdqclczRerNvV6aHJD
CFmE4io/h37Jwqe84erglS0UbaqS0IFnCoCwbHlwVPJroA29qQG11GhXC9LSrXgJ
AzUw5kcV9+GvO8Eqm+arUe5bno90r5VJX9C+cqUvXkeQkf4chu83JKnPa4BIIio4
+ZdhI0PiXq4pBvCvLsWdLpgapxN1YqrrMiQkwNGaFV6760JB5RMAgELLl/ysxySR
jrU53y/e+Pe3CVnMdZRe0QYe7fDlY065PQ9IBJuZZEwF7ytPP5w8qULxce6+5RMi
2FzsTblLPJ7iOQ/JyA58ddShtiCqfVuHz+eXYAphM9mAxFftmH3DIO7/FDtD/AqB
qbj9EGl3mMVcEdXde48pJIGsqbwDOPyRkxg3yEi/QXau1+D4OsBP/lk2RcnhrWf9
emLbH1MEEzWvHhZuLdq5twqxxSDve06xu7MoIq/FqKMS4JcPXMd0yGI9HWK6FKgL
HrPXgkqlwOh45mmYaplhh6b1dd4+c/IfkAu/8JgO42H9k5Hfza09Urf4Z/6WBqJ7
uW1TqclSkXVVn7PC99t3xC3NjIqozT2I8xUbogU3hunrMY3urTXns+uIYyMQMesF
uhWEUSjaS0L7clKRdSWFroSNTBtj0FJitfSSesftpu9k7q69LuUDXLJOYgqJ02cc
EtcQX5bWi+L1d7rv5y/CQ5Uy9XPVW24MaptgVVr8JN6+sHFA3f5AUhXeRP7EAMW+
zbxcEBgD/YiHTjeflbHJR9FcxHOZ1NZW6R8NmwsawILzecJjXfMBuaLKxUP7ewv3
5hCEL+KtMqaY63ZT52HEbXcoBpmlQWRVAhXADUhH7q1/XligVoi77EHdFVCyKRBC
/Wg1kOI70auUCAMH4aQfgt9tZGwVUdPwJz67Tg8eaiy/CF9LULz/PAMKghzxauw9
iHIkgSadwX3o1NDU3/mW21fYYiCMMkI1Vi2WMRzEYAhwkP0ALQo8fiADB3dof6lo
uMLUcya7/E27k/1f81QjWe/F5c0LV51eNKVM1VYKGIEBDe3u71cvtupe4P82J8Za
W2vwvOLEpGwjo7JHIgTgTB/cG30atUmuWuvfLmfkpIBmxahplXAwSWBeXscxMQD4
QRYhyp0NTX04mGZv9gWRGlNVa8Hp+gL0z4ClBiWjAJSAiP6/YjHxpiRbk1RuQEXk
KfBFw0b77+US4VRLVShRoT/gYIGmnu8s6+LNfBMAIzqDBDQcdj+r5NSTskMTFj/C
xNaULhv8QQW2xGIpJrkV8ak5BqM44ZoYzU0AGT2yG1LAUf3nIVNffvTuSZv9NoPA
6+FNRI/VaMY5pDD75DwzDkiLCArE1QcTgp4fPvtdCAUGgf/qSKNFPJ5wpUVzq0JX
QtfoDUy2opTMtzc3yToHoNp8pnNK9PBZNsGf0H4bHlWmWytpCRpwyO8Q2wqjSZOD
S6YrMTwpubBlXMPphI7hI81p3gLX2of4d1+9OTZ5KpQNYa0IcfhIFq9/59SLvVec
DIhHgN1xig/bwtbm7q2BW4sEbK4xQiRZcKgT2VRNeKEgx0c5Z7mBovQ9CKrYFj6h
5b53yU2TJmklyYwYedmG7Lk/qE0UAULRpjCDMsM22sUOSNIG+vXY/Y5kv+A0Rl9k
qUvqcT4LAsVn/mxtG7x2Dkp/kInf+Lg7MMCHHuVtIVbZLoEHdf4Kjrb0j3mZhq3F
J9oOJ+psHnVsz8Pxb/pdVg08DmvYHFWexafcEetlxZ8oFEtttiiw6Hd1oqLZU7G1
nCnMf7sPa3GZ2rKg29M+87VOlUNDDBXDun5T6EpK7Jd8T3GWGfU38XNA1k1Mzfvg
V9FdD81S5iLKYUVHV5sXPnaXw1wcQwGOHUQ0Brxe2laf5T3Wr1inEbKv7soSHc/u
xNZcLf/NMCyqId3wdOvnQLO1QAaiE5D2xehnDvlZq99k5goJVbdq6u94G0Gb9ktL
U3EZuKPVW/nReA3xCkysYzsIK46IBYigJqcNSVUMu0FVBhMIdHmmU4bJfO9gZDB2
HTGwZaMWzW+zDNwLSGRsIFND2lwdciYdxub0/nTwDQVFN0aeT0fqV72AcDiUZieV
NyVoSZW/GcDBVjdZMcXsF/PbaUGH86dCVlRKGVRZAqjnRLuHpbG7XlZXmyojEYxG
Y6BvFGbbLAVAx9iWcTC+9lY7esVaUN6el9feLEFNL9T12d8OhUXwYGS9R4bTsEEG
VuQWhUWWWTbEJDI57GdR3NN9zirupnI9O8+x1RFPYNOhYOJJBAvXeLoAElYpeMOW
VctYKc6g+sI16M6Nitf8AKZHZyWlCyM6bij9NXobARqOCQITQaYDb8T+GAuHuWi5
xITpVnBTkmeIE8yILZQeCTcb2j14g0wmMK0R0lX9XJUGTHpUy6bQSuI9qQlKHaHi
NcZOczbCNth2IBY12BCRxaJ9g1FzZCV5SToIqKu3jyH1R3/ny0DJ8wSXVvFRK2x1
avgdo8Cn8kZCk+H/qoWVhZK7mE4cKThHoF2kGtUZhwb8Eh2vg9oXFtNCvHIRBjZl
57/u8wjYCaNcIOphlq5whQGXueD+G7vUqxSbjCotA1iojwp/BEkUSk22LEivjM6N
7epg35UhxYdK7CS4kLZhAxQtU8GBj1+aSztaw1IeAhHNwyuf54kPffSL9LJPSo3X
CNG5r0DoR9ZVOtLJiPM90wbAcNa5fHjCQo7jL4wYoam6mmEPcpwe4FjGcxZXMwaB
IEP8hnVOTnEnRxhC0h87dg1WlV5PTuuT4y1o/IKTXX32Ok0ZH4jp9tGmJPrRM0Le
PujknAefY3OrQl5fafOvZVmtjlg86iSrxok+lTgi+5DS1DgsytwZsd/M+im+Kpu8
I73xMldcxaNK0fh+UhFvgxsxToMh9JhtuAB05PHAIdm70hLYaqv1FNj+lO/EGfuE
W0XU889bnIzViwvorg+tML2XEXmmGyOmhMTlppM1E7XzefbJiGAUrpKT0el1mRg1
8L87tQa6uOnKly7ZmeiD5fLm6FFzw2ZV2zLGlUl6t9dfbYUEjJsNAtZp57yvFty6
9pGVmfY8lUaJNjBfidpkrB6OLDC8Vxmuh0kSG5bPWLrK75fP1RoZbUUBHjljBVWe
kJ4BvKBxPzQxcWzrhCAq3bfmTLPeFBCyiqXDmafHUQyCa0V5CCSkLR91yJW1gt6E
1XiOpeH100Q0MErTSIrwe5kS325gUGtVKaRyUu537kpbM2W+w7auV2wv6qGx4+Bs
P/Xu+5S8qEHa/BUZhknJ1QEUA1F0GNYmnAopRBQUhS+CY8ImVzs1pddQXE+YaC8O
8uoQ4/TvKMJp1HVnM+45Yy2m04U1iJPN8mgBMyBJh4B6uGW9g9rnIhsuLkkcbF9Q
GoXygxF0scywflWA0RHE8l5UP45uJw01jqVinoyBLas+7z52Uqp1riZWoueyUrED
h9Q50QuhIB2Ry7K2+PoLfBO/ZXDV8u8sjTBLp4gh+Kv5yrQSuPOHrFS3fPnIu792
w+495ASOH3Qo6IBwLqGT09kV6FkcfED0YKpEknRamIXSG0L6t/QSOarlEAA686kw
QbDskz5GIxN8sDL8xJiDUSev995cw1ishw7eeqSMUGAmAprh05rs3DfOzAjhVXIS
fPvqTNoc4HW0g5aZaZ0IWsXlbDqVGK5CRxRtcJGGrslngQ4bLzktl6OQ/U71NAfZ
0n9GeLZljHwY+Bp8gpHIOB+YO7LsPpwQwEfqLLSdtnpO24ZKvrGY0qE1Nrva74gD
9y1gGHpdK3m0hNNjJoR2elrKtetv9gLt8roz1K/lXRSZZD83/RObX5d15ygMDFFi
b4wyYqb/JcG5NoNIaSVfvluskEoGhKXS4t6H2tCRV3J3nyfVVeQnZ/Z6lDh2fofH
r5t1OIp2X+rnAL6/1XMfSvnSZTvIPAHk9n8J8yZS64RBIEnuswxUVEwbKIy9fxVc
R5DjqLjShUXjGdiEI9c8tuOd2D8VkFUsm8TlxowIJTQ8dyBiPPjcNUly1SOybvpw
Txbu7tGbqXoadoZMAlcRJL8QeELLEjH5G5unCdFZVuXVsphzHZgvV4KdxV55uKqE
wOWPFH0JcIQwjnuLb4aUpoTpNZlJ7WdsVXjtSQEw5KwkooUv9+/tYCt5gr8KEoEr
CknaI93L+QcGUSbBJyQ4Xy91oH/MfZutFBikQe8+zdBcehSMe5oRGAu2ALmIdY83
2L1MsgRR3h/SfFgREyNQHI0ACf0kUgk5+K9xQfUG4iihRWIezJAcmf5ViSyVula4
1K4+7aRPTXhfzy64arJD098GtoEdGxx7DEKxETDi9mePiMLNGuoSEbyzzqfQqjig
nr682kq7xixngoHHnn0wzVwJc6vP5nJNHhQaDmVQVYe8IO7iKQr5WAVR/qbOnri5
hZCjJ6cuj0MCouyMpysckiO+XLHmoB4wSweQoht0ZOevx4dGOMYL+MnyPHAqVD+f
hLN3+bloI97TLNKr6cFOPoQ1bkEmmgLHhTY2dKwWHMkx3Tga7kXzerv7Ncl8PJm4
RPf1yH4A7uFoHSF6KQnHASnRVJtURfpR9xlyp4MEXyDupma+2p3MdYV1N3p34LsW
tlgYCdrG3oEJxzW7pphWoXC4/vM7M8tzbIVaFCYJk0xpRjN+NGIGNSGWiNh6o9WM
KWxYT+0IndoAt6xU2i4o0SR9bh0Vi6s78e2vLxWm7mFLne0LFXjxF0IiHMU3pJcn
SA9U++hxXpChghmz0UsU4NwO6JB+ATbQ5iqVhAmRecFP/hN/WaRfCm+NBWdkzn13
47h9TMzed2reRx1pG6tQMlAWV1mmrbV3XganM7dIE2XhJzM+VHkT8pZ8WjAOydfh
/3oqJBxPWK7+vdLxH2JRCDRmfnDXhtbbPeoFU14x9VF5MussGh3f5QWF7HsZzBpk
8qpny4vpJY8Hwj9OhF4QrHg9AkiiPek0qnLPqQc8Tmyy1c3t8JE8OJY6UbsNm41f
sL9mGLXBLb8wgKzbYuQLq7XAa94WK5pWemxFGqTyAjTfsleb8bu7dqL4zKUfn4Cu
EdprFGpGVQpKFwiTIKd6oY49sYiCQ+c8vmuvpPmwBzhFLNbvGc4uEJV5KHrcYhor
ntE6kC0QXsCjx+NvewGuyq6kHQH80tyJ7qaVQBWTuZjNTHpCyaw0oFTtPOYlhozj
IUVDJoYPuR7Vln+W3u4h+7agLecPGxsYA7TkRo/7PGWQn7Cu2x67dl0Z0IQMM2hy
3f528lRUZJvcXP1i00K///Pl+ndVAlJ1b62CJJ3AbC+TadBEXJTH6untAeVpIH1N
QQlhXIfSVtVO1YafjcHpOollud/1rMvwFTLQI/IUTqbzOZKipTLn7MG75D1UJtQ3
O0ZeJMQ2X5zdqnwo+1UgFtzJYvivViLP5vmw+gxP9n27kgNuLLJGRkAJdzdA7Low
18KjlVWrxbm78qvd8gscCi0lLQIXIse3pyURVxpyJt52svExeENiCOGkiqW7+LwJ
3cCj3Iw5lQYtX9JhKX3rTYxN3jRBYqx0IPM0hRjpCTPVRk/07nYV+7H0q92v51OD
e55VMaISiFezRidadYW9GD/8LsVi+2BYUVQMGD6RipgoKENHTpKV/PBj2GW++RUa
/jBAlMP+6sPncGq9TXiej28o05jrRxwi8GGGitUIKNOGW77IMksqwNLua0TLcA0M
arjQ8MgTNYC4OS7A6m56+2zmVlJ8FaWH0dzWIRlSJB7/ysJwUclQWCTy+9WEvHnZ
7tflDvozFjwpYJ3NdtbUj+ld+c3dGokCqnGC9wXGbGkXSYD2MkGSVNSJis6An89P
4gmG1NwOOQ/is8/USb/tTrG7/PzOo+PxL3xG4b0GzIVhq52yL4E/09A/fsV37ocw
uqu0efcVOzp8jeExxbUJp2lffq/ZUQQq/ZkOQLspzcNeYJZOPzhoGj6b51RLqiv7
HwUnPXtFQZ85BH1DyiESurdm+/QD8rwDTEzSE9b0FNaHgN8gfKki/fAgJZ83Zor7
7POVHRHC3MPNupNbhKrP90iFV/FtoB3ZXSjg55r+BCXtQdAkxuzC+nJWA3iW9LPX
lon4LAhOuRIRq0Q/c4qHoCJZh40F/Oip9ZyKt0rncvNZp5V4S6O4izpLfa2Sn60s
KHoKtlV3bQ9taecfO3t9m+xjCOn7hEoBC3Ac6gY+TMvAiL1fpTh634Tv7LQBiHV5
WrbmQCHHlwx6i7n84/wpstfanQflosCqXusd/LCi+7oGIcL45i4vU3G1hjKZ0uNR
tMdYnaWXjnjmTXAgw7jLOddAT0zfzh034C/ezGqrX+AH3Kcl6NTI2IVlloOdgU3R
vxPoGFVCpkPbOUR9RuD655Ljvx5lGEL/GBZb+KmhdCy16uNXy+h17smrGI4B0Gkz
Ed+q66BI0hOEbW8dE9uwHa1tT5ltu/zW4VmrrgLiwbEb0XPpvr22u3eAriO6I77l
ingrHsDt83iVqPJYqga9j0pTMYgyhAvank0upSHJUMI8B28zzoaJ8igeNX/eQGAV
g9j/aOIuqwUE7EmLmrg+1xMvkxi/d3mkoNlnybEMtF529MHSfZ5q2wXhdzPwPV1W
XlR7RyeqJ9aULEWuo2E8yAiDChV8nVNEPykA+1XK1+niuRhpFUGvcS9wf3z7IMDh
LC7b0Gw1b/X8/KF/pac4ku6dwdVFa4F1ZPOu4ZxVOEsYwl0z1QEvbDlVwxWSGrZj
jk9rEmSs4dlAK/dVNYg7x3xS9j/XIVJAdqpIIXn6eGPRJZ55hiNp8xXjJcvOwS/3
/5YSorBUGrqJ7/xVyHr9aZF0zLp5WaPYevZv79kyWzaR23cEBv40UVIx6l3dJ1T8
fW4SjNCJ5XYz3wCbtKMcbcF/MlaQ0KY02woO8gTw8D5zrWzBNzvexY/qha/7blvS
evqxaGQH9/vN4v/9oom2qmkkplVo6mNxrzBrfnI05JV5enddpAnwU0XisMwl42L8
99u/esoFvpmfNxbpHlMvvbEyeSZV2nrTAOCfsxWLPKEueDFC3OlOOj/YMUVeXkWr
lsJF5bIXrVBqFglkH5IbPWw8I6xd8gifR3hzWuu5DCtZ/lVbZaMhshLxa32flcpC
5z93+/YC2ANTh4pXU4dqd+EIuI2TwNL6ZKYG7ggqGeHfBu/K/VO6PQUROJd83VuU
JRA+8Bdd9IyiGq366ocykevR5jd2QlphI8VvB0tYi98xoSGl0rqYcKPxpVcfJyza
MZG7CaZqotRZAu6W7QwCv/xHY31FCuP1WzS/BFHXr3iXhOkBFrt1rdNRi6kPYLko
oy4+hZZLAu1BroaYOyC/uaQat5xBqJn/pCOwylHblnVzVYvWKkCYvf8s6JR4TzDA
jDYV4QVcUA/Pw4ZDYKsD/+THkYIv9TDXB56eM4RBR3KHtIFZLpnw6ns1R75gV2d7
FxA1muXJRAlvB+hdlPRQov8EiYMsV160jakfS3e5adi06h+Xnj/pJP8sbTNmB7ST
slM4nEIRcUYe90c+s4NFv3gTSLYKpCVYFwe+iyLdOsOav6MdB9RdEtwET+yX8y7d
Ux35b4bOLXWybVNPImV+ve3ZjFbp7/isxwoi83TzuN2CrCIWumHubIuO2bZTC0Y8
Z69yfUgbzcgEK5BMo85m8G14HdnUBrJUMw8HEdc0Kv1RfD3xHqMXlKA7jpyP8zc9
Ncn4lQRqw+ptQSpSSmXJu6eW/w35QXtFVy4sXGBrusAE82f9Kw+dt7RUJ870zIuZ
eUzHbylzXlFPIrMHX6y4ulTkxy0dGejxDSyuXjRSJmBpKNYzVAgnA0sbu+aqzjnb
U5zfAjJdp/U+C3MllPsxwPbW4GIyBUA2JmqZL+GE6XCaHIYYpGST/WZ0G+2dLU9k
e0Ukt35Cp38B4eZlf2+crX/LcrJPRP6zmzp1dEo+p+fSQd+xuByM1O4+/gwSqOo9
X5YeySITyr6n+IadI/X6AtOm10M0OPretXaF7HQw0cS+L9F4bClr37xyr8qKfeha
wIOhADwsZh8n0EjYlehLdx11Gpl/BP8wAyWdIfB3gKC4mnaHyVJM5b9S98HuxdLH
L87fWsOiLDSZsVo2FQ3+Pm+Z+uRYTpac9Id0TQnN9mPmiO+yehkBypYqUkG0nNHV
7QAfwj2y30wemQbEKaX3NRf991vCxU/fc+PsdgTmFfdZKu2uDERBJqA10M2LJOpY
Vz4TFTyhwqJfdfW46rgqvz8wIVxqOinX1AUMshgvVFPAa8giNowq2y4oUbmHqjfv
eTKZg9C9JbMCv9a0BgFS8hU4pDDaR/PPfugwEhZZWdxQkIavcAAGc16udbIvC349
oM5oRmbDzyxsq/ecpP2eQRT0y3Z89cXvNgz9zv3GL6kxYNFk5SYqih6Rls5OR7yB
MUvg9uEEQk1ySB4JiOpDmHfMOlwoq5t8PjVlwUnD6/rJRv3bTK0Ww8aG6r7j7LZT
CUA/UX6UtoZUvNM9w5FMLokRI/3d81HjgyDPw0/GKZcX4Nnrt+hXnJZ1FB+B2TpN
OurkOxDjApiR4+fa8oxmsSTF0I7i3rJ5zfiWCnH2InFYeA/pmeKhbPdQ9H0FbbBG
k5xwJMlWK0w2Rq5ZwOdXekomkBu2csfN3ZImVStArCBf/un6tMRePWXFnfBjNCRB
VBFArQ8mngxSqE4VB1zoaaGfuAPA07u/lAC0KXPZBD75RkAsPjmOyT37CSf64ZmG
5CWVYHJPTqqZlzHfP24n8Jv+VzE6j5YzPI8aosGuHhOC8Hg+BFsIcVBIuE1luHAI
wD3AMWCnesKR372pYkEeyx6BiW9XGSbLp/ZIFo6egmwjwIWxjN3lZHuVI4+oZu+K
cw1OY/UDo2bAwLQ9cyuoY+E7LS/8IVOlondLhoiiBu8Kp2ww/IOYn4EYQXdLmTH8
mbCUzgX/RPwz5j9SRHtCug0Jze0Hon6MK9VemLDPIUtAqBtU4Zd/brNRJSOoZCsk
I31YmqYaLvFDeeh0dxp5MLjNVRU3vuCJHueIeXmF1e9RPMb2qVPPf2/dTTgM9caL
PWso0gaoR3yqdanOhedC56rJEOPokTHL+Je6mP4vxq68+1SPPjiZBZKowEhaz4/J
IZlLzsQrQ2NkTpLommYdvryzACDGBtTWcZx5uJmF07iAgOePE8LWE54rBzIvBoL5
dMQHakFa5HkkWhjH5Gt+tHLzVX5UCaQqB12OCS2tKUp2FW7PIkEcmZToY0YQH1CC
C5MOCdaLPLWSf/W14FboloOIkr99hi4Ij7y4DXX+1bKk6sOsHIyc2oMPVQW1kUbr
HBPC5nqA7B6h/RVnLoY5j0a4fRi7+iLureDxX1xCX9ADnN4gsrN6pwOIUlXI1DGN
nDT+SNjCmne296xH2KHk3yKSQFusVeR3T+e5PvFv09YaWWzA13XFq1FJYsuzAgYg
IlldWKfcThWLpKAEDxK/taB6XUpnl4z8+R+sKqHjQjXjp09Zt7EqM7zCGuO13ngC
SZE/swVXdI6Ts73EEUjZHzk9/YBKeRyB2zdTWUjviEolEm4Y+syadOsSYsqzEK4A
Iq3Yw5P8csIpkMfa7KBkukFF0esABRASwst0KVBhiO1ad12hT6q932Cg5pZTqdhy
FACuMshKSnfYuKynUHWLzVayDTjlQu2uP2iqbsBvEUCwZJYYWjIkKsuDsitM+7mk
EEp2ibCZZkI16mJtUdTRrrJkqD49Mvs/M8+2DiW5GfJgk6TbcV0MJIanu1U2UElr
yP9kdLiH/W6Z+EhWB3oO1CP8UNE0iVelLNckZx4gvvqDvWlS0ytWDjfE0/baT6pM
nsoTF+QiljQcTkA9gUQv7hx//kmnZLdsBk5+LWroI48kMoyXeWnwjLWXRlsbSvCY
YTh+3A3SHjxt1vE9BxgxbdLhZm1ap8xiEw2zZszjLWQuwMM2/6dxAJoOwT7bVnFf
l4sDGpBmeyfYpPvKKzDJG5rGX9pujUiC6jDkMU6a7wnke7MY5dbQTwd6acpW2+le
diZrsUphV5e1gexFPlxcLwSoRRLDDjvtt7+rb+nPegSppGUSoRMq4qaerUpT2gC9
KUYF2u4827NOirK3eKDzctcuZhRuI3kehSDex4V9TEdSHUAtMKxYmyaCyB3AQLKh
d9X9h21OAqlkwCftFjAG7rbxWf/YXxGIxTVoPlXHiHAc5ktyh0XxXKqORRdfVAxU
9Pme6wsrOOOFgI2IhjhDkmUzfXzJ9SjAZoSQV+xXqcICiWdNK12ehs4+qQOlvjyj
HBNPSLB1tqj1bDZqTNYB2JHa2Jx/EVNb7tbWbrg4ytugSi5cny4Ohn/aW1ONTuoQ
kSkL6MgANjEjV0KQAkjeHuWou8+PCBaSFMbMZ1v24zwcmi2xW/KzPC5Pu2maa7mH
9662Tlsn1yYl8Hv6OmphOtssmlIQMuvZoO2GLk7sRYDAhM3fXWJwwm9yE9gPOH5k
NHTTe6IBaOvdZMsvQ8e6qu5K3VWBvJukB9HEmkyCj6K5UI1fPx+Ra+X5uZmo/g1h
EMq3+tM8QLl1QJvoPGKQiW5hoaoYUikF6OEoVbjqVWPrPpmbB5/lbD78sQ6zlIP/
7Xa/8sCxba5lIaQRR1a3Ca1vxsBI1J5Pt02XePu6M8itUVSems6M6QaH9bT1+kaS
mb5S9pNEC0YUn4DOkfodr57P2dNaSeJ6mke49pYESoXaaoGpChA/X9KGj2QLIGKr
93nPePJT9q/XcuI0I9xqC+KqkKDLoXHZo83KTUrA4iq0/QYt9EqW0R3L3LiMITa+
s26tHcf9GDxGYFO2dcb9wARYcEYDL0NSBj1O/G1xlfuun1RdcDQmBSIwWvGkDN8t
CuQppmgPs9vyhmoHmTdkP6vJov7ArezK/56odm2iEXjfLia0WgNF7XJeah/MRXQx
7jjOuyquXjBzUpg4H/TWmmH4v0dypAVnNeeaPQn4uDxDAgP+EhmCETSHvBLkAzsH
KT0vzSxuEmcyuIsf3evLlzevoPiOhCs0FKzyCY3WoyaudRsnKCgNPRp8o4KafYd5
fLiHeZx3Fya29PcpH3xHeCOtZeiYsXpOaNWVbYZv+Z+L9AT5zn6jYNu009AONwf7
OAmfCSKNIyqa0B98AHVGQ46BRSWb+xS1gBcXmWApFGPLaNeokoabSKAadpPPjkyM
FhOuJecRSdkA69lofBhoJwvdpiDkoERkgJuDTYuGILnun9ljQRNSM7AAczvQJGjA
rJa59nhGet3ITgDO2XV9fStLvN1J2AqLZG45lknI+q0i872UeUv9Pitldpo/mYjT
QIFHns2kJnXwm1u+A3Qq4/gc01RWe5fwdgXPlxlXOLAIaPnLA0/yfj53YNjHB2kp
xnbUtGYNVfslc+vZomQu/SqF24BTM1YXTmNjE0ztjA8HbqgQB/+75IeJHpiNNdo3
VpbDBEHsiObxbBIl4baklANFC/mR6A9LndMTz7/SruRmhVnBMS6ICx5+trdjri+t
d6Myc+42juwH+NOfuDz8KbZRywt6TmN4Tib/PPSdanKIcx0fu1ItaCQhr4vw19ar
sveJVUfL54Ats7KUn6au+g5iMch8vuBOqgn/jb2Ste6axNSq5sFq2uOxmakMlFBR
efGk5mmoE04D1yndHpkhAiFE6BON/rjKz5zPwAbab67gsZRVYc2y28zc9in2YeB7
q2NkPH/Io2yYqP6Ed6QFXWh8MrA/vdVCjvMd2TTsMRQZ0S7Q4r+1ToT6F5z1oCHL
XFgvMXxgLfaxPbgRUOzmdoX61x26Qirn7OO872c0XMMLBEPEv1LNVF7UGS7hF34+
D8yJmjX61Q29O88FdlNsBOsN7aD8ESYXAZQb8dzb4B7SKPxtlQvPEDCF3GMGGto1
sQFsW2IgvzHNjBDI9m8ZnGEr6M57URfgdC6ghSyF6MXeV6bOW5mVZ03ovjhdJdzH
BcOboKm9JI3ivCKJ9wnQCVx5oBIslzmLN4ReCgSPeXUPRAgWLIHnS0G2a+TYrNNl
zL2WMzaTqQZfgmaOq3MnT6i7pWbmjlkRdVz0FjGAgrQJt3byjBS3sJNb16V2aubG
Bf3pLahOEV/WRnHBETY3sxZ3NVbN52yNeupY4hR/O2S2X2kyLnxiOyO6zUaMQERk
R97l4BimVKeTNcUsqrZjdDgoFy45KPOY0VehexTl1vuVfjkEWFtnNP2efgPv4MW3
iloeAKTzeWy0SJzfb+pnZnjIdKW2YGHTtugi+MlET1HO4HOmBsyZs2EB/fTrPXEZ
ofxlGldBXxYJyI3b4r1Ea2dpnr7E90LtIm2z8iiT1VL9nfzCGPrOavUDb4ygVuGp
bNFRY46h7S975g4H2heH1VufwpClE8Q6qH6+6u4R7NHe9PXtmpf/z9Wjozmb7sEx
d2Xd4aFCJfFyM1YIm9mf9pnjeVKK85YbN/UQX4juT5AIoid7NEmExWwGR6X61CsX
cYVgPnnOa1tPm/EKqqHfzZtMI1N+Qz/xGmSKu3zhKvscLlWCeiYf7+bNQf5LxTHL
7RWrN0BDjQjnTBgbkNBVoZLG1pxvHTABBVCB3F+iOc3OqQoABFEvilWONFNDDIP3
MQonEfd97TI5rhi754M7a20qezuXixuAP99opQALhi/UJOe1nCw5GfQukuXDbg7m
YCs+3ykrJ5G+GGtCngsUMmhOK4zd6isobhpRjaNI0Jtl6bu+kfikDb+3Z184ZbaE
UaaNJL0X8KGTK28Zf+fnVYk+cLQFc8sCVOQbhnkt6agpXRLajodVvYd2bEbKdlU7
jFrCAb8QCkChDR3RNcuME0/4X3g6sbGQqibZ6neZ/7RO+2xvsBAJhA7WAajefw4p
QCimoDQWSZ3CHuatmLOrdhFbfenJ94RvEQsqvlBza1JWh+brh+gcbVu3kfOCxh6t
yWXuqVboNjYX0vPkIRVZvtkziNgz555mNl4SS8mKNl9rNsLEte8Ua553Tzx0wbtd
yrO6Mjvv8g2SdKPeIKtM9wr3SI0SN2JsrOar8lKHBeouumRV/HiO/2eZGigwyoKr
wKUvmHa9ldIkXHgZeaksbHsrYZajLtEXF0tL3DijOY7cpt+f3avpsS9ruYlSzXM7
d2rdBGhRrKj5wIPNBfHEOHc1te2/mcGPLk1zWrcSOS99FHt+VCbzaqFnIk5JmFX3
+jtnh44Dhy7/p/50rWoDcUflv3NXf2oMxD3npSZ+E4uL+cF3by5ihYKQeemMAAI+
1ijAVHuXhW8lFzHOA7OCmWfP4k3NBJWkFm1NGLssbDm0ge97oSmG7Bl/Jucqf2iJ
WBOQ+PJsooVxy7ZAR+t88eLYRtYPu3Yt7cupdCoWLWUo54ycQBm5UO/vtSCNtgC3
G6OIg1FRXLbupeOjJctAMaJ3BS853wNiRIn+Bn/qq51LnPd3UhI+U3ZCz71FF8wT
FngFPCKjecv/Vouh/Z5jK/29lE8HPL6we7Lko7+eu8b9J1OsB6JoeUwidHSTRf0p
lcHbgdp5YVi+PnZfY8IFa3DlkwVEIj0B76Bmwy3zcx2ozRqJ/YgjBpid9HS5VP58
kQK3MNQdxe0ICipQ753qihW9CwaLCulyYdf5V25zMozBSSKv9Hb8naNqB1bIfb9m
du/4+Ji2utkqFcW3xAzDKc0baBpMhT9Su0FWk8/csc8kzymst1rEpI0Mx+RE+oBb
bwxCLK9POtLorJZwV9T0eUHFvGaHCWp16aCwtETvvRToY9J9Vrepr9UDCRVu49m2
sxIJGiZkiQgvB6Deym33jKhKd8JSXA4nk6pVeVWw1/rWC2s/AZcEqzqEsqGj8RYE
EMdWLMA9jDpyEop8OYfK9xyHvBw+TnWOn8Bhaskf5I5vjmDwiDGb8coYqk1Vj63p
JCYpJ5gP/FTaew0RtUcEwOa0DgJINIDMtRQ6GGGns91fz7l3SdvXqTeD6oelMav0
+GgjbB7J9kMcozsp37pYqpE9ZqXYpKEH1nwSPck0W08jzoDqf1so8gI41im4E9U1
vivHjzbxuFvmdDJEfDZ0ZuNNLj+kHosYXHS4uAcpx33mS1mzFiHzOpxnlgSMPitb
cp58IgnhaK3d/W8dQcCf6Hb8vOphazw3Nh+DU6Is+r88Mir3Fqn8sDtq0SMQBzEJ
G6xkbq1S/79Ljr8h+chb2xhBBCGV3sZN+VI/OVBUUXX0fxXEG9w7Rioq+veM33NL
t9H/ghJuMoi326y5s7TKcbC0AHwCKaPY4rmAco/lXFrIjJ4jAKxGJFPk22GSwCKf
zVdyDcSqqxVnY1dOoCueyn4UMEz8bn2jPbvDz05ietib1YhciJ450BkGQcN6Ku9N
mkCgEh4eHwgnVYiB5bKNeN9uqcKb7FYLEQFcSucgwtTIQ6vwg5XTvG3jH7Alhs7D
Egy0IBXakFpL/ZoOWln0Zm3y2m/eNVuNcLD+XL+UaGtiaJV1VMalH4cLMUe5PaTS
DJWJsBbLLpVVU/3/hlI9MjT5LAOa8ywUfn3FwaKyinNz2OF8RFjTnWa7XMON5duc
mlohRMXH81kxLufou0ZX5bd0lLUB04Phe85kVuXHIxi0oXFvFGm/UgNy68L8WJw4
x4gXkhSYIHXhNR2qpQhiONX/ycGWNOK83dYOA3ervDtJhHlAZiT+aa/f0IpQcCoh
tg2Ru5HT1wLVnhULKUlno3F9Uf8mitMhR23am9lBnvRepTxD3YjtWahtbd2iwa+k
rn4CAzOP7ZH8KFu9QUdEgyysIqpv1Jux0KKZUNy+8OZv83G3tcNXq+9CeSoJlCTY
MB+3N7CFrdBpbU/VquLV2kA3SQA4wu2UU1o60Vm97QHWRZqrov8ZAsAz8afgDsNB
yO80qvT5sL7G++jUABdVh/2O8eCjU8qDfqht1OcLYlx5meyYZryimEClXLsOWO8K
RYraZe0xt3Imk7AwEHd17+Qqx82MfQ4SJFdAzsCYoCVKPTLFz/0MlM0cIe5UhFQ1
j5rs5pMHY18iUAqpvt/zkbm6lv/cUvHbx+HThyHIcPM9SJqGpUguUMhbNQn9qe4I
zmKBQ9d0Yts6OwpJWTGcTqua0R7MnnT+UnVx/L+FJT9PV+YkVu64/2XHkHKo9NKM
wpVZbYv3hS/pHPfmm9SZympCKCuZH/ntHAi9yhiPcSDxBDZZ+NgFpEKT1RDtuM43
BsENTTfl2p1DMXXFoH/KU5fL9JyUR06b7aCMeuGo81OHgUtXbxmd6dLa/NP4uy7R
dkXCtk2NmGuN0HKJjhIZMsZKhJ5kSi0UcrKLeC/hyYETHMUjJAFjRvySGKrjeQGr
lJTakvwK+ycjpGwsvYeRSS1QQ5bzIG7uzL9oCtV/NeW8QINT3fvfihXtB+rnLC+q
Nd3FL8ewsVapbEHBvo4dsmypn5Zhut9azUQI7pIK/dGvgho/+h3H4VUbfN3vQavt
/wcASHF3Rai7B9RvrnsNWuNyhd5nfFq9zGoTzxLkDKWnZpZ73XE0qHPIYJlmABdT
5HHJf8ldG0Gn6g2uD+ng5yNwJdpG1bz3bjI8WzasIzFYYTAGqlzXRDvMv8fhnLUS
EOOkXDgFExWvzenAVlrjlEEvhrc6a1PYE4qwxZSC6uXr1HdNungGK/16jPoKnUf+
955k9JRdHc3MLME4MSouLk63+EWKWmKA+g375zym6uWGKFNP3Ssw8NR98Rm5g4GL
qWo7fmBgHKxU7Rn4Zsu6g6WPt81TM/yWb4JmuFqFgG4iUd8N+uTLTCVVM6vDdCbr
3SGiQs+0gIJPI22ik92Lrto8SYK9cRXKILw6G2Yaru8kT5w4vNU2F5E//gKr7iRh
cIUMO4LrTokRLSgINCU8lMG4shsKUwvwmWuwlZHNPjSuubfdCOChuebgELHVEZgf
iWxnU/pl+pWVIkP4qZeHYLRnf03g2yvHMBNm2DtRUzfgzseSF4JMhTDu1np9kYCE
UGP38fieZ2kT1/WVreAA3momE2hms/jotzXociKKpXlFkppAoMltK5IdwoCJ9ZMf
lB3zDoMJWHkQR7PfdeqqV8JW7bsy9SX3XXTeftCm2wkNp2wTfenRTJlY/iUYcSOk
8xwB+aX539vjSqnDqaq/iRfAI+0wBOYuBoOnKBy7URAfxsgw0qMAp0g/jKO/aVWe
sCrBhtSyIpSs8np02rcCzwBYoPU7gzleaE1e13gHvHOP9Yv/uj5QWx1csdyCsn7z
2xQ8n1LVaxbGfQo2ePE8QitlPsL7M/1nabHal1KGU43KY82bHe/xISgMY1N1PpYL
XCHczTJJPg5gGg2S09XEId3Apw0coXXrCGPqZIiNT3D1tK9O1SPjkhj+6iVnsNsS
UuH1k23LVsnfEM84WguGAWILChGZ6OaQGSbsV3xCswUoi6SshXbKqbsCm1cY0xKK
DoGN3VFOiQrWuCaEfaASvukN/f09h9T+mdt+heEN8zfFMiegvdP1eMibj0v/hk6W
O4KJlutz/tQeCcZuaVwwDH083s2feBYmuhv79iIXz5nH35QhrHoJuF/HvwyuKTks
lGPSdm611EsxizsqjbrD4MvRH1CMAOtMYXphDGRveXJcq6HH39y4gnd1g1cGB1cZ
A92s+Bq9IyE00d0g1sCplriCER2YCJ4UJPVGPsjYgCQ7aT9oR8VGrIoXwSMs2cFP
sE+XqQNdj2dLM/4nH4npz+bckxkWzLAF7imxmLF1NoY4GwySL0mkX04yGRR1CyU3
3c6p6blA6RuQnsghNUfiiqurkc1aDQokzKAxChsSbjevBbNMdPwkTNwSUJL6Yma0
TVeL7Ym7MhD9QfUcLD47oTMDcTJ/4kR4nUXHs5lPIlvNCux45P1KKc38UQSE9Ho/
7X0mrxVgr/dGUsHFk6XL6sPRpsNAMEuAGmhT3ofN80XEBWyecNaY1JpaVi2/J7Ko
RyhQwdlLJ7Pjuqw6v9Bo0YWdt5cMcbgLCBe52Ukj+2vS89GwJuEp9wLChGQ5O4EV
48OlwakR2gSPNPXl1rMkXtMHDt/wjZohunptTdtnCmhmGzuGQU6hGnHkY03EF2tX
goyAeWPor/5cLHYGQ3PqWsUVwXShv5Wqyv4Wlhzn1yRiIeuD4NfQXeh2acCucgC/
TxUEScJpcqVggb8glQgswtqN+SJ5qFB0cf9Gg4xe/jEVt77usj+/ccf8eIg8+J52
Nc5vAQwUlKItXGVcDkv77iIQJusvoaCqt73ndzqZfLA/xQTX+a7f1ELiPspjG8Jb
V4M2Tk6ymJ377RfCx+7Pap9O9jGkyAmx1F4nXqz5jvcbQaC1YuXniJYJimBOpiOR
bMe5JFQsCyt+kZlDOuipnrCYeuP6iXtQeDn01T2oW/bOTS/pEpgHQMz9a7166D4H
Ph6GfDj5fisaNy5cp5UHAC61uiNHAGwVHhGRhpURxokdzDah/f1X/0/Dg8wja7tl
yh9R7HRooqGXm/MAhu8nrSa93VzkFcVlXzdUsYS41IamaLq6PJVwZO/ueg8yu+VC
krpzLa6Z1lB+mSxHUVuz+6730wQWJI8B1PRrfxNgXDiILtkts6HNbuPnjWtODY0L
VVt9BYJw5uDU1vcf/ssLeVssVA6FkFH1PcMrXl/7/N0HClFWBlA50ZRxdz+Bfb70
U/qH4pXN1nYeSkwTkjf22sYBP9LutGU29O1t41YmZdrz6WEmhHoRYrfGAvIWQ1lM
jYf9BcXtEluZ+6RJme857xZR4LNAPESnOVWsaSHiFcgbeY6E9yW0ThI8tukAPqNF
ngJ7CXyuUAxtil22s57eepA0Km6b4+bNntbZxEZ7vjxRZBbNjMXe6VEsrwWKHaDd
3NAD3C3HDS1zDio8pwNeCp/sS4sjuiAjPuvIA7ZIwMzD7BFR/l1ivZrwvbFcIVwm
MhrEWjB1MlSJ5Zem8M9TTQPl+lT11IREcQggiTfJsudxNE0uN6mu8Yl0MF00vdOg
zTXN31wazgAaUHbjzFfTKM260+wdgE3RypZkpTbWL9gCcUBvvFf4I85s85lfJ74c
X2rOcR8X0tYZxfUjYgkDsOWfbh06PCTbojm1Z1dPtahewQS3WQNP9sJhevmWTPEQ
Y4zlwuMrFHsNyp5zi2P7TaJQCq4SRSJKNPK65qpamBNQRvtuU4vx+qLm1MFu9mxs
wJQCdAlY23LRnEm/4Odd4vY7SfI6MrhIPiHs9uFyk2K9BcCp/WCkV7mXsxGFYnbv
Vp9jTbpNnvWo/2mD//lFPD+ecIXFHV8LTStS5I9YR/xL+khNQOGBhgs7qzg6f6Aa
DZBbifVzi9iCA8FZtuvmYS30h1eEiTh8/CgvMrjddd0DeHVUN287M6FpcIaaRASB
0xYtzu0cvQ2Un7HEPazxPkVJr63QxxaCCwVllkuoy3Us+bpgIHGlelAUU6lT0UkW
sRCEJ8k0uDYT7SEhgiZT9VdR0RGil8dh0Hc3Dxu1qx3cDGNeeue8g2zcbvGKO6/O
G1jWzY8VpIF4rvPh8OLzBZsZDQCd7G8CaZQpLDVl2LlKovTXidAj+eM3EaxdQgAj
gt713OvJeOLSq+Xt8gW2FnHMbnoisGy9+1pmhprxNx8FLzrDsNSTwicX7a50sYZW
EF8/KxNS/Yhjg1bg5kSoLZeNCZD8GcFL2c1daCDm5cvtkF0EjzyiQyAmlkRPWmXq
9jeF6C6Fqdlf8yznzLlu898JS/2GYDB3mBNicwZM/hezNP9BAti6JR7XOrLlX1hQ
2Xdlx20h6AWE0I3ebzlRVcWWNI8R69LrzaoidP35Zy36fiPaUVsqVNTSXSyfxRJu
jtfw4EYIwOBB+zubSpwFBCrkBZGYboXJjyajmKIq16Tp+H75wrC08BQbFGDwwEYX
GqydM2aZsEmW8ztsg1diLulhRkKa6Dy0niefwc4+f6+fAT4u/6xwltqXHHOAAI7P
E5l5ZQfIiYjuE0gI9ucX6cnhfxYlD0oZ+odFI4DhuBLaPP9YvCdQabYfpkdkcAU8
pW7o6xiLYgO6w7Qo7v3WF7RX7EqFMzTtYgavhrKKVBKR+wZcacrzZRD5W/iP5TAS
FJygfAyVezSH1chY04gwEoZBSZmYxNlAoKt4rx2I+9jyy5enWNXEwacB30m+Is3H
j0GXYPNOEqW08SRb1OCJWzdjW8HWKoLEoUkFExxwqIjvhZ3Q8dpuNkdi2LMU3Ozw
d84uAVTThjLnixYuEAtHNMHZ9byFD9L0/00pqa3ulUFP/5LSjhcBQSowOcLtXOmV
wlnbj8k4T19TxMuIQNWYbgD5cKqVBDeBhUDJMzfH7ZlwMJV2ezFKvJDCX7AFRRIH
8hu+LH9fJrBf5AVUlL1emNR1sQs6EY6Q5GNZggcGitdNcGmGQZ8dLlHpj8jsa6L8
MZLCL3TTNFkxwDmZQSYn8Ewra8j031daKfIwD9N5Rx8x5yPbPmqq23vIQfKnKvRo
sB8wDMnc8LbVCWpyv4ZcTKEdbuM0/qsd1Rk0RXZLo6EXgwDtC7NtRX9kKO+PW+Tn
4aPLOqIaTu84Kfrr2tukUFLaplg30QA8jW1iuskrQRcWIJ5er6cCS/YR8p3n/RVb
rmBUzHSKIPPNlz5MREyzbUA3IRwPI1RuoQVkNWRi/K2RQBbskJP65mMBKaufbtqo
LHERXSaEpMgh6V0yiJYqGGBUBnrkc3LwxXCE3xnuHSEenuImrQKRAkDK0KexzSiL
o512M9/BYWaLjKuYw6o4VzNlE85CDjNlUI0V6ec9G0N8SjgtnMvfvhPtAwVRxI4b
4LvVa54dQSVuC2xA1qaSPVFITGHqAeU9zaL7a9YaIXL8LDp6Q3hIPHwEDsAmPOCv
Fj6Bw9zP2H1SSn7lmNiz7FoKQeGRtuU8BIpsq9bnEN9CKnaLCKCY06vYKDMkBpzM
h+1sWjIvo4IBmM2/0Cq0gwgvlTh5zKVo3fvuuHdeWzqofFVynoRdwj8njXVUZ7mQ
arJdum53JxrzDSAUNOJBbB4JdUf+PAvjuonoxY2TSgQ5NXCX+IvTiEyJo2yhxoVw
8+zrsPbP5O/1wwlwTt7RO3RX/ntgtbj4K+xdPBe3RC8RjXbkr6HpOsDwFQYH/VRw
5vVQkDIs5XB0CTVzhG9tmGiu5O6CIVgwEVfQ6/aGjl8x1dUF/Tt2jfzxwltknQ/c
LkBI/ctRA97LrZ0Mh+4MHbua6iAQSRmDqyPpoUrYpbPXnw9vmPHNLXy2FpRCNGwT
tJdDt3bZ/HQaIzijhZ57HRmS6AIcITE+QVSyv0vQy3rsZcesS+zl9Bu/ccP2tUnj
f3CyTHLyeRlTvVd+Rl/+b9Y0K6u6eCWLQNFMgG7mS/Myu0Vh9dstEqMgLjQA3cxx
70d4qOEfkbjKCB13uYSJEURSs/2bhkIyJUUw2IB10AyVhGxrW8YOPGUFgWx77lRA
k0MQKxoyts7QPrJC7sBoJ9FlJzkdCe8G7kH6Gfy1yccdFNgSF0HHECqqTM6VN7++
abS22ZgK4NIFm+icJLMIZgUowx1LGtQ4dsMpkGxKeDZ3pzLXTD5Nqa1dtRojOBpl
71XaN/58lItGYxb2FLOXLzOAllSvukiqmSpOkfxL3oiW6PW6+9aRWqS0U8eMA85P
skLH97qT4xOQg0b2V7sAeJZqw4Z17AMve22KdyJPAf9/35M3UmfdiiXugxVmDGWu
9WseBwlgQYcNje4Q6kpl4EUkW/xuapUU0/G6R6i4B8co8GrnFxp4iJBBpwR1m7FY
mFiJPMTbjnQf2Tur1faJSQmPPqXQ8SnUIUAhkXa5EsbQQJjthtAj4l76HCxvp31W
ammV+hsclVTVsemIkEAuQ6e4/RNC66p8WQiIm8783gsteKCbAml7zltgCSrtiOwR
yVaId6QLWF66TRHaoinbs8MiLMU1SAivftv6QOioCV9M/ZZcu+d+C+kl7TgkqZiB
p48tDYIqXrkp+JImLPjVtQ6Y9fdEuYRtUfjt4OXT7JYWZnCZUAJnULw+Oi6F2eg5
EaU6eK5JsFTgJsfnk+0ekkRCa3bU92J1bCBPDRWzyWIS/LItw5tEHEq/o3zfK/4L
A11qwgkJer25WY7mKo0AQh7aToS0PgJWWmF7+oxeONsrKgcGhNbYIAucFojbdyJe
WvMau/hzhPS4YgNMTT8qvRfnDHfUHZXlXFzqXyTYtTMiAIH5DjTGt08r5r4KmN01
U8kzkwP7EaZDubpiUAIhvDk5SZi/LSIILHQhcmcanMDb4DC210bsngYaYGgQ/V8O
QwqYCGEAWS+sdmEAXICGl4yGklXmrB+WPJjFoJ4MwvnrmUVclx7Waf1BYmk9nyV3
XXn6iaTZNwIjF6sZ+6pUoGZBXxr55EyzB/IUyn34IfFvz8nTZtbPT4vyCIEZX4jC
KW6Q7ND6kL7us+oY31CFCf8rdlvAbB6XxzLaWjMApHCxC7v/zANA/PnN4ihohZtH
z0bFWplYutpYDV238MtENSD/tj4X/GdYtQEEoKYxlI9bIFGZMDOsYWkCKkM8nr1/
3cHqksbc2+0pFOVC6SDKuDieHXRy28PGFDcbAlc8zjX3EXjL34rCsbT0j3qs6dZ1
PbS6SNMyJ0I/K18p5wqbodMOb10Gn02+IvNM5JMqdNxZrilSEfZ+v1jarnnMweZb
03SvWCm3RIR+3lSlZpu1W5gn9rQrUYr0CpAs7DtDV0jRCnbJzRptthDI8eZ3rXbF
Sqk8YOVAZGEnUbEdqn1LrOHqbgj6FEKlPha29HVwA8sGxaGcGsxnJ4ONfWV30WVa
R8GJ1VMQckCKQI1Fi1Ma32F9W3qXX3Abpn4Os5s2xC6hRGU0kyyKbgSUWQxUJ1VZ
JVNo9zghiZuONhiVEpLn5YrOvmWfVnjmmqtrgLdF9qQn9xPMsYtRobDTG0xQ3sHP
axp5troKQlnfVkVS0aru1lpixbmheqpN22Ciwt724BhJUEUDQeeketP96aMVjVzy
etdCPXM5WgCqpZCfw0nAopLhHukzanIz9MdC4UFT5O52g56iFimo3D3CVQi1KQ82
mG1viCPmLHG1H+ZBGzh2Ywnk9ZhHvzG/DzyR0/IQ3t2aXIlZgFHFP1lJ+PLm2q4P
chV/lC8D1k2OuB+Ploe7TkQ6Ma+9B0vrqpzW5IzCVliXSpAredzNgRmAuh3ddLX/
LtPq5fYWz0AB9sWUcRYn3apOdmcGauYTMXw3mA1Mm7uc64MY+FmiIs6aGdjjxk6/
GfWCyayz3FBuEAS9vnhA/wgx5IV5wcHPyGMH/CZTkKsYtITOg5N6eXN8yEVA5V85
UsSXsT+U8DC1Pl4aA3vX6kCY3CfUwx1rVz2aPbAUUpCxP4GEivJ5G847nAi39i3h
DwEXpmvP7ksUtHEIdj0qDpuiI+aW9aOPVUh4QsoSkQRBj/sRQt/BXY6xMkmY7USf
tk8A5CS7fj5d/5R2CtuNaqxy8wjl5im6e+su7U+EBTESrvq02/rrtZ9/cu0Yy8ex
51vlMD1NZnHwTL9Nt26KpnPhQRanus0LiIaf+VYIOiq6tty3n1wH59Fg91dl3xNJ
rV7FOs4ybjaFBitsGYwbK1YU3k6AYaPPue/5N2wacXHbl1LS/trs7ziCb+Z/9aSE
LN04hC1eZe45Z0nS6ofhMEAKLJhoUkRDIUjTA+JviE1h9AT3xgtDLYN52VjRrJY5
kvzUk+xPeTb62HKx9dwR1VBmRLDoMRAeUd/SuMsoOwbvgoVl3Gdppo+XlizUhn4C
5lA2iFTFT+nygxx+RYK8KwCmiCxr6zoQefEwZjz4vuDXABWC+7fPYMYDaA7NzIA8
xR8AudSZ7U+hvSYWg+8V/qknJFNhaWLzWJ6fYwcqyIBEXmtNQkZMMvYWqBKufKFr
DqOGDCDHsNdJggcz1t42YdvFBqCgo20zh+oerQ7EgzEItTRX3Nc84MHRWVA63/TD
crGHZ3qwZW8c4HobcZPgBpUHV8rGb/Jy98xCbhlg1sRJuiFyDgNztvMmAIioL65W
mINiSGrLzHU2RB68pLjv1bp8RaBD9iDuO4Hik3NGUYhY7BJEH5CNXkXOje3dqf9k
dArznYg9J7QwouczvIyiF+E6P8T+4+qCe6drI27oWUhKtVLT2eR4QRoYdV7KZ38l
NmuRpwjodQxnx6Dgbehpg6mA9mcqDsiVXpRKLgE35yj2XW1IZ3IRWqfOiZh1MwDw
WAUGEOBlPdGKRxR44VtTlcriO9si5zIR8y1f1vTCk5UKkzbXiJHYjTO7J3lOl75+
Su8OnzZ3ppNSpVxfbrkv/dMbR+DE/xT4wQ42kVHiORRF6KErS66OCFJzOkRC9UDE
IcVscwB3kvRv2+P6nvOF3v759HXukN/cRjlFLXEQ/J9i2t/KbJS/7jHlrqB24ZLw
Zz9rXGumGLq44XInYGw6DuOUFqZAhGaAhLw/anYc8GEQrSq4GxVcH/b/T5T1Im9e
8QHh1XPR5qvSuru7AwDMyzn0le8intxYqUFBhUqc3Fz885mFGVXTa4RTCWMb6uma
NHIhWxLHmhl9uK4PJticHqRDhG7leh1Z3umPBe8A8exuJdzDWu1v0W8uQOGMoiFg
KgjqNIKlRFFRtbUNNRuCCMB7Eh49Fmx/ocoNkdDGbnWHdzJy4JHst+Jcbdr9e1UQ
cQP8lLCI0NTo49/uHQq1JI99eiL/eZDHHl2hbzqm3eBS1TAe/4ry/pO9HPuw/86d
G7FeZ4v1wgtYff/TzTFefQx5006hKfgJVXy7QH26gHMi2kvKZ6+tWibLEoedq1f/
7yUL8mSUYAnpH2okQyO21ybCw9vUogQLUD+gVzgxXVNeeMn+2UNmVguaOK96+t0O
o5vIsC3o7CyTgjtFjNI0SKhFOx/qtV5oPXzFbmLXtfKnCJSsYmVF+G1dY3ZEddWA
9kSI0VQ9OZcyNjNHn96QNPs337emZvPPa82midfurMsuk6OWIHgMfsW1lOx8T/bv
tmaXgJS9FNPrXgIw0J2zjF3vQGZtd2SsjhHYGwOaaqowaRTZForcwFa9I8tMp3Ro
yENXdZR5jiAfbLyLInq23TEKt/MnT3L5LUV45ofUQsorNcxTsN7MVsWpg5TzLwMs
7xMUzcTJxC0+ykWWfbAMqwF7C02lX16QlYFZuWGx9XPhO1Y7PScU54jdz2TctM47
s5o4HfkDFHLh5HLdRN9ufAosbw7fH6IU5DZ+ccxQ47vfFX9SHi1Q75p6DxS0WiM6
xnlYMJx5qLxXdd2C7LUDk/4xvg1jvuQyyH1Cyfg6WpqjGX/qFXmLaKyiwWGiDLCl
QwC09D7PTsWRaB0kKgo+JUiHu1ynh3DXAZJWd0TScrSzlJlGGIB5FNYVkFlSNFSG
zmk8fMgpbpliRm/6bc84W9YMYxesXsxDJvoS7RCMBVUyCNH3c91TSK1Yflpfhp9a
owHWj9P1owsVCXk9FGFIZ6HrXjLgoKg5SUqM9TI7a8ciHU687nl4eSgFMIjUfysu
fTWxB5UrsUcUVQPFVsp72YtDEOOcN/06Wt7ghDRG/EwowL8O1kzE1uBPwysOoO0L
+JrBaIgn8h5kgyk/9b0W6848CnITiJ6HBNnpzfBJM2eiRhXGyN97zFlSCyfcy6u0
fiQHb/XKQhkCq8qBM0tvKZCddwonK3FYMyuPkkW/XmAaPn+IyfoeyuYTVlnC6wOE
zR1M/JWbyNM/hTQnJR9PBu+98RYIRC0IOLifpMBhxc9wG3F3KL7lFKXdGFsSfGEp
/AjisWmZ68oRQxWx9dP7hflQXCpjc6XQIIoTGv/Jslf5KmWYK53UooHx7oSncuYg
TeDZSwI+3zr2//DesigwOstN2sE01tlKPJzaE+VFs3oH3f+M/SnW3/wZSCh1QEnb
+A75okrrsLWIZ1RBJdFq5zPv7JfJmEGuCvrUpXBMgcm+I/5xg+mJALdH3Vw5WNXC
Fg2t1lFKTG7PufHZDikN3bQCk/H5y+V9AWfP1J3SNXOjZ8ctMB+eh8n8AWUWvDHG
EmokSMVxfmfmtvL4MICGAokCzauxnSY3JNfCYsOqcaF8tcJAt16wfznP8EigSr2H
BVNmdnQETz8y4W479FgbZrWHcPRA1nAKFCgy050UqqQ3JEsY96SpbWF7vfh4Krcg
iWZWfVvB5LM99LrFeM2b2/vJvZPtAc8j9P2XRks03P6DKIOw0hGD/wVSM3te6j1N
5MgyBcixum5rtmFFhxND6p7zLUR5OtUsamWHt1G1D63bzVO4NL58iIh9p6d1Xmy3
qeeYailEo8GpaJKnWq02lrdTxgck635SjLTDZ2rApSKb2ymLVbBsbU+azH/fbSWW
h8475ye84zinAfdp/fXcMLmHe7JOVGuYV/xbf8iX1E1p5AngIIy10csk9GxfTipZ
W1hQiSmw4fZeSM+OgocgwjhnCylMYY5tC8H4mDpmfwIDhiDed13dBrs9quYqI+vq
i2Xjx3vhTaUtWYZNRhl1RzO/E5SFbTozHXIdnt8th46ygC8qJuBxnh6cK4xvqqKq
ehrLDsVOE5qinSYF10ps/VvDlIYr8qF+xWgwNFE8N/rGh5lVHYIbyLvTsZcGo7Zo
phn1vdQTZJfIF9CNSKosXLLI5WYUQHa36T2yPiBPA+KVgIYAFaYyKYI5xMM38Jv+
njaeMdxPnSQYIAfdOj5t4tQvbzfqFzkiVjKvdVzKgCATk/u3dN1LjpECX3MsTT0q
Z1Q6m6+dxPXPJiawwTSHZX0vc+kFo7sBu0NjKeiE5cwv2MilUv+Kh/deufTarS7Z
DmhcKoy6cXLd06uI4RXDust6igSgfLUgkkx2YcyETmYIJo+GUrGLBgBA8Z/E7WfH
jRl7xLXF2qHCC9Yloi9wM8yIyx0ItFl9HW57jsZXD0jdJRdSURE3gW9FJOVCnVnK
FWgp2OLiQvL/bVpepcV0x0nCi9EOec8JwLh2zHBo+oreWY3DvYNleJiHzVbOKw6J
FGmdpX/l/UuTbsIbZnw9ejHSQgJjG6U0UTmUuNXAr0MtQbhvx/Nz+nvP+If9tu/L
w0jLYyrFv3bsgmyrSybnBxsXA9EN+EJ1cKN0KZY4m/ac0t5K6xWhFZQHoHo16Ylp
ICKcbpGEoU/4HbAQlEjt6e7w/NHpOH3WomP9BWfAkkayz2cEObLxt7jsKjfJgCOi
FUwAcpa3w1np/Q+SKu3mJh8A1tCg34lk6UL2fqBb2GiUMTU0w10tgr9b1UXNWKxe
TqX9/50qtucNJPUgck0Ah1TX2XKry+Z2N6FWKPyct9YHGaIbGJF7wUr5iM4aOMSU
KWb7GTex0cU7f97P6GVELSXiwV3k2pE08RypqHUh/6zakutSbymJYuebVa5rkwqN
av5t0tV/8xOlOLy1/puSmdknZUGzD3GMaGIGnMrEZrgzgbyng6CgfXqFErQM8bxL
1/2EXggbcMpnrgs9+JtZQs9kRle2DmKH32ZpXAIDxmSM8il208rmyRmK/RfLa8B3
4cfrOQu1NBl7aMGDUaFa0av0Ndh77IDEpYkOuTyJA8U73diIhZbjmNV6PIqqFBU8
sRR92Atb88DYTJ916cvAA5QFoN9f6hIlI3dheDlGM991i2oJqqZM1JggNVSQp2UD
610Uuv/NTgheloPZv4X5SAGiVjaYyAeWdSCK49A8pxdn/DGTJuw0PsOGvnVvcPvy
lNtbWkdqVv/uiwqC10eY2cY69OZ0bupZgGWUDwrsHEy48BX/4cb5+exI+fLGnypU
MLTU37VrTHs43leqy/vDdlsN6poLSDQQdcwFk+fW6/4VyMp38Y3iF1Zegh4NY4mc
MgtqVdNy7ZoI1a87zpeplUBnDg3vMrZHCQ9ctlYeLf7rkefQHne4BPgqOVp/8yMI
`pragma protect end_protected
