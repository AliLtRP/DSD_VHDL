// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:30 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qUkTad26yiCzFATVe2umGv5+69RdrIDFC4RhMc7B4gteKyo1vdz2ADz8PadT1hv5
+5YfDfWoIalB97uNnRbJpPd/rRn3ejiwO+ca/O7m5aUhvrCyawYkM2g0u6UpdBC3
3ln7Lcpvs3bpaTlkKs3IizmnoiiApTEFcphRGCCO6Mo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3728)
ZGsBGW637BFqBwxwPcpyQLmHks1p1sJcqdeC06xomn8BNP9XzRb7O6LoNS/RgMNP
w9wUjRsJjG4PADj6AD4uL5LTmtRGKnCoQvjZEoZdTrPsszkohqYysPo49v7fN1C0
H5wpK29bVPhK7Zidp2W7p38dfH80YD4AcmARPyZcGu1Swgfdexmsd7OVp+RKqFUn
9oZ6IUT52ruFw83XwssYFUVSFhjgXCgIlZqn4hYysJ66VzBevXmIrblW1v9W1hYY
rD4D5gPcUM2UO2S2yC27xCJk4uT8CAm0tFOSI8XlH839jHm9EDrX0pJHJ02yIV38
Opel+DtWagU6ajNwTRSX3nBbgDutb6ALSi/+sImt0HU/uVmbn8bCyEp0MiosRWKT
9OZileMOPimN7La6iabE+77mbdFWR+Bpep3n1T1yzgVOM1Nr7KVIVKVvaEwlMHSF
LrKIoa3YvY3mcJ3ITMwqeMMsrGD4RM6Pb2Dm1XKwQrPE56nsuAWxZiq0LNuKg1Go
30FQR4TRLDIK1ZBYx7sow/TilFM65lHbtOgrcyFdTzKHoBgsjoYMiFUUfTBmet8o
XRPMtXXehA2InE53KehcgULnvCUSUA2Ll5zXzWNkV/mq/jC7FYJxD3oThEQIfZX2
SMhuR3wTLeIPsLIsbQM0chV4kVi7EuD8FfzFdIgGjQblnNSETvC3EB8gYl0e1SQE
kYWbQM2JBAyuXDzV7J05Apl/26+wVFFgfuEHw5JgoSrNpu5cVBLyDUqlHsDjh/Ry
OjTGEHX0IqbBy9KBw61OsbD9S7h++c8KqhF7bXuxuT6QkumppNQ+xjsPdRidUBAL
keKLJMqgrQIiLaQjpOT+wk4DGBeMbz9kWkmKHyQy0NwZvRVxgfNwf/ybqRRnCxPF
VJk6LX1V0T3PjY8CsOEtgRfiKDJvY58og21ICrLmHo+LeXyhLylaUFsFcRYxHNUV
GfbN44s6b/kG2P2nnSVUNpYK7pEDMraZcta+iv/QCzfCu9fa13+kiQSrE7oiO4cw
vMsv/s1Ljp23AgInfPphlbhBkdErgnUwWF7C94SbC/fhF/2EuaX+TW+1lsDPdf5d
xzRSMAh4euYDurVeLw7KvQ0GCO9GYlqt9zltlpeYw0BN7YpiFCgDId+SvhPQR1iD
qiJwyGW2RPI9nlbFkOJLoN9iSe1JYGweAHShqE3XmFwaC2KGoK0gyCB8UAzMIjCz
Kj91Ka2t0VILIY8RyYvR/bKstbMdqhreLRr2mXhUGiwqJqCgJP+cdTOIm75viuLy
RDWOeUuPSGICY6CUN4uOCjnqyAfyvLhXy4eHdm64aiMi8etFaLFPsDhH7UTgUW96
xviHJToBSIQd30GcIAPXlMQe1Q/YX98SDZJIDl+a1wopKMWCs6Btk0rdlNm53vxd
I4y8U17XojEWUcdmYgl7rVTH763woM3MCWxEYDUlVz+wc4aQuSGQoinfYp6485FH
xJplLCwgVdT3dsIuITC2yVOi9l2DAuaEaeX+nswSTU60+TL1qZ3dbax643eGPJNU
kV1HGYl68nbA3bh11T2gLe/MjPwP1i8phGFBcoRVkRdvfyncqEs2Ne3+JjHAyWlk
sLaopDLEnBhsNM11ZxKWJPL/AsMmYDuQb4KKJX2zrsMH5ZigsTE2ObGZHvITMyCI
TRWBlElnVhXA+IeXKauFW97mPaJf1lkNDDasH44duWUksqy5y0sBcKHOfiqKGX9z
uI5fkq4aXV6Lxq+r/T+GgkPe6CBOcKwpw7bVVKKyRTy07Qm01wf83VjKQCZk65Td
e2PfJwptkE+6ekLjHf9h135clJMPkPrc3UwCrI7iajZIXTF5HTsEFXmVQMd+gVcK
n7KVQVTBK+T1MXatjOHcd+uGoV1IkpqVDlnXF93rcRLQmFuFHz/j684e0BOaBqSQ
pSDLk0wi+2QieEnHlJ+6N9dmz54Bk6sE99rnfBpPRe4A2iRc48RsqDWfnWXsJo0O
MNJKbULxyjSSyWn3r4VZ4bag1ReXzxL6KDWHjkxoXkQNJD8m6lI4alvsJvovsSyN
xmkMNpJgEmQOYdlrgUpjm8zQrO0WshQAZWvW5Ilt4jYmE+pkus7euKyG4rsVl1zL
OXYoZynwrTvZPDPqJEvmH+2RkEXac1V8XDkEvnJr6dpr5KKu8OpTjnTk8bv1upE4
sLA86VEEL4Zri0rg9bQxJ6JFjPRAxRxQn3xM40VFmVn+pesdGANHwUFZfyR+fGDe
wmPhc3cxj++3UukMgDgdm0n6ScUxNLABXbn6pmgBc+XZ2yuhxwFXsGKtQj9qVoBx
YUdy48szmR/4CF7Vlcek4dDBRpvrS6kRX3RfGrTGcB0nGTnuD4wN4RVwX8DUdzjm
89zdCg5JJ/uc+HqMZ1tgvS6R7fthMjmkEu9jT6KOvA3DieocmZJaYrxy4gzKuFCF
fZOC61fJuKDRVvvPPay5rUGlXM90n98LDjqxDOQLXSwLzYWDrfAPUkYIH9jJUEfP
z26yO4HXZ65E2RkL8c9oDG++vQpXtbAZXLjuDUcMUbUcIy1TzgW78ZdUAdBHqND2
TZtVUq79MCHfkBTOILI9nYC9qTrj4l8dn2rY9Eo0t1kf49gDkoWf79cVC6IEMnrE
6n4RidHfvVViwT2ehFp9C/1A4K12h5vu9k4TTxMF1YD/SokWgrcgAtrWeh+WiArM
w8fvt0GKGfbY/WkGqu37mf+P+57Ac9B+Ba9+tYIBkeT+Id8yvQBRK6lANCpGTv/P
tZlIepDDJ6BT32+PSAEq/1/KZh8HOUKTbVUzahP5hD7vGKwqjBdZTH+kyGg2e9SQ
wm+sqtxXRvfujnYIa4+XWLfLZ1fHf//9A4BC+6fw/FzDCupripTn71/mWn+iZvRL
QWw8x3nlhVtLFzlTXmr3mNvPv9xT4hrY3vSRXBH42UBLOLIZ9u9uSEkIkr7zpvyU
Sn7ZFFjRQA8XBK8isrpW0+7Dg80/Vpv2tshOdYsUdZP7rD50gb9ICsgqjqyVuTNf
6+t4Dxyi6+D/jiLAhsO/3EnHvkhYUX7wtlbCmjZJWI6Z4wVYY4qapLPdqNkcDSVg
6gnbaJ3w9JVneM0l3qjS55BxgzAqAVBeruZyt3ZfWla2urKChCbH2iq2WN0vYHmr
/onV3+X4M5BpdOI+a1HkGNslMjHWLACDvaPyK3Jdi5IHOYSfrrksAthWyzP2veqg
V49hL3UAj4nwCU0+wONgHGUb1AGNRSAZENFLpACcscmBZbxAfQ/VTo1c3fNYYjjL
7IoOOF+SKJMc4+JDqUCIR9CE+nlHNTg1yeavfHDQcYp7/9ha0mP8Et1kz7cuG61G
ZNhq2f8wBTiosiOwd29sHuo98iU7IQTDOPiA7JA16LFAUgrCuwfG2v6miTev1aAO
VstMMurYkWKnRIwO+Qkqd+7hOeWrDDaQ7fU6pPYR5gn+HaCCzIfsie/8MST52Ya7
HhXia5GmPcgxmjEpwIFGJ3EFQCpc437PJWrDav2ACo+aRI7jPS7C1s6rAPKJKCLP
4zqR+g4/OV0GzCcWd/ppLbFkARxHTtkuIdfVNK6wcJeGIh8nKBMCEX2tQM5Yp1ze
SbviGYK0cy+eDP7He8C+MjA53uK7S/Qi8EDI9ewmkDH3/0lzE4qELqo7rThzOZWG
GJBbx8btskFspt7ut7qtKn5h83IeWvVLXvUF7AzJjUoQF5uJSPekd1FXhu7aA1tk
1A/Ola8paGZNl2oOBM2SV6koS2BfBFnNfOQF1hXR3ggrJXyNSV5YOvFqh3YgzvUp
AuFxB7+Ub1ZoYWT7mG7l9vbfOikgfE+GU0Ra4wyhUkZKLRvYY65oPazNC55sHz0U
P/3jPWZ2w+jTzoppQnFsHIEErfEMk224yAmoUNdnanSda3XYpW1c/9vy89Wg/10z
e2PNUKIYjntgswNcWPLm1KdGjbJWTsGvdc7zG+6XktMwMYSx09RBTCAVuY4dZP+1
GOIyloaa3YOkuhdcQQBeIJ6U6dap9p8HQpZpJ2TgOI6t2OC59a3AYO507oBl4ng4
D9xbHhT0esdo+7UJXxzbXVHFcdM+M1Gs8f+jshJUbZn19G03ZiueveZ9cCCmCWjC
8930f54+waRsxVzcI188vgCHtx9xLOIzrdglyfDcTWr0RJ3kQ1hYmxwbG3wELMJK
XdmuTZaEklLapRpchDA3ulOQbYkxEMNX/J5EZEwjTjzFUh2LJR6PkVDV0V+FDH9Z
TXmWJH1FABzUzjAr6bK4hOOvEJq81Ut6NxF24LwHkeqSHBSNbrSTv7PY+BRqwlRi
On/xpkuHKUotV5WPwWFrnK43sbwMtGDruSiiyob3yHq9Gt6HygybVpzYmmlF4koo
2d9DgStj82CXncSZE7d8woI65quht4ydQrtIPnjXiewig9iiC+xDbgTz6w7MpWof
hvAOl8vbKJMXBZGtmmclu394gtDXKa1tnZLQiJYiaHn+yuNcjVqIi+oTIOmoOodN
KGsOWfDZ95uLIXC7XZemcCI0UXqt2NsZgLDE3zKN6y0DnzdO7AAMl2AYxaydIcZE
+zPJljNePL1ZpUyDdQooPOjiP9xroEaq3Pq3KVLMWOP2IXnaxfWj0cMga8Iez/Vo
t45UT5+k4FIOy+PNPcm0WlijiTwr0p6/KIdkIese8Bd0gKAMuZ6hU/yUGwb3DBlD
1slWvjP1w0rTwJWdPMYPcgDEmMq7g2sYm/w9nFC9xE4vK+98fhISdUCQAec0Lz77
aRPGkjC06qSGIZMVRkhfCJCdzHUfZ0U2ORH5cGWRgnjaYBFTF/jZfezugak375yo
vPJZMmiFo3zDluid8vin9r0RAPa3yRqCFKBN3rrLtyeNguLvwqhpmEanusFOHYUO
tef69MX19Eyp6j+6Lr2izrUp1sPX177sd777W0nom9qQ34d6aM0m971XGbOdPYsZ
nJSGkBbJYxhaJpS3Tz/5kf6LKQyu9a/qKM5K7/Gl6Cs=
`pragma protect end_protected
