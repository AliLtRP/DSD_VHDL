// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
lRdY5tgT6dP/B017DpR15B1c7X1xk21bbwnaMQTVO8U1eczIWRXYwRQdr9/C+gyFOmKc3a9kSaiz
9arSQM95wvQ4YFYSv6z9n8BwhG3cT78WooDcVZtrHytMtCW8cyMFvDNnWvS1yqJhx/GSLmlTVIVs
8Me+aTp554dik9hGeS7h86JvnrtmQF2iDCrlfDgKRSx7tglu7sa8DYp9eG5o3eAWRRwpAIohgsVC
Zz1x9jO14/yQ9/Ee1TB50S6+/7ghY1n6RF2M+kJUxKLA795qeTdhdD6pYrw2WG1THOiUCPq/dsMJ
kaTjG/tVmA3rby/ObpeejDxsFQ3z5sJv2Sm1Yw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
gCAcy/lMBn9yy0DXkTJ3+95ztDb76Kd5sXfmeZqJHhK3VoKkUwtpPLtz7GiobF91lXr8GebTL3/i
2BVPLA0OdXe3R7Opvy3VRhisg4f7iZ2temm2pZ1+AjlIuA/Z9xz77bkU8cqMFRoAZYy5V1cN7GLx
YmsTa/wnMMPBUcXW5lkD6USGO+y1p1/9twNSaf0apuGSBWLzoXuszLw/3On1nu2J1pKVWQnhVzeA
BasQ49LMtxt3VJ3m75MFkh0I9bCpZ072q21IinByPRD7UN3yjKUCycyJZpV6xZiRPqhc5yTfoV6b
AZz4LPBYEN3tiq2JY1x3hkh94FQk810UMkhgvutDcJ60YnNUXY0ze8Om53BaVWne5KWGk26P2aT8
aeTi5la+ovW7f1HdQonJGLoN2okJtmi99PLeuvoc9PgoteuiVzmwcG+CJTXv3nXsQkbKcezwlDTt
udrnC7B3YunEhui1f0HvJHI77Mz6J4g6Q+RDMNk23wzODOfK5WiNVMhDxw90vBRuAFyGqACz1ov8
J2QJta0XrxHokkEGN719kUkx5OlEDWPDQfsOBo0p3U+EYNTwKKkYoLJIAp7TQi+TY3I3UwFd9EH4
xLPLvlT3fOo6K1ST6LQ80IxKFVyCS1bSH23GShyTzDUT/q+iwtoomvKY25d+KzQvEcYst1l1kkid
x5TPgUtYof0bgzsroYctwca2rS7EVSAH4V78BS1Er+H4cR0h4GAAquGe3noMRmh+vZiMCV33J6F4
dHQZZc30S5bRjfznLYt1jD/2vtAX81azVvSnr9MVJ0x9+kTxIzStYC0ggDzOS0g6kUBVmoKO4zAR
NK0hK3Lx9c9WtxUKqXsrVLuLQCGj84FrnopkdK4SGT7Op55hbZVtzc/QHs95tU7EqQqxGnWEz9Z9
94+vzK2o9q0kDhDnNs5j4glup3vyqWhGQ+zBclZer7Efp6ppPdJoWY9nMqiVeJyQsvFgIb6a2hxq
NlR9G1orjNxNOVTsTtbxW06rjP1KjGlzPvdqsqSawnYiFd0C940xT0sz7fPDY4fQE6maNh0+2/zE
Dcbn9uy9OgMxVNXoeBKp0qxQZwxWuxwwRXc/OAnFO7+U/gWU3hFxqTgscKo0YtyLv7XIK6r7poL5
RpdmskTFhqbaEO4muMHCv1jxenqRo/73XMlxFtkW56I5tDSQ4KzioPWMm2hcPmQeWVK15tiu11IL
U9o0vglqg4I2YvlzQWHjWl6GcE9Ipdan0CVo49PGZLuRttw5kOwAuDAZ3EOOzcoxN1doLvKuq9wL
BX+JhVVaKQ/h3rdym3CUpN4293KDT36YpgwE9gR7gRbDgxrqCBdFM/2LpPu8mPQaQIf9R50lY37b
NCwB6RMxkUhfG0TAyFcetHF1JaMSzWgpqzKFjH1m6e5xRT3FmLhuNQjqc6rSKOsprqugSSW773NC
prS6RxF+NRB0fEH6ud04l1uAVpevXPYto89+MZyAh7OCRuRlVEawhLWleJHF6YPbxCslZv3YI7nL
Lyt4El8mRyZFP2VVMBjrST7ZmiaLy6ChtZ3BKdB2M9TKCGO+1Sq1hd7FibYa4hpckXI81mSHV9fX
y7sxHG3QndkAKP4seb4M8QyyIHfZzejBLs5Jsk/WlzFsCWxSbSXB4i6QD2XJygC4lEAWyXA9/VGi
ROZvntRsUaz7APM0TZw8cAjKhzRqZKrFMHRcXuN0EdBjT5xaZUywDubEANpY/5fw+WMEmW7G2QZX
df1vt3eDqyYkBzo1lrOwpATOxseZLA/yj9mUUNYtnv/+zfR7qsoHKMA60zJpHUcCE3axK8sJtSxC
eIUClCP+ne1zSmLAC+4FtMHcdtQHrIYvhA8IrS/qOxKDTkp/sf6Vk0G3s71NbNItzrjYXZbSlJe4
tHEbepXDwtGwvxBEQJnYBVYTdoBuffREDDIgQOO++WY+y/WlMN0a3a7JZUGTpa5O8nwHY8vQiWsG
Zg+gRFr79QDfldyKKbf/QBBw8FftYTPq1LhWd2UiWwIzS9cz/sExqlLbqC1YVBg0vpBZqF9N8+NF
N5hyp08JxyNeUBMkDj73hXOthtNw4WK+HIyw1PcBm3TqPnklm2c61qWJbxHa5CJlqJU9O4F4UkdK
xTQySplOjku2x84FJJfKUkQw6GooFsmwdv5jtKcPEBPHUGLfW/LLtONP/R+MeOR8JL2vprzDz2Z7
GJQ3/mKzGyTfuD6WPhOo3r0nyFlVS2CUC/VXK4wgNx7KKs0zYdR5swHubavEHtnEv8Fwl0yYpe38
O8wLqgHOghcEHkUVHD0oZk/QsaLX0Rki2uoydcBoYYJmGXIZECZJm/HYIp7EDdhR14RDtW/MidMJ
FOIibgEwpSBem7ktkkGaKY3SuFylhm58QLsV2kzWoF3XIewE4O40P9ulZryKcG/VP/OVQsLcyxbO
1jr0Nsmaf7q12CImykoubYo76EtrYtG9pl4iUAZVB19EGRFjkSD0TsH1SivWU4md34RWp1trmb7H
+3GvaH1xgPkXyrVbu2Le1nsVPk1k8ZgVbFuM5pIlUH72bgRKwA9P5Rvde2qy5zj8/7OdeTn06GHJ
ooaPVPSZlMXzML0uGO5en+jjIA8B026EFRq12LfAGWyFjoH1sb9KtsMNpGfjG8NOHNoigQBVA6FO
VoW/x5cg4kB521Cn8EK7kBuba/fEBrOhdB9j9Jdh+ORNiY+tWVulSVDQS1kWE/2MixOY5gmkytnE
FsAJbDUefCv0hexcN6TWUu+YZCM5hlIF2Sd5E7ltAoBic159AffJiZkgv6JP9NYamuJB2LwVAeMa
+W5NTiyj24x/uG2S9N2JADEMpuDg8lIBrytx+VsTC8yXeZIeIFiGabRVaqCzJo65STFL7z5a8PKn
FG/4CilhKCC16Jbqe5bf1428Mp5ICVKnC28SeYjeQyl1S/mBgAb9Hde6djk+Rn3sYIuI5Sv7Ttku
L8HrKLGo3wkJZiJmx3wRYsyz17CHYxK0zgPSYlC8nn6QWvW/F02KcFbK4VmFEalUFlze0X2tdFlN
ftWeUhjwQ0cWt8idwlPzLAPJrOkkNlY1HXZLxFjDZuDVcDqs/BUkW9CUc/kdr6LJg5jwrkfdNaOG
60OCWLquKR7Zf+YLctGAQaGDFXJxavWCCX5w8dQL6kLEeAsJc4FtMleUtm9foRfo8P9e+xr6BJHu
gINyeB7xi5oIMaL8Js+1a/rasU1xSZP1uT1Dt/BRMgSbaF1D0+JwgXcw5rO7vP6HdqMLd8KCVuJg
4HicpcWlmCacu9HSFsupqolJ/ssef0l2CfaEGkcUiWEsUZV6Zh07qGKTS9Q88OBFoMZ7vSeGRw1b
YgTtaqqU3HuqpwNDS6Niyxg1CxzkB+8e6Pp0nBVsFU5/LMWh233pQyhNcS/w+RkjJVy/m3s2TRdX
AIquxSwGZhn7eFA/je7KYkd48kByQGMpJafxjMaTbueJlcV0tZsONLKJUsbf9cddykwdgJg0jctu
kxSSpnyhAi9T6O4lPMW9LB/NR5p4zMLsOAeQUZOsroh6uLhsK+bG9laIq39GNFD4NFfSxrXktbtj
Iplrhd4c03TaCduoXIZ/44r7EB5kztqWLVqWWsRAPC7d19WDWfGvWwfIzU7ezgHIymCnerZJML5h
AxknotgnLpi0X3uyG6HTqPuMEQvEW53rd057tmeyYUDQEyvk1mL15EhO5jkABKWXYSh9NEoKbB1H
jKKZyKuBvSrBFkd93s9wPoSLyxMfWSh436PXCt52FtMte1i2N1xS4RI9g3Hde/vzw4V81S4U+bLb
44sBdov5XyiRfrSFuHag6ybmoajycsjEJLghwUJtlFyuXqdEx3gM6AtZXreiAfnd6d2XZZfq7xTI
rv8shz+Wih5iq5wP5kFwYnuBVz5Dt6Mwc9WWgVenByViQ88IXW1P5Ii0VafjjSVttNuT4X8+n4KQ
Ele4ANhuSZm+gX9tZEctLg4ZJeiM2kLRlhTtLD4N3UvM4uQDwGg4Yhwwj9p/TTyQfa/LrPqQJYxX
dxk+Kax0QAp8Nf7g+Qa8qIjyXwKtPn9Et04f1tTqHLv/5vKdVSVheVgszPj4QzK3BIIrPUiszNPQ
edM+4xcgQrGctsCvEzg15oKvmJee8YNFfenEp8v+thqGxRBhVPG8CtDFN82djyF8xnJs+caQa+Sk
B32R8zZDg6uEM9QzMF6vzm/nGbYZuexR1cpjjLspZrdJuYTlpw3iHCQeJ5xMsWyi+IxXa/w2pN7b
JrsoZXXYw6azTnANX4uhmnGijPqr8T6kuZoiUZWYiBF28YLAdqB7b/ByS/s9zcHwoVDyc7Bdh6gj
DV1dMYXffhoTNBcH3U9lKcLSUXXJG5WvepR7TbgS0OR2qe1BSNxOpLDF1FyqGu3qhFZkrHdGJ5ts
gkFF7Rut8BBdwTxnzi3DHFtubKIJHKoVKjXPUORLq3b1Jd3EqF2WZfm2FR//lN4EYOxm6LqOrKfq
VYD+fxlcHCZqar8WYm9ye7OFdlo50lE7s3lVPfRGuYeVH/gnzHQivgcBe5CmWoEEapCmiIELHSM/
vxWJwrfLvg2JISdF1zUn/w+PeTbsGsRu95HzS2Y6/lIxUDx7zSaBqH8woh2Gh8nBKYbGU+kLbNSo
VoYcFFAg3dEGFPgu8z9OY7/RelfdCfEix7VBWCzarM+sVJaw3c12rAKT3P2GGXfKrsNurSpHChIf
DTYtraij7IOm8nhA03LFRp9FvO/LRMe/B8brEQnMnDR2V4aCNP812jl0RaKNqxqLhrQ2qiFg9E6C
hbkrXs1+Q1LE1aLm2xlKNvNv+XzIBunhvTRJuhsGpA8M8GtvSZX7xnB3uXWtRzbjkjKACjXJtD5n
+Q4P4FEEYoMjB6I6+G5Y3AyDcgksKoH8eCVzi470I6Z8eXOqqj4jPlCFC01xCRDSU6Z2bk5MPXrM
K9kKxdmpQQDxnRXUBQ8IHQ/ugH85xX3mwwDkVwvT4zZAwaOvEDGSI0g+6a72e6iPz5d0WQaTd4HD
a5v9i3kahqTRcCISOQxTho/AP2JT8ON3WNdZRTLhUsRE/BAozlQnTN3M7CLpFoWolLH1FSDwH4En
yCPWnu+xheEXKr2gChWATCyrXoSb2dsRG4vyzR4eolODhklCmNC2zhimK4dUC/BzBjQQ6EBwRhfN
e2i2lIigHxvUQwR6V+/ADAE/DKpHNV8COREcKQRmo+KiMr6fAztbFl/QMs6Vt/iJK11FakFEXKQu
EwIkzW6QwvhgSmnyoo96RxAWaSPG01R9Jm6Z+04oKI+DB+3bmjTBuMBzkc7j8p8jC7NY7ZVlh4cy
w7WoCp7CMe6qKRHbtMEdz6ChQt66xPEzvGRiDzFPX5FVNOPgx/loWZ5x8s8egeRYE81AL73YwaNI
Lsbhm53u21vd6aKtU6K/L2mLBWJiJhHjOy5OI+CmfBxtUS2YGuAd7UanMv9vqAmT77yswJ8TNT2n
RTCt0q5py2aOYu8gr7z8vAPr9g4dJItANQjH/rygNNlDhvaMKxx7/f8PruL8jUKVA3r7cQ0qCdvX
ybT/RsTD6+7SnSt8mQLjNx7LI8yGaWH7rXRWCptMEb9vwlQuKzcW/CxlArGSmyBfsFhXw6nE43Og
Uy/7UI+JpKmSprYrrc+XnIcQEoulXflh2BHB7gQAldcsJBOcAwSNYgxc3ITG06Altw7DCzcpwRly
8N8gOu4OmtlEuMGh8O5i1HcXD+SyaxIh0BMKS3s5GKA1yneSQ3SwNW/u01SThjSXlAnG4pbJbYI6
v7RInEUqc5rdWIoWQkW8b/2fBbKKpe1ffnUtRPtx8t1ohRkIPQWdiC+lOe0iFGy52cJp6xDsY1QS
Setxamuj3WUkZW/Hh1MWUb+5K1sAcNXxhQK0n4w/OaRMrjYRHTdphAIUuXIHoVWfxfhmmfGIUkGv
cR5L7YDRPt6Erb0P6EAKFujcAqEwQMr+FdvNDneifqGdpldetSCXY07hh7Dntiajwjjc6lfMhD1D
dfAO2VsAIVNoHAOvvOwxSoNKf279EC2SfTTEQUI0Lj0faZ5381oHkkFD2DktxS8Wa5z7zhroaq2E
vQtvhY6Ocgz3DYH9YzTW5kYhKaEadTjHrQifmUFG0vTdCteUYYQol5yk/x5dPyQR2ffdnNA6z14X
WaKBllzmWwk3LxMO2LYj/wOo6Q73L+bPJJ9YrbFWgiUNIVeILH/5kI6Ber026Fei1lPdzsA/JW6W
T92zylQXL1Yt9Csbq4sStJoW+IU/PL22QCm0utgizaDKvufDISzbFV0kEhJM5xkL+trgfZ07t6pv
8ealjaCGC7asPLz+yUPSh+wTMwGJ20CvmBw2nPiOAxpV0yFNHq+Vq/cpXvoa35Ab1jbXnLBcKyBb
GzzUPzqzxWD+yvjDvxkNB/6GCBvf5G+O+ppyZR5US2ENzR9YLA3/hUTxiXMuO36LYCN0yXqRXFZZ
O1coQmWbC+v9aP489Pfabk+26U5GOZ4JaYu8A+NU+/JC9QuoF+F/miprjRHGG3mCwdnIiPvmDwQ3
jCR82EvUlQrYOhvS1sbo41qWk/1Op6Ve5uM39RLNIsw0CPtVLT1YbFNO7AgR4hU18Ko+I8ZvyI1Z
w6NqdLag1Y/WpmFocExNTe+Otnq5PqMkhf1kwU6MO8w+uVEN4nB5TuxZLOefm8w1IJ5MnGrnOHea
Jtd7+kWTAFt+Os+ypoApE4j+M00kQaXY+Bmx4A6F5BMxi0LEVlV672OWaC6u1zOpdW5c+tGAqTy9
wn400Uy/8e37WZ3fKEsXNDk7jFe/u8x8S1nTFvHlvegH8DjkgPxLqFxKVcWMdpGihiV0Bm2gkmfz
PJMZnq7QJG3UwY4gWr68268nOooJ0g8LYM9TbpV/rIBthUXnPia+KndDNncpY2305kEMyLMeV6J2
UGdabzcp8IGbFMpwW310RaFagwZv/XHgNrog6q++DdmPHgIng9MflTYvNcd1wSWycNARlH2mUQvq
7jF6eirOQ2lMLzsjUlSaLA+1HvR8f+KewPEqoiDyAAOVh5Ub8gHX/ws9jbV/PAZROPA+wtjas4sY
FeOixrYZHM8tlSyPF8RnYAfvoCvLgPl0eNaeV/ssHBWoS/2AoepCJLq/pnY1k8km9lbi8X6RCdOs
2cEkwfuxcPtkOZuOTmVtT153YELtMObmc22s+BubXDpmhG/AWlqpAOrDUUSZrtBUPD7yM88g34fA
BaPJsb0ZAflI7EJU/sbm+tF799ktpzYfQ7WsT3x6k4KryWHTY7KuxEWxXAVnYFtUemQcJtRO+ZHJ
q33RaUISrpFlXDfU4yopkqvkgdWsI8KBk/IHRsXCTHskX9WqM/l+taYIcBfIiifc+RL8GX9o8fbz
xbJxhmz4TXxgGlJNiNfEFVFhS6nmRCCPj2Zci0k2m3yUEUehvC33F5G6ZGCAKn3a2vuPXR4BR4BR
CJlyetXMAtyQ75J839x7spbSQ/p+55OvkBGneK50dlDUbMFmSJ025+3vqtOXjWAvBDEhrw4jxwHT
eBH0aXuaml/0DHWjqrYLHGE9wpdQsscA3ATdNwWhf2DybxNcsj7bgc6hx3hj2DUrrva7qJFSqiA/
OVZKanZAY75sWgsr/4Bt3B4daVhLUrZggPTAT/4fhelkLFpr8uFNIhBbMwG2X9sKoafGsoCzuN9L
M3Fy6PWj7zn5CPQoEnHPdXgn+voexsFKsMDbp12VYDJla5BXylHWZe+7iSu4bOoKY2gZboc5e08a
6XvFXyNo+9LH/D6jeLgFmDDg00ukMQQF2igmq9IZVFYHOEHzcqV25/ov/f8RRhXW5x73X9zgx17t
xDfBtz0Cf6NSp664c7NXJI6eNQGfrAYNXRJ3yZpBuBmY38DrYW/dm7zyLhLACnPSlGnpfPcvvbS5
vyGuTGbLY6PvYjI8onIIeWB4VyqlbK4RsfwtrcBAb2n8fx/G9gXvyMCpaTuhYBvIP+EwACtZJP9r
pulrk6YL4U+xoy1MX71VFpJYBWCqvqG2pIGqmHOA+Iq0YihbwhqvkvSuDZUTnX4EYE0xKKE4Xq9Q
oXNc0k+48/oA8zL3lUjT2m87KS/Kp3JpRe5e5ufxzp6J5HgsvmKigwElz1CMYy2Es0YykJGDUPRp
UzmHD+1itcu5FGcBI85/dr6k/DF8gPfliFhmBMg74BZtqU8fEPz3wZChZhX435fmy1vHuqf2DNs8
0TxtqjHgt4qg8tJ9B+0w/ue/DxrcdKNxiIpyTR9U5CJk/O0kRYK+wIo/cgjz8rRCkteRQsnT/YZx
0KDPflHNqOiFEdQCI4BiPO/b22j9Eghw01nD+UNedYxsGku79vDfwfzGjpIXI1j1AGPtZPIvVRTs
rk7P9nULR25OqrP7ocy+7Vn1FBKf2cCLxWnUO90rbKec2z0d30yo0Q/LixHyGBCZ0hmjugfC9u/T
71rGSXwTIft9OEprnjp1cBYKtVIjT+TJP13tDMuw3lRnORiPkcRyHk2+Q85VHzGrU9KSdcwRQf+8
4wPTOv90LoL+joybwM1W9XldRn/pVOX03xPxlvqZnebZZoM+G+RfS7yVnyONvFMkXol0BZ9E0CSU
QaYs0FFlkUtw5pU6zMc8Gxm3eRXSGpAsax5bReTdKf8Lhutl6tbjzlHcIelPhaeIBECAKXr7/PMQ
BJ+uAgYtql/ObknAVn33yteloiyor7ZE06dfRXy7FhL/VCd+LJhNk0X5MwJvGBfP8rP+jjnBIz99
J9JpK8SXlLyfVnURRsectvBPQHhyK1ET4rJwXeAORVNBgKNRseqRKpQf5ecyKIF6q+3lTzhP8Uvz
89n8mqFFE/CTmY8U4KM5A3VT9Kawb+VLfZcP6pW1PJjrjpOfdFoRquSu3FqgVEfpFRi6zegNhXxc
5sF4AcqMsifcwBnVpY9yGgGUDXYGBZlKKtsQYGg7tixXGI0zmHVg1kUYn+daQhQfrxKk0w5jreFu
M/Tcf2gPn1YbJipJIwPyUhIGzP38gMSGUG4nKA/3ehirpK2l76nxop90mczZECGp9Jg9MmuiMi9B
9nyH+8ENL8E3wrKn4h6E9VsR+Jfuu0zkwylIG/V1S6FvciCX67Dpx4NM2xrrr0ZaavhAr10Z8KAp
d9BCpQ/efMeYgf61NZ5euER6SM5sw+SlgIY7y3qnbPWWkwzJYvxHIluWuRGV8eJSkJT8ALw6/znR
McMzlP0Dja1F4T6gHPVXCmu1P4T1UGubgv6x6pyL6rUH9I4ChP6tlLmbTI1QAQ9gYk+WnQc0Wb49
sz2ceDwyu/wNC70YgdEuRT5sWUereZRh8ozkeMUMYKLV4JhIMLNyqVgy7Bi+TrPDMuT7l2N028/q
e76OsJisWMZtw8dEowdLOlftE3KifFxmCqlisMy+AxRzsx++rwysanXj3+mhcIVdTVVnY1+T3Vvq
3FKQbwgjdPo7qxt6+HUwy9nsKJvfK0QjATzm9G02JaMjEC0Qzf4RMPuOvKo1sKB7XlPWXv2xN6o0
c3pQuLJxUEOhJMhG7av+aSoLAqsBfWlR0QyNAqweG9oNG09uFAb/O45eNM1YHHfkj3SX0TQramKk
vrNvi+Xw06b8XPUDPfciN0fohngZvHyzNYIBuQBvNmuhzgKEdaTQOKwNjqftRXVO+AqDL7IB+vzC
ms/g7xfYu1sswFpLk1cnt4t161Wyz+YuPljNma5AjaA07GOxwRcbQPYf/byntqZn/9gp90uCvTED
xpk8r0EEV1Clf3Mv3zM/wwj6BXne4QcDEkv6NsM4G2YjQhQM7WCq7T7zeuVZnKUXnZHHLvjP1kNm
6ytblYXhzOoC7cmEMlT+JUSLuPRfjCRSIBLlsUkyA8IvtZ3qsBqIpsuR4RkcfEcejDy22WjDw3Jb
aUfrqZeojbKoY6rdwiTP/0089M+F3YpOdJPq9NS9/r/OcrF8qyraXQuddABeL/wrFjXWE6xHBP67
y/HiVa9FF6d45hgTvEWX3vyw/v2LUENvH1okJcSAgK7bLRCD/Kqgj1xLLGzqlxYoFxYuTBQuGegP
xYdRYfN2vxx/vz0zpMJefZOVSqNLfyACbxj1GQ4YD4jB8xfxyZjUM06kZsO+yjd7ieSvYpZuzNO8
MfX6+Y9WhQEE5I4lvraR1wvYp1deDDdBoGBm5ZOF9savf2gKVHQ5wuGA6lBk5DS2opZ8rSZ2UorU
n8kq4L9q2PcfkIIwkiSZ3rr/i9c4CgR/uE/9e6bn3K84Q9bgCZFSrJeqg0LfeYnZN9GG3p0luFX7
IV4XhLU59LkP1ZTmPJY3CTkCbEm+Vktby2DaKwsMQnV0c2SduUtE9Li4Osd/ymESrYtNajUea8s5
SS46T3aFAP5k6ULLd1bdKUxs5VESLS1TKEAFESffHdRnHvjPsAtKm0+IshtsTG2FoVr2BeFfCjSH
WFMm5spax2B0TXVuq9UAtw3A3ZgZuOV2edsT8opHkB9M88FifltoZ7AHw84xIIPQXxbxHT6Cd2XF
zJPyfMAcnarbTusMR5ts1HW/Gw6Sfra6+dX/BXmYpq6MgrPxEPLDnOcN9z9+bVONQTMmzbFzv0wI
Ha8Fr27yXJQBcCbnMV/2x2jxbtZCdW5g5uh9qeexuOy/fUOBjOgz5Befj9tde9lFY8KYNg0kSvCk
PNvjZW/zxSlP5Z73xYeHlPC+sUkmrBhRl05rNK5bxe4vCo/jraf5rSvCB24uUEoEmKpALxmfjKfJ
PUoYf8xJFqBDsJ7xqos0fe2bdVj2V1py3il+672MWuH3iJoY8giIEvEYbjk9GTJBefZAf0iRmXir
S4njdHDCk/d3CAoQUByw2QZTLrxm/0E6LdX+jXzXuvbg+8acpUUZh1s9jAmc4NfHsQhW8PpwMJcO
U7N+fpi+nEx/wUPorQpOAOo2sVSQ+HdmwyzNyFCe17fOSHeARHO17Jmcn3xdNGrDEC9YX1VUmbcc
M8lWj+aDIqTcY7iO51UjtLfgNrhIm95CumagkYbSfsLZ5qKWW/qGhEWuiRSBjzpze2q+u3+6ItYH
HhGsdGKyp8/dWGUwd9CzI0/VmJQ07fNYDX/2ikMuUoVUPBkWuBAJMDjlibl0XRBV0TNaQUJiWxhI
E5qq7FN/f4OgKKhbGHYrENGeTzbpOeFwarUXekR5Q3ZLHqfPLR9FLFrOP8scezoYqLQLhat93j8s
CU+K2cw/YFuujcuwlcqpqL04w6YdsT0QV0n3uQkbCIUoIO8BudiNLiSoX+ZJrVPOuQZiYLhajZV6
JwBXcUeeV64JX0Hnuob2A4NVQ/l3ZKKMm4uB8HDaTIEX7AEo/bchsU0eoxnQegxtWQOylDK44fne
c6ajcnpO4r/KxPiDWgM6L8S6lMIcuM97QI/z736QAlw1FfeACBVgqKjiWgdsGWIMzHUah2v8f8mk
cRjpRGByRB/4AtASUfBqc/u2OaMYReewN8D48Z6JmvX4Feqb9TCibZoO+OMs8BLDl7EEljiJWO2I
DvcQyRIYnyxqTrFsqyjA/5wYCZOmfi7Ezjzg4XVRbyH1HCewXcPDtTAR37bwYyjqh45YzTHXt8Bv
te4BJbS4PDcsFVetDzZmlBJKPGOhz7286IpmCeJDDk4k4KtOU/QFBxUVQMdway0IrtkfTs/Bgo/W
3Ym2Vg8ST6lR0EOlaiXy0fCrGK5JpQ1GNu3w6a13IRinQcLCTCLaI2Ft6sbLhXEVCprgwpO04+Ub
JYu5Wuk4KNStXh7uWvNzN1tIUMAN5zC0gUMTsbu5ehXIYyqVGVUSpRWMSmYvjLN80fXp/qqOYqe3
LR5NkgTcyhTYztdEg6ALT06ts2LZxEspm0Tc2oV2iiZYYR0IfbiVjdySRegAJnW9mGibnaDvYg97
FwP7I87fkXMckQ2ZHNRXU6kE5aL5/R/h1JCL/jDNi35kdmphdzzsRT5g9FWI8wUhtDCjWNHGVNze
fp7mMZ3i3EX9krO9KZbLNQSNFMlhsCpK936mfWa9iiDA/GlVZQwpo4V1cepV/q+6KrCW2daxkuMY
Pu4MknExh+3w1JoD0hEzQqsdEmzoU8iIGa22leSaSN5MfAxhRdpC/rDhxiSjTSqVLTxDAFtFAAQ4
HU8zl1H1Vhbl/gxZ5LAqtoKV572C2fHoqCNSivjCFPq5lSdtqjqreQeHWx3yI6bFf9n6Waaj6FQ7
e9PEIY374UyLZm/HnVRqbYyBmuYENGaOroRGwB0m+OWgrNkXlFh3kJYgtQW+J0fAsWK8SvWP0Lso
gr1L2tMRt4htDZEtA/NMXIFC66SENu0oguhlutPbyfcj7vJ7FrFoRrAwlPMiZGBecwSTSmJtA2w9
pU7TDOwEyDeVNOYUQosjlHqUlO4Hv0aAd20xbCjvbQ6pNqlPsjCccECyw3Sgda0B40MZ0lTvpra3
Sop2rtApU2WABOlMwtKhJeAZtdPO5IRMLhzBJiLk03rWXyt9xV5nfC8uxx7ZirHbun5d8qZ2WkFM
ab8542wy4rPvD1Cfn91dMw5cndiMre1iBiGPf+PBejwl6wtxM4BCktWtDF9dov/TqVI0w/UFI/OL
X/5+MXHSn01uuoYIG3FRv6EE8MCOYIT8X3UaHToTxjhAfM6nRGsowpNxANHoxI3SQvHzO29tQcY4
MgW/JSjHUpRwUlMcxpfNHBFN6s+OGkWwz0qhgvpYNS+xCEYwB0U5GGqTJZW9EGEzaCDw5qaoxQyQ
IlQqnkrNNB+OPjUj6Wl4lqelWNU88LKoWsjoxt0DBioBwjkRaOASIXd0HXjwWMPFC28TiTW41iDX
TMKbc59zw+nj8EbUdMOaf4m1AgcFCOCohaPtL9ohKCwlPWOjisPVLWJoYhAwyc8pi9KWWb/2hXh8
YHy12iuIN55rwShnkCYZ/J3PWwNPw0Ex3a68tlkH9pq/IaK005wcizMZXcsxyBOgr1p/C5XoWeJj
3LjzBP9zdLRGNBv/yJQ7u5agLdn1NYEFG3YWxX8YDKFMRKWGHQgK7kjkHFiLpg0cI8PfE/11GylQ
KURSJfFSB3/ZXtoW751WVJhXmUiaH4qNQDMvz3r/uGRT80aQVx+s1fy6ni806+G3LOtCl8kAqfEC
GTgKU8HeobNL1rPRqnlbO/iFipdNzuN+GBaxc3NfYXwf3XuYkRuP39mgKs55QC+l/Jj4DXObMFhD
l3E86IQukgbxOHS3hJ05sMb1tpBEWPL7Vn3RQpNrWy/OnEMdOxZMBYQxgBJ6klbFeMy1gdW0zGA1
X2ZMCd+wmwNmosCNq1CgXUnnZ6cEqyj5o8Qczt+TOaOzUyD3EA8KaKie4Zn+D0fAHk0nE0IAgQgg
88BD7CWHSVXFI/vc8Jycq7LVCc4k3seO/3wbtk6cvoo76Ww7yTKvO33wIprVVVk2imovnBy1BTLK
YYGvG6n67abuE4mL7CnHYAZCw0mcLSapLjfyNphfJKCmso+gxIsN48oH9HbQpF65+wK1XXz0n2Oo
Nbx/tmhNyUJzWEelME0HnZfuq0/YnpKPU4WRotv0X/7kvdl8OwHJ8xhY4dmv3i2w/z6eVwwYMHqn
gIyACBUs/tDjmfaRVqLT4IfEYQeEaADIi4BF2JBnW3lEUSOmTfncproRh3bwoaVkla5YKP0Ut2Mk
IV6UsCrRNjHKpQF+VREfAVohCvG66mjYaKPDinDk0lSf32HrxEzhb2v8TkaL7mAjblry2Vt72XZm
ohfrsn3Hq9T/9aOHYPVmO8PmLH979kXxOdYI1OGAAO+nPcSVnSUf1TqmIEVXLACFH5O72hC3Wsr3
YkaRxsuLfRrj3TAQoYq9ZE03zJb51cphwUBOQt1y4Savo7lfKPGOmd1Il7L4fQArd1klvdn2oz6b
pYAKStX/ceZOSWWpdYWDL4+q7i42UBn5N33gZGcYpB/2rYo2HW/BtVZEBwUL5e5WDUxEUJUgsw4K
QcWqj3K5UcAvIIrnlK20QRbEqaUj1d7FAuqoMJrdnmBi0dHRp3Iz19dpyZGBh3c7xJuNPRcGskhC
t2rYCcErFNuRSXBXgc48CFffnN/JklWuWptiBURvxoxJT/Q4GTz7nyXSBCJXaiuLPwAVf10TLn1S
dYmivWzX8BcjhrOs/A/5dPFaxvTPyKzLFWnBNLrtolarD35x91VnaHKLSovbyl5e/3g3uZiutoZ4
OMCrRONM4qBq/djqdKp4OThHpKbi5c+qaeWk6CrJIq4Tcmic0TfBvoCCXVmBAwaNnrBgBCgaUhzv
LpTSmdDu4YbdWLnNQRwfg7wDyaN34UBfCrNWqlA1D7OEycs3zzLYOqamdIHqOqGs5MFzrIZ/db/U
ZVSTaA1upqNamcXhbh5ikxBftuQrG9zwqQFXUPNZOhtQon7aN2quFWBCXgw00YIRFF7l/lP4Js3R
CcSOkCbbRGrFIiJzB0dDMXoqipqEZG68Z55X6V/UeDbbDpIhGInM+VG/5p4e+ZOTFP7prgH6sRL1
xCj2tIVxTAuJdE1CLxTpflh1A6UU5VeoLCYIDo5HRFx4kKT4i1odKjeFuAdNT54Ody4BoUa7fn8i
l982Hb27xc9CJO/8wZ5YVKoW6cSDCGX9Qm84/oNflbBESXEk6F71U9yVYMGlZTVPwps8mwNmXk4l
NI5dd+Iyddh6c0QKA5KpGiY8bsihRo1hE9vwG59ZRsTdOCoxZ+jJXxse6Slv3mh3jJuSiDzF4HB3
US0KWd5O9v22AH2bgRs5ZqCEnEEy8I9quXmv+RfR4SxOhx28EBZbHIhor9GhlsNChMQD2Ldgo23b
Kzfq1rqCTmDJrO0+3h1oxP2/fmk7YKAjrFuZQV1pig+G+RZly7xtKXLIZonCarbWYg+DquC0cFTT
Vj8wmzryZQQhg6/Kz3oPipT5d7Ver8ZfYSOpobc02F4co1+aQLeX0xFss2T2+ahbjnlXPZ0nXZKv
EOysPEHlpvrKVHo7GPNccvPAiQT+Ev9EQMS7e1BsmaVu93sHq/lPsweQhbXWn7NMrLqUAOsOGiwM
54rfEm2letW7k29npIwf/mhyY/VYGkwBl5oqXkMmibk1tBN6OCLpg5OWK7hHMRI1bF+Dx5sWLYrx
mpip7zi1OcLRwpYt15qhi/kLJHrrRSIyspWje00TnH3cs95YYPP9V4qiPra+Ztqiz2uj6lLjR3he
DVaXcvTXMRUcktZys/cn5UjucYhTF5Z9kbPHVKvMK35YsenqZyMJtNEiPIJzEsKBqKO9CyGvsxk6
hSCNRqV5UTBUPF56C6g83+sraka+lO/0eQyL5hjNTjFF4NEvbi02c8N2THxPfCqzarLwW59dn5UU
tx6cEjPT0n34+5G6iEe63m8i0zxLFyNRyFTqwnZk7u3KyxU/ms5Xn9zfZyqmLhUNjNKjQixjLE3m
sqZD7JRN9sUkVPWRoI3bLEgS7mAuHrUARTe4lChzDrajaI8RxFyCVqpB6p5WDpUpUgR/poOe54Dt
rC9hh8yRXkynv91XfIOXUQF7JmFp77+hk3jMv2ZmTYPMAsPMkQu962Q9ZNhFR+itIpBieaFzAyQH
sBXpQJ5hJ6pbn6xOaZXKCR/5xZqtXc5y2K3uDmPmQ1UTxgj2JoJodBlxW3fDcoTmTAi5orxSwmPc
wuwEV+Kduwr1iyzj3wZPcYNEZimlVTqfC2v+ykFNjbe0qJZTd7vCO3JVO7yN0/8mSqfzuxFffKtB
Pil5O+lZGst/xX5ymVQhf+pyfDOhipSzFZxUkLFtv63HjtFK+BVPFLShNvWPp8YK43mFzmYd8O9m
JbJ2juikySAzI633/c9zxivTl328CjdW9mYbNvVurfajRCx5Ec9C2m2Fgw8pQLXHZqyTrc6CxVnP
2tU7+Xv9FnNGDcZICDaDCsyXcW4ZamesX17cHRFJWq/Tv57SEyv1dLoE2jC55oVr7cK4JgWx0uIO
2vSJCAaUl7eW+YD+Al1s9hvWmfbd/SgKnevRJZiFp8n+bLL7dxy7oCfrcSETiaCiC4VxY7c/+hJ0
s9aLhw+gAxAEtQF9lsmFrk258eqNecwxK8J6mNGonvWGcREkPhOuuTL3tCbmNg996h5XNyIR3Zd7
NDRTdaTLMQmCdRdd0ykwJKYJBXL43A4dxMmNy53WKb3DD8JC8YO2NgslQWm++ncqCRidXdoNxy0C
slWfHi58x0mM7+XZjs/Gmk/GZPgguyITs1jw9yydYbqI0N1Bg2rNugaRtG4ly4/wITk3abD6MHM6
UXBps/zwoGHtpYybRyoPfccaEVLZBMaoleLQ8X56SKTiURWsEAyZ1nCCwOux0kd97Yb1Us7Xv6RJ
qHj2/LoEDoELn3fkMXDcQ8GIQGgt5zxYAXbmAEPEZbxoT98ZAKe1Bd/x6fgrl0c6tVU67FvbVqI5
RadgAizqtfdWFvb/+o6e58UzlPgmDOpHig6enNs1hGFMcYFTecji9QVaD0g9yUaR+xO+La/Ry6Gs
kdffwmMYklJ6km/G7H/TNf0LPY26mDmdJHrdRApiV1LR9LmUh1+tlMjhbVm+ng2KkrqH73O6M9Dr
xswxlTD10+3DpPDHvMuAr+Ruf7P21wN4HnL/K40GZG0Xu2vLVRQ2PleyqfSRosm89WH7sYp3eP6m
YrtEz+EPhiqQArggTI3bsu6kKf188LLaSIgGYBkRNkRXRPyl13ljuGO8aldzw9I3AMPTZOBdy3Gp
idHcQ6dTf4uTP8N3EAXmvdHfg2UbKZkKP3ONPwc6Pv90CEbl75obSVKnGeChaz4XOmNii8Vevloj
SnNtsVUTqjv0M4xqTUbjDicUA5G55gb6PLgMDgRqqLfkBMt/Fy+mbR2K29/5VDC84oVuWDaED3an
2QPkHqCo3S4lwFkXcvi3YVIPaesSWltV7N5ikMM6d10KZYRNcMv3hDSWLUbSPxirhk7ReXjg3UMw
sI+hVZBN7XmdGjgaCeA2AoTN5MpKxBxK8INny8qPQqkh5blw21VfU4yJGrOI/b47YkDb7ZWSMdub
A1EE+mBCucO57DSnRt11nfBFGaEQ4bbjLmvNwgnjiU8rtRX4nDAJ2asTzjhFxtN1ZUrTyZznEWtD
dy+uQ9DpSoXt/kZwdiWcR5yGmSIv6kgHZajv7QeX4sXKhCXWZ4JvIsanj41Z0r8E1qHddH4oVxEG
DqbGlnQUC1X5tGZaHD4xqoMwILIJfdlRs7IsxmWDvO/WnKffARMacdymoMONGJZKChWffDSwukd1
tptDoaHC5K9TPuV3UAnbzPutu3DlYZE4lsVujQi+QjgQI5Chd3WmTJE51Txl3mS8+FMJxMyf0Owy
irKKWKm/sqEyFKMD8mgmIHAcf6kaSycKfnJi36XqxKeheab0fu934VSrdPxtu9KfNvlCfT0BFeGK
H6k0KttYq31AdpTVqmePlXcl0RRDMogYIDUDq25U8me1EMiQ8ApOI0bXyR3nFS0zJ0mOK0v+qFBQ
wOnXWHtbve1K7MiRtIjwAle3utLE+MA/G/Ho0VA0oyjDvOs2NqSaDt3o7iQ46BPFR/K/pROgPEyL
KaxC3w6mzVRBvyEsiTj35ZlCPnO5F7lcBoH44XPDYf2Wours1hhRf5YAov5PR+s0/2DL5R0ekbZz
4M8aDVCeuM6nGvZl+osS2wp/qI9f7rFK/QdUUUWsewQVOZwUaK0BZm1hkMAXnVhSbSA4odzwoER1
liJNaq/FS8x6dstk0nnHFu1BFV0hzHw2oLJVfxTCVCLnJ9MomCR9ja3kUvqjm4Ba1v/puIn0dv4l
8e1hKO33s+DxlFQiUGDYAHjnOli4pGDW79HptljltBs9JQjSgUMnIHAWFLJVpb2AK3ryglbRkX7y
g+VbDvHzAA9aBKQj5SCSxBqNyGBUSUCnzVPBfpy/YrlzKJMS9TBbNhWdH+Lg7R6SdDfbRxpT7WFB
N+CwhpnDzbKbQWFgdq+oyM/l/OZkOnAql2YruFLwxd0qZg7hY+M6BgCH6j8xxJ8uaHtGsFLHA4C0
6OiItZN+53mtIvZhIXpbLfUSzzXVloTUXoULJPQtEEnFsXz4mDf1QVHcFRwKMFggs4EVhUymRS+1
nkgg8+dlsd9B4O86wy3HWghqDV586bFEHwFyFpCZPgVZG2JZh4rXPz2kNVgZx5TLD9kU33EHCX+1
bSubXF/Dx2l2P1spJ0JXJD4oa7n0zfUKw5megb6OaH3j7JbFGAP5Vco5gPPit9kIK3CZRVa6c8E2
IsI+IvLMutOj9xK2KDRtIrk3qfZYYFU9Ri8sfcWXxZ+Usx8i3VgrwbV0RV5TirHD5BCh/2KzC9xF
jt0HBFRfYowTNjmzTqVEV2j4e059n+Tf29efd70djyOI4ORtFkmWnKwGfGAcEr7W4cbIufgxasKZ
UmHXHABsLCSW3AH0Nhw8Mg3W9nQfSDlCsqGZsiLkwPGwRS2Uaqq5+zwNVcvROwmkFRvkkYhTsOEl
++Bf1HrsqINPFdc677anXINh3xmnCfPu/YRodOgAe4bqejJCodKzBGMuEJ6svVp/uRQOBoZ0tKqG
lsQj3m4fIYxXo+bC9vWiX/bVIrap0Pz4HPe/TJ4BX4pGEs/LUG4no1d8J/dIURSCDu7OuVr6q+Iq
7XUTkACJ1SBOJ5r1+kS/tXEOLh9Ns3WpQJW8xLRuz/2c6zgJNUvyTK0eOfBFatJLUSzqHmy6IDDx
kYurpcFk1U4F4lw6CcgkTIPXPo1FxP42aZe0qyG8XH8oN3N3tCOdhrDnlbeMq4b59JPR/jxjUPvO
gftfuXjDUEgVg/9R+HyzvUHmPPwJ+zvLnRspzYcZ4xVHMEzY7ms1hoNmFtHkmC9C96EbdGNc+n+l
CEVBUm8Y4oVcV10SZgw3pDDEKgvn8WSPnTcoxv7ypE27wfkExYSOh9riA1tQbUKsm9Pe4yUatj7E
GwfLgvp/Ua89UKB/efy9l6HoK9hPYMfARlo8V+NThMAPeNgySEucy0fjsc3f41dD9ugvcUpk4fuZ
GskU/rXBJUL9AHOhJt0xsgKQZ8+cniqwLMnPCsiYp/B3a5zXQwT3yBC+AkyiQmUFn89miU5+s+CI
fKsJDeYnIs13Yz/Bov61sRw4zdLVj8hwTT3tsauOLd67v2O03sO8lQ5Bs4ndS3BmesA5iOn+Gomp
Qr/IdCcznfvOfl4o1vCPOylN7lVxzK9WBFKBNiE+IRbOserdq3XQrIZ9xfh4pryuUgaKziTxTd2a
b3Ip5Prvwina/QCo+fPZZAihm+YsS6DbJ/1tndsRRgC/+B93/+9LZeTbeQp1fet9EASyhyR9IvZ9
ZUank3AxUr8CUVf1P1G1vkMEgpDEiP64IXMNMWIpC54nq8+QYiYL/2Esazi3izv8WqpEnfF9+LF0
ahKiLX1KY44Ci0DbxAgxS+RSLPm1Xnj665KD3pHc/VpvfU25SPy4Yh2bx/Nyph6jEZ75COb8ybNR
zcGJtzyzGcd8UxY8rEx/mnrhU6TIR9dlNo+J+02gBGtGXeZac4/FsxSbKrcaBCgCvM3BNTlJywOl
1d6GK2/R3vt0s7aB1U5EjDqOC4/xhAO3nEuDSTGZhV/RG9QlcFfo1z81u7+punBbFpDkjm6JwM+C
ZTb2tkjOr68bnyp6t2xy+HBrQ+NQUTxw2gCjhA/+8dBIQT4+6QTLRDf4ppa5hspYw/Oq/JjhnCR6
hkVsfo97HVkyIJ8ZmnH2tF0zwK46edwI37+oD9J4XzifB+tuoHBLJ1Axwx4GNrsaT3qAPonvfK5U
PMoqDUVFQ2jFBRISW1HVk3pDcldZlfo4ahUOW+FOJLk2fvT31UWZyZfTkb4NsRYSx4gk1s9atI2R
OtU1ieXO7f4qYeVBzmMqHgbmOeHR+cZHxkhq43YHn0TntiE7eJNn4zeFg7plxAATcK7OAtQinb+0
R9ppi4bAhfCt/fwrWZNE/ItuMd8VNPCRVATXYpHR2skWGQq7jFv8bzECStG2ZVqEDX4FIpEP/lPx
+A/uk13cWtkHXIcK9cWio0CGfP1BgbuVeYLXUS/tFdsfQD2ErHA9Bj1YHLnV0vEH2zjJ16dyJ7F8
vBmI6C6+YBCta4CoGEG+CPb3iT9dJowFT8YKMj9pCmvaMJAWAIj/VoNOQ7qZZLIVcYixzRbg8Tok
96M6PiF2ai+aH0cs3nNLqXYqBD6rTOMTenYV6lh0SPF0dS6pYTzuuaCESfqbZOu8/ER4wLsK3Vpy
OwA9YuMpDpA3/QI+mQ2Xdaso2q2M4FVSXX5B1iob+GWeBVaDUqAriMvRrVINNVkLC+saApHodLDQ
Pfbou65aegjftArg8tzvww+tCsv5BNVFlYR6P5BVzT16TPeMATySs9QUI1wfsszdDtsqFHme72tm
LT24u+50uPzecYYUqt6bIGKSs6HGMofhGUmLhkgku0VaVLdzPFxrSea/oSbx2NCLlkejc8J9ontm
J9douv4lPcIf6rZalqmAcQlek0JqESgNM2ZdNBkqo+uZQWCpeSt08xFhXQW6fMqdQeHl1lWbNTtQ
EW36Hap3oVtVUpPmnmgghebCoQkgcr9TWh7MlhS2w1f4aovAJivCE97w2Ub4PvM/+6zHDK5SpXWc
JpWUSocDhI2fl4hPbBgTKedTHLJFMxo+yoD3zIUjTJu4OX9PfcQKV3sCD8A042i4LB+ne4//X7m8
y63yosbpmPaaPT/wZNJygMsoStnL9pzLxAH9bBGOYEyOJHKYcfBGDSwlF/KtsElzyDMkq9jQ5mse
/pO1Vp+95MZjMvpAhqFaRMw+tY0drV1xXfiP7nTFBcEuGRgQ7OMa7jX9y63sisS6khalnluLv2NL
xjeM8cSmgOudNvN5rHo1wzN/RKAIjfVjHzhKXvsGY6WS/NJy3Lv2ZkXeK7J270BHIIogu/UfAmwo
H7zUMDOvCJyoHw4NKioYh8UYse+eAz0CsWqzT304o1pzrLEWUGD2JCWlDsw5sL3R1va/T1bYmBWJ
5mA3ioJYlT7ft4qPSRRJ2HAt88gsSKrdiUD890/6WrRekNzdRHmHv9HlBRy5BPWDfczgy5Gx7kxD
WyMwJ/o2LVnSrAWY69vx2hRdpBg116/135lgOhpazXi59IaTwcP+tIE82KncKan5n+elaY4gIk1u
kRJbQSayeiUEHKkJsrTkFrhl8VsYcdoaD11l9uL38f9B+bOliuxHFtuA+WBsQjMSBu5mMIg3nEGm
L8U2C9LsycxLZKGoLFAM0j7J0ugNQ4DSRYTK7ociQwVloNIGqJkgEIhJ02FmxcZGoxQdoBV1AfrA
P4F8JkUFJU4iK2pCHTVlfdj4f6FE6PhGxQRbJLCIoVwoSK3J4/pUPv1OxoeSHjgwn7zjv6wGYTUJ
BpOM23Zro6/iqyi17pBN4Rmn0T2hze9mDgcnu3xRwq/GFkd3Os1t1noiLZZjmNVTxxCTPjQsZw5e
mPWvphxsD+nz9ZmRRAanTT+7G8imE2yXawfCPfRjJlf3mSP0Y91iCiLXsQQK0YcyTQm8RSobF0fs
+2OMkB12vPZAXyPOCHu06Jh0QsvUYQ2lbCOYCR/JYmbrn1t9E/5PcnMjsXRh+2Qb2C7xOm9vG4FZ
KTzT+xKDsX66sTqqxYk+onjjvyW0i260veSUzl5a+y5K0gexIdTf9apoOXkTo6COrIQLsqdywiod
WyXA5GD5GBzP+r31mt02Mnr5CbNhx34JJXrESVLpcHOGJvpKb7exaudptraP5N/FRzUSZCxBncu/
wvFbL+Yr/Nh12++lqkHoam7RRd09T5BhyYhwk7rgrOM90HHc8sj4CSbD72xtOtKWWTt+hScriAa9
bcqz/K8SGtzsmziSvjB5REjIxyrRE1f7kzT/2WsmnAo5aQ8BcAFQ2gfWDxgd2pQH0pm5yY9hZgsk
w8YmiXekxAPjJXrPR7CZVpvm2ZSiclkyo7vQ/9J6G8pxXf6xVx97WeIj4bIujGiXZBYb5kKxNODK
UYsLx6dUpT1nOJD13uPGyyw1ty5l15VySTxZCuC9Uf3ztMe+9ukhSGdkSMST5pKFjs5mrLveXGKK
OBUp4OeGD3+Uo3uP+VIdc83yyEPjc9jDAwXwPRzN7JjFm/Al5pqMn+pt0zNR4NQr1RnbTwDFt0yL
9jIKLkSSrOu7DKZw8qo23cUs+NuNHdDEQOc837QC9J39ryHQiqbl4E+QSZ28FwjDy46u+UIwLlsC
FeV4yblpBaMDr8VdGgmRROqRe0yPzRY6X3raswtiiHvWB4f37oxlPw5YZZucIw53hqltiKjaUxi5
0nlFjiYkJ1y+1PmHgd8/Kg3GdmJNn1Tk7kUA/WZYtY+e8pgyqEEYyLSyfIKzbVquKuXWnc5C602j
7kty3IjaAoP1tnPzbnbcf0AYaMHGEs3jsX/VjZC2BpujtvGBnV4+60hJsMq1DDu0q9Cunt/EN3AP
qvLbUIgi2rwLl/QakqpXLto0WVA4YMU9T/qhv67aOR/w5APAPKRvFxZjbK8X77l9PvZFfi3alfJj
IRtDsvvv/y1A2lVCEM3c0Az5dMlmsq+WxrwCfH/jH48yCmn4nyFsLEGUSltSGUVTI8ITqFPFKtJR
A7a0a25isoMPrufsj0NC1o7dzrBuNhaFX4Ejg9cg56zNsy3wYHeiBSEcWAYNWv1hFgFjViLNeU0y
mHRsPi5nZ29FtqK+b1iD73Rt3xC6StCfd1+biu7FoSPyViXKqHyNGdo8JzXwlBpWsuFlOXJ+NYul
ZXlySCNmWE5dQUOfXEmryortMD89OJhhxj53xUYVIqH9mAIHnXadUVftlZnP5oy7FMy0QZQqxL9k
bI9CqXUULtsyiUBE1QUWcM34NcXHa1QqhXFNhW/+YKt/uHvKJAMbTDy1QulhRhOgIip2cY9JUI0z
N0aCht/R011i3/oxE+VWVcSXF8w1fyjRHHRefbFYNNMurDL9UZj6+lqNO8iJAfakoOeHRCpgbiXR
tcglWr4l3+JthcIhN1EfFnf1ObNnjMF8DS0UE/jQQWdOIeaK+4XIr8++vwFtkEEd7UgZ6L2E9oOU
baxkhXFlqkXGo3Vh7MvkweUn7QUaYX4YOfgNXNKY8TWGn70vALSvpdIVjud9cckKUMZP1/BgY5Kk
gZsh0M5yAvzU/B1H1lohOnhbWJdyv0k6AcJ+cip1TJ9nbaSPwsdjckjehYlHv5Iot16GIkdBjjRc
5Cc81hlDD0IpCbrxW1Q0Y11pFH1VuyvrDi1R1wDOCE+nadE6coZ1AK4keUyxOrow+cXmoSip/8Dt
z9H9LpWLhpTzCzs9gvrllIfrVHeeQrYpjY0lA7E9hvsefXSXkzB0RYjHFbkdvhiN2okVq0rRFtHd
EfhbFFR2l32cRSaMhxA555Dh8rFSl28zsYvDGZa5GUw9Zf9peiHkcBzmMv+Ru9Q8RQ0yRFoVfH+S
AJ/tjNVhFf22jILmxFc066IVexmXI9YKHNALot2YGgKDZU4WuZm+SpMZMrUeq4vefSYPhG60mzPP
Uv2lzPL5m2eLKLK0gKATRtw6sejYyjqeJ2TnSQp9eboWI4NLsSr9mLFxWxPObUurooHI8j249ZQY
IShUG7LBMr2FX8kzug6t+XDuNlF9crY2Z8zTFl5Anbjzp35hoGJH9H5bQXJv5Tw3shtoCyndGeWz
64kDhUMagMZl/w/U7J2vhA+eohuSYyR4BCvLTzv5VNE0d9lfitR+Rhp8hPd43qZG0Og4FTzySpod
HcpWTRbW4qavZqyR8wTTNYiZ5emcKIjR1+9mmM7t2EpsVo5+G0hvftX4F72/9HvGQbvFR8LKCHdo
R2GOqUWXTz43LIvx/XlMDz1IyRYxKDKSytMOYZiyzQBrQ8egJIs2qn8mVtO6dtyqlDaUXUnalsIw
lL6nic9AH+1qV6Euzjd8dvMPdCzLN/9XYRXXNq9YsNBHwVEXg5oqrK8bRAHjNuZg5c5bN28FsufC
hyQmEupLR7HET2kFwc4sd+2f+Ogs1HRIV3c62PwUgFWAPc5zk38w+bN6zglmgPTpPOiFQWHjiyU3
gUVuVrozXs1jl/Ix6jIxgsfn75I4OXEMIiSwOOxtN/SQWvKfsqvH5bGB3trF3AIFGNdEahMWydWQ
7L33XC4Vv6OqWDvkmf4xBJNvABzng1sNgl1/v011NBG7D7Igkbf4upGBXSqjygvMQV5mG6xtnaHn
mY0wbmmvLsvr+EY3cWEKtj0GOkFtHAR7gocdHquTQBiK8oT1fX1QZ/Pssb01OdS21hCXlJ7q/2IR
vW80ZKL31d9h6S7UPPV/dMAdxi1a/Imq0bnmkf7J8a2yzsg+Fl0URT2VD73plXQaDQRGkGgXdQvb
9pZrdEn6MS4nrJ9E0/NRY7ge3GkzNbdKUeP89MOpQiolg9lcCOlvtHxy95U3XZyGeQCN5jt5W+JV
Biw3KyRtMK+Ugxr1bNNcaFf60AUT9Eic43k5WTZVM07X9A5IStCLlOdfQ0gvDljNG8P4KtyeEMMy
AA34FAPI7/v7o4eqpr6e9CKaHNLZa+kcZ3+SeU2t7fInIgIrMP7Tca5uJHr/eYE5/JF9JnGOclYF
+8hbyqNukURwKFbSdv83ety3b9cW9RmcxfmC59ZQeS+s/34+XO01TWF//n3ui4XldIjZhKOivi7/
O3ObdKOsv8m65CPkQ9/VksayRoHwzMPiwc9QmICz6o0wXwgUKDyL6B+jH9pI+0E5g1tEwThBbeDE
vdljbXi8ToL3ebVM1naVr6eK66TNT8g+bkWTA/I4fLC8pXEHBFSk6VayrcZv7i6HdnSc43Dt3ixN
h1jwo2RnaFpNESL++CWQpT9yn2klXUp7hPxZvCQyNIkMpZpk86Tw+A+TWk7iT1PvazE4Grz0fdXl
mrPiqzAgLYxRNqlrQJ2NjLyIf50uzdBaE0Q3E6VbxFkPIYnu+CEkSq2SeP2HyQ5nNo5g2a0+c//C
ko0n7zMisSrty7hkc2o7/HDrDemHYVfITr34lWt26lKHsZMg9jvfZo5pLL/aOpHg+GIz5KhTNLmv
kjOETt7o1fNIg/X+3y1JEuiDJ2pXYmFHTZhC6xd4ZhGV9YtD+EUuXEGT7EAeCWDjb8gZk4T3eMp5
u0D9Cdk+nP8TLygBswxyDjpWodSdajAC5YiX3p1FgZHifzRw7NktWx6qWT3l7yPklVz8wdRr8yap
S9G9vVsFO6AnbtoajRyCmcjX/JA4Yotl25puoGGy2FkTq0rSne0Qx6VDPCWnOcMnKDD5wfbJc/j8
irCy5KVqcAn/uUAwxPVXlTnkmdEI/q2OgaIukifzplGcMZbO2YruLipd1viyCVCh8/G3pfb9t5Y8
7vgTr5zGsmr6os/FEWk59+NkgSvQRfJrB1+Bny8rBwX9SaoWmTdwODtYWKLKfU52foMTTq/tBG5t
xxbmMUadpVeI+E9a4EflB0Z3FDTwyy1YdvvW8T0u4kvt9uEWWJ+OkhrCHTdNn3uKVIrst57/nA8z
rb+vBZkjL72WQTPnhRm85qO4xHTIr8lzGE5I1W9sMhJiUgjzHttv4Zfbz2bTIWmbngz9sTQTPh+4
ZLu8c+pxc1Ar8o2GDMXxBK7bkm1sdeZMy3sJmbWxXiAwFF2tExQabyg8jSuT7LKoTJwqly+4yJRR
vLFAwSeNYaoZwLQCG2RY5CDAqAQNKbunf3etDbQ8ymkYqRyO595CLDPlGW/cItYtXrQlwwlWXlId
nbyLTKMnU/tZDJW6mTaa4e8KxGZseSjKKvDMLV+hq2oNliX2E6T14VZ5W1bRb2sGMlnIVgwntlBZ
wJ/ybqRFvMoOcZkdDzrjouLhw48Ow2GWTVdaNiWVyK1d4TzZJuJ0A51OyDjjpom70GJEiWeXhVuM
lCaqe9MvA8k95zZNAX81tX8hpEA3gwkOCtuD/pKwmM+Ha4AtvNGi+TItvK+pvraUYAQQzgQX+NJ/
CQlSt9bSahTr+8yo4+WEuQURRAY7uPDiAfBC2qeYBMBrmC92p6EIOp/lwmwhdZa6eSIpgxuGVAJk
SdumE0pq1q/L73TFXqWAiY3qdGcUS/mBH/WfTxtU2J+izXvCTD7vkhCaXTEilMA54yieUdekYSjr
H5/0HrbKzkdnae1BBjAMPsW68szjg8S7XthLzwVYShf8l/mrhboqoyYVtpkPD/37IZ86qWTzpf/6
WSSuZW3eTATIlDgw4vTuFItzjegfeFub4+bil4Jfl/mHXiWSjHu/gUjJo43gnNfOSSO/rk/793bn
h2x7rI5JWrOgaT3X/hvbmDDiP63hpnnDoiuGhhFUQ6uupZLCw+SlIuZnKPynOHLRw/d1xKpOcIqr
6RJX6uslyI1wQUj0Ht9RxHgVskC8Q1mP6J8yfVbeYncvuL42JpPadO/VQN700E+OyGeYQlXqOZLb
MogkkqoZL8VT2rcBILvhiHyITogFGXoHtacXlFtDUvQP+hfSiwXjT7ls/xRZ5xJHdOEA6R93CBrQ
/Aobc8l0+vdm76cWRdIE3vYEOJ9SqEJP7yPcdnI08w1xnYqsJRB+yIcYhmpRXz2rpcWmAxhlnoIy
a8HK1LjpLI/SneJRFO/Nsyn3Oo/Q8bjqDrmiJCyx1TKqeL0kgYyCL9mD98JLzjW1e2o8/c3Qe4Yf
yhdmtWQ/l1xgKvOos2AO1q5jTolQlYkK3/6ith5KcO2dxJaOHkrF9E5lwXJufloRuxhNbfz1EmuV
K7s6O4iWM37Y1d48Ja0A087rGoK4Ur4/B7Y8xjGHirJ4kA4btR378Rt3CcYNkW32f47TwPVUCOzN
tAvKiMRNfPVcVGC+F1w4gSPzL10gFXXTTA3asiLmF8CcP/kvPNNWHrtFYkkv4Cbq2juGBZua+5p6
XiWc1D1DH9bASQX4JYL6mQDK52agNN7FZTo/aazSSNNtRR5Ouv4Nma4RFKujyScAuGiNLc5NhC75
VIJFTxBgsJJvUT33eH1s5gKF1S6iM/gIyG5uzD8m+sfPP5i9DX8P0agxJCZ1XTSHBMfpkeJWDUTU
BeLie3eDwjXNG8HFuz5ivs8VhoEeMe2qdWdpW1psyoYwQ9zVSjopBSXWlAlzajaqgiy8CtnndhbI
aorV9thh6/jaz0ag7aq2QSaRJRecSzj54q+XTvlRqlvlLhEkf4XxHYgYHTtgacx+jsMUuSDANxtd
tAKanVO7mKPa2K6WeczGAGCcV5mpn8MDV/AaCW5LW6SXt9zyFURMjXaUnhKDfveOz0XnxHb2ZgRj
FsXeAoBSqjnC3nCe1V73r4J/0HZWqwOcgEJFJPf+EEe6jVc00A5gvj2vbpIciH9gB6uyGisXxF/1
Q1ILzVUdd1ytNEYCeypeGVCI/ELlTe26KKQWVtqrNJM6vkzgvWqiJEsIwn+DPCoMiVpEKKkz1Ysk
EZYiVyDZPsO7wFym1lql3r6HcXCBJrTKNKGZMXvQ135sIWXbhcAw5hHBHAoF3vtzODrgcXQPM2rP
WZObWfwJAS++2S2kv9/ihHSUKFQlsufI7Rah89hVEzBJTHlzjS4ikYQlxjfz6GUQ8Q0tBaP+iVQ8
BRgkshxEe3pgbMwxSKlsVJS3hZZ4jjqpAOGBu/iEZsqmy3arUmgHhAHbfkD3zDnwPEw/pZw1pDZH
swNBasj3IangHQcgRY4iizagpLGI+HFMUcQWATwSvc1g8cLXa17ltKLgXVUq0bP+DFD5dzDTAIkV
UK9mt6TfmoiQvsn4Hq9xA41dxhXV7FldiEPDy/hKolYyp8lp9ZkcCOdqCBZy1W5EJVxtgTL1S8rX
MmeRaqr4OJsizvPaC7T6iuYWQOiltyDkFT1Dw9IoKnsaIVKpuRGGxvCg+cfXR2HDAJTdV7dpednv
QB5HWrC8RKMNQYEtLGB3OxfSVNi946oaWc0P5SAM4TClma/kacPItCTDf+PnF8UA+lk0diy0NGMF
Nr75lcyy3pewwk2bJlzhZ+U8Ehq02idAL0lYZKyDn5+0jWnttNg9LU49CBhWtlmSQ9s0YQKCveBL
Igj+ZqIIpxKypZpCZOdvk3EgkJGsuuEEfhMuw28QJYBYW5b1/HujHRWK1t5LTjKVouQwWGbM34cH
oY4pO6riNDLlHmRfS0WN1tQPMcAF3beYYTQFayugVwCCKrzPbmh7xqfXYpulgOfQArgfJq7+6DzJ
TE3aak9Ioz01WOChC37I0k7bQUj34QvbcUJ5mkjhCvjkYzNLsV9APJpQjulCzj5GlHOXnomBziTT
w06A7bqVs9gwmCPcrtnFzsOJOqSSrIvsfowWKhHwL7Y6UvJCvWUjsiGSS35V0ioRZQ3m21pZCuTv
FEGXroDbz2RslY3xOmTK4aHyFmti7Hx1BEqDOellAFLCQu2wfKVl76PnpaAe41McqSLHRjtKZZ4F
x2hUhub1QRntKl5HckFzO7pkmoqVrav3xYJ/qhpBlU0H2lKXH5BDjLoZ941QZv6qMzTJRaWYxYuB
44IURK8q+x3RjiCfQt4El9puz0wdYrxipqe7u0VvIASMOOWt6pkAmUYdPEv8r+eUK0fxjMx7Go7W
mCZOIu5mHnhk+Kv5hj0kl96Ev1KPwowGOh2VNZso8e2MGN7wbdRWCsksPaQC0iNon3PaBHjmqGpX
/c4xHRdgRRefwae/FdwSfsp+s1FStJA/76AkJAUKeqfxz4AVHDF/e4i38sOD8vqbFtsgv3KDcLdv
KkEEzAAd3D1FKp3XUWYUe6dHBaJvP2v0VpNA3eg2RskWkqefQkGaPWhLqfIoYe2x8QwFq+EUP0oi
JklcDbO0GmrLYneB+fnoY5I0EZIJBrDuzOLqis9zH5GhThxzHR4jnBWEVqlrixdt5v1G68CpQjJa
3CLIa63dkD+6hTYEEvH4ZXeibXlh9OCVaZ1ydssbwshfENzu9/K95lRve3+WPtq2F2dSFp/xMwlS
ilPdlhiZlKO+siVDz3+l//LZvU3oyJU4ZTg2cDS1pN01ia5qvkOeXpAQtQLMTzhXYXHCsiMDDKYN
d7TDr9CigPt2dFzt57Dn3tNLErsCKtvTx7lRvZOC3bESeR2NpsTRSYQkBDz8bX0RjYf/8RRJoIh2
ErWFxZpnc7/bgZlz7kZQhpKJvHH7hF8txyRFUXiL/AUp+/GYge6+aJ01Ao9H7ZBwaqAR0rvnG74O
P4XNylpI3lI/rsUgphBn6oGFNXwyBlcw3g4vxiRjvYZExooHiQMSAFPjRWlcKZDW5SGliLukmb/R
DzOvZO2TXkIDwuXdf8AkPW5732g/Xz8jO5RiFkAj30MhQZFWLUsAyYQHUh751MBpMNIlxtcdIoV+
p+r6m0tuTaXXcOKp74k8bD4OZBudeh83ilRfP5nJPSIUH7j8nv+K2YtvZORl5LdeZ+lHE2Mz+RWN
dpXXm73aVy3ATP1tQs6cIKhxQxPC1q8R0VfhsL+mLF079EV8/jyueZ9nFtY/wz7aHHi9ARrnJxj7
wi5AzmfWKTuLfuq4U7EedQXe3QoS///TI01p6VQlCiuEd53ic2+Fjspr76FoxpzIWhopzjHtpBLy
qKyRVJ5krpWWn1tS4L3QUP4ZD6VwW7AQMJEQ/BdWAbBw+BjLSozjGRHSSIlCbCh5rYN3MT06Ij5M
kB/IUW5uRTficenoKjxmtHUxMmYNos8jGJxB37/yaTvwAmyTCEsuHiIsZWeAqPsDjYq8P165BZvZ
L5eHXnxzIDBuzz5UYwrZfBlzg6f3KGg3yashNMx15kd1fgzZ9J4Fyj2BBnP7TPg4OqejrOpy6t4L
yFgaf3Tmr/aMATmz2Mf8NH5KB4aqoSN89Bvg5KjUG0C++VPKnmpvpExgswnKTgImbmNXW/AajZpC
Nxtr7d1o79nyXY9Gm7H3Kc8RPU2AgunFo2l4YQ0ACTxZDUriizvK/6a8ZH2yP+m2tDhc6Yvqfas6
DfhfqDe59pw3Q5I5HqD58t9Ohb3/M2/psqPjZGhuln6dAL6tHZSxUdx+L69K9nnMfAoO2prmH3VQ
kRJVEX+Be95vW5valPkSMqeF6Mnozn1GVsWVbyoOY4x2Ky8DVV1o+RlWtN4AAC/t2t3PyhGrHehU
bWr/KP55LS83UnzdC/PRfiQQOH0lD9+5JfJilSPxb69Pz68dlxFei8o4FAy+dMRnHzhc0dFIWKf8
c5fJ9nAXdq3wA+avONTk8/4lLn4MQ2P9UHNTIRSk/OmAeAYKu86QVRUrNKflBozmGeJuKcO7YNvu
2CRKslavyGrapexS1A0CQ8cYqp8Cu3wBS4CRuyxh3+/BOp3N05SLdOKEnMXhR/ElStaFwpA+JWrh
MvVEOBg0ODVJ8Rbqzp6FzP6zn2hVWnqwhjVufDs0B19Livazzed+V438+MdvKOOLk/S4AFj6mxTr
G01YTAxFl1QrIyNQMShImNDJW3LPnaHglxhtF5aqQrt7vmShxfnCQrkZbTNPI8gsDFJaNQhLVyCG
ULQZTiUSiJMmF8lPrR34CdDqr4Frr1gVhn3FemNstVnXlPu9wqIaJm+Ema/TfmHAVi6v8wn3t9QB
k8ssPBbmh/K4CiI6p0Tb3mmy6rjYFSeF9COeXDAMG/cSEjImy2PuoO5nQV4pkaDZXJeOwkkYbv26
Csn47XIAh+m5R+aCrOSr+nQVkLf7H3/MAYvVgll3uN4Vz27txfIWn2PP0/RmS30/bLLCFN84/KeT
iQK5rWgUEy24knlpQK1Y9e2jU5B3tgZl6wS+PMZXHwjBxHOWul/Ff8/EmBW5lI/HP4VehptzytjF
czQQsVxbS7s9W3CNmLxSRUsvmrbgqmnL/Z/3Fyy4yg9HUfwFDSXXmH3lx+UJfGWOJUUhNFhIDSkb
rzAJzXJ7MswaRvpCpc8qPsDbs+cCFR5JDHavMl1WuC1awrbFxIvWy6Q5dlZmy4Fto+BCXIe70U8Y
yMcA3TT5tg+HZFW/dGetjlCGUUSrzLGW5blxTl9EY7DJRMCws7KB1HOxlWXRbM2WdnF8L8tbwRf0
spq5B+faHu+hJsU/XudDK77ZlbRRoTkrWyYK10PjkLFX7nQ6MorrKLXCWNZWWabyJSmhKXhs960v
rfxA1Qnrf1/Og6V2ZLqif6UaiXLGcAtgPbcYwmIK4HAWQXLTaSyBoZ3vX7GU0IeiiA4IgZwHeFrG
IUx2yF+SUEC51GIGEmeiLfkWvVS7WwiG/h8+ej3NlOB50u+o9WGdWTd1IA3vAvXCht6aN2WzNE9b
QbdAXBS5NFh9bnvs2XJ+PGoXRL0F13/jRx74uGja8cHu9QmwX1BZxpALmqqm75XJl2rcRmoXGUez
qGJaOvqUpUFrGmq+PFmDf6QI7kS9ZDyMx6LE11vztAFHzCN0lGwzNqLrFyycZrky4E9B/OECqkwW
Yw4I3KSm67bHEGTi6r/pLUOwTglAvrr5ipJzrGxo44wyri6IqL8sXVbTCR1bTG22ezM5Yo2+uhjA
+XLxgXoC1FI+ySahqjSap//iVMBkOzstQ3ikAgKU3xsUXVe8jg4lUD2Q3LIHh+yNtO0onu3YbB8w
4h6vfIYYPs732zszH73YDkt+r7j6JmZ3nxdAliFDEez5EVuwyVL6dP9UR5YVtEpdt/9wwNIMIMyT
R+9okMrpD/9d9cnKlq3jgUL/fbvCoDeEW2s1/a6h70BGhOHonBGIhnwxtROt39Ty+fbnWyguH45/
RopeJsnYtBeOpEDBKBMnCBM0DKPfzOuWR2oAb3ovVrz3Ys5NV5uQWS/IuM1PAlbSbMvRaKEHfs99
eLCi8QMvuzs08+uxTpew3m00pfApzvr40sKV3XIYyDuwUi83aV+qCjzhpS9uLBWx6+BXMhf7AGg3
AcKHtfRuE3N4BFlFPR+YzlgSMJs0Y8Vlfg7D44jcA1U020eKc3+oT7HC8ltoORPu0BCFuDDCfYQw
CwzIUYxUZX1kmFgNyvfkG5Vy7ORO0dEFzLaIQ2AZKhBAKYmCKRg4QtLqlE+cZurtiVd9YbMHksLr
ikA7CGSwpoQXes+p0kMIDfvKmZGEyLAI1E2JNed0yIZVIyds3NKAIa66lp0stzBRvl9EYNu+PP8i
Rk+c9H1KPp/z9AXY165pTXgESLklbYoBZ+FHj3O76JPD5RnP2noaPiMw5p7hPJm0s3stTsxP2IR2
WqDhhnfYPn5alzUmzmxuAdSELZoAk6i2FPxKEgp+9psWcnKYFBMFZUpVCv0ZwtVpG7HZHUzNxA98
UWO6FbgK6m0bUo/UEanP0NXJLelJmY6qpLFbetdBkQEhBjHsFqvzcS/sXAr7d9XeJaEJkRdlWdbm
1eTzryFQIpQOdFjfIq6TLkNnkPFlW+QXRpxjGEfDcsdz4kzWMAkXwrY+V/cR3qRRf+wyGKC9j3Ds
IM1MokiRHqSP0oSJ5KsR+Sf5KgtwstVmE9TxCNxAotTZ5wAnG11qbVERDvaniIEWfbD7ri1cuaQv
7UcDuXgaurY7FyRfFTJBieEHQHzE5RAq1QtBUYWe8hRzudqH/zXR4xf5cBxbkTx82KsGmKz4KlBA
mulKDcFhpMBXcFQ0AObtMid+WnyP3wnKNjJBlOgxFyiYkWN11G79Z17VMxkK+mQEp0a52sWf3aH+
gKdEPKo4wUgYmOPiZfDOdhaBWDgWYDU3/lQ8CiBdCz5JiJ8H69eqqiCPnG0fQy2RO8jJcY8Le1fe
PM2qXYpvYchaWZPoQT3ngFHScXk6De0TGWNRrJkMkajJtKcX5uvMmxQEzqbbkrJPsFMSM/+wdTtK
fnvZN4MO2mfVFAEYnVD1F88TBvfFItqufYpAl6TW3Mr45YMsDsKq08AaAhDU8g3oA03UgNkTUDBO
9WF19wK3CenZdjm6HiFD5hTGvBREFqd3pDr25E5m+aedNFSRPrm9MErr/wW6hu8uCbvFi5RjurgR
72Tl6YwvmdQMWipFOrLF9g+K5ZMNqq1v1oFV3HWtX2hZ5QzPqkBZYpxc6d8MIVBsZrBhLWfhoowe
uJMenV9oDidVg7rEpVxCtamQ7/8gIENMy00y022lUMi1IYjVO/8KQWHiE7LMnt3ZwPjUqdrapD+i
RHlSSgcDmMxFZynBNDF1k5vMdyMCa1LyU88DRW6Y7fX+w0bZ2yT2m5Uitr3MpbPNUjul6gTfBCX3
0wPXtDjx0VIdeilqYo/J2fWtMTufNBtzNHA7AUh63GW6K8AplXz/59Di++xlgkI2IaDW1/srnrKr
2rXQyMiIeDLmoVsQb2fjMSIDDDq0GPuVlygG2MMOv7W/yLLB+cxlbbQWVi8avpLdMM/QqJCilrBQ
VKtTs2NfZC0WgvwyVdP3sFWcyTz36/SJ03A6EFrJGR6SqX27LvXsrKY3gQ/Tu92m3G95AU2T2Y9l
z7INbZDXrKdJXkgpkDyF+QCucroU7FvGji7ysLrgDpwPpoiMhectSJxmGQUNFABO4vdMnclC/YdW
z9R8iKzSpp1iRIDAUoz4zTeytNRgLxXPJDrDe7JhVjg2SnPUTtfKLpdyBby+7stNx3axCJaK5Bc3
+I7VQr82qfPnABLLYUqIHuhLwqhLQOAxm6/naMaIBvF7sP2ZkxObfFs8BjOMOKzysVhMx/gOTPc7
SCmb7ayG7Ofb8o9maXuV/T7r0mLzQ2Fw68PZTw8EmH9OQy1JTTweQuEc9+9blKxUgZjZkRpbmktQ
ETcbmz2/+BMLA4PIh8mIzxqZfRW3iohTVInd/rs0fvFe5MzRjnETIB2sxn/MR/HP7uSaVLofvch2
8gFgy33H0rqAvHiO8yZT9+8f9F1pxzYXbZP0leik+BuhnK5EiXiBr8SMmadVbMJbJLudCg0zZlDZ
xKFaMUe4HJg6SUA3wA/3kwpOqo0v2B0eY/2Y4d40aiPmgmxcmhpf6N2NkIsgjoavj8E6gbhSDwg1
HB1rNs/tRCuRTg9CRoeQQvH53T7GMnEBjhiLSF3hXzhfL5HlkCwjWnOJsYujP4XVZ3KSxML+fiWx
6OUj+caB552KMbPDYHupaDfT1IhfkHadLAh9NipIloCnnrOM76S1Nu9LGhJUqh+P/uRm77byrxIa
lzil+fs2g0BZbp/Wkt44tWa+CUjgv52+lbrtl9zW9ObbwyEoJSkhaXem1JCwE70ZHLZPGbotTwYa
E6FkmIatP9JD7D0jkP+bZUpOJKqIilN7aJJYaWNBe8VjWbT8lWVgon/QYmbAgl9awLIAwGWFcP0q
mjLF3D7hrccQkOp1F6YXgHI183S1SZDgFtZ24ZItggHbLQWKtxnITVKlhnotgmz+AjXoLudQcETw
ECwHjh2fUGPY4xDT0D/exKU0WXgc+TgjJ74IcaW6GCHdLSFWceMVvkhV8ST0sznFoyTmQF3ypMxH
cVPFjxNPUn5OpWRE8g9agVComCS8jzDxIBRQTte7ZDHH+Ahl6SL2Zb4nOkuFjgmiDad7Ksf8g3nd
9VodUp5O6Z6IEkIgqafcAsdzei+4kTG1904+AGPzm86sAliUyBNGZqC19v91PsXAPLJ+d9lDV+yk
qp4XPSbGuaV4VVGdMvS0jajp2XarI5GGwrO//zV47yY8G/BlJKI0KL/i3OFmQ5RFnlwvmAUMYSP+
uOr8vW/k4JjADd7iyQIMQK5EKsVNzm/eM0UVPFlqX/mrhrl3Mxb+pG+MRaPGkrCx4QfHT1LJoinH
5c6idjnOrqlWumgM9F95qeJKJZytJIMUDOQwb7R30rguFZ6Q/RVr/fXwu9YZMoh8ZJhwJpFxBMRT
WNERHi+MVH33u3Wieka9l2efQ2mMmpYRu9+MFuFOVvSxzS1LEKvpJASTvXhNmFRRlI6UO/n09QmC
0b/bM8Dpz8DHiKvngy7nPwe7i7colv3vbfsKrMzf78JrLo0N4kh3WSahL0DPCo1OX2/S5wxcMSVp
L+Hfz8vniqP++MFflyQjPuRZ3r5FiUlfYWC+Dmn9eIWGY7KG3K3vq/x63ek017ScfsbYBCs73Erk
huvDZSRhPScPfAYQX4tAKptvzRAoxb5TSv/M0sGV339wlbTMrbU6jTUOKBlDpcoKkNdFdKMhInjy
DUVkgfteTRiP0U5k5yLJlu3vlyi07IUq5J3ELltYkhSOc+ptUrwAkMwRtQ26DPPF6Gx1LcBH5LeF
SRK5fERUW1zn5214VIs24mD+HqZux6kSkvQkXn1vyp7Rr+gh/sZzpTuwgNZWq+gaKEdPw3hwVkm/
EaiHH3cX2Ls8UpGEtojzIyqAPHZWrGDpAycZ+nHpO+xs70sRfLB26V1yzVgRwNzNGTLaS/mgNtOR
GFPhPyiFcQyFRJaVeMOTv5oQS4/aEXp89Gxezg6KBB71TEOZyO4ddq34cy4mempknCPBIPbHnPwd
bEXZEKrp5thJxS+2SFp5uWJtX70U9GCtZc00aFUv6PndgzJ/PLkWrxqz3Km1Yym7X74YJuR1mH15
7dowY93ae+S+fCH7wytzshIMCjhqrQZ6EIKc55XleNYXuYdlHhMAMzJK9a3/erKaoLD2bgwR8u5/
qytqqd+dIh/PMaOlCsMNXpRf0svFA0P8dj2S15JDAfugt+DXJOIe4xhpOLQrDuCGFQDyfhdRp/A9
N6cziUvAQxf/5vRo3uXc+BZ32a2am0wrBGX/eMAqhGvH8xx3dymt++nTrEU036kd/cUJMoOmoIzZ
DpmwKIlm141rLeOJqtQHya2QedWAeXNDoy+8tm10lPLyKrWmxuy194BhSV/i0ixMQmHebK0gmaOG
lbx0PkZEdQPeaHFaJj8y00duamshv8BSYh4w0KCtWI6inJKcwx7xgyce+UmL6NX/Z+NujKHf0g5H
SzIF4ry3tTWPE0RW0ebu5f/xQIfx7j4IsRptIj6wMj64oo3PYSHlz1kLuI7ueBlnwNPEFw6bzB/L
bnpW9Cbb6tQ8IPb4Of6tjTT6szsJeCpW0/0XHQsFDHv6elNcdbUMIYYuGFRsujzbJOckrXmA3uF6
Q2U5ngFaxKXlZ0dbViAYid9BI3AsdOSYwYYGv4UFO73DhlQ92TSn8v9tUidXCCQXTcyQkikZZl/1
H3n0L5554UfIwF0y161km0wSmUrT9yS+PwiWuNPS9RtwlTSjtbyzQCxxzyCGmn31OeqSvhy5mq1F
5BRgSbc2xAjQlpPdCc5j3q1evaAEEGnqH6Aj52On+nfFSN3jbrCXAiHVf1bM9eGOZDAfyHM7/5No
/XoiSOwt9wloVJd87JaWOJxafEIMqENGGGe+b3MnVv3Yt/UG4rd2d5h5XQxWcqrNBN/w9lDEJ9JR
CoDHj3tkzabdds3aAsrsVhp7J/Lt7xyYmSmQouPuZHgQqvkBK+HSpj2UrovAgLsrgjdwX/H/qEE/
0TO76cxt9Os3UwjeEKCk5JFa+gW6pHdgbMljTW5i3U5MMv0iQ9fGun6sWia6NnhraJZNxsxd+NfK
kKZGJID3BSa5ZGrySd82AoFPSHLc7uDEjhuxFN6OvYgU6l/rVJgA1ydhwGRZnbOor0wV9QJM3CTO
9dpbc2CVwP3zT4GsY3ubcm4Nl86tc/UahobNcjHCuekVowa1hzO/664fXvWNWcBVtO75V1ZO47cH
8tceT00mqgLD51Lf73icLVK2B7gCr23HV7+uVqOIxmBL6JZEbHZhx5zSjLSJSxtDfZZdveZ53hMq
WMmxbcXQ1G+XBc0mHrIQ98BnbWA/s9X5ieJQt6ucoL4+/MPDWyjc+/6h636fzjAxk/E77m2qo/rB
Ft7MVskybMmOoSxYOuLe+aUVPDiO6szVh6KJhqtNcbLXHiYBAt9buAviSVW9cjpEhj4V/zp4kEoh
pp2xPUtGWykjmAO3QgvOJ1W8DKYHUNWno48oS3JVreXhftyDGUq3VB+7kQNNfTHn50XmPS8Ku3sc
cDxFoyF9ZtP7uFXHZ4Z1ZVWg/oRikEjCG69ABOBnlfTx69mkpEgelaqyhSyP9PIHyY/k9psBYE1n
69upur8KaNa6zD3rX7mLn3To9+2X4OjEzk1KCR7QR15tfapjY87Nz2bganS/29hDxMD3D82QgPh1
Ih593++81PMAQH1Dr2SkqP8+FbobuySGoas07wN9RpTtLPMq0TooABHPXFbKaGmyCkWvBqfib8Ih
eik5Cx0OhAB46OfA7FSRcu/wztQC29ClEGFrXQaAAUKU/bhE83KtxiPNYtlOABeuN6cCqodmPMac
GCqJaIDLQj9J7O3IZ/pND+crGPzzvEB6qihnN0Am0/Qnhx9UcYztUYkagkPXUs+0jyIn7YtystOC
0tmhm1hraHq04/XhGFU6iV5RJVlBTNcGEhxhQyCy8qnAU1FNlvO9VweSnW5KJicbVsbf4j3zGeDN
iQXFTmi8wCREBXY81XTPFDJ1RkVnf1WscGHvVYuC/AG78tG4HSs8CgPgrYbp/WfbF/iVpSk1fijs
efxcvn55qmTiN+KxqfBAmXboqhSu3WE4VNwJGuhi9/KiCrb5+VlShVI3YGzyz3XMM+sFPMn4AAg4
U1zuH3r2KkZDQkaaxJfOljODMuwT2DCzypQ6jf+kNjsKG7MZww8jkFhNME/NoAvlg9O7P0bOf6qS
TMVnLPPOy1Qt6As3f4QgNIqeL2IgKMktbkpBx0hQYUhgyDavfysjkK0h09/sYsXLSTgiY/aHCDVg
FEBaXPMvDfw8VAyKW2YMtVth3OgVTL6sAj1MmnP/ZISsBXCUZB62N6oXPbMKjHRcXw9q2PxcVQc+
U0WKGoY6txlQ4enb3xP9jQe47SrfHlHAG/AeJ7zSflcC7KZIRhvRvsp1wzSp3pP55viF0yd5kbsc
LFhyGYJm2FsFxC3pEKzOHRb6ypVWoGMZYk3EL00hOpkOdLK4sTZ6DDfQdcFyJojmLsYMXtOaJZVa
7kTPhprgcM6i3hTSTcf13qrOTRImUMC6uOYl322RrXEGMIIjm0b1/SgqDvYdfid/riZUW4ss91IZ
VOfkqfiEPoPB86VUr0AtniffRVnqVAr7yOaC3iZyHircID0V+vO0ORsEISxzmPpe8gGM7JRsI5hF
8pIVTxtDFB6O1DyMP8ujY/N4Fn2pdFLh4YfgEE1NGM2GdvVp5px5A3UtSqkJRPEZGwKDuXz6XrKg
7uEox5rOBquq3i2uw4R41isc/TqKT1fCz0Lq3GgU4NluULM3vJTSZHx5dpMkqMXw9xytJBamjaaW
BUb4opeS6pDfWZaodbqhBDGxD0vxSGPJeXUaW2FSkBYI4ah7VokQX8/OLFq/ZPlGxf4eE4X7BXiB
ge0eoqmyQD/P0g0L/eN4bxlyOgIHDNCfiZJOeX4Q/d7wXHQrLSOpCt4YxHQZHivaz9sKPqwP0OWq
XLrqhwbOhfiBfgNEDkcD/DNjCh64ElBiQsZlAc2L7pZxiQDLUG1kBh6+6C58cqKzjnOmKBU8sWcK
pAayWeKxdDupPIpj32zspwZV90k5h1ecM7cpY8jFFYYy6M97DUIMBv6RTS1i2gV7iHW7Kh2ksJFv
RF6tPiLkK2p3kCmZ5AN06pOBoftF0oa9739K9TwxlgyozNY5K3O3iYA2BjnKpU7JrMlXorZHtCby
V12JZd/0jhZzlmhqbl0qJ7JrgvrCf/xu8PmPwX2qqkqsWW3UCVudKYWgkgJqU2TFfDFfxyhWa9Cu
0Sg9BGaCw7kMNMg2/JIhGrL1GrCz1NovAgVV1IThp1xQr0TCg63tidNU8VN6/6fZTKWck1wH7J5t
xYNE/T3K3mVj8L+eUYiFIWu44Yv9+/VP5BxAY7eaJjB6vXfL7yaOjno5YzNKHZIR5pwjieHgBG8h
dscuMOZ85aLShR/x1GlQRMJFonSZKvqeXAUYvrUUo5V2w5pucKjTywTqXIZuwuN11ZAvAeWCnb1a
ZG8ph9hHCHKbKgeHOIs59+IcZrrj4Nwhp8Vk0JHnWb6wL7NDK7MtJ5GaOaon046ySLH2QRlr72eO
/+6UQHmkHZZZQLvXshXACZyF5FJuD4Zd7TZHv9cOK2MBBY20MIq/fqYQ+SsTrlS19VZuRZySjMRp
PXbPArn7FJiY6yQmq6AWwJKNZ81oqdBuv1xmWP+1WM7tcmcOZ7jr9//McziNSH6FO7icECbKxLhq
oA7kDijVsw9chYzKDu0iASsS4F8ZFsKHpYhOW8iIWh5LPuMu+72EP35BjJ2CEaOvhH6yTSLG9mNs
9SZzUU5u76YzipEzLqtorQDjfwhtZs5S206XuBKyO6zIzV0D2fniTyBdO8Tsrb3ji5XL9dIzWeqW
iXU31mxRsZ4tnkwN6GLOuuq8pewsgVTgQkG8isNmhUBwaT2xyc99vswmWTUAiJbaq4PFa2/g/dYT
0quBLhIG2Q26Y6G6EkHL6hyblaqyM86OFcLI3u45cgvrOzKzaTTUdaCRRbsjKicInRDnId02kMXf
6AjNPJglkSTUdrXXk8gZ48LtMfBb9ilA1SMN6IP1fe5qJg0k8z8B/99clKkQ2AKBASmEEksHEhKQ
1cbw2P8u90d3YPTtm1wy1+L0t2unceRnvjer0qrxS+jBrE3FVREkfWSjeCEc1fQDQODz2dzX4P0m
8toKeFzDe4iSpy87/IH4iOskXBrUOf3PP0iAqxVGm4oDDC/NJt2GQw7fDz+zUrMUAqW2XrZQVBRu
ZWsxfpDSI23/ApInKGg4zUJQnr7VEqPXIwXICLmFz8hbQIKCJqPJGgg2oZgVqoaEROHEyxFGXuBs
NzLGS3zeNZmftEFtv3L++atctY29MhHkOtjwAI5WUi5kVrkV71PR+ySi26vrvgt1uArNuB3XoJQm
bTN+S4SzuUDY9NA23Nhmzf/i0VgOwWCkwpI2j7Dc5MItbgLylvwSfyMWnfs4LVlTEF80ntPnxT4e
NE2kp33YNcoYp/+E49t+DmHkvX0o3e2sPELFG0lXGycDh5CaUy89fEZTrXBlqbvkLwgUd/ptEe6g
ykQlo2uDJ1nxeUgW4mxUkFbOzwAthrn44ltNDQmx+6K3iY+GW9FsnbYNWhIhs8T96xEtvBvejd7G
qyxxO5ZyuwJh5Y2Cak+lDdwlKKdhR3qe7Wa/eCvNfBcrymNYdapm8RQ/WOAoGjlbQmnRYNb0a9YI
Nw0/MdSYL+sgh7WSF7nDMVchzQIvkVao4MWmDrmWPuNKXDGAhtkgloBU/D18VwW973dhoYw+YTS8
Y2Zi8egcajdhZ+UjVltnNEBlECXaDjwso/N0ee+3dB4fkkDM/CXK8acWDzkRLGOgs4ggnqtvJurz
YChEI6zJTi+XSa4DG9SHKsp874eHcPUzra56uueUBBzdb8JYj1cXi6TUMB/IxV3P81aLJg6RMoXK
wLEdUIaS5GKcjKxlRIAeB8HCRH15KoBbBukl+zQhQ6P7YrOfHqzUNVUJPpZ4wWKV9UXuWAsU+j1a
w2E677dEJRgif6cR957rZtQFUhT6yHa3YQQ+4jLIwQ166NERhUmriSKxMYtulz0D6bnjzDMgxrwK
M3xf1tgkIWHdcY6o3MnROqgoG9O50U4yoM/9IF3xiS5oUeUBsF3wIHtWQKFD6QyOOs21+OH7Qrsw
kW4+6qvp4Xf/pHiZxiM0pQKm5C1FbABDFep5hfU3CdF2yjzPBPF/vMR5uzIRpAfpTlWzQLs1tbA8
YklmmgnhbSacFyii47LCalOn67mT5lwW1QSb8XTT3k/eLiFrADDpEtmR15r/oDSSy5Wreh/vqYs/
qkVMlBpMNGRQWvGcOiLu5iEth5N4iGDq6qIdJm/vEp/DIVX5rhoWU8rhJLzYlrgRSL4Tkr/h7nEf
19ek+ybh6R0HTpX1928fkO5nrUwUgWQp2wMAPBn1mMr2odhUE6TiLDfJX4BvVNfZBHEuZ8WSyJR4
6u6I08ZvBxVrBsExWeBckIPT8t+mmFiGrlBqqw1yA20VqnSAR92m2WK/jPP5Anv+yrf8fPhLcYpo
I3W3/q+nPtojoRMd/5pY6+CD9yTZeTB2T0ZKarpSCcpF6MgJ+9otHflR+hY0/E6MtNJTQLt0I+ny
GJutbsdgWgRNF+ma2MkVY33hdjWL4EqMzVxbM1QKkJcmLGk2xB6RM4qdAU3gTt9oiErk3ckMjVuk
d6vbfSZ85nSWIdCXbaFMZC+SOM61qvifje7nG0LcsebgVPvmSWCnfon6eS/cvH5r6HU76EAok3Gh
qU4y9wNYIc1tGWsHW9IMz9kuRvwg5M0dWePmQvsqgnZfRb39xKiTX3QnFhn6uuDIYvtFarNbhuvC
pwoveraA5Ee//rip4rML123dBSU5SWjkcoQ2GnyqMe4X8zXdN+HBzajRRD/ehhSqmdygnFA8wF7c
Ps5LE7L/fqwcy5h+CYQDJHQJvbe7mh4s45RbkXWbosHuibbMz1YVbRKAlRlmSKW1duQF1mKFQSAW
4bnd03jrvSMjTdI6z1ZCMAug/U3iB9Xs/tK2raCUGX+SaJyJtO0dgH8vzAN90S0SYa/whOC1d/8K
RrX7Q5Nlo4XHIT7zvyw5zyzdvblrHWRVQkiSme/2STusfg8h/BeNCCn1udDEptWQZO+rHtVTl93I
4zfnqUBVSyQ678bBw9OZiI7cyyYeUiwr1b9eaDX60hAE4tLYQ29Et55HujK8j4anyHvbDNOy0Orz
4CddT16vzwjRo/hFNumzp66j+5RDY6KguCv2tt72L4+4v/k2l41VoxoTA2TDnwBZaob+OV9OyJPn
qGIXhlZauBvgUXvoJDnRKMcg5T7TOhph1pQ568CTBBrIcs/KxuacmRyF7tLec/lIdSMpomXpgIWX
bFIMKMfyJ7lsrmSmM7Xzkm/HOZ3Kqax3UsVc6xoBh1Cdvw71bsbtzc0TooizPQlsx9HOdbF1DsJw
D+J8GTY5awkIyzlHWAxcTb1qIpwh0TDr2yQTkM9j79JuXQwTxFQOET0i3v2HB+Uh2Xrgha4HH+xC
R6vAz8QTdoONuZfw1uszKYMV4sbJFn1LoWY2XkhyvEOflMxje9AUz1XEJmcuBWG+77fKPgYQZIyM
9J6sqyuKFo/G9Cy/sVF92FzuqmSfoHV0BeAJDKUfMYkL6hqV+U4nQWI9sgawuputKHZ49Rj0Gua1
di4mv7b6XplgXQVSkntRfh5kzq0UaD/SNamrUamjHhUDb2/jXQuiEqtymle5t+hBITaWEr5Bzrmu
XMZLPL9Og6Xk4555+qQ0hUUlg5V+RcscytOJgyxtqflASWr7sh7WNNmGmlxox7dh3T8Cip3htfnE
fejHu1eBaowK79GNh+2SIh0BDxsrcmh0yKnCNul+29iegGh7DV7iY7YYZthma25OT1yMFvPMuLcy
mZqk4d64JhTY6+WzahNzzaDEnDayQ3eSDP6Kip+8YHk3ScWft/IKSJTipvg+VZtb5rikEkPjN2P/
wbB+X1xYlCWGAcVJKsJk6CECozSh/HOdm5dYDh1gQ3bhBrGr9P8M2HDrSHDxraWmixYtDlgAUC+r
hvJhaJ80Ae6Lr60hBCE6UoYBVSDHgUtLW/uExwH+XkQubKYUy/wQ0pZYW90fMF2FnPuJBOziCpLs
y8+2+Kdb+TPSFHVpFtlY6AtHRK0D+AX+fKU9E85JQuU8mhfKMlsOYCZ5tH2hDLZGPYRg/VQR55gX
wNd7XXIWUIQpyux/Dmt7bW37wGEmn4zph6Yrf6roH9aXRbPM3dyANj7n1gDxPdcfx/GHmiQBPx2q
oVKufvq26jZNFNIfS9hu+eItyOxdpG4ERpXNppQUTKlhjR8CucHIqVNUhI1P6AD999VzdG+/PoJ9
wN0Vzhf6+qrNOzDC1llgSPz2F+aq3kBNzOxNsQAOOf+renhA4V+r4JiFsjX0lZBEIIFNB2ioGbd1
MsramKYN/lNE96BszA4dZtRs2Tj3acxQSpJsQl7KMpaJAEyGG4UQF2bc36xlP+vJHUakKYzZfAkG
lf6oA3iyxWjHyCASz6+qI4RqxlrEl6BylEWsKLKGZMPovSSVUw9BEZ4Gcw/MXybSKffFGbcEciBC
PfC2cdx0cYiZHAvSF6MPI8mA2nWio1hoTMp0Dwh2bhbOx4nEAjh+FjlgQHmPW3tV9kWyJif1w9yO
JbXgV6skcLz/V72XTYnnypBwdyVtlDY+TTXKTEXF0HD53XEmpvZbzNZqtHhHkx54eBXV5gq7hZ7e
66406WGcEEqcLhRQ83Bs+LanFcbiyfdk5J4YFkjQ1ZHhQMDXNGaFR8IkEey2cfXzlm2DVly5Spnz
u4088acmqL6gKeWNSJvh2Z67qy7bRzxEkTMch8J3HwHqRhqYzmzlKB4LcowbxLyNlF8CHv7B7zRM
u01iFzYGenr/JGgSlCKTD73SeyQpCZjRVrgdZltnDoZ114z0vr6KuzPXSx+o10ohmhusrM4HEHaC
FIZnbrIzjzLW1hrJvSp2TSS+Qyx7iHRVJySCmd8s7898hdbV4shAxULsJ0f+5OvcJNXb4pjHLlVc
Pc/4n5fPri/elZzwTjFhPzhDZqZ2LX9wSPAitZq6xZpKEkTSskRKc06+ppNLMaZ4sCj2iNh3qoiv
ofRHEnvNnIfLh3CmGFzIXCmARRwSNSdgKNX8kjol7MHnTcBZmYfGP6M65ceX8mcmqxT6AsGOBnaO
BfZ7ETPOyl01TZ6X0sveCDVCs30yieHHlLDy1C6Pbn4Orne3+h4GkP8LzN1MpCjDugMNqjyoprxO
mpAgHoJ1r23zeoeUZvsp8CHBYaSRDsD1nTFI6KEyWiXhYrOA+OmI6rqD24GX55nggjjS0ZHxbYo/
nfLdo3/BCmLri5mZl67Fa6Xq+mIHrLLPqCRCQ9ectKOQM8QRut7RsAnl30CpnKQDKK4BME9eSveh
xdDyvE7WQxyVtWZBb/aGBbTo5v9k+i8tphzoxAsemWrbEMtbtDK8oMRBWcV4GgPfopdCU2smk5QY
xYO9cliOhyqAfAmY1QHymiOrQ4mf7cfZSWlF5A1JcLkgKcmTfdAYqH2uoCL8UBO9KOXQw4MdRpoi
5TpP8VLXKd12O/OQ+L8AR+FlIcrDEYdD5I4z83Q55G8qQYGcq49S86JOx5GG5ixNGCNPmqOZgbCc
83IPporRhE5IwFgaModFwL2PctY1cLfFZ5Qh7aWf5WMu84p+j/32JksQdK8gShjNIDk1m3PJj/rK
qq8LmJiT17HQqc/we3JAf3E7EJ4zuvdwet5HM3X70BJYcwNzXYMXUXyMDS219CadUIDxK0+pSKOB
0UN6+YMriXmzpL7bkVq/dmTt29lzN7DbwQRzMxLKpbXun6UG70Uh89zqSudaGZQ+u/TO+DVQoM8F
CvFh4DADn264L2j+g+0gQb6WO5GC4dYJmvK2wZCG3BjToYwfblR0lT3bF+iW6/rXQvvhplmJKXDj
wcFA6iK4JA2TCwEGPTfuWxLshNslzu65SsDgUrlLN6ks7yYqkqs5v6aumq5Uu28LCO4WZDovo9jD
D0gPaCVgyyjAElP+KcArVYKCcZ7bTJRM7tFok4uFwJHVyZFlQBinAhtReC1UMssvWMvBbt+vVsaA
pJ9g1lcyfQXx6TGsvCo/783pU56py0KK3OeXx2PRAKx3Ew/rNSh8Dj5n7o895ifA10fJ+DL4lIg6
ojl64Q/sq+VHuqWbBUTi6w2KXggm6lL83HYECFfa03l4tch7vvA2suU0YtxXteYbqOJAjn36uhJ4
2Pi2ZfxNZSxilrO0l4QGmI8cDDPklhZ/4ct/h0tEIKW8MHAsJi5F5TjZ8eGP1BT6wMu4Sx490Z/6
LPQ08cmEkIuc3JwnhuuWOmURr78biUfCa4v7IfOwlF0z7FOBai6ikwxPccCWJcDAHgJOPMVb0szO
3ZRI9raxo4fw/wPDr0jsLCUw3ZE3FdjorsaIs7MJ+U1HSKzCKOv8QkRXYuuqgCUA07YtJr2MhOZ+
1aII+h29t122lxLEUzVMvrgNkV1X7huBoJFXpjhLatRThfiHKNeIeZOleGKKteg2U8tuOdHhvhzo
09b22sVYNizUqjsvKKMSONfJGiQON1bFeUh5j5SNvoXYv5WCS/yhGU92q2Va01URMoTZPs+Fe6oy
OelEQIEm+h1ua1sqo46m6hJ1ZYomOiQ3txmqCY2OuhsmKri4vu99mhwpwwNRmtMNFNSQ1F/okEPv
mf5Iz+GJgj7rcm86BLK/ykcHRow/Q8VmgnRPim0j/NGtA8nAPEsNehKI8YgsuQYvaPjpZ/nvT/v+
83mV0/U22RlllDwFLOD+9yoHZwX6jhczWdS8Fm9o69eUBC3slC6ana/BMcF1jbvpZKvIvHK1ON0Z
ekvi6XXgAXnwg+FNFjaa0TJL2xSQ6Rl2UCvocpDZX6Kg7oYuTvVwMnoLHDMzrmbS+2xEUGYkuIk/
IAfCtxHZ9kdifS90tgVWwu4wxYfuXIg7XuMsqodMgypJEFRI1547Q9W6iCcg+YipnrdurlG5P/FN
cXYM8eMehW9pxpnBEejIWWaQwmiAnm/WlLdSGGt6YgY5aRJWrw6pVLeHxNeN0LSL+48oy6Ji24K9
ymtutinvF2CUKLJotA8nTFjbrQz9hrQd4fvHbVLH6s5UztrFQW/9nix6vsFUk4mVTlX9P5ZS83yF
BkwlDTAL+KZoh5UuwvaJfDNP0rDyu+0susl/RjleS8lavbM8mAkv5kjFufnbdwB2zEOlpez6MJgZ
vmWtY3jRc0Ih8oGkpqiS3gA/IjBzqZt0TgrVW+OpfpNlqMmCsRFLj5hiVmdeAQw+BU6xJPF91OXw
yjrxXphvoDcnlSZDMTo81TEqGflyY3SS6cJXiMkqJ4UmKVUy/h6jvWF0W6BBxpze1KpK2I0tZH4p
IN4nD9hb58K6uUvHEQPThA55XSzSdUYgVA6/NCcnIRmr539eIpj+eYdgagcv0Ba5phv2iEYtU+xU
xe0jhVN40h7EZ0p9nwIgPycOrsU+oa20qzypkkAn1zrkPSA3Rcr5dRwAH8po3SGBbz3VGL/3bsYb
oSS5ST/x4qiYXaH+tgibljH9hMp4fZ1WfHxOowol5+OhkqlNOzc45Y7XiAIh8xjA6JRvj1Z4qzKp
VD46U4SsqbyLPMMpWXrgSlC9sM/NVmPeMEORqVSaP6cBvw5rN5hLXsHmJmNyxmXYIwwjbWsqJRma
1qe40qgJlkw8vysPFC6ftGXOxeUl1b0SnZcvAyY5qWgH3KYB9phWT84tajcXT9aMf5QXf51MV9ss
VlpKzP/8FdM2/vuAaMIvzpG9Sdv3J7BeGLwYc7hVFV/+Ozro2S6c5ZtYn1rgaIhoHaqNmEkjITDM
jqZkpSziKMxlDdbVAzqLQw5MYYBoGpGmVfRyoCEG+dCImCVUiCzf3tV7ycEdbzqNRKIlwxRfkDsA
qVhEJ8NY3JXXQUPY7obLcAA4t5zxob0zJ/BDh/Gh4xb6P6gC8UeA1QkETv0EhK/aZQqm0YMB7sYa
Ld3ER4zbGGTwiYNJ19Oidu6DCsrsOLGzOZkemqXkufWkXOGdDQCJ2SNGheNzp3iVZH2KvX67hG6C
fw2S84ZHDxTe5qMEDwWdfwYP/48XukgwyxPpHZEZyF2r16kYPAHuZDkYE4Xd7syQXk+rsEF1d5LD
sK7dREGQYXO+1NDK3Umb3FTVok6hr3CmgCvLCxQqXcH/U4cZmjUuStjZiN5+scHBiEUr565uwJdI
Cfj5kRg5rEN8xX9s+hvyDS+kZFUkWFfrX4WUsyyzefKi2blrSrQp0Yfq0xwT9DFjDyuUvCxNTVIh
w6AKLvKMmVfU3hp6oqOD2XZwIFcr0nGTcfetQ7ErT2FfcAOvPx9Qhb93cvjzvdz7HrNZDI3NxgI+
EWxnBynyAGawT1B6hBnD7NFnP584P2MBmjsj0S89OoZQOgs07fHPXpLWkA959hphoRU/F7lBhGSN
r8vk7sqeSU7MiuOKAq49k6fsAV0bVI04e4RikCwhBG6Jhv1RYfLlMIPlPnLgU33q2U/u6lFgUue/
/o3339OkA205LWX9nryzq4bhKRheYh26sYFkjY/GYe/DSvLfx8f5EaUdrggH4ySx1bisF9362Xo4
dzjKQYFkMF3Dhl0qbUJzbWD95ufbmHSDDtBO9oB6ppu22Xfb7xPd82f4bzJXcb8MTrD0w1MexIzY
89YWB9Rii2BZHm62etw/Cum0XwmhEHDQ3Tz5GNl0MbWaBNkv80Yep6Fl/XY3+80bZTEWdoBAv/Bl
RgxORm1tHm5yx8TXPv5zF1ZkrarGiCt5nj/pSD4+NGFHxEvCaXzhwu+95/xSryu42rCfW//Ecq3b
nnKqISS0q/xSSdQ7vtu31lm/vtIrcLaBCFJ0ZYNVsX/HEazWQrjdbLS+mFZ4VojWlSMO5ghEwnYY
lr+2VPknupdgeeBexhJMHr/l/0Me72Vp5rYRRkCJuS/25pecUXuQUKGnJTqSYwtGHcAmEyfDWh0r
fur4o4GR3cHQ/AzA3VPPcpgc8iCf6Mql/bPyTo4RaEQWBP0c2RlMEtV7wvmRUK2/NRmuGSDRBnQt
5grClAkKlGxMKcIan3SJ0DtkwPn/mWWkk4UDhUqqy6xs5YZmdx+I1GbpgQNKdEkKUvmtZHdEy3E5
jyN+e+BDn2Qm4K9hud3DU/2jKNU7BdloIqSTWczLXuqeCFH8Mp34rfg2MnMb2/+C4FK5x/yL+jsz
BloiFCLCg3hQnoQIomlqeYXytqUw0WxDg/KJH8txCYLMwFv2rnu/YYbQi+gCjtr5Hz7TVrpw4VSh
gzX6YOA8qclHWOgdcpQwgVSJ64yUhVr2B3a2J+05krcJGisGyCNtSUce7bw9lsK5ohHgcAJm3fq/
EluLjwB70z7FtIMN8aNd5EoUduuqOML+stxunkssk84PkRWIn0TysRdfM231d2Cl0DYrOUfrNrfM
VFjzGzA/weDe43Her1v1qR7OuFsEOoCCY0L+tnPekwphZXpDdLWOd+ktMMyOOwybfqJjVhyNJW8G
FlaDcpkwy0JT23tPmWrdpJvggLD2BTnVkTyJaamcIW2BoDlZUWv24hL3axhskrDB2WvX/1xHQu4z
tv+AHlsTZ840xUpmKaCBvaGEfcd26mGTM+7DuJ6Y7Krei8gUs6XcpZArxQj3BCpGIDnLE7nyYVfd
dOozOy5N9SL6ZGTs6OUrh2JH2RpsFj4YB8ogVZUp8YQH2b9NCnjgL/EuJ8rHjF30Gn2Z0zLXuMEv
48kWb4UYfk52U2/KQASaNiyGKPHvpn0NLsttd2DK85sLvPRWZCNKqLo65Sk9HJBI+7oGC5To7pzJ
nTZhQNOA7/Lb44AePG60CPWDXmgiuZ6POcUJZNAwjTKaO6BlyNtuHLXu4GG9ERfmfRkZ477crj4U
bKfGts6WdA0CKLz+GmZWRKLqA/x2f0yWftJOTQ2g6XkoEgnwk0atoMJ9HVAKAXsFz3EFyr36zZ43
4Xlp4Lu40muXbJDWuoDl7o24K5d9wl6nEi/tRYzCfVKLnitxxpBrkzW69EBaf2tOpTTH8jXEKkfM
RI2RHfEJGZ7uAtxf1kmy97WkAvVPPgf1QMAxGfb0J4DdcTm11WrXOh4VGX3An1yq8no2VsEPH2VT
hTCcwlIctQyLU9lh9mO5L5ojlXdrbCgdaVmhj1vBA6GlpTyAMcJ8y7UWzqoq65qUdHLWS1YVu/r8
miSuR04yaYotPmDwGE+uzTmndJOhWpv6Vw7HYM5p7kkRC33y+izfMdU+4nxZdfORUKdnA2nioe1c
tZuLb02wm0Di3DTBaBGuIAZEFJMiUvqA3ae20+bbqmK7HW98UkiRRf6O6pzfPf7uOnSVweMi1Fnr
vcUGlucHcwTvypZjfmEIIV9Zcym3d+aq6bdRVof390iqfwnmeTcRFXBA15cf9/7G0P8EjpTj9zAH
HQpYIbDaLzMSzxd9KnG9BKmKtnlu78nZnoytAvrZ/WKkcd71XVPwGNd7xV8CCyAKbdEzED1lR832
FaMvvY1vYccY6OUUWbMl4/Vg/pTfNFr4QQvtbrBgl8dUjaBAXDfcyKnHMcotIQfVp/Eq8PJrSWmV
oI+KqLFL+hgUwWtKxceCRYLUigCkh9NIVsJzla9uaWyVwoqE1BrjsbKq9dGMx8CYwfTzJqkYfEh/
gTLcthcamQDFe4S5QjkaPiuDC/8THEk83k2fseuhr5Hq+37W9phhj0ATiY+x9UH9FMmo1bBy606w
uQP1KQ+WZkP1+Xx6+0S7Ic/ikEw8kbyIl+oXP/9rolNUuCAsulNPXEx65f5mje4QpimCTGk1DIbp
FvbK2XajZIlgopY0qb4PvfTAWq8C5NVrsKqqbqKCbYkQCTtGHJM2sz/MQ33Ou/Te50wKiO11CxSv
VCcffc+w+smeBo1KpSmdt8vwPtNfbAa0raLRh72FC9abtCFObOpHA1pmfihETLAYWWW16uq3VQdi
LTd7WOI88YuzaiAFPSmmpvIDxyMvxoH+FVPWMXGQ604d+xuOpTlAsaHOsljQhheJOd3aRg801MnO
J79rbgWh9hjvq2L+upT82UQ++gjzGAqhIkBtoQ+3QFds4QHVaZvt4h6rP2p7M1vLoLAqSpeRbpWd
wbBQJ0KAvkanahlPokGmezHlq8UnURBtz5bTMZAPiw980800ybc7oIykOtr5qzm6OSgu8dQy2MD5
+XnRpLJZ+TgGMRf/e02v3CWbTTcF51LHUGZAL+MJ245l/zW7xqol8FTWbu09LU4KHJLqFRL37Bdw
O/A37ghP2UWw80NoVL0CM/OjUBHEVmJjaXdDW1FsyekvWBmbL10l+3GmvZroj2bPh0a2hk5jJD5w
8zsTIjCC5RTn6F6VkfLeVAtYtvKmWVg2hdQNXY/72FwL68c0Jf/FI+s1Dr2w74tvnxXttxoyV1sF
GSojq42aij95+9ySs0fXmtDt+x0hrTncRX1Q+zqeq/LjUsl9eYrPo2hVZQIPk9f8sgA72inIXbHp
L9YDbA6bdgUBFYf0T3LZXrPBok3Aaqld1DBAlMTeIk2XJon9SnRnGq2lfOuogyi2jgMtReyCBYCw
vJ/E9czK+SiBo7OW+t61v7Riy2ivMQqFqbaH+cBigRj2I4KF81B0HibC5jZOP1/+hXpGS0JCEvEO
kAsiovam34X5I/A3RUPrmhj2LKzYpGj8/32cQpjUeGlDgqbLIQqYxFKJQmES5OasRaidxqkUGZaG
L6HsA626JgwCPA+jhR45CNJHRhsDWnSjG6USBwvenNMcYqNjH1DeRCbRTILIikPtwdDYwVipXjXD
n5bCX/Kw7VvTJfiTPz4SDZBWCJwjfA/BM2NKHoT3QD+Bw0xfXJl/EVCzL1J1FhaiGoGpOtWz08/x
cmHBi4nSJXTj8tNkOkQHWzzZrhE5s/81XUnJEO0kkd85U/h+HSKfqPwpMYQ0DCH0io1oCvZMYlOR
AewZMFTnO90eGLiRq7W24ly45pjrK1h2GQBF3AEdrQqe6S5igXmOPZA1NbiyECufDURmoTa8IFzr
250p8tbOP5d7aJB3ury9uzS5kfYNVSWCun4DmWLWFipy2e6ime1O5vTB2fhc4mTIksPoawPohlo5
hg42CTa+DejEiiSPD+lZS3pBY2Y2IVIHUceaBIPSPq6h95tXVSARjxjGSCCZ2fCCdya2i8opXfHJ
ohUwHTTiHCR9+ixpHmvWxg5Xn+iAJInWGT4GxTHoUYJd+75CRbbHjTiTUll/RBLTrHTRUJkIRIi1
E1N2122Sb9WUjIQ6QVrbCHpnhnpiSbSLun8Xd2yGIEP7+khCdUvIEAkqSN7ZMsF0g7+j8yPuoYN4
n5gJYK9G/GlcL+D84EhT+1Ww9jGonZ3/LmMafEWYjgxtdaqENBAwYTwqEcqY7YNer/S5o69pjlT5
tJQ3VRMVxibJjNpbm+yJQ2BiXeeyd1NKtooX3P2uV4IJNe/uY11Qm290spJ9rLFGgi3vEojtAhSU
lhhGZfwpCpN7hsIShYu/exfE7lq7E+SK7sqf3MGHaSESDrN9ca9h2ofrn4WA5nsAV/etPJi5ZmWE
Wf0SUoBRrL+PXNSCFjIaLULcyOJnsLXtsvbmGFkC+hMjf9588vS6UN/1Nybm45JHlTm7ayZawtAi
Muq58ynHF/FtXOjsBQz657K8v33JWfDuv92SuWFDk+mrzcqyulHKkGCSO3K5kZ+FpBtwvBlY2H1E
7luF2MBa6Cvr7K/bvISZsqgTM4oRhH+MA5O6W+8P8MkWkXY1lKbxrm4+hrV0vyAwimRI9pM6GJ1U
EOhHcqvLBbTQz7jFrYA86Gr9mreep8PVprpA/hAD/3csmZUXaaNv9pAYT4kmPs0NASExOcsr1Qlr
yC2RwV65wqWX0nNNhPTLntaqZDotXGB+xuNMHNFYU/zk1/ETvOWKPtG44xUk56Y4QgZTDAm7Jtx0
z/cA5nkRagToVrBb7dnmMzVQMY7osXxACgD50En4vsUKlE1BPCrx6caFcauuJpebOhM3+XKc/1VI
FguSe/xUHbf0p1i+eCR//sp83FXr2t3aRmmXqBapHO4kclrZkay84jin1n1W5Dh+QdKbHs7CBETr
CXFa6nt0kh1iCh9uphS0ujTmmyc+kIXZ0391u8KVp6mH44h4wmgTMdHfdSiEZ65ea5hrmXv1mFvc
2oQjiQOuYgFbwE2nmuJMgPSM/PwfdU1P6tQd1rmZJmL+C4K7Jh0qNmlBlhkGoXEw1LdCOZ8bRSOA
DiGDfUajSheDL6VgWuSB59TLWLx4Ar4T7tvkk1cE4IjVc5GiY0NqCTMrwn1QruVh6Pi+CjmdfmCu
ka5nFvjLttxA9ytfpWfggVH9ZWYsWsRflWLttC8hcf+vZrRiyfyYsimZ+Cy4gxNzuXFk/G4jz/N0
bVP/mPVwKeVNkFj26JMwEct8AlgZ1eJzyvWdRX68I1noQcMMXi/MMXTf6Z5aSzmtcu+r2G+91FPU
aNwMZXQckh7ZRF/SPQI89BOxBKNbrdYKhZlv38E49JIx6foZTdBkIp1FvVnYWdflNKIEpcmA22a+
qVNpY2msXLo+tgAv8b6ReJYOVYnhqUl7uhp+/ytCXom9VKuSx8LTlD87VhtesNFfIUVfKV9D9PvN
RPdSGsi5lxuqscNtEE3Id84pS+H2WQct+Zb320fB9pEM89suDs+nxwGiJ7MJWZ1e1vL9Jida0mIb
NAYWXusVG7PGbr55orQrpK2fthfT4FHrZXy3U6Yp4HeeXDNQz09haRugLsWaZWgBkdCsYIgSSRLD
xs1GusyBD0u5vMFsG79kfzTh8k9zNJwILDsbX2WkQxoXn4wCta+4P+ZZ1BuVU60lhbo1XzLifznS
q7HYPoe3LZrZXy5ESOlvKaWvESUiTFMw1S4Iwh0ZmQmAVPXCXSJtZ8b1V+eYr8g/vUPJw3tLHLQL
L+dFl+wXDK2+zn+ZMAhf7cKgnew0vzyBHWH3p3S45MNkZ0NR6oziH0KETfLW78rNyiZ1FdPwHv8p
OqdJsl7laqqtD38PeempVdx3gUqOeg7N/xDprDQo9WrkumkbUQtKNTg5F3GFFA3wKv6F+0IJr8Qr
uXqcY707GeKP6bQvhK5LP45yBWm9yC2zmrLFBugxda0KLCF4YzIbmQYVv0NHvLhv2tvosJK3miFl
7CxDMHNl3gq6Fyh7U9Ym+m7kFPoncTz6hXEvh6EtQ1+R1vSKD9g9/SfxrspZj2/YhPYgXtdVQLf0
qkULHFHzjtzIkZcti4ddoSw4BGsZIwfXcuGhZya3rdXf6D43/7aKRTVQWZIwA9Y2OWoQF1zO9M20
6sU7Pcl1KapnqYIopCvNxuYHIV3gCfN0xUJfqoafgzrXFkbiFUQlWCN98MsENJyfgx1Sz7Q1IAXc
OUIAuZ21em5c5KUMvkbzeBkkWIGB1MYuAwPyCr0cceg6i68NUthO9Lu2x98gDQh43/bW0WDGhFk7
ZL9YjUuay9bwkt5/L10hXoZ8VpC56h2yQxNRdFIGjC9E5yqPOZX8sf5pYa6hCSSg0G9c+H9X/v0D
zGaZ3alp37zQXpNeqOAxqTJhgq1iMm2+kOJcg9KVDQgw30a+nCjRNZd2wp9PIgftHyUtAgdHG5Jl
1m8lhdYibznn7tQAOXFb3ngIbtlJlQvuHrAxwijpQ1gTSDL+jGeF9HRHv+6YQzqAb/1yUGbHXfQY
rx1pazHZu7qXgTTx8GfUcq6d4MTioFP/8Fra4hf7iZ+0L1RgMt1x1T6bGIPpoeXZpz2YFHapsBjZ
6MpLfrrjYeihqw+Mr4yUuUvz6DIOC9U/7/33inICZ+5oRno1tdVi2TzZDbtZCscvxAXk3iXJ0nxQ
eHWFISezuV3puBwfdC0m8Yh3r1XsoqaqEulXFhvDIvBPItAxd/O4S2BiqveJvXZWkWZQB3E2qLlx
IKUjBPhi7YnR87ET3UllMxtBZM+WRQglsOTyFs0BbDoBfkCCzkRO254zt58XzOaq7EZiM2HQd+gc
3TDeg8yvbbns0SzzG4c0JjDHtgrozv21ZuaLj/OPsdlbv9Ieq/cQH1iyP7AIx7y8mCxHUvtDASer
rKQg2JE4tBSKqx6WSNURr9lXsv2cjERx/K3ZteMxq2RKRtfsIRnfY7Vacl6WmfUnIN5PXwDI+VuD
OPcSAJfy9ISN57Cih8QrKq5Ha4FYN/peyRE719I8YcSQRyf4cBfOinP4PtZa6XZrI0M0HZuS9MWA
2fk/yNGKOiJgP2NcoL+PE9tB7Qa8ljKKS03dVAKXfwD0x4uUCP9qpyxxC0S9CV68rK/JfI3YrlTm
1uDGk+yNIMCRx5KaXAnUXnleA9v2Ag6b6s8fJKfjNad+j7x1z4x1xyFuLv1/BCyUK6Y06F28fBdO
5mVPRaqA0raJE2NXxMpX3lH6iThAEBFS1b2au9In+3jcmeD9QSLDoBMh8p42/mAOqhCAM1PitLLs
EdoKkI7g21jvFH1vGscB14gCVWYvpTg1th/XMK1QKRM7tKbVEZ1OyK3/uVlGlGr/0QrfjUwM5a66
oX10C1f4VMXliE3KzUnyks/LL/U6PZARhN0qilWOvCCs/rlA8XQdYhCNkZFMeRf8GydysKFuvvYN
2u9CZzsnUQSQgyenXvAkl3Qmp+EgV2SSIHu0uC8clAJQIQUjIOf0PsMIG+55GQ9rMhX2VGj5iOwn
idqsIhTmAQ6LxMqPyaPP2kJN+vJLXu8BVv2+a8xvys1k/U+ZLTjHbFwF+/yMJC38xhVzxwu/93dP
4EU6XKZzB1co2D8lP8a/UABk9lZr74Iz2iM8cUF+UV/nfOSrzGTSakIfhtyN79oKETU7QfXYW8RC
W4pllgUdmGtM2085vKbxU20kIVo9qa7lYZ5M9j8+0UQI+V5ksM5ydahWQxb0xhThWodq9MItrvTc
JeWODkrvQkOovrluj9oasa0E+5QQX80xcuJQGtzwAgXX9IME2JECnsd+4GPlK7Wk/5nWJ5Ma74BT
3nmzVL5Dv7wFXXp0JhggwOskxK70AhNYb65n+IRsrG0Uo2lHlkrTciFElrJANjjXN3IXQb668quW
wXloTUTv/6zhONcLv6WqtcgiiolW+whmWUoACpUFTwOhO/tDGPBUHPRPPosEajBYkcKB83GG/+nT
KiLgdvVqHOA77B1PtNCsIXg+l0dXPfqA7SGUfuDkyJabLBsUH5rQxAhrrq1rgWNty+nZtYp3J7n1
aA80yTFRPf/g5CFlodMX74r/8c5GIynWZyEzjzRdiZWJ4WPNbqzFPldrz18jdJU90s+WWAt85fS1
OF75R4PFtYjsR/mDNTm9BdutXdEpRkzEk7+mIlW+0LuoV+RHeNjIgsOt7XiksoPIchmoOjBYcvOz
qexUXKCiS5NfOPvk+XDsQhlf
`pragma protect end_protected
