// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Qq6Ky1FLuH0/PYX7pP/wFvMOxbzhvGopgjp9rvDEC/lb9VvydcNNh+tnav2W8s4e
AtqwUihUHxDLOmDFCWIxU8tRmmbxaLeoT2Ek05eRK28i3tP058Gldav+3PbistpW
6rfg2W5ZcWC8sjJcJgYaxJOTjFSmxFGVq7zqj33bbjA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19872)
aLKjbJwONMeTzL5ff0JH6WRk8zKZW3M2gBHTtdZmt0FWXwiQ3hvUrSXhX19URIrr
zDLXKYnjIDnASsxwkRTRecVN6jMvUepw2SfDwjSSVFac59x8UGts6t3k3mzenNtn
KNTApTs3G2Iy5Y9lgkMUGEs3rsAngTMMb0FwEwvqyNKgDZ6fMLYI5EQedvuU0DRP
pv+pFGvJ8nKXJL9puTW/Vb+lxTf6oYk8180hzZr91AiGSz4mEWGj2tYGDBteM83S
2Pn7jEw+tMWACQajG5s5TyySnqRngEvc3OzP0xTcanPRsL6JSeGoOMzwB4Mpz0v6
jiZCL0uenaB1JciSlCG9COOoVKf61vZ3pxtH9bJkaB3y8OMoYRNOL33c46uqCU6S
r9BhqGarDQ7Yw2vqq/x8CVeo7Ykywot5zP56MCHSaqzUnZItG7U+zjZxRt1KaQAR
TgF2ihw9TnPilqoJLcKVyqxo+Ifg6eJCcAps8snlgSsOzdlo2CWJ7/apaZFlV0nb
iE19IM3aNMOmJiuNqaWYLTPv9WhFFyb9M6xA0WHxbeYjHx3zHFMEE+oyooiWjYlw
7JeakRz8JeTboF7RSJCY1YgmSypmRybc2qoHG39TLvw0TXQvjINNOzfjhq1sJq4e
pFclpprILKdSMnrCaO7isfp1RULX9ETH0gAdHF232D/04Ry6/0JCHYjBjJfJv7Qh
n8frteKzz5fJROT1VrnSsCrNn1QD24V+6d8mYN4hUk2PC87dKRW5kYjuGVJEt1ax
2z/eQ3mppcLovsuH5DdJVdQMKiqOVtvm7HMuGx58op5V1cvSL0jwm+H1mxaQQVmM
2uufgqN6e//w7iTYCkETr2euFuqXApFs27LAErLffTH/2j2CyKlbVVWE+lCpp9bU
Q/zAn8ZEyZIrUxiwLSB1Wii71JpqbLlS4koxOBk9pznvklHx23ZcKFP0z4NMIJnc
2WjmolVIK8H5PDsWjch7A9Ebjd42NeeaixxYeK0T8zrkaOAGHU2ubXJ89/7LysSq
IYq+V0HrebrPLqGihzYTF0fuB/NtnkzHJI4A641vxXB3eTScYo1p+GU7D5DTYzFa
S7rh9PANHpMp+tN99+/J1BjSvukDONDmCO1y/+hh4sgVgVSyn3yfyF7/QudUpHuI
tnQV6LkbP/qQk/3Ppu0AlpbVTDefdYiHUkjUsYIHSDcejt1yTk+iSJFb/WDLSOLb
gvU5hQwfG9uBBOxtCbM3tsTzrLeJ42RApV8v/NtNNj88SFzGUyVZOkuXUQ/KaPDp
+RzbZzoba/WOQzy3E1C016Ak5OzrNUXNd7Lzz5JwWl9SvcBrUM/ytSB9S9xkO8UK
uFpR62DkZ0hA5iR+bBhNVwgX77sa8DAF0Sbpm07+QNqqOZmwzhEcdRM73qyRMwTj
whGiexyVGZOTsq5N77wXBYpTc4QUR1mzMjqUhC8/xQpHI1mFSFlJf7D5KCsmWt1p
t0Y5khID1pIen2XlcV0BPWklkxMVXHkmmcVmq7l/QfIMcNHHg2++5DoTwt2YqNVV
h0546KPkybZO+LVjXGB7Z2pSAVHY4fevVwHH6t9gnYob3EjwHNH40Ss4hhKoxHYW
T4kwoK/rJpJi7qT4uBV+fkF7LFPIMb7Cs/1OBMBq0zXoCzXh5aozlmDoNdC3GlOV
pfsNXOLun8fvpE+V5A4M1qxtIgHLzQPN9EsgLCotM+glt/B5AzU5friF0+RWZMZp
u95dNUbLGPsXPzOrUlK2YOQ0B5OF12li7Kc81bD7nzIW651OzA6rcqxM2JuB7Tov
qlWaFxhOsGBi4QOqXeXBdiiDB7uC5n6wfhZPeR80O9Gnhwz8mCL1PpDg2ObaBC7n
CEzU+zFXunimp+XQE8T04603ejzS1Nhi/9sUvBsL+T2BnYJbwNPmpJ6yRWHtAUFC
0itKthYE9TI+A+xbxvC44RQfK0NVuIATwscLwGmYn3kWw00RF2P41evhgKbFgvlE
yL6zPg+sPXhB2y8TdzVhwU9np2SsTtRF2swrxShl5GCWsnSZ2PCKUxQK9wMR7SFO
x3tBqy3pbsdIXEWPj6vg629M5FDAKn3XY7Z4o9mptzMVN1nwjZ0a79BuX/AuPZ9c
rFZAgyh+UF8Ay/+PuxhbLCDYmM0PaMx6vIwDe6Yh7fm667u771fr+Xb6J5AfMP8o
AUbKekIHp4vcxbpgGiUcVxs7Vgho4ZkISxP0XmE2Vzki/W96QSPWae0smGQXD4TM
6vexm6LmitwL0JUiyGOar39j3rbsOaT2fyGN9r0ABvoaacSMyUPD4bwrYX7rLNtQ
rpu5sPQ3CYHoN0yntE2vjf+oeQaEDsSfzqOP1Vg24LJG5ZhkOG3AVuBz05xWOUr1
xavz3toyfbMtEQolrw0ECetyH5s+RqkCWIfsST93728hNmY8EBGsn6BOegqk2SdD
I3Nb+sQPSq/v4xPJutZ0DgdEeQSgkVGeUrmOsofhQDxFbTZzu9NMEOkW3iBNFuzm
Er/3aHkggzJ7AhW8K+Wu5v/TgPPyGGBt1IzaMD5I0iaTA7dL3eSCyU52BfBFRFRs
SQILXl4q2IngU3uapJ5s7wAO3YMvN5Ym9rrHE4RqztssC33TjkS1ehFQ1FqZj1rJ
S7/28S3uCbMgxn6+1PDL/VtGik503dONj6FS3JoWM3adfx8gqweQqMs8n7bjH5kE
r4xx9SJqimKE4ExHwaDuogxBYphnQVsEJf9sVMzHHDj0mgHci+2Oiu/zJs1oO393
72/yEhc2g86T6YpovwVE3c6ZuwQnXgVLI20jg0k78xu+gKrQFaqoHl6KmCl094kb
ZbfAdVWEvRm6lpaoVKtc1uIKnJi5cay58jsPU4DKiFuIusHmNI39EM/JRFdtK7Yv
H9agLoMzncWVgSI8Smq9K4M5WgNjo+eAhpT15JZLCKPZ8JC7ntNXMQw1OLOuUZSf
+MdUS8LrXp4Q4zdj8UyTfYDuxvD9k1ZbAf1GEA9PAe8gm3/Op8tZ7QBzKI/TXUNH
XVwXR4n9TNb0Z7BS1Mga4cZVaROJxp2j+oHNv7ICTCzk8nI+ho6Amk6QJeEwgLzU
TnPThQ4944QtFR4dL8qGEJw+0APdn+F37/3dtnPYVNSAxr+gdsc9q3/kdKREqmlH
q5u/tbnofKSFmoSiLoca7LqlT/OuRdu9/2QhQQGrbf2GRQKFg2JW/XoxLkrJ+f3b
u3k2RluiOMcvifUSqSJ+06ChhnjntDFzHv9/nyGSxb/A51sJTu02I1btAmXPjUbh
/7ySFWeJh6jYK48gr0tX8FKWhxFH5fGcBptDqkl9mbwOnsLsX49DySSm2jaKlwFX
R5GxGU43SuNr7pfw6fnVlP6bxtvJjgT30AGKM1SncNbzxuXLlMlLWnm79cnR/GBR
uSylicIk+KH6s9mUdWennIaArqSpYmWZiNMcrylUXKdfkvW9D4UIdk9Z/lrwvuQI
uZdB+hBTh7wQp03rEv584AjAnqWx/9yaPCRcLYgcPapiSbMSXkIssYbVg5+isrNT
/mTFxeUzkrzzJqsew7GIEAP9fGExZJ9d6G+OcIZ7z8y8HN6KhvdZVUiKjfVX2DGr
XDEjiQjZ6zG9is4uggwaOTF5S73jxzeweS0rgjgkdwSRSB2dWixOYK2Q3UlQA2Vx
q3x6tISSB4IgEgfN0jDNr4FInJVakR+0wRFsNqcPHQVNJAOEFq8IdSNsYpaqRXG9
I0vOajP+Y8xEHoezh1Mdd4tRY0bjzzqZekDRbDMfj6zbN2kA5AmMJ+PnJeRdR23O
3fNH/GxnDE/JpjF3S7Hk4H4xgnODVqzbAAsj8ilES93/Axwg95zhajsDjV6ZiERi
k8cabT1QIJvOj9qUXtDvY/ZD0XEIHyHcXpwHHRUkie8VaE+I8L1F9QSRXsNQUlZQ
BWzeXqFBDVf736uUmieDSh7VR/5SN7wXHJmZptCOxhd+5FA84lzbEF7CSRLE71cx
k2TdrWtx741gC4TcvUXwELyAu9DcBOfhrhjR3PaV7+oKTSWb/r5agC1rmNjKB0Sq
PGMckrQlp09nXJsU/oq4Ym6I+v4wdM4ucq0wmTSxf5VdqHKYr2wRxMGlMtQboPuq
dRRLNpaeTIiNfHNe/EKcQLDhgRwwyq1WRF1ZDxVThk0epo8/TRoHgk57LoWrSqcw
RxpDofRo45ubP2bgtUzKGp/9ZP/pDozIH+UXanwyvSa2f2+M4IzJztgCsoI1C995
QQfuosjJbgv/l602opO0wAqCQ92n3nLuUwuJF4HztuiB3I9cfZX4s6HuH28vv4J1
7eLDUEKFeLi2DjM/SL7qh0dS4mnNw+xg788gg78/0iZK/c70ejV/0FHdUcNdA9Ud
xn9GKZEmc/murJqnYZHpK3KQQqix4oKgmSrMvMmoZ/AENosX0I027h0NtQSWG/Xn
wed3prCEXhsOePUXF+FUvqdtM1czUt1xdsHgyn8VZaVu+H7ONf9JR1t6bwWQenGy
GlmAcus6PQFDh6whIvUAPQ9nyfTzbCoBaSDY4t39La22JRZ9rf/k4g4ms+d/ni8J
HfEGpGv7mZ5tUsjFhIHpTJ95qjfog8xCa1KHSdBzKV84LBFpICtCblibR5j2EsXB
WVFMdhzsZV4FCmwvVH3l0dQcXKcOwdE9CokL6nx9AJU8wK2r9LvbvRbuoVE2hRvl
e1DtatouZBesRa6s2vwVyuRb+ydtLMeT1RV2GIifEsbpiyeaU5FFOiTQ6lLcrwLS
qfQoRX8LU6ccB7glcNXrSLHNVSOuL23dSiG2Q1dQsC4lMZkXmlKUU95wPSWlG2Zd
UZsvqi8GOr7s4FfKGlK+Y/k5r/GT+Wc71UVGcB3KfcO2p5NIgMG1o+IK+D0wWSOg
3916LFVEVuGyy5q17p/F3/jxuWd443XZ1akz6F7l/Of8wA0vBtMeUgvafVZdvpjl
qBaDNUZRzOiKRTdzURLLEg7Lw6EB6MDWWEuwxCZTP1/gwyxgYnIsk4r6xrFjhvMt
QfBLr/g5xADyrekeABwJ6Yl4+PXA01/udxmR9W5ghliflyU+dhz/Rz2VJLxkhqu7
M/iw/XxwkTOyvTk1vHlqbFCKOewjomHtvFymPKzIXUhwkbAGviICZ3czE6TWC7kU
rUNlLygdvZNLP9E6WgN36TX1gUKxw9CJbNk7eN1Eu/hsHYS3uFV0cahPa5lBh90i
sKIC8hXU3ptjHpamsY/TIchNM7RoHy2CDbdbaABH5HgApl2AG5ndqHxz6fs5jHG9
6M4JU4CEmfx7znfwmCyA3K5JvxdOht82db5EeRO6hkK9vz/jqTx5T9cRTtNrpaV4
VAxYIEbyZnxPBvtulS0BEsio3HwzcjSyYleFIXVzMWbulcby1kuuo6uWUE2KC1WR
sXIfM1ozlInwlrcUfc/ZzsTt+UNjCd2Q4rO6U3SqqSEha3tDeC88nlrJ8VNfQ4wR
1w39PwJ6l0DbUpa9RftRSp1y2zlL2NK/h3C4LfcaddGCn/yjf2MzyphSVmMnuF2s
c73ckEp4WXW/rSc27Z9iXlqWkaLVgAEcmpszHTBw/jZdVPJhj1KwLxASpS/Y3biF
oZ6iCb2VqEPkOvkbpzVx6L6SRX17tXu81Mu8toMAP3mGjVgC0kUhIm7+aj2NxqP1
r1N8jpHy2mySSvoz0Mh+OuAk1ASTf2LMOKbKlpnBPDrF/6dA3/h7tFdGXmDrzGbL
V9wHsTzcFEFIUGeAJISX+6/dOfWD1JyfYdA8u0fxGeJd39AhzupTVcRWascNTwaF
Cq+rgTKyz60AujyamMrhL19DJUiZaS7cveryzs5qrIYnsG0imK7ER574W/Wxnskh
X93ND+PixPCQ8Swhaoaw3hyoPFVFd90QeZ/OSyjPJSgVahCgwQlZU4iuiwVf60gG
0o/iWlHUEJm8v+oC3lbaq/Zgp8G1P3uQfWKtaQqrvBd6lDJlJMiSMIH2nWGJfPD0
Q06IjChluspNv3IUbzKk+A5QjZb/UXahd7hQdxMqprRzd6Hhy3dN5r4GOxTaXrTr
2hKWy7cAwR/hpZDaaw8gHaqJLaPXdIkLJ/kZMNc9NFb/7hoIulgCC/ZuCWae4BSN
T0+m6bu613kinoPZ3azQ2q1wJVqv7Fju33JfJKKJ43PsuCZdb7E+6smFetgVzMll
Iet7pQLm7QCthUGtxvNdkPDIcHDmEZklPcyv8qU0Mwac2cj/ZmUFxdSuIQi6KFsJ
pitaAjEpyow4Xeblo+dr5EUSttF6uUaT9gzCwJeiEytXO1A1b4qgAhsL5fA2VUWf
Dsq43XaXMwApfiv7Q/I5TyvYAK6GByERk9ZjORN7vCZJh8RieMb0j6f+4hUfozKu
rEIWh7+WDw9jT6UYC8icgxnb5AOu4Era11t0esFaO9bL9fF0y7KyIBkUrTR0Pyla
NxPAGanBbGd99o5EVE/phyMOMoemV9V0ZOCpC/7/mB5Jq+oiHaG2Q2rii5RvUoAg
Ekt/7dIZ5+7glpq293u3OdQJDsVyxnZFtl1/kyh5odpGVwP0AWPk4erkZZ/e48JK
NuZle7Ve0IgxV6wjyLE+A40SwAX7ttCn3z1g1mvL2u0Y+JHy+/Vj/vaarDf/u6jD
4050cWeKxXnfbzl5qRLrP1Q/zigF1sulkWSqW+ITv7TJqkmGk3TDo1y69xT7R3cY
Xr3RbmkOxxbywGD0pNS45ywSpUQaGbSLnQ+qg7e6z074aGlW2v/TrbFpwKp8LTgc
A3HElKVcr72M9WET7g+vonP1WOpcYRgM8UU+svM39BWlTDbESttxauOnvV1PMm1F
VXnimocO6fGZ5QqJJ8DT49+l4/bzW+FcFZTIyRVQ4z3dPsiIGaA0oaQm/r21tohk
zkaWhGmWK8syGmstFoqTDHN5cDaPvE66YRZb/Ar3LzTpPtWCZbx8hDPzlVTwDNTv
BWJWm90/avh0IzTPfbG0eiFabwbMTNRgTbB+shjDFqBqJ6rFuSNpHWTcVcP6Xs/B
UYHgDHBqy9qQ4zlor1IyA9ciALiB0SFjWCrpNcank1SlbQzyPFo2B4uQs30MFgdn
wORh1s0yJeCVn7YeoSEY6yCNE3rFp/a6ovDGVFqs+8hR08pIXy+ur2T5wd7SDMip
ijPU4M7J6naOoR2uJ6KEIDnDNtIgbqhddy81tWnASo0YXX4Cu61Jeklteig8sOWU
1NL2OjUXWj96ij0R6UvrJJtzlX2FlOL03QjiOq1DRGdSCslKPDjJcN9zz6lHg84b
3rwfjqRM0IbnsTe9a0iJhIw6K+D56sJpwFcIZ+5AqsCdcDsU/4JvrwQYzFZyUKJ2
yqGuT+PyCUeooTePbnUbrhuqwbgl8jZNBlS6zX+2ykG8o+1rEJk8+DHYPn2L5ry0
hYsi9v05XItbvEl3uOvGxQz6RAqqfo2g8UENDT7P15bA2HI/FvcgOeiVwdx9iONT
9U5cMP2nw8dab0r9Q3VxcRkBNC6bS1+wkmTOHYHXc9oTVnCWxmlU3G2UAyDyiUgf
4NYcYULuMZktNUh1WSdngRG6FWHkKL+IYQas30vTWjcgTGlDnpZBgBJj49RP+z3x
FQndmrqNDm6upFbWGPBYLB/B2/O/6kXUHCE7/L+eBvs3cwdm/PZtIpTZPicOCYJu
FosSjf5l8FRe9e53igbDCaBzGr5YU9b3udWUF5OK4K6UVhUFbw0JKEMyoJxkH+43
Cc9dqw/eQjKvU9lwrF/y5gstaZDF/sMcODVtd6Ti++uLOl3b239FjBg51Ad8MYNX
ArCP1tmnDcCoV8sv4tz2ro/Ov9bo4UvcamVuuQlPlXqtEW5l2G17SIpzGHll4g09
4o8LOqbbQRHmOvTXXukXCfdWGC1RWBfEGko0/9CD60TCA2m2KYY+mdzbLTBs6l4H
0sxmjat/KRFb6DrDwfvFdvrO3WKggM0fATXEkOAouORO91WwVf/9q9vzfv7UzHcQ
SDSLETGTrOQ3hQ2yCOtLduZ8DGM9kwoMakYI8MZUb+qUHfT8itt8xAWhuYl16ep0
bY1Sr9vRUP3vkZJYjEJ5MfdnEkZDbXiyUxxFu1NqPbt8gwFXnlAs5DbpH32+UTHT
UIOvUlzTTDm/hJb5NzNxB28Gx/Tt4s9FWSIVKAfnNdLAXmGYQMthtWdPwmWPrQWV
3gPqiHYkcKCkWTCbn+o6YfguhZHw+w1jGIyfIFibd4xHRHNVbvf5chZGNY5Us/TX
XNfBeN+1VQx1HkKjHJ4aCDHCssridRto/bUHsFUlaE+jmgfsF2pwGdB+nhjkHavW
fCMcaiAnwUpVrcfX8wnObLYkl6sqeeWzBQZZMXhE+vAbPMMxkPUCqhCkahQf3hsz
qofvfHaOMLZYDRvI+fvPlTtCGuUcO7SZio70PDNP89zLVsWHVGu2sZRe13pt3Un4
Tfqt7454dqOaG7c+ezIZEXYHZqTbq613EUmKM+FG5OhO0m9b59fqCv2oyDifvCeF
/CUexlzDrcjh5wVpsZPn8vGS6nPcyOyuMtfqq/WaZ7GiNqMFsh37MBgMQSp+WgKj
cmq2FmrnKWYkF7Ys9cBr9IhJ6Hu4vNGnN6m+ejCkm3lMvANTeUXerNQebx2N3uQV
Q2LJxnpuVW/umRWdt1djefpm1UggqC5zbNC2VvbsMuWOGojBhqCKNCyXZlihKm7N
P+EgMO+VLOn2cOvgH3JVGA983CS4drvu7DojUvjVs9D4cfDAHK7sD4U5RW6Vgs4h
IhVPEJnD9/fkdotbKwCa4Lm0P86udTSyzQvevUX4y7Hk25gcjagT3MZRy6GIHrrh
JSoEWVW6K/erKZ7PZWegH9uWvRcMUKQvaRvKl6tFdpdK+4Cv8RkxHqnTTmRPu+hZ
E6SNEcnMGulnxT6s6J4bILVk4Bg9E4UBgLK4Fs8o25kRV/YbvU4Fvgb9V39wiLQq
vqDlP5XJuOaqMG4AtaKKEybZCEkRLg1Kmu61CmSjnB5WbupIGd8Zosj7QZBuyYKH
l1uSkJaCX8GrDwlBqNKnQPO9Dw1KFnMImjqBXYtaf15czYKLc6pXTqCtYrinca6s
5vKOTd5wlsgXGdC8RziyJKa4d3N72SFzsn6tHsjyGA00KoKUD6hPgpicl8MUDvRy
EVdvsuDf36UsCZhrurgP0tp9QglcecZe7XLIWWwNXpSAyo9n6x1GrAbtyKNOFlYA
FP1VaTjxB3ecv/EkvnQaXf6aiHz6LtqBX48aXWas3DC7gBU9UBiLZAlsdYQWxQLH
1TuVWSNzBxUepvJ7yNI6vy4NQn6jkLq6l8XfHsVzgI6OTDQUIJJbMKukvQ+KeT5V
EgDyoZJRa01rH57vUejrXunH6GZf3MuxWCP1N0FW3VDqDpYaadChxg1OY9FFICax
T2t2TWb9a6d0p8JCYsnTXLSsYRUt9hEGO0OU0RHZd/9N6kWP3oALoKdtGBRV111x
nr2BAD4WQ5hA/Gb189KM9nGk8JGoK+VvR//+XI431QHYrXUnzaOKDxg7fpPyhgNN
5AFOjZ3iwxIIrkMmgQjrNOL4FXudHdcOcuTHVx2Zn4PWTx7tpD/U8MmzxP87aCeJ
GMIvKGbE+vMJj3TmEpfPBfbPHZnxTd+NLJP651WIJ8F66RyRP/1Ce2iTflohNx9/
NeDi+C6kpnUCbbHzbxs6MGkHGsyxe9oDtfV2j7r3pI6rmnQVA4RcVJ57KF0474WO
mbye4E/FDNghpD3M5VkOjE5iovEWdg5qJMVey0yZbqfRHY7Vx2ktkczrek6HoaxN
o6hvuJ+hkmpmOO9psBH+7tfBxxL7KAny3rSuM7jyOtZDjhSdL/64KnDazAzDCUz4
PEIUD0n2L8M78hyaX+2ZOWKJYRd1fG7R/kNggOrqWfybLpaO3504IDSw9A0To90W
97/6c+FBx6ObtfJwcDDCiz//kshNN86IRqrWjB6BAQtgmDRSFdPN+lUVqLjSgcWp
PE71ZL5fzp7tjrIyLWOSa55gM8Vsjq8p6rjeza2sW9gwZVNwO+87mPVQMbdYNlSo
Qt0fO+wCbIYfkEHQ93de0x7E7g/u8RBfgSL6x9KatsrS9jPBlz0BuPpEU2uRVJtV
Z9JD+YiPsNIFDk2WxnXB6AyT6QmvwJ+3Jq2ZXNJmJRZZ8dgG9ozihKL25+7bD5X8
mO/qREOKMew6bY1wEV4IUeNV1sgewc8DiQSQfpxPbHhaNVICdsbpq+qYR/dGM/7V
fkZSAs/SrgHnt8jwJ/9xQ0uqR7i5jcQBq370k+tl9KRm44tl9V/8eXyHTJADRBVC
ZZSl7Q7kAdKt7jDSY3L5BqlFMredcV6Il3eDjmtRhqOCN2ZYHmHBpVO1lmsw5BGp
TryJrcz+MVmuippt+XqV5tQQMDL0EUeehGr5qUk8muYht8S3wJ/0m64bFFyyOw8W
/xTGRqrZK/BUdkSWiQpujgZpW/5ID5RhHgXWobsyksGXWZRVrfnjJPAePM0LleUA
SvYKbUxKXvpsP+24HnQcRRIJtsINTQk1acLT2HxCDGU3RWs2dU4WwboLxvRlxoc3
USTGqWFwiSAKPwLQWpj8qyhNbR/OVPfgO1Uyt9gGYGCX0twi7qKWYTCx2pzyTEsl
r41Lvh+Ahic/yBYp3HsmuYVkacPvR5c+TrBL267tYEJ9gOswJW6y85aMFoOWLzpm
0BOVPAlig5+js8c5KjZLFfmcbHRMbKnygVpUEacb7iHFSXX3zWhVLroKuho3CZ+M
SPAz2aGcJMUTBGWsM/mzZCEsdbikQL0zVqS3jjfFa+2uZB65o0RGUoExdeDnqiJY
aaK3qu/Qa0eQQbkKrlaXj/91UNQ4Fn+9BDZYBfQ7F+sH4ddd8nyJFaRpjU9Jzwt1
FDaGsIgDTlvJxqfgf2ANH7M0CoFnBybUkccFqB1Ec6GEQTEJT6ciDk5WU6ra6V73
wGgg3Dy6tOBvlPE9RmVb5CjztlGnGd6uwOnR6wt1WxHB4JKLXKeU9uVQP1V1DdE3
GLFz/s0YwoRIXMA27WSf0NnSbnPX8TDfR/6cYhjtgCMNynn7BIVL+8BDr3n4VtDa
ahNSoerVbExjh1+zgk9JLjfV5ABzssbrlYp/c9m6P+YRctV917l4GL1EEi0Ng6tr
up1umIKz+qlmoKqkT9XLZriQCefLWsPxvJYcfeoudKHFVr4DnIP0t86E1dxV8YpB
gOcvG+LBWtaWtF6Nd3aZZWYR3O0LFpowA2JzcK3w8cg1Wix0vmjuDmkxeBgEWAGk
g8WUyhSSdeo3IJ3iOxtpmTbqNJQnjCm5xFCfr5JqwXJHfQHeonypUrdwdIbv+jDX
AowlYTJF0VeFvqULvMCYME79xleJRD/2Ta7AuUEg8XVVcM35x/YfG9JQkztC6oHf
JxRfsgVSC8oyKt3ZvfN6yZoyfBBQYFjtWslwchAwsFjbt3PFOj7cDvyGqCwRBA4a
zkNAFZ8lpQVDSi1TPlkJC5LZQ3No2Mgj5iG6XTxOQHHUBTWaMb4/zSeEz6mm3+AZ
KNjpTGFQbSe8BSP7U1U8mDbssVcnjF3JwGxADoZWxZTNqrVof40O2lWr8MMlB43O
e214Yzmcqriyu+6zZs64StWNvGU72tdOTRX9FNqmrlhyBlxvWPrEcTsJz3u+8UEn
Jg47Q9ray/RhsiQINnU5nWoD85fOxQfX0j8/Sa0+3wjgEoZLxFCkkt80bDS2HUN8
2VPaqp7s2//m3bYxhErkDo/5aWPRUTUMbsthn4zw0aPYD7X2TKsEpJKORgx8j+vl
dddTV0m1vAAh4lM6vBEem4BgFMcwf/qNkpYB6KkZIQpX90nnyYzTAPjaNO7LcjeF
YX8QoLMWwquzbpFMEEeJ0xWN/54RYVj7txDcevYtC89wC4A389SXy4zujRoEZBSS
75tzcAmyqK1NOPfeMOde+kU7z+nDzo7kXJ0OtLBgLAujuNIk+h2Dic3l8VACpi1O
MDZ5bqY9bdTA+gXJo54qu03EgzHrZ1ki3OqnRTJU3Z9SEXbooyDqEsvwUOT2PL/T
Y3uTt5y/fsrowFGKSywlZLJntXhxO4Dj8EJXiULoTQfemfBuDKmQ6Zhp6mTrERrr
YwSS9Z6U6lZ+Q1DVrG/D5ZFSWBV9R/CDcEHDM6skqee9u5nf6lhmi2R+jPNg7fjY
nJI7cDFJhi592AjLYvWv3ce/sFIKhGvU9OdhY/l8BvdzVx9fWIU6GgCKA3ojb3nz
pIHI7vMnn1x8tD4cYsX3pwhJ6KkSy7Q9fGNBb/0AVSYxYksu1FW80vqo2HyMBxPc
ehZYI9lzJMVsnxvjyK/bLnnq8aCM6zFTj1jli4yC8jCnZQSiGY1UBwpXkTxfKNN3
9gYW/QDtBqMq7g4J/MwocQ8QmPNzvOQPjGXXos9bz6kwEePlMjG58utwTSDd9GvS
ziEmPAGkKjcAS0zZFZo7izzM/srztmaQCJTKCdrkZHG7ZaryMe6nYOBQJhHTwZ66
BX3oAiJvcIpX/ETqG4dO65ccA332Pxbkv63hKh/11HcJXE/AFGlCgIt0STJuq06W
q4IXmONFQoKYJql8uc/tz/clkfd3kB6H0rsKmjtTlva63EXb/JymuLQn/hMvWLYi
1EN42I1p/DdJqK6fohh3vv/z20QpY9a/uMRjcfQbQ2QkwVZqJtca+5gvAVheQ6Cf
JJQ623Yu1nC/N0lOtMhTklbzo0LoRM6yTna9jjVan+c944X4r2lJw3RW0mENoYjH
UQ0hsGQa4r5vXNoJS4bzjsEuKLpCK6ufoQ2R5Q0pMZ8t1nEGpc1SthyLmOB9TsVs
2aS9rg+wICxi6WQ3CBjhpH9hmFdfnzu5/lNVB5HiukzAxEDoy9fDSziWDRWwsdoZ
S0HCCguEE/0B5dKStGOjqHpRjtAB0k9a0sIlpf4gNYAkn368/xKQidOzgXIjSqCX
SWFPTMoht+0fpdjBoCdQqR9S8fOe4dIRCoyuYSlc+2PqAvAl3+Vv7x0YpX/kM9Wl
blvNC9/B6df4+Kz3zzCgbvVV7zVT0ghm30TiylsuTm6zh4U6fHJrRZ20hQV6CBSY
m5/C5ex8fhEwp8fPrjON+NBPfX2xR9oY6MAq9YvHZgxLzGVxM0ln/19Z0Ve+eAEi
j3L0pczbTxick6WNQlpTd+lmaz/Lh7Jujr0UFYMVt8Zvn8AcLnqHoaA1/WOl+NGV
EAFwIYxA2DNh9xMtbTPw6sd06VSQWZIG+pvKqwKGq22f4p38WtwjEdqWqmaEBNlY
7M2t4eUvIDZqRHy1N5I3itupwjA7IkhNp7lkSNirEfoCVdIcL6j6ErcFF7kTBae5
Xrf0WclbUFW+sIuyIzHssDDJRrhFqZZAe5jVXUUfSkvvViLcoP0kaAgfoIz8Q3hl
CvxSnEdUX6P5k8doh57ON2YK2Aq+iFWmmssIDEjxovobUDfQ6UhLNGQa4s1XZ3H+
RLFkAVbAuT1c68k4rj1XcfLbxpr3ke1kce5jNbpLzVaNcTJS3NEA2KXvVXgHzKJE
J2Rjffp4CWn8iY9pwHELwBvZ8H0PceUbg76hj6/kfS0YX+g9NJHEYnxLdAsf7WMI
Pjl9wXbkeZsEp+VSpapfs/vyyNzfpqCxT8z2JoufQiwwfjIcF47i8RopCeMNbXES
xB9Ayg762DZdIQTNZTTg8ylD92J19o+aRjkaP5lTdMWdCJrkfF6jFaqaZx1e1dO3
zJOXNHa+3dNMkkVr8sU+HU8Z/+DkOJlKsj8PbY9xfg8Ey+spMjPKh6SPVWRyq9yg
wvDeFlNkZ2uNJqmplvAzLlKiKrkg6D9sARm4xnk4mlA7ID+xKUAdqcu+ZcmwnDmw
V2qFsUPAJf370D7bKjd57YOzeYiS8Iv/VXCRCLim/0WEoD8NvErZVkefXHefsmE2
Z8B0O/Kv9nNqh0vCIDN5DSiIWVZhlOh4ZHuoF5pn9ra1rGl9xpkQGFXM7XV+HsAk
G2z3jwohI/Q5A9KuRwll1HeiXPhDM/+zXttwnbKUYC10eT/c2y7PEXS4LSu2wkxx
hTAplQ1tceml19Pb3wDyIdRdyeK1bu70WsGI/l+31jbZwHcRzmjodwlQB5iHO9sW
hXcF9JOallu4x7z55lbxfDbgYeY/kHfiLUR9Rlyu77YKd+5BsdjRZvjgPkIDrmTU
00/HJvDxCkCXmfNf1KPrd68in/IJAMqzd8j2UrEk/57xnqaT92cnY+Om8y1p31m/
57FMswvERWzXlawBCQH24+N+3FPB7Pyiu85rZVrR6JmzK/YH9eWY6q5dHfixhvyt
35u6WhImrO3d7wFbWkJlUbQhka6W+G9Y4/YahmvzHPRW/02/O3/d8zHncU2wD0OR
qx1ZOWHbAn4gcmZBT0nFNK2NDlSymQePYiHoffCLDt2HkT2mpSy1NG7qKckxfxmg
45jcNFeSSIg2uXkZANw8tpjgXqHtr9UZn1wBvLkRfKwEJqipvQfpxCMM1AC8wfA0
Ik3cZTMK8xJHMp8WiYoz2BzcVe7nEXtaPeOc421uy298LEiaM5TdUTLOxhyckGjt
t58Qp62DEYhpsmwtpWO5tsWaJbtqPABLRkBs15tyZmfxMFnV2yUO7a4FxCBzf5ft
kG9qkuwlCFT0xaRD1EqRpt3m8wjdczMJA9dwv2TtsgQXQ0CgBElyLMBLPxmX0icH
bAfrYYAs4wCD+MKePYWzf/vV6thlKwHiWAAWv7YY+AwyJ3+K2tbJbllDV5y+XNJ2
dGHxQsjXIOhyz1Wpzu07pxSbHhCHsOZ8VUxzTwK8/a0gzH1ra9GBz2WoJTGiUeCw
UwoZwtvgeycqTplqwlYGJ1DZQmKv4wL3HAaV47CkxLDbSn/whRVA4MrkC55j/gfI
oUT2xn9zZRQscDZmfY5t1d5fMSEHPbAgYED4YQfHaWQP928JPmEUJ8mstWrRGDZa
ZNyh4GzE+z3M7BvnasInPhBYb+ca5vdn9XCrfbMc2rb+4wHpeeAPNXATMqfiPsz8
FM8ChObEkEAV/cBaXMzBtNRnphDNGxUa1CrGS4QWE6yLD03zS7vm8O+Yt52jdKFD
GQYrtV5jb/+7N6tAYS2JQ+W1meqb8biw/2+KS0mLVqW6KIwewmlUXps1mnUgnbgh
wmcEA4rMWm7bTIyt/r9VB/coBIys9XSaaUAOooitXLzoGpJVSb8/QLFlevAwM/HJ
tG23CAfPpPHKMBH9Rg2qzZ3T8JkjzL5U2OrfI6rXjoWhdCBiDHSX1GZfWPZorMfD
nZ2qIHTShRAfgri0k8Ryu5CWhCnWUD9Al9TeT8vA+tRXTLttX7IOwnQhb7FFjdEp
zru38Q6EMPqH0y8lD7Te3tBjtge8ulmpAZQUsFoeWO31K6ZoeZHp1UTXGY0PQbl3
5RU8AUyhZfXpkAW9+N562+xTLu+g7HxQJ3dXEMExRST2O6vM1rspwOCIr8uh0jWB
JR54Q5/ZpnvtNZJrGBazpYE6PRekNYb5PojI7groTVva/xlSzSgWKSQEBwgqSirG
vTVkigABoBktSDqtV7cisJ+eYkmCCL0W3TeNMLA9ETvA/vcYnU+iRGUyg2yAHotO
k9Ie21DiRzOurcNZDsD+5DYCWtNlKnkm9tkGyi+uG7fyK9BNpz3t+8PYlXXVyWm0
KGlZNf6SyNEs++lkHO4jHSUAvtWhg5as4Db7gYCB5xmiuAgRrgHOjnmZ64siEn/e
A/eC1dOVZWY6NqDtfXszwL+sQ5WcxifQlVimgf6vwsMMisb3/CPcQW5IWkwlZoLX
OBEA2u4vYfzkPOonJPbp8EeMyCjh9oJCxdndn8IQrrBmzjn4+Lj6sNzyeymqp8Jv
wtYiiyrs/qsIPd/FBRggKKqHbw6bjJQ2gIY8AYZSqa3wppbV3t/rROyQ18axPiEX
E0uC8KaaAioPQmwqkWPHvPnfGmL39791UMmBmdPWnA8WXkszvuv1gAEhhBYOUioz
21Uku6AAwMuHZSi++oGBmVToXWyOwI3h5nJogZhuPpqmavLA1v/ySDJxs1MC+DNy
Sr3yatDoVu25dXeNzDOulOOiE+ubQ8TGVtbSVbS6ZyD6I+1ct6dpz6hl9jLoASPV
cu6VULKRkoJeE1nxRqi72zfYaVZ5bklQFmKIhUXy0a6terPd+peFx6M/g4yATdcL
DnXJjVIKAaSYVNglTvsoHALqqxoAmPtpK6rsZTQvlcnuxMifWGoYyaLLr4ytvaxO
SihmzyQX/ougsvSODJGzIVT9LFCF1jecVLmNGqnIerBAZXq3kip2cY8PKhgWRFGV
zX/EyF6zaP/ZEjDkvoK+w+RHLfSEsqOEsH2GWwsbUEfza4GcV/9E+dJWCqD6zbjD
9MbPz9UkmlQsfAHQgxwDNJ+Izh1XrmBzgPJ5DtjL1hinb/Yk35xhwHz/lj8/hgCg
FTQeOYEo1Xm76JoxNTXv25SqdW1/roYm+JCeOj4XAaEOOwtu6Yt7RDEo/gZuev8q
bZej/F95TJ5ZOIVWgOddIrB9wwC6SrWZf+ZsJEwZ8jI0pJaG8us9WZPh5bKPJObZ
rRbswbtJXtzXkRAakcx/F/KYR7DAGDrSd95pBrjGQL17x57VtZxLqA9BJm929Z6Z
woYtyeMdxkemJIrg4yw/ZmNLAeIPBdq8V4TZ8Fum5omhAXYP/v4AlyhpSkWdE7t9
Fi2QMQXtFKxzTm2W1M2OxEmkU6eCPgocLTk7+J/voLPObcuH+EincXW9Qz0qBVdV
mRJr+30bhoFiW3krwXP/7oVj/KBEFH/Mk68He05IRUCL5ta/ymu6jQTz+E+Wqi6Q
K0FXtKlX3+YohajfqNLEQ13H+3TedtI1JlFWVFHkgIsWKKYQrAQWJy6l4WI4zEVN
nWve2OxbJU0FbCyulpI3F+3JRDZ7OTT3lk49PCEuof+fP7sfoRan6ZsYHXoJOxvy
0SBdYteaPC/jYRVSnCazR+n8EZQjgC/WjuHiHGuKSGtEVz7xGg3dkXY71Xh+Q8d+
beHKt7JSKQiBAB3gElgUrU5ipxmOfcwsmZrSSjr0U+0TGK0Rm1XagL4CZiQVNHnR
7x6NUbL07GoneIwVDkfTq+2Gs9FSVei6g85A7jXPIUsK2TzjzNE7lyZTZbWgWjnc
FRBf9kp8gGB6541fIyQcbfiyuTvtKwCnH8meWC2aGT5f99Z7teqr4c1RfGdTiefa
lF+01nyIToWz57KHMMv78sdFACjemhTf32D6NB5GykwSXCE88kzXykU15JF7aGy/
N3dEEPlZ03lf1qnwmcOh6+Bv+3lzP1p7upEp6r6QnPOFZs9Rh77+prTPPnf7XfKi
qVyjk2djpXp71Vvi71lVXBVRsloFI3yTpiO0L/gXbuLZJOzt6dwYVB2YdzPWHvfZ
mmnC3rt+XJOjfsXnABeGJInPq2z5plUjgYP7Xa2zrVvrcnjI73Wg0wdEKUqg/lPy
VzkqeucG7i3vxrEI5uj8RWb+pmuDibjxjO4IMCBNTbmlYvHRU/9t0bM0r5yx19Ph
S1+8BP7UAeYua0kYj9zZpCbLGFAy4yobL7DWG3HepavxC8D/vZDKV8i+RTWlhzlL
/qyjU83Q0zMMRphVThyCGjxXZsvMSmYletX36RpEFc1HuutKf3R2PG8EMWA4hh2Z
RQIhNvZ1a6qMBGYyDAryOU6bMLdUXN2iFx9Pc8kYkGh4ku7Rg3TLNCcM+akUvy1q
dlsAV48msKONZ4thtGRJq+x4CXZGiwuyUgr0XeouNgo0fIuaHI4vdJ9xfWOt5QoI
c4YUu9bf5xzg0i6AdvWpsrtn+mdIB83ocmf9Wm4fnvsRDZnQBwiAsPSpTEMF//TW
aocDZM+/yyFA9//MTKnZ+yMgjfaqXeugJ2H3DZjWWA4X2vXaMRvPLBnXlkRphSRl
5WWj5wHJfYaAcKkrWyWrdpgvU+uqtzl5wvQxii/H7ZeJQ1dR6OHObb/DoRz+lJQE
L1Wyvegh7n6EJOeNs3GLODfmHAOm6Wf3vdmKIolSwzt/7oV82TmWKOif2cvrkRFQ
UShcxJgpYgb1VZt+2VeuDd8ByhaylbOGwev1tA6XD2BK/e0O9AYoHrJ6/X0A7RSi
hSH098LOSXom8Pn+S/yIcjSlgkJrQVR6CPZxRmAB/r8FW8UIb85Ifo6MtpyrspV0
NBqloWgs0+3hbnUULhHsXbAI0bp85JxQCEAPtbBTyT9ZkZU8SIRDL40wANeD5fKg
z2AwTHFvyJVsqIKbJulUs0wCuBQiKPl9PCigsb7to0wsWoHlSdyr460nJCgFSf+C
Vp74J2FevO0L8zcC98XsLEbcgWxn11P0z8AyqWsgCFySNmeuPGpnsNE2jn3nDkDc
9gJj6vkuLUlC0srl4FQGlxEEceqaBwL3HNonOU6gV9uUpuDM9OLBnHj4X9r5wM6V
jQzDsSkIAgwGmjm1wD509xuOd3QWNvqp0gI523iKkP1QkHL37LqFqqfSiBKPB29g
f1F5FoZlED9+4wJr+jCHqCYpoxdl+kerwO518WgFp4H31ckEYbmSik/243+8qiO1
0Br0MxbjvM3ykJGt7LctVnrTA24/8h9vA9y0RKqMlGkNqKk11K5VxvuLWhXrOJ66
Qxu0WdcSsNHe+liVYA9W4HGWYOy46Tpp1UViZGrg3xjiIJNQeoCovQMSELdqZ7Yi
0h2xKnEssimEBHRDVFDLsdETpvucuArxA8PGuiDediser4iR+UE8tRM8XeeLF7tm
sDLboAButKT8/uuB2jr5IipT5roePlSQ4nE1MBoL/wYVcWWMJP39uQeXyMkTnXkA
nmdHCHuoX0MKvYDErN78w1B/1WXQe/F5fw0/NU4thYyTXEqci5i8kNX/4xi8Ol1z
hBm45Kwk9HHPdviVzRSqMFLgqCyJQW7rv3ZIveDY10MOObQcvoX+znTNq+3H8OSg
8r7JeQOTpRCY1wfNyLcClzFhbKbw1RrWxCheyNNGn8aXXZAETKXJffCx55Ftc1IL
teG48qnTvn0/wuN0JIyPpIzoNrEu6MMKKVvaiZfZj+DiaNJbReimhDdeM+eEQFgS
UMgsKKN/FyGN0+65fdqhhvb3vIT/BHlqoJtiz411S0xMFD+m6whM5R+ORaGLje5M
2rPbuoRgsMrJ11vekvqVAfAp+ozlkDe74FFWtAsnt0IZwEBsv6X0uYrdtaDJbp73
yZLJHwQmdGJhbj0k/9y2r8CJbZzpky6RlyrrEhE9oUHXW+C4kRVqLz4r/SSC95lW
eja+S79gukYPfgnzVZ9ProXuKRFUb2Dz1xRzHjjMcWcW+Bg7Mb1leEoLFPhJjwd1
HPlTm6jfeIpuFckMwpX9f/WeInZ3w7PLr0Bq56OVEztfQmwOH8SoMr67y0vDljgI
nxHmS0znu7fLN24YPi/o+pcwDZiorNXJrmRxWv3heblGhlKCjJXL79ddcGTVgTH6
sMc0JSSf5ArpU2amgN08bLVFzhOEuoITOlu4nFNwK+gZ3U6GE9JewMpbIlfMhIRu
QOVVsXOZbekaOV0xvWcwOvna+4D08VXXmcJfpzUzlJb1ZjRYmKYA2d44F3QuCZyt
VrfTm0cVq3//naLQK4sv3CWQIFv1fJS+zUHRNn+DLqLZnvrsUMvb/XVv2vO2EFbe
eGv7JjHjoxwS5M09P9uaKXrY/TNss2Sy+fo+MLagw28AdidkaR9ROZ/cmrXAnz71
x8uURSY/EtXo6waBLvunjdDTWyGp6h+u9rP/KJfrHVcjUDajMR/5ABLaMtav1938
+nbAAavauNyaMiUGWVqXC3gBO7GXrlZqD7EUlaBtLTJMYu3Vhe5Tv+vJVkdCxjcx
zhtOJT2V2WODHE6rCX2TyCHmpGvdhh6bPxpSlEIHQgMtJvE2iAup6SaRTyFHwYiu
7YJg8ydyOCoVm5Q43NO+vXYxXgRvZr/pt28jqKIeC//6rnXLVCiEQWGyIW15jE/T
urtrEpVxNm2vyV9+DO/jYt2vLAepMgfKuPDtshl45m4mMHsE6OSluCVGZWN6+XPS
YbR+XbyxQytgGRPx7ZXBDFFg3BWbpt6QF9dxRW3hQLSLUg2Gs45lJP5UqGiWUiOd
LlKS97UYxHOK8VDa0Xhfg5wffylflTKDRv7Rbl2b1IINcV1MpoLpUtj7XNyCuYr+
D0BsXFmN63eF1lJGuPEu7LtAa6aDE6xa5ZQmwsPVyAJPK4/Wy5w0VyYfgmDpI9+h
h2iyZYe8aE0MRzpAkDrLaAWspLpl0re+iKFpv6lsA0kH+097j0Yq9zymNB8ORX8F
eCieOLn2KtgKLFQQbGsBV+7U5bdURhF+jp/moxtk+fhPTHf8MmImvhViZxbNNV+Y
bXpbW1DK/vNE7lzdgB1CWjpkZwXRtTtZvB0G5Lid1Nll9JCHHO/16RscH2lVuhpe
RrQkHsT+uCA2oBfsRV18yWZT8jxmXN2IuDg5Gg8GPPrgHmqESr5UxnlSKabAQRUg
UBJHxBNfd048laAxOit5Q9I/SwYRyXcIbXKXLhIW3zVK3OrnWLOgXJDPayEdHRh6
3lx4XFs4e4wGvuIvjXly1FzzW6JY5HvQlSX+tqZM946CcuE9Kase9YzEcpuUORvT
WV3iA4x79Qz0Rt1KQhgxTYGI8DX78UdwChau0/gUCu2x3+LJ55onzBbbGuMwYviQ
M38Wa6VyHkgNu5e3IkWZY4EDxWqL3+G28FVXyp3VXoYX6rFE46rdWY7c/j8GZkuD
4unj5eoBzfySl1aqyK7soGky2325pliDIBrzE8gLQL6qlj7dycuEz+W4IYF6U0lQ
Un7oY2IBPaNBoYK565SYxeKI+xjvqqEWEYpSkEBGbI0d3Xxm5cLy/NLUzhq1OAjn
dbJRb6G6hcp25DN9f+GWilYboimsOXQxLVhA+CmyZIcS+QTSWmDVZGi2+HRqrwly
JInsI1enUT7ZT2j50ebifvP22+D818Edd122AJCOeUeiXvVtxE5qNQRWkrGodIHP
kiw2A6kWdehHhlNo6mIMzpsuYCXZsLbmoC1FcBN8unWJlEOnDGn1uqn1E7PASvGC
AyaRPuJ6DcWJQL6MCDiv2DF5BegxKiSax/LbJOwEx08B/VXV4Erwkp+Du4bmYCEq
i8JAK1x/+D6wIuHgsn64gDU6GW1CtY7oQ/ctrFc6+UiHti1LIbhA2F2m5AP3aZxA
o0UI/r8NivRV0NBwHhdIfH33XeIERYQOGfW+D8vMew2E2eSyBlVF/V08WnemzT4H
0fB8dj91CV7+c9D6xPVWmKn4CJfVmQ3lAX0TQpFlXlkPDZXSXIocUEEFWcWPq2Gp
sAS6rSSfv2WsJGYikfI2D4c2NfeKXjAsv+ON0dZ+ldXV2gQqR0PyLbwUnqwC2Dl7
FKSvN/J9AP+s0KVQjXAizNzsUBOUZtJ2GoNvqGCPsPN2jlX7/IctauTRgbefa4S7
ZNcQgD5vUF/vu3euqdouzq2vMIdTtwuVH8/GT9hwyqTesPkgbHUyqq9N+TDnfSEQ
8SgTZskbMkZL9RKqQYM2Aj+mN++g8qi1zK+T/IfRwEtfQIWEsCq45E6nviMpquC4
BbQrUiGg688P6D1e/kRRsoaLQpu2GjdyEHtH227XUtzuHygOpR74dZIjwF2gKgoJ
FmuK+92e4+lhHjD6ORFj0Nw7l3XXIAkdcnNMZKPNu7Fx96Ac9qZxEsH69RMUlCZA
HSMJwYgVEYsDBWBhSmM5c4mXrCUtqiKvvWYKfcH0e9Ct41cPPHNYE3//EeVVMghK
8jyWJ/NF2dLFZwfHZC5fyKsS7hdYTej1rxbs+lCxmvqWZdTCuFmCiy9ImHcRzFSU
JpvoaQuT6Z9AqUgdqlMG10IyCbEYTXdR3ZMm1VNqC0JlSElFsOWJ75YuwUbuTLf5
4+kOVmpDRviuAoLvyGfk1hxKLw2hsA99HcRWZYcKeBLlp+vzgOydiYFgYob4i+wb
W//pQE14GQ4wWs8SRDsniKKmn6bmC5iYz8VIx5zym0LMTRpXRrDj1HyF6RzUmC9+
SbgKPm/R08QBl6BXoHqWV1hv+RYRMs27PqgXgBn0KkLjMSlACUJRAFTbWvyB/UZY
3ymNYif3K7F9i4TjLeROl5uR3hCznetO9Jiumic8Cey0rWEkIEvMEAZhgzogW0q8
M5KFCS2MwtpgELAba3I0G7FgN4javdwl0MzzZmCnznZ9QTU/K5dduFpT0dDmcR8i
XYW1jGGIP3XViRGMAqsrJHcPLYhZv/35pHg2SrmWQA4M1O9nyLlvyBKTuIQbE98j
F4ksrvM2e7jmWKPG6R21AB0i8m71ayYA+konxJ5tJ+J2diX1Farhv2l8hvvUAVUJ
U6pcLXfgHafbEo7Mvso/CUMy6FDHjwFfXAfISpEOPkWMaiKzsDAHdJzqolGwY0yl
WIrdpafRBnTgNgOxaiTziEdljtkllSttclYGEtBp6l9pTjI954V9ODrY21/sijne
AYIOJSkY1khlfOtJ25JIqkCbqa2vlPYh9arnnLQK4GvZ7FekYWzX1jv06dsAoKSY
HIsouAPZxXA6A+AqOx0J+hJ/UF15rOYYRd/vy3s7SGP5cgv8BOfo1VWoqG+mSG8y
lBkTK5e50jTFdE4Jo4LGS+yst0QJMoyzNquNvU6PmVrt2WtoOJ6rAtwTSmXHuxEW
hNrKc9jr7nuyy9Dld2968mSvJSeXjjHlhkCXMQww9y4gzEALfhOgnVw5VspNq4yn
/u950AM4MsOkPB55JfbxnDQRksNW6rwctz6eqH1XD0/HPFfH0HEwy1i4rYwbjbyz
UO81AZaBc1sKm/6YvD5Cl1gq0bwIz/l4pecPzfbvCihIoDp3CcdlMCOCIkAYUpEr
Vkg40BBxTNVC9D4EB5uAVgykIZwnF2ekxm/8PvutMhHrkJmfCYpCf4v1k5lhE4EJ
LK1VDuFgiaILVbfRWVjaDT23qdDfKXMWIJv7VlddA+Pn7O90eexLGbahK/JsbcZp
8tKsemzb5mjpjHqwwIjUme/wEIu3u1uItGoeVcS7QwssoGO+1j9gaspN5mZPyAeL
frMBDwwb4K15lvBQl1drp4jEdmKmqyCRu2V4DcVwWfwfmXuwVqnvfZporasJMtPM
exvUcjUFDJYagcN9kIYuKZQfDWXQR2Aq08nr8+hq5kEMzrDjwm2WIU4xay/hjrxN
d5luOzwQIcXlzi0PAWOpQVUmIV4DQwmAVT4I3sbZyu9I8C1MRuz8SnZ+c2/vOdzv
6pdNczAEQhA7z9PxYL9S6uGW/5T/N4eWvRYZ/JOIo8oex9kU0zas5ik4L0l02e4k
ovYBveSHjIA1vl1oc90Hu4/C0A3qM8rZ6x1yk13HXzZ38ziuiH3WDCYx40fIjGMK
cKtN27M8RSWQGDjMkm0v+WcjtozCizaufaGCXetRpSzyBvI1I9jKaQgJFlRux5Eu
aCVOUuGV/a/efC83dE/iEw3fuVqTuIg1Tzx+qTPrzjONOwqG6sNNU/AFCPqxPQP+
SvaJgBIu46pw90cUoKc0Zdgm4hf0jJ0m9PWu3GXH9URdreodAhRAn3mdsaCQHV7s
fgxEUgP3rQ3nQ7d0jXzykTFBFF2NeZsMxSahI895CrxcEx9Z7DIpWB1lCd22X2HG
EQGlR9cqeNdb/bjNZWpiQE8dT3nUXAD8Cd8Y5PsHYt0fd/M4+V7JabzbKe1d2Kaq
tPh3Ms6IImenMAbwlIzCG8wEF8ZLlF6yYillAas64ihIc0opSw0ieBWKusUQBARG
ClTVj9oSANiY4NulGRbZ5siGLTidsk1EWiMPEBrqSRSewQUS1SUk6N2rRFaItOY0
Orbhj5bOqw+kv4bpYJbsTR/zKPTIcJTd6OTrnSnIav3mq5ZCI9fJXgP40iqT7qeo
m9XrnMVNSag7sTabsIau+WiYliE3YVL9W+vPZiumPeoZVdHtXN74r4PgR70k3EbF
Jvo7GrUEJukpqGqBGNtlAxcYoKx6lvDlfV9aWAyGGOr2rgMdwsue+gx3S+aqq+xV
cwD4USzu+v/e/WhCPe8lRyRnOJegE/gcB7JERUceanpPTi2vsnlpI5iOCAff7Urw
UCCZXOIK4GJmERowffHuDMOM2/p6coN/DWxolhoQoV47Ayi718sRT4QkO/vqI2sv
w+v2FaOVPrcb8v7eV9JCEYukWhaslkY0fV8hIm/Y3L/ScKfYFBSM7HaSru5jBz05
B31aMhcq5KHX4Vw2kF51yw/GjkVydKF3OABDWGjlaJG23wQdKKpvTan3XZ2c4T9R
WgZjnURUbWBUG0ZeAtauSMIIp+D9CpKjHXLjoIhbWorCY6M+LNdJRSeYGWe/p1rO
zezYvCSGaunYtd1LU24aAGhkVHrYsvYiMTv+Ym+88Scb1mUFNGq5PwYJT10Sbl9N
MPvSvYeMJTcfzUgT0NQvnUtPyBgVkjvleIgBgGJwubUJZLeEi4hyLpAkm9R0+FI3
ysCcJQSPuwb/nE3nhmgpGOifVSBMcUYnOrMG0FqFwe9daIC8UF6y+fOgtrWLCxCD
tQ1wS7KOB4wMoxBvxl1CtKCLWO2wyjFnev4AucWs+51FnsoYiE2Z/9MdvSs+8cly
JoQjPksA/wc85m1HWPDYdvWZ2fMV6S5NCLmFJQ0QcAtPg8w8d1LEJgHq9NDr7BnM
sF6DutqmQDpJMtGwFf90J2ghmLgnOA5M37qz3QNNEu4LvWl3038BxtVC37U4y7vc
y2+DYCeo/SBn+8vq9CKjUtHneqSMcx4PZdT5bYHey0Nmr7d/P3rN6O/kgT35GxQZ
XFdm6MuHXJcOLE8xZZFnOcE/nUyFwTeslaAvZv8j4p0I8yukoPcFHkzA17lo8Eii
xzPGEG4m8P76P4Yl47Hzqm2UtIh7u1d81eiPzYvr7XKPKozV8Z6EnXs80B0hCyBT
bTpjequGvTg7o2JWS2fwYPDhdsNXsNI9qlc576A2e8zPMhKj25INAeLWT0iJHPmT
IX5SDVmVqFPWqiaji0Go+awY7SBQkSWumngblirTVqMH9Hludvk44X7y98igajC/
mm01l/25yK1QSRL99Fsr3Pay4agpBmoE2NG1z9sxTH/48Q54VUtV9jSwuPaWFR7k
aErexsMqVfGJAkgkrpGq2cnDnwi91YMbBFoj2w8tXu50z3mSY3NbVKUH0YUDk56l
N1Lyq11eJ+RcAVDKHONgEnukFOnokxCqXVl3NMWnQiXY1dvnl6IsqwEMQu/PU1D9
SNTo1cJUUiYNgOfyIST9zx1/fTyO9kjsVrdQG5o+My8cty2G8KyMxRTClRCMsqpH
5QlyMqNH7XGlfke/ZyDFc5cZSkZ9S6HKplGlEUWDG1ZDm3ZWq9aiuca5ysOWBhRI
AJTWrG2coqruC0O7HmQV3YkZCKf0fwh9qpg2nPCO+0WmJ15bSunEnRCksIENO0LV
mGZzR0Q3seN4sPjFoBzH8iPQEF+Kk54S0qF8Mdbm2WSoRtABGsO75N3fgxdHrCHM
Jp3O2XRHMZxTWH9KSueat2fOYl3/gfscxpN+k3VcC/PqCzgo77+3mniXeTeGAxFb
QwnNy6oSzt/D92cvVUocbmC1Ttn65E3T7vN8CqDEPow9kDGzv3dhWym6jc4y3cXw
Tdx30GkHXyEGe6uNZLt1E+FbD9fIYr9PADhLF8tZY2CCRZ2C/Qd+X/O0EGOGaBOB
Cm7GplSdkqZ5lNHAWqV4ztUWx6okh+60/skx+OuvZnfMpvwDW0UrDOvKNC8LzK2L
xVA2LQufjFXslyqzUdYj88lPvHFqtXZF4v3QN1wn8M/xGPhDGWjAmL2jo3dKTKHU
N5BPYU/9w6t/NcblCmiIt+DWgjo6BiLzFT7BJfjcc/VT4gCOKUu6JPqp8gCYTozQ
5xOfTu2JubAYiG4GuO6IDLUxPluw2L8E4ooFRTVeOxGhoR/Hp9RsZhwa1l6EIzIt
A5zxntZ4rl/bbVKyPuXjHq7b+PWr1HlkrzNR7vqzIzTsNjUlOKbaI79cfpJUSNQE
dER2a/OxaxWLsZfah38oEjnEnE3vUNXodaMnFkNH0rV9FWreE9/7vx2k/JeM6cAL
WlM8iyHx4aHpaKfAmxCDPIxj4ZrTVEMe5ga0eXNo57lC3TI4Gu3MnQPBJC98jl26
dvcbThdtGCrjJI/+Lu0rG8C53Er3FAjo1qKCmRoKDMg+t5S7EfUVfmeayiavRrYq
Hma5Tl7O148gjjFBGRxqouSKc03FPaI9srWULgms2hqe/OtaLcrF7I2UAc9sv02q
uD7UeSWymxUl4PbEpDY+BIED4vSNoHBRhLsh4jYu9c9tQXYWjaX6MkD7lOIuZxUl
NeGcJcngDZe9uLSiLsGBHGjuliKpNN4utXrgsqs9lysRE8CL/w9XmSXGn73O9mBs
jjesSn/L+1yVff92SkzJpEnCel91Ag6qk41UO8z4gclLY4ouC75lB87TPgqyHknB
d7DVpKIi1v6hkVRc8qhRGGPLLISsbdUAyadvfeJ8M6x7nvob1nCrpdHSO1G6UqcH
A5fdi0Kmbnn8h1jo6LTkdlZwsjS6UXamcrxWohhgTHuWCHEMiCxU8gs0NiwRolX7
Zz7M4Pt7xiNQf5EfGytiatIfl/JTPVkNBtOGMjfhyXc45n0/LdYOfuIxIXJ4Uxc/
`pragma protect end_protected
