// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HfQI9Kao1yi9zNyp9GNYPaRLB5pS1MyVCEs78I0C/PoWvMfoGnJPFURGFWL2AWpE
NjR0JZr+f4veWyXBLQzuaP3QHmpNGAV+V301sgYGZfmfABHYPMqVUS/m0QpKBtTE
FaFDviy0Asgi1wkV++8kaN7bpyqW+GDTq+44kjJ6Aqw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 90224)
gQjcFq0DV84DTC6kTJKv5wE3J96rol8ZC9GruP+7r6jv3+GzmNke+eEh9YzH1fIm
FjP+VEYbVEGUq1NYU3GK3g+t79+fR47S1q6v9tHkevOlqKlxYeStA3SbTp7XtAP0
dU6SH61BTWgGp0s/p4t5g9z1npcqybLajBcvdWE9GAqtHcM9e9ziOI1rQzmFfK7J
BpqOtzHvvsAIQsxCPUrXzkNj1HT6oWczwl9jZlar9F/sW54i9l/lM51J+lu0n3aN
/ONkPSRn48AbLBpzRdKcGVTW66B7+NxRAd1OcAlYRlXbTDDRzp3R5OEEl8J+DSKc
viAL3kW37xv5S2WMxc7d5f1Glf0kVqjQBSCXuQCyGbHeZv3FvIBQimQI/D/6DAFB
M+7WVI0OiW0ZqxrZ4uve+NdL0QmSXSKccUVE3+SSroDBrBjmLLcKfmLanfgXISMy
OaHPqHpl+WewBqLIgcu2LCeYKpI1Os+ge/j22oyz5kerSrV35cb4q5tOCyA9fLCu
mm7Lgz9ceT5Rw+e282XXb3XXuSA46jOpQZhkxNXvAj7qOgqlTvsP2Vp150Ig7JCI
nFlLAJCb5ncDdW+OToD+b2hYFjLurlwIBwk1NIm9fMSS8t52IEEWrp05OZOYlT9q
iveVMFBFXTt2I8KRIeSTJflCNZfwrVqG8M6LFspNMTy1EYJqhEBb5Qu8Ry39eUGP
2Fc6pZc6BLIm8xz2Y0ZaMDlgEPz3IG1YnqJpDvR1pY3cC7X8ICTCrEbRe9yZeEtJ
TPSQads05EK0hV0CTtkvfg19R1mVJ7FxIB9BoERBDrVvyglUd6JcKAspEXJ6YLOG
CTd27Dbrj/YeHIGpfJ97Tq0w3/Vd2l97MEXV9YWG5McCOyNJYfflBHLj8Vtn1MLP
OMBFzTB4WuhHC3uz16rgQVmV4QzK0I+gR4tBQDY86+MGpe14cUuTXF3r5K0PzSYk
CfVbAme/8P2Y1+ZO5qPA/7IYN4DrMFVnw6mkqGhJX9E83ZCZ6B2T8rFtGmcaFB3w
wp9ytY//BK0EErWbKVBhCmV68k5c3JwLoY68yp6otIqxAOuSBLEiTGFsN3JohDYI
LT95lxx6LDvGKm7doCshmESSuEAbYDMvz6BvP/12DlGY+Kd5xo4jZCrZOTC1tyTg
3aDmsvdNApqoL6uhYcZjFD+17UaFi/fVSmdhOQwQS485YgI17alSe/MBA8XYX+VS
ukbW1BMX7Ypky36TAVLBc4HMFnQn+z/ybTc/0JVXZ9xEMbj/3Iv8oOeyhdJv3Mya
nj0Yi6gOzFF/to2gsaVNqm9q4bQU2dSOPX3U8euCTIcX+jhj98Ks4vAHWcyFOY6v
Dp91oUn0KScR7d7UPgXO15QQbXRtD8ga5o8UEMdcUl8fFiHUMsVgTaVGZvj5goRx
IpILBs07eO4RxSXrbFmOwt3cPHrKZSI6E62ez4YyHXeGKHQwM3ZeLahd6FARyg/p
exZRQu4G0GJ6e1/VcMSYcJ6A51po6RjGyxQgtFG0zjQFY6ki5nPCNXSIgm1PpD39
LGG5MGJJFXI8as2efxjqpgRCF+M69TvteJPF59zZpzb2YTFtQSkTTmqgLBcT11Iu
fmPHgEtIcZ2JpHwR56uRLPGsWRWMk+SVslW6bdVbhE+PD0T+/PGs6bhmzC0L/rKG
4T2KUogFyXsgJu6zQzQaXZM+ySR6tel35/g2hmb6XIoxMrV1oc0qV4lTsWPZV4ZN
idGTlPgKwDNVfjBfOXctHPt96457Qz1xDrjex64EnitbsuBRqbE4cn1QEGGCHgJh
P8/jygI20EyOKUD/3rwQo6tFPKivRhj2WpS4irkAjmFAdkx77lFvysAqqG2nJkUn
v+VEJAsJZQdNdkWo19lyNDFWyadaiatfIYoBFoTLWu5RWl06oxUiVaKZ7ZruYyE7
kBeMEWw72e4IbfbOU1cto7mf1BNPp0vcScOYgFmVmuuWRtGwHiwVnIHypcfOc+hn
NyurDDMSr7BhsSiXinCvTYtkAKM7ixh7h8ak9AOMfA1Q6f7ngYzYtXUPebL67DSr
nf/+xsfQHjrpcm4jbSeUuawuBqtOg+l//ZUd8agXTPBcwH1MU1M7pJdP/3eds6yN
uM3aU3X0qg3ggqj6yGMAHw8QaEOYHeE/RE39Vqt2XJKdgeoliYfSC+1MyHQzAH3C
RlmOh+CRKJ6EKaa0XXEVirMeHa8xhbBVHvnqpddGOpadyRq8GpRkwX17eRrr44f/
Hq8LuJ/HcSWesbtW3RdtvhK8QBxVOnqNvivlGA6eHsWQ8LlvHbtFf9xcDVFpeBh0
/FHFfU1FWX4Tyyedq+b78LzPikMjD1uwI4dHXCW3c4QliJ489H/3+i/jJp9zHNQd
ChqGo7fdm/YIBh2wzq6DMZsWHDEHwpuna1gV3T8ShJYf5FWcdXWv9x/65pBAQBh3
OBeLv7C9AuTXqqJwcdtlFTxAmiku4KMVA2Rqni02+IurUzJ9kzddSBVaaKbzAjvi
jF4gCZXAA9gMInGJ8j/FXay5FVVtDJ3aKwa5TjX/d3BJymASkKmVZdeuJ/lt8yQX
KZugbEl30Wu8MbmQOW1hYH3jxPrOUWEJwMixQHueg+5WcVF7ypBLaxsNI87+jsrV
iJi7vwLiQ9Deaxz1JsuhMVvl3f4/G8A/OTjKVXG29o+nbyhXMLF+2CXFk7WHJY3j
9kodTsZ5QLdVr5NsMxsosPXOXBd7cw/bgT6NBV7x0Y4JdS6uSJsplwOhKQ6yhusn
1Mny/sfnxHoCVmNmofu6xlpDMvraRu8oo1sU37fr+8tw+Ahtc2EI94/GUrr+KY5y
53hhIHxap1EJmra/s5S51tyGm6+J76uGCNN02KJdmvTUmHUFVLBEptMM1A12LuW9
QTFYz8XT6Fcs1SFUHRpp7/Tghv9VeAnDKbcBNYp42tERC8r6tE963ovT4+PY2qTO
RR7yrhfQbvPj67TLThO8jMybmhVBvFiSMkfDZkqAmHJOaxp91pVkDhYJd/bN4W7v
470mxGHOp3Wc+xt87bNZ2hhRlLei0FPXvQvThaghIfGrkNKVTBwNGMy+VeojEWTT
KiD6u9ELeRsdU548pI+qch35xtlJrsVo7IKvCT+dw/rp7dUJ7rRsus2Cb3euAlZc
KgwTDTshrvFanH+P9CI5P8GRodKOw3gii5bHHyKhX9t4xSZhQQVdPqBYMjscvcLX
gdOuKfculTB0t9WEf53ZwAsnLggwLocKYdmSBavMaK0fmrWSBKbBR2t/hB71u7RG
8BU4Bb2vUaA54JgnvkmSgS+Gpg9QmW13UPNTLfE73wCX4hTxbVtN0pfhZaV+Uva1
l6Lm+oMkhoSTkq2s6cKL7/hzlHfej/tI52LREUy3ZEVLQuFRr2EPDQdhlmFpPOUy
t79FYkZpIVPbtBbWHuw/dMEI204273+bYjJ4Mdq5upBxlKLevj1alopaEi4PN7Ix
3nV2gy/+NDZGrBnCG+fKE+ZbfPG8xumLX+O48d7D5hf3/bSxoMwXKOf5FgkvZBNa
ejOl2bgWR66a1jqo9afeeGShuV2jrGsMRS7Ga9eL/nVOnU+xMBL7jW7bpkQWAqm5
38JCH3jNAw0suhD/3LQWbNVhop65hWweGaRT5DxzoVP+Cvil+/XGO+jjp/mdlD+v
CnGYYJtBvrIDIZ0NXTHkZajhqgAsym1eIB+3eFdi76XxaQrDK2j2ooxWW0d9Ht5K
lXgt0Zbas/OvVFPNhpdQrEi7d1aADDrkBlili4rBnTb7Rk3+fqn1dbbpzBt7gKkX
uxVJH5pE0di/hEq/4O2TNLQGmVsttpnqlSqGKG4miEID3hYT2HkP2CT68OFwqcB9
80gwxCOw7YsDLi9IbkWO6fQPY/HI83NwJguyspxy8O9AXjHwt+e52oBhi7YNzFvl
MHCIgGMusRl334N+pnsOG9D/0lYAGfNvYpSTZwkwV62OdUv8DYJaHxpoEQHoeIaA
jA88hQBYzvVT+aNuX+Pcb/ocJVqAY17m3edfi90NPMmnXMgKU8BZ9+hGQvhpd+U+
nblulaAN1LD0eU8QqvXpAV5rQTMwtyUX2J0t1aKaGhVnRg+C8wQmBLkq8noL13kV
1qb9ZuTg47wvbanR5THWRr2ZZG+tcv/YTj7j4k3fdPmlLUQ6SkzTBn6gDiFrInab
L7c5bDPuZ5/inGxj5jEsF2JCVMmT5XBAtL/01LixywPqSRhEDupNWpFz5joHRR/9
3E6wXXQo3LHOo3PKEt7aYGtaKbkwAqtiW1aujFLICMWR/0eM2Fxf/maTLuytr7N7
BYUCAyx46rJHME16ekpGHS3EQ0LEE/E8vzuY3K653tRUNO+UlZKm3Y0/TDfj0rGb
Q8lt5vyohC+1n7RpINpEksR6EOeGboBBgnGtnZNcSqW5flXWxUSMHaX7n41eXqoH
FnU4QfrQBmkGFFEHvVuae2iEK1CeiKBtuhbNZLxLq2cf03kR6jVXUgPAbcOe/WHy
U6QXF20THAezfQEnOc90KrRTVpOLHFfyENUWSpz/WbMQenehjrbwvwz9i3aJ+GVg
gUUO4kfBiuRROPFF4ytGBQyJKw9o0GZVED3q51J19XJGwlPC3/D9cXHZdq+uMwiZ
9xN/fJqnrkzDBVFdt+XbFMHdMADmrH/mAX2TpquZsWjddUtp9V1DsqQIPIuS31XH
uDlbTAhMHUaj/BWwfoq1K3zL1FzFyuhO4PoBVf0BEuk93yYwSqbV1RvHeuBeyVJL
jXnFkecgK2muVb7ZFrPt2t1j3VpOHxUyF2VHExa+mYtK76egecoNRIw8j+8g18o7
2CTrH1RlFc734AUG/hxsjvv+RpDauEOKpawpcEtWfFxwgRJpC44LbIwMo3vykPz8
pPbAWEHJhAbc8nlf8mAPNHhIMxXoeXr7CwLfODgfWRmMcLKdW9GBS36rPkckIBm9
1+32mPzhJ1HzUhyrvdE5zfzJHaaIpzv1kY/6OWcpGWH1EpEj3xLsozFhcDQLKLRN
qvCf9CcKxakzCRGBfUeR7HTUl6CTvXGgTqhZB3k/+cmEkg+SLUOpeUhqS2oW2cp+
jkuwFDA69bgE4nerhCWeEB8lLmPDU/+P60ruAg6VnCfif+78wSdFOJXehtP6Ehxx
Ea3F3u4SHCni6RA3n4RPQiw0hQSJi36r9gmix1SF+HOuRGIdrS8UzVGDCZ92AFXY
88fXeolfaid7oxk9I2zI388d4NTYsUGJLwmrIRbMiB/JwZueRsfDYqhadplSCF2l
2JJH4CS4MkODFS2XK8NCPyhqcAr4hK/sjIs1L2u7ceo0WRy6rX9BsiUQzYp2FmJJ
GZTEskpli+S79HYRdChqETEByy7AfP/w7oGURlc4ALCYewgpFo4Vttfrt+3Swocd
aKllgSQiUWNloyTa1Yz1qAgSmP6cPoRD7PAhm4fsshuuGzmiAbXIUyvDYt9XqXgj
squVETVUA6WBAjy3GKxHe+5+NPCwjciqQhHtUZOanuPlbYbqBjfD63vMdYUtGJTe
7nwqnYzZIqbH0BBt37HzALu5HppvKaxQBEfAdyhNZt1yvE1eKTLdDM29YRk0G/5a
8+SmPWeEzSaMSwTkJaiVzPqCJImL7hfZf08fJAoOjli8vWs7vwxM4QTlXay04lqf
w8W1MiC8B+QSU7EWhdx2iNVupWsvbHkPIwDmXiMHie2+8VLHdz/upNxxIxGxNRZ9
h/pS1CrY7irx1Cwr7/iJwjTgHeWOMq+E6R23VPaE+NeaSX4AIiue7+R1UZC2xA7D
yeIPRUNnazMvgQtl9JIGfNpEYMbP40r99dC2M2L9gLq1V+sTWYDYLJDLpO+aUb2b
R1LwTvvu1NfbqTW+4pirCFN7sD2tbnazwWjocwPTiVKgWXouKhGQl54VOogK1igZ
zZfFx2a8/VvX892TSR2ncahTIZvxDyZi3jkYuRuGzXavj5yA0BkgUyMP9blwG59v
+dSO3E7BKjbHnFrtoZ2N5etPE6gCbud2xA74c/ADbSvy5dSqSw682xUfWkXb8dwY
xkvoe+fWeRVy4faHaeD5hOu0jBmknJ7ePR21BDYp48Zlfc2u4fQ3snHroW6GQ2yf
ktn+JmSFIgsRRRf8qMffH+O9ES74bAaarOzM6F2Vq3Q4vA30rLgIFHLH1x8HNNbA
I9acldLc2r8fMyXCe0v9oEfnFG4+Y+vL9Iqh+5Y2pk2DUKG+q3hFJG8C/xJwtk3W
hoxJCwdh803CdwaVLewyt0xIUh+HBiY/71nVvVAHO0N9RHsmFgXAslpE0YGOI1tJ
wJXvDhfrxxuuzV9aOTsCekcphSN3kecDuL+IWl93/9kuzCCr9QlWqwZlM3vjAgzO
KBCYPi2ehJvfYjy6BJuQD5NfNA2rFtXZU1XXd0Iyjs4ZMaktLeV2w4CicrysCX5Y
uS5rU7piST2v7rotAN9RsIUymdxzaMMAdByRmSnqu5EixreH9ntaGXHioVvk7Oey
6H7FAnm0JN5luCMzxaQhiI8jInV95P4Xo5bmWgLlxehXJJBcZNwF7tHiKPkPoPiY
zGedmbJDrGDvS5D/D3tnwGfjT5krNjxEB800QwgQPN0ojSbo3tis1jtC7VyBcurt
kKuBSt5SJY2i0K2jEWNIlDRoBA9meuHpNdE/76lPM1N1dE/Fsek7oZeS5myJMXUB
KxRnQvLkBAGreeVU1AFt9JDJkkFGCKNoOkmkWbxirxUahGjVgyewplRpuGoSOmsG
RIn/OznZUC0lMTAAyxta/4dKSQUdZ1T3iKXRn4kohNGcwxB3+d35a/NTe/HXkXrm
cmUjFR678KkfHa+W8e7ZKMTv+Jn1ecnZBiPdhAAVhGdfdIlNqrn8Z+m/Ive65QkP
b4fSg5Le/FSST3HwIwy/sCt1d9kFjh0J9D/ROdtGVGwQDeHRqgwU8gGzLOkSIsXS
Q8nC4zSRsoTwdSs8fCSVHmNRsa/7t3EIUObpLHIU+jtRHDN2AtaBGSmnoTgWtJeD
p5ZP5JWqNQd80V03rP33gDkkAgpvLzjw1hRpmHwoZMPR7DoG1f2142cAWqj1RQtO
0fmCtgAdndTUs4gdfxUX9Vuwz0PU/QwPuM2ws6FFt8/OE+jzItpxndZyHsbOVPWG
30riGDfd60uOK9Zgxw8pWsk5cyBFdI1zILX36+W2DCC2BN3R5Exwc31A5GAZyFbH
R0M3DNUAfDRi+gSeymEZEbvK6dJkVCvIzOf13Lu7AGhfDX3OkiWNk4hgCfpeQWY0
N/vUkMeP1NvD7O0r6RjVjOE2s49zB78KSCzQJEQ/TQFG4pszzr+E2aB0LWTWi9i9
iVrTjZrKj0CI27JNulMpZJ063s2XIVqNnnNjRqhvbV41IcPg7YN/aMB5Z82/acqn
RqNA+D1r3TftAmLRT6tPbSsWsD7VFqXZWJPrzomr5xASuRoEFwuNoZWOOcMGC2LS
pCn3LJ0V/uxet2cidzQx3R2H0TbSdAUOqJWGBaCldn697T/Hm8ZJQ+Ry3QFWtEFs
bS82IO52+QXHYzfE+2pSD5KI2/UyzzZo1hWqsa5/SLheqPI8ZJpmHI+GwqHRVcJc
cslKvYdXpOaNd2RPW3mG65gELg1kcBo1Q97wdGDmEiHDgzHg5aPO/0aFMB05ll6r
b/evNC5Cir2XXYWUlokEg1nrrsb4h9zrN0XpLPWEFt+vgZzsgYo9+GFngzNewWFe
dNxzISO3OZoUV7hSsGuYwINc4M/FXtCUZ7tW31Wv85At08DmX4I9KSXlOkL/B0tt
M8D5Q1NwXzzSvgXf38SfVWgOK41Mkb0MvlrgHfFJJO9+CCokL1bLwxKXhJuTPtP+
nT8CgQ6MTYaN2syCFW7TGXfZABW1/Gb4nhaYXyyeY7ox3M3GceCWb/1UCsho6FPI
t+b/KQ/ZpYzmyJw4Y+hWzc7Z57dPT6YXJnx0dnLRkyBZVVmldTreCE7+fVA2D/ma
Ufiuz9ME2POwkrFabvsUfd2NilP4Y4z8aAQ19hPVM9JYumrxzLJEkM4EmV3uXjep
V0r9G9MCDUrcQZF9pOtXsX1Y8NobQmoSZbQ5gjpVpc4t54Pamb5xvoVynz3f249l
zFlj956EPVatqktyqyJsiI6S/QX/UmCsS6kZ6lCIifMjKGci83Hkb22H+NcZA4aH
unpMX1c5/RaW2vafbgac0cReRT/CdE8PSeSlI/4+qcxHnMtERmFYaMYHv4JNCrRh
FI2oj8p9iSOlUxzdQw/Y0HdVMoByFewx4xXgeVfzXg6HJWBvXsyXh5iwm/6634US
RNNR7TqlMqX2dIB39gmyoXX3NcZKE0ZCaZ56d1jdeiCxr9lhVEYKp0Yuhdn6nvKW
L896fYetVcdaVEMW7gMLC7hNAJ6HIqbq4cmr7gq9o5MKySeMfqUq4DYnmccyK/XO
DzDC+hcsBuN42cLkyewkYgIEfingB6W4+2dNOqjvtvh2qhBaDlUM5VcbGbArDKxo
d9fZig2R0APyM5fNGbxwsaroJEU5nxUN8i9IZHrVp7r8eG1HwDMge7vLyP+1TGa2
MAiVmSjE0iXPwjMrHdUkgXVVB22HHqiKqWo/yBklSoM9waMmFfDB3/GRDQweZI5c
2omhDBbOmP1XmHCrN9+OCmTMojJeN/jI1RpCh9sgYR7zFlhio5oyBDTSTfixKgUs
WpfMmqn8/HVZenU7Yj752HE8AnnNk1eHE+W3Rs8uomtQtq/8aQK1ooATF9plwT2c
MVIXAuZ/g34UB6EWO7m7fOyXVAswFpYMJH929Xvx3hUZpW6+aVIYkNoleJrklokS
Nf8GV9N5GqaAZ81LiL3OeLvdsd6/RGjlwmvhWPBTADkz5ZMUhSgT53lxudTHTpc5
Ws3CTLNa7Bt5LOVsDFNh5iYzXEtqFIyvl1ZUmsThPD97hG/wdAIrkp5k+Aq3x4K3
zK8PxC0gIhmVh77C405zwyGQIkoZdAmhIjL3tJ/o5Ys9JIG0Rj92+YBmWsvGQfPt
/LrW9SiSgUVvMV7A6L+i5Aw+wswsEU4kfcWCjQwoiO24u4XmXjRZZEJv9MRuzb/g
2JrIDPpMSTrZh4szefjN00W8n6W2ovWqMBnzjGM6zx1ekR5np7tKFQ7ZEYiOaAGz
e/CuBnc/jxDNEsDWbCuV0sD+B/aG6BkSjjGhSzKSLPR4Ak/GEfIMwzWPHyIDN6W1
QmnWX6k4LoIXFVu6V8OMhsaLRoItz/f6oMdJaC56zhFMlnb2upFc7oFHPXYSEB2f
yGPy5j7Wcd/Z+G3Q1U387/uqpgp9sznb2HCpfIURnLWpzORFLEtojMsO/OZLaH9d
/5S2Hc7IOWsKjyYnGAUGyvThAgw7swR3RzRXJxKmW6lHArmnOeu4FMXj3jNnu4dY
wiTHo1/6Zxs9qsocz4UYDrKXEOsdTeYmWFsPHfmV8XF62hja8U7/T2HAeKxCxECW
r8i6o/9642GNWxF5zPvcy9k75hp60a1Ki3PM1z0k0qa6SzwA4FZBNewZBM/nORiV
HHdEig3kLuyutxhE64SI0SfpDAol9x72p4dZ5vWCAHJCYRjK5XdlQvTv3VviVV4c
qFbjcKQpKy2VMCi6zmez/6BVSigm+RMBP4Sft8DYj8WHXx7fX5GX39rUtT3wxcpQ
xvCMst9rCCnU+V4DqwxXDv34DNcKsw49Q3phZouO7JtwWU+3gZgPFu6ZeVWPBHUH
X0eJMFvMrcahshBTfMo2n87/ZnMCV1Bk7ZSTXanAzHyLy0YT9RJetlGbCfzdpUR8
mTpStLWWEsGSuZmxY3bc/hF3XZONHCxrrOJbeL75JUOIwMwIR9Mui1umVFmL4A1M
3ADd2DCZrjG2yEz8QcmVSqTx/fLdPOxsLwfE30agQlbO5ZC6GNeMhOnivjGmIUwR
lq7bc9uHo6/JGVvL01cX59xsDhMp1X3RH4fHMbBD7O2th4VUP1D8zEmyP7R9ti0M
PcQfy2gsRk6Yqyeus0T9rBhfqiL0OggHeVbc2Qw2uKsEOzusBLXqXylqL7QLbmg1
M3MjLFixSsyGxyeruph7dB3BcGh5qrro44JiYoKZZABHZytCksam2xGg5DkMm4Zh
Z6p1nWJMQ0M1YN4AxD8HLqjJOgCoO3KaXfFTXLS2sbhDNfAnP9Nvk4oZ/L53prK9
WjTaiEzIGaisHRIPK1pE+AXgLt69ZgwxGjucNdRA34rw8y/EVpGmNGFPalF+ht9p
dV9eQanDG43UBc3nr4cLr4eClWznhlnv+sqHHdXp6OTVva09khyOT6PXbFy8gDZX
2joRhNOIBrFArvcEPNuzSPgHQz8VNulYul4KQwGQXocGYrSzP3az5fvozxTCXdO1
OYo7xbU2TU1Yrnjh7LV8s80HBupMH+BweGGNS150yqC6bJ8XSpln8uL0ip2jp/Ft
NvhnkZfQXqVgRDAxYsTgsSZtjUFbeUYhf94ZV/qWMDlytvMNAoYO3SR+BN+0vgSe
6RYggDtwXwSDM7rdhUPNMagEiAiWwgpwZqj6IBawOIX7hhNAYIalqWyWop1OkskW
Dl+ySfKLPXeYvw8lZgoUmrsQgCnVWXkPzrBJVzNU5ngP9PcDqOKMhtrl+N8Om8jN
cem/h4TMcw0pvVb9zeVPzqfI+hPLtHP2XApN6cPALhDbuEZ1YFqGTD8zxaCEpYOo
NGsqk80zbRgm8W313QrAPKTVnFEaGw22cKElkCbDqctSmuCRyhaY9GelPgQ7gQoK
3Zn0vxmeIDWcT183l4kwJ8NTsU9/h68g8O8bROmoh+AUYdDRZrRCbQij+QIWFByN
M0KM886PXYs0raN2X20KOJkyXj+Qt4JDnZnq/E8DwjhB7lW2+1goatIVQEmUJBlm
g3rhK9Xd3LdcabobK/o4c7BTmUZgu+h62J1yOe/fuOVdfqRWK/maPURWOOiutc71
20I2XBe+Cwbyr66BVcvvp2uyatqVblbeJV3m5VEPm6XJUr9ro/3Z/gBynZWG69J9
bF3J4pCrgifyjPb4taGp6pPtHYsLJEj5UsVZIjJniOAR7WfAQcN11R4jfxZLuFc/
c7z8LcrbP8hFACmtR+/nyq2ZSUUgL7hVROfUleYiRUYsaK8PzgZcp5suggAWNkFx
yMtzWBoBVwXZGE6ZRl2pe3+YPatFLszBKOP/gQupqETwGwGoyI7TgEXxwuZlkyjm
4RuC46LkFWydze28YvKW+63RFdFOQIx7lQzrB8O0kfqNHL43ATX1iQWMgb88bHE0
eSIRGjZtTba+EuKzcD0QspKfE/mdmtsybpeGO7g+ImvIEjymQJP24ase+gV7iXmY
hz+YXrcisNYhe5ke92qgGJXOCThMenx1YjAzjbOk9k7kd5I0lPzGImPBX8jJgywh
/8haTEcWRlIndln8i/YamN5edwK2GQKk36vk7r3PjlB1ve2BTT//CAgKbPsVNxok
Hy14rewXcw9zn5pwXeaqvu6Dg3rxOkE594EL1VlmQa2Th1HGLivzAlwU50Rkktpl
KIgy3Uwnid0Teh54FHKrFniDNo7u1ISB/ZqrZQFot0HAGnciToe3PmWCg9Maq7md
LjhL84X1FILZYHXf6jt3wCwf2mfyoBvfu89u28BiB0245WaltZXTNGhz9SOyzj7B
jUbtKpo0xxSo7FT6K9RE9gDNqAwU7rTaogCnyt4zelqERxmUpV5g11ibk2ZVxptX
Vc2wWUPHDyPlx+MD3pKJf/l8B0P1dNiSei97hSA51COlm54Aq7CDa+19vAa53zWC
Hj3B1LqFNsQ1Vlb1HqPA0hlVh8qLgv4FJ0AlFJHv+jxBl5jDjdU0j/C5l6SJs0jM
sb0gQ2gN7N3LMpFopEMkQC+45Gw4WpzCiCc7xZQB4TEVD1irVEwyVw+aTT73KOk9
Wq2I9ni2SHwaeDG+CBZ8JHh1MZzOI+44VziiD5aR/W8jJuCC8VIW0OuNXkDxocPw
NxSgMafIZN0yF4y13t1tlS3SoOjom1CaHpqW0xEfuI09Yh7WQfenOy7Jdq/jgm+E
mu2V948rlAM7s2LNtDaqGHOXhQzz2KUZWgGghuQkkX5SlNeJ7L8rdtExqoGG9Eaq
YauepKlQ2scrBOGy540fBG6i264Hgjmn6hDGHvdMeTgv/csR8f5ZzQFaeSeqkov6
Mh7zYXcVib8XSd8nNAOsl9EZg7qTcQ1QRvYXT8kP7zb908K7z7zAV172TO7i+smK
RUX7woKCJxdPi3wMcmvWTphR55KhmrHwZSeKplUlhOQ86B0PlbDkZ1XiprF1I1Gi
skz+AeZsUCgWIawNM/37gIreuQpvlgmu00Yw33ECCbiKm3nHz02flSXA0bboOVcA
jfk695Gzt9+TxNaV9DE2xJL7dLuq5TDkVkifWMZs91YLbZOm1wic1sKXzEf4b6En
XNKwO7iZNelw0bcood1MxKmb5TwiPxcVOaU3yWqQaQpd3C76Pp6KuZpNwF522eOC
pKLoi32GMACnvZ8zo6Dnbviwuq43lGbAEQ4+hTuJ0OlbW2hHJWwFt64ZxRhB21R3
s6pBlYNf92/7Q83gVdbtgbMmKoQkx9XEdcCOb1rWgig5YBXiFD4UJYA8TtTQX9vb
7P+5BJWmtyoRSbOVbR5ph5RjuUBZF89/X632emLtCNI8YZ6qTP9qy/bQuUKthstb
nVzRLm/z1YeJUvnzNiSoN+1GwE1NaDJ0/YbcmkaTJWX8NtCcQSvfvj+U8TNq3ysC
RkKRAGJakkDsE5i8xPDeBrVffgdUV7zhrL0sOpwaA9X8RT69+IJMIUJOKtqVBMyT
fUjl92o/5KE/7b/WbcPFRCwKthmlLFud6+VPVVXQmkxdJcFYDvrui6DtUlp0m6ZL
4cJi6mMcTgclklhah4aWOxTtE22p8PfVdpLIE8kIEfK8tJqr6s5LOy6HdMXb5B6o
Ds2ulpbHg8RAzMhhk6csxxmxZKalCY0JSEQCIXDwEQ9ZwcgFLD9FbfwUHXXwmMC/
faT0y8EiH2VRt8cET+Guyra+uuH3dYA7lBfj64DrymlmFQhvpa2uoPbs+FXnMylS
uxlpE9Uz3OrIL0QiQMjyOiJedi7v8EVVG9A5Zi7mI9Ia7gTCAEEspfl8HJ1Ha/5u
JkydQWeoJL9I/DxRjoZeGp5J/JHi9lyx3w4zt9bXLttMvn0mQIdT3ySMq7NwwQSj
zUb0lzCpBAw4rxMDShXeK5Ru28oYFs+JC2iHiZSWokl2DG7vzc0cQLNrrkKsl8Bf
hoWGst/6E7gMf5pZT/4/6HhZ1lE7CDmU8Q/WljVNCei3oneuTGzGxLWlbRXA8CAe
vflVgUuCFSsQXYKw/QVoH7Yxs72znS+HhPqsYS1q3309IRyJW/NBxoUOcijWrSzX
g7+ZsAJOoDi/+dyas+x6zCvOdxN6WjR5yoNiUgetTzryMyLAs/G3k35emyF55UoZ
TQHesjTaGnJxad0PB1OiFBgzCAl02fpIITaIxHb8u6JXWq6URh5xKylVOAKzyP13
W90l+gpXXtewbG9HcNc66Fz8w1HlN82sze9bJR2DL4YKXRRl8ZSHqQhruUgA2bYX
pQk8v+a63FXdCMgIQXtm3uykw7YZJUn+udGlsmeVY4L/5XwMN4SkMnfYgX7aLHNR
MxJptFtx9szYWPJ90h28Ndbl9t28wQvr77aTorUkrJjldlPAzBTt57xdeNf1z/YG
lBTdre0P7CTYddsuRamVR3F0/TlOTQTitkjtUeSR5l4RBEEBlWv9rACeRz3ljfdk
kTDwDD42hIRyil6k923dH2K3khoqrTR83tnFR4fAueFarSuRHw7lqjEHgKLq3mm3
JpUvcwZ4QiAQzORjOq76sXWJxRwC26QKKrJAx46oRAvEEYJ+PYqxQI3LJVf3OZq/
hVR7GlmvrnzT4CrAp4kcgbbWhx3icb7ApcxBPc2mAcTHCNxIYdxbypuc/fSv+UHW
zMcD+chnU6Ow+FtfcvuQbhW+MYKquO0f/rpUYDLRRPuS4T3aeVrQ81tjIX01mBTu
KrpqoYePW+K5VE2Nnl1SV2gEvTcQUxKNoGmM6m/YFKO/eglrGYgdUebFflDfMzei
1aZivBCSOfb25+VgUqFfl1vzpTFt7aM3YiU7kf8pFXZTggtZQJb0Wn7yMey2LI6l
0dMv6/s/N0oPADEQnafclfjloE2fTFjkq50D81BePzhJRMQ2t1ODiOQlMgLfXjFy
acj+SNcmNtRSutfPphVgi23nqIH89eRSya+AeIRzN54CzsYe0p5Ex49RYYTkwx/c
+ov68kBeqpXoqzpDsaCIPKQVt0YKa1tsgJx9ZPDk/1tEQyWh0Qhl2xHGBdIaQXhM
lKKYTLXGzVX1OuKD01ffSn+BQeFlSIcbNIhwPZ9j0gKVOlPD2GsxMOIVi/qAg55C
mjde3shXqGOEpIpJ4YSL1665NRY/H01V30gSrJfufjUVVsBx+sRzmjSyNOw/5GUn
CfegDf+KMJA7zxhhKC50bZKUEiyOQLHsnfUJI0kXRJeAFI+Drfyay/v29wzZ5vVE
oy7JreVCacxcB8X6EuagbP0SOpYzYUUuPZPcMvEDrnEEJ9lgQCgwXCEZG2y26ifA
Vn35pyKmPprt7E/In+uhfkKLLaL0HwXMvKk17/rPk2NCA4npmIAy7gBQ62tekzK0
7Y1kD2A+pjUEYFCp9IfE1af58eOfhug3ZqYWKgYOIWbZhQH6fvTECDLn18eQuPdr
MkfywPSwFrqWBzdYW6nuC83wPvpjtxZyy9TVzuswNFarLsddPPYsVOq0hNWX9P6O
pbTiybLZeGcSh7IpSo7ioBFGO/lc3GmSz48sh9rPeGp6alPHIT39Qzw6atyHT8Kd
JAcYdO5pS38jkyh0Z7N6PSblsuEsPRAr5YgynkFl12jStpSHPq2/vvW1Asb5b9pV
7pR5Y748CrGExBbGrO+lM5KfXhDXoePfYmNLQH7BGwMA2+4B4fQZYMO/Shx+BFLL
GZASYOa+acY/ls7NiX8HbD6mjvUhP8r9MfCBOyquNUbXQo3ArVRUKolj720M8FYZ
v5wb+SRUcX61T2//PibJUTSuLPcAIYYr+fEzT+AxzpPKV58nPaJF61U3v2uyQR7p
RUdW7FVjDU1SYNQL7wCJLvWyFsWRShZtzM/z4vJys3sMSSH8fmFCdvPCiW9Ge37a
m65/YqoWCMy6GlfIb/Bhb6cpsKXQXYgxCC2aNIvIv/SGOPeMIrO1/ds5ntpm4jsf
t7ejGZVKN/p7rzg1lHz0DQz0bhI6HqGwXhc2DT16xTtqnBhyz+7RBO0y3l/1rX0q
uWWNdxZlf8op4CGgs/vKRDhp52dPzY91eafhfl5V2uCvrlO1js6INc7FVyGBlUA8
bXnzH2ki0aQ0HSsKrKPHN2jf0dYQlQILXyF4uCfVwJGkAMHlQW1huWKQPBDlAu0c
eTsraHQ0hnafioYZR2zR2T4x1FSgchFAHJkVl1xjvoijn5K4ZqiLdp5fjU2gHE1w
uR5ya495XEaA07rl5GjDQoDJ6yxr7mj7jLQydHdFWYbj1X+Am1KN4AhfSAgyxKNd
K9i/+ALVt5s5KZFJcMdgJQ0xd1J5xanuafVqBqBFjJATA76WYVss6/r3lym4ZnYG
qi6kTIodThSiHLZZcO3uDQFLS00Y93/Jqhur3FyGvYxJIsRG3YAC56p8g626Qicv
5KFnTome+Cq6TlYxuNcKZp6EF8re6mrAyfjbCc5tzfM0HpAhCQVvQx6mQXLD1K7p
aZEnQXmUtUZ4epS2DLDmuFgzAOAIBroDItAqjCjkiKOMkPSD2v56ekfiZXV85hcY
zVRB3P+B0rKv575fHDdP3V2OOc1tysMS8WfkLG/hyc+O/9nRvWkoNWGoWufZBEg3
6dNfpdvQRL1qwgop3HKJiGcrTxZq1Qdsh+XJhaWmyryB8Th55e9v/TE5HfXYQLa6
clRNfwtjBOTo13ZV3/XvyD7GQ1ksff8pmeZJTdloQKY9pFKI0O11bdxdICWSR7CQ
PvqBFbfYqV4acJ0XhQnDWJmf5EsQz29T6svI3Ga75kmmSILirfv725qpZwUFr3XC
Luw2Fpq0CEsSvu/7Z1rTWnd6/93xvt4iR/jd6b6zrU4Ysg3y25qPqHULH6D3xCF5
7rECVShHtFyoqVnZApsQQTeJv3Up7je3FDna1RsdEJ7PomrwrNfUP4kC7oNXbuAw
oEbVakdxh8tHL1q8sTBLeEwYXmLMZgfhGefHqbFWVs8ua6dbj473zS6dXZqKGUwN
KOBA2IxN40G+vDld4XsgdK5FaEChmwQT44R/mmYRFCCBdcPVyoLLsP0xbc3gr0UJ
f8dBtN+uW5JXHVPS24+yAKK0OYG70izG8tK74bHGRrUx3XzVQUrZifuskJlcm/zg
N3I2txa2u1N/d396roYHWdL4mTwqa3ff2GFcK5RrUzBkH2pypfN3KCn6BAFsgfm0
UUcdWG1wxzLDsdg+b5/52FFWD3nbaqv9HgF2IQdnSZQQAohCt0lh25Pe6OA6Fhwv
t8XAMEtEJRZuNkjoA64UWEwRrXdbBBbfVd5+NiZwYRIB0d7f+BrImAuFWDwS5w0a
ezfJCX0kX1WlqGwlMCLik55NpQCdRo+hWexuJcBMza/Ogbvb+WHLHiGkpU3+YT0j
09qLFuMdVvHdgOs+jWhQk8hF+WXKEaQeNi8gxb1wzA56uhzn5oMLOP1r5EiYg9uB
/7mBcJ9vVgbP13vHgIPNayGKoCd2jzxfT+DBuVObwlLve89BppTHod5MgGAcXOB9
hJO8zMi+PYoSQhjBCKwxAvU7PHdGVGuJc05q9QRjiN1AnWuWNYWNVboHrB9HdokJ
U/sxMLtEaJss2QNezeebEPWAAQROUGtzv/X2BdvpHBr2iARtWsvFV4iNjmiR5L8K
YdsMu5Vng/snH6UdIfCaSXLLzuFQvB9UTFkSkQbmzAWdISoOqVIqUuu6wzV6JilG
D9G2Skogy5ID+Cp5qH1HhY4xghJ7v3TMY4PEq3puH1aVjm3sA7iuCTBmdGAWL6Cy
O1EIW+cHVHNayQ8wO7IKsy43bmMBz/Yc9XT/3nCUmmDCA7Q5oF4abYjP48YQnlf7
610AWa6KUC5WNGeU73YJ6GJu2LeKWucAiCIWyL6itlElgOzJzUU/FkTJXYSxJvkK
uG7O4joiYW+3p5BEtAtieqvY8+HXa7dIAj97yocgA+uA9BoytmhR0YBCGRck78di
OE7f3jtJOIyNS4NVysQ+Nf0dGSs2kL6M5d2fFFcC8P5apeQ2Q4+9ifAJrwjpWIsL
unUVV9JFu2c/2Iuzm/jge+dPEUTNdFkMDbsnO/d9D9yfbf64zSo77XOglV9l5zJl
wWNuusumfYNmm2ee2XM1OE0RR+x0y62G+HRQ59trPr4NUAKf+wq5dpRAJYL3AuMI
S7xpc4OLVk0A0qBHS0oBBAuMLEOAw56ztg7SNIhVMI4NP+vlCqWNIBJIudB5jvzW
E/sldLdHpNZPOSLxi3ZJrBcfrkqk3RXvEHOFAvKNuWXkBYgj6PzcGIbm8CVOjGPQ
NPOF6alvz6xN1Ln84BqzN4cJ9ZoKoOLfTBX37n7iaOjPXYnyArxEYCAV1SRs/mfv
XGAcpAcUNEDCObphtezC2RInKvvnthJV51emVLf+OpQlvpYyiej2znQCOwTDKDxL
O1JW+Vrrbr3Fy6rSjvmWvfs1dhfucgVVcta/I8dyFxZV/UWSvnpmuBQfJjuRJDQG
EU64wDPx/o6cFQTcqsIdfhOaEGAPeJg5wgI5sD0oqaMEPG80c+DcXTPzWTrbr06Z
j2cBkkVQHomDggVYkTO/So/pQjQh3+7rMbkVbU1O1K+IhZifgylqrI3LGsMzNaXA
XVkgIOxMXH9mfwFB1nE8nKN0sH0h6tc33XsZxZ74uyMPewLaymMhArWmZnCnMo6C
Zqdp/ia7iQuf0XJ/7iigq0N9swfjeJiQ3vAdrrtY2qHjK5oDZ7ex7BPDvQiDvvsk
sfq9yBWXHV+sax09CEOnZoQjhhL6J3NV4/8bTrDpLcAPL+A7xMN8Mtt+6vZOG43U
zOojWk59/GwYPBflpSaXCRkixI1QwQxCwXoGQNnH0Nx9atqYYMmWB/vtNG3FD5xO
d/TJ2xTDOTFSorWNJsQb7hV+dPBqt+y26CxmS+pBKpksj3TsGOnhK+doOZxmvZ7M
H4pediqIB3A1iLcDqO4sRy+rcyZNS2id8xyg2t+E5FQCm6vfHhObCSdDquaU8ct5
D4fGh+DpxTM+AkJ6anmEjXF3MjhYQUW//mFBDFJkSoTmjCfBRUuqkc7XT/k9owlG
Y8G+/WE45pdt4DhzHWouL9LCn73cjz/+g/9Oz9fAobqXko6GNJLfSLghlq5FHbB6
hhRH2OeROK2LYd+q0OVdD6czmeVonNSuNbetB0XNgjSooilL5y7Ul9QSLjd3Zsgv
abC2wnSEy4BCtZpXPkWEeQ2xCuh8Ig423DzUMNw8xm1b+PT9tCcYT799Dfe/8WGW
i3tOsgX9MwcyZXsYOBHQMQmKga/tMc6sGO9gtZmx4p9tZb3NNX3AjF+X28+M+N80
pefp+pa3hFk4ORw5BRzz3tNpNpiQEDvWOm7iMABcyNJfYNqZVF36wlP9rI5aAzH8
W0byv7dj3mdsqa5hmoW5QeF+Ys/saY+Q+gccJGt19GlTSSFkZciKFlc6TPjJDkZp
xGhtn0haSoqp1Gp6BmxIbp2M7/EII4+1U1L12u5j8YVgOgBKd+ZqIkRLeVGohTdL
OF5krL5lGKu+Eq4ZmHSH1OnlSZX18vf5f+XssxCTg3hsroovkHyo2LfmBG8RQ8ya
KUZbGa1irzrewU9bm0KXaZAtnaMlXA1ZG/r1FGqv+NwaQHCFGoWcEbau/WjvqYOH
ugnFEgDFIsYKYYRY6K3sa9qfrTzjStsDDASW7F6ZQ2SIXwiTDQu0KJNyrYpSC9tL
6beEFsaZR3M6a2QZ53P5+ugmUCGYHNgLHh9WLlFG9Oi8uzw2aT87plhxk3w1S3Yn
DlI7K+Ulz/ONiTM8nvEBC/vBL2yXt5yqABRixeZFVaYnhDW3pEUZRUl5ybdWhb1f
0wjYsVrirykpsh6CSDQYzz36oX1zRSB73pCozXMAPgstxI5hOOZ2/J8l3Xg5Xazf
JZQt9l7FkyYhMMLO0tomA2DA2CDypVXNCLFL+6nCAf3YB+pyRg7Hd4jisQFVrybm
Qkzb/kokNP2WshxI0rdYWrWptyc8XFE82m3WdYmPZkiVvRYu8NV9kEkeWmMp6XQr
BRxq5xqQTrHMFNkeyvUqa16eBLehGfQ/8Hz00ZM9PBpFR2qFVv10jHj3bhyR3189
OoAh5h9KgSOGy5qs70GLIwMA1Phulizq6ALC7CgLnu9gQ56mgW3w7+hD2eFkJQTX
QVZxR+gGG3C48IIK/sH/m5XAyswZzfpPUGCddjEtOCzFPfgmsAtVWuARHqITa2s0
Ot/4b4HFzH/KrolBNDcqjIPATxKWJTRV//x2SBkHeMTy9u4WkiznKZyPGgcVXTVr
R7CR9buorB6ZOPbn9pdlZ5uDOuai02ul8sxKPMtkqkNGs9DQwnmnxQ/GDMGlT8eH
xhsrNs1u8eImoPS94N/ACr290CAydfShT+GqIWzsbHQspgD/AKVASF/DGVdDLx2C
vwLSw9zCHhV8n8/IW658GS1zyIJs5J2Ss/ZXf8/CFG+/J+2uy+syJ610IKCr3+2h
wtBu/pSqiqURug+t+t/EgifGc058bKXujZbNJQSko+AC1FDPANTyvhoCzognXJYg
FqSryj3sHqa/0xHmjdaEboERFe7DPhUcYi4eY3tjQ6DUWfJdvefx7p8MSYhKv0cR
A30QMmmp9SUOkUPvKrF3Ad+qMJfuDstSmiSbxUaNvLmkhpkj/7VHwTP8XSCQkLFy
kMKUPVd2k4NeQPkciti9pQ6PM48bMEVE5Bk8Jamme5mo0TsRllyeTBEkMaqDH82M
kuxyscz3CFy0bo5BPLKA6hyQ/mdH9+aGrDguzA349yF7aS+Svkj5EvLN1vKL9RhE
j5Qa2upzOXFcqRgnazJf1K8XJsyMOYDtb6pDZ0cQlwHutHxlYerLPgYbghHTPgNP
OTQEzmqURLb1KIVZVdxrebyFiWIM2QI5Sgdbs+daw2vltInGcJwQ82qILn1w9up7
cOwT04dTBl6GzfGId5kdZTPWM3ZDnx7fMGkmFEwPtfg49ocSEw16PVQiHjhIQGwX
zt6RRXIe2vc1RfUVIbzvaU1n9fFp6ssHKL9IYom+gZ3IzgOnzhnt/kXUXz/rTgtH
tA/iTXjmtppzNUu7T2qMeHMWUSYPIxfOkjf5pJU+Zc7TKUk+kS9hjLBUf4Po+4yY
CvYePcdXkJROobtizHG2sDs76HEhCt9q9ZSKIjZIgjcD39fZtarrk+uEJgj6VZ3T
vAY4nWGw6SMxkTjif2CtLC6ooadkZgpcKaDahsF8VoWvwWp3WpKNKnd6kmS6J9fp
GWno0ZpRkOEEGm2wDQQSROLVKaaj8jFC7iwaKtx9HjZhLJQgJkEzb0iEDNRqrnwo
hSDIMRhyd7i2gyZxSh0QMHIy1o3fgHuDby12WxW4z9C+2paFBUJeDYIGCoygfrCJ
DPT2Dr7N0Ct7ZiVsYKkbDWrem5XO/D8cFX5Ga9dSOxFNi5LvdCX+cdHeh9VKFsdk
EYfZaxtTyl/DA1I5PIuM38v0OTVFZvsmaFHDE5Gp6HzgJvNqnUeHiVYNHkCBxnNt
/4C2ji5T56ztEdcX8zxBQXmTczRlMmub8wUbbQgFYLaK6SrjiBoLcOJYrN0S8ZHk
AFX+fslHyWtiaaJ0xh4TXp4Mm0jo8oEqAtXE7MrTFDJrTiMv4Z9wtoW0VdDSKETa
vbMw8L+6SEEsRzuv0+CLW6sY8ov1mIcHpYmtpdhG4TRzINYjrTCFIIDLsBS5L70d
T6PR+yA5cyzfNI9qEAM7sefw/ds2k88NNtpjv8VoI0dTJQK7WI6yea5x5OPT0f+c
SpgpaQVG1ChwIyHWRlVCJXxTswoQY2Vls28nuvRff48avr1wwKacZBrke0zBVDsj
fSny7yC1JB4tPkV7pr5o9y3qLnXiiSF2j3L+wti/tZygHxZwK8KaPV8lVojhtNNB
6LTnfTiFK1yoedh2P+mG5ciZjF67DmI14b7RlfJc0bdbibesWYsfrqJT2cQ3AK0K
44AqChxEPJ++T73RKGu8ubrk8elata6JLH1PK0qKM+23CaARqImJuOsZ22ZxTVT+
w9uVzhud0uOJwDyMkV893P9p9TVo45S9anOqWVgcHkE66HiaM2/FTo2zWLOVqzpm
ckoNrXpkjzdFrpRG91A3jPcLwSVzhpuMRMYBGtx424dp9g4Q7i5vGvZrELBcvdpt
hXi3iduYiXSw0YZ9JG5GXplUbZGt6J3o+dd7AMS9qNoUmGCUMGd4P6n8eYyFQn2M
e4W6KDxph5aVWz52d8WGcOmmEhK9lUoxz0SDTXbatazoRX+8g66mZc5Dv8BIOH/r
DOaI6X8jjlgdvlPW7pvdDMPjmczLtYit/jI+5HZFOR+qy9sYF9liWagidbt9RwYK
5RIhpR+M6sCzZOAl5wk3WZ5kJWZLLfHnHA88RN2JhNPRORwe4xnL5uRAws1wwTow
FHT0MxwNinuirTepMu69DnNyUCglgeM6CVywfnsW5YlaMURK6T6Uu8pSsrdtd/AJ
A97Q5XYzaU/Y6rsb/Svp0pVtmj3HslZHcAXe01ga934BhFff4ssz7JarR+jYf/LZ
rD4A4ECfjK0KazfJIDWdZR5AQILz4kdIAngFAS9jqnJ4+18kKq1kD9esw5krSpl5
Tp9815+8ob1BIaDT+5U8giSxPG1SSuagGH6kmSxiLklwRoSchcCjWXzM5QVjCXbL
EuJDDgeUoadsPlE7x259Y8JS8JLdyJXLv6LNKCqjOm2A/tkRITWD7ziZSufJE84B
sw08gKOaODzQrYsnQvWUuk5DkT9g7ozZgiSvonJW1OrIPpY37GVq49mcYH05zSC/
mVNzyYb9qTpEW86B60Qzv5ZuTf/XWKk+TI+RLYYhNNLozNzpXQqCM5vr5WYw/uL6
+yqHssvJp0DOqDzT1JEQngKttJnqEhmA8h5n9NEXYoDm1sh08wKAJ0xhZr6ma7H6
SlMjGvNCNUbbGOh0CPoSX/KavI+NfTJlJoDovRFbLgTtVOcbQAsWhJGj7M4oC9KX
5hDoUiGaaQ8TLgIvd6SZjqhztUJhU6RejmokHZiypkoAXIMSN3DsHH9MW6apnb1t
W6D5uVwIWfwm88ugK1yd9LA0l24hqHkR/lT/SC1qsoln/w3uZO80NhQsqja4G0q/
gUZu/3YL6224ANluW1Y5bt9NHeAqoOEuWZ2vG/tFnqm0H1nuOt2FHTL0N7GDYB81
JKZ9Rdr6UWcAzQDC1aZS6GWv2pNRC3Gxe/DGWjP9yMFIFEwT2mhO3SWWHyvKvdyp
1HzC5owZIt/EWEfOCGmGavfYO29nX/GCx9pF86Yn+MCw/WSzBcePbmcsf+LvGALn
C+P6YDOYFkD3SFpf7D1s05bH5uA+e36/WoX4L9O2GmAWB76KRhd30qtYZKtHQyOr
/nEGmqUpWSVi++tKl01eGD7YXmTLyinBIj6nwBRDyhDd2O+3lWJ3PdfbIninnEIZ
0KInc7h9v6PypG9qNDKZFSiGgZoWuHtvFHp/E+m2EeXYWRR3XZOAGCteNHCT7SZx
rZb8v+TYT1Qbu8kqUlqhXDRx1+y/i9cg/1vplfI1fp6GLwvcAO7Rvr1pwyy+/wEa
OPHLjpQw5cheOYEkW/ewRkc60cW6Cg34NejaKB24qNyAonGsAIDthR9W+Wn4rhiC
+PT36LJPz/8RU1Kttzp9Ya6xB8vSemOHpL45R7FNEp1w/D9njhNJCWkP0J5OaxXp
QA5ef1JBrQUxv47b5NMTQBPx/c8pvOAIu+CoSErCHV1/gUvDrCePsfnejWSjeHN8
0F58tYKarMyx48m7XQlB32c6D2ZN+oSHhGsE4oYTxjafo8u2r7/5Ew2oI0d6UOlF
Y1hC/853v15p3jZ48TUANBGv1ar77hrHjq9oiw1BjLQNQLgK3y7kh6ab4mm6txX7
kg/yljT6dW+7C5e5aLbbk8p4QEHSan0fpRfmWjCkwUxTBuI6l03t2OvFnCSJoib+
uMMVQWvOy9dXSZUc7I3A5gAVQu+0vgyPVlYtOMajImMkHxHHTESsNGi+8WVG4Wrh
Euk0X0fs7h6mvP7RQMIb9vne+hCi8Lj2ygm+toaCR3SjAzrUDNSX+7Dh5p6GG4WD
o44YeXf/1Y6kvnsSjTfw52Fs80yLAZ+y3qfcjpPJRrvBOSSEMtrBQhWLl91/hr5T
J8z2euwG2vxxcujUOAxmLs1upwKcwJkeYnOzQ6O9J2fbPQ1w7MmpWcopX51oL2iA
t4yUCN5E9fbMQo6crBCOfFYosqZepSCGuJ+6X4n3NlgyzVA6T3ROUiQKZhBNMaBK
oR+MnxZB84s4yIiUPdEF6oz/t4fqJN0ElSN3vCw3nGouvXKTmRn5LCRPhxS5k5xD
eJHDIOlNO/GqD99DbzesiuxyXUvopk5tomf3Ibn2RJwNVSsVaU8OwzI/uqdUWbg6
2nR1k0VtGD9/pSn6HnDv/xus8JgzkEYtkHqQd4XqDkPHJqxEKgn6eaMUeq7Fiu7H
3dapOeFAaaR5ke5dqYmBrJ6QNGmC50mjkgv9Zj7rh9n1AZFi7yzRJ4xEoFwbo5WZ
Vzfj25DUNPDhlXYnyMHz0oKELUWM8dIRgTgfe8wWxNiSGSPI7wxKH1YgXWLEX/bV
g/6Nej1g5YDzUuL7bKsf8xojPvn3uf3w3AgzduoDp20eVcdmtgonf/HJksCUAo3P
zE/AmJD4iiHqIuCEChm9iMKsocZfKwyGUmHow+t7s43wtVYgdWrCIKnryuN6CXRv
Mmk6s8PHyEMCAArWKGA681oy54/WG4CEEPeuE6waK0Ob5LAN5e+xeRxR8kNkFSDZ
NeugAnPd7UAldA0CmPM2uRQ81yaDJVPuQ1oRydFnCq7nrC44EqANcUWxcV1aweWY
LB2Hp7P82UO8bpuG3zrQ/ml4RzWq0IFRswq5ZRcWcmctjx2hoSpskW2c9TxfEaxa
2eNuKsBUY/DaplAhVp9e7y1AMHDTaAL4f0wNtJmgE+AecWCQu4xpL4kmINaeerug
DR9Nm5RyfTGMHqq0JjCPGbFx/HPe8zq6rP13UcPq4mE+661niw69mMW2UnXZrmXh
qiDITGjQVmRJZk6cre5+OR4twIJmJxRtd6RyCIGWHqKzHUn9pLoFjJYUld9FzXBN
u4GIGUkxIYAZoY06lVMHw5hY/ne1yFlZ1FgBGmh3tLjR0Pj0RwRzjhyNAQYVXf90
FKEIH2MajvKHRkKnAzJZvgkqRbk4ePUmWzBU8P+Pmzcn0oXxyrdJgRnuloEDfVPS
/+HowDkv5AfBwo9w9xnibfTri2QF02H9GCJzGFQQdi5Bmb90GGoQR1JKKFYl+KQT
smA/+v9euff2Yx7R4vhJCJWMOhGKFxec2e4p8K4poGdpJx1iGyv3+NTKv5JFwLbX
+PfRTt1gXymt/ANUfnLzOc7g5v6kDZ6ik7NbpLqw7NHeqAl2f0ksG3EMy925OwYC
f3bUhIeZhtOr6mlfPKlnB6VxhL0oC0dXW0C9yJO52eN3DPYlx3fvfoQrV/dZSmaG
DiLNdlfpDZAolWZ3jLQZFtmOtwswiBIjIzVdmAj857YOiCLGL6n2Hdy+y74tG6Pw
JaRMa+lPShy2PUL4shGkoYkLoGTvUm1+YKbx5c2YhOMEph0TaScIZDngyqhM03Y1
UkQ517TPtQanmxOewxyPaEpWTdlGvjFshLbEG14nP6ArVTuhq9j5wpAl6DtYcSmk
bHD5qCZKuupHbXSBs4ijMfK8GvkNCXixAjs1p+z0DgujQuAf0Z2xpxZHGRtECJY3
3RDdqqW4pJhzkwkWJpp1Z9TGW4IPpOwM9jOGsbFqw8NyGLCVcIm1y+g/7crO6CoJ
WiA3CS+A2cik9I1XOHeR9YqriyD57dsaJKcKny1SAjzGZRVMEdVws2vIYZK/68up
iAy2d9phqjZ879bROOux3YePFFSTlPOhSSBkaHtm9YJEU32MW908MMqPk7iwevI4
b2KdLQyI7HKysDJQeohhmgsIKDbHk6J03avWDwJFV6FWnB6ot/o5Dixu0nuxG80h
yDNTeO7YUEJMBpbapdyNAoo/GYs9Lizz640igt6yBdtP5PFnTFuK7b5VBBgOm8Oc
DYlant/PHQ2U7gNi87ovQSfA4PeifxzoXbX/NXBDEFZsXCKz9AdfIcXvrt1nXpp7
3fx+IAj4Ah6sfB7gpQHPvnKr273I3FXz/85lb7e7/3oSINjN4TERg8YBMFqIQhHi
AxQS5uWBJvy9dyMpzPtye44veYZ/hs0pQ1gQVMGvhaoTvTpUF54UqYu5InxBCzgT
93FvInatBfPlqFhTTWcdpQWLSbdFM+mpNzXXWmI2t4UdX4QsZolIWCvcefH66O/l
ErVy2wbd/Cq7Vpu4W3I2jz/cUJtsmQ0//P7gjItaLNWLK+OF9JviBRaYhL3NVslW
ozbYQ17Cy66tmy1KvwrYHpPtJ8mVSLTKb/3Wk+hL8N3VZNLV57/tkUs+I/XlsmNb
yBA/C/0GOse3ehAkzZzk2MBoS0C2UZl5qjtP6pc4VMH/s6y9KdAB45+v2czrO/+p
pWUlOtAU16z5/lYUiAc0S2QAZSu8/iQKnWymBz7n0QB0WJLkRdaziMjyCfOPX3EQ
gk/hxzGDkJlZeA74wuNIuuT/nZQwOZtTJhPGUmskGVZd2Jh62/qxurFyf1IEZ7QH
GlaMlvKT47eaU8jtMuHr61YWdJjrU8s658adAjSINzGd19OQDu7DoOomFKbStCbo
W3Gn7uowrz+EdaB9VXsZe8UpxJWcOrf0ujyAZJgOsyuRtNSO+K9WsAIlmnQlw1/o
VmKSH/doWsHAkuuxpcYO2dm+oSdZAUzwPpj9AxgSiIXn9xbRPqh1ti+lU+myUYUV
oUEuiOsgzF0Iw7XnSSR9mZczx9GR9e6MSBB4/kb0Bpiv/ytN+3WB2SB1MkmQaOlY
TpD+3M93gtGxed7BsrohgRy+z7xmw6ldFsHid3TFTpmYikO4TKxc3TBRN1yVc4gp
vjmDyg90uBa5EindSBKEdN1IqRmmzKXdxERrD4w6ZS8FRyLFY/r0EpDuEbd06kJ4
ISyKtHSNdSsOaGANY226mYLJyNBrh9aSQQ8hlJDObKv1HWbdlKqOoh4t/vDd9EbW
TkE6pxpNnoyKdJl7q7I6B+jk7NYY1Nk63oiXd/eoW9h+sjyia4+VFWAmkXIQYbrZ
o4jAypv98hjq8pSw9TE5yH+WRvs5vGhIQ8GiH5pucQ4bXYhAkH+9Nr+gEDcdmPTe
rr3e74INqZCwUuLfWH2DlY+j5Xit+pyym5AOEOLY/IHOekn1VtwiyFWWowUUuuXg
xUwt1O5C8tS9ST4LM/6pguzVMN86oYJUGxknfmdIk6cqRgt1c7ujIrk8ncvOH/KP
GdPeE0WWh3R1cCDRiyC1OYFDsAvDNSS9zhw1scEwgR1ovEkconqOV0JxeaZZ54go
AwtGtHURyjj1DXv6+RwnLmnwEE7iPTD6r0GfTsQahvId8wwTdHt7K31nw9Oc5mjq
22WV8rX8RjHYIM136xBvWlcsEIKrTnR87ogquObUuBKt58V+nOqqMCNZnrY65HZ7
DZkd85Ls2fiTkLf5H+2hzqctosxKEaLmRwI0hcZ3ViGhd/LeqZkW4Ddcmzlx3SVd
PlaDVjZyxBU+GUmnNNoe4OIHt6bUmH69PUib6U1sj7NH/OZBFHs+SDSukOCc/eLg
g+bBgL8PfJL5Hy4FbUlWCu/SD4dVcNv3vqh5rmqcRMhUqwiw7N4SDNYh3cF8SrlV
WhJqJ+lDV81u57hMbWHNwLh59icL0b0o5ljcHN1x84f5T4ShCj6CxyPCr1XC+1xB
yEl1BonH1ivQSSVmftC7CsMKA/WeI0kfIDu4Ep9p2IJFX3rkyF1Y4UyYfMODb99q
94pyD5Mq5kOAG2BilAKo4+QlopIBmsXmE+5XLG1zeoYNFUK+gfbNBYIZJ3JGEdlK
sgv03uuplj1GOze+fBvNwN4sT/NKPDtnwpDb+5wRbA+SqKV2ywz0cMUMSQkZ0/+S
MPuKJFRBrzzltiKPZHGsr2FRrYZbCFYVUFbmUk5TGlIWSWvWn6v+5dLG4/0hjgb8
awtAY8h514eESvdprNlUC9I5E11gx0jPuXcWA+6Q7TyYMCtmIqcnMzzzynsfLlAV
+Jn9l4jMRNKQUXOxyY89o5nOo3nBvZFvdzEGFinGlXBm3aj6tq1V13pDICE8MVql
+FbW7R9oLgblWH78ebnCsxfuiL0eHo7HeHOeLmclbnnswpkJZhq8K54/cfficCds
L2C3WUVdyGuEW4EucQAwME1+RUSNmnXy+LQtEHGy4uKN5LrWtg1KvtHsyxAzMG/a
udOF7SDIIaH6q/o5mx4P3ApYRq5r5axJlNAkhNrOdKhCPR7tFHK4sfg8QBDux+fm
TOA6xBQQ8OsnyBWQrZRLVnc9UOlrtQQ5SP0FHvZCVqcz8eK6Sq++Fl2VVLTaADTD
BfadImBa8jbZIinZ9i1rT9cYQ/pTD0mtPHyt95ZfrT7f455YJrWAnMuv+KQTDAgm
dR4ktU0s+muQme3y6N1Pp1NIjwn3AnAPdLPDumFCFffQx9pe0N0NVEqQAjrrUT2l
NhYD8mOeKWwkK0jzceCQAdbk0OA1sIkvTtNnxfU5zC4gHuREarQeYi7BZBPnoP5Q
9Gk9PVd74RXW95gaCSTycUVn4UEQYMjebs9C26W1xotRQlt69RnSBJIGX1i0UF7B
vA3f7aK8hvDWcUMBFwPahTasmthiNT7CpdFY5phUThPhfCPZS6UygLBFSs64h1K1
HW1tvOMfsl6mJ9nWnBzI3E5QWN3w94zaPZQ77UFUh19qRAW8HfxkRn7iRha7/UiW
2u0zeoA7ve9ltuFGM/xyAy9Bd3NCVwwG82TfoPWrjTKabN89SvtjDsWkr7XLYeKG
06LQWigmgjcDQ4/P6Dv5yS5wae2JNj4z/6iHoZKHKkM2D4lcIaOXYC0JPfAeebYB
TbW62fvOIN6BgkYE/cVXFuS7YULIFpd/InTxr93Fj/vdgFthjHJvzE6Y7MrYB72y
p67YVlXBAq/RzUZgtPUeVahkD2umwWFpVv2Xc6CowxNythBfwulVWOP6i0kIfyWe
qrsXJF5D+uO8C0F1+sNOltIZVKg5KPkE7EOK2f5eciYS3QN6seCnsf7bZA63kYyZ
77p4Y98yKfTOWQJtp6NUg6tjFByf0oBAUJYPHebhZouOXFiCJRq6YQtK1pT0R4YF
Okbb8V7vXBE+tk1uXX2rXHektHYStsZjZLkwXOSLmmt5ktX0/+qWiE/aQWfIUt7b
H56m5kWqYmW4mEywnIEmmTg0/qjEeDwzLutPkg4UHPPK9nnb4mcGneooMBZt8I/5
VXzlYN4Hg7hCMq6rRAbCG0Ac5y3mQ2PPWnb+J4qkV2GUyrfZYXMhibHG4CCW5YQ4
cG8HBkRq5jRpNHR3Q2ngXRl+XADRMhLWNgaQUGqI9rV7na17FAcW/nb1eD6dCDFm
sOJuBXRcjtmcsqkzywK1Xt3o6BW1QCGaLE/c3EeFRz6cqxIGeLPxQfCoLssykAbY
K5WR0QvH7JvVuZJuSNtusPMpwSnNhIALd76zz39jGCgIH7L0dQDi9DQiqLwgA+Ib
Blz6VqC2+y665x6n5EpBnptw/KO+UnombzecWcEaIuK3SswsLGXHCnN2YQQ77mX6
S3jkvB4G2EZiWyCw9kyPMa9gsSf/iB0dVucXjVI7J1aTXtYGvCL+ddUjnV0qqQxD
Utt0mniCjr4Csnfe8AJIylS/71Y2FvaMgMSgzvoEBctr9vyEQts9APkdC7h+PG9s
YgQI9nAdoBxx303cOgXelG2+JpTjj2ThoCwI75E3vxY81zrnIRx3FhdmV96UxQk/
zMTBJV33wvW6w/hkyWc2VktD/3ltxXKSP2tBKi/H4IdPe2+gAFviHcf+7aa5RsvB
EAFLvtqsB7+rRhbbcVoAs3GwQcjj4cUaglmrFXReQ5tuHYPX7Lqyi9bIjHDsxzui
XOm6g0VAni3T4fUadQ1KuSEPmwkz4ZmLCP8BPe8pIx6P8WaBnRS02fKnro0wJF2H
vPH3U+FekEWfXM53PB97WvH6wOOtuP2jkGctp4xoHX7kxPkxWV5NCrqwyv3Ys9oz
13OqaZord0hOfbI7dzi/bIipUyq3Yo67oaizYBtjcyLMqsDCb8OwgqgHUrpJxmvb
QG7lQhxljcI7uf4TSI2NIgkzNAZIbxPUBDzpR5qUkcm8AJHd+I4qBe0HLMUnaSOD
/3q+Hd6SRl8I+QJbzNsVL76zto51B3WJ94qoOiNda1RhRxiFfXwoTnb6/SYh2B99
gSxS8to/FABVL/WXnL/ruFXuHRcS6zGn1gu9RHUKbUlXpgZLh77SrXyjqD9+VZEm
FD6AIblUkT6NS/MwwlGObhc4S7eZNhHNV95IIYVlXY6FV4Ec3cWYebEqSGFNlCgj
VHzHXJ19zZom/JaZreSzEPIriizFstBNoGL/emBhzaxb4SCtvdcEnvoYA/9SN/uW
wHmMhaOLE+hPMmqRFpMa2Aj+NEoz3LcSrYlouhxSVdngQHDerLfW85WEOgANsCZt
uPkB8kKQyPXMrpE1QsREUBbYOCf69GsInhq1fgQDns3iFIcIZBk340TVFWnaiuFU
D16CVFp2vt7ojPb7byJRjnH/EGIBCnyeFe0Nv22/rdU4kpYGyF6XdeTuO+fWe2ez
Br6IDb4UEL6FmCvljC7lgizjCpNg8hY/2wGYzAZUrD+NC3skKAUWB8BbjDdk3IJL
YI32mFM7jM8WAuGJwLBIKCG8d9w6QH4gICft4B4pMXdJKriIl1PPP3QJbDef+/qL
4hm++a2lbYVIK6LlaQhDLm3Cszw7pwGxR0Y71eF/mwjN9/8dRRJVC3gPtP0NaVBF
f7WUd/4d8zxkIU8FE9VmT1GfOZAi9eAEsE8LCXtSqIuCDM334Y18ycix0hmTfBkB
+WBix5m8XFdN12aMAx1YEAaittKJD6kwlVpJbK12iX6ijzcLviDx+vGtdO5AWPBa
bqtWnD9LQCFbw5rTKr01gwM0wmUFEQqdDeFbGEQFB/n9phqDaXomxXmLa89UvEEO
6rvsh3kI4g2lXgFPYLdn9KJYGuq1yFoMnY+NM/MRJlfxJtfS9nsZN2wvdevJIb7+
Rhh35/4/gnOMai2/dXhxAxEodkr9gmlZ2GfUGcUwgDD/mApqWxOZ3mvBAU2Akh5M
0Fd92d0erGRYWh+B7XEMwEXHj8jaMIZsA//UgfiDH0+CmmTM/Rl8k0ydrd39ESnN
vZp3mTWMNKn1+m3lFbU4/NFhyYkGtj+heAI7QnXFaIZJkHt+g8avlGr/B5TI+LZO
v36XIddsPQo1stSpDe9yYgJObh9zzhhtcyRd+p/kRKmaJtBwfSanDcJkdFHMUsMi
FpnqNvZ7wBTiItKQzccGEfAz4GZQ+RgnGStqkxRtH34tCB1fWXdOBYXIDa1nbw+D
KxpfDk579JyKTUDyjb1CxUCPKxAtWCUeVSMhtn8o+6e9+gB28U5aR8PUJDLPcD07
r4Y+5JKpVljZIul8MprflNBH8mcMeSo5IjEPMagMOzmqEwLWJAGGOZNtK/KJmw17
WNJqJkhP16u6LBKAWxXMi4XF8Rbe1w5duEIt0sCxwZagUligT2p3eo/o0nIMJBuA
Cz0MUwuWStRIOaptgv+5DBk22nsc4htdk0Medo4SORycZAGQ2tMT2+4lFUvHqeKf
HhFNno6JAn77eZm9IU0iBuTgSk3RnWkl8Yo3HqkkCfWVbu4ZO2S5J8KIk9YMvHKO
IaS8RZunNBFD2k25Xivr32I+bBWPik2NnOBc8VYFceH2cxZSQ+o48JHLKHFqDhsd
a1SE6stdsk3kQrHRmKOLuro1x5igLX1vshqg6mpdPorv2EnBmSTAZ43MHxzsUFv/
jPAuj7bNV6YpKazqaUXDnYl6p5+6jW0RyWmKXXFUJ2cAQlGOkNvLGaxuM9XmUDI2
HLIZ9+8HdatmH8bUFtBp8UtDYeW8hw95xythN33uDM2Kp+g9zdqbKRC9IoPxEZdI
bc8R+X07zAQu2I90FfjXOVDATwSyO7BN1x0XXxqzaymQznZQWDHRCPc6raAcR5IR
zx81DwfuR9CpKapfJ4nLpYHPSd/x3bqm5mbkGLzJT7mLc+qgaKNZhELkxPyP7IW+
0lBUx88eLdkhjOkS/m5QSoT3+Ue9GkmHpLjvC68f94WOTitFzTjBiEMWjszsqHSS
AevXBsM1lhJ6ff/vbnLHFA3teotr1tYCoWev7xRiihFkoomoydQKEZDwsE8/DDyV
QgXQDNXcWHsfmS37ZIuFhyYDVYg2A5At1MjTvzWdq9qLE6KnLhAtNJcGYQuiimIg
PD4q+HZWeqxO3IGLzOR6KPkFFqSr43FdqJJZABNkxVioW5Rv0UKW8k5JWWUWyUAM
pNfZAMA08qEvYLsSkg7t2qrMBkKTvAl6gc4ZF1mXVVaDvvUoVi+7lLmnjGB5ar5X
iaI87eRQWOneIEmzG+IyyABPYKNua2Kefm63CN4IskhzEVgcn1BQdkjZUU77tu9b
j87XwrdYas3/n0SOLLQ34mxKGoXuFoKrVnK6EKVhGv4uKcPG5tBtbFvq/gebpum3
W/z4NxtsLMpCr3oxFqF6J8EVt2OH/NTFq2Etx6+huh6e7Q7Tu+cNcbtvFZqhWoW3
8Hdd2UhsWOGBZCv+EHoMQ7EBKi0zDb3Y27sCzq5wCC6zMs8OrSBoB9MP/jEBboQc
hTWLqpabIcsaLciJcIhN6qBIaqbLdOyMyh8+w4Hoi/K8KoDpIsX72+Du8fwt3ush
9+jz9ehn06tziozUUyH9jAApQO3srlyYOnHPBFbAcOy38UFC+0Bk1kvs3M9LIxI/
pDQUzqUysZE2iThdGPwc98ioS2Rpa2oqL1V+Rd4fTJaTU6bX7ffv/VxNanOoXOmq
wl2gPQG767+ZHElPQDcWmznDYXohMvcXmZmNNt7dK89P+l3+hWB7XdePxLSx5NRW
rK6zjF9KyduGZE0DQCa0AiZy0K4JmdWQ1M7NUWl0FElnv9zuoF7Hk3dCGxt910r5
9SuEaVoBbgNHsVKNso39389VArFlsORigJ6HhvckROjA/l0I9FCLFmIKiufQLp5b
pwypzVAni0CpwTcfg+RI/qrlwjTYbblWEyhZRerfXyf+QAX/bdLUdU8Gv26sa9vS
iQFT0xr6nwHHzxCbRHSCi0Ng73AvwJDDc2XwpYcaMLpVg910/dNBShMFi0O/Iywt
Ny8AF0iTvyZtrh5M2fnvXQzb6k+KluD43hXFHwV5cLVQvUCGPUpvxbK2HZjKMT2R
vuq0wPWVaJETew7KLVGWnFQ9Ci0pZ/JgMYVXElcvNryD4RV02Zbm/QY+9RJO0e/D
kJ9vUnrwYh2FiNzp34SXe/4CY8+oJBig/VTJng2R6+JhY4IPAqwCjjNjGzfK1heU
xQIz86OpNyAdiTzTNLS95KHGGXVV+ZSkhV6tSXHtyuFh1re5dzplu6UbObSzwSTb
OMCPMFwWWMq1QJx9+cb255frWjzFuIhGRngFScSGA2iCSfalF9ze3mRKviNxf1/m
JTVJ7aUF4cJkB1r8Vmn+/T2shgvU2UjqUCOB7j2HTYVuQeH657KiNej8rpPrGG3k
vdiXcI055dGCNIDkHdLd9/7cHIWR30uC445jvkw8aE8aTvwvpIcJLJ+PGcbMaJTh
4kFE9z5NTzbCMBJ7FXqJjdZ07aq7q213aeg3dZFlra3O3VpNxII376LyQrHytHtn
mESY6UX9+bYjdgUNIQnhrhR+RBHMLM6VyC73LfcEO4XzZb0/Wb4kkl3SHemijT2+
dhf7cKDIKct54cM0GJbBl+Zu/oqr3EPqPmxJD+ffHTC6m1/rEKAzDUS5RBjRViW8
U1oniySyPqsSKSBtWapHUr6LAmwdvTk81LMOq2ZvXHR/vJniPzGrWUc3eBAMwEPP
1crjDB3XyrC6ugHuVZApPfET7fAyzYT0kH52vRYfIh53IVUIH4dPqcZ3/zAEs3D7
LU0fgm+jqn4OrLgN3/+cqRje433kpCEE57kOLJoTpile+aJsRqBc9c2keQcTKkTV
fVME0MxDJuglYtDltYzfXYuLN8KpUpSnyYqi/MhMrtP0bwNmYhE5yfLmqHzajess
NwK5xGo0GNbOQvoiyOaaJSi8GRivsaE842i9F5QvF3pMmyzYIFwnv/SxlcmpVrOs
aXuv2prWdz9mu6XIzC8ZsDiI2yqO0v4woDZoPlWN1TxuRRYxFBHwc0pMuUQfYgJl
6g50AGNkhIWqJmJr+p341inh1+bn4l5uw+mY5Uqu0jML+bOR3Y/D2g7aY2gs8QVo
Nqxcq/MRCikA+qBAYxSVycAKeGi87KfDS5JPK2+Rw7Z96NqqCkEWsDSRBG7u9tB0
RBnN9GmCtSf/t17GkEyuhelfLAjCaXVUbjS0lQfGGdTEPxWMkZWp85mg8W8qeNi+
C/kvM6B2bAV//rPncdLzPwgeMBIKFoRkUEGLGq649bIw/xWyFHXFrNpiy6aqONpR
52NUloIHWJyFM6JIQgRXV9eQ9X60xnj5a+WUgY52DBVDMnQqsJgSU0Uf6rYEz+kR
YeRLKVR2+bcSyOhtfaqwLSBtD4IjxerUhVaPdLIND1wbVE6JYdttzMSuG0K/+qmg
O/CfYQwvR+Lva8XxBF4Co9zUuFcoz88lT3eYCUGQiOfn5ahqB/6SDkNpqEayDYxn
UmwwYuEJOMYxYMGqdzJNNx2VzaY7ewae0wmRdhuDlYiz3CDSFr+8eG1Bj9Fpz5oN
gcQDERj7eUgwoRc/HnGykNr2MzXsj6WW54e00bIc+GDwwcXQMrS5PYO0nZudKZmh
necg9vi2ghMo/zPW0GzG1F5pqlHIhqspIPz7NtLiP1TPidnbnRVEdmbD/tw6BceN
nq80Z1MLEOlcqjNUCUwTe7f0B9YumHvkcTZ4tiQh59HEqwwp1+zg2UiG7e0GTgPa
5E5IUNC28Q3YRZng7KLosw4f62F3awKYAHenLojJ5NfznFrBFAXuAotfN1F9CPCG
UDetu0QyJJcXYPtuueI9o7mGK1yQH4ypNzkVhxpbtSlOsfBC2KAJZIT5f4/0gDEE
kfCXg8nIKbv6sleplwBdpr8mrZCZfyt5XzyPFvte4LKuaQD5qOuE6775SNWYbkqU
vTv444M0abC4KN3TxQsHOvLF7hxCbkX4rEa7bvNzN14YF+N/CgrhF/+XtTiyC96a
4Q/2347JO6pdLD7cfA0Jx4hEn85ZpdGDv9uV6Ce9Tkxni4xwwEuk1Osaz58OtQ4l
Uw7ml4j4VoAovVV6+97mxVRT+gmsXjo3IJ2+I7SWNfIb7jmYiCeDnl7bPYqgbpfX
6VcdWq3+QAKXQAYB9v9ORyW2tNOFi5763CVtMhYAwyXoKAYcddqBXi1L027OrzSs
aLRdXIV7+TqpZkvz4JNJ8tCzHNUMmmm7VK+PAITNyu0mGLFLP8sPb3A2iHppgXgN
c4ZScJFTxyi06kK4I73pKtrQy9giGGQRJfPli6lthzAL1cxxD3/zAopmNRn6Xfmc
higoW67Kfer9GHDdlR85lwPEJWUGBt7DONQgXb55c49BU5UzHT2X2OlhR8rsEcgF
dbd3oO8gZiuIHk3LI3Qlj0mA6azhNgD8kuZH1njrOynaGvXy4dn4CcK7Vg+Fp84j
Rn0RuRmdkxIEfqrm4HpkXhzH0afHYzjOkAWgUGzEIQuAR6BK/UJFccA31jENE+sG
jrkNl8sdvGr6eAHzbfvwMZ/EMXaIeZ9ORIPn2KhfmeiK4a1DR08q533c+DSDob97
2F7+33oh91Ha3+LO25RMAdgPW1Kjl+bzXMuKCqAl9sX0cJfB6vxInGBBAfh3hV7g
WljZai+waa8+9u0ExqTBg8Z0GTr1rbv7DqRNbSz2OxS/rN/HDwrzDBmzpOKs10Ko
AuZ9mJmPKHXNh6BNzg3mTrnUuUX6VLLCnRV4ymCn0saac3jhVyF/n9sz60XUL6gn
c0Jr8Eni5e7AGIICVZmefnR4DS0t2m747/wGix2TIWJX+4ftDmNEvfkx/w8Z8Dzy
fy/iFJxsJG4GIG6J1kPQZlJY/91oytg0+eQfUhSNGd0UXAGO6nvQTn9akz979KCw
pno3OnzItCIiV8cXSm3h4VrEqW9He5B/TOXLidNkWnCl/ccDxjF3WP/lYejU1hbk
zdyW4//gyT2Bg9t/0qiYr0YGpPN+nVIHsG5P8qzgA/u3FlaBId71of2zoXHN2CIW
o3q+Un0VKA4FQiyRHFBnOVdosS7Guw74BflPqKhmeHtfMRwkhN+9SW1ec3tcxMME
apNu4h4SQ3ynr9T0hIQkLqzudwHOZ/+iJck6mKpK3eqV3/18CEddyVj8YcXVaBhb
fCA19wBqeZgiSLnmnIDsKB0SSuLFd0UZiXTCAtryrcMmchmnDEh6PoSSfehocrHM
dN2F9RcjapIR7cAGvtcawKbqD0udeeLbxdzmrSFUi7rQXBErs0Jynn+73v79tXzD
j7P4Vm4p3TlAQrQ4y6EVIicz/BeDZJ9CqR+Lu9WKVi7oFKrblOmgkcr1Z3IjHmKh
PJ0xFbzEOfHigPBZvkVJZoKXi227vCbjJNjbnDzWlRGy9UTNVuT7EzqUZAbfdNU/
jh/+TNxSgcsEhxMmOQvJjLerEbt1ZZB6Hcv4wa+YR46YW+puUz+oEcfwzVWNSjvm
FzvL50nfjbveJljpE1YKy6zpg/8pIxcI/sr2NBS0CulEXOD4Jh+bdGBQhVLLC7Hq
MaDZy+RCSUPOJaIgZKOfwOIBUpu/tJLrxxvXjNCXz121JasA63Wv9hSDAqGrt+3F
It4xwqyXZGgVnUEaGhb/KNwJVCiR3Hhu/bLNCidBsVJf1A4nhKuv6wNxRzgqNKxm
MNGcbkxfnDp2Rl2Z8RdkY/kxxKDf2FONl0DAVGd+eeNtpa5aKN9L2Uq8z8SMpJf1
tfwtiCJg1pb5F5ENrGFonJeEhyNTqn6TkaX6SmWJUo0eS2QdwOu8Mcg6PLZqTm0G
1UfOTe6EnOTyUS5D8xMIZCIpgy/M07XffmQqAUzMHYotA1fwRtMi5vZNKeanUiWd
0TOVbgVHWs1srjuqgNK1kGWVnhyj11iLFV8JMdywLJG9lWkJ8zVLoiCW7bDtvOeH
GnVMK780E/uUmUc1zYejsS6IsWXbQ7HX5oyGX8ki0Ana6LJ5UcFOfPIJhPfQ56pR
FyAOJmzs5xXNRLW+WAte5nRCyMsU6262yUSGqwMDYlzIE1vWXvrbXlE+CrirWUTM
7jqJkPjE35Ut1uRnRTsvkacJiE24stPWLyCVuRODpFRgdSYGTaHgEj3WP6uuD/S0
stFsBp5qVmopM7VQgUIq87jIUDZkfF5QLMNLZmsYhE5OS5M8GaFMyo4swJi0c9bX
hkYzPL8rT2u+2KrTXODL9gpcyVug625cRElO+hylbxaBB9U1zr48iLGKTsTCmFqX
gLJygf5PKyzjU3vKsuaPKbjEa5XhgB2m/9jInqtHCUB7J91fw3rhoBjrDFxDGiAP
ysF8C/mk5qEF1C+neQ2dq6Zwv4N6fHPgXmKn2dYjhuGy02pCQmjxccQAGo8qwf3g
43h05mwn7oBZTO4Hfct/SA2u1W8/E+QSI2oSAKg/k3olFMZ90ryjWyRak7M0nerX
A2+pHCsaqAKiyFTQ3XZ71PXxBfSxuWxJkvTwpKTLZqZpJKLcZ7g+KqytvirRUBXv
OkUu13hT/7I3z9HUBDqTkfrR47susMnZPjThzlWmmZ8X0iGPK6tcVyFGRzI7V4L2
9c/PPrc5ahZbb+kAXwSdZh84xaYPja08iySZsGDaUUuA2cBV7H1qcKm7ZIwWCBOO
oZ4b536YzFHyAF0lrdTzr33XATprgYplpBjbuYCEyFA7oC4hsnKEdtyqnlrYqug3
jYLU0QExho2MiJCxCCBbIvc/XhfBIa6+qFRVpdB+rjMSPuD1guJd+ditHFfPx6xv
f4yxFtYAVD9Pg9BRUtPjtGcEMuSZh3+uuKCzo/eNBl+zrQ7htFdXz9eXTd6gmVko
wUs70hUpL6t99Mn68GLMfBwaKXpsmcUrth05djGziz5/Fkvw0YjBx1EpgqQgVhhs
eWEu4gt2Gdu6HhHfYrVNqIxiUduVT9M5SA6/KVJYAxKxi6oDEPOO4Z0K1j4WtQ2j
8rCkH9ltnEWwCOFHP3KYqxGESFoKct3Z0gqCF0bsSe8sFiPyplwe4HYts0Y+4M98
UWnWmaropHcxDAe3ZLtK/PKp3bE94GFTDT252S7DXmhnCYx5JnCEOb9GAmMnK54J
wpgOsvvm6fLVGpYKTxKjjpGxFD/sRmySV8lNwebZrOBDqyDdBd8xy+T7CAwnMWIZ
DTrzzaig0VLTsPgePAbZG0plCcfN7eUPJS++GRmday9HpHgRbFPzfSwPoqT+rFCQ
qVo4W3kKuPYORWpouGvrvxNTvAsmBAfaRTGs7cg2RFyRn9kTSeaoAEevl0RkHlLv
MSrDho9+QCk7019UJ1SAC+gG8oB2+8gmUqbqaCgWotveMonkj6G6qsfj1CP+Yc+7
evodqpdqOd49ApvPfWShAbUJeHFtLpuCJT5xFZ9UYRGjm0b89il9DOPzb3/0hPU4
9xSkMz/bt6gf1TuTGMhzSITt5iIlHGx4EVxDsWJMWwWXCVqZWB6gQbnCInZDxW53
pJXWQZSkuM060jg2feEArY+RmPR07JrIPcTVdxQMhMB8SKnW4s1zccifXhll8L4B
tHodFiyLRKQtvkUebVfXWvEz8oy8NeZLzmUHiS31QkR2io45oM6hxXH0QbSVsDGW
lhej+oWwdEypMHVWzj4J/48kHfOCt3Iw6uREmZoV7lRN3LtTiNg4LMuw5dhtktD7
+H+3SpkYIhmt4Y+yXTp8eZGhYlI48rgBVa6lK2P/1LKtehZY8ICINZ5MHh1WE//K
LuzNyzZ8/xtE3KDsfBHC6otJT1BT7dXh1oK/DM1wHQwYeUJy2VyxMT6RgZxsnrBK
RKSF2p8bZt9IpaqdC1rNcw55CPQxETNBIfN6i7OXYnSkESl3YIaM7OgS/EHDghLm
wuSOTrpW7XYfPc3uYwFGQl5uNKw9AvWmwYTQSqDe8J5MX9yFlcf9G2k2TvmHQCYw
3SBWtgnCKN4ywTIYmyAB5iCqYe2/QQJvc2Hkuc8nXmBjhBFc2rua4JXc7actmG+X
IrGvTfq7ecRJu81LXUszmZWqHEBUyfk83cT7rdLQzATmL0NVFEX0zNQMsxic0JfC
tqnDTUPzDNHojV2kKOhPMc4aEVWkfBW8h91q2IXd70mghrW8P5uRjImFUg2Ace29
UwnTsmwtUjTuv18CCCNFDhjwXfmOFnmT/KudwXw+fRmCFonCeT0+qIG/2/YiRSt7
3cMjEcfv64IEV36ws9vCwegb3m4mz/gxlMHp6OOgeJ146GpApFhRM/RyNoJ/S4PD
WtuJqIsJE3Wu1/F9fivJSKWKYFZ2L5PRg8747avdvxG2jO+KuWDrXzoE6lKmNkVc
SH856SUlHZwJ9khvhd84p0iiO/JEAq198kR78SpQcRSKDFIjCKL+Gptb+wDtvXHv
kgZqCa9TYO53bthNilFsOjPuYDOLhMgw0pmBx0Fgtx249vXAhHRUSAB0vq2EV+dj
cEokMhx5jog8m5NL31rNmwXP/rgPD0quxMjOtYziR6FCRroE82BGNgL2Qlj+3/AY
FLjH7xPhcHRQhVefxbny1Y3h0P6h5ZM+L1RNroO17+fPlP8ocwKmSqlZhcWcglja
jhdvFS1Vnq3QqfZ3aSs5H78Sz9s9YPibJYK0jvec2GzXPp0aLSSJ4BGbzTriRnGQ
1a7Jvc2+7byy51ZGtrKRUmQnmquFKoPvU1vwiEeEESsOtAax0n9Lblu23inVCjpc
TcITfHNRMdsOpmpIl0OnaxZlZQpS5kLhKEWTQnM1L7MB3HAOXwtF6QV6eS6sZFi5
p5bBTfvR+1bL0tw4vQLzlTx8RFKTP+m+46mIkipFTfeLRG8EKNFPZVohm8Cg8qo6
FPoBgVzABwJmPvUEMZD2Wb2b1Pp2/vCCnC3qKri6qzXFuAXm/p0geSGGnlSUgGAC
W+LzNBUIYl9w+gZFjewa+yhvkrRF7DBxCXZu5Y16o5rVfAkZx/g87itZrlPzjCxs
YFm2jYCIzr6HqEy9ko8SRXXEIT+rX0auUYV9z4rECvBxwcLTz4Sa9q7O72ByyNZp
Lnn5dQPjzw+CfvpQ9584y5NA3TCOWJwNM0EyYl2yow/TDqYInJckQlov1HGsMcll
xeM31dgctSn3U2Wl7mFM/C++eJKtAjxnDMe4VSm3/SKKEBg5Jxn5h/xjcRt8qnEu
RPUT2R3183SUtO8I9rv40ezV3JALnXI837NQq6UDX1qcRJSeBHy+rklUhGSun0Rq
x6fr5mrXgogGhOv8ssMreGVCm9tUOpU2ju4cKTzw3shqPahaL8/wQNOLTiB42ww+
/Kub+JCofCqgDGuahv75BCjhju6Zf0d/WyqmEtXbQVlZlsLQQgLqBkFs9r817aDC
IEvkEJN6nFUYD7oWMhN16pCRiOu9YIDUGRZaLkbE5v+g0+/jUbTLXYAkfdbby4CK
ij+aAJF/xmujXjFzg/nTpU4cz9nzRLj10wFv5X1qRDgqbcKk1GsgXXail2luN7Wt
Xxl7/Xz4IcOsjwtol302k/4RZu2cnxYz8aePxyCAYDdmUs5c4aNszw518RliKnWn
vjcGiqwhYWGgamoMxJJnBteMyKzgyiw4RQLv0PvjvoyB0jlgTyYKvQ5aw7lpU5v4
b+VHiMUoxskQ/RBq9Ug2mN6JvJKGOJDut8RfZtOzd3P2vrs4W//uzra/+rQebFpX
GIG+GWzaG2orsIHDiR6S/DyPPI4KXzOFl6mXO1v3G9WIIjN7ggPz6vcfdFmyPRqP
UhJTAmpGpDIGHzAS8t0UeUJlNBqzEqlJnBl5YemdmVJL2MoVWROeAn21x50IM9mp
rjmgUcFGES0ojIT0q0ssH5Y6sYdSs5jtiYugJ4CngdM5t7Y4VhLPdPl7LM8HGMRU
kBj1+AhVafbwR9BNWI+DMl83UmyNenUIHZ057JMSJnYH1XuDAWXoHZwcN82oTcVo
wfye/T5DUbrybVFfv4S9ihYtXRYuj7UWjb2Myg8HCRGbtEdwYSz+8oPewZr29X/F
V8RnoA3nZr7uU4zh4zYDsR0uiqRBSLrQmFnjtllxw6i8R4Vg/qovkoNRFzRFNmvJ
EC5RgZJFJYI9tBLRCCLpAJbrYxXU6SDJOQic0XZ4EaldpYDXP6O16SCRjgFkuwat
SekjZZPOC5r7zDwpXx+KcbSM7TW01/ORXIVTJrMYlUGb6mtozyD6sRAfNmgSY65d
NXQo40QcnPA4Vp8qJgrzgQG0srqPDhOR3/1BvVjz2gp5e40vOen26Fzebr0V03Wy
LxmLLqafYXFPB9qcRWUD+TTqlBXYFPxMjTv43omALWu76mOA5hxYNd36FSNPUHd5
KzXBE2h69rdeeu5/Syf9r2501sZlGG18cEhSw+3uJEkeal5xPaA6YE44QC03/q2t
p+j494A9je09Q4t7LZkaJE0+aiC+eTqtsbk/jOW4o7g/5NtAd55O8V9NSNfr/4hd
qtYPEDxhwrei7/4nbPA+bjumYaMR++Sc621KxKM3Vh0C2RJ+lm0fjJPwa9npAGkx
Bfsl6C4ARZgKZQdB+2AoITDu+Arfbja6IxYnBeaGhiV/1T5S1Xn8U0hSerQZvHTC
z6Gpfhr3KCYdR3OmAcQWvAtTpZwQw2n1BOEqXYVappnZgwJzUHzEXTOfXfJQld4i
n/e5GLiNxGYc2t5OocmpiqGEgNwEwdw7nqdz9Ft1uJ8w1+jjyRsdVmVwUj1sJn6x
2rGrAGpw1bzDODQdZNOFggTUgsx7E8sgEgQFrXmZNJ0tHoyzh6KtGbP35nTrQuWo
UhVlE6O6XRMfAND60nh2h5VKKj6BDpSWiEmzOc17zjIJHHlnJoOkSBKvr1wUlviT
yoMbUiPdSNUnAmwoKyr5qUdCtpJ8P89GlZ5ib1mvkJm2BScfKydIXiZvC2IKO0yl
Cs3P/tISH2f6ZX4tqYqLbyexBziedFzljEtqmRCqbP8wO8h87R2nEgp09CE1+hZn
zsfKtug/VTzdemUs9uc+sglcEj+qYnN5TCI1YnBrOZx5SHeFuRN+2az/hG1ZpsdK
rxA42oHfg1PiUt21/nfAiCPNaH8Ct8jjKRYXnBwVfeXft2OVzduRSqdJj+ssEqFM
2TwuDKzzISn8PxzKIdiWUm6C47YDNTe+i0n9B6fwSJBhstTXfm2YrmnBn6mlRQaf
aYhJO5IKwuEpS44SSnQR3eoaFdbFHlO38YL8vK7OGdtEAq6Ra66ZxRMxIMVy/SrL
6jhaJmWRXGQcalGUtgmb5XwiMqnGQ4exIhHdOEdiOLvwyvg7fo3opqmDmJa4LMUS
t9rY3X6IbuHA0laCnin5S/lmNbvaG51s+8LQSmRsXu0Alskd5Od0kq6F+RUvSTVq
gBPJumjfK1Kny98OsHK303rxxdy2BZq3aXP28FuqPWbj4cNHvWXFJPggHRlHFzCA
UIa7Y3QSEQ/hRMVoLEKRIsQyvrPeIwthF8xV7v2FVxboHo2aiM4FZ4zLQgSUjfXX
2YPJj/PcuD8yXY1umjJgeedOdSa7LvEt2yS6Zd+oggqfO4Il+u0eC/+Blz08Rvmh
UJ7Tr02kE8CSsbHW9EFwpS2ifw0H8Z4ygxJ+cnjPcbDzp50wGviBn/m2bhG5Pt/x
8ZsayfNObVbGb4WiJzVQ0V6qHyRAZURCi0l/89ijJD2gzOeyD1ILZ2gv7ULsOmz+
0Bn5nc25VAFy3wNrR/CALKmDGKYMkma4Rw1rRXlz5tHReFKuOWVi9keN7TbUPIuy
KF/pigrHH8ZYBj6qw2AiFFR8RKJrSfFMxW//eTXwryz0xDK3KaxcneLcuybI4aGE
HfpoCZ84hyCY9lM6sW9HwBjxdmM5vjsnaA+BvQR0d3JQNJs1yPyl3RlCRes8jAes
bcJKn2O742HlqEOqqnmOedtw31dnOLCuwO74nbINJ2ihIC+eq5NjQauHQ8H6MSfx
s1AZZwUWCUt/3YglstGKjdZ+WtC4wDYxuwr+lYY04NO2KsopNWrYvLDhwWl5po8+
iqVkA5U17tWscnRmd3kgdNyIPmmkDyXF2HJOxXEQ+PblI8XD4eNzDFkU4V+ynrhJ
Gqs+htHk8VfTbpNI2Yzq8zymmlKwGi5X2D5haTfgcq6/k6/hm/JiHJqiVna9A/kw
tqYEFR4xAR7KQdVfIac27iiZMW5P5m/KXC+yGDGYsSUdwWVYr6k8sd1J/saI77Zl
V/6o2935lDeIkjyACD3ZaAV9vaRSOdhZjZLlmMPRSi5w15p/UWuClxQqwT6AyXX1
64LC8Kt0MbzkQ9NotzJSifzNDQ3wmZdiy7LV5zZxjR5G7juj8E0VIWgrMN/yn/Ll
BsenkQnD27lHHSZl7Hvg1/qH18TbEQpgyXN1iVl9CNbMl/e06/koihnhs2/ylm+G
QVFHONC3WE5aBo6JbDv8SFAXgtqE0G++HHyOaK8lANmhMUGNHRKwt3bhZOhm5ti0
cgpJVWk1qyLJY5HouX4RnInPZPRL2sgr+/QAEITt3lea69SPCE0dQXKfGed+715c
TIh3njoNKK+wzOSazn1aP0Vy1BbjLIZzHsq/VjfgcrZVl2VLyNd9VIuvwkVVy6wj
vMth3aQ0D3IdLEjHLbB1O3rX81qnJLq1UbHx2YPAa1bLITA0i7y+U4oCTFTEkmgB
mKwllSaUSEGIeaCOjOTPeVn4Z7Yvniq2sWxkioxOU3lhdTgdYvhtFro3NDpk+pd6
F94IMx/MSc4IuCeLyE8NIdQc3mIEJ3BwfILaX10GPWVBCWhs7oUD+Lz/XhgXgFVf
qvkNoNGxRFxDamFJX2loFxEcxERPlBiW+Yw9xv15QvQlut2vwU8PGH5vC8KoaEx0
rfevbWZsPjDQAnw51SNBCvS7rrnAXm7OwXjJYdzfIFYMUkl/KVC2p0bgkf9nuujc
/Or4Hc7zzSgdQoUaWFRrARRzKi3+EcNPEGBqVeKauWuPTTCaBgjJYhIFphg9lk8p
cEHuaDV21xAvE90B8cJIAcYRUzvH4frgO4PEEXRKDvW5bn1HL17yFY7Idt/7o05L
toDA3wSfw0MOWnm86foTDF34sW8IXoCaGWt3h3vTJXV9GTird/iO5DukFrj0z/sr
hYPj98fSjnGZDC5o3WnyPX0U+LQ5jth9nnuVWNZAIBvetrxIQeC+kYe7nHNOLFqy
bNvm3/nFn9heBwaFg14gnENmNOvxNL7Q7XZFRI/VAVWCrHW2WXDIFiAoXOe94fBn
l3tG6LdSag2+mGElAQ8S9JL1EZmmdpFEGHEUqEbD/5y5hcZGg+xXlUI8BZUwBUfe
b0UoMgfDCnL/kaMeOglYNd7Nn6MH0Hj54mFskIAHkEf0pEg8xNX7DbAko36pB7RD
NRgKz4dN1YQUh9NrcLAMs9znT6MFKdQlXEuJWQ3PkI8hMhcCG8cAKk49C25uRfQR
nCQBU7A0pA6Fyh/jTmwmXMD6amZq/D66yQ/hp3yvYFP+idZPG+LKtNoJIQ5ix1/Y
E2/PsHFgev6/Dh+gy81PFss24PbtksmubYubdtYjsz2/4isJ1sdKzmiIbhwtkS14
wXe467cK0zU4d7JXg7xkBxiu2fenMgnH3vw8dt8mSpVX7gM5AYPBsY0jvk5YNNKP
lXpIBvMCl/PAjfdWuJ23CHqfA3Z1rDo8jlUyvxTo47Z676sgwKVp68Kx/3ceIhmN
Q35RWDlnjMDyezqkqMUWE4sZ/MCygeMxdWvzNCudYmlMY5Vx3kAGLPqGRaMVy5Q4
c15WyHiQuf4j/6Fl0Nsi6UmyOt+r7TVI0QwzdTzTTtbee58ljca1TrW+deSMyYUS
yHO0veiOKBaWpHvQVnRtm7B/AX6md/GiVtax+baJe7hQoeuX+CC0iwwGhYkV/r5t
Q5lULtgiEHRBTIer3eCAw8wDa3X5ZmeVOOQyzPsqSJOL9A4C52Qc+N8kVhTHrE29
4IOAdGmc0xkE5Nincpn6DYfqv1e1PRTeDCbHzUIzSWMGTf1qHLAJxWGgcDpn8mIZ
8Y2b2XVVihAMqUG2Rm11vgFd1nrjA9Ommu4PhUcXSdKTgfSf99IKBaXlkVptO6xg
q+acfg9uUwJVmq9wMHKe7PkvLb2Mw78A8/1y4+pTHXNVrgsp4ziOlQHKRaBBYDmR
ISU3dQ3Cyt4CPjyj4phENjmsO+xZsY3P2YaYWKvSlbK3Vr+ZZuOHeZVFB5k3bERu
o5FTMwvnaJNRxNx2000cDkZZ0E9TTIQFoT3AG7uBvzijfY09kv/sfGQCbeFetwe4
yHYdEsav/3RZLzBwgqWueJah9N3PZ3OpdxtkgM35XlfgnI6hCpzD15GUWRrQ+Zz4
uBS06OrRipMfNteGefZ2uSAicVi83CHjOiTVYjTfcogwD507SO2e7bfBmXdwF7nY
vVjE8R+AwPf54YtZYeV7BOl4DBmvabB7fQSL7edEddtFD499XdUbHLYxrjynh4tf
JR+7TXMGBP8SZknjJZBr4yHj84qRBGgBEVaSSkeRrg7Pd9yJCBHa4/HNZDVUlpat
U0Ojxgq9RkXEdk0rYunG3xdA2AdOuSQGTaNbEj6/fRVJkfNsOZh0bl4HWfLnkbh8
GAfiIEzL7QTzsgyQ+Ejf3ByPu5IORyTUjTOthEmYf/GHlNn9GsC3X7u2dPNCf2Me
L6UUHwUbY/YCJnsLNp6hOF1RC5ELQDL0HinUTWOaPMqtgv7PnvClhmnZX8u3re8q
9XYdr8sD4n3V8C2uTzEj0shuOlPBEasfg6QXuYKv+VR0r+Ge2w30S38Cp5uNScno
VDbGnjv/qcDGXkVyq+uMX4A2EKQrFZiUyHJB+znhjOmw3aMInbkgOr0QAgUIC7r+
QN3lifQ+cBe57HpEo50InGe15uRKXbi8MN/dwdCEVGlRKs/TGMX3f5/5s8RMEQCI
j7ACRzLDBydAW3v45cloPErs+bw3ES33qhXg10nNugHEL/fpr7Ro5a+W6frkc58r
FelHJTV6eAxTKzEsNagX3Ky6L5NTCa87TufGuU+LzlKk/Qwh2t0IkkKarb6byX8w
JVRBFMeGdN0zBp3crvH/hCQZV5H1X43B8K+hzeq65R3zwTOUZ2O4d9J5V3ZkIC5K
RTxwKRgVWs1FQhIJsPTh3XV3V6OtdrKcafKpowDjsydzTIT/ILE6QJor+CS3aiXq
03ge/nPEtmXaUZ6ZUFb5ciZ98iU0CkxubYbJW9RSvcXmne6Zyu2evhPCfHi8iWb6
fCh/RtUAHZrEAzLkzs4SPuTojRIJzcbwedOjL5Z6Nzn71ogjoSI/1Htz1ouqObcK
KfkqXXsO7Jfm7DFgrUpeeohF+JDEsCtZEcoIZQhubDQiZA3raaRpjGsjxM9vlF49
dxND2wSHPSFAHpWRq1zTRakxij0fKWx1QpE+weU+zfeFu5u7dYNs1tvwEUH+VMHk
DVR+bAWc4dAVh+5J359/fvxmsk/M2c1Jcznli1jow2kewXpEmOzYOafZ80jcxhNv
r6uFdrRjpOu84Oi5BPj+CLfedtDIFydmCSsAoyCkuUjXdHhq0mLKuDdkfslMHAvV
9P1UTE0Q35Ard9yCntHWcMGoaLuaLI2U4S8GvHHLCvUpe8+VsnIo2efAwADEpeTO
3zCmUa5TBG1Ju0OMvj6hNbgm2uemcgYyQJ8IJTO8CztDF5KkOpRavItrVbA/AsX0
BoJg7MNXgz2EZ4SHnMdvcQWwvYk71DpQPIFJZm8H84CnGllSOPPRBgm2CBKQxycy
dkl9HB9N1uOswa2rnSFIVeywAQXiYhGRUAyfHqFC71RGZFhrYrSSue+wV98nPQJh
wTv6BWs7S1rE0Ni8rxLUDIV+A1D2OtF3hgJnhCZLXe0/MM/r60fpXnfajBCjIpQn
jKp+T2a1PnPS5riaw2K0VLIJwKbwx10SkpEqJeePCtJa31x8bcqnkosVqYkX/B+D
vJA8MadR789io2Ar23wHo5/2IC+1y27vQ8IGTYtCot8uMA18i54tLQxs6Umk5ITM
KuA0x+82iGoiifWxVqfDavcSuRySmZ/GHoe/Jv1ZHGuDTdDj8Pv/wNpBF+LN0rZh
tgScxBDuk2UyByVjtLqdTTHO08len9DxqiyqSe3DIVljqjMtw3BctmVM6mpzdJOU
MTDgiNWkYiC/sQoF/EWxUB2/qk5vi21EEdVmZzljGnWqfPL39AoWbKoJI+/AKndo
q70pe6pDVxfCLcUhlea3X+hZzZq+w/HnnN7TleGWhVUEfmgPyzjZouhlD1MN9E9G
37PxX+79enGxYQdwkTMqCU7qCC3fZT1glaZvmSmtgStOWua3sKqmj8uMt8GrDoyd
QKEaOeZfh8DbuCOWG6aRovVq43ZMisX4wGXATdRK2/bPuLJer6Mv9QFs6+ypEt4c
1HsXKAJ+7/s5k75/+s8tEYGuPnv5hmCKwrzJrVADkPgK3htPGpjmbYin0aDXQz3o
7gKBtyQLD6ijsbScwGsz7yG+mHU4aaQZhTtwQpOg1Ft2XaheQieZPn/Z2nRSkUnL
AL7QW/bQm4vDxTEHkeoD4hXjjp/VrMO4QtMxCA9s5t+ulVUj8TNiOuwZPd1/SyAA
fY0d1BbAtqypmysSy10ev+5l0wMJjrMy3SJxAClxFtwwvWWglmFvjt2+FJ+RkIUA
m6yeT2E74yrn/WdbQqg/QggvL8Z9TrZyKl07pnKMsh0IqarP1aHo7WoyLJ4puUsv
UvBPGdKOrl12gEGIZ9ykUVBA5I7DhLkUvWXGGZwGBgA1EtO5gnIi62/SFpWPlrqx
ZX1QNUOyyGgVhGHJF7+LUFDE9Xzmbn8CQ7ZtD2s+p/yt1sDbZ5aAOIG1Zd5g5Piy
TrUbI9Xs8fI2z/72UonAZCsmro9ffXIaw0tqQuwOL13NM6SqvOBSvlBUUuCuNF6x
+Ghz2PAeDxKIC4KbmMEH4UzUtwQfXHUA8PoOADdkJvAvOLWssgGDFuqxYEh2XVK7
UQCTgC9TARY9vE85KiPKiMsGn3y5NBw6lbsWQTn6t6aU2/krvN/pr8Tr/AzFn6PT
i4bNc21Th3ZE5+GAhVsEWMISztCHf0ePc+uyNOziiG/ThtYXpBx/kRJDqV8Jcqj8
WjRZExEQGf+P0wXnLv+uV1t/d10cpH1v4NBwH8ZWpH20eoZs2U2YHSMa18JwK5Jr
pmXTC/hlylv0KlbcKinKLnA3gfL6DMhHHaqt4AEFJM1Yhb14ObOR61YsY/zEcLZU
6gG/JpJBZ7fKmJmiL1jbzIjijoiPlhxpdReCHSmo1k7A3g+zhzlqMXeakLzuEWkT
YfUulebOTQgmRmdFfhb1cFKHk0EdBN6LqpyKrViUqVxyzCK5JvVLI77PQJYSlKMU
zWLWD3E1GpoE2kVeaE1g/YvwUXhVemVxZT898oI6nqmx6bOxMhqRdhK06I6f1a60
r/twM58ZJVMWOqgA47Snj70Rc6JDBjUEI4n9OTMjpEfOcXMyiWQ0ZHCWo14TUUGc
l7MHlNa5bv5b8FcN77ebh1SSKrh+j9oyv0mcpIAeZIjRxt775rDnzWse2C6TK3Z0
h+9smNqNJirvvJQ1nnXHTAd1XFvWs2bjzAq7UPKM/xetHbwQWOzkN74BTX8Atjof
AngS+R4yFtNh10d3FVfk6dagXDN3gbiKnA9wJ9h/VB+oYg6E+ykxj/yJsxSoa2Ob
xqqm/cjQLUIe0y0Ubx8y97RfKcFYn+cdnQ94EtWRiEFPOBmKsQ33JUdGXPKx5w7M
6KOkjX4C9v03DKpSIN9iPlLyRh1wbxWHTpkbz3c/FXgbmhkYw2ve236Rz+Pdsn+A
qJd7XbSNKAeoRT5waThXpehrIca8GyaktDoyl7HduFSNs9kSrj3qqPPiJFURA6yY
5yQzrVmD46Gy7tQL0RUPDEmRGYdc1+olAOnXbH0eRYEXG6ny4gc/wvpXZWXUbfxg
bh19reAEuoat/F4KURH1DaG4bjCFIQzvmG2RcnQsBfui57icm9jjJkbURe+SgEJo
GGXrFm2z2flmmGijq0+PAM/ekNeqVVCXLrzCfvizGm728UvPtryTonKOi3ooHb3m
i/dZawJBqmPEZua7wRuGKd431dcvAJO+p/mFOLU8B0/s9R0Y4IwOr7Y3EqgjGzM7
2s39xSqw6FfvQ5w99EoeMFedQiYrbGvpP8GIcbUvL8hIiH6t4+48puua4ERSb7lB
D984KXLR0z0q9jd5+zpp5vFMsH8j9sJEwuKKwtENQpO2U3NcE4irkrCvk+CQYqos
U3H77jd4oE6sKZVOmMWCNgn+GRt+IT/oyu+P5VcBDPwmA4uIEz4QMY8IyWw9BZbv
C94VYh/+mNHvxNgivpN1rjObHj3K3DcRAJGkSrXpmXMKoZDGo10MM47AfbXF7m4m
pWsczE5viIpadtuBIN4sfseSYeEg4m6VOA9rvrX4/HBDsytFzVD8gPvpknS2Jb89
Uw79MwniCh6GGOq5au/JF5Ns5XfoPuTx1uE+PF8XYGV9zBRejaLKGGkIPdpeHO9r
AaZnhdLzXRq3pjX7HvXlJSAPk6kgRwd85Dy0tdW94uC3KEAvDE4qwtN9PEuwz2lw
moQjihjpDw/j71bKhwqYd2Cz5UKIhVERZ2LsaVJTMTlJ4LFoSKpamDXojgOlY327
MhCHEtIosqEi6ZYJPrS4XdIvI7cNBfDEGOxhZ9UleqXtzpB4A+JHwUQs1KD4PzXH
MZzQXeYOQYLqY2yz8pBGl9Fn2bbLt5Diw82g2mQUORL8PE5xl8xj908hoFFtb9rm
82G+vak6R4BD/4gs6TKrGHne6AQ9cpULj2fj6sKSeUwNqeW9gkc/IKbOtmaMlshV
sgS/qD4kc8e3PSuwYCyf2RLgh2t1ElXSlu/J5EpeNHkwtI3XVdcZNCg5Hy24sDKC
ANqKhru2hc5j5OZyL2H45x89GutP/4mw7EDT9TtTI37h793qafm02OYCknc+x3UK
tOJWH/1LczyPoBDvr8pq7grL47wmA2U/O26sdDt/lcXfn40g+mUYlaf1Am/A8wJx
gXYV9fRH6MBLSv0wojfil2oh8ac2fVDDmjZadAZgBDY81lvlqWrSmwYY713HRa9+
oEKVkPeZLl/JwMP6RXKROyGX+mR+ajURlKyekjgpNFTKShS/WOeoOFUuSvwSOcjN
OEvUWh/bc4C3BFKxz8lH+hrCMQKUF3UbCghLskPftMSDXqKXxahugdvecxMH0LeS
9kZZjG4qiEuL9EGks1JK3kQhqWeBgMo3k+B3Z1XiIoqYqHAxIrYPd+C7F9l1v/z8
Be2Xp9KzcewzOll5mlB4MQls+etUKVSqbJFW0dKWNpP1LRmBplFq2lq8UDxtqMnm
Y78BRqDAe+UU2coAyoidxHWpAeqQnauyknzcjxY0kmfhe4OKSCCFf/x+GDLJxDN5
viKNhyWauGnTGcif0ZMV82b0H/2nPrA396i0R9i125UiWkTP5ogWA4ww79XNqfSS
Jl0Tx6BZ7CAwg7pGv0mBY/aEfaM2JjfKqUX+r+2so2EN70PcQaV1EkxB718za3sJ
t9lERQIO8NIyTvFTcMx+/DqsZEpzYPjQ2dL4xPENz7dTnvyVJZlVNTisizw29ZZN
6soUPWthiqFiUsbeCxVdWPXwMQmKKhWbih0XV30JIxOLNvf8TgbavXQcU/XW4HIH
aXk8fysLtkbk9vsHn9Rk9hJqJ2hQ/ChGZzZ0G/Teis9VjvqRNfS0bx3PZF1+RQmP
sPwqDcFyOJSSBtuzdJMxwopLJrsBfIyC0YDsFpXJYAVGn3zLKYnBPsuVADc9n2LX
k14FEGlYx8rXdknrsF66wxjIDzuE18t/lkDhEFk7V3rGbXBoSZkHEp5dCJcWzXh+
URiE/EejypIJZyOomokaAXE463UVnQJlQzyEiqwgTbADNMU6QuCR9w1SWfvvNCZX
YnWfTGus8OZFdcomW1R2pXG11SdEeWMOE9pNk4DnW9oCQTM7bGEPeS7C0ReBkuG4
rI98qvU2uUE+atAZ4hGPQTEP95Jam+MBlR7YpYojZ+qXXCT0Q/3HNbzkjTwr/0RA
Ljzf3ZwsLBTeQvQd/UmEWUkGJg2f6l+SmpogUxRPhl4X1n6h/GQbuBlmVFX3Z43d
ZLHMXaKBWlNgrxrcSZYYnTK0mavSbPtDfdxAlyYIEbFhL3CHwZHnNkTkfQsnN/G0
KE4jmXG/DA4qz4Uh1sj+nwnrb2Gh5fhx2uX91PW06hwotKtiOU1HbZFu94tsFa4e
K7DJCPwpwEstn28QZ6HcIeTx6rDUmdMwn2r+wc1W1VvXjAC6e/Y3DeLpR5QNL4D/
StO0ezdnO7/d/nRcD4/F05JK422mBOkQXKxWqsltGj0WPd+REyauXxksxAHjZLyh
XlcYWF96Y6nj70Bw+jSpNBE7bUsZBkWZbBceaQcfkGXDEbWoR+HrTvG1P+LBWhwB
5iSOgRaqqu0j+Hrmf/rXJ8Acr4QsAAavWbDZGRuko4rrbCdcyCOwfzqbUvRZcTHA
9K8eV1O/5M8WPYUpt3G6dcpkyOTHnAKRk2OAd+EpfwxMaSJDJww+KbC3rResIVh0
L/0qS06tqIWMZZ01ShO9YLruCXevMB/WGUXEkN4xiOvMQeuRurYc5WvJqJvBqDt3
aEiuOahKoHaZ6ZTKhfYuBWfCZQxfPuQybO0qQr+KwhtW/UYeraP40ax+QsuXPHAS
w0mgkatJA1qaXPRHzjoAS8WiswMvhFmUKt7/Ifmk81i+vmR1ZWN3pDnIe1JUOI81
tKdzZm4nuzQDPezMfMq9hBFsJKSQnKOKjQ8WMefwoTlxVkkzTxYJAXT2SKgQzkK2
4okf+GQf+hmrSYj/km/TMUAbANR2CYt0ixOKj8UXZDCS0UgBmwkyOujujHmRDaXR
nYHAOLzW01e1eUdV5wzUA8kih35liOtca/Vf1F25LCI/qM3G+4rYHna5IrXcGss1
NlE2YE9xy/zrFhzSbkmPEUC3IdAffkVA/Xp8lbevy2B1Tk3+D4kH5mo7P2ST9cgk
vhpwHeE4CjdBKbzarbdonkmvRIMCQuGZkG5F5Ekabr0GlmTwtIVT4GUXKt8cZ1WR
70j29eSVcqBVfIz95J225YWDZQPTXn1Rp9k5itgpm8/7s8i/SDKxS9yzh5PyaE7Z
W0RGjXCWRW4nXc9a/92VNJALiLSHFaAMsO5CE4TdpAJI/v8cXAmxQLVNsGg5fM/h
Q2VlykTImfwO2jWu9c6JSWXRswsY3M9De0vketxFCyBXwBCbqm50tqqGtN59D7A4
tHztaG5aABaxcHIMZuZGH7rTdds5gjORJHzPQOlTiIFI0jk3VPAvET3wmSreVBra
z1tLKbvVlEvIrTEtxquPZLLWIqG8PAbP9bh/TqcwDSfhCqPPr+R2/qEMwk08RrDQ
VEwNGUV0ok8mL9s5bj8sJPFZlcR8PAAVryHUg9yjyQh7wj4c3ZO2k8nYaH5ntgke
VtEqp447eS12jV14xRw/I59AIN4XwRvtM3NwRw0ce17G+PCV5WYi1/XG2TdBPfi0
lJ+8ZUJgAdjbwIEnFnGYSY3tMV71Y65K9+ScuP1ZPkcds7xhStDICxpQ+vyB8lP9
fQmmhULaeK3xTdKUAZz2tCLkWTe1ouCTj2P7/oyWBDU+uRvAbJ3Rt2JEJqyycqw7
NVljH+CYQQP51EqkZPXbWd09p4bY3Npa61v/5OvOZvAGHzLRWQsKDOP3PWZWjcNm
i+HSnvw0uBqL5MqVRWncxrdNWF+pY+CqP0JwQnt+y1Cfsy4Pvsma32hrAlf2zC+q
iimHnU2ozKiPzyyQUIBhgrJu3tdaR+ALhNd1kj9PVTXT+RWTdPCF7r0zCEkhEgKn
fWjGGNcbf3A/5u+Avxl11y+BUVjwKmnVaT75Ne8jlnlO1QexfFf90oe47I7ZzwMC
ymIbkr7mOcfUFde2erEBgenfllOJTGvv3ynlu88O6X8DlcpU2PPNEyYdekaQltt5
S0N1ajMMBVAYwmfDW646DucWSSolYi+SgP3G2Nh4MzJHkLkEs66fKqHLV7D3eNvL
yatL1N+jOToQ8HQxu1xGGn6SWU8tYq8n3kLIOxD45H2nHDQqvnbimPW8OUZi2xcc
1WSi4XwZ3Eby1FLAiXPuwY9yvkhe9WlnGEo6CdDFfddY2TTtmaNGchF5Y3CBDhjG
h30o5CEUsl1wPLLyHZ60edYwNYr1Te3c8SClHXV23nF89ONOYsQN+oqQ599TdGv5
A89sblDDgHnKYs5mAd01m1Fpp3EDN5lZXaPdPaJsHawxrp7spHdxke2guara3NfK
L4iu8Oi9NYVXGjGU0VDE61U/UoyHI/SAAdeoFarXyyPcSkgLsZzrHjYUvZj8akwb
wNS8kldFUiAH9ZM2LVIN48NnjhyB2sGMbubqfG2DQYYA1yfGl2vsMkfzbAeCjzVL
2RunQRvsCRnqEsz0LC7Xi9Dd98M75S+mttfSBge/nKfuG5pM6EQ4QANVxWriHaGE
r+yUznpufuGLL7g17YL193aitZzPwqG4E523K994NOsbj4en6W2MmyONBIsCl9iT
hS7mZxn2c8mCBd3Osz3FdMENNm71P8o7tRSuqqdBOFKO19KNiWU/bAlxXSFbtGNG
HX9gRIpK0BeGTzhM4h3O+K7jDDVhYyPxKte+tyDUXXH1Gs1Me7wvb0pFNAedzB20
3zKmA5xa1hYOefy1BJE+c+8khbGVLF0b8de6SBaAHJilCJbH4B/8EZaMTquoEMys
klsv9p03ccIXEHmYCm+AXDcMIjRe+m35hDwCEOkPhM0P6n75i2WL/vXxnM5NMbHI
1PIUft/AHpEriIHfhJGY/e7PtMgcJRquVpM3v5t7kBm0LoEsBaaWetR4Gkb7kawI
5jnc1fJMK912szbgU7QoDo/PXRrCFDTxmpox7tMfTwf825y3R/Lbgsd9ijul1yRb
tXe6qUIMm4VgmVwYJHbIARmbyB24ek5E67UpfaP9enf9wwUXPjvfzgr2f3YhNnhA
AVAxOn4MSxC//E/H4uVKfAcVLSJ/nYXNZyzWkYLU2sd0tX3c7+o3HZIqZxf526xm
V9iurYq6KCduXxJknOcuok/3QH41Nz0pctuvK4L1hPA6QXkRzixiEWVLn5zrNRLW
E7zLNGEMfBsGmmkHO+9tg7Wlp1Y+QxNcn2m2vqCrjIvC5V7eC/kf84FN+qxkkYfb
KbtZMAadDdLa8QyAA7Y2eVUs+lNzv4NxfiTOqkd59wsr/JYF/DGL4HtNTBqSUvDM
OL2iV1Y3bjxtXaC1ywYTJwofhoWqpmBf/qjVey090/M+Yn5s6EVr9n/WsOd2wQ2A
AZul8t3U/Z0UeFdWzFrwogKljfKGayvopzuBluNLeHY1AJGIGe+ZnhbO5WNdj2df
GRv8OzELP7uCtjCejpLbX6JT7pdvQuiOAC5OCiZAtpswGRH/X3WoCG2sbyynfFYx
BKR4uePXH1k6NItIv57CzFaat7U8BbpkCze2Xavilgf9/3kt5PCLiIa4hVV1qYMP
9JF5pvn6DJGG85FKUqcZ6YhK9Kk4mM4AACF1MMoERJobQCl8u5NnltiD+PIo7mZG
f9F8uWrJgbBGcpT5NWxf5dThq21yB3jMRr5ESK9iz7NKtZO9yEE/ZUwv7ToVEIAz
IuUG94Z6nxiDkFRrFn2cJq0Rq8oBTTo2k5/jrraAIbXBjULgxP+8aeq7Ve0lev5G
dDXkZyX3law72Wz2eDA53QxZEzRIOLHE2xoPp2QqkbeClkoAUm6ZuITSou+IvfJ9
vL+3FuAyXlD+skBimo1MefKEEOuLi042g1An59cJEyBBCiF+PSIv9pJDjqwoXIfd
JtublGzM90Wk4EnTD2BlRJuZ8w7ehr0Yemnfy38R43u3W16KbhvJCkl5wze/OMzW
JW1JB+rCpuDanAQ9I7uEwg3+K49JKcdzrzCvvCYiITY45cg5hR47AuKtR/RJxo4Z
UyPkJ8zFfKM7uxdwTpL8aHfT99oDRRNe6MfQUbGJg2BsJ+8xg2WNRO5vrmCvRXZO
DxZ+Zd21gJQVkADZaQa9P1nk3D86u7/fJQAMq4qLCxPEKKry14yWIR2nRdTQLd4R
AcbTxVuMg2Y7ekK5Iidxw2Pjh/irk3zVcH1+s8L7e65YnMXWy2z8YuWQMwd6RU3p
4eiwgL7m8nUABb7PlGGdSm2h2fJWvn84FGXBrUPmbiyFTXtPp6QtCRUfb9uKoOFx
kio2qtfuN4lwzGCkFp0Vpn7yyi0v2KI4ETSa7pS7B6SiZ2hY+exIRLCXaSS4YtfC
GJOtVfsY7oXZ09po8WyOo6AUqCscU/K0Lioy15ejrsUi3HRoZTfx0QwV26ergIIS
VpgzErrW7WlqSkYyk17rAwOvFpuoIv1GALz0YpZDSs+j7WgtSUCX5o3+TSNJDa+2
Kr4IHxDhl5dHG5UI/T6GXHq5fffPBhnEsQWcFJHSz+UhtBnw306SCasg4HVqdnO8
aNgw5TMIX8n5ZdBhZQbAYHNmpHl7N00hoyY2VCRKfjlK/3IJ0V50ZX2Eb3IZDY6e
OnMRJjLw3hx+4Pvd7dxVnRfR3LLV/Fdc0gkvYsV72GYrdytUf6cFeyeTOF8owCVn
oFdi4x2mek7VCSc13GxjvCwCMq7d0OwcQ2ex61vAzxtq9YilSqsDgPMNGNzfIx+G
bdo+gE3YCqishLJl+TfbFsDOtaMgVcBjoeQwmTundr9lRBg0bdjXRvDHsldaLKUf
3JMx6fIAaAn4LGtmaWKs6S7+7cmdsZuisKBajodj4pbUGawEe4LlyD7F2I3V85Es
bi/QD1bpoFJsLveEyjCzcIk4z87KDLoQajXS97BcYOmpg3VDUQKLupXswjv3CrTK
/+APzCo7dWbee1enWNfsy5i5UKKoYF7kea+gmcfBoF9XUEAmoefUnk7EZJod2+Hi
kJLf643fMxX8t2aihzlZcjFrww9YQli3w7/M6O5pVa9bTqtyww06X0FoIPWCA+B8
SQCm2glWfRykmkxJgxqJNRMbJxSJL0x7WqRQP/aZ5Q+ui6MJ4b2gJDzkKh/WHaNi
jYomCkW4/rI4OJYmmPJLMr1o1vLykdPNK9wqj9O5rMqa7khn5JbwVqkvmFmq4gFk
zZzonNAqyfHElZ6JqJBi9SmVO85jKPl0Srm2yT27vEB5W29judeIG1+uOlRWqI/h
zkpKUzWNjePYp7t9F/zGI7rd5p3izgJQcDw3QD5hnL6HMW/Tie2WvhxOwMV/BpBO
UC3oi3ej8ehn3mVuvY89srVm3SkE+DEMYJWpRfxyg24P5IzO1lfgBDjZPmnblFKd
3QSXi4rq93HdMhVqnj87Y90opj6TX18zO9iMOzjdIPDHJzpFxUUq4TIIvs40NG5y
X26LZvi8WF5NziOSKPNcC09NI4vrn2pfhnJAy5sZQeQDH6JKeeoHKCyRLWVkxmFZ
4xwTDcV4B/kbe2qNrMlkx4AYvI7OOpMIjR+q6Pba7q98gyXw3bL+aZ1stoNy3SCB
WT400M3k16C6cMqI8+1KuBB2NpUARM2Qz6+l1HJr0+IxHqE4en/sHGK74k06XStI
hwpny8lU6r61CZeGeCQvPr2td+B3jHBUGngLHoU11FcE61ZF+jy2fraCIkQYo8qq
NJEFQpSCNZhZdN4jsuxZd2Bdk71DqVq7Q3TtsX1RecAsTi5UsHN9w00ou7cjN1kt
BNyE+ZQxZsMZADeIp9vK1EwJcvQD7J3hfxmSjkOe61Mj4OghWE7i4BiWY3BUNz6i
VfVQX3BBr2yIwx3lXo93GKRmGdoWxQns2JuL6ydie6yGvoKCrntaFG9QcUygLrR0
TjXnFopvVrvpp/YrVOAac2J+9JXITD0NUrP/++XmgB7VYUau8fKNKhqKVQfCk+Cb
+L5/Ki7kJAq7wDjWc1oRNH04NvU8QUYwygpo8z4UVHKYdrjWsm/0O2o7QAoBenHJ
bV/C/vwTzRHPdkdWBfP+TiyoaR3/KTIwy6H3CA/XiWHH26zt4T/A+TJbN8HMhyu0
2LahiZVbSUf6tdDSdqwoSuS/8gV+QVTfjvnTZIpX4qE+nMkCgpx/NZRZZDQKtjmu
dQOFEipsI+BKByk3ONWFGamClkVFqkDcO5wD8BsB0M8tF8VmSC1PLJDJfQ5ceI61
Dp+AwN9QIQauJEWYAn4fWHdM1R0ICEQ3jXh3ESI3jkPYw1TOjDq4iz/WXvBYtZ3G
pggh24ZASuGU3wgwxjHXfqmhHMMpGVbr5vnq5FrXMsC+NafLQ/OTAyzqWoghWtZs
ocmstvEUEIO+/2HieBekgfJW5XtEq2DWSeoSSqiHAItWj12Hut4E/i5LThwVdUdF
EtUBd16bQGpGPX1/37ZScut+YHaHgEK1oeectKj1bWVs8fjyEh0u85C6+LMJqzYJ
VrVodP6wk53OfA6SNbDZbzXKjgS5wVRhrBqAlwwTw38T/EQWblWdWoGqfTrpnUt5
rqULDpZZ+zEFluOtVBvWrHGesr4VreULvpzB8AMu10nYdqlZG2IBYRFWBD70j2B6
6S58EPLW+ehyCso8ckP+ujN+mKbHRHFAuhLJgf3DxKOCY+eMwE+i6juZvfUz6PMB
lsEdpaXstc9rxgftLywF49ehvR46Ks8JEDFQgjyqtVxB+3zuWxf3DxGyQz9JC8JH
Nfo4du54oqEHKCK5RsqsEN49vhNlPqcoXkT4BfIGc6dmRWbAGcQUBAGn1WIlEdEs
EdATm8J6tblAGPqj1UtT5OJ13iBtAHLn4jRpqzVN3YnOmS3JVlKbr423YNUzRbaz
VcFC5mAxJyryDN8yDCACBA01Go1QBS2uhJt/dG5OHl1UtiJuik4yM9KMBo0FZScH
t/UbL4RMskMXJd3GPHPE07zSRATRo1y8I554AA976DwpDeAr/TfbAbI4WLvI3W7H
XND6UwtTjJfyJcLl4xBEPWoeCDr9D4Xsbwqv8/RBqRKvf/UcxIEIWYG1pTrioJZY
7aAxvmBnn6rjNvDObTIeyyIOWMSzyhe68/KhalPqQDnVrcZV+Dw62Yrzk9JfxK6o
BucxR9Db3CT3mro/6oLS9wiESKzncbFEW+3LnApiv7MVAwOSCh1hnMqbjcNV1VCy
rTIq5csn6uIP4+OybiRJCqLQUSGn+5AxE7ge5zJAJxe7elXEbpUf6UqnB5I4mc7L
igdzTS6rjPRyoOeI70VJ1hV5g74joDrbmj9EuE1gqsLePCkHj/oDRvQ15hGIIpwt
sNGHH/tMbetaZN5ENzHx6/46pDMUXhu4hBMEDBPyv8WWwFYttA1RLSs2gn6NvM2c
St6FZu1ekJV/zeCPhT8ZeJXGkLsvakf0MTisl2Ddil8SZCrHTrZXNCWOFxjpEiuH
tZFrQeyN8QTCqeXPQ1bP3+apq+b5HBC7cHNCoe/tMPOkd1bm/EviZGW7MXJ68FRP
RXfILpEApqgWMuV2vJa76vjIweqY+NxYcjB1rTg5HAiY3vmirn4qmCv8m+6ArQjQ
/WaiV8S0xl1FXAf+C3VXfG7NYXSMe5Wmv1k5AlcVtGxWOMJFRex0pG/FtAp65iW6
F0a26K/D1shXRXo+jIX3PU+G0oUB2XcSYvOFXRDA7REPD+3+HlOBsVKCmbd36kuI
fCbZI982Vvgi5hrd1NkNIfqt29/MW0LvTdF/kTIxPt7vLOpSKvE4tEpZdps6m0o4
J3xvR8L+918ulLioZlAymliOx2nL6hFTxcPh2nzK+qdBZWK4eMFO3KTdq9WhYali
MJyruYg0gut2wLoQb1cX+IRAETzDrhUb+glyJve/Y1bHkHUZz0uZlU7eCkNVAp7t
AyeBM7LfGMSt7zVnk4A0rkufE657NPz8P4/mbBBjX3s/k9XERKpZxgTk/6DO6f55
kUG7m1IsX8GrxYva0RzEPP6jL/v7Mucth/bhsJ8+tU2kvcKTjKKru5KoTe/GkRgt
BrGUVGeUc4avYuyZs7PB0DxAg/t0o2S/uRElWQWbIwZMGHkZFwB0ms3KL/GruFbM
IB9klqSjvu4ojDCDnO3EihPFYGEQWdXPpjEVCaY6N2Iu3JlNsXSZshRwjhvWzBOV
R0wJr35h9C5PIElSViBY0hRITp1YCbi4XRp9YUVATtEKmy0MvULqVpxXNrbbhRXj
tYUAFdqvc5RjbD9KzfWIspoNnCQyJPFwSb7sVdsChVoL5/wUKovwHSn4WaityXyP
jxIScGtNiOAmAfkbpQOteYt8Z91Mhvhjq51VEzEIy3/gjkFFNnPPbDrJbNeNVxtZ
/EIO8+C7sftC8zjkydzn0UPPNYWg27qvIgDDMeKHcRpI5PosUfFg66DhAoTZnRGK
pnJUC4B+uuDqvIeoPoZ9z/k270T4Mni1oxdBE3LCXcGNyXqhSk4ktqJ3FZNm8dBt
esUu3uAC6kFT7JDXlMppXN/AZFpDwqO5sL3sEowE7hrOrPZH4bGexrfUaeihFbFA
0nOw0a/XFrUWToyy/CGdwTnIzmjUsh6wpHFy5eWN8wUwN383XnUK5fcfmc3OBbnX
yzrDRii42ReHy6DJ8b10SdkMynF4Ebcs7Yro4FAVQFXjW6s0Gjfm3zXt3viINvr1
UhdVaLzOmY95j+ABl5S4+AZPn77eaoGicKEi4zFB1TkpCYWzpF79v3rB5+9HTUDZ
1olz0eDoQ9KDLiM+gWgBHRxh41lpqWv/mjTwv0beqOtp4GAtYccTF7B2dVA7mECy
CqBotnc8fS5wRkEIybLdHF0lrBrjyfLSfo609Ky9gH2IneFhSPAD6zarFNlRa9Ik
Br6F50fVCtZDWoU2E5r1Q0NIF8aDyrJLWFirNF+UV9fNbiT+AQKuxb4+j6nzUpby
X1dsLDXrj4T4/xhgQTqXsCfQmh8zW2UJobjaP7/eMTheh+VUe+0vCcqC5jNtJt9x
+Q/cAsBSwZ9xweIyj0sBI/cdasyK6qwfAKc8B0Pmfsjr4KJkMh3VuNGfd0IOgXOV
AzLot2mgqvophvkhKcbKMYYvgHCVrgBdMesnx1ttRqYoiEBxVbP30MJ1D612RD1b
OM1sWsRK8NWKX04PDMV2yAipMta67K1oSChfB09scybv8xFL65xiaJfKnupRWgZh
XhMsDFHx26tR+55TnI9zQscVaDxTa7ZJsFocZWnmUEOwY2b2I92ooQQ1dCsMwaei
PFbTDOxhPbc4i8YoDB1hj2rXOVDt9h3HA5bZYP0z11MZRffm4SrwjH8yDNEzknVu
PC8Z3ZtV1Iuh4tm4/W+oTVt5bozZKjmv2LGJCIW26Wr5ihwAZLgqBPoA2iyuwwJ7
bHlftzxpjZbNjklJhtLOxqIxLw4wSlnjQBghe19JIGSpJeM4eBUe20WQRHH+F/oY
RiuG6VFu6lOTWyke1io/3C9B5hT9VJqsVF+ijVda1JwAoGSk4Te12KEbclamy5Q2
0xa3P0gmACaMiyLLq8YkINlV4SoRqwUxbSVmTL/6FoG1GU1Yv3I8ok4N9A1KsXDH
3Dt58qdhZBGiKXUJe4zm36I/Y2PV7ekGHTgsYRTxZWbajiD9RQrFUibBkbwbgfca
L/gq/OhhxGe7WasCIkTlCcX19/bdhI7mVe5t2RzfOC19BGOmu+e+C9quO2POWo9V
A+Wpb7wEsEfCmc0uQxvYa3EzYyJ1vNSwLTWHbAPGY/1sr0+FG1aJ49hLfgqltHIE
wSOREnlp6riVxJ3xnDGhzzX+sOqvEobuagT0eIm6oY7yO3oB6/CvWfx+bND0Gueb
fetJPY3Fq3a3zVH27PPPd9oyMwl2bwlO0IzJTRqfhWPknvRDK2lBRLwwrS4XBoHs
HImnu8dSe2kFUfPUqYJLdaQie4g4XLoBbojoZT1CCxtgqmCrX4J9F9HRSe/1ubBZ
2219YA1cPl1NKVnPv8zVbLKAvyt68CIvEWIbpazp6IgImAufhZoEJfDeEEpiEwuQ
Aq4k+K/yBqif+X7ChhaLbQViZGcP44guN85l1e3aBNgmHhDFGCEZ7O3OB+p0Pr/2
pQZSDRFW+UenvKXa2IhqBsVtGFsrDdumCf5++n8GN7EC77FHYwKTPo6zScHdrZiv
0ptXY/a9mYvFsfeSwaD6miexU0/7MvpER66oIyqylPPWU2Qeb2mkmiPqKW0AKpwN
42bOoB22WmtJaKjoMXUjB5PJideUgD0CF9yHVSEocM4JieCm3rCduybsG9aF0cdV
7gmHg/mEAkpioiK7JIaz5V31TYRBbKlL0DVtdSlieMHpYAqyW3smcK80wCwWU6q2
HCEQ5SoLABVHNrwLAwYnH39TjCKZsrtvO04ncHlHENhNzQK3mE+g6lqb6z8vFyg+
/q0MR+ZtHdLUJjp1BnPw8GuLNRjzpRUw8AujOsDlaSAaPyniqZXUhgWwuJdneqUX
bT65Mc2B/UgxDn2qcGFlCRjpsRflwKZFY3tJPvg4pBgDj6EPl2qn+XUcKzjkcFKl
f/jXYXVl6oEyydESuOlNd/kWIllke7aDCF4iJMZyfvPBg9kXoTQIkAclJ69DkDTj
4ojvH37J2ACiRtpo//e+Jh5KsiV/Q1psC1uV2Kltty4zF+7qR1iMPb6mXm5j+Nlu
T/TIe9Km3tIbU8suqOALx9HEJrw4RUBFM6fD4UULvu4vlItChGPkNxFZIYNHpHk0
Fzz9tu5trsc8z2k5J8B/UeXeGL7J+VkwGqnrm+EN23QIriE6+xZvrjWznkApSnVO
0MTe74lrALqDYpIjLz+xUPnEDjmGGft4PfcJKtl9E6eMm2tDTPlmBvjc0P3jL8DP
l6AThcG6JBI2rz/DZBywyEt/ko42IsvWIggyUt4hoPWr6Morz3QhBvVsz42jO8LO
ez7xOrt/GJ51/n15Toi9ne5x/2DdOMFsJoVZJ3dvDcTvOqtiAE5vyPh5JwHB1Jg5
ghTO5X5uqBTWWAC9Nxlm3mkRB21M6A8akP0qTCieaKm+AIN/NrnFJbSqJwG5HNRh
tDZvYmeImIUBA5yz10YkVlM+PLLZd45t6MJs+ONZIF9h8sOtFxf7PVbmTeJTjGcr
UsuOW3MzELRuli/CpEaOh07kPCg2W3blQWd/Bhjf5cijam1pnKKeu+TnSVx+2wbd
VpFQa+2ieEeTSHhwI8HRiGwa7L8qca4p9KUUBxc8/SJzK8XqY1OgegmrA6UWoCZH
vL09LJ7z23KKcJ8Ky6R0wIOrKmB6mShxN+n2as0AxZqiF3FW1+/Rng1an0sBkMNU
V3ESL7PasTSx+z9DMjKxZalVap7Enl1dqfRL8WeX5kQS4A8U+HJhlFVyNNMHWAJA
q3J62KeVkCmO/VW1W5p0uImkYe5UVon9cFZ7alLpHUjNU/sO3G/gNEjqiBTeNjk0
6MRMp8lAxuMH4V2VIVDEnK+A3da7tgtOPx7Tt9p20Y/PdjOpYfqf9becEAIR0u4a
Yh2ixrozc9B1w3hef9ksh6Oa4bUlyC0R34ud4/AZLjESs3PNl0Qx2XiE35GLgOrw
h6Tz5Vhbid/R7b6wDbn+DC5ssj0fYPno0MpGSYekxEHq7z/MhMqVjusWa86W9D5p
j+YCWzS/XffVeE5boVAiCMOmdIeuVmmm8GFs8sWqtNZFR8ZLx4mG3Lzf8glnqO5v
ONz1VnusXQ5LdB79T5ULeFrYaFxvFTH5SbF2bwbv+VcOId6xVbG5YAh0XSbpa/h/
g7JaNy1w0Q4Iu+UE6bj0rEcMv+CfNzGnVB/5vNZ6RFHsGu/IDULiiRmpXW9wJvP7
wWvfiJHC9NEnbJ/tCE5C1dLizxUMPzniDTzhFWUK0BIChLoY5UA3HIE0JaTTD0U3
JXw3O3hMmfPeTwsh+KK6MIWSpX6DEB+ejfp30qWTY7iHAPIQbe6GSQgNrVpRTZ6k
yX7GxAYqyMMr/NK9ProvlpXLIjUa50NBLdrRSIvZrPGwfWVHCQH8+HVqapva6Fqa
soD3HU69u7H+Z7WXJSMTTX8iWzwR3dIXAUpg5KJTtfEtuCbeAAzMK1UohXj027tH
cKOoX/Ym8sF/7aypBQPiU3OUTtrcCaqQAoYXD5VfjKQCKi0mXmPjxBlR3bzdZ2sX
1xmwAYwOjxuMEa2xI+KFwc5ADY5T9iQrwox1WgXkQBsnZd6q4LcXBDrUltui31+H
e6Uboqt9QAxmZUuDkQlQeJhrS2bGRB1OrqDQMdYfT17+BLOtI8SdsLl9R6rDp8QA
WJ+193XtQiJIjVCD29eLvd44GUPHe4qHzytp++IElnR8DlYD1m9vfOGHt7+iB0AH
H+sA77I/9yxGQIa5WtDJKv5d4/hN2pSafz3Al72ffVKCl3J3RE4meXxPKaXcwX3g
G/yb8uJG9d/Lza8Ij4X9gx1L5grzus6JoZi9gGG9F0Tek7yG35rcjabtoG4O0KsI
EAkBDOvM4ldK0fhBPGZFqaxQwpjRwN25e2Ot6DRKtitXV3+/U9DXor2lrDtzNFKf
HlN5UFtEsFdTdLwx/4tkoW57I9ck1W9CS3OYgpKWPCYCsXasP79ftwNSMBMjm0ht
FivBO17Kj8qx5GIQpjMvB9KeyXYgUNOmZddIqZgw2qR7yZKca8Z2lEKTeA1X92ho
LXLtDSM9hDZQkDtjqkv3q2eCZ0xt0vSSj010rTQXU9Xa/TpPrQMU+1fp8KRBVvxN
oEzM2jWwdgO+4SgYG327flesirrBBgfDg1+yDxyAe+QmAqjs5HLd5fgLqDfcv+b8
cyKhsU88Tr4qBKU72w6alY0j/bGl9Qpg3O/hQG2sY5NkWUhfhfNV23rx3BzvA1qZ
H2xPWF9x6/tWwlDbw0SAWrm3IWUUnnLLo4Ne0FiIUPSBEb5vMQGlFNoD4LycKx+i
DaApCN1vtNZkUGiQgWR/btFJ/luQgMCyCT48sjKFzAHLuiqavGMXGX6AlQGDqDI1
8zXd9ueMF+g6ZoQC8ily89m1Qox5IS6FR5jAL0b1JXsa0Q/aREp/HM0UGG8cAXF7
YTSKr6SgWA+sYJ1M20c0t8DLoygsYbRoPm+/ANprTdRkGJYzUkZn/MjBbatNaVHr
eYOeqdTjmbAYdPqBXdp0N4tPL760vgdgowVu1lSKPqEzhxoi1Fhw/vcipEaEq5mF
OgRTM8UnOoBwWBxT1flF2dB4N2Ez47ZdK30s5a0CQAg+avBdbtfPUvJ1eNMLWiLP
ZVHMX/EehFb5hDrGtuaGTG3qODArsOlcTn7xNKzX5yA5qFTCvgFIoO7/RK4yUcaC
LxL/W2MXWgBgKGVMgGOxCFlQCW4jEsRpOgiPZ8/0ivfKD+blRo2+e742jRYk2SZb
nkEA/et8hv3gU1RT/u8SNGPAGCh1H9G9jgx1TBEyq2yD72BC2tboN6eRl07iG58O
f0ZJoqIjSsOL4wxF3LHGiBINoqZ1yxoiJBZcv0rwDzzwveSu7NAbB9tbhCDsHlKe
p3jjFmc89FA/onVIJgfP09xozkTiY2NJl2u6HT0oZXjMlW5jav46LFUvJdh2gqiq
VEk4ZVrU9V3GeXXZ+Pr9WbrUvx4K1iT/zk+4NbhgXdEsXwnbs+fsBFIGojNNUilv
EwS1vv5otujNIZdyw8C4o51VO8NLU60lyi0u+aH4WZaP1dWjSB4NbBoZawoTLThj
vJKpEKSoxoeS1qkNarTaq0ifVSzmXwCtifZVRndiY0BbVcSKgVURlzwZd9DvmCe4
bx9/N91uDkG5wU9zmfSf6NmCNCyaMX2/B5GN1pNDgLLnvDnLRbYMwn6gOthLT5Vp
k9gAkiU/3yVtslAGIi4CmYoC9/5t1WJwTBTKICSEw4iveuFadnp1H5Oma1bETd10
qunSeGptHnby0b9m93rACNFnt6NmhRz7p8KxJzt3yDskJ8ZwPsd6xSo0nqzXh4PW
/mDY0rPFOqlmgs8EupzKXoyb1uguEUFmekOnsWSjY42/I+rG7pooGLD7eECCGCfX
ZVoMhNwz3ZcPpNUkj3Upvs1k1+kMcWIKctSLhMCxjjvOTs+b1ub7d4GRj6dW1DJE
BSc1DiP7VTZ/xtZf4E/yMvYzNTA3onQc20jUrwkJbrA3bmpFMSnwt0ZfBWMvooyv
vEZpmZotJXz0kqFgAgqMX/0X9hZxkL/5/uw212KgQx6xf1BwK+u4dd4dTcONyxnV
3S3tCcUWAcD12mM0vldoGnkx1Voj9qiiC9hBZdCJv2fHlT4AcJOb0PUQBu+a6QX0
0aDbvn8Bdj1jj0ow8KrcVnhPKZqZdWzfVT7OSXXLceGi0lDekPsCnoBWV55ReMMJ
R6+ZylIeeOiO3uVZAN5+WEX1ZPbAdEm200ff2SDjbpSKO7bVEmDEKBonQVH9ke8g
1X+8b2UAj9jDFBKRp6fcbCwNiua/O8Xw0c1UpEq1Oe3eR650I5l/j+F4aS5DZ4tu
1TWdHp/LMTGD805PsfqeQnWEPLGIpSni14mcxlrA2mrvFilBpxz78ab52ICY2N+m
icuIuE+ZlYszg4JNHqx7H5zAMjLBk2RnVr8b154ff3BMlNgVFdfnNg1kOdBN5WzT
U+5G0WDNuq9lwAFiksIoNh2gIJAwGgZPPbarHQSMyN/LjASBO/8IxVoNh0oCCW+u
I+DPP9K2M9YV/2hjZfkI7bcOyA2tyqGvA1mQkBi5t30dzakxE5ifeFs67ZhXvd8G
jMgatGmEb25MHnySd8lOtdje+vac8Mm7Be0WLYR0zgRPccWreGA/HHc0UHdOozon
eYp/44+pcirg3lV42OlE0JKULGjJDNgWUSibHCWFxZtUUPM3uDrrN87V40/bhYIh
7tMXNN/KlP4uDfr0vbrUfkkYkOY/+5DctMvyGWNwq+FxuUVfQdq5DwZoPbFtqTcf
b2g4AKfhVl6K1woW+qaOflK08B5267r1ctuZiOl1n93a/tPkgV8el0/SxWfMR84v
3JdS8QLPpmkxh0wnjCSTNSbMFLg8x9HtMo2W4Jk9v+scrGpglCfqMd6/5kH7+c5E
iJe0ydsPVJVSz0xEJ5sDWjjnzZExr8l7PoXjtCllhgXCfMy7OyJ5rq9Hb+zj3z4V
Jm3UskpBTqOs/n2ARVckqR96L73MGRNZDmN/AxkCMIOPfkkVlBcVsF5wjgkDBaK2
o/LOsOLfqAab07k3zygWcQVv/ZeSn+sIPoDaHicKEIj+kj1MPCdigOLb++QoUkDx
PNEPZBdmr/iiizcgLLGP/s15cxwNUfn8GXfBCKki99F4X5YbycVvGfQ0mSDAa9rr
G5JG+8dkU+jnIijnxKTW7gUbMZNdvz05K7INYR5mv9si/2s69FI/u7Yyv6COzPsV
0liTHRQ1s5vzysV6WDDCXMSpsIghlc08KZEdd/M2zD/sJtVZFrkf4dr+ysN/uuQn
0G58eTiZirh5gJgUROowRz0mzBeAHe2EnwUDH9RLS6tTwE2VpR4Ioy0YowpIO5Qb
bg0W6cGtaT7km5pkulJDwMWqM8G1hgb7zJetEibfFWpgPHa8zgzH3EeaATjIec7b
5mfcD1daAJ8rvUV9stUS/4E/KQzk1s3rq/Z/7tHJdRoj5SRbT+mizwGUdkaNiL60
LjE8kkLbgLWIqSSTB1JTrpbD8mKl6Hg3boKZxq944BSs2NtIFKymz8QT2NGLDmND
58z8HWZ1kwnBlIePqkq5fjRXPlVtpJ0iD940YprMDlHyYwMon7EVMKyq0+24rdzm
a6GHrG8ZVeaL+CHMA4vK03LLFEjGq5Pi2pG5WMVjmbzN6Hcy4dbAppresiWeBFni
hV/et3DS4/+BZJQ5x17RxGK4UPyPtVkP6z9GiZ/GK6K8I7rxShrsIe2oUU+P5Eux
wP17yqtHZaPQTf63vDVeW/i4wKgpqzrKqkt8PjTd3o+9P82c2LGqLQPXD9rlut5W
k/C9Qp+OHBupuBvh0i4NIUacL+lhEZotkOHYMiw28aRZoLtCZ6aDCIU5k1r4dL4a
cIKplWIIVfodYxtNcxbFoAoZWC2VCrbqN0XA50aR47O9fVHM9x7K6plz3wd5Q8yn
a4FF3gzi7eDnIX0kGR6oCd2+w5DMuBZvVyoQY5tEDcAz4ZbYVbPFynymLhSk0ejW
F9velpzTUd/1TqfEMEbgT5blOY4cXEs+69ZZy6L2ULvAUWBq2a8RAPh/h2vZeoNb
DZWxCS1r9eWvzsLtNUjdzJ72AEPT3bBRGz7ewip27XYi2G3U0AWbs97cRJ7xK8uV
a9AL1u2jH/EJoHXRD41fgtrE1BPrcTbZEcwSgwQ667Hm3qYOikFSFaM+2tYJb6Hj
FBSdRQicSw5MUCjRMP43ERV93Q/yphw9p8ZjTi8GNsqxZgPIhL35OFkGOPRZcCDu
/AErCCzmRmZ1R91eX5Enlp+BDgeQl2/aTLAY9Ctahl5zaQCt6//818YaWW+usjfv
3o2ntgoX0/D8ey/yOWvhBGZJmWjRWhnIZ3DQykj0RTCY8CKWj5EoGCAXS8C0afWl
QeCGnDpOW53RcR7PjWurHwpH5bg7Lqll0bwtZkubFxzjR4RTA2IChie+sSIw3PJk
jPtvm+EQ7ySYuXRlxHf+lTeaidmAnIxRc99VJOjP36uYrCMoJko5KsPGRnkFcD9b
Nrvi/5rjOvbMFFJ3Gm16dj7APaTTN/kvQxP4A0QEji4EfhwEkYLI+Tv1hw18E3CB
IVTWu8GnjCuTrvHJEmLbQVXqmAS0qE8g+XFLYDPvVRUzBACPHeHU8qnIGFjJcCby
ICmKgY58WaNwMRUGqA5sowxffGohSmE/dxGO9ifcRsgvR3LuSe1MrAyqksrDkkeE
r/TkHvwD+UMy/jphgtgJ1vGo5xpvi956sOCsC+Q3VFy8g/ba8QumOK5W6ArnahTM
fmsuRzRo6/CaswQE1r6VtlmInWr77bXM1bQqRByRr/nT5DGiwEem6+4O9V1Gamr9
nLeK6F0CSNL4MkMr5rcJJXugy/fcvLyQRmEOzi8wT+f1uIppfxc960MDiDMOv5+I
ZTt2ahXbKMgThdNPUvmGJjeXaGjEOmVLWS01+gUnx+gNdupXZAen/7cWBhQMcKuD
Gt/UbiGruI+yP3vEv86FjMHGaZ2TG/0S8sEOCIcDcS/FPqs1gsv5ogpVIOsYzkeD
ksFyMgjJs64LO30n9bqApSu2S7HxZpY+OoUBaeQBO5VuDmBoeGJaum1mhN0OUqhW
WpU5/lZjfm4Z/o6mwssnXu1IVGrvaJg/NgmJ/Q8BTzbfuRIJ4sJE4Iz7rexXGAAD
R47fxxxCFhXvhZHz0E3YSXwlnCLg5XN0kCReyMsGqA0he3MEOezxVL9rgtSFd8Yt
7+U4pG+oQxl6tPETgdH42Zbk8jXi0Tb3tFFfJp2TjlL8KmI87DfnBBooWP5rodWM
RCvXiD6aX0X7eYGqsGGsMFaxLtTAo/BtPZNulGFoo9prrqJS9e3NrJO7yWd2poFc
jclRHDo5++iiZij89lVTgenHwL1Ch/AT7Plo+0HsaYnDm0RI39jGQCXaKGtUM7y7
0MINMkdfpoE25/lWUNnjiLXbcWBx9NWWaLVZK7MNtDh5hIMRz+smJStWqa9VOWO1
8nECY8nUKxcZ+bplkIHb0fNesQ9e1EtBEFlBau16ofMCTD37RT4rHOV4bhk6zRHe
S+L7I6/d6tJRSp9gDlfCe/3t2JXyYHmkVR8vMonHVTfN7knKG3bvK+gwupiu4tgr
jZV8X9s5ysy4s/a4w1UMV5Eh5hILbw2K63VPKnowiUp51tTePvnuOkuurxwalNu7
96dGAAWzW++9/CU4hnu4bIbuC8UUo+3xC1O8OyU1W8hV9EBf3dnJca7YmH7PVjn1
sI1Fwtu8WwmmFj6ICr/Gl5Zu71VXtrpZr51jVhmNQOvTMBtClfqZoPV1mc2wT4vs
kFoZ6MJZcLScfb+5nLrPjUdTrgWvSjxQ4K9Y5hcitvhS2fQPXi00jeo2XFgDgaW/
ysR6xNSTaJoizEdkyX5txTAmtWOXX6EO1zuR+bq94SklB7x3VOtQEST+pVBBWiYw
nBkrRo/G7xNQeR/rVALR2WhDlJBH3IvSRaD7TtgPeNc05hN8sXxysRpoRZWct3AH
iK7jAI3+XxuZ4/meAU/ti4iel9I3VCqF1cgyk650ZrPI6erEev7whYcTwMzPo/Ct
kn9jOxUAayyt2Rjeq9ElFeFOY6dvOs2Cj+WV+bxBVcQPpaz0PZGz8TDG1EFfswMW
v9Ni3QjpbNncB6XNftPr18vA3YZfJaP3wsBWhKb6Yt7aREoU9ZzWeLv2MABCLM5+
sseKv2k/SvSlgioX6dkTdzh1sANaUDNvzmUmv3cBVP8EvXPI+ep/O4bPq8U8JLQd
ddFxdfQCyfFPahp/epl0dzn93vM/3EoxXlRsVx+GXTP86GBer2VgUcCChu3bthIz
J6CsUU47KdUn0x4URpAg2rozw8Lo6Z4C4ijDIimAKinFKMKoFu0Bc+1RmugeBc9a
xFAjuhcps9Q/vFVIVNDgu7PWocTQ6j9ytUdvxdSU/i/ExDsFX1DVXKyLgo5SCNod
zLvpAAq8VrRPlHlLeOPXoofwcfLoIbLgacHNs8QzU+MskaYe91vdRSjP1D9Mn4gS
S6JESBRWDYaOFBIDeojGLbi/KntGP5imNiDlv6yJS8dsgVBAbk0uh6ab3M/QvIiw
++sASXKhqEoVOzcbLhX5QSs/RlP++8wiinXSHGdbuIO0PT6Pt9F4hmItWS/4Y1Wj
Gz8T+eyJ0XmeVoVILVbsz68J6se8BBMk5/PJoVVIhcMvR3m/5aokxHLY2VO/J6TK
x21FmPQGBXaQLDF4bVgP+EcuDowDzgdQnBcac4hDoovGASp61jTAEJXCY0HpV0ej
l/N2OlSh0wPxzvCRkl84q4qtu6Yyty04mqeu2s+y5Y63mBTVOa8BfxDRG4fuJ2XS
ZZ+znrhHnzdWauR5GOoG+HkaiDEuTT0uufb5m3wj+mUI+Q43rtZlFfv09thAN+sl
MwYCPRlbgoa6b/FwHXpekzhl/5OLicItZ7jbS3miocfKnNGP/hYUNfJ7RvF29ztQ
gF0/5ZzsHC6I34rBQbkLxCtk+G6GJxjGrAyNhFc0uU6ghEh2DMxh31VFdA+uJE2L
ZXtEjPg3PyHqzwk4fXnYKv2Pr+wyI+bwC8fZEf45/tM50mnLc7+K0O1hpKij8M63
ECx/cZbgaK1qqUyEbaRxlJ4OPi4bf3mIliobsGkbjkDWXrULsqbSUlGnen4NWHYv
QjZUwnjxVxoq+0ond8Q+K+vaMnB7UF7mDqsvTs4VGvMYu56k51eBqT5CLGCB3khl
ltNe382uKyrYo8Dx4kljaPlr+UvVEzkZdmIzX9PJXZ+HAiqyV3KfzcawGX7LHhtN
F2cwdnpuiaJPHPik8s5jt/z1c4nn8FIVlqT8re/qCnrV00go1/xlSfw67eFeDXRM
YL09caML1aE7Nh8wHg40GZBVw95C9SaaHD7ghcEJTf2DijCpPEpLHHMfyNiyRAiT
cZRy16eNRQLNEHEfq3hKV+6Wcdwq33vedRCKYFgXI9XMyfqRVcQaHwvyjDeUYJpN
bVeHysKt0OfRr6ECaQEHKXEl9EyifLA865G/bz3IJngUGYLF7/jNAapHtaaSDTOz
mFVx29JSueDu7TyJrKeo9wu2QtZoVE1Xm1lTec+kMtULDd/WNc5NO+IJX4q8nmmH
s0sSkflcIbEFZN2+X0K4/AXBTwhce0AoqIkAYBaoRfyq87mghJBgSl7V1wfO9W4P
e0tdG0nPi0W8bN9+seBP5MmqBGC0VcLRIvwR4RrCKC9skSN5V6chFsfuxsMb4Sm8
v3rD9XCpc56PD3cysb3ccM3nf5abbQA5ei+aaxgEWWig6T5xUBQsOW8Iwi69K85D
QXlUBtS51/F8Uj6NbSArGW0BPuIwKbsOGnndxojuUsTtLy8+6MO29b6SvqtoPJvg
zbO+PqHUZf1ABEWO41HctmyDkyorK6Fq20uy4PZnwceWRC4Q5ZM6MjR2j6TFjalV
NyZC8xwSOhZy0wwvHHclK24I3ZZzSnCUzl0M5fNGgTVC4R8Lt1SsGuipnbwiAs+B
BZdk8JW7osgUq9e05ckot0U4I68D7B/OjxyKSaQE8bp4yWVbHj4AqxUqGlbcK8XF
csuGMExAFMZEr+qKT9/Dismwcd74TvOYZlnWppKcx6eDd/4cKsTYzZAw61tyZ/3k
M4gS+uWW8a55jPaPGnqRVebdXgRLVaSCAwNKH8wMiK9tAQwbgs/u9DeRmdHu1/ff
kvhpYmbhwBAnWHgPTddsl9yvtzLr2U+RImlvntWtzEwynyN62IoBfACV8RDtRSea
oWmbnKeM+Kc3KxNYLGd3SbPQYyeTEGP5HZkvvqAC6xzWCUYr0RlR7YC82RxBs/Tm
zNI1r/0paCYPrxUk/9qHyicVjT1fVJCH86F8lO8Q5kTqYf+UYeh6V3G63Qz527w0
FwPmkHP0kh0APiH9KDPTqpvYt6Yc0K9f3L/H4ukzm8JCn6JScYPsdCAh/rZN92Ao
ZUi9ko/QQDUtJ+Ny73w9h2YB5AyxLCvxPFF5rSNxfO8d8iKckHn19zCiFubvaqxh
hvsahi1ejXo37Jrbo8m4188Lh1pYp+Dc1r1gV3bTjaoiOQRf/CqZ5c5uUDQcALMM
P7Cmt0L9UPCphEqtHdVOzhpnSmOYA4MyErdlYsJxv4eGtfj3iX/k+92yRItZmqHZ
FdCNxDmCc8ahu4TjtXf0COtEumjkyk8R7ymUG42stmJ3OP/XD2zPUb4uyEWqpzOi
mlhbgA7G6pH+IqCTnIP4gXU1491xUUvTbrr1SC6HMrVOxAqSQIB9+NmRdZ1tzlAG
GbIL4KRYIs9sDLsixcJshb2gS4wWPonyL64xSF72V0jCbikalentDNuRQjJlXlgJ
hdLAAR26PpgLzpREQngLRq+rKTb1nBM8ydLnDLQA+7IDQY0aRMUgrzB3UbyvAsqR
yVjbRAc7cD7SC5pCQZEdAb0vWyDopprbu43VC/Xn5GQaANzB9mAOidNClrjZ0z6v
+eDbbRQFPt/yr1zAuJGcqrRuaLfRt2MskO5nJP1J5DXk58h/tLnOSSQFBDvo7HoP
C9K+S5P5B2r5PMvnwyuvCHISddRNbiX9G4IQgDg5Oif1YqSxTRC4inmP1NWCSSeO
nDwk0io20EEB23rMh9xsesAQprnyr8XbApAiWpBb/RrsKmSzePSzu9ozl3kkCBHk
fjnkeqjv+twlsaipJFmHKpuoD8iyCA1Vr4MLk7KhBxfcLHaSXWrPa3u8Ogrg/8+E
h7W/aKhrzodOsD9oPq0KjUxRsxDS0gcjVnyFGeSoecfd5OL1NarHEVuH+qZqRkHo
cSvu7X5x0ozX2rfOhfx+NkOTdlR+CjR/3/zoXIzR4zD3mh+tPU5bOdw2ymB5beX2
z5EntmdScqbr7pWVO7c5/P61X4BPypFuxVlPW462hy/Y2Xf634XTegT1yRhtk4l7
i7zhaEYMVblMMJN7B6YMwfLhMQICZHgMz2FTw5WwHWweVxreS7Y65KHsgddIXtoW
FLi0yUy2kyjuzUIC68+oxbtgLHal3HnBhJAJqdjGZNWauEjx4kb2noHPL62o8sEy
2sGbdTsT5kdvIEirAmfeExnIlzjV3W1EzP/LgLxZJdKEXsth93IJSLbxHsST5OPY
TPaD8SNkQnH5JSE98tZCb33S7Vu4JdS/AHoAdCLBufUg190iWsrxMsZn2FGCFaHS
o5tjFzJc2E9NLZ0lIKnOdwpBx9EIHH44CNoK1ixDzXkILDKgm7+gaJ069AHOVERa
ygcTqv7zs4vXDG69wYhqb5+PE312GlX6whGSNpcGr7njpZmlBfye7Ca9Qhkm9KF+
UbX3peW4Wh5J2hvuF/h2w3A4SQFbsgspKYztyTdaH6drn+JIgMM12kadFKa5gzOA
FsvcrSJxoUAPnFuoBxparHgn7yi5mqG6/pyYZXlfnpYWfLRxgeUO9ywenOj8khs9
23JTb8uGQn6fDkrp99lEn6WDGZl+1nJi0qNNkrEAZDHBDQt3FQt3aNjzYJtb/X0O
BYT5qKP8HxHTpm5QNGFBIV/ezmAjLtJtdLLzAi4bgMuV2fnMGFEZf9LEe+W8WhHE
m+b1UHFbXKKsbQt/etzPxiHHUXIz89IV3jMvjHnBbAy87t0xXSz+I0GjcMiN6wCj
jxTwLckx0LBLCKEXpcnurGYi2LaZK0I3RxTAyBjRewJ4oJv9mN882xBALwMPdVkw
IjpiCQhTMdXdOUscX0OeIWkV3RZTfIpr1KGd81xrCq5QELaSAtgMyLYbLqwEQu/4
4/opQo8W3Pzu5QO4DHB8Ud8vzi4UFslT/xX6OqRSn/iSdxqfropmbfvE5wj4opVQ
MRtV5bIU1ulJyqlIp6+ObEg76sZVeAXyiThi/KE52L5x3Mul/gTUn6Pma+URYvCg
qMwWo7Xd0wrS3dBEvtkNvdXozUJYrsGuxruMXU2poqISbUln7Y6TrRb/2JXnrioI
JIxlgn7DKw+x3ggSJlrrHlwjkP6BMs4i8Gn4eeqCoIGgNO1G7eacI6kqP3d5UvAs
f92SbYgB7YZ5qUB1Upd4BA1x+bAjFoGetxAjLqwa9kR9hC5U64IbPFZzrjsOV/1y
JsOs/fIdcQ0OuFLcvfSSzzlfgbT3gkJ5ZU9KPdQglcft66x5h4O5BzuPMVyy9Ow5
FCUi+p2s+n6T8i9h+O42rGz0EZNNY4/Rh0b3iONC32grm217b2x6ehwZFQveN6Hv
0uonfoPY909rX9WOKobR/VwirLpokSSUh2oDYGRKKV3gPuumD5xoRCP9pJE5wW1I
WsHt+dD5z5Wgi4BIH3/9eo/dP8fdzy+ZnlUnX6bhVpej/3zG/uWjYj43crxidzuE
b9wkYNPZnTywsPkU6Pqzz0WDUvPf6F15txSmRU/gqqLi69sd+hgOMT2z6PNSAaNB
ebAAr8234iKvHc/OCapGx6Kzp2nUmUnslZXQ+6WO7UyuGHkhb6/k9yfPphEgzt1L
bP00Lsz9zjJOl8qfHPZIWrYS1TTXbnYghTnVuu7+M/CNm45GRxmrl92Jb0AVdXSc
4w9nJFE8tDVIIRWnscFdPgbFf91pJzgm2bKIM6+wG9PGTbKhYtTc4k98V6DOlZdh
XPYGtCWNVkuoTQXy22y3GMx8KrJwGhcfivCViiTLCrxR2rq4qvvG4R22+P4IGLNM
b+J9V7x3z2KR0lsdzCsLFfk6DzqRsi4/D8+UEcQ3yo/VBUu5YRNbcL/kip15J3Xb
fnaKrzJNqlXE7mQeEFdNKfWTiJBtCd6APPdD176Qgq4hTENlKErVO5dmUavQLRyZ
KqYCnZrhZEwIpe9w2xzQWtHyJVzbplYUE5kA7uglJOv+lMQpvNUkx1jvbhj97K0P
3xRmV7ndOG5WGhZOE4Jlp22t0OXaXqiamqbj+vDWlGN+nMo9hJIoP/5pOsrfsWuM
4RUTI5Xs6u/FmRT8XWS6PB4uMYBtZF+O5SV7QpEryQlaxLvkqrx0dT6xowF0eS8h
7/hkzS5xu+/aY2/iYUzsCBM7rJMNhN/siRVu84LCbaj/BNR88lazQIFbpDv7PrS6
CghqIs4ZCrQLaeF/jnl6miMGlgUGtnQQxS0uI6SjcfVwZNUOV+aLVcfA+Q9r5QQv
y1MFbvLowDHBvbnWwMeozRG9ZO4xeBsCh/8Urau8Bncgn/CYhlQK35n5AGyfqJh9
Nokiwqf2vNOpXd9RWIjzWtwGpdpwVwE10hpykBiPLpV1kpeboylPpDZQaLjz1+u2
zp2f53H0NMgYDNTNS3Z+dueXEezDzl4eb3f0aUxikjt57APNSIokUK1HbiBDffNK
SEn5a5oRP9AFoXOO1FyG6NLZsZvJGrjKcPnc6Jdl2KHGvIWhTP7GZpsFzutDIs5W
HC47bin52pSTFchg+Za8cjxm2NULMXDKZAwVMCiz5/AD9hYUu4c8+Mpd3my6VemB
eQ/hPRPNPjXi3++0CXGhkDkSSBbLOSoS6czAX5XwLzI6nnA/Xzq0QrBpEpEnziEw
whWAX66w8WboknhBMGGYZgp3Qyp46aBy01ccwfZrKn6dRRvMY5Dcle4uPm/4YFcS
XkZHbInaMoujtg2Lm5othX80HQowuTBiEZ0InAAgi3M6z5wO+Bg5bcuzniFUo6L9
DRdcA3app0/NQ6yYBcqgApLXwhwWbX/QGSgBd/1QmoIVd7Ak74bThxEfsQoCq784
frPokAi/BsfMyYvU6xnXHgJJfo6ZNwbjZbNCL7ZFp0ER3xMLObblNua0/DdEwGeb
MMwPflCk6fDwM/yzwlQqOEOdi3jAgc5stqBjDbPaLiunpB7EtWpTAKGINkbTMe5g
rkXAEUNSuCbJ2gC4baYS99GrpIuelocrU7KXImRpBJqZJQf6lZuNyT4W/uvIyQpo
DwjpCsbDvQbMIg3OGO9cBrpT1o97d+wNgnR6ISPoV+5AD6aouqVtm4MXyAhIh7ff
alceIifozKZamVBqwjvAvYapYFxuez8/Jt01Y/4uyNFyBm1fywwl51Uv+7Z+dwqa
Wa0ITb+63oSuW8V1PnqYy0Oh4aExrwl4a416b1f4B0ute+kLW4fLHy6wsyfPbAxV
ja5ZeUkaRUkDV8+QAH26xP9hbd2asb+ndKFkiuhCsChv5xKzO1yZ+6u7w/5DfX51
cCbxZx6Yjobby36HKluj77v85YlzICZ+6Udm8ekX8smmk1YUb0xnt7bSJPVbcmXe
FxZkgCISzaRsXDe3yNnOSeLfCMK4U+wjJyO7oJ8Ah8X4tmbYTF5lEeeFp3cMhWoK
TRf/mHe5gSpK991ukrwzjGXg/JomqNFYgeLnLEm0/2zynq5tX5IKn5bi2KoKhaCb
9lapIcyHcb45n/HjNUY1bKL0MpPszLeeuNwvQvJS90GpLeKEIIjwDi08jeMqg5gY
J/CkMjulqXI0FZoSsDFtGhg9pqZdnYZC8wDqyE65XwSd5lHGTROnzy7UKEsHylii
i6USRI/zPgDq9KiyOElLMd2elHdtMWO0/N2EXp0ujyghkO65+/2letgyUtJXSb7f
xHyFvykKzFRRJ5CP7eMjeDqSYfqtNTsCq1KPV/yDbk+QFRJZ3pRDA0OWq7BmcYvE
+gHDUk2iDv1qr8N3y20t3lVV1bN3hYeluWEVfo1Jnqk/rd0T5vg7q6oPVW70ByHA
2/S4iRvRbcHguoWiqQ6c0bH6yA1BZsLZXvod6k3Ews9UCK72OuU6lJz2ck/LX1Ml
PDtVlT293PUyEzFBB+y4V5g+jKGAZaGfZC1Pr7+LlVfeIX7JwW/nccQ9w41Mygow
Mh5b0yp+N4P9XM72fhqyrW3BpsNJ61If22huo+UGaGyq0yI5dYjJBGMskFpmKDw+
q2PyoEyXfw9A1MzZgpN922Ib1owfiAa89viFcjuUNgoD3zP7kUzD5aThhsi+POhI
OsD0WqdrZV27cjSrlTi9m79+OscbzAl1yiLEjTmyuCdfWNJ7m70lNirSBvicASMg
gS86capelMhJPKon8QM6r/sGd2alf1DbDj3Z6YhjotWzVf45iKYWuodyxoixyGXX
jspWvlRmiVMWz49VIs0uaOpvaubD0OStm6KN9gvsmLDVdQT0igPbMfq59wo4MaI9
yZAXUxKnMofoId4f60EChmr38gw7NbRyWbguE/mqfFE7vTLFj00uF0c96MuPG0XL
42S1tHr0b1hvpMWCSmWPfLUJEl+F9K1uAIgL9PPsZVJxGXcR3HCSdgUu3QOeC+TG
3Aeos/k5L27mnrgrgeVAuaxH6wn2/vQcndBvAmGiEOo+PIzQvRpJg0LHEA9ysP72
wzPIVfzgnFAVuLy0McgTM5SxDPENBm2e0lE5hIPk1qhQtZtLVYG4rxpcae4+EshV
ecixFabVwVKDSwmANaDlfMmfChSt4diCmF+v/kUlsX376onRw+SKRnD9wNf8nE+b
4izoX2bsNdqiQnz2nvaRvL37JmLPbguJxqc9NP+FpBEJ53s0l6GvahFAG0EJE9M4
FGLtpgd4ngKI0JQjsHBO7iM6JftnM3ftPaLOnwo8roxtydemZF9m1NjyY3aprNNI
u2VraFDTsED2JF+YYjhPCxgs63bpuaNvw3ezG6Gw8uv/EpKHz9z9BBkrClDbL9Tg
jSYX4wOJiFzrzg2q1YBXOe7yDe0ZCrPA2L7gnCW7g4ozJsvi96XoCqHtf8rNGb3+
VNaplYwsVYbO2nOyD1/oOFRFAoYwwpzM9ujZII4HUtE17XtMKjGaG99plRRAy8q3
S5Talnivg2GHoOVQV90w7Dtqj3NhUbyxNBcnFhwwE693hbEZmE+Whsmr2gB+7aPZ
QLPNx9ZkEULckSkLHvg7ZHxRbuuIIh8ie8OuLFmB2ne9dMCRoq3QgEklSKGr0u9U
svKwV0AuKYQnI4YDZF5gsmH0dd5Z1ehXIUOjJTIlnKBqEC9Qk6UlGcNtXgqUQl74
bN0xlnUmD1YIngzfzG/vl5VaSobZPvTNLJL2kuTAAh2y4RDdLDttaYGV+8/B8V7r
ZNY+6GgunOuAftkGOQoSQh4OiAWSZb1LlkvKR+di8BKEeuk1Kt5eqTTqoNk3RUYY
ffYP9YQEk51kLx+WVSq5LQ6oFPlgf18OQJSnErYfmykWs6L2ycLEI746HP0VZj82
cEvf22u7G6GyhzNsZ4PQV+HOiS/WaconCL27Uf/ZCUoF+zx8tHj40P+W2YzZXiQe
A2kR87XZbA9SIvAef1XtN8HL72snryOtUdcY3labi1fmYp6VpbfGy8akQXD5cL5V
hy8HO+RXnueTDoPHlNO5vSEOkGZZAL26nPX5mAFGB0Nk0LjKsS4qYM7cGWOD0kv0
NyAwZ7Y0VgvnTb/6N9Upz96KYYH87RlyfqLOXohrOOayREbR+uzskzEh/O1EcLaL
ypejzTxJy6hdtYGvcbq8mGMbNRsNdhp16oQZ2Gf85gw5jpWc/mDGa4KwptITg7u5
lTPxUOyCV+apCkgY6ySZ5ffUBSTm9G8s3WJksXp7gbGt5DyuynrtPu+BE5YScPyG
rNdPzyLV/P/iA+bba+uJks0wK0xMj8a/h/ophAzKP/OlnxAgYjRPKwZmfiRHDNFm
Id4ongj5S1ucd78ytdoAsoEocn3vS80js1Ml79n+kUAX72zIVhO25QJkrtx/SXlT
z6j+S3O7cOh/FnuSiaOZ0eBwe7WnaTNjIYp6KSTdgZXLea2lLQYtWM5XJF44rkKc
SiI/EgQwZ6on5wp7qLfxz9uaufZWh2ujt/+9WLUV+6H3sxbx0sygSH7BhVVdn//U
LbbrKRy0G/7BUHYyYxYCS/yftI6Xcj+5miHR7uzq7JimTNdQw1QWEUpkkY0ydJQS
muaCEXFrj3zVxmISvRphE7nPH87pC4tuSqeoNbNtbAtqamk3zTcJDXn89/6ihy1e
dUnP/bnek0ANJU1J4GNbn14pxihTNTwNg15DoT3nU5DvG8gEmyeQkDBfRkQR2iQ7
dsBFrKnJPTPYBWIIOCYcL4o++iEBurCKMODvBzjf9wxkSOh/OUuMTWSIQ5XoK2gl
NOJiAvDFg34mbM64Z76By+4ONLtd5MlErzJmOQVCA2QT9/W4vZ45arN/U3h4YJHN
gD0FIChJan2WLJaz2o3okvehdBJHcy4DU1ge/LaNV7DXAUU4Qr0W6YT51X/yQ+WL
c6aW2iOD0XL2TjhC7NsLtDSR5OP/AhZ//faQ4BNbVO13FbOJwVnC23OU5GHm3itm
MhJD/1oRZEtRix3ywNcTAAGDP2HLVLC2kCEcblPRWo+H+SLorNsyYbtHQsxzuE/+
mZgsD1c/ije4Kl04EsxcWIobjg8B9r2Umw3QRm9I+G6XJNwbT7bkXznMiN9OMwMB
M7/8vrw/jiTnKhz7cD7DNG5Apshnf/EC0Me2gIy0U7E5nhojMu8hBNqoGDdww7aA
tqL9MTRYor2eKq3XwSGISWsaA+OXNW9ed1bYNHotV4Us2JeSoN1tGYJBNqX6L/cA
5xg0s8vTl7f0jd5P7r4LN1A48HyS48HKtz+M6xowJaVg2EnQnem8Z7oR42NeDIiy
B/cFMZkDJ3BsjOwmHnMaXWkPzKa5Pk0TlVG/VTIHdlYRhkyybkzXsIWI3dy+SDxA
0zgN+1lAkSr8rr5kjyZHbdZrSE9MBs6j6nOgn1+KE+beW1eCgLIs1YDelybel74g
DdoEHphmGtjVSe+2yDEm8Qi2W+fYWr1vR7eoz2g/DZzEI7UCCA+CBzVyQo81RdnA
Js5Jxo1hWOfs+Pt7SdfyGGM78DC6NKZtUQ9u7rLXB0jSQt4ti7KwDNZxGUN/7+l/
nezAT5Tia+ESdeq4K+W9roxzKdbcqPM/5H/fDuzs6cGW8KrzH4Xk05O/mbkpjh7X
3OSenNsjuAiKhhMF/uVFwQgW+DhLRkYW/bgI0Q4IYKg9rihOKs2wiCXtN7ZTJ0yY
6WdaUA75l0tC5TMZV2D5l0D0BVndCj/WEh8BWoSxTJku/+POL4Hsq7rQuu1qie7l
exeCFNkzGa+AzJE8vZ4wa6LqDBwFJhoVEgRSa9dTNJ4TXn6nJGGAr5+NkMxDbAhx
thiIox5JNWgemWE+5lpBNr7fMzxJJDCXCiOelIQpEdBzfQJweSx+m9Eg+NuHhlAl
n4QLlA4bOtWZVF8+r+mYK0USu5Inq5F4/fj3PB8oHzUOxBztxNKwEwUZZ4gvJThH
VmhbliF89W5i0jik6z1BQROYEhrmSBaTeUdQ6fUiGFMKzGmE0jc2QO9wAMCC0Hmu
u8KMmL4JnAKuMmsPeOD4siuXLaQkLcR8TQUvnRAuRywKmXS9ltBpSYbCe+Fvg07z
qpdomLHlizoZI1ZPrO1ufgvzd6YyfzampSqKty7cBoLL1owI0ZLeGSvc7oG6p/rP
2IsFsAfh3RUQZlMmaGzYv7aQ6aJaEHUd3n8DVt6jh73TmKRAd5soxpqwp3y01ANK
Hed1ACj3gmE5pCSQKEHdokzHcoEzv1N4BdD2hu1s/wFWGIUt2Yo6vqE1Kkvhlc8M
xYyivNuzJ+eAElw0jG9b1sasEnkwkd4RBBzLTuj2Q4dSFf6Vwe4b/RFoYlMuHrGt
VpoNk+1y7+M0qbvkshfW7dmKtCHLvFJgXaGyU2UIZEJzsWynsXSgHYViVbh6usSA
syjTEIJzblWNRERY/s9hbmArYJLlUT1Ug1zGpyEiFH94YYXE/sReBwNgrzIJUB95
S6kZCNWj4FroLGa7KzxCBunapXQJrM0maqmRGsJuRvcw8kYUjC7NdPUzn1Scc9m8
k7r7Hwxeat9CL5R6obCs9pFiT0+GeWPysOcUm3tbeDy4wL9ORY5KJxdu23ENXDYD
dljAWVqN44UUYNjZuwixu4mSBaQihLuj0EeQX24618BajrMMfiEIT2ZM38LRyBTr
QUbq6SDgbu/440i6oVYkSGFK/LWTTMrK6OegCqShFAZ9Bt5VKfm6dJnnwvKOMEtM
PnzUIEAVU1tqOsE0OdibR6OrEqQink18i8DksbgYRTWJOlE2CTiZFtp9KiBRXW1O
Ur4ltwU5jkjuH2hqo8igXMivqdGA8Pcz7qUOr8bUNVAia+S6CF6Jox9UhS2AOdYq
1Xok6UFLt8nuiE0hUiNaAXapIE6gnozLIED+MahqcM/RrOOjo8IqPfpznRAHMHKj
W8zVrc0av1m36OyEn5UkmY1ckDULFXD//YDE+pWywbLmJNEwYNL7LoyP1rcatL2F
8eHQYybsBgtUmmbcbitb4o+aJJFwbXF5tSVkq1mc95t08wSS1XeSKxeBfmuAT6uR
KRjDP8IE2703y5zjTPkM6+pd78EsPiIZ844NJDEsBNMrYNUAbr1tvEtQhnlC4SRq
4NfcEq5jqTLWE0KSrCZvaqO+8xWKqmOOTpi3IMKSSWcJgIIH3oV7N0OrTWWAJPBK
scBb3mZBxXQWFWwX+nQihNidfBtDzhQwJdP5qRy85tvPW8gpdHQrl8NG1/pCOpA4
loK7lghGtzWZkSY8y9vQuNmkOZVUxSi6hHH2xiACf55Tq114GUc//qjrsEaoTQXm
3AMZvG7U1C5vUEFk90vcK3K+4g3CHd3rs3MCNloRcQ5ZooKm/8e6kG4z7gXQ2ChK
F5y191CcvR55VhGLetWDlK6gyDfL7LRFhFijN0Rz7KDdlUnxCrEvkVcsUFo5lXD6
gmpXjR9kBvVcrUAEM+jGB2GJu15O4WB1qrUvzbcyVX7clWwMlqu2W3pmCNMuppdQ
mVZJTZdu6AaOT2tmyL2KLseaN+2UAeK2ahs/KgIZl/wSPwmxSQjptAPoDWvAPyf2
L0nF7XhNfOqKY0sFd/ijBRbYGQZaacmNtap0Bm8mje+RSpCljgXFUtgQ3NacP2kT
6owfD6JXRuqEKwO8J2+bB+DwgFzJyqLz/yVuaVdWghUQR+8SMLu8yZA/FM9hdw/H
3XEkyhbNJ6ZwUZO5b2FlEHeTIIUWh8GsAIbm+6IM+dTbq+rpQ2RQxa/pFfS38iWk
xTLiV96LoiOfbkzUFKunF7+iaIJxOqitYtFhc2ybktvX2cbvO0GaxgjEw5gr4QW0
xQEiUaOqtx1g0zP23XW9jHDvX69cqDYQtbkFu0zcdkNvTSj65bpiCP+5fAMF2hpF
WBQcYyJXL8ADLZI5YvQfsDhjjuj9xE2+vrydfMUWdf6CUX7h6Pviz8zkdTASUlsj
RD22cMErHB/5XyQRt6REC4ksULweysXKFLtet/W3LfdrpW16DAnvYtQ/BFOzh7ir
h89efQ/ScQu7beZ8T4AXtMCj0RVh0Km/SQSNxHENMJJf6D12avtg6SOS0ZSjEtpB
Gzrk2ysN2p1tYH0MUsqhgwKFYBkzss9VrTta49X9zgeKWPTzdPj/Z+qyZR+Ud3G0
UNtWCbHkjAp42gAvmk4ZEcIbscsuxt+Otv0jOtMAQEM7TrftH2ep4Gtu9yYc3Zc+
qeZvBdUfQeB96XyaaICSqACsFkQYD6UGIMbq6hBQG0u151+jc5tYAQ2zTr7NnzOP
nhL8ZpUgQe20j7aFhFmMeDs90qgIhVRibQVdxBGjTKUnhYSmJsVAQOR1ihPXdgLv
b1WWAMWFH7cNG/sxlA0fZZzBMy/FXYz7MSYNtwPfq8qma1UBEn3t76HCXHc/+K5W
CFEBg9jg5so4Gyau5stpICKMGTarJ6voFAHm+JBjPXaYWCQ4mBaWQA7wOs5lyQee
wlekh513BJ5qvJ9aPHjWU0vUE+XRe2uxY5XPWdiKnuLkq0evdhdfoZYtAfIl0n/B
Tv0HKPaKfE1TILPKo/d6Jm19ODa4dpJ7KElV0L4UaIEShECoxgEL01Q09n0JXPfE
nAagRn/lZBgjSVT+GyDd2/Y4vjjZxHncM42GGG/W+QiSDhBTbMfGZej1AyadVRKy
33JU8zsyfO8/q/UKGXgw957QmD+ZcQH9qpoED/Uf5N4Hzzi5B8HPBDNVZ4cQRKrb
4R5mCi4hYCt2RTbLXgXQvDAF8Z+d5U8Z907yjEL1aOX1orBVYmeeAAZezjy4+svm
dc7/wJI/yw8YqyajVCD+/8aV+r4i+9wo7jy+MfqHD2cSRY1igHmSvO1FAxkbPGuv
ewN6FKClICNb7i9p7BJ7vgCLdnEDXzPOaIoXexx1HM/3Qum0Tsu2s+NdvZPdRZiW
hiVX0KJbeb6lmD8Etpw1xhRYVZtHpav7NuQP/yQyZhxjAExBe6v18v728DYZi2L0
SSBQAhC2ihDICdBvM3ILOPLcpp2RsO/2LBbWgAwadUoOZeDumPSfsQ6cmwcAFSAV
Tg5xLKm0Gu8b23zoxVWOe4bDYCCmJVjbmmRQ1r9u6ce8gefo77LN+DyYHw8Ye2BH
3awFu2sZJU3Z3sdQbGc/bSbRtCKtTK+U4I1GlHAj79Y7LQwNJia0tMM6ul3TAEst
JiJ7e1ja/3nYiU4gFnkXHbZwrvZDcq9DPbWH0I5ELnmFQzcBzOl6D9JiDa7H0SV9
CD89zKtLyd/i4GtmXV3qDXOmQrQcCrfPxfI74ShlgXH8Ijadua7T9xOMizuHIUg+
wukMG8cpxzj41+/banUFziulK6ye+CLns8jWtU6Wynq2d+06Q8FFxPC4GDX+rHlQ
VwRLuxOV0Wtth6zCq0LcKdVtmGDLixYMG6LE1B0mn71Obt6t1bFu8WAzfVFHcqYU
nfPwKkKwI9t5ukiZBINi3x1V7KySfBL4uxwQjbVqSJwmodGa3tX3Gvrw8joORjnU
1SdWGL+8gIMEkbKPtlWkDFeX6mvJ2AsSnfZqbXAbFpX5hmDcMiAVyfzvQMsnKNS1
aw9zKdShNBF0XtXinJGrHPDtAKbvuCOkedDYnJ/tAEQEPC+6/2GdelLW2mNEriVT
RUTRSntOTf5mvTQH1hfEwutdnyftubXD1F3aRdILKFzPNBzR2FynOgMzTm+oww/C
jnvNhpGFEJQgXX2PYpTsE2chjLuuTvpt/UgGL1LKNXj7DzX7oSZpsPqGBxxmrkkV
gwLtfK7hu6cbkxPcn6vWpZdNtD4CnXbn4zh8hf6KphiXCqiqHBImMkqZxNFO8IBG
+sRYm3XuPCtMvhRQRbERvzzRja6lxfyICodfN76oQrXf1kz8EGUxuHJhU3UfFDpH
LPzuKyAfJ7fIxHuMKIHLqu2eBwncnXXDfJwbUbsah1QwFWFm9MPwIqRWh7ZkuG1Y
QlmR2l6HbjN0WUFen9azOp//9j3II/l24EiD+qqVn6kPpuLm0czA5eaT6SpAwSjV
pzZsShrK1O96IcEunJnzw/CsZ4qCVMrt7IQlQDmh2LO2tmfyBfskB+JwBl7v0iKl
UJnRoU0vM0aRAouAkVzsLPaka6tNrpnyhVqcO3GL+TDOC+nnVkP3GYPC0iDpZ8Na
zF4sNBTEq2XTzj7G14zW3JUNN0eynko1lXAj3iOXNn65vCFDSeBlTZqn0E9blwea
jZOC1kX25sm8bjHjTl3Lo3itjC4RDidyziOrr6T2cDjFsqd5RcSrZv9AsEL00YbX
NtZstNZLuBHRqgbIqLWAip3roV6e76jeqEDxOT1WUT5M/zwL2lVA2lj4tvTS7p7N
Ie6YwTtRM7wwTbbybb70vnJe1zfoLuyAlGgQnT1r/rp9ys7xReozd85z1JTnWBpU
kmOPF3TYx5d4o9aL2Hi1gqfEudopTIy32B4pJZXkDkMZeLVPv8Jrlzl+HpLSLNW5
Cge15RrfEetAKgP6YRiIy5gOmMe2+QkaBG0ilYM8wFibxM30b4wKRbRSoxYz6CYD
miX+N/k4rlsAX6SzAIwNYOQ3he1ZrcKXcezLqUrqT0I/FMlMiDX7aW31aMnmPXji
EaDKsIot1FAHVyTrNw2iIeUxVBxjwX2ECpbmnSwELIOJ20aUA8G40uP7401JIllR
Ff+VZaSHNqCoTU50z/CmMNT3iG4xqAkgazUVbJtLtBlVQL1TRCEtUmiTXzHCu1H9
3AtozSLm+Nla2XbfsPbX/xwCmphE/RgfEPBmGGvYIPb1diMcBFtNehiXUxR2gTJy
n0li6LwcavvvJrTjYojKvUP8Q5DEnfE4GNIZP9gdHtZmzYXAo+5iyEua6kBcZkff
1C8yQmMAI3wfcMpP8cZ/DdCB6OcpVB63tMeJsuLr2c7aXMWuXihFlmd/LiJjpn1w
bmcfA/rNLEfjQjHU5mdeZLODqw0r4ORL9dTH7Pj0T6uZpViQIdmMmXXW4N8rwgJN
y3ScB7S2B12qeRLuFIAvvNAYqTTdgSgzzxT5gRlWHMvmBozjneElG7D/lZ5h3uQK
UTEkyAQtuQSV6Kj8ri9YinHi74v2H9zAKCDZR1IyCA2adrQl1oOOxxjzg5Z8//uJ
h278I7ZyYWme8t1s6IO6PjCUbC0kB/0wfhxK8Pr+OJsCjEw+TgHvF/X3Tgmgyg0H
kI/0vDcWNJFog0kGcnX8WiYOv5r4DTEuOZ9rB4zpYGERg4OmENSR6rDyGsL1ZcDp
TYUOIopCGlP7UAbvaAI4EssISyv3Oc8XIxcGWnWowl3D315V1LeW60pixn7+W20x
bHpPsbnGVC05IUJYvvggQIdOfmzMSniZcxNhczWySOdxJcbgPb+VQ802LKa4Vbs+
ome4bH9AD8cwJYkRc7V0kOb70w272EsI/Au7Y6WCKYwtmQC2/akjYTmergPQJ5f4
/8n56nQ/1xWBpLtPVqqGRUXh8FuaITJUIFysEr+PL0UR51zji1RS9ZmlJgUqoeSn
VbL+5wP1wk4MyI2SXND6SeBBKQADafPGDlMpI4XpOq68QOMP6AQrK6Y+Gm+NVb9t
RJ/Q0SF5rF86regv2mOOh3FBGyVJdji0pQsAuJUysbc+p8VSxUfgwY2u59hRzKz7
oJNrk9IzISMD/dFdllZKnSM45WoAqA0dk5KH45C+9r3upaP/DvfIFsDDW6p0et1x
Yg+U+EcaxCiSr3obr3Y8XrRjuVMgnAgxjYznMaxkww+3pSmW020IDUMnVL4UT11J
OCGVCyNiQABgBso1/qLFOyFij5KrjEoNiO2xShW2p0UuWxaVcRQ258LNzc95S7kr
NGnEapxeVhdwu3uuUSitQ1/2NH+EIXs6klHLbBoY/9OnBlPt9TrxLkLdyLJP40Xk
v4mMrm6tAeQ9U+XzY6VIyBkuotwtwTA28AE5uiV+q5YAx8/xklBpZAlHSHkshZfC
mPgTbUeQVvYrchZQoUpItdxT07wS57Fx5e3HVQ2zbLtr8ufiK9BTxaO+I210AvwI
qnczmgzSCNDt3Jo9l+X3dMqXindoCAqw7e0cxck7SAd0QcvOkr5dYsAI2qUo/f74
5ObUuLvpsyawNyblQyHMN4zxw0P01HZ4v0aP4HMaJvPCTx8zaE3hqHTWCsnT/6IC
J3d3gjPAJY8KE5gSQaF31gskOQBYvw9aRsyMm7nTyM/Rc8SAShBhoWk4YL8FpCpl
oWpI68d+AbqJEkHq7DMYFmi2vgs457I188tYSsqAaBMfnIYPjT5sx0NGSmC0I1vv
OASdWidUFhzmRFwqE1A5VL1gmVffnsNpqHT2VdwyikMGu+hc68k/iFqakR1nCk9m
hSqi7fS7FFW1sLXVpAgoIOMVGDoQ2TfsejfPG3KJoHtW8Y1vCjlk+XHTDClqKQSV
O0hWICRq+OFK/lBDIg2GD4uOH0KsWQWRelb5+5Ai1FrrQeZWfsc0pAPlhO7a5TB2
fB8SF9fqvXMpZJ9Mr+PUHk65/ARqcTAEAgcUdw4TQG9hBY2+ikPRDUUtu6yC2dwm
E3vWMgCqTYQFbnNOOj+ena+68APSicG6fCG3BV8lCzuml+cpQItKckdhyoT8+vW3
jFZO7VhDvSl0BwULgH6HCGhqNwvaGvzoq6K9oq0k6sJv7kQAiysKFt42F08o0KtJ
sYZilAh4guKMnPnp1gRD5ZHjO5qDlZt/EOkF0QU9JZvKOgnW/viP6gVcRVzEk+FB
vI/Mor9CqBbYdOfOZSLAm+komMUCtqCn+rRtUjv6vsc/1X45+AZznxuo9BTkwdlA
VkHb4NzRI7aGFopGxHMMw5Moq7ZN6Kl/AkK+kUj6BeC1nnoo+kdxGXkniGI2mVdp
u5SyVTBVPYh8hyL2eMzpE59gZAnYVOsfzB/RAdXsjDFMeFnoyk1eJiROnvbsWZWz
fmNlMr/SNuHlu6HS8nUeMoW2lQxMqcRg5ON8To/SyC7XNnjPTMr1nrzpd/vfN29x
p4dNg++/RAeN8k/DjFSuWubByVvL7cq18Lv9gUbT7ViihTMJUjS5CHgV7JSkuhFl
Nj+40I95X+wIEjtLoufnC5PEFkhH0ZpG66jV/Npd9jM9WwHJQjsi/cYEWYgOcWf3
g1S/IhVdMSUGi+Me+2e2knvJxE10gpM1WRE7UYfcOGj2NICZLhcMoATYF53uEk+a
jp9gHrZ6al6SRDv2IUyXBpYQ9/2gq2BeQbkse4mjofoCDCecBxAWur6ZJtgnJd6K
KsEPpQQP3MOpmWL0Iu+FlnePN8ZTvIqWqTYXUAvyMLoYnEOcvd4KzvwUU6BI1Ud5
k7zJCGpCteYqEpuqhAmKmjhqRN9b9FbnP5TfIKL/wiFWM/dEA0mYysX4OvRY3Evt
a3EQXJkNd00Po7+/xnqNvCSeJC8lsVc42AInWPKMUgmAZ54LcdyuO/z0c5xD+1Lz
NlITuOCyF3UDjoYH65p0y+CKWKBdb2EGRom74zBU//yTOpyKy94nq0YfJfWOGA4b
eI1rhVxaWzFgSnrrqdkaIaWT1A1du1NpPM2d0m44xHYkVYYFZqBQgdwwfipQlxgY
IT0Nr9MHoYeSTt66umCEb+j83MI0qPdAbCqttY2BxBKEdzU4uthkRL3K5R/CQrlX
mtuFR8ghQjO16TWkJnJvIFR+qVYTcWCPnascGyq5dxBu2NELyvkfOo28UOvv6ZWR
nXcA0akKb7GAqAJ1KgeWW0AkmG1xOlZ8NeSVnLpHTm6izZ/ovsSk5gu7kq2QQivN
sh1+xgDrTnOmn0Wsj6OUltW1wX8BjdTbB/TigDo+TIWWILKkyJHxJcTbtnrh2dWX
vBZ4U0YfVFkfjRM9yeML7wMHdLoHSYvjS9JLHRl7CzzNlvXm8XYE2gTenNTIBy9g
png4VZSWPoHgN80nxJHINrGlmqYgAvIIMkM8bAxc0xuUn7UqBCzWjdhYuF+UfmMa
yZKmPTArh4W2JFf1DzIrRvaXYlagij2bch00+zDgnQ5w9oCsf9U8n/NniMfemLym
ujygXomLFGT0PvKxeJyDB+hmuWKbJO3URk1HF7vEFUgPl/VhsYzidg7k0duZtOQF
nLZPssEQPXgPe3nwv2ZD52dWSDuNRU8bNPFCnBTkixncU7eaPzAcZTk7G8HscHB4
HuMjCEwTWXepxRMwct7lgoDaJP+2tA8IsAwFtCuGT0+mY385CX7IPPeM9o0s4v8W
94byGr+OgPQTaYCkAx5gWQxIRG/aWeIPaysK70MqCOuJcygsdoaDHTBL0BQzfiaq
O6iThRG5LZyWCojF3DUfEGAV6VWlEa9SIYCmC8LDKJwAvzH3eYitZ64lxwnqiZHE
7wiqLVRSoYbtrsv83kGT3Atznrle+5GbvCQI5f12E0ARZIcnl5MjImnp8VmJZ6JQ
JQ1GaelPHVhHdio39fIlzt0am7j40z32PBtdp+I1FzPyigudOCn3DT0XVRlyeXnr
HXEPkkTG2kZzYLbB4xn8W4uXt5A8zuWjQsf3/wQegKnyIWWVymbIU34eQfzCElJu
vGIKcqNv/pJ/5G4mE/tbS+KOESoabtD8a3g//kHDpGRNZCFK+AaUlDelw5Uq4l5G
lao4noc0Ufy1HKTQRxsPJbeHZQ9wPFKDY9vxl2Gz8v+oHsX8XPmgqC3pKC/g1Cc3
tD4os07Z1dd5s4cYYvJAP97ChB37ULm8RxN22+/y/KNYoNiNDMRpPUNghhlpVvIu
ZTuzuYbEcexP24TfkPJQm5TwEkS24BaUvvc0+xc7QNGB+y9CPyq+7QbJoGoxbbcL
+nlZ5Kwra0OtoAx+cMEtmKq2Se2xX1mvR0Q8xQB1BA/Hr6TuWgv9jJ5sYADHMiKf
mg0w77fPNGXXQ0JqmXJIQLD9U0lxi8nYU5fyt+0Cpzvt1hku6uG3+vZ+qQhirNOC
FAArSFUekXL23ymX6LztGOUc12QpgDnUaHrulm5hUjBVF7QOlsL3gkEi/zv7F2F7
Ls1WLTcavFoJ6XkTFzN4zlDFqxBpgAdGkXF2lLM6FT56esvNwoMmvR56IcfX0m6R
gfheRKQgJHrgfEbVMHI/WISexpMW/AW3FcE8IakguhJFTZpl/Vx0uVU95OOl8Ahu
fy6zxZkSWcJUU+vGQshhNc5JuRZwTwTkQoRXXzJSULVsmRl1t6l96PfEVaFFM7yK
W4rDCEY+9w6k/50bMQcKYcba9igOujIWoDBqYu9MipryMM9eS5pUtn8aWOorqcdQ
FxL/NPdoiSmufNh02I0ioynl/squz0jwNxBcgehCbek4OgsKPVYBFH5UY1ps1mY/
Ax/wrjSz7SpF7jdnKy0HnbWx/aKq8kSWssgOu6yq3d7gC9qfbYSsnP9Wl+pamx3W
QaSYQZ/fSbmiqVpO45MhfciC8s8gcHf/eq3FfwN7+EGnMw2iCGZWqJDKjcHCWmGq
mZnF5/t1kFUSn75s20mE2gF1nZ3pgaXmpZnnzn/FipnIqElaFpmsZ5qtaUwMZgP7
8aFePf+7C49JJoRVMkDhdJnl/psTyLN0jym5dQ0Q7MGGZH+8ZduXPh06ij8BUe+d
L3i1MK/s4Q6/biqWifmZHQnS9uehhpWZHlm5aVON3OrpgfvKar81e1ZoBnqIgB36
0tx18iKmn3xrkbahtLjWlF6XD9rfd0mAdjdZvLPG9zD7mXXpXISV99IqeD69elB1
PAiJ0yPEnvwUQOUrcRrYSmFfCYOHsH1TG6Knp7v/MsSnbAmDLL6inwsPMUSrlXuy
Ey7cV21nMACyYklQGyWAxeSTgaVGLB+/i9XyKjZMDFMDmOpDewLhhKJRyHeF6lKk
jjgwyuzTkfWApB65pMbijO/KtxCl9FiG70gZ82KrG9cppD2w3M/NKSzivJUCNWxQ
eLt5lo06qdwcS/3nVEgRtquCbUqiN6OBic5LkkM0XzMLSlFu/Ga2/Al16RJryLcI
wwRs+qmtG3OMagPpUvdfJxJ2F/9ZG7rvtkMrsPqiZMLVxlpIl6gCsZcayrq5Ewvg
UDKTnUSGT8XqXJHeI7mO0Gfn0kkt64X+gzVUip2Ywvpuwj2XertWlyUbU37VtSI+
Mu+9V8ar3ZbuRQ5KNqNEa6IgTulpdDRVUXHKmhdhmb75TvNfyCPRSsnrJ9b/Qz9d
evrv2ks4WridHCYkpy5m/fuDkffOHX2SQ9Z0hROGpXdmR+srp/Y81L8tyLwKVpND
PIPdFvU89wM5y7u+Y/lu1cowf2jAnTu/OfMIjagHcWj8R9sf+iP8r0SZGmyrGxnO
xUEFFq0OYlEb0138UCiOtSBQ3DEJZw9Rvqerhd7BIjhPfmG3fSNp3xjcqFSJh3PM
dWWKAgaIJb+E+GB/gY9wqDi906pALo0zpyBKje7wMWM2pZghiXxfsbb4Z60id2S1
g5/yO/5kYiXQi+bFZxlsnD4ynaoaLMct4JyhqS/PmpOuEzwgA1QfU4ETU/xAzqlT
MddHqfX3b560mQYfTgUsGLpKD+YDEY+FPerfkOaOHLx5xVhGov7bE5aBoxzmZWwq
Jzm06HflfpNFBVCZuYjpu+8ZcDG1uW8tuI4mMBcKX1UC0MtGExw8OYApeg0P4GGP
4zZ9G1sQTIvhjeWxeZhnXdp3EGx+geZaTHLZGgj69aQ3PPaolfAAL/jERnDl0yDT
0o6Pik+uz545cSfOWhdoO0teRAK+NaFH+GDh6nHvVuz6zQAlvze0GZ/W0kjrQi5Q
vbGI5kbJf2GPzYZzUoIFxfSI+AIJ0vl9Vl7aptlY3txET9hu1AiJZfpjqF6MiFIc
u1w3mtHIo5ZM8O6V0K1TOR41KlT9TNixl3/FvunCY1z7JFi6yOOgXgJzKTPI3cCP
/vm2II+E0JWEA3Dv2h/kw3BFibVC/oeW7iAhYdxu9Hp1Q47HQAGN54Cy1VTHdwil
CXNhyA3d7JBcmzRiVXjI0lMFwwg5MY6MYlROxaGqZfK1wVa2pT4v83qfATfNE406
BiNsRe/u+0YjJgP40oqR2oq1+zcQVsV20Wd8HnmMkY/B0a4JNn+DycKrvyKCFWs9
VQdoMNx4piDMM5tOCxGdfvAGkRlQjlGXkLLCHTJxS5A/FfgYfpP9JFPeGm9zPQDI
dPQ01YMRqy2uz9NvSZefAWn6RNvE8iukPou8ZYXYzqudajb3Iq5sTd+YohDmn8jS
cDmZIYzd5b+VKIwGpi7Nt/YRs5F2FzZYDEErn5i/BYJ7KXzDZNMXKU+0P6ltMVZe
TVZ6AMqflAym8ws4yjgPPhzQOZJR0njiHTyGvGOMRNdX8KJ1KYv6iWum9ETeTZEg
ZMdY7R+hvvxJttsPTPb7vaGbE5fqNsSRotf9tkR4CmTkflILvz7rhTzPtDkZZEqJ
iU1Le1qtw9SoLyOL6r0V4iwPP3GWE9EmhHbXIhFS6zjvkbj6xU9V9Npo3E5YZqqL
hq7lIgOm9gtTXA7L5UuDNXdh6HIu84THz1blAu7dDIPu/hCySxMerDc4t/qzsLWf
KW4mzHh7xTtKVARkGm00JxeeAQkvzv0Q5tIrGoiekjIcKFpgh8wXqkipNcPgl0Zp
o7RakdmFXQHNgitHq0z5seB5ArgFAQQOiytxbu5U8e5PFUYZPJaffLdHZs0ceIZ2
xg8bh+2skqby/wIq6+6oDl39oBUZ2I2Mlj79KhxQFd2mhjA4GP9AfyN3WPtznImR
hDnwYlhZ04SDqTGEZYoiwlRJcei6H1a37CbWjZYXNc0e+v/3iMa7w+3PAiZ3R6n0
ajXiiVtYB4NE0EAlfM96DKgoE0H6qNRU7a6l7cGtalWbMFtJX9LqID2B4LSw46lb
qgkGuvfMUrVnpyLox3VATzvzOS8AK0jZaoC+5VggV6d4yRYbUxy4Ik2Qr6hpmP9h
iCIBSABi0QUuYdBFAGH4sCLsam/yzC9XWZuQHfrl3dCACuZeEBvGH7JxoUPRicHC
BlaJNcHzAku8NTdw98aYXugtn5PdLGgcaOBorYCN5o+kC0W4bYBrbAOoEyQ08lsx
6ofu449Jnz2RcV1oXchS8mE9dbDEiJ8W5lFADs4iNL5uiCiu184ZC38n4Qk+A0dY
WkFaGeXSYro9tNJLOf47k5ehVxF3HL0AywoSbbW1jYNpcwKjWQG/tpa/qAlpGelQ
Tg5FI/cMXAZUW7qZgvu5EaaLrYAylB7pqn/ZnNzo4iYCiRyzQXdbOjPKMQenCQOo
wmvwssckbne9ol2nmFxEYnRkFpCQ33WUE6kcfGTcBb63DsQzSeIquXwuAbfBNaeq
hjCHZ4dKgCXKLvHoaLiy0GVH1cyj24s80Jb+27YoA3L7X0N5skn2BYoIgSCLO3tn
20mpNFt/VmoC1tpPN4CxFhg3Dd6ZEsZRf5lO9VaERU8Csb74sQIYE4S7gD9vZDPX
22ziuO76va4P6l1IG9L8laF+Pqua0GRaYsbRIJ/Zr+oWyxGeAHDjN/qrxosEBAHI
XAMqaKgGdTqKv0PVaUJNL5NMu9+4peHM9rJFNkvqg8WPxzxV8o6upxl/a0fwMqLW
tooMYxcLjDWAx1692jHPXLe0aXP0ZNSO8WPsaXycepX7NK5/olu+6Mpoa5xyQAiN
BDmtMXCyZPZDtgBrxui45N9aHJx1CygCo14QhBIiaGysuJ8yOk5er8Azb9roHGhV
XvNTg+2FXU3drZRz7N6O0nMFtnIMFUFkZmps3h+Tk6e4bpKtojcmn7vb/mjpxye5
DxzQ2DV0b4LS4lmdqZt8bHuWLHF/P8WkB77JfWDejCbQgdIe3iZt12XAK0q1QlJV
ED4vZ8qOmax3sBee3z7FEHqh7e7JWgzBq0F/rD+2yPcMXAus1JuTUUkSHCYDU035
EkPgX3CnP3CE1yzWMQJGFqKGASLbQpO6yCnUUkOAh83H31XR1a0+yKru0bm6wq8k
N/gTYQgkXFH/gDee6E/BU8YojyVotIssHRuqAE4q2hHwXKmcLQPpPsA7KO1EyE7a
BVXXk/CG0AOjLiZA5Ehk+cff2av0Drp08hLyhSx9P1jLOVTpbpYaah2+7QRlC45a
Bwp0Ov0iMmSRI7p+w3tRu6ABhjvm/RJxReRuUAjdSrnow5wDWVxw3Lbi3dCrD5X9
aEu5s38wfx0gj2Y8zaqiokoT0d0Y76fhi3X1gKGK57Dzdnk3mI5rk2HXbOxrjE4L
WkgrgxaYD6E57JtfFajHgLmK6t0HGmJDnIsq1j4h9Gd8OV4XcwsXDGF7aoC9UdnU
n4zssr2K6zR0jgyGAppvE8QoSV1qsaw+4pSAYGhqKD8OHEbM3JMsbfspYGOCQiF4
0oxTwaFnxEuoH8NG2oNOCW6V8PUzyFLGtJPmx2kB9OopvhdbJcF0KYUWzX5OaulB
nDhA7gD/cRwIiA9dRZ11aletenoH9eylBy3zn+gU7flIP2sd5GTfXauXxqzd4xrA
exVhMQqHVccpsVS2hFVCyTW+FTPq07BIKFYPBB1ix3x+N6h2yuPouThtKdYkCLDu
T35P/SapG3i+I36TMk43yaTW/pn1WP55i2j87Ue0PtZHbjOcZY5tF4/P3Z1hjSaE
SNwvmJkmyX4kTnoK0zcV/E9UZ+hFW/zaxPs9drOFu9lf/G3aXszet4iAy3am0g0D
eeHYaSSy3SqS0W2Dd0OqDK/7xuKaDddFMh+OPEO28tE6T1OMdewUHcbMa0r95V5V
MY8n/D1fJ6r+T2DlRpHHkOOdnxcCzXSyVBC1oRhfJjal78jXfSgtOTsJMncxE1tY
8lAAI48+UFPrf10+EhClCmVv671lU+T4AOe5E4OGpdGcEuQ9HdCEF+5Wfy7GFuEw
TKXPOoiFAWdbJq0wVMLdPKgaTuLez0Q4r2e4tkIp93U1Wh2NQyTfuelMq/b9Nal2
3e81/2QbPZ4NVENHELRbPT0AJbYQiA0rO06pMeY1BwNTIarnP7KyRB7gMmxcXLOs
rOSgm7tSuS9X53ard2hA2Ww3TiavgR+v0CmDqOzZy39qUquH9dixOI7xSLWD+zdP
mUvfoBFN97zpxILmA7OKorllnxEosHLC2vz7HBANFuZWokmwrrwuj2pQDFlYwt5n
pO0uwMrUL284aTJnMCwADa0tx1r8hZGa97Y7GGEcYUhPPPUka5i5MjsLoZVa02a7
R+SM+84AEqLPtRGCuhKmNY0XL1aE1QJ7csd4msqDamtg8Cm1+GWWV7pb3sPpCdyx
6ixCcxbH617rMjFr9Qc29r5oPGruWFFz9VmWDNFazrNVdz4kZKBJqNkgZASD1E1F
lNzYLAQb5CdQEFCQLaw2pBGahK2XEFm6izGccqvD8nyjBgsrNCEOPBaJfOihVHIV
SqGA/0C6r8Wbx874rjMeyrdQs0IJzFJ9s7fnSIT4tLwpe/LCvUe9b5vy6JROsgm3
R/ZfSxGX76ItUs7UKA0WzjdDQhwremHxY/2mcghp0XtoH9Q5Vwy8ksEH7IOMHt31
R8wgbwBjFXuT7GmNt7vSWSMWRQMKM3vq4l+muNf72jgq2ScAEs3WMw9EHDIzjY8P
zsKLuHxLj2hIMB4cdLNIzu6c3bTXOdccGZUmQh38okTvutzWSC/aq6/peH5hYDVs
tjuOnxC+vPGd+FPax16qNTJJXWNENrDotnoGcGvNxcO+Jsf1qEqfBFUHZD9OqNyc
SiKOiore/HmI+803sBsEJfxklfmfmS3fzmVDKUG9IipBpPiChiBOI5FVp4H38mEH
Zib88y+DHVGn59J4is2bhjyqEGY/6ANYcmXAOt9tmjhKyg+kIVc/nchn7vWYL022
hmC1bhk7S9jVCNlbQWqv/rO44AwYhHunqcVy0qAHmz3CIrLusZ/hXWCuc65oRw/v
w33j/BdJdyKhX6OKIfJBHq7LOcC2wlvLoMywwxe8ktZwqFMlf8MEvFICn5cScyaO
mkckfuI7TfeClaJpNv5EwvnXD+05AreIrI9f6dq4ws23y0mgbtjo5IJPGPVmGZEl
5f1rnKu++Utu9tJd8eyWUZ/ewRrT3WQQais4mwcQPm9ftjGt3PI29Q+yeWTwRois
i1KBcm59MmqJM+6DImgVAjYSo976U++d18HyTdOFq3sch29uYFJkv8vJwx3WQr1y
knjpFQjwz02csQXSOmbsKruoJ4FRg3h9ZNXTkH1FAgFiXKEtXmxTdhb3fc1UrIAA
lqfN5RxCS6vv7I6rJe6uc7FPfu6s/LWtVszZG0MQICuMS7YWP0lAzxWvK6D/bzTf
IBRLfHmsOiqIkybYFxk5SxpZ4dDujOZE9R6CG+pbVQia0l2s3lVZ5SywuRsCLQhO
sPnr89K3UtJfIxmjECt/TOcnZXbpEAHJnSenI+PrgyQeyAZ8iPHO7hTMvmyQcuJv
6zjsiaJIDlmN4BeUB0+prok7ntAjjyFc/fprrAfCo6a+THKrJLFCZeEWTWDfv8Hq
iS/YNLB4MEgpDHvlZIW0CcA2gOvsvDop958h+tGls7sWy/YoH1knr45nn+dUrB1k
dtVioT4OD6qQFPwH2V3MVVJjpLS7NpRCH9HLZYv+abWgUP/bGL86Q9HPUBt2ZGIe
RBdcE8JW7xu8BSrSBDK2/VNj1URSEKisOIcoFJSG9M1Wt6j+h+ACTF91N4NCTDks
4h75H/xfqCpCTRVlzO9btgM5dVzmHyCvO7UJu5Cz4+mTLRMX/2kIudVxGj4VLEr3
vmbbTCPv1w5sf3PDV+Ft2Ci2Hy4l9C1o+Y8m8Yvzt6hinwh+UCxXae6qQBkjJsgp
3m/V87tn+TTRk3/lQBPqfrIdw00+zvptkeC7L7WanyMJ5AGxqoFX2BheeOec7l2f
SPdST1QfOlCMdKYfIvuydSgYTsktg/omo+Ny7bhj/RZaarrGvjrUV+xGgOYdZxIQ
AeDD3XXBV/EbCYmxqZj6BttEGV51y6lJt+a+UUPYp4gD6yDZ1pSq9BBo7mF77Eow
nRTNp0knE3HA1Rsc1atfTZcSuNWUM905r56XRtW1O6Ze3qA8N6PGYW2DPKOQR1rM
55OMv+vCtO3AAFu8aaVYKB/85HM1m4fifFw9vD08z99wfe6dg5iFonkB72MgyBXU
Cge+Yrnz5mGECzuwZMIjQqG5FJaKVwYpKaSmGT5r9gHWPNkuC0ZwVKy+6yQmjfWj
Etd9nUC2xgWSMJ1rTmHbyEfNAn2V7kzg7mu20szWcOzBqg/aikbm9xviW/9U9ouZ
XLj1nMzZ0vbGCQnI0Iht1sy6wDinfczFN06YxQ4zw9lzuO4f795wrC5r1mYoMTqQ
bFbHOnxi/io7MvfnIs8LBCpzcBo2+SI17yfFkhglXKueL+g0brNjMB4Nud5t04io
3oqGgoy1HTHGvjAz9DdjKGbQfCjR6xi46dW9WXMf+KUiifc3sFkfaogbqgmZHUO/
Weypam8Qr4tvxwi9dC9gDUIUIaVQO14bHZNM0KAn/mZNFHV4Y3CJznzBQDq9X7gw
JwmYgvB/Bzp9y/VZDSoe4E5QvsVIVTtWz8JA1O9CaF5ohtyo+JiIWafEALhuxmsO
DOItCFWtCNhN5q2qkfe2PcXyiZlfCUI/4RwgJ1gwdfg0VoRvdhPQSmW3iMt7/VsA
VOZ6pc3rI3e1sEOarPPOup5eJ1FmcK+KtAe1LfBUzXpz0LTUozCfs/nfklx6PSGm
bv49743HNnP6YpF7Y3P/bUISXnOzt7XqHsTlya03usx+WATbg47VEIg3s1poJTbr
rcC05bS7Z7LvL+iS2skfMVzcxqKc1iPdkG/gwozISoaW0VlFo8KdWyGxUpQ1merQ
D3SqdkbocSQdHSuTRrhx8G3WN22hogu4KJBleym7Q6Yzn4sHhlS688P9V4gySzNf
kPRo/a/e4vnSwHTqkGBySOXMOmQV05fJ0nJ1XF95a0QVzIf6DS08NhYe23cJj7tK
5WvSZJ9e6RVcgDFM5y7psYUnWZ2fl+QGTno8ZA6Z4l7R+Z57DqXwjaWnHO6o84I9
yepefuAdZzTdBsj9ajp3wwPN2H872/vd2gukmQGY/fsUoBB7N1fjT4KkP3QhLtl8
y2hobB/TEEOXL65EYNoV4JnD1BP3RAJWNItrtxPNQpTSCxFbgwssW2ETXpEMfUVG
GcqTu7okBJ7JI6KLvTuv3WvQq1ZgZwJ9zKOs77RDEvgV3P0QNJlQelbFix7CDXlI
Um1MnsB/MxgRexV0DRL4z0UCLKmnl1+6Ny78qmj+PXwUHHCyJtjIHODIBjs/28DC
RfUkAWJn6rcFS9YgMIXgGMfcMZtiWROw1ZayFKpKBeHz6s6FlvAeTH2X58biwWT1
PsEHQ0RREBPO8QHiZU3GThCHWTZwexONSgnSOu7+pYqdCW8GoJei7p5pNYTSGUVr
ABFOJRY0+0/gGyVvvDm3cGStYv37JmwwX5DmYLXwtlj0HmILJy7abiH2SdquFN/c
mYiXBmop7YUhfSYBgwNxM8szRDF5SAV6qtXWY+DB8RcRu2Rxb/y/VbJ0uG+cLfFe
LHBEy7ApTMnutqtbC+5kzlGJMeuFFhR1VoJyWrGSdDvnPi1xBLWROB99Od0j8nJK
8CQay6OaD5lkud2n6qGn9h0eHvnA/YcqeVvjmb8L28MdyN4P0XhGtKlGummiPsBf
GDcpOWsRLRizRqqwpDzZLVg8fhpwXoaZnzraEtXNs/THXiZhC5J9+X8QAAyClj+J
A4gWpWrK0CncGiHWiP+vnPM8rsd7GqFYgBpMf2WDiI5ysm/6WYH7wc9AIY8bBrVg
p6A0ckJiRKufq7/5r0+7KahV9AUAuLCwtARs4uKGd9/rZKHjlIg7T1O9LgJGVCTi
MQxzPXNAR4P2tVYNIIMWQHGdI/blQxihSywQRAxgyvHQ87lruq14k08d4pcF8tQl
9rlo5bTCES1yPtRWOniYOAI3SJWPHRSQHQaYevkDxdInQhsecgeBCIevGgjzV27C
WpfizvR66wD3gfGuXTNrRigOI5B876odgE6pTG+8ysphHRiX58Scku89t4fiRofb
j0c5CMe9TPBPWlSHsipST+cFgWco5fQOGBMCp+NncY6/JNCBUB/7GzuX49ZOlPKw
2n3HXxUQm/0aIqZHjOIYDDKonyoOCfkr93mHPOqoFw1ArIH6vFzMfpPxtbb4s0Ny
OpgCGVYJABII7pJwmtvu1KlgJFfyBfs+BHFD6CoCBpbv6Pe5wuE6vN++PomzL2Pj
tIM1llwdQ02xdJFS0J90wPb1U3aX72es4SyD3stpUh63ISViUa6vMP2tn/M2L5Qa
+dfrIkL9UcaH6zD8w2IFaDFznH43RBQRuHCqMN7pu5Z3DTTqzxcFiMd8suCvubVr
Oj5rI6ZZ0mA7050Ioiv1XV50q9+NGWK/8WI7ryPYr94qyWLDWjzzYyLo0o18qSlM
bhjxKB1Mb2iLArlFwLWKSWlQnQXYgp5zcrheQfJ7n83auPMY6whlFA4X24ZOAu0X
ZL8X9KFqkdfpFKbfkt7aiXKfzNsNyxmyia2krshrg0W+XbwXlTZ5PzwLEfSs8Jxp
DvmnR54sueGcKrz7hx5Wk4UOHHTSbbh/uKN+V95+KdOAIb/r8PK8vbqwfCJQoFZB
Ux/+M6x12+9NzNKxY0bIIufaNKwPfrAlAoUvsDfGb+3EEhqmbanc9z+TqfyhZJ5T
lK/IMXDUsFUW/WLXVD9V8PFhYQ4Em6WclSd3S01ryLSnogNqVo0NIcEmPAm4rcRr
elS2ktLql/gkrkOjZsvVZLvXd9Tcv7aib66bm0voD6MPEC0NzDYxu0f8f44MJPRg
vcBrhhHoFYxPsmdl4tt0EsFjFBhZ8Lc3bxwweyJXyBwMrVj9lxzuuj7sA219AFmq
7PZyICQcNVqchj7ZE1Iaf4Zx3wpJ2A/XLfektUAqwzs7YSzmSdhxpPt9YQW4AoO6
rk76yW7WuCsg322Imlh/Er+6unTp7YpovxUcVNu+tXm+JoHFAjlpbNBJ8JT8nmtP
moLHXMQM23qYgrMBu1H4hat1X2ZPMpdB+DFyweTPHAQgTVhMf823aWA2fKlTi7rX
51N6zthQ0eb6Rk0q6Ceix5O5cbgL+PK70Vu0clWxdoYeTiprRdIuBK64HQh9DdYd
kHHjwJz6DqteMa2cKmDTBTKPc1MPbKrpu5I+XtKdy5CXATWRFVKDWqbNAJya30H3
OUFz8W9dFRiDzqEBSREQJM18TIKLIOz949aNsXZGOHRIJkOnvT6nrtNeBDYZfoXX
Cv22XPzmwRGfifZxHqTgkez/3a0R6IVbOyYDtrXyAsK7jYSySYOtuExN/MAae8eN
ehbj9Wk6X/GHorFSr6D64GzgyLyXFYQbgTP/gcGFXbRDmU2uYI/ah0OJYs7d6CfM
pm/SWhm8paMEdbxWMdwByPG5FMrp4C9ABVpavgMomMugqurYi8dtVfxbahC7qm29
O3WV4LP0h1VwtnwcmEzTaoeI89rBDB353eNDZ18HFy/VE0DvYDrX08JzVbjOgczn
8X0x3bZx8/SPh2J70BiOV8tVTCRJzeZe9VdzK4x2kAFNp7O3J+SD90J3cjg3Cg8I
3BeAntGaJJ1CCXuEwRIogGhMQ8X2HQUOMCcaoM4CNH5+4PfZGhf0yS5cAU3obNzn
nVbVCCTttJI7lviYDtF9cBkv8k0BpntjPHISf0XawEERXFAUmbekPMsDUBxv7cRn
SPHFSAF4CER+vHSGs1wGNCUOxK4WFT5Fv0aOuIt+w6pyWnwjvKLBjrQjj0wcekuP
rS6jcSC6OX2+zVKHcjxz6mKmbcjJ58QssPYSG4xeCMj3A7172kwwMqdVbnOmUCNN
4iUKKf1KFWRNa+ODtbjLf88rX6h/rPt12JllglyVRRIQxVQBhn7tK0duCaL3g4xz
BTwZ5qFCjU2s8aXNjtmzSK/v2MeJx0Vfqr6N487ihu1/v/epf5GcHzmm6fmo60Br
hVwniVKSl8F4Bm8ArlGev++updIzzJSZvoTdCP7lUCOAHWEBk2V8O0aP7n/Rh3q0
UtxYOybyXCyodNhVeEuo9r+9QYwNUsu0ke4H6WQhzbEhAYQRBr1+Xv1EjlhMkK1T
xEmtGZnsUkz5SQ7DW0U25gYysBNZWY9PSVSDV+J7ydcs9h1NucViRIdZottNnJBv
fDi52N3sBFTh6nmCSvfqN3mLsOe3lT41I4r0QJtHTfsKToo+mQMP2tfHPM5Dy1pz
cOpPVwy6MvH+yuZLMKdEhmlC6R+kqFZjOlD6MR0rs2wI2cUM6ruS+6ISf9FZzzK0
wEni2R2M3ZZ8QTd7f/BsACZcD7idqJbnfyDv5+EXEfeotS/dWL08keDOkwFHTzvG
hmB+sFZdUYjxuB7uJ8ItQLwQGGGHYJ1EWpCzSlkjdHMlglLcEwUidOYW0ehmzggB
FjvP62gSgCmrDHONjtdrAg1HGi2MnTKhs3lTxReV35b5fhJz6Iq2h9zds8LAaTdq
PAqL3KwHuDMbK9X9K0bjELM5C65aOVo3PPGo+ox5OqanbHD0tIXgYVuR0M0TVg1m
9v6Z6QQUDOxFKpQTwyc4OpMY7x9rilWNBTYeMsA6pr7qIu1FIK7g5jxOeDvZEYRr
Ql1vzHda1Y9ZfjEZIdAPvNlQDequBRwiLyVlkxHNx4WlNUggw97W4W3JVKAybuAB
u0IRb3fhGBE12rSnNTkEUt5d3C3RDSo6RWUz0HjC+3wqltOsjA8hWTtI9bv+1UzG
crMQiy6UJo1IZSiEdHe3UcJpTtiqVe5faWzstB9U43FzgAeZqDXKGSBFXOoWKB4O
nCnh0oH3qnfva8n+rRMw0yNYDdpsm7WZeHyY0337IJ2CPtSjpkZmA1IQHkq7Eu2+
ubIhM1U8JTLaU3CFKktMim+wtcRewASXOV4M2y5TkoLzkl1k4GQSa0g92ImfkGdY
q2rW3PYRyqhdvChw15VZEnh6nA4HeBXhORAlLmY4C0FdGzf2HQ+bzHblPwztK4bE
+/ElwWc9h7yRvzN+OpzK3YvyzwIYa0Z65K6u/IwZEXXyuiYGLdQ1eYFw+W5UoAPu
vxvA2bEE0YuqJAOceDDHKCaHFkpplg2BxWz7fkiWzmWnE3IjoW1PcA8LIJ+wQ1bW
qOa1ev6RTgvA1vobBlhvK+1dgTMqDhaB+ilVzyMYJe2X0O99TFaSkhQCr/uc28l8
I9Ui8d4FA7Pyb9OPsidgohcnYm8i3iBmgG2d9H76Qizg4iU5CzkpwgZWuqFyFziS
Jc8So8DQgQmsXvBLAgya2HwWOXwpLGYmBcP+xyPPfTqMj/3ElHkleMzlJBWpafKZ
oqCg4JMsmdBOaLfeSycbBE0pkn5PqGzBv70oVsf9UxoK40BecRwGPaGEkwO7SCuH
9vaApKgXnps2FWQxqv6IC9bJ4UtsOqnYuxU+0meDuWNbOdStgOI21grpBhCUAIdP
FLIt2NU5Fvw6nA/yHwQTFvbjK3+e4U6P5L/YmZ4nOsNXK8bHfYflqVbmL2gHQJ0C
jz0FGTq+WO8hlNin3MQH9476tDxcYw9p2Lszsk60QC/aKwv78hZQP/8QpwcbR3XF
X7vo7TkSWPbSOepOwccJG2iHKiXrvyDb2IbbocJ5Y5IS//lqrss7EyR+v165q81R
R2cqa78+rSvJHnsrURpFsi58gXEs9Pr/7EaRF1cyjDOF1qWAwYpejYJwOmhcxrOL
ROl7c+wWIrVwbj7DWpQ6+YAIgaCCmyAJqtrBPSY3R4speOnZSJnpuQZo6M9ub1aA
1+FofGXDRhElEXYDDr+Si8Hl52iSNfAWiAOr6YQ/lHIrz7zkiPiR1VGoh5u2TtWd
4II+e4GTA5cPaeww8v63WcVXx93TJdIPQ/s+z7dDMSMYllmjneaW+BBmlE4SqTXS
shXCQbEfthnZzdsOxrVeatWT5egEBwYIZSbpQpgRRgBtlJdf4esxSuAq7eFUEHjR
i5nxv3+b6HdVXLVPF4yMCBClGhbCl0sU/bs7LjdLEgn0R5Ai5dlSKffK7Qsr1d+U
i/IwfnQDEVPR99x0kGyOeM0KxZC/XIPPBUBeX2frThS0SxUF78vO77Yf6wvdlbM6
L6KMmWP/QWF8GAa/f/xggXwQKl/oa1xEXc9GX2FkjnnBNGaJP3saQpgVmvruaMCi
OoEN/HrYWRt8MZ2Bxag492vSPhFaHyREHM/sTMiLAkbb0qCB6HoBCsGeFPiSXtA5
3aOZjCpv2bHr9LTv7aCPF2MAnXp/+GJOEzaeuYU5OiBIQrWfQBZd5h3UybiwO5Ia
sprsw9RtZFzlf0B6STsh7mk+XW/aZaxMQsJ2hCQSzx2CgtWtBFRFN1n0usLCfFZ5
9S0v11WRWOk9S9lwhlIysmHoM6a9/x7of+Px/dTLX76TGZ7D/0qU5EFvOWOt0LWP
dKBehyU7plVyd20FJPpa7PuhokK3akQUetBqy5+xTbmD8FlCqNAWwHMsd+1a9l2M
uWX/u3GmLPP3NJPpyTQG+lqHAURv+8KkZLQ/OeGMovNmSCgzHXgSP9bFN2X9rGtz
BXfWqJUSuFRXa0rnR9hnLvh2DYLE5Etw5fH0FfMVJz6OaXfvT7tit9lGPG4CeZNg
GoANcydBfUxEslPkbQ6+hH0dOHuYJI76rlZzFdDU8QZFOtwcoOw92iT/z20APE+8
ft3UbM/l/jOIpRyHzj1LyLRkyHgfncXtBRCwFy7kDpKWKSB0+azyWliZPu9Bph/O
gpfm4QCkyrWlfKmvHBTvEVdbEmRVZIRybNIr8rpcM42z9D0QiBip4+FIgeAZzT0S
FBSABikCTNH9olyjrAph7snMtaibwrJh9DqiqsR49kCrxywITdPRJrNg5BCgN0hI
z76FG5Qcb809RMbTncC0VXU3hpz98docFXljlwBCfKlQV8LoNcCke9eQYR9buRH5
8vt+pQMN39g1Xl4tVMYBokSeLZeTknoM8F1dOY/IcPkDtYxrru2wM5Th3lLRJvkV
umBQTLW9SPQ3EQOqNdU32Jo3CHscakyv+8nuZplbMZTBrA471coHlV48EoJmurCF
wNmW4RX7PfjxKklBhTZr3VoM/7iATckwGI6DJO+oBkz1KLk0r9te89Q/dANk7YWt
el9hLLA5vev5zji/SASj7dECXAbvdd1NZY2ch+CTuT88xmQBL1rqdkqzHSgkiYOR
s25dORidfibzE54cDnv0ofUf+FQLr2YEsGMKMOv1t6gW/TQtZp8eX7wVWaQI/kLj
GyD6kOo17pX/Do/UIRfEiPCt35JmIDUhg2bCrcJtPKZEnf1tprh4rUjUruDH0NW2
/inkQj4Y8g978gADhq4TDu9KatIfp3lQgS6edo1jwUSrlc/IIkNbXoUfgVvBOrL0
S3ZT3oGiJjDUrznQ9eVE7zLhpmRYSUe4KnyoGINe8lAa59AzDvVHR9Um3wwI2qEC
c2cp66XyRLnt4OEOGHe7NfRVvzD3XLCC/yHATv4LOna1K/JTh80j5GYjMom5BKRa
FUykHarmNzsCgRaMKi3UZdf1R5xaLAZYlAs9uKEyN/H56jqF8esStRFyoE2kZhXx
q4v+FI3h220xqtfEPT0WzHOxQubqtl2Ovpdjb5DBcUJetumxXGZg9pXWehv6rbfx
ZkPkiEwYhybjAX20fbXQO9GEywSudIa9Ck33Vi8QVil0fumROcmKMDjHZx52hOix
i06Z0h4s1xpYaQjzdjRSwbsx2qVBoVAY6LtBBNPcqWgRTo3lpJHU7awWh0O6Zng4
K0jqiowL95ibbg1ObWkf8AV3qzkyD988vrGJkCmeLHgPv5hFs1A8NFJMEU2/qR/n
y7RLZCbO8t/RWGpJm146tvVohyXK07AK4UN6M7qXk61F0ik/Iij996vTndTrPNbU
/0RphflCRkN6vvmPejuSXRCkkn0wyDPhc4rAo+FsCwbKyLtU/GfBvrif64q4Zmks
MZ13hqCOu3Ct2FKXS8fu4JxQTk+rXH0PPXj5Dbh44p/pgr+bFkisp8AeF87Me2LL
9GjwOiruaOB9lGKGBNCY1K/b90o6tp/+Yq4i4hxGIIgzMze29/0rBmU6M3A6GAWK
WSXuYD59vSzipT0RgjJNo7n9K76kobDnE/83sC3zuYRVh7vg5seYtGFk9/IaRHWl
IYP6mglOsLnansJPx1oV068klxyYM98Rdg0tgX0TUjwzaRIoAbCz0sFINNpp9Sg/
v9T0uAF41UqCBEFiYASak5NNx3q9k8WrMjGx5wgbTZOer2iaQYl+nwnxcjHmBbGU
tTHIKon5JB08YWuP3vjsOzrqqTaWDBp4YtAFZuvd0iKR4vJa6u46UqoOszlTSzcy
abPQZ/UNwOvUkTrE6E9Fcf/CpbXVfT5sJSJ7yK88Fyv1spVUHx1q3P1tqrTyHDK7
WzYDlwuWN9Fnl2h6sAuBq1lQJ6HcMg/EhPyFLAR+9aO3McthSTXuJhaqYtc/oiZ1
1UHaTRTqgJiYv58BQzjgOvlOlXBI7iJQqG9GLiV5wjbzWzjuyLE2XLoztKChq9id
kcEFXcli891PskVx6lKcQDeyZ+bZZOdIqogj9Tu4aaii/hU4ncOwU1iZwx+ln8ib
Og/BM0FY755mwQk4NIx1eAhfG32c/8Y6ZcW0a2jmPKAP2YFaWv2YOOvErWcwVnJ4
a0O45noBeWcV+KCIOQsbP+Pm50LB1Jg7y3xxlBVOys1eGDA5RtEBK1M16vKITNmf
yNlPxpdLOcqhnqis//Rn1/dwrcEO2Hq2hgZBI1dhJWyyC5UdGlPix++zsi2Ggt+l
7+WSx37bXTHYRodSVSciSzPDQ4uzVqAcybWEHOVlzYI+3m84ObD555h7g/iNs6p/
bN4uZj8Unac/EEJsFxFtRhtQe+qWwumfJLMcmhRMcl6UVAbd4+zOpJG+0zN3Kvz8
MWp3Vt5LOYR6wM1EaeG42aaZNADr9r6rmZUFcW1nfGAR7kQ9Fjm8kTQxBzC6nXUx
opEjmqiO4odYNWFWYyU84leds4xD7iIVx5xCQ1girxX6w51QquxI0YuzGGxPNaCf
omIcg8h/d+Ljach2iy2wPB33+a1HlQfgJTjRKZ11LuPDXRCLJUiC32QbEJLHXLg4
R3n2fbVmW11FhD9zxUMUswHjVdH/Aq6gENW60F8w4wk2xf9glm0MJipAeNmwDqQk
iKqJhF23BQGdwp7eK+A343O6b6kYBPQo4ZIlcQ2uNSTinYA4bYY7KSrjk2PoFKzt
7hXtowDUDhX/aKx0aGoHVy3+M5N5ZavKky6hqP0rdexCwrFq6JYmngMcGQOKHtCk
XnnNs8wK0oUIIeZAwtC5ZUWMEIOKMZfYq3NAVY+Q4nEdiCIEB/M8pCA9VQS6wpGw
r24tUy5GRcYy079VJyiM2/iAncprataLaIarUIf6kB0nr0dwC73pdBbbX/OURrIB
m82w+5A8dPjW39729WiVII3x8fkfYCz1QrqMJLAOf1cYQfV+f47bchK3chIenGXG
B19lUi5UPnAYflzUHEIdGMOtW5zll13PEJmEx5ksObRAPd7FinUTIlpVGIFF4hsr
KzZiN2hw6bR6hVZSy75FCynI9/2kKC76UAfkKXRnw695aGp4k1kzQldO4oObKy0V
gJ0gbtE/3xRKCgBPdMZy3baR2HRmtM+MzANyah541IqjgNeHr+EPX0bMY70+TMWR
lArmznll9fSV5IAwi1eGggHuxfAsqeDvAwli8ekfvI8ENpZPiMV6IiX+wXZ6H9u4
ZZpaeh2VUCZ7OfRaWFhZFr6IwS/ni2Ol92dQ0ZOFvojwvTub9I7vafoYYPpjIuii
+0P8BNB59HqNDjMxf1piVyvgJUmsrDtd/mYyPxubTbDSeUMKoNJA2v5JnH3nyWnH
bmv4zTzVZbx5GFAGb6+0ujoNXuMg4r7rKr7ZxwTOClAz/JN3JMSuJV4xEgCD//Yh
Mwhs9c0fE+RRcKIEn+/ARW1gxpl2FJVwFr5Q8aoDdKCZnBpHJ4ywgiG0NG1amwYC
Xvnf1RUzWZRISJhJp5/0MsO8TzBEyOzR/tjAWqv5CKTJemKGBoqCDMpzbhPywhyb
xnEXyy/kGQ+F1TYYUy/nV+YuiT5Xr28dBUMYZ+GhDyHrLweOHjcFqi47j6N3AfvL
UDH7ouRGCeSt3mIztYk7O3Jqp9y3ulVdL0+Fsc1z5n0Xr1SuHLDYFj05yerKck9m
VVt7T5OrV5IiYD4ONAMcOZeeCQlBnFEHeUmdukdEQsXMc/p0H/sMllinChzzf8y0
YtWGnVy0rnf1JaDv2W1uaOc61FmuPND3StGrGjn/KYIwQp7IzLFrhSLuCFJb6VJO
cRMPlJ3NJQ0biulrnzxTX+10YPv/SJJ35R4YZ8944T0iL1tJvGECHFIGIkh8HtWL
Io2xqaJmShzXTW/GwG+JNI+ghIwPx/KnXHiiEuY/fAvDi9a3zXbbYiTuXMeVDOdL
lAGeba+FRl2jAo932S2HOEBm8fwrMANlYikngFpwHBbX3JWhZ4jTO9kvecnee36E
5eeL6Ch5AuW5J8otWAFYf6GFqWw8wowpfNpPBjXKYRYn3cnv+jJaUVxMydbJxzbc
PWG6INTOl9j3xLQO/iI8PvC0VfK+WLLGma9mq4WvWnDk8BlDpkGc17MKBS3q7Q1G
/uUPTcWoGeC5cDx8xKezodnAwZ6mIaFj/g+sUjAVG/8WmsEsGF5KkuBY6Pw+B7sB
C6oPWM3p7xLBaEleDRvnLCxCrUCv5FPswj3Qcn31daO+8GktTtZaUe00ZOtjHK7q
BuD2X38jTeKlm/PcQuo8bX8tP55F9rQCDLk+548H9IcH4Dta2xS/nNSi3RD3JJHy
+YnVMciV2fkRho9cpvyVWAnviNeH59WVFxognoLXrOmAtn5Dyya4nAYSpldepZu/
vUB5Jz/wh6GJk3K6k50F2z9VefDHjieeCffXP8EereJg2db3pOjH1lDq15UFrDYS
1gyZImpb003016w1qPyUxvNaqihWbMWkSvEcvJJadJxXyg7WEDF3kwN99IhWJvxr
pzMCRP8FO2mKXoPIEi7vSaARUjfxC/f75RESkwGmK9DNKgTYKUi1zVVkAZMfaZOW
U80WAgZ0kXBB5VRynBHq8dNx6zNTktiySU7j/YP9qDlDzb1mLGiA0kGk7jjfejSF
XUVaigb9o91j76EQthbiqVU5q3cp8zPjt9yW8yyQj/p9wuc+x13dd8QrKfpzdEqI
QQ7nPtuuCcLWfHfkEopXPT7ys2TafC3rgsLI4Tf+JqtA+LKJHSTWVN7LbfOMym3f
8ozU3ey5uuyywsLK6IY3couqEiFRY5qTx3wV5H5zxT0kL5Eobd82+P9+XocqXp7K
NuawLxaMtiJGxwSnGfshf3lBVYcnhq7XSHy6dzB6ayXioZ7f0HWZEq0O/9cFDsOK
hJwzzPKtWfyoeAYfhZ/HTlCnlAvOJTcEgPSSES67o3kjsb+72ZbR1cB9f8ffaHnD
vG9ehyhmp/7Pr3RisIOPWPebjvLuK1ylhNeceI/CCWUGDFVNQSH2OnrBJPI7oUZF
2t6K2AGK5NWiYNMhIjb65tlekUOuGQ9rKFfXGFsPGWQHlh7bPCwdn+w6+zJRWfah
i1Ibeoixvp4D/dFm9zrdns7dYKvoihgfXfvAxnVvK7b/jMLcssPiFyJDpNP0dvDX
U0/7BKw/yxoPeKmxPMc4RdcC09+litstA5gtbrI0/xNdZ4V8W+hi4U3hBv3PLFFm
X7ALDIHNSL+A8Vft+vB1740zGaPQRAqT3hdtUFM/gENMQ93qmHRjs20G3+fcJx9c
p2dXvSvTeUavoQe5Agz0Wszct7BUDdl/eYsGyJRZjuFVh4YH57SGY/EmdEOzfqzf
uO8rizV4lRdP8qaVvP6Xxr0ed4gDs9DIg4tAOXBdKcZ11dIBBV08pVFXHofLWjJB
MH39LkgdUyuVnopMJwMrv6TnxyEaq6yFua/j49gbkLaAg7Mn99bnHJMit9hEuRIf
sKuhHz80sTT9H7W+YWrTv3lqddMPTGpdU06lJthkJxszGNcdcI3phW5j1uN1GmVa
KYZorNCDX2ekOrTmpy6oTzhH3aUdLm66xKqTpRmLqThmXIOf60zDpsU0vg2+UIzQ
mDJ2BtUXsQdfz0JPwl3U2846zhSfqNKuFWD+NK+bBGlXixTmZWQ5tqhYxGDK4TV/
yDMz0iSfgDpBz5yA0mDRmhTD1ncEKZg6H/moXMiDYxvPYSZDhctABBPyy9nCvaf8
3ImSO0m0SRyW7HVJisWoPCywbIo7g7xlETJJg7V7HdFocDpebkEN8vF6ixKWRxfa
tIl+0KYmZylKKbyYjmZJZ9WpYfVfUi1L12gnGrt2HZC8Kn2B4vbiiLl55Zk46eJL
TDcCR98hS8qb7ZQPTvL0wNE+/OlQ2W5ZO+/R28oqqlVOkruDi1WbRL+njYU7+QHq
DMHD/iN08g5EAI6kUrXSnjjvbyRiqUQdZUIpPwGYcheTGTwv7UJP6A8rt9ouLpis
P2tkbTKVaYJOKX1mrVei+8ml3IhnW6yxXAN8ot+9xr6nFA4/rNiMgOzjJullU4EG
uPPpRAQMJ1Ll+1qRPw/CJPR/6B7EKg2wWdM7Q4rU/2Ayevdu3yWVXDWt8qITVTkk
xvVCnaGMYOHFzp+2PlWFyaAF01Ks5AfU40XjStIQ5gmcR6VfT8cj+V//gcEawO9I
IY04rU3kEZEbAAHE7aGm2H9e73p2wMyoRzLSOr0EnnfBKAfFjh5O2UlpBmKIgdOi
/T6e+4kymJmFoc5ya5RzjyXEiw/BNzippLFJAdr3YWuEv2yCbECDteHo7I/BAJdc
oVr5PPDMnAXIDDB/5AeWS9/nPrwEEMEZdEl1u3SlEmyh5MTcm/4I2WS9EZfn4b8B
OJMYXTTcr434bBRA0L/M5p3xrnznPNkrKHkhHKUvVHCv0VTVcF0Sb3RmMCd/P130
TKYsQb6zMzPBVcMf3ThxfgYBYlL+nSAFhrGdfGOmlsjEWNqFrOgVSWJKwGA9JirQ
rQSNa3JQSm3UqJVcvZiqQyT4l1h+jTmHz7d933zmF0jcTGiKsjQzOlTQy9YcKvFk
1ZQoNXBHwqq3ckNHejUoAq3WILvikUIp53sUkK+caqIAyRO8eGQ6Q66vVHR4j9uW
BM7jQXr/21DXiM7You/ofCaXuq53v8EWSjG5Pb/bP0JZJHYHKmZKEEpEJLLrstAS
t8UEPQC8yGfvTD+wJjLd7H9PUnUw4YZPbbQTL3de5FGOpaQFHi+4SfsGU1MlpPq7
77z4kgxDv+q5SSNwBgbH+qmSIvHD+lu/pvECEn2Pl5szryrQVR17DfApRwAas4Qo
P3zxupGZ6/wKbUmbfvrU5N7z+8wsprR1THJj8qCKFkl3sTpT/SlhG4pVMZ2YNmXa
73D5Wqd06DsLHMNE8fxjfXWUtcLeF0iJJtCt5wDGdMoLVYsZW+RSYFkorwVijPak
gGgln28n0AVxIyRg5PHvpQyx8WO9EV6rjjtZkuyARUNhxrq+MxS7KNo6viy00GAH
tzQpKVFWWkjrZxCFSZJUIRGjgfwfmBmPFYU25om7K0/jh9pTjP5jW4JkNMcWJoDI
7B9R4GsyOiz6ZhTc7jmW1vRrynQZepw5iO/+e2baUm59PcXIcmnfhEki86eN2EI9
LsnzmXeAADEE6oqdZdC4wp1yFDz0fsGtTl7prJlPHcGXmFNMG5Jc7dSIC1RGkKFt
HRPBVnTsJxfvvhYbRJD7+I31Wi2G/sO8ut0FDzoZrz9pbsFjOjR7834Qj5mvbdHe
40dWQtP1MY4K5iIT69JLna3d5jpW0xuz9Pjoq3wXPqIC6T71AwKx9z3AFy7rl05Z
/qxFpb08f3m2JbvWVxhv5AoW9J/0fxKqhpH7W30WKJa/98Mb20ixlEXOD9uHUE0s
nAK93AD2jY45gxNhpXZeP5GLaTyFSntlcEIOQ0anWfh6hZgOTr2BMyd3Lim7qrgV
Y2RNuTjzWi1w2iAuW42pkaqHSCosTtTRE5BxIVZspB9D52sDAy0YWD4RyysNbrW0
+KiLQ/MfeYC4WH7547Rrp9a0XDVzUFfmiPuWEjtVqkExOTT0jYk6+eJgcxyaq2Eh
On23wDW+pkYCH/o6amRcqyNB8I7PZFNrpRQxthxygyNUttSVh4obNGvjZOrTS55O
vEsooEu9sCwaYt9PHsfZk38B3LPH31GJqeRBiwnQJw1ohFvZRUH+wgCzZQegRsP1
mJA6xb6x8+b3qzk11B7S6Fpu9kPq4RjZRo8XWZ4pQ2fUGGA9SELgNOrOA9SC7A9n
Ilw858atTXFOJOknxK1ksXVjI3gH8EuV9DfZedKsVGYJP5XE2HT2SKhQtMWf9kik
tfFRX4zdUkpSWXmR5RdL0x//LSbxhKnvKBvBy7UPzrn4EQLzgb5zJv6oUHN0aUIM
iNTOwCZU5o51d2kmq6m40yDSisOSF8+KJwhe7n6Pf1O/S9z9ev6H/3onlYd5aiVx
aXfTxfKtD8oq6BMjoDDKtJkUqlod8AUB7SZgISVUGyvyc6kb1hwPsm/FGY/puvsW
vkgMhxN4vi7gzn11gcYvh8GREBsVCSX9z8hgkna9vwTvyb7uiAjBFQhctOvkPChq
dva6hi5dyfxM8JNDFzoHpmBj2t9XZgDgg+cVh5M3kY+jWyM6lR0Ahg9SQ/tTRox1
r2zg5hYD9iJvdziD1OwekbeYXqmRrh6ZpMmJwfZvhb7WsAT275IpD+EOrcF+BW0l
oBwPFFhyZlDH9ryLEezLf1j0RfcNqs/u/E3vBtAlxXq0ejoQUuNvmd1kJUDKQsBz
GMCdCuBhV71HZBYWp7CirHRNpZQCVkybRpBsbmpmMNtYksdKoRzog8QjQR8ad0Xv
uiqWfAJuJWIkD/7DA1jY9DRUrO5huLnWImi7TkUfdz4alip0L2FLTYJkcQSBL5S5
PbLlhsPonQEbfqeURCrDuub0RE5jx5bOBsddYF7sWcqoRzOTqEj9jNS4YUDhNoo4
rZ5ymugNz7kkQjpXX27ZDnYAJ4SgYeR/T9cRcF0dAY7fswr2ay1EXFMzEqTcAved
J3827pMUWbmF27LlhLibB/x3d63M7lYHH8YKHyt3RThMgcR2Q/PfcOJCPFiYS3Wa
8aFnNjBkT5tJFJu+r4T7Vjtd3T6KVBEBm6HOTnXF+P+w4R3UZjb65k1ubNqDKdgO
W1QDhkaU79clRGikNVraewDQmtX2RPxNAyBjEJ4VsJGMbPu9M7PSOJxQdOSBee7L
+jMZwjWqU/ZQSPFQjDz3RFV8SLSI3Ri6eX8ZIiBF/eakw8NsMhUuBOb4BSbVtjJ0
9NS6cxMcQTVmvONI+IdehkUWzP8QCSsd0qY2HaMcqUTwSrliZz4LtXMDOoRy0utQ
tjYj9+AjTH8rdsb70JOd1PBzGhnW8wHdPYP3YIgu5kqrN75yW6YdMlW0X90xaPod
nYXLOz9EIqAHQeTgKYXu8BKi2oVdjiCUPwJuvKdBlYRV5DRS5RNdvf6jHZS1iOpa
bmDT9jXkoHd6ILzIXV9zuLoe1929Y53DupGi0itGGLQifc+hiZfb6ALjG76aMppw
pd8JemdwUPV2CtAZzPV8DwU6yKhm8NkD8Q7dczN0W5g+93I0zwre05rcfwpFrNZK
VEv/mw1508b0JMRVDTor5YoPgkeU18sKsG0Y7jEkwJLdVT7pS04ytITNNU3xNEu6
yoUA4WfjqlTMbnCM1+vnj3soVLIfIGG68OqSnNSs29F2ZLjdFscKqEds30sMprbW
BHSO4jEdGsOtGok9euqPbJgGxbvFwTIwpmeuihtCMqPfKegEx201UVnd/ir2sl+u
0MWRQ7CMisoQdFhkjKK0ozrVL3GQq9d7Ua9rDflhD8sv/chaWghRO8ztUmBkgIWx
5ShswLF3kzV4wMw2sE0YILeKoZEDrVtRrpJ9XcdyVKEdaBy3+42tTFWugLeoJO6N
FMNKfxyCbGDbdRRKY6/WiizOoSqaeybo6Qhy9xqIIhZnt76q2+F6xGzeeyYc4m5d
rqApW7zZJJNGNIsq0wE1+HtjDbx56S3YQIt5VCnFXonAcOIaqm0DHr3QXcn2NHAF
p9XT75GuxGGtoTkvUMyOCSZZpmT0nmM+Wqw4zzAUgaoo9Ut3bQ80KAc1xLhoA9Zu
W62COlPeiEkI/CRnY9RGIJDbTz6Rl3pawYUPOdNlsv5Xo3kfjxvfRl/y10dhZ7dO
Ji52vzYugKPC18s51nOh66BmRQ6KSukQ7UYyeuOyGA1dX6LfgPDvvC0Rc2NVhk0w
de4apl/u0U9oLpyCbcxWn/WRIUtKHXxwIrr3+ZPJgHJQK9lojXOjpZlCUGniOgA4
Gh1O+1bZv6DqgAd/N3GkCPaxg5Yq5/H6kc3aMplR/MYF1RM6T0GAYxcswff9FCcv
Vb0iWswF852+TbV7MnSKpVxl/iPtp2JAECeAmzOSEpYKmHGZPdd4GmjZ83+TCNsR
s+yqk5BRsHPLRgUEEtH+DU2aouYnvK7qdZsPYZkqSdZCnULk4XRlYiWYys19aJIq
Ku6ZKLmpI7VW1laA0SxaFykGryoxOTZQ5blHRrut2RG4j9x2ET6Psh0W2FBQPFza
xh5ajuBBt9aeeVbnydDlicNcsjXcEUfvqSNbLl+Sth1b1V+9+caL4fyn3IFJMiJg
JakAU2YFmRFtEJNAGg8truJIkHbfS3gD0A/RIbm7ZY0M3xXHaWWjoxdHhpot8hSn
a+el9u8pye0vzsny7vUcpgynBJyUx6/MS4N4IlwzMylJ4IWvILOjX9itjqmwFnME
XjHr17iqGceCP4xUvBtEZ6jNjApZwzaGTn7Mk9FXJv/CdwBnNGGPpyTTmtig68XK
ezTZ6LC8sK4F2Wj1ihPpoubNxPlbGoj781eLOQAsLDQPCNEhIeIkDjQ1OS6SuQlJ
Tj2dPGNMVpwzgxRmF3fz2gSX9vEU38CeWmwZBS9g5lxupQ9PsmzJwLQNyE+Ysi0m
/Wo0hB+Euo0QThCOlc0kOBuskljH8p4mBRkBSklHWg+jJeZ48l8u2Sd/F/smYajL
cN9XXycYDsOsLsQ4h9iwqeLz4lJg+eSp1gYplt6ltSk/jjJhDNfU/OjDpUa5IAHc
O9TPgaTYz/pWHFoInjMQK5YzzRzXT4Kg3PrHyb2W3TWoSvuD/PZHzE20ZrXQ4NyQ
/GrEi2iF+IsG66uN2cyl9fG4uCHDFD0YoLVmhUZ6TacbR/dudVW5aU4U4hmPrw6T
YLPhxbS4p3JBtOXfdwApX2yf0ZqNv9ERREXrceUr06roNAZTfO6oIaScsgZ/bfX3
WUYnKCbPOMnfHFAK+aptQ367cmxv/apGKTsPWjMxWlx+1kqQE9lMRWGog2J3+CQN
UVr/7s6WEUI7LSggNH9OGzy+ulJrlFom3lfvkchjXUZTwsv3mFeH+/jsvI19EZ25
eJ9SpUvEHZtNsPgkVeHC36qCD6mbTU5g5BTgM6pWq2Mna9mqJfhI+3cBpiNIvpGK
zMB6XCidqNfblpe4ep3y1Fz/b5KKq3wexkUsd6UrQA0SPyrl8mRrh/7aaCIIg+rb
Sg3jnX/57NTTzXGof3j5G5NdtqwgqGc5zRQQQ4eU49N4ntt8F9tWaUpghAy3+6xB
l2rLKYgtVX/svgEU7EQSw7sp4zi1eGpPwO2SuIwjYsT/6j3zkTF541QYTeZLxXSv
IEeALbRAGYHmwMv9NiPddo10EcF+Mi2evZFsAgiDZYCAnOT3t1aChLEYAMogF63j
Kky7toopc6ODN6v88DfgCg6djNOo3+5RGfDVvGl9YG4HVAj1rgphKWnDD6bHjOPv
acQWK/TYDWIu+TcEmgoLF/bVAeVaPC9BEovxnfbMcwrphR3B35TdFAFz+/HR5Xz7
KxDwloU8dvI03k8uc9GT6rnylXtz4eLZMexKo3rDFwWcviQ+DlAZiTjgYnLiQu8L
HRvpv/MXnX+aifMxdl9eLB4RsKgs1t44RdrMJHIgjEHYCO13mfi+EWpZJ6r6U9/x
S48SIT4TR7IFkntexQNHEjgLxRR9SMypKIR1WonquQGwMS2/9h+ecx0nSGUOyGQy
s1ukiDh4x+xHZnTfFyynyaChYZ1/HSzU8QuAz+BfQNpm9LuOeHPyvZ2dT9wlEJh/
U4PxABzPT3hRWBdTXgibdvlIK7sQepFXGTnH0RFvU9QAYWtxijKEVJa+8McAdAPm
VxxXHI+AwSTK5gyZwE3YhzrBjiw74PaIoiHqAwMQbc/8JapBILEodoRI6XBj+tdM
sAsL1rJ5kX4Mr+JZle31qqjPiLH5/bqoGqec2QY/rXx/0Zg2tuNBStVDcrvMLdKG
KoVpWJLqnDR7EYzn+difhPKGGhY9lymMEVCIMSZqP4WYpkRnPwwwMnmwN3tBLZDn
JdVkTCt02jwx9NJqhsKMncwW7pZpC/qmqkbtqfrqnJvZXyP0BN75AYvk86B+dCR4
Nj3InWMJPdJ11GsjD762cLvDd7yCBjD93EU7ZWr/f8RbQ4HT1a9VTx1xDF2hGvSA
0hSoCsZBM1Mx7QbvNkCi8weGieX8T6babrsfVn/wa174cZZwzg2Fv8lzAvZTMrRD
BRtul/AvehcnIiKrtDKuvJe0Ae6OJ92u2PwKMYYoJ8zTPT7zDSNOtlYJlDF6xjaB
37BPkUSJKpwqkvMFhJL/jivKTgrW5+SuZuTOr55VQ9o204hP6B2bsBt9KBv2iQ86
n2JoQxgM1MTZbpZxnDo0Ki8whle1jh3Kz90XXUrwu/IMuCBNkQyzpVmL25DSv6y1
YaE2CaemQyN+1t9tDpZCDO/n02FXRIMH9jXnM4CdZoIE1AqJNQLrF6w/ri4ecPTJ
G4yGtHtf4W05P/n1Z0tMtw+W8QWfaeXPwVRx+RZ4Lu8e8CbH1+oKg9iKSU80Gdtg
6/HNVr2z32CcSSjfZTw/l8vTtr4aXlgLXTioyHoC4QCpkE/yIn1Hk4TqF9qz6kB2
Nc/SxiJxsqPC5GXU8Chc8jnehuzMlbM99hN6MGDppVdqb6JXZ6xj51uiau3UDYU+
Jgtr//56cJViqnEVahL62keq7B4OSHZ2zrBmQ+EUg24rxvyXYE2BtwGHPaAzzJp9
C3/yL9VVzbzuXye52bGh9JRYpjO/toWPeZ+gxwFZbuASeihW+DGoWGZmNYhIUkY8
/acFJbeP79MK8u87U6sT4gRZWgNug6lXusPmD6gEADO95LKUUt87yrE0OGjGC6iA
V3QP0xyUBZKhwB6Es2tvgL4ZlWv6bDedz3OkO8QbVJ/Z6dyTP38fAk/XvfW+GK4r
Vp8dKNO4MvFtzZTIPPxYYhxad1oPsQcjTwQlyNelgB9yR7aLkg15N4syVqzsIo/3
zZwH1pCxnr7c7/wk/BUn8IXvLioSMmoWB949HrFuxwWnov1Jckhbog+rr6Ya6LkU
FzgL4neF+jbzk3C+6/0/1YYc+1lI9Ry5yaQciqleWNTdIpM5+WdxZ86UevRqJBdC
+TgXnMGOqgr7nGMi5TE6A5OZiYfFnC79Qs0LYUcGj1oEg+6LE0TCM8mgdCLGLowU
5KjQfzKZZRbCQpd3tZtnAshmZHp1Mw45nSLHkxyGHSO89Ye6hcqoDZ7IRCqPAV+O
VWniw189UOHHGPV/WCV6Y5k+8x+6FAPlxURE8MUSohrMGuvzEJ+ksGvcNZ3AFql/
k2ZhgEF4Zaou2LJ1ckl4Lvvk9DeXeFrYcBO0MSih5zsevdpmtPiJMlR2Gjf8LHBM
orpMkViTirvLN29lqH+Jy4pOhI42hb8uM0YA5Ngh4a2Bd/sb01i6FtdWXyv0AdFn
FRM/y1rBSm3c4nLiisi33z4yjQdTpQtKW2gOzJ/OfWQvwjQAecBoxL4hbOXd6zRi
H5hI7mshDEhQSBMwdNRwancGPrVGIsWSVAPybOprCFwfb8dJeM3wEY6Y5iZkdSWx
WKs/dlj8FI17mIVXamrHCA3VVIAG9Nm3Cmuk77Spqjz6buVqIt45vs5RHVXB3Myr
1IN+zkHuramarxpmv4JkL+76IKJsGKaK9wLVZbxYYUHETuwG69d7mxPGEB/GSPSv
hWFqaNUayep27R5GZeEqcAtfRIgB8Tph3TbOZ3Z8Z+5GJF/XfGAwU0tQNW4uvUoH
9sfAKo8v2KkxO+/oYasFlIWIVZ3axjizaRPonUEn0DMEXDkYxXmCbVQSTvlpSQT9
G31EN9Xk/Tlcz7Micsq0fKTpCksbPWEqf7AyLU1T+cnJEZpsfxSK14tAQanst8tu
dwK/O74DeAVFpNMChwZUC8Au2diOUrrqFj5Dc8FZOsjesBfQh6GjVSvdzpJZ50QP
H+y7j/KIdSfELYJNvu8SpnTy9qUUSuCuhzkYy/oDAT9D+w0aBEHkE9GwKx12VbUm
v2+D1BBOHZkBqJXur+1ZlRmW5Yp9ctNO7lQmAKlDJTO9owCdm0hOxKL+RsuU5ZWF
pg4ocQe64jKNRoFds5MxtzvqjH73nAzDavFdwMdcjoP0gaOLuofkbkmIgShiobdI
0D2+jK2jHrgBqU0mensgFBlltoZ41Nz8t4FkTyeLfayjn7JmUBvATuBRCgrnqxhg
waqbkRx890gOVNEojN3Xc8wOH/htMHjVPLTjyayVxPikhX8eMx0iNg5CX7Gqn5We
TuaoX51a7qHHhL0mAZwdo/uUwKZELzznxGAEniMfyHTD/KimpxcXv/cT0X2mwlO/
kLgZBHDu6IbAGMv3d5Wf0QRDxAIDpyHPjULRR1gkuG1vr0iOjDUAa8rpx0x/w1Gl
h1pn/Ww+jenORq/pI9Qromcjw2eo7yAilEfw8mayXcDc28juKVSgqQk32t1hCWEw
kVAohCBVq29i4OxhfnDvJpejJ+rT4KLc98zBit2Rh6jBQPsJMrzTqjrHmgZrTDb4
NM0mnRmpwIa07yifFEiDfIV4bme4riJ/2o/kjLqwFX0ZFrLeU2rqRyD2a2f1bVoR
LCNoUDX7HGpUkVBEBTF9rUQC/t/ou/X6D5XWOYD1rXngK6RAZ7OuVdnYi2tijYbN
xbYalZipcsF4WyE6fzaAmT+X3o/DTi1PfjlwRqF+vDhjCQvBcfR22YuVQUiOsHGH
75Rp+sqCZ9bhq2V9fmCN5C3uWMQMV9S473eiA65ugYT/zE2HDJQoxZUr2/jqLyov
7PegsAgJ39iomgez8ayEdrZ4+Sl5vjHdiD4yV3+xdQRrnUbG6gVDvS4MNp/P7P4z
V46BJyn92MeIVcSTHgNEfCrQjQPOhdNEF8tcU4mGx72riPS6wPDeYCZdEPa/lGAF
6pm2ToiD2TTTaHz3eBA29EhRDKFH4TDCPHWKqK/NZsegpXvKhBeb2PX42n9ylbRO
EUouSZa0jynYf6eATnPmB+HofnlrbxC1pDN3GD56OZVUj5wp7DAhYLOFK8Hc5OIB
RgvyUbmtVLlebvEz6cjDAzYFw/ePHWXFUeQOOYe6j3vSU2LIA072eA3AEKwinRab
F8Zs4B4EOa4hvmWB9VCbrN6ea7mASCz1z52UVjJl8o0c99MkMspMHUDI76xNoNCP
onOFKX8yYS6VuCeav50wOpIvvt3iyWnpSTPYT7/z7gSi1CSX5ko2aYFH+Y/jj28x
K9cDPdq9ERDArIV7aisNV4dGnDstaA8ZegKkMFUy14C42W9v+RQnbZZ3hM4JAjxA
bGxGs6lmgb7KhodLv03g7oJGMMF8ZZnKOM/8Ig58152epTgXfzQSN/EyZkKd8XpP
q/EZmucrhmjKsc0ghNqhGo6L29dFR9LJNEoRIRwlTomE2+JOJt1b4pEs3I2t+woq
vecliAuLdD1fXmDtKg0U742XECFFrLOH3VO5ruApG56DmuuoxembH0YJaWorDb4A
6YvGD6QEZDPwKZnClHseXhZl627wihGaHihxI6xd2DbaPF3Ili70iQka5qCkV+7n
3EUWUf1dcIWKsBiRjMPKRKnJNI1jZHCvpa+kS73ys656oD1G0pbudENa+bNsKLtO
swBxSf7RHx2daOO94W0Y85J9/9+67SVkEYAVZUuf/RDlVyS26SSuIDi+tj79Zj59
K7GSOCKC/7SEyMSTg1X7L5ofQLSjsnVkCSHtHeX+EUJ3tTppUT3Qk+GtnlBVoy55
eVz78v2FldczfSbWjWCN7XHhWlqNasUIBbaQ+wIJibOi7G0rmRWHY0d35jP0UYUj
hkwXsN+b5BqSL8V5+HxMKPvcBV19qw5bKDCMhXF/iWGrVMS9pEmwATYdYxsX0tdU
fRtp9SgyN5fiYfB9rYnEUBUOTqc/DZPvdSExyPP5i73wgUHXea4wZH0gLL83Uv7Y
tUtjmlQhZspNZ6x7vmn6t0x/UsY/l3K8n0LQdisHG+ltX2y8ONb4LhIhIMFHhIG1
jtuH8BDEW7Kk08S/01JYP6jsIPfuKH4Nf+Q9pdp9+t1d64gBz5qt8HjevDdz6cQ9
cxpoH3BIOeAv95gWEaPvGE2IvzUeXiu+3p9kVryFlnvNiS+QvygbgM3CTQDryG5V
BUDPXYBEFVTtep61dKX5BaFXxSR3ukP+ZUN8s9jDHvVzx/AypqF5GEXCrZynpS09
Udz4IeYcFHdcUp4OVWlwxb7ARg8tDAX9OrO7mc7T4GntRPIJMr2zqmpR4kwQZtJ5
9iB5C5fzky3teq6zCowHDsDvGSgDj62oBYw6cK5GAYjlOKUeWgbD/6B0P0tPjAFQ
XETqCwNKkat1t5G7qqPjQwGsxCp2vlQJY57+DJhg7QAuqFK/+MVcyh4FBJvzKl1T
t7PnoIzFYNnelZ4A1KV7Ny5jqUTu55o8oWnyL/a62BgsSd1mEpbza0enh5avwd/b
98D9tuhEkJ8trHadCiDfclyxC7lWaWIdQRQSomtDpsnBhF8AR87mNECmHr2tXzWx
HybLrQTxi54XXvW7xKbSCEXRnk1VosIyZ9987cuGVMHM2AxEJOa1vQJG5Q6nrMoQ
IEBe7sSGTsif3aUVUATyxGpTAMa/elmLejqyD+h+uoHmAwgbfa5EPWJ83MYWcwXk
IRf42wHBmUoeCI//vIReG1T9NNKytFgAJcNI3KOPh7gRk2Do+8c18VOsm40zZ7Ny
asvKhDCELamE2VLgEemPyW6mOcTKFLikCiaKPFyLtXqn+2TbGJN+bhzKM2oGy6Yq
X7Wqog0HV6qA3/eBTALoX8VBiIiacTHh75JHK3bBuBlhV+sWSusvvTtFoUdsFRbI
jvNGTOsTq3DK6qEHlpIHADgqU+IWijR5spX8z++3pB70T1uOUpwzvlbym0RAuOtl
nlyVOyMR4sqio9nVtyCDcQVWQcIwAh3FRd0AmF60ZXjhS4mtk6/OIM0DCb92MYz9
BJqgEgKXn9Or+0+JSZ4ZB0IVIO7XijRpbiDA3o0aDjTf+gea+CvUWXEYkU0bScSJ
+SfNvHq+91oWFOCy6eI4wC+TnLEpYhGwowR7GPxdUbn17VeO15SurOYKFz6+vblq
dIQ3QJCslNHxQ4GA/Yvj1bNQZNF5Uwk1/EZs93P38L7t239sqbfLIdPdRTv0ffn1
5aJSDrwUxBf4F6lEOjDwfeoUaV2ZTgjSutCkUNJzNKN3Bg0eFyGDO7RWOaJhHTqh
W/a7oAuAqAnrk78gbabtf2F8+nJDSKKy4iDNi24gm/+UKlO1VqUzNm/B8F5od8b/
G46+TdL1mkDkS2KvlELfVzChwIO9H+U6XGoeMvXYnPEICJ+kPEob1/kCsR5dZTUO
dFEDMxIbIX3EZKLjEGET0umFgnvrHHUsgK0C0/0tfbIEgHosrm6HYW7h1c4jvvBT
KQoTGARSVYiX9wUbjI+FSc+MU/yjnTzvVXmdPcsxae5aAWUCnCxmVgkmBwtUV1+a
5WBHEcSEqN1zm52wlDhW8xnujeRAnLB3163MPzjBsvBsUXtlbF3TJfyGpAWh3GV/
CfT9HK06UqvnbWmcJy4DI7t8A7q5TUpOO0mucxc6Cip++T0NsqHOrf2+tl+IAhHG
1orG8bFXMfapn8MCzUeDBHwkmL3lToAgGx7NyixbDZMtFhUnh1/2DSM2l5W7fgVv
bvtztjDpv93Walu95FrPHxmofwVMAyPolM58UJMGohQ/XuYPxyV03AOFGNkV52HH
vHzxApX9uI7QNYU9S1iMxngkEXqdqTODaXIiDWJjpAmcggYZistxCmE9eeVAWxAO
+P8qqYSeueQL/mfO7MJT+b1M28QJyIyrr6idVsR/gnYu6bigMduaO3u60oWknbp2
rW5CY5a9jnTgMFoX++DQy8tOI2fDE7ytqhQ1qoQJGmrvohpRJYJP4RwHezkbzJ9G
pNdFTuLsiuLrpaBM42NcCSGPR0WktrB7TXCdnHrqJ9fvHbp35Od++iKtlBJ3B6da
B/dy+JBCT6MStbsQJkXBMXQyj0M3IVGQr660yaI3jYd1Y9Av6azifq9csrmarYL7
Bl0XU2Nk8Q3eiZfioTOzTiqAjIEFi3FugfX+1AYNjjWf1OcNts6vA+w/JP8zMIB0
83i4oJpCW7Jg36UxU4E2UeCHZpHFB0CzipL2LImGRfuY5eYjwObejlx7WMxzL42p
NxaO+P7iWtxVR2VLc+LyfPnLQUZK7KCfW2t5EPWtHkzB4/znRjr3ocU85LwdKwmr
1/gH+jpfyvn1VBtLZHIbEwhhFmJp/IkpGeHwa/KYEhfRLUHo27kpCJjRRp0CG4aU
J/lgPSNmeQE7BQBDn8vqVBLnna5rFg6wCu7gSgkZPHS9A+TQZ2Q9aBwiur4q6YJ5
82OjCTvCZjxuQAJV8AuEUTqZJhUkRdLsuoBbefZKiCj5ZJmntkYoUZf2EchqzHLu
ZHajtjuw0ks7nBGkBzXIgTjqEqWJHKdReITNBCylbILEzmc/JijV6eSm8tUV9JVc
IUVtMssYujmU0xX2Zv4rfn5xqXGRFWoIJcHH/H3u1AtbZq2bdjUNmvMai2xcIrmU
w877vkrv5W+AevsmHUV4HmLG1OEp2P0tCxxvJo1BIkD6tABITIZBhV5wmKT5GGW3
v37h/usxPlWUY5z8qkgPXbpM8p1pZm6F9yPAfsreOhKj+ALs/mB5Axn0AleaEHYv
58KCg+ZrA+yzJiJJ1A4Mhy2lOWHgnRwk+348LRf30NeDKLOsOSPmMTbb6A79c0Ls
1GTuWuMQV2o0s60Yxwk51+VdKv21RiZpuE/qDMXKIxgw969hJmjphviUfvvCyHHm
rMoyOdkDOUQ2Zqzcpf1SYvAMWkX30vWXJDK9e33IBbuXoaOw7MpM6IMoGrDaUufm
no+uZtDoUvBQxLoJFldcudLtUNsOIvHQP8RFyTfy9zVi83yL+eaif2nkjrfk0Db9
3QUwkZCcqm+DQIUe6aykao7B7IDPW1MpTmTRa7S8rqYEVsNFypoKvtDDGx2Ueq3o
tZAwr6x6IIk5VDL0dpHoAPcUOXoPYazdlV0eyfRZGgkimjkStjIL7/hSH3vKbc8F
npfqZUOQ9wX+J5QG2BQXWI2kFogDzx4NMlBTZMY7EHsybbsi7hemloMVPytRd4op
OdioRVtnqKEhJ2lJokaaXs2vVrSX7BEpsrgjg0pLu+rpNj9MCOwEf0bClZn8PKXc
Qa9t2MDp//OPLfHQ/eH7TuO9bbf05Jifb5us89NKHew=
`pragma protect end_protected
