// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:17 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ly52j1MG68DLjofgP1FKMMFmrf6ns3hE2gi7QcGiGhc00/pYa9j1QO5weZSyuqDi
WQCqYCvcwEV0Hju+1BLz4xrI1A2Q/HZXE5Z5b5KGFlLDQXHTB6hTZpcuyshABJD7
1iDz/zBZZDwFZrsu2hRdHDpoFjFN3M+sktk80r1iyIU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24112)
jS3TUtq0Q7ht+CGPOTSX2+THfGzKQVF8ZkKZYODNcqpmgQsI7BgGeiROeRhx0xbt
NwcLykfULIu+poaoDGL+/+xQIwEhMGsMV51NrbKGtm6r0QBdnMUCaIkkXaPe+XSJ
k0uTcnFmawNALjSvBlEjjcWpGEoWRJY2BOc85y31/LsVB4i6WycyOHcmFpkjA2KR
nUdcl0DpOjaSuw3hc6XCoXHdz7iaEzQUmVURda3r3Smp1vSICuZxP7+XMsnFtKRZ
/93kur1dTebPxtRnuqEvAclOfB7n82lAd83CUpMgAvjeg2A21OcOygT9h4pSmNmv
ABO6h5QmCWZILtLoT7XwkdOsXlJf4lvJBimEX9PaitsUwBTqOQmo1TCysmIdOqIJ
xsdWWvAXDktSWd1g89iZ+ivof3+FQLGvXD0nQsusgpXkfL8moQG2GrhJ55Kn5+FZ
fvasvQaCh/n/8liMBwhWzLuIoPLr2857GFtRyMqn3tGMo2XcbmcATcR1lb0v9Ca1
/Ak6DIjSUbO47wIGwwIbO+Y6EMuIHMPvRYPJ/3FFVwpQPB1Zid+jHDa4K9xyFQac
Elu3gIBB7sPKMTi0HwY/+EaoGHhrEWEgF6J/2v1zs+NvrY+X9fDOeRUNE1Rmeq1x
f/DyENLeZSI3hpNJ3m79/L8r+jtmS5CdhZ2kHc26TxYRUN07L6dtfYa/oeIdeM3D
KAoU71Z67ntmw4NBu38Rfy4BVCGg6/a7UVIH6qKZ/EWycVFpnaZAk9JzMGOB5O7g
jU1nYCD3IawOCo7dJRgXTt/v5O28jGn0R6UNIbsGGgGgZMPxumT0zFYjmHrDbjTa
gc8c0T6Ca8KlFmsLYo4XP8R/OHj5v/M7IHHQDCk7XabO5doPSxt3qElr4U6Vse7z
Dscsye/iYbpTFETpH7Nd0Lkb7ccmV5Eh6WBnhueJ/nuPBpELYXQIBi15MGV8HYh/
gFu3c3QV2SEeO8ezIHFaWp/EeC+37V0By9nr+qC+SyRXCkzVILkKcm9e7rzgG++1
nPifiX30zw6/OXUOw3SUM+98FLQGtPlus/lDK6I/HPmQnOMrXlGkfMklp/xIWFC1
xIrYHP0Wa0oLbuoIUY++VF4B50P0G1iyYjnwouGuwhpuxGwR2JdzX/bRHeMRoza6
N1EwYCufF76OD4ifvZk/jfA1tVV1Jhi4U+CcVsK2POj61wHA4n20bhCKPBUfykAZ
MQoVrEw/l7eWKI5D1HYx9lI38Uusz2andK8lklGrASbZFnD2cCksDTgPbSm5/P22
AqdEE2k8txHWMNkpLrbittu/9RDX4iy/mENUTqC0TBrY7DihfXWiPQ9QK8biBYE2
1d25AKIqD1KEPw1O9rW/h35PXPAq5/Z8OV0kVABAFnXsa0VEGXwGtE5HrCNi6ZP9
J9Uj6pUFvkv6O4epIUj4qIw+VjEjy1Cub3L+5DsMdJMSR0P8sgOaSTtcIf7OlIGx
SZ6AJrph+MIbBqzu0xw/96YsCAzrFRyU8vskzDHgorRBv5eDiIKaMrc9fjpwcV6v
rxao0rxJBiEDdOiFcxaJ5LvJ59dtbqtG+Uz+966+zAimlhdlP6+1z3RMZIhF2erz
TbRckqOoMp6RXcQtwnZ4v97ZKyZ2MC6p68G3aXSE1WRm8qEnv78fIJfoNxXMTMME
RBTinhvYeyblbgdkW0v6IaVzbpivqtA9zhfusB0t6NEksq7etcYOfLY/cWDEHiHW
RFLFX6HxhNy+iKkPq58d10GHWVwCvkCbP1Cw5XqPTeZVgX761rWiQnokKvdkZkq5
u/969xb7FXKwnR1l4jKy/43HziWeAHHXSyM/Apsp08+zr6rJJfdHibtvg4PQsvLz
uToHSRcjDuyRKTrRJS1TKLWo6h6vZNXIAQHdPgoNNFYd51/8o+STsKf+k+XZG3Lg
N1w/PxB/cwPcdHGJ732OWCUyugFElPOKDdZyy2FxjPRUIO+mvAFWEmMwCl09++J7
8sTq1u4Xd72mfW2OXlkHbKp0jWrERusGgPbyvX6kAzL+eV3IOHSXVhAKGxzY7eJP
gYeREU7lIQDLzgRx6wiov3r7PkFE4jpi7wf/pbcZvjFnGZNKy3SpLLvukQjCF+VI
qo7zqProO2OHEDFuWlaHPP4WSbX9OLtTnjL9KlQexsfl8KSWj8aBcA2Xocn4Tc04
yDMMoI1ro68w2Huqxgpl8+fkHE1DTT4XxNWKBJ+dGm6kOdbXkOfBIl3cg6XXM/jn
jUhlJ0mzPhHp3Ezv2TEO4ABj050hTiQCi1pDbM5hTcpvkl9SyNTLNF0s1cHDt0Ob
BegLpsETJgTwK1WWElAtASiCb28C9I1eVpzskdg7olbvWqKPyOBWVJcUKeH6ADSg
mhw8ZvoC07mq74TkibdPxw4epzLnj+uVjMYJiOn1MDGOuGlOT082sX0q+fDkf1e7
Me9tAIf0Ae1tNqjrB6Dh/ebLIF+ZYow0gqk+HJgINvR7YMDs5u2U6tR3eA5pEdDn
7/ajZNiOXWJuS2K3yvi3PmhHRyKLywxBTuQOhgfQq6Z2r4mCo5fAWvV2OajW7Kyu
1H6Bcz1f3sD/OD4rnJOs7LJmm0FtA8gsB4LMX61igJZJBQu9QPbvvwWjn8tXg7gx
AunqT3RiTdJFb7idF+HCChTN8xcXa1G9FWxO5LTKgsZYePYPJ9p2NXhiaR0U2hKJ
xXdrfR0pjqaLfFSOMNoWNw5UnjYWEyhd5WBFMgoyuNNZWfIsq/XtTk24xx5Wwnte
++Rw4ddyp4dQUhdBi4jeS9xTkBOhekYq6GYotEjZlMV0hbjEZYvFBowyECMVA5Yc
XpNf5v9u0BjZfYoBaFlVRAGxVUoXhRQhJwgcx7RG/SJaxPC398v1z+A1CmoB+/cp
5ZR5X5BAfIzUFsOrp+ioDexNdtMrO4BWmhbAKuskyzwQC29IEaklrfYPmDFgkl8A
2hfGdrxdOlR1VaRszPjiFhJhmT4h1z3FrD/fFDIjWldKfycPQiPOqY9F2bRMPa+c
/QvihIy7VKx8eoenGqtTwB7C+hIQO4uMouvNFM7Q+/2cwbRLEqWdTr43oyrpuQr3
XWXHKxuL6UxvG/OtF9Gm3KauxIvxyq17AkcranVnQJemBZ1pgdRjTSw72YVFacv4
mMRUJE1oSg8lr/eZcsB08DvoH7Wgf+uMH1uGxOL9OvlJKstTdhWtBQ1D/iHv/sR6
/aEx40fS1pIaOGh3dJL3pmUpm7ODOe8fm/RqyVXRhZryvTDL4Y0vkJhZwuSuqVfO
qbyy1ZHcVy48m9/NxrQbJmphyrRFiHhO0K5vIgmjCkBicnT64mRCALRe0SBnFq7N
8DM7vXNCRkqqVpJOFunR1sBcD8l9JeZGlo8ZiI4TAMMO10PCjgwE6gqoyg4krCtx
QfUxbEpti+3vv8zfh2/IJL0zHPNy6Szp1bhhT754IpMQkLJ73vbk5QGG83qNPsPH
gbBxhB3b4q15Shltg5ic9cuGV38hDH+XVveL/HmokIi9Y9QKEVJpINfHFIsxUNu0
nvGnROfwtsgNi/CRKOXF7V4/kCWAxDAzVwO1yqogJ7iil1y044zX1if60rYWp/SN
O5CNFJYqLWU4sqDE9jCuEu80bB5gAKbzf9/5IxxLctk7+O1GCjYqDcnzK4cmGJJV
xbOeb3UKPoCJtjzApYliasrdZ6jRto5VshKFLfEGTyTWG6QOZ409aRaR7wQPySLV
sQnDzKoa9ARvdQfbND5iHXk1BZ8z+zEURQIbqECJRMcsrWRl3ikItkIFyWSObCpR
havM4WKajhEFQBAzNNl3sIf3AhvRcTOy/2tGgYe6Fvdnm3/Wy/DrU7ARVvIV4ELW
qDK+LeTBEhihLHOWKbxGeC0DVWwlH+ANLHefo59AZjeXOHzt17WLeSUChqjJQnWK
DnCGDHoQ9oZjCUrY5aXXRyJ5NUSBEd94tpctMsvG4jnEjYSSFecYQWi5uP9DuK0n
e5l6K2ct1Ea4L+TDib5yU/MvNGWFUCVDq0YvFZ91lrqeL32J63Ytp9smuzztDooc
SlFL8tMx8Sp8WFYBFxdIk3sV2CDsftvKmp0xuMkxch6Q0YXp3DIpkBz3QrbMJ57N
IXaZa/RcuZDcz0xnkwceC2gFRgytXXXdl5sv3c+d4WqMSQWLqpUtcYeUGXqyKRl2
Mm8hGASlokIVSSW4KEb8VT1jetz4YeTLJC5eSqKsEljCxtvbyPREaQDojGN+7rKb
b4ghoD9Huztit3fwYlLzPc5FBuLIjYEDBHX9fXkwRxIU0knyFkO8BOHg5q6YbAT5
W6NFC/uH8Llyd1L6CyBlBHXvpGYHNW57EFeI+y2dzrz/BAZYOk9NzGLgnsrJNl4u
PHVydtd6IJo6tW1kFaQabuLPdVy9izJnO56NW7t+Eey0kmnlizB7KBdDYPl5inPu
+YlZ3E3YPHRGDLHa5xjXvkuLQf5aXjwc/ppLw6kIvV/n9I3nvFwBCjtqaprEbbfH
OaN02/G3RMKG/sGk++qA28fABzhO0aWJnJDSgAOOVIgtX438Ww6+jfCl1c12+Qjv
pgdZQ8qMEIXF/R10tFrKXT4P2p2HQ/IeLCuc4udUquGazEkmHcmArodeItkFVRO0
W48MH29Ncck8cQb78Ofk+ZTM2ZA3v/mKhGiYiDcXFN73pNvyKiJSJuBG60MU9zRg
LVRzZN/8wt2xdyrradlzU/xHMP1hiGjB/0+llK67mAIbx7eczVLgpPvzOIUE5vv0
NaZgamGx2O+tI4UkemTj73eSVV963iPsDJcztbMW91tIzSGlZvBGBmkwOqq79hao
2+tMbscKelKwsVzUXGyhZuJA8NfvbDD0t/1xeUN2LZs6NUr50pdsZYCOtSbIvn3p
Acb72OLT8eo9pBGUEcVr1PmmCKfWJJGMk3uI5BGT7Qg3G/rrIbeM6dK/0YgkMeHr
N7dzDJpDRTKlKoaArZY1Dh4fctljQwxT68+/B/QUQaZpFwCevDmqWttkn9kSMAys
gvDey4c35wKYzTit6/9EK8AO1QbkkjxydDyu+TqdTTewh5en4fOwkam7QzYQUPyG
BSpfVR23CJB9BV9BR5jm3+HH/yrl0grqrCh/+YQp+n42FHJs/xyBC5w2Gm0SI+Pi
Af0TB8qN9BEDhCAkAvZS0YXNUskIUn9LNLgtOU+GF1g4nrG0H96UlQYcUd9OAmyn
6ANO4Zav94AZZ4O4NivA+f2UizpSw9URKJVBpEgtqBBtjy8w7/swOg96ulSY/ZWp
mqgi9bUxfOFlymNKL9HEUUu77crCIV4fd+STW2R+Hok7HD2KFWu5ttHRauyCCjK2
u1NVTjENG6SxKS/wEXUj9ykKE3XZs5jU+m/fTWkNXGE0ThYVS8ge9QXEAmUxdvoB
N7EEOpTdcqBk1vRIgJzdVGri797QI/OcEI5jl53Sx35JJ6dsawZH0Z2YJK06z1/V
it1Ih2UaYEJJj7jXDMm546tB6C7XwvdGwfEso5P/T6UvQh7C4TbUl8femzbjENoL
ivovFqd/J+gFeMXhh4gStj/JZkN5vkIaQf0LQe4fuHPn3eBVibC+FQk45XY3RD/w
XMwXk9RoC717vVDiA8bXjpJK13ZEH4rOltqOiLBcNnu4QyUUoRNCYLZ0TOiYS+vT
H63SpS6x8hNbIHKhZ/ZAu+eM99Ofelp6ibHw1cgaukSulD6iYl+FTP05HmqNJWr0
DPM1iLdaoDVu1m4kdm44YcRBgrC638n8b7CGjLzj5oG5Gn9EPHZ7TPyyVQU5AazO
EjVZhvzRsXlH8zPEPK/MO4xFsdkXCNaQAfmpz3FyRSSV+Mj2XuMmvhJyNScB2B3V
v1+iyopkQBluTqRkw/UmsyOIcq1PpOJXczldShWkCdL58J85hgBBbxQ5OqUvS2hK
xEtOrVfE0u742Qqwk1jlWky/7PzJp3FDlBHc9kyMNkD5nN7o7cnbwkE7aV0dpq63
ukVXf0dLmlrW29s0mE9eYM0U96SBcoxnTDOX96xZ0wq0uKyITeRwUOp436IbzFPW
ZW4eGYBoYjvZcPBNZPb42EsGFXffQmTAbtGCqBQ77PbLWauyvbAIhwrbP3wYbVYE
GiLq8j94D+TRuFt56W3yw5pam5cGpMHuDENRIOLkH0rD5NxbJEn/pR4ngELG0BAs
IKwY0jBiwdEQKRhzZrbdu7E4M8FoDoKC8z8DJIwo5brTD6YAJod8t2jwq3Y1Z/xw
B/xejIhzTOoFB5AFGoJtLivL63ARVnAdV3MDMeitDJghLoFtlw7TDey/Rcc+WWGO
unOdpwTqHzuiCpuQKYOdlU5UICOhVJgGrKYCZVQlRrvApqL/VTSV2g9tOUDD0ER8
TdmU741cvBC5YgtZzImdTdI/wYn1kTCUzzE8xrPZLbGtUf8PJGRaPBBkfKXKSUYL
ZFx1LhFST1B65MhujaBL5Vju9YeRS868RthRl6AcGSh9g21QnrhN/NUUm/Bjos47
StX8Zv1+NYwV0DD4ahxw8jXcmip0tAZs8f7qT+wV309fB5wdNdcQWutxg8YkkV9F
zZpl1lK3ywTkCsa0GzUrT8//ck73iXOWA38qVXzbISPYVohglgSm/xOodWpDru7b
6tufEPycRczAWbCig08fD39nenQkg9iK4XDBSRXx7XG9YTosMzuu2JH22UHoWd0R
KUzmT6wZCHIY/TWKNxpJCJ4ALUwRt/XtCziRVfqjrXFbZVpUIFJAtKClyxFnxnHf
dv8agXD8ndCw4l5dW2+Z6NmB6/0/oj5vd04XMbd2g8gmroJ5P11ZRM0b2tYvMRuS
3kjPZpvCwxIaFFyXXnBkvNFyTa86aqLIPgWqAFl8BZLCJJ2ki9bIM9iJphio82Lf
vMoJC51kzIz+Yh8gDxRCjDfWVQinuSXAb+tzNRIzNbjOuof6ea8s+t+bDb/nBA70
kNxAKP6N7EujhI0Y8chDljZyAvGIOG1PiPwboz1dTaGvvlrybUlhgxSPvBouM3KQ
iLn22ZGHdKcn4FeR9oAtWJRvxVFbpRuh3bgQnEBc9JjitQhdoJMOr6FaiJ2w4zjE
tt1LNexNFwsEQ4wnwAAcRiqHBJ/mra+NuYPPJb2BRGRkxOtmldd2W+Ny9hKmdNyT
5Qap4GQFkz20Ri8toB/y16Xy3XSuWuR8KrFuEkwC/bapcZgx5tXfvJbXalvc245F
Pe1TB2KppZLGlKXkvNRNSTknm3Me+hERyLkldN4gM03jrX3CUH3JrM0kBHkFaeNe
CHOSDDgMCHNKLgevEtFb62KHQdKQBpq6iD9GLtkGMA5WnO4JwvBJWhEho3t5cVo5
KcRSzKh9KnEt1l/Fz6v9Y05E91oOuKF56JkNJwSEMq53w1EJONxfAToDEKVFpxz8
N2cFRI/5xZ/lZou6zuDegoxHIohZTO/xmOT6akcB8vVuIyoE7XbfT9YDDAZAaYQ8
awzxnGzHpccpSF8evboCWp9as69Nb9HS7dc5DXfX+embgxpEL2w6u7j1UtC0ZsG+
r6Fqq/2rO2acMpSG+A1CSFjkmSnuulMf4ebHcblcgCc101OWrVISoy+8N+ubaatW
i0XUQJWdfOR8g20WoD8QO8nd8/C7X58HrV5qqDHs1r8gXB73pb3EXRU0lXkZjAma
8WwDkqb10z/Jeeg2rsGRbejT9X9PmM+IkkTRoq1BtkWh8vxuKyk7izzF/LhQ1cuO
4nRhraa+M2OEehghXxWdzV9RIo+zhuLLLllKvs7QWz3qm1gnlbXC+NVp/hsWLvk9
/U2u6enwmi9JrA/Wb7u7ZoE9fs2MvjAimQgP3YDrZIa2TTArf5XQYcCF8lFkIenT
bdcwLm0BlI0TPn/yke4xd0BBy9UnRJlYtYeMDe2No9oRzn0Pb5suIignBsMDSQCe
rvZHPSLUY8CZnU0+JFBzXI+/4Cq4OtkgDEvJ0wWZMrRxTlnYFZWL9VxlFHyA2Y4h
Im1S852dm4z5q87M4ruUqzVfaZEZyMc3kRmKRGm9m1uMjPZRdiNEwNPaH/0ePQ+4
4Rc5fTFgStNhyrm6Y9mL6abhpQMc34kUNmh6dATRouQ77+5VShPvwVRtJzAwTDcz
C3C57PgwFlt6ktmqkM/HYrRso/u/ZxBsNZtugriv6sMNPIxPQLsIYvtJK++YrssM
/vaoOFuvXPlnFphKvQFMj+cJUv5/oQuWyFCbZ0G81GohcDaCTo078At5v4Ci0USi
EEw0VYkaX89FYKAbbo0Ie+Hh0Zyg64IsYpujwN2lrn4K1lwmrz/kwG6osF4jsPF4
U/3oFwloqp29wAZd5OHZctFHloSWH3hzeJ6slgrVBZn0b2P6A08kd6qH3PxXGIzw
k+E+5yaJ4KJla8ge3CVdPiuU8JGJb5PS0tH50irwLn53Ji4Fh/i7wsvE0ruu43hj
oOQ6VXYT8bP3Eqlhz5A979w3+3laxkrNkrKa+vPJHtcWNEJrFfvQSkb0DzSeRyDv
Z99nJW3Iwf51M2CkCV/HjtlmmyjY/tOZNS/LB9ZR8Wl9CjqLkzS9WyVdhPkbKegw
m6rmTiZMADCA9w3kTK7nqlVL3wn9RS9RvwvHMIn/KvesddrpnSEaU4JfNpbeaykS
zHqEDLDIA6KeQqfBC/Fvi47USuGonLx4swJ50aWYlSmJ8xhahgd6tvbF5l2/XXKY
2VdU29df+0WHH00ydi2NqGr/WfZ6o5G5vbTYmvx4O0dQxl88izQyM3rUIQKMDhsQ
lrRF1mmojVk1RjzVjb9/Wk3tMBcAsmOJMKKv3ZZdg97XaPu9NXqGVLj3ptxpFvlQ
WhpqxvZkLoqAOeuyVniBDgJ/DsONIi258Im9Ma3FmvWA/uaZOnhdWgN0wjXCEntf
lOGnv7KpwHgX4/QQE53dcZA810AQyCV/YPzJefIIJs2nCJN8Zrzm2GivZrOW06hQ
Xm86eT6zB2xR/mTzsBmem1UgweMd1N1o4Xo5kAn9QaPvsWrx5IF4Anz9z8xknhfS
lo+hgr2+9h2CUvY0aZbKuQ30XvnsZkDUcL4nhuQAqLIvZhg/GLNYkqR22I4f5egT
W40M0B4ONrD9alBbtVOskgYXyNtkB49Yv2ot8oud4cnUVfotOsGUKnrMM9z0TNfs
fkB9xQuRLWZRpnikSr/+EdMxwQuQMrNPptMckUom0cYpRNmv4IL/byG62u0gbrB2
3JB+Or9mG79Jk0ADa5lgfn/wdVRY01Un5UgfFmxVs5CUwtCKvGNsQ6wmvN8DdjTd
6pDQa7GW0/GTwdySIP4ndsX6wGVOoMBK15JPxyZSQrPsPQj/dx1xSnFKAhPujGFG
hkj35668XLxmzdyKwbUz8MKGDcwbPCNoRbBm+sbdDaMKLLVE+RHqri/NuueXJ7rp
+jNI0HAEBpT7ZECPNBmgaf59/18BXCMsWqTwMpkR41ITuRwAEVh669mibDFIJQK9
G6/FiLRrkqesQf2PI0FW5aeXWINiLChqZkbgijWhIc9dk4Xo4xzGoDQz7Es0tn+I
JTSczvXubAtSwo1rldLjpPb+nln2VLpS179PMxu49MU4TIURDr1tKps/zSCgCPIU
uxZ/7tB11jTmxfKQMmJOczUksIe9GCA72C3aqJRXxrF+KvbKbjLehJ5AoLJF8b1e
dIwmOMjDBa6qrYRAKdiOrFT14/gbIlEQhCENyUVEE53FTR/8PgDS7Vf+WPWZKk74
mjnqHsBRgoTv0AsvET3+0omgFwUZ93CeafrmvAgqk1wXQjCvNudkDAK5Sl8e9BkY
zOQ4ryqE3y4PWfGqCNrKavvV3TbWqvPsJJGrFnqa40N/Y/32spjo8Hpz4Qr0hmai
CmJCP8JsElYCBWBkDbqWU+hBlRMXoPnzL/hnFrt+5R7xcii8jpAkt+Hh6dsaivnS
DiMLPmvPLn4cAUs9iMWDhxs+f7AGHbOlgA7KCX1FHI7DMkZIJWPmJP7Mg9NdzjDA
G+VhrgTfieEWiQ9HeQhS+mcB09nbqvFNRiGstiyBanfsGiHkSx3lmMI5ZYrTE0N1
WEVFCxo9t5q7J1M3E593ngADBwVm2+sRqoeybg1a69PGIf3AP4IV6FnP1FriXzMm
sIjk5TVhAiZd6sUfoscFvAkipSmSn/UQiNrLTN/+6yCJhNNu7KYPOB2JSfoVd0Aq
aWhW27J8FETqPhrZjd3l8sLAulznloDVsM83DuzEOmp0MqvAdV9e+TjIe3ifvy+u
Q6I03X5ljez5Hp33aNEnujFxZvOutwP/jJ4/XnDnAmKGZISeBfRWCoD0vbk3so1K
R2At+Jvf2WHw+h8uVXsZ8NfaVlzzHMzT6mTkWKiTLMxaevO/xgvrzXHORut+ZfUE
Y3e9c72Bz+eOgIZulUE94VxeJjh17Yd9FlzZdC3Ctnq2oO3+7yxcf4oew++vl5Ad
bJPQAeQFO7kypfl/1yPEfI6zBIVHkkpjoax9zhJHq+DUTNH+3x9pEYRY4x86rkKR
VOSgr61rLAryF2gf1rjVqUiyDX26ml+pZSfo2NEpffo91G0u3KQ+zkdFL1090vKS
uAutuQOdtpK/k7U9c4sIgC9GHXF099d/8Y1IsnVK4uXNyLw5g5H11NFgyhNTsSyY
hhLS8qBgf2cKORwvOy8wU+hJYu8N8l6+1LQ2iq1G5FrMb9EuDa2w1chTOfvqVieA
mBb85MDYLUM41sKbd1rGyI4SWJ28gpjpNzk2sB60ejy0acraqj39poDxdxnen6Lu
oMd2SRFkhsdcFruUfjX1ihhwSwgBZcP0lVkTbkl71mJrYPbHwmb5zt31DnR76k9+
5lyAEdn0Vhb0w6Dne5VkKgkSbxmguOeZauvCh4wjk6n2r4iHCKeNLmntT+5kUIHn
T5vlRc1EU2sZfsvDVV09P6K8QNev1+QhFkms1NZP/DQW24dcpXCmmBuqY5e1kS8z
ZYRZ8gSC1aglKxHAykHfOvY6LplDC1lpMbLgCX+GueDskAfu0piqLNRu+NedXlHT
Ffq5sJUwpMnskBH7cJ36ud9gci71S+PI77zh4esyyUTlDRTCFhQXdTmp3g4gdedN
ReU1ZnDGPEfy5Z/UsKfhutaXp5KHQzv6mX5Gr4XgqCfzLqxdmOF/qsaVstuJBF2v
ICTaNcv4zxGYHTVd0QqlCfwZHD0XgIKp6crbtCO8s1xdpiIY4dFypnbsCPsLwa4P
aICSPkK1WO5NlynpjoQXofWp/YjI7HyrZoHOXKMQiP5E9qAWA22ET84Cn/KnemXV
a/A08+wOYcmdLmBq1xHSLRGFvZ1VOMoVLySQM6T9pKnkrIiPmnxDlf0Dho58nnIC
Hegjw2wRuqpkdDF7YTjOOiJLz1F1IsLeCvb55U379EOh7xmTkCBGFhcZ+IxepWz3
z0aomZXetfdKXLMsDWW6LGZZiGBTaBFdBP6B/e4xA/qq5ajorZrvwWxGlZSo+Hke
rX3HCCFsnsPtH4gDsCFse3y1E0JHWi2iEe/hlxeK6p6McoY4JWtfw63RuAduE3Zu
xpMgcLmJp1rfXeKAFBJ3b0tJmrAfrJYCOxZUQtVjhG9II8ANSIR2+IY5t2CNiiwj
CDllHQdufZv69KyHCCZQSj/nrmgLOOYHhfqe92rAv/PguekliEQUvENUMF5f8GO1
9FmgFBlmMxygZN+4H/zAYa/KYrKOFEEJnzCQMj8pVg73aW7ZBbcDwTXd4HWH0BOF
JlmMH+BMW6cR09AwD++Aou7Q5HLsA+f0dn1BdE0hoy5fCd2eksHHssNTADbQFpSp
jxgO/IWZD1eO5hML3uK0OT4X3uNR3+xvMY4geKeXU/kqtBmMuXc4nqdQMegLwO2I
rKqnjQVhl73N+3NB9t7G2Wist+mb3MTuWzwO4O3FvokdiZktnJaup2q0MNrkYrbf
M5hXZuYzgtIdB5Cfp9h3Ns5+mjZXcgAG3qOkOnWEtk2BfC/BuHJ74Gtn1gby+Srj
fHHx+KG/OKt/U13o4mgsmTk2OXPzHZR2OpLwHJJqCswMy0SBHbXdRQEYZbVqQsX4
+mAWGhpHQC59Lxg9emI4uI2XSURW/42BOFiHrajXJQou1Cirg1rRmljAnDkthNwd
+cMgaFda5iDq8XHEFQy05nLOtNka3MG4eXz0yA5NPT6LHx7uJap7XdMAjZMWEODb
PlbA+LnxwagA2YQWyjyLLyQ6r0a/+eLnt26MHihu4hAuPVZvY9lpp/J8Ui02NR2z
30+q0TjAOwwC+KWWsrZ99P9Nhi35Buw9ofsoNVhqrfY7zsdxCk+RmEznIPo4Sr4H
2kaqttIlPe+P3b7rEwS7/OgLGwAz/8tg3Ns8AdLcXmXibfBWh4LyGLtaaJSO/xoT
b3O4sWkvEVxc5k0TtA3vueSBY+ljs6swS3REgNv4bUV4OotWFqG5paM4dOI9qoWh
bJ8B7H2TZXNyuz0w+oehnqCYVTgy9r0xbIfuyqcf3+c+Sd8jeiz9wga2Rx3Nuey7
0oeefdHafmiX26fiiRLkaksb7ggq06vGZAiWwW7KT2MyudZ8u5zvolr2trZblZ6J
WaceR8QXHCwQcHuCTlLo1FygmKT/FvTjCKhzEOTggUn89olPBuroVOwlt9sA5I8R
1NE0LnHv/vz7K/L2wthP5vBTx6hbT2LzRsUWghlu61FXfvEpRnEc4qG8F/MO9zHG
p+5n4MR7jXI4bOtvCkIfmP440zwEioqC+jqq0KSmiRYkPiAMHxRPBx9RB2rSrva3
RuC8DfTMqMeF6B8G0T+u4/+X42zh/zmmwtyByymPTQryJ4F+XSuVumGaqEqjqMVA
YGp90jN3421A8UCOJte3bgl8XfOxMi0we0GNW9HocA2bLuhy5z/wnvwWtv0AmkYO
C+7y4t8ItvGcNiA3TFzTBHtyvqR8yZf5tlHyzlmagqq51giPFlRPJZReeM8eL3bN
LBa1KXkGPHdMjvhh/9NwHZT7BApxfUsqEwKqQFFMQrBsOyapZL/p0R3KBzBrzY4N
qNH+6ATnVpvATk9M+3qHKQ/ILnDhReRxA29o9sZxagjA8Qk5RC4y5F3oNgRqaGXm
X7L9KBzkJkPRF32scK/aYPed3P3gPmewn5pr5pK//3QhE9KR0bE08oCmnGLT5dYH
eQ0TwcDtzo+55QGHORKCw0bAY4QJ4aBbV/6Fm/RR2vEt89ckCgogKhEIuv5M28Ft
dSZqnT4Zs8aS+quQ09rd2jN/SyaJ2eH96BFK6szHt9DsB0hv5SZv5g5HxAQZN4vL
kiqSo9bQE5uyANLZb06mSxSgMhdsNIiAP0ylTJMoZlqeRKQ+ZSBszACGQovVdkkd
R50n/fXjjT9W1AoVKXcSk5NYYLrC+dBPP1heuLLX9r56OieEcewsnrjA66ua9pUO
rRRofAIm/CNoCyilGVU8GjyTl1kD6oQkF64ZZEICZy4CZeyowiG3GvVafoRCra+R
3bz+lrN7gQ+nrObROAQFdwqlry0sDEdiOFo+8hAWtoQABYvxEqnow5n8z+1CH3lD
z20csePoMX4w1h1snT/IAZyp5ugzh75elWOXk/h/XZXJyiCKg+XU6MzMtWBAilM/
SEIaa9X+mWP9rzgtAVUWFJO+Jwl0muOYvwHDgnl80b9OXKLrmS1p3ueHoLsT/wkz
+VIDCCN5vVMy6LF6RM9lvb8sZYg4qv89mHAECLb/4RpEmb726zvTU0EC8IcNVnVH
xfuMjjzJCK7jxk5IPxNIRe/RBaNlI3JoEr0EgM1bVKojBYIt/iV8cfBTsrhJyFcf
fAL7lagrKPqOi4n+aggQOJT/kBgLEp1zJY+C9dD7Dzj+tBd04jxN4Z+N9axkT/7z
oQ8cCQhu7kl87cRqwoNcvDroE0gmX8X4iNiKKAj4YldH8jp6BFi8LYnxRTE0S2fM
jAPkadyq0/iooPIeoj2sij7DadJMzoCCBr7Vhhm3G4vmx/+NTabyq6o9zUdZkHwN
13xJsWUX5gb5zn+2+713IU0A9T5mNai4p/E5wXEZBGFweKylE+sFVIu/aSEhbKAX
9xtBcg3EV4zNgZfnZi7z3bQdCsd3Trd8HoI7FSENQcq1CEM5/sgiWCu+wtwGlB+T
wOtaJY0PUVWMuegvqljf3Yvya+Z+/Vj/JO5svM0hSU5igS3tpGBCLrW3g1cP54MV
Wllqq+07fiaOz9zqyWPSLuBZSGc5vCACsUok1UNVfgPYhBghLkq3LMzetgB9xoCv
md9+jdWhqyVr02s70ak+O+NusefIJ5Zpv/yOFK+raPZUZGwcWomKOPuwGvD0zURI
GA8tpnmOZHnpu43gwCX8x2JK9UNL/8TjaXuK2pfFIhWZ1OQmEyKPyt9fk/d0gncV
7gsGUblO+5qqLtzw7UKLQOXseeNuAst9kxfipF0nKha5lQDE4I4naMhwlzD9xQXx
OK+NS4hT0JeVQYy+KmtRvHPBaXyvzL7aopIdYHvjqwzZnX65qkpZhJyFJb9KGC9f
2rajo9a1yVLqVzCvpjJ9fFq4QmbwR9mKZab+hb/cHwUA5Fc8hfXwFuwEHElZuzVo
5xOHBE5Q9Pqn9xoG5CILPWt3mbrW7w39z8DInmFbInfuWO6YbMnp2CrbHnrkTXbY
eOhaOvy9HGOvg3Xvn2P9u+bQnfRSWltkQee6w4MbG3LEoASdEI+rSvrCdhv95dX+
Ze1pI+UsiU8EgvSGq2LaS0U69fAwTmvX0LC3GrIz0ktdLQ/fHHPdgcM4g6sVEk06
5uPlXaZVA0t4L2WxLI4JKojwUPLg6I/9bdGiNp9dfFZpPUy8gDhUZaX7f3JyU10d
EEwxrYYCeXBXHHbuHhEIJOpt1baYHYs/T9lbQvQngSFxPuATopscJiCTl+tgMEis
Htx43+gpo3I4ZHrvyBiQRlPbudZwvfXfx0a72hwvfeOYZHvwDba6f7sRVrAnt5FZ
LrGJaJtKFAlsgDw+kRFBWV7Fas+ANu0JorC4R7MpNYxTFBmsAca1z9faTuXXTb+O
TDoRHjajWj9Z6HpS5xOFRkXxSElFzEAq3Qh9WEcbNO+BnSPCiKPEn8hjIDY5aq78
NV/S4o7ify2G+hvmSiVql6t6jLzoaTtNSMSV8nhH5LgdeA8kufZsW9UXZu1AGEje
HQwHWIeDQxUq75VYgq+A3e4g7IkmZXLp85dQDBEcTX4BYMnLgpkzKWMKDPco/f/x
96CXPvjoHPOc5Ue5ySVBlCKZut1KYAimAe0CD+1J/S431Hktp9UcYLAa4Azhqyt+
+CG47+YJiwAw2PKSGrB2awCucHG5uq5oNEt1bjEA0c/5hDA3/g8qhqzllD6S7Auv
98DfgRL7ubFi256P8L1RBwYwxsMxrCe2+JlOXWc3hO734YFEG+PTZlG4xoZ1nkVr
01xBWWETF2bncDa2OQ51g5fE6ZUDZPxgLAvcnFGqUraIBfZhHiQSX6xOE2kOL/dd
+1cZsLcFAhteTfKvirZerz/eQbwh3C6X4xifejxc8knOl1EXhJkdAZPCiroB4108
QzzNH5UIzrCj5cpfB0+z7MTVqyicQga3O8UgLCsWiaEK1EU0M7jVnqXyWF3+2Lt2
9VhpWgIQT4gYrbHsK+p0N8tQ3hHwrIRgptG7KbUNfjzjWGDwy2AY3Ocdkg1nRZAI
xlszJKu8X/gBdDhfDhj9WLumY3f3v+L4DDZ5CPhaeG26CCmIAkQxcqBCYKGa6BMK
6rDYr+7ZYLKq49zzFqEgNbCf6xou+kbT3p7ORK/c/npnsdksW9sTSWXQRfaOEEw+
IQ6qD0qI1zOWJz5zhavSxhkyZnwvcFqddnNuhH/zgpkF/NnK+PF+hu4hG6+BJXOA
SkJtF95HJDKf95GU4K20OjIH9CtwwG3xjVVK1bkaUOw75dL6xvSS11iz2Hvr/eys
5dnwXzaI5FpSbJ1DQmlEOLhxSOWcTFP0HFa7wU2fBx+0UoGu9VyDVu7yIXupGQG2
JkVbz5rP3wsYw0So6bzyYjCOAEZu+sbbDBE6qMp0FxVq+ocUClMGRXwvcn+SKUoJ
Xc2TYpYQaQtDw7T2BCmarV6xyAuxr4VKPD3j9zYaCk9oIWBSxdL4VOPwivDM7GPN
KypuqPisf+Rrle+PAT9K8LJy459UIVDiGg6NZ/1rE9aCVJ7q7WFtkA/53z3qNOQo
GJFFQbKmD+om7DYz/O5Cy5CLghbV+RUM6dGSAlJZndsRx0S3zPPkg6MegzZXJvCl
TujQtnnob7cYGkeYTGe6BVb5DH9h6fKaUuwSkoBHp7ufaoaUkDfkfMijAdmCfQb6
XllZ+AkqTAvebwAPCNB9iXmTXeJ15Z4kgJjuPkaJo6BL0M/B9z5KEqbZyOC1a25p
Oay3qcY/w0qUGxbfs1DNcFV6Wb9ZTwxxWginB5H1FWofQoKs6y30Nl6xwxeRRimb
pThml0fWyGNUn13RVernk5iFq6fuimZrUU3rNqJ+T56hxaj7LpF2Y0XXBHzryWac
5kVADlgrLc8PAvYBfoa3YvO9NHgQgtnXqRBbH6c/RoI3MsfDW4eSAV+nFsj8p/RZ
oXRhclEunDzL4EWat35qGi1VQ0CfL8TeQtDa2j0ugKe4fpR6elEVrblQ0DoU409O
6mPthmWY59M0EGFQAEciKvrhetExanvSQuxTf4oibTiqn1Rw1K8k1RpGALcLjj8x
0TMz27EcILNkQ2RgaesYgkognQZ0OEbf1T5Y+/OkCCSZMRV6JCwgLYTWuFNDaUgA
5foV/aLoke/HPk9smtkSky92eC6LbZzoOH/axbBdL75uFyqpE2MUl08b8IGJ7/3F
/hXaiaNObNPHdJ/C4lhZxa93TU5e/WWhPFalQXIjxQ8DoS2BIxWyqiLA9VBgyeGA
1s8jNiWH8TzhfDPrACay5IOr21PsoTstM1kXkGGs9DzvJRzamNt+fH8lEqIWN5fe
RDf7RBq1C1AlpH9Nk+U0IbX06OsCs4xfAaS2S2g6g2YdGxRE7BDfhLj7nRPyqSFF
qjWRkZWxin3hymR5PXxPVHeb2jz2BII6ULrSeXDmZOFUdPn2x37kq33xcJPXG7PI
piE2STn4JZ0bITPaKY8d8HIp5M5uhSLejr5bRafOAoa5Do9JjlD3mRQsINUbbcWb
XQRPa22hYof3e5j0+NtnW/I6bcAgW4jNSBAegUne+fc2qqY3BlEnmU5k3Z1XEYDG
gL2VGgxBcnEyLjmetXYsiQPPjgEJh/++qZ3wkUALoNR/pqTee1QGl9pGEs7Tn0G6
wykhHR+7MyYnj0fLevNVoEMRmmXrNBWmpN5LHswk/YtBEfuWCqjVgrRYv9gSpvp6
oAWCdBAjrxxgJYguBW96jBc0QtHAvP7ztbPTAFsKV/LmPvUySQhexeMsdnho3md0
k213ZVaXUHCvyesj+8UcaZmEE/wGF4Yrs2oeBYYga11MFVSVcpA3L87E7EDVc6mP
oN6m5LXtVpXU2eQCZlgLaffqNulWvM+BGIIleefLmGvmJFsJAg1+imDMm3eDUPyr
8jq3nJUzkoCsb4FO8X2cigz3IVcGdbCc/JF6chmw3Kpaj2XbqB4Q0cDgOgcSeVl7
i00ENgsf2wdZwFQxTa+17CE3R+wbOCHZmDzjIMuynbxJCfc65gjxMpVMr10aA3n9
w6bnndFi+nXtOIdpFGm75s5hC9i2gVm3nK4sG7cfBFJ7u5Yp70z1t3KRrqTS/kSz
clcCNi9POBacow2QKO3Fnz8mNqhA72LVKvpur5YaEtIJjjalzSaEQx+HW3G3vZPG
fX+yCvmtIDIFjACmVcwVUftRJnsnU9dLI3Hu1ZJHoq4uN4yHtW8GXQYLd4HDQquj
FE57EZIFiX0lnOLyLcc3PToS2cCkOGbEd0ZKJiRb4TzE+mqUng6C1SsFVoB9eP7z
dqaFMWY4ukW3ZN9rXV41ON4fh/kDVLxWBjChUp5K0rihgW9F/MsTFmxaLr1LsTlz
gImezF7GAjH17FfYNnAqruWHIGuCfLDnyyQE+ulObbAMMpycX3jqJWUIa38jGQE9
lRKckiamY35mH9jCUFU5J5OFEw9xNttxLqVH6SEBYAwrfOI+iApdctp3UfGmuA8N
Xu+CBlwKOkO49wSHo598IoF4oyhxrJOAA2yZMtJZ18xK09/WkC5FMkPQPo8NM2Gr
9PWCpF1NehIEIWjKsEHzNXOCfVUKjKphlchTSe5kPyEkU39H8HiFS90Vx8OrYbdN
8jeW6x3Ul5/mZOzzk8mQZwxuWWtDWrA8rP9kKPZEuWfo/SI9GsAE7Y09w9JtsD80
L+3P5B85jfOdapmwvLbnS7ZVbOSn3DXIIt8ycSe3ZSlnRFXLWZnVZl6b9JuTA5la
fPb4efHwgUH61NUjmMO0qaHNJl7mBUsPFPTh+cB3Aj2skKOcsMxSQMLY+tLSYDwt
JyjFTrLinJYCECj8naPTYQuxNTvq+AoIkJKjiVZfooJPriiB3UFjzL1awGCM3maP
IiKcLIDjy+9rkN4QMKDCKSIRxbu6hi+1I//R3vj4+8hD91+ptgzsiaGctYulr0MQ
mLSqYuqs7OUtRrc320FaoQ8XUCvZgyiU7lhnnggUc+rjETS4uZkOwGSxnNVi55kI
OPXozz75j8ZtDZKHHBk0ifNbWTQRFEw39eE0QoC2xnWwVptfWWQDitOrh1zgn1Ib
735VCWPBbfRX4EiUW9MRh9JoZy2yPWH4XX78lt/t5cXXVZNDqxdiUrcmrbvw/oVV
5ocodEf/qK8L51eBuuvvxauiYk4qq7HFsjJUwGUpj03rN5un3tLWNzOHUhDAXwmD
ih5WWW3iA+9WfUhgWDnbA0ghXBjwl5q2xF40PAGRyJ2/P4jYpJPku46YtQdlRCcK
YcoJZ4uTtqOGH87olRdfhuo7fEve7MRVGBrA9qNzzwJxfUQq+zj5Xjvg4SnABjEH
0PsJPp2HNd13Ygaw17vQCWdC1sUEtDDhtYdbbNZwjgjmHhquV5efAeGSN0BlCMdS
19idBm/+tBoGmBw1q8IfnJ9QDWO+/tLtr3CHT5ViRHOFxDJftzuHK4l1VmgY2fXV
+2BlCBciPXj8nBRQ0jMBaDWWSiKWVXeqBJwwKJivZQfEf+nfKLOrkzXfeZ3WrvtS
xUToHhtI+WProbDDrlUBoCnDakGpQBhVxAXRXHtRJJCmtdi7STGKsjl2vsUOHGv0
a80rN0i0unfpOjB3De9/YI4maTzmLNCTdRm+U7ICsJ3CLJiEVwCn5iGxfXNPvU2z
+4K95R0PFqojpfuoYUZUTAmBWhz3ZgzDJQset3ttjdFVYN7zft3CGbfQbn0f30bX
G+s2Zx0KCDNPe+Fv3IQtt80Oeq1r9WR2WR5AlstPFK+ONemxON8+SFjHmxgrqyIW
DayqTRBNqVOXcw3LiZgxMCP3if0iJ1m9WLVUNKA6fp5Ow4dr2WzTXduuFHl0NJIJ
fgRNFlCEhCY7LJcnDXWw+t4tChkkLQt9bkPbIYwcBLEnIlc4HyUgxgjkg1beepPN
bRG/c5Rs/DGeeuo0J14cks4BAGFai2qnKs45svC1HsRdiaJx6IsvTafiCwwdm7K3
qyCKy0TnmSx50UVPk5tzyoInt/pslYnQUIwmlZQN9SlqGxxPrrhN3D/D2GCrKnlj
25WtqW9cs/Nr+gjt7A8B/DluS92HIW1oDBJQq3KMjmXfgDG+VDGnJRK8mVgoFwUC
nJD/xsGwbWmgkGzEW5a5zxzYH3I4vLGerHBD0/ndYdanWEcgpyan9JLMwzGMH/Hj
UUVxVT9TJdOZ15lLP4e3WPr3TKrOHwh1v62Z87StF34yOm/afwRbeIwJYw6oSlct
KZb4VO6TVvL2ouNuL5VbBXuMorPfbyiVK4JgKoGHvcE5EcPFiLrsOhA7wObCAwpP
G3jz5Sc7TZ5Q060v0bhCd3mXQ42fJbUj77nQYI7JZrY3bm13QKlNfvasEzuDJR42
nTsku0C9OG3r6HwSmVYp1o5oNgmguLynBApqZfVgzbD4iO12WUBvIU2BEjPu1We1
/eH66g3rOvUNNdJeAVbLwl0ZE+mZFyM+ht00DSnkuusQjWbSkDuRhW+3oeHTDl8A
wlqL/NR2NpOEYrfDZytJMGAX7CZ4bLVSK/RmCNllVoI6bO1Yap6YGPZm2to75K3L
zY7DivG4XLcJzcj5NkzQzJ/emj4k4SNo16RM5NF5H3vywcbQJiGZQ2SwPTlpLGgt
KDJSGXOOJraQ35KXNPj/9XofOScD/Trqc6V9UaOEwp7Ur0iwxsbUIMJbL18e64m0
9K9mpBmZFObjUeqPv0ljJ2gBsyqdiUEXO+bxLBXWVOd0WLOkL4bSxbpEvVzjvBvw
2er5FP+zs5TuTm/5ju5yHpV+p+gsgenQf+8+XvtYOoJPYvKPzzCw9rEG88eDeNSh
zXURVDrQFxhnNn6fXHhIQ3FnMvQahbELTtHIkiqT9Hl7H4H/H3aVBKVF69yA1isL
ZkERHMf/NUuFAOhO5j8YFub4ILONeW9wxE/bqNoV8VFQOjVJSR+KgIz6SgQ7e4MO
EGHxa0uRFWd25T87sMcDb/4q0xSXvj5JkmFPW6Muj/CtR5s/b+jpHSr8NyDEWzC2
5OiohlT9/b/5M51phcgLKJwHXERGWDvOi9dv8d4zQ4F1x0OodduYqvsTeOuHBbMz
91+R9hhGTree6YQABCGASMFGbiriRmLoMTq/OTnYnSeyR6BzlX6IlAzJDadpBfW5
Keo5IzM3wW9g3+KXpSTwkT+m0qa1VGfwJ58enqtEb9HRrMr3WsWLtrkVROFs2uOO
ZQUzA96eq7XeruV2xh3dlzrsCCtFBrnIrB4dTVz41+MPq3KaSwiia9HTlNsimA+M
yEtNy3H3C9W1aCO/p7Dz+OMKPgZ/CyZklRHSp0SmAx1ujvmLqiRTqXX0ksq56jvj
PQLRS83V2BE7KxGIv8zPE/1c+sLQF/Io+baOh3iXW/0GQYRdPZLjXdWV7MhALADQ
Sd17bkzhH8yoB6qA9HzXCGlyztbR1dYj2jP6STyZUna/Sv/MU4thCPPumgGnHCMQ
0RZi2DD4L5smi+RUYq7vqSiDhV2OQtcOCy+HkSAYLdUC4acNrTTlz3cYRhNB/1n+
dJ/Gm2wX1AUJltPua5V5CIEzkS71RkjY0/dktkOkvtUKmIMLLp9/Ermgiu00RwV8
oWyQvxJtIIHhK7+vmAgg7/F1l1KPdriwxM5q/x/mVfUnHh7XQM66afxgUG09hNfu
32ZCaTfByfZhW3sFS4sXyYEZN6J5v9HWUWfEpJOJ6I3P3gkLyjFyxt/BxX4Kpapm
cTG3sD4cfWzbGDLaAC0ZrPRb2vKGk54My+nGY/YAZwIeZsldK5HeDh/q4rf7QRji
iQfuMGGzRumKl3s77gIAElVr5cS2Gy9dGCLIWabZLQDUmlgrO+TppjG1BE05LHm9
+wAmxM9yXclrMy0tog+LUAM8MU/vHtyE+rrFtKSt6ts1xEeF9WWcyh+ZX3XPSOPL
CEegRmwsPoUhjb6PwBSxB2Uzwyb9xKdbkgkDswB0iKPDsmD5E/kUIw4oU7FfCb2d
BsBq+t/ya2jwkDLm2iC2H+OLAET2hZSx+6jcisq0wNTrmn8eUBLH5dbpMtwLUUM8
M8WueHSsyNAXRHzvuKds5Ed2nBP3Ik7wPAoFqTZHMhdi0NwYCYzYGqwNdK0ai+A6
q6e4699+tXBfvh8nN1JB21ZdubPrqdAqXhBO/fqkMXWECEMSWUUs9Y2BthfjEfkX
Blmow0pa+GeQDD/60ZWmszd7ipYEyTrAwRNKBEjKUzntAlOc1bks0FA3EzxtMm9h
82YqkGKVzLLmupqIkpQ/8ToFBQesyVtA2ZKVnnkp8gTPSQgPUQuSYheEVPNYDLKe
iYyBSvji670TIHWz0pzGhdpMi2loEY+ilk3HCsyJ3N951npH1+cVBZU87n92F+vz
gzOH2ZIyGIPjcA04ErYuXzDUlnbeWhwm7RYx2GyeAXIHBtusmTBo4utm0BEE6vuw
u5dE2LukeXD8JTxFM11rzkd54uqFKSAuc+dnPM54zLGNLPTjcsw48AE4DPcfajfV
I3y6uLqA3SeEEAK8wE8Zhe/H9nZZpn40IxmU7S9vCVGDulOKi09LMjXiDVA9MGoV
BOlDWX1WKALM2S2/0R06ztUSvrEz1uMCRTItqPt977KOHjoxOUoSJM7SOWCvz5Ew
iAfjOGMFoiU1o4XGCB1sAND1Nb0E1Px8+MPwQ/OKma8pKq/1GVE6VSh6V70iN1vb
J6ZdBEX44zKvTi0m8ksScgwcYfOAQkRQSdYwhm81IHbRIyHVhVSRcqXFkw+O6P2a
E2cD+b1gUcVFElGbWmNxbWLKqNUaM1TpyEGnaI+JBFOgIw4FkuuOsJPq7RUbW2PC
3jrAPWpWDU7+B39s+g1J0TLLhGlkI9SLp7sJwaQ0OICJpajTYe2hjxttsK32lKyx
SVhtM2ybTRCgpXo+dgdkGigJzi6blJkNSAX7XQek7gHsGSQv2Yy9OT0KnF+GnfkX
gbUzsW1Ifp1fiAivfzQ7DJkBGJFAJTRnZQDLkOSKD7QuIL1vIKjQjBHL8cB99NSU
rcigWwt3CgHhAmmrpnC5WWXSF5PsQ3GnmAM0WmC1oIGQkYlXFd7+xjkYkGaP9qUf
ozVmdH2EUl43B9deiN4gynYCH8ME+r60q+wpJuDsnR4fkI7nGSOh3dc7ZRfQ49An
S/XwXSZGzJpoZvPx3N/PhyUbOBmvgz+fNrS3nI2vlhkjussFm6wFCNe5dzjT3Jo+
AKAjylSoRnKEAjBiF+1j3yCC1Ak8F1Jmtk/e98V4vLq5NYXrwNXE4egMWRKKrcDs
kK/UjppXlyzruWAG+EiLYJjl318zszKy54p0YGfR+qxHnfFaCA35L2Hn3sVVtzJJ
u5JMRhrTixkBpYzKadfYcRlFnQQS73Ciw+qzkXcrW+QhWqAycQgZpL3/l9d0BfOh
CXVptNRsbzqRtG6updoGt/yKNFCRTzzLqCmw+bR0511UBpHWGNG8qCIjvxiUwBPw
jBHaHi1uB42tpnrABf7SfDr/JXm8wvbj5udoIVpJnyXrwn38k64QZM0Caaabt8fv
mbCOTUyLDl+/L9oWW7W7rgrN+Ej9RH/FLGNC4UsnU+b/+Llwv6ZmNrLh9NNKDHU1
9Pd5idCMHFvVP45wv/VQYHDf67RAluyXbLQbDEwP7d2/Y8VMCBE65LieRuEPteje
VDsrDkZp2UDmRWUzfOrCP0981saKoc7LCbLQwla03iqi9uDw81Tdo+eZ7m8QVqZD
Y1scJhkPVYiDOThIRBb+EpJwNTEeXBWljvhVFwPbl9oD+WVykB/mWbX74qKJ681g
AG/XzMTJ81AeJfjZu8O5igg9zzC6YoG+o5AmnG1GkOPQ/zNWtFswUj8n8dmVwOtU
jf6qBKCbKElfPaBMiDL1r8iAPyOTjgCuTl8U5Tb0oWbh1gBE9Is1ywzvHMuYUJg1
F9DKO7txAAuBrPfI+c76gMs8cJancfE/ezzK+vusL/tomDhEo3sLiMEBkk+2jr9J
G7GjnXBvQHp26x6isMMG+oo08G4U5WAWN4grR2sD+X88J5QY1q4TQ80g+HudJboo
mhXJm3V9MfDLduHM2FbB9QAiFXCUcZ4WDivLTWv89yq1oJoYYy8U57Aq3Dh2wdgU
+yCuI3zY+5tkgHOJ07G3iw573546pFRRYk1P9r/QiZEaForr7/YxFYP20G2WWM/S
6TATMT1NP7rIiKGHGmqc04yMhhUiqFWUwdS0iFEApFv8CzXeGFUMFKeVx+uTMaMd
LeVlQn4KIY8dEZZ2mVZh2kedwe4iWikmy6FreAX0SD90NwuLuoTfvLoDbAM6yqZw
h8KTJHxhHLVBg8cyLezLjCxMFR3/AgGFtPs8+ymOJgrFQqdWqgPa6U4Uyt/gWtqy
wIRJ5gPaMlBSGg1XvA8DW1/dt5xvjuAqFJ8+ifqZEeNVSpTGIT61pxCc1Q6AWCL1
zC+b1wc7Rm8b03u046lCPMxSu/79GKTBa3wMhSZyl41k3MMPPtaxajgdUaCIqy3e
zOSlEuToszeLR9DNSBs3RQPOV+JlOmqogRGRQQEkei2c417Fv0Ec5Ul7vv+Y0RGy
ywPERJsfDf7Iy8Ok0iNBGsRSZu/NDgyXgGY+A2v4F/ovE7vLutkZ0RXZTwLVF5wA
cxs8To4GuxDY3DUK2ehjjU7TiBwILMl/VuO3fwWSbXwmN18/LzG72nHuxH4y6TC8
MJji6fWrcvoe2CWsgebknOKVQz7AdWtlN4Tusyz5x1RfWt8Mdvn40jUU6WtK6wh4
0HExpGP+0vH42JgqDWehSr/1AkDKLwfor7K+UPaeqtGadFc1JafimcMR4k84X6Xa
g7q6PqKusxXtlerwAExgK95ZDm9l/lHVRqDNEGFvYqqGr2MjdNpK2d+j6EvLBNqd
cAXfs2usCcwvhx4EaRDzBVlW9hgzrMBEtjpBwPY3RIxHQyjeW3+LGn62wuchuzBS
kO+dihghm5xPB2+E8brIoT3QygZHAmlBGqL9fGOs4GLdrwKErSec3jzq8FZsR6rc
L+MMs7rv7cohUnnzGWTjt91THNtm9kU7Th7TZH63vs+yhLIE0AnqtwCkUnYPYRGD
kdJvVXG3p3o2yxe5v/3IDGnH6zu+taV4vr1Ln5mLVy2K3AbliaHRKKXYP59+KEnl
OYUPBXDAiTnr03IEGrGu56ndNaA4q61CQqsw3EhStZ3gmhg+bnIbyc8jZqrWDxcu
UedZ6yqvoNHe1R3nK2ccs2+L2IkpvBqn1kQ8qTLdRR12lU9vKKwHFSe+eWiiL1Au
DJk92o5Vy50RMz8ZQfdoFgXrDbmIYZc5Mz9VqIllyq1LqWhrHshs6oMd2Jjp7Eq+
d/lt5kfj4dDU3HPpWj1RN0y8zFTIfYnj1Wp56ZnBrGF5ovbSlvGSoR18VMkbrkJJ
k+xa5wvYnbnjm7OgtReLI+ZIH5pPvK6w8ekvATHhPrgbUAx5VNmtslF3GdZW59Wa
qfFmAlteFlFUBIH0N8OjOlWDnOvnwKe7VKggdWuicNqkP9zkIblMiNAKJG7W14RN
oQ1hgi32AF6NJP0+CkQoaw5MnnUkJloy2u69PnxXm3mCiRrS9X2psPcsTcnlsKTy
FQH3LxpOHtPdFr5e6vBTJL52TYgQ1Gwp6d4w52jm8MAmXPi0hDKd/B/mCrsFCBHi
ISmwMiknnM+RwIZ20OKy0UchRpBZ0i5N01FaOxgIqCc9oUoDoDEitds7sK7cxll9
JVAVJG1R6O6RMG+YD6d+bW+Yw6DlG/dqmmebjOhlDWuNTG3XLpBaU+VnHYozOybW
ChH4PYtUC2eVm6vO4NwCnYG7RO+NdYucbRGXuFlf0vHd7gZJ1TCrtDG+hZuyrHDH
TjuqCVF05wVtFVDUVBmTZu2HZ+gmdX5WLSQW4PfV8PKptF6JwUXztlEWnNRsxlLZ
SNlaZC5r35sYAL8ZOIr6Xx1zk8IITJsmtXnOf5wwrCeZcJMtk8a3/dm0QsG/9rXl
/bKkHXwR0wm6+wRvxcUwKAixlJvPm+U/8aA0jef/VZDaWgz8WrCLcLMnSReoPqvW
Ky/6ljxV7Rtfi5GuoEYUuWGpLjvFAhNLLXRbPoUCSqiWiGPjcrSEozBzTyj/ehZi
wSJCXdt5w75qgMjvPFrnSGqDfZSsj0S8Q0yHxZYyEkrVqHfu+njiQ0X11H/D5mHG
I08T+k9jA3c/Lv5HaIefhWci5f0BywD4Ooo6i6HLvZp60hdVjyxyYpOWX9RyooJK
XDFZhkYKIHoi+HrCCIdm/oaRwQ6Fhj1y6yWH6yKdEtCJxFkr+fUWrdgjxwkDNJce
P/oU6KvaEXwi3eRAvYeLxejrwTIYsAqL7EbDqhWMSclDxoe3j/HZAZDZB/8c9KCU
3NGrSD1qfqo2uXDCftWifQQ7Ns0T2KgFHYXa+cwVfgauOVfd6LYMVMJDXzvskJhy
g2w/xbEB1Tqh8xuzGxvZdisy17J6o5kpX4H1zy5rxFUG8hqtGkPWtIHKqmNMM8JG
MqDp1lB15YZd/2AmB/Jxjzxr5KE6jxtDATuJlH1nvQf3pzDU9G36JG+OknPUOEjm
P+Un5Z3yCMU1tt6SpJqbtZO2Jh/ZmBJ1UtrpO1/1ZkALKTyapppcgHqBYUYsq9Ed
YPs8/e1Gyg0IawO6vBhQHBiyCvcy6r/E595pit8gX1UZAmI/OPDnKe/5d01wEWpL
ovSynLT16LkfuUYeHfV4F2I5gwPeX6f9Y5C9Xc27uLOhMttFotdDK5SIKZl/8w6u
9cTGZk00nDUynWz4/NcJ2q48dN9cIdKYxMgVYUCE0v8sbDS942tYqVn3cKb4uqu/
1H+nlx3FFTDTHk2PYTRXbYyXphRPNQnPFPJPGB/CDdcaIcwHA7ejkieNbJazI1R0
MdMGCpMlkMkMK+hdir0n7NmeKlsVJ8g0i+U6LmKRJ6SSP4mD3Q+7VOfKaGae5YQR
TRpqf1rYZJ3a5RP26I0qElkOZwtFck0b1EnlnFyR19hdWVHzj4884dVhsFQFRtNl
YVojGG14uhdTZ++XZuAUO2BS3x2aXniVtHzeMTr5K9FeHX5QoqjIJqWIa0+rlI+e
LEmXYZvkvV7IcCgYvtYwCdlvinnITWHqcrB1V0/61+sAhxxK/fhSUNYl4q26hJML
j7zkYA1D7tgfwSN2u2KwawVnAkndGq25899TxH0G4Ktvsy/okXYnFnRsj2woaNR0
AeOHyp3+YUY48mC4pN/DUmQqb34Le69oy69whSLx2y1mhj3aN1F7aPlN/a1DegRg
DUvhePvxJbxYCXvDMa++iDtxfbcmmaCndPoUxoEq/eLtpB4wfc6khueRF1JOCbhA
TalHKdDYrTXzBLJ871z5YPzwEKT00G3crR3E24bwhRLd4SOAeMfw18GUWB3deXki
FsTvUaqBnOVOV9M487lru5HVO/fKQtlxWBay9TXycPu0rtZ1ttr2jcBPzsTiILne
Y256C6ONYkHselvKd4w0Ma8WEAh7lmywmaEE0bhDrScdNdtVck08gu0Olc3TwAFC
Z7r3xV4n1dDcKp1EQn1+m94IT3xIo7zu42yOAfvxL+MziZHyJA9sfxAetT/kgeM7
YtvL2iI3p0647qtKx3SdajbEcpgfmKJdgDXJo2bz+dg9VuX4DF+u4xEMN70iRHVd
8Wp2PRznyN6QLC52sm0fGNzPkz8CTpMQfnSmuXh9HQ31tz33ksW8ZLabFAr/Ks+V
300PwJXylFKJ2/6UE5NCKibvM81MSaBJPNwbxuWm/it5A+E52SVHO1ElJkXV5os3
+n4OT8oWEnnCkrW01VS6d1xT7S99HXBmxpPakvch+0mr234N0HZtb2rvBNGn7Ceg
hgD2NYJIT9rpk9LsjAS548WWppIlKx4nIeH9yzs0RN9SnJjN6eG6ex41yRLQepoa
qQ/50coSATmN2yDtbbxiUEjXLpdSaVW5U5b6zo0yeIinzpKOpfWIx8If3PUM4hSm
uWotr46M+gRr9CbczEk7sP8dgE33Q6shF206+MQDGct3/rFe36fNc+WKlIMGFujF
OCmdnkbK4hsU6trYsgRLzk2UgHeju6zRz7iRvVcRm+Q6TWSFTV9K8qykBBAbnLb2
MT7Vmf3sv79YjjcpNYYIbsZurMamFmnbHwK7Xn7OD++nAnZbMsDFnjgrVEiljbEK
fwkOygGVXJisC6OKqmZ2lbR7g3cnxEukXBExPcibG4Ne02Q5jsb/6x+lnilsHDez
2w0JAqT/OdHzkv53EVAQY4PKN9T4KWfhXlxDFHueFtEd2otD7YC/5f/KgbsccZBa
qzXK3D0NMaEfyvEg8V7br+olNMWRFWtkO3J72ooBGMHxoXK2uhvapAHwKlnOgEPN
xrUxXpe09gkSrbRHsQiU0jT/rNz3+nipOzW3PUiJ+bzHn5+dIP7miUYOBpCdTdqW
HbA8zF7wCOJi7uG1N8pPDeT8L/vridCqVZV97AbqYxokFoxSgfbFp3ztcVWAMlcC
MDWXZLrc02ekRCkMNlRlx7O8J4CtmwWqroQHQs110fJOVIeUWdunwrjxeKa+97YN
aNYKPuFkOUhxgnmBNyaVq1EfzY77MRlNwRc9iUaYB6/7u/ehMTCtMqVUC9rM6zRn
RzwTfe6y3w/56N2vHDliwoTYFkzUEFHAd3KvtCVhp1sNMGxeGg+y0AI1p++q0O5G
ht4CqlX1mlBIttzfKUMe7Z7Ru3UlDt6kqsJzbxtNO3ux4SoVw76p9NzOsYJYhqon
k73n88yIKENy3NWeBIz/JlTpmyQ+C/rT2HrjomGK0SG36JvJc+GPjfDhEuZR5eoJ
/H7+29lsPx3/kJ4RgwRpW7YcAfuMdmskY3XVI/0UHAms0ghOVaVKF4DYQpasEeex
0geT6oMmKs0StKtFtZoNSgJRRc9rzPBX8oVDHyp0JxC0GjXE28j/a0Ldvknt2zPN
O58+btDDNUiuB4UBkUgE+NKfqYZIEU2aqK0GJwE+x1TuMNNiVg03TMrAJtguLuPi
ynaWtaoQ6Npyv0UE+n8E51oTsV7fTZ6PMna2EO7nuYwRLjxrEvu0TvyJF38qlEjZ
VsGKaxAzS2ZfGwTlS8VDhox7gegYVG5KWnwlU41h71KP3pU0L1aQtmqWbKPrv5Tl
+rKYCWoUBbe6AJA4/rJdYHYkUILU+CJ7IwYkfhi9/VfXUhvZtmds0kFmMhUhpxa7
QfHxffQYMj1nLC+vLMwq18vKx7RDXMAHkppWDg9lqCanEuMLaTHrd1rXIvALLZO+
btVYwAUcsOfa67aF1orVYGH4tLm+FFKtEZRdw784xMX/cVZqA4cAl2ncetWB+1cH
TV+x8MGd7Xb5p4Ds9RFTDduCPol+Y1FZ/RGARFiREis0EUpx9MLwrNcAhVa09pPl
opz3Wtb/vbNt6YR+qJU0Dymbe3wJcNCTvxT+qXDpAPHVg4ikTFjntVxpe3xQPJie
3dCV3CYyVZhMyl3L4rpiz98SqJN6u8U7zsER5DZz6fahlN28i6TiphqkPYg236F+
jiLdQ57jb5FUEl/7NtQfwo458YtPROXfF6q1jB3Owz1mgM7Yuylg7J75QH6xguoY
+pjlkNYHD5LxZt1iFqYil8scDFcnBh6L1OUm5QAH7VgckBux2kbHOcUjW/64N3uF
S1rahF/AFVMLyth517pPNXqjMKP0sGbU+h9DDTSI0so7bIGqjk1C/KaYF5qlQPVh
QSMR8lbyl6t9MZfVPoC4OkQMwfyztJRgglp6B8nPzEtSWeKElMCvPSFtE6aJf2Jp
a+xyrXIxLm6ssLjG9GdhG+GEquQDJW7UFiNjxWu58JH+YnXWNCW4mEhHHvCIKnO3
qe84U7R+RXbab6HbZ8vnmcctu3VwgjjUdE3bm3+QtYxdxpDSrcLY85cAHLnOEaEf
tDZusZKkqSCd01SEupPdkpHMWrWZmqTJA/dq2pRQj9agMplPfZ1FS80NsWKwJ/9X
tEYsBBWj261dPo33qdj3D1YaGedTc5p0tDn3pRC3CTXZx0EWh5WUnMOndbeIqdum
aDWWUPIdrBgxW7cGzW/Zu7X3a8PtWcZzLPSeV1v4CroCEnwd8KV7toQrHawICDaa
Y9FLJjhve7pRIgSRC/k6ulwwjRFev0gkuXTV93q4gHRQsrdZRu/3yvCz5YBWezk6
Qd8rYGCFQweE7O8JQUQA1ovCi9SOTTHQv8SmqeP9ICnc1L+e/bWF3Z3z1r9kedvF
y0gZI9EhVt/6NBHL5BxZ0cKjVH8xIY3RaX3xqmlIKL66yPncKh21f8K+ZHtJtfQl
zi5wwCtOwYnlcdZyOLqvBbrrxbYLbM1+N5uBD/jfVXhchCVhGXP0c+EpVtxQDqEr
wIeb23X3QeAKHydvkopJZJRkscp+/SanDMZYKGtyl3z4RlpHkMt3g9V3VfC98674
6nd3YkP+s4ali66w3pE2XnIga8kLXc549hNi7/nDrRJJ+d+q4dCGftgxeAHCl+qm
xexrMieShqq4nsA9Wjrxk53VRTSDsiqWeIZU68tCHHQcex9BPUXRAhSVEDjMLa9k
foE8qCmCJAIGTHsCNiBw/AGFqrPZFIWZLpxL96/WQC7E+5ZHI7C7S3R8iGYuq4X1
l0VfpMP9GXJABUZQY95IOyGOmRrDHl0+012yoy6673IHm3ps4V/XGkXZOhKp0tXo
TBzTsJvlxz8DvMUOkRffYs8bVa89AI6k47xCZ6KscKtXiGp71UEVosJiajlNfNnT
iBXNMfiweJpH0lREDyuuxAmTWe4asBeEzUrtv3ZbfjwzMxz57Rn0V8j/sgUoNQgc
nKXB7uE9LwVC7b3cMYOF0icg+b7xDW6OAi/Mb60NUrAgE4gkeanlGCqevDmTlzSD
CB6bL/9A3mfkFrzY2iyYZFtG1e2J1kjykJznUrIdI6+jCWuay8V1k5O71g/6sRJp
yOxTDLjIzaZdjd1KM98/WJ10NjBmS1fIbUKvucUv+V2BcUSqxhsENm4lgVmUsrH1
O5Nd4RrPQKt+Ik3NKFpIbfmB+J1AMdu1VNWXFQutEOPLlZuHMwhstRNNPMgYmIfw
fcYLASXnS2/4fwgjq/JtBVMizt/Lqa6ZnaHqYH7Wy13D4jbDHOmshWJUoewX9ChX
7ODKw8AiL10Uq4KRlke9hbUrTUvPAFbccnKQ5tB8TBeDd3OkTBLYUlb/CQCMRzcq
4P29/tZRuk3Pg0AMNe8Cdo2XnlNt9s2ee3RPT+nR6+9r4tKxh8DbPROvG7EaDBp7
tEOz+wCt1bAE4/mw8GFZIJLcxL5xOkl2mUU5sgNxJZYaIu77RMUUuIKNrtMncUSw
+qWC9pCbKY1mCl27xzgeWjP803PptMNeUlSrflaxcQicfNF5qwTiU3JMw0eWRqp8
LAv0xkrIUmJZdv8hVBN7mGJtsWMBCdVlv9aGtsK5DQgAJqjwgd9G+4DnwsNlOFVF
SB7n7jWqUhO6gIrvOzlQDO0llFRuTk/7e7WjDaB5FsacpL8sbIOwCB7KvM2I0aH9
OW9udghBkIshtUEfKt7jUJVLHwXZNWUGEcXlgzkiwfDoccbQR/XHp2YuhYQEebzi
ZF6SZjVyWJ+Y4hhpnkVyFT0DS7DpW3MnrnPoSgIh5iRmMRPnVoEP1tfinwczB6mG
tOqEKuAVpttJAK0Hzp/FVSiHgRKBzddiW9uCqUdZl6tBFezjbp2NQno6wXAgVh5Z
C8dV31JoWp7+U59IgPWu02BTr/P/PIQ/9zYp3CvxFfi/btqRO1Rgsbcl85JbehIo
UpRcjnjg8WgPg6OasuRqev0kuTNZ/pQJp0LijzP5bp7fpGHE+2K4mOQ3oF0JU1tG
4W+JJCy9C6BgmoV9XsFQPydlso9N2HUbV4zbHg+jbUWGD+BNJ/DcKp6qzHR7KfS+
qdsFudysRE3JVofnV10zRCxjvMI0a9CSqzWvUVPohc8Ti9hdg4UY9orPtQ1+6zoq
CLFv9eJe1BlR0TZAyWiL3z3TUXBUJhgXIoWEB+8CDMJ2dWlZEYsQsc24kfvL0vvT
Wf1/WD/vqqyPShFHx4t3OQmjT2nDjPhAur6W4mik5Q/+6f+Pg7BqrdzFYSHFCrVb
1rQFE/uD2yU5OiEBCWnTPa4UywwyKBgUPabu/vHhLgHKOuz99qOHYJSZBTjCbeRK
kUZaQ/BBAg3OUTBG4hs6+A5ogQfdsJtl5x20BbzRuhup9bdsSxgSQDxKSyVwXKny
ERty05sOzl7vnq10FgI6p525MbLz1sD5z3/lS4p8cvHeTNlFimo0E/S02QwLEchi
f5CasSU+/f+476ZZUPV1H5UgQbUzeffP9mc0nysFaPiHKXjyvUgG11wqkC1MGhm/
p9dgVouvji9owM0Dx5z98N73NPzSUbkMIVtVVaxCswVkjsh5xnJNcjLKhRFKJvd4
h9E2o4JYcOG5OQqGoOeXRq9rpMB+yGBboX1K1d+52Eh7zyXhQAg1qnGZax0GxFue
Q7x4eZ7Sv+XNZko0le8P8Ef2XTtYLlad29mcAkX5T0y8Rat0k2cULW8Kk2kXbsS1
pcQ8s1vB4dn7dktmElE+k4lWPGb+pKooT/DaUIkMY2uo303QIFFDK5gLH0s8ClT6
5ZgJo1AiAtp7QMMTEYg3flHsbWwcitmx5p7Fgdxkry95H08MoLTpNx4L3o9Bwdva
N4Ja6PWNyGd716PBeyVJNejn+lR1Xz70v1vvHpmgaj72Igu3WN9DmQbf+zjY5soX
+ZhueBzJaPz7PdAO2siL+w==
`pragma protect end_protected
