library verilog;
use verilog.vl_types.all;
entity decoder_4_vlg_check_tst is
    port(
        y               : in     vl_logic;
        y1              : in     vl_logic;
        y2              : in     vl_logic;
        y3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end decoder_4_vlg_check_tst;
