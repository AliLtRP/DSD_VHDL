// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
C7ZRveVEbAManWsmrP5qw905VhS+MAGrYOfVufqe2ByKdtF2t8bu8/DA6Bgq4DFkec0TtCIw1TgF
S+leUJgiptwUqlRyX13f9EQAEFxE2lY0sN1L6VONos7quEmW/E5cJsY7iQAjbNtpBcC9li0PNL1k
Y+uKaHvHMsfleEUGnd9aGypcM7nqFzfdfGZTmMvvC2C7NQpcCMGNIZoZ5aorxVv8uj+XC3XDhwI4
tNzvH5Iub8/VEam4hXnU4izwQVwj3NWZ3DtkHiG22GcR3+22f6+61caBvxIW3V860TNE+HSScf4T
GoZuAhtyW2tjLNIignji9lBRRB9ksnAM+JJzhQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
TexKJrd5TBghJHtcHLRWjrqq8juCEkecekhN9w8/3YPjAm/yJ7WICkznUnb1UNr8zUca7Z5uz8Rx
qbwdYmxXmKrR8TIgev5nrV6OU/Rx58KKoW1VEVNuEq0gBImVA8aaUlCbBdhm++6HJP+6z8N8cXrX
TqXOawibdhCUv5zn2nFr+Vje8qfHUytQ4gU12tGWir/i5myHRwtH9cEfH1BMlmsXf7ZaLv5ltMCL
68UbZXXkILlwyIv5lz7hJvvWxV3vUAzcIPdc52QgR1RCOKyK7mloS+eY0ncmYTFmdkz6eDWbo/As
8pUGiLDWKvj2LOKR4grs4kIaQuvKO5KxxclSz/GUzKFvpE9FoQzoT4c/K1x90s+vJ1ykHdx6Cm3J
orca1FdKXwZgwtL0CjTpeMz+Ym055VCuqwqyZyCknY4SvkxpbAE/mq7sPLDNwX+j5bemvPa28Qs/
ZyRujCJnSyXozI3GZKwIbBgpJMTweFUUPOKcfhJddLW3d2YmLJEwGz1EAOPZ601rLCzFUDKs8Jw9
+/1s/2hs2m+37nQhwldV0//mqhbCKxskRlEnWA+z+VYP+6I2k/mRZQcMRoOGJB/+REs9wm2uj7OU
GQ8h9NDm3yDIMFsEid3YP6ephlWSqrK91ToT8dJEpg5tir0vZgYUutu2P/QsnccoJxKFc+i4wqDj
QD57ypi7zT/GaWFnlCkLhaiVK/mld4CawUDEXVRls5IDUh4vo8ddaMSgEVR6mPrROoILVLVSYD7J
/Le6FPWKzw5TkKsBS4QE0olUF1+OdzReke9bFEb2GcH8921efQUsBKZvJwhi5uP46hjtm0gTK6Mr
T+LxsntCoPkicmtIHPf3DNppHgOfe9xV4tE1porDYPDhlcGveSTu8oNAGaCb+dNyARsorI0vpITZ
nWX5AR2SmynY/NtIMsR/y+4v3OFaf13wkd8Rlx3miTmZxbSU915ISNOUGemtxvpS2+JmlLtnnpgu
1zfsyB/CRtesCrBeBcwfRmqRnUBrXfPju8aLAEG3VP+4QTUr0iytvU3CfllnGzX5DY/rfwqd+A6W
upqLDhECk1v8M88hE1tamaooemSJdhEQLM7mbH7XadmqG1eyQRJV5hCbZknI1Iu9o50Ofah5u6vr
vlxm8CjiK1aKBxkKUiGO1BAHCIm2zrxKUB02utmPBOo4FhOD2+ZS6kgce4CSkbMvnI1O2V70oy+o
TDg2XanB5Kc76jwiNxC4rWznL28YbjWZy5teMFpAs/Cl2g7TCmMZCzO62YRZyxcKMQR3JmFhiy2i
Hj3V8pteceLPgcy8uwkrzhD1/cF3mexRY1S5140YwO2v/ob1qxg7ZQ6F1ur2m/AjTA8wi8Db5bar
AcSK8+XkCBh3zWEbG/FbAHWdNCMgzj1tmPtaalvMsapyjiHTs+7lsGT9WYxs+DfCiF7vWfIj3Eyv
7m9DZ+fzP0kIoQSVsYSSu67gRQ+aCJceua10PmtJ4VENMOuvnzoPGmi/uEcZtxZtULPxBQNTRioK
VQz+H0Fl7RPCOe/dbcN6TdrhNeVbk3NDTXm12DxjEp153/8batsmrND6HEMlBQGKOhkbv5zQ9/6R
NWN0cv00PHbNnUiHNZJzdTLHMgq34iqBAhA6efRuTn6HzJfqKECtNHp8cAqfGrlzmJIMufiRrDCB
ScpZB7LEzRlVoHygDRUuEQ8U+oM7SsHp+EscNsleoNwQwPwlYMl/x/AuUlXCXYE8FIPxNWi+JxOS
Bezv1YUaMgrMLsOoDyVjHMMIBQxMNNaspU6gj6pGN6mMNi23QZpMWhHHW6CWtVtcuYJxnSPyX0c/
LR7Nq1KDiEn9UCPNo0Q/sabBzFeU4AtjL7rxlAGyHHqChWxpyPNgMtOCFValRBCalN/qE2jSahA5
r+U30TK75AgK8ZAov8Ml+9t2XbhJVpg//AMog6OT/2aWF4B4MXC8lvLgAka8M9Uc0mwOOvo7K5yL
O15SxeLF9MlvRhz2/vNbGlwQk+9KHI58rI9rGHuwndMWsUYTEJ/seTIKuF85tJnFMFcWkPs9sOIU
CXTcCsJl7GYp7oPomNM1gsQPrLpWhAeiytGINAo1S1EHt5MkTmRIHSKIfZttdS83tz99s7p0gXSD
1nC3lBe89cfA6z6iw8LvHiQGjl29vVq9jBdXmWWBIOjrMml2n2k5i3jdVyxDwCyMCMuo/tzNzaiM
SzyT1MK5slroBvlM85nBLQIBz3oBSSzMj3D3tfJlWGhQQDPzNbttBq5Ipge6sgkm3nNU0Xrc5c6d
0f1LD0ENOjaUcmh35YK/RSu0b2O+k2EZZaT2grCYtdmYsWLTLlM0oitDp/M08Cl/yJZOJZuPnaWe
Vxp8BG1AQkF4yN7U7lEF8kqeBctwOn6C1wZ3N2G7DG9yrYQoLTk/H/T8TyxDkN3/h9iAhoNFums9
uuC06YE5tcGkMgNrZ7g6C7oIcgPCP3ROVBDLEGU7qLUIiJaCiJF3fMnCp8xpQ6m1iyhV5ylRDc1p
GBxyrnZ/XosTR4zhgXDN0ASfnEAaCnNARp05xXCmP4bHD0oJd6hdH0nZI/bu5crSX4Xb9B65m53K
xQB3RvsB72iny2e5904WKx7qJ6L0SalyhLp3W9fx1kUqT0A6T2AELI1qYxvwQgB4/e6ArGr2+BNK
WaQBgnaYtFuhLAstgu2iKpg12j6hjD06sq48UduXqeQtrR5fS417n9ck/d6oZUpUReYKmCgEq2gC
zw/uiRbowW2hevHKVyxdnFG6WrX5xGjYrf6xOUNth55kL+YA3JvWxFw+opb8/gkiGhzhrJxiXjWG
5XyfMwCLS/ACWSR51kDYSpPjjeBzXhR5sg4NhBxP90XlzUZ/kPDLsfjLeh0BGfmyLbO0PWVh04Cz
bWhYP4AehyhczkBR9a3aKlMIAKSlCkMFfmJXCcftKb9Aeojq1m6jXhn3PYgZXjP6xsU0kTUaPc66
eN4qxm6L9uDUM9ggvcFDsx53HU46Zs4CzfBtcZWbO5+D+/rB4J+4feTDQicYUrHJxmLrhE8Kh/ym
K66uxcZ5hIWwwVAcu9vzK/sSX90tppwvKxMpUSuRIG2rsWTadTL1nuNzQfvM7/3ChEhAPqLpb8el
RfZph0s7MIuTWRKHR2f9i39UZ8HUJ6ZBGD6eCDduzmMIiMs0lJ7ONQaXeW0jF7Slxlz6fRp1l6tO
Z7G1e1+9Ma/e7vjuC3l6qFXVeiuUdLiz+4xz9XY9hD/RY3jFlAdHBxIwaeSkRjJ7HF+yS0FdaRi9
aPFn/l3JibvMWJZh7vydvC2qZFSrZ6mmN0b96JymKqNNTIGpWYvkd5MhHI4LBBj4pSWm8rVvi8Y9
6RiIyoE5FxoeqM73axgyffcWukPs+Exg9kqouCVZnGhSmR2sjTVyukKFpqaaFJgSvFiAZgChNtzV
iSTzEnssr13+XE9UtzStjxA6yGRXE63GfnC7p8ierdiLHxT9QCKaFKMVEhPiSkmRgCwXnM0LeFon
exLW8l7hUxtwHF2khmb4m4Eq0Og6ZJaHeCNTQmaAMGW+Y8w/fbn2t+3C6Geowq3O9G8Sx9HfCzyW
IHhda16t4YRjaAy488w8eN+qn5pqsPlXkAjehyblfzAi0F4AwgdaL1zhjrUWZ2IhgtJUX+i+FrMG
c3+/HcOWq1fsrd4p5mTxHQKHze2pjBAqVafqaagG2zrloP7CaDqFH6KDWy0We+eKXYEpNkRB7gkB
mNsC98eB4JUlApnC71C+LBbUE6RuFHdLi+yVZJ2efObOETIzusmmlQnJUt5+UebTLK5hybR1Ml3l
0R6xuI7U2lL2z5bHzfxfK6L627cVBd432WhftWKm+VS/pdBH3nokqsX9r4u0kKuHsB54mNAmsrcP
ZwxZfi+M55dvsQXs3MKeKPmQsvIuu+uCkpDLBW3e0gmpatwb7HowNR+Y4YjZ8zWO4wl18kybvu/x
K+5wmA1O+BhG3N6JI6f3nJN7i3eeEuzJxA9vtQRHTyygslWw5cMrD9SeZQ6qdYa8FlORh0rAqJUX
/nvn/O+Eop4zaFwdJ6u4rU+3pEp6I3u5IC/jrHnLQ8c37zTEk2GTfP7Pv3/1Q4aVjYTH3zuPJahQ
mmaa8mm8TinViYWA2+7Pdm+hsAYM64sfrYMIk0QDDFrxs/43HGsWLERa8zHmBykelUqXX6Gsz8lQ
6l90DEpmo6uMhMIGR0VAlg5Bdpk6BRH+kNcwPrqwnPESF97Pl7EroT1gPi1FfUmd6VNOTy/dRW+P
IIzVSgKwaRs3H8dts3MjzDqfBwI8rgYdOEuMxKQswi/b/14vSdq02jac2V/J4jJycc33dh/I5HgH
Be+H8th5dr1VjLzI7PRsK/RZxm79jcVhNZLB+ShggFul41ZfOe3EpKK6r/srxgaLzymTOdZGJfsc
wnQ+F/ww3sCkKGjyo2jkxMSGIFXImtnqGyKmiC6Sbi93m7tBr8bCGKLbdmt1otUDv9T0aOXOBaOQ
O3WglNfyEUnIzGlHlwCu9hqXvH7fABmSeJ7MMnSh+2xtlqWVvdcrQqpc4ltraC7KoMDv6aNZnu3Y
RuzN1PVgrtgvXBy+CLK8Dn6KuLPIgUf16oL+cPfnFMS6GFqxJtQyIDbMVU5d2ajBwrAdDnqmocI0
dRwtaN+L9Wb/yTRoPMkwPgNN2K9qbrBqccaK8hVgMN2kxhhao3+9/3gmlNir2kLPdIt041auJJ5W
f6kD7vncnaSZIO/7ZQ2whalSkCqIqd5FNb9wC14kg8mSPWsGFpKY1/QrX3w1jXzXBTghqNuSaB2T
2820JEkZ4a6DheQ5V2O7CSOodDP43D+TYnzTAtu+zjqxY7QtKexRI469lqboYXhWlSVcJVvDAa2X
zM8rxsVGbXXN3S9WHhvAo2UB5s2DArfR6QcKwCyPVqctgAvUBq4jp9EAL1aAGh6qXTGy8fZcQPie
HSH1QJY2U0DkVnSGcrwcFOW9G91tQLzIzkkrwstIu3Zzopb6iArYYBgYbSa/mLHBiUgLkTM9n4A/
DjeNjnhd/wmBszkEfT4VVbS4yehzrlNP2vP2LF+Q34qY4AYiEdPbt0LEdnsU9SBEBvk30I7DXsVJ
3ypCHI54KMNjRmHiB++81F0HKiatO+/5eUfrq7W/TG/y+DU5X4FSqk6rXVfkYp47l3kV74OuI9jx
IaDvU/EekN126316khKKFHxY/jt3j5/GMNhxRvLP4MqW5/7JqIzpwkRFWpPn/FpjejryW49e56wl
xuRSc4JHzhuDmEY9ZqxhfosE63rh2z6yOHe1DzrxQCirUNCbmq7/+cwfRsRBwSwURPouVVKX61kr
K280dr0aLtU7nibGQW2aTR+dpOZ1HAOGjs3RVnJjFG3l9LFsTkrLtkTJTgFcIxcAqcsB41FNmZim
2r5w8O2tJ1+0Yz0kJlRPZVy6LRdkWDd0rjx67Kdm7JCZ7Xjvn5XU2p72GiKXdxa9PvSiljKcXrCb
7PkTNDLEif3TfQc6xwDGmUveM1g/8sVQDNOrnPFiLFGABKVM/MeVkJ7Kelm9biMUHqqiw53tGSI9
ubeSN85+2zxcGUsI7VtHcdQvnARTImtfRrdsT3iYp4kpHvL3o67RA5aedID8WdRczXYxDYIdoDyi
KyDLI9mTb4xE2ZvhzdHPpOtyQ52XqtJlJ94gul+9CwR6+uu5pEYGEHY+uBDThJKI0saBoi9dhEuq
RpJYdS+XuEgyPSRadKOkAFQCYyQAXknZEAQ4rE/pQU22uI+3XMMZr25Q2YtGfWmTrNpbFZ5+hewc
hAtuYQQYSND7rokOMYgBcfFiqnZEUIFhP12wD5LrlTiQyNEkJ/hEgNmsVxm3ZTIC3+okcIzr3snc
yZrUy9v/YW5oFF8ANjTFfyy+HuzBqux1rslPfr95v18eiclt7UxiQG88zU3K8r+o++KcL7pND5XC
LyvKz800M2ePFRfBXVOClpNWusvNSHaWja9OJQx7iiWN3qqA+SIwl6LladCS/ONUczsHS8S//B2z
rsRl3yyK1nYJRwiZzk7l2Q4XRQIOOIfoARTufSEUxhSBn2T16Ou4Svkq4OJfuNQaEM9Q1+JmdVLQ
lnizJ6j16GRHejDompPGVNxr/OihsjR3/a/Bf8qWbfiL8+c9j41gyQX0bmAEz32YCW2pF9iCl3uJ
4YaestANmzhXtjZQa2SAIs5a21pyRkdTSwhLpnQHci4vw0Wbz6/+OuajytN8ZvwoCUXqDMiQZGPv
FqXOXmLTmSGkc6boXtWMn2LVdpPug6zBcN/UIn3NfgrWSVdcO2mNC2cgCrI6T7JoaIZSzeGlzgo1
Rk9evnJ5vfyUuXnLTmrDBt32bDS68yLzQJ0kbogdL/fGna+Swn1FdHKnwE+GPd2UfFHKud+9ejm2
ewjtRKdAB0YdRHz7Ne2K2LAtJ6C6dXsgpHHmBpXEMgB+qehwCoaVxZ9mjukZa0anDQy7dSqYkRea
FkUQt3yvj87hTCM2ScwAZVZN5BdPbfB6qdaLDJ7Jm1GxZ3lDJwKwXjB8jE4zWScSVqhVuqSW4iAC
5RdeKjW3k/8uqExaeDJweFemHskQIr5TTNV0joQR9WFbmlZIla0kKeBfpfuX21TLV5XIcImn4H1e
X/KEdLeqn1m3xRB2zUQOQ+j0HRmmE47gIxkSbD4zDLi19WxvU913OWOF6lrBmsLJtKxuKpDTJ+8X
9+GukvTBhiaQ/ZKo29T80kU2DBXcfRLCJkT5r02BgWqDWUZuvuBxexlgWZbH00c5Ytq8m15gkQk3
mvsW+JQXA5Y+cGHICMu0mjGBnoWbV7M9dofJES5C6x14c24jIupj3p29JV4GwiCNo2aCSlQ4NYXR
gr5Anj+zYIKydWc7D0gJqfwXBqgz1sPXqjITGDTlpx0NgBAPtuvRTSpOw0vRe83+mfDt4pBrHFFG
Gcl7bKU8Up3f1vDjuy4b/2uaDBXS/Ey1o90R4+q4BVcdiQ3U2yXc24sJQNhF3UwdC24CAl74YFUt
MYIk3H5MC/TeCJB6MlFsf5djuWWGMp81QD71RglwZqgoYz8TvcjzbyWk+QTRaRLWkBxIvjC84eDe
Rzc20Qv/+Z1lHftFbEpiwek1UdVrdLeRW7mucQk/Uv/wcGHDIUMKPLrvYJRWWH7gY6L3DLfdesjT
5cduUQrIw0mYUFDa5X7DDGaG4GQ0P0yRVnyUcyq3GYQf9C6LxB3mmp8avNVpNGIh9tq+Xnyi+HXn
M86SP+G0JADwOEC5mDf0CwqXIkiKD1KhKoGSRey4ZatIbk0B3b+w1eMnIf2cK0+bBFEJmusLzi2O
H9k8wzX6MdYbPPw26sXvbFM9EzxVw4TOAANyxAtcRAntVua4FR3XpDlJEzC1kjGoCg/iYJj4f/ni
Cu9/UzORnc6/nckFjgoOKBlS9R0V4TSSrT9t4fStEMZwCoeyDQMXcaG6aCYH/w2XiVZxUgAmZ7Uk
gDKpgmZLPN9xsEnwOL/iPcxSyhgn67QkWiqjWSFsmu6e1TLBAPFjWKuV1/KOPqyX7bbt0KNhIBUB
gSwRjh1rdABJ5J14bYCYqej7BtWHQe8PPNDstjMcdbj+W6+NWuTrQayxP0S0livnRWt467CMVVDX
HYO/8p6SPWQH3J9HJ7gKypi7Y9hXwEMntfANgAsMLP21wIF76Ob/gif03dcBRsBs7+8owUGUA+AL
/bV6hWul57iY1dbhRseWaISE0XzJ0DlB1hx5zsO6iZ0NdWyCGmSmYIzhZ1NQvBHC5aUMqoSXQYGj
MdNms6h349rQ4D5nbVAO1uE7KzUjzQeWhvUoSoD/yzdeH6DH0XJsQcEZT+pamKcGsnY7s5ksXqeM
2lOq8fIG3BF24NT7jqwqZJXJqF9IbT3qY3/Zt+vYrykmX9y7xGgIcUxAXsg3gjLwrAJO+D4SLZtB
IYTxkYsh5tPohZLb72hlkVsUK52VDzOvOO+M01nzXFaoYaIf4Hm2uoTVETZ6FacU2yWSK5FizZFY
hi4Jb9Szhnj38UqkliO8r6qPbhjK9ZmpK3WqGlKwvbzqb+r/uh7uQv0E/W7YfjRqZ8D4TU+e3MK1
VxPh4Msgg7dmCFA0quRdsoI4qZuS9QDVxMeGKwjwKLr8SlKH3KI1JjUMwPrG4jEkeGl1dB0cd2Ui
fVW0Un7e37r8eUb315/xO+CCeYZEfefPSkD0BC1uJOWjqArmhPH8sg/qK6vVN4XT45SYzVEi55iW
IHnBnwP4p+hK5spaRkMGJr79sVCVuQAEuBLH7Q22E6DV9PlAvewjD3gxYnToskOXPuq4FpTyaoUk
IMgIBNr+61B/GdP1h3n0eFryQzb0m198uexRpaIDjwVAY7MP/GJzuGuy++f8/j1eYSMyiz5X8V6B
b0r5cOVeqA4kKCwf9WAHpq0oydZcEreC05p2NkGwhKZscCKp9lbP83gYvyRaPAzc9wQX7Ufv6uqj
gXKWOF4YMQ+bD9KBzVtH6eQ6/lz6pVJ287clxQwZvpzUcsLM13VA7soHXYgyzuh1W1ereFKGc4zf
adOpdQipxbFsjSo7uD3vq2qKWRcm6461ptzcJPIsdzAYBUopmorhNBV9htOKSiUeBTnWhrDWQ5Rq
OaGnV0GaietQh3YhV3FoX0fGkJXAXIp++3uv9qj+0DifG6POAlq6Tc44yzbpfYY3ElSyHtm3Hm92
5a68yW6BnYj1h6hhl8PAvEcJ/d29Eqj8JvNPbjMjWnW4vuF2XKc23iqooNOmHXibZ9yTwp+ntDU5
CANxWeHzsTq5V0+dTtUYdBpspYYuN9hBbNYvLqTu/qxYvE+Risa82Ue4PPXeW5ojU44zlXhXYvcC
mS37S/qngoQQTAskg1nl8kUaC1TnXlffbKH0ItsjGdg4PVdIPsbUQwYz5gZn97ISEJpN8/yfViTW
b1SZACg32LhPzeDoG5x2w6stWO1RIxcME7gZVA4WDDX4RkykiVY8fosteDAAXOmrDlwR2X57oIQN
F3DwHiiv58B0nB1Wl3YdBIHW8XFv/2zHNW6XisV3TBNjfDuw2R3ZPVCCQiPYQWWPtks/+c5xcVvC
baThzfeMexyNJHIvzD1MPBS7RWUuhFbYIbGCQIbylAWIwyniq2uB1vv9lDFt0l8I0+aekjmjaSM1
jS/8XRk9BDGv6ZhBOZ+owIlg/HXsrgAArBlPt72PTMGvqPgC/IG7TgxpykhXyDMeq8OruT0gVYlk
RShTsm3JnmCBtmvQlt9LRr4R2CRswRkc3CmQ5GNJtrzEeKUODleKgI53ujjQaKR2q9hQMg3RiDRT
1DfzeC8aelaHXpXSfLxZKt1jS/CY2ExhmM4kZ6Q+LqRXgA/LdpoRWM78cyAhui28yyimSKgU5Y/a
f9Rg2VVtASLXafruesQ0rUtCK1UN1kPQYN2H0fkidhwp7Kfb7KcB4QjluhaTOjPSnW2MEjt3fVRC
rSFgrEZLGb0NmDZg8O73irqTwOCSoR4ila+VxE5qdSXHN3Z4z4J4nlepz++R7dWBzRAHBSYUCDWZ
TRxnkmaWv7G7VLNdPqbQRmy8JCppfUt8btwehCM72QHpED4Ldlypp/REXKCxGpBWcZQzL6KhLnx6
kZdpBWH4tKqbwXjaiiYSi8c82iT20DkTdp6ixZt9XAc8RTlqzeQ+hZ8A6VBSMtA8dFuqcBbo9YKY
YwMVi7W8vWIwaRgobTvyvTUiNuXMfYwnsWJ4eaoPF2RYsO9Xa7U2lSIuG0oMa4ks5nYn3105Jp+4
MGqJR1VAChJ7f4xXjMRfI7eVDM/nFh66Cg9GKgmeCUgHI/TvjC52aUtC5SiI9CJPPl7PeX/Hig3Q
Zu9fvcMtfAdXyqN9spbrfUUXdfdS+/dggBaAxnZfssYIOcbjL9fXE9x9ZQOM3Y10lsy/ou7nfY7X
MSf0K1xqZzDf6w0pRGvdIQS1xioAJjn6fu/G/h6HTjn7LMBa7PgVe8gKzCr119wm6cXixvnluvpA
GDNCdxZBYl3/VdhQ301lIEwGkPt5z9zMfxrla4OSOaW2d/GZUPdvql2Au+Xks+gvkosJoTZfLptW
8e/e/UFkaCuehrU9otNJWyoIf8olbadM87w9Gy8aPEq5Ntr+/7IPW6vnZwcwEBUXAAykvXk/aUkk
9dJzK0LklxOE2ZSukUTW/BmNgCwpulXlVy4gTovpJQGAxFra7yrMGcDuezBMrKXi+AftbaOQFSJS
qKv1tiID9vEStf38nSv8DkTD9Zix3dSwut6P0gFDCvpvX/JMiTfDB85cx86Ahd7GnrGovxxE42hY
/2EcOtz/Jy3ZeZp5Yj0Ga6kGfAEiispbUShbjKdsJTPWdT5tv9BTcJaiiOsa/+rD8kp1ty+YdJBq
XvFQHgvZpKd56W7uYk0k9TwfZoDZ3PJlMQHWUCB/O0h5bWNI42HzMkcJBzFH5ZBcRASjHbTj+qrf
10c6ScHe3sectzBHdFsLLb107KQ/fhiUZatDKWuQG5dnXhHFhEGncE7oufKfl8+9cLr8og56sKph
doN0OY15wm67/WhYXH9NzaDQTsEVTZkUtzcSGmTmK4K45899rsUgo/fomTRfbZSjTzRIL3cFD7IZ
ZcClx3Cu7eVOVLQ9rEBnE7gc4Rn9o9bOOSy71hyn/zflWqLQo/3HFO7HK17BiKXckBMq8/sUn0vu
O+cerEP+yITT3YdPw6DPFitcv7yF0QFhbREsS+8FcKrbbWBom3H0qJF9Cz5OeOXkqK6YDezbgEs/
TBW6oHT6ARkPUw7vot+pK9NvgtYOYepJNh4Zhy5rK7klRCMMpPvn/gYVjBLBzInpOixWC8JjzA5b
cUuHQYAp+bD1RUjjH82SC3NUg92MyPcEiMmyvpHWrT9T82b1xM8KxO6Rsv0Qt1ZqAB3JK30vUgqk
jH8ehJTOjCi8QYlIlMImcCPfSl0TcPN29yzH/TBqB87plWj2m0mMqoHmqOHyr6hfjqxc67R1FMZQ
QroeR9z8XgmqmzmH6xSEuh8wW1TTPGMPJijUfrUwprXrL2+8XxMUrwnpL0RruNjLrTQkGS0gS2Do
KIDcBTlsgq4FPBf65Q+syooER3CfBQTe9pFbj4/sQBQTgJ3ag2lOwc4u0ooF2rM+5CJadPB689Ky
k3a6bPRqUta/4jQ9GZTfyE33P5Q3AoAF125wDlgDvVi/Q8KAM2Sv4aKy8ACIBdZFdkdWsV2pBiuu
NP+M65KXVZMjE8d/fK/dzeGMM3kzUoOYCfhpz4HZHa8q4NqOt7EhPVZEZZFCUPXOWKlv47fGJzA9
wjVq67ppbIjkzYF6+tOVnrZjy7khzZ/C8Vu2sNDq/NVfU6+3RWZFsJuwuBYJZzsAfH8vwqxE4m7S
0GIF/VJ5ojGjoFTk+SNL/xwJw2t1ox7ZohkqARfAIHumI7o+Val0dYeUzrobjJczDTf/Ajs24c+O
tcIfMQqQAIr1nxiJyWJYze/B0vn6xMUdJ8kMgdTYvZv/r3ADgqSlFZAwWd9qAgetMt5PgO+u379k
xcqDord4cjE6xELh8dxZ8Q2vXg5pqajRHfyeJyvUUh/AZ5ESTUiTChlHrodmigW/RcIYjXl4jMx+
DcWHymcq7umUCWu/VbRNqBHagJ8fI8P3/CqOuuKrGQdXZcPelvlmOVxQ9r6kWI2yv2CsHprMAUkY
rGxxgXLBKEE89vylk+v29AAb8/1MX1GyktQqMrW1S6P4kSL4t37xzOnBZ6pi+p7IrINsz4Pf3zgI
5h9e15WKuLCr69Ds6DH6GR8v1cZiNrOZPr3/2No2gSMDcEs/VVj5o1kmMksUnWosCArV/AANjiQ9
JxXn20DgprSfT07cPjR35XtYtnyUn1R77GtuC6Nzrujo9vpmOnU/nq8P5+6uSMDoohl/825w5O/5
xgFirenqawa2dhZoRHhiQBsmpNxjmM54FiBOvPaI0LWt4dooReL4Tg36QULQPqbj8nUhxowbZ/BR
U4+iOLBsd8iALmXHJW462/3c3hWNQx1qZo6Pex7FvCaFsuJb3v7Glua/X7Nv5BA+dEoe2BmFreFK
It1B2IzYyH9wQ6bdhAZNBHAx6Qon06LmIXRaDgJ1W4mNJ/P6iSBHzrbdxCbK60X5YEkcX/bjpTzr
MHR1eKz0kWJEIxKhcyMzK8HoDZ2uMgn7xwntlMxOnX3WHiYIkHvQvbaKOjDwHLnHBcZKS4r3H3hQ
w0KbjR2TpQDTPiheeyXPLpCs5BNAksWURTtgJodLSF/YBkOUeOsMN2ZDm05s/IpFxpQUOWi5fNyG
/DWaBW3ccx4kAcPooQ1LRPXPthkCpxd9NSJMzCk69OH6weRd5WjoUF3w7vymlPMepJ57ytH4cfyU
2hU7IPZklLW+IEskGaSD12QPqCbkmXR/iNQAyJA9XUjpt6QwxaoRb4B6a78MIXRbB57yJ+z4jda7
mjjfGCrtH3YxLts/FQixR88OgNvLBqzn6N4jkxUhCSPKPL5CoCT9cn/n0q3PreTtGESB+b/M5aDs
kZC0YsOlM5e3euiNGCuN6c3ZD9pLTgbtC1mCl2CpNJUbBopDfjSLYZU9rK2CWMnod3h2Y0Kmw6Tf
MxgctdmMiZx/D6Pw+gsxQkDLz+JeMXjwfMmll7eYms1l43UAqXvVoAlwHLMWv2UMkltwlaxt4H+V
8lM7YkUWPj6C2n8Nuh7Zp7JyriG4pCktr+eTp/3SBBR2aGzugvAz5cgZGSdrtxTYu/n/mTlI+rFC
Ik/gICwDNfrSKUGwCD/bemU78kFbhNkbu+syZnWtX/L/VBEtVjbD3zmummb73bA3UoQE27l1Nu09
y91++eMtiTdnDqC/oLBKvpyuNs7rae31H/KYWDHWv7Pngs58H4eNHgip+fKC5bN2EPEGoTGZxOkD
ssi7t3Zbn7a0qGit5HAViHn5qG/XaYssxoJJvVhtYfA6qekjpwxqUu5lLCWgiKlQQMdht1RDgepe
WD7lKyuPkNwOfD1BKDQHPnjtMSdV8W+DzGyY69Wn8dMTXnhq1hy4eHBhkNlxGfblrB8QLQuDoJxP
EV5u7K04yrnm6NP1BIDh2J+GCgLyR68NHl1XzDqrSpANRJASCpIzlANw00dwV0hKfrXg1n1pZU23
L5EAVsTA/1NS2Acx2/NMhkdZTlRJfEJ2Taqoi6qdCO0+dt51olyritL6+fD+TXDOcfGVjwzeFWUx
UqT0FcLpCHmsMZ+ISpl5p6xsgwSN+nAPiwTMnyeB+ydLsbZLyPjAZUG8jEWP15oAXaF3Op6FPPVW
wOxpL51+U+e3MYDNg8IFL37P
`pragma protect end_protected
