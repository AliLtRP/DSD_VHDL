// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
G4GXgDopnuhYggS8Wdoz3kRrvdEZEywP+ehfT2xHRsrcWsYP+P418aEuC5jIMfQV
JuXxGpEeZ9/PjK/ASsTq2VI+fgp518ew9T4e14za79Qu4OxFtH2OFLuhSFW6dOe4
LdFlfJHeUswhDvu9YNglaqumfWGc5hyrqL4gR+SBh4Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6448)
xzNPolzTV+GLUlL56EVlxdF8RNoGt/3NU5TRhfn87a6IZYzmUhONkOPOUhBhckfm
RSIo3AC/BQtLwu7bd8WxKiA6XyxnwfBrOe78gK4p6xsWlgcQuXCR5LHHuLh4xyGC
ZNRuCwZZZK2UrRjejCdRat+ELKW03HliBFPaH1+nUNs74j+MU0+XdjxGjv2SR9vg
EuBdrpFdczD7GrV1z0ghD/odhBQY5xROArUOf81Kk9zKsUuMPF4BGiWVC+29NVfC
o5l4W40eoGksQ4tIm/VjSdIKkxU3qqH+1nACh35QeyhI8i9ryw1H4Z/q7NdW6J1H
XQSWZ9iqfMHM2yUZx+Izdia6z/0iUBy7evy4to0MMRRuHhx+C1sK3oBOdU4YccFF
FV3gqfSXZkqrPg84dF4DShFkSWTLOye1XtAF48nqXdQw4ZI0AP5qjth99yEFGDPU
xoy9aWxIJHjRyMpLEp071FqnpH2bmLWu/WxpU+f6uS+suVqqnYll3MPZiJDIzH5+
4ru1SOqtZjVt+glwFel9gn1hm8YwpRpI3g+w7oqh79iwLyXmZ8q8CkLBEfOcQTTh
UHv3p57fbj9xeDb0AfNu3ULXIHZIiH/mAJ1/s3pnV2L51QuzMf/hbf9ofwJC0jBX
2tgVxCwI5mxsrAezF4DcB4Oj+S/jvuteJ7e3gPrglYH1SS6cMOwEODETUQUD8ZdH
4yAchVT8jrUsZdneDGzsKztdIRXVXkra12zJCoZ/H+YMJ2B8JpgZL5X0H5EIZaOm
qmEcP8H3zAQFhClNNdrAcbaQ2QmR5ZzxwA/wFayDfWQSUoCnUQLl1zfoMX+lL8F1
3E1vFIjkoOFPg/h583A2Bw98KShkHdVWpVG/B+d2ZuE9RxCqwrh6szin8KPtDUr/
nYROjOk05IabWqEU7DPGWoXo+oqCqRpflcmdClYy+n7HQkaGeaTIEkwlCPqj1QfU
osE+uMN0xqeKdJsbljTuBDdyVyN/IYPlEEimGMEvnGf29XZ0Z/Rl/wqM5Y5dZtAI
7UdcTZxmMrAyQ0I8E+dKNlxLBXGUkmB97iglk904eAEXysTdlIXZvCvvJ8SQurS4
V8m/QMp3X6BaYPHb97Xc7owJN5OLVvn93Rmt2XycpvQZDjGOEJNZmq43bZ/5cszf
uDfMxc5MoLBARZR+xFsVWj4+KkMriwUFOf3EI2hFZSsc7RSNNreHt75rVUNuqyFM
J77m/FG0ecmKGVgVk/QqNn0+U9hLnx+8vlvpnQfuIvOfIQQ+1u6omXiofKLcYQ/4
QLyeIBNAum13SZWnzP1i0pugFcTcEhyxk5ELvurDU0uz8ugdo2kVl77F8PoHAmLt
KhOwGMz5dZ6nJoHwbcE7psSbdCuCO9/z6jHoLjMk8Kl4vD6DxpgzGxqhPSGMfYaP
SjCzgtvoS3CxiVM9btQWlIIOe7yCOkJl+KE+jzy1BM/o+mFRaPAG7Yl9/SS/tWEh
BtRRxtYLmbf18O5pbsKilmv34tKiRj8t1ta+NpUWibzC15XOSS4BBVcgY1qLhEEo
00bqO6/SUPnDM1zpzf2GwfEYNqsXO1gM26pjOATbZV54BAY9BpXFRu42lBxnOdkh
ZnDLW9fcXSYSMrxvalBZUvKWFmVYUBxjrhk8SE5Fpubc9GtpmQ4JKxP5crHapobq
xc4teLvdsmdZ4Vl5IWXvwcoB9IHsOrGXj9BR+stU+XoJddVW5OiHO6iMbsOfad0y
6UCZWDCUD0y/jkg/KUmNAbPvlCmyFJny9+PlsWz26A+eMUoLHDPUIar2BwRU9qej
FC+irfuc8aUYPa77bvS428qDJvwCgbgIOgxBOAyKkBwftbLFvp2hjyjYB7BYV46G
J7Rp2yW+mR76q/jMYlY3ELzDbxQ+VolAIe3LU5FT9z9T4sTiYIiMG9SPudWiJEk4
nRUqtpszqr6KjmKv526flBvZ7kRpI1y08v/dOJkBe8uTJws2AARXwc1rjKEPnJiy
POl3thJJS9P1IPSTYqG7tGb3KPF1m7980iyGnIpC3ynIbt8ntJW4xQqgbPaKT4Bg
SPrFBw02Bdh6iYpWMNR0Wycg9kjuhnTUGOfJqW5rQ5g2HI/w15rga8Aq12PuDtKo
/Bb86VRzjd3QMhjJcI5h54CSsPC+uP80W4OAp7/pZxXXX3C08D0i7Qxmxly8vHXN
devAbSnn7g2duUvbdnqVy81QmZHEvPEl2PKY7EYVTnMGE0CxZ1T9Gg+a7XADhyo7
Y88uR1Wxh+ESFoNQT7U1sDdiuJ++x0My8Pizufm5NYSMiQ8Ye2EDjakzkMLOzjDC
5Zva6RVURam0nJ7c61jwM6on/96WHqMhabzHlAEepeQ1CQdeqHLFJZu4fSSiMFmZ
i4UwW3DXWP4ukuO47XtwoNZOPGM8domsVKFjgXWTzsCdhnmbn8in82uC0uIYTC/r
9Gl6o0XuQcjAx9AoODrjq31col+XdJmqBjIl0GA70fVlBm/rVQqS/oN+3j1p8rE7
UOJL4599wBUss4zp7htSmGZ2ITybRwy6xoEiTIDZs3e0GA+Nhd2NlfWHvC2W3HlZ
QYcMxBtSYS81k8Hm60zv6viXe/Yo8LicXNtZHzNoc1MoGT3lngz/dDG2uGC7M65F
ANfF9i4VKC6+5RHWbbp+jhbEDyVhqNP6H8Z2kfnBBTpW0/bLV2WUT8oKupDJnOSZ
ZcHxHzbgmKywMBUxERZFMYLffjQLQwBFXlfGy7eMdxoBnmsZekwq6mvB81+dglvK
fKDvG2TMRPWQ5wIgzIks7J+qFZ5Xc17f1b5VLPmzVFLtzKHAnsaG0Q0BCda3k+4q
3YlvdIimg77jjWy6NwLOyEsN3JVvGSAvlvuSNu/kHAp/W8CK5cXoySJNyO1R5mc2
KUh15TaDnb3wWD/u8nWpWUsSzKZCQ2/WXuJ/pVQl5akntIE2EuzuvTTXYTaQrFat
lZelE2vTZID/Q73znP6/w4zKflVbJxS622G4JUyIuM8E1xGjCbB82VKsYoAJ/WIu
VC1GqDxaFK1CmbMY1cL+E8i7poYrww+OP0/hSNYj1Ebm3hiLn3wmfdpdaVCfj3pL
GHi/wX1QqkjyEUAO6iCGn012TZl+FEkVeAQs6Sqg/E39ahGL5bGwvX0+6+2+HCuU
N99JpAUjqURRyEZ+CkDU5cHZ5znibocHQTYXMCswFfiSHYhxZnDdQ7BCfiEmjFJN
4EcXZ8EQS/jRnfRHZrXVfTJdtrX9H6dgKmTULYDDUzVNhrLNpkd4EYGGJiQHbjGO
k3pgT0NCTNzZMQj7/Y3sqgntcjTWnVkCxPb3GaAVD7dwfU5+lUiJ/ZyeR4jfcI59
nhJ9FJmeFldGLEB3qamVCDZHMA/WwyHc3/4B0p4yYdWMrgc7cJOPCLi/VYpiZ9ER
FahBw8aohsVybkFl+JRQmH2a8gtNVRn/+k6UWCJcbADZsHFk65S8jVhIJGlRXeFr
MEHsMeaEaG3qhikjhSInjot5aVSLiTscELJt87tA4v/XycNjZ6OO2PxUC2o6Pw49
m73GGRyyMNmn2/31h2yBeMUBEY7Mm+VYDW6cDZN0VZGRNgXr+T3jT5YObyQHpaAN
+CGUttEmpZaAu48zwJ5xTGVexFSP/e3QKjqzuPJtaVCM9HcNEEHGGyRUnv2EjEt2
Y+euzmqD1X77qfT6NjchutCmb7F6/ywg1v2lAWcs+nET4uK3txaW5RXZ2v0R+CdW
t/A1hjaHO+3Xun0Twu8Df5ebRsAMrqMBuUThqA4zB8V8C+9P9duanEDC/O5a2hpU
Xjnc5W5WW2+BSQSGIdbgL7xC5BgOYfxgXowWs15wSAwy9/dvd9cYfRUXJvIZ3eft
ZSB3dS9zsif442u/7jpTT5EzOIsBBeuevKg5jzI0eYVBPaUnJQ4rilDOFGcno1iS
d38Fla1xGwI0CFPBAvnktq7zO8xg/x9QpMatASDCA8jvvFwPKQVq9Ul9MAQGOe4b
qZuTCttIwf159KpRyvXk8pMIUmV3NAO182mvND8B1FDpCd1CsOnLn7H1gLj6GYrL
G8v7fGj3oRrYSL4py1gXdELgT86oRtnS7R7jHnyIG/yiwZXRr319nQHeuYrU07XS
MNX89G//B3jBfrFsdegnmSCk4wAGzMze9XXOaJUSRelqDBAJLY3G3Xr3rFl2k3qY
9dCCPLRxVKrMqW2IB64BGNtDJTHkWuB2ZKYvHge/ro3CzPOiLR5QIvG7yfuLC2VL
9rPYM+dGd1wh6BxVoQVHm5+33uKye25cA0Ccqqs9ZaYjWTmthX48Ayia9rFFD9HJ
VRSrVtquRMzjLzebPnbvS4mbEB/TgIxVRfze3X5QrgfLuT7X1aq4iSErihFWKiFc
8DNJ5ZPhGR1H2PZpgSxYPBmpKjtnwxaLxj1xOT+S2L041B2k0xMIeSNRG8wWiX+5
RFXIsvrH0TeHukh1qgUDuo5Am2X5XPR97Uv0ii9TNa57+PZUgwh7AGO9BRSVXTPb
Dgqr7Es2AD2S1dnu7w5PmtUvoTN9cFJOXVp9EliH7Alz5Ix/Xv8ADQKHyxTG2TDT
pPCuWPfHOGOorNtQ570v9Ur57J+QJTVKLlTg9bvqDCXzBe9/NHFQZwymNIRCDLCR
Mic5KOHw6/X6F8eQ99rSzcY/+UtXPO9E8jjD5XAnjyTKygUIj1WvEVcGDwOf0I+J
MMe2Y2RD73R1lS80X9GKlpJ3njRrRJokHH2Yn10zVYzhjLiP+eDpPXiPxBp3VN2v
FLJOwiRhmgj5BwfWRpcpMnUPrAbN9j5h8KtEsVF0wG0Hz1KkkfG5nTztpazZGpFp
sx7vOczoVSTvLTtV9BuV01U2I6G7JZiEU+vqBF8sqOFjqPol6PnIZ4ZeDD5vx8Q7
dTOJ/U6cuoAAjeXn/assIPbbeTEFXdnhPHDvmtj3PDxTU6jnPr9O4d2VxnHtjZKL
7lvDMlZAcDFBh0EgaBtP1K91wMSmi77uQYnmRYBiwTim1tzZlCFgiZw/epfrJBg2
BIvEs35xUTzmhPta706KDyWTteLdbOEXpnlgpolBxSfjM7urEcR7iIP6erzPdmb3
CPNQFCuK+ciVEnkeWk5U5xYYBeP7jw2qb+bjq2YzGnS64Gwz8bTc73kmWoad2SKp
H6NtxzZdbGTacxRdDJQz76w/Rbxt92TtP+z4tgEPUhZJE4yCBLSp72iOGMiTqgoc
gMuGQmGhwW9ZPeospLR2fGnS2lP7DTF1vaBdirlsG9RRzGWM6HRkB+NfeaK+EPvJ
t+fMbDluQWuFrUY0fb4wNiALZSPE/qTpaRe37fHguI20Y/GGsCnW1JCEnaUwgBG3
oHOJ/WTSgzP6gcRY6Wus4fpbvz7ThpU8QiDDZsoodIgp0W7D3z1ClpsLtp0O/ZP1
CiMjZ/+IOd5Kg06r7b9RWf23cfYr60jSr2IHfpSAZ+tCYErAaL7T6fJcMoFd8t8K
Ck88owxuFeiSRBVmBH51Gch7KroZCv7x2j6haxlxnk9CojcwtmrfgcrUIu90bi60
zO5O79vlc0zbHdrNMrzhs+xhJwCBADNPCrl/lmSJfB4HWA4np+lsVuEYySszglcD
pb+m/OdDMLxWMFfal3UIS4e+YhAdMGUF+BuAXwcCLjU1bqCWtzrHI0bnF0D01axV
CKRUg2Iw7utQTprB17StqxzBEgJCbq4ja3XRxOFsOcGOnZSJHO7rmsW7SMLLt/ki
fhlXIC3RKVXjpHhj0a71MPzz3HHZ1Ig/uYVx4bnMJAxeHXn7HX3sJZwaPAjSUZ29
uXNq5DqbPU+FqBleLanfoB1vWfNC0RXm1DI3SPq/Fbho6nPLyMG/RvZjtuwy/BZy
lA1OMdl8aUD/B5DglQH10suXusxJeFxCYhwWngdw9mweXoJUevSZPLH6z9jV48x5
6EcyFqA7Iby16QMQCeKwXIMQHTkKOD+ByTZFJ1LbH/KBerR+wizwFpTIqelATPct
GvcM3qQYRgHIocdbNjj9jTyVJCPsxKZj8Ep5ughPHK6bHX/y+Ix+ClgO4SnbdDfA
vXotIUVkBQfcrSHXm5vYj0scue2/zJrsmDD2hZgXKQDfvUBtunaClTNi8w9kZJ6r
AUrdeq7Irs83h3fzPAsk/jbJU9Qx2aeXahtI29Zr646TXxlcX7B9Qp/8JAq91X8K
InPWvvpdHPWdEssUn61vHXV3B5tBmyXK5pgb0r1fK8DecuW6727Yaeg8M/mX/3yo
PkxuNngKoVQkpMCzyap4l5mMsZQAn3MPk9hWZUKsc0oyanLThy3spW2b54seRw5a
ja2S7OXosYZs/J99uE1Q6UF6cFz/Y91o07aJIVqTpqRtUqK8YDLDwvtxX/iaar9/
Bp56LA7+HsHL/F6OzGRLn0HZnLBUKMjOeVxgWRcxajdxsU7dAeeeWXES/wa9QETu
yh6klzhCh5v6xk6HoMVJCRkb3cnXSCxwB3NjJ4G+Q/qj2lAzd5clpiw/JMqAsF6/
T2L6KEv2w/tOilYwedFtuPe3pX4gP01UJBfCaZfX27NuCpQ0bmY9y7RIu2xJqzhv
h6DEvgxHkE3i+5KTHT7nClXGH/5/Y2MF3Ti2nRxMMlLZt32b5RuXXuqxqQOapEPm
2defgmZEEmEgHIdZzzuy8wLxjL3kpmbRb77aNHS9jgRNcKy++BxYWvnuvsDaH5eQ
d98bFy3o3o3eWuN+jsatMzpL+GPhrL7aIpBRjsiHV35dYN6AmuhVtithaclDMpyU
Zg48U6M9c6LxTZLcb/0k5xXQ3aLfwl2WAfTou5AAMnqr+w6vEYsFEkPbfyP8v8uy
6eEyZoseEQnP8nJKSDZNhZE1zEUjJKXanqsxBYCgRebxrIJGEqYBJoSO7ajKQPdD
oWK2Jl34KNO9Ib7ppD3omc4YjsYnETn80obwQrZlL9Yhj3jshaZPc9h9pXqn3YJp
+oLx+9bmx4vyqVnWwotEqnZwXXAtkWS/wRAiAcB7KrdHE3KRDSkLY+ti/JrHbwER
yp06OI3ABUPoB7hiim+g3JBGvpWxYDC9sRsHw6uZ3AsjjSoBkdns/on8Ck+nza5B
eTOWt0xaTCACtmLWZ0kNzVptOwIDMTdNhyQp2a0OQK0yeFGNWqcBbbHah6KwWfYI
xdEXPvLvt8YV4GMcOoogK3EBLDJlDJ9qjXF8BKGZEEelbVnH/Tk5oiUywx5VAzAi
/RZq4ymWxv4uh0pWaxYxeRoT7RObuu4arML8Kw3OVoQfJ6OrB8PIZuBOX4Q/fs9M
bwc2K+1MRn2h6N4OVjybWDll4b0BnisLJfuKEJmqvQdWGgMULQkpxbz3Xyrp0Xe2
iGldOoXPCEKSftqyLvFVlxdGyalDFjIQEzVc1UUy1iZTqnxFKWINPgnzGixOfRMI
MK3eKrtWTIMiiB2e5I1ntn7pi+m+LJxyUoz+PJhFbZd4ih8ci4fqWtKoXdr1vL+N
W8ovmPC+Ck/jH7l2UEKXzly9nvG6V1xn4bHj7tcNGbw9HEKrtz/ERellWS+vEa8K
4RhcT6FSQu0WO/36QlpY9fkNFvXFy6vmwWjO4XS+J1UiMljm/PYMdV8gPoYpBinO
0uIzWB6GAEmSNwIi4HLSpH5XF3ZUd0wUFI/J7tO5QX3gxZ2EHHHJk1A3ioCwurqv
CtyKH09Ly5lNYPrGI+ZfC6DG0LjcPmzefMgAUxW5pToFeS6PIbAZEyXGC5kM4cTh
5jKusmaPtUVIPEaLLPu9AUXCnTTKZFCc9aNLfkmJm7/99pOfdxrMCN38L3SSpCbR
b54S1NNoqzxCknWEcVD11qx4UO8nZcbxaeYlTpVwubnlFK+ixkZsZF8QaxpqbnQI
zGkbGk2Q7QkytNFAaV+Slz2CFFfV2QORnwisfNBvVtVWFthmDWLnZv2zNXCCHGdR
1Q/R+abtvc14WaEkDdDnvjbiJR3Y/8em4lU6holclMWndO7VZX3vqVjRenQ4GZ68
n4PR70kGcG1nDFW9aWqxLAfQQHvoWfAJP4bzxXmB2TMvmGl2mRm45XLV+/nsGnPc
GXOBIcIhbZZbhejwkMY3ol0b7/+woh3z74I+ZvLQA2fNs4s6asfc50MHrUWJ+4Z/
BDE10Oiz1zFUkRbXpw7YQGarsgooHppgb9DqJ4dVRb8zdFcpfrjWsfwiIYKpP45M
JyQHX7aL6LtSxRlFizgqXhw2ny0Jf64VntKc6cAoCeZh1pC/OokIzPcONtiyRxKx
OKwp6pvxgj/2k45DapgYXT8MeInoUyR1dEYsbXtpKLm09ZxvcH5d6r71gGBvGjN9
68YXv5obIQLyLXHXUvrLZlPd85x4/Bqhu8oM00Kx155O8dwzwtyCQnC9bHhQjhZ3
xPokbJt/ZgA8sWMdzGXHtDLN6939IfnUlUTdDGTAMsDTnjio+Hrh+FwWDMwunWTV
gPYqrYEpNS4ARygO1mkU9tpuBNfDaZJaaNp0YD5GaTM94pvLP6ebjj8m+wEqi3U/
7YexFLMdUIiRMiWP0x26x+nLLKcv17PtrsBXKqqFjgYukK66DkmXp+G42tFtXm0X
as+rDgDPuI7xRL4gfCXkggD95C2yan5Ui0nqBDvcMvtxY67ZBgh8yDiBtmco4AiJ
FlWIauRZyBP9WBAxrK2MVg==
`pragma protect end_protected
