library verilog;
use verilog.vl_types.all;
entity one_vlg_vec_tst is
end one_vlg_vec_tst;
