// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cQ9ErjwsUiugHkEQqQNmMco/dbP9IYNL2UtGMgWQX6BTo06nw7SX+zwulRhB2CF3
U8xTRY1Jq29qqCnhJ3eVYVEiw3A+9iAF4hKlCkSJqKi4ytdEPHgjRcOZvEGGxjxk
XDJvcg9+igi3t5KMdm3pwjfPFXxlxDr955fid+Jjk9o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26400)
FXbFFD9h7UhlWDUtLJekfKlTzigxe3op2psKw/p9M9yJQp0B4GJ2iJzJ91dTQ0qK
AiUVPKwGjU42qdA8tDNJgUwzxuw/fS+EboE0zDv5njBqZ1H1Eir5IDF2fZshUnDd
SajwWlYkgEZIWlOnk6QdXwRBAw44mFO9zCW30v883cX6OJPTpoo9HDtlIk6SLZ2U
kK9G9QaMhZ74CEs4d4k5VR21pGMiLXL0UXv7BBpHuF6ZtKDnKtEirfBpR6BOJsYn
fcZ2g8p9seQ9FUApn38R2qwO9ALp/Aky7JMIC4oVn1LQrbeIqDSbNKKFmQFtoW7U
uegFiQtkNPjE7e4W1U79h1KIzeBv5cZcK8Nt2l/bFGj7/glgw16TpgwY/0tpKuR4
JmRIHcR5ZUzSw6oeGFZv9R4TqgYcrPHSzblMaoU6xcIEMxaeHD61iqCKIRi0RLDL
AYR21LGTcCkpEdc1uZ/7sd5iRHAOdoaIYVP7e0ACWR0VhIdiNv9f/begGkrYI28a
Ao/pFNyBGssST743xtp3YEJwyV/8wiLUsIuGk7nRtvb3ths7m5nTnb9slqtgT+05
hGySI7WUywJJZPxYigetblF1mglcEjB2h5Web2PraEggyz3G4E2F640eZo4tGny6
xF36yR7dyR96Bvs2FshMF3QLtJMLFwJSs4/iLbrw8J3ig6ywcynuuV7K/2jeSpsU
DV+H1XCM2RDhhZCqoaWT7S/I56jdumBW6bTLFZNsnKZU29K/B8o+0go81TgRHKdF
CgiDfrKr83Sg6qHkkGMflKUBWw3Hy7at0Dut50CWEDFWKBA9nLN5JGDcty+/2HRB
1cSYDlbsWeOXukozOAdd6VpCO/L1Cco//vo2U9RZHmw+OzzvtDgpsErvEMQv37tb
vJf6TVfMarvjZBF3R+Q2IcesIpuuPE8+9yCcwETLP3bV7Dghy3wi0ne1MmlEdrFV
hlAd8U2ZgYGJcdUhGKoOlq/rj0bnEW17H/+oKVpza4ZJqW4BJwodTT/aGdgZIhDW
ksc5yczAXtugVwMLInbTL2DxGihwHPEixyAH5JMAYJpgRBPM+osWkGucmlpROE7e
KhAi/FyYVaUdfhocP3jn38VqDpJ3sL8TEcZz9e/ECX1MPvlmLVzzOr+Y77q4ytzo
hLkCiv2nQXrLL1ohjkCIzVRFACSHRTZnjYqM6p+mbSzgS+ZXlkKByIJYfc6IpoKh
XITUrKZI+xUYCaAL6Xd4k2ipMuTjchhhvl1aL/14VEC4L/aVcH0o7YtDkcTmmnmR
o1x+DQ28FMk99clus2nTAB8kmMWyEWnaUil2AXD/Q6pTPh45UnZWEHET3j27fudn
9IBG5djyvNeoesdpquYsLMyySYQCE96AaEhmdo4ySZq91TIGUQg92IAIb+9s5R8o
SGMUqwB3dMIEfu4nbsgA0UdSjrcs+OuWCAUZio3LHkdwtnl4M3GCtLHovt9HitPG
+Y+UMb6v29Y4gaNDQdQ/hysNlUkBTirAIvJYJeFvqU7DAm5eUraBDSEgMreQBnW4
MhfXsNd40hSPObq2G7ys935pVuj5pj53pN8p0TghQ6OYsVnnB7S49J5PaudxsDXr
nrr6pjxqQxcUpyCmhS6WgBcnlI2suKvCYgbF9LdnPBXQZz0Q0V2LnkQOXdySmUjN
3yugwoCGpnQLVk1us/m/sM4TrOrs7UqgbYlEX1/2HB8H2aKfjSvxLUD4OIak9rek
ac5ZwSMgiJ1jGCgPqZmOOvXm1OoBfKcZT2W/k4r7rIi6hs9GtVgXzFPbSHw1d4E8
grzkq712T2Nml1/2GdN3h9LcPKqLFTJyiMPqO7xLmxhRCMNMsIzRfly9Oj72hJuk
LahKWIvxTM9d28r3yu+ytlNKj/vNTHLvYJOKKC6N4xcZF/tqKlJsnBgHxfZndnis
pqsfC0qRtmkh21fh4QZtQ2Kh/rq9cOeNw42BcYghsR5POoGAeJcBcPC3+xZ/HRq8
nshFuvE+TL7TpAwl3IQzAY1lt76qzkRUfd2YqTe8L47WPgI7/oYKxQhbxl7q6HwS
0xu4i2vCzctrgqvecdsbF0Tnjpj3moEOiJ7zK9pFDi6t6xED/Gr2qOGYVp0z82Q1
4KxIMaDRqEnrm/0olWX0G8bRHtrJz0ZOPAUUzHBThkitXhVhL6p/UdJLhWCR0tKW
HUjp92d+q+B2woBKSs0Q7JWJk/nnXs/puSRZy+y+0+U+1Ho8RXZdVljak/tOwghU
97tsvEMqbIk6n0ZjDQTBMlzkwOySi0Kow2tLbhdbDCck4A/e3NTIFX7V0oAMO4Nq
ba8IV2JKRcqwCLVP4GRRO7teoLJ99ZuaXrlo6RlalxJsMB5DpJFiYGs6nVpAA5OF
y6/BAYgRFRdsB40hbrWmelipCsQ7fs5A4TNbp0H7eoODAcqW/cYeS9YK2QW2vUfq
gSatEpJ5UCgpk7BioKeQ/5UT4FEvxdwBiqyuJv8JO7qck6noGzBkONPuBCsxpEnl
c1qtyjQKCS3sCJCQ4HOSf7vdgQl7BVY0OuTjFqDb7t47SduThkQ+OeccxlRLvj3U
+J+GSo/vBiapK/G0vTAM93BIfzyvffUOsfFkDquqpwhVMy1yn82e1ANrs4phJN+q
POwj+qTFkcKOztoLBxq6tqIw10o2V6rXPPWsaUe7kHm5eBYH86xfAGozdrE/XajA
TEhYIV5Mr77K7pCwGJeKd1HQdtaNhMAosadnmi1q+M/nr8tcmdYTvdWpKFe/yze9
rSVTGUlepwOHKESxhJePxcqsih5UAZSU/SQ0K40bscj4z4znWAMydpVhaBkZ9iPW
mHXMqDLLsDJED3jxY7i2J76zWKNku5svfRQWswdBMig/rkK/49feB5f2EtVo5V6N
NuFpdfUk+lViWd6Hy7pP5qDM5GWDSeqsEHW6LggOgZX87GPZoLSyn8VSDJXnTmId
AK7lThaiIQ3crJOsfv8nUNGcgYkPcgvxx8c1/6H6ItKAbuaAA9KTP/WpVwuei20l
ARjekrxuBFC9V9YYdT3JZFK2JNHPV44xxcwdStlFyWM90+/boNDAB+Qk5A07FiBs
R/xaxLgrQIGUjR2nV6HCFooOEedVSCbs0wpaa4g3hZ5CQbRTURmwWGGwZ6cXFzyS
HfmyoREnmli4RSRbu2IcDpjP2frKqBGSi72dYKZfVI14JO3Sa8I5G7n9LnEA2jl6
ZuWk7LOZoOP74Xa+6LOLa5Gs44dHOZc32Pr3VGVktVeCnoR3cCl5PMO4r4CV3qwd
6UUWeZrR5U10iwKLUwAJl/2glSbHxjVoe5bxiPYJtGrEdBe7/tyM9kl8Zc33FvsB
kkTvRLh21v4GVIu3f9kRQw3hxpDI9f+z1zCIQlmZ4egVeJaLZlidmraRPbItS8es
rD3XolLmpkra8MVTc35We0nRkHlRRIirklfBMxHPDnzlFR5oaoV882Q06oDh5NvT
yLIIDYOGk8EcdWjdKLuicsKnBxYEWWxKzFXsqTK9Yvygoux8vCs6hk+bXmfZ0SqR
54xIZ58fwt9+gtQCP5we0b7UQpz2MjuSxdtxsAaegRt6Gy9HUHBzyAiMS16/znUY
0/VFTg8GfRv0rXJnvgiQU5C65PrrypZ8cJkyMsblc1HjX9adodZlQBrELurMmC/C
CQC3eJZg/plExipoaDdZYou1Um5SinRBkBdO8mWVqU/PFliD84K0F+820HzWvfsa
0hJtYtscOp8e+yXq6NhXgjucvdtv4uweVbBZKnLlsbeaGqemB+McrgPhN9jzRYf2
SxprLo45n5qZox/BcQvRGZREc1QL4dXZAJhM02y3eFsQo1G5Ffo8qPUOi7HXiN++
zVCrtVTdAUn9sE/7iNC6hgRiVx20B+lMiWJ8Y3enVhn5DhslG2TF9mkQWvObYtqp
H3VuypXjsLf2FxXO0bIzUrJa9+lQv+pe8Lg+YAPEQp6+G8i3KqhZb/iOf3ZOcu1d
9uttURJOfoTNu2XT+gYkSI6taFWL58bQoxcD2beUwOT3uqKsak2psN/dIHe+44cX
09LNCuQJ3YX6cQON/FH7ox0HRsXSmhG6+9zSBVgNRtyAVcEQfD9HywETaZ2TcRcE
3Bdmx3KW3VM1yA5EsJ455kXfxW4Sepi7YGU+Nt5nfurmdKHaDHCyyBKBzmJICn2M
QnWzEmlwSIhDXlzEThQBezKEpThJmUWvJ6BsQKIOX5Mhx0AYWOASFmwtxijR5kRC
yBcVeqdJHHD2jHKlz/kwDf/ob7mwGnRwXIs0qjzQ0gLTtaYmewZnZhtu7+Q1pK+d
WsLL9zhFJwXT+z8h69gCb1dqXre7Zh6FZvFKe6gMaMBmIhv4LM2v2DhgAQvrIROa
nhrOr8eKcAqXSYeFaGrDM0Kenunl3yetkKEkbsUlPDlvJxoaPHsg+Lm9Qvh6nCfa
5UnK4CUXVk69n8chzIJsvevtNtFvtptUQubdSWoiOOaHvVvGLTD1+sarKt5hmduv
HXnw2VXwq/p6R7J5Ywmh8h91IZCNyc15B4RUy4O6kO9zq8o3J+fihzlGIFLjIHew
cB5fATJgtMhQfrpZSdREDlmJCqu+j2oXOlsZnp54K3tnggAGNMnzwmPB+VGt+XAO
qjCHvJfdZTmG1Ig8ThfABlCtjB/1Q2IoIY0KwgXgBEUFhj5GpnrA+Fwr72M4mWE3
6ZbNsjTz37yOaPI3HuvNg+YWp5zN07t0JeKzWcgA6hqSrijrCWNZvotRjS6hIpHV
UxJ7XNEcs0nZeuMKgobBh27t5Y4YEQUrenlCQX2ZwIFLJ66bCGz8NbxMR0yfNXFj
18Lms/Of73J0LHRNK9fOTz6qW+9sSfod5pVzYJwGvQl6oCE9nGJXjkIRZ3WRGHQI
dTNf81fx+Ksd3TX1+rc3H5ceMiOl/GrxPFjcfElaxT3zpF+4oV4rvbxNaM1vzo5g
q6hfA7PctSmlSEUTTMfftmDyHqFXKMgtqtESj/Q4/uiCcGb+7Zt13nhU3CNWGBvi
aKkWw+8X4kDSw8ff+Goz/j7HI1t+0GJgBG2TxPZ9YgK/Zo5W8TYh3/+IszCv8rBB
5UBe4jPuk8Va6hYzjahxiuiUNa65fdkSoy5/yDC1ZhiuW5ScqEY7UCpA7kJzhmsx
7Khr81acuo3HfvXZA9Rxhcv8YGL0ZjAJihLh4sX1ACpVOqCZmuHaKvzkso4eWorW
r9BjljI1GoilhMFroDyqXpkRK4Ola1aXFvK1onn8khETcJN4fFOIcB/eMYd55SU1
E4woPZRfMN/mKdDQLEyfloT06ElZtqeiXWtfc/6bKEEXVqgmywbQquiabTyW1z6Q
pMb9lnhD4is/+0EKtsdasqDFgbMij6l0QZX8VHejhrICujbbndZAg2GOwe7Pcd2r
D6tctm7pe7RazocmRx7Dl3jN1ZYHwUGv47mJpXUPsfUIUlcqHcTO/Y9QscxjEL+E
fcziPPpWWBQYsXnPqqolarD3ukzdguQg/Kucf/9OSGF0OW3yRgTX+sUWD9ZnTG3v
jAebjv14QeyM1HBTjfmbfnctBKhrP89zbiXN0zp6XuEuks3tC7MyW6V7IZM0eq2e
nb+9wZbvXvzdr7uE4TPqffY/JpyUVMih6Qhvm54QzLPTEw6rCBeuc2bJ2HCLG+Rl
5n/TM17onFU0VCpgZ7Sea8yZSjAmTD3N22rUhI7jbmOnaVmA8N+OyqB7YsbYW0WZ
8MiAI8K4M9HNiHaYURr0bqSabfmA9EDiHl98yS72p2in/Ik1grgE5AYMij7SkOBU
/r2KbAV1j3XrzB/uzdQKJODmBdpy+JP3jXbR+NxsabWMD7s+oTYV7KEGvCLIYYZd
T9MPFbhR1zRyIFVWjMyFeo+CmdUeIk57r4gf6+7+5fRm4I8u1D+nPxbuAvsBBC4q
kLL734Rp5UjDgwGCwwXtfa8DFIEcbDOkvbOya2IVKuolD0P76u8Y5DHu8OcLFAZT
1xEIcKLy+Z9yVhWXUSL5QWh4BSHrN4pzAC6zIfmtEa/z36OJ7wFEsHhkx/d926iB
ra9cxiB7j1pqEFf2oiwg2o6LwMgnQ9+mKvdWuBS+IRo7JPy8zLVx35nGsC8qlgdN
ks31H+wN+miMIVR/hUYvWU8IQqNIGMzHeBw5kLL6CseDjvRK06Yu9TfifqcugdH9
fILBTx642c/pexnGV0nOnoJUVZen/MCm/o+eNarR51wEheth/dVAHx38yQtZy8bk
PMVUcyJ3u2ZPIaqVYZ5mcBhd1k8Bm63NOHY6L5u1ANRyEWoW9M4PW0XNUXmAlcBx
mQ0NNh4/KiYuQEe0h/Sk9vPTW3N8NSgKaJ1tLIvTWpUs4TMzrqOjuC/mzyGWUppE
SM4juWr7fN2UXQuurQlBLOcM8xPEkVL/+GwScU0tSrbLTHizLnNja8rlj59PyXMj
Dfb7znWB+S4nx1Sx3LG2AalsMCxg/h5uUhk6URHBhE7LbXxxk+ARkf/l3pBTJgOj
t7FacVHaxgIseiIHPdFzSQybfrKYYC4084aweOvaQ/qzX4D/Kp4hl5qD/4WlFIVN
OucNoOf4qjAjKugy+TF0z5fMwG+nyKhMbRtIxkh0JDFAwM4qYGMpcpHhQv2eyEcE
0opkcsk1dpgpXNSbeh2wkN/dsNE0dUKcFIUPVSru6MVdZKilZr/eX1eKc6IUoBXI
3LA6lgDdGXpqYZvtNZmUA5Lk3AIYb8f9aolEcZbNd3fWJnqmaXHgWQFrosvh6pK3
BXP8HE667sIOROLNRTYt0QVT0i8DT5nwB8S5bFPXrbcd13BiLjwWysNJbkl23I+J
ULUkCPP68BicGOTWtf7ogkPhmh6dh8Fa+a2eNMWoNozesKAPHee0nGMGDZwvpXf0
xjmbbUmsVAxGqI1h1x3VudOPdS8WswIHMGkTkaD75wUwOW/9toqHhcfal0++Hr7U
2jbvjavPKv7BwGYZ5bRTPsm8ZmCeZip5kbCDiRs5WAPz8JqO6RQfUl/0ProoMSwd
H+XD4qd2f8tSYvNcFLojbfARM3yZMkTu03C7F6d8cDdyNRnCuu5/5s9jp0Zbb7Mr
uzpZGSFQWMmdxxOXNNJo/v3vW9eGQnjiHfmaKsbVnHrqYfkomXPqsLhPomWJ8j32
niLGFTSXyOIawusulHB5b707yhHydEg2ermBMhXh91YPl1tG3teBsdxzWBFd6kPB
q8TZE0JBmRkJmN5Yiyww2/7jipzlZTKsKVPI8VlEssTSiGmuFqZCwxOKGGUVcSJ7
iIYvtWiv2N/TePg18WFEwGSrJSmdBFWcHtl/s/8OSQnxTGDMmdLU45dZEjGd16mx
8jUPZRuuMvzLZOh0bbmqYa3RimyZyQ94feSaalgmjAE4mKF/Pe60oIjSTkesX9rQ
oM2ul8kffaVPLHdP5uJKqBbFVNPNoLGEyWjpSIJk+/g6REwtue3WzkaEMj2IqlAD
GzKfQS0Bx8mt7rw1Km/rAZAmJ7b1Y8FXKRA3Uf/LLJH+GELYB2yuxkXDLeiXao7c
chbPOlqcwthvlF+Cep7pjWhaY5yGnjvi0+3DDbXT0hZnaHzN8U9uQvdCCp038+cD
yuIHlbfJ3mhYIRJyDcZXd+zb1yGIzv6DgRPkTGc5PXZVq6XOLRklOUsOs65ZoUvV
sekXqy04Sfo/qcVLa1WzM6zxRCf3dR0h2CUDomF0xee9vJbgWn9LLTbNOnYebTIP
KBL40XsOlWVrJSwWiga0WaA4p/7GIYWPtJTSrN54HawDcIS18861KQDVdlal12pW
dNf9YRZCOJj9B5eKI9PkW7tb1mG15+AxmRDlIAt8/mzVPZ8nQXQDjIZQk1b99L6z
Yq01DcXWfXHyBnpBW4rH+svDID2G+bqHIOcYE7RKat8SJVj/TUcCCRBJydvvuW/O
8u5HLKoeaFDCs2zWVSZFPI+OOOmzAgAvyvL6ZH8ykyK+ntx/aw6vUfuj7az1vq5z
Wa/0EYC2YjOKe79a/AlK8RotsKqbUEpQfePPPgkUjUdmGrXgCn0qpjtfBYjPBAdE
DMbnlFMlH1bMbk4jCuPUB2N1PVHVCt8fE/BwugbH83NYWaDlKCVVwjmfHVtgc+Zi
6B4LfpVte3hVKyhvdQNjNekNszEbzKaZLX4jSCMEXd71VL7GQoua71+pFx6kJaEJ
XmsDw8fbVleowaYOqa3u4Io+lmvT8uZftnp3XJpOGWJil1W+SH8MLZpBUA8461KN
nYiDExgLaQRKyRG/knD54rNkaW8kpxl0yCr/1pHdqTVMvBoC4DQGDOXQ54L4CMmA
fWCSWmRMQ1cfR2fVDdStWGmcuaiOULQpXmdEkNSUt8WhGXsbezmDQEKPmKuP0S5j
HkIaRPvZv8QPtqclhRONcpcoJv2kxofE+NApawKppqus/E527eW2o76HEQBWrsch
uyx3f2UiCox5ADG746G9PYEXqd1yF6T8VJEGkOdxfxzYUUfeSLDGZvMpzere9+1C
veuyt8e0WZRM0mXdxTC9YncSeD6uK3jOXajiOA6oTLrpdG4ZntS2q4eQpupwTjfw
ArNT0u6JRaKCvvZYx/at/mBZ8UYaATNEXiGrA8w6k4LY+pbIgcPL0viB3zeqd5ra
9JWLVkWxbd7sxbmgnui0cmKtFjb+NkgZmXHfBe7T4L92X5TyYLIwkCnLSyPPn0W4
dTR8VpucIs8fd0otFS2dOITt4CWCIJ5qNNEO48tN2ar+HR6lhVRQ2MMA6URHcYfB
ZXMCasepNiJsmNPJcgIhZvlFEBVSHtsNbYUHNGknInrXxryZt2N4f/OWFmuo4pma
PzdjM8aCDr6rNqw7oxnQHC3f92slQrDqpM3HX2z3YljDGQ4cNa5tp/k8aF5TQFDj
lSWLsD2qGdQDpz0bxOmdcF+/Y5QuI+rhUGVT/hF53Lfa5igbQ4sid4SSOLPpgOAL
J2vO0unf5z+n+FL07VKG0k1kv9Tv6xeUVixEyKGjtWTEitWGXmui0BEIwi922iEG
p4rrzsJpunIXeH90Jp4mKR0IfcImuS+Ona7LTrAPt9U4phbcIIhXUjARluUfVpo9
ZAfQc1jaiKj2cfr8RpLThA/n8FNe9WB+eaAjEoFcv8QOkQwWdakhrrOWUhlRt1FL
U54YMDl/KsLYYqpe3KbkpZ6KEXjenlfFbQJTCX5jElZ4cUpgC9ZMhbNV3Jfi+dav
6kO/qhCiKKnlqkgCYNX3ftp1/RIOR79l55IYen2h5aq73KtN+TCmJpaHdeJMCzr5
aAVqwxDj1l5Ahklc6GHkL/LLhxod1dyiscQtbbA9b0UmPyFjNMH5msuLlpaIgy82
yXYiKlxmLCSTcxFhWeyec8Sz5Qd6xFm7g6cKvJfC7VEnTosZw/wdhHo4pdaS/rlo
9C8f+QUgGAg+gpy5Eu8kOO8g2yCaP5zTab9V4De58w8+NHpOvYFvVqy50m0ciExU
zKNFCqorBSAq75rWgoUA4Zi6XWnv1EfiGzURsrtU6zHeRTAsTI84mPR3Q/ujD3dv
MEyhMB4na96iULxaguy6ncgMRTKFZ/zee1f6OGn4xrapzalxJe3WvIEIRAhxTUN6
t8prSskWCtedumNyLgL33cRGNvAn4WWhFlV4p+epMJNAYHhvVH+PuYjbs6AOuXQV
G/0UaGxn7y4iWk+l8mMHAfPA5f74KEoVtaB/f4DJlY5rkSyECzOwEnz/7TrwovLg
NRI4fGpwDJpWU6EURpu/ZLK8EufSydBhTcoJzMzRr4jVTgTcJCjLvjxBfcp/wLS6
Oo3pY9MWF/E1KUh78qRwQRrfXevl0IgbswMW3Gimh+avp83x8vMBRsTE7K90oke5
A2CFTTlGwz8YbpjGdd3lbt4nx/d1FGnZCymclwOmlboeenpTnNE836/ABKCu0bcK
FqHe34mqQmCNXSHoNiKG6H2ad8r6a792W+ZkG4WXKde8Frful06Y3gx6zQ+zBbrL
fP49ksGgJzcmpKAZ1XWAZKYkFOllewmPFCYM4lanoYrM8PDYpKxycjnaYggzlcpd
+EjfEJGVc/k561X0OVLwtSb4dCDl0l/888RgzRx9nO5++CZpewmCdfwxTxGdME9a
GXQ7PB1jcjgAWOxIuThEeERv/C2NameVzRq5ljJ7npi1cKN+1vPqD9ohLuy+si6E
2zu9BF4WxqDWA4YDupaM17l/BbAThvxw1UF3m5DzWqFciPJg7P1DndqCGGjPFZn3
S6HhPz2qjhfkuRdMrIxuCc5lR+xrNQXqRMi+Hw7Y7WyIzZmHFCibxO71yCQwkWDc
kwqrPJ7vmxHnHPu7QNZ5yuXlkFBO1zQFm+rOKuB3rwG75ss/1xsp9EKOUNCt40Xs
VrFriIta7ZeiCtHS4t13DYTDynGJLKAWNF1/E9pxhLFIJF3PzlYDmRADsE9N8835
4SLkqqkDbq4Zqab13TiwMCXPDvqxkk03t5kwgBhVE5oS64Mh4Y21RS8XUCpbMYRQ
JamFKk236yKQZl3eGxEf1d5YAslEZI4wBAPpWqpK5GrOwhkzFyOFwGBcp+VGFBg+
s3AVbAjXaypSe2UsUieHVZmEx3UO9j27iU+hyUoER4qP/HbCahhNll/jkSdLGZO3
SbTnY325jnr1YXMLGdtWYvFeJrK6A6WAiKzFMjyQucQFYo2T63V69/dNZ2btIrEm
unNcmXK51mLc+UYcZJCbpbhvtIwkLjdgFc6u/faIWcKLIidei+bz98JsAWDZDPly
z4y4Me66iWHvTcMMsQRRRIqThS+aIYnx1kVCcPO51vrCE3jmNh+nmM2Eyp66GO7q
g4pAeNOAwcPc3PX8N93CX4HAV6SIU538KFR/cos8LmHYvwZ21KAJ1j734+zuaAcr
bCmrrtQPIqMMjJwMfnXr1Oln58Lp0kIRQ2liJf96b72ddWcL5RU7GG3+brh4ukMm
Hy3bm91+e5EZUhcsXU3HAUr2lEnB4Zg5c081ur7fhEr+AuOAUiiwxNtjGfX6lnsW
HNVAOxwc3S8Y54PyrZdMyjBBDTrVNtsY/6E4X2/7srrLqp9qC4wCP/66rL58JuZa
nMjtQLRSJKX/QXqucI96sT9VGaM5tmlYdyO76kh8x5nRADqgMWmwDRdNmzpBf0C6
ejBBNA5/UNUam2OKK2wCxaShSfU5zlEJFNTTmArM0sVlqy3lg2DmQdc8p3TyWFn7
zLwc9FBUhStUju/17Il9dtioEUVRGqiYIperydK9FTIfocOemyxzv/geLHk43blz
qE7r06IJ/74cZC3Bcb6cuebAVhhPKbaSeXVm2fDiv8+GFcJ043yjEJ45CO1i2i20
yF8+GxAl/xQTAf/UcWpsR8VDu+x7zs6k7h1lIFxNWL3LaBRGEGFHPD3rBmmwTS5j
A1GO51CZNiMXCcYd5av2npbya2Aha/ccRwCSQgzUdphcZpRjdbu431+LRKfkroge
VJS6utJgCPrF5dMxRYNwY1MuRPbNGZ9sW2z9uMV8SKREcX1tQo42l3Be4GrO45Po
F/iwNexCALeoucRT5TLo8fuOnG9cc+YtnV4NMWdrllvrbyOUK3ruXSFTXNEbPW4i
X/t2Dtb71mRSKOq3rSD7uC2/ioLVt7MtZqqHqYJC12VS5pDLKL7AO3F6i5tOSfs9
bjQrDeIFKtuyumWcQZc0jJB4FMlAeRsTw3UrKWmTVy/9DyWGcf1wrp7zQeqiBZQx
ksRC0R39c2+RDQVyoDaotc5OCKQ5E98fsqr1+OccuI8+qlPwQxKodYJVGwlWwnmc
x2fH37qhKjWT+/A3Ua+dEvuFfoeE16pKIGDddw8z0skZu0D+lpDpv5ixQWZK4kWr
HCg5iUUENY1WethMAv/3gXKui145gZ1gthZTqPgjXxyYqJ/8TxxMpgmVOKUyUZ2u
tLUX6/1fgsB3U2tK/nzKWOHnY9EdaVjAyIXbiIA71wIflsk05lwRc+9PSx/KgSqA
kqK3XGHfCxM/zUsGgiHgFefHnyK/xdo2I+Fuh1f05bvi9+DHgvd08aUc6Ic61s8c
yfyZu3MAsLe/ecChFkAR8HwmL9yxHtmatMNLWo4FyILfVTL602lIAkfDkh6ErVn3
lpNMhW6tpcX4wkz2h86w5nBNKhBclQTpYDq/U29RO2W3e9TyYRFOk+VtAbVN2w1M
20SGroh0XB/9kIcqHrVV99bYQ5AchiuNKM0kvjB+wJiYPdx1uRZudqUgvPhplUAT
RHSMVhPpO3vZcF9yd1xx6sANfbptWiOBtk2pb+T8RIChm77WCHg57PS7Bd09lVU5
HrVvvDqXUs2wGTPQRWE2jjSrpQH6VQ5dEDb/lqkWFWfhNDkNNiXPH/weMZ3gL3bX
iZtkOby7bLCumGhBs78un/25GhNFroZ1tiatbrX+fMttw74h/NH4FDJA/1ev5I0s
IDTcJvWamSu5UQ8YD3Z4Y4ScNifrUGN2huoVMqonXT+PxQdXdHF0mTlpaNbgARVW
UTFi/vQ4Io7Fe2IWdnJ3tz4StAeYrVPB+md5r38LWwjxcnre7STsrPAir+RqHMAY
R2IVRJjGmrxQdyqrtUpN6XSq8EIGSAas6twAIyGo8Chn5WdfPAyF6lJsoEuHwr+2
Cy2fFyVFM9WdDZV1Abv5IErKM4Em1zEJi3+ER7B8vqDxwoPu1qHg081k0SQi7Roz
KtgaSHfviYxO+c0z21jCrHDh5eCW3kU3WYep3Px7ccQlTHveWcNlarXuO23C5Fxw
pp8w/xC3mR7H4LoQ8JWte2HsarTWpgA1Dy0JbqdQ23CE22ZYAXAithpByvHnDQ+p
YovMbqwYQtz47Exq2DxgRnS2WPEu6M4gE5EX3yaoF0gqDBDOG1uekavlusstYBs6
Vh+dSL/yNzmPiIbwt4IXeW/aXArmkFxykgsL+2eOnOM8sD6theqw1gQYix+di853
j2OFLptaZKhYH47Kj3aXC1f5pvbm4Ybhwt2FfiyqZgR5km5JJLog2RhL612NQ3iJ
sUe55oAvpl0Tx4D/HIlDq/Wrbu5GDSYVTMpKNireqGa36QUnR8cypCozyX2bxeN9
/JP5VHCbUlO4xSgMxqViwA41M6fKevYdejRCJbihz4nU5lbDT7fxbw1+WSLrxcAf
l72xQpVGJzu0dDNuBIdTBK73JWx6r6lEAJqgsLim+Jhycvksen30WFMnfkA6tVwj
SS/agThBNOyBKsRIbPyNTqLx0V0CXklTfibXjmUkX7/EuDj0pJHjmTqAD9RSLDtG
xACQAif7bs8H06sxiVrk6sm34DZEJT/9nzuf15l6iwD2XBH9gcbP0JwOibM/P3X0
5SbmUj5nQsKCeOO7wltm/wvUgcpCxhJ3je9xIaSuua4fHTt9tGB+ZCuDR8OWLs7N
nwoj4IGHd/cswOFR/J4URLlqAmned3il75V1mM21O5VZ34o3asnYFDs1XiI+asR1
vrkGsiSfbLGRw3hhpdkOoo5oQrcBVT1ccKvWYVpvNdPks83houWtyD4oXttk95zj
LZdU/LqDKYNppiwAgfHUMLtfqWLynpYCVyOvjMaDB1SFL40E9s+YEUOZIGa2sKKM
cCSDGaJ6NWakXTIvOcIKjXV0RXD3XLbTEwF8NB1/JR2JafF8+ex2h1vrQ0hHaxel
RJ65zYJ9ZPNwi6JkhA5FrgBlM3WA/Dcd8xtDLZWbWAp251FXh9T1+7MeMDGwvCf3
WjcAHV71z06TWpB+I/F8iuJKcyNrh4qEF8Zeq/OLnM8ZB+5OU3icCQKZpf6tDCwP
WFzEmOeDKpl3jsCUno2r/Q0r3d0aaDA8LTA+wZ8Feq8H0iz7ufIHTOiTW+adfFez
JLB1G4WQjLXiEzj+fx5H4YZslJd79ellg5bbdNlvP5MceQpYpHQ2/7zfbg1q6suh
7cSC3EC+Y7275Tzne5wAFF7F9Q/wTvI4B0lfOhpgLAKalnPF/3UTg/DwFzB0LVvq
sH5Bu4cSFOK+JjbEk82kC8aGKgKfptl9fxeIBjObnh7LESKOwyaNBQmOHm6/j01x
GCfD1E24/geEu/2dkx9/mtnHUFUlqscZ09l3dyWuzdJNu8wPS8+tcPnpBAQTE99e
eiVIulJCpS6p57rwhhNaCfFyCFiq3sxk9+YRuxnKXvdNOO94DX5YXyuV9yKweUmj
0pMvkeZOqq0B2hAc4ArdM8d3eqdtqVfZ9ceavvnmNEU/9BNBmqRvlat8HKAXxK7C
zUY89MitxPahrucvcHlzan69VahYBN5Jh7RJjL02o9mFWdRjRumL2RoRMwAj2Zb7
vvnFBOar1N0sF+pUx1bU2906keGIBARIBSACYu65xomp7cv3SvaZVoooWabTpKEu
A0ZKLqNDF9VsLe4Dlnhly/6JL56rIt7cNeIWX1Tdvy7gKtyAPcZfpMcbLbYHfTqW
dBm/Z3Mx8vpZgHFgxfOLQTmmi/d5q4cP6yA/ehwflAguEGDkOl4T6YFg5ZmeIpy3
CW1lNTfahaHX109MCsMkLcMpCq8E6bpvZqjjAVDzItMHqAtegW7MUIzoZ1oeJSB8
AVszgwdrBuw+5rO1sJAmr3nk3UbPWrrlG4TmrjCO0ZO6j1WGRvotks4jYApR4Stc
S/sgv6a/+mU/f0IwC9w4qIM05yzlgEemsNuhOEGdqEutG0QGIkIqJb2VFBLRk9Rj
ljuznlOuXYmQgm9IEppwaniXq7mTcxUun3e+mzi89+Ck4ZkFiEJuUqYLR6tOPFpE
LJKfGRgT+H2bAOeUyvyO4C1kSERFWzx+4CKljxXbnaQl0556vgqcc7g43UdWHiZR
qeb9/GBgfVCOIMKqkdNvwJGJXnclAIwEwMc7qDskUDdY8e+rdr5u3z8CpcMmO9wb
DVE1H8t0fGVc/R65ubpuaZVS7z7sACFDYIliLDgf7x5q3adICHtBcuGDBGEFTtbz
pDkQMgC92SLvNN028lqN+LFFYp3YGRJAVWGvHDDXUsnZPt7hgMcbzuC45IdKzY0P
REaPvHaPutgCBmq66LKnB3ubqONdUz/v6QQwnn4Ii9T1QcEZ+/1VJMC0TmzRxeGt
Du7wlgyt5CE80+mBo64MhbJFTtSx+48iHAeiLEy2WtUnBwNBVqXmNu4FMww+TVuX
0nLFiDsxW5qKUEx3FeBz4pL/ycSJcgsOIttp/LlUwkncdAW2rAVGjSBcDbwUUwnb
QNA0LJde/7rYVskTYSNGWaVzkDZfsUQndReicxr9vIC8vvEAPV0lHXwA3AxghJkN
2wjdk8iT9FiD6qSlvY60afSF5JRgdSR/Orzv2Hyh6G3rd2XFtm7G5f3481lnGsC3
JqF2m5NQrhc8ad/mSFy/Xyz2pHOJ7ML74QQnV21PNNxA5Rx7uhI66g+KOJc0r0Jr
eznCV6YPQ0LANNoLoTLkgRv3/SbjpNVsORN8qzhN0hHFvmDOodyNyONCodKaaJ7K
pTn/J+ySTHtrQaD90LLDJvTxHVpP0wj8s+s4OpvMHTg9j3+4e8oVNP3O5A1BbIN4
NOXgYTyCStjC3qqNJPhGEjgI52AlQDoPaVKqVPzb7nkYFhsi3jCRqeZL6EE5wUei
r7NOeIWj33Ly0/IZxw7yMKFG4Ye6hSa2E7AqHZqYEdTYldZJnICAsVazb+ey3hHO
eaU1JUCRxlnxPXDrU09uQK+tNT3xT4YBJi3Z64ArfC9Sc8rzKwyynOqvZIEvUhBM
IElP7XOrLVQbKqE9NaLRSUnwXYVohKZns9ufguxv9htYH+Tx0QhNqLDWHr5Kodte
luVGRYva4hVnjMBl8lg7Yn5Zn8E5LSdGttVm0b5PXN5Yifg+8ZfxHKQw7zRxQVlN
oPQZtcn9AMFbadHh0pZsQBveFkYBQ1lf6yh/3Csu3BhjKXwlO6LI/nMdkc3OZDTk
cmfBFzGTFqztzWWPyDnZ+/zk7h3yeT4q4A8OZKFmH/Gqw4SX7KbcIqa1Z9rimyLw
c+B/bmPV1RU10PM6pqokncLlo7gGkpADMzdtyCcwLflcmlp63nR7W+M6o6P/yzzC
0qQ2QKWLBcR7BGdlhSMGxT7DadlzHozM5lqg6rWCoGdBP5I7aKN1Z2QzHzWSJt/a
8l9AnzPyAWAWLweHJfOqfJNQqgT0NjkFkj/+bvhrjEzZZm/Iy4ZP3u7m9rh2dX7Y
K42iYxddkMUVs9cZjIDqzX+C9JlUj9+oKzT/O1q1cGweUN9px6UC1JjbiFK9HAGz
mhp8KZ4yRGSSBc2Xsl05Ajb5aP1oo6KgoTZTEGWcTPCO6yWbcUfmkn0nFtonYACi
cVwKOaHLfHW9LEWB73Q1zMY3GtyLX4jarOlORGy5CX8OByszqHypcL4AjTGHu6Oo
u2z9B1ienW08gTGBhJ34hda6yqO/k3JPyvzawW2IPK9QMrI1RY1iJcNTej/jc8NB
9mej3DQpHnaNy5YYLYeaWMfCs31wfVGsVzW28jx2ObiVsxFiwGvUJEF1J82pfKF4
Z1dOtuDKfv32Z84R6RGQaa2AzFZIFKWQ71nZ5fsGWwbgpChpbEcR6JuqT5v961f1
X97EUf3iNzVN8/Bgi9zwl2WeD+XOENnxNMsfNL4NmCgwcBrOJyUEp9a+8L4IhV4F
qbXWt1ML2fvhNpvTlVxMhinGmolkeYwesYWlghTtSwwdic9GmbDankUiiQrBP9Cy
OSBLNVLVcCaucE+X7fSXJqHKMLF6cNJTYrrjCfL1zCKeTMdHUx38qQnxuIoFPJIu
ou29oT8M1SmGYN/0Dw1MEKPaZmzYrRvoUIXLcbrSsSw5VN+AFyyVl4hxk9GwcATV
dchEg/z5awrS1vSVcjAbywOyqN4XmcHBq2EyQxlW3TwLgC4sfpg6wM53RKiLjNan
9Kb2kCzleBwVQ9QoIYmWdQIpU9ernmdqsqBr7Hg5Ywp1U8eBPeonrTndTLCveE+3
zQGRMwEp1A0XKxD3AVJxXeF17oou/235JYtD3lzk7XDdhzRiCfXnRDK8ax45334u
q4F9gzQICtGtkYjRG8jNdjcpQL3nN91Um26V8MF6toYNvHoqVvlkGQK6tv7mlX7c
tuJZnXBVoLobIuZ0RjoQSlJVOx96wqB0mjTxD2Ns2X+VgWax/ezclQ0x6eEY7/3F
LKSdBypGvJlD5FRHh3Upa24myggpmNv0WPHDpiBCAwujKOpSdCeZ3yGojmcWqS+a
KKn0FTLw+rPHkUQMqdVrL/IF+EIbGGdN142uyBjA8wXfFxZSy8X79kUm/waH38m0
tYYEXfsOmae2rZexGaMUGA3cohE+z6q9mCnPqiV3+GfiXEP5JzfATB9zrScgKDAy
F+/C6FLn5BT1uTwteoYeeReGfO4oxAY6JfUUGuU7RXvzJrteIpv06BBtYZwz9O81
SMx7+Rk1TJjtYOWp8DAZFAAXVxIULLBYQ/eLUiy3Q+IdZHwiwD1jV83GBdL4pVuW
lRufkpX5p/L+ZCGQJN1jwI7RwZyK7BFIuAoLc6iNJc5cgsEgjr4zE7rWG8rKDreG
sj6rWny0gY8SZpu9jn5z/CIsrHUq6GlxYod4gpITGDvOqdB/YTOnlu4eNz0aAeOj
A0v29eY4ppSPtiKmJ5PPcHPo51ZRDatFHeBEaBYX0O0nrLJp2JoIIZii8DlVjjQP
2IABPjlGmTYBqDtD0CiySbV6Z96eOlSA2upGVh6mA0CK+7fOpD3Je0j7eg1dXFAh
fq038aa7kzUYea7vZYcZ0b1RfBklDgx70qLLBZuYht5AYIlxJSBlG2OkfLi6DGGr
YLayfOpmujLFTIfabytrIF4mQ00mdLgHyVEACFvhKPUUKcDxyfQTGK1GJDkoHJqf
i3O/JP2iaS7O5UMSIdL53Az/ao232sGF85c/DnL/+5egi1Nsp+ltBBZuKhq2WmvD
54e+Z9x0XV4JWqN4YBwGrTAjaCvj3upTfpRHeqLvkgTrT0seVDQ2NwGPVqOz2wDd
kcVnn+XpP17TXea/zrJWt4lBlcqj/vzj+fg+gGcvsuAF/l3lQ8eFVF0IszodDd3d
BToGPh9Ng6MAC/uELYeoTE70aWI5ywNVnhFwPfslMQON2TWY/ClYUulOhW4qQ+0A
E2V/sG/SYaXANSEFig1qP4MoOmhvYB+Wd8IjOKyvUCmqAWeLj4VxICibiAlXyies
YKY+I5UHM0cMrUwQhD38GfjSMp055NWWXSz7nADXZE0nb3e2X341NOxLVzehwejY
wyHxouB6QrQ3GGWsJDPdYAud8RhAebn9x7ceWAfeUaZydKUHXJu4oD0IG0F6DKOQ
oslaPIwni+7SO18CKEsfQWeIySTFXxFRdk47HY/3xs0/HPdwlf8hPcpe42U4TRj1
6cfJBB2El2vcOZFJ+tshtJtniLOBg2UDK9B0+fTtadEKJpBgeoE4GAVShVRaQdPe
DdtkDXL0QK23HsdUiJbFXDnd3eiA3K4ubOYya5y+6tDLJT1xvh5JbVDyZoCQfZLT
7AZG7etdOMPd8eLpWvIeAlZ172JXggnlwvBYvZ0GKBZ1bo76GyJqMOQqmThVlQQT
W2LhkjyptgR7OKVR4ndoAjS0LHOXFlrQ8YWxW6aMS5md2qbWBGcumZBBEG/nZUZ5
IJhmcQHx8XFeAvn+2ztM1zNRf+CMDbD1kD+6NLhy/yWM4FDHEso+CLs6D1Yi8kRc
yGOWzRYX+0WBXYNyqyGqXw20HqT0/USoFIFmu07KUq+PoVwhqAeY774syYlA7yGO
pAC6ogj0L4jta1l+ZXiTQ5WoErhjgriT07dJEy2mcPt8c7oAPiHaXaClfLYiDTcg
XBu7khfsZItcDJSyqpfrNNh7D1INQ7qPgQcYxUS6vJtKoLdX89/si7tywBnL943Y
6IXcFwIESVJjBmB4D/JHgRxjD04Inm2OxY/6rDNUBDwjo0FRMiE1TTQxkTor4SpW
Ql5Bwb01G35HsLzNKEjQ2Z7D2vpMl6tCMa9t23qsRoebSL7uv+sjtablseBcY2FF
d6eotuHIaeIR/Cw4lr84kvq7UJ9ML/yusfNo9JVy5TwRV47869XXoqVGrtQGGwq2
72GNrQ7usZb9b5Il5dxPgEAIQzxDksva+9GZ+hi5zLy46fFHs3HFddbitclmr97S
IIwTEXgMfqnV5TF2oZb4dgD/IMLx9nr8mXNuqxwUaGlNJ3j9KCBh6MDgN6tBgWSW
NEzJka1GJrmeVSIB2NJ010fi5/HHoMuIkYPvpjYWYIRsWBJm2PAtLUinTIz7M6WK
A9uLblaNiWT5a3Z0owH6RF9e49C/HCOODIL3lEXdY5e2YgRegmEdFNzfN+PAWzvz
4/q89EFvmfVpXlHAkHlyp6NnRmXOttn9B06Ilg8nc+RhTx7cANBl/T77MzI7j1p/
4NGa+iP6znkQCMuAau5R01eK6v7rTXzSVF+YLDKCr7AKp+NNiceQmgV2cT0/7b5e
nevyGKPndayryJCE9AdfMiW9nfhu3DqROVLiIkaCkMygI2UrFCOXllPrXff50bbS
cj4sd2iBwTIiyKGS0OulFzUnybclPCPslyYWRXUCBnWm16u6TZfCij4GGMgrdb7c
ixgZf9VWHTich4U4SLGi8+t/MkLgd5Fgo9uzOvuYd7FCd9sqZDDIiFu7qu1fIuSN
XnyM2PjAyai5T1W+uU42tEs6AEs9WpDwfFiqS4Lg20p7QMlTlbJZoTBG42oIjdRH
9bARZqLVspOUlIraNvNKQd4Xmw7jrK/8yTJQObe+in69/+shfbeCiZKsLGT6uagU
L5Gp90LaZk5S/cGCusOUAi3aVcaq3T+kKEEwMS1rWYA021uhK00sY7GZ5P6KSMfC
sG/2fmBaJL+dPnNLaQ6RX4NPuuSyQ22ZpXRyp56k7KF9ViLxthZgXeORGL4h9GDp
+0i+XcGm7kdvgsmvNxQ8A+gjugc9Q3FlDq7xcta8ax0HlNKjmiGdM0Eq8SCDoQ2O
9fb6THmjq4Ptn24b5sifVlX2Wph+9XNfNjyJjTHzZHkrC3948GTBluin4eSu9u6s
xAG21E+EhF9kpTBl/R+YcrmeKAOX0+A2Hd/kxXNxtxaXSnSOHGLWX0BfGDcdi5Ei
lEHaHawHTK7tBw0cP1N85yR+QtyHau/DdtYdsOugoheIJgifKlu1jYKo9X4v9cTt
OzteEKRgxAZywkU6ljZ5UzCNct2fnwOBMl2k+AB/1hANfx/xt4O6FgiGHmxV1AH2
ss+ClbVKgvxd60HA76l35n4RNR2qbbbIKyd+hAmWcHsuFMoj/GcaoJrwMt74g7ka
66nK5IxaZasScFTBmbAshSll0XslKjBhk0XpWAzR2Fal9Ho5SuRGV8+T5YbFbyJX
oH/JD5KP3KhJ2UPElBhsEBvRJE+NnBeVRy0cyQGFLsBBXfW6b9StIoDQUdk4aP4g
OjwCgFRQ65mflrNIEWWn/JA+249rvdl70mtbKx74juiJwK5ugQPtDyud6rbuXcIm
R2CLKgjW+MpzOwBDCeHHe5V6bdBP2uk8wq9Y1K0nb3oWZG6Zg+eRvcSFw+NA/i+8
wqcGnN7NHgkzJM1WCnm6iJSlkXBd0qmaWpUETC3Q+bFbIz2pQMpYaFso4/KSc+AJ
0sbHdQhtV3fdFXkFVlpPjzsavT7tqIY0qhNAaRyUZLJbUG8mSrFVSfV3JIQrqHMP
WpWJcQ3tZWMpZfAnZOgcBaDFxs/U7YgXcQbbCeRR9NSCRE/TzuR/H8jgx4qbxShU
jVKJMayg4jqWxY4YWAQZOD5qQ36b6YbUNZ5FuOzjH7kBd9GhGiTsPZ1k65Cp24vI
G4/SazTDqleceIHbFkqNNpT6NYT6dedHm5SLoh9LgTJAZlIR4Vb6Gl7ZBRUiyo3x
CASTgpKM8+nNLij+MOH4Ky4PzZyu2BNVIkY6pE5q/mWLTM43c0w2gLKXdTc/UQDB
gyd729arrfBNlFWVt0Nae5MQq8bkmQpPA9otdHkgSFQLdaQ/E2aCkZssliYRMdDT
imKQoO1fwkQ70A3Lqm2joAGHWiYFqA9gHdQ97DiSJ+7X5vxdgUxH6lLDowMB08V2
j1fkPswFd7PLnXlRKuEzb/j1RiVQ97LNQG75S0mAYoWp9iaDV/+8UKcoAD9AnZ8Y
wGOajWOYKRtFGEEUAOuLuYWdrZ2HFbp8YYxDjSmIk9b0grOEtNAXYBguDiIY0VV1
Cp2GaMwG6rwnHaPwkaYKzGYyN7q0YKA0pvJVSt9Tc4qff1ca4/wmA7CwfenqvotA
PtwlblKDPrjfWZxch9BAPaS5ib19QB7NcrLTH59WDyALWbggy4g8ef47s+HDuLx0
nuylj6Z2RFnpaREPYmZBNq1thyv1TlkPVgNNWRCwgoa1e22t+otmUGGeuPBg71/q
X3lzNTZsIgOQn76D0YI3FV51ylCmotRaSTM2H+3unU5XA5LPFlxg1MG6Usa6ucI3
eyQOei+qUvuCLXYCsJ7undC/OHUI6e6bJ6tp+J7LeakscDggdZPTO5T0UXdFWCqD
RFRdYK/7rshNw7fT/xXBKP0DcXtIS46eJ0N+h8gmZd8j9cnAN8uKwwhTZMoCkzm/
7nRy/JDHZq0eglJYcnCeGjF8npfkwdVO1Ug95MgaWPcMMf82MXE+Vs9x7cX6B+zJ
s/tmDFeMQ1JBfRgU0iN0Dtp+oWGGAjNaNzaSLwtp9x20P0Jx5oxrfE4fe/6+eR8t
WUoaEQh8i8BbX0FTPCxmdJmGlXTf0ZY4eli1g2Ol0m0OFuUIQNKRshn1YUXJbXvi
EluJeIpWkfT3LKt4LCSUjYXDiJPuJ90QXNLDxoa6mGapmr6a4QL8gD+Llex/OrpM
jQTxgDAjrcXBG617sg6d4j+Uib7iti3ZkRbDGwZq1G9x1H6i8uQmH0Rc4JREOAu1
F60tVXcm/UmALZLMINcSJHqtApMiMqMm6vNAk6MnnCtxtvSvjBMUr/YjCor+u0eb
vqY/PlP78EDn2dJREflN9QKJr/bDjIPmZ3I42zdhJP5D5yr6ERpnAlCrSRKi1zW3
9ILYdGgxOvMLfr8cIibJn34OyIASiZ5W3ozMTbTSpWhF5FwqQrvkMvRlpk2AjKpV
yOga6Z2e+U+WX2Ihw5vdC/6/Q9UciYvEMj9iOvzk89CX/c9B7lphRjOsMJEm3hWe
FfZnJ+qeXiyNpW/IG9y//2B1mIPhSBMF1R0lLeMJlB9ysYAa7vWGDP7LfOUEnBkh
3y+r5o8ABq9fS1DnavPfF93W8JrXW7CkMBfhdSDcvVM5ckTyV9VYJX8vbt0AD4EH
MpUUQEXRSKNL+xm1hhUEG5kD7a0EOPZG7Hd/WoXAIAPT5gdMP7uNObavFdrMIVbT
gQSGqUxwVgnWX0IeeAVGHt3KvvPeMhOWDNouNX74Y8N29Nc8iiko/8ZPYb+S9yn/
BukE0VP8p6+YKjUbA1Q/TGySJYiurckBM6Yxq1ufQnh/szDcRhBwCVEq84NM9sCn
jJfwEEsanRrCjDp4PzE4c31VLXWFylj8wqWayeUgpPIomq9B/wP42VG9JPmiO4ni
hgZ73a3qQGuqFvbv2z9iu2TurKQLLQ9IW7ylQkvYCX9pDN1Em0a0SQSGZyzN9c2G
/QavXhmA566sTnFcjPaSH4q2I+C9lNX13OZAOlA2pen4KpCzCCb5swQIxUqeg5ge
6mmo2fMVnw3/xsFaHWUbK7CtToGTxB0Mc0U3JPfK+wTGWtxkeXb4gXSVXU8Hj/kQ
HcKV7Gq4xNXmdqkQKVNtTMybh4Dl+PFdsQoYxDFIzSZi8FzKqcktJrmFXKPvEeOh
zK/ce32ut4k9YcQTXeFpXb7pl/1Lyxytjf/OLS9CgL5VIepZhwlvnyzrfkL0uGAF
oXYZ/lSa6vkRs26B2PBpK1a2t0P2ep14EL8HZUTxuWMRF4xObt/pUKMAgHLtz+i+
x5u6VKxjaoIIGThL8NRYEzqbe4U1n6MmxxtQfx8EyXyrYmIVhDOOsiuQddgKkpTf
a2sPo/PL6jnJGxducAtB3phzASGB9bQorirAXSyoZFtRQGB+sfUKYGVh7QNSWA6x
c5M4oM4sbCy2ZylSYuM5M9e4enlc6P1IOib2WX1w/yxPBB006DGnOxv+JfiMxCQX
KdXUpKt2E+W1T1S6UrFc29l4xbZ88fkaVhy7qOwB4MZ/VnVODqLVPyTmHdQAwlMe
31cjvymKBMKbALe34EuCBFrEOCyXCHdvkA8b0rW5O4/BTTcN/oZnds48uYbQWa7h
+y7LcrBA4RHYyU0fDgFrBAKZGSLhaN8dGUx7tFXzMbA2WssEePAOO8JfbXA+Nn6T
U3S2hxFXqtbrS5HXkBuQo2UvvSzfekC0S71SAeCmwEB8ZcUR9u90mTL1XlYvN4gF
rTcwzDluH5U6NnoDtecOeB4WCtMob/JkXxLlX0OoX0OJ+DM1pJxAv5i4+GCVdmbR
j+avRWQk32seGJzfkCsgvjIa+MwqSiZ6sAXhLdEyUkIFf4jH5i6Q1MkCgc/O6nto
sfXBEYaxRJHjumudWNWqJM0cTPxDcVipnDiMUcmU0uEd7NBQdnBxxzgwMVvnNTds
cDtna/oykyWbAsZIYcPiHJWt3rcRErAh4dVaYFsJiRI5xygY0xldrrntN+CRH0ui
5LXTNFNHg8cZwRlOilfqzE2U9OdB2i296mtRpwQJLF+50MeZsEIlxMJn0Hkk+r4M
6LRGQcKw5WB0KAP3sFsJEIYy9nFzH/YZMhHcos+mmCK7rBn9WjLKEkClBsBN18yC
G+E9hr8sqLdDV0da9naxyq7oqBkQj4mrWAnccEP6an9r48SDr/T+80ky7ClerAST
9mxc5rvApxf8SD4dIf+dWLnfoCOJhZAQZ3kmNSl9yUm12dCD4bIKUimHg6nRvUZm
1COKdaGZTIChvF9GMbHr31+4hVe3H7gIBNOhC0q3PAS2rWCQUeyzDSUhVK48kqBE
k2rD+9x6AWEyGKDOuxsV4f4IyjyIJ6x2Tg4+X2WAfksyax8e5SrDY1ipmBHl3A9k
wRu1QBBLBvucriq1oHPDrKsMkROcPoT/2pkYArW4pyichCU/7d/QRE13DeNp3295
R7AX59SjNDJYFCoO4UyKJuhi73lzHQfaNJ415keqpTtIiKtQvTkTH2mqX0C6162q
o+3RrQkItwh9JwF1VwsljLS78iXO0oKweQYTkpCkatqKDRJxXcC5y3YthxCIYDL8
Q1PjW90PtddozTop2eF+kU3h4AlaDlQsBl+vZ9GTuOj6ytJG7AYId8VCgvAM+tOo
tY7Nly/HbzVQoGyoTMjG83S4K/zT8jcZ3Ju7SWRYBh4FeFVfoitDE1AXq25lVTwt
fEXnV6qbVeUE46xT8qbskM4JxLkvgmNhvpROdCcm+RmByoTKr8FdDKP5E1t9c8j1
LVb+t8gYkz28KQUb5kkwecyAxrfZNOrxzDovBYhwwa0HP5sgGKOGkTnwKcd3z203
Ed11hqTcrOitS/zKnfvmsR7VU5kNjpywzr1eAIHL/jYU3h2vJ9PugPeglqtSL00m
diRYv0NRfIyJdfeGHlSmH4FuyDA9sf54/zNoHLgFFKH7qrS0ixOz1x/iJJOFBR9x
zodVIS3P2A0AfCgE580k+5hEoZMSKeAEKAClhx+VYE7THjTjKRO29Of9D6mjcyvX
haclBYD30lDq5LmuBO5FnP0T8X403QTe0V78QSkOx6OAckAV219CUfYNrGDACW8P
4ISgmePS8mmH3QSWYKIUveknFdXam8WKJxKNfyeYMq1RgHDAUbOa5FAchSjvZSWR
uYUZqfNU6VAEcjYhyxu81sANno4uPVcUFtiPP9dL9UhgqkNm6hGWIROkIcDo9NG1
sUUp6I3mtda8Q0STb4ei8f+6hQLpvM26DN9FbDvXvEyjHPA4S35Hffv66nhMSMAD
l1hzGvK+wdbSpFGlV/E8FYAOk2O2uCKpqEn8aopP+9xhO5H32X3E/L8tyhMJJ0fl
g5iykXZtQWMD+RIqsppQeHTcmRuCqF2moEWWz5126Bv141BiYIjZW7KGTUyVYWe+
Oeuc5EAbUqmwDo3mkRlfmukgQwQRXWfOuMGmb7SDqL2tA+VyUEaRpFdA9sNQwr0M
i0hI3OJTxzmXL9QYKcP7xZKIv2IQNW25yB/svOJHGMsn7+2rhp+H2/jCx0BphuKr
AERez5y7ZwIdkvSWl2uGuxhPbabifmdUNr5goMV5oGdbIf3s87S6FYVBvuEC6Bck
IxGZ3851V4YLTCs3uFKgF8CpQDJxb4xwDPPLQialxI5Qrs9IHfbDN92fXYRk0upV
GRYipQaM15447wuDycd4nXFDyCC50dP0IQF1q5NTtfu/iY43kIjMrR1unRgw43D4
/ZfjHiVmn7bgg0Yv6OQN/G2Od4+GKVUlVOXNmjaS8fB8eY0BCdww0f0244LOcaBs
Y1t7X8ZCH2Hv78YZXk40lyz0D6O28yhmwPmAg1HA0cWFRM2zUGGXaCnATwPLdqyw
ReBvrvlFqJH9bJ5LaGWPnaRCpuWHQR7TIIyDc3Oj+CJhcFTLn6BN93WCw6nbACNj
OwxXuIRpsgxhkTeAo0nscIoMMxN/2lGgnIfGc8QrV4XasPFPq9F+AKxw6ulufaxK
T7N0oBW5gLj4695sQ4eVjxMrgNjrQnebdmMLh4xz9CzptT0cqbp3KEwnyxaqEyhh
A/m1q7j7UTTNd945d1zQdDFX0ioOAOSPxFl9XmheRaRELTHlr6IBXOFX+3NypCR1
PHKd1xJpPEi1E8pWTGlUSla6+lku+3K2R8AZ/oRSNq6UnJ0pUVVX9yL3cOEOjt2u
sKH6r7iImr6bEYZ+fqh5RWMQSzf8n2r+22X870SmfM2gPamQaviVNlcxq6GT++LW
0yB7TcLEPaBV1jb0a4951uoVatBEU3bcCwoaytW2qYqcM11qIk7PlymOjXlCaEnx
6zokx0NJ+VunDHowZ2Y64zkCdm+X5hjQxVky/QsOjceVuiRRo+/qht5CresZ+cPI
ee6/qhF9yZBSmvNnAEu26+RJ4GVqQttZhx+k79DiRX595pJwPvNmROUp6d2sK+1m
P2UduAecCuRaNb0cUM3sVAnXy9wQ7Qf7gHKr7p/pqX5HbZINamwXMTB2wnlJIklw
mYCeJs4JFcjgdPzF73W5+21fWhO+Tem+YWe99pkKBslUnrPqLjR4DZ73nTWUEq9M
p9DdcOKNPtWzkUUb1UQetNClfGC/0Ur6xQkzNqiuVL7dm2Oqxi0ioQaGzWiZ1p8y
T44MKhZdaAzWur95VcVH5o95qpWpwe8TirBqapugzHQjISBUt4Gk7fr4T5ByLs+d
i21FZJU61/SqRrlHPyVGmb9rTjAjhsQsLIWlrlvIcndqrJGn+7VwYxW6rh3bMbIK
cK3JGxei8TpLHjUv0ohDN+uaMeWm55o38QUjP0z8trBZD03VL0fnZprjHZkX1Q7H
f2JDuYszopH6aH4exHfF/hUAwBI9+sx6L2kZI60rkEWV8HkYYjs37pwonGo5AHzX
plZToPnBr8UMQdObmRSfl+ynw9iJXxLXfkkq7OBPGb7VsLBW8m5L22fg2KZdgJlx
IeTpEzQKrpbv6gxp9jJSL7a/sM801TJ6DR5fmMjVYL8hVdnE0arBXiZs+e/OeCnI
k+UDGSp/zW/ApMyuO3zBI2SLncdwiucqeoiAbwVGfW4q08sYX4N04g/ZeSkYNraz
uFkLRVW3L+ygBMJw455VqgK4EMO6EsrQ/mxSQRLsfiAEUAy20JjwtrdG33j7dnqq
bcOaugwsQDEiuNYZEwtI83j95rhGWU/YvV8oebAb49G4hU9OYWDDx09C+ywctZYS
NFTjw1xQu+9lHG+YMnxQwLRRso7RLR34hKS/fsTonoUhBeg/jdMhhSEdZAB9X9Cf
DdTa5ksET81kJhcGmGz/vWFTp9lLSkm+h2dDbMKypWzZUecpshYFXsVRAK/5qVUt
f347mipLE0yj9ZpP5gn2+1kAqUW/UZbxiJmqNSsH3wn0CYklndBudyuzl6ij9g+O
e/qy+GVJPR4PZLm0Fk7YG2Rah+u4XIo7/ZZ4JGYoUT6csmWcKjEB64vWRfD0WW+q
WC+FmmuAEiQEqtxBc7GfMAKZCUAQeg4U8ngGrVKhP6YQDRfXB3qF1GtkuiYFfpRV
OuQRdkPClffWbi5FUyzuKbnwXfXPqPqODAeCL4t9co6FWlobxtZcpJIXJ7qTs/wr
c24KzekdfEe0dCBg/LpMFfGiSWIIx4Ssuya7BT7auwr1NxdS9kI0Zia0wJUUXFID
r2vYY4N9XJzUXQMcs54aMWMZnBVRxPtnzifNeNuX8S4QB349daibW6/DBN+nv3Wv
+VNxokJkcqEp4I7uoLatYkxcSrP9YQ90vMfnHngpDst6Iwsy6NZMePfn4resbhuB
zYAQN6U2JmgVWlPxMWAZHhTLCH1q2i3JnE9UIKb8offewBELBD4wxJ06wl8Yoaf9
tCSTuShGFRNUBNjSG2Qypt4mNr3zHMHU18esYUurPXGQ4KOOvUl1ooaOFxDfGh9k
qjBWNSV1vX6n17cxzHnYOCR/2gpr6USAOcEbo6DnX4lx5BUcFNXKHR094UthOt0N
Yk0uirR1evql1NaTMqEpZ4KxxBqCHB+muZS2AYWQ+wDu9Q+AI9q7AB0lncGQ951Q
oKq+MtLy92FKcFRLvqaxKFbkHC8dWZ1TFXuL6egjk/yXN54b3rf/8KBr29PVlt3U
CmybpkKuL62ng0XbYkiwJlRuts/oprvt7oGn4ZyeCBHC92sMt2hH77ygpKuVEafS
ZkYjAX7qZupMwaOa8eFUJmPWjmPrh96fJMLbyD2NsQKsOgek9ccUFZOVfe7UxuyP
O1tsqb5HvmHnEz7/A7qg+jRcRvgCa7UzUyYlY0pY9yFp5/uA/X8y41Ga6BsH1dAC
onIfJg52f1zUULSRw0Qh0q4V/zK7nXCGGAgxnnxhaqCY7ge7paP4pEWu4cky7jIY
XaEClNQF5TWowNnWONfpx1ezIeLI7zBR/0HdhhFy7FevlQOhGSJoMJFx53nGGN6b
wmsTpPYfo8dzciV1vC4GeTw5Vzg0hGtWMEhZQzloj4DypH2PAn0qZlwNG+VtYdLM
cA2Z0CLY0oLlHJp+Snj5m5H5loxE2ZJCMtnJW+Z89Y9hmip5FJKQZDqjoCAEZBG2
O8gZfeZCLtxKpG431nb+cLleSzagmfng9qDONlH9q7w1c385kds4QdOYAK6bEaB9
NpJYXcsaiz8kMCKF1Vn2MAWPPUnI9EjhIGJqNAQodcUyQ6V9S5fN8sjYodIG1vCu
z9C8+hwqLEb6DRZj0VNC6CHgaupGsaSeBaJ3ijb8TZiEddnl3TqnqYMBz8/sJbLv
ZQQKN/Kxv+qWnMHLf86Uco5CT3/Htq7IJCIpaoVQiRpmozD9j4xABlCIk9Jwc25M
/MeITfGsh2CGboUfJ6o4fY4mHte19/keKdadfBjMqOFT/MpFdX1eEHsfF8QNB9tU
3pqH0PrSka2edxRYjdXbnbYPOjz9pQSKzauhCCySLe4mt9cOgLpzss0VXTw3s1AV
KvU5hnK+6OnEiixOUiamblQkCpZ5952htZYDor12G75Y9Jx75hMybamEZbB8cvt0
53O9paRc0gVkOU53pN5W9Vd5XKYRbI7vD9xOziOlzYb7HokKxe+/pzCg799WU54/
R3dqqn9RZDGMXMRmeKrkqOV+AdfwBgL2NgGRd7bnskcwqKbmUPYo6ExWHC9fBRkm
znVYdUCLO6h9gSIHd9qfjXHXe9Ro9YJQoX1Ak6X71U++45tka+NeJUNk7ZINN5tN
W6aAMBMcfFglEAyAW05vxeu97vZ7lKiOBqu2xN5wTU3sM5bc3Jy5/Qdtb5uaixTh
ihwVVEn+pf2a9iJp2V7zziikq8SILt/tNgTv2Yr+WlPN5Fg0w2K3EE20HXwBgHbu
7N16H+DyE8o3YQL1J4ps5T+K5xUwuojARN+kw6jAuYiZwAW0Qp8j6no+LT9menV2
3TbGSe5Hn+mM19SRMdFC8+H1p5c+T5EijclBJ6Buc+nlYh+sI27Rsq4mnyHFlTQm
E3QSV7ePpAEXYNmo6LAROnsUJWmLk5BnLyxa3vOEk9tcAa7vkyJaS4ZIldk8YuN9
euXeyymMbHULw9xNhbgpNjTpjEiSEWRDh/yLsCYcFowpnXCyjeZyOuhuczcFf5Qr
ovroR5HOjv8jP1tcqF6+nfOetP6i63IMfJ5KebYvbX8sl42imW2BdnFlyhrARt7t
V+2I4x2axa82AtPNruUoPE9l1wmZyWGuoSNK7LzPWz2dKXpORK2t3rO4yPV2+yKE
rJwO3iBDpcs/z5DUVSjycneyuCHv6rd2GdtizxxPlPzwK7lu9cMCmLi60n6hXrSd
M5B5DSfG5/QLW5Vrtvf3oleXfjnFtZGNGj2Z0BJUFqBVxAEhOM0jztt8/Cohgqqp
TVFCgLcFmQo5k8ngKzjhdI+PE+YDCcIRK8bsmR2rZ2yipCyfCfX6WXBS2vL4eHSa
WFS5yARh5NVN8uNrXaymtMycJYULHy9wLBWEFPcj8UXI8Vw8+FpG8adVsCJTiB3T
ZvmDIOLFnfKu9XqbyYEyCN/x23n9/34fSxJGm08a31RR4DDEuBBGVac4pZPgOUoR
GC2IlZb6ljPPDRsIzlnZdT6J2h1m6Mzuo3pzu3xpSO9Utgsw/6jorvCcsp+/8IoK
4tpCoCRKhOlf2Z1RzBgvk2mcqsKN/ai/ebroLj/dv3+vc++o6p85bZ5tF15lxdJ9
oDw8E5/rFm8Df1pvNUbGdaMzh87RaKvYjCCDsXa2O7WUxSELt/yLjq4Op8+xipWu
l6itCdpaiBMfKRa0ZFzk7LTCXEmt5tmZFDdK2hFBzBuDtdDTHlcjwZJNerO8UNPI
Da+cWO1rqiDc75buaFN09zrMjFe3lJIEqyzF7yQnAYebom6xUwxoVdpLlDPCfE50
aG2FvTFLWnmYotUIZ2M7Ccx3vSLPjqI/4PpnKV05h6U+1PkodJFYmhufisyOA9jH
/uN3zEzQXRhE6AqgM/er/wlcSEgaGvIrwelN6vokYHeAt7ldeqUtvNZefKzZpb1S
UFS69SQKRptGUuLMsR/+/RRTU4o7tUv7xgv72y9UEAHzBhkWKmQoDfeRYDatsvMs
FigP+qbaEWofKm0t21R+3dy3kM4JU1EUXqUEj776QVKC7x/yCnN58nVIRGv2ooLb
vlflSWoq1WWNvadMbn7b3v43PXWpawz2P7Qnvk7C2M5FBRqQx1uexbhnv7wfu1Cb
V5briuiYbHrZ1XatwECVGdwSwSwg7b1G361ge1lP1TCh6OlxuG2Nzj6KiXoMzQIw
i4wc21pNS+G3anIJTKbeyBDDAwwv43kW1p95qnAqWIvegJ8d3zV6yw5jXkExR5QX
neoKFskvhnr2VUGoahrHoBZmv8Qs4kvhZSE4JGe5C/1GUpBbhuPjFKJbIMl+4jYr
7kpIOCbsLnAmGq94TVXiXDRjK4WZN85OEwzg1vjTMzJKNdDRIPxZjOWKbP70S2ax
dPh8vAtn08a6fzDRMGNal61991z6CqqyRPRvcgkZE0vEoELktl29SyesmXqtypw0
C+2lkjSvifke3ome55frgp8I6gDB+RzWavJk9Pv194PTPigbIqLKUyZMvs6Ml21z
c8nPrnFb+x/ZeJno7MVpGpkAnK1cdCGu4eWgXWyRg2IJgSzZPD/TXbU7AJ+ScSHr
NazoKmaIolthynfP59gki6J8q4T/8RQT4Rw54R9FEhgBb5SrYnwUcirCcJRYhUEx
YYC9NCrXa9/4uWwR5i1jNQNrdw7QjTXQ+AbEExpb1eNL5+4XOiHGTtA/YBKQxF8p
Pslgh7ZqINZlOX1H1zU639JkWW4I5L71KT91fbFSQ12/A169Rc9gKP4vBi7c693+
dYsg8ux8aZUwUOxImsynY5S7LSGdMYpkS0lfGBCfmvfj/O/yekDX98xJWN3l+cv9
RUkf6q2/CO27otaUvz0JCDqi1i7zBeisGE7KZ4ndwqbVE1V6EBxV+FFUAWLqxJNU
X3GQ5UgTgCJD6KrNGFsS3E5TJSDvqhNd8107XXrLzYBooCq4p6BvDABmwYRM/g1A
Qiyue4rDAp2VcB5Gjv63ZGk7i3THvdI+As9HFSIDmboIvjG3tRFhZ3Z2OE+dyxkR
zxRMGkrQZn8O2ROkzGEDwwHM0J0n9bG24NFgAzprEsl3DpSKVHQqmKHN5OFF3aEh
vcFWQRH3Ub2EjsNM0Ecw9UMVirrPMkSChUF+clH/xLuQRVZqtCd+J/bZI7PGOrWH
fEfrFDgpSWRYj5It1aBGzwn5OmTWs6j66y0ctDH2bz53Al8a0AQmTAbQCjkq6jeh
LVkw7RfeHgKK/Qtn0LNmhb+XrDXcD5e3ftjZ6c0A4z6OKYioHMgGrYQggmnCAwub
iDkOmtQxePduh7iZzpWWw1zymb4HNjVjmnrvvfK77YrUUXCAYy79WQJKZq8YRBsw
9Su+Ux0LiZTtFywNm0gub9uXzKnf9Rr8N576c0ahRphKKdgTs8BKmzFzXNSTpBie
mBEP148mv2Arh5ZBJJuM7Dx4oFE4US9G3EWlC+4uSXSG/+BFHoUJgx1NDYHyM2L5
vQuYy41VznFTg4lhy2rT/qpHAY3nTf6PW3XUK246nuPY3+6TBt0lrta+1hudOJGy
KLxktkHGvNj96Tr0DNxz03iOOb8FFSY1wKremX2/SwvGnbXIQJEI6CuE0pijlPPE
Ria0FwRdc4ZjlGKRaC3qCA/cKNfSS4Z54umvWIui5IsOfbjo89bijuVU5D30Cd85
nRvNRPzfMyP+WkWXDskUHl91WOM9UYKVJyJ8FVxKGVM5eRnyg0bsQZy9eOUBHy1w
9Q2FdSZwddlfm5KeoIUSDYLSLK5SaKe7Mp/ElCglc0eKGjTZHjdHkzg3rMe6SgYq
8EMZn8qrWRsJWmWm9q0uHdoyVs/iCsi7gwIDYRuZ+6Y+ksHqv02Neoz4YJtNQbIA
64OZnM5+XW+XsqYOowWakZG2s32ShFdDSPuY1jXBM6+I20BkFVyfISQGkLAeaeJR
YFCLLQd0V0cYqXTScEopb2mKnn7/ybgxoQ+ofgiemGNsYjDJacPY8gD+zLhVPhW5
1qBuL/5Dem8okG1n+ECymyKXxfK6LhYGkvlmm6rnnh95ra23fAuZtW9n5cG6JebR
DXvxYHx7j84J2o69Q0xE+S/kpk++ZH9Xr9I4pv5IwEyaZNpjnUmRPCvc42gS/X+s
BIChg1M3SlTiqXM6cF4x0ZkKFPkClbT6JnkqX5J0PpDXEdwwKUPitSuUhQiiLhPf
wNp38/mwNSonu+l0/lFnS/dCsDUV+S6XkjGYceYZyGdkDsnK3AUCM9DPgySI1Ita
0Ki+Bfa+vr1gqY6cQOxTYnfp/wYrwLWZAOXIf+qvjCU2WN7XgYb8XndEwMq+BHDJ
EsQXyCgkvjEcsJWbZG3BW+RXJvjWg6clCgNUzrsf+pnaZ9bVRMF0fnoGHDY2A2av
SykH1iSdYzulzuE/ZutFJVJ+qipmhjn64DQtmRFLtNwkFaPsRaKRFy2vCcUg6/lj
4KvPHZQCPwdIHIE5P3GdrjIZAh/BbK6u7QrW4ImVDEhr+tQ0W1pBzdY9pAfYyWIW
o6iNrNsPIQS/777WYPE5q8/TcLW7WUOoCWf9U70X10bJXnj7PJO6h7lPtHix8vzA
TAtRFz5vlful17jug62p0vdQ2mYlhutnO/f0oBThM38QOcNIYRXDUg9lBNF7Jj6s
wqzV2lhr55102nNYIH8740bQnWALSCZA4ovG/qgjVeM6COqop2oh/QK81bfrw1Il
acyWSq1IO4U9Y+nEkJcXW3fFOaR5MSXKHjK7cPhMln1K7rF5EsDWRC63JWZwx25S
JTPo3tUbT5gm7YE/aVBscIs8NL348Ga0742eHX2pt/sWiK9tOm/FBY8euoyCj/cR
BCNyxmpa+eah5V3MqK/lSo05aA2oGiWOABaX4/X8fRgtT4H6SPd4I9mUDwSKm2e8
oQstGCE8tRyEpZzLEB9iwX2yqb/iEJu1BalDdj6wkPZmNz+rpAZbFljIjpN9TPZh
ac7Lx120UES4XYoVxEYk1yudQnVwLLUwqaLOE27Rb2hbDPzt30WKpymtJBvuzNJa
jqG6jOUtTssf3tZvpGqws+Aor/ISDV6L059WWuV9lZs0bhHOlkUzy9DDcKBfTINI
cmbeYmGqaI45Yybo4VrpZfPaHJ5Tuoyktk3qomYuqkE2yXj25Gawu326Jj6xIHS0
KYz7qHjrZt5Ta9ywFSr0rgw0d3IA2gNpShlCrNPzeSuDSKXnRBB0ayR3q5xw1XXv
1KqAzviW0QKy7AChFbn4XiF55o2NJ+2gOmWQNfkwauOo18IJtwfHGeXGOdOVha6h
jEsqxUs2/ONoLPaC3jP8nquWcvX9EskmG/IxNJKmXDmFXTSRfzzVRI9jLKP+0iFh
Pw0qjCNlHGZ39Qyg1TKWi84bk3Qp9zVX5zPqWxd7rjkvWNk+6Jve0QLP6c4kIIGS
6j/UcLtUnxl9RdnrugjYTxP2X+bw7NHgjLGPKsuZ/PDt1qBgfgq69cKsTuJsWBik
ZmrUFXOB2nYLjVQ/4fy6H/20jGPpGGfSiBCRSt23HhCogS0cJKu9HBhmlJ2zvDhN
A5K+Fn3ghvmn0nsxe7aFLapfdSLMeslUEQLpTRaRsbuo+WcL6aGy5PIZhiWQnOgI
ALxeGjoZfmOXkFKuBpOzqGp/xN+fjsw434x1MF7C0b+i+t3T08tkxoVamcGSvcNK
n0/Dmjsl3M0eBJsFUacEcT2HGlGKS7GMBoHILTGvyviFUUPXYBoJdUb4vi3NsADu
PVdDaK6UrRGO65KqQtL5BEOUatdn13jcTppQIFbnXBSWDuK0zh7ku5PGdKBbPYzu
cjFfDLHZ7pUL4J2cGKQGE0UQ2YB15t6SyHTLT4a8dwsstoVwh204olqoFP+02V6R
aowgPUvOgbLswgcJUjAdf0y+waTSualzTszIYj2pUdc4x7Cg+E1sBJ6eRf5f85z2
I0wewj9nYzvpbIxHJmVrK16EzerdHxFs69r3OC3nTmCKzY/2b8F7v4pDIB/ng0nF
8qG93rXozLjFWQyLXx8WfMYF9tUkAhsdHM4F3rLbLASXoTKnQ7HKuLowmjLSGlO5
YtRgmgLjQ9HQQALWICc5chXxOmhI3rcOSg9d2xy/mtMppNq9kVwib1v4v+neMSwY
hHSinxzwwxiZgWq0cyHdEG50X3nkAi3zM/w6f1ITWWkDgd0VtEa7QEQN/+O3fP/A
luHuM8pduquY0uP4xQwyNsQPMzYA+vjhBTz+q9V/KmWNZnGqzKWTmsKzjXjOeY18
p7gu/aGzVBh9/hBooSne9nK/3kXi8DQymAWQZ0zOTtkBQoHxMcQgl2wpfUsZsMmd
2NWhQhZVhWxc+Ov1aQ3YBLJKAH+ALWI2x1/3oXtMQRhgxuuuWwHOTaZGkAgAT3eR
SFHB7IGqxhO04C7GqhZcqgqVc0Yt6WHbygUcRiGhatOGjEC6rA40X5EgB1NP75hZ
81f+hupmMPvPJXGsJy/wM1ty6XbtCxMb+Gw43EfBIsTXNPsyBsNML58bujCgat/y
y3yCG5F+Fo+Q9k6ncZVJ+tdXWQxxBhWan4aPVwvLOpBV5hh9Z5gZ8xnkXjPGq6U3
qSILNjfNqoH1Km9Pse8p9z3evEQ1dF4HBSgNHQ1Unw2R1CA84JmywZJIXhGC5MWW
1ENVh2HoWpnBzg+AgJbOPYz6wvneW0xwpwNlaAFtskKqxqA2040Uoakx+9EJEUw0
T4ema4wxAi0f2z8SDWNVk82BkgXdLRUBlSjxtrG5bBopGFD4u3qGaqQMn0vujme1
/Y9/xt0qbV7wtMiSTfajC89+uGSdo6bFU+I3x58jaVZRe0LBpnGbtBe3Stx/q4CK
GC1RF4BIzF1WlxQ2n9Gv2k8jugUfrQpzwamGp1Hh8aXxMfKimrPPuuhQzXkOosBL
RI+8lp/XTKz7dc47HPNWRW32q7suwIrXW4hHaJP/t+YnEWwTDvYmjGl0AAJBERvX
5zaEeFbxCO/CQmIGHzo0krZ+fDbfd6JqZzmO5mX3oYwCmnutwxFqJ9FKFpH8eQHQ
BJPvZX5DMvy1Lnan9A2hGX9MzsfoAepFXTUpVR53sDkdSgCGtqgBtRRwqQcpCuSC
SNSxLo76qtPBmW94zzQy34KIiWPGcPT1EjmI1IdycqYPA6REJ2z/bhadTGr//XcP
hHGcKtxNe9/EOBCVHNNRp/0oGoWsOGcrbk62HYJ38t1aoO9FBXetUMdyTggcVht2
`pragma protect end_protected
