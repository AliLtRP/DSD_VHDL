// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
QoTdVAVH4WRSlvcdwIfRy0Ud+Zk2hmdmm2KInD0P9jKseaCkN4GLfZqzB4NGtnVIDtfVRGJlQEbX
r3GGzh5O0V47wwI5EBB05HMdRy1ECiOButuSXkCMAKKYpuebrHFVZIwiXB0Aab+uCcBeqEc8blDO
C0b9l7r4ovAzMYhN2b7zB4ehh2CM+8BCCdZ1js79puDOmvJnKy36AiHpn2eO2Bf6YS7UGVOFj9px
+7cwfoLrgGolLU0cJ5WThoZ54Ok8auptgAcf/aWe0efgvQW26go2/TOJkPluKR9z/z3aHwwtlmDG
bwreVPnpA72K43WE+3cx2waeePfK94X5qkVWjQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
YoeFP1LXpwKijzdXS/b8vYAzcX80elF5mEKAt3Z/tYm9NF/tlICOtA4NMapAOwZLnujmZShJi6j6
kBfA5bZx0OYlcA2Pr0sG2lQLu1YlQTM5WgGkpSISgSIaTgXauYIv9shmXM9KF7PEton22pHD9j8s
ooWRr5rSzlwGGEQ1+2ejrOFoS9P337J7nqLINaP/Rj8ULzFK7zBhF6+iE9MBRI8DKgQLwQnQ/Tk1
iqoJ8fcCcJornCzzaOp437yOBrGjwLX3xDdMQKLQO8OG8pcmUPqFQ5FBjziD14oA7v7l8G4+w43L
cRvIDmuJilWm2EaEdtBV2PO5eTQnKvam3fE5bA0PgPQBEuV/maRA8eze7C9YGKVNv+KVP9V130PO
/3X2dZ5n+vqhxJbrzawhXlmzW1OUt4vR2MIJ4wcVT5C7713jZzN3X1bCVQ4ugZLOgxwfgdSElRwZ
eNQ8WpqWjRswsHKN7sOBJHd8gIZ49uH1XEqhFBQp2bsmVgk/lZR1f077RQK7OvrK7Ai/NF7mv2eV
D0XCC0PTRpZCJ0DDwZOB5Q3o69QSR2ZujlyJHg+R4G9kNkaLef7GUbHeD4mQxRdo8jXtUuxWQxYF
zgWezkopehorEglOaijA5p8wFIDrlr+F2HxLPFQL0JAvsWW5HBCyt7NCoYj0WY3EE7PC4XKdyRs+
NkwssKpnFoTCiNhHwByg3SK4scwQf1KkVrG3+DZjp4b6CfLpbuokQh8rxVN3KxF3CCyfbNhV2koh
kdWGH73GuFbn45lt9ekMZ0Njx1BNRyL4M+uRpaiL5zvr491M9VhJ4O8bgLZBwmdDho3UDL+xStO9
W/su2ewVVjM4tsZFY0RMRZNTp5vOp73/+b9CRvxF1FN45YO6leUx/x7u3o8zGfXCDR1L+FkVIbZi
OFAgWzXJziPBQbtCuZ5ea4hmyVoXG8Ip02kD01SQhfTIXHSt4+bqJfhMu1n454XcxKjserhPlidL
Z9ghjTZ2uS34WKufR60vh39ibTPf3tnTUFTwIqvrGfee0S0qvYTpSzEeKcSlYuOqGrMUivvrbspI
r+RjkMmlxKJtWr2TfKiAQRUaYZ8HmK7w7JHI/yqNriN0kh1z54J95LO/bro9Pt3FPwjj5U+SWciZ
cHrqBx0k/lriA3RrAia/RgWOG0M/jGm/oBvJw5pnruSQkGV3rWo0nEt/a6XBko0/UW751yZMgTza
EqjtsQukAN8f8aK106DivWvSeYudvWMBlLFxpwQfhpW58PNU7mh59189EybbBDETYk29BhceI1z2
Ibx8ZW/f780uZzMCIVd5M5ia5GN3jxdulKrdE9h2V00ehe/lJFm3ksfkbKpWFmk7wxE3SWnfXjcx
DTfhVo+vX4z5V0XTOsrClMaqW9ZqO2/Fgy27ien8fvz/rRSEXTfiQ9U1C2efU2Vdu/l6q3Fu8kRy
Ua4xJiVI7CA2SADml1qMTS4Dkq5QuGwr5fKCXvEscFgM/PIgSjI7ouoSWNq4Jual5rRl8IVrZEDQ
BK8jLr9AJGHTTSrPxxwme6pcJ1NYHcVzzWeqBPzbU0tSVRdd79HUH6D+sK3qZ2w5FOMtwtdDIoj+
MJZsR6Df4te0sqkA3GyaTg4IYH3lDjZObKAQ2PYBtJEdiHRMOwcZhiMgfrIjSzUsKf+oDuidrYbv
tGLkBsqh9fnU0RfogJb+EQtffd9BgFYGZ7o4Nql9F+lp+rUkJ3WmwtvXVJcpFp+X4xynBN5bwyfK
Wv2uAvXFtyS0xsyRGIaAr5RkbFp0L3xKBTJfRjSTltXOZ91BLGTx9J4+7/F6lRpHjahX8Y9pHY32
NlQ8Kc+kK/ucmx7heKs6uAHhwZn3Ai8uvZZ9dCW3jhCcZmYaoU6oY4vkG4piYCI+RKNXk9iUVwJP
n/N+xz19T+OFRDReW2bufZ5HXX0c4xIx+OL2tBYHvzk5zumv2hUCXSp3Mb5hl1sFtLkJp/EvT6jt
9vV9oL4DH7RT71QsVDrguIMWXIxY2IC1Iwh4fF2TTlTQrL6OA/w0OvCmGpTigJmpQwflrbqYDXg0
0efNA6GsqJkItycSJNSQru0iSJD7DkuekAh0MNqwtptl1IWCqssAhld6fZtICGfp/LNfoK1QOuml
UF4mm8cjq7AIZ2x6ep/PHK9NIr8ONDHbs/3OUkFh761XP9RyFDkttZSziGD4ZMzjzM5z/s6X2o/m
+orCJasYgMd/tmwzcwA6iqTOueQvtUw7nkhkgySQZvRQMH175CrDjvv9uqb48kYBTKeXUM4U8TE4
4P9SPjiJe3C8mJFN9VlEnExmeZ6TqbkGs5c1un+AOL0szBEhVCQVjjZKv7yPBS/RkDHQkPdyJUbL
T8YgxuWrdgPUUkcq1DWBUzicBwJitoOn5McyOuUbW5zuKzC487UDXFhnNh+6TKFgHFTW9GZUId0h
pWcBWWbJL50bkRFlnODun3apBY80VXQmlkT+h5jvry1Ff62dUwfsXjoCHtN7GIHXm4vkw/kbsmFC
QCpbd0UI/WMAd2CeTs6iGEPbBbb6vUurGzGF2n80QhxrYXJqoSzqiZfHSUMHPqBdwgTs5zoNVzfD
9iUAZl4+yD6SEG8STX2XB3sJ1drFLaKrBibawl6/+bAQuQJisLKW9euGzki9hi6vy+4TLRiJ5ljc
HR7fOQaT1tL5hsId0NeMFAUU/tvbDu0EYyzBC+3H6GAtrX6pWUjVjsXluy6KEfLq0sVuU6ef9HLY
AbRFB+8PQTcFrMycDYQ+6j64RA1P3QfU0KiNp/GViSyBCaeXKYmclUmjF6CN+TQigwS43pGWeAOh
Qj2PCuwEc9mK0xzqynhgtfbXF1qGqnXEauf6/BwOTvSkl3DMbOT3EwJHPKuvLYIQhY7aK3JX7NDU
raUMgXaQPwvlxDNxBgEWdPWZYuSnszY9r0jXU3X4vBW56+icsqYC+PYMcelspJlQAcJN0Ck3V8Uk
dXJHbH71bxF90HAVcW7XJqqw6VjwsQCwXD1dIYKU76tcHjQnbFhXT+S6p5u6dzLMimGCbkNEB+Lb
h2xbM9E0LuK2dXSq9Wvs4C+3aoPtTMnASMKFwfB8Te3k31y1JehS5DYQadMKsHO+gIe/wtZ1epwR
Xt2DoNX8TRmRNeRuBnLplAwBspd2SjTt9c023k/SRY7EXW+CoMEyXTqg1Zbb+j8u2m6VaCiLsXZg
GfwPoLRrBzTDmRzU+dLrBq6bXdujUtMz7tV7k79OWCwlQlNPFxl4ioy5YqnWM7YeVcW7PUoDUh2+
6IcJ9637I+LPP1aMUaY/O5tKuM5MNSyfar3W/0k5QUvUwxgTmTfDM8MiYPu68Utl698Al3w2rdRy
+bEgynV0YPoHPfBsAvE0fGqKdkptRHXlqmLuu6suFuwf0LN2ZlnfQWY6dY5wzSZ+tkZLcLMq6V6M
Les6SrgFUQfoZ3WJRS6p9r6sWTwpLK/Imwi2hs/jiYFZY/83oCdW4lm2kv2CP6VbPNSGg7QmeklN
l47i745Oe3s9cR3VWxJ/9ITDKdVONA4obn3YYVpzc+rXH9QzizcupfjrKSnDsBtSBeXC+mBI00bB
rZNg1sEfuydkK7fylbBJiITJxPMh4qgyX9aObjyANWy+hgFxrGeV5VwtmN1saJ3isn9uWI0FbCpY
dy18RbFA7Ikx8kHHK4yDtCt+4+A3TSgTGFFcAROtZXwmgwyywFXGfEz/vK/ww99+hXhW2gVY9kTu
TIFu2uVLrOBYyak2ZTEBfj/PlOeYZ+jWYy2CfZSx8JWIeJR/ZbxjoBFButqKCwhOB2IrLDtpmz6Y
GiPoE9cSk4Iv/xbHtABNZCwkoQKdBWS8l9BHS9x8G117iZG2RzxQfFUwzn4tvara4RAA1UBxZsWw
DdMynjRMHZdYEmVUrT5m3PKprAlntHk5m8qnltbD3iZ6zbvZKvsAhxDQDZByJmlzDIxrOVO74W1U
tdyBW+LUfrgW+3lvpFcN4EtUViXbd9PdzCF4fWY1MDQNY3TbTQ016BuNfHFICIX3j3weMn3mKcKQ
7PwWR94MBa1ZNM+QI7+zJSvz4UDIgBLGveRZ/d6Sr2jN/hnKGnRnPTwJtcXvlB6pHAdwq5QDYPZ1
llurijoVlUERkItILrDv6qDIP8pnLvo7t6zld1uGC8R466inmL81sABeXqynx79QV+Jd0nv/AoEi
zB/ftLpZLBveEllRC2IAHhbIqDaG+AC7+ERFJ9saMwm7UijrH5/07qxRePSlYpH5Wxrz6lsRyp97
GhoW1jqMLYuNGTPtBUCLUC2FLBLhrY/kZjBZ4i7wgPLY1BznjTl+9GiaNI7wsti6/KQM7mE+Sh0Q
IRfQi5LJG2B+yz+k5bIyC14GaPM+tgWwhap0hcDl38MndFKYiIf17ojI0CqV6Tiam56R5Vme0eWM
jZM5zgYEr2t06J2yxlbYpYmHMh3mm/NksRw5XCGWCjMASuwholzINI1IJlWgiVJMejJrdXo6Agz2
SnwVdWz9VTe2bj+tPCP+ZKMqGd1hI6H64HYuSJzMe279mXYJZk0VZjzD10qHeTOVQlSDTTPMHEAW
/lgyfn5JwpLEEN6/accJmC4I/1w/AKCOYgc1jEnT6lH+h7Oi1oywJnAyc1ZPd704PmjGha53ZHuj
lGyp2SEVF2af3Gp/MtvGehgH/Dmo0T/IjSUOfL9gRedtCVgvjhee0+byv+ndPBG/XE8iUI42CBTj
lyYxPMmVnfZv8Jbo3/13SeOOIO0+ZF3zbfm54Pv3FCGFSsIbjEIDKTqCTlgU+doMlVDEKtnvc3Ww
Km5x2rDtB2Wxqvb7sJp+4gtvBLssaVIAWxelCUa4siL57iZ0aiINHP5N8jcxXKSt5OOBlaqRBwa4
lD4CRIOnSA+cDJugP706UgZdZfohN0SB8dw1hQSFJEYj+Fcqi2qAk2cMaFU/FA7WYGK8EQneJm04
QGCt2JNl2vlT6ZHFs/k/wMDvgGhcA0Qz4gZrBQnVFTJbYhDiYGP21gDBvDfoYes4OLjMVRZtMWEL
d8z3Z4UHKevrD9bqjxOe4+P6W7NODVbudRb4ZmE6wcFP9zDEbJ4c73+LjrBlYrfLKVvfNFFNEjKF
lUZ4TMyIrC1NloFLbGPToqni4KT6pJyX+7vMO4TWPzYIwk3NC9IbvZtyxcPioA4cvQeOe9E5UB3O
cdALCZkJZGqtAYnVaZwftrjaypQqfLsXbXOQ0Z1gEMmFGCmuljWATK0bSjxK6xer+w+hXyh/c5Ek
1AZ2T0OY8bNatNhX44qFyc2iVFIB/ngqKESfhUt6/VDL/bAY3myg8Zu67l2of/8fKrEoOVr09h7w
tsZY5t7utUNxOA+9eOYQ5apKlalvjVy421Gngy1HAPig1NmvwDju8YesLcLp5O+l7VaGkXHcxhpf
ozHv0RZL8JvKvlD9Nnks6ETxuNYXWBC7lxybYLxTiwqhl8tR7hIDixC8xch4QOiwJunrNG1bktdk
d8OA/XAX8cVJyvkvjOgkya6QI2pYi9X3yf79goxBFDH5ON9h8Cp9oXQSiE2J6834XFMK50Qi4KBx
VlCSIzh1LRy+Ue/ZcKjwXipi7XJ0HL3CIcHx5Plmeopj6RNQAtA+4TIumlG32ngxt/nvgxoBwGPk
kPXweVn1uyDIUfaPNhgA9JblK6qPOBhQmESPlA1YT9KRBO6iS+a2PqUTPVxBIzkpxtZ0XGNU7TR9
Ui2tpRmY7PR0bhewEhTdrskEAkZo1PMI/5NOQCOLorlMIG7Jpv8gob9tuPtI9xTuGdEln7c3gLKk
ohZKuvXUh4LzosDTKFP25Y5rfKu2c6GSxp9FbApYpPKh3Y1A79poXs8GH2K1hlwTuq3NHVVCCA5t
AH+InM2lH0tjtTIPZcW+t+FBLlVL7A6adl8oGDEznSrGfPPxUagF5xfUh6ZtFNFpotoNAUNBj54V
/KpGUHvdDqFGlc4Q1SqX7vsQ40ent0R4PZkmry0Vt1vIyvbNwS7HHHNRD5zrOZHEmLONhTGJy0u/
snkY9TG+uA40NwTwlrXBDL+xwbjYDgG5NWBC6YWAkBNi+T3uiTvz2nM2gh+k+VCYkFFbcC9rFNTe
LmEkoi+ypeC92b3YGm870HI+CSD2tok1y8buTiJ4ozL3aoOaEoV2WbfHBHKNf11I2fJIAEJaV5oF
eLgn9+2VdUb6Sf7RXgdabpdeoIZwaXeIYBodeZ3pz0disEKz0kusC/vm7vxNiaQbzzVmXsTtWAXC
7nmb8pGBgGEhY8bqm5q+fYnNHRTYju8ocMP3JcAs0xA5qNjcKXk8MRF8eO18jJTPNnjeg2+nknmF
2N8Wfo37qlsM0VWN5Co12q57IOlxYTSkOTBM8aFai842QVc7vhnr0ttPL+dVoA2g9b2CO/kewJJQ
Q/95ptVYn2v5fj6PqGfM9Fujee1Lt72WLx72k5AqE8Xi1CQOnzjCHeH9KMMTKS2y6Wf7+p/gZ0wc
Owv9K40z7mgpp15U/Q3kvHuljZWXH8MyaBUfzvUZbVwz3Lku3nM/EfVR8VscobUXIilPTETgJhjX
BeXzJ9SgNjdal3n86eY1/UnEoLtqPoQtyYIOGQ1tCxo+k+y3mNT0dBC9rTmznUipdtf0lyq/6d5Q
Yv2El9QtfN0FnkPYrDYCJk9Wl0aEVz3MDZKJqjt7KHeBmxxNhtd3M316TAcOqEEFIwKUAjAlGGYe
0jFzI8qNTd2x9Fa038FrFCVUFHlN1jS9gwQ7zRMPbky6//Qje6VgF9k2ns1q9AEm6/XtZuMM2wUX
aEcSvsHfY6102Oj6WXoqTQvCrVJfBAEa4keXdJ8mpBa5+0tEI7910OtrSoXAHEMz0FhoCxziWPVE
uLyaDGC2EM8RCOaNM++WOEqynqpFcxnZPu5CxHh5RAYlqVdcc5bbcxNEPkNNTmR0mzQTldVXPamj
dBbFNS/HwrBGWcetxNoD/vffo46AoswxkGawdijEOtR7it6ukvKc+KPfbrUk61F2C1UPc/LCkFGI
KyQv84v9bEZm+iwPczP7zSSbTk09AUzVh05OsiZZtHS58VwFIqQKbypxNO1wD6/txCzddIF4yMcz
gfofDxHuSQdrKdRv/orP3MPTMgXlLQc90hoezevcu30WVdz2AMq4hOySNlrhSn94tsFby1fro1ZH
Qxn6dK1LjIagEPwJPWB82cyXIljoE6EBIJF5oovBvKafkn60iJuMPAd/o47ON4h+rAso4oFPSUXZ
PMTpqJ7aP5RflrcwCwL28NGlYrcleibthZr3pXxneEJJF7BjNNmXGj0msfncaouaKGpuuDsyv3Fe
9ac31ReoxsQV6z9tzQkVNqZLabTTvHG5EeFUhx0Z/Ug46Ii1uQ4zmocFjvfYBkkGGuywtqkEZ/KT
KxG9Xlp9PAdlMnvUALY+mT/7cK18f2Za+1KJkJkzW4rGiP7bTffaRDqHjKsHRn5cbzaJau7xU87E
rh0P3YkN4oYJG50nIo3FRSCsJLfsCC5yCd4iALxcSrWJGHi2hzK+9MZJZ/gQB4PYSk+Cv1OVky/X
/y2Vyfxke+U2k2jv1BaSK9Y2JCHIA7CeEieAsHK0ERe/IfR4gAvFmifdRLzHzX4jaZmSb8jWonmm
zYKehSG53sYF4egvww/9Et8fkKG6cWd/yMWx/gxnxatS+gcI46eenzBiwTkhp1/ttE7m+ydZ4q0V
7hLGsF6XdUmgg11jEiA48URQ1nMjPnYqDv90IAlk7Rm14KkT2yMpiZb2ioKApGmSf5rY6Nu+9Kn4
VjAic5JbLPPkOBGiyqyMxRiWTrzbBxA4svXcUdWpYIHrecnjstYG0f8VETVp7jlQuh6srebTeWdP
yUXLMCMWTVUi645saXANN3zLl21BJwg4dIVCm2riTs1WN5BR4GfoZVUq3C1AUs7RlwM3whgn6sMT
7NeJeHB7B+Uy+IZ1baz+wTyU3pFfZYVbv0Rx7AlIwtbKSMR8K6zM7JrE7NzEMaaSOtMICocPBJdP
JLLeKZEBnf1hHiGwV2w+UZv78GpbmAfvIl2aVIR0qqGH80vPpHeWswio7r/daPYDhaQJ5kwxGh6/
AThmyCPRPtd6bzIkdcGIOjGUe45UexuKH62HSaXzYMGy2UYZcEyAS2MtGL6tNftzzw4oOUp8PxYW
afi2XodAWT6SJKWQET0yDefprDBhTHPdD+RmmnNDCqTqVKmQL3ye3nhQ5HZik98KonO5A4C+7RQY
LHRd9F8JyUfVHOLHXVede6mMFvZqO6kZam5brHHRkkx8EebRe2o7Ae6rpvjPn6WE7lC5g6iO67hC
r2Qf6aYPiyHxVX3bjW6Fco5UGroPDeUWTJum2aMnfPyhZzGX2/Br5wkzMAhpwfbq3/txO3HfvKCY
x7bhw0Ao18WQib/IPx59UtwKz1zo7LpDOLm8qyk3+YCIPlaPkANt7xfN2FQGNAxgpsMc2fwFTa6O
hqrxxLgN9X94CeoFKWwTMulkmEj7thjIKBOqk0BO5YfLfBYlellFOZO4jyR5HIFjJOJaw/Cg0XMS
KL5Tan00p2Oe7LQxSkZusG421CDE/hzTuHXTIWoAqaCytt7uIl0FHaxoJqJCm3vlJ1J2zewU6Liz
nsZhnDSDgeNunzWWXJevtaLv4ZO8OKJL6/VfXGgychGr0UEAQWKQ7xZm1SYFcCxQYgiV92fA5kPZ
oJuIUYoBf/hdn+WNNZh9p7ufUsqO2tnpzQK8uZBqNOobagud9quCvs2Vo1/tBYf1zvK135/HTEhr
fuXinRTADOU8+A5h36JhgOLOwUhO6h4BXW8RNNcW7DRJO8zvQAF2ZmppO7lAL+4oZR0xuyFz6mi3
Fo3GlRDCz5rO92JbwrhrvQnoY6tsIcggTwc7zS1S/RZxBU1KEoSUFhsy7/XVrJZNIG/17H80Zs7q
9YEOQKRiYgtp6DIIB8PZsDhVwTf9rnqjScj01wF/0lbQKb3mKloPjUOyz+uQpSxg+sPVGIfnhNFh
uyOKpSxa1F1EbzH/c8rCJCUjZUGVkijbAvTDGhhVwF2VmRaZBN030zQe4Z+UF1cGkSVe8QFSCCtd
KEgaLghXHKG5v8ZIfEjSA3AhfBZTbznz5nIyItyHHzxSPfu1936EMM6LxowjkVErV2Nlh7L91Ikd
Cwe5ZkGk/jx62jC2NBrBIR77sf6WmPExMlJJLZbtwUdsyPPnQyD6jr12i8HmQ8sYgDO7170u43v1
ioL5PVwwz40IJ3UaCobJRoFPJTyTRoRgW1GZDkvSTYoPoFamEDppMEKhVLsPcqiTUGr/Ok/4eXlF
uMX7roeQv/jGtiuJsSn5Ouo4UAYz7f7k/q6pu0EY35dWTMwb8r/jLgAkepmt8KmrKuIe1QOD8hxy
b9sEzTSFeCQO6xZ4onExMQeAqJuI2xCWrlHKMCwIWwS2vI4LA0O6HregIgpAzMPSn8HiLRb1ApCY
k+aXmQ4kpCKoKtDLRUobETCxO4ad+7O5d/2wh+gB3G1mKtkAF9gp8Na10hXkqhS4obGIQPZubGN3
b9ZUe9J8Rp8Umf5g6yMtkx36R9sTHkp3lt+qMluRm8pBGva5nse2aFs0f41+NQgFdnuNfzXzkNUh
KAbWBD74gIereZlPCkj4ShvpQfKmYgn//i7gh2aAbnydXn7m/c4dBqbPB1iVTrKFySkd5yG2BvXm
h02Oxke4NYDgosrU5Ew5B2Sm2ds5SR42Q+mk8LXf79X7s76VF8ZjRZ8YUv2prut0VGeczXJ8ZoZ7
4ZaCHkuHOzR0EZIIrU/f/uGH+CHie3ElqsOy66sZS3kKgz+AyF32XYCsWhVNCUKNKNVdSHwe/cj9
Qz85qquEHE8lqUMlvaDVihP0QD7oTESKq8omb8AoCXGrhf9L5mWUscWLI0Q+cGwpqP9K3e7DYwzf
EFSSFKbVfcVMn4xamVgRe0sqv6jp3MxL1aRXJa2k8K2bqCXabxV3ZI23KGPAoJPiumP4MYDmwjnL
GNTYHnD/Knkf8SDGiiYZkAqxoJBytzgPQQlG8Wz9atlHZFjzgTqRMPeJesi9YFUy/89djcZae04J
f2TTUbnCRcPy7FR4GUTL24hbhNZsOFA8sIwZlj8x46xE/B+sarXXCxauAD/dTNDi3TVYgSNSWiQJ
HJYQSopI+1Df8IpgVxLNOmTH3Ee0lEud8nsHG3WgR6i6aoscWFtfxrOgoZbqqr2BjMw+o35Wiwun
3vHJmZxMqdvRRbIxUbaOy+Z0PHPtv7Gj7X5QKLeBVncOUBair9Gey/F+N5eS0jurOH2swXkkXEsv
AmlCQtrZ7ID0IUkpVLbSxeTbn9CkDrtH8e4puAduZTRJjRF1Ds3F78YqeGb5vuWxAP84QXsp5L1c
wafeSbT+netoKASuRls4g/Pdx5ZLdAkA7LsYMlLZh62KG9p0gGoOf+7fKKGA1cl0Dfh5h3VMScxZ
7uP2EZwQWqLVk16tyxpGcSWaLB6MTIn+ZOnVQTRhfUyHCs5HqT67XPTXqcaeRYpcTA5XB0Kp/o+Z
ssoda0c1L6QHdLarCX/ihKeIJpsGKC3dyqoJ1WIjh7JclAMGc3n5SVUguEp6VT/i4ok1mM0vqCYi
2YNdcD8C6QQAmJrQqxsCkK+noS6e75OQD/vp2ceR7zFPOsRqTN86s57f6KgTVxaSSxCpr+E6dD8g
lsC8H/8ImiOrTnSV2SZHIDFPlfNluoi//COlUrqpTW7bv0muXzLo/nN4U8LNN9XbiRd/9Ak+VkgK
fYWrsm9LZA9W0hUUH4d8dzz6tFPzup7QZZKRJwQYjTEXT80dBRSVFWnKgr1DAaboSWMiWbQGEqv2
37ujEziqxAqcebrgiz1Wq9kzrhBKjm/1i75AmVtxaKSPAb84nTXUm8J5e87WXynzR1WgLIUNYILm
D8NDp1l3WacyKOFA/9dvsLBeB3Y1WJ/wVZmBQV8H1VvvDJlqEHd+uEYGaGfmfSn9pXRF5IV7Z6ip
5sTAdBuOjyNzyCAOzmSF9bY2k5WNkGN7Dc8o7w6va/cN8oe4Uy954EDv2Hx1E4zCJE50Z0sRuuzF
JrMqUs2UbtgGQgkC2Qmc0ss1qSM2ffQVIEZDFc+U2menLRCXKE7zhN+duA/Tru9B7HfJAABIkV8M
e9ouUK4is9ivYOiLptSr1i34dtWzq/EuJjMZH9eKtZVFkyTOHN0iyFtY0GLUOcyPxnb7/bcWPJ9P
T2+ZooxjU7H5ENo+tHnHq0APv9VwNdk2e7AO2n0LPPUl/U07hAaCzEiRKLnFthIUuxC/mTnPJK2a
qjfr66mkh3MtytATHHgyxIrLDwO/oKLbKW4La0mr9fLLo/hyFX0SSo3ow/xkndtZAHbB9FlMnqRc
vsPvTTJOCNGvAMOJvlKuIpQkW1YGs5hytqZRzTz/FYoQbCkoClbKdy0HkadnoSqY5BKw2sgl3xVt
S4m2FbPUo8ARRYv7AoWmmGoM0ddgzbL0y2KQvN0ArVrzQ57IdVQw3rAlMRZg+USOtBT1zN+U96d3
FT7z4xkxOOsgC0S61xxpvJDlFVFo4oqvGnaQAEkTzf0nfvws67sMyNjAI80DD4JqsC0Lp3Y087Eb
gnfslymEZTpNen859o/yZ+WAXewBfzvKBkhbOHq8gchFYvQQhfzQHMV6w6fx/m3iYgkZFYWaKWVg
3FV3IqjFa8uKnLo72byGZmF5ffjdNrBOvCVXy5jN3dvchx2SsPI9UqpNDkxGqdf6W0lluH7ta4Ok
sGfqWaEVqfmQjHkVTczpsg/1tgzLOPG71Tk5Hc9tWVIqH7dCctCeJkN9DYZgnx8E50NnsV8Jw8F6
pBuHsRZ5tTsq65qGW+r+DGReLAv6j+T88HDkRY6SdU0QFxevMQHCdCX81aG7EqFJo9YaefC6eair
VL4ZLHZNw1o89U7ymbvHJGElSelyVgp0gVU1yIiKDKoQFtblvfGSqOKsWWNtIVmuXAltIwip/qQh
L7FnWyxUOYhQn5CpykZ0cyNDLYnh8QmpS8GHDStQ1GVIWAdKHZU+FBJNedoQZ8r4gdzZzxBha5pN
fi5ukdk2FU21VfaLFMkY2gEsXcZnU3Jj+THvXvFuVrFv5c6X7MMongU+7dekwpv4f//6zWiE9+5V
sKXxUzui38HGKWTemWc9d5p1Pu4vViJevUc1wARrnWMG4ZleqpbvM9p6u6N4lcpd/TSOGbW8/cw9
ts6krgfvo2rIMGW+9aANdSdcB1jnu8//ZVPLQX69NlURY4xBWD1efnBWaH9XPcYq948JuF+8WXnM
RvHMLH1bPddv6xvUmk9aTeLvjRFc1Dn3FaCrZ8Qk/W+nt807cbWrwKHbWFnESKc0JGOVpTJIrqBt
p/9vdLHAbAUdWnu6qZVEuT+2YwF2+fqRU4FIIM3snYoBacIwOZbi3d4rcOpv/E0xquEBFYsBOlck
x0aY2fxTetuCtGNarjKm3bwwm/q690HCYClQLRPY/8S1dXxzghcY8sOZOQNi9RQtRI6nbN6GJrVW
pcVpJ0LWRszOI0luy95oBbiJ4ypg1lY5hTXy4pkc1BYoxSEMaBCRjTPmjIpRdMlubU4aBgqUKrTF
RUTOr3x/nXevAxhzYSxtW/vQ4BQfZsBglSDL1DMp5uYrj3O8OFThr85GNWiXSZRMnR9Qmiw3wgv4
LzRvigoWWOhaLthTHlFIWSDMORk/4lc7x3jKlXgH+j1UUVs54xxUbPpGIkZl1AUNJ9hRkmjGSZ45
5Etv6LRuhEvB52Det8ZvuVLC1b8E6Y5DV79vCfBDj/iiQXej7zA/1G0Zt0H6wKgt+MXQSHAAWek6
vpHy+XSx7+uQTKFdFNXqlX2PH6fhU0enAZpYHlqKCJDPtvjZzxuOHjP88DshbwXnAl5kMOdFHpyE
cLf1T1PQtfR9NmEo4OfMsWXex+VoT+PPRL1ZeFPLtBj9MbfVX6KOYEoI6M8Ho0JpjovyAXI5D+0S
2G3t5IGGKgBxxLRRXBzWVJQVZfQuLdqUyE1qfxH8mO17GU8mjAQVc1MVjZZfbHwpjnWfaAbdruq1
Z6CzRzZkKZwe8TByzX0u1sOot4148d6Sz/xvx9X7u/PUhwDX2Vh3cqwMg1xl+VIv1uVXzf4Qwf4w
PGL/r7/+J2Wn4L3Y7v6gqWaKNyr2symn/pxhnpYnhIg5t/rcZlRqS1wTmcL7bO3EF2AV7pkIQzIK
GYjsND6A8aG4OwAilJq3VQnmysI/Vn9I2j+ecxFudQgnnvmVfx5zvXdROBJzppGZRDd5k/+TKzp8
Rh9gl83mQcCRe1E9w9K2DDYtcCmTN093P/YjmTFB2/3EGniuXc5o1hqthLwxMH0nylmGFhDY9TwQ
m0daRpnlN0xUvzZFFCj3DUjQQcPiQIo64kujOBU2nOkRp3cLPKOytqZzUx7zdIS+wpubIlnL0xnU
9MbMl/mglrInR8RqvlQCOJKYmSc9Bjv3T6qxZ1MLazZ6F0yCN5CbYvr5n60OclLdnNyPN/umEkJH
obHiQOqspwrBZphJQhyaInS+8+PyhVr7adOeRNlmZ8j/fZ2EByAHTVVMTDvs/HxoU8l2HkiUuNON
RkISB1LsQRxeanNoVkXfjEYePAEcskDtu3PcrUxfcmM5Z6j7sDKnPbXa0YL7r/r75VnEwr+4Qa62
KRwbNsl8O+8Av/izaw+rS9volybc4DDL+f/127YipQduJGX0DzbG3FqFv3f9N+JHPMr61L6myllV
rpFz1vOMkhwC5ZLxWI/j5yV51g+IzwSnzytBSL/0HOgfQG0mYH/bwc9hiNkPym0LGknr2j2uETMx
++WgdQX/vRh/95qnBIGPzJMqRwUzRWMfsyvf17zE2ljoLHxl/F/TVEpb81q2DwOg3oLePCDTxZO0
88oAjAT5wwHIs7x1neL18WisYmJ96PxTT9iIY6uZT0g9czeKKmzoA6brfuZI0CKwhYqJ2QcUEJS8
QuWVSmxnAHzj9JzwB+0pLVIFBtSEwa1nPjKkLjfIz3II8Yi8vFZ2qmk4G7fMtd+4Nr1u+QfHMG9U
koj8S5VCywJCb+XsVUbgiNqHStHcd3ABwdQke7x/Km8UcgLI5SJztMCfX1L+Zu/EbzK6nLZE4PRn
Ae3SKSJ8DfuQBwzKLBy9DQ51AZeTMDyOJd9BxmCwUtVMi0rPixG29SOrYinIdhpS+/4lGeyziXiz
Ks6Z05UYO39nKIdKX9MO4XU5tiSBPEPkAZifxQDw/+1Ca3/RHOASegcUvVoYlpu4q35eInAThPas
MJ6VBFAMOdHG5tSWFkW4MtC5i/SOMR6/FgbnbnHIzEbL+tLaAHuLAWiCT2bk+EU26aw/WHH8ykTi
j/BQ5EO3UPSR9+SKKvoHXuV3A/TMO0WTi5NdVVcYhyory7XRr7KARoij17chtUmHqu8lydloibj7
EkTA9rTVtEMHPm8xdO5Ssd+X7sKb//1NvgSfPnrtzPR7m/0oBFfRAnrcTsg5LtLlDbwDGtTY5YEc
2VkpHf5QhWarXWMqEMW4hjN7mb1pbnG2D/Hc+LRSDHc5+PxBZ9yJR6WcgpR0nQ5x1lJ69kF0nWq9
WMIYyEWtPCJUyCOoO9lhDiLZM6SS8L5NMjkaqheAZeeOvpl07PPeI7j8H8lMn54WZBlBT6l1juMw
VDIpSuI0GYShztBYmg2e8toqSm3wWRPP1NuFaSdaOOQOkBJAuDpxn5HwMZGRHlxkg9Zi9XBVuM7Q
6WTvOj/eG/U++vO0JA5Z42GnG9mVcsvbcjbu8B6EUp6CnyfdMfwqhKriJxVHMVLo4lg52ns584CQ
YMaEChcbPWB1vDPs9CnfnvlKenYCfsvYKPdRY8Yj0y5hW6o/NLlqR/+sRjqu7oqX9m+8Ww2hp5sM
yzctREfO7peCqWuNtF1X4V4fsZAnxbm72Dr6XApbzF3rCQv7gnz3o94xYi9KJrKgu+dK206YNojA
5YfayGVu7OLZyoVKGB1YvmSwDrmq/2Q/5lZWFjDLWL4RHtkhx/bONUjwWkKHn0z7Qearr++8I+pU
I26X+PXzybGMqvhsxSt3jMXqfLlfxCW/aNloQybyKDKJEzSw7rz3Xw/TMtjocORAJH3eQpbd1wBr
vk0LY6vAS5NvVD8/2MJf1E95QNxf4ckFb9KKRy6/4HaabA7/sSFJP3/WLfiRdhAU3FFYuf0YdG/k
iCJo0fqx47cr0DDLPqQEUFhMvXehay/Xj1ZY6vvvHOkyzo+7TzWqEGL5z2x1sj82nX988SXQxrWd
jzd4R0VgDeS2S/RrQiHetRsCZD4YjE6Iw/rOD1ZLeCe92mDd6SDifNN/P+smAA6zbhtlnGGvkSmA
tQ6MfhNMBljS7xE06Z6rRET+1sB0feDWBQacU9ciyb1mYLvy+m2LQURj9K36QA8Rr017eAqzXe/c
OvmIIyvsvkwiMQtE9HlicHrq//q+f8uuQNE2MSZ8Vpj0ylC575JIf+oUy5sttLe4bP8aRgWqPJCh
M0CaEqPLDF3RDFWy485e3uEup/iyQe4ZwmDqjWctMkJgQbWnFmW2UDsjz9WtGbOLd7njloN0oeyR
F49AF74GjYYfgcvErdbkWc6JFP0n7WfyhYjOzUTGyMR8keV1N/ncb+ltZk6Zx/9bV5eJ00P6vyp/
9UUj4++9S9UOprnhgqrcyH8IYUBDBd8ol1nmzrO77WzWuvWKr0ptg3E5kxnRAh8jDfWDNiBH61PL
DITwqDKyuZ+ntOM4/MIPf/msfnQzC4/B+jKGmrPMEo13e/nn9dCIBc0ire+oxJhxXdJRcycLZM/3
EPOwh+uSashTqDpUIeBL3sBmDlCJTj6d83519DSwlacYF7rGXdp4MVWxB56Wd416TZT80FbuKda9
J13Uk9SRd57wOIILIFmp3KX4qaHw5I2c7zVnmpnyDXSnNXr4kyAM8tfW22TeUSv105sfi4lOvuEn
P2fnItZi6jA2kyexxCYYj7GIeTazhJCG2SVl4g35DzFovOkuBzhqU9iGazmlIC+PH4WFvGFHt25a
DwrsyjbwRBudZEN1Hq+RNk32SBCzyBchAFaN6tnI/0qB7wQ70HKKxk7sDGOXvzsqhQi5+cX+kSve
W20YGzyVSG8vyc260t5Zoy39JlgkdnZTYPzJi26JsbykRrZ5VkNxleYuWt1c1bdIUgVbUZoWUG3O
aA/iiDt13/4tAdVoZlxbDuWwHa5HEF9hz02wUK1q+JNI0crNaic+JECljCzxuVhbaa5XxGgFj0yP
0PQmgyDR27dE8x7LRyd5XpjASUZZdRbcAqJYct/KmLykWtng5L2h5G4/6DwdIB+pvhzevAjTHElg
HiYCio50e2JECwHdNHyuyT42Lji4JQ4fVAj7YUi5XyLkhwdLp2EqZ1tfYFkAhlYMZ/qHlnfjsYMl
cJN9juH3KTpeBnKhq4ZwJ8BxmW/e9n7CKn3gUjAatlBwD+rjcKQ2nkoMhrff+khP20WtOhkO5hCT
O9aN3ovpTiGqK3xGsqdWhFr0PMU/x35QzvxniHwXKCizqyT88sULCjpUpqBGH+raf9GGEq3d03HM
6zurzlx2eAMFbaZBaS7nXPwatbNSgrwyJ80319rYLiYD73qsrSdiaoGR/azqugNoJbDfMrOwJ7+9
bu5E1awK3QXZlLNGijFeV7YClZ1Roq/OMgGw0AfioIIQgliwjX31X5el+nvDefMCfjXFGWrbNkie
J+anOSjScBjWbgrzWCIEtaLTX56snXicv6cKzbG89tm+MLUteAmoQ8CfVjUZ0RrJ5H54dY/EYMFV
ikx7w8n80JjUaSBEV07dGkHNGUZO1QAG45eN3/1kvAoFB95ubPyqJgeqrVqjKUkacbyLsiIh22ku
Zes1k8UTM17UyAWewYqF0aSdZyvq8+UXhp3kkGR9WvUipF/flAaZwLnRmrqmK3Mbg6MSM+G+sX3g
7dK0MwTg5CoThsYJuO7IhkNQXgntl7WI5CN+u6B3s5+MGTKWo9RQNiBsrZJK79t0TLrYE/oxVCyW
V3l4MFXNnNUXyHSoxxhZaQqqYMG4/Rx0x8CsQxR65t8Ej8+nTcOgJ7iU0q2ASqH0xaALyZj3Ysdv
s5mzjMF+T4qYYSost+6+9xtjxROXa/WGzezQUyH5t0vzchYFDiY/Lx54R1rWBfIS+yR2KEn1xOWb
3MWdqAzSEdRXYiXZea/YZHqyMna1qaLZr4yxZsRPm9D2XEiXk76usjju13fXo1fovRlnAFBx5aLo
U6cXV7eaWP5hBJFegl9oa+I/oEPik2kzlebi8YDZLQBNSfToS0Vyc2rUX6ldBhbSXxHXpTWBvoSE
9PvLzXBy0zMdGjOBDKzY64vA7ALIoN+jqLYpIM/Dn5UyPtAfzceI8vNlPjaSoN/KfCZkpKB618Po
lQDrz14U9tME99bgJEmuLvt4fFZWD/n8ZwKqlQyziSDjCz3JfLEzSrIXdxrRGfDZKW8LCUOT6Ma+
a/WKhK9AvOHJ4n8tdQn0X5OgI+pW48BGaXnIIMsw+ZdMz9FmT5CYn76iKJ0aeEgNQjFKvaHi7RQF
+MQIGBhg3YTzMDQUBkrLDZup1e46nZmz2p24alwhXih6Ax8Ycu8Nw/w2/lpCZUuMHwW/kyJXNM4I
xJuS4njsgRd6zM2z1LxF9FCDSzGqtyR9CRzEibPxd9naIRJcwLVXBLHZAJF3uhKaie+9fupYYjPd
cyGUxI+7Lx33laTVoH7z42m3hK6r0g0ZNUMGSh8ohllnoDCzLPL6wpkptNHDerJCKQWBopLDhef3
PfPjudVfY9jjTLezGyoliLcZhGbr1+J6tqoq+5vZ9VUMveUyZV4YuqDlzJ2Q3kk/ABXEXGrmYg14
2rvGLg64HT8812g+/AptAGned0LOtPGKe8qaezLa2nuUwCjsDdM6TRUMHlInNZ3zU2qOh6EsiOyu
2WqDlau93Vj8sPrDqLVWrqO2kYQUO1quQNj3zFXTw/fr2TYki2Btg72ILAhI4dKh0joRsjNVxOuz
ZX8V95gKVO8YHNd5uvo4x1b1ksiKoJLbNqZUwAGlD02PQUhQsTnuYIXFwVVjkoIrZd8FBOYTNaHX
7VyfEAN+7hMnVOhfyrwHdOukrtrkntVKPwDiZOVviLO/1cq36JttEtFgvjlrdPDOw6DFblk6KAHU
l3Zgo71tUzwyAlFyCr0SFVYmmJbw/gx2aQUflCeHeftu9IXITppk69v9t1v410ShmbRbnmfLG4kx
jaiPQGONgPXYrKr/xD6cNgZePqVCZlmUvbyiq1HDkBUze/H/uneI6LeH1UX4COCW3vvTw15foYom
`pragma protect end_protected
