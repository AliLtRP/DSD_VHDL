// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:02 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Oe4AvdWvbhxKufGlBVaNRqqnKcV40Gdc0EfprEQiaHciAvIQ+Kn0momm8P2erzks
pfPSO75vz853PYUHyVTZU1RD6jNZJow4OCTf4tXgZ6XcmA5Bs/VrDdATqcdnXwh/
mX7NgYeBAgFUO/tk4YK5+euor/RZCj1ZhEODDn7+ku8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5712)
+u/2BNWVc0rDZ0fbqYJR+3ocmt1acOjee0fTZ2d94gFPH70miBDT+1PsLNHWI6DY
MnY3r0I/wRmuqH2gnX87qDr9HXlX3h9x7FPp66d459lFxujJ1XcVGXWieftrW6Yv
ZrjT7htBeL7qB8VKkYSZ31ehF4R9UNkOQV3g5xFDQs0r1t6U4GbzE17HK+Gp6fSz
ACUNt69NpRrv2/mUmNbqRlOLfY322PnHviDn8hpRPIK7nFY6t+Z2tptK7/njm8LO
qn4r6cHKs8fvbfOEaTUQHkD37qptB6NOTHeW7trVJ+YBqy8MjwVpTUNJztjXWLD8
ORZaZ3Q+NxTxLHvYJq5Xp+7RRQIvdokK+suOUug1ynF8H0k+ZenDp6T8Ip0Vjl4C
HiTO/5eZxKXDl969cudzaizSaQRi97QEs8Xs0FT9uvx4wDAue2XTfnY/OV6kTgjn
H98vCKoW7f241+yQA7o9ag346qRinyX0MeozaVy0dTvq+sKwRwEECbVHy5RBfK/Q
8RKERAHCdqYw6RYvv2a9MeBv6NOeogilDSKy6Ha4GfnsX8dCDRTnV0XO0qrWSdZb
g1SbYJFO6OLJdoYZlJmr3IvNSpyNay/WZAdE5GtK7zSO0IDfmTTJF/8ts7bj6Uel
WQ5UWxWTqi/DTRxlTrbcAWU/BSEeVjesostnyTe2xohdIhelPtSBAPEuTeJ6wZx0
POaFX7cGin0iNFJbAF6hdpoIcxRGV9roWj64DwPE+k74c5b4z2k7m8/4sckRwXeO
cY6m28p+iIB181TSE/q3eLw44LLHlfUi3tUXnBTYbS6eCEneEYIMHOgTDSPUvyMm
PiqbL4dvdZ6a+dPN6fWfr88hZIP0qaFsgaeAUjQz/y6+8RrwtWRw+DVLxldGu73u
EgmExvKj6S6/zptphUBQp6sfYyXOUmYxKmzjc6M9NxPvzbsuenJFoMscpfNgry6N
kdxHm7Dc1Nn+eS5mssho0ILxkMVIiiPR+gkE/msy7RcTbjRCBNqj2q+nCwESDGho
3bq1S0njHxLyRYcnCrefKt/B0V25RumgsVHXUIFwJ9wi9duefwDAvv6AKaEcTq6s
ghsIin1hpuz4Z8Qm3W3PQnfgNQcKKuyKGAWpya0Lcectbyx5AGg8zoVM2gK4UwAA
VpOd/AxungnwWF8Sx6eqbzBvRm2Mri3SWf9b18FoqOtdPY6JokFIJzBlcp47FLzl
5PwcE293oDvDHVLK3Lw1BJJNcYYHNtC51iqhi6alifFLiErcku1Y+4ji3thnOnt/
dMXvQmyrm4Cvh/r6uUoU+ihsAeNAluABgBhCiXxovDrS7xlQ1qCZFdgo8txC2I8A
Di/S4+2FiaPLUs54U9sf7Y2lgTzTJc7DspTTaelmfDOBcn6+Z3XHcEXznlujITFC
5U2nzqcNhZfeygBCoCoeVKmMWwtH0rOxzajdVxrOL497PPHm8cznN2RglL1EHV7V
rcEVol1/dUBbQQK2gPcP6V/ZUmEgYD66j33/km29qTl+wvbUxt6VlFAStCWj9S8m
My14rbGuzLxAnHkBv8PtCikzIEzR08ZtKkHeP8OxUuwE99A4eIgDbpXyPO28qLn3
EpcnTHGx32FwqWZtNRjyz+So1EtKaKU0fbO32I3y5b+YGX3poLoFaRvycyu3SnKo
Xw+s9gxSlFBiFAC7QOq8rfl0Pa6ZyIl4PoR/EPB9PBRPfB0F5zBhiwF4Ob2zB43R
PEX3+hm0bw3HW6sJm9bvQupXwxmmcA6lfcecMjeWVBpDDtTZ2xwAZw1Mr9o+hCP+
6tgp7oovL9OSlDtlSOcaHT5WcDbNYgfBYs4zr48RMkyvi7n+USYdVRFeNSljsrgB
l/3QXJpuoULm+6yqlIv/UlDsLdXDuFc93b+nOVsz8J7j57gUwxfDFMs4W3f77YEV
XeQL1Ou6Kr4/sCHIF0csJVm4bma19VNN5YWs/LY92WdreiZwao7t0EOuhhRa03Lx
imUxv4vEz7jlFw/7czYexR7VRIGxbvZgMECmXg2htwKiwv8Uma7FW5FND4Jnguf8
svFpsHn3PoK/bAIXkHyhWMXMvCqt+o5+oWOOEcwLuGwlMoJceaYUm5k4zB7zoLCR
yyaPMBc81c+bjFDZtNy/NAR45/s3mNX+93aijVYaIQwtWK4j3Q2mBwMI0dLEIW+I
GGm5MBVd9lX7Iyznq/Zo1KyzOwdrcukJuig8DyZW6Sb/sPyVjTPafnuFGZxfRO3h
mtIj0K+pJvmplMtsNL+1rjEXYa1/kixflMwsye2MxLse20QpwMWVbNYwno2FlCE+
8VHvkjphA5le2DhNoZEncUEw17Y1rqZ9005E2tADmDkFR38nze1qNECNx75oBeHC
l3QS5A9EArjMJR5TBAhMSbUM4Q65YZEr6j6LHCOyfQE+8fnirIfY9z7BJcfPcj5f
DpjFspwDxpAwEF1S5+EbjkIZ6QrYUGMZ1FCdSjFgFeH/IBa5uQYgOu88DvI+Qazt
16tkn+TK+T/ZBmBY80Ux3RPss5RDxseu+OIkrByPfx8q/oIFPHGd937xJA4I+h6n
vMbUe7cTVwmRmkurLibUO+a6O9Ue+xqoZiebeEFL33nkehSPjbX3nm3hHfQn7p7j
S4ush0ifqlBNHB7j9vSz5aRq4JVf0pK9AAv85HINv3runYfJExkyWLyms3jYhgTM
9YncbYgH8v6nhzm96Nygoh0p2lQOCXtuRrkU5QqkWRHzz4tbN+4owHHCew8ab7d3
UJeUhO0Ns2hmgqnJgnEjzPkw2QO8meLN569gha0tLamHak2QsYTi6OdHMhG4Tbqi
PVA4H5xw05AqE3IHtfPKmU5xytHMujLRbBeh/mAhhGZ3qqpYlOkCoXbDCpwjCTNU
tJ/BwIt+QCM2u9yh+8XTUs1n1MQtR/nXY4DVswCbFS4xOCJNO7uVcA3XvswdYqcY
uXTw5lmqFogt7YTQ7w/XYuXQLK1ageTDwSbiz/vWF5n13+RckcnGKls9sGOQb2w8
1wc7jPlB8AeLDIDi0y4P+3i9GVYEPZP4Q3KDVAycr4y/hkcHGNJ6o0gCU/rXe1to
hnrn5JjhMOchBf+WZ8IME5KfGLqECEtdE8e/JGPrHkbWJAUeTKyC7hit+TIm8jYK
URZ6S9t0nAHGnharH2tgZMWAgWBjo148wWM/ronnXHtY+nxAQkjsWkmwM5Jyu5ZH
/VjypZdbsEWxB9SgJ4mZErNi9Iolm7B9pJGUlMRkSRXN0tg5laNgv/S5xrgQ+yOh
tFgUMmzbZEu3qES5ljuesUaFqRFEkXdux19yPNUo/Uh+Vdf/Darm5b1fpPm+NhXI
9vgWAJj8LJVXAjTGTAUNQ4nTL8O/9LJhhP7oE7iuY0ET3WxpqD4aFuN7MvBW1IY6
Prmj3AdZYBun+lch3VyhgOiqWlWp+FeOJtyJ4gXcGXivqivfnapuu2KPEnwRt94d
DfZhvnIXtft59eLJVMHz/HAi633R0izWcKNujABhYSjWPi00XAdow1cTKSmCjOn8
q5iswiBwmggrJagLIhV3IL1+4YOElWELTxeMDUz+kk3mWLoC5ag+C2xAdN3a4srj
qX3l8n7Vtmtx3Bmcs4KlB10lUjvIc9UwR38bc5KOMLwPNAX6VYfuK5P3amrPOdpe
V1mI1ggNZlk7A4hF9g9Mld/YrBPUgM3ODMK5sxY62ZZW7J5OCP7IYHgxTpcsojjE
2EmeeJsGoUQGEnss4wgRlwzPRU7NXq7fUl0uM79Za2jEvp5CwxyC0xr4TiqQodcN
+K0FplvfQQCc/ds2VZ/gksLUs6WfEBdG9U6eVI3GF72uUHUrR+vGeqnqM5FskQiu
hTnEsRcgkkO3kgQxSZpsxj/pXie2B8nWlppXjKm8ySyhYm7fDgGwAVyR2iCc2Nh1
31KBtdFt16VY1GozO69SMwv2skAXoYe0CSwDpn1AVhT6Dk/xQxKMtN5IwPGPQKzq
K01lRMRrqj8k+0KpKnZiOEjZr90PY2bChbJzOQRwG7X7Oh1ZUlJO/Qcb8+GSY+vt
eR9BFUeP39dAcNl5BmRQACRxM9Ynlkc88N3Ihnw5wnQueIrZ325ST8rpXZXSo+GM
1C6FZ/WiaYRa2j2Hvc2ct6Bs+v2g8f05Kvb3Qr9ROa60SwwaPeSJo0JX9A1MRXOU
LIFqRNKIuYCMV2GJWrFT4VPx1jJ40yR4qmI6pxAssA61FrpjpjYpOOpxl5nUPwfr
awVHRzyHaAukfoobAdLzwf5hiDfo71GloGikBmsI9xtmJRiQMSA58i0+pRmHEdBL
MVXraBzViVqsLWe0ETrPaLf1Dq0AZ5TEQuG+UWhejSCevedMZqMrgp0ntLiiF3Na
/NM9hG1fz/vfckxoLHlMPQVN3x4I5mbur/PG3ZvrkJJptiPBcYjWoLgPFjhnUyJX
AcQi+oPxsI1PAVKgSO8F/549Ilc0/0DXc8CfbixppiITYTlddUi8rBcaTD7ePCKx
VO+NYPPt5sk0uJsRBbHFCVouqKnaPdoHxZT5HyO6JKABmP0Z1fMPyWqF6VMGtD9P
JY3TEghR3bjTu7KPKCUDzUHzqwrV/IVZ+ruDTrWejY9JiTb3wgDJcKAJs97bI/P9
IWxkQlND4Ii+IQJXJ7ZD0JYWfh3MS4DQE/TIbuGs5Rqf6V57hRJr0PYAIzX/tnln
x1y47c4WRR/sPDkWeWWWDaWE9/uoDCV8abN1rFqSViIUHqnoXA6GtDWztNqHCgzV
C7j9xWYLXhzuCVWJ+ZsGBKUZMU9MUv4d3kJ/+mQkxGyv+q96ij9vniGp/kj9U0WK
uMyn1d5JqFWNmE/DWr4c1nyE8eiG3f9zfGRPBPpaLQnwJGfBT/TI29fKKkuX+NrZ
eW5TyTb7rk8RsTAiDdwYvMBLcgva6l4SZAXUZBPVFvpnS8G1cxqPz1vO2CHdbbBK
oz7rYnGTFAPHd0tCeIHHAtDK8sWCVguKhBJ4j4ZaOBvM4Q/GjYH+M4CACGZz5r6K
R3qhlPWv+JKXpaTRX9TaM8gEVx0Ql6bG0NS5XKf4KpcZ2PeeyiDnExkq0N0JMo7l
b2IvWbmt9eufm+ezN8zFESVJ9pt5PYgV+71blmaWY/BasWk+dPZ3Oa6hum6bcmw3
NQVFxlbSgFKPSjNFrpSvDpn2a5zznITEt45+kdgPC9ntOodKJD+U5TXGbjKtYJex
dZx1Tkb9tsf5jdTDhqwgcaUeNUm3V9SHWye3C3cNUOf0Dm3LZvYHNDK3dYBeNvZR
ebPpkNlVBuhM7mOUeewFofNP72A2kmN5jSv7aT/QqZdKfQU53RarRfXT1aFVKwsG
T9Jzub2Cw6jDBWNFGpfHesdjHHwXh12qTPMUSJUfFNEiIL9HhY3Rp+aOPig31XFP
+JC0bsxBDggDWtJMald/EZ1mxfy/wLumeKs/2ciZMORT2PeDkv2M+87vrRQJmh7W
c10ZGvXZ4hoT0rOhp81awKm8EDwLdibgD29tV22uEiGlVQMrOvrp1bSUARPges4w
LphBXGlwS1BKS8/8NRPfz0rLQHXzuhRIhjRG6MoGD3CBYqlyix7BCuW3wjI4vtrn
y5iJ+Vlg1rei+nU6rT40WuJw/PhYJbaXEmUZ8mOVRhumQqdGMOnNNF0RpuWC7rLO
H0Kid2e1TKM31/gGErqch5BQhglsATOP8P6rQvq0nKf0ukT8VX46R3DBqqtik6tK
dP2/BLv+KcJa7xuApchXKN0iyI8sXA5knviQNTUaQ67SJZlinEQQgXvf1HmSgUwv
FzqrpR1lRtaT95g1XzX+mdfjWoti/yk0RB4ZrOzLUIDJzsoi0Qhv/ovETCL/kpHl
9qqQDwMmxHkutDiaayCV+166+SXahYr5OFCADl0yMtpICgZN0qv5ImYQrqAOhruR
2gIokSoh7WbnzwhTxrUIYvjPlYCPF8Ts/S0E+h4aZksFW4/x7KCBleB5EWOecRjv
ISupVXcJdIUIC8gBYICESFb2jeqwUEALv8Pnbm+ZrDqHqMP+GYLdkXe47/zcanY8
5iFW6T9AA5jQG1nIT7po5sMT7N4z+ijspHfU0rn5XErTnZQLycplOWFFPBMBEcrF
yxSx4GfkSZpclvFFijZ7LtRANN2SgeZ9IodC8Jux8u9jz1lIICZUeAZq3saPQXA2
dzLlPcc7iYKolAIFhuwjj1zbbutZwBbfwhFimDfgH8upMUTrLrOwGPNRCRZ31MbL
2+IhUVCEY5T3u3ILfPsDKbCMYzKVJNkCaTF+Utg1CrSt5A/9kmBbD0ngh6Ce7byI
whKqpvyoMuX4Ef6/TcA/yFdaqG+rRnxTalzh4PstvzwiDrbfFLeIo5jnWUP18cxU
q3c0gsp53dLLz60Y0XkHAp6SqxWBCOIaoGISSAbEjF7Oanhyh8UEN58EuvPTjUKI
OdhxDb87Gi+LnrcY1sXlqflCQ7z+BixuqiothSfqa597ISTpWEnNLR7toOFvXq3g
1mshnGyd7Ys4NIqtnoXF6EEua1PAVHPMvTGw4b1GgIP1eRBHcrxW517re3POfSwD
G2WXJaSarPW0WVRni0IH/tslTTY59qrcldf+YSUhGWUFw5xotLJuDN0++1sQ+Api
SKh7SMdfoXDSumSv7B/qybSnI7IREU1YPza6mrdZD95SZMYSu83lMoaaJtaAUFhw
aFAM1gqiv2emG9+joCYxcvi+TTJPvPIadRu1SPsaes8fJOep7QgM+l2Rd9Hg7s3Q
gi6EtpVQ7VsZm+cbkXsZL5X5moYLGjBGAIbpZ7vd24JALwPdjnAT1gooi8bPoB1t
wvmPFMZRM5XgUea56nlvFgvnDzb3NqadTYrtzqykGWsuK/PBgvEynKEBXdiLz1ju
qaNJqAWH7ARwON3TwJ73w1AGrScgb0QFnoSeDavL6yPo6TaY7qiYq8pUAq9Xmt7q
9edGj7MpHASSP/9AxhFdPC2FM139UrZufP8qDhFy18jkju6mB7LHBZ9NPCR+ZI4/
l+NhWDUta1pmZZtXa54kCo+CFl/EfJtZugon/XY/KcKAGjxArLyUhE6hV8gcOhUE
T87njFyD0pPFZEqQCWmZxGq3Y1rWr+lIx95HF6V5gnlOfPMzRKg3yMJr3cK1lHC+
B8pXnic81qu1O9Tcsy6YRIcRZjdibK+iR2/djZDOcSokiAl/Q7w4It82PHR2t2yf
oDL4lRcPzvjQEj+3r/PW+9/M0d+mMsAnTTYwRdnGnVo+lBnoUF5KwoLHRllLOM7H
TvRkzMKHgCu5vPyv4+h6iiRfO3ctHaSEsk3ZrvoLmq4cNScJcf4JLs61hs8smdAs
LCTGCpgPsO/JwSYoXZqYWBPqjg12Jo1c4NwJUVU9r5thRcP/kFB8lPLSx5vTZWan
178y0/eu1bKdoAo6jOuBdXldh0dsR0TGDw31mZ586n12yTfbeKAo2llCA0xCiFtx
SCywtNyEFN4HILp63tuF5zXz5cQxnytRm0TXrYafFFMLXyHFDgLbwU/MaJc3bSQE
LI1lHQ9EtIqaq22+42lcSmiB2Gzsbr2KzgErzRNub4cB/ExDm0n3i9ddMA6zWWM1
VCCCH3uX1whAjQiMeIxyDrFcKwXzFOobBvi5tGSP+GAJjE/kP5W5Y0MFASPuXfc6
`pragma protect end_protected
