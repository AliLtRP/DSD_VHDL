// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:13 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lzArVuS80cvrLusFSVHBAbFXqn2EnM8UVp9zLUy2rFJc9p6BtEeijSDU3iYPxSff
OhD9xaHA3jxk3dd9nNp89CVOQEF5J2/zbp5kIyGeWzlb6coOTWnq3T1qt+RACq55
GYkOUKrWe7UOC5LSyb7ivJBJuZZz/2wzedIkR/5XqpQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15808)
lNCMnW7wwJXaSRu4KO0kcXhMpjgw/nBBtwSSXjYea3sld8UxPPRJX2C24ahkpTpe
B1fZ9iFwcy1g9mwjYcWIPxaOCXZr5kSCrLZomH3C9Y7vRSX9M2VRb/dggPmErJeV
7CCaTTcuQ1UMajiShazXRLaESIln2kut7Q6cf1VNlNfbx7yvZrXh1ps6TShEH8LL
H+T/B3nBj32mVU65omLNBOL+3PidyasOcXCfxDUV/+YcNqryUTVZotI1onwFhJD2
b5VRzPTeItijUWtrxfMF/zxKoRkmbnzO2FK/ysHnw0D1FCnWF4Id4PNHS2cMpKfG
0G2ERIPpUhTATfee+PjGUKZ22/qHMmppCyU14EvJK7JX8YhHPqZ6ay0/U1/lAP7z
FlZQXDxwqOZK0TRTR+5rtzh4JOl4ucHeppPosHbvchfKR4poAm9TE1H3muopsPtP
rOUOCm0nIUJo3hTwPONOciJkRYwC5EcLQN7HwIiKHA0vpKC97j5tJQZ5h2uOvPHN
+F8GMBhDRrRcy585k2y4RCg39cb6bgEBI2J6+ARjRjrD0hMycBfZAsPV04ruGXhR
pCm0liIGLusZFQFZrckuFk6fG2vGhmm4o5C6lJJbrb5rXf403ULcqgknocIVrFPS
Lhg6Mj8rtJb0pHF1vIMsoDV4yMaAC+PCkTi/UDt2YVrf867FR+CLISJwxFejoFfj
S6ZC3tn7gOBmB2YSyXxu1I8ZVAyLIkLenTz+k9OpeGa5shaNY5oZvX6KT4Rbdgl/
Ol2+zC+IDhRv+22daA+wRMvmPlm4HcMj7N75sk6ftgJj+fmm9GtOy0N4BBAiBUPQ
wyxD3T41fKfCjWV147IjmVFqIzphblPoxpTDrd9k2+OUEkRrrSONyAZI5gMzicoJ
Ne22fb0PtwZB+iIPi3Ikl6voZcHd4RCEPsO0lFk0Ht8cGFF/lcLtyeTxyyHh1EBD
ABCrsyun+aUBOi6fkKNcDtWquU5BvRtIBoQQ+CcLBpYtjCF7zFHa0Ss2vnXSxSa2
8mtmaRz1pCWG0upnWXmqtAVdSye8xhdG0/IVBqccpYoKGoR5VKdU+844rD+A1vuf
+d4nzbmSnlIn/MkjtlIOmAQkj7dDzjphJ+9a+GMpc0GEh9gnepWhiWoLTbPu/qLC
4HPZGp5Qx7aZ3AvSl7gG6ltt8bjOYDX2FEXYAxWvuWzO5Q++MoNsVDV4NQ2vXwBl
Lc+jbU1PAvXnApicjuWbLQpn+ecVTk0nUxFzct3SIXLkHS6t4qL1uVBzqRWhj6TO
vXd8EMz/UB9h2gSbRs4wxN/cYGGD9MTACLgZkXZ/ulEdlCVXAl2bhwdLWIh+FcMN
DStjtagf4b4qO/w8Z2HsylEZTbChmWddf3iIOcgoJVb0LPRMfVI/JZ8Ud2EMS0ak
u94tZs2s70jUvMGiCIEq8X2ONQ/wmvd/jD9YOK6OGX3QueqzgR+21wunVVa/tTqv
1lNw1G6zXE1CX70Ae2UlNONROKQ47FC17LxcViyQM5VLhiqwbpnAN8lWoiIkAo1T
KFSGH0Voi4Kk/932+d+zp7TG6+1j7Z1cLubtngPTYSIIuG9xWaEVq3lzyMV7JYKo
d3qbrKNcT0fUVUvxFykF+KZkpN19BMEtlt3x325YWtZTWgM3Sy/lrpzNtPVZZP7b
EtXqaHJL6IPjXL4HSbbPbVhVkjlexwHur3ArM2KTYt/Sdb6UK3LqrkcOF3zamSGW
D6vc//+LQnKIkT5jZA/M7IbCVusjXlivM204Qp3uW8DRsdy4WjLyG0bFvbASfZeJ
v48bfB1n49J12RDKJLShyK9y8bjEOeurATwkj2kiz0cFk4ZTGxj9RcCyMAfepaRx
6p2sG277EU5QRJ5TI1WJcrFf+fpQoDb43S2VYekRUY175KFx62HqKzByuUwVotdm
yM5Sw296JpG1170c+FbsYFQx9D+O+lf1OVJoEzY+CMZRn+yeJM0QtlTfhXzGZqfp
0dm8q8+6EPCtFG54jgVe7Sf/iYQhLGdwTiGZMdkkZ1vmPDqV2FmkxjNeLnlRWX4M
bwMwOdo8s4ppjFpNY9DnJZ4xNqJBG6kBzCMGBXBB562+mGYs8gqK/rwGeuwY2gan
WqrCZ8fes+FELG4PBT2b109qytf6ArI+qxG63Cb/xOwSXkJmPkEYuLruahwWv0h5
NO2Pm6W+5J6jyRSLTe5OPdUGvZHH9v2mXktogQSWu7/G+0BptgPp/ddg5WYnZWQh
Xx8h+2SBPuvgLFHwJ3QWRGdmOIGMvYmXeB4iSHxP/DqUA8OaUZJfiAAd9WR3v42d
K+DvE+InO9PGLYvcEmrwmJpUG9pq/BPLk+HYtxjO/GjqpeFbdvmUeDgyXterUSeR
uSckvgffyvGqy8TFPBHDsSlWD/DF8oaWL//kjBW1oEYZJB729A9bO5pM0yHU9B6A
pEch4pmRvlJ+PZZd+xa4GdrPC4764c8N/XdNR86FhpPfJliM8/FKcezUH092mra6
pmf2nIvEzdQsNB9Y0ssIh+hFm/FeVo1o/fOAK8HwKjpOe3TeFEqCjByEkQTWVlTq
ToENszQ/nqqAqvw0sGbN52jfUJ+ta+r4AYTM5R92QDokUP9zovuFAehVJIX7/gSF
tQcuTJ1fRddKoV/e2pqOjxK9KHKsTy02d/28e8qQ1NZtxf0fDIguAQZvNqvU6CLf
Y83HtAH4c9Ds/p9IZn5q+D0DXRpM4i7/zRVTGMYsRlB15p6sirGLyaxAIbeX4vz+
VWNy46AFNInNASuzulTcqAzzcmV7xDSkRbOdtSnQoIe1nRhIP6DHtm61elMVnnFY
P0UM+GJWNS3kaZcg++4hFfkNYyr4m+bfb9qMBTFWiS/aY+thLpa+pdtO02FGwQNz
GAGUh5dsSI7IHUFv+D/VjvpQuVO6KePDjHZ+R6jBaSQAuxtwi+vODwbT3PG1ZZU1
Cp4FSaHhh/VJ/o5dXhhW7KmFJuevNF9QE8vIvoDUAFGrr9dZUB1imh7Z25So88X+
n6ftpI7AwJIF8D0gAm6ZkyYdA9LC86ImJaeHGeqIMn6/aZM6abYwrcMY/xicIACr
TJid7UgWU9lK+4NNi+ytIxPKVl+x1leJu/3NQVn9swD8kNrDrN9Slr1lC5NUzzoL
cW3Gtxk3yZFBfIgFEB9N/P8Dfs5SM8xt8eAtBCLNA056b6cxGDEVeTYRsNJQdCxM
VZSrmUJZpUbts/+JIHe21qZZ7IXZ6xQEgMls7fYcdQNv83bRd5XYuZiTDsV1J288
AUFCYVEBdIGr8nxRfRnNxnJz4/g8PjzrMMRGH7iVPov3S5fcgRT6m/XCMVH6x+OQ
8FRlndHiXw7AdyA5aGLG2wk806Avcq3xtFD1duKjTdI9FFHuFC/uH0OkcLqI/rw+
u7PTRYWpe5m17icC+W+Cjs934qjuzhIYmmNZnziwBgXCPAb2gIICgV7DWrZs8J6W
Lu73TiFE4kbB2yPPAJ/R2efTZ/EpEBqZMwqg0i0HJ5vWfqicGcEsqZsNJ7ouFRAL
8CnuxogGrE7kEvrmBNMM8YrdrEjm94umXjZpeTPy4AoGmHFQq1dccKVTICznYHgk
Zh79tJiGnh20c8R6tR1CJ/60T/RzEdW/MqyRfkGy6EUz0RTOYTEQdyti1/BYmOmy
TtU0LGyF9t/vEen7FX1Ng2yjJLT30DBAf3jKJ5wmkQ7dRhACPQWUFSWUz1vOSbmo
iMKkUaO2sjjhGbv4NiYWtc7Pzz9L8tsfy85XE4ddE99k2wlg8mZ2L7Ccacjc17ZA
gF1kqsjWpdnXwVrlSc4QmJj6d0ldzZ18mNmh3xUGB4MaJxW1vk6X7Ns//SeiokFF
Q958vHSNJHegV3OmwIgSQN25tEpoGUdECs5wfHy/jIytBRdYF4HcWn+yUfKMxOYb
FbLdqOMMHwAk9ue6FjcNw7f2a/mD+7IzyQ1EzE6K59JCXZjFHyAja6sDSxYL4+DZ
xbYUSVF45KRQFYSSul565LrI26V7sMTes6ZKVXvaq+TMvf7x89oWQV5Ohp9qOwqF
dqwJAOSqaVXOOymzEuGqQs0Ik+XZsOC6HLlo00ti7ooSwL+Hts7iV2G8A4JDIEOM
CQwJpEgResqYPH3ipoAGTr7V5l7YZC4B5Vy0vw6wlqXw/zbbAEFrwn96up0dpjOk
DeafL2wnWrYzLm5geMYd3sMWQlgwcKD6XKiN6Q/6Du3jBNDkawFSXYwMWNuItZuB
j9CEXMHdFxsH7ffDCox4KOy+75xkV8+6QpFjgCbd+9a0fC0cAG39n67i32ecJTAv
RmqYj5sNgJA18yYbv9adzvgRBqOWW03GyTCqSizf6M4k9Ci2y8JbJ97uN/1UyNWo
Z5ujuqh5UFO0iWIaaqV+VHramdhRPtO6VJrF1ksm+losqyUoFB1YgRdRBOc10LUN
WzL8y6rtrgzkIb3izxiGvb1XrGM6/dXVSX5DAlzeCbm1UKRqEU7kLD/9blZZdLMr
rzPWhPu+EZ6riBIVqQIO23uyGCK3+zUTqTcSY/G/8MVCxh4gd89CqA+zNGbj6utQ
f//20giOIGrpRUP9BP7IkJzSIMT5rMZFfkw9xq7MZAUfwOSWMo56vZxaOcRB5HQ0
WCYBlJjgezDOkZXD6+un+96YS8ckxWRrW3tuNpNRXyTYHgE3nIUT5wRKu8s5mLCs
j1ANxrVptZfzrafpEQM2SvGf7HSAa5VtJy/BarD+h6LhCSjrZEECtW2quKdrMOFt
0MIWidLb78gRwx+USr48uD7w5jF5B4eqVNlRb52VTkJldPVXxLrSM28K1qUFkIid
c45gfP3p01btwQuWzGlvmR7eA1cKqxAXO0rdPEiQoyjcmKLQt0k9yFtvFaL+gHZW
N1ncw7W+v8AHM2RVKwgGZvsiWnU2ORUCU79m+Xu1a4do/qPBggFM+H4ZM1qXjV4f
UZiRINrrpXr2Xd+4LoLaeHQmOC/ugCeM+iQd4m531tIPQlLAQENznGrgZ3yjadFP
IvYiVg9L/nQmrN4dLnuy2U5md9ItnUyMb0N/t/1SLHzkdFUda7zs6yWohNoaB4GG
NjLnf/B0HLuk/6XQqAgm6wHV52G+CSFEhU05O9d0nuujlyeTztrungaqtOb5kPPY
+hY3d4DdPh6iAe2HHoTUFuQkoyXgzxJH9Kzv0SANx9P4Vx7M7WPnOE45V9ZVFucD
xmxef/Ix9d6yon2SEzXadm9pnNK1pDzTUFaEgSCuc2qAk5WJTHjrmYosB9Xn7S4K
z3NPbr+IyMQeLy3KNciODdrEI+cHwwMUhxs+e0oIQEGwBvGf2F6POaFAE4ihUqFJ
YguPGpuJpJLaoVkZ7i7ZVIUMtSa9wvNOdIeFi6EXYfgEB9J+b+R6bhvft3oqoiAZ
XwsUXEJmjS+dyY8gcGcr9qEbFxGRp8TDCNPcAqUTDYE0PGzf338bHV38R4NAIBIT
yArDIh8ecBnjS/UjMriMHbbBvXyg+O6b8LrtuaYyocM286nEU6K2sbF9+Hjcg/+2
uVtdHGqsx8i0T9OR+Piq/fThjzCAiQYpOkqZdPMAlbtIAo71Xn1/vgtvbFoTIcCT
G4YqatYWNiQHD7kPOHNjkn90N31qH5T+xyO1f5Et2GvmeW0/3vF8RYnjuctJj68I
ttE/26+daRCKb7Qxl0UB0938nJoh5LYQVxtDZRbz+xToahf9ImCbUpl6SFb5eSFC
TkTH2203KKs40PPPybwUwPivMAf30Ox7GtDmaSWntwkjH9JYJC2krLII/hYEZmZ3
RpJLYkiDuXuvtvaFdMO+Q0VGAzjRYIIk/dK/jESptZDWadPeXwZGco4OZflLteEU
kEyuwzLV9qq38wvIWj+ihOuC3PhJcV2AvLx++1Tz6pjLWXvve60brPLZNMj/AqoN
ptCkSC724Jz+FcE3fcd7ncQlzlQTzDj4L62PeNTcwTvY2X00ytvOhMBXiSevHfpA
S1CZNAimPc4h9BFY9bru2vH0+SzfrpG4dIOW0Dimlhg32q7ckq6v84eS020R9kxP
VN3cNzj4n9sEsy8XwJmDWOTyzwJOAXPncQuweO5nA8p5NKYG7NoAvTsklgXzhixh
f3Getkj5PiVxco1tQ8wqhPdLzNlGPmuFRMThRMR8lwWMO4rFE+IkWoO5GRhOYDMW
vWFjamW7tfvbztl8It3oiTX/WxWacMlfF5WbdnDdo2DvC58Yy6ffnF6kE5437mbK
uUlvHp6sn+J915KPZPl710JZs8AIXhDRh1xCILe78ve4kjadiqofVTwQICJfCzrX
0WhSuasPC4QTDZQTNBPEbCVDYpSr3NTPDpHF59l2inIXtAcZt4MJAqEvdDK3JqMT
h/hOHV5Cd24yYykoIMF5WQYwk9CI44OhVbkjSyZU3qNNez0jOfM7/wuPuTTrUIaL
GxR1OalzOSzTfCxPfyyS6IlyXNyidprOGCV1aJsQNlHFtxpbKn2lmfnjSjylGTzw
NyQaUhAebC/1HFNP7L5Pl/FR8paH0NDNf+57AHlmaWqnmEsQxTJJYRer8FD8xriv
NoqriHdT0uRw0kbjI9kjdP7IWeJvPg8y61KgTvf64esG9YC/tzpUOyQUcJaJFzD1
NNn8i2CDFqjCg2CUm3ufF0cNzkCb2qDlRFCe+xG2z/flPkkIbz/OTGtkK4zkq4JP
LwxABC+IjlzHrxOcckMLiOiw8ETQxCYm9+A5xbp8YxBEzW80SL/3V/atPk5hF8Vh
dSZKAG3Vs7nPXPMJ/nve5hqKCKnmky/xUAME44g6ah5Oq3FIPjPvEgBeAYBQgHxL
nS8mRKw8hMsCHjYL5Ftc+YaDV0ssnQ0zwE7BfszuUGCC93MhJSvcLNbSYlxmvSSN
Gqxn71DSeHndei+M/uMrM9y55LQIBU6wV0RZpLvmRROtQvt+7mzTas2JZAV8GsDu
gv7g/oCaQc807GPWx25Ox+r3PSREHEKoS8DWG9y67xquksCdaY7svNQ1Urqzu0Ft
esdIqGzPHQ6ixtzcq2j/Nm4LT/6SlkRFH3hG2dKvWHs2g+YyK1YhfKWfCLGbvuLD
UngtJTFc6a/EEY9uAVjblWdt1vEMrZyGouznEpUsojqZcUg1dl6E3+24UhBI2YlL
w10QG9XF9/wFME8D5l7lWGwzW/Zt17FkbB23TUXaxwU318mReR334bSupe5k2IzL
K5Ov9e6JYOBdLGv9dk1GD0WS/rLR+BFwc/WJbfRwzberH0hLFcK19cgfSD2osoqH
5Pc/oDAhOZv8JiV/NI1xerW2aeMarWX5oACG/bW2AdYUxl5ucg9SqgHo2YdJLwDK
qoyL6NtyVTOp2CM09M1/gDkmntKFqfF4Sj5RrLVpDhuPJiv3bGjf58+iGRxu7Xjm
O3qW/uDiAUsDkOf0qQChsn7a8dgj01WKRb/LRGbliNEWHYDk7P/3udOyeNMyw0ns
Cd2ueLVsdeA3Ly4W/1XHZInQc5P12AJ5FzcpNraOP50iGO8KqZDatRpw3tPC08Ju
GtY4OADyOrhmdsUrlqZdDZCnC8El3RpgWMZhRZu2fO6nGjRbOk4ofqGe8FLha6WO
NgjRLyH+4gUVSKP1xH9Xb9+G2r5kX0PYdAxfwSS/HWpEk2dYObdRbxsCQqMIOgyP
AFGh/Q6XKIxUo7NXzHTDhGbONDDX96c6YrvQxSQbw73q3LU9J36oyYQq2Le3eSpR
laiujjb4Hbp7qfFoBbLbsF3qkD6mD4pVq0yGO6AhlAb4xB8WxTuuM5kpElSPYtdg
q0FCXsvETVsbYxXL02Ur559YLva2EMkdkUAGjv2jteK2BVro1lBzfOF7jJqBlzwH
Ph61aO30lQ5P5MzBiBaSaWiWfjBxxTJ/WHKnpAA8K7aq+j24PaT5U2BZwOnCZPs6
NazQ2gM5cXUapig/GMqt+sTKdWELDw46jE1u6iIW3aSWRh77OPTPgPDQ1eDFDP6G
mwZYvpOFA1SIUSMo3T7qNgx9Wt8LMGaRdztQqvmOGh4aMm02HNf2uZ50VhwbB/Tj
5f7WeP9CqtZl1pCT7aaGXVfg/25fgscY+fYDMOpiadxvm7ERc/GTsVhfZ9IpyCr+
ZnyODX1QeZOVcLfE6KM5JgWlcv+rpMnpnpnAoWZzDdRhyQLP8j3G/0eg/LpGoCmo
SJlH7/n82oAJLFWvUBR7gr2UwGcCucLMpqitZXRTyulcTUsBmaT70DovolstRU7Q
A22pJQzFRArn7APaWGfUHLL/DBeQ945/J8zN5TLGj6JdtYP/An6qtnS3BZtxH9UE
FPtUstat0WeDG8EF64xp7Vr8G2ojlDes2UJy3Y5Ymsba9acCfk7TNLPWHKOB9tgq
GkY0/6YjrDYfz1T84HGhH25G9gcLNjIb7Ujt8rI+MsZh8hymha8G+00P52awYGMV
fTWPXgAL+ZXoK4FHK2MwTJdnmXzmSTOy1Wn6ixkB/zYj4NuDIztcNUO+X33LtEFm
OJt/SNfB8ktvriVc1bIDcZ5KkkG46Iy8Lq50tFyi/F8+E3muGCfqsP9DX9JGWVQg
D+5IV2xx1PPgf+1yBN+4tZXuvzqhgYJyJ/Ldaw1jNe6GlpAC34N8sQy1O8n5+66r
YhQq7pJW7Le8CnMkJivmnBN5vLLMyobdHM+5tuZQWQvGet8fuGvgEGhYfUHfpEkC
h78glsgkxVpPPLuawjXN7RPqhG/QOf9kwoJuOkThMA/Z05+MmtLQxBj+M1r0k/dA
zN+E0NPW+nZPgKctxLmU4jgtGdihxo8exrggtCN3WqmAGBGBjvmtv1jCY6Xqtexf
uHlWP64eMqC+FA25GQTxz75+jMtpu2XppWkGG1spzWdUycPbhdDhlNTsFFeApgsf
tAadlIV+zp78XO6HzboSmWUTBOCgYiTVrbSrDmcwhGSoaUuxsOaMVf7LpsyB5nO7
MfGqVmbmnXb0DZLu+OmlE86br3pBaD6orB+eg1Fz25p87Is0m4W5aVfWDurtbTdw
pk1zyei7tzCq2npN/cEXZnCKn2HzNVZxe6PYVcYYrHBPtEFU0alFDdDF4deTbaKd
5gPkFyAmlK1+ivu5eN3F4nRG57Ik9YT7LfVcD75SJqOIQWhLo8cmpHZIEcmc5XaB
dCXS6VIMK+yeB+Zu1eo9q7u1Q74YoUrz71iMbRUqqGlKhcuQFGXvayW2afxTgFIo
mZUdSruicjVG0+CI8j/DJBXmkm/44gq81uQ81EF5lRYjP2fy0jBfjauz7Vul/9Qb
1lHH6AVT8QPsP4BBrDev8k5Js9L0oQXYAafNT+EwE3ecVkf7G+URYNpogxdwGd1x
8ifwaoTUDmIHy0ttPRbOMJ+wzdL+pJBHBuAv4M8zyqOxtvC03NYlgCcWFJn3b7vi
d+t3DZ2PR0Plj5rnuqWR134T7bXsAXWn7xQ+CIuHtKnNUjVDgqKbLRDL7Q9fRR0s
QsM2263+fh/4Q5cxDiThI6EXEpJK+0OcEPN1/dmeU6gIhNvfHK8QQvR/7fa21GUB
+ORPzml6eRez4yWA6GzKLlLb5/597sQXGOAmC0mDILTOb+Okwx6O+pacZ25eoTet
u+bHcB3CDjsNnKRKOulWxVDyYV6TRxmNfLWH/waVD+i8GOXU9tEU+pWao4/gzjXk
bJqCBxqJh+EMOthJBiBpRxjqkI/y6RKXd5hqLuEGn44kRmeYxlDCjIwWQ1nRSHSL
Nx5n+RHVcIVxhNgGitFd6NPeYq0HXxG+8tmN6Frqk5WEA0ziU0x6/szWEuB4FmFY
HH78jv9lkyADjIh24lHGcQyFkmaVgtwklXcEnwQX/15P9TcygWhKtIm/c/FuZ6UJ
w+1cvunV2mr15TpFD0EMXbGuNT4hSeEW49DBCe+jGh4TAw1DzWPIdzFboRvgW9YV
vnS/T+DIxo6nV479cE3m2e2OQN/G3iQ0/CsEIuY2bzRxKLBWO3cwJ2Bmrqpp+nwW
VofR8QOuM/0dTggscPMIWhwDauykGaN2n9IlkC6CHi91VK5TUoyqz4zS3LphdPU0
adw3+8SBqRNuYbKIQ2Q8qsZu6WllvX7T9auubp52cjsJcZ//bY6yziEs0CTFM5cW
79LGArKLUbMfc5Uq2ZOGq9jwSM0s3oRVmnuAHgV6fm3KfX5usZht37mo91wm68Ps
rr0SGodBuN6Ow2ZMMn3kK8pgAGWEjM6xoMfS99e4C0gVxOHSWzhzkQWAHyvDZcRN
J11zDcZDzNaeJidPQVW8f0VFO3IFOyBFb66FT54kv70USsYSFnxt53SEKIeGb4NP
RTR6wex8mRc+ubzqJOIk9wrR+7uIyOp+pK9CCRRnrhnPS6Eww0ZYg0oAZO6uFbxO
SK59LyXybLd8hSZEF06UN0xikGmo4IhL0gmww6mcdMoJK8yWkUMe+PxWgtGX89JI
PckNumSgTVGDBVJ+nrf312or7Sc782++xdJgTbHedRS+UXDq3c/kIb/dw3p2Hq9g
CD10ihNg0vyQ9U8itb6uxw+zFAsAFZF0xv+9iRbfkdm8zJKNSbPaBf2Al1qJbLr7
wYeOlcKlZEzLWmw21EC8jcdaXANawdatx/ElMqGM94LYX6HBQHebuWJVeNX6L8XZ
7nmdLmKSh8+ss6ajf+9jhQvoD5NWvNaa3nhfIpBUDOUPFnEC0i/1E3RS3pIR+1ZJ
8H/vA9kkDu4Ie6CZEF9+NFjaeBcDdB+Jf7RhGGvyjdRARfH5WRc0ttM4HoDw/eQG
GV8YGN21MBRSwIUYAwjUNLtSRQSxUg10UFfeDJLJr9J0UmH1AgYIHMufWU0ORyLR
/+rJ8RX1bjChFoCafJPUZVvGvibSsjvmpayK2c//rB0NWrnutpcS192xQgy/Z7Qx
YEcD1fFpXx1riQNepWS7/wav+S0FS5YENeo2fnFFU6OMjrCpR7eRV5oqCkAcaL2u
3w2Kz24QxUFOG/S/dSd+ftjLekPs8iW6iRDeRuz2gz8nS2JXCZ8N5kpWy/4a40Vy
+izYdvhHOBY9YhC4/XKC0abcPk3BvFh1bWaSh7ixaFVEZ7nNTB/XKYumUjsqrgGS
/n9q8g+c/rxJpT4NujnzqEXVslLOy6pMXUsl68u3NUbTxYw/zS9NEWXuH6zWfWF5
asLRcVs97vQaUaJTZV6Du4Dq3hGlcM46xlwHlgDA+fIRNUNt13JSrCBy2ZM0/bPZ
Kw7rClIn/ykKRBQp2LRfu7wMs6APULLzj+Lh5nhor8eia/bae08cv7pUB+uRbRZc
KsHWbDBQwOx7mBYEs9WmC0WLARF1qSyX/QV1SAcJ10xvNXLhygm1s/Zq4PLWpm3B
VXyeCUCpiV5ECjC1A5HxN2PgZhP8VjpxpZ+Pa80AjpbIxN9JERIwWqAKKxXbCxc0
NsSOXOstyIX4xV8ztkvIbE8M6RGzRqDncw+G7c6QiDQnfb5cdDEr6aBFeCxJtzl9
qloI+s+YuYK3gdXnjCADElkv1MjkG3tf83bSagWyk1R3udsckI52OE8G8NAJewxw
x+equK2KysMbj1DKBcy2yqNUf5Q/4zSVtGmijQYljyvXnh5TMWPeSCVQ9DmfzhqG
J+0YFf+dhWVY7FHlIH/QI5UfNILooQQBz12+aSBfPascCma9rzd03DsvC4+keGqh
NGwcyswfO0HS82x4WpkeKVWsi1aiwQJ/fDa1tqjQZ8JSFUQoIeg1mlp57rdjncAL
niMKT6KrvrwGf8izSTYGTUm8x6balrRYXypwLC+fNA0vIrkxL8zH59hoM54Sm8+G
w+WpMMhMYvqchtvWn8tyFbtR1/eY42allXI30JFBJ/1kkgX+uoerjHF6XnWJTu0+
4bsvO+03r3fjr44p+PsfcDYrvzUtIfi8QDj56uh0vqBDzxqXq1tnz0KkNMd/u82n
5VqE00UGEG8vuLqziawewN3UZKEqA4KHIZW4G0D2J0hL5JP5uNAcez8/0k8+NgUT
lpVJ8IjLwbH6NB65e77i2oGwzI52OkPjFuQOLIGXw1aLhm4QTIyIKMx+ur55rK8T
pF6iNoyBZ0iIy4aRKfYY73Tb/8OmUzKLPy3hsnyQ8qDqFp6tHUjgSnsjXw8srGoY
u1HPWGhmUVhte5MCnytmPEpervkA8mANyErrGSNqV4GOe6i8UN7JjHqiGw9NYodl
+sjZ7ZzhGfSF2hx1lOORvjRvHp0AHCTwnFw3MfA+jAqjju8HE54ndSMdQbaa8Z5t
QwqRnC83zMQw34/cOzDSxlsyHU/abfDP2ENcUrsGpTBKeTVy+9/0LIQDyOBD66ou
+GRQJ7mLkcNamn8zHdTqyKesQ1XhmiDL9p3W3gMRDlh3peKTR/TsC/yNaTMZ5vXj
SnrN9RpRJHxFbISHl3ywxWmyNkcxsqlIBr8mmvCCJ2HkfOY2RVfziVNJatVhuhFk
Q/JV4Y0gHGSe9ghcUm/c/FISvaurJkMHk2AZ+JxfC01CZSbo0LgT6eCL0PdzFV4I
UOpflx1sG/uVMS1s3EyI0Gg6mBgemvBfUyLY9ocR4752dPpi8uZyNVbQ/PVynE9j
om/1ZLhesw3oK4obGKd5kcYJueejp8kVlEVvyf9XGtQAp+QnE6aZ9CiNJzef07ZQ
k0Qz+x2vnV0FfG2YhHj5HDEkUIKLiMYSPB2jkKaE97Dr3Z6ZrJDwUqgiladfGzn7
7Bdt+ve4kJdpJVdN12qyWK3t7YVOF9UcNBx6P/9o43UE9Bdepm8sbtOFLjtF/Uom
2F8/k2T7fxQ5dPB6vX91Up6BW0z5FD07hFXaYhk1J2lIDbaP0WjnRWHEaZer3LlR
vqGhX93ah0+Cy7yLzdD50tWVSChideS8lCidk+vNBp5IvhRw9rm/p+stjgU/WGcZ
LbEi5BcImDgx+E8XeVhh+wqDqcv4902tiLpLT4yTa+x8oIfkK+y5y8FmypRwsety
vDbn5kp2J3htzuCnU17UHdb0OQpa3Q3vHOddzrQHxeCrkb5z5iZKGQxJKS4GQ5ST
cHkPpTX/pFRRzuyFH1xm6i54ma97d3qb8KtybI5wAWqm93HZ+hI8rrLq+DIfxs7J
0GxK6di2tq4VsUfMNBRQRv++6RzQa3+GUc7+SSQnDcIxXycLcZOVWOfIU91bfbBv
rLuzErItMhXsqJLRXJRKWCS3kmp8UO6uOxTTE/C4+H1QoQHgRnO2kQWqAFzVPZDt
BWtAOiAn1lAd2wpA0srSsuFzqlifzjpZY9BnqDI5IcYSiPOKbWZGcuibc1oeei4G
XCpybcyX8FsN8rNesot/EoF3CU5dZ8GpoKtl83L51YAh4AZIRWEswQS/o0S+e+pJ
UHwjtFM7nGd+xJduo4ThVunwhoyUxvv2hceyLG9SKgI2AB3ppVCaAFre27j3S/Ps
TqXHzmgC061CvYifh6X+DlRTRYe0jI1Oodi5YmXevfzMWtKNZra5eLGZbGZ0jNS6
52L5+3SZBt7lopXSKP0ntr0UGwCUnoeVcq+L5UT5mB3YgheS2fJ1xa0yagzjtmfq
rmZlTdYeuyauRd9BgfCOZ1er5xHNvI12pbs+31h4NH+32zDZEQCJl/uZpc82uYc+
My2TsenLWFz3rgIdI9KmlLVH+b27NHy28zpzd85fhBeEut6MmzuMg8XdgK5HTtTZ
B7CEZJW32UeI+x2TYzQnyReS71PwJkbU6EDzymLBNEcHl/oA/qEUWIVPVz3pCgDs
Wdim1bhC16fR55m2TCudR4eYj1uIAMy8mMLWulrRgO/5sFFzyTSDsLAL57uaMD02
kk95Zc+sU/xgmlCLbGdzgiRN11i8SLmwiRhulj3nyi/jPX6Yp0eEhsH2PeGPokEw
OcovAIXHXiDwkcYL5v48VXFUi8t9IqmU0arVGJMLQEHezy+lwJ6FOCpHKVrgv+fL
92BgykLTFkvIS+sLBlBYQmcF0zQvhLqOrsPdSKCk5GUCvJl6Ur8sGe9NSS0tYMPl
pM/Yegmob5T05YOvGDwfpkNXX8VT9reSmry6gMqAUwlZXcjICYTeDBvewbaYekBk
Tr613h0xiDwKJW0YZSVxk+S5GnHlDUX1jTTSMtnm5lWuz5xy0+3S6nSIB+bvZPpm
w1aPmA7IISoJkT3IOHeFMUN2d3P5U0s1fYr0sFR7NeWFx8hyjrTjmbw62xlADLJ2
B6X99eMHmBefnAaQsVd3gTqZmsTR0YKynStrYOjRzFk5BJqY/9XSXipsNaXD7iGk
jv8NQkuCd88usEiyuVD+0hJv492nO1i3O9hEQWbtZbNyWhfuIUZTg/g4/y/HXZ+D
c9AUHa7BHShcWp3CiwwspHFbEuMQVLHKsBT2Q2uMjzaynE6+yKsghprXIUMRs0rb
t7amaJsul1ltpqHiS/am2BHMx8QRQBObXBQXRqeY2LxNswGxTCWmKTmwCW0Xg8qZ
BUAWw6mRu6kv2l1ptLFVHLj1tB5Vunczbd0NqdkZtTti/MqUe4JZetqc+whQHiCx
QoAyhY96c77TFfFc6RMrTewKC/9CVlmeMBdfMmvDgRtLMY95AZ78wToWVbdxnA4D
d/kjw1EtBW0w9XqimLrLrrp9gDGFuKDFc/x2cUEaKms8mLFdlLHpfbUfHM6AYNu8
xc8sjdL8d2okMjPEjhiBE7XpuoytxfOWNlyb62tIr5o3mdogL3f8uFMNdgNGXD7W
z8m66uQvfFobT+48vlO7d26vUMYzKw3gY0e43Chq8n0rswCQpbHnbYbrrqcZVeYN
4BMWAcTGKX1PbU5Pao1HtSwS9cgJNVxjE0CjXOP2033WOADmd6OUw9JQSz1sW4EG
0Lfe02NKKkZABSMdno/0fIr+arjS1/+WxUlSXSt2+tX3ZijEkkG7oMgqU414EnNk
eDPxwhAOA1YOFQcHw/1Wb6AaqEgT7538Cs66bg6u0npXVOhUOjC5CGcIvrHSW/LN
xyvjz31YmmV8RqHQE1MeacTPhpz61BZWysWHWc13HzxF+RCeWStumS1K+Bf77Tbb
0T68ttqjZt28RtDzOKaYca85A8T/qgSCmGJoHE2BftgvfFvBBz3pDNMwNqoQ3GCS
BFej2A8gEDzOW1lUARMW6/LM2H1I83OZ2QTl6Cbe3rivFjGnzIetLsOyUuuOelEO
enMQrWBu0qBcgf/4NOGfHZDeEMngqOhanfJIKgTyWAwlLrZgeBmdNy48UP/BsrK5
yjej+PpEScTG1M0ig6Eb70HqEkh/yC1ygzioq7LsTYhO96z1u3dvfKeq3ztyiC39
KQUuPEtsg3LEZqBpDiMWNVOjj9Yv9li6+AVziF+q98HyWddqu41W+5cGkkte5Xs8
DSAWk0ftKW6ayxtdr+F6oUr9JTYKoZb/i+rtymOPMH1iVgspd0ekwYdPNZ/hEmm5
HVg8Z+ShY6yajRkCEsAAzjWJ86nvdyga5OI9MziTQ5Pq8GzfKN699kGlhq5Qy/Y9
rSGsENGqSpOMjWzTyWVl/QkrIKbUECid5q3M3PumtuYoVZTRfVwS9WOtYbBiD8Ri
6MyDCpPEt1dRiuY07dDNvk8vO7hGiHkoXtX9B2uVRo0gX6LgnY5DVmLLVrQQC1RJ
svWGa+VJFnTQgdxAkBXbfhNRB1O+2lfpQivERkKF03hnxmJwzM1EwjCMuQLCGd96
HrUqlMyN3mRGh3PTJbgkuD/LCCjaVasDjEEz4a1Q6JPccH28O9ZnaYVdp+rhjYDJ
U8qJRoz/Tql44nJF+giHqtd51PXFiETzWvom6sxS49ONbxGNI0C3DHzwv/C86tV9
2f6QZMTMQ3u2PYphJl+TnyyJbezvlHDthJLXJONQpbpzZLLrCEud4MsoHhrmJafJ
DIFG7JENO1y7wKBJSNYlONGCbwB4F/i03IwHNBufEcbvPnClEE/cFMhvnwyaLYW/
lwQ7GamEEE+yXHdVGYZVSWc+8WV5o6HQ2k6NxEXBCqTXG3F3Ud5see84oanjArbt
hjjCrppziKVGK7uEbq88QHedLmtNJ2RlC5LpL2CZ72J7mTFvDOCiV66XknyQ+n2D
7LLlQyvZPuH09SEoH3g8S14/+pdMxxYNT/af266j8FlBkeMGjs3vu4A4F+sWqrH1
5mRdm5QKOEYusjvnM5sodN+9rA0rXt+rU7aA9tqRt4hvHXgOvHlqO+2uIHpKTv0z
PhqgspmcRUM5IPighgHGXOp8/upCw3F7bw73ubtIRn/0MevokaUAPM2I8N09u8wL
gFbsyM+CcUQH9+jxvdYrzoDp5Ac9q3L5hKk4Qv0JB2EFqqVz8dsu1WQ5Z9tZT67D
AkjiBMmcrXnSmXC4ogwCq0Fs7A1iyQpCFT0GBM82iDY2ixmqmsyGW128Q4E3OC6b
pkNnfXyroP/BzLntO4fHgiGHSyk51Ags4ruew80OT6Q1a9Py2EfeTAhWcCx6Zp5f
kP69tWbC1mmpAUbra1P63amoom+NLSm165a/w2g+GX+ZYi+P8q2497ajKw5bgrst
DTVjEkN5MpWSax5n7Y91t9IyVXce+f9cDx8a7BOq53S+dnakx3l7pmj89dYNmH/A
ttXTAMm59JeeJqlYL2/g4U7yq8+7nq1lUfAMOuUh7cPx5mdes5Vu/tu8tVW3F95x
IsSu1vptiCdAh3/qTEXCov19qGprWxhoMJMh3QsWDI7EBTbazAFiMRioHb2nQE8s
r7CkFn1vBrEdd0M5TMKChWSUewNz79xmJXnyt46UwOB/8Zyzsgeeb+k4oqFLYCLA
APnLgTqVO1eYpbYfFCcBmsn5b0GOUIOeKUp3Dv7mRYz9cBU7nrvw1vpvRFP0N4qV
5uwBgtvBUfuNo3w5accbSDqx4XalyM8EImlLkDW7bRRWQuUDLb31MCsIgi7ImsXK
i4XQtQB4xJf3o4mJ7ESk4RziLcDhFq8WeAKELY5iewoClBD+VtAcFHuIsH+o6Z1O
yxEtk7a2aOzi0Ad2rrwxA4GuOsn6faMz7aflDKumZ9sc4UiZMGTLw3jhskkKsJdO
A1DaXsFbYdJWnT2GS8/u56o21QcaMDzh0EVNAkmr3pxlrktMxQgiQBbPXOkNbes3
0hv609SDp3FKvihRvrQSDhpDj8W3PApTSQBvySxNmHWtiEsrKtHbssbNoaT2QtjG
Wbr95mhDsx5ktevtB2B0GLxNMz8A8xHb9ktq131kU1Hu/lsagWxAddlVHwS5teMr
RYvJSeBz2Xx2NLrEm+4yerxcJHwglPo/lmG7z4MQjdK7HcrjCc2s520LhLreoPLN
awAaSc1RPcxKGoHQ6ZqecOKSQyqCxqBb6SfmC8gBcokaeDX+5VHtffgmLa5FZPPV
KyhjxxluyKiDxN0MXV8CfhBQ1cD3ffS5WAHXopB/ZI3x+ylVO+dpOHMrtIZ7VoQo
z3dQZOP+lwrYdrpTYO+3pmxweA0/O/N/fhjsNO/MO7PiORay/1GgdE+ZzNf4PIbX
h0uI+VPahPPdLO7mCkwQXiI2e5F7wn/ua85UADzkj8REVtZ+wLNnK+9W63x+WGbQ
thXGICLsyIXoV1SF5HHb++g29+LKIOEOk6493kfaPXY9VJS+rpZtP2HZsAjTVrOR
G5FFJ6eLhqjsazaa/2E+LaPCIsRLOSqK3ySM3jVoeabas9kX6yQTdIJuUZ+81BmI
QCDZCrdaMTN3QxpxALFkoXNMNg4ccqkrK2eltU7HAFHBPOVYqbXNXO6keKJ2XRIc
BJHzf729wfpRkZFmZvP0KLGFHy07iTY6CgfKBw6K9rBgHc3lzgvtxhWMrBwsSgwQ
v2oZfAU7WPwDp/42198NRm45NGf4HKsU4T2aSARyeMMOIfCX5rZmBV2tgF6iXAgl
dUQ92sKbyQyovJz7z9YwR6GfSzm8gkVo9a+V9xEh6eiPlaK0TJBBKlU7mDumweXC
Dk2GlDHG4DqOGgrZVz8fNfXAFE28XV7hK9qjsbpxjyqnotWqPZla5whVKNGTxXec
8RN0G5fUuhxSWF+2MJFy7fsLdMjuxTXF6vl3TFV2yA4k7oUj3eykgJzio137not7
PVlqDDVo/mf+wUOmm+Xiqlx1qK/hOUq7PiRORM9cCpnvAYp+5/RHPHQIMRQ9GLlW
SzZKU22A05juumIofSPkFHTffg9OWGdFwlyO2MZMTse4dD398x+HaE0rDgor7gOY
eLJ880NA2KfAzZmIkVpKIsreGyqqxFrqzFg3xkJgsf4Vjf0iOKz8u9QwkcEqB2l0
616xjkhSM5xedA4pUEOD4q8G7r9iqVCkA6YTXS/O/uIm40Eomtfi+9VyoCm5TqH/
DFNQTpcGUQHHYWhgtxgVz/v4TA96wbZSlBHEtTYl4KeTXReofYtJM+CEIAKsvKk2
eaNpYRA0n8TotUZE7ArWbmD34lj9Un+XqwBEwe8USElDMxueAepKdMSPI/mm9hwt
mND23jM9uk+WRMAYdXw6da3KRrLjCdD/GoZhvgyfbTcGSH87T9H1ECxEQz0lCAvn
C41D87CiDwJT7WTpl5smo3rjjluxv32XghBJLDSBaEzXeF0liDG9AW0m9bwCRX73
gcxKx+FjFprCHsmbZJHxC9Z3dBI0J72Lup/0y8dlojRMTSsGtLzSh+KxAUNtc3A7
hQra1swf9qB2ECSo79LrkotedkYKfRDb+EeqtHeBaRhVNC02CbU/4WZD6JAKScGs
7dcf0DZUPh9i0z/nDr/wcgcclZtO/iJrffaIKoqMmH5jRvk+Utdm+S/EQICGw7QF
eeofQQYRCbtupEts/P18XTDzMxlOhwPtRKLsjkQlgMIdasHEgWx7ZkYKjPoMD+yu
hQUt1XxSCdaew5XzIESRhzBB5R8QX1UODGlsRmb4sJO/reKSoOAy1qCmUiPtiUpa
fha/egbmIawGSUpvTLSKn63cIO4xd8niVUBICrR4a0lUMG7noDEDYFP9uE96a7RE
4ATd//yiJ3BVND6fdyPH5Dm2EFWBB98h3WDu6NtQD0XJoI64HmkBwFOpdpTGBYlu
O1bnielH7+FwnsbR13mdDRryoMzv8JrF8Zq9yx8l7Jxhls5tvdraASWPt6H0kLGP
pQJRrP5aA9fRZms776b3mXFFEMzhWQWd8PgjXyGyYAVz0cfkVrEmRRCPD9Bjohtb
rbCJX0Dw4OuKT2hvO2zWsmRWazpI8MZS3DdOjiGl65W9JJzNtT0run+s5kMFl401
b36WXt5M0HhwYm+lKNgYeUPjXrre4dxZdt5ThE5jTYdEQvH649WJs9h3DELoxqBP
S1Fu7UTEmep1afgy7EJsVcHzLD44kQyKo+Md4LNfkNShTpfWM41DxkF3iOl4veYq
9SRz9n857A9hri4/p0VULjZa4Q0Q3CLhQdHNQfope+B1J7buU7ByD+pmgk+xR5jW
0uLdMaGoZhPMfUaq7v4jCZar1d+/TDHIlKVhrRkOo5JysGkXpAgIZiwpp9wjQM+3
vUaDZn2bXeTXfhcP6a3jqV2hKVTNx7lSuCc3IDMpt5icMp1wKljCQEeiFJt1WQ2N
XnlnTbmsFqkPy0dDqZ7/bcFnq0q3bASr6jOM8XKZL7L56Ow6i5rmEzJe/5UANxw5
wt4buvG0en10Hz16oPkmUQwFp34vtdVYLZFtXE5Pc87p9/BRe7wRERggDYYIkdaT
jrrD9/jRvhM6jpjVWaHiczwHzkST0slUabLk8YA0X9jBtKked1BX+94++IhF4SCB
c074qBQuNT/QEDVa70V3eeYQruMHpXJbv/dJzmvsJXbvS7Bi1S3MAsf6BU1lfWxS
4cSconjeLWbqCVl+Fgt0XVjMgHfoAYpdVK9ps4rSZ3E5Ak5IpQMBg0cQ2C1dTW0B
OTkc+YT9u4VZtx5us4zqZ8huWqSgIs96toq9Nd+GkDw8nhKMWPi/tJ+mkFBQb2O2
oDpuItkSb7P4O8mumKOSHHaUYspwtgi/hPGf8KzmXO6KceAk3H9zAqTwIadHLSI5
bPQFT6xZDahcusHcFP3h8LXmSJrcr5KulH2YiApoizxRI7Ej6ZvfALv5DGpfE3g2
Svcp0PhfnEpWJS9zYxtIQ0rm1FV4dH1y+BQdYSjCTB6nOkwHPeDH/GBHkZYVu7cV
hRaIAelfS4o4HAplcLBFZa8l9aTL/3GLwFPsAa4si59kisB21RAzjoaqRlxCSrzi
K4edSFNIbqtebzaLKNif+elOdfFhvT54C7gmFpXcYcrvgGVsx/B1jDFikwYdIeds
aPEz79Sao5KzVfI9Nt/A/WNXUEWZ/c+p6jg6TonbMJDeZeGfnlY0ODQjlvL4yBbg
5hxWq6F5Gm3zcMPrpAcu6g5ds/biSh9s2QMvFRMINT3yhnuOkAhVKV6VnAzysT3Z
Nm1mpqIcvUiIHHTQy18GVmeN7jtIrD6Lli9Gpk5hwklLi1/48rnlCMVyJZWHHLkF
/2W/vExG4VllzHsMLZwVYhuT5GbgPZaEW8hxSqbxrnC0jjCQyAoYytFbE6LfO5im
izwJJ817SxCE/A4KKGbwYNw15ork8zFdYX7jvqhlm+lxRyHQNXDPeGi+tvYFF4pZ
GVpy/b+y68bs/T1YIF+2yMZh/9s4+4A+2qoTRBWvMWdAHiixeBr3kPLwsEV8lObq
mZK7zG+VxQh6EFQaYxTimSCSNv0mpWlCxBrafTD6JFBspQgfu0o2SfEEbD3MeNMT
bJqF9uBa+WcmYH6gjOTpXV+6BNLZzeFkOE9J+XPCZcMYhnPhtRPbpKOlYK8sa/xa
pvpOIJ2+4Y/AolWv/z54cWxLgzfLSWyu9OlRWl9NOBkpbPXxZI1BK8HHDJplPED+
Tg3iRQCOsd3Ha1tQrvq6NBs+pR9dmrBQpXsqu4urVgvKWOrmOYbS/xm4Kmo1Vslz
yBCNbQW+X5HcEBSI5TcMc7FwxEn8/+5ZWYywNv2gsyZw+fOWPisrIb18t8htM7TP
aneuWD6EwI0/OhgEgojhfHuXVg7pe/MLcyvmaluhK1/zjrzE/0lV0wJN2b3Bk3Lj
NNSrHGOw4Ez/Cyj0FHbuwi8dR3uHEukS0h0rLmur15Xw8KSfbvgC/98Pf4EySDuy
UK4oi2tMM/1oX3iT4oNtHpRbT6jydA1YLwwPsowKyGUPA0YS906Tv6bQ0IiWNsbt
VaKDkJrKAF2XpLSvGeNxqiK6CcDF2RzHwhrw1j8KOkmQndsEWptkzrq91Fe/SArw
zfO3Vy+U9UPNjHxCfMl5DA==
`pragma protect end_protected
