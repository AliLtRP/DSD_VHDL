// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
K4aEFNC8KzmZ77e7qbf1pdHWElHcJqcEqmwgHsfIBEqvMCZEIlUtl5gPrmKFNdK2F2uumUgDTjJK
A85F1t35G9BYBITpZYr2B/cinsnMCqZ6jAuNnirCjL2o/vMjVne0lby35PY2oxyzq1TQgHVRCOBL
09hNPboP3gTNPMy/JxYPv2BkijxKBoSAyC8pbY9nuR3pwvKhGFwcjESKDPoBpmKHlzU9+gvpIvoR
bJwqy/a9GfgzGrk4g82aqIowjU22vUhfom4E+xgWlfERvG6Kwuh9o+YOq8L4WaW22kO9X7MlRBs9
5AMJAagoJ6f6qPsP717VmrPqwv1Lz2LyykZdug==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
ny2OMbOMGHkapZFoFVeuJloayhDchQJCaXJl8jAlv9cn72TNCnR7KeGMOP+zgesk6P+VmMLoNGnM
mr9LaHWx8FBEzscskG+ubxGOqYj+inWESnaJa2xOBSOooZ5ZCuV1rgBoAYfDEWpOMJYROzg11QSQ
msQvOIA+xSIMz6ByKYjO4QKz0PyHpTQx/faX9eN6hEcaN9sVWxCKSCR5y/Moj368CNfFgk9c6LGy
nTtsp+wUlJJ45zvaA6bNHT0GOZdF1ury52fsxgefe1VUcISuNDb2TOcdzwrvZ7yrOWf2/DxHQ9iz
gyM1SL0+y9smy0uPanFZ+XRoVBESBCg1bbiZ7eaGwTRhX0nEUnDZV/T6JNO1Wds1aEvPc8WT4B1K
O2faIBFEHRscV8sVojEgoabeMsC9gzwlJShHIjJnlWbZ06lK6derNWjwvlbL206iC6GT3phAzOdu
4jgclx7cuCcHxaxLHHvr4ueTgkfX78ojy51OV4pg6EFRQlHdoPvzKYXXLVNRd2lasC6rwSwRSqZX
KSPqGZNOtl63W+nQgHJM7uxma0pKAClQNEtutCBxtdAEgklGyR9LdnSYpF+sKwu8H9BU93KF8cQm
X2eSxFQwEyRdAfdgDEK0TL4AOijk9lKjqN0MPQrWzODGM9ffvnzdoU0jQjLTCXkZ5DelmP0ZotWR
3px8aRlTtSn60mG2k8NRd1FI+b8TCvtVSYabhgMp+qbeuqN63XAE34m7vFjS/XS3KFw5Qr3rqpsH
pMwD4R6UdO+a+q2l48IoopIvSdR2ZERDIUGBVkyLLmvQfML9HlJM7uiaJmuOfYd18sSFXYARdNpl
0ETF7u6fXAq+6fnWAb1Dg68VKC4qfuEJRhlNrQjz+zH+aD7QKkUV6gIOUKG4YpdBRZKV7aKfgCID
bzQuNQFOUmXSQTRtbMMS5cwJxIELWzgOIg7jIS08pAYQlBP2Xdh2NkUGQDWpfQbIegm7cVo0oHAf
OjPR2RW/RAgRSx4P+dy6pxCxg2Xwe3K1Phch3waAxkbhidXeqPfMfduLB3DQ7ASqCQT9Pb/B8QdA
K8IP0GJTlL0D10LApAFgFn+fxW3nAwc9h+78LUJ6OxRIDpUYXlcsRTQcSOZ9zOd2h/NF5e0ZLSfb
L9k2F7KaxQ51A/qAm64etDk4tU404iqZYvdgfAVLKh9K+qKHh4MNV7F5f0OuVo8ej5hoaWmlov7x
sD5VW5J61Jojp+H+NEYrixHS4KPQzdCJPmC/77vxqLP2YV1nWkc71fFLBnQdoe15hXKWzWkz8Io8
zgCGmIt3CwCFWUr/N1ZYnMcxEo6anZWOi/llnRonJ9vZtSxASKuThqWaVIsaeww1EnAU6D6ySQ91
aXScn2KYBxs6b7/xB3VXdcUaP+tzm2/Kw+F84MO5AUSMfcILIZTYTRACO15k0SnR91/NShxIkN13
lmBFxxdsEToKqRV8uuoaa+uCbnETFqBs9QLtYWwZCwEMa/YcXsSWa6Hygpgti5jTcNCo3JvJDGhv
zLZV9IInvbTBHZ6CJc+fi0guhKm1P1KYmSr3a3tC8UC2ZIPJ2JcHubNZ09WeawuIzv1EbJSUvp++
IS7SVyYfY4f394hYbr/v+mmgnwkBpe4fynahdH7Zms/7nQ/tEKQR0DV6JYxi7ioWu8Nk1DW0X5WZ
Mb6vWmpgeMO/fW4KclxuGUhEe+4rDJ1I6l9rTzDUyHYECpAs11lxJKWIZM/h2dmy1GqFIgk9sv/0
bzdtSo5ElVMkT6eSFJihai1Ae5s7uejfH3FZXGAWAOlBGDkjy2e3mmYSguPwrBxGEMjVeHcN28Ke
DbhLfxYLww/VlVgTe3B13SEelpNdOzA13t/zN7X/n/1M4pwmU9bKnNIuXLaFwSxGCAepbJWD43i1
SvT2AM9QsKxYpSf28HRwAbOh1fKpT3F6tq0bWop56O+3krlrUnv8xTjGg/s0crZ+1pw0QRRMV68S
thtGig1yeOKmsq5V+HcOo9M4KJ+1MpHTYm60mq83hdF+iohc+AJF/4Fk66qVQS0Hh6NL3U2Vp5O9
MP1BYTU6NoWEHWMMa5HLW9WvhpT9IUFmNfA+hoV3w+2PtGsjS/RXRDzr4O5EmmCxmrVMk02EaBSA
+6dHoKtasoC+kr20kQJ7E+2E2fEzaTN6WfXbtleLHRaEOxLUWCpY1ToBG5o4jpl6SZLOrL4VGPIs
O/tm6zy1Q++QRIf9JJU/n3CHlq30OXEjTB5hsxjtsw3CJFtMU9VCyLD9tCMefZPmdnhutEPuTDDE
o0OUusyaikfsF8W6LaHWHWhLUfYgEPmYtZ61rADH5wyvWBW2EYLNi5fclSUCKdUM2RcV3AQKNKLq
IV6MC532wDqiIbrXjud6j+fRJ7k0NA6RueH7tuq89lqy0fOtgaK+9Dq9KUMN+fuRtQb2r3f1zZDM
V7nVhXNOrmUfKo01M5slecz6Dq7Pv8j9EBqJIlRq36T23FQr97gBg+fSecWsVRvqoOn6YlX4u+mC
mbK+nmnwo9LArGEZVKAXy6lIqlMz+ToVNv36KFKS5AjS7mAFX2mMSRhhYitUzvyL4mdCJweeGzjT
h+mqEORD8eObs95zy9tkoCtzjlhcptVcp28CR2WejdAq3eFGIRc56jCQtCpt7rk9z9OTMzPiR8Wo
QRSggJP1QR2q6nSzYiH96anqRcw1Ddgo6YJ53X8xIZFS57JzRMFSmXfjful+SucF1vwzYGfPt9jk
CTZRTTbA1BW/JchvPl3bcve9QauAOuzsO7n02IKXo9Z3Fr5FhmTQ86wHsHGDFBFHXU2HexKl8V0t
jaSV49BesaA83NFS0hQDfYAJLcu5mB77RTxsw94QT8lSARryme8EDVxcGb3HfjAbUZwR0SlQjWZX
yBf4kHNv3R0gBynbxHc4L6AVC9xyDHg5xRhHie74c87lP0Z6V036NVpW0pEhfAypUr00l/+d91Hs
0XpCXCa2YvIApXFGc0kecGr25H1iKhPN5bL3CX3AwKz2uAxW5bSKXyPCUQVVDQjMtDB7oTKgW6s0
bgj+Y/mU2kW/AGuQwPtWyhoGGK6yHdngOlZssBEpNbr3WtTZPWcf3NuChj+id211xuEgHO5RKQpM
1e9BDmR8d9xVyL1HUod0rOwBeok805tyrmXbALje6R8ShY16y0AFDV8WamykDjuEFXouMKU4zJY2
DArdczMOuATc2D2dtElK1Hv5zaQ86FQsvkZxsQ4eDVBYvEMXPyWw5JFN3m1EsQfKL352qmluFv+0
QLSLEXKmvpOEoBh21BHCrSoqUr506nb5BpvDKfa2FIQZdFL0l+9nYSmZPngDkFyA4hpSkIKfj2+/
DGH6YvmTkucLUoUDwDQbi6WEbLnAGzK6kIqMqtIdih9l+SQGlBdUrpAtjwUbvx3WU0DFvgmreC83
9HIbCGx7IZjLrWu3HiFhbXJjj3vO4vPbIH2/yheGQriHwMdUFLwVqegZoO/wF9JG/4BTjPzPkRIv
uSpREPEmZbhv7WER8io1a38eQ1lrxZnqWvVkN/+vADX/gOFMcFSVNd0JlUorNoY7RQFRlxHzoSwb
n0d5yuFyhIO1SgSiCNPoDX0Zes3j9GSd0h0t3Em7/CRdMYApVuUGHKxOxaR4H1dK/ISeWDE/Se75
0Q99XnKpcTGjrMMjo/8RKrTtPIQSvZQN120A3oP5/VJ4tNpWQghe36023lFlKJMbqolVvY4VgZ5h
xK8zj4tglPc+clIbBEtBCJsOmELT2FOoCcJ2LBLvaihf83+GxziYZ0dqxsKGM0vrUAs/WsAp8faE
S98drPy2quw5yTQfWYPnwPZlzvKzTrR3X5PY166qY2o61vkU9T4tA161fZUNT9q8Q+Xevbo+CP72
xCnA0NIW3lCEzND9qA3DxuDe+rgif+H3J4A4WBYLC3G7+GDRIDXqdOEQiPcimhvrMzOn27PgUo9s
EqvJ1WkIGa9hLv3Uz8nEnkQeOGS5KgcQydJOGyAKOKcRzNeeOk9bDGBAGcQ4hxSMaqSJDgg4Ljtj
hGDh0vhjxpj7cKG5rIjc6pIqI/2Sr0k/IGa2S6IolPAAqeR0xFmbhCIX/jLUPI6R4qQlwa6Rvoh6
J84TMGcsQSo7KaFKGZhhDSkz9qaVi/jrjy4RPyGMR0IS9fJTjzjt5wgGvA0+NDBGco0cQk3ygFjf
Mwx/nz7hHs5xMKZX5epdZrLHAGGR5N0u0Dxovdz3PfqMH2ZnzzOXm+vFqAt1uQerD8FkeS0Bb9Qk
gw5/mOHGjKfB4kSntKlHY7WOyhnH/Fi32pl1Dkv1Moo0MhbgF183qTCLuc++dDZjNMfOB7cg427j
H+LMGwV6Q7iA28PUrBL8hXn+LNWgaRvusGv6h7M3xHf/E8zYqAGfIHInKS0yo020hRfQf0T+lf9C
etZeLeXQvydNAQlz3tJfBMpAwI+slMf6pHzjXu4/gTRy2m/OAyVdnmXC/21J+pRMoN02MqyTCLRR
b+6ruPr1RECryyhy+1/lzkRQvoVleqWmBSvlP91uW/50btmgS/HJMv/zzFZz33tHyIN89OFcIfj5
YUw5grasUgvfBZJHZaZ9KEQv43Y3OjL+NU1eDfnucQxw7x8gVRTu1vfb1M0z+eIrFqOpaf2bPB72
eiZ1c4gx1b120Je7GNhyVlfLaOBcD+Abuk3dR+HZAihKFdSDpCTwIWCwqYNFi5dyaRNyNstjuvhA
diFIvW2ntuMPXx9uwOdEIkb8pYcTrnRRkOeqrKs2Cx6SwzOcHS7CNwTARjr7jL1jAr/hZFZuITp5
vIhflFjZuSANkUEg5XQTgiSi0q/zUorKU69YFHPDmlSah34/b0YisvLxCWfx7mzNsGrP7DyxhkOO
LNLq4qk/AJh7VEnG2H3P9YC57bsuFnpJJmB6LYnU4cCrXYUgkKX2lRt0MUgr14JTHpFkn1aoIJ+7
kD+jcJAl248IyNDELF2P1EQv5wCik/B4Cwz1EPaAGrmcmFOC+LcqZbV90GuG8RYJStpMtXOhGX5k
fLox3iv1DV4+bE1wtJlA31uha2XuivDSJ/y+UJGHvMyKsfuQ0+AllvenglDLAkpOCq2M5CgUiV1t
TdM7jamygKjA6+q81zRndDX6lxHIrKVvYrNbmGNw6aim+rPofYuu5XXTmhsQ5C0TkNI1BOhxKgp6
ZRljK5FXaS+TF0FOoKJgOPPvIo9x39PQzkvr3/trVIED/kZ1O5m4LZ1BA/eVOuuUd2rCRGwLh3+d
kokVt+t3SZWv7z0JA0+bAeKx3GVvDcZhxkp33yZrPj4+f5l6jm35i8gLTpOYYVgRLYO4nl+M137n
MHUdSbw4It5AQwDs93OulCwBeaV9k0g22hluqvtZaRYriCU/ZrdLm8atNOOQ2HDo42e9VYr39WOj
6wp+HzUIW3ByL3BGempqK8ZAM3ZAGCgAtQQmtwsh43R0VGqVIMKAz6qZ1MPR9ef6eW/jY3/HGyRs
e53vCyL1m8r/e3yTitchh4wVqg74WuoJr/7FNICSeuaI/a9NHi4LkNt7p5DaFtkHeyqjrQH2GdFY
96smU72o4/G/vnXwfL+jQ49vIAOIEaSWMAo5GNav90l01VVAhoIxxyRxKKwrElKWzZrS6A7q7Rex
60kkoO6jXQYYshsH1HnyfUPdA63In6EIV2Le/JoICzjV88kF24d+xSdWcDG5QG+koD/8Bj5NFfgz
shA/hgSiBGRCWHe8nvBg9pSC9ppvN1s+qne49NsoHdEJQC3tzrcCwiQJm9oVUMWqkqRyMv0da5eM
GMPuOqJdm5w2afSqRlelxvaRocfaQHtK2ni67yqJ2cmfvwJt6qRAry2vLBAcJuwQdicsbs758CZj
rCwXVYprOGnCSGgKuVeqM0OlOj7Edf2LcHw3ao3L3J2jIYTZU6Ow4X2u0nINulDRtjMMUsOe6KLR
2JsH8/aXAPMukQv+X9STZrKj+Xr/LMSvpgaOIWexYLWudmbRYbmZac8qsxgHZXFI72pMwvIN5RKt
YdxAqMIGGeh9AtPMY/2Tq6wXTVejGAO3jq/Uc3vi0JQz4ubSGKhIDVXzVwvcCPOSYL40DyURmJZA
h0CmlBP0ZTO+nQsfXyvWSjYAhQT3nho+UHJaG3moiy873lXIdZfOTQlfY3SS6aWekLlJmhtLv/v7
FUHjh5hQM/cN0zBGgPrgIJX0TZSKjI37L9sOVBe9i95j1OrOdNDZaP/pYE9p+9H5efp+sAbnJTvx
H4uXEOBxbe9lksbUyU9LN0cc0glfCfwRIxItKeO8UO0wJ0VciRxbnwn/PvO0iRJp3sZZW5mKBdbc
wdyj2AcegY4QkpIZUqxOWsUm9+pLihSbLbUkdTz3xW8UsrfFmMlu0Z+NUWs7VioQoLN+bLPEoBC9
Wm1TlCaWTEzNMmwnLcjiSyH6U2j6Hk4zZfeV7mDNaOzXPPzE3O5lJwBdCWyMQ+oUVzs72gLaVICh
VXtb3M2vrIcY8kA5kp7cjV0Drd72ZV1KnaAc0c4QPh3X9M7QOtiJoZL7yFIqemSUsi1+gkBg9feB
tRPVeKAZ35miUozMJq2g0YTOo92u21HyjW0/pYpWdiu4VcEXdnObhzUiSFjxEgWeVoLGqQxSkJC6
Pt82eoVHZomO1fV7C47m5lJA+2T9l7eVmnEMThoT5rUojkSUPaCr40QA4fnuHveF5TC07AznKUN1
GrBVhjSNHO/73MgDoRIktFBKwA0QTl55qLAxz4hkp19C4/HfgFOGPbpokldZFsAefY8mKdpELFMP
1dq/Mke14eiO803dnk92VEAl2PXpUtzqVBiZys5fW6z2y5MRvH4888RW9Q2Kgk16us38P76aAyn0
+4RVWMES214gwzOa6INHvlTvIDKH3MsLIDLLcIENCdfqpMHA2y8HPzRh3dDqT7O0cweotq1P5kxg
pwon2QsGx2hNxtYB8l9cwifKAQ3ad8iMjNHj1D9UvHv0wSgcrr6Pb76Biq49HKYUnVgpYU4ww415
p+f2auXAWhhZG6e4RSR83bzg3tU5gp+7vkA6x5EN6aM3WvIeL0OiixUVDI7UxW04X3OD+ftBpY45
VE2RUMSOn7nMTV5Ry2BVTwAO9NdsbNC00piTMDPRhGBpsP9ZqVNNN8JfYRNd8jorTfwaEjJIk9tp
qVr0PK0XSuH7FxSTvBQQ2tFL0hkbV91Wlw498M0og+QErGv4DPdHsq0HMYgHFDgcslvE4gCde891
VvojiVVL4k07kinhuqaOdZ37kAW3Nghqb/8HToJavRQEscV/nNAN1vWHSHXhkhs2RkPQHv3wCq6w
zDdD1z2v9Qlqog4ExZymyff7j+b5B6+nr+r81KonFfxv2xEpbe7IsLjdVsHISNgH/t73aK5eQPKa
FodjsWRJAcwXOZTfGGGw5IS4QzFcY6P3AJfNxzlEHuUol2xzhPfns63D0mcr/SGV5CRqxN5jn6eX
Pqjw+x8s4Li0g2ad0dJAhp1XMKbPxjgdFZkXXPwBKAOYHrFnNNbAi7J2rcVqgbekUl2+JELBp7ed
Fv1qdPpzcm7mEq0yfnXD4Vymhybrgzmx1nYktVXVi87hI8qZYLy7JzDZvpDgLCjIXgzkt8LIAkUG
mbkghlygXg1KxQGJzPSNHASrx2Y3DaVNaXTeKShb/AptAe0HtKWvz3rJxEvQ9ubQGxDwpsf+ZkRe
pwXi586PHL8JZdibQa3DuivU2FrSLJAMpO9qPrxxyChmrpG6M0+SHgvjQ+yieDJhCnIjYnOvwXES
nujozHEHZLONhSLRTCC2VKaLkvGnnVD4/DdtLeBd4vC8yAznBt0ZrBli+UWiDXnQ2tRkTSBLUzfZ
uL5JumoFaSNWInvtHbSBHclEiDQbEmSQjMBkGHcT3YlLAIbRUQuBg2KnlCZ7PD6bzTk1L5WSttLc
Y7LpJaZ0ziLIB4Kr3DXshevSuDSQlkZcvyuAYbI3IseAeGv576Yh8zh5eSD+7jXihfUC0XM/TC3p
QuUhEMwW3oyX8pTKXT63bWmrXnpZQa+h3dxl+57FiyVi0QTBw9AX5SJoq2WanKfppmw9htbc0kOu
G2RClseg
`pragma protect end_protected
