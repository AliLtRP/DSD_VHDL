// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rhru11LnWXf1zvvFrC22VrHFaf6Cyhp+C4fhC9BgEsFawu79ZSHkFzV+Av4Hcz6T
bOkPuNtbhw0WmGScTtiYMoeBGS0KzVUtwgUAYlDL4IUtFRoaoYnyPRuzRAZdgh0F
uOAJ2PV0/VjGDyPWSUb5q//eTIEB4pPw7/DAXvWCuxI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6816)
GlQjCRIgXczHIhi94sxSe9L5GI03tpWLR1hdvup+O8yo7jI9kG4YowCjXMn9Bg4C
JYn628pk9pbJe2EClqxrI+NTOs7IPHvQ4W9w0rVrMeh3cmR+YWrkTn1/Qik+GQ6/
JWyyrp75deAVfkSDZEuYz+9hQZ06RIE0ZjcBSThhlIkfXfajBHMj5A8VBpvDF7K+
hiLljr49Wr89Fqj98Odnjrav8O6A0tBlUEasVdy19dPw0FtyuadVPC6j8DyvV3kc
sTXfn8g66YNeptvE2WzQSz4eMyBwMEOOV1hqDJ8YK0ZfEIo7BtBSGlW4YZ4v5PQW
8BpYQ02iMAJ23q5UdAEaVMJvmRz3eoYaAfp+xuLPLG0vQ5/+aAA7Iwe7rkEVzgo6
FzHNwCq77jMmcJo7bJWkQz20/fQQ2RM7iu4w7Qvez2DmSBxbHv0c03u0JZeDQFF5
FjqQ1Ckos0GhBbkjtcwJljBJMhI/ARoOFh86jjT9uE5LR8WvzQ8G/yCK5vgGGboi
ODAv/FbgweTttZ2XNt7LXohzZkeBLOWtvmKBQ0F3Yd6UqxT3t+pD1/Sq7qDOfVLP
mMAFd9PVW58HRCfiotghNqAoGcTGzoq44A7DJPlVC6gS+G8iiRPrlzCUQqfCzcf5
VZF7PQcKwwAuv1NrbeMRUrKBoDfRJNf3rkmTV+hYk3Uw7EhqlH4V3b1ix500+7Ud
k6yVne5RRhkIxfqxqazzco39xEyyHU+tkse5ly+V0J31i+9rhfbeSPnSb59cGQfj
4wdjtj8Bpsu7WaTAXvthaUpOUVpC9dfjPNcW5Uo5WPItS42vR8/6zNV538Efqklw
llciza8Odu9vZJSxpHHg/ZO8u+LnhG7vKamBis5bQEYldxRqTUSB+csTXUk9C/uZ
UOCjZkrR0TIuufu+Mpysf93HVcCDRkm089b1VmiBRJoqjB5P64NdAfivaGU7P2Qe
eced+U3fB1QQi9j9L5ch8Ml4X45ecmkgqi57EeW5jYwKOBVhoyvDf2qAmRkjk0rs
HtqlFbAs46AlBOzvZ4Vqm02KTimRj1DjTU95RsQ0ekWDYOr4f9s2hPCL2fxAFiQY
FwrZACs5aQ1d/wX2BFbMg5YRzNFuvLQmZtGBqLOLtIjgZiAsURGEsD3O9oCV2dSA
XekUqOtVVNZ9ePTzR/avuz6ZiGHkV5tJ9f4eL4X0deTMJocUkCro0O36yLgTfJF5
dUvqhhRmb8+4ecLHwqYFYCQvOqVF6JCzh2N1x+l+97T2QBiDb5ye0jbeo4G1RHB/
Vpos0rj3KiqrjthdnutaqWgXZCmdlPjYV9vftJHVa1SoptaK/AtFIUybt9kDw62W
nOSUKYdVv0hDi/iboprcV0esttn6D0MW3K5NQC0LciomRBw98ddb4QXPEc/+6SI3
/plyLONat6ft7kVfh/v4LgETkolROC8CKImomm9/abZYoZE1qQZSL5qeHaSjBHjy
GjMd8cm6zWVakQutzkTlNWk1VIU7r5ZmOcE+J5KPrEYpMHIF2Z8PG+aErmsG0Ebv
Z2eI+WJo34SAYv9Vbb6FTdTOVhdHKRTFC7ghx/MXT8rlkR8gTfNwB0OnHFSS6s76
cW2RC20Z5fWxxZbDv7xl47UszUdzv5fjGB6pWl47zxNoxXg8E5aXaQSEWNVIcz89
rn2N63MiNit2THBYuWcxYW0yIKiaI3dmgkO0yeKWMbJm6H8zQ0Xue4/z4X6r0fOC
z3N7RYndOVvt85LmsL3F8fidq9eNbI/mU5YJHqF4jGqzm+jLQoXK1cN9ityLfT6L
71u2uTwDp8J5ef3mKVoGdeY295oK1p7sRbyck1//q8fuqvgB+5XENxCLD/fSqmss
eSxSin7iG8oMM/f/23YNuf1S6sVntZDDrmaeYma/r0458hpWjt/VIr7r0ymxc8xo
nG+z1BsDaPXCsN5tjrOyKArsoVCckIV3QdAqYYFLfhUbn+nWIO4SD6W3WFyXWPoJ
0+BkKONro+ZSoWB8kRza02/msQkhWPvoeY5TxL/w9LKBHtBsC471JBciy1uznspQ
YtIJHJA/BHvObeLMCIr5xFhPOAAQueHqjD9UgKjWhEFr+0nssECVggpWMT6nQ130
+SJAqOySGPTQAaNaphsabTPb/huLXEhpt5GxcWTMWQYjCYbuYeqZSyqGusq+68ly
mhXp0mY6nP5rRlV2MfIum8xAdBtMdZVHKjwWikYr8DLclx5wCg0RsqTzDzJgpRuE
h4H7a+unW5a0EXs6OdifuiMVRHVfkMub++KvCXOuCufnvb9cBIKPSU9oukyomH4T
KcfRe3kRWfJtSeDL2/37YCS3U7boTEfabzO3xf47iBCSPhy5ViBSERLsSLsOt7Dz
vQ8I4Vo4Hb0/z1tdurks8xoOFmnLv5qdlPXuQrVi9Sm1y8Qn+hT3jcv6k2FKACAi
IbQimmSMvirmum5jc1HwbUmkmZEjG/tTBf1HjwD8uct41T0UEk5Es/dxbmg1tRJC
bljK9NIXHQn/j2brEJYqgvujhvZnEvZUTNokG6HqAhwuwSUF8ngljM4raNc74ejw
Uz5g664dCYq6L3PFUKmt20xNrvVlrkhtqB9BDTORaProHGZejzEBLfuOPNMEnJ+a
fCy7K/MEl4oqVb192nWqYkilNsJcvwL+ao7BQLKKYkp0Dv0Hux4gANp2GIcmF8Fc
cXsz67CyMzeZ8i/qnKqdomUOGL+tt4vZ52nYLstdP0fz+FuZDuULm5wLlYKC5eTM
i+MN1vLPRLo/Do+KzKSCtiDG6M7Agoq0+kL9x6cOPaUaflWE8b0kYAzIk06GKuwY
CvX/S/t5i+nlhUbP779/j1qfb190eO2VVnvXiG8c7S3MkCkXHpdFGDx42K10O8LC
NnCDmB/tZAf/KctQppmVQFuxoZUViur7w5gCVgLFBPS2EYuf8XTmDAKwRUVEVOU0
x5cRnQVVNv42TPOxyd4L5cpPWU3u6vxLiyFMOpO54PgaSipkNBG75v1iFRA6uD4+
Qg62iP6y1aS56rWkOFSl/8mvF5LVQiJIyPSrZBomN+yjYU3pCTCdTjLtrfXO9A9N
6mYYAO0W+vI44w+fxX+yc7Z8itO9tzjQygiqEf+rQztnVOBFVGeWR/fFujn3pp/b
bheuTRYQiXuUk+uIRM4UVOZWl540yPJrmxGL/+GNdL++DdVTGYXiZpCLqLtyprHM
NZxYjWKuOOHT8UDRBwN5FURIFlDfCD6Ea5v1iri/xz68P6SWVfURcmO1pObfZIcC
9Ok32VVEzuh3mjtN8TuTprXHhmim8SSB5f6HcbIQIk8YQ0A7KAVVvbB3BW5/SzA5
ScMIYhJEs78dTnkVlKwm0yjfDb07FfOQLDoaqDhVDnM4hau9epthx9Neqv1DQrFY
RyUhdIdfNceiBU4lFABQvlD9Gk//FNvBWaS9LCYeKBtaOm/YM/mr7ySCfGadl8/+
hqRRxINOmsCnKEgekofxVQHlP4RAhzQ2TY6UpBYq4awEGEXxYLcDcN7oihUxkYG5
Y7bLchST0Dg7ajJZqKnY+IzoBZOQ5pxzYiQnrKNsYZXk2Ek4JxYucyI3Bt4ZC+m6
fViOCmRV4tWCXy1o43Ib0179GaxOuxp7au1ySMJMiZ654KBUvQd7Jcws0mDHIW9R
rSIlLNixejde2UrFVhsyuXJxDts1ktP3VAvF1Znec6Ycs9boMO3R9gcvEf75acgL
eIf4fcCd1Oq2iBZxrdo8jNPhJ4pifU5gEnjq84v2//p1Gu35JTd7TlPuOhjhYE7P
10yBZCBG78s34k0bkK1vItk9lrPXWlECIMtIU9LsZH1929QAvfpDn3groQ9QMz01
0YSQ3jSODFEx+884PbxLRUtYdfQo5v0k1o5Ucf/uDRCWxGbLKBSaht4CGWLVn0sT
HY6NTwFqVa1UwBMUihI8CguUAsRPWFMpneVTD4/+1GmUP1nMrLumqynKb5j1qb1E
6+PUS3pLo8kGuJ4kJxKvld8QAF7nwmelB4x0DzOQK3u25YizIWvvJkofKQOlL7Y6
KxwR2rujIClDysu393RZlNIaf7mvTlfDw3Jl38FKdaynVZ+YLIvLNbUv0Ph04yN1
3slakB4run01T79vcnZ/e8muGNZs5qGUma4eKC+4IUAjxb9uANxZIjKX/sHmYSv7
pZkmpeo7fLV7hOoejdE1pY6sKeOZtrkyiKd6sS0dUnkKAvY30m256AvLW6D5VUMw
Hvh28g7F+TA6qKC7i+ykjV91TwIl3jgTKPxz14WBpzKdrRB6Xpw6XCw6wssX2G61
HXOcbj5AwUx5Huufb6aO7MYOMMl4duciSGyl1z3E6tlXShMn9ipnc5+H65vu+wIe
8jJDNERmHctkVTSOokv9R9XXGw1tBSVczR8+sdsoeHAozNvlI0oj10Kp9rHlYyvU
r7sbR/hOk3D4gXWwEmapW9LI6nukpDs3PDd0XnsFyk41ZXPHlzNxX5OFokGvAgH4
vmxnLHVRxfjOkIe/plJ1A04VDBwcHVFJuy74+Du4H2LSvXohTs+RvAOdF8RP22+v
klyj1sNt7kSDRjXN+JY/8dm8F6/tscazf5RjejTMSVXj+x9NdPS9QND6cFXSky5q
o7Hgmym+iY2hcls8Z5aKjYgOXj3cg1K2fwSCpIDIXWN4ePTWCwKLfssTxY3N+r/N
BgBdXgHxvHzqmgbRUXjgNKvsOA2J2vMm2VpL2vk21HAW0PGmkFicvp+kwgvRD3MI
gVtn5ZW/D+HyVag1kd4glTCVrmQNkbqK5PTsApd2LCcwJJqxcX2hKSbxfp4HN3Yw
QPheXM8anCGOIk6aojUNbArl71xsbmByNdNLI0Vjahb08lMZhmHLySQcs+LaN4jk
T5IjqjJWzzJE/vsSQKXmbkvrfP3qNyGJw57Oy5c2dQ33aJAM+O9iOgWQQir/Y7Q0
rHtTyrQWcwxb28AvBT8DDdIIIYOmes5pmtqZawab11M8UK1CYnDNqCU+LKrrxLij
SoJniHMCkWThljPHsHj7TMMyRiT0UIWqgiLx2jKEdt445xcdHDA/IIt564Or/8ja
zoQ1psVZCDKfpUiaAoE0p7HDicO4NUkKjn4n9JUZGE10djV6bauDmY6XyqEtusol
XcjQSIQU+9EgxG9y78IMo8+DgY0BxcJHh2k/8x0oo9o2ymWRYDmZFSib1lVoSV4j
W2qdFoRUIVARx6vVYQtZ2j2kfukmP9P9fBCMq3IWjG7WWccaOLzZEx/nQTmkmZxd
ZXTCBfUEfQc4bh60bujvzjhgVEKAX8SR8tdQw2bELwzw5GqDXPx4EXmQwcP7NG6L
FCdPwxYHpIGvjeVDaTZkB+zkDfrTfzbs606uE1j2AcU796EWkwsfXArzfOhWK3nL
MPEMwdjLo/2HXNl/NNnNIJTed78hy/QXqHMprM69FSExFRM20wYAn+88FBLP8uvC
LYWrNxskrhjrgtmWQIA24hJLu5iyimRuqbiTNARWkT5cXo3KUWGSduu7XhVTDVkp
el+rdpsV6tviJvfJDubKWH3vdG5VsnIt6SVEuC8A5XzEkhVQvkXCiKpe8CxXYxzc
ugZM2Yp9aOFHqCTcUVrmReOsUF+TknjBzLeaRipxGW/bw0oXhdl+cN457PJm7GKT
Ufr5Nr+Vu3LZTnei1oK5xvkQ7l/bGW1rFMTArKZ/+0KajegkvsygJ4GGuoc/pGbC
aaOnNZfs4OLVMV2BWI4/7f1xHzL7GdjP1NkNqK2mvyYQELqYBkAK5KNVrmu7+B5/
2fSy9KndBZ7q3KLYG2vLObIP1Zw9WApe8jiQPr4Wqooh+uClUQ0sExuklWe1guWu
joTyjHvQmcEXgNy5snUn60TWU/tEr8Hqde5oLuo8hn8xwhV5+m5S4NeP86Zrx/ZQ
L6k1ucN92PvkXjM8FEacRnlMI0aCUvv9Z774/uIS1WXw0Irw2WIsuzHfE9Xq1He8
p9DKBgyH+2VPg4dMGB8o56lB89s15mosWxXd7IzK1t7c9oMItu+3rGbJvHquUbkd
afJopldl0ig7xBugNmjsxfB5QSTEXne8fFct4pSiOLQaEJKQxkz7iLuMucvHGHlL
TgVSeWh280QetETF8VAqKP+w9pLReOSeuMrvi88dv4gQ1JeZA9QwxAwJnMuETIsk
5ARF1byssMqxYmTTuF2thg8Mr+ord1RJVFDG9vBf3ehjIlgBSpmVUmxrpQGDMXQO
QIsjxJrpffNlSlWkOSpBygfbXln7E8ijjKDqR8H+JeyLcFF/rdogOuP98JnRDPfe
7gXB0HpME192y4MkL1hC4xSLZsHtRjYuIYmHLRUmsGGKdOnC3/Lzamv0JwvfICAR
8on+LU4SnleH4RqzJzuJ72DNeSCEURfvJPigC1643f9hNjmEUv+CupFKNEqXB6c0
c0IIlt/8TFNtyqMM1xf45V5ThwdyOHxhJpwiiFtrpmF38zGZ+csmRN62XAJjlzLQ
wXHOSl2+WmD5dDOHv9HfrNumIswZIosuFLCWsa8PVZT5nJ6wGgbMFdtReJ9GVHLm
EH2fao0IKYunK3beZ8mPmqofquyNxRlH19Gqu1mN6AB2SR6BKmtGsuSmK2pSMYmX
PngmTnD5oFatqAkcDW3KqUF+wQWOk4IRASiIgk8Ja3NnzZH0X/tHH3Da+Y0towh/
tBvRTu0+GEQWUoLtR+9SFvo3TBpEkILjqmfwrdfcGVdMlwioAPQKUnzT6ye5Ewk6
gmim/C5Nr9zFlgfd2bGiqPmGlBCTUxEHygoY8QgcjAqTnZhLjXks7DhSQVw26hj0
Gxi0JmLQelE+yvmFLcUl3LTPIlBZCdQPWE/Syoo8F51+SnmDSD/9n9ZDSwAsIQHw
Qs9830yS/7koukCE1V3CWmHaXDdrkuxCC4E+p6RNXFIXx10H6RJbKrnm3+PVhr4y
emUZhjnvGMqGluQJbaInzJl0dFux1uFBraJ0w+tBsR6ntHzJ+CEznNbIFtqG2afR
x/d2uDHvgXXbf2JJKyf+DqsRLbeaApTkakGOYFw5BfjNm7YFFaRhDMCY57VNZWUO
ZJeFB/OmJYBNFo18Eq17fTggf1fkgltfudRCqVIBONRuP9Gt/X05dQ1tNy4ilD0y
/JnEM21Li1sYiFj+BhBN2W2l7YgmS+cy5vTUSdc9zYPyU1IjlivRzCxcC8xupSzC
j83uPpuJR/+oDXW/ZCuFDx3+YrrGLm/yAUi5OefWQtxS24QrpTodzT0qQX8WSpgU
fidfMvbUGSgBXHnf9G561gwOJNcqTd8I6oCzQjTxEknNyMvPSyVYuZhSRgPsfx/v
AANZL6Itk2DiRaD9XybT3Ocf8p5AHZxcdSHM9aFe2Hg5ucvz8DEMD7Pj4gdpqaEO
ZpRi3CyrZ5nRlcsxMlrZ6ijUEeoG0RSfjSNyQ9q848Yy0huNeatwVA5/cql5T0/G
12AVJZKDO7tEv3RSgleJPQVICNxb3mzlnLOfB05jBBXNmHpjEgalUllryYAAOYEf
ojwMFlxRtUpiQfUTne1urWpgWGk+T5FIxgU+0mvIi192HqQ5udMh4N1LPctObVeO
mQEjig/kqm9H/xp14kOSs5gqneTbyikjTni51iFS0YItMuix77bK06zmoWey70JG
Bchc9DrQGhpPdP6OmYV7Bd3KKAdcCfiBGMfvfC4H60RLY1AubLomkYiE1hoO0VLt
OIrjbouBXL5M+tkUBDfd7iGjbvrW89xcYfhfFMeHenYxTUBif0u6t6js0UqdK93H
QFxPygq+5jcm+GZTzZqA1Pw5Np5eFhyTm4k0ldN/oPryQrshwP9VM2xqCWS16/Va
hsAnUulJfjpzd8sUUperXtDpu6ZhkrTNDAGhDP0397GF2DiSI3EP7J37zrYlQGPi
C2F44usgMXwgVIOX7y7avME+m3sFRgpfTwxVHkezZ1NiFXnFbGJ2UlNpkYpW3gUz
wSHHsOvE2Yf2DMAnUHSYQ1atTUm0e9E7pSjWNIsd+7wMrfLbOL914Q9tjdtr65q+
nAb8BvcFRXF9NjGnJj8feS1uDguD/xijui/d9q7oceT2jXartP4D0DbYcYuDon1s
aLGUK0MxSg5dLLY+Cd2pjOk31NbQZUmHM5P1tI5UWghR/FS6n6NRQUHBq5MsvtC1
+zK1NH/PBmcsQksEgQGu9hnrfE04WZLQTIv8UOBrGMX9GwWS5lmQ/NAN+ruvmJ5P
90aOaMIKU42rgewqju+0l7+kqdCZjvx+f6qzqGWG96faa87xMxUGGA9+To5q52sc
qflCnbdDKLVHtYtBoTJaotafGvmiPFeu7ORLba5RBPnGBfzcrtkkuODVXgIpD26x
ZoMnr32aQ2+7Cf/hUfbsmE8S26zk8A6iLeaMQyRVIlxn0s58qTglo+PwDmtMHMu/
d39UuZQxdL+DaM7OWdulFs25Qxz85PKd4JiTrNRPyw8MLhCivvzFMGfpTwp5iD4g
6qdjxGDZpdpVU00MYwZPzLQs0cQp1Z2kh6nDBal3/4B7IAofpEBO/EDzChSnaf9a
67fydsNIfaQAaX1ICpQevhSt06c9aiIQghtRmRgFkZiaNb0fDU62zaNC9oNZJqsh
rRKADgPw8BGv1aTi/4iFGaPwM1RX85UZytN01MDvpKAj2GASX78rnm7zKowpPmBt
CURIN8k6xHr1FQDuu2Z8AlXV7epDDKicV7NoB99UZSAn9co46826gB+C6Fyilv61
+wNLIbMgFMQpPZvB/G9saIV0QYsUsvipTqUExPWpgoR2NhYgiQA6LJEhGVKsr77b
AiJ/VmShPWxGxHeaCzLrZEi95j9K0etFbwDgjeklMn/IFvotmkDC30SxuwcwmmOv
LKccpI5itIlxMYOH20x3iG/PqbCKgD1BdJyJLxO9TKyLfXNjqSzbtU7+chOJnyNu
hV7gsXhBbxBCRY5pGH/9mxo3HHFfl2kStTue4/deSSZK35CbDqoC/8vdLNfs+dDG
Vx9Fj0zMSJmAq3i5/TN3Hqk7gt0IKVtSV4EisCGKZpLEBl34hwtPFmSJM1zx1ORy
VOz61n96ii/3xMmih27Qg7Ypy7R191STPCiQpKHA+fR3yddlVxr1xozW0SMT2Kuz
`pragma protect end_protected
