// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
AN7HsNQ5mHIgd3Z/q+ZXMAaAjez1wiojoc11REtqxQhOg2mFUFsqdScoYAFSVG1mvWk9IIME+fiT
P5Vr0dB2Qyzo4woCrDgLJtdKyAm+7NK+MYmh3kHxyYCEC9gwLIxoMVIF9uY1EEg8tDy+zdGpnjaX
91L96RAKelo0IV/PTFvkHsdlDHd9gat5G6O7551i8OJ3aa11B+gXo64KTkj5T+URWL8yaUMh1g/q
qMkBlsaliljjeyOz7WNKQPSIiFYwaQgXZXw7lFVF1iZggIisS1G2aKAHEB66gjJUsBN7apd5F1ho
oq+kp9LXURqnkoyW045udtK7zfRhcb6BwzzrQQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
p78kaBOKpaXKR+SxkHV3f3/6FiGr8NsnHdtOZlHO8rLNac/Qd4/XvdA+yD/b2RkGrXCyO0kFvvFy
zfpdtcI+EochXkQ8J3wYM1x6q1Yx+Nkg4ZGwZ6O5b3UJybRkqU0TeOB/7emkwvrWwQSzNEtIp71v
GXuXMduJBm3NK6odQwCCWYANf1m4vQ1N9/2ocH2SWQMvbxOOyR9gDQ32wLKCYHYbBjTysNYEeaM5
220uv9HagyRiXdYpSOkD6mKIOdlolSE13IQ8zNP79w1BsJWfjkrcXsDrma30zCY0FLyn1Vth7U3x
7AMrD1F+p9wPXisQMkV9uqJDwGqhFfn9bxUTiXluLosIADi9HHRCpemXEATPeapi7JzteYRVN5g5
b/XBJ8lsFaKcwg8Pbj+Mi+sbmMfhUzaXV3+gg6h9Qk7gNc8+ddTTdg6Sf1xIXe1cv4wAkFC6wR6b
fVyPW53RW+xNkLeeGgPX3/ipmt/BgWhXB94PFNU7pNjSH+iCAjPCP/WVm+66ujBXcEB8Y3hU1SkR
dxTGqhLy7nnupcaPEbsKn+6FkFb5ZTEhVmVx3K7nm0yUdAl3dOurvi9ZFCwm7njCOaRglwzEVKEN
tvFiX+eoSksJiZ8yoK7tEWL/SytdyRZGPMFFgUJ0E/54SPrEE8xoQMrOrJXGCmxcE16lgUrGg4JC
6cGHvDpne+b7bXeQUiXrBY78QmhE3msfvAl3rQo+Mx601T98v0mJ3x6Ut2H+1TExGHHAaWdWOO+8
czD/uqPCM1QHhjGvL++6qNZs/VZnznnUTeizxXK6j4wHIBFwjvzSUQfoG84Vy14hWsdoAg8D5fTK
YDy3uqXrvVY3M8HeEYGyjSvwdgspwNld7barIdINkpKWTrEFQIi1rOoE/4W96lNPsbp3xhK1ejUN
j55iS5X4IOXYparibPIUSJxvR+5yq0IwqjSTvSShjByUK7vFVSKvb6RfUNC+EwQI6DKBCh0xDbjN
ODcMhRCwRUjCqWrDq8VmL+qF2kWuXpGYb8J0ognTfdsS409J1YCc9eAqQBxUxK2MMtn0FbV7i9f0
oHeVQEsyr3FqK/O0NQLhfuI+2uCtwIJ4OraPb2jT9GNwMzxGUMYV1LsEdJjuIOsLqjYN8GocW2UL
Jz+3FW4y1G1JerL54T6muCTIGwE+wyoD30ecImoVVH361d9qxVzB9PExc9tbDwqY6vli/ikmSJJv
vTGmyvUchcp45FX/n7cMCuPXNRJ+P07PYZriNQx82m5Z7/KhbD7kUwBv423IBGb2VJwSLjKCOFlf
gxwV3S7hPHyRte8nO01kKgqCHJ0Plvb+4coBSJmfPjlWGtZ7nqpC5ss4o/pnmf+dG8CtKtlESpeb
/cx/6sizsSF7GyxzOPljJO7T/EcS6r6V1yNkeiIbnixFFL8mmtN90t2t0KQZKHdnMkU386FeW169
/VQgdB5ucjO7bbnCs6nOPLaC6vgK1CLp3s6v6nKBnxyAIZ6wkcGp9B/5eCkGC5EqlRBB7bJI5DLW
OYoR04oCH20QOmcGw6Mv9mlcb/u+eAC51FAp+vYxzlZVTZsAxpjmWuu7ZTFmrKrVksHRndfBMVek
sO1Bk/anV9NtoNjIr2ZCeY8rSfq89JBo736Q5OY//m2Lr3DqIXnLb/iwgQm+3jZ9+ICE039skB3K
lkWSyJmlz6BZOQNYcHnmjclPCVoAOaD/md/IZVIZvT+mlaQlHWHCXqOBu8FoeFzO5gyh08soF+b5
WnFUkFGiuyfbfvrh7/UlqUXBsGGrbptxWOOnVXz6IvsU1z68s/zdfmURt4FjcDoTAP7O/QN8Ac2U
2sChqm2BFEsB/NA5VZjLJzZl5UXGSnXGjHNJdsJtDIkYXqzUCsaEQ1FmdtWHe3qYnn3w+8kBPmtv
xE+PpR3HKDwAKPbf3WwpJViF25kARPPXWPPczKJ+hiPbmoQeCw0JdOBI4/6Jbb5DLVTqQSHIRftU
TkveAe9UM+aye+Lwy0QDqGwt7sbopt4Rm34DeaA0Jgb/9w6GemhA63nMKWcnYVXhHp9Q6FSjY4WX
ke3uOM5JaN+d24Ubbhn8fxsy3oI/gKiH0e+XwRRBeidOUQ8ceewY/IERJ8HC17z8m6XqA1Ehhm2M
qD5aKF3PFkR5uImllI0PsPwylj4R3O0UPOHl6dpbgNYb4TXN2SxJjS/Q1TPqbTX3CBNW3HnsMIOm
/fgH9TWDKRnkS0Bay1K7pnBo4YDUxZ7EindzMnenu1o73p9djEosscBX+MYMOz0k/9GuwAerlLkr
n6pSo0cJWD4G+NxafrhvihZlHkEKz3+BkmWFeeNknzlAfzgV58P3uMqjEPQ2yZ1CphDnO1ryRF9F
oL/m0ksvPNW/njUvGDWlv/Wh+TGDgsIsS6q2HS3QLVM+jNniVB7wisX6iqpfX5LZRT/kEfV4bCey
eY7W07n+7qyKC6bKcCVnOjplSj6xaSPnXQICQoT3BworOLdiqjGFF8fqZhXF/pzr25Z6EVhMZyqI
wA3hNfQJWmoplqXEhmPywl/21MyCsrA/W2cJtGRc85PczaboeRMI24XyX+Wwri088fcjkipWQzag
HfOi6Q8oyQtOE65u3SVWN68oKk4VKvoUEepFvPf6AQ/zxGjokJMRwWXGUD8dKSSOFzm3zhYwfp++
3iYz5sSqJlnFEsM6vaciAdVNuZRI8MN18y1skVtmXl99M8thN3sj7rYq3ld3c7ZSSPUkErJNO11l
M/4YwZgqA3aINcyOniT2fTZ0pTkqg8MWviwMoCq7FtR7uVyWlruvug1iK6rj0B2ILOeSmyDiObLz
RB+EfgG5N57jn1MNQdCB5LWDUMDHbf66b4eXq6GerRW4BSLEZl2EGpo5jXrfNQqQ4BeLchtfFNLg
G+e7EO8hXw5e0l9gXJy15NMqO8Bhc7TF21AGOewz4EamtKBJIHUrD3VGv41TkYzYejAk3hoq/9lS
5NlhchkLF1YCcYyN2HnwS0h74lUZu62fYL7VP4VXmCW/4liCixq2OAFfLFeeuGJOF/ObhQ81oCUR
4vPvfqMwVWEc4VPGPRAU95t1vV1Fbsh53z+zdvTIFxHKeWXM3/0xMsFtnaCyIYEHfVGXC2VP64Tl
y6/4/2qz/0wipZWH4GYjUSJwuSFFk8bezL7+ZsHTs8w+/zkg9WKEpbremxZPoaqFLZf66PMirVhh
8/mQEkAmL9m+YLouYVY8DbyK5OWzxK1xqugAsBKmQIjG3VFU3+R/K5TAyhasRvlknfTE8O9W7V6y
KkRhf1I+3VxwYCvhNxaY5yrPKXjIh3GXt0ZSJcQ7UuCG+L9k4rzqH77npTzVhEwsXQfPl655xFwk
jSFy8qUDXnNxe3n8KZa7pMTqGNUdRDLmTDN/cyZAqWwi5f9UvZzgwlFcRxHDhFdn54ejX28cBSM5
7dXe0fO3xZf0advboxzqMWn9fl8yvZ7CNsIX/4T3enSi1heOO3X/LpfMD9mVgJfE6GlovrEIl8s5
yAsQMQsmpqYwd5heWSGY3DcNKqYS2ILuPFTUurDtp1FxhePvKw853pBii8eeKzIXVxzw/dPXmtsJ
8SCAFXXeA8VHAF4elZGoj9GlZ+xupUyLwa+FOe6ZYp2uNEIC2RmbfBbKQZASKWfK0tbzg+DtInmG
jVe9JBr2nQT9Aal3vcpje0GAg0Pt0gUbN467k7z4PCDIkxWK9pLf6UfROaOEEUS/HHjArHzmY+xt
baorJYMG2+o6HR2mTsLMsmnZxSa2mKIkX14QdwWNFJx4rsd8CeuN8F/RNserKS8RFrSGUuYUmYJU
Uy2Gq6uNausf28JorCkzq/VOtdgnGadHAdY2UiMPysiuldtzYt1NfYBBR7vxnc3zyLL6zl6zDmHt
adAdN+ZNdLWlqos+Q2xYbo/PcfQwHs40DwzooSY2ew+7fO3L1THjZezZLnzI5vEpPvL41ybS1Fiq
61Asb1laXeIDsAheJAA4yqb/ZsVlCQOiAUTABzzqUJFy6LNZMowIrdBvqnlUhwUNNaDHGBULX3/9
fgLUvDaSEjMdXutQOrIOV7DC427CNGNpCRpxJ+28B+LtfCs5x382Hb067vb4jA8pnReUtHv3P3Sq
nofWyEwQ8YpfjrDCDAMFcaAHnkRyoegjO7XcLMq6pfp+physydQ7kpDCxa6Wg2KUNUhi+3Q5N98w
i6gMekmQNZ7YSqbuifhvxSKPnaDzYTCsz3/MTW/HVofIHuKORdNHr0h7Xvs+7I/ZbFRH80Zdl9DA
/o09OsYJlCebDAYsMtmlk8tglr3IoBbhSmHnmUEEF76/mYeiWJuHcnbw18sCaMEwJolBoJAxtBez
4BEJZ69HO9fafiV0azb9CCSpq31SUJzvuCef2iDHhtScLP9/JEclBVLodLcbzJdbx6bInCqxf9vC
i1HKvifSib8H2mvS/vfEmcKWh04fXXnhZZ5u6kdAg+Hfu/ZjJLbK/7tzXJSOMqZuYXMEoj0s9+En
BErwtBelbwzzmiXhqAHiE3XHmW8wVly7owVcGUyQR9koK1pGU2joYzcHbzf1ZEiU0W5XekFx0S/7
aMMxOiP5uDnnD7vaFDKXtyKEkzBmOdb/qvmIM2o5jjLKsTKEPned+yJwA/6ePkjgmJMuOOUFyJaz
bxkvenPbAjM4A34lyzPlQAe0kgRLvr89fm4i2UhTCc1hW8z977sXXidZ3VYR6uG0wcOPjZqWwgWz
+TJMZw0dGVMOVNE8MiSaN+QIX9233XepLSNf85JzUwbwXYJv54FgZ9PXiWnaunn1v6uVyyiDRLAZ
/gzbNIY2sQcqnVT2LFsuRu0Tw+ht/kt1qPN9NDPWXqGE/zErLvZUsZgkCNADXqzgwAKjXvmy9UZn
7RasGSOaIu2HkzQ4W4ZaN4VYoluD06sWjSKzNbluFv+FMwOTVrngN8+gFPXDxxcnyrB5jaQDndmz
y8NXM3rJexIGRv8plHSdr+62qlsxvQSPQwsBYJmBJC9nduurfueyN7PovXFDCOZbKbWTncTntEwX
zsdZa2YpTbolGhCzIqAkYtQ9Mp4dEfiZ+QxzJ6NwPHcivCQdedJbHdEeOPLJ82UWZjEXQxVqgCc7
3YHp1579mw+N5SgHaQiXfri9hNL79MK36YXYDqsLV5+UDKg83fYIO0zxTtUpwvUBpbm8BoSVlCD9
O2MHaUxVAJAzv/fhVS0o7RHOmQIPn5xWkhZ8xeGzEdn2H36tEk7c86NHEwOzv0BtoP8FVCer38XH
Fe3jIk6hjDKSe5HRIRL6tznoxqTaoqlb4Vs8fnouS/ZXwmfJgQnjRfOT8ylLZHaU1SMH+djZpP6M
nHv7trpKALE8jBjm0a6xx/ghkct08ozPIaHXtNHlHXjIQMeUxhSAXnYltB6gU9Cfz3m3d1jGktyF
pLmpAqD7u2MnlOHgyAYO37G8OU6G+BntXqiJenYJusQQky87uPCOgm/vb5bvNFFJJuc1cFFuDdvV
B3V4NQWzPmNn3oetvLHv8din+osPM9LqOCCkP8jfpoywkNF+cX+Ja6EGzO2ep42CwPf7YyUfYeLY
Btr7i42COiTz6RUSeRlJKgcFM5q0JogHVnsOmmNPHKA6PzDGII6fNwFUSC6fxhtK3ZdvNyEZeL7h
wOCjse+aKN49KANxblpi1IXj7klzPcLeBdzlkVOoQXfqGf5WS6C0vQRky42bMggwj2WMtZSCoH49
Ce64ty6m5A/QgVdhP+iDnB3fLEUVR25+Mh585Gu927xuKPfOuX3fZIlhq4Ca0OookQiy6gkU+Pe9
xRB5MnsAVpAlvSERi6ciILvf2ZdP/rvLGL1Dc3mN/BCCm4HpUPo5pHRBnyaBeru44TOl5yWybgcK
qV8CRpRbucYqrSnC9DPvGMZMbMoWPUOUdxNC3oSTL8+RNgVxUB8rIUYOgmwR3pvDjfCDzWFC3v3+
S+yVl37bp+L8dT8bZt10U9FevUamJqOEl5O1/tH5EX/Qn49WoYb9Yl+iiwzny6tjTp7BgoLt/FKg
ryMvkgpwp8A10CStssSHrkDxM5l2KVUBaySoQUlD9aYtTkLdYXvo2wdbqQVioOWRb6uPHZ+dSEVA
JDmDhI7nU/aFtGmLxALk3NJp2tX2iQFn7ztXHx1YGp+bJ3JCuqtrL74lFfZJEdfBz/2taoc+gnan
+to8vZa1dYtHwYdSvqfVe96Mmstwk0gCfTUBMAQvZU5UFaKOlDz+C/MKb+ORGWJGnKTnIsG5AxwC
mRXlwndp22rq2f1WVi2q3keMq5QweVocT/dcsQIS2R7ijJCAwyxtC3yn41ybP529zJ7Q7Y2eie9+
K2+DiV/RezUVfpwFgGB1ezGePh3U2WZrr93FBOTR0NKpfvnGV5pY8+oiS5BFsEEyiLlVmw1RsTna
hZeGN6sPH1ZPcUZ347k0dHACx2u5KOmVLpGCILIEN7jt/7ib+Y9iRsAMiZ2e+HCzuQRzAzxhzL0c
9WndrKlvHFq7rlvyybG7ii+L8WbjVCjLvOGEheA+a9FcuCbZCGEpJgPHonmIsEPXr8ZbyRpvzaQv
Sw8nmvdYtVqStVSpuhULzDQZoWzROsbPMF1uwIWLbHwdLaEWMLj0W1ZlL4f5MjEZTX5LJ/pMzi0w
w4+AqnySJG2k8PRr/hB/qxjxW/4NVDc7LFppmvlY6KykxEK5UIKybJnq9JVAidnW+IXKc/Q8r36v
T9uHrClaQ4zuXFhzVpSQpkx0jB7agtMbSWvcpiu8NMdvcGtbc8jno1D3snIxDF4lR7Fp6++ue+BT
nWYpVemcQMZ/2qpWVQ9muEezLz9tgUlCZjyeZju9VAe205FqxlZHJKNK0/fBh0oYTL6UEjjXgS9u
Mfndun8QyPlcZ5WjNqYISBarE+huyDM3oLx42+jjUgy+zqJRTWUif1aX8RRJ61BnJdZ0BXL40zoC
ctnIZjRJDVGcNXUalRCnldsPUpgKickLlXUxhhaFrQw0KpPHdDF8+LDw7nMf4v0gxw5Wi1jsbOL0
kspzHv9fPBtQ+861zW+6RSVrtgVo37lgr/YcA7EWhWEqW/4u68XivEM4SK3S2bJJKKqQpeEd1EGD
ngpzUoJHXxslaIfjl4n1udW+wPHhpjCIDNHz1nOM0oanOo26HQN0qyu1mVjAM5bVz/KMlCFT//1d
vqTg3cgKVhiZ0Q+1N1jX9d+cUARHKvamlFRFD2TATaMmx2Kdj7SmwvmmyLRQLTezFatUDVvFGybN
hU9p8z/J1NRkU9U2VbG68n95jTHnpjzqN1TdY6h/gJP4golKPEg4RCpL/l4qlS7IObUP4S+Q5mYz
TL0YjNgWacITJ4Nw2A+qrlPp9I/EAlIy5RF1+6/BsEmNW2WA2+hr4gWU1918uvakwcU87Bzpmhky
KwzrD1XMEpxPP/tQI77nxv66pev1BuFTB+DvNBD3dI/8lvPFjC2R+VW7sJEO5LDpuoGe+flm+xoq
cb4q61EbvtMcYQPBvT+TNTjhANqJu3XMqCpS/Bib8fB82hIcSC9KT+GSe58b6ZFnsZvqm5vY11LT
l+tx6r7DzMA6UupnFV143cCBOxQ/t0y0z2p4ENfqBNrvfo46FT/8sgLXJacWH665Tnr23CeRWQjV
OIsOWIbbEY+vdSGaoAfBq8Qqo2s46/BGs0VwJ1JJweUS0toUWC8gTTI61Qb4R5Dm0XNTc+XS12KL
68/FCw4cqjtdAWbcYMzipKsldERDNpo6hr2AAoeLCQn78b/Y0khXf4QKcs03cSKOInmp2oQ6+AWn
l8jU9dxd4RqHPYURuZv+NJMnpRxgIEWFHFaZMagpHZQtj49YYYrrPxAAO2639ELAl7UoELZIZtue
iafj4q40HqIEp5GF/xOyv9amcspyiUKVJJQDTHMk2bmy11vgQAN27kizBzaeeypLElef4RITXfWM
gSx87s02oNSvjuTqbefilemoeyXLsEA50+9PymYQI/WWMLd5K8tW+ZNXwHDVvrNcwFOVZGS7YECq
ttpj8ouLzhqnx1WZoeLawlJEPngV68IMpUfdtHJG+W6lPNa8kkKb+OzFbpwO4nAw90Iy6F7SqdDP
/IFTAUXQlb6gwZB0fh0javEOuLClifA/hqR9y04ZxtOfPOFTnLuCfeB7qLiez/3s66fbR/IlY0nc
tiA4luCVML3mMK6XDmAWYwueoMY/e3XX0cfpjHTLSzK8IxD4hfYxMK6tYF+hAlMF5U2YhqXyHAzk
kjHHwLU0Q/9Al9eDrjQ/qIJmJybMwHCcf3MUpYbOeGGGpPgHk7CbzfokfJe8bOdSeF4VkmeFXVhK
gD+uAVhUFUXvXR/IhpvY2nOmyzsVePbOhx6hwYjfcKNuqmqcC4IKkni1xSHkTBi4Uw+VQQ56X5Um
hXyPkUnN1+Es3JCzIirtdbE9P2wV5FL/Mry38MROCrvtD02m7pCYobHUTaOgPAxNyB0xE8Is/9kF
nkpd1+CeC4T191EWQRhZmIPNjcFGiheikz3I11jZYW1r5H4q+2U2GwaBZvVD4IQxrEMniZ7Zfv3/
WYRuf53ApZCNaizRrpHMnnRTA2kRSiLnf3Hsqjz0vxPamWXpKy2RZMXnV9sWahta5Cw1qUKlm5le
JF+oxgymeEvdeGVWz/MAzb2ovXFboW0aJNq6UTTyXWKTzi/DoP4/rFmEpdNxRpGP2GzKVKAeoWt5
XhU1qnqn7T3EUxOfLn5asE+3OweGcJGqaBg6yEqk5MIdvDvsU4i4wg1Oljqj2VZgPthNPCQTMWUC
+X7OvOKhuegZPfnTo2MFNIWK8ROeiYv0sob8HvOejv3u+6drAC/I83v4uWACTXTt0S7Gs+bKDl7v
tRj7bWQTuk/4LupV5PLJ0igj0oJoW+lfBzpH1Mvq3xHVCjPnuGSzHaBOnKMhM0LFlOqa4oy7KMTD
gESVWIG/zU1joEOavIKPwh4Ghs5m76XXffLFGZ+sXcByktz2yUW6rz7u7ccDZrl23hFiFu+cnp4i
dC6yrUKp/6xOt+QMubJJ1zCGQTS23GYct0GKhxhtYn2cZuGzz6irJIGbjyXP88hOt/T+XqbBXI8M
0WfXHZckFrjyvFJ8AFT4nIZgEUE40IyoRStl2gCuElaBEseAXezdQ44D9qJc14F5Xa8iYW2D8ETc
rzgbV9M3J78se3kpDH8Ex/0Y2W+7gIYCior9wkWpQNKMPBvbqL8MXtLvqxgRlk+58nf9DedLF1TA
AgqNKrxkSdQjbF+2b7ZGPbGlOWIEyLzU7CWFCq1ElpZjNMqo473Jch8UUjwXGcij1cjBJS3Leg4W
uQ41V/OA4bKaIG7I4PelOrpd//vhzp1NvC0GQzs8HBKWfnOEgIAUZdKtjJw6drOiI5D75rhlkZoO
4mdwtXh3Zru4z+h/i40Sy98Ff1iNE9KBGQvVxOcl1IlAy56UIl83jWzhJfWtXsSypwKIdrOnlxWV
O/5xDZkAXTYYjgowJEzfFgYOC5kd7mUuGum+QfRF//9fF1MByGqkGcYbb108R6HVT6fAwG6QbwMJ
PC/3yRBHyxeCqmaK9Umltwz0lZUa+gO1enpNrrz3i22swcsIWPPTW+PC3anjFQUG085gMumhBOKC
cSEaRCo1KcrkEpxQqpN2ZcsGmgpf7+P1mlM8EOPmOpfpmTA6IdjJOCXukpU/iDoJeyRbuM75YDUp
webrCLyyNHscREPol0uG/tGYFrmR6iQ7x8BXWs/jJizmmka/fOzIua4eAU4GwBAI7lyL1p0QjhBp
rL3mXCLJtg3d9TCpEBWRLSS+jeTzsbmVCdt6F3TMicY1ByO5vH/VwRjAOxIbO9Ezb3W8YsyOzj6E
Xt3NY9htYjpELBPXox+Q5NrqYiEab4MWn0IM/KbKzQzqzucalhW011XxM2tmexJznfwZSs6pqFZc
xONGqvWfLOGQkx44DBAKionvPjCo56Ms7fZGDLO13yBzf1YFKccyJ1yAMlamgWr28iKLsd6M7CTA
9U/JX+3CdB9lvCkWVr+WO/lf1zM4F3ZBkitoib3bh5UxwtsiR0ZWiUDed0K8l9j8p0Zm28kE8kUH
23pp65upvxANWDXMR9ieKT65JB2b5vLRFYvUVtldwhcIm8E5Id+IjxGEe3QzaVhLiYxZMQmdxSGs
SUsuZU4UDPFDPB1hnIpuHsts5U+xLMjKAr3RFjwOzDDyZxlf72FGJcb2ZVjabUYWFqkba57paENi
ue+ScgM1bsynHX4K5FbeUSlIwpSQHAWUgXb4qGUs6YNEIR3FvGdEVaR0TiJKLT5JuVKQZpGgYhfn
Yb40jb5LeSd35TLbwSiYy6hZZiW5Ll/Y/R3eQlm4USrq6EfCZ41mRnZMeTJ8qrw1TJD0+uXxd0MK
qWkaPOHt31wlw+MBPhf+q4tFgWBCOV/qOb66SxrerTP3QdjpaWJKbr5+pH3hEiK68TvgjenhT744
ppIIVAK4HHJhMtT1guyhuO7/kzQ+ZwkIPAolZOioOLwtMQjEAdBckYKO0f3Vxmqh/61e/eHkZLS0
OdPkXI8AESc8rlWZ2CBAn+IHF9ndrhjT3z/C5CrZ+DGDHJzK6AOS2IH7ivpiex/yR/cVG/hmOcSR
vhOuT+fqoKH69IBN2VZd79ok2L+v0ne9a0osN/sGEM19Ccj/k9RUv9xzNgiI+uc6umjs3++FmaAI
XG2t66+IZZD9vthGgwqeSfIEOa2K7w72MMOtzsplV1OCSkIYq4QJ18NMcWANamxfuzYSYAzONiDG
GgkAHEl/VN+sgu94ml1nHoSWxRcEGXacZ103spoAtLbT8M/YSxktja8pBnvb0e2focfrFYTDGjH6
TdSmsZC/r6HI+CLICaLxvUO5snRmLVGP0XfqdkOchHbVx/G0FWUeARFYRBgdBTCIykl6pmSGfKCg
ehPF2kJvcX1eHuEygcnPtotSBNhT/4pq71b5CaVhLrkroRYr8kLoEA7IcDJY/x08FntAhh2ewSvN
LcpqsVw00oKbRTjyghbi1WC+X1XQsyFXRQVeTuLwDTRCmp/Y6Ez5/YLs+9jqcLC9j3/j/7k1sqN8
br+E/3jmlZWE0G/MqYuozeDdy2iQtO0ZQDnEi7c0UNe2BGXkwNEWwhFwMrLWZjca3MJjIZwYZExq
GYAOde4T6Sjppy35mTHoHvEN60JW+f7AQcXbfIwjbVg6FaQna/T1DmGnFgWOY8w0iMVLkjafHp9G
nLh6yKLMiCMR5GYkUXmKZkKBvD4oZlMfjgSLlURaVAK4Wr7+HdpnOkEXC90ICcLDBHa71Iy9ONY8
tF/2tO5NyGEeq2o6Y4tcWT1CkqgOOLqh4Bod5T1hKwIgxGKEAU9bR34piy0EGfI8aofmxpbTMYaU
OFiuZCoKRjrWoGz+PaHlDIdLoLOGs//S14XVH+x/tLmgJ9zaasItV4QU5uARkOeGoMlRLmLnJdA2
oMvJhFi7cRpJvjqcEszLkdZOkFudhk/489Z3zpfS+QXJTDqDhQmKpJKIeZ+Tc1RRpulR55OEjX9e
f1udeALGg7zDHiVRDaZxH3Edvh5DNGib+n0ei/33kXxZbGc0PKP8blbqkkoP9WXpUhnmkkML7XTk
/rchfYpOwvsCuuI+WVUpdQQrxIBOhyU4mFkYbGcwt6+pv6Lqh4pYFqQtlrT0LfBFtuU77290NMVI
RTy3fmD9rYctgY75NpNBPsZUWaCmVVgZY1jMgBV3nJobztO85l4Rubr0mvhEntrjZGGwWIbxCFAM
VcvRTDI9f6RVVfVP2ZzcQD0BE5domtQt7u4g9DMnzgL5gQDiKyCuvJFj1zwWYpTIsFUgLF674c4D
KIVKgw40ZyNFzvqClQDlg0aCd+9Bkpf4aS+Kcie1b3cYsLf23tCU5+8A9WgM8LoPX72v4bjlEgB9
xjHElmsdq0o4WXmnpULqBZBSbwsYCPSJ4OnkvXZUbBxCVMl9rEgZYp1eLjtoJLk3NXjpSYO/Rvbd
NUXx7JaQbeCkO5HWGwkteA0S7a9pEGs/8BHcHNBCy7PodyCOTDP2qDLFoRsIDztaZyeqcrz+jAwz
Z+Dfgy7oBhfO4wu8COTZXGYp11zLsKQvlQTGRWySdd4mnS0CDqTXTFo5CL9mc6ZiM/chrXtRM7q8
vFnsWx46I885d+hWF/eqsxrDqjqz3otCEJxc+8lGKjbECEEN8G1f9XtArLHbs+aK5KzqtlSIkQ9F
nwplSrEELGI8Rsty4DWDQFhgJlrAtnFgXwLIrYxEitIATfh3wxWlswbDLWxZPTzU9BWWoyH1HJ90
Ro+srQ5y5ZK7AwXmoJsPcvpFTjbul/fIZjJz/oUA4RVp6O743dPB5dhXXJc4t6JheDtb7mxoy1rv
VWq3iYpnczn0BVU4l2fP/gB7rqLla5dgx5JDtUQ5WdSImnUHE4QtNRxNrUgRR7NnXJkKndt4DWT5
5NK4tTDphQWcu3THfKJ/Xz95Mf/Lqc8mLzFWR4canlo6NDK5LwhWCuWcf940HRJbACBw1oMeUfrE
IZwkm4h2+uLI4T7m5qIXrwbMHDXpS+a8vQC+xLT/grbm719aWy6dUEatEEimi6sv5/qxCY2ZOL6G
MwTPI47Ghi03g0iJ06JhRfQuXk/zeOgQ7X03duUy0uJCYpMkQ9VCY+j6nHWlnDKOy/Myg1zReACL
p8hft0uhjZ4Ds1k9Zzc1BifvdV3wlGUKB//nYUdujOUVaXgbRNjaaH+oxUxp3SewSM3qbADPERBd
s19b09lbN6840Q94WufouY3DMJA6q7Dp2VkBqfy+jelkAU6OIHLW0MjlD5V7W0cwpLZ8c3PeSlY4
L227a2Qqk8PAKwgFt1b+xytauuLnnpwBG/r31nK2ZIhXX7s8YFHnSPuv7wISly/JTp940zcPx4bP
JnZY+cheFuvXVyy4AL+GzzFikhsaYpMDh6UNMtS4ff9sf8Jg3A36e2k2K7hEpXvc/ff8iIr00eqs
qzC7NjBjY+wtqDnvqwOCNZlAJ8zmImUaYPF1E/NBXKPYsV0t45SuhaNLQopFFuT01kQqcYnX
`pragma protect end_protected
