// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
piLPS/MLpJn2yzkhvgtfOK4nnmxUEQ7RQF0q04C8Id5NGqIEed4R7+p+58cvcZn4
c1T/yBdDvQRmS3/GNGBiMTWP47q+qr+Jikt9HA0zvadNJ6IpLdXmgC7wC2I4CKFf
wqHVZtKN0QbdB2VFu6IjoeQvtsCXHSXl5USVo6bREwc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8048)
ylYMzfRPSmHosmtfqigCSc/H8n6jIlACnk9V1EglMQoPqOnN24Y3tKAS2G/Y4iSU
tXdiMN8FQLUn1kVTWA+eik2rhDpptRVlP9XE71PIGwKOY2sP2vplBryatKuyAADJ
u3oSI4/ObHbtE98jiZtBs4VTKRUUGQUPGWTVEkDi2EMG8SVCyIW0WAHraHVXI9Mi
vyc8xeJckFG1GOmrLeEZN11MPhMVS2oKwksAjVFpjobxFVEmpIczSylDPR749yCK
7M6gGvyreArNKkzIEUPolbcp9a4UpbghnEPZz9T1AJEcLmRzXom8sOvbeLoS+CPn
vIAK3YRE0PL63EyB227GY/CVkGWCD2dl6dNiFjJ7TzckL7cGVpjryJXG6Cjzkzbm
nUEJqCunf/01MfcEllLRm7InP7LuUx3vTu+48PHXTZf1l+I6zWOo9FYk82wxDJcZ
G/6RsC/xQ7dfLtRdGosJsLtU0CRsbXFx+E14pdOIFXn5h15zMauA+QTL1B7FDHZS
tBjBCMNBlrbV4aM6in4cyCVsS9QPPB5ucZszUu1a94S+nnaKZwAzXhE4Huu5f+wT
hte1Wm6yYBDo6Hho8d4t4ov63jzWtYDEg/v2qj5tkpDwiFM805v1PtlvUI1p080h
QZycIg0ySvLjFWR1fAhNKsrBhwY7jwP3T6VZEdgx9rPKbmOema8EaCNUqqyWnu+E
6PNTN4vL4zGwfiRzN+rt6hIsu+30NMkUYcgDT0yIbDy/sKxp3edR/4e00FolSFGd
XKjsUJKLWNAt7YbAWEgIPjRZvMTmU5oB113n/zmin4BeexpkD2eYY9QqxFRpKLDc
QXPiaIaO8HmOOxH++rLe01lebwXFKWi+vvETUtxXkQmq1DQB7jbC+k7BonXKva0a
4bKy1I3B7bNLSknSyXtmP6AAjb5PKombdmtgOQx3G0MG2TCSCcgZi4ECGBc+pu70
HdNUCdgDQQIz2ZHQHgniydyrvTSTTuhfbtxLUDpDKTzowN0FB9+KEjdP8hhnBtAM
q3KwMozqI10RpQt3I1ao+swnBhR7ZcayWL0GOziCaZwcFE5P3nGh+YkNWbkq2xPX
7pFGpjbHS/5gETSisx2aiHdTeRzAXwsL29aNUHiv2EwuY6GWdeV8MNxOkMtu95t9
HpGf1JoXo6LSUNCZ7wBWNOYDtebNH/yWBndLDHTGXuJl/ERNHe3yuLmcPYG6ak4+
SsuSxXIsezaChAd3bziNiw67KS+c2xo59oRvUZzJqQ1QRQWmpugBhP+Lh3QjN8xd
qFI5GSRaPyD5CuUf962hjUJwpNu/XtEKDhtouofDYWvvPPNHOvSm80gbGu3kdg5y
bAmCPh59+CQopPRIPRdBzdHVrJFOaxSKnHM+Q0nRySvkShh/I02mHN1fMSTiYeHM
h01I9bOfCA9FLrIxP3YcLraV7gUoFl+ZIGASe4KbOtB9PYfW5EVeJZE48PkxRKSj
E71Ob2MlScgcy4oCXfx+NWNXEnGBIIOJS9euLM8ey4J19XNIDme/HvzKIhpWoHpP
e95CP2bMcwq7l7VmpZ/D8yzq48ra3KCo2uP46W4LjoV5EUnrmjq1cPjWgsj3SAmD
eJoX+7P/tjsMFdtnjq8KFb6YLFkK3cCXKIo3OAr8PMSWfwW5//6ZTeLL35zp/7yd
BWfNWgzYjXLd/goItDX5nzoVbJDVRj1mhX4HdhBa8DmrkZcqerlQqnjqdXLUZAxl
m117n9NUVV42a/QU8gUkkLToAIDSymLkHj8oWs4FWsG+l+domBQdjJeUBq0dPiQY
F0ML4644NOIjMa+9b1pSu/gzS4hpsSamPtGJGmhNCH45jbsQEqHk/Xg8lMNCe/am
GN354+O0z75WgyjiPB9QxO3kXi7cDZQ1JT59u/VhojbHNbFfPVLzMCYf35cF31KP
OyRzgwHtQHDyQABui0oOV4BIgmg7loch8ED8KN4gs03jCI0jIIT5sSjgTdjTrY0S
oUBWrHFvMfiEIbQGR1cpp+3fO12rr7gpQm9G07toHFrEk/NuJk/H0oiS3TpqY95D
SUEJem73SeMHWo6un7lwIl25O4Fjgf4rso/ZTToUZROtwqoyx63sf+pE5U5s4eoK
rB8+jL0c9hJlRnjOKzFxmhLfYeseaYwabsy5S3yRwFtwAjkMsMSwK7XEiPWSd/IT
mezWLwFU/FXVGLAR/Tt0daPIzlDhXvj0DB4y7UmF8wb1u1BA0o8QQZ96IeGiY2Fo
mD08qbQvhzPPHWyffZzn16WkjG2UMm26AO8PjsdKvR8gp0J7Sj5z5Ejpcxb62IgW
tcrz9mtpnptlxQ1YxkoLAJckyidtW5m0w2AdzB2rSrdHM5pJn4+jYfAOx4K0GuCU
YaMv3IXRY9XWO49SzxSA8my84gXSXGXJmqYfdLxmxP7odwboekZpfNDxFFdUbvTv
Le0wg89HnRbY3Il0MBU3rvHC2JLs2TNp/OrfqFyJxkY2uHGTaRfCkzwX3C4LBAY4
4wr9KXbF5OhI4V75S76WQdo88GB1uFNXPpxsYGvw9zd4QUEj8CPik/aMxSNFlE+v
n836WkUlHzU0lYdsuk+2Eti+8PnenSKYwI4W3aSliMrcWFRU6cJogLdv4cIIJDad
efCYQ/5nmYS9IPuVMxsB0nK8xUyZ+HTXrOAeCHfiFF7AYgFAnybCc2LXuU21pT3E
S79NOlIEH8HyE4vmXgGsJwcQVfAfOv5g3jiuclJGjoOJZJL3BClw3dlbwt9+gTCa
l4dywXUrGi6k0cg5nF/XOHnGAfbO6NBJgwbgrt39V5CC+aV0s9oevho9paR/3Ynt
gCb8MK2gpfYY68Wz6zlzr2ddlNWrSq+SoM5iBNqAoKw8/s+ZSJr/RgCyNMqU6unS
10BQT1gmeGEvl+FKKNWFxDV7O77OeJvQS7Jh40Os5/PkBv+oiDntbLiW3hIvXpRo
dmRFtT9DU4P5gYxBxPwq/gJOIVZyB/q5YW/fKHvlCpEHaFl3CI7MuNm4bvixgo4F
+ic8c1/ZA3qd32eO8hzN7YAKLbh0nWcyBo4xfUBgnQz7gCKP0XBaPXO5d8Oy1m1K
P7ZJ+Hj6mcRWvD/q+69NQOrxgWxvSBhPDwesfDowU5fPYCNvnJ5oIlPThC86622S
GbfVkAew5R9fzRP9P4R7e7T8fI35l/pNkuO5hU7bl3L8Wr5UGdq/Bw9y89Ii8gmE
CCIbXMr3f0pEnoMuIJfyd9ZRhuUYr2/9BbyHV8awzPnZGuTNjB+LlFV3SR5ufEbE
WcNAH2VZ8FMV26P/dLP+z2bJMPSDglptUxEID1fBvcA2HwJJmS9RKS1sUd9vGWQh
gWGfq1h3z13pOCXN1uETcMzl+XmjwN5nSXXnfdBCXNOiNcse2Vu+5YWP7w7NVTEZ
YA0zY7r7LbgykTLJXryCMz0hQ94i6hnNoxeyoi6f56GG7QgGPAN+0oPkRGdRdSvV
AdpS7BOq7LDnDt9FojgsiIA0MZswiK104/2dgLcImpwK98rltgHKpaSLqoOPKnW2
PQizJnLCUHwB4Hj9FgIsWBmkFe+hUuU1X7FkyxMXFvYdkK9O3uSyzH/dkuBcydB1
LZI3F4N+rZ589UclTZpCtjit9panpFMwVaVhyiqG9eeUZeEwUTUCHkB5Xi1Nzc3s
VCBZIWDfEbStVnl4QgtekVFsKcRGC301OHJInayx10s5maZjMDLUd6WtXO3yH6/E
1O5NYtDVweNg52tTXNFaagRYQ5d+1GclZtZhEdUeJrc0LZF4W0WVnfV22Bg7OWCc
ELbAMapoAt+1QBj9jvAAynTR7ZOuh+A/MzwNHzvr/2m5Ccooy3/vq9OoSUmzEByg
S/Ik5kFX+MqBGxK3Nf0vACddAYBCUU9lzRTFvKIb/ixMnyzUQwMdCumsHiXFnpjw
V02khmU2HoF/RkIf+UkMmQgOuNTbHMgVvcqUlKNh8tjybYtEnLwlRjWi+xoG+AzG
/Jin8uPyZSRMZmBTOoGpb8+1sqGJV7JLRqXZnqc6tYdZfL0nmw6kEPGTF20CJDFG
wtKK1U5hvYMs81qw6LVyDhdSQ5YOM4LiqzYHMLl98LCw1ki1cHKvobc0D0Y/n+rK
zFbPXQqjPCDM1etngB0eTOvOemIoCwPJDTJ5ZhhAIEuFCZewQTVQGDGHG/1QiWMV
2zmeFPLxKmaFjuepqb5uF2WR5fMpDxHBqeEhFmGAb8PZQD/dU2OF6aIcglx+Whvs
+Xc2ilB7zGD1KLDbtvO/MIkKESAcaYJmjDZkIJxKSX91Gj8xwQeod3/u0do9BYD7
2fTYUBBpD1G18NLarhjUrbK+9Tw6dx9mABWqKZBA5DUwqeASb5khOjiqdy48yJk4
TmCgBPm3U0hzSxlvJZkTE7N0Cg2J9THhU9a5JDfRyRdWpfekpZNH6TRhUEwPQAFe
8u50rqCFpIbV9DoiYIxqXTzPpLEJiOK2vHwR20/L1pc1kTJu/qalVLwcMOTyZvEs
AuHATU2Q8nQHTw4CO2hUOgaGB85xjP1YlCMl9OO8CK3UhrKjV1MBMP4Yvsvoybzy
fwGGLskPd/wO3ZKeUlWs5vHacn0boJgIhcwjJI8Za0610JQmnYidYVgcoL9DCzPn
DkCjeRUbP6ywZOtkk8yrNABELgUsL8rqw2Xmf+P6o9CmdcRbkyb9eCTSe7ykzJc4
fTV5OAPDzzejzF5O2hcwdtKT1CzXt52gAfp3Huwn50Tobd7lSKnjsVmlRx1scxPO
mV1vJaXrEr+4zYxwZ1Lx6bj7xCI3Ke7kLSV7UYTV2o5xFWZf9furzrq0MZ4boSum
zwimzBXEheP8b0mmO+x79q9iwgGGql4TF+LKWX59OHkoIZqG2bTLlgL68/g1hwvf
XbDyK0EV0FZHHONDpO8tuSjQ4uI2KLzClf7zguubjxl1CRQ3BRJ+yCeBDw0YmAtN
vYgbIOmbsZYG+d30VtRgGhXJjpo52ekNWru2oRTLEyssOFfLrT4nzqp6gFw6E43V
FBsEHNwD87Ko11+M1fNg9RhQgv3noEimKc6Or1NIEzfdqGji5lIHrnf/jCbUfL2i
okpIQsZhbSKnY5yxzbhpfxuJ3wyzro1K0fvy1bgKBL/7ky0pgFWOTGUB3GPrVXhW
uCnL0fM15Plzh0SkMO5K18iezFOLxzORBYxCOtG0JxoqHpk9lp8Ph5IS7+BBmd3i
y8n9vKcoGIwn/xRaFaFG7KAKl+uBrrS+6KGZtbR5geUQ1aYs9rzQJPjP17P6+6ZE
kk8FhQ3UnH/3gkXZYqAA0Aatnu/IcrNBNGx0xwMrJTBPtupuZOZp3Om4ltj2+he6
x5MEMn166eq1anzJ7/pkI5D5ci24N4xKHEpEYwxCqtnvKr+qNw6JWmVKJZkhRYAG
NAloNwsoT8MCfEAHytRHmFUWbXlW42pxHnyKeBUkXaNELLe4+yDcj4G+k/2xFuQf
1lGXLLGORbt4R+0arNIqwtace6xpfcwk1mQIPzQnG065GD4yDoigWbgNQ8TkzGbe
dqJX+vSrtI3gMzjzYssh0+WIcGjP/lHw5QIIrSY2N8OQpJIOd6lriyuS3VbSYS7F
hjwbL1QdEbzUFezGAgunU9jaeQubxotnzce9dPpFTACuKl4zXj34m3cnIyef4XOj
OoqxgJcQicZx3sKCLRMUY04eDODKptpwe1kx9fx8MtBS2yGAgPZZeReTE3ViGQKs
Kvo+RTcLapXM/+t526edCmrGfqp+zzC0alYDNk1EYXskCKQbT00fi2sxkXLS7raV
8KO0gYhHFOrcjWEjgrVVrcoiNK53ajJ1U7Gj0Vhp0E00TjX4UaHHQRD+ksmnGDjR
0+5U2ZZkgUKa/mgIu/WzZFr7VG+3GmWDwl1Q5fuhdDiSFX1lM+uRqsTBlodkuUnK
33WM7TvGIQYhcQRpuTKcbzOkUm6D+yERPjvSBjgj0CsTwzu/gA5LkC5CNfo9stbd
4ifRAipw9N+IOLDrduK90MDHTfVyG6NJFkNFrdRdWhb8jFcJmS3v0CGGdgTGCUUf
hIt7BupLpvFxjsPXkz8j/Fkomogo9TLokXpZES6zozLEhKmDFVzxSnEL+2SGEi4g
KfUG+Oo4aNW7/B9qKlmUCPFeXp+HKNYIEmh3rs5c8m5jlYEDjaWZB0EhNEU5V3zr
tE50J9EQvmSaPoylZO2MtSRq28qW0pYTky+H+21hjW6b51idFgUltBKc5ufKuWqf
Lxugk4iLz3EgQXNqP0YZjzdiQiPTQcQTlEbfZwgeZ/zddxAJBGobZQoNGq5ynwIL
bE86ENzUpXa7xoGWnLDxPrmUMnBQD4mADQMJdiBK4EW7fcf0jhFCvcUweNK/gpu0
BOfmp8azqk1NrUSQALT7kXUIj3LgnpnEMxud9yPMianwAtIsKjN0NECZ9bSWWyuW
E7vrCC0mW01pfzptkMXGk2CjfDCUqcYFuwa0kJNpbXYJX1t5/aPyHs9GhlEZyrsp
9gcVVzlFUCNfoulY2EBUx/A7ZSXAE67H8ERFjDsgEEJdD9prTuKOTverH7/8R5AM
BxrBEpZrNMn/BnkwlEpGz+BfLHsa67QRY/pqFnHzez6Dw+jVhVVL68C7gB2OwKNS
Oa0J0YOZ6qMOhVj/LiTs1+r694ikXqOjA/rKu/9WeqFCWhEH0wTWPlfj27ho4IlY
z28Q/73PmVZN0rOGTAYNp4BRXbXZhT0Seu823pvwO9tq5YblmkHviXXhHf//tLI4
phuIPrOPdirqa8QQU/6mG47HWYj0MZpKdf6Zlqt4JpMBna+ZQGZX1G64W2/NicyK
xP0qEAXhva30twaPbvuc/sVGTJF2fIo8iLEVYuOBIML0RWxSpdrRG+GA80pljzZY
lM9jUhtgij8llqY3zvbgD/8+dXegVr+xcGXn5jrRScUg5ozq9w20HEmak2bnJ2ZS
HiwJRkRhV4zUvuz2BzQenoGd5UpNDOI8C6ngMWOBYpWje5s/ZEwqx35H8R75DNGl
U1btHfx+D8Jd7Oj+Wr9F5rxvFckiLh+0ACXKF7eh022BRs6XTlDPafkpsBOJ/SCr
hKZYOhgQGpJbdFtg3wtn87/Bdc9qZcqq5ju+2k+2jVj8gvBW+/CGkSuOJacBpomS
SQSJVliPchqKZNrHm97jCJzaEgska8zrQPUCZLBfYG+03WtN5/f3Mhn1026ETnzl
lpx3lYNzsNQw3+XJRGZNrxudjcRVgu981ZPIcQagekKec/6E22HVkF91ekzKud/Y
p7+/RP11EU39Emz7SR8vte8Gn26XDbU41Ff5Orahahsq/Z34PdlQ2AxrEkRVlDnG
HMQI6rGTbDb2oznv2l7YQSAqWs7/ZOuMiAO81Sv65ckvm3oM2R7OmunkpHshqloB
AzSqInhaCFy54FRGr9J6ohuxtpBQe+FVoWdvq7Ed7c2D7CzDN9cFKsXUN6rEyMlw
7wU3freWjRK8iRxuwi6wgGFws9QEpLRHhR4v/mJXnQLuaNooa/YD2kpG9cLcy02Y
wJTo/+qFbt+Pfpo0MIIZ7IFmZHQOpEkV7aK7J6Ffm+9TLZSVpXJSA2GvFj8SqL44
gfDU035ZvdCv+bArdiV7tfbAtEH+7CmZWLPp00GfHHXEnRKRHFVsXNvLcRA9k5Oo
5J+yqUEM1uyrCFPxfIE+S5O6SU1XHNh0OsHJj08XPXIuGygKJOYHV9tnopNGPHZ8
HdmvtaFKvvKQI6xC/jZQcAgTlhtxRS78H4g9GWVbLBiYX9oLbktOyK3AtW04kYVN
yfY22YJd5LuxKNpscA0TqUwzznJdLjykCQTsJ2/wUwenf+f6zQkKcr0toSrhsZo7
jqgRh23lGnei6cVLO2pQa66NK/48aDLo62wvDmcJ9bqHGEleUWusII31pPZ0F3mT
llQfDKb5rsFUkA72wrGhHl/6Fw1XWi5lfl2ZiGeea4tzj36grgBZqqwRP94Dw40z
tVVDNKiubRF9AGlWrLKQlm6Ew/xen+e7/Fd8DFsReiA0ZswfH1uIrbpGTc8Q/2sC
WVpstC3Xc5I8eW6TCLT0QJeGTR4C05mvaIWxjmXmmFlomtLDYJm6q0XADT5CGqLc
8O/zYrujOebpux9bi61r1Ea/zWSAuXT7KmkiWJktG3UQnIHgHBRV0FBqeXBf3Q8K
D9quyPauyKBjhLNHVF+DdV3Fd0FjIGtROiQpQIovW/NQDwOOeSCZoqkRqouyTWFv
Ok0izd+hdB3D5E+ilPMhs3NpPtcdagpAoilMfuBzE5VS4ABf4gZ/bmvToStc/ic9
BRNIMH8T57gfeboIOSr6QnXfZbVXg58YcCovHfmzfBdR20w5BEcT1SrXRndhIQvT
vn9EFaySILeuAsz8NHaRy924W23V0CDuFg+UKnNqac5pZhbO/zxyFSsEhJybtH4M
gX+RK982WQKDP2t3vss4Rf6ficudI9nnE2HJAWEMSG4iAdJmM9h825U+YbQwnfHo
uUJTcM2Qz+ui2sWDfaKy/yqAzlk28MLmx5A80YADV167H9hR5g3oE48WE/uV2kwS
EYPoKtcYYSqdhEFPIqBB4iNVUA1nveEWcD7Nu9ROSGbIB2hMVhv5dR5x6wvdfgBN
MSklQOMfrYLiMM8Bzcb24vrvQwzby5s5ZLwy+tpoX6pGLW14v3O7d9JxL2xlkJr7
ERgbnPNrFcETHwvdINGveO1UpaDGuMpX/ytGciukJRAYRRZZaXzSPvd0NzAvnp3w
wVcz73dUrGMtFzma1k8kA2e/VLbcgRpbSJtTGAC7mr+CDl7stNAAMr4Z+oTjqGgX
pzIXyD6rjhBcyWxzLzLl6v7OxiYnjeKYahrgPGzrF5D8TIgoK/rAFubCx6NxIJeu
ItWpuNBEpZVjxS0N1zGKaOh6XgGR/gIAXwKcwD+FAeqcKjrPzKpyLVC8WVJnZseU
COv/8ykquizdQQhEzBjFlMmomhm+oAq7ql25zaQB26dEeWgaR/qet5LIVA/mVD9m
//1pneAXsSHFyTWZalQ9hU3Kye9U4zbXDgXWDGkgqllpivf9mGschXmHUNt1Ydtw
HNWgFBuOSzRiiNQGw+JmNTnbizJiQjY4TFjKzL9jBWvNfVQdUNCv4AZviRl98tWe
7sgN7ArPMSKRF3AixMIVsNYTlrWF6O0LxgQw1NUeEj09hYK5FnCrbBbH+T8Wz2/F
isFv6IDidd5D0ODESIL4fWQZ0Ul5/bTYgQd0uIznS5sLNER62Zr8Hq3ECi8x6F4B
6jU214osGAtkAg22XQ3Fi76JWvYeapCb+YEdExzjtIB8Qx2b2c+pdnZJNYp8kTbU
2zozQxwy46XE6pUg9G5JU34GYwpEPLiEyMNbH7o9WCWgbswy4qYfnW57g6c2SaaM
9d1Z7ciCy85CJKpdliMchhMzspleLn9TyQw+t4Drq/G84ky8xF+bn7qVJ1mghOGE
VeJZZ5TDr0dcZx6Q4aFDV2IeHUodSIfz7ZuhzPFSwxXw+Vh+UEVSGi/316hi/4Uy
EXuGWvTfCXSvAuul30Po+MwZ1vEqe5eUo3XOW7NqgRhcSOlmdOQEq/65Ao/OTB67
qRBhFasRMziW0hPhztih/vFPYVf8rhDtLg5SzoBhjBKWTlLntv2nu6yUHB9Y5cCX
ZyeHmhuko/qt7S3HXslhOki3hRTZqQRBES5paW9xLVcvLLeEvgSLhJw+3ynNHCr2
QVxYoPjpv7kWff+o6WQ6Xv0k3KUwpvyaYm1kL8E0b6NeyEeu1g9FGEeMoi8H7Bqz
uOr2ZPweHw7IBelZZohIrrpGym6eHKwF+/RW2/pP7l16nUb3rF0khVLgDmetdkd1
iBOzuS0poau+uRO+py2EU+o37KCWvglzUs8kg5cYu1d/Wfi8rk4Gggx59KXHfUqA
2SHuHeqJjDt5QRwql1/iwlqJailuwbEoLYUI6UMlIzm7dKcTFBxslxeacb90CbdY
LLgfdBjfEyLEAOzDzEQvnzsBumjPwzzi+qAm/LgFIZ/bKrJRQSnzlk6E3Cj8bO3v
9MhltdqQUU+7OwxOaVRGJTYC/cPxbNk9n7AD6pSHx7HoTlBIF9TUDILsTTzxqRZY
KWDpe4uJfYqH47/ePV2lTDmeTz3uqlO/pIfDyWIDWJ/4c9AJkIhV73Ybh+v+wKUe
qqYZXznQGYnLWAs5+Lw6vk6LJ3uM+I5SROy26G0+RF3+FVTRVhZwgGgTVjEUNV8J
DvukwrPs6vxqapEuKK+S98EmYLSYDVQD4Xnzg0Xm1M6t5Bi57n/J+21zW6Kdip2U
tSkjqpgdzidL2YY+mu7+MC6YYG86Wi133Bv+mNjQyPy+2ZfAEKDwq/J8duEZHuCt
xV2nainRvlulrzLjqjqIOHXUCnv+3xmx1+6W9Hsm/YedHzzITJ3//J6OHa54QND6
AHmPkrqS5R6rYilFMTxPUUf3BGhYU6zpbzoRGguS97xWWizRhNOgwnXYO11VuYdo
0TaQ7MV5zX46sPrdK1+xR0Hf+ai2tjeLusxp8JFIxAQwtwz6PjhKcaNV8JFqOVvO
AZSr+GcP1EYMrR60dcNFP7qmSOL6fyWBl6Q/BhlfLL72+GfWa1exmcG1BcBiVOki
TkU1ahNcIOFVItRTFQ+ZBibBRLKXkohaJNM4I2Pozpv9Y61x+Y/hYhfl8ftzXr+H
i0dqRRnd/9d0gJad3eNu6ML/C//0tj5HR8HmL2bACqOPu0vJn7DTRHxBDhlPeLOp
VmnPTi1w3ctXQyiERQrocfJ9vf2N2SUYFbzUPiZo1WI=
`pragma protect end_protected
