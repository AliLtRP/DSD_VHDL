// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hxmwu5NlSr2e7BV22seFBoDZxXv2aAzet6Hu43alkNwRVisOVnpww2bfR9I/JQvr
DA0jGgKKUwkEfKQhybpG7xYjisJGyXXzgMK0twQRerbTLq/OlqV+65/EpcP4PM2T
zSw4tOweK1jRfpmzJltL0TOLxGML8OlUWFlH+gDY1eE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19616)
g3fCCkk+aKg4SywvPmEd56NhR0N//TfIwh7HwiVsb/3HRFaJM4FWwpLiZWoNhVYE
gU/gmW7jTFJZKu19tiKePE2UTW40ZT3E4C3vd2OZaciTydcszOSr1o4Y4x90AWpH
ryfcNaPwB1oVMUXvj697atD9b0m/Waab3gNSd+p5PIURaP084docSVtJGOC7PDxz
NDTYJP2KZLpVgrnNiLSs/1boNCKSDJhZ0qmZm3XXnakKKVKg4RzD/yagauyUaN7x
OC9ZQ6AAoXio664YLvi2U8gqZSlQH/RVBzWXEKPBTwdddm5BHpsSOEZKQypwO4LS
CrMxKFkJit9OvB0AcT+uXI46q2tnUDUaD1TJU4NLpm0DpDBXeSfYseCt1KSRTJkP
sq+rLCOdvN3O++RU1XWRar/3u5OLbqN5YPUBnpKwe+6ng2MBBilmVLaBcKv/40ds
FsVthKStMv59D6NUVTx/Xx6v8VAJX48zFz9kaWI5y+5phBGKLzbW9cFrvVt5YsWp
ASYWvoqmYKQGqxaUXBN+ubida0E8KD2ZsgnbQzcKY+0DNX/OFwdf0oDnBKzGBUTg
3/O6Wb26j9jaT1ITYnn5FqoevPFPM3yloOXVPimRlJLqPU8K89LzPSGzdcNYZ6XZ
JxoV7KJZyyOj2IFKPmWL468xLJ4MyuIjwp0+IO5vPrDj3P2Py7E2CelMNmM29cOM
209AxZOrinrxzq7EjTkeWfCZFH6Ec16k1K22r+jC/muCxA20szeVsbU+WmNRN0FZ
D8YLPmMFCMkS0V8/FHrZtjdXalY9IZAsr/4rXiJb5bk9iIO9ZskeAD9yAq9zkVYB
ngfg5T9r6IEooqerKGFfTwbQ825v7FBz3U0AjfRM+naQnPA25AE36tOuDRKIBJJB
VN3HtxI0ata6MtA6UxHB3mj6dHvbTSfjD37SqW9nePTCVVW80cDBqUT1X34zy5qg
yGv5tvo76JGnE73Au7dU8HsLYyk7cuds5YIe8tslWgtQc93UP3bJe24rOO69sYgL
VbXa6S5QGMrMPsFVNx1zkyKrCZbeNwH5OYtbSVBv6DWD8/Mn14Sc61KZ+VOFxggl
sMVq0BrFYkVftrErYH0PftUXYZysOR/ykzcWzB1J1wE+G+ZizZ31ZmzQWs27NjbR
5fWLARtWleu11QA+0V/hgwyFhjwvibpyP6U7dvGJ+zabsiLz0kJwuHiJA101tWh0
JhorfNW5ayeQglh4SWTfpdy9ihWJBKq6EQImNYFEWXdjmAD5ES3/AN8TKYWTTvLZ
wlC4Vy1cuR3Pw9iSIR1nq3WsFM8cltEVx6ifW70kr9RRarePP0byhPaBzoDkEVGE
AIscKuCtjqE2oc+Xg1Gm39pEfPOJhXNzaVEoJ0q2dvc84DKvwPyF/OIjwIV/Y55c
d1+VCfQhekfk3m/FWpQ6Tfo0CGgtb2t5w40KAh50YwstUZNAcnfj8J1RcbkgfCa4
MIbrG5J7p6vsYrBAXmFh5EVZ+wroiMIISbKI8i1+ybXn+J7vWqRe2s63L4hMq8Ak
pBowDrh76jhsSQjknvAqP1M74CVb/GepixBL24fKOjk4VgjgDqgsVXCHKHMWLe4K
P1SlNgRIZ5SC2aP97mpD35x9vzb5E/4CsDLe5M8e4cBuWfDBZXzxWjC+Fksy1c0c
QYwiUCiF0WP4P+mVDbPwB1nQ+pEZKqlB0aokBHE1d5q4L4NkJ8ZqoSp8P8xaoRxy
AjW5Zfq7AT8y50wGmZpX675sx1AT3mk7ITojkyt6pDBkdhmbViNgf8LunegJhb9R
BfCDN2b7VbpiBH82YS2Wu9/72EaHn3hktDdGaDT9tn9XxizaVpCJDCKY/vsaZR+W
I2zdUWQZBESdkLTPJZ0EeWEymhJ8bKeRoJlhj0C3OEIk/aTEj6hUU9ORph+0Bt0+
VqK1m4xezKs2cdWT+Zfyyuh9cMf5e+oAXzpWX3v7xNc89+/8m5PlquhaqrHzLGuF
K406Z7OHu13zCylA4M+t87dD4exPt6P4Kz2Lkxb78yS7M9gc5mnJ7jofWuXCAvbh
JsdsMCdawm+1vEwUwTn+jjFbwwe0vjBE++szbUhpowWJ60Z24kLszB5SautiJH3Z
hfYkC1epMPAlUmDYPyvV0N1JW/6t05vqlvUoUK9KUvwBCk6BKcKSyfIbrWmNFV0A
Av4zPXAsWt/Zb4Risv/ZjXNHoM30WmRHQYn8K/ChuwLz+QPF0AAbgBOojdKssU8W
eXvbaBy+/vPEuo4LGu5lHCIQ7wpQEmy8NQ/PSbEHMyydSvgkVLJZuMWJYz51LfAW
I84+0Nld7xnW+JXWoSiq54Znt7lCznjeMKKdCUDTOdGmGqewWHtsKoAP4zB0jGvI
9JQH3EQQlGQ8zoWEWEyWQj+kQSJolEzUoqnnOSZstdxoG0A4vZ410PLYtQXcSzbw
WnnQSHdjgbeEd1Phnhgq5jdMkJDGN060cB4IhaseGNtCGSqwEw8wNLrgew4nvV5L
mUj+eNRzBMCycVudAeHUmMP2HE++sanP8eCu2CORcxwFf5++ez84IUXZlUZ9yaSA
2/dfr877xHtozv5ziq6b6bn7p/KVpC90zQP9tcx8HngwIUV1AFBCsa0Pp58ZoBa2
tLxovENl/Yt3L8rUXTh9deL54dvXZusktFj/BGY1kIacqRkLEAzpwaAjVu7xPYae
1ouR8j198zzcetmwHkc8XI863l6p9lARLitbuUK/9a0VOsDlFEeFGkdRXSvfanBn
cA3ynILapkiKvYLqKdyIN1GG8STqcV9yrx1GIb+xTdDk9FR+jXTDHL68bNj46hzc
DFkKUFclPRNPnYdjV4bc6g9vsgLqIviUfrY1su2HDErYm+I+7WXzZv54MhuOGnFh
rPWKYKuaz26va2E3EbksOXz0yMWJAmHtNtwAO9Ui3PFv83u2+wFtjAi6TvBOrWR9
ELp/kvqdkVmcoxi9fEO9EVYtfywrR0jvZEowkGVVxebYoIzaVbMSOkBZN12ZSP5w
78CYao0A1bICKgeyZxIiisN20bqJdOUHjzy6W1GdENwe5Mxeaz8lAT8YuAJTmURQ
tmQnv2i2UfTXfi+nYULT6WFEA8kz7Wrxpww9jKyxeYEttxLlwurTulBbZc5hrc3A
+5cLjpc+Bt0IjTi28RMPI0C0YlCABicg7e0qSxqTXx7oMtXNTeayf/kIonZdq1uu
9kCHwW5kTM61mQtcFDaeX9AuRqOoIS276+Kz3uxhm6O/lSfuNCcUlzrxxUndM3Ea
Z+A0qKPemQtxnFLvUKtx/9OgexYYvydGSSUjviWCyCcqPDWauHH9S1kTv0bsLdeh
w9J2unaYgIEIvS4iRzHCx83U2Q0hMbwsOB2EZO+jHDTcusxZAUAZ6Z3FgdVWBd1U
nZuRn8rFdeMxfUI+IbKBPVA+4e3gpFZr07npcPJukDN5kNPKqiBGfCst4HHD3ArH
poQSCnxKqjzz8hgtxIukD2CJWIPgr95jlQ9k7GiZaSZiQWsRiXeKObysfXgHfLpX
gP95DvYA6YZq8fHuKvrakFRDgkAjNJMINjve3SJpvCLW+lOht2qIxHt0BxLDWhRA
Lac0kn4S1QK/5A2jwSOYCo0PpEquYKhlssVuiiFmTt+1cS0CQP4QU/pfFyMOYGX3
aEclGs4Y+HXU3isEHhalM0W569Y1gU0CdlIKOhZPZfnvOy/Mkk+ZRuQ5Lv0tssRv
TYE+/uBP6viNFR6TnYi36KmkPrlxS6njdspHlVp8TqhFb+oDSd65hkmUExe+Q6Do
s/eaDiSzhQ5lKEeCpSh2r4BY5rfll83atGe1o9BGsl0uRaF41c6dYRYy5BUG84ZK
6TfJllHErXyKodib+XxLgpXoW4cplgWHOFDVYxedlyS5i8Q7SPVRGGwmGvvmpowR
unYefCVSSQhLLc5TU7xIAGKxn7bdRN3Bu6WE/yrNUSuyNYaPsB7iHmU0Lcvzz9ZP
FuhRPJij+Ov1xWZsgPXMrGnrzhjBYwkPEcQZo1XKJCMjBgx1A86RbRWbjGEhKJAn
J85ymO89ullVD8idN2Wyvg851b+NNJMLaTwNKicIzD1axdbYZSbWfz6pSrGUXwa/
r7FpHeX5Ja0k4ZcJ+S8e+/J1WBtsRLeGnP0mrxE1NIinN0Xhja+3JBjpJNkGoPfe
sOaO1a7DOdU1rVRt5yRE1cajiJ3uOyy5BSf59D+AWOyso8o2nbvMdzcjZ2FDE+Qw
vn93FKhmG9A5/Wwsrqg2XZ7rBlA8lpdTmKRaND2GQ+wiLPSkD2cUrqUPNKVmlq/N
5T69WKDsUnSkxkLh85NV4oleVbsGg6AcOu+FwvR1y5Gzg6NCWQUUOxWC+s5ysHnQ
ZuYP9gy8u4neIuVyn5Mj5KGWXKl0C/FiZq0aXTk6+mfoosDLgKW5dHtmZNcWhIQl
P1vqGYs1FhgMMDjVEsDdLeBgMHLwEZkESSRMWGPtG7ElF6CvTHGrB3GiFEbpgcur
uSvGReUKOgb0nKArLXpWPP5JkwlwxWHExtLgC9aldmUsKTlN2MSoh7tSpnV5aDm7
SSeTHO5psIRKHtBU499FErEshUBLpJKeVmbBnmwId42fMo4MzADs+2GOqjynyOpp
sPVKNz4FA/vEoC9gSsRMCgv+OW6h/XajK1dekwDw125RT16YVLzGiDkvxy201Bkg
+h82CX5h4EGa9zotFqmTdjkTZXgu58wVJk7fJvOLECRHN2YKsXT/py4BR9wtMsdr
QNvjER/km3+P1xSG/i7ueway9wG0IC4nswkWTC8UFQ2Y8Kl3zohxHfv5ptCRyiPC
CwXOrpXRgMw+yXExUSZ0YwxSttgRbR1ZiWDdx9CMK6E/aCCebhvDLA+0ToAmufGK
8rZ4s5nzbND6RH7ypsUttSveBLaEBLlhCwPx5UWTX8XBJjKq6GskG7SiPvrrPmBw
h2gy/zl9yZdyXftpBWHzbnud5mUXdlKhXeh7nXGi0FZkbbMynBnK6MlpmQQtQ7c9
FqJN1mSCAuApCs6nr1c3qpVIWhm/VnRMwQC864ERZAxxnaQjRAM2t2rFdp/qclhD
hRleqvf5dWwwDcak4PzrRtl2OK8IS0xjpzTKqpNN92oSomli87HVyROEjo7+e19W
oOYx1zqxe9Ej52Aa6U4K29XyDxDnepY6S6yJ3Ip2qLTISegHaskKjx8W3oVNWPqU
WOgf7O8bnjpWas6qWihCeQxDy0/jrlJd1RDzw9zwahgzMa0WYaje1NLJVkshKlnB
yczfPzcmaSiVov6rawJ+NfopxZ3WG4CMnZpqM+wKOTv74TXBPiz30IpCTKx+wBao
JDVD7rsweF1GOwxdxo5Q9ra39XF5MlRpDzItqukJftCBjpUfAQxCEvSxxJCumhZS
IgO7MD4L8NuaTnyXTs8xtf/vglGgGq02XFVF69RvM+TU1oK48kZCkP3e1JddZuLS
PxegfBoeRBDf1bq0mErwzSbqrPJvrFGac+Lt5S5sZS8rWtY1vWjZe0vBTxN19e5V
sthuPiz78mwgruORnRWp21uM4cn+hJLLB7hgcupW2Vk8a/m+YGcrS5mN8daD8uXA
KfAJyZOgi4/LqhseMUe3qzWy8Kx4ez9wu3j11X5rVjY4gCiTvQxUMfmUKqbHu4oq
b/TSb/bjeb1+DcPls4eP8aBpjG7T8SCjkDdYrCWOCXMOSvJ2ELz/N0I01jcnQpJA
n5CtupLokJr34daNwVR+0pYli7AvlmNfnU/gTViZDMnUIP3lDx0fvkLhCQjKoyp9
JgxbMx6VN0/a/QsM4EzO977TwSKeSxQwTH1+du8JnYmO4pxxHaVyxblhdZr+ifUR
l3GpQEtxvqsEwhbYhVHIstJqSkDVlKnmO49/pq1iFalYy+eMrlD9fimoFys/56VW
jfBy+ZhYwaCtQceaB5u8rT7mxeSrVtzPiu8VqtE3IXIXrh9YF3x3KxvnwEEGhX/b
V5uIy1J4Fm7guhY1gEW2LeZUQ1YS2W7fn6RfAGkqDQMdCw2/x5O7eiyLaYiWtr8e
FwrJcFC0Gzn0kBju2kxNu4r/ZI1pjEBCZlJ2O4mD+D9uLltsNKegrP/gbiZMuwIG
lAAlRFPrpWeRzCVlU6qP4xQ0BFP4ecLAWYbQPbqQMHdxbTZ6kYaxlxkcp8P4RmwD
xtzsNbMnkZAWwT41LP+JoX9vOHQ4iPh2sBer2VbUtT4vqk+NliMU3U9By3VOUox7
PL4A3XxS6V5+Uz0pGqxLFHcSu+05KAH1PMuIYQk31JdDH5HZhilrxRwA7ZvJ1pU4
2zlgY17LLgkMYLFST9d9veRujlme52j0xyNHRK4koWnY66aDn98c0eHK43vUfTJ9
Q6zvxFC3vaQzd/51aiBNVHxVrvNxCUHHZxX3BQoZPzduxuqD604oQKACBhMb9aTV
zLeT07DNKgXmSUD5n5TfOY5Ke+o8c+bCNjW1MDHiFrdV2wkzNEETp0LK4utAxGAm
BrEg1tnuEuYLmUjifHX5HMttdr68gfSkB7y3EKKSI61VO6K4FSxLfQYfZNB3JRc/
DArrUeNqZR4h9De3jlgLR7QOo8d4d4bM+/6DF/tS2ssPQRQXR3ZjcxH1HDrgqRtj
qPPoaXvn7tN3hE/lD1wnsICR2Gax91ahJLBtq68YClmidjMZ1RtUl52SYfWrHH6T
/MCqnxDWqKyQsL6ejwuMyk8JIbYHdoFV5sTVQA89WAjlXBHsDPERghoiibS4Tr6b
PJM9VVsNP5JrxSvR7VeeKv5jSr9bxAKyFyJVC+Y3JNoL+patt91DYuQ+V9NE4xAm
akOvBEWVN1TJ2kyMZD/IFB5Kj3nW+01SiQvK1XH0xMFThqpTz8jnKmWSAVzm53Ad
uqElO7qR4Ronj54oQoVTe7m19oyF5o7Qn31oQXioejVyvld4tHMkhOKcP68V/3l8
L8QShCm3/riddlJdXFQGk+MelRmGE37SCkbJYlUCrCeiaSSbORIwynyqGjNw1FIW
dyYVPLbGwmnn3J6GJl7wWNerOQYGy38vvJYDBSGQoNpq2eyocxt+6oHXoaZ6b0C5
GfG3uijlCXXepxjeI7axRnsuXkbHjFMrtStp4Qe/+qn0b8wA0hnO4UYoNt83S0j/
0CBs4TCeKkho+hBwa9fKpdweF4FQa8RaVwLKPWj5AddQITJO3cILeF4WG/lz9yev
O6YH+BM0M1Sv7dFLGeDMkSZ100cAaaMpZn47D3UHQggJPtgi4vT99U7GGxgfeTN4
LpjAVuyuQ0kISAaAFrTR4Ru1Kk+vcTE5BSTnfTBoEhUz8+soqSQvMPSuEbyUZ2rS
udYAVNkOYPMCXiQ11ra1E4k/E+U2IRIl4HyuMIHxqMfarPvHx1U9+C6n7TLueVAR
GVt913eJ+IrQWkJdnII38HPP+p+WiBXsSFI3Vs2+WRU/mThDkDBueHLll7srmhjC
JWukDzgh/zy4IaYiL918Pf7SmJeWdMaL2TnuoazoZMyRPrEhGBakEavfl9n27kLb
bg6z7gCdSf5Bs5rwOAAMV+BmP64nR+9VlUH9V7w1UEeTIrfoJhQieY7yw0zdylFi
P8XXDWVTo0oq11zimwbrFr/8bX51rg1yG2Mdvb8jhlBHt2+d1v3K//327qZNCYbh
Zu4pdGFFP74pPpgd1m3IhYeJeA6ogN1VyV9+eUjbX7FHpbJ54qnFSeAKArQtChqd
ZKz48I7EBPVngDFxXlUpbFqMrL6Mo7LcJ2qEJWAhE0f4tQCJoLzYY/emijCxyzfp
AwxjsezxPYqe/Ap0K5inUqSNOWR53Eufz/i1DAc+gTA3fvQ6Uo+EXNzSZrXuRsCP
T91r1rFq87zQXfPXWseMpBeePvcJsgO9l/GtXDL+931g9kRkGF/lksAx7qnyQ5Lc
VJIIZmAnODtNQNAuZAneDnadQGvWDWHUk90C2ifPDfs9gB0CoKuxmEGuAWl5Rz/Q
OTLsWbxj0fGIkQzYocckryMK5zGq9mfVwqJ9NTuHycpI1tpA9G2u+YOOGIbG0m32
t7SdNCgmOJ3tNyT4e/srlv2O0SADu8X60bCDagOKP22/gQT26opEXch00SDXvd6p
kvJExCofTpXo6lOI1a8Dgc4pf4CsYpJQx4XBtbyh8rhbYiwHX7xJWVH0FmAgSbu7
BpzyfXGITP+Q5uT2l/iBD1aH7gNK6mzQTnkwYkJ2aC1iRhyUGF09ivbukoDLz7T2
B5y91J6ZJjmk1j7lDm91Ff8FmsOQNOg2eADbqSe5krmUEo/SusUctn9it6giagPK
UFew+y9Aw0XBbPWQmmVKnuOsWtT9UIZPiHYl1vuXiz7gT781ivYuCkNfuVEMuNjl
tpY3S7oXM+73Qa0RUXXcwJVnDFmUPN9pOzx2b4VBeWgMRH9dggoQsFJvcNHeppC0
NSYG9Lwqidrb4BWRXgaOxGJkr83fP76DMTsy9r44qDVqEhlx1vcYganNdmVb8GAy
cI8I8PuBCkU1cYs0aHVX9DD7fM/iOsu7mt+E+EAIDORoTuPXxJcJhbIPFOzBwi2v
WTmHHO4+uo5gOfN8lZg1w8hH5OKsg4KiUYMCai97uThGIDQbDZmg4BswBfJ/XFRR
Jd1s4sg3u++B0q6z5JC3+V/dHAF+rRB/UjEF2a2n3ecMcN7N/vF3uO7mGqv843vi
CZScHf5HgmtU+ardAl6zWqYRBDueddZ0AnTgdrWQIuFbfOEl7lfkQVlrMoQ4A7Ri
HSEnCG1iCJjFaBRQaznygkjv+7H0kT0zHjSZ90AEHC/z+KUHAAy7zwM/C5CZ/LPj
sHoSFTGwImlTVtYPSPVthG+lusEDK29iEP5PTq+Vt4Ja4l6Q11OvLNJLT3y89aPO
N/iMohRGQPL3eecWzIl80YUkvVIRZVLAckP7a446Fr2OXptFbyQzUag2WvCkEpcA
dHV47URQPEtlTCx02OeUn36s3sF4d0W2weGqEumtfgs2b6/zvQHhx3g3hg53O+U3
7ig5Yg4hFJS0VrrXIj6xKETjLgGD4b4376qYfcYEoot593vtN5GYY83pY1Pn+GcS
74GcSQX7GMNl4cXB+a7occgw70ZXyrDbmdcIPSEtNMxt+bZym2zlQCScfb4w1qC7
5flqJ26AP+s09XiVVJHgRb5/Qus+q7bpMwRYgtHwGI4mrLlbXvUq3mWozuc7TKCO
vUTRCMhoQz2eIJ+Yh/XXXSsGJ54a7gsocFPMFVsLUbAYVe9L+Psff99BDGHXIhur
BJwWGxEUJImBI82l3Qwyq1gQjWILZORzPCfFggIDSsbiMPRXZXyguFVAwrewh5LH
Fd76zJq9pmuQKHOVMUsjuKq0Np2NpEd7s7bDOln9gVpA7hTd7ig2zo1cOGlitmGJ
E5QI3fl/GUBvDabmlrg5lISzbvkvRUk1MM1Zzw20gPGVGRywaiNIF4tDaAIHGKVs
Ifm/WeJXOQQzAvJoRAKK4guurxCxsDm3xPtMr/S1VjB20ieiTjj+hOFedtNp+82E
r+fhRJ5CYHQohi32qBgI3ZgmkKYqiPD9OZzLWKv8tYy1BhvInwrwqlurPIwDhpFh
SJsgmDBIJIzfIuppKxYQzhqm+3ORGfmDfoImTJTCkkHp2j4GDxVZhFsf77QLyna6
hgF/9zrKq3oszdpyoVZL3YsDiAlbaSs4AAFDaNO3HVnyqSH5zLCP6cFoNM5jPkHh
FihXX//V4HJgf+v7p1KRvheR6bF1HnBEfZghnxlvGrUpqKxsD6rxINntiNYbn/yo
FAkVVQeyPRRsf3uwOibVBT54n4nyaV78C4Sn5GA+CKmeqF1CWJcmWqNdK0hDKfrK
YrrPLJhzRmWwdATrjG6VBQKCswtBu+kA/n2z2wv8F9ObAZk+HGkdzQ0u6wsCE+gr
rza5bc1TAB5nWyQffRadq66rHBZtikVGEMOcXWt+fAqJq8vvYD0q2j11CE34N7sC
08TAJeHp7LXcgwOWsyP8+jn9L+GN5RN8SzRV69+AwqFC9rv9gRMi10MiDPAfdI+b
JLPShVpZV+qVHSyxtAeUuyNtFCNTzyj9uFak2bf0GFZ9CCBmFFDAicM++Chf5J11
/loy4xc3WNxo5MFmP7Plm8173htPIDCYVJk2W/+VHBNSn/rGQuhXRap1rYXx8L+R
ZQCFW2rvjRZwe19a2xFMPGpRLM/eAMHykcGGsFk6QA+fLatqX6fEhkkelzwbFCco
5ZbMeF2ZjmwV8RACYhFgS86gzJ/t9jjtpPtXXS7Z5s1EW8YfCaRJvuPQJN55yVDX
vkVn1bkdMDK2X7mB7N7hnDu7s2xy2xb6y3/F2MYgna+xl26JHdrjdtDAyseoGFCM
/IA6NlgVgUswhqZFHxGIGaSSfTirQ1+0P7GPE8rluyfOl/JtLwVow9d4d/k6d1Im
qNBUYWpHzPXtmThS0MaTe5q6BMEyocqdjrVg9dza2YvlWapmjI8Ng36sprb0RqZv
qFlRJ4LkgthbyjZVhSfP2nKXwaptoIS+I/+rWR09+XPq/aoS/JckoDz9VmzVpdog
rYT+HDHM3mPvJ6iccSlMIIJfzpjDhGauUZm+n9uX83OIxD7McmJaLusv3KjdEWjx
2Qk4u7OE1Yd0X6DXbKpblspbs9ivrnrVgeBz5z2pCkp2uwhgMdPK5JyQMR7Evtd6
zDc9gqRyphUSE/Vmhht8bw/7gL9G1GKNW4+xSy9CLbeW37UrCtbyzM3iG0LdV18q
ScQMf7H72HabEo19kfrTwbPXzX9jdLfcmTFWeUskQV5G2yGBlcp4jkvZiMkC/1Nr
/0XsLo48AtgpWh1XoehA3TdvPKwNY2l84rE5B9AZcExt+hPIH5BdzttIBOH5NUW1
2EhjO4iJw018wXT6Khegm3KMBnlCZP8qP36c68ED+X48zoFlXUBHGnGE4Zl9+feJ
GoayvzsV2vfWCWawukdHH54MUH7XoNv2EBlXnaUChTlOP3dwBx7aL7nxmSJQbZK7
9ir2bW/NzdSOZLffzj4QUlEYQbWejG5gysuRvXPBfkZLZ63BjODcN8+QNaZLf/lm
Nh25IgRmX5H1crMUky6f+wztJ6Zr4SKtOEnmIlCy49wLSXqh42r2eB/VT+S2ZLLe
gRhMzI9ftArwyoeHPODb9iMdIwpYeGjnYDBE3C27F6aIqFDLw7a0NqBbR6ntCZk4
Gu7nuD9NKWfVFtaiHAEnQ+JLv68b5t1y4UJQ5MVj05S+GpAZ4MF09gbRCdqXkWgT
sjTxYmuVzsOLhRm2BgfRKIY9bz/e/5zE5NRVXXyQVE4d0uQ5xtrYEHSF81/kxv29
z8Q0J6hwe5SNZC7tj69Ef7Ij8+NL6bICsIOYuN69R/h5CN93Cp5kh9Pw6YouxgkT
yBz+mDEUgOydnJqwEC9Y3mLIULkyU/4H5bjOwvBNaqfhWyO1KRJqI+6Em3t2l6xb
ldndcO92Wf7hvmABg7lrkd/gi5oK8FOQ0QXo+DCiTxr1LExoqcoe88orIkhnd4V7
CwBX7fwF/nbWjYhHvCryYO4sMo55fo8k4RBSrwfgcyCBo8ac+AoRKzygZuinNGXt
tNVndx6Jwxy8mlLPl4tfw7Pk7lROgMWWEb2sAjkNIAfrUa48c47ySSfCXyIPosX5
j8gP2/NuKhgOrF6WkgUIaBXvJ5pZEsBLar2XMceF7e8nAP1IKuFIcx7XQYcOeWh1
pjEfMD2gACJSQAEb4Frgm6m9ShhdyKHImwGobS2r33WWHwcN0jgnRfRccCVfRh1v
hDXgC+zjbHkll0ESHgO6uSEbFk3NMUhWtHH4GQgrTSKxoMcdB6muQz8vt/wvtFC6
n0rjQJVqNwMXZSD4zlyInZkeLpbdG9CZSqy9PdVNqhXj/LhFCe1oN91BQGO4g4lu
+p4fyaGUi3i0PPCra9I8SpnwsNG7Xt1et7Z4nM3VGO5HEO9wTTnazjaQH4IMjgN5
KdZzY1tFHsEwL3Jpjoeryxm8S5jaq0FpSqljVyXE7sLruVqqowc0PXfXSb9tp9Z3
X7WpK29AAO8Phg2neWz/NPCOvdNicjTAzpJDwPXGMrfk5kN+HN9ky1dY8CoSUp5j
5KHfnf1vyEGB+ThF//XY2OUCgo3hA1SSc+kAKLYH/W5McYBY7CTz2GPsAkilYEf/
SpUv7usBU17E2lVVvW0e0jYgVN8HFVDLm2coHj9uLGPj+QOSy0jX5OBUDmnBpuXB
8lGZS5bxCCKyUu9yB1dRgGLREirReywE6GoEGIzSDn0KUV3Yy2rLILZmLkIimKAD
QJet8datiqa8h6eYnvYcvs27c6mVKLkxdCfOWt+gDn+xZDwnQ77Gp4DusRxMJGQE
mVSMhjfMWSyxYPY4ceUbBeDhqUfbJ4+yCgO4Cu7D+IEHu8l+JE1ZXhONZakpU6QX
zkV9fbhY5wstBF0oP1Vtj03uaTgKO0SVA5xHVmFP7m3wjdvfrAOnl8oH5IL8gFSp
RKNyOqXuEcro9QxdbXnj2//BtIjGu3OaEyqHfN4YdqFfdF13rp1MWZotWwcDs5mo
7TCn++CpgGN8zlk2TzAPLhsvTPHKgyF401IIeAgRjUNSodNP4zsbKf/5rFtXRPdn
QX+n/mYc287aSDS35xY+gFI80/CvQfnJaT4NtagfCl/lYBv+VgM0Q8PpNRuu62Ii
C/LjSi1pFsxGA/fWm0X2+Ye47eWftNXARzbTnICF94UMePxIO0ZasXNrZtJK1gQt
EIv3l8UK0gWNkhan8REuyQx2bTOhKjGWNo2b8OqKxvEnovtZqEuL6glo9dk0SrE3
qvTjw35v7aXVJPTagvkWf6dwkTnrZy7uZJhDNj2wmbX+P/LYLA/DD2MMhGxfyQP/
A3oG8m+VFEFbIxOttrJhKsP5TyMW//W20789B5aziE9PeXp7SFcchoRcckegoPZ5
vFy7Ou14Z+rsB5SRtCZtLcWrNQ/EFIwFX2NLaCI+Ru4qTYSnFbnZ8DwtjippeH6Q
rBpApLY4KECGvbtrUFGT/RJRhhH7TnBbHCDX4BFYYEB9XPekwbMGdBQWr7tstvzi
6ai1aRf1p+MU0Q+YyCKdNabzJiQ+C+u72H4jY/NOuXjDCqu11E6cWU9iNCQvS/Xt
59oyYocO024nG8znHapkKSgHUnb8ypXF7mUPT0TNuscnK8Wvq+hnQsd40saSKNRF
cVCkX0F5L2PEcliLNQTQXjAvIoYsIFA1IplIfj1QLNTmFRLNPkToYBodp6UtlmtF
KWXasWU3GsSQEEffGYzwc6KyQChoircNjgtLbqrKlp0lbGPCdMBKSgrvmV8Uvi3x
mvKXwDhhuqUVFaMudNtM78+bFwe5gUbtseSaBbd2iyljjSR6LSh5jfvL6XoOKDB8
slhyBWIi5VsYWoUgcwzmEqfyYZH5skENlt5l7huK3z1XV31h1S38pH/CNvmmYPKg
JiL7WNwUcyftaz2xhtA769Z24oPVG5iL//ajQctA/vk19k1XH/dTON3ZJf8jGf6j
io31FBrS2BmAsztKwoo3l6WVqd+8Y6vk+mzXYesnDqdr3uGZyR2AII2CMOYKn6Iq
vqXDQWe4VukbeWzeOCmDeY//dzMZq6OfEq84nRqUoopyo+uo0LpldPb6zHsgdTjr
kiNrSs9JCMg7Le5QFw3A4txcn9VpgIt33MFaOyS532YfAKdya9utarSqQpdKpRnT
h33dDJ/5aU7ma63OpF6GYbpG462zCA6LFcW+gKM4am9A2skncUHK1E042mG/m9xh
3UsztjUBzER50Kr6n1rgueR3tzSnthlniahTYaAJXLm78eJ9dx9OAdb5ekMpoojA
MErXb7zNDolnivhBj0lpJTfrekV4neCBMEaFjX0cIjO4KGIQUB4dG+1PRAoMf1px
mfBaSFUUUX4i62STmKx/qPevjdD9Ytapm+47Xa0dP0odfcLt4dBwPmhEXE/lie1H
FnlGrzuTn/xd64ocF+20B4xfc4b4WTgwksAsqJVn15AUuQVGhpmZKDQ+jp0z/4PT
DqkW1KcN/Gda/x97tXcG2wdeaN41vD4YWKeHvHesjyxk7iG2JU6bshoglVcP2vHx
RkrYvBtqH8G8f3XSuvusA//dhNTl7PZUbKQotTdyo51aPW/eRmjtOtT/UHm4zRnc
2e9aBkeuYh6zKCLOk/i8QSo3y2Koninwg0PUk92kRHZeBFhKG+1cwl19E5z9LEoV
eCLu1LYC2XAqkpreJKNCPGAB8vAV2WdbnrrLXnpNTM4Jr1SJkcHBTmaWS54jDULG
UuYLaB476RvR00W/Kr7Dvb1hMKaC1ZD6dJXYCczWNgBQwbrRNuvBJI8ylsD23JGD
FAjeRK0pqaPho3Ew7yG4GXpIFKQADdLCclSiDu9EBblD1TMQZnSlQ0XQKiWFcF5b
/D6IJV9l/UINcZFOZnlyEq7RW3oiWDAz346QF0T24Sk8TPIkiMmb8p8jsdaCwMzr
nxGgagQH/stw7N1FfhAJzXWshkD+LVSRzsurK/E9sdk6AOuwYdUH9UXdru2HcoIH
goAePr5vRXIKHwchwHiK90KZZD9Wj2CZyKpZ1xq6gVYmGXAU+gnp/KZkoA4tq8oi
PZlvjF4QmBYgStEqrRSnWzOzt4+RSletabrDm27QnXLg3mXXdidxmLf8GQr+tfTk
V1ZAwfSv0L5mUs30ynrtRjnaZRFrrhujtDvWtLgVNbI6uA7dJAQ1TejDj7WesnrE
shO88dAYdSEZ9iq7BFtjCrfRtrEt4XxEcSvPqadnOCSrxT4kbEuiKqwPUAXYfuQX
9bMU5b6C9MuHSNpdmQH11abB5rZDgBVnd5N1EQCGFo0mfdOulna+X+3x56I+rZvh
96KCxkQFFakLloaobAtdX2+WTesas7HYwG4lOOhVcIWaf3Z6i6UMpSN56pu0qktF
EVnV56QFDzjfU2MWRgdAgzaeubrkjp0N127BRNJagtFDnhBV/JLRdgfvE0b/ZKVI
k1UIi3QXUBV7K/agLZE57avMgvgLta5AAaNiNWXUukMPoEb3hWwyiwK4ovXOp2on
7qETEvevmOSM3sDaCYoajsfY6na1Kg+GlbqW2twFnA86Cd4MgmILxnEdFj+jXDLm
gtR89BaThBdrd2VPo4+vHrPKkW7U0Dd0Lp2oC3u5X9SN5Skl1AnWE/aXfo4apO2H
krybRQRql6E5I4g6aouOgMLK0F7N2vljiTWfSIuqJwHr3Ri7AWdnJ6LftI8XhQbu
/8WZDnZgZbyTBfmPuE7gbljcKMha/RSH0++ng1RxnsV9PUAhXNYRLfGPMkKvG985
EWj69SmvUQXEM1VBCGup19w60Z74/7xf4ypD89HwYKbHj0HT7q9ublEIvvHR+KPg
cROpEOuWQWxdDYRbHTFD53ADsOJHbp7Ms0zZixfBOv8olPWRh+gCHaBSmCsMk9aa
53gVYVKnhWFxb681Q9WiwV2hbFLpPQkdwS9486HsmXTzNHpL2RzIXVqKONbDsChh
rhNLC1abYaVK2zOupE4bvI6cb43KTAzBWaKthyHP+c8nlEPk/qLpDSSgXPi8LoyE
dncZgcJO6uA/B2BVLXhvpVhRXXLVOAF+ZAtDYGW7XpUL6QhX46ANJkTo9niCuYDD
gRHmRkizTMLTbjKCeJGIOPUwgbmSplN6xA3xWHoT4RuwqgUc+zje4Xae/t/lrOIy
r1Kyy6O0ifnH37WyUMWDpunWXjWlCMimSvAapFgaiQLzOTrr0DzZgFBX9ogrI4bD
4P04PlWI+eLaAvgque6A7VP9daA4uagNGzC2xao9u5LhL2+XnQIrJL48U+w3U1ai
FmVzH1+ZnljIcoDaLq9eBcaEzIcyPjC2iJ94NF2203PZ8dAEwB0zTncAL+K8FFUd
Y7UHVOA1wlBal9ko2hkWGUxmKf4HQTaJECvC+kSgmc+2abJ5znoTlzvCZSGraBp6
dFEOUMYlxd97ii5i/+aik5Cl41oJ3Z3O4I5xeFuTWL3NXgi7/RHLlYhs8DFj2s7d
H93ZvHdbrAIaLFEAEJKiQipCerEYPld0oHNLpDHpeTnuUgg69n0MjoEybUuyRSZB
R3nIbZCzfLhNALKyFAD5Dtbi9YmDVi334TLOxUXGc5XE/OQp1uPuTFFA7KtFXFaw
V2OzHIN6bdmjE0gVne6ylpB9f/kvof7rCuVkDuhEBMxdJQM81PZmFOIoybQJJWqs
MH484hTBy5Mgfafe6wuxRfjujz7AaHplpxU4hhIClN8CWg2yTIGe2Mnz2g3chKd1
6Zbse/NxUcFqypeSKbboHBAHEMXNH8+BaCC5nmlAkj2WXKb2BE4C7E0j9ONPaULY
lRSUtF2G8lI9lfWpTeTDz6aGzE0tbNaG7XNy61++kDqN8dSU4hDKodboEQYDpo5j
CrS+zEAhPH1sjN9pFA7hhYsLz94XU4VaTIQc/ur9B4eDxh87oa42wLwgw+bCthAB
CzME55UJjb/6d11RDWInA+FBvCgPg1F45eGbBRoOamPxV7W1ik7/ilSuD/5eORBa
TlUFJFx+jalwjoeLSlRdVdhNQehdrHFhmTRDzmpe9nk6urNpq0ANWeNFJ4+Us3Sz
E3EAhgVaPKajY/hoB0U7poMBPQ8nVoqhukKf3J3iG1fYQ0rghzWxgwzB6T9h8wom
7D/cweAqdpkpIo/rZGsdnaTxv1BX24Ab5Hp8cLjZqDTNJ8BH7JBCKRtyT86409QM
P6jQ+TF5Co12o8Cd4HLHCQoUJlSW4KHwWNsO43lhzWoouysB2GAYOO7qCzWuCmtI
SOwU0oX+6mOyb5m/Mmcl+11NEDgvy823l4DeiHatzcpOEfotMHIyC5BlPvka/Yqf
hsW46TNaDKf+IncVVDoSkGsHp7I0lwt7xrRMdjhGBqydeBzjDHr4Rvelsf9UUdZg
UYtIxvTPUkjsAgNAjDfdcAB15dYROKqSonhuYK5n6VYbfJBB1SjAPiqHL/pSk1yl
cuyxjkxT1IVst2s0uauI6DYEEefOoTHD0izxSaFIz0MJwv5gTRU6NRlvd9T8syjv
/6pk170Yjd6xqeV6MpVaHuO6fPiMFwOQ5L5yvoiSiwwaKwOzJqDqkO9vvbcDRfHP
6JeFVU9KFvXBvAaVd3Bj/4hNF/Pc/q6ApZbk8e6pY+lbkWioBDJM3cTo4NP1TQSG
6kmVLpJZVNm8dXu5BA/f2/5J+r4MrrE1UtkqW5nZxI/8baUM7KBbCd4nT8RT0Qrw
Wph2AnfZz8AhD8npo+mmdn1gCib86GsP99xJ3E74o2CoSM3J3UOGZeKvpX30pDVM
Bh5OTOsFJ1M4iTn3cwpBNwZ+riBnQxrvumH7nKkSW/RvPI2NFAGpOdI7bDngMAvb
oUL9Bwxd9hdIwFZrXrEomkBn3b73TOWC19l3UA+UBrJZjsR+YNgLubw448xORRhM
XPz28eWSdFjbjwfrf2kTJ1UgeJ59alSj1ZslUvll9IGa6Xh23H3SgId3EwDo492n
M7QzU9fH/K9kWwGQ+Lpo/oSnDsnnG/pnT0A87JbCa97w17so6dY2PVl2Jr0zf0It
4AQQ7VD2c14vmTdsxMxuUt1La47VAhLEPs60grrI1h5cMjfbA3Kc8ce5gG+NlaqZ
dNWrYx+vUv25WuH+BoG/xpc4lDLRo/d41m2iKoJMGuBTmNdWlbBDAtd0m375fM8f
YXuzbPH0i2A0DXEzTjaFrJ9D343kXgfae8W2vWjdVduBCSboDfqLhNImfMkqILed
u1oTxHBKgbIIsJwEKNfdDdka/QFQS+7NtD+DZALSaMkIDpFOIUzmDTfhQwRCF0dw
BWLbLPbMZTpdDHs2YmlZN3cFUHH3hqV2JPT6I/TwujOtTdB9E3X2otW14N0ecaVr
Ca5+U2IfFlqHw+a0V9fzijG2CNOCz/Z+34XI+t8ocUUwIwiJrfioSKnSp63Kc+JU
/YBKcNysTjKFPx+0M8iEqQRD953GUEJyPnpxhiTiQH5q/FgFQo7LJhOiYQqJe1qa
6JteA5Vy0ILmJeoy6TqDpgNxgXSWvHhhJk5ejptA80KZ3cNd2z5b2qjCPBdQhJJi
EI2q7GCTb0K6j9ghJz1PCik5dYqc1TMs5sAf/uNc+laqK4ir485/5REqkNFOb7xT
mHmd5XPF6liKu77P5aNi+bmQp3Z+7WBNjdG+fZNSl9ABdpBOUcSEeNNB+ot0q9BY
ef9mC/A6+xierkBeQompzjSoly5rWcOX4Fh5dbH6Lj9Uc0RGJ2OWcW0I8CGCpkBX
ztDgdrh5Cd5UmgZCvlypo6gCNbzeQCeU8s6mPhYBjjRcrNF8RxlG24oWRXBhLBxA
GhZkzOPpTiOAzz0aQQ4qNxDAmTxRDZ+350qlKk/oS1Uero8wjmpbUeYKQf5QxHc8
V/LPWUozGDdK6ePed67teYfJT64i62SpEPgZ+Z+TTEO68MFa+hQNkLeCIcB1m5F5
nrK3nMWCbC4G/XFp4RAEWhb8pcGUb6GZho5D+hlpLOEk1lprczewmpk0x23aL5Im
oIVNlSJuQPfUYhdX9NElp8O/MhFl8uEfFgvpiPGfm9eGvWVJTE6YDnQ8udQUh054
j5h9N9SYWH22Bh8iYA43EL4Ytz5CjZwhW/A98ggD51pd8e/n2Az9snKdd+7Uuoop
UXyczhmqXppLxdEHdED00RNgfWVF4ST2omHGeWmXkgNlSkB3g+pGzpYVKXHRRczb
KCNLqBCf+wwYk5lrJnqa64rPwUl8YwJZjMoaG+3OoQ9R+oGT/acu8lGgJZ5eTzGZ
rwNGjmqlNcUmVgK8cxSWFCV6/H9UE8dqIeLAO4a7hTt5FOoiUSG0fUHrMcbnPrwm
vsXhjvsONdwrU4vFSogKLKZe8jhuvur/Vwpfj7k7esU8DmGJC0on3hedoQwAQEwR
lwVVTrhPnzkQmcQfcgwgGuHyKfZr9FNcrOqIdP72cIekcG9YSJ0sBwtwCehYPb4v
QNejpnhP+1n+03liWiZ5Suo5sZtF5lE4wvzN7H+ZZW90HYwNiNlZwxUkb4+Q6GuH
Xpdv7ixtWb+AGwIJsYfA+IODY06elUB+xjE8Rq0srGf2AnEZNCldWjXi+IKNXe3h
BCSNb0Jb9PTgmsMpFB7lcHN/zknFc+hofJba4ypCYKB4AbHk9tx/ukfjkYaQVIfO
DbmDEj6Q5buZjUMrRfGBLbkGLX3jheYU9ethWZAG+/n8ibT45V01bdQeC18Rtr2J
mEoNNR9XwgbKiQXFr1J/EUpc88vpJAR4LHfUw7by0c5EfKhhoj+XeHPDRYhsiyMG
hipKNWCI6VRQTCs6BWypybiy04ue2/7u9/4yQoqNr8D+/Cr5dTXrsmhPNkA8rz+B
wV6+d/gkQ2E3gbHVXv5aMpfethJ2ZelfnPAtQ5CHEliuPdZsx9g1TBsGKuH76ibB
ftypCcjsRt8WbSwK25xOZUMJpcltZUSYd1lLv3l6+pbNNRX1dMUZhFAOvbtMKwm9
DJ2EIsYUbJcLaXihbUyzVdcFzRGMPpib6xDrPwRwuH+HafpGjAjVpnV2y4/XBEMJ
L2jZgi3D+meNti+2jjRXlrSG/OC6pbsoo+cV6KeZrkGgl8G8OMnpMmncv9UIgGuH
OnqZgSfPDZdYZmPtXK9H0zdEcxFE5OH73aICeKDGuiqDRFkYRZS36bHR5P0UW2nx
YcLjSssxIijMtfKForSL27W1AWCW8hI6SYe/dtwkNoRzX+iB048lUyUhju/Of9Fg
8xeEoHGck6Ck19CMlh53/7fzyF7p7PJ9CVPM8vuMhhePvVNzjwGKrFoD7ij3nbAG
HpNqJOt6hivf5lh3FuEkMBZB16oh+kJReDQ6Huu4m5d20AUBiS36lo1D+M8r5DqW
tGSGiGjBJZ752TldaR1ioOEZ+fBeXE0vQUd6dSu3+oSacVXkiE3jR1YVXWsACjt6
yu2Ho6nccBhJeelmYuBIftqELkN5fduwVBWHkFEL+Y8XskP9MUo3Xe5Y9iV4Z/DA
hRUbzVnHrHFTpCSc/UTuPeHuytfpjiGp2ecg4kiMGXnEd7iHQWW+6JU80QJR32eD
YB1rx0/S8PLJ5jyhx+aoPrxCGnloXGP6XxZz7TySVX/d7X8NJ1dJxIP6a2ckYsYZ
No/FE0JBdaFOJSCUeihScWpxMpzu7pVEZNIGLFwvbaxov3sikXTHkJkPLKCDQWo4
cMaIgrublvBZavfQLPZWvwHqIW/TiIjFw/Dbn3pMTcAXbWDCU1EBwcq79oMjOZgG
aAjE+x9sTv4Rrz9j1+Khm8FFxy4kFWyDByX8LJdX3LZ9rGeXa6XG+u+lF4q5j8FK
eWHsL4JNaQjsMDOGd3oT8FRHE+O1srDV5j+KK0+R8/GMg6I+otlgONjNfCxlla97
1SOEyOAVG+p5nM3dDo0InqedqnIRPvJq2vLjHdSWl6bT0QVGAez6WGiiv2+Ejp5h
U9nPZ8ovP6TrAVFghj95QoS/mulbZ4/aA9WHcQtaDh/m8ryA81JGx5abZoCSS6BC
koo4BK21sh3nGctG4zb3k85xEb4/9FE6lf5AcgFArRSb52opNUrzJgY6BNNmdCMQ
XB1d7v4ECgvG9+2fLmdBXdXrMrWvCVkpK5/dzQTfBV9lalv4VWK0/QP0AfSUBwj+
cW/HaJ5h3zY+9VnRD7rhM3H93LXbzka4Gp1O8EdEpLz34v5K/czpT8DLjpoHwOQG
Vw1TSrAWR6KxHIDA3wC5QO2xFdMA4xIkcVBLVuWlXeM2TIkVdBzth/NuQdlDDdNy
txd71Th4mPwH/RXf4BUfU1RC2enkmADN+Zwdnc9/uA0lF2dCSxX5spsOJ5X7XoJ7
4GxpCEie6bmpvRtDOzh8kSBbzZW99xkANWGsMWDfKxBOOLwj8flTp2i1WPiBewrs
FBpexEC5Xxht0K7UMKRoalSAU7omT+RyLwPqTvCZ816DtFLpsvIPNrV0xuq4lLLQ
0jzO2U712hH8gzPtpfWMMTE5Y06/OYo/mexzNoTG5AGPWiW/xq163ZExlJ7UdKyn
vMNooQaTkWMwEqei00tjAdf7AD/+lXOMo1UpGguGKy1Z0hw30mkuE1JBD+CHrYpI
M5MzEg/2Penv+MJ29E7UfFlai6t8n0zcCCAv6xmbpag8QtI296yfzLrI2TdQNSzh
N6ETj/yK22CLNtB8URGh3ZIb8yNlbYJdKceb5jMVmXZwu9y9E5AIuzjayAltTT4x
Mukv6/tBfTNMg7B0B9dsK4HPGXJmVf1AvKIQw6z+zaxRwGqzbYoa22FsDm1JhWT8
V2F/xdfH3he/R7YJVAokC2Q60mucMlgM4DcctxxIXN/gd794UkVWSKqaQ6seny9w
lwWyOFGkOQffRnlygvRGvoMB7QVuwwGrMlwZnVdGKgz2Nm32KwuOm+JNuo1elqRI
0WZd+ywj+Q2WDmU+fsqP0QydgrI8KGaHnVvlxMzs/dJSTgu1dAMKw7Ae5+Nb4ron
UBWghouw4y06QTWUyoq4mQxSeTqPqCdZrIp3Z54PVviZlWSBc6ax0WWFH1V2vOmT
qKT5FMS/o3+uaxNRCCQxnW9t4IO3A/UeoZU8I1ffp6mgAcagl7F3Zdvfb1qe/Ri8
2FRVsbBfZncCm9bhulfJJT0/5eTn2G9czg0XuwKRAPTohvmpjXdWchX5aKSZr0Uc
WPk7W2ItgE77MYrO6pOlXL5AAp+2hI2mA64Ib3SZ8BifEWolcSgnDU/cIgBn1aMB
/+2L0H1YvIQML8UTICbSh2pxCH4h/uuoPlz11bBzNmh5oR/kSGDJg3P8mYa2H3Fd
VipRPQWcH+RsdpsQknVABIrubnkb8vCFNdlsDrlixe4wruqIfV+8+qcrrRDZvXp8
lV+ix/onGs3fbebnRezyJhv4l3LCSqzOdgGH9G4iNLFYUgNocsRrfe6b+Z4pvsBX
H/+VcEM6q73GuRXoIIOpXZwJVgk0p2mflWPJg3rwLPW7g71frhI8R5WhCqUVgqNl
3OwJISD8h/4+T+9REIiWgNE1foVreJn6iLbb+MOnmd4IwH7IeWoAt005l+2sZh7O
s7tLwHI+U3vxfbG9umub2XT4rVV4UJj+v4hphrr/JaoOqjImvmfGTva7vNnxSVhU
TPWkDdV4NyEybd22hxAG2vWIkeJokkLl2SkqavcYkcxVMTivSNI83XTA0Sm2P8FW
XLKVqhXOjejokbLzi901k/BCGQbSa/CvCssSHM7BQqFPnc3hkB7VLPkWMgwt97vd
JSqGIeL2GdIWypZloH2A+w95kjGUeGC1Sq3mOhITr7Tx1Cmz/3YQebEWzxRFV77V
9oiqEGhPR8iZztYbD8U+ZWQSm9ypAxFOci625U8rGudu4GSw+IOvMyun3kcqvoOA
NP5ZSKAPF0uF/CpUCrKlIDmGvaBwybUJC4mnqvYqnkJV5ob59gtnAcOQXahUtbb6
XjH0OKi/A7YybUB6k+qr5LB2DUK708uzVfvMiaPCJI5l9ReMh+lo95H5p1cB0BkP
RJ7/vJwb4L5NiPRB96bpWZPogFQV/u1c/Pc9bnx9iXRXT44C+J22spCw0SUbtn1g
xlgwHdWoiM6+pE2NpylsXzu/l9QzNTGNmWn1eSmA/ukmFKptBwWL7wPaDCVgnNq4
qcN1qOVPnp/xnbAbFNTMBR9hduQyBPXxl/8EgCJRcJNI0aExqzPLJ4b1pjrdhYrE
Q1zNF0i9By+goRrbCoHYa2XimlCKGootRkE2canm6RIksaZ7TtOyqjS30X+xFRwi
hbEcbC5ht1rub8kYMzPHtiwxtTLwF0dj2pRW6lst+YAD/sS7m5dzW/AQVfnOcJXp
7d28DUO9w79B13fLaj1k1VP1sfI9OvhsBOZJ8i8Hw36hlQn9+j+EaX+q91/8NvFi
IfrKNNzberoHhjIu+G1fRQENfzGTpwULcweMFe0SiSiEUlHJc+zc2ne57LVa6MOv
H/jeY2bIHOiLOK9Or2h9f2tsenGGfgwxfg1R+5QVF9A2DVwu/qQgITyqTmEahQmI
8FLnDDhoA5L+LU4gI0M99QqwKB0o6kSGeSPAzVPXCnOgdRw1mrJlHL0r6XsLNs5e
Js9aIznoxSTuqrrow+98JfvSbhE3uSTl3HOrHCM6RmVULKNbZjTcTqWzQfiz+eHD
KeqvSgj7lTkv2q6bQ6xkqlshs5eC4uPLh3k/tK7smEkTA4ssbNRlV3gN4FMvCj3J
uaevjLvyScVyky74OuscnwMLddDqZU7Y2KhWlyBGf6rygdNVWoUHpVZ3P7oFEqi8
4uM0bDwkbPNi/VGQL6UWDuWVGOQmF1KECQs6IzvJ+mxELp87uHdntxKymeAeOt61
Dv1TTcMQ5W5J+fsPNwHWezFspO0PqnCT5z2ucLzj/mpUIXw3i4MOENO+OWg4uoeq
RdmJQKLYrzYtGTcxObYXPC2BQF5s+uw7vezBaLL+XJicPEC36VnrnEJ3GxAFHCCz
9feV4qZk54TYLzWKs9qKO8IQF3Ki1/vBEYrgFdwLnSO/Ym5B/qccYdHdCSFWigSL
Sx6cxgk85rqTrAlGCBu2B55ggcQyHAopwY2QDZPp271t7QgbSp6ODzLxeTRzVLpe
m9zxdWAyMJ8WaQPVOEhhdg8aQ9dtZQqZodHF5BtBjoph9wCCdeBWwflXrsRv9Cr0
1Oyd06J0vKW+RiEKlUUu664Xm1+hsUDGu8GSJLfbbrt4p7OWvmsGflZVEKPHx2u0
QaijLpAurcxWTB5u2W+N9YpwwQIuv5LC4LjfIfguBbyCwcRtZ67O3QwBDO/KSGSK
rUCovG2kqyN6BBrxEcrGH8/OGten3IY5Tv+ESSoIgEBm1pXAH6RTX2aDRMzEjGh3
jWJTRLMt8Mu0tWFxn1kKZz2+QjugQGPVK7S5ISz9+2Lx8h09wEp2PhDUEyij+xuv
a4RQEZr5jpfHCwreIKeHueT0Fao4eJyMA29up7BgrXLLKWqQIRy8yPGUQ516SSxN
lYmtveSX2FyNUH5wqU0rpAwV+5tH8ysTmJrGczTt9hIUFZQnOJSqNpTu2n6tWhlK
4ld7sF2v2qSg9u/dt28gN94DvK3RlpuL0vssSKW1mGOzZDFZSuZJQ4CPEOSHpsv+
jdBrxTn41QntHJR8c12xi+DW4Z6hMdL0oAk76RPXNfxMUkc/Cyt8Bnm7SbTzfQs/
ppZRAcNo+H+cCUxLbBY3+TIwTKnQzaUvFdGAZs/XvJ2vIQXBDMVT99mGZ8K8J5kr
830LRhAYalCeMBoeIoeYWH+Gx56YzfJoBIrHsyeL53vpHFurZlc8JVvuyNeSLqCv
lly97VakdCscwxdDj9mY0H2vzklHDMpAtFMy/5Ak/z3L5o7V1CFR9jPBm5DuzXBD
F6IZ+lvjb/B9rDEOJoBKDK9dZ6YR/oIw7XquqZJHnHVeQxqP2nzYTKwL18vyN2Nq
e+scEk89M1RYWzc4KH/dIjYSLR9YloBrTHtlDhG0g2ehqXBwOzOUgYD27fjgz8K/
O8MyophLS2cWTfhLa2WCKRS4RPwStHY1Jh+cJiOLg6DXDK+UfCQvwaTWC40KWauK
7SlqHz7KFrLQmD7k2aZupE+6ChedPr60V6hUiTDbNA5g/tqMZKp05EMOPsaPAHr3
bnvG1vJK08350WiQAE25I0DFAjQbN8ptNAawe/8q0zysFje4r8CL32vieVc6A9s1
7KgHLQ6YPyOc4h/O2NAuGHBSxUHgQKarwFNK/7mhDFkph4FrE2iUQKAiM5r8r7pi
2QSX0X0EufWw60nadD4fAVOVeTUCGe9wasI0dfHjWcu25aHX0Bo+mUsQeDAFZ6uo
CPV53R0voBhNj8duwGQuEiNKsgceryCCgeh7j5CAiDGl9u9w8+0EFmsovvMm/t+Y
5u7GfwdvAK4GS1MJDDSdMYsJj6Sz7fUM+VrFYd/pK9zQCIaONOLew7dI2DvlZf34
FzMXeT5zf20rNA2kuk0eyDLruRqrRXRQapZuWi1ERTiW8y6U2XDyE+kKHx+On8vg
aZ0w/GVzYbThLl+FNmrA9mQy6+Xme100+F7lmgPJW2+jwbDmAkkGrzu2Sq26uQAu
OMY5JpWO2rNw3WpPdTv71s1QALTVYHfMX7btwPzR6StPOzChPffne00kqZJ8+OWg
QDGK5fINAVlupyk0++cw1b3S60oiXyTnNiUvQdF3nbkeBtbnoqnnktSSJNGQHHfO
hmwevPGCAK/Y1wVPdr39YTfMPP+/6zMNw8aZHRBu5RMVBgJnQu127P2eQLwP3OSa
vdJJ8GZRcI5Y9saawxecNh/wjfX0XlJzr2SLRdrdREEDr8oPS+jcdXzAhexyH/8K
8dvOwti6MmxbV6iDmqP0noecvg/Cbphfa8wGzumPE3VDqrtsOKSwSH9EQHoTQU3e
aWLumrGBsDD+yfEREXBtr9GZ0fjGoR2uGeoubReDaMKrLTMvs+oQBQ4uJ22uVpbc
41D5Y1Eh/9BicWuYzms5G8yXDYrQwpI2wn14JeO65vnuJSQ4u1dp4aApilRvEn0T
fc7HHN3cjxOJ1TTSnDdU9UIe2vhApqkrDjtFSUGmUt5mmps0Y47t+dUcW/2piB9/
0ywLk8GMiTzVZ0ix1TmcKqlZNO/2pXYkBRQb2cuFFwaRhZ4Xn26LJtrFkE1md+bY
jboyNvECOSoJfkfWST3GZLjpd0L4L1qTBYYlLb8VWdBHQ64NQizXp5gIRC0VxbL+
iPwxZPapSTjLIHJ4LsK3Vb9yVBwjvRRShLjBfg5JxfB3bVpYpkC4QLNW1QiV4Gom
+x8DERe0zNg2jhi4eBG3878eNl69yFUGpKk8bDP3uColYDJZzF29iWUrSMuJ/Lgo
SRNUyNS8BN4D+W2cj0Y4PCzWsiNAHEtljM2mgLaRTN0EZrMJJ6KMlTTuFXuTdJYo
+ZWXbLxnKXc0YSSqp+xvkdQMBuEdYoNxfMKMO+/mJOA0DmnEx7FFbGZsRCqglH9x
BrvjvFK+GuW5i/puZmkEFMm4I7aO/QkQGL3tyyXw8QqAUIw8TsfMsUuF/pfdJ2cq
int8Y4MJrVQ/M5SQxQ3use8Jxv40YhxLi0sCd+O13ujJRrQyd246TIWsJJBrxAoc
ZZ/acvGzeWL2SU+s3w9dds7ys92QcDX66F6eoPaEMUQj1iivuj/aQgRxbF4ufMRs
O1btmDivSoqDp0UW4kKXfhnsiwP6h5Oh0lFV595gf4vzEL1RhJzR2clkqXpB1fZZ
bbwdvk6u0tSHWtNSm7WrpXW/YPUogeGczS549nUYyL4=
`pragma protect end_protected
