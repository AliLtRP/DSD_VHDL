// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lpZZ4thu5zjlMh1iD6Rql0beH1JQFzd11gBfibYlX4+BTBvwy2iGLq8wWHuucepJ
VKQDy/iUkQsY8mP9NUnPFCIcmU3ropkWB5Xm7pFEoktY9cBELGeExQpeLAaOLs2z
BfmeBwffTKjr6vJDj91ulkHk5lfCIGSyF76YMvGQnX0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5504)
Lcz/EBjSYwGc34NAWs1fTw+PepQCQVR5VajvFELEb+xER/0KOjXgagG6TxKzB9Eq
1awhxIiSM61DpK/bDbMMHWQA5es5gjZ63vIoLmAAf97z8P2t0GPb5f+u7zx2MQ0x
S26jgFSktStIj/4MurWINSSKPbUt1g0pnEPD4lrZug2T9QLk0Z3iR+A4vEevPheU
S+2ushGktPqNrwa0RDrXIyEUfm46c2ftXKJeoyk6qOkoTy+1wUFWkhL3Kfl+yUWq
aLcwujDFFBjpmVLX7mipMiL5SU+26fX/HKLx5g/V9x6K0HCZS6DzUT960vHmHFVv
Fa0vVmpCgPxZc94G5cDfIgqfx/5U/Y94rFpmCXiRktZsI+KPKRngnZg9VH1K+vCW
oGQqU+gX1/qoiHy8R+YkDKtsglOJmeebFtY94vOH09shcB3G02TwMfW3Tv87sRLy
2dGKo0m6bkOTCZCtSHo5xiD9Xo5rTbKQNEirKhkjAIKvDw9pk8LIRIjdmzhsaRcX
s5A3XEoIM/veAIxCePWGEx+vlMeFuFcVt518qLSwD2uaY4q3djZF+DbW43qLBgQh
Rfz2YieLP+vSQrlvW0vsqZ5M08YarBG54E4uk+GzKweg2WrAdweYJGcpVjFrcO5u
Ce9PxXrqtvJLJjRewI7RpKC3p7WcdRA/eU/+STVNyBS1ARY4f2zmLvUD7oK0ibuL
sKq7gdZRS1j1aY1s2ndsTugz3v0gFfLEUcSnYmnaVVZ75CatWqwhxZjukG39MVv+
LKZfE2auAWGQEyLwWUW1oN6cMT5PymSLtdOcToQCQOLk2AptYCpBwVeRjuWzOoja
0UGekO0UFT4ln5ZhC+dBI0bOxZ0BMsxtoqXRC5HAEgxqfB48k10TW1K97m4Z0mZA
YT9lnNIvfZDlHV0Uc5wKASLZ8lPugXUyp3Ind8LeVEfAvsHVA42VNFEWwSferwfk
ddCmhbCwEVuKG5ciT28SFNiopT03+XVCaJRJ+iJpSQSCNo3EvWLpN0/xB1rwse+w
73n0gM6aeBaV/I1/jtC0ef+4fAbLzeRncoKcX8O/V6tt601+qpH9/S1LPGAObOaM
oiI/fQCrMHCQu5GPAbQl9Iy90/xlIsbfMVNpMS2DBO3B5NfTdSbX8jLTwKSFgw/G
uhYGIE26v9ZDlLsipVWpj7Ng1fOGNETrSloashiAibL8toUNPEb7Bi9kmnc7wq3R
ZNHw4Rx6GrP9KhhrM7QZFjusYuZFM4OS+xD659zSV4amILczQkvczyTwPhSwSoDB
NziSPThuDWb/YAF+MmhonGiLouLbLvrrhtRLpPNiC7mLabgfl6g7blvuj9Hzg3Pb
sUkd4AADIfxBmw7xtnIpg8LIxhBNutB1c9wlX8l/wtkdKRtKvjY9zZ7XQFGShHCN
gWjpvOEeyfKLlIxS5XQH7jqNpG91c9Hjfa7eps616J0STt/kymWL7gBmvBnptPTg
HgJXVEtBSw7pUhC5AoF+RVz6e+usVkligz4qEYqgqfesQhX3s+17iUJPxLtiZqSe
VHh2TrouB4J65ClVjXWMqwPHsnakIl6WiRrAxG+db162wgvEFpOMKEkYYy1cpEJ1
+WqZ6r+EP9deH9Hw7RevrqZzCLl5SNG/EjQVZcMxhLC28QXSaoBDryhBCYEXBd4A
d3ZoVZe4URohzRRcbGjdzB3SF6yRqqoZhiAT2jT0G7vUxqvmUhMyeWE48aiNfaug
xraMNYPsCdPProSqkoZmqLH6gIulMeo4WBeEkUdTzX0FUexgaKiU+EsecxEpinrD
iCAMZFSy19SKu8HsW7p/RRGCLv3vIsPRW7qI0k+/Pi5J3c/NiDxI9Fp7wK2y56zl
3+NOZk4ZheLJXbnusU11YvyS+4IfBcEonErbf367H7PabUTnAH+oDKE8Jwy2y2+f
tvQtcq7tkuYxOqSHpN/8a0eXR9+Xb932/jnJ9JBpa6MklW9NlgxMJoBbNo6YsX8o
T0H7fdoBrMsGzVKxKuaUmPJ+nPCqS9WlycPVH3vzEVdytPJHiLIJtELMV5JCuN2r
Md1oe5DbyYlH0jf3LhHf2p+bC+rn+s8yx4fQ0UaLm6oo9womyqh5Inl8mJtBhf3J
WcYt9dsXMRZYxAzn+7BEL+EiYXDLWHtEpJEvRresn9eLduyAqjqzXQjSDM6QWzd8
0h6DZlzLYPPHD0N1Dta5YpISWeQTAJzNIuUuQB96fsuweTzCKRiMssNfAKQCMOpG
0yQQNdhxxM5Fy2BwcYK6YVmkTni49Vl6r84Y+nM9d3q+1SPeM4wAmhWbYyNfdm1m
eV6mdxvO1ZjzpQxponMGFP0maLqAwJNU2MOWtOJjW/0Ukc3NDditn+Ix9jAvdLxO
5JeLAP7h/ZkRveY4OsbOsZKNOTLy7QhzP9TBc3zvB2u3UsX4wI2MN+Zju/ZFB28R
C6ZIWe7IKc/j0ZWBWl5qROpTmp57Uk/WQu0QXGD7TG5vjXcdslLrAoUvfIU07Vxe
8aLwZWw2BwTsXb6lq1UR5phaIbOuJ/6ILXmFFO21cWx+aLgUUztVYaAO+FGtGdNu
T6lARYRvMy3kdagC2qXrOBzyfmOeC7uXUCfYejtxRE5eN0G+aw5zpwUjkD3mg3RM
Z/IlLQdjArRgZ1c7x/lz8mnGhMOr5HujBcwnXZfe4q3bA32wSjlIleUNBFaHiA3B
eemucF8sRxieam6UGM21egfMHoMztgHW3GUnmL3SijSnmI5PdL21jc1dxNQ2z8hL
Pbt4LwW+1D8x4PM1FYvbzwyMJD7sNOu9FrtNKoyNa5OR7gIbWuU2860FTrpzgvs5
oZMgqhVA1121V83diW7O54AraEB3+Aax5uEhvKxayCu8V4swQGAYa+XUa8Gu3NP/
dM7JfaJMTHI+JvIb9OZhE/5+OnLx5PFpOVcMk0G7XGDeosxJ10XMT+rIcFg6WkM1
vlGj85VfMOry28y1rh3bJiCTH7PqJT5ml87rsA11cyq9VDLir5U3X4daqdpTtlOc
sLB9kC0sMq33NC7LYSh0KDrusGUFfGUrtbwlaXCt581FdA40InmHyNzBluOrHcWH
5aOxJve+m20QWr7ZxjKUGD9u8zXgEEvUOZz40kbIFIOJMyA/PfhlVrgOn6dttk2r
rq8Cmd2fhouagvYZrw55PLM5j++wo4j6XbEmF6/BoAtTsrnS96cfcwYQ0ipTfMni
2Nq7TdwKzUUM6Cjp2oxAlQZVc6n/6sVZFaamPxfJAqRwnFEYBPPxxKtVX5IGnkNO
AFZS8RQkKKs3XWPugQRKhbtYvQTGz9iFF8Uq1ODCsm1OISR6wrHFSqcM2Jx1+KO3
SZR1dIXmZ7gXGQzeP1aYTw52/VI19Hc1zeI1SypfB7Q0NXvpPw33d84JsHSNkinc
++XwsIgg9ZOBtnoi1yEbONENW5LDMK4lPWVFI0wcGuzi4iKqufc2KLhF0LHhyEPi
BqVSrg+NTJ8ziHpP4V2UDOTbTf04c1RWemoW8juG9IeNaJP4rTfTL6pnYIgXzYK2
x/v+vVobo+riYgEDL9Hx+qyo9mtO6Oj/A8o8pFpyRqnnuVX/1l+VfUJMGqd9/uwO
GdmAMpPDSWRS7ZzinMK0+mIp34IoY6ew+5xWdNdZfp9JP0p7iAoANf68RjBeGK1D
hgReeug+KGMB+cgmhmeiGhq//nQZAHc+0+pvt7D4y3jto1nQFaG0XjQ4JZgi/u/+
mhNP/8+wQT9OdJHY+mUaQUPKKYYSm2wVHiHYHJpnECeEOKgSomCBrfUd7gtJhKMg
yobzowL8/BtMQMgwXIn30pN+By0zsOTsOYeNaZqFwFX0Gn/OEUfZkPx/4fsQMkH7
d5+YOkZ5Ps2S0e4b7kBiStxnO4bA7TNxysn3/DfKuO5JGQ/4sGtPHSSsXpVh+/X+
5ExjlDk9wxx/m/RwgmIg+DmVbsljY1olnKmKJm1OLWYL5rvniQW2RPoro+LsL9Lk
92TyWkSdaSsjUdHgmeGuD612qN/wfO92c1FSXvz2Ju+RdkJx2qvldZXf6Lan2Nkp
oDTqR/V94TdGq7jZC8JEIhf087df9Gfg95V4lNQ4D54s07ujxFcshXUHkDHYM85u
d967ToGTS2py1aPIfkNWjrnqky+Ghj/JLIcXpSGbCLmGMQqX1ZVZUR7eyGuIUO3g
UJAulkRxV52u2me5oVakPjkTUDAQ5oGYHG4E9x5X2SdtBEirsf/vATg8Tdbr4ty3
4bwUQ5126kO2+HrYa6yLSzZJyjnKlJ+J6iFJTmJfwN6thFZjYt5kdK2QFLerjRov
gxPdtvgvkkDvHt8gfQFp6ICxGMitxJT+aPtb8l95kIg6EJJ+mNkmU8XRKCb2KdF5
jx7StPBnaoxppXMjBLIXSqJdzVUDxZ+6FLnp5AOgM+bKx/+8wSTcVgN2p9pQ87Gk
xp6LeE6dGCXJm4Xd55J/Pfuj7+Hnwg++sE9VOt4Yi5iIPl0mjdNFMGoJGT1yxR4V
NKjMu8o4ZrWXFMYZlbODC6H+KgoXEgCmxVLjPvhyycetTgnp94z9AbEZTJHJoW1r
zxJ80REkzP0QxPETYS0KeWwfrQmIFelbi63CcGdVVNI8L11TfESaw1MzyERR6dCp
feZfyUbeOOp8NUihVTIgZFA7BPYVYd5XVd7N4IkSdNPa+Obrn0OwAq/P474A9tPy
z60KHSNocHhSaRivWTvW8awhz4X08bLJixSJ1C+GMPwOJ1eQf3u1Juuu7Vea9iRp
7UKP60ME6/uheVgCgtNV+u3u6rIz86LzISJfsR+wmiQc52eP/RcpTUn/6rjMwi8B
WUAXUoIgLdfmjwrVc7joTJd1FNBj4TUBuY5s3zU3XjfwCknPqv8QUsx23h2YoXf8
V3T29USUmqlgiz7i0j0dqyQ9p0Zra5XLSX8NUBruMLoWPac29g2iOJo/7b02D4Uo
GnbGSyIcuEezTuplJxZ8rlRMjBkCcUpA5fAlor5/TckpSXtnvyYbsatEaWNBUcaB
g9fAZZygKPN2tfNlIRlXQEf/3eeKBTq8105+PjHTbX0zMOETc9DUFhC0iu+77w2m
q2z+Au6YUO5lhqWSv5Vtl8ZDarHhBBAdU7ODnqJ+fuf4ppJCHNJ1m5u0AopvOMHP
jupdhLX3/kqgoon5ZiXomQLiUzZqOvx1LvbGhP/pYIU4IXvHrDm96KlnIkc5DaD1
gtE1MCy1dFiPsD15362NENeh+CFsRLHeYqzOHIqxgXlLOGcW24zIcIDCw1Pcevje
UWwM7Bm7Zd6SExZ/Aa9ddy3n0gWiH0TPCDl5Li0rXdOHQX8kbWypzLPbpb/kZkPj
jfBxH/hhvZM0Blqe/ibUf+mF/jYP83PduHwofVnhe6a09o0edH0Zk/Vw1am7INNk
WQ9N/o88ipSXDkFY9vl9kmuri1pNAmuM6rcaJ3cYmSisdI9FcTh89xzgs5g5Ea6w
/Hu9E3ieU3tWjpUm1MFKtWzZ59uimAcMa2P1r93MDmW2hFtQYSRRZIqLGmO8dmze
ds7ks4iQM/dqv6dyNMJo9vLHo/wIclWa7K2APQINPXolFnqjrnn2ivmz/1tp+TF2
fXnaMeO345aq1ul4ROCaBSQ0ur9UEXeOyd5qGRHaYCYywRc3GPkRz8ZBFiDOS9T3
79mZfzQqQRTCKOu6OvUhGDreJiIGbwVxtrTj8mSog/YIN1KdEiROtnFy+1egnIlU
uvEm8vbkZPYC7X10UxPKP/BhlF3d6pmMWyOr7O/M8321eNpucgU49nWx3/RhCMWa
ddM4hLDoBJbq/xJBR5pt66G/o4A8BsAyoKdF/CMBhYJksSM/h7CAl3Fu4TXhaAg8
82OQB4Kmbwg4CeelM45x7QIgBukQ+hNmqw9g4Xrcqky6inNBwjJXdZelMR9EI6Mz
EJbNC7v6Lq5JFBBd60e45Ga139uciWzJ6rLalrcfnuhf4nBtm4umIM3MibNHYy/T
NT2Un9KusQwweNm04DGsVj9+f8MGvOv5Wd8uNJ/IgUtFUIq1ylAwmytc7G0qonUX
IOvRlnYoTfU5iqKkc385DxWNSuu4EpSdYqnvLRC89lRnpz7ogO6yUq6Igk1j+88Z
PkXmbp+dqmqTzgzyIC29u7BH10apqAPBEgNIm5OKrhZ49+PbuZwkU7y3HvhedCQE
kt4Kf29Z7t5Jx1H52uWJmKODXd5rTB4KxySVii6A0fCJotq16GVQBIr0wN1mJkmV
GPEfX8PdBzzopgxWBy3Hhs1LlB6HPMyeYEX7u8IQJqHOjb4BAQ8v5MM25YgF9q3K
oRg6hlRTkFtuts0Hb2DjZaATYaQpn8tk8eypSwCgjclvcdqxT5tn9CgGXgDOPWbI
PqhDwS86DWPzC7w/6BPp+Ni1I7GcDEYxZvCx8UGG4Z0NOp0NEquSfZDAU2Ug2w7y
bhdKxZofpc3RlNlvUju4B8jip2aAITT0WEpFfa+4A2Sy2LaruAzVrnWlENgapr7c
k2QmCHQoGdDYhuY22F3aoRkVljChBrtIcJNx/M5w9H8kJl52AJ7ON0c+AYuSHdWo
VyACBFDtxYRI+LRiHxR5o3n4Cu3adbCs9Wno+mtVhqr1cBbbuzwj4nqGRtoAptBV
p4cq+8WeQTqlvp7YPu15u66GO+mJXZxRKH48pAy/JaYq3D1wMyOv/Y93X+vqzN0H
8HB18wj9hc3jWn7cCsjaAIIY+zsI0iX2Y0d76ENepP7CRx1nCZdumNR2PL9CFSoC
cHbeJff8M52rXwYKtbVXrN7ocoSZNczd9Gt09LkpUeGg+PLovltykzPlhup13jo9
N9WI0rCyMDL2hfZ8YZhgRqEL1HGHHxqizjPdZi/MQWj8QxprBFhmX3eckTMVD2na
Zp96ula9ZhIV6TN7wufuAN0ZHonxBHtj7RUkpvOPXl4zbliOdR9ZcV+/HZToBlWS
voh4J65kMYAeq9xZ2Yd1bu0OE84m0CnG2vlMB1Gyl3AyFu9y0YHwkIWrWsgW8l1K
evZbtV7fzAgYC0DKsQW12aJ6vx6w2zZE8foEBPdlCY3NsV8nSDeBzvyNzFln7ObD
GB7utKLtTVfnYEAOXDckiD8Pzl6dzdFTJ7zgzi+CZSIwYRiLyZX3cQAe/GiBjGo3
oRS8zdDcBBmh43xabrAzWepub2P/nYvigz6lMjWEyk0P/+J8jU7198bXZHTFkHAy
CSfR+lLWRYvlk4GEtSyqX5WxT/qXYcQZz8gEOX+sAxtwLEhwNGdbA78iMw0YjWcD
IVFAKNMIurBDiGh5RKKYtNXIBsxLeORXC1hBTFu+sYmePyTnmPhZKZZK6QTbavIV
V0NAh9O5zpt+yrMgDdTZkmkHbnLFNjCDQ6oEfaKvhEk=
`pragma protect end_protected
