// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
L7bkCxwMjxVXBgkYlso2N7bLXrWGO/3NrD5IhjoMeUAn4vUC6j4bgUIT6fW7FcYqezjABRNwQgXK
jz0vgBzQ28uZJHv9wijdiARewyyazVvz51rpvaiU6pD0DctNnsM43d/95ksPr+g3Fx/fXkPMPzC3
3e/X6fXHEiGe4/onMwQg+Q1W+9dbAkZREmUTUDo2KOoZTGXK0vNI8LXzhiFqUFvrelQt/ghSY73l
fV/ogRQmgOQ7Ow4nzP1qB7dcZ5j6vLAhABqN5MsdrbyQoMBEjg1TKktYknOjTO5HnTv1ww10t3ff
979etRafY8C6gw0V1OWid3/ZDYc6R54D42tk9g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
gv7wBlK2PHJ6+JEU+UmglGrTeQibuOl7pblu+wrnimRgviJPpkQw3Swbrru9loAZRGP5bgmgg00Z
onJz2Fq84D2kYbEV3AxC8I4HXHYlyt612WPMtLTlaRwODb1F/9SlyhkEKIdfY9bkXZ7JUp+ZEwnu
P2Cn06mwwnTGOFykcUMMvdAJLWXZzPgAKhb6y1WoNMkXoH8d3jDMsDvhRDG/Th43/eWp7irJa2iI
XJhWwIFbSL65zrbo0JTqpChZAE3xOilRxQSzw7sovBUq0UTJJUwEvWYRkNYCUdTwfnhgFl4lNC2A
BPRiY4REfXoEyrICWRKaVSiBUIOXVuI9pQL1Ds51iQskBcnAn7L9WZaZ72V2G4HBf/u87eozsjXo
VAbWOU25ShtRAWylCgDaMvwmz/Zk9qbrDba4x7vV4V7y7o2l2iwwnyOtEB3b9Lf4uo/6WcavXs7x
122jN7J3r0oJOst2kGWUdbODVpAaZ1BdC/4vIQFC3arNVzTCqL7hW6Dsy0TmDz8C4XlnDd0BIc9t
Bpvqecy6uYLLou6n6YJc9fT04z+jYLm2fVR44upsuULXaqEPVMWL+br4rcpkIVzbBCoOocN6w+0O
8L4k57NDmUb/KX57v5qOB3AU2PB816EwQotDWzrhrhwOyUfJoV+Ln5lckFZp42/7CWpD2LZ0cU8u
RTBF5H8inusx7z3/XpW5/O4u7JZAsPsupoDXTqpEpjr/AuKrW0fKTW/BFvgBgQwRZmcxY+WS9bwY
4VyDz+aGLo3eJXanslMPetEMckHdzgSG6IO7fxgMwgXxaXy2wv6tx/qcZFHMqC05klVrFFieaLLb
tQQpsJ/+SyLaeQMiJiCe18cdftV917jFuJQp0yKXtpRvY0SwStB08cunPNyTI9/xLdH7e6/q5MT4
ChO/QVYB5jvSx/ZO/EOFgM2tBK+Gy3Y0bM+DxPljrSOECzm/zIp9LZJhSuWCDNbr4Oytd01q2uld
B2/YyBpdXKenjI+nP51pi4wYqvAmd1QCooCpvizv6d8LSbAkHyFvI8up1HjFX+cWhYsUJxlGQckO
Em9cfsrnFRhMdLHSBCsR1AvxjfiEKOZAKosC+CMpDSttAgC+spkEBrQ8iL7X4snC/ZiJTP9bLJzC
K8BFTz9pvh6vpT2qd33PlTIPEC3BLa4BCF+1DkkNo04zbV6tdWDLymAAJCloDIn1imXvcXNFFVgW
xizLNSvVnYfVToWgvTUCgs7alQx7uNtwQLf6LcloILtwRdyXeIKKRR/pv/YcZ5VtZlmxNtwTpoR5
aZqsjd8FL648IPcekU8yLN6GvbFlJzEjoB/itkGUURpK4ULJ6DmW9369lluZG/viTloDw3AR29wg
epDxcpDkwTTFf+7FD0pnEZz5VR9P09okK71BQ7tlWS53lxKDsIasgiQ0Bi2qXv7OR5oDnlz8xrBP
2SUhIiJKLi6F1+YD+5gShIzItBZRlzDcwbwwJyXEOY+WjRN+yz6VzgCJfRxuTlapG1xC2REdirR9
7Un+R4xz1feJuVaL3cuDcLKXCe6rlBmUZ3/f7htez5FXSKuzPSCcFxBHygK27tvzo2YFdF2PjYJo
jLXcX8LShlqdPPZgYpTIXlLYa8pB2hwappIDiji+mum2m9kXDOiqrpWels1R5nqEnLsX5qlC3nMO
zUa13KCnUVo3NnKlm9mrhszfLPmqt0CViX4gZ2lTi6kPlKtMkRapqYGbjTgs6t+cQQtonYiS1RJo
CFzeDaL4QERk+kSExlcRJQaunNfPTmDca0wnlCksf0mlgGEJjyl4RorB3KvsOL5D+rc6JgSQUO7l
ST9fV/t/l/zWecO2bMY6AEp1q13qBdGlqLTj56Jt08ybMh5+5N6RqS5R60fmmnUK4j0PPP0zEE7j
iq2ooUdcPFtfM5mX/oOcE9uUdKsTeAg8+OjnM0atpJ7IEMCCuo3/XPjTcXQ9vrKVFHqsynzbv62g
zWjxT82zQpfAGDULuQW/++TesNQtsDUzkyPA25cgWdIsctlfvGIcSjY8ecW/2RGWc04jiYfZ5CK1
hlrLQmoUoH0Y25e3Shvy85aRqXY475GnIs7Zj4bkI3PssGzSeCED2sU7utx2v19Z+U0W2WOrnshR
TJgb2JRTycbn/f09CGn1EAxQ/2XVn+51u6zClm9dErctHWLU+tVS3OK2OQomPAAhLPizZA3ptKy5
ngE/OREsm+MGXr2Ss4UvKWsOUQIFQFwoILGSjH2mauUeJBCwOaUCDTYYR0/KZsh5pttPftWgBTOp
4C53GWWZ0m6QQsqkyBojzOUBp6rxS8iKdsuXa7KZt8S8zfUNPBTzcPi0qRW1fCzf2f5+a2ayMWEn
1gYWYa456PFCXAZsaiLPSotbmu3iNVsxBIRFNgBSvTvV8rW8OvE8uk1i/cxq+ea2bC23qP1LMkr0
NE/IVFuVBZjFVjN9u8Cv4dbl/v62z40OAW66ygTgB0Kkc5aoIHttyLUWHcP4SxlbWlSN00rbO+Me
Vi+nzMLIL6oLxO4dvAMpDJGNs5snGRqgmzWbU0rBatikztl2JoM5umNychf7nHabWriRwcrr8kdo
pbauZqYU6K4jSW5LM0AKoBCZ2RqGcbeK8tBU9mBg+7WNdIF8ApLp0ET8/Xj0KRo2hIRTbkNP86nr
R2ITXsFNIX/67TipGVGfEcddT9FstQFXxsiJaMeKc4HKgiJjfbUEtqnwoCQLIJzOm0005yFauqEo
he+MVj2dvqAsWm4AayCQ9fkZaZUv5I5HjJXcJBOdxF50AovH9laVRYqycODRVpN/iq10PSS4arah
YxvomKvapLJZ98fjRZFHLdWtvLORfQYvlVwJhZxlFOTD23/uHaYWR30bCkOau0t7ZqcAeNkQn5Yb
uDiBGDYAEIQ9U1VEkIZdFqL2JeNBlv1RD5pghGNXynBIROJgR0PEqALPec1HdLHElvtXIJMPKezB
qHE8+mHzr8QB7PdbwPItSMpqH+k30/2N+WHpeh0yo6uCoknXYrctCpw5eCLmV9ufDEehN4Vr/DRP
W9n6zi9PW9IpPQ6zss5wYccRNXV5cKttuial+4VwdLWdVfs+yIVaABGDFkLubfLLcypjGPpSpWpY
KO0kiUJAT6bU/M7v5cor9iTs3MuZrkJwOPXGiUH+ei7zIyBQnqsn8DqD1m1+3lg2wmbJ/2fvMPJQ
sDIPpEFjwKE0QBGAyRdrGX8soh2x2kWoLFlzEN4b5E7oiXY6YbqHhlJqcy+Teg9MieU74DbrpsHu
3FAqTADZLm+fZtW2Cvm5ojvKtDPXbVyawevIIZloYtO83t6MTu0qYxHfEpUjIWlQepQPqI6rR1PS
zEpoKuUdlkdsMTtBVBUk4LkKyi/CZE+Tx50wCzzdcWuCV+tfUe9ojjAar5nf1IcYnIXmxYX0yQUi
ZK3Ca3bQrdGTsYoBOATCPni+FKoB1cMX1P9R8rO8dCTMN9sK0Cg6LIk76QiMXy65p1e4X68ug9rR
ffn+1E/p4cVTqQbOOaX4BQEAxz/31jsntY0pYt439THZlnGkmZumd79ry0i5Mtp1kSdh3hiBHyKT
RjS0woCUScss72G/mSPGgCcddP1Gx8J2rWJ4YZZCnV0/q9JJXFoFClBShoZSCwPY3n+lh3eQReWn
ekN/5skZ+WS8ZyNbmqlGW8/bdRtp/RPE7O1zhjQ6r7vJA8S/31XR54KZHjvQBjZI3Dc0yX5DZIYl
U6PdqPM0++7b+2FqUCA25QilxcOU2jlCyarfkC5AvQhn7CZmFftbsAL8gOgjNnoLGaIGNdP8h+Kg
fSOuer/t7BoS1wUJuDHAtWzkFAV2d2+s/760rNo5EbCnnIhZiz74U36UDezLyoWc4sPfcBvS6LMa
2ReHMKnSNz3ljvpSpenQZFFp1AvqEHNNWTGb7kCUB2wQ472zbvb3ckJLjRWuAEWWITYMOCp4w5FC
V1aIs/5aweNs3VxuyUHZT3CaRiynyb/9UYHNy+2AhRK0qgxLxlIX3ts4efMOL+P/p1sD+peHt8xd
cmINIoHpoVo+l8DNMJVHwh0wKr8Tygn89laNWP3g4Tfpw9qU9qcetGUXj9QTxWXBjvw1I5JflhXw
sZVdJRv2Qgu5rgBArpvmfdHywH8ao9sHCdkBiBXsxnp+BeZK+vuHJwoN8E1YFa4e2x8vhwn+L22n
EU9R4JppYZnwlZ8vLd/G2w0SvnJZ69seW3o7RM1DdbTa92t7X/Zv2ZAjiNfgHNogovdlfERSAWNk
7HylYDeWqz/WWshZ0ZFmJ9x+3emUucK1LdQ6S8s6XVh02cd7eexQuUcWUfnf2QEUsqFSnluXERBF
A+BDfc4prhu7mNFr0L4Eh1TldwX37LWJQPltL1kY+p1kuAhVBseoItr1wAlWdoAD/BUR6FnPS00j
2vrX2LqdTIZDNOoB7G21QoMz1lpFKkW5T2iaNehlev0mR4vi3JyDL3wkzK5hNTRGYyRCogWPoXbE
v90gcBMv0LzQDTyxafZuYtnBhbK1gAM9yco6WHPER8Df/Uhugua/W2RqGss9ntcE+I+cmhF5eJvZ
DRTP/Kdw/EyurRiEN3/2+jVmND8yMk+SWOfaCUadERLEhdaw1hPCE8ILWZ2Jj+TW0Uzaum/hPDEO
q8X4wMcU9Mr9OKggnvcXUzGKEgo2Pl48eDy5dkmG0wKfyXStPow/72FJWChugDw/bXMqnl+KTKgK
CRVtZyGRN1q99xh4z0Q2iX/HDc+sC9KVEU5c+hYZWTxySzibPJx9f7Y1mTp0S2RzMDtTzGV++TX9
KphKHnGRe6Qw7ykl4yDfyLvEa0H9v/Zh4ADjrOFFJ5WSrvi4JnKEcznTpE+YDxQvEc6A8MOi8ivd
HLA+bj9XTcmldxbXc8/neoU5ToRV8FxNFS7ngtxWY4/9dxnyhLTZO2qthieixFUglqtcbcLk9Vuo
uI2ujsghp7XR0cFkfZ65KkqWj7YsZJuZ8MpdbU5fMc9mOjuGDDW106QUjkik6TvvETSiMk9/MjQl
VQskYjWXvJx+2GZjzH84hIyji/Uq/uyayRRR56gxDwjfQvZ94O7SRJ1SIkufzt5eCxOMpa6Vur4m
Ax4WO/C73KmRSGE8x1eo2M4Wx76UyVLxAXvCKnsfDX9xUNozKoB4volihPuQiGa5o2kCnxvwB7Ey
Z9dqp3aC9hoajEQjNIA6yYQ+K9BOGW2LoSNUlwk6kzi/X6nV3s7NuR5YzevSXb9ZBKVBzuVVI/31
cds6iM4TjYKIfbn1hUxWmIIYFVMB48t86cFD7Z2kNykHHzJIh2Omw2TNEza/pA5c4n1xRqMl0u+B
Pe+W48FXVYkQmn8RQzNMTgIU57MOwEasBaRC0d6Z6seBMfwCWjk0TZUXbK13VPHgo0jWIoMPYsIB
3UwjH2A6ssKoQKsYprKdc11jgq6HqiPorMQVk0atg+CAEVmmgqyhX4GCIxvDvBwaCoA9a+mKWZgl
jdUjx1Z4oVu1/2bSNC6+t7m5x8qMNR/S1GqUfqri6wizhxuOmbuhd5xQQ03ON3dqNDdFFRG4vYW2
6h94eOr/TY30Xg00LXUkk+SKCS1Otl/zmZkP+01/jsXvD5GL7bhODsq71jyyWAi/qve1MgjEoexc
vGmJl5M3BFFaAJ+ao30d2WK3oAa3/JCxGAgj2DUd/yxdB2PjNpsY6qraaauXQpn1FCVRUniqmZqz
zdFJL8/TXd8HBIwa+0K0RbFPinsebCGUM1zAQdc0m0dqqc1XMyrsDh4CsuZGubwH9txsKNTevbvp
R2lHwiQLP6+skqSkAmc38oX9Z4rHHC7SrAR6SdTjmDCinnwH/XW2uQQ3er1sFSQOexubpZmLjQOx
uEgokT6TjGV+pE9i2ud9bTxTdTrwi2TeY4Gj7tar8iE8TWLt9k33RrpWmPTjgc6IxzQ56Qfu1RyX
jgPZpYKMKNmjlo6IspehsMseIdM4jFIYMsNXXTaCwZM6PcYNJ7zhE/zhe3YVbJlMJiqxBD5pk6eV
wAu9Y5gembQtVqN3s3o6kof/LOXBbP0bIAtWvwHZ9+/kddDwiW2ybduIrVwWFIOtnO09xNruosko
u7XZpH6ypwTJU9g55Vij3VXPNDAYbIsLQKMku+HOBmhJbbPSamQMo0bNtgMR9wiUl++DOQDLwUDy
4DPrHS+EVE67J5tlGR9L7x7Hk7U/mfkgZhTpicTdJVtkWdK+h2FQ+8CdQDJuoGwr6Pp+Kh+LMjzt
KexOsuE2HvtZghDeadZocawChgnzj/ZArcw1ZSwc1WZDQVtM+yp4EdbmnJIF4cogMDCRtzb+RuKq
6M8Fu2kX8+NEIGq3zyh7LWkBb88CfCJMu8f5qhzRXrVgqKslhNB8NwYY34J/LY0VF956OPu3yCAu
lJ2mq9OFjLVaC5xmcHXd0uCOeXasU5pRSTbf8d1DklDxdGW00co2VzbPZRqBwewOfXPDAZj3IHev
HI1bBvdf9TG+tb38hE2CT2D/hWu5NPi2ik1VNB+2qPJJLtADRLyQqMlwkUiJ5Jx3ZCH9Vg/9sweg
DRRVIhqAFhYpf0q/BZ42f9HEpu5AC8+2cGYSWF1+jdbBzE6F9Mptr+LokauH0HyUuVVhhImrsmlI
KbZ/8SDnQcOOATs1PthkVE+ymuNfmHmmqzTktMKHr3DTxCrwHq59eEnwvNgJMtkfop/pECM/d8uK
ptHA/UOpl2gGv991cr+LoMqRl9cYpVrMyMzjGyJtYQkxMxsFas3DfRGfCxQpE8+/ANiABliw3dqm
vv6W03dmb9Jy+MR5CgbYfz9eId0ap3XpRo8SgX2/Z3cB/Mi42GcWC36eutMNO2r4SfQ5TO/VuPQN
ZW/M4cbKZQZkkRLIDS1HFq25uFMalE3LFEtkB2Xj/Eospmikd/qF8+yTGMYYzQMGFkRQgFRjuoa/
wNh7x4d2VZ8pATu3K/HWnjNjEDpuvZTSRA+WPmtymkglToml7WJW8kiDOA/8I+c/nyNK7CouupeC
4ltPH7kw+YHVzkzvT4BskAyz14qqh91ZP3EQ0TdTQmlCXWKwNSU869p11WtDqyLv3ef2705xSwwj
eAGXsP37T7aREpIpiAY1ec6vRubzCWt7DPo9CoiwPYvqPdQe5avFffLDU2TwetM3GeAmZlh9LjGd
orgyS/ejaOKDZvB+GLG9pnZsAHd0/s2rFS9PX/rjOlJ0k8WzjQk91ZtFKd4E7gV5osS6xkYsHw5m
czBeT7SZCQkfPTFRyU0n5tQxFeK+SDJVaSLKOXrINsR1CJQJ1oPbKdc5MrWPWErsNMPhKWCiMIwg
vutCP9c1XnOQdwp9r9kVTdhpUWgTCJnkHDeUCKofXN3QQsCGqfS5PUnM1BR8YrzySWZWoMj12IYw
O1q6ovf9cm7dBkVojERjnurpubG2MvEgwS7AULoRrMsCnYfsgJ1nOp/ZzCEeW770xpWFMYw/YBdD
INj7E+cjmdsXXwI1xuNf9+zmlABF9CzzSPBk0w5ImEpxchgzXFphlpAiiec5EFZIojWNE9FckbCl
PZYlI723kOi1FUxMa5zOVOXmU9m/RqU2URDITn3edssM2zfA8NWXYj0ZMtF2KvWb7kyErEsUv9KM
vH4Egb+y7SIV6Gq8P2a/7ThHwxh4p+bf3PSMyfFZ28DEPQQff7euzIBnzbX7GhMThcpAvh0T9cIV
sKw09J2FLQKiIY3UniHWqaREUqO8XiaBLgcF0OVVh1jN/1UMzjByL7paMGB7zaOO94mB+3H8bvsu
rAgmbCxCwV5r8SrIHkZjMi2nMSKOyEmulQnBmezOk3JHu2HbUJZrDPbORG6Eayu16PDYifTp6xGP
O0LtVrBImfvqf1Gnbf7+1Y08BwEZoQqqg7QuTWJUIw1Tzz6I2f3vX7mSE4q7VpKG4M8TLObEoS5t
+eMIigzufhF6Fu9jJlB/t4bnZ1x7+hFdcBtJbufNnT0mvEFkd43nyBrp9wcu+zMRJ1BCBDsVLhWK
bOIrcor8UV0tUqvBH4KDCJy7Y70dHPJ0mcU5QXmYi9a/GrixX09QDgRiKatUbNVTzBZ1vxenJEob
RaJ7ywJQhNaMLkJHuuH1BvyykA7Kqo3VGBa+GsGJngQ749Iql8IBobQ4zMpFd13IUSI49NJgH/aU
Al3aTO9SsmA0IhVF7BgMePJC5AYc6t66M4eSaAMEeqLA6dPvjyGEncjyoMS1MuCtvnwBtpKpsi35
Lx6WxpaG1z0tVIqda1IF0KnsExWK7jvRa+snZqPr4GXcVY0eO1/1djoPgoMGwm3vDNZcS4t4nvAz
wn14RQtAPNU2wLFrg0XShBy9/j3ZewZQ94lGqFItE5Z6RBBG4DamNJRi4rFVSlV42qmxqOc/sbMM
YefK0wxSTr8RpU/h4e58kCF+GVev2CYBuqk3oHHbz1K67Out+ZTxn4v1kC2GbnJYv8WiOrcf84DM
wDWg1K4QWR1Ig13Qt7zWGJxMtJSltw8UpGylDh4Fl4f1A9IqsjTXBZM5uTXHNcyLRcGhhCzmkmRd
TYnnN64CueIQCaYGfS490/SuiicBjAJKlK59o1PxRIut51/A7DH7xZ1Q77mlkakupOijrBeD1q0s
DqFZAwj4EOtWXrYwdT4wFxImXLSJVTi1JE9U8thhs4SOb2fN/ghuVYglUdTfnyGLe7UvpY04l4Z/
s/b2VCCNvJajEQ9O7iVJ5hb66lyi1ADgAd0huDOhRmFh5+oHH1SEDLNkiR2xjwY/mOnFoGQ1OFq9
XbzE5+wpIXPysXdn40HzqO02CECnalFbbSpIGc+wQ9spqY53gNDLmXb58A/K66jXJbG6O8AX2f6S
YM4DiOP5oMUdr9yG1wkaMkoRiuOA9BMk7xDep7rHmmj27w5vhsyWOGABSfOHWLm6ErNITgliHRV+
cqJb1ZG8BITnjOfP/7mSUQ9QiqFSfyYE1C0rKhvAo6YIRwUk9zG8nwgF/2ijPgmtJwmy5cbY/FxL
w9mt9zU/8wrSxYwdgNz+KbrFMBJjb7/zBbH/me9To2FZVdnq3SqOKNguxtraH5gyVYTbpbX97SUX
3+h6afeFtt3JLH7shP2hsLT2T6E20s4sssI+LWif9tQQsA0U7kt1u3YkM8I60yS0iZpXmykp+UyC
gv75AceKKWop80lvuItm+qC7VeeCi7dKeEN2Uu2ZtJRWgH1M/Gnp0COZ0H+2TdgpsAZQx2YNyVDU
+84NH+gj9Io06BmonzmfS6ylP47Gk/w0YWmfxpsc71440WHTF8g3uwvUT0LcA2MizrnKt335+c4M
ggNzOKpJaL1kcfw7w+CijCD11G8aanGxekAAvLiWCd0ZI/ckLvn/YAO4LBthUO8f5eYYZAx7Xy/h
Lc0cTFFrjMzGkVgLBJOZXCkRYFu4d5Jpe4l92+yKDhlrcpZnE8+i7I3LzSG/WgVaU8ix1Pl4r65M
pLmNaRBa/D9ruJ9o2SfZu39eA6IT8N9pFciOUJ0+ncQjAfBPN3IMOsWg/tyCjPb9T5pBH7QuWQzI
VjCOkGt/GhrQKZ1cBmeEAHETpig3JdB0jjdjJT2PcGF768RvHqmM3xwR9bednEUO1VY8S15rAVTk
zHhKFZTG3aQY4AuA9weSDkaYRSvs/GH0gCE2C617izjNmv09ul1r4klkVUqZPR6yk3vCHUtXzP2W
d/ZbyMRh8zIxbCxKhVbtvaAbJ8Z6CjKIByYLjb73VF9pVpeRjaS8XVUz+y8xGvTqGmB2qiECjriq
enZlnSqYkBwjUSFC7lH9kmiXjOrYPSnj546U6trkA2a0gQhoM3AndusMRkBTZ6iJ/1hraVI6Z2eH
lixuCMrMt7BVdsaQWA5rjSxVE2GHdcmp0+HLVk223K0tSTYZu/lpZpmoca9QN1PHDuAomv9lVJxB
1X8YtQq9WfHQqmj+GfI3UtwVdz53t70jcKOdUR3BrqqaqrpTw6B+DM150rsiZvb8Bi41ucrjFf/e
IAAoOjPuv01iN9SGW5vNmUv0nSloI27ItIIAYgGdteDgwuXiWRByelVttmkRZLDJCT8MWYdJgrwt
hYfUymid1j0+rBpEPc3EknHay79dfFh62uGoOd8cLwz2GIGuolS667hPxHSGBAjibP/CIDBIAAT1
9UWRSafDz/7wTNoCYfr0KvjmKhiFhuZODG+vR/pCl4I2zTRiM5JrLu+LXOdja2hIbAUMjfaOQPqx
ITHvvDHgHlQavcL3qnBzOjKJnEzfTqeeNfzUm7opUQPFKv/WPmC3NT9x32/F9+fcDCE718M4sTsM
mnWZLyM4+lashWNQKtIsBmFju4c7G7QRUNhGQZKpEg2MyX16ZG6JHLA+YZbwR4ejXxz/ZUpTseEG
KkVvVNcpRVH008DjWgHgAgMuMnHHT8KU/dDZ9sz3i1x/oUfuVjR5OT9vC1FgIJnn6iC1Go9E8juH
2GPXlbRmIjwydaAVUOxGIfeLZm29MNCLLnyP4JmBMWo+aoZNdD0va78FA5Ur1gWdeYlysKs/Xvpk
N3XYKhVHGCwD8pNFn1lI9xdil08kjCB9qKFe+mGUDLWXRrkHhAvjc3AnfZHFNnMFTcOpiwReo18i
o7XhqK06BWmT1t0k6PnpB9whkf9cK3mJZxZISqoB0h/HtiLF6SrkGGZhf6c7RybBSvlJsSHajI8A
OjHU40j+ukydTzbDb/Bmfh9ZvwPM+wOSWhN/jLRJMRPVahdT2oi0WQmgqYjDxWZCGAMHXNdY0cgj
XF4f3HMZsk3lWwCFslj/4UcIHxBnWgRbHc4DELg6/bTj8syRqR1AM+FN4BCSNYUaDIoZBg1r+muh
4F8RRY9hEnr5DsEe8WyYBkiTqbON7Ro6P53N3j7pWjlpBp2F0cpanfSYWSl5DfLshLvhZB9yWDal
XBLSE8ksDbqIN0OUc6K/pO/MerzM60gfbVgDHhBV7Q2u1LrI+t6klTOszB1NGDpY3fHD9D/jFXeX
Gqpfq5F1sQoWzoJxmBkYnXLbz8nwFG9FnGSeZrIV4vJ4VZE51nk3nO7+qxYJe2CDZTjn9Wxv6OFm
KMjGqOTY73GhQXLQqApsjPnY5jl46RnVHBcvIM/fh/3pCB6hCUQVhqyI4wBH+NdguehuAQ2K1Fxi
Cw0P80Z74wf1GhehSH3dwF/7VK167Ei/Zywrf4yYgXhB6YWzw+pwJayiNQrdjVduKhTlZSJDuLsy
QjFkSczzPUI/IsRyL6PymLiJ9Xf97HcrgwztNTnU+GKH3veUj7zl25/xH8AGqg0xYAyjdh2K5ZpI
LsJDF2YW7Yi6W843GsxiJ3A+vmULw0cONAOHftGJ6no0JHxc3C2B8shzOyrsaHU0rRhcVLEo9Nzr
dEG0S8h8amjkXO6MMFwpXRtkn3PfOUhrPSnwRA3v3UZX3Nmv+cSFwfJmeNzABTszD054JdDViuWe
fNSy1hhZ0uRhPVPdBZdFdY+DwofvtvLO7vXRLAkxGF0k8RiWSY8D8YoEHy9Vd5pRwcsdy7raQL/h
qlayhXsea2ZxeTLwLs5L7kS/ql02KarYYuJ5kUVgIYNKsitCAUG+EwfT5uWaXykRNB9KOcIiSOH0
qpw1nB45F2aK7KPxB8Xn7Ua95INODp2jJVi5RWw3/m4isHFRvkKYdqT70TUsgMehqfseyZKjmCS2
HiUO3REhYwY1yWCLCimyd7uVtIt1hGS1WN5jzwuWSQnltM6Xs7PbxLV/8+YtvPbckaRvSH6iUg+U
e0Pe0TsXKbOxeWDMBL8fqCFxuR3csoCTmk3dDa4769hmw+Pn42PBlINlrw2iqmiYpt5A6k4YV0Wj
2BsUXNF1ab0I5VagozeRpTM1xfybpABeKNeKOhj02cVkLZerI8zn1Hv+rURWF0t3FiujmKdpCxYI
0O7/hVbdvw+Mqu1eflq81y3jc9euOMgaPJLpOrJtiRt0IK/VsAOEG4VQw/7QJg1TEW8NjAk99u7s
suAsTmfgdxVGdKHUAwSrWvANwMV0j4tkSeREbVMu2SB0iOkMIrv+Hib7E27dROhRdfo1zTghZ6Md
HNjg2OvbmwYMAz1fumYobc2RZCG+VTWRTXkvgZiVHgS6nWvLVg3OCHYQksyxwBfBb3QGuT/QAcHc
PoqXtkgK2WAUslIREQeqhz7KBLp6U1B1M9NQA3Z8D+5vqXp8hRVbwEo4o2wk0SEA5c0vBfNV7WAB
XJqhFrQeLym9/ln6sutZs3tJuECpWMMEAj+7UAUf5ZR/N8RJ3GxLVwWQ4ZqkoTvLLdH/dXNlgkmB
L+cO3xRYysJVknsETP5Zsl+1s6xbfJz4/DCIjqbpsCBwoJhOoZBYCQZ50GWST/eb8OIu4Kd82E6+
ClCvgD0euvJ6m03BXoR6FEUI1zS3G/aDN81ckTHxzBD8bqvfK0cWLhZzA99wOpwNolcX4mNk/drk
T/zRR7O9xKF9Y/loxnSS8Vm0jGitrcTzmG8qcRKAJh3jz2zDj5xE4lDt178rO+coymrrUe/KT3ZY
+D+28ClFlpl5AyQrHSzwVuOU0H1DNtwGNs/Fp+xEifUXiCZN3OvkXqadMiYBvRiewsULZCGTc2hu
OK2Jiu/Nz2m8KMKQVIkqolk9F3MlI5aeuJxDtuyt8NgrXmtcqgLXct3wL4r08imkGbj2RYhVPPmV
mSEDV+g9rcjn62lIB/H61fZ64F1rQ90RZlrW3DycFrSa8yJMEreX7pJOFqLpITqpk/0tJWBahDB2
DN6nhX2j/1pqotR31bCPRyZIWUP8+IlUQ4egDvdzxHaT6URnLzm3tda2fVcvo9eCZM70xr52C6t+
wlJGukT7Ks1UQUK2gvvkil7NSZMLafSOoN4U9wGECrQfQU/Ig/rdnLyx164ApjyJQG97Zi7F5Lye
6VuVljlXgtsRyL7FwBKHIKQOWqeqNjWL+X7IxOzU2bdN5/A04acmxZH/MkEHVq2DMZF7agsRhp2C
VKqL+hZLhUVVKJcumY3ND+2Xxs3GvJaYvDGmo5VTZ5F8umd5TFVS7zqvCqjMk2UIT7wCbj9cXgDR
tqP7iGSdI+efiWjZlGCj7Foe/6JZYJUgvBMnxKHZqd5CAE2+lL/Akr6THLZEzPLt/5NBNj+ay4jR
Bfkg9U60Cn/prLLz8zW2mfbpHymiiwFcj+850o56oqr4F1lEZvVdbmNDoL9JFjq3KTc8e/WumADJ
i+o/9J+k3TbMrUe5jJOgSdmU0GcewQ3Zdj0SlFQSX1qtfKtSV2BuQhiqUFVDMt+Vag4F+JMEGujA
avs48No6/Mkk5yayh0zOLfIUkg4r42KISzKDQ+0yZKyzFC4HQeZNFMxjlNIyqQlu33ZTmzZ68AIl
vWLy7C20pzAaMz32VfEShmA2SXQ4Z1IZx+1OgqwmZN1KaTjSt/SOh42kLWrFrwy0p8y1M+0rFfSn
6idIR25Td9kxY2DeCpRhkyaLctmPVc3W3QejlAPWf49wkBq/RbFtQX04Z++cphVE7k3X9Bd0AmR7
x4BmlCGsTzaBpUe++5cflbR2AkZ7P3UvMu3BC4KUOdu3bEkFqAgtmQruOQmoEQu6N9be9Mgjcr+Z
sjqmKPBPeZsWHz/VELTizalKQixUaoLU5RKXgIcy1OV4Vu3xGGOGtWz+jEZ+Cm7u/od1C59AdV/I
n3ZkIK/mdn6ZmrMcnyvctsCFV0qxCZ+KvfCxaGY9/ccMzFPAU1UWjSdDjupY8t2jzN2DRdmOT5ko
mrbuOxRb6q3vpzzhFrum7xCuFNtyN3e5+1ukpJ9WbC4O8e489BzSISHhXNi0vWiOM03NBNbUBKa+
Z2uz+EPKI+jNGHuRtH3Uc2KXOW27UP/w+ZpxML1yH/7PK96lMHyBJtmFir4poTXqBjCvQd47/oqx
vgHCOtHfP79EBPyLESYTqigaB8a4JPu84Q3nHbawUkbNB3aKRs5VU7hX0k0dmlrgyZpmSAm9bkJV
NkdgqWYMi+k7gydjn0jsDCVTUl4WXGP0nWIvQlBwJW9+SoewHEbabusmZ/50oeDdAlU7OQAc3OiT
MJMJBo+isEumYNAJdCHCBOBRKCt08gTR1GMZjKgIJBsi8s6sKEeJLCH9tFu4GabcnSv/SlwDagkm
+IbjrxA/YSVbIDQmpziFbArWQzmmTXGuXt4fw1KbGnkLVJT27h6iorKQZnuA2O79hDsi9R1ECitj
09y82sSMJc3QoOkiKvHHiD6h4Y++mlRwnP7agAFL8YJGQ8s5o++lmksbHMYde6pcZajohy6ust75
9vSQxRP83bgUYU5s5Ks6TrMdFnDgeklIzMnbIC8SsRe5Tlkt47P0+SmkXc4605RZrXZ49kvCpZRc
SMAxfKTAC4ZnxoJ9dDH8w0rK33ALwKk1Xkdx4aAYjIyNSQizZ9f1Spv2KfdNhox//u81qV/EmV6M
V0wvQg4PJwB4QaE4llI2vxOpH3rGN6YvgPZ3ll1sSF0fvXYQX2jLeOFkF1djNyVPUZQjVjIZ2UQC
WsAALdyOBUzYhrx5PYUH+fV6IgpFdoZ6v04PkzVuheWKmuBQtfjA6uUd9z9+HiCgFIOgTVbvITbO
RgLl9mt+3RU/Vcn2wYsUzfd9N/lPIdf2+BP5sZgZTjMrvrZBaUTkYdFXtXcNCim/cL3WeHJxXddq
3MEX7wiOXrGXBDPLirlCZSjzX348wCqOXnhGu93awcVskIY0TzNaooxyK5HdSGgK+B7vE+Fdxq9p
/jVs9HdLMwSdAx886AKDKalY4deK+hOv2Azs14XKB3EIWcQ18B+hmBmKsXDqctZ4UwQYD0R4XWy6
lKNy7nP6N5rwdTvwCeyDyWgdHdzS4Z+/WfRNFqv0NDISvrPMfHgNURFg17dIPKAc0NPlsHkaVihZ
0ECtlCdNnAG5sAZQ5DXB9Xd4kKtRmie8g1ExbVGPSyyYdE+H33uLD1cX3LRmyHfNMVnd/B47Wu4Y
MJfhcZEkKWuwiYO4S9h25l0MzMC1QFZ1tmJn1mDsTkBgHyieBfDj7q53NWkC2iVHmkeJiN6gtw2A
0S4BHhkj51miojV96iUUyhgDkvM5P3YJqy/lbUaagPnl062CX5xy1/7ix9aQhKyO1VT6rqVyawG8
+faf6tWpCf7uYUD7hN6x78P4v6VkgZOi41DdWdFz77JWPSQzejpwhGeXWHcplbLYEU9ReoomwrWZ
X5XEiAW4VJ9RcULZL4jFs7iokze+IayfHe66Tgf5bl4TgeHpw/rHj35lW/KrB+E/vdVaA+qsIU97
MtbWZjnfu994iwKpSXgdVjD+S+XSf1ScdXuKhGODRqWBZd67iApNkE0+m3B7Akg+01L5IqH2gLJk
Ug5h77t/tjXy+8iASco1rQlSord1APKIljCfSh0HtVERP8RwrqmebWz6/VTgW86o565EliQL/F5I
yesyYgl2En6lBYLMgXo9mGY6TsBddkPI7yjUtVn1iFCA7+nJ600A5xCjONrwLeDu6bGG2TXM6ryD
Np25GreK3Pz2IZIsaUMlVMYAwonnIxgA35Xi6y9E5SzcN14VFbGcPOp0zf3vii6VM5JL6s277bRR
KX4qVxrj/sOJpY5O4bDdK5sSJZbv09il29WnqeDrkwDUtX5wYAS75NLK+DB9g3zjafk85pZxoUBD
QQQUrp6aVBXAem/n28pIEJMD9TOGlR1TbxUMseMikYt11KPuIxHfwTxYuzYUlY1GJH1JHtTPMJO1
lZE2PtbEEgWDXUIFyOYFBkScW6HYnYJVtpRPV5y5sAbK6jpCSrS0JhuH1Cl5jVPdjA6rYm62Lvlo
HIJw9pxzBjRGirGAFGAfMJvmu5WTpjfZzhlbXp7vWupvPAhWGp5QbjHla/B+F/FlfICq1/f8rdaV
`pragma protect end_protected
