// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:06 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rp7G1gua8ddafWthmbDGcW3Ndt+hn4ak31HLZvLYF7BvGC3ie9Rz1mUSxOWc3VtR
8hwDZD7kfXrFH50Eg4BiDr/TwoRqQsrMZDy03AbehOBCNmarH3YlxvG4NayV4yU6
1DDbOGWnkMAgl3AIqxbKaMrvpNl/PLUZ7cid687p7wY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20992)
wrP9LtNKxHC/OpHEHRrkzWjpljEE1of8HxZjfjv4vgY4Bl15073U0vxuZAh3NsOy
123wMFiZEkU6EK2xeJyTYX0GkV9Q0/7daKvQmVAQr8+yhdNi8RMtFQgZDHCe6Dwj
KUoqqMKgqCunFiyMDWWvCaGlxzQi5QCPJ5xD53KphSm0lNCtRLexJgWrOSGkpu9G
ZPpFfFREIDrboeh1m1uQ2cEhSS36V1HFZ+5ayPjdXrJX6JwuPUaZQL6GMhdnPMMm
2vAZaBpGaNW5uqyeC6ruw/1eqMZFNiyk9SKVmjeAlzBTyTxu73QaF1farkPIcxG5
YtLe+H9g4W7aYuw8RK3l7+XUg+WRYmhQ1fD1JpUZG6n90ZrAXXh364TZIdknJWiO
tu+j8/67gUBOiA734ZHK0QhUDmaVGbckaSqXXo/IbsV8RE2W7qjxtqipR9/yWCjl
tALbcmVhcZwFQtSk0sNBJm7lllMrSk5DIKIqb+0+cv10L73Kzo/PtEekcXCEd+Dg
l4hK2cma8+QRxp83v9MDkhaz0fpv6+rHHB4SFy55czLL07zrzKLePeVgqG1v/n7b
S8ON4WzU2vgf0ZaAR2UPvKZXYiX1+rhu54L7kXZJlEqhIEIrtDQzFWzjrkJGSaFj
ejLH2iwr5t851DmuMwbLND0IO+AY0d5B1Ozwak8m3pOU4YJMZEFgOJ3gcOca2x0E
bB+omjsTqkpAhR3sA3Ts1aZDCX+xIVQXIj+KXrdiZuHKSKSgmXThxBVuUJMkXTC/
A5HsTwrAcv5U4gOJlQQZrbWE/S0U8WnFI+E19DiQvkodoz7fTgmxp6dQsh3/ymFU
TrBXvSY7GlFh5y3vXU4jJ+14+qjNa5Q2V1q176r3CmrF5KgdNZYfw+y2c26Nb37k
T0EOt3OpA+JdgIVWKvtbld7S88+O+DTbXsbu2w/l5iTs4Bfa8KuVeLWpR+x4Azru
v9AMN5N19+GASSWuwwkQudggfEZtXDwp8fJDHcfpJ1C7EzIFO6xBzlE5Od1Tc8c1
/t0b4gZGLKLcSdTrQ302uXmJDvMXggWOzlNEZfpinLz852nHuIl2UzGhpT1Qa1AP
lWK4QpiPc2G7c9o+GvZGemweCLdBI/TvBgVggj5cryfh46GX5zu2qLiO7BNkF5b/
5HDBw/sRKZ+cWWby8u2Nk3wyvoUgScMvEe1pkQIk78oYUbGTuaHV3RD+/YnMkSrG
VTGlXULNKQIa9i26NdLOS+OQc+MWwrnh1l+Nr151I8Z4ffXpebj58fqqs5XUsP6s
PbDhGQXtmved5U/Ofr73XZCjF4+Shcasyq5mZaDmoYas5psDbFL+jzpyzp56uFXn
5GX7Gchf3HmVUE7ofT48PRHmgdA+WxR0kBh4HifSwgpHPzuP1Y8HKwy41SDVDw84
mgSCkDL3oE7Z429Qn9+mcwfH5MEXYuba/Nfoh/zKQJj1Ra8CJA2gsf86hm4o+9Mo
GePFZp+OHhNZUXHUNRd4W+0+TTHnG75vC+j5kULiSYrfIbLMg62BT5JM6qe5LL4F
nbCUY2rol8ACxJWSXb85WTPdSyZr0QUUDMXea2CFgi0nQD8ZGMws48ls632IBhNK
qAtHTsRFHxga8up5UVuu787IsgkzoQGzJrwWcpBy/rXOfepihw1cvKz6CSgvpDuS
H3Ixf/DcrIz7+iXHFCqK8xkG7R9ztdRGRdalbd/TyPYaAMAFocHXHfDGmOPa9pJN
L7E7UIsX5Mw12TolbjimIcoBeYZUOlnEfrWDVjfY55o0lDKOwKkpSlwFUkEcWOgQ
uOOBUQyB8WEri3vrs8ZBBKOh67TDXu07QzKi9eboCqbwvZ1XSZ0TLWQ73ndql7u6
VjhDcYHcdbLx00QvxZjIqmrKGN8D/IkYxMcHaiy9kkt0owUBIuFUd9ByrJM5WYgc
61qX9KmLuNGmIE6czSMS1JESqVhLsqZF9PghTgtfTQlJaYQYBi+bKMcXKdS8hEB+
7DTmAVixSYI2V2HembMFxpQgUFhCJ/9VWsDDru4xadq3qXVkLQXx5vM93Q2HddSv
6eVFcy+zI3EMVssSaoo+Uqq5oDPgoyuRefG0N4rbAXx4VSBNfjVrw1E6YhKNWCZr
Zp/d3+v3u/xw/n2jElE39W68zh3cjMrVM8z6PRsONRoh5zBfwnhu84I0lq568V88
g5GFj42S0u7GN3xEvkH3vZhtF4ZKM/ruLl7rDtt1TZ8E86xh2eeoik+QQIM/HM9z
oTkP0C4fh2i01fSGI9VMRAFWKg/j56N9aEZ5PkE1vf3txqaPttbJiXTcRQiemXzh
NHN3Te4h2mt7YQXxLpgdDNUvCg+vuo79tvrAyuxLTCxaQl+f+3KFBs3Dfy1I0BPg
hrRW2AB6BcByD1qZcepypky9t8azsQwB75E0QeBWvpk6q5yqSI40qU0GeHfGMaXy
yDSOutIY4roZj1jRfOzVO+hn1npGuA46s3sjsubUN+v+o2mSl6ts23hl8O3e1b57
7J/1v4aVqpjfizONhGXPkWNOyo9IcYdS9h5ZQmdqf9Xq7aUFFjFpeiIPvyYrXuje
58r/0hxcvB0yoHAJyohDg+pF/gT1emoM06XFvpHUyNhZbRK9WLGSlhjVoJhHPzeG
2/PMdUeuXvt9gbqxkle8KlSgPLOsOB8qkP/k8zP4LeUIxc+KBispTAnB3BPFXlOe
Py4xrkG2O4tQk4cbSN2XXDfEMEbMfZwFCAfLC0IgokF3wNZcKtPEYGWWbdUhIau/
mpjA0jDtoCVny8rIckNGy6S8mGJRCXernGuKUEaAkbP2Or1pDF2FvQDV2qqRRJsr
NYMMSC2GZuRQ0iRWDNzod++ZqlH8s3HCWbEvlLFgyJLYMdIDMS2j9jYCD/qsB6Hh
PX8ElNfsCDDGyDiBZHj0muIMddwi7KmySyyK4dAoyljL7S3K4M8Kq9WoxwzVN8ZN
aj1dCiqHK75CWrTSqHb2Vh1Yt67J60kM48F6cuFKAhHcuDuUrLNBjtOgtjtkis2j
UyYxvPcH1pLv3Cpajgyip7DYqPmeYhPgBib4K9ybZVJsk5YNorUQVZFUMB21jkX3
aDQdZUAAO+QjbEJLB98a2YqkP9bMWPjSuqEbOo5n79GqKW6ZhciU3x5KBDBhsREQ
J8Nf5PIg9hMl7rlhsa+Q25EEpQhH0qhBMbkw125MtBoFBLZjkrpdMmKVvbQWx78X
h9fae3cEMpHzBUxCnEp15VtmtMmOLfGnPvjo2KC5R5QjRpTTElAnMOcMdWg3l7lI
isZcthCff4U90OtD2K6c4gi8GHFhD6/b9hzWViYVY7/Qo17X6GmD3vbN/q/r1V0f
KHxhjhCb4r+QodMGogarRWL5irppw9+jcZn16Gkmoq6F+7Xx+p/Fj1j1PNPw+V0v
O9stfbwBZ6OSncaEd8DKfIEgxvjG1B06KVMHpi9/5K2T2gjJZJjhOuGvvmzEeBhw
YMov1X5yaC3/mRcqr2ditp8Hzbrgfxdh6U6Ny8XQDHw0NPsT4eBNIxkddG8ygJT+
AZNcqZz+y9MPyxT7E78kX3K8oBmJe9M1B67LLMFmdc93kCB/+9Vas9udXQ4OutrP
kXd78iUerksOtTYBR93sRg7P36cSEy0aWg+iKKxIJ+E8lWQuWY+OBLzqQgcAaB+Z
2ePb/JcneqPlGFWNywm66V5rCCiB5uSfk04Gf/rV+N02dBlNv6KXF9Guty2xPMyQ
Opc2NnUM7vI0zw37F08lNcrj7sIk1rtS8Z1IaejfdjE7MQD4hWCMcpnwj30jUbFI
+vxg8x0F7pe4CiiOYSRU2OUqcjn6yvYNh48vauMyBLamxp0CtyUtrKFHoVy2D2dk
MnPZ5avREzIm7NT8w8/aG8uV2GPruYJJtQIs7TxahGzLyO8BqsSRNdJ9OUOp50+J
ZMOVXgQfhuJI0/nlM51dl86OJlpA3LQqUiW3j4TcrNPQ6Ct+lO4peb92NbOatGVS
lCtj5p9C6Cn+IWmkuwgSJnjFTmrEmto6tpHEUWf0TCXL3gySAP27UNoxAsAfKl4K
naOAbyvpceAJ4lH4pO0c4b7hXtO6iX3Uh195yMwGzbP+Wdq9Pke+a26ZsR0kr77j
GxVwJ8C/jnygHXwPeAH3Xpq1nvMB0lUbbXnTNVyT35uk98OIPFhSIJp6szHc1SEN
sngkdBKpmTq065EzDRX+hamYBDNoSYYVW7eL2/XBhnQPBLF3Nu4qdid8Qh6jyOXQ
BWCakZN3jOLJW5NPRnDLr3FirhPT5+RNu4qd0SlD/fe+/MmQwdbM8YmDKxbyJPDU
lqXxtUlmr+LeFcaoNcp8AHyATaaMa5rDgYpvXHvU4u3HJIWCDSDrSIUWVG3W4i8c
1mHdvLD4BTh5UfaGN44GwwvZTA7oBlpxVZrIfiVuQxETf/HPDbcTY/4p96LSv8Ws
eodTc8xsQNknAybjRxxWM9Ai8lFYLma1KP2m3VXcS5cDWHC1aY9LRo5bKgBKde9u
o45BZMuLPNS1Wgx/583oE/vUFbAWfgWJK/epHkjO55TwXa3/xr4M2fpVAnvfgZNa
iwT52YKDKmSxzFhs9YWL3Q+QTfMbeCADQMUjnttCl+g116rvTERfNGQ0ZMA/kmC/
Cr4AADFfOLmAmNS5ye2BOPb0T5wSU/S95DaKFgwQpWI2ufwt8sLMJ6mBWzuCS6gg
P93YxRfZKoNXcsH+2uRZF1ss07zw0J4WXa6CpKq6q8LKOTewAgM1DVFiyV2tJSmj
D6MqTNla0otj+u+GXbhkCHCkRkbHJtmWBibLjqfI9N8Do3ojto/9U8sQ2qqBb2oE
GSxvYquHdpQVJqmlFDcwpxl2nTBUgpWSAQ0Cqwqw8nm0WCQyiVfVH3IGxLQzOUn9
NtCZHIY/H9ikfAj+dWoENRi6fyloal4wHeKj8TjXZ8lg3S8B+jouoLvmuCfUrAVn
nmd4bAfwfpCgg+K7VMdrzveDg5u/3xk2H3iv/0oysVG8qaqeZ4e5nbf1mO4wn3K+
uo0D2LTrGRkn8klh+kiwBZOzwUdITLX798UopalqLQAHPnC4AcvZCmXglveqyvAY
S1+jjZSCbs+bX4uNfG1bw97h5iuNUp9FI4IjYIl9vl+JyzVfMIOT2gDQRzpWYlhr
1T9W4t9OQ41A+R0awAXxBvsU6RloeZsq1xI6nGSuMlsns2cAd6/d3s9n8xv3qWVJ
Uxxm9gbioYh4Zpa6KKLDB0cAXgc+omZ14ucJtFOe2D3heEORsOR4FjkKJ7+PoTQS
ssYRuoFdH0DcRUL3dv0XYtFXYaoWbS8o95jynsZ3m6cRSISA+wTIqVKxezKdaUNF
wmR/63tWUvkCu3f3m0WCz6mbY73PPQJxGJ3e6Bb0fGxdjeQZBL0mYpWPCA8MEwvu
3k2EcGYrTuVi7aIREJAvtXKmED50ZJMuORYwh8mxE4eGHph7W14yRsoQt3XAF4Db
WTGiQRX3fPvhZtvh3OpesGResOC7glU/gPU8XbDWQmv8jCaaxxEOzHTaNWKKW/SV
wv/gJRNcKDjchua7chtnM2Iwry0FUcwOZWoxp9WweKPE56uLSMQijiN25sjiE3X8
EnVZ/wDYGsMJR6si/+gNrLaQNtP3gwR+Bre59mo/tDZLvxFIe/cshF086iRV5eF/
nLj/kmquB9MNm4hBCG/zC6xPtxarKWLHoSB66PlVrf3nlcFDmrmHuZXgMdmBrSI7
zKZE1+G+GJMO/2Ausb/bSNCu7p1E74Ma7NtHns3hgI2sXODUYtObjL2Lg75ny602
dcmFAasd2FE83tYLvI0vtruSy6k7QnRIhqZ+EjHRy4wlOpxMQs8yPvDWNlWdK0kc
Qs+aLZ+Du9T7p4/YVif/rrV/xNsk/jALEj+rG54QuGGFOCXQWmYatZIOJaQz9Q8f
Ggt+WjeId9mi0N5QC+p6nhK2BAodLYPISEAMtip3eJ596auBiOK1p2Jm+2lGWwjf
25DGQVBDGg40i7iJSC2roFNTSyS4l1nef7N+zLzAUN1BK7vGYo8Urikdpqn9/fY5
fbnr+VJydlxKK7V1hCOWKxEEbVbTJ6NdOGjcXOuk8mrr1M9xlE+/XwdrO7HdFm5Y
BUpmU1dDB6uUHQfZfx04n+cmm5vK2YCXNSLtO0QKnD++f+TTKOutlpH6+1uxyEbj
nvU+zQztSAbLG8+ngWDgrq2zU6tHZdcT8q/KTi2Hw/mUy0ut+eK+OZx6MHgbLh08
ibr5qYkJUAntaoVzcYyJ4MX0Il1E0xmF6U2b2YM9pR3CZdnXmbk84+uurZrxsJE+
nJFaOxoG3Maq6QEo4JEe0ZxDl5FG4FjHjUoHlCiOq17afy6n4PzIhk9qc8xLAkyL
yvEUfzh6rPYEYyvm/FRoiEJ0lEFEIzl+Dv0h6zHs7WbEHm/PyB4Bx6d4N91zFxXO
fkyzynLOUNogzdWpSBrCqrwjfWC8Qz4CqVSR8DQORzaJ6r1xIaVETA7DSS4NEMLd
YWjCEv6S/+YCu90aC0Kty7S5cn238kbJWm2ix8RwRan69eCElcgQsHNAmnNkLQUK
mT3qpPmcSd1Gt1TRKI0nt1k0VJ4AyFLUfiwKrxQYYD+5Q6Tfpbn0BUclFwGsfvEK
lIItxOSZKxdRiO3AHjbVhauksIGTYGipKjvBGMOK3T/T2Rx+hJY8K3GkmMQPN+WN
TPurx7BnavClMNcH9dWYS6YR/MsAzjJN/m6Frs6CLigA0k9oQ157lL9jnttr6sWE
2Yf8uh/Dnj5gMpTYeFojnyl0aBSOfxavIuM5bL036toGJdKrjZ/1OJtQIZH2e0nS
mw0W10yNXLY5DbZ4alyiRlKnSWDtLmxvRXM5wgqrgvRhU06e8LrByfpT7aQbpRDJ
ThqyQMcCGLysdmYdPLBLGH8uJDL1MMRBDlRF8sIlk4X3sybi8YinPdUDQD9YqB4C
Ckd1gJIMOErA+Y+mkm6d3QJn5dtRs5PbaXUL0mlttPefMGmJLAoWCDbNEDSYqSwd
/qcCwcdbfDbvfzJe5+GEsALlnk9uo//jUkM/o3AaFbB+ly65fUIy/079zCrEdrpW
9KHp51tr/kT3rGQvX6Knn/CClklpSVBO/x99iwBPTXBTEPNYPWqo8QyRWDjddMVH
oRt72Cyvv70ktknLeJuuX+lTHCof0JqdDrP3FeJV86U0SQBTuebTI3ViXZObZWDY
0/0ChaHZdzVpenHZHOnm+NOcktjkTtvV74by4PPiDazRtEfKUJjEpUHbq1+dgR0O
7kPqWc/D8uPQ7jZiiSovh46yUUQlNdPUBina3g4D1Zq0RsqVfKGz42vaK7uhxQAZ
d7t7ITBjgJcDlPfKN1duFHHefD9NMajDiCXsAJvQiMw9Bu1MEGeBz4mzr04sEWwe
qBjMj8epm1A1VkE72CDcETxkezPo7+wMeUCvAv49uqYgY/Dyc925/g3Uxsw37sXM
frjF7A9TJ7FicpibyoUHfGWaoSCTCSWZjOi00jbzi7wd0ohJM67vGOa/rwRHYYIv
RMV2kePoRtzg2/GEYHhLd87c/AmlFJfJpAjd53awxYZFY1CS+lOT7tHxjdKhtEe5
lrT8EGDz3tnpKzqk4thoEJKbciBYeUGAiewr6cWP5fh7HtReli/uKHUMmRkGHtDP
8Co1NTNO+s6lpM5GaxuCZuk/wuG6NHBqw3aq3BblLu0/mxN9Fmavsvgoc7mNQlZZ
jXYD1D2JDScP4BO4gVrpKqtCDSV3xbNn3RO3aRDPvcvYj/bpRnDFabuYo6qp9ONL
mc+KOqQTt2inesjOt2dnrkJxta2qd5f+QbtsCpmFUe+CN/oVMC0HgKOJhpd00T7p
zYrWxBtbEjkFqWSuVNZHVYxSdTPjUgtArI/AfylWR19fMpS2tEBWZE3/UOjI1etI
zdVqK1T+krA8LkwitsKqANiHcWPhSU8se2qvVvkaTNYgOw78VKqydI1pR34ZW4dN
pby9lWihSPWAIEHwv1279fSOq6g6HCstc7of6/7b6sya48XKeKE2/WaxiIbJ7jBC
Filp/EZmFOszDxkjOC8jXYcqok9TQsNlsjvhwLVeDDfiD4Dvna6WOHoBkxKSAm0U
i/buqTbF4RrTC8DFrFwo6N5ymllhoxKY1wJRVD+CMzBmYRNYnx5PjENPgwemhuJ7
/LInUZS1nkL3mu3eCKl6xI8KvvYlsVNsX+WNil9X0D5VPcFZJUxZssfT7ThLWvFX
JqRC/noL38fYPlD3VmHNLkqhu2GjMH0f8+DO/F/Pmeg0Hu5NLV/HvwPWPXHXOP4m
4cSVCU0hrUN1oq5FZnYu2R6dSDaaB3GJTfIlMaoOmopsn3d/vPq4vZur/URf7n+B
YRKAR4X17/E0WRo+8kchHQqMzEl7Sw+zpitDVdN782qbNaxvTZyQTRX6seqrueDC
/W/sGK5GG9Iu0g78LjdsVDiAtCiSzq3dlgebSVEVAYUQTg8lijkrgnGtaIAoNfND
YWC9IF4uRBsbVazp/iVjHgksQipLTnvy2JtUnfeANKBjYggJeY0Bg+GwjoL5WS9X
B87uOe8NHoqIUMchGyG99zwuTEsGd6hFfr5lGuSr/mf77c/nKQRfDef4ELKJdFTg
BBjPibVVPIEGkvYS+/7+jObX5/vWrANg9PVZxOqCijros6w5QOQh8U2VIexkdDcK
5ujuQEW46kyAewd3zBlW7TB+zjocv/vPLhMRcA280uPJ1n1K7buxLWnUZu6H5D9s
i1dNCs87tAgYQbxBZTamd9vvdIT4baRLFXT65MaELznej15egVy+G8gw4VKyFlgX
CjBnbZyEuxMcee44zVdxQVhwZrXKydo+LJgz4ctbxMGIlOK4NjpnGrF0iCW5Vu8c
j2BctwXTTQYpYn0YJhGfYIg6NPuRoFFq2svQALA5ZGuCb7fb3gH9MbLYq+Xegj7+
nWa+2BrMc+4eFkOvMtSgAVcr0y3m5UXcvlvCUdYkWDw38ikIFozo0mhaRViiz/Ex
Ut68FF14j3YBeWBrGFlu0l+mx4+dBV2VQw2aKbskxIZ6+5DlDD0cJqlRLsqUhpUE
N+AW+bQwL+zYsqa+wMnuhRBL3IxwO5S9sjuWtszofDjMVinFFXLQv9Q+ZuuJPr8l
Kg96cdM1iLZqc+NBiGXNXVhnOIftPITRzGyK5vlmKySbsKj+e+RmPT/vpb5h9E10
qZoepbl5Ohbv3qC/KqrJt7QBkOtU6GL1VSvEiljqP0b3rzbebsUbhE1Wze0O+TaI
0zbgRC9W8GACmcExwV8c6NUUEA/kel2Hrni3l6IeiCrWQ9XGgNwaJtwhv2OJZITQ
ju3mh15rXBA+UBNjTZBfdxOhOO01dEw1HffHv8z00pv0svcu2dlGnpriYgVv8/yF
XdXArvyXKd1l2fl3oaQonqd53DYhYrQz2ZMdcJ1SmEEgJ+OxKic7Zc9pYCsBA7lR
fBp3V/gQ1f0mZKzT/BGh9tuvYXJgjFQYgcK9J3Vqfp1zRdqH2E6HkpfUCmxSDkm7
dyk/qg5IFIQbMWDj76OPnw/H0IdtzMi6xCyn0fJmDRIp09YDgZ1gpdK6FIJjDlYj
9m7tRNJoD7Qo6XwQUJGSvHw57sPeBC8tNBwG06TH/SX23pigDK7uhvpi6ZPh8U2V
eLCM5n/xggp3LA99ac76vzSgP3CyKW8wP2lntjCErcKBkkSY8ENqYvhngc5tAeeg
Wg7VdQCTqHBOtV+hegN6bSkYEeys3gD8gIcAx1g55tRnVz1Qg2tDYiInE2I8WbmL
GyhWW0N/SdeE4V9xkGgYXo49sDFqjOr5sBW1/nQsytS5jbi+LAIgWywjWBKqc28k
Quq/9SMcsbV9uGjI6tNN3cKK+nTYSR0bs2mIkESUhuSoyrFbyXLgwdWUrbFRdjQt
SQ0UxxhyxK1nX5UDspjayCSkXaCamkubsZUL5N21HTls7/DwMJxwBwF/VUlnYUuI
ZsUEotW0y1P1b4wK/FtZnodQkhfIEtTXiWvCtxM9HxpZw2EkgglJocMhvkuClXS+
toxnzBzVC2Z+xkeWeDcWEJc6goE/B57MiK494PmEivt+BlhoitZhqRbeEpdwki04
+Ov6tEtSgtdiaBp+Fu0eWUl4+ya+zhR/d/+ywkric724n3GHblB2BKknV4aF5Foo
LKrVkqvYhrQasnAc5Yb68C7h5p5YWuYvyWzz4+lx2M+xZsGuxtfQ4fIj0iQaebse
GrsoJfJa2zFvC6jI/pcqFyfg5QZt7lD0H5/aXKchZbQd8wCXlT9cvvA5BPDJd7FQ
C6HcTGT4FVPKs3ZonBcsf2LsUoB+grssGplJxsyosNIxuJJjLoYWpOZKMFGDUFTc
+/L5IrftnzV18d9pHswmxNzFDN/VTKOwXCYnKYGHCWxRl2btiUoeexYwGl9BdEWg
/G2+yWgJEQvUQJHgK8TJZWifSNr14BWR+08pPp2NEGfxh0Mn2IYkgTti2mmM0Lf+
7sKko72u1/nXTVo/LwrZOEfwNbzhg//Pz79+nkne0AYISIkgdpZISb+JHPeNFUIo
bQtA79u3iIJhPDUf8A9AnQRAAT2yXX5IcsVeP4T+ExE/BKHdh23eUB59pIXm5Q0Z
Y2gbiw+UMUd0/p1D8A+Zu8Oh01r8Ql3fu6m1zozxeT0rbVMHrFrAx2e/eYUWFTXP
M0TGV17CQUqCLZceCXGuGJlrloBYp8N85WUYDCsI+EZG8Hrh72MNcs5+7nSI8/yL
mg9DYtXEcorsEJoKO8JcGefQopktcWvxqL3DRjdqLkyixDrqgBv6NP4wUmaivfy0
2eVIjtOj+d9+SguGW3fE7AIM1xT/cL4n5B0cXqbF6hN/m0h6WwX8uIe9IxTKvhEF
X8+fTdS9KaRkTL59Br10vaBKprA3G69O09YQfEukD7Z3+2QJ3zqgxpPwqgTUHdgg
PzCAtMdpfWb8zpkoz/HjpwG7hTQ4ch5iXqVGvDaoNj/J53DnxuHPjPrszxuMfqoM
s5aD8HM9jRpfmEHnnvgVYmSgkr1sgfenKFGB5OHt6fYMIWktwF5k9YwqW3wOMrya
or90C/ywju/D3j/DTXxNRUwFJC39f3E4V+d4Jvxt7qH+rp1Tz77HXweesPVRZKrF
AzFAs3kwEjwSJKaZim6H74AtUucFoD1m1hLveFz6rWBY5VsWKHvmx+RxAzXyVNoT
s/KWWXiB+ugWs/q3QU48yW3muDCkWQfiQp792XIKSnMVSVONGVJrUEXu5iDTj5S2
j4bRfMxTgO7oX5ir7IQap4LOt6LlhthDsrcxhF6mbdp4bnAWSVPBZWMpedg+JziP
6x4AbdRV6xzg3Nn3I4th0DdkEUzWpQEMA2c23oW1GKUpxNQgBaiUikqOq15vF+EC
C6yJj1pQz22WVbQwmm31UGIrcYJCmndChpXFcNeM2MeP8n3LpC+sJ/G2uyWcJlmL
mHrQ7/e8c46Y+UHqSvhGdcp+LTRsYAVtvogDMrUoHXMf1/jg3HcCDK0XoXtkh1yn
LorAMVsU+X0R17+As2dll7cO4AIXrUEyFlZbkKgmMDh9eZdMZIconZ2vhLiGvjhW
dQjz8N6P0JFNUZueax7mwW3DiQyQA76CfjqG/Kz5bdHOOITUoMqUeSjpBLu2fXf9
XR7VG61tS2KVI5EQBaKk9soCB+AZRpGu2jgNT/Ap43HCL/GD/NHwFI6D7Kkr1a8U
hr9xNkFMUHD5QdLaGp183WaehQUg8WBZh9HAwHv0vcP/0UVSrHmYh6zT6adnXQoO
7zYXNREKJ7c908eTbV8Z9donDlFW0hB39DnDMyAoNr48eaq6tnm3R0x45dwzCNSt
BuzCH/+r3ZrnVM9Ux+4NJPPrO9zWIbgwkVMRPmmzTC7zyqHR8uC+MvmzJ533M3q1
5hCbDzmomsJV41HFFqHI2Ohq4l5iPIkDwNbPDea2tuZHUv1gmF/B5iveLqGC+e67
Nmr5tuDitW79bW1rGAFOy9IHAfXsEMPfzsXM3SOIDp2kkLf1NP1vxshA1QCVcL8Q
UeA9zJAerTAAHJ8RPYeIcbFWb7IYFZ6bBWZImTtAVq/HDGn3l6c58CI3gdeoTI2B
Itwd9JVii7Y6qpWtQTWAImbipz3H8arST9+dKcSH8BvPYt1wmpnQBZ6dUh0u4UI5
m6YNpjIZP1OdNXcaZ3jTh484lgPjuCGXv03Oi1nAu79tKo61D3nLlUxjS4LagR/G
cdZsNSd/bHxSY38g9bMVurB3EMTVHM0IoAvpoVdZupyi0oYgbbTIZVwxYsgv+uWx
mej2tug2A+xWGhPjqWjFHXfaJNzaAcwmtrMlyjmkKYXam+Sjfb/tgkSeMjYG0WWN
9E30Vtzyg834QHftdY9Dod3c6B8KRUpkFds6vY9mTP0nzRjNYlhEX/itNfkITZ7r
HLXzbM8+4oqzvzsMOe0SG9P6UT1G6BSAK0OxaAHvxH9V0Dd2oUjKXZmumRU8droN
cW0NH3EOuvpkWRBmi4oobMH0bLmJwRc4AmECurdF5rFb8zsgk76R3VACBiN1EmmC
D7w1yLKvYLP+s0Oe9w6UEIzQ5HVnlm44RVKK/ix30j89tMarEYaufs+J6j45PHbB
yqMKaKM02xLcop2WMndvtdNmGrvQBZRHbEx0RfM4AjtnriB8u0pcmhEqZyXGfSNU
JrlPnaPsrIIMiBjyjjPC+11GR6E5eC3j5exEIPlU3b7nU2nEs4npqq+OAgY5C/pB
POHewkoiH3eTjZPzj7lcI6LGQ/pugUXf9bkVJVVORhHwzlSeHGZ8N1P26JZB8cWv
5Fkv5xesewBL8sMrm/VcJ/91xpiZVNwmGIjpXhsdkkjcdwH0wemxd47F7AWbV/5f
U5nGezOJH43dH7a9DFQzb+ttfZggr5cOe8onE2yqR/sGzGS2N4Pg2erLbE5Cn4VX
qRulRfOOcn2QQsfQKvtIblGyVcgiSmNnxT7eCmnH09g3Mq+Il1b2jjl1U6dvqzJH
0kNWnCz8ksMtpq6RuSC5qk1tTVvOq/rDRnfCsWL9KuOHEoocgfNkWV1DdvLzKWpx
OSjW2djRYFw/+sfdNhR9rXVeD1avnj2OKS+eAFpcDAFmDwKE0wxUqdEUQD6gjv9z
kwXDmTtykpV3m7lyadJQo2UqpjiAJ9LUbgZ1KLxrtmzqgRnRqR6frh4raXtaM5wg
JQLppjfgVFZgOthbVB+m7D/PM/bBnAHB1NBlV00zap0Lwl4vQ2ZIEwnC+ViqoSm/
w6GQgT5Hc2JNeZKU3Scnm6wA+ubhPOCqjK4dcyCPJYI8D3E60x9t8gC6ubHRbRQb
t16+PoKr9dXQ1aOm0aZ19GDXICYTUaWg0mfxPx11a/VrBU4H/+uHlExWmAijuwvd
kqbqKHtSSa7B+qaJxf/qhmIxeJ0LNbyz145AnGcv57DRW0jytmGTZDDdgiuQpNkw
/AHA2rDG1X5HtJ1n0VEUaMpmIGldZ93CdCO5XSyywp2rHkq3wYtwiUlxI+Xrj2Kf
1WEOJpmK39M5+wwWLCZeYZZXQo2S6gCJ+LGQsN103T2gctSRwFdFQBTbH1IjT6oT
DcHpy/288lfuFEru8p4u7odArD8qruMoToidmWXpDsDWqXfKGoJNT1cCnQUS/gj0
B+NvDM1yJPqR0kM+1sEWdZkdi3dbOOJktrglxYmvub0qiE+VkHrs+7Sxracq3YVf
e/KwcqLNPjdJ+5M5WsCIpdt8uN8oJHfozbLJaiZh5gaTwxxF6YqQm7lJ4qzk4wGs
9X/D8UhCXdRKYtsLqZYoDwXkqagLJI00el76J5hdpXJWFC6bHYDnmmsl1dGHqpNS
/f8D2sN8VH0P3mOzV9BKpI/vkRh95vAa2q+wjdeMuKseScN9ONEwGkapr3igMFzr
jEhvnG4BMFiaQeAEAbqDixp34MTrZrstLOy+hlMo3PbMG+DQ1KL20PEBc8x2lL3b
j2T8cwlEwXcb6fN0rnQq05zZwwCVLxCQgA7iyAGgnXckI2ak0SUYR1VqkxElQyhS
B2+WPWl1N1+GOaw+wnV0+0lCng7PlNbMIEuQ/iCDiK0NU9N7UrZdqRseWxLmPgkn
1KaOU3FeybAATzj0zBNpDmabLXVMPfwHJm7GnJAW+nAGcMqrHf2OsXuJJ10lx9ld
PRnadppS4GDs4i9DC8HbX7WugWVSSjFKGXJYiboc6rDBVYw0AVhATxvDb0PynHTk
f9A2e35gO1sjidTPCPuHpkEHsS/2qR7WkySTupkR7NPW+a5lnSzez0klFsh08i1P
Exd3bJjzK+tgVPezcwf4582A8+AlwcHzP8s10jGjpqkIlwSwNzEycRFPHxDgP93q
08c/GfaMBJQZsIQ3ZQYnioj4LIqlKMZJ0DyICflFpPRLhMwDXs2/khTT+VIXewNA
oWoOS3onuQ8DPUoCn9fBaXK9e20PUnn4VmxuXVT7oGR4aTHR9q9TtNQnftOkFhYj
hicpz2VpyFrqXetTFmmARlhPW87w5MAhNpGVlOSlggw0TGFQ4ZASMBtbWdQ3D3ET
PGBuM2iZvbcx+pvom7uR0v2Ojp4AeTDhnm5NnZSfSoTjP033s8N3BztLtALrJk3S
4wsQi367krk5AuJdpnQXOffpvVLQyO5aVnUmkvw3UyYaKGEtkN9SDb7ijOgcmlVK
PGFjbTPrxeZxPBoyDD+AhpIJcIPq4l6msjbZ+we2TSTnAyVmIq5s93HSrTjyd/Yg
qylDO3Nl2U64qPB0WKxJqwk08Gd7HcpyzFhyftbl4Qppo4Ixs94fou0WMwldqlJ+
JQ4O4PYItmhKs2R9t2mRwo9v39zm83IBLHWZ0ilOtC0SqnM0lK+lF7yS+lqWd4xN
1SqeMvJCSALKi765JFjnLlDoOo4Br0FKZtn3V0rL83tRgcmhi62wYerwVXlISzUD
vTVzYSxHb6SHdWSm/e+ttJAMtTO7ciB8yvVOiqTKwSg0fNJS7GY52pOADC+LUypF
mhN1F8js5PWD3Sx2GQJO4NafNoVvQdoYEAhIycnJUk6PmYGxs9GbJpFdUox9KNp7
rLSuL3lilp/TB+BgNkPD3K8moYxZbdMlqH2KZyecUW5AQha9/PKCvxAyvD1h5Qth
V/ahf9rUcc3b6u3HyNXJwbQ+4ZFDlDp+zh2Dj6ckIT0V/K2nK/Sh60y04pFYTnpX
oJbBlmJiv48LZgyWte+AxIL9OJ98iquw+WaQzd8RWIcW3ccuQ7hIFJHeiDBpzDE7
BzmREivPgp1X584K/cqJBcFb7cRSYDneAEY/n907218IY9aMYaYNSzyr80vQocrR
AEn+tYm3YMkEwB1OwdJBNCXon2M7/uZ5/k79UlROt/ewPV6SqdyR67cBiIZmyXai
aI+mZYHcIP+KEeDs9r1sa1UmOF4ehvanLCoD47ZDUKt1gnuN/9bdIc3bH2/PiKMg
X+CfOwXCYbNoUeB+cAh+b8ObsZj76olV3hHK4uIeudoY0IoWScL5WOotuWVTC1Gd
bN/hUZ/34OXlcajXKOv9WfkAJGtSE1PAmrBba4swnvd4DVlZd1p+ncDzRekS9sS3
fNm6phJ+K140azfCILdqPEE3z7wMdIFUPihO8HdR9UXtaQZbD7FnuxK8bAmg92PU
mBNb6l/OzYt3AyJGthQh29n9fumKtAx+UzBnF9a9NVdwHoYhAZ6nlhb5klebd03Y
IxXwBaHK6CHiyCLs7LmxxPLGOoSP5TOg7/VEP6vcyDmOfe9zDgXCYxa109+u37/J
jHdA2mZ2uGXQdb8AzYwYoHu7kPxzTWmQh/RYXKBRfe6sJkV25SEQm23rVfazFLhK
lJwS3YCbnJk5wlRyXFsMEqV36xzfDofPbU6J4VcxtuLlxUQSlBzF3mniQZ/UrbI2
tdeJ7eN787Odp1TtSLlD4VyFCc3aGFT//vttptwk1atS0sjYY1/o6N+/bJhRsWcI
61HaBjRg1eF6DILPsRq7YpxY167criY3lfyjahHJLDX5w6HRwRvZPZEiqCrV3FmR
P5TMADzV4TUzxLOoDcj0l1ZMdqSc+3sCNuhWb5N6RhZB1B9u2gjVFhd7XE9P1KSu
V7D9EwbqlkwJqVySm0Sb4UY/yrUbE9ZsMM4prpVr1VIgiu4OPCtMJYF79GlEa6wW
CWcjF6hin1mzVWD2391/MsB+5P8HATdzsL0oLXFNMLniwuNX1W9hXXPcq1XLkhXM
BqmfUi19xoCAaJ56TrbbLw93ibAXbySaCCbfncgvhSdbdJ9QIOiihWHyqo/Kb6w/
iD9tR9Zsx8NZMTgd/4oaswIJCxm3YuhmGPAuNDHEdqwGydVzdHtsm70akxShuZae
qRZw6rXeH7MtlyEB0ar2tS5t63avxE4EDHHvR2OaGCT4VYW9jiO8SZKZL8CMqxDO
WtdRx7OAcawQ8JNgqtRh0g+mqbCmaaX/Y5lFp35C1dqmcJjWntio0VFhuR1IQbvr
/YQUxj74a+B0kjqn7vLQCxoMUwfhgeRqBGNSt6wKDj5cnaBDsi12y+0j+APMyUsr
gxNNsfgbhn7Au3gRgYqsiOYGfqem6NdOFvuvLZGB0vR4SgRVGyHIs8asyq42e/Hi
Uq4AscPtgOdL4aQzQFTlGAnRJ8P8uUGrn7655+NWa3T23IH9bxR7awjwQU2QFZ8l
Lj5h7H05Os1HxiJEGjsdUYTsAhZv3jiE1YnMaBVa+f1PtwghTps8IsqQpe+Cl2vt
wkUuahH3E42+clfkGeLDONyYWP5PQhsj6Lq70xOkgerGw9BixvqBYxN0HXlZXKax
w883O8tR1ODOiuBa2IktTU/kiEIIER0DMe4D91lBqED/qi3G4JFKDxO8Zykz8Cp5
7yCfCWSNnPB/FRV8sbs17MLc533BRSSBOBFo7A6EV4UB6MNwq7sOYwzn08Tpj/RG
WBz2Msk6+xFRVGfzHFXvenH+xAximHXogO9LekNkdxfN5ZFtMvKNewlry6KW+6NN
PJTaNFWDRKWrvKy2p28fu/Ps/Of7AffWKRqlkiAfD8UT3B3GXw/e0W2U1W8pJNZ7
qHIUY+At0nHlAPgVjgMU4DIzu7eS6MRAE9kxTD7G6qQvDif3T0cALhb6CILlCQld
hSuGNB4f+zRSkg0YYEBJJGxlDij3NYinShVfpJFI3a3tIH/RJKqBvHkzghNcShmY
urcYMvSS0UYz8ZIpgmCBRgyp4IdaZz9btX8Uib6qEFWNNwLzQ1y9uaL5FrL1GrAd
ELl2ghSs7+dzdU3XBKnT0cxdWQCRhce2850kdoUptfDGxcoXSPLF12BoTjlurygO
P+1Z2MKYSC97e1Y1DM5oIo+ller/y8E4u85Xr+Y8sS6OOW5o56JPGtWA0J3fRyPg
ZBnnm0dkiHljSbLg7XXbn56OR8zWfhMcVxZ1PZNQ828Yrww6bicShsXDAYIRyAxt
FkaOKQ7kBrdWM57AsEXafrn91bk9BcbpAHqaXfwhTY0F1sXlpgjoBjahho1XGj5X
B7AHyYTrMkG531ltObgPd+ToAlEcHmfGO2TuJnMIHS7BLUYJf+bBpXUubRUs5Nxu
DHkYkENoJJdlWEzrYIWouhBz1EbJ+H2uB2MS/QfS6nuVoSu6UKa2PmUHOBconZ+V
xVEwQJat20YfuE8wemtG/TuFNj7wrGku437P9azzdCm/c2l7E6NW1+gXeqmXBlWZ
Bg+j/SLJ45x78ReTaP80LvJfbwKYj6AMZlafgIdoh4wFDVFHlPGa+cbMYj54+eHq
IjIB84p6zEEOhCeBKpxSe+T/pnXTKy9U1xIa6AAkKesqCHf/Emp9v9Ew/m+3a+Ud
mxk9xBy35VlcASCHjNusFBkAe+1A7UQNPMd0xRE3SiE9vX6c/KO48YpfKEwmW3o9
CFZPf7ymQvorNrCMy3m13fai0zTckzoEy1YHZuG//+sH5gkkpH+8tFGe5e5iz8xF
XT438OXG928S64HpEo4rlVd02SfJTW4oW0F5kzsEIUQQuUJgJD7Rwi4k9g2/5s1a
toBDFKilKlSoFFnLlog9FcjVpZ1OHY/YGzPg3hd8+hwAdsuqhZhodxDk7mATtPLB
qwb6ijv0JVHKQqE/VyEwrrePgVOtEMtAYTNdzH1RkQsShXWhsUxnEKuihWvweCGj
SSChD2s6O4g9Vnwosx63riFKHISqS4FP9THrroS+dsIldi6w0Wc2VHjOpQPpAbTK
Hx8OJa3lk1DLYYNwBE1xiMQNYV2CZDQatQ2VNyKVdfS/daPGotji8y1epD+rSFzo
ht7kgWK0kHmNSh2ScjLmo4xnC72Mu9jKH1+SqP/qJXWSesUMj0i2Qlx6oMUagvfs
N4WpZiOtLMMw1oJIKHZlnNl2WNlX8FFYAP1BfEjbuYYMijfxP9kaB8t2GxZMUEje
sud1DFpwKVPkDnyNzsa2qmCn+6KfdHWNcnR871DRKox0tF2DqKM9tGvqmC+PSBcY
iTObnuiJp9lK903Ax047xxDd5i40Ie7lUu7+zAYhfFo26k46dwhG7ppDKK+jPmFV
MNn3r+B5CANMqi2ExUi/4x5ztvL/DHJf2pkZ/gODmx+etxlclwlHYvSn/83fOG/a
6x22EGv2krfvxj81kuHbOoJWwlVCxGIX3djlI2AecnmRgnzjunZv0+JYzQ00jfFs
JhgKMPt5nfnBP0ZWveRi97+c3SWPvYJgWhY7uKPklwBGogmkUqmPJauEYwXJVFV+
Dl5lhm7Xn4JumEMy7QhUBmq+SVSFuFVQt/ZwyuwL51KOoN7r+ksUrRirv84xxmaL
Js950pieC/i+Wsmr7FbINv7RQcWrMoIVGGc0gtsr2oBhnK72cYsC+MKEl1I7Qtb7
/koORdFE+xToH3JkkFfVOb8YYC/795wuud5K1V1ONN19rWXOtqGngyM3pLfuC3VI
VFBGo8sTkQFW9zwwu5v7XLGLbikl3nFkQDBv+cd25eh5Hb0XxU0cD6Faq0oDWi+w
vLW2N7wMqRCrGtPpIZKg1lAWhvnDsBkFPyqRx0/2LPzB14Y70HILPbs6QYj5pNin
/OQAImODCR6J9VaQ6atI/fZrBwsa7b8kYWwmDUbupjT2UvAE8+J6fGaWMnlQXG/N
4SSM5G+3GIpvOVZkCXtFwGe3PB2xEX+eh4VddACC+zEkfYTSbX6roLnvAkp4DZck
VXoQQyGRnPjYp4nZEoHvxwJH0VqlZD2UL5w9JpWlTxMxiq5dTT3SZSksVueBjeaL
HhnlJ923UUEjSFdRgLPThTtCClf5heZyyMbauKdHd2iU2tCGB7ruH03BAp4xuNfm
J/0brlD0ZBeSVsRl1Lfuq1EnN8yvBdtp6R7Hv4UaKin/vfm1g1OuNZYwrAFgegmz
2sLBO7PpaHCG+OIynZAyS1Oxt2ELPUqaL+SBDHd8DMrhzr/2GBU3gZzhCnR4WiMu
KOhEWwgOnsDP9PiL21xMidX/Oc2VioMS7iAytmYAQ6ehwN1UeyOcMA1R0uy9PFW1
vpyOuYZqA/qRq3gvxTZZMSxhGFaIsjh98qLtjgdRob+cyQfdkutZh4Bgr2a87+on
Pro9xMnTCyUDRiL5NP6utoFYrMDC8h3dt2UzeQXjg4FeUn6JI8nVxt4NdFWuw0YE
xo8kJeUsyhU9fPszY04JvFRcZ6KLIxA/CmChGfY90biRuB6MXT03OgXMpqQhbbZh
W4aGeN3oqoGjrQ1vrTmnWoeMuEVT2OsJye5swkmtz1YGKRhiEXf9f/da64lePd5b
tXijd8z75XkOYT8YpkWVorl/k6u6f3nD4JuesnhQRI6KsORiEQTSHdoU53Vtct1e
gomrLGe3a5CwBHfY0ws131evYmsbN0renefxX8d8uL9hFn4kUMQ0tpMQzkRXSb+J
aiGGFds9oCK++uDzhEX4XDGuTnWazQlRH3s1eo2nBqZSmJd2Eh/5BgRBd3QVvypj
u/bb+GEBvOFrwZu69mgWLbQQShR1PXMuo3po5dnygItt4+F823ukOgsA9WTjwk42
svRLIZwjEYSgflwpAB/1Vy2J5qbdQvTvPNJBRTCrcJehFrQRsJlnidpIbsIuYJzv
GhkHEvWPpsDni6A5Vj8GOruiNxv0yeqG38aLGK3j+6JewptCVgzTWnClMngG/iTs
E7+7VjUD5A0keoiHSvCFBDyrBOfIb+cdZAIv1cI5PdOnrp0b3lNjT/Zi64clZRu6
0Z4sCROBbeJw5xL4YRq2oo1B9zyzoadqyT37GxDXQsgyktUAwXEYC2YrThyb65XN
EvW1UEsriHpB8/xhUdFzBHT+Wk7znDtEso9XCv61MpAvN1H5K+3icSUUhS7XlaUa
XB2YR7VOifUAA1peRQx5SDvGlt3Vnx6HlOmA7zSwUFiU3LLvf8ht7u2NA9XcBUdu
GERHKTn/5iTgQh0Z24Ll9oQAJUzqKTmUqYGFZTPNpKdhjnXgSQ4LzgAtaXOUCOli
G8qqzl9BB0CmpRyBDQJSqb63V1HekpiZ05QrHoS7ghMHx4XGx0fVs++v33v+SzLu
h1+A2O9jPbRzXcI6A2+OiqvcAeHAFnvTwkDJST14IbyWztFTOzT10WWF8gZC/tdi
zRL5FoL2ffkot5LHdTxvYHqhkazyKc55fbQ85SUK8AXNFDsM92sL3gXGJwi5BQJK
/hJeqIi+HXlyVBQr5EJyHc6qGGwU6DYLzhgnprRLsnRW9OI7AsWXhf7CKw10ImEB
rfOxUsI4i4MvkJpU1D/7QLFzFJa4tWc1Q2WYXqdBBcbJWjVccQtQuBALXO77zVbu
IzDQHHAX5A35j9sAmVYBPYGlL4a9fCmTQsqZLpU+2t3u8Iej+VSYK/EjB/QpyIjH
5XZl66kGS5+nToo3jAoP5KtvE9mAfpMESM1xwYjbl+hiHSDLZ2f/47v+JTaTkpIs
wB8avQ/zArVdSMdTTwQNLNWHCCQTqfKH7qHK3pRo5iMsWsYoSSM1MhmvjAUV6M6o
FbCYyXk3hT0BzxWLiTMZDM8vGbNfGvLYVqM+HtM/U9ru/pGpDL2wnbtewcU8OMJF
+BfiD/x67MhSgoWKb+st+jCE2eUK+FLc3s08wyrK1N2ft4abTy3DZK/XEi0s3wKv
7VWgE/+yMZ3gAuL07OtF02CWBYcXvuGNTAFxMLXUi+yYWtnefO7dDF5Zo0WOKqXS
QWsr+i4N0/3InMV1zuoP2ZWCRP7evTsI2Mh7JM4HcE7RkREp7mpvaFMJDzuR5FHw
qeT9kryn6ARsuKj3a3VJMLwW5pGTsEogahPeqAquPIeXLkJXLf0CcO8NLiDdoFcB
JzFPXMCRVdpaSBlikUsJzEhrxG/ZapTP030s1DK0+FMWZcVsZHwK7yrbEUCwXSEB
VJJqc9DxbbicjY+4Df/ZIW7L96NUCtcTEIHh2oN7hcpy7HvAKEk+KTNBZ7n5yidR
/eNB5v+Qp13aKZSZ+TnMkfeIV3TdT2ddKw/a+EkwhIUXsDqA5cR3EI/IN0Z8EL//
cpcC6Iu6mj3J5aq7D5ig0BTjkOnJdzHqsfyDQ1m1O7iTe2SQYLupo6wrvn6ixb0F
l7HAPpa9KxMvTkWQ1mpwP7sjUHljU+ZbDWC7RarOernFWsHhTK7JgJDgBLwnjblQ
13112xiYzOp9u3DDLIYheDqkxjCW2r3uYy7q6ryjDIxdPhstxlHdkS+iwmaPGZ7P
aLOLV4+de9vkxi1u30H7sqMYHzz1gXICZfiSdxOAgroc7zuDDUdX4q/ohFLtjtfP
N8EhfWPduoYm3O1/MUimZFD6zRGAsS6AfcY3xPituTWYowaLpTzzYlb6HT9GdxrW
t7jRYnEraYK/iBZFN2OvEHgeZ6XOvMuBJjEqoSnnYITNvE9XmL0V3+3QoqbRpoz5
ZuXBhJXOWOM2EAlBffo9N+bgMJxMM19CeroEe9QeV1I7qAIsbuNVbMCum9ZK2lI5
/KdfmtVd3oxd7P5LvnNTFpmg0coaqpmMqH9WsJqrYPx3hkZBvJRizor3KKJcmgTu
b4ifHz0Zr9I/LFKHVONb3rsueOIBW1KUcYv/D+c2ebVXDbWWTc0SwJ/4alHojBvI
isJ3SFta5H7Pnvr1LqsQw/DGOIN7Xwk3zbiPao4SXrqMiLVM8TaHekyG+jC1B112
Kpd5pIevtRBD+WXgp3Oh5cjIS6VsIa+tVUXbxgN0tCeeI7OdRhNDVlPfNG/iK5df
iMM3pThdBFwTgvXbzXnpclYfy1J3RhI0g4tbU3/pW2akPGm0k7GfOtVFPPy6tQl6
gZsdFuea/tjrS8LiXUut6LN+3BJigIGC443CReoFXX9JLBuebI0ku7bO7Z+Nhe0k
zOLVtv9yvTM9eEhg/pbKJvlGxn/3h41MO4CoTKemmGZUvU9enpyk5Kl91ZSaTsvf
R71kKEEJLooj6eSfyFGRFUBQ7sdugbP73f5tda51wWJukIG3v+WTzycAmXws5dii
eYGN5MZYv+3EPGLbo2Z/zJMJ4Hu73V10FX+qWYqkij/aHUa5sEIqMpHbd+YCC1/M
ANDa1kOzVWROiETKaOxBgSDGBAAmMnnaCL+nu+zbxNDEs3qXxvtMNjp4XLlZjsMU
3BB86Dv3JubAtdaSk/0GIzEOB4WILn3cGvBI6ElW/fNOPYV322bQOuAH/G76R4hh
1cTmql4krB/dnSo9jO9LNNHnbvbgURJ/IrtUdN4Za2aPx7yL0kuVbtUqgY1eUKEq
PMGhzY8UVrtO5as7c8Y9+5lOvQcJO3AgDINHemIGhSjRJVp1JdDuNEdLksBOCQhx
NL1Ey5MZGUd+clPUBn+GvG8MdRn0ICeGXr0FHFtrM2X+x/dI//amJNMA6A6txDvK
Ay+LD3KYpAdbL1nw7Re9nWCrKE0jEUZHkdyTIbctCgz5S38PWCAfv8epHt/84p3E
BatK8+M5YQUl9MtC5LcMXr7gbDhS8spIxnEtLE36z6CHREGfZkK9Ve8L+uB+KB/0
xMWMJCvyIIWaVa9Ernu/w2EPjPoxRo4Lvi8KZ8rqw3gehyPI+2oeADFqlCWZ2tDG
DztrEF3ziQuptzJb3pPkQDtzqh650OyRCsbqgFaL4Mmv238sPza3N5LAWSg6mW6M
tBOYKbihenbiALOOD0R8XzaKJhOyW8qQNnB8DD+nJ2zhHcKLFAyuXxRPDkIHydGQ
GhAVe22VKN5UErwYzAyPbk+odyqlN+mRmJAFTJfHA/6caY4FaXZaVo/QfagcnFVn
F7y3myrct/FmHohlRmpu7bh61hAzbQ+aZh0hvqPJgpwA+w1TmhnAeevkiSvS4Z3U
pgxO0cOby9nhAq/l+aVNNO9V8zyNYtWymECgvW1t941qRJfYQS0Lgtx5cXfWFuUG
rmvrsDD7WCKCMUUXSZoNx//5PWmU5KhnUsPSD5aBcwMPTMB2mZzUHQ3tzj9GUyU5
Q907eQE4e3BzqAwG0d9+HBDRX0h9qsQlPv75PfblW4R9TM+jNvHArdTbdNOKlLZZ
rS/HT7rRZBc7lC4FBU9Y4HFsyFNstNhN7dLiwPKDWFZB7TDyo9Tdz5bH/seQZV3Q
nWAGN1ezk0j5BTBk8fIrAecYPxgQ4wjR8oFR0VpZjGnLXnWYK1VPQYdmY82xBOOC
Na9Veu16jPZyxG1O3tmBDN3k9cg3FI0t3KAgCuB0Hqq0jLBHqaLMqmVwwtbBJW5G
NE59HLV60JmK7+9OrVWNH2iVuAWORFi1ou6gKYFp/nih0bhV7dnkthwpHH/zS8e0
d7M2S6OjOEwfE3mLJr/BVP3lHYxLuGW+yxXMuB7TZ4mtdgmUDv/0iG2pkd/gage3
906DHzE3KpFRZT6BDDKIZ24NUDvqElBybQ66qUPenMwgZmShg6o5T0fTHhDniawS
6Z80v9TuCq8qxnYi9KdRdOIk44/ukNwoX+Ymm3FbazBr2e5NV2uTrgkm5BxXhQH8
4fG42Gt0SzKR93NEP7hrIVVrA8fftYayJ5mQ+mZ7knH2B51L2TGptfqH2EFBGt+r
RN2Gd3gBApE5NaY8RsI+k1uI63HBybWCY1M9n0dd1DJiqiISx/0KSIuadfcwdgqy
zt9nLfx1Hl2N8JwHSy85kXtsAokshoYadRxllh6K+1337dvC45CwC2rDu/v+07F+
nAU1n8qo2Ie4zjPz0/a7l7HfZApLBqwnudqUG6qcx6LjXVGbaZ/FHB9kXQGTEYWM
dzwddrtWI/UkZj8NHpsOsOHyC3j9glCckco4x+amCEPolDKZg1cOeRGWMIuCWckV
jLRxALfh6An+VnRCdhpZM/Il9zxptVsztry37OuEv5wTe1uitjMnzupe8s1DslBY
LSEIwTOnq1rW4NIrLc8V79ewqj5OaOxF8oY/RTtnyQ94dXRfc3PVaiQ9udjj38hC
VwabSHdxEhvjLCMtPw5Rxmh8Lm9T9z4KA/NlNsFNJ09zob+GuqR7JsZ9ZFjFs4tw
znaNvnAvWMNubhZh1E7s4K2MQrdFVPH+q/AfQ1rggkMj9MQoyNSKTrFky3Pt5k42
HG9SrQBh/P6srvdBas7ExWzN4aukgrWKdtUYEFl3J5ElZDF42CNMtIWMSQ9GXdSh
2whdfyKg0QCAeBDg8+0vF3ISGeVfZgux0l4W3KeV6XcyJ9Bf0Bdl7YSGDk88e02A
b5LG8CZsgsat/N0gQINLmTM98HUr7/qnANeBxpa5x9zrE9zJPAzug+7Bf9Xwtp08
w3+WAMgA6d/PzvU/dF0rJRKXpG1s3Prb/3YO72Wk4eJc+k0y14czcYMg4+7SUgl6
nIYGxnclkIc36G0urEMs5eTgx30sSmP26KjtJQVDbZjDR3QqDc7uEg3UaQY5sViV
XEzD/09flNMnajNq4ESQM1SCV716zUdOI4xfHS2Fa+oZT5dow3Y/90dPa0rCO6Fa
qzq2i6XC2ADYGdxa2pORw1ZzmvSx/hxt/6aptVnOHdKZrOt+g+kXaaq2cp6olbSk
xIWZje3oZvyY9A+ZolRmA0xXWq5ymbCV6n3zh1qE5/xobEXZW5qdy7p0fosBITYQ
85zuiXAXXmuDKdX4lE7/A6jfetQ4fo3zAS9UtglIX5EQc4YRCeqB9o5USKdGCY09
c5rZ+BHvuHgLVZjX3X1+F/GonJISvRLHOScS87bvt9u24ttavhT8GuAphjcLpoIC
kPps8Q4+uJWCivzKL+1pmu+Zs4my/VX4FdX1D5pK6gelZhu88JCsWg4Ujs3EVwIO
nxeAO/6Gca13hEU5QG7bUpECwrRjVjDjakNXx5+vIafh+zeR95azBI2SzVjuVYXT
YxmG09SK7LAAO3gBad3ig1fnW3Gw8O/kFb+H4pOL4L+NjeE/eFrL11QJ+42zfBSf
A1+WUnpLg39R9Hhj9LwNxFxVx1ujrSPXyk9X20t6c1G071oB7Vo1FFa41LHcmyQ6
YhlJDI9gy4ihPSZxLgNJ1+gMaXaAHMC+vSO11+wUy51qRJskIObqA13+64AvWLjP
Bx/EjQAZ98FcKGb+G4yz5rDUT/XB1MbjFUY6iZPwFXXrGUlhV4p9d13bZK8lJ0I1
DrzSeJZjGyprx7hCHa0yNgsQloMpbg/4SizXX8u1cKReT5cw2mXsd7qG/SWgdZ4E
0Ghef4HXLur3l0d3JRTQjarEglR8RjhCEl1ytoH/P7uFwG/XU21smEZ2Pw0cuWUJ
Rc8zAzIjNPBApfv00XZnmetJUyakfRpYP/F/SWKmPJL6XRjdGscDwfihU0iXSAfQ
BEk2hoV/9eSwmL+hs8/WWU56TxIgjMOuAZULOHqVed9lbHdCqPyyU0WHRIDPVK2P
wk6TF/nypin5mYgMV3GadFDJAizThCWBf4bvoHZcWa+ADICYbILjUQ6FX72Ncy/u
Q5RfAlVWWrXKd/BBeLCfShE4Qs3Y9BMU71vc+4uteYXuQy07VUNBTHM6QnAN6g7P
CmvTR4esGp+jw6SvXQeQyYiOTwI/1Oi3n23zPqoT0AMG8lVxGMGqnfYi0SYtFwlE
DrJIhJRunaNpBgonAwwx6CbSr6Yjb1GOm+QF2PEhAi23+ccqQDaso0We/bXHiFhf
6zVKlsXufIFBaxG3ODzgVyxeEVNtmj0zr624hOQgoSIUliF0UfGdh9mkxWiFE7d6
+HE1Lfrp+i+JQekgWTVDCWgaQdEXkQGi8GLghOOZK12BrAnDJc+sWclWYE/IVxxz
EF667nM1oHZCrIEYt0AjUBZv8wh4pzxwHAXa6h1d8HVnJIVf2VQFF4S9/EchZ8ov
CA0ZSyZtr4cGRnfbiMNbzUqOOLIg82oFZ9ayQtqaI8uu1mHY0Dca9hQZopDuKjqn
wYDIxg88xPaM+jgke551oKq0lb/kbVhUOpUkNBHqXsp++4q89/TrB3bUCpeDNu39
tGSoCK0XGFIBhZCS674CujHgwRO1671pk5VLsVUZVysJr7+uT4NwSOpdlpXKm2m6
sB1AYTm1YwsdewsprdUrjv/7wBVTuRitNzOV7Rqk+0w8m9HXcxExXmoMOdobjPnD
J54FcWhCZiEQp2FBCr5qX2tm3mb6jcgddkFxcUmJbX8aiAE+9Jlziak5DnhID6i9
4C1S0RpMMZUUPDd8EN016ri0EHJfX1jbfAi23OsgDw3PfuAmoOajED9QjB0qESDY
kCdZ4cffy/584AzT/5X/vLM29H8PfCfNBfbfDdeM1ZD2aNig1tfUyuDOrgZ22s3t
Uh+w5thgIkE8wbeINsejcVeDqodEAd/VAgLbfgVSfPFHJ0L2mNCh9S0mWnUKX6H4
M0LGd+96Fqjkht5smZm2Co96FwOb/dkYH2M+88vUGA5TxeIYvifsjL7RJvLU7J/S
BVj08Gx6mbeX8pczQbp2jWBIYTr9o3OEpHS0uAGaasZDywWbX81Um43jzanC9c7k
H8/lHYXFNd5VbB2O13naarYsAkpD2IiKJA7k8JLF00GF0sZYY1al8GCBSBRWqzAk
gsolWfoJkCEDdPu0+eC9qGxlxpgHDj89fCwxYX0RzZPmaTmn4BNNJ2Om1mv6FQUn
VaqZptPYNRcsdy6ZHONkZwBD9oJvb34FjzejDywVmUYG4xwZFGVDGozkK07l9zxI
MAy9qZHU4ranA8eJ4aRPKQeuqviLFE3eewr78n8VKkuUSuBuCocGcyx+XyDKQVci
ByqgYxw8LZ9R1gXmIeM8KJrWp48y40vJjLzjmWc1TYG9dC7BpDwKmjUWgRO2TIrs
rSamInznjI+FaznhCuvLs6YIkvFg6o+8aGPqU9OIPtX5BMFP5dIT5epxHsuby79N
o2iF/guvJ267uTEn/g6BQe3gGvlm7ieWzXT72LoW2kuS7SXrwiuud7MIj2CgWxnA
05r3wQ9hpPG1XYu3K8Zl6wMW8YgiXo33Rd5gRBuTff+RaxGQ+ATMMX7KyNT7y0UG
ixTh0GbqflX3xrOL19nrftJBZ9Z//nSPx1EgjTabHiMadCJCLlUOI696O5Rrz43K
Lcc1Xb3rRaizJ3VAsrGLAl/TK09Qja/JumBGXKULZzqSkEprHcSRf7WJq7YcUqUb
HFN+5GcASJxZ0rEJSLfjcVghhYzS6TAmg2FSk/6z1s+MRIgp+xJjVw8Zg0g2RZEN
T/JydjOzc5rxr3s16YrKkXJ2x0wJaStSyqOud7wAXTUQ70u5f1Cv89MYhq75Szr4
s7dWX33ch/LOCq2SwbOKpLnJBC61eWw4f3EojEIZKoZipxDny7in0qkP/iHzb9ZJ
gfb7801e0r/vT1MKkybKKUiXaTamRB6/v7S3cciDbFf4uo9SsiElBLRMrCbvpKYJ
ycdZp55uclGi4Go2UAVFnfoYLBu887Zu7r+SQkqFEisb6T+w7bF3cykiywUmCpDc
fhhHnwboWUkz1kKrQd7cACNzOg+I1TTUECoWKpc1sPpq9Rn/Bbcab+YXS1MEuo05
ctDeAh/iqwClEWnIcMova4ZHsTD13XKVayX34DgmFbujP9SVF7IND3SNl3X15mUc
82FXJVja4hGvKK0lYXve7+VFye3YIyFb/ry/EiTiB3dLRerYhpUbZBGt/5VzIKOm
gLFIYFGm6tFyvVLyV/92IVNZPbpunp3trdTwpoyWr6QRjuMzSOpTeqEJX4xHcAoK
CfCC/WWGUuddoCef8MPDVQ==
`pragma protect end_protected
