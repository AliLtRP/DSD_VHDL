// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:16 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NuHzxCsrul0zvbUIpNM4jOIymTQctXMa3U9a2wI/2O/M+T9eLz1Kr7mKKO6d3I7h
XXjQZ0oWc6gH7bvWWn1CXQmkzN8mSQACdMOiZoB5VeRncAYLmpOI93ZJlCyFTBuC
XUSxQCuIxt6wbrdHW7dtGj6BOpkEXONyQgRh9k6zPZo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6960)
fH/9gZl7z3POgJvKodjsV61En8jge3L0cyh0M2t+c0eSs8n02Huyc0iR5+VR461e
xZfMPnf+TQyB0RqkzsshTi+TM/qTQSjdXAAaFWDnx1u2Fcj+oEUqpGfWYsxK+lcQ
p1S3Hao7t3GhY5IxdrjEGrVjPjD6IXkBXR4XznoUZkiQGHXyj0cQhst/IhSwlpKT
S7xAOO+NfoepG9bxy+EvO8EYPunjctA7j4cq8vAVlHfsxPgvzNPj1vQpkVyze2Jn
RwU9wqJ33FeAEeXCIYU/3z4sZd6nZgQuHp1MaardNtrZWHSZ5nEZ5OO4okdHH58G
zgM2SXW/rVP4klC6Ak9tx4i42iVJ7jtC/JRzZ8AfdW4CG7ab/TfFwz4r8WS3iP97
ZxWoFnRGRNqHL+7bVvVcCUGE7sj9KMG4y7SCNw2ppHpQV55waSNFhhKDogRtU2mC
NzTmzg1CW3GIIToipmBXiCl4s0uSswjgDW8rj3ezoXJ8NQMEULzk/IISw8u9jZL3
WFEAkrzx28wcjjqHCX4kguguRmsqe1uLwSpVq8Bug7MJGKvI9kovtgDHYFprXQqR
ht0hXHDe/6ef2QzMKYliPQnP9biSfeaOhXR8mpReeIkqh61rq2cJUBwQXZhT6xhR
QkDDjCl8yRMHQvGiToxheJCRBsXa8ET7AJ2zqOgtmLkKjqQRpbZTAsoQrocB3AF2
qmMh3kfYuEUwECRe6Kzi5588iKDkeO5AfYfm40vlxzvs/4zTICkkw7aOkLdD7j//
R/FhMgd0t1U0TSDCCo0dyBK9kjrRCLVXFYD3zW15Jf/lrwdQ5F99et5jKzX/oyln
YfxzRR57ch1xmJOMV2fsGmMg54unyfsBTy8yRqNCecgDRrivUVcv94AXlliig4j1
jBmTPfdYQml66qfd2Euus0mUuKcTHI4OA3qRBeTSdRMKvpz5jXxVj31DKocgaZoK
+zK6//TweKdkGBrhgbRgXo0Gmk2rKUanB/XIGKXXHKwYE042ypZKBLHuq2nsgAkc
z0f8HxdnCvTppYJ/kVzI+OV5UxR6/rwLoco4dI06CwZugOnvVSs2JsuU5oGYP/mk
Jz8DUO5OJ/CnIXGyMv1PW+DRBQIm6kc8Adm6Cc9FRWF7VDWZpRH0AWxAHgkpa1Vj
b66QFtjD4swBW7W4XHVzqqI8NJdoFiraygrO4YXmOcbSx7J7n7jgDRFa1qoiMuxs
zO0qx04A/JmYaK2JmYbLBMA5VwI4nPGY3wgwXLGTGAI1Mmz5kGQGn8rJNsRHFORw
LPQ/3O3PdZ/3fF1RCkte0uByD6eFZxE/44YAZCyxxyk5NUZaGkNP3+X/4v+Scpw9
rVXC8mjfI73l5LASJboDntwtuxLg3qq7u5H8CYlVIQjEUiAT7gr1KPpK5mo+YdOv
WdD/azCtCfobE3nwEUT5n1ynmyLdzSB6G1UIwTlt1LOrAIgQ7gvZnkbRyai7P0TG
sxan8f5JW9B4gCIUc5lKYcK3aIbp9dQeN25pcf3HrELN+RTyNgxOjnb/keWbA+Sv
sSHRSW9V67hwSgBff1LsJGrSUn0NMTNCZKVn0cnJDanTawgyPf8/vSScrt6e4kmq
GidxGxJvHiFu3ChBv6IIN3N2rB5lcwROBTe1FuQp1rScdEcPL6RiNABFPxl1/JyL
M3UMC8GM3zpm/yJgdrFUaJsFBG/BvoiuBIcC75TijP1ame33FwtJqhr5wCPZHrxP
akg6uX+78jm4TYEEfgNG91lBkWDPzskLDnfb9CEmc464CM6ktvZhcy+hgcdM/VSn
G2p+KVktyOvGHXrjtfn0BgRE66n8vPiB5TPCHp/X5f+0X09iSizxcdhcC2oydP/t
RMVLb2t6n7d9E8ADOXbRy7RyROUOG3lgaNFHPLJ8O2RBzsMUO4V5Ma8Pen60QGvU
/d2JUZfS+NbUwRhMP8H6V+GlxPzZbsYoWj+kmZ37ppos8Rv12OCr2hAXhHRAdKyh
wXCFpZM5n81zcI3Kx5MUzdMjv8OwnhQOWIccfde58ajGz2IQMGan6kCBY9nkuhMq
WygWb1xz6K66tmlheEvSA/i1nh/MbNiWZQbBOe+/07wWGY85w+P7IPkyfOmFifN1
UfeAi9koyuJsJqOGn6Yan1Qb7NytpSW2tDtn4Q1QvLM+nURLapMqIY/MzK0tjCDD
Tri2NeRRCAgYoAqwS0oOFt8UCZpuY/OSUVFXuHgdxmUuQonV3J33zz5uGVufcarO
zP85A4DBpb8y8MiaZ9REDnfgGNBNT7W2yNzHvzRd6xswcQ8wm31eiwPU/QBlMMI0
uUsPshkUlyD9bEiP/6B0AdIhhoTSdIu1c2De4ESaMuHw4OsH6hhPRtfNqPNtX4eR
5TEcHnHc6C2m7lI4xjlxbphJAA+TZ76ojQqGJXgFuS5Ho77QmHJCGdQg99HGfBoG
41ByNCf4AwTOBotctaviwEubyyrvYwqOFRqgbjIuqEWQzrIG3fnX5u8zWv2T9MlN
oda5tNsy0iNzw3DV7VkOD3zOQ0l8o9L/RWAKPMuFaxA8iwgJE+1GePxhZYwDPWTX
MOgR/ZrPFu3WnFxgLcP199EYqHNy9hw3PxJ99etscWu/Zr8k88Uwv0LSzNH+Ztrp
2uygTgrZfMX3DXvXVY+nxFWzOYCtZfkrF5QRGG7QjDm6LwHwjTgrUA8tWjvWk0hB
89OAIrpqsOtBJL7EbvNOLrAIskFGyx439U8QEJodNLt+Kl3iu9Hoxjc6qyLfzh7R
T+54Jh6FPw0us1pGiLLgU1rwyPcLGqWFXLYX5oEqCV3JosR2PbxEaYKB/vuXdlD2
7B9BiWI0u/sGWh+n1nFCerKfLJwIkBYutH4LcKryr7FhW521KLUl3e9/mKV3gU4C
969NF5LEQX03lBirY/vNpKpNXxAdcT1vQMsdazDrV7Nk4hVaD/UXfZPmJrUeiKUg
vEcj6RhO/kqm0JQymZmtg/mzy3ztgYBuFRSXE2SZ8Nn0ZSfEnSkKJm58KT1Wj6XE
XK4R+Xhf80eeK5W3H6UUitT3ObgWMCymv2V/PRwRPIKLFTwb21n1pdDeXSFgntDC
XoBnRA7KeJWE7rO3gkqlpUk9zBpOcQosM1V5qR22mCxHo3aOCyEVVitKve4ktCs8
qzRpfRrvUpwKKVq/NKCxFbjRAqu5Tm4rWWPDApTPBS7RMx650QAAqh/9cn29rlol
cnIYnAcDeP2IkiRdMZLS8pCK9QNHiG6hTa4/+wnhTDBDB21P2yxjn+A1rLW/r/4+
tOV82R6RcaAOJeB1Re8wx1zlIJuuMm7UvDxq6kLqvN7b9H5DOJdi75XU4WiTvEJo
79p4APV55KLWASCPUtkgb0WDrM5w9emo3o2Xh7DLdaRjuQfo2QG2RSmpqWOfb/d6
FfUa9aYshcSMEc0SXDWjCknyTI2KqY9MdohR6hummLnE/f+l//HCzeP0Hjz6kQZT
4woC8mXk5VXWnEc5RJ0Yxk/dMx1CBVp9dX4gMXyIS/3c4Ne1mJGUVjE9YrfyKEpD
bKEVBxaxQcWNUQI+lCC0nP+i9lES+4yjYSSsEbD+lSzN9L+Gn7RWfCWO0eggqhsd
FIvNx0KiZepho52xqL7cO4z8UegI+gpJiRqT8MwITVSZdPdeJYwYARggZWBtbRjr
rWdjAGJFbUhuFPyQGkkuN5JcLW0/uH6Ss+g2YGi9eKDJWTM/oAv3jHBeEUnlcuxs
49up4qFmQUC8KKl+b4iYYbcDJ+Z48vSD8E7QdKsmiZMbLXxjBxyYaZQNN+NxShr8
oBo5wxsXK0KaB+Uwr5bxgC3QJBELDRa5qxosqaRptUII1sa+BHerPV88zRLD5xrm
zKWeVqJYJqpt5bTjf88EKhQfIh/vqZDGddD3L8GkyH80AVS4kC/f/V4eI/6VvKOO
UNeQ8G6zgJq7X8bYn0nN9ob/xj/6SZ9lZ2Hr4vpTLfD00X7YL9fKepQyh0M5XFVN
RJ2o2DlMx4rgNApzXu5zIOv0iBXG19rge38MSjz7h4Rr7Ko5qk5TNKTDCaXDJYk0
h9i5WP/m5beFYSi3fhbAe1nFiFKifUM3qVd/NCOj+4NegPPcRMqEvaf7WU1D+Mpt
YmXONxE81xZjNmj+efKYnnAC4sxe7r14F6DvDBwXxlSK/jcOEQ0YiOY/6/oCf6xV
ZELOYC6UOKVdBm16JIKm2iQtMCUkszORJNjVzT15FuKl+I0btMxvIroYBUwjHk5R
heHwjGS//R3zkLHMw9oWIaunUUFAnacfNgqIfcV9HmPuUyECLmyjvw2JK4jrF7Py
ipkslcKLUrLx2Ti0rWmTvmfWN185MpsD/ReiNKuWJHK5x3YW+W4SFoLqjM85kStp
73ZzLB+ydky/Z4X+3pO0ylYxwrEhBYoreQ8nu+KTkKFxBW07OJYE298Jej2QQpw9
yiZ+YSRQ9o9vbtdnN3aGInQh3HiDyX9NRurw8Ak9sOeE2YfbWP/ikxlW5AWMnLfm
tlj6VW0TqdgQ7a4nZqq+jAVE9KTEhD3lO7PsTwfsmBIO9hefwMGxgnCiVrdm3xLf
GcMFf0e4ObD9Gy86OaHIC/JDb1TLSl22ZU8NCGJrCq1YV2lQleaDTUHfjysWT32n
+SmMKl3JXjzru19v/3oW7sSEfgCJIf2+1P3XRdGTuSWiVzreH6cP/3IYpAzcPpDq
2rfw3/NzvWPsO+DUqlnkZDpM1cQTv66I6obhCYXavduFdyxfdwJ2WABEcw0e5z1Q
CD3rpHJje0ouRMnvz4hzP8n733T5y3oZdmbB7WaJxBFc3MRQxNmh8ZFNifibVlk4
JrNITBgzTvgNamOclDTrFEaSd17zV74pwknCQ/9QyH903Tew1LNMusAnjgWPthwr
JBGzq/m/8tcSrvf9uF0BBxIugdAY5FuUrd32HkyMIMArJ0LnTZOlZ87dX3gP1TF8
LX+XMMs4F8uoCx04v9Q2ABlcirOOq0jwcPs0Qm6t9XU8BVwVDauZtLlsMSMX2auC
HGOODbgs3qD1Re8AGOVBpVCFXWvad3VidnqZhsoCdZZJS26QT8Lhh/g5EIql1LmH
rlwiXsY5yKG1Lj3eOKi0NcvSiQBNmSAbxiq3BocvAwm6NuBkYbn8FuijgQbt1QSm
ezeQXzTwLrQ+uKM4cucJvpjECHidQvcUc9DWaRWbhvVvuVCAnfxxOKYV1DO/gqIn
ymYLyMXlP/DYcDjcDt29LB0MjAgIUz88+9gYSMr04nkPXzY+fRmafazNv9EVZELx
hQpQH+lNNOCEr4+7iipvN1UE8itEyioT5BgP7+3VT06skFPb1dPT0+EgKQEathO7
rQGYL9ZafGp05Rh1Nfi/hrDuv7UlCyinkHQzs0m3QJEyEmntuxVEr+rv4H4LEYty
BJX7VLIzWooPSp2WAQYql1Rt/f5qfi04TFPw5KWiD8MzEqc7xvjF0AxLzuDIYkeV
YoerJCIFK3SGn/pXIc3OkmM7Ds4EibKnCA8NVtKURHCjbEWWFEBCWuMt5fQMyv15
5Zq5EsUpVKEwdjMgCwq/LpnMqAdVuLo9uE0n3omulQm/kXVJz4io15nc4cPsshXc
feJu34XkCp3i36YAVu6CIEkKB1W/0VANUyWklTqBvyklztrUDTpcnVOElPPLq2fY
bpk+l02tXJRVIjiF/JRPmph6aoB6uwub3YbQPiXiASMY7jkR8ag6fbZgMnJ+08SE
33epvW4ro0BxeHM9eW5A1jihZ2zDVkNQmuZ0ogF2dd7nagNuVHc+U3Z3zZdn78Cl
9BHodex+1Khif+oB0c2mKfiPDkIniX2jb5olEvQmSzzruFltyAs30EQJETArUs38
CtaT98dO7D6e4tEqM4CO35+3d9nxic3UGx27hUQFO9rU8KfLGRnNUpfRCZh7LWdK
NfJVbxdDKlH/lJl+0mLBsYaTGJo6f1TmjAGHm6Wj4T7bGm2xZRRISk4cg4mg4gBZ
2YVQSrxvkCYYiz1n6W5Wzr0UUghQUNAZItSCXc4CYuatSb0sg059VRkymb422T/3
LLna12Ez71B4LNjOuh+5jl11tIQV/fxQH9UQa1mDZBgaOq50ZOhBtZ7bigUBKjPg
/Aw6XNdMA7qyfdPeYiODiFNg2lzou+T1B8YsCgrZbN3JhTtNbmsGnKeFxkDeUFWg
wPmR1idG181M6S/t2+JpSl/x9TiH5hChGVpZfWQjByDnrH4NfVlHjNe50HIaOa1x
pMN0DC8EPKyIRESP7i4yTu5dM2bF0XOPULOBQD+nEwGyQ/x+X6VmidZ0ooP58Zaa
9DaTtx2Q+KpR88HhTTwjk4h1Cv5P3fozaRH1rb09a9Kb4NreZ2hPQkvL29ySxzR3
0cXESX+O3VU8YL67eRhtaPOyAdOnlpER2C94V2YjnFtBDujIBBNOFI/d3m6T5kEb
BsVZ9xUPzf01WsEuC+2bJDSiBYW2SeMjVhsBXaH9b1ryHpYMw9C01dxVxvxIdQ69
NW02yoWgXc+ILjGt3zy+YPwo9SYgTpRp4Hub77huCuQZgUWfV927H58+wVPXJaOC
eSDG3xS3+FmXg4wdY6UYu2FIB9FpAgoxnr41EUachN+Jffl6uYCpTmYuCbAqDvJb
SCUerOR/jTmN9FeE1PMtlmfWF1ssotN7VXQmhPle/u8CnnuXaGMmmioB6JYWu6rC
5YbfQR/gD4F4HgTWeoIKF/5+DUaLxLNOm3DAe5LKpXas5UbP7UrjY75aK+kpLOw0
DeGoas5CCGdNCvGh4mVUQe+if9Pw0W6SacEzDUksAaZOZYkXsrPGf2I9mIUz68wR
UN2//AT5mqFAtOWQc+Agc/UbwJ3lfEop0R86bFkGT7ZwYEFT2jgevVzzXmpAGPOx
Gs+bJUHZX7zi2qAIKYUTRbuGE3eFt+zwrI93ZN3nb/Mu+w08JFowEGr1S8+3vKzZ
ffEKecNm1Az4M2HgWQvsVoRBlT5Wnc7xGb/vWrO0Fs2sTXIPHPfavtAZsJPtWhNi
OTQ80444aQZ/hII0cshIVlEvLZkGs3cQOEC3y+IeCoNiOPllDT0YHIrfD1ljG35h
kYT0e6g1aXp6nKLD+qwl6WO6CtftIWqiEkrcLxDwAIAfa5QlYLxkSgrkcvYEIP2M
k3CKuU3jyuuM7IiqwGJvI6cLS4GYREf3B7dcX+iYPwkV8KFSEsoogrkLfdZMFHlB
UzkTJSi+8lEkZJlWO7BbLf4zEavubriD7PcnwCFOaIK6OtMaqfOYZUuj8gASRV/f
zq6M8rnW6eD4vumwvlK/8uZUM4pklo9Yo3mIaBY0dpRoz0ec98WsmyBK9zrvI0NW
Ad8JncoeESL+aXoJC8g4hXZ2CvtHI72OUfnrhy1oLqMIyqLaE0RTdvNE2stYures
v+cPhYygEyGCNLEw2IRxuXmzukJpimIg6iBw7Z5es4MRvaUf79FBgryqh9iNrD9y
IrHHo496sKfQ5PZznk/6INbc9elfbRWi/7wRuKonTeEMLEZYWZxDOEhnzPCFnamJ
Z777E2BSV86ykAcUKssrmFIF+esVwCeHFBi0BrA4mD82G0b5lNXBajx0AngW08Ko
0f7q/OaeTIHiI2IXmz4dP/8Tv5le1X25Qk9fmTYbvItg5jDbqY6WM86p+0cyblo4
n9f9EaihZuHIIKjVFB9vHRfe4nwgmpqjcemcfVbz3fNM0VsThP+Ci8I8+eLN/y5j
1Yf60/l22PPAKpDa8rdrSjbZzZpjoUEo5gsCXmofEG/rVwLZFdYTQJ/ufFRiKtZC
Uu4fHJxH91FqGV4Gsewoihht/K6xQCVWsxsxQLAlHyXv472wxmdEUeZx9z01awKw
MORUam/fjZgN7QQ6ZMQumtvtJ3tpwp3eVLPXMsH61dUs8uncAlqB6eksvNBczhM6
ucK0nmgMr/qcXgb77EI4txru7bn0X+H+BSiwbg1u4zwbx+dVCEbYS8ZSd2OEBFaO
2Thmwb48F9JSWoc3v5NtnvZUB3zgHCcTCfrBN4xQyuFbEQBR9cdR3jhLfrS6OIxH
LZVqw5Sh9g5JtZc9aK3E/GYS6q+nXV6Xqfqo0jbpvThhLIHsO2CjH3oHfKrusCKv
GuArydnbvruKReCkqOOyavpYn0HsnXXSoONUIz0mB9doULw6EH0cD6r1qZHeGK27
sYoSwESRHx9AN/PzlLMThCdHzNeI6w6EHOPuda1bz+b/N/nBIH7HCPqDhiP+P6W6
nINixLt2ahA9JkgYI6XTEQZ/q799dlEdzDMwtH/YWdo92zQs6o3jPGKqTWk98KEg
dZsJs/BO3r4No+8sKHtj3uJslhTUCEi8ZT11XtkTluC3oj9JNGo2oEkatLUJAQdf
KOvssUgrhblrqGBwPB/ONuhlICYCD4Nm/7kvMb4geptBFkQrSoZ8or2JLHZybVqf
ajuw5YLpooR5rxjne9BV+hJzY3FLP8JI6DOTpRerZFPfDWrkcKqb0vDUvO1Za9zs
RzOHPbVLzihCx8wRZP0ajdL/fa5zYqlJg5CN21mk1UBxjicjgLyLU4EhSIn4S7X8
X4YrcO1yoTIbFXOurjQjgeTGeo5X5Cdxf4C50dsiar8XusoGS//aJi8ktp59KZB/
7Q+VNMHStCKn0T33JsJxpJhq2KB6c26GJZBk4rqczppsenENjBs/eUijOGi8LI3y
GioNgKf4YmdLyXi6TWH1MBBpt/ZNZSZaPAWT4vUkNRrnIQPC6nO8PajJ/qE2lQ6k
2qiCIqFBOoFWKeeGK2R7+FhaF5pZswhnPCoBiYk229qKL99Wt7qirhmbQL+0rJ53
RKeWQiO2RuF3e7+8bEuNjCRp9+SVZJWNdhhMp2ToSE7F/9tyniJAP03B8hMuWsAx
O0Je45l4QfMjeqaAe/HBrNKGdQsginlm8i/EFkBqXHHSoD+wIzBfBiXiKxFD4pPd
gTnBYjqz6tdMjxNXN7YW7DZ8JeVI+iIcaG6uAOyzovv8P3Qz3M5PjAmrQTk+0gb/
OWlSlbikI74SP2vLE6hMYpbvZn5gRdrikiO/6vSPMPF+rINF8MS0ZAho2JGi9PTa
avbCIskep8AxQjwU5WETux5UZ/dBuHvBmG+liz5TMllKiVJYFGtH2mwYO4C4UYdJ
S5U8e+J22KdHXt4SCf80Rumf0QFmCSeWlj/juPGY+1cAKoG+aPQPMQw4zZQyIugK
hvYlRx05b0ihJGnrJlr8vcxPbk9Ybs8xHqN512fS9qcXFeydyoy/erqHaQhT2SvQ
8GlL7H+R+eOBy4jCqjJzDbcqvmg9PFJ67tvHpp2sRo2c140W776hbYNwID90SWPQ
`pragma protect end_protected
