// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Io87zRVumN6w9fVk5oG+7Q/Jq+XQU2/mBf1hK30a7fOV/g4337seybUZeE2dxNRl0bEN1Nk/7uqo
rZjlAdc4XdBPziyn7YJiP8MfBfIHLGuIpa5p5HEzpL2lsWyYTTurpplbSYFy4WNpTXIaPjM628g6
l+SYVpeskatEc/UCTCs3O8dB+GfD+OWME4HveTlW3Xi3qFeZq5exQvhYy7cDOdcltzS3fSCltgCJ
g+3u6MbNrxKNIGLnTQPZ0G57t3ACwoWr3Z8bvJEs4GELwMrERAFajMF5h6VjHidJSW+y/lEhY1LY
rxKoCmptyVxRE03GFr5441b2+8k1/WgfGBOSwQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
87T1Fng+QOHNqU5SCFxS7EEXNlifl2ZOq9RePhKM7P3api0TsKCAeMzNSyq5vKu5JFgycTI39TvU
Ej3/nj/1FR1vZ6VhXVGdYWjNOJEWiF9MYDOqQM3HaNL3aWKUa03wkQeEqUt3E4+6expfKriCrqHk
I+0KmniZzPmAZPkCzD7/9euLDBJT3bCe1SI5sod5UO2GladOGgt+toV85HrtyM5JmzKdNk+wC0vM
FtLumhA22khC4HIs/wXYRU8FpiCYgg6RwPq2n2fwNZ8DzZr8T/YrjziTr5LP4gMBiqGW8ptYr433
gVu1ZGaCNiCaCnjvCXwMsuSGDuD2Wn/mcb5H9g1LJL6qry7P5ONVPqfsOT8hHk7Q8PHJjsnrR0dT
aPsbuLFwUNAGsJxIP0UwBSOii2OzeSBrrssQriGkBRfcRocVNCsCQHsLBeWG5fAZhV38JiPh/4z8
ydjur5TsQjpdYFgBYFr+ygd55ChEMObz8tgWPbNEbg/tmc7RNkuF1Hgz9+eouSHvAn6Tl3MgA1PZ
4iPvmj51xfWlcwLUs2sJCwom8YWwCMr4y5+Dp/GK/hYWEoWSR8LQMkW+PfivehBBNJ7LYbxu/Wix
V7X2csFEZDxAqvfzJc37KhX3k5uYclvaKzxSd0ukJnF8f68jc662aBQiJ8WaRqgNj+4dZo7FheS9
jRrc7yZcMOh6ZBK0D+1FW5oBjUJmiWlTdgw/CO2r5Fz5l35Gz8LHDLt2+Q6Z7w4YO5fMNyUoeHA3
BpRpkzzEroCUT8xmUN23kYwb9zp7AFBdGZ/cESK6O91unpTNUBpDQDtKVdhnrHWbPogMa3+t0qAB
JpPmwCW/di2N89M+cqJo3TnjB2xxZc2hoBM92g7STDuXyEl1pedjXsiDhLVKsLy26DyJ7q6qk+p1
f7P8QAuh1jVzECXhmHvbAvoMoXVIIuARvgGZUhJmfYh+/z7alDf/LWVD+gquTqnR3MqnGfXDWg0D
C9lI5Vc/MeVSQPkKLcjS2ogD+oDvxMhRM3TF7wS8uThgFEX8hOBMYDrKEqRA2Z9lYy1gFs1Fx3DP
DIhOJ1TWa9XZHntsyYTfQVOS8qyA6GGeRvSDw+oWbPW7Ybyt7KwHyrq55wUUoRVeG0sxFF8UwHpt
l2X++d6n7Qv+GhpAfKEeQXIsRr8V2QUZukQE+8Fzd1Heab0n5f3aW9GlNuIwigv0DmFCKcP35hKD
czFnI5gri3NYZ/ooFzchGqC+mtbqFN4Ye2IOyUOQ4RKk/vpCSMw0pgB7Nu0Xoo/wjErj3GUCmkot
mguIaQjiFrQOmH6Z2Z5CangPxqoe9kf2rqxeOtjCgziKKafT58N3SRvheH36hSa8JfA3YmJTGn8U
6ddgl4n/EVmHcjQxeRYNJBZUSu6OpQAs71c3xnRFeXX6gEfof8aqYYJ/IjEnLiBrHOE7qrZu1GIb
P00vszdKxrTULWiFfV7qYrEdvatm2k3ffhf3QFFpVjmbBV4AT/kwzb6fhaZbHgB+yOp1IjsdmiT0
IZ29WoSct6he+VhsMG+bAIMeplpNXY4BEAU7kBl0OemGln60ZLX0O8AyCYX3oGUq61svwJwxQ/g/
yZvEtEwP7cDgghtI7QHU7ogVioq9r6kepu7/1LNZRGPgp1lU5+DCaz3YGdtrr47ho+wmrHXcpmZh
pSWCDznwMD4Wc+caDN9bgYYK5FoZRaow2MgeLUPKuB4abr/g5a/A3oaOjXPzmD5rVW05TwB3NYjx
rJXCPdUBCwsEr4/bNa49HbGlCG2lkWD7cLp84CKoYebxvLT9sVskzgq+Ihij8jGsx39pj/O8z62T
ijrGPtLcLAe5Z3lwtylL0b0nbqQiqRPiGBtcDaaEYzYP9t+hFTJquhDhaLfAbyDvBMb8N+oGqXjO
0xYUDL6M9RaH+TCh6NehiyDg3EqUAOPGXUbHRDDWtx3z4f9NqGb/8lIn7ImcwbWymmW7YDpIlLOl
IH08u+CopEWA/UQtD/uD3BR5g/NKi/ENko6gmGrH4LzOgEN7wmBH1FBRWccc/05kzOvzPfX92NTP
KDDQG6MBdQaPoUqBCE6LlBv3ecRH/NIfIayzMxwzTJtq9mQ6Hp5wgKpVSW+AFcrQ2tE72wkX/8JR
Z+AWpzmq83zOxbfvBMewQmbkpH/19sYLHrcSioQ6PrQ+4yL4xE9KXrI7TvQRGjsrxms1iXyFVdz2
L5/ESx0XPl9prXBn1fE6V6eM6PqpmhGeXBFhaHuA2WB6ukarJHY2rUsskC5+s5AOSmzYmLurZcDx
egUXZ//t4EkYBSbSoDpfIFUjDPijxrXLmea4gicyT9iFm954U6fbc4MRvvtGqIrlUBxEVORkiRjt
0eFDR8x+6jC+qXzA1nc6nIfv3gcRPL7LLIbfrC+80kLcBB1RJa3bT47vPYLJrV+wN43hkDmFculz
6wJh7t7snL75F8ZOApnJRFUUDafIxzx1Fx3ZC+zyre3qSoTJVIHb/6693HMjMBqTUNskwg12qzfS
+AycrpgxX2Zag1/sCTDy13jkZguuQg0NeenNz+6YxLsBt6gkwNqwci6ErYzcqxwO05BHzmWZH7it
PtVhadz6qq67jR5RlhUm7vnbx89cecxlyujiU7VacvT6oYRSbCVuZV27k6KkXO6t1j+KbQw6Vlg4
c4RCI0/ViZm97JYY6s6s/x7oM5pE1RNGWdzmleV6+s1Jx1cssuf8nz9DWQLiPvvO4R1Bsyvz12P4
4QDzG5bhLi3m8Si4qbIEptzaslGiSY7YjILYZG1lPOpkpF00/uOdJAV6hjp8ISIx+kiic7HNWj8Q
aAP+XGUiJx8p7HHd1GwFjRhtnbOu6/Hzr1cfflciJg5S62smnusX4V2ZBJ97P9pqABVwziekqfCC
LHtIXlcHZ4CRGdtZmVsM1kvL4fGLY+i0fB9rhOL2XNu2w3h7AbP+F5cR0N48kcCwguIShmx738r7
tj/+hqDSQ60xqYC6Oz7qUnT7WSYTSwhvnQ8mfx9dEePefue3KK9Pe85nc2eWBCnVVtheb0O5NH1o
X4wBqHtwNEShCdGHxMbm+9H5NBxGZXQElQ4Q+oI1LIC6kZFc+HnqofZYT+Wxd9Pkqw1m5dxhvmK4
ILgxJ75898ZaCBwcAigvwECm1i7GmJFMtSEV3abh4NGoVTp8egEuwEf2vNIVxNw3PIMqglWBezU4
Wmgt7Jy/C7osaCwo1RvwD/aCwpoDfMRNBNmIhO6244BbkCATHIfGYlWL9a92cDQP2xGFF3Hvj05p
N3zvwovAqaKpj0+oIQB0ItkUebzYiX4UxeScZMnQLE2bziioj8Viy6cezInBp3cn2MzAEV5voxB/
+Nig4pPTX0Z20l7q6mG4g9SAJvKl6V2AGNS37KyLtpL7VFLlAKuaoAYltPq53NwRjs7N2MExMhXI
k1flmIVjR5ra+oAw/rlVnDpnsqGQYphkN3FIycEszBuf0dzRo8YdOeNY0SX/l36YIwvnuVBoydnE
RWi5NaiNTtdQXJlTo2cWFpu/iGNlf0tEDPF8Ja1Dh3VlosAkLWelklkrY/7ouMmt4KJgFkgVb5Dl
qDIzTIDq8fFPaGyQwrG4R0OJkw8X1dJYNl4c9AsodlZq++z8YTed0zR9tRF0l4kmMmLbEXZTxky0
LzswgCsbBH79sXQulHQQNr5+zzee9RXDKFo7PMEDB88qAI4mBhfNuxJZ+bo6T2wdF/+aJi/A0qjA
KtWOxRdFbx0jJnD1WaRXOIUh1UrefXeP9KPfZG6MQHwxjuJ3NVOd9G3TS9MMF31wEYzltQEHDjQa
LXKFVYk04W44HP+juS4yzaMpdurzg9z6pIAFcwdHyAIgUe+0lq6Monu60GDBOs9UHN/ERVTXw4YG
YwehVxh/NcU7aSEcuW9h+oogfdR8qSG71LZn/r+1xqDMVFv7N3CLKuEN79C3xvzqTiXGrcRoIBAH
9ShCxEcA9l/cK2ZX8XP108U7vS9G+sCPI6S3EWsebx+GY5BnLSxj69rnCqgz9+IwTI3KNiLQ12hR
ckDzZuaZ9aO1gT3xo6my8bnS7JAHB/o0eMie9AWJ+IzJaYJWn3LG7olIt8VfkOPJdq+cRQXtnO2+
g/Jc+QDJl9cr229BtCzAjx3iuzoaEqFeRT6BVr7OfFvV0lwdiFr/JuyZbKtvX4/93YATG8JZebgt
M6T9+IqbFd7yYUzS09ZqHi9Sj0VJ/5NGXb0MxMoyIzvhoz12eYQopMv2A6gLgZOL01X7bLUTHz/I
ilURqT+OKoaq2Iequ1t9Z7WiaqEv/6nUZtj3Uvz3/CrZRvnHUWbI3EuNq+i2omQ2Pgg3LKwgFtnM
ktDMMSpN6vC7CdYNdsVc7V52sRz2Vvx2CLNAdZJ+/xX+Ekd0VzQHDXjVJ/8vDbjOpeFmuLCG7aW6
VkOqKg1iEd2o02CpRU4o5qmZ9YRZvM7em87sE54c6Mqe0iJpcx7XcsdeohDVIdJern0Jv5RWnb1u
zWA/y0Yc5A/scBRr8bLIoijvAcQ8/IJnrYLcY5dwt8EJNApU5kbUTJwiYHmV7qwMQ62Zf/AwSNtL
yA7sGkgfr/GOCabLDkhQp6kQQwFr8CLXa+RYIEooIsH6EtoNRLrUpeKBiaCnkaAxM9x5jpWyw5Du
cuwZkJatmE9wGYZ3PFwPPnn4s2FXfI3raxeaWPdd5vXnnekt7kkSy5zqZ1A91MxnWUrQbQjjaC04
7iLSIlSUQTbU/28o5IyJUkO1FV57lf/QJMQIkTXMwHL3HDKcFnkSAY9bRaygArvjyqvD56vS/zWa
gFW2q3LKMxwHqFr13Oo63NeYh1JFCDCeIq0Y6vdAcdEEIh6BxprA+57KpstfG1CGyLuixIDNFZ4i
9JAlH37SrF16p0bIsNvhCD2Dbdv/sn3efZbcca5EL4mWR0NR9038jG9UGNPpCEUtltmylz7Li38q
5bxJJlKRoQpnm9zC7x5IXcNH3r/K5Qf/U8Neb93CjwrKAc/Gey+z402NJhmfx8hOj5D+/EBg+OWA
genrXGj9xi5/kzy4qPGogtWcZOWEOsw1+sxVBcVNZN1QYnUBBs5bvbWmc2MwjH8VZX4EVXgsLGfe
H6OEt+4VN/N9FFOumEEuqheECo6tnHLaa+2DsTBjF5TPr6IVOBoh8nvd1zJFQSP2cOo13gIa+Id4
dMMM6QWxJdKULjYm3hsnyVbdPuZ4tGnBpY4Q1JIoqOYCsx2uE8wUz1RACHQRwr5NvdvVmzEAAIZe
Bt3bfFL5E5R/9UMAwxnZNA8rwNtg50GDIN0V1Sb9nhOkM9Ona/F0fVpD0tkk+xEwQYnXrKiHuswN
1KFvlo7vlQq023Cg8YPF5MyzEthiDQsWg3iOg7JCkt6KYqPmxRyKpDGNdTSJns1I3hd+v1NH7AgG
SImpOPtKx8YVnGCCrHj/L9KJUescRtdRLFsAQadSzSFaTbYsnStq1aWtv/aCuh0DEP0lEAGzFga3
rmBh32h7BH8MaodMYd7Tbi7tm6Gw3Ix9rg+4THUcgXL9kBwor69SjQyKx0IrV4v41kQePDUTm8mp
LbM/jGFffyYGFd5XWRAd0MsuRJSGEdxnsAmGwph4xZ5wjHlI6BncZ4SJuorsLKIOiyDJkqgH8AMp
5juXshYAY5/RUfWsIX5JmINijGeGZX5qirO4Ro8kjARzAm2c5AStAxc8TUhNvSeQcqO1/t1S+kJq
FxrkpuBy76rd15TX2wxpeaSHah58lBsxWsHabLNfNHJvsGkhV6kGSJ17OvuSSXx3e0pdiecCGR47
01rTqH21EmOSpYY6qd2ykfi9G8ttJBL9g8QD2x2iMb+KHb+UZSwvF5nIntLnzZvuoa0KEmihKOEH
7o7JcLYyqEX54Jqh+aI0Bt6DcwUo1SBi+JJvFpRuUE4ZIWFPeQ2/e/eAhOW9Fg5z9hgnS6HeF3dY
SPJ86p0QBTNHnYE9mDYhn2jm06vJtj1/l1hS9evFpKSJ87rlWbTlQM1MJj0CtTsmtocm7NDJAMF4
3jPpi5Sw8tJ66281cNgMsQCZUYiZaEf1X0YMyO76m4V6zdG9EOrrtFgTx6wNBxTdj/2sjBWxH4w4
snEFRTFQYT3O9vlT6jp48nQutMeP0AUk/XNAl77s7afkkzCTGj2VChc2PavWfwZ57hr4BBOvAxBc
qTRv4UzR+7J1OPj+oPpLPt9Bvftf/ud0jdrBL31/is9UFBDKsH6Ob0cRgDp+FOUFauUcCm0/1cv8
zlwap/Hh4843g85/KWgEXPEr4aKE/TY7kVymAkoc3Udt9YMCHpb6vAMa04VLT4j7S7UAtX/1nuMT
B2oqCEt4SnMfhuny+JYh77W8fzhzcKnbpmurQ3/Yvng98E4bWarrSmShi4Em87sMHxg/q/vDel0S
Io4NVPwgpJCPIidfo/l2GHsXznaY1AdTVAu2wZZFsxnJ9Kx7LLKzN9oeWcLfGoyEYKE6SiPg9672
sg+rSfT4UnlUTkOO4a6g6S4URQCjWza1O2ZVrgrUmHnSyg/FSWOygqlRluTppSuC0uO1WL/71wtx
YPVQc4aLHjeHC/0yYV2oXRa3nRKWzCeyFV4GBH67gXEAMoKyn6wXwh7MtDPMPGjc3LfoNTldsctX
0FnVW180z+VKUYW0J+rewPbIodeTsV8oiM1nQgLrwQ6iVKhRafhJ+JHnL2UlBmRu4WaNjH2LYqBs
M57Z3AWeHNu4r95ToieLqv0poyMuQWp0GZrFzYbDa0/Tf5n5LSMYsVip2e/wMf/Hllh6b5mUBgv0
HaJPgeQSwxFPtz3tzBbJocfU4I7JAS/JXRTgxWwkmwTLnkODHzwCIxquWedsdT1F3fXP4XIQjEGO
wt3/09Btd8ZgSDTRF0DnskEVsOmHUJmepUAC6soIJoF4gNtcAI4yAoByjoWYVDaWZZ8I8ilH3zwW
hkkmDClCvTBXn2Uq2BtchH8u+UxwpX7aQ0pDo+HA0DPemEuAx3LdkBaf/xQGQ1YyBEvTtcnZj9Nj
lWQHb4z7FWxjogsC7r/6LnBQudKnnxxFIwlZf4aptP5a/SmZik5X8PmKaDZosmGqkhfsf28z/uXr
qAbAcgQz1odzL9Po01QSD4ObkV/4VHVxAcrJsQjWGlEAgd2tiSbWGEBfT3LeJEHfd/rgKX/PlJvo
PrOLjQEnlC3tBU6hPsAz+9fbkmPwOfUQZsy9b2OLhwtGsAnxreoagdP1ngcW5ow9/GdqHALSYXgh
kzpOyDYfiRyTEHZR5CkEUqZfuVL2rR8uohIYCAJ7+fPbDSM/bRDDww1dwYILIipgUXHcDXX4Lkgr
g2j+0mXLnONfn3usOe9jffik+HlJ1DJ4QZrdu//wN29L0Q7AcTn+x8QyylVGlFSwzYFnU0Pbkepm
nwEmBu3MaRYYC0hNlYc6d8v2/WwElZN6x1YdeKcqYwqYvsvZ1Jj6Y0vQvZiqupiC8VA8ck9U878l
VTXpE7vooo+AulwmBxqxjaeinmlJUREzTYxIqnv/4SkExr2QpunMkXL0qrhTf1tyAkXfHblgWXVO
g+c+4EhtAtLvjisnMUCwnGkO5dMC7ZQZqIvPy3DeAX/0lf7F2EhlPFEc8L/6LVIdATjD6rFGwb7P
aW6y0PivO9WTAdOACTIMH8erW3M3cqgj2e/SI3wNON7pKw73SNkck3YGqsByv0EVtWmIRn+CqVzj
TA9c0Mkp+3sAZPCEt3XOnWgYCH0kBNuZ70K4/EY/WKis0teSlYxfSo3OECQulBwla3JOIQ38RQ6e
drX/sjKA7cLrl6VhY4NT+UrrsnO0DRzz4c5Qf3h2EJqUfdJaOC1WkefLsxRBgPczckUAGdNU7jCM
iJwwLE4SCbBKFcYCZrrQiiVh4wZV5pBnCZPs/l+4egxVuWOGnLVbQtM9dpabT9UoUzv76RWE5N9L
kecWyXZAPG9acndTRzMXZUSypLRBQcX6a0VBTqRq2opX4gQ+Dtt/xqqt3CGFE/2afwJzB4Ovo86U
Syq+PrJtvNlYViRpUdML2XWSXfZSKsbAsdEdqYPJJXam0T+/TEpos7AEihd0kXG/sG5QbCKjUSNO
wHQIDjkqOQt+Xtj0s3A8ZqJqbea/rrS09hJfhU3sbXsFzfQE1HzjXG55z4dhYDsV4qAlt7kNYrmj
IiSD2Mb65F/1gqX0ANrc0otxvDumUxVcGWBs4NI4tn5Dt9RwYoSwQXl0JLa6ltQZ0Rg08cQGtB3i
QA9/hEzK+g+84D4KF0hw45pDtTqwe8AVjZoyetK/viwmtFmHV80kjsz8v8yv+80R0g7gyRVzAmLS
7PIEcyQfrhxd+nw53wL3Wrouylvd/kMCnjGhGhbS/s1W//B8myIvfOP/Z5xNk2uCoBe1YhDU30m5
uvb39J/VPBi5omVWpLu6okwPm+lkENJLSlhGSQrOjrGoSWeNTg6QIAnt3BvxVm8MGEoJWSQrcvey
z3DpnhODfcaaWd+o6+zq15IQr8zmnO8WCx2xBDnTJdsp5DP6Z9oCeX/HkIXHg0DuXWHvFTtr00PW
gPlR6BYvqWHLV49jluGDgMgiwrx/QOkstjgnp+skjHBzd0u427gPim8NUw3C7nrUv8grIEC9hLoT
//QmBpOmtosiIksFVg5JZ4D1jWN0D/o9XgOvvEynZCWN8pJYgMdI57Pbz6Faxu7K/QocDqO7R1JM
z1NRGkNYMxqNue0afAHgg0TOxTQAhZYVNNjwiWYIA6g5gVLMefzOT3GNeGJukHArMQT3jzCRUreC
t17z3ZxbbKLXqqE9RmRpme0rebYQLD4g1NRbXdWbOw9LPvB0K4dIpu9g1ibjbMQTAqi/o8sNkAWo
iLUBRh/IRlDI8z5gzzkBD1XGp1MuNs1ImHs6UI/eQ49ctvlvXN8N+k/utgw3k2UV1JHAaiFAKuFm
Or190BN2ST2Edjgih14ysVrtF4V+SfB7Wd6zfQYN0Og1NFeZANdDokKQgqKl2PGFip4UDkE4OV5l
CGrk8qs+I9OCAVP6OJFJfFrOTFD9hruLzRsYILg1wVoQql0mniR6S6bM2V4k5BQJcwkpCYF4n2Aa
qx6dcDrDA9dxkA5FFTcFf/3h7iz9klgglnXMbV0ZJE56QO8aCfxvik9x6HGZJYDwABPh5gGOZrzS
zpljf0dIWgTa1coR3qohNOmvrGZd2dr1vLJFXpudpCiorYXMla/7zU3iAKNqYZkzgNJcAy1b1TCO
9xBKcU8s/Ci/rYKJfn+kRjc7tLJE5z+8hqD7xXFtRzcwR0R7i03zyiK+1C7hSh1TJlRIYTAFvKCp
JfoMa1xE0BN/BCYnyJsK6534kq2KGc5queNfHGpTLcIdNAN0lL3z5XDm790KHu6J1QOt07QkEOfy
7FpyfJDGsBxRZsuxDeo9IxensiU/27962AI1V/59J3mEOvqxyHnbBoR7RkpKC7gPsweue52NWBNw
vRlm4zG0wkJo37kohsq6yaiZlbO5s5Zatw07QPHcY4zs8vwEmt5NM8MHoMuAGrlAkb7uHb/LvXnU
G25LjF8b5AFNcANvzwJSsBXfRBHmmDIqcO9jkAwPJmwAxzIUinfPngadhTGrGSww46mdkYNLr67w
ik962z+27Tk0bTpw5WE4Cuq9pzJ8lMuu+ifXkMv2+H32vjyHb45BxGLxOgJr3C2/R02/QXdz7mxn
uyS9q3mMtidH8j+kJNmiBhZ1Nw/traSjaHgiWu8F6J7fnfcJeYvWY0YmqHmc7N4lWVpY06QBour7
+5tcp6mX+hGHUWjecmgxvdIGC1X4Pb4PIH23TYi/Wjo+Je3/qCEbm34I60MCxf/VuWpyUJkZKQT4
UBuCmlVLF2eZVcR7y3Z+cojN1I6nnm0P60u5HGpoCH7SN29MiQVVGFrJ/BnfXv/gEWaRLK8WtW7c
lV9xAF4G83wDtxh7JqZZ65JYAP20JF239hnfHsX5S8kiw67G6qTy1vupa9iA7mv850jI9GsOi+UC
UvYidvxey3RmcJCW/Ubp/mlNvYP0vTFQJtQsGZGIq+CE4kuiQ1gzPl/KQ+pZUAY+hb2jtmHlw3ts
KeSVAa7eFp4alc6deQlgWVjdVbWzl3IHwmne4womLJONATwnkYJyjLjcxGz3ERS3vLhZdjOj+LSu
yfW+aIoIVr2B3cmTxItzhxIEcKH+PG5e14TaiTqES3it1MkByScotvmllVFvrH2DsXrBtPEKG4tG
D5UfIcD8M0oNf8J6e6bpJNGR2/7LPDSqBwe9FfQyEfMo4pF9wksaqukUGdBdWuPXRhXHKUQjrw+2
1GwECy13W/iE2alGqVdi0wXBNJ1rxfOHiXIHXsFyQhQkUZ2Ke19IRdZgsQOdzppWNbWKADqitq8c
ACV6KeLebKU6E7CVc1tq4pLY5ouJKBRAaaC/4bIIJuuaNZas0MvAjCQWORQzdGQBt4BtBzh/9VNJ
/EV5J/Tpc7fSm2/sZWTD9Amb8eobb+gCRlu/Htr3OpcZ1aLtIi9wkRh5MXz0UDEj5YbSgxtjIOn+
/2AOEj9eOQSlqnO69N9B04pTe0OqNZfy5AtPEOAcpFYbiSbOfeosHUUsQHYCwKkxS8nWLsYb7N6K
DZhEtD5rwBQDN2GJxFpIV6jnZQa5vrzzQOyuYEOAowa6j0MgtwuEH0MVW8WkDJL8b5bpeZJDXvs3
0URa8HDi/phLSGXJThSJrmb1VsxTewyJ5KgfSxuvoYqYeedsDCtSL/kKs4/WfAzcdeatePB/C01C
tigeBGiGJT+xUqYRGe4UM9J3nP3TdiO6PetUZgjSEHp84cEzNWtcGNkG3L277pr3axPLwxvlurHj
kDThYZxGNc/NeI/1t5VKGuhsp7xudJ4qQe+sZhJY05glm0GIHABYIekW0AXHF14Vg1f2R7NxqEXt
NpL22QB0f34YlUDrCbZAorbky0WfZWans8CMQxYff6u9MtboKX45FEWGrWRNrQgZ/OifkG9rS1fF
lHpYGSJ1+PRLUkpnMxO12u7UAwFMp0xm4npRNJPK0H4XHErSdEOrlKaTJbgU65d10W2pzPmbwuMG
xLz/chJdWChA8YExHmilHsHyYdg4VYhdMBYEX6ntXhfRGu5eQlUq5t+uuUeqkDTl3vNd1b/tspdZ
Dd7PVGOixJ6f8oZ4yJjVBnfBkEyDXtYQmh+qsrwxP+parCAOcmflm8r4nAI0AWDqhzvqppmYGgvp
wQaP+sq+qgMtgVcIo9HCgC1crCjLLwZ8weScG4XQa4wY200bfkeXHbFfJY9b/pMRDLKCCBpE7WjO
urP5TqrryGm5JsX8FSK4RLF0JawNThF64QDsUVj3myAKnfYHuvCyi/75lo1mYDRPXRqbxQ/xEpdP
BLcSrobWnXvRZDcMicp1HIDcmn5CrrG9Q1n6AYgu8Wx7yDGorFECsToJL052KIs2v0W1Mrxg9GxG
ZsfTH8X9PakB+wq6HdQnDiqSmMzkVD1Ps80G++FAAQfTcEo2WXT0G3zjNftBlCm10sZ8nZErYgnP
AG9rDJHwkJacxkzoFAUPqekn3X7Yiz8zla+wWyWw5S4xdNK2TlP1yMkjGLDqLP9a9EZ2pc+HnkRb
WK4sT/6pYzEgys4KIUU9/2rDil/akPyK00vkz/KPR6YOAMP8kFfdn/bn2i30XvMG3lG0Jryi6RZD
L4VSTwnrg0O+sGWpRbHqnEi3cPnz0hRt/tNxSPJF2UjJ3TEbgri9Fv+TxdbBuCFhn7EYqjxxyDR7
l/ux/kg1Yia47NMfUS4qjFnOM4p3hm4J1i+YuKNd5FoZAxS4glRAsPgpKY65I6ypL0EaxYEbs62M
2Hyhs76dnLNVo5dS05cOgxtIXIyTvWYmgc2rMnl25qmxJOqImdjStJhqJstxuleg/pIzwqYvfYcX
vjnhRRZ252aiTs2ONNHhIPz/jqAciPBgv5ao5MfAHB4XIU1GEKWMjaMob1k9Q9Q0XmhqnZim+f94
ReZEjpyKeQQ47dTXdT6oykdV7jlnOjbMA3oeYqoQpouk2Yo2KG/YJSCU4/tGGri/Nqh2YKEBDSVJ
hTY0wA0lwJcL70qsltxzF7ygia9Tzfp8SBd0OnfXGINjlbU3vIQtjAEtOYk6zZfMHjPOhxsuShY2
Pz9j7wcc8LbcnrOrwN7YM1ESaH0/gzzJLzXtL2OZsf5BXaJR9G5cf0ZaLkANQqtpIvisAVWpPz8N
Y0jEviOfWTATcf/M1yPLZeXm8SPLuP3YHaAreDKn74jFPmWLQdzQKwKpnRnxhLSD+7VXROFdlisA
bSsIkSpw8GcsQVnlumpkvPdDoNnWzhFk36BmQEnIcTXQpWT0Ldy1E5+NWeZWnh7CJ2K82pzwdhNX
nWcRumh/DWUNVdTkeLlSVIUCDnlFh169ty6vVdVh7VE4EyiYKxwM5jJSkz9fdoJlh/S2L9kjYtc8
o60R7QZYSOXMXvYZ5uwHmUaCYfGeTk8A7f+T2XEpOhSSwbutcwGRBCurQ/dOdexkx6a2dS7TD12c
K6COKpwaa3eyvKi3O8hh8sp/XGplNqEJdBEb0JzsVrzcYb4mLxvnHuv2PpKJlw5vo8SKCDNdsv88
s4bkb+bOcpw5rL+aUrtEwmswv50hxgAqIuUPGJbuOMv7RzOn/ZJkbKm74J8izPmp0Gwdwyzc0Tub
iO5nLjPVFqQpGk7ZnJu/iYngaT8UCZXcjWQKIOFS+VsPywbCi/I1JD5Gj8j+n9WtcNUxX8OojpnB
CwwtYn87BUdkKukXloYmcMabJdGmJxdqRZrFUpT+1EiER1+EqxNNX04vIwERd6AXsRFovMEb3TGn
uQNm3V+egt6jfyI3z3AY/LXDdkce6PJifCo5KgvwnEHfW4I+b5KZ4GJRKz3PexLNz4kDOgGeibCp
ZcxXNivc5I/TR/n1mCEquEzgd4/IBHtEXRPOvjO8/u/bFPHPsqvh6SKDMJ3R7aKwC26kLUZ6ln1N
RMeIlTZnTWjI45er0XqESNhECxVW8MpVzd24GqjnE6DsBTigE1i8oTQTVwWgyZa3EjAnA9dcu+jg
5hYOfNJTt8LRVNpVoTbqPb+2hkifgzafM1WW32SIHK2pHseD8cO5OBZ3xTO3nwnHyJRJT8wjJ2Bz
dBcuF6tga9o8YuDcZrCpjLKm2j/R4tbqE05rhO4f4v9Jum411nL+cwpxT4twzehkBRq+DVYBMv6C
qULWZTeG42tuJdudoxvE/omqWAMMYBzJIm8ycUt2PMJ3W9CSqITEMRN9Oo/GtBkE6GnUuj/HRkNh
meUJLYx/lO3fnslERgAVItQajbVAoNVbkwOMkqxRbtQNMdRUCMNuAdfPrIcuvCAKtvieaQWAekUa
MqWs9+2qhusSGamiCCTZWHI5uCHBMaW1qsxMZ8uiC0VAK66KYmlR4YWcS+0ga08VsNdTxu0/vfLp
pqsKv7u2+9Jon1cAeKNxNGFszABmgjxPDSStnVVlYcgXMHPHO/rHcUg7BnP2gZTXgUG477J5A5/T
6a9CEfksmNwOZdj3l4MpRjkHjIaywsUDJTbtzspHxbuGlcCFLATIcNvwfL4x94WPd72Z46Svlyhi
kU+bBmo/08sdfLAZjq2+xNXPlZ0IU82Kd4zSK6aloOkxioKfmeQpuEb47YEI29Q917QWw17UqFWF
oJ9lcl/h4cYLcTg7MoxymlCmxPPHIHS5pAx3LgJNwrR/g8+gFXqoPou5kZMiWt8hz6dipJq8PMoA
G0sUYEmX+VgCIU2YaT/aT7eh7GcToixLnbGEg/gVvSia8I02g+R1wcGczCosFe6hBoYYGk2Br/Sx
bz21SiiKEJZ0IRsIS9j3b42FziE9zg+JizhuyNxHwhUhUlIGXDuVFjGnyjwPQzgjzUKOb/ZfPcKR
WYES9RHcm/LRAe9aa5Yphi2xDvwMM1Szlqkzkjo2CPlfPVBWUAKIXkWjZnbidiIhi7kUC7BjG3PD
vmFMqVgDbAKPZ9CUo99Wced9fPBiGUTEWdlmMjTVFcgxLzW6/eHnkx/VatQrOaudnaS8zVTSHgUM
Bkx6bnF9gKj2Fv1ffCUWIdVhRRt1Kjo1erJwVvEeTa2YkMU2tGFQKko5aLDqeqlwn7N8uxhbxf44
vanxXGhCso7bbdASMDk8r4y9WULixwv8wn5ft1SdNzmqa//+hPP6ddyWUmjgErUwta2WIpJgPDKY
R8KIcBM5AdYNJ34JWDlvVjEMjfFXbDOdysBcQ2TCjd8+QAOiXlRjCVTrOyjZiboEB53iPM4Pv0US
2dVveGTelCiO8AHLKbAVjIrtsU5RPiKzyY+fJZRhiWpy9OVZsJ1NhajFh089CWu2zPZ5evD/BFnn
TMx8vKJh0bQszvYf8Zxi33yh2thXvIY0uqac/N/BrfF0+7Spi6tOQqICYe/pCzN9Hngsz2akp3rs
0nAs/TPj+hSCsbSCtLMCJAAn1r7esF0TwgnhE54eEEEF8KgbApDe4Ts/o9+YVg5Duu7TPtfp04Pq
ujGfpsmZBQduskHUjYAW27jPkRXPil51/HtkLHr+e0KaH+8mHslTP2lQCPjU83RrT6WRUlSGyqqv
8+2/Ce+O9EP9D1+w1eaft7vovYmtKwr7BZDA6FmxeOoiQ3dbwUwdHMyALT1kh/IKWyZdPaQMV+No
X6H5Z9/lrHvotYR5gTrWMViAymp0JpLQlmWW6rjoNG8tKQzLVj7YtCMdwOx28vlqDJtcSU/pZD/r
XhBw7ppJSfSNz1p4eE2E9jT+9YhUkNBilXR+opWECwQbdCiEPCTp31wejZmAgl95y/jmfah5sNgD
xfBispIAgSKSqH43kTv1azMRg4E3ABgnwQz+tMUklthgzi0XN0aA36Eg6KQrN2zt078zIV8qufW4
hm2tYOR1Zri5YA+tbiHqLTKi4zd+9QZixenBvMfL4HmIeNF/Xpp81wxVqLXyqwL2hcKQlI8whJI1
E8X6bBN777rcG+o92GpKDTzBFUcJfhkqD3ZzbLSm0a597I2E5lwLugv4n1cebJFvSWtJefBWthTk
+VBs9vsiGzRnxo1dWZwnjkamg1R9e+Emr4F1Nk9+iOUZtpA8ueSIB6nYiQgi87rtddQFEz23b66O
G9Sw7qu/1e4Gvyc92pv7VqD+EMEe24ly6MLXqJwRh2OBt/EcRumBS434Ht6sfUx10SXxncbCeABf
08vWXfhS3Oo4cm1Xf6C3dgMJ9RS8K7IrQiwaxxWeKfc0F2ceSJyLq21F3o0aAHi4udo8AEmtDKVT
DQw4HFSBZOWsFlK1rEk6OCRTTwEVNuavb90XawKJejmY4rJJR1rIFFG4ysoJeW8vSNXYj9CGwUVa
4HM3iDm45tsxzUSxLzKkMmhOo1IBC7ciDzlBtUHVAhiuhoYYPs/HDxHzp/41eIwaiBFr+9LwlVQL
xqmdb0Jl3JYHkAEu1CsO7ldq7Rh7hUsgIibwxE0SRqw+3oKJFJPkDvYw6hW9B1R+hG5pwztVRIXA
u06hfFiL1TrSD9yDvWGqe6jGV2lGfy+Y1//o7+2r4o6pxtbZmRl/1W3emo8MIkavdF4oDaV445v+
z7zuvO/rQdo/G3DEju4PKkWOWo3QoiiWntiTXMqq60gq+Kg72JN6A0mOlCYDT66MlmttubX++Mt1
RwYMV+RMhjMwFf28JEIpuU1o4DnWRHHVUtdlgHa7XIyvJEf0M1X+m1lC7FteN6Dg2Hr7MuCE1PqY
YDdiJ8NfVUY6fntF0hfaiqkO7wDC1rT2VG5yTvDNA5vOPMRfRaL1kgXLZpvIIEIzFnI0ayg8DmKP
82pW+FmsA4aF35oprKLrNC5UEa4WGHA+9g9Kk5radwkQm0HodHL9AqZQdMT3Oi18mdTro4C74Gu0
TDSlnvJInJpIN1V6Tf9kkpwYl8/ZQQc3RVKFQTunfrCaWBJCPMHGJArEOxg8vK+nvdg+dzFd6vge
njBhVGZAf1jPL4gdfWwK9f4SjEHVzQcLDDLlLznKpkIK2WawWUHkflK+ihIxLlu9zKa6VcP3Hz8X
xUGIoJBwm8cYSn7uBcs1s0fX5oVuUMcFLf9OO8wKXOE7U8BBSBtZT0xJOm5bcR38leVDcSH4RWrB
uaeRrC2bQaqZ1JTY25tsaqWjTEH+k9k+8YVQszJQbZLbIRjbM1PALxGP0MZnU129X/QLQl0+av9m
1Jc3brfplODCFH/cJNqgZH8DEfB3KPV/4I7ENs2PB21rlsei4kJ4SiDdENktSjOz4DM4K8Ffx+4B
YiCr0yu1s0pgMBnj7hw5wQF8wIYlhwugH0Dl+SrokFzU7UnHOCBRgyxT7hnXyTgGMpGBukvCr3Mn
t9x6nl/lRVsuz0bvudHj+eM4lH+inNHf1GbUnE1TKb9MKZ9O59wX0hf1pKlFRR3u+I9qfJV/S1Kz
7csd0rFnIqIhQn83uscwIiXe7bfsrABOwX3uwjdoZafvuDgaSe7zp+cZYqUhLEyyQ7YkEukO1Ckh
ZR2zPn3n6k7m/HzoObWs9lPwR4FPuSIXm9f69UadMsFpncYUU8Mt6qbseswoFJHvTLaOAA6nxwYI
n8XzMgSkRDgAf9BYq12THOd1dXzH4kUHYBS7qPO6CVJm945/+okWnOtlqigtP5fv9tZJW7esZAU6
3/QW61xnmOOSGzXrSVCHCwhdvsQl+jdJSrz13h0/U/45x3fE/ce3OL/MSDn/dw9wK3YoLOJLM+nI
LWSdsc7HXhSQ2Wbr7I3vIzgF29VSt8d5QVUkyH8Zq4HotvvTvczTmygq1ka8zrFNU0C8RYKeEL/K
6dlwj83m/WQYvPEBGVvgDlWAMIrTUUJ1YBu7ZCNWroFm9eHo7ArOvUu/qNgt95wtz0YRKsMkYiBy
hs2l5OhkV1nliKgHVPP0IvnxUCP/SYM6MLlViGEY4ViaFLY/SJCVRSXSJdwA9qWQ6O++/CS8iJV7
DCGTPjk05LDXdrrKch3gCNSsW4JDnupdeMzgFpUjpfIhj3oMyqDOLo1IiPXUMR8GRVABp1VJihQR
EPY6tbAMRNw8729d2q2NeFFTUhffV7D70gS2BjhX6wSpxvnR38b5zSKmPoSTpAwcCMoiz3ieduaI
YpBpSSkzfBQrWCfk5ynA9jZOPsy1SJMRWD6RxKsLcsiOgyRy4P6XGDaY73eQ6cI7VVbS3UD7ThOx
Kj8bWbU533jpIe/1wtYCArM+wzLtCQA8Y1jwpm47EhZm7vj8uiTMi0K9KCgiNOP4xUgN6AvgYdbD
UpUUK9Op/SSQM8YI6BJSDv++XmL3o4C5u5cBpqNKoVXiqXULzo5EJq5pfGl4kkBPDMfiurd37Ym7
eaRd0A/Rf68GEe4eWiotjv0PGLXykEc2ry8jtB6LC/ohRdqFtIEa68f1GANZkHJSCnQBS/i0Ec6e
lsF/hk1l8eMryjC5cFV7RBIGYG3r5LW6ySZixjfs91Aiy734uvhDJ7WR6beyh7QmbvArfJ4CaqVG
v6dsKXGQKUlXG6uEsLWnuW6pO6BNZREbZ+JZQiF5JPGsbydhyfi/V/vtn5MIt+9eb5mV8tqu+/Lu
LreOvDIDi79p13gxbcfH2+YxXueZc2UAOKQhgBcyhIQ3rMz4a99OszXxJVRcqireeFjoQw1GcbJg
UYWwwylIDKd2lhFNFPaJX4vE80W7378NE6bxW7jBTZ5XMp5CicsvGse+pr1UHOPNArCkCl0z9mYf
2v5dqeqrwCQFD/3+1b42rolDaSA7t9lDTbwVZnSovKB+OWBkQvDpJDKTMcxWr24NsoIucW7kQPn4
VrzcOkSp7Z8iFEycrmqDVQOcxKafCG1yB7j0mAc2B3Z4/eoYclhGwGvlOGxbf1giuK1PmCArCzNE
D2+Qawo2FBO12T1aDxWkaKoBWPklh6Ms/Sxxtw4SXsnzu/P59vg7u/KdzrY3dpLv9oD14Q0gy9+e
2rMMcuRnsHinkCfHly+ze8TlDe9TPxws+wyU+zunrPSEkWW45tUR/PIEN+AEVkwnvNpEuDn7ZpgI
aw8ovH2HIg3SCSxIULcSubFOPx+0ZjsFsN7wJDevapIHir8pYxIZDhIzrXZ2n4exEwS1Se85YOa2
NtVVaRIpzGnBcohjvPndt00jPxhjmdRY2YXZIHF+M8vIQLpmi2DZ0RcHyg6wgJeoO8MOaq7q9l1l
yPyQqY2+wc3Qge6D4hzJ8ZzS0NlqB8mFafbRKZUfblpskwispmAu9jOAccg8JF9IKb6llAJ9aNcm
Pjd4RVwaJhHgM2UZpW9Aeo0+SQX3ifSJPOTfulcJjRofRzfWfBRJOiedh2AgCzg9TGfV9zBV8II3
IFwCcNJ9TyXOc9ceVQvnJL/vY7I8JrBo2+HuIVhNuVOeQRwqBFZQ4L3KkzthY8VD9F3wIoLXvhc+
hATVOPuGquyMboOAfQDZ9/hxReTqAKzMtjluFuf06JWTZ+bVTLnvDL+f682evzlHUQv8KSrpGj5D
O14cxM0yXNgpIDX3ylmTHFTeHMLGk6mim6vkIv5W2rwlKKsjDaQufrz9pGDdMIEob4hjEx7153ks
1OYfAIELHbt7g3cE5W4JMgvHr0rvQQYCUPYrWyry5D5fOHzVpUuELTiB2RB7KSqrWvOtDoZVTsk6
GeX8bpKwTDwEg/Nt2AMbBMoD8j2D/wu8jYfNM0FVCiZZCHjyvKMZUTvKK+1N/bxd4ViZNiQE/ruJ
+5jtRotwu/uFj1tSZpbeuqfVLcu5TMg74v+cb5pM/fjXFpGzVmlBoeR2v3vAqow2/RMv4byBWYXF
JVWYl3O1yYM1uVloEVu7ThnY1RdR30uYX8NB5buIwJV+ZccaCR19MnwOIKtU1tKZpTersvPDLJ3K
SLyERZdcvpEKNxJWr4KUW8RvIN5wjA34RKQ8z46+Bv3OAl+l4CugZSM6vWE9Ju7jPQPRj1J70aYw
CkpWmnTGOtCwIcd9mxHD1ZBib8y5QvnKwWNf9zZUB6+VhNukEeCyyaqZzv6VTCIFCXIXjBGYqsuL
Rq0dyT5o2eIxcX5sEU/kSqvYfmXxZk71zws5G7sVuaOs+rM6+pl4KN5lxXn7DyNen2PTO1xJ1Qbd
eZDsJGKUUglok47wZ63yZIem6Yq7mN/HRtj3jRYT6WtocwYQM0DydQTU8UvuEwFe4MBgL0ULT+7g
D1KJj9C1aGHFj91uo0wY/eJ5gPFrlWRRD8AQO5X137kAdY1ogWmfOoOaeGF4Feiy5ocpQfpMAuM7
wjGkJG0ICsaRSBw0JzLGO+Om4bIW5KlKzF9wVzfA8kPlljVtRo0kO4ljhg7Nso64jdP4mstYt9cw
iMfSyju9Mgsf+pEaCrA9TFucGKAnspI03S+pIhQmt5wvPoIcZlrNgIAxXcaGkBhCDghN3i6uxz7w
oEfNvzxpZSIH8hwpF76k8agdX+G0sXH8j5y3RW9OYFzg2nMlkpAXkOdOFnbTvZFZnt/e7s7Eu/N+
9LtynORHoM1Vczh8+Acqi45hlaYmY23qcrfT7knpxfH1SDB3jECc3WzDKDuTilUWaO+vWH0DPID7
i56j5gIqn4IjBOLg/wIeinVe7UbAgvJYY/h4/0eM3Q7xLWEbp715uWbu/Q+MMVSbXhHN5XgkzZUX
Stp5wJuObM/ubmaZG9BiE2P+583KRDW1QFcA9YI0zAv6w4ipp/dG0BYgn/xiA6N+DhR/6WXANyrB
MExkRoq6T7+jxo5jCMlNYuomz3J+ykHfwuOKcn5+MN25lhuAJW3Ch5b4nIJPNGkOxILoiMq35tx7
M4C17KDdLnjQkBd2RwPLAzBTYBri/doeF6VYY6tAdfKQmvBxaNY/KHpdRXRbrBR2W4BdTlYXdb1X
sVV32safo9g94gzZE6BpKh1ecMzFgto+3lgK03d9x2mnIYJkEs5wC9ulg9zin3ULofxK/se1jPps
FqgzOjqox1bn2f+DcmMDBp12Jvhko9iaLeEhXVf1MnxIDGPFBJbNDiR3iKDjgTixpWoA5ig9mxHL
yx1hFl49++6U4rlvlPtYgXxwhuOO5ELixfZMcwLuI4HYod09pg9+AUW8laxaaRCTfSnHbZJ1K6pP
Pvx5xyiFrmM/M54gwLZaDFJUDLb7yD1oTRY6CDtbCeVq4fu0afjhgq7vPNej4+4RvcQ8xcSy4Az1
qzlBQ3VwNFqV0MBtaIu6EiqTO/cb6e0k0lOP8bTuMkQdyNvm2FMnbPA5Ry7WrYwHH+sCI7VGGiQD
G9SwE+faX/hlbXNwtvwESQX102DMZhsJsLTTZZGmmurQxI5jEOVl+d2/iRvvT3dH45xR6DfuUnfS
7jckN8brmhwR8WoLDtnBMQS6bLVJe9pm7ce2P5H157mQw6dsMTECvxihGF0K9V9NRJEfZjHcEnR4
B7uV4c7QmUU+cYG9s2/izOiEnRBn4ZpP4gou90vb3HxZin69r31oa7KURZ6XlootlGEdI0RXX1Ip
eT55An+0XqpFuklo7E8oV1q6D2fdIWkWGnZL6kqkbb0lkS0uubDUMDdC1h6A8TT1G6hhESeZXDNB
jjkf0Kw+XTD9w7uGp8/46cZ+62Ye/zwrB8XxXXy+1mFG603dvqT9cQHgZdIzazWGOlM5pd8JFqKg
/ciaX1J5iSZRRnkbNuWXlA6ay+seRi0sH9slCbCVhTFxHEheQkLhHc/6ayI2QABztMQzhBs116gG
vvDyR0Ly1uuF25FDzoco3HlTrkFGzHZvnAE1FG9+/9Hn4EjP+xfaARY3wKfSFQDRfrU0CBE8RJY6
h3+6ESLCaVtVRagIk48WtrFb707C2DVupVcCDGpyWJWruaIrmi++/SHLAUOlmm5jRi6jKFWJNtHf
FHKQ64u5adbrI1+8Lq/Bns776VnX0uEMBWIbuPkEjhSlz+54ahyvbuem8d9mF/YygsTeVBXwfceK
YCdTY94xwBSbx9+v8l6QsiaJ/rI2FZ/2f9yTpGnn9a4CFdVtxY3DEystJ3IZDZcPh9wsCZRfklCO
9at4J7H/eJ3nq+iV8Md241/ygI25Dg2OrOmAfAZUb8YpUUnEm6BfHBduHuXX/WWg6FEjirHGIMqy
gZyM2QM+xA2cDrJPPKm2DuXiHclorvBlX6F9N/yHCSCI5xDMjXViPurDYzfyisUuYcG7zR7Q8p4M
OPmILMlvxBKv+OXrzj/pbrZdpaguDnpzNhoL/V5zt/78SBm8pH/oTWi7JqZMEzY8aqZCijDlDKkB
2V2xa00tBC7YyU4J/7c3ReZCXMJROhmvsp0WhETfTzPna36fL/r2dIyoq8fGUYKemLiOLqxlZziu
dgr6f4DVsSBQUYC0PkbPqwbnGOA4AGjla/HcyfBw5RYTDk16fMU8wm2RdwxMCrIBZ6KXdehYZals
+swqrgRm8l3V4T07QL5aA48Df9COznKEaPl8NL8qWnp3vzldxwTcjeuSMoztuhPBv5nVuqwkJDyU
D2QOE9XGYLj7a19fIWKpLtolUsXybtzNRztuR4ooTE9f3PWYgIZC+hXU7Tnd3R7ImPpjc5Mg1wFz
pVY+/mSij+AlfTJ7+n4dV1Ck1aqERYYpGKtZXyKcsaARSgbqY13hzpKM75GwtM9Enulf7DPgBILN
7o2Fzx1VNh/e0T21lKocJomfOfMlJA9fL70KHFbmWCoRVEFQJVmpuvq+8Afo9Yt2Mvyc6PAPRonI
8Vuzz7RjWzUxPDFtoN4rRgITKpHQ/D1/3OqWj3GSee8TbQN3dYYFe4Pev+mYqiSpQDoMF3isGmYx
n4j1Agrj0/SCjDQNtqMEFPWPq5fVlmWq5ARLC/5Ze04oyIf5d8rxJoudAHYMs9fJ2ynKa/pwP2Ie
ZxWed2b4nTEPVwmlX5qfc0+LfNxNoc7pQFaOCtameHoLp/iEuVNAEonDPQlp9ie1NvE1entBegVc
lyKrZRf3AaN13sELjGKhLu6hNwfHcyyEhAl4knz0EkwqK6VhlCtnRYlDCtJAzdx66KvX8MwoGTlX
MUcQnW5paIFioyyyi6yTU5ZFUwHMmR4SYP6Oz8dYTww0t1qS5kkX68OhunesRiF8qPmpUQE0OCmh
lIed0c2luHvKBNcl8RkjCUg8MdhVcmhT+yU7ezUQRgo+jtGN+vCjWA+QhH1zpAUtgOq/0TMB+++Q
PAdnA3fjR5tSQuzmXTR59MmXdvd4j1gLRGgG6resu10HYIi9sVD0EupPUPHyFK5n8unKfmviTNqi
iT57SE7f7AUKYeLdl1n/Q34q1xIY61L9SfrV8YEj2WLw7WtxK4Ks5z84XD1GMWpdkM7BoXuN1EmO
68guQF6jd0Mp1kXgWjEDLMkzvOxNpNYGiuIolfDphVTmBf6NWjkuiIODfsrvb+Dj9ssj4GxZfmfZ
rzDq3zsXtSa/pQhS7Azi0f9qcB1zkX5h1x9OV7do7VjG3hYYEKtnwPEOrwmmX/IIfz5E6Lamv+H9
DEMPCwrkQoNTs3qhWXDAtDHl+yBolPJQtEty2Hclyz8SUJl4W3iioupO/ZNxbFInlJoqsu5aNtxI
sNXZKMOeFUxhBoi54ZU6IZHXyVQadR1IM2kF+J85kIGdM00q0MQJB20ZCgTMFgz0FW278lNCNq5f
ia49hDV4SM6PkZhzNUIPP8QNvKzuiq4W78eP0ZjcuXPvynwBGubRQGH4IuglbUBTdlT6ZG0uV/pT
Os3SjkuKO0yKSSNZ50XK+1l1PUys78SNd+pNUsw9NrttLDYxQUcLxEuK7RP7rg1cgisBsyOLh24Z
WAIo26LRJAWY5W5ckuvc8HdMAuQxsEsFuyt62dute1lDJLjjGZ9KrgQ6hlCirvmH9rw5FtSk615s
vBtq5MWfup47YcaIBBjkC5LyUAdfTF7Fa5P6zd3vK0v47QgTEzT74m9igjOn/WqD+eJHS8zsE3ML
22/mwnX8BRdfjujwQeaV0+ZDOrSGxO6fLZVs6vTMwjYt+BG4l8P4CImr2uoSu78kEhNNKJsC7tCQ
r9YidifTe5n7SAa5+LKoL3O5QZ8xOadz7MLV1Me30+20o+/Yf/5/toXA+A/lJhe4VxU2KW/NnM8O
ExuotGtZKUX/IBpK3c6GREeXLnjB8yRZq6TEWQET6A8ohk8QBCG4+9ROtg3hAtj+bq/MNDrwYSqS
aSIoJCWpnvzpcWU/Df4bdDXDbH3HRVkFMSqRJQ3HprO5ef8OJYqn0p95KZWdfv9nmDDeZMnK83BH
pOyv72oIsj1HdU7Ay7PqffLXiM6VL/FPEok850lbvTt1eaZ8wrb1mW8iza9iMX3TR5BQw+F0lacp
iECDfnXersVpaWLkCllqyrP+NMzd83zMuKmtKMjFHA+IYZD3QswAOV320KbmNZTh5D3lo9MeqNXq
vMRJDFxROgkOkhIWNDQw61dGDHO7UWwt1Blh/gNSswoReY6daJF1GYX36SRDlvbYBaRyfX60S+Hz
9hfGZ2glE50djjDJRr07NAkqU4GLhec7s+C494RDI1Car6bFhVtZaMRd/TSoBh9zB4UMr3YrF4Re
j9bqsCiIj3hyMccUTUGfbnrz/NJwObyjdklamNBywMjYq0Urjsj9gV9LVt0ftYVmVRdd6DtjAs5P
NAzFOt2cLvoywY65q1X6p7WjRs9o04QjmcxcfMc1hUQe1ZY0KOVQIM2U1YD8rxJyg/dEEbL96hNG
wAhY/Oe0jZvHWT6SAPXXxyKmb6JekwLlLvFOeDYO1vaZSEzRmjHQbL+PuYrP6cnfB+yos8dv7U4h
aTR74OXyrzzg0H/2g0ip04HkmnVYlakz27X+mGl576AR/GZL5h/y85b2Hp6rEVr/r1LycmWKdr1G
a5+2FJrc4WqyNnT2en6i6KN6sL/K7tyu4wHyFB0KDHdlOuRq4u5jrOHQD6F2kjHZHWT75LhmNBmA
+JxYXg85c3gtR1qC56UEIz0B43+OwXTIIytF4oCL4sytAyhBjLlMMiGM6WbyteRGDQAJZFnRcqyn
w8yLzUI904GubkzWuLUoFwIVQ9fM9YqZi2CNMmS94S7di/Av9jZdiLsC/WrnSGdJVfoQslfT8uX/
b6yAfMgwjEM1LN14e9MyvgZIdpPob2xnR6JDvPXXalHO41Db9JK4o6R//VhwmqSIVQW9eZKEkqWN
hZkNwR+CPDNjPMEg09sbLLMlm683vpUCtJaoq07rifL6Gd7u2TU/2AAJy7l+rgzkBI333LGgM+ca
fPsJTnptoEUYPmQapDM0x1tTa28D7MLB7EL/SyF10NLzVMRC53CFNpqDIKf7hNPGK67ZAji1j5f5
5YqzdkTxWuxKYRYwX+ebE35Uc+IZbMCwTLrWLn+oM3JXzWaLXqlhiEMLPrZ01RdBXtaPL0HkAFi9
czUpLKRYX7dWDkASld68JGwYCxt4IabWZCcCBvm0mrK6Ww0I7m+IZRklyRvLNIGKrPnEpDgrUyEY
YdswcqpfUN1ghvF0FbSwwtf2I42RckHiBCxNWwWmVFpMmL1RXActsPB8R2M9ahHh9IHEfaKuXSqr
CAd9R2lYeBwjf3edTrSxs0mj9e50YaSmyZBsSwD9BVDslBRz5qVxgqmMNZ5aKcX9InCVbPSB0pk2
gA8PC6IM8jmW5XH5zNczmdsWv1OZahd2ila+SuWW124YWDskWrBMJPa4DiO7yF8k+gNr642FMSMK
ck06zLmkmmjVZmfyOA1u/I1GZQZCS3IZMQ7aiVekki/6A1VFTIyeYkf3oLYu/1gBL91GLQy+fzoR
iUqP4L8x6RJXIO+XDikT/tfBUka7DJlh3PubNapWRYbqHBMK+Ih7XM17mrwvTxWyeRzwysCSAbnV
y577D1tU7KTnkwMmsjMuaxHMGbNaT+St9yYoMESTYQNwYCDz5UC0UjdaTzIOqoKuHRPJKCTVAIPF
JVWOb5wpJHnqLpWbBKIB1B/LJTgnxQZLUz6v6S5kyw8eawE1LFkVEGHQ/pYt+OWH5tpH2LSWi+LT
yB/YxmM4HSE9N9DSwFLiNdsBM9lTxmvuwRwtnYNXYVba7s37SlPDbDYQyoV9wNS1Vytasum2ALUJ
N4a38SkKbpho41ZZp5fb09UTGSLIDAbQ2QVOWHhsoiA+gpq3UDbvm6LVc59wGqNpc1rshcyq5Dqh
jM1aFUr4DixDVFnLF+irlIEgnrO13SVZ+p2t/jQUmNLzviQB5wlZexn4yjq/fnHv5O3OQ3C7sRC1
v2GkysGMMFHJYndwZGfNP0DyhUvZSrPDFaeQ/TcrJq7Qbd54vlLEgQH2cQpa5NcWWsdJhFbslQOb
OiBYX3rMkZZD4QvbZAkggRRpAoSwcUjbUTkMHne3inReOEsvc5i1oIpWXdt0lgpFBrCqh7SR4XXD
eyq9e469yW7TO5v6Y6EpoT2h/hLcRFq780kAQsFFkNyg31fn4mjVEg70rGWepT24YPo0gQfcxW8X
UMgjn9VzEw62YCcW30oaaAaLgb5gfLPSsG00pWY5fnPvlD5Aq7YA+isTifhQiKJqATNBFfZ2Go8+
SaTvxdZzKgX14W7CTymFlSPtUc8EmLABVW02Oq7y7HINSHU6L9aM0BW4Jlus7POO1GFlR/0Lah62
y9Cwqmk1S/FCPUPuwUQdvpnPSUO8mDvQXbiUp9KFOF4aZc16tlisZrG9WYbYS1nVWQI+tvkMPncA
MWpK4NMR2AEYn0jMZfJ6TwvRjvJbrPSR8PHeXi7XrgUx8M6pzd2jgznpbH3A46+FCEEc8YXDC0hA
IYp7hlmqIO8Y5+7j9ygwZzhbPJ673XuBTMDKdq+rU0ICafyEcn2kaCCMh0W2nN7NUYmKgAoJO7px
E7ElD+PhUyiuDo91cEZOtAZz7yXAD+yFSGOYRMX3XbTfnjBCxBHrf/IPxUfFoa/VNAm5iWaHC+3X
JtezXQfpzBmrci/FYyEp0MUwIg57liqVJdMtRdn6SwAy2se+N6PZ5lOlvxnTyjWXCW4axZWa4ZJW
zi9Di2hTBp/vOjrUcAnHE0+82sJLLsZEL4EXHkp1gPuFV1A0KqwH2jsciLPPSN0uF6DOtbOWhDMo
KqNTn5CO7ryk9e3fVCDEu/CUALtXXHJ61OpenbuEapJ2kuOkGQEJfrdlAkqqKpyirxsGAPTKbaL3
GsYUkv+1wGNBaAbZKQg38vvRel3oYbHkM/aqWZKiPWyeVhtc9cZipScvtm1iMtkoZgP3v8k3rZ6G
UGSAEG0SZhWGGD55L+jSsK7YQvqSKxqDrMZ9Oy9ZhCDXu+eocxnrsvnaf7ppuzeFsuQL1ZZAfHeO
f/bdL7jmWdYvlKhpeJkzXri4kHLqp+2U08L3vzyyT94fWi3WeVpX1jfk94C3EBQnf1HawExYm9Kz
E4u4JOpkB1kv2lalpxWBrpNcVmM9eEg9GC23229rnaDxu/mk53G8aFZC7gbxZtXfj0en48EMSfKX
ChTyYgFXEKPlQ/TrA9zBG8y9Y4nNqAYTNZmGgSH3ENWJiiVJ/yVMrqoVeIDOWgRdj4pFnkwKA2FX
O/CMFFYaoxITvIfirLA1NBwCyr9vosxDRYGSlpuglZwn4O3hxtQjCnzXnDR0EMIcp48ZgRHeysMy
1g+5eI2wrgJHG+QgFpJDzkqGcdr4cU2/DoTj2UtqWbkFNpyQjZxx5ZjfssE6wAiBAzoAFWugaooJ
zCnJjldCLpcrfoOlM1pkQ6KLVE6i8O8xcmYHMJI0Cf8r4UG0Svmt4tcT3zG4p07744JDta5cUYaU
EQ/rJRGRGD5ZXa0lHj2r+N8/OJVXwtem4Toa0nFE6lqWWoddHB/Fw5LEUmxxEA8G7XkBEFNGH8ig
w7S2D+NFwrnycoTNAUi8BA5WwLTMi6Tq+4pRg3+JS7jkpKsYFUmxkIxwsgFWIPYuGLMIeRlDwAsn
NbV/bmJTtG1iX4kw7EgDr/B+7OqlO0zU3d+fn/i0kxbsSTkX9maMokqPMGBJt0P/B0PZ1yY9p8pQ
2Ada7zn34ZqFJFvatX9005gD0GjZX9WdWIQ4IX15/YdtQddYqXm6it5xFPPkrWSbB98Zb5ih0quZ
IPc7z34zbJWyeBuz5YHYQMw9+vJnw5JjUDbKKcQYPRDcuSC3kWgaAJXVrivJJOPchTu4DCG4guUV
7Bw8sXaAnU3DB7VAFYFUlJQxkf9rXPugnbOppfdeq0EOqQ0tEVRdS64SVFmJyc+f9fYTPs4mVPmN
pgDRK3NGPJBGBvnzk8dcJLNZfngUzojRy1NtzbG0cpra2D1owR0xkb4VIOioWVXn+JdDsRavLnps
ajp7kQI1dUKETLR2vemIBxyPVudn8J+fNQFBV1mRARuiSpeD9ORdvGXGsZq4uigWSYXlfPGFpkLp
OQly3ogGg3jBLRrd6z1tK8jc/2kx9HaNHBtMjApKHbh5ebCdljq9vYAjNUu3YCoun+SjkMYY5ptN
edeZJNEtQ5he4PP9V9cACW1x7cdcNQfMgCkpw6QWW6PMin13kfKy3Fb3f/1rR2Qi6wF0tlIzhkNv
5f9q7xRAuhcOrIAAB/x1BhGJvZ7S1pPdr/bQ2enDk8q5PKOWFUZYZOt84ld/Vp0igzf8a15mBY6B
u4sZIAM7FzMOIbhWNAtNMhfmvxXQkKcFe/UMtikOXMJ9mlEDeg5DQ0hmUQm4Uq/N/y2C2n0xEFHW
zbO97X2TSKzKLWfezQFWnp3TxdVuzQqu6HSlVdiiTVdbOj0eCf88g0UAaFBL7+nzK6pZnwl8w2iD
WoNt6ZvS4+YiFvMxJ9fevLaCH4hzeSslbtXBkZ3uSA7nNzTdEkAy1dgAkHfS3/ILybUi9gOY0YIk
aUdfw4njCAht5ylaakZR9yKXNk9G0JKVgZ5Y7T01vksyq2R/tKLXW2ieDvm7dAqZJljdb9hTSjtK
3WfmJDTi2/SmY6SDUJirvMh4AgUQkU5S6iMDo9EjZc2IcnoxUuJpwgJlLDDSvyo3l08Ich8DI0yp
sTtBLt7ts8W5fIVQy+dP4LHbljXqrcqKe95G0MGVbThrFiGkiLrCdOit3qKibexKNt45kO3J2P4w
yMnho3zQfQ/K3Xd0yDI2YMxzViLPZB+bSk4aKkjQ1UCWnj0IewWrIvLitKmGPkHyVE8A1RX34cQf
sXOU7fgLzfiPsA+KwM5IRdXoW9o8cBK4LhPt7SC6AkCwvm+kAeHEIYaYPixtYQV+FnBsSXwmze25
3nSSjXgHnABWoSs+stwmZmdRJjg7K2lzpqWhaqWR6TN4MOdysE0ajO6xPVIofK6vzSlQyYrnGNQK
i8zpcY9dZtLRHRTwEmvh8jP/N5eq5yGb9dcuYist1ltuZYUmVVsL0fEzY9atDQcs2caIr6PpQm/8
XCthTS819en5qqLmZl+DiirESZyT7qzdDoVbZJb+SLjfuIC18+k77jny5Oeyc139gVtG144cex91
h1e2FKUAmrosRhANnfKb38Bq20C56S3GQ9C8MwhAyZitrhL/BMh0H8ly9/+csuTgRmxodKc51xGt
nX69NKpWdBI/LrkswMFNA4iWMW0516iU8G1mQP59eYusXAlTy8lSc9ZC238Swn1yK5QS++YtXEa3
0bwuhIDd4V2FLotA3y0iIfyKPJAK3qbxUQgIdioWzw54hnBe1Uo67QZb30gjWAstP4+jhXzhJ/de
q9P2REEVFBGq92Pe8Pi0CE84uUXHcpPBlBC8eMCHeO6D2swUhZXPH0Z0PMjqSQlzyPfObaJEhLcL
FoRRaCXqWShkq75UBqxhZM8NUQJLAUoGDDtlgGNPUtMv7Q148XC8JK4OWVuyH2hRYJgD2IvMwMRZ
qduUR/d7+/ojmbAE1g60YTKQt3U4TCsyVQclqSadg9nGbYP1pEHMO9AXFqd36ov9MIbL82wJB0yT
ZwqVs8Zt40vS3uE4hVdGqSvCvS2VxfgNFG11uxw9dL9eKJRQTJfyG7Xnf/mKEBGKacc+WGZzH4tM
wbMz/APw3PBe8CTAl9yfqZPX8xq97rX8oV1Ah2JU3HHDP/bu5tjj5r/5tm5SarfLRtFuOISIMkLH
XiwddwJKO5+XfOEqNBD5asFBTWYUeZC2lsKLRfGPyCvqJfvB02JSixuk3AzY+DR3dzQpvaliuFk9
4bLKujBhpyQgkIxoujh0SV0wxa5M0QaBlHdxdDdRaxr7LxpV2+baIpyeTACvAanSTQ0zh2MPAdXU
JLtC3ln2AyBW92n4U3zuDKdZGJK9ajFjYn2NKVUkzGzSKguO90Xa+doi97DBppZqOXu2epDl1LJ5
Pbr/LfzYAgvUA+zuQt70lg0tQAv6Fi3umxRHl6ynsxa42+wvYH+ACKDzAWwVAipI+QXEBlJ3iYlV
Pgmy6mXB5cIQOEs8lo0X4WZzEJsm+cm7Biy3pxoyyRilhen8Yzq0+D7lWuiO5uUX9wW3dOe+OOEd
TijCSqnYDwUPYzPIGyrMHW0oJXdztCvQD7Os8J8IPRAXFgsOn1NH2V3uXnb+LNfp4iO7fuBxM+4Q
yf4UjT0xhu//YRXbXK1GV6Vyl2TKNPZr9zwJziOPAEupr/ZM7ORfpBkdWTdfb/H3GIVPQnlX2aai
NgjxDpqZbxFs26fNh+gV+8qMtxeV8sjxTIrXJ4aEHPRNCQ/VR7uAtcnaaP83wI6RGQylnhUhCc93
Z7r2EPbFs6xvzfZ2Aihkaw+NygLhvvRoQB7DX3UEHAOaS3oxZywh+My2QtFWRJBVnO6xZhYwNSzC
ffqjXJQGq7ZH0ozbsNDrOghJh8jeQzyC63un/Zneu6RzRQRIcfuy3eQ1YO8cTDvyQvbfXaD3NrnU
fQO2Oz6v/qE8C41gv1d53P8+C47Nusbefsf/AnKqVW6602gdEho+kjyhnGzmJ13Ijr/S6UFw9/xN
bZFWkP09VNbmXK/1x+yMOca/AlCXGjTX02ULD7PzvZyLCXDNNW/OXpIrHkev4W5Meu15zJiMa+Qx
MnIO7NNjp8foxSmh7QyhPZiRfEuDbQAIOKjU996+G5rhAP9IrUx4kohPHx4+HgD2TAVN/kPAsl/6
Vih9YhEqn8vuljzf1p7E5jrrbykcFSiVdP0lT4x98UB8Cfbs8HX5QwSKZSE/dR4hi3RKsIeHuZVm
7uysL2iqgwgN15XV6OaJPkVbcMYk7k7TZApEOmsgwqkBMzLwERbpATk1eXnjRivVFZRiJmxjs/q9
DZNRXrtnHEJEO0L6scuoUXM5852256oHPNQiwPJi+MpZ0kk/8z5WeePocJWW0XWZ6Gt36OgStfJh
ZwQ563B5ty6/KPjI2c98lAFkffJmnQc88cbsYdlOBKHiBlT8yd8Ns4M3stz97/ik+P4G6BfN81zU
8Xab55Qq+R2yaZHUaxchI2DnA+HW8Rq05ka75xEkKyQhx1lEyqLCvYJNfacFJAPS5ihqFT6Z4CTx
HvTvcv51RgwLOqdvGx4RzOFA2q23ONnuM9Xdn7WLDHpWXD9S7vy9CtunslVsKJjXAZhMN+7X5JVS
vwdXMPN2ucY+Vk5e525w/FOQie4QF+E/m/H56VtFdJKPq48ZVfGCUN6fc1hol5Crc4xeWjLI1jaQ
fuBnlDZZNca+5FIJpBdVtDIPzo0mfnlXNBTuUl6lY61b3YS35W4TczLcPfgD73IIMiCggT9H404I
cI6MGtT36Ypd+DZZyN4lgmEtpSPtHLKnbhn1N+xwv+stBiit6lzkXj5EzExF3T22W24FkZQVt5Ak
u+9r3gGOVs0KjhE21/XbSMYgAd9oYzSl23HvyQnx15fx+vKDD56wDjWWKPmj8VpsHAfPDon/sX71
TbDquAdcWlO+uxjNv3fp0R9H2VyY4kA05I/W7UXl0+6FK/MTHOgfquwraxPj5hWim1JmvySZtSyD
b9NNEBSU6v2JBq1KVEPeNcKbA/qa0HkVnxfX/U5MZnRAcXBFkLmvIaH2WXRdaooH9BraGZtBvxBc
5ioGhCHrUZt9ysouRWPEpZQFfwOzgxWz/6c+OEf3UPdFOO1f4ucSr1eB2iGvnmAMQFrdYmJ7Zpf4
98kNUO5IYyWRUaGvTW9qG786lq8ZoZtUiiDZsnrCm8B3BuSlRPciqnGhnc0P4XE80YaF3rO3/4/A
Y0ZOYowMKVVLHPwfV4uAF3FYzlXmHZE+odA8kqklbpsgjW84eG6XSKeVFQyuEUBFmUqkcF7VJ72p
NrPFfuMs6ursUEmhQYGrdit7be5XlL16IUIrLxRdyLqgGldQEVbJqJgrSQAxW7PN9ZubPKXtc9DD
nIUkfgGsh1Fn4Tkt7jWGScIfyYWSGUi7sPJlnD5xQ+Cewk3zbtF5GqEuXHjHyIW7iN9k0Mtp35a0
OOwCdRRgzPzcAl90JGT/2HlW8i4saFfWUKpuea2zPLgOn6sR0bHJsMrgYLR7SfWHAUYY8k+gNUvd
TMdBEmyW7q27WrBRQnentqH/ERFJnlRuFHQj4gNpFOYOeq//wkgZ4OYHsJLZZ0BXJ1F3DaTBhW40
Pa2PaP6DBlazHsZaW3FgEmBVo6X7DFNp1spz0IwXY/VFQ1Dog+K4rXypBtwrxEiy/ZpW25Xuhp49
RU8n10qUdKH93RSfarmBnEKF0U9SX5dgLVDO8QCIPuziVKL8w74Vo3yKoznv1P0e8CAOZcKE+c1c
+/amvV4P3BegH6vqxzUZ2tKpYeJmUGU/aNxk8xIB1puGjlpximtJVnVMKPc5qiL/aH3mZis4JAp5
BK3irKv4jhGcq4oRmjzOljw1X8kVPP5PLMtEsLoxURdq36acC55yVhGxJLdQzjgkMh8fF8XT4tkA
QPfIHfUwSGebO8czqzu+IsGsHXX1ZUWDIkYkqY/r+mrIeXanZHP4UANX8wOOkcl2wzB2sjM5HZev
5P5gdICFLJsVixiXcie6AABfXhgpUbUa51pRsJo3nAA+2CcVBrTI8FMU0QxsKJGgiEkDG3Zzd4wH
acwGFFVx5lQsJURN/LFuC8j6b/Vbwivc/362mmqzmxr3/P7GugLxUtY3zbyHupzwcBvFj1cyjI/h
Bhm8mnlN00EJNDm+5AWignyh+qvGaW1Ma+s55jBLP6JCtqFLTtweRiy0OMnC+euPOMdZHgrjrHZ9
m/nlx/KSGhpgaxsoTLmppPDcO9H2e5o8rXT1b1diN83pkC32duuFaoOOJwP7HhVS040wQuzctgdo
mbxoeutST61U8BZnGgts1PmBM8tQmchT+nRXm3xTLXiVTn03eHtWIRkyDLxAGh2xW51r8RfglP3e
OJPWCAcmOsnxtTO8Q/zOgGtX68wr1uKaDozZ5qrkkHtdkur/RMrkpiJenojjMgwkaHC4QtIUiLRE
/2UR504yyfS0wf2bglxyz0izLI0lnLFE2D0+AMcGd999MJmqFzcqaVK96uW+rzrnirH/8FMJehFO
ePZynockE6FMXiq0depJfI9s6Wg6f/aORAUr1xlbDs3BsH87Fump0ii0e3q3ZZgKKFRdisYLRnG7
JBO9kWNxXcWTlfvIHFzcXXaey4AdYs7OBFdU2pJ+4ECAWyKnfJMzLxPPGmlbKd/W6/BDLivADftX
r0c/vmshWTt+lvhV3u9kM1hPnPe5w7oWMA8VXa155oqIQoi3MGlVBvIkmq8xiYZzbW3T9z0FfE8q
guF8Ph8au9l2NFFW3a9cZDK7Cct+UNOS5iSJUqI211tI+hU9XhmB61+EYWuY8cs1gQwmI7uHQX6c
RjSN/uAQ2URo8dsREYTZuucazqDR/A6OwTtxJT94MI1kc/P7edpOiWk0+3NXXGzSLtJNJ0Tgk9+z
nkSkk+018mxqMXgJ9Ozi6Lk91xThzWCllKYLa/bvu22ekniok5IlaNOwOxcyQH09GbMDInAdiAdY
ODo916/Tc/GM9qeHon66kXVSIS85MgaMGdrW2o8Xf4oMZ7J5/APfJBbF7e9w9srOtEcpM/XLm217
OgTZXrTj883YzbeXNox086lFyinGwA6K1rjb8Huz65FYixE+cghh8wrKQjRWD0q2WoqIfvBUnmwt
0Wj7rJX826uDL5fhbDghMQ6qdlpTHU1GsuOzReZPQWm6qm3DjGGgApgRtnJNgP+E/2DdkOcucDmo
0UqRMfAp3AsWdHW/zbqFlJVDavB3uvIWzIVv1BGBDuH41x9kXfpQ5Gv0ltHauDhO+yOZaKaf0Gsw
9KhZaV/+2FssjbXCZy8/7pFE0+83b3kjMoj9ybIKDs16ENBx4gT82ubY/P72UwvlbPsYjKadk+DP
JAFp/0FLxpG7wCOcD0X/4rL5kkn9c2JjmIbl6N75bUSLIUbgnM/6gh8teMYEtSH5iZRSuoqRcTIX
RtvokZBw+IcaVk68WhD/mQF919FG1UVLHk/r9OTJvGRahLtJZsL+Tm5rZu2aecbWwjkdIwCnTTXu
CHOTXrpu81hzPk0o318lLfpWmnmDJ/61SOslyGZcdSaCVSSTbMWxltnAB+cpZz91KwiuLrgiK+cs
t9mYRqYWE/pEDKJWglVVUL4fZCU+iozilzyaIx8KEFjOGskNr6QZ820e5w0wjAGTGJLCoh9AN74F
RZ7gwPOeXXNnYb1nor+V3kFgUZM7KsCcbJijvHd/NmTdYbHOtqvZUyN3DybrzlTqs3DpCXRr8eRg
9b1snEF6FIA8E9CND40/3unKim52RPUkHm9pbJd2u4wu9TVxUQ82jnzMyK7te2+ZhzcOVh/VFngc
FyyILIF56J1zcfTN5yEx5eI9346Hv9bEARo6x8xk5gAMxRRGSAYJkMtbqqzz6weozxS6zYhUzGrv
+qclivmqFL869S8WiBHJ3ih6sGHhAJ1yWksIw+d1Sua1B6I5+O20q2i+fV+19PKXgPYWTm1P0oK/
UzsF8+pht6ldZDdy2Ie8c2nghgH1wTy4RqyGkvE1jI237X+Xa/uPKA7eWzL11sJm4FfeWYEhmEN6
V1LW3ab4tSz2I56s6CD4I0KT8EejpWwrrSYQiZs4IofDdlvsXLlrjK0wvk7OHraQJ9bRUy8dg24d
G5UmSRTGpcBmmUiHVSnkdR6ydafdULbLTNmFLfidanDK1qVHYU1ZMPbgrFr4mmEtaZCC7AWO7gls
m2kEXrGVpH33SyCmM+q9eX8r0ho3j5HuUcJU4Qk56HHGo3ehVGgrkBBOe1U+dE5rIq3dgrkiyLrG
6CncSaPbHxVaAmrMVYH7CrD3vSoamljdOOCleNX29jW8vKttJ1Vefbjgfq4gtM0jFo5IYWC2gGCF
MuuHjnSIRXI63uDCyRu7FZ3l8k45lkc4it2hoLvuht6n9B7EKCB4owAPLV3FoL5zIHjpYq1GyeO3
SUHvr0Beu/7wPJCEeyzObVKlgRzrjdL0BEtFpK+9AQhBHzur5/yOVlqT8qI3aSRIyeCv0zPGMqb0
cjJAVGO+5dve14Spon+3QjSI+9V8ChC/ATAhZufomgaf6B51Rrq/AT+Tvp/pGta9b1EvnvhFVdw4
8WftW9qTpuVzQcucUck/W+BNXHExa4rzP2yBwmEsOzTUxwzAzzXd57tFXvqXwhBmo3QpdLgPaDbx
+Bcv+cimHuWrAcMAEsZayky339wvEuV6h14puHeLszt8eD+7ctQGC6qXa1H7d6H8wRpg/NJj1yN7
SCpVIYVoMIOrZSInWXFPrKmzIDwoMr1PLcjAG4PCDEVLeB8EwbDBJDihUz2SvF6hqqn5t6jbukXC
MMsRem3KbMkL3ivESpPdfQdVYlbB7CRKwshu3DNbeH8sqJb7tnoVasM97LVr2Vr2RxNlI4d5EyKn
ZYNwHpFSrSNIB1hqNUm9fhyI/8xFByWFNSdo0Y/3D9Isvot/TAZ+XQY5vFJsKwQ6mpepZhseo2aJ
eeIUvwgdyjIfqzCtnCUQbdZzjt1f0xn+p4drhI0JU//LXqpf5HgeBh0B+oCi3Y5L85Vu0b+8fVJ0
o0axSqri2r6LQNb9jRzjbwSApI/W/Pdim9nR/YE6rNAKV7T1zmGWrszFy8BB6KplOkg5WxdQvj3m
LYFhOGu+yRM0HBJ0h3GGIUURE8w9yZJb4mQOU72ZQE+6gH/t17vvo81TpAmWyg2kwRhztCjHa6Yl
L3hjwHwFEGzhnldHBTeV7CRAmZcx8fBlwSsjZWUpSyBhSTJxHq/+AVbk2Eyx4i0053ItsuvZdQle
ZP5ZAqkc4SHOnLuGbgkkM+sEManytVS2NELZ5z1WfCHcYBDxuGQ44ahrLM8SO5DSbBddS69njd++
J8t1+zS8TQOAbDo6K7tET/TaVCuJ+OIOU0rOJ3KhIX+9O0SgRW9QwPoZrbgelGNpySSpuUXrk4MP
I1tCNgFgTdsJ7CqaykgXXk0KOz+qB2L1OhmCut8mTtnuDr4YrzNabT3SLTGHVqyBxkm0R4Ldw3hV
w+jLWxo6tb5AdAgT0RR4ScOpTUDyIagzFLbuG3cCBeSnlJc/uPnwrcN+GIKQeFslUy3p/Fn4jizh
KNxQE7kH/iSwsfS2hSMMoBIzoMEKp0eovQK2UNc5vzodClUQxQ3Rm4ztSxDO5JlFh/hrlH3Oxn6d
eTBYgePsRpDxmFDRkxSU6TLL2/qN/xB+wjDoFITusYOeZuy334RE0d8VpVVvLz1YpFnXj4KU5LUp
/V6fZhlYTV29Zk3GHDrPSKTZgeQAcaccUjsw82Hui/UU6BlGKgl2xvDzV+FcKfhpoeCxvLy171de
C7CG4ZkojO/fLSQyVTIx52RuFWUtbc6S9cTdPAJSI0s3HYl8fBTQxz8NS/Qd78ICfdjAbw1jjWhD
Xi4ev6q76WGY4OGpwzEs2KGqYGY1/ZGebY8y9Gv3DU4NazBYJ3WFEAQluqgd9XF92DKrHNQJVkGL
+OtoW/9+rd0WWAXcqDURYtZee1tVw4MYSebmN8XS5By2LxSD5lwW6E67+W1B2OAbvz+7OEFr5JkA
CY4hjEiOixVqj4uGA8qNHzR871SpY8D/ye5yp7c7Db0yPTVm73Ov1wPxSVBdPsY7P+jQ7DVv3YQJ
OjJab0Hbxmwu/0uh3jgQU2/5UqA29vnOX2SUjjJoYhYlQnZVgcTQr/a8WFsAx2GIm0MuGt4O6pY7
Zi1ha4ZOUo+KOVsr7HSzju6YuWIeHqFdGX0mKwRerg/LrzTlybKQgVnGMGXSTvKbRHOpGjJxaM8G
uStiAQjTR+vugn1ypvB/7jevUM/zykJ0URnoRlMm9H7rE90xBvgXw+ViJRLnorhvUI8Goann1s5o
NocAp3SxbprzjVZmdB1L4AXbp4ikHV8T2KB39CaiYf54zKz+x40mi4/m3YXFa3YxOp2E19kvSSTe
/f9rRsfRauykMTjN0pNM4wAChlzhiB8knM/1OfqA2T7fZgFalNx6kfntPS64Uvtjkln2D2acGMWU
rx6CSXUFb1ei/hA49lGx93iF2z+z672HN8COw+rVQBu/VK36KwSINGTLuyS52Zs0BMswVTGMib5F
1lRVo6C2uHEy4nJxhhQEjFvirSYXMqRfX+zuwn3WraUQAXyiJEXNH6ecXDSw9Xd8Ri8n+wjnJE5u
dvPsPJkeRKausBfpJgJOxpAUxcTKz9YC41d/Jo/ts1MHHBdvcMv2s10v82HMXBs2G7ZXg40RxYoe
VobkULLZ2nTG2e70SpAbW6xI4SehmPBsrOIoYhXkbZXCWwwNzOFoxg+gbBvryyd3VVR2KwP9QMSR
E16z5Y8Jc7uLHw8gqYQ3nFo1VTXncG5MwGMWo/yTBagRkpm9dGV5yUzbUmGu1bxVmwiuObi2HUmS
Lqj3Z/oQVlxU5tfp//K3wKdYCelvl9C/uo0wZuwZhDv4107xm7dY6hhX/rDrjFBkdu0l/0wjLsXQ
3p3DZ1vYKogdBYKEmlNGOiL4lDNbdDK6boZy4sd7F5dqDGFyLUEImiOG8UJnkhIuOqRn7f7m2/bR
7mWD+1GuU7myHODBb4Zt/KLucSoSZNxxZ6liy8VyD51YtOMocgf6wGW7WmfeR9hsz2GruhZ70uV+
PDtxAHRlPbsMds3VbM/YPtgtaRHEIE+dfvRv0U/reyJ+8q1hoQ+DnH0XYLJ/djlHp0NxqSgkrj/a
eHbiM7fpFIwa3PvI5KZYpaNQVCpfh+CuycJw6ufqmX/QHpWQblLMPg6UcKKbZn5ct/BpS9qkZUts
zD4psgTkQP3GwlbW2LXIWBskomr5KT8R2ir5NfPbgC56baxq3L7v7W+A2Xe6OWO7krfF9N92ivYQ
55wRRdxLkQSF16mSNafGXznZbw410ogxYvGs6781BpqaRV+7UMWn3VFucvadhhreGF5EcNCZr8W7
Cxp6G+rvGB+W2yFyXQvo2Mk0f1sTJRfCijKg5B4uVWfhYPfo0fULcycmeToEwPfswz9hxc9l9G1B
SBqm9r4fA0leFmYBpRmxdvW6A/rIkG3O9rF2AvcNYSJk2h2BwPmxLbuLIQbvyC0lKNN75G84EVoH
/QXTkshVCQzO7fntSC+G9zAyMMCMxcGN8h8RActGmuHihkxri/j2hayG/eKWdcNIYgMqq+MtoHpb
DC/2HAa6eCFm/HeLUmZ9wwiL5rerSd/gy90uBAToAgn+UDsx1kRAFeVSFlk6IC/RPISA0dSFBxCh
V6ywQ4AcIBtMo4ncJRWIX4qUDc6dXJnBJL/Q9BmgZ6hGdbXTkWYuQdewC4wUP2LJagad4HjFDPbH
ATfiP4btgrqaREEmDpvmXbV19Wf3AgFRnJt878iOP8l2/HXuzDwPZo0BL+dpFDo5+bPHnhZ0OT9x
lmHJU+3ASObh9GU1neJAJozvArNTq8OqK/I1L7Iwjy/B3nPtFtm5Cd/+fUAKtFKJIHp18pgt7zmS
yXns6Me7XvK2IAo2Pp4J6mNqR3pPIfLGmW7JtoZ6folZvkgii3HeguCfDiSxRWyv9U9ROHIyEXg4
CaYI+7mcOwXnKY5zAzz1EcVzY3bvV/AetNxMtMv21gXCbuF1gCM1jt59ig+Z3a82FNg4AsuvBj5S
foxpLsTaUX6ST2sVd1CP3y1VvYbTHXzA0D9APTDqpEmq3fVP0KNL0FN9hIbFSW2lmUrh9g+xu3p9
te/OTZSHHWqJYVYy0azsKi1LgkRK6I4vUHzimseoCDC2jVLUjrwE/hDF9XyOCABi7pGqe+WbHTrf
O8xSziLa1txh7x0hKcQEaHiHAtEdpQevBZ8OTw6vadXk6nwnSVAphZc7xjFZ5kGYkISztj6OU/6r
s31DQYGfMwMso3CkbyzzDjDIaRP/wFWhhWgR7q7gt4zirKLjlKRe+aKyc1zYoheI5aCvYnk18p/7
Z/XTXbzBXauWOKExqZa2KXxWWyB7HfHgqMJP40qMPLPOqm2PzQyQQiwlXAEz0mUdEcqj4wfe82lL
nh+tH/9OfHcDLSTuuzK1zivQP45FBim7dlyBbLZPJJ8h5HWOqhp64bfu6Uzw+KKusoCvZ0oLiulM
Yy4n4VgdALJdaQRhXF1GPPqqqgOIVr9fHECNzngIddZQXBLGKlj4MaPMp/RwUbY/MVOWnqKgUjT3
rozoY2XRKIhX/i/uDApr84fJulOlE9/Uylljju+RdoUY/Irq4qLSoZ+VXvTJs00Czrp145daffqD
mdzkjV4g70QFxOi0FSyu+kBXWwKu1YSsL2g6YJZ6fO3LA2njnfQSWv80QBUCWLDXYGEj5LSgjHwR
VHtiv0RNbFx0WnFXbdM59l0buO8gti3e0U0mZO98b27qKfYirb5lP79qxFoizdicxKkB4b3XtlaY
IRiIU4NqIVCeq1O+BTHTJBaunJI1JfUA2aTapN5qw633/pkmOWCS22oQCzu/aB0TZCgn5cWsQRcF
snj08NZvaaTHXMSYqgBzHJ3hZx/sA6vubwHswTZ5rEY2RSF5TzPRvUAhwNyGPcFCKlNcWVZwggfb
Gts0cVNq25fMvlxmcRRqg6VuQZiBgRax8Fh1HODRwgXvESdgL5REnWbAswRqK1n4pl54WO+TTLks
bv1Xahh3ji6OihRrIWtHBOb7QQVxErnfopZwSMXKuIL4PtQdpFWgMzQhBhFyzL7kuI316vgqHFYZ
tbU+g04GoJtEOUHWnUa6XBiyUd75UuAUceQw05eZ4zFF217veam7z6xop92+FbAfMoUHRIJAc9Pj
zpt+7T75pqXXFd0xK1DQKy0Koj68iJQ/i0bC0SRAz3XeRj36wzaKR1lTFRTwnT99WamLh8O1IUFz
iEEGgFcpCc/dRHHFAyf7jFz2LqoLa47nMULsyA1cSSv6g2vrC57J1OjUMWQd7nG3VtPkCwATrF2O
tdtpwUftBjJwvyMEJb1stfpXNppjFs2VnTfLZBhtwy298EjCeq3BTC+X6SuYwCLon2peFq3rZo0h
pZwR4gU6w9TBNmQD/IOBosFOIAFi9pKccw5Z9qAylHIfOgmrjk3kfa5uuH+B+VIKPguEX+Wn37fS
1FeqjdR1b1JKUUgY36k8Z7ZyERQgLcsE/jZPyTkXwxditCTHjnhVJ6ScEAQAhqXAliwOU89VE/lK
ptaw9ejamZs87vbj3XnzdCPvDnEVyVXZpWtVSnym4V56I/qzAJR7J4AnDuy7w3KkUpyYFKOhCMyi
I3iM9pLWYQWpIZpbRtaYUEfz5Vk73x782DgQl4nqjVqwOfdRhtZ6oqdIQBljiqaI0PUj3u8VBsFB
2/3013XZ3ZsduGuTQl+FHOLuobW5z7sgo9Aqu8NWShle4Fgrdx/mbO2+uty0pIGfklmJ0iVB7yYZ
2CaQmakpMD0DcfOS/eIvG7lP8zngo/RbB01ZIARgAtkWDHnOZHRnfhZa8FHxxBGLFc88iB2aOMVI
IeYW2mntJeOFjpEQQO5QvHHRAi83FbAJxwnuMaRBUL3S+Di399Xr+blhjELuye7+4Dc2nhx19NHi
YEO/0hHjxGKkUrm6qMzrIjlPQZ1+JaPQDSlLHJgEaW1sEyj5HSHJyCVtkmA8XggZXxPld237a/j6
lTuGwNKipL2t9MJtgIyZJskFOMG9wZkDT1phVzmnX9n4ua/8zkeazGDKSLthwRviEI9sY26lofKN
rz9gX4Hj1mG8CwkjWmQ4/F91gOzerUHxsKmqzOX2VPJAxkvKHrgm1ZGJA2aHBGW87gkkgH42eL4m
OGysJ2CupElwGTLsNG+onWJ15wCSRMUoQOna3EfqbGDPcCg66YU4txNIMOczBe3FIyGk4VJBjneR
n/zgkr31a2YWx0mcGKTZOIOWU3q+J9JSJz0duwtn1X81jmLmNhf11deYahyNHhWLFJ6j8pJi+Rcv
G1Yx0aJMYxWTTuZ4l7Fz7DssGpbvMmR2F55Vllq8J1ZV4Ytu1fO39nZ1BFVW/+sOaZwF6s8FC3YU
Pd1F0KIvMx6MCBypCGrntGd94N1LmxmVqIZQ8EAqdjkyCp9VwX6I7o9C/XCykbFPO9s9Ntjo5ciL
yqfjgvFp+otASl8B/UozBo+Inlcuc1FpS6f3EsfrxLgHYBLLGFJHAU31a0fzX35oG8c4HH7Km/6b
SrtKNon3HLXzaryJ8fegiixX0aZho575bZmEbZSkDOXlPkl/nTUdc5yMcIV1gxCwc8ZyLYWzAd8I
GnSgnEms8/hYY1IWuD9acShIYCUJQE1gYy1dJrQLCxbAVL0TmH4vKGERb7lBotogDqoqoQUoSxIw
AlbwE++Qgjn+HryVNrItPnKvgf4eR+PJ/Kn01nYBDHYhy9Q0+3voGApvnGbHvvK3GvpOYv/rA2ly
vicZvDBXi348UN03OYXtTKvjA2jPasEK0nQ6aex3gLddZc03CSvNbbx+CmXHCIeKnIjXi0sHhyOM
CvCVKypNhxZhcP4XBkUExfxvuh/N1U+ncYOrA2RSs2w0A0uzEmSYoiVFEX7FfsJmiSxEaXZf0mWd
rgOw+m2Oh9Ah9Xsj5QNA2EVmYC3NMSUZvvzJ81i2zyGhewN0gdBqec9NQJvqA7Kl64ZUORupW87Y
/GPhYAUYZpqyi468NOZ1/ULM8j4FuxT0roGY3bQ4IL8tUX+wWvulbqlgIk+0ar0zfQnTqhv81Shm
ArzxbqAAhdtKVq4N3lXmn4rxh7I5ygHT9+J0/5VZT3J3HX5Qu73byVgWvTINlqQRwIRysK/52fhp
cAV4Vkp5x3oUCp5oCFQB+HFevzlfzkWNIOfpwHSTv4yQxOWM/XymW6YUWIukAw6MODeBSgJFrQL+
ET2BYVHe0JW4J0CNcwfiEXI1H0yCYoDJC+3j+XgJLVmONPcONmusyCKrw7UtHWxRbwsfmXP2MTwF
WtvpEppCZYR2J1EwkTi+hvqmVy5MhwbunkX9Uts9nFF46KwMnmHIu56IaI/FZD7h4T0kwEE97HuJ
XBafSwHsskzovSbHxUnUnVZDmUVf9H36yoDVl8OfdyPSTonmfES6HZDkC2TMT/t6Ep/YWcJc/Ovu
TJHu2SzhWYMdvlqpvFkms4wWGRvDdH5JplVtIjAs2B2Yfe8WaqwyUwMLN48SdD0iXWpocONyMUg/
Bk1kSt7P9EtGAiMJFDgLAKvJ3a51P4hnnpFVeJcp+1AhNYi9CLMIdgHZhC2o5reaHWYkCHiXBCAH
j1uun/g7vhTaRQQen3xXgL/htWKRfQ8O6E3kA9JsNQi3dy0ijx0e0qno47/8AXYTP11Gpy7qH0Kw
VMQ5/gnn8QEruGWamSdNyCVpDiPom4uNwQ4LZIGgaPruMq0uaXGFwr/BgNJc2ALP9VBx6rGp4bcI
b9EcFbNbD8Mn/ijp2FYCNppWEbXnZWnjcYFY6LEBYN4mznxKAg+a1UiWc/s6/AB8KEgt/or2Dd1i
OXZDqJPh5e9gXEIYvQaaXO1cK2vORdDNJITDwlRwYHcOooUSoW0kC8/4KPj81Unj8THa6X0M32Ly
xRvs4dASUjwIdWOBDS1Q8godnkdejitH6tt8hqgOBelSp2v68uDI20pX3Y4FOKW3uE10SdQPoBSh
ifECLBCxPVK+MPF4GoaV5ZA5QByuFM/jWcD5Z9DnBBtvOT/xXK9CgOjjW9/B3l3DSzoQEZq/9Zsy
HtmZAQ2cyCHbP5Ndp/rmp5QxNacQOrLuDbDEVINhwEIOj4IyyLvNMWnu4S2pC7CzT+i3kG/DGXia
s6SXsd98ZMiyF00W4Bz1PK56Gj96NbsUTs3raDn0WNBRKs4TDZeeCY6XTyR9/IqTGaRjY/oCYqN/
bZz4Yv7xVh3pz/mgTDKyo/uI6/WGpqFvPRGQxp+wZlzu57r1jN44856Bd1Kt7dC06jIaDk92pVBa
BR/9xzAIvZG/LX6Ao8kqEcnLn8QH5mS1jC/G3twoVVAVqoAJyfpqqC+UFMa5ycnokVAWx7P6unzG
5he0/HR36SOKA8zF7/WcjR7FJ7nPSBnZWFGEHmfZPKuGjCHMSBjcnN7QFc4mCVYc3U06z33wA+mp
5t+iwiWtQB/CSjgDDZFHwbgqMroM3iy9dJp+4gQ179fs27KYtIOdiWtGnRA1iNscj3w6baNggMe2
fa7LmnZAVK+9oWpXSCcGsSSmkv9Idmg/6sMsO/0rwH7xSMdFNLvx/dWdUdSkWcTsaKIQcAsHhV21
7vSX9rmVTspSXIB73ECfwNmTcP1mnKklcFi25Js+cTo3pIoU15+eRtOEWqctNuIY1BrIOGbCMeMr
Ixk3FasdtIXLUR83ZRYjYSJgwXO8/2Sm9g+Jehf57zbneEstCHNIKxpIqpEdwAStYdMuTTnBvdB4
LjGvJtPAL8/9PRPPMDP1zZVfVFZ03x6Gu/pkX6uXnmNK5LJHZP8VKOZNB8CnZxVXFdX9K70oEH2L
9uxVYWhgM2N0DSNaCC400qGOvCiPBtnDfmvabeO4/Vlc5W13WPHUHgKwB013S17hLPC0gGGx1F/C
3B0gy0+umQx6g6mpsbI038DPJ5m5YmcR69t7/oTwnOwA9mcBFpRgdtuwoPukzuWuv7ZADTlnQ1/h
+YKecolWgEs/8OAOcmmoE12Dc1F3SXZkjdoaT5KXE8kGVdl0zMMS5WZjo+85uaVAWxqRdiie4jdy
xpHtB3F+DzvgzDPeUP5y/ZnQL4XfpMnM9cLVQ2RqfpKyMjbpxioxTiBZ35bHV4WxgN9gyFptxqNW
ylMPg3SUsiTYhgNZ7LQfB0FJkUFLoTGYsbE1tjI0Qf4JQro3pzeKyvPsmDblR+Kz6n0tK15kHQrH
nEHdQujDJNONpO23saSjloNC4uXduYQVIf/cDFrSo2WuuHx/wAwUSrcWxrm+53PRRWQsQEufWnnJ
gqeU9w03bPC1KNK1o3BzDIgWWRKydTSJb0NSo5Bsd8aJrWtf/Ao2uEGdBCo+y/gBsNhHdFZhuzd3
tMbn05u9apB/I2rIdbZJiL7+uLZR0fi08RvTYjWOYxb1bC35I7GYfNnJ4SjAK7t1baSkX9twWNX9
1PaIzhDMglkrvheLLCIVbHLmsDNRXKewucx9cD/h6IvF0nOeBJ5Y16kyaMfuFUfunc6VEkuECqsr
Jna7JjxGXLE7yUj12NkH9rhc/et2rsrlLM9R1s8IWC6WbCupvvlKZpFIkg57QqRQXiA5u1IPcvnR
nEik3Yr6AE0h5OvqAKhUf6KoS7EDDESU2W44Ocua1e9lrQChh6MzSYD34ogXUa+Xep5eZVBPiVkq
N7Lz7DgfU4fpb/SjYLxqY1mDkvmZukBH82a1NIZ/PY8KEV2QXQlkJcLN1W+H73rsCoSbhtOVeiJy
sEpy8L6aH2c+Ilw+QKkgpbSjx9drB1bYbwkCPyjX84mVoiEcnr44DjQevLH7kwM51+i3g/copqJm
/RfJquBRDo3rwl6OCcQVCamoCKzTsr/ZPBFO78s614ZPKug+2c43ykvxDVP8ATCEBNYBxb/7Jl5q
NZtdCQlVre7Y7qdKxQlhJ5AvkD5AkwYoJuPRvCRo3zqlj4uPPVUygPLzae8NcJZ5C24nYNtudUVq
gyxToRl8fD64xpBXXue2iyGgcdC9f7SL6LbhGVWRN2jiNE1kqO15y83EmHTDvYYlUOytb8L1mx65
6F2SxF60ZySNigBHHYJPVL0ogaX3ZHRIJe4eOywq9lYH6967kaa2rkzv86Un4rMiEfm+fHDhLh4j
WP8NCirKbUBOQipckFJzkSJb4zodZulotUjXTDpUfs2sdS4zqbXmXSzBnpZ0XgdMN+WWf6tdKQRg
ZdVAnOiQwWhSynmMjTvUzNdhSpbreGI7FdJnm1BR6mAjDYUWE3w1hFS4zLt+AeJsH8SOcbbSMicK
/uGHknX58KfCJcosuUNFz9iERYmvYcSeC5capItpeLRQKkLov+HnzYaDjVjiBGkHkb3217OF/vwP
RM5kwWxzs9resLEh6K76MIBAAXum7n3mpI2YPZ0U1tlNgEJGOfsDvHl98Bhdek3acRGXETIJNeSr
dfD86wllpGWMrtn7NCLLMInbTbN0YFSuHMyMIQNw4cdDh+jAoDLSaOEKLMhSqzBIjvaMR+c9zzkS
P9XChXlozg2t9ZbKG0hc69tywgOEpPSNdAG/a7zOpuGtqAl/fDvKYYuElBE3eGAnPcqK/WGwI8aZ
i3q4AD/z92liODCsmU8vfWmm+nksg55CGmT6PQZCqoRM6DdRmagO23oILZ8bJ40lwXYxQj9fahJL
8W3rL7MezQfvrd9+eBCRl/fAyWnNfuFty4jqfBGr/xNQHlYmEXLiOnpuIaQP8aNnaBxAbAb/FQwa
wNZ7yRiBiG3wJjakk9grupO2NZFb3De7UdgQDoD/aQ7S3nxnvb8/0EgZhXh/KrK8YhGd19RyhKIv
QEANQmI/jF1poAVc6V1cU2qIv6Z4hMlh2dmpsJRQmYFLGyhafMU+IjnglfeB4AtVvmFVSnX1EWon
56L1yDhGPl27o5C9XiCi/NMP2JW4b7IvVDyg9RvYglQSJBfdX+Xl7fQWULA8PZNG3iP4jYgcssyK
XA+sBhFQPgsy1O+NM1h6ndnx4kc25OT+lxCebsKRBnK6YAZFNBtRJjb2sjdGg3yNmrHlgirbLOuM
rXp+eN1y27GQVrcuREITIX+Gom3cd3Hq5AOgtelFSgM41WpdS0iJeBVrNf5jomfF/+O+6y2kjH6r
vH3eLZvKjdTy3icdp2DgfnJY76gNGWe/fK7ywABaRZMF0xfT/j9n4+vg/FzUrn9DhaL0udtUI4bJ
PRiiz796hDjL8Fm1dlFLrSWxObsBpMd6VTUVZKOBU3v+dbJKjPUnKv5adh26EFtOERnFZqCvPjwO
Kcp5tKA3qDSTWaZVRFpDfg==
`pragma protect end_protected
