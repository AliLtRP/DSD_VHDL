// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ECgGBdP6RvQm5By4NpDV3zzJSnYXgUuShHn7l4TcYAYS6h3x6BEhEbtPXRBrz05C
Qhr0wOagqBwuAKDWV8FgwRwOpjwoIyUPPDbEY9QqdS4lH2pgLejusTciW+dy6oVN
baEJg6+EqfhFO0njr0EAMW0Sqq5vXK5RgNWuOCIHvSU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11136)
rYCDTJWzm0/GkUtEZp4zuR94UstDuQQBmxQfKWyDetvhiI7mKmzmLiohHL/OizeD
m7l/I4/ih+vFj5kwy06AI/EmdV7LwPskaHyNfOiY50wr7v2plIL9MAO4zSBi7wcb
R4DAnZIBfHBR59pnc9IafZ8mnXdCxnfEGaxSA8a7y/MO79hbSXL1gS695vVzNjsC
Zh5QqPFd49W3nNYn1FNKmTlda6CcOy+c4cxQkNIckcneZ+OhmLZEgrHBnML5mjbb
pi7OHliw1W1ZbK+ko1HfJ0yeEAXq+QNwIvUQjKPP2QemFdc9zC3zwEDaCQ/oYDuk
qw7OwdXyeL900jhZmJn/pBrHan0osGCabdgbA07A31dw09Ckj0iOaXq8SkaCYi1I
LWVT06CbBEYLa8s+M9gzH+HCjSTbZlJHax3gbLTfGcYyulM3xjcqNa7eLIz6MwiY
DemUKMKIlfhPfWMa+MnzW5NydDuHHotH6+4+o3GcvFs4fmPJpNKGXL2Z8nGRWwpt
7MOoeNa+2s+bEeq5pielQE+E/QiVXoyviTRX5CA7K3nKSn81/ylkLUfoVUiHhf6r
w2x/vgpTVjeEDZYd2LuYp5kK7205QLs5oRZ5Inu3E1hK1cdpjkiFtTugklJzcImY
oVhAoPhjgP2O5xnKHloSsu2hunkipNgVPr5vQ1rBz8bngqJn4ZXsGZp4/1r908Wp
VEvL+A5j+J/6EYvWpNxRJnQ/E0a5yC+tt7p7DSjcgpK8reQrwNmQ8RhXbImdZEvk
F4PDxljR4uG5IfjuTUap/BXQ6d62qT1+STRiEZCehCfhAf9juxL4CbUDooilJdKV
tTO4uD6Mk/x64dEISD63sNDyFgIRwe+NeGIjpva4rlXFhoAItgUuEblj7TquxZQV
u8v2fSS/MNecK2/NyeWg0WR1dAc/CASEV7kCra9WMiwNxjJQyeocoDhlSeDcrzYN
m9iin5bDRNccIyktLCDO0HheJW622BfKx8aMZ/FiflfibhuHadV7aTn94660yDnQ
HHLgtcR+c4J709YXYi5KeX5Y1fgkhiq5suLCw98Xb70RpMDfwkBU6mP7hBihrvTb
4miqIuqc+z27G0gAVfWYoryaKN6FlwBauRSxjtolEAMwBOM6I3lbDFoQjmDkhd2B
oWYHkV7LX0PzgbfWZ2JnMLXtTW2LvHmVuZgI5FtsorolLCrEzNLyPajwn5jQagBY
hUvIVxZXVF+xB2unJGAjH0i8qlixvU9jmJ+JHfeTbKgx8j6QMu62Z50FoPot8bOF
ZZzjMX5XTE2ko/mXnmwyCxO41qgW+6cq7MqWcuVrA+6zT24ld2JnU31HKWv/S01e
W05OMddTHVh+IyDUWoitTjJBNss8fITBr4v8qoTnOBQTk5ALHThn4GfzQOxVBVbS
G5nzg690XSMYrjjjl7YbFrPHALRAl+3Kc6Ueia44MUc7b6sJptz/nKBCiRj1fNov
CxCwPD5bIxj/w41aqhm0CVDj0UeQbgmSReMT1gTVTnkNTt5tZN6on3HxXLRW1kzL
/+X08a5eVA56hf9tApTlm/1IVZIOhP7ZRXXn4OmZZQ6tQq54Xcrc6W7J3iRK60Bk
0E6UF/mYKnMAByVE8/Bxid+QNXvRcaQXzGZDkXNHu0jIv7tp8HwP/QMFZnPdlKDH
GdAJLIZtEaiEQ7Egry+wRzriQIR8fC27VFbIkE3OS8Yh5KmBa8r/OhcFtb/dfsbG
v5Mdxtb6frNRTshi7rnz/vq44HqSZcB9IGlRFEDOQeyV/RU4GaEkx0bRH/Tdd2vN
7F1U+mFWcpnqwOW72lGth55Ff6vFdl6JsDnNiLOz17FP9RfvmCNz4pP7Z2ysMlHw
BEUlQ4ISA6qtLsWeH5H4j+gjl5iP4KVI0n8w2aW8f91qPKkIwHOq8lyRaXvEcTkT
SG8F7c9r+bJIdZhG9PVUjeDL6TPbP8P3xBPo8TI3STqp4AODZa8q4vGbZISYFVeI
w/tMjfSgc5vDdEOFm5V4dtDTpUKLve2FwhuVCST35s4nQIcg8GtpM/VX68+YqnFF
CYlWRSbNfGItHbNI5SphMMWflwdaogmtzVccZ1+bZTisvdKAiBdNU49tlkGtHbpP
+FwjDoujD2Pg/0tVj7y4pTvlrmubeIc/eo2nNhhzrutF7vILJEhWFpWXOoIHDp4w
rd5yvqJVOqI7M1Wwt1AfCPTkygaz/hE5CDdJ0J9qkDHpDHPZzdDUlE2ORksKiBpE
/Mx5eH3YCfQ+USVxbYTpO+iK1mVn51xQ0mCGGSnJl8/f1VqaV4Ig7yDFwCDtKUPX
IjjHXck5NEVOe4ek8djci09cTr/qOL1yVbbYh2a/aT5i2HMu6e1ciMUlLWsEdnaY
JdXh21iW/WgATUIyawx3Ioe1lOh854ZYofja32jdgH/RLfuyR64bkaTI0tRApw+H
sGOFVsxDgKJAmdoaS3SHKm2JEFKuzDV+LN/TXfo6NsDj39+kVy0oF5mUi7Sz5xe+
YWNlRcAiQAq6hM8Y98eehcfgPlwlzeZ0wEgI+fYRo4K9JSdRo1jgPN/vD8YW8Y3d
1KmyvQVBnkm8AnxvFvw3xOtBl/850SsUVZdArnzqeB31xrEuchK6oLka8w2KpJ2F
ApZII1K6EACnm0wX3m4ptd7rPmJy3OHz19/EJu42wjfbITYYrBn7Vvm3906ka/wO
g4sAl636GMbY4pJT3yhagAoRedBgMB6rjjGxZ63gkmdRUBXQAoZ8dTPFm3gqq4Fu
XY+gj1TY9S/yxGOr5KVCtjCnocPvEuREIvwmPMMcrUVBPCk8BrWoJDa/BRXTqoS6
Pai2oG+ewPHc6lTc9Osuhq3l0fUgVSQWGWeo3Qr4hn1dfswnh8wW8qGc8eCTFJsb
ESxZkIDMGBLVLdSWt9itkngRJkEb9J69nGa4vGY+l+XEBzLMqB3O3oe1DM2ZGg+T
gokR/6fs85HZwMLVJebtUNj6nwRsY9UIFcaa7LlYuHapaQ6ZBriyWX+2vjp1btnZ
J8PkdA/dVb4Qz8o4APResEuoq+ztly579vPNvgt447AIrnEuBt6SdOrnjB1p6Z3z
+3nx67vtig/Xou8S79DVzmAI/MUIhR1GYtBGl5bc08zKg8LJy7TTWDMwV556fVUK
i03DebE4tKCE1sSiQsrt5UXioOkK+C2VvpVLygQw9XvU3KUOdK84geD8D0ZzDEDm
QM6EnFdhOhlJ+nzM2VepQysSvlRsRKR3SMW6A5qgN0cdPOflz+DUK6QF83DEFXML
8c59MFrXMN8RyxeojjsrMy0fjbfqC/bWoylKSTRRliJCye9JmhR5cDxqESttCTuz
bX05oW371aLLVAZpkM23mz9vzZRN3CHcJDo3I2TmGLgd5TkVAXsr7Og+EQjyVS8R
SZW5/H/eSf9MoRocyJHZ3iRg0btStztl474EDdfFWpz3yfR9nqY2wsbCDXDbSlS8
rioJ3cw+K62yEwsLjEf4KjVLu/f+MAq00JbXAkJTcWSUocYPuDYz0xyMDoias5G/
Hqc8FcvTVk5AIIVDK1xMtS20dS8RoEDRb85pmBP1q9OEuLhL5kX6e9j5vjIHvzXu
+vd0LJcCPwlmqUD/KVm9DMV+PmD1cNrlJAiyGGOLltyqEK2IPDHq+1n6PD09E7uj
UGa3IvVVBHKFF5rhmCtDOYTW06Nw7nPD+N4B2ZmvrmK9uDyJL7UO7ZNO5ef7CtYn
NLN/m0CSiKQfB0WI91Mn76yhahsPVmaziJXFpLmPJr8aK0U6fgndQrSD414hxOKJ
XPgexX1jShV3JzZv/hjeBeD7xwBlwSaVu71opm4il/IFGha6Yvu7SnNhxSS/XvtP
g4EFluBDuQpMD9Zj5KnnQMmkHrksFURFQUOocNaBKOkXbnvrPdUchJ8OVMiwlliy
inMuPs+ulAM2FtIZh1zAZITfqwJLgwvPDH9GFLHDb7ETSz25JdQ90Kvb1s6+LxKw
Gk89mrJcHucd2P/nKCSDhSO3mYTYPs8csFnSouCkO9iUX4enD2PeJTsUbMiA05Is
1DVHNfQFVfgmjIq6kvtYvFMe5+Ya55imZlzaPi3EIjgQMEDQAr8YMRFlwpPro17B
uPIXQsSZlIfeAhIZCvJpU1oNYmzaLBvtFWRfvoiyXLRZ2MflCvy6pt1RWzltevHD
fLnQp1aZYRKGuAIrSvPPeqaZM+xJteju2N4oJDB+fKTsAxIuCXGddf/A+QBKl7zw
6ekU5JV7Kt+WdV1uwIait28uQG5ltW0rqJH+n79otAzIkKmZXeF9QDL7HWB2wEKF
ACw6+FYyWa1Fk2JKSje47ZKwRo3uwmlqBn2M1BDwAD0yzVeizHMayyM7WipGdS2j
2QNOoKTD3ECp9ki5IPTfC/yBk/AHkA2c878iEwCibaroh6Oj4kNByxmJyX4gjpko
8HokoBwrc451k0HVrZkzgU9Xcq+23UG6F0O66N1XR+iHgGEa8wlnpsi2l8Hnqpjh
QCP3GaVU7t4dSIWevPILmNnAytkv18hmZ7s8p9GTiGTl02h8/9F5WuGKGWABAcC9
AQqJfbb4mAd64qq4vh7sJ3gAopQ0LSsV7uVXOi2grk3Kw/iQM8BN7kcdDlnFGaW2
5fC9UySDbPBfTh8Yk5xrJN7WionzxcIB2HQMFW77/Wz7tVie+ETMi9eoLKeu0Hut
rGVybIToB2NmM4nZsIpGaQ1vYBihN+mfTsWn9hxShetDETHIAmxvSMnLcOtb3Pn3
qhgSZxVqS8uAOnbCmzDkzvxpEDNEwRZU5xct35qeplvcTmD5OhetWMzAe9BJKt0s
Ftbi0TZHA1U+fzwbl6nUYHkkmwmDRQclp0xlxkw7pXKBf8uOB7geIMw3NouXmVII
z6Xp+8EBomD3obNC3f0rBAgMr17P+MC24v+cQQSKsRuw1Bq2vc66Q9bDcZqdjXlp
qfHrpVrUcC4Kf8K9u1KdW0IsBMQEkJJ1KLJplQVaxVxhnDhrUMLeqvdNceYE0hqG
WtfTBbCKC4tj5SuitMjIBdcJkAW14p3JKSG8Bwd7Kvx+dmpyUGDu1sA50IW40WiS
uL0ppzCCIMcXYsLhaQITdPKVQUelgWTmIZ90HmeaMPmNZe+tMLnS19siFAdorYRV
VhygDdNTwncr7oJjz5+0I2daCkVtoql/63bu4BeeWgi23x5te/eknY/evXGxZz/5
v3/qXE5/pJi9yHO9GQ+4vkflIaEkcYbIu9JCpA9aav8Sp8Q6o3jKTmseXKUYd4+z
un26pJxso96ABDzF2pnsu2lhKrzYS56dHuLJYbPfWV28mVAu2S+7YqjQ19ypU605
5skO+c3h5NSdBF1bPzIbxv1cWHavGlRPRGNSsF85DpSz/OML3z9xVq85CcrlfNBF
yNSJdhu/xusroEi3evSw3720vWqhwyo5LuXBP+9DkwY0hzJwqzFHoEoPcmIBDUp7
hVchybVqCeYm8B3FSKq3en0AFnvyaekDGjgyTV15IgqXesNSR6Q9OSzU+kTJzsZD
6zyXWw2Fr4p4ifurMha3QuYkVx9lT/6SJg6/DDg5H5x0UtBhcFutcmhloidA83Jx
70eYZL5GZX5/5q7dO8FesO/r0aq7OvqlebZVO1LwcUz7lvgzd8y3h4HCeY/mTyAx
JtgXOymwFjF0HqjpuDII1qXDZp5yufhg70shPSjpxhswI9D02q4LcJImZz0yG2hd
fm1qcaT7IChE20AKbjOkWgaeVxs4XdJhyOitjmOTzvjy9ZcqqD84N/9PqpTICl8h
eobK2tuePaQo7Wd0uJFSLTwuTu3a7gMJhOgoTYxpmwsDomIO8TLLJVDZ3RH2s/Ks
bclha9suh6ikMEIS1jDn9ZSuyUcZp0TD+GfQhSDl/odTNuIqN0WTi7x8jp7XbAaf
SRU7hj3shHdAGjwCv/fY2jWt73Q1xXnPpfJcwgnTIqZ8e7WCOLwGVIhNJLIhm+mR
VvCemSOIub2dQUqBtTtKpUoTggm5qov8jtCTvwpoGRt6a2PGwK2kmwsltiuqMSqi
mFlLsnZh7Q+kpVpRKh9tiyS31dH9uV90JDQZyoeCWaokkfH04SOe0WpRzbVIHv+R
Q9smSJjr/9hQae6LFEYpd8LloWjbazke8xqCqk+ShgTf2eQv/RZY2rr0RRhMYIvW
t/gNcvpXhtsPzKr+8AmXNA7/8laEcfclpyoCR0oO9w+toG0zagthmS9nE8PROcoN
xdyicdu5ort2DOXC//wlWknINUjzgHPz9iANgDs86sUAwoqPcAGuktl52ZSKd3Li
ClmOHyRH62q+WtWoJiTURNHgNIfVladgmcKb+Br9KvYLgj6dS7rLFt6Ch+UWpYpP
X49PQrQQfNAPyhSoPU4RUujlVM3WcIAC+jBmvA1zf1Y5Ct+cnP1Sz4kRZmM7yAYA
JC4xZ37demv+m+uUsd8hGSbRk5Gh7A3F6O6+nUrofmzveVzFaOV32bdxyARUrk7g
F1VpY6mImaQ94QeNgRdrr/V7Fz8DHFunoxxsIsQGwnijqu+hK8+2bbd+LUu8Fh9a
murMWD0bDVwtPTiikaT00BXF1s5QipBD+Fad4MR1KmUQrBLGd3AWal8u1WtWh/Ck
KC6C6iC8/suEFEkvE9i5RB+zewV1nOsbdOFeRpLrvYALBb+Lo8H8DuTc27PNrC0v
19NSvuW7djh1k8UZz3m6Hp3ABu8/NO+EGQqEKCbmS5iFuWkzxKMn44bmI3krZzMR
lPgVupagux8qS2gW267IIx3v3Vql4czIQ7KMXJVMoQmiK3vmXcDVCsnVHcTmEoj8
jAGG13jP1ZBVq3B1zYfLKUZFyVkiHhVH0pZO7KK7r+TI+OMTCqkmfnAzZ7u5FiRe
0r2WJCdx/y8Q3amDi+risLb/Y8GG1yCnS7FYlq1KEdm2DpF9x6YIHgIGh++A5EZ6
tqTeywevsOVqpgqYIu1/0iTFyevDNwf0AY1TI44bM6yRdk2GdKn170z4MaUOUAVN
av3MR2s/NwwglAHTbTO7+srKr31FhEJnE2aMKrIUrNac9/d1sBAwlfyIwoRVcNcr
j7lYEtnhMfM9SxVD49xrrQeXrxZLanGcwKlOAPYMsgnIfPsJe5yLyKqXaulfOQOK
wSqP96vwDepdyiFX3+itv/5kspBHNVX3RbO9q8CPxsVF5yddhmdhY4PR2Tv5LlXt
mUj0klrS1jF4cumBcj4GnQerLHNyGf0xQMF+vSGwdT+ogpDi78e5J3jpH/h1b567
JQ1EvonEeWDoSQ4SO4hDPEDBxlmKI54sz5S3Jk+ATi6Rx4VT0DoSU/ODmw7apRNG
pN0+iOPGD89KLAgSxhM4jcfxEADL51kSiq0H9ceTloYib3FoXQ7SiJPG8RUsWCmq
TDgYJUbYY4FpeBgsDVN/dVBc3cI4mwS9xiMPoESTiCJt/paMHHpJen0hJArkZuPg
nuD5KYf4F7qVzeIUXsU2+1de6J+adwkAPaBl63JsSqWD6/K5+rnbOqLuc0iWxjzr
KhgEGAhiMxdaR4Cohb2wCuHUoUmQL9ddkGWoEsrDCrcpxSxpUSCIXQ8isihS/fXK
70j+EVkKdznQidWZizbILnhBkTsunHwS2X/xRBxjfpQNPrxpqYs7IVFBPPLDCRiz
aELH1Q8ozaor8CXBNkBKQ/XNY1wuakPCgUGpV1rafVtcPDsmpbXHtmav+NlYsOOo
NP7QM+pmYMD3utyBRRUFUz3rwLzp6Y55Cw8WXS96h/C701Tsi5FE7m+5XohPlALD
+5GUFEGIFKlatZSKVRgUksYZSW1rC0QROZ5to3KOnpHmN+2l+T40ywkHjTxsFHEF
72knwEWEvpMSLoUSromV7HUfMpI50r01D95+nwUcVNBdI2R96XQL4uiJ2/36iJcY
jcequ78Zy4E6REsUJHBM6UoRCzKNYGDON/4frkg66tM+gj0TNQz0BLVUEvNe8EMR
KIuqGXUisQyCrSHPiyjeo8bVmfo5TbhNI7RhGRziSeEPRhBaJAQPEHJOTncRagsb
cE5cA4rAVDoIO9kVOQM3PjXNKW/YJumgklfGex37iOxMtjsXuRfq4Fiip2inzXzB
SxCKQ4wha1ihPrQozR3U2AELyHWr+bLbbcqbYdQCA+w86/ZEtIsTtKTB/ZeDcVNj
HzlWsakDGBbyoHwiwoWhKhawEZg1E9DSDwkk3i9zGzciBPHhfJefZj/OqJTPELnb
y/n0s/s4nbecWCEzBICa+veGGYYk0CK1wKxiH3KQA63y060jsVcC2RMalD9omG9M
QaPXSeoTtBuVFuG05KfUI+oDauKXdQ05Z4oqMrWepHN17mJPMndL6y/o/RO1II41
0sQmxSRjIVixJiZPRfXj23jJ7pKmd+Lzn3dHVd4nNthdZcq9uMxGH37qTs35Fn2t
Vj4qv3uQfxF8w2FDZIgKhTvYfU1g19PH5jOJrBtMulxn7lg3a6h7mq1MkG5tPzx8
49txkxiYKfS61wbaHVdjV36GvSNhEgVPAyaCp+eFQAh3E04/ntkAsYFc0kyDBHTe
W78LuNYSGlmwaBKrFQLz3+kTGAIu7omJzyTy82FnOtWIoSmMObE7FPcXm6u4r23z
4DxQrDtJG5G4sCOKmzT5hutHhrsxdSiPpFtNYti3H5VkN6j+w92220jrWpNJGhOl
CV9EnJUSkFmhQucoLcQpKckI7D3pemA4jegWAJOoDur0E6ovoCaIcxyTIIjaPl1s
ExPpBV70UeXEWtIAsbtERrRWfQJcwBZxN9jK0oxvrrwUXhawVUB0bYtVicryjY6E
SiodJ+Lda/InkBiJZ6Eo7tSBg7Yvh2dDn4kYhPQxYEvoFiSA0vwwG7oE+5sr6xtK
eR+DZLRjNs7gjSjVKVtFi6qyCdbhO7pfcH0GseFJaT1YXgXedfLOxko4xTxp1ElU
762pM2NM21X5dspp+yg1vUOZyHIfxT3JUsMjuQbIS13kE2SutZeJnO6X+/Ij2xIc
MQUL+9MAtSdrwj/hJjIZzfUAGmKOavxHLvO6K4f5pMauqJ4coWQ664dYVIZVK6tT
sERI8llo+KqowR7mXOG5zVZo2KTIm9JpLv3/nP1a6ZPJa4wN/7J0H3ZB8TaMirgh
VvxCqomtV42+qaUBtZZt/Fs3OidY9PTJ4K1JGJv0FW7hdIynHhGl2na9K/rIHT9C
IAVVQdfwZrrh00QX23VX1/sULe0WZd9micu0TCjIu/kn1wdUCcpYdu9yA1WiJfYR
d4Q7nBRySK8AigtDDQX5LgmbE2D5cbEE12ygG6l8oMJnHh49aXlyUZxSxJFeL3wJ
j9sLZ5ZyI5eXo+WkDKP/u6yzsylOUkWSZkrac6XP3CBcSu0C3glkxZf9DkBN2mu+
mNkbCC3xcdNEvHcft+XokEmQmPLBpjlPofDUJZBNtvztBloCSp27oCvvY0F7/OuH
/Qz4DecXvlveh7ewmtR28aItQwqnk21L44qg5l+ILvWPaM9XSNLhrN2MQ1oXdYan
C6wR6KfrhF1s+7o5+xk744Kl5DQVbMiEwC5C63b6igfKuvIPLKiE0dqPDa+GJrm/
agK0+x8gwaVSCSYg0sHRopDTk3a/bwj3y+nhlaj5x2V+6uHrVpavdWaESmHjkV/W
bZyb2U1lf7m3CZ7aZGmWbHwH3Zu2ISVtMIlG0Fyyivgl034EV2toVNdro38gMBXo
ScFIWbbwySl3vENKJY6FF+2fECDMsxxFVh5+zEVFkqCj9hMPIfcAHiqyMnRkY/Ae
FPYQY61ztsy5FVonUbdzfPfAdkRnPRnpqkSusq/Lqaj6VWv0LYGBT/OU6VmdZLdh
i4yvOgvyr1fT5PiZgPLVBlkKXPr1VupYAdA5wE664uwZ9LPBgm49ZtgEerFxoaN0
VOWEWDkIylaslS2zRK9XBd4Gf6WUMhGjdcQ0/h1s0LkQyKofdBSehLCUP5KmGQf+
/cvz2z4Koxb3LZcIv9/7Sgm1RAOxJBg2Njs7O7GYZIRn6/pZe34mVRbj5bbwcNRp
kVx9C9kAKDygkPIO0LblEEe7qq/7cJ5K13AT3qdgfdBOEdOPSquQrz4VaXmTD3r0
qoDx3y+ZZY/jITlYwDRBC2iT8hkdSgvVZNSeHfwW8g9k7Poen4P4Xvr4X9RycZoC
scZsC2iDVrj4mIf1aYQ0ES8ErTJSta+MSdGBLHwfFIy9HQh7tFS2KLDSRxkSa+kF
EKiOngl4vQYBHu/neEO5uD3yy9+fZRbY5qgj9qOcdfoW7hQ+6zZBhPL75f7nliY8
f66TNPQ1V+vu9yl8irs3ryyXLDcNob/nx/xKkAzgWbSRK4oPMeE20fJQ5PkH7M3t
cqmCUfUrxnIs/4rExKFKOUBO5cd19bgbe1i5PwiJDa3uRCD1yQH2R/hkTm8IGJXo
nJmfSDXGLaJ8hzhaANwqffQ2P0bQIOIjQFx3EZUVcf7BLav3jHqyjmcMRihLvFJ6
K6w5ety1QMtL4AeeQ7fyFfacknfO+KqOr/ChnYTOlaqXtIwnVFSbKnQYoz3mWAc8
XwHRwczP+Fwa1WsdDmhzC+xRLyIqY3v7GEQ8BtLl4i49tm6ef2a3WojkL/JTIi9I
oEwE7G2SrdDsfbGAkiMwOnwLw5cqmGdP+p4EJXCrcKj5mx/QjBw+ixsXGTEr3oMK
KWX90TQ18tVs7xv33SkiAeHeRhP7gHijtwN3WCJaWEoeuhbVSZZBCjf9fhQCuYTn
BNAfuM4VwOaIAlAGlhQ9TrksJjo0k0YNaK9ofHh0Ll0u78ysHFcKxSf1Qk5gwOSZ
kH/BP6lFeKdupydMc7PCS7Nveui1gYA+yvdw91SdYe+ORgF0QEOijic/beR31TaY
D6eH3Z8eCsF5CfkCJPNecnW4rfL5g01Br4Yj3EsBiEAfwbUjoBXfgIgdwbX7Ug+9
DTkR3tXj4u3Sn2GKcQl3Gz6MOilFdx8We0CehXIMoVENNMGeGEgAlIZK5dcaxNqR
X5OId59IfkMK/DiaBjo1OwinfCHb0iXt1Uf+TBDFlnUHIaEAkebH6cdNo151vxQ3
+rnPQ0y0D4r6CVQHM0zJb97VSmZM7GsGjU8VbPJN1b7oI3lFuq7YsagPggiHNH9z
9IW+1vPeoJMIG4qHilfJpWilfSkmlI2ULRAqr5yk17Y16FESn4qUBazEnSdN9Vg1
zDtTm8EQyPOoZ2HzbtFvKqkxAVfooLjXVWC85oo9czaH11uBBmtr4Y0QWjvxPS+g
/3m+pPfM06pysuQYaPlIy0vxm8tf/uTr1D5291ghMdLD0SbwOBJcHrfnGgjPo7u8
wac0Rwub3zLuDQONWwHb00boD56Im8xWXzhmokMCmNgumP5r8/1LKajWLT9R1Fqk
4OX2YYf29eq3MN7L1ByZg8ipjZ/552GJMbI+vP8VrhnqNKKk/Xt7qKhyEgRGv6Gu
q1wn3aMLZ3J/rqaEEXelQXY3VseaAqujfPNwkJF7jqPWfML2K5rQhp+tAWx21MrS
4jl92XabbgHVJrU/NSwHHDGbsOMCud+z7mIvVuC9tDCkVly5/wE50E2yWLnS9zT0
YnsALxVmSgkCKWqXjXdD74V1aTp1IeiI6bKdMxm74NIKfbVDTXHSVQE3pQ9dPHMe
ZQKuWV0cYXoYgu4kssCprkAegQbSww4FcNC50FruV6vct151AYN8F/UKedNNdQUX
2fBI6v64mBk4bIfXLZjk0eJs+m2qW/vAluVvYhihkv6EiOW0RUADP8L4Kefuq6a5
pXceNvG6Kfx0Hig/09ym59TbuhqPtSdPVM2R5PTWmmgZ9BPXG8cx0pk3UTsVEk/i
sPZP0ovpNKh1qCiFeL3ifgyKRUpbM4/5dC21REP9YNV/SQ4DVH8ksM/2LHe08jKK
/aJN9OdErywcCDKbrWxvkXhljQaOgWcfLzPDPRM2vGDwz45n0hyRO9RTc158VFdz
E2OC/yee7LNh68HIgWRjvct3ioqqXKZcJXnmfXTwEu/fUSswFmQpaEq+6zM3csgQ
QMNTqFAGn8MGgDX6boU++9T2VA/ZIpYZRVbGPrd4E6zV6H9XmKKCnXELM7Mn4J88
x7aC+EYQXo1wQl+zKnuyZVcWcjK8P4GdgrV17/Ua26aj5UGZN4gdb85Inj0tfelq
fBvnuhW2UVdY/qyg6LoxsDi6DY11roUtb3cS173expCXKt4P41CO/9B1CpNwI/E2
C/mezTLRgM+T0UuE9O+jQn6v9EcASLxozwlZxjbLVs9/fFwdKnRxUvtv5WjlPsD4
vpHGzs1PwlIwlRVzAK06J07xbYBzr9o0BYXKnyOmlsnFcbFZMpET7zpwgll+qhFt
jvMEGzIO2Kafuz5AmsgXs8l/g+mhqh/7W46lFdBzg08KYHgsxE8SdmTHsxf5dR24
zMNwo1mVup2hQj5N42G6LChM2r3jLRCJjKEfE05QMvsXvbNWb6USwqLaUbR2fJWg
y+E64zBJ3j3jYNJPZl9cBwYBso8HrPZJWfTeC8E/nJK2Ic3UXOr4kAd48XdKpKhr
oHMTLJS5WRbTnQIjf/K5sWpwEhqsYGvr0h7bxNoMjuAOaAUOHa3kbrUjTPSRIn15
sWoZ7sbuVB3erXep+Jyf0b5Os25qG5u9zuNr+ZPASstyiPUBmiKywnubjyfwFm07
YWYbiapAyCLzF7P7aCpTtXok7IbFlDMFUx0NkH5ykUt2u/YyqRSSDCjJb8ieObdf
Xf/HX3mDQ2m91bTrSiRdvLz3uw2aeCN/+CLKGr79h0MGmM2fjkOMnfA1jEjOgQ+F
wNXzB/dkeXyITGmWFuO97RqMpYJbyWLlkyMW12cR9HYKaSLl0fUoz7VPHfxNCIea
6Tboq2EUpPTC9zuLbwnsa8p0/CO6HPXtJVPi6LykL9r8jBmDg1UYthuk8uzVHIdn
zsgfBTfcNKtcpR8MdKZSSUMzp6HEthlWDMcinqnz7oANlVLQAPWHwNLrysnC+P6P
TlQ8J1JBT7KZTwoWrdnTrBvM+7UXOsiW/M2l2iHLTK/u5hYuvmyFykMvcDxwP+1b
tLeBN3YMqD+lAE4/EnhrbMFS8fGmEWFCCCXvDxppySgAZk5l/WxvgZc8P6DF3r+9
f2wf917sce4GtywYraRyjx9PIaJuN53V2vTVcrIpdec/WrLeB91mZtGyDo34qf4T
kF/RMjPM89APAdOCjRNgo8gvPXWeNG1BALjTJIGsqpkIfd79/mZcsJL+pRJhCChE
/QVQiM76vI/s4FIpEiz3cGBAs0XPvF0PYaqwShAFQ82nED0wt2EpXKJ6XNyG+0A4
fdpjoHA8j+JdslHIfyk3VgFWRoF0JqyqDvj9pIae10nKqcifRQPIPiW/kVDFiER1
gG9NO9bB0JV4LPzhsTcGGQYI/jki/0ZjSclKEHDLBaGFC2kOzgeNbksQzgSkHH+R
tPFGYy2Vom0zr4WEFobyYBXFgcZZaSVtHSlI1mDDgn9hFHyBWP3CHzMYA+8nj/Xz
+RuN+M9CX1OqTYabXuzknMneGw+jEcV4opVCzH8vN5T9zelEbbYxYGvm51/LiIyn
8cD4T6gG84BrM2iyzKS1G636dWGxhxWOpWHcThMp9kJ09CkU7AAt20Q40FC7Wdjb
IkuhU7M2QogmR2aK2a/11dUTYVCrCSl7/5sHUWoWW9V9GzWDgW8Ki4My9KGwwAUA
gQ1Sp4Q0sMTumpwpHxgzBM+HDEK1nANacm2ZyNPPIdCHCu7nLKk2JCsUm7NP8UOK
puH7263mc6fLabs3s9gyeuEPr976bbSt6DaGh9iyuTp75KxsdBkerHr3ZEcg4m/K
9ebcLXqb+tM0dWqEJqgD8Rf+NgOq5lgg368PF8oCGIvtlB0USEwENftrXRma+hwZ
kssGal3LZVDzvzwwPy9iLVVqJKP1FhLYNGrhCPn4H0zkgfXIRTG8pVJRi8Vdciym
sv/CYGauUK/nYEUX+PDI0A8QMb88le4hurq6lr4uTXWGwgXx5TGrFJOnQkFNUcmU
LZTfDbqPojt8ztqN7XwhHPQxf3afsTsusdXULp8nXgyCl8Orj3C3UHXRJGA9mmtz
dBnbTExHOD6EigvnuXt3aoE9MCjKDInX9vNsj/hDSZ9L4o9MB0bo0El/tCTkQrOJ
B/2Iv5FWoQxt/VH6LIcgNP1buERAGsIntt2OEN03PgqFcXhRaomjw8pYDPMVasr4
lwvwzuvQOePdL0FB+sjb6CKdthgOj5BNZ8ERh1YH7Pd7hRpeXq0A3CFSd4ZbqiEA
RAZJ99z4G4s5zGXZ8BLqpADRuo/mIeFGg72qZvtYGOuSZK7wihKDAsblfdK6krpr
BxsuByV6wexvq8OoqD+kmn+CWsEileGpBi23xkUJSNfafzXfsd/o9TBP3Ik8nnOF
H9tpGosaK0OCDmieF0gYxWji53YCWRjIvNnceY6FLOu2xMkAxIdNJeB62tErMmbl
e0xEWrvarkCdKPNFO3kDHG2W/XUyEYnN7iV14INLjitjpEmoxrQzMVkFfGOGVFWK
3Z5USnx7oRIEmYrexdZd0MMg+aY88910v63P1JMxBu/mbov46CXEg5Ya87fo63JX
XpZ4J0xivQrytLy7T3T0t4mkJa6/0uaM4ibQWjzYikwbq5SEzCnlaCEeABZmIV11
EyJc8KOZeiewxZjMYF0ld84mrRDdJHgeyaBF885wkLEtRTykSB0yhLQGsiJyUhLY
jUNY+dIdLjKsgHVja0U88qsOmjNVXbSgsLGTv6LBJlyI/sjDhrDr5mGu/pe8Okxj
e4+98WmxqgD0KdT1eI7yZ3AMQocYEryvu2PioqF1MLeQjf9G6UgjkMefuR+uSNRz
ZWWOMP3aiilSGK8pUTB7X/fLemlKbw6p+IP6pIwd3Aqg2U0DDS1tMIoASLtASCY+
`pragma protect end_protected
