// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:15 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Yd83eqyQXoyiQiTWVal/RzdkX3iPP7/JldaNqMBfPnOPnJfq1vscrAV6rQ9mvUGy
A/McprjpWscYOJEgXZu4DcPrPZNpzfcaCzfRbk0rAO+1zWqFOdtH/YmOZTStlTAr
OG8d8z5GSD4e3Ev/SsoFSTqwizSoyxr0IF2qhgO5zds=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28048)
CZSQd1bYCmQqjIllPmuv94KmGI48tx/7uJvz57k20WKxOmAQPn2qCPJD0aVifkCU
rrIRyb1NMqrKXpb7qN5TeUy75pUWcGk3UzkAmRYXPQKnVJuilv60GTwk0cWioCwV
hLi+3YPVkRc2mjgelSP06NRxcJG5hNWiVZj6sO/kwaVThFAhTGBcHGMJoRe7gRcV
0u6SFoxpuBDXmNAA2nXz3peEmUc0y67YQ34DoE/BQVgmnhPtE9X1h+wqY4z/WTrq
SL4LaG1OAC68J+EIS2ffUbVz6mTjeXeVJfrjMhCAOSu/8b741cwQBKRt3eta7P/P
5Xqtu3pT/yCR1DT2bwVfycwghmplN9DhiZi/rjEosDtleM88PgfBMK4FUYIk+86r
l4cwQnCNgMmtc3OyIBmpf6XlxPwXZomzIqtvtNL0/aiSQrPyAOhPkQh9FibeUkmO
eDA7uPEd9sMgbtVZh4xedU0E8sZ5cbCuxWBqZa8wHsFKFEKva4hQOgx+3jJ0dQJi
viNwZ2GITI8N9vQ+ZOEt77PvG+QDdGK9FvV9e41cbwrDLseoklWXfuon28NTPEUL
7sCb8KueVBWHCS9HgYyq+YJySWMqSsZ9OLcz6lTE18W23UhPzD7HAvkOTAUweJxp
d0zbG2Ra5CFa62FnPM9pKHv/6tfsWeZzHzM/VLg1Ygkk8xV9Xj+12qXWFm095sCK
sUZtYh2UxWdF5nGjxwW4/3lnSkywD+QQ7uPlr3tw2WdN1usEGkcQnu+ftjWXiZgb
y9IRtOpBeJ7fblzO7nQHZejf0cjZUnkCbM3y+PgsW6ttaDdnrr4tx4js9JGsA1id
Jv3rVwqLkeezIeneZpLtfq+AEmm8/5EK6M4k+1xo1IJTN93lym7fLZp+4G3dMaPJ
rhqwZudSMhz2JvznAVHhntyvYmf2k9Am6Vjkn+ikEykSxU3Yh1fET5TspxxHy0E3
fb/o2ufPPV5Ho/gai82ZMLZqcvpSt03NdTanzWVrJLWitQRSbg+q9sdiBaBMBuv7
KC1v/vUCwd8tzgEymI/DJZRlyTevWmkWW7UdBY1bEhkjnvhOp0RAQLBwvI+A0se2
slpr1BowVVgs4j+w6WLe0ziiQDk0nsxjfGkV/FQCW13LI5yPkSzJNmXl3J3AJuW2
UZF1z2YGosRJAjJtflFeibfYdXG7FcXjXQbpGqwlxbczggJBMKmZh3Dp+SeVw10J
yPkaZpPaZHe9BEBnmPUpnp261sVlmr4/UH8IjI9tgNvWOjzRkXxUbUbjDYiOs0Dh
ANSAtWKttNBKx2iEiLUYC6KLQWx1dUhAAaQ8cHH+gBduBHLKvyL/t5lEEKvwKVdp
Ij0PsCI59qpbtPgBC6dFNOOkzpVjK5WTCueexKFw9O5L/X+KjawDq/Q6TxEkdW15
22D0/TjUAtrdthPt0EKmBuCoUSJxTIM49ldVYCNG7ipWxatTter7ypLV1XxgRSUH
MjAANATo4SM+aOB7/a2PLXGfto9R2vEPFiexRsU2F0+bolpks5EbENevg06iGHOS
I1Ix/EJNsRHLSziIIYj4UymFUfYmvcA4aC+eTLWU99+2xa30jqq4WDHcgb1/f7/c
lv6r/5TWC7IN66HZ1uyqaKR/1/VcmYRhajXdwP8Qr9Xxz2+rcaSTx9F+7KKhfkr5
MBHGhKDjI99tM9SWCHplfgbl9tMtJuqGylJmxC+nxgqw1VbngOWGU7VJg1C6HMtC
r4AelU4qh0zTCL+tqLmTRcUC/dgFYHbpU8bEeKFlCjnpSBGcxo/ELc72ax32wiZC
FWPgN9QhxfrDZdGJ0n9MxakEWMo527ZGAtDU9lzgHTq7t++eZeOZOtfZ1zMTDiDA
u88UkQXpX8PwzPGCB21lDoP/SXOJLR6et/uWWcW0k2BdDysxVGTfyPAIsDkgLfA+
+kjZ7aPtdDORpcNX7UDPLOAv1LrzjeEV2ffEbbguHP2mQ/SOEA1QtpIYnJqWu05r
O82YXN9OyO//BmQYm5/3WKZqIwv8xP9djieygfLUjZU0rXA0IQ44b5+3/SFAFvIr
uyEx/6/j4fxnYOQY7FY7AG9cwTYyN747i9dPP796X50wseGc9spILsq172Lt+PXN
X/XEOovnCy7WpXbpF7Ob48k0ceijaKNPkb379W911jUnWBZkHo5w+5Y09N1ul2bs
RsVTU9vWh5fmrSQjM3fpjkGr3XMNMVFPbUA9aLl5vAOj9IgmJO+UeUtoApQq3jh+
Eau4p/PXEPZ+GdAlp0vyHzQTz1hbPqkPvBwR1chh2NUqFbf+8Xf+gdD7i5LrNQw0
FBghtdqIMQbFnhs3oww3OnIzs00B9dtUzWvJCF9+QgGCoBUj+OGM05os0Kw/0+rd
6o4vYGJHv81roKsTmEgmecDvd0b0/EuyQwkMzGVIqQRJRDp61K0H2bWEtRj274Yq
uCNn8LwkknWOZGUwA05t51EXDBi3IHXEmFV2NXDPERHPxyZ6i3KnZB4+72Aa7X1Z
p00Ajrs6F+r8CLYTHZg8gSBl/5oEcuAOpnY9oyYRXwGCCZkZ29y/eASz5ZCU2wHl
HZSEaCiI8l9kKmLT23rYp/mbrsufOPFLm7GTBGCzsM1P4nPwp8t14eXVZFxyQAJd
S5zwxtn+Yt1PUpo2lgDk3dNNjo0QzVz+daH0Y321FVH7evR6csDnNKEdlRARCq3h
epkUapsBRhSqB7kgnhMRV7tD40St0RcJw9ZAuQtXE+RCgye5tpnwKPu6TNPIF1kC
GOR0ab2ZWGHHJ7IAHixI82b4TL8+w/UyEF4fhlUgEHUI+RAe9QSnmDb4qqfkQ2th
nBCcGZ8xwTJR5O0khGTJzq92I7fSWK3OTC3kjcqIxRK2UHhp6gIE+dieDeVw9ImF
/iRsDPunrhF7a+ZDL2GnSvytc6Kel7IZH9qeM099lqMidrGB7l6xX7dPjt0gmdwJ
DM0jEZdyrzBnf/g/gJqpiZoibYLtel8j1oxHiGuC6Xsoci0Jwvix68IT9N5hyozn
OF91Qck7WPvPECiW/AS3sR/U42cvF2QbuR7hgZQMf7dF53hJCmlWzlAy5S53RewH
GgeLBLpDgg7LBI7Juy0nUGr665toZarK48dqMLMcYbzH2ylet+SuLMsHlaBgcZvW
HvcW3hTvztMa5KqYp6roWhRtW5TTzyEDbD62C1cfXPjZpv+fFzUm1c9CufD0cy75
V/czTDftHZ+cVScfCP7N/nzHatfrNA5T7uMSLNJRTW79q824QK247MYqOiciPt/a
Z0i6A8EwZYKxfjVOx7IQdBxXv2at1T7hmYOBfyPVhBwpsdpxIFrpzQ9NapNt27a9
wowla9STawYPONeSxomy8wppfY4Xa2G+aYq/8CBpym5rC+vycIYm+sPW7f8JPavS
NK+XjMWaRS+Wopr5jRYW2n/MVmXM5TAnnUhO+UpzcHcLUOdKdv3epRAxoovsnN1p
Y7aYMsTLj5Y6RtchbHoJLXY2vL+z7I/4RkfKy5bdzG1oQ6WKGmWRrDorns4qNH8P
b/d1/4VI59Q3mkNH19aShIgftMRIQFVZ+ucPq04CplYqlRrY6pg2q4cjrjNOdVmP
LRC5cYUvJ9P/prlaPa7jYfRuRH3tdtgqXx2JH/q2M+8H8wvsNUprBxdWSpV6lW+i
3p5oFJ9uf2/KVEnxL/CVEl3mgNJkV3BJy7ug6Ksc+UdH8dpElPpYUVHqiAwVydfE
a9fwTPXc0BNsFZU0uEfBMvmJwyO+AZ3DYwereUDrCscWKu7Ym45/CCz3+4Omhfjf
fgdphFJYGWy0I+NPYLKdkcaeJF9z9Q5s2ZZJlAxV2KTfoXW+3LONv+R0HAryfw7L
+xck6agKThz/QBWvaR8kRZ4buJpqqMEgz4YH8nPDU/fkqNB9zQJHLQnCop7KDjA3
vKOcxlVPDuqXC3BuuYrOAsqrPHyQ/mYOK7pIzVuX/cGoxBcncUvRweP9S9viqpRs
gDup7RRmziNBVibKrEhTvv+qqBzwAHcobcybK04l/dGijVVkdNMZildzT05WNt8f
wJkSYZTWjrlyPHMmsmYPtN2sRoI8Pyj6ryxingcwzoE4udowCPC7OVdxM+kdGfZq
NInv83PL5gZ9wBF0ebppsFFxLP7lx33xNF16TmgG7/KrLtg0c4PAze/kmb2cKS1i
OcPtccXojYF3PoN/xzqmAe0F2KsjYaNNBdYV6Gge9FX4kw4+yyRyaZAD3qMDdAwU
GvTQVVddRX4Ye6gySaxuXsnorwxeGtg2o+rAHJJm398hcbcksjVp20r+TMcgsd/i
cFGVoQ5hsHtVErS0mrQIPfA1ympo0dVbgy2n3qiSOWR46B1Fw0R0BVoJzrgN2a39
2VLTtDvb481dghV3gXHYhmdUeqgG3bFQ2xHf91K8t5HndwEYb1BkuzPiEi32jad4
YRdnonavlGuHsGveNXu3QX8UpA7iKPaj9dbsbMIq+tIAiTp6PqgcEzbGme29uvva
cysWRmx+do7pUOa8pAEcHfyDHTBjpOVGuwh9sBT+aweWGbrt/fYNDQ34kAH+xsuO
BgIdOHSea7mJNjPgEzqVkV3o24oiGyR24OmjzNbq9uneW7jCfzVe4lPkwzkR9wln
EU7Ck4vBilx8OPdpdXpwYg4a5jnkE18DWiyJSjcWx65nfcGnYPr7ibuoDPqe6KxX
UiCwPnHZ7pOid+xVOFr1nSbuPwo//cgOVTnPfUjSsCtqa11k3Zst1MyFhWn65ZeW
SVYtxqBVsyYadtBWIg4GfcX0y/7SYjgyf0Ku2TFCjA24vDU/UQdnvhi8e0BWkHc8
Vhgq/bQaJ8c6z2KWRFKM/lbK/tmNWOboXsdmTvmU6kAyxqa0iwI7rBV7jTjs2Cwv
7mAGVmGWiB9pYlf05KRD6s691k6Pout9rK1qo31ITNHshExvKWHnCCEgOpDrfVFM
yog0xJANoERCep2ffLoj3D31g4g+HVAN+a9tAmNHbF49kNE1L4eLQEDOFNp63yGe
vgjBg8YrfYXHZyqrG6IUA9O9Q1/AURzhTPhcXMCe5m3yWJ1QERLTjLGSmDrW7nMp
zy/4MgsTb1W2wMuMSM2KnidMewEbQ6xHNH6pVEpyx3zR0b4//CbnwAF4b8w2mnNO
/pSLOUArUwhSn6lvJtF3HSYs1x2X5ev0wmbwcDTQ+dfzAg4eTQpdbFLouv30IHcS
oXfIuipmIHUltDTCTF4YrULW0GeDFrAxXu3BUjxBWFQ/NErfux4THv/REvg7cw0R
a3BKOUMNdHX3YKSrSrs/jDRpcrd89QRKVeRSyEI4XX1/DQ0muRj2P4wAlj/1w20p
y17WtGMeqBeaEl3QGyPQkiS3fmir/tkJVySiH4PIXGDcPrrP2bwK/qMXfTG9Q1Wf
I3QMy2wgdI/1E0J1YoVefhFVg93Y2qEyh38mksG7TEPj6SqxJkLWb3iVXQ+bh63g
K655IRLXVyDPT0+awGtf7aVjmRxlIQQ5TutaQEATfAvRWMxXkRWWJDvfJofQrkNq
3G8MGIIYNNQlH0JWLYEkzDySNNPzsVddbsYoZ48y45T31Qz46jbTAie4NYnT1W3C
ZsDLLap1qCdEgoCn/jSsTHyeZQFkX26iIYirYmzAi1LsBlv46mx9fGkWMd/qstUb
gjMbzCqaX9NPyzicCcDfwleI0vqHOv/EYKXWbfLlM+krZbdjvZAVn9+oaWfaAvgE
fPMvrpuY2xaD/C0KWOhFZBWW0Yz45UdA8aFZFo0xS+LXm4KIOn9qT8yIuBkp0YGe
aeP9kLXf0BTI4rsiy1FdkAw2O1bnsiWVrZ2ODND/RlwV7rMAqGE44nWMsZC6zZHm
PR/sn2bx6wby1wwQWhQ5y4fE8JWvxyb4By2nxS0wUOEvQTH7EdDQpSJOj9WkXcuA
4PVBb1B9zMNLdiJjzjLfVxl0rdh1JgR2j2YHjzd48gahysdZ+ew+goxEP6ZzdV4V
aeJWLR/B/UaaotoRLHDnXC2z99wjGpIBLwaKTFLG0txFjvw03dJrvFii7HkYkozE
WaQWO6UK8fqvLVCVotaIcC+ksNMUeencXjHNm0psgSELyX+t4FS7X+0YJ7/xj/Nu
rhrNzn/POSps+AqfMG+s0dYaaQll9bVzjmwUrMx0LownHxyV0VW+nQuBdw2LVUQQ
xFE9mKlQZND98Eh/gDceuaD5u7qCnNHgzy6yu0ZvllNbSmjjfRvdhi9TbKtW+B6L
efWpyiwkSfMmNWtlx+WJQcaoJij1nFqlLa67ZzhFBhfjkuxbmNJHw/PTIhD1Bbkh
xBvpkrbb3daf3c7Aaz6Xv19lrsZ3mrae8SOSq0tzdwP1HYkXcgEWAeiC4QnFViK9
97kmtTTvg3UBnS+6wXite3PSC/Kt7dsyR+zMZ4Cq9j5qEQuii7WJpm2yTrlYZUrU
UYVIkprcArx7xYpMZ7bbyasTVxOZ8BkfMCb3mQTHOww0vnDXKCF8ztDmvVDh0uEq
HftSpdcwFqdHAawhPfo4VqZRP7DR9jZO8zJHNciL0KMIWvWQ7h8+2GVIQCXcnggJ
f49jXExpmTcI3dfNdYWYGh1Om2lzP9kRqTsdbl5zoT00mcJThrgRn5qcI6P4BX9w
V1+XVP0WGWQqMi0XlLmWyeIBREV/nJLp0e+fkexcIdvujK2g1qiaRA6QfZw2CyHY
7mctJb3bUfLZpJ0jolBu7hWCD859i1VXEfxaE7o7euWUmU04m3HwF2QtJGsS0uXx
3mU8ZyjJiVd7vvPaMnKeijCNpJ6xKFpVTidm+bn0uLO9uOZ1cSBN1VQI7r7jCZTW
i0eybZyymZwlijO8/Tmi9zKvuMCHaRZRaFssR/sDuHAnZ6DQXGlLLPM9YJtwUalr
spgjLI8R8jcZETl1ufOloAU8dlMvI0+ynob0YfALhiWYMBijXzl/RxF/IM9a0l//
kJKdxhGkBz3LtuP+hV4MsPQhShAuNVisZO99TMGA8d82b/0QhUlnaQEgUE9qm1gr
vcHIJVdPGKNrJF6KzJnTdeJebryxZ8x0bmm8s0pon5/1IkzJLPTeezv8HyEZlgTq
ACqauxmyDpeJQvuqjq8X13euq7yCEh5eNdYhowZ2SQ8OKZUD7Vgd1XQvM4ytgkKd
KKSETd9pqLlvC/p7O1RPuXlzUSlIJGJsfdYiHw+ERoH34DABSFF10jctze/M5VXh
qUvwqfQs2j3feqwfRwOTP6wRPPqTe5y9p0ykLpUXNO9JuFbSB+xes3i/ZaklsB9B
W0dcR3FsatHEuxQyQwO4JGlsCDK19JwAYBuB/tz+98MRi/u0Sf9MQw4RJpLxQcYo
xWHru2L/7b0md4y1QUu4W/SmqU3F288ePGLi2NSPPXus52wUK0Jr3rR3iNB17UR1
2djTeqN+bJ2SKM4CJi0fPUnWF7bFAIDcBzlSmmclnEk6VcZkVAK4VbfxcEH9M1ix
e5r4ZQjCvNDtVTG4jKxg2FZBAyCoKVS+xRouw7lh+Qc9AHhZ6FcQbE1nA95SuYf/
+g54OFQ1Mo7IDaFAWr1ZVH+U3VEeeAbRzWeWMSn3fw/VtVheRoXg56X6kKZYXuA5
FpXscNWOX/dKXEXzHs88EUL/5uIjDM7JtIVCCqeowSvWG3RaZHlVTJuu6jbhPeTV
W42nVhnnK92tj31Mm69NYZCLWcvrLihc4W1FfjKebcttrynJ1fTGVkLjM5J0UFwI
AiaTqJxi4x4t2ykUvCgLrm/b+LicvN2+ke89eA/KSESwxfcBjYgeioeCaox32qTB
ESPI0aGEFRhaM6H0Fmm5bxdsqHvQWd4rBAdcxe7QILa2lhQ9IZO9H4+WSem5WxJM
+Ozyht//ym56yR77jQ3gjdXwcw4LdDppETCRMn3Cl8pRoxD2ucXH9ixEbXKuze8B
NcNIvQ532DrcWuNwxcpord60tHupNTFjXmZ0+qXWf/t2qYi0u8G17TLrBloyiATw
xg1A2CZB766dGarRLqPgaqbOijtwrelpwnQ+KeGPMw3OLj3akfqU53cXN0siMEo5
GI83Jieu2z8iJn6TQeL4tGBeRsBp+iBy3XZG99zdrjxirGkmrFZenCT56PBMngpS
hLTOoH2TvSB/oPW5RSAXd1eN83DAFVx2Yvl3gP/hUxEPc5XimoIYcIc3GIEsfAT8
mefCo7glsA+F327pQfmqnkx9Bt6x63OBLhzaoIn81LKdyXlw3QCOzKT5jlCfQMXZ
PiqDnUdhSTOsmakJF/SKIROX//bacRkMHvS1Z3caCbCZHGabwzY6Xzo4sKzbnsOF
kYpYoBoCEyZw0j42p+Ax53ipJM2mFPN3fVgCgs2+p35NQyrEl9jxgIZdZmq4GQp4
ZFBMe3SzrpRKIKtlYI2qdEBKOoiL9hbsWJuwayjs6Khh0udzUV5VKs4wYu3Cdjsu
HY0gEh2V00CMEfg2RN/FCs1HouLBPLwI2KLgPWAw+/2uJnUx4VCsWvVUrmGDkvz2
4mqhskGLDqIy/O7qP6N0mcKRFMjaRrxkz9SlaAQ7xju89DfTwvls0CHlb1GWLhtN
BF3Zdts+3lg/AnrCm8zYh4kYxCtY488Nt31qMcI2atbwvYuLVQik2V7n23nsKuEX
iOjvfbkz5ZClG8eQNScnskzTuL/p1HdVUZ9+OiK4W684Aa84yZJMmZTjMaE5SjYh
EefCPaNw3Zoc67rGFAI5FjAroOEa5F86/SekoVgpVjOVIzF5bmxIThrjcRV0kxXZ
lntijbr8pwluf/7EUHTvXj12TYBiUrJ9WLsX143sEMDcX94UuXj/oLquw7xr8X8b
XSwd4rRTtBab7hf0asK05GfNI5d7bpc/H4v7tUeBrtpNRKzjwAGNeR8yZWZkM9sy
s6I9AhRUC5k7lH5rHW8bDATFMGuEBdS0ERIrMcePhZr+5qvq7N8SgGopIyyLqQaY
m49/1hNIhIPmpuiGd6lhMjUQxVekWfd3esg8qIj4XdTq9wT7qYg7eIlcljwof/BP
SKu3PDykSHIxsbVAED0Z8ANzQTHDMOSNarYp8DK2tNzlu3zC/vK4HWiS4jEBvkYn
vlbhtX0eKJakFKPNd92ZjXR7VnfKIXhkCgmBfxFqFHA2H5LbSyxPjJ+ttSmRAnmu
+lyP5mhT9YQpjua98fC6bCiFPh3oxfaJuOTNRZpPE2hVKp24FajTuwgXLU7n8U/m
Esv3shaKF0aGHh7h/b5PTim6YVlviFAyd/EIjrvTzUgS0F/7yixdpaM+808cKLcV
Cwxett6RKXSoYa0cnpCppS/NN5EDhH6Fmvx+ElIE/jpkBksF7X8Pn7GcE41ehpcU
rOjh9X/YnzPcT6fWYbGLXhpSY0jvKgwVe1WxDqk1XEMLzY1IPZso09RmQChppjED
vYxJRNVxzpzW6UUKXCAI878cR5zgWgGah/4pFI9D3SDKcIO1qxejKDNy6Lm2UfQY
f+cAa9tMI2zh87/mSYwg7WcdAvWGmpkXK/VUuf2MtagfF9JKPttYfxtwEDijv9VS
V1QSi3ZMRuGwoc18aUVSa+eMlG2g/6PLly3Id4Iq37wMd3IgIuxkotm/oc3M3y8V
MNAaH1Fx0d2qfksvLAThuT8CA/KRvqiM6PXN64PrhSbTQcY7bDWPhU278AblC4RI
LgA+jHExUxisWyTp51W6tlWDz7DWBemmfARnJbSd/YJLHqdVepkMCHRvioAzQ4HX
fKQJ/nVG1Enq0E6X55KxDrSdojqvP394VgUnMoq4NyA1t8EnDgVkdsLiy2A+r1cJ
k6tQSE4S8x6xiXITmUFlIAtw49UEWI4BNXj2A4YIyU8jKmIx4SoGL2GV/ot5XHTb
5pp/pAEeQL6ZMBL5kaZy4hgolx8JODgD6BzAj1eaXLGGW3fSUJ/W9aa4+Tgawl3i
rWg2aawEKKFhmyorDNUx4OY9xIMBdtswIcCeDh0WJ4CCjyDY/i0Xz0WN94BQhKLd
IyU7f/3mP6ZM5jEEWJNiLVOJJ9oPxdon/+W7MhcTfZmxcIw0tkJmfrJLi6JkGmFX
yWtcAqCcYAl4FhnZ8crcFXR7DfxaOagfDpBxFqepl1DqhemZ/bK2gtkp3NHmz3Kd
mH0IjbXVrU+wDU227huiFRc23bwSPvx8s+Mml2NcVu+XlC5A13/tC8G21yqXGnBw
DFOX73WwE+Rg0dfLP8GuRDYmQeq4vwukYJOOnMFnSVuETtc76/GNckV74OrcILXh
7gQuFEPlmvbPyH7TnGV6b3wRcrnXoHWg78XiCAuImkHsAU1rcjuVXbVkObYvZJhP
1nJz+tQ7zjRcjUspUL8dCIT1djlr4z/GyBfBy113AIMBygjLusuyW/DoCs7shHLx
7iBMOAF3oIRB+Am3MnhEVXkSDm9OROzxTCgKMv1ZS3itDh+mvM/Jkqcre1ZZANfE
6uFP1T5oIEDT/r4fhYQSxpJwa5irEmZ0nc/VMlnJ00rbLTjxPsXcHz1h2NXDAOmH
6A0yGq3FtRIdWH5fEcd8r0HD4oWLTJPpNDBSRAK4XL3oYcWSdfSUOteNPG6NRNlh
wRk4dWIQ1kQca8djh8eZT57Nu3yw9s/ZkAl6YuCHeUQTkEJyZlnqMJemSZ9kOEHq
kTlmxEF11mx70ZO91faOGRS4+5uNNDszSMqzC49x3oPjevpDMu9uXdb3fGbN9/QS
pDBmx4Jt8rQaKjmzodqCmT/2ZbnFCshQbzHJ0Iytoz2QAg09jO6rzkVFaInWJpKi
br+A8xe6+jOeoW6BLmEaR/W8BccVFVj5X4q3+ZVuWg2hxQlQfc/MTzhyrnAlgjW1
cIaZNvPNKIIpTC/j8CjGj9tBcJveuVAk3Otf5rKUODJXYea2A+a0B5d+HcYaUTqi
YqQpc/cgh5YNOTO4KbUcpPCxPclGJlf0tGZSNEKnjQsKKci9+hXyQXeXZn3oeA5M
BIYmTQaMPLTighGsej/vVU65QGMhaKgDyyjCTaUi5OFR//wndqKQKYMd6TvDfl2c
HaL0LTtTz0GxVNrzUHnew1jTJMrZpZ7cr/adaZw9c5du+suLa7d0hpNPG4k2usLt
6KnEqPAYmyoFfL5RpxqKQ5D4aVU/cGx13hwc5aCFsbd4xCZ2A/+C+jxSpUC6xACV
T9Cd9ok4ZP2+Hf3itTWeA37TXupmET/YJ6fzFi8Gt3rS4SBW4NcxeCA+iMV+qMuo
AgsM2A03ICD9olp3yP8aJq99s3kLbK3LRRV8a6hb5Yt6itw4+PKLQy/Cx4imcDgh
698q+ua3GjdM1ylQhuVkmiiMbwj3lU0SPKU72eSep+Q7l8VgPYkwikNcebU8hHEw
KQNYCc/c9FB7ZWx5LsgXuL3qywCPdvYo40WGWNzTcVwkGH+7g4uSCR61WGaM8dDs
XfwaP/VBdEwGsay0s1IuwqFsWALjs8TW2N0q6aS6z48ZEmgIP70xMtsa0L6pcE61
meqq5hbB6M+9xYbRcuA5zBPEpXoLLC2GH3b+gc528zG3iqJh0lpPdMYnTpzTfvm3
wzdXYDPYW3ksAC3j3y+sJn5p7E/juOJQ9fpYj1/XMUoTy+5WryXyue7qkOfIuqaQ
5kZQCqFZhOf8aWF8sjlxWelipX7YtJ5pEzMz/nCcKROkKqGqD5ZQ3+Z8z+W2x/Qu
z550bKSvjAZaySn3DgG806CbT4NbiEezbX7+a0LkVwh3INot9tyc3abRUT76IUH2
+RYki1qWZR+5QnzbnEDQ8NO09UoY3iz0O6qIWuIn2pS4L8eszK1Uw52mDa9Gm0s0
Ng23wttwqZUHmG/uma9ohJKcTR4WPc18Ww5FcM8LNSGZPfo1xDU10ZArzl0z/Lk8
f6SAZ51qolYe2P8U1vv7U90GLLwRQPWU3vLlfzg3Tvh6TP1P57kLzbxW1JopnBVK
BPPWGhUUhCxsNcxU9alL1+qm2Y9iFxWB47aO2qsA64VSQUsa2rd0PnmpTwiCvBEJ
oKnnJ9WzLasdSilx+S4GlgBussDkaXsJUbYvegQt1KJxI83PeOVEnqZVfk/24h+V
Q9DPEu+bUyXsF49EWNbFsNHPPKkXazvzSGlTAzZri9z7GmcWfJo8Z/z75NYTMPtq
ojESzB+z4QmInIahZgCuqbh6wd+oWfRp+8lQRmmuCIq6EuRsxskliTCXdpNvXTBO
lF8jqHTvZt1sHRNp7WGy0s3Q427yf2AGorJJ2Xr0fMoNO5maqJlT5YYWNlz1uV70
UmJM8YoctejUmEM49qhL3P5A28SZ+74kNfKd1ilrgW9OSL34qC/inuwnask3DE3A
tEhP2+qagRgRqgojw/92CH/ID8VOZeMPlnIW70QDZYrzB4RUZGtcNvSdzylAXLo1
OQCZJ+CDmcSXzyaMftDKGkjPUXyaBcIvD2ou6HA9fOofiXkbY6ElL9i1XQgP1/hC
gDjJ7NIzN+kVFn1N+iCmt0K9wK/bsN5xD03DcYvstR0kpiS1xJPZqCZdII75lzeD
Oyr/Xgsj0xgFQbuGKvpHt0qz+EVK4cj3mhdjlgxYOZR3TxO+tIY1mEDhbrF1fkZe
iwahHCubHxdsQ8ByeSiv8ttDYf2He+DdsypztUy+vSS7RGA257PZzFXum57XcTtv
fVPD/bUk+5fPJiaVEIryImdUGa6sYnl0+YMnwmTSeZdJzXbpC656QEAMdYgYJBq+
2rewB1BhmMqJAvAXaED+KHIAqndjdtaFzLrMr15tH8tpadQe4gLbAJRhVgRWXwax
jJAXrm0vdxpvBd38VAJjc4xfQWJv9K+HCsRo+gTRqd3hs6C1wnATquBAmShOdrhJ
k7uD/2uvt7AXx5tFTQzbMH1uYLOoOVRDD33sGmUtPz56HZxvgQxx5C3yqTUuNpTH
zaEh7CE3Rab8je/4RBNu+TYxabaS9+IJrzB6JSUMp97PQ354aT6Vhko7+k6XNuYv
nHy65EfrC+BnSeSXgNK9zkhkVnIYsa5DAg4UdYkTrbXFZKA80AaFEHqPSfWsJrsA
ELLFGfbNeGTock5WVE5o9orI5GqL/zpFvRf4h9COZ1Rrw8RnKQFOBH8H+EcVpZLH
rq/0RKL2f4dkxsK+by5dN3EV8PGCZ6Xm6S6S68v0tQt9bOulaT9SsgP392LPSk6O
UhXA+u3iYMgLVypxhhoz8Nnwed/WEnTI9aAcbYRELWgoJeomxCaEa+EoETbzfAm0
OqlIPGDyZGF4sEEKQuk5XuhFIIRmUMyyBu82m/H2T4Hb375bkq2x8p/Sm8CIAOQP
z20kzaTkIE1McbUDW9QBv9M+MNCbR30SAFhDzpQzzUeAPbUqKzBYGj/cxYC8T+Hw
jPxbY+k3zb2ZhbS/0f37bg1yvVRATfdeX9gK98vS6vgh8/G7dMuL1ZCf6UrlQoT/
vP2jM6cl+a3F84wFR4/PL47A+7IRCkUe25KEf6HAOHicPreRg6J4OSoxpLqVNiNK
Pi1zkKywZUj/pQfZhbH85nZxK52cK2Nd/dhRe1qW5gjAsePtvvhOP8ngfVyz5LfM
oCU+0SlkKBxp86toLHih5l3Lvd5rzg8JzTNl/wcRHDywvA6wLlUu/7BOewBJyvzu
j8YZUiuhFezZy912gjABggdCuwsyrUyF7aVMCS5HgYUAJDXcbtz5qFo6JhGNxaGF
zst18PBcIpyVGgnNmjkxepjjmcWcM1/IjtZfYFiaBk+TCAFbzJzvO7yNxwEaBnO9
0pFb25YrQH2Vea+Mkecmfytbd87KeXyPxdejT9Q2r/Rs6wAna3ALLC5vPIXd0Gtk
KjYuOco5ovNsmLISkXDvthUgtlEW6qm4Fwt2oUUI1gYiEIa66qMcHiuFd3+ZM6hp
hzNq+n8ewZGflUCg0e7P0B8Wz637sHXUama4iXiM2+TALvGIVEna9+NfqZfv4D1a
WaAAbfMtvBpxV806XREAN4WFGsbtNqvJqsMzo6O1C1m9S8ttkmkRwv1pwJjmjKJm
Ki1MwG/izfJbBKQr6Ocgrw+OsV38dMDrjoBvD5uylLKdoICT76bo/mdfVAlbLZQh
+pgu4FkDFNt2KIA/f/twOtwetizBSu2f553Ua+qH+JmWTWmQdhz6h0q8yBGFslDi
zCG1P9EVceMSFIxva9JAzZXOC/EqZBBvWMeU9ObcRli0kmIsmBlolkqVx0iC7OJ4
LKvQJ9FL7sm4QO4kbvuhwHyfCZkH2IKzvd1uzqJ8fNxnSzUDAi9iXv+ueKmLiZxI
YnXf8Um2oLkIVJ28scLYc+he/pcYUs42I6buoXwHKUGD7F3gAhQaHFLoEAQLqaRs
czFd78OCfBMPNqcUTmewB5KN7u0W61CoNFtWbkma28guoLktSUeWpBPiNWmLldlf
o2Wm84D8dD8ExxCnW7m3tGVU+myvTj/uBTaE7dgrPsqNdJpUfIr0vJix0+tAxgYS
f4MrQUioOd8/j6XCKYtSzm5hMAmjoyW9z2gWObMKKuowesWzl22p4/Gz0kp7Nt8x
3nh5oNoMGIXOGqxcEVhqIPzc0BUJm7rR6DoO6y7nUzy/fsgL6FlEZBMjktwiykyn
lIHiCI2d4Sf72uyz2w0M9vZaadMBUM7JVNz8REoYxSLiWGxE54u9tcqhnglH3svq
laL1tt+RpVKSewRhG4MWfpKRrs6xYZ/+ectJ7IKJkfT5vYSY3N6gwfsI7x2B3i51
5/lbJ1vpIVjUAfKxUDFjJDOCyTeXOyG/gkz6Qwy6MIiS0/p/VrhUgYKV7usuWIii
hCdcNRrIROD+AAFJvgXD9vnTZ4+S3oskMjD4+VdVRFrHA/kp2UDyZ2uqcB/RcMxK
x7TdWUqiS++OdfSVhv66kzlsqKK5kxL98o5E3VASIPRdpe6ngVzpmg+zMIaxZpwP
sg07ShZ3sEfBWEYJyqM4m6KBf7xfrwd7gABi+rNWgML9t/K1VMaNiA3PolpmXAzF
VpC4p3kr1f1X1Sm4Bu1p22dkud1UCw81KDxeL4SbIKhr5Bfm4m5Eozh2Bmg3d08I
YBrXRixKc6pCjK2yKRASwBEjo8z1Ls1qKHMMEBV9YhP0rSo/CIZisXe+5d1S8je7
SMy4EdHrqjztwlocyrqvfOwsQdjUKZ4Fm3tA02vg5ObHVOp/bMOmNaQ5zM7iQJrk
KaWr8DliWFo5+ug98w0bsOFoeAhNDz2gpX2eH55HVSrBp1Uh41G6G2hDaPwWk8Yv
oqdnMgFmmPGQhY261RfrfZYbPKg4+0v9PwAnWbBhfqhPoA26q7lxo/iTBGWFP41M
IEO/xeA81L2wVBWwV56gggDQCMfFG4/MuQlY88ts+1WzN3QdnF/2L71fNxf5oUM5
V7F+tAtZogOClEIbF9hz1tvGEUEN79TnA4DU9tgILjsU/ZC386ikRaKE/bkOsRN5
dmsfWiic5w9Q2JyM+3GR625GPVNmt22NkcsBBernRRtndvcQDG+pxdw7BXRnRn6s
V0NDUu+dnQQaeke5nbzgsAvGtFjrhcFbxzz9b4bMNHIjg2Ltj+oDKg40F4VJL8sW
Fpx48UTkWMM+z1XlgsQUizHH1XBu/wcew58kzXl1B2tWydLi7ETY2WP7/b7Qa0+9
l9zk7dZNYteZE3ctcl/yTsxHRBhEb0pmmB5R4owDTmbM1Ka7YxUGqHXuXdz4bWzV
6DmvgIng6ZyZpB+qxDQ3Oz2wD6Hzv3e/U8rDvce93wr19qWS/Vri9hx8VbNG21tj
NXQ2/ibAv67+mNA2rD0pWlI+at8GjZ+AkrzQXnk864WzZpWGzgAwemkhj6CJuL2Z
5RghyqV9NiavyICS4C8HeAY6nI5UKu+31WknJrn1QL3s555rhVVVMEubnXpJOkZr
bxCD3vDiIB4SqJT3rWDlJwGPzCm/5LueCmHCeSA0m4daYO9/xnwbO80feOodPvP7
ln/VnZOMu/A2hY0drSvP8rk5gAa/DWZqMoTaGLqJn0jERiVtBimemDf08j2gq4d8
96LD1lC+Ghc7TiKCOqGCgFfCdzhRyiaKxRkOI5oOtCJ8iEego2q87wNQl7xOxwSf
qKpl682lVomtxLcWY86QDu1sqxg6nfkIsfXAvoK2FvQq6m8zzISIqM0xyFzjaqOb
MZjpPpQsOj9oMjgwVKp7xT17WcJkBNtWQoRKa08nyOJzT8/sLzNPAJChrxcB+c01
nL76w1V9VkFg5msecMjXBsqC7yAKAB1+xCF2ktrQrwV2usHNb+VVl988iYieG6Po
IAOOIK/FmIZdST3wtf7k8QHEWajpas3cWXKyY8Mg+XmBeOC92BQnvG5JbasJcu5W
fPQSeKVrZdmCUuN1kHNTltyFIXa4x6xx8+a6tS5sNZxtVZxwquGXskMw9McgbmEc
bdmUdKQfYf/o71C869jUpyRQts4t7/8/v2tdYto2+y+ZahVuyUohD5wC6hlA09mo
UN+79mxmCErAgOIo1OeGmaNb/rZTnFk7xQymFPitgFyyBQ9kcaM/7wXHTB4uCY5Q
u1gtqql+rySktcf4IzIX9Iu8xejdaqQtSNVtG8g7rHz65CuGS05YWubGifwlqlNk
lHM460g1NHOwUIT2LRs2Vxy5kQ2F6IbLe8/dypu2zWtuw1ysv7L9eKksg1AjLozh
RUdzhmyxBX/WKhsEfpNOptBi8DGi4giaOFtVUtt7anzfPrjFZuHP+JTXeOoZyLZr
TIT9OU7SD5S5j6AgQQMod6U5ldg1I4Mql0CEeoXTzSLqbyggcjhcx7gjLCt4aCDO
2jxYf1WOLXIcBnvBA+WMjgdZuHhyR7xgQI08YNt/sEODjckFjIv2krtQ3GvgRvBk
VUeyrHj5FoGHBtb0V+8fnO/SzZKwxxlbStOO+J/RBqiKXYuPCoskrbFHo9iSpPIW
M8tEIQS35c4T4W19+HBKndFieCeCjqHXdpkhATPcRFUvatP8ZNLDjdZnW4Jqaqkj
eLSScmOs2Nbd0yRw1MhwqVBlkRo+yYwUUNmjTcZcwgOvZjaLkEVEeUa++LX3J2yj
dOedIGT0whv6GwaIfQgTUqruBBMK9oF1WnoqkbwrR7Gzl1Qj7ADLRGpM0r8IHfQM
tbxVPBv7/Ushe2j+3yYLab+kf5oyYUz/lErQhNt7Azhgx4uzC+UmtWWOBwc5WgRc
uOWlLuQ4rvHpkHYmv7/Zxk29o3CRo1WfWQJocN0HoKjEuh/lGbAHe9JewHMg4oGk
Po5DveB/0FiUFCRHwwqGvJvjWVVLcov1GOJPjL88iotElj+yHfFacTJ23UhUsGHM
thiiBOSNgFqxIeiF7KTEQ8ywrEJHAwyb3oiIDP80ElcargZTEkGC+NuSIo6fbfqu
rGwOgtXI9t3ncqqgQGn72ROba6gb9WZHMkjepU1GBlw1xFRW4B0nV8/cbbDuc782
ne4pAD0sGY8nMFxxQPl9jrJxWNxvf/wt1xBHbt2WUoILT0cYklOQrcq4be82w6LG
qwz7x+1ckXoG0ugrR1xTHz0XhcsNORKX+Rc1sSgaZLH+UjZxSASjoeUelqLhFCjR
7bjn8pzUprEtTgiuFOJITwJ/s43r+MuhzY0xYC1bR6JMvXW77vOOm8EexuB0xHPN
V50xdEjZiIB3a8lTMhf+joVGKDscXc/sgRMEdhcDxMR/HWBSRCjyWHkZ4MNUWAnK
de1WmEhT5MUYVCqQby53stQMB+wnC/lSKVj/TcOxhc6T+fXhpZgrAxB2fXNZ6595
JFXkCu5rIMCvLDIZWrOXiLljycyQHZgDkdSDCQAnPwz0i4GJlGi5eyhxSNr5BShN
bAPjWPFI9QjDXfVJzqtf0RekIjR2YCPyx1WPsQUIZfq2P3X8I+VA2Zye5w2rvl15
hee5OONkxilwGflzzhvHDrs9JE4CI1uS2UgY97sHpdOsmn3u2TTYfwpOiXxhnsp7
JIPh75roWEp+EBrsKHAdF3oUh0Q/knMXDLfX6LD3lKLnGYtw1RtQ8d+kfa5z4Vfy
EImmkidmYwwWdFRBP6i8tab/+SMoLsYD45QapAg9qUARdHEiCK+IHAA3ZUxt1lxh
F63cvY8MwycFN9KDdppeP3tnfp+3apVARq7qUsd7sAPxGEmgWzboaSKSGfVDz7io
I+z+tDeFzz+864A8R5n9HPdeR9RUwiZHyezz6Ns8UbgH34yWBI0g5lcXJQdG+6f/
oiwE8ywXRMSj3O8Ds+0O5ZXjL8W5HZngBpH4nQTby+aFzPOjipw7tJhW6xLBEhTb
4HuQkIKARbBYHftZcdQJ/hBRhn2sUlupTen6NekG+b2ody1yXSqNHDZWojxjeNQB
LlSVernMbLiL1IlA+ieFkwIUmnkivjPi1WuJziZV39gkTIrYbrNkt+cXGV3TOrBw
PIigT+CZYQMNl0bJhH4pVxeYKWsaZE7YEZWysv3cW+uYY3jC1zROKPAyt7mNJTHP
Kb8eury4ncjOxO+ou2XBztQXGBdI611ebTHpg+8fkjConrGtQv0/c9kAc0bUdCqT
bPwn+tc292edKtwPBusCnCVsA1XTjtzrPHTH95mjCUK/5XyHxOYtT1JhGAlHQ+A9
ZluXS3eBa8FskAb7OlELXYYJClmT7eovQHUrHT4MYpwtVsr1+aRZ/didlNg6oX83
0mitjRxkmRWphW30pS2hR9VV8oySHD7xvu5VJ7WvhZTy51HF8e5pTBXtVev7ndRC
a6TbQXaxtKLj0pr+0bUCbaRzEAA9XbkBYaagK+ZNdNSI4j11ik09wYdf1PRzDpuw
Vyj26/Zlc22QXlODISn5Byo6pNYUiTqiM9Qn3A1yXJe1uZpNr7J94vr4NhctbKu8
Yq1tOhHXtt/urd1Xtbg1ua1tlar74Sh5+hng3xihg1vB3HL4OfDcCyvUml/6Z4O5
oa0qh2MDEbzjiSnt7KZj3NyssODEJJJpXTZUDNC2Evm3zOx3S7JJJokSgJ5m083v
fAhJ2mVxZ3NK/kbFNBH7ylWRcUR/USUwZWtpVjujN87+svWYmwpkbg0pyoKbQOlF
/bY605aC+g7tItbgmr7qICmxqQEI+FLP9m0HYPGVeSLQQmDAJqm6V9LdXzl8CEvJ
QoQtuLdaaFrPGg1wENs0+KuovSeBpmv/uzosfYbXGk9eu4DjADcmGz+2/3xhze3L
+MnIT9Bdlv9OPE+VKB/kWnGMwec55SjBP2DeAxWDqIMU8ITUnLT8efDQING1/gU/
XfM72m4LXaO466usrDkIaSH0+/Mgakf8ACqTRD2WZAdfxnFzR1JL0XObtQLbGQiZ
vIyMzGGZBzx9JE14kNkywq5ht1KGvpgNO99JCKLRMFUFactANRsdEnreq3DIr8ni
/Z2WTKjIMRwymom30Xttl6onFrNTH2oULINWmHaEVIk6qV4HcN+JrCIgDlPbN4C2
RlrngcIeUk+/XWMrI0Sjl3DAZft0eEXoyxqBSFUHeA0STheQzjciRIgQFQ+1sZGC
togMuwg/cMu4k7iM2xvdksxP0YQhT2LK7FelNREgkDt50zFTS3yzazHaMcSQOLKl
TIjEz4EaFwutQCA4HF0jKutkji6L5Gb5K2V2AqNaiyx39cGKCn4SqInYytxMRZbI
efCFMlTuB22f7tEdMlh+NXP8QQZLahdE8u5QDtjToR/ZWpVtuatRR3I2q/tL0dSu
WhTDejukMtB+xYJpEIOqjHVtavXboF5TY9SYey9zBMi9nonuyLkO8CIOIjx8+IZ2
LJrQq5L4xbe48rC+ZyCnaON4VnT8+cRGIb4i8RO5zrOQVzxh2R+z+cpuAoXImxdd
9ArsZsd3pOLqhqd63LttnibtILury1mp4qVzcgcCHsxA4uIpJ8Pb0NLkJOhcjhlj
gJU/DdUkEMM88NInKWZC6WNfrXJgkcVaokJvKburQm33pwL4aGUd9nF1FLmFRkvd
GyKUcUViLdD9wtfXvhRY0n3UFybvKfDFqnYhhdG85IgZoYSSOrAqLB+5zudDzHGI
RDxAMgukYDl8LRLNpmTXpBCdVzPIiMqkuzKrPfK/7+sF9oKAAlXGRX98ZJuhUtPS
TzKDq5FVcnpx32ZrtKTZidjY4yU74V54xlNu7bySeoQFoC9he6mY12Iz6T1DwXx9
DxCz1lJ2F+FvQmz/z8E/vWXhYcUdjCsLXLXOE4o8axrcifKlAFdpZNpcWKqH+00T
XoV4Zja7FLcLTLaZgRiIS3pxzBTZ6jI+LRscdZx67IHlPibC6L8CQjqeJhFl+5Ck
w8qtwpAgi25ZasJSU9Z/vuc7ED6B4wc2MfoBWmIaL102aGANZq33N6ktvTQkwHqD
qydmvFE/02EpsnjUgPzraVexJc8MSyIM7icpSTLNn3AOWfc+W2/UCvzfFXdQsQpX
FGm6BoFeCBLrHwaGgcJ4E0FfcRCVVhxZMDi45Jp2e1oQ6GuOhKzksbemra56XxCW
6L/2cOghL8khnpDvQepJ8B0BpRv2rVSSAyPAxOimTPBe7B/UGyBuMtuXmMcTrl1g
gTfmZvZ5DYJxEWvi/Yl34z1fnNYEWXXAoy8Jy0IvsyAuVz1Pv7XMrpDU4uDgXiob
XTJaNNMYuM94i4PmZRswIRe72U1i4Lih34Wx+wgqdRjSI7dYGU86kWSFVsrzFnSQ
+r3XBi+uNG6P9hgWZfrbfh42iCmChbMLDnAbBGIFEUDQuF6HEx0+l6YCcvWgMeSO
qwA+I7LV16mgcd4sSqZ/USR7/DKXvxwJ2ZUVc1ft5KWY+bkZbvavlydu5p7nXMtG
mTFIZEhRbobk2TyT7by0Smgl3U132C/tTFP/8ONGtXRMmSJaLgiGaZ1ZEQzlYc2v
VhIFXcA/OSv8m8JP6vF5g/rEEKAd88d0D182FpgTMQnTlK9sYuqzkGfqqFLq2b7i
9ZqykzybI6Gei3Cgg5VuZGCEb8F4AwecwMTQWRZivC8g1mVKTFKoKWdqDgdhW25d
1mUi6wjQfK9/LDkEvgHgiZDV/F40kNwJfvKWmFHqNjHqU+8RPnv1GApKnK79RtyB
nNrhSgRG7M8NebnZ/Dsys9vujByCAPk97f4aLSUueuCNjTO7AyUbD80txXs1BmWb
vID3Z4oNT/DJGGFo4eEdhU1dsl7AyGQX8rJLK2kG0BaliKAiIv3slcvv9JZ6fqB1
6/aRfcMieEQmTnUYGQ3fw4U9rF5PL0B452ECPD5ExrZm/8aLYRXFErxdzJMH8IQZ
HZoNz72T0+K9GeFiFJ7rnOft62AB4iS65Ecb1Si5VW0jned63xA65nLbYz5n7bKV
N6eIwRTi88BSWhuwiTRUBNO/aQPb2m5KRP+xMpcafY36EL+hX5gyvD5PCjFCfwuk
hZQN2Pz1+OpvBQMqFyJ8wSG6JtPAKU16nFKdRc2OH/QC1Y+uueV+2o55TLOV20Ps
F0CeFhdq+1M0AqkVzVlPc1WD1f03fLG4GaCicBVwBpixn8qEn7U77OsZv0Uef+SF
4+mZ3cupY7RvaI2X+oAEfAbslkjhO+qNsw1I/QzlfF95weS015CfYhxZZvRCr2pH
yfL79ohk6snhHpoMqkMaAg0B3n2/hfdfN8xsKuyldaVq3Td2QMfBs0EdmRL/hKPk
Kw+JSAAfVKnHb7veHVpc55hnz+k2YlXSIeW8E26jzpdznRmiimbCwo2HLdzyxyTB
c+gEoAquVvPu+/dC9TFPSaarOmSuExg2fHol/o4kjUo2K7MMrU3m/mWrXQTHWnJB
YxCtLnFswrO3ZxXVg4Wq6Gwq7+LAZdx8GMXDEI28QZxK7hVheyxNh6Wwsi1QKQdt
ziixEAZd9dT3RahKLwfTU1W4jF07kvPiiE31KrXOkJkqCqpWnouLRMRAPyTLgBjR
8IWqGMSFITTjYO2yfQDDBw9NRRaFvxAfB4/Phm/Dzelpj7pVLCQ9lioqnw/fideY
ikh//NWOfgQCcBPJZ14MCkxNMPMYpZ0Q1/0F2veuhIiM9aKYBSXqS7jimSGfNjg2
I1dJ3eBDSya+NAANgWGwp/4GsA4GBSwFMZqb2Ny/8kzqUIuaM8vuV2jq/KmSuGVS
8GuCZsj1qnGmTCxNrM5BwQVxvGpSN4i3RktZaZ8VmAiU6lfVQiwOYcYlzxeWwfV2
EUkybHDbgReOVfX0TInpyvHyn7nJTiN5l87+rQ0ONZGb6KmoVFiVSGgQQc7GxUfx
YeLG3ZbgUGaXUp93z3VVdh5ZcptFd6T/ttlNiVh4CmnO+c/HqHTOpguOSR618abP
XIVsC+LsSbeaSsLahyb/9CXs8o1Z6tr66BfqM4b0ivoHlFLt/C4J0Cp/9wf2k8SD
8JKotLQQ8NprfoKmDMlQ0lt2A4jEtFLvDSKOSH5HHYPe2bOoMB+PgrVIUneAXLZ9
cL3p6f/9Wx0T/EOHlol3PYsMDGw0Ulez+IfNxgtzXElPwVQGZl1THodZFhwutxXP
GmPNcXKJTmgoHb29d9mFeeMleRFbU52Q246NKvAFBC7hx0uf0nzeJhkiJTZFrR+0
LK8IB4tqw5SUlWpB2BEpb/+wPft0ZQHmzUAhPRXk56PlmQxK0NwF+uqOnwrMvMbH
wrVN2xPlthByox/99NLzYec6SzUICV8ebFhfsE0sr0ailk2hmZ0FQ8ydrjxyUQYa
OpQcgX2X2HFeJ07Z0wJkPQ55UJcCvGwjkVNR8jPO+XEuYwwk26PamqWFwb0lcKiI
ccD0UurdakQAluiZLJF4NigQUWv9uwbRzf4A3M8n/4dFV7vWtG/ryiWVjZr3w6lx
LzjxVgSqjjlDCfDn8+jUMwkAKy9+ejKtdbzAz/+1jslaN9VKyOsIzZqBCiI82qyD
06n7vWo+8ViWaBhBxLjLqi0XEiuWy6gYKE0+wL/zXcR8PjmzsvzEeY8auwcdFEPw
0d0Fal1bG7U3J8E+Y/8C1zouKGIRzRyIc4GlEirMJfn8ATqc5qqezbDoMXCatcxv
deZaaxVJiAJ7nBG8lGsNqccQe1MIeLjRvLnSKP6fjEuPyQEDQEtOIM/G9xvQokWB
k4xZG/H1yrAXFUZZLbFx6ZPmPqVjPh48qRoBaVbS/F4V4JaY+5GtfOf+b8ymGhi1
wQ3qsGLehZRFDYFVKsJthtpNiqrRbJHnBoe/QgQ1reRiYLB+n4H9mx32ADwPkt/c
lX3+OGFvsKkX/5HvOrCNSBmaG4Ch2wdX456w4+4qte0BeqX6t1WF/QA0k4jNyqFA
75eMNTCT5yq913n2XmNn62dLhCpajK5ng7t0+TcUR3KfE14Z5mbZAa15B5iGLIj5
+gkPQT9uymw3NgY0pS5eLV/E8m8xi0BkQCV4w2zLQOg9LkY/GyhB93Rz6O+0AGid
VOMFZYv5snRnczgKd/1CmC1XW5Zo+8TIpBrLZxY3GzuNHlvi5gwKAyTUDp9Vtvbb
Y3hiM96yqnwUo9lKBWYSTXER+LPgIgzPmCYHJ0sZMeFSntHSz+8BGnRr2PfzEX+g
vhGHlFSo0af4HaJ78vZZnjRvzblBFup25A2mChmoGzVFcixSSmIkTe/evVGge/Au
dHwB3xklLo3N5fkWlNCf7qNCUiNhnpEJmSsm1sJ3HSUzMa3Kcu9B0G5Oyjexq0Kf
eCOiEZk2Ku+oZuVm7kcUDKw8msAT5Gx0SdtylKdD70xFGeuyN0r6Ev1LQlhed7df
/clEnKoh/hbgPEkrZgTDFrT6jz3zA23BexJiQtlQLkBM5qTwMF+fbBFpi0zw4Lcl
y8nIR7pGsJz/+O1A9JTQZ2zFNWZse9BQZghb4Hbb2XbRd5/7Rq3PTC9dC6CUGEbQ
xEVDnIyh/Q9ThjUoDgSnx3bZnlsM3horAbyMHNIdhQGyLJSXFMJFWRMDV5vklvaU
Cn2/pfBkF59JnXHeMYzSdmf6potzDV+9Y4muA0udlgKSXnJDy9v1gcp1h4ytJDj1
A5MbTeTD1kDUcCxxbC/ZgXm5ClLDgf81eUziJiTe74CMO/Xl+ttm2fgQF4hqEHql
quXFFvK0MI98jj3rCKNc5AIoyc37vp/uFg8SQLH0LeP+HZtIBgX5xeJH2aT/6tuA
oBOiDHAfBUJDNfwpIITif0a0veDOWhV8SNprT9f8p/R4sSABQQIFjhzlev6Mltbk
gxCLeuFoKUNqv7AOXzQPCyHaAJrIX3AYeddO71YSwO2nIPyd7REb+93GrzdaOMYV
6D9BJxtDNInqKXEdxVBuM3fCGJw4PxbTCC7py4vQWri4mImLJUWvFtaGkyjz2mtn
ntE0O4Bvcs3yEdXgdMvFjDOxKqmHoOOJHHTFkviFf9Ge/Z2WOEz2OxU6b3bBFwiL
DHCBKZLbuWEIwa2oBYfb6+MYE76Pp0lN4PTL0cIaFBK0iLxwM59DPLvlPD1ANNfP
yE4bBP5rgmStD2G2fCKBf1QBlr3Bp7U6XmHjJKMi6ST5Ot8GBhp1Lf1mpD/x7cME
FJj/82NoeHY+ypIEYPQDQnI4EIFaD6ElTTET10rsUk4KAiBdZfP/8uwcQKbZG/d7
Cz8LLhpmJlewREPlqpaBkuGYPS4pqnnrNIkBEZLM3WaCElWDT5Dz1lEnzFiktzdb
wDsd+hLkRUilZcX/lpYHV8Ru+nICV4uq+6ioZSiL26SNKbPLzzdV345Zv5qbIJh9
BP4i/4O4M24e6lB+CYBZ1BkvUsTEUFC1Y70bLmgZuNi5PgYR96crW9thzJwtHy+L
6fgGItf4C5w1zAs+9kYpgJQGh6OKCgrQc4jeLxLeLIFsFzeagDM/jpjtvbG2siHH
AeqFL25lpeZo1A3XrYkKE7O301HPSluesLgLHOTnLsbkVDKlY0iPt63ITZ96+VJB
R4IHu9FB5Qb/+upnTVy7VMiiSUy/5JhFrgzltstUbzUAnGCtl/+hCyJjp73zd7ES
r6TgT6KRz4igB3abQX203pVq1CfEirAipOYLWjZZC0TJJDwz00dYmc8MnYqw7qsn
vgDoNHuiu4emoxtKksxOxOQide9EI5JM3BV9lFOhs2fdVNTsUQruju6AWkJ7PObD
JXgK0grl1Kh2tHRVujpH5VXv4ExIfArvCoqRuyyFKFzIJfWvBpFX3p5Fzmb1QE2O
yiBL0r+KUW6TrLVBvpyWv0BYg60tfzxdLZs212FLNHkEqj9T2gDIdPnQiyW7AKXa
t1IUqnWjmCZlvMYp7E+ppnwOPSMfsnIRtHHQu7B6Gimw7L7mx+L9+Sf0nvB9znwt
LX6UwO7P5H7z+6uT3UL6R+ErcJ3OIOxD66HmBJhH7gRdSjcv0NpLVHfvhkLbbAA9
RTrlGQfGcpfy12raWjK7d9YOGGY3ELkngdU9mEyO+/JAHt7izJjFZua1wEWiOc7l
2ksc6/leJy8EWdjFo0QyXxKBRX1sYZvmpUg+zNULijm+YQMUuLQtVJ7BE9/nO5Tu
AjDmO4wCrgdZE4V7Yz+WPAWAoX+fH5dmt7GbxtjQhyctl+nyn9JbirichM27mduI
2jn0QhUGlK7DaJ8BIJVQzh8oln/W6lCocq4exvww4toCeIZBBEbsDnOJ4HrebhGN
73x2srVconwIIKXi2iQNN5MhJRW++Kav3uhlW7NgEPjIQnogOO4gs2Nw9fLFXZN/
2w09omC0mmxttkqgNomW4UbIB8rI4lo2CmdQrlBlDV+pGzpaGlvBOzvafKrWIjwu
KLen19enxvH8drTu4RXrhlsw0547uLquyayGS9Q/D5K4syN/eiFoS/lfyCveZqcP
SmYBn20EsE1xZMN72j2+5Dr16qp+asteyhVgvuLZ0rFzCQHZejbuQ/o7fvCgHtq2
DvKNajWxxI5un0pu5bjCK+mAvwPmog7lPiJM1B0rx8JxRc/Tt+6sZlM71c2WvdS5
mb1SQELcx5h+PE1Y79G3aL6sS9N0zHvDhhNSoajBRlxXXvTYX5QROJqk0i8TWW8f
S5PwExIUE28PrBSsDUsZ4+3HqxHnJg/vW1xbpCuz5f1FR6qwa4q3WjWDhKoKSHme
Biqh69gk6MCkjl1RvL0pVkhvrWHfYR5WhIuTjCboBJlRAotLDNpFgANrFizpsLJr
yvFrX5+zDSNVwNsjvXoaTVS257RAcNZGQ5ndD115/HWi1jUXEroXsQLhXvYVkJct
xbTNOGC41zlLE8sNqZPTV+ENbZHDf8TPGKG1PtySIII9oxNQo0F7HEztVoxSjlj8
KDtwiUP7o8lKV6oIirnf9JBI/HaRbRdNqplGRkWY9G7X9s8UGguD9RG7+7E8wZ4h
P4qZLgtsYpN1EKFGaypZH0899X7WuWbTlu0i7qqhEcZ8XPtnhwQFMcgVqTr6vRBG
kZl/oROleS7LqJkv9t/UpRHyHNL4W0HwCFagSsvPo+IxPWBr6NVp+X2+7oi69NUR
+rDPnSS6aXy+aJ9D3VUEb/3wG8ggiHAcEY/HjYlSOeAGLVrFLPZBMfJLeD4+6F93
WX469Fv3gPKguieh8v/IOty8lFixoz9EtWgXmNhpGCSI8xb1lFSkViwtKEhifWjT
yYa9AS6pU8n1F3SV5abB6R1kvDNgSmaSXrUnTiBKk5c4iI8DOd4yNMMAe408h+Cz
auIEMMQVMmE70mAOv8adnj7S5CsMUigYBYJKnfr5aLgwKAvwdNOe60P2bo6fQHq5
AXfqI6fj9/lY8DFoTP4xvkqZh1bA5ym+OVtUGICmkdLZZWWv89s0Fh4PviDubWlr
+LQlhx+VPodunQGBSllbI4ezcmDPhjpnItPc/Xmx5sn+uvPpt6QvLK7lGr/UINsf
VO+djpwsFFI/CtHVchr7YabEp+lBjgSxYnSvoKSqwdBpVHVuDgt3Prbv0DWUHpnV
jE/W6UER0mw35+chIlAvVToP1tjT9K58gYRLVPETquDJlNvBa+V5PEeSyahElkj8
GUHEDSGnbfCdFVaoY9oNTDKIwYOCz9zghVmq6oOIZX6x3slVqmxq6kNbWLVlDdvf
3vZkrCgl2e+Q7ldCDSHnQd/uTQOaE9XWymmTUYZBECIl8N+9a0PPUVr//lZZqQyN
2/9A2e4TqoJ2HBqPha1HJYQUsy89DXHvVKVv455vjCEmEWHTyNkX4iGBOxm8kMqA
70bIuE6xx+r67eZ1GbEDi9rDaPjXxQBE2UoVOhEIjB/2Wheg0NCcuy+BQEtXz8uK
KbiCeb1TMQNyu0L0qkZpSTaGBd/qsHDvt3rYEPkCRo9WSa5YoSVF5PrvC7obvdNd
RuiOjCSUVdvENuE8K6Vlj+kZVJl44bcBp20T1lZ2ZSYB8PKsCCtH/sFRrkH6lyhi
96n44rT/4q+WGOo7R7r8UdSF4avjaBLwmIVD19lw89AsUo/wt7IodeueIc9M4/AG
1kVD45qgMLhrZh1M6nvf0rLJg2f7rb9LiDR0OePvk5YhpxbkfEg3Psin3OOYBs+T
MsHAqI1kWHtGLte0tlNyiQpS0LAyB2WEqWUHWL9KlyeHGPCwM8kIU50LwDuN/3vB
Rk8AC00Qt1IjKUutC5B2fP+FL4zFktrMMpBLvcJop2nJhLBKFL2eAPIhjrrRePhK
r4GMOZdA9OuHnb0GpugDi65SZDmh4QSIf0BPiMrSGc5loo6SGvYMUH0N/yDL1OMn
bNEyVV1wCiCL44GQ43BvCDDWnic8boorliM4yDOFujqMjEx3X+rnaERyLXy7Av+n
AMcLYG92OOi3mFxrFE+boyYBAfteLChvUg5UBt4RQ4kXrNSByP2l/Ri9ZJUI+GWe
6xwfnGMOEnwpfkLRBmzfk73DQZKYf3sYQxjkYBht17z4GFaQyKdzz9lHHbEkNGyP
pLGvdA9vjPFOqWkpjc1SqCp240AcahZ1ivt0Tk+P2VcmYNBI6mbVNw3pDvNtgdiC
1UrayxPjrYUaVSYp95AGj5gaPDcMyi47yxdxDsILDpDhyxFCjFQaoHSY5f7stH2/
VZNw6mcZ+TJB91y1C04X0Os9dvyhpKDBf6K+ULlcTdtRD0lgK3uRLRsxcUivBo3x
i/V2fKHX+VECXltWezlU9cMs0E6O0p00zNpp8q5EptHj7PiQErspvRlYbzp9ujh9
NHxhNeu/AD0L5G0Fgab8s9tx28Bd4nLkYSgA3ayfqKEA9jf8LpkSgbALmoD8uFLQ
1RXrP3m0GBXHugHayt/Egg7hZFv9saXySF0sWMWHCX3k8VFcSqIziC/nDQW+NSR8
egud3JpS4NFARkGxdVLwUhhaQH5bOTMoRHSPzz50NOHrXqEkznoRSVnEJIcR/RH8
OWqYUuE9H5Y9jofUWRCFgq61pNzoXo38ZuRPRFCeysAT5WLC//06EVgZmTX7qr1i
xXxMDZz5feNfIG2cfGCM8vfdl33CQiCxVnY0VwGO5W5+WUMtNqvNT7kiWjZax+hW
YIIoYJVFG7yg2KHeibxS5foRtq1ZPShxSluGo13DgU+gyfpizTRrcQZs3eFSNOth
s/0CYnab4afqYnnY9nUGTCZ/z/aZnH9X5Yw3l0GgGXmGBCm0+RWZ+PLCrjNegofm
sNkDGkX2nHEv3PQE+Uup0GIkTfCRxxtxogI7Lc57LL5DJWl4bKsI1j6onssxW+H8
Piee84Gywuow/zH9CdsdtTpeP8FdO7LdIyKynD8826ds//9KTTDpI0hKaoztom9p
0XBFcoqHg/ugcyPvBXel6HVj31l32Iu+yJcp9cVIzLu2M2sHer/W+pwiR83mdPTT
3ZSG5+Izm99028Y3byAFy71mGNW13PxTXof+kTurxbmZHX4JESwr70YM9rJFuf+X
pHCl5R+GEW3MPp1wbOOD4Oyx+Y6xymEUpjDmVm+N93KoWNx0w42og42wwQEZrf7h
R+/+4t09QZJj9qhtFm3XTrnBrES9CVUfNqqYhZ5R64+xURkoYHlGIkTNDoyGPXdl
kLcTHHwn415VReIVwt4Ce5rr/xd2AXkediHHBJC+mwD+EXW7kN4z+wvO8aJSGk7r
qFFOM492IbvmLIdUnAaU6sRoq02WxkpV2YXsLgHZQMHAMW7BeqZNUVtSLQzSdhFn
/OUVSYoh4lY80WkgWC00bWQw94rcZk07DlogcZMWrkh05lYUQpIVEA1eefxQ5PDi
Q8UZvhdaXPNlp4HqxZ1JFw2TaBrXNDNSqbQZAb8ItgbyaDMv8285Kj7qSYp2owNh
UblDS9FNtSvDzcpRc+mxY19CW31wOOgEsf59P5D+3ZJjT/zZBnwtVFU3O7kDY2sC
Tq9t8HhCkdsXl1Ux1gFiAB1Aj7UH7aIg62tI4fjae/8DrQAqKETfvUymtdtMBjTs
d7R4oAs+vNtgCGVhxVA+bX3hsPn0ggJoaLlFufFv05QnUlJOe6t5adAP5JgEuFxd
HFrzbhaqVB2qgXeDRzT5vynatdxHznGa1XFveQ7DH90o1KZDsQDQkq67E7zgnEBs
QsCH4NJc5wccYbXOh01v394u72ir+YtRikenE7YExGn0EN5faQIMR2A+Ojg1p9No
/b+k3V6nq6f7iem/6nMAj5037Y/LWPnQftjx+4z2CjcBI2wEynfaiCRNcF88/S16
oXKP84EGd0aWIhtutkUEWwIPFZweZ9lMitzxZbn3/59KkXNFVCUN0TMCLd6YulHf
jKsq08ehu0Egq2iIPpyIV5hHWSlT43auv95Pw4ghkP1wb+k2XhIm5nivSqNiT9wd
4fXFMOAoVMLhxAKzEihxbvuFhM17UUuRS7Adm9ZyedlMG39AzkH4FH8ZAhtBU0QF
n+WmMfV+Hk3fVsvml5gF63iMZzb5ODnB++nMr0RHrOz0PtVmnHOlgQpvy7Y9WDix
SS9mzKY7PQMhQW/BGXWgV9k/7arcu1r/9U7o0FnasO7B5UZ3cMjVq1tE3u/mSoUK
l/G3U+JEMCNBkgUcrsgbJO74bFAtWsMY87ln9SNhxSqUiwJN+2LAkZJs/wSp62tk
ETGT/ALX3P8txdL5oAPn2Z6X3PBjU0HVG5IVMFoQV/mkmm/WjrRDthf0VQtJwL1z
vVoe6lx+UhhYsr1tuGbVW+ILp0ZW/u1k4LHDchuImRvalQsJ4DvjUIUpRz4Dt/yx
vtd4hHC1Hg2R7u+d9/8KBekboAaGJ9p/cmRFzQmeG75e9bAmfwGAlN1DnbdMFB/g
qwDlY6v5sDT+pbRCEuXzCUZXeXgYxJAWjwIjmxa712IBECnvfJuGU28gbgM0Sl3l
QfYjzPRb1fAzlBIKG/yx5fJbETFuu2dLv5FTrwuILmMSOIDjqyuSdDXBVtpkMlHm
zi4oRBHH1s8pKamy+tAk9mvwbwJX9RRgn6aIlC/L2hSXW2mTFImxwOHATYD5trR+
2JmY4gH6Xss+dOc4epdpXApTNuYBXVWWBjNPDu4/7PCsT2GiPHO18AS5h+sH4J1z
DvHqmxJ2o1th/c2WJ/KK7hhwR32Lf1ab0eXKKF5PnBr/uXCmoa6heaJRY40ZD7q4
7HIYlrvJ9qYOFqI612ESzEY1xLgW4Dri08S+gO7MFmOCRfAqbtcbcVOQkLnP7Ci7
+iahTyDitKbslqmAvcfXdPh6FkqDnWSYhr7X3vrl4WI+JQSM/mloRC5GKwNnZ99D
UKtS886gNpkdMgxopti2VPr44DjyIulguSHG9jpbrTOaHuV75k8sNNBSknzpndvT
ElGGKyf04EzCCrU8UKRD3ONJyW09YuFuzvAoCLCMG67Se80M0pMkwmHqW5WNgUTy
8Y+suQnkeqr2zwhlCAQ9wCxGU+xNX0hG/0StzL5J+5TKEhkB4dYqdEw0PQxpddRo
qcF/Zz/JGGdXbA7/iqFB4IgOg7B6cMJwPgMaqXgXxIkw/xhjvZ82tlCSQxZ7/UM4
/h8VZs0uRh0QawrBMVSOxAGPbAQql2zSFnpaP/RdOK0BZ4osc/lUeqO0OZKzOhCo
Wcq47BMTmuvBzTsWFrAGjd+yh+XSo7oHRV2i0VnxyjOYVs9rUAJ+zHVgDCawoW9r
An+nFSVvI10FrT1GjFTXQwOMcL2AJEJ894dmD5t1veMv1ZTljsaXHVYmayJyzPFl
zlpN0T3qMNLXXsl+EEuuruoTUWS0KZUtM29JquclRdpEP26R1G3tWXER5auVF0Uc
G/izKKlLiWLCDSwqT8PXkHFwDoln4Zl9ZxfjfWImHUKWdtaQM7tpRmcSMeCMVjRw
fJD6LuuoecamBXwgzu1pBJt5ujWX/e1fCLsvxdVuu0mmUp72rnjFvhW65AuSmMEe
V+/6EWSDA4IlysYrwJmveKyZG72XfdX2/nzOf9Jd2TJWfkuaWvijoSgzmpFqgjwU
utkPZLERHKMqbaUntPU/CcdTJa20c28OeIGQplsiFEJZ0IzWT80yVSC3Hj5hwVvd
EtmyjDPqhyyhC3J2EtQlzHNnZnT7XMwbUkPTYD/idWLm1WXdy41bIk0sgkLaaXH9
7ANis0z6hjyhhre7AMrfS78uQpp0wrX1CNYIYftalRwbKAY0yDd14jtnlzfEinHR
K+MGOSF9tBBfs25SyTxAcQSQq3l9izy7jdkE/N4Fe4pY6L5zZoS+AzIgbkEdpvji
qTVI3xjSRKxK74W6NSXtsOkwAtB6BICvjSfFSElLUSHlulKQ4WacfePlId60W8jB
OZk/KPRo+UzFUV/KQ7QDRp3Y/W5+EfZx/CH86N9L9LQrM5206r4aP66SlmFkhrNz
gJo6Rs7a225rN9IGGVbveY3H2/GjN6mT4oFWvBxzVeiE+vrGE6+Ryao4hINiJuDV
7ln25JKHFQMepbSEIX/hZC+GpWuUCpMoihNmhY4aZx1vIoRFav9jHjEVTmKgBTUa
0psuhAXrqDqEMYRZmc6tHxBeLGvOXNxs3lV0OUgckOxS83zgdR850I9b+fWBjoqY
yq2fu3PdbSTDy1gU+P+YBOTWPYHWmgLzwNXXMJLmJKuOfMpWDQ0uOiACk2gL0wiQ
e48rRxVCZXOagcQ1HhN3Qso0Xj4kpE7KeiPVAvLEKohCKqkrVh3ZuyIeNMQcqB7P
cMfyotDeZo03hxDY0hupZwC4posHzZ1jRmoYI7JjDYhO4xdFBMb1PYieYYnuQI8F
uvY9K40zN+PBU84TMNQL1gjcVDKrS5KKwK8ruPyJ5ZAsUKvaLr7jQ93BiFAjlaA3
8xDNtTIYlGH+WEAE3dt68WjkR9P/Gw9f9WhYHl6pfAl9lgyP900tTuE5O3flwK2H
5g/UJuizHw8ko7qYOtQ+nLzXn1odHFnkqzgZpiWw5zStMCffeMhKjW/vygjGrx7T
NCOgQFK23fdIKiXDUebV3wp+GD0lQ+86ZNURlbQVtK7wFkfXyCfmfk5sUqNTLJNV
F3B9QnKVWeaEqysLKt92YL2eWwwTnbHlpqwSyV6tUkJpfKN03eFcIc0ry1Wrl4e3
2+OSc39oJPofT8+7J/d0vtoHm42V05blmeBREER4cHpAP67O/QPA0YL/emVlcZ1I
avFD2F8wU/FAN3vdf030rWz7+wFpu8Ztvi9IopLWgVdDqIJ5vKx8WtQPi+IsC53j
+ft4ca7vrkDuCZWjynKiD3jeBcx6Qj2LON3y57qGnbFREdJGnF8YGanEcYqZG/k4
ITofyIWffr17EFuMzTZbDIzbnxf2kvODN0HA4eR32gwj3G8XU9ly6ntuk+ZpU6SR
5U2y7mNYBeYijtRPXxHz6c7RFZyN5DV2F0Nd9BGoG2OxknkoIBVxeC1bUoNMX53N
vLeJOXxwbBCu/9U60R/X2PP+erY5ONjCroB/wmxOBb17PJLgf7vE2Bbg1fd+dkXW
YqOtBVvA9HbXmODluuvmUktKOZQztmnJrGD0JMGvTIrc86zTb4b/wII/+TT63gAK
3eRed5G/bkU2Js1hzKfjolRd8iZDyR7FbeWXYTKF30KraPYDzsZP43+QmaYAWRjN
MBrIya5rn+C2IMNs2vtEME2/6vGALkbTyUfxumZ7Cr1arEqoU6WZ/acpfI8PxZMs
5FBK1ZOn8YOmIvf5ON79r96R3z7A6nTQIrGOHUGz3ACBdMLj8hqeRmWMfKq5JAJp
lLlWA8ixPTS6pTD7LDI8TLZR+7AorIFozN6XQME8hWqZPknrnwUOjoIIc9Csbxwz
j8MTgasYtntg1oI8RKwfF9sOVTZ9VIEwuusoTwv5a4PDOPzgxxtq6704v7fxKD63
VY0BTqhru87LDpMZI9aQ03i8HzaXzOIUdQno818wagSPVnA4z1XSGVWnWQRt0/z6
dw7DL6LgqDFiYqID/MZivp8iNm5s5SGX83H+USSGoG2A0hNOTw49pXq0Vtmwp/tM
vGlb7bEUw3bq2uhkcD4VlOI9Vfg3zmAaBNrIDv4fGEp3VULgVV0sJbU8ARAgmL7z
cStAbEREeJhwfI8ii1Etf9zKzH2TyaybIDYROWfyZ6vCTD4iBLG58WQ2lkFjEzVY
HB/ECAI0oX1hy8rOFmFAF+gCjuPcx4Uvi3CstFub3sm/sg5r1T0VxdAJmgSlfyf3
+2WQJR7u1IiG8S62HP+ctnyUXB9wk+4pZMR2qTQLIVdHgr0Bs5wewSyDeu/WlKZI
SrBsFGj5Mkye6l9E0yz02H3Bomz2tUIYpior7DEfqli3Ci3g4O9Fhx4Z5ckjNMX6
c5s86+2lbh+RgZEP2pgJu59ldgZxW2gYenfuELpa1Qxq7B4e53wvNu8sLf84fKD0
yj0zQVs+1DSBEKrAwrq3t4GwgWLedVPGSNuWowORmMbnKjWxiRElGQG+KtKkKc0v
pK7zOHXbg8UibZTxUOb/rjTDXsQCqv+AgQ6G8w6vcxrola6z0D92Il18DsOOm7rl
7q/x3jnpwBiIDoFGJwhm775v7+FiEkNYL1fdGotEFwL3BgPdkzraWAW1ZtQhA6n/
HKuwadJKXbwuwikqjQKeMnLA+o3DLJpcb6hUtU2p1p691Qc0LQAjtHS1fxO6HeO7
wl/2pj1JvZNgc2T0w997cwJ5d7opP98Gf9gO/VgmLdP/G5xP++LUI/C2OFUvUXSZ
nHcHuzvb3SVnata6WtnhHDZTH5GfEC4mcBU8bhRyNCFbtI9gHuKy2Rl7/gEZfYFU
ysPJ6nqGq7voFsOv8HU21uK1N+kLQ1QMKbxM8iTwun6Bu0YDoDkhsaiDV5huD4PX
Fxk5s0DikolbuNueJC39y2CFgBCpJe7hZgHIHnptuFAUcsecic/Iw7ksmBKiwJgC
gRebBATkRllxXRX8J08rSvvKQyJgWUuICYhybDOef8ckQMGdx2ion4vwrIEADxeB
9/QyVUUzts4wAahsobvSMS0EZzJzJ2pgk+ED+e6GY04avs6MbH0r/KnvGoSzVB/q
iPvoi6Xvsy2R2z+6cMCCfXq7ih/XixvCpNGaSkcCxr8KPna8EoejAG6RssI2Xxmj
DUI+YsgL8wbqxVVL8CwiWLpvdX3bnRmYrCGkKU0Dgosjq5fUuAJ/4CyDr0MXkH/S
YUOxfC2kI4I0xAPVWkMP1qqYQUNii6jDhoA2YAD7CV/68s7KyXJk4oGKNFva/W34
Lp96IQCXxKnYpIxsMazpGE+wfcressC962krvNB9w2wdjrLu9qfKGotDM/LDqGli
VMzy1z9Gy2N33pu6CgmaiDNFPPpQhqfnSA4WJxAf/uhudaO2bWvbKLajTrwIWqRB
pw1bgoq6XG7oUhTmNH2SEt1+k4vqumOUgC0l13v5G9cJw6qbzAa7CdnuT9apqLzL
9WRvr4VsthoVoyTTbfrOAOy7N4B0yr8oGXGeTQi7D/7NhTbNHNdSWxLDa3jwR0G6
AQ5kzjhoFWjeHHwuL3c08GRG6lN0ZCGVWaKeh4xVCbVFMUsjSykEcB8sqvRVMEda
WN+4KeWrfdAlw7W4aR7g5OYP7YoWZS5FCfakeortC9IocbXrw7w1qS6VtPj6fFMt
VRdZOiFtbzngJDgUP0yU3NfVxcqN0oacjCK/vhsM1ojHaceKQckwiacvXZnKCAK+
vG381/uT6ESk/Eb8ip8ln5hDY0NtgZStdYqQ7XhGWVSazXa+CvAnsRRF2VErOiKY
q0JFnrEkKep008Rw4unhwcXoTUyYJVCpt9G46b8Nl0clT8+O3TdTPoaDi7WlG6HV
EAETS2wyxwutdn6BDQxiJGuip77xLMEzcJ9TOPiSvT7n6ytxzXNpw6MHEM2LuglM
22fxZgy/e0yWVE/daLDwTtoL5yMAr5+bCU1WNW9Qje2ZvvWNbGt/N/qbQLn0bx/u
31H9YG1kUL1O8kQHyrDQ0rzZ6YAotWcnnKh/S7gIYpQn4kOjwEvnjeuTZAtwmQ6/
oQoFI3GUIKH4sxSV6ihBSLYaaTdtTjsKcPDJPWffpX26ARpjl/fsEp1pvOdq+1un
YFMiyKg71PpBO5R5VET74R0J+0KHtHVqEaiywNyE6EZxmeGzcx4wk7C255nTko1Y
aYTeNvhVgQ+WLopFONfEBA4KZYOpk4Ws+4Z3mMiuLGR47uUCb75MY9O/ZXJsKiBY
NmvRI7QVnNlI23qXSznscOyiQKz3c3xeqo8zIRuaSy/97Nbw2A9NXMq0EVq9LRJs
Ao9iCL8WwgilO9d2IPvb544FEARnBfRAdd2NA/aVYisH/6tO+/XN8B9ec/WLyFl0
IBgE87MAmgLqh4wX+gJU3jHtQzVEWAtBOlRN8Afha73b/+ZfZN6o/XttixE5GTN6
3Egs/Iv2mONXPujPE4WXidC6HV768T6a9zl95+s6GWCPYZ0/eA9rffyypRAnzmt+
f0nOBGEj8QnNWRIGHJFrTKuMv6sJTVBRYB9MTJEzf8VAoWcZ0upG30cPA+nIGeq9
CO28bdlGycfpwvNnvI/8S0eVQxAQGfJNkmnu2LGOe/OtV/PTCm6wl2wyG/2LH4L0
f/wt1LkN1/sDASpS9MgDabnfR/Osg+lOUhwQfDOKkCTUeW/4J+dLkDg4XuA5OBuz
M9jb3/rwUrdIGgMWgLTlZ4Z9Hq/90c71BkAOKnfmjRUzRy0HLQ65pmHmgpMUlTat
miEqtlwz6wCc/eRiqT/c/JUXXeWy4M8aRrbN7gbXqC14J2leKDehAhZ51gaZpdJt
+I9o0IHmdAbNV0r44OV567Y8WEN0HEG3l+tCKdcgnYDV1jzWcq6fCKvsRhRb+Pho
Hey/kHYTKZYXA8mHexl29VOlM/nutL0XGeYa8CmxNRQAaXNeVRYc3Q2IPedZcsQY
wXoG18n4/QCfqRrXaxJnmCrqUdRTdMkzbM9szPFn56zX7SmREKX/qAjXRGslJl2s
TE0Fu2Qql7UK3Nu6lNd9r5S9Db09BkOdgG2Ew0hnd4aWSPoNIkjDlU1FqhpDWxHF
ivcSwEKFlYMrWfQFQji9iD4F5sTteacyEi1iNuMaO42ezFwSJmSMbdt5HSOwEcT+
/Z2h/8Xw3emNoBC/bxIKeFa3paZtg3V9Q4B2paSJ1HtYc94IpnIEJl8pAshIDShf
W7ymBXJ66xM2XVAPq7RDee3WzUgpw1fmIsv9lhjfT0qpu0QYW36PG+kfa4+ybFKB
NZQUpRAnxpxor02wMKdiSWqOmdIBR8pGycyXfgGfWvzAIwNEUUEZMG3CsH0kmMEq
AY/Wt4CagWLNCCsTJxofG8lSFlgKTq7muA3ibyAuoJklspr+Fxul7S8UHatDhz3z
m9Mj6t9mnvlmqLEDdL95C5sBFV/HthmiHvAkgiPNbWGZqhqGzn8dSYV0V+7Jx47N
STxw5Wwr/kXiZWdaZRUVFpM8H2L0JHiIz9O3s+K8LfGlYunPXJPE4oFcHfid1waS
AAHF7pRWOeaFnFQuWQ2rOO9d8so3XdUwmYVibmGEjV18mdCe7Witn+Ym7IV0B4Xc
3vLkfyM+lnk40GhdY66UmaBzoiIj962DUgtWA6tLLigXgdjBC/xzjelKslYtGdH7
1Kq9GlNfAGFWPVIyT7uCEvAUZYraQuAAPa1PVAtBUBl6fZjlaPZX/RiZM6r599Mt
LkmK68ixgtqi3E5dzEA/1WnnamPlXoet+wk2iMPNcQ1BCAYCWZSob3pvUF4npw+k
hcR3XHrDvhvbs4zPwG6holH+5yQrAvmsiw+ELj5/qx4db90iMiBY5EtJ6huKwEFl
y2rlVj38X3GkPte7IXPMjKPT9KQ5fi4oaKM0QuSud//EGX1RT8fH4M64QKIXax7a
+RzMo4US5QJjBzQJ09aYGDiLyv7RIUjXRVEh7fpyzU6q71cXthPcfkbolDmbiP93
PndztYToE0mkImhA3f6z49YJqoNdetdiL+rFer3IPvMXQB99LP3ZIwCWEy8eReRa
ASkYjSaDBe6HN6gHiWODo8+CsATp8YQY7/p75VFMuBITucYXQ2fn2E30828yp/NH
vLQN4KGY6Eko6UQl7rV6S4TUfbAhTYfA9wmhh4AHzdJtKSS3uwCvtySEouLNQZoP
o7hGpjj7WoewSK5mLeEKUfBbJEE5Et3JRY5bJcR9sh6tZXI2iTZVNxKlszJP4dUT
QQY7WZiDo+vOvMpEqWrVkU0LSAJ5/fQjETBHvm2a1EgE7V0yGZN0OqaFXUIMRlw2
tPKIdeEVJWi5Ra3fDjjZ7/fXPOPKUZgGErvW+kOIelTEyYttb9J2epUCQydcC2TV
JA72JdH+ZV8XuOxdLN/0mkOrRjdjl+WkuRdh8SbmVuXVAnCU9qTGDP/Hhw8NK3ei
lExqBCBVnD9s2HoCDb7D/g==
`pragma protect end_protected
