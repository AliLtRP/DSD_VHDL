// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:04 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZCbpMgwZ1b/8W/pBlZqwkfj+KYGSVUHFXjbsfd6cngIKzrKKdUl25aL8AaZ1TCRq
+NKBXKhp2l7PiIYP7yOxE0aCR71FbMA2DxHy2hxUFCpoMRldiI7CMD0PYUXIER9z
T8t5OvuEWUi9eqHNx5CS5xAYpmPqSUERYfl8Q9f1qwM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13600)
7ryi0d9B6ePERKCypyoafxItTHgS48tpmZcJpD15m1dCAHVu7GwY8z39KUkoPJSx
VQjUN7rxbAw94VZ83rSCTuupc/w0RDehZPm5vES3vR2plPQGVtqIVv4xEC/CVvbP
PTf3k8+gL7QXYTQeVJ3s3Tqcwl3+MGvrbihzZ0iYwd9g6HzWjWgaZZZFjcHZ+2JG
ucvUuYrwaOxK9md7hlgHdPSDdXbn9ov6S9TZSn5iXUM0cM7wJQTXiCs07RyGQ3mB
a25T3CJNWwO4/PMtKNhxq53NzLe5cCdB4cUfH7deuEXDqKNzrAxwK87Vx8/f3YTg
4mpnMJo/QARSnep9aOAKHT2C1TvPxew+PmZQ7yJyrTsT9pSDJm3zRpFeJyJP7yJX
GnnZIc0T4iBstVOOJA/RLt0pAadDgWAagYfN4g6+m9I1vtqgLtWbzXynCnv6+Qyg
KgtO8VXbYDHdz2OTv0SH0MbrbT2hjzp9zlHsFXiKojGjxsFwv77DsviwPS58/BNN
tl9I9GVrd8ZDjw9DqtpY45+Dtm4OEA732oAdfsxBy1LNmLsDxg0Hf34die8f74UO
anrF9EFEr0CCCPpift/7PvqAi7OvrfYV4uD1xfMCkyDjwzDclEmmKH5nGkM8etNq
ePYaNWW0QJhSJNdIwVgUwuoD8WK95hsWqaFpnuNKN8vihWseBl1YiyFbeV98RXEs
kxPVAeTPLncyXeMiPcAZFxF6ao2LuIDk3kR6QxyqB9OVHpBZ0zACzg9qKjziZsEv
n1PXZ6s+ZBXyTnlqDI/sy/TFgHJeVewcAF1ILR5J+zPTjBZmXFysuUZj5ZV+CSiL
bX+cC/ZjjxTpRWEsSs6nSH/YkN0I2bvaYiIcawcxVpAtLAyqg0vzOSAt9EUjrPqI
+Z9Cq9CHYJ7MgefE3mv3wvrSsjTvApsQ/7oH5SxDDtm3zo5HJgFvqwxBg2LjJNZM
+dFooV4yXjxTV+GlauL1B46eYV02axhAPNTT2I16cvStGzKlovU136JTWR9QaGXI
qrt8pDjOlAHPrB0K8u0VgHHfWzbvrRk9cI2JeBox861uk3SKIxfYtm3ZsICabeUm
iSpY/HFSxR3FupHWFIzNtTRbf+/1KjnrALUcxjwWJgSyu+kKwz0+nIIoYa5reuAZ
qFFQRFfWWAyPyRwyhnpPq8XzypKrtjxgN0WOjL1eark6t13JGWNtZggYitKjgLNZ
mLves42KeLejueLaH3oe5Cfx4l7Um9nY7zRtEhBAQfn7SYMLekqsbc8/Sflgn81i
OeUyrbEud/jdeFbSZQiS46rRW5np3MOXTR+akJXbzcc/FNtLbfkJTUDnZ9OjrPfm
pB+216jALWGbiefPXxRoUMZFEWy5Jlk3OgQzx4ND+9Dbl5eLP8wB3gieKmoVBRic
MvmdSDqFSAJ+LBN3x3sgXjaVL4/uS1W1V4e8/ymFx2TBG5NCjz54yiS2nVYOuWe+
hY0BRHMBoqYIGUmLtreLWetK07hArQEaiT3agBinmY2zALfcw4AyDiTjMK8VYlVQ
iWVgWlw51jnzYo1HLXqozVGrz09a+4sFK5njc3us3urmCNThCcEnpBaZN+L0FPoG
YfF3LMn8NTtKxAi+sMfq3G2kxa7+Bz6UZqOZfN+2wT2eFU4aujsqpi2LDPShu/6+
BojV0IpuB2sjscRHqCdzUCvRAUp4sZt1yg8EiK6pVnhS18lxcUK5XU9WDm4kSQPt
k41xc7EWGTO8R9qghhjJyIsknXJkNa7spzrZh72kjjv81HuMz/Rg3tdQYV8FUCmy
ZErT1BuWE6X0XNSV2XFtVgUAinWBlvQEY+ZwPfYkaoLNXbltKmdm/PB54zKpV8Rh
v58kuDuLO5Q+UP6lioEe95/T27XAmkF9f1Z0ybxuPBT7j1oxgGr5fqBRk5zBjoTo
f/TjKU011ujzPQ2tRcVATZ8fpBh5aAkbwfD35w/oyq4Buyy6G2R+gLfqXEktN2Oi
K5NYVgVeymtGxgl0DmYFXI2MBjfu6WQS6jVWAMAWpwIfXszHuiCzW9yxks+AUnhY
fLAYF/6gbgTr99XmlhqIGdtnnyhwuNSOXay0cJLG6QddNQtGA2Q97azoltmpNhl0
dSqfpM7vM0+QzEgUN00RFs3yKzzYnBmV85/v+a9Dmf1MD00XHu7IhACno+BNa7uo
IxiRCmWZMP6SF0RbNJrQOgoMCFd0SG+yG1sUWYa4W2TdlzJg/XPNA/Upg5gXLSnp
pel/DCYmoHeaSx4eFxHTwCTT5qwzEpkA192KhQrkO8szWIRjo5opQMFa6mV92PWM
jkj1Ue8GeHlzvMyNKUQOU0jQQmZOCFsGxqWRMh1+7T4fG4BwPIxoidzMj/FACLa2
/1fOQsXXStFY7VvDtgN15xZl/V7BkU7SJ3Yt4y+pAnfMVBKCwz6vKeXzIKVs0wZE
VdzPXIJAV4931vj/R+dM7rxUetAnO/rmHF76utMAhiw0Ri0ALMdp5tnsEn1fi5q0
1rCZPHUZajFvhnMd5MGjvDJdYSO+V+pwTZi9+g4nrIB74VF4yjH3QtVVGy+1Px9r
AbL1Nau6wmqMsMZqJFiMTnW2bhzz8xGJTdL4/ZG2TS1LkiilUcT61l1an90Yt0Or
8oTbTmFg/vgSp8TN4pqtx+80tanG0lJFIlRqnF/kvexZANR189dJViKNraQoN4P+
ea2wWIpEroQ8HoP99yfaiQZZu0Wo5uYa8Xbk2s+DMUsf1eNKWvsgm3MQWTCWudDm
nowv6kwwFtFWWMfuVfEVL0d8mB96qacIt6kom/m35/k6SSCahsR+kjZBNlg2knQI
gdk9dgJp0+NgFJMYbonfkW39bgzgzv3TTTaYmQkmmOiMq0FtfUY16Tauh9Z/CHWU
f6GD8JqOwpQEfTuRb5GwtxS9fsfPVjn8wUveYfsE6/JQdjEKSwk7km7/2ONGiWZO
cEPScfpv4+HQV4ewjOi6F41vpXNZoTkC5DQXBlkKyguOZEVv4HY/6y28f6biyxoK
pIqKxw0ahcTxqY3fsqXTDORvYLp1tEfZ34bnk37/6/YFX05XqrbySWYlGlbrw+bD
7sFPZ9DNEDK/J8g65+zvLExop9GxuSUjUnRMERl2Ox4vkUCF2fWlDMCpSbE8iFSr
JBKV2YxmrSqhIZtJSZ4Y1DoDiGVkBERN26k1Mrl2SRH98fWhg5X5XTB/d5mflkFt
wDicyz41E2fmJbHmZKhSHeWGSzHtErca0w4/njzByU5rT7lNHgTVAq6WCxooZMtl
FwPwCD+/CLb/GSlWi0nreYeyfw/F2J36UDEAjIc4XvtFVA/Q8r46X0F1OoAJAz/v
kyOLlcvpqwz5ffHHr/SGxdcB4Rqu/ZtvG0sJUGkOax/mnpXM6RaHij+wqdckONrP
IyfMjWzZXO1CZ6V55KX7gYc4A6knindGXO4uW3EHf6Sc20g0A5eh240xWVLE0TP/
tVY5KZsRcLbG0sCOH7xgT0+Hr6pJjl5x8AAKVSCjpSpREGsQ9cCyoZSR5ta3Lcoq
cw7Rs7jYHP1vuzCZty8DN7XxKtKGGDz7tAK87sPdZvuvQbT+ZLOqJ/bM2yu6it4Y
3/ZRPPWEmn74gtcUBip2KmYRlAMijW2PpZfP3L+CUYXUvox38iQxFto49FCUFL3s
gV7I8hnQBx7fqnNiLr6CJALoOU+dN1V3LcSrC9Lfsl4xjwnFofaGfRafhjsJHtFs
eYxUCJIySbPDFysHmejrARL+wHb3OWSL7duqNNw4YMexBmhegjIi8FOgiiW9tfDC
nLcNdeRnhULs/VZUfpBHb3Yn38iskrVAJgcUEQXiSt+ExvzKS+4owLSwB8cPamtU
/W0PKaI54TZSfpzg6pZmgG2g5so9c5athQxxLRJnWlAD7mA237uTvkl+LAxc20B1
VkfmKJvWWlLk4rNi2MaZOcly4rjmDfsXlIUP2UCgVbjZLFAhO0r/Cvfpo4j28HoK
4MNsatBk7Pz/JABPtfuf2XmgTNfhfsAAxRb1oHKgdec5bApvZlpY5jRtYXnQ/qyg
tJk6yueFCSoxwxoj+ckXC50ncmkk9q+4bQaYEZdZ6hUB9E3HOiYsV7C3D6NitoIz
BgyCYX3OH3pghC2VGkpLQOJd6umub0gptrJ8UHzB7sBbL7Xh8BLrNgPv6MWHQZ0/
Gokh9Atsm9aoCpMipByqc6In01CsoMu0tisRFyUYOZqR8XwuNsw40LU3J3k6yjWS
2J1mpsTEChriQQkm6OqSqtGOSYN01kgMSHSPnOKjIEDm2QMZj9A5UW3bB9xrPBR8
7pTHoNM/fQZw+JUj0855MqNX0xJr3VVma90HXWJRrIVYT5Jpp2XW9hOXfDk28Gs/
ZRymz1eRIWZ6OZ5Vnisvplre2O+lONjJLXBnRWOIHhFHp1eTh6pUxbyVO2Pp87Hp
vqDMNac4xkOb+0nAOPC1eeGDuTAxttQs7WQns6OMZxn/x7UuizgyM6qBaWoudXw5
+HMN44CybAdWSyVq5TPvqeEIpoGRbAY9XvRtPnObj2E1Dia1vHUwG6iBhU3NCoSQ
lAkv73HzN++gQm7OOZjXEN1YqpLz0eTQM0it0NXmiX/Qg/vDaMlvqzOba3iwbf4S
OjZn89SYDpm5yMKfBtrkTVwFRuXLO4svoqTqo2i5PkKakwVfMT0RPfANg9ISx3jI
yBYm+gj64YtO6MunhFPrmzVvsUsEhdtkcYiZtkoOcH3K7Af7Fmv96dhlE3MC7Dws
4A7fc/8tqWx6o2ZrvGJIVEt+XsD/p4vM+MXUdPWvSoEtRiP24fZbm0eNCOZyGAyw
g5nMUuspQljD/AlZBWhQ8Dp4Qj+2EHGIM6t0YclBuPuoJyKMhoBOZfJ7VzSlERyq
Ri8Ubz7SBm/KAZfAx0vhHGCxr/MFbhYnWawplJc8FqHhAIb9ZjY/NxgQ21OgBXCa
tS+hXF4Axgv2fuiLAMUhksKj5CrH79U63kst6u7FTB9NB2vcKQj2KGAZPl11VQ/g
0v11zq8wc2WiYixvgQvbf2BzOuXsrReCsSnCFEPTB941UV5avKfyVUbMmrVObamB
DwLhw5G67GrS+mh/KJorKOt3DgzE8Ea6AMge0yiZ7GFstvEV+aFmoN5uVAQr+55I
0zLD6kWqD+kg2WSjxImvB7JyiJSx9EeS+H8ZP9i96vLXozddurU/uI6qhItnkUzT
CTl4QOwgPp0Gt5323fri3/ufq3gZMEY4gfjfK69N2cmJ+GmzIBzp46J+cP6PjeE6
X+2jCEr4/hnkHJx37nSqMSyUhgV7t8qv+WJ++cQKpK1HuX9zd3DgYWe6soR5gHq3
iea8dbkFQLg6obCnQjC/8dC25ApnohwVGM+LhvsgVptyXfsKHoyFZh5GnNkFkbpJ
cVKp+J6Yx4MlBYhNTM/1pRRe+13YEAo7+aQgk3eyCOLCO3nmBakr+pGoN3HsP4gD
HDBQ5iS0m2ssHPRAj12mpp0OSOvEkj5/deHEuAVVqC4Vg2Df3RGdIVpgfJHtJy8h
j/5zxXkm8OlslF+gGPSVDSk3piMy34VrccNcMB+7A8219j5FdT4lrtffg98MAfuu
vMmjdcttF6qKsC/kNDEs6mRwLw8KbmYxkzODppwD5dWMa7v1ypuYf7t7v11sA32J
ZkxYH7wC0ssXMGExRtUNcwJ0T2IOR4ZWqi1u0XHjeEzmUdfT/No4FLPgwZQyfCsq
oZo+AEZ2LgKKHJCzaSo0R2SL6bLNzQ5i2Vq4rIQpgrThIT9ThONAwFsxF5eCQcN4
E1x1AjWYt1rEA4V7L76IIrekK2pJNPuaaBreZg3C9DHeeaGFWz1l59oPUcvLP1tk
O7kWJqyeWgyyyvWZOwEdj1OiaTCAxWVKLIKburlT4mNwzX4kwlxzSLaLMB+LxKfT
xOCG8ZkA6s9Afmon1EHuVvred+p9Nl/7VpeZ7J3P/U5MGKoPIjgMJhiosO6Dfyi7
K6C0GpBG/1CCNU5MlcE2euX7pmLZON6+WZlCyF5YadVWeWgCVllwxHCh8dPDfa99
9/gn34qz+CjB2uGsop5UfEkff3l5Traa9rLZP/OWqmPBQEPy+6Rd184KnCdjdOx9
8vFcVSNCj5QcaQqsVxz/Dwqq6aRRR2ofPxyynO9WlARkXW6RPNOemaZvTkBdG+Hc
jdNMPuYrm/iis0/TWaF9wL8NEWL341OeUp4z8ngSR9PyRu+SfZn5n3zXuCtzvVsX
arIXy772B7KA+MreViVXCL1X0vuJGfc5YUdgYfqTNcT56ZRwV3JTMNPizjBnGOQw
p7nALEcODfyuAKeLzCZKg0aahM+bWNhI4I5n9W0vPXhHNLQMwjOm8ZvAq1nNpMf+
2t226JsY+9eO3YtE20frIQ2hQxFNlfif+QvuQTWX2B+kRfgKftaUV1hkvVwzAYw/
X+1SI7CCn1t9yGgUQ4SFhr2lQRCklXb+eIbTLPUT23QZPlRnFJJI+AA054KGhDB+
R9msdjE+IgWT1pl/MRLWvKybtrERnJBVVdxH6injXCU9YljobReDjLklNMBTTK7J
pIvFCJ1NrnmM/ujnK7VqK0yPDfJTrH6+LVbs0iVvJOwL1qpKI7thRu9IxHP9ZqgC
msIbaGuyDhQNPXGbjtHvnFkSqrebFwrvIubWw3zfSmpYSOz2qcqEnKBh/egIBDB9
/ta1xkN644v6YAjo62YSqWCD9t1MUFEHXW6ls+Dnt/CSU3zCQiKVFopsAuoWcF44
UIfq85d3Zw/dBHc3GEXcm3uFFfXIYR6kLLrVnL6j4FqQH9UZ9Dt7ibnca84tUM8T
lpvsnFYHF73CuJWBu0BqigPT3ggVQQkY8QEqCBm5pzsG4L6DEzcsN1bMvpChOUWI
EFo93fNA+PfzYnredrMrMCMX8q43WNPN/UVHQ6QSP4NvIUcjl8MdQnPr+KNIQdFl
4JmKkJJfrNQzqWg9vQRhGkZ7+45eQyefZjvpiwh/NGcCu+KPOjBe0qJDj4x5Cypn
JBi0JIVaXTJTtX9baHtv28NZ+Ig7W4CgCEQZhxfiURfFh1YAMOiCQuF4MihJOsXT
9D9tARWHkEKatMIfoPyr+b1mH/IU3bulvIfd2+MYNdWwW3tM1/DmfEs4lUYZffH+
Z++Q7R8e2b7ZITmxtUdfKeP9OPy8eRWKJ2riLR41nNRIRPVLAEdIk2qdDQz/Q95i
KwfxDGy5Hg8CdfkfgHraFqGye9OLVX6F1T7KJmAcZDR/qTjcw8A/sZtAfXXibmj5
7SgXJ1eh5d5TlTo9jkjDjVxKtAsRO5Eiz9LsRbUCS6ysKMKzUcGaVu6cTy5iLiGh
YYLdcbDPoYsc/8ktZvnWqwaDvmOi3jy8TT3sltypzRt+nTi4/fj3+CQrGldDwIwq
vcwj5luInUb6QMgeb2HaRVSOHLPvW/+xDOoL03H9ai3vyH+BpeKHQPAYCaJR6Orz
YOdMHJmypIu7FOWLwMs+p5FdzN6CPrznRdOR6a2VAtU2IgS9OA8bs6WRrRjbC1A/
HCF4PkBuIaaYauH4HKOLAjUrp1EUtq/0fwKgLXKDwpGu4r4Tnfx6MHiTiwbNQjjZ
n6TUl6RPwKTbcqbJ8H6174a9rHbrSvY1lbkzVZhm2dnMOc69GSnOS8oCpaiQp+yV
Ov/8m3lICbTuwqiG1v+ozolxTU0tKbVvf0nyzEHVA0AAMGmyrBQptGsJhdzkSqe8
XIWKa6JvvVlJB+UQMTq4AUzpz4AKovPWD943j1od3QQuZiXUzAifcEsdN+j3bywa
eMH3FM7xAK0A4tHOvRXt77t79kHcopQM50t2ID2dMSGsPcICCEv9bv47XZWRsuY0
qjGahXXW/KaQ+m0CL4SpGXRKhdI4yKNmdB0iH2FrCVzdABcJXABDaUGK8aIkSm9c
T7rcuKLxT1PxKbKcsTKQCrB3/3nq0KBTXgxDm6zu5mPV0TmZ51mwzc6sa52vNmO6
yB+UYKoUuOQFd0eMkK8qWyJvTpS8dlNZ9mO/x55ew+IkT0EEsbpC2UEhdRFi5aoj
tyyis+5baPYNrM/267pw5PkOCmqNI3OxahxQ4ZbZVElTXvgQHo7q+gt1jN04+iyg
fe+PL/GoxiqacTkSWBhzPU6g+VLexYUtOtOvYp1j7cEZ/iYV5KoJ0uN4WgFVvKdT
Kk6LrBy1igvsvIg0E0T86kIaznIw/PP3I/ygm9o8UYNVGISOUJa2HaT1kyj4dwX7
iVnF4fCzbEqt7pyvgFbVadxJtXKC2f+3EqyDICZ4cWa9MpdqgJaQpSAbzo6kQ7wM
zHefFuY2zeDbEM8WXlwjUK4lIJCvrL+SDJQ0Y9fR16cdSWOMBAJDOUCXJBQfqeeQ
1evJgsDZLcmrqVbgnj/j2bi859wgCY2qTP2CsXSazlATFCG/rBmNRNtozUe4N//F
TIdxUysQbKTEmalMpIM/QMxaC861Gc/YwBOn5hFACEthA5u9w6EdLOtOW5/yzRuB
LzFC51IMZ6/pWqtllirSUdGRrbHwiRDxyUittiRImiZLeWK/qIq/0WIgHscEFA+V
KkRscboBNShcpJd5qdIcsik1Xh8KlprN74YnwRli4tOhaep1PesnEVYf8GyyhTsi
8Kw8Z1uAoK6XT2KeYdNaj5aNhd52ZHCw8/2h6jKxX11MH1HUIvh5e9jO+CFN17m/
qX1P5nzAZXziavpNcCFXcY4nvWn/Xbb046im3lz2/8qYx6Ie8Hyuyc/klb/luo4r
0wgRC/B3r4iz3yKr+tR6n5SF0YjeJ+nmgJIuv3UTguU+fM8n+0U9agOvUxhrB4kD
m7/rf7N9waRhu3e0rUjAta4eVZU/ed9CILKCV4RZZpVEvlqdnTu2yaa6f0X3oUc6
USw8LfvSvbUPwtdztgu3REhrj6G+0JJU/b4t6LUw/VAylf/TBJ9Wwh/QlVcQr/D+
L2j+jm1kihhRmXOVkHPggRazU8NCH2wT7ck7tMEaHwQn3PNaIE6OoDWVYgo1fFlm
hJcwBl6ut+vLmtlfCiBV11iOLJvqvOA3bgaA2HPhHFPY3Pat+4qPfW/SK1QyVZl4
8cT2LwukCM3PpIArgPMIcOKcfFWUY3sqwNszgKuayQYXbEgT3LfDd08Et/LZ9S9P
SOrfZnTR2XctIwhX76/TdfI7rVXf9j8j0paHRaCxnDpqdyrkB5Qzggb9mCnaXcZd
3EDFxnncRO1Hj1VFpR0heNHzXypJT4WS1mKdNr09GmxK4ohy5Z0ubx/crNDxIAVr
Cs7qi7LhMBAEtKKSs4N+awneCq3BqcdezFLMM/F/3ADJNW+iohgfSZUGNFAA+uDS
E2dMv/gFkJ8Pz9mJ/S2W//CbhX8CSUhf3uYvuqT5VQIB/vH/LDaBmDSaUQkKO2i8
AFcKRecr+SAmtqoczY0htMsSciIo/hAdeE4zeYjGxlKtcAdZYmFtu8Bc1Xn6A7ee
+PSCi0lDR2szhU8+gU4QY2YTXlz/XyHlLQ2TAcbqs2DJ/3lq0O5jyZYJyQ8ELtVc
5oWHDQjJFwpV+Y9MHZXEQWRJQo2TgQEDqB60scHb+uj9Udoz1/+KA44VYING8AM4
nOfc/C/BCT+liggI9CgguIra9IGoUoF6oKPeGQG/XucLAlov0+mIc/QZQPvKA4nZ
2JF5rfR10x900i58FoG3JsZEVcH92zOEVYptAJnQW38nrx7medIt03CU0YvktmTW
tw4h9SWeOC+7jdYVwaqnnjKQ0K2a+DGhGG/54acSfU6sSd/4wHCq0Ee6JRP8oAA9
ysDj3ac4V/NZw7JXcXtcd41/zpjBPQWhkwKQdJd2T8LGviQY4yKAkGX0CwIrMVHQ
BIAHYjqjXsB1oKnVDv7zj3I+lEotTJx/8/wa0XCrToiuzSmPogz3TtWljAnwDez+
TVus3StKqWT0aRp3tbWYmVgWhsEiOGmLsrS5iSuXuhokxh/pSqY5ij5xFqyr0W63
H28S3KZxi3I8daKvk8M7oZxQ+3GuczXEEKZQVPQb5c5zGPMNuhTj5Bmy4cALweao
bZMqN1XB6kkuxbSeD31TxsT8WbtOX+k4ushN7dAQHdGu/DbhvrW02eQDsn0BBmKx
QKLGEmiU1BqdlgCwZ0l7A8vrRj/g9GnybsxGFWlQrNuviBnsrN+8ykuibJE7JKOK
a0EL7PP+0Vrh9oiB0S09lbPNqUuizmVF8YihTPHRbyQ5i6CL65ng06stDn42wCrG
Kq+phPjxZyi5UNh1yYfPuxcFWjIzMMbdpwqELMVVcZPp0ZJemuuwRNXf4lDohsZl
Ywf6nttgPFwSKzg5Y06aIcNtGXDeDf7bi0xMI8YJXb5rxQ9KDEw6iDQf1JXfXT4z
wcXmGMY1yK2RcPajl2h+Vq95CmM8N+IMQE18kQxNjbayFyfuAZQnnowFR4Sh+Hud
YoLkDOZLkJcLfCKGoPZ3qsvQfo5Re3OVqmbpctP30wCZm/BeKSLNdhKAy8IGhlL5
JKEtd/C3LW208g+imBhMtjuvIkWxQH0u5uzAhBIDt3qGkkKyrwdI7yIxyd/1EnpM
juMdJg0dOESsKz6j3tfoWNX3cGGipOD8MfUoDlWzZF49WheJPosPO8dwLa5eADy0
xxnMhB/KbQj1m3FplWaJme0964uev7bIrDnrE+RdcOxM7rd36uY21hTlIFayrcnT
5/9gEflNLTukZk8j4XteG0gh8c5h52VdKvnOOLUNu88Jz5+T/wahdQDBmtd9TSQM
dwbOxcWbCDIKtBJAHYA+GfrACpiNAun5d4uZDBBBBsyWR8XNFjhL6EyVKBBzitOu
OKe5fT0fZ9kHQ8+X0zn2SXxNgaooEFWmSYvsz83LrVNaGIhd/GPQUwifG0kQKJaO
4OZ/8Ucm9m6XHTeVTfrqw7OXDxsOU13Gb2qgoEAc8fj1CSQE5gylsXYi35PlZfin
1R75XGk4BbfZHeeSunPT0MPtnqPUWuA+s1R7Pzl1BbKee6+gRI+9SYdEdvlpaQ6P
Kx3MNHi6KL5VPbwqm80+s/DW0nZh1ntOXReUWPUVNo+n8ZKo6WiickWqCiHhqVr/
ATXggBsVJe20kxqHkG0Q8thZ6hWl28rPr4nGig8W0yKfs9pjKkQZoNIeSr6j52sl
KeNtKFd7z/9TUB7h8xlUXtMdl04/07dzDJUglBoTsnnU3sZ6rEzVNyb1+pyvc45E
8sRcbfQ7ZngfWUGYLTHQpOi98m0d9XHImUIlh1gxB0vpotqv8zHp6StiffH8KH+p
v7ZjMoqRkoB+DsaPZFMu95opWiv8Bmep6GRbIVCh8ruPf71dn74lPkgW4J8dXtOd
Ft/kdZb7fvv5Kf53hmpr8RWUl1RHQhC16oZXcG/wyI5xZBZJTtWnsMX+W9E5v9Gh
fhlMlQ9wy3YLsfPT+cR+zyDcDlgoZ91Ckmg74ZoGAtrAgbGoVeAq2FbSC7NFVLbN
SIyjsu0Nk+xKhkXTn3Lmstz4KrBbuGu6kIPGsB+krYNK1qg5HWd1MrNuTYhCtzIK
8RTvdbVwTpMbQXtGfQXR0oiyJImECrJPZNrSxYL2x8m3CokmS/3Aip5nLIRuKq0n
l0CM0gtr3cvC8+PK/8P0F5sGOa6QAPXITPWQ/KkmvMEtFT6MpnK1xrNLK4tugGiF
jtmKp9s97RZ1Ib436UHOMnPiWmuu45lh9IMWM4GBKRqEoaTFkVNDWPIyV69FYEZa
CMqeT0H3OFySE97GR+NUAroWSNFBEYHjd3aMUepNupU3tM3VoA+EHfnzDvX38rzY
IneXt9GEAvtSEbH3rtkW10d6rvinw1XrFjYSGf14YR9bACh7RrlLQ9TFAa4dfHo3
i/30oHWUMpuLd440iyWDmbLL/nTNPnIF9zxmUGqlOXTGfwY4ZygIRs7vW4kaTOnt
pMeF3nszduE18UsJXNObn1TvBaH4nG4D+B+k0gQDDyzwOETI2g8Llqp8PnRA0IOt
rLcGopmQ3IFB78sc2letfh8lrYn+DWoYhp6NvJLcpKgJitn9xrHNB/Ou75NOkWAU
u/MkDkddbMlg6Jcbr0Es/2tdNNa2YGqzNxxLodHYlg4e6HvUMF4XNoGfQTbkRWWT
opw9o5YAAT1LRqxkx1pz+xQuXBbQXUEJzNHjO/MFaDpEca4IZTP+nOIdOct+XjtO
yWvT0iQLZx+uAmosL1RLFLn9xv+ExgTKHiGHxjY3QGdAcnW523w86Xo4TFNkdwL3
ZSgkxy8N4Qqk5WRpqN1uUno857r9gQ6+WFEKHtAqRYiZjb8GsJabgqsOf4CLroYh
QyOlQRX7nbdw48sR3803siYaxBRj/d5klIEwgpyFijobfKalWl2RBfU3wm1wGr4k
Z0E1fjiQ6mcY5L1Cs7Py359wfyl3YX1/G9shaZd4ZzAAeBme35i2+t9AmbQdnp1q
Dd/lAsdnS6QvGn3jbJn9M4Q5aisDcJtrCPAc8aHynInfgRImqX53VBJY76C/6Q+I
SPB/fz+RGO/6OESPU8zNbjMco4HJHOAeQQ8ejL7NReyPNxKxkM3S3pWy+lk5r9w5
htpCIXx1Hv4Hk+T2a1AwrZBLfT5HMFE8CCvd86WGJY4M21LU7VVjpe4HxDN6u24U
OJwFFvqD5XKL4oqsGBsIo+XZJPFvNy1xRBvbod1aLGxCOM9Dx4TFObVBxxfx5fcP
NatlhapItlhQmzVISiJ3Pd8Egow94sM8GUOHFKjifax3ibAmQY/2NlpO1nM37woV
YhuGWi49dY7cGVumyqUfMdMk6rnPqCInF47AANeceuUdrWppk7W0vxe9FagWKRw9
I+dnMnxL5WqeNGk07J2QgTLrGdTrxcc54QnuJZDr14KqbaXjFDr6GkUEVrzZBc7I
4ERhg7PQX3hAc0VuDoUtH716Oaf68iwA6Yt7J39+ogwPUlbc/PF4R09Qg50BEym+
mWWdKUZ45sX4mgbiUIzWHYiMhEmuNJ6P7+RBlzTyBVDXD0KjLctfkQP+Ut0O5YSe
YYCmslhdbW/6GjAsZowMH3Iwr4+Uf5G1AdDPPDvVsV+aWrgWhpjE0qUdq50+C3PI
i5IucaXhPTVeHCCwEI0puxOqAbgTGrZR3w/a1Bwm42Sp4bxXY7t+tHHVNgV/bYr6
wZL3tYkTI1w/xAPuf8UwM6lrcwwNurJVfJvw0s6m9eYU9ovwX5Q5Pap04bwwYjw6
Q9+9ADt89RWedZc9lXUHkZH1I+ICXLWzC/9oVVF8b2Fpq9M/lEkbM9Ff1RiqweC8
g1qY+NPblCHr82WH6/uJrDwJP0Qj99Q50DjgKXIgNXFOOxvD7bxkaa9YRYWo96Ma
2tvZT9iU8r+VKWbsfOemMQtBFu8GhOzIO0j+9ajmZzPTkPB5CuaMaY5Tyi7uuSAR
CSv4ZbkhluR9/c4DlcO3xEe1A38xEMRJSNzo9cXv9Gf8cMjBsCEgvmJXb09pSE1e
ZHjhiY9NKVKg8wVTAR69nY6P3p4I9b/YVr70+RWQsz2UAOyrT55+0cF63AyXTpME
P9Gu38hNR0CrfAfySZ2JqWmfzhwULl0f/tItOjPlG0uABsV5QpMHr0b1qE6i1k5C
U+Kvk2JLsFX7rK+EXI3D9Z/FJbuVffjpLYiyhOVmlah3/XApUVFTX7lnxe2huuVK
2XwPLt3C+JALZ2Czw3P+MYYB5OXKg+uIq/S1cfo+wY3wTigPY8G2MoWg0enApS/z
2xUN80MNY1IJ6xUKOIOHR4Md+NV9wfYtT8FCca+LAhwpdix5NTYByLJO5pKh8JuW
kaDy2QWvXfjfGLWzP+hIRss8vz+ksoCyXsjVM4m9GcHro/pFuc+PvM1svbUrmRKo
O2StQDK7Sa4+Mx6Wt9WnnJUCwvsZ04QO17Jmk4P67HaN478EpB7VS/tX4TewmT8g
XM5WPkl5rldwOIeLdqJLRJ/qmPOXzFHcMamy7uTV7rXkwGT0eEQiLE9FyPkf/dJM
5xlnByPdWhgHcOIvNs3XteB5Ul56SwzwcsmQ0CUDbHWiE1RkFrD0P20DzxLcqwI3
8NUQUKTQt9bCaVDShnGeefyBfZTNOU3cOqrxr8J7bGBzjjWVJMlXAoab3zJRqcLY
aBGc1TOgpQxppmbehec2rT4eqUqNrna8XaYMh5lsgqGLUTrDhjrYQ985NH+2ITYR
TaouWtUa0S8YdAvtRtqSjX6gKamynPRQ5THcFZuFQV57yCLDmpc0Bd1d9USXMLmT
w3I+df1GCUY9t18SOT70IpEJpZNdlBXRJBSu+qri5VUauLLaUbgPXJhJeW6c66CP
a47iVJ7yZlvEYBCAqzGg9On9/hANKW8rYv9SHINdKjFgtcre0sAFXwnxpt0wXUUG
1EtN/jS0sJQYkS6Or7Dyi1Ydr2+ZvKvQhKET3omjnGWdy3qM1ujBD0ieW7AheUPg
Jckm4es4jMqe3yjTjxitqwOS+jjVEpGutSx/flAjRbeS2xy3LrZznpcgFYypxNCF
KMRGndYz8UKo+rTlMn5sftHvPZ6Z/wAqXUQ1g8Qag8JPazh6Saxn5DBpmc6Ja3EW
EO08NcdbOFXazTpP5+bxwaqqd4+cFzpEXfu5FI+fK4D/ePpVf8iaon0g6h9MMNgw
hO1Rd1y2FrQVIdo8RWV19V6RD2PWf3xcVSix9jBiNEkyVrVnRf3kA3bSkIjEIXDk
KpnbhIcnp+WPhInKiBS5XTxMnkfTJSjhmIwoFt83I1139532SbMd3JDV5kXN4jiJ
Qy/dSjOTvgjYhBXmdINHwQ2UB+UnLrq0p+wwGp82njDVq55hLmasxT/pcOenqOJA
42mqZNXuPSl5+AknxLI9wPjLDlL9i0tSvnfnuxpzGU81IdDeKqoFc1p+JP8Nib6B
7pFNVntLbcLf+bHxA36m01aqSTZ+B0XKEltDsFxHQCKH7NkrdOF5wD7xAhV2YblS
q6ab2B3r9QGFxqVs2hzdv1LGJxFUBwtQkDF4N2GZ/Je1lEQkmRm24gKSyBjOb3wT
3Vmeik7CpOQPvrA1IPypp5AlotmG6m4l6/ZA+O/MSXt+wJq21yVKfVebLYtS/le4
lI4WCTHKfiDYm7Tv2q6yHLVPCZ6vM3TlUqo//Bq3jKYC33heR8t2FOyXG0s0WdA+
EDswgzxa+kPi2Abm35MWxBjjTPlxHiTi8+nMnbjqmys9Cf8ZjGIjuglHYPlDAr/G
0xyaqDT5J/knQy1//vYJcM2XlKXkPLk5rkw0YvcIH8jopgMe4Fnze5PabmF0+Zx1
0u5dYIF9nwf8LP13xfqKos7M9+PKBpgkUJto8V2TO/EVbN29a43RpsKFQeVuXXQX
N6RDxMmOEYBTWGdsjKupTS8QEtXrLmuQtONMSOuu4VqBaU0UO0QFzDxOjb1JdBfO
zTjPGsEYf6qM/tFUNU5NtNWXQp5nNGYNiXZicUddFf3J5qK1qWiP2Uz12AH9t1Zq
fnm2cO1Ot2noEnF6Cxxywch1N0HvI8fi8V8OEz9kQqiF5u5HyBp9xf7HDhbPSil2
Qx8PRR838w/xhu/381nDscHQ9ibQct57cosM3X+hxMMCDJirOaCNXlspboo9OvHZ
hs4Ne+2AhFAgVEwTGMF8RwlOJyfY/p4ObWvVc89yzZG2iZC0FKVyp8iUBYq06U4a
m0NP33kf758UkgnQWWesyF09NITsBvdz8NVjcWrZvqPCTbWMYGapSgYME08qDU9O
8NrZtPASwK9ys7GXi6kShatsjqnwSJ4SmjOhZwYfWiYJ6+oLqMEa8/chx2Uh+Zgy
ON8DK6fBJST3GNs+Zy6Li46rzvld5fOO3SF1KzUgI16X9q/8L8930F8hqfYlbixv
Jgdgq5z5YZA3wRdyjfaHmgJhARhkntoQfvEsSkzmV5/JE+C0+us930GXYnSi49Z6
EgFiFJ6vHu5mrae1rgpjcyCPS2rExotot24H3L4dW0c+C3RSo41la/GTWFeClqt/
hC2IbSegZMX6yIc2cAOs6zYJjuhFO5h4i8lwtf/dB3KXtVaxTRITSEC/yv86g6dh
g/uayxsx3l3hqCe8Fer/wFjHHbfy3LmZdnPCjNDN/UjG1tAYN4tBz6ew8jHZTHu7
spDS4L6IptDVSx1kPLYSn7VS+Fw1TbFuh3ymX+Sw0XoaH4TpWOeJpXxu44RbCO1u
405wj7kHLperArrrlTvB927YxA7EVBnC0xUnsTvczqVrEqLS/NnJsAnhU8GcqWIO
XtjCw/+hQ8a7v7OkcJviw+XpkidGvEhOyMBNy35iiKgMz2VzfkBx3Lj2QhxkszkT
hJhq/dAkUoD2klJyv0RiIMGYhSwq18ERVcxMtnNoDwCmn+u27ESB6uviszBLbMIx
GHl2CoOrCSMQ7fyN2a/cu35AkG0MpdXjKyL1Y6vYband7ZIdC9znzk4O2In/+Kyc
Y+cXYodSg8nJ0Ev9N3lBlVRmhAH/Gjj7HkXn+wYSz3KcJte3pWyEpBAwKPRlb4u+
LmenSUUTUrbsk6nzvFv94MRwztngDqg3ilyV2nqDuGGFhL49yFR8/PgN//z46vqs
ptiz8g+GjNih6XhYaARvSkYIZgzT0x9jvzF0lWjzrakzS/zO09m0LeC03IN6P/8w
r+maXc2VnX3QlssYeCbWDB7XWqMdX26BX85cPwnLqqd5ghKZxZym11/lLPlBXox3
qum0QhI+YRlf6NmZz4zEZSKSYSAdspXCBRfzI/hw6Hl988oM2vzLWgkJceAbt6X/
Dy8nvQIp2cMdAHUmX1Dx1TvhC82y+sNJhyIXJlkm0VzfGTxMMdklNQX7V6DOS1wy
0Gfizj3HKSimy7L1qsOATXvxBzB5bmyWRRodEha05lbLoz1IQLvEB2/7CG0a+nt0
s0qybareFN5qxpRgp/iq3SNLrSb4c55PxfmQ61qSHTpv1zoXQsGc/PRh+Sm/mWAp
igQgNi3Xtn3YiPdkFXOe/rFCRJzYi3GyW5uzSndL7Mp8KvgpAtz7uzTOUVOvXub7
pVSzlA120p5TEGfAb8Nh94ycftGUEpCP4udm9cg6dI7bLTrYyKwr1NtNiMHzJZNf
3VHICdmij/1ZxFXoHaFG1u5m4glwd3fnSDmD0FsBAG9XObUMvPvYXTKseJVlioSQ
wXNro6QQa2XhwQinurBr0qegntRi97W5Ld/B5lJUcF+KSSZq33SO54KI8lSzcMHH
Yoq8Nd22HyndzGq3zv/HTQsPOHOgJJk0jI6TS457725X7NRsVjbNsYeqfQfezukX
L9+wdbpTxRLSfhxl6wHhiHoEdQciDTlmQB8TXk/Fc/sCJ5V4vn4GV6v10VbODUde
5PXhsZq9MKFsqgRGAXLwuAoyVLlmU96rob8948CaxALBbbmK1EXZE67VdRiNfyC1
bTfx/dnKr5BuNUT65L+CoFQ8E+QFrgx30T23jGPKVcJutKUWpGFnAcBMJDfdOGuY
zrQpdSPf4pcAXU9g1CU+RwYe7hpjVCOhGto8ESUfeP2qydad8vV096fknsNvd1Ju
cj6p/q9tI+rgsG2mGu1hPNMyCiBc1+KDWTFo9JmsAoOri2seY737ZyTAooxLCJd+
C0unSoDrUo2fM3hjFgZwHnfyHQwym6bIs0G7A5UEM2mkcMu11Z3608xc79t0F4mV
aj69WDy5N0RMDhbIhCpf7r02G8I7PwlVDCsOQDG3C8J3b+dKkvwq3waG99FAL0GB
t3apnByjU0J7IeSzanEC8mQEpxKhVu89zEJCv5DzvGmXYMWaiC0TT3QwQ/+/bY1o
BGjOUglK0bzEWrAVu1Jj2aKMVB4VrjgofHCr2ocHPYBG954SYQvlQFsokjXIPOcM
lF7z1EWbx/dKzpCXDzsbUYGd2IVkmg1GcmLbCEBt1hzmcxS0rN91Gl8x8/PYqCJv
QCv+bcKaxIBkwriWx4Eie3bIUDr4k+lTrQuPekTwFhVTgIw6IyQh89/aDxLjls/t
iJ23j/yX+Rn+y0Id2iAoIk/MPxogULXfirvUQGC/9X3WGFxOFujxrAc+HHIQErwA
Sd17yT/p6dLySy1ofNAy00SLbr5Y1dj5rjUqSbvLZuKI5eGnysDPW33f3cIpKxFE
J3wGhibUJV5OD74EKhlsem5rPWhsa7IRkSwwTkkh+t/mrK4MSPoVRGn976oJCT2A
xvdnYzvO1mJMS9RBJ681nlIx3fWre6iMKvhgt2Fl+VjmlI9H4iEvdquWBJiaqs7o
6TpdG7FhpHoQqK5iBDCO0Q==
`pragma protect end_protected
