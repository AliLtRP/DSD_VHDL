// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:46 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
j3HjDp/I51dXRxUCL2We4jBBCYIpxE3RD8ZqRGfKZsZaAbIJmIebGkKiexqOL1Tc
V3FaIz28jYN16EQ8ZyTLWJ+MMn7ChfhjVttpyL60zu5SOTbleB70NG1XJMET/eH2
90WNgxTgVRetuLqaTDHZDBybJN42aECyKgWQgb709vw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 43168)
xPHVjMwtK08TKlGhvydVrr/DnQQRDL40Gd0610RhJidhjzfiJalDvKok+7dzib6b
n2c1gy5RYQrd37Hwdfve8tK6od0JVjD4kTNz2BdaBAy61G1ENEVaTDTDBsRJ7v3H
JVP1gmXC4g8T1mnUPlxZldfzt99LFQD/dA9MkWdyfhQXB7BsMmS6NWIq3Rinccb4
N/aobgCYm9QVYfGGFzGxfhYibYACwU76iT5mKi5mFjWuMJuiv/hpui/9vpuqe7IG
X1zEKW0Al4/+Y28C1X8dA3OCD8KhMa9qe9ybaIZf+xxB/A1Lyx/qK22W9prbw8D1
SYBiF9uNwBa2dy7/5QK4j7INMlJ7nAPDZ2NisDuLeacxiEqpIqaWUHs5RID99e/M
2sE+V6ENK/8b5g0uMgfR6LH0wSlpUYAFFu6GMfxuOZHR7QtYY1lcPFhfZxqaj/xK
LLJWs3nTJCEFcIdZYgyvWUpVLI+0H7BKSc73CZFJLxf7yw70cM5fVHECeTD6Vvsi
M11FByuNymyt5JurGecyvsoxQOh8Gh+sHiRIp7EhK0pbLs/WxLKUF/D3ljkMqiv/
T5rvMgMA7FFV1C0gKpeu0pf4I4ti65yMbd4uGw6yN6IPSI3EYsGn1871rnmdr1Yh
v8Rmk71plQZ135bDuShebVRrKos8sdUzRd6IvJecKmDn6PZnDBkfyq0irG+UctTY
igyu/wwB1h5P3l7wyKSIepjQuQ+ewfT1EBcAQc4w7fFsNpWiYwgfVSn31wHjQRHd
PYzHSHMH1E/BdSayIjV5ADF8elatD3Jugts2F2FcrL72jjJBG2l99r+BT2XsKxrq
HJmvTdnvSArsGQPbTb9mpHoJPhsnMGjtXEYwoxOx0W07oDSyo+czejDAvSGaLLpd
1EEw6ZBCNQb1nwRpV0nfi1Bja5GhkEPGqwfW1ljGfOvZD0Cn6gc5PwOSPrG1mtJJ
DOzV1DU0FDubeVEfuFq1YZoGLGmyVxHRIGn76hKm4yWEGAEso5nrvhBktiEKxcbz
kiRtGWko1ph7TfyBpKqHLN1vGvxB51Zb3PDMGEFjpAj7pR63KIS5Wgb9UVa5Peoz
5zLUdIoQOXY31YryjaQLkD2z2tALlLMCWtPtWu33cN0Aw3XmAe8pk85ez8V47gj3
1sY6Q6plc8gcX+6y8yVsWBonAxheOj95NajI2uWdo8Izrr6kEtiAcUXtiANz11oJ
YT3XtN9RpLLlPHaI8/YxrhpqaHZLDaLozi5498zNCV1vJwPewnsluzY6eRsRgek6
ka+aEUe2g1X/jRr5jnDYXAz/U41889FBq0RHvIfbg3Q+VVaQgZQjgtctL5GpEg4Q
x73cTrWlqCy3LlxmvpVEHlI17CRzEmEMpwMOHb1OdKFIY1bEbnsH17+yn9bDzHnq
CIdqQ3IkY2Kve1S9FTp44ssJ3dSpdUOdZjLK/peIRCRbkCl/UmrL/qDodphEh4cp
jvLE2V9INT+BEiVj8SfXjcwZK40yxMbx8+7AdKRB18VUJaiYaks2IFiINzWkugDQ
Yv9dHHWSq9rYxfi52s3Sewg8Ull0eFWXF5MRokVUkWpnUxgTMdW4GGP2LUKsCKhE
gL2ommShYw+Kfx3buI+IMWqtBnDBvOGNQjN4rT4zIkJhbGOfcD3SdxENE07vQbbB
0VdcqIGbY+y3tWSKDwK2Ux9NFL/WCMs0MdQ/j40xKgIrztsS0pGB7csJxXzoteaT
wLmxHdh2Crt4sPcMFtULBnagvjoVGVFjIt88o79iK7zvmEyKXQGfb3Y26qUcjLR3
Hf84qvgGlMNlOtX7z6lg2uzHmvoq12Tmf2U1qekEKcO7FTm+9D7PSHrtkGrt16aS
DHmx92UsGVBHZl31aiK3uUfFqOSg+AWRGphC3ZiGxNvORQz8S9tdWnncpMnlJUa7
X3qM9UW2VlljiZXfB2mPnayY0lvKhOqCk9WCQs0cnZZ5pvCBt86vFuItK7ittb7y
IM9O0RYvhy8375ddafqQxYmshSfTrdcKzfRtmxoeir/hMt+H6lokopREdcYYoUwr
yPAtd178BKFWboZL5PY3oBQMDohDnNHgiGBKYEU+desjeot5YQBpH4NiFAVEoPyh
8YoYnIiKqZo+pc9F/0W5bYgZNe13K71l6DGGIbLAsN5DklGv8s1XPT+AK+WxUlVG
28bQbQIl6uK70CMaVtgjPncF+ZvUnLIQT+jhS1AyALAWGQXWYvzpBtNgVCeAFcJ9
zIvn+1fy8k4pBxYklzSXnKVDh6vnLil+kqPDUmJg94hO3nSwZqZAWuG8+X+riP2d
fcibopETSxflETHz5GJSkEaecY6dmifXkDk/OG7WPw8gdSE4rYJ4GcCGXJbzN17d
pypf+HBBHRaZf9/TSDLjokOxthMJGnz2VOfJypPvCifRu4XY4Cm6xZXnbq4EVZzc
IsmpaPvF2JIkWnxRdt7YT3nU3kB4sUv2aEc2DkchQUYfpWj8hDlMvCKfYGMdoTSg
TU9XaJKY27nEISNjTPjuQgpXxPsGni25VmVoNPwoKlDNEWaomnzCpkevs/HDkPyJ
J49FyGhqC0HrHN7+lSnHUop9FXlMkgA+dClcEN7GZig83841eTPjQ1hA+o/5R+kT
XTveBoFcABYx+7vH21JSlMXALolT5DmhviPuQHdlpy95RTMggcqpZxpkUOjYnqmA
d6xB6OQwDqeuiYJUvliuFfczJwSxcSHir3zsspB95uqymzLpOvKi8/Nw2wAUeVgM
swX4VzubFXvpVLQzNhZjeRntbwTAJnoCwsCMhTslg9/7uJYq+aQ+IFr41kjvacY7
xZbP9WuAmVPSuJzGgCRo1lp+1VpgV4kx6aJF66Zu4qBIVcHtNEzhrV7SefsYqfaQ
GgTXby/SLg72VhHDnIB9wed5lyF3Q+xhcndfoJxh2fmwKPLih+LqznZLuJRP6sJq
CioPwAblMjD7/Thf1G2OIQ2UTP7mltf3ArEU3Ek1RR7vOoy7RFkuymwsdYku3myD
10Ib2RXQxnNbmssCicTbd4TpWxzzOaOpedIBCHZl+OCD0D1Tvk//RFzaFK5oJsPr
QUVT9rQ3jwTZjG+5cy6K32Z4aJWV9/bHJmwF8+8ZQSCqQxk2e22qqerWl/uS3UsO
qyc5dtXlVbejzwm6niBdPvDx7u1Kr4kbfJGb+Nxeihbz7HOr29SkOwZIY/cglSn3
Qfa6DVQ86i07FZZhjoNOYAjxdgBu1jEFVAuWpsIBg2TXaOpV/bE1ZfVoMg46A5YG
brWiLMaK1Lexn6ExyormpRd8xaV3kQkMlRmsTHpOlM07/xudwyiT5/zPa8nh/nLC
fHLEh75vQnQk/qgc8pdiLcdOdY9mQGHuR6Gk+WgHMU7lHyL0W3XE+w4RyK+SET7V
pLk2ch8xhdO6PD8/LJWvUSTfrI48cps8zY7wRQ6Um/FjDJyGul8NJKDovDkoVIul
r27+4aewQkXJi/WgKcQ9fcEHfz9bL7mhc08Y1di9VVKGm1D9bj68r5T0GATobMhw
jOixhc5ORfq1upO53XWPJRDM9lZAgwqKqe0Vn/K4+qdCM0w//6axXFoAQw7n2BxY
ua5dGClv24/IIzQBktBffWkz3F8yYX2kQyBLaE3De2SZnU6ecfTN0jWqNWk8scQp
SO0UR65ppKhyln9K8Rca6MXjBngtMZjXhjlvmnwbYsmb5712aJrs7udaT8vxrNrU
Rxi0G8BC7Ou+ryb+LZneoXoyxumPxWkfoCqhHqezqX90bnRAUNNHUY1RK66aWau+
07k9NffhbdgZVI6LpOJgzSK57bM6j/WWTqA680Ma2FNd9ce2lAK+iFapvoJI4Cir
9n4vM8gmxncnCHeU7tIpHhKwD2LzIgWJ6vPFoOOgPWnP2CSdl4PnHpWxJF7v47Aq
btcQDFOUjmvudynLhn1lw44IJsxEMq8Fcewi2uSlcL+pFTUhy+xnOmLZDaxVShdU
uc/BO0WuAdS6J8+2oCci6sbk6JKdk4VrlOtdGvliHm2yKtyEYLroGN2hR4EVE0pm
cMlhabChFUQ+s8q+hhSi2gUIrE5n3AC8f/ZLlh1eFeGThYYJ6I/2Fl23sR6asDrA
4rGUhUazfhiCVi97FC3ht0ac9cSEU5nAxCdg+kPUW9jYDopHzeCnk/x/O+ucs3H2
/CzTQhI8liPbQFq/aylOY9s31rIfmssQu4wd+o3j1QflFZu15+vBu7E6Z9+9+qnv
YQbkQNaoprmzbwj9kmKaNg7X5/LGIfEppiyIhLaFjfhSeQ6vum4epCS0XLov75eQ
fC4xz6ZDqJMnRbt/ruOF8QRhjNKXPhHpL+zab+GkExRY1Mbnvw2HK7/Ix3dU/OC0
fFrD/YheD9Jfoq0cEsK/oWigj72CS4plL14SHoXChyWDfAyNYJ8OWAUE0vf58AHR
Qx9bup9jSBv2i69GfZorWWh/6i8POt6xpIDpLO/JLp2xnlV9nXb04qdD1c6WAdlR
9gvdkdf11wQLf4gw6M2S7CfwCV2eaA2HALrjrbNw0f8ofQEhO/EybPDSgoJVGbag
rtfa9m23PPFee0I0FI9a8B2gKZiNCaATKTxSwobqyAgH7zEDR7bXSVPOSfUNNk1y
MMQ72BnthvVzO72oUtsNql7r5stQVxEId+Mio3RNEyfkYSpG69sFiwccA+C918RB
VlpU9Q9LHU4ddmcQRXWN8azNt7C0XcHCLEgYP/KIT9SoErfQWvTnhrh/WXoWXvsG
5jkXbBLUKgBf5wh1eMQSr322fuIfmER8UReV2qrxVi+P4FahZYSDmtRdL37hu157
eKyDR6l/DDFmsjx4zM+s96/3LDMYy4lYEfXbq28tpK8+VHDdvu4qOLpVC9Yz2Uow
WGdfOylaKyXlNGVCrW5fR0g+9dZYLs2T9TV0+MaMVrrWtMYm52JdC8ZYPqXsgVjr
GLRSXlq7cghIssQQeRWzWGg3RpWe5t/ToZ38Juc+1i2O4LdUA14ETDcP2Envi9+K
El1b2X8ePCAFrFsMAFjOyZ2Zwjxg/Rsu7rReyJD/lKznsNwnAlwlzzhm1l2s7osa
Zvtbiahm+uoGU2yCydhG364MMo+KMSSN20eNNQTvscpGBVwPTHtkxRquyqbPosS/
NENC26H+RsYBd8JrJnJ3TiLdxn0XSHKmkQA0OayBqhzRaZ132WeDY+j6L2AqGIsz
wMQa0wwwDRtIb4LBL8FHLGJayN1IYXMBwl5yHbf/23PbbKYaxphEsFNr3HLwNTVG
uG5XammNOP8U6x6ygthQdFnZCCBJahnIoGzPIgvK/Q/r+BFuPLCTYOm5Kj61TdyX
VIO/8y+IqteVjeRYad8IwiR8hDJKYgaBItukgd3ZISLoRlXsXLw7JcDOiTrUesGr
Vw9YadUy3GmfSgb98OcTbmv49ogWXPuCAaIXQG/OYHW8drqw4RWF9XqdztLXxznT
yGO8DGVVdJYXCIyiobCWE0gnHCp4CM7Pnl8td0CDeb7kh4DPq7d+WbKactvdjm2Z
2m/kZ6/DUdy2IHMg4oG1+82MsPVW7ndMFkvP0ap/aJJRazUoBe+VQBOEwFwHM7Lw
o1g8g9vlU6SfPZC5tnUPycnibotzKKsEXEW7Y/O51FZsihcTjZKmh79ldksmSYSj
gflH+D+5KODHzHO+8dtDfUs3uMFB8gHJuaoAU8oluH5zDwAgbQnGA+/uhhwGB7SS
7sU9B86V2S0Kmo7FR7t7K/g5tQlkv5K6GvZu7OuaLWg9kKLqqJjSqRisvqVj9DWQ
5MC3xCb767AEGOOfFNC+muJFlQm4zbDazJ2t5sD0qJ073zT4D73+O28Ta+YNi11G
Mi0Mp01s19TC+sWAmOZC4iGRy0mslrFnIvYToRSP8vaeZgy5TdEMLOhYH3tuSuZr
XYJUO4es+ojV1gIrCyScCbetXoommNrtQLzEFA+t288j+jLyHiDl/d0S1d4ljOQZ
xX0Ir5nSJeJrwgojlglWSKhL0dMJo58xTWmlHHQA5dozBDaOq66hmsuUNPGQ/iVz
oyMYjEnPf/Omj67mYIMI9Yif+9fKF5vA+Jf/PCVpF+d4YKTcKKgXklG3Z1/ga6ky
uWC4NZEr1M82dwBsI095xDXaL97yUqfJfymDfBFYluKJstxyYOHgELXire0wWW+k
dRF0brbK3NKBRVhgW7OLJkMK6aOj/MdsqNFlnS8fsiB7APOXVczbmPSstY85o2mV
/AwF0qPPhiSbk+q9kweXFB90GXG26RrStWlcubZKFPWu4P3B85ed6Cyb9OwCIjfc
U2qFGUlG0s9eVcG+rBsOzW/hlaapKA8jmnaoAZYoZ5u4hX0s8WT2CXkqHJq7XMUQ
styC8JDipjfsCwc0ZLKSPQ7+LCCdJlOCak1j9MTSsgPfRDcRnWLGMMJuVSFhzGrg
tkiAsHPIqzEUouQwN46lGNmodxV2ysOq+gCaQ1Dv2OJCca1naMMvqfHsGrb7jHtm
kmePHmm1NQ/ugnmSIbDuXlrgT5+1Aap5wrXC3n7lwNmpAUKCQWFuwjSXr9YMdR4E
2oOOfU3BwYfZbViwvxFTZyQM0r3go83xIL5xtryT81ygPuQ5dY5x/5PKT44yU3Dc
HkwLlSKtyShoSl8JQlgsUNZq/MqJSnYGDW/Orw3WYCrv0oOIrDn893SxrcBIFrB2
+FXDD3Q1IX3sZRnISH0Pz42bxh4feEsHdVHDRMKkn6UoHAjmPm9qCRdVP904+qLc
RuYs3hj7hWPHFZ1puNXum7jRzHLWUWpHX6UjrVzDNebReEbt/pKvjbEpKh5arIDV
KNnrKB6Ctv/9SZ9m+OEOavMVgKoL0VaGXAQSqSWFMfIymFRQJcyUWk5c+o7FXE5G
6/fGIzjffj7IOeyyvBrZa5iy2Fw+gttXAy/H2JitCCJzpjjS62nxG5jKlj7d3ZyM
qfKLEFd0db1tBnyu8gei2biT67kzQSz7NV2OelD5uYAO5KB5YWlQwF31gxT7D8V5
HhNADg/G5iFxjVP1vcmrTUOdza6cq9XN623v+EhnvYkCGNucIQV3Z0QVwl1842OQ
tWgN+7Tdgt/gf+JcXlLAhm0KtB1DXMJ6vtVJjfRBo3fl2mNqY9n98ln4skqCkRIx
UkmMj06Lz5Ltc8mM5Z9PLCDuIgyuL0wIrmfzMf82ExqkUswBI73uthIYAYaIdPA0
ZB28gzZf+kywcF1KVAzc05ITsy4zFtNffSbCUd1loeOjknkgmeXMhHjmjyhiGSaL
WusBPrIpULDGl4pUROc5rJZrUeNqymiLJsoNhkAfgqC2qmEXXArvKfcLRtgGdh0V
IoVDOZG2R/+KqT7d1hujYotLgjbjLF8JAwe1m5jvMI6TacGy6jU5pyvwGaE4X912
TSp9cN2FSaE8IlKgi5Hv5Sm6003INyA5Xa2UtVBuID9wUkP3nc97l5bbc/K5bjC6
5Pc+41CJOeMepV4cz9RVWxAabxy970ijdhWQrIwtJ4qw/ZaUsHnwZSQcqVO193j5
JoSKUFtc7iq7G3aq3RGQAKAmjF0V7QaxSaSmcLqQa9A7LDnfuJPGJKYHRPVnjAUY
22ZpjsnujtG9r8NxaYuAFBUysg6pnqg5Yz217cyJO9oShXVtLwkM6YLSfQgjmi/O
4I/4aS6MY2f1B4zvaEiriv/wayOafpXFDQSfJKVDgbjC3KTDBFYTAQi9VA+QLSk1
70PZfpe6IawVqJ6vMc54t/MYe+Y07+WFVeuQAQ9SbdRv/QTwfFwV8qL/vi0z+D8K
VsougoY79hk6UZ2nLw1jSUc+JZPdneNlsEgAXQWAObP2rQ5qrMerODIHoLLCtuy0
1fm88Rvo2Ej/Et0eAGGrEodzzphIOz3w2wg39gX0HumkKUQ1fVta+IIG7DFG2kLw
vVnMkSClJaPq602iT72ZY+MHoeNPN/ughQK9yoW4TYeDxRN7tNHkAv+NKkdPUteN
V0a7O42dAXL+1XZJWB3LpPPHdrbXJDulddZOGJxKH0ItzLsrHTGLjGV4s8MjigD8
NXm4sV+1d2HotgGNozbU/KSXCGb+R6KGJJ8anIJQTn8jN3Qz5S6stDzGgeoQ4esT
fYM/z34ynISbC2TjAff7LJvWtad0bUEKfsqfrIA/CigQRPAonfk+Aaj8BG5UtkoS
FVWVJg6Wn00VnZwfMLEb62/8Q3iIoBFqYaJNjknKyNb3uZwG5hbvN8CRW2XJRzQg
87f1jkf9YKEb/PHXaBmqpPNfDyQAwhaPFo+6JtbYMbngdPcLC2zM298vxKwLxb6A
lnyKtzIMVi70uvaeX7id4yTG0bRDzoJm8ldJdWxVlSzJ+WClvBGo2K1j9b/cQXJt
iXN2oN9sVGn95avhHz6020wRMGuocCA7I9K+OYgm3gFJB3ejZHU3WTXtxgC8uEv4
u6bCCS1fXon3HHoLkmhy3vfMXniOt4cgEMHpTQPFZx/MUKxAHMCDqLL4DHlAlEbj
jjr9ndB8TQ6Sz9E0+3QFZTqq+JBmTCQk8Pij7M74hHmy5iMUbPz+hauy4sVTS6OO
ganEp6Bws54qOAtvyk8JumKYHHO+OuAKcSBP4qfz/pUPlUtYk1ZeQ5c1SPBAOHHq
UUdHTEyKaGqk99O6w6AND/SoMqDG3UqeUToVTuq9k7XvemOeVFv+TfAZtxRNdbJZ
lbzZy0yz/RbErZtqMcR9WcpwEiaJ04vaTKM0CpDdlOuILoy2kDb7Xx/85wBrm0mF
72d+MUf78fgjZpXj4f3t4nZGU3vR9XDwEwxngQt/IuFJpnkmWhnRTBug2awsIzoL
EMHDQPkR7PZKAVa/4JT5pDRGnSf4I2T9EE7P5m5mp94qbmd89m+fB9IwSfl0mv+8
VWizYl0zshnTha36vPZE70Sq4EJPdgfeeHAJt+k+T126UqDV/rnj7lREYSAPq6fT
TwSxEULQzTmcAFFymSnp3vfFlGK+GiqukQa685FK2lPiw2fjP3uNe0s9hzs9EnYI
yU9ilO/3ZVskwj5KjrRXKyX3QiBngQGfagDAKUY3GFiA4vMwNBI98tV8+1gYqk9j
9qQaxksz7muax9cH1aPivVbrYEv9kRcOw0laQVk8NsodS8BfI6t8lCxIZrFZpA9R
o8xrWo26jsOPQcA6KTt6WSCSDHXc/UiHIzluCDhA6/ncaetS9Qk6N+zzu+6/wIRY
0+C77uL0ECMpQrkR1ZRzi4kexM0clHQjT+9h5VGCdbvpt65YlIlBvFu3xgtXgY7F
VNN/SEhaz8vWlTRgN/fy3czAREC60feoyegRAV4yawKIA3uv6ckCxD0olDD+UZhb
pqG4PlNNqGOGGxBl2v4dW/BLmbFxOnF985p1N/EK3ijV8GYnDvQXgZdolY3ipw7/
TFTsg4gu2+1doDrHGP8eZjZ/mtrlQK+fJe/PoYH1euVjAU0RxCXasr3bc4NyZHdd
khMt6DcxathiNDZEslUCSasDVJV3m0K47bR2m1GChc5504Pp3fo0K7KjTW3zv1hS
ufmiiVLezPnLy3G6uXkBS2ZtEbzKKsdBkZe5Ph0fsa9UgqP/qWF3C0zvOaTRun8y
cXAEdnps7N917BA8zBC6zUT/YigJktT5jkbRVcZqF2uRWfaYiO5UmF0GdDL2J4fp
vOaxy4YBnNqMDWo0tJYxRNKIGPM5w0eS5hbCaw1lmew9975y2qPfwihgNhWBd4q/
7IB//oa4gVnjscNthg9+f05jItbapZxS0vswGUWkIUYvmE0TbNK0oKVx17EGbImH
0saWwvZdk7IHFdN0xf7mTZ9NLk3PdUjF7NXB/aXdUQ7/UwHlIpqi0hJm3IGNASbk
RdHrsSheBK0ZsVii4yGFUP1P+dRDmy0Z6ZdSUS2OdDhJYztel6BZ2LWN7tmjNP2U
HGUOuxaAv+ZDc9yG3rpH1YBIEhDlLiI6DqOIdb5dxDL8ySxBGwMSCDqqVmBu5dcU
qGP9d6DhAvKRR54SAxvQHG01fOLWPd8gf4lI0rZs7FQPKVkW7F+ojlJ6Bq9S6/6N
8/M0Ginc8MIfoygT35jZWcyIvwt0i/gulu3Z4cb6DhQq7YYIKoFpvmmxqlsjoqdJ
hUAiOrql/VxMesX7jhazgkIIWTnJzfI/mW2FptIYE0tUpNPBdnXlbEQv96K7ro91
10Oza+1bB9dE3H1IXkantiPzIcsIlYeVmwgeGobGo5Z+odb7PpMHInfIdbmhm2RO
A/BBRTsFBYEzzuEGvvE2CaUS9jinv7fdfqkhSzKtSfdsSx8x5OEhpob5IjY3bPTX
FoQbco81ICng2SKKnXBmnyPLu7SkEZcH+OXhQczpJbbxq4SVlZXz95p8jJdx2fJy
p5P4W7o1vLJufOVG6vakFIVSbbwiYR2cElQZPCVWuso01sS+WMjeGfa/6nAN1gIk
sbbNU81wOpEAQMEZV6NMgQcf9fz+VmmutJGObTtXrWJ5i2EaVIDVgzxpsmW5tO5W
FJ/03JarE0pmLn8ecCLKi8Jw62mgv4SxK4RH/iVGrkeYMpBeMnhd4DUQxx5xu7+d
jIE1Dg+NEyxvpuwsoTku1OLK0TXlUunYeOPXEIqbOOQsNH/vXtcn/ePFq9AjUR1h
o/xD09TVlCeazYCIqpFJdUqknNPEvl48uW/JY5rdwY3k6obXHNqouPwaJppB7eFp
sCx1MuAPylpz2UEap+EsVWhSpiWpgQOVP5pDnMwt/fzSPORqstkNy1VkB1dL/VzA
msaAILmoFS+WFJcUXFE7o7EQsEU9lNvwYlG79CtokSRJHRbGWbjBMPPPgU7HiywR
s4UkqYJ7ISTn3c9p/TN7gHsq+vBs7Lx8FJPFFOir5sR3QXEf/KNs0kX9daMMvrlM
RNwGxilq80iwTXQ0fCB6qrvSJp4OAeoXsXBLQ5pRwF+u5PiC9TJxRTNuhDJfLO6O
rde+3tMTT3ii5QL6YuWpsnKcTC4tSwm1CB/tgpHhzvHDKSBa8N7fiMIeZuaAjs/N
4aDZovvnsau/yUkrDckJSBKLOWDr4efUda0LW5IHI8GMldxMFBHkorMIJ0bOyOgN
/mKlqWnfGShfuqADKfYKMZbmkZ/COLahVfzF1Apb9ux35iCcSWcidKSPmu7KdAVU
MBE7K7s5Hjd64/9Ci13eIYqA0zffprcdNkyn6vwK0fjL+PYAql/DsC8/gYhOKwqC
F4fqXvZXqhadZ/SA7tuXCBoKT2lVZTNmqNEBpnPWlS+Mwq/tdDFfP+l8Y8kXeVTw
tm0r3+Qkd4VRQAtl3DorHs+abUKjBpaeyLlZjFzY0562UaVGCPb109YwJ8NiOQnj
5rClA6frulkwr2R0p9ppeLtHIep/4d4OCj5ke7Q5LoE/kGYs0ffOIoSIL0woUVRg
yzXnIZ4BpUYJfDaiPfPNbTetucDtyKkw0H20D1Yf+nvV2OETidJd/cFMP8MqNMdo
OjmjqGnDeG8OGg2TiU58NyqV5UeaiiUMHf4tVu202Le9pbsKIJkV+L9gT2xnqRhq
4aILeC8JlEJKnhH4TVsvjO2pLYYCC5o9I7dlKRf3N8z5lAtrdWs8Ym+sxXOSZHgG
FTuGIj11pFxZRX/Pu0zSmKbL4j93Ai7HGLxEkegsm74fONOxy5804BeweET8h61n
2+LN/2sZQ5/aajPBsUOFPPBkKfyN5hMO5tBWAyyVYtfT8XmXpGjYM3sh8+PaE6Yv
iobDDjj/RXTMG9tiBldZ8d9W1+bGqEy5SbbDHCCryKJy2LYWnfJRF8V9kf1rqABB
BJMx1iB3yn23Bwv07XgahkCEMBwd+ACsLfWTo3q8nODKNj9DoD7V32TYpEueFN1l
T2cAnOYDvzDOn/MoPPc6skhuZxyzp8RUqmpEqMdp4U0WEDU8RX68/yPvBz/l7cFN
RpRinBbLv6CJcia3sX1HR03FCqssL7ZK1Xyu9JURnXv4H+hWPyWfUxkJtjSg6rVJ
J7sOHDRZmgwuaRtjfbbp9fsIZGyH4FSJsm/Ng6PoGslTRSNWJnwMoY3mn/UsEns6
CcBR3w2dVNNMFFHE9qJ1s0IjwtnWrYoIl3ex4UI9Z3I7bL8cF3CeQ70A68n51peG
MlLmpRMWYiKMujOyBFEjIJxQoCXpg+vi+b1XP7sRyU1/PBT7DNispqBrTk4kIU7f
Hrq9/LC8wbNpyL5GhWY4zvx/Eefy2unVt6XFM+sDmla3SZEJQ816Mhfh0zdwVBjf
9DbZksE1TpB2zfrADq+mA+YkiPDh6LrUxRLQ8M9hTS2cfBJOI49vzU+XBGOzJJ0k
7CCDp3k+ZPzJ5Y63Ydc9CYSAYTsXtYbzGjF9M1AdcStKQPLx317YJiLH7o+zJYy7
OmdAfE77hZSHVA9ChN5rUc69/5hhk2uLV3CetZej4k+EfJi6ptIM3bSHvhJiHfHA
D4efGA+lmuVdk77FqPPdEW8PEB1pkVnQ1DO//T/L6Vy0+wFWKBN4k8FmAanRlvsV
ewm9n1Jb5D6esE5P1MOEEZh93jckIhK1F4iqAmNeyndUUYm9A0igfTLtZQugoqw6
0N8Ke42IPbniMzxfHh5xxZ7C2ovFTTuvhIH+vijDhsq80BVgWyQoJCBSaA+2vKrn
jOY7vd3EsUwR1+jaZ4StkjmTUuWCmdrMBbulNfWx+36SRc6XxtxIQ5ql43JA56E9
fc0vuRKiexV4LPqD8LsyUZGTNJFkL8MLfCCJqqi66ccT/PQM7U0Q9K8UUmF8di+L
+GtOYyynKYEMBQmHNEvch+fDudl/uz1ncGbSD1+wuS8jgTJXBSYnl1XMCGDIjBSz
jecvsmm8iN5tse73Rk4Z9gQXEmT6hNJ24SwoqCi9VZ54nFOOxVIDhWlXBAgJa4fd
tiOqZwXMEabYL0VrcEFcES+9ZpGa4Yaspm33ba7QktH5/LUd58S8nSZu39RzyY0B
//Jm8mC/D4PBXEwFtp4o66zwp9Ir65CztmzcFzFHXiZjwzbMr93yyq3dJnyUGRe+
Id1rFOPRvbprLyTERtjVdQOvr9j+Dn6LoeN4Q9HRrqkyiaZK+kou8+32dcawECr9
IFLU8+4+q2vu4rStV/ze61Vwru+Q0sh8qUL5OkxaoKxHZKUKAtUIQacPEJ51TMXa
a0Zhd2Qq66SuQ7lRmgrwnAVVhWNNZBQmozrOndj4bgMnT12oWBROVfjexIISircx
WZILrFBOIt8+v+9DtxL+NVoxxZCMfDDku4e1kMBZrt6lQcv5xeuu+INzgC/3MlnB
7hJs6t+5pbq0pocjXmpVZd+9wAN1GewGjZ0Sa3dEHObhy62x/SH0El0BQuoSeH6y
CZDXJQc9yoJcTaZIR/FPMaMGWgkj6uj/5UYrdSIMqAno+LFr0zg/i5zdW8T1fEwE
TEnGXc3FCz5XjVbAtPIJFK80lpqT4l1MUwu7iLaNJEpkVKEZdcAxmGbDCLXNt2bi
zya565Z+5/UhV7hRvt+TnHB1x2Rabil22AjWivRlx+FrQNbs5juWx/V2tZmMj90F
QqTOA7RTCDI8crneslRaJ40+UMzYI8ATNIeTN3js9gkfvcpt6cOoF16ivzu88a98
7k2TfzG9jWiL4wlp29RFA0ADwxyK9TNVzTrx7TE3B/YVx+HRjZS1vATC/fidDHez
s6ITQd3Z9geKCGTd3e/tbwvPlDawt6aFx3ZIwnH7VscUnInpsc1RRs928No4XS7I
R/V9AscWH8TJ6lzixaMPvK4X9WNl5Zy49esDemAtlA3M3XIriZe9fMAOqRh48z5y
ApqUNYjUCt3XKvYYSIpc3jz1E7Hl6qCIXKGFxow7HhVOUnby0leb4AevyC7m4csK
FogByLaO+OzR3jBzOOjDsbVFdHmixAq8dxDYxMOvE4s3e1UwdRFr01SywdFxe90C
i602kKqdBfYAlcnkWfPA6L+QyUkD+YoYnI8XaDU/gjC3xkTMoRpVMcwq6QmpfB2A
RPmr4GrGA9ayqYGn/GPbe8VWTETdC3byPj3eXePPkphUGmM6TZqru8Ih7RTHAL2E
2Wg3Bk6EPiwX45IF0fW17y9AxOl0THHm6getmzkCkQe9TRVsyTVrbzjETolmID2m
6Ts4yaDLrIqQF+QNHU423azxjIE1YIXuz7S+TJyUfGUbuTh1djmI6q1mhiwyVlwb
effgLeoe55OW9mvlFrycUVy3NoM/BKgEF84RwB4s7WimvR7SM/VSLJBMgXkytevF
UvWje6uCH0nUyyqfIkxKS1+fWoN8KRW0vTcUgiWSB+zpBpimdnuASoy+2lYSu5WY
04EN3hWfd+c3K82kA92v2ZR7Fibuv0wmXnUJS3SWbnwoQWLQMXeXstduNMNAyVw7
nze2FclFtNwhFLkd2O3YOqXSu1TQCX7wz4hps1juVOEOXPGxbq3E7Vrxkt4SXxt3
IIaPMFpIeFtOEsByvp6CKspcZjaL0bOZlx+kCvzB7Hmv5TxfFYddg2eEfkvBu1OJ
rkwInajTvq2IJdGB87I7pOh0s9ocAPy7bJuQot4GfqAMyU67qtYtNWWDxqhj1nqT
3NM2bcpr3j6xvYFvPLP94HGySW3XDwSPTWglwN6snxRP6rhTybg/HkzDzqTg23Rp
rvQFPuPdBeS3JlcGahDh3cDPdDRtlflYnFu2kw/+5Oeifc57cMAkabJHM7qPeVJh
zm7HA+W52CeFuMQiUX0Nmtah87Ga6AxcLDcQE6E8nnIbL6IVXq8aDcYVaPWnzgU5
6bTxX79/g87vfrFojvBkbC70UpByCixf/tUcss93uUP5KCbtk+r4L15OJhl8oXOZ
fDeTn6j9GvR9St5CfikEurip1wOJanlCbl3d7yijhT/eR8mnr68EzpGVLKGz40Tf
xPhLPxyC+blKZFwe3uTHflJL8vdspy+gDy/CrZuizWE8go2yo3kprgxQRYUyWC/F
BbcJ/XGMiXJ4h1+wLjtpbupS1dHrqwg1b2HqtubUfkpZmspVyh6SDkrnD0aFdjWG
zbynUdZJyCkHj/rVvolR706O1pTHw6jNPmCBr8YLwJAXRc8cScCL7T3IYUURHJRe
mgwm7c0iheR70Qw6joh3MyNIiGiE/k+N1v9jTLktNpxiY1pmN2+eT0+oBJN67DUe
4OaACtQNwSjRrru/gXef9S0aVPXKnqekfLpZf/kWdAQUzX8MGoWS6csuoYRmoaqe
SHzqgcjqq10Yt1hMRbojkSSBPjrgtyxABYxrtpwjOdXL44OkgchTVvj6KxEyqp1x
dMrwcYetTmVeHPULlFweIgOqGbPHBQmXTHM/KPlYDj8oKxYYh/3sua4ggg76nUpA
i+KAmcoWWJ6c3FoZV+QebQ0XavAP32PcR0VYwutbwGbg8DvCV3VrSfzenW88Qkjg
zwcKk+J9ynNHlp9iU5+A4ZkO+PUGh7BxRh5fpjS+HYf5utEaj5DT5PYRe+WwzBaf
Zcv5csBGavKsWVNn3uYCy6fWHuXsdxCpAJ8nlGxYOOqwoPT/pG/PDDrpZ/98tA1P
ZHrcxZoDaDKPGK5ihn01zoEt7+CMDQGIN2wuZoSV3Iit11Ok0+4FvLt26R6HcVVO
POGF4DVxvfvs2JoP1YEAY0F1ou3A7LeIU5zKtY0UTU54ME7Ug3JyfkvkI7xui40I
h8Tto99Mx3ceBFZWhBysLatAtubfmwasnqgRlfQh6Muh/EM7gLJsAIqJiZMUqNgN
8SRxJHMw+Lno/sZb+BeGnaee37H23wKYr1WMRUZAxNOxvuV6HfkeCSuPOS9V/U+p
LNAmxmu0YKbNFzcOZBKbFWABTCuAr/Fhd0g+bmVc6UZra7d8QjmGs5nJgrPyBaOu
tqRihV/zkHwTeP/scrxAdk5b5y305OWvh/eOHrJ21S31blANdxeVNisow9RQu58q
0IhukUIoKAAk+6UfSrlUKSBSgatLSUrskcc1yjJCuRdp3gpRVvXrlIBP1R9c34yG
NaRlsIoHVbID+8Ku8bcD5top/k2nKimOaTw1AGiZPLfSNrv79EiS5n8YjcLbcuOn
vCHc4elvn+56wTPgLbcStneJ4g05dE2X1T+5pXiF8YgFRJyrfK/fqius9YE5a1qL
hxSakZ9P/lV4xF4QsFNmywmadhtU0M1xLngBeKwlgD134YOjLgdJVbjQySnz9PRS
hAUsKIYSHInQ0MsLGUmH5hHnpKqTxnVGiqqmmDDo0edvHFp211hkvTUrLjXrYh/Z
TRgvc40cGqDUBhBb+Mdlx4SF0fzXU+0x9DvaR0v591+KHjjYlKCKRYPADoPgvtD1
9uAdZb84x4JjIJhuLZNDoh0iURWwJzg0D9q87NRAIJZvEY1fWYuJy7OY/LD0whn8
o7k/1BorMVk1vO2Za6PXrbB3SK+Q7e79VUYiHtMCAnwMp1y9lqyXej1iwh+JSrno
RwtAigrkoz7v+ExcPFzMRQeWMoBxbwy7nl7KWqhDVeXJWpXSVmYDptWvuCM6ruDs
VsV18LdJp96Ssfo1tDV80mhI0nyH4OUaxtCUm5U4yeQjpwDVMHNybmV3DF2VZehp
Ogz59P//aouCGvCmUkrnTN+yMmQ0O40KHb/7T5A8tn0EmOD407MKQV2/H3bf27Tt
kPtGU0OdD0sVpS+B3cotkiXlaeF7gzwDKkx4Qo+tOIeeZwkJfVLbOGDyERllSvWY
uDq5iLmgO/UUd/3SeE/we3/0Xl7lD/hmpBUCshKeqgs/P71gh/oAwyoJMEDkFNEi
Y8qbOCZ546WTlATyXqpmvO/vMV2bfNo170Q0ty0BpoPxUtZrp6RTTmBf3p/tZklY
ShE+PVuwPmxCzn7//35ZSYBg+TJuiPaRhCcIxwEYP7zhKyViaS/4PmjyUttgkXqq
2OTSngRSKYRYYG3gfcd+wWdeUdQ3IXuL3ZVFDjnhKwC+p3i6anv2GOz7pKhuPzWv
WNbPpg1ZkRcAoKrGFb7r7fgOBpmZxm9OFxYsLD0u6fDn8pzMGpCyTmgUn6nJ26u8
/OuDYX+GTt6VYswDdAOu40AZUPtUKBKPEYPMpAybf/yRbDuGGkCFg3EcSCNbbFW3
ckTAzbpkeyFvvVCRecYr+Z/a88rMDjckuhe55xTehniJyx1qmWB7rXWuReuOEmDW
hsM6IPRefBeUmt5TOa8wQ9+7P7acgcxc79ZXJLEGInPYy35phwk2VyuCllx79yT9
JY9IOSXPpZal/EhO+TpWzG8r00v3n0Cf4adZujdGiqBw9DIieDdfMaJxtSHI+4Zf
l+XYhPPNTuvtdEV5Bl1KNLCY/j0kRDSTVbvCCB/lt+jhOkwYA7MPbeblk44qBzsj
xMoPbrPIUWQDCk0ItL72scbeR784OPwo6gYYbSI70Sj7Jb6tnzuQgMnEfQPB6mBy
3ZAV2FTUT/dioVXrJ/ic8UNX4R4fy/OeRrawP84xTewRJpLL5f2xhCtzjLTARfyR
zDg0DwsA7qFV1kIscoTwHx2sJ5yn9Z8MKeuPdGcALzARVZhKIclrvvfUq4LaX52B
iDYdbI1HhgnL1w1KHnZZM3Sr7ETj/4GvImtvlLebVSw6+r1piAlzKJTdgdIbjdjl
0qacLmal1XsSOpHSq+EMXvzgK48O4KB5DwbmkSbxomuD+3SCJLg/3ATJNBfzE5ar
uG5nAZjbNlPfsIAv93LfC3tICfpre5g8mhPxwCso4Yzh5uN8v7IG5FubcCOkisOt
pC3e9SpUuDTGGTf4rR7BIySoXDGBVSox71aIT9OBy1wXyt6JhBSpteF4GOvdSUoV
ATqGHUw+tMHbMai3d1WBOqED3J71CGoCLpTSRS9fRhdsCUSJ1gps7MinqZBav3kb
T/5r8aY+4pBArIOw98XgQ7uLM5cZx1h6TDuDMwhrasb+A8ERK9dh9sOFjqaQJXYJ
2lQVCHZo65YJqOpGens2JgbFpN3R0tK3+VRtn8DmcpR96afXIVHmgi5+Dc4E8uRD
M88FzpqUbtT9utvAVzE6323XEMuW8Lyy28UQ6Y5P3gaqG++zpwBPc2aIAGNklMu3
vIkbW/m4ohUkv5K2RKSd7gJa7hEBqB3OqPH+BAV6T2/YcL5bLhih5uZXzLmTA1Q1
lAwqN+J6fTJtaDS2ST5Lgm2EMsRqMMlMITXneK46tAuza3zjBrUo2opx0hBIN0kn
XP6MXVIIvHdTHYldllhECd2EI7xojhsaB8ejzoSPwBLx2UFesgED0FWqQKadRFDt
wFY+Hg5tsuROl5KdHuyipCm1QrojWmIflRss0WQP6YPAAOsBhkEGghd6Qn1pApxR
V+M8DrBD5Q1K81HtpoUuRNZap0VxIq1TaAbfN91WzlPuQ2pA+h8uIBvKwkpXe6Y/
Br0kOow+bOx5QqoIhxhDqcSziSoRPdDn/y6BbsWqETx5AVWJczF8msX0SeM1stMY
LWSIg6OCYtsjQgypZTjkeTkzXmgEThoWG3CQB5yYPuNVLrbdXZPmtxRoAZ0spi7s
pAZLAb22P97fdZDdHqyXBLArtTdrLJ8UgCMkyblpT6TdrfvPGFsgTXStGOfx9V6i
2mQ/gpgWttEJ72esmmD7iVWcCMQl0WAIZR4t2qn0uITXNPEYFyLdLcciSCARcj51
/GJdbCUhQo7tVd22T85G1ljBydriCq9OhHi9RYXFqYlrLAt/bVFJMo9ckrq67fXs
U+/QpSUXiKBpXH13TLK8J4HMNyJmGaVq0UXv7xCB0NX+xs5gYB6wtZaj8gG/J/rV
3eZmmc+VTzpMmrL+nhseqx+FDP3qNp+DOhMUrmieIvzaY4mWqjYuNSyzBEp0xWad
V2vRZ7BFLP643cIMvp4LpWsptztWODWTwRDPoNI0tSiG/Pm0UIdlJo4ND/9KW/j+
3kTde7YjHWeXl8O0kmRKG8VZ0U+FkkWQvI2yoayCn5b2/50yExf7vaXGwLtxdhkh
G1SG0BMKbGeKXRKWznlm4VEmMa+l2VOxBykn+YdREndA6s3Ocgneh29Tm+comD7l
PRTmr/T0tUQHIfTP1jUsg8Kcbm1fzet82C98RGxputih3fvbUyGd/STJNFeFJh2W
bhkqTMsfGfpWnhEZcD234MtNQ8djJx9tYVg4gPrfIhee3ApphGc9JyX/t9UrLSYF
XOlqlfve8X42V7z1NPDm+fczmn7tI82xrVePqYcKMlLYFjgqkE+CLJqHB8m+KsnM
S/KhbvoKDMVBjakO5qbLtk/izGHUzNyvPfLkRJ1oRRulgDSzwJWv5DcR/pPbgMqm
yHuhJ9+0oscM+vL7HWVORgQkuKgSAQTeMuIVoWu4OpbYUHl4LQUP5e1taicPEg10
lXeDi5nzzYF1+TCfGoshVIWjkaekozCIoUYL9STy3GBsU1RN20cCIbeAAKwxmk8/
lCthfAglzRqfQ+6AkY2vBcu+D+dUgdxZukdQEedWiz86GPYriVVS0WidIXHorxVb
sABKlM7DeRXqA0/b77QMVLaAvX3WDE6gviPSKfO7E0sE/YdjHoULj1lePorL2m5j
n60Kx56wEc88h+lHPg9dvcBmhLt25xFfsVYtpLMrKKN5cJuJ7uiPKmU8j26tv2rx
m8WTCsj9/UFICV/jlvYx88SBvt0ortpNV/MoWLCzH5uiJl/suFOaG7oyOlwWP7G7
VyK7Q2D4Rkms9/HzZURybqxwmLuxAiViA4BeLhIctRCqZbRF8bZckuCqVZQykGJx
+p5QhXUCrFYRay4kHUWB2kLylmKPeWFKQSUiovhNhBPqfUZ4FFXzVf6h+CEQAvi8
qYpF+u1lKhcrcz0x1Hjp2Rierdt/53Hr5ETnJoT1SQPMDzAev7FHdJlugOiJInf7
uek98dfXNZw/VZqiF2Gkvzp3D1TomgI8cVcrRJ+gPF6T/OmdDzRwF8GVD8Z+hsTn
n6U2DlIW4aPW0QJidqQ3lFki99PTLsqRJ/PS7XH/do5+JD4J9aNg/zvQFaO96UHt
Iki95zipUkzZTB15Zgtbx5momsEtjtDaYdw9VEmSmbPsAmCimlxs3ikdoZP2E3aQ
ovRHvmXRG84yxVMPvCQgxpFlwF59Kr6yX/4YgcbM/XJMYJEvirk+KPD0d5VZDAal
Tf6/ufDU8mfwNAFQQTYqGphhtR/y8FsQSF8obsDDXATjE/zA6cl4HHtviMA5OvW1
Qk8rSoCDmYnhmYyVrFGOZLV3k7kbt2edRcvywy/utEybnnLW/Vn4R7Qh/nxvjsEp
SHlWASndnTpOVGkazm+UTprVwZe5VzAZolPHGfUt8NfGHBqrHUkp2zIC+DwH1obi
MtrDSOgguXBfVVRMp/qrcvBgsHc4yRDiSVK7eNwSX/AwZfJ20jdgA+rgoVdDV8iT
qPC6pT2RiIXMIcu8g67G4gugbjM//P2kk0lFXKmEJ/tyulDLJQECpSSBnqVmpnAQ
R9rgl8kELUYSikwn2Z0hjeCf5tVcc478fc7gkStQ0I2qKo9oQ04UUaU3/1yknDD+
uUq7Z0XTs7jQ/5R3+lPMvW0FQlV7H4/XLnnPlwP8qQT+jE5UOx9txruLZvb+NW6g
qSIjGylqrZ2Vw7VwHgJtY8Mgw2hohzrGtO4gbRrCzwcFCoLk4q79U4ojHR8KJ7Jp
LJoCRhGu74kuSIaQFHeaK59Mpy9cOpoiHaqywGEMsE8cOaAT1OMOaA8QLeyCUmA2
s6Vg3WIp28Krk+g2+Wk2Aw6bBS78S6QFz4xf+uvuv2EV9S0k99ycQ6pleRJcz6W9
A+H9irORwJsQf85lWZB8jzLfRWRFmARhZXysS0v/2pZxNf7BO6QJWdDunRlUnRU7
bqJ1p5eJGAmE4nLkUEbjes75r4MTnT+kuJ9Vo6hsRpraJWE9KkuRdArfpj4hxCuT
GLdnseZ7HydNPljzJXeOFYIDQVWJn9zHg22hlRot7m0rpJ8gMc1hzA3exY6i/xwW
owhirOf9BuNk1BxiGmiaoT/tUQxdc6gBls3haAGjEs4wQm+9vn4vs/KJpWzBakOn
c5pGtRw6n35i9EaZXsRQSeC0+GXEjuis8vkboODFpc5Xa+NaB+vG4Acb2Vl2Yhqx
2iAPjblZ1540eIBjCZCRjHVO6qSG3u4k6io8W8qkmy66HM3FAevH4iKrBTWzlK3G
yLFm9FyqE2xqfuUY0G2SqFjnwsjll5M0hWPhcU3KyH9zNjPLJ5uot6bRGUcLlldX
J70W0JD1lqGfHxRHjwvCi/ONvt/U4P1m6Hz42OiAVWg+9p6FbcWIgNwDjus83fqR
t4lPGBE4Dw6IHmGp0NEVFuydhYEQlSOlEubHJtelnl9On6QcfJ+zNGsF+IoVvbSo
kY7qTK2sL4eXtggAFbnHKFxXwHfWUCpWN94HgeCZsDB8HjuBcS4Y0SqEAjc11KN1
tFENgJwVH3t2wkR86sYd8td+jI0lPsEFrd5pJ0CGteL4wyFqvRxbiCPHvzc7io6T
fsL41I5uvy6wwhCH33pUZFOvaU5/dNn7jekmqblJmk+3f5MU7N6vJ7ZTo4n376Ai
ND/61wylKChT5kc10Ut4xuyynAts3nJc1dYbYrv5S41oxXiwG8dkfZBarGPYZeFP
WsPGDX36NUISGvgGw6eg+bxig5SvtXWKn83/G1b9Zb1vRXO/naUkrxQqwW37M7sX
CmDo2tEjE/9ruC7mf6yhXY7wDV24saYNRa6nBBn4a78T4IofmYBT0RfFVWH5RYa0
tEJf21Wp6x4KmksqplcDwAJRlDkmwH0W+o7WscsJd+UdpnQe9kzqA6MVPyHOrCq/
jOxQ5ff+4CD0XtW0KopPcxi4pvvOLXMOEZ/53KLwkfg2PZv9BWnRfeErSMrVIP1C
7gdegnUAaNtKWzekfGu9gWhmOuTgjwUNbiDqoPRslK4VAeExa3//g2hvHL3ITEiz
JaWWvV+CW+FpAhNH7N6R77DG4Mp22nxW5UNrAPrxylOhNNdVfDaUwD+sfeKeBg0Z
EIeRFRvwns7d15GcBQwF201031l5NYQkfSe85z/mQs4nW4gKz+8vUGSlWhfxAGpJ
MFuRHeWOJ2QPs3HLu6cvQBjC3d7oaifbisGd8Yh5ViPKk9IESHDf5L7SnZefjGV/
5yNCow4yKeKDqwrboKpeYvcYnXomU31RdoKDB/NY/n/e94tY15KY+TXkNg+cD75M
3mrs3RT9xNJVYMCxIqSVO0KNN/AaMZ4yhfcGZlnzKorTDbvAGqKEHXdi8pR6O+N1
zL/Zk7yqCSML1BJPAuUT5Uftoaf/eWkLGBglGCYGQ2zBi94FYIN8J9UKpdDmno7z
HpqjejaXKgWdUGnJcCE52MmEgPMw13J2+QW1i7D4aYSj9Ybnils5w/Mm5Crh9Peq
+DbpnpaSc/YY+UZ1kL76hrVfnzdpUTpRaqIZNQWSSGAykKx3pwwFHESDzvWxDPKU
QCB4tMUssfh+tJZrfPTHsqiFOQ9M9OGgv6Q9jrnIP2/kWJidOXBM7ab5hftpP9Cn
yeRzizThfD+JGyeLbWFzg96Aohx2aytQMoXo2TDNLH7ZWOfyzPxfJyhORPphrP3x
YhqiO1bJnSf9HZe9N9it5HMuZggumQx87mkwwm+oNpjXSzrNHaUV0oLOtpc5LIy7
JGmwXmC6xNJ+vF0IUjpMkE6gNdpbvBu25qCBA+IXFuBxAoBrYWIlwtwqR9zmz63U
Rvli8Fdg2e6zfn5dgnQe1fVc/Klbu82e1bVafTwWdRQTe30c70SayK5LMiGelonJ
1A3TDAR/oGW+xe3dU4jnKRTu1SRiumxhPs4zSdmwOkT8GOmduOjWXIHeqSHphoPY
zGjoBPewlsOzCqYRxKxmGS/F9G3cjfp1fygnrPZbp83D/KBEzgFeCxwTaz/p6/IQ
1HMJBzgOIvsMvYpdB64vfKOGF8lMhJI0V5pCdAzBw7svWHF4TW7btNWWx2Gn8quO
VSAOLtbNdkh80FOQ8oEJAdozmAxj+KE20HhGMG1ClNCG+Q7AkimQdKvUMowMzmtV
zukM9KPnA9GYzck9q8iu7TU5wpcWHNdy49cJOd/TlZ2u1k65M1xowrNGI8sskr8f
TwsB9hxvSfWg8QHRPhTmdMPMNHnjDi+ZaSBcIkg61pjQW/dwqYKa4fs6Ie6ybkoR
0mxzVCLZQ3lxMLDhNseY/cyjMezsW+6IwjJE9ZKclCuhhQDT7TFQEjaDPreMTFtC
Cgn9/HSIViydbNxKKIoVMwUz5rtiAWz7HULo6t8klBdaWmGTbCshzJl9vN+sJTd4
yesX2dz3sGlqZMvP+bWCvFzN40/MWmgJz5gU1l5lOKH75EZJeC1Q3af67nq5UL6l
iDKs69BWBboxR+umJtgBdg6m6rVJRkaIEK4frtVA9rNekNsBzSJe5rmMONhbD3ky
Ybdwh1D3DD6G89EOdaMRhXjciFR0QNLEtJsiC0aDHpS0G8PuLOyGpTmU6TP0TWsp
/pumAOjrEmB1qPm15k3IT03sJt7IDIpvk7CE75qtH+zX9XUNKpDJGD+r9iVntZb8
NXiZvzrxfaYJ1oBFFQyiJvEmHsNIU7IeFUawMLCtzGXY474+QpunuUAfY7iD1g5b
+nQtLflAZqLkKDBAKuj33j+G5bojz8ZnGtamxtSEA6oTkRfIQd6hQ58uZObHnalD
PUN4qqMmw4Y2OnHR63j5Qjbd3GAPEaTkPnZQ9tga/q4Ld4rFSgb26aldjx9JC5yF
lWorU74QRsM9Nlqg6ct+xdNXzv4Bjh1qbrts5TjIA/tIchuRwybvKbtvNv4GqkIv
vzfUst4ZO8ov4YaJkfoUVEcnpe37AmHHeqCQf0GkrTy8VwPi41C2KHkTVoX9p7j5
xuKPIwntg1Ogw2FXlcnN++rCxzWJTYS2XR0GqQsn8njsq4jEmDeUbEAb2Zgt806H
wrHYy/CLvARGUUbEA4SziVKa0hr2YOAEMWgvSGhgUC0mvn+HURysowDFgPFtXcB2
tNv5/PFD7zZJ4CbNgj0TdDXF59SFHb+QlVTL27KXB3B4yzckYS5AMU9Ie5KMk82P
1eRm4JKXXcDSjfp1N2Xal15jIT2ytCdP83oS9gjTifTsWc9RLhpkoIUyiN/FTDuK
8HRS4l6x+8TDC7cC0IoweZ+BwAm8CNMbmozmuu7w4qjjjzWIi3BQT3TnxrQVSkwv
wFbsZUp+vtORjY8RdgxwcHDpcCkk9lOpuNFgx7bd1JCW/ubyRhCBiwUFtZe2vzWH
9gWNwO6WtsG1+Fu7LUncaf46AxAj3OKWjsZ1EteIPb/djY15f7eSyY2ccMmmWQ7W
SDVv/AymZSe63ZVs0KbGNOJ/fzIlWSjJcmnJ280+lI+oBDgGXB8A/7givylI20ee
t8DquidyLApZvAMfq6EP/px3QNbvUj6DFcOO0Z+2mmOAZAqVu0CNau7q3ZFowQW3
2wOdBo6BvfxQDX7zedkBm176bRGa0XZNY4iPRA5RNgP9Bllz6fUFl0E2EArzTkL7
KblN/RGyHIPUxFYKfyw3ld5g9FDKjCGCkG7pZHBSfw+kIK2arRscyfeibUT+r7Pi
pZlp5Vq6sDqey80W9aq618jkkvSX3aXjbOHHk/liYdzffDmdZvjZVPhOGe8cwCJS
e6VrFSeQy1nchRLxW54jiSvsekBWstqgCqRwbIQOOHbb8SoRdveRdMDSxtOsQSeG
cKpHvlgC5c3vfnrB4kfdgCYORCuKCR1CiImsnkjKK3XrWPEKWFs8w99uCqX77XpV
ZqISOdy2Bdx9+g3kRFnxOp+MkepYCAyaoxCP96+93w0p2mBWrh3WwRq2JltR0Mro
1wMbBvA7TqvHuwNXB7gVOMxlQpDqM0tC4Bu2d0/ItkNYAxYQcgXRIKsnIQbRVV8B
9WH0fnR257KoSH4cwSlxuE1pHdSOWEwfroKVCCZhXYoIbFdhhl7qi3EE5mggBkCN
wRUbpLuc5+HmksZKuKBs+CzdbRn0ni+eSftFDsgpZbHML4sGtM6C61YAbzQzP0S2
EUPLNRgBAyePshJHbkm6qGmrNaiSgUYn2M7BPREJ/2HibV6jC4sjxwvEeTlrDXi+
GUSLyJtzO506AvTKyKt5PtLh4MH1Ze5lvVlDP+0Qn3haBqA/v2HP+8BR6p88u2S5
LPZVQlLLC6WqYRTbQkbyjivzwnIEtkd6iKmHOeSbK2MAJQ0IKpIe9CpQMOH0OHxX
tS/DG8lQ1vcWFKHu2nzy/Rxdpv9IQwp+CwMH9AWUkgsnFu41HPkEbUg1mjFGmpkL
HuNGxtDWAJV+Brz/6WNkv7WoAHBTeRq6ZF9Fr3xB/aGnvwZ7OxrXmyqXuFm5gFlo
Rjwh748qPnDKHbwaZsbMteW+qf8lPlILODk1I79s8C2ry6Zymu/psDgdFNIAeick
oT+U63GNrXE8MoGTbm6+Dlc0vwFAmfU/eF5E0rJRpUJ9+KLnvfM90LCBiTbvu+Bs
eKKm/N9O3GztB0z5l8uhpUo+04SvPYub9sEx4JE7uYPm7EbvDfV4BhpsKa5hyW+E
Hy8HsT0UybP5pVS3BRVYSPEVkQEjQqKIiE5wUbsZ31b2xXwLQXXQOsajIa3K79L0
mla9mUJMXSEBAAZx53SibgoTeMeHUThIFwZzgWTG9qJ+hizLAOYhTa0+3a0GUmdx
bW6oDreXKf7RsQMLgnn5z5HPy1GZEJ5RKp+PPqK/OvKfTNTw6zaNYovZoavDEgGv
sIzFi+XR2M8Ko7J0ty6PEfwiQ9RNMtQ/b11JpLiGBhG306X7OAOwocHjWZ/+aKN9
zIHUM+zSjGBotwEX0U6A29jAzG87lc4oJFtwHXnHxihmvsCEL3D6+dqTd2toMkx0
TawT+3jwXvx/7MJS4x/kSQ4PGdYzIhLDDR1Dy+ZMQMDt25TAarowO9vivBgzUl79
+XSKJ2OxKmd0Xuhz8punCeVrVV5w9zR67VAKw5F3XIvC9PcWidc0od08Qv5RbYQq
9qlIpgD/wDV9IFE7+QVRN+/awKCQ+t/rorC9Om3fas5ED4dL1RDO08dXlUuLIcWk
7B2YSOVZ+Y23bGUta5akMBeMYHG2ZoN04zgtNpPs4lpkYcxEzowGM9BShB8DTj1O
NBFGjscgwg4A6/fwAa24FfcqVQtvo06txU/un1oNqo7WqtIN6oL8rt+pdCFUjokQ
AHC23x1cHS9RTM/v+efSuBNj4LQF2Q+PPLZWVvHaVlieER99yJfGuz7fM/y2gcJ7
v9Cad8on476T9T87CuMBN40HQkwZDWIJRGoY2dvw1zZZRwCMu6BBuitoR9ERYkSh
hEL/B0SwHOu6IseJqtYoUm4HArJ8rlXtZxIu/l2wL3sWbs1RsjOYV7zJhAmS4Z7j
JJxrHCxiUXaOCq255PxfiZJcgLL46NF3wLTdRwsszVhYlYHt9v6dkY/K/1GZ0+Bm
9gWOEBowkWMPqfzJNgDQ9kzzsUYJSnn/pV5TeT5N2q6iN+54NDFMM2kEtauEkr2h
NjWcIwCmXTj1zVG/RZsOAkTxzBshNmeRUJcsmXREoEdgWtikRmMv2nP4AbkKjK4R
wxeWDpx9RNFljj4nQTxmeKzE9iK/a0axX+9VuVJSdykgvw+lU6eP1+KZEg4mO7oL
cok7S8Zy0LVMhPev5K+mLxNVcXT1cLHcKvqVLtA8is2OPTN2T0GT6c2MLsPGwn/x
cUU002HNqILZPDlBZ5Q+6AASzbfxr9egGqgzZmT6/bevL0OgzP5R6N0+VZ5q9511
Y8eQwU7CGNfVxCIAFO2TqsZ/xccgnw7IkcMUC0SCv/K3K+LMo/QEXnY+MTUwTK+1
Wk2txGsf1ZxFmTnZ6+tQW2x5hEDNNHZTcdqnOYVHXPOntagy4HpKfwOciWsaSdPR
JV1yxZGmjKI3psLx/M4pJm/DD8CdHTDGyHQofNnNh9v7vlgmkxX+IYHKbarDB9B0
n1VRlpVqLPShTHXd1wFDueu2ZPoRjgYgf/L+C2aTgzFOvCE8sxJrq65K9U3qoGee
0IU/VW5meE7qtaCmYh9Due7yYd21i6ZfVjP6TARybxw/OulitrrAQ4F9RJPbokU7
sNmKFtjL+Zv7XL5E4xupQhovx1xkpOQtpEEpqngi4Ee3SgrHiiRTkBC//iaVKqOF
pakiWGzbPdmQlm8Mar0NEzxB40cCTOU+RIy+bQY8S9WWZTxrF+tS1CK2GkquS/g3
WWH6KaA3xmSxaJ7fYjCa0KgQvYOnw2KWLtEX8G0E2ytkeJ/ZmXGHfW6entI/HgSp
l//hpHTdYdEbhMAWZL7TSbckVzMYjsxYggOGCw5pICGDCOzI4KELJF7/9OcC1IOi
n6tY74RrrZPe9lRm2Su+XSpCrhmSTP3bhOSZ3E+wMxMbmg6PaZGL0/6StHZ/fB4Z
Nn0m5gwzCNP/mDGY619PsVbjDRk5QyMGRiqIs0CYZkBif4sFxd7JyP4z4V5m90Zo
GeS8a9V8O1TV+mExiHjIW9kjBJ1WcTvTOAn1ZiTiv8l9opYuvuXoBqDey0JAsdbi
MSmqTjzO9URc+5QmPNzyMYRTlbMrK0d8DTRn4cwae16uGFSmMaN7rJZEdXNmw/4D
9h8bdZR9yMnMXH8MwYhvS6HDrUwE7z52UeIs+Oa/YSKFk6RqayB4TCJawx7E0eiS
blf8pcHd2D+6j4eMHVtUYaUZj/aumADf3dwJfj/T2PHOUaJxRxU7s5xtRHu2U919
YMQfzwIPXcNviBLVCRDFZQJaj1maLw8LRKOmtJpO+b2w1hI9xQZ8LlGioXqMjQVo
x5Iqz4Xoe3WNEfR7foodBOuD5va8TEmUUDHBjwpuXKJv5w9IDQWLLdJAsDO4pJAN
5UMq0NAsZy/CMgZaQHAQBk2varD6cE+eziJfsJ5edTXZV3d93+ykEijssHPGeI9/
S5IVpYhxrU2ifTRqvTchiDcRsy4LgdPu6vor40TbjZebdtIgzLDX8psLL1u4xYpX
kEvrq207PHYC19+wbP2qx7yIlc+s+RHb2//sXE5KahZ4jg8vWkbYyuD767jHAQQi
Ts0ydKIFXCl0cMXunw5EpaQaxa4o1GLnmhLb6W2VJdWp9OZ/ZXnSGg4Euxx8Tu7S
2CX5X0tWf9Ijzdn0JHfPVjggrsV8oA1ghUxqfcNAslQIB0inzYnD4X0lpC3hhE8b
DqgUXzoWup5JT2mlZ/1yHMWAlsgAQhGwHf+pJIXmgjSObUycxcIH4j6uNLLbkK70
Wwtog8WGABJwzlDafcQNU/nnddtkUxbgcuzmiNKyn83FRjXz5TMq+ipltAVsvase
bMJJbtbfFyuQN5hdvkmhKzfSDwnJaTTbE2DSCXqKNOtnhO3A4+CY0OBBi3GqHfXB
m8W0CnAYveGGTqwzPDHsWCChcK9fq4xIB8q+bVG3Q/ALlCj32ICUMeR92bU/YLBS
/GKIbvGeVTpsW8EJrMT3GZ4u2DfSdFyrPuBAZbdPpbCnMYU7cNCbuviBePRCPwtk
0Sp7sN0YNhqlwB9umZDSQASGQ4LRDndFZ0d3IKCK0AOzmPlEGg8lyRKdEI1nDtUo
j2WZyrZWbKsboStPzEpYgtw1iXChuLGC85reljazQFD72fdRuzIHPpDwK2VoG3J1
5K0gksCd+CuUs4kFUJxd8h0InsUPK+ivxpJWKMfkERDma+IsF8mGYIyyVZLPV9Jt
4uRnLF8SEVnAAXcrYfAjOaLIh3aNiaT445PqYEj15c5Ar4uPSZR3P6hVxRwv6Y+b
Fzk2oFOgBSSsw7d1+t2ra0f41I389sWChQFN6ehPconOapPFS/8BUuk+enFtC95P
VFPvS4gDwwKqoI29Fq5DHVITvcbwtcg647bchQBuyps5JSSHKExxNo5gefBi+dlk
5XJCEu1bzO85+frfS4M35No8gvcU25979a4rewx5y0nX/7cjrSxX0og0wvwjEOPk
xsU0jntQ56whz3pORYYSBG8Rlv4HOGnXCmmUxhr9PwY2VRbUf8N1S2cT+M7N8sKO
184jYG4muDAtcuB9Ule8O32LFiHR4cmZEbL9/NyTKkwzvRECDNOISq/m/N5VolUB
i1rQE2rqfW8QhOk46AZaY081tHMbSb7zYSMS/38f4yP91hFJpcPleF7hIjk0GCiE
UTkE3paXFuQEhD9Mtnh+1mQBF59Ejz/TncXtjLHM4VmrlCMeNQEGHIHrH32c1Oys
VFVGWnqe++jxKX8eZkspeQP+5jxV35ZstSJhas8gZ5UOJFAREfEk4mFfmox3vZIM
0Po8JEPU2RIBsLFJDV6zDHCOL8PU9q4+1dU0O6gYlpTG/vJbY01+X9B+2L1kWy7R
NKrUT43RyQt6Cq0IThjoAHtWw7w2Qj0QnhQzcdMT9A9gEoxtyOquWp3Kwdp/t9+9
eayi7jxTmLk/sG/75jtJcXXrkGJDF+3Y8jDW8yBcNC9RVxG0FLHYu/ys7leQA3tC
WcGhLWgfn5T82x86uxriN5/8/Lt7sqvlVCZvoQEGhS4FV0/rakL7/lAKfmPv+R1N
QVMbbYhdBidF95YRBsCfjppl6Xb2urx7tRro29OWBmg89RoUo2ri82c5SIWFSIec
GBSYCHr/Sfwd2+xqwMxQjYkioxE3Wz9kILnTeVcdiJn31nIVo21OvvlT90/spTLR
Qw2aSl4ta9AXQ+8vyJFwWdSuZnpAbqkO0EYGmf0EimmnKChBz6jwNkYk+oDaH1yE
1mXNdaPInzOo9Yvv/Gsoo7tcEhtuqUWuEj4HpfM46oufZu9rYBoWBTzHQgTviHBq
pfq0jwK7PY+CfS+Q1xy8Top0A65xXz0CGIpWz52mzS86F3er+A7z2osj0Ug/D3ae
eiIhPmJnxxLAV8GLtYEyO1k3PlDliQGLSWZq6eXI6RvY9lwCHC26Plw0H+8p/Gbd
VNUwZYWNn7NIiZirR90aZpgkose3huBdxS0lRN31yIrs6hkS1k+IepGXR2pHXxJ5
/ZpfwF2zvI8+wLT8hVEsYD98qF5dvJUw/dBdwHR12rpbxhedAFjaRLDSsM+uQ1a2
eopFCSSnGiS6TRLwCZTyL4pYctU1NCZhBWg/tskF6G//Sxja9KChEPhzarAfJOto
xGvyOR7SLCDulla632Fho0beIjom+AYIsj5xaRofx0Z4sh/pCM0KQTrPquHBtQ1w
IUTjOYqh2Pi5E7GsEpbSIHvJXP1WrRVcjSKAaGyfqIqtbPikLx9N582OdD/YE8r1
2pljfBct5+sjBmu6/l88d3iX7MrDSEAzevYMkBvAZuW5f/fWnMrr1S7VG3/cTOGD
ADtN4T/E3Uza9wH0pxxJPyeZr3HeTesttYCHzGom7jXxV5RFwUJT79Kn9XofrxYe
CUVmOjBhS94utpDALXvSGm55xkf61UNKTkG3h7Ckv6u3L6Np43rGxvLqkLPYwBs7
FnUXEg0aYLj+lrV+zOjNMuvNIs6SbAclqs7LHBtnQSQiOM0qb5xWawHly6NVaOiB
PJ+7Bb0b3LG4s7NjvSwDdYja/p7z6FxICdZZf0x5kLY6NAczY5Tocrv1D/WwqLtG
rcWbmZEbg638+hFsm/BEJVmALXrCmuIcmy7NNftWURTXdPp90QY9S/oXyPlcu7xf
hzRDNGj7CdcOlidWcVC1HUfkjbxAQhSSgavLiqp0WkjIrXyiUYuw2ofUKLviS/n5
jF3SeJOUwehfgluBOcaT+SQHds+lq5Cd8xiI4R6ErjN1VF64lP3seH0cr86ECu3y
droOD+fANG4PFM2NSqGi9i84obvnejr/Q2m1Mi9fG8AT1WfBoCanYQyuhE8gCOSn
/N8vVHh4IcxvRDMGvOXjkyAKadp1VfoZEVLw07BgJNUgCcWMDkBnr9dtFAaoCAMO
xVcIK67kJv57CwtMgb11Nm30sGav875ZFoCx1eEh6RdShc/KQ+jErAHAVKhPJuVu
U2mEGtId4TvxPizsH1PRWx6zDTytFSKcMGneuXve7lOrtD14TlWEYeMmhIWysSFk
AzaodmxJgOFBWhP30R9J8yVpuYWVIogAMX2FaL3FJO0VDDWlG2+TGKU08haGbcQE
cK3IxaF3G7ZbH9pHvMyPEIbwcUYMRrnqX5xxV+0nBB9ZB+plshAff9VKZW9EIUi7
qlxo8PEB3ut4QtybaEaXVOCA0YYp70xGCeI+TrvD2RxCvDCVmPP1IFtXXPTBsVIM
/qVAgPbQvxTJpySofwvPcp70z61YQFjGMDzRhth5heqklxM7Fab9vfnWT+ia3GAM
4KQyzU4K5ORy7j2Pg3Z3IkdiYYszMZGZWFdDgrqK0MUecuy3JU/inXW3e7dzwO5O
OM+H+9wdzNctlDDGA411gKJCy19I1uzoaeJYOHEtr/5jtcS4buFd9bCF3iSZjQSJ
1S77PW7JrQ/DPFDaH42MCe1DZBWnn5vMNw21u1F3n7vkVefRMu2q3qTs4yenSRB8
NAsjY0cMTnmFU4Hc1Vus6Nh/cV+eiDqvSMYSm22krIysKrJEvn3JZxdoJtWQ/kPv
5uFaqor/4VWiOFJpJdljoWYgR0hv548RkSBV4YtQJ1wAiOCQTOPshOqlbIG/7FqR
JRB1pJYtBeMfgR5dsEgpeDjBkRxo2m7Ao2OuuNVnKzymPFdq3ofvIff5yY/PRS+a
8DZnYfico4xBc6N60Wr/pjADkSzHYpdgxn89p1V5PT48SEc+zsv9TR72SOW7mD2M
kcVVps+jsXO8Vb+Xx7kJ6/gr7++OcSZTZ5D09LY0/ejqhP/IAbdf0iMn/E9pLDe2
XM8FMOH05trYltBelytTpNpoYHE+xjyDzn5YtIpLPZmmAbVPQ9kmfx2OALjuv1qF
1OaHBZ0Bav/a7xzwCNuqoj3Ikhb33mVY2RF/HU7g3dZH4A2ksoZbGkDNfE5LesAp
0PXKKpK1V2x3Er0IlQ7qRIcAAUyKEymple6kCv8V6YXLxYFW27XXTzCw1QcPJoXt
QDWBsviZ2Wnbf1/HiebNmL4fg2CB7oa2K6cIlvd1LQ9IotCbTq1e9rY3ZrZx2Rja
+w1ke5+16fOekEViYbYHBZCyI73cBj+vEozmoISk5MoSu7QQvycrgrM5h1HlRy7Z
QwpkZczw2Pkq84rmVuIPif2ttBjfwFe3ZSjQPHVQrZ+KoPIcyUJ5/T0GtVZa518j
yPMrrjlXsFltTYvAkVixGxpacxkFKvzmBZdRVWSmYVjZ4mScaDLJ0vi+/y6rFh4R
80pYeaQFfiT4/Zh0wR3Zdcr4rUIMRR9PfjQNq3P2ClHl3s/wEjlB05MS+f4vRV1k
qiybd+ONHcckb6a/MkQEAR1WJzmjzBWSUZz28mDwHm74emITub9bHgAyFYIGMDBP
MMiDrlu41qdeTlOO7+7R3DBM618Hg7Yb48Rn9XcNAdcsUFLjDuOaLNhlbuRTunYp
bh5bTwTYtfXHoTXatUpcJ8yL6Fxx0HgBYsh8aKmJV5hpxhmdTNVzebI85SrpXh/6
X2e7TTcLKwbEmgwxJCL6D24JDFzykcDwwCRPdh6e1mSRerVPThE8nivEnIKEurT0
G/LuBNbbdvNbNWD8DC7EqC4mLvj37HubyP2x7LwuzV6FqxkZDN/8GYHLt5cOkA0P
NmyiatCkOIE1lvNKUIBKfbVJpm6dgoj6sJqVjOb/7ONBIh4Qfep+3d0+jTXRLWBe
G9vzhjlDSSJ05IH+5k7KLMQNBNxHHXmiEvvAYNd4Kmag6DjkJyZBpJrkJ9+3H5iH
3GQdagXkL07w8moaPjIuPefBkPRFQVswYo0QMwngTKl/oR7zL/H5yLqOJC/0l594
brQuN7aZju0ZTmD/v2AaL4NK256ZkhnIhyFapwp3PrO/LFV6gVPU21MfZkN/Ei2p
lcLQOoEmdSB9EjSlxypA6hPLrXMIohBT3AI5artYHjqNE9Ba6I3SEl2OXO4walWk
QNDhWCN29+HwHfIz3vc1VHxfj+RtkrvEJp/WkuBIhZI1CJTvslW4CKGTz2cQDYqN
DTDFbadCUqi/nbY3xGdsQ9D3+i7F3A/215ZPAtqDHyxbg3kLQtdNPfZEIZS3nfYW
AkoBIA26r7GXy+WrMdd++kk4fVubCfQMwX+/qz8hFES40en4VKKaBklHctDflZ6n
2cX3lTPNetXIS/WzP5LiatT5mrQsZjMWz8UIquLi/YNiiM+H/mJBPurFmpXgah1v
BE5IdAREd9WlsKXsLweWxkda8dbPJwA6CVGELiX+bFkA7IBeY0elvGdaGWQ0Qwfw
59/DrypROtUK0NcyOp0CyIrfqNqDNvD6f0iMvzbGi1n2J0S741/kzm7H2jRS40Rf
UxlhwhVpRa5w4RohSqaaNyMSWMvZFUjqTJdULhrt/FzSVdOQijrQ1E7aP9mO6eVa
ZQAJJMafIaWNIpw9jcbID/UGPXGs61RQVTvOTq0ufopa+n/o+BDnuPB3JdeezVsd
PBz19h+6WSmT3WaaQSQdWKSw8uN5F6x7Ysy5YZHSRuwaRnDzAHmiSFeAyaXshlQR
6LRV+F23+/rzGKiCzUiQ2RFAF0wLfrQTIo6BYjtcyycAj1Pgqx0AtpBzVeTTiufW
DN4GA0v/JBgR4bOn9jQEDeYLH72EAP4pWEUCPwrYIhem8Kuaup/+NVt/VY/LiBcT
1EAX/uWakCcnZseUsPxA73VjgEUUnS+eMS8tErl4ragFCKx2nXTq5tcephgmznco
BtPjRqWjT7gmrh5PCatzfLe45zD1v0JbCUz6mvjw+GgCTiRMAy+aQs35TeQU0Vvj
n1uP6l8oTwL8OmrAKgVDZ4crcpviQqah8F7v4LidVXdrd0pvx2SFYxEA0s/MK8pf
X9iJ4MfoGfBO+9b2niJMx7dC664O5vUwfg3aUNzBe4U8KXShl2sWp1NtjW5BeWNr
ih6YyPFf4NSacXWK5v3L0JcESWnaf7cyGVU4xEAc4tdHvw98pxqaDGVsCpUbr1Vq
3eaerHPYAInH/PtfAa5f0zyAxOUQqEZVwYJN7Jp1eDGkwGJo5vJMpSUD31BaNP0l
o65gq/Mk2sPE5VacxOI/edN5XIIkARRBFiod6aCmAON6lJR16k8oHjycrTURR0FB
nHjxPRvA32kbNfdUj/cW7y2mBU6++aFcpsB0fGv7t/azIekj/pBNkeMdIZ+d+PF+
MVLdZy5EylVefi6txaJGhfTKPnCJSnRWDx1keyv1S+X37+p8ZnqL2/RJnki0WrZj
1GYndJwBPn6tpZ+rIiVeINWZ8p28aXq+2oENjb3MkzKQW7rq8/kWxi664hl8TJUy
qLc0ol/cla6TNZZ2ieUfESsD+Ssr7LoOosf2vTRwn4KWBo+h1+UyPqVUfnh70RPZ
j6m09TTjCNdGLBMq1GpHxQO7/y79jzpf8jPkTfuFN5YR6nffBbuCqxNBzcSSnGHM
DK9hLmTGd4Occl2l89rz2/2zJs/gfJocDmqge9xO9O59mcrKiajycphWTJPxzG8S
DubSDlkmYqmNgSwT0Ar8kR4CFrUP0DRinvzZ/VIr920kiNXlegbUEXPNMJxlldGc
H7/zYQCl6omo/HIPn8XbiIjXgn6+vS2ujDldr+DL55lAb4ZwITLIe6Pjy/KQ1dtf
magOa7kOTdtWlv2yYO3JMI3T/zH8xSxhaNYXd31iFjphBw0/6Zal/vYx+alq9zu7
56eKdT/uyDjR9/7dxcZqMOzXjI/fuHLf8bOt6vtJOx7GFo3AhXAseRUbqyF3FrBm
w8RDXGVeFLd+1L+4AvxZz9Q/RTp07xqy+jo/ytCJVrFQvyIxsLZbP/eZ4qXvQK47
QnIxYwgj5kee7lZ40JQStcgayXFBVOqu6pLgpi5V8qKL5kr+1rOk7b3/0SyoeXt0
4QcuQNiKLyw73C0kbTN1jrtmX7qQaHKokNK3uBNeECnEACQkQNipGQ3c0Sd8zuBA
rdoyCdDOlyDoGvLz3hcjdp04HA+NEtILXaakO1JyQ8ug2xZb+TXTtLXmnjaM3HXr
zoZu91jPk9usemgAjAgQj15Wve6d7d8sVs5jx3anH+cUhyNN69w7Gm4x3qTiV1iS
gk7aj5iEdZcLmxvtvYJ6h5z/o+5rT4K/hFUDlysdJsbP0VSH1nUHTazCD7L9XGy9
H3ikoAVt0ire44Zc1NiuDlFOhZa3bOlGomm1u55t7fMZkqYdZCaqXcshAnXNfyAi
OS4dKY36tv8qs1h9U/4KdrDOwpSjkwT6v9n4trV31ETlUdq/Q6Fp91NvyHqzavvg
EWbWmvPDh0hKecpPOcz4aRze31vaCry1MTwAxtjPmk7c5woHejcsPw8/VRyezFfe
v9LQkp0MaM5fSFj8JOJWtZiWvl42E9PHUaIf1QUKIxuvpTzw997Kevz6niY0MWD7
+jkKorQv+7NEbn6ffEzoCx39W/UXPfW/OBVh90Ti2Ae9sy/IaJQB0PoFs6mNff1e
HAF3kT3XM++OajpnP4VnHiH3Lv5weTpzWTXWpDb6rwxR/gf+ZlvOBxmypS5rO7jN
xrPT4eHTOidB91mMUbHoXBqHM9KCG3FQfDho1PGUakD3/zfH//Ias52yQiwDlA60
2pNC4DuynYZXqIlEW+0PJuvQBxAq1ocd+TgmJ3oiM2gVpbjM0rjD3zm32r2VmUgk
2mT5WLiS97UIN+W0Mz+oxf5+gTrIgtXLNGVsE7gKMNzulmJdpyfw4aGaf7qJaMO3
RbIoPy/Fuy+WvrKk7mVdFfwS6nAgVNBAa9WdKEd6+6M8JvED3CESSrdPH8clBWiW
+nIr/wbyXNwzllLuReqQt76xGAkeQo4c5C7taqvloPE0Gj/I+dxC+EZ25dd8tEm/
Yj6N87CanFU9mhBLroO3YtWNBy+ZKcD/eYrnYx/71si710HSKB++tgsZ6XqFNzS1
9zu/qQ3qiXSMs8tENCxLf/b+R38P87stM+jG1RbIAnTG461pUe3nvvCc4oEEB6jN
1FAYHbxJCwG+Px2t+djcArA0K76W54/WW6i2Su+f8vl3Fdpm2xP/up6xr6IikOt5
m80hqQhj9Icbgg+VlQUqpLDNlg/lQBqWExJO4Z0ok0H55ga/ZzvjH7GKqjnR3Wix
zKy5AVMS5GuKdmXaOi35cw6VIuSgHikRCwPNEV120NsWlJ+VijeE0OtgUCJeD24N
xp2MAzSZ1wqjTvZrvT0EkSVLhTN3muT3TJkhlqtjzpqq2qjnTenQCtGgZLaJqBiR
n7FcYHaaRz8wWFbvFX+K0Sqw91s0pIh5wtmC47/rSRm3/CiGIpIrpCcQ3Fv5fViA
znsJxjcdSL0cUx3Lq6iiaXKT9hFejbC7f8NXf/nN6MiWcnBMrOIWh97Nd5Z+vY/u
e+bgrNIjdHpcC/1Srla1bR0HBlGfAmWJZn4dZBh0ZyR0/Fooh0lX1WkfqIz5VTX2
0sdyqwzyKtfxxkbLGPKMgmHZHuqPg7Qn/uwiJvBWsdOhikDvA5v33ROCR395Yp0W
WNYV4LEj+e/QWszxjQtPplFNcSM9ckARqj7QWemaFKJAYN6+pXhQivIEubeN1VZ3
Flt78ZGNylpyYru7QyBTljOVxYvMR/h7LGq+6UudP9gQMBAp65aTuN8GjPXVANPa
cZQYLs3W1SN6QaPbyzFshyXk1ovpO6hMuVpSt8Z02OgZPZ18EERgCbJiWG4aiXyJ
EAT9pgekkUGhyvY9mvgIr8m2QJvCiByGcZV/wV5cLkBPMR2QzCncSRmPFM+ZiKA5
dW4TPizKL79dEX+VeQGsU9iCkHXnF8uwhPCMrLXl3/3UrDDe1QNuDVKFZQqU4cwu
G0aR4iZfezKdkv9VRn4rJCjBsT9a7offHwkTP0flUlDlAxTIHdovv8jCko+ZP7nh
7kyspjzpFs761hy0z071hy9WCFoTW3A/QvE5wMFGW4H9SCI9Xus7whfFCnswh1/z
J8T0GqDPmwbClNgRNymIHaTZSq/7zD3Z5iK+aLOPbK7y9CbQDfu4gADWTK6lb6A2
4r3Afcv1EZIFmiq96UMWZnavUTCOHQIyZWJFRx/RkUaxr3oxVUKVSus2UHb89dIS
URqanPIjSrz4xWL9wBC+i5Bifz2RIAFBvsWpJdfl8M7X+y47HZZrKJBOjo0cLbmC
BL0vACOYoYtXMJV/AGmFDUiBpIBzfjS+X9p/OAkc+ovpxrg+4FGSkQJWko768NYd
/i2udr3TxCfMdlU4+YWmhOb+Vyq6YIKCQi7q6EXmZ/aDiHIIvCfGII/ceXmdPIQJ
VxJ9O+lW47DN3N8RxYBNyWoUexqX9HA+2/zUJE/7xzb2SYTxWX2GIn9t535CA3v+
iTVxtS7bxNbpC3r81/DL9+HnRMfd94wkNJfMeY8PWkUog97wbGKuPo5sPENnqjbA
hVYxq01OmHhLu0qFTNJVXZVP8G9kC90nUihAe7Z/Dcs/g/2/UxscQcwiL52D+BFj
+MvrX9QGUI+ojdr+UhfxrXTJH05LE/KSRoSUGjLfUFQNBLLg1ZdNtYo+fGNSjTAJ
GF3TgVe5Yk2n85LATeiRL6YFWHPexRl9+0MJ/BhBxpP3Sur786hi632rFg+YqeOj
sS35rioD3xU6384HvcU5/mU3VtijVUtmkH46MJkrd3ueIN/USxdGYfdrwb9ozDhW
bqxRtQflHNNbk9rP0UaxGQcfL8Qi1wb/TskoxIifrH1dY7iwaZq/RbouW95wfU5Z
vwQGjbdujx8g1Lwd4tZ8HiSY5yIgDGThNNv3NLnca5qrZWs5FMFpr4tERbsPhmCu
Jz1WDty6yXw8a0neuBSyWhJr0kQwxyWu8WnO9kz/esFW5Djtf9ZrF9C+0ytigKGj
VS720Cct6ur3eDB2TsVy2rqxfN3UvzSbK3tZTKo7RK4337bmeHw6OZ01BIZa7Xzh
dGcTOFTN/609MuGwbzCfsJEeVRSaAB7O7l796Yw2+e1agPaVFbTYPm+DcnAn2K6v
Qpndlz4cI9hsl0w5FrkvgvpQ44SjxdWIPdp0czB97+tdMchJ97sdB7ThWLKVIWzs
rtkPo54kCznVn4C7z53KnP5p+mHmzrY6oTYV7l6YvdYkSP9oljCPx5gllIq+nAT1
u3ba9AhAXadPCa+ZXBMUohIWd9jYu7iTjiyqSPBDV3D97CovLlec+9GfoIZU6PxA
JnMIOsYaI15l1d28p5JyklNVsyHUC83Jb9wQqizL4uNUzeH90qOfHMnS/0fAzFQB
QnWSjlsE5p4etMRprJ/R18ix3ZjFugAP4Y2lSIms0HPuwazRrBkwev3OvHMuAnG3
oH/TKay8R3q+It7LkFZFA9+QkSf2PoRRJEXhzfuDHzjOQBvpQjTS84rsjfXnTXph
+kJ5vw/Gz5ZiKLQh9Dt/Ogv3sWkMmPN+IJirryrpWLkk6d34Wetgt4q0ujU37M+I
JIqmh50SV/DA2UxxSRZ/Yet43AXqydNVxHkvuXiZ1xEjr+AP6Mcixt5kwogTskuY
XjDyf7QWiOszqsqT19MOd/gMGerh+yvVxI6lVIJvLvFXn+BbB+T3wizo0OEs1vjy
X5FfmaSAC5TWdsE+ZzOS5UbTkaoL54y95eXqEJgDo+6NEXGZmlI2TGuPguFmgl36
u8Is5uHI+byvbRH4Sjfbi/USg+0aj2z1aigzLuqKoknXsYFNsihgrPm72tQl5ecP
WoGID2NhjjVibx6EUvQ4pMMd54gP0kVlNV2dLmA3UD0Eou215vlVzXT93s5lBPBn
syKLmJ7EkMbbKOQH/dbbU8/mlEPZo3DTbpMWqpU9hTpMIknICa1G81wuD7yZDHUT
nkkzkm2DT0d/XTkqMWYn/mBbIJH2fUH4D1L1oYwdUeB84CGphj+S3Ad8rnJX06ve
gJWY8O7LLbZXjW+1jjE1wCTqu9ZrMf21rSe6Eye8XBNOYRpq44t7rClmQBeKeosN
nFjcHtSMQAXsGhmqw8DeeFq/h7OuSO8kRXfHqJsKbiv4vS1sKnh9pmhtXxSff4E5
j9brIRxtAuSK0WetX8AhxAza6GHYd0C5EBXfTzOoV25EzecKjsRGL8AciNr5dVjC
RllGH39oAv4h/L8eWRSURFPCiYF/YxgueRjhEYWJE89QAeYyOciTNHoWlTtaCDtg
cCTQ4sdpEKRLda307R2ihmPwMwJRKG6yUMsFSy0aVx9PToU45YvSUWoHB7Md1Zx5
F/qM6JgZb7JXpJ0K201y6qbGNcyjsd9wruFrpzcfKAuHOjq1vQK5xzbROYNZJvq0
fnjd7sUtv20LhF2j3tjVcaMYj5qzzdIlyE76/fjUOaCYc3enN2Np3IqkuJHl7Kkv
lP5NUM9QGwct1qtTdqJfw9RGT0ayCxWS722UadnleqEV0drQRhqaEKoMLBWJ1kOb
LchSLLlaoLx9+Mky+WR7qLXukqBx6bEPWOktgiYYycBrvWObr34rWkTeYPZL18Pm
Y4uJmoEb+Wicb4fL30MPHyWR4bQalPf9vu1f1k0L1JTb2zyab/5F8cyCVxWBSMF2
80FUdjhNV6jtgOsZFfmW5UjVw3svq+0zzk7o2lHvv5n6tUSvloJFx5AZiIlRMOl0
B+n9MZF93pJ/FfVwnRnmkmmTSN6bEtTiLhcbS0YwtHOirDFFethCPXJUmMPhrK+D
F/gabJCoAE8M2508XIrGs+6MUtdcdeoM0kwqPAULnuxVjKUDDJI6yjmhIgTCjfjO
R8GtB5XfcgM52I1+B2oZcpj2ncQ1DeUiM6yQZAoUX4JoH5LnpmnNbMBe45FQHoVY
Fzk5aJVTXqBm+o+IAznUEYsM9af+hAl6LB0tjpuR/vZFC1yRaE1qXJ+s10gLs9kY
XelLt6Q3nuBkNzw6ojM4p/8Af03TGHnJfivdkhgNTdzls+rZ26Rvk+nHqCZSd+Yy
0DyjbMBUUOnhdHG1HN75wXCUK+35nCG1w37iN4t45gAIqS9GYCO603BqZcnzzGL5
m7llEddtfKNbF6cy+fiKYE2+be+b4F3wMZBJB31Tzy9havH/BG9JYgP4R97dJQnO
llolIC23hI49oQCwP5vSY9RSqY+47PNzaV5ACsgk3tygoBZ+yY9ns+4m2uHsJYe6
/U+/i6xfm0Cpar2krPZkVgoKxHv07h3DsVupG1hiiLzbwQ6iyz8Jmk0ENonn8z6C
+9j0PYN+uF6I2TG/T9+Zc/1bAHhuNKutNLVChk7jlSqHvrmhhlzWmZsD7n8kUMFQ
+HpHlPxCUVpaCZneu81mK7aH3tQ19Hd7aqpcG0DsipDKQuYuFE2q7D7nP+CCTx7h
k4K1g9O9UrRiiw7UAxSZFTEecjLTufWd0TcKOJ/7dM5rlW3NEDtAlr6UpeJhSBP1
OGkVRQtt3PSYJDss2ljUHx7fhlyoGnX+C7+ZjTvVKISmSv7vca5efdIVtiPlp82C
ibBIJ5s1FX0ad6G9a5AH0hsFkvJ6oT9v1AylcTvT2wuY4BPWsdWZsXd1XDOhQmnr
dIqoIbpUVZLwNZQJD4XV7G6ShyjxNzjLain/eW8uhmaL95f+vTdSV8lnSHKAdYsf
y9mQHeNfRrRVZvenv+L4/AOpfTGqpd9C5mwFAM3lbsBukHDgu1bMGn9yX8uKxIGy
wBG8Bw8Nybk5z++ctvITtfleuuc2ga9umviknCgH+PFOjyb32vzhA1j+vXMf8ES7
EzohPVWZTQUruBBkz5yNgKLKs/95zvkCfYQ8ZE5AEBB3zyU3XAJn64ml7/kw0ES0
OwrsiBwRZnQwmgQSLe3Q16wZhyI08nvnnXFPWlRtV6wfOJ079aZ+xaxVoBBEKOs+
VTio9+7VJZtcGF5uM8HGUr/f1qXzjGqXaXSH86ONBe9q6VOv02JeLgR6/ISq/QAU
bxArbf2gxjzaMqkapd9aZRsgj0sKU17FSd8+sMYQIJbydapJFkSLqcgtVn5ONNt5
oaamjA5DHCxJEFUg2M71VspDi8Ia90QYPDuw6C5Q30cgOvH8Y/aCNQb7xpbtMQh4
IzJG3wD/+QB2SDzJVDqImxTY8BrjFbWJAJndfuxoT9oOX+8Ec6scICjsv+lgbgUp
HePiIR4EjGPCzyP522IopRv9fz0vze4wlyVv5lST1Tb+wz+PqwVVFa5L8JNOyNhq
wRWX/VHhfqCOjz27/x/+yLa7sqsMzIqm8Efu4m4aSmU5XygAIV7w7aDgY7XbJxoR
w6IW/1BsSssW/A48uAVww9ItyjoUs4C9ranYf96POUV92BgT6m5GsTTM10DTy227
FwQnbHw5lAEudTChaE2DFaV14nbh1IrXFLIQuCAgJOENMvHlOnBLRYCfJj9oF/27
871Ef4TMYOZNKIWI3cl2SPY6qRUWccm05jl8nWkfTetpAF5ONOfX8W00w9NKpVTc
BYLSWSKVsDg16IAvrrBJ3D9wluoaI85jiVzPJlcwnkGABBzF4ItpOjBLge5XXtHC
qEC7bYY1S32IZ0FOW2a38RKG3uoVoGM7k8+hMh573lA2oxbiR72upyWNSWL11WaJ
y1h+KxyS1/JCVboGrWLJXJU/swoiD0KNaKn6MFa+aul1GY/3vsitqOFqBjeP2TvA
IPNgM7UHZTtPewGNacixBk4hyp2petNewJczPwm+wElkfonCshYY7qiQcbOgowEI
CX2SF/PC1fl5ECy0odCnqoS7gU/c5zZI1QeGkX9EBnRe1nCLuIh4ZZANF6l0iopT
bHaFX3DLEMwg5pDsWLJzWQgKMU6AzQODMe5I7PGb/iJevOWWkl5yAE07BnakjZ6+
h9pdDKkcz+wZbT1PSaCcIZz1n3fUTKgT37OTWRxcfuyHJBVdv5tb2a9huVi8TFDH
j+TlEGWpnvyARyhb1JQ4YARweLQr4WDVBHc4OS2uRkNwfkgs0CmxPTfjigQmCfBe
GJH69hv4h/a61pNLdLg2vu3NmPT2X+xoUVsLTWFrwJqm4dPYpCiK/ht21jmi84yt
82pTPFlgFk5xT3gkK1Yp0BCAQZsLC3p2D/D6dotuHBO905++iuoa0ObK8kFtbA/Z
OVWk3yzsvF4lwWWMU+/nDp/hNDhgCUu2/8Px6DnlXfrXtY2mxtWpcIgYaAHSBtID
jHZwjAX7oxgHpJihkDxQI0PeLEcN5nOkfy3jwn/TMjXeClVxCifffh/OhvoWUntg
IA9kqACrR6bh+T9MWcS+IjnCjnyC2bF7wiPkcgKMBkkyAXHrrUlJoS+fKgEo4beg
kl7PNgMPcBv94OGw73B0B9sR3Pq+1C87vgbdkRFISbJ/k1V4yeb9bOt3fJWYgcsY
m3Hsw+kqAQzemy8BNnIqtQ2fcYsNppk5DxXgScGKnINtxLqUbHWlqcvvk/DWdkCm
MwMV2LvkFgae5Q7isr9gjGvn4xxOOcKk8rDzYJkCVhGUZDec0mN2QQ2+dhmTKbrh
yaPwxhRRQJcEp0gSE84H/i7l73H57Ylos9HcxwpsdlnwpLGVVXrzATxAUZpCSnnz
J0N1Xujba2dr4LcYQRDE0sPeY8GSNtsk5lWU6S89S5eQRfDZVFPN7+iJmBvruwHR
5pyEd3vG+ClwR7mu8vhvrQpRfT7mLAAtuzWroO4N2BlZabcfA8cQvfB2560Oq38+
ZSS/IIQXnOvBB5YBgdqYqyzKsLoE99ESGRqqLX9qoEI86DJ67kmUHHrdMaUUDIHL
vOnPOZYL5HLhlI+nudfsOrPo3JvbD/PqZgqJoHlBszJfovxQh9wveW9RUyJEFueO
28q3Vzz1DRXMO0WG4+OkKPzvsCxQDf+CpuEGZ+7V6zMtxvWG04WEc4v/OMyZWN7Q
oRTryM9E8OvycOPe9xmTCT34QB9tLKRu4Js4PCUA6f9bZJhlNJXvLgkBlYlpOUJw
ixyhdXBxf8xS89pLJtJYK1j08QCsPwWeYTRQdtXFEvBsMdbRfjsF6EKJdSnV0ipu
fusBIqMqdZ97wCCM/Fm/rhxFTTeyF4wYSDJDZ9gLu5Awxuz7d9WBKY2KgdTMzrDR
K3z30HmlVo+T5gwLM2GTZuh434TfSgPNC57t9/KX6o7lwEFm0Z6WxnmQfHTkZKBF
OSc3JCYhVOs/6KqmgUi4vlB4966faBCFCXTr14+tLwJzB9OOo/FRnzfHN0HBdlNX
DGULf4eAsUoQpPpy7xBkJ0UL/EEX1wS5tGZZI3yhikrEjwdo9KkANc2oXO5ZDMia
4NNeKHqVj4vdVj9qxrblJQedFtOY/aKgTgTKLcQ6AZ94OpkYO/KL+KJuGC3xyFaw
uu9bHkcqsbpMrmXWrzn88LtCg9ZLoRETfbVFjx9XvoNiLVLqJuSaJYKXJdho48UR
BFwXZsWY51+/5gvarGtqHTBdGdZ5cl+EZkxFnkE33xCVY/ZXZ8mIaOW0GdvgVX/c
io7bTojFS76L2vsrDK9bA7mKC3jfASXx+Tl3u73sMGE1qI6magXrktTl6mta5esF
DYGiVqiHOEKSSLqvx7Eov6Hl3DqGHxLix3Gr4nFZ8FdhHEex4N4nz+VXsiiEglUv
QhNpxn9gGUWL8lzLcPGWMj0n3MxsQ6NkM+Ri6VcO1Emsaja2Oh8mzwmLW9qB62Mq
av8xxy+mDnexRJgBTwRpS9ZEMojPjKeP5lGpZ5/S0pzFDZpWkvLTr4KksI+bnGCP
xc1790fEAa/0IUQmOnPCeT9Bwu3rAAimwThANhWsJ+Y1F9ZQEHDn53iHSmTflPyD
AuiOyPWPbl5ZaGjPRgqyS0WP7xkgbKdSViVvX1W9smlXeMH3Dt2VJB/ecqhJmcEt
v/O1uF5KPSZbO6G8U01mZ8OZuYkj1zoqeXdYya/ghZPefT6Fl+j33Jl9unhsjUGi
aftC5oNFDQGXTv5CXqMDULNwHYokAx7KT65Nok3SQ6Yp91GcWYOQVEybT46iGlvz
f9q40S8HxBc05SY5JSTfBrcsGEnYRn/yHsCOiyMxfpPsMOVXSQ6sNZPQfdebm4Lc
VgACLQ8s4AYDqOEYcZGw7rChHlcHSJKEY4OYfwG/+hOP4J+/jjN/i8aKMnCpQ5Zt
e1NlitESKRBz8Dd5p7zWOvZZlgbwgphdlTyBK+gOKA6lok6BNHnkDSXf6Fzl8nPT
C/S78iEjkdIBomWYxW0NYC39MelefwCPHd0X4oqkL76egHDMA+CRhR1to/GosAor
KMyyYYTPE8d+6ECLodmgFtoTx8XLKeSwd9Frttji50AfxxdKVpAV/uOj7v6OraBO
TauUNk//yG+xYAM5EKcI2MAJ+mUYPz8z4Oh9BSj0f/XaQTpUhA4UfccMCNyJ4wbJ
HqhRHu+5Vvgbcpa88icQ2811Tk1bvCRLkF8bRIgcDBetV1kjEqoqes51E8oHkaK0
y9FB9iB3k+7cle5bzDYImkm/TV4m4Lrhs56WerN4ycJySgZDNaDD/lvuSs/h9x6b
L1PNfVifG0YIp2PmWPogDdXmTeZddEM9VptQ/u0ndSzwpIASGOgF0DWvptQ8v+2b
eqOPsOo43j9DmRcGsaZNWP1L6IrL+N0EYYdr308Aa3mYNkTEvMY40TP29w/7GzKX
b5mSQIlfHui31z2YseK70qcjSLp4+iIAsctrWx5zckAJozr9rs33h/ciYjLwc8wG
AwTpPJRJLLHk5MD9heOWH6aJkEvIs8BirnGYHULekK8ZDVmnZdJQ+S2dwBgZ791y
PuGGSQqb0aRr6Bom54qcNUBlqrRyeJ5Rq9pMq7YzLHvovIkwghdl5KqrM6KFiQtv
W8V3Gs0GAVEqm+d0AT5C9EyBFxcIQ/nHSJWZozVWoAzSiGv/aXOUzVBRlE3cPFsE
YVMNRZC5M7hyrI6aBzG0IVeabY++90sgiRYMC3om9WIdKHu65eJpxYgjAJ0rThiG
FFNrBz2UHTUmf4U0s6XvY5dUuvHlsmlhYjDtciWiwcdjGXlWLV/pLUS8yRYXPgcW
9M3zP0mvDX7xv4739mFXSKA0L2TGhr/g6LomCrMArhgAMXDccp9PvvMfYl5O4beG
tZxEZDUzryfYclrWnvzYlXRyFqJk7JaMLIlsVnWDb3wS8ev+QF65yrMBzhvq3ApI
Y+2i/vYgKtPGyc4QSGgv8MG6xVYW1xZ+4DiMslcAfPc9+ls0en45zbbtnE0dbJOM
1TNju8EH3mCiCMPWpAOpCD/xWAQLl28Hp8T0Sj6/tzBWl9RlMc4Ocr7BY1/B13Yz
RyRlHxLHtZTPnwmijN+bOtyN0bS8lCubdBM7onPql+tJtaLJs7L1Ql8gYdu3biXe
3UUET56ZXRBEtCLi5I1tfwY88eQNK0yDZN32MlwjlWdw+Fgwn7zp4Je3DLr8JAcL
MnXLW52rzICNjlaXBQfWIKCwnecXlzZAzdMP5xhBY2y9XfQkUdBa/seSPvYkKcRh
+QMoWL+GTkXRH5SH28S1H4bkyIOS/l2elVi1oPmruw9YBMyggxUtIrELm99EVPE3
Efdl8u+7ypU0g3XpFOoJigUgdevnrzjLb6W27Ugnk2/mhUuUFhRO9kqA/tVvNPIT
gHam/rSxK+0axydzfIX4akDC5yAPbpE77I4YEgvXYJNOhjlfrEC6i9sRWu+Wvjx8
INSyhIzSSpK97dFUtMHoBDcQz04D4EP96LBU4yN+xwpnKnmhNopYL8gmvcVNvwyr
+Ef3NUcUXDOa6FmMgJ1tpKy7Yx5y9pbkNIrYZ++88wZf6z5FUPQI+h1ZKbCBS2/Z
YOPlrtnCXCWV2zUB7KKdC5D6lxXdQJN2XhlhV1+Pi58na9btHOfTkWk8WUSeZXFO
FJVUcoiXTJodeE4GCU63hjmfQSBsaj7eOg15uQ38IoW4eHONy/FOrWH++FiUgAio
0yCsvY1M7NZGuT2uKK1RdtfXKJgBKRr8xjY/P6+cvfuvFCX26olMq1AnqYkw0X0Z
BJc05MLXAUsv0WUrc70EhK+q3PDDnmmOR4l42cUdw/TJsUU1ECZdxvVZDMeH3NlN
cqwvMOHivrBtg+QyI9JTM5vLSPFat6NV6cGPvdsmDBwdqTS+cD21KqA04TvDzRex
pD/pqtpJpv+Aed6Gte99dNZEp5q5RBBhDf5sSB8W1f9nyjy1sLs6X6Dki16dlVLS
H8AdW8ocsXsj2/yWWdaPipcc28zrJ5dihHJNH4Nq/qYJTQ59cXT7jCAYX/d6Gag2
Qm5xTbiBUMz9B+m1azHR+j/Ky9HVyAZXqZnX5Y4Ij6EquaSlA/RaXT9EggjfB/0+
E2+bDOcXVfhRIA1rLNJ3nHZLc+LR5AECpo8Ol1+spSxZnGxMB0gIRVDygo2rFb8M
E/30ea0JqX2757joRMJoR12cB3CojalLC0xEAP2KboKVXKent2Vj8qEJDI6+djSw
nEUJAEN/TE1Y9xJy1hF28FroOP3bTcXp1D8FRa+8gCytjEzTzjiYDSUKVyzuyYFQ
7sFI1v+rPFKbgvrrDIrXuhdaS48fHuX+4r7qvK9eIvGE/cpG3vrhobeGpUfDy0+4
fojolMyZqkOKXy+5OXVrJp7p0/XLXX4xBo2/BlEYTkc5P+b72ZlMhAL21/qk721w
uBC5N7hncEyxtpBj4zAhqcMEoDZlHURivuj7cC16cHxrRfuLD4HXKQxxsHEjkU0Z
Z9tA9QBR8plbItjNlzMXS4kfDqlRbAkItoLGYel4huLqoIba1dH1e5Zhd/Yq8/cH
QLpkFCJ9Y878t5UpsYctbnRXoOq+lYIPbLYkLPhxKGC8rTqqQ610uTLL2zYVVj7+
HdyIJW7AC2krRvBmsBO/JhnzNSdyKrXZP08Nt/+lqJdA8YXq23HWO+aIrbcww21C
Man4+biBLVsWfiK1eoHhXZBRxw+XWNXEGo8XQS5X5UCJ2iqxmNbXSvHOLSJTNaDD
JeTx43NP6+uskVQ998Za7liAxGSBgsf+YboIJkisl98gB4cNMqUplPTSp1i+yls+
/v+raqQkLWiOzyYlavDUKvV3efzeLSu8io7sK7Cv63TSD+hJ5N2fHQEo8S4xNLys
gIPc7qJtFbmIX1wRY5LKWz71pcuWgjhkdZkh+2CJjT0+PxteqBQk4lIZcu9B4WxS
5oV3DGwDp2qTSyd7VTTtY/e1rYGDiH8UacUUdGN0Oa9UGmAQeB5ZWUwvrDPaJad0
lQ78EQH+JBIuCfVAfRgGgSTuajkMbKpDpt+9/oTK4+EiOI9GnLZe671I0O6Mw9lL
jQOx2YbVjtG3SPr2EuGmUc84q7M3+EzBi1LlGCPBJaS6saYYFqJGzAewAHp0Duso
tefS3of8rOfc6EAv3LQXQ7OstY2WFtzJnQd1DmVNPc1BkNOagMmlYhycgxTf2vk6
nTvb4zNVgMIVjpb/qX42ptIWYTXIx4XYLwcDlenzCMi2j4bNNjxic1eeyztAyj4u
PP0g6BWTyfZurW7LP/EQDx6tKPuoy6d8B3TFkczuHh2i39dwXF5TDFoBaGY1Nw4z
EDe6uu7l6lJYnHPv9D+BKYwcd/bZVhh3DT3J9TPUIgddneV8gKbY8F9gumJrhgId
WSjwiQUkMIIibQZfR+UZYHMOmHAX+LoynDHj0AIALiZgNDp1pSaSpgIt3bGVltXZ
lG4kMPUN15o30a6h/JoOOUfUQfvthChnzaKZ8e8jXySxrjnHsGb2dvWCQ26j/3HI
8MBA2A3hVA2/QUEg6yvprnlFrzD2vfOr7bWQ8a+RuMDIjf0R3RbM/hVuDx3mFKuU
dPrHll7U3vb8uA9xupWzkImtgSS8BumePI2a9xqpECptt9or6Q62LNnOz68ILTeE
WzXjbCvg2h83YWsGdGTstuhwZkwBJkyGVPMRC/OEuKizyvPCUu/MSaqRfTxuAO0I
tH8xXx2UG33RM/LyKJiLsHvuGvOfwzCWOBOyl/hhsLdRYZuBInHDtfwNcC1MZRmb
gzjCpxOnpU3p0xDVKZtQRt3cxt6cE3pACsCtK/1zei+rAe2Uf8OQCwmFVvwR4bgq
8QCkh7EHap8eoCsJp+S2dgWPgKJDCwEDk65e+9XyH0Mq81/a+00Thdq5fcKhl84w
8iTW0BIkJhFWPPZxwWjN//h4lEf8rvHiAUZubJyyscNLU0BM7tYTHg4J9b1uqx5R
ypmKrmjgV0NmqYqLSQqiCQfV7JfeCQBoEvXVM4FWSLZ4wiSbo3jmXXKIRt18rBs3
Rt0tkmgHg0aZHwtpupwas1QlZ7osLLKAi7tu2lpzfpkhvuknPwEu8uuTMf/QvUB0
qyeKvyZ9cKFPbI8wPv0A9gPDaty2+OBr14wfeNl2YiKOHYRJagHmQzz+ym0fZeMr
fgqUHlRmCIb5MKePjk+XgUnmJvl8osvWjz1SZ2p25PNHiUTnGEl4gSJFebScn2P5
25qgGi2XRWVzT2y9x55fLtKFOG16GZ4YC4+eApoWeb0jbsY+Ic9+RCK8YtDx7jkt
W99XrzKxEo//3ZdJmtS1Mnr48rOZgQ/FHwIHpzWIHV2iIpDGOY1WTz/+QV/WmKsd
5HbuoQEL4wNafWs27oQIqkXpy+5/i6TRPdz2501S0Ajqxex5wbn1l1grTOFbkgjd
9R6lGA3izv0kl9pbAuC7jtfi0O/dcMq6ixtfqoro7GqfDpQ7NEwyroNKuL++Gh/v
zQslz4C60E1otNlo7M1kaScixCzwywJw3lEgrv20tNk/WMJaCmXyv01q4UKJy1LW
SADPRxHVKWOBFUnI1mVmbGDUZV27Pfg4akjgMsTi/ns5Bww5CU90e8eGZIqcNJZu
PJaRGtvPPbrO5q20LTc1UeRlL17bSnSxf8yhcDWeTMUqMHCP+GEo+3Us+vmm5G0L
Ly4qnIVdxdhPsGa4IiPomwle4YzyR+kViY7yEP8rO0+2CLY0PhUHhxA3PPZOMKxx
grmtG5+3sYoKlzcBBeYi/WLEAcow3oUNoAxaWhVpEdpT42MxnD8DeeTWRXa5Ensl
TEKJi3g1EnO7gHi8TNcyxgCrkV8f8Qp6ZLLzEOIH9czEeLBkP3aMbnR8Now3WAnK
oAm6NBHIbbD4P1abwanJKyp4c47tzvHGHwFzQaPcAfWhGzKxcb5CprcGnzx5K4Uq
zcnIzPKohOnUO0iGtx0f6IbarS86dCT/2DWMi52OXKPRA7rYlLggOClnFmWw4QUM
ngtJ8TOc/bbBjkL2zMYPwE5yQrJbzC4prxyoXNg1TxD0jpCLtmVkeJHc4d/QmslQ
iZtnRZUwntvuy3aiPQ3q0Rw3wk0Xm6Hp4hO3zAVUjMpWiyOTxn2Bt/Z6y2twQMpw
/4YxKZsnJVHOZUyDBEtXT2u7+xU/rmK0+9MIPzwHjrehfqc7o0X6E6j3PMCMl1aS
skbxL44EEQeHCWF730WBZ3iOJeYeagMSsjsbwv74hh9xxAFNfOSDelhz++j48IRO
fCaEMd8kvPx3mGT2vuQK5CzhOb/UlCTMXpJrc4hL23yDZZ/4ihVnR+/f5vTVLdrU
x8roWmegIbeLLY4NnZaYK96PkaeyEbEcSqbI+fjQLwLylLFNpuHZu0H4gT2N/UXQ
+zp0yXoRYS4T2sO0Nd3pKAz/TbdlnLaz8OFKyj6AaawCUnCe6xRhMKwPkJ+GXr4V
corTZzGYZgz6lp195LvrL5IJMihOiaBMjwwgMmqxTZ2xhfW70Qo038ST5iqkYL9m
SkSm/iZrIfayjQx+Jtrkf97kpNQXXFSFxaSkXAodH1vFbqWqfoVHxvbjhIIqz/rN
EsU5Ovk/qAgdK1O9StGamGXyiepnB1/dRbdHfUe9ldHaxlhxy7j6omsoxjIiKgzI
8m2m77PmWTbsscHZhBJ72nEi6FJAX9YUDCl7Xu+e2xrCbPl3++Yp6B3HPt+cabVl
Te40DDTs85j9lyIzUUb9NxDwNnfAy1HneOadCyWyMbgBja8t1FeOR2JTvcmic96G
jhHz1/wuOummk4QKAOuXpxLCS2Udstblu40lGaMO7CeWKOIqUhZVZVPylEqkqew/
GFe6qPALPAleYifK5syy4KOrfx9vfbCiSzVFyCW7aolfQlkW2YLy4+t9gYSoybex
gPZsUT5YrxfHyF5eWB3q7Rz2CLWINm2hBzpipAV9Vh+bPR00NbT1nQ+2bFdnX4M2
QNoHoRIjMao+s1NvXkIAtkel0/C9YWHZYqEMqIaOBrc8afi0FgWPaK2XMx8Divuo
FQLdrmQazxMcmDgAfNnYRSe0QM+2eIh5rJFrLUReCsgGi5Fd2f3myi2HhK1Mregm
n9dxjOZG01LNDiODlbtOSX4IXrNbAd+nccnoHxuGrwAfRVij+KjLG6EiX253pqPF
Ks+T8WIt0mu67Dbd/xgLaMYpb5Z6QiGcZaUQyc3qWhneF8ylMRDISIDhLVzTXD76
fsXTDPCITs4kx0gGfJJtzYNCQaBpMnBpqhNTXHQFPZl7Y/ivXgoqQJWPk3MC5pao
CZtbWWJtEff4KqnQMMJDIPdbBJfl9giFQP6sENXn6eB1MY1c6tPpEVJku9nU7AEK
D/f2EkY0AKxOQoKWardYbgQAhLh+If0X/7RyS7qBRr9BbGmYEnNxt5wZnzXOnbel
zN4tJEE/Q60AX2mpkKy6JYbbMuCtwhB7IrtvATdp9Dz+EVgyzmVldZntquqxB5b0
jkvtsc8a4ojmhI4LF65jnYpoeRQNS+HqNuY8ypOHLV07jhfIaARw1dbCiJCOvkwA
bJ7QCchskM6Ac4+OhKEt4aeLSl0YsVTHDZzfYhvo5D9HIZjKgjA5pg15lg2Fodwf
6dJSm+sBx5MD6c29/ged1/TCMwU4dLqfWkfHrvTtCStRg8bed+teHFKcOvhWqoeU
FvodU19pyX08w6hwe+5jPMoV8PDEalXCwb6cKF7VpvGWc0xM1GjX1bkC8nxPOKZa
KaD57MmjoeiowqIS69ngvuyLx3XfQt5ZE1KcLOp1rPU4dhNCMHQQ9VCE55++66Wg
o8J1rSKOBBnYROWIqb9+cUMbXriX3JF6JiCSWt/bdCTeZl3EPlQUdAnWOlsc/HdS
UTxmrHkHdiSZM36nlElmIZNep40WcehVrSV4L++ouVz60qDo0rSOud6nsSJkaIm+
NOg4REt9P7XF8ibPJhO/V0lJzZ16j29+f+pNJFFcUzHX4SKczfXpK4F/rn2wWA67
8MfM/ZTwx8JNlgmvX8dL/brRiumaYtIpGALKvYaVAeBUU6RgF8c6ZByqmk4yC+Yu
Pn00S6SNJkCIZXo23WRWmr1WufDWpx789ysdKuSuHnEeIW7q5wtMoxnHDh8NnOtU
U5t1DemQgI2a5Pscp7D67d5RUjVwP8E/0AM5jrNqQJRC7UGWUr2jaSN8jXklaUNz
sErSlTf0mWMQqv5ccXbr2AycXxQJjJDyQ+uAQ5XLXFIB8dXl9kfT09qtXAFUPg5N
4freSdz/72JR64SLDSLmFfU4+ll4KLP/CB/sARUEFLZ0hlm1W/Aimaijp1cfM65a
E2swbVjD64VUpasCGmQjvy2XeArV+SJfpVLH3NGvUKER35NXqhX5ehNHnrVWv75M
/N7tL3dZ8C1EnT7PxqNpDvyTUdq9mZRVvkr4PkbhsKXkXcUr2cL91eCYscPVbhNw
V+2wFLMbI4r7wSqAW2C2zXyeAU8DQ93hEVFToYMiPlq3XKzMCKI4k379CpjcUgEK
FXcH/QJthaSjDyZ4AGlBakmRQnhSc4DlUWO8KjUhpRxcpRSVVJbKCkEePERddXEH
HvaXpYKaaxrEal8mn8JSF3cOo6fQDPv7J/Dr67wMKJLghn/JocgidY79BDv/Xo1x
eAENlMeHjt6P1Bg1+tcobORHDzlZnk+lJ24nyUEaK8riircqV2PY8mboZWgyCkWs
gov5pq3EIC6DdJfosCOE6bOjLFkyrUSWoSChXoAhJB6+Z7ix9U1+Yzrs4jaLY6C8
iK4KFDfpCjPv5iW3TUO/lMJa0GAJcEdEc2H8Kn3nhzEsoMG68iaYxuCqLQkNN9KO
jrfd1HjHnAht7s54IP5oiw2zoWWYJfSo2bDjc1Jh7oeX5qIn6lPACGIgJzb19Bkb
Kf2GsHPYKDwYJoj1WD7x3uAIi6Q1VEyFiyPw4bEQoSJh7ue4uiaV7f+9fJYZGvgf
a47WLdrxpoMrD4j5YS9RpPZInH/RdN0gyZeCKytLPcZCALOcYXCnhWhJ349wYcaD
WBZrJYBSGPepEXCvHoLPACXE6QLeKIN0tGLbz0eLElH26xf0l6khoM5o+j6YVPlb
kIY/TRIHJ5aXtMVcJ9k3lCXu52o6qtCa9ZMbdvsixkgRrwoCa24y/kW/1FSgCWpO
ZF0cRnwqxw7Xtc0ev4sbI1s3hJLaoRG19/3IbgpYQ9Qq8ssOhXGS8HyEKalOeHWO
zt2aWDCKZV7I4D0EpZIEmGDOP8ujzkYeFHPhJoNp5Xcc67F4111Zt07juJrgzuLX
FK8/zLMbr2NWFzeY0ww4Ibs/HEa88ib41FHT9hbHNlq6liAiypxCMoyQ99DGDeg6
h3IeEBIoi70d6R7lvqkdtz1zu+Cimho0IwTcan9PzYTNECLNzR1AIqCmSc+FzjlG
Bj1h9ebw8+8DIYV9UnVgxsUNXx2OFtsEQ7yncQGtdXYBh7bhnuh+jvk4J5d3TeHQ
1rPpXcwX5tSPRV7DaAQJE0ub42+P1uPXbYwCO7S3ZXHDnb1IovZWl8lIVDZRTBLU
SAvpixFE+ZsUnQ9ilFFczsEQizj6Zwx+OecgTTvoiIkuxoZNHQ6wyQcvilq2/eaP
F1xOG9yGnaeHYWVI3ZpSjEY+AzJEGGdY0nr7U4+BTkzYeamMER39zXrmgTH2G4GV
qj8OAhqeKVQGn8YmCSSwHu7nAmORSiCugX1vIbzAivzMHN6D+mO+JXhk7C6MRl8p
58bfulUznrSke91xP56GZKcXCaMltfn/5lFFlM0qMBNj7XRXJVKmVQgojsxP/agG
D3IF7oJllM+EH4qzNcdiYmHXFNVJZrKwihJufk1Tim3fYHtmCXy2SdRA95+pGQiC
auW/49AiqfChbp/eEe0WKR+B2/Uavmf8Vb5uMNezx+bukn11ohSutOx6KdlVIe4D
6ElnZL6G+osd2YsezqThbO8LvmC0LfpQrwElnxZJPbXrPOAjFwXVxULlSHsvyRLO
QziM8HYkPcCA/TFOemx4K8UFLr77C75SdFxtxS0uQy+gJCKyj74un028FEa+9e9q
sA8wDODgp7ra4rfpieTSHJMCMjOzzYZUovBMgigk1hVTrCYnHhKcCPgnzP387aVz
31WnOoGM1177nqHqlar9OFrFpfwE7ocdFVdI4LWY7J/5eLxoOr0kXrE+W9SXGqs3
LqZC2jq2zpA3FeVIj3txEWBZrUUGdwHIu/KKQpmP68WzZvCn4cwDnYykGcE+WGoH
urlXnruUUa32JG+RXau9eW8T66u0Js4cQ0Mw3FBjQAHGOmPiZ84kqyY8HYzNevL5
JMgD75EF+AxQk2cg6YN/LJuT0QAb/ctymrKLeG8/x7/DU0+RxzBGR1Dj6YQ5OKK3
YMV8W0ZD4X1h/455CaregultyPBgBgFSCWT/B/ld/lCVcJlEWg2gRraH6byJ6U6l
JEh2DBocbVPo9PQmnE/5VdOG87/06c3j1CeyhwttXg787GhTp0gKqnCF4yTXYYX+
cp2O2uzljUe2n7iGw3c0NTx6wnsrVBVXkK+jLqAn5Q2ArnqQm4+1l82bdLGdeKhH
pYc8fE5yQgs/vUkRaRF9eSsM/RAxV9cxkjti4Wqs/5gBiKd9f/YA+nESKi0rvdj5
zhluBL82gSjcrCC0JEEO28FGWV8LxTdOEPeyyebGVGQZGJUKbI0sstUYKdKjl8Ye
fqvPU6yGKAi5ClsMOnRt9MoylFICF3yOv9UCC21aFaGMVJ+fKm25sk2bHI+1s0AS
h3cMalViOwZMi+VxrZIHlABv0/vDBVH8VbG09fltdHk98bsWfNBAf41Q2VdvSdew
KV3ZznJViLbaI8c5EzaFuA4RmAX7xk2dJMIsx4CiR+T4kZU9rf3AdvxN6qnjCs2q
Mb6QIEn0XYkEvzWSqsyjnjuHfwTK3Bpk1q51Ii77wDF5Cdl0pVZfHOeCud67Jq6P
EOeWRptQsy78PV6pYm0ZwNkOMqiGKH0RQ4eqhwr4+TJvSdHsl31TZ8fNIxA8MWfE
J3wnmeDjgMpCW++IXE8p1b/EunuyhEQf0F4KIOhJEF/AVj0ROtwt0rZyki2IlcKb
g4bZCnlBFA3he/Oegs9bN1XWYqLZe+q+ZzJdSqfm1vE9NMg2aoabukEz0Rf9RILj
0nnfXglyOsNkWZVZzHzPDnUD3dQ7YsGlo9PahNM2S5SEOiwjWofwieS0ydHWpdrM
BZ8ErVs1jNJqqs2HhNFoJI7zl0H4MO4G6TGwq9s9PtEdN8+reTs+4Nyu+P1qaQCX
8Uxby7ZJLGOJ9JqSn6fTKHJKnQEzPfBnvo/hhfDzMBMvSoIp4NdGbyVG5iaan33Q
bbnEGO54RImY2WGyi25pWdJmlojUSlwbCtTBbVp5iK3I+KcXcKK/ux2SBGZ2RPlO
MSVK35lKx0QioACWmAyCP2DXjCCWGaDWIm0M2FLztGPz8imqEXoWzQbie25RYCHz
XEgKLLEpw5j4w9OOWxxRT+fTQqKXb9WI2SjSE8Z6RjyuihsI6yrZ2K6ZTUNj0GGv
yqIuOQIXhYQcWh5UvThQzQMd0omEH63opcs3wCbLxrEF77ZOX09XynolKEDsxaNK
hiYOBpPPLcY/LAFPC9fK8nYdb3FSyzlMbo+OsSAAWOK/y2bamgoqbVjjIm8fZDtF
iZ9Dv99UOlaR3/3LVWVUSIuYewsSV4Fi6yD72kFrFWBa8x8Hez4S/ZquNzw2NpBp
VKZyrTz3/S5vvDE3grBMQmftYayrZNyuvdR/yJHPet3X1VycFgAC00k8qSvcfAic
9dUwhAL44Zkfz8ZJlvNci/P78ffgH2esfXs7qM6Pksus009MFD1/Q/RZZ7GhuqaE
uwTJ0lK+ogauiW7W5GysUvLp0kLL0c0dPgFYbAFpmqofzkh7bRnKeGeukkoljDjZ
hQ07aD+M6N7ZWdOPj/y2JJ5SjJobTRlA+EhTirZcLcJfP5HznCws+jnlHPnV9Sgn
xfzJozXT17Wn/jPSQXjIXs/Mcb8dSqf8gBFEU3EpiLZcYGjuiZeaBmtzEvYLNYRG
tOaO/ikuekMetCJv2mKSR5AJ3DSpxEOp0DbFU6ZxuOZSVlF4wH26uuydaTN10t9F
dsFlgod7+bnOc9uTC+RYJvAYIvHziWFBYMWTOaWPmM4NGFgsSmbMK496ofI23tSl
SqtV7Onq+SFjkfxrX19rjQ31cJ4sEeeDucUVxsCpCTOwI25KEZ2/qlGWOF7d6+yY
xFet9UYupjp1Qx4P8JsALfDcT8MTsZryAMd1+OJdP08DPWKyb/OEIdzEIMeE5cTW
ENBj45JRAP0khD32+VkviAGa4jYfPNN/oDxLRi3eWxm2WRgyPqWv+ylpCPMxJy+I
0x9HthfIaauXmHViAU8joRw5QbLH0OP1rTFD3i7E9KYaEKa2p8P3zXSub56PYaVY
53adWJC/1CAbNs+p3usJBY3TPWmyO9hnZzzWfz0tOgGJLXHuQJUON5n5KDvp1BFM
P/Je/PCBh8LZ3ezo/zzKOW0hisVXCpHf3Izh41RajLGk6uDC4UOjS4zcvk18wmit
5oX076j4HhqMuGlI0UnUVImP+Xmxr8eQLthz65W5GdR62p4voQf8Ig8Vcx+zExan
q+EjSIyRVCyVMvFUqlaQT9pSP458LVeMKlQC+wsNmJIhQSEUDqO+fMLe++EXcfG9
oeNP62kbpTDxt+Cc+3kv4NVc1Y+DbJgF4hORrYrqxOR0JHJz4oIjne9sNN6Pb4ks
YMjeH+qnFIWnIBbxaQFKCZCkXRGHVAknDjFCqBq0SKpKcBF4Kv/DOmfaXACVOvOF
+GOQIKZA9ThXNXDNDtB7cNro5uiwfL2Z1Mt3oGumOEMyNxfFcz65hHUZ9k4Yf/Wn
+/hjrQKKwzUNmJvs+VROIllmNfMiBv9qQJPVeJOrAEIskGPAlzj9VVCEXTjMIDCr
v671tEt7ZDEkKom/7VIxENSNl2+YUEyIPJBkfnxNVRxdo4GGHJnGUPvrXPXQp+J8
n1182vHZ0B0xbjm5raHJjxtrsIrpbCrsSVqThvi6GmBye9T5fZzPVSxUQOdP3WCV
z0LUgcteL1++J5LxO5aMyCr0w6yXGyjwBNpO7zGrIPw+AWqhnpuNzd/wY00nF/UE
qtdkyJV0qJ6uJIYLajODgN2fv6MBgEzKUUo1/CGkICdljYk7W8AXS6OLz9xkWvJB
uW54XemYqxtIKjhhPY5tlnU8VDFq79y8jRg4zd2BE/4lolUwb7XzrcgXC14RnDky
QseKq0suLMqZ80ZBvBs/mPkkQXA0lU+79bu2esu0i1e4lq+xwOkx1WMFsjbmA+27
gxs03Cp3C9wVcAyrm5S3oK80yMHJdBIj29W4i7E3DLKaLbMNThYOwqxNsJLK4AF7
f7hk7sUGMBbeuTw8/KsGHdiw+5SlaM2CsSBPqnmgmMisUhSgheku6RO92pQXsB9d
cNnKBdsS3utTVw5V0yrdXTvCm1hTVN//OkOThJ1zWzU1e7dGkFefuyZ5Eb62vnL6
SW6kBrDwy5zyad+AAQZPk3MAxzPlwoISINO4tOzYLyF9KRJqGER40WCBVHdsB6+b
7B2O8L6beovnCINLdG6Y/fQfj3/Fq08XMcb5oZmiSp0D8RE9dA8mn1h+/Bo1QSG5
vTlfK3nxkC6s0uY7kedX6eeesziBMOlZCAGu4nciqaALXkKan0/xVwDqA/2EvJRC
gcZu/6WpST+s52SQqMp4GM1MEPmAmtwMUI1x9JuhC6K132pzDExUUlu3Oiy6bU2S
BzjLFnH6Z4UUrZMjlYUzVDH6cqvoU0B+85HBu7NHnPjNrUYSKnFaBGQVIghezyx6
nhvtVoHNC3Asawa/K+xHUnsClxZNtAkHNXVxFEzcBOScVR7jV0Tzdvcucb+KfgCf
t0UhDxWrN5AHEwrFDlcde2fjyJUp44OsQ8o/vWK6Yb9/oZ1n0zIPSL6AqyW6gi2P
dPcZcdXxfPtEpBTGQoqa5mckkEK4N3gFL6ZR7v+0lU5HYp528cxX7QQ6k9pX/du8
JzrhX1Bib303zGP8tOKwgbuL4ZrysvRHvkNiEA1rNp6nO1Za4iIxu+QwaZHP56BM
OxHkAPy+YKMTv2j6/6/wrPh8nqDpT+X7UwyjCT1ld7wKPNq+LFuM3jVvMPy72a29
3307u1cRwUBE1UkdNDRfqmfSoHPgD7/l7284VQQERuFDcfXOjoxjPRQ8oefDAwzx
xlGavzduR4xiYXckxnPIgdZ1E2Rd84u1UMoizO+XqmDb61am1lv0/sOnl8nXc6K8
DA6S6CzmQVVLsv63g6/fYp9M8y9idHM2aAXdPlaWNsEduJLqOF6htSQCoWOwnWaO
P5J7Z6PAMUGhVkSoIM/J7ohY7Mw0xNpyzC1ye6It9j6q+vZhXuMTn3mhG3hRyVZH
bSUS1EL9aBibn8BL1FYlt5ygihQ/WwqN14Bps5uoOx+akwvxVKqLVexQNc0no7Xx
mIaCUZtxe/p5mQcHjaGLmPXffPhfBH2D1aTAfZq9EIQO0mJ1nYO+Ok81boMSKGrt
Qi41+lE9o/QSWWHSJW2o/jeZNwgK+HL05u+C0iqKvSfmCeUEK/h0blfCsV7DMpen
ipxyHsSrsqGF6WsklqZfpxUr1jqJeLho/fNeI4VKcIQVCXZh1xD33oi9l88x1Uhy
jnV6YnOqp47QZ+Vvk+wLvvqn0UTddQaf9Tfv6nx7zUbuQQNzsRmJ8j9UusEglMsO
+upYoET5HE2M74FDEd05l+buRPDNiLVv7egBV4Fwn16iw+4buZTDLY3qkvlMro1M
8qRJwAw13cy8Dn+CHv9kjw==
`pragma protect end_protected
