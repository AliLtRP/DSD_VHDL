// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BUvsOCMkfruU0HMViCZ4eqiW7XVx+opsWJ6awFGII+b3qY4v+8+N/PkR5hvySDxz
Ye5byi/2df+4Eu1DByaBzv8r1qoVN6XYsmeSD1UDWp7Yn5RgntzvQ8+1SpNX1Sfq
uFNkTcjzOiA1l7wRJrrBquCeHI6nc0jv6yU2WZJUAyk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5616)
bCmFgu5W/cPapBp5ZnledJx9hp9NNOh5msa4MrO3koOwNx2ThwixvOJLMnjizjkT
RDG/hjF4IyhDaSonDLpd2BgO+eelikpMHXKbf62e2DR+nWfKvKvEiqrrb5Tp2Srh
LMZgVraV8fnt6QNKn2hN3iAhX9BAfP6QzfQPNxUOfSc2pHRbbdW3FNta0fZDfgKX
iV2DTLrY06/HZPVO82tzT0Fd2gUFpqfbix43vbYWO0xD0oZxsiFU0ig/XRc+cKa5
HGmwexc9sS4pMLptvvyreuuWANtmj15U+e1nRQHKsdGmlLXh2JkNQAMymzFHMskL
UUDTCs9ZsPlrDzAKL3vmqIHvoOcrElZwCB/esul29KHC5f/qSbN7398HxwZ3A8gg
Bm+st0XdeAGUN7+Fpdx4+is/kiJZPw/Xb0ei9tVckSZXMK+sc6frf8HrdT3mlbCO
SjbikJeTDwbSLSmi9XQ7R5ZpyGb9ZgsHgOWsPdRbvwkvSoiFfslqERo8butmNP6w
WBmHAZot0EJNraKsO9+uL8y6d4Xrv6g0nhohFeY4ZojfI4EO4shx9B+YGZo2NyAb
C0IP9DlGhgW4TU4DfEQMD8RIdY2Fqf0OzbwTShIkvfaovO6BU8oArkdVVDik3HZ8
muIW3Au109/oQFWgs7HbqdbVUc785ypxnTw3keDdvMFTwhCHQaQW01bU55viQOk5
69AzUH8483fGD62nn7gK1K/Wfr4zZJ6/E+Db/zP/vq02zJAxOBRzDF7CVpyGTsPN
+v2rSCek1rYDhCqZx9lnfmKWHKqIpTVLqX89n1sdJIg/y6g7K7BXTa8EhfXmkl1L
F7lIQ6gMGySQ4/CPZ/7whzrLF1Y96WtgjrudDgZw5ZdSFRqYicaqR6uGlLHVS2DH
el0qPUHTE+GQtSqu1zEcGRPkSjlZ/uoKbx0DLJOSdsL0ukqY3JD+HI2PD0XmU9Oa
TWv5jIFKQm76A0PrESHsE5hTfqa+6qfht4Q6zEv920Kb7Q5wCR4hSttQjHWnF+BX
rJNiXEtQ9XtJnJ0wJ/wpp+RL4cd+ZfvP2yLyYYw0uWtPOQEQhASMq8QTukschjEY
EDzQgqfVtiYXmxeVEeM1js2yFEXa0vDvpE72plCPuebfsSEeqaPA0lHSnvOhUD7W
2BiEkld7NaYPRontfIfQN/ZaKWCAZ3xBhSCI02FChkyjl7WYpM8LbbdVAtSKpE4k
PSgXrDwUn597SOIdtEmAyGnRaakaF8zGaJLf+YKX7c8l0s2RBjvR1I6l9h3T0zCs
tpw+ClKOPN4FOraGALahHDx5aMfFre8voh1/cf0IPNrVM8MxUaOKcftWxU64vNnc
TKfhFAWziJOocl/htcR2HVbffzrvqurCdsYUBvs012EfUWUyQtnL+883G6xOWE2C
zQP/FElh+V1BTgNoVlJ7g7RWAE/C5HQSzu44qpQ+d4/1DTV1ssF/hK+OQPEpvITf
j4i0qMRFdyd5Zywm62yMx1PZhygRSfb0cYsioCZYoXc1KF9ElNYVaYI8Zq+mp13f
yOioGZv9UF0LjV9ZcGMbn+zvEhxpGN2r++q+vtLncJ3we2W4dzY2zdFmrEgeUrre
x/b+dI/9ZlW0il6qb1twzsg9zWzynUzRxlk9BApr6uq2t3q4oAJa5Q99QGyoItm2
dvalq/TJzOrreJ5hX1NR6XjrWri41ZI5UKxZkP16jxFVh/bs83CC/x5ZwOf5zNHE
KYRvW1kmwwTqPYDTeNtPdyzVYN+0CNm4m4Nls0yI5v/nTNA5MJwRNky/+NacwXAF
WNtTH11BxcUdJLjAsKpuFLcZ7YAQY8ksj9s5172EcRXjUI9dMoYS0KlgyLM/HjTW
v/dj0g/Ph/GLrwdR2u8zEYESgt5X0aMoBzX+U4/KNzWONW2/AzIzRVyrOCc1CDOW
7jXSLv+OWTLLlvN4KO/jDTmBN08JcElJGAdagxVZwL36T4b3M1+jcZvP7un21MmX
TWlTggDWW+aqiUGAbbC7DhW9zEUabkVERWhC6Dr4GCDKkh8Q1tI6nqtfXecU8H7R
pX72HCVYCEblO3LEuLKcMP+BQHU+OL8S0O1RXWEuHerrlGX1iYzsOXNRUW85GOK0
wWI3C6D+PephHxr6Y/hT6fTNl8wjlY+4fGeMXmdF8QvCnGwVWheUIhMa/EjHz0Lv
gx4yuV+vMrE2W5Njk/7RlHpFS1t3r1YHsqGT7P3kfvNxlCtDjmFjQOT3vorbKuP8
0QvGWUSA6lUsp2xbrTsLiwJrMZS1K+dWSPmhnXA9NnguQx6cQz9htWrNogVpp+Q8
ABnQky/0hPPCpWH85cfzukHqjHICVm9wnPl+Sf6e+xxFol527Wem3NcxS84YnqeU
B3t9WIvzlBbKMrvZAHb4uSn2/8yCi5W2dC04zl+ibRSisGAXQGwsKoTeDLR0IDsp
LU4y+3DAB5LMPFibQweS5g4iIR4dc3vu3MCFBd4IyMNWD0nGFCGNcRd1cUvhRgJP
gmxmxkYrljgEwxgJM19g2lfOWYQ7lJ9W/tQbqGVAUOUd+BQv+Su0c/DzknnAwfpr
NJtVIa+Ake6aMNgtpUrtnZG6QoiuyYe8G27gItOnszqTCUFkZzAnI8zoEH0XhvTa
oR4DHsyfjEZSMSFT1TNKXLYdG5E4FL6vN9J52AvgP+WsRARVKiu7zFWpatiNd5f/
/b//nysSBOuO5CalnhkRpxHbAg2mO1G77vQgqvZAj48w7qyFDKdCKUedhsIv0UmF
TL6ErNt/SCHzyU7N7GJ4pKwzeSe+mLtXuf9kk1K/9XAeYIn5NFMtcamBFy9OI8if
dam+rbRvczx1admvGjI5A/nwEbFQZ9YICH0iwD4+bRuP7UVhaf1SNNalLHETkP41
O2e1dLTEOWM3gggoZ+RignX/sQkx3E8QT+ca+9/QEKvPCeH4gyLgq4D9emqkQFQZ
AnnPmlj8Bo3itijSVRGHOuDlAsaJUVj71376H6F5WF24hYyb/reHKrLArhv+uNxB
0GlSo+M5HSzEVSP0EUNZf0z245JfDN4TdnzPWAd/ACARijEjUXOT3fBzrKRAFNr4
ar4E7d8RxSaE5bWY4/tS43zRmtSR1/4u/acE0ReflchsJrp9GNEImqjwrSiOqKiT
kyAYcGj9mx5hsdYkZeQ8RbKuUhK7VZrejE11QXEU3xFzM5TS9+hpx77db+wjMYgG
kKgfpjFr7TrI1TNT9xWBYG5LAkvDsyvgHaMJ9GRQbOesdfExHZs8WH3uwkgGIqPX
ouT1XtthmsDkaJ38h7VAwUkLlM6nawMt7C9kuxmHNIfHyLY/qLiHXBY7BvWz6zZ/
SWWjdrMcigVrec8kOsS+0Xs75MpBHRM3tshioNT+2GGEg1xKgkw1bQEL5f25o8zG
nS7wxlpqsVvnxUFj9KoKlWC3WtmK8RGSheruWjS2K6U7txQnaikDvutB+nQGV/3E
OH0gbA2RsV23+YRrHoCrHTuwYgrHVIyadEd4Y8yCSQNIQoUyqi0efqOvef7mJk8j
nz3lN/Sghq6hFuF5239W2RVhNz7z4MBkc3+O1IxhLFsnkwyoh1EWEE3hu4CU51mT
hQLVR2dlVA97t6TfVFh+XLC78iE7kDygba5qYTyFLgbhLGEEJp9psmyCEG6sLOM+
+hHnZkKtNX0kHy8BbXqN5v6vYisz0XBu3VCOHp2hny50nEHuZKFLwihi96YrFkEL
/JDzN5dT1k9QeJqRbs+1Hd977KaX2OdHaBc0SkTDX4NzPFsMnyoSgXt1mPSKOQvG
efN1p/nEvVcsJYq0wK1Vp102/yuWPT22cwyGspqTig7PuV/1NkVFhHHZjVHvGUUN
LHqiYATdWfABl0pjeiTVIVD00foh94DLcGod6gxEUkSVOL4BKIQk3BqBbf8MSkRP
OuysUmwfJMl5Cs3Dx2DKg7cw/A5H2XYBv/uN0mFBN0A75fUtWGXj8E85cuco/Al5
Q/VsE5hrCXNK//I+lddtnXTRrIDtZeFXvYISge1vZZsPb/OAHluqaIOPW/+09VAq
3rqzGY+crGt4Q7PFagbLHN3ZrUaDfdNj0FDRl6+/EKn3jcapamdxMGvOrCC8iNAE
fcezafSWaxFq55CkwGICdpHLu7TeJ4TDtDDC2eyzfLuaP2FsUEmZlKg4C9ko3rTj
/0MAyq8X+E6SnZsgIH4LDZ8Afu0BainYDwVkQQqALgHfPhd/q55AjUw8Vbe+AlqJ
PLhi1aPHveS/N85HkqRUwjBB2Z5uj04jl/QeVQAa1CNEXLLqk0XVQmjonpcIMawy
ymI46zY/KOJVF7MkLoEaOBpXYk0pakoxFUN5X9BEg5JrAqi2b+DPODoyob7Laj6E
Czomu9j8ST+ctqZ68jhyAirjUp9O5svN6YSUu6g3LKQShiQouW27nm1U+jQ8QB6o
qXGnUS2ffkN4ScBRplCDKuG/O0fdpM3yWiPlAI7AKOPfJ7WuuT5OoRZTjm7guG6P
caMiCIrGhbIxYyPHXQnJEgYVobJBF8XuZA6wO0Yp3mg2ZU28i5Y+4n2b+fiqkdkE
W4RaKS0CWQFrvho9GtkVfhPxASIIqlDuCoNAnH3ua/DwPS/xAClnLKvqVt6xPNsU
ouuVBagfwnF3Z4++yjIvzxl5+0BbGCaimMZanMiby6SP0UKaW00VYC15qsuDdQAL
yg3689w8b6RvIuXBtn8AtDgWyNMjlev61TjmaxfHzKkbC2diMx/pq2P9RypiUFGK
byBCHCIbUg40MSZDUabQNujvOYV1vb93sSvVboaGVTat1sctsAQOZTNUfnysIbGo
6ucKSgcGtoKlANAlCP7PtxkzJQnYc0HSYuYaoTHVQrBqDLV6XRPFcFZuETaq7i6c
wUZVS6vNjo5/9u2Flpa+XikTIrY7uUKxZZBGZqhS3MmywMoWQQixrDdtFUunMCNx
qKlZaxxAZc5ewvoYHdBKFjWGxgv2zTXzvexDkFtsSOTLTpKxCgR8oTQYePnb73eU
+RwMc87VkiMRuV6NsIvH5dPY8NufWX60UvKfCEXWJygSh/Kg2hu9N4LyEk19Hy3i
RNTTGVIjZrUmMW4NpouRm5d10XPZGrEuMhCZtLyR3jAPtx3K+KPsSAeBYloPiqOn
6Ma6pGXGeBG9KbTvRcebwEiBfCucqkGcva+EQaLr/QM+VQVtV0R3hcjJxdBsHA8a
N2F0NBm6OdkBmB4W8fmRsSACCrofDes01AEF4MRQxA2ALgaUBmPtGHFD5EQ67qK4
85IVP6YuYOnYU13XgNW7Yh9Dn+h6BQsq1AfhhGr/n8ZIzPaE/qv+ghRpKvpAEm48
16ZjPyiyqsmC7CHBFpk6tbu3WLE5SZv32/Fwk7Af5ur02YlWaBW2QxZURKqW8A/t
TOuOnju4jOuBfRiDH1VBRkFX6deUmEsfEuO4PusQguOfVbXNqFrBGya7365P2csK
Xuk4xO+6YtoAZ3ojCuLKqyX6y6o5ez696DPe2tRsrOBxayzDBut134koZeSM94cy
zOVSNa4Gh3k5c6Uf5cN4LWkK2GwCM97uMZN4tA1t1rml3DbfDZ7tXAqHUugaFjIg
xmjkkGXGpTMTPXiOqEnCyihNGdyy9xpSQnFmBAD3q1nsFyWwZjEiP2hIrv9vw+mJ
sdVeUB/1VDGS+vFz4B8GT/QNtCloBLA4+70OqDcYczEdphpvCr+QLNkCcJUcQB1U
oBlati6c8PbG6EDC/qBK8c4NMS3nUjlPgrZvZSFfzxU8Xmo/Lg4UXeC7Hhax7HgE
xLVoOCVxkTYAhDNecpw9QEhzhn4cN+BqcCz+CfJ00nULyQx8RpPNLf7ie4tPIT2N
PO3oyTceafj6b+Bxmaed0wK8fNXxOsdxb9X0HB8Lgi6VuSRTamEkagtwXxSJEH0Q
//da2mCK6NADmZs9oxtzyG9v+ztSvz1XjZoGDh5oIC3MYQpOtZAbZdgApVuS08X6
e3hPtlR0Hw+Fwgc4c2F/y1/jjcWJgKXxTQ6zpvN2APexmTSSYweJfA0LI//TodQB
rUBNPy48Igw6kxMJQY43MIJNQ9MVVS6RFcvTvC7KIpiwdN6GgYkH+TGcyG/eY8oh
kjZujNyBlmAQUyCnmNwPJvnBIwMGB2pu8hjbTTDl5J/mHAjRiSfLj3Xsk5H3qAot
DlTk4u0fsaYLCDYOzYeVY64Lnaw8iB4xUkPLlGJQP1oBhQceh+fk8F6oPL91E+rp
0gHKSFIqxkeZlU0qqbE3YVziLPmHUMXEKu9BJiNw4ZyS3BUUm1meGqnKcy+tm1c9
DOF1eLPQ2wUYVL6zlIbm5+GDLBf0xE+7ru4NuR/O/z5ee9vH/hBN2cFDL1ZGXwqm
r6PJbXHaPKFZVC7GMnNIg7OjuAFBcgwXn/VVfhGFGXyxKMLszzbYNmIJCUzzMF4S
PXZ7c6dHAfsw2jSPUPWiAIAwFDMirUhluroOUWtnc372LJ16mOIKENN9W9L88BB9
mWDFzolYdNCuDNPdQMd+Z5mhhBgg4pO/dJTLsEGT78kYJR26CJWbnXOsONaPF1Xr
TCAVLs8sOhjpXZuMzNQ3/kUwptvkOFa/GdmZ8siNhL7+8Ge2kfAMrMIbswVIQ3Jy
EAHA6HghR57c3t23K/tbLwxc7WOTVOVbRX6VnM+ILsMryhCM8ef3bcFf7PILn13p
tm9SaEfPDhSFXsRd87y9CWEPBHpKvJIhdlAz1NMQHqMDcZsu+0YmLUOV9pkZEwVF
JnnywT0qgVvzExwyR8MCL+8OO24Csk95U07UkyY61BYyu/7yW/EHC9nWV9WbU3FG
SUmXR3gCFzgJ3zEyZM0xVPfB2g63nH5JeI9XhkOUs/CNvICCYCJLkTv1gSVaZP3u
Qg3bhCftTdMNykFRGJ5SEV9CRlmctvEBvHaR/2vfLICVew+YV+csMGkDF/8EpVG8
cV6aDtSMjHS1Bi8zLhHUrD1Z8sZ8lPxXBESRDJqXczw6oUC7YW2Yfpyyn7hOlvr6
wB/UX754O+BSf5FE85gFvWoD0rOYl+VBwJEFlpsdT2P2FysqPJqKM7b4+LBaLFPp
d3fImS+YAQPOPZ/f3NjFmuJjmzn1QEfZaMi0QW4UAxmLntRjsJ6lGZwrkc7V+KsT
sNaSzZq40BKzkT4gHydqFIoCeSfctpE7tEFWNEC84QcD2shk1vLMJksothuvLJaj
kuW2FeClGCxBgQwNC4LI0O3KQ7Ap/oYF0B58JPhpNhT8NjZET6ly+sfgKbWhpFOf
qpQNg9UPGaFtOm92EMjZBEJnMSnUvQ4Vrew9JiM5TwBtTouwMQ+bNIO0JKVHV8V/
wrk4tqR9+rRRh7HAikrrChCCkJ2w0wBUHcERUPVnX1LzKN8H7ATPbvOJSDsu9Sfq
jBQg5Xylb5i3SMyvfJkRgKJtM+weqCOgIx2jfdYIxdc5Lyg9NTNeg/vtIdyyYS+O
L6zPLPigBuk4jx2HJMY9isTy/i4stRw9JjteSucfCf6CGX9PrHjOmrDvMuGzEk1D
`pragma protect end_protected
