// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
YL9BJTPCW9gTVpE95DNsemeIv2j6bzW+ufrNtUcdEtuKM7pXImb6wCgw0ciq9w2SqIEadp1jlRF7
lSP+QaKAjtmerrQQ8XApLFc7t9HEzEyeawN78DvBFu5o5VX9JfRQEgd+yU9RVUDqUN43SNiInF/b
2MieSpvarL7i2eyeqxjc+FPjbautUIs0burHqlGJXP4mmODvfa1Jvzq7Jqc+7dRAXA9mn57GyKw+
hAFyFpHqbu+yQWbng1t+oEigNauq36EQPhTttKawILSnDNP46qU3N7SYD4D2W+/432S+dGRy/M+H
7/nbAudHVZtMYa/g2nMUrQul4a4t641Io3wZhw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
RqG/rFyZp933UfAYTAYKRrO5VTCHOsCeARi/LA/DoSNgEgC9SuBWZyFeoWY0yR6AlJQGPu57nJdG
gLdm2xBubMDd3oV88yoLoaTuekNtCDIYcSyHbD+d/ewv0YCuAA+ThTkhxCtIPvbI/ZK0LApmwPxb
A4QekciWzm0EEsOXw3u+gUvzozuygjybd7k5vt9xojefmBU4BSHJGuj9MrgOeXk1fdPxt9Gdx4WM
B/iXdg2kHDZZYTcDD2lEcVvzisFBx5sDTXMrUllPimREH7c39GhmY47Jfx7Re/1N2Iq40Xetc2iH
VoAXwhkexgzRJkz7n7xFqvaS8cBWEbUZ70ckheiIly0MTc13jK3JLXutqbQLFEA9scbDxWz8mO9o
Cb5agifjWp03xudCL9WKKXnsz3eIwKLkSaFoDKbHVKdD147+vE67qqqa573djd91qcqa0kxafcUP
A+ARUjjNQtvm7Ic1YPTWdjaxwnvVtaWanUhbmQAMoImInmEYc0RGWGkuEHy3kgywW9yhSmM0T9SH
BFrRfF1180ipG/6AhnvE5vK0ZKhaxoIeWkpkEtcBN6H7Ubin0e3p+/T9o9g8ipIaibpEkrpC9k/w
qZyWu1mhGeiqKvK2J202/pzeQ56QEd67ZldQM+Mvhr5H6EC2uaDN8G2tJcK3YlWHp6CsFfw2aAlI
KuxtfoTXV7fUBzzF6VackEpkPGZ8h+VO5opaHEAdz3Aa5WSXdltPeKrD9WIPQjRHTTeJD37PPE1Y
sqdpgRvaeru4glE0CJt9KN8L1HEyCMfEDUyOlSl64c82MPsyOk6/A2CbsNfioaJBLdk1RyrhdKIF
pFvmkZS38XFt29zSTQ0/IEDp2mGo1HhtF7t+3zCxZ2OfaUPmUg2pFK0KY1phn+7at+xyZP4ZjQ0g
G6+0dmVVJvq0WipbEYa+E3x5ub6uxJppfa0LgL+GX2/EJ9KknPk8g41kCQg6Bflp2/onQFECdCkR
sNh1mFALXxtHIfpscGTcx9DY8yQ5hGI46kZVSlt2FPrtM2qrgV6UDjE7U0hVWPQmvGVwlY7xQSC5
ZkYyN6M5e1ehWZQ2LgXgdvmePHatufZ5prqA3VnENQ5AzNYEJpt2HO2BnlwLcRce4hMryE0mpFeH
ZV+es7fxx4EHXfVRB6dycULIClhOaxdoOQN1OSo8DTvAa41KzvossZMB8oF6Avncb5gZjK6B+fpS
bF5vjdW+V3rdc4BnswSwdLSXpeLCBxsKTbZZSxcHkIRNosz17MnzIgJ6mNLo00WQ+MWJmp1I35p+
bKKtrhzlCkNtnSUoRtpS4dm1SdOi6ZN9jdWCubhzP3XU6RLWq5Zipjho26OkqrJF4ZJKBncr2n6q
tDvQfA3DxmlHHL9KbrNWckpZ/b3FSQemnSEVcyCQqiqtLoTPF24KBK9oDcFidqplQIWub7h/ltHe
eaTp6Vner0JI7rmvX9/5A3b/Qz5OPrYnQyCSfB1rGoGfbK3cp7NFB6On6UUn0CRS4l768wvU3jZI
wVtAIE5k+DcrXr9sKqqhwHTCqoWq6ok970ncYIvE1nmyxjiRbTjeKqSRa4Q8je/zzg/LxcriPcos
GaE7CS3kOH8XrSWj7rLclj4DQY9sXoZKnhEB7xBt9bSGATnCbDuxBxIM46gmBDZ/ZCniU/W8vv62
39cayK2jbXShE5pcb37WW6r5mTCL/a4parjxBwkPjI0pBbijNumpMuk1cTMbXNIP8Dmv8Rc4hv93
VcCl3FgeX+jBsv8vJOj4Y1JWLd3DYetkz9Rj/RQJMTCrbNMq0sQe7aqMTRUnmyV11olSAqtox+08
6GnEdkXw1nLmpjpbH+dz+cQuuPSaVqcay01d1sSADBi7m4OC8h4CpUHk/OEqFjJ+BTgFrKqWHVix
OIcAYsvmvhPLDGVyahokZLj154bDrHfC51qxWq8lwWulz0Nq4mAjHfvdw038Vj0M13f6lZRCCpgV
c55M0u+zH0QmG8wZi01bWeCE+kulbwnePbkeu8dDqt0X7DjuKupcTSwNdANh9ul4cGnklk4flJJR
cwVlkUSIyaC40LajIIGufVXoytZwekvK5sPe3Ur3CoujJeLgQBDMtdQx0LrujhkS2KSXqDSBxOUQ
pQkJOShjHonnkBF4FjlQvUtu1q60XWo5UjQUKDC7pz8Qa5pGWjyMm1FvaC3dyum02QY6xtcdosd4
lQwawvlSNa+bvEZPnX0GvcVEAKeJAJy1hQMLjq6jvWGdHTwayany4WMoS826pZqYjkUw/ZBPof6Q
AMHgu3WWr+VFrNhReibK4kiZQUvDn9bhq6dKNX/mZNSywhtJZcGZ+WtBLD+YnMCZ9E/8kvfZeHU+
ZTHZ0E0G4/GgUj2gdAHi9xW36KvwtTXcr3ZWEDZIJnZhug2YEaf+Bijg4XVD1xbB9QHYLoAB/oet
L78zWCIXAvB/m4LnCA5L44SkXB9xoizm4sQRAR74QdwEiLnVhbMZtBvCY92i8FrMOjMwWjm9eqT0
a+ehtfWAQmZbtZXO4CpQj5yZFNFSNJjYg9hBoEZeyrMMJBUd0pldpITZ4fpArqgXedClAgkBNEbR
aRtMzIVTHhAojk+ZOhLyJ09x0fzWyebItoGrO6LbmiosKI0vktN2OyKwsfIZ1gCzIe3j52kGrWZe
4R27bgbwfDVLGTFGk37HQnCb5r48Tozoxq7b1WQ9fffOn9LP6XA7SrH+IwMdG03kz5fqI9HtohHz
Fvpgj/pz44dgUo1iePQfksHwBViQ26tL82l2g9GWy67KNImdr7qi83hdKmPzQjAA54x0a6VkJvoG
auM/ynFKdTjhH/P5uCuWxsukVGKleIY/nDjngLA1ziX3+LU5AS3UOPhqBhThk7FrKaNY0GjNrvTb
zLfJ+fTqI1O55m6RGc+ed4H8QxOgb2VI/7+tSf24132Zbz7zIv6uo17YmCjRJ9Xl582laMg/Ivtf
xxZR7ICY0ny1kwXamVuNREOTRWGLRTpwMex4uA+QxVdjURBIMdALZmvFSDewwU/wR7IfWdTfg5Da
jFa13YBFVdxTSsvzSvIXOg5gk4sIrp3Jr09upB/0Gxu65y9zKP5OyCpVSTG9x03f7CFldssvrdHf
nsf69DbZBMhfNynFuTPizGi2EY+0yXN3mL5XKF5uMHXgv136/FZMQiGwdkl/w/t3RnVVl7LqteZN
VxwEBpUBUMxUlVwR0KbVC7RiSb5JTF1Jxir5e9ZBikTIhm1EJ92McVgNVXkZPlHYVX/PrbVs27n/
j3mG2pf4cCsFxHShApYQ48cf4QDtr0oQh/Y3OwFZaEfk2WkF4172pb6uv8bgIDFXYpaXWT7PAMnR
kD2+4F4bKMtR3cvN6DxLEbediMB2sQ8ZSr5FTk4xwyqXkjJWB5z3In1Ka7JgctGvz74mOBbVnE0S
vwZXPRW0H2fG2o0z+Jd7hlJipRM2p7qz4q8ZYr7YC5N1PwyktPsHZr2j3w/qBkfNqifQWrlFZPJE
afcFUVlgGpas/pnnlFQqfrsYp/38fvackpZJQkisml3kUVeO4IjzpBeEqaEijZUSEWqWyvATLrHm
3j4xsNx5/UdP9IlFndZO9ERy4qaOXRBSV0yjTbuDXnZYmf4xkl64pMwQdGudoFSBIj0/HGJnhUjG
UxqbwZKg7nEg2me3F7jO7FX4ZuS8Wd5nSRs2pPTTrKbWzS/nhi0/a8jhkG1Wcf+PGcOljYFuZl/E
wZF2+bShkI6pGYCtH3RKH+sV4RgDdip/fVmOgKXsT52oCajd4PFRIucChZAwCTOxksWErGzjvh29
1ngZ50GOI4IhBiWwPxHk1Y8ZbTGXJz2Fu1nFPwaNF9JK8ycE4NubmEHhOXO20jWnIchIjaCZVKFy
Dz16Uoo0WFgvgpuCixYHzcQ8CAbEmOBSoHD0FLuPU0eBlZLYg0EZswP3ZBox6abFhM4pF4F9WeKa
fAb65nUabANsGL4PrS56CcoUGGtEgUwGUtiPctYKQ5sO53zvjBXY8Y0L+Me0u+3I40LkfhSs031F
qqBYLXMMMoP1kSv+tPqEOwf1kddylnKLQ9VFmNqNOIFvH3/k2Oon2HKqmqSU6qtih01lD8fAOcp7
PVqbkhl3Zjk4djhlG4cr0RTWZbczHNttOgtMZoMqCX/hTgAOTCo+ur0qHeL/pGMSrxvKHC/JcEu7
L9ooL1cXbRdiQxNZZkTm1JDdt0qFuCBASOSHmbMkqJCjRSrqxHbB3GsXceS7Hz+OL+ZLVaOkFX0w
MPBLfGH/rUAnOrQeZXHMsMf4FkxITcG3V7HqW/20BMM5fmAN545OHhakiWi5+7zWlyK/YL8hLGqc
1h2UdrcRiRFLXrLCMxq5rrqLDPhNv5uZzjCNJw0NAB4f5B0i7EVHSaO04q8Do0iqTzcsu8bHVCoW
wHO6VxHCesPSqtsb8np7Ua2Wkb9B+f9zk3cV8PTycIEYpvSwtZQaEydP0hTxk+wIX19TbNNBx8XA
wj8CR+br8Rbxw/NWU9yDBhJ3wH1Y/Ns/TcCDEaiyY2pODuzahGe9mKgubD8UHQd3Lq7H6MbDRHNm
XBFcZmwOSSWbLzWZ4i5RjUvwEbxm03eFBTo6zk8hAstjMclII1QiBnivLNRRu5vlTqb/OgZeHHIu
UzqKphZAY9OHDPiwnZyi9/I0w4K5xFu8jJf7GT7O184yZYIwkgTCl3eK149DS5oFSGV0R5HjvW87
7WHwW2b6elwwL/gTzPiQQrfV8i1gWqKr3IUsyv2h1PPVeDH5GNSs944GYxZrtsyYRJdvGmXxgWn5
44Q8B4XbVaKKpYLFfGL8+AnJRh9JNNcl+h0wXmoDkqPRYP2HUQfODLVDHi4fk4PVkGtNSMDrnE1E
GbvAjfJ9r3MiIfSUUsOX/B/Q987rGJin6ncvCTf1E7w2I1LBXZ6PDeFAKiXkmvDOudp/K//tOTr1
/hiYTg5CSzm59JuO3P+FW4NjOQL8JzQTkjI/preDee3bmiX18UQ3tXxzTFVw96F5uSPDmMVPtrwp
+BEf8VE5HXtU6dPzg8nV3BXJo/0ZWbMDVcn5cegV0Bng3+3qDBtcECohtkOiyk9haUFEXmYBdK8e
cZi7S82ODDY1vAbtbkAUiX49tFnvrfIVpwsBDunNv/ocsS4pJzcKUpZW9OcDxP3f15RvBmx/FcYR
ja+XLgf0y4M3z7JydyepsoYketa347FF6CAZ3Dg48KpI6gogGXgadedIs2BjYEyJgjWYvs9x9DPM
m7P4vmifA97WKOVr0n5kXwPmzmGODFmOxDyRHH+Ot1gtae+tMdwta4n/1iF7YlByAwCBtc9rp66U
gp7UTdTM7cZh08/Uhl5bpRgS7wFBWQFtayP1atfXbNYBSPrDPtZhx9wRPhz1eAOmMB0+uyWEm8oR
FVRYj0ZdyOodxCdAdVICQKQpnB/mctJ1g/rPsG/A4/EoV03bAv7UDw70Me894HKToP8zWVD0yhxp
q8qs5FwaMw2hB00qGD3syxxpoK0oC1+2t7Att3QcFFCF+67CD5CzL4Rt4TuWV+ySt3ljUdCGpidi
DuYLRyWaM1qBZRn4HgoNM2FaU0ze9cSP1srSqi95iD6iV8CD9wxwVTjfk87IiVyp7p+IkjeYQqs4
if9/ShJsJ/vh7TQOVKq61bo1rauJz2p1A4jQG4JYvIwtoi3vmhkw6bX7lECLWgYfhCefGcKTV+FD
v8jYU2YHdBRx4NYHGC8EEgfVqLcijI89eiK1QHo8mKZmf6cr7hQH+WdXGJlzyMtM1aF8iwEI+Oln
ihIefRf/1mCVOSwq5rYeoi1NpIJTMtSpdK6rUQO4Rfgsx/U0vXPNg1n3P63Lp6o1sVie32d2QPog
7eYSmBNj34JkOWVNIuHORD9GjFwaybMIQZ6LapkiyQlTl+g55jZubfnXxsgcSucBlXZ0/INxtASb
NgSorijEIaGTTuIaGRnAPIvP9IFzXMgWPu9z7fUm4KKeSK0u3rkiMgb2C5gvtAfGOwBzroScvs8R
RN//pMq/8SDHfvBVwVqyHFRyzhXtF4j774Qf58RkAQ/OPUADC893ltcnr4o1gLzjgYvWd8csxacC
HbMagz0zq2CdcSkkLcSd8KQxlpil4k0ovmzurL7xhY9ETJ1HVNwylNtgV9iA45bJNy8wxQQUJJ/M
iXdVxr9n+LwzlLGNjuoa04f3HRvpOAg2I+uyZI6XuXSAPIRrOK/4e+/9FacZnSX7PdmyaMiuqx/b
0h6Av0VRnrNprYOzJ+UdXn0f+Kem7ag6TPIm3eXqe/zzyjtsvCP0bJwRbAxjdLaX1KjQ4kkm0d62
Y97DmbJKn2KVrfcdskkbRXgoCar56K7Dl3EAhNGsUoBzwMGL4kOa6UO2XtTATCg/UgpOyFyre1/6
jXyqlCUAb+ICNmgvG6U4Zp2gNBjo8nDnmYbtp2lxa9ipLKiFNzomertpfDUYV5IZmEQ2LvmxoQRe
LQNHnFCx+GhcWMlilIzL7xQkroY3yeZWtZI1b5tsgSsDCgX+7Mev07Q4Vs0Tv2HVjiIdm5bELWTp
u9RrYNldA04AzZd9hiJvsO/AhLna1SPB1Y3nh1KWgBz5lw1PQFTvf0VbQUjYsb0rcZ5XOCEl1613
E/WR1gUejkDlGdOa34lPuiObJ/77OjqbOBPTI+u7267Z3tSzyihATHJycjL7LzhTp/XjZ1/KXrr2
ANdFIZwg2JMcljTQoEJ0YspxQM3R92fcqIIbcWkrsEp08oc+CtalwMCN/C5CqLly/Wq9tQRpwEXt
NZzq5JR939y3pjNUaN5aWTIK5jj/lioc2/oTQ9AEidL3FgcTISU/4fqeRMb0YeObDuDYoT4PJNEb
YSQgbIq8nrPgJEE/cDZheI8dlwb4oXaFK9aahrHnjzRK9ub3qRzSiMN1yLUce7hrWFNzgTGr+qMd
wSUq6WNoycDXNmsjM6AZLhtU5cBt8AazQUmgIhVdJxmaORcFqiARt483CEwV8Z8Pf6XeP7dVWFKY
fwmdEryCuFwwOsVWlKevB+gTH2BOPnFvkB/DlfhYbWFCmBgNYwe14GPeTp5Oj1Qj0GMzLEA4ea8F
CxvqR/ho5s+2YBiQOnXTq3iioYPgnEOs86IjFLm/U61I3eykILX/2yJJlELkis/8Nw865lWXVpFr
sEH+14VhsnOjfbf5dsRqd8SdmnyFjSIGYQOZAoFkLpNJEMy7PJAOAO9DPkHpFNBfJ4/spElEXIc4
tEOFD+38QQ5eIPLBrs2K//7p/xSeMRChUvHsKedh/DK937G5g5vvrusy3VQ6j4jKrxWFrjORFAB7
jBCE5Dpm0MjVvqRfb2UavRrzJstsTbxxi6WdJ1yf9eNSQxokM5l1JvC9l+rh0ZhDe3R9EhnNGWgx
GsdPAX45hfZqGN7TdgAcDLk2Fomfs8bNCq3a6EfgJNUnrHUVL8jDUDE7Xe9rtxUNZFfOIkw/PnZw
aaueuadCnrlpt3iDh311tcXytdOv2o6Hl+OfYvZVK8X8tsuTwt5Rq/mduUdOT1imPR20JDeXCPJL
QFOds28fSeCbKIYafumqQNFaf6EOE2PqOIWFtDZos3NZBogh1+0bXE/UPNyGH0/jA2d4CPO8G+zN
HoGr+R5G2Up8w4WdFIzNCLWLIytY7Zkm1wnC/4Y1ZjVjYQnc5VSCHdHlAf5l0IpjzM1x1ozbpFYh
KCMjzMe5xfx4XIdhNSeMFTk+p/38eVl/w46E8vlPgaJCUeUV71hD/I0QfMcvJT0/lP8uqyVDzDWw
l0nwfhRIJmXbOko/GBIDSSoXBzW9i1en/HZfCmXmlO59A5dmTZntyoF4Pxzeod1T4yVTTNPeLyM8
BvAwObRvWId5x7LyQ4wrXUsstK8CXUcAzdIxjth+w//Q+vyqxFP67wDfkLhL+3YanreaJKIBzXnB
HPgY9quKZIGE6YUrOBcD2T3DHNd9BHmABGJr8kUwk1lK/uArq2g9qwgTXti+Je7X0rbKWd+Fi+1V
S+jEa2yKUAkHlD52igXHmD1vLYl6wgnvXJhPmvg3AOtf3b5iT+K6yZZBMoi3xcGmVrSoX1780gfG
0ZK+bV+WKiFByEDXezehJ2Y6YjiP1+FjYxxVMwp8sKGOzFQ8A8hXUuCCTUWnaBuhZn2/5+hXgJF6
lPy5KdGP6rdNNp8W0GpstIYtCYftF/gOE2w26JAlNjJepgxpdBbsZOTrXoxvCawkosCLCwn7cZWV
kvW1o4LlxQ0s5N9CTE/eDHWVPLlKLV39mDnZ5hMuqv50PXwXB2Dbe/akPvdJ6GJs7X7dDp/332MR
4wkAH4RAkwrouBqcSqcYuC1zdDwXiKuht9vYbRW+Q7tTn/4hZ1rVU58R9Mt+nuVt4XRtUTmq1zd/
L8hsLY5CjWREZWhspPv1LdADFuJNdLICofyitLblH5ou6ADEFoq0pfIRYTleIv+q9QzaalntcjQ4
hPW/jnYmuQe+9egUqPjqphBME7+iwkr2P4boRqo5Yhr2vZwpY7eCechtOjqqvX2Fyrv4giHelTYC
FXpQw9If329KVgFqnCVpaCym79K3bXFCGM0KG/py7h830fljdmAPoxTY9JyvFzl7TFGmLF89akLQ
NtnsPS4HMuzLekBkEUjDb9XYBJ03VWaAWRvI8v0huggGy3tYZgKimZNbx8ZJpw+O7WLyg1JVcYe2
0bwqdRxOZ6RgT5HQX5HRjSpp1JnuODh1H1AwSEbjqLfFr5oerj7ad1x58dvS0LJC5GN3hPDfdm6W
zLh09w8haZnFpsvtNQEQ/p+llCBHV7nY+riQ9+bdcEVki8zZZn98buCeY5g0lEIT2DA6Hqsi+OJe
8IyIQsFpNITk4a4CWW0sv33mwJhdo116OFvicl3ssMstYgZE1/2wx+O4mZtLgLTix2ovC2Sngnte
jxPG2La4Bt/ZgW6XA60nAdWqfbedp0L5HuYPlPPifwFenQ3O5l3oPRgS5zufBXVu+9Hn9A5TfKDS
2oJolGgtM+fGqfwRHmv/Wj7802wjRb/EZve9EoS92z+ihMYUepKw5Tdz/pRkAqiOE0eCiklsrA86
epsyPBaLPA/hSIfdUdu7JXz1YrRRwJuSqbEYMq9px4BW9n4YwHUaGLGc3deUT7vdY2gJs4ckUbcb
y1DIQ0bOqIsZXe5Hm2htf1oXM60vru45/XWrf9+pVg5fieIKW/h91GKtJAYn/PkLfSRy8N6PVit3
WDPkrl8nMvmJZPxtTCkuRW1S8C1BCkMEaVlJaYSiH0Mwa/4in65XB11/Au1niFq84IQyp0FRQba8
WftLtzliRmO1Twq9iG4ZCOhAtUZeh7dCBiv49v7dy+nXkcjmMICDJnt4DRnpuRo+ixNPliISJGEV
mCB8CC80/ZMm5Fh0wCOsS+95Q6r55CZ2TK1kqFmpAHylSg3V80qnNgw8qJTASm2+Qy+6XK+xVj9M
YqD1ftEql2D8JhqTIdFyiaq3o51dLn9ijD9HIuj/ix6aXfOw7/YWdeR2orLONuSXz6LHdZMnFrNx
T96eco8v0sbdEndNm+7HUQzqjXrcmkqVcTWqWS/7kxl7zJUUUmPPlU0bqhYPSgAL53T4eyB+/ujr
qsTdZ+4dk2auxVvTO/id3iq+6pQImKkHQFI6M9vQnDDvCE8qfPnmEO1iMpgkWpoo9WscTHan6U1u
SxgoR0y4nqfp5m7TySJL0khd8LhHgn3TKvEFBlZMugAJOT3pK9yz3nQ9z9AQzg0QEk0Mkp4pZ2NU
W1/1d69IEMwqISgl2dOA25F3wN6czMamS9Rl1SkF98AQdnlgmdlcwo2hXqKKBrXD+ywuvYMDjlUW
WbS847qpet1u2fk0OVNHt3Y9/o4hG+u5oop/XZ1nG4jqtO3oJmzIB32e0YONMrf78fROW7olLqOb
vhGSgM0qeqe6ZUuOHQXnaoQeIOn8IVRFOsa1leCVspT+Er5Yf75bk8lvzTwb2nplDLeNj0EaxZ2I
6WB0g1ejeCiRXtjW025nuRlkuq2NcQ404lp5RFT936Y57WWvL4xuJDoprHdMe8RSfnOo7DXB4GX/
napbvkqXq55kZ5lT1+4Lg1HXVZ5yvhMMIIIM1ckoCE0PnU8rXW7L/jcI4EWLbQo8eXMEAKEwJhQS
QYHPms9cxr86zNho69v1n45LiPMkvGO1873iby2B/9LH8gFUblpKteLg81iZoMARGi/xp+BAJUU5
rq9JMrk6TMQh6TvhtKpc3ukBfAvKGhIJZFRBFug+CFLvop5KMJ/iyNPmC2pFkDiCWvCGaW/JL9+H
E3ZDlMW3+0sbP6mmX40wsUvUTcaAxfETu3UauU7TWXHbf09wD/MzB5WL3eubDOd+L+Qh1YqK1CVs
9XpMVqV2/9GvqUDeOjDBtYzCZc0GOV6389W3Z5IWCXF05MD2YbGLfslbeU0WL8Rd5me5OpHJp1LE
JWjw0VhVmdyefRcGhWuDlRJEfzsZ4EKLpf9dOzWaz3EvixrkvSKBINSwflC/itx0hbR1CAK21aDq
93LZ08+mrOCGftlAp7BuieocbOAhO6cBx6K0tBZi2H3NE7GddyyNKFJOt1JCDdAkNo0B5YLmdnTm
FB4ueJ2mf+4vh9GbPT30qpHkUIknz4JI55ctWNDrBCvKweOEQuDtaHJkM1pygTI9BYQ+JC1ji3n7
TYD4Ilqq+g0qBHz6Bep5LsI3Ca5mKUJJ2WpFgR0UJ+Q6NIcFGE/JZsTm8KhXZqOgk5coefs84ww+
Z0S+LfrtiVROj/yQ8gANBS9sdCAn7R9OXUMyulqzwJDNPH+NpYaNnENTzf903LdWJpS5bKlNnJWS
VheJe0U6mbiVMSKjK5OZdpA3S7OZblDOu+7JCvJif3LGFvKv9JCuxrBxdp7541p/VvECQ90aYrbB
EChUoU+HqVKMdOHn132snuWOiE307tgBMJ6ui8f/1nDpZUIF3vvhlhK6v6wM1wUusBe9qC2mKfw+
TF8iNhqbFryLrlym7oJzp7eYJfh4TZ4RfdDKRcEQxFdD5R0zFqBUkbavVGoX+Iuq7IIZVtYk+Kap
V/cRvdEdLJ66FmkrVYjezrv9OQNJwyz3dPEcKDe7CZ88HA/R+rhXtgLhwYPu+5oykyIksZeF2Y0c
cvlDHI/WovTBsnCWyBs/icJmAs8ut1rj8+koLARLlF2qe6Qk3RhJpdil+AgwPkVp9P929gZjEPVE
evUk5GOl406ZgwbYwn2521SqIGg/DkOCdi8C7wsP6zl8glrU3+SGM0DIhFCnY7b/EJcdmUh18dVI
hQHKKCFoLLMDB5gPSaidMdA10mvYtN890jhg7FOwkVFy8ayK+77yfnoMNVu0qBBmVNxoRzBTHRpz
eLKj1nsefEbW1AxlOO/zqLyeCQZhHY5bPULQvgNSe/fdax3K0SHIt4qYHL18bkm8PegcCbwgElbC
4jS36UFB+aVHJ836NQszXcCNSiAWLcgrA2Alqd7TVG4iD1R8bbr/210jDV65+7SmEVtIUFHCFCYI
T3iUIQo+RhoChJ14VmU5GldS9nhM/mY7KUalTXPHeegBa1Nu9OAm10pENK9Hc5oN8BVTZsdnA/MY
smVHEMmVrJSQqPyfEPTFGdiO/lWx3SGhNP4PJ6RRzwO8sn7/d57QSiHSqRlQ3cDMMQhxiR01uku1
S/Vmute56COoIljupC1T73qpAupARh8ZkIsxEMZlmnfJWOv+O4ePEj2iZUhorjsLWPEPqk4unIIc
woczv4lOuzicgEgkd+nQuzSD7kHQP0E5OY2SsX1lbf+xCBp3g/vhoe2ttMBLh2lur1AGDhpz9JiP
+NprXAx7y5gawz4jvbBDuEmPkZ5uo2w8jMyUySjWt/pIv0tLbeIW3uBwe4j4B8hUiZn81mDi7t96
DgboqA==
`pragma protect end_protected
