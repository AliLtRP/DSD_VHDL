// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:54 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ob1k9xHaAhiae1dNNSOSHnXKcAyHsfjTtVAU8ZQT5MJxPkllpUfymEYJW0k6mlgV
EPtDhHpWQYuoeY2oIMFmMirqpDfNb3ajpfoPb4FALyPSzXXv204pdppxCtKPLO9I
YUX+lCTwU5qNEY6Dwim7F43x9kUp1AVm5oNZ4W0gRJk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8560)
eO+tQg/HtHykaUi5B6r4KjCbeskPaM8RLdJmxtUS0Qs91lb20Q4vnLWVqrdIh1rc
WprpBzkum7bgpMKV+mrRqZwsgakqKg0ipPruFjkljBTN3uaus02OHHNuQtfOlFnQ
RAZOe6R1eOx6mT/P8AXbGcGnFb3xrxG2st1/2bz9FaF2Qtb2+GGFvF76EuA0Bjmy
3JO76mIreESbdo/UfV9H3YEeOpJiDbg3QDUf3/U95/H5UXVBvyyN/KnjBXKvL6LA
rP7+a0HkC2FcLqdWTNV4XFvh57Awee4D2UlOf22sio6soYlIWxBCMrIQnV5j6GbT
b83Qmb+E15e/w/4MU6NNvwpnNyXGsxAIrnUJIStVr6I1FY7rW6BA4IdNKjKtOHb9
SW+wMTeoSBRgAU72fOdRHFZi8PJQHDqDvt+H2F6v5sFEbuWsGAqOniU17rDe0sS4
PdtMGTbv4y1FqgcUJXQ6bc9gk6JMbR1UBapwch7Ot+nxJoVmtUCzpxnHLwCwj5nb
5j2Hq1kyaTyDTFvXFXPm87mr4dRs7qAMeyo2vitKGYow+EY7aqQSrcsKtWOLfSn+
xN/Dy1lJL7ipWwq8bWxEbITLb8ofIU2xLUREoQhhNSyJCEhLfrDnh7MHSouEBeoU
w55lEHiZW4lGX2f0lh44qzvCuAXiqf64+CMDQtANYxJABXTOcaDuiteJZHZIRuRd
9hW3RqeBwN3OhWQwTOVzr6DPojWgYHthGbubxhi+HjrQ779//+OgUwKfH3yxJy+H
3hYIFTwHhFNc4WE3vnjXiDHM483Yd9+3XVkv9H5fOF3paR8DHQL8W0x7Sh1SCC2k
xjC7lAVg03kQHlOmfvAKm5cPR9ei1Pysc4nn5/ONTC2CrNvkoRZ2XR9Q6vJtyZKr
t1+6kLuw4euBVK+5G8RT4/jxL6AhVnKHmBDAhDJNhdqP9Ox0CBRb7FQ6ISUyMlB8
xX8Ijf3Rc4+qXlVEB+m4050RSJAUtqFN/XrIEp1IhfSbc2hUW83FiTLTt1xBmLky
sp40P7kqtwMN8+X3sIXHCNi/tzAx1bNCwHuTSa+x9wh3ZCOhqISWHodsoncEEaNl
WX7AkWItjAZIzldKuafsPZFt3zWNBJyBiSBLCwzNRvVhTfiepv/EBGWhMJPVa4+J
8zchRNxULZzGxFZi5e6ljnDjs4XCfFDIoNKYendZCVFFtZ6Gkzhfn25587pvxrkd
U0Hty6cohifM0nnS9+AK+e7bnXswnO3KH43uJs6WPveNYG74QtVAzlSgiSmsmL0L
ADVFLqQ9jGEv1cG34uNaUc0NVfwNtg41f1zDh98KMSGMtZ6cTIiqp34GJGfhywcI
9dCx5U1kzUcvH7xOeU6tBZTv01TgXd5hnh8C02GQtyhJb20CrLfkG+acRYGXIGqh
0og1W9pEng+4PqUhXChvJ9N0PDSgAC5bAaiLA+hiqI5w+SgNowFSAMa2AFTS5BU9
bcVKl1v8AS5BpDdK8inevp6ipM7WVP+IxFU38+v8NUfOJM/1NUK4fcXoNbIyjlDf
EKLl3KYytCMvrwozkOq2nHCcXNn/7yJ14mdS7BEettG1BnxJ/pQzu2aZPonvw/t/
DucjE2mUtHTJOM4w02OtTpQWEyEbO2o1JCH7Ck1sNNmaYQ+Ngd82SQx321K1wL+C
sTN/NtrudM0ZgnzCpTDTW4CzVRuQp+kZxTLRNtnRm4JSaDRs9wDg7P7l/oDx1mf5
UU7gQYrOcSGBB2/UB2LtaksBsa/6tQkuySQPMi+Mj88MJQQ3cCxGcRqPE//ul2Xp
jHIYpzvfX11nLiASkXk0tor5b17DTcBLOrjmlMCxvDjyT+s+jTYGM+MXrvpX3aC1
Odhkv9ASssdEDPu/PhPjtLUhNTAOkC5dexQREl81GJO6Tr4g3V6rbduL6eKhF+QV
6L/Lh5MH0k9Er4EKlsKGa0J74NK2Z0Gq+TzKvn+d+20VdiFIQCmlnPW3fXZsUdCe
89kuBvmY1F7pzLeF4CpKjaMdEKurR7j1U90BomAKsdC735Wxp4rihgn1s8Tsk8FQ
jDEkXIyiAGfsGWj6IKevUnmndS/1FVmsoZAp38RaHP8eZ3xz78yWKM+3n7Sf/jDX
itjTA6Ym6hi7cspypMVd4qtb8lZsZOUvcZJmzCWlkw1rBcDIYvMAO0U6nzqI1Tg6
dKYErcygm81HJufLYzXNXGw8W+kqRdnAu0aMqnQ85Y+mXJoBX7vuJQqb/t5ir5LO
E4zHyL7Ye1rnxtIm74KwZtHoOcOMts5zRzx4DsdOK/rVQwjA9HOiYLzpkLt2pBeE
j27rsVO+lpPfwszonzTuBesZcTyaweHm7AWFLnHS1Enn0ZnDsJsN/QajzHi/rVlp
df09kcuzxkUYEP1hhscf8Iz/KI+ulHe5AiYFpHDq3PMiYIxt+8pTtzy8pHIo+ca4
fA6cj+Jvf/a6sStAjbilldC7HJM0hyPbWh4YdzuStkvDtWY4o5hq1jNuaGnpxwVR
Lth59QJreVfeUKqVowseD94x29Nn8d2HfX0+kZKKSKzJJHUAqjwlKcjXIjtQ3Va9
nh1o7calooggL44dROxiJ2RrnxI4PNJSNBue1fUTBO5GkhR5+41plch44ihRZbY+
+HXD4QLUG1tfJNZWpZpVKG6UpnR/PJnOK02QO/9PFDr2qY5mHPb8uCfEGzt5hSm7
2EKwaTnbEkF3s+rRPDnuEcjLQ/T5F62YsoiJquOKJlCF+IpriE8v+cQP1MkL6gqa
ZcDlZR867iGPTY2KinXKIV+g/pEyvoUWnB+zhouvzOq19rthxmNQWRCZCttjbYIa
Iyd8oHWd/1tp3wiJDv8O8El6dOeoPmy2MldRHRHbXlurscvQ8xVAOCW+g5y4QjvG
9kQOxUB5mg6zwecvAwf+J1326uARbz53yPaSr/5pl+cxDPM4lvP+8QNQK5+G89F0
4/8xf9GVadkb5ZHR/Ej/tN1TdDTiVyijF7Iay79HNnzbOVOlFtx4KMjMhpRxSL9t
a6uMjg5lrvPMVAOg+ZwzdqKJTGChbjCVfwDTBzW1UWWZ5AuDcqdAE1ZqkE5tCARR
/caFw9l5IOqUTL5RQBdtglyvxqwt0PyDfF8GgAFNVu9IqXJGpaVzKfPnrrZRY0XY
47/nUWOEl/H+ZsDEfY0R8OMy9tIa40QVgYufX9WnHKDcjcB+ffMFp1BGnZVvzbCg
8qpHRfllRiBAmdQ6ZZfA5XUyUm8Y3J37JtmElxdanEqyo6wh4+ZyHHz905OK1+ED
22MqqxBPMkDnltput0zQOgjJpFPZtrHHR9QOrrqHGcYBbLXs8kFYBCLt/8EyZKc6
2cGaloGLoiR1X+XvSbXINJTPFlCCc8XOYlzI0c2tB6abNxBv+SkXIrh03FpRMGt1
z4P4FU8EtYoUIoshpkeTRN4cNttvrgnBoqPmv3crEP7n/XHa5lnLXQyoFQK1DUQG
O0hjBiD+COtqXdFBfAtaIEBRtmdhDH5sksC1dou2SJRewgusRsB1x4vUPOLVCgXM
FPzwzmfaCO948R3dUJKj0ynGqyWfu7C5bYaW1i3LPrJxY4P0F1YFSlsES7ovzfhw
zCVWJPOTV3M/Yv0nDXYKWZsdzarK2cN3pH73un3blPqryNyy3dDfAUAp9q0IWfex
SRF5iBzWnb5Iojtpy0dH0QzlkC8uAQBuGV/soQlDPMKXO1ONnk9JWb/JlsvfiOb6
VklYylh75fwcNHPqwqEF09i50dwO11o1mxkEmtkSPBa2pNMpysv1JHPllR2g9Luo
yPhC4Tq4HTYPef1nVCMpgNmqMAj6xvKzydhcXpOqfloX1Cunze6K7aXR8aEffBUz
lKIQQybztHnv5QhWljolNeTHEgp+dpxupKVJNJfwfv43SwP34IieAYHH7YYDFB0W
79FPszBzeCUTf5MDvtip8VqhAe7OC3MeewF2n7y5EbuNDnMGt1wn4AzDwXPPXoeK
Xow0OFyh2lapuYE/BZUuw04IOwJCegjOAnQNRn13f7lcOXC6ncJxYrGNo/9xn957
1JVIK0w/++nDHW6M4zF++EtX5+WeEXYRpimg/p4NDq43tOjpUObkXh05RvugKspS
u2HrENCKut0SCzAyFSa4JnHQNn8klKAOHPPDwn20SPbx8uYeEdtH+Rpwsw2R1jRp
qIdsfuP/YfEfS5yTqrqpTqLDR3mTXyv+UkT+okJJKD5VsuoV9IMg3gUQJjUX5ySW
ECYgdEoi+hdQ2+NQe2+lrnAVYcS57HNKvRU4HoME3/HGcWSF3R7g7J6srFByAmsP
TZFcfppTV5dsUwIbm6NZRU9sCne9wzE0VRsWRgiHG65lt+8csO9TUWb64Itzj6Fu
qrzW8b+ss5eZ8pSBgF2lCBlDQUzClxuLGaBGMk3cgcIIGZ1weUIiXQOpEHK2hFAM
BngQ8dGm6859I5oDD0TBZ30cp1QyBSyqU+zjuE+XI7Xs2eDV0ZWA5thTvH5NycB9
JrsLmzCMpLck4Utc+ajghgMdCivRqgEVUeVrcKo8asUWvSI9++zIpuwdbWdt9QU6
ZKJZhzKu5wp4xmyygM3pWE24c9CUjL6pr3sQHuzJIv/4d8KVC5zbM5WFWBl47hft
TI+JLR3cp/YYYJvrEwW+kbQXHp+1kO3hNNA8bhUc9b5xuZfVKlF3FSvfE9rsPBRK
6ECNfYTA4ZaxrsYbJnjEADZ0wy/rlhgUgaCBCu4YvkpANO3hCWwEZO4VDleLl1Tq
XTHSUe/1XHN8uZr0+nuens9x0d2PGI8ZQb0EEfY35LCLbc8fhUItEULxFVOfwyAz
jdxVyz0xYltnt2XU7BmmZFGyCYG49Rbfl0ydPTEgaScT/PnD74vRuOO9EOD3UOjZ
zuJqn7kBAYzqM6LtYYIddOh8lOgLz4LXlNSaM40JZnpGdJM9tRnd4+PfrjRBSfUE
7W0ZzT7i7QEFUovNbUT8dVDKo8ynt5hGC/RM2fcvaAQ7t1xh8iIYbWJJIIdQT54A
iuVW3m8Exhbr21VEfR0wc3xA1NSH3bqOL+Io4/dXrpi45kH4F7V2DevLRcj4tcD2
8jdskVuZubfZc/6oakC5Rr+kXquRoPmYcos+lF9/mXXq1TMm1Z+ChKH6K8JEhXOy
FZq8/PY+d7nLVbwB7xsCd6EsFmwJHBaQzaC1AEbKrplOGZU/+5bElnG8Ry3GxChd
8tCqcvVpge8mgVKyuhQWHI4QYZp5j9LSC9RyckHd1hrzZ8yfoBzU1OuKAnx7irTk
f0vH7+8q5Q5gjjRccL138aXRo8t56Siopm0vWD6OzvfNUmuRJ/otMU85W4NYaHM6
eBMaORE8lEWWqrMA0GGplkdrJjgwcG0os7ULyiZGn+MrZVetrfSlF2szniFKDM1i
Pcxw5FcpXOmPg9ZyyLsJVGwQAgsfl+qm2PbO+a+0OU4SL+eOe5As3e9UNtrOU/Z3
YOwXsmtc67kvUt3w9SgIogmltQDiCNk5OdbsIhQccVGvGajC3w4xQWdejs2LEc3F
gBEfQ/5GSilsdhi+DpyMOIU3HwtAHO38pVv2GDF/7CrR/dMuOFkCtz+ilHwleJpg
zDjaSx+tg//hellLK+xXHQ23hXrrAkDumq+j5pOSB8dUFihv40lU0p5A5pXtIXUg
53p/dOcLW8WsKzEVm4JV3r/IlFyoc20gm0seTjPXwUr0iEEKDAlD+eMeaewByanX
irlZQOo5FlXHgKyFPVF3Y7FCWMctqyi/JE0v5mVEMNjsp5eNsXkrn/D1i28j/D4y
ZilO7Jgc+t1wzmAsWwX78pYbXxsaQa/zYRWrk6SroCFac0BVi4pv4oI7l/u1tF+l
j+t1YZXoWrodwkkO31ucWSeFbSBswFUkkhXxf047QUBN6ohf/drC9jIhZzRiBYmY
3GthfcbBsxMtOeRV+mMahp8mAROtzBS7NbG27LstPltng43rStFINMVtri5O/8FX
V0lximDjZ0gpKhgnZFVgXWnCT797HoABwJDTMwtD/1D9URUfRDsw9tipYU8K5AxV
nQJOjDdwHQlGY1ETH+9WhhUAzhihGyiyyvrBf89z5SOW2SzDD41RdrbtCpvpKulm
+YJHQFftnu7UZ2FUWdOZkGOs4tWBHF7jGNKrMiTNJViynAgqqAsMIuIWbqyhNXiJ
v/bYjhgvIaVFpImkahn56SkXd71HA0fTKB5zrkFnLI++pdgLTrljcl0RWVblGXOx
rssNPJHBYOW65uYB8bs+Ytfo1YQ/Ppgb1eLWqlEiPMmGOwA24csOy1OgKylBG8bf
rptyEqbAV0R9btE+2i4XT+i8WPDr3HL2pAPOA8GrJ5nlXG0NJQ92xGn28j4yenJh
LN2fGdmJCmt+aGXwq/FhRPh2He+7WxyxveYkG/jr7Cp4MS4cj73OyrYo55U8CGQo
Y1lqZY6kZBFMCjtVP5oINa5geMhN6gZYo89hCIF4Vjzcdw2L+5vnR2cU3tkOHEZu
HgkfOOR6usjKkvu8fDqq3nhph45CCyrxN7Knk3AGCFrmo9K0tZWcoEomC5MX9is5
fitglTaLVVDjN7pzyFkqsowpM+jggn5Jc1h2HBEkV4rdgyePbKM98auGY7n1MMOF
obmBulDlwq01x9Izd61O/t+q8/gk7gFrJbn0TkoqqlR0+kPnvAalARLgtocsIfu3
Fs3f68JqPU94FkAvxklnfGR2877Gc4+LIWFSy/uE/QvFKoZhg7oxVSd7e/Jo7UqY
qRSzEO8xYoN93GE011ynnk/x+MP20pj5+GoujxvBmyjcMPLWg6UYDlKeXgPQbFag
2F7UBPjQS2b4JzGWjSECRbDIHJl/s4Aov4l56XnOl3vfhDCNjHavtDxX9IguuzdX
OXipDUQdYDrzY5wnkKQOVk8nJiY5WdZq9MV90Iwr9+sZzfLi6JQnqd7B4E/K5VIs
A5copUj6BFivhyd3GniWq/lJMla144sNT/K2gc1nHlaEcW6kR2siQSC0o3++zJjc
zho4fe3kZhV5rb3tKLL0INfB4tylXz65iK5CLEJkELLSxwGf1c6CxROwoTlyUrtI
/EkweMOeefkNoiR7Sgr0LdNsLkxFs8GZg+3ir7dk17kRAJ/96kSdS+rfoG5T7Qv1
ReKaLksEuzLCGs5l9Y1b+c+2rjv8OEERt4hie1Z/0zKoSSVl4JbeEe02IISa/3tY
A+VWqWQAebYRXXB01vTcCz1YRJPGkYCQCnL9jeaZDYzwgKDNnnleBlwjRtvatQez
pSfHaTJxVsPWXqm92V0z+ByRJ3wAGV3CsTa/qK5ZVuC2zCul5qSt+E7K1PxiuYmS
ajd8efGdo1fovRwwHwg1wsDItOmnGioXhy0Tyj19A3Eh2Le7OhiPAoayJZ14EWxS
GfALCjSCQXpZNBBscWREGcDr7f1UTVXfVprei1P13UUvIG5Ftl4ZZ0hA1HZ73Y9/
WG9IgJ8CwkGZfEFxTD93/4xRm7gOYCGwplQVxpeRpS2kjRTxg/3NsgOy7iZOMK+r
I8uqZ8Nvk0m7iWjpc0Oo4wOcYHHSuOxcE9DtignwncVTuEUUQsMdoFszPSf8m81r
LUbANjzkwWHmQ2zngIsxjTI6UoX2IEAAbg9OHxBgDQIaF7BRIHD6Xta7p/+kWr9d
DL0B9UdnpD0AX2Uh5YD4f8DdwvSQjTFAVk0g59MorQOI7LkUJSwm/9Js9/nSIuj5
m1CEajz3DRgKk2X91nRU/U0/DQ3bSTp1/QNEs211laDG6CidfZ6+FqcPaFaobwEj
V/EoWDGL+AB0/K+8X57gazSPlVDi86GmPmypmpm/ewIOcWZDi20vC0JPS/l0Ozp4
RhwVj9WDBUAPwvZdjLK53s1I7QFNQfEGul3bi3Ddu4vsOi6zHCaPTC55ZqFB2zKM
vJMcg/XuA7j/0xCScT8HTj5LaZXnbTpQpoE9d9oSD9Gh1OplX70WVNzA90BUOE7s
6z5zrcBdZ7NGIckG97MeoIXsr+qhSjp9HBDzveTuFkL57oTHNvceHsmIM3znCDB6
9sIX0LOaXxEtGIwRJaomhGRuFhoCayIxhagTAZuq/98RXfcBJOnOBTFIhBAj6GZf
PrtwOgXuXESt2PIpXzqERtTwD/Q8C30/kyfQnwLcLmrPnyBkeupi71ce4sm2tH7u
wRGs32jvmJbtUV5rfRACQWuAdJ5rYxIeuh8aIA3i1ujKKVWfWu3O1DDaBMkvG9FS
l9j/hGwLBDPg56X/w9BabL3l81DA0Wi2wlutuD4pchUsXnevZu7CMoAbA9vih4B+
K48eRdjJbZgzmmP6NAqWHkQoUynOHFj8xYD3xEU5Fa1Axhf3vKJ90Jhshy4kPGGJ
rVz3+//n1exkX2E/uEapjMulZdKj5jZP0NRicg7H8p6WFwNUR8q5bsofVzJg+kDu
7dFFxvqO/hZtA0hJ8JM4NUhohaapsVhzF1uHy5zuwBPZMazMtdaSIbHDtyagJPMI
RKic+WZkU7/xL5k4DwZsE2Nta+LNSdhxVgMDNrUrFv/QE35n4zPRoUhpkwz+cIW4
y2XbVLPfR/z9yKNg/XbUp0QcwPbunpbRvqanKZaWhbOTeAUcapj+KvIJv4zzZ8mo
v0ABuEKsEySXTzm+7MdRbWkNzVUW2JcCHbX0W5ZekdH3Jg144bd1SnCiisKTFFGB
s5KZdmj9/2mrmf0ly5b/IrIXBXErAgXHEu++noBBbmoaMyrhlDX69i+hM6TAvs6/
wP2Loq244hbQMHBozlADT8L5Ld/g/C6b7wB9juwtm24xEseB9UV3cOxUUI0QFcxa
znFvvdiYLcCjs5twU3BLKkrDz7//zRKaOVBhY+ak9bChmOawkLrSM5CX6NT+zH9H
fIvta0UYuOj6OlsT0FEgiepiDdHVrhHo7JUr++38m741ZK4YLYz5t5dpFo8cEFaH
1Ds++XAKfD6KjSDzMmlgqiSC9guL0gHE0VvOS4LoL191mAf0CLCm+9SNmMtQtCLF
rfGX4z9l7sNkPb2She95kwdoT0Bt+lYxQ9ugyKCPGCoR2o4hQkcC1uD67INgiN3S
2RVaT1j4XhOue+QTDxvpAYOB8Bfnq+MNSU9rxSfMf1CkO+KB5ZLU+9khdlp82uC9
FYCP5EOn8te07Fdkdb0TPCTX5jO8SxgwsaBhl5LEy0c/jiEC4yTDGnaH7QD19S5d
lVbgzf2+GfTnJGOz88OcQbKAxusedAF4XsVCzPA3QqZB68OJaijJOz3AKU9TTZ5R
+caCFGZvP6lXrY00Ticrsmdxa+ctWL+FNBbE2/nY+jMDex3q3lPb6N/4jEn68Vu3
MPOIGFW4Dhz0FkK7u3SoqoD2BmwlKx7+ORynL9zwTlnNh6W9MjpyG3iSe51zNbIq
xPniPego04TZq3ahm9MpMawGQHlYFsMyP6+wLPS4HrG8LL7OGK7BvcymBM2ABeEW
knVLx1mBRzwI0zimN9iM0WhEZne7VjhKRw6NMg+2Pdd/UKVQsNh6fPhAV6+aK8+p
v1oo43lDVx7RLNBR8Ta+scyc/gY/zwf75pe/EvSJ3viveo8cr5R8uSx1qpTXH/Wp
+u09Gq/UHfBLqt49Z9bW2C1fR9mT6mE91itoVnnSDfmB/h1tFzWctpiW1nUP7I08
s9N2RvILGD1BlGZnOEspfNcTQqlbottGE+wzY43ya037uYQcUA9cAghzyU+ys2Pd
0VgeXzh8gcL6FaiG41tQMexOfOl2P6ccfY0qf9HC60X/2QEq6J6KEefWieqgMCYj
c4YaYc/FkIpWojR0cXX3vlpj1djAYTi2Ca8/S1QVKUWuyiM0/3MB1rXzKcS8xOBI
DsksINvFjzIGosOAgavcMcHfT/S3p7WHrNERfuLGWy0FXknAT7P3y44RHITx411G
pasMXe9ViRBLhw5wPKt16+4+gVVgNdoHocWTKtNsFvDpY609JxL8QFFzvojE6OtN
CbBTcrvbkzpEw3SFUIYii2B9lm7wBOOSYTdicuNry0UwwioLxgucL1wn/lPmhiJd
vzxUcLRIqoFf8ndU3SVtvBMzEM/7/alRUMLhNSXHnseNsa9HLiP8cI2NZEMQKCqD
r2DSyscTW+oGZ11BQoOzn+303SqjLeE42X37k5hJP/xgUH3eJBXr1TuteZ3doIpq
hQcH+YrFfrx+vm5Vo0TZeD601xzuTRXaIwbdR8hARe6IeUDb8JdWby9wLrLYYpjQ
H2CJr8lSNdkmKT86tjgjHHCCjrG56afCZ+300V/ZPpCfmTeipt/meK+O8hAqlpit
rymHiPqlBuyCBDOjHbnnyVubYb5nIguWGcqkZSdmm4jBl2569Sf+kpEiIWLmdmFy
/5+OKHFZ8L9DBqfQV8gtN5XhdpHkG0ZCdSRU2CqVjsBoACItvoyCKAbZ72lT0AdD
9odrKBCWC3SnvLES2h1KyFzt6urnJAWY7uuy9tpmcweOhG6BtASdT+oHf/r+gbLp
Ibuw5nI4yP1/hBhfKiwOgRhFPe4zIo14o/Bscp8ntkXVkECKk9cRzhWceGBmM5At
J9Ub6CQL5qG2IjyCBDHf6+ppj0lFlkExjPb8R9cTE97I5uBG7d+HSUqt5xUJ/Vs0
DAgA4nvycf//4EdjPBm7OLMA1SyVg1UXizdkelQ1nxEx3INkIWVHnd5ZbJI1H6iB
K+X7UJkbpuW5B+1hMxEYB735ZzOktE5o7XyejUEo+b04LCtqqFXTSTELjdXFjKWb
oi3M0o7xATT9c1FNqidXbJF3ZcF8EoJ8BOQ+UKz5c7QwoTS8ZBeJqXyNFS06UoON
G5/PLf6qjeDN32ZrqfPyVH2nm3LAFnFJvOJOK2VWZqNFJzH5v2m24GdQn0IYte2T
yMI1EpX2U4hLuvJaF/1mzryOGJsbaZ7dLPl4D2NR/mU+FrNJuBUWai5MkdPfFJQG
xy8CzhoEDZYR0vVZ1ReJm3UuG2+2PoNpAvWUjCyhicx7MqGrVZnzR3cNWiC4vrFV
WhrjRTPSxio9im1FzmCDYKBhB9tJUx3hBt0KjxafTpElueqgrJk9l2Zqg64Ihay+
9Deumhb1O7eyjqSvQ2lLJFxkoxUzRbmbR1379WKmgZz3uWheFi99ZL678gztbcKW
VCMaNGQPeKK25SQ9QQZBUaremarNJVJRdhNjkziaD9CRyoVcEAioXDCkAnM6LQPP
UqrKc4PSWtmetxEsbK5Kp31F90j7OlyYirVaYfOH8aKKEoU6my7ChtqcjV1uVzS/
QitT5CdQGf5KcIFJR/J9RdgP57RSXtTaONI8lcnzvDeCWOrM7UpFujVDk0bUVFQn
6OqaU8TgbLCrdX+sgGSLlfko0xLrm/IVdpCFK3u91x25owlu5+M9nazLktGfzG/M
kJB+4PkgxtFoLIpLUisYtX2RRYnlTOdnYfAvxw81me+K+rrXwdTcnsfPm2cHDZ4/
axfxeiZcwQe/H9LdZWvMDw==
`pragma protect end_protected
