// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:11 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
A8L8/YI0kTHxECnr+i1OqAGD7KxhL9ce8NwSA0YT/VS7gdLXR1K/PTRwddf/I4cR
/vSrU43DRPW3FQ+8T6PP2dqgwMvsxStHoxdHlxThU3t95qM4r0/CAnT+cJ6PlQJA
njo40dcRz1ZqY8ZPShtbD2hIB+y6Qx+WG/vWgiC06hs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10000)
Y7A5zQ9EBpW7X7jSzzEPj6RI3siN4wzLhb9jPNnc9y1ArsY7NyeWcdVJnXtpBjAY
bt1jzGUk+uuCRCwBYPS8FcIfAwQ53O0X3xWCTB5/+FQur7jb8qdeJk1VknNu9PPb
fdU9euWoooZklhITLhE3+k0+azpydAsH11eGz/aTM1G2qtRzyhKOoBgEk8d9t5xy
yMvx/gtakh5EPhfXe4oZwtl0Z7xrx0amSsLwmMBllwwzZRI2q0ZoeDO+qCSXlSV6
6o/DJi3XeudO5N35494GYa6Ib7ytrkUPBf8YafehrOyp+mN3ZbGKEgcuvQyTXwQX
vqhJkGvdN3JtRJbYt/iOM7nRzqtbUIyKDR42+QmrGoNKteY+7ds9T7lVl2DZDSUq
Nlky5j5ZlysA0R+2gExxpEIptsskdRHESRxdywuN4afaQHjV+dv5TACNlGqMgCpx
SzzwJ3orXtWwCL3UNd+VR01Uim34/0JL1VOHGolYD/SFTSZoUL8DtUdI0uUnXJ7w
C4jDsGu9ZXosfisXx3XyMemLQtMBMcwxUcPmuz8G6oLdSYh4HLfTY+b3BaBNgUNw
RJbWZ8lUJWrHG2VJYB1cWBe6ClLuKyos4NrFD9c2UqIXCwHzb/mtOzNMdD4TMbbt
m+zhfroaOzo7Qj9vJgfKtupz8K4BgkPG+jpQXwuLXg0sp4Gi+lGzA+dqyekdOnMo
qT9AUTRGhST8VgblLtFfY8zHRbRDr8Zp7B9l3ls7JwTaHOtj3ANR0ZQFOe9yQU33
Q9nDSgVlKpdzrcdac2aZSJLQdFFkeDJYfQAgkZIQmAJEXhUl9DVbKlai03k99BH5
IiqMi+hFfPOxKkfAQTi1pl/Sdk9KKjbG5QVQy/KkhtBhoVFgYy4AkyUaizsRpu7Z
6F0a6Apj0TJhJPAHjARvUEP69bG2kLHY7ZJYb2XhjDOTL29MR51e8KXi7mrwyTVp
U2PNFQlzL0g+UyNUibey8hY+CTu0JddL4I6h5coUil7IzplHHtgMJO3SJ6A2iLJT
xOBD673mmYKxr5lEDoIxLfUAsCkOeaBgf8TZ1HGHQK0cO2B60xXkdO2xE5gz9dd4
mzQAmuGgUGo18WjtRcdB7cSMKgTibvETwfhm+MOisgS5gWQOKf+7RdqMeq4Oa69e
bYN7SfTugNB1/060AYsFWzAnKmqHkXv5o++ZMml9b+nJ/oKk7TJDJZRTQsmbdIj1
SbZNIlURghkvl2iRcIK/E7WqRe1ss5Ne2lReDR1HZOmmOOoK0XuTNwTxyHDMF+EO
wTN/tKYVII1fG/ipYwejuHCi+BBYe4b3/LaRpb8KLy1Jphtlij+CGPyBJLo1MuY8
zbKgnahlTFrh+XBfei8MG1elXBEynUUdrNpKT5DFUW5V93TI8UX3LSmw8WtzDt2G
5Ws/3+3G5k/1qV3arCnUy1jy5BeYwfR56UBQeC8ktIBc19m5cTIER4jm9jTgu0zn
M86aZAKMl/Wx/lZ2yBVY42CCyl0XO3L4CBEQCs1iZTYMN9uIuy4PW4Yzu0yBTjvS
l4U/HQMCnRc1v6+JykS69mokQFbFr77OxtQMd5Hzh7KILDB/nZfjOH/gfA7nKrcC
f8E+U7hPPh2uDxo/U+i12P+CXFRetGmDpJaCSvunctBIHwXtIf7Es0HkEBkuwK6M
uj5lp56NeldWbzI7Ar1uNiloD8tVHX4K7XnDI1W+brpVqv89locxBAhxBRJCWV5d
EgI+4f7YLg9kobJjRCe7S/4SskL4shtmZf2QZ38FUaY+FMhZP2sWjaZC1ua3Jt1y
VSWLmuS5D/LlM8ojwS+/0+riva/VjbBjOu322NpHBzqVTX2MJy8MxmuOmc427zaD
loCCCPOZlaO/SH0rQ8W2o5kE8rs2zFkZu00vpu+nDDROlDjaRKy/ZHmvXfeMQQhn
2BXYwUnNJSpjfdW+1NaxzQSVQpmIyNp2RLDeiVeZz+SL4Dgtq/BmWH4EjZ7DRv2P
AeHaIVmb4pOtejaPMlH5vwTw45+9iJ/WRVfxfh6emQZ52DTRc86nYgaaqt/Tig3/
9ycJVPooSfhlFMFhn9EsWVPbgEBZNomVKPzTztjdiwPNYVFuxMyDzQFUmzliIsdt
CK13samI7OA0f2TR47XQkUcsxGEhDGyUGkrO3s34xq1xoYDCqvxDvod6gNEJ01ps
n7qVxgSVYMeDITsyys29cEHSCW1blXlvz4//Nt9ZVEAnZ3+4XtTdkIO0Nf0sI/yk
nVQRZvfDPbJogCAvOr+mUR7HvoXScKI9D33jW98AImUtuK1PN8y1bW8+xCIY4tMU
GLAYHckqzL/U2TvnUpmsPvyAsqLvodjN597VHXgEw3IZmbqi+0vUZLPRDUlobxMC
82hbIAdA7ffenV5ZK7dQQx/TBbiY+LmLF09kOAqaMVt/SDi0iaOO/InOW0bQcMwD
OgB5kAoquCyCV0qnia+GPogHzQVe+eAs1iJ41Hrk6BPZNz9kY+2UfxAbe/Nt3tHY
KDUcKCiNnsPpyf2CyYVr4hB+YwbjIA5gxz4cLdKR2u6kO7q3gm+7TXfGQAlUFHx6
/rYSrrJ1uBYQmmoOtAThTdWo1u14KKfVVrPGgQ5YDhYmjrer0spfTkbgsHrWc/uW
YEPB6U5axAiTJcPM4MPfMlvXFriOANzOHAaOvQEkWhXqYsQQRqhd+aJipcHG6g9U
3TyC2MEwABWiAo9uubU7GzO3XvcNq9XSdqtCJUCLvzgey4nzC+Mbn4tz9wDpJ6fi
tCG4cbF+q6DJBjef2FvVbXepkitgnBzZTSTw4XXI2RQl1PGPU+euOaIwZXpdAYNT
wzVAx8QStZhtqJvZnO/iM1EZn/ZH/hiX3X2SKWHKnU+ttC0H6zZMkxR2+UsV7vjG
HnrHm08BLKSw9g43q0gG9pHrEj8HFopU6ryUYe6yAsXupINt2Qq4kKKo+wBwKp0h
pJJNlLm8bQl5blmNPFfjS66Msd0Yzk4uR07huUiUidO1YkF6yycpmcFEyH33+kJG
YpL/EBJsg/1jRwXqZNKhdIJVmadw0f0Ecl14tbLHzOiuvmMjYRBqaZRw59COGOp7
hPlbMC/goa1K+eqYQBVG4Tt5aTJzt0xz7zD73BxKZ7rl0jiGxo71AK2zobuVEFZL
WzfMqw3VpjGxfF2OPSnWTRdKH/l8jC+HK0R1dYPH/HaBn7DOUfdmvtbBtjXMjZ4E
noEUadZUAlOuH1dyqxRoeWFrjdhmRgK0GK7lvfr7eVyOP3cOx0wpVlfir/BJrGMt
lq67hr1/YU1lrYvwO615azbXyg+TM8R6Fyhqtr/T02j5JuNDB9JFE3VdYL+ygbN+
4Di7YqEikzB6BA3fj7bvlzqN+TOnDwmWt39Je9UDO9NP+1vTBaYcXiqt+g8bjfMj
QY/wiMajLt++xWgv/yNvukRjMYsIoCi+ZZ/Ln6kIIzzjHI5mUZT5/7MIfpY45Yk9
uxm/iqbSNj+9OUg5NdfLQphq7Iu6JGF1RMWhBkW3X4cLt+9Jr2QeohG/j9NpWBgI
73DpodKZWMyDbMc8shG3F1l1b7fJTDqMrIloGuHW4gD8wkECf5lH02S1LMteU234
pWlL8O8FFe3gC8TrDthSyRHO01gtWj72ScqNzr8HJE5SbBbcp7xaW+AW+JG3ddQC
DmUIJ7WQ8VY0qym8Cj6ORkNjwTA5bfRMfatcqHnpmbMZIM+ikvqkVBL81O80LHfm
7ZHvRBOX1SV/hCWA1Tl+NFAou7Eey6UFppD0y05OilSvfiWLRaRGmyCNnpJeQyrG
TUq0KSZILEEWemfrO8DWwF6pHkMO3ohgkHog9eN/DEBZZPmxtsTqj6n3UH7JMB8A
wZ5IbVuLbzDyv+oyZOl1U1E96H/ljb7TW4oNqw2mX6pWh7480EVG0Io9To/7Z3cy
Q81JRtyyEa0lfyar4i0yjh+jZXlWrn91fAAaS2C3Hhc35XA35dBry3qM2Oq757BB
NYG9FkbrbYyirqCiZO+m9W2fADHCYjwMtpYNFu9V/8ADcysW8YSP2mwNrXBN4WiE
XxQeaqnNYC98zpyZ37VLc+XJDaZBRfE/q+bwke5yhkYHNCfe0sZhQbjNU3i4nUTb
iVqXvvcon6M5yBeqIQOLyPyMTS5b4XfMoqXE7urDWZJOhjXjorIxrt/Ll8Stfijx
KZhBqmu6pwL4F30Lq5KQA8/yEj0cZS8OWDGtSJkBHON2cJM5zgZtB7gam2rO0GzX
EsxQqUS++lMbNTDvMnDwC8pkq1Jm4SFNGU7afSiA27o1FmJ9mQRmsgKNXMzi2MgR
KVqsN5UxIzC+jZfVopSOG561ZddrJHI7ZCq9YDHCB6fb4ibgd36qs1NbvHFDeqgy
LJ6PTtJM26R2wyPikGttr7gkfg/nTWqXt/+zeM3zzGEXhT4s8btur1/aaK1yAytk
ShdA3VXiiY3FmTAO/6Zn7eZa3LEQ1RAyvydtiEuTXQD7awyZsM+0sY+YQrf6bDIc
LZw/PLi3nRBPCfJSWX5cFdjg5JBiF9BvbtlLMq7niBbIf18NPVU4fNKCoAwgqxQe
VlfZeP8hedkAV7tI0Hl307lH++9E3RfjDsaYsGAGwAUw+ChkFAJGg7pLa0cHu/4E
1TbolqDToPykTwzecRtwFu6dcpwU2xyPLMGaT7SlTvOztBhcayewxLxh1W7XVqPh
vntsG8FZCfa7xsGVahcqTL7piFBYsRBSnoGM43IQ1KFirZUXmKKb2JG3WnehKFVz
pBToqobgQI7RqEuMMOxR6GCE2QfQcBBsR+U4u/MJZdMKzZXPV1TjqOReDe1LEvmC
Hx95IPbgyne3Z8aUzJ4JDFingwZkoQNz/NElZiPXWgbNKIXu5iWs1GOaJY4tZpmt
CU72BSghqfFNlh6m21GFs9hXSqZr4fATCmKodTeBHWalXFmK3iAIe2liGXIEfPbH
w67mV9jwDx5+lJa0Q2L+xUU/Etot5ppEghQviOD/Gn1JOwq2wM/YfpIxXjHEaqmx
ThBkg+85dD2m7PeOae9neJ4R/QscCiBSzPzjhShl7j55wPyxC+1kC7l91Lg6BvuN
m53t3sDWfizdK09/pWVbPAdeixAIMU4tyXnBAnDESI8fFflGw17FC53Pm9EB9bDw
sQanW8zBm9mjc9uX5NP5FiS8teW0Se/WMn71KfVIj29jnVjLmd/cLHVvCWMUa55N
lwUGuU+Kd2DtP/sRUw8lRyOA1ElnejYonW3qLLkS7yK1zFgIb0YJOPOymShMo50+
Kt90VF7M501kafLLOEEN4AYSAvit8DeC8hVbilgSV+AcFY0sYlOMsclTh4zFrLvC
cVU+B2gU9MR1osZjJfrFWbE5fYtDgc2fHYut/EbDxxQwYdVA3QIBac2Yhj1nzX8R
Wis0wykLgPEKFOFqmcrJU7IfjmE93DFPfHVj2JXEO1xCAMmU3gRfTydsjFmjUL6B
gyBUSWkf3xmziqWwXd/p/eKdDJDwywBgN3Lb71nvSn45B6W49wmyET9q8DN9euIl
/Jk53PknXrBL0MiCEHcWEk2v0IX/OWlv+6hq+27Geb9ALoSH2yAYDwDnKSbqPggQ
+3hauUJ7FBvETNBpAfQYIL4DYnzEYvp7Ya3TFAqs2O6THVB9Ov80ySU/QrEeeXvm
doioWV01JX6AbL86WVWaThhDIi3mDKALR+ISckzAzPmbV3pLCeHKDVLf9R8MIaFu
OxgChDXJbYsqD3AUtMugDn2a8od/DKdjakav+TYN5T6qzJburrJyDtCuo48o7j71
T3XW4nCvT1YFSF0czwOgBua2dKhAnFwADsrB/PIQ9NcBQs6aRxczrEK3D9yGpD3l
/XyoviC5n8ntBdr4Z5eKGTq7PkDoEl6bPD7NsSoBgMIjKdebf4oTG/J2YA49Cezu
PuF0zXYHNjPuWo09KCHA7oTYaHnwiZJtOLTQoa0Pe7O8DcX1RUKVS1cslRDYeb/p
Odmi0/2jOaS0nq6+o6hKazFzj/KYZQRZhxm1jrUv9CDtpscnOhxgwQRMSxWsm4nQ
JpVpTnwtrdpt7AtwtZ2/hiwZjsVBkZmuxZ6dRWWH0Thbrg9lgodqoXRQinij4lk0
fB1wIXRcXIHZVKyrtjWOqtzpMv+wyAROuxtSe7BM5wp2Z85oZJHZ7tNJViFPgp+9
26ng24flYNEpVdH+bubGyq/VrrTEbLwi6+zxbyRlPD1sqdjVbJFy9e2wzKQvx+bz
gU3xYH8snId0MiSTmwCKq1xoqYbLeQgkhZ+5Y4loltZXTrXodMOBCxSLW2yJ8XlA
DnimplNH2eMVBPdoDDMw3XWCdM73g60JfCAKh7JBj4dqXkNsIjuHfRWxLYHZBke3
CM19yXXUR9P1bTy6lAc02gYemHtlodIeX40G2LbqXq3YRSMgA7Nsd06fQljfHH8V
bGKoirUZg1ih8050OJi6g6p5vyKcdpkdwzMV7Yph+VqJwJnI6lSHR+dL7E8a4iqm
FBk6WmSBAwaHarnS10eoMa5o3lmvNzG/RmWU9knKPFHJOiUiwurCeH2JIvJaof86
S6iRng/+/LwVYmY2gxp1rYn1EFme0pgIgrv3E3r2nTdD02newwd5OvsRimNGGb+E
jJJ393bA+sXfzlt9mLTd5VSfugz+LfEaHCVkWR8M9w/CYr/FN4CIac1AOtZiw7iA
UnrQ5Ftp2gjXuxTJJ2qw4YVFKQQTTeLCz3/XY35Vi+2efXBmDcMm2W1V1izHVEjZ
p2WRvrpT76fj0eRdcocR1ua1seUj+C4VmVVyBOBpiyKyWvGO32F762z5LnpMYD7A
xbEpaJ+7RRyjJ69/LHdGXZmDrm8Shy7OP+av0FGYMhYwNIlQ/q5fjcSRSi3r+i1S
bNV11uhw+zThPc7WU3jRw8sIcbWzBIQtubqpbWbYX/zcHvd5Jn94J+b3CG8lWLlx
SOEGCA1YesvRih1oOdMuS5loOWI4qO0ZbN7y663HVv9lXuc8eVW+Kb4gJx8mP7Pu
93jEbQivU1L1GuKqQM68sppi4gJWyp3i3AhE/HEPYCBq/wgQtNmZ/KDV/FsbZmQv
wSTH8Cm4S3z9FzybDSYEUYOaA32BY9iFJXXY8qnFIwHxn8Ajw5+GuqmRT1GCJPwm
ePv4ivHILjPjxG3+NHSbKVVC27miNjxgerotIHBBCekFs13IQznEiAAg9vyiB5tA
P/Lz7g9GKLTLrkpa13LqHD/NP8yypniYOv1eb39MW2yPh9LSx5hhAQRMUDsxg6ow
z6OmFEkQg1DjLIRySF740wQ+TBKAr0U/WGBjw/JSVwoXwXBrBG4H0aglfb1dm0Y4
vFhKlMX8EQfQzjs+QIpwKzCOAP/SJnaZqhalJuJDQzLca3kCqyojS7egyM/p4zX2
FZc1coziG4N6f5xdQJpVCkNCTwLLAloZRvt7s53Mn4u0/6GAMMrvcsZYLmZ4Sv2W
uwnyp4qLfzBKJ2yVh79rspSy6ha4w4W8O2VYjpsKYwSyZzPoXnZFjpDtVz0E9L+E
ku6JFM1lLO8t26polqXN3+Zh1bi5zNkyT9uXnbhWosJN9fuigCGV+arsm63yt+4+
2Fwl4Np/rb1QerS+pfdhQkhmN4zHAP1ylHv2kVuTpp/AM13luRBm2xCMoxrVSDIy
UZUw3V+81x9W/oG5KhYTHuXpDGI52Ir2A0ws3lT7Um+MU8yWGhPXvjtyQbCfvZZF
VMHE2bYKQvxUB/c1WIkGE8Z0X/0CrZNjS/9aA3v9JxojQ7jWGq1A50yFEBWwI7XT
RNTGbtIIriGAjXglKFJuLZRqOlTW3cmto2Uixv0h/vN0T/SHeMYEubrvSioGxIaU
YnQREq0uKLuFQ4C62WP2FrKt4UkjEajib1L32LhfRWVV5SNvaNl3/EKvmR6IiS/u
qNIS2xupBKrvG3xxaEXururN/vGdkjfxAiwDICbr0TDfSGzKRmVjFb1tBRcoNtAv
WzLubSQlLG8UUJ8aqcvJqbVLN0JRQkZT0hrdcpBitWYBd2NgG5+f6Vxrdlil9DIA
7z0UoonOeBbBB5qf0BI2qo8lyWh7751lbpb8sRgBnUtotiiGcIY6mWZEGFdgFl1e
yHkHNJh8T44sXl62+lOaogauI9RajkEVJLAz5EirKgbxlAAk0lXcUMSV+ngToOEH
zqqEfCh3B2uaqGH5fvg3t4UlcCM1JC7IEOLvVv++ta4kabIw4cV8Y6Gy18Y/cLEY
3ZNxwrZZg3zDjnaCTYgK3B3vt3WK6+ba0kHjLMGv73qe0PpFdTv2iM5R4XXWh5yx
AHDg0LnKz5ylsieSSQLJkPet/Ej8tWpS07sYhjflPYsWvmhBIUZa9VDFStX6et1N
dj9GOizs7RU+JG1+tBOLTg4SdDG82HV2jomZ5GFXmQk6q121SMpkfF7ptWuE38hV
cJCN6GWVN93RwZQtDQ03DK5D2PsV0Di1fGyHMff7rzPMoJDwblewgugnpSgbpf0I
fgUwfeFfCM2MdXzP6CCKFXtdFWrGatBx7K04D0pGnu145PJjX7ljs9Vg8hHSD+i+
qNnUJdKrtQh6B520g/Yb4q4QnE0KD/lJQBZmF/CCR6bbqmg0pAJFbScw6W2sSNwK
4rSL6CU1cZrfH9WxXBAo6YtKzSB/46PTMUJT3WDAqYmCbRJJtTccwczIDU7wfrC6
N4wc0F+tYAaAnb0u4+mNgxMcvFnY0+Z+YE6sWELBDzV70niR4/AflahKAJGqXtM2
KCxvXd+uBVrCGJm2OULrpHSMMedP05NxxpnmX20tH+yxD2mF/435ZzyE0xEljxYK
COGeaotwyO+dKGlGd9h9/GdpRkyklGcfODySLmgqElpyCS3fIs0laKwC9sChJf3H
MsinJmCuHNOocwOdFCDYzZ8lWC0hBzLh4phvvvI8eIGlvFmKsWnzepGd7W9GLic/
ikKrKu+v5JwuaXjfS1idM5c0rK9occt50l8eMACbCFiYdF4s84X+XEa4D+cVs5DB
Z4/mS2qKQXtvWuzOQRNoZToyY+Sxa10S3A8MK6HGD2Vw+Ohi9Eb9QAM1tXlol9Jg
yWD/mB1wb7rSB0s6lXYDyGXRrSYya0wNj2KbPGJn+VIh4FrdZcPsUDh2O5SptosL
jDHTjB46gfPlSPnYvF+pXb5+F8W5V5cY/G0ZYuX9KDt58R0z2DX+1uQShsR9/Ni8
mxx2L6CixdldjCJmzmTOIPfL2y/VIlXwnuOcKvuuLNtm+CH31CSFvQSZ3VhrWLim
yOR6MvgPfg5H80bwygarmgXFzfSUueaYi8fNIlYEZruWyNhWP3GIpz5g9iqJV7R6
XjPXPrQcw/xMK+SNIkEMZO8OhbAhINzaMAMNVyJ3hbDlWV8grh8aprSl9+jmYHOD
Aw1BfkQB6r5r2h77pyPEAmhuTpHlkM2Lk5kEWJxZTgKGYm14x7Zm8iiUSn7bqhPn
7izOZX39l/61oGvFZRQRnGZSSGp+zIQd+GUuVeLol/Qch3T54ISbwaeybki1UqRz
8wYxxaZMk1l8iml1Pcr8cJdNdpg52oKHOxw94keTpZovVK9+t7RFZlq97J2pITvd
Jt0Ufv8iFhUZBkNBEeXlbxhCrUshAho47eC1BViavSA1Ljurm8/mSJSBfxJ3ETQQ
GJl0hkFoQ7/pxCBUxXTFSoNo7ywD95EgMNgHD/fU6uSfNYY6X3qB3SXneqWiWcRz
patLIXgAUgZ7+xJIK0RSqxRAVcm8PEEfzvRlhx2l0y14CeBmX7gR5K6ptMPguzV3
A1+C5Q96yXGSwIHVDsxt7285VuTySU5mJdZtk9IUyRLurQUOBAYwFY/a/v7ydzvU
I3mvMWIEwqZ7zwZtsHmYy1FRDk5rtVl3yy5eZdM0Uwpqvcpm2Y/prSna+vSIkHGA
DyqPMjNIbX9NvQ66BFOBDF/QyeT6o8AOuYLzb1O5lHKDqQ/16FxkMM9Ut2qd0dRZ
gzPbwdxY23P+XBLSDZFIkDGk1scgEMffoaYo0YnGv3AksYFD1E0FkJiVRQuZKaWA
+YfBvM+ETikDBL34ZmUQCWp0rwmQvpmiu3OaGNEQYnyCLBKjR6ycSLwK+GPh+OkA
0HFwK2zPUH0DyO61JtgRTqurd7k3zcxkBBg0eKspoE5FE+T3UX/sMFj9Fy115cb3
bxJOVBOUq25gkrXisYTprbGBm43nQ5kVHJ/7wtWtofAhyJp4wmli6J4DNm15rqM3
6YdH8LcgzOSDUDS6ZYEY8YHb01wVyLb6KNh5MoLh2Lulz0q0yyzYqZDn1rcE3g8q
2kbMTt6rIMVlYKo27pzbA2Rkw2mmXpvL+Q/x3+jfphXcw4SdAB0TSeq6S08lLcD9
55OzHfPx/EeHSVZu7tCKrTfNlkDmLvnk1+H+vli8pkIeo5hR1JCLn5xL+LHdzvnS
bWm0zWv6/Vm9cNWwhCwSX9879SXsHa1a4lZGmFSlE/q9Z0GiEWR4t0+b42PKkPqm
YX6kpNNnOXHNN8uEz3crgy3aALty9GyP3eBKq4WS6n4+OK+k2ZHUhH+b381X3I8Z
39b8FsvEVKwhBjrw6d/LVpxwWGglfbaKEMLJTU7QX6cnj3c+I0K65muEau5FRS/w
sfoCWvWbkqVdDVJ3UCWKjLjW5hpPdgsJ9b51Zea6KTbZ59tZOR/7yME4r8sy5lIj
uwMxECpM4zUr+5NyftdutV8wmWdM0RgOO97nft8yCHX1/IcqAHBxDgXPETIklZ34
kEBEnnWlTGtYqg8+LG9osiI1A6M/nv952WwxsBuCWToaihfZFCgDDuYkUnCfQ9rc
UpWnBH51mlyhjpR9pAzY2RWetu5Ra5xY+OS6bL/O1gmknGkpJy5ahRMDE4E3+1n1
iUFdetQb92HuOQF9xVK0gqCoGStdzxJv+RCbJixNWDa7cKhohTAygm+YCxU1gFBS
ugS8xhkjiKNI0VK4cCF+htbdTqtJSN8zb9aXKqyc2Y6EVEKQhgvekuxhjAiq1PWD
02kj3kMU0lA4v0MROijUnDlIYsh3XsxrCkig1j7LiwzkVhlyYLvcDrA9+3eH2hK3
GpHvMj0uQh1heb99aitIxsOJepMFc5YdkQEqBalJTvoAMZkAMK4J66yF3t8D3yz4
lcXOAj8riIYTClz8BDc+njsE8s+HfdPA/vF3P7X4jjGHgt/f5dg0NPIfO3Y6NifT
OTy8NYUpecAkLoSEld1cSc2oUGJax8JwXcRUorSO2h0StVedpMdgBDhThtzFDzMZ
V7vyzSB2S5LdI24spwmzlSuGYTmXl/i8L5PHZZpe1IYyQgTaxYxsEyL8cERUWuzh
J2HZfQNCCVhNkXDzVVvwb0GdDyU2i1a1JqcECqnoio/3ZYkgzdzH1+jHOeUIBPy8
FfO2wz84frGbe5o6D+iq+mvBxOZvqw1NRbGojEXGSVqeV7EzoGUhaSDRihQRsM5J
Z+W8jGMpZhILdjZdm6c5bT889mXRGEGPrUe8rQoxpMEltWZxbO68LRs+MmzLkY3s
NulEJY7zuxECSGIHo+DqcBhPcRprAdaszH3/+nkkzYzVSEBGS36qREg2Ufni2Uha
w/dejxO9LnTdrKp0RNMDipWWx6Cr816AramS+LKiXvW0vofu/clcSib4O+V0Zh8n
TxIeMY71rZobUXtqLbP/GhF0wWxtIb3GaHmn9JjvERsklnOrVXnVPtUzflryfM6w
jdzKbPd8zEbc+4/iVhs/SEmnI1zW9psrDeLD2BQGJCpBZcojJCCnY7Byj5pySQVl
AoFMaXkWMMdQewWbJ0fVeLI7lDtz/uTzoSvWfrft233tC9FxRwa54pQpnq7DtCqI
yiGdKqOETC+SvQTvIIHOk4fwkvE3+TzyuVhDeGtoyoLIUMDUeP4yuflOyYxSjFlO
6rqfSjGYlqwqnbzNXba8UKspT9J4KXHRVyxdcrATwxT+V2Qj/AoIMUTHf+xxatat
Tfmex/BcesCM2HP8YI5u3F/3Y99h8cM3acRyXwruveiXMTuh8Di89RdEhb23ukT3
6EiDsbvLoBwIjxr60xsRsxxzq7D7ju2up0hRJtqVwQtVSLJmgaBilm4tIejwSskm
W6Pg6rG3LXXdIumKyckQZD/Fh/8THwICISW/NnJq8+2t418rUEhIH7JKeG/a2IuC
tVO4o8om6sBqVXlMSC/qsYYbwMBjEjEa4ccx0A//NKUZhI3b0RXlChE1qDqLIEfs
+j5NZKRmdwDRKzzTSqkO2E2unuOndrjtCLJCdJ4P6+4B7terVN9BN4kax/xk5zwD
iTJxpbADaPcvmL8ImleA2fKGnFJdW0mTsAPM2bnEkZ2Ji9fPP8IPsWGW1B5fQ+ui
0efop4MdiCj1nWVuesjeqa7MqaqQPo6iLty7GZOyK5bhGEpUIGeXGVl1SdmmJQUz
b1bo24MJ6jsESwIGOsyWaXFl4D392eVFSBuAMP8oPnnTEVgIp6ilTAG2sO31LcGP
mftqzuVl5bNtUcl+DPbTfADDMPLm9fNMy/DNVIE/qdhIG8oGkonZJIcsaaw7pnva
DGaVLE4PPDoElWTSibnaRT1r3mKYkO3kPofGsyVK37ZbdX69p+ftYT+QI+6B0Xhz
apYdsTYIN9Mz7FAsQbyadmctbdIWps8zX5imilZLk0V7pzcWqHilw9Fh4IFF+mB+
PTx0rgvTO6gK9E3bhtY5KwRgnoz6ER+/Nqa66VLJ0SvMXXz+Lb8KFi+Fy1s+KHzM
+QfG0GOdoHcl182tMpCzFYm1mAzKQJgYKYiDP7R54K6LAe/Hy2jsHLOR6jLoCMeu
xBBCrP2I8/KbHrzA6zviUkLcpavY5HDOmogQhlBQQpyLokbJZVWZXtp6LJSwgA5D
SFX+tvHKkal2vgmyYxUHnPZmy5A4afRjBakK2lQLMhwnk7Nuqz2NTvLdX8Vn3J4f
YcbvXvoZIw8/zm1fHorT4K/gd5fWouC53N+tctxPBtk2z+OKkXcyemcsdNVZeYyH
1rfzCjOwE9z9rEfVvRBmBt+ZGgTQcmx8hpNX5PJvf8w71k9qpSPSVBuzwhCccWNf
S1oub8CYF4Qm1d2s3SnvRISs5t2BxmmGFk/q4m5Xz5d6V3WMhFwGZrqoGvQr0CRC
rg9fVdmtQRvX8pKx41R1WL4lK6g+K11ks5noxE09+tJYtur6TKPGfCBKIIzxNz/O
u1F8XSt1t1ijrlBOIRXevFglAo8+YMI9bhAXHLlg2JV1AkyxJzMROsxSBeZ3+Dbz
OQa3TlGSAMShq9tc/atk9E1Ohvs5g67fRI5/P6CE3+T6LMdSS/HMxsxG8N4b7PVV
CrGg36L0F5FDDGnA7sDklfnnNHLgrH0mJZ6qmvE4PkCF6wilkdSJ+8x/UeSzcsC1
IOJlGw9+TxNRqPnGZqKVaw==
`pragma protect end_protected
