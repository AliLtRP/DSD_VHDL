// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kRyhd37LJ/o5HJN9ouJSFvyb++Bhxd7RFwbP2ARUfE0ooxfHNoGB84NwCa1pBY+g
g3LaRKTPyYKKuP9DhqphPrLZk5VEHY9XDeaO+e40NmX4IJMBPlEh8MyF3SxYIw13
fW6JT1Lmlt9YAYG3bOtX+hy2ttLstDSQxismahMb/z0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8464)
INJxPItnlkO3Fwg9yopPpNAQZn7aow3bq52EAfpHEA8IyOQzLloKXrHySGm8Uv2K
Nc6+ijguJMLQO+oy8Iwi526tEB5piUHqs7alotH4Jd5+6cD1Eqtgv2FSqn+FFkzx
dHPXLzfsZ5aGgJsMtE5OetjJb7IW/kKDjQvMxf1DJJkyZ/HmoioicbzNBPYDAxJB
yu8Vm+oU1mopQgwoYjlaaTKI/2pQbBX+ddV752TqoFc0+fpvpZWj8Q/0u4cj6jMe
UPrld5vNeadp6ORYZNhRnianqSPIcLZXq2bH8hOXfkCZeBe0S9cz6EArNX+DEGQv
Fwb/52N7JiqtEEzJiC74NLfuGMdWbOk6a8oV7FyDrtICopuD9PU3GJtVW1PrWOX5
/68WSUiHSLMmsjEzMVp75lzjuTbWN1Z8zuIHDSLCL4YDHNaMiKdt9mjQj2FrwUYt
si1TqFuqX4IG0gI9gF0Jr/VS9i4tPiSDOvnUphFf8fwXvmxZ9t7X9QOMRRlrP3WL
Z5xVehlwlp36sLLlntCUP4pOppSJXcYQzB9nzf8L7lZT6rfftccuZZni7jgKVnBa
nXAakLP/rsV3srycMM4UY5efCoCv8f4Q7Sauasw4sKla8v/BNVUcLP47+kgaS12j
sgj6RAHdeBscJWE1k7zIZ7JFMDBDKX3BfrJRDKjV1susAZjTrJcyosWmw5LFOn71
LAle+o8+DZFFLmRqL1cvutYGuFIw74hUYEeR0Gb/KORVQ3LOExR/BHGCJBClk0YD
nqUUqz0NVrDe3F8GmmVOr4hEIclfqCv6ot1a23umHPBO0YTeQl0U1N9LgcOVwx1u
SD+wtl7bNJQwGhQoo+bs/ybRg2crYYww0Nc7BWh+xgXn3v0bM/zik9jQmaljRmQL
ZcXbf9e2l/5byTS4wSTyHNJubJHt6748MXpb6rAAspp7WVp8NA541MkVmzgD7HZD
wcWkg8/CTFvhM6BI6FcC+NuBtGhLs45E5Ix7GYCymAZAwXdDknwqYKpw0x+KjZ01
+cnr/3Rkh4sLctF078OuWO/URMPQdP46VOW4mmj9MC0/ie5DG16Y1pUAW+AdCxB8
Qr5zivQk4c8ivtftN4yCNCfVmm2FewpXGR7jPjMGplCI0icd9uIXZQr5eYYqpNiL
pkWEamD9Fo+GFihK3SVPhoe3vmgj0KxZiWRAObnzBYrJCMULsIpk7evc5PJCBzB4
xOnyUIsbzxGXdCsTD/jW5Z1NIspM+3ZqSm1GIW2Ct+gtMQKn0tWnJ1by6h+iFzbL
LViqHFSoxqJsHwj4RRXgsTohzxyYQ61h6SAxLk5cjFrhpedWbbcWqh+zes2AF9Km
AJRoIzUOds+5vNWOaHb9yndrVhM+QhGdOeVR2tV4PoB5nVwkpm46adiSa/NUQiCu
NkxBFALtMpOFpa+Wwr6kF+L6ioEFJoVXpIYIeMAKlqqJP8tvui/2BZNFGp8aF0M0
XmTc/gIml7YWvI2I79rFQ/2j4U/AQTn/j21JGE2U4AODfa7050As7hymcXSl1fh9
4GgEa9EBsfa4H0hG3X/vwSTmHX6ZXVBNBIn9NLud9s1la+Mcvn7G+Ufg8OrkHmLR
3lOIqW4swq0p8FPk9qGohF77Ey/pMHqbYlIvtf+ZBM5rEucxFf4ACWq2XN2ZHUUr
idmUKY8Ht+3o93odKRlI3rD8BwLWmlFnG4yw3rq7RK9iBfnaMT9G8q/NnXk/17RS
lS+flGLmx85BlSw4By3Sm8LFdQbPZximZIp/HADmFiYY1qek8gCSwOmOw96VRTIh
7q6NgVdoSa00eEvXN1qH8Fy7XrkXTIBDSZxl4QYGYmgn0P2Pvv//K+3zvM8kIGaV
U19nAehUM/xzgBWiNyq3gIjWsxqqmKswbTO7bbNODi0FenlQGIXf3EuLAL+lsTtX
wjxTlZ2tJClZLIYmG6zHXKXTOgPIg4Q5WGVMOYRR4+y7F+7dW/AqgbWgMTAc+bYf
L98lLJXkyTMeH6/hhC9T0OtINNOMX258+qeSAjLir+gKtrrXZPiTD6O5RcTxqoq/
CnCMbOod5BWLKwADHe0z6OYSiq/HsmmqsBqGj/ckD+O5c7Z92FVO3G3Z4OR6Yn3j
nndU63gSIRFemqiVTdRsuX0m+KT59M0lO5kFa7q4zpBbOO7tt/GkmJhCvrak0EDJ
8gMjgzKIwLkvZf9Xe4mVvdEBORq16E5LPpX4tfM0yypJykhPqtAUproqScwVzOZV
1XAxVgCXl4hXb64O9zMFNXXVeg+oK5v35KviCikCv9c290IOFlJ9BOZOOdJJYAlZ
95hfHeib180gDELul02Mtda5F81CDq3z8RELH04umOusI6gr7BlWqOnRauadsxG8
miLbPx7wMG2IZ+CbK8PjF0JGIrvZqfyKTbeXDbqNb6EP4bCYcuM2k7Rq0l7E6Osw
aAoy1dT9By2kFhKH/K2mNSsG9T0i7pUAAMzUhMl+ldMQ3/gZEIVD2YKB3WwVvHuC
ZqLQbkFW/kuu6Df/j0lFnYzYo6tvCicpSF1OiZE1VOylwc8qtJ1PG7r/aD3gmVB9
Wb+wRmDQ4J+BSEArlxDIEvhDXEY8SPZdywLvS8+oN4xSH4CEyKAetYWVC4caEZNA
zBAm/4OhiLiaaJ2eXhPLgAL8KYmwXZAe73DHshl/SDttrz6GVIBzckfD0CuIG8t2
/qOTIZWvnXvGMSgk7C80uBnMd9Oqp7ITiXW3xIxXIV2/eXx1MltPQ5OWhdHy7Ai+
iSD6esAVscN2hUd3gQ76cStlorwVpNTZswhLHN1VeZ4YIqEw0x2p4g2ziOEXDHEN
8sfi8ENkakHYZ45KgF377FHK+EH2Xq+j1pHGZiPKYd/cjE0O0oLOFzHjZ8hYEL6K
gU+crQYJpFYuR4m3JrdDWQlvHpYXw88JzM1XG0V775VsChAyVPVOxbBRg13Cafxf
Q74o5kkRRyt8iKtDNpjgEJhO42trT/3hG9gf+qM0xKaGogFBigjUELn1xzwVFKMD
jvgejvCeEUra0qQQaFYF4wbjIidXaBoJk0JqPxKrtAMXgtKHxJ/h4L+0FGHIh5pz
Ms7F0F4SZdfNegq/xodM99Xa4SXifMUJ3LIis5My7TSmKvE2xcIBJ4Hh5c8jQPpi
yZQEPrzrY2+9d9w5lu6iVzGuEGGvrb+Gxm3BRlmlfItHPPXeWZpr9JkemO0ePd3f
T1bP3zoi85mPtm7L10q080wQ7W1jrmDcF3vGRRdYNY5m382wYlwApu9qoJID1181
STvIzEo/xbKMjSsecH4DFEOSoHAFI53bQqqhfccBnEc/xsSf6dKt+car+GSkVdsF
OqQ3xyna0Z8YgzSXmxVvRRvnMvYeeoDIt0C7HDoXj6n/ZHgbq9NgsBO0HIdWD3Xe
DLI+8AGrjAU3rbTuihiH4Y0omMikPoImNjug//X7v4MILl2tCa7KLQ6xbXLYET78
O0sFRdtSqMUj+vyI0QJEnTVhH62NYf56R2ae1Kz5v7hbP9fzSzzSQwn8/w9xhta7
HkIGxCPVQLESfcCnkPrjh8DwnZcAH6K4NvG0ekKP8XNYq1CPz7ETNywmrhLHr8mo
1HKmnKrZuje+mhjbFJW/AVoZZgo6a/CA1k4OyqqQykh7jNQKN31Cv0is+dhMEmAO
u1woYI8XPXeip4YdVxqPT6Qp4qBncffLThPb+1V/CxZ3wd6zjd308eYBzdap2Thk
9kv4CnPxCTy3fC8D1ikYicGb+aj22bvwkz9DafWyTQ9kSqePB8ZojXrlBEaBBQAV
2q1CyvEuv+opmcosBCm1jVJDEz3tzY7TJXLKLinoe9e9O8VFbHWEtsGmmeCYh6oR
V5yeJN7KdRwLeGxtLsaSkODtGjEPp6idZdzNpjcoJygQ8hZ5crwGk9PnJ6MejW1b
pox9fhAWQWccbTSmDvhdpiBtWbroJ8MWiea9x7ild2BTjuhFw0F9mOhR2BAx6gv7
GHXNTW1PbM1J+ceMdF4j9/LYzqT40hZNxfjQ4WaN2nL7gI2dw0b6cCAKjnZZZHFt
K1R26VFwakbm0MFexIeE4/o9d/T74G/1PlcoC0j/P3VU3aRJa2qZoWV15yTqDALT
uT97JIowmQKghCWKvPGDxUVr3Qb8eAdWAvhnXmigLybnfWBv8fED+FmKAYL/8qoJ
XWX5ezbb5dQcvK8x3djXP8/6vyWOx2h1GkaAsz3cWUo7nJbJTk1euNlmeZ72ja6x
wbL0thhMMlq++dP2suXg8JfFwiawonT6VIISA/h6aLJJa6SLRWBDRdC+6yn+F5Yv
nXKpqkJ74meXC0WV8fIBl54DlFp4ajvIHqzis7urXdOIpJBSBBNLcW5d0FQRbKXg
uy9ypuyY1gEqhLyyH4gBv0UDfDkcc7SWBRmhJxMdxkQEFvpzqLDBWBEW4trtiWTI
iCDZk3vs+pwiF+jJkTFoWnOW3B0lTS7/sOLfrP/ugYwgsNm2HVaXKoTHxFqLjvB3
IAf8VIJcuVkwa1ReMMeYf5I8cTDtVe47qSesBs+3xKAq4cTaZ3QIWG0a0NaCA0UF
aEc1euE//erw2PKt6LZc6iDf02N/NDNilkXA2c60y6u3o69rhUkK50WaXQIv1OP7
PKaP7sQnML99tui00f4x33vh9Kpsgt20x9x981VPJbTIgnXeRQxhiIsoJ6bjuj4S
Nm1IPVGxGyoddYjnCw7VSlXSlki/j+2KDrS0lY7rFFz8qTfw20R+GO6UgoPV7tni
QchF5cYZ8S9rfeDlDs83D4hboHtlIOWmGWPpjRRjMb3VDmlp2QhAkt9SApn60/ke
wMbjr61XxYVPohZjE2nhkDQLUuwn5v/w0HWbNDa5ZtoTqpL1sk+1v7rpQwD0TdJQ
ugtmFdQbd4hcSW9XHHAN2NiMNY0d/D1Ppbwzfte2nZ1UnnrGdvqQuEcPjw5rpxa6
fTcBI5h9bu9amfZwndHOZpgbMw/X8CyE4DilFGVN7ypingHpl852jxdbhuNQkbt1
bTuMShTci485hDSnraNE9/Nhr00YeDoj6NpomZLp92V7EiO9Ra9WbrNdr3UMCVxX
6XI+u/8UqTvb80xZB7HhoYC+hjon55RoJIQZHTIJmyd56RzI4NN0234MMKsFjI+s
BntnCimRohuLKHE1pfSZNu4vEyGfkLJ41JWs7jB7yYAvEbDkt8qFyRBjXSaY7Gq4
dA+mHX4e1wCGUY+HWvi+7Aok/+VxG21GLrdsoaynFIVwBRXR0JSOQVxxqRm6BeFM
XnsObnNMcoDOrPXSeMjcLoInPupAqDpo7vv6EwO2yo7vh3dt0HulZI8OPR+56ln9
TeU3G60Gdu2VEgieutmx+LLb/IPKNS6RfkcE7Z8UGCWEDxrh0or6NXyFyZIQJ7wx
1gxjaProPMbauzMS+ln4XQzyAMiwzo8DxbD8OUm56sf7b1hkEs4R0frC43gvqPjx
CssqTC91/BQ+19IojC4OqAwpT5xTXLvYhj4/SYXO2mNdP8caiFSVcbI3++Zic+lG
xoheWzQMbfyyCGAZcNF5l5eOAO8bIIf/q4TuTHlUZANkE3/nPzswfMKT7RHY1r1s
6iJdUFJX7NSuhWngSY8A0LkR0ibvsb4jlmXrqU1axxCEPi8HVoXirzjN48Cz+CLD
s97tpUkLSghWGCZCDy/EX55E5PC0k+KMB//11MIM4UZ23GEPsUQ2R9iiw3Iuhs1Q
qQfqHFSiVMuXI+nZuhOZy9IzOT/QgHPThGDAw1pNdnjT5ukFiHGrhrBPto5C3Zx+
3rncuiJnMxJ1meeLX6dl0c0v+IfFSSlYtDUsJ2aqygGY0Gw6cdwlbvFyqtVCs9HZ
KCaiKDvNmpWELM6EZ5hKxDBnaw45djTg3js3Gpm7zCPEGH/AvyXrRbx1rBJCnBWg
DKhj1/3aJFypd20HUS45UJ2qFxjYcmVIpX/P6iqn6ZpEFzuL+Bki7Vai7jh2LixX
UtJ0vjrP40L2TkMFIWRsLQ7rQoMNA9znvFUD410NgOrr7M8K19YOh2VzVG6ygTDt
I5cMGSVy2LuxX/meyvJYsmoznUX4Z4JbkFlf72Jn89Mf4nVgHNsRdWMhiWyhb6i5
OBnwn2IZKp4fL2wWCAKaQo2ZYXdYluONMZSxlrUlaUaMCIvDnYYmsPKKVOiiPxRR
WvV8cy2sYx4Ty05Vz47tpds6f5h6bTRu+n3exzT1Ef5GA+MFIU8JE4vWVBsnjd23
68QW/1tb/gDh803ZIE8LyCuy0zMIgcqzjI5taoc4u5+LDbBJr3YantFeq1poJhNX
8nMoh9/V77yLR2QNga56sKGTNV4jBkskjuN0/WjTJo/Uu/v8azhu1UG1GCK/SpnF
8EDBWB7DuMbYjz1Sm7L4/tPtVF97bEt3Sf6GhUMlRhXKDFsF6g3odtxgyZCUYVsu
fpyJMBRDyV/cRGK89IA6QHQofbfcOiE2wnt7FhRuJiY6qakoXRfNygsFkiM1AVq9
98mdrJBThsXwrd1v5eXjoehsGyBIXkKlMeZ83XY+PFQbGwb22gd0TrzpsYDKO0LB
55rrxq0g7LSyceYXv2oyZuq4yRrmkNZcl/OIxZq52mr+auj7Hm9sR6Q2002HDgeE
0xv2nD7jRkQIj9aJHF6Qr0d+vdBy5gdQNf0K1ZWEuKKjDn8YgZxoUf1ydZF3Eyqz
c54oide11MulqAiyHYIHw6raSM1tZx7Nru1mJ6Qsmbi0igXEaX7oeIMJB6+/KmJV
lFdQBQHCCfQ8bQ5O2J84paSxLNFORgH4UxYxyHzXyF/qFG8CMgwLLN9AepTyEO5Z
ti771xIMzNiHy8KGHaojal+mfu7EghnW5B4gW8zX1ev2++Zde+L/u/gVDmzgdLZC
G38QYLvhfmq4azFhzVau5cND9ezKMfgo0rsi+ABNVjcWgWALJ6NgWmpTzch07JC5
ENFvobRtvmB5vxrroWeTKjI010AN8ITfCtLBmuTxSeOYt1eH9g99v5bPPMZFBDMM
btdnI30XM+cWUy6SeFjegi1rpid4urLSu/RZpLHgd4gZoDyyoio38Xx9RdAOqGVz
L0KvMm+TqN+fWkLwTpx6vOxVxCdiCoKTdkyHVW8yA4b4XFA28hQ1bxH3cPkoxCYs
rQeLLOqMY+780sThnfK5sx+E0xS8MMcn9IDKyHpvPqdD92PxlPkKykr2STDQ/jox
9vPpUR/+BhY86pb3R001Pddl9X4Q3ijteXwbdmGSjZv+QrlbIMd6ISNYEOUMPYF+
S0vIxYpVz5kg8/0d6TpbvJYcJtByMQ6LWmNNzYb22dA1StDp0WC1ufCBBRhZBd8y
ZfHsq5+iQJ1ZUcZK7HMwlU+8Qmnd5rVOAtkqNm3jpAU3dwy9fChNw/8ELIhSayBS
1iF0CkCBsFSR8W1GpXgOyQe0oEWdGgoZAnzPYySwc7Pkj/1CiS5j8IbNzznVn2c1
i/S212pORte6RNDDLRagLg2PK6Zd8euFfRYtrNz/ABLbtqqiVcZXIA73ceBTaoE2
FXNCGRDzWf2mBHpxCXA33P/lOiy+Dh6oFp3FaVKSrfznVBQcjVotynHQNp3j9jd6
YeZpZ/6zngdMFpJUrIlAJidC5JftZy/mvrUwoORDXVYknwsBaZJUpqZeSq853wl7
0OTdryVzaV7R5jIZFO9DHhqdVrkXrpgMVQ6xJHiWFpr6Bzt8T9uO+J4YoGFwQNjN
63lm2rpKei2D8mVV5oEFbDQNxViquyvS+tYd8ra93vdRzL/s4/DNwuaaK0aBfwXu
PxajTxAPNu/NFflgOEWyfomFcKFSxcQ4mxUlGFHxERt6fnt3Njn9I52Fudu4IPCb
VtOHyUZL9kTt1KBNvpYjPAa2JB6NusalUJMTscz7YwR4rq2HdAThTO4znht1wSgt
exwoiSJsdNz/K/bA7+ePQOM2AWHK3UdtU2LFG7SR38lfZO8nrjmXtZTlqrxOSmrB
N543ahPpQd0JqQoJ11DL0Ch52xXZxrj2tfRw4LVqdKzRID0IFpsYZuXOmXxhTTXX
0OI5I8LCOHTn7yR31f5jUOXqbUahY7fADQbdAjFGxab5nTy3I+GVUvEtYi5fgbGt
TvpWNqOitFpbbXPmHKP60JxqZuM0N383/RROJf8ElYWw08oI5reph0vwR1X1jyEb
vpjDnqh/5EudOrsXoCZthnNofMlDbQ1BVqnPVvC+h1myRL7XFzrF9S6eUZS/XEK8
wIhnMqmEUYk9gPlY3F4DnnORStq2uBVW2Bc0ssfjOKbHiJX5M7sUXPCBNqieCyEB
9RU2oI5MA4jhMAn6udOjAvV2lSmNnsBBDXK4iezRElDeByRMp2SgfgZUomnj0T4m
7fd4MaDjbEIuw4Zi6EDrztp4DH5vQmt0zMjiBYZ3tM0rsyKdL2jn/sYOsoI6py7u
vya8F6B70kKfeERuBHC36qtN2z81uL4M2xGHFJuUiaAr3QywyqchqOdOp0QZpS73
EjQTeZPj5wirDGDDD4aG9PDMXlnv2LT/e71JbeN3NwM3DsM7m9dJJD0KUHsP0PxV
ABuI7WDmFiWZJJDq03MPuFVbDPwuxvmOyE05HKbrt8fI1cKU8JRN/e5b2ZE27Mus
bvx+DfV8SUOZhvrv1DYHycm9RBPXnsWj1UUtyWpD7U7gQdCKFreK+4/TnRk4YLfK
+IwN8UKNCKEZDSFrMMNEA0mxmGu6APBbv+TnVCGTFl7EJ6OwSVwoRn3k4GxcwId+
GzBAsbRcnHSHuvqei1Zt4TL/vxdcDs7u7xVl6al9fj2Y5oDEA+u9FqkUmjOvp6Ex
fkHgloBiujSgXXgXpaEVI09OiLcWaP3CxoPlIiDZCfbDz27JrOjK197Dfb8SpVvV
AN/hyx5Lbhm/kEzJnGjiRC9/Nr5FPJKacOpik8CHI9RL2tgpGpU7uzJTFDqEWw0t
58RxKsdSA99qKqpGqqplqZgEoKCjQ/4gfxkvquJy6wj2krGQO1ai3MOYEfji/R0G
jwIWQqz8R8pPAvrLSHo9m74jJO3pKU4WRP6Cqp6f3OJXlVFRmZNO1ZYyCAxW4MJ3
t8cNOG1rP+4UBpGg9MMg+Ww9myEKU2XZOqvQo7Vxb5HEoiZffe+Pmp4Y80W6c957
rbtnhi47nyas75y52f2JZJtRHiu58gCyXBukDRCSk1Jqi6yhzqcTH+8CWtVEgFCS
baQN5d3Bu/4Lb4wlGZcLYrJeQD9iaYZXgUmvTr2cL8TJxbwz3wy+ugYGAikrU+V2
ZG6QC1qA1bgxhBKkV+IxWl7kKpBw2QqFJPZI4UhtINdntykamjPiCHuDBnj8eMT5
kL7RsdMLzB+Gj2CoCzrmV2F+zxx2Zax83ODkizIwO8NzS7hON028BTgcGfuCLQT9
BwlUZKsWQIbr8kiNd2a1SNXVXR9XwDMqVxk3yMtDTnnrBrmi4rOK5Ad+ScHH6Gk5
g1Polw9y2EI3zVTHDjWCPza50zXN1pkuUE0ivDCltMoNhmugLjlHY58chmeeY1yG
UlU2o3U0VmtRQ1g5SAnt7qhKQ+LbHiI6D5nEd+k3Y9HgmKNQIpjOE12WSnLUsZW+
0bUwUHg4P11FCr7guYJ6wihPRRwpq2OobIED/1t7KFJsHx+nSW2P/YuFvRZRBCtf
J03O/1XKw0UZnrqlACGof1iwV2sdsSbr0B5YJchrGv5xW9TJUfZfeG1bfUZoyZFG
CgkA/QuQavwmRPCCfc3NXNYOKNVlzdTp6BcjLwyFJvZpMusdN4XoIoFeUCiicfSr
O56tYEwBmQmLRLgYgpf6Tcf8yR5OnL0oTUqZN6xDAqCROPqbExxZbboZnwwPrb0C
e+R+dkOR2fsaz5RZJiguraMl3wxIpdSVTdBmbOQ2IkvzwPW/Ih6CGQHTZwQcJu4D
pnnFHbsV9gLTU5sMmwckiyTgSobdL25kZaBVlXDPderrdyNtbN1NSjPXq49eLSak
mp4quihevtgqTqIkqgnM0jEW/ZX8vlWx//1jzCsr1BODkbHSFEPXMRn8qr7hkdwv
pinvlQhEMPgXzU9hxprkIjiloqbDG6jV/Tvy+1ycWpF6W1XJiT5x/0eYw1/Seo6X
1M91xUMqxpHTNrlRBMJS+gGnTYjNJE9rZRPDMY9vM4E2LAuuraUDYbrhNHyax8/y
e53qBslDptygqu/Mdg2lodQgY4IfT2q805eG3kqUXs3R8Pu4HdtGD10lGu/HOlln
QNrM2HEiJI0so4yOhOiZcVYDMCXJ6b1bMXPu/XWcrPK3Z8/uwn/q+X+bLEIU62Dx
kZYOyQWOQbc/bQ86mOjZ9CgLtSTp2SuTKanQt4Fiy1vBEgkdEhFjJyl9OqavtsXf
iEzpnziEqpoiW3xSos4G3MT7ErHpbBOKVRo1nRqHP1qDOwRubf7KkyV7UwK2udJ4
rQM5BoJQ82nsoWQJGJ3s50WNzofi/OXffIWF/7vQcgcJCd6Bd+ZRGB1sU0sXkFbG
ZnzPvvKByFxQXtaKKo4E4v6pDyK1/cDr2odcywD+ub3EAWtnfvxSFZ/TYi8xKrZD
EignnVeXk9eZE00C8ZhKscrc1WZJaPXXa/IuSSfBMb/ErV1fgI6VlhaixyWcaYO3
/9r7nSmeCu+koxhzxTxGYz43IULxyigT30vpNoD+IchOc4xwCQh986auXP3rHyHJ
3Th7Q++bJTdNjIJSyBU3KVIU4z6oiIhcygG4/BLvMshrwS3t7AF4D7lZXyG7KM8u
vHrbkoAqwH3verGHS0/EKnsVIT2Kqn45nntFXwaJMmmpBDSDIyBOS+jZfARZg6oB
lHLn3BEeZgwyEJhDuaJgWD0EtGZSAYfcNtszvRJStKGOeLkFFqrDYQLyfqEwWqgW
G8CIg0dQ8eZ+EcZeWH5Umgj4G5QpA4O+jnnduqdU87k6fpg7ZuTrUuXQbcFPM4Fm
4x+bnWYdpOH1JFbbwqP+Ab0okskHxIWf2dpKQ9A2oUHi58PSpp1wZsD9uRU3Asgn
3/LU7l82aoNxSnTlEjSblDZdq/1zBLLDnrPnvQfs0G7sScGwwtzs8X14mgvoEb1C
IvRjGeR3xWQe6piyXa8CxCdbtd4D6S4qjpQwp2wYHQaFAvPtINIrty/dxY6Q22ua
0zXDCnSr9lyAt0OxwSG4F/FPqJQpEk8tvW4mCoY5nf4bWLf29jTI1oB4ePq1QiMU
CvJA1P/LED6j4a/mNHWJzTRHodwgf91aVi6KBMZX2eQrbDFG+lj0pLyluqQyLRjX
4XGNaUpP2rNZFqrBW8P0ZHHmA9q0y1dsEBE4xQwpsOYSGQtEhPNCGntvi8Bl6NYi
wFhe++TkRCKUlp2btSvW6Q==
`pragma protect end_protected
