// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
FdEEwgB5lHKAFop4B+5A7oLsN6r31BNZK3cHwl+UZxM+3olqeN1tmzLJxnl8CiXEUtrOVN1fUq+3
FSZFfEtwhiJWCFQNIc8UOIZpFYZPonJNH+CO974oN2rBm59bDBIVr13q6vcsUWq1UI4FSM5TJvhM
nYNIovluHkehQJtPXpJv2y2/x2tibbMY38fgeFwx+Q0SYWjvKUhRcJ8YlyY76fbmuPcehImv1vTO
dz9ePasC3p+LKO8TON6YAp0mOBJeB/O7IanMAwCNSpX11v3/mUduysHsYPeOh6gRoSEaG5Hao87Z
L00etW0upndfJbWcJvn4iItsrKAHBG61AQLcxw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
XpHnFOqfro98cNCB7+relSpUeqRBjB56UKWFxo/uV2ojqFceI06UZgfz7Q5L36I0LGb2Hp0MXwSF
sgoVDLl4m26fW5IKh7SEGeCxnGHwJ458Tw/eLX4eiDoFHny/w+7Ry8PhffT8vpmEyF1RHiS6L/tE
rANA/O24CFn0WqpOP4PHOAeaqiCT39SQcduWzswMu/QZS7eBKHpIvX4czsZxVvwkUg/EKYKYgJQT
1fxC1nSM5ZoWCXmgVXcpocmRySRSRyqVMavgIVodI5NRl+AInMsTH4/RU+JoTrCJ3/0njgWF16DE
Us9nLEaBI9sqGQ1xwBNAEhI981DjvXmfjH/P1/q8G35eHUrwG9K9rVrgYpPwqsUWQZuc/HdSwjEb
G/T2W9p5NhjBtODWwGjbKkM0tPFDtlR0Ydhz2Jh/jCgL4VmYc8VP8UlG0AmZQifVw/ChxdmAIY3n
Z9iC7w9Clu8ivv3FR51hWpUdGP/nBBZUq00wjH7Z+gJbZQpfsAH19WQCKd9vo2ickYdyO4OgsDLy
QAoEwbNpN3iaMPDINrIWzHOFYylKBD8cjtDVShClLNaWEPdQBrYj6wKvywpAjw9pLFtfYXPSeVL/
9HDl4cThnb0TXsdOW0RLXCp2kP25qrr5zHrvDmUeVKRRJFZgyOEdtssOvHGHxeqV0Z9L0bo8KoAc
PZ4nBROuMbTc2VOpoA7lRHDtUmR6Lz6ouGSSWxJYsXiseH8Jlse/H7jyPPcbA+a+V/6nvuYbJAjg
c9ecmJsLLokAK2d77+AdKd6rrBAnGubrBhWkd0Q/N5/RQnNqE9dWvkBiImX3jPc230IWfhJtMfvH
Wq3RWA/cB0vhdnmuaKNsW69eMzx4VRy1DnbFgCCcf4go8to/j1GurOtTr1F6ZMPPSTI+lWY5R/29
JHKg6CTPRHZ3dtQPst4p/380SEwlSXYE866GKe9mBHzD0hkA8FZpHMbK1xI5TYYVItSRhNYmR8q2
fAkrQABXanb5Q+Sd64aU7ggiVYdHUeIkHcYRt71GsruTZ26p/rdvhy5ZUygX5QkJnCUSRYstEFBN
aRc0yob77xkXCC4PzCq0qqgMH7UhdDiK4E9POzf21UQYjjYAGZtJr03Gio76HavDJ9k2tHR1mlPH
om0rFhNbWVFDYqURZfhz0i3Yx1y7nXjEMenjn9HU5LWXkZgxPTF7E3hs2JCz0sFyiQUxhQIbqPjL
1DgoTrys0KtLLsOdEDs/JZZK7cYHhpPE+k5oFXdGggXt1i6DltghQFqahcuGfr0iMrgTMSQSfZpA
Y+9bHOKfNg2POdIQkPkI5zyrpEKVp3MMP2t5C9UmSd+6rsrVFyOKIrJ9+ekh/sE4Em2tPQTY0mYO
RBOFPfkX064eD/4lm0M28lLhKAwAcWjQksw+SUCkEx5g1Q4tl30tguSPq57FVk5RUC/Y35Bg+FFy
T6FMYxW+LDpknEcaqPT+6T8+nO10YQWvWYD33xsVEsLbAOJwcviKvYaxP3OlGHkii0a5kbvS5weh
HJFJRgnfAFL9lz6tFdRfOm8Bs3RHrt3haVT053FK8x0o57458B7XW6kB55mIx57nDhYFUssfqHBW
gdJCGpR4kkAsohFeTODMMslWqmS3dPUAwSU1RnzylNpQxPXPNzJwG0bAr9hlFQl2jCS/BI6w4W+B
8WPxsa114WU9WAbAyZPPFxMPSu3UmXrVbkEGlx135o6Kzb7m5ckH1KE39Thq+RICOHIFwm/ieWyw
qNE+TSBuE/+PxUgp5jpJdQNtDT1DWwmnDjpENbWoikr3WBWrRjrSL/mgBRUYekWz51mnVGDckeOY
eehR+g9UyQDDhdSfnE1+da0nF7huPZT3XLLA6xROKsKUheXIGM+KkTpHezi2XpY7v9G9GKJDniTo
n/QL+V+4/b4Hsyyyeth5Ma+0SdYMrASOuyb5WYmvmbM5PA9Hj/tkuoJkozjlLT0F+/V1/oMLoTci
qbnbRt0iBzHectABnuuieeO/nJYCZaRQRf+5Lp6DPNmD0bsoSmLwqt8JBdQj8wsL92lCAolXS5al
Q6fD36NFV0JbFlhcU9h1yq4YN4fbVDkxbGAwrocTbZ0Oe3svBiNRtVxU3min4bM2t0V6lsMyUTsV
NlDGjhLSq+0oVweb9bYR2bTVCgsyC+BPfFIcb+PYGbWrlYMbCdf/bwg4n4YBIjbH8cR1iZqZm2aO
0FEBReWfQ0CtXfA4ZBfhEMTY0qXvZZWJ9ZVrfY4RRqGKfN+cHD+kTqZVhSyXEEpnKuCR3almV8q3
bg3bT60SBlZwe8YzM0mWnbLrgQKTKl7pl7lANyIH7TO24Fz8oVSv0NXa5QckU6JRoZ/NmgLXhAz+
yrS7SxBYooO8kF0oVVOfbB8HZAtcw7E2mDuZWwtTJU0oAEV/hpZD+SGRH3sJiY5GMVShURJZ2yQc
tfItzy2i6YwdL8msWvjhX2+8DsAH2FjrQH9JNWvOpoFnUG1NnZg/mBxEbP8nmvT6t53HsBwCGrsP
qFHGbCYPIFEyC3t+6GkJN/1FM0KvFXiPoAB31FOFjpc5QkiZeFZFRO7hVIVrAgAThOkzj6yGEZfs
d0TMAKtjkB3Y6H3+JmadGt3dKESf5RtRDrNeM5YriW6RgvkOw2jfynJdSbydO4mdtWr+m2Ucn0u/
yMYjIjo8M6NenzJl1Mak952vRhe56M7mJSbJVLUCIyyi4L7jRIovkH3sKIRgovdw/tB06HWBJTvQ
nIhG8w/mrOcAn9hU9eCcDQRA+eBAc0OlWh8xrTcn0R4twSlgfGGwott0GWLBRTWeKIie16CCH5JI
2amXdUgVbYfy7kSy7q/ruwnopKuM6vFcwz1zgR7pAwOva+Z602XnckVtdFbXn5Y8BimnmfYWg4hK
trWiUG2e+mNOg8ko3qulpzoqyeCSjh/amc7lWaWb1UW88P2GhcDQKDCRrmR3sCwoMukRRtxQhFTi
QhSX9wmcn69e7sVtNvSb/FvHiZE7BjKJd3IZXB0WpEAbug3R2JUSm/MO8Zlvbqd2NPXYvQYsh3qB
wxm9dpK6eQJtIVYYnxmeZwVU44mIhuDedP/1mfOaLVcghumtyOpmZEcrnnZ4dehpJv0a6E3exkDv
bJCT2T2ODihECoMBQqlk3CwQRasPkPVH+PFMoZWtRWmgA4APE635oTlqZtNdNx+kt9kQVoBkxHdJ
lo2GM8rrPSbzBCSDBDgAz397w9brUSfvKsj4vOHWJpBnDECJGQZ/FsyelwNRMw6i6wnyxNMD10Ww
4TaGiDdK2XZ4scDQJgAdYMXE5q4ka9XmYUYoy8iMXSRHIEJ0ZyK17dHA4hLDKzUci7cFNl/At0mC
RBCPE2y+fByBH2xLGBgk8Y2qOGVAelw8Hnq7nxXlhCAvI+zOF7Hz7wuQNq/dfgwiUAiFVZMVus2n
5D1I/RDyusWMpKjfnh7NVonoHSghyFhYp0cG25XcNrdADqQUBQzE+2R+ZJ/+acSaECL/ModIxtRb
NILAXpflCSiHl3JKY08Flxd0MPL00KkUSSDBJKwLAikG29EawC5IJUzoirTqwbXd27AZN/5J5iWd
gTO7XNzxkWAuq3LU+lWEPqfYII9RswF7x9BoA+YgzG31EVqx7yvxIf/HW8WW66fGqk6xZxG6h7dr
Sgf7l+GY7hDaYnTFv6+Tg00x2sPb+ZKAHhPvabjIt1HZFMfERHJeRwstmSjerTlwno3vuHOZgSmp
TxhoxIWgWhlOYEQhvekXOnjph3hxMdsAQZ6Ju0QiZoiexfuIKjSkRIzlc/ftWeXs6Lst7HLi5G5m
FgQHaijASESejW2uPXEJfTc1nmC7+ciyaIpBjEtRc4RRCJrH14CrZG3DlddC2e2M6dlPFi8xXp+u
pSYoisiSE2Nx5Pmy9oQSmRDLqdX+1i48VRKsRCLz0oOBhR4Ha3S67eE7W7RUGYhhNyRJwvo0tobF
GcFVADSPdNP0ZfnYd41QrryqXKlylGC71/J4WicahC5n88Q4t9Hbb/BYAjXw/uuso/m7qmljr4tS
KPxfZMZCrLwnFPKQT5pyNNbGRVpV+NoxT+tYoTFj6C+DM9COlKP4fZXJhCkQEfZVs7GQFBNp9F77
fZKsek0hGxVy1wkGmxdcnZHPcEFYu6+gxapBlcjHuw0QibpgudHtr8tMRAb3sjo2Bzlneb8oXk2Y
/ZBBBq5o+FZnvtg+iwxyvyzmkq0T9qZsJHFT9zxXZNhAgW/25h2Okp1TLKubtPjhvd6LM19LswoL
J5L2QwjSALhgKruhRCYSIkYH/ohqjZSUcZOwofEDfDDQqP6RrM6LobbNuK/8ffjbaiotai2jnZnO
gFXigB0Qw/2bVSO8zKZamFYQnh9Y671z2RdGi1RaU/f8RQqo8VM3L9r/nQVrB3S8zxUbYhTnFULG
T8dIAtXr1Gt3gEvqSamMdKHUXlPggS+km+veL8g/wfZKzFWKLadVEmE3ZWZeIPe+tbi907Thb20n
jzt/vpwKlNcBlj9aQ58Za0KzU8WHco30rEZlySPl1X2cI4Iv2kdIT5eijTpD8l2tEZ/1pqvVv6Om
36iarzkasRIq6EXr2d81rvk1EdoTSEl8NFp9KM4vDH5fRbrqWwRFpbSLxoMN35vkfhgt9uVAkEdj
YL7c5W6GFW0NbXKD7jXGl9wJdHcBlKTDBnztLROGptbefVo17ZmKWqIfVEP0JjfVTR6dORCv6eFC
DHg4eAs5sKA1S2dQhj6GG2yjpqaTkyosFclkO8wcM0EjSNPDP6TW4njpvmn/52L9lPEKq2kgdliA
7UjMyPoqIDF+K3Zfs1/7cfpvyfZf5kPrWnfIVCvjx5i+0nP9OiNZbm6BF2Ph963driIJKxXVrspO
8QVBHWGToj59XI5uUWdWeDYrPLyk72uE1VxoOTDTCYGjiSRUiYN/l1vslwOubxggkKxU0qPHJvFM
eugs/SOXWvhJ1AlhhpUj8I+NZt49DbmQ3HsgtfuPLq6RkLVo5cqK1JlRGbFfi5lbBqy9nOL2TAdV
hPJEInR98vuyQrXRb3QxvDS+BkP6jsCUm9I3NmzjF3UmgLV8AEBA17iG+//5sSMT3sN3puHh00oO
z0Y2QaVnHvbzLqDk6TmKFGZGymq5KCZ99T0GYXhQ4ztazC4w0yRcsOnhRXDdmyc/UUrOoxNgWxpK
oGgn9Seh1SWzDkTsc+bhcFHGXhsh+mTKYD9MZaACZksnm7tu9S/wPRCWf+XrkLv0MXNc9RLfx0Rj
vrXQ+hPmZdFKg4vxer3mDxN1lb001ARpdNADCuBr3TYVHzCsWGP+8fBQRZj2uWm/19Dh5ah9RJ21
u/CceQcWUynsQooGxCoZj7t/ZkQguCHIA2MhMc1elo5ZJEo+G14pZKOxs0Iu/XuL08hQZRQon6MR
VGVWJAOLKET9B1rCFB/YesM1IrGdFv4dleShBVG60BiWb57wFIcKpAOhDSgh4C5pU5+azpL9AHtF
43uXAUmW4nngqwsnZrmQU7QJmVDWnr8r8CLu4nF4fQlfgT8Jnwtdr40YFjbNeAEZJlpWKj3HEU41
QcYWuq44GuOrgA91iqeye/HYKIQxODO9sBGZv4Vad/+tyP5ja1sX1LaPixgjMCRAjJJ57kxlY76I
5ryrge0a5CtJf+R06FDnyjBlgIpNSFLYTbwo+rc3yEE8KhCIPIhRnR/xGLOiDa1vcVU8Boh4kN22
Aou88lYdGNcu3rBaTJcB7YVaSVVsYFm7fZMjMcVc4IMmrqU/9d4prOWK4u4V+U989kJqAiFk6+ga
sPeRm+LW34TTASZ39USjC2vKi13rlNJKG7KtfFxyNQKT4f7jRXNDmfBHbqs0FDhmCZLWrEzoT6/u
xOIc0+UeCG8BgPAp4qOxTeBq7KFZCNpOy2Gosib4voAlA/I6zgJGWR1CH+yYfNmBJLu6IkyNXyiw
LJo3unZlC0vs0M/915/FSvfsT4UTwdgr/u4h83M1rQ2+FzOitjTJrPhw7vfxNm/mo3LVSwx2FI2+
OvviXtlz01l+sE+4um5xO1mywDDDPFKIdMFkjj6RW88Q2D3kNGRTcy5S106ezGoVTXJuVzmOnxKP
ApCuluTJ9oe2KHtxEKIbhordeYL27wsqadAfKMGORieDzWV9FamcBJoE+YDimBpMDECiVAWM9q2P
LkZMU+93Naf0JC0W1GEA00jPXhTswD0Nu+EsecgVYCTzlEK+4w+EwRli3dM4yeNlb+LVVF9Mt2aM
YJHeZ/te8ldW4r6Xy2bD1M63X1z/U7C+t4GJ8gkJ5+lfF1xkqxNSIkGujH3q5cp1FNYV3DsfjkJt
dcRIJneLUyjw/fkMlNUsCfiBveqkbK+K3SIGYEFZnyL6jhfGMhwF2ENOirU2OdiHSa/WVwyIO6qN
xR1d9EWxgTBfuQ2BLtxYpO1XZscaA6uy1KvP5IUzEtQJsCW1DMTidW5PatGKvHq6XuN8wuGXoARv
PiQEOiryvEZ9DHwUh+5xEGunmHWBB2hYBihnbZ0waQjCEyZS6SWFshpssJdelqCJvPB58LjBHqcA
x7bnmhfAPtK8E1S78nV+ryRW9gva4oUD0mz8s9tT6O35dOR0qP7W9qqhLqVM+n8FgwX1/uxfV8H1
Zm466oLjozzFdipHXAXvJqFPcWXctIMyMkqZG8NqIDFYRVbBqaXTi4tABHLiuqccR97AuX8tpRvJ
xMpSnxiyCinlb8epxWkupe3aUD4Zm9LAmT972fPISF6EmcHO8SO5pyHZzsYKhyDqMgcXs7BZePWN
rVdZ+pvgPOLhmkZL6JGwUpJMRhyH7HUd/y8f4zMUrvxL2Jb8P6NSyhEJKhOn4GVIuIXO0yev16Jh
JXBBHX4rGt8CZHrK3pKvvjRc0nXwHwky4AXOJGlmUl1wt4R3j1RHEz2WS7zyvy0ag2EhlGzUyopW
RQmazKFTy0mb9IZcY5TqxnsS/FRrapXC228mRkznwHJSqyYnK73kviAzvZX/oIktwprwBfyQByVq
s1xk+EBqyzkQQAbYdReQYMxIk2bKTZ5XelRiymBguftaHeeJTO28cQMLLcAjzyvxHYm2NBrAD6ZW
KumTEbAN2oygwRIfx7OSIlan+yf6RDyRJPGhcPDoAL4rrCpX1oUehNDVej0cBBarK99o1fC3ORjr
R/csXFEVELhNemhjzR9y/ZI0qfBx1PCIedKJFTO6T021Ew8/IknLC1XVxEqcbAdIkZjM0nrNHSXE
nmmOq5QY29tYONDVT/d3RiJ5PNF4LbxWWVoA6vM4BdIMK7Z6IAeJa4vviGoDdCu9e50k3F9LTbFO
1dP7NsNm+PrB6MTrt3yrtQ8ZdJPEkj4YpFFhPilgc+BTHQY6t5+LORRGR6FW12SrOqkZsDHwaHad
MJLg2SCaCnJtDVQu5xAHlSeDr/mcbIFP2LkDajZ/rGYVQPLr43ULt7kzhjopP3UYpaFqp/3y+Kl6
pMvWwro2Aa7kBWWXIx7bNnOrKXtdEuF5SdWlnv9gi7l9iuubPxcQFYJyGCh9VCFcBc+6HMyZ+l38
/WJUUHQst3waPjv4xT2Ab2+rXFybdS6+jezD5OlTD84tzuLmi9psyFeOi3PRs6inG9zllkQiWG9t
eR2cEz+xDormdGYIit0tiOs5b2tO4PR1El9hoQQBHl+JMmWnZIkPibMgvut8OjaLT2oYQ+nF5pNA
lT4i8vho+iDbqq47h/kt+pPo07lQ+tOBp9eNxcfnrgltALGJCTg/l9McNw2OS1hAhWtfb8InwRHK
vnZvaHUUeg7HZa1Iwa6hsEylvVD0kPzSgXbzUPitEG89oyk6XIZ4Mgb+nlun7+fT0UQgXJyr7dy+
W/qoGHiN8R8fEoR7sxGhwe8zOgTY4wMT9XcjxW8wfIHmPDS5mrXHSSKtNQkUyNFwNkn8dsRXO0r7
wsAQ2YYYCeWYxqMKSAzT8NS4VD16/q1NwaAGpWnpw1bXymW2Ct5723Z+WdbzbQVj3QZOpqn4hkRE
puKa3fE+J0MG2eqpuZD3m8KaHNLqg/ogANJoFnnasHjxts/uSu94GzqoWtRyXT7nKOKJ5yAtePDt
liGyGtsZM9EZ+fIWlwUXX+4SsXTzRXVyBUBTONMPQNKblSinQi713ds3dyt1XxWyo83UeI8QSRUw
B4Hz8mtgLD9lQVfAN1wdu7Yl3VZDdFioYd1K1UX3RUmkcwmO+Rwwz2zqyYxIOLs+9BEobq4A9CIJ
vWlSfHiX+xU5o3lAqWfutZKCOrInNPRwK6wgCj1MIqItNCw4i8RVTnzNvaheJFkQ+LQ++GTAKeyL
uzM1TVnGtUWxUqU/fkzIC9VR1DGGIQlSysjXRnL+UV/E1HwvEEdx68PW+nZ+ySTJEdlPiRz3pExx
Xr47zsGOmQQ2s3KQE3bNq29B47A8ZYCvLQwoovNePf9J0uOCCmlklhblFTNjgFZ0FLJ1vBrG9H/y
CQhUgpptMwqzdjSj+beMRKa1aGrnsEJfBaHkD8IXrfIhQyE02QZnr3ly3bzeyJYfuz3H4kvJ7tGt
LcCCOqZZ2/9GatTNWjar+MvfST/tMlt+MZLX+9eprdmnGxGZGR6aJwciZmfL97BO7UQc7XqIh4Mp
yZ/zDq5k9E0Ui40xycHscaBEhLNxCpE8kV3GRIXNmh6G6RTDNL+z8OMGfYFPNlZFquIpl5wf2wcU
KaTK/tvwoomuucYtf6o9RuujbwoSFuypf/cq/bpz/ytnduAiIXEFu4mUiCPNIXX43xKqjazvLvnA
55Gg0/S3xlVEvYMUR6ANEYhcYEBbESCaby7W13Mf4SXK9C7TRiKM5d0F6J8IyQXexZLqpLFtd89w
KT27eRhqilxgMqpAYqD6hvyflZgd/UbsNsNXDCGC6ZyuwoTetgIyB1k2h4kM+DT3jGu6OaY1K7Ja
xSckbcY4KV8HIT8ubWVZadv3FJcnCgOkDxgaNam31x/Pk3lhUvwkkS0ZBgJjLn8mlwr1xbTJqyO6
xF9WHVKGytY3vMSj+iZWpj09VQsLgUlctwLDmQ2Wy6Tl85kkFHZ/Nrx9+mZcHCi89cMiRenTa8Ok
jqRcoMoxXewCurn+huIP9gfPIRTfPqQCfom/tQKBBUuKDXrsyeKkTiy5LFg5MjpxAzG9haOmpi89
mb5VDtcl5WlVkORxs2VXiGWophC76fy2oHyhxZil0Qnt4kwSbmumYldEtTnUseM84359mSIbwgpi
+8/ePhUFt1TAa/ZxarLguEKT0qOUfz0C0AQvPCrQ/C79cJhAe1i2aq4LYffJXsefN0yQRpY+ZbvW
ZHjjPzhq1pQYku611TE9UoAfr3hyY+3UxMMOeg/+2GuY/KDkiDi5FyG72AtPMIdmN/oTg8gIY93U
r/DOHLw5DA6HITSsuppBZWm1ao99eTO5WY+76bWd45j1SWzYGsrBI9yIfa+vIPImIH61ZshkGxl4
V3ImFD+Wjq7JaMS6WxFUQwEUlNDSEKAEWFoTGpR+CjQcyu1YVixjTNI67DMd1x+D2EeiZG6myqJ9
Bc8TqUs1dqU3EKvRc4ts919NqStsDcZ6UMdXPomNUXs5ByrHjjjALlUnBGvvYJRxxRq8LnaW02Wt
QGW8iYJz3xUsVZxLBEf0AD9QRTw/hUo4DtEozQ+n9wQaKl0q9gOo02QRVor6EFknCwVxtHz5kfSH
BqHFrc1XKzcQxtrxvBrGgZystt04RqDESbYisxST3wtMQhzG9MJFvgrqopp6cfvJHVpfZkV4UjId
19KIfcUWKkWq5bEVn/pf8gXwm6Sj3AmgHGD5KuoYHuGT0D9C0l+jtSjaNGhYJ6eGKiJW+zMnhOsd
u6ZAMGpiRT627YMuTtM6e19rEai8EM/ZvmcGCy2931GTrK4LjRNxj/XvjpZp7WT7tHR0Y6UaUef1
Ut1732uRdseA/ZMUbWWrU7q2SagUFy36SgqETc7gjB9vYdk2mF9kl/6Y0DOlstsLs3DDgh0C0hHZ
uEBgJKnEnTso6d09XOoIXx4EFANLoEOBywJ7OFI0kxkr85szQbUU98pc86VmDiGlrtf+9XRF4NdP
ZeAfuuCr3FNnJZR5tgJXFhrv5hhyAf6hpf0beKuCJnma9gzRzcQ/Jq1n0L1zjL4YIlgjEifLRhsk
W22Op5YNt7kcrytJUKHbUoOOIC4dIotLTPYj81AfICHjG1a5a7azrJ+AP7eswxDVDuCmopjhJg+a
CZ50Y9/2/E64y+m9N7KbgZC61g8rTXcuOP9qPj/8oq8CcyhyNRoAhgm1iOuuD73ggI+9D2Nwnv4m
5PQVyoJ2ciXBGLer7eOZSvaeIR3ziuR/QhhkFL8dviwdWokhHK1Txxw7U+AbbjE2xNsan3w7+dfX
GwxdVy7d/jCg/9+75a/kKAfBlQCyDR5LoCAVqe5fwzv6rhPykvWtDsJLjmzMr3qoCuVfGmIkwR58
5rUt/yfMiT2JbtPFKIUKM051L9qSyGZnLi/iTlhBI1tVnvBkTxAh4gH9S7TQZwi930pj28SkDf/D
qY2qva7PLZf7AjCHcLfSZCyX/QfW4l/aaQLeAEDiTeIJB1QWlF9aAhpDoZRUv9XjL5GVvLkTt0PI
TjcyDeDnpSOF1EbE+3rBy7esE/z7/MUAgTieAyMruhcEycq0DyAXn/A29DeZqwCiabGmpe3oQxBk
JU8XhR6hI9saruOPni3G+MFzIK23JZTZN0zmIYytCJfvEjr4cjHS/ZlXe4cJ0ffKToJRAqqq2n1W
CaB6GiTfkyvkKUnHBGVhRf2P/ICYrQc7cShPZwjtwEHy/7pEeeW+uouSGQBbKZyOP/ulOGS1E/E5
DMOJ/3+Y+wXesznU/FJYd4xBID89k/UtoLIrlY1PCZsWZGqB8mgjBvS1hHsJf9YnJ06BXcRLdDGX
P8PFV+ydCENYLSr2w7nBFocqYuI4GukkGEnD4d3A/ZbHMsa5wIpkRrCIYFsJRRwmVmrKj50GH8z2
bIRWiClkHHzhddni348fTfNHnnWrkF5jJzezIKgShBr/8dWMwm/RwpUW9+ls4wc++rrQ4os0B9i1
6Bgm1HkpiurVW2S0367uo59a/hsurQXLyQs1l4HbPFh4iHmscUAgmUNrANgQqD+4ZSfX6gpWEdeq
pTwC0WSa/BAqBzQ5WCaVDiovxUuDyw2Wm0BkRqRbK5zfzYZjZHnYsJ+DkX/iudJln/YvF4PgVsFm
nNU2qigzQERayJ4c71BGs0XcSnhvhMN03nfgj8b+jl18PiTRVkLeRIHePfGSyIZiKFlhF6t9fjQG
KGI0DcHjtU0AZ3gZ4kg413nvLA5gQO2ztHP+usuwCIKZSyYgOTc7fAb+pRN9ZCTF2xsE2eB3Wjtm
FIF5dCo6NVEvN02LIO7zHbqoVi04QsDcVEuF9HfzGsF9eb5k1YRp4Rq9kQahJH2wkHvw2VaBKRwo
/igbbUNA40/L2cbZQb/gGgMggUeqltDXndAQB4MSsqo+RXYzewdKayjemBye+nLcdmcsdIANV9WV
IpFyJ+2fckA6GF66ZtLLSK3wUrH/2jEkk8vc1A0gVbuVh/umTg0FK9AMKkx3a8Lk+PLWZEL9oCSd
xydOCgOl3E6k08JByBuSNd5GS4vzNaHtMrBEyt12sAVlPSWRedxBRP9cJk/hdY6YTdEokMcMGY8a
YpM78SvA1BQ37x2KNsOhO2YdnW3sf4JvZTOBqvWLkEZcnYILBxeC3jx9/P9GUBxRM/BO2orhxbgk
MPzD/Xm0oGEnburZQ9EspLTz2xYXFGNRNeMur4WlLAbR3d8nMFEU5HgDhjhnUbOZx5X+5wllIlT7
4mgbayxnBjht8k4i5hjXSSsvKRjgI7mbIEHpVEY+S/6P2bKACnpr6CzE7oIWRoeoLjGTBfkoG3m/
qfL2flBtjqclK/i49IlZ+ZogocXNUVl1FBFMTrKL49GaGI3GvlQJ15jzl1C99tRwlkqPpyR/uW9I
zkDhtwQsDolwyHOPDJrCqA0KJHJ3IfAFIjLwa/MFaTlW8lDJOF2e4VJUsFe/Oknxtyv3onC7Epfr
o1LSna4//3YDVhvk3QghNTaruBz8XJxy96jbCmtfhGt1Hw==
`pragma protect end_protected
