// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ppwZ5cWIcuqRvAE3G9VnqUXXIFlFbZs+yvMGQgHik+ZKtNWgfSMITiG5brPKbl92
5NQrVzPguUi0ydRJ1Mk57XhV5wU6xe2orOHrJDMcTbJj8aetY5exsH21mYC6otOQ
lFsWtq4V63VpfS096OPHoHj8xWMnouCCCuetZJ750LI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3200)
FWZjSdQiUd/8nQEMLDPpICDV8cnpXdmDFWh9qPKCqRhCWD8yWgUp40RGIkcOy67C
EtdhQ1O1vc/aJny9ZuDb0c5Aa1xdf6ZZTusJPhn8gE9gFck/4hLpy5doVbyKR9+4
D38X2NfACvC2TLBhAibyMKGY4dta67jxsVwGt8JPIB4Y32B1b/M4DhYwlzgdrQkJ
wBbJJrsaJNctXHI7PZcRNgMTdTmILbLu2TsD4QSEqR8D9b86FOJqihfl02kQrEZt
NmXitn2HsT5wMvU7LTKeZidWWyH6je1kXIDLmnLVUoeMYOkuiNtqlbpv/x3L2Fdd
FlIdi+Z68qtSykRgdYenW8iMJ8CAfBIGlGYh53QaZFkLAGV4voHC69uJuvbclnY2
UZGJHHoBTMGojy5XSBfOyg6CnCa0Fhhyqqqq5WSHYh7mauS0lowBAHiQ5L9Wx0v6
W7KHrz9PEGJATs/Iwg0Z5Q+TT+XJu4IJfKWxuIfDbZZ5NsAoDpnN33Kg5ymikKyf
hTNGocVXHrhfFAu1EDogbeRDpAMn34m7zdfxiDB6+6JcbDPCrJ6k6kdhm6MrRMEX
gAG4yxTc+q7S3TGdMv/UH0YPalGdbLKl3FsL8CUQELxCy/wgaFH+Eu06MTr0hJcf
r5hUORPKs42zGD1HtRoSVzBM5MpW3V/BT+7+ZF83YV/eqQFsiYknPvOgNO1Z+pXG
MvB/BNxCsGMSNMiEL4xFvlfhfBX5CPAftZyjXGykAWl048HSC9l72MLN4bh1Ralg
tVcy0vvUOHhpeYIDzn5Uhq6cyRNs8TrALuvCEe4eTKb5coM3CB8dB+U8lU2R54D/
HTysS94AU1/lbjgQWxwYhbUS36HYBwg68nWZ8ju1iuvia832+fbB02NqJVVQqMIX
sfQNU8+0KO5HTXniC/D3vprjkEUaxa06nOBirLl7/MckVVylPeK7usTorCYINeSH
Q+v/GUdggRpkwzCV3cuYpEylkWHB5NTP6R2pQJ6wWl3VLv+k2nUDCxwC1eTmzuoH
v4tNkvQMwAI2ZZAX01svFK4BXgm7zBNpgn7LU3blzqPqpSU4EH45aX5KmyUVIbLx
RahKYff8rJBO38u9PEr2ZIw+IzttJnKTJnEY4BkrRmJxLEVc/ZO2/aC1CtDVwgTF
lh+X90+WDMdQ/YDyjeCJA9KoWR9+j69Qr4iKifoiL+jrQPV6zW3FTz9kXawvIeAP
zxM97ywZDa0glEHwVpdn5ytPiKu3a0bGwcaVSYCjEX4j79OoCOjuzPwmEqCfd7Oe
ST2pzNMBMS/HW3GZDHnlr4G9xD8CKarYB89MPpFzoeXYGqUDIHo7wNNfBKamTFga
kFZLsZcEOLf8sVs/d+B+/KGsuR4QnMlgcC160SXYR0f9r5/7RTapMOIphAfDja7z
QIiS2gsQ53ZmghhSA+m+p1HzgM4KlJP5icD/f2leRw+6M+HNPIag+zqmbVn+vPRO
cNqMp5xiO1BkFtq2Q0rBmLctM6pYXGcDFJf9QV1YFpD8Sv2LPXLK4j2dHc4zYpdQ
yxYAUjKm3Uw1UptoNJvCaz5dCUj2DZLqquLiw/tOrIFTQ6ytRmXmPosCXg+kBEC3
8pylrFuArzsgAoROdK/aJb+t7eU4VqD8OqUtqjq06qD3+iV7KxXNWh2J/KfnNEpv
GMxbxhYyQDGTxCBIdHFinxBR7hNHGOf9xl5BSboX76lVPUurROxtXKhw5uJSwvdH
hqASUNElG47xO2PZznC1mJDmpiYG9DQXKi9P7TraODamPXSHjvvU7wEoTOi8E0um
r0vYq48b7sTfk1FxLOpKYHn2mA4bqlzRsccfCpS076+aLLlVdtpZ7EpslmLeNd6S
meExbmJqN/q0qlJYk06Yo5briSxVTgqaMRD8sdiAk3SWuXBR+tFCq9pIE7k49H4o
P3zoU/RKvVKV1+iCmvf4Qx5fsXf6HatDTDwgarKnCJ/7xKtmvSHE37IPBhaa7zVV
P/1+nxlzOlaHUjGR7saMZVYyFTy6zy4blisZGcF+J4J/TQcn45NoBjXXAYrdEtO+
ae38FFJ8W9+Et/QpxQB+L9RYtmYVO1H8tzZy4MzboGzrGIuaG7Wu86k2QtH5/MWi
Jm5My6OT+s27AV7fgmHv6BxqTQCjaTWvB1sccGOUvDFgfy8QKvtF4Xl5Sr/ommRe
sC9rl2Ad5aniVHIvALpyuilHIg2am7BGZgAdhCEy7sMZ8eY9TAEVyNPlLq/7lL7t
8id6jPFMIjiWpn0dH71LR6eCcXSpENumXA5ESPGFjwok1wV+hngG/+RLl7NtnRS9
dbSA6ISpN2GGXy28osAJkD6pvrmt5BWnQpOmSDCi/HOSyl+G+vCpL5uaXh//3Udi
8PC+rDh3pnszgAcizGZbfX98w64e2/G60fmlY6AHptS8gG3PW4pcL5n2RIZdLrY1
mmc6/o2DNJqTHbv7nNS1JMrNBJx+RLyhiKaaSacAOtV/F4cJnFxxmAdrGYiy6Eho
wsZ8jF0OQKkG/6TXqo2y/aK/aIPvFR7yt+RX9SzlvSjqhqnL13LDtz7ouKSl5t1j
oX25Kp9lfaILXFIngRwzClKXnZr7z+PrqpzAlajORAeUEP3+j0R4V1a+ptpUs7Um
+2X1L4380YGy4GXuMr7KGTx6CUn6AcGWr6K5Njm3OGEPGxJOGAM6NvqXYxzAT3Ku
ksQDzMLKCtwu/uK/aEtDuesKLK8QDYxl1omto7ozo4/DPBIn6GFIhaqGshqN+5N0
MxQ3kOozhzgvVuASaX816Ubgf6DmToQjhQCtEZ1b+8vj0CqPbpvWaITf122+/IZn
x/zac6vd7gq5NMNj9HCJBPJtxZAqvqYmwewV0zuIhcUsEd2wMvOpTUw8vGaEJtop
m53sV0saKOQ40cUOiZvGt+eEL1P7tmUijo7F+ETiuZg6UUxu8kjU5qZ4iES03G2y
D32lCoanGebWFl79qc5Fi9Ahj2u2PxClgUgeOzjhzBCNbaEvGq6yZcGncGz/RdAN
B55e5xdA6BxPXbonfqYTEIrRvCZ5YbcSLLrU5aTEnnIa6fxIgALPv45GRb2kSzMy
igDniQXdGvKw5UAUpWgEgl4WpkUS+OWMdl87ZbHvzfT5YM7gJoH2A917zVXoC2vS
atrYnfOl0QiszAF4ZxTBF4Gp2y9UPmHFulWRLLGEnZe11eik8QCLNjr3jSVUGAbs
ostjCD1zFwYitRhPxBYWwdtbikKivsgbRpXRt2XEAQd0LdGbcF8buKz4shTcSAmZ
Wo9ppohpb4wTUNMyApohOhFSBjsnFEKSQZQw1Uwh4xCE+Q5wulD6e9yrwToqyKSG
OowqqXGVEnTnd1ePm1dsFdnB6wn4VI2DYUJAIpTCsy+7UYr6vGrw6rej4SP1tktQ
abBmVDMMTnvkqv0/i8yy6CyAhIFTf+2KsRZUI6rKSHCEfRd3DslskbUaHlqT2IDO
lvFHTJjXUXQ62v9s+6T/5Wfb9ea+rjoTky3W/YcGlalEauJvr1DIcpkAVp66icY2
nMKe6+1+wPdO7Nn2PmbrerYaLtcMaL2tyMjtJpQvMqFbxuoAj6Ic2+6wgGnj80/5
4BhzBS/8AKBoFeZt+MCbD29qE87ACb/mD5baeyak7T9rvXhLxjOj+ca9QFAsKnra
vhdmRLkp3HXuPN9h7YNtUDptUw9D25DX+9gHpWSaR5Ki1NQhdC7Ae7bPHNYGIRBt
15zXvYNtYMDXL22va4BpEHDXbh9MYhKRvQcOGacU/wYm2B/pNrVtTP2couv+kAsm
UF67cnYveZnLlA74DFHKt9+pXmQLISLR/EfPO/i/N8JcH7MV/zWCnUF+eFqVYmir
r0UOvoel/OkFnSVLUE+5/AywsDWw3oF1dQM2wqLpOZjzUgiambye/GonBGuFuyw5
vAxFLf5gZQboTuv8hlFJPu33gyNLnatcbFQmhdgf8C562YeQzzNAkDO7AgH/xi1N
E1NTn2o8KxVn5Ub6tufw4EF9/eXj36dLhKa6WMwb5sh9Cez9nZwFTeScn715hO0y
D3z+i5Xe8/4DcH8lvoQ7e2arFeuWMghj7jp7Lvlpc7mNMF+/hrvP/5F/T0BB3mlL
QfF480mLHPLgCsRYYsJW+O0fJVqLNjX/UUcvTKe+Llr4LH0fpSlBS21XjIXTv5I7
hxMDCISJQzzzNBwCGamDszcvA5DbAFAn2qA0U1Y2ff72qIdCIbl1824BBPj9k71K
iYfP1PY3rGnGCEmNpRyuX/4VfV4i2A6P/cMluzIwv30=
`pragma protect end_protected
