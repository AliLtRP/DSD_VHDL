// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
NKcauN6q8rZR/mzVxW23FuyPMSbOjYhieWDbQz2BzZhXh0c4WwTcDSKOzh7f8kbAf9XLJ1754CDg
xwUMlO+iYF8jFWqcfUdTrruu9ywxIzROL/L+xAFDrzSck1Kf3N5FKCOqrES4dL4y4awH/CkQiG1n
Q9J7pFYh/7C+RUiFdjDNCiFQo3njqVsOsRamZzUvXBPiyjvF7K8lYoG7tg50rU6BUoIz7oaHaBwi
dh8X/xJYLIyMxqc4zIfIOzr5bZ45cMWpZ82ICFlh4aMO9AscZfTuf/EfhO1SzDKbAv/1tzr0JeJX
mhOPTywi5StNWTeEdNWR7v7eeU5Xqgjz/65tVw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
N5uEjhQFS3zWGx7R2SXu9VSXR7QUY8k1Qx2k7MsFHLcT+dnGnNPg/MUUd8Nw0uwCW+iGQpImM1Um
mYffhy+j7b+J4Un7wLsF/2kYOQa46cSTGxLld/Qy0Y+2R17f0QJTT5cmZ9R9TVINCZHgK3Ahyp7f
cK7Cdi85n+7IaXl6W6ObulzumJKrVS+kEefzc021mh3wJHu5m0jODyttJRKdqvuVARRVwdptZeN9
3ebmEZLQI0ktp7ZgJkMbje2e/ypKtzVzdzRuNc6H0HhFmNNMIsdmbaNFI4/DLSJVPGo9vMEi5iv0
uZPP2qVoTjQLwZWeOevTX6cWARpHHDPdteuqxl4GYb4FsBhzuccN3UlYtfepo2gz2iz21xwh716v
wSiFrU5R9eLy44Z4Xj9IQsznhWoO2KSScBZXeA55MbyaR9w7vLjZV3re5R6sfFegQFwpMCiJtQcQ
AHNPoyNcBQzsrJfjOMFn7V46d+tnKWjAUBnJEEIA7kh3cCINs3HXGzUsLIuFNflSB9JOGVYdMf0j
84iisjl4o5XpWcDJA99srKeWR0aPWCEpmPJiFIYgxPhbPJzQ4AXFtacUbb17nhcCVPXjTqFQFFhi
aC1mp1IQ97jSqyS+nXIbbZrsDx8qYqyIlIzTpCeKjF+QSUruanyxaucVBscKhASH6O//eQF7P8l8
iJ/ZiM2dxljkcnueFZpO2MsOxBOrb7cSm2xKipQosQIYe6Q3LZop3QxbWzijq/0XBu1wJEkD+xqR
q1mRSQWegGdLpnlpLiaiUM/cbreWvuPTi7e54JMZYhXrByfkSzTy1BCm4KTZOTlpPN48W2IMzPOj
Gj8oi9WWqJbLPJ0rrJVS7AfRyxBGQgpbXsDOtoAjsitFXJYuk1FlZjQYi7e4ISixgfQeh8+8Vx1h
RVPLfuJngQaVcrQHLf9dRh1xYvaBDFtH1MshhgroGVdSYqqXzAUMtV8Mcc8RwfNAAcHwbe7Of4xb
TPOHbfwXUK1zvplm2tKSigAU1KlLQC9IWe7MVJ2VCz4Q1CZlYMdR+xK7UmlfTUK8ETfSetn9ktnf
6f017pFZA/H+at4RyNDEyPJUuj+WTQu3YTdTDTl5BDlaOR+nPVjqCcflPJMViF+3kSlU7sXQPxGa
0k22RnS2AzxbsFNLS//0aUV3t9Ge9yzttXrGBSLP2pFU2NybifNj1ZRd6yj0Wul3ttnMMR7frJr2
zF1hNhbXxCHnEBZt+CoD4GpCp+oRtTN1FbcNDw6vqYJC5c6fBvo/5XpMIl+R3Bjz+Gmn8otNBhZn
0v4uTqPldUY2EvYfFOpKm/lyLM70xuMXkPMHaEXP0VOQPXTGoRw/CJYQiC0ILzSQ5tDMBX9m1byr
n9Ghl/Fet0qBwH0sZcr9OLWI/tMyJLabKaz5I7fme+hIbElivbB9nd/ystrCOxbUwVcYPmOu26lZ
3IcSxWw/fjeNHSCiAN0SDDxpcYplaWyXz2NeVl/YPw0QcruWg4ToQSs4PZYPBuc9FlQ4oawxAp8O
E8uowbXhfcz/SuGG830DnPMs65wIM9CnuDk3jNByMRRG1i3Hrs7mOomvuuWduiTUbZzuFb/XGW95
WD373efWsViapKwP34D90romV6jdGQzZ7HOoVMsB0b5F+MzalrA4VNQ/YnQ+lyVDpp9XflJV4+fK
yhX6Jq82RZiPaJdpPz+PSaG8B3cvWMdoDddmIF8CJZVbWP0wIg6vgDBGXOuRVpbazjuQ9E9f4/mu
p6oG5/l98wPE7biv8VIHi/Y28Uq9ut/e5QcfDWpBYrFOIkowzp8tS5AkdBKvKAVD22YlkVjuFF2x
dncd0R9nZmTqZF8oaV2QJqqPm1Tj+jgIoE59y8VfLulIwtMm8S2CfLro6/RbVIh0TS9uvzjRhdIH
fWpe7gWpZukTXzVBQaGIwjSg5fImyhZSu6SRsoNi37wI/L1nN6KDKRf1ra/o4RiJokhStFBO7k3L
Fc+pXTfQiZDbHeL1huR6g8a1h1hFGcFPJUPjo3S0DIw9qZ3Zc5mrmF9GHlteco3IEU1v4xfI8ruC
VJZJHQmzJzHiVsjaxrlD5UdJEHJW3SwnBgGkh/TKigOO5kxnCgd1gGjMwe9UPtofjfOU3+8dqCXo
zcO84/y9GTEIs8AycisP8YiiTNVhR4+Pw1lbh8HZHo7zGffFxUQ/51OvdE4x20U++ZvaXKHMrnJU
u+ZzWbUtI/1etSNXFzG+rwi5c3Hb9kQx+u+TK5eS3gTsKgtLm6FGVAbVSPx8I2LmvZ0J58MQZUu6
xDjalD0K3fAY7N8A6EcvscQ1cbRQfDiyvm+jdDaRl5Gmje3PLUJajH3byiT2SuhMTOQ3OyfU2hSb
ThlHMeI+FZ1c6OEuhYku4zINYdQ1SbyJFksaBEp+gUl9YnFT//iivsd24lAu5ubQXJYQJfNsvmi6
zShPmezy5EBIUkW/kCB4BthFXVJbcmvk05ac/fsGi3KhLLU3+2oRzf7NizffrgmO1MOCcV9Gw27s
4KBVNidQJvoXlPZI8I2yJ7FBLOL/JQEPdBxTHiJDdPiEp3JhgkpmAGTWC/1Rin7SQvq06LrMiSUp
xtFRUyrlrHU130PWuPoe2crcyudDowoNtvl59BOJdpPADQOMiqU37Fi/eTpLZ9kSP1vyVV4oyy7Z
X9gRpD45ivkEL7rmRcP6J6DQsuLNTtMmqH1h7TQsAAxQyajGGQ+n/UaReFIP5Hi/wpa3LnBoxoqC
ctk6GiWEZfGqRAZbXZHuJ8mRHyQlQTXPXF7nfOSRHrKZyXwtXhSmhZpLXyFep399IWrbYuGP3M/X
V77PBBVwuiQTogfBswvollq7287co20p/TsWbFVDwvWktJ7jQY9N9RX0JD6ThHFkm888vkqQc7Z0
/Cr43x0GLVr30wf2eEMkpnv0nxVZ3xCEAhLbl3AYxNR7e/zCw1hVmjB8cyuMrTvaYzslq+o2Cb07
hXGQqcQUhmsBH059mLrNoAOH+buW57pIG8zWKLv0DMtY9u/nxC0DgUtJ658Oz+fow7EO890FSlcb
4byXEcMWNSkxmslyiMJcV8Pb24m/YZzerR2Lxif3TG8h0qnidzLJgxS66BmR1DykVzpUBKVdgWp0
wKi01WBkI5/gCgbVXp5myrZyFvVognQnNI+Qen4kD9B48+n+8o97vAfZeg9qeDBSYmpQbtIPJhyd
ql873EbW04jq5MI+MCKhgKG46bnMygBnB1ETtqWPWDckiE0hEGZPNlmre1iTZcpUOojUjZBPEqRm
wgSEhc6zdwvO+nP+C51Zfdk6nPj1jvM98wqafKMU5yB6vI19BhvIa16yIuFX7W1NFAeHZauP+A0w
/2n/aXL/ScPJ7Gtc6qnBfLn+2ZxyQSOPFxFVkSOGGWYZsL9XJKk4s9qBULDTBNYVDuJ8Sq67iczY
bQGG/P00T4Xw8zzAJji2/sdBho7SEJa10XFI8i8QKOAUyR4GJ7oVzFgefqsUPzZndh6SbWghJlyj
uwrIOP5L6Zso2R0FtXA5uR4F9YppaTAtkyl7D/s5+igaLfQKbNDeIW42tVdDPJKD4QcJuS85F9ul
Gt6z2BsPW6wko8+yvhVr104Q8q0Afco/olkoFlOPVJMCF620MeBTN3CiYPuN0iN5jvOlY6k4A7Q/
tHojtG/B0KsmXh/atqoGbjPbulCgDMv0SBDPkGrm8d5313/Brm5ruE+9hHsoxDr+e+du6JgcBkaj
wGY3cxqCJCx0M6PMmGpeAs8yZaAUk9Bt3TcW7hLT3tbaIFr85QTrFmztwf/OpKkh9tV79lIf+7aC
oVX8n3hFg+CyOPT5m8+n4oGY2dDfs5uwujn6iYzqA8dtMHCgmHnym1r0N2YpLqFziOExLPUPr+NC
CK4n1dVu7Li55lWNAnLaLsltisSVaUPg4ANs5U7csBv4993x7OOe7zGo5BOM97eJ92iedpNICPcO
6mdQ6lsEmu2CSmWhXgV4dvnjibNf5aNnIXbd+8xuFaoWlR8surULL1oV7SydqOKR68gcetY1SaHp
Kku2Q6dnMO8TP0zmmcSwTApb3qZRUg4+KINWrHRysIZRKNDzg05tCrzeY+u73LCCI+9Fi/VVTsEi
HdusCrvjOxTmMcN2vePwNMUCtPEIHCmKHfX1n1STj40aSWDTv5dyDcWI/uQoFrZXsGncWzqV+XOe
RY/jF0vPDnfevQMRh19ypr9w8pMTJEOKkf8RwpfOIa7uygRhC4hBPz5+S0eC/HEjQNB7h8wdsXnl
gvjQgsuoyX1gMcQGieKKuH6lYXggHYTJGDjqbeXovT4i6+KLzGn7xhC1C8ThcV87nEPyxRVoOHFZ
6lsOFYZUfgCGN1pltQsqROEs4cUM9I76gA/Dy9rjLSbgtNFhLaTr8ai0eUYJR4eKlBQrdUnjMD6I
Bj//Uni+3wzuo8gDdZpq3nE23+IzuYwS2sx2lZC2AiWo2+Kvn+ezE+0oUNkogbEkfRyf9RuqPi4P
RxXqZ/5gj7EDNmue5XnZ6vaqedZ7bbEG0Rhq2DBOyUwhdW9/WBbfmwyr/aUZqufDRX8WPSLwa1O+
7kgcD8BWAaXq+1yebs2Wx4wLgbeOOTUEhMnd+zLib+DttARf6bi8OCcLzezRNsMNN9lP5Pr0nDyu
xrm6+wb9yKqSjyZa7tdcUfvNKwQz0V+9kZhgwmJTFS3sNqUBx0AB2J+DCWpUCbP+9zA9cqKb8Xvw
9Y1C3uK1VWxIc6XEvp/hxZWaGxdZzeBhypOyMD6fr4rxdEN1sFcHDu/ReRUhUBCKIOJXzCkux17r
XAhKo8jeBH/rhWaucK7LfKzou/0C7aG+rAcr6jrUShz0hT6/tIpb4E67xuVGh+xMCRnspx6wMytW
eVCvIBRi5CAAWYueOGY10e+vr8QL1BcftE82aGxiMt6vWvbq0NhcjcTQckkyRC26yLRrbQhJWc7X
H/sFqtpTJirtkAcg3uzu1Dxb2PCmG4Xct3nNn0K33TNwIKcfEXClUwf5oGBJQmmjW9Dm+Fzwvyuw
is8cGTgiskRXuW73PH777xfzhyrmLtrKzD5LiGwFD3mUqbNdi1vhtGbowbanjui/oF1XtDZZoPyc
f6r6fBzTihEJdN34PC0fRY33jOAAhs4DUxt7P2BO8br7VJN6r14Hzj/g96x+bPrSBaES8jne0Yq4
4DQUx5x04Tea6YWFYXlovzvl+TecKOS8JiHPUoGTgwnG+HnLswauCwt6tBoayjCE/AIREV2TYiBi
kFMjZtpAU8OL/Cnq+vrEKscS72PmxqmWFrUmE3/TmwBk25oi+MKREXSpFBJsE9f1FyhVHpXr5M3J
mvdu9gIjCnXO2Lv1iyJPbfqquiQH682MT5wvF3aBXSlxo8RT0b6Y5EehKGw2Z7sA2Akcs61YslzS
Ubn6tQB/pDdoY8EeP77swVDrbGPLY6pUPrNPeg7fdk+suSvKs0mMm0AXM2Cxkz37bxm0YejDQDB0
iYOMT8bO4MzDspTRgIHRRR1inuFzoGwRCsicDN6XaDf8blJnMFkPzgHCACGAZWcR5xUa77zh4bC9
lXW5DZPbBa3oX9pEyZ74yb1VjwYFDu2J8B4PywmMEOpzE0zBPJtPXqMIgqX6laSjzgbsLswK9Lom
HGiu79tD+xTWEhzRmQph/+EexrDPTXqd1HOZfJ72hMgHnwq+C0W1RaEdbHfqwmvcHa5K7P049gPQ
qtuLRPuQkGG4GFt3LQGu8KKymOFkMCs4y2ylulugNhDKj3Nf+Gn2bfbuwy/2HrO3ImS2LGrKHRiw
pweuta0P6M2RuM4SppGdt94sj2tgW3ehcqsACe34iHFn2mNJzJhORl7zZXaAiLgZJ9tjtzRJqZ/I
12Q6JeRKCywDpnfqciGQvLov3Lb18zpdXbWaXCgWUzKQVizw+ut6MZBNnq+FWRERMfJd1wG8Esch
W2+EaQFESwgWv5yyLG7EbIxFDTSprGd68I8bhInH/taNatGGNXOvCSPJJH1Nvv/qEyvhbxlq/Jol
Yep/UfZPssboiW9rvjgOqp3l15lLViKnMLWdP7GjN/TPC8MDnGfNbevACwr8Ik5Gb7YA1V5JG3xq
uKn6kX5cdLgeNghciznNLFqy+CQmQG6obRyNd7sidQarF+d8ri1kwQE1zClkTZpKOGxj8IknsnPJ
AuHgGdx0Apis5kbK6quLW4hfX3evXQKwEO9phmY1ToPTEOXvqbRLYUEvEuD/mAJ8PpZSTSzSaiQI
oaOppvuk0YuqpE6bCulFmLGOWkINODipdUVAy5Nr5H0ZOVFEL3tVLL+daT8XUDnNg3lnmuyXqHJZ
/qYOAIqLk5gwiwhvGQI4TNwA3yTlIWYsqYNqE/P5dS8skxX9M3i9X2ZK3H/Zw+lQE/i147GrT2E6
NlAWUjTNEpMk24lQpibdaBE4cjmT4ohYqw3jJ6jObWCuL/ha9EJGXjHLzGVHg6eN07N+r7kDPD3R
yKzmaEEr1whmZjNg3tA3GUGY3tfn8BBemncrjJBz4t9bDWxK4pXkuJ9IxFuRqzwkLY5w07N8ELwL
tvfSycRx5XmjTDqfb4/F2jQJ94aKTJjduAL+Iex3m7NoLVOXbZ+qq+hqI3fShspOLDRoNsJ65Mp8
Ht0yjxiJ695+8AooBELHlGWqMzCns4XLeVWBOMXKRxg8WfzQr6TL1k7YDFl4iM38VF4N50qFxp39
Jl2MqTC6Bugrmg6bFXl52OBN3f7vFdI+XAejAk6Aq40A9CVI+PNSAkukEYzILouEen41I5/Lro/U
6DnXwMILlnRXE4Z/IcLcsms3dJty3VL6WRGyNPeGrZc5Jrn+6wMqPH2ZynIRoWIdwlbCqbCZ9QFc
HvHIIh8ZDTSO0oqg2gLcjesZ/n3uMfXIk94psPTZXQEPRgYB384QRivW63Kp3RJ/1yWqgdqlH5so
UOM08ZJF+Ta+K9kGGbxCXNJdFxtHP47uFbH4RoRlza4MpDTK9SpU7wXGOT5MFt7JS1V5dIpy96V7
9bEO5z4O8E52K/rZ49HFpr4eAprEjotkgzNbcz8nXoMpeBAI4WcEcStDMbJQOhR2dwlnQE2NF4sR
mk8DJy667FowxCc+BTgsMuSmftxsKUq+QB6iqhA3Qdabuw4cfx7RX7X9KiPl+fDJqGgynV/t1Ncm
W3UOPYOiTADuQltmsTQdGWtMGPpBamuVQDn3SATH/vEc50InxtLvxwU27V42E+UadqiUgkasp65w
Y2zB1wO7HGBt1XdJe1S3RX4lVWBeERCEs4pWmRCsocUkY1iRwCDQyCTAAC4M9S4ylaLcWE4IAqWJ
a+MiazZAdq/dJt+9ZPtS0OElJmUnEtm/uW39gZOs8iTmnf2oKylIfLBPJrh5w5aJm0AD18XfAX6j
GpDOO3Le2jzP/W2olj1Nj5idFAOX8TEEuCeP89gUTYQ07Re8q4pb5gipsJFsEh3ApG75apOYaS9+
CR5nB3Pm5/mcZsO0a0uDCMCtHoUeNuh6wmyzij3mUfBgr9lZ2EMShV5n2f+iVaZafu43NU/vE682
uCUtymrriGwPzbGAUmkxxGelAr0LapMcw8NiL1LhxxBzuHJrul9e4/UqCogEw+W3Jk73KgNbS2qL
uQ0JMmEKeoLKa87pG2SHwbS45m+oxar+Ps88Qlej1R4mb+JJlX3mSoYxqRUkh7WOwnYlY2i7ZZGn
207uY46sKVlgDehlFgNzdU+LvWJC22clfQ4DMGp+IUkWmoWSmOzm4ZFJPKPQEep6FhORI2tChBXl
tWWlvpXXzUseZwZJsKjMUaTViywxW3Y+k2KFk/kgLnmb0+iGvqIJ2Edk+7NDHb+4RPAhlwYVhs8G
aiSQAKtBLad5/EAQKUxIUU6DeC7oHqmmN32q2It/qLLqf1y7SPC1pXTPo/PJZbDn/PyOZ5AHTLMD
9ZynGY5RW9pkn9Vk+QoD5xrx2hK4BloYOIy1tRAVcKoZacThgn3w41mo1kK+dSePiXMmYrB/Vk7x
A0nC2I9yScwqj/X66bTYNsv2fNqDMxKu6976OtsC/fGXrMUj6H+SiTStUgTfb6+Iep/yzmlm0q+3
m61mpnY9B7HsyL51oLuurI+NKPZRRUjbWRBDRySvR4TTguO9S6fUk1GRVfztrjqJAnocwqQ4igSB
HCi//1Pfe+ekJoEswEjgSJ08l5E4QA3wALI+507wIaYvnaHDfaTxSLRsW8ysXIqwTpV+cNuz3aHi
wMEw0gJfKZvt1ECBuBuS5JL5aUJFeMzxWCvejQ+rpCUXupPrlK8PtOYO2/VPXUlCWKCcRpWWkUNi
UmFwiKJ0PJ94hBzA0KdJyD5dUN6UI44PDgb7Q8kAMY6bQEaawN/WCWU1VhhrtL/UH12a0hdFCEsZ
1Q3Cuksx1a8x7XHTSWQt9lxTCGCas3ickW7zJYW8Eifh1AcxfkOX3BeuS87piNWQM6WhrIDhIMqG
rXigwwtwI0s8V00MS5ZgOnJCk3kNjUfWp3ztg+DbGhXoksUppbPeIgtWnnRSDa5F2YK6RiKELO7l
kGFP4zlIc7STVzAM2jQcZeMw/2FsrrjuTpmrydQYeZ0QWr2QdB950w9zdhbQTYH71/B7rJZiDxCe
9Sq9sBhDz/5LSioRjnaemcGpis8eenI3HszQ+JduyFIy0zbriieyoALHXwfXrO2GnKRYXtJrFF1n
8ZJJ8l9vQNI0HpPddnp0yDPIq59qqCfwzXh6RpHVYPY9/+dwPLfE94KCvOY2wcA09sr6/Odc2jFM
ZlrmyTiHvKe8haZI6Uq77m3F3IDBvWZWsSaeg61uAbnzK50U+wcG7fzxS5jbaqkia/3eYzwSmTdU
6d90HChUKvZ9AwSn5jM/9MhDWVfeXqGYVpjbXeuwtbVjA5j3K5Fn/w8lz4P7G/DedDyj8ZDkQ9Xg
RjzdswzSGBtKMOe8WOfaIKyMEmR89sTQnRDf5hmCXZ4pgBbl4yLm24bHW79mqNB6LFDshl2AZv3e
szJ+tcuhPekijrBngZx0oyJohCmT2cgFpjvnkLQTAk46GfHNGfbJdpqTfMAg+DDSrkFmuLCLr9k8
oMlCMlzHs67u3GsQp/4uEb1J7jZBnC2exdnvDutgd7xark4a6MAglt2FbRElFc4aHy0+cI4Tcr4U
GfKNuSGhp+5C2r1dmg3edfoSBBhtH4carWS8QVnLbOQUsQrj/S6+ccVeVG764Ke7xP0ful72XJ6g
kmaFaLrR3LmBc9XiIbiHHTDIsiTX47DTF0JBdiwOooR9tRqz94eJrrr4J0DTaT7VRiIuzzzzomk2
6C15rkVPwBoxuzAqdLmAKGiBCcPXpJ/kq02NppE4U5JU3uRXu0aY/LuGIhkJTEvSPWm4Cl2wVHm6
fVPQTJKsh8VIH+ueJAfOWVn1UDhy99zII+nADkQNGozKv+pLGNqr4/BuFNxY
`pragma protect end_protected
