// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Hh7lLBbRVFzJUFdEWvURipoMThMl+tsb7KTIw7JQTL8f1W28v3JGybvTM+fgGP7B
p4d/FniJoDEWzymnO9TiHfCyk5Z6H5IlIK59pfo13oqWaD06GVLqG1wFqslwN5Q4
AzkenPCu7Fw1Fp3J7Ux2a8UY31npE2gS6E0gTPzJZwk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2240)
d1a90GI5c4BVHbGvKqNYauC/9+sxGxvIooLEGL7Zipp4VE0Bu6GY91bZjdaAL7Ox
Hxj3alGv7lO8wlII5t7Niqdcut7oMqRJvTSUcZvFbkxVE7/FyAcSir+GWRJOeIO/
bCfRQsAyusD7zsjoiR0rXVlQZcsukNVlyhQDX9SnTzyFNdSbWP5gyTLF6GIQRGfz
/ra3W2ilx3tw6ZQBPEatm/JvFyXjbhS4kcgv/YdZU/OqipM5ssGGJFfle3wCACFv
cJjb8fptmrmzwKWkwXRQJdzpIdC/qW2gH2+YyFENKSerBy4660cwVRTR4frbL8Aq
CRS7J9V2iIIPe/S6fqqwQ3IP3+sWZwIPhLMv8BGQqOUxE7DDIqmX/iccksfWtky8
26DsWAor8HPrzPBPsidrGT0gTbQYSvZuye2hXe1UWCvmcz7HKMENT5hIGYrEkjtQ
0ufe7/tzdg6+IAyhpG5zXT5HwwVA4Y7+H5LFc0b3iGE1PIxMHGaztkYY54k9GGfr
8b+lU8sZzhmep3dPIIsLBj9P0JCPTQsECg3h1J/phXOXDmhrjVRYlogoLGPzajRe
dkUm1URmfDF9TJwn71w02ydI0z361gznTa5wACtm8wwbUqRF96EUwoUUDmHeh2az
t7Csz4Wf4Si4ePMhiM7TXOAK9en1wR61kFhqF2br4OqxDdNGZFEoqK8j2JwFni3C
gT2CE+KSDDf75RntKh2jvTTDX9zASMg6AA0zenLwMiRcoRO322rkrSia4IAiQhR4
q2bkqyXUr6Dy+Uih65SB1BoUhYuwcUyuAbtg1OTzTZ/mW21NV6e1wKcX+unjyH3H
Rf/rPw6LEyrtnjX4FJV77nmlApHn/aC6F6/K+Kh6yFZu2NNMT9/QgqAktSYeq48w
VaXuRGmEQTvMYhT6ISbbJMD0f5Lwo7IVdoRodcHweoWrBLMUM3nXjmBYoyMjD76I
10NlfskNlPd1Jt7ngkc/je4P1F5Shtj7+GIWEO1zyyqNb8Hww5hBRi/vrKergthU
vHsMtgqKUKJwnBmEjR9Y1un2aTYffc45+hMzHeCVxVRGbF1Ech5euFXqaWLebrNm
Zu8QhsdfQSE+PUF5+pOrXcQnEs1HEWxPxJlEgpF6g96JOF9L2QR3YURjnqikZ+Vl
iVyz2fwAIvzlXLg7EYMTmpzmMEbpK0Dp9q2i2k9RKOnUS04lWI8H3ig1Ln771tmk
CWBsL4Z7wczanXLpZXOfrUBPh2mky1Vx+zAbj485f6UYaQShJ4EFQ3Vju4wV4SGC
MQz5N19G96qsAysCyZ+7hz4bwJMRBu75cfbBEg6mqH3hCVYu+/rmxKi1SeZg6Dw9
r3PQeff4rR3hnWir5eYlgrM2m9AhFQCA9a+AoKhR0I/Dz0OIJ/tawtZOf9H+x+Sc
OefPxLDpSoWdhcsKrSIzPHgFpcO4okI3BQmd4Ymi2LW6n6mlbYArYxnKUl8Qdlv7
I0owFG7P17qtVccm8B3NI4fC02bkBzi22hO3n0uSSY8H9eE5uuD3/PiYEJbX81kh
DY3m2aFSmktgsc518lTbPMFDtz5F/dpcWb4b55v7zn+OWQ58H137xk/G1FJgKa5w
74pCuKR/EWYySRCYbyYIM/3Px136sWqVxUi+VF2MNutkFIoqfPqe4DF7htrpjPOd
HlU4SoIRRHKXG44yo+mPPX/1aTL7iSJzRc7dsCFUpLpyYn1fPK6bIlEtcf8i18Yj
AIaSvhU8t73MwL4K2hXRX3nqqRJcgt+a4PqQD/rgopq4apb2UqfPr6Lej1hLltJR
9KfW5DGPqD2W/TP1sZfgpVzjtNC9nTtgZf+z7veB5WqX6Op0k0Ss7DoyKiyIhFv0
xWOgOf9V3KFU4dPTEgFxi3NXB00N6vxdssAE+nST8FPttMcw3pibLqA8G3RxZ5Zr
SPV2/1nWFyxaEC2FJeAMkBh1ttHX+mGuzZ3oOT/4yl4TzEhD5Shu19EPO0otB/oZ
trgbBEnyTVnfg29SQBWe7nxq0k/r3A4ACT7JzJn9e0cHhsLS5MlKitQAdl/1kgEs
76EQRqMSs5JDR/UxPY/LxgNFwLKx/UV69qg8zDeCrO7mq7qZD2eaHqHyIuwaEVIH
MieCqNq8n90pIZyiSMujbQUpokU6JdIgbTYg9a3fPtPgqXJju0TVcq8QLHs7uR4H
v39C5HPdNaY+vum+/Bj2+YaLv61joQ2jDhdKsZfSHB6TWSzrJxHbLiSPKztumH4b
j7RJGO2FAzGedvuWb8QSKs8RUVTg3YlH5o4Nk8u0UE7cK/6BtepLVGNo446E+ChZ
kHKewBKDc5ND/hxLBpD02itvlLnl5AWb/7ppH0ZC6u6hMf5PMEnB9mGS7B6/5gYz
ePnQbNQBNRHBThMemtPRllZkbmQeOpo5gUzsBPmj7mi/SfBOWB9kEqUrhb4IH7pM
EbG9nRR6LanzC378fqgOzBQH4ARD8b+0Pxp6HZYVIt9REnXwOpDi1A6wgUEZ+21/
DEANHriT2aqi6Q9zAADwRxEjaVZwSRfAiAE0Qss62TgFaBxLFCdOm3o8QdOwsF44
TXT8rWRu5z43WZM0IGU2PT53j8ZedAzHpqycRX4OK9uO9ncmgXwRJvlJXUlsed5G
QxhXyAP5n/cGR83elZEgVhESq2Bex02uXuUeqkBHXXgDG7pSLG8B45P1l3fCeWXr
S3UMcYwedy4TgP27uVl6QDpkbW1C33DNNPChC6+I/TqgRJygicoC13opvq+iNXKx
BPihGWbTRaMar0gkpnvwYqJ903PSR1V6pEq5lgSP+8DwDi0Ah/PQyd21KgDIC1fD
nyUxHW5DmWk0IOLhTbWnPF/8XPE3Rt3TbTiNFdWuQ0TJA+WAeTXyJJnDYPm1QQW8
wMY+zDH736Tl4ub39Yi49NuQhGMJ695BeYg08eTOSZye+KAICJ5/MEG6Jc1x/qBH
mdou/UNXBIPwEYYSuXOMxBjbBHhWY6j+drr8elyK7jw=
`pragma protect end_protected
