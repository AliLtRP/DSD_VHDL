// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oYRUG42i0rIMzn+1lZWY4qvDOry60fHadPlrqrA0uk2gOem6zm+KsWjq6yWHORWO
GccKGiWYfHTvKtRUnD58U1ZlP4sI4aDc81Yre617+cgqI4MVBOaPzuTJpb8lDnsa
IQrEy+ByxDz/ODd2lmzoRNUTaVKXk31+SrYOlFX8fuo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7408)
IeKk2RTP1oOWnNNKaGX5qhUkUOx8KO754NBhGe5jW4CIZOBIWezdJ9VdeXj+35nQ
n7KTbqNTv5m/60Fp8386mfhoJHcoD0CadGfzxvRj+9Dr49/XrF485nXxw8glEEuQ
3+FhYg36G/algYfrL5gbjFo8I5si7Ah6qB7ivvEeAjGK3HmCUYIcwrbV256/a/AJ
DfYwg7boE+CwPjOlkseBuHHhnsgD74BQo8TFviQ4npTpi0pIDpsZLENeXODEBuAx
lwdjhiKFr6lEq8IqqssGro+SX5wFHCvaFqjDljqiCHa58eNWmrTafJAWe8FCKgOf
sQ+qwaSeviYvV7ieELTUEAJx6xbC1i2htdrque0bSWLF5LZn9EmsmwJmqb4ewjrO
JN+Ne77l4a1CXSgLgAJvudAG27r7rPKA+WRNcGcaxebfOjl9VYsSXRSvVjHayXvJ
U1/quSKjNjtyb19ehHWOOhsWVvWeZJn/xM5Gew6l7eA0czhJn2Y4pJNgn/2iKcJ3
1rRGHJ5cMPa6PPEnozLktFhExH5HIS8nSJQ+vghgrrH2xklWTAemVqO840/vdAPO
3PDBOuKH1hlZJs5NJbnY0vFHMLeMS+dUy8tpeB4eSDi1tFyDd9ImW6Rxh7kHtH1H
hi+/H6riKocM+7UrCtBbC/OIY1SeJ4nGlOf1IP+hlZ3mtR1ZCtV0WKnUevRbM7sW
9Qr0GSB0djhUT2Zpf+JgD5SFEu22lnB9TxyAK/5WTfg7v2N1DB0vkxTvno+rsVYN
U1BVN4sS5s6DLWknRU/Z0kAURfUI7dvThEVqX58+Edhcfq/mJ0b6u62SpI6x1mGT
HhWK/Agz+aj+oNfZHvJDxfUME3b0y3rm0kAHbg2YArxUoxCiY4YiN1s2v/3MSO70
MqHT0/Lmyu6bKHVzYhmpkRGR6kxQ1/oCwjqGp2oFjCUGLZeGmx226ABYlcp12N7I
a/RCKunDuaT9daWEoQyqMdx3MgS6uMF5YH2t/hlOZX514NilusZnJchV/N1KtPnB
VtiGO00ulr3GsqT2y85d5kQmh3f1zlRGFN039vfO7i04H2yJFafmjDDURDiNZzTY
Ylfxi2hkjnMOEQsx2FqX87eqzc7aVJBq9nghC9pIXrJBDPu/I1ROM0UJfH1OtvC0
EpHL/4tc6n5psnMTWuTYKSz+k13pXXeMAjCd0muZRPxITdjJ2KnfKEWsnJa9BL8J
VdTzBtlbxkZRknSznieCqFgMk2Yq9m7goFI45TBvHugr1/P+G3qDcehYzNxfoO4B
gJv7/W8US1xQWN9u57zhqwwmTjy7GsKOi8KzQs0IwSqTt4roGxVVVOZ58Qf6mTc3
rHKKjznhKMrDgbAjNjvn/XhCj0RON1hNokjJGXSUTK4Lbb1vPQBL0rCkbtRiogBN
Jm+7r3Skx0RFElABuNfE/eNDf0/VQy4rnIPg+UDQV4sy48NbBvncOuC1uMPWlCms
zuUggKRBXQpHVjaQLbq+FqTMKeB+fWSLxTYm8LRYXtU7xtujzWbgTLTybBELqGif
AwVNtn+73oRmvm/zI8cTiLV5nY7rlzIraNAStEhV/wYBhjBBAwAo1UBeGeitJ6Kk
/jKUAxACQHx1i7UAF+QF2Ki3LUazXLFSMa05faSjy3YHW8U2Zw+BhF+zdTSL/tZP
LB6mk+via5GkuVJN5eGwfCONpk343U18N/ZVVrpFM5+awI6ZME2UVr5oIMCtYnTk
7nGrBiSQDS7FDcNDMuy43AKS7S37A9dakX9QTQm+1aCa6gAMd1OGRmM1YixpgzQF
wsu+nOwdZoniaUR23s2O5gRkkJ2Ph6TXuvpQAauky2kzljVPt6lDHjuZmELG+1K0
8E3OqTerzCOfq07qfeimMnq/I5MjDEbF5BXVEgpL4hcSgTU2F81Rpc/jsBgwEjZ9
v11jRKXlrHaErA48+mAA40Z1tKB+HkKApBV0IAtXB73R9G6Dm17/BNkxFTeR6hhk
7wYrH9e9RRbDenbL6Qs9xvCizpZrByoAiJ53Q6u+ygCpZFI9aSsLfDIFjO3MOdWw
frNDNny7cmmAqJ2nhjW0TamSvaJJYV3hMIxjePT3rjE8Mxo3JlEXPQpLEknmBwc4
tRMktMP7z8szmTla3t/qKZL3BJ1kMY409bpn1obA5gH2PqaVulbF8dcnnrFN/wJ5
ehL/7VtHqgwQy6ArfK2yGD2nZXVq4SmJ/cQ61B6OMu+7Kh/k4C+nMfqLnasFsgNx
4dz3fS2gElux6xS7vaq9/GpbGHGL84VLkpa9fcL02nn3y6xscPAehJlagrZ4t46A
Qk3rdyBv/P7Eft7L93Sc94Y2O0EfgAe92uYHo2i6ZmY9yRm8pIgg5mfgitqN++hr
GCAjGwmoGJvw9CFhIYYjVESpjAP2XSK0UTzTmWgTxSfaEyYXCxAk7YOtpUJ7BFyv
tTnMC7u4SyCvpvlwuLRVCAOV3p73rB1TTBZby1+ydLWfqFY67O6+U0x8k9AYIMOo
yhklJD8/OHfKB/z4hqYH7yF9VSfN71Bs39YTkLVXTjf12s69V3XlShg7VOPQghv6
17rlwNEtNuXVBUVmr2iwJrEuDw8XKfWA9uM8C5G8D9X6JnhLNGpl1j/2RX9M8/kZ
lMjOMSCtPZWo8DBbdqbjzmYWi+dbSleZiD8/yWZPNNXvpyOhb5xplJtCYtLf5jTS
u7Uxh5G85c83UMUxCP42yJ1Z7ZzxSpLdgc+E1iTehQDOMtnMkA2ZpbbD+UwZv3FW
oKIENVe6JwRbEeu5wEyLWYlqOO7q6LyiJSRmnXAl+4sn17mjXG/gYL59UP1K8cak
TxwQvxoIu2KFyfOkmdrcXVBiqdF6KX9JjV0cqX4xnvyLAYECd1+yB91PgpQXODbS
sSf58MTKzgpqsUkVWPqyUzzECF+iW6IvTmLvWSMaklZLdgO3ptONDWXxZDtd8k55
Y7qKiI+8UOQBmrDgrPNdzrS9jJcnNE36jfsE8EF9/eeXY1Oe6mUSiFfLdSXc9f3s
veSed6IiBBL7vnNctxmhFsCF1RydPNwLus4psvz40JwYrQA7TMNpZIvXfePT+Q54
MkBU7zEzDKEuH/CMVsVp4CUyfQCwyZ6x5Yok5W5ghLSbgpuLwGbV/lU02tE8MD2x
mOxSisGXWNJbZYFLjOj8ok1FOxpb38g+GDCIhyifmzmi5zMJMJc3gA83RNWqi3SG
Kp/hFTAfTPLGE0s1Wo5xbJDp3I46u/xvYVtq8iGlF6FBc2wXA8Hw2kN37eDtL0X6
8gL/MxxTPugWSRmoPoM9CrfY6ss/5Uhp5nMKv7G73yywhRSoS6kgV1k+LokgV2vp
hakKxHhh0TqSrx2yJuJjgSCw+TlxqzkobGGZ/vrd1rDcAp/4o00H0UuTdaKiPpwP
qFwmR8JHqBXk6vnohsVfFrpR1vHkK9E1VFPnUyBVADOj4C/3XvxbCD21FKHibgh6
lSxQ2ZjVl3AQIgNX7j3wel22lqCyR0ZAb/8ETZPH6CxGCOpBqbjWyPjP6vnDxo11
eLUSEfWa3K0tlsRfRU2kpz2tVWc8rAZy7DbGKG7ylGWv1BgifIpckwoUkEHqEn1M
UC5Qrr+/2eGt9Mp2rcXUDxpcokL7NNHQ6nVPKodhAb5ngehSxO0029P9U7+DCVAF
8dNIzdXYmZRGTmul6t5kIuTaKwbDXB43XS1IiZ7VVZzHZt0JTOQWtk901kri3Lby
DmWRCkFcqfabcCOAfIApmJn8UMStR4/A/xFpRClfpfHchC8JOqIFVcGtTIXUQWg8
PMAHUaXd42RM7hT7R6ChsXw2FZe/jkR7FxePNsb/AvDxo0lf3pz1YEKLizZAE1Kp
FuaENRkKEBaq1jt76xM6eiqon4VHJS24guwpcXmKw0oQkThuFgmou1kfW9p2+EZP
dFbNkBFYW//MCQNmLPlDfu+i92F+E3LOd7jwTablwJi83s7CvJVbBtg61WSAdyOc
lbPMsnSYnhtp80hgO0sxHzaLSxy/qAyih0M8U9i2euPDJ7rZ7IxbHCwR5jqVCZoY
7K9fklN9262vOeYuRbQguboaAsCKF+nrY4nbrt+54laFhox3dEj/Btfp1HZMsb82
rQjnKh9Jrl6z+d2CpJsDQsEsFMlY8lmgyvktklJnAs1K/ZrIiicrwraYuFaKS8wg
QlZsjjyqL3kXmDZ1c00pkP6mBONcOF+5DHBIFDetulpbeCwkCp5R0C98G67OVxBl
g6wHncJlYcSw2tqy8UorY+iNYr++/5thjvHZJU3LIlfzRQ7VXs3BedKDH1bkvS7d
NS8+r6Rv1JRdeZD5NmPPM/g3NQtoS3CEy9r1CROUlIXg8nNKkKdbFN3xM9Ei1G1B
Ni2sRhURaPeshLh9Kf/cWsBFb7ZPl7P+xeZX14fVzOj06nMuQMDuyimrKAH5U/yo
HbldUDnOtHKKBRndbGOL208k7WgF0sRuPwIkPMJwS96lTkdgiLVg2AZO81gDAA3B
Ph+uUPEoVR4VlOG/jY4FjUCsA4ldKSreal7ezAkMZBG9KKVSxc46OWIOgZ96IOiY
7dB/umfz9ixS7n+5Z3fOE8CjDdva0GU/MSEcCWsowO2Ymd6mE3yQzv5OPNS3ufCB
je9rjRFNt59VztxbcRkMzQBWOiw1aby2+5kq6FVnhvvQCGKMudnNIrXnKhhrtZE8
H808QAox85nlFbasmkZ44fBvzKZMpLZVww0DuyDQDhDSNpKQXVJGGhw5BcJT/gvk
1oy1rHe4VxedLURveVoY9AVdvgVnxI7sixf3d8NSZt1muYi9xpYbZfKR+KSQnoU6
D8Q+JFEdefJ6SOoNycGVvy+Q+Y71SysdUiPtWpQYa3yQFD6+YUOGAmsMFD+yYDFB
n69GwQ8UHmcPjIk+VDYXXCQtg41Y1Jg0ieq545/+9z79RQRVLom8NHiwTSg858Du
sk0Sh/w48WtF3Y4x67676YQxuNWPp8hzRqLFAuCmmiYqszaNVVLg04v1IsjLg0dF
GHwqeUaVa8n5001+2chzVhWf9pORoSB5WAO5tI/iot6iV1hx7ffYIQBOXtfGmGub
RA90men0D/FZK4Rh2Jyw7mL4WfhdV+5yQEfmdyuPP44RSa0A6jADnKqr+Vl7/aO8
jh7I/ckesaA+ul6gAAINGLUkQ5G5uCEh6Q0oZ5023hk+YTkUlw2g0XkHabfXqTRc
6FuaQYlsD18SKavhzlIvqHOtNvK84sqq0/84+lIhlW4svPCVlrTrA3B6SUhjC0nm
m5Ir8yhSRxD3JY39TC/ZoPjw3gp6M06U4LHmfE55sLFD+WTKqjis1twSD+2Qr9ie
pAADO1JOo+rylkwGe868ePa7A1Qgz2CtcCChGHMcfBMyilFMQy3TPGmKS3PRsN72
7Al4YKudmZmtS4+F488mezngs/6dTThLS/T28oiv7Giv3R4N+W5kYyo27Bxg/IIH
L852U8MffUJBfCYNwihfbh6at883NXdHJ5PkLVh3uq+/1Ww/lc4brC8XIMMJ/SiV
O5gSFxWmtOSIivp13SFagu+t9rTlr+JJsY0qaMtvQMmB5aZUW894oe1IkKMUtQjz
oZQYsG7pO+Cmcpg0Gw+Vhs/1EPyiEPqU5fdfCj6FUvpRfjE8HVb87L897LUFs7qI
Vsmg0s83DZ6A30E2JJILYY66oDkoDzC1QAu7ys4g3AQG1EIYUS+xgGfj5x/RNzhr
EkSB8Qh1BuHwSqKGLqTMXJVGNoGsIrco5MqY+RIzYY0gv/6W/vMZRR3wYBMnAMAU
AYEYmBFDhjypzJ/afWtBZmDmC3WanN9FgmjeIuufwoFSG/csUhqYs96jZ6lzZmT3
5s30Ab6brF5dVrB9JCPNu9NVXhojvZyr8XqpfsQl+EfSfTGh85DHsWpfVJolznkJ
JWx1ZILFmF+8Ccd5K4NFR/urNHmb/cHom2oUuruskHUJfKFxfFuJfjXPIRCVaPK8
SkZvprZx7sZytsk+uCY5eg7+KAZfEw54d28jl8TwtRnQua1r13nwTthRWX7a39AY
Xh+J731Mu/q2XjqMTFoxuBub2YybjGOGDtWGuTDGQdZRnf3vPhL5CfmA5Uy/sr0L
SXrsikCw3S/znGDFHj2MMVG08BhsoShYkQgoFxJHGzYO1LzRBGthvxGO8DBr4+rP
79SdGcDNMp0VIQ3dvx+TG8/dW7o4jV5WtbDehnv8LV75cDqRzoUq/+VAQjXKG5tV
AOQWMXPlx+bcVAFPMpJ/S8RrcVulEYlV7PmDvx4EiLMxhCBoNGmVCAqnE0RM94Ix
7Zr5/dvmLUtfCpbh9+Yj0SrKELJ/IxFEmjaHNPvjjr/UbbuYjDkKUm9u1nOOXXfj
qbdwiknxFI1wOQvEZvbznLB2XT2LdwUFUsMrFDeG+G7hh/nU8W9TbsFUVjKWpqlI
bnReXQ5aCOBmmuJCPWXRvzDVDMl3+E/2ttm/hygUMhfTod8/w7zeVXFUCNZeATXG
BT4Z6XOwazW9/0OaT5Ny7c86RJEfgnsWuv7JVqMeFVKi8pS6dlTekgFUz5S4OIxh
A8R6gUIiXSx1YDsnD3wktIZz+kaQF56NeXB3/+dQ8q5Pn34ZywApZpPuUWuq9WKH
KbJQwOTA7rj/uE3gC1+55PkkgE2P29nXF02DdCxfi/DDKmLE9Q5DcWwkWV8h/6a2
F93xFj7gx7/zkqgjuLOU3AG/ViClAIeh+pL31yw5qbPNSBDQ1ccp/Em7hK0RICBD
Ht/INl9nm1S5bUPKmIfMZX4JFHs4RfyDasRYjkuzP44vOT1AYyOt55GYsxEBIBLn
mnVjRXicb8cEUEw9jGNGCNsBd9hicSvnFHt3pK0/F0hGRFxYvGodLB9Q2UeSGbcq
EOjAGF9DRLIFYITZyKxu6OaxW5R+xJ3RnayhXSgNrhtCf7iPOOlIkZty/QP2ucW6
7oQ8bV824ewTw3DaJrhG5Q5b/7NBV1GCqZd4MS+d93sXckZLQ2fro3y3M82PhPgD
aG9VBFdrSam5DO1Svch4P/TUXNTOwLuZIanv8uocXleGd5+KLRiLv7XLveULljvl
vRjpLpZlls3LR6x2j6f3rGUrQNptWr1HlVnSkfgzdudEUIZrIA6VrobCeTRUJZBM
j1rzkGeZ2MmTqztZAtLvfSt4Rjtdzj6wbQQoKVjw24BGqIdoA+pSW9C1pH7XX8LI
fcWWinFg2fqMv/GLFRT8UH8BawBx500fBuUzKrA+bGetd4bsNAMq8nVNmLZUHr89
/nnWzA+YtaQtcyzgccRBfL3nDO7gWp3RycD1CQZx8tQaUeRCWucH+e68xLDFtsNZ
W7dtIuu3+ipHjRpiuhgxXOAKarOda+l2Wyx38HWOxNsGmdcaZ+hxzjyH5PRRwVZV
rdSxXuJkm7fBwhKi4rOkSCxO3nuOpru0b5X5DMrRS17Sbsx0K+UlAzFZm+KPIw3O
s/cG5y1vFCAZEx+lBTbX4f6f0qKrix7ZtyFu34LKfUZTiDvhqO47zX5Wke5fDjHL
PDJIMnHnK24prCfvZ0x3CgNxoPzjc8bCKcZQF6JqvH2/1tMV8Yru3soS45xp5e2+
LcVcOI84Q/HG0abaDqmR9KUq1ejNSalLcyULiQw/WadWs0JeU5PHpM5GXNDavAHT
zQW+RXO79F8bOQK5cQpcAU01JUs7NaCOTHTdAHr6cKleDTcxhTElxeHGuYsLY0Hg
lByxelXup25Zxpi+VZrIkFt7qlFXqWaxPYm5Rp2nqIRoAhQU+KdgpYVN718dyHg4
o0q32mebuXX65N+UD+Y3aMA+oGknziqb5IKspVED6vPb9skUHh+/6QiUpHxb33Uz
0shQo1amKLd4YpGdKl8TVXeksaTdWX6il0BW3YCdkE28qzaoKQJNq+VYk618XdRq
PBS0nhM6+pAz48Z1uA1KoFa5BZY9s8bf5A8LcBpfqxxe0grFa+oEAvfgSonie7kJ
pX5A89U84WwOpJicdQzAo1k7nTSzrFhZ9cv8sUXlsbnhPW7oMTV0ErNVm2QqxdFI
9GLDAkVrXh7qZAIhUONrU/WU/vWQ87JirvVfbbrByN+TT3ppk1CkMtW+Ag+kmadv
CxD+yTddiqUR0zi+gksYQmYA1GmQXpa5lSe1kqVUO0iw0WiFmD1OiFcwhm0rgTJN
Cqr0weA+7BcCfgJWIkGgKvhIz+7W7h+mTGV8mgq2+0itTfuiZF5N+YXAJczG4Lot
FumEjC+4zxP9s7v5U739zU0O86soRojbMZQxYRduzttj0k2LeQNNWsbtxiRqFhMM
lYwlgeoa5XxCmnjoPnwlx7Nl9wkldHKmP58uGwSZWQYWyONq5L4n67u1WGTsumH2
ywd2HP4HmuP2Wft0w9bS2tln+STvfXGDvgQo2J7SraNHw/GDyDUuHX2bXRb/zoth
MA4hyX9sexpEpiQN27bUUl+7kanpcd6Yqp3dtsfYEhyo7ImcEyAdmhsMGYVWosBX
okgvPL7sbsWIKuKoUb8/tBskwHmXkZ0GJ0Hgp0JKLtm4ihpoKAduf6qDQCqsUMZ2
hKh7h9hFchlcoV0NpG9gPQT9RYo2ySZ+6u7e15Ra0Z/Tm7681HYYOjfZ9rJzGAvV
NNgVF5YleafE5Y0CT4c77g41rKgtYrfRn+BkhIMDDwdxFuMO3Z2UvNP6FdNwGRZd
wrmiIKVPaR7deHBPP1pyOcNm5ASS4r3CWJ8jgOG3tiG81xX1OsSoErGPAMoJl0bf
fMbiY1/6opYOJgeVyAr/OE1/VKM2an5zunMOPgIk4pQNulI6j0l74SlCB3B6ggzr
yEZQn814z8/g4R8oZ7LOel+G4vXQo+MSB12H69Elr+ZiZ+QiUk68t7UMfwYySH4w
mqLBrfey5LB7yVzE1vhmErXE99atnxV8dtEuuSa89Wg+6Z85g0sGPpVa2lXZWPqs
PoiNfwoNqFdDOopx0mCv3TO+05SjmIa4jbSYGHvXGuWbtbAIO9h0761fPELPKLR3
QN4ULhfztnYCuwj6c5vz8QJdxUp0YMNhIJD1/MulocDhZoQ8l8mJqVVLTElNsQNG
rUm4KeEPd9vFX7wmDUatbILVcgVthtImWX8uAbKpPXnjmsuP72wDF6xUTBl4CCPA
1xwmCp9vL+QwMQBvHThh31mYv7RxYhonBVVQjxRI/8jYTmPqPXUofhyTQufUH3mJ
fTBcuDz3H5voIK+EGt92WKoI4TM4xdQG10ZoTAcN/aVzGiundCOj96ZmBivAMVaA
/AQKiayO8+cTbHybKLATZYpvfuYZbGTv3IVo4z1uKwXsejvuS+1bIzyVEEdqG4uH
2H57mfsY/wCXXl4kyOJb7AZneiTLw8hDeucvfKZkRlOKISqvhn29ccQ9mrpPIJ56
+D4X6uh7BNvd/xAf912U8388uGXACx7AsKgyK5QlcaX2DUI7eUbvTW4cHWB+l6Xn
9J1uhlHitUJE9yWSgA7W7fCyOvomn21/GK9xPRI/zT36rEmaVlNSdU3YKs2/JlHb
L9lWB5YuEk/ETjnIB9KGA1rlTRjXcpMey0gZKA0BKKXIewnO18lPwX/CZz8eKl9u
dLhHGj8bRjTssNmNclYftAi4XLAj8Bj0zhUkbPJpoCNFy2FTZ+5Cvot2pZ5c3ujy
BKK1Rw29OG7xJ/yFojnB2A9SEN49zIMzaKY0qfJGXi6C5jaP4rRm41F1L+4H3UnU
QoZS8CeyXCklJU0ybzG6eDQQMZMuDLQAN2Ky+c8ghdPSvv+kAQrtOPxfhURc9htX
lG+W8+J8XV7wHpDcNnN4aKRp4vzVypLRjRXTYeLP4QNayQfhtxQCZpedSQr1jLcX
YWqfP2FYFyXuoyAeoNHXcImoLOGsjou6U3W+msN3CAuFzkpho8rxfsMQ3pZiWSSb
WJ5pA+8d6oT/+7VFGoNO1A==
`pragma protect end_protected
