// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
E4g5AI1SezmX4GKcJ1LuvJ1sXbvFA6s+yymM+BsKaDPiDwZIwxPl4wBUlNIdb3714rL5MtqclNM5
5Rb23+XrLvrabFul5ukj8zhpczo6s6t00VYZaPFsgmLCA8YZ1z+Ws25KlG/kMkaawVxayT4Y91UW
Dn2gIc1Nijs4r2x0VakwiII4qyR5oZS7R6oTAomLImIz2MfVU1nh+qLRYkrZqsTNXfllmQi5FNjn
k9kAVBADOfwq3r4W2bEo9/scPQ/+flv6eRB+2iVYCu5KSoSw1/eoisPhgVPAsybnNlbHCnQMwXz6
OFEz/QeMuLg9hvoAXn+UAQhi5wpLPltCEsR7ww==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
MuN/Fk7VerDqMvgtc2Uv1tYKeeVU4205v92D4SWPxzpNoTzg3ZrygtYrL41iTDnN/k0PZd80hYqg
Fr24Dw35TDr62gSyhJp7ixvMpeKNYcncS/S9Hf+ZLBXpZPf3y9+trWPZ/7My/tLWtC0W4i+Dm6Mm
zqex1PitQXS4xeOenrMrxCZxrqdttHRqlBPkgI/LtO4HVqu0n47cM0Q1zoNGmPNEQV6qJsORbRet
dLgI2K6RVFaMhAaRDP1/j5/6wUYHqoZDIxeyLof/bQ7gZZ4AbwbkCvHdLJAoovlGGNM9PYmjbr3d
2z4rjPoBmq8amGXwS6gPbq3n2Xnh8M2uPHnulX7mPN6ERE4QRvvMCHgZD1mLO9/Nx9cOPQJk11dy
6JeBzk/6t5vKA/AdDBpNM1KXPfpBYOD7nbVfs6ElurPfdpSgWgCCnlnyRiWsBHcXOwSIzSu4O6Sx
IKpT5TloNU7WYOjBYO5AHSrHcXb0F7+NOWIvml091/oSNakJDdo4uWCK8utP9aqzjG+yg1qo1DUN
nPiSWE9Jb1iC8riDqOI8PYG4zDym6OAHvuqLsiMSWcPxAZ865lFjhGAUZZnowbsE8Y3iR3gb5cNk
KA49zWbvGkWqT2mS4VF29s1yLSIIiLcUd9h4YBl2ICfHh/oX9/kaz42VtlO3rNVMLNUE74JHew0l
CPDey0CVNoG96ZDCalh4HXmJPHGJ3Vpeo32FNw7GfmcRAkaLTs5CVCBpyNpNI79H/WpCA+ljKAk5
62ay4XgiAWQ5w7FUCsBhOxDJA2m4dKcC6Cs7pmnUQMKgUUYCHGM8n3D0+Mo78EwBpk8FZkLOFfEe
npN3GVuDHhu1t7zARPTkh93wF+uqf6B4rKx4YI002XDegZo7FhGxVP2YWufOYghqZ0qAYzsqO3fI
1f6ehJlzY0yIpV6r+ZqRJKDCQMy9xVJ3iTkUhHtqM53AuRJX+GlU2GaeF6opoMPBCNecZEvQFXCW
CRz80rA3qjCNeiiLaX+mlRKxHBVcWKh+8YoAreUdeLGckC1Fw/ZhGrlsiqj8y5sz14CKnxoAwZ9T
mgfdD8VIwj2rQ3tV2+3/zlbmnnYPXgZex7fXcFkTuNj34uA5n+H1VLB+FvN3jNOwFOJn3KgmqKDA
PQbjyQ8s8v3zY91xROtg9AotIMTD2fa16qXCQgXgFH3eYzYvg4fBboM6Jzg+o9x1VpUlTPYnCfH9
FVXqg939JpZXcwjpAx8R5mfJTB/qstv41lW9B1juhr6Nh4oG+MkFa9kgQHOT9+yRQdsIAFgEUbTb
IGDu90dM3Gd9L2AtCCUvaHAjCFhCt2eLn7jSYAu5lKc5mC8I8IAvTc2R/NB69m1kiCG7n+jFTBfm
gOLvqc+7S7RXTgD9X2btN4E8ubtg0ivWwFG9pyEMziuwo/TpoRlTG3E2EDPhPc/rHw3eXRfxzFgE
H0kB9J/0V3gGu+y/f9UKwpbpQP42UuUxHb1TMfaZtc46nra1D+Af6bK5+HK3l6FU6vWa0chScpo0
/jia3vUSCq4c+CY8H8YO78WXS37+s4O0olJ4qLvubKjUaq9GsduXsOZ9ufIh3yhq9SHcgothYDxT
qcsZ7nFbulgN8CmSZT4xJ9LpM2D85CbY03rqSljMudT2R4Ip4hVgg1bV9Z+COFBYnl/SVSOx4E9Y
HQ/xAYVppEXPwHBjNK29S093Aw9/Y9XxUbzwUCBekD3dWBAiuqdTIY6fx3vKbQp048hMehxqxEpk
FRqalHiSvvLZdgpGXsu9Q5UWLHFGbRyhT+p7ix7K5K5u6vfmBuloAM2wAcRQHNjONmEUTNy0ILNU
e88aDErgsztEry5irt4Bdfv0JqRLz+sZVH3hZ7HlnwqlETbHHwKPdalIvAzntwbL+f8f+0UdE0NY
Kn0ro0Z0L/d0sfNqM68Rs4yq1sb5PAbPzmqrL4HU86tOz1PK4JG3ClYigFq3BeB2HdS2Yyn7IaMk
6293ghPSx9jq6rQGtoKehVDaOo+5uqTV4cZZKUhE0Eet391SFly5V5ZbR1tZBmMnh/Bb0sknN3Zl
pzxhIrKqydJ0XESJx1PbMIZCcQl0L20xlHnce6OvVt1LAwsnkzv37VfXjOvbeeoKGpd417OZDEvS
Fh3fdFqlfUX2OCLtrcAOju7FtFAbT/f0YBKIJWzVlhgoyAtM6un2lEIol8qW2as96UdnxwSRdbE8
h60LLEOICTkUcwCfCz6Q86UrBc4o1SUPKAgA73v56zKO8WCsvD/w0lxJEOUHaXUNNrn4ZEBQVkig
+/AlItlKNII1s9npnwwv9uI8lbG3MBVKX6hXA3aKpEA8ECaCC2Dd1pwMjGLP93crEkG9j2pHlfX0
pDOOHLBnQFLwT9yWrB08I/xLW6AoUWsiH1tQ/2hrIYSFAWSXh3vsOzdV1nLMyln+YreBNs/VmvHi
esqjRZN+aK3/iM0cne9unObCVqgn7PtvwDDkcD3O2Of+A6Lq/Vg5FO/np2V1Bpf4GWI4Psnkbpnj
hLxVdsk2v6GuTuokbKO4J7Vrrzba1z851UENvX5eAkeY1EQcASFyQALwg6+UwH9UGM+d4kYZiPg0
b2d0OvOpt3NNIFzAGexYZeIKTg+NLsNNAjv1pnI0dMGMy2gbIEf8tE3bvjLrcbFj29Q11DNSBRH5
4muLRiXxqVi+mN9eXq3s0MN4n7addIDxIXwhQzRpdxrShs/Ai54LbjBHT/tMQEtJ31n8JZZG2pvY
GZ1rNtb+v9ErDLnrK1I7iVQDd/y+ym3OiFc+vebhXypIGI9eIy8yYCQknuQb5iaqDQRAx00C18Hk
Uff98BbhW6k9jY/RaG3LvOneFITIwc5lW5janzpnQ2+z2cVPPzgfIcqeJvqHkzuwR52Le/a4HJQ1
f+ysEyTFenOBg+6Ose7h8B5rW2nkGGp5cI8JnVqRuM7yP1rNA2fUtBf8W8ir4J3LgpCwsjAqMacO
keHYJujaqlJ/k4+Lc9cMD5RENz7QOcBMq5D0s4Hqy1u1PKOVDnfLpJzSCMAkbJepdNqaeOLhQLsT
4w2XtBNNH1PuARikwabhd1wudrLtySlAAYzfBLt2jlPVqPNw31bHjFSrzDphqcQGrjjA3q049NEz
IXIf0h8Jgav3RBVhTX81Fy2TnUHE79I1+eMy1hBK7zbOi/IoMAq7lWOI09MdjCI7VoWeqp6ZxA74
V3idQ30qK3rwBM2tkLUsKQPJk0t04b2pLIxt37mAUJS+pvrYQLofMTpVmz8WV4IxudKOKbRRrgqD
6K0JRpxqibF9fIK1nSObRbNJ5INx5egi91uNCmJNm/ALPhv1ZBvyNACZwpvXBrKjUxF84m2QNcvH
IoQd+mafDg9DHtht/fQ1yotKYbB7uipwh9hUa9K1HZyO9pvjfxutu6y0sXC8i08zVF/f8GWhKA+k
o/NNEwl5fzleiwGAHg8qCWXfGHDRiyD3BeqOvlmMmgm9gxS+JeS8Omt/XOMjzcu1Jxdub7LUN5CP
sB8wkwDYKiKwbJlnAVfsO9m96PoP92Zt06juTgQWTIWdGXu+kp+HBMgUt4jMTHfju2pjYCbsK8gQ
C0IVWf10QnlCoAiniZ8sEp+zkEg7d7FMW3n0qQj1OVuOTcRc8cm/EYkfz4LT05OIQjOyt/MFF3X9
exmf6Ifb5N8VrQzA9anDCjdG18h6Fht0OvCGI3HcbRamNtrwrZGbntPH4+eLp2eBXS++ABIz3KIE
9wTGblD/0wm/2SDacXrfab45B7K2KQTgiqTZtD7yOobYqlVdcTMoe9blf4olrYcLTNpX6qbWnp8A
N7k5jP7RsHZCrsOTmkpch5WgAUG0LS/jPX3Eezjamy4bvrWpjlQH6w4XUdSfJZWdox9QzP6i+O01
gfLQUrXThOlO2f7rTsGr6p2pqzGFN4OQdWpNq7vxfQm+eltvtpqxolQFiiwfaNHCNEJkgmfgV0v9
NcYD8x2Z/y1IoNeCH08dJBJ7MWokABsVFDH0CcXSFJGbe/AeNsf3XjPeVZrZNNFP0dRTTBtJqsPt
ibxY5H/ssru9pEg3vVI5gaM6ga6crVeLPGuYbWdFELy6CPhFf8t7kKOchv0y6lffVvh/QlnRXcju
C0cfisC/DJamCC3FECAlpS730Zlb6gua23QO9iUpH2CvUMrGGnocqwDrbupv+n7NlZSpg6MA/4iS
4FJRDm81lkfZ2RghZsGzIQ5iMaxzB15iSb6aLZZ9M5x2lXPtbHibP6KXTcOJvP5XjhdGe0TC7D4E
XB30FoEQReiJw6uC5W3NBmH37hJPeWptR59Mfl8ejpbwjoUhE+x5wJ4uqrr4+ir+idzbz8K330lJ
w64XScuQNmFaHZahynKCRYRJ798y9Swhr6QRUC0VG/H+phDAx2vWjbMdF4eplppEEjy2kd+PgZNO
+BHxHq1bd2GRmhOd6vPOm6dIqrpXUv2J0e6Co5nOc58UJ8Gk5v/6C/uEUkZVUfNd7ou6FesDQOXT
sdlOfQ2t9IGS2gL17yJCV16CSVCq2qGm8cTLdUR5443L99cj1jiWgpZ8Hb3t834t96MHElIUeaDI
C6iVUetooJl4SbZksnu27jm5JoHWNK5KzeYfR3cRBlo7kDVUNOrIPiynUY9DASq8kBRvNcy1ISe8
x/raaUEqMRUU3nTaZgRI7S9MwDQw9olwBKdnp2GlUmX3f8jNS6CeGszTXXywPx0HP5/SSWjYRNz2
eBNG1laJRMKULd2Mi8EUtFf+dfz0Y6Sn3cQvDW/YT3SC1E+mnlR3VdPpfxmvyobngs/SqWSc7uLW
da9G/+Xwl20VLHKbpYooAeoBVSPlxP5AWydJavRcAibBoyrLzpHCUBm21jI9OrPoKRTWs6ULNGl/
9NMUZYaBkaLqiW7D7dRSqBXAx8+/CVVOVdoSq5sQgH2dwgHqtUZkqXNtkbRRI8oIDpiF8FM489ro
0WtxtLm72iFWhCer40zCsK9xgcERMGzlyKJHG328lCwZWavTics9Ad0ZXqUiSVlNnnXFjHgDAYaw
4dEGjKP8/HWGPkhFugEdQBuqI6rbMBf4u0IPmeqdnhuvv+xwT8gC3gnMPwDCvScZZWXLalpwkLoN
T0CL7coXNkoVX9E7TRpKiJtU7rmHabCSVEdHiDsiJTQInvgkhp1QAqs3ofHZtSKiL2UtBBSdKr4z
F2wOcVGYn0MhOb9RAFrxQgHwAWw/j6LwtiB5lSW8vWt3b7uwyGkL0aAGbgvEOlzHXRFGeRmwN4HW
7Du0iUX42WbTkpyYvoy6UmLf2yloYTJc4oebyed279ZzEh69mkKMgg/P0v8GXORwXOzL+L7PDZ20
l46uYEYSyx06gaMRPFTrFhoqdtw0BFRJPc5eJhAEruE3F4I69C3ZXL8wpOwTDWFC0MO9YPon0YK4
ZJN8g9CqupNmegqg02qVtE+HTsWBtH8AtndomNKAM0zsId6WAXDuG5GQTZ5TJXNJcDlp6IME3yKl
fo2kDbip9zBDywvgmJ9O35BlolXu8O34zwPgIOVz+lH0m5qfr0kpNRh63BqdNOspH2zOSa0kmFPc
GSJK6gJ5WxFQyvI28zsx6onYCOfkTrNiNyKdhMCbysGuzD7fRnYRxA7eEnbO4doZ6rm3xkmTJY4c
+RfxbIlS2xMO4NLTtddRrBaIGM4bTe65O+iFVVYR3YiAzLFLWOxNc9Ph/BRo5PfzBf4JmUE2p6dq
F9K/rj8LDzLpbeqDM+gtlVHdiB8wRHQu64B3585eYsinAhhOhRolpfmbwC7fPTqbub/rihWC6eop
niNzKsBuLmHj6t34On3SHyqkQQ2LomA80WqMjs1/MFru94CsTYFbRwhTdd5CjdfLCueT/8yj8Lae
NIuMTt84720BEfXbPqz+bj1bbShJfl16HRyrsw+eOCXEuKHXhPg4shFAljkZsa2Zl+bppxy/mU5Y
uBkUyxXXf3hA8QWWBUM9WLW+vjgqRFYHkd2hF8ms2fuiEjJAKD7PPZ7FGn+JK2qOL6dqnlRxiir/
HSqoY83oH9uzdFb5BiwrF18JY8rm5Dg2g06OMhVGWqDmk/28M3F7YmljOxHpuXsg/fVRz1cRwMuz
hBZHw08w2hz6DvAYWB5jGlKXb9CsQ2vlGSrGDr2zCF8v+Iv21JVWGPM+/FypErK7GMb20igVG6mo
g/ikZiFmQAxxUMs3YGyn46Tez85dq+CKDslzEKtJhRcnbtbWWZx45VTrVsysXpcKipbUJc57uj81
KDQx5d9TGenDg8actp4rzHX9TFQ9GQDtRT+DKItIKR6baqWoQg6CuUeHQcvKIaCo6r4xI3iSfX+F
Hd/ZCRLm4Y0KYKlIJdGflAK/80qbY2hTMpLpx/cz2SBT3Lnw2prOUwsxReYRkeF5C8X/6ZEbBlaY
IOmHepF4gPtjv6wkat303uBYkF7nMQPKVq0ux7Vo+rv+tGfrUHrGDi7kXheGtgGOFdbGxOwK1Aa0
0xEctL4DaBlNMtXCnXah6NWXYO6xfgExYRM+CTihCNyKASGbvVGADoi3dWEehKsYNj6FwreZf42w
rW6oVXPUMvFAqwf24ODuSfdmnTQPa4LgTTCrmsEXabesyblYjmCXsHajJsOMSTpy/ek+oAjwtdFi
tgyIEDbNq4UHC21qJ7cCjoWfhGqR91zdTeLN4c8t0EP2YfWcq0+NP0XmJdVcNj+ne61dYT1D35BB
R/b7uS9JhI0ftTmN+sKQ4FtkuYN5cI4kGodRv2R9h2zdEMTtopdgzQQWw+0EM3gAsTp3SlcQb/2f
vf2z1IhZuI36BBHpaA+GpUTUza1G1bG4Gje1F7PrtqnvE+gyYblXAh+TEnhQFX7/OHQffACrKpkw
gHn4rS8OYRQFZ+ae9iHQWyaY43RSMhiGbZ51pogbc28uGXmLyNEMQZExzOWNRaGz76zT0ZyZCViM
ENL+GuURLsOSybFLnm4udqGYkS1xsg+UjceNnM4G1iaabzhWXBB8QSZ0HCHI4TVevI9FOBApAA7U
TTcj7NduoVZhnRjbQn1NpKnO2loAuMKm1UHi8hCR78KCJOH2UKwBr1bAPIl5rTMWtPLdOw4ZCS29
wheVNGkJHM7IcZ0rPFVAqEzv1I4N4A2yJ5WgzdfxFtbLj3432jk00Fc22FRoCjTymDjJkWvnosfC
IYKFeYxtRdnqs1rHrtJYCDoIy92KwkFT9tP8cGEt877pO74cW3h8f9VNi+eukgXqllxp5GEX5zW9
4E9J00EyolS46WaWutCY3dZRYmMthNzk1V/3SDy/1da3NeI7YLnpGbTmKfR5EOAJPlbWh5JQqcRu
44H0uFPoISh0Xx5YtzziMXwH32FSYby/QPfnjpRmbfmViVmleKGICxYDcRLvcFTYOTARn4ZVdLfg
0MtVGvM7mPP++TZAsGGN4dIH0y7etgws4AgwMdDkIScnYNX+awCTKLXnw/7USrqPJITMbLM+0ESO
F3NEUnnGIeT92BhUzlbPncn76Cp/vIBppRa8tBbt8LF6tmaIZnCIP2q6qfnVeg==
`pragma protect end_protected
