// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:16 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
U+EcflmR8IMGSEFT/XMucDZg4NWkTCwtU7uDdy/XRvSfomqlqq76NGr/lCODfSBU
Ey/pYOJ5dIJEGjFe0lNmjS4Y3SDdPMW9lZQVRbH053reCmO9ZB8sKDogDAfuAg/+
6tCSJr/iXttZ0ZY5QeRrruurA+6GDcXrwNPmmJXPMhs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 68128)
0SIzfXYiqBqf173Yi5Br+h3/k0FzlSWVa39nKTjLDEirsM/eX9KBIeV8aXAtXzSw
GrgGk3LrkAtZT+VJM3YmfGVM5pc0xF+MBfLLqXjcDrKdiQQnPAfyUPUVp1BxsAe8
lQ7WVm6tcK21LSewV6TLMl+e9/bhOWlvmglC2Gw7r1aSprXrfwh3VY2cducvoo1c
C+4JNCaAuYi6vKcfQ3lvFSVcCwSax4dyaDui4LW4Lmh8296XlMS1QotzV33u9PBk
UGLbVHvE5Y85WxMnSftyF+QdSz9NEZTUEC0ohrB0jsG0ysBk4Fe1aCzwsH52KEUV
byj0+8yV9p3qczhDGo2fEsPJIy1iwCKvjUjgGrxRV3R/uC7f2HjQVx7B8uV9Rto8
UPFVhJC+2Yhmxr5k9Gfa9rTIJbmxXXjPGV8jNcmcZUsIBD9bL1NxR3H3vM9Qcsaa
3Ejf1sdxBGg0OtqGuhssjt27K0UFuVx9e49JLYHzuQ24+/yPsJjaoMm+f1thXHXs
C21+5rG8Y7OJMbqmpIL+ZpCYsmKBOVdK43MUJB9+dT+32Bha/hvobce7sihol1VA
1aNhZlR8bR+gsNjLwzB/SWl0vgI5bE18NwuRC245g9Wn72jqqnZMJDN1BfLPC7Le
gosum31qDJqpS/VGNQ8LnO8OHHJFlaGLTHscCJeOozBDNFTHj1lCFfmPWpEueZu8
6mI1SXxVgegz53oAucnrlQ0/jHaNzoZBb8GL7yVPUGYFfAvrru8xAdp8PwIj0On7
N3ygRwlFloBa4VAoPngVa09mwSGrNAn+VMp2isllOIlUutMbK8TU5u9KbE4tfPId
Tk+ficjGp74Uea0gzys/0eVfJe8swdgq0MrRgAQwwq5ZXQ9VMWgoMzqO83QN7/5H
XGMSjcUzDBKUjs7YIFw37vxQ+ew57GtgI5LpYtcbndolf4iOaXNpuYcVlYry7O9w
IYxxhpVq4Y62bcqdRZ9DAkMn0NJAmAdRzJA8tfwXWHpZM/Nk9kjCIhrGxUfAPTP6
45cyC0/xCL3Ssvxuy7zxGf4xFJwno2/OD8RAouMnTC441GCdhYcqwtXqfmOaBDje
94pDgGIjPQ6Cu63SNw7qapBVOExwNAJBl8nPtUS6QafhozyjKOJBGPUBD5fYRuU0
P3BeoopqcpDcpHmapWJy96Ce/T1xYgTTYRdIHRkhZWzZzAgFd92OoBITSRWLm4eq
i7r2o3MN9ZVByfcQflq1P2TR5a/C5QIj04ioFa/WIRZPxY4TA4C6zFV7msdFysSC
9P93QrMCLsSPbe7IGPiCvJzl529NFr945xQlSvmtX2Jj8lXAri1oBP4z7nprUqv0
xD5hIxMCBfQgfDnPftBLrVkWEhwFYFRCKn94WTCF8NsL1vi9wYkzBaqK+gBlsuKJ
sf8/mkALvPjriFWrtxR1HttuUstnsppSxn4Hhm8ShS13JLU86CHiU2GrTRvGpT5T
bbZrex9cJY+MfewxfSEeIuTQ9UNz8iiuG/ynbX6SDjLTVSv2nRvKsU5jbInpLUra
6Gn3UIWeMsP+q9hfhgY5jwXGLlYggn0HKYAMwHguayf4bn6/MAPez7Sof0HHpIpp
fl5MrXCFhS/1f1r2lsIfPyfZ1rW4v8EEdibIMmY0/D0NHgrCWjglxdQGOu7UXCZT
H5/wcv6L/sUGss8yMM+5dVqXUC7AZvyLhxv7APsLedcPTWBiBaQLGxx0GdFOKPxe
9dSQm3euwMuUEtq3r3Z5oVlqP9BPs8jgfdpJcrAnL65T7BuQTSZqeZQd3wEG7Y3Q
cNCWCDWCgj33ngcd3ksJNpXH5baKGc6NUziGZsKcaAFSRpVuPnxSp7JZjQeZAhl4
2zfzQX4u+SGyvg/IgtC88tejTV9Eg5vYStKWtLCkB9Q7leZizHZTwLw0JmWdvaT7
IxwVklRIaQW+X+MsaNmr+HXxmYy2N2HVC5BTArVt57ScNo+6rVq1wWPZMH9a8ZdH
QetaABRr6qPNlQP6RCt8ugALWwGNMIe4+K+cCpCTwyFeqC2ckuEp8cyARU602RlU
7pimsW3E6LtYEpnM1pFkeGwfYY/TcyHr8RCkAb+a5coQcEcoVEaWNS1uMmQfMah4
Hd2MrRKpdDs79uVYrVEqyE84+v69PyVJJU87uiLANqQw/6VDZVrVjeOgo4NqA7Oy
EAkaBwO/vIm8YEPplGiYaeX96UKSWN714VYIQEcBxFlvHXPjil0Bod4RHYxyAM0L
VqZvxelITEszlpnsYb/KiiDkFjF+aL9TTNpfETrEl1wcScrh780xta+yeu/xInVJ
v72FYnHNJnyww21fPFwBppnjcAfAiTtsEp5GnVGT8WK2Y24yzvuruiZCX1djqPh9
LqlBYzaTjdOJieFodLztqjR2v+MsOtbVT78PPPB2qfomPRVyuDFFyggjKBqHFCq7
y43/2WLZFWNJnqCuxyJIxZZmbPSXMbI0CT+JTv1paB6ENHDVqLOR24O57HptbyJv
hYn5QJl+5rK+Lh5j/wVXkNyuUS3KsUQolpSkOnurxQVQtJNaedmCwnUFsqR5m/Qz
x97uonMAr4KZ8IFkD0Bq/ZAUMtilUQIXI5qUpCd5tk115TGmUQlEkZpipOVodm0S
y1xOxidlgJ9YTR/XU5QjbFvBIoBSClacpvK52AZ6RBbh511kGjd8ruwnTyuMVQkH
wCV+7E+Echj+pJ4kBdT6Vx9crPBJQ66mz59+xnlKY5Xumk6AkP4U7CWBhgfYvVQ7
AeAYGzZmNjkT5cmOcQg2G+c2+4ldifDCzUwuStThOOXl25IB21yPvDRq5A8d1GuG
djElcmBWaVqezpy3OKku3i73I1AN5ck06xFMWdXk5Pk2rRtixrbhWZqMd2yWTNXP
rpT/LfU6IW7pg3s2FtPru+M0gJgn9UeKk6MBTWPqeEpKFJ7SxMVism6KSxbPZbYm
0Dkh9cFA3VqtYwuZfXlwGkyuoKN2f6661G0JRZmc2nCFHOEOTT2kD21OWu40OUKR
qJTU/9c6ZdRGo6RYlCiLh8UOrgY4ek722CTsTFN5DV0NnVzw52JmcguCTCNyDByB
lcPrf34XA+dYBEz5s1+JWEZk3xm6wSxv28o5DUI9U9xhq0vp9diwDV9UtYMKzrY2
HzOa/AACAEjUdXI/OxDs7QeJPzAvVyd/ksuX6XhE0b6nB9x++fIchj1WUEIEKYns
spEzmoJPUzuyWKtE9i5CVsBK0gE1UkH6QVfn0+z+7RyiKlb+UrugndtrhIazns6v
83N1y8q3VVF1c/FG9njCF17j17JLnoTTTEIyFfKDD/bpmnNvb81W0L//LZJWgCGN
Q5Mbi35vC9X/clqq+RwqXAgH4uqDUXW0Gpyl/Syd7/eYJF81Rr6rH97ldGQweE9q
dRaH2ySfKQNFXd3hvLEubLq5al1ya3D7KEdYX5QTpi3EsK2Lq2xxkS5pTW94N3HK
ITO+sg7KwuV2Ijbs4xJmDOGnJMiv049cegT5m8kmmDBd89yY+iG8aOUB6y2yHNCf
Wk4xWTDQIu/312Pvo8YrXsnLKxBKn3+kOsH/vyIEf79bUtXuzXOBgdF8ey02ycYp
2Qx4Mxkj2qI2bJ1AujqogdNlo7nX+4YDLshrrSzuoSTb9kMFdaC6zNxRPMV2LDJB
I1R9cp16XegLEmfKH6Psecy4yyTUBKwFiS4KjrWLNjVxVuM+RubiQG1so4wHglTZ
u9vFasxNFbEyNJyZlqw/7Vdv0JCm7MqBCSqhXdtBvyChlk4WFBsuBSGai4WSgQGU
sHdSzRaibxs0BEM9igAoMu8ntfkMAV0aLBfMccKgsOzysi5lWazjHlP0Aiutn6T9
gK+xhRz9gv2uXMY3yZ7vTSAIXoEMFFnP7ZSKK4TslukOFaEl+EkR+9+XW1YJyC5C
Qi76L25paS08vsYoG46bfW4eOeyLQB6K+ILDZk6sMUG3Bv2X1SG3FcqclMa2MjRe
Fs7Hr7w+WfTQo7jU3380/ylMryrf/JGX0+D5oeThPVLRw250mBX7RdIg1bomdckk
uzGJWSuWUxHOBviWXde1Mqky30DeXli4pMCNwKcLtavnggU8s9OBEXu3HjEgMQ7p
O1nOvtPylvz3MyKL8ntVldXYQ7Z9U1He574lKLLwdd1fDDztFep8NY79PGuW+qtt
ehFGoXduumWi2sz4bP0xiMJVcuIX90isZtA66/6cWDE4UEy9z/83LILX6LroFii3
nKGpqdL2KoWa62Ca4j2KXWLswCE22ZFnUtH/i8zmXQazwge9gp8Vn62AjiXiYoQ5
7O7umWGxUdN8JVyl9PVkCaQc/ATYTYaTrZTny5oN7hpllVcvRBnLXtVCy2LNHSJr
eRjbmWhkzXAAxhZqklT3CMU+0H1XGYJjrLI7C3p/vHXjeKUFbUj0gu4LdnMmA5Ow
8rKqAZrIlPirWfhLCWmjeATGcnuWBIXmXTl9VQSRBxbFOOuScC0iIbQlDwj9VWtZ
xGF7GqAA2BjAUNF+he/XKLBFK1ZgvkX4bTaSosJHrpg7Pv2KPFQC/FcedCZTWeRb
PBmNoNbywoAyQ0IvOXeeEpgAStTByJ7fJKk4HuleP4RoWuUGiqOGEzdzspZVnftA
3iOqMoJJeIzjfVYLuuWqW5E26MpCEWJaJllW58a3RI1x5Nkxa38jhJZiJB2e6H+w
9cQDxRauosfUD+ffIYsHTLMIoVZDBp5we2B7rucIyQmgwIrXrurHdmrtSLtUvmBu
j9wV8HQeaoQkHDV7uc5KSXrZ1FFF0s+8KajxviQwyPC8MIlbLUNi1fahErGJNAWJ
gHaTG+tWprZ/sGUedZZ541Pie7FlQ/d6ebywpmpaLMp04qBwIm/KlDHO917ZHD5r
09vonpR5O8gUkOkqQ7dxKXU9o5+0rAxXvRLNK7eS+YUKKD4+bDurbX+KhW64crEW
ygipdeIiY681gdR+C7M93MtGUmTtQKmD3df6iaWq0SfcPPsDiUgirDtTa/X5fmz9
QLuwKdSbITia4UNVTWx6u/4Syw1DG3agB9R5jVixpbRfhkb8JIphfVKo2UiVt+0A
x6cUpApQr2Ecos0wf4UQZdiRYMALU2JPt9LFyvU5jjXakdgTXA1Ieru6uVLmsA0m
I6fjnlqSI3kHXi31Bbbqizp5LNXJTLe5Oaw1xIU1xrQQ1uWbkAgq25qMnTpXPfGS
7P69CKp4cculN9peg18kXUGMkZDTjildi8hLUJU7rq4VHw3CsFVaVDgXMjYsiEr6
KozqawswoIpXxYD6pf+p9zgPHJi1xnj/uxjZpR6rV+8JGpuPG3zeQDtrMkwE41PH
VKEbflOqgSd12A3RP7SrHTX8lFzTg3OPqMZQVqnEjsJzIDoiNR+ktGMuyR8zQS1N
ENp+RCmM91bAD2tCqLN16b4OaoQe8RyW9HaJUMoB0qKNqkz1csgYfm68ebpZdg+O
OzJ3ANhBYxcM3AY900UEbrrH9atN8nYVvGt9Elt57jaDzjfxL9gJa8r2ySLYylnt
dyLq/FlqmL1vY5U29TDWH/FtYwttmpeYyXA1VcoIa+KkRwxsaR274TJ1C4UjrLIt
j9lY5LLz0e/UhVumJp3cMJAlrBV4asQsQCP7dugWmrg9i7zq7ciwFVVXkC31sKCE
AC7u6dcXY7k7mKAyDP2WjHYqV7Y03cOum8Mm3RQVJ1iLx5q8YBWMXu2tOWBhzKnq
Zxi0yqhfU2fm4qqfV6+bn4RE+QC6jdvjCA3LL2LE0sXKiWaZEk3rVo2Otgz4D/6E
kxZwnqqbWNQlWUYRCxc88tdyUPOAZy9xBC95SXpNTGyNHFn2720Md43XgCLutWzE
IxPxciJ+8GjXNCiIVHx7GID1PvDj5Di4KEYF8avKlpYvngIJtov+MjtJrHNcGe7g
9fQ5Mz5XWQqxCToAUA8w/7dRd3cuQsmR+D6U01ZA0B4Buvma6RisIiJz6Tn+0beb
rPCGUTaWOXLPgAlEze7s0VDAOsEACMEpq2pIJBLjpHjJyN4F8j8nYXEymnXL6vat
WcwlgqfJWXpR/oc3XlOz9mlkC5AhzJrmlSKwRVmVok0eSGMpQEOywqrDifHhco1B
/E4EhIl9SRq7XiWsIdF6GsqZu3h4Di+wn0OH4coHRZpT04XgWG7uh1l5pah5Wax5
miWQN9tWIlH/5PwuXALJ33VfT29CwCTkxApmQhm3SeiJb2o22GrlXUl3S/1sCEDW
6H+PMXhTrftv6A45ZpsPjKFr0Qbn+whFBivwMqFQeiQ526irBZcUoJUUwKK081rU
gtSPUDGtN8Zdkpd4IcBdY3HPTe6M7RZQT659A7zLpdhGBnnLYToV2EHzCStuQqPB
uFRGd5Y6AB2Dk85Y2xorF6gHE1QEKBYP85G++tRXQ9s9qkvl2VEkTi9D13qQCs4Z
cSeAV5aUcJoXvHix04p39CKSaMjEYfjgnYQeEWUFDGexUK5hMPHjylhxFpZxoBFJ
0ITelE4MX0NJN0koZSpphIpC4fRlHylQ0Egvt5tQ93tociNIA1SNyPNE8zSqH1/+
aeuwWXqPEXDYylZ+n6nyqQZtXM8UF2tGClCDYi7zZ5BWsLoIH+2RbmXjYdYiDbX6
m5YIF2iUzTrMZ+o3v52qYFvhNjEPfXBSXKDjof+BHKunep1QUEa73jkD10VAiHiH
AcWpusrEiTBL0ySSUqpCFvoGPlPlrskmFF0n8aXBrfDjqRAD97WrtF+pjWYCv54Y
BU/AySUVUrx8s4yyLoTi7GMG1pKG3hkN917SL1uTTFpVIBS379isnMvHHOmWnyTC
BiBFfzuEmccb2dFXlvB8BtYk016dGrgZaHNrwYX6tPu8oK1PK6srZb8bL4jyAaDT
OJZgq7GC+tgw21pf/KOn92tsSAs0miVWQV2pNwdoUP8q3qV/fRl6b2e3/KOL2V64
fQuwqg6tvXunjWONL5AmAagb3rmXzh01iYmK+TfgyWlLLosR+KS9aDG67ZNRUiNH
DAq3bcJGtHju/vs1UasS0dIYiZ4GYh8ubdAtIdS/73bffNKRSTRENS+v2lewdRhV
ClH8vpNzJN43spSrurbNIr0Wb/nqxc3DpZry2Ok6FucvpoA0voSd+hNeFb/1qfbP
l9VsFMMJzF7uyjTlB+EFKQgEzw8c/3TMJeYf0KgMD2qjc+stPD29BC/H0EtTNY9+
UU61Xdzn3wYV6DC0spt1wSVwELRh3y9lXATWETe/j08Vbzt0KL4Jh1SKyhUlTbcT
A+JGJIeZNphSwrSZD9Cf0p2AqN/UEibLP4EUgkOblI5QP4lBbEJpBRfzBD5zz5vA
2bKHZsQyppgQGBQ8tDJ932K65KuJaJsAbUgbhEPxBkAWyZeXb4N85ZBM5m9vhEHV
yVuTcQV7BHyMogrC+SuGhonPEd//NZQE2on94QGSxCIubfodQ1Dg+EkB5astMeCm
2dHacBnpL58hYjIWek2944arPK+E9uKlbOUhvKJseF7AiskdAsn+vvbGgIpbsn0i
ct9sFy1qu3DVbkIAq3aGZgr2ukegQJtwIubP3bt0OBV1QO9REtxwJQgZkWmuOVUB
MQ/pu7KA24js7XNXWamAkoh4tMI0Kf1cqPnKjE3K1Y7TFDpyp9dnPYcoOYZ6iof0
j+R9Hx5s+sKBtesr0OMJuDzLUhcfY+S7roB9ocT4FWY6q1qBT7WPj0x9iaPkQHhO
o6ZS4wi8gTXYy0+5hHNqdgK349yYZNr+52CvldHfH+839uVr5/ucQ6KMGiYtdP0i
gNHXpqB38TKa06bFdmTtPOYqDJpyjUrKA9JhZ32O4tMT+nDO21nBIARf4hAbMV0Q
ewRioPy9OcPOyqin4AlV9RlXV5cHn0vCDV8LQgkTyiJxHG7OtFM1zv3phH8wTx7h
DmI1z/uEUXUuKVn1mGtm6dcpOWGz2x4YRuvuBIyV/00i5hKGMpo+dhyP9wZIUDWq
uD8lFjmO2bBo36MheJgnRLIwOWC+yoKNlZTwIPqRK9txb8tiFBCc6WXIOcr7Ll2p
eeMK9PHXBgAOKisCI0t6s6arqUxTX3uxd4a48xECe3rbu6MpvOjorHwYK6h6pdfY
PNR8zOhTsRWMwZGxDbQwIsNSjwdqto9u6WYdLbl5Vs1hO1y/WaHdvgIg63Jn4rOg
Em829TMdQ2QMweTDASzVMvj4q2W0ccBsiP2DBfUrSyBITHgllzykHMlSU1ScB3Mz
4ottHfvl4QfIAeKfl7Nemfab9ISDv884hLGSIVY3+QD3ojTaFKBy2kGv6hUxBriz
6ymWhiR+PHO2CHJoJDpK48RMkEp+vieXfRGpPuLENp4RFbg8xHoxQI6NLGlPAZm9
3EYAVA9zgVVp5V1YLIezD1DvO2DtZvHKb3juOhzIySb20hJTw80An0wJMKAYkK04
JfpIlieqqbxcfxjY2+pZwUp25s+Ix3h1YDsr78Rfy3Jap7En5qz2rOCKz99iNn/V
RU2Tf9Ss/kDdZ47obsjqQM7xw72uCHftjSzKVnCEePcag43a2qzMA400hB+3WVJU
ymmMFTOWryvgqHP8aZM9RpB1nJ/HSWsPoGt+ILa1HlHYyvGMoYAMsvO22kFjisqE
TFm3wky/uHPziXOONsbuNjugUjGeLpmtH9nbduCykCI7fV3LGs08m7F4/BNk2cef
IUtcmXlU3JrT7DcB9DKt/UiaKtYD6l4cWnLMeUJNNwpO9rUvXsLTzF87plIUt1sB
rjmBpnhGP8+TzeNwhuoJKxV11a22oFvUtDKLrhwHZca4zIXHoJmSmqaWKiJ2vJaz
Ht4MdpXettzpPsqktxV5dMNngd2Pd7I6FNHvVfx4sKUrodUygV85/3mojhbRlohL
mJoPN2ZPquJ8MiM7EzOkVRBhPMo7heIkptHwpwnTUsfvNi8xizzZmFfd/ptq/zjp
ichtj39EYOAJVzEX5HYG2LSGdfW5r9gfBPyw6r4SXmhW3zuCqbDUM26+g5ncuCTa
YqD3GC2qKYIya8qvXBTmhe4UjJFWe7QSBfZnh81/l5iRjI8PHZhOUoO5BrzBthud
dZKDv87iFb4fGwOJH2iJYrAu+EEPyiEzj7z8v2+Lc2XZdfE7jUY45GZ4oVJha4B/
Zl0V13c1+BHZsaVEC/hu94owJY1Q+NKo9SLf39Q7YN+xZ8JL9elg2FCs/8zMzNDo
RQS9LiEFnu7yoF81ev0olDFWxaH1abOJJHMO2gRhGqxB0NHYjF+YKITHf0uaBhs/
in4i5pR3tim3DD90GOhrAOMBoQ+bcxYFwW9pEluaTNOOW2n9n/eOBGPIJ22K26eu
U8usCK0UoeObdp1aAGiMBdKyuxJjQB5pzuJCizCn6YAx3YB2pt2wm7prs+jTbHjc
tVPR9XkrCuXaJ63YaT5gvf01qgaisDwJ31BE3TtE0TT6zKPgL6bZq/tG9+Hll0r1
uAoZifVw6cw6yApgX4FwOzeILUWHfXdpgR0TQK2aWHJ68U4XX8P8h6yKJqt+eGtJ
JUlwhtH0ShtxlJlKrTTCFMM9DTO47QWZiKYfdoEf7oUc5jeMuDbYI2FWnxuYuFD/
0SP+nDt5Dc7k4iPPuL7r6HXhglXQkwP/j7f5dLW2jjIapINvA110MifUclbz/5Zl
s9n3kpT4D/RUWVWwgEJe+BxD+y0ZKQTnUsaOPwdiqq0sZfehBFvoYyOKDV65rkqq
LDcv1diOneK+XckZqbt+7q19dx4YQM0ht35mJWEHzbw1UUox2yxIOlPzZYvWI7VT
CHOQNYxKbYB4S1lEXe2ZPrurBJnPobtmAkTyL8NgCddtJuGAqmXa0ntX1CQqeVrK
gWa9Iwj/6r8PENlLw2Ac7s5Wqtxi3OFXNHg0oTE3FoQCfmBNHwAy68efvUQnfCVv
Ff9hIXKVk0WvPEu2w0yPUaaTUR1v2G3vKMBJgP8bt/+dTRLI63D9AwudwMyl1Ml1
pB2gS1DZVnUmeTIDuzAts5VY55oIfasMAbMKJgiQWqBS77C1xJ7SSfd1lnjYgGOq
cSxBMf2UjMiJwJe5wrKue6OLudlmUGzdIROofX/vGHmFsmp49XxxNgcaEbPcyibY
yHBt0S78ipRHFIBLcQHIXxff4ZMUEk2oUseaFoR6cMqFFA2Ea4pyXwVQ9HdI0WNA
hoX8uVHDgr24CW2kb5n4Hvu3EZqbAlVeqXymc7DQ2CakOFPW2uKcmGrEs649D0Ht
L61QfnXsTXBC9syjIHxoIZrdniSoBCw7H6ZeFnvJ12i70GSXSW+2MiT62nwWfknU
vE/mF1LHovzEE8g5RYGd/f4KawjnluZ1QOXuSWPC1y2CQBtJhPTCI5zAwge15yc6
9FntJ6CuwNQH5PQ0CE4rU7o7BppKZsH4mQehjmikkLZnppudVT1qlF9QpplWI0Lw
qaQizqgcn92qNMFrdNC9bcfi6+VpOQsX/9sQ9aicGUFhHGZkkkZqJFyyM6pgWU/X
Og+coIjBtg2BOMYcpQqk1PVbNCpx9ESEOprCoEseuSFGomndlQ7zNBJqtafzf4g2
RQqeQ8rpH+lQDJW8muWUhX0VOhyQBfPqZpL7lLR3YtIfza03J9QSzE+zEmCDszVG
/IVXKr7+h5/b5hPsen+yiP76D25LNqG+8RWUyeR/PE0gTV/g/vrH7DbXj+1wZQpW
EuyN/DfMZwiUBSUJkQwAYXKCXxoYrA/PqWF15fc1linvcnWT5XL9BNGtdUoV1W6+
VikzEzSD4AS+/aqdIZm1QVx5Gf7wAjcYrQR5WQzQq7w5LW/OfVCGJWQgzhyL6LEm
3PQjcsUPeE/Q5+gYM7ffQFRrAgcqFdhvpBFpnGDlUc8ghYIXp7Tsyo7q893wyFxN
ueaCJ6xu1wVvoO0ZBIU3eiYpRwe8UOMWjryLb8xYFaetMnlYQbI/gKhpnPwBhde5
m82TS5YcqPyhaGImfG3CByBvx8Yujrv0q9ISoNQjJeGlspO6CjHNy9ItzWBKofJ1
M+OLD/Hh7Ib8rN714DiEJOET+ytZDBIs/znDVgm1NYpL8W5HwgoZWHppoDSozFd/
a+NrUpr3nOiKiO/E6br1M8xwD/8I1/GdGzuVT8+uTxhtSs9zzbVFw8fbPCvPWF1O
1iZEM6v9qnStDrpBWul/inC9TA4t+y0OPoIMooHjNaAHHGHPfnGXb7grvesQX7rE
FlqokLotH6P1t/8EywX8XiKq7LsF0BXDuKKzlCjjUaLNnLbTQ6sNGKl2G5tSghol
MBp0HZjeIzwaC4QCBLrDwFNfG9ik1E71NRhxbLiei/rSriU/lg2RX5XcmUqZTNQT
ktu2GoaXemIzksIZN0K/PppQMYZ21+JW8RD2Vw2c/ioAXzdp7NK8BX6OaSM5xLo8
+o7LKfZIXsw+Nc/sR1D2po8uE31Sh0OHYwxLWxyNgmh4XAPW/c4LEaIIrIcx/ss0
oAil3zHHUHwjALeh88AoJZ7Yx9zlodgo0PUvI+ZMZcQFbdqDtT2fNOKuG64NC/gI
M12wGowMByzp6y3Zll+PSt5kSEHaFn1PupV3kEawRiGoZS2hiJzUk3ayjCmXfTwp
bKNfVQyP+nDwZjKTkJRyafDVqSecS20CC6o19/AkslNMgXIBqZ9HTjpJW0xChGyv
ZHJYSYL8061EAoFt52oprf6nQycCRNvUGvtKYq7lyGaNUaInjfzyX/wnl27O9Biv
rwpWeCYgG/ZQgXSxdJZDQJtTS2TbcFhPccTj7cv7ZatM3LfwbUVWlw/KYIF6405Q
hw0eglOD5KB7/bva5e6oRLVQkzdKu4AIo3D/XDcqJ1bv2taCNp41vFx4P/D3S9Ah
/3n+6eIEj9dRZoPSuQwtFd89PYz9ejWxsR8VtlB31nMSysh6UCiaHwaFaSKcE2hT
vY/uVbNKyyFTpb+xhXLf47dxHxRbKPA7bOlPLs3KKsccEXj05yD3v0p3SAGQXu9L
1uSHsCy9ZThLB2nQi4o7wDxRlOk4C3ApvD0jMC3zbDme2MWrCkz9qvv7LYP/ZuxL
uHmZ9eVWummBDgNuogId+S9dTMdx2vBWHvqaCqZvMzuYWhKqzq9wjcDBTMtbNUOH
scf5eZBEfmvGrUuO9uAw8L12cLydmhsTtXswHG60CyWufFHUxxyT78CPsv4tTU92
Ia9BTQ4Y9WPNDhGFwd0hcYy9EibudrkHtv9diNQfCcKxFPPO4w5Onsw6dMOSmq9x
Ap/K5s1ouneeIRZ+GomenCbo6slmbC8uBwOI3s2GM4RKLABwtUi2XElhfHKMOivi
YwAxlrD+FTyvo1YVZUtmQ/3f/bXkEPJY+tiH4PjkVuDEJ81NKrCEm3bdT2WMGOev
QT6RDjwWfEQMB+6+RDcogXQbjXL1qyuc6/5dySRL9enS/GkxJwBKcp4aJ07/SL7K
ZiVODBF6+PfjQAv2ZVui8T0PTKZyxJ6+ihASNFXJWg2OOMGhe+gD4yhUmt1Uapoa
EadhMMiO07z2dAyIhp+/MMqbW+XRBIPdHfZmQpnoEEevO5P+reDhHpcNC9oc8Nj5
RF8lVGHkg6r4tozPtt7EDqdZz/hGSe63vaUgDdIOQUCXuLBpF1MzoH7JdsUyPzl1
9HlqEajhtR2GrPv3MbTjI/zS9yRlzKdJQdRkqGaDix79N/GuZeUvq6k5HKNfvvci
zqvV4fXu6e42IdqtsrF4FrtP0kzllD4zhgNh9KpVLz6gc+rgxrJuZcrntAMGkUQy
5BIb2CQcfxkpjGWx3q1XFMqo8cy/+aWoTTEV0ikpgk3nURDerBn4B8jTZ8Idh+OE
KJ9ITmgWwS5zatxpQA9jDRT+HyPiYxHr994eKwlHJ/ssla6xPlN4NZ/TgeYJZczq
ZozcOorzSR8TLQYSDMH2BRtxQt2Uw+0j6kkFf5cFn0sqUTAuOzEV6HAL1uSVfnyI
JlyICJViR/Z+kFd3yO/gHMb6BCjFZnpEvCZLQLPvCoIYHjbpmVEZAZbv6x1bgdhc
7RxeLGy9X3TXWlQ8ytfdkXskbFAHzOIAtO3gECGhaB2jq8Uv9STSLNzaj3NLZiJs
wSv5/CinRISJedFX3ORuw2MfV4552HGboydfnRZAj8ADOMKmtXP/ADzxczDNCsDC
KytuYPCm4MrJtHyQ2TdQNZRDiWxcpBXvPf6FwcCwLfHU1prJguj9Q9tuOxjDfht2
SwvjoeZw8lOY2n/kH9ceBzhlBC3AglkbLqnSn/3YLIEm9BOXPmqW72SK3qdn6R6h
hadrG2jDbeAWFOjxWx2Zv9mMp+nJIzlraGIHnqhDBC8OU9QdMzcCbUQgHcMCI+ps
BUAze+s0nF4vHU8SIVHSMtKKlzmykuZGgSZNfe49xnb+0a5oQgRpIMZ9tGRL850U
OgSz1Da8afzUenpBiWhXseCI3gHuWiAZcsp1UqAetJ9JsqMmkgSkUQyi46D+atUy
nlbHFuEVjvDU1vlJuT4IEYm/6eJyaAWa+Nr0thAiZ5IR4HGSF6dZwvfxDqMGPShX
s+j1FFFgMO09QTpI8gyA7VwwgK1epkT2n4kNGyV5dulkKfT9WlIyRBCx0LMiAmnj
goarfCpTwfnRzUG6+03EdQU8Xhez9hZeNc037tGs468GjEWcxdODXMGPjRQrcD4e
BYi+Z4fOqmdt7e58Vv/dL28DQHgELW+cn5RJH3b3x4WZxYeYaK/Gx8q4STBXuC7c
uVKS7Au43xX5uuZTiNGevhqP81RZ3NlsNIt0iEZZbXniTaab5xp3NFv8CbJqwwUU
WAwstWKk2ypOHvitg/Fqx8CiblBXVqNla/mRuIiRNrUduKeODWvbSwp2HwafBOWB
+9WJtf/vCzZun/oKemZJ2ALC+twyQSEKbHyQpDvz1JuK/0eDsBpynOFvUTuXHDdK
MZK9PgbyNzVc/UJqG2MRU1FGpUu4ZuLzWMp2HKA+6X9ym9WDWAFWFPcAg4im3dKS
ER3u5PpkxoBLZIPmdLlvlbvwH6HCo1FqcWqkSJzVsKu9whM4LSxMG3CGdxy8kfk5
ytLEkDcz7ld8CQUeOB02Glvmp+WVASsm+9NReeGPtwuceSw9oOTA7apT5/TKil2j
DkXnPIBjvu9R/a5GTkNPZty9plT4IxZsPmgFW/+ePAv0pwdDyQGLS5Apn4cnQVgk
VbzLIGiD4hClr3WfLPVOXwF8nt48cnR6AkjBJfS+vdzjQXbw9mlVD2T5tosrbeDX
B0JbqY4sc799AiOCMK+axxi9JE5Dy+BVM/ei9DknovQd+8IP4dbQBxkRAE3JPqQT
uHXzzYfxPNHFXGchEJf9cVDX+OA4c+X8hD/SLfdqBW9V4WB44SKI2tTFubaW5hVY
844uiwP6M3rYiHRbDQRGMK+djNpX07JU0Jeu7rj+FtdP8TsmyVJhGykP2uhbeVLB
ENkGrgI3Nmm3oT1sCODih/CDgV85cKvb5+1mW5gG6/6DliRLBMFx/CPQ1/pG8xmM
ytQifBb4ngO+tqb1pLOsnLDRdxklfVOLoFpzrTeDVdlAFF0FgOKhg0UAkfAy+8a2
cdUQ5SOeZqyT/YSgLGKMjf+kf2PiY6QffExjqTkGlmJrQuLQBWOew62eTQDpeh8n
+GPt/2rdmEdyU/6bKwWBPH8UC5+7wZ5iJHjhctLjTMPizK1MX1k7pd2DhEnrPyxp
+CW3l1l6kCGQbIQIZFxDN6ktv64d86aM4NQskGm01e5B3Y1nh7dLjyHwXc4NZbWg
C+3f68Pmp8ep3iGgmuBkEb6oOnKli0hBXJ9YBNNgG7Kl4TmXvaNl6bBWw04elJHg
qiFLBdwvi2/+oStCJK/tITFmg6xQMPzM8Oki/S7HN48w9PY6zv4XGE1JsOtXVTnJ
Zp3bpsd1Dm8BU+AE4bHDRMeOwEssJYlWEdcc8XFliO6akNwMkzc2jWNXAGn0DdDn
XuQxgIPUv1uxRaKApBGYdKFszcTDWjB6hbBWaC8ZNPZ82RANwdN9Tp8C0x8Gm682
84vRgkprG3IGvo6cP1BW0oKaETKwwSqcsYL1lVaR7FvpAIDlqx987ur0GUz+cU8Z
U7YfgkOc1hbqCoFtqV8MwPXDkQg+0bTGUgHVz96HaFd/aGSZ0PmAQhvmKhy9pkYz
LSvrPDuP3fW/9hQeS457yg8fK2jq2vf01D+pB8e/HaRu/+u7+O8kr407G3by5W4L
IqkuKR9dhlj+ZsFOvalsP+GWcwufzO+dlrictoysQu4/0mpR/zUWjFplFEaInZ9W
0JUGuH0w94hi9Nx+hVrt12B2pvm72Kq9GxncDhRnQbttaL+h2mw/le4MUP8+dq1L
6J+aYGez/IUkhs8h0/faU2GiGxuBGgIWZxp63LhYQCCqXIZB5kpvkj/MNkK84U95
62okDNQ1fX5yTD1RtoXlGPZt6lVuDfifbyeINJBERtujeRE2K2+JZRGGAxAw0h21
rLKjHFQd5vslnlhmqwZWx9Iur1JfMZz0f2hcbI12/tod6VfXNJJ5aLh02icfSYBL
1MuY75dgQlkRQAmd08rdkRQbEAtDJn0OpQswsNaxIwhJ+i9/xXWvR3g9ldlvXtUk
AJ6Z9+Z7C8ikANqvFCRu63MkhWL67YldsvXPpZFqnONBTJwTceTqQForOfhiOyA1
vj4zX0HoNiUVNOPjUywCKy6mtawiMnAhXKl1YwkiQ2S/fu9gmC1Ko+lcXFbbBhNu
GBBYqM/wYN3XhG1SCZ3tbw5CifKwea+ZzAjawJFhMyHDs4iFjrIEUdF1a7Xwc5Lu
ymmnZjZaKReijKh4R6+EpPiXQwfo/ODuesglAvcQz7VWqJOVXFflwbjbFOb1y7sd
HplikhZ59PVZJEiO9Eu8xbp3DtdBsONBl001M5MNICOQkvbN5BCNRXyA5tyHn51u
M6lrfogZm4CtjN/eSOgF4ozuSb1aSUdwwjiTHLZsiSOF+NJbp0gG844QaNjcB6lj
s31AteXDfi9j21RfFRZWdoBOrvdN5BGFOxKAjDnN1Kr0gBat6OKZNOvXnN+HHKRY
Kujo3XX/QnBxXXfNC8JKxo2Ok9uKXgTkSiRI2p5hu3pu0R2q4ntFg7mmzrTDxQVf
G2h2aKs4QHcyUV7GezI8LSk6+86oVILm602uCSv+0N+VO4B/uhBnqTkIuu+Rh9wF
QBPr6HIKIbeUKbNe29saF+1DoF+ZhhXS9u5kL3X/VIHv2YMsnCeE+bsPfwSFUEYZ
atW52R4Z3Gr6GPcCD+Wx+QnMbeF3v0HbkVn2T/Wwc+EqJHU0JAWUBzLe5yJdLZ+f
59qVbfxxHIJXcb5R7nigKgAbeYOWl1jgLID2dfnqgJU2RwLElJ4aJUirgOLK2X1i
VeJBzeBC9857j5CFDpsFPsYnxhec6qfSiwCjY1RGg59o83UubNtjmu6Pvnmn+tTN
yMi9vPGHjv3S0K8hezI67NK352Ogv0BsqJjAfem15iFeBNjDZh5+PvbvpWg3xmmi
toYnZHk9rjlMXHxKsedr8etd8vF/K53W0eeJfLu6FJSx3ujsEeKDH2UUcRmAYFNM
mOiJAC1obXsWxz704ESGAFvylItvrN5V9wF/iZoHX5Nrwk4ZQ2emiRpfiFuw+PcM
m9zGg9ha67pdQNUbPXfbRbSikB+oxYIWn17ztwaEr/aACYlPIDHofBb6AfqZKctr
8EKAiiZLVBsKKR1HO/UCCqPPy57z5SctxyXa5Q7K4WGJp6nT5QuzGNi1uAzj3pWi
78j/7lDWTAOfaTBixSbfUmlwwzcHRIZFdNmVPCpUC4mMyqvdZCnM74LVoO+xGfoR
FTFwl5RPq3+pvwm1kfBa+lu1rDnCaZ4D8Sb40UNB9fbYYDiEo/3VThTc8D3PQuOI
dHGHCNbE8pJ9paLaCTF1h3+Fg184coSMUjX/NOgEvNkKuulECf1OLbhuZDMnZYjL
+qybXkZk3yzLM7dsT061yEidwcMULy5cFZp6wgwIE40lFy1uhC8kauE+DiTiNHnA
T7rNu34J/WHPrSSB1Xl/levGEPJhqDz5qm8zNgMeAOMWVoWbjtBh1pbExKiaJR/Y
S984gC5eJBc7QCR36n28bJo8WmJDZHRasb1kDWTRkZHqZV30x3jn9ymx1F4KsuQZ
bSn4OtnIytnbbqiPJkHEModUTJfm9NoSp/JZpYTLKUT5Xc6U3ZGiKdUK0ohDIGx5
mOw5zfUJBGq4xRCFaG5tNFZDruJ3IxMJjJDDk8oNsSjd6oibVHu7Cl1sOyoPoD3s
lRUGu3x6jSOdIMg7RpLluMcL6NRnDMEAOGRcbJNq1aCtzySdUdP/Va5IH6arl+g6
x8eA1mjjNfEvzthAx2p6VqFdzor+L+2Wth//tdISdEz/yeZW/htqMeU62aVgaYb1
5H/gg+Rd/HdE7a72VdrLOChSIEGjkQQjm56h1FGMU9Ue5dVwQ/ouWYnsAtU9oxqS
BEKUteqNqhGP2V6a2G8xxI1g7t5ZobJjQroSW6f6OgDpdbGaHUi2wCgOyVZpaa7G
XCDG44r+r65rYP4kDZhkPGzoDrx1hOdTLBCWhMH+omnJPxFi+YN4Ev5j5KN3pybZ
5m0LOhl4QFztrN6/DW12B9qNbqDdhnnQtv5k7ZjudL5wMHR6FYDVm5sJ4u4gjVOx
M24l8RayHHB+Pe4FgGAK/xRUH422Lo1191Zm5jGZOLHhayA2dy0QP7CJzWM07Vvl
ZqV/bA8AiMhb1E3r3xxTr46rPuq26rZxH/Cl8mDeRIHydEuFOOqkG6dNPcrWSqUR
CLSJQx0hL9GvpIPl+HwYNPsJSBJBaQzwNBK/YbzmN8D118C5SyIndugYUxVTWiOW
xoxQpYRSXSMZi6l6Y53d9/Zu73AQBiJ7KvJec6AfUoNejo754HmlUU5zbXKBIDRv
DVMGte7I9bfFjeU6ckHjlLyMW7kvzytTnb7e+CmJGgBurR3XkWXzppfySCHENPnp
5XtLaWExmngVttMXKRlddKE6EEu2AlyFnMtBxFg95NhsG7JjUodvw+ZHaqLPqW4F
3AtMrj8Cvu0dTXaJuRKFEPcM2eB6CIEy9WLYedjKEyciwNHSyYDXX8zEWGjK0dGU
clICdI/PkiX3fUygwjx6nXJiSUzyhoGwyTHZxWHIB9mVYHp1UoqkhfVOhgMxipku
VrEzs3wZ0FRc83rM9a4t0H1hbYSh5aCnUvSObRbm5FHWwX6qU1itVwwTggRG3e+Y
rweMT1idHsQZqKo7+7g0HP73va/d30UpjM7ZMKdA5y+SHLXvr+l3cxi4+FrXNEY3
WKMGCMns2IoNDn+QMa1Snt4eA2huaHT3Stk6J26URcoZn2YYGiZh55D+wo1969wf
llqu88rIkr/R2tw8oxKm67uVftTEz1fcXQD+DQhhP29vo7cyDaUdjR0ZkMFzNZkM
yVtQSvLhKmcZ0aATQb3mjvAHmZFuSg2fvjyPSozkPae5fIZ6bCjdO1n1b7JTU5QQ
q7M/9vPpFD5Qugxja3yYVL0Aafm2zl/Hpp5zun/sC0EkrCMVBtsnDYiEfJD4rAxt
DxfdqxSM6bqXc5s0a2FZ8hYUvhtB6K8Qvm82ylMiYgo9cwpDSbBHPAbxLtN6fA3t
URXfmFURfaPwBre2HE9sxARGgpz49f4h8n92385XA3y5vjvBzNfJ9hSWgFlBvnKL
6Ay3RrwgvilMCmCpNrdagvv/CluhtMRIsvWetlTxHBQ52o5fcr5mF3Dm/uhOINWc
J9dnKRS1WF/MVfMDZmQpCh9hFYo6PKiBKv5jFQneD05dmImwrAgS2UmUrEZujSUK
PR9R8/3v34YA+sjeGr6Ci9CTFsOwYNfdhfztUM8LDCgaP0ErYjKgzAztlLnnzp4k
fg9DeswI7/NUR782nugrcl/wH25w0gNQrqfJ0bIcgHMlptrF41iQpHaZkKuVYeV0
HCaN4dyrP6iHvp3eMGz3Ug6xXn9MgEJ2qCAitEmdwAYuGGo6XRVCBj+Jq9zEaujB
N50dKBmNlRR/1VmGOTgxYOsffHy1Qb9t/VDBfaHksXOwrSPn98hStmsZ0yQPnPYu
0jVOw9FM17K6bfiCACiP6o819dpPqgzwuykB7dBPlijSO1n7w+k3h5VtjBHNb6fY
3hjE7SQgNUMkI9jgW+nTd4DAdeAAPW+vRQR0F2G5toDpX6weQjsqeaCbEq96LOm2
lYFBhZkleYeIizhO4pPGypzBGeXM+ZraqMNFVTdhHzz+AJpiducOVzxEY9Yrsryf
/dK3znhXzDiWHnWY8LX25fcTImXGI8h8qL92QYSbLbqbsFpkhKZI4lAQXony74/x
oBY8CDza6tP0zWTZTI9zJk22mOyixOwa7kCXJcaOB/m+V//Apwmo4wenxt97r5PU
ZX4bjxwir9HCa3gZvNqRLYer0ya2McPdPZi9s9dXDpJTL4VnVWrYBPcPNtIP42BJ
ZaW1iceQDcPtjiofHauT5Z/O6/CApAQ+HxfWTU+/lbZ3KNIr5VBZKIyfAnk9BGRe
EozNqnm0dFpPFvTBQg2KkeHXXbI20wPZkBEqdRJVibyHFD7C2oFWl9DH8SjcnpTo
8HEN8V51TjgGGhxRxb4B7bJytZz9cZfRzqrAiWNtJznr3YxTxnu0jsg+DH3I08TX
jCS7NZBboOQG37frh9m9bkeOBG7hIwiBTb0gOZp9eez+fixeD7ZZqx3qleiQJwkW
4U+s3EsoO6OBBbSNQmWXNVE2RDamBlsmgFbMgoxLHoIokYH913WobxcbEkmQHUQO
CPQHLRWxvLCCQw65HuMvfH2+jv+5nUT0FH9nNEP2Q0Xbi6UiRdYN9oJ0Gp9IcdWi
GZYGMr5SwLKeAOGoHz/rXLmW33gOGb+N2tbYn+k+1pqvTf9U10FUB4mychVdA6W3
jZGAMvbrB+7wTi0l7NwCV9lz8xoNkufxdxETWUUA8iQS7SkwHiS10ce4zd7Wvgz/
xqUSzxTrR2wgKJU9bFlkBV0c3TQD0+qmls5peTRO78vhJ8oixT29jGHvfrn5YEaz
pHOt+8GAjNSXgyIdSVYVF1pJYW4Nzl0kv2aaVKToF6vFjxcqs9rLuXcSuCuD4ZiC
aKCZjiF2HzVHxDAjV883qx+cADBRI8MUBscN3jIOhJF78Ez67dAAVIwpO1cdSGSp
qw5z1VdVcxx4hStDtCvTUQyZk79yc58L31YpBqnH5zoJ9AuTd36LkzfA0KrtUYC0
0F248YW/Pff1iB24J6eLWbBCWIt/sejbQu+2LKxN5Urolr3krTtio7fAiYtpA9ev
tJO4kcHF17DYepWaiSbtaabboHezbVVFQTNIOs2i1wP+sqGPY9uyOxy/UgM7N4Ka
jbomcjg4/+Kfa4R5+ITR+a8diR/wjET8bYhRSUnWC3cbsnCiSJFhdi1YFDmeDVWk
IT31FwnCMuFXMhRbjC0dI0WS51RAwY5urXQO6RWpP4F2QEMSPVvbTmJTaaD2yCn5
Aq6JNMMZgWuxKzS1lAUQ1wMBDiKvuN8csPY3fvn0Dvxa+0J8zhyrvOORuANAJRTJ
Dsd0UfVXPwMuKX5FpM0QOKAwkPaILeCflOm3I/SlF1SBn0uo0D5BiPt/GZcZmls8
lGII5rkCqA20SaMTO5UfWV1+GdBuNlNxKaDqH1P+MaQ4Q7NspHuvGDD25cfia9OM
eA5u01s2OUDdQoS9AEyOKn/DfXl92G2vFtyX2PgFJ43GlJ6RKhvCfhc+lyshZm1o
swqZMplNzlJ52YoLy6BuHHncBXol8RKLUOTQo0HDGsl84mQDz0f8XXMnFF/pP1ZR
xGDfzZUIaNjwBshvGoStJDGsjRbd1Ymu16WQBUWkOEz2aRp6NiTojZh6INAP6Uaf
fGpNud5uBsI4dYnNzS4j9/ucwnfyljs/rjDlqxXCoVB25ReIYCW8g8ZnesFHzw8Y
kEWfPBHHnQs0mF+8tJnZk4xcKjqnavc+w0NJ/6D97NKJjnHg9odCiDHAvzIrJXjD
7HlFUZrpBjzLjSjsBtHlTS5U1ukF6gX03AogcXe9TwBHkEXPbz6tws/UdBHK0EgB
cKOvg/CWvaNJA3jVBDAjxp6J05RC0Ee7eFWSOLFbB4x2asIF9weFzFtef3G47NBk
MakgVaDA9nu/JXRLXha0TUWNT2WidzGiDPRQkJK2rpyBv08ehsY4gVUFSa8AUo0M
SaO7cRoSHYGmbXcZtdeCtsxzV41PRxeRe1ySKx5QLZ8wdco+T2GRJx2F8ZNuWhXC
ECD3D/WRyO4c1v+aQZoQG6VIdsjyiyFyx5/+oyknYlb+JFtl+8c7i+ZoYhsaNPxM
O9UWNX9CxxnjNHfOqUEjwuzVbbPJYfuXWa92h+cAi7iHoh/LGI2+CxwoLiKGpp2x
UoPY7UqzSHVyq4ZJ8GLo1sH0F25n3OZxoPU2bLkpyk2vBV7WFtwKarqMl6jHGlZX
ZEAbuZFXI7pi7+HuW2HkvpYyu0rED5ABbtXFOvJPYzy7skpifuRpaSfqgqUybbiz
C8L1dy5rBczIWCAntYn3no8ZExncCejH0RRsw3fMg9lgJ+7JDLacV+dLlHjw+yXa
xcQxyAkM/uR639T5Vj7G0J+yPdpX6V8smGuYT/MxmtfbnhCGXFssUzR4ONomCz8x
bM9WnDPXbRvSHvPzwdISihJhD6mVIC+dFD6ciiwTntBdTkcSKDimKjX5H27ABGrb
KeJ39vhvUXUbcCEXF55JYaMhaJU0fFEY1/7ycEfqZeLX8kvUTU7wule3HTAKmLpe
/6KRAAWKMTxKNuJFvnQu8uCkPKuK24+eKSUqQGs6nalrfwYlZat7KqPaQZW5grRU
eex7jX3YZ8gJ2p+ZJQ3U8+VRXjhlTrwhAnnLvPAVQulle3wNLHH5z9mt8U826Xkg
dZhe2ut16iM/OJw5MThtRzzFgAsiyfrYbZHbxiDJDP7lYHXwatro1es1kGKhjCm2
o/DP6IlJbyx4ZVifToCTmphdSqQS50w0+nQ53SHOVoi1E3auxWaFhzVRcvonC8pc
1evJeUfHLulyhtWma462QdvvHovjawCIHHYMPgnPQ12y5bcA2JxDu8eOkY4XT35b
oDPWB1GsPCwENVZiGh63UWKfr+7HxX/5Qhc4duDfwh8eQJgqeSWbDSgJ4MDzPLX4
hhGdvzyEP+Ex5R9nrpN4JVDTiOkEJZW+oEEpQ8pVYkw1m8W5ATP//eqa1GB43G3v
Hu7+N46L6hD55QItdXDhpPGgfKbJZv1lJMS2GWNdKyuIy79gA0FuUFrtOfyRemFD
iputv2Cb72CcPHgHD7UFz2bZ/dMcJNmUgoL3ogO7n5Sq1fs0+wLv1baZvp1tnNkh
6vrw7T/pm+4x8M28n73OppNdgaMBub5dV917wgTQHtxIgpWx8FtVG3LMWcAURr8F
XVYhpWSCnV5r4yrtzW012cSix4bjkcHlgJ8jkqQWv2mmXKZNDj20QRJuvXVUOkbv
CPD+hH8YseZuwf4jOdBd39CkSTEu+n3hRrzhUI6PKcE5Y00JqsXSjUmlwIE05yth
NYzcTLmCIoDiA8E9KDInzlH3Z3fhOcGm/PI5rB12CbyFCRPwEXpSHv+KPOQIsvZf
SOsBmHSBWb7b4EPRwYGWAdVR9vVBIpYJCl3MLLaH98Skz/+hWCR37h1APgs+e1Fx
cDk19Sdwf8gd3zgczSdt3qj1IcfrNfrvIp/ogcTpbew6pg6XfSIlDKRBbxOXBnfe
tso0EMiwxauEiLY4lwG49ev3Gu6tGsxytzq8koffx0qEQ16pbv7POGfgVWfVABTe
LZHBWCumQMMn+57Mf/yje8hQzFmwodKkNawKrGB34jjWC5JHwwmx1XWsO4B1DAqe
Ik/okaSYk6qIShT8ke9EbrGStl3hZ6KS/jkyb7IBb9q8mNoPQg6MT+Dliskdd3zu
n6q7xa9mD66tm25xM6+33ilt7/lBDwMgdJFLJI2UaO8lXE7QGR+Af+Yqxtjerzj9
fpXLh2kunmZWVdHoWiLmkiZlISRh3X79Kkrzf3BZCosB0PBgEBPI1ZLBOZtKIYGh
PbrVKfH/L5HT2u1gywQvwE3w4XvKkr1nquSRxHL68RyED1Gc3ndn5atIbMvNeVbT
kjBPlrweEAzmnx4iJuhWWMBGdg1L5RaidBNFf5KnBXpvws4W3eQsCdDYwQTQxU12
J4z0i8YSR3wKxiAI96OOxh2eSeZu7Uu1YMSO8P9gjp1WCCqPETlo6W1jkzkeiw4R
SSEZVftZ1jdQm+mv/S7M0IW6eQgAQNQO6xbl50uHJSW2Um8umNA0PcYKObqIHRBY
jyr5x19xZCycqyRtxR+bdSCRFXFDsMhhHYdkwGytfSohw3nQ97buyjBkTgHN8i9K
4NgZceRusCFbpjWxk/dhnKOplPth5TdsQq3OIHXbvnXKG/3Krs9nvmyn/AxnfB39
VNLTm97upUcFC3abaTuFPipQcTPgNZ5Bg5deIOXefY0xVJAvNp08UmWbQJICix8N
Q1dQB8tcG4wQxNlTMofggrdeUiLb8TslbmITZHHnJTTQMwJQT0CVr4PFE30aPGG9
e4+tYfkzn2hVSgi+c+zWqX4kWRwi3Di+Kkv4f0Kg6wU6D+KzpuT7RqPpKx2u0MX8
t1d+AIgOR2mPR8cYMxciPDV1u6TAsK2F4uMgQRPpj4C/x8Rr6GnSrTbwYb+8lnIq
JxouekeGlc+0pDgWgiYl3DMELtw/O5qUHLCYp95DTJjcVBWj18M1Nk/3nyz63ktz
jpE3x/J0KNtVA6GlwIN37FGDynlnP1/asTVmGAVf+uRO2ClOzOHom9EnTQ0zxT1W
PQGg0jxyf8Z0JNIpu8OHZzTULqxRN3NAT43SVp5DGsnAMfRDy2TwSUCF+84to6te
AYv/aT6LryTn5IDLqJngRExCtFdr8uP7SUFbezhaF1QqeiTzuMLCUAwzaD4R82LK
B4r7AixAVd3mpGt3mukzNIVcou8v8pk0jS7Ojzmgq8POOmKpoX329KqQo3mwZvR6
Fbk6HFPbQeAta1C2nPkLlDKnq0nsbBlWiSWcGgS83CX9bn6czQ3XCPFA7t3fZ0KW
IDQXBYDBfhmyt5LTdK+4dBBgtFPQVNmaKOCXOGbO4F5WQVEsmpKRAHMDEGFFk1oa
9GKe+2KPm8X+Vb6EqzTrPmaih0jc8Ca87otJ9L+QV++5pmQatbHViH/b7UYNsF0L
azy5HB5AE7ncve/wJo+1scoYxemaTYQGXzUUGoqxbHs+G4sjHDiNJ7XiYnciXZEB
80lRIbTarDFA8+/uxLFb5VokswhbhGN8ClQwlgRTLnXOPEgUXBP2xHbEH5rlp1OH
3GR60k35Y5a0VnnGywIko7mpPMXnF0XIVI+aKc8f4TNzizHSaj5Nzt9l4g7hw7+L
fftNId5hq9QpzgGEGaSE/9Sq8SM9bRbBEcM+mld4ThFtYDXBr4EUV2DpcgdoUgz0
6Thq5cOlHUzY8BN1i+rmJnWssBmH9kuq6t/SgEO8cKpEPHO3CoIaoWSQv+esTOcW
5C89ZS1uMYlHHMCqkVx5ykgLJ3TUdno3rew8OY/xSoGCuo1N+af5Hfqf7hd/JU2g
ETCCBN4F0W3f0iUuFHr70tGYBxqIhnuXFwK36NAb9OIBgXwcfvWCgAT0OOzoRdki
0buYVKcsgnUFkLTBoiJFQLJKYlQhLp1KoTCUc9qureGrhYoxjKrhs3GmsLnn/4cU
0BG9cTyYXj5IshMW9AeS3iWShlExM8TwdPxAx0eyNWvSIZXdjmj+W1nveAEiQFHD
7i9QEYt+CB/lgBkMIZglvVJWcu1pY34g7cqphdwc5sTG6BQLg72ssSjuJ0ZzCB0s
IBcGZjKGAu4OC7GUoCdg/HoOBa1b1OYpp95qFRFApaE0Ei8yO580x6rFhj+YYmft
fVjZvLpj+oASz65aaP75pz+0eVf4GkR/F41Bx7AGQYc7ZN8ckKjPEqp5UGHtBai2
T2e4RLVzO99OrHLG5g5zhgXLUO/Ti4RTKeyfMpTzK3nZYLZXpEcxWPSutGkxsRzW
+jw0f6cIRV+YQZ+E93wxuRRlnQAbKw/YXfoGoLy3/FwuR2Qbnrip+AhbHmUIEPO2
Nk8cC8LXx1Ph4kM270vWgJDO5Wi6VMvNblYDt+0jYOqjBHlUZG6EcnT8sPaCHZyI
vVZ64fm9ctlymKAD9+mxkMkimnbQ3VLimwctVIXEkraBdN3j5Xwj9+iTnIdj5i6Q
bj4npQmHn/4g4YOlisMotQgp0OzLLY4fqYlU8iFcIDoR4eRpwI+VxzYWFLOvYqg8
OBHONdaBdSh858vqBjXQGhiFix7yvXAtYb6hjodrjjB654C8lNHDZ94KJ58yhhs0
gJLuBv66xPKN+SJd9K4AvKETHvon88DQ2juH5sxCYGyek+OJGE+bBKY1Td0H0uhO
IbrV218KUhILGnr3qyD1HlJocpKTXuj+qrrQzucYC25nprws9pqDyfADhIRhnX0H
zUqBE2vEJOlZ0JIiLVwu2R+SotW0PkvNcWUo9eXf2NXPRrakSGTnqu6ci5Et35D+
fPpX5Z5Tkvb+4BkCh1rAcOkNrZi3pQyMnB6f3Qv7eAHTmbwSKb9xBciyRaghW7Ar
rBE74lGm7hh7IsGfqc7LIUbBuklmrBXMC+OsqVu5G1U8ul8ZqXCCavfZntrHJFEU
AyJDjDHGbqVerQG7PUMA86lKF9x/xDAsWapvz0MZBEPPotdfWk+r7/rVeY2F53uT
6R+NRMs2/4+7wM/vZEoGZYXBmrahgoGwzdunUEFTMePofv4CzfV9j3FmuEDl5ynT
hRrK/6/irRAKKBRGbN50ZTZeo2w/PfXfBkNZqhRlSEifL2YmR6CXXDWCXVJWkYmi
k1lg8F/yRmps9Ff+7aKIOvjduzxqMMhnV2WmfE0jLFKvyGs7G/Pps4z4mhEh/yUf
Njv/2gDSFVrTY0U7qLuHkRhpn03U+NjFyDy0pfwyCICPTznpCuNi9s4zCBlrNiLY
Krk7KsfFgyoe6n8Pzr2tbYYW/Fr/LaQSuW0WHlOyx8DmrKp7o1DsnGTklGN4GP6P
TcvS35je05JtxrFBfkIhBcdf5zdK5RdCx4hAICTym6AyZeSSoOe65qW3Wx3WLK5P
8507/pN0hwzzLU9sxSVbBWE7Y0C6i9RtD5TzS/7CNSA4vlEcPSZLVjEJQAumch5C
Z9BUWgn393E8to5YBdhBf2NkKO1h4ywAFwztsRmOnkTcQFODttS1PhqlkN3ZAj7c
n8vFenw3hcxc1GGiu36cuU22Lz4xlB5lR8RBqy4uM893rNNrkaAkmhz2bQaMQ/ew
jv1mHt1H7k1mEfvB1CrpWxltpn3F0/9UE6NozH3uZcuVE4Mm2bEP/VmiIOZUWuWm
rIZWs9t/m7BHBxeHbVV61NxDKuLR7f8TLDawfeqJuR9nI4xsWOzqp3I/eKSljzIb
ze8rS4kUncHFysqoX/CszwyCZhOv5q8lGhhR3L947leJjaYKB0/opPwed8hyKFgo
XMmRz9QV+0+LqpCtV9u5Rle3lMowxEwo8Z3+up0iH7e3r8tTQiGQ/RJ8hnUaQ+pc
5m3uZ8YClZCkAaSoPMAYOpyuK4l9k7nxmwaar1uXqD/kj/bLqqpS7qFGAJb4HJEi
yxxKXcV4ORsEZKeMDxkXvUoSpj4K5JcxtVB5u+3upyTP+y+e3/85m7PL1Baw2C3W
1Nu/EyV9g0LV5PZwZw90SNcE9IbkANgzxJrSSkSwO9QM+7HesIzwnYV6G1rsJMgc
8h5HNW0w8VN3rmsJqv6v1Er2NrIm3Wd/FmgTlWuLwvSWiRXVIJIhVGSZh7ULYohS
/qmHJECuMCvhcEaK8mH7kEKu6tH4DwBX2PWCfTO4mL1qoscq8wSn6gJW6YTXbBOm
XTZODHxOynGVNBAQsJeBADkA2lJTmC4hXPTNyYWDrVXNnm++r/WBwf/kNhTkF5Ac
ms+GW2zl0Lhq6x/2XjsWqh51Wi+/7Ip0/g0279Y3YBtGZ6QN4R+rL9dmpiyxeZXk
1rCHHLeR6k5JrpQkBfXdoMiFEw5uk09lQa8BZimmhqtnPsAu6c1JXDeSJmFPLX7o
BCo33ywfCkgBeE6zaBzv2co0/HtQnlyL/t7z9q7zg68noQRsSiy3i7UKoB9DrIwF
dLzMEFcJP2boS4HF6tjogYSccwh7JOjlPh+A2VdRnC3Mvw8HQemxzC+f+d7c8AHh
claXVScZZkyC6jYNEN/Lv6lbDjA15tqyUunRTzmxqqQr4UQLGM4tvkf3HpfnyCPX
JweHUklgxN0V+eW+Bo9r6xiM/2G9Ly4nKva42tWSyYymeAV+ONhI7ll9fTGkq6JN
sUwI3im3f1GxJeGrYZLDD2Zdq+HyQAgi/Q0jIiVa9nlpovI8oGECi9Aqdi8rWzW3
LP55VFBMw3k1y1i1QSynBUOS9qn2Lg2mYQTuFtSsDNYFKdR3wAwN1MmszLhXC+xy
S7q0+7d+A18MJkbA6lzoKyxw83h3O/vEJj0v+tbzwRPO6m5le+xRHhIQh9uGv8lu
JkurrDRKAg/TvphiyUPKaPNlMmQlnQzCdG8pTBhfZncQNMxVO4WGTBmoY6AysmQ2
45yHwP62jtgCSQD8Opk4rbdr+628tKyQJj35eeWa7pR2ymFu/upy7vZhFeBtT7Zx
d/PkzISINmXzbU1GP53iWmOqzqie7yvv86J3dI+UvQnfSdVOBRSZLUY+h4OQwGQm
HPoqO3iqfdEkDMJ9eyrray37LVRafMKPz691fNYBCOC3Tx1i++eCaD3AWBOwuwoF
Uj1SRMeOK0ubsu/oiwo89OqsbFG2mabYjEm1u2vC3pjC0LqKWCYCcRCCNxWcDnt3
rLxwdMj7DZjaSWgjPM2aKipIeFjJJLJRkHZW1ejTOashft9H8zWdn3eugNg7Wt6A
s9Qtk9ETxU/TKuXqCvJ33iL3uo7Cv/M9NySB/tUkTFr7f/k13weiENdrh+BBOrI5
gHkCFtQo4/emRfYTV2RLk+LsJI4B5a91RA5TZuJZ5IOcc0C6ASf7g09m7UUCWT/B
nMO1GuI7wDkOkBcD3nbIVKWxtFoJJllEezTO8vNUbdWvbh2W4rieSYJ2jJHuZH8n
KOBnYSnZvb2f2pJU/weCQWlovV3/o1QC0p7Nu861SgLH0+KmawK6aNfGHIbBr6W4
Q4pjDXf/zpgfEBwGBkGPvgpmUWHgkjYIZN1CLvizrvyjhlLejHdrxjUTyH1E+aS3
KTvWcIl5pw2VVOC6h+GgQwskRN19rFr63I2aj9h69uqCLkGUaPmrR6/PwxdRD5wN
ritmwq8iv9hhov2sRLyORHFVhhXIak/25l5b2qD1KRjuoXt1+jG9dGPI+o8kVGul
yO4mg6dWOaUt7KSnoNtONghDaSKmXLrE6jlr63KvrLkfPcpaD/gJaXQAb7PKI4F4
aMAAgxfxhFYUDa8SnlxfcMkT1v6EW0LpJVLPMGnlY2+SCNrXrQC9MBhtIFof8B7q
ck5tFA0jtL773WGRMFkR/e0Jndl9Jvt4SZPR5gp+UpPUWZUxjL9/kCn/DE8twdj1
vg6KbKc6qIoiv736mMowCT4hT2VbjKVdgNaaqqfiMvdv+vJxfDebXnDVYjekbk1I
CPzfGYwknMpjlcLfz11Mq57eMCLxN3Zu45QMJEzQq79yN9fHPvLR+no+K9V8x5Mh
Hhx0HSsGG5wwe20xaSTyPqlmGXtZ3yizPqCxqExmrbThG5hboFEoL1xlyJxo3c4q
5yxRbP73MZdpAl4kNqMEnQzJpEF/04FmNy0INBLypWh9BGyU7j6PnteKKgjjyDur
yFCj8qfFJVCJKW4ZzAQePp9spSq5k8mRoDNx1voZmFIHwp0cRGcSidKJGb3ebqHq
Dr9MCtGiBeJ02HWBJSm677uCK1AiB4DTy0CaY+CRQEw1WP8xT7kaaffplDhoFY5Y
5RxXYKXqu59ucxpj5LGmjBLAnpGZ9sIkMkLaG/M+jIVDT13s60LG6Sh6IQZwExeq
3efqAd9CDBHttHkXgbx9Grq0W4yQEICbgGGW10bTaJHQDYWLUt17D7elxEoTlOZU
l7FXUXYiLtFXU+3BqbR3eW01TM9H943kCGa248KykPgBrfNahJ+c7bPmIvSG+QRQ
cAS0nAS31L869pEWe6XYiSFBnb21lWS+UJmvHmvnmGLDbp/OrYNVinbD+4avJkYn
ez0GKcakEhmTKd6HYn+3RueYS27MEa2ro/BwhzUXNx5t9AHjoPxDA5bdq8MUb8WH
iFubf2hNx1HXWtTixCDiVd38VAFGaugu5zLuL2+jffSt1du0QOnc4BN33urnVgOi
4emMmxdsma4dp3SkQ/OfprK45VyeY9f/v95pPqH+OI02A/L6UBB9pBgvvk9ZSszc
xGgR8DAImFkwWYF+NfMMVYvrt7xv5FgleG8Aeq8tN3DNxZkJVoHYfdLNDQ7donCC
Jr4qfcmMawUgv3mX9AfOgIM9Rq+WlD9a29FDIpRXb51gLybqUusqvGwNHOkDUw5F
Fz8VJa4UixibvAXbbA9U2xXxxmbMAIFRgwY5YX1+68l4qMx/jD3vQz39eGn1UnOx
sJjaMzk4egKgKGwFyEwi5s3j0CzgeTtQhSoq0bVQaSk2AHbqx2krqDAGbSN8QeWd
i2M2UbkAnurBbzEbZC+hXo5c6xSlCzeW0HMnrIn5kCULbJZgf62erSMX2JyO/e8u
4tbmA1SjTb0aELV6VyDdmr8RUFVKe1HFcN58+zvyK1ogZg/PWf/aGrvECqAnfxCL
Tqv2oD6rznThvfJuleIQpkKPupCeSI8EQ+tekztqhNQ/he4roHbHe5yT5lvrFN+R
EOnhJiIv81FbziVgdZsNTXMdRC3y9s5RtUzEeQAFuqyHgaKFM7TDUUpynPvjS1gX
I7ouXVWnYLHIsn/z+MzNjQzMPSyO1AR8LQdbtSeK652M/6pn3f8iSNSZVGAvTyMI
AQv0Fhce7IoJUcjSBy5+OvAwe3AZnyVJ22rV4N4cFzzTBoG7QyPbxSlg3VwXYGr6
c3dI5gxaA/msN6WWr+dzjxCYZ2sdTgGyYUoqhLvY5HHG+tvq6UCxflSWwVLsABDQ
lam0V8QxvGKMOjMXj7/QmOZDax0cTZuYBaYluLY6fHR5rPPTCQ0w2P+v557umgSc
aZ9J4LiuleqiKgcIJCUUJTt4JBoyOzsM99JuM8bAI951EZndeZKFv8lG1R4D0eEN
IKIz5+xrfD7BRHwS3szG39knPUMkRA/f6kHoRgZVVA5KfUMtzH02SYeLaL59ugTh
H5h9uWQKVyNCELLwD85oPxvkvyiSRPnyV2p3xmlsKonfFYc5M9AooyAx8L9jSHKa
0FLfomwi+dcpok9CXiUlVlPhUxyJjYoqj2dQ+9Owbs40sAff6B0WI9nSuMYsdAUI
adaWN1Pc2V+x4YPWtGxc1DbSQh/qA+12zXi6kjdz7hqaYUNfygok71GSSpQUKKN2
m6pKI0hCSxFB9KKpNOVVK/CkMnmgOhEoMS3er+VsbrX8zqqIXLRJn4LFOMFZWWqc
WoTu9Qk/yZa9oSsARuCG472P3PGKIbyKwztxg0Jy2mpdJC7m5yfyz0xltC4Dh5y5
wZrru2/k/TEkZ/ezp0kH8HtM5ZpEzuSwOiG5+7uqJdmabmUClVXiMso21nR4gN9l
9C4SJYHfp1A7osd0GdB2Riphm6wtoqHN5tWDoBsULfjSkb7g3fuRx+poIA1/FWR/
r/vWc7/u0yqknCUz4DVA3cNc7KR5c3DAllZmD/8039HClUBuBK94NbF8SjcYFgRN
n3G/VYkOwxZu22JS2DX0iBU1yxFAKZ8bAKoERqSJrKIUmMyjyfONwSiZd3QaDvtF
elL6npzsoykrflrWzKPMmBt5At88WIobyvH+FlLfIZshpsk3kuMJk6C6BKgAXFhm
vLdt8Xvb/8et8WCueI17tCdQq8YVjer2546xp0lKavqjCn8w3DSeJ9r67MrLwVrx
a7RiGBjJcH5LC5eDSWQEpkqlH4lzjxksvXBA2mdo7l12wXHqqxsld1cw4kjjWpxz
dVZ4rm37BEYiHQMlEsDARHEvbXy2ysHvTL8kiPlrDwMJOKj+T+Qp6MQ0gOVOS0Nz
YFcVqY5s1t03C/wXgPOAEzVj4l8FwvMP0kQiwk94+xKmBXJ9O1+dtfj/RdPTBKKw
MFocZ9APnsHRstNtfAoJ/OfKXuHJJJmWxsNTVH9cnoI1K6u0HRpupjdUKylKh62/
i58vxhTkQ4721vWdc/ZkwNKww/v4p1pPW0eCb7V7WE0dQog9yo6iytgZXMc7buIY
XiQ4agzBQmbjVNJb5Fv0CcFPFauSrkzIdSl1TeXqANS5zN+owtQwxliilt9ldrTN
7jjVgZy0C5Cp5GAuRyRnQe1mf4hDsB28b5nhJqqTgD77f4mY/M8HVwapRsOyPijZ
9c/Q3VoTIOClATSuzltDELRZY1LxrPAhKmdqtdlE0hnK7iXuyrLT4PpSMT3X6aIG
dIH9HdRnEjGkNQHNaCtWbVjITNP5MAkU5BrS4HwIaFgBMxqgCbOV6NnccyHn6vnK
Pers6GrP5BI5rUNFFZBJMg+byA7eKvAXG5yF7FOs7cJKFCY4osRsHzychKIRjY3a
XFtVII5qsyflwdGKhdGNMhJoWpNDNiSVbV6GQeUVBo+tRxGEBaSc8CiaSj2bwRog
uZ+C9IcGbvI+z64wz76qXPbuvx3O6tApcjSqdKXPnP6Lc3tLAjmsQbedWRLWKbqG
yFrmCrHQoQ9WGzEBalw6fkXvlh1m+0PMmZjhBEV5R4AKOkqJsbtoYEKhvRsbUu1b
+V4vvGHV3XulE4N5jBt6KIVG3vK16SwJAiOSjaPYMfizzrsFZKK7PVxaGI5kJYe9
ZLlrKnQpkWEazzKpFv2CsupM6dLUW2diTWaP+6ofTTWDaDKwxtOy//pNuEfBCyvR
XfORVgoHwLcUhzfeRh/80ooYQs6S2gwkVRzetAXW+30Y2U9WidojNWmOiuPhVHup
FLlWRwz4buY4pUJc8yuUJplWYr5V+xWU6ePaTmxRABHa26ZxfXAJoZsjp1uhYDc6
KVSx/0bpBcRrMfoE8hKO29fvbo4pEdjvOZoQXaPXdHb89mrbO6fJMb2hYelfc/hw
0E4gNsfPNLki37OfB13BeYSyWScDrkT39iRXYpueMEmiCAYu2mgADjU2WOvZ3noq
6TRPpL/bfoavgwbBtKhqGqzh4TQF6PqHkSrGyzdB/s0ki5H/CDuid55XeZ228o4L
72cchPMvpkVcRDg42zPcyROxypxJXGtBaAlqoJiwlVPHz3VpE+UgmzUp3TdzoeSL
LOO56bvVnpFF/d2/IaXXowtskctYu375f8VrRGthYcbePOa+1l4zUZEMS4wtSy2G
5AwD1XWZxMYe+w9xVZdrsmZHR5lT1oHndrYdMcKnZAa0Ikt6V5i3g5ZV4TPrwSFI
TZGclr6tRdm98UDKv0gz6t89/iSZP6ZaSvCyAXaCLcozplJAe9W4XKNpL3IX9m2/
YjZnFhzz6MorLXIo0Noq4CvfHM0ATcWIGGBEfjr2UgKG8rbKiWgmX/pf04N1Nk2K
agpPgusaNtpppklXIjGzLU6/HE86L4BcuyCYO9n0vuAx38pxM1m5NJ1+nrqvhwlh
ejj3noLwC+YxFvT4jT5UQsP4pb37xKvYKsaxSqQKYFb7+WeNa9FER0lDC0Ci4hMx
ZKEYkvkETQEKDPmN2dmdgLDT1pHtNzlWscnvalg0c4/iQrqtBC4VDf02flNOUVlu
JVQVS3ZPwJ3MzVQAXDvheybWOxwunepJHTbgwwGh0HQagkg5+cGZhKGNMDqXaxSD
cdfNzKL5a43HSZJD+l59nEXF7J5AdSNH1+7sPnZU2kySHCRamp6Gp+zU1XS19OBv
l/vYO6WI3zvIHgFeA5VB9eUnXb6aKV0wXKxSFLtuBIHnePNYyB5Npk6S8Yk4MwQo
rT7oTOHVAVTOedYXE6e6Fs2beR6tPe0paVV838MLEBotAbw+UPyOx0CU9l41m0kH
cs+OpqDVAvTHNoC2p6mH0+TdN4xTgzOd7nehuBJ56tN+gQeIg+t2qIPzvzWTpYBs
DP35Zae/bORiglKu32HpiViMieclr17hTVKXkKJKzgt1VZBc6cBkYWcNpFgM1AZY
cIq5ps7SVyjzGN/Y3fE6Ucz53ZDAWgcZCK0tz/RjUSk/4a0MtcDOTfNqPIiw0oYJ
lumTilQ+TgXImBRBUmirKMsBxG/CLxLkIZaA9z/58eABwe0K2rdwpn3Qnjw2T3Pf
qI8TvrrT7PO9otURIDTtHT0dKluoIqxCIjxWBg+nM0g+lusQ/+L3J/3Tin2i+BtC
20v3PGpJZBTEBK9tWENE4GCNK38szK3HhhndXUNRg7upVmWPjhPNx9C3Wt1KNzMR
UmMdNEZPmCgSKY0MxO3gDu//8GwhXRTNI81rU5IOy9xCrO1gToIp/Bo+RGI4tr7I
o3tge8JT21C7J9isq2qInGVJMRSwS6FxLM0D9o3EJFzuEhS2BVvJP3WHPFD5L/58
mXfbZzuT4+BbiEeTM8dsluY0XdN/LtFjkBv3MG7LZkO+kDiwFkcjJ2Bydnu36KpY
4bT/BrDSvhByKOuTUui+5n5yH7new8PLgcvuo7rOnDMhW6TdmaBag8RWJanOXJXu
SnlmLoJ6EatNzAqlN/pDalEAUJQhHG7OQc8Y6ZPxeLHiQHfyUHaKA8cZOQTMg9HB
pcyl+yN1EmLoPmOWqV9Nh7RKGB+6VZMNzj4RgoQhmZCZrujU8uHtnjldTmA/9XaX
qh/YOHJZ67UudSfKiTNM6OIO3/pBzU4bjEGXMTqYpQEEIziSKim1brPcIdddEZk0
nhT1RXGuqmx9oaunyMpLH3Sr50AH5D0hC1XBqMdYjM/3DvT0ZZOe7DbX92bsuQR+
EYFSgCQHbecFsVDqVXs5/Id8g6RNHOkdj0zz+NnveTsc+RCR0NYx30wLdNkW7bX0
WQd0ORdQ7zHtMzmaJDb9MxA+yKMW5L1VV/a15OeIqP1LUIMsz14Uu7y1wglq3QiM
nRFzmTcRQgN1Y2GBLEG4nc+7goV0TbeBNOITz8Tp4zv+QvHYRP+sNL2uWtLWKPpF
Cz1KLSekgL1g+irUNfpfohzwtyot0q0VX25M8+jOaPED6h887SNysncyaUlsoAAo
vJIkhs4AoITeJU3ZL+HYLqPq17p1zGYVJsTUBeJ03J7jBbiwwK83kBbwmeuqY2VH
vkZDI4QXFV+zIue5iXXBwS/rmHsesfkkWTYJyQ9EIjRkFBlWsMYcPaGjylKoEhCv
1KRm0TR4QtSzx0TldTI/JXA7na1f3J3ZyodR3b6rOTqfYEkwgzLoLONdBI2DPq/m
vXiVEhhvimFLtM6Is9y68roU8imZVGAnBLy1RUJX93+DScnEGlWldGi5NToubpGD
f6wM3M2yPEGOd7yhfn7780+1sZn9nVAvi0lqzFjlrPpcOY4VIFEqcWg9MijXvi7r
iSJCGADzP7iKA8cxM6mz9lIGfyQDvA3Uz7n7p6UEv3gkKLSEDznR9jmtiG+yt3/w
ccgDmIRaOar1flMdDiEFgqg6gAtbLW2vVpfRayZdGQ7rFAKpO3ZxrhDyaQKVJXtn
8lsmL3G12csd4YIJdHyzjF03Uo184ZfSXFoEb237hw5Y1Z4GuwBjN58fIcdkzbD4
NylWHr6iQyq3JKot7bXiA+qBnnn5wKbW+kKnyN51bvRtosnoxOF+cwaNuGg5J0RJ
0WhP/K0ljX6bPRrv5eUqL3YU9HhOvd+K63yCQvR2JoNRFLf89ZjYqlqH1jmarV2a
leaZFLMVilri8LtJGGbL/WfOFMag9+q3sylfAQe5RzSVGVKMdMmXfCfdN7hqD54u
X6ntMc8kfelVEjedrOcp/+KWkhdUsa6YLF2NqCN8pjzbrPheafCKs8PHKNotgBbt
PflfjkdxYSY9oU0exkkOLlHfrFeMHoC+gPjdQn5MPbM5JdyZrQQ3xi7BMZiG8IiD
LK8Ijy7ZTWHxNtE6sjExz2/gR1ewnMK4mKFGeFa6NS1cRqJhGd8f6NV3IAQpnNiE
S/UuVe+ucCxZXN3btadEQG9DgmtKGtjeMqvSFRn25Xxb8sIkxwlZdgG9YU9QlCjB
0uz2Ek2B0d6hJVkljhIrf2DdJ7/8A5iYhVwEUtTiH8S1KMubUsEj98BokDhtLnsn
/TjqhFOpaW39o2zLhS3zjW+am4hF4iERpNFaa4xKRItMFB+rPxQ70/Z09F7l2Vlk
NGGqTrAZVBXe+AE3GsCkZnFn8A0oow9IM8eYu0+LB1vRpH+8C2+l988ND5KCfpEe
9infljytcFcTFsS9Svcii5NCHJMnsWtCkiu74wzSPM+uYcqRiPmqmrfHz4pPc2VG
05sbNdb84WUvpI7/dbUT+MGq216NGesWctzw0P61u9PI/ZlUPbOKAs7VO7tHuzfs
Jg3YoHOVmtBoFRnKOZCqBacsdvPmrP+fP86vwCjXfrH1cImOQqv96I7HaVWmMczw
jhbeGbZRjwwKw3Xi1XqMki/1L2SR8IC40JIZ11pTSszk/IS44Yy9oyYM/JTpsUfn
20/vDQJpi3Y3G5Xb2Vwf6CW9s5B9xuMvgkhejEjWfTVaCAKt1KOidGtwMCE8AlR8
wjHZypiQMtCAt7cmkqJyz0zguoTDC7HiT4qQ7Un1FNnpYSPVm8mCnzHokDeOJwrG
IQpaPsz15NkD6rBpi+Uxq/6AsmtOmmrguD1khDbKE+3nykM8Lfwc5wk2jMWp9hKf
jSDMNTpfDpZpQ6araYaaEuNc2ddyBYUP5D2Wl1BgpAqlw2I4stUga114O/RaFmzb
KCViX+/6XjD9EvYBPYqgIArNyrmgSogsY03bvvPIDXYtFqYTy0/1O2FJWxtA0KN7
HgPqpGFbv/KG0rmrbegI3lokwEXXmx2mpumCF06vg87RAr6uEroAJSUcpnL8xySt
VFF6YrXuCHIoChA9tdP96EbIkm6gA223ahUwlTvJZjky2AJIfZv0wt/giRz6K1H/
KOaQd8N+LpcZiDK/J2W3IHswoJJT/1ZciiF0Rd5+i3tfsadsVHOUg15SqME9pvgj
epxW1Nnv5Ws8S/LIq1I/8dSxl3lmuigB7AaO0/YrpNscbrMxLnsg6zkPBTUrcHI1
7in2iIvFERtnQvbIeUrfk27XNAou3y73qIkGUBY/3TrUmz5NlZxrtpy1ks8bqMKz
zxj9HYBqEfrK+I9eSBzJV+rh47cdmV8GE72O3SAOyoH/Y3MeI2Y8a4uxXoWP1plb
DqTdvEtAJkqSX2yMsmiCZs6pw0h/6f0zarvD8ForY9nKyVubXoHV+GQ89i0uNtg1
S7YSb+PvaFiTVYSRxVB+CUeYbLfTJq1wdaEkyczipVN/bZ2XR4DmOpU8gghUo+Fs
HXjTSCh9PQc+kge3v65LzHFRNkAe/Q5HeMEER+JNNgPzH4CwnmDO5dBNJun/3yFj
FO0yDmIPbR//Gp+kMSc32nVNygtiITON97JoNc2ebFCB6fsEMv1tqlu/3o88YAlr
qGxltzW9SnmNYjFo81VYbxntjBi0VM6HorOfC0mrzdsxpw5DUehm+ijX/N0z5iKE
iZ9nU2YBTmQc5hMA/58fHbd1EPbAexmv4wkd5IsZPs+k6CkTnEAJxPkLKYJP4gJD
duYZiHLLi5giTW+DwTBi7XsgjDCGeFYCrRciQwllYGwUVivaXqZQs8Suu6fkd9PT
I/8LPUmCT9Rl40hZrly+VAj5WECRI/nFyoCqqdoOU0m3WVoumA1OgdV4aorUPNjz
3F+WFYzf9POmsdg/yt7iOgR26gFWvSwq3a2OERYWJ6tiLN5/vmZQ4vD+AmfuI0EE
Qn5koHM3LU1tDCbrLDaZDCrqcXSWO8T10BCAxBBeoc2brcXVnHRkALvB56q7Ax+5
2sXJbb0to99228C/6jPCrq6irOtAS+96X8PfUp4wkxCPzK4pjWIZ8QPzPHFieVUw
d14HQC96DxoIPnTvJy41t1h7UppbTBDh78YY4FlWQPXcr70z+jrd14eDkQZYB89r
VJ2Fuuzs32RiB7ka8T3ZslIFGsjk7SSEO8rAL+ukO8xi1nPl/76zEADOwix8068k
+lAuMiEdN4weXDjr3UQgmwEqgTrNVk3F2xrAMuRb74U26JPqjMrZ49a8bAj27lJ8
q4By3AKP+dCoyWFQ2U2e6c2rXB/WmrEz9fJnZ+Dw5wC3keq8v7jylzaxd4MoIGZT
OeLpVvFYtvTudkGKvzZ2zXrbcV6ue1YnaZ0Sev3u8iXtePR6J4MGdee4ZvvAIIFk
ZKGTtySxgHF+CwKJbCBhNnwPnRRrSDGgpM19F9xjBZwK3XDiL7S9erfv/zgBM7JO
en5Y/ynJzSudnQlB4GFa919px/Icb4eQXdhvRbo13jwNY8paCFWXbGfJ1vgz2OcQ
H3CKcveie1ezVNtJwFMfnZ8vl729iSxEeNl6YsnvlkKCqSsR27KQpkGSrRwkn+AD
73Vk5jtiuYyArDYVIPDFk3JVONC2TPZPCxau9Hh4++L1PU5wKNxC/4OvL6YriNaV
SUzHEKF4Bp6MxhORqPVR3QTu1r5e38c/WnopPugEsyhKavaZMNV4RORkoRdromHC
Vt7WMO3nE6KNaeL8Qca11fOYIG8o1QgZVnpfQbJkeTSpShTBOu6b4d7bkpyvtcBV
qoX90yfvMRzfqLkDkfqcEBxiZrKQLFoF9G0k8VwJgnE8325yajyUBEgb6V2/A/yO
aSdUcgAIBG95k01RzRBfWASLnmLO45jSHyZqaBt2Jm7VIQRQkfoEk32+h698bpRi
uo8m1o/Skn06XZ1j12aep6q4a/wUZB+j3DIq7N9MCWq8stteOszWuLT8QeS33rXZ
1NINyeo0Gdz5hag2KVUy84DMzIx+jPQuyJ6JwHFpBVx2ZjO55KbVLd/WsoYoDowy
sHc6DO+otgxYHrj4D4BhtmSr2JK0jMvmfElcUIfqQa2RgpHCdR78Ww3xrRVN054E
60Wft1AzC5dOF07s/Jbrm1ov6lh76avaM262m5oO7x0gKQk47iZ6BQVQ0eliQTmn
eYwPmD7TLkCmD/9upVEw/iPOTYIyb5x8cTBB2kbnKzh4JvTAGyy/yWT3odJ8KklM
p2xRE+GfaQ1NbSO/IqmJkM9psTiIwJkUJVgMCsIXQ4ZYveaaFW9rBVtGAbrDN8CX
oZ2wgxf6T5cqkRmvuBhX3WvODXYoSf5zXtgr4hX1TFpvZ/Tg2ivAxz9gNsSVi5n1
cSiELvbTm7h/XkGDrFPVxuaV80sMzRH9esDb3+NfekHJpUX4/CgZr0g7YKM2xbrE
kLRWeQwLZRvQGgn+nK6qxmK2F6EUGuRPafm7IeSxIwsZYJ9s7CVzO67UD4lSSNEC
W+8fVMDLGhUriPnj1LiM2yCHegjK24mnzeORX11d0U9o8u+aLS0vWYC1MEHFJEUH
9p/OPwwDwGQPfm76ZoFEZ4XMpSrZ4EifHTvtDsOx1x1T4OjlJSCensAlmGgUW0V1
RM1uPlcxqwig00wy8t4Z1j6Htsm5VlvyMFQq0Z4vMfS92gqfFIq8lEwnDp1dDU6R
yqkocLEeFjh22xRhn1xnJ/k4yCTvFyIOnvTxCkkRBJ44+XnS9oDBu9y82JiCcYQw
HkYo+FhRLl/WnfmxU1jOF6aAm7yNJsonTrXPPPxCwOU2UWQ5WbHGYCC1l6Nj7Ux5
DgPGPP+AAojjlxBbOjx6e/AbB5+p1AgM+713PfTDovVokHe0TjhF5jNtO6sexcgM
bE2+W+aw4e7gSoZp9EKtTZ1PvEDvN2MYgEKhUoZSS7j20bK7xLCIHFczdSHIFjy1
Nqaq/bkueJsLk8S7c5CKjb6xkpaZo5OkLXevo9D7Rb6YSt29/bdnAXI2BwzPxpHq
SPx1Nvn3e80Rm0G7akK9xUZQkU2Fv38cQX+A+fEIzonyb+fT00kCeJEWjAsEzBEB
miUP2cDvdI/0vuyR3zj2sDOJ4t4BTmkJ+1xoJes1O14wzhixc+feOaKmw2d+xw0g
4WR/r0cPgaO17k7dGgv1RFLrLNqGfLbhF9HBQIJtd4M/itTR9YjJnxk/UTrci7HG
zt2cOZu7biDiwqTuFwQqA3oeIOgtE7Z9F0FbrJ4SN5XUxbZ3F2e50XQ1BcfVaUQ7
PGx1cvGfC7doOyI4YotqC3J7APKxyZDvbNcscLtUZAs6M3QdvRO9wFedmTarUySM
Eg+9Ti/bThmMg/yjm/604PYXPCugde3a1RDt9r+40wkg+G5IZc1x9QDi8Ho0T0Op
xIOOT+6iPsJVVLlx9UeXEDojaVFdg5E9x34y4ZXsalaNyTGNIa9x4WxYmhGvSXVK
0fzT6lM67E6QnSzjTrUl8GjS9A+W3G73d/1uAbq7FGXdkeb5ve7KBAnsTsLKVz7Q
1TLKDjXBFYHMkt8wAqHfVdDYlvHB1+J9oqz727iGKxEKq6dDIk1Y9WgkDOKoBnp+
5ufK7ofNc0Hmm+DPzIjaSrVM/SrgjWVSyZFWwIeuuH+Hpu8GK+Y0G9M1tFu3miiu
Vmi5Y/J44gWPF+VuIwieqeId+aMBT5kqsVTvuVsQ5f8oVbKEkW7MSwwHP7vkx2SP
IWcgZiOwfxCVlk4fw5NY0yzy2wCkUQTKY58RkzTv5FEKsYTsbIBTp6wRQTGA+c/h
nUzvXJaagwiXfldO+Bkz3sXCssKLLS0WdzMgozlo4SnCtX6f8phO6gQhmt0ISxeV
SqTt0Di7h2J9wRjzLXJai/rRfLV09v3YaFFDSyUM+74ePmppZJFsbyu6UboU6g2e
5qOvmKud5N65MC2t5FaQTOyTngCrS5abzZgafe2Eva2sy7MWEtNb4VauufL3asdu
OivpcVKEWvce6oOeymrEQvPDhJRJOXStGj6xSRU0K8OWI7D0GeUb8CPtfErwdOyP
ZFs6zak5MJXEVxhBMvkmW3lKLJLcfNhmwLTA7vQqWkqzJK9B7p8g9q/1mpW3kEky
rvZ90DryWyK2QSIVj+EHw6oGmpSQDhFjqaiuNAAMXag2Vs05WoIRzYWGPm3l9NR2
OUEys8hs+vyXojN5MMgcDyKc2aPpUXJwKBFmNlonoQaecsr5W9+C3cAizNE/L34f
pTLKwvmk0OLo4VQqhUgoL0nd4JAIqG2YQIRuI8Wz5s54e3acfx36MiQo3542WPuq
PNZ5ZmYsZj/ERo4RpfpdtT4f73LtAgQCmmMvKSdhJtdaMnKuWw7dsO4/UBiPNVgq
b6ZOf6abS4oJPqXi9qPA/53U/+BA7jB/qWk3CdkeWIlOwm/J3xDnPbTnK4pSrEHO
AEapn/AB/GjilG2/q3J/WV3hWV5iSjerNGl9hJ2OZcJodKojOuXkwWeK2AZXQYSC
X6fTIFfHOtnLT5zv9fA6mk7FtT6VgiVSiYQWscTp0968PPrbfe1/HAr3JDjjuWHs
kw03DafsPHymln/UTKOb9INXgOPcfcXa+ovpl2KgeaeeGkWNvZwc9q5b86cpPa22
XrpgfsBjOueWYQa3zdBP8+fah4Zp1PznAfTytbukL5URs6IK/Bt3mU0pstCdITkw
rWzojnhRte3IkNPEuQcAte98VfJ8zn88n6HWZ4A6t0DVpeHFdu7ij++yO0skH/qr
tlnN67BUSfqTXreI5xlgrlSCiE43bvIvFpaJc5BjAo9cjN/UtL1S9eNw9Ixdq8JQ
kVEcYTdQqLRbMzS0M0x/e8FPYyacQIQivWSZ3dJ0U+406/ZwcI31V+0cym9JP0oB
UhaIU6SzBlQChKkpP9VZWaWqoLf7+4a+5NWN39wIYcBm7isT/aDZfktR7E6wBFAb
EHf0BPD9ypn3DrITORPPelZwd+oY4RRdUxUcIlLEu0FpruEUaJoMd7poPlqfT9+u
bIkoYGuZQJfUSdodb1iq+KGAuQPTO6oi/80tZVAxmAdR7UK0olTU1Nfzf2vYPOhR
th1EzOMl6SQhMcJzbBuqZ6fS9ruD8vWHQPIwt3RXMOjM0X8B0HG6r9gVRVSM322S
HcNaRVhTaysqtICmBlBudPkkdTmc0OTPKR+hh8RYiFO8Vq2e78TWGIU3jnjrMvyE
Of0dPtDeq/96c1oU5PncZHIwtP8tXe8jagPR08X2idflCjmHicLUgI3RTbo42JYs
eWTKktPBlQRWaP6+MDccGQrpE0qAWP8A7cMfthXwLg5JcOs2g4hBmFduQ2mzWKqs
t1Pmx7MGg9ZcnrgGep2NyfiWhRClOYfzusyJBvLAnXOCA4IRmZxw4QWUDWKUnFuG
Xv9gMAMsT2Aw2gAepv4gnnPkkCpJ+MxwqILzV2l7XgKMT5TXM859r2+Es1obE+Wh
RrC/7qY7M2sbjUR2glUeDd9kV7ZDvrAvFOWGRkjbwvFiHimHSumrngs4A0vhdXwu
2rTz9vhyrn2Z70kaiJ3TodcNqh80VV4CZoEszPlhMnmknIZr6SEHy/U7IL/K/mPc
KTCmuRb0LpVxcYhb5xAjBcoOXQtsrsGMr8c+qlei/zDY774Y8taE+CYXu3Owqevn
N9YbV1i8XIFmWtHSst+xey0sXVOHi63dXxb+VbNLEuUWbI2VonF1denih1+xhG+9
oQ7esEcS7WvLFVUtam38EqmFEM+IuCRQ0HqvnACj3YNjp/MYdUiNZ9gUBvN4AivX
8KHkMtxfKifvWWpmAQ0OCM3rE93rQWTE7NtQ/Onf6jgH/KzE3dspdJQRArU801rz
yhPj5GftTKrj7rFfcUPmnOxZeO1EhfsOmtRbD/Frbv/5uycD3G/JZODRlTegBOOy
Pi2ulGRoD33uvQzDwucx5TdL7+XpDuf8/J4zUO1QA3Jaa6ApvwK0z+1bhFvD5C1g
z8+JPH9pfi7DDCXjb97VPFTuUN7WEgwj8t4k3+YRYfGZQp/IbzBUWk9SaHgfp07K
no0cuqYXfFPU+GVgKhq8cahHJ0nN4wsWrw9aSJtJVFekxld4F+qZxjRilyIl81bt
Un2A5mc9DouCdOlhm7KEBNndUrSViDxguU5VTIkLzc8U6vh/8rOtieIj+GsYh5px
X5KA0DKFQNzZ0kDsmMaAr+CDOx1IFIxsDSm4m5dzFq2oZNUeyHenv6XSfH0VePIH
F9o4X6ux1MxbZawKlO8D6j2XfY2aygTNDFD9LotiEYCSEh5N+2pnT+El0Sgz0CVb
KIuty8cFeyz0x56J5FRQsekEEvc/esX4Eia8TAfOwKvdid376CRyB35fU9FsHLXQ
dwU5HxNoQgd+AqsP/6/XkwoPfRmnRYbIgsj69Z3RaUHK4Ick4VvG2c0CXjoLSvJd
W/JFESKLrDLDQVQK1KT4pQ0vxjI7INiS6qrmwhNlz+8rVUYPiE7Lr7sHsKVjCLIm
Sbf3eDZZwW7yOqQdv8ZmxBTo5EHbPX5eWHwv6SVLDPscleOAn0e8oQ/ewv8W6rdj
RngASNrksfDFPmJk+fj94M13WL77GAt0dSK/FOwURaQcIcbSWvqJPnCxGXMlqvty
zxbeyYCCFWyMS7PKI8RR0ABGQZCdRKN3rZdNq0sqhzBJ7MBGPZBfhLT8sGkYbr9F
HnqissFv2RdKhfP/rLyPJ50hlQw/+O+Q3gy5N39RCB6ndKJ55iCHckHH//eYgg0x
OHGPAKjmvLFTgYR8+3XMR9EUD1o2h05cVn1T/MqhAdYEy7dsdgoIgyELSdJKa81w
TInyCARgXuRkQdrtdeelnf3n0LJTbWr4qj+SyrlsAWgwHXHi0qXsbflopCMxHDxp
VzAP4zilr0zXIOraaHTy2UodfUY2tbo582CUxMZJ6/WU8khP/yHdOWGgZoEut5QD
re2prlOAPRKipGz1tTgnGN9Gf9KEgwwWHpMKN3fALxBxJhizHBLXV7oboIHT4XJC
gdgGTxEGyYWCDvhNGdcCkS805yzxH8dpA8T2GAhmUsffUiH8d1/2t8kxrNzrW4xA
jH789G/7Yd+HEm/RXpUmu0+o0PEjNvDAgDgX1oRHKAIfU2nUHbBQmHEH/RAAzTvU
0GVLA67ATNFQr4wq6liyZzra7zyKaMy8Xg3lYMTgN4oO8LJ3D7FjBYrW2tAitGAB
q7efxA5vSQFqJEKiT/cMlLjRe9DSRw8p5gUgyDBV/7BkJyBN9lz1PjjKmSZS6991
gMaP9Y0pE2W92LBfrPbvkA6p+MiLfv+pF61XEcdmpT9S3B/w0JGkubaDepvWJyCB
VHhkTDLWDatYRclnH6PhbkxgcFrzcJnN3n64NCq7TqBcHXMS3zCCb98qq9YOsJI5
6iC3faxegu2zrQDhRaY+2ziXgvqb2nXXHekAKcR2u9pnAsXJLjFD4OqfS0JjXv6n
thGg5B3WyylCOI5BJAv7X6ZVMi8tSN4dtv5comAH0RVoToTPGufLyACibV9dVZg0
khP6YoariRy2f3STQ2FaMqeQdyRv4KJwvGFz119Oo0xLqdlSZTxM4fUdzfmk2C0b
r2DwBVjPSvI67/zrADW79DIo+xYX9WK3lk24xu5GjJagCsYhnIVl/TjnPE0f869b
Ta+nH/CsYIM7VevPuGMoLexnmZ2wN5RPZLKSU79kcMl/mOEcfw6UjGlf805qcC8l
U5FZY0zrGz9x/nUdp3QNywSCE6Z3+xsvAft3pM7hpGh33jcroooMSDVfVyKCkywf
LoQXDTLHbte1dQF1kXTTV3IiOdx4SAE72KkjwTBM1OjZ3ADSyN39Lm3U7JPhhwyk
0ShJyeOdbIcYEdPJ/sDknT+tWhXqoFe5YGZPfh20l+NcsAMZRSn1+0XeLGwQ0DXB
O/uv4o6ET4yNIARnlxxxSODunGjzPMEle/wuL7ipwcQZIqBEDHaD1REj3v33P2B0
xTltuUyvYQxT2JMvjmEyuBDpku6FwS3wTmgSDFR8js30vSt4NTaUAIlYV0nUj1ze
Bnwse67SFRqUv5IMHuP2E5Jmme6XAb1rKS5b14JpxQYp+h6I8qyxP9JjHMS7nM2O
NSXVtBdsPd0Yw5YkyVNRHtNQPYLHjD4nm08M4fguxu494eIah03aoVdMHz3zhRBc
og/BAD8iF3xUQ9RTykHufHJR7wNvNWUjJkfBBKe6d7g1tjaSrKQ2iJqYFeSGuXHD
bfPE7rHI1wQ25ZaGXyVn480/Vyx5MaXLFcDFHN12NQjUgfT4A+zHwK2fMpAMW4jq
nIAgyLV/g4oMPnREFuIm5/BwTIvncdHywcwHX4Kx0UA5AET8ZRH/R+SwhMPjZtYA
SdMEQZg0eQIJ5yWrPqz9uslIj5WL6FvxYJovdDTlngvJJCmKPHKrZXVKpZClG3IV
GC+LrqUA9Y6tPiYV0SYvGRAUn2FkrT6wN0reiRI4h31rzsSDbVIM0TinMcw1NV92
3BZ0n6VYn812o0Ojx7CLNj97K/v1KJJC4kV8O2IKkmkABHcX9mlSa25VqVtEpF9n
uxJzm7GtCKfz0IAtvSDGtqFmmBBc3UFpZ8kfQpU8vgVz2sNv0UEOv2vbAg8ujYOi
Trs8LoyydeG103sP9bMVRDkbQz2jp0SqM9Ab9fIlvfvyKJhhG68YBHKFIR2BbUc+
OZS1ctWsl4JzSqzQQ9fRol59TP2MZhJtY27bmOWaer3SNG1Iinhvcz60kC+CgiMQ
02TFJwK4y268iNH7eTH81fEt9EAhpAhFrqMvHTQEnCMp5fUjPSt3bFgoxTz2492Y
Yfi8Wb/WUbZvaYMZh9WCvIMP5n9oQOklDzG5gAskS7N8U8nO8B2dC9zicgrR8jtf
/hi3NXwfDu0kneB1bKc+n00Q+hjSvLwehyAPci2x1/Liw081ggSRD0Fba/UQkVuE
UO324jxcMMZLNqjeUql+nUOgZivUI1q4ZJW4hZuHvtp70pqz1v9h/3LBMlX0lJA2
nQyU0Q3dZ6k7o9nB+OzxJ1earsfrFAG5Kr+r55npbU3fxooZU0pDxvA0dCsj5gRj
BhWg07jZXrhSYOGNL9dXCHd9SYudNZ0zBVPmNxum+XmC0KNWY6/rvaVoi386oius
wJBfLcQQi79XCQaASHdzFMnY1GwRfAUb0SfA5iEZLXsGB4ZJxpWDxEVOCjMf/H+b
Q7bBadUh7v5fxkbGYSP7SoIFd9CE5Aa+9nicRh6IHdNn+PPTLD0H4cgYxi7ZM+5J
oYTieinduerhLnDPcm+BU6ZVuCh4F+cwBI4fdGfuexn0LfM1EDoK0jqMI5h0abwg
g3r038ASjE7UXecNYLyUdnf3UxToZ+pdmbjwHzOqFdggj8wNBXeJrTTzdNwXHOAn
AJ16jcyjdqBPWupoHUX2py7TcJK9jdJ3gyJk2LmuCG1oYVfKiEL90ONNGgLeHc3m
9MenPQcSsKqt4ikMGyLplfdBOJf9EnI/n2NfN+bncLWNmzV/7gA6/1fiJANTBYtt
gpuxxjgvzYikA73r72nbHz9wjVPvdNhWprVZrEKBKd8jNcwNQPunQcVs8G5X/o5Z
N239SoqJi4S/ZHXXic+6KE6S9u5srDXDHccXm5CeoQlHLhEt5WSEk4cowrLGBeoG
zgGpiRTP/K2qxyXPoSEZokNgLIjsrrVyBgUlxtEbf/Og+VMGl9BAciP3ZdC6cLWm
VUms4DNyZ4Gbv+NhAi4ns+uub1HlUfsLLbn4KU5dlsOFO4Fv15s/JwDFSZOl9c2r
Gj2IAwlH9SXDtHUbHgaf9HbOjM1JUi0CGl5MHzRaxW0KZ/sg/0obHPbNyBHYmZP5
gUQg5CJKtjMe2XOoesfAkjinhiEEOMR/hNGtUgVmpAWHtwW/m5+sbwZDmMIyPwT6
x/wAKrHplgF+MSzBI/S6HTbiMzcV4sPNhfFuvNkgzyUQEgg2mX4N9rMNMBe1Y7y8
fMIETD3yJG9TYJZaKBRRXkCx0cFZUoxtckbwjRs3BgmhtzhIeBR351KD0XobPRlz
Go4zxQNRxTFYuSg1T/sudp15iFymnLwq5r1yGTuY0dEduHxNmx+dPaBccn1qROU6
p+SdF22QqNabERpUq2GBH5AyWdUdHjPMVxH2UtuUBsZvAqNK/LhcuVfrRM1717ZW
Rfbq4eU1TKB0p67Sx5LctkXc5iXtXgmf1KWeME741WwoznhCd4Brd3hcGrtt5B9N
TecPcxbjQKP5JfoOyz4j41oKpYseD2JfyL+EJiLrKhs3g5dsvHVYGY/mlD7rmqD1
r6B+7aizeQTeZwHf0DJadgzfvE5jWnzL5odoP3eJwQV2qwdifb3f50fLjj/wugFj
Ep/4/EglfEPBv3trJ74GUpyFXtWLkdF8lBKB9k6gIoqgstQ+tTmn9oa6QKHPqfr2
u2FilEl/ke1jKApB82podBdPZGga06oocYAKODJ5HpWDsowSkM7ZT/0OzD7YpNCc
QPGh6HinNcJQT77888TmdIVvELTSylE1YDlPiwbr4CKa9EP/IToEAvmS4r4rub/3
JB7dvDvj6U2ij1RJsmfpZujIToiTK4BbCaydwlVbJckAfPooa8nuZJdU5VgJo6px
II3dQGAp3h+bK+KpGNraFc67NmpMF4sPM5zXmR6onklmmDcJpGzkQuKfXhZDK8On
8rqzwin82FileCthuoUs33bSnxsM0x+JLchV5y5rK4/0k8VnddvEnNap6oQCdHIw
5870cWG9VNEyTKcn8mkUmx9itPSpYd512PdACuXWs0srN5oT+6hZkhVTOsmQKzdM
7/DJ9LTETmnkesoW82/RZ1aD7EmeAhL3v+6gbkS0HNll9I5IddxMhs/lewsgvEHW
xMIbKq3ubf685q0HjZyZuLYUiZVUT5jeTWd+LpwgzPVm6ZB3qiWKdeurVEpQKNhF
XLfXB2id9v0byp7eEsjJyXo0l7SdCCdSDddczvbPw+RNpGcMMb0FcydRe8ofusk1
+XugNoA2VzF8lwFuPJDYdAk8DE67Iz90ZUP9w+4UgmV0kTTWd8j6GJSiWjOTsr3b
1VQiaxczroKfw7p9cykK3ilXLv/K2419iG82HWOGGYVq1MqDdIQycBNEkP4zNcav
3DuhNoAXej9YAhjxF5eBX2NalzH9+wVp/CxwRsgJC+q49YV+X6t9cajYv5Z5OM0m
eWbRXDDdKkFxBfZOc8gDcmuYyMgaMhHl74IOxbDL4tyIjNtENWVAt97b3H7Kv4eE
kcwV1Uzjx7wRwTz7/nbq6xxYd5aXq6JEQbgOVcqQghyZuDkYZt6siQxH5hfOulZH
jjqz2FCLaMfwg4ureOZp8BeYTJozvIjKBFLyCJ3LQwyUIfwq/DGYGW+ZKBuAxUm+
uId1n5bKIo2NXlFl8ScOxdY423bFzkWjaImUBu5f2GvkTPvQwgGnfDuXTYUYUf1e
T13uhLpkEeDilXyL+h67wQ+EIWBxTCxcsDVr9x/rOfPcPcFC2KmFli2BYS7u9aGT
MTXun/Msn5U7Ywo/u8h2bSMzKFhiDTvgtjPFj6ilMyMovlmmP5EcZUK7720z4T+s
e2Z4r6sr9G5Tg7VRyOKAHD06fm+LXMw3DnC90MV9leLScJoz0amZ/I0jXcJ0aTf/
Ot58WTtos8BqQ4ekhO4DWtWbOPNcAq+ewgKSnPUEDO8kXmYJam/cYtWupMkRrHeW
3NhYKCuMRcvQprz+z0I9+pVfxOwVKXp6v6LqczaxHu9+hDjk1qPucKkuYiba9fMB
WsA0suS/Vwgl0NzCgij9SxawUr+eS4o0/aBjE6ID+myvlUKYHPe+DH/TGxF6t4yB
e3qjjfa6OtkBOBySrFFcSl48g2ONp9kRMTtMfnl10cfjitIaR7k+vRqF0BbjzSrI
YtV+fviI5QlgCM83DrXTIa7mkCdbg8Zqa/7BZLqG6kIMR2QgM64b6Bm2Lvjt5bAp
6wnw/H9RUdXFxpykklvpd6mwQiY8m8PzMcnesG2t0XSPbJijlHRP5iM4WHX45pOo
2/i6flKoAFTAhJBEGQS/bzm00/tosrWOoxCqelrxBiUz0D9klM5ylMJgUA8FmMP1
DnympC2u82LF3DdUIZeqny/OXgSe+mHONfz78TBBvGJOAFtQWmkADDl2FU8QMb67
SEJyQmnl6GvV8OO2UtVmcslKB1xi+SVst0Sy+GdkoW4ATET3l5GMOJjmOJU8TQ07
qL816Vn9fTnxYYk8KQc++A+5lB9RvQvLqct7VCIBdKIZoiO6fN8HcbnWdR0Jkxv0
GoZiFpa5EI73X/yieu0xy8JTSrGlGhpUUameQiwRo/bdkIGYUs2LVaH5gZfFlM3h
RjT60ANGWHMRFTH6xFQmqV+cXlxZcWCmfKe5SliJBD4lGeTSq+STxp4weyvq0PGH
hgKeoWA4RJGLlLD+T7+OVR+LImq1wW6sse5AMXYKy/B4EywpRi/UXIe8FFh7NWk3
Hnda3sGr5+wuNp/kAzHMZW/Smot/HdLpBeDSANXW6i9e8ng2pmbCeGM7kQXBXReC
4EylcJW+wBVpJVlC5SEJraR5tzfE1aK6qL8xcyKKoWWBIhphuToXPUXojJp6hdCG
KE6/vF4ZfIy/x8x+0VG0lG0nSnXNOGc1Wdl017RSWCLOe7sJVtPVz8GUonoGmfES
G85ne6wqbWKBivz0XafFFMnpkW18esQos/hmlcr8ITp86ZbFPODmdnBWHvtgVd53
myguk/kaUCgljXjOqpW3HNEWVChrGFyiKT2KzcygWwOpqHUmP03nUBNTaR01qcC6
al4NsbGb/HUEPUjoME04aqum8DbQT3tzNKo7QV+e3eohccEMrgy3qDxGJFflVkKX
S+gLVhJ/lcwttbZD10vUnn+V8f81Am/icLQnT7h2LiBrZ7MFNPt/CtmaiAyfjHfX
nf/KXwGkQJSpK11b6njNadGa8u4+rC5qYjGS673is38Z7J42bwmEjPowaPiIunzB
2Ya/YnSd14k7nKf4JD05iM9SvyLKwTzesKaOmSeeH7Vh00pCAL0eVIt9TMmLyJW5
4LarZ17TambfmQk5uWKcjMcj6kFB3gbTpBvCeHTwwX9di2l415E/h3U32QONjKox
u4BTXO6FRCgDo3sDJ6EnYTH5LsoE/A7NQjayl4Sv3fyAWOCBNwZNLjsEjzvDIkFl
ORcsE0fYIzskAPlCetttHOe7WqAz51VFEJ3q0WopLotj9BklR94vTEUN1DS+gc8t
/qIJkTehH8oI9xCRxnwPIg0AlqngAs3m8J2XEvOod868oInF6XrnezoZ4ZhTeyOz
udtxuSxJuwhlR+5q7naOscqdP4Zj51JnEAzzgFYNvlwPB127xGyuKGHbDNNzAT1a
vtj3hiit+ZJ/4tgypJLvtFQLp3k+wmiYU9DFnLbZZGsVCWWesFDyIe0Fv4EXj+Y/
npSfZCuUbtCpiYxB6WpUpEziI8T2zZuMy315xhmGZAXsuz6482QCeIFMmbYEctxK
3aQtYf2Pae4bgb9S1I2RCf5ZnfkRwHF+yEr9K7m/h7y78iWz/6qVsCfVRPmnrQ0Y
u3JDqpN5m+TZcV2oufsdF+8vYMLpCtVtmpv+BXPJHlsV3C1JDZfXmNwB5lB4+pwi
kya/A32+VibuRBbFdxncxDB8lq9N99ZRuYlYMTZGk97E2N7SJmoJhfb86vI6mO8Y
Lif/r3madHpnPXLTWqDVbjHOQey/OSEQx0aU1qUELmsahZFWtdaaTcsB+mlFDZyn
/qNWecePpKBuV2nWntJ7thbr7GGdfWOl7wN9P8CLpNd/k+/EmjPgd0lxCMhfPysJ
vgOQQ5yNhdVojK8MeVXxNLXwyk3z34XUX88UskhaNdRjMD/tHoDO3zFUZBC0gsjn
7ebF2bbKPBjfnzbyewY4Tq52Roejoq6VyRstIDkmR4RP9D+UIn3cI0byXyIlYTvh
2Gw40CpB4VjdxHZI13WVgC0HpqwzO0gEkZJiNW2lJhJOYPyNpCuUhJUJrx7B+R23
dxiXVfVimFDZ7RucNnackkz7Ugjht/dqJn1L7CruYoP8HvtcnqX1rLQk6hvb9yMP
EsHly4Kc/AxGpdmRooMAs7d4gADbfgOkHDh4VuoQI4X/U3TmhqcapeeQ9PclNBvZ
w3VkhjLPcuERDwJynNKXwu1sYjJiEK4z1ZGGJpYWO8KV80cdR97pDtxZbBBoHN/1
nXdh5fkzxL6B6yoHBAxF0SoUze2LuQatNvetARAXXPbcmDMzb1AznhWPfsn+OR1m
eYGfQKy1gtnmJMkoe+imtiblOHG3pxIN8PXVFUr+22OEkrsofUv8LvPef243bRFK
9GpF8cGCa77P6siRn52gMYCXGjNdyP00sxYKi/OtZz+TFreR1aOTSvK/WL1kLAP5
guXH/FU7QWLJRFT4D0jJ9hNyTfb5KWdO0UJT1w3A95sJwghw/d0gRP/CSVGeEQY2
5kfqjDdb+C69wzUVTZx9SC0BQx969elc/K0CNdXMNd25/FYoLfiETKcOBzWilERX
PVVRVphWcv1GPnRhFmtKKAdB0wBQ+qA4Pf1mKYj/fGBmIzPQdz+0fHv6reaZFL7F
FQX6m2QRtLysGx9nrKY4k9ACpMctXKTjzXgpAzp4Xlixst39Yc03TmkUg0hAFuws
eQ8PiAeSuN1ja/9M/1e5p7HeVypeJdpk9qtUZ6Eb9sJQh67BNs2mk4IkhWML2S0x
3Ud+JUScLRANpni5FYcN4i+2oowwB8/HAHNWz67OihRWgKYebcGq5rdq6iYBGxJb
4giiQ4rcmdww7d0MsAnPXUHdH12A5/TqdEOsW2a1xKDm2mArKbaUmUfuSTWQFkuC
OlDBSMwFazVaVEDZNeT3Z5pg3DHnRcS4OC3j9UL/+ArQuBweMZf6nDipeasQh4MN
7KNyZdZ/z9gVRFjyt5VWlXe4GfDCXjqkyF94WaQGGISeuwFGNz83Sa0sCketrO/8
Qe0V0SUqNz9R8e6VjTTzRG3+qKp611p/jcdeeD42yb3J8BTpN4ezEufRAi7ZmCZ/
73tkUegdDr+5UMa+BGMGX9ukV4N1GHl1qHCRs0CyrK43gCDLF6Uht10pE84pfYjN
81RSczJmnpp/hHYxlCGwx3qDaJTrUQiCg8VcGt5xdafZNU6LEqSv9ylPvE0LxaT0
7JEUCzrxA530qoB1BhnTfYCzAjjqli+okIfB3xoz9wLFxxNUBFPwtWopGjsnb2lu
tyGtEXRfW77UDfFf8h6UmDFE04ViOQylUb6bZqa/zTu1Ukw8gwcNynteYgXaPt0l
0JktA8UbE06+j7/C0OAP7T/ObFjMONJVjrjfYpkWrmnD+AmZ1xPeieE/PzyePYDW
ZwXW7y3GXqY0c7VfaweglYr8awuU/L7Q5eXYHd7hyczd0RRJOdBrHLoYJydY7Ii7
t4RC+40r/6bbZFlbtJudVEHygsCvmZ5lx3O3XHmxcelRYA0VoWza7vGVBk3LeuCn
PToTy8iUEf1u7lga3j2II77DcYjk/VS46pQID1W3vTxoycfWKa/4YRiyhVnIZoSt
OcZsViNKNjJKOGGwYEQTuEPuzil5dc6ajeTn3QVWgfUq3WldoSEWfK8wV3HHVGcp
Pyax7rBfondj8zRhGtJA3iGDR3hLOHjOhZfEvJG/3bIkCh1vaIgTJvBIU8Zzx/k2
O2m+Rx0V0qFZSjSjT9/o2opCm4zlOGi0QpjzeKY7lFatXanFP0e0aMD0IjjX6yjh
uY/MnsYKEpt4NB1wV3iFOtF0g99avuLeXB9tVeyRvuKr0ch4nsXMPQpeYavwS7ae
O/pKQv5UlMzzHm/fRWhRjjU3EkCoefprfSY2kRM3LDgvImVi8p/ksMqEX97WydMS
8RPzbMTpmWG/8D2tFdy6tIaeHtRX0SXeNckWLwZvMFWm0+qQYPuzBiuVk4Dj0Nw4
cKrXUJ/Rpd1QG8q1MM3idjBjrDedVX4aV01AQjBn/nN5NQjLagTwKVWBNd3L9j03
CWVZU0QoK1FXXKcb97K5IMUy6fjnY/7SYtFg0yPHMxlS4AFBfgtncnKkOdJH8/M8
yjQV9FligSipBNvbmTSyAUUPbQ36WCxuXJ45Ivq3CO/5njdCdeF3VleJ8XAiGlg1
aIUn99N7i8FN+aAXac1DX7chjd/NN4APnxiibH5Utp0RTdHQ5XO0R5DXyleEaPA4
4cCitXYvMJtPzhc80E/8tO3aav3M0ltUAHDVq1X60xWJZ1UFHfZkaW8Uq3dpQ0c4
YGvlcPBkX8M1TBLM1pnYcslfjBeT26aVSbiTX9SeadhT5dEoIXVYUjI8a1tHSyvN
4sZvcclbrKwhhAUHquStm2YElIuvrDJ+pfyaeQ7gcsUzThMtu66V43kqTwZZKO/G
tw53EByz62dfLOJazOstcq67cqN0npEYi8zeaGZANGKtrX1Z/eh4lL3Xl45y8V+2
u3ZWwZRRI9P7j54bAE5LSICSBxVe26hHrpqRgYJHuE4pPg2/CHrJjy+pS06jxli8
f4oajh97pEBTNtte90N1UBcLS8Ed9SYsCBYmh/9TX8zVeHa6KBrr0YChyB8Yb2NU
TJhfoLrXaBMfSXzU+YImUlXOmaZojF0nx+XlNxV/9Ttj43F0X5rkw/V83d9TEY1b
o6xVsUkZHGlzYpJe6KHqY00WW0pzgG28CGHvscvANdkKic2/HNe8Cfqqk8G1D1Xp
746AEjUeILabHl2IOUvcMB2wHppBKcPSLbwHUIcDAI9TSVzNwa3yGNWCixuoT7gU
LXvRS+Pzxn17KLnkMDh0ryNJ3hFCU1F835U1GJCxMVGC5VaTnsSLPpcFQ0MEnUD7
FlQzalK33Yq4MwHg3YiFy+V5VWmApTXu/wamAnnbWsTJURsRix+n5p7rXpq3JayS
1oMUhTHDgmU/9E+WcHtAlcBIXasfM4DPHjhJ3hz2RGsuu+Pn6U02EvYJr2FaTkKj
gXMvj9T8+FItg2qX3AX1jf0xcIvqjl7s5E3U5XquCVnhPFYiOA7zaUc6WUBLjDWw
H39EZrpBr9phwLGJ5opLgNFt1dElmoqfJU/Bdcj4E+EJwrejiu3IszMc2HJU9ldT
4NMccSr4Ros5Hd1eW4q6QHixJIuWs1TmZ+mfXdNzQRufs7eB1kn9dVFbrl7fMBYu
92MIW2qsvE+MrFhvrXzjmhiBwYUMLPh3uS0j0yzFZIEgmZ0b/a30crOCwrhQo4AC
GWjeZY8pQDGB1Bep49XF3fRfWFyvTjAIQYyuE408F3EEUJi+20r0+9kv4D7U1LEQ
VVFjlj1FsTzkpxHpwhqrNU7ignAKPvlk9jdpufFY9rLnxSiDei60Tht9z+ryD+eT
Hfhgm5sa47TGcJUSDSeyYl3PqEyQAWM6gMEB1lPwDD3coY8KkvnX7mbSeajZF4Ll
d3NFrfkiH7u63vtyMS47X5A1ifiLepv5PsjleoF51pMgw8l7Awj0/2L6bdZ/LKr1
IIE0Y3WdAjaq3unxNm9VCbUpONq8XQXvAmpog81jUXro8o6TtKInMI8pcwdtZ6Zo
hDFCqkRlCJ9ZNlyYHspKgDs5Hi0sbEjAQ+0BPQrYI/8He665TtfYTojcRelUhHFg
2lEcf8Gyq3tOLHz4YskMm6tujMHh8HHzEY4d+mwpxQhdPzTA3iwrclfOVerRye55
XONr3hvaTW4EMLA+1wX/xlHg67kZQtJyJM4mpp1w2RRg6czZ5tcw4dfWVO7tzn1y
VWHaWMiGrmv8OvEGVDl47c+FV7v3VIh5TTzHdpRmPRSFIVHUUFjsONTqaQaVzCsl
cEffEDxu3Vpi1NDktfihga7/GxClc2A7bCvAZ4iLBhabKNTHnrGs1sSQ1WbN8zn5
awbDSzhqkCw3zeXm+SUQBdaudo8k6UV94+4MGA3Yu7g+LeycAlvrRZgRRaL5nRZf
XGDolfarHPf5t8fUEt2OWHGptuht/oWpkfegxQYUwTG1LhuWfyaSehHuEAEPaJb/
98CFXfatVs4cqnXC6Sl6K72s0wMQgr426nDoZS6n4u7FEi1tRA5EyNkXAT+omN9I
YeQlmO/UNWrHKOmMByM3Ed4DZY3zAp8KnlfZPKQdvVv0vCZyrH/B199NaGySEjd3
7w1g3vi6cJfToWDKPeyJTkg2Tzg41Ly0mI7hZGoDQbaQ8L/X+YIF+1P6Budg7S1k
+Xw00ADCKYw53jKvt7WHSsJyRPTkmCSMF+JsorbaRGFwxKAMNjHNbCtHPt2shPxX
v17zjGW3BDqQp9I3knhrtSzw3MhN+iQq8uEOmSdR4iCuoAt46IQ9E3uCHM9GXpEx
ePo+qwwDehJ5bIxjOZ05fo7QCgFRdb/Dyps4BQLNneEmGBncgrogQZpOGYA/KM/J
QVF4n/eRGSXh9kZlvxBCfpdFM5IqWd6FpRD9MH/bXPEvzeqm++th1+dPIX+pX6Po
SKJcDGQ2ydqziqDYBMRMOyzuzGcjMNWspo/VKCtiLUfbu/UMJQWNP9FAT2aAJblC
Z4cZl71Rj+FlqGsSgBgOnYQm/5/qBYd9zHwvlvl2xhA7odWirdLS44v9VdvexzNC
F31DwgwBmMT2lIEe9KBp7vqWtGx6E7/BLL7keGjLeqbh7IS+rOXRszwCBpSFzuv4
oYhrDc8y7RZ/HY9ULGMS+EkMb3cEl3MniuUduWnN7NO0rhGzwnhWSxc86xxMmXtA
LEt/IJuLBow7fkeATkb0lyAhpzforf020SAUBbGcpdnhZ6QaYaX6jVTRrORLcQNk
AZGnarvdzRcHZf8VY+MTDSa/Lz/rKyGWaa8cBO74S9iR7NIHWTuRvKVn8KywoSO8
zkum4y1TgKLkcZEGUO4OTn7YFfMx2nYCJFWeFI34mTj96AmwqBpmo58m4kTBGHtx
F4ok7jWlwG40zo/mFKG0Fb5dKQ68+BIpGdOKIhmspBdqiT65Rr17QYt5zOlXTm/K
gAK9p/YifgXcjFBXUJivopHZJjwHRScRApz+4ReJso0KvoB/F5YyUUo6cAMZFrX5
mpaXYV44ZUUfXwQlfeMgB3sPVUGoGjPbAf3sOBphijFev0MM/y0Eql9PYShaEaDt
BlRgSriNn+eQeb9HR5ukpkuqU1bJeEwitqRM1wKcWKgDQ9ga/xpyO5tZ0zRQXwM8
tlRzHNAfOSXhXBHnOSB6btbFU10VFmsIXaF2PSVkV319SWKWMMqknET59QN1k4vq
vUtSxw7yP1MV3i5X8NQSB2mR4DlbRljk9KiC6OQ9NgYq43gQdChZEV+3uU+N0YpX
wllukxaJlIdFM3YBHPYWEqOaVFavDMUZnxGBf5iNEp+02i45kn6V4Rc3kI7z8kbP
+Zn8HOj+rIRF0YP+EyK2QGhcaUIDn9QSHgirZQ07sddV4oJKAD32JHOaLsXkHIkF
dSPGPc5uBZw39NFpCDfHGEpWqXedraUImVC236NFXZCAVS0PTIBFTY2VHqDpZuaO
iyyQVgCu+M8OmdrN0mhopLQ2xe+yZBmKP0qcy3eNKdZ0gT3hMFKrDoDjvj0B5t0H
PkB8NA5Wh7MMEou011F1G+CKCf9twLwOKKr8zMLvwnjlD9cXe6gekqYp0M4YfAx1
1hcGBMvK2izQPe5EDk8tMS8V+TiPJa7J9G/xhSk2YHiXt2t87AciE7y2EALUy1Gu
EXuD0vw1fQYSslPFKzhgt2VPFFVWhXYl9lUAG8Tue5o79chnMygEq3W3kD3j0XLv
nlYyo2BzwqIM84EszjUaBrz8nu7bTQbwdz6Kiq4dfpuGKqNIMETaLBiPAFBUXyGO
c5P2CVtfcKGKkcxmTufPl3ne8QLySPr9upq6goOiCDBHB45+NPPez7ZXZGzlh4FT
QPVbDDMsS37fmukBmdj0cpUfCor+TFWIUIX6oxLS6iU4EgTZICY6w+fJDHHBJYbm
OPZvCOSVLOHdR3v4KastcwubTbgedIbLorKDjVJy7ns5v0eodSAicLhAL5h4UThv
jNp0tOjzavpaPNpszJ5cLMEHmdYaYxPjMPQMzFxRisEHR2N8B5bcAXxf5YWX832g
o2LCGlI+FZcBEaEHmd5ZyYPIrDP5o4/IvV9e93YUG912PaRHZkxJObQiIzyq6PRw
Ge/fN44OZeaQH8sTYADMdmy546v0hyXJqwTRnctnSDkH8K1pyZMbeHUEHbCDCboI
+/j8XwO0+X/vZvbMiO8papXEnz8anWtinEVW6+ZcN675FuOO6+rtzSE6mplpZNhY
V0JE2VDfOG4k3nI98XP1yUPzRITZVmA40+P6VoiBDTQZSz0dweounucG6aXCGLca
goPQC/i/V5hA2PxdmghK8oWDMdMILT9L76ZSvmOlpOe5GriF5WitXK0bp8pj6WLw
whaxyqaj1xiS31V1DqwT0XieD3Y16FI2cjZ0TZcsteEWApjiDJOMz1+L9gXn4BVM
+doCwZ5mJ0B12vAx10eIC+zOXM6DnJytkpqXWx9V3+jfu3JMhaQKtivu+TsTWJUb
YKt6T1TGutjGmHNzoS1IWohYC+zGQQZ3B+VUdgJwf+jp6OHkA59mSIiDbnxaADBC
h1AmXWFP3N2HJ99acrSVJ4POwqz4jeaN7w5wcVqHIJZU1bX2VGuWSoSrNsBPk9yj
LDdhEFA8TBgJnY5U/f/xwbjKuoJfE7Tccv0UEWyHLtH46cFO3Hce4aL5/n8lmjJ1
I3vTGnuzKSOLh/nbG3LVxOjSpDcZn0F9QC2YC/WwLc6yltKeQVUHgXdDe6jZYpPo
b8hJ4iE53/rEuy44niYyLMF6x1DYqqHqWqDj6SLWZVX46K/q9Tvb5tnk16xmj8Ib
/Qbg7u27j+CSzp0NekCe1DmATTY0ozMOMZi6wI5y9nS0kdr0oOZL0sr7hM6HJlXb
50D2/FCH3eTA8d4LlJ+Eo8lxGoBwXwyr5q4vTY29KpiVTG/MkPRUsmLHhKP7rqki
RXEMn8bUSmkqXz/dY1gO3OB1pYyxKZo/aZo8YX7P0RxG88j6D8Z2hy7JGi4hBhSt
TEAc/jueVyhS/G6Go11Ab+eWYgty3FTCTK/fH99bu0N4E7SSvKNUmO5whvuAWWcT
q4/zmBxCvuhBSXujmxzCRqnefQCYc7lbBhiPOOhh61zF+9YWWOGa2BwnSNEuX5IA
56WwY2r7MC13ztWIuezW1t1ST5601+iG8QxOWlijWUaakRKSopF8MyD+l+ZFGslf
FEZM9qnVK1g8YDJrNsnT8g3cyMMvZLEXTp17Dc1fCIOOegMj2T+GNqf3Bb/99xhK
ovgC/W9AhJG7Ve+V8OqzjKnZtChhQJhKUcI9R6jZUfh/sX6Exf5CKQze5BV6Y5pg
caUW7UjTcnJ6aSx6Z5ur7GsnT9k6I5CMSL607yB7d1cQo6AZK9EjN/+pHoGBCJFK
nriKmtCvkzzDDeGCLuRCzSbrh5GU8WpIZHl5jMJRPWqOuBPGzYDAPuY5WXjoYDl2
NsgtkmWKTu6EED1cgF1IPfBbSi5jjqUh7GECPVMr2gM9+kYnTQvEy+JEozhxezvy
+OZOvagJxlnhkjY+LzTeipDgASir1EaakNEAKxqB+tPGL4ynmbbgUAI78abFHftO
IQDsLyI9ruSZaxo075Lj0z3430pw0111rC1LhSDvRSEmfecB31MJK0rWHsiL8XhQ
CzPoFuJb6L6fgL3emzC75d8iDx1vAtCXLxHdQYGCur3qE3m1Ih860X7cQQ+kKUSu
+aixFBS/vGZU6Kia3zaql74c1yPDsf6V+8ry0HCCHIRmrA/585lZuoKAqEcTR/Rf
qizDHyQYm2/qL4EkcfGVZwCfYyXWRJZTs2INGQ9+Jyr2RC3CCIwhwsCzKvPnSBep
Ec6Zmbjb7xOqT9u0T7hwlRhHtL+8tOdMQ68AoF3imxMDAUj9jRx8v2lEa1FMqvd2
kyec8FzwDyVl2M65d10GBV6ovInFlZP51C586fmA1PZqCiCngSmBd3/SwZe7Kb9Z
NLl2uo49WAh1FVYygCwR4/qsuOd1MkgI/cU+1yJyyZsVkMm94vAR0bPn53a6WLoQ
LKjkTmfKDLkVrWau6dgOuce3ASMTi8LHBtAtemxbm9e9dJpw2KkXg+VbUI5O/Okf
YWoUTgo6Zyr4NbD5mZcuwvFMe1aVoHo2qlEo2TpFvDO2nFDrXoYlLZQbdvoCx36R
6OL82aft8zXyrVzyb3yAVW32Y7xwSwn/XCkQG4piUyoH9/9HHG/jHTZezAiemphJ
B9YV9/rXQiuY51mhXRixPwr7fBwWSr/Kk6BKf0qsJKMr0BDR0v6a5Wcpa8xQUwQo
sVV4z47KCBqy3qHVPeHdqg0ZokEkQvm+4CUVW+2KPHnUgUVrsoGcYvCElNRhUv1M
7ifq48JY7yO6ldM9IhybJSVnm7Ece5Zq3jECHCNEjTmoDPuTipXgpQ/8iMMVUvZV
/uZvbnF3QYxZxBR/fvLG6N1EX/A8r4dPQIEfXd7hgegM6Aw3ak+b7YlCXjUORO/j
MG2Oj6AXbu5v52ZkH5dyS3aXeKsGWSsFtAgLaqeDnll570jMct6umROWewyOyqnW
a1/BsOtcZhqqBk4rmvAwiUS1bLtUv1I8hl8KmwiGSU1/o2DOqH0okMKt7eEOlGON
l0aaoxPaZqh79dGyvpH2KTVjkBdgrfN7w/wS9jAo2Qy0qrDQF7n95Cq1djAmTehX
u/I0QR1Kn8aSVXTSq+zbTVb0TZPeAxu4ved4Q0QeSAOecCE1/aDAtVetbkHwH+L7
4W/HfayF5acuTzh/BxouOQpmx+ZeqSjXM5ShTvINHQhdrkZ18jnsOcpmxzL/5oQr
F81VIz9y4RI0vqyas5QVmfwOcaYq+gcIY8Tu3YTJzS76PSP8OrwvfokPID6cyLSe
1A2fo6HdE8ohXSIrjz/uLTlyRJ7B3+F5bA4OKbL8/jRT8wdZzI1iLuDoOT82OEdz
/jZOaxv7VT/wPirDcTVRe8AUi4ZEtythfVru1KqLtuClYivA/bHcFkEfugd5pVfY
iRHZZR8zjb1t7PpUcDXXTZl3ZMHM9HBPGWFC4JdbJ5erLY+Ufjh55zoVQUeg2Brw
MVrudpsqca+8fzfjDo2c8kX/NNBsTZS6Z5gH2SfTn5OE058CC/oHk4QiShNBMToF
Gjc86pDANbDFWP2B9iuP/CmhDf9xi7syQicL9gvjegRlOJ4jGTp1R7rwX9qlLVuT
0y4HwSc0YIaW77FjV1ml1HisEItijNOGuQfWicnm3re0Wzq196aQnCxT5sQF+vDj
s680vNet2UKTpOh+4IYY9wfQP0b+K6vm9sq4Cd4HtsNm3AXuveMuE9IYo6TxBo8H
s1rasqsq1GkOpnk8Yo977Od21kAAX4dyomYZa/bhHe7KMls+OaZyNotCyfabYubf
bIZdmWRiLkSFIAvBoHI1dFbyHdFjPALkMV73JuT/WQWMjSJue5JPvjtxP4+4/LvC
rcKQMkYCdLvlar3ZsTex2dL0XJvpe/h4NIVOYq7a9RzdXq3ZZ6Mc5w4O6hCS978q
7O21xnD7dwYYFwPkASSLNOAOqLYXHH+rxO/H+MZh0/FojkVG72Axa/ZNqtRoBKEY
DdSTRQHx5BJZNXRx0G6T7Vkeqb2m88YUoVALAlPXTtzl/AR6TGMriGt89/a7/0dK
3vPiEhSkX18KCKrxbnq8JGQ3VwY0ySTfbZu2aS14H7IjDGDSfeFisiXzUzDjgoEa
hbV6PRdFHbRQa7VX1ZAF1mzfws/n01SUtN4xKkwiP0CamfNakWHOCwebyWsfuXZW
5jmP+3heUm31cspsVOsYMd7ybSc1wcE5kLl8so4+P6GvAYvhYaLw/euJjwguRX+c
r3HkDXDGlNLv047cpk1isCS3QVQLxRQbwQOQBCioBMbWbfx0UB6Pn/rAjdkZ/uPc
M49KmXV53/sRK0qneN8jFwTJQqK1Sg1wDEXuPD4WNM6hMbcexQMCkh5fSqddcgzm
lQ1FzNClPEMg8FtTGeCmK3PWRru4V/387oQD62okiyWiEmW8klBrUlxrUpregtD3
uNnBodG9djny5As7JWt7Gm77CWfmbleb2Sezh9e+3Mnmer1R6vg1iMoFucTd6Jai
RJnvIeL4LbrdDzzOEPYDCg19PABkGcPyu7xus/sIbEtVEK97pc/EoG4kARyowIpz
kBfDFjXWl2OVqTLnIzNrksQtYNmg7DJk9soQXkGTiaM/ESKhTzWNHO4ymfOf9Fan
SxLJEauI/y9QI1oIx693/jCVZQuttIkkqsj/AKMDKmL02T3yEoCTnIqonhENKLUU
aaLeQOLliRyz8gI+LnI5rQlwWCsyvOW5DrmgI5EB7TsQW6Tt6Ik9gH+RFn0plPkD
rVfJiMfpXUkOdsVL5f1Rn1JArFo9M6L6mYdlVVsKkaBY/doLAYJqFrf8NigY8V/+
F7pBFkg5h7pRtyYjL+5wyIgd8rAGUZvUluCtt6O/mwi3sMX77IvxA/UNhy3qnLFi
AalyD7IHPJemO7q+EHQXjL45QpQASM9r9idxtzCnfrKl2mlJFk+h8HK0hktssMkD
feJNAyHc4eX+DjthOwgY0qzXdkLpoA1q5ZjhjAt7KJgDgEoltRVO+6RhVh4QCewr
wBGDMqoovrniAIK1yvkR3REkTcp8wdEoSuduSoqYU7xlwDlaqwwb43ibzLxSigr9
mxBFhiihn32USL33X7k3cn+/VQBu4i9uJKjYqQlBVN4HcIfZThp9asmJcgGO2nW+
NxZNNxYtHwYoNIW0+K5HvQ2x5lkmPoagtA+KYWTDmNIS23bDCEKxyzwCiJRCoJbv
d7e8ksdVXLK7QjASD8CYcxx09rA28kry0G9vd/2m9Wa0V2pARDpH1hOpjyrqf5Gl
12SsXbZ8McjYn/iUKEOOFMC2NTLis14fjEOZ3I8fqSwb8Q6VEObseqpeUMx1pmJY
VUuUqH2865Yjpd+83P4dr9i0lrwp91vM9ydsbyiq7dWw0gmqPgdYmp7qsHD7sRNG
CbJsTDs93K9XSpjWOW7zcCjIekOFpVo5Y+NVV974oIyXwS+9miPWwMev01915t36
MeFMXbXQnR1TlYuiAGRId/B6AcWa+h0mxvpCzW+A+aUucZ+7efEE9LR5QFT5x5mR
2khRAPGKTkJUZoLam3HuZ8eORqbVsBQUB4ykrhbNzP4HvfciHuLnzkkPwCykrUri
uCmVCWQCJeScJNkWrJoRrqZHF1X+2oG35ZDCFyLCALJ3sHfSSjNbX0c7uWJ7pnWC
jyhEqbmMcpOlR8q507+NJ1+4SZDFGB99d+MA23crB+kfSr/hnq8ydqj3dYPJVnbF
2czohraD+QCdFla7NwwvSeeCoi6BbsYctCQx2LAd9cjlDUVml7R77JOy0KbM2opF
74a7T7PzyseM9i5Jvr/Tb6A0JTJjyxeR44cz/5zQt8Ep9q8iQ7JnJZNkrNM0jaYa
XFFgcpvosLZzCzYR/97nP4HQ9uY2Gn4xkUcJjObZU9puzBV2b9tPzpUdwcGJWzuC
dmH3/O/c9tLH03PAaKDESiPLkv63cKMsoIPlfJziTjNdK7f+fjjF3XhcFQYZo9hZ
CNxXxmfAjrIoi/xxI5K5WWU4Cq73ih+mcw4rdwWx6VAolRI++N2NfZh3XggvGzVL
cZRVDBP2wGURJF9P4yJvr43iHrJ1RAZpo91DAZTrj+ndO8NrKGztGuDI1jABwKxH
9zUT+qqng2Lf1oii/rdD/NE6QOz0+tRQ6E6zaEPRebKOKY7T4WOQyqZM6wQWKzgk
4SvxQcSrMA6ck7yBJ6yXkBIgNmVC7FGQMdBUCCfc0xEpRm3yIvLVl3Uy9VIwWh2h
w89PGCc+Nu4KCDV5x1OD6s7uxfo0es6/6Z/xvMxZqwC/dXqC25o1TIUg+8SJkAQe
LJa9xrnDzlwRHN+M6XF4x7YbZRLWRRZwxdMlsMo4IcJ69oIPhNsqeLR559NbWAOg
9RWcwaSUzzoRzw0EZ+frOsnZyqgWoBHCE9Up5oKrsNoKuTGNgT/o1QJ60H1awFH7
rl1RanoKhf2Zbud6+PWp6vleVl+yQx+9t1FZxKHbiv5XoD/6gg+Ow0qts4PMhHAB
QS+ql2tUt8YVQR3PzJwqGH2OmZz1qzc6Z3HO9RFlj6835XaJjYAHOWrZBHToZXDG
osjJx4rxIXil5VctPhE7CuRY9MolLoldxV6FkQTHJpnW7U7Zi0hCeN1s14sZ7/iq
nt0qgXdMoeadq6Pp7C5DyxhCVHJgr7jnwt9M0gV6Gv1BR/EXLk3I5NqOfYPs5Bit
sjpDbC7ivWpd58ozOlEhdJK0ldT/BdAuW0SHSS2BAUPK7+1tptS3lt64ZZrM43Fg
yzY4U8jcX72hNT4Lr1t1gFkmWu/hjNozGHuc0ddCbUfqyN3XxfrcyJvwUL4rTndY
KfHkYwcA8A2sSXi+jlFEJWBAbdtGjz8nyHLcyM3FCgGMxfEjj2kPBI9zbMpmtKlW
48o0EnAsvqH0Sec5MwusMDoJSVwtxgfhPnA+3Z8f6CN1gLBBYh7BQ06dp+qfreYN
OhYUao6qDYX9G5y2p+uXfp7V5GJHlvCK7Uyjj8s42IzoK8i2Uj5AGDDjgkt+vpYS
VjX4tybTaNHXbj98XS/Fptx04/6MO4xvYqHyJz8ERU/Hf+o6KXMqaS0s8+Abpek/
iynXEixglDZxr4bs7QD6H+tnP9N0TrOw9a6nrBHCz1acAcFj2Lvqapkfv7EvWiIB
6FpKjI8+GvWYihNGFoGRNMjtkSx17+BRjv2G7rqiBlG9/n9TBaMlZGDIVip9wXj0
2XIn10aYeg1YnfO9oJAWP4w20o03o6lGOL+JBIMl8tq3Aw9Y9L0sYUL+TFn4OxCU
FpxNi10sIAkXlr92VOd6cC2SW06yjD/kj+qLfjec9/H4VD7+0I22JO6YaB2l9iAz
HAiQ3gekhcO929m4G6D8LyPdFz4oZdJF/k7icKsjTwx3fmw579zHx7RjwEdMvI27
/YiS2UrD401uTkJJI/qvrDaG6lieqDb+0DmLI9l2YbHrvjVEX3kppGu34Z+igFRg
bTPE0C4t1cwXgSjkK0t5TBd39ejBLEBOxSB8FHydIXs07fUwkDMZHvEk45T/zMfI
Bb+jWzf3GoRb+IG3Sbd6Ux2iJKQ0KyLAf8syovcmMSSdAuIpQqmKPazz5tmiObl6
lSyUKCSkzZX+w6wFIvg4vXjk/GYjbD36hVoL4fYFDO1FqI+IrHNDXlyMbse4/Tx0
0rNPGF1QKxhKw6YgLZnApJhVkCHBmbhMa0xWIXRor2mJ+z9SLUpziKoZxCVI+VUi
CvxhtZi61LhdT+XwbtRchCaASlcmuP73tR9wdkjQZIim4EK9z+MH4naJSy17QsZq
0Un4pYt6/RotAiOtM43wZPjyRvTx9XnP0mMxlZZ7ZrAGaASUgh3eg2nLCr3yUY9G
aFYqktEdu96lzmPkidWgyb94C+a65rw6lU4cRuqem0daxnZPw8s+3ZcGG6OwlO/v
DE0asFfKY3mzXdMQKthVlMcwhE4/p9EXk2T9RLTG4QyxMsimoqVETsbyMSXuBSVq
Dqorm84Es9Cpj6QyEL359TrPONvouZPxVtRDVY4qcXCgOvLw9Hbn4lypLHeyq5RV
kz/VxiHbSG5E7OjA2lWHLK5tw7pRP0jRsl6GDcLaB2WffiuhOrXU9V3ErBPG8saB
pbfYveufrM6HXnhYA9DaeoWntw+83yoeitcRzuSktUlGPBvV+gZYEw36XrjSFMF2
AzaiAIip3tgxzQwtQc7pooviUNEclJZMxuyywacyGlpHf49x0ndMojdPLhPVojpE
jy7lrKlsRDtO90NAs5HXmVaXVrhUsPSU/yTAm8uwuRTuIDURPbre4niZrCPnitx3
wcSyh9k8Mvk+8QYL/aqa8MUI8VU/f3sDbn/dOf0a4PZBQ07PLgXxLMkhJATazoVa
tUwlLOZLlSP9qIw09xMdV/VdKXY+dzxlW4UGchfh8s0O15NhY9tJ2NtUjTdO/3df
Dweoi3xl/eWbeBwT0X643HEoxYUnkFJEXuQnZ0YAi6yhjrkCFxkT27QDo4hMyDH9
pLVg0JmpkYNAI17383Q8PC0tclPEj4zmZVWWF7LjXoTXEmp6pBMU9kJbbTDqHRe/
nS/VGupcfiKsJb4JjyPWxSMadniYKFxScuQ2+fZj5GjNwBRgl08Qpfrk+Quozy4O
GmJQ0/hyUkllcZcU8DCt7nfoUA6mfbFEYJGvsPPAPimKcUhoX3jFlc/t8owsf/Eq
Z8EQ1sHwErrEyaRZUsRWg8mqulcFYLMr4xywpwYVlKsjpTXVlGS//Cus2G6talvL
5SsFUNIs0s0FnfitmvKWUCV32Voe8xq7y3AvNjlYWCrxnXTaYe3BGEUaGD49pkUm
TJansaajhkWkdeKR6Ta0QHpQMeP4rS8rxaUutgp7Ug/0oN21Gsst3wi4YO+TSdLn
61WHv7Hf8jwVXSWuFRW27XqMR+/fMypC+FIAOGoYE6RQ/HxHBngqrIapIUbLSPl2
I/15PdwdEeM2jbY5TyXnwqHo98FX+vcXIZNQ71LK/rOkWwcqVY+dVW4zgo1ezXsf
vrMiCKZ94EAuXKkwqioRQue7WxQAVqrNEzQsnd4HBSkyqVRGQMbBcY+CkYSJxvol
JkqXMIEzTvh/LAEzxY0fhac7LPMEcIlwXaDfw1Ugd7jT+DwG8YS6s8ey2vbB7CM+
ygbyWAP3UduYBEDclcbzpGlZBQ3quBMs7B7lSwL6czY+39KoRPSEmBg/muCtsFmA
L1N68WmVPBl6wucUTu+eM1lKrV49rk5JGh3Q9aUQ5lUg4palXG6+wbCQuzzKvx6L
6EANSg4yJ+w92JuZIN/rMmrwvGdzBGt8U/tO4ip8al/JITDJlUqZGCHMGjUkTwOj
nrYXZ9s3uAh+92r+BSx3H9zxwNC6bNIpibHsTAsFdFZUy9ZtP5tK1/AWBWHdAPnS
xYSi6l8I+Ep7ctLnFGhdLkZGBrxgV3q/5Vb5uBpmaKBOCwi+rj8HjQR++lhwKdyS
ZmH4K/cLjCgLGfbDFA+BYkjUpAoKHzwpSvCVYJCju8Zl/LsXRRjsbAQFSMArfRZu
keQyzyj3UE4Cm4F0QZM1RtWx/nFvKXVq4cJuDA2UrmwM9jadPCqN1iqmCVob/VqW
5v3jsQb6ePOMrYJSpLRk6H2CJBVUMs2DfC6KxTAnnmQ7VWcu40vSV2HeOl3yQVC0
YbA3gHhM6ZoqX3uhMT9LVkRNo1zSJxF9BA+xpjqH5pQKadw74DOQBtJWz2DQDiFp
WQWBhNMUFqW6wbbAIwHGWX97RaC4hgd42PPx4K47Y5Pjf1KrifPeBhtBkvGtBvMR
hBbuhttqCkTMNQ2ngXQBOMPx+/lhP1Mex2nVTAxSQHWytenWQSExgqPYwOXLmKY+
g850IubKYlgxjQJd9TW71JgC1mKcZEc4l5b6HJyGc4mQhUQlAlFCG+UaQeVP03C7
+ESc6Q6y2fNaBatJrj2Lg94eLhSalBnHZ38nMmhcxMaeJ91LzTSIAOyCFejwT7Y6
vqtTYR8nKtxmqx+IUDvJxX93XIIUoc6Lr4/W/qNMVietVC0nbmkHFZBtaKxoks5v
ghp+UNnEtcvFGU8NUThAXTBQqramsCF17wDeVjw6r2NKNUWdkW94jKPAIJ/9mKKa
jJkUp7cNzppWKzQKciZST/WD47zQm7SwtHKQkydAqiBg01DaJGvTSRQxbuuhH94a
0CGwFpDp+DhP0VZNu6wVbyPXKbxFmAv6pNkLL2TeMLNrG+P0Gh6rxn1ci46ElLd+
7SbSM+qpsHO5mxCFnKzIuaZWiIjz8CbZwYIM15usCmuxyLqGJbCr5eV39L3VGdKM
Kfc6rNMSGZAw84DdHwvTiMEWZLixGViFH9WrpMpCiC71l8/wo82IebjHgaL+cZmJ
S5403ZTEg+efVsIy/zp2DzFLEkF1WQjzjfZaGNUkOEdIgLb9KjmjQAGRd8e6Y6tQ
rGTjzt2i10u7xaq039ke6qlZcm0f+x0tBrBuXde1BsRNjwtomE2FPLCQWEkD8EKw
v133RhD1w0vz9YKNHYiQJsFcRy4Rg2E7EUSa3CnOhUO3NVs2ID4YSUMQKu3xSdNz
xBKy7OQfA92w8ZbWbxR8TRI/H1sUbh/OXILA+5V7zR7pLkmJnuEA38RXoy1m4uuj
Sw27xwZEhN40DykRPqZ2nQtFA3gV4XQ0txoWlWiZIwmiy8APxKi7j/R3pZ6yw9Sa
C85Jj3da3lVcVkR2M+H1R+lNnDhTj7lcP23SqI5/l/wXNUmMNmq+U6qdmcAI/ftq
pHUQxdtreymDa3ir9pJn8cFPowstUKt8bxtPH4NL+STZKSAuBIBj4CmJmC7nBy7r
YnYmYHTbKQMTNe7t8BXhJIGu1+X/rJbnl6ElbTFv0y+jlvWyNJlIk/GWRiFb833w
6nF6SU20k0IPGnThNkG0X3bsprb3X9jEDCi5u5lV71BQSv8ewYgWe1y3RQbiOzmv
Xiukbzfq6BLUdb6UCblWmAoLb/Cv7nFYP4Og5I76tMRjl+vgWomaCTwBQnlsxrMs
OSpAPgUGBVfj1skCs6pM+xtpV6UKC0icRC4E2X7eCZKKjVTFT+iYbazMFZpdj3KN
tQ5jjSl1fqXsSSWMGN7bRhbjtxBFZ3TCoi5XTZrh2p9OUwMkN7ZPZcLoigoy+8mw
vo3lwoFhNXASOLY6NtoatNmmHUCnqwW5ACy9ADXwaggbOmCqOuhOMSVd4tlAgj0C
WwdQdOKiIuzvAqRiShKU4MpZF8AQrx6YjSdxsZ7L8Agw5ZjVzmlbWcEBSpk+K85b
h2WSLMOxAE+XiiokvS1fVv8ABjvK00NuHVzWHGR8TKS46UZ2n58HL0o+s0FFGPqt
Aheqo5ru+dEJbvj3D4wfm+qQsfQyjHJ7g+GD5lVBIFiHcWvOtKgdCU7AvwAG0Bp7
5yJTwBpQ78pgtC7J/Te6kJj663zzdrTEQxwnsPGPN+5+p+XIw8zOH08/VrtQNDWL
Glodmmx+NuW1ui1NnpXUgaQil3G2xpPu8yG+5oO+Bkj32A0DOyj2s8n7r8cOaB1z
UNROLu+OhtKTWeYJyS/iqukhXB/+qSTooCqfmn49K/xE+f/2gL/lNRBFpCmTACzQ
tNBNRKu4Tj/8zR9qHGQA8olv3AN50ENrTkGAbM0APNiB3NQImGIEJDt7T8uuX0xo
omYRWH7H7yZrewsWjQNSiMz8rGXEyhyz3LgU2h1cIUHmOnE3Ba2eJNeJ9RWNYnHH
YRK9Eyd+PXSLYtZfGtFwlyLQI1pZnUGyyEWbeN0M0P6A5ICgjbAG/w6D6GHzFOn4
hh2UM5YuQfivu81wgOt39imvWVek/+i69TjE18SmsFtBXS572IiFy3Phsu3e3QVj
Jb/aGebQxVxfXgfxXNbCtfumXCV5Vz6OMdJ3v515ERoGiPilLcpRLJ85/HCk6iF3
LwzWOqv7/Xi5taW0T9hm6UGnX/BrzfBQC8Tzo5Bwx405yYVs0QnP4lYu/WxFq9Nm
1fyobZy9oGH1mgGfMCwj1BdeoXllw/r+b3ComqjdMO+1BYL075IgIv2CJ59pjNSH
YTqa4uYuPH3ZfZ4NlKbQq3q9N9Bpbt1kMCWTQ4QUnucpvmeIrkshQZ21zRMurnVp
qUatP7ZWmnK6gUYcUQsEH+wZa5yUp9JVg90rXJp1QOIULBIVdXiIkhQOWAVHyE8S
fG8qCDpjqtESHeXQzwa+7Xk2kMU5NAM6BLWUmBGjqTWNZSAugjuKlXFMwSWa+Pta
uzBDmsPOWFJd5Y4rvsyuTKfdPbVfnp2VS7YB5IpmKuSvWiUG3Qe+lWcCnoPWENDs
m7wjrSfWC365Fg4C7tdxOU/lvLJXSDD5zCFyQfkfWXhexuTftR1HuYLp6uwXbmin
55TwxKI6Lx2jKCTONdqA4v3bo8XAcFBPwVVYhipn31efQfia0PXsVH/3uRtHvM6k
j9kb8ctwLeZeZriUKGwrCw5Z7kMGhH5gyAcPkdquf1r4jGwEdQkLkxRnLH2p/v2U
iZPEB50U5bOWWpY9sHuDrdpgINRRtBS8FVk91TVm9OMP08DhUjcQLymon5wnafrG
h6IVtnXcPZYLg4uYTm+tW8K4Ql3gez2q5+4QNbkTX0Dh2jxMy2sis77OskA/9FHw
bAiMLrRVmdUHDnHurpNl+O3aNp0gJCctc7a7bI8nMC9tumOgUEXGP0U2tdHVCbGA
HhzreqKwbNlnwNI1S8JCxWNBz9AbwDY0kUz5FrOrbq1lM/2s4hPDjl9Wrt3Gw+8W
xtzfODKFx/vK5/ZOpARgPI4O3LQ7VzdG2OtY6nWJQrIsWDwYi14MNGbuJcWF3ykp
aHRjqwe+OMXgWxnYKArOc74Xxkn1feII8ks/nNcbzwSffMOEK36OOAQFNxk+Dulc
HdX083Nw9GpypbDQr1w8SOGc0tiCfbb+fbhtMhOfIp8q5EGGzGtfn1ycuXK5LsxA
6fjz561rZ2VEEvY4MC7/jndBkkg2+UNo2yPIgqlTWmALdkyos3kL68OJSSbWF8CO
P/E+ZLfiS+1TDFkAYjhI+7AwDAFIm07+VyBC1CCIgbn9LAaM91NFgcFn6+iH0IYg
VcxMm3EDpGGJLZWxMvX9YbNGiZ/vs+JxCGklZoGakvcXygFABGOkYDqI+0dF9la6
opzVRnlGhWgIEgS1mgx7XPUXWDD8dfkXf9kONsTAe8g0ain0hntzlsx1ntEW7OHe
Rfb0Z77lp1+WEZ85kBdDbVH9RvaWdVE6wCv+1csr/zoiPRdQVQsyt1HV4tJHYT46
r5vZmGEIy6JiVq+2bQ72ttC96l83qmKvs43W14XdQbnqN+UtzyMdzzezsn1Z6U7J
h+vUSukkWoyr4+EYmf9xJ0H1seksCO3IWedbWkwG1tYU/u+yFME2P9M3DhbFOHLX
I1YS/3vSRm4mikvMZbeWo1qxYVp/xrXCkjl1O8GRcIgAozydh5Hm7XCFqIEWn3Fy
8ELyOvAwyQIUv9IM93XKa5ucgh+oWqIFauio4l60P6k2gadDd7H/6TqsNFEDT7kJ
IZAYxc5VG6LZ1YbtNDneBtpRtAbCHl0nvbHRu4OQxpvQ60bROi7naaCsHmHy0TFK
wnwy6yVShUhBv1r6Pl5CpvxJVQy965QmQ59V1dr2DfogmUBP9ijPN/jgDWsyylBI
isGZqCYkh0hbyq1LHVqZP3jGsjU0UpTSwsitsUI133EdJYRnX+X9w1GT0j8mAQ2c
dkSHYNO4JWYRbL9TkTNmJgI9/D0JK6wEMTtYPFVngstq9T4gg7mJpPWIVh1QcOG6
oRahDhbQWFmgvKTxFR+z/TubowTzyU1WdNnp9bHy+J8OmpwKNjx9cZabFC4weMrX
d3q+e1G95LoAF7rrfZb/aNeQkOBlZB19RklADV2RTr3f51LaBiUJaLBhWSjH4OPC
n+XszEm4NPUwZ8RRmTRKpt3gsRr1gZNjCngDMoJT76cyHq7zsexwCBz+Wlerq6ww
Idm3foy4GRNyivCuCX/EFmp21QKiGiuqVgS/xVe27td09pGxWxBakBNoqEmFBIF3
KOzvHCS2g6PlSO/Imtb1F1bJ72DQM1mzPyXfjpHKbSfX0yA7Q022FfJUEkwiN8yB
MohcJ21LKodxlWY41n9+Ohu6yDTRmGiPQCAzFQHCDJlWYDHlbPRfS5VR4f1PNkdm
Q6fVh08WXMzGxShcqYrWYVA84NPc6aVAj+6w9IyEQz/MC1PEsgyc9iXpAF8KtQtR
MwOTksN3++tTGqyVTZSIFYAMKTxuJ9Ncn05DcE5HjxIirjE6of5GDgPzJZhpumal
qDLLodVNNlzcu5IH9kJnvPiiL/4UDTe7wgNzpjBwtvxovbWxbI/K37zKQ8V6h+jv
OWVnbhbceJBkBY4mgGI/LYkdLuEGf5gLKbqvc0WZUI2T0w+pViaROzWz+qtdMN6y
CIVf6bk1MvXIOIo87cUqI+MjCFIJuXoKU0DvkkCYwB9i5++f70TZD+DzmD2qQxHB
vT7pc3FV8ab48lovQZMTahucIcTycwsXXtH3JU4yB2t1wkRNHYQ6+XWRpnhp3ZHz
p+1mEOmvyVIxTiRyUL7inINT7TkM6wwpJGclgqA6IBhnia3CxNDy4y7OBG+02KaB
Wt6sbE/eUgdu7SrIsHS9ALrUnH6oJt/xL4ordKDikjw2rrsfBsPNRW7uZZ4wLtH7
Zz9Q9nHanxosp6cPHF8IRrmeAp5IVTz3/UKrXY88dpDQ44WnQa/KEi/bIgcHii8X
FryHHxUU5WesnSciUewvqQczOmwcirvRs492nsZDYeptBXFUSfEFMMMvblUvb/F4
TcgduQIHmMJmXnXJ9ofyQldiPSJ3G72ZZq2m2sHCtzNAsqAj39fNr/e1pGHfRenT
HZe3aGM9WPgVCDYmb7EJ3ZJTjkBZC5kT8IuA2xDLGxcsgH0IIzu0Ejx7Dr2Lj8AC
hAB2t+MwW9h92T298TnGrw2sVH9JiYjokad/6Ao459zfqQouq4pZaDqcHRx50Mti
IEfQVuJPZX5cl/sVZfrw1ItzDiD3ZqQJtEkAE0EV0/IsKkQG7MFLeBo/OPhTpsvG
iPYXD8b2j/sINSrWFtK2M3UjsLjkfe3+fsJ357HZT0IEoIn9yxBHvB6CFdnYyF8g
oUdVc2eVzPMRXabMsBMtK+dSmT0H/xYiYL2zRU5EIN6011eeVjDCTqih0g5JHjPs
P93eP8QMvLAWW/QD1//3H11IAarUvg93wvqyVmVfm2q5oel3p4EqJHTCZEvAaQw8
Al4w9MAI1YIvAJQW4jirUay3q+U+9oz9jKInxZMOdkQ/J9WlS/p+diSoGh9EP48k
NazhFxrxdW4vUJGt1G6AFuOEoMcWu7kXAf4/XTGjkjwjA61du0jyrAV0ZzUWa7Pj
EKa23LZ1+pwA8Qjpqt2Ifp4LXFZrWwd/4Wzc0+1G3Px3XsMWEIiulKgSaFfmUspo
ancGyoomaXjf4+rBpwa4EPkRepwhksEh0yW1ZI5L680/uMhAVOJQVG2Wp+MudVt4
J3ZbKVIsP8027XRCnQriWwOqaTCdugUyyigi4fboNstA887jz3Xg7fsQean+yUxb
q766YFDo8ZXE6T6TSdYOMuj0P3lwlsTmPv2Ucu7FtPQeqYj9ykXKqKQlJCixNUa2
Gsnmg0gJnHnyjI5Ir3sdeNVdb+iAUmlXTk046RIiiOdDK1tp2EJqp2wzEZz6k2xM
Zp/3zcucIIL4MmrXTRUDMxrdG02rm3mA5UFhStjn8L747OpKTd3DV8A+47EYhkA0
r42/ojnXko5U2qdsVYJ+2nafSuu0I6ZACINHiluxIPcKKo8xYA/vJNZrKkOUWkT0
2vNnFczKTtuWm2ZEOIb1ykCY/srNzH0MOxxx6F68JkS6QjN0AoIqglpSw0D8j8zL
1cI2Ux+tqQwgllBfi+jPq3ymX3ywAc3Tnntvrrpu7DA1ZCU4xx6ycaKKN+8AGXSz
XSdN7RVpn+Qlpe2D0sQy3GO9HSPNWBefCx565/k5xsEVshpl7OTtZbERvEPTXWvQ
Movda9AuGWdN0ztL8DCFBVuaF8oG0OsRr5sYxc8GJ7e7gqEadVB7Neh7s4ia9VyQ
y6uL6183kDiystM0DBOTEN/zgDXex90r7wRM5haNsN9xT0HC1wAiInxwyhc/mhMr
zGIUIv7AnlbQT/l3sbYV6A15MgBmWKIKAtMVyK2i32qAeugB6ZFzUfXiqUxsEUiM
W8xbosW4SQC0yTBoq002+x/6j0Vi52jJLZbLFqBpe+u+gPXT8DZmi9X217XK+QP/
hK6fs6+WZYPJFU3zSJbdCv1cKgC3Mqub/5SxRpq+EZ98mUwIvgw9Et3FsRjHgCGI
NgoRBCIwFMC4Xqr7zX+NRY94SCtrI2ZQN4EuO+lsjMVuog4LJczMPYxrFQ4v+U+e
vVtMZqlyWd6ppvCM9zGAIhEnLHVGWh4WPYI/UNedQoAdQEb4mtoL/QFOdSjetrMO
NifH1fcxKj9ofR0tU/b6D3EzSUonHHzt5qShV1Ks4ftwuBmjQrSTQFuAo2EEdJ7U
O6s8NhgmnpwZB5uzqXtl6CegXz7ewyzAAkecKoiFOsHjjcyOi8t+pN1Q2kw9j/Go
TFPuLpEn1zwb382/nl7F7aOqEvLrsD4+EHw5bh5EpAKtpqt0YP/mToHHkvZjHV1T
oDcnvebmeqOEsJgO+b2I4eHiTYgGPYgOqJQAfNvY/LD3OoJSbYzf+WbFI0BuTd5V
6+YDNcdKDWIX9cLf6LH7fYD2ztynnxbYMDlZQXk/dYzBzR9C0wSeFAA9BcHAd2Iq
fVahNEj+QO1WTmaGXv//gE0LuqmS2YNCfqM79a9gCKSblktDrOqbP62M6TFbsGJL
TbXCN3n8vO2xxi7BlgcVAUpZyiovIu1DiYZV7XTymtxinjLkxFzeTVXBzk5O9Ye/
hUD1giyAqQ3L5i8FsWAgw9ayq/D/ArD5mYi2nJBBr0voubPV1CRaTdgiuNxBNGRR
cadKRZFfPUpNmWZ0h/X4ObSMYPRwt5wNoH9OuER+PqoPzuxU0K0RGKPRCX93Xetw
IecfxM06Btn98AnfnPb7x/kBGyw0QY6326cLqptZQT/D8bNiLh6b0SbmvIEq9z7l
mpByhTVPdOE9D6Ad37MX5GcxvKhBaaQucD+mCBmJvjvSXg9f7HHQhngrh20VHhCV
jaFzpngipk7YlBTB9PcZgiIqM0YurMAJAyNmJcWBUQfK1vqPd4S6k9zLQi71SXr/
nP4/VN80Ll9Q5dWtEvpN1sz0gDo36VZvRAnGMyGAVdIUVQnqSYxTwniAoA6RZ5cJ
1MJPDR9oFZvmM+Tk1DE8vQdnF1aZ+0xmP2UNQ3m0nyxpo4GfbojM7j68gLqbkzNK
p5frWsMg1TNoLXTWZLJKoDUzhapxuo/uk4oWnf2AoxlpARQ0cA9qZWU/YYZnsiem
QWhTfn5wOS91iv1DbhzXEzaqmU+UYZk8862lQo+03OkDBkruOMkuUPTxSrcAcwK5
gooHpYfkz3yuJ6rPZDgcMB8NX6muIkKOAYOrF78h7fDdpl5UkbhEZSXeENWMDw1M
hNjU+fgVIlIT40sAzInQGhlFYC6B8preXlmUCHmIUeUW6O1I/5pV9jiwjvHuMGZD
qY3UWleClFxBUzt3Zq752J8HGDmXNa7/q+i85ICTNlioqpL5vkp7WtmeLgI10O9j
p7Xy1gE//pRyBRxToz5bPq7ePShoCZ7c8ct0bsgyBUH8sclSQ9ElPv3Qs1udd6Qv
Ns40DsTpRbFVcY+SaIkGillN6YKKjV5GSpNC9iKIB/4IDnC+R5w/0+vY3m9el00O
TrhLVo1OTcYH1zGfUhzPdhl72ROllMOUuR3C6jNCvNw5UVznYTsKcNlsGg3R6lSQ
OVyuZOUVDA5h5g0wBZPGqghpqPkd6XWSVprZpjiCNz35i+zA3c8kcQOm0c29IEYg
xi7qrQ+XXP7FR0S1vWnRQAoiPhpcWdcS8lvfzQKV/KpBfNoop8phfFd/Z9deAJmJ
f+9eYNUR5m26+FpzoeMJ6XpPreUj3j2L8bVk161CPoPHvrYd4vRv4Cr0UMxFr/H2
lCEyxI1M5reksoh3WeO4av0IH0FiIgn4tCGj1wzELt3LpNjuuAOLEamQwAmHsA84
tXVd5uSiQ7jT6jpwW4SORV+c5sZBs1kD97dg4Unnk+z6tbqqq7mjKDcwnly07y53
sR+2s49CmHHHISig/bWpQLZfVUqhlKAtimWehtNonl3i+0X8nZVwaLKddNYX7tJ6
sTJHFvuzimzoQeYpe+3RDCvXi5neiay8TXJI/wVoo2RcFKIzg9ZePCSWrmksfs7v
FfpfZIv8QiTbFEP9aq4ytZj9Y7vTdehrBtk30Bx6RKG+6iVrjKXgyb/l/RFbk6S0
59X4L4u+e75PyvWWuTK2/F0il+bMCmWS6B432uQkpg1Fqc5kplP3qjkLoc+EHyqK
2/2fA9y8JWo4AAVBPZt13Jw+CBQrBDbmtP0R/a07DSGeQO91EfExp6t3EuswATB8
cVmydYtzzUBfrmy/HAwCMG1OKsZdz0N2KNWiGaSZe/mW1Az0L1yQYczmqwegqROn
74++vvyGjfA9c9v3EUBuQqobe2QHB17FjyeJHM2HX6hbjjqQK0yl1i4UtXKPxXOS
7qpxkgwQ8zEsAbroZoX/OwgtcS1JVvqJRmqH+pKq01ZT0lHRBHWTfiC1xkVTQVCu
S4CuE790ms5P+UG2ycZmuh6J9QWyhEwwNz2yf5Y+jBwei8zQukBFHrZl2i6LRWiS
lbMtmieEFx8hMMk5SbiPZi8p/u0VE1znENsGTL18Frdt1kwSA5RpRYomhYGRArHh
Z+vKNkS/ZVkMI9cZqAetiRJX3pcuVBZY4pd3CSt6xh4M8qf5i7sY8RfLHXyaCkMF
5+QX7yIRHiZYncQYiux5I0NsPrfmc5w8dkI8gRP/HojaU/972SzkhFKkoimK5LVa
5PsKzwrJ+j5i/RYA4mLSI5IuKwsUimLJja0p+t2rkXJs3an8LI+J+fIuNcnhgkKX
HFTu+VvzYETHZWLZ/jAYDU/ov1uUfckpzx7TeMPVD2ognwPlCBsNdmABjNFe6zRV
mWOeGf0ZTO+O99cY6Avdfk61JoqcB3Qq8Xvcevi02nNRasdm1JVAfo1RdEEUKlsG
gSA9VBK9yS2d4Jmh8L42gB0QgWRnT/0iU0fVePAwZbeD4cu1QDosOKOBcB/l/umq
SqRwDYYQvaEHFfx2v5+LsF6byXP3dMKhUfdNYhCze5pg20lwjrFFxLLNq7kcQ94t
mP1hcVSDtTJaK+NIBc1dLRzsb7DnAubMZlxhKnZUscKnz6tti9lhpzf3nGYMlJYE
X70DYxiAqCKAZ39w2w28vDXjSk4OgBPW71fNQcID0Us8Jnro/K5zJJ3F1jEVZGHQ
DvIwW3HxTVyAssuIKaaPthfrneiC7gJFHUKR0Ow3EOzLPldR7wAxeW/Nw142CZAt
E4OjBbzCBiusRM490eUTsaYVswzmhwj4TBFPcF0gZnUZMTTY+1JOve+0hxSiXnDG
+hdAEQsSBp273KiRd9x5od0+AW9eiDh6koF2bJ5rr3nt1r9frw1wYhAOLz3v9wdC
eeJJH2rIrF2MRSS3qXstn4oTcQBt7JqUhp5N2T7+5R+7nbmIUswgfcH5c5Ajim+n
aawOeguFfyY4szFXe+DbqaORcnzwyXHGASmYfVhXJFb378Tz8Lic9DCnUsaAc7fb
SZ1GyhWNFnPEgrnANVzkpCWHE0w3XuuxWbqf0QkhCSqun3KX65p2L75SUkoz9GCK
fA9DAabgremKsKbZYv8Lu/PwlWXym08GMNLexV+0QZi3F1V9RBW4qmc+cb/a/ped
Aw6clOztDD6Pr8M4v+wUCCwmX/rF8+e1cvc0M9Jn3NwPXtEkpOVXhwq/8oL7Ufi8
b/UhN6I7bhmQs1/yDV+NwrRBgeOaijTfRkRo0XMOuOXcsZh12Tc3u1Lw9uJ8mXeu
iNhSzUFkNhy4LcLHnuaCfvrrlRRdX9B54FTJpsN8sg2PF5PRrbDyub3ziUZVmmni
YRI0FvyMW5imiydfY2ia2/fKbmKSm8loVi4nmSC1vZNfBp9qX3nbPjJWcMHL/KKT
a4xj8f9gaKWMUO6FpTuCNDDIx5hDi8k9q8VrFyAsM6c/1wLgaVp4vVBqxEAetchL
DAwr/fHH/01natCeFJX3XIqDC3kIAqSoBWw4FIHTD6glUr23lfI1yRPDQFQd1mvL
kLcDdD7G1psnN4DDRZ7ssxjTEhGCV2ogQQrYkMqA6CU/3q4vojNT1O3NXCmjDu8B
24TeTdr90RYySWlBh8UdfCDwxSKGpSShodW55b6yiAkggf3pgGgBcS7RNU3aGIyb
9TuP488Zuru+wv1j1YDIA/KrRhYqV59vECFJLSC0UZmph316uquiFqqYdshms8/K
RfNBQTbCHGf8kf7zIQar71xSxFKfVbszQT/oDCRzEDnabFZ609dfeHSKAU9urZar
Yo31gfyTfDm5fAYK7E9R5kN3WxBV4n1Fm8qDcLhyXQJLaGT0nZW/SW6SGKThWLBl
REkZwtaFdPLoP2Bl/YxJy59vMM/OfFTXyLrplh88BfbN869S/t1ItiQykSjOdzE7
blH+w2yjuart37vztCzy8x98WoQzjN+NOaOxizfx3fi78gXOGZvmGyy8KVM9nMq/
4qjynMbMreMeKPsFLqU1Ru1xdrgPDMbVzjecrU6WLy5c9Sei7Q7wr93lJfhPia45
5lOA/OdV/a6nsA3PyyYB1l9gCPkRcsqMGkxHLnXh52/7TojD7quo4uB9ABEndi2k
gMKk44AqLztGYzH9UQelK1eVD2X8Oc5hxfDVSBTOfn8mNV/YAqgiUHC3h7MVoj8G
bDDdtiF3iASsuEV9ZBpnKYx8lsFLssbyaIYKEbiHkDcfAZmNILkWe3Y+K4aZqBkj
Q0OXazhrhDeWWgPRgyj0ZsEHAt1L4eZGjdYkpliXHK4ekC2LDTsNOpybhhYfnHxT
ZGnmR/pEvkgeOuJl/2h3u+9eYnLLfMIkFQo24o9rV1ejtLmHiG2X1kdhoDzXogGm
m6ncZSXvh7V0d4rWBAlLY17Eg7ae2Fu1CjOk0hBNn+lZoZzld4eJx9c9CddXaBpe
2FJKAc/Wa1uDIVjzyrndKWyo3q3dEarJ5wRzJmJMdsm0BsPTqgv8yTFQv4qgUOKJ
y+igUDGjwqvl45OKV6ggFGbzDW8LhiJSsd1qtCimyX5ZG9HhEdrinJsaTXA3HHHl
/ZquFY3lLzanTj0P2qlkhR2/fKvp7uIzW/Ov1pCxyRcdDs5J+2/NSG0KO/uNHAek
g4+XM4Ensst5sRzem0TlLE5Rg7sajyYnlzIiVCweGJGqBHUbWJYPY7aRXtZ9UEfK
YOPT5sHwaHc2j8YgIhCJDEVFK6VHePJxk+qGCleUTwxl+gsHMOL/namudR3vU/9f
t7szV1p8B9ins/lpqHIBVSjDk9HfmRIraWxMrjeV2i3xRIJWcdfFgYKkDY+JoMw9
amCEfhWkwb10OX2v8+pr3mT57rtrN+XqC4o/CNXelnOCPllm9ZOOq6K6f2j5xEav
1EBd422n3gWOdX9P/L+aZnXPAEmhtugkvaE62rPMi50JdnIrmOyhVw/0rBB4kXln
1zVmKHPiucLEPbX0du31KH2aIjL8fe4LYD28LKws5R4B2JILQu3aLho0A6JrwsLz
J4GZzdlNvFJYVVRWs+TGd0SwHjRZlMvMsDbqpppRD18tUZTz66BS0mAcWjIIu5PL
qQdRsHmhBRKUxw7dC/tjBp3qGxWio+djo8dnOhCdya262BzmfVEeNWs9Gj8W87M5
H16HMpAAy7UUEAqxsn5gKdaiAr+6IX24Qn2TNpWKWw68Ef8hxHX9EnVEz1jNsPgw
T6flNhUqvwv/xLNUc0YNJ3ihLosG7XjRV17UFM0qNhrsLNvhpFv5b/FaECtbUsFG
goKkUEZ40ZX4lkt1BOXlbnu7BzmS6afAi3GpI4FM5uD7LR9g5rZ6XSR0ewuXsZ81
r+slnLc5czQYC1FeNq4cGp2lxvrcuVh9rXkpVWMGVfHIq4Tk49PbLFNvt/gcF78m
+jOOqggAa1yCT6ifAoOszcRjaSmX4Y32p/s+BDFA7G/P0h1+1QDV8uYeaBePvPdQ
/JYrdZfL3VZofjcF7F2auyTOMULkX2E0ePG4B63ubzlKpOYyRbuiLyJeYh3VhWRd
7gQz2K0PiHTFmtuOk8dU1+S9NBKsn5kjsbildrUL3uS7/ErE3fVinYFQ0MY9BCau
pL4gcbV3X5Ph2ENm+VYtybS73vHPB9NsxMCif/75TjA71b0CfFYZUAaHzeXtLoyl
jyYbWbOR12FoWRPsrO86J1HZouRNvXXShnzc+oH+s9R6oB+guS4aPrCyViCPDx2G
k/T1tlgYKZMLJ54S5c8AO2KaoB3AHORqB0HULOHpRFpeNzpbYcG6nP7Gm/Tqg5NE
YTZeB0sN2CIbfhktYOyr3ig6AR3R9KV57mEEg1cQ3TeuxqOT2zFeOMBtc1qAhaiI
dpTzpUQ5hRcJzOCKhk3SzUYKyWEChtw+PTEaBo7OQuFTd0W/8oGsaJtWFsRUbPVe
bjCbnRaW9/1nmM03mc817EVScUC4VnoMj07ZJPwhwZkcOqCH+ELmwWW/UMq7i8Qh
H0cE45uJhQyM6VtvkzE+g08jYlOjNzQoBY7xdCsuQeeloqRhsIHYCUs9HPgeaJOw
D6w9cUTKBsB48L+7ptPP12bapzgYHlFHHWsNdYkKHUGaznIaaxf6fqPKq3DsjUri
wPZUXodGifJXZVarKMm7egctD5+EBcA9R/kjh/+fNHLkCkLFlTon91WZCGt6lG3t
c+Xt7yE4bUTB7HxXdYVXAb48vmfA9lDpmMENHooNwdhKEqfFGhReAoYOmilhp2uE
zsQn9mp6KkEd9i1eOM2K/1f9lLvMcoUAIPum3A2BReCoz/h2LXMiOIptheICo44+
HYFEmKePZWSRigiwdg1wx0Fq17hLW4+VXMVIdXUFA9azOrkQ1XHzd8WeOpWyYgki
AJ/zQyJ0zEgIvskIcIsTeT+jjqqf/O0WYUAw3wZapoFPJuseF5RAMcL7xThdS1Jf
DMtEPfFucFg3ieou9FZN1ZJGJTBNWJNfygviQvHUuw2r/kV4rPCQj6pjKNIEe7wl
8xQgviV92Q1If6nje9ioem83ezVSAhdK49yEONTzXk4kYtOAGzt4HSgj9l5pPJff
D0wnzQG1ZR/A5UvKratPlEn7MJBVQOggSeNcdnu+YsH7B5A0BSwCTsb70sNrIC+e
rOvl0H1r5DVPO9+9O5wpWs7jWoA85ZG1//7eQoLXT+5Is7L5DjJa6kIkNp+M3Dlo
QF9/O3YVb51mODQeohqML3KU474lmRHdtQFhiQJn/ybhKpZH2K5VX3Qek2ZX2V+R
UFun+uoKHei8QnUZ/bBKDe7oXUiVWI9izdOvaIPoazKnwYsVO9hm3c4b7UJnQnEw
eaEHvvJl3jzXTqA8YiX/o7B++l420xG6OqfK/aVxIL+7gWsNgbu1avRecqvP2zrR
dcfsbaWiIyhjQFEu0EmTgyGQjbvDm9+QAkMuhi2xew7A/uV5LZo9pzJVgVo1hRFo
IXVvWuoT44aC5KWOs6GRojWNK+y48kKcoyYRV8EvY0suLcUzi4TdJ7NgBTGnLRBd
J1p19cEqcU+fl26JBOIDlwN/ok2muvdQULh0zztBRs1nUTxaX1/8QxaKoKVZyWtg
OlvwVsRAH4D3pmHJrPN1WZTIa4TRlFkbkNgtBm7EdmMngopuoEbXBgZs/knheJvv
6LzFg0zu18Pj+hGCboMYSRncnEe1RIj4GRhRjnI9WYACVifNgLR83EyEggvDHTOX
F6czLKSJ3j5vBQnPrg6NXjQlCRz85N4QZoShGSKB4tmelgQZuB0r5FcOWwGUKoT8
mvereC5euDaxGLjw1bDCzqmbMimCWEGJfU9pYsWn5jDHjqul3JpFWnoX+OVoR+wo
WyiJ5EtVkK+BjoARNAJzZGShDTzfqH5nU+hi4PhzfF6SR9yvQFlDSMafb6l7qkN/
WIPqjKxFL2JpF0u+kYrKEPRqu8Dr9/1CNXO4ZAVIl3swc3xZZdTymWcb6SYTd/cQ
i0xgcsC4M0GjnWVlQz830hDXxmBp+U4NTOFgVScbBty6UpYncEPMmLD9rNgi0+BA
Diy3z+wuh9wxVwNyM/JYi1eDkJDTLABCzlWLLIq84p506Cfe1OezKzRg8FWwVtJO
HUUJwJYQeYrgvEYCw1qXt+mTVUPoG8yuRxrcGTpqUqzcIGHbhSGG8unCxQbwf1fx
cxg2hNItU4fh5zcjMY7MHNdlUDChP515gGAmyhscS/bJHKzYZ5PObLrbzELye84T
cj41XltsQfeep1EgKFZbnxqtpyEbInFo+8qJYSN19JYRC8AauSHP4GipF0xMpiT5
FhFNPD+FhBdnLdMeItobjEjVpqW4XLJ6dlgu/eFn14ajSe4TC/pyFcrxbDiX5B8e
zY9Q0a9HTwkcj5mSTFz54YOYtLCQQhp2taLgizCIBClxy4JxXBZgTowmMITh9JLa
iJTn7c+sxVJ/2VhaKzcKRutVJp5CQxYeCBe+gm3DKcUNQF8KZAM2xI978UlYYWgd
f3b9ae+GuE+zXJFXftLrQZV1KBMPbKMd4cB11oGYi2LAeYa2rTJwLnz3O91A0vIS
rop8dWWzJCHRXB6bdx3Fvrina2EjCFw8icA1babkGNneTtI1wOzFuU/DuIW1oSzi
BkyQnD9NsDLjFUlSG/2fWI8VHedkfzkZ+xWMppxe6picX+iNE1gmjO8XMJTZovLc
xpyXMbvlHBJ6rvwMQ5kcNqc4IV1IkAc7rCpHkr/b19ngL2MKoq+NE2g9Ln/+fEIb
2z7Z3xNpT1qN6fGf2iCcFzQ3GJ3nkuwngKIFPhH8ROfueHmYjoYgY/AbBwB3PZEq
vzMsAkWeFpuQ56WSnGJexfzWHxZcfE+OVrj1tjR/yH+jYUSkNzMRvLxucPxxleMT
76Iv0d9fpYztjF18KLBWMOPLYSu6b5d8CiCLAULaYXtFFRftYwOAoQR/mETmES/N
XtFFYzIVMuB+yhoDlXiUKt+LsNmZsP//DT+8RJPEOZ9WgHXDvG8M16l4vfVpPnBC
sjgI48g7poORZghDmAc7zfIVpfL6g+IHuUfYMeOxkQRYmq4iGwMMza56EPZJtAxu
e8mN0xQu+enPPXkPgiNheEu4VrqoZ+Cq6txSToj2mWa75i1kK5PtaRunKA0hEf1L
szi4r2jEHno7Z8fGXrt5DFOPiyUk6AEG9ZMMS9nPnl7cFo8D9lVNKOLupW0yVIw6
jYXLY/VMWvo5fkw7a2azvU/eeURU+LpZqbtMalDicZc3Jv9shQZyAKN2DtJ6dl7S
+ewyaq8mHlrvVvSS0B3B3UuPV6ngruOzoJlWxDHXLCvxl9PhfsHtIqqPE6C3uzYi
1Ga7VKmCyBEcLMBCqLKRxsTNCjTT9aOaznSBPe2eXvf0Rx6gZJuhyhgEJLcfbCHB
aJesLZ3EwOpN3putErtcdkAJ7ZuX6Hy4q72M8a1pkDbADdPlHPTZYuBFIT+VpMiv
u8kM5tSVIjQ9QVm+fraXC+666CNifkeP5KcZDjdpPf2uPrlwhW8nYX2QSxYEeeHd
f/ADdIlxNUUQre3ObJAYvP4GqmKJy49hROT9c2pPcnUVQyZ9W8XY7O3/8iTuqaYE
i6uiRszScP/k0RoBtr52FhjMbCWVHJh2/yexudMzwEptBSX4tyjyW+KX2NPhrk0r
wBq+SaLIbmJhZox2ztYUHfKkD4OGOqqCATJoElnEJVfVcfDe0NYA4Shj5B8FDN4Q
Y4H9hbZMgQk+kpZJ089AjScfqtLu37thBV4w6mcbqvlQQI9iazY7kXHQZVRWQ8S3
wJU+m9LJUcehHQIIUmnDp7sHKpG1sR2hpvpjMMlKE2eK0Thf54ojxokCCZC6zoSo
e61rQP68NqKXJ7PVVJAlbQrNllz8WM3+z9t1DPPcNLbVP693haEt+aYvG5zToqNZ
2f2BTdER/RKHcCRmif0cVqJZKAktZsUzn1xrPmssPTtL4lkvZQ1/SuxxfI+xkzan
isIV/2+kpaPiuGmch28hdnFif270TnpuJQobZlpQYbB5RdO26mHOeysSPhv72u2i
hC4vaqJ9aauRl49lOWqZMAVUKcrdTt1/fBF9UiT1UeFBGXFv3OF1YluANwRHj7FH
eTypT2Q/3BuM7DdvUCmYkihGQoZ6RP3KSADEl8oBZ8BBocEtb5PykD3ZVgfmWRas
6tUr27eO5KiKxWZH6Inf6gLBn3BbUui/ZBz8PUGQGyn5APYW3LY3IOlF6U+v5xlb
3So9iLJsZ8AJVyvqjOxbqglsozFiWvBugYljO1UP588WWmGAxHbytuimpmcfYK7p
03NbWT5usPJjt4pMwD+SOgr64/Fa+r0sv1FQIwOcww5kKw+PGDU14M81KQcjZJSR
uSSOUDg+a4chwJYemEca7iM/JptHwFhTrQO+u08yuIUpAL1xtMjKrBt6sWpKX06z
4lbbzh5DianyI012Bvn0IffO9hM94fmwS7zBr4gD/5DARF7Me6quUOydETmbEALQ
aRptWQKHxCXXUipUtQLYlP+oihKa034jOWv1kVwdu9qvqRsSDA966kbIFqH6GfRE
oruhGZtHyRnV6aT2GRK3Mg6wRkzFUKBFTqUK08TJvylB5W0ogb1akgkyBp1pLVTG
umo4nMIx6U3KIU4Pw2ieB8tRcOMupHJ4Hf1KI+wlJ+f2dywiYlWinxClR6FkxPm4
HU88SKK3U22eHmc7mvTgThxFsIjCLdj7XS7tY/X6rx/kG2eNvQUckM/braojejyA
vpQJLg4j+RIOvRGiCaG5VSBgXFzvCFwVY8y5ipycbq9lroY2W+eyXDkeO/tfpTJQ
RQkpsmaYUo00PyhbAk6iHLPA7eYog4UFPi6PgSILiqhJPskNRhcbJcCAF4JqkSfQ
YXo6GE5U1qx9Xm9iiy23k5LmLudlSNoBa7CsPmtZonnVibNsF3keT0+VREr2ZO7f
UVWBsEczjoA8AG0ILN3zHwEJvIM4V5MprTQqeLbZ9Jq+Al5cjsSCeYq9LJlB1Dad
ADIlWSiFJNbBnAiZ/V32EOSPdYDjeAJwcEb9WGPP6jDkPkVtiXAPXLiRAV4KtlEz
wBja1ZTduQdjwsU0a4+iz6T2IjDvnHCAjT7BBSywophfAqoC2jiAzM1M9KzGBZT+
9UWEs08Xe8tXMIi898QidIviEgQGQrIBmrrmGprGbW+frGhA1ilmWxJkgc1pTO8k
ymWI0sHsq0IAx1DQJmnqyFIm18B0HBVZ5aDpvINDR52w72Zva2vwh+zowPduIkEK
3LDigBGGe2z/GI5FlYT3S9vsIxYgiW8pNpMUm+hztEsTNn9SnPl6ltyp4ZuC7j9t
2EM/qKB6Xbnw0CsOp6V+C8kN+SPKV1SiEtrEn/DitMfw2BpWw+o5epLQ4QhB7tiD
bZQhOrFc5c+qN2qdOfHNl7VgWmpDS5uzjsa1oJYtsFwOK0b0G3uOk/EhqJJ8qYIU
G7Ql6r+Z+qsKRF765sPr+fTB1tbVYxqOdbyq8h10hjuHk71ZGmy/ohOXS0uj7xFO
DzR/smhkxZX8n8lqZm4DTmzPEI6R7eN1qvwIRgJ+cGKz0qfiE7v7YCEJdtmN3+ti
Q5S2Hp+IJ6AncSkxNDAmZBZ3eORtKeNesCh/jGDexdnI5pqGo29VYS/pOHJGzusy
RtnrdX+8Nz7oq+t17Md6QTp/nRNIcXGGijOroj7ZrV+z8cQcVDT6wRGuvqUHyPBF
cTMNSZEQ+sfe0VHTteDkFRwofXGtnVsQMO0PKjWm4nCvMrArTzzGpXvQJ9JKaTcN
JxDhdCFpPz8zaP6a23hdAZGe+e8+hzH9Oz+O6UY/2Q6lLbQvvfvRwlm+MnmjWmUp
vGkkisCKX7jZ5pciYenALqWcc5JPZIOT4XewW2uV+JcYKsSukRkyTgj88mLI/94O
Bd5Q9wR8+Yah7f/0ow/noBysMwQQhZjed9Z11uovkrNJNV3DbyKgKQVh1151251M
83Y4s6OP2NDGxWxCj4/L6i+CfzbjTIfpelMN7nW/2AiKiPaxuWNuawsZYkqpDxUr
Xrjy/aSq5Oxv67K+jQP0bRYJaoaxb4627TCy3t4WL3f2+wuxDS74674LvP/Od9Df
zogk2crP3evc1s6w1kCuaYBxi8umGIay/Ospq0HQ9IxuMjUMd/+6LQSIJ1QG0520
zg5WUZGzqefcD7EnvalImWw4eglzouIYDKiDQHJofftIhMUFHbISgmcp7w1yivbM
R7rRu4/HaM4zg8/iE9IdbURaauBnO5ZfjgGSRkGPMCrdoqIqXqoEmfi8Vc5h+Cbo
L9vPWI8hyXrZ9hzyjW2PsR8Aujfpo0JnNOnLJSwp+Ps0rEVqzr7NAJ/Yp2l3sJuZ
9aaG17gwpF4BLy/wqq7N4+lyYJbccn4TtGYzkqPAi6kWQ1H8JR/9upEP40MJrz0f
MQo9Bw7JhEJRpIoXBSQR0tKqzMuuZoOurwD2TYtO59/lDvvJ4QEO1xbDjGwHLLBF
FI7+mpdHpLaiOcjYszURqX2XkgUyf7jvw5/ZSLSyL4mn9AH/8mACmSeFmT0Q9Pi3
FnZ949Ade5c+9bp15TLKzb6mqkGG1LgSZ4YaEcbP+891I7duMpH78wGqXa7DIdrn
vtGKZgmkI8Qc9dYaHPaF5ymDB2mCGQOv+lMhZDzBvG5KyAqyi+p75RwAEULiIZpd
LkOJrJraNd4ou2xgliEcEa9h/Io7j/WY6rL4C7wFRjaznLdD5sTSjegjvrUGqepD
zgyJ9NJ7aa6XUQJA9xzXa6LGeOcVOHxT6p89B8DvVR4rWKMfGH/9R/QU2BEpb6p9
EV8FYDFFNfQxKt8Vb+4VBTxiSUk1IGG3L4xlYezReuk03tqYWGH4vf2++5XX/MYH
m3QE+LuGgnqT2PGJaiCPfDDYX+4gIU9BAaG6WxUAjA2y3bTmZvkYKmCDcewUdnhT
wq2mrA0YJq0zsD+b4DIYm9gO/8+TZL51CgsCP12HWm5lntTZly8UcfamqUCBxFwG
/gqdms3T5b56oZpzWDLFdpGf83ZvnQH1VfmMi8Vfk9EiO19wzFmkYzvirbCkBc6d
YD5iRVSh0QZZPWlSaP1XeOl8aAX9PjdR1BmPDvAPw1Pms/NVgPR992DPJ7G0OQ35
RtPdS3xsHzCQG26hrQSws3cKWvI0MxWS5JtR9VP9FsBY14AOhWI7eXim11n7HSq6
x9rp/8MuUz0NMYJ1j2RlmdABHsXTsiHxRLVeqIO3NysGITQ6cEmsZ3WWRtJE8K7G
3joC5qan5dITjgBdDcT7JzN+IQM51TR0rlIOMncyiL++kWd6DJVMSzQnHORhV3fY
zsrgLIBbyfVDCvo9FPzp6xibRW6IYrDDbRLEmfCr/KHYsjvw8vDb5I17wAysDRMp
mcTuxbm8KaBtLhfedB+QZ2M1aSCr4qldLxtphlpoWraHbkJThjrnG7oMVx3zMtKs
eRqZO234DJuJqg4gvmn6ubLDE9qAM0An+/mIaeU77LNywXkcRWNRlnv6kZPvyFZ4
sa6l/pakUEgsXSdWH1EXZviqwsdc1/R4OCGx+mkSGyjYRAPSRjT7tAWyagnBcXXn
xjbSAAilwJxP63HY1BOp1t3LJ3G7YQkGYGnotDDgwvfpxjCxlqY66E3CfvQvDHLy
Vv20VM5NHugkzs4SDffWMl9s3P+onPJ4fJacn6Ws+rnB7nAkL+V+qc6ZAppBGfom
+Ydkm7w8FyqW9hxVHv4tRUSaOWYbDfTcVFYRfs81/2eRY+imDDTBbDKJ/6hTjTre
BEivUw9VNibL7nIRtGoEfko9IwjAZeUiliRW7SmpBnuj7lDtNen9yv9U+7wD5es4
fxBKHmtKC0vP9yAVTR4I4pnUAAkbDzRf6zZOAi4pMYaOHx8fLxWZOQv3ly8n8JMw
6LI7eJBeMfUxVEDtLAO6vd0+VQZpGNwZ+3TMXa3DmLUOBqvYv/F5JXFwL0QS/9Ta
PNEClLF7rFdX2DsY2qvzmsI91vixWL1kUS2RrDp+bpxdTXBpzztYM77bnxLK/Wxt
rl43mkhjxaNfT0zIDzNMq6/y41Lg4JQ12PXOjcBF+91IiPMVj5akdRgNzwU0oukZ
8F9/3xw3aNn3ZamSq+RIdXF6IxU67lVQrZJrb0dlmPGvQamxAcQy8SEUEBL3+H4a
sKFNAJCmbsn9I0f6V1hOX0Sd3UC3KqcBWnCidxrPLkX12pQt2ZsFXWkTRKyWzkWN
/F1xuKelsaUb7jduvVA0+z1uZbCxatlRWLtkx+cH4COau86ZY1TGx6yd2Um3FNP5
DKMJIl1HdtTn07b1/in0oNBUGjKLFY5artCqjobMNHO2CywsrlN+l+ezYDCPz2q0
Y5KGSVAdBVT94F+SRvJg3cCJB8H+V9bhVOrZMyfN1g6blOrhwoHoLfsbMwbWU/XE
nPwBww4X9v6ckygt6IJX5egEDqSyGFn8pYxu8ujTIoavJJYPBIoCiQRclyDex9Zf
X/TIgoJfOXbIBJMRwm8tWgDBrOxPSsCRTeSLxmqC8XkaGIvNmCEiacW480VZGL2R
+d34Q3EJABsd4Cx0Ar02dQ240jFQXYhs63/Q+8vfOACcjCEsOksc64+sTtGwN0qn
SzYf2l9lNaP+vmz++vIHn3Xro59TY8Kkg/ICTNR933pAhpBCzLmjsjwjDrtzvAuF
/VWkxo5lf0nIR3w8fpjIw59p/j13OSrKMpvX7DHYJqiolficuPWYtR2Cv8fi8Kko
95lxL2gHtOxMt7scowgw4MYc9leZ+N6BDdYTBElouO9GZ70QUL4HhzHdCXTFXV3p
QHr5yRDPl3qSS2jO/um3jqcvSQ0xlIjt101H3HnsZzt/qXfE2jSBThQIABrXlhEV
YwAqCYrAe98uYUrC8VGbHdLNh51Jw9Qo2YAoUATSmmluidRuu4kBjt01sL2bX/ux
DQJXM8LkKnN3yaZpjdz+3nOAeZ714k0yN1EuxaBiULFD8XoKwrZV1OYEXdC1yVSO
gwdd2Xok9cHAgwBNOut3JDZHLToTprMQk3roWQuezW59RdDRw5E0YqDe78JIjPIk
Rc6zfZd2f10Ku4IUR05b6/W45oj9G2sU2Z1Dq/a54qcbDRy/uI6ADVDEPUkl6/AA
B8N5fbznKshnkN0sHsZs8117QHE/fsiYVm7Ksgps8coeHnZbWuwdLMyjaknINcY8
kr1AGf8AdaNoEqasJRBVQJaDNIn527Jtxx3k2XHJzacgDsYA6sexyEa9MKLTThn3
xPaCuBzMUFjSGk8gH8bgiicQnSqYc2rYCyB8o5srS8u1oSHl1f8j7shLgKyprXkB
MRGxceGMotK5Kt0Z+11Gm0Zdlawyy3pO6jQIuqADEYCOX8R4UDj+fn4vFAcjukO3
D2A4e/dFz7esaL8n9uOnBWaSVp8if/nkyJJYVkBana55uYgt6F+rJvaDDHY/bvPT
HxeHHvqCeh/X27HAu29D4plOAI8SU10PrLfz+o/RutRZpz2R4Ah4yz0/VwhAiBhQ
zXfnWEylkjaSahuPjovKJO0DUhg1KFPfzw7AIqLV3ewvig+KqOQ6rCchtS4MYKWz
ts6ecY1peEa+tH9Yu0XgIteAWlplVRvJlctzJ8khBiNOGtJlVixM0n2ctLaEPptc
8as7DTV6BQ/riKQ15sMtoFvBazTDZzGSgKL/9kpUwqvrHr3V4QbG0hR9ekKjWX/6
pV2dBHQ2RyV+arQ5P0kaHUPI1a6bLbN/rzQaiMUVBnNb8pPVlKNr8VqPH4CkUkes
87oEfps2U4LRG/DaV7/FI0VWyEfjMv5mBaRLomwC2hSRQtux+1slVgEynGPzfKaY
GwDkTxYehn7sZHtltY39jg4bSHkvZVblUOb9OuTiW6WEQEUoJVHXaNYf2M3p0R1X
2YjSY5bf3wC3P7LBlYOjmR0Ow/ksIGJ/T74MGHOQBatDRXRvgjf0/GKLizcr2lwc
RNvEPov+PPYpSQDtoTHcQkv5xAm6QqbntPSfHqfcUMVsiTxvtawKH6I8JpuVlCkB
C+UhLcuMt0xyvdNLKBFucxrIrgHmmiaPxgmHWm3FOXXr4G8bn3N2SyY6O0MgrfWE
nSYqfnzLJ8d2NWfM7jCzYLUA7o++EIV33bw8t7wX92dlOZ7Qu1QX+6j3e+p1IHLu
T0runGipe5bbxxiqGZTcptEk08CAMA9k/LifgeyoFpyjVNM73i+0y1uDWK91zXjx
A4Iz3cihhvnyJ0XUIiYeuLzhjIVpjjDUVOBzgg33bztbTrwRlGOII78X5GTIzLJb
S5vMjrXRyj2L3qg2b5oOz2Mukgz3gCRaBiyWwVUnpuaABZM6fyzkjBTnL05o9jgr
xTifzno8vClM+SDSQ+pDndXOiOyoR8pqENKhzV/ejLoyBqMCE5ORWhcs32Hdf1Mz
DTL3S5wk2k1S8y8j+fYS2DfKUxmqNZv0q7IqgpqftyDqC2lczgnmGbaty3nkAfdY
stEXGT5gv3zIKJ1/QbonHYljwSGtRvrYU2nu+NLrAAf29Urw5dfnLL9PnQfgS4wq
i4vzlh59TzRtjY0bsGon5CYxQ57vnNQNUc5QKzt4NvATPhtH77Kf8quVMHXWkAFP
230SOOWzwrbS3BKYTRclYZY5mQzD8RcKDgPfsx5dfUleFHw4EwyRGnC7q75s17WV
KUmT4tJua/cq+fpk4nHRuKlHmXIYzMTgcSwqOntRUsoqILyRgvR9QT6ziYJqkiS8
EFk7ZNX8t+z26WshBQbxcG2OsvIdau7fS+rVJqwauQLZEGOcpxS9pXuJWjmcU0eu
/aBbL1T7S9H0ZAFhyYs1NNsyYJckPVJ667tA/YiXvKoXrFQabhn6Q7TSMx/KHrgw
Xu5rXBjmXKMkG1HZtuLkLCVWleU2tDUfkyLmSrBY7VVZWyG5nRg39+OOZ4Dywy4Y
FlIvzRGSajgmNjlZPO4+YYw9MlqugbpB0rM5SawBblrn3yCZxk8uvnikkBS+b8RD
7nbxmgxRV4ktfUNz+ZXjoXOKHhG9c1IxS2vUARa9vhur20O1mEGzBdBMUNcpOrd+
z63yAwT+OGEOM0E8WYLOyxfU/xxnoHSBXYGTg7HDXqUD/DKyouhpOtISK8NyZACS
Qx5hhl0y84M+g24pWaICrIMTMijRBt4jECEiyI4GMwxCn6KPCY1xhjolsYByt9zE
ERsFzGGazXbbwCkcugA30lY1eBaiuBw55rxiTLcuIcDIRnP3Ssr8EyUVoikVo2Mf
8QfiCP1VvbF3xFEB744TY4ZMWtkv5O32evLgez3u7n2genJj2o49wiWZpQF9I4XH
XeoWY3oNDVO4AsH1hlX/gBL5iNAX09H9OTuD5K1kY2v4XnMnDotA1UawY3GXa2cg
myxb42RcqQ0D1NrPLumaGEe2bQTbH9nhtrkVdfPlxWl3r7AKK1nHnRY7UrYsS7Hn
qePv75gL2FO0jG3XB3yw3u2/5jhX31XCYQEafsk/RtLFqN4kzEoFNtjOajixxkJY
wl0LeRHebpW3Yl24a6SIOFoZH7z6cFT7K/JvsnotCUhrVGL0ag1Ek7tGFVo1d5tx
ETRZwtr8isg/1oYx6WCVSzf5fY5Bo/lh6QzXc7sbbNFDxX7KTPqImFYGkKCtgNDb
G6sBQmDE0GcHW4Ukp4scnO9NUI5aY69xK7D0ygSGO5aOoLHc0kMz7WA0rmgkINKo
5M2xqOAUXpe9EJiMnI5LEn8zPfNh+ceJ3hsLhViQQlTzddPjrJsC4CfcfpeOgkf3
ehK3liQY1xf9AJHl2XuBZJgegAqrNWg81VkarMBRxD1QiNAOHrDLvBBSFyuX1f7x
ifh8/x8RAHgr9qa/ofylwOPAkQcgym53C0htiCDul9TmTJE4BfVp01tsPEbMZsiR
sCTvsjNeNYQnFMHmqh6ni1IPtpJxd0K5J1FoxJKIXsDY6RZ/RfdxV5SqsYML+uGg
y7cgLyhG5riOZ9SFm9TJ3mKnT/vr6ELj6F2e14A4WMHdZKSoq8DTkXnMefdU/94y
7+Xn8lzhsXE41bYR8fMkTobhpEkrFIV2z9iev81EzwJaTolZ6FjyFzCZnG5kpGpK
ye/GnDkDatEwpoe0kX7QaqGgaOnQZwoAJPedvxY3M4MdM8H7d11uRE0oIz5Q2ZjI
H86nK1gNKLiXS5hrBlAXfdX2Zdx5+Qt3DLO1jS3Sbo0/F+F5bEsSLgv7MF72o9tq
jg6l4/80qc8CAvSGN2DUwpcd/OnyH/okLHBNKnIR7mPlxNA96NS/btT1mL6gKZTP
ZKFQdRQTODYKhyA6DfSFXLyMIQCwM3KVtwnqTB6+Od3h5k/EIuzq7yLk5kiBC0FM
xX2XgT2MW1wsv3SaskbnRUUKI7EokgPFUhRpH7kocRBY8hQAkCr5iqiSAu5ll52P
/LqkESvMJdRcs4PUe0zEOcF+o4IvQwWp5lT9aWvmDWidzo9Smahma6gF2+DIYNey
u93PxPOS26tFn0dPr/2UCgweWgE0dOBrkDvh9agZdfJcWMW0fKtk+pH2JwqZuB2A
9KwDF3M+UykmVTLe3Q9Jhivqr/4FiudTH0glF+3hx2qIKLukviOac803zsrhJO60
Ygwvx2QTCOSf34j5FOpVVMuOstr45CiQ+cPY/uWi08kumdfKCWFY5BKckaYZVshD
8Kjymek9+DWMu2xuJXUbp/CpOm34+kfBG7uf05Ut8yTpMSnMEt9CJZvKPCS747o7
Fz9XFAVHsvq5PDXwA2mzUgonQvb0mhHOWCGDI6MgsRHhf10XkdvGiFpyZyYtrHUp
4P/OskRGFESqrl4BKoc/lQaQ3w+TJ/RAGo0GqoQidBwKjV7/jK363zFO7+QETR4w
y/B1vc9IlXfr+cRdIYe4R9v5YRB5+Ro3SHHVgEuQmJx4RAd5DKcZPbtzN+sNCCis
2HTFqaQuHKzR8ER0xwBWaWb8CdWKGTJssWDN85EB+D39QT7D7E/8OVSrXsrttJJC
BEh75QP3T+x2Ts2t2frJdCzc1TECdCGq48LBvLmfrkD7DsOqTqGE6mu+EgxQSjuk
Gaqmi06Z0byitxqLMlRef9/SsXvPuE/WWusf5DOUTezpS4nNNdqmhGtZqxX4EQVl
wep7GQZSrvSLqaGtTEP+A3Hv6xQS3sqhDCOS5pSScVMm+aIu3waicNEMmxDiwOkJ
dvZmMEfb1jJkulFSmTYYzzMJtEvNTRzcLDMh0uOdhOpeXuzaeaCv7WQsbb+NBQrG
7l9mHKDpe6v3phul5HzGqSPygAOn1wj4HsUZeTciAl/N+bVRvrX9eAbgrA+dKeB0
ZUh4hgaD12SN2rXF0bevmiH3WlAnvU323Zrwye5G+rkTsCcG0UTe8AkwWK9KkDYI
9I6U3hO9tDXA2YjvjSYdSjiJ17/BUTeTnUaZ6lqB2dDF3zRv7AO8hMiCg6hELFfA
2KIQwYjOVGXpDmhMBwqOQsLBpCquOhf2RcIk3LqVX9GocZvoNk1+iLNUg0kO1zGt
oYnsjBlUYbw7vUOJq6Nl3A==
`pragma protect end_protected
