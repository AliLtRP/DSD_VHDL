// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:08 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bKkNo32vxvbIp/REyO4InIvgyLt9xdFtm77pyLQweLv3cYOwv59TpPbsyD7GgJ9W
6WvGvAvTS7NbQch5SxaRpQSrdiZE92Q9cZ/sL9ZsrIhFdl8Q1IP5kXg1rgoKPD5C
zpGlvBB1qW+zTfSLPx/1+74VsLbwE2ZbasXpop4M9Jc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32976)
2VPoaa0uK43e/8RJC4bN+Xw90t2kVzo0zLaeF+1eSdhqetshbTi6PA5Lknh3auzR
P9/kv8Bb+llsljmM8ZPejceoHN7GCKtYlEBvGEaUY+S1WxnFyfvQ/A2LbINBQ1pM
qyVr4N1w7CMaqqgG70zfmCXDIbyWy0UroKaaA3loxTuJwgm2iMwRFecUqav6wIfq
PKDi39vyIr7hbFLwqQGSI/PdeZ9YhvbjGuM8aUILv98jaTfwX+6t+F/QgfUFSCNK
hs4O7DrL/6+PnWhFISsb/fNL9aWB9HfFGTlS3GkCki1JdJPcTZuW866SJP1rsCTb
LJOb6rM7xJs3T5qGBQGmsga6XlqVX3h+YLVCUnL00KgqSNuwIvGG0aYu8/OEBNje
ZMHG+tPwSzR344t6ACFmbQFywWWMWrBA6KxBhmSjBA/h123fOW9/2beY8YPAldQl
xJeQ1TenIJl1ydh6Q9/SUrEZpfkP+XsuFyrPjp+xiKz3croM9LuseEgjofDfw8I7
dXF4yykV7j7ewyyg24IPrOSJjcVRjOe4avdIXJsNVHK/j3obLayk2rMAkHFBD7b4
SpBG2TrlzIxTMXmZqwwQiX4Am8bYUY59x6A/8QlyxhXbUl67Pm4+Ni5tP9t2djK4
W+ajP1HsUQKv01jFJ3wNUMDZOMrL3yPNnNFtw71zvgUcaQLPLVLpqSldTqLMPSec
j5QZoMmCK13zMqFNtE6sjJtO1NEQJoBFeK5UVgFOQ8D3P+YoURLBaEFndH6wqnvw
gAzllpbT/7VGMpBhvAo7aOX3KCEwwGvdPGitd9Acjq3317x+j/Rhth9b0/8oAxPY
4DZf7Z3pm9xnd33RUbGy36IRvni+t3Y85tG7f2jGRrp6EHyodZfIJo3nvrEivdV0
MJvAc8ugLtTPujsEqhHSFcUS+9CXOcdSIW2crsxJ9RUnvndsPAikw5u7D51a+Xbu
rbgqysAsfE/4h0zyfi2fXZiwKffxoiBvMFCcV/BRRX+Dc5Y/8T99TF5ulg6PWeJY
QOE6iNq0x4fPssEHy/k+6vcledMIx1uHy1izpcwh5l9jtIq2MOaJhfNXSnNqGXg5
n09MTzuaICuScInGi2nD2UXV88UVdP/oWRIcwm9qLRd5mjxKsf/mBbB2EufGzZJE
/w3czls17LY0u6b7OE2qDGZEePQsEkDwVevu5+4zPJDjdV65Y6XChR7fPxIPTwLw
laZpQVDlDeej6JJNGe+AkANuiii3x3e4dYWtPv9xLqYZBbJ1g8xgw0UFZedn464u
bN1FKq4DvEGUJdPJHA4WNmCB921PXQSVLYB74acanriiQ2CvEzycHRdQNWjqk4Qs
xODQ5EQZh2En8f3dmhr7LCqJgYcoN5zGRZlMzZ6IWZ72y0NugjJg6xwONR0XV2us
H18hLT4N9j8PkTR2I1ufeElV1X26g4YjbySvnrYFEsWFvXPmp/3umlo9J4GRiOHE
pRtS2ADSNt00cYG8GXR8Ln7ewThXQTGbp39Fsbby1hMcvh9wNVM2/VbMIAu4Fwb1
XLXFcjJGX9ZVFS2I2D84JSmuWNZ5+wBo0RQmJQxnDGfruyvKBPGuT5w2103mp8qC
cXZyqCXkRofyTe0uQ0BqB/Fb5pjoEuuEOiQHl9Bq4/NU3+qBr+O964flIooQuShH
/eradbc6X6RmF8PiRETUSY+d8CvhyzZKcwhSkxx/jvAuqGLiPW883gR2UyR6h9d/
tC5ljvKDCA9jUZHNEDY/t1G3QmmSP+dBTkQspQX4my9eOd8UK25Tg10yjZsZ/urb
mAlQvV5vEy3f04WepCP8bljA/3DogxUcuUKSuKZ0EEEz7Fp6TOIksG6aBzmt2yoG
PbWX1frQhuIlgOi6C2CMVvwDvh+8Y7vY0CGsBE03JSH8xXI7oEGchDieXqF6W6Pt
HbfoPC74QddDjURMYoX7tOhLlvx94armEZjc6+vliYRVLnPMjrMuxEAFwKcQJpov
US3FVTfMR+PfTd/aXgpQL1B6irtF4Lh1ni3n7EfkkRa2DMG5j7yGmmKHt9MwGEsc
HWc8dSM36k6SYIAiwJVeFvFw8mINIA0KSdccjwIt7Yeo9iyea7om4LKFIkMlOfH3
OiYgiMDPm7Qk7u7eoRJnzFb6zfjO3pdbkTUE05suPdQX1T6WWuujFu/R6YDW7JbO
X3Fe8HGGsmmTn+M1HHFWvykPKarcs1Q7IcCP9Ks75ykO28YfZ6rbKLGqoweGZelZ
1/xtVGZTY7umWhHQ5TyqLi6/RFaFg1RWC9E7u9XABVYspNBLiMBSHvZS9Q9xBC4s
yUT4dRD1guSfLm7RDUyv9//erRbGqf5wdLYcnUNA1DfsyzGsxOdm9au5h0AJdhjs
HD8Z1dAdVMVLrMztlnkGcbhsMBwq66RqMQ58fAdA7MVsaYmYP5EUvqO2eGJ1k0SB
fiBoigKV9ztLt0OX8YSQRHPREEiWb3OfT90BdEY1dBJq15vYQ7X3cvqbO1azRTLs
YHIXHFSjW79MACK1XOcRYerwkT3b0P7F7fU8iV2KFmzQXpKiltYDn+HLHP7A+kBp
gXKAT8IKd2FZU7mPFSisf+cbJ5Apkyd5hQPQNr3TtMIy44GJQ96UtI3r/8QP0hyo
OaxJDBm+6FWxb8jvPJ7QU0e5yfLAnq6xv9+d4PuJQ0l7dZVMOo4zcZ7hOUPJJ+tF
3BKyV+AXNfQRBiNOmvc5RTbI3CnqZgH3j+fA8H3+E09lT24oslM5dVEbArqLJPnj
xoE7XJADL8KRtKpJ/SbJFGkkIL8dsV99kpBsSbYaopgwPhorjsMkvWXEfSjp5Rxz
WYPh49YQjx1MtVZd+vp/hC9agg2teFNuqhyd+WSAvESds0vNM42KrFxumLB5Le7i
OTW7Qd7WlNtnrKzwWvqzbnAUWhCpMQOFHxvJN4APMVGzHzU/JIxf7g9eEKM0pE3w
SzPBn3U2LkCLqjLHmNyv7QDXb+Kvz7TNnZW9+saAdFBg2zP7UTTfavtThpy/tBb8
KwyE5DSvRatCq52eT4UfpeBjhGS9DkemGfkqlgtEdrVBElbSJXKt+L6oMum8DLG8
vpUHHzJ+bcbcwIVFPEBzyMp3dal/hMkInM0CUF62HTJNW6hplnoU46wcacK/5Jfz
gAo+lZ3X/gKmp0s3y21rsMj85+CCs+rYIswag6YLjsquum5GOGj1zodvGxAsECT7
x6FpVb7zeoOlq9pbfhlHGVcvlfb5n6LPL1WAP2YfEa8mb3FopG/KBiq77bypaZ6v
g0ga/UEljG2FxrktL+jJ+SU9ySzgalMES7dukc7R0/ejUjCIFxRkjUUxxJDrsdd2
mWHfN1u706zshIhXPpynXveLdoSHk4z4FRqAzj1sEjRC2qqaffQ8ljD2J5vD9wNy
/j6tl0lT5hcCArDeEKJwu6vqXcPB1+NTbQoscutQGtn+1QUafszNWTU7nfx5p9ci
DE702ABWXC3maYFp5ucI+hlTU/2x2MFvJ5o77D5pP7gKMBILAutJvQU+3QtjeMCw
yehbgI4ziHZwSwMohsAK6agK22jGPNgppVCHx65jQ6+Du0ZiZq41vv/lrogYjF/K
2s3i+TGPzOA9uN78dStsJ1jWTldRzG/U3URD+pe3EggBWO2nKpC+FOsm5Zkvhh/o
wLYWGhQrPdXy2F9FVcN13c8jjbiHe57cob9c3hDq87p4T5VaL/X1Q+Hk5pPsP0R7
OxKlK2Yoz3p1BZIJ7/BJdQ3rXnaaz4LLJvlc5FtlyY0iOHWArenNXpAH+pAQpqkT
4LxWYqHOX1tiMzfZB5Zut1x2lvTolnTmkq3lEhEHoepMUJAOVwwyUe1jGG99Vh2V
zPgJMNzofewG7BQM6Y6QOlARzrZHdNIcR+c/AhCuYkRjgu9a+su7dylHceymquEB
m4fHzYBjNjHDTBm/iDXEjG9nfW1SwZwTMpiqbj8caQyFusieNcc60bQWjCIAzBOI
0shYRB+SNn6etwLWaORYllTcx+pckt+EaRdaKYCuEyw8dH4jmLHN8BKQJAWAYqU2
di0X45e/7WKcHa3okSz+grMvYOpEHR7sLtlU0PBvmme6COehKDeHUZwsuIFbW+Gp
DmqNjsWQDtrVxh8ZgtbfqOgL4eIYMA3MhYuu/CoX1BbpyyMHmWlBaE99Hfc/MRrA
y+r4huDc+ZqIq4MNL0xNejwu7csMtaUqRYLyCiwBDoqsa5FbmFSGGwUHhahOZepB
iKPRjhiBCxI+ocu23jGHfVmbSxqHb8aIkJ0YunbzWK4vcy6dijjUW1sppNynaXcO
tXSVwTrrKuVjzqabaZ0F4T17dAVFTkAgOsQ7nDnODcTXIPo97Pyus72g5RXsu24x
2CpAgGz/uObsJe1rDSvRBYxdNRGsBh7yyNCt4EgfeMXgz36ioHQSiyIw0Zx4JK6c
k+lNyhJmqcinFy/AuVd0zoL3YSzoAGpJjJeJnX2GdZUyZU+gAeyhTmkpy7zIYLBD
wQ955PHoHPxn0zmBxWUWw/VstrnxNxzBuCHk841yikNpJJLGuFJ5MUaucOCZMuUf
1fr4AxIrAWwV91HYyinsn2Vg4ut9VzTArJJWBWBNpN8K++/IX8jYAbqXUyRu+BU7
WN/J4OYibBzWXgYZtL3S2s9qw/Z+ezHsqYA5wpi9FnJTy0smFsrK0xmmH1hsvGBB
wip9Yct5KrIfYOV5w5Vn90xehMRK6YpyLEWSH7WhMQTOYurcIU8L80yuFt4z8lJO
+RVGMA554p9YwUwCaff/Z6czpDXdmR9IklVcMph9Ng+rjAPYPOMAdns1r5pKYKi6
5zFdo9QWvU6jll0jFgH/p03SBU/3tOeHE4z+3aFR71tiCoxRtqG06JT3JRvbtAe8
W8ap/1NFgYk0VqcqoHXaqG3kwLZxMYRTwunEA/wtCMndquCuyVnS104PMYlu1zzL
elowDDRVarkNUAFkc/7Ze7CzLSke8K3L0W0Y9CXOSNSmgsXQZzrdinZJBOGT8aF2
AGfXGExdO2cJAoyVkb/5MRe6YDACaSKTYuKRzdkQASe5rRQ22UKDrIHNgiAgGlSe
d6xzqkE4LK6b/Lt0q04I6XypcQuyGGogJ1Fw3vYFtiuvpfoNwzES/PRxUU6JWx66
+rm3kbK3VF/ecwNJ0rrS/OLwBDMxCp6SRpY8gG5ykgtKDGbRiGmbBsXY6JQ7n18M
wB+/RWLB4SY5QDMxtuOG5KiyE62Fbkw4xI2yn5Uqxwd/PmJV5dHouVN3StykrhMX
VLt5rpFalCFtVzE0M+mxWo+G9CCf2js+wU3nU1Ziw6uotGAN5vBJlP7M7JoULh8w
5BjhR0rrd9XNDOuOfo09B/C/TsOJ+BGwjmibM/Ku/RHNMA7qPArB0RZEf/osTdvv
p+pG0oVdfsVVJK+ZHkh0x9N1x+0lSQtuRkZKmn6Gp/byN9Qg5a1/gOgUxlj7mQsS
N6aZ2b1noTpci4UGneMdliLeGbbLuu/ZgDRvybYhh8yiamKtWbxauDtD8q6aMYyT
ZJnGZYbALlIDvzKn7C8+AU9qgTZCtqHO9FFKIrtS07wMuvHZ4xGJ1KWRG7HgG3YF
G3CuH6a+ylwrQrtbJHVmIVxi/vTmopxBj2NSYPIRMAVdKOVwU72llys5ihpXxOv9
Xw+PUyWPJqsRo0djuDspD3XYCFK9wqhRcABPLt+6l6nfqFIWsdK6i7vavoYbbdCF
Xj8mK6xuft/fD/gYUkZ/SLVy8WGSLEdNo7xmAYU2bhJRrgX0P/RGEuIHTgbmG+9V
Xy29RGmI1hb+OgK6WmMAT4P51QxwVsEzqNr/db6ZlA71tR8vlAiJXdrPVZSoXFqg
RQv3XfkFL+TO9JArqGXTtmeTZg0I5fLKC+io80jZYzpIlTTYStH40dLTS9ow1kZ0
ibpwXT+hgm+tCZt3fKOesZ0l+J8J8n+BPfwSrIgXjlqiuC4nm13Ym26VAVpyxUU8
Ln551QnPjc08Tki+GGwTlPPaBzJk10LkA8j0XYakUlZFd+BwZfolTS0SqARpUTpr
pm8ZEmILwEn1+sKlshQXYlAmV2RmDxg56+yEtJ9D06cjF7ZP/jdCCNjc/UPriE8e
FItaYku1LUKjldEa6rgdbO1Evo2vV6dIxGXbORaLP/L0O9Jxou55B63AMpbroXcj
D7krO74hdkB0id+qV8XWOLZGzO4ZPy9Uz+e4KDQb4/dYzQPxKXMHQIulNhxsOpL5
jmoevT9lGBXglVlB/yuOEQ2v38tSM9RSIbQX3tX/zu/6K+w8Nor2WwmExo5kFkow
l/XOsSQpNA3bKZRRqkquc0Hvha9XlPxXPwvX309D3mfdKrBM+ONIdyOUj+SZsQoE
K/ZIVKqWeRzTId2xgBWjxWy2qI+8NjIaCJ02lB2V0K2HyrsQZTn/9lJ9IH0JQ9fv
rn340Kvf5h/24cxe338x38TtbCuMzaqSWKgiVjRp2n2Cenn33Iz6s8HwZ5mk/rOy
rt0pBlkQYRPdx9yl5BZNM5mb0cctoNNm5kmFCNUwVe/FrCyngViKosXl6rrkrr0L
kp62DyMoAxyH88LsESpPI8DD2KP9KIbFldbCUGP1Rqz5wAtFiilrFaJXSY4JkTwT
oRHaFEd8f7k3QQC/S0xHQusvZ3lzwsDZkr0FjaHWybL6cHhQQmbR+BHvkZHVpEBX
wkvWsBzv+VKnfVowhKZVmD9R+mNCwNNQ/epRI6LgNGAJ/6wtPE7LzL7PK6Zc6Yal
vuAwiJnqTD2MAAD0GJ+NALXbnwvPLblMUmfOpLQV1K6cfcK73k23lfU5zTr7M2uf
0FRxo4WubSGIqGX5FV6rMzkg02ICcAjqEg5BdJWXVhqkJZ8RtZH/K8DaXxor628P
uY3h+tYEqwjl8R9S1GQGYe9cqzK0Syrx8EMeAymNlJY8wlD5wSbCVE8jgupWWWWY
VCZLpUGZwf33g5janDz4aq0f9KKGRlJo92b9RKw2pd93ciZrxiRtNDRVnfStbm+E
t7FWE8VBHsyeoKZKRDluFk7NVFHrKk1Tcvmzuv4X1BZm5oskaZLvjBE/Zbe5IHL3
s3LWS9i3MVx96FY73DQaumeCGgWyr0wcJiIkYERqbmfgedNr4LTc9MU7LyJdvjUP
9+gOT+mAHotUEo2d/fQ5iCfXIjiuPGH2sEV34EjT7JsBYDd9nIkasRzBy8OaFwxY
TpPfP6+gxDDMW15XzDEbJWloYGo63aHaTwywSnxHDK+72gMfwU79kFvyFfgjOBCB
GUTSChfPkUHzKziE7zN/LBX/KLaiCQs6JDWfUfs1GaR1Gl8rcXUImvwU+8+L7qw3
WQWgQOt1FJgjI94q4BIqhzhwrO3MVYltU7BNGoh88Twa0PQyAkG1gAdC/E74/4gV
Sv1d9/Dy0oq8CO9k2RO+xXGs4IgjFPOhknVpZNSuOsNpniSpbDmOImGCCBi4bnKq
Ujr1w0Ow5svyGPERP6/ArwXqZgGjI52DZKybMlVdviQMerpbPM+ksR53jEmU5WlN
a8aqS9xSgtTLWPEu5OfvtZyro+7dlB5JguPAo1XOND+sXeaU8kMstVJHJxggYr2T
bfuMfgA9bacWwO1QNBaiBf0bw5mCYfKfXVzxshE7JE33LFGp1EVmxgk3eZVNVf0J
+Logy0wRsaHGUtNyCjeztabBaxJd3gq9OqdWDuWXUwsgtEGOTD843/EVaSRCKID4
CPTjn1aoe81N7cJao55iMTsQ6P/u0ZKleAFFitzRkp511J0zV1z1YjkLzw+9fnGx
ZWMALSDpTMRBlXkRbofAdjqgEMJYBPzAk9vFrdQkuaQZovKH+yll8bY2ZVe50VLr
PC57NAxMq7WQNfb+ZmAAGVGXrIDK1FV188tU90ND8EsLTHzOhdXZAelamZlRjewP
UZJd7zk9iBCniBycwMuOcv9kPzfELgWZ3pvgVnF6NxlhY2DbXxeFI+n3FKcdvQ5R
7ejMSoB4Nd08SHvBX4M76GaBR8pbSVu3OcDxleZad8Aw+dHeZK2eEcGlQkAgbk94
JDLaAQlRsFU4DMJ0E8sAMZyPcgMk4f9iA2JqXDqWdJ/yEmFd0/6tFQw09mBRtuHL
S5TJezE4mBXDDZ83/aMsMeGovKyZ7CSASGTqkgKTwouT6VScHoifUJiPQcMsFHAa
TliyUUnzuf3MFlFn8Kut4BUzFhg/MSdO/Hklt/e8OBcKtZg+oO2tneAPJKg8VnDt
g+MnFz9eFi2YFqp+DRFKbIqYA/QFbasdxHc2cm7AbvKQHlbbLOfKeGCqtV+hguS3
oSe2t9jf1xaGMoB7cjS2tB0XLsvwVopdpme95CyVwA3BOtwKmcFTg4nwagBnJQIy
mbEm3xeMhPjNUHv6kXKBEYN3lqRoCnDZp//yEYZvgJNFHRFU+qfcT+MOzgSDkigR
hZmAfJ//CSQvctcQWldcT6s260M/zzDdYJIPXzt3CDDlyTNzMpBFhR/n3Jug5HPD
zCJXCyvksyYSFt9M8NoI4xehMPgJQDoWXRt5wlIq8KQLcp72dfMRygefzHclSWOq
TGJY52i30TH6jcftA7VCte5NtR7t73jbmjUy9b5h75+KTlPWPb7znCgvTReHK1oX
StqfTZFsqV6SeLnRROpqXEGxijlNM+ImyMs6Qvw7T/NTZ1AW1mN4VztWfecHRGJi
Np4/xpTCteZntBRCFdWCS8JoYdUQLBYWSbdzKz0JEgm7ys/j4ZXQZ1u6RC7jglEs
xPMRbGaSfTrUtKsbRTaFYaPQNzdufyOrCk2OPiZseqPz1PESTewpC41m3qYXeZwL
NMY5btsYN3XNoGquCntsIGLg0Wu1YVTuNY42AMH6B2IwcY/TCC4u9OGkJrdN89U4
wiA1Gg5czLVvSw1dxaDv1KrI6hd8liGtI5ZOgeL+KV2EGVscmaYr7XzaqQhO5QjC
PQulWNiiz80oiPSVjnwZzzI8OC9tvlj+IiyzGM9486SgD3EnPAGQVeEcwleDWvF7
mOM286HdRCiPoFENtnAwUzyO+fySMC93CeL8HQ3kKqpDCsoF3bI6ME9NH9u1GhHi
3iboPVOAj7viRCl8nonfI1D3hfT5yoeF00uGShCNzvocnZwspXfkG4nOxykmDrtW
CeILlBujh3YY1gmkVmDCPAm+L+MnA8aCtCLwZySdbLQBxVx9JcpiqqXBC4zXkOJm
fdZwgxuoBLnez0TPhvWGlIJnmhb7JzWBuveSds5/pFp/W5WP9VFtKBaoVimo5jrS
s1XESGKG2zhF/67D8ONE7p9Z3dNk5kkbgBMr5YXT/HZTlh6up0d3cAongiHP0xFM
o3faClbRnykfzULk9ZLUWYdv1d0XMDnc2WHTp5AEpn7zMxBunQJypjxTQsfqGX46
LJrQVhAdyT2UYXbqA3qv1hjOwZcj2Piogn4b1+uXT23wn8IRdMGh/ZCplXXwomBl
5jEZf8Gf/WfGToBys6P1ou+2IB9xccX9fjGtvfkZ1UHPIjRzsICSDn1qZIB2Rb9f
2XUG2TvJdxfuqIrZe/6MjUsvcyzZMB6nZyE6ZRkm1vXkY9UdkrvOd0aW6JM3CBKV
RiFhxaqouvxf/LiL+XnnWOOOAUjy5q/YI4ZES69tJeADOkO0S/BRN9HYFUlu41V/
OEu2r+NvsII1H1H+SVlh0poqKghpgpS0gtUI1C3YNDDNh0qCj4dcXmYSA3FPbzzb
yRImTZ0DbvkHAQA0EIPd4otUybrRPMtqIk+K9JQHjEcPNLHE2GOasvXKx9S5gu5b
zMrCREQKY1yjEeDhDV4XQvcarSn7kj7mKdtfk2ubhVuUiVsFq2U0A+fsHIQ3Keft
b7MJMiTIje/reugYiBAOA57dc5TCXgK/8sVCXFPZkAAf07KuwzvxcFsEM8y3sZqy
3M/DQn6BEEPdTCPLbT9kNdCGI4GgGhT2cGKPZwbjMf5mZjNFJrAMus6S9K3Hu0jW
0Vt5PNiAfh5BpFco82rjSLMMS3y63imfl4mkxnfgcHy7CPXXMeRNqrzykOpvFJEI
awq2iQ+klCzX3H2h4hxvGKqJxqzzuIyKaAEGofXbengd9g7sQ8Jdztb+cLTc56VI
i+eJbIeroft4fYyebfkNPQl/A+1zmB32CphyqL7VXn4zvFezF+qf0t+eI1epKF/g
jOhOIaC+fiCGAcS+1YaOcOqKb9O7n0UGGex/XbzTGhAxOtobcyVmqTEMjz/PHyHo
oLyQu/A3OHHudKriKHW/AfpskQ5ym/oo7fMjNe2OhAw8xHXuidqgK6mjiVFLN0Ru
zPWi5tyEVpFOXhqV1/Fc651e0sv6hDL+qB6WaAWfVjayK2Kw0q1RMcXgsBFaz4nl
OHjcsijZhJqRCBU4e5CWS6OuVCbOO2D7JYCgfRMwlwQ9mMmTZ6Ubs/p8ZFNlEN3d
G54vf3Z/9IsSQrm7YwSy3m+jsYOYaiSLschAU7lcU67+gxwtqkGtInIbULT8pyeQ
bUD6Xffl/uR93INfYPezd2bBEAsqAKY8x/M0tVP+Jldgivh8QQK7y0a/tZzym/ev
sO9biOLVCLmN2/DEeYwg9103j7EY76UNHRWrxAhJfRaNQnTa8L1BNCINczQ6bJOg
2H9L2RQyB2hhV8e5929ZvlLE7ur0dTzyrldfeaJJQpRgq1l5Q3by5Km0tvKlm7JN
9JInhg25kWauiricBo/zVQHPzuWdXYXDr/u2dDiu2VY2+Yc+RpZqp4uZTazG2f2d
kv4tjPxXcTpd8n7jDUDdgOzSH4jbFxxrS38fvvsDojJ6o9+FXv0BPfSCK8OrO/lf
7jK1/NoSl0J6j6fcWBkuF6dNl8TeXVfMvZ0fRVmCV+k02Wco5YAqZYPqAOTctz0w
xCCc420a3f5NgN95jEV+6w4dnSPvHIRO/znnl4FKW0q90fyvgUjawrsPfVu7ooOi
VIrtOPdA+rYCEJmz77BnBS9JYu3G2E7BBNQFfzCRqm1MZ6WlvPKYKCgE9AFyNqFs
v36rSy7JEx3UCd27DobzPUYmBW+VjDTNcyIiLhjBj4+Smnaw5SABbz0PjvBA9J2u
SEZJsJUrjf+N2Ag165uXIZGnaqoVXc+fIiarfwFqvjBTkx3s0QJtwLLWrwv5dSsA
8sFtoWuTNUZP8OS/sX5h4F2zh5bdD8LrKbNnJNmRYel1/CSMWVwaWytQV2IvyzPp
h8qBF6lCSKBFc616LXc2xGTkjhRiFHPhdElbw8RMGIJ/FufMIrVzri8QaFsoHVSd
vW3acnpJmEE1KiPfcVfluXnqT9/aRRP7AuQop07t86UZAlyCc+53mn1c4XnJ4WSk
XSgEJaja2k9uuwDdkIUdUfXfR5y0kEmxLtQOehvj96LWpxsEFR6vcTdI5Ynke+Nr
dchb6RYxMm56guXyx+z/XnDKGdQ57Kli5IhY8FFDULsT/9SG73GlYsYmtE4XV//t
+Af7A09vKEEIiK0UTm2e3m1nKn/kzz14Z2LPh+16PDyFcO07fBo5OZ5/GXO0d9As
ETeZbGptxr0qiWp6GLAS3TeCiGSivTB5KrPRSeU/hdHxjA8frKdlCUKMA0yq4oS6
WDSyLxlFsOqc7IbysmDLlJerIIrIv2Y3v/Wn3flT9m/GsFXB6Eypy1XUefU41RyI
Wz/aI4fS/oharsaC9Fm1uOA/7ACzJLa7FWZc7fu2iQNWN+JwfmwxxnEgxTF0MbmF
5yU8a6EW64eJAsArkSzSUThOLECgZnMH+dItt02kXwoNNwIIwOB4w8u2WNZJOVsG
oyAn1nI2EyrzAL192noi6QuQucs7ntVPbmR8R28xC+L69mmUzet7OtZUY9FpMLEy
4al7TqYzW/AO+X52r+bDYl0OSEoAwEAY8hxiKf1/QFeqt/4zrVda0AbyqsKpFavJ
dIw4BcBqLq1qlN9jC2E+aDKQvEFqHHVMHyr31BE+Bfswiv7srPHAGXqXE3uqgY0r
qdpFDV90dtUmYUsVeqTROfY3wN+ua+xL1S4fsobOBBtNHHk412/4Rf4j9J6sShI8
X5PbZtCftAD5QOrnms9HUet6qBx0YHvpcxB3JdLXC+FBSBMzf5GhmS69ioR5/Tjz
nuKATdJlLhxeBLEqhyYt6SXZ+hCDp+9NEvcaUPurA1cnhxX1nh+1eJafncujb5kY
eorypRPFZiSAv6vie4ajMr2WlKq8h7yeQ4vYvFEKwaSXge7sUarihC1EhSlTqRvY
GfKn+29KmHoHZlu+cgTjqr2y4GL13cTTzJtv3VKb+bf7Zt8Dll7W0uuekiXyDVYq
MqImZA7N2HPpCe++HFa68xEGtXtx305eU+cPe0M3JnPoP72Rl/DbfmcW+JaeWBbr
+Tc73LAn2WLS20a1id0vxYmaxOv4dz/mdoac9wyiTSEo1e5/6vCM5txzsH8mw4dy
GhOT+oHZivwgnKAVGOu4FtH5ex8v/EZstJ/F9rfeXfbojxo/MDChgUL/QLJIAV6l
C2tn3g/s5flGJhKNkJX2FUfW/b7r6Y+4n1JOmtOJIYtYxu7tatOluDNN9Xahlc5q
SJyvXxT+M7pvAxOOX5lkIhZYuVYitD1wPbAniqLaNs9fbPMBIszdfeU6aA+qYG61
wA9SNS1vKgh3G8b3JmiiV7BV32NdN5wvHGb6y+69rf/vn0dHf+B32PNgOBbKlyXl
wH4KxfjvTFAheIpZCajQYA64Lyc8ejCNNJILXrZO+Za/JKk2V9+kJ48RmPsFVb32
M7isb7vu0AupEAXYE5109e5qaO4BSxREiVpfLVnw0fEMIj4gYHTtwhrlqWNbOkzL
eimWRR8YFdYbEWCGDKS+BK4b4r847EqLOlLLsTFVIBwL6iwoZq3FrJ7ioRe27iEB
YccciWsQD26kR4Wu+W4zVOmwkcjK4xAnk3MokQEriXUVN4Pm/y2g2XoUQMprnJx9
P8nV247WNu5f4GTLmz3yAaNCWPUH/pIUrZjpLQv+SLb2NJa2cfq2KkAUGzJr2j8O
//kvgJyGDTlSWGWOT7iuugX2s7dUILonfB6WN7MQViboJBecT8Y0vPHG0P7S/Kod
XRgeEud3WSF/iFCv8S9aEikI9Br44KU+LrYvTz+5r6z5jLJNY7/7SW2sHvBtck3K
HVsuiapzqbAPMmbQ/I6MwHKsC4jHNV5sI48UHpOrE11ow7wiWdWoOs/dDedIz/h6
bPOuBAXwJmW3QC1vK84nAklEJYSD3EPhEkzbeFVsUfXJ3jUGUfgnQdQo0a/Zrk+o
Cl2/pLbZAO/P4fbCzpMHhvbFdJfJj81ySK9BmpoCNYVUd8exjFLxrhFxqHL5tJEX
K7QHYDhntLlU+hm+ONbTfRF22vld8asekruB3DOdYXoO38iRGkXrej9JRZ109pfM
DMuZrEhDPi9+6XIv/wAel19x4ZP0r/mG9aJrVIgx/7cr/RY3pGGdxT9YBB8JBRX2
cOoPpX3q1j5sdz8E5X8mrNti/VfKQ91WznfsxuMbCekYkY2SUX+gFvQGu2wo5pDQ
WaqzpXfKFZHQ81QDYpV1rvM6t681QzNuIgAsfjqMedo0AR5a6gx8A5HIqLOdqdZc
kHyCJmxItj4FVETB78G3EP8GUy7Mk1u55Y/7IQk8mFK8bDATp37IqirbyIDd08fa
PV6LM15tOHy0dwR1OOlp/5WUNed0cUOqK9xazs5Azp4/JhESQQ+Qa77P4ey9Pa4f
32kIKogQC1OMI25/HL4FT99Geo4KmTalesYmZH2rO/VsTjM7qZ3+QsqXJv8JrgWy
TKsRi9aFLumjyoSTrOlYvmPNpgV5X4dSIpX/SqEtVuRjWWhwIZOZPdK7AIJFeDtT
x/yXzuDH3HzM+DVWQ/su0S2QLt5ic3tL/3p2gB75QQh2ghxO3+QZvuyRTRj+YoHk
mmajhc+FWNfvSCwcPJ7/XiueoDMQsNg/7y5yipAulfijjLfSaLPJPTv4aIiz8ujh
i5umoTpcFBBTe3aysFpSL+7AcZC4NXmuIkCsJgaB/ThBoSRXdhVjialcHIL5CKTq
Tf4F7VVTQ9XMGviBPl21+a59CXiFeg1JWsLTl+4bacAMtmXkyEbqz9cwFbflz5sx
63HB2nrOYOHR/4t1VPGILzmu9NGIjkKHzHiiIpKCBmrcSi7wflD9uqeJt9iKIapV
MUIeFSQgPPy6m0ebJYozvfSpfMAtQV5wIyURxUJX0aPLEVn2B1a3H2RZ1KKX/zYU
D70rQZ2U5etCBNawSQNxg9XOmLh84B0I/x7Afaz7Gc7MfCkNZHA4rNjjkpC/DFNW
BLEEwU703IvLvffFeJFLWjB6vfNrbrdhQiQJ4GqboSbfgwduuXY79bXxELXqhl6d
rQ2hNyoSVN2cb0orDrN3fpxj/Xu9nYRpO3QfiOqeMkJJmgCoimvcH2AU6syzJoPN
6GJwnq4T0rAFsjYQYA9BbniqlebXJhofJR7mXgQvPo+gZQ76T3bRKE6xFPKzYlwR
SZppXYMXQ8CfVEnp32Zp11tTc3X/15czCc3ebu4CWLQqqzP/8CMjd7tk52owr8Ol
opbsNlTgA7nKM/5bcO6BzPfBxnLDtVAF7EMOCUmPCJ04TlTAvLjzEToUUSIQjt7n
yLHN6dla/SUkVmz+XrDuGLU3n0Z7+nkBjdHehveMsbvDvwkFAJIT2raalFIGP9ei
HYXir67rqEtaBATblVsj1XOZ9LaIvLYcBkhm3Kx2jL4PkW0vaCAfT2FV1KyBpDrl
U5iTLOVcdRs4u46Eo3f5Zs1D88MsNfdGZiMlTaWsl6JZlQKOYOXE3XWFmLUuxw1q
5w5YuDxAYNLfVL6p4cnvPk+NwuxL37zW4+bQi5PQEFOMMDWWRNpktDBM8bPCp2tw
eTUEWyBUDauKqSDN5MFfQStQcJ77c3X0J6TG7DIze/qrqwr1LpyS2jMX0AxCDN2+
mt6yAmsCIlZ6RakQk6I0RUJfaNMOKjNgEcJejdOidnVIMWI1rzfTrvFQ/hSIOvZm
2RevpNJ/uJk5LdlJ38S3E7eOj9Q6VmkuAcRwRH1dqecMtcwi/TLUiq4XYbhTN/Lk
cHg4vgbUUMQuCR9XzKWLAzmxd5K/S0i4IAXP+sNOY6N8pytSV3G5RaL7gweXFkAj
gw1zFVEIvalVMzcMP6SnRNYTWdjYQT2vSM2SwNWEqLsde2RQ0xdO1FmRalZhaoqV
VZmmUtWBOetyb7vm+ATK0QkWHS49bxecAHUDts2FgSWZ4xXKwRwYWvMm/cUlsNWq
mgWaoypneqP+WojeipEHAV/HutZ5jJypvnZ5CiHHwZ5XHRakgZUNusnyStGpLzvq
t6wHEbHec9id9qYfL9UWwdMBpxym/zeH1my1JT8cY9OeF+Nf2XgcDdLaF4Vq1kyy
u5uuT6ubWNFT7fzLwprbvcg2k1kg2qys+UzN7br0CXXEB0BUH8A/69NXr6ZZYVJ9
fyrH83U40DTZb3PDAdzV+ht3IEKpDf4ps/HP/Q0nEy/Lze6qvnWsykiuygJJRo9F
uuLu5JJw0ZLWBbL/65oswyDPuFBgp3EcpddolYNiR6Y09OGkoZ6/sUGXJyvsETu1
j7sR5Hft4vnZ4QE/+HZzSxnl5wVkqRABg7a8dvlGkdv0Qf7J9LKU2zJH25J7733M
wBR7dk7jgZH2T4CB8rov3U2FjzpBYUKTTbnjrkxcOUrrcrKeo7csVN1lIDhv702z
5fF0lkVqhwuFaMD+5qjev/wxRcQcRQ8mO4ZbbVT2ADZHxZxVBekPMjyTRaKIPeUY
V0DH2pRM3Y03Hk5YA8V3wm/MyN1WJvQMxobsmPGJ56qGP3Mnkigjz7uPdJ3dkqqo
lcztA9yxsfs63JHqSvziZxHY3sZiWDgiyPGDFZtDFPEPyFk6Y4rHyrrgB7ZypGNt
y9tsSWIIpibedSt1DS3ELdUyNr0CI0J195EKGQqD7tOXII8J8PBJEDLyh42xR0f9
l57om6gZ/gsy0Gvl9IP8/D6Co9WYEdvUglVd96vrMGusPBgey/VKxgOfdJVPXwgr
dRINkdcFYHjSm336vnnwqG0H9cD8CeW/gdpSuMIT9QE9sPFOJtS1SMwDNwAT4B0T
81BgNwROw7IxY9eBMK3YfdAm0Gw8NpkMeuRfsLYzOoQdqlyO3n5gubZiyGPOLnC5
QHGPgMYbwUcF3S/geomxPQDyGXmyFxTsbiXt7tqNv5TgrfnFBigFaeOw3jtuZwrF
JuTrxe4hZxtZEM9aEz/SKe9uMhMYjQAOC96gcw80zcfH2DtCaS58rfGWye8W39y6
kaFLWUvMo3mTyWe50shq7gA7NQP/yOaIOpXTeCmTkZPQdHcRc3//EVSmb/bS1hQp
Z108f6QIQKPNQGZq4r153GsF1/V3PcNrn7FF2swi8IRp55tJXkDXrlSjPXE7Wp/6
u98aqjPCZOmmqBO1qBDIqN4pQYL6qCoDmTEglrtcc4fuNvoy9BH+VEgcX8FBFg66
UA05YfR0zMuLVxuO0CjPe4Whjrjn/pM23pKSd+bPyOq2ymHBNoyzX600VR06dA8d
EIc3m07nH8X33BJk40EmhB2aVN7aHEptdBzNntwXl8atpASV3gV+1y7dSVX3v8vx
u0fc0+/UW+c/oxvNCu/M1/57jdWH4lEpAMGs+NKfx0e2k/WtF+t3GFyt0DKwTrui
n2Pr9BWJ57Aa8q1jKVUdw4w7dzMgV8If6XmdnmInu0RgDnO+XzMF3gyxnODWXW7m
2gvFxrME9CjItGFaQEvGaCy9I3J2gjZLVUUTC8TY7Bfep4RYPcRdI1kzErXqbD97
oS1w9kznm2Bivg4FYvK8TD9JfbjFpC+t68V6yN3LdUBxdH2rYemDkY5QtRURzrhE
t1Z+gldt7xZEZTXy/7kTKB2U5q9+2SBYH0yponCYhqAuL4N/fEG9fXUhorsIilk+
unQo9mtLneHTLvoEl/EM71aEVyIWbiXc3z1Sszli+EWGndG11QFHfwEJ2JVZDY67
PLnkTIJduXKzFkiYhdmGExSWjcV9NGPoCB4B4USllnmMG0P2RWkFGTrOLPovF8sG
HcIhw7h/TcUBROXJUY/mBj4GLD01IO2KgaTZUN/0f5m3wRYR8tsqHdZ6JAuAKLDG
IDGBTA++rZDe5cJY4BqHi6u5RTZlmeY1R/jVfPYxb1fCUZLv96ee94+OoTNhP7gB
EdzK6L46gXPprDorUGG/KeNgQBurYgTEarO5OB3yZ6qpdyZ/gNgmu0GxgXz7/VAK
Gyx0PJ57FCgk8Tuqmod7ByOBzw1eOUr5XK/VvF9nCUq0MsTHvBrCf3T2w8gvEPch
Y92RYQweUGujU7Q2FdDcYowh4L0hdBOQaFXAJXcvggObTSls9Y2TSeNTNzHs37rE
0iUehZ7LwFzeprEdNOO9AbEIkJFLAQmgsxB01ykTCw43MsY7tbk3BbIJz6yRahXS
L7bbWyZElXoSJwghiMtw/NeYs+TEh1GWiZw66n9NoXrJWlI/xAxYjeaq6nj+Eltw
xQIKR95hcUtWnh6qKFgBhbOByce+Whhkx/qtnqLLntlsANX6gQQ1n/+FL2j0d4tv
rqhBrFRoMF1tqnGPiAhg5RQG3bmpKIc3FIiiK5Y6wgOyLiTOsdmWrlwV2Fs4/w4p
9gDom+h/xzpK/2ojQtP/wX49Tvi5DUu3mu7YCj9L6US0aYjGM624FuUys7QQo74L
1cGqbh+2ba/6fGM0Adx1qV1EUN6jMO5W0N1lOrsI9QCM8y3qjQtus1luHLL8ItW1
Zr24rz5S8S2ZFCuuUX5xFylsk+cYf5HSHIhj1hKQ0k1hgEuVMT3dV70fFi3i6R+B
H5xRqc/jKXrzvxf7lnqeqbXOHSepXObmmhmDF1cINYam0edi8IeOfMgklhbzJJnZ
jcJe/gbIxqQmz7xy3bOoKqQ8cah0S1RG/pZq2TZdrPipi7Elg+nL27bi/2Cxo3Vz
7DxKnzJ31bA07+FnsG5bymOazOrxY0B8uAv0lu1yYkSP3jF5vgqiiG6I9Zh+aToc
XGIff73otL7dyQ4lVd+l0HOR7m9IIT3EqvEFcZzVFROijTjlSO9UiduMgS3HerNI
ubCM+p9npNJMbDZB45E1Q452UA6Spb8V+p570pA+KTPj4DsE6mWKNgRizR89SOuZ
kVXKS+RiC2ACBVxbdKMARd+BGg+OelSknYGHuNXqblTqtcgQhvcJ/Vzx1BLTviWG
hyBnPdxf30Srl7owy4LEyBg8+dPR+lLi5XWD5C1PtrHEV62b/iD8uPZJgykcZFTu
MG5QpfYUb5dBdeH4jfgycmvarz5JwxlZvYk1LKOKt4rQLIbKSi4CzwBrLBKuMTrn
tOH3lPb/TyEXQC/nZqK5f/O/j+sBjoqHzwSE24JhYemgtQACqEfNN5+B0N5VdbMe
YSjrKnoZh32TFXXtv/g8hFmNW+Y1w1K/2up40SOcDnvAFzfgXPmVj6V2/9VRD/R+
5O/G2NswEJxCt75+fuhwksxPdhrLdR15aluZak9x1lAHllPRt9M7k6sA/1TiYtGL
QHFahgfU5iJxHRi91NTJze3dnbNysDU7ZozYCLVUBbNHP4WjdQi5i07gliRfKnnW
kFpo/0jp8iT6u/V89oChonX0mWyQOVexy8Q3h71Mnf0Dz81uBB88KZAfwNNoginD
Foi2EOc6w7pomGTr2XCeYjwvm8nCMVik2GfFBz8QCXNpIHxEN2aeiISek/wRgmhC
FgnwysHELIAJjlhvnH2oZCw82UQ06s5pbyzTl5zelItuZyrBD6R9rwt7f/edAR6r
+E4PU5dwG5PEf55QpnXV2n7vqE1ldyckq7qiwzhIkpYmLHpTWGCaEAvfSv/EzYzn
HNtaBx8rAw9l4Ieg3OHpMxKQNIgTtfhJP7byCb6d4RPAK9yIHqDyVYfCwIZJLi4E
10urIgGohyJ30sgZzAsj9U7wakgL8i7jy7hYVu5DruiO0RzelZt9NvZOHUEhr+vN
8GfqVl/4BMEk1c/BTL5rzIkbRfVUmUyJSk+iBKQbJy7z9iM80cR0BA6yQPKvtxcb
B2vZT8qd3h5A0ATdBjnwYDg6xwVfWJaV3rBoBtxrGd2PENTskv6o4mUt7I0WMv8U
KTGP2nhseMtDFZMTsvJiaBy4f3XlJ6P9ZVS8FS/MQ9LkbkdZszro1mS4YbmcPeDL
0MQEH+JvFlBXxTMjthFLE/fwivy69ifVDFAvJOOKIDZi+RrV8J45RrvfdErsN2yt
ns6V+rawVLBlAuAGwnx25YSMkfSUdOzIxGJ/h6LKwVmnnF/U/xYW1Swp4Veftvjb
j89AR+To7zDSIOHxEqbtYBEl0W64aSEynfZtrofGkz17cwewTEP9dSzWwokKKCDz
eufOdkovUDXS28GMW0SijQl4BXLQPBqykB/B6szQrDU1BAA74ty+J1PTzWXFnTAM
hj1qINMN7Od2Ucf4G1AZ9qm/kdcKMk0nmaCxp6/8VR49isBaXoxL0VUAJZTG8Iy1
2/bDyofz4KLX+m+GtClfQRp8zeI3FKJwJErb4qCBVFX76MRom0o7waAUNVXcMXv/
uZXf1JSwHJI5wGhwVLjcV0/ihAZG9yMQs6LzDeVkf9TkhBNpigngS6JAN3Ez+fJT
HyInc32Rh0Qzi2w5U3tWsCIMbXwwf/xDgO3IA6Yd7i8TGDx9LwED/sZLxzozEB6w
t8b3OyZZK4D7tmom6cLp+yQT4oh+xl0JyFd9Fg6uLaLgKlvAJZqRcH2LX16iHuVc
OmOA0elZ3+qWc1jizwOjGlCGPf8Hv1s+vAUwtzQGD7Fg4hzMcBXVHM6lxxu1DY+h
p+AoKTPftvQeQvmPmHzgpWznksNfBFX5t3qhnf6oTJw8OurRs1+MwUq3Xzc0L+MH
ZBXndkGsdapxeqic2GzL1VvwVy725psxFHUH9yemD97nDKiGjAnuUZhQccsiDTtJ
Ex29zQW4eEtR1JThXk6uR/W0eVohpIhhgQTa5d1eqqX9SPMcF96rvM8xVuKOHunu
c0HXZtUquebxbHt9wc98EdJLiuyy4uPvhCHYRLEqmTcRPeCV3L8FogkMriGCAA0Q
NUGUcmzCmAEzWZnGQzA5o1go9vg6v5MXIhPZg6RFf/SBpPdRT107bw5HFpUTl86M
9FQ2D3DsPqLeiBe3GCQe9ieljgihL3uEkzCBYlUBX3KWYL7f4JnXqGpLhEott/W3
mGRASHvMhpPMkNQ9DBW+AMt0fF6EFshD7+5Q/cZRojIp9CWYFFTZbZE2kKjk/qVB
hWLJADsyfRM0byoNYN/cvEIiM8wDi8yIz+HnanNzX1vRSW5/DNxHDdZWMv8NkrB6
BQLa8lgIfcGIpu68jdagt093IBpnkCl1fBBPZ32kerNPXhc8Ll+e8OQouKXNuxKw
sF9nt5gTdQqDrP8EoI96fgsmpav4SFcz0cUDtDQ6m9yuJsdGErx/BepwfHYwR2cC
oWYjtBditFxf4cqQTH8SScZb7m9HjWUJsqwf/yz6FmZY5HI5qGDrcT539UD0wfMa
QPmq2+g3hdq2qqoi3vnErl5fbEuikBrHSEy91LaVT+0HGeF3pOvv9/18LO8b+rKo
jfbvjSeKHGpfk1ufGIR2IU0iy1S9vmclJeRkckymqzLZ2dyhkFMcoYqd1JUpe6x6
xqBBm4gTjLKdD3sdcjd8mG2RwuyWkrLsfyzmlABCm6RQ1XO4+yfnTWUo5MGdWrRH
GJMS8O3etdGFvIK6gt4IwWF+KGVqRkMCYqXtwl6thb8ZABIVMmrBYJpfCvJ1dVJi
tvZWLHd9Jnxsc4V3EtutljF/VCCriQpw2Sk/tYmVh0PCoC7hPwYyl2ATsXtIwXM4
C/fO4lm1Y87VTWLGXfJFa/geUgVGs15jTTN3jrmOVIFgu2yFDc/qQY/KOxvTNRFR
JuRyTAB1na0tt3PrPtDNveNcHQr0cI5WSmfF+Vc699XoCOCkxC9deqRROIikCCxs
XC7NKNKXJ45h9khCgfDM9aIaQWqh2gndUIdJBP6DEGFQbF6RoEfoXuMWtx/tI2yc
9lXJikD/AEHa1H+Ml47Aa/5r13XZRteXWka7ctIChQQr8cjjhrIEJh4gKxcLlvhr
45oXXAxGAzsyDvULbzWxZS3LlAhY0E1jBPC7BGOMdKR6M2A/AcAQ1eFbFEw1YOUJ
SvVWWMACk0IFMGyZfVi0tN9Fe2uvgeVkQFC57brKSEYZLmJQ1AVD2LXytcoQKP6A
wIAC4RG6bbyJz8nsb+J4oynfTtWnRSDZmakYky9LOrnveji9Z8Lg06gQHOu53BN7
809on76Lw4AK15QQzW8dV4ATmkipGUEFt6MplTwT0iyfQTrocq9MgNoQpLP/LSsb
/KJjnTCyzBUkdoMXlHVUIt19hv0YGFo0I1wYtB7Au0e6jeovXNR0W/SwZCrBYeWf
jRypKlzIuH9678Bmtma0QFzDGQnD45uIuXQVHL0FK+W7x4SVZbdSwGy10WLj6QK3
efRQyVplUrZJbRBtfRD8b+dY0JTcbHCj3za8eHkG5FDw1Sx6b8HjPvS4uSiip553
bnW66r0F53r6z2bjlB5u/KGl3PDXIFxyvkAyd1qzugkDWI4GQyanz8Ua2eSxO5M7
6SaEcHwghdVlfR0LpwRx0PPlnPQb8dfB28a2edO2tQGxiMXf6oCS526HzgA0tKdY
X50490z3qHMlkBK5qx5PACh3Q0CCnLcOBaOPLzH4+HzZ8XnG0h62GMhUdnc0ubYH
Tyn83kZMgzKF//JZPJd083w5u7F7Qa+eSi2KPt5UsI8BES5N8/oanu/IJqtaV1SA
h46hTw/YFug5Dgd9zTOGmfbY5BtiiVxm1ICAeBe9Nq4sMkH01yUmlfgEXQBDv42S
NZdeXvdLjs11tjex+KyoSkb0TIMzMiEGwU33uduRNrrY7kHvluLr9MbQgLlyQ1nW
7R7xH2e4XzzY9Fzd6wzo+4asfSQoeTyAnJcGXEEMi4rntXH7fuJ7vsoisdtvXfmQ
HQmMMBFJbnrDpUF102kPoS45/WxX3OMz7JtKHNkSwnn+AypIFdbu1BnbE/hbvUXu
UhRm1ZOGdgFUkBKJEFlOfa1S0e1VxnSnP+hhGpmDaTOeVeXWnFNG8c90LWoZXfVQ
lkORbGiaYnkuyJK9NQ6S9d+QJz1EygEUjFtxfaMN3sMnGWzWlZifGzwwJlcLVz4k
4W1iNyOgXxPK+5TgYFs1kAvMOGFVCFPVpiUIaeylOqsTbxOcGzCsZGyzkjf5RyvQ
Z21Ih+a6/6/LpkWuBm+/Y+vm3PJqGPUAoeyI5v3sZv8+joI1Nt2EOUeca4oQ0xM9
k2eEZTqwNN/TvVIt97tQVe0x2gso0tWRKpgFQzKfM68AUdPGORugNRf37HVPp3ie
UCQIINBtAwG2hnDRgau1R7W6WBdcPgOr2QVAZA5lx7+dV83HPVfzZxH5UgZWJfdX
QRucEJYBrSc3mWe+jI8PVYs11fhc8sfKOGJ6tK83TVz2X+Cksm58PflY8f92LAzR
KqkIJDiP2dqLiipVz4k7rLJKx15gn4ElH7gnxJKqzcs8+LfjmpHZw5CeVu8Pf4bW
f5hOTv2YDn580f3VmzF4n47oKtrIXfkQoiypHKvtA1HY4FaP9sRRH/Ru+xDr23b/
uVktUs3JNH1VpkPBsefhvBv9S/Sncjqn6tP6Xzse/+kQq8u+pP4H0P+xVnsrOnSo
D+m8Fq57kUV0A88GwSOlJHc4QIHHFJkbMCPV62UBWJYWB9x0hMU9N+xtK0/K++my
eGpXnNwz2O6sQOI1/AAdqMGWFChELk5cZXLayDpPRbiYqcv4o8h2p79AJJbwMWPE
cw699QEagFoyg1OWnb46sEhTaaYiBUk+AG4A5xbqLJ0YbVE/KVLYCeoH3c0gzvos
6vF1KcoLY1JxEdBnGJ9xnrYBFIYiuj/7fRWHNmO5A4xDQCdfRWei53UEjaYEg8gz
PyqRavytJ5jW+/Qq5rX7/uI7U+SKYZo0qkaTjDPTxnRwqHF0AA/2Hg/rv3fdrhY5
AZYdeNRPz5XrOkjWbOopWYCgeAhxrGN23jD/Av5EVPfTT1BHqtS91u6lIbUh8AWP
vNWx3IGt8jXalOtdMdQvlHP0T6WEQ/Yuju/PG/O1GqnH7Qkom9z3afrcH47gxShH
BMEGEfudFoKav8TYMVKUuhFIU8TQb4Si3u54H1dYX3BXWxYYoQiXiMzE/SSObXkI
27nEYaUjDsgJSMiYH94xq9pW3mKkAXkBK3rvS1axT6Z9GAX/rn0nm9bhZePjSdaC
dZqfdDncHg4MFw96YLjcCHa5uWCZZGCZ6cyPaVei0kXNdOOWapyLlpdqFZtp4MZv
J1GvkC12ysMTRoqxJ3hiqUVzXX697FZdJBtx48fVu7bwoCE9ZkmpBcCHPmABq4Yc
XIKXBiZdF6Xr5tvAjgutdtN2tTGGDSz1OKv0cM48dT4ActLCG+REadqRhfteur2E
LETYFdwEwZjTUgCDQN0s6RLkzMb6jAKdPQTNNhACqrkSJBYCz+lLEleAlpoZJBTM
QKh6S/XihCAmRD/GhMvIc5Du6BliFTRP8KiALzKdNk2eVAhHkmGW5bnW+jADNBP5
oWqAJwbe444O+h+bckYK0d1fTH1M5I6/HfK0h93EwGK1wfRnYPG0E0xPZc2ZUQ8r
Sqwwb7eiilb9jujncZSyrQfLokzvH2AKxzyI8/jaug50dIsw7gLgrMAx721E2rwY
Q/gxhnYlQ3+p/ZkKbEGThJ42AkkAQdpOueXaK5+peZXiZEXkl86PYJWkxBmXJ+2s
wdYy+aJ90aDGQWLvLa7P6iAztJviDUNL6HAfQLgFLFbjHnkFEAjv9hJxcRLAMKwM
aqA/Llhx9CG3IffJheHR7hQ8qu3DcYqu8n5eQswuTwCyMvQKc5ADbjN3xgEhleDF
oVT7RubzhlsD0Gp4yTNmlP4iVUc52pBT/d3O3DHQjYcb6M2U8o2cmyPYNuYdjxyM
xTvugjQZb6udC6fCNhd81BTOR77FT2VFWNb3b3OJ7ruRbqpXdJqBbTaXbkftKf0M
5B0FBiAbWMcIWFVFMuFaMlS+FzlCfLwnzywupzy0sqs6t67pqPdx7vMWeu0dtFQr
GrizSHlQ660oQZYxlcfkzC6Xj2CmFXFZtzMWSDJ/166QjjxcgopMj3fvM7q0lhFi
ppF+eE+bU0MOJ243RgKDlzXyVraP81vKmhtFowMbXLPgCqsDZxNdXXsymBi5FIQ/
io3t8UQN5oCFHFPcfp/s65xuTIg+hnzjHyONKM1EyYZfqJJ68pShw2e+2LmORbWP
CYr66o2Ag2SC1FCDdymF0CB6FAp77bByMP0yCbv8h4eKcY2nW+mCWZfG7sKwCvCe
hMXT5jc35DZajUNfa73BAEKpwUYmZ2ZXzUkBs7gf6cixuoNHlqolUkfJFFbnnBod
7bL7rtMCjNVWUyc65yTUlYkTOadpe3k2/qLiMkwdecYumrC2X0uwzKkt8dFfWZ13
KLOgLqOzP6qeKEcXMmWeXrr6ZnUOBkew0wfv0MrXd5S1PelV79SFhZ1I9C7xCGhZ
sH706+uTSJjbtdRAcJQTeZU02FkBPkafC9vzgSZVT6gGQHYkxB/hFt5GKb+XVd2r
gIydCfC8u8bWJZPFQA4LgrLLxbfdAq0BfpX+FiMYhrO63UEHQO91P3qk9UWuJp/x
++JUdfydQ/YAYzIrEhFQrWFR3qnfaoFHCxn+cMwpeRPKsFXTB89iVrubbEMiJpWU
nBbPEZ0M6p12C6krZB3l0XQhck7UamvEoxeKasfLhPoANzKLXkmhkKkeO9XNJhpz
r6Vbcw5e/ZYzKJeh76v3otkMEHldQv4VjvRti0dbX0SZXgquDuNx5SxBNxPrPDDV
2rlUrbspNiOId+WOC1THC8bL44vffSeg1szbfRLKYqx4xFxqndz2y4Dxg/XOteth
64EpQ0rzxRQZzxJaSs6E8HwkozaF80BYyUybr1MGSEqBifvhw2oC2y+JnRhJFMxZ
p84WLRzo/c4p6Iaqr4EbUFKiwoznqOlHDr5NdAEbC/NlwKwNzmu5+LYt6NHMWd4h
dksKMzJBOkrv5wvmdIdvZM8C1lzJImqwLlfCrOdvGjZaCoKsJzoZth76ZuSZZDiI
ncCxdW5mLMDxESfFlw7M00Hz/BOZUg6Eb6CgOIThGOL/t0FbFpk9CYbjcLV9Sxhb
pe6ffXgKSF/7LVh70huHjIpdzq2XgP1ynuXmq0HAUy+131ZzxC/ZSLysL3UBg+Es
N9ZD4ef1ebcMEiqtXo6fkAKowAXrDUJYIJZRsxr/xYH4njIx/pvrzZZlUMAJP+PW
xu4nyI/qMknG18LDK9RXs5PPKEBD6m/My4df0xJAGHwiFxMwPMD7siWBWpcl8o0V
OKK+8a2DQaHhSa6O8cN0Mtiq6hmZxPgX6zXN2Jttz9yPEDMCTIFDu9FZx3hJjzno
OmmWzCWR20vUvVX829NsQXt72xmH5Y6N9Y1K4yIzpGLFY+B/UHU9eA2yGdkeV5pu
Pbr7gyRm5M8puecJfUbSj2pikEwgD4+ZR1SpMwY0t2EVXjEDK2tZ+1gjBWS8qRAH
lFGH3FNamr6Ot+V0ddW6GTBBfpqRJeZxWXDItchwgR5chsyIEF9C3NixC/Lkx4Sj
jMXcqIxEVer/26rzFBn2pPMzOZ0957U+I7mLCN67sGqjJFmEsiIauAjyclDpFb0i
zoJy8Ec6QIXu70gjhwmET9aiv3dqGltI7Q/NEr7aokfBhA4kTle+J8E134WwRlE9
2xdEsVgP0wQOnzSD2z7YzdcCDjUVlE5ueaP6jZedASEk3HZ8Mb2Y/Z3xVMVUmkV0
jiJ5i5Dos7X2jk7odn8fIHygIbTcwr3Zt/YM9vXN94QThbK9rkN8WcCwrAya7BwV
Wum+sKG0bDeRVc+oNLgr2DN9vDLAYsYVIx4VZvCuZxyVuRnX9RfHRyHgETm8NSky
jjgBQddOeWmVp0nAEnTfh+BZXD9wleocMPcYp0zjr+o0JrBt6iYSomI8P+OAHYJ7
YWcZyRXCkvOu/BdhWX3if5HoFSkDPg83x8gIKIIQD8e/cVZ9gQu+6vC26essmXWd
QTrRc9wy010Wb+fJztib9e79HocdkQ5gw0xZKhtFSrC1u4O9YNA/BcgECwZBN9K3
TvxIF7i8Ll9SMHXvaa4pvvlbT4Yfs3dxoEy1CEWgPIZKxVsmDIJeJ399DcN6FT74
50kOVOc0VYKlf66WLQ7H0Ga846iT/fL/4Kb/TNcdQ3DXosDzb9SzdJ+ppCqFUyHe
Uz4CS4E3Yh66hhRC2wBjcGXlr8fnx06kRo3nuYGwHcfgBaxnMX/v4gdjAisf2gcm
MQLdxikfXO6GnFI7PLZc30hBOTRV0qGidiDLbDRWDnkfZvflSpxh9bdC7NQXCtJh
v9O53TZ0Vz91k5YJpfKHGMF7geInQ0Quurlrme0gLKBfZXhxd9/tHMaDb4VAAu5g
k6QSqL1RYAgU2TMrlzcxUjgbjuXwQndrycfyG2F0iiFPb3a/HXb37zxTMk4Xd8MO
tyfHDWeqpAHA9WtAFlEsWghf7F0JLO0/0ScJRm/ovUkMYMmEIKG3ZIdVZNnhlEd1
ha1x5XYAgZYuqCVYmm/qOdwNC+DZ7d2pMN+x3FC5ywHzyTVY17IJjRAVN1kxVTaQ
1NQWIijE1kw3fKL8p3fz0kxrGDbyvUIijEdDC8syRsAlfzpP8md/QULX2IKJY/ny
p10ogQZVi/ZTMOQFT8FxRuj1yAoijiwA4tSiI8soNbmtZdp8KJnZcw5S9HjYiqAO
9fKy4s6WTPIyoVENxyIacKOeiiDghwyng7nKqSa40f+uf+/t/yqYO5VitGUUrw1P
5zt+r/GfWB/tOIg18I2y/MLap13/3IvvoxYLevt5GLwbFAKTjQu2IpqRw1Uyt4LG
oN7ua3qEnELCsGwHNoDUOfVWqUIErSlbJBS8PwTP9TfMYpyg13+1H8AYqL+7LZgW
pW/RyzSsKdL0kreG6jY4S7Z2H8N5axeckFvo48DjqVH805K9smia9FT68yTh/rl3
FITyNVTPI8iRVdTkBCWs2ndtmBxh17i2Qvn/6OsbPIKcoY8DofUvwfBnXXo6KFgq
6vdIJNxv6CIV7z0BGRJ4ac3NQaOgGFcq1cKS/NnufoUmuddFGzLqoepNtxj2ufVR
G71XR5J7LgbijBKjjjaGc7aL7eDcYMDNEfPwNYNerueuPNvtopIe02Bii7lsWS1L
7kmtNUHsMbdDzhqNF7IssnFW8EQSSuTKCgakL58+0bWP+UsT84Tg+VQmjlNa7ZI5
8NOMmhjxs4xwmg9Tr1XRyJXDll+RZVGH+qzpr4fvkdA92AdA3MMQKLY8Gk7tcZkG
HUIXHOdeX7LOr/vfIcbMWSS4Rj8tavdMRoQ5XQ/vsbiboqwixma2W4zRu4JlVSCB
Y22X8bOwO2zPn474UzpGd7scXDci9mNTkYc8CUXvo+7D8WVVL28hGQNiSsZ+C5Ty
dn3aqZudKKb92g7uZfcfN/h6NEOFIKdl9+FDmnrierhNljn1xIan935AKGeSoi/C
m+3oOeJUqTDkpq1N8bmdnj+MlmmcANK9QoHawQQSlAWaZFOE7Kl5vzjbYS/hA30t
KY9/4BKzOlZwVF4fks0tNH/aSu2Z7ZNt94AHw1z6LAmCNH8JcOBCq7qk4vY32OZf
yQOFt+LK/do9ZXVFXZShs8v6JRlbPtf0h6vMXYvmF5E+mm6tEHT0APkdARN2p5/I
X2Urn9wqmpLFy7rnMPFgCCT52bJ/+z82FfJyizK8ojSvfgw/lvU0OKtIrwI92doC
djyuifwvpdvayMyr5NEsuGuWkvag9jbuQU9nM/KZfPUzH28if9p7e5Ulor8wyKpS
vSZPGMM2pWs5aSMNnyR0bHgPTFPDbTLtKXEG9kx8vVtc0wEQXQOVma9TTCpYadLn
CJzXwtRSdQDNSwlEwd1Czi3+pVYby2umt7BDQHj2t23l2bisUS8dxrEBHv+id9FQ
AeIjeXygiuAdZIuSDm2w2mdxK8GFnH28EKad6ZllyOAO83TP7DRHvQjYkgWeqKgd
jQNxOkQHwBRLypQHzEtyOSkhH0LuluaPyKiAxX+dk6VM0qfueHNOl0gjpqOzAKbj
IcUv4RQilyTQPlE6H7EwpE8bIPzAQx9pk0u22ywQ2/4CGGdWBqNP/EpR57UZ6ej0
mSnJnuHQI3mQttm1iHFYKRqx3C4sWlgoxfiBfu9W7+AOn85GcMw185IslS1ckZIp
f05+68Dwol9bZrLkG0Q+/XQiROmCIwv3XszoZKqF38xGQ88SYda1+BnBfcePDmqA
43gEnLJojNyVYAoaMV0Dt5ZFobuEzoSzgabZDsTtLJykI3VmydJLHvblGD5jk29c
7b95fLzuRrNqBMmjn/l7KFZRU7sUgpzFL77h+ZhC1Cpn01woj6c45lrE7TCJQLk0
PWw3ZURFZnrh3MhmPrKGlWScdA7yK7J9epmy6rGY3Gp0ZItWjuI/VTfO9V6WTTTB
skxcl0BlkNIq9W/U1+CQeHVD4I/f3cOywNVzvMmT/Ns6vEZ5v3KiblUDmT/rb6w0
T5HGoey3EawzeTzuXBrYgGOsFBlFhIXCMscVuGFrLRMlce+uyDEvRf68fRxJCHGu
oajY88vJgtLdEpgt03HHkkl9g6/sBvr2ymyYSWgMy6Lk31uX7CE746gXA1MUnKn9
x3fT9qGWl0FmHSJn2E8SZg7NATx+Zx4hr83507c5U4jkFfJuTvU4kdYflPvtpzUU
Tswvv8W+kLqi4v1UW6n2EYjeBg9sao4s6hJ+Kh+vQpgYdIEI/7pjoYbOmVL7lxms
SYohhl7icdfRWjMbplx4tbR+R1dLyrMWUEGUjimVdI4B8Czo/hCWeohq1AjSNrD9
OSsRWyZ5GkYMYf2M8ikX5vAnV+rl3OpuGOlTkortG03aq1yq1EH4ryGB80qj3cTL
pyNKH5+nAQ4VjrMe6BG+/nJrKSTm0ZOrC+7282hpYqoLmqSckGl5024hWHZxIGv3
rRIdeUCh5wFd+YXSRwiszc/V703PX9hN3Lg0U5vzD8z+Qtod0H/kuljeOyRNzhc0
wVjCLTLQ+t6O3sAqEeQNs/IuwASGCyiD8BS3dvkCLVIttVhP+8MKdYrIkeqdL6Rc
96Y68x0K9sAXGv8O5c2PXJ2yjm+x7alp+9Gm9zkycboPeIeY/oqTkDtstM/eLT8t
27Z2ZApDIbyu4kPPfpdzQjbjLB7Q2gI0U0yb65C2f0KPWyK+tkeuhf+hmLuiw+oH
LsIjQ7ji4iZ3VMmdjRpo57ba4ogNIrA1US8UQACj0DSbvAAVitTZScGnIEonliyF
KDxQ+yLOagirYpzy2NUQM3kbOwGiOqMeMeiGGIUUYgDwT2sWreMJwg+s+6yJfgaE
HwqEXMHKqAWnMtm+Jd6kzRMenPB38lwzUe3PJ2Yt5Utw9Zup1TKIB8Yc4t44VShS
TxKppJjBllVltfpNJ9fSkEd8DfaTqumdOnqh9dkityAbInYa+FkMaddTiLNhrxJU
kqszupeeC4GvEdohbTUL2PL4dk+GKmnWXrlKK1SfxHHc4Rojvvz7m0vIRaRr6EE8
kCqSGjWgzI+BrbzKhv9PLycPY7cYs/6hXciFLw7iVvQx3O7lqMSaQ40BHBXDNYcp
Tz/sm/GDXFfo28s2X4lfkgRqWUuKGSCQh7+a0gyRPxmYaqWSi5mMcm2RLlmMF8wu
rvoWvMJMHMQNFl++c0OO2ulTRK6t/cvWPLC3Sd92YbYgPV4yguBlZ+ONGExnXOXc
9E/WP3XUfaDONbXBEdgI3AlnXEMk969ovv3pjybWaJn0Ug8HtMV7RcFE2IMOCbIq
g1gOTL8oEpUw/XJyv2iu/5A0DDNsaTg8PCLXKcpLIjSySp/35NAlX16eorMLaRey
nVL8gLZ8MA5Bs8RsNCcaB9xZ3wcB7tVrTo/JCefIE4T/sOrxiOQmZDtwcB70jEP+
n3IRjUeJsRz6ToEYTIOroJHwt6IJNFn94ZAg1GSzaOOGpvDb7F2iy82qcLY5bBC/
CaWHsWRIaVvnFZOVD6NuS2V+z/LyTJRsz/pV+IKovR3EFIZ0gta7zfU0cynRS7tz
gZ/pvjnedtlkmLFb5aTqJlDoAwoGKKpdq6bhH36TexEIuQ7akQrZhAyYQGBrGDTd
UPqkNQTC5PCBxM/KCDsi8eeIG+kXxPkPtv5hbfevY5GffT5vEotsfgcoYP87I0Y4
0bHCxXWoctde8cXCLNBmNbppO+sWU33DCahOYErrjjHL6KnzlTvqU4yiId/+fppI
jutcM59cyJNoJUNW+wXDxb9KY5gnMzkkHuwnsEMrZ+ziLOPoYDw+wkI5Je0IszqK
94rsXOno74d4uHi8w0OYPvUXpM6iah2mOJbQ+aLJ2/aeHy9PY0oru/0jKNo6UAuA
YdviZVnEIerz/dj75gXRGK01LLyEuBQLihr+rK01Nnwms2E6pCupkuEUihOFMU2x
V513dXXddnIMnIEgt4bSmTaJWoQRYZLT54WNvBM/33yNYcJHDNRHZGa6YnnEucij
Pn0j989phATRm9flGP82P0FrqO+8qH3aL3dh2nIQJqLN2TJKdJk5o2ijMpoBvYu2
SfdA3QaMSpkZd1gAVPT/LrFsPrSkjsQPbrXU3S6yLE5If94fnk7EnD+fy8qRYdgG
Q9+tk88yVCv2gKQg2Bg5gTJlgO/QuXzx90Bm5VgONDwGbenx1pbMzXIcsWS7tweo
h+jpORltEzdbMptdWKDI+ZtzPMB+zZv5Ub7wEOgG1AE0b+FjHY6pKYeY0ZAUjwLo
ZbIaOurWtBxInGUEsWrhbLiaanTXG4VXhTcd3NIqFpYMsvAw3KvTDTDyUMra+GUM
MtysJguUW6nsidYflqdGx2Oz4+iYdYM1JJnWPVyrV6BwGtkiPhTGizKr7rROIdWj
ekUGOvpEq5olZ0OrYU3uacSYzqabRt+fFT/pIzHLEiELpmNIzSC31Uty8nSKn55h
w97NPrwkOp64WGwRb6v2tjoLHGBdZvliK+l7SKQ0NXsccwf80ZbaxpAns1FqFkK9
PVTfY+gE96x66uSPs1xTX8XpGZUHiDHseGziWAUiMezt421L/GWvlBKw0aKF06wp
vzhZ6I7MWjfwUpKccrRVLjKWbaujEoyBzBN0D2ZKf1s/C9btiOjD9HIP4hpL4sM7
E/2kjBOEumppfo0gy911nB5IORm+5WoHeiSR9VGijB88E4QtxUr21x/ihixucrh6
jMl29BODQ3QKiG/QA5RVAfBGbeu/JI9/o5R0cAaeQN8UF1uJOrCrcCoNUCouy3XR
AYr4DOTsPlRcTtJxRjx2WSwKf/0NpvKXKu+5LlPvZrOVejHCGirfrC7GKRHI8yOJ
4hpoAHVmMqhJ1arJtVHAU60EGPPcb5SW6bjjpNb4bzoy2xVltQ/G2QAWjq/IZwXN
4KWAzTFNrc+VP992Lz6LYqIHXvsOlVFQWAyIbuDXRX8KGbcLFOJHMYC2rFd4k/Xl
BABbBDlnQsqj4CUyY1L/zM3/FWFsSZJlO8zKdvpunu+NWa6WZEEBWotA/8uDyiru
v8nItwoL2pZXFlneFlk2vkeh8Oz/V+fiLXguI8YrBZefsP6vDGkfi4OoiBMuUWkJ
Q0ygliKCqu0WpWKy4djJRjJWiJErCaHch6kxJ2w5tA06U78yGhxKIZ6W0xH5/tDW
4YeuKIdt0dilSBs4xdKRBQlcNmVyb4lWCRm58UYbj9i8PCSXFlqvfNhs2eFjk2pk
z4buybx/OWirZXVtkbDrBlP+PaqvXYuGRZSoueSNcosQ9SSf4YYvIvb0s8AVyl/F
AxGQREkWasuYC/hn5ZDKRylWQD46aKrKgESMdGkHDgM+J2/os63HLiv27oE8Q+To
NeMPW6PXAhF8yAnuJvz9ArGpawRCZgauxI7pKLxaoYaIA/YSWkXu1bi86IFsuj7b
sKaWYdjhd78QRcl4CSEt9X+yrhp/Jw27b1XNSa/9U2eMo3ODk+UMtMUXpCHPF4fu
3zFT3PsY6v5wf+zE9l0XDRuKezz5uNXx8P6J3sYuBxjxU+tR4uV1xAGo0qPsMEQl
lMExSnGgTQwgSBF6I8ahvEa8cHEiMxt4AzSWRvUqkhuBJ8oCpTJ7Z6URzc9C0Lv3
1AfVSoR6psmzVm4jlnA06O9gLRxPnLnNtwnpQ4kHr1ct95sSCut5HbbvOttCj8JA
1UZgmONZaJESTWPWebs3xaA1SaAb05ANcnCUEJAbk6sNXc1c9yXt7Im4M+fy+d2+
XXCpM0lW47uQdjy9oFHY83puLuClmbrhcOKnTPYUHzcOwPrcKI78G/prh1EIRQtN
TSm1BjbmKJODy64OK6uKrzyQyJ3eqRIEKKcu+CK1+JUqKCRs2LrpCkeKkdaqvA/R
LelRNp2zRK0e+6GZdTMeyGslzYoElpgTxtv9TEjPcTdzxcpzEEb0sprNv76okZ0O
xf7hEQel6eCGB22PnPYclkmiG+08Q6kJsDO91JQTT5iJ9yyvMEI6zpdHvsB9cudY
vJ80R3gN+JCssUrO/UHi+sUeUD/R+JENO72eGm3AOqgUPXddCGVUSsxjYbtVZYCE
JDHnblyXto0n/wFTn6D+cw409BUlomCysQrc8xSgFHN51kwPwOALKoojgJVGI3yJ
Kl+v1jwhv3pkv6C0QOi9k0gsZwa//jYWv+deOPs11BLdmGMe+CfYVEQ1AeOjZU3p
CrqNeeHO0RBXm7HigjJaFMB8QCxFGmStl9+z7991tj02NN69ciCZ1hnhKwgr8Fns
OBrOjhx6+3Q3cZ3QttRKWGOJc1lbb63bBpB1jdfUcHs8z1FIjL/Gy/7XxS3s/XGM
fQsJvi0YbDVKv5BtfV2fqNZTPGul6dAu2SNqGP56NEbhS3AJWivzTiZ/QxcfU436
20knmiAqiip2xT5brDLFKMm3aG3lo/+4Q9b5MLKO0WCHEE6LGuWEX84v186XBquw
JYiPg2olsyA6nCfC1d0iUBrc575/HKs0v91FS45mac2IZdJx8Whhnz8u2HxUdM1j
UYlLuzVMwZNkJh02f8rRX6wrp63C3ZUFrPT2StFM1QtEkDlkLKSanCj9uOKn4fbt
wd+XkJt+LcLsjwCA6U3xLxf4YShfTjmcWtMxq/Xm4LjDQnkKEQ7URmar7ZxIBSAb
KVF6ftvI1hEbHqr4UVdUlJX5yJzMUXu8uR+2tyZzFqBfdM0TP7L2yJBZEUigX0IL
bJTVaXmtZrLYxIJx0Te+QBUHQH6H7jAVKdxafn6MwzWjrRbP/dN7WLN7Ls/smR2j
P10YN2D/y1QLlIoSW2yKH3Lk1dCH3haq0ksTBMWg7xRL12m8NOBt0hQfp6Y2xQC9
6+03fbr/+seOhYIJ5Jz5/zISDyM/V5SE29sTqEtzVjTTFV7WWIDs/Hs8h2w/25j2
uvfKJ6Rkfrt3N5vHmgvPQmWC+gJjnEv5Y82eNmQEQJvbjgAOn0oaGdx49bFSt5b7
eIdIYiQekMgmwo+jlhhZkGPssSHMgNEZxdd4WPFBTVQT405oWgcZZX4HM9CHnhy6
HcyeuyGouUBQqJaQaGBgEdWsm5MLsWPPjuQJkdOiDN0FFHkHBVFJqTVmUIH0xfrG
4iPxEtKwgP0dXzs7mcRZx5A9RZ+4jr0yAGcz2yBYg8OMeB8bZsW2SC0lBeT65wHv
OUibx0hoVWizzsFePLfPpwc+lZrmVk99wjQTDstzfem7fTgXX4t6r3CPw5X5/tC2
PpTWcCdw2wR598La6euN6uYRMMwUjRMWGuXLaA6YoRoCoDOGNDIMSbonH5+j5lAa
IJapNkHzl5U1mhPBrK1R3ls8hpNLsIz21G7lGCQ5RXQgmKWjxyBqxZGPHjWgxGHa
2fa4K+j494zTzCztLz8DNkYvAjHgEYajYIIBaxWk5pxXnfyzDNDOpJXd7uH6tP6k
AF2N2AUS4KpsVVEhWCk/VKxfNe5rSk+S/FbL6bXigRzkenc0O8w/+gWS5mTNtoqg
Xg5pnzJbonjVJSW/rvjpmDz3XcHA4hZn1y8DPIrDQfcWJDf6XHtCyPchn/RgsgpW
JvH09qUZq89wPd8mjA9u+ATth+2K8A3raXLj0wF4K2npDaKFPqHupsPNpWZ0LUau
uW1IyQo2ca7yNajD8NwjIfY6OoloWPBwWUQqwyR1RVACMCkhJSiDIjJgQCdmVdIf
tsbXeDoCZVJ7TJ8tCZSpdVvri4BPCt+Yi+UTc9zKo3ZtYmZ7LbxuYRLckDPFkKru
gUbH1zGRuK7Jv/XNPELJLnC26Jep/xzjBaOxgp9YqTNEerxvVP8rK6LUyLG2Wsdv
GK3A77gvfE2XlNov31Ketwn/MUrcvJwgk+XGR73APd8gFccZwoLJrT+We0t+MMeA
Z2X971gC8X3qsXVt3wT5vHdcZmHqZYr/RlpKhwn87wyds6JjgXLC7wHgBEb1AczQ
v2NDBkbZm2Su83a2ETYVWrddQ43w/1W3kz1v0ySOF/VM9mvnOOkUNgk7h0Wpk3b7
KKTAVb6+U4O9Xls8sDpxhkgc4v5pwELGPaPvUWhsI5hj928FH+pR9vy0nL2PYpsg
rKCmlcK22V2HDXFo/slSsqNAl+97gc76Ly7ndYx7qH+OXtJdHtEdzygTeHKFPaXe
05lOJq4hT86udGHV2P/hrdqq5pNWuYO1KlH61y/wH1e1DZ4aaGF36wrY8kLIW1Mw
TP5gcWhamVChefzP8trACb1fdMVpf0F/6jok1FhpyE+QFXJBUPzh+t97xCj9AQFK
BaVVZAAOMOVLP4xVZExbdLkzr2uJwmD7cHWFqIGvtr85ZyzFZ8c4ipMVTn76ZvSs
HVvxp2MdxhNfhuuV8tL1/4b/KxDHIyftTY7wWL8KMUcc9vMdJHq+fJuHeM5F163Q
YLXL5oNzkmJIrjzEOcfS4KleQm+WanUMVVte7Im00pJDSP1akLyK0XYU7Zdu+UOf
9eURYNEmNxIEKfrZ5nO1wTaNM40idKdXq/nvJbr5+6KBl0YRc4nvLU4Yxm9ZRRba
qswD5+uUO0Rvo2ioHJiTezGT/iOVSOrt1A3QsuOSvwtnmW1jwmTCqX5NvCCbi+RE
F2bPccpjedSkqLrlBlYgRzn5irQ48YWniwVMF2WrrgrcjgWF+4TeApPKyCR4MfCl
sUnPIA8eszj0c6Sabx8KTNRmDbI9O0P8YtBfsGMlrb2HFZCU3t/siQ/iTtAklKrs
lWzn3Tjrn6UoOx1Dkn0kmIGqiSerOvJJHLfwBD4L+ujHQZqWAGFEG1uRLkJTsOil
bZFGrSCGHQOpJUuDVBAgB7fq3alOmRbFbyVB59I/dADU5zF5K/vNN4hmLkSl3T9F
+fq35XoRZT8gy5h3OlwCe0eqpaBpF21ZJGTnqK/AeJmsQ1LdDEgsSJtngIjuaKuy
08+31hdt/IzISPr4DZkdBRP3x9ZBlfC35bxi7BlBpJ+YENgALswxRtYsSQwzOtsY
+gxfMJSa25ZI9FPl90rQI5A3AFF93M8KUEJuhFFa9u6N51yuyHZe8wKn8NXxRa5V
g64Tp+4vdnrAV7ADi4foIbg6jfA2h8jqlu3I1PVB8k0yMxm0iP5luhhYXfPTVxwv
hm7AUuDWEeBTylxUOwsvQ2bsjo/b19C4KLEpCV/LPxE5M61UcU6MCICgK573zBzc
ZkvLknsMOVAMrVw82Dq/yZeypRTUv3WGwFsvJCmIVxjgKovzxYSzy+YEExE0arcI
QvEd/zji4MVwYm26OTIEPLXfrTvyf7VPXC3BpsBlLsGuyP76z9/fafbyh5l71WCw
i1m9cAPF2yh5MZe98lUOh4Hm7rdr2XryggFmMMMQv3Fa/rXV42Daq7I4OqQKAXyu
wGTf3We32FWaA3zPd4L8Bv0L51oivLVKzUnq2eCxT0tIOj88aDqCcX10rW4VKXrR
cf2DxR8N1QC7fbdVFOlGWUsyGGaOh2eGv0byeGv2nujt+UGoUPeAxJVoswBu9x+0
/abrVInrC1A+2V9r6GkJd/37bmw1cVKrxstXFAmtwHvosadJomHR7pOPRCa6UmWf
Ke2KOhXVCGWVnYrON2U4xJa/mupZd2AVtWhKb8BZAvsDuUsX2wXgWUu0zxbpONd3
hRMtfJDAUWj1hzhaYfoE8tLRYtYKGcYl3PLEtUzxgZkwXi9kdd4U5x8CiHLJ2ckJ
WAL1FDkaFN0jDL/6Pq4Qpg20CnKFAtNfdtLaC6GkMAA+FNIX6vwMwR8yaraQMzNx
jiW7BmszyLu58jt+7Wn4H9WZR277SI+0gFVPKfDIuAFEz6a1wdc/APGmQ0FBfV2V
7H9Z6pzs4zDcPQdPZ3oQPgC7jswLtLT9lNnCIOhqWSbJnIgX6di+1rfhZavrdU3E
f4zGayTXb02VGsvfobK1ed6WvOx9+ucIv8Iuhchq6p8V3PCjMRkxIw80wKMEUpIZ
7AiDP57tj8hLEJKhu7a9qDj6NdT+Xtnrohh/Ccn5Bs0On9onuSREz3t26ys5OdYT
s3EMiMPlFhKtA3+1ReOZD4oXrvduJj/yfJWrjkGXxZ1ydTaudTFnq9EQCdeFITTs
APW8SA3xsLOxjYhojb/Htz+PLHTRozlxz97jYCVcCeZTSGj9OC1486KUU5pBcbFC
6j1uFRP+g6TR1edX18A6ZEjjhU7W2Aggkxum85SbKv/VtBBdt3KgTVWOslmIGO2j
hifuKeFpXAy9Q/zg3ifPz00kS8IVlr/fpWIPPETCCu9oG+VvrHVNReEK1KcFIkor
+8NRRXytzrluA3q4QTQF2WAJyqcaquD0k990k1U9evn6ya5vPYufwhdfAM4gSY71
tzESQd1gpm5Z7Jc1DOKQeUC4IFQ6IW9UYjjX9I+UsJoM07sJlSpzAoHGt15OcJZr
pbkuQ55zHYPxos8rfe4xR1tAXdG51SKBiqxowFChr/vDYzoOy4502ARPL+QjMUGi
E9m9L6XUkxHHYSe0g4F/VDgXrzgSSYvVHInfLuOVBZbNjxEGvuFubRfM6FSLrxhH
k9MSXrLU/PeszFy/kWLkrSzKdF3A09NiAkcVe0jv3QnaziOVl7WSCqyMYP9lXPvk
kN1xOWdvNl3HPb1prkK63oef60EMQxDSBaUmzva0cxbIYnC1WONaihkcw+QNTI5N
1xwFXVcf7dsW1PwThnGlZpQkzBAfxr3Tmc+O3dBQCkUh0dIxPwCOWj+44iRP9DmT
vl+pKhVn0w/CRcbigi++D7AlVMK2icvS1LpjkQoXQbuv4QSQj7p480AKJwKdigc9
8BJNpgKTT8ouG0yzJxgm79RutvEIM/XcIz/RSb+YKF+oZcpH3KVtGUr0XP1Me9hK
1GJlfafBlCU7s43WjkIt3ND5mVaCbKkdAYBgLaQtoj5s1qf88e84S/6eKuz/vbKv
NULqgiVpOQEPWo9jbtTbzZLq7l6w6ZH9On2n45TOSKithYtFQ1lvApYoRWf8Za0m
f/uEzejoKfCSwBDL2EPCBfLhjgb0/6vzzudOiWzK5y32ywyejqhrahxFCD8sX1YF
q6rSRhBiCaJjmkm/Z1bmk77jugphp//MM3yDjkNyaU9YuwC09Dayp51WTyoLtwV7
A66o3AxwKbvmbu3rGQ+/F+yBuYNEJl2tsg7K0Q4kDVZqhFniW6b8GhtIMkgWD6Hg
sO+7uOK9bYyc4jVcRwqYAaFsa4NG3WNigKB07eM0l0BsjlzQ3Wegumc9ZIsF/9cv
HEilg+vzuBWMpv+dNNtEI6Qrh8s/7AcyTyGAf5NdWMW4Q1hd6TaG/BSFX36w+cXg
dNdIBLwnnICBQsHSTJqajXDzMWJhBpz72UtAC81uaPU3aQDKa4zdtZrN48xYuJUV
LlGsBo0jbNp4nF8kJ/Qreq7AzqSueRPFMHcKYddJk2RBxJGf4NjtSfXvNBuRD9I7
R3AUczUyNqwvVCMn5YKYplwo+/FSZ9ANd768APjSZhr/foqhcL/hXcvxx7mjHdJA
T8hqgYcOFyAnEkdH6amWXaTbQJvCOEvkzUViL0Ew5deiv29Hp7U/bkjtO/OVIzCQ
t1Cmy8WIuCSHySy5MQe23HcAp4OveqXjcYqZCd4czO7hpKZ+wKvuR4TczfPMRd2s
/9Kw0w+LGykc2xu9AE3ypEFoo4P0DfkRszXsj2uvBTEE/MVBK48maUMavjvN801v
t6iD2RMadh2OBZDCtRxnGBFOXx2CZFLh+Br0L0l3HuePdaONmGs4MrK8OQj1lRWD
W5ZrAODR/rEcMIpO9L7qSCzWAYwD+c315g2+gUPEiVbE3yulyS+rsXnf4ve8r6k2
7mwCQ31+pmbXrjdK4hVZmCHdvQCMJPF7hMhAC3GE1lnK/zliGXVSQk4jj91fns1V
GicVNSHR1gTkpNo3r2fv2Zs3PFmfhE2JCFMxRRmbmRMaymKTMuvTCvRA/C+O9rcU
yd5iZUH79ra2S9HBy6hTDFT8tgfyFom5UpLApK8veb9jmEpAlq4cJkWKb/RfhK2R
ncAB8ZyLjSUITQZhiunVXjowvDwqu/zVgeX+6N6k+m45eAt7rix5zb+hLPQ9Id2g
OEz5vYRwOSjx/f21M4NEiRQTxNpgeg8Ve8gp4bcRhjS2MOfoYQpycP6y5kO+H1Qq
U1seaTPdKqDz1L56NFOHumY4AHNIOR7vTyCwcu+q/a0oK4poD55ES5soZQX1ATgH
zeqiTGJh6A8J9vPEbUF+0Ap5Ko4JCuewZsVEIVNtt53UlmtQI6fn9sYATsnd4rjA
3ITiaLe4Mdrdm1Pu/1llDjEtVgdJ/Gl02/Tg7bzJvj+dPsaGjyvTlMZhmLhPkn56
gvQr+LViQftS8BGtDSv77+Fin6K70GjvE6uSmGPSe+qIEPkaz/5XlPpAfzfL080H
42PvAyxJ7aLJGW79RJ2QP8EuaYP83a6g/ftBM5o3rWemMLvumxf7fBb2VuMdgkCm
wmfOfi9KAiNYXQ90Y/WkebDw85tO9vgleo0NlZg0+1a5xJWQ2/sjCyouuTV2iVKV
KeDlmZtahvspmWpvhmzQWyK2cGCS7L6UlLpl3fZpARYy/HcofBBaW8e2tjptPEdj
kMf1ZxaZqB7uTDXAaM3AWkCQXe2dXvR2bsZlYo4YCadq8Xc9QukUa8rt9o4z2j2I
TkTU9VRuxlh8mFZbigf1M4g7AAg97+uVSGcNwQbKadeCdl/d3Vw/tJu9VvoREKhO
VvplFFKXtquDOGfagXzxB2oq3Ylm0lzWjkpUdv+nY9Rehim0CskGP0mjhl81XmGD
kbkIDBdlAKhS2w75ekWjM/oucg8Za9zNyIO0XJ3gNUr3GWKKevLjKI7T+mFNeXoc
o+uy1QTJb/vnA1p+bUP19fD2THbaXUzrWY3RGaMDjtrTngShpQVG9Wo/Ci8BcvPZ
EpR94TQ6gI8W3xiDkmezFZ/ySYdJoig7wrYFYcgoEk95p7ysk1Rxhjy3sN6GuGxw
oNsJJcX+W4TX+Nr8fYcQotfp3vIUtbj1eRF1xz9XVlSkBEYR5hpkrsc2pE6mqLd2
tzbEXKAWUCPLBwAtGA601Ts4Ifa3x5u+8Le/Zfrbr7w4B9h6GeH0zPCYbXE/jLqL
8rY74Y9fGhRYWrwcSN6eHgwR2jDc7CEUMxUtI68HLONAtck214AGoElPYVUfUpEr
zZ1S9GF3+XWudftvCuepXmGI+KZSi06iO8OioQtQ47tYPSvkcaOX1k75YwrpMW4B
mooXxeXqGWgjKNuSomL4aRVM5GMl8XlF/KiIV8xeOH3k3vmdErxUQ7saIYWZs7d6
R7YkewYiLcTrFnDDp8VyZ66aSSE9BmQ4l5avmvpWMFqdVoFpmyA5ZjCKBJx/erp4
a6qW1fgQ1TGVntpgFA1Kmj5F3tJHA4+6Phw1LDsDKo6IY8fooiq6ySOEQZNr1UVV
HDtoW47i4n89E4JjJlevpiZZh+pLZ5EUgWiArqDGKXbt2+5yzviH543201h1osuY
sv9T70c1o2GFlVyzdxFTWMyOHjWiTmWFWgbZnSwyeSmXMs8ct580CMJ3YsjN6pgD
Gz1VJxYXEUpFVDXVmNO7mXtbBtzoDqYBQ/P41uj7vXuj0odvCIG5NJ2vH+WcI4qz
iPRuZtM8a3aX3wDwEC1PbLIFg5ylk+BeJ4INWCEHEM0iNwBIZomrylY42De6THMF
GHGGDx5pEbnS2Il6L3H0lmWadrDv3Zq/GRiwIYq/iVRwDLuuV4STTwcqzv6TXX7l
gjWrqkdmVZJ0VHWBL5N2nxeuJYLRc0qrx8i67meLZCDawAlL115qQ2PoOAC9cu/s
B3GNp/YCegqgPEVpJtRUMh5cBKnp2XrfcUSkYXc9NoSHY9V3LeDflqURkhZeBV2T
MLmFXiIYAoIyIADHNJenclsYD9OhCsPV/X8xKU5DlLPsRUJ1glTNcdMNxTfbZowY
f/IOj/nnp1YvsWcRbdoRm1VDEcYokW6YqlCZddf6dUitU1SJIxJqbEW6pMKv+bB5
5AvW1qhoM0KK2b8dgum/VFpto2TOQXwjHAn5erRylKJuFyq9f/D9X8BVhr0+ahEA
jqZYbK8WqmaQvwJFVDWJnMsKPzwQ9zzRIczh8Cwbtitc7KmbL6HA9B15/YSqU2Se
i+1VBzv3Xc/+Sd2tc0ryyrgKofzjnG317EGI4KGufkJLbanuIfqbOumGhfZUe4w9
WTO+JznjXQPv6macC+0U1LO4erov5Mzfqj6SJs/EYG1G2eJgnD3FXfIGJSWVx4K9
4od8LjpGuGXmiDh728vqLq6jYdqTFniJz1mpXvZ9wiEV5RYRGKAai6WhAiJOwkAf
kiuNRy+ie0YXj8xhy0I8ktGoCGGnQcGUK1zFqmgSziyALqxmE09GnWZMyYLhNeRH
DzPlQLqstcr3gpTui3A/LE7h93etXEubc3tMnb2v+Jx1YLKXMbSZ2bW8LGnSrgSH
rcDp7tcdbH2Cgc5NI2iJUg0axwy0Z5qhkCqatpLn0VRa/zmpPJN3/ZfpKM0BJzzv
rPyP6iQ5Y0MNZjmwOsf8/lATTp476IktZObcqhwDwHGLvhluIftBI9diZ+OciEKD
J2fbYuq14WRDFeRvQqABRdE8WkhZLEuxsa6b7BUfmCS0OrCS8rkMfpRlzFqDjZ2M
5c9jrXDRH85QrHtoNBii06SC1/hbSqI6+5RbRsOhYYDm3hr34iNR0bzRgJrM51yy
3HNlUNMIKqyQitUq/jtEzT7dNZtyqJwa7kohw87cI7sypDg311u5zIgBbNDGZ2jz
hokQMstWbYiBeCGdOFCJiaSb6+tocZwpdNzRR3C2LwYCd9cIEAMBuOAwwccV9SG8
JZ8BDL+PFpnral0I+Fn65OudVR1H3GTn0OZSDuF5UuIihTrfdcxHArtyJCvQGZip
+u80K9B3bAhne6ZCm45nA5P5Cv1e8pfM0KSOwO416mcmpYIQFKpfm3GHLO3EVNvr
HL8HDY1MXoBJEML6nenxAR0uxNIPnVCACPuZoY9kAgjLcyge86nozNBky0w+nK34
bvtAGPe388Sx3h440uq63UClX4mqswZC5seAT5mvR781t2DiFDxlO8xXD7ynfLOy
8aXaXRU/fhaqMgCF/HXVSzU4kBOtFKsUGkbkJUY3cSWsOGJBJ8kaHKstJ713Nf6q
Sg4yTm53Pp9YOOveZpvnNO269R0/hYvgpLR8ND9/BFNA27p6kyph6L8HNUQqBRgB
2Nu9t0wjgxY+G0xrAT5O36q+tTqHusgXZ2i7j2g3pFmR5AK+wRlQ1v7J6qkBgVbT
qrucd/TfnX/DllApwRbv7J7uqebj81rq+4/xz7p0yJJPZAGCNdw9+K+MVEWTRzQZ
z0X83BM/JBKspJxw5xFr1t6OsH9t6YxhMcbu4Jtxtg3BhRsSLgUG3Gy+yRTbXYDO
6GQ0FXLcRTEfVduAKc1+Cej6Iz1TOwZXWj9gpwdn5RCM/dzAGCKJy0iPKs31YK1i
hpAQrhyMDjt+1EUzU0GdR2zBKqWFIrZ3fEi3K8kCCC9dyN2z7yjJd+EQmEQWB5bI
ZJ5f90w0kPfwDzpE7TLXmDKmo0wqim/CUl9hD+6AOMi84zQ0b6t/B7jsR7SM+1kk
Q7Ib4ZEWUdFzYTPdO1VbIoxRRpU+fxBBL6JoKH3xPkp8n+RgI7PN6sPKEIemJ8mH
/S7weZSNjzkYuNULempb0y3C4C6t8RgyRLTtLgwGSk1TPv0O9lmLTDCgw2vG0oT3
eE29XHUpUX3XhCwMc3hfZwIxo+2xEfoyYsNSOftco+1KWeRw/29yDEC4NIqpLpr3
5IjVXEgw9QnGazZGYQxpA5u6Rn3WBcAQvAQeUYKBEzaQqP12Tzp+WQhv+U6gtzI+
wX4WFimov/sL/KZty8DcaXaFmU9G9f/xjZZe7NvXzRJvY9iUxVdBGK0WAXLGtmb8
GczwZ+zIQMxvGl0cwIaB/AaU8Ng9xGQFcW4nTPXffGWSRHafX4che8L/vpTbPXfS
MdqkEgTxzLw73LIrMS/lfnuwthI4uf7mrdcTM6qr4JPPTGJ82TaZLOEPaZVNxwvT
xKV9soL1KI3wsj69FbdjkIM9kTmuj279Z9ON7FMccmpoao6oTnJFHvJab8ejOY/q
oO1SsSS5D4Rb53bE5hPyW415VDTK+viY134r5fobqizp21e4UG3kMzL9BCYGh0BM
TlbvlOT6PHn2IoyC9c5sIGwv/JXXlT6BSjOoXd2Ns2JmdZHzFkQ45jy8d3Ld78Iq
VTUOrXsOiYMIkLA6OCh6f2frhF7uLrxeXGQ0fMbeh8YVIYcTGmt3mQH7NdjqsXk1
ceDSU7v6XKNcF3OdJP/qFethVl4S+wgeyMrj6e+UNZUWCHobxBiw7fwVF0r/vget
o5SrVIMtni/XNRDK11WmpqNqK9u1YOWujdqM3uIODOJsLo/X4LQl4efvbJFraR8q
CJoIKYbRrKXG4SdChBnGixXuhIcODLoQJEsQx1j2gDt0dGYftXpQqprGarIO8Y6Z
HRyaIHe9IyaXqs6UaGPYSwE3DPSEwECoPHhRBRhJwQV1QhC8VW+ycc4O9ZqgRPIk
783DA4HjdVNpWN1+dz6BMvQeUqUrp9m7T0NzvlUhA5w7fInH0o6SoHDxkG687DKJ
h+lUgGeFivIT7yoBPDLDL6NSxT1vb4YaVQRQ81gdEdabEQg44YvZfvXeL5MbFJ7q
qJ03aAD1sN49OgCl6ZsAj2u2F3tn8NXmVQxkZC/Fgp31RecfZFg6TWRJAv3QRG7I
Nkbv1Bt4QXljmTcwXJNZhGSDHQBMiokHMJtWtl5bt1J+CEGUIZNIUKDMHTCfCyft
zSq7zXn7qwvJsqffYbyFm7XOeU5d3N08d26v2OsQ9pZQqWcRwtArySqUrj4GhyI2
HlczHQpWOKm8qKhG3kf+2y/x5LW/qmhbLbKZ/U9oxOrR8EUqAq429978j03DV3yn
oXlqNCsUOdSosW3D1kBf8OJt0C5hwZINajOcjx31pBxW5A6X0zISO0CfXfqO2D0T
W4Og/TrPZphIE1ugHCaMkRsHifhp6fHVax6UEiS38LrkzPz2h2Z6iVkwHAnmgvr2
82pj37dzBRkwfVpgU4CqmFQYE6YSFAyg+FpDAjMDMOSAcoVHtldwz7gh0TZucsxa
b8UJ7SbrmnW4r3yVOW2Uzaur6TwArzM1GlTbPeqLBnbXRY9EtYbP+tg64b17yG/W
SYHc50HcmXkW1xsypOT7bsdJLrot9rC8FEh/AYxdP+1s5eCAkQ4ce7mf5Ktg7jkt
RIhVJgN5lg0qLrJ9zY2nFy445WOMttLp4qAXcqB6uveHrRq9b54Is+VjBDP6qSKY
OvHfpRR7YHaRaiosP5EIAGRCw4LC9br56dlRzZIa+a4WnURSb5jKchhPK+y3e735
aedKDM8yD3x2jPSpWTbWLaQhUm778ItQnBAav/A0Ger2zb2580KxcDiWtfh3Ctgv
U7/B6nzAJDK8SqY+kAbkqy6uuWLdFLNnTt+oHFaWkJSRBJ3egYlIU96acfhqTnOf
brfjXeeuCMOEFCJey18NxVRAU6gk5o8C6s6zFZCWsBg1St8DTLD8Jniveoap7bkR
`pragma protect end_protected
