// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
jwdjzffox4fXhI4jzt9hrk+oWfeKX300ozJ3iX0NE+1VUPzrneN56CbPyzSrj9gZW14Xz9c+AAu9
TVd0TNgdRzWIt0Pn0qdp0Q91UjIbxCG1KuLk3aXCYd7KOYiKb3u2Rbftl0Lg1FdVilfWnXOqCpUa
jlIB+FKyifpgX7nfKqP0mjim6MsEZ+IH5gFcspo3y3ThwxpZPSQW/lLWZERAjjR0i0I2jwll+vf8
UmKh5Tyb9sxPC0ee/oOPVR/xCrhD3egzFqdWHAqntRFulULRKTYq92uThPCp5AO5K9sDmQuHAEPa
tkV1vlV9Iiip2h5SnOlSOuEgMoJi+pu0ZKHKTw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
Ne84GpbKhdlZ3imRSFxOu2G9q1SO6okcCYQ02BvnaZont9/Nb22UzGZAiZWlPh74aCnnSmM1YFXb
SXUZXIdeyJTNcLr/8AghaIzyC1T3I1Pg5x2oIRS0fUblZk7PHe6vKYmwykFLMAjbNfUIGxWpO+PV
X4QnikUJ4YfHCOmP35Lq7PGFK4qxiSQUma32ut++1uLpVDST3gDlaE40wwauQBRt1JwJWmXyLKGz
BgaRCZhCufaoDlYJdRfcbOJbyRnRh8Vjo8KcvG3vn1zKwEjcWQDU1K8bMoBFPGNx+JXYj9GV7FXl
3pHFTXlp7sXJt96y7E/VQSwXkyv0DpjBPVUUuNekgxeKNOCNxj3dZ+c8aypAv4Ch1telo7GvKjI0
td2e5gTVF1seNsYVmm8XzCikTMQyEfR1kiGyKEJh4Fo5CMqmuFqH20kU9aJL2cP3Rgv8EVS26EBi
nIdzAZr5Lug7VHtVOmuR7Kjztuo7chTVGHfNwGar1OsVMvLXOcZ20kbCq7MkbTa27TGD00Fizaia
WQGFa4i5tqAC4D2hl3AaP1B83xvKZcuCF4hwQIYALZyi6LRFAnHCbxjT+eRUX64xpkVhORGx1iAj
vnMYUvDw+aNHtjOsbRphrle9V1x/WjpH4S4ZRJHUdsanBuK7+T3KsiNQ79qoQ/GMFZKkffBwYQQU
Fs9F8hIkIxbOo5CwKW/3qtL6WQIFqrw2zTGZ1rJ/CN4Jdok9A3pefHFsDASJL82hZHHlTqD4+DYz
gL5uIeCg03MUrPfdcNxdFd9IO6EpM5Dw28IWKDBtm4b+7oWtUl0rXVOef1y6CG4At9nXRYUkI+YJ
GULRcl0qO5zj4+Gr7ulWvD75kEdTgH8f+D9UIxhIhZdwZPc8s8yFhi5wskgs5zga+rgnj/2l18yN
HNn631Bq5l31yN2H/wgVp23wx+bleiyjXmSEXFEOYJbMSSe5A3QSU3+UV8KqSkP3qjKJmYgz2YxK
rMPZVIRqO3Lr2pbinQlBy0IT49qoPtwkFzBkv+F9KsRvyxgVRzGONXFWi+8WJh4eUBQQktXaicdW
Qjen/2rH2FzlA6tjxQw6m/3W8Xi9u5yLeqZ7PbJKVXVusqnfIP0om65rsbtY+Chhp9dr5rsKw0Ki
pqR/jJDIvfmnm4k139Hgon9cspxdIS+2AkJ/lj3XzqjW08/mrHoaCYn/U/A/zVJH+OLnVL7TW3zv
nBSzSQlzOBVww8Z8EfIJXimiOWLdyOkl6WG6MSN2d+ypVsFVhT8HgGLj7inPbWYxbEnFtx1e0+PJ
Np0tmlEzHP5fg+y7ae4BfobGGFjCGMRCt+Cc8HzngvIF61IUrLGiP4OPvNas7OjIHHD78F98f0XC
EBlGmILNWyjQuY3sm5uQ5QVCmx2DqMcxGpKUCZOVMN1SNMcOK93VZiGpiMJXmlPfqMiXNvOGzgUe
sS92QQ7bFwDKLpz6fi1ZJMPBG+1g83skAy5CFmMw6XFihkdiPdmgr0Jfm+vbstBvkP8e/evJCUkS
FtZRJ+qcBbxHkv//4PAI3QB5td71fWJWizqZOnwg535eDOhpbmFve862GIaW9/00zIpWrOOYhBOe
0mkxdp+tds85GeaJEd6nDAvWxz1gk7kWIhwyhc48Uc3AjH45C8KDL7ZcYxV6Z03eMaW3+d2B/T+v
Wjvt0HmG6ftlAekVYXyjBnfUypnM62XKhB1t734cVYor7LSb4nxf6BnkgUBOtIXw9EBCJM9oVeJZ
4uyvBcBYlsBDAAw8wOTK1GSaW5KlQ9Q6e7wAyG/v/8E/amO2XijUmbWRU6RvkIjGB25ZH5iMpc5J
FZJs0awNSJr5gUF3yXvMvyAtZbXyBtzNLj2e/SD9AkZ94dbCG7PPQgZ2T5zHwqKT4TMf3amki0Vs
Vfa/4yOmz3ddIcL27GX1XNdF9NWfZFWrg8pqAJCh8aChx58rIBaOeMpbunAA0HwRWb/iMhQenKdn
/Iht+pkCwwosSf8CRfj1r269dp1wnelvAj00LAhDgOQaGL33dDBpQBZWsUdrGr7eANRB4jIDWbN5
uaosFWVsd0s2drqzmkhGk261KsJG5F648TFs0DaGIWuBnT+YvE9ij81HlJT6XWbCNPS5SsB/FaEY
VXRLvFuN32ENP+8d+cchChaqOSvxRnuStfiN78Ei1GfTvOm3oUxWYHrypxgYCYmeT/uc+atQYnCT
IG4Q49bRLQZzvWWpviD66X3Gzd+YP9WaFeOk6QY0+7j/g5G6g0jP098flKJ328Y89hLXPbLWJ8gI
IksX2IYubCXBQGICN4i7L1ASRbaTiWFtQU6jL8FA2tWKzVeWvC0pqhn6l3WrO+G43aQVEVfAP6di
Dil3g74O+ts1T+2aM6cw/23ymCp9toHZqAo/L4VU04Wf0EyuCdT2E9+ODDD52/6wK39JiQ/9MANe
4+xiJdrvMHHnTItzd3aQ+8RLBEdhQoD2HbA+JwuAPu/KipYEiJDkTkZRshyKP/8UDLZn9IjDtWUT
0GAsm/1OJRW8QIoLSK+dIv2lGtYpxhUs/+tqcYvSbr6cdmYRSA2DNGeRKSa2/H1x3/CzyhUilcEf
P2wNYx6AYla0ylGrAlOYiE9bd/BjUOklSl6nHAJaAVCFmB52nZrTvwLF6YlD2AF8uB3AGt5y7nhW
+JrmAxuenrGnBoSYoJn0ZTvlEThmhnNWX5WZkE25JWGME3DCqGatWPFpgvb9CehhDYVDo4Cp+eWo
5+05wSQ7BvmaUFhCIr7O8ydzLCUiGeUoCs2ddIUvDfWdipJGneNQNcD1nEdnILncXuvpkO9ZFDzL
02oiIgN/0bfqOU+LU1mnEFj2mLdbv+Ae8eIrqWBW+HvUG/j2L15ueXJyy0pcINAlMWXWwDFCwmqo
9FB6TebvcT8fHuK9bGyn+CHpt7SeQ1ZbGDVm5BhoT8YzqwHfo8eNMVAe/yGm+AabPCaMnueVyIPu
LwNyNG+UIaaGhawTDhin3B5XIKjB0VcPJ3Mm0B1K7jnXeFPQmLg5hgt+7GK3pdqHEe5JpZ2543Dr
kdO7LbTjNLhdBZg1XGGVOMZrrtkpwuho0ncKRw5pcB4GeJrkgtu9w2PltvMxJ7wB+IiZ+ZYhhdtk
Y5xGya+pSmUI7EDMlHYjku4KHHUYdih7QxDCaY6Nqgb5Z1LeVeqfrD/iAAQtd8/tgn2KJ9adhSim
7Hw7oR4/mVfqtDvRxyDGUZ3HQZXkW0BNLFCSFBhm9o/cR4y4oeQ51jfUWix2/KFQUWFMVvzMf33o
A+Ek6xiLzyTfEhrz0V3Ph3S797MptmqPWQDWT+G2CYImL+X8CKLmk0IgHFQWTIbrxQnnaScKacoI
pev2EwAjlzDuFjSiPNjHA7oBktvAREiG9uYVgnzXOyBsJf1Y/sCW4iDGcK1CjZzifXIsMyQe0R3t
apDWBPOosKpOoPc5NrIw+dfTnQXWu/+w2ncL13FL2UPOT+eQMQunZIQicYplyjgDRKmEu+sAW69g
U1yj3EjE1OgHFjin7A/ZDZAq8DZpWP3sxqsxl54pEmsnC/kikKXVRJ4fBra8DvBRx5ZV64OnxST3
lYzqrngk3SUnYN4jfeoH6EtiNEEXK8ejfoQ2oMP2qvJCE2OKmd6MNwFIR8/QUDGTqhY6yryibIHg
M9vK9YET4lU8xCQZ03xGf0JgBrHA5vTTcQeBZmIu45TuIJnHngFOreBukFpzeKfO+mHpxKYsirzF
QIBiybV4V2YKYkdsdAXmd17dXp7wqRqbDp4SZbWckHW39RCGy0PctV7QGW7p3jibMkgYNNKqmj4U
k2geZkjXGUIyO0ABgWUXNVBMnkn3bESkLrdT5kRxdocwmBbNkeaL0kxGFvJwQUNTBNEc0TM4pVQL
Vb5ccwD1LjHx1EaTEIlMSM/NHFvglqEwvSBFWpV30CyEX9Xggm2b6XOqB57FnRT2n3UKt00ieRwk
rwX6OMUguTsQWCLqQDamOMqSDeBqDVyAN7kPnnBLiqsQlY2PXvW9VUROx8rj5wuieYScEXNFLz6t
q1P2G3KKKH3LpLB9KHa/klk+7+OUGW79SF/0HpLLPyMvN3Z11BXNnHwT940JRdKrBccN4hY9WfVl
SyPa7K5eA3Ll5FqDV6ss4BHMe6mkEBvNPL0f+QMon+vjcvnglDrPqJL6v+7t9zGzN7PmLjqBROOb
gmQDKCK7v5anzWxS9q+Vpiwgg9572TYkVWt0s3yyjsNeB56fca/FmJJjhcutw6vBAcQOoZ7ZqPy8
WxC1S+qUIDYKbENfo/JXgrTlF2+s0fcICODbzEyYhg2AtpdlZw+dPmgoa6bRj1RAuBX8j17SaPOz
jUlMya6W7N+PioBpZHHQUnHHxJ8zBYgnKjcXF1wcXABLdWgmeRyF3LAqzkfVXoMLy7UyY0pnA4Ku
k8fwjE5PQ9lHoLKQcXZCxj2fsx0GRSgPYhwTERshtwOncFYnJ6kJbeL8CEFMbIPLyxy7B0lD0zcj
AacgZspjFQ95X/HdtgQ1DpDlTtpXX734DUKWfUrU9KWslBSOkUkx35/eZGSXUpE4j8nxSkNgSaFl
A6DBaYvWVLKjP5znDLROM9LTabaKg3OLjRUkdwvQg3ItfR00WW9OkanT2w87oxswOUHRVcwmixMN
axDekP6j0IIPNzbPTpgky8MDXOmRXrpy7oTWeccNIY32Yy5GyfZhb0LSgYExjySpdG484W9uYwL2
QxI2u7BJyyGA38OliRzpjC0tHvO3aCBhJahRTB7RnCfg9yxnJzWnVQ42691XO2MXbVQQD4yNv5sr
hjlpTBjWF8usmYgMtrYuDZi4SwIdm1WcatJBCg7ooJ//LeAMdnhcP4Aeri6WNzY1L+UHTs6fQwVf
zfDxV6tKpL2GqgDEcZ90e55Hm5nvxHH2Bu8PqIG5isrt11g/cMLW3dbD7Giq/IiBGvPOyhee8LPH
Gf3xXxWrVr9WD6b9nyheVN6jaCXuKs8IQ19wOj5nZCKkHGz9onPC+JrgrAS74AFMVXNFgV9FZEEc
JdFfjVkKpw5zUgOlXMSf2zPIpQvMqMxCzUSUtzHsJE43pdCq753Ng2ebr/X9+rPXAOImQN39oUCZ
3SO8AMPPDHhpGMeJd3+qhT2GULVklnnE/vLdN6xGTYg5eJEKzgefsHfVrKnJCfSJ+zD0eJ/imFZy
xOXCsBmp/7mOccoABkJ6DmeTMNa0XvUuRtimNysOTb2+DAzQS8zpktnn9iPvqnd7oNcAeGz+BLVV
xGUkNqgD7gWl429n9gCHAgaocCu77nCtDx4vebdmAvGXeicz1jTUvGmKLjQiAkpzmhzJoXH9mOjo
D71ZJklri2TTCmaj7soct9lR9mVjGoL9QA8OOH7ra+AsUEKbPHDPwY/53iOj1h0A+CqjdjQsdPmX
BGXG2Wfsy5XNndLgfl8VJ4Gi2S9ThQxTYY0IQYAhveXm0w/CRLTyNtmUavsTx56zCSs/kWfsA7vU
6ADk7v92z7yBSnDGTfiGxSfcjGdo3lsIv+GWa2MJ7CAOTthtmS5zk0wtzWr8GH4aH8zacSTfXzju
++onyJSZz/NUqetXMgoo2sPaBfTB7zdIUBjCo+yhiz+YTn2EPo5DdGfrpLPF5foBzYOHRjMFsGWP
TnFGi8yckiYCdf9tXMHeBKawbyo1lh9JnISOUpP6/Nbc3YQa40ElnUaEhNr+MSOLugUUZsYPP0lS
9ubJq8aoWIKMy0QRY2jNNc+ddegKXbT0Bx9KWlYYgxvwiWHSoBUqyKpHEL0IqbO0LUxCc2tCexJJ
J2dwzRk+lO68KZbuHRcwhKzafQLTqaKtHb9cYB4pwWnBDjKolTxGrQlhrT+5jf1mALIWabd8oM1A
7WvIxTsbyJ3+upNgZWLieYOYL2fymifKYyGlGj3UMROZSvmRvjkSiGVUkY0QXn17V2JL6P57ef6F
e9nCx/xnZEWgeSPDgJgjAlRVMXaM0PoRcTrOp6pJyEHPIUQ5Ckp4jlfW+yaVaBC0ZaIDV9oGWUY1
9yjERnFjzzKFX9E8G+WKWhXhbVUrbx7JARkDRSP7NNn070QZg0bSwCMdmKcyVBHmsB68EaH39DV7
eD/Mv6aVMeciU0JExf832aF2H/w0EJTEz0kAmtYuz6l2GbpEqI9WrZYdcITeJbPanQUNT5Ot4kk4
a7nINrVzTmGy6ZykL0FDM0YP82pk7M2uAW2TdWSKRZtkkMn6tGwxt2HffYZYTNVeMZwXzqF0rwgO
7WeKJpeQGWiMTIyShfQyXE8zOjs0USp4OC+2nsqlYVCkpe7MbSuvxjr+nis+qXxtpainruLUUzfP
Y+XMRfvCHOiSedcpUU7fQuUpF/A4t+IUB9WK8Jaep03rVzNA9+3BzQ5hgGWY/ZG32fr+Pn96RU2V
qHW9aS/9+Lxf+5EejH2k2SNR5k3MlsXe/ZlstMucFOiSdY1CWWmVObhqcf+KxCEp2rFuhWu8JL6E
oXIV3Te8Jw+YleeAKlXw4K0Eg0uKS+009aEFvOeo54ZC3woEA9lWDkZP2BnDgEiiIDU2TRLlbmwH
1j7RWHHG2/DBeQbXUhe+vRRDZrAshNZvs4DV8+lIbN8nWQTxx+dh54Sjd/fGOwQ6I2wx+5ulVpzG
0+KtkWeHJxzUwRBesFe7hFR8vdseVwuoTAY/9xNj+gx31l1eV0UddzhCJ8wIPG8/0Hmlcw4PdWjd
OIw6sLlWzZO9lxpUlZBsW336h9hK7QPnM/Iat985VxnuHLDo9BVv/RbOJWAlx38ALxjAXatrHGdW
OXC65Wla9F2becf49CanpywwlT5eGD26lCpUV+m1f/ZeRL0fYj7qiNTsTUiTuMKmjzhGymA+tH/m
lqKnblV8eIzcPIEgQZtkEYNwOKlGd7IpsLCGRN5Oo3WPIGI7cCnd0vtSIgyflpZeORKOLerb+qkm
p3ZAzwqO9tQ3zZYR/ussLmBVDYKUDRMg8byVoPXUeMmDHlaGoH4SP976PpSLLlnlnQL9W879Vtur
4pPRopzoDllLUUA1t0PTjDAq0B25h2wssNUrCR1t79F7/yQLCR5r52Dfh+4bPSVrXqN5Od0JhKmg
XYHEZGOIiELWsku6NztUtTSN3yPQtFme3zNDZlQgJLXq+9BZ0BXAeJemVfsZQ6fy4DyWjBc03+Z9
PUBSmBb2qU/JTZ2tJ8qgPA0JLLokKRzZz12pzUO4bgouquQk+56Bj6G1BYI2J6Dj7onVEBV2KLJk
01x9Ypxf7EkhBsQ8K569vt+g2/Qib/aSLdFwCpnQV5RVFe3mgOjfyVEQrRQI6sSeLnlr0oH1L2cd
GOHE1trWGnPd54Y0Nbxmd4tlRGisJR12f6jT2KSprZAfuirCMlywK+Q6ihMLZWgvmpVzI1MJn50D
eNYVMmILqnEyz6SmOq4CBie+UzGXOWsvO2ozHtUkx3UkHuew9ifuaUTOYtqzbaw1+s6Gx4lHATGj
JjsY+sGX7YSirCD/9wet5+fx+FuxoRsud8PLAL/6SLLA3QvwxHrkyOtRMC2Hvhm4vjlBHuKnCO9/
cmQthZNakJXc1vBlIPdhIvdZo76wHjJrrsU/EIJ+IAZ97Fbrnr9E3MpQNUygRXPgpqQ8g9KWryqN
R/Wmggh5QLersCBhncdH8KQeKUATaGwDDXSlHAEJuZ5pYQEkvkalT/KdC/XffhESnxTd5dC+6RmM
o1Y5msD8ibRq+bjFbiS3NW/sqcb4I/daGpXMZUDoUCqdnqeRiwYRWbElWzqjoOielH6KFCGGBKyq
A+73ArWQkq57kyP03rPJSQspTemBuyrO3DBTecTnqN8EjAPPV1EqkUkBWwGqm0M97EgTOcqbyc6p
BTAST+ELnMBXAqVmovZ7Q8glcvR5KpkNDP+Tojql40rbZzO50iemZT3v6+6qZNmpmjGQ4MpU8VoC
W58G29r21MRhdX1EBGBfmbpdHijw1wB0tNmA7f6fh9egBBw85ZB79D4Zo7YlM6btadzxIpjMj1I9
rV2OW4l23yxohzzyENS+zLoOwWmb2Uq53l/+j1sCOV1AX5SEPmzN88CbPqYkYGBb1MfaOvzpjoE1
MznXmCXOL+NfUCaUNHzCQ58DUvpYy+Nc7TRIxnvrXrf3HhYxo/+53Yig1vrmNvXdmiz4hEF+zWGJ
QTjeNx80dsMkOPcom5Yt5vGUYi24Zv0hRsDmWb7Y+gWW21A7Igk/11KWxPHJ+zW0PpPxYw1BT8EX
l9AG5mTJaquXN6xyDP0wCx7UJPgC8atpWWAO3EFyDhw2SyO/JRYhgjJYgUlUy8MAYm2LZ1Rlea85
285nMqExzqcfqxYxQriodlygt1W+rDLQK6IgE2HBCgzh3VTLe89d5PEBoTOQ0By8xMPtqUI0/lZq
pDRsvNi9NpUk5TNzsnprsf3PAnRC1aIpPE8yumbR+wiYWCosaPmHo8lqFj6A2/M8s6EppSIyceY+
2w6E+YXldIWcO+ET6pXHykY0bD4+tY3uCOdCipiH8LZfwafBoQi1RXAJI6ddDTmTVNlVAerKvumJ
R7fxq9sfRIYgeTBjNqBElVhHzIDqRQo7+CZPeQK/mJiF5pQUJz4KAtv/i/+C8YjBZU/treA0Wx2j
M/EdEBqDYk6VQF+0Qj3F2PWeQ9U6HnBhWRotEWm4wty6fMqsOp8CCV77aNfs2OFeJystB/MOSvC6
0HdHfPmxl3E/R1V1zOCr0SWhjrxpcmewpGYZ7TjKReUmTUJGUu0q61hg1XTcmenVAgrFby286naD
NZ7TJ1Mq6Ph6Jl1sTQ3WNYiuaQC/ap7odBsHUi4BNP3hf0UQNNjVnA52gG65BuShp4WRd8/pzFrD
KXoxNmzJ77Rv85Bac8LNgKQn14PF1pY84F4diVc9Ef8/EQWhqCeTYleLrQkS5inG/k02ZRI63btb
lzNORbsOCPeMK6LADX/ffFLscT1+uXAH8IFeZzYg5lvaeAJOBlYWrjuEgHejFRgKVfJImFeP2kHA
yxXPavdP+tx5HIkl0qWez4duxSVVeo0tZbZRxSivFX7gwHHCa41FHWhSEQfuXq8uNYmvI0uHD2NY
Fd8pQgZr8GEsrGxCoJDlGTslGs4/dza5/Quqcrp6FYqsjA7wEvbMbwrNwk0W+zNas0F6hNd/0lNG
wKRa4ZU0qsfKgqmFBT59NBnb7SwSjclmrR7g0nbbV05d5+ivT4RknIKfDeA+I606QeBjCfoQ22Vs
CIjk2zVbWp2l8XyURPPgTLaz3Yyho2eAjlJwuRQomw4bzAcBpnu9cM3FkrWpCl/hc0FKk+yCT8hr
tmIhd17I1+mhVcSPQsKHDNPmprMu2A+1RHpMajf6qSsjTy6aOy3ikcMRsbkA2tQo1nr+FXXJbcD8
yijevGGyr7NpkTaQB5UCHznrIL1uMXLQo9d9e9fcx8hINp9b6FzcH8RWLRgAgIR+Gb/CJI7mp7RQ
VTUaV5X8BIP2/wAmcI4cZLEwMVJ4K1mY06lyIr68hBURvHPJEIlFK6pg+/Fh3Czrc3XSP/dIGhT5
pLER/AC3Z8lnbelZTXuHo9iLBcINLEYlcyDLxguUYhCmZFK4Dbha7ZW/8wBbSWjt39/Ya9oKEI2X
b/Adm4C7ayCa1/GszzaBocF7t+ADuKi5uMkfOuUGm91cFuIq0hfvliyZ9+2CrFFgqJdYBiuLONqM
RudZZfBc5hEvK/styHrxaEgNnQcxRB240k7KswyoFK7r3EuhD2J8AyBnU2HjT+Yqu7YolXiMyIYy
MgojxHTT9LnFPU99rLw9MT0NdbhfHcom/SXvF5YQtrNnuZ3nrxogJM662e+trafZ983hvuZs5nQS
FNdfxNwE58m4HfkcNgqyJ9+Dl2U5cB3HEwBLOxV1/XBdX6/duC5VVGM4CxV1BhYGVj8zY2DEDyqs
ciWu0U/otx57DZb8kV7iyhSWEdE2Vf9H9HcUVpddU6OxEEq+nMWt8j4rPOsicKjh5N9s+EEAzkw3
UJt1QSvVAP9l6PiLuNMUaz/PA4Q4RuEeyFNA8HUppPKevegun8kvUGhIteqJxQszyEa0MhcdnyVz
kX4kBds8hMz3uZdK66QBBYztRHDelSmOZCvY2/RUF19kemPgfFUT6vxncPEVfyrv04/byNgjHGtF
XRFZhs1BWBTettgoiLmy5ByJKRAeogLQaDOf1S21kPF7u23lzILT5EkDpPZAIxTzn5zGpv9aL8zs
8XyCQrLZefFSv226Hw7GDEP3miVEGqysjQ7OfiBO+HXxZ0OqiR+0j6cVQ0d4nI3ulBwzPVTK8UE+
X3GpWm4ctfxbiNHcqpDFTIjOakbaQu05GqCMBVyydAMHWCtsJmKKUr6CfZtm0z8RNdMhorcqmjlN
ZqhFnlf34YCKPdnHWvVyBkZ42PexFEJgBj27MUYr6fWNMWPN7RgsAdJZtUqjBGxnIct66yVvE7gz
Bfcp50SCpFMfDxctyLNuKQRLjIdHRG8g97lhk7TrBbw54wwX1ST17Uj7X97TUMjX2dlU+dJWmeUH
XXP+WfFVc0bBXFggEz3uJjc4b0MwPEhpuOBJZzc5e7O8tnNz7LRE9xXpR7KoeDrTCFe5qcHbyLbf
f4qKw+a2erctuRZ+RHvlgjaRzcgHHJ9v381KA1DIGcmjJYgPflVE3bUv+CB6fDQfmNm+b+nKdlZn
l7lvViCcXJHCQ1QtJyMy+s0IJDr9WKVop3UAy07gfJfPz1Na/bB0fHUQV1JO4YlEpv50dapzGlqj
Md6+5c4c3q3Rm606oUHnyb9z4sMDCNkgtUVMCUB9M3s99tjgU+kqfGZ0UHXQ6jtisKhCVMGKJn0i
/si5TKwvvWcMC7vK7pq/twzSQIhDwybSgf7uQMElm3UGH4hciScYfJGymABw+miN3TQBFwOsclZj
PvHTBXtO+BF2esXV6VTG0lxdcRClVbbdhZFz7xIoB/IfjNygBQ3RB7XpvFbABtp3ZnGHuQWtAmsr
tp3FodRAhbRx/+RsE72eKEMbfKzgzfyPAU27sK/lzkaiJHQ5/G6AwfZSqA500pCxroz9rQXsal2d
lNVHWIncPYQUf4TsrB16su7TI7SVBBDTkU34Ev3ozDv2qDCzNIk+9LtB14P7IxCryL5dOritIh4U
0tHd9qYCoSXQz0Pg4xy6Pj205KHoYlrGBOIqHteEeiw66PD7LBeX5/+L+TOhpIA2zGeB+fRLp3LM
tLILKODOSXW9fmQPjYhNQilhCX4EnAUOdT/+we5B37foL5HMaBp2i2z/A1jjCYLmky91tuSTD5Ks
XE2S5dJThSvtQyqnNTpNJV39gNdFjVGgd5flxCC1PFYAkDszbY+ksUlsFa1Cefth/AlQOgul3/Mb
+bBcHrFqc9pDExTfkZXpH1Qvhu0wXbKz5xm8bGuPAJ02wlunMFn4Cw8CASqWI6AyFyGryqQoiJ3h
jesWMZUTlkCwqYRrfmASqovedygdFhjtW7acVYQartGWEGcAnvt7lY395uvWo2+W7MezpSOcgp30
sRtKWxyh4vBh27hzJNGr8Z7n/UdA6eRQePKCi14GIf+z5mkyWdpXQFw079iyIEG8xAe9Vk3XRPeI
bKd4ZY9Mt9ubdL7sLyHdo6PEjyW4WcpADJiRxaSMgGr+YrXPHSc4JDAupT5phwdJKQIlnCW55+o2
8N+8k+Xa0VdltJQzPKgmtkuwm7oL23NEyE+bPpliuH+xtePk982ibtIt9T1/C/HeKXLQOnVQ0kRK
+0KnI8Qzm0KifHeZdxpPSXLlBalzBtZVw4ZoaICvdLPaP84P0gxE17C/ho5GVk8qmepNU/kgTece
OgVwUlYpt4IXIDaUAi+EVDJOT+YJl3YhsdoGc2iC1mieyzXDfcmhwOhyi8IB/BwyWCphl/UKSpc4
KpZ0YYx0aJzYJ1FnyHR8HbeOsHuDQwPRVCj7VXI7T+5E/RWW8ck48mbjGMYpMtvGzoKMOweYkoZo
Gf3jTHVIKImtCjBhYAmphNb368WsIPP2nQtyher4cFLcx2JFNoTyk6w213Nt6xaAfnU9GreWsSMR
n8GQc41K+c1905TUTZuAig3aAokDIN+22lfhiAtoAQ7zKWuJP3O6SYZNfMRjgKb6N5JilXau2iDT
mhnv6C1ta8mp4Nuf6+mTrbS8ZmrjJeDXGEi31PfAf8khr646xpQ0KtXBxVono3JtBZG3mkDOfPek
lCApeOvsew9NUSOLUCsMHaKykFlQsbpo9LdcLHH2frKleh2DElpRB95zCrYDQfZRWzY329tmoEKt
zybS6OQUbxsKPgG3u/oRKo5e8Hq4NlIive58SOfWGjW+gQ1Zere0kLeW16JLMF6pEXrNEM7/jxha
zPK+urBX5B0wbVAuxwxIrjg9Ptz+zR9jZ813dqrcSFCm7ewFdIhYpCFQU9RGT8UxCQJu+UYd+7nC
oHtRzXmAaEK2/7B15HiH6QT3GYN+rB/ZYM56/j3m8dx2EMEt8yIjitGiJK7ussl+wweNUiOsa7lK
xfflnGfIDS0Y82aBeWryjkWOJ8HKjc0ZE23HPMcZX3MUh/a6CesFWXRXXZXgAs2wu/SLvBSaJb3K
qKO2zly2u4R9ikxY0pKNlY04yFYL0vsCTYDZNY6UdJatNWxBN4dWklwEHFK/6FXCUgdocpyF7tE2
3Ya41WAaBkYmqqO9AqLW2qanIi+G2ymjQotn2nQN97SWXOK9aoqGuCb+WZaZayRkMLJDWJOOdY4w
Nfx4MFCIHR7CheGaZxH6SZTeVzFE/iI51z+SavEcxeeZ5N5akhgrfga8NNH045aJ6YUfRBuc8cO7
Zk/EbMI1YNYdlfh2B0101518wHpMYvHaLHTr082GhkLfNt5jUk5E1Q6xadSxJ9AVUkzOp0BEwOb+
IiQZC/lqEk7g9RywgS4JQz7I1E09JXA0w3l9cHE7Vrcx+tSmPEgR95solgaXJex6KV7l+k8oVWXp
awAx5MWrVAInxwzrKUgDWygExKMTBvpqnXdmxo9QXVIdWb5YO9VlcJPAeozZmfqkryQgzk+LN7OF
r0l5/lczgz7sOEUkoZumgUdTrTPeUHMvCh7/+9hZyYsupXTE2adChjFdNCuE8PTvKvz1Hx5z9jgC
/JeYCVGkhiHKNh+O9oEFAyhiH/LDEmc8zZ82lodvajBfFSMp3ObQQytbhjyHOsxICo3iQ1KSHVLb
+QmiSZ1ZG/MXDF8zQ9cq4c2UCSTb8jquB1EWF+U6HeDOxmJL+peNY6xlf/o11LFFui3vvBsi+gbn
1+w9NqgLtsb4GOHOue1m4zQwisjpvAdd3xZG0qg+sjmbUnmktHq4aSN8VlvKmo1EM5a6zOPsJwlc
lWmWNWO95QpVZlFeyCJPPxXEINPHLApmEwfkE6+HFCobava3mMgUqMRm18A6v1/puEdqXT7vToBZ
aS7QUCLP3f3l92n/PqJvINNuCBkIknMvbYkRaVYAq3oUi8gJ5R1KQkWMx4SmRIK96zzamz0phuxY
7p8bdWt4SH21feyQlMRNijxqGbeL6Uvzlsgonr0H6iJMBlO8XFvyvfTCjBqcwmwkUBk9bz3U1V8N
VK6sfX0ue5sTlBS8NYyrYGTSOrkonxCPur6i70JXni7Qwz0v2HIUExkY+wIVp/tIdQqUaG423ENR
ST8VAPsq8GMwEYUbY5haiHQCZ3AnlvDMkQqzKabFa4ZYlhuWZY1GO/pxyEZdANrOhZBZqx3V15gg
aDkj1cVymaMg6LRBpPuD/qlBzgynbERvVuwhcrFyvH4S0yNXP7GfqZxx+zSxju0hVhCibTPj3O+T
xEx/cjMnT1s8AfyYOvnj3EZTVyL8z7sIl8cNyN6CquJ6NjDlOB+9jeNuPew6RXt8dKHQSMlAlwBm
FnTLxhoAeA1cyH590f6tefj7PWaQf56Yd76RBHfSaPAFg7aON39gT6sy18Vh+x/EHm3iOTYcJ0M0
zf5thXu0Axm5c2AgUrKBut97qNeAN0FTicT/f1UrQj+KcutyqfyGM8p8Xgp0shUUPRpML2OK3uRV
2uJY5OrEoUczEFOJYTjfcl5cFRf7oRpaWO9h0/2LlBKYCfHWtt3odB0aTmnmHeyoRaAbJTmVJDg+
kmPjnreF+xoHpDyzMRQ38X9d+9LmFphZtmovjuyY5uGBUfb8WnEs9CJAal666IshNg/97NvDgyBN
RzqyKEp1b8QlFSIZnGDMMVBMamAl3JWnf54nQtkgC1y6GB3f7/27PSSKLPmKrnu9wKNxvmW4yl+X
1+sOV7fzgzAHiCCNZ6FBB3DGZxQwufM4xE4cPQ9YgVZHt9LfkO9ACki3ibmMKLCxsMnABBp6bT/L
wP7JAjVvdiVlHB6O80TcBuNf+nWvAddxpdNe16BO570YlI3JWsUSwvr1xXO25U8arYCpb38fKYaT
TC/mJLLI9AeQeE04+1TACLTTfmwNpJEj/fxzLKVjt4SEeYEdFbgW/hJAt3YEVGQIIewBXoNsgobp
gr8GcplHM8ljuWZL8/Z4pYuz+A8G4b5gY6zA4fdTprPmIEIJsaLzZx1Ip9UINe+pVXwZobrtuwU9
OxnRLs+3LjuNuubqVDK0YoUGtYbZoSql/zajkH96awdLA7shZdgzIAM+A+7EarqCgtK8/ASWBhdB
jzktBfuaRtYHQcRkH34hqWaVmDba72OuJwYaKvVqhm0lLAStIODDXLB2iXMjeUM00mT94rWUZnrm
XVgPrTOrM2VsXyfKyMjaGETMkSoip1Kl+AJgAkkjbzIX7F0xRaCakiLk5fpyiRnBEjWy20PmRDON
M7wq4O4/d3cPQFAWgOCdfiLF4fAg0s07fH8kqOpx6oJwY6iRpWgFGusefX2UMHbt8uSzmrpO/J3P
ICKveBwqzGnAUiXQAx/lEA32re7xsRZKaG2uA8ZTArSd6PGZhVzEzKkr23uO84Fo4swXedT43+h6
6fA2UmoMdvahdzpLmpbVRx5OWLJ4kwHizUgAwl0OeK1Cfl5k4kyAf2i/8ycCRiygsAanY2p3ky4L
IsGev96wzAwTuJHxSvJQtZBY0NFhBgdR3fafLSAN37jF+pvH+P7jaJKY5C45j9UDXF17UKrgBIJe
72qBRNvDpuRmt8yToaCvxH0qC9hNY+/evaxDmAHYB5KVevpCzOXUHg+HLD6pM90G9uShHkWyUNWk
ARM26mXo+ipwToT0HQyS8t5eXEFwUjqWgqsnLyH32f+orvZ03Q7gn3HKQYX82YCazrVkya+vCVcy
VZhuD6IPUgrOUiNb//PWLqKQqTAYkx7Tx0JV6+UWPfIZu+4fOmc+EP+fnaqTiuPRVk7GZ7qwB7q+
5dfxZDdNyLJX5It8dYYgWP/Zz+NrWNtJEF8c0oY2Y0hLYJXdG7HPsIaDaICDBAeUh9eYTP6yZgP+
cw9B04rd0qDkfvq9pxMmNKFrp6Qvb7wG6Ts7v4AwqcNriR/x1NAozpYhwl6QKvlcs4MdlM1NHQmP
hJOCnSwr+mpk5NIJj7UyMx0Za+aus/kqw9VJRiCRUB4oQ1tzTP+Wr/gwOUwgnU6HTy4idpa3Gnjw
5Xd+V1z7mbQnk1keL03LOu1G0eI+9Ioje7/V+rH8GNAHEc/ZoblIdG/Vb5dyar8aEAu80ddVw3ZT
uYtXdlrMLO1Z1LzrbIf/2NKnyrLYTYZwXF3GbV+Rm+gLZBN/aQJQ7p1tuPt6AiBz0/LmwJQY5fLg
yXl4KeCMtcoGURL6cknTgPr8nAAsgc/awQx+QMtDcSx5iXrUHwbT68xjWRXlmXq8pdrCIAQmDasj
fHwN6SORuudSjag1Hg/64ULRNMWeyZtVaKYHyV0Ya6QkkOM9AnfYdIAK0XSRWX2UWAiZVlL76g5b
MZEkdpTnPD1HJKWAfUUL6sqwqxCMZH0tjAYv5ehVy25rn6fjnIfMPkWJ5cqQaX9mXrpKf7q8jHIe
GV3OScac5OlhtTMmxoWw+MOtZgs1PbmT97WwNauQzYh1gkBcF3P6GiBOhjI5XOZIkGwmdqD977vJ
v9XYK26LKwFFK0WMxEEjo9JgaRyBEFpA6Q/jjkQAQw/BgvS0TYQUI1q86gmFvZe40i59fN+BNiO9
5moXV/drs4QFd6yZ3f+4QIpKiTaFffWlRDMURRE83qI+LLT0xOMTW/GV6+DEWIVh0cZnAzC5PxVC
IcRPchiaEK/RmaskD9BPdcTy0q1Gqq4sZBFKKbcXsci8Oj/t3rBkrsbuGyCVyb9BM9wUi8MSzGrY
2qa+LwJD8czsvwXoaiA60BWcWQ7Gei/epgFpXzGICo62/XWCEBZaH2bfNGs9SZYQiPKvuyXUG7aQ
UOSUkWPGzpq9GEeoE5Uhdw8K5dH6u7zNAqdbI/YzWp+iIdq8wGUo0UUcEmRIa34ylAFb9G2MhQMX
swHxVgs6bFrK4ekXi6GEnyN9mpMYwPXZxkU4lipZcXqApQbyl5R8KhelPJO4WfasL24mlXx939vq
DfBy+xDtdDc19r/mjrRgSgOdOaEqda+dnl8p2IppmFoFMOtOLe0ehRiI2tzqubvcQDccNsvyuvmy
h2CXUbtMmmCb1MKwo81zA0ab7/4rr7i4nfkWAR7t+cvIs6pP+jdqOE1kHEu2t7BwgAR6aNhZIf8r
I28KXYSb8uFF2RU3KyJRW/07N0To/LFkbGrSyDPV4UojHeGr54/zVlh0hiSaZVaf/Em9fgn8dfqs
qkK33lmWuBwGJerE7NXN+iHjKUn9/PUyju9OxTz0t3CSJQbZOzdbP2/a1lfveOKgp//jj4XkkDHB
oaGcxxrahweM4JX/2Va/+lmeCWR2zGiocPt6uQmM2332+tDUAjwk4zw4uKMkdRAPBnlzscnsPnJt
QiraLyC9XPPKiTcqXfDZPRdhFv4ASyDHP8ucGwnXo4GhmasQ2F51rRh4qqj5CmU4rnxsdbUA0VnC
KS/cTVASfVCJpK8o96vQQBoPhC5oUB3HDdZxNZfwEnO2LTvs2CzVPZYrqAbrtYgfIqyrf45fVpXQ
ohYaoZ88ExfkLCvsUKQknflqia09ymKWQycXJp63xzPESoeF4uqCS6wtcwwYSaYRGo6JuTtALzEd
QvRUI6OYlmP4ryboUamu8qX07vNa8aAXAwQYgVJ0rMjOOfouM1J36bqa8osSWRynG4yP/v42fLvr
G48dWXDJNBbrLJSUpSYosHvIl/Tw0nnZP5QI78eXuNq5JmhfMFarsTDFudINrcq4ok7VjlOwMwFt
lQPpjhZZoRyWb30ZrqWjXpIYE2tMnEsNKWD1acZwW8IHgL3nLOYaul2LAXwhiOipu1YQ36syfGGt
PJ0hnVWWzVV1SXJ+MzPZXKWfb8ZLTYBAk8mf00WZje+rm+ljnX21M79B7eW2COMoub39EeoW1qM9
QXtDczbEcRWBO60zOP3Z7in9d9QbbiKx8BMCAWKQIJhl/PBc3B8YG8KEbWSD7j/YkktqoyrV5TlV
B28mBnyB8Y6cKnkEgVxKAbVRsZf2+yJKoZOVRAv6Ob67Lk7/abnwfTZh+tTWUPCDMx07Q//dRYLw
94BiB+SvbxlOE5Q8cM1KZs5KFcLN3AUAaLKkKDIPvDjaq8CG+LSwS7C1lUsTr0JUzS0FNa7ZBmM3
sov6ciFsplk64r/ti0uBAsH9W/Xak69dWXhvaNSa9+PMp9ENqxjAIeD/q4XWfDsGVwKx6is0Phd0
jxpUnHlNz7/Yj9bVNFDKfAxRUViH47a0DAWlYwqkcd3aD6/KR4k3NtRjzraRy5Nf/d34XoN2hH/e
byoF1HorIN2OyrJLToZJEXMEVELSLNLnQYIvewz08Iny8ja9he8aLMmdtrYqZLf3rEV3XZLDotS5
Cy1kcB+qkuZSKkHpErHjyzUTZpysYQUDGbzNA6P8uyL8Zcj3iLDEcJ3r2KOrEK9R76AQlpY7F2bJ
M8w+D1Bece6ucXggqkx+Vbs3ExWFjIH3YNzeQPcIIwSUpgKFqHEAjdGDUmVhe+Tzdassb5NbdUmN
FxLijixaG2ItCZV+VOWbYIC/FyrvkFYaZubO/HMiDa2OJA3uE+upvcPUWBAwRcxifJ+tOWdy9epw
fGiTfKZbDwsL8dl6H2IHlJBN5vY6c4SpGO1VkzuUjPWvD3RpjeHKl84z0bFTrCB5i/zXWMZioiUw
FD916hwBQd44X+3rFOzN8BCeHGzf59DrsSF6grGG2IB1J51uoM28tRxDcYeWt3HqnoSYyZ29Mm/0
SpufiKu389GuFpbrsP9YQTuCnM6V11S/15El9xGzTUqMtQYO+lSFKa6+0wPkywEFi7xz5rRrUude
7gKQVf41hzySGiMR5Y3QHAeJW3xQHgeBomRlvU1dnMmvvVuNAhQsm7BZ9hKLm69yZIZ2uyzeEhkR
urzSg8MEY1j+qRNXbz5+VSD+P/G/ydx6T0YigxldSiV66ZCIbUv2bzO15AEkCj/LNsEHuh/P+1lI
XmQkJHH1AxKWu+yNlTwDHw9X+dXCp6o++KHJ7FfmjcU6lPhs/RsTHim4ElU0J7Qfk9Mv4sEoJHcv
iY8Hf2LGXYeK4ef3H8l8eJrcqzxxGDBhNvfun5QoqOsC5c44q6C/cLK404s0cPpy7lVUrVtyE2pQ
1PWmGmfpebS+SNrXG7sgR9YZ/CjfT/AiBkw2UVS8lBYjgXykwilU418ZNmDyuBFBIHoE+CQghYDE
B4BTelD3tGCz/H/Y8AKm3FsrOEMsHJTgvZFA4kL5I3XBgOUrC8FrmAcrZf1PMtXLsntwupdLRfb9
DA/6vvSLjq/iFwpae7WDIvk2y08Z2+LMKbawMS2b/pji9dK4kAeaTLSoyBJ9OyZtvCnTSwyoexRA
mpWOowXEfnU6A8wiBQkeFEdauNzYuoodb2KrNMDrODouHwQNoEtoRKqV2e7GhVvklmAYjetoIM36
Rnrz8arN50OTHgoU+4gNXFm+mZM7vP7D3xMVXGhFRU1GGxqPM9JxwPL/D3c0AQYbzjQHEbRjHp7x
wa4zywo1L8CG+XVO9EOeCcNhPspNoSueBRx9FZRCSKVoco4IYz0RAGqLOJg4GehiTQaPEdWVUied
Q1cUT1c8kEgSXukp3V2uSHi8j/MyiGSCIGphBN/6RMCsRBvboY+CghC+lSsNmzqQWyIVsxi36n9Y
r0JYROjjZU4wEXqhrn0y/I78Ti2Wtv7FlarqMevxTnk6VgraarPeSrGdeaA15Ju2WrBKm3j7oHfR
v8TBIDQKEur4WorMmWvTgiLVQiUuVPumv9XVOjl1NV/bm8ZIv6Q+w2tXhTIWO3v1C4qCjBc6HhRd
KRDjoofc6GUYnNGI0OZ/YIhYkpsmqXEfW9NgTF6Kui10u3QPWyc6GmgNiLV/GUVEAslWiQ+b/KL5
otXtdrtzIVM85BmL7W5kbUX5cYUFDb2KKJKaCVXmHFe9/u8TiTK8KlxB+X5JzG9aKzWJR/TNC9ru
3rgjonuHlPfYkE2phgpih/sjOmXOZyRgUR3Z10CqbzATrh8iF//0mDolhxgt7+cDBPwCIXYBdwIY
fOZukc2sNkPtM8yz5ZCUe2nXLk2jAsN77hVKWlnt/RP8aJEQ/qaNfarR1w1VKtWkUZ/eKGxYd96g
euKGm6HgAvP1q7Gs8Fo8ANUpP1X38tY8eJCekSld7iFHmFuaRF82sTp6iZBddo7JyZHUr8Rq9wE8
J3K3OgmvTpm0ZD7Kr/hkM5sExs1ynLojYiXbu0/MEkj451gKPeez6BqsYdflSGXPcIqIx2ag4R8/
7vYM0XEyqnn+4PL14fbhlCTFrSg25YyuhuZjGkL6fJXRC0HtKZYEzrBd/WdFMhmKXx68RaBGFuDL
kSfnhWMUKXPzG5nMR28rz336PosyZTNKZRFNjs5BERRsBxXdxdSB5GbViypH2SIrX/ZsXWLMrnY4
8i4YROqZLI8dSYKBhT9qNkWoYCZG82g/Jzu1dHaDLg2vcsEKi8GA5dUA6bpwvPi03U8XEUdLSmFq
9e1qh2nWa70lYRykH9ue7gNtFmHPDC8LftdG2uVd0QrfbaUpTJmkjfp2G1u+Y6DILwVpGvemTR8C
cVcUUSWelyUBvDR0KulatYHRWPGGWzDCIPoTO90MyRdnpxWqrSVaGxEGFNfgKNwTRDS0Wmua1wbh
SsyyApnHZWyPo2yaNDDiiWWBt/T6Jp/EMuUyiGFTQl2nJcF3lb+tP3kO+yzCZ7pG9eOLCIpEjmEj
JkMCdUMte2xXwGFtrzoEVzuqG9BRDDSb+UZcxD5j0uwzRAGKlgpbRxoA4oRS+twlIZijiGnMow3l
zfyYBdWXwqYt0FtrS70RNtTBhjn96JAYQH3ZN/wG9UtM+A6U8vQfGuBebosJf8/cb6uBFewga5JK
ingar17WOQMSxiV4W1vwBOadWkZJXw5n2Y8x+73xP7cLXEyUZG3jmG9s0p5RltUHZB7gmXYcTa+l
uzeRKjMBq4oeSclXOfVK2dY2s2YuPnxr91MtZp+dG/LPf9RtugKP6hwpzXV+dks0qR9KDw9UV016
k+SS2Ez63bcH/b6hKfLBgNOb4h4OYHLEb8T7Z7H79W6AVtZsBLCcF+1byBEQV1Gr08vg3C1gviRC
942vGsxFSFyyJX3KWe5MTK8GPy/wLihib/VyB9Ud+INtVS2IJJP72AZmzezELpM1+5fzqfXmJopC
HZ8Rx7qeQyPQl1pP/Q3Sw+U6g/qD5nswM2oDyztK0eRrR+FWqXGCrxfA/J5wSOB51MzmPtpb8VqX
LLpNyL1sd8bf3olCu2km1QaikKb7y2+coqhRYQkHONE31wDAinQRTcA07GV4vcmOKCxVtcUwlZl+
RWwZK215786/ggxVaz44xViTKgjctHKSHJ2xUdToR3Dk1t375sCCRtZN8uVJ1b/aIK3MbZr3+L+c
ZH/Fi22KHK5r6Di0AkU8QfXjojgRoR6HavMB8hUa4JliiOtgWGPvGvJRR2PqkLPNfeVzSKwmOxcF
xrerJzQyt/kgSKSD8h/3aq08UavKidKTk9LYh7wCQkHigYNnOVeoJCQkN9EDAvbCom+T+5kwqwZt
KbQ+5sEbEgdgca3JhDOLYEx1hbLDjEYEX4TTqACtUnpuEA4v1XNPSmCn/trYmjx/qCgtuduwaczT
47FezVj6QemGLnDT1uPHZ8hnMjNax3EMQJ0drMRAhfFxdqfRk1iw++MV7T4Y8qrENPGqMHa6qJoS
e2NMk3av+kDkuar3QSDtURv2cFwy8gN2EfvAfZtZCDh1Xym7sTdQhAdfE+4MdbKECZ1Do7iZF4kt
qXwrN3HYaZBcZq8j8sFtoDzpwGk6GwxJ/iGwLuGBJ/54l8hBDnVF7S+d8PocaOUacEEKm4TR2EDm
M11eQ5Oa6+QGfBnZNK4UjiM5ZpvmIHS0+VHZ5T8rcbCIe2wrh+pHmRmioLm1KxFsxK7j6h1qwRde
z/UBfU8h07ndmUoI3dTW2JKsUC/htYkuoiV3KOKqyF3adguvsUGGvSCtDIU2k2HP+9kqxm2Vkbmr
mBYDNZqu1GtApJ3GjeH7JJ7Kxk6v+H2E35GsvEdm0A4TsjSL9rl5tke5Eo5lROQ7iaOliw8Kr8h1
rWu/lmATq4AloiDH9uj2OW6wheCZNVgKeMA3LHMHcaHfrDQAg90wozIAEmx2OP0OtlP+xSNYxqOE
CLSx3MoaIBdR1OMCNgYpEom9Q3oHvsgGDnOKZVT1v0I7zGbmFBcXhk2Bdqjm6cByCauZq+9erp3v
oqlrKxOlyCyJ+tlPB3vAHZgHFkySaiQfVk3/E+jJIlZzkzAJcbCThs75AxaAeiy2VvbMWDKKtUGL
3QIviTG5Uq7bCNOoOZI9p6a5UsgmffM/Z8pPyXlkmIW09CHXNm6RsbOjApI/DmYSfPbs84s847kv
6nSagIBgpz6EgSexPvW6WssT0kwMMkIzfpMmYILsfXuB4SeyWWJtz9q6NyXbzMAYGAGgG/BtpBa9
ux3zs1G90u+tRNj1PDT6OetS0VMLmraw3sLs4h4+01ketscuKeNZ2iP6OM2YqhXDZhZc7zlpubGM
uE6VEpgTINxCR5SYeN3IMEMO7lVkxCPr4iJFx4d81fbkQX0Au4h9gDapYPMtHZN4nnu5D8UnX+wX
DM+27lmHZfcJwQzbvjBWKY7OzwCiL0RTvlf7V/TAsdQ17QmRKbSm9QAi1zZw0NtrTIyEMz8GGi7r
zZ1lZ05byKTvOFSnGQjimRJFkjmESlqkGYHfqJxsHpFSAOlT5WoeZKagZMn1qrTElkFTxgxzb6pS
JYTMiyiSbbgTcMfASp7BKTTQowR7QGy3/7TIeXkKT3l1UW/BelvE47P1nvbwmThDhd5uVqKopiEE
oyn2z//syWMMbcAxFhzzynlE4Pfgp3dp0Aj8yR1OjVgaYk9sXRDzYxlHb+xe3W3ea/zrJs7qD7sY
w7bhbRpFjBiwhPfNdr/iw/x3TxlDx0BjQZ78C6HZlwCsXr/Lu+h1svyMBUK8I65mfyPEosztxMji
jOh/hXIrhMx4CW/4ZCOeEMEndJFvVW07uEzhul98vEG/C15MI3PMCyXzmrP8sp69WT3s7sZ7d8i6
Xj3ox+EWTE+3cnNZGXncMaliWjQ5RDqu5m/mdKyVzB46R7DqU30+NwMojrnL1aLfHDMRzQti6jU4
jX2Ma79xxZV3qY4X/GuIN/+4lsmvCHjoq60X3Njo/LVXwMYRtBKc4t2LXS5tvRl0/Yuk+OC5uYCd
F3zj2HM7OOb92Tx1RaPIxD9FIO70zD1IKZU6G9IoZrv2sk2Wf3aTlI/932Br/49iGsX4iP+v4xla
60zgjIsSurYLTywXciWqiAnrngTmGUgahx9D7j9IufzP8RW2hJ4im8xPKbz+KvpQnTZ3F2Oz/OAA
5PA0rG7xwWVKERmzd/4C50LctNjAjhdMUE8Tus7/UUDm/AFxZSyLLqpQ/GfAeyYCcwB5aMpOY/DP
nxwxsFWQYYBD0RUPrxtfuBWNJ89cO/biVra7mgdeSTqatCsLLrYoCjXwH9lGlo5RqBras82ZXiNX
fYpekQEGRik0fJMMIg75q4hP9kzJzLmlA9bjL+iyryfvvy/Yvt9ga7CWsZ0an8k4c2p+ERZ1PsH8
X/ZygmXyH/BbZiOZPW51V6q0qzsgp5lcUEnKJYJtvblgpAMDMa93acPOd0aIEPjG2zai8uC5KA6C
hYhbt9hdsOUtzfw8nidUq8j55WFfzfaha//4ZYcCbpzFuZleBjp5ByKU+1PvSjoKFWqO6NDR1bBp
c3IrpTWpFRGjWs6WCAbSvdz4oZTe9d829zx5wEKODohAuIaReh3b1JmqQZXPp1VFkOsnVeVQ3c2p
SkRcz9meNq6ID+yv70QSMJT4gr1H1GMYKor+3Y9Bwzhy/DMChKpK4vhhLnKb/w6JPyXpH+YxCFv3
k1OIlzcqvqTfuNCDhDyICPQE4Vf+eE7DtHy9R+iYrR/c0agMgKayq6as/le8SC4cQ6XhqwnUv74A
zHzDVGTyunCD5xy0O/9j/12YJFZLSUQLLX+AdTm1X4ytG1vyHlfEfhLrqd7iII6WuPyzSoWl9Xri
vRKYUqd9DgNEZnGY3foLF/L0GSl+HjH63Xf+bOELkh2AVOoHsFIy1eqV+oPLboXdGiMop7lvlVwb
FaNMkAZ3yuVkPoIO4go2d1+lx4ZqHNItNdRZMV0LUHcT/JK8zoSlngQq8mpCy4hINkSFNV+7ZbJH
mbtPuG/3qtviAeBD5k6dC5Vig/rDLIq11bh8OQxrDEGFeuOfApwODLy2C73czpb3GcTNP27ZD1nc
naGsxdFMD3ZPlZ6Fmd8ZOFjfhmRLIfIfX2Agp5dGub1q6BJLMsgMqfz54Qms/r14GMcKqCY5RdBF
XJNOtcf4lS0Kjjl8AcLjqi9ulP0DTpx/dQoAfvOh1ppECuOyX1dWu1ViX/b1Mg7IBmbh0iENgtgA
HGbo2n+aixauzhfXA7iWFSd/STe9E+v3amYEFbSQ/0SUC+2RsLTw3I5QCS4qWpba3nFRjyxo6AiS
y4/DPc3i2N6o8rHBrbaiWWYTk352Oe7/RIDw44+DxGAGGqqM4ukmyWcqR1EVqXvF5QoQOuYXxs+i
qkS7FdC4EpOhKu9JI5M4t+4pHQRxU2IiAy4y4956Ta34nDIkunMpzD4lAYO0KXEh3SfZwLJQOMs7
x58PiQuogj21yL2+BZgK6ae+QjHyu1Lo0A4SHBQ6mEa3jwqlXYVTu9LksDhcGZceYlAX3sS5WRcA
wuuXbJC32TAshTdM2BleSPBYSqHzcpg+fiBpHQ6MRuOD6XFoshPPxqnFEduZYZ6raKYMD4px4Exx
dkQRcWAc5b0d3vOxkK+G7o2cs6guWfE4GL9gdxexs9aoYRxKh/SmOy00+Uainn3ia9mWXAi/kNPw
GUly5SmgbUDnbYOAmMEeeE1nABFtnc2hiWg9eZ2Q+YFordZRj4MIFMFSgolIZbiE7ud8bKE994rU
1pqkodlhNuE6njRxkek0SMnVEf97nh+uqg7K/0BhWvYlZLgGh68NnW63y4c+hMBMLl6Ip33fyNqz
/SWcbsKDQ8cFU+Rw4MCnsyru+5yCpIYmTAiJGDc9I41vyZscT0laSUfSwmw4pE1H8o1iKtdUFr81
5Vi8eH5HBPlEYjh2KiOtnZri/ojKSbSGCRbBTrnqi3MtMoFGR7aeoJqVhwLGF5qpJevGIoqW+Cmv
RpcnlkKl3yMZEYvtq0R6R2AGMa63At5oVisgP1yqtMk5Z5MGHR2JN8+TvZr+yZWcUCMqkmdf2A3v
kX06J66rlWHxr+Ja6hbDbogZ72nJaOWtxCq6fIfmd4Zs6u4BoYgZeG5mZPyHEPb6H4HVhMqCWlWg
lovI3EqB0yTY1tPEEcgO3tF5tNOI8zZBvE94mvD8J0ZaEw/uTnifIymR2wscr3hA+K31x40Eianj
6FCMo7TUdboz6MGnjGW8YNKQBqCUYZjUs9pfp7eoazVMrCZZSKD8aczVjVZROie6IFY46AQ7sFRo
QhUcQptBPG1E+D6gdNh6ZODw2/7FlCY1QqvlLSYrUaxzpaLsjrpbETI8WFE4RJDS8ebPOl6Ijrw0
JWRzA2Iu3UDoqjyExinwK+pm+O2qiCRrd98cl13FXd8goK65NVOpF/FTVAliEmX/GNuC8dY26VRW
K1Q8k4dha0qOeYbZ/y5io06fKKL4wj7QepnkgoXoK4gdRyyZDkeLH94WutR6bkXGXTg2kSDTrTsp
r1MCr1bRH+682Atoztp/L2D03dZGQxIXMuv1xGOfOXiYMnp1F+VKxafs+aRjm12pk2WYVDiM3jXB
ZsyhDzrY3D1oMKsqeR26moE0hN78OJ88373Xp7OwEmF/qm0DB2THoccA5D6wPbGyl4M84S4YEjKt
UR3LPww2UHBTOfhC4mHT2FcrCh7/is3U6+JD2CZf50XbeMvm2WUzrJgG6bWxILdX01L3Cr+9lx6t
nkK6NnQ3BXsyoHV6cCtabuLzE1WzGR7wwC5xGRYYoJskL73B+eaJFn5hioxE0QFnhXtXzN+UiCA4
3CRjHL0BcuDhWWGoEJVG5Z/gWA1es7kWcC56aX9Rs4HdcRPYne1o2v/j+xGliRhgf35Em9JWoc7Z
5lBK+Qvw9pi2+iA9O1jO1ge58ysGPGM+/VrNlLSnzKRr1NHE7sH9EtDjEU14V84MIUHp7xKA6Mll
UKYIAIPEg3G225JQV5Z/2UY7PK4819fo3MT+hMJnxhypktOytFtDAyzHCu6G/+rI7SnsNhrA8fE2
KscEq2lMzWNKN2W29TPAYRVfY0EhDOXlmrwezHZdN2hH/qO4Ng6gcyEiTcE/MS5tjv0ePWRYF2or
3z+0v4SoBC64qwY7W7dJy8JKaFFP+axe0kxNwX3vxf75FvpvYCKZ0xGsR4demxBLjWit1fJ9E4hm
nQWbggbw4AOaD1whMawNqftkG8SXa8F5uagkGyGQXczjrr4iUqg7v3fjiS/gu+XeXj0jwpcQHf9J
Pr0zi65g31esPNKwo/uJUoOkUDQas2YmxN+hlrwZPXpMvIhIeta+U3Y4Ic/lR8uevwaudFD6WKBQ
StBF1pH7Uw8iMmso5ebAzaDoor8mgrzNFvmm4FfNss9Pe26mlnuXgUUZPO40HdMbrzu/hh9OsFwi
WN19qPzjFgEzLzqTxG4jjA+fSx4ePsWnxJJ2i+3AOi/lDSQvIZqpSX3Q08IGG9GSViI47FsNOVD/
abtDPdTka6XzSSRO68hzmCrIC794rMynEco/aBPFONmL2ZJnDVYWrHH0WfvrE+oShBR0uulqUHbS
w4zSuOKO/hzUcag4L6XPkRDkjaJ8UagG4Uve49taR9bCm1RbYi8o0WLSoTN3yNQ3InvHAVW/zSLe
5eOKAv0U6f6RXghVkTMAet5LLtRXnNOzIqRgFLkOYJ07K8VRa20q3519FBOFpAFxlR7vYqd0G8aH
Quo92acj7Fo/f+sb4YI3+Hz2Y1niI9MgeuKCsLfcWECBvLlvfKRglw2tC1tX9Ctts7sWgxz+PdQH
59rA+/rX7rskvWVNUa0DK1jSr81/DM5EiKK9B+khsHao6JoFMPqBLvzBijsblGH6gCxksCIrqKSo
Qq3BIrVbOG1INZECM6dwAbtoAXQS+dojSP7tLYME6VKi2RoxJ0SUzhUIutzvq9mzG3DSF3GIvjFe
qrbAiovyLZ/VyCrzxqo5pOmIUxLIElqDpmU6NRhtJrXUpjjawP6yUa7HKgEAQSzSOxzf8W6mvcUU
731YgS4a/KnHMneAkLtRZLRovdxcApE+iykBUfbYZjogSmR+5nx1hDpr5fm1RngtpnwL2QUiE5KS
sxoCN/PbsjuCMTOCcy+avh2zc4aojV1ZbPG2CoAeeDm83rCeGvM4w0PTRYP48QtkABA0KCU92TR1
ZBcRYlKX4dUQaMLs96T2W9kK4tkPsyLEMqWmHI8/3u9CiFphJm9pn41KhQqRuPIWN+o4r5/Gb62F
UBinfvd4Rs8KhTTsua6UyMJyeL45i57+Y7ykyjF87L1igUiQ8+DoOg9xNCjIBn9HgPjFmR4QUk1b
OrBe3V5cY/eDuP5ZoWcrXJGw+AH4iF7ZjQQqY7eVE1zRPHxIHNS/zSXOcvog9PX/JQV2Bukdk6ed
kOdW2QmR9FiVXhN1LhH3hSt4PvkS9C9WBQdooN0zf/ZvmDdtXVfT9u5Dfc1CZQa+0QsPM2+tp2AO
qM3mbYrR7fDD9cHYY+6lnu/iGhoim5a9T3JLOYYEM2xTdaEmm0SXZzy8Q+uJ7TYrDYYJz6N9y0nf
/ChvatpwVc9ZKkGFMaP6gorJpU00P26WiBrGbo5zkpUw+3eqcbDQ/kCMyWvtiKrV95SZU8zAPlDa
+yjI3L/mtbeLypgpuX7mjL17Znsy3x/WBFtpZNZDZ74vJ3BC6I+CRC3M1eYcJextqZthufcKk+V8
rmUZf43T6SZ8Kzm3x2LO4LesPi7UrscLKb0RlrG+YOGMwfbC4gfkWpdzI8JIcmy336dmfTzs/cZL
H7PoLfu735RBfUobo3rsu06e7hZB32KvZvQfepOJa4Z9SuTQQuHIyZzezWivFiyVUlQX/wV4vnZW
TYYiu5Q3vu9Wl90cfNQDwdaSwOJUBLKOgcCRwHyK16MeLdkigSbuz4AZ5cWDLYycosCuAQyRaOvW
zPgys7HDML29lhfJI9FxNPQjS9wIiguSNB7c7FMDxDxn9bDVeaKDRVjGdln9uWHqch/0yTDtj9L1
esJG4LypFugVYV6j4B78gK3ugrhvEcuu76Qgd8vkUjhoEKBwtmOHfycHK7xui/uaQNygnd5fJfzT
ib5CXc5/jY5mM/XAeQ916m9XVgsjfgVnPmgZf4J+qYGNLmZZBAamgi9M7DMLN4+DwcLRcdbGUCFt
39rFXz1EabxkXZJhHy8WlHWgvD4e9U139AyzMvYftisehL9y/qdPPWj2WrKfvzuyef05Tc8u+VWw
jCxQttXtVCHnxzCgeId2DVJQEDx+WCWQC8yhMEGi5s/EB9cB93ODjR64Cve+qCSYrw+JDyYppMRf
7EPtIV4Rgoo/ZVQCTHZu7rJJUvstY04QkpsG5o6QiNaD93y/JCl4P1LQ+M6lRdsYZ34nHGiZU40v
IrFNEA1Gcq0qFY9zqLpJ18yWP13FsHr82nzs8vNTG1akZRJFOTWWELtW1sZvtY8xoHHPRnx8YGx7
ubGFfQMurfGQYv7l++Kd9eNrYzxRjLE52fW/95p8VM2JecpsOO33KpUi9So2Ugw2HRypdGZNlZ4p
HzgX4EDpmCKMCAbKbc/J/kSUmGjCc4pWy6ESxkg+QXYEBOmySu6P+jGIDqXujzclqxy7vqrFAr8Q
JScASeBqY2bVkNAz+9hL3SIhETNBBpbTS5fJNlXsdvjePOM+ksJzc0QFfxW0yRi6MsEHeDEBrRSQ
vhtn/g3xeuFz9aBoJyW+kuxBnN82lQTeyWEqelxHEvMxK0NmUM/608P7mK9vXAFXPWNejhLD24VL
fTMTgtZPe9P/acbcK5Mv5S9v/3oIK8syD7T2RLIOR9aUEAdupgHssci/fArmu3HsndzPWyD5JECL
39fIudZHQIlm3W5aZNiHWdmod4wMR78K+RHiuEjrmOJmAVjmtPzpU4wZyyDVQWCs3sb2be0IiBBC
lmzBL21Km3KgWMotyhgMFXBRTlA5HGXGkAcI5KwstuG+M0FbsXHqaForBf32Ee6kug6fqNHiWZ3u
NX3JX0Rp+9qWsin3dMI0DCwZmNMbMK8AAH1FbdmWlG1PdGjTs/x39esLAK4gebzLr1PK+VQhM/Pv
EZfVdv5uy9TzLjzIq+s1txii7NUqBmo8vo6kBP3YH2NIagYuECTI+HZ/S+NrVdRGMY8CV+Pmhhvs
Mfe/Ayrv8SF0rPmtx9DhdjjWj86kD41sRd8rz3Ptc9mKashpbUwmn7TdDE++rrKyKKGOI7tgY4fE
f7BO5Sp8a77F2Vu1qMEmiZy+Mf+t65HLn4urk4DXqNT4WTpibMUCROmN4jUC1yWr+v04coGrzCu/
qjy5Y/V1FI34ySue+N2S8tTTuHenE5ifOTkgpQUm83vaGIx//n3zsOoZzPLupQQOwC4mfY++gtw0
bWPCHk4hoLFT4uD7u2bs4f0AiIGUCl95rqqvrtkaFQ1XZeTflSgvubt1KoiStauUZpmIkbnKgu7n
X9SEuwwXQPfF5uvGOOuJHwg0kxaMvK9w4uOxJa7Lv7UbOxsxmjTU0qaH0bscIgmyCHV1vDOgGRRp
jaQXn6XlQCMoHddT9adLFBT2nqKzb2IM7uETtY+kPX3Pu+8jK+LvhrvzEtrFolsNaLfrK1TW9g69
50BZnIwWKS8G+a1SvUnJprThqsEeodNgbLjG2pPx4Ba1ij9UiY43KKLAkiGycmavEhYIJlIdvEto
kGAUQubVyfaMC9jkABuQPhNH2yzs0LMv/tWe97nFgFUJWxJEO+8ugAaSYESIbTC0j6ddaVT1J30z
KbnpujLliV6lTVQpQlHfefxRcsE8C9sXq+CWiLPgPo7j/m73+51/szSewsCEGz67B/W2XLyYHuA0
oX2ZynA2Yuav7c9/zIEhMO+wCrXfKwW0emBmqMs9Jp4T6z6AsTbup16AGbscKw/dVB0rwVnP7ye8
/O641N4InpezX9JNCZ7N0JzvrBS/ByPDM7xTcIA99okTRt+sd6BfYvrVr1kZQtIkOdr1gZ/xQ8al
ErH0CXqtSkByNr90HoFwKW57xoKVE77nPDljZUeJLPeoPjLtPwJlm+MEJJM3/MnHpzeYztHPbqfu
WgUFm6GIrrv86NOnME/KEvV0NNG5Zfz0x7p3C/0VT99ZAHeEDw4PeAqtZ3WEzppK4fdkH4sPDEcO
g2lOyBDpA6OCfBy4XwfRXhOP8yUIFXytXjdUTpaZIyXhtpJpc0Wnbv6/p+A6vmNMyJw8VapT+gbn
Z0J2rx9g88Z8OXaUKIrDEO0F7cUf2Jj82tD/2RzRlJI5UactEPJFfoMSlNx6X3i11IPCur5pfMTL
upELP0Xr5/ggh9D6B9thqwg4J7EQS+aFCY/OIblJZTONkOyvGh/W54tC7BcPACVCv/ujl06tNlVq
yU3u7HLFxtRzMoiSRKQEvpJH+R2Xk1gr+Xd2rafxaf9Z/BJOzKfX3KkR0A/Z1vBFSfGeqXcb8Vr3
tgVwBpDMlIBKtr68G4pY0IZXXmVbPQ6g0UoppOPoko8m/wgW/SzevviFjQrO/sg4xgBB73PYSOTl
rCTcTJEX3i3lx/B0jiwKdQQpaACPj9qtscJ1hOEWHbDRfhlLQF5YMPI+YHfIS1wnbihuoxBGoKN2
M0EejPyzxwgyBSAvAo1lsvG0li0XArfotNfv2VV7bZFQom9f6IuvYgdDNkoM31lhAe0D2P7x/vFi
Q2aXIwv1KVnsxqJkoP1G8zRiPZ0OBno7sWkSWEbV6ZVuOWo0hBO4uM8xi74qXvjOV6t3KU70blgu
YPes+qZAbtPA1zfATOKMYLC3ORZ/zV4wUIVTOlum+2EfsTIvLPOhau6cc0pZUU2mGzzNdZUWl6ys
1HSUUVS2X+Ftg9G8dc1bg1o9jjZbsMYOTXoMn1H8BbkqVvOaYzXr/euHlVEBPRNxbrpe/6emz8i0
57bPQY2xW2FfSWTpNJvwuL1WwkPVJV7a85ImZA+2hNwqph1DwMPOZdD7L9kS40CfKe3FdVwNOXQo
SMu/sGM7l8PfTnigEGgRa/Fq28mNK9QafhLGbrXhWyh5mLP/dO3T2HROLYVerfEudTqRP3yS0n22
yyOtQs2ldKZICTLe0dGIb6blyDNdUhS8yjXpBEqQftJudcJ+t9+5zDVhxhdXPgp5qXKYXmsnoxzd
hfYVQ+TY/i7wC0GV6Fjsrj02ZmO+9GvbhQJlT0bqBtfa2TiTFEKbf6HPWyBF8NL7Ya/yvGOA++GE
niR/WwBFhyPKInNNEObbKjwj7T1a3lo40zm4V9CswC2BDNoFkFLbA23NmnhZX6pc5qz3b08CU5x2
JnlWibxH39krhxp1l35vpau+euVn4OqHexwNLMPJNsXFSYfJ+VJQ3FyKzi8/todwoG9LSGRp+XQz
NJvsX6b2d40Lpkpmpdzh7zoqLwMLpeO+M2sr7pK7Dg/OcW17IFbQecZeL3ehOnEdyjRTOR6nzrMc
zUrtrdaRfNCbXtqgvZcfB9f3XCXK9qcPZmoxL9g3sXdFRKi2HQqIOI7pil/xwRcnnWhOnl3gNtBM
yeicG2wf+F7rbVC9BCxrGHX+og7FDdX4JspENN7kHGqwrcwhZMf3JVqcYOXdTkj6tnPgzCCr2W3X
6F9i3d2vIsGUdY0/UwBfJHm7hr7ilNtGCjUz7rSz/OkOyDLm9/6pQ6K2dRvUKWdG3AFnS3tXe3A8
4jWDMn41L0vaEJpXsI/jvPZsEGDEgK8PhNwqglB5PsCMQ74pHEsdmCoJPxqz8sDwr0j3Y7zwURN1
t8FMRPWQVkLetXtlUKVkOsE83M5OJn/yDQu6cCYq58TqvzjH6BGSuywtUurQHxWJpiuzbvC4w/Iq
aCXCc4DtIblrfWDMX3dkkX00B8gt1fNqyCK58HVCAsYqcFaG1hYPmaOU/MOALW1GgGpI0FJkcW7W
lkoj7OKHygbt8gb0df1AEEvDpnIWOHUXHKWKotoBjV/K5gc+WYQ+v/sJp6ovNDcDEWtzXb0Fa7Ue
68JQoIAmOXlzJcLidAH05vSYETn3/1F/yP9a0qSyCDhP3rxDV4tqktONURlhPHM45Xx39eqH4gNQ
zU+TxqHzoXOiCmeVrd/YWZdX89QHGEhtfhCTQAXJXIXcNS2ydqphTdcqLsJTvy0VPaUOeUytTNZK
jC7wXgRVlnNIfRSgDGaGbZW0VzpLvq8KOKKqAC6K71DIe7vXKCDGh51jIAbEddxhAYEDU66xkWEW
G2rcs5hxpCFMfgVYXKJ5LUtsQ+cC5RR9sY1+IEyTOv55IPRGgmhb1rWDv+5O7nwHBjhRtUBGC5SF
Qp+Tp/aKOFzaV6zDtkv2mNGFqlmMc3Lk+v6y2tlOF7LgggyfdrwCxRpATQ6yKrGZLLh7IPkJ21kv
IJ2a/L1Sf4sJCx/ZgJ8nwNJ6AXbHNBxfwhXnYvda7i3ZjOnZN8uLFF4AeHMZLH9Cuf4uzPz9/EN5
d8NsW3p+8TJosbacHDtKVwiO2wz5H9BoUun4JGrnvQZC15V3CRRS8C6Z0KblZGdxnBH5KDSgdEFT
o/OJfCGZ2AlY1fMtcdEfTmmL75JI6rMy9lc9VfmGzAaBfdDdE0X490HlxUXsru5Yz0B/cJe4RxSM
dVLthU/IUdFoYfn78A0jBEfhwRYoiXTdMl7Tewtqt3Ucco1snEoOuUoVGdxMUexUDLdE0GEQaXEM
FxuObJFCx7i4/HejIrWdCtPp7faGB4ahlxgUVprjCVOsyKf1eRkSizN68QsPl5Wgf9uodY+JcPef
kyy5Tl7DydZbUoDJz7o4AzP7jUQsk810XGru2uqLDWBxwbEOkBF1h4hX+sE/UwQmijnw4mEDP9v7
ODIZbmVHzL0U6cBvNwQaaZZFEvzTMxWVZAPZjuPKw+jnTKrXYGXbRAn7dA9JS8ZOr3+s/7mA+6hd
W3Jn5nyha+yde/9NY7OL+XeVprIHdjChomBUWY097+HYMgMF9ayBTQWaXjanFEvUjZ2SSapT0g86
BOsj6qzkN77aEtL3OajwS7NimV7yZ3CWIL3b9HB1rimVoIhX0FWPLSEDgijXlc/CncwSfLo9J9G5
YMs91QsDALlQz+Gvm2L8PRXQjC3aeOXHXj/R8ikGVxGVKjPh+k412cYu/sbWk+hAWN9fg+P9lALn
ETmmB4ejmq58dc4ds+7lSUjICvA0g9OkbB7WZgaeMlLLT/yYPNYjHp9FnEs5uj1b8ouzvQgDielx
vT8ml2qeov6aZv6jGprU9CNF2pFIBQhGJT4kRsunpN4C+F7UqI+Duuddrbq3+zNhjqnSvC7LYE4P
a2lxfWBJn6p26nKooSkxZk2c8BotA1QmwUNPNEXxBhx/3a5aO7WYMHP63QmCIaVzgMuXcSowXZva
hL+wTGl3JBqgb4CCFrpP1L5ND0vpBrMRCrjQDE6pknn07Nhl2xqXwYnf6+kmQbILTRkJH7ARFJmR
N1sNxQh0ffOIXNMimuhM4EE1fUGjwGcC096tGhLwP2ry3XVR1tfmkL6lmhPIiCfMkLU8jCLhFJNj
+z/P1Rs63qlLBs5I4/2MkT1ggURmumoM9ukZbJgSNylx1pkYaFMkh+F9jk4BezCnKCYq0wIfvSa/
Ltrsmqq8GDmoM0SEOQrgefmjcrgonddjFG3DFnie96guVVSG8jXBlvTTppSJgIG2M3klJUJcdoFo
nOmEXB+ZJtj6TDEtzjyCcpMe+6qJOtdriqlkkJbtQ4lmkZY1TJ+rVa0LADeuhmulfi//sPEtMRL5
eMjII0AjtxavnrHnfsu8fAiDeMEF8nqW9bhwYR1yL+yHo1xYsjJnsIW+Q54nNMZbLFPcHDm2QwLI
FmGdAzOmzv9ugUcv4ExHAyUVOVszN6I+huvbqHCc76C5wo2c5JtfTVJvSK6fC1s/pjlmFUO14hcj
y3sC0bLgaxLJXQd2FgS5hgwRPRb4fWOJGsfhbcxDy8+/CIGUw5rCgvqdtyazzGh+Uua3m/Wit1Ga
RKmMC5MgK51Xhcuikngbon87mIji/dyps3q0bzCsu4Ao+CsKqUJvgaTY2LVrVzw+kibGT5HXmHnD
vnwEQZENjoAds6COVuihQNY37vvsAp4MpQcSomtYy/F+RW4HLYxRoaKmct3+XG57mXzhIczC7ifK
1LII47d9h2JJSOBcWEdy9bTiaIAgTpXTyUtTBR12mrupX6YlKk2TeqlILsupC59wvLluqKEcmz2I
8rfU20rT2Qz1ge3d96HxJMw9MeP80W57h95Qo86Hl1v5mN9g3AAjmti7tpYfpsLm4qMf+3Ta9IT9
bzIrkVekNmmMbFtXuiqLBrHrfNX+W/HaNVcj2refUs+BAVg8QkhQruiM3YzNIPsskzsEf6utd9nv
GsFchDpQJuyMoOvn/EewHlvihEHrsQwGH43WOZ1nPtSlk0ZTXBFpsawc5JTmt1tyZZdnSPo4S/aP
Q1qObijYOJVBBemUd9pQAGFMBEKjGpgtPygNNZfVmh9Xs5hGr9dvVPOD+WXmbHoU0Ze6RUGjY+ko
06JyaNlqxzCTffoQX3ztXZQpS6jPXJuQf8wWcgoge4jNqtwjkz4UAhmsyHWv+5RDEVqFyJMkbGgC
jZHLXvpzdbg4DpCWRhjUIOx6TaMsS9+tNjMBiQOY8ixQS7lYsvirJZ66WPiZ8HzK91xtmYtUi7Su
G9dt0+QWYvF0zsujT+tzEDuXlpXIP3WDk5cL4luQUIDTaBWm+4YCIrEefZEJV0ZtJJ+mfoL2HTMh
oPf08+74XRp2gTw9OkqR5OKWjWc1FARJz4YbiGzqpuYpASglXYsOqFMLrt3HsamBgbg43mE9JcxL
diWy1uAQayFBDrxyHxsk9eNqTBLFmwXUEaDAfvqh4ooNTjkyKvhbrsJgUVLBFKwdmi8uKVqXLNtE
yyhY8vKO+ivTb72DwzYl0rVfFKQorTvXjii0xkRk8BqT+3BWC8XeEzLvGANm2AogQwt8HK534D15
OYePJgpR9YppYDWOPvejHT8485ULSJuma6OFGSOIFB5IrFN6+RhaJARLAy6rQy2SePXALi8+7g55
fIa+E8g9+etnvONgb6Pvzsc3kLPEBLqLgrInnuGpJRMTSN8PqJu8nrSk8jkt8a271N+WfR8qCjET
ytZJjdyx4cYTVARHNaOB2zGjYL4Q4Fy0VACxPaD/tbnUl3BfjLG7XfUGVOTqpPmWK/GAJdxTZN/W
eC8s11uifx2qQTgbX4vf/mLhHRdf9RteZrVJC/PqwqLw4yy05AMHF6Gon99fUzYTLkzk3asUrgjg
/c9iAtfkrEZWDPN/fZAZ/n2rB+dgEfQ7ImwNFFcdxdkzTwAg1msJdWPHsLe3hrTfyRsbUgRf4v1v
3b80+FAq96q49HGU3WS1qJsLb7LRU+RuTEHfxB9btnYfUVwTjoS7EIvJPa0VgoQqfus+OHdJCSDL
nbwqqZ4O08mB544u0vIfwWoP6mlYSHeo961N4mk1swARTlthuanTQYPT3mVphpEF6dxN0es1FNA7
ykbAZyN/aZOLC6po4/7SKcyaY3UlbOk4b5lorr85hyRZ+RNsbPcsLW91CwjtLJkwp9kcbyMm8YWu
uKwsTsSHAD5gfkfRyk2fY2fabVuSqw4jGf4TbW3AwEwlvZTCHREAeaPkVRMzYCnj6ipKTwJtGFnS
TozP3NKiA/Nw8MyeVZZ6Z+V5fCeaf6KPPginM1vA0WYf0DLQQNrn8yDzxRqihfcdDY5oWNjxKlsv
JDTYBgP6dx4fb4FUzKgfioFG3JICAJLv4Cw1gHtkAk8AXPcVRzSGltxDLxEDXeSeB2h/0umoowHA
YcqgyjC4hnwj8wBjkuoYuBYgjsU0NRQ48nk/DyqONhGnCp1blsMB6YomcOYkYsGhhx9ZqsE49oDd
hXsrNWbif0HOPCTNTaEKbzHFEq+PJKgGJ4Li21pFjMgXlRDHdBod4LO86wOGpCxIAUQvQkXg1ufQ
wivC2n0X8AkaDRJQjeWszCOALTPqtLcmGRGe525g17nKDQ0FjhMEhtpkp2S+s2Nzy7lp0/PAR6fK
GdQCYvJ5xGY0M2wv1FcBK4WSA0mCHcxYeEgHxcJ2LVNrzujzXh7rayeT3WJ8bG55x7h8XAumt+5U
wZZyWzeWsPrjeZfC+VswjpWJy5EhSPzojEqCskHqFO27Be2RHzq4QGpHM6xXW5WAsfJ025fhBLO4
tl8cMZh31qww7CyOM1nPYO0DuAFkrZqMzhMZNSdk8az1K1lSJH9IlHL2dFZw8Y3ozwRiC8Fsj68c
wii+jVepPndo7x7NYEUU/Hv+Y/mXiWiC1lanlf8VinsmpzdGKWz/V2OLonCPr1pA1syfPjhixlBL
/9S5IGGPcHSrsNKl19Qj5QBrTFSNUt6EnxSJt4U0iIC8kZECTTPzqKOWjILbeCVnE01aFv6hsGu6
ub6Oa5A7++HW2fGn9OqxUSO7Jnxp2TCTjxYh9Or4M7Uu9UCyoS0ltw4aUUN2Iqv5yvy7ezK/a49m
6C9R+38SrgwwKo/z72vHyAe7QTLgRaDkMHt1ymkiUK7e8FOLnFb/EULWsFtqwi+zz0hw6KmAmjjm
ZkAzRkJ/BtU+TjstMxM9/kxB9h699/AKcCtoyHB3xkCGqLrulWJhiCmpX/hEbrHsHcQCO/pFkLFF
jwjySM09fk304BEVUf8Pbln7vMdzXB34hBNzSAfO8b82hbl+bhMD7BrDNDIzZDycYqnCN1yrInG8
KfVm4imD+aZgzED5mJB2q8mO0YWlZ96JjdqOCK0JVpseXEWZWvxQxX1AQEyMAMTLjADM2k6Ff08J
dbP33+dCSZircEXuORFKGmKfHV3IHApLbH2Bzl0bvsJ9iZOZpgq7Ic6nsEitPFU6otOlCUSMKJDL
/PBWBmIkRfsn4jim+2pzpVUDdijyX3qpCT0KU+vlbCq6t2/pdHFOWlqyMtDR316b0le34dqnVSnh
Fh6DTn6aDuKQKz1eAB+OxrlwF8FTMKjujuLBdplDMWnEJMit9n6CdAyo1UDyEQ2QSclBNaP0B2iN
x/Zy7kOoYk19xwVqZ+mMXwDdK3NqoAf7XDYfdzPB1t5zgDgS84u4Ou56HrQQwMMOyIqcxPe0/JCO
XplTWUe5Ih5iu4z0SFWon4+P2RAzThj+tJK2bcxrOwOjVRO3DYqWXQCmPSvoENBwdjFwDVCKQxkW
4WG2TGKzyfeQAPBXsmD5SOSO4yEClidlgXE6AA4azmH6ZzzIHGZlABdty3wxiv7mDERjbInJFgRN
kiOxFA9Nl+AyaSEWFX0wN/1oNJLKGS/JXFnfQPxtDypSvOtDERhqrPnTnRZrJjMXh5i8u7cvkhX9
S3HzRCFSDxFzCMIXp/Mfx54L1GHc9z7muXaBABMeqQ8+ZFvjZOmiM8r9rh25lGMleK0k7M0Bs+a7
JJLuzvxbroNnsAcFqKTIhJiY/IMqf2dPODpMoiGQTwawwSWaykgZsL801gA6B3kS6A17E6Nwp/u8
/qUq+tvPGNj5dnJcu47RUodjHjQ/MqMmnYAAKuUBpzUT2p5xsEt/5WAClyogVgTP+AL64oPQ1n8B
eXRsT/UY/H2ztAWzWaVcAUcjV6cTdsQCmGA7BqHeWzS6bKxO/w0572cflGjulToYEE1GKGMkogbx
BFesn7mtfGii3dhrL3xJnPhgsnybtmW0RhuyNNeAGEki/qZm9hB1pcjlr0G2kSGu9QZylz4z5yyD
DFytYZdC0xKrZg4Vt/b+lzycBlMDz86fTAMi9Sfs6s9RZtfi3rZ8f7y0vYodqsfoIy2iWdV533fZ
PDcapVM6DGQIf2B0yU88q2mXDk+CHqKIovuTr6OYexD+GmRAuEaOaO+8vlcrdBHlFrvM4RDmeCce
mrydcDauISPBiwsPPqJtZi/2ffGDYz6h2BWketqEO7ZVEm3sMjU+Bz0AFUHy9QuXl2AojRBbt6Mx
Yzrebhvwj2rFYtAxvind0nZd8FBBkd+8s1VWCaBooHb7VMGsrdPwWPHlmpCmC6WrMmbAxy7H1VHB
GZR4FbLPPbfCgpD3W2mcV3Yhj7TERNwqsKLgRvIXbgy0i2FXNAuC5DuTrEo0HwAfUxVqNrjG613+
2QO1fgbGLI/ueOttlZts3TuAq9tn9Wv0gFZHtJc3RiuNUO4jclAL+TNTEtSXztb/Pb9fdy3IxIIX
lzmn2GC3Ta8CPk7wZ5eILC8KWf01BzYqm0bjcQ7dZoBM6IURsCKPXEyd/ErzZawpjLkXX461iC6D
od5iDB25fXS0xZngJ4uzNzgdOu/sKByDmMI0b17qiJuyNvR39nSXGC0sphmlUcZnfzraz/uQpVBG
J19jUfW65GfcTxEj1D02J0q3Dh91yh0uLdO/l+0m4CrOs9oeJ30cQh/c/7hiTlf8dhK5+w33ymEO
V2eM7bERRpch/kshENXFFapnleY7vU5YGV4ikYVZn2lIregnUaOirJccvjk0s7YswCQtxsEDos+i
n0oYuWjCcBcRUhnmvHadwZZld6vVTO7Jtqhe5UWds3uLTKGJEPfk6iDg6a/e/2TmIrN2bQMI/i8n
p4n7iOMcElFQ4pEoM93sU1LrN54iNZxmkiYAvaTTeGzzm5i2ThiXgJrJYYe7no+iU36VQll1ODF4
qmsSh4CIfPJ4N731q0Bl3gpNzvT5+5OP7QSh592hCR4/ZDWa8dUxJd40or16YMmaOowitK9abqVT
jLTeDexvjxpx2QrgYsT53hUyFxhoJ/d+kIaiAvpRcQCK6RVwR/y0piqO4plitYPpYNel9oxTL/32
XhmZCeJ9IsG3IxzjfPEZri7kuJzyvXph1Qs/3riPbNyFNkBnLGrf9tYzwrnhMT9ojAEgjDA6rUv5
nebAa/ArLe+C5yWtQStKs3s9dWcI20lWenF6r+jY7G6wKKhfnJdoxoaGC/rVg6erT+ZBfKeNjqb6
FFao37xrSDTG4+VUBWRRp9gaonF/LCCQ42fTI7A9wBkiftYnjhTGz7FxXksXemMGCar3Mv7kdemf
1PRggJF0d134qTi2f5zlqUCwo6rV0udvQ/2OAWUfgQGM6gCef/pt/e6nvfhiiXRV/5UMZx0QvL2X
ULVwRzOVb6m6ft5VE2ReIpFpxZAxz1Y+u8O+lBlAx6ZASrhZueNYde89S8/d3LYK0jj+xqLyN9eU
0rlHT/jD2Bz7yiMHpbsNmCz4LhhUZqbmvGWCumyQSvACwfD+dovAiXNozOLorfvXyGewZFn5meFL
7WTEE2xqYs/RChMirFeCiupYVJoZvt9QcfUE7hg2l0iNkXqhSY0526OojSciPCkPi/OIH39M2g8I
OGpgtiI8PW0MxGwqrVS9l/lo3G8bBzVL2JVxPxUvWxGBVUpappDRGtwoHD07J1kkUFxnMR2zSxsi
nDkJ3/cNQCwawuoxNylNbMdHiDmJVPEXr40oB7ZFg55oEDkSzS0+FpAYs38AyYp2awD8BwwiBfK3
HZSriuCQ4HMsQoFxcPMIHtuUQfj5RL06THmN8IIuA6rs5vwgKH1/3kfEOUCtd/XecTxm+HUrPxld
NL2CG/w4kPmInPlKR4DybtT8EQosFQ2B8zmRaN+KfCfbqJhvMOt3faa9EA3tV7U+LidpYOTbVQmC
k5L2Za7fDKCTomQbk6/3arKb+hvXtsesrv7C3VX9IknutfjjZ/ATVv950FrPWsgcbp1hwuwnAiU3
gnKF2yQA5qBzOBoxqB+b4vSUUm+ytaNPrDZP24Hqn2VpuyGZzmwGt+8hA80LCcCUoyTuedzG3TvK
H5XmHO53BHeI5HNe0v6ChBoagmOzOXBrN69vTr+XkZusQgmhvStMDaRJ6iYk4dhYsHFMlBBqOlcQ
4QjlJFMuMYWFSy/X6CkjM6Z4Tbkp8lgkQoHNJdxjc+cThxNbdBSKo6Ap4/DHUJq28t4DVnbCbC99
7OVEYCMs/azLEbC1zpQzJFWoweM3L2keAARPrdt5uXzkeOazY805PwnbDhbFWUi45Pkds9xYdkUd
5xbuzagA/NwkmRQIT005BencdYmKDU3hsmvA/stsUSVJwJ7M3++HNwj+Ed8odPm+6S0vEHIVPXhP
YKJso3HzzmdtpmHrIDVqE6vKVfxgrwRZhRHkSmZ1xPwCqNOgbmXeLUbynAJSxI+8LhJhmqIh9+5F
QWYuXUDN3W8U6EfQ3b0QUcoBxITXIKnHs5jZ5MIwgakL/PLyZ2JbTc6LsBn5+SMmky96oLX4g227
Oh6sbDRVwgtWbkTGr9NQ/uNaSo5wjDs9V/phwS3/JBENStH+0sSY5GQeiirqokLSsURjpF2V6+aB
/nrrQhD9gvnH6PE3a0FlT86QEm62n7pxrrDQaNIe9dqITDS1UCnuRU8RJ9KfmJH2jKICritGDF3Q
Q3IwX2eMPsMrpvmbhFt9pUDSX1N7YXie4zVs8rKF3yjMCzM4+qV4stiyoY/zxMjQXxOL5c0swyY4
eiUqL4WGlCqjC3FjUba0lMa5hPY28n8NW3au691nlxP+LMF3s70v7kus3CILxavvImX8cvJJY93N
LSibeOv2HWmi2tbeWEKnNggs9FikmF5bGDAcn73S5oTta43lCoIwAwL7Bk8FPliewWJelHHJrvyx
BtQEt0q+ybbXYf4uzqgRTdvwXUj1rdq4XkCMcUWCHbBLUC5ckXX75TKWvwhfrGllXMOvx+kzfegB
i93yw0piwxEqlDqsxgepJV0P99LOIf+GFeQ+OokeeCETp/JpcA9lOFVD+Jd540pU6qYZpJpgpvj8
V2HlMtl90LpNu1o411cauSaT+3GtogSTYAq3iH0vaoZZdvGVFgsf1/oBwN9wnSERqqb75YGp88Qe
u77OrL9+vaM7weReIsDkVtrcaWURQp6gWLC0T7T1+bFUixm729ZN/Xdu6He9Xv/mL51QjkxDvD4h
ieioeCX5HkcUUjoobdoqAcsNCuEKmMgVMPwZlEVQ1l6OZ71m7IYUg3JDdWXCJ1mFju71bQxWG8pP
/weoUuTQ6i9wDmiIZI7g/rWhw+WSLfd8mK2uqwY68y6dVlOQhRcaIWudDuDh0OE5P1dK5ScuppKV
08N7R7UJFUa0aK3rU3KkpINb5CD9v9sBt1dUfmhRfirUO9ldcfkj0MvDxULQMqg0EBtdC1vtD+wZ
Faj1d6W3fETp2JHcuwr0PQrx5A3b5x3nd1P1haU/QIQm76G4a6ZAEF1qFEm+JVByxGUJATDfAH3C
1a/kdKInu8F5f3WVRMYBz1c4YgsUB0OZ6oHnlIk4QCzuQ8uigNNI8/e4T6pktqN3HX+z81m5ajyt
yqn6or33fSBT1KYYh3eeP8/TlShYrI3kwy4WklApNLOwp4x+7vMvb0CPp61wysXVOUX4cMXxxzsB
2u8bEs6s6nP/OwaSo6ZUMA8CJFZJNz7jaTHjPtasRiO50TczSCMKEDimcDUmKBVLO27qvAqxDVN1
V6fxZmZXUgbIRjQXesMzJcz3Ca+uOjDZ5fgzJ1MfBCXsG+++k5rpdK1yqbiS1Pqrov0dg9EY1bjR
r+VIUVvTwwyYz/e2r+Ifv13LzLawnZaroaUHNiyeurjU7ktTdFUw/6E75Hrl3hCa57ImQ7JRAAUw
6Hvfb9qnrCucVI8mglQ4AEASj5UCpMqm1HcTWJFUh9BIRWbF3W/VrWdEyybjJRgfSTo6z7LjVlIV
g6f3iuQxRTvGqsP00KpPyoCDp/FMblDY9HJXKeAt0PpE6m5WKtfqMfLD1gEpH17Jgf22QLg+8ykk
jh+UnDK3t+A5I7MuLFKwmVqgt3XzSWb0O80LG7wJx27yaz2yNhBUinDWfcGQ0g9vsBOlYv42Euh+
vpS3sVprkZCsLTvsHeTUunzY4amjTbOy2ixgMn/g3wJE7RC3C9kGsGM61N0Ewg34UFgSlDjXW+mO
ylofCKC3k9xIhlP/5ZTgkgDpcmzeEgrN/QwWUjz6oHLLXKiccWdJC+doN/CgJ8ltcM75W0cb/JHq
+UmyB1rGQ6zKjH4MBSqolVJEFU4z9/eUsNyX70/dltvpD0uXLDQ9IdnKNK/BrIT5+2Juhdi8l8Z6
07F4r927yep6ElxIENQbzVpJNC5uZjzlY2LWQyz2SV1DAnpUBagdz/o5LYBr3bHZR0+d8bkrF9QT
S5ebB48VjtyzyBOTqh7eM5tyoSE7riYZIUlhwGMb4X0lUayDP848N/Qp1DYmPKK3cWgWNVSWgfOr
H8VyVtLB6bJLvKfSde0ultbekkeuemIiWM5nslv9lre+ewTSzEJtwEQnmcnRFrwC8UQIchFLSzfn
y58wbb18YqYKR2E7kKvofSs4KUi0IDq2vXqefopgHJShfvGXC5KJQUaPHcy1OlPzR4ESW1iWwjGT
nBN1aDRP8gUCO6g8Kw/MUK4Bzcqf3lcZ88ZjurArGWhCB5xowKM3uwYtAeDoxL7hX83v2ouIRKfP
jDgRz/MSc2Ir5AsHqi0O+5tV+Z3Rq7SXQkw/prQRX0DqODAELKI70cR9YSg7uEd2rNbyBKSMK/NZ
Hl2xR/M3tyP13Io4ByH1cIqukauiVjoeFuNql2vnGqz1ReTn9PcdzEP61MEouqEIBR86l1OsOF30
F547TKGtbGlId5Uf8AgT6m/czLMpvXxrjoVA+a19EXxUtzJnoyAEsZpbkttqNLJ1AmR+i9rGNaVK
PwQxI5kvuvz8zbvLlzgoN5ritVpm5N0BidUp/DYhO/tyah3xp5y/FvGiwc1pBXR2cgSXzrLWvI2O
75kFUkvIx9dIPV15Es5cpwa3rBagWH6paWAtVB2phSHn+2jF/Q3vGc7j+yuU02NkUA0WHr0GZ1UG
ZbYZLj54MPU0lDWSDAw1LOP9JwTxaTATZbxnjFlRpFhlOT+MmT4gLynZbnDDVPx0j6VbpwrcYVi3
yRnMLlmN89Eu95x3ng0VTGQBqG70VsBcRoZr33HOHXc2hUhltMTqFrRHHqQSu0D6LhfjknCWfdD+
+SoALcq78zLZvIqoBDgTSeNERUcx4Cxt0/vZgXFQYaN5IjNOxz4Eq9FYef+LFYnAHO7msdEhIwA8
o+Fvnb8LEECAdIWB2H4ELMNojuoW8AD6XNsGxbFNium77bcWLtkYchfMDISK/ymYOhq38AchfdLJ
wwW1SNTjOymYcvwLBTi8JLRu3LlSQ9hipT2G5EFnnkuvPJq1kJIX7WIMCO67nCEe3BDx2G+24nln
keNBtqZ7dVkmsrgujnOVx9gGCjn7Z22lbYp+j+DXrGJDPfYDyCy0XfCZUqx0wvQsfgtd84NvF2AK
dSgGA5rfRRMpPjhkLhTYx70BqYKsAal0Hz01eD/PeFoBwGmuAmxlsyeN5oxbM/29NWxkRQ4JVw2b
jfGPwZvjbHgS9hCLjj45iSQkz6auW6BXEN2LtUlNTDOIDB/X4R4zwhZdZMVCchTcc7ba4ySGSeoG
mPtKm75l0WRZJavYoUqSZqqIyYyCQc48Ahd7HuMX7RT6jitTDVDfKH4edz4OJTq377bMNJ8oef5t
7Mf9Kj9VadlPL6Frs4Hz1coT2TR9bwe2pocx/dkInUFQoXz1mEpYrnl+0KtcrnkuhdvcEH2tfnI5
/PCPboUfKjCyG1L6BIkDnKTh0krRsRicwosdrQw5Mib09u8Z9QOxvmHLO7F3NfO1DFfn18WLXEZN
+136czp4ZSzdQdPLMgSVYTRydFhYm/AJsyjv2ppK9AFuQepXSRBCLCPXkF+rZYTqHFCXlx/L5+UB
kiZRG5MNjGjUtDkYz+OyoTb45Q0EQvidbWTo5Hxo0C/VhNorjONA5M7oVufmsPVDP/PQgVfGS7sZ
sszZZChM7Apdp4yDJlAnnokByUT/fhUKFxZiAvxMSXx3rMikNygCwnAnZxTkvefz/sv9cs4V6iQG
tV0ChfGy94Prhe5QBfjBzVCNE1jFL8l7UFEOlIwjU56UzfqXtnUBtaUheZd1eUvjRJusuGCmynTU
rXGnIUjRuAe19ngEc5rgbyRFxPDezT7fJfVxnIgKSGuFvqxFpVOBalL7+fL82tKokultx5GeS3Xo
V508AQQ9U7EAOv9FjiukDffZJUp2ly8OC11FVi+btAre0mFw+VC3xeBapUOtBtgWF48vY6K1w9kj
LGLn7bun/mpFelxykMQeR0N6H6XkCkpfrdFtgmXg8I2Ptd9FEw+tY59hQxRjPUDFVJazt6jCZmN+
b0uIlTKCZzlDZU0sieRcfXAe85uJiSRAE1n1singZ8ComQe8XzSXbqBd9Di1XaaOutjHVUVon9x4
CKNYIALW4vfYKDtVoYuIyrjj5G/7bPI4eEacPuiReSRwemkRQ5Vo53YD7AxWIrcEWVyzy2Z5VR8R
QDTz9u8ZgHzNBW/8EgkjjkC2v/7g709HNuYAXqWsAVDmvXIcejrXuXfqArLR5NaN7EWdTCirgQzx
vaZHzNZIjPDlEm84MoPxQXVzyM3RUhJcWWKmgXJ/0/yPzXWTXxWkw23yeYXLgOTVG2jAF06KiyGI
sCS1fpPWx1jN+EPvk6YcEkNlZl6W9nznMOeyM91/6tM9SBsVFS05Zyj70tHHsh+jRy6JhNqzxLbe
50UagKEcGGqkDONaVN13Iw6Huqt77OpgB708KYFyyeHnq5hsiYmQJ/Tr18oHfP6w423Nk1YlKzBa
spAWHCxLyouKEUQf0rLyWSU724V0lrJQQy9wXofKrp/oP3W3g5naIIB/Sr2d4qSzFZJ/dBvJWOtz
cnOLsOkVTh84LbHLqlIo93Y3JYAlOWLH3Nwk0mWJYEH3DrwZqIPdRFTkaxxH5TsiAkyqqMXCitqG
38PI2zDFUlNh2Mi5GQLR3jciVRdj1LOImhpwiS+as2i7GnakkVgjVjqmsHmqFy9XEq5jfSxBjoSI
dg1cl6Nhmv5F/rh/kBFzoR2+ywCxQWUJoh7g2AuSrl5ZuweCniIg4sDGFw/pswc/I9lHMhhEWvAG
xEdHWP1aZED+a9igAVnibI4rZasXDKcU+YjF895w8dU/BD679U7tMobSVdOp9URqyyGaxBeT7dU4
d20HUa6HoqiwYb/FOYQrPBkmhSIHzXqV54xCAe5sxLoch3RYFbOuOMdG1LzFobdjPE4fV49IUqKb
KY6FdgPJi+4HhLIv4jX91dr5rTArfZc2SrmRbzQt5e3S9sPc01YzlKhCB+R00ZqL0+WQ3q52upT+
WfM95EAyoLFj3OON44PcG52sNRyT/KPOs1BFFcXj9usVCQdlumS7ZeocfwI/7f4LDdluFGEdo34c
w8fx8mgkPNeaqq1tCYVwkwa89Wa5J9LE5xD+w43CZ8iIW55amQYCW8SXRZQyi9B4VBHNKKcD5Tyl
lrVTcfCBMtxJ4aigN0KqQTjX+uKGjSUr/n8sdq3KdRsAIn0JW6SwSx3oApi1i3jnzncrqI/AdVPO
X9uM8MeqLc1sG74WmdZgIeDCdOcBqk/10PDrTgUPEie/it2fb/drR0IiwPapOCJVjcO0mBkYcS+R
ReIr7bopKkFzLCFLUAV20V7tYTw8CB71ixCjhTIXN2t3uK2o0ivLOIhchr820Nxj/tInRiaCZJIB
U938aHsPpPXrNxLAaWIwvIYgDRyimSYGc1S6cldodFEFNtR1cNN9J5Ks9TGtA8sdQgiiEcwGewUR
JNODIhNk6cXXwEOVyM+RMJZkpM2+fVKH5Aa0FWpKUtM8SHoD9U/nPpKSg2JV0ygpsCqXjuwz3Qf2
CIg8jQ+k6vFPdoxtmppr1BdDFp38sB5xrFjn83mVMIyCuXgkvAh4IGYIm8izaU7Kj8sD03bXL2uI
xhkYNAOQ6fndFn67J782mcrN3XgX9eUMwvWpqt89QLaDF3KOyBIsjwI80pzbITVQF8gsmQm7B9tq
yQKULDuKxvC5QpjkXzT8pqcRbCMmCwxDyDNXklyihjR9AS07Ajy+rCpovr6jRQPspK/FqZhnp57D
oGqY0ap9OkzZmzT38oonEuwSXfy9oRoQTC7VF5SO5ab5vLI8UbnCjeli711pAIxXNzRy9s4eY6IV
0x86/r3CfEyXIHVDQxaeVDakKuA1tL9N3h268CVc2VfIjK/Du6vseVveyrl34+EhUhonNx1qe55E
3woYqjQozGgLr1at/epG4qwkgP4gAfgSFpo0UIAoc7kLdIPCdNvjEYPzwYFNuCLtRx7PKgyF2gSo
eTxiTDOQSXUs11FUplBHkF9a1yeeU5xtgTdqfpNEoGb7VniibfsO6+HIL4zAEuD5ft9O4mZEauM1
Hy6xYFi7Raurzul45Rm3JXVykJr16wyh2PZMPSWT692+s/KdCnuoETlIpL2FHUzsdzUH3WF6xbIO
TJNiqhyFHcwOsnjpBWa8Aa5f4fJJ8j4CaNw3mWVvKVfEITHoolxK3j4rooM6YsaYXlFbqAS6xKKn
rDSJGletYFRDoM5WQ4S28hOpW6LbKxo7MopOBeJOXechpQw2bfUml7eSTVZ8qYjkMAW9gy+Ykhws
vT3X4t24B8Ev7mDZDblFIDc4d8mmjt19FWaX6mNMauCoCTSDXnD3/xerHSLwQxh5uIOOS4liLzJB
S9vqE2Q+P8kqkS4se+2pzfYFggQkYoeUIKauKs2WXo9K4tXjA/6SL6Im/wew3p21tOonbmCxiZhZ
cuH8o2a7e328TSOcZFjq46q8U9dOssVMuzTlxYkuO5vIqdQKKYRDtc7TztLm2qX14qg7m+DnglsS
rG9xXe5HCqfAbRSTjNQGRGtTtqNJ1LSB9FdTNnqMemT7dk3z0N02Q1BvdaDe4kG0vsaVsB5oIfEi
9ocMZpPxE3maH44KrOcmx8+vQPLtLLH6pzyZJALQCUTKTQBU+t+RUvx8DrkqUgEe9UAv5mfXYIiz
5yZQ+n6lMOJBUGSbvmD82HDfQLWkvPGSveLHuBA8zk8m4MSjvi2PIJItP51O/O2S3aTloZaCePGp
tG+CrNgJWEJQL39wMTShCi7kT7EauMpNv8FLu+NkZnaI63wMwGzC3JtTQz4T5HbNfnC48N+jhCN6
NjV2QM/x4PU3jDcS488FhF6pZqy8s88jIRSh6+6wCUH9dhVuB/XIByTVLnqrjhSIsKP0VmEKA5iZ
V0MjrBrXHkl6XQPH7kAerWuOQrNDoQyULfjGUHiFRluoSu8Y4AmGK/yWId/YTvewileXt/ynsM8a
Dsod5ft+0sPh/5dFXtZcerG3xqvdEl+6Fz0pBjEIiDnXDy9sLQGt5HJXJrRh6HokRjE6gkcgsHPD
tPBkjz98RXYlmZO4Q/ru4tnjlnEuaHIU5c5KSFmOLoVXiVdmFN314VZInwVwkN9V2eVCOFinc7FA
xc+197YTdxv64uMScaLX57gNMLobEDy4fi6495C3zaE3J/9ulY3D42awZEiA/Xe3b+8dD2EUK68+
h4AM6YRoctaqsoPetUmiU1ueP398ACSw8jP90ykRl07GO9A1qUUp73syiDevl3d3S5wc5LffkJcT
her3S19nb/mB09l2ZMPvXeq/xdmjUbR2qK9o1sPe+rYXxwIQs/HJowkr9FkyI07rpgJZAwnoGTdz
tBdLHSWQSXdhM3vReGi24CKHDKgSb6tA/YId52VOB4nJZvNTTwX4GZe9MEHRea0iOvFj05WXD4Bl
i27ocD6qL4+uuB1Z2wnHJmXGXidYeF4DsFwIBMeFw5O0FDWGAzhSxHWELfsvuJZKkEdzYmq81OYc
5hlpaQy2BCpAmrZ7T+2Cth6wtnqX6A3i4x91rF0LZlAGH5kxWdel+101WmWYOLh4hnrq0a8eklfW
fPp3F1ZMSKyHHE/fVG77YhdAzgKF1PcYIQGeiMfJWwGsq6TnATVlCBhy0s9iJL3ITokaXGfi9iXT
x+j2XRB5BVT0R7NaEjZyCjIo2tpACYx8X7BSBAsInuTrJtmESfIaY7ougqgMrD9TxLzZZkWpkTeT
vZtokaV+dOnDxH2fncMm4KISB09y+0vEie6K9Q+mbP6A+mLUbsEWrmjX2LSIO3m8kZ4mdwOXWkgJ
qjE3w9IEKlydY6PnQl3N89KPuccjZADEzYcWb+r2+gcg1DFZ/s4HhKx3CuQXBilcvCkBiMTTgv3c
1F0OuwJvpUUunUKcesbg6mb1x9WwnsqvbNTubOEhNKXwVVwUJh5qtQ/lLCfKzPYu/dY2rKnkZjP3
zLs5WpXjU4z287PwzWg3W2nTSaVCBNC64NLkwnd5o8cxT84tXKn6Vuwjr7pKbScBDBR1Nmt3pZC7
92q7mWhO8XEloFrF3IQvekc2/b+UCrnVSTXMCmMPr/9glrXYT8lEwteNBXzqeMnX5VW5ro+jIbQ2
TKBR3qxAwyeOnAWCWInhbobB0PX6Qfd6Wo8tUoqzdzIaYGlel+w+DU2C/XtQHCQHfdAoX+Wg4XcM
uLHjXZGrOMA2f9YndhQD6at3kL70ZQ8L+TGuZIxoMhz8j9gb1dzDh7bO6ylVFbangHsiPOjTL5SM
QrWMdbvzwqPGGAQKf2nS55eqx1+NW+r588y83oEFcwq4B2OcpoZOfb1g7iAHI3SCVs2Vd79cIetX
ZIQr7x5UMcaBj506UdqRnX7yEK7PDRxG5lNMs8HkcV4VQBEQPKb9VhtOPqGgjG87LPUoRpweFmIn
/F1WZpETV8DrV+yq9S+TmSY8HVXJUg7LvOpOAabIMwCagyOrVwEGvLONuSwvrH8holbT/5mjivbm
0a76e7DhyYtShnrdJe8wbbmXnFA2/lF+jXYDqg3unQUSQN2+LEo6P3ZZgxflQ4BzGKoozL6UkD6H
u3eMgPTZPQyvVEDibdEqBYbb5TfY1B8cHODX+Ov/SHwcO9rlNdy0f2JI0qcr+XgByVYINNvjVMMx
fW/FuIBLf857/vMfvZjlr03vPz3ACHvE0lW0KZViMUfERraIKs3hjOPX/U865DxEo64W2ybFuwsj
qZn4gJW55bbNBGG/hY8WhgD/g6XPUdULBzEHEUBs19Q5tb8zo4E5JN38Z5pWuTue+MsefDIN2yXo
NVWlQmPh3kGU2aMPg9lXwDkKrMrx41zflqL4XAf+NxJC4HUUpdVXr+UTLyXDs8DBkwM0sEbsC0dv
hwsdrlBBJSU12zOyi9+s5+Ma7zBVuBUuLoA3WMcU0xZvGFh4S31X8TTU3ZT3hXQrcyEcfkox5xT6
IUh0UmH6xNBIhGECKIekStkTDUVlCblybzdmXgwA+tjCvODsywkssigZB8y2A/TrKrAjL9R6oNks
uqC8V9ItUpoG+ofnTLgPPZ5LqUXlAwCCTV7DzAkee4ltY9y2wIP086cIZnemyGVTcvenx7LlLq0R
oFX/78IMely6dXjgW7rjMVeruzLpF/qbv81ReneTArE9Cl99GsRNULuvsxLdQ82S81Ip/e+HpLI/
8AWVmYxNynifYIVUQjS/EwZwk8f9VIBtLIvLB2oy8jMuKO3RdgqruOg87iM3b2wc4FZjj0yEXAId
K44pfmJgvH9JDQzsEjf7KPrhSPHZ8j5D4lcsZqfI43j2O/cZNNb6Wh2E5B473KJ/0IWVivLgg5Dy
7Qr4HYZkOooXfIM9tCIQqXgFAGpHJJTywLCSEmes7PDhDF93bFCgkgVx5NH8ysruMgFETxi+LB9z
OFkThola/ISBS1ZFxhWjmMywBxsFQt+F0SltrEms1QrFnw6WvxA8FGkZBSXB1A3XxUFRv9jaxqUe
NMfet5535lwOEGa1qM9jjeAWV9jmTgrmrVSiEjcbIL/VqN0CE6kB/5fN0M9O3guBH/M1O9Wkubvs
AeR3yP3GmT2UO5dHdo/VNhOvxVp2vat2dT0A/Iwe1cFPrQpU3koehIQc0LzErLzz47XaryhyoaAx
rkBVR1Wus6mig3JE+1TiVJzYp+urpEy1ep99HIIUA1ZglvDk/1MEGQHTRp/GwkVq3l8JGVoVb5bM
09hF2I1noYZc10PD8biyV6d1haGJtbnugIgFK9Bkihj1IkCWRtoIxwUjEXB1w+Ei52pDq6oP8nk3
Unw4q4Sy08y01JJAbORxfJHE+qJwQctxs/fqUkD/eBxSuJXEt3W0vf4aX8PN5g6La7orfJzlcS6F
c+/u0zyjVotKD3W5byehgu83sYDWAw8lONEx7GeRnajEUgF4U4JIwy95dlcdIpQz7bnbNRgCSxGY
0VgiLzHCJjjmsTAJiCWAOddPMGTFO1IAxA+389wQTkQwMqvthpHnRGv8ytIXJ1zF8YFIWjkaragu
zkoRYF9oxHgGZ4u1rnHgV/jz2hh/uLfSWnV+s89ETtJm+czJ3zDGU4eaA+P/TUuybeSBdD+UDv2N
PMj5atLNQXVWFm98ijwCEyYijnNVwVWJPsCUprwoZ7lxXVz8O565Noz1dn39wi4vNIsHmQ++wnJk
fXV/I4tpDPS8Bo4zJvjUbPUPns09lkACjQcJ6jpdY9Bwf/P34jUlkbsLGf+rpUxtjK5wcIabqDDq
DU3JCaAWlVK5KtiQTNXo8xc3Hg8U0DSOE5Ko8Ui10u+M+8h3GzSkPQxyP7JRxt68738kfjgs5OhD
LghzYvG2kkQbXXJyPv4mwO2i5nrN8q0iXnYnBAvUhhPHHn+Wpq/PIjJmwHvKCcccFusbj5IuRgJx
6T4CZ7P3ULyNxbXaCC/zr5WCOaTuUAeBWCAMkYHAg8YTirMXoFFL8j7p/uba4Kez7ksbpElQG+fP
rHAwjgnBFc01UsfF40rDJ7ZaBObbrDDMCsihE629G4mrELlrEoyuTPzTAiCAWO+YkxrQRy+lN23N
ohZGlINjzTZLVG7+tMuVBzfQ822ETBHL5ocMH6FpTWawTQeJ2PMR9STPydNWfVfts7jOqTJJ9Bch
NuXrjJ7bLcGU/CVPyp+MT3RodlqPPvoboChcHsMIqDMAvvILivJ9C/a2h+YPjeUdTqezsfwu/hbP
DEGW8bFK1Ql/1o7zHTdA6m0WrFmYwJm1qmarw8aWX/n5EKtYzEsa+tPP58mTGG27iO53p+UqQFil
qaq877H9TbU+mK2eKYkaXeGq7Wy8qyKfNlhFVn6jmndtHS9k5SMkuQTuvzBnAvF9l8F9CrOyJ3gq
MQea749UPkLsc1HbCsXHaF3mYfxY/YyKPXV8idc75cJThjhFkSayoQAqDWCfEF8of7a2sc4TQ3xm
6Lbkw8IJ+9egBbdHkuXrqeI9VlIQ4yiuKcReBWRWLi1kSUfV/VtQpOqJoM3CThlThHuHiE6O7hq5
i//QXRjSxu+e4aWT0FJPEelzT7ctkhyPERXGct857oShtbdQ0X7Dioqopa2tO4Xfv+OGurjSMyqO
6AL83/1FbNLwP8cZNKZ0fksmlAy5fhXO7V5/jmoygshoS2OZy/uAEKiQ3NRjuxhWNI8t5Aiqw2N+
pBP7+3JWjNvbXNyBC8oEMnS5Og83+kz08s3IhOTvKQRnug7MVBlmKoKjDq0SY739M8Wbp4HpRG+U
O2jWR/2S8+R4wvI4DoBEm8XuA3KJrigq2paAbVYWiUhlTgqdCFUeS0C2Dyc5dxnDe8H6fe8G+Ybn
zCbhpk75tVUFgqi+hBhFZwi4Y+foKPvFw0J+gV2JSTr+gkIFfiylyAvBklsh5J8TYgqBC6UHiLnF
H7OqUwXSnk9d3dpEwFZEtKQnZCjBuvJ6AbF4LFznK+RB5LqoaeCr4C+JB/IIPAfMb6G3BUk6R5ZG
7hZx94PTw15EQmNmOxsDrXYliOH6HCWzj2/v3Ns153YgSJB/4By4RhOSogxmQoqbRLx9fk/XQ2Qj
GWNDr7X3PGI58erqzpZ4EbD2qYpr2yYHnLkdCHtIdRoscsqcvXQgDOLyw9lF96w7MOKEO56S9ZmZ
GVNPaEpMN7LnmSZroD9AboxCFDMjSDTBYvWI0cDv4qYYHJy5HwUBKQUx1FFAKym3xozLGrD6erZf
LPlJJPPojoM/4CCDBi+9QzHpCN5Y5eFICJL4ZmmsUb+zmtF8D68hg+l0LY737aDCxirb6ZM9rhbz
TAlorQ+kO6unazfTfYipVLRZuo7fbvIu6STNptFBMQmqzYUn+po6sRW71AfdU4vcr9YaiH/6+zP9
uJG4SzVoMjihEnzubwuHTHiBBV24SUSUOCZRvwSWTUlukz8tKGJ8UEpFC8vHUaUBpuXKK+XSTnl2
MF4nT11VG/klhXSjte+oimWteiRVtrwucYp7mdutGw7o2SAfi5Uj68H8VE1p9WvXX6kSJUThRxL+
6iwTBCXxFHUrpBPVGzEROK/8m/fzKc2z9AGZkXUiEXOpZBq1k04XfVz/uMB1wC7Qmw3RFKU85+zk
qIH645Nlxxpjlnu3HLO+IGc9J1iFNk0Awu5VPaPAmkriJ0X3CYseeLiyEkwTnKD2oGW0JS+w9N7d
744VhbI+ZmAYMnLRxQ1Syy7rbpCxfNVMTVrTfAB5fCt2uDlOKGF3ifd3+KydN2UJCh9mWLivh3Hf
Whpc7xOPp/qCAbW5Jh4Ufqyjk4XpYHHXUnnhj+i3d8l0fvD4amniPy+1q2VFLrKdv8jLf9TIZVZK
ufX9NsAe406WMEYmfF2xkOlK1HV28n0UceYaQqjwa/+2E0MowaUVShY7QOnhp1qKobKJAtPe4TLn
5HiCbf17WW+ABu0mPgmVMFJarNoCCEloXfWQNSe9pv8xpCjj/xN1eG021fHuJ6th15mTqaxZr4da
Avb1G/GiLmXN63qdSMqxubwHwREZ5b/vvG982KSWRZ5AsMWmEBhfB3RQH/u1OVHjbnMkkX0wvoc2
1xTG8NsZ+6ovFCs40UnqXEY2qHhGrD2Y8nUdOlFZomH1keiFBg6LcKekTMmHfUg1XLlOJF/+FhC/
0Oo9QLj2sAqF4reBYEe7Rm+GiJqDBZ9HVqffBEaG3rRP8pjZJUFWuUJWtfehDfTOrJ8zlH5qS/hu
8tV1ry3UV3uUpx4hcWkJ7U008uHW29CldAgLbr1rKHD56Bu/ewLleGk+IcJJ5zKEDERW4t65pOdX
eYWitPlG/1WB3NYrRWOztkgQ3LZW4GPs6dv8qpG2LvTdc0mItsxkNKnCVyNFx5Cv6uT8Qlx4cLR1
DIOh/MXT+777BeSotG1vnQOOvgm4GRigjpg+6dw3s0VAGhucP+0SaY9EgC5b1F3DLTreWk9uEq+2
rc5kq8HCX0//ksjMqPFc6mJadAoKRNpIVr+r+d3FWfajERhfzRBPcMml8/P284dF7WKBLxPkTQFr
tpkMN+1mkchUL1fd7jFrD6fOLoUb2/GHVXwrnK6QEG2ghWgZ7MVI66qaJfg353C+j8Uakvj1YvdE
OkZflglI953QhmK4gas4xj68g9r4WCuUJNeAt8aj2t0BSrjK4y+NCVoPzuD73HgMw+wYLiydrEOn
66qhQ6r9g7mn/C6fPhsz3DO/HrTc8Gx1610auVZL/3xwf+ymMAWXsj693edOBpU/IiXh1c5WprBi
ncl6vwov9dLmPGC0EOzFzZtdX7ECkPBCXU3IH5NE2kzy5DHJcDEtxZkCfAaFJTYPnfgG72zdNhEu
tQv+8bsAYjdRcj5Oh26RZkMhC4Pj62UmFHZj3zsWYoVFGd8O6EPDtmJM38pVZqZz5nlZf6zp6q2o
bmIkkYZvn5O9KWO30XMGNyDX4YcDYf3zL+W1MGS8J2S/7bqaB1KIHgQb7NMZRUZ/0tdjUkjRze9j
xYocoxjwtI+zYyyM2pkoVLF1Sji098XhtJujwvNd+k4g69sfq6lk8UhTxP4riySDkcqfSWTO1jFM
zxI1flxE7lzQLO9yybKu1YNxD4ByIbqrPccrvtm84/K6zP+zyJ30/Y1hzqK8L0wHzl2NePUe4h/7
hedM4xU+ovrqT542ZMcOq4MzYNTq+YC9WcFL2yItVViIMS7BHEOXfMxpEupZG9pB6qs4H7Is9jmt
PAQXTCdB/V79FoHQcbEF1fX1Cyv7oFLUr0Ha6GzP8edkaJHcCpsS4RsIMUxAUa8lEpnNY4UEQ8vR
hig/Z5XG2YnJWqtouh2pwSVd3oL6hsE3UQHHDdXHvMUjoyC+gPafKGU/Vdf3k+5UVGfmDP7/OxBF
recCD0ThVVG/9AiWSTS7QCEi/RCSRSJQ3I4u8yLhSIywi9+2nlvAgKmocQhmAJwF539MktnMrKRO
FVY9afACZkKqPAgHMq34WfpBCvzG8zjRIMlOBmO/ArzJsdIHZAQkQ9Je4d/2NIfjqaEVz6yeTv1C
ImlhFQtAsuj/d4M5HHWs2he/ROCVcWbhd6qqaWljGti+T3P81Wf8IVge07g42TvY0JaKj94EVL+U
TWAT/5pexEdJsUHR387kiGkjSnZ7lp3MMOrmvWaOmY+oL1OZkXlOYi68W0xelWDRBJhvqhhLWnsW
2PQUioSUgchSMX/+eDYjCd9FJJbNGsj4KujZCmAN6rddvAoTWqLrOGUYOLTHQ9iJ6mKZPpNrWKwx
xSZgT2B6YhWsaTnYpAdla30y/NkMEyQmgZYYt7jZYvV6NyU65ppT1xnTbIq4SIEqYc/T3x7fzf7v
sA1jgTUP1+ECg9cqC07F1jhUtvxZfSFAzfvPk4FNzdP/F0P+PWSJm8i4l3tP3X+FOAWYPQc5zuvb
K3SXcUkdN79XPs1Bd3LrJN7MgOeCf9sDaEsztg8iiOXceAgG0Ym7JSqf11wOqzr4iFZ1d1Ms3ZJ1
BsC7oDtnNI3i+2FeBmW803j71Dk8fzrbhg8wZfqjlH4uJ9X62t1OWpOVIKdd9NNpbVs8KBkWtb28
bae5dGF8pMgo6EtQtrciZLsq1TTOWHpzjkqnTpUCzg6deIJL9TW2E2fbkqJcNO39EYvlymOkXnI8
Pooa040uyDc5jNezBZN+cytUmwXDz0X+yKUZ9VE+JC4vos4UjGTE+hnuIO2JFk3Yaaltp1WzL2DF
lE/9PGYNUVMr7jfqXjO04n9knjSf+UJL/W+NOl0je7IXXXTUt8qSAIHwvEQGX+dbbr60/n8nW2Rr
/XiGrySG9Z9Ymk2QklLceNGrjwhHV4KDWmv8d0f0TgWjljk4OqH/ZNena6djjdUo13iDMwO4qJ9N
fYo15bU4UFj1rljVfEkjuhqBPN7GSsipTxXL55WsvsufHZvcQ73LNsyaAy46JqLkejtWN9SXPQco
et8aae7W97lLEk0W+FZXTTc66IfC5a3eqDnbaLqtUJUL4qL56A4nkIoFrlMgzwwuyhumOGbvbOhx
FJRuyuWPMMadqUrsiqETW6KGdHSSPDe0I0wlRjvbw3RUWHBWYM0zF2eTlDZRagpuXf1RnEo6AUGD
MeBh/duqy6ZN+w3qLSOIfe72rsm7vdDL28UXvf/eaX1tSa20428yNuNMjZEw6QMFGLInaKmTEgNO
qdXETqmnBnD1ZJarIaYFME+15qhLsFbqpdIP/s9Ad9zJCMiS4unwadRsD/nBdDp5OBkmvoo4Q/N5
AOB6pQA9624yYSUg+0UkviVp4PhFlR8f059iTKJR5irjNmZPJ8X9jjJ+fw84jEbEpwhV/SQ4gM3+
lVpS7O57i+3jO3PSpF3wN5Jd0+FDTzUoBLFCG1o48l96EKGMRuc2FIOJbkkhMdEma3ppgIH8hNp5
DxiS6gJihUvFzdlAU6j5tk0FqUaa6M0sxmecuvcJom/wHaA8PXm3F8bvPgy8lLtmt92lmYXMs9bM
NRf4QTO+kMVT+NOdQrJGksA7wriAGoaxNu9+IDLhNgaIdyhvKNw2VAWS0PDJn4CLn238ep2lDsqk
IbD5qhGO7AaFzawKfeLYT+mc9Wvl7xuoqMgi5/nLYx7T3I4o51SROykeU1vFOt0myDghK8F114tQ
jshzOBy7RoKCDAPEgq3fP4kwy9vtc0r4X8KJ2lK+xzTaAWcK6Gjw7bU5ffNLobbF6B/QXn2kCjiP
msnEYXvSclbPXo3uA8HFDfnr1RI78J+n0sGMPmHBL/3S8fT4MvKQVvMhGQgeT1UkkuLW185IQmVm
6WFH+bHnwfnREiG7xF3roSQiLtuSAKnscLlKbUIlKFZoPO6KNH5CKWrYWf3VyEBTTfWMNUhLn3N9
ZnS01u08GF3uVSErjvwo0xRbq0fUKFyuU9XlQW+lkCeUzFxcYTBhr/5KecfcnQsyoTZE2vt3954z
Vv19eKsAof9zvQ4u9KX6X7idW1kJtgOakjBVbCmEuptJHc+ZI7iQ7HoqEkkO7LuXyHO8/o3zdOsh
+xJNS3PlJLibCh1Mo6meXAeK0Af5v/RlZ+7TocrS2gvuQ9JzhwJTkN/pcJMDcf91+b+I81WFKvG4
P8nUz2ROm+WTA90qSNnT1/qhF7SWnicA4HyAjouMHiMHta4oen62n7WYZ/elR/O6U4RS6Ik1ZwJR
FM6miYxpDFnf6ZE8cc8BOTtBLubIPmWyzGhyyZ19MS4saD4DjAZWUCdI397Ln3hfry1r5ruOxn0Q
vDPPkPwH2adCzQVTYc4snhlnAjOn3zE0Sgk17j2PyYwA61MzAERgT7+ZwkQOvLdtY22MmOsFRIoz
YheFr/jCcQ3Y3wgq1rMsXU9Ro+LdHJTPsqM2fzaEMjPueFlEI6Gz7WbXeL8TSPVAnsTWbaX1dt3e
G8aJ3BRA8keanr1DmwOAegEO2Oh2m9W4QuddeEcG8+9uXWfI71PL3/u1KQsROJ0t7bFJkJcCsQsX
HhO7pCEiQxGLG4m1wytcJuLcgPHzaW78xofWAZlfZoSNc6lMbHtE9fu6QOgM/JOvZPfQI3gUIBJq
0zcraTHN1/pvAh/uTSaQUvV4VDqCMauNmkD2Oy9OdiURMuTo4WXc0hS1W9V9lapzscdgJs844uSJ
Wq1zaVGUMmHETnqa21ntCGIvSuJh40bnYF7IIbLue6mtGzQk+Kfz6QPVyssYDUqL4xyULFNFHD+6
o0bpt4O4KZWNbGgzYYs2som/2c4iKbeDJ7Kn6//ze2DLF/6oByl2ZRS+1/T4YxgcpmmDDC3trwNQ
k38sGwy3utZCKUOGkZWM/7USTonZvyDJlIPyjrtefaQW/WdYIHz9xsLTpe+e8Ly27lcoZB0ybrUI
lAhwdsbBo1d+uvoFCueaQ9q43P1rBJNARnWEyhA8Jx2PmCazf3+aJIBzO5/GKZcvu6po7vnyNFWG
PWxE3qj18606TsikcCnjIh8d8ERFwZxV45ALHCQ0qwr/J8/kMdzv/AsLAzQeT1QEo17Bw/n/FqL6
t88yBTmeDNDMSRk+BbORSyWTu0nLMv+x5VTJCqf5VGG1am/3kxF34j6ndC25Ei3REXbPoT8TBPzv
uoJyrLLpEWvtfhS9hFej7RyTFbFWKonvoUgwlWjSMxEQ7D6W3oUUD3qryi6ojzGuWLKb1sitiTcJ
fXrsei8q/I+CEV8srVbwbXpif3opsEvKt8fw5U+mVitTA+1951/kR9N5Dzkh4fNs90xpzz3L88bR
IKlSYwwrq1q7DXyeDrElX4qEltw4UC3xuF/vzUPcB2I90qQfcfpCW7hbqPAfGDbSTdB2K8duew6C
YSSaEVdWWkS9YpX/N3ObeDocoiWakp1boOlsVineoIW6UtQZDIVoanSsPzeXMHIPuFHHnUglSS/b
S6V/xs599pYL5jPCrUENYRiPS2guzIa+wBTJDgRFycvys5O85DuZ9PEE1ANKbl+thSpKqW0QPZlG
lsboCSNbrawYlZv2CXhUluotBVj/pFobODTD1oLECNDGB8hJR4CYMDUK9WGdlRpZcuETmApaHNc0
rVTg7Lm6XdCRTxUDuhlzUp5lbO4BC4krv77Z6+BgWyFb3kh+4DBnfK+jKpUy5CzTjPCShEBcP6bu
a1zvpN5IGvsWcylIT8WvWKGHhdO9qrLKlyK5bOy33fqiVJZBMfx7X7UYSHb3Pn9gc/yOpZa2je7+
j086OYnLokMK28pgJpT0D8S8dH7fqMgW+ceI2nzYtxypi2vsDnV3wQhW3y89yKNM1Rq+sMtvlbfk
Rk5HijGxP3J1OWtFzQSLfGuYyy4z7pmj4PXrLWm5UHiGXBPgaNegmaGxQr5NA+QPNerQCCc2M7+H
GPgCBL9JIsUxQB9tS910S1u5nQOszv5SwVajTu7p/UU+d4vdYs9EFRAybI3rG69RWVNZIZGUeSm5
kyv2qHtUZ4RAUTjW8qw6tgCSSBmfZ3IHjcJwz7YwzEM8G6UKwYrUsUTsK9L960t3m7fcHf+e+YAq
DEvtRRhLgWQjHvRkSB7W5D4C9GVnXo4jVNWg7Iae02OhYiTUJ4XlIzL9Svr6ZKQ+lIYzDE1Yegfy
xLpREtKkP2Sb4AKgAEcUL0NPMOoFyM6Tlwh5xqLRAFrMNCdo9ig1YP1BdlwYt4/V6Z68IwETyoU3
tODzK3pIjYtdqpkZwmfndiRqcbGqaqbuvnhcvosjjrKArf2csYCMf4QdrlDx2lJG6h/63iFgH6V9
p7c/YCJeRuD975hSGxzzXrxWoZkgiLn6Zs7bULhZtwmnKSTbwyoI11t5RKz8OFUTORMbCI5z+10o
Zf+ASGoOvctlsmS4Ck/+6DxhdGDM2DH22p/2J6dJ+ADL0HkZ8r0fsdlOvRUn9t3AqKOeR2Tk35e7
6/b9EqewDXGItsM5v0D2FvjfPWqnyigM455oG3mQUlDyIAMMnWNI7ihgmWhKHlF4ZPFj+piZX186
tuXJ1aSZoQ+mca4WIRsjzl0d5bz0f+qaU6mXQX+hPj1YZNzrIHsWl1U8feqXddDVHxzRG1VpEVRW
+lmgnfnOqCKxNdGivvZOo9EjG6DkdyQZV3jUNuFB8TzGuXFQQTqENjRdcmmOpO7bsbA4BErIZWpQ
cJTWBiQ25n7StP+1UG1Q5YPiBXZ61xrIac00vmLs2nggThevebB0ngCOECbggtjP/XUbtBQlANHt
uBjjNn1ob2oKb0zpPmaCkdDIo6rFis4thv2X/79TxhO744VqIl3ptBeqUbUCh3qYLnNc3JNBqZpc
qDgeiBoViYhKet3YDfo3i/zZXjuPgg5lh5t/Cj9xc+071tVdbO6fQXd2V7x72mwpmobGZrXMGNWx
cOWqRY/yf5ub82SVFtvx0zDzY6Rpe8C7IWJ2u6OhgWVMO9OV2ZqqthTN7MHuugnw+2/d3cckPzdy
WebIrE+G/Gf/kxcI18dK0DGsS8suhxG+rAJ3Wq23W50srCybQbANKAhal1u8qPfAVkPiyUSb8ooM
3jU7SaJlyUPVmFMQj6VJQfNwsgSaiJZTkjid5+ilek+8qVU6ha/Uf9NNGL70Iq+GyQfOiXAgqaJA
VYFxoQt07SVp+7GzLLboEIAAElNZaJVMFY0/j2nNThY64RtivaobUUtoXB+LLZttitpVkZKmDr3U
zJQwn8KyM7qkUcQt+QAw0gqIgb8Uc/re5ciW8GuzIs+IWwyAoMEsDRIaAxm++HpZwdw/WUN9MCxq
6244LTOU9ornwzggRWnNfT5KHuYG+/gDHL6ISbi3aS9XLfjU3uIwCMwA2EHWRfhZIzhJ1WLsLv/s
o7tH1QcxjfzFWsmBzTau9EV2V3OZehlkgVq7NHEtxIQ/HbPRror1N+2dJqL5i6VQoTYBcSQF7JDQ
EkR1P49BptwU3Tynajxht9g/LBWbu9AvpDbO1KGxEUfdAr7CL6Hbmlnucz+APJh01BaO4HD/rqCV
dTCjAvZvlyj4QuOIy2j8gB3GdPcu9QuJoavyuADsf+qUrzJRuSbfO7Dr0qgf0cuurrk8efnI9+Pm
45pABDsCMmOvyWwcTTMXZaZ/oszFByBMwQdbo0V3gWY35wD7alzdLBCUCy+B3uU2NS4q5xWkPSwo
d8++PjC58lJoGIVz5mIbQxmAkKMA5QpB+eXkKchykhfLYQJJuVI/Xkku6IiqVORMJ7mXcDMadbgc
+69kTB+lEJy3Nl9khaXR8S1GX0JuoCE5isYxa6p9xPoFXlkCq0hWqhL3FRcEqa0oEeA/SQyZwQdn
NguA7kkp6tS0nSccobG84Tdfi38bTGDvdS91rDzV1qrQhz8N1jpJ4hFbuozX+RcMtkNRFL7bFhrF
Zmw1AEWxR9BuXFmchp6yy7P52RU/lMXtLKltkC6wkNtM+24euRtwPjEuZ/5IyRRxI/ewk3I3iOZu
Q7R9W6VAqVTLIY8yElko9z8GJtpU6UvVC4LNlbzDcO3yc8fbJY3O/OmQGOnMocWwQTGbqBOBlUJz
Gq0mMLySCj9vhULLk2MiDBEdfAcOPbsnIFV8EY54ZEWZbu1g1GwuXytSzyFEitKBmDbGpV/e3iJX
fyLVdPclzFPw/2gL2cKCq+MDow821WqJCN/kE9UYVnKOghwqMWd62q08UrCyiTg7XB3+nlVQZUmh
zxUBkZSIvVLm/j2chW23etixcUWn6o816TcDlSOn8EuPwVC89u80/nctL7o4B5sG23L7DgnUgY8g
0UJXvlFdpG2Ck27vFRNA0nJ2BwR1Q9Ts7b6uEo7nEFOFr5HbW5StznMOkGOlk5ZM05q7X8NJJzyE
JunJ4zULb2hotYK2oYWcGlzRyGo41yuRicHUK6KOkeyBi+HHFVsDLBZlBka5Ymfnl+NTPS06lTz2
U/5o5LlOtKAQoiFZsUztbuBRkUQ0MX8L+SJYOZuFCwkW9ORSbZgCCWrAF0tukKFcHnMf1dCWghc6
0pwVUmuupmkM+3acEOAMwfb+lvh4Td0y4sbDzfCjMyJkG83Zu4ex7D0gsVkAlMAkP8h2P3bQGjvZ
brxDtuNMRFDL+99fNbVsie6LkatHyYV9xNtilvGmyNamak1bUcu36kVXmI/3BlH0fMXvYqqDCPP+
qe3GeIBrR+LAH+ZsMz/+9FohdlTn43KT3nH/RGt50ib2hwpKiUVY3kswyGR3R4W2TqoxrDWKSvGL
eU7Ij6XtXw3LktRHoZnC7RqUSR4dbJTkJ+JPg7rK3bltx14HkOxIE02NFG5FFh3r9DtSlJWaRLPI
+K6vwoQfvh1NxpuZBsE8YgY2pXGnL1/zbxM+g1tmGmWjxdOnFWhBFqG/hDfctVubD54QcAzn7yy3
2wzQeiLUHHfC7mALDcRIUF/UcCfEwvdfL3APg3Lkt8XJ4wv61udxnaQVEfB1DOjaK7y58r6f+Ln0
aTLI1vpTSXCvLjane/uRr7kZ8He4oorm9zuz2Mw71tgyiWLU1QtqEEAQudtu0R7XjUpTFAb6KHqc
L9jUWM51KAoR5/ArRkEy6ngHybcXeh+R7fho3jOgxYVvAQdoyEGzUXp49rs9zUFAGBhGoJKlgyGZ
HrsRpkiZGRPdirE9tXU9h9NfkZXfJYJF9JjmTCAfLj7Igooy7tF6s9UEa5Nj2J0sCabtZdiwTrv9
XzPGnXjB+ccQ99wekIeWeqI6KinKkpjitu6660RWhwD4KVbvAJb4IX/5qB7kjTrp6PTOit/gGySF
hjsT2VMoLD4h3Kp4Oc41gv5sjaqd5u/Y06akTNisg9xDaxKEBXLqEQgLv9EAgJQxCFj+uJjvE502
IpVW4Gd6G0KMuHw4sp3+e4kQsjTQSVAAa4jEMjQO+V5xFicUpzIRWxwX5yqSYUsZxCVTWKlmVGbu
9isP149IV2TLj3m7m6WU/h5kT6UKtir5kstyKnmbkBn2Znp3uOeYE4swFpkoQMikhBV0ZkIrpN+M
FmJ+MU6gTQaHUFUkdf98sTZyAS5+KVZPhDi7TwuFwg9trXmJre+DS1KLAwbO0Pabo/5DnLCz5bF2
k2fJO9QLiKey9+2Q2qW+X1G7YM7M598XCn89cnDmZ+JbiMjok1nvLV0B5bTjchX0zXJnE8IKzzZD
WnctUtXSKQc1zMcF5GJ+dJq+AmGV901trU8m70W/GvSo09rj5hg9B+IqMv0nFpOuKAmMqJhJ9fa1
7E/jyzf1NrZDqjn1JYlGS9Ijg5HH06t9FwjN82+DV6UHwGvQe5Avr83oynXwNopW1sdFEJCfmsf9
bXfi+IDMC7vafp3LVEq8enxR2vMYEAkJLCGJFchu/orUvRj3P6vLouRSmtBPmyf/BeT39FRX5A10
f16pQzmNtqJU9EI7JY02tnBjrNytDhwdakPS0IrV1VHc8Mj2N3lxT0KwJ7moylejUSIUUYbLwfgU
OVz2yQFLUMgnzdQH30hHV/CAbr7ZMhJwo2DnerbFdGHz1QqXYP4Ex6oxK6neNrXqFBkF5uKp6yVo
FjJtA+simtIhyJL41nHUhqnZiWZK01qDnGKQ0fjzKxy8XQyweJgYfUiSxrvJRZMF18GP8rLd4Giz
xcCBt2NjVCc231uLdvplGADc26xNPWT3pfdbGLKH5SdT7Q+GFEiNjt3oSiObXGWbIk3sJKJswy/S
x9+7spEYuWaKzbaFP97/yBoG2NMc+hWX2aYCw4B6uVokp9cepuzabOWHcQKDu5CytxliLtH1ZNBz
BPny0nlyCqBINTXnNBM5SJll1fZgWpzbS1VE6NyyUi0zq2dLyi0RnwnU1Qze8pfTznItcoxR7hcc
MZKM8kGxQpRVMsDNN4D0OXTq5fEnoGN0HX86eoP03XmvjZmOwaoh2ir4AY5MM9eZ8HzGVmIgitAY
PghVUATep9pdZSxsgbPmSOp0domgfDDjQNuyZl27SEADZcVPRGq14VR1AqiQ1e9qJrY2QIwmRMHE
vprlZVOgliRBfWU0DSzbvZf1Nl8vf1DAbtz6D8Uy5jrz4UdE4DBnm+rUqmYsrJ9VkbjZQHxa5AKg
G7kXePS/Oh8aUH3j8oy/PYONuxfniuB+TNApMbbCXH9VgTpjrvBariudH822p5w4IBfF5kBiuC7d
8X9ubmleNEfsQRG7vtrlDN7qMw7ln945PWuix8pEiXJbhXzUHrYr3dUPnzWxIIJlvnfouK4a2h4C
q0OQiPjriI6KSNKed/owbrhNaLcP7Omu/5W/f1cL9oqPwHtIYPaeTBf09bWR7ncYKCOsq7slq5fD
fvWafQx5XDBWu9d/QeL7FOp/gfTGHB20OaOCqnum8QzSRsXgQJG2zAr96fIeGy0PdcTXbK0ggTQh
EHx35fWwTGDn06O5gyNCsa5aSYhUpAr63CShGTd2OXs4qgii1n5pmTNRCAThXU1DTX/hr+8H67Wh
LDagqxLtLOZTrPuV8rxsErc/thH/JAVKDzYTjNYlV+56vOHB2o51MKkOixa3EJWxO0xhQqfRV7vP
ahKWYIjLYDx74F+WrLfuUVveMnHfC/bhHNwkjPQdMC78pKUNQoxQjc8uQpc8Bg3rXL76hI6Ed6hy
Z7EoVX+GwQzxWe5UJpMYiFqK6PYLSFATTlnTeaVkqYh6KtVgqB9MxDo38JXLEKv6x6kQspfsgq1d
sA6D4U71M7ORI5v+/YEG1fz7ez9h8pF4GpxePmQVlhZp5ZDOgoDRf3XJZOoztvYyyXbGFMlcbKid
eWgCUbBv+jBbr5ee5fk4rPw3CAwnFsKoUWtO+HmfSLNwZVYV+Idsw5njdI+ayAW2oeBskcMYM50Y
e6xkHuuAvV4HqE40rTImUbLSCg/5SLKx8pPLcuBpW+EhbvfrB4GQQgh6FI3r9nFJ6obDpYxzuCmf
DYelLh7cR+Gy1S5Uci2hbTBzV6TmZmO5hCcoUQa3pizGQgayzP0uXbPpeVQRMxGutfQSLtQ/F9Vu
UHwkMOorW4oI9Lp5mgQ6J933vWvQsi1PzpIOMkrdKhvG6xLTc3Jhfmi8YgageOElM5muDpTeUXFV
1WPPzlnIINGvVmYQq8E7nZHh8dS7NHRy88yFRZ5FA+6E9k86764nTBDiU4lutYyEIiPrDZtbClKh
sV8h9Oy2ivJw9GTsCWbJFPC4zhFYSd5kvIsY+nIDqtR3e5MJDnDW1rHDV0fBUAT0SwV3SvYY62kR
f5TnnpescnVB+UjIYkMZF76o8hjQaXSxCBioet/g/N1p3ImIr+sNk7JHP0E8oZDhV8DDR9urYiwg
tshcQqeaerbtzl5Lvog1tW06r0vUpn1LLKVM2nZoSLA88rl/K9doLcU6Mhqrb2ybC/kqBcm+FvG5
24qUfOt6KDxqz+MAmaSvrJrk6d2yAbBHnnspDZ3osKJ5ac0xNMdh0rYtZ63Uu7+8u1Cvd66Iwuev
l6W/W2edawADXMHtlD4Vohx8RiB9QRRwXRF8VeUjBR/jt9AT9ZOELiDMfaDkSPh7KUnsDqlHg9wa
OYkqOll2TpryVBih/KkgjjF8sUrpYPrwSRF740TrhbcwCbEoCSSleo0ID0l1QNNtJhD3yMOScM8R
sfh25pcOqNDMHM1FJN+EKYUChM9ONxvBhoBZYrxINahvaup9AznOfOAZurvF/+SEr3FqnkiqqPkI
m8LyhAE/0s0QyzTZ6i5k34uc/oT5GTYigTF8VeZMnQIEZNY15unGPqa7ESEpPvt9Q8PkAjHXnoUg
NGhTRZNDS/Ceb6nAOjz3pi2TR5dOi8TZHX/9WLxPgZhZyGgPHSgATxZ8Bnl3VJWvccdEFMF4+w49
0uucn+0vnIJdi3Zci3PCvJoBbGX8aIPHfotp9mD3aYZFs7cSU/7wmDpSSFaRPj+6W+GQgKH0AqrQ
m4AwVG7GndvfH2D43JTxs4B4VckwWvwezCbq9TfH48CrymL6hGOYjuqWySN21hfy/R6CWQHtTQ9m
VkRIqTw/K5slTQ+efuuiEl1hVsJn+tbK5Je2jKnJFbUgqwutHokKj19MCLG2TFQsqf2OCRcdgWZP
6ZL5HyxsO7GazK0ucmzuf7NWi19a1GxsmhZshJj2xS0rr07XbRey8lDH0dxeryRL9j/RqRyN65Qi
YsWgOuJnD86v1MHgVQfvLIKdQwKBfnjDtjjsB5/shGN6cw8gaulL6KDIMKc11ms0oZCiQogHM3UW
9LM5aNAa+sR+HXWhTBL805LIIMuEccLzM1Bci4z/zbIhmsHeKpSU1e1EZ5KzdXDgpuDZf7Iq9pea
b2LJxM94qnaqI1jgicaOlciyl5QBxHY4Yl+JfXoCd0RWUmvTD/HudaURlHRLn1aOKxczqLRwrrtJ
bdqAWFUMibzV8BL3f5Qr6WOff9jd5DeAPPlpc7SxovuHPVc7kNOf1bIrR7IF4lPJyLrtycKKbEWm
mU/ppS0O9MFhxK8XopQjqggpHtIFcLF08nV3YRsK1fL6guREo6fUKotZcovP90kroWx7jhXHjOkQ
e7EPPrY2JHv9hCoYl4zu0cDCUrmh7u+ARCcnPzOW3mNqukM88OqopCxprsiMEBby7uoo1C2hErOw
NMs1xSbyDzPVjlXpC6YW7bvFLk+3pEhI5AQ0ya2xSgPyIdcOOMRYsKKx2pyVf5sO697H++EV6v4U
NESK/Rq45lci9/LkoVrElX7vfjSk0nB6SsAQrR7EeggpKG8D3GzgSZ0fej5j2RZpARuyabKyryum
Yu1Jyax4tbky51/DY/f80WLJO03GXf3ixs7w6XlxNNWIpAddDz3E56jq14nDPs/izmm2mFxoYn16
FRqYFyCLDVs5FjjfDJiVOC3TrNugjRZ1SpicG5aukwXXJhnU7rEJ8qykCJrqxjpoZGQLW8wHiVwG
Jt7wONQXDI2ZUnKfyje9rAyT3mRFSa2sAi2/uVQL97By8qAR4keiQS00hW5dPzDpEZmtwJeyp5nr
hay63meB7cTZz5ALtN83DF2Z6LMB5EOifNdoJz8sx+gCEiYyKvpuT1IIHe6rAfi2HnBgocLdg0XJ
EQj3ifFJNPDwOeyzrVmrhJwKoAl2hSBk1pA5XGcvi6gUtMFSA61fEDMhrI2/DzhiIlrxfYwPBzMB
+t7yiJm8razvP1z4Bd90eGFlaLWB1vT8QwmyO3iCRvkeVCecd8fgOF4KYoKzQcobmC+lPjT5w3t6
FN8ZFOPituTMRkAQP9Ynheu2teCcbH4hk8MCeruf75DbR/AoDbT2d1xqUKh0gQTSIpA7m/UJQjre
zRZFcpqyo7uK+yHJfIqqSS4h/WR5sWcNGKqwDFIRleJMNiHM4x8cw4dS6DW0CYrlLwRDv1F/7snI
Jgyh5/ARVSCIPwQIo8gwPGYEW/V1P30cUWk0s34b69u46cWIwTvLnhn2rjS4Lysgpn+qsOz+RwhS
l2bNzGM8j7wE+oXMV3Lk7YjdcvKvu/hBJIMiF7i2kKLTaiv64sk2YqPROi7ZNcU4Oo1EYaQ1y/HF
SENA3DjEcPiaOTlVApwNSkw6uVwvjkK+yST5u+HiQb4vy+p8hSG3WaaOZ9Wa1t2Fy9PLeO7ceRIo
T8YKvmnmdnQMcZ4wyt6KysS7TJx+Rej2GGYRvycIC8+iEdLiLQ3HfH31aeo6+1qImH3URk20sWIv
3BT27FuX7inHJR9RR9B6vqbRkJ+Lv3mdt9C1EFlIVlJWlDQYOn1jI995wAPdu/EWWrAmfigKkuSU
2MgRozQUFrdcs/Z/VC400PXtEQ4Vt5liv1s7dFgxlfUtCujqY5WU0GLL0SlIJesM3yhYmLATVqtO
82gQJ1/Ckr6SSnJ+NHGqxayYo9B4C50oZNJ2wZr1S0kreNFSxdycfrMfVytylsDu0kxSJqrgaxQn
gLXteSjAb+s9dSCKu9zqj3kG/1WiSSxipL1u/1vqjaWrLtc2X0fk1F1hybimCcgKB5X4TtNvHstp
e9Ma5KWECGYsOlP30sX9n+5K/q2FCPTBOhTFPGIk2XkFe7n7NcrlD+1U8mVcbZ3B0mC0FH//FGrb
FdpGVoldQWFbTRv0jUPZs9Yu0vub8m6QeQJTfWGCAiPlGGxC+u5O59zLXf2MspuGpodAYR8jJbqz
1hneIujY2SZhBgf1FYCfTJAqyhzWvroGD2L3USCn5N4ITt0cljJ7qanASIKxjHlz4Qbb/gTUkAn6
0d7snS306o8CsWU7Tfzqn2z5OpIvczhJ+CUov+4nyegpNJQvVmO+dhtRa5OwuXNu/fahAo6Fol/u
yE4LA3pUuNzJ8IveVBLGpnAZ5hMbX1vbxz+Kl6Gm2bLwL/Bw1Naz/nmD5bn/6f7Hs+6HaSiRJs60
BxLTNJd0CEqaw9tAFjigBVZXKoSa7m+KdlJAgST42sUdtK6DwTI4PwREdGQI84VnsXEIIzIQwR8/
/wp6zy4P/rj0N6QQmFT9tQXFjxIQq4K1IFGuSPuIRsLGrGBDCkeSfAWP+7tF1goBWzpGBEEa/IGI
uh+W5vLSbSSwoBLdPU63j2dWPNkGfxU0HSJ+jMJR1DStx8y3/oqfKulpFRJxOKqR8ac2ErGnC3n1
R+Bmeem2G1geW8+ZmX9U4L6EAux2JD5leXz7x9jh83KcV/wzIIZK9k/94ZXlVZP33qI1eCiMCbDG
RyEOELX1bdnzWAquHu7pjGqUJB8qo2xWuIJmuHNrkdeK2ip0r5RcM2mBjpBpk5OMKug3aa3h9lUr
SX+tjZzTyClzfGfF9lT3/0FXjuM9zgwg4Evy8QonEuNWodf0c4Ou6d5MmU+wZn4CORX4KrGlw4FP
fMwkPT7kN31xfxQN+doM+kcwC5Cax6cMHgEsOq7NgjXNHBR4klMUGMhjEVlTA8Vfq2D0Eg4+8F9e
FVp+etlBHRv8VZWHKM7UNs0VSSdBTo9w3RMyCTNx0IgDGWp7D7uvQFrJ5OhaAb/HvHQm75i8UqsR
VZuKMAB18so1KlnpUPff+ckbs9zGB8Bz79L57KfVmqdtm2DQ4M/FZP+N2+ngy5SZHe99tAxwALzl
QELY0d/qk+oHhjzFUaPqG/0GQRy8hGPyqjTgBuLpRICVBUVir97qJVJSgGrP37GXQl2FSwXRfhVm
8ePix5XDYDP/shKPlKI4YC6TWMUNytNmtTXucrK1fvggpbP6vSmhO95KuJwhjAOZ0KoSIJnG3n2G
pKXmrMhOU4IBdnkeHjO4Va8ekOuMmwBCiRiK1AhY0QbD+Mt9cQ88VVbOipEnZcTouKrPTf5xKdM7
T48S52T/0nAbYKj5aHe1U8C0vxEm2I2wRiaDEgdlmTcHbQzmP6YzZFvqyN7jrVlOM/Yd/OHrcHR2
L2jdgcqc+p5QA68FaXOLId99SSttW/VXPZucFc3nF3z4M1yybuPL9u/WzJcDQkZkVS0LD8ILIsHf
nU3mTSguNzFZPabf1EF2+Kkpu0zNuNVGvgyGOTz0rWCGCWugKh0hXP2M78BaM0BG5rdtXLJ4Do/f
CuYYg/A7LB3vem2sbmcCxwS8EXqLOK852ykaDmFueWxwqEzkeSURuHVJV28CJlP3JzXSyeI/Nx9M
XeRNRfQtPAJhgtw4ylwYgqBmMewgnj9sX9u39X+y90nZb8a1a+uOJ7LEXy7/PWvCE7uGxUanmyji
ntELCyVtDWymOw9rKZeYjUaQEUzG/ZfFr9LXXlAlMwD/IymSha8hL1cupNvVmxoKHj26EesbCfl1
mvoX4KOvTvzBl+smC4SYjrLMbhVq2RRaPOFsG2SBRNBeELxrSChlIpnp3xxoL8SIUENfInFuO23Q
6EUz2gk6odjLI2i3P4hqw4Jm7q+FzgkFLf7eGYRi/gY2tvgTOxEVIp016QDG2R20DfEnkpWSm9Jn
ZgkqyBJovMnF5VODUV/Vvgy/nnbddGqc6TAvugDVrYMm1L0e78k3QtLa/LnnBuDNXGLnz/VHJHP/
jfOjTxEbFJ+3ROGJMVaQ+ggdMMBOHtW9nrMRST2rRdi7Wz/2KXimQdUGzHFQTDXi7NH7JjBB5ZYW
Kf1OhWitTfHQk4c9RiCIkHp8RUcEkSboxnEcWVuUSwW5eXdUjDlUyF5f84RoNwQyDRCerBdPkIWs
m16Ul/DoUjJW97/D3bcwOX8RXnOW0XK3Hog3YKrRuO8IaOml8wSnQFnve0nfatpYEVrq8foJz/ql
zplhCuJwyuCO1m+W4EYgFdImYtPhFxGrew5eVbcnZ6jCDtd8F6CEehZIfZgMUmIDvlW1gvuUUGD8
9LFZTDlzHddjmoP55JMZiI43rrjgJpus+VuVWZz+PM9k9P/Utt4VicHvoK9mBKwOB2Va/06GLUEV
RlfHqmc/lrvFQgpfYXT4RrcZZwr7PHC68EFU657S6vmNDkIFIiiXoAt+bbq/a+JIiuzfv8CzQsj8
/s8JClpGndq9Y7tf+3O0JehYtKdyAnZoOzymSXFRDhotGufuOS2r30/uZceivMIRY+M1b12XwWIq
IAHf+sql45oVog4mxe7eANYNyXIHSr15FP58PtENNgxD5vRINBxlkbqcqgWCdXi4NJYisTzKnJbF
rDJhMnNtRoAj47O3C+K32aKH6RUptfxyLOXnKCgpKHHqM1ngaudcK4xVrtVZRcfmcZF62yM6oOHy
csu6Op3r0ONEfTVLLjlgOUNiDRBV2FbSIZ9V9mG11sTpJHMYTtTdpyxsDmThzklBmbiBuro4IeWr
0Y1OZXlGbYC9+VHZcNQQKOwICTAY9NteItcKJghdSEAQm90aQa+YmcsqlXyQTDLu+Drru2CbgfiW
ttCLr2rbdu+FziO1swRkKCybetAFVdC8dMFJLQEitJSNUxAF1xGf/mEikeRScChZUIImHYQZ5nLQ
VUeY81J8PDc08cv3KS3/Ke93fpFeUOJaXvTIZwB0Y0HOrt+pTMcKLFv75w2oC6tE/DunPLz/N8tf
mRh+9EIjFunTiNv7WdH6MUtoztXkrMcxprDXa9bBQjAfFem4ESxjJhARfB+F/naEFMRZGafHWx2E
r9SK96wlsacIOYHQxUWJZv6E2cfUlyY8aLeyMdTUOPfFXWdIaLfs0XbLJo4yw4BxQ0Ql9As1Lsdo
JSlzggMP6lHFGz1Cml4NsMyXcrIvxhO0YzzAikvg7Gj0yyvBD26zPrud3Mm+wORbVnGdw8Z1aZlk
Lk0+v5uyIx0oNcvRXt+G+MwLnBHjDdrgRCgJMmuv50WaCPfTWu7Tbxg23ctjbXm3kqMxLsBOcqoZ
dQNdDh5i/j63vpXOuUBJxUq5t8doP/dNFtzhkuorvhAHeg6JKAdb4IzuflDchBC4b2oJhH1uF62k
LfesllQenQhSvAqVn5B/SGQZK2J/wbFPTmB0mSkjF7ct4hw9whAACas6TIPRLD+TuKtQWOm/a8Bn
zBLx9OuVYk3L6P/2bbKfGt8Ab8Q02Td5WrzhGfaZco3qk7a4eXwrht+BHk7qGGAhZoU+xjNQGkN4
IJQ682Rn7xvzULJqjcuYBMkH7uTwRTRu5ULKGbOawJ25ewQPfYXqBo5F36djn/9uynkgckyTCfMt
nYw6SrVPRkHYHdLE/TUb6eGEY342yBqQD7rT8uH2RpoGfc8oP2bufAKP51ldwLxHPkQJh0iYzo5h
5PcBPCQnyKamz7jYcgFHta5E3s6RvT0Eq98+ub9MMoVhW0of8L/GGYSpBCFiZM9dzmIiBG/NJ8ge
gZINypAf1vrG7YZWOyPv7SU5lHFfo8c273Dg8HI/NVP/BM/wXz1IGUm6tuvmJ29f9O8qvG1SJcui
c9a30jyM0XdDjCZk3Tw8VaIHy7YWr1WOpFxFTQjU9eypftkDBaI8uGhAN2WITVcBLrKVuDE2GClb
6Kv7GMBa0TwktWJ4TxoOH9ZlgcWt6mKooGUhqVWonAlg0uniKsn2CaYDJ4IPu909qOH0yQ4s64mi
FFzTFqnlKV5jMWPoCuea4DoQY0SMEtTe0Lw7tPlg5rw32MNeF+TtYbBlM0LLbp86/bH5GItpv4QI
Z4fVyGgz3j1taRt12HxvRL7d7rK/pvqmwWNExCjQYHqSE53g8wo9yWTXzykiKy8Ct8XyCwL06SW8
XaWXlrbrmglMKF5Kptofb2uNiSo3nWovMLX7PDNMlhOuv/DuFfc0XryFl/mdmf4dyh5WtqelMnNF
Dhsou4/o09ev7Vq4mJZ7AqcCoB7FHR1py2voJMD7PICoA8Iilqm6CJY7hVQyQqxCNnlmMb6gHEO1
rryGzSgilIa0LawnXzmKXC4xeZdQibxL72zKkuE4ZK4gs/IQ8kddxA2mPvO5a6XXr7wpCUhzeTdL
jSQl/QflqmgErMNnPZlJ6agCG46Pz/wgg8EVCPxm7sErqfTNBCwoKYLgNMooghfs16FFijD6Ef8L
nPvMAzFqnnnirrH4V1RcCqJ2rJ8gmAxHMTisFVM36NNMEK8AoZiiGeaF2Fk2q7+WfZENY1q8wVZ5
vja3Xu1AXRKThbAhLRI9ByMJIkElQ3X9pjAealWoYjziFqO4wTAIBd7L78Hs31tBBSgKrOKrts59
RHCWhgyVXp3a2SY0O8e8NE8WBfom8bCAlycN7iiFJuHwEZXWipQEQjgntmbIQlk+zAawtB9/T5ix
onvegW8uN8JyKBiOC8nDE8Vzg7basmr6uoVs/dNWJVo6U0qYLNU8paAY/3f58Hu+7Phee1mzInME
GXlIAs6+BBD2ciW/dW4KGb/873gz0IyiqSWH0zPZk+syeuM9OvnFE2HQpJbGrpId8EJTQqS1CsoP
ja6AMYW51hubguMvzL6A5u5bSRLuH9XulFMtjYieqUjyKHxSKzu4tKy2qtxxrCZcq4Nw4rGM3N3q
7kCe/eTjjKdqprn0m7KvO8RCioZMx2Z276RaScFDL0Zp4GUHGRYu/Nd4ayM7rWdqLqWw25Fb29zK
y7LNDWvUW0TIVY89FfkPLZDYNfo/AKeL+GAYZxwokB+ADLcQAmRiWQiejG+tT/gC7G49MZ6undVJ
Ov/IXAKRLzVplEsDleEwYC3aaKcf54ypRMWM7VnFO2yqz4OMBbAE4e3J/tZF7cgKYXDiRTt+C47U
8uI+jrkjbMm2vjrnlMDt9aDV1fwXQfxp0DIkdG3NSPetoWRSDmdwNTurrERyV0CZWKNK0sLup9hp
tjvP33hKGfULnRc/GzNxM8OVXbOwQht0HzFoQMLKK2uouHQ0KRY12WIEO/2UdKXtEh5D47+Hsmb8
ybEP+QMs5OGPT7hpQ2RBC1lYgDRMXqo/2SQe3kIuZiVNjL4GWKiNGBdImI5RyHllg3CttldqsAZ1
oJnBkKfPX3Zz7M1ZrmaNi0BGJcDstmagGD6CBcZUYYdayfhv0v9OgSPTENZoqh4tXzEkOrjElbfZ
m/foK4+w3DaS/Px2f0KJ4A/ZNvr9Yj2kZFs8KxWhV1yWXh43Rkn3TZQAiTEbz4RoXMwKLCyQkNRV
lqrNG/Vs9PmUSoLyQc/RYaBkXwydbn5g3noF4szFqQ/WIuhgQ/utyvHPopYVtcujA6mO7eYecj6n
UUaBcjXmctSOe2n8eix+6Z8yG3j83RWbmhSTJnHFf5Agqpj7qj+ObsVtxBTiE4qPFoWWCgQC73hw
xonGxYYDkbozc/UaLxYTfXaO1Yc1KAIvW/Wrq5URUL//cynOgZZn4nFNp7B2qcdQRsm/EvLr4cfi
WEKPwiFI84ZFYmgX7E5RFqaLNZiaGvzbi+mPexkzv1IwvJqw2jowPRs2ky9m4lPwvcvKiYPATqtD
m39wsQymOqM5GSm7zCX+2TvollxLmxABj38C5Vep6SiI2K9HXdiomj756MWe7WQaXEy4SL/6G/0/
71MK9kxOn1bTQe2dMq8p1MSFpOfNY3gXVdDGqhoCAYV3Ls5O/Rr2V2PMaClOLzeaOpFgt0QidkkK
c6ejdV6gycEGGLyh+jR0h8zN3CWlstzWrtKLY7cxmvDWh0voKwq1MNwUIfPwehfHdCsyBv+uqlqe
KNn1hxngIsI5rRIJZla94+SpVGL5Hel76y3DohOuobBXpEmu+XzNjAgnH/UhLOU3Sm/F1/SMVMSv
ih2aYMjXn8Geu1IzXbo7PB/VCp5vjq6jD8uGQntYKdcq2AU2lZic4yMcxQN09h3Iw/5FbQ5z+afF
ixTrsPCcwN+bt5bvvnHzMxbIlPPq/pP+oTnP1beXVQ/6cduVHY14iLgxYRazW9pweo7m439IrzZ4
EcotGhOkb2mSyKRz84fNLwYJfFH1HGiu5CDZ6FAcBQt7Niuy4d1WeM8FgB1SxkKeOLCbg7d3hNXl
BnvmpG81irLol2drh7VJS7cdQmqeMUXEvYEceYd0U+Qu/XcPaoWKT4v9LZbiU7Z066rac1C7OXq8
+4xvcfihDBWnG6/bd/dMffrQZHD9wMGWUNaAzqGGTiUBBN337nKaTe8w//x3ohUNnEvBgyjICtmU
VuYWP5TCdpCDqNFbjPfOgFTZnpzvHFqCtaGutYYazHA4XkEmO4Ef47H+IGiQ6fDkrcKb6JixO2xr
l7vIvWYgIC8BdvUWlVCile6rRlGUeDa6DUmjhX+texjqgowefmK/zNZ76Orf2TH0J7M12/vN5L+o
HU8h6zmsgWKrKjuD66JCduWTuH1D+kp4+3DR95svxM+4EZPSMz+dv6E93MVkUlsOqu67cmyohqF4
CZzkbaGYluQ05Y9EEndseUK3KMq7h7HUrfAjuSatwAHbfFwgA2H0aHUNVvhwC+e08Ocus4pU7wyC
UGRRrUDZV8Fzu5tGG+BI0Tt9/1TSpz6Ztn0KTrw452dUlrrU2O/V3xdFk6DhB56XuxoGHF1xz5hA
EKWEQM/Z61YMz2F1ioYq+aefAEoV0pfT1SBTK5YcUEXxAZtGx2Adtc7BWZx3TET50cmLy5HW4MvK
4F1iukV8Q3tdcFUUmLdRUXs6yFvAtcqd6qYc5oIqibv63rTFPcc7W1+0LlBONnVIZtDdGDIR8bc1
J6lCUKnL/DAzoaVlUsDNnJ46TMLdv0BuTP+x4dYWTjyveO7nv6nusmI4K5Y+naoTvgkyPOeePSaX
yeTo0R9qWDlZ7MZsJsorzfbBhehdcFHvxT1sSP7fhDx8og/R2PE2aYjqC9ykcZD7WDKxCxee9ziR
Zw7OyR+rtKYlqjRSJANuK0wsfsy6iTZHPqtk+ix9BRFd/izBT7fFNh1twCqpuym+zMO+EtoWc7gC
haUUHMcJAjEYYYvBB4mvAUpwTDs1rOHER5gCtbrJ83JLYsXvxkEuoZiQkDTVLQdFYmEQWEuEaZ1/
xvRWJ97HIUONdpAUAv1WeuB0gQ+wl96FrSdHVDA/bFQRTErUuyKXfBXhiIB5IOcjDVFGlYe9rml4
RFFRmxD7d0g8c5VhD+ryceUMtQ4pq484C0NaORYS126T3X7eFt/Vk+WXprUnyRatNJkvaKuBMCNq
2Ph8U1JegFXVtwv56Ar764h/E6H0kc9Cy4Fp85ctvmSqzpwwUbIUJSBESTPi2yYNnXQme6+ZXV7t
+chow+kLaoQOzaSxX3jfyn7xqR8fnW1eoTkXiKyZ9l8YwBEzjTuAVmSuk21HI4eSUSZq39zeS2xg
ET/zak35w7OFKEnCO9EjRvm5GSTKwNumDKR+KtYeFNB5E74jCiS1JmsKGOeU+GxO5M55GatlXiiF
GSkQVLO4yYUq5/JOA/G5uxP8vCixqpgvrCE7FtxW/yE4RTrF1aS4f9Pe0ugjria7aIQ3hDfd8nyM
m1u54wS8jcFlFMsSSLAt82ZW2h1VN4XUaMPGP+T9isj3EWhgDcLrHFgYyCFQ1uvlgR5DJy9t39Oj
EB+jswnTjH6PwjspK4XVFHgYLKO6LQcyLKFBqh3yBSBKVxXbOT+GI0hZZMkMnVmuGjV2SqbnZXpL
CzaNOWtPTjFKA6dSamqlSliTCxgKrla8YC6le/Z35psndtYohxJSw/jSmHRL3OVPyOcs7VETV0+M
HEwOvANrdpTvajcCC/nNxVVALWq43hSKfoEFd9hFjD6jXJ0Sg8yBdMAOdNfKTy+hXAafLrVK5wSa
gHTTkRsts1T1nUc8wZYWfgvSRpAcQzIg7YD9hF0hUju8SYP8yQCvxYxhjEMnkwbJkZBsGBrfy9B7
Auensq6ISB+RpGN+x3nXWOuu4zTzZU2lKr+xnlvK83YltgTHcQofdaGm0mZV6dFKdCI9RM8lfQCi
dpsDdNQRqAZypjP6Z8rqafJ/QkmS6LI8vnzeor7AYk7CC4XHEVgFtW42B0F2rNjU2gbrBE80rYP1
07WGvNLL6sy3+yOJ0nbP2UTeHfAQooOxqjmo6Krh4klvPNnJY8WToTDyGR/QWb5mZz86omEgBlwj
dkIqFheJK1LRdT0xPxvaqbzhFJL4q3ZbinhVqYX8pB0aPdphT/CWtXGGzrhuGWm6SP3ziw+FPwPj
pZgh3H1CN4PVqSKDw/ICjHMBQxvAc0ViSCUca941JFD+CO+dA0zYftcw3MjDEHNY3kx1IyhGAE34
EhaBTqO6V74OPdVdpSPybsr6vurQjrOv+GDS84boaWo5dvHb6BhGiZX6YkWWZwlr9QbpIODqUx78
/IIiZvLu5jlJh4aCQbP48lY9/A9EjbcwG92+gaKjE9YIBUsAaDJ2qT0GbTHQ1ILIMMFaJL1l9w06
UjkBPBEzglm1ud8fZ0nHB5ZJPRtfhMa+LuZrEL6UIYNssrkIACTbVZRt0G30+ehhIzPe7XDvqGId
gORsJZEeJMUSzl8d+tWktbjRgNPxfU272aZrEqeui2N1Q0frSX5xgwXXQg1nOxuSENAXyW09/GKS
ZoEbNhVWaXT59kKIiArnRBxRXUIm4sqSNhBc5fb9nrVkx62Fwl85AZj0ZrnKEoBR/qAMfvLUoTTN
b8rnbFZdY5kd7EjV5xI7edSUHBVTIH4C9OkUSk3luMKf/1hjQaSxlWybx2s34VN+pB6TfAYJPLxj
mJOSWxFKYlw8yuDwtrkB1XnLKmM5Q+0LPHNQIYQWxwpaN/a5UwFMU8ea7atGBxHHEBXm8osufjMQ
u+oyfQVSpNz8REbfGsPQUL2TSIi7bl9yyWAwE9VF78Sr3T4J13vOTckDcHLNPL3XgTPFJ04kFGFj
4935IkFwn+ZiXbA2zVZ7P6ecUDCUg2DfFR/xolDX+zM+1U+z4OIUArQohDlXAG7lfXoVV1M4RFS2
JHL6lJxQGna4YwyhrQaN382K9WlXAjBC2UKiMILu3/Hx0f9y7cXlYi/HZKBcb8dfSQ9MpvoyyO9C
yWDPnJ/h/7kXY8sxh0EKnUFo/yPwNycFaSNiCyxyjaxARJJqKxDmcQGqedgK3BM3XBXNDzqdcgc+
xYY+V+hz8tRkskBvdBIjrvE6bgxHEnH7DNmb2IRZBDZ843ybwvIPwvE4bL5oLvUetZsNI2ZKb3Zz
L1aBRs9GZJt6WMkV8FKWLV5fTkqei33f9UlywkD1O8ez3qtzY4tnBdAfyGJrVcmFddKD398wIcCY
d/b7Vu6BQbLZu8j4042tXqxUQyABoee3KJWjwcycc0zPyidPssrg7m1FnkZ2203+INUPYiR3IxLS
hsfV7o2BoTU9S/fVYAJX+tR2egyZT5xvluzMS6PrW9LBWOh5ZlNWXrdn+XQJFWyVAtBlvMIhjSj4
YweZitFAJeJSjXqTMyAAWsYDHMUY7/iKZ7jQzfYOPfv2eDU8LAEHWs/kptNiIlI7i6BygWEbAYIl
7MQm6oLR6aBUx6z7LArOR6JIaLAMGrasPS8TS/SjECMeprqJ9NuLeDUS11IWTqdAvtB4i2r9Qbb8
p87LzONZZKFcFAINV6zTXrrYbf5GruBsFos3VRs8kOBnNpfzyQo13aIr9VuRW/G2NIcB5JzBjvSI
dcG3Rw54H/5vLqzDM3h0PJSi8MOk3N2TMGasMH1G8w5v8xN2LiqLHjgch4PMj9nGOBlcz6xqu8gP
Ddtyu6oFm4LAlPqmCtMOhlsPmWf9yqlxG8ATHyPKaUZes8s8xp7HH8ALevz2RzHo4yrJSgrmoUeD
RJN34Xyd+Fp0zaqq1bf1WYno8jdD6o9VM3nzg2e/D3oOsdFbczCjRvscGvw9TBdQiimhq2fuGx9J
FEEKoVbX3vC17rc/F5aM7r6uXNLlvJekOdAK4ZtDzKqUUzWAH3yEmgfc5M6OjbPwOMUhW+DEH3PR
dB43WefBPot7teLwA9f4hYbwBUvsZbh3rIN+tFiI3OdDmHxcmlPt3xGCoPMkzQ9LvgszCUIDb0w6
dNSGiI+/JhuQ1BpFIdpjXP13Fadq5HmWkdEa3YkLWqkPwzWOo7wKxh63UlUK21mdgMGWhGi475Rg
NdKEzovZxsxnyA3wC+ceqGgedXac5V4klpNtU749kCoKruTfFX+y+UX2g6lNAH+BQsw8TM+cDs9M
snIudhSYpZsn8vC3+s6IXCMdu/ZvkFu/MuquCvyBM8QFSeJ0dGSMdE7RUznok/Yh4MZnvqmLttkH
ULoXV1FTmdyiiDk98+CAoQMbpRkg2g7fuvRowfFnA+4CDsZPhlL2SNgIjBEPkegY+Tgw5xZiGoq3
75lkPdf60BcnixV9uqM6Ss9Ux8aiNJAmrOLV/Pa0mjafvTbvIyHnTbKsODa/2JtY9itNYU0E/v1d
JdUeccNX6nuocYUn3vnu7iNp8Adl4x6EmYtgV46KbqLdcfsV3E3mKJ/SXKAIY/w3gF/b2YHxXiCE
mlTofNlUShpovKK1UQ/LTrR5HFg/FTeRa1E7vbct9uyI4hMhthP+iX+Rn708PqOh4igLHUqnijGl
3LhU/MyM94Z38SdR9ufJBDOAgcU5VfPC1t+T9FDpjv/kpL5R5A1jp5S8ylcVHPeWPJCtdowBGWuN
KX8Hu036yJVOE52tpshFH4Ws/G+NSi79g/ow8jc4KUAsjFltEAPUFZQkQYJ/bPidXCtNC/UyGbqm
vPzux4qZGZnKtz8dt71rf+fYf9lIdWixSpjQH63sAG3FMeY+rYXrhkHGB5EplRaJMLYdSuLTF7E5
upTubecL7ntow5/z9oTI5Qw5QprrjCLYm1moDgNYIZOuYxG+Un0zz2wD3JPLwyPeluX2bQZ8aYLr
66qyU/qawzHfhb6e5F2Pc85uhhcLiHJ4TW0NHXp9pkcfL6ynOoj4Sxc9cETFHE9QfgA/MHNA1AEV
0tDVwsivVu73AE+Fc5wGeF9ktFVcgBoCae1tOpyu8sLUwJencbZSQqN/HgNHzu5bFQ7VS8ujyBVm
5O2WNi6v64lU/UpFNDwqjwZuWWC4GaOcMe9rmEcKD4wwFPbo6yzcGH8NteDWGbyWd4a1rTYpZ1LA
RRY2RF3ICu9ihAKvrdN60dQuHGBg0KfuiVtMKJT6aelgP4sFplO66ISSd8V/fdCP49cRaJVOdmZu
I5JYuQ7p0hxHDkkN4hEyKpV5FSeGsz3mMKdP/Ybovhntywo2AW/dR36lFwljsYo07JiHeBUXSzcT
ZV+reAsJHoDc9ukMmXKCimzlWh6G+XLUzsewvucEPq2ZFRvwDNM9KOwchVBjEaB2EWRz6hBM0X7y
KKw0kRIUAH3vu1uCHThaGUuj5PgXslVgoP/8SkigGrx6monzgs29Ihm7cJtDe4SEJlWQJ2d7u9BH
jXwV39glNatMo0ldQa9SjKpuAu/HKM9MBzyWTGIR7KsHikMvEa9vGc8UnHI1qJrtiOxa34S1XhFV
oz8R2sIyUMbwDYHupkcVyMwPthIsdbho+OswRrRDAqQOnD22XeCjJrxHC43MG6A7X8WuX5TPvVx6
40O8D7say1Dbv7ABxn0D6Fo6RqPFJ99DaSiYcgnJxui0yhihXtIQCd4iQhCEzPOxRn99rKOZhFVY
6i0w0WEvUaNborzxqHk9MvBhdDudB0vafvfjd+Hkh8cXB8TC5y3WIdqJz5wD72T9ttNC5GSloRwD
4nGnts9Eg4kxJb3j8M7Xs7C06SMPMIm5BfdJjkvJegz4eZjCvro/xm6QN59hP5WukDNd8oyj0kuk
xBIfDszPGpfFJUXNNHPKBsgM0BTxZ9r5IkRCrALFsbGDFJx9Us5Dj5IzfPH1g9Yc2AkpsROwGpG9
AL9vm0ltsuno8Ifz9xXtvi5NVG/VYRMJl57XhYyqIzc5jCVWy1lDQLXS169Nb6QEdQI4R+BwdZtH
r+ThcgdjzZqcBJZWyNCAkU6Zho/QQDVTk9PNDztmpTfxbODTREk/Pewt1pFNIyG+l5lqEGN6ZsUa
31fYId7GOSNxqQ/CzYf5B238DRGzwGmdoLTOiSwccJ8nfnEm0jt0mIspuY26B7JfKKhReUUewbdN
Qr26bmNqHpUWlQLgvoPG1an9iXexbgAWCFLVaoTCytXbhW8FzpqIliDbITnx866NCcztVU7t1324
fp8cRcJZQjbnjjOKLELolDOOedyi4rWGq1OLKneWEauKyul8W1/hhDkcKs6IvFWEJrvGc9hxGfo8
nxJmA/cPZgqa4J8YSH9fC1xiYKlzIhIYgk8I9id+iO9PEXVIS8unf00Y6migmg3tNE0UT+W2im4u
ar/rjaY4+H41Z6Z4ZduEhYxeeos/P2dy+wQm1NiC7pG4oZc46NWyxEC78RI8Tqdia9QaX/DFT1qc
lsvJcNg8CA5xrDMyGwRYV5bvdT/5XKHgZG/ZIwR+R4OR7Y8OoutEJwDkbjOU12JQpnreqaDNJSyC
y+KDOHlyfJbQNxeC0hfHjMyMYb3+IpfkfSRKzzzf11AINZPoQZo8Eey7PMzacMrNZBTSgEyAaPFP
2zov774XWSoB/iP6LNs/RYyWM2XICCXcvz95bky7fGFqL4EcD4576W0tod651ny0Tm32oI7AlCrq
eMqelHFQnB7E7AXCYE2yyDQF62n45PZpPDfZea+wTJN8+bgU2G9ewnHEsOUpuXgIbp7WQWeVjl95
0UAFyEZ9ev2au+Ay8Q7GUG727CshO9/VXaqrLxTkd45ugvqvJKznub/lC0LIrlI5rN73ElQsLO0h
hc3GVv8TCoCj0c7n1b3fb6w2wG1BWs6qzG1vIcMwGsVjBjDQgeTo0JbMty/Zz3Y8DlFTaH21AthA
M8J5p7H6/AQCIWRe90ZUefbeHBgrEKxO18ZLPPU5dA/pCIDSO7o12wvBI/emPdm+8aqHxjkEGqHV
U+fIUKyptjwb8AQttd5zShTZNMU71y9DcfBFPR8ts/1U1cN1gLFj2WbwJZZt5KL34v2CNkfC4IXZ
5E+pZpC8eqKOO9RFdvTQ3zmj6TNCF7sZBMVf6QyPJZPws7W5yTWbFBiNQa3os/rFMjeUMl/Xmg2+
BVNtwlCXd7WBwah+8OTZQ/3/NQYb6DRflQrfGVnV4y94jpE9tQNzSDZAvk1ODA2u+sI35FncLjmU
Oykt1haQgrcq0YWYhJzqR+ww+xDPCfG6lYp3rd4ffEvR8xOdBCZy0dEBgIRf4AqED1yYRekUZKxi
rxg/232u6tjCEUjPMgu3Fy2FLgWhXIk3Ilvq1ufyxSrFzrCJDi4XNz9UQQbk7RhYfLM5DcEOhItP
5SzZHCMDM84OWun3UJ8+NWWoAoYavAFNfREFJf9SYftjCxUiq6JYd1ND8ZtSuTAeCv+E2rewHrve
r2YBf/BXvE6vizynpkV1O0IfVeNZ38A1pECOkhwF/odK4BBUPLE+rceX3xvSM4shvJ32doPWbUWn
sToSn7/Mfgr72xMqM3Abf2yc8k2VuPI8cdbX9zGn37akTzg4mJIvnT1kYQg1rs4STyNoTbEYiLyG
dsZHGn8+9zQUGyax3ueTSeuHJ/D0D/X0Dubuw1szQdwzvD62t2DGPiUEyltLCl6r11JX+Kh884K+
m6Er/KlUPXAyHMbWQaPHAI38cLuhfOB2jVx2XGomRiovtD8vrggLKIg4xgDqUhYUJvn73Z8H5kji
5eMsgsTMJJ3HSwPxFFd9eB0MaqOUeAzD76jl73ABGtPoQ6n+1ffY8qIwVUefh6MZ+4QBRzfLya4R
rzrdsAIoWwYqeC3cV0Hdt/7IA2j0Z/yRTV2Qohh57U92ZbJYyMbvldgJNMcZTlkIiSkuun6HtLZZ
+6Ise+eh1yurM14CcvmfjO9wv43No3SnZ+5L5r3ef+SLPtWAOGAG/1AKTzmProvD+MiHX7I+yCd9
C8ZkvRSEePMFp9FvUM8oTY6LVlv/YGlvnOBpDC+OsEXgsZPzyQBLo91vDWOTl5l3wg85EOTzXGaj
SWCh8+pDc7nLubnoj5/iG/I/MCl+k6YAl8fvmA4g/Y0aaE0flnk/l9wypxgr9GFyMxSPi+UZ4icM
bIyIsK0qVH2Q7MgYanZPAkQDmToVt+EyZfVtWzxDLUVS85XDswwRJo52hXLKOcxcr/c0UQFzdCFr
1/N6sl7unSTjR6Vl2Rrn9fCodtvVqpKua7SI0fDpr43N/WAsPPggHiZ2JuSbR6yFqN8TieLM20Qz
Kggn9LXCYr5TjKPt/cGHuy1tcPdWsLzxb/ziAVEHeAfknePq1+uyIw4PT3i6AbgDQI8OU8FmZ9lA
I1p2Fq2lqw5Ubd6XHfaGnn+aTpRn1oSI2zXjfzQP3RGelxhaXg7W32WeNhq2yk62sXerloB8K0H7
HDrXSkgkBWErRu0WXobuUp1dMBLe3rkP21E3VL+dJGnAfay5ruvyxOVQJu4eNM/z8397hMYtjMjM
JhRfHOdq+81EK9y8tf69NKc4UvmSmDIRuC459SF76pMWu4thISgxna/Z28SC1OacUPAu/E3oZb5B
s5PsxvWKnjIf/HaHx1GxbXkUNBwbl9VSwgvFPx6BLVffQm3uIuvpLkgypFT/4g4H8S/MUDkJNTk4
TcuMel2gTFZLB+PjeWhQgzpOer8Cs5G4m3w3cJ2YJ3+TWRZ+cgTXchIwTwpmUSJ4X7PLv9mErMLK
tTIyGU/zB5P3RaBw+Fu7PNsAM374HPelc/wHoj5IsNJfquzo8cSE8CpmbcJi2LvxpQDm3yhpNlCc
V8ICthPUidxegZYJ9mz7WGAPci5hNSi+N0iMI/fBvw0COWs/xi9ZLIm91NTbqAUFbc/EWv/h+XWZ
84Vh9Ob91tiX7hYhFqfuUEqvk6Uu4hhVaVs3yjVvpCR0XHtatp6o+TsXN0d78sz6l5MQoMLuCTot
DdwMWlJGRW35VLBIEPJR84XsD0jX1hbizjJGa0P8Vl+f2woANYCfDR8ZRMlMs4FoVvZRF1xqyho7
ZuNL8PFlEHT2Y27gxQs0B4eXffva1HmbeEljyzXWUHL0DwPMCDn5yHyiX49mWIOLB9n0TSD6nxs/
l62mNxIl5sxI17UTZkl2FGDRi8nyFQLFYu6WSXE3vYw+kOJPkhlKosV7/dnK9stFZZ+IpLrbZhw2
wvYx1AydTbLhE1SsRG1a8WJQ6sDEIkJVZWLDn91SIBl/q3Nswgcoqjj6N9KAKRcSe3tD/VzqqXxN
NUHXPURwrNAW9MIaEQYXB3CJg8DhwscMW539vNqj0ZlngncXAOPfWLeIukFSE2Ju7Tvshz23cOfW
+hvDWIOjTr/0XRTNJ4xBQKaK5Vi0uUjtz/fm1mBPeWiuo6rN4FM/KtD5poOKDJa+AklQK0uNv55R
D4/8qmeHCY7LzXQvmPhBPbVqWtFtCs4U5xVBdFZcw0u8ZO0ikPY/gEz/Z4hPjLA+P3U2AV5jyGor
JzRlPWFrpCbOMh8MVLNqREHaqAjNKtehtZUvuMUEkrx8iGqochbVeQBY2cNvKbPZf2F/FQxJWf/C
6+rPGvEIF7HDRpbNZtdKbRdVl7WZE2xRqEjw71nbFR22BeZQ2l5rd1Y/tFeFcDvb79/AMMCMjCit
yutyL5jGi5MQflmE3gxCvY8aNWTwVVBr0WRaUfYM9bxSFdEV+8/GCISw4Kw991bmeydDJp8igbQc
e+2k4yGmJBbvlQVqnkF9qkdd7AdP2VVq8IpshZLkwayhKSeWFf+AoWFb0qcngkBrluF+k9rMn+nM
YgwjhnIUDDA+SGMPBz7AfJSbHXBT7nfdFG7PTIBVzIhj+6obqZCA9ON5kxD6teCf7xuea0TqOOMc
i92HB5E+NEsIZqdJSe2noMxhw2AcxWJwKTQ6eDurMKIw1deU51CcUPMeJXGRMxYLYRa6l5/jxJql
IW56+DlXAOXepMbSsmc2zXiqLfiN0aeR8nQgt7bDoEMUqHisRAZaXRMdncBWPuHWsIPc1xZh5nHS
FXcpiglRUDts3L61sGydP0dvU2w5zKInx3pl1t9vVRazfrPrZuL+YtiTYy66+Z8xSGZ/SPx3oORz
/fJEpomaZh8wQfmG4664jiM2Rmx7Rsuu0IxDttpwx3agvn1NheBH3fmOa1WzBV8up96RQDyeyzJ1
TQnkBcdEIwmV3y5ifYdTVRbLJkfC63X1MbBTXQ/TJUpbjvcTvyxN8I2IVBrmINHRKDwONEoY2b3A
YwZ2KxFd95qum3J1XFt49zthdbUfq+Crs7BHcpygSXdVMQLj6yCW5/afjolb04Oz/A1RCdgxLJ6m
MYtbhKrXgjTzrW8VU/RCbrVnsWu/BIeNccryFmyHxirfCbFNvHmy3LisjHFV8M3T+tCMBnyf0Wd/
Z2XB0ppWRJ8EiHH1AU68r7POxmAdOzLEYuwT1+Ja0mY6Z43tCHL2NpEBxZhgjKNnx3klOgKGAFp/
YKJR/gWSYRWlq8jh6w2mt63H+mreHyS3haqEo6lBcuexG0SMK3dJsRaqkmF96wnqXQUHFZxHFXi0
diVO7Uom/p0tcvoHm+k6A30Pq9SiugkAE9NN8VX1G5FSyqb28BHjO+cmYQLXivlZAakQEbR3XQX+
r8THJYEJXi28ZSJ/Dzh2APFq+d0YWH2dYXJdueob94Oee6QQUHKuq1v7RyYiBDeS+E42bJmboy7o
2COcuCIVsIkFeDE5GAQ191gkAq0lUT76TTR46uX6aYNHM3mHY6x2edNVvjs0VdF8hInqXQ7f/Zb5
j7bKrPogXRZNseJKxixt/sSSGp9Fokl0lwU+6wa1sBogP5phlQFR6hGJLgbz+K4hke5zYDTjQHpE
c5XdXOfugOGggM8T1ZtFf1u3KOPRHou765bNiVwEPO9YWwHH4o57Tqkf7es6oBh1TY3B1EpB58c5
7qxUVR1Q3BU+8+deKcqOhoqhEUthHRW8IPOvOZ2aH5JW+IuZhyH/bRWOE0L3zamvfNjBqJoNAZdB
S4u6DFYBVZfCoC1JRhNOssnIikv8FfyijVhJzmS+V3lFG4hYzsce0+v3iR2rfyWFtfhURXOZBygg
hA0eZ4+EXJqVmcRYhB4UC5t+HP9zCRzdbnb+0ZMNk1zIIQY+syPJ/u+ButV8ilUGN23SkXZAjLXz
yQn9MwjlcfHI6qCdBZzDhvE17Fx7vqK30aOYPouaRJjp5MQaTGul7zaKNCfSIQgkKV2FlVJmt8QI
+QmD7ngt2aquV1ViSvurLdru/jRf9SNANtVCfLrUgUXU/+diGUG7SLXCGCRwC9bgG9yQ3Awx1Cme
YZ4OcfxVdL5jaxlJtGUNBrXxbvuUEzAS39I4DreDudVziBRESIdb1aXD6u6OxGxiydt7u/tuXGIt
cp3fNjwHYoHCR+6Wt7Cvlq/osQUTonHFfhwDdm8EHPuLdfyEa+rncdSJoQQypWhFMqYh1GM95Usa
4Yq8SqG10jRArJAPecUMPtvPjaH6U3THOSTplVvuvUh2i8LOyB7/jO2eaPdpV1YNV5daShDJJZpI
G2rnUU2lrOi4A5uC1//zmfqllyW2zxMAPMrn1qdothoSO0z9wOzfWkn9QNbHvJNc7vaLiZF4+Bsf
xwYlaAYVosWhmjfBZHRM2iGJillwxc2v2OT5D2XF5zF9kkndqlivQJlw0HrDDVq8vutD2OGZBUdK
UyHkQKnXD26BwPI8enlAOn8DMBPEwnwPkTrpJyqFDpaJvMHDw0C/rEeLKruvUdDAY29mF/0wYBYw
iie6Bt9qKIjn7MPGNcRM83QuONtyyZfAxXyFvumjRASinK5O5xLFA9h7fQTimArM+asjlpNEiUmM
YfeX+UR1NGollTwe/wp362Bru33kA0Rpi7rTuD+ZiT2Dv3Lyhd/7Z63Co6KttUpP5OK61Khevm4b
3X8572wR9ddi/AbmW61JSMuuEVSbBRNBWmxdjKu69hpiNWKfGtyQYTY7L4sWBJFJtUaOL0klyRPr
zzN4GplOBRgJtyxUuzRRVlVaiLvoMXJRADomf1qVL/Rm3wk+f1kn/LOGps53ocIIeSrewDjJEi58
nKTd8VJMC14jmLtekd7i//U0Apc+W4sFrKd+jk5V5evdycGdxljCCWDev6GZPgOZai7RipmHClVc
NQS0Mg94fZ02ofANV1FBc9YiqPiOcnQT18cvpgYKz6aAqho2Vx3YzRlW/0zhSLhA92iIIX3Oa7E8
zQns3+eEkL8laO275md5gykCPH5ZTnKy9oJu5R3w/r5bmly6txsnUyOnKHIxdCJ9bOit++Qzknki
9FTusqwVGcaj5xcSGjp3rG5x2kWPM0E9rSOob64hWQFtzqB4c/wdCDk60aJLyJf+oSQpKF87Jg7U
9N1RwoQfW7r7+1FfgcBYT5desfkbS0IbhHU0PA1OYG/3x52GvprUeAKRm93pa/LTI+Sqt8Rv+p4d
xmYzpYGYKsYw+mpfF4JOC2jdJ395PmljWfG7jFsES19nw5VfLOLPLznhh7it2YrrQoitQecpGh8G
dWJXRVAnI58+g33dGERVuuhaXWZiDXlzDbFgQ78Hzcz8h2NFGY7pS7XQVmeWqhqgOoSw0fBrnI3W
KGZ4JZQgyMmKkDR1/EQA9Umk40etc/dAr6D8XqZCV9QIfU4MSqScYX03mmfVTLSVLqYaua9viuH/
C1pAO1hGX0NIp4SsFKt+BUyv42E1hDL5QTLMpeozUu/ukxmuALgnMEdCDoK8hpA6H6H7OJPeq5KS
ef7kqtzUpXKCGD0Tet+JLW92FMlmvMoVCevwgNwz5CZ2ZOayffiVuCz+T2NKcIk9vcEw57rAhrx7
/QiLWwKYca+uoHV9c3dHLTlikNj9n8oebmacfA8gRJuway80VkAaPKLp1EK4K5c6bRt4rh61pC4q
ez7Hodleg5VsnMxbZRL5LgjyfPSeA/5w5UqoyXeVjLjFjvf8TMTNQDzzJjhU1c6B97Uhyt5+8/WI
7CPpOpu48ok77cIOBicjuQHkq5QQZ2bH8c0+Z3pZm1c0XvCuZsTmxh4H5xd30oXiCVQFNTIZ+J6i
Zh8wbsW//rRM32t+P5MiwP+iIBECiTGVHVvieh+3A7MPz15c8lR8McGoJP4wmrDeDP706lZdkH/s
NzXRsCIHCJ6/s0aiuoH5yfyGUlwUSIcACFoGpUs9UVyUUB7OBT6VxXoLX6ueR42NV+OWmDculEJ/
f9jpY4zomdricDCG1E/U/4izxnhb1W+qlnna6Q1hjaTIwbXwBYJ68hekuq5yoW+i1lIs/8XyHlZ/
+7R1/eSVizs/cHE5SVESl/EzE5ebsT880eALIe8dT3P20Wq6jnW0+Bmt+ZyV0iQ6l0kwxsgjrP8/
FaJrbnzRrqOTtGTADoGvVoo+xvI3ya7kemGJwWRT5r80gAqZJtPd+dydvIKSYUJqvoE7MARG0QNn
eOO4vL0gJPm0I5vsO150ZeOTw4W5bf/LHHBnQd/Ow4hhxlxB741E7KuG3V3gU1egOr3/wvCvyfH9
RkWZozBJckqW0CekKR7zECEkgDF0eaPTKxx21rsJbqJ9GlcBWddroXp6cAqmvSm9lz6H0ifwTcZA
W3Fq7YlxAHIVNFCRj2xqOEj2WuPB2bBKYpqPqcX0XeWleY5wPG7LBcvxwITBal2xhD5JUEPFO9fp
pYWEM13/ccckzkTC+5xZxlvF2yK10xyHp6NFWrqvhSkeyaZ61vAjzZasrNdpZX0J5RjsC1o2DHG+
jVx8C+BarBvrk56oqPnqdShJkL5tOOSUrpxj9d/VRwDK0xmHdfADNnb1S30Cc/iJ+lcVAyHJWdHV
a5zW51flgXkvhyO/IZdJi2YzK92V994E+Cx6Fm60j0oeNwyJaAmbPhbJWOpuPiPDolFIeQL8haK/
6aHeM3i7IKIHGXUNLJCZjEIIrXZ1xCkwLtWGS//8Y1Ba+G2w1CFdX+82ZY8FcNBZWv/8NSLQz6me
c82gmyMVYxpwO9okny4MFXyx9k1UR2hcqKxnOM+/CgQSS1V1JGKTVU1ZPmx+9HqUKkdHt22iTu+p
SUHEugUGSA0lNRFrvHFTP5p0dtCJUQjwBNT7sLK19iIo2aS+U1Tl+iJ5IUZWsFrR7WijyI1x+yOr
/KwOiINBNkzdWjuwC/MHkWUboGXAznS8hTdFzCSrmVV2CHZZinsuLPXz9MIvQOLUroRqHeb8mG8H
6ON2N8aUPdChqttkx/JD5vozQoy82H6bsI9ZZhl1DZ2J4Yu2SeF5/vXPMyTvyibsW4uiveinvAO3
M/zoEg9B4rZxCFysu4Vp9vsuaIiDYmg0E8DXqMZMzd0X0r4FLk9ky3TrER1+LkRTK6MgJAwArI0A
Z6eTeNdXJb2RfKXJlR7+GaVKuhEaTvzQ75b7YWgBIcFo8W4VQ0q6PTCWV+Oy5ff9DfYrCds/eMwc
iIB5aoXeCMA8Z7vtM6z9ndiC434Mtpklee6U/uwPtN/w6dtibwbgjZUly990fjIZ/+slEYrSEeVb
Y9jyqxMu5yTPTXgkKYfpNEBvOacgVOhgNuLcV6874Ns4qJdDA2nGiMjoEk/FeNXk+qPrETLQXQcT
gAyQH/ZfK/Fz+pOqxXjpbKPBKBvfDTCIWBvYgNJS78/1vE/T/5UOA7fkztH3q5RDgozNZfVQTeic
zVJGb+zd50Xaq8GA1xqFgySNEbRQpnJAxFDHEUBTdIjSCq1CVWoqw3BoDwBekHMO6eXqxDoP3ZSk
SB4zjfkRPOC/p567PmbceAJsTdW2tCFvO2dKrquIEAdhqbmPuo2kWVHyFROEyfrekPcKBZwckpXy
ACdOrTUtP0MuNmYDvrN9fBQ4LISdEDwWdAVuQ9VQ4ML4HSf8plulWtatBDQJBakSq8iHxMxnyVk2
njXkCLPjLCbc+/YxW1vGJC4LlKlPW+FssehxyCPVaucYFyiV6/9WqGXMC71qDSjG5XnzNJvpue/D
YLUJCjWWd+Y68FePpwjm1q/I0q3Ty4vxoNKDLC1DgcO6MrgnGVeQYHVh28X0SVNOHzjbuXjB0vVY
8TQYwTGNmivRSMh2mjrqm/yDQafrnISEd/oIRiNFArFNXGasOSWwcHS6Iu5V7p4mOU8RESXspnZE
UY2baFfWAySKfrxhKHV7gjWa7tAFY0Rm2L/5JwC6tpvlp709uNIdRTqd1O23VXNA6QSl06OIjt5c
FCqtKA1eebfqJszDGzKVB4WGu9016FuZjlQ/Xt2m+ohxx6M2p1UOIjRjMfjKQ1TPiWtaKFR9BhkT
7O/7iHpCZfeDfHqRLBNOg6DG5reeXset2T5uCZEPpNBcgXB02roIpNxMTVaO+j0CMsf18U6FVb2S
RgmL07BnGsGwPlFaiUIYpoqw59jgoI9xKX90JiYzRUumIhTPsmsUaKkDFty68aY3h7fkC56zOIoC
wApVGrDflMjeak02qUDSAS6QPzGoaQZAUutBdduRnH4yR7rlyGncKLjez72Cj9GSXicXtbsDabdU
OtCYRQV6FmygD5EDYrZVf7hBbyulczDS5yBvvvnNOIWTPGORKi9MJYFrJUsGoDpZbK7PHtdcWuVd
6SgzWb1ycx8tcGePI1hGqUx9SOheYx8Y6JwG23VSwdK9xUg0w3UkYGtfgoCSQqyIutxwoP93S0im
FZynBwemp/2gxrpHQWOyn4+NxWa1v+U41c0LO9VmotOWCXSaJV4Fn1QhzyNJUGJ6pzIRaMpDbxLO
tn7XAR3FOjMgZkqKccVDQbidvv/7KyoqpjhZJ2iLmeqiQioQtFiH8JBbfAPYL6gF12KT/H1TLQR5
EmMmVJrU8YGAY7cCs1jVYLv+237vNid9f/nozCENFtpzFYDw3TqXLhQphQPO8AW0gHeH0rSk81PN
F1YTS1X2a9WqTv74V7HahG4Axo3NPBHfWVSaKDMGe37W3mjWxc9gQT37Oj74QoTXRjur58smEjhU
4NeHvO0VH9rKc7syIusAjL5J1xVMzxNvxOQrAYZGdeDXUb+rUYh/cngBl052hRtuAXK8kHA5bW5h
nC/jK9jl1DPDXhXiLRxtQlAEkTxXXx4z+SRclH0xyDwDAT8ZKMaPCaXozFrSRwXLsluOhScN2fOO
tycll6Ee0DDNnVkzmDxmvfVbLPv9ATkqf3Rosl4gfc5SIwa4E/0r8WBrWLWmQNpZtghoE8WG2uti
g3fD/gg8ICQAltnvzDU+5kLx+wTUWzgkPtradl0AvX0MQwblQvDyyRsPP+U3oglXAH5h1RPYbbn3
8oi6JwXX/hRPnmBolFUWiQVjnt+Wda1e62pUQwMO84/gZAQhtoqm91lTWA/L/ENQsbzP1d+dSE3F
YxfWDMwphaLnuds2gDP8K3WOr3YOqKVCktg/Of7jsrxeuIFnmP9ErcPAbxtLdcYqswBDlMEkgs82
3GsZDHXjb7qWojKkxvOgXDADCFIKlfA4u7Fml1x2Qc1N67HZzYXdpftman6dEXA2Rp/PlSNyh6nC
tJt4/a7K9HNm0Q0omckJpwSVSrmTCS2DCbTE8wD/cqAqDMr7KMJ8nr1MJ2eqkh82J20Ct8MCmz/D
AAOYVq5ecSxSUte67f4l4gDIoCBBzVLHQa9HIDkZR3Pto7k4v9RqtI/SfVXT5jV67jjO+v0c77S4
09J9gXJyH5ukFwIDMKvmiQ0Q/SvEZZtYlB4LpFF0IyuOu/CSvpic3ibKg8AonPoR/iQcwpjfnPJ5
i6XyaysV+O+sZdwdK8jBCT7XcVhkdQGpwnyMfjMq3JvAi8GCYILXQfGmGiFN3XCZHF9CBe3Acg6Z
MkgtqnllGdIMpyaFxbrgGZMZRiowARetW0gWRiBXZ4XO+cmHiHBqQfK3XxdXct7DGUnN/savcSRa
BBAZSDGc35bBJnMHQDwVtIbLMdmvmaEndx9qj6WvYVFkhko1O/M9hJDx0hSgEoIJYxhKhzwK1Qez
kVBhKHb0TcTv0CFJo4daa9nmS63SgGC6Za1OTpy6YIgRRIlT97H4VaQE0RMhR5it8mAvMNARPn5t
uc+jkKObarjS4h0y8wPnyy7JDbsI7thHZZJ/A5jNkIRfVovBTDBtcjutQpTGkZv3V7zsXoV5pCfb
7tuEdjjN1EdQLHE4Knq99wIsH7IMTWgQWOfOc3IWJXNyZ82/dN3wdVY/i6fC5tTDaaXdSKLFfv2E
oGfcJKHT8RuSDFxZU59/AwKNcsrzahAMkD2RoObsmN46jPf/Lk1A5/+xf/pyEQUMK1xPD2V9VBSp
Xzi2VD3dOhk4sdI5JldU0NmSf+iJyNwF/tBbPz8ObLw02sH0z4SC8ZXbrojwJ2WhI3QR+nf8P6TP
7z9wWZD0IKC/Lo5b/oxB0NcTQOX7FvYTGO56t9i4VRz4xuf8Wb4DhuobOSniQB9PIQHot1yCPiWa
5yvd/6mo7mikBUKF994KPM1zih1AHWIENdhHL3MH9iL1h4EWDQ71tazadYOPQ+IAaaf0/v1CgrXC
2xQ2di3JCj0zv1CwMmbh79hqS2CAcM+0R76KITrv8ud8DRT+44fcQQkdzaaHtNzY9KKPcvunCrZa
DYlDKYaYPDG/YcDEAeQK2jrvodiAD3OcazV2ON1ekRLTpVDr7Tg1aQVwZekGP4bew38/jjdFKBaR
smoXctjkdJbFYHRDRf9mVINZwY2LalpFerZa5hpHSImHO6yvP5z/P96fhQXuxwe0Muxge+db/5kX
oSuN1qXtBkoz76lIxPSHUUr7tU7aYTsxWxhFzSQggaIPN4NdmqPFvDWfzmwSHTJZxl/e47JZjpyX
Ytv71g+F6QR7m2TdQDWz/xlvOSX+9PRvFbOtrGQX2qJhC1zOnNq4Hsp1iN8PuTBDv//LTg4KWHoo
fRwhntwRlX/1mAazzLWPXsAZBk8wnzraO0JKBWxyj6Qd8+7s/pS8IfRTCn5pLRYzA+EPYe8M6qFq
gfWyJTHhjiN8XxYyJunddvwqOj1Mz17tRmST1s/dDAXPUEwEHYUjp6VyvnmN3bl19Y4EZZ+9pvP5
L3f+r13OV9VoXDxpv0KwJKezHeV13N1A0vsBuNxrfk5w0K8jFxXbXFavwk0X7OgMRdIrBrWEpEe2
y8h5NSS5gdtpblXAlJ4k2jyuo1L4TSkj5I43YQWzllKa9jZpKeSypreVCl968CSCKe+zXzyFnQhz
E0f81Hw59Atghcxge68FBdeejrkX0XQR8YEBQ1PPYx2+28z4uFLcsNjJPjFass2kAWX/coISx9ju
GPwHOMFY3+3sDsL10slpRoA37Ds4JOjw/Uxbyt56+unNv0yvdfd2SQc2m/Uq/FUrhHLhdruYVBwz
O02OBIlGq18UWoCFoup7J6i9EMq8oIdEz3KlpLAYx2V1I6BLe1qx/sCu20dVt39PflGUSXNuWlk2
OzqFrpfKUPtwBqcedsl9bW8VVArh5Osc+nl+PaQZ+J/E68MvuDqcJaUkrdTNKUH+g9+R8fdXdB19
qff3e/bleNCQsXt6ZIoNEnJ87ekMtdwE2frga2LbCImj2NfmdEfERfPy+7eBYLvqMzrPX6zDehk6
rE5SQUD7K1M8LNuEkWUEK3MHoMDRpeB0W0GloJijqoKMOjpEq8C4DzfeKc69fSPSSViAgvSrlYT1
iChENonMK4IZAVs5WwcQNwtJHMcFzQjK6ADC+cKkpp1jI2jgsgGIlsNE+z2rIr77mpZkg68szDn4
OlXIlWT2PuXc61PL0R51O+pkesN39Xiyu90PvmXn+ZfjfDy0Dhc3ImndtUuua3IOVtDkJb/Cr118
TuZANwe3uPwllqIwiVZOc9TIrPRlEZ4RLqlVQLXrV/HHkydnX9BI5jjXpT81Tzc8er/YnK4FTPd8
1uk1qojAqQCLIHAWqsvaH/q+wABfwExh6thrQjhwPdfU5tvc4G8W6pzIGlcNA89vWUlfE+CY53K8
klCvBV6mseoPUAckbF5WuWiU+NKhMFhWVtL1nY1kZ+ETJGrc8uVs0XUxdjn25ND3TMXkieCKWNFo
S2f1DgfQUe6sKWd1PsGegxVsieXQGwYxjgd31XQNsyoPCh78MNIf0dD8IKp1iwjv2ktrqGO/yeJ6
wc9m2ANpISnJ0W24trAsIcLPPzgdSo4aD0uaHSOinHAIbihWWy5Vn8E7NjDZbsRgoiEUPWDsnxpa
MhjXLKHZPw/PS0OTLwnxZ86+wO0DcIbfQ5TU+hjESwtElQwSaBK6G1XbBSVtrExAfdG6cY6LnfGE
IhG0VqHa9CDHLFe1E6z7qPCdeIOiUI2eB4IqPz+whqzFahiW8AtLno1OPnb3fKWwdgUvFB1mfQx7
tqazRpMnTi4V0GjRqEg9NabgDqbZQ2/kZUuevJeRF14Q6FWwRvj+Ix3RNLZ0BSf/7GQ7my1u+ADK
EdJmsOM+KG8pgDBUpTWzQRDjZ456nmxQy0JF7M2JvLUucCDuJsG2jdyoNHB+BXsyXrWZSfkqeLU+
CT7gJ46pPdM3ow+03oHgl9Aki4iI5JqaoXntsvqQIu3eDRNGUDg9nBc6u0YPRvzTkcTVI1/llMQk
xQIjzn1UB2yKXz542NR9t6pLIF3FbOQ7R5S5PDWZEt1wHH7sNf3CuDjM8lOWxZxOJrq2BPNOHTpX
i1Vqrd7fgo27399aQe1oJjviDKDilKxXYUfEFsJpSglkkRuZB//CR4y13lLDzjwrSmZPpGfvc6xf
TQxjeNJGcdhJmHc8X6kaeWKVHPOoo2gMxIWz22Nxyc9w8S5TGZq6uyiXg3TVKrvZqwNVPRITDaX7
2WW8lt0JbJ5hjXk1+wpwPuLfaawtRnUnzgaBgQryM9jLg/FQBDtskWI1dm1QP4RmGLNtiX6lGBDm
Sdluus6zcHeNI+8u8CqlweARoMSr6hOyRhO+JALGj13DJg1Tk6vRDV+x8P0/WaePoxCyrAupxlJa
hv6XKW0WIMca8l0ep44mdzjPS6NyBLgtCnv3jCdqH104u0tEkCEizMWCo5CIJkm5rGwzC0RZENQA
gC2eldTQRii4pm3LImscEVfnJa9kXsGbbNzGV5Lbkwa7AWpUFZQCkLrhaTt17++rXX+izwFwy3Gk
WfZRRD67+06eN/QZ2U0ud4byrYKvsBk+/lahojhOLQTxZc/mrFwnah9NMwp/t9dAsks9Pw6VYrrs
D9eXnvfQL4/kzzPPMTk3DNg6noIig+t4DeYDWIMM5hoxbplNHlFJNubT25oKr/vQxP27bwd7/Ym6
FhB8gWYRzJ2jK2UmCl37PkQLw3c1geD3l1F/ZpZAg14bzaTToDrTkEPfqFbox15V84eM0f9xX/4h
oN4Hx22LzxwCr7h8LG4fjrcsZAMFAqe+HYnlrABugZKLMh1180c86cWGftLP3339uY0jWeEduUs2
97OQSual+4sb9kLRbSzmJBKswy56Jqj3Syqo6B2Y/TAqA+fwEyZ42DBAminbke4ecKMK3HeIKd9b
E6YDYoBCtPzKBkSFW0GS+0W5tl8LvhmNzhEK377F/d1QZLauh/GH4f4T4yWDzuvgfe6Vjun34s3M
GZpT+Z0M1owPhBxcEgrrqYbHLxxKHcDsn4+3fhC6M2xxabgnIt3CgcbCzaFFwzB0zvQZWXO3EICF
uO/gNM70dtuWwtULhjlYCBriWSPzHItl/Mc2/ssSMDrxlL9xhuWoo0XjplNTGLKCvlNcZxqCbv99
Y8F19V44E9HqtH/1kSd7VrDdqeamE0Oln/rAAsG/sy3tSD9PRU+L4uOUjOuMAN0VSEbgJgUqaJ7o
fGbUtvkwEYTfVrNEiJprtNP0zflx58ox0wqzI/8aUUSwtFwy/i5npeKcCx7NY8fT1QTxRu+aLsP+
bfGmnQnwv7QuwObdny+yDVKzpFNEgR6v+vzmoAdASTvghryVYH3SH93d0WPTb7ddM+/r7U4haXkJ
OzLuTvGMzemm/CkhbKcjjp1kAJGvSddPspIxp5FqKHvpvsXBCvAY392UR0Qn4xs40wJVZdgWINSY
BwqkensLssy/1c1xKafPy8WL8IrOcmKmGG2Dh0vhzbD/mtqLSnMENHoIsuwD2t3E7Zs2SmTLoGpU
mDO8T0p7BAcqVNcFYRPzhWJ4KueshcZX54EA6THk9vpDXlDRPY6OOVLuFJHPG7GQZiX5ok+XPdI/
5HPSHQ72iiKHewVpbwDzZjzTg81YJpFxHoVyq0xLgl3FUN4x6WDwmXqVesxCIqB/WmkV1USIxw7N
0XpRxVrzUX+9zIkcQBAoCX89+G7Sbn/VJJnpweY0TWdnUqUBa7YeGg3P5TU667NOUX2h3IYusqlC
5MCth2o5kZejO3xomMF/2tBDbSYCOOOoc49tVH5Gbk1uyILrQIirzMF3VnmIvEDeqKB6L+DqKEQ3
LcbBNR7IfitWJndSoqvf9Ng6dNuIrg5KwgbvSXhh9HejjBa/z99p4vaG1VN+S7f1zEhKa9UhdKwo
RMq93i2dPviKu2oHxe8hnTMTt+gRn+Px0X+ocZJJyzv+bqoXQON0hgrJjBU7mdRCwnuPADiI4bgz
uHN10FSCdk4YOnhnOhofZN8b+YP+R1xJ/IbENbyrMHQJ5UucLo+E6m+feKYrpFFsuIMBFTJMGdIV
8ebP6jFvMRAl+bv3onp0tm5reJw0gcFBvKlGMGa0+b6edsl8D8f2cJXrnB+epd0jJ5XTYqROKdJ4
SC+YRasjtlvHKzhGBstmdAg4mfP0SArSXad3+k6mGIdveMw1CQJysWkpyrN7uylWHpgaB+DxsSOh
Ml2RGF88VlRzGWidNpTmlrbu1oKqJ/FluJ5IN4xufg4j1jQ15v85e7TH9dP3rNmlZI/LW2c8kG4H
bI+ddgEIS9k7y+CXQI67LyGQ+cGGiSKstVq5Ry1I7Y8eVATVJkdFV7I4wbjt+VLvu0Etx+5cpGUD
nGZpQ9ecBvWSW7sP8/gfEj8pHZ/J+KSvGB6DL732WOaIb/Tb29LbU0J22PxxLnP4Y3NhGJCBwxNo
7tSRxh7dCQiJzggDZUefO+iTAYDPtzBoVPNZjc9VgmmjlqSuetFOfEhZ50m/A6M4Mfl5Nj00PzNv
dA+RUoYvvG/cHTxxz/U81IOrJpKvo0GP4y02SX/8RddqyqBi6nu9a2jziaGlWfHQZdu79L6N5FHD
WmUKJZkwmeA8DqqUz/DgcG8dmYkoclCZSRulvROn1n92f7+Y4/phJU94pG4q+SXNLY30kM55JtT8
lcWwdizI2Uyur50/lvpKDhcb6cDggJKWvEXjQDVsQg9XTtrK855wx5jT+hIgj6W38WyO21248fEW
LZxtSdhE5+gLZt7EnGQril+ey83om28mVYYPAB8xDgq162mTX2P+suVMq1OpnRPWui132aY0Zk/m
Jk6BM2LJZ74opVAqdyt3wrM5Bbmdpwj2dMVG0tObDy4Lg1k2FyibpT4wqTjAG81VVRHYHmvTHXsd
z9g/H9U24XyCuLYDX/3yyoWAmIgXY1WpzTCwcagJfJKHFnrSwRxc+vaX3O0viwfY/PTTj0CerhgC
JVqFBjFlaLhosPyRyRpWK/axchhNGOliOXQhEOC7TjMU4ayWe0UYw2X5x37d5P5D6KXpZ0tH+JGL
REaikzVIfVKOEY1a0u2M4km4q/kqRR8i9hoZRQqqCw/3v4wpM2wmcI/2cggAw+xd/Gbs/+cHxS2w
Z3nk+ADE04NRqM0l8uZN01NgaZHVWH/f4mkNNXkz4AZgJ5JnkDMgwbk+W8xZ8TEm+uD6JlZRLuwc
xDirAJAc9pfjR2wOjt+gsDI5zGGp/JWdAOFEam9ya9rpdTZ/MFvQui3TIu0YwbvET/sZ7R/ZG3lt
UrtbccQpQk7zE7ttkKjdqvK/FiEaX8oSKj0f3E+h+nbI/qZIRRl786yAU2RPgV/V0RQgYSG/BUeM
x1kTwoLYogqRrlV0gVhoaCb7S0l13sBUF6TAvpf++SeEQyY4Ncqef1QCqQzP/90oUriXalcLeV4J
mSGt1K8SVuWA8GHhhyI23moLygcP3MS+RKbFw33MW3oKKEIdTCjiSnemQh8urVYoqvxesMro5Zli
ssQ1DbjBU0niEDGM9w15/bVn0J7jwPCyr39VwOdwTXgtghafm7+FWJ+uI4v6WT+G6l2Jv7BkED9L
Y2RKdx/6SrQAlWrbjY4TnhYfS7p4wAU+XZHV2DO0PDRvgUbsjAEzO5dihL0ZJr0i9hwcZ9WXw5f0
JprBvSkImsmukWdezEcpDYOatTvOzMDsrvQ8w89/5iuk2WGQ4RxiNpcIpht9fwKw7fBqqkVD4Y1n
CX0fbD5xl4qIm72OAKxHOOzXrnbTD9iIbIi/mxTszaSwWArRn2Ub/ex2Hk4wPaAmyv9OEkTOujR3
fyVgYPpap1Qxk5VvOjc/1I2NPlIjpq2YmzZLbdKiifYLRO9CW0E41reAcb6L2CGHeqbcd/PpSEVd
AiOZdPmw1MRt9iy/vfhgNFooUoWPT9mk1rz1FVY7Nff/42BxFHHGRHJD1dLg6l4jhtsVJUQMMi+C
qfqu6XhiGXRZUkDPNhj6iMpKO/DBk6EBzsXfEM5PdqERP5imjXUkzDaiUoB++tXJ9rl8yV/pxwXx
kCiMuOv2pwducpr9viIDsfzjOIimpg4W6BOdRTwkNsEh0dlskbzLZb7aD/P1frD7wCHTsQFRFadu
RhdG3lzTM0HaXxpSuTyrlo4HptWEUmUXcV5DGZQmez5/oo3S5v+11YA/7S2S8yg0lLxOmP+ZeEG6
dGCGA7dTfoRw09fgSqn1rh4Dwu8LlqQ/N5tbQDuHeNqzqBtF5nNIq1PvkL9uD8XgqDRBgi2h1M/B
Kg5qlHHi6iiOnBLnb1adew6H1NT8O5K9dKG7zif23HG8SAUa+M9e8CLabIgyzKamrIbxjhlYJ5YH
4D/aH7PPkT5niwUVOumH2eu16F86gllcd2+Jx2jswaFTH3Ogz8gvlTKbGWJPbCthBulD4dDYOoy2
IiLg2GdZnz181LsnxRleJ4AFZD6h6GHCxhsCIq+67f0JyEgmkW1aLqF06dzmZnx9zE/SdJnLZANN
ahDL7OYQs6m73ny5SIMnCSgAh8EB2+xI9DTAo27FpIzqnbSFU5tfVFTWlskzRNCUZ4zYkC5jX8Qk
hZtge93Oq/COFfI/sAXgENu76xaIHFCv9mlDdC9Tx0aFRQ0cdLni7SN4NznovxIN7lsNrdrrOPKX
cLFU9Sl7lAd/+UwDdBg3vfFEN/MyZs1YcDrfPJfUPsRv7SZrt1BEsRQMJGdvsN/EfAoTbEw2yRuS
s8OTewAsHNl2IffpixHfjekhZt943RNIjIt6mRxrBaFNIduuG+ySBm1ALujbPHqFmTPK7iNRuH+6
cEVNHTrV0CoSfBflTCZjIHF2nWm4IoJXNA1WoCVLCHn/F7B1udi8IuTg1Ly38xNhUMhxA8oZrLIP
oPvbd1cOEIyD4m2I07VaUy+t/iU1qWop5eynKWWO591mPHtUNznrrfd5/1loLWvIgZVijnTBDvjC
1gthRabMTBBrUP41zrd3hoOxTgtAj1F9BDK5+bS9FDYH6iEcMzwB6sB2TCGhyL+oqn2gLWzfXZb4
LyFvK+zTMf4OMwEOsZ28S6iA5SxxMDJr4yCLjuM+u0+MnLro5xlyzUueFqpWQifUV4aBisfPBqCZ
DZMBn8s8jWxCs3KnSQun7I+k57n4csQwQmetHBJXDjPWI8+yEDut7vXxfIMEZc1UMmDmz0tGUwNP
sQCex+TNEWsoekzzktxlDHFPuHZe4n8ZlSrdLhuNlX9zPE8Pr3QQpLQ1tvvBdMa98mfk4ErIOdbL
j769sg+Gvaq5nTaMutFDm1YzYkKtSjIchY0B4jV+G217aTb68kBU709mqGNHrES9xx8PSqSTgtsy
pp1LgkjJk2GA0iWfunWlYulaLfwNrxE5Hrlrx5TlIfyY05z3C0XnM9L6+GagMzzlaQUdNWr0x7li
GfK5s9/L+/sfiuJRHQeFWP+QeK68SLf1RWN3+d7ej+GEuS6L88gI/CFaN3tPvhsqRNE+wJ5O71me
sNfPUs1Cbh2HtxMgrF7QwLd++LrYemcnRx/QqCfXgSRVXx6yS+jjAr58dg6essAc/6G9LxJbdIAZ
D/aKlYgBY5pCIkF59ZTDIfKGVQKvdnBr4y+/UPVM9lHVPpB9noVz4RIxvkJSHwFxoFTFDj/p5IG4
ZMlDuwOqA9XFJ4z9POm4a1bD3lHkED9VGapAryL623cXs2AeySIMFJ3RQa+VUb0Px2GtZBX4snXx
Qp5QjtZXVyPZ0ZS39ZYHiA134IM7UD8VK91sqYpcbUwjnp1tTM3hH47xR4wcMoLQ/wpmmhCj+/i8
70yGHRLN31+QgC+mzXNX3P3gcsursgcPAptyzP5h2BwCpMUCUZdW/YnfUGqiLNx7fG/JC2ZbYc3K
RcPhFH3bh3wvWOG+B/6/w19l9ZYhjEJmAx0MHIqojTvsT10e//9w3+nbzfHHCLJTplcp5NEHggiD
C7pqVUimCQNby6jdPGoufvssFSD2B8hW9jOArdgn3/ggAsqMqjBhbryHJbb1CxkqqcaU/u9XI8x+
l9WehtFXFQwoB9k0BSkDGJA+RCYgqSkJ+ZL/K6aUdcxXwdqnAfcpaajJnvpXJbyzZa4/NUSpkSpB
xXZOguQ0UhB723GNbxIJ1hxBS44tf3wErTSPsOe2zCtfksrHl3G/DtX1ctmMjEjJvXwjsVtrjPJ9
sN9ucMfiYOLnVIr287ykcSTAEe92jjiOWL7JjGFYh1KcfCF0eBL5k02XPJODRar8BwICAmkqdhYE
M+glZ76Wky2ItD7bWQKxmITZfexlbRPAcTTVQLFAQ9cC6ewjJswrGYhO+nHkdU0IAQojCh5gcOSG
6yoJ7an70mZJaLuavO2Wy7M21j12NHCYvvs87duBROGha4xgfQNXxQhsylga8wsAI4sQfvkxUj6s
betW+SF03V35h2aUXefRAdkmReeOiJipK2Ml6wWY+dL0yj+BquU6X/l/74h30oALJzsJ8c4IQWaD
6NGBCkdf3VSye+DvM5ZWSdM6DtxIVj5EWaF+qRcZ1xcL/mAr9zmEZ8s08Gh24wMlp+ZDyjTprAA2
m1xk/ccHKo4p/h+ndbq3RE0L/O4IG1HyQrB/5e9U1AaUCzue8VV9tUYftVMJdNriSmJjIeY7KJIS
S7/b+PWIhG28youAUA+2Abj1lNsLKMHhbEbTVlkAt3fiK3Wnwp0l4IniVeFmwA+RfMIruZxrL2jJ
obakEN9o5t96X5B8SIZAEcns3xNsr9Fqxc37Nm6DjPoyjUmf7YTEAO0BaHPt8J13FT4Kfn7eHaIR
7sdYs1DULMmsSj1QfE61lCioIIYGw5HjOA9TDALOZE1ISwRF2uJoiJdoAAl1T2ayeOaKc74UaTet
Z7lbe8tOz4hkp+PJBt6UV8dxEB+wmqgliWIdgTr68lSgRA5XseyH8L3Ly+89aQ6mssw8Ylza55Fx
exjeZWgq+wxsLUR9ucW1NSLU0h0RNMvJcnLLkhAEjbDFYPAM8rr5XFC6kmewQkKAB3u5bwI82oiB
g/uOs6JS2CicYEjzW2disYuIX0vn6lAgBT6vNm/9to/9mxm1P4NhbwO/52FYm6ZNWDiWbmdcee9k
Wxhka1KgKh13mXL/KT8f+iA2X1oeXFUF9xcdzruW86X4txjNRsVe/sFIuMphotR/36RW5R7ihiWl
5zMNLrtUQbeipZnQHJsgHY3ZtDY3QoJBlJ1Ma9cqwNSpNpTCRTaqoJKbihfCDr0PQkYVLjwD9Khq
Xga3RdmU9tDi0b+6qsXfqQNhCzNBycoZDy9oMfaEyizmPyeKQzjprBwE8RBCQ6dUW4PqNcqgA3Gu
/QiJie3bZYqyxnNkNr/DEk04ENfdYzrUJdt8xM1mqofpkYqTqMfoXY/Lg2/ZFYRkpG+L4DnI1D67
gOaxnDTI9Q3+/XC8m3cWC+BOnzoMjOuhi3HfPkZU9p9DP/D4Er6DLGRSHYsCNQOh6d84j2y4uXvb
jUwgbcV7weGybUJX/oSZ5t3uEHi7/pGoX/O3O1ajrqB/IqYEN9jO1b6WuQevZk1auuSGTjJIthku
uCE2If579tctDMeIxZQxqzC6E0wp2e719cXkImMWSSmOzHBm504YVH8KHARBjLLidY2JoCRSBsED
KRpunxspHvlVf7pVKGjYxOihMK4cf2ogm9rekS0F/s419dhMt8N6hAGa6/A4JPhudGs97FepCame
KPFrPVgpo2vUO5UgJHB3X1u+UPwfLqbPDcoZGMn6cgzYp3TOV4Ck3eOsLvFGEE7F96YOaC1DafEh
p/BPWth029nVLrSPoK1ca7cBk9fwWEkwEnOZyq8bX+CBjHMNV1dUN1y9G1QHQk9I/Z4MedQ/7qiN
mkSR+ARTyE4HMsVyY7GLc8Ze6a7jgI1HudtQP5CSnKoLzdmw2Yn+PuPUFPUkyF59TMYoq5PCVwbN
IbPurnPokNzhvzhjbl3AhF58SH0IwNWYxftDwgxAuOnzCassddV0O5tbVnMzxTiPWh6JlxhVeE3L
Ko2h1GfVeK64Y4dNvJWKGtszd87/F+xn/lbsFv1Qp21cLkJRNarQxnfjF5QvUCL9gJzTmw3jcJ9x
S3BKKpBT5Onr5dktK2NnyTxqObo30IMVbs+zvOfdMrcv2Jp8CBoy9teNT048dSDXfcyB8/3Bo2UY
FjrOxx9w0nUNOxutBW+sNNNo1hI90CTDSVkYAskhsMsBau9RhZHaC6Os4SQuUvM9XG1XVmfg8Tgi
vrIRd42BAwxV159T0atkPsOtdOn4PQhxkDOQqKb1gry0WK6JnuHX2LaWxUY5lK/0G+UApthoCj/Z
zJ93X/NqicTA6raCGvPSgtJMIrka93rYi0KNO59x104gHFf9cKZd5LCS+84gxsJ64P863KdRH4lo
HjgaW7Ics2ZXu9JKbnyHhavvSThcU63G40qYlvnUd7giuX3ZwrBexG7JY4PIBNEsv9CHUpPrTJg7
iYFzwqKz/zbMDZXbK7IxlbMY1j6fYwN/dT565Vs4vB8kbSJKVfnvUzccsH7tIXMPulj9Uczj0U29
gTtFrGLTh9IA0rtvw80rvs394i6+ta9xQL3mjG/gmscEWRz9gV3hHiV2+BTorWb9E3EZZYEzIgC3
+DvF2BNJP/B1tmHlKkgiEIKI4ImLYgkHVmiQkhv54aN4UR/GLPwCspRGSv1RXqRICg2QyZEueri3
pz1/RcZ3GyQEBqxqK4myeDGcYNEhNHdDkdhhjf613zHFrqgfZBg5ozO7ceJlFGJn+ybUn9B4MwnE
p0SHfKQLva0uyb2q0pqmOoLq/B0hwcdjGp54m+VLN2yOZ+PFDEmi0xZPRm1k3DQQgnD7yySUbVWL
fRYGSn5jr+jSJpr7wnW6mJzDcZze0UhW7HpbmLlBK11CiD77Zn7B2/m6MxDxL+jnmUqHwo08JZYK
Z38hy9e4KxYCHb/cPy/Gjdin3mXuD33m/Zu6Xkfh4XUTyx36MO17yqTwm1+Io7EqQt2J46sf4KtC
2xnSmJgi2G28uHV7KV54qzYyKpfIpstfQRvA18KgGfY0JQa6csfuRKAJCPzAfTMGzrUJpeHcVgyc
0IgMy4h6gT8241bHpS3A5prBl99srLiBhJpP09pFE1R5eG0nboDoxOoRISql9yaBh68tdVQA3xf9
OAjFVCb/uFfFuovRDZGfZIytYQaW0tPadfK8qdy8SS5tsFmv+HRC0O9GF5aDUvZTWHLzxAtz6GNA
/Q3ghpt8iy65xIA1/MKLcrd4XlfCxxDTY2EVDO0Ro0EHXQetGQi5kB8ka6tNOvLhyYHjTeDOCpkO
mUJRMvYeUrTyejrN2CDvBy6clqBcQYlLOo454CuphxHwgXiUe3Jsj4qhdBqN0ei6xBjoFAY0SkMS
bKUuJ/NFysPEvpGcMpHXkqVeQS2/+HYXAOrr9U0EIaNskZWIt0vG2inM88Y2oCZmOAHCMkkbn5Px
O+fQ0nmIaICmUO5q3Wv0mXE+TZ+aErMlB+3A+1MXJgn7T16q/RQMtj3o/jHc4CeBIBu9odtu+owq
jBDxxNS2bMc8iXO/wXpJl0PxkQY0MaKf5xO7N32Hr8LYdfOqdn0XYJXVbo86w+T00TbE3LCqPGNd
C8on2MVo0gONKA/sU4kST1TFtp2D01R3169edR65ucMflbyW4N0KfnSMMH0vQ06QCkxsKGysGTtY
S8VkBE+OAxCNGeu3MQ2I9zvhqzGT1qKyFTvn1NrWD9ZYmfsj5veO7Y/75UHXk/3wRH6sAFNVhGcp
6FpgCNaQBKD5L+F0AC8I7hswz1W/cE53/llFTJGGdA7fZlSgLVba/9tntndQZDiq74z8t2Tx4vp+
x16UOSB0Opp0O5Q3XKaZfZZWRz5wUxp4beeXy8Om1L4NDSEnvFbsoPeXices/aB/NORtrwqjTPPc
V0yQeQkAXVKzQVXqsd5tncV7Rbn1Fo38GKE22Pf6p7MNgXA0iWT1Kobg/MzGKSFudg6IxLasbX/f
FR2GOGn6wxnGx4vvrGRJ9FzgT1rBJ0Hd1oBS/4g4cN5nc60edN7nt0Sc5M86Jl3GKtOUUwuhkxk9
CXZhsfQYFrMGRkCJpgOEPvkogmRwoenuYOj2vLE8qHvks3nAFD/jt9uSrapj0ObqrFgYYsANy3AD
BjLN2U+34COjMVIrMsn2kS/ibLfhyZMejZFBMBJLQtHS4pvTGuz1I4x3OlsukzNnal6tgcGlTgBI
xshHoa9PMM8qFa+aGWZ8DP5Te2tpmLBn/7pMvTDUJxigdK5g5MNvvmTjmDDs68oerVoK/0Qj9lXQ
e3LoSP884xKllZsDQsTXi3H3wBcbd8M6KYf9G60stGia5w+878U3gOltJGt07N2L3k+qhlXEZ58e
re6+T/gzoSysD2VBODDN1viE4T8+wo3jkWUWSM+YBqjSUs9Dyhs28l+NKRTOx6A6nFs+0HWwyhJP
4NEENIcfJXQV8uvRtkQbQ5squVzrDmzoDfMQjY9u1+L8he+g02R6l/A83KKecqClVOPSa/PWcTke
T6gazoaCNCFqzqFmLdJc/ZSNUmJc6wXjy+Ophaa9PamrggdDwfB0ML3LVbZbA5xtEnbhny1U5Qwf
nDPVaxzrTbfz4sk6pYTOr+n3zliIWoNRdM/5y+unPP/K7KIC95RRfSknznJsWhpvMi5qSJVPVupc
qxdbJtiZhmCfLH6WmUcHEZ4aYzYw4Wju2nM+4mvpBrPZOr3PQL6tHlEs8VqIGWcypH/fU9Ybnwxj
DYgNFzeBDoaxLcx5kMP2E2g8fUB/UTcx8PRV5Zc4JU5ICszwx2pG53dj2YWC+Hq7zQ5Ig4RC/po/
iwm0jtfAvxhG/orzeWbO4rYXaTYuTA2HonA7IeNH28PCFRKSElZDMarsgPkOk27GNR7ybXNoTZhE
CBcq8R9L9TCe/S7iFg7DovFzSmkPaQ4gORC0o2YsJN32OOAV1w+3jePdHQjFy4GaIET8adqtolVN
vb0YiwatZC6RTDelw4+A7L9d28qK/iSL4qtN5lfajPtW0oFiBuNl1HVp4Yt8ST03iAvZRtfQIxry
pFIZsd+oNsQDkJcDzaiqc4UyEo+VlNNtcIvftzKUWjXUKWDxB3mp+8aaV3uFrwG4AnU7xeVcKaCY
y+9puahTLcGifKcikHwOv3p2LN6QP+J4m3MpLODjUgE914toMG+HfOtLVMVrQecYg5PmPS34Wvrj
nUu96qDV7AaFRHqSAI++4db/n/siod0uWwQkL61HR31CxOGc4Q6/AbfKWF7UlTGAdMcBF/tpy6/A
NfEfxAfkW9wW/5w/n62p5S2EnX8j7tUhKLonyvICn8qhsOhmLBxbJB58aC1t8xv9bT30tDryr/mt
fejoZLcTtdWE+RaQT+14ozjDecVHEt/OYXRc4lGzCsJferBDZv0bhT+rh6YLW1G9FxRIkY4HCzww
NHMiASK809FX+gv6+ippGfSLI4XWqVQ54cHr32fILv+vZj3O/gOxCrFzh4KSCirCKfY9nTN0e8v3
duNAcQn4YencKIvLLtjf0MAnI/ljyuNserBd8m2fov+1CLb09nMNHOKKEM4IzWf7BloulYk4xgE0
Wh76KiAjCu4YATpC+cLJ1lGxBwzc69qbh+YQtg7uL8Tk+mH9aj6EgmEnHlY0kRygn0nezAQw9WGS
XlZEL39rkaddYvGnQON2hwgohapCM4/T+BWhdB2iyi42wEWzwMM1PJ8dEWsmTp5gkw4QLYf1H5Xl
tr6OBxs4hy4mMg0a391TwIedMjnXNwd4ANpfUx0bCyJ2P7bRuPwOv3lwUjr3Yn+v6pArr6cDSibG
sqa6WuxuRphSvo0HvqetKveCBEIjPHf3v90NRwD+eUXpSF7hH2qg11e4veqXHtWMvDALED8/SqZs
RZWH2010vusVv45StnZKqm2ZzfcQY4YURvIQQQSJz6kUGx8xswll3VigcsFfmqRFsfhduQwOXcyE
ZOtzgdfunE/0GJx2PxzV+31VNSKSxpxmj97eAN5q5pjKfuWiOs7Dpzxxlj2v6x8d1tN1s6on3iWN
sve8Gidy8ylYQryaeSGdOPvygKTcbSmNQroiNXUZOoZqAcotus9D7z555hvMX/3bECP6GpSiXjKR
vdS6c7hEprqHq1HbUfGlJhi+//4Z/3Y+eTLZ+HxZnWzxdu1Amgd+z6g9iPf+97vWUcrM/1mY/do3
40llAIEUBMDuPQABH/9nNXqc2QIrZDj/m08fqvwNE/hrN/nrjq5i1ut78N895rNZUBcAEj2t1hzp
Kc4HsZS8vWK0WeWlyrfarETR9zAmRW6do1rmMwk9rXPRmwM7W6eTorI1fA6CTYC5zmWhdJ/VaNcH
v1wxegW10DP7mrmePbaLdjxgbt8F5ZpzuGH5RB44bBPH7WcCmtkSb5tdbKSpxzZqfj3G1ynYZgFM
K+o6ElTiYC0nq7IGytSRGCJEP2wbvSXiZe+XwnzIQ9U6nb5x0k1AnPAzznUn0qqDjck4/ZQd0u3G
sfBTIk+94OwMTy4uK7qhS0U8TA27i24htcGNczi1H4LOn8wt16c8IwrjeGSMaS25W5WAXYCGs+As
G8/lGtKRJyo9Z5GxNP8JxRl/D0zWODuh5WVsKEqWR/BtToGVmVsv4LpJ0nqyd3YyyOM3tiCUTIDs
nVMGCv7a3w4wtKAXmw1m5JmjL81MPrabRZsfhRDaP1rdJhQaegQy3+1U7wik7ox6OVB8GNX7lGFU
Gobrl6RRnxtanhqDEasiCxUmJ06zlXIUNiZYht2kmX8V+QDrwo4oJk1mYe3Wt1sxLSq3d+P6UpLN
9spwtTTAJgxhwcUk+xtFLg2SA5idKmvTM2hU5P5XR7ObfjgCq7Ne7HSbJFxQe6wGlsBBKjavzr7z
dmDX7wW07xYPCLNR+4PM36rM2vIBUiyzYmADJgXc/I3+Ori6IxVBmUu6tn1z+02w4H23viITZ7G6
SS0Z2uhpppfP7dRz0uV8WyAuN1716/b8LMM1jGgXSSJkVLJYdg86czLdPjLpZTExP8nyjDlXPsJt
U9OWjG4A1REyj6sNogxKp9ypcCZGKbdC0VUN1FfJ+P/io9QHn5BjniUzsH/d0ZehKbfYDGOKrL5v
Vr8eipjGFmduMnSbI8iTMv3Zar/13AXJb4ouKDnm2Fho1i5XSvHaBpg/vOsWydmA3/jAZ+/bsN1Q
4u9Mz9Ka+TWtekc4/LRJqdOjlaHSgwhRuS9pvnnguJBR++yggmRRBG6Dsyi528MOAC7i2TsEezVj
Ic8QEbyXRot/XkKdYYNJj+3QVFFAaOmk5DrOS6Cvyw5/87VNx6tKvC8nVXhVeAlSCKIMspF/3aes
hWdmHYrlW/lmGeyJQ6OaSuU3BhvAuM/ixabgD1Pb+8n9tMhssez7aCndkDvKdrkDofj2+xbF04ux
rCSEmb4RV0eicW7dmH7Gkt3wU6kaQfDHFHUhoclWWkgG7ldD/MeaQHmruQC4gnNlN0nIYme8fml9
IPOcjlP8+uB+8Eyb8Ys5wDkznKMGm7TQ2g8MbGSeIpfo/mWZ/iLNrRqMLRvc6Yz4DPs6SlPwaMlq
nzhbD2IbV5f5dtWQr0/KaJVhQxtdMTgxGcLf624rXbl2Ie3JFaPpMz8AxJ/PDSj0HskVlUr4kCiK
pdEbeCq4pj558Jfy/2Av0ieDO7TYvRLhBimSkOLQHTSJYbKixhmRrXxxCspdmYobzPmSc8/tMdQo
q8wSfTCaQht18S+2uLz0bxXjQt6xs9cs9X0hgNiniONXVixO8q8HSbhaTE1zHxkIkm0q016nOGn0
Mx9iAF08ahkkgH8KxXM9lFpOX8CXiZ0fWgQ1stK0MODiVI9XNKlcRD8clBpMSsysqrsTl/dEahqn
4ciojs9cF8jso8pwfkHglYWU23SbFeVB9eRyukmH2SoUzxXhHXvcrXtcg7lfJeg6cxdCXW4BtAUD
YGLDc+NwdQ90Tx/irAsAhfIjAquZ1Hbk7JbteJxTIuPcvbb4fT8dvA23h4bYMoB66f0V5ZODt96y
CXZ8v4QozZDKxpnxkXif5X4BSh7D1jr+udKeYYni7wGPXJLx9zRHDRCZwB/HRnOXCprf1y9LjWlE
q4bUrOWg9nU9mMCWeaHWTQv5smZYQ0a8FJHS2Q/S5CnPmBw8Kq421gI38KZ78Ng0Vyr4sSCB5Geq
6ogwNW3lMepdismkaQFUUpsNMOvQkfq3tvfK5cObl2cIk3K1q4K+NdRfcqIcFGm/I0mzLMrABpes
7oT+fRZV/8Nk2X6w/0lU0arKAwWDvBsxaGrPydBgXNzQ7QEqR35KI2Lw23BcFGWUJVSZBQRg+9Up
JWa+PWvUOf7aVo0RCAq4xiI18LmQzUEYsX19PHH/dpRdzslhWptpW7Lc3sv6UciibT2/6v8/+lr+
eZ911CJ7SUWnqEK8evsJv0gf1R4Uy1/bX+hOGyXdor7qdkt7fUjfbQ9BFl3jcdjF41gcVnpVcGsW
RXWReONXeCdNgvt1qFVbedMl/+SCaLlJyquphji5ed+9Ubz9NXE5Xws5oJzmSlenazuxrAGBy7+C
+fpjcICNIDRvjzDIZ8XeQVHZ7w72wI962nEAPeKHIvUwv0W6wMHkTcYecHuV18+H6VCIWwKK8Uvm
EjWZbwcl9/bSecl/0bq2hdp71pN07EGujXjmf+R5UeGvScw9vjOJ5y00UfBJPOWPdncelLaWRu72
FUyoY80ZftfNh1wkU+zze0c64EIqGn778CVPfdC2iqAnm9imdDEO70mfjeMillLLdBsNTtCSU7F2
E29hDtS6aLpJ6TkNC3876wl2+zykFfwiBhLOtmeZ7q3LLZyobcTje4x9row2CBZKa2wtdzkPBmZT
9hVf1UZplpoCJmRYZG9oyd+ozcQSr8yFO09aLpVBv18/mbKOPZJ1tbM0KtMQ91vgJ74H89lYhbAE
yCCvGmC1dGusRuBmbTA5toXNEII/ETnYvEfdz1fWOwxndoX6Y+7BnKOMywXeFsHO3D5DsMS/4Po+
62yhGssgO14TBhWyJ3N7FzEL0vANENBm0Vcu6DHh0GEmy1UQj6WUyivzcvFnhEQEepz5LhFmPjE2
O7jPOo1DFwEa6/amPDDOX8c4QC0rewJ7ksSADzhhmYXnS9Q3JySFyB8HJv0+xlJ7U/ndm+lhTq0o
xuKkZc4o+O6ULPvoQKCx90Dn2YFfhcBuGaVkLQ1m3F1C4pmBAmd8fCtt6UwgCEJ/zqb4SDNJ9zxP
9MR/0g5QBR9dP7EklCdu+xP8SU2eJ5GZ207FaMaaYMDlr3dpyo0iW0zNeEm6RHVmuulUUpqRBIcB
DOmW/9Fu0mwpaOy2g+cKWy+hX7A1CRFg6yQFzYtjugpKpmtjlVlnsAYj3z9n4MynBy7ufnvyC2E+
TLZU3s/C2x28pY5yWkLFvOEVW9nGDLwLLGObzFx7pI7QsHr30Midxw4Xw1tBHEFJ8lTAMritrOpD
gML3FLbP1gQUE8dTiuvs3vTUUXt6JyhtUIz1liYuj9veYBwjw6kXY8DtsuW1kRCJDn/PNYfRaEOV
2uPtO5AFGahbA7balE+EF9kv8bl2MvVama/yV6JEnV/OZ2wKMkXgZwV0Pri5JJZZwwieBM/GP3Dt
0LZ8ARxbWW31X1m/Zw3bPjuIxQnn4HlAtGyCHqZL3RpaafxhQHMtHdSG9NlfSdM9vzJVEvWF5CIe
GoiuTfKiOwPLxlpluN2t9ilSKYyP0haMgd6gAlpsHgoNlrGmyvjJt2C/NdMsJ1XC9lGuoEj6+zvu
3Xht9LXpRbohHyz6xMCgG20UKFlrtfAMij00Opve0vKRCFp0n+n0oWFCgsXK6H8AYaDXC6sPK/3n
tlR1f0zwFVz/8v73K1Q84DU4//ArqNJ0v7djx4tyGnpNk5JHy7RuAn/kvel6bni+wDfQ5khy540B
h2Uhtkm5xiqAVUF+yEauRcQCRp7zSEscd6YzoSjZF1jtgCbWtuuZiR0T+H9i8+7glV951VK52tmN
fnTY9smnfP/u6C0x9oxgrEvvZGyxNjKl+wJxvQTKRcECdjVXiD4dWagx8Sqv9UVKubaoNisU9E4T
Epu7t+7qVHOku+Nok+W6r98LpgrNW82ukRsOTJ9NSiwasTF6uB0IYqNL/TMNEhZ88MacF7pFYQ4A
sW4PNlz+B1GKExPM+nbvTA8sGfpBab5KfFrpTa6XhdEjvs88HydJuDXJtnJVrCV3dSkqKDZCCo+T
KSo93Ucv6E1af0/Ei6RE16z9NcSk4wMMfRTYT5YSjfigz6r0LACu26hatgh+pw8/xrFvhBNBClrm
+l09kEW32G7s1TSLlMRarZfOXjYxIjDfVYp3GIE5PkCNl+idjMYHuzeerkPWILEKbcVDdcjUx5yU
qnh4Ik79O7VIPRSDveGvBrEeNjow3rcqXkdD2cNXGcG6TbZEBnmOXfkehuZVQWB1RnhjsZTG16WJ
pv7FCk95m0JZ7K3sGYrkyEnaUT366d5Q3K3ofb5vHkKp8aLn0SG/pnj7jMaCtAKPBNY9QylsYQfV
OTq1TOYWlbeeET5m3pwwRlTfF4VGmLxuLJe2D1qo4PTVnSavrENl65I+CX+c34YvzY7CajFXSTpo
IFy2hfMd9IrQf6xFobFNgLxC3nZajeWgQ5/2NP8/AC2u4MHaXSB5F4+JozUhlRx9o7QuwhksTULx
1f1y8UG5gIkN5ofCzoed/SSUbpwz06g/qvEb7B2DklyVRtj8Jy+0j1bKBNkxIpan+xiZ1CtXDiNi
/3ux+RUyGR9pEdrBMb+nXhoXag37AiNfAo91E5dQW2iRVc5kX/be0vzB0wUGRS/SGvqy1hl/TpZw
mUJpPvxg+q19IqlhT/zmjt5hSiks5mlNATQye4iG8TjKHNPldaGBFztEJcwH+ctg8ag0HS3mm+4U
5n0suP0uX1Iyueo6ugaBKoZU2bc8dIYXQgZzS3rJlLFCWzMmze/XMxrN+/ShF4piU2FYe++vYOK2
IGK0H0hUCs9x4pLW/tLa8+8ALC9wM2/CGpRXwxUjAAYUsiR/St0fhTGo/QDJoUGKtEvTrEXPQIr4
qcKMz+g0LFJg4ORWNKlZ+y3eFyNv5sGA/3+EbDIKGFINqpd/roKzpymV+/nRDkcV6G8gmocIifDA
tKz1Jq8tjyj83uBO5xUu+kzXE9YxW6JcVzmZZeLUqLFuu9eYxlmJToTYpZkv6qN04aIhiEiooHIo
3zYHthNb4e1CA5noOvK/ooiO8w7BaDkkxxEKQTyG9WymU436Uyk0T79pBlZ1E2LJmVKUcyBVsFUQ
FQm7nhAuQchuOIDsqb6Z5pqHr8yZIFVEEDACIMa75xl8mvrRHEp8WB2thx/4TIYcQ+uo7erAqjWK
P2hL9lKqb5HeA0U0LkcH/E2inElkT/XCOleNZdhXlvj0f19iIKPFrm0+n8RlAbA8PpSU/QSV10nT
S6DOP9VEoW2bbRpWd4xjc6URO3y+mG5+M3M3Y8Iqp/o4DP9qcA/vBdJteJzwD9oig/dyN3a7cWdy
A/tNBSHaGpbatJ8tNcxkeVOLlZLNn8fObHRH8UeQeHjUQQWTB32PygnFSkT8rMpdRTV6mJo8ceEf
xCKu3MFfgx+ggIOq7+qE7QpHl2Vj5kE9wi9z7shznhKz2a3sheD9vDrJdZL0JP8gYaK/wWBkrBSM
g5qhGhBHezHNRB4uSFrmF7sV7Sga37mADuB2zw77xMZ8cAXlPymY5KGL3tCJ99fU2xUbIyVSUr/K
+Ly+rjjhVstBIESC4AgdQQ6HF9tuExnKpH7qqx9OF9GErEMPh+DbKRlDk6kUNzewPnLTVaCaTge9
MG7AZGdXxe3MoudBCkaQ1eYkEGLsYY1ORNUSqb7NxYrmrUFJlQE5nr3E7ka7kUU5rKyUt2DZIDc7
UqSUh2MYn3J++X06l/R+Ip41x2qh0cWx1s642f0gV9LWuGvprb2Ctv+idZba/Q8CdDheDU+CFToX
5p1Rap78US/hkdB8kYbpFEVtBQ68F42MR6MEjVvHu0Lpd+vfBpuWFWB17bAqWBgcYWHiML4PjwAt
g3zhAUQ/LchmQuJSHCd8/9EowJVf/Bpqfg2+nxfay4Htj4PrnmluyLiBvJeHv6YiRRdAn4pPprAI
0rF4HPasqp/7wGdnfqvSIPSxkGkZpxsXvSrZg5K+lMcOvHsonN8AeCAp0nI2VomO90YCZcZcFlMb
m4ePueJrrBU8jqbx4YmxiJwsnjXxndn4cdRaqCgsGIAKq6yuhgEqjE7QizcZ/nHV1v+D7EUFZJ8b
L//tYJwNwOKL0K7MrhLF43MwE5SWPbk5yFkV2JP9GBcm6lwCwZgJKKa2eSECSrcMd6yus6t1t1ie
FcfZvPOIJ80u+ggHoGSBEuCTqeZX2ijgt8Ii7glODg6ZpWMOzLYsG/hIzxDjIiSiPj8k1cQSDSXS
ia0nwpz/rjRLgp2cPLPh6oy/IJ047I5FjDXSaEwYb63N/m4k3KSN5WF5wp4fhZS7Botyd6ZKO1PA
AyETAF+ZF7KmW2Vwo0gR1hRbmhfU1QiBhwKYb5w3Si/O7F5/GAFzh0WEn/JQwqhw5P8EJdMo3S2u
CGSRmBkfNRJi3Qjq8qCEc0nETWu0rPQ5U2PppEb7xm6NQ8mxORYOH7Z2ggpFHKcZJ8rYR5cvaBW7
MKYjkmCuuIv+l1fb+sb+pq+aOCVf+r3cfFBbtJswwK+3QY+qP6TtwQFt8v7y7RxyvnwfcrIW41au
1HvXNJATVQDMl7LMnLB+BSuqPGCQ8hkFSPmd1V6OpFmyzQORrH9QxIhgKoKuE9icJZ5AAmm10M3G
hFPuM72F1Ei9Lz9d6iAFRWmj17s9piVrKqO9Lms4MlyIPVwfEVyE82N6sc8bgld5/lszEYJrwtEv
162B5/qNqVf7LGkNqY7DWqoXgOHPAKQeiDXnAQ2oNwvF7cHlKFqId5bJbiKiNiKWPJup5341Xgc6
xnbkjDIpfPMgQVOpZxdjFytDgR17YMAZe0ZALkXt2ukFFwi1knABi0zjmJTVnUslzKU61CMinls1
x3+ARMpjw6oy117ApddDO06RM1ow4NzvTEjTcBHrXNLoa085YdS5XpU8EJNIS7qMHQgWq/hnb2DX
F9l66jwuf99/qioFCLKjxBxrpjpv/Q+jahDbrWbtMIZgkj/MwPZD2hUXfGMVR939PSzrfKiVSW0s
QLoUm5I5rfpIewSUlDM6EHib51kqQLfdEjaWSYkhzjkNHJGxSzLqs8VxwWX+7WJGxYUdzClOcoAn
gnsFC0Cs9watr0I0rTrV0erN5AcIwR1F54m3NAQ7xycq8Z6x1ceJrGIySp4lPZ8s6/6ANZjIb/Pw
ualtVLC9Sxu0YJlLxz6yQKbAud1bPH74icC8mwVwRBS4CYyT+zCjlY4XIH32fMnkd/9+DKaTQPzR
pnFSmA32U6/6zQwjdiUutNJm1eX+WKobcTnhUIdOMwzlGISub6hYs6xdDRoRIg17Yht8wNLQ8eN0
0p2F3WUvA7MzAsrbPl7qxA4Sm7Y+UxJBRYk8oQI+HzJejqmYlucHpFDRPLcjfP70rLdGxzhP/WfM
jYScNy7m2r/WrDWyCZCyprZ821Jn7ZXwWy+BUGMn1NvUVVvsFciSVFXGsVTTAS+RpwtTzRuu5uP4
1PHn4q9CrASquk9I1JILZDL18PE2/FFIzKb2nNlHfdFZyL5xDfInx3p8db6WNXFxIc3KI+c06i9/
3esEoXQwmii6TNHj4OSQoh4Hlg58zMnmHWFR1/SCR+nQVMhoE6d8JIGSadS4Q8MkFzORk8QX5DGo
SfYW/PEKPhB1l7jK4knTQJje52rgv6wu1rQBeYLqEwa3BSiGoLLKhaPv0Thrzv/GSIWqXdf03DmM
FkC9AumKUUyPWCQ+z+nzOCLxT54a//gDudgHFDGSNzvnrXRlGGFQcNZVcXt7QtgGB3XnIa6vsZEt
U+IBOnMgzDS5eQ1OBddInSc3kMJ5nGfUE0R+fwCNkixa/FS0wuK+UqqhhNZWciNf0rkw0Zen04cR
kdrMxUwfmv1Kmh5GrT7vpZo0e523dNLWkB3v1A/SBtirr5BcnJky6fcAK+Tue/3lQtxNjTfrCOp1
nVB278WYcGS9YxNJWCggJXsNsjddo1PFVRrl7pJrXhjCjRYPfP4JthpNCCXqUqOOiF//G75IYvqs
d31fFF/WWe/+irZrCe8mWCORwAY/4oxZyMV85WiAe3hjhPxiCh+jdHuXEkhKaWfVmQ9OoLMrTyMa
PKzsx38w1HdSaKnvG6pn8SE4k2XBmtI2Ifv25O4A7xkhIGDXI7sWrwLUKHDG5LzBNI8SaR0czWVD
yzuGznhz9T63AwSw73PFiGu95aZwziIg1cuB//y2n1bhv07LWG1MSWZUagYmT7dTdrmbj3aoBD5K
Paac+Zf3A6KH/hAqbtyoDvKPUPVJCXrrN1kjqZ/eAcPd8b/i23e1iKmFqrWo6anz6fGfxLM2rbaz
HCeqKVY5TQsXFoxp7NK0cjb5W2m0NBBTzPwEE5eWXiBcSvr8ivv4OjiyIerV1LAqJbNvT18ld1KY
qtXi7PGHsFfycm551oiDgxmO1jaWT3IPyehUImllPP5G12OL+FFWyA71ItW3y2ZXAdi4k/ZM6JIq
TgqurtZFZnD9xurOuKI44UAcjaUIG/1Qc4lM5EPlmV2EvNdt/0cP0+U7n6uPx3S+zb/xFYEM93Vl
r2Tutgn6A/L9O6wbE7Wb5oOuwFCXUEVIOyWFQEorDhmyxXXA+OZg77BfFaKn8BGhSXfnOVBC9u9a
ADFbyIuMBhjMRrKVQJS/wfQXRWxm3DDObLmeT471W1SlCnUwyCM71ewWrs3drSf+tqEYjf+8TP2P
iWI6IkXwOfpTICXBiyMQsBs85xVBDSJct19TKKQnEV69QpFfX+D44OwOiyEdVhfuoRdUvj0cmxf8
WEToSJTw5wUvGp+fGNM4OkmQPT2ws6cK8RTEHYSC5NyuuO/BrQZtP8KqzNpN3HZeJ6eFPiEaicXw
bh8+yasNDJrYTrzXgc9l0UXcYKUszZNEmiwfkgPyNHDMQO91OALMcopqE1Uy44eVb8SioZWA20/O
bs/3suWcDxg87bYN1vj51+Pbf7EcHBCULVaDIaBwk+jM1jrkQ1uHmbYCpUHzCBy32wBQaQPpMDnk
kxutTNwTjvL+HorYrGMtgdE2heYjWFN+u+YYIDNg5+NeYWJ/O4AeXDQ+7n1SvMGX/hUraDtyysL3
cIYDN2vLt8DXxoZi86yyg2eWTc9secpaNawBXfUdQkuNieMiOUZ0W4EZ+oHVbrGOxoevPC6E2bSA
4jjeRRzUQvaMp67auMe8MLnscCDLzRh0MZHONW+/+Ir2Kb02c+ZsH9JZ9y7y9iTrey80xAv3MBgL
Cj+F1VRfp6mX9IC678p8rlOlJYYKmjV46yQE+LarPDDbURDNYmH3b9yVFjhhG2osm3k0KLa5vehl
IeeNmb0y0tZInx+I39qVkX+COlpVvctFtpth2L23mCL5pAuLU27J2MK9fzb+hXi4mQ3SXArhRLOq
TvwQROJKkaRJ44IsKPKckS9718g33Wg0Hoq92NHgO1nWrd9pxYjI5PMiKYMGdIDAon8RXCUsRewk
CGK4qK7yH17MpLZyIQxy2HBSHq+wLoXJ7GDRwkhnapvkTX0O1JZcwvNlGfSDVYCme3tnAvG9PqAY
OqAEuJiwaUeBh8ydtYTA+U8Rp+d2N00R5I0gNjs+KYTTvkjR69bW5Mocf47MQV1VE6ak6JhFLqMQ
pVg6ZWGODgTajDS58m0zCy1O5gDTQk6uYkFS21TOuVZyf9E00B/8vUaUmPY5G/3NOfR4QrXj21fk
yb6v1mJqWVn/3EsBey8/nnNdCW28O0O7TneYH0rfdCp356mKZtN9hBCN9+I5q5mdLfh0JSefeaah
hCmeebYKNP1LvYaAOWa/UlTZ2W0UmKDcKe3GGUifx156MTravFqz/iXmzf9sFM7WgfsMZMq0UqJg
zm1KUovx9EUbhTsYLKsjPyMbl6rgSWq0TF4zJEYRS7dTpBBsGcrQIg8Ylo+WxcSEtQyJO8yNt4/r
/d/+fBHk8qM7TaZEzoPfV45qmqOLVFUYpWcL5+uCPzEiSpMxUeES8O4My9JzbSb9tNCuvvvhbZbJ
OlksA4M3OIvGHFzGUtvhSpovqUwfVHTzgNzN4mz1aGjiTFCmmNfKfUIz7/M78XeH07+wHf9K6tU3
8r1GsBqMn7HTaQhkTrpz/maRkZUjROzGzRyF+lNvB+xsFDYoh8OO5f2cebEuUUpgJ3MOfffF4NfA
2V49jAdKRjpcQrvfRr7VVma5DRjn9KgfuVXlBv3HisW0Y7UjCPT++EtBknERJzXrXpoA1WcSp8dF
JoGoTubHCj9j9P9fBYKDwvmDtvRgs+vbsibJu/7mmh0/bOgGS2kOvthxEdrtViXkIHvbUaZdX76N
20kphxY92s1h2UiOw0P6Ic5xYfTdOq55bxR5I/x0DyD6C8831oIKUJrJovecQv/rd81tYhWSZnqj
oeMQkpya9k5nP4MN+WbgdBR9c3oYVtbhebJ7EUxOio/B+nzBIKJDtT6+Qy86//hNMg07ceTMUMP2
rQVe2cP/T9Bju2pI8nxzGF2Lc8CC2bLRA7OXGFK8LR7/1//FQpXL/PZKXWNwsCfyvwWse+zHG5gd
LQ/YvA9qsoA0++d+6bkEa5+Cmo21hZo6Ka3EcE/qpKeV6Si4R+Ip83bC1cQ/RIpE0xf8TAxvAImg
TEZNbOEVoV7WEjFfNyBZU34yZ+5iMHks1sHPIU5yeqJplXZDBffbxaLnJwdu0McBWqSNLDBS9IPV
1aNwlH797jCZ3PipInMXX4AeEUOL+xTpiWf/58m73W26P9wC605Wiid7Nls0O7edH/LtZblGCtWA
qZTuXWJsm8mVQDYVl9CppXfXLYRAImjpPXHpbX3US5Y009OVeuiuWmmRqGu5J9JjNxibKbliOxvW
a3QQlUDLDrfDKndHYIYIsMwKSXm32PaV5O33brZdX6fv4UWpyMAW567ztHOcBAK6zLzVjZ/r5NZc
1oNvQBcPa65nGaveIytPVAQVda+nXq65whbokpmNk0DAV3w4vJih+kNBvaRAtLMPnpYrd+UvQgRE
B1imTEk3ot9KHHENwS9K9rY7MRtrwpSnZ1pg25X9onruGKAnxIBItCHbXTBdxYO18hPWeHiLsd59
BP0PQEZkesvKuD7S5LkBAJaLlGAjDu1CjU+0DqOWEAFO7dD/BpYJ/IJYaewkFTfL6Jm1o/rrz3L8
iVA7jqnqXEIezc/6+KX+MzQDMiHOI7GL18MYxXPybDjewH89xkwzdwu2A+qQsxseDDazssNvG/JQ
vqBqBjwWK4QyTlOzTfmPiQ5wGL/P6eQAFUH+aKLbzq8Btot5WOvTyceidYWQO8M3lxFfGB6Lpy9D
aue3bDp4mK5WDX78ym69o0LFLY0M1bvgrSTDRSfk2mpItp3DuZ4xX8SRqmQAcMfZ8UJ890OlcR0O
aVyZaMZnqH7dsJilJ96NJ9iPwDbrKZe7CPThpWX0d3OBbWIi47VtFhlRf0Mh/PeT08GZJl8tBmEJ
ho1qhuqVo/xCfdf4ReMKCpddKgIQQOjZ55u5MZxniU5mE5gasQJufD3tugjP7CqpcsYlREQ7R6mf
dDvPWfwjMblmM3ckYsqhr3NkrNVUUMbor5kTCGRmg/a+9+UT2eM34J/Tdpk9iUCTbAfrfRIc4LL6
Q9HDvqhAzPoiPkW1bVLntW56RUNwZ0EoDJvDCqSk/XhK0atWi2AO3pXaHp76Sw7DPSuwtddq5tv6
8C7ixdZ3dSPDU4E8662eEe9ZblnkRpNxkdeeay0Rqu7qBDsYTOCNX1t/OMB/RR70a6JuzaW6kDTO
ZaRcqNREtLbrbvt59ZgmnAc88/8bqlxo5zPG4hEFnlOtCJSNJpQnw7Tlk7gXrlSp0ogv6LipMjAZ
D1PHJl715xhLUN4y8lP30f26CyhXN5zd6v5SN0UehNswerM3mO18B2gHQYMwDU4m7kH+q0HeUrKD
jtJ8tDa0ONukK6+0ETWBl8SqouRPxeSt2Rzb2h0C/474WHblx0MwtcFXLbGPHs6mUV5MLx4xQDvq
gpdXnCU2QrTBQcbAc+OUEY+7/aLUygbTesPDBagPMEin73jLphGgfMhnSL5oUfWcuOo97xzWeyK1
ld/FGY9szUPnJmf/6VgyvjxXjwwMlQD/cTvOX1tPW71hEYD4I1mXZlJOGh40mxKMbBZaae5LEfGP
mvvNO7loGM4J0XEUBXm8IwxlJ3uAEX4uYx0LodXFBlFhrpdshbeZmMLYHfPlGcftY/npzicgslbo
SFMAiMMXg1yzjOP+Dk80oxdl2pin2LLmNqAZdgGKhiH8G2HVyWM6FFCUqmS/aRYsidQr3yJkmM/j
CSrQpSmsav3Dw/i+vQnCFQdyESmgEldhfnoWVCdL2H+tg/KEz2gPEyG7hD4vEcCjEoNzqxl9r8lV
VxFZcx348U2bl5eo7ly6VcmC0p46aI9EH1v0erxadfVKlJYsMMPhsInmzOFSIwqnfyi28+abHWvM
FduUpvISK6jqM0egqxku8lv9QZ3pu2pMPUVRPqvlCRTI0eSYtGF+T0km5v8tE7OP40+caf+/uuO+
JrmyNWUDN+Yx0850Qw3yoTLyqEiri5wkLbYuAK219gh50jgiwjFYAZwBMskpWuIYuCk/x5D0+BkJ
bEAVa4rKGn0GrA7a9YqEqCHexVP07TEZXC5Fkv2E/FX2wwGp+Vz0ZoszaCk0tM0s8R02NAnLBwLC
Vx32GostTr55MEDtD2G3+p0rVvQJ3EjH3BosVs+sDAz2SDwwwBMLdrUtbdAfHXLfxUl1SNSKVa+h
aJXO2EStKwnu8G9MmQzY1FqFnbnJMqMjWn8PUVmNTRNoVBcbuGhVy6YFSuCZgL1HLI3Hw9LdRoMV
OnekzFutwH9o/+Q9R+S+Qbgf7GfsmJdxiEo5w48pso0RNTJKc9aS1ZOnYTD00qberQpY6vVv1MYb
OemMaSShoq/n2vjFHnJOA0xB3jHS1/msijIhhOJNkHKhu5N0AsJgGp4qaxClVwLWLwX7HHiZVb0G
JvWsdvHtfS8O8pbI7k4A8M0ZJIr3g2VDxDZvsVTB9x1d/bw5aW+ZBbP2tEhV3K/0F8NzVrIPQu2K
poLQCWxLCfzMjmVEjbccS3oJhcqaNTxExTic6yrvf9M5jRuBESqc3KzykIZKTd5OKCErM73uvzi/
5wr+t+ES7TvqCp5b9KMXxbOamwjJkEM+wrY2Cf3lQo/RjsLo1mllLUc7C+XLLMl5syxxqfhMl9k/
UdNf68/V6+xYR+LVpgS2jC7M2g8USYqY5f8JCDekk/RLWyvghFGrpfmnvwHJwwgfqCAvClYKZhOg
HoTac4Drq5g9i3INJlpBR8xFxizHBempvxCSK89qweGHTGclNss1xjndQSdcahnFLHDv07nGzm+P
vyWkg99r2gEr9z5qdH1Gm7GQDUDwPBr98nHsgrb8qnEcVLnyx+6Ut7vniAOhDwuagMCcKH0ZcGdI
GAhH5R60nw4sUamvTDg3ED+L/OV6DmNUcBvYh3BHOGY8Jx3GisizkD3BwRDdldFw5PBFNmN4Jm69
HrOjui7YzvymVbbpe1Q3s72SH9A06BCaEN0bH0UTM6B3Po/aSl3Gg+tpKzH6PX3Mfi/pt220AFKA
8xUU+/dshYdz5RAAclZmG2PynQi0sd/DU3UHCIc8URs2dNIlan+jNaCPn3TyXD7/ZWQkAMMLs65B
MwxP1/rIUm85trJt+Rzlv2RHv/+21Yb4dxmFP9D9RQ1lYNNMM8J50Ea7vWZrPSOsqUOBADx6EfYW
bHSj1WqlrrejMyR3n3zjoSJaK1uSlpouyj6T4QRuHLJI0k5cVUsyL2tNUsnrv3tzxERVwstj3jBV
qKcGkY41aVgd3Ok26pdotqsCSdF4HCP7/I1YZILyJS34ZzXFpwAaDlaZemNwwatItHAu8H2PwnjJ
JSVW1TFSv+oVrB1Uef8iuiTNKz6Qo7qDRayHgXo2bjOb09Nx/jofeUehkgGcQMnpdXjZ5S5NFOGQ
0XE7jEr1IB64bLPGN3+h5Jg8R+kgrfhQZ2UpjZcePikdvvZKBtgU+Snm12+PgkDp2GDDIFw0y+VH
DqzRZns/5zR3IsnhzBfMfAOfs3c1zJD9+EFHcIOFxkTLF+EaEr4kmk8MgEC2z4eI2bJER/KbubmZ
6qDTIuWc3T5aa+WmmmHFftBBKbDHhKlS9cqMF1xfDYJX9woT0eCq01sr50h96zAC8McTQ2aFxjSm
+IVZ/LYS1KFs1DM5r/N+AxsDX9f6HRG8XXK/Y/xtFnjvEIt6PHsrVEs+Cj5apFmMrU16vWscj3Hc
YyNB/bvB+ocIkGxd6rMTNy+1/xhu8yumP2sarGCnxjflEYBJsf96iHXtHz4MFJz0+Fc12b+oLwOY
fpnmvZSw/EL4V3riReNoOLk1Lic1B4FUy+Gm6StppbJBRk7UcRDszl+FFjVLUNCxqdR699Uip815
9pWVF3Kcj10clPAuGcB/xdhJYxIwfdpSXaH+qzQMhU1vp+51lNn6sta70wATcPhVbCKu/V7VShLY
4YzecQBzJTaT/Z9kgjKgPIgCwb8jYGwULib9sxxDEY3oTiu0wvYAA0Lum0b1ZCtSn7C6ve8NiHJW
CQ6mzOUfkA6RfawtRgojTUDs32viHezx57zp4fwnQl3vY5zObOrUbSQXg9mMx++Ug0jhoEhxy3DN
7+EzbIEx7Wa0cP2gqup7N1AZBcT7sxkJRBP2Cggu8KVpqEIO9Gk5DN+6+KPzwwUVtGT8vk5U26ev
kwldn6F90hrySGqci1d92+pza3m3gQt+d7dfZAT99oEmo47ax/NccheOMBMF0OF8dlWVoQOCMidh
MG0XKgVCqwwaHatA55xtVdkBcwLkjygmGVK4Eynw44i0ePz9xWXOwJHOa6MhX60QicDCcd3Osuqj
MF9ciIciSFg0Yoeg7lhQNXcvV4PDpTIe3CAhR4f17Tj6jHhe4WVjSQ0svFTWJqw5kTGMwalD+1fN
+0H2cB4ByVuW+Qe/m54q1a4dM6X89agSoXFG9rdCHA2NnoxwDxix4UkXlPqEUXFmOe4rkPYGIX/r
UuqgttumlJcdFXfxsSckf8akXLrTfD9D3HTNXe7ze8wm0zRRuuQIyTt6X3g6z2jyWgA7E13oEhE7
waUP6jjoMeGouLnLmN4mIRkmsksuwDlMe5ZZt33GjEKrCTdrOlPT/BPQX6+bjK6+k3KI3XiwnLhz
xA5NiOuCrjigBkP2N67XZwJZkqEpbizDIVXeuivJVPchHSEYZuvnOQ3xbwN4IpLq9n7asJXJn2eF
gHtNDaBdpO0G8mK9EBx1R1aw7/KEOwYt0SKoCBe2AwrKJFMX05zvdta80v/g4uRE5f6WXKyLCxoT
2SXUCcgpEe8Qo2cW48LyiqEZRsQrfWLqJVycKTa8bI4nqTm80Bdj/NTaMcXuaPr6PxiXdjPnBxpD
AK9GlVWDqotlkJooowF9TmTIvY1d0bzWJdLlN9/vD62j/fXxRyHiGnxWyD5WVusr8GQ2KRwS3uze
2803GvjJnBPWSsCc+/OwRNKa78Npd2BooI14qyDYh11D2gZ8L5R8MC2L6+TuIyPP5si1wuWOe9aG
37jZZWZLzytUa0oZLoDV6q/AdQR/yM3X6E95LRrnq+vQbhDepqDXzKbJC4COY1Wl9C5oyw7B/Lgy
Jc3EULWeXWCWyEy0mTAlH6QqvvX4zaoymerOuM1DIfNGyGLMtKbx7RrpmgD4KYseT3QVqGrFH/Ue
tYh4F0Y93B1SIzfn0eAkPUdWniQCn3XVYz9PuypB3+QV6B0z1BUjXAcRxAw2I0R/NMi+xGPwC5Ya
o6tm0H9v97eW+5g++c5wvW46wEik+4DKXFCuHkwyfnSRLQYUvNe7h4TpTC0B4JVHwieOWbnhBxES
KkFx9STLyXKLyZ5iMcIMpIGXQqW/WpBufEvCQqdzA9PFV4qMuXjvIL20cVA6ELcKBFWubAwRnnf0
Z89o3419FsG/RfzqXGrKJl41V6VRkHZRDDk3GtS47TmxnGcWS1jKaY7CpXGMuWoziY8rChGqNXbR
Yfwg2m8iWbs5dGSc+W1VTlG6sq+in9NL6N7t8ahhmopTldj2+YYXkdjwlCleXLdI95/DXQU2VCxb
KvXOd1By8N9HJGPIlXqK0Vul+i+li7DxMbrtPlius3G9YrAvZmo1vSvZQCtjpnpQa1XUnJVi11Je
3r+S+cOEhWPj7Xo8aZeEKCQRKAzJQy3n7jFbe5wWwrVi1OVJ14OS2IKP90X16Xcwl1FnYWZUSjVy
JXNKK8WjxwaHoThd/fIASMwXVDURX+1orStiLZWHHSXxvMjGoJXRmqXK/51KCEHJcQYXut9Y9p8C
YYoBFF6o/ST+jo4/dUjuzmhdHCD8bpVfjSdtyPUX3j53i/uOiayRBFE4Sx9B+8jduxw7UjIyv7eP
0OFlDzLei3P+D7C1M5NJlk/dlnkGGhLjlMhE56020upz2f9hwhW4xc0VUobwxLptERPesftoVVmI
epOcfVNvkfLGpFeKwSQAw/Zs1cWxla9IM37XTbX46FVfoMHpvECT7i/UkE63TcNROMJpYlbrqka+
+exKI7D9V9B5PRjD8rMGqvKMxymp4O93xRpmN6w8a6mTw7v15C2yVl+pfw3KRDsM3en4rIIbhr4i
gMqKe9KXcaF4Mv784wcIcCKD+FpJRtKjdYRoVh3E1tQG/Bzfzl7iNR1Ou+TliNKtULu/eAUbnbKw
dMUQT01RoghBdAZL6+FmjX9TqAXXLLe7SazRG1WdErnyZg3vi1hLT2VNclGr9Xcmf3doZJcCRRHk
PbkodDmR77fIuoQMfdwuHvr1GgQ752NB6G62ClHcl0V7AY/gbOIC+5ZcCEf89HwqJr5BtQBkl+zH
vv3xNB4umRUaM+CVQ632cqAowmZwKD+SnjbRfLtdbsPAq6H553mxX0PxNsgsXqm3SYrPXflS3vqM
MgUNZ6UDNke2iq/NMZghFf71Tf0tZsoT2ALWlGAvhEf6ubQY35Y98ZiX9BojfxcHVyXt/s5OcGq5
9Wtvya1k3VjkHjmoq8vomPm76bW375chPImbfI4DLfpTip4I3qeWEI1z9MRkl/7qZN3dBHnrrXZd
wEYENtKQ83WNqZBzeeZ8QDNP5+U1DH9w7VbWXS49hsddyNDIs4H+TqfsBw7DOGbQnAEtEKmT730q
T2EfNC/gLqsUf3ftxU0ypaAlGo17bqwwJfixwUEO8Q1O6uLislQihkZfvJycMCBn5AK/fnla7KyA
WWWLSzDyG3ghtrLU6j/KHZbkW6JDNIl+cH56Dep3xuHbXBvIjbMgLFa38bPNOmtsW6nwIbbpEGAg
b4brG+ma2np0jjA0bdIHhyBX0WieB55GKR203MyQt7fv+K5wCIPeVXrB5s1oLD890w2qVX4Mbw4U
nOEu+ceoNaNA83CFuqafZOp+hv8xFTt17s228sltnULo/uw3u9z6zJaMcJpFSx3it9QLfraLCa7E
Y7h11pEG8Thj6kWJfN6pTQ+IOyw2uANosKcY7uRqly95xdzhacWDErYj/MxZldXFd4xV0F53eNnL
rl99yFgmfYJr2TWjd44FIOWpX0bXuIa4/5O84eK+K3ShEOfozx0u1V+m5x4a4FNctrX11YKzghJ3
xulqHguPhBCNs8DAk6tCTUUNzg8nXLndbV9uatQb/YlhYX3uIyhybxce1LBSQphb4dkZlFQGzKJI
moumh478vPJm5k+iYsmMo3YVHXLvBloCslQL5kzrIWRt4Eiv2bi1i5Xj5rW5H78IDBH0J6CAmQH5
f4S7Fb9wDnRPTlgcLHXxXkbHL8D9frdi1T5jHWytYlNGWz5zFZvg6seXd4G/5qsx9LxE/vIbilyJ
1xh+Ix5WSm4e8taaON/I9QORx4RyqenYkp40+Olie68OnkrBIP7AvVPVNu1bmMe/ZnssHgdQHRla
EoBRUFhlviTjjnzsfPNutOAPdUhcgVHh8LXSuUoCJM7g/EszteXOS85wN5mBsp69T9xzZ1zsH1wG
B5cSflcYqKNzRAvOD48UQHe97Pcka99OyszMNwwYX7s42OE7wmIeF3XFWzdThNF0VGyRbYCrKF02
o424CjcNLnS24Q/hQ/ikNzKXIawinMO4QB/dA86vywlViGsJqAbQMYbOP3KNOn9gZ6G6IVNHo4+7
Ak4fLP6zdaO43cNANMF5v/JHXnYTqBF6TQILn181cpHbAO4Ktl7mSiF2BWpMm/tRPCols88286fX
GXEHqGXQfO9t/lUO/J0yYtDJeMyQVi3xeMHLEsZOZrtf2swEGPQ6K3ex1xFYZoRw+CgiGcIwdog5
rUkIjAMhezMKxrzPL3gVxZCTw64M7IFctIP194ZMH8rcMXPp/RlVG4EzttWAW9oKYzN0TfplSGJx
EAQk/qnGggUld5RaC6gDZPRS6TXr0oFSrvbuaEhP35vcnQyrbEEh2yEv6toFWlLP4QhM2kIztK/3
xhoo8k/dCPgC/0zJZBWE16rI68hDt+1+A/MxDu27zbOXQUZkFh93rd493HK50NGMUihlMnLIkaYY
S7iDGoE064FNml9WczCh/9iMUh/j1JzHJID4TR2N2e+7ecsIf1htvo4digBUVKMG4daeeWObP7ug
YF55lpZIcmjZs3piWb7cBMXhLasc/8S22XfzO+AKb+PYgDaOn1Id+LAa/IZz3Bj9Dhb/mRPESzx/
RibSO3m4d2IK5HJfPHHa/ywuV/3d2f61kCyrm4Kk1cyh+n4usFRUdv8Sn6K/SS45BJq+H4XBoKDP
XnwMshJIz5VA0hGvpxKTqJsoGNkdysjp0GpEsF94IUWE3iGP/kcVz/QdvzlfG5fI3u4dcCc7drCG
z1Nhsn4jVcaeGSvrtjXdu4CLFjHAN/Z9Uh/E5KpgvihHwg0VL0Yj47vSzwUdNI8ojhVAlImGCdWi
FWhtTvoYdirxu9P+m3uiUdXYlNzC9nfCVn6iXxNJoDcjkJ5aUdJZ979HTHN/8Ie7OtAWoutiEts8
cxoQvsC3EivCKayldVhYYFI7Nh6SBYbNcPwdiUw8ZbgjirxOQnmopw8c80J3C77NIc+kXoYcOIkD
Gt0cvUUEvTd3Kb+XJci/rZFRgr21SXJZl++y9OaSF2EDcdYPej4xm17FBprznsTe58zLFMGE7Ctb
UPrnwEt0g3PzMVTe3xqoJrMJcrX4oXr46c9GxOcrF/Ksahv6/0BfRhz8D7KWYC8uDXQ9Cmd+TADH
MnE6nGkEzzUUVjjvoFD40OWLlXoVh6i5T6CbwOdLiNxWISWjbuqjlGeLNQw4MT/UUK9cTlzO1gvj
cEiJvyFlklKITss86AuKeHOBV71BAPHswOPcHLiwapoCALd8EpJw5GLvgR3qEFOaKuConwb14sPK
QGdn+8T4xiaLg0ZpEdW3/k0IDMPoGtlp2oNwzj/6is8hWSVksWOLmi7UAaq6tvYMMPiZgjkcNQm0
glthSkiOIZJ0e/X6qL7MkVEnffUNqIKOzjfaNJlaWq6E7nEakWdrwj2ZHgKZIGnZOlzwyWOFyitO
NapzGrMyP38FrEgSqQkM3SJ7fVrVgByg5PbyWZroLHpFS2gPIWFq8DaTrKHx636++5Ot8Iftm3uT
Z+TxAAdwfsqHe6UPE5DalbUgG3maL9vXzHlfkZcktFVVvRD5bqbHkiKJ7BvuQcNFeTveDlhn0+At
Ju8xODKIDgrWVz7p+XZJ+xt8yLKc1uZjUqLVSrhrvK58jPpHwKnlLI0vHBArVKwBU6ZP8ejzWW6m
fV5pSoQTxdLkP7UbDXkKvcAJKLp1N1LvnfRJKHydrvzL2YM4cSvLK+sUbnSD/DMz+kAhj+7bwDBN
qPnzJ3LDpQKNozhzma72hHD60yhS0/sK1zZyvUBqHyLIhWLAKaVs4gvP1Cmv2rVUhs2Qe3acCnui
O3U22QrIGYUHHbzaAuR/Yzmhp1VIAQK8oa1vQrc+PFoY2PbroCdpjjTxmbX1PdCj8ZStF+pgAv7W
6Jgk6Jn8vXKlSfiFA4NpS41I+6IExBWfLxxw3kHWDhfnd/wm3U3ECVqf6fJfiqnmuybw+qaPRNkR
ZzaF3mYQ0i7eq1VY9RWnnax9+KhQ+CBHGw3TZKBiNvX2szUidsdJ2dmqShheqnoE8OOeKTHAzNaU
TzGQtNXtgKkmA+5+/i0PMblrtALd6efgOapNqMKMsPsWRlQrkIV8X8jIhZeIPSThF+Zce1HA9jzx
hpjppCnikVghsmQdA362DM43G3Cx/G4qu0GSBPQXACiYOSn7SIQMXxtOEMq/Ii29UT/a0V9MPcqK
ZSuxfS1kuCCwD49OrOjo2Y/g+hT7GCadvYVBBOe49DpVmGLBKWqKl38bHeEQ7GaN4PPIeyKzfjfy
nJWHze6MLamr4OxZZ9Q+NdT2/HOiN3jYrwg+fjBIG0SnAJHv1WJdFoQ7Ki0ziXIoOQERCAcIiz8O
1fpBYXdvrFaMQAEbqM1BKFvu+T529m7+Me9usSkVUQoGgvaOuPyuJTHjqeARdEtRkS8Yv66wO9CS
QAXrnBkor/oFm+q73FhkAzDoDxXtwAOvxmP7smgVnyjz+nPsQPDG7mUblfOVts4szo5AIrkwWfBx
FSoHkg+7fGeZAFnNF3VlUN/BxyPC2EyWWkU+6Jgrvm2xXrC5taJgSitqc2G6+2QGNJ+IwaZ35Ty1
1cFceW5cNf1LdCJZ9bRyHqT0FmQ8duY78VQMxWCK9rdQ4DHX6ZQz/aNTGJ9DTMdDeRAPDcrnX8pr
za4FYwlwnzGoMscRNnPMwqwUVhxRRIVRV+3I4DPQhBQG+kL0PiKpmrtBmFW5RhPddzBdX7XjGgut
ARotKpFYOEERM+r6tjDrZcNozau9X1LLU4vTRWbnp5cuS7cNnoRUdxlzJrYLg2U0d8lRVHiJzT2q
LXcjVVnsa+EPSAtnO79Rct+G40viQAdod7tDKsyW/s+qfDgr80p6nEe32TQUWzt7I9dZYsG7pgVl
NKmo5e1MZYXf/H0k4EM2oZ4Bgpv1KA2SS/AR/bsBGOOIwGQWKsTLPVxv2lPs1CDaeDNYekivTm6f
rCxp/LYj4l5jZLNWElFkpN78tplaQFEXWANSSbhlqc0jiYKT/KMaatTrP8KJrhayIr47alUpKWLX
qApfXZTd11yyzr7i+PfipKrc9FhF3QRVxu4Q4zVSh5ZFoqmlk7AvmggBpOoehzFGtQcQ68eIUVsQ
igchmqKExufAIARcB9wWyxnk0m0RfHz9R2Z7/UuLLbC2TJeMFL58i6fw6IEPwxjE9V8QagonHtsm
2Bw1RdvuYY0EbTNlBmHOJLzyfFKGLhI+Qbw7fcrLcgTN1LXmxPzbNxzK0+JDp3l2dC4PN9M1mgGL
khtUt5jkoAfYJ9H0cXwd1j9n6S1DyowXok9flNr6WI69xpvAsd4NIUTsaEuNQ8CChk0TjAV7x9Zd
mGIFX2RjC6ytu9td/h1hay3EiiFU8mj/VdqA09l830pS5P6mogIcgUM/Vd4B3LaFrGX0cApe6uzc
Y6O7mi+SiAsVYHGSRz+tHJkaCIuJU8OpldKqXP+Cptr22eNjmotDhDblK54BXbYDWgevQbPzLkUk
Fv1duqhEERsRm540ok63huzlcl86ZncCcfSoAwEZbRTJp4eK0OkpQq3j8ukxtZjrC238fpZ/1m0/
PiXgusWQy5vRpI0QbCthL2WOcByXzqZYCJmjS6J75k/2sMv1CTlr7aLTzaP6KMWdV+Y9oA18369/
TcEAOb/bJ/h3cGtAxJ5NdHKvCRlO70nSMr/J8tUSgUsTNiQfFewUM/cv8YkXuMs3zsuS6cMUNSZy
0znPOiEYPIu3tgskQuMJUmoJ6XVTdDtsPbLn47iTh82kvUQj7/vWnFGCp6Hr+S/jP9WjIPP7gRUX
buko2UMlSW/F5ogGCfqITKxSMUrywHdbBf28amxFEGLeyTuhffXRcBuFsNPsnE7IaJpBfakMXg/z
mZsb2+WMmCoA3Io6PQMnZ1wOomtpG/6JJNkLITyOU3hWS94L7lP9k3uFJyokA50MaXavE5I04KYF
Ypx7/7ApNU9I9j/v/I0AC27wvyb5UXMfyFvqq4Xyv7cWdq6yezWyN+GQxOjBSZ+JEorawW/2d2WH
JtpigH+iDiCAKSHNNcviACv0tLXpqLmerdw99hiOZAnMSYmIPP5tFxIL2GWOboL7aZ3sEnLv78pE
uYgYYBNIOxMOivX/PNm5LAVy2DKt2Xh6rynC/BuYqyStxvpV8pAIGWSD7PTJU+n76f7rLp3HsX+K
UhXKMS/IE8zZVR+pEFNQ+R8AYuo5CWZN04CS+LteS/lnwl5NhQKPDNHdmYOseyi0m3MH7t/hegB5
YdARSRyduQUBxL3csPKtrHSEOBbgc8tsQ+UyqGqP1iQXYi14pfeit7n1gcM/mCn1+EvS+g9qxkmD
LjzHnBFb8pgeT4G7i8/9fhc3rPPiPdNX7aCcWYC0bys+AJRribLvQyaYITw7pdkGNx4BkEB3LPCo
v9XPEnXWgm0i+E7+UWAEF3XD7EugCkgD55PpjLbGBAx235DQdcHsS9VwErvXNtE+XDbPcL0T+xef
yuidJXjLfhJFZUyLLvHE3kmHnfDc5NOr6vtt+WIjbJzfSniXgBSOc62phGhLG+y9XinJGgPnzAAr
mVCeYbqC+1Cu7hLc/Z0X49sbGOjagbtg2MoaNrQ7UZA/taJqCZZYEgA7cclCwXhCDDOSc6IoZ4Sf
VnreIvGTZdzd+9YkBWtjFD8xW3qXSun2MTZp6XoBArWjwUZA+CZ0fZTCfX+0QUJm+blSHaLaF4sb
QeCUvIT1ikd74tkIfw9nLUrCfqZoitNISFy7/PAC647sA0lm0T8HuPe7Qp5TKEvw5xMQuiVTVvCz
eBxKNhxNhPDMKlmAARlcNkK1BnJ/pt3mokxoYOMDM33cUEFQjbQKeWVyMu33JYEF8gQtVXnHYg6r
MLfu7OOEumLRlykOVUj4rX2LB4cDc6m1B5mwqUYplLBc8TlIfUq1Gt+xMuPZzk/HBpIPXn8ONrgK
fGgfyNr/u4Nuuzu2udsjtQK32sdxyabPSFuoFTFujpYk0lYLq0X33wq6bk6sPJRKukJtVtsQpqcc
uuQFbCAW3Y0S/LdEA1koqAAMA9RPEkwl+PYVbdoKiPaMltO9Egg5nQTM0bcWS3tJZ/Y7kmC/MedM
qjvEe3uS0kbLs2iLcDI0FGCch8fJXE2prA3luNBIyfDSBuIugAM56c63m1SmkEG5g7WxFy/fvaUU
Z4F9qMfgnmC2JYy1gkjwa4VHTs6QB8gxL3imy8qLm898eRMcuU9ANHC56vlguzZEKLibS1crNdRh
ockZpbjT0tGa+wCozBOfRWISRl5ZHU3jEOUFT9g3S04oHyE2GPB+kLTZoPxCEfCPgzNGcWhveQI9
iFvh2yelVS6LQm0y2wD5dfELOxnshWj8WARvpc9pNylwe9K9M3nt26TIx5GeaHWanr1crk1mIZry
g8FCh+O+iUDWHzad10K9ebbW6tKlLZJxFesHC00n56xtnSJ0EuRxOJSaf2wOB0l2tiRWCjlHOrjW
vAVFTLrsJea99WRUe+dw/5iv5IvMyGEqOCDh2Et6EJS7FH9pNYbrX2m4Hbf/lUcu8uLgpH2Og4kt
zJqO+Gfl3W1/TzegTwhtL+l80rqs/fmWKmJ339xIywlzaSkH/qHTGR/SC8fSCDswsxtpnfqk/nX0
xyPRkFgu5j0GzitpuUFLeGzFaPM6DcvHVPkGMpc6VVsPdEi3SyTAkcvbXNuv4n3LbdH3RVIUuNYp
A+BzxFwnw57TK07HpbDvuC08ns5b6jini5oiapS+wNlt+6QwHfgU/56EXROClTAI5P5zVa5eBOGC
nMcoX8rO6lNv8l7fw3BKsu2WMPgrZPql8b4uXty93mXOsbWZacklClbnkjMu/Twmin/crrgxVmZ0
nLA5h8WNaFZ45Og2/bh/jJmfcDJDJD8AWeOqRcP3zKo15iIB7cSXcrMQjDiXi3gMq44lsNFiM5gG
o0sMOE3jE71PpdYgE3xPvVkYk0a3/PTTn8H1w3bkaLpFPiHEezWdrqU2CImrBjFFJpieHQtege+O
zXoUAseCETiHNoIE7VDEg9EtdwG5tzY0wsPKAMbURK1qc/WTRDkI6Ga+lWJPYAbw/5vHq0WOnobx
P8aIo2uLo+a92Vcj9e6xg14JPIoxpaFPwcfdzLJVyn1FWSAhZVuUgY9G4NNpj+0G+4LRf1V4PglK
P1yPIWBI5EJO8Y65MWBPVJ2ghhKvoDVxWFVp7TzMi1dGx64dKhNjyXSAeKolisJxNtTrNzFVeUde
He/GFLPvKVvp9UURm60hbZ+tmaozu0eUKX4bzFLJ4w1+DlN6n3JxsUioR22lzA9twe17K4H0UPVm
kENj9UmChIOgsqj7oqeQ6oQ5cvU0JsdQghbIHlZj9iUaNzNwXmmH8oEbdhtbCNiTcBjA88HXWvww
LOY6brBD/5Bu+ZEa3trkMlIsWDHPP3MVrpslQqCbMzJb/olzJ7idCKteWqF6V/KlJyYlRBkKs+ze
uhqiL3kFjDYhuECnt/xLnsYzLd63khjDKgeQLOg0ZVslSQiciIh/lF77oJkJit0h1GLmqFV/fKwA
A40XxTM77yci0J+67WfjABhTeSVxTf+wJcCPVY0VGwswbN4JXq8IZhjLvHcaRSJPG+qvHJqXYAaE
E9KBuFkbj1EWHwsAL4qR5ojlhlzZyyd2pvY5ym4lS4bi/WfSzeQGX9kL98rjmlODqPbRUQuE01S6
yD5V3NNKBta++IYN2WWGOnBGxPaw/mqxDJj+oFgny/NpmDzcbH7xsu++CuEw4zJd3PIhsbx2yUKh
yNhVBv6PLJiTLDywtOFsbHvgLCK6dHMCK3Kvfjwqah8hCAxVNYZp3JYgC8Sy4qwtbiugIGrghtBB
+VqSvf8p/+Si9rxR0kXg0l+kr8CFxIDoRoD1Us7hP1oOD+O3Go3M4FI1WUB9D+GawRFkph8XoYCz
qndQK3TAkC5TMq7JUj5B/Eb/hwTvyzsI9/dB2TWclxMHm9mi2bqmZHVNTqByzomhnvXYF+ZcbRku
mpl9DBrAYQf1oRtM2jXWJHA/MJjQIfTQ6Cz8poa9BOYM8fSTw9D44SKONCdvH4UmOGTKK0KzURB5
9GUkpxNcBNkGCFO74guhkIi84qi2FDpcl5UOy6WFTfokWvznrTpJsbTB6qwgTR8amfcpMQ+5cccM
CcUQn4LRdar2qo++pSJtDEZSH4wCsVuQFyGnnskCjplES0jNCsLq3R4yx2UeHRxME846ZM5se2Oa
hou8mquh6x68lew7vGyy0YS3KaVrnlkw557Gl+NbwRuFgh/sRnl8udd2nCbsGHWJ1FFUdsx6GsWF
NRDg+O56O5+opg1foaTklljBMeNsO57sh08tkLK3NCnh/CC1X/vYfElF+MhXlMbdUZKs5tMilfS3
9nuFUK4JfBEQIzSTxRmso5F6hv8HnjIh8lfx7/0xcWHM37pHmnSyGABAKP8UNDThKYRqsi+tv2GO
+o3hvyVFB7l6nDYdfQLAYKD+5fzodegZWo4TAXzdaXhGX5mICfVS+xUpm1tcWA5NvqooThfbGB3Q
PDQnKzlhgASzg+gYbVz93qm6qxjmBbxOk9TqOYsAt81gpGJQvQOO1KJf2fPIteujRfdclKqlO1JT
hnKalyu0b2CXAhBw3+weMP3Ozr5srkm2SBlpWCqKz4ki9LEw7a/5U8HcTeuPC4BZm2ILq7r7P3FT
dt2wS9r5O2qDWitY8UyF1DYGx4N2eSP0PAMlRNrM0ttUmE+sRHdXPoAt6DZ4NPYe5lfNIzX02zCP
Iv8s4Tex6PsG4iSe0Muk+pf3Cc9kG595sSOKE9uGDchBpN/K8kytrTq/CJSdvuUyZyaI9mHEQqMg
rAnXttRyN4dckSxnAK7i/n8v+qGL9BgSw3ZsHi8mY4XMAkXErTIhI0YAqmA+n9Bfv9phIvd5LB/q
0yzi/vHBuJ4dPFO9+31CBO6WLmJxjxm8Fq2GqQVr51Ucgb1/H6wVcnp/l3sUgasQViSlKyvFgQIh
Nv4RB0RrXn8YtMadazikEs7Raa1h6H7TLk2ygJempqd+1aN/HEyd9n7I66H9bp4QYTyv1P0B0/nN
Ec6+t5nGKItAK7AIT/I/jbJlDndAst+fw/UPojXy+C8ookBuSK3mt6sWMWQLVIyYapVwd6s2bDab
MpT8DAwX3qNohI5kJ6tYXmcLyAN/ZW36POhhdVIT4AvJIu96d0o4X6gCDKPp+5T/z1zkYKPVhyFw
OPifqO/GD/c1pULQ2X2P3gTuneG+QTbMYJ9lepfAT5SD3eqnYd2rEgSjw8jWc78iyv34q552/9Ro
MO68PqY0Ck94Wc1JNDH1dQFlbhiuGSJ7EGhX78S0JGtfgBxaM+WFzvmYlbEoQYvVzxflrQqPedZT
Gs9G8Ymr25NGjcfgvwCxlY7XB6Z0tsAuSNORawq8brmT0JDCZjg/NmAobxBWs1Kzyd6Zi2YPzyJg
3GwxqcnhptmDnUaj/9oFYviFRgQtFIXEnShKmeJ6UdLYNUk7ayepadTWKiEKUdptN2X+MEveB7a4
BsyOhHdtBZMr869ZE6Mq6ZI7NaNp/HuRIpU2Fe6ILkaeLTFPbVRIfCTwk/kmS/uQI74BQtyB0MzE
8CB7D1CuCs6y0z48HWaiXkXtLLxb4pER+vD1GomudBfUpjrVQU+Wog10RY8Ck8Smmu2XVlFMSpfr
V1R1d4mQVReypfgV8upyKM4GoMuE4p+/u9HJWdfyb4m/Fk/YQcAGTwgudVftOp//pvVEgS+YnaQ2
cCXLZ9Wpxr6a2NxqaP6FbqJaauGPgRQ7/68QlrMJWt7xaV+5QbI+Wv0a57dilB1cjMFB9nMvLFpy
F2Kv667sOQBAiiqlBbCzAipDWUdMYZoucWmX+L2nuf1HalNCVTFlC4mkTOT0pU7CnFkY3w2A72zO
WsxH5OpjqlS/gHcG9kR4UO5zf1ubXPedIsbvlE/bD8VnCDYjdQlJ/QB89m2WN2GHTnmc1wWuTbB8
yUoJ3HohAifr8HfMrWXrpA6pRi9PDmHKdBf7bCXW4ioyfjKEm9SPtp4Oaa3CZl9gJPXBoLRtcQyx
ODAWj+626dOc+ivg4cljO8L1sY4CltNLk4axd6uT04moqemR4MtrKwIrvAnLRXt9G7MD/sOxRHMW
RRpAU6mLXGTQUxgNflcNpE14D45B577tdh7/7uImr6BFFe7O57fKXgeYOGGjgIL+ipz7jWebxHEE
CBtNa05teWqketcJDkIh3ZyK+QiVZFVF6alTAB/1LaB4pdREw8LplNvqX30ZxNH81uDiDoYvUn5+
f5t3cTs3Nq8tQIvY4f7wnjd1sSQHvjR5r/+Gu3RXiyAnVKLh9tljZ/7wzEs4FIcQWpSR9QqtvZJL
WYpKTaGhpzfmbvxQqeSvIREBs3gh2mWFxjLSF+cGH2wu6+UQo5Tmxi1bEuJ1fRQ8y2A/79Pf0aDo
GzIZkadIS8nbeLmOmHMNeK98o9+4i80O6svJa5B/slWFtuaLykWMGFGgHDclVfyUGJbtcgURzLu4
0SoULRdmr0lq38zQaaXRAQ1IxflpKZMqquKF9mfJhjzMV5eHOBbj0O9ph2rLxvaGVYBTbcDyzXQS
VaiDKP4gNokNN2tk77Zwc8vjq4PGHM/gyxi6Xj/qOgvsz+EcgbNRRR2jQhAZYBiT0O5XBB1WQHZ/
cvBafqxYMtcfRDrSRNvhUEgBlYXI3oqpfwrcKAYMr/WOJLobArEA/vteJ3C4Fl7pGRxcK08Ksl8w
rmLMbL0oyyV685ZR2+EWybZ+00M9ePNTvvQC0W8GmLx0eG6NkCIjcr4+DmCesjBcHfomLqKww/rf
nKw3lpura6zxdqYxC3dpmnNnyGc7T/PsfOFkzWUKKa4v0nWzNWA0DDOZSo/FW0vCxUwAwttIAWtX
3QVxHjiMzyFrDXbxcUMHMExBsJFZ4ZNJT4djuExgUsEjNucfyU7mpkLXZAileDbSihsCSSXomQr8
QOCg5qxWz76dju+VX3/98rN4NDuxnliKa+S4wAnq7z5GJsrnPB4CDxTLmHYJjH6eXqPF8HUsICOD
9frq9AO0xXJsdBR29UdtrCZTY7D9Kk8hMpw6zHj3DyTWl66Zq+qRJ4hEEvlst/7BuZLUDWsFc+C7
Z0os31pFphTTrYYuhav5QIrUcDvp7mq+K5A099ip9mZIAZdBHMUp6S2crIfNgjmSjrOjqQp37Ocj
IOcEyviXQafNHlZqkUSe8nGUwM2AjO6vk6k+9ldon1O+TxOPT/HxCuekeqFGxYEzrD5PwFjeo2ob
USXEa3ig8uwBgM/Bq9azokwjGSRw/zNYvNA2AXlVabpg7vlHfY2DDjgZMUwH4ddhmf33dwRAcZ2m
YNzcb7ZsZiw+dlpvKOSz2r2nmJOMEJI/1r931VyLo/4LbKH+jjVoAoAHNsWwkfO8nsT920Mbj6M7
gNoatXzMPZpr52zaK+XK7hzOjrln3Nor2uhJOCSfX2ukKjBYA6xmuGvU+wczN5MdttNTw+JtV0dy
fhgeLJe+FdVHgXrlyqzb62vHRpWlXrvDDAbs3e2L+vahQwLVWholuadgnToHPY5ubKaIGZCtFy2/
pHV0KwMHvj1VNvQ9PU5DDhRjXBD5cU9fmgASYTnwylcUqb6NO9AiJqTw+eEre8POdse3n2vcDJfn
RZqFpxtBkJoAQcMvGwm37bsNG824kJqDf06Gjmo6wG2/X+JnwRWeBYIzd3szAaeqny3zFTHGtdnC
baOUaPllMfDoeq2N2GIac/ub1Ee4feZtfIYGNgkfVYQaXEluQt0V/gYtSEfqCc8wBKtX+pNvtiOG
gTQ5oOdmLWS8SAVaKb1sTBH4D/KTeaxd4XjCepCGDnd+W1evDiY6A7N0izzHpTWdro3x9i0tWVpe
Nse1+cxZ9Yzzta1IhtZ7phDjzWFzHTG0Vmd5KYq5sUbx7CQ1z3jBSFLd6VCBzho7JTg5+OwCYNzu
Kr8FEwuEdxUG3Q3lojhB3XRIndj1FzeKUz6KIKwmiEqeAZXbfhzjmTvd14wNIkUmuYAoTEkdKD0y
Czbv1TvtdRRL6qzv/WStM9mkUbfz30CtYObRgZ1njXv8WansBzvs3i3fFKp7mSnwCkQq8RsUeL59
tY5eDUswBbFKtHuMG8HSdJFdjnphc4DCbxpl4g03qiBK1JrE3/wRzWIgaG/fioABRsJl3iqODF6X
MbOk44dLjSHD9Rx8Y4gNAhgKD/bh5wdM47f+BaSPPTKHlk0tyEj2W+PzUQxy4HWnC00PfWz4bBTE
1t+cmBF8r+NR+JfKLvYK7dTZFKgb5559EZiI22ubct2hgpYIEu94epSjBX33/gqPafL64ukf6bNo
qVkfzJQ18ifJHF8VxoDEXMZTNArz/xn0cibcivO9zqpc3/7ANM5o4h9LaI10ZYGvWwgzPvDFihzE
PkGjkjsTFPPNLmCrz6KjhDPTDxWL+h1Muy/2ZLPYVZO1p1Z3UWM7Vb8NzGu7NQYvfGdMlcGLSVvT
SSvOgdXVvoM5JHel6Du+fntvSmmgXQHR0l6VuIaEv6I6rp4b7O1JOT3uijr6ZptxvuK0BQqQVO06
Vt2KH8/8MVGvzKqHsqibUy3+PfQyGBrjucywvNnzfrJrojoQOxBG5CiiqjabcWDAelRyby3oOSLD
R32AIdZcy+uIgrIQAp7m9aZhrePbRhyytUHZKDRVjtN7+1qGq58LTaSyChiKaxFbaHNXLg9B04Qb
xxg9a18cC1D7fjjS6TZ+wnY/3YdC+xGeeZ5ddIR0tUKy3G1nTql4id+2/NWCknDSBnmJFyOu16Z1
uNDlrDmZ9kSkpOqTv0hthV1l9UwJAAfz5NS99jK7ZXL/JhgBmSph21xaOHea/xkpwLQ3tim6oxnz
Ttau2zPiF6kIST8LjxiwdUzZwX/ZzFmSnX6fKoKDoBr7U+LoYuv39iGvFjCPozo45KI+UnylF8MU
Awwb2cIOZf/t0bufVpG27r9RLjki0lpxmx+45cNH9DEu+SokeFYymSzeu5VHL+Z1PWzqJSlBW7jm
tymLPlI7aB0Q+Na3hhP/UgAsAdHxWtrmDajkZwAcm+U94I24i1aIOR2vaDbQdVvmm2UfmRdLUygQ
ZsBtxnJ2RWLo4fd/ZRMTBEP0ZVQF2xZ0RPt6dtBCR5OQcJT15m8gp0j4a8EmHFQD7UuiEx3ltuOP
yyiOLdH/mV0buvorSD3wUWI7HaBHbg84OiXkciksxmtjwRPwcK3s4FLl8nULX++fDhY0Rus/xFRz
ClTiEzxmry1wYx9SVwOC4PymEpLdJVXoXGJEV+LkX1sVJQNoOiQhX/aCdcyckN6AYn7S/udjoQu+
yWYBGj0M+qEhK6sVzNL8yfuJ+hs/01dFNfIzW/Q6qPCTEhu4okTzfhV1ThoEtl75q6Qqhe1Cdph0
uJVrCkrfKYUYqKAJXI8AGg656A8nJSfz++c2XA+7IMOFqHxw6OFqel9ZV8P+wwyYJFYgxvVvJDO8
8g6wk/tzZGShoRAYQ/yrVJoZr1ldePdP0c7JzBqn9hK8g8/kdpKnn9FNjN8wcg7T+fH3lszsCoyS
JoUfAb50fns/ewGqmVPstEGtzT892Ny7ihCrD0WDXWrFx4VWJ3wy0r0wl2/0oPzeydXhQOG7Gf6x
+jfJZTQCNnN63XZgWWRV8h7JgADVB0bFCNgeif0USte7TLwrisCZB0AwYs4aL/LE18VUGltMexvh
/mbCjYW+7xGI2bXr3o53R4hKlUHqsRR10jEVznrk5wWdlPNfGspB7DnqfcNDRFiUA9z4ApvbdUZ8
gR21RmOdqKnlgzzP+CiAJAXC9aJ2Kp5Fg030gKBAW+I2IkUc+lxnF3N1Cl2jNcYSI383RVt44Dt5
voE/PyHj9h5AViz8tlvQTmRiQ8Bm1VnqeSYWsm/CDC3GiykYz47R4nl22G2Zm5034UIBtOdc7SRv
zs6NWYj1cKVq0RvSSpIhdSYsLqOKb/rtEuuCvS6sxQfJLkpDoRSY0OoNe7BgPJYekyEjvrEW6/Dg
Hxy0On+cJQYo3Lw70gG1q+qYXGZ/4KINuLOYsTsE7kigEcFHPR9yr9T/gZ0Ps8NZdPGz9u9nS2Us
EJoquqa7oIBZQy2eH+Huq27cuUYit34PjooQj1z5Hg8oDhKfFcGVG92qBjHTooj9MxHxIfgz/Yr5
0Uk/3M1jSrcBEyqGMSlG4VD7HVvNtQIMMS5GO/IWTgNCU6xndiHETb7VehcuUSyYgPX6OAfDm1Zw
ELh143TW0gssuZsMBuArd26idCac9pTH/Mln4hunL4Rz6DfOkGtiFpkVqLTDladv8MHitfug101R
JNoHl3zvQGgpLa5w/YRHE2ZSaXGoRA9tCTF2zHZ8XH0WqbsEnwoYI0YxDkQSD87AvqvcjuWjNNMp
jpsOSSufug2eNkKA1XcodcxJdd7ZGx55ngTd0I+R1BKaH2A7JYVT/rT1O88G+3mMahzUfTK2TlCO
7Ff0Jvs7usxmZmHPsA1Yk4SgzXExkpp8GW/Xa9cbvIuC09ZFby0DnJQT/92apZhw8RKxfPh2xORj
Ctx7aSxCcTSyJBV1ELbrZ4+op0U+24CLsBhc8GGzbjiOl2e901Jq4pudk2QwyGCMxZSBT4znY754
AIDllsar/Bv9eRxxMG/JuwdLwHXOqEnItzZR0pJ5mwawOIJZbpBkY8zEXgZDpbdO45Iej/wzB7Cb
3+84wfTCUOIGFYt1VpgyJGK5mX9V23KIPRjvKcnaSmJkE88nAGEwhX8sPjOcCW7Y+JfOe5UYmMmk
0OAhsD4P5JopEW3DHxwIWircYU3RilX5EWzNJ5gWhOolTzfd1KvObLMzV3PPk5vuXE7ZcwZOvYdc
GECe0LO9VEKzFvHYaQ20rnupmF4VZu/kTiRWSHQcgn8mYT8+5GG7kuMJnvpFFzXKb0DHrZmZYQGI
lwWTTmsJ+mH2IKLX3ldXYol95fa6k4YpcCOYHzOlbHSaCrjBKi4OUWEZKUW5BmsWizNgK2cq6PwO
kGN6R4iZyzUSpsTjsVIl3YuoSMhpwGOVll7/ysqyoB9/+OTXFZYfMd9hu10SYbyBLqc9DLlspsU3
5P+hryUh1TbXsL+xbhIc1Yb4LsjbX/fJf42qePSgkWhiBsR67vE9j++bRqoSe3IEoTWvwgN2OdCi
Idpi67gPhbWaC2YhjtZRfbexc37PzEmNwEelqewtUnOaI+wAHhTxhX40ukmH6XFAaGASSIIBp2MN
FbTRn8OZqfr9Tc6vx4rV89aur0rJxgwkrm8kDK6TpS4vGSc4NR7vqP8jj0brj9qID0v4SHm9yrRX
Xho4LL4ZQCBF3Be0q21n1+9i2vifEXHN3tJ69zQuiJiJaRgwgqNm140GQtJwX0ehDbFqk73FTx0+
AfXnsFYQFJwQvoRmvbuQOUaYmdg/4P4cSBjD6vNq5qktMrFyIlknHWVtC+VSO3rMZFc9ljF3YLXC
g/jJZJeGSv2L1O6Jsdk4rIbmMMNmL1huo10fcBWC/myOgWqsbZzO2hot6B/fldK0y0kCXvflLTvS
aWwp1R3WM12U3R1lT22vlDTGQWigQcQNOzwoTWGWuBp0Il08Lfu7O8ECncwjQJEmlkfM+/V9+/mU
3yt/Kqhdyn7EpBGEdbp/1dvJj2EPikX7br+1Gcm4GbPcsNFXRYUIQqTmVgICEjttbks918X7J7ci
a5dIC/3CKbEeSq9ZTrKwIq/b4lohTdfHyNgr/18/oSxhKGFdCTNusUQN7gsOl2bhzK1IMHyfKdmm
3FfKgdfqGwsBD3wGsebja4NOw5ylx5qpD8YV2MFZGdCfTA7gv2tOZfGBT0paU362gAyymqpREPKN
0rPuCxSiaPxH69TBWoOoq3/lE+PkYH8dMQOdVys9q0gC6YsjTxcYKJ1hKUJw27h2fnrDiB0pX/6z
14xmRYSSZGcvsKZwxHeGhFNaNcnOnhlbn9V5IR6uBv9LJQZ16ooMtSoz8JIcj/MxoBSpa1bfExHO
tWj8cENknCnTNNan3n3uJlA0rbfOSMQXMmVNSlH4yECjtlc6I1T9jAb4SBhiUhqjdW6ccYFFgBvI
sf0yRKySk3VpwhjNiqsHgsA8GKyXyBDByhwkUfGCiPEXIe+IwDQwoOQ4jH2F9Rq0N47R1ZqnKa/J
KudhKeSayjMX5iy+IPvUvm7EwR8gelS10s7u3hVzU5AONcMlCl1aKA0/5E57k0B6CLbIwojIisGD
aH2mEVQKYOFIpEdO0ztleQ8QTeM2IPj3a0O3X7Ch7TgQYGnyh+KrbIf63tnjdEUk/HHRmXdpyjdK
IpskN5CbNpDXnidYTYnS0hn0CoqImEEkTc7gKZdEs/58Wc34HtCzZrD2by5hpF7PSTdwa3tqoquZ
Q+MzMycfIxzGedqzQ+yud1yfbRnQzzGO/eZRFBmJi5H82R5qWE3gv+5DRtCRUZiaizKzeRlt+Jd7
u9J5S8YBxGN5WpbCHSV43vVeoiIOuI6U2AOXK2plh8pRvQCt8zegPxAOi7GnxL8urdaGF++Uz2sU
ITgxlKPSf0LBBeOSBmiXCm45gpNsPvhBWKdN4VrQnegbRhteMw7HOr75bUCK4Udk5BjdQCslkFmb
9KoSZjFJGofH2S3R7lqxtFG8slOnZ21DQSVhLiay8yRWYcU8wjj7heDSdxswjQSsuALTvzhwwBZy
nRBHgaBmxOiKfZ1z5B0gL9dgQofHWG5hvTZd0emFW+sk64Gmcti9MYyqGfMCpFZuZ6nXqN4apNk9
/oiFaGMmZ2GC55zZc2oGtRnEA9kU1AVjsoz4Fs26pQU+AM1xb6HxIFasVtGI73pePcuPYAWaRB7H
HUiS8Ke7dRtcbN8VB9UusIfh7uMBDj9BBxAR7pDY29QwWD0LFqgccjE7EH77cpvdQm5NfeIcqzox
FsTjJG7DtiNy0VMv+SODECH1FWodxq1un6tTQjbNw++++gG1h2I9tUyGQvLuZoxlfhHq0oOekomg
PnIR6KHI6VNMRLM7OTo4RtoQetEkSSy76dT0vl/aBA9v3r1W8AsQ6/yyWjfRO/mAjCFSSXU+cggP
hB68ItGyAKKmMMPdKOsxWIUrdKj7NFI5KklkbgYeoaV1IUacN0qPIWRdGgeVCfzdUOPUfgzFvgN0
UJrAHk1w8Cb9wVM+KFJC8aA2Bndk231RdWQBMvgZUUeUMDgn5rmVZyyriA+623N4iF1vyl+0vjEn
b6FdnRkS6hBBB7MO2TaINYNEOPNId98FWy4/n6VCIN+oD77D7GdUGsRr92bOGt1Y9rd8TE6AiM8w
95KS7GcxTWdYKB9l7Mph2boz2Uh3ym5FGzdC9cqkRmps2y1OkgyF3tb5xtFZp+MeDMTmweC3TP1+
nv4sHg0JAM1AJZ2DG01+VpPuW+Zjx0OtECIYik9kMOc5ViHK34BD3Br+jTd6vJod4ZlDJInjluBC
rnQMgfTF7xp5FnC11GX/mNyh7OW8civod5vH9x07efDo0ChCQuZKzYKukKW1w9L7Z58Rj0JbaMtG
mFiR5Rn44VoWcOt24BF7rqrsm7FvRGJCwI65l2kyTkALp2n9JlB3LgAbVR81L0dcWT5WXM+0ZgV0
3jOg8LGXUOQ2M3z2bGPLLOo+1HFAEooERSlsc/BvORkz9wJC5u+J9ZDOs+Io4x6TEIryNuQeKP2d
NVsZoarBkdVEl2AHF7ZMmCxvNYDfNjARsFZ2xWtnxrMMMFO8kQMKj/atwjl8PQQDA6SkdN+V3U9I
N3HaxXYYkBa4uUJTlqPzCy9O3F98LTfp1UrScwE41I5ZJrj36DJkGs7tYvmGU/KofPNKFRtkJ196
qwilbIo5BO9yPFeRKt/nD3lTe86CL4FoGFxS7kOkBilxUGxaO6nHxa9C0kjxJ4YyASCoNo5FiaGW
XTDAFjdX/94SIOb+qDuVcb+hDafYe+nNf/y9HKM3BXhdm3JyaJlG/10/WWg3kMjD1q/YAaa/GE5T
sGHiGaZImVmgRKR5StdZMC97R2+LYoamUHRJVCGlc/ca4IOOQVNlIBNQeycp3XK++36x8uEURllM
KXetJnZAvez5bW89k1ccV2gq3PNYiZ2ffCjT6FgYnGApUanARvS1d2s5dU2+2SKlbwLs9gjd1fty
3IdXZMrM97fk+yJvX8zsRNBFMUOHbpllEcYPSnnatIZoaIR4j/alaPjEVfp1VGQPVy/mYPjgTBRe
SiriQL2cytKp63k7Y4fJaeSSfEHhoQdfRE05lc8hjRz5EQqPr5CPmjqMqXRIIkLH4LxHlkY513dw
RDTWE07xSL0FQjMPJRdUqdARS+pVlRmSH/0G+0Li8kmZYzjuKjonDvkWbmx1Bir3OzM3uML6MVff
31Piqvo+HQ0txYW2DFinsMpkDGbnI++cbdJlHSqODJbParP6t4rXFQvfGhpkQsLRhfsP5dxhXz+R
ATJBQAL/d5RlrBdMT8s5AWYNxG2AK1rdqXeLGbsXuZY317idtuNncJPTN6zCziB/gQEJuAberqIs
FI51d6zCRd/KqRIpaY1t8PZ9ntQqVZkRGUCQJuhyYavxlY2OCWA7j4EemOiliMU+9PHx15ReH32j
EAPeUk3a7Oy5oHyVGM0r3pmSlaXICtkKkNeR05ngSK4FqrragsxcmGE7ZLVYg5kJZns3rtR56Zdz
bMwE4vkvoOGebFael4ec0dXSdMemUGpiKHDO27irJicP2OI9zYtLKkLVEjSM4BoW/plJAFc79dMB
66HMuTsrSQNBTEqzhaQE1e+kheou7qnzZq3GblN9YYD5XLMocPF5Pwc5wKm+/9IPN2ivo7KDxTsF
1IRKZY2FJdIgiLvf6SJT0cf9qkQtDraQXInfrQpf7HDtTjTRsb4RZ2h3avGY92WZgwa/mfLFQxku
CN+rElhJEY6HVwomOZinsaIue3GwWt/CZkCJLZ31QTic0RU8r9m/jsYTPiFbc3tDHco0g7OZIEO9
Mn1mBuTd4GpqpvDFr/YtLV48AGd0SSktPWxEXZtNgMBwvlnXb+0PwEaTaoA8td1CPS0KLDGVSCJH
+Go69TcmSeYUr88SAN9hhrktzv563+qS7aiuQoe3ViGUqse5tq+PE/OETSe099aTUa+5uflnXhaL
crquEI1UfIN00p4gXEI5l5okn5Scz5R8RHJTCM4hjeC9mxH9D/7ksNm7JQbAmj0qBmUaeXYOdgc2
MakIm4tWIzM4KxcbANLkYYNf1njcZ1XXe3UwwUfcew9R7HouBsEfPUZKPnJlBf79jHW2orNWwgFw
xdXYuCUHlpvEwTMETc1nAB0b76H9p5zPovWb0ozY6uX6Q2wfeaMGWaKEh/ocfSFCI2JYKRzNFuv0
SFanYZeP0TGmITgrXYvimKEmj/LGxm3VSdaIPuW9yYkF8XbVo5L8U4mQt64D5PvcEP0zEVwk61cb
TQwsa5YiI928nzsyx5nG20OMSd/nRaqDeN+F109l8Q8qOfmiQkzOoq2OodD59RSxFuIjAGyvGBNQ
9lApBNB8cJSeEds5r28ulFLN7aCU2dn8+rIfyORq1t5PbCkgyajXOuAT62SD7lFjjoCOlLJnxn1W
Gx6+uDCr4b1CHEVfVwU3r1iaDetyAXFDvHcuM4KIJ0FVA5VhxQaR+LcmRmCI54IlwAThEUcB1onr
tUfRJrz0T+aONwkGfDH68RD3XLD+oemG8zMUYQDvUQJzdO8uKUoGCqT974B8sV2d07fxYTRfHKar
dF8wEJTQFsgum5ZP6b4CpYnY97tBBZYwtsaLUchaC9J7kYAAX3/ENaY5ceCykF5cql7xaF9/wtAW
sIlJhNnpvgzDAURDYoGFx49HaJvgUNd7/s9U6+5cgdNdNF2qbBP9HZwdm2B0jTB3MLJwiKqLd4Iy
7+R0ALiwi5J2cnpDxoTfmRZjHVLsCbcCWuV9J7xdmHoJrAU1imYTA7M+YpGhiQic4HNwopZVwScD
r+JyUnV6mC4GjvTlPvOP1aeZb17A9EQnJCuHYPZJG14f5gxlO7/mer0a2MDFn6eOnfSidmnZbuJ1
173H8uY2kuhjJfA6YTwCNlsd0f8jX3lQVVLXkdTd1vLx+djNcayDyqDS3EXnL1K7/LYEvgf6tjJG
dKkwJZxSmMIYbLmburBO8x+JvcDxQCXd+p3Qvb9se0twBUU/cHRcT0DAyWqQQ2KoUytcNS/3zSap
P9g4OeXfiRbCTbmxECfoJj5sanAVhA3wNdQb71MS0Xe4Gjxpl8ABBUXJZm4CV9Yd5B6UtcS24t3r
SLbg+DRmnyHcVJJ3pnzOZHRcNBM8f0uHWJxET/3zKrHtsUpVsbCI1SPgun7RAGw8K8lNo+qxfMSL
mLpGokc1YX2FXGKIug3+ppD4R+fqgpO1QNgTsIJ48hgwTRummcpxQVvKIV0QVFLF7D5mvbf6B3gl
C1PWNTRNJ+9kyZegbvHQ9xDPDF+BJt31g5ycOGTdS5M4XluhTOhjz2LdFaR4D9tNNndSPmTTQaT9
sfmOJthlwaSBDHAb4M9bjagh7EE4aqamO5h3cCetYT4bQAWbnLgKlJSB86ocmN6/+dGH1QVLcBdu
zagtOus0TW0pHWZLDdPdZYZjNGMUxM8kCjCY4Bw7n3xQiMT1SglrcZp1+EgjwXAIg5DejpClroab
lEZsgyOk46mnvpeL7gDkHbHDARXDuCmnyCVZAoM3vRtu41fsbNYGc03ofveSIbxTTrFYDuAy30Xc
UCTTva87qbOfFP50e2OAeM9SnbigzS0PlogbQ/0JvCz0KkWFR7o87wlvaToM1T1MkF6J2HNpkxlP
sGjG4wVu8aR2GEaYEj/JQ8P4KSCi96jzNj+rkn2FVvBVXtZs1V3z09tHRc8dltaFhgmQzwQThaQA
FZY2kWgAJNZZ8pgC7v8T/lSIJNAUQ9usVVHq+LsqlDjn19VYlP3pcbOnsq9x5aS1R3ZCk1QtY7av
cnujQikkkwss+qAf17xbGfzqgDK61hBtwbUDFuM0dDGocFE6lzfDK2MrxSN6RYA937w98w8i06Q8
fPBpPcTX1ApYVEFFfOV/5H7oWJDrwebzkVCDnXzY6QEtY+m2gJu30RhsC4FEO0GxmPqOw6jOpVWK
0eHGIv6aY/HyJkwhAf02VaGa9DXkb69+1FRqR6Zgae44WnB5mn+IOueLu+mjmJrG9oPhDqZSw5bM
KYzSUnrEWM9Y2+UbFpdIpXrvz7ozI7ckU1BuLuapbvV7izudUmqB6xHiPqS4HG0K5plol4cQcQ4A
H2e0mhCu5CHID9yRTaB0rVgK2SIBh2PxtYZv/ebY/dTkaem5IjvfCC/sHu1xXig6QAkw4AKRZxxe
hq35tbs/P4BsHFtEakXOV55MPVtoao4qS9suAFmQXEaEquMbcJRSzf+B7DtBVgLkGpz4glq+3UY6
gsm6CjUTv07u7Pb0aSc4OKfYeqp2n8awqpdFLBBUjgTmGaFSraz/daf+Wuf6OVm3KgMykfU5vXC5
y0fUTaQChXwLu8n3NgheE0qgt2GhfR0qHHldFJJ2feXwmUCdVsmRW82zCm5XZoGaECqyXI0ngnVN
xUwlrP4ncFLDQxgeLo1V1X6LnbxZLtpfw6b7U7Wh5a946p6/Z3s+aWqq8YlIarTh65Ag1ff0X0OY
ELkfBs/YDfjSpImjqS5z+uS30ByIJB09pu9ei+/IeZCQQCsKOLD/i3a8S0pXryuMoEWIdnsaDW5B
yg0ojT8ZzE7jlsiqaEkDwbXEf4G7pcobcFqY56tfN3otXvtFYvJZGqvPcIMbyPf1sNfzCd35wldB
x8t4PEpJvpU8u5v8pJu80KBgaX/57P17xYTPrVMOu1Y0fBiE/StsiAu25VafA8VDv9qsWx+ZJdmx
Edqzn+8cfAF303zO/dsxfGKO9EojYseF35t9bffu/n+x/wVQ3VdBvpzI9c1iwPiqpM7LddIebJ5g
s5HXoW1XTes4cJRPmvINDUe4o4Syqrlf/+B+yDGB98lSZTOmj9f543pgd1vlMQI43/vk3KfKfDlA
9DmANR6GRcCr4LqlB8aSPdMd93FZLbvdSr1nhAP7SWiu/IUr+ROyER8osgwvgJjQLFxOHSQezYYb
+A8zyRFpzSpg8z0TfftS47jU8p39czCk13pGsmLSwJWL/pN/QAbtskT1wq1ygt7v7mSsK60oIGzG
gV3I0vY2mPxsoLULrnJLXmgei4UOMmlFOQZzkM29zJGBvEOicgxYEaoHjirF+lmaS70QmeNvToHe
3LYJ6mAC8g29wSQB0iR0VZJv34/GqpOoLrqB8kdgrlVJ0jQAZFlJEQ/g7Qzjy0YlxXpNRLNeDqxl
hJ1Sq2cySafau2WJaKuBYRkCfyufMWrIGdzr6saQc4RDojqor9lSiz4mE370mIFFYYTsqUzN+2Wo
qXarvnb1A6kyvBXLNfOO/iyh+lWY/FL1teeOAci7m+Cgtmoo7hjO1omznbV9yp4YoEMT5L12vc03
VmaEINpAQgakpuO4rUAsccfF/WeFLE68beeVeSfqNYhfxksZass7vmLn0+C6nCOZObyfbVk9AqeH
M68ImSvXjV/8ZZc7reTRASr6ZREpM2GbH68Dkrj7oT8dMxImHCD74P4+fZbQLGlh6jxwyYVSjgMM
KqcZlsu8S8k/MMSvI1i68rzXWWaSrq/KX467sKSuCbZCNhSXNRqXQ4VrYp0YLt8NX3okYZhyywpL
zcL6bLgBsNVoSaueC/Hdi7ri2baH4KC8Kj3igZ4fRfmtdQ1jxyeH+DuRDJacMXMzMtpGxff+7NqK
neij7dUULLwZzUd7keLXtPuZ9zbC6r3bazrGnXL+8Eb6lCQV+qlJEzhMaBqQAFlKD2tjrkKc8r1u
JPzhiaj3wrw2Og1cD9Ne8BOrgtHbKaUq+iGAj1SXJIafXSX7GwUgpUU4r66PI9IbCDkegGQWA4hp
QFGrdll/t2ctU6VCTToK4xdcxGNri+8ihK7sgbwkals4EfHQdwrK89TxBlJudURImR8UPnGBe0YN
zD9z/mmW0/KkPr/64vE8sWXNrG04zPUMvLdEDoTm1gnszeyb6WXlf0DnbqzpJdKnF+DD3ngSC79y
s9ZzK+++Rs74hZdG/bHNtoL5fWNaZtAvMnjIKURA/YuDW1sqhiXtESKSipa/40kDzytZn1lekpM8
TO9XLgoaKKmriw7K4LaAZNXCTJYbiAAi6b2wRi430zjAF8TRJntaRfmXPl4OIMJYE/C6GRUukLot
+IYIItgTyPcnGbGM72b6Jok1d922bwsdcC2eRkdlNVcfGLl0U/E8CxUAgWE8+dmicfGzpI73NJMV
NL3zmz8WboREbXXS7pCeEhQaNiVQ0vz3jtXFEKwiHQxcLihHJQn0LWJFN1WfHrI7CzeYf9VMvo1M
AAllwrh3yJHLZFFk4int54nUotr02VjT12VJxSmZeXC24DW+44QX0jo6vsMmBbpMACWm92iyAr3T
YIt1cCg42CPdIQFdNInWyxeufLSAiqq2AFtn8j0Iut8tNSeheDi/TCyGiypdi7kAQ+fQ0kz053OJ
rpeJ8WiRnsgwXiGhvs02Keu8YXNSpCaGYyqhHMQOnHhbbQW5lyXbjICuvEqe6jZyJEXI1DAVjc/Z
yJCDOW4WC3MAfkZjqCg+diMnf+zseXeee7Oqclb8pQVMggZi8kKxskAguRhELp3k4tki8SGR0YE+
7efVaeC7WBUJMpQJJOjCrPMSqcuXTHxiRDKKBsVo+opP/lYQpQb7DaY0dWInrVVnJUdwUYbhBueo
EgmtiwkiTViLlkPK+uczhJMy+epnvq0VVhZ3nPtwLAHrr6QIfeWRBT9Q6P9J2IQDVvVazeocH1Eg
YVvGv1W84Cm7g8PYDe8zs38hWetjGEq4LzL4QFNRtMYFP3eMB50Vk5XDbZhDOHYBzalnT0YwF6W5
kl0+TxI+FPgNTAbNm+37L7JqWIEeXO1jqaRy8k6uIX1toLl6PrQTowZFhXZIPNKfVx1bZxbK8t1+
bnJkZ+yl3CwTAEED+5kIzAyUHp9xBy/Hx63VRuphn/vdaHMqqQQ4WkcSlg8lktutfx/Awz0lfOHF
iofYb23qA27scl+Pl8eBQ7UNGzotO3h7Qw4o6Y5c05Fnc1y+xU7+jMmumC2YoRjdLav9xbH55wwa
JnaeE1CFDuefCv8F/1uDFd+ITZf1x1wN0HOH8HA/dItteqbcbbayflRB0IOoED1/LKT/xiby6r+z
+g4LCF0+c4f2m8eGxF4HnVsjZolAI2kDwnTS4preI4tPq9O1ANMRQGOuoEY7e5CVRFtRk1psXHQt
72UPh8wKHH06pX0GJFJz6BJTguPJHaQJgLJ6/5Z9A7Tq7IFNqjR3S8kAFB4S9GU/Vq8VkXPRyMVq
zrIjZjj/apOcFEV9pSv7i6DZX8+uNJy0sLe/5mMNKUK9SmQFE8Kmf0WkC7qIELxiLNMY/Vl2Gj11
wau/JIUY5H3uIASlW0W0BaiuBfTSFMe+vj8JX4uH7kGNc65LimC4tq9pSn3dashd/+jOdDcG5h0c
9mekDaEBeYUnYmu8HbMoRn/rZzQau0+t6wUHY/d/pXVfY5cwhVjceEzfHT1XwKZxnvHfoiZZP8Sf
oFiMjksxFaXE93IQ3dDhfCNYkKGmqUI25S9abE+r6GS5oqkDZGsZFoQBonqE1In/Twey1De4j4wq
yh+DTHhNC/1WnxkRReyZcyBgjbcqCOc8i8VTpN4b+dGYGP6sp3RRu/SYok/Vu+bMW8RJ4n4h7IFG
cjJZEgI3EXm1KxCB4Vc/vq8cMLwad8i0CGFptk4nvwCCSm7W2yInPK6Zvgpcs1+oYjtaORimrxLQ
6kULJl319uVfym9MlVeRWUrruK7kvyxAa5HjlUohp65+s++3jssdTkkrXuS/yAOdGS6gDEHutti3
PODu9LeJVWVwLfKzfpYoSXKGumidismhez80A+gPdwbI2plynkYRYKws932VBdR7hFxSuAjfJqnU
DcQ2+ymKlv6ahZCM34qnHUpF5MIRNJx7nYSxBPJ0T1hleaycG1jC5YA9ffLhhtnZEjomz9n76gbK
cNBLD91DGYP8WS3YgPu2+2pFX33h18JxtRPrTDO0jlm32jbS8XW4v7vI81YPaarxnNSkF/EwK3Dm
2J9Bb+0DHCTXobe+gnd3i2PpmyrM4ZIlx4F+93HtVMBulpGbcxfGAPYc4Lg5Q/uzQLYhC/f5atOC
sffmUR2T8JoLMO6Tr8VpYw7Whnl0q3r6e/jzkKKj8oQiTc5PHACevbZeuGubb+uNRxum3vcg05q8
FIXh+I1LWHKmzNfJYRZk83GqDUT63uPTTNBnBrJiIc20jzwXx9Qpwbj2Nfxa7UQs+EgmuQqZrraw
GQU7n73QT5xiN+O2VWgr3cThlU31+HKv7MivVhtzW2AurfKNG/WvTEYYsf3FLf+XL4zUDH9Vpje9
DmhZ2/h2YaHcnjFOEtY+Sxx75Npdwxi0a9oIo7k77JvBN3Y3i+AdRiGvjgA/Kek3unSZLD/kh0fO
G1jWFc9cUD6GrAOI5aX+UiqOOg0MM0rGx6EL+IpeX7HR2f0q0MhR0c61ChaIAjJ2xs1Q8WO3jQc4
qFYJOV6/3SZImRdMuH5ptLbVNwoMfqqxVqb32nvfMHiBr+uDrNiGjo6jsidxqwFTKDwRM4lyitkC
iKgXik6bWu4VzNWVJuD6yKnSO1cfn+Ivb5eTrPKy0aZZXIXdrKTFDPmrXB8Nsi53cPhKhCOpv5ds
I8hh5yhAg4kxwfhX+llg+b9Tma/mXadDdcnONK/ZB/vSAFoyaIf9e7KPeuR7GjEdqdoOLsm5yKw2
gQhZDCumPghr0T5GytlFVZuZ3tRoLzFdvjq30GGC26JeeKMeXean8F0VQJKaibWhSdNHYwVpQld3
jVgHkt/Ro8yU2HTY0Ax/FJrJP3n/zjWVcVNxG3zU4Jek56z/3sWqERxI9kldriizAMFhTdtxY4/S
oXYFcqxCtEGXLUIewzc2pwOH6J8jtTFbdkD7qiKW5HU+edZigX6HwIaTxuc1PGrS/QSyWArykFRa
WzHtfgOoQhaJXaFVsOZfm01WXiiR/Pr6R0eDJskigo/QBejJhcVODRYwAdKjiYlvSEeB8lDcD8I/
f9sUWgKHtIS/ab50tcR6HnBDdBrETqg5d32SfynOtFIKBtOwLVa6zU7GoyHIjMydq7JodKx+ZSCp
MsA/TugG9+4rOZAex6ywRINUWfBxb5MfpDv9z61KKLKpYQ3yAGZvevTM6wd2IzYppQscD0EuNMW2
JbySx7JkR/8aO9PzSLSi/3bDhi0e+AoFvuwlC5g0FG152dLDgwtRdDyjRJY3TNlu+dLR9Q7rRh87
OSTR9GqYfgTLB/IY9qAbU3vIv6VA0OC8ccoslaEf+Cqg4+YHFPPw+dDbH4Qjnpn+UeKWAE1OzxT9
ji65bDg4ePWUTQ4dSt6zciwSIKRslAN/GZ0CvHDHc9rc2gMhvE1r2WRnAsedjrDoR4WZd4/HXRkb
BtIDj+LLD12Iomh8AotqEUxtx+sdj2txWnnHzL8QmQrRjgbRp5KOxA3n3PGZKNK8CexlM4GoiC+o
8+aduzOLq+Y7I+bMgyS62eiQ/r2woXTOzsu4uh5LSoVtZouVH8BClQHccGr5bq3OWloHjB2UfR49
J3Q6NMpFcGNNDtxcj8YzKW0PifT/JRLuLt3+56Xcv6Tx+8p5BQ34u1RE9nqe/g/7rRVhshgkLqu/
WUA8RVuOQOUDqCE1IrX2qUNmyz4DCvPI63ny0pOAEjjQftqDS7RWYGMN5wiRmt9BsircTdbS7ATT
M14v+adR+7zX6zwbPitivMt+zB0AqR80azUbghUlGb3pG0Pcy6UWR6aaMnkgk7hGMqvVwjL7/hxL
q254tmeQDwaCm21vHxQQu/RxQeDdt56bs9SMJQ7X5O/GH3qIrE9NDmGgrpUgBhR3aNGpqJHQ6L0X
rukbznmFFwx7Jvsq1drPsusnBJluVAiKCmKCY+30Wk+Deb25nILzQShmV7Km23jWaTLb9sjuUb64
yz1y59lHGqpKHYEt4Plma8rw+Y3jYxX8QAqtM9eVgE5r16Kfz860FGySAlJRyfft9aagN3uXBctu
ATN4r81HIkAt8o9Tm9gBsHskHSV+EvRhsmUfXcV8729dA8lADmqtZ44j000i3m1qqly8JtExq7GP
tddGKFo5xNvSC+7d+5apiGsNckJ4UxBw4s4ekZYKQHgkjLWR13rsBzOgrZoi/CClRCgqLfWxGOPo
4zDe1l+WNGBaZ0Us2fzJXeFX2w9SeXeqdwzN3MFB7BO8eSmAQqIKYdV6YS4eG9a4Xj4gpjJXd/96
50QCV7LyI3dwAnY41gOg3I+p3/gBYyN8t5PnLiWvScnynEHm34bK25AMICRRjV4sNPsPBdc5vbDq
PCiyKx8fzKdTYwVUu3iEcE33Ae46/Jga96q1KHF6cTsMKZ692KhNc9ug1TGloXrbWBu0Uu8C22hI
uF8oyMumuwo4tA7SZYEXKIuZdOkHfHFymIRzUBGplSq3wLZ8DEDIc4YRGIPCdvEAsJCNf6ZvY5mv
OReEIZAjXTwhSbQFnkoyc4C9Vph9gS0p6F/m6WbJiTGsJpwJU9BEMC0FPt6y2xTzshBSzSwiEeR+
j21/Vs8LBWj+TqTgMkzxMyV7q0b4ekuAyxfKFTOh7JSDQNVaq0WIq2Z8/Eqbxh1cRIeSqthX85DQ
b1tB2SYZnrlMjXyvrXY2NTK/ih/TCvhQZ2W9WKplWm7YJ6J47PRLTrS2gkQH5y5co8GyGC4/+Hqt
dChdKJf9mAE+zBNge91VjKOkn/6023kgbvGBmmnZDzC8+B1Gk0Pw0RjTZ6D2cdp3eeUSRVfuhj5T
rVjPPiSxEG32CeoCoLVS+vd9lx1KSK7tcuEpwBrkRtXq6Y4XcmyFF93ua6Xc94S8wHZsq+Ec13Fg
cq0TrJA/d+FLWjpAogLJPbQ8z80MMJZbgik4mRq1czBwiilEtOsrnhb1Zg/D6TG1Y0bG4tCQmiwA
fwjX8/DTc2tQNE3/Uyw2T0+l3iGGlZeeMTIIqUKNagNo7PmApnkiWzGVE0Y9B+9iOQyuwnwtS8EJ
Uz1wEmTmKvUCS1imKGPqsKiHx8u6y6irLFIJNz03J4JnQ0NqkeHXOGQDbao2OUKduHqcsZjwwwrC
l0N7W+XXvZlf5mZqlvkyW0dEBaWEIrC1nH94JAMsF7zWMJGaniFRhTnPhm+Lcu0R/4fqBl0f2Drn
0f0r3BTOx43/k6v3hyArGgcJgnU8ET2ooSZJrj1Y2+nBYF2oPtBvfu/uvwwgpj92g4SczZB//Fjb
OeCVp2j7et8ooXtQZRUhSe/yFs0epZT6CWJz/VWEyW0RYSwz+SRS9yDlvVJWOZMUu3kVwpfV0xQR
4/29pAYrdYvS5nFSX832IGsHqYmbTTV/oamrC/LiF+WiiCSSNu9JIZkCAPxZMqUMhurWFp+VfBto
SqpoBfs+4PIgVI3QXfArRS4QlIVl+e2gc2rOSOfPaBs0sXFu47RluVzmFhipYri3rNfxxOPbGJGN
O1dS1hR700fltIQscLzzCA4cl5IBxlrnqAJVlfTXW7snyySA3vEGD0HNYxXeaCyHxM9tzrGywMdU
+Yz3Dw9wIXFBUBPcrQXHckTkZQey2IUKAb6mFjKrm8GuVPM5OiS6/FlaAa8agC/DQzrRvfA+8nMO
TCzvBleYQiJFfonuuRP/NNfkAyLvxqLNpD0woLPxDtpPS4P+Dp7ZyKDgxcclOQDSwWeZgGhQPu/X
uhMxMmDlurHSqf2i9L+o2kmCcANbIO9r9cBDhzo4naAU45+efI+IRB1Z0GJwOv98cB44RIX2HqaN
kK00xkH0W4/eoYpuvHE0HJw+qSQwDoV/D2gbDLFZIYyoJ4aDP5jV+YDcEp4Jhp8WGYeSAcXc1TxH
hjb2uhyigu4LX2nA1DJefkIVZUktwWdIgLUr+dOIBXe+omLt3IL1D+ZdGJLmdHuzAmvgPc9bVUNB
Xxvevsh5ZoGSAVeRw5gfDvxDc/NX0G5fsAWgfSVqmuP65AXQEgGxmLvn1gGUkz44KXNCwciWOWth
mu/0IQmG/bjpXHbgZm5B9nL0p4Ya8c7yb37k8GoYs/HkzZhj+EDhEOoa/uUNzuipzQjFBYZVtG87
+s2z6OoTZOnNfTO2RVK86zJJvPKl+FhtAKrtLfY7Fc7mAlmgal8E7lvT2gmBcr93+tkELrAzSI0L
1bHWM9tu79zw5yuIyx65MqMEQGz0+Dod+/fN0yXlarwnWhCyeX9EXgQQ25bDxm/ne7mBWiX06abg
lBSSi3E9AtThVMy2oax7XzZfIDJvviP+panAXY+6vkPwvdG9Swffqf9MhI8a/SL0MTiZixHL1B85
rnHuO/rEm1Fa9EtD51LVJJy6Y8tBaKM00IIb57U25sldf/GlXfCmA8dMwFK+DZ2Om/lBX/DCEep8
pJj7FRp3Q4Eq+9Cu8OVXUxFgeplmKm2jRjzgs7Ox7LxxbFV40kLIQkowT8oLKg9V9N3frpe3tGpV
fXe3U+p91ds6PRzg2EOVJ5Kypw3BZfuBk3Z6QZXwN9dk2ROqywZ1v6/XnzgthCIRQQ7pAdhgzKX0
sKaaM2ZRCW5JLmmZbQg9ueYk2v/XouZzANzKljzYLNmNndbM0g/SS4QkwyaBXmSsMDCB10826425
lIagnfyZK2ck9pcOHuLgz2vb5TBa1r+mWjFLLwyff9oukzaJINqZr4nR0njDZgZatFm4HFVWH7f2
tOb0OA1O6QVTZdpbSnQ9pHyMI+8K25+sIBNKmu9mIl2GnSkfmJ+zUTBBJ8AM1QhjeRoiULvt7U6R
Ar8FmC5eaY900h9yhSDXNSjcH0A33QlZSLovh7pf+otf8dxjw8YOBlH7o6emZgDGs61GQ46XkRog
FQHgKEuGgCJeQ1bg5idWsX/7NbxALxlrcDyNJE0eODT4MQCA2UV9GK6OK/su8h9VqwaIPKcJVZGq
/iRS0htDMbS80n0G7lEtAt63hmQdKfeRp+6O59Z+6wn9pjck9WJlsk9pksvE5fNVbxaM6wk+DIkC
kbu5JggHEr7yIj6aARWcY4y9oi4mc2QVenHSm/WYSvjNZejdnTdYT1n+wmICN1Vs4s1lMH/cvGDW
N1MRJGSlOnAavRb0mye4ITM8Buj06+QScld0labO02+ZNvfB+vZGhh8phrP/wnEk7YOLncpxcY/c
lLIlw1OUsiyODRG+YdXYX71hl007j7K5tup3kYAjLoheGgPxROc4kW4SubuPURzIJuiSgwAltElu
HqZzW3NJUXX2C2l0gb5cq6unWAwr4YXymftHONB1EbiM4h7gMmfLiYcvV5vrArrPLaQ4A8tsJvFf
TGQezAS0Qy7g257Gu7VupH7JTREkmhlQf8/gNbnxcrQkTQoPzP6iaVIXpqQzzuHefj/9V+y6BfI6
x/FsLrOEN+C2eme3jjG6tLcnYaxvuu91IniAnTPfxZGLx1i6O/g78KOyaym8MRS2UC8XA3wyKDrY
4nVT70Dyh6PqUkMBMCAIa9VlSSFASe1t0BU/hrDcMCidjsJuZeZMEfbzeN/Tqb/It0xs2bG8dhIR
5WMYGsKVvId29PzcNFSFUZb9oQcikhKUJQhfvTw5Exxka7Ks4v8+/QfxZZcznKDWnzSw8KTr1mYT
Zm+mpsek4LdW8cdzv4HKL8QKr3XoNX1sNWzzB5+DX8DHvlPV1/8SAlcQVdmgDnAE4OQ56zTKWkcF
9ramefr4ItNpDwhRv3cjCfcwwZdCYPoZXZbbd2+/uzKMVeGM/NWvMoOP3H2hF9dLEBa2ROFsFUio
hwWhdX1Giekytpgt08nEqm7qm8sbDQ6DBg4EAnmr8mGhlQBn7vNNGsg/F2nlFVDvW54RX6zhqPxL
p9YKbmwktpI1eJ1lZguupv5P1cQlp98RYZBEnOE9AWQPlm1gYd71uj2+yphNT2mkl/qeh2dpRvDM
Z0wfH+AlI4DYMq2P8xdOYi9+bufQ7H+ugJnjYyQwj5ur2uTBBelCR+bvXl3HaAKtK5TE43BhTeWU
NYttrJ18timceMTaJVoY4XglOcQxk/6zyAtWMNDOG50xFeL3oZtEFXFiNct7i2eeA9WNuny4X7XC
eOQZAL4MbMt16Uud61g7sF/bIuypvLQmT+Hl+H4ureaDLzufT/bFid75GwRIneR+uZTIMhgY3suh
IwNkJniA7OcQR8/6DMKOTqb28e4oyBB0WW0QQwf7DrNJOXKxJJR0N4YG8Qsj/6SA0G91nMWY1gZ0
1bgwVCnA6EEWuh6+cOem7s8es1exN6CBitlZUiYtlqW+mN5AwrDShzFu46n8SKa3tByrF/zklzb9
IrRwQSdEjBHKP4NOTcdDRpiu8QNN
`pragma protect end_protected
