// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
qbDtF2BEqWYhltqQ9GlXxF1+0sa8Q0sd4Dxf+cFrI8FJqLvXa6+bQI2TkVw29iC+CyZUeXYnqofM
45YDPnOrrrBJAqNaced5FkjZ1P80aAXOaxyG323whDmLBZQBxWfYYo8q0xI8HAtt16iUBuI5iIY8
d7p9WrtOWxvUIodo7bodrF+iKVfN4JIxyno/C+b5B/krPPtL2D2wZcw3Zu9BLCqe7DRMPj0tqXy7
7cqVUDYOuezL1NQhd/M71LLI41SAef60PAAsrRvP0EfXdw2TWFqKM6ISESzlCjpc4m85eeVSePRt
dS/j5sBUIIHCTfaI2XTezBZ8AcK3X8gZiq8GUw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
6u4wnKZiJhcpuCFHFH+1LmM/f2yVHDgTjrJIuih6smwqVsHHKlRP5DBckdbgG5QjKZ31G3WSv+ZO
ocbSu4m8DiplbwnSadjTX6/o8blIlD80WzY0zlS+w7kNyPRpDC6epgY4xBfc4fkD1Zjeq7lPYve0
BxSlBqucEWr3yoHg4KpA3UcABySYjnJ2BWBM6ki8zIWDGF2Pi/sbU9YqjSODe9YkIPG7yBAiiyWt
+I950PNfq/bVHN2otCosfIdnR/4ZvRmYAq2kssz/qN9T+PesfANP7/h3njNdHLzdWTIwkI973CbV
QrmG9k8PnOri3hYK/uJBk1YWqc6WmmbduymzoMyWgQFgs4eLBHO1bLIWqHEA3vvOOkZ4XXIBhkAX
4ayyAm9SPiEBoy6ddDBGpcBju48VO8QSqUyjRBnynQOTjNIDV82daqHHC9TE2WGlDMFA7sK04oCh
4v+m3RAgyKl0snaI79PfBOJWegjuW+MBBFF0aMCUtggbglAUNjL2pE57bdXmLAH00EAqsi0iIWoO
UQ76dNLOfTFXvEMwZynARra6YLnENsu700LMe8QWuJzcmc1UUNguPFJwMxkdlE0oK8i7QaHOHKzF
Zhpgb7d5XKVk8XPvTtkeNPgUlOvyeYP5w7RmBulYtXVKaO4GctmX3We2/DCXyHoW1n+/kcZT1o4J
rAJL3Jv3uEqNSZDyyg6ntDyf2bFc7zdzV9bwH5EB95RsiKmgQ7aB7Rh9Za2bOZzqwHAmY0zpdqRn
IipSov9Hcc+RHFKJdb6FI9//lrumi0GmAcnN8PaguAalAsylsUiF9aYQ8elRr4pa0Orns/PfceIC
e4Nh1W5Z5C/eay4TGxOUdNtOWLCLdMirqJDsn7FdfvnGsrh+peuZ8BNqad+UXUrfP8oQ2WpwT3n/
qm/ss13bQ/5i16hhU+BARFbDo3r5J1ZW1DVpkwf4pEFx+R1NMNzVplii50Cmt0RUFJx1PksS/2Er
UCE5xlwT+j2p3w4My6diIV9JjdiNEqnsCOIe6kf+tx0EvLd3NMGMpwLrXRmr8Y09yrkdpc96EzIH
uWQdxOisrNH/p2APZLVa7h6LxklVsdXJeDHptJipqz93GpqWY9OM4daj90Qq2y4BDQrSSGSLsQQS
XVtoG4wWD8Up9xg0cp+vNVfmm9PU/Se1NAXrGRErtXTRO6cZgxp/4vH1uUgQzLUC7XDPpOpvy3my
X8gwxR8EaZdYL/gRjqLpwlpTTnzuxKgF8fRETAZh+glgA8lWC+NmpH2nCqinOZrfz/Vgsan6hKp5
KpadUOmjmgat3AlVGhHi9EnzlDenX6b6G+MhEazHgVFEpENYCWfkKK0V4nV9kKcFK4WMXp29eMjJ
v4AEM5u8HPyPhPyP4+PjMgo5eTHagPxBQHLq5uY95pYpi5YbqD5LxHB0M9BfJP/wbzeznL7EoKu+
zKDam46ULabi4DJ1eRKH30caa2dqqfx2y9BCcju6o8lHD6wFyqqKrZSWzcy9MUNcpmHh8uZVsYrj
AwiwzUmkRyJkbvy6c8VJj20khMVrFUs2gPUHIAft5WY82pYHr1WBnB6aV0LqhRRVomugSpfy8iSD
Kz/eWVlnV2uj/dSei1qRtp87tqeQ3NJR/N55iIXn7xfnTAIMOgMj27waZEZxlIqNIiGu9VaPPLAs
TZAk+m+d/fNpUuXTWHYKkLRspxikm7awRmuZ8qpnQUDvvjaWD8yUGTugNkEsiPjXKOyudGqHma3r
BBbftOOP+6SctwSg8hybVOq5IHWi+yxBEpRDudMZrfU9JjJiXvy0hg+ItFGYT06NYnG3D7PuRvZ1
wCWe7KbZ7n60anIN6ckPrZrZTYwoWVU69XhYewZtusoT4uh04S40Rcqw5G5shxqfbj4YPHnA3pM1
cKfdDCCnvi4yt3cEmbbv49EJrCciWS0DcJVzCt8lzKkMria+GXFSJk0cMl1HqIC8X7urcHnwm4OT
F1N9KErppYDuOAIEA7d3RmxBgkUmcnLwySQdObVCKSGurZ47pVIFWEDB0XfXF4l5mxq3YurI9B7S
1hy/yUWUNoSw2jfwal+9N1oDLu+wlPzHTKwpVGlq6db1JfK11XtNMDdVxYb57YARsnWDpsJbuMJH
SOBOUpNAwDnrZYgJUXhBFbH0l5smqH87firIXD1YAA/N27i+7Fz+1la0dZ1lgxJ+igC8Sm0SZ7mD
R0T3dB58HY/5Dt6g/0o/wDwAr1b5qJhqIxZDKLLyIsfleK9Xo+IXSF/F2UT+EbqOswmSny2HWtAp
gMjx9+V8c8s4k8nOw6rpJhYO7IZumAEZa9L8XblGLG1CYCzGwEhLfhpO7BmrvxHY3pkpOe32n4Ub
LSVrhE1hfZjr7+cUJjE5ILQIIlj/IL6aAHFdbUc/rYkAZO5YOXoeKU0H8usOuJovluHqalOeiWXD
zHWpsXxgKQyyVCSHbSLO/fQB2JrDUAUR434bGD/AA0ILoV6rVHPAyabfsvxdLgIgOl/868usj6OP
2OToIy7z+XjS8nD3a1uLyaLbg8HcBXqdpaj2EGp0XGsfQNqS6Vi/zGW5jV+J+l+ovjefaqA0dTTc
vsBuL9pl2E83Izxa5pkyo1e9cCgzrWyTyMCMz9B16raIxg05r2IPEKBQ+hsqF7hHGV4X42XQV/61
E0u5s3pIPR9C+KfcQkNh+nIIu+1LHXDEuZbbdTRxOsu9JZ8MnApWUOnXG2DT1AQ0DIw/FzvitimX
tSRmY1JkimsuARWBsR9wqwsLIcIhcvtd4gDRxEdWAI7dSQQ01UpGnctENAzUfyolsM9e09jCNn3a
y2dt8Lxr3YbFhl5MYJgAhlvGo8V6CVAtQbFYY2lYMap6eR1ixcSv5aevtWkoOlPHMxYvZTrUl8yr
BdjKh3TEg3wkms2TYIhI+KdkPEZBIogfBZmtyC3d/KnpWJAy7ZxoMQ48TS84pfFIoWZb3jO98ITl
RRZoDAjRMeuAD6SHWHa4TeCDEqXXt6VbQ0NjTURulaXqn65vJsSuNXTszANyoOhYERqaszMfhQfR
vVP81D6OQ8teR208WsKtF6fH45xjtZt9ytYHbrcAF79CGepqfV/jo3/c1JRjCW0lurYJqhham+Ph
oPLfgwD3E9AWUCZEGEOvKcAzGhBO93i9TkaCl+YYupKaCjpRiijmahrq3fmKtMOFSX3GxfivQh08
JiE1eq8K+epHA92bgRsbIbsndC3eLUzqOOpUJvpi263pQi7W2iAVBTXaoHn/DVZZF6cD4Oe2ZC+2
ZOcPUZCJqdARFX6eqtfoPtKSkmOnKIc1nfX9Dw1Q8JwgbLWfo9gKXK34J+MA6cCuIdYp/XIV9EKE
AY6jXDzsvnU8SmG5HzuhRuXKHrAnwQctmZta4Kp5vQGHbN3M2ghWpKwKKFZyjP3Ov0mrc0W+LOSl
76+5idYhHNFRgk284qWeA4ie+R/Y9SowWrhEE4j009u2GFc8NhLCTCAp68VSYpyPVznI0pwxgJAs
c8nLWZan3s0Cbhrh6knWlIDPMCyIFK6/k8RTA9Je+mq1I0NwwlHurjQ7Jd1QAff1P7WehNhgcDXk
2SAgdJ8vsUhWBgwQQ6B7Lg9FP1zDpoGBWNfJv9wM0i3YR2UMOtDKyIFlT+zdAPlBFdDILV5qAr1S
2x87a04qBc1EUf/5zrx0kj0tEQrYsn3hKJHCYDG3t2idEGoKf99KzhIPZ/x3vsaM7wnfGr18hMZu
OunvAgqfLWJfmIG3iaFJjtHzrTVEHDAyyDzZ3XSeTtltsKuRtYjmNi2GOOrOAxnuo5X/j7qDjtMo
ofpA7Seitv479NyUsAHBGawcytY4FJtshiKosOUHAGoOhk7J7jT6Bt0e1m5ZK4aVNvAHeKOj4NRo
IbZUSZYV6yvQ3tHOBWfs2/DAZ4W59ZkQWsD4+S/R735M8Y/G+apz1FHUUYS+o3V6OTIzCtWuoD+h
ScH95PKY97lY1wHSkJYe7YGiZQmN/OJFIKoO/GplABEu6N5DVAla4zsqh0aShdBLCphMAcGCQeqn
s8eeqbqiffYFBpBstrHW926QhqctEqiKW5QiAqm37yystIhxmQoWtlm5DvSVJBfkyvisFSlHx8mP
BsYiPBIDunzmt6AOqZuT71di3I8hHn5KCuLdffhbEn4V/Gwn2lLDLkxf4RKymF3zzyz6xOSjnYrG
Xu6bS5LmXJqMTMZhUPfd2g0srux1k0noFrDHDLlS6m56voFuMAQ3FNm9leFFP5pdZvRYxwVDglgE
6654slVURpmydTy7auKT8GsNDLJuiOyc9OKqnHP/8jZsoMfZOnv7Y6Y8DxljTM3v/qSqTIBSdfIK
uLCYNt+SkRsEfvr3lyzknj3uddEFMSRQxSmKG9ynkC/Oizs42ozdH9mXWj4j3KEuhCfVWDxBJ93Y
thitj5HKwG1klxF9vngvJV/UsYAjxI+RXXYskHOpH0Ml+AUaEw5QfzK/E7oVild6AeIbXPbq9jWD
cdaPDHUJHejCboxeTla03Jq9dSUq73Oxt254JtPJtQ/ikWWBFS86K3qSyuFLRiMtHvUP4wdZHZUS
lzCG4Yu1iqbMESYB9RHuAsfqEfpssuFa3XkQ46AvvOZdO/zGURMw/GVfKytS4ecxypR/tpgnjeKd
NvDKLGlCu+NvRjLjPg9Wndi90bKbB01VCsswIV18xtcCCYsmFS4A6WFdeMI0Mq1GAlB6Y6sbkkzp
x8IF6n9JMt0TaYL3axMRB2sc34qPKkJhRex9rAOdzdMTZxDIB6uPKMQmjLTvDA8Fx8bcUTmq5Rz2
rIaxphj+QY0P+MFnYOIV2ksTHgAgkqwxucXfkjlO1yle7P6XEl0/3hPeDqgjrW1NyKxOd5iHLQ/b
vmTio4MPKoWIk7uirVRE5FP8LrNuO2Dp2CU06P+ZSIHm3OvF0Uo/2CLve4yv2kSvFVQQhnWJunxf
a+h9GapjDLMMYiwMHM0VnsfjnwJxwQA9qbFdRjAj9fc+gEvAOBpl4575M93g8J8VCRc1THmJABey
yk4BvevV0pthjtot7GKSS30aoMXX7Q4GpCPrSqeQEov69seEDJxvWFOP4QAhd6oGsUZ2lQhNo9AT
10gLwp91ByL7/N8hgmuSq9TFAa+emmPKMRfMYjVUK8wstoiiHQeaRX4sJ7Q8XRQQ9QtEDHKlbUUs
73BA715pUyEB2UHMXbpU3SK9EWXjIPgceF+WrgC+dfZJMCxbpyE6yIXkqjVeK/Re6tZsdJqLPzTy
tf1/ykRXnYkfp5wBvA74l43r62DZHy0XeuH3SB5V3EkcNyvVt9gCOoSYH+CHq4tf1mWmeO2nEZ+T
H30QNgeVXmslcFB6etcQhqBAyZFLhaETmR4Pcbu7cBgYR7GlpiPlrvmgaSKamnvEQeq+rOy2C8Za
8hT26hYtbyvGzrui3K7VfYsqkJQg7t/RkTgQmz0gbPPs/qEFZtcd5DzEPWLZqZUapx3vlIypKHPk
NizzOY7PejPWf+ieFq+WsC/83rYkMCt5Cqa7leG1wVUSL6cHvIto7WQrT/qe8BBGgFJV771JJd8Q
iL+56Ua/tLuA6yd93QzuLnh8vEOY22VUETgs76i6e2QXCEUDWW1xD0VvicN9keDCmDJiC0eqv4kC
ViRGK1ysHnqRdxaXcLXFkPzrrIxKI+xEgv9AW5TtOGvxex3MKlKCCXsY1GWkEsnB32GPVxaAHvrT
71ixdWhhHFjy+BE/Nwpq2uwt5Ksc05CMDNvdq2ug+mh7YtrQPg/wUEC02VuC4OtfZ80hcdvONGEK
cVO3Ifx1fCV+QbsSKMRV7Rmb2NuyN7KdrvHxSw1+ZBlckBfFVoV0M+KCw6HqvRjqivxZa/Br1N5J
22Pc8ZeROGCeL8ONuTGaIQ15WkfomP8N3Ox4HYRUioANFWtHGFtQbYv99poVwe+g/HXvFYweqcr4
bNYFzSAcFWGwam6u8dWcw63wi0TTPF/KqUFtrKMxMWTF2QJCzkHpLcn5PvAUfoY53Tzil1DRK6aV
dm06qv3UcfO6K4pEz4eMggnXdfhd6Fd/kL76fOZHHZy9PufvCvC2GNuXtPEzwiofN7RtMydcrceS
1J1NU1rta9tOhyKzv001yxNWF3JC3ACCes2DQ+jCSPJajnWYBK5F5TEcuRoSzCWjA+TxNQwzh03a
bKEf0teVv1cq2ZZ5QWlvkbXVbhboeZkAEvnYN2Bvmr/8TLAUBSBhWBrlWgZyFiIIchATygpXC3oy
9WQPr38lkIzlx5y5g2ZfP5LLy/KdTTYLMHWRoJRnMuG7eN+0eXCqAOE4j+F2alM6zeb5D7gMHu7r
+8taEi0lui5Xe0xjacqvq8uYEuJeMHoaYYfBY8PMugV4fBKsZ1hjTHK2WMDiwLXXt5fzeH+qDNwA
4K/VvAxcBLztuT/9Is+n5VxtgL/2mYdIbZcjkAzKfGgCf8K7aAzszngSqWpNB4s4oXQGqlo3Ijyq
tKDpVP5q45MLuGxZkzHapO4Hme4y59mGzLLSE5+rxzi+mtnhyHXZaMfHXD25LSpGPEpLx8+b7JBt
6u96ZVj4YcmzmwdngZO7CwpY8WpG1djWpa9Z74ephtDtR1lznuoepNAnLXXQ3Q66GL/XIxCzQdLJ
ojR27o8k6GBhieeEJ29iNCOi6Eif1hEPGQAPmJdbyhxLvcEucpOs/og9wQZLyxqECWjDWNA2dhdR
5xEsQIFA2gOUyohzSWFkC4UaPds1VSodkL76cXjygHawIOTKJDfk6lo0yU1xS38fJmkU2IjL+T+s
4mBA7v6/gwjFTAmQjNpVRfiwT80tFIk3i7RsTm2sR5OU8DIJCL1TrjFo05fSDiD6eOUvGQ0vPR/u
6EaGVYvOe/8GDX5e28NxEkA1Achwko2TNDHUNlvH3q73pLp4f9mc3MjOJFdsXJvVPosoNXSWyTu+
8PRHqOJ8y+yqDYhyIv3GPso5oouxkVWoSwNohv6BuTAyEyavogW/vmhqzMaB58pzjpXxJZZSr+Pc
T2AKwOHPQztobxZu2F0L+iS0fol9OBPwd8S+8z5PvvU9HKPmNJbt+1vj2CyIYxuqaSc96myRGZPc
BWRT3UC5qdYTGhls4IManIDd3un1ovSiswFkEeEcMV8CL2n8jmVaXGgloYbUVth5MVOs2YlG/A4A
DovSew1PH4pdewRgP9HnnFXr8bNXstCmptMxG6xXWEAHoYtLuKthF5NPYZpwd/GDLY8/5YsRJmtC
eDII13BO7v+iojXoHIxVwZEL/AXF8aueDDXr2HGs0hHpWv0nYU1h1ttrRDi+z6KZpk+eSbrzqRml
I8x97sBzessrHhNH/nEkG53HKNoAY57IieofoXuE3mhWFKjxR6phuaKVwDjvuvqlZ3iwgGgwkxjT
0VrCQF+4Z7UGpZ56t/j1GvkV+ouwPq5BoficjB9rXEOJezMHvOdBQy0QpkVvZjVqkqvUQ3Chgenh
Rm8SbyLvQHUN7byzIFgsX+y5qPRm4n++hQeai9G5XWC67gmEUAwQ+DUXkqg2BfchqsQLBojLAyIQ
dlfQTivnyMzOoq29/6aMz9zg4HbsON1cLuwEnuEARHFJ650pQgn6wkytVsrlY2TYOMwgqvHr5i4e
6pMrgcqMEUk9YcW2sB87YBtLZgf5Ts/IQ6R9WwJldeiLVKFNxID1Fs5Ny6FzxJznRug2ipdxsvQF
qMcZ8FcZMMfNb9WmXn9y/W0t9xgIe2pfC18TBRJ6UkRSVDJhw6PEr6heJYN+oontIR6zfb2dIL9D
eLI1rHv2IZmdLqmzA6zncknFHyjACJDAcR6j1EAaaOxAd6HOJZoA5+T340a0Wfz9BdXIFznqm8TN
8wzld0wlmsX7qRLZqR9Pa8oIOr2alUVU5h0l5S6wlAyRYzhRUbjP+Ch3SD1kkG/bQZCu6JuYVetn
Ehmvje/HgiMjO6JfOfG5EcROcWM6d53gL2jvA3lExegbjhHj+uLeCeo6j9v0nokKkC1SgrNOGRbp
F3aFpP/iqMpldiAOX7OugnzOKihB+P7GeW/b4wEsOKdeI0RpW+Pm9TvELTSXkbneQC2DL0z3CSjn
CfZQCA1Wgrx6O8lQgrwxKiC5IodtHSKteKcAQ7P1mYA6WS3nShZoUEY9x1Xm+Rd/m6RUKhiJFwEb
FftSzNsXCE6f1qU+yROCVKZNPqlH1qL55Qmi/woJE7XPVKMB3OshOsS6vanN3jpXO13J7GmRqejR
VVDc/S2lyRrjvcj3BOlcGhMeDettcBRVRTB5XiT0umKT7EBe0fYu2JrB5Qv14mRFtmA1tTTvGbfS
0BxwZlWlxi9umntP920pgeszvlRY83bGn+wWswraGmN3UsFD62FLnpq0jrlEEIAsMeKvb0N3bz3c
ofI1LulEd8aT0PrWKY4Tb+PNLLld8KKhJxHOhnB+ZNwc1WAjBFI0eQqWEdbuV14EAeFOHqAK0bek
cI63SwX2rFWs+rtAeymZnCEeAEnE98lZMu/hbESdh1E9wsGiuJ2gSMj8Lo3xmdHx/s8lMDRDZ+Z0
Md4FZB/4jXFwFbajHC0Es+omGeUOwBp2tZ37n5bPpc884n2SwIw83V0P9K3mJLPG6VcgTwUWt+Yi
zw9j3vroJ/orkO643nvqVIhYAvQNC9+uLJZB3aGNZArGv5Iv9QGlHxZLUPHYI+1bwGeQUdLfpsud
ZwlkxmVwG6d7yrgZh/RDgm+G83EVHqxiK8SeNkAKxGyEJRkmiXqVQmFV91SHskeofjF2ACUQvEsr
2xwtPz/T8baeOnlPomJQk2FVEMTINEyejXGc2Mqzq7ZsP97xQ0BoUzl0dCcVbsl2yzFqp4GeO/Qb
e+ntw7Eklef6rKu+onWRYhHVQImXcvyTv1LViLfUbyAx08MPNd+kf0z6W7bN+tzONCtiPjyvjImz
TrIA4ASIDHJFQpjkCI+hYYC0CCOnjrajjTfYl89go5MrvaDK/LsReHGsNyERYhZYaTlQY2gKsfr8
03Vjk2XYdwd3YuoCFIcZLgquUtT7dbqsKXtF4bVEdXmw26un2P1IVoZH/ImG66IGTnxs/rbv8fYV
HRw7WC1WU448oe23yNoi8SlAc3yWrTVueW/Gd3+0S8Rc0Fiz81hl2PDRNXxlroJvZHPQ4O39KyC4
cc8w7wjhuLCZXESkLMBWW/DrSl2THsiTcM4dcfQvgOiwiYGq/M6f94Sr1gW2gzn3q88WJk6lmsNH
vf5C2v/BZ7L0/KbdQBzXlC5LzKeFYyOusMH+S8SDvGpDruf0WPezK1DEyR9JBh2N0CuWQDxcQFTp
ikfRfM5aliJc/d7FlqxvN/XVyRvMgA10SVKtyXdk0Et7EDCvCPxyUUzerd+L3GI1gTt+rWFmrBi2
g5kfoUvrqsGwHruoY8edqru21cVYrWKe2FNV9CPG2VHFHwk7bNHm/A2vCqS9ZdDabgyXcccT/J74
VYNoWGTR+b2cmf1tPB1+QoHbS2vdsm9HFcnaLBg2dqKlpvwcyweHiGR5t35qzCkm137WhgC0B6SW
VxxmXEeDJ2EUhLNcWYOqx9I6oi/xypc4rDmW1HYxP/4zSkE2XYuWdkH6K2e1l2p6ug223aHjsykM
rsUrlltw9ROsSvzzvtGf6GFOjJWy5OFp3d8P8373gVwcJsERNlRT3Lq0xdDUGQEA4TRZmF1dJl4p
LnZYF8wQlHjgd/T8NE8fKpd4YPAvsDMc7cOku7rt/ol8sp51LW2Lo0JnAJ5kUO99y9cZEQLBL3XT
wPvU9UsjxcybGtH9xfEKj0jUcDOLATEY8PmY04JjQiEeGEfYVNJJGs7y1JF+vLb7V7LE8NMapWmX
JKjJ952x098/2kktLK1lK7hS4h497fxx4sb40ME+nZjXhIS03h9J0Xi5IwZqXWK7Ij8B2MKsfW1S
CtlrLCS+QAD4lE2FA3pRCd4+FkVh6lKhlznIs5/s3yvnPrqaVjVMYRLwDL4gG9C3xY0nzGLdjBz3
KrX6EfkjIEWy/8i5/X1UAgl8MMd/FBa0NQvGQVeNLTycdUVKOJURSOqxu6KI3o+VkCgkQfSfZMEZ
KflNvjBwJplRLe3NcbMlqURHg53r0YLP3McNJcpp7Q0Z342oo7VDRfpA4wgHfxzDUj5zGxowJn08
GHQEn1jur/ZER8uscbj4CXiskucbiDDvJlHsvxQccBqMLiy2NMz/qf/yrOmbRn8kXESGcoU0eWG3
ddR6XotT6Y8mUoKUlfLnTHGB+NrvCar/Z5Muzixbvmiy3qLvh9KXgwocIw69mHRWhkO1tYOPTfcT
IK7hjKDq/b5V/G/X+cIZTcPqY++Woesoae34EW5FwD9dL2Qk8o3yvzoM1cWU9OYball5C5zbl8Dr
i96HS9LH+9jo3qaIpypqbrraw9r5ZAM1b72u69twRBexUmy/ez/pwgG7nLYsJRaIP1xc9o0zHA/5
pt0y8GzrTHvVrGUYyjjlR1WpERb9avDu2Ljxd2zjCDGAQk+6q0TR1OXc8eKfW/vr2CnVeOdJq9s5
78oiQcaJAwrQUjMmdoOyxAFb0V8T21/pKRRfi/ktaLNMm7aoq7Ky3ItlIZddXb71i67hrndi+SgK
/cmEvTTFce+eNfd+97ysoZEG7k76lTZfXAWufbod3u8rkCJp+Uls8psTlxtma5mERfdUSVOw+ALe
3BN186FB6ux57qBgumK0WiVKR3tz3jkMMBLzEVRWk7xfIQMTTZcYX6i1nf8Gr873iIrSudCFIcPu
w1+/WTcr6W0HNzfK1fVdE5IiQS6Z2Z8XxUz0BKAFuhPri4fDVJoxnICXGn2rirRSSPTaG7c46k3v
TE/aoKqsnt/Oqi75KGBjE6IGrwXBdPp6lCrXYeQbH68LiReN6OwHoB5ose63I8M4u3CDlhHJjqQA
YOJbbTPulIiyDSefeV05y0J59itJAHta6+/+ka5PVRTTPENl5Ahb2sUZZxJ3E8qEqhkHk7bNuXnS
kBdwqHpStTeBWi/S7LjdW1kOddI+yotpwiOeV6G4+/lXG5FbNvEOHf2Cre3CGEZ3PFyxXAqLa7V/
P5Z8pUHC2ffki13/T5vpIYMjukfn+UOuEtl6enjzxN9y8W2ov42pF6H/L4hs3qlqI7gJFRhkj+3L
MA/4XtCaFE0N8mXvWxbz3qhAAezYEgqNOkNzF3NCaWHm9XT/A+CG77bfutU2ah2C7uIn4meub+OW
NJqCQXPrM9tnq/W3KhJE2DwHB7pHeL+PDLj+d7Qpt0/BUU4dMgrrC7znoeC2KUxZGocxjgQ5dQud
9XfYxFpK/8iehCfdrCZ3pTGJDlGYu2/0d2a6IcApz7AetT/ZULbLVf5rE6P/i34/GpA5WX7XIw2K
7J7E4vp9cdylCoQvTrrnT/gNGmU12Y4M8eKH7aZWw5gsiMmB06AwpDdnxOKBPvcBlpiHWUMfq7hc
zBOa1hU/ovuwJ/0hhjDQ8xIhh/XSriV6bMzQpVA+T/igfwHB6Rl9Utifm3F02uTxy7VBv60Iya8P
C6E01kg8SquaADQo75mti3E8pr5sDh8d6W55jmM7PGPun1YpNARxr1JPb8rGFd36v33B5cDn3+kG
uduwYA9sMcZO9gfMuPQYP8doHBsLAef/lgxqMfTJFEcVhw0V4VU36Rr4jIkh9QoImSiAVg7pL3qv
l72D1nKHb3wSeNkhNWTwwVvcmK4H41FsaP/xxYxt8CswloFWa1HtYyoqwpIKnf8t8SwEJbN2cJIr
saLkBQWe2o1Ii/V1+NFndso8B255g1bmVVTT/bWoomw/jnkyjmPbDbYZUweW661AcXH3ROQLJgfJ
JVyIN75yRVty5keILAPfbmYtwJdTdQNHwW3XPcqXSWQWXXeb3eJxU+4eJm8hiOIN+gtxHqrifs8d
Y/I4pvtTJPdsel1iRDBBAidaz62FjNCyRTSOhx/4y4nz164J/CkFP2Fa64nfVl1tFwYLTL0h2SQx
NTOzCITmydxKGLaIsUlaRG8oWbjHB29TJdnVZTPcnn6QxxxVhL/uTJs6uDgwnE0xjInqSWkPD0SE
dP2tC2ojbVDNnaeVj0vnuc7zFEnx+a1ejwMiubadeWlfdy8A2XlxVWHC7mbgh49DmmSsQuirIj+3
dEyBp8kKIWwCzp9WP9tTDJNBkasNj+HikGNtI3XYLE097ORS6z5nfKQm2PvXA5DwDJTyBgluVkiK
wXadCVHsv0vVlR6F4Hz+zZ21mZva4yAsSAWQL97xY9/8igxtTI+eYEPEsEp4p658VqYvaS9FwKuJ
0EtB1leCczfa4IwqPJ7dO5X/O49/eKuTISMJG22Wmvoon9QuphBfCzquhff6ixnaCswt2Gg2t9S/
nZfw/qdtTtnmEXXCWAZmyV31YHM1cOqut59L4lhWqh5YJ7iDl6N6Eeiq9yPiEBFhneCeTOzGkKSA
YJ5eu2oSprJMZY1fEjzoWUV4d7x5mXXJmXJ09Zcb/ZHcFtPMu5pBrhdAKBtIzvA1aoauREPy3AKV
qL8DhTpvpbz2cU3ERx2k50ChH2znQjutQ4Oe69rxdaaYadHPv+ioDyt+JuX63eRbx8XJdMO7v441
ZV/nCkVNk4UIryTZoGjbR3k6IhuNiiQ/ttgmW3jBIhIRgic+XtgnX1+exAtbdni2msTCM5byLEMi
dRb6ON1GUYwJy3pgAypcdg9DAu0DMxFQtT16OkDQOyx4TKd0OsGxYoKdQxX39KSzM+M25LeHedzw
/dh2WJK7zFRnr+tgjDgOfnKHr4I0P/7LWM11HM9iM0L+Kvn8GV4TP8QGMFLjnETGxR8Cylie+b0Y
Nl0ywRUXyy5pNV9grU/wl+zrQizdRckVfXmjdqnVEAy1vp1pQEP4s531oqILU4GzKO6QAiG2QvT2
iddunwq+culRSXiQfSRX53n9hvLi80m87Bs7UA/QNkEX8Ozfij9Ozm/ihDykmsTTdbY52yHZf1zs
X6ChgA/zRKdMo3+2/gc671M+Jissnaq5QLs1gS/FoFTuTy9UCPGkngJsCH8ua+DQA/adWH0/skZt
OqxSUYa4kkB4JQ8C16LShibjpKsyA/Zw0AbakniAMpTJ3nv7AJL7xe7YT/rmPIqTTCR/B0M+pl6n
QSib3fxfiIl/w4rWkbFqOicWVkp+VqB1g0aLG9tNhHCtvnCN+7KaGdrhTsH6WA+XKH+PzSFLt5Mn
/MlWgLjrAnKYAQj/Q9Ti9OH6def2tEcGw6WUU+AdIKs6vLWEVN1Z1XLtQnOvB0FC/nbPFsbQxZII
Qfl9rT+vGxrTaMnvpJapP+iekPQz0Y6IqCU2gSuj0rWMPWO57WitHDmqzs/yVuWLQtvEf3JgOLfa
pZIMJfxourNgzx2VOPMIoXMAodOr/Tmibd/1W+5SRCq3TbZNoIAl/tUMIl03VPcU5P0Np2UuE1z+
Dxq/+HBu8cBARRozCWHPRZyfiADkvlwLLIgACvVeW30VslP8tiTWAMsSEDwhocNzahj1Y5ExELEk
4K+uvhv8RkhQCK1utSHnVIcw4/6yyuEIYnjGz6yXp0RLH75Hvykkd/+RRMh4ctv1TaLlCyYABqir
CALQmgjq079GVtYAoJRlsPL7EX5xBJbzFWcTqD/fHWb4r0PZrovqN4eNNW1c0graxCyJ0Bw9DjX8
GVX0wzwTwEiEJQp8w3KQ4AOo7LgGTXhnSYMy/jLyG5hIIwzZwyOwpvtc/5Kum8TWDsUthAGV7KHS
EcppshRkRYfG4EYT/riOdw85+NcxMfEsKjQo/GcXLjH6Gc3a7mYA7GW7MkSzgNvDf1iN7xttpiyr
w2Jyab4LIE8VjXib3ATUSMQ9gk8sgO5ZEw5sR4WnqSGMHJ6bvxmVxwy/qslZb02D0FQdpve7jnU1
9bywfrHV9kUvlDB8VtXTNvzIn43UAqt3dQ8shH/cAUCXaPOqo7BfEOFLePWknrpNBx0AZUPtjs4/
6Qx1NlE6AVEMVtv7zz2RpO2Np9jlefZjc26PbH3OlC6GL6c4KcVRQpxoX7+Nyb3FCcsGdxzwvvgx
Jm3Jt6ICZAL2RKpRezYuhT0XZDFezuUUO8cdJ7JhjYZ0DEW+fYYXnMLz8xi+/AeyTGzlhmldXC95
XbWo92Zi81bKiTooEKQT2TLNVHfEQ4D5jrVTUXUtg8pNxnDqVLVsMPT9VkuCvvj75LT/sxz+Ktjc
1bVDEQnC9getMbzCSedGuzvKsjDKEwHhxfv+41bXyF5ywaU8osE7S3Uhm0TqpsPF8I5KX+8ViC13
0HCpd6QVoz3BRxbpkG5rtRjjlM6DaikAib/8pj7eGUeoqYA2WBtun+0hxnvx+TQLPJKjJBO7rGq2
820J+QQfuYp8sDmyLRyeb86Lxn8PSY/opjzTFfwq/qPgaUwSTCe+XDnBrF53+YB5Ex2vePNvRQ8T
mcnkCoNqeeOhQlqZmwMoaza7UZLvXJOn0cmhFv/zvC+H61wmcNraUCQ+ghA9Vwyfnpnv2wq5S1NI
zUgWluQ+rYWdSHKuqWykjEEg/kZZ7eRXf0901iz590u95DBC1AYKKlX/au48qcjhydDLhqTWRY86
biH1pEP8pRL57gV7EhCemn0kQP9rVDESoUsTvgNIuI8YGW/QrWXwqFXR+O4TtuKpiKQLZA/Idx1I
3uJ9WMAqCkUorYefG5/wpx7iYmdzg708nDUFebZTU8TqDVB51loprTu7N9MKzLhxdnmpKXoQALul
RbPaOR4hN2DKZY9dmBidQkZjsdVCkxQd4uX159dE+7aBapu2C78MWDWIjhJBUGG4bIUUiSAI8M+e
zWMaUmlp4feG2MwBx7R70jKfYZVCwlEP659NwaArZuNjMHXYo3ZY24mYWs5I3acIpsjLzLb3m19h
YTHapAmRUSJy5qcwqR+RE5W0HyBotKADv0yTq2lQjXvBJ2BmNKUhJnJ/o6tYFJYIqI4V6onhpco+
/sDsg6HDL4AWtYva2JLawK2OckuZHxtFCvm6mb2LmRUl9zRv1Aid/FjfnsWVS4gvwbPA9NNBr3qe
OZlmfgOtZ3p+A3OcTRW3UDt3wGNlNKlmysyG4yi55GsTNE3KU6BtZeM6Lqm0/UKzObka81Z1Qsp1
0g4U5V5PlpIR/qqrlGgx36wlH7kK8a9ehEDfKLP7tf5iyR1Ti1x4+wIAoWUG+S/36yPYF+Ck/juO
sRdN4HavGxh3ygUEzy/L4jzb0qxVEoyWHyBmofU3rkWzRG/o+r8BdWiGtEU2jxdWh/gsur5neY2d
ukqOvZTQwJjhPU0YVynUtkYOKw8g8oj40+zdLWlYl2Xo2eKBtBeSS4XfQTLqcfcHjnuemmByn+wo
amCpwIuERq1knJb5STkA30vwjY6byn/8VLTYg089+9NJhirUZj4xVy6EtS6vMx9YJIZ6ZdKuQu5g
u7y4zTtCpadLJHA6cb32imegfE7Z0p8ciw1aDufAk8xOnN6IHoRI9I1xKwnPDlPlodOqLWapxlnc
5VNepAplmatmK3tcqdKomDMnkAKqp0z/o70/8QP6H8FINYvK17EjTqoUxaSz+C8AnPt1jiuIHjH6
0jBocZZJQjSzfy76v/cSnIi3cQR0MaVbfQzGM4GeJdGpFFuHrNpH+7nCHD8DuhcApuFCEZMsNJs1
c2aa4kPb8GS/Vru+cMZkbKhsA7zuWXzpPpTnUzISjrwBppgV2y5/TljMPiIhmuxPh9dL2qAZYer5
8MIK1lK5SAubwFlBv1MGnPTUnQmFc9QPZ7zMnq3qJ9dCOliqrR/nKqp/JAv/L3yoG5mHcV5lywZc
TC/OGor9uZgPLC0QP80TFD8TzY7MjY9h3yPMVy4DmhMTedi2FPJBLaCi+3OstgVbGZPHsK5mWlSb
QAo+etBAvUjNgLWs+ogDMmmXBvkODCl12DYew+QiCCrwzYDw4M+RnFLBgxXX52qXsZ3/3cI/+AqL
/xz3lwGJtLrg1w/o4QhgG2+Vj5zSD1mR+9e6Qak57ThqZJGQsgzx2ByZkgs4gOXskDTykw4JsDKp
wCIpGNDMd3pS5nzPCNVv4VyMKrfCzGS+xrTPei3Un4uPAY+zOmDEEp1Z+bli5RrgRtfUsDsWRs3E
3RZg4XUEzcsSfex5Rq1hht9Mt4wbS0WxwG/uj6hlrCrqSQumVj3bNDrINSqHak1z7r1lHA9UOqR8
fWCZqMMqw/AGRR2dFDSdOJiu13GlA3is4PTjggCB/PUY8bjFUG+hSqru3urhTery5Yz2JoS6YF9E
mFRv+bhe1ZJGLLCiLpe0hM7oV1r3RFQ7WUpnYOA/do6aFJW0A5adco7Qr7Qoih48DQI7MYMs8KP4
gXOEoJRxlZwRaQP+u5T4DSC5bOw30KNoK6HKuTPPioePUmd+iWTGDBQhLdbpkVTU8WcbX6+Xg3/c
BiNJ3EXusT0F15LhgQbsE2s9Q9T4qPunMQEL7+Tz44dvjH01Rb2rL6gQSY5C5n+Sud12ucTtxmqv
kt78u0KQgMejUuonSUr1+9xyBwhNBYNWbRdMItCCIqA7C1nlMdp0THfTWlnRey5KhWD8Uk3EXWUF
kLiSyjXkOLrqXTTB+Fup9PJuSDyhbgzlom7uoizIpXSdTRTQTo8/ATb+guiehkDh7z1OJcHVnveL
1+Cs3qIWqJK/XWpfpT55n98U1qSekeMjN/fGNpYd1tZBewPT1U5SKDzn5H85FjaX+Lvcoh+HKLt3
HLuEwF6Fx84D6XFLD2RIfnoLv9yoRqg6top7yCFWCEtTjG8Sdf8yNGKfEsu3oqJmRet09dcJFvcv
GJhYAkBQsN37TxB/0HgzZHPa8ZF/uRcVJzq9eOKez94/mXAlUGk6Rcka1IaXyUJ8N9CJftGPoqkh
xeuzVS7LAJYKScOkzYjT7Y5fBqkuSDBHOovZAcBhQauSHgg5QwvRnIhK5RKkm0KU+h8MTKfTqUeo
qHLfkaGu5z8UgfH9RY+A3ZB5XhfDZsYblxPSZ8rd8vpaJ4Z92llBXdiYJQWgO8ManoPtVmm47D5C
7199rX33RpL9WscIcBkMclqvYk29zORJ+7+wUgey8yVO+HwLPI+Pyigt/MTQo+T2rhMDgfXt/RP7
7fir5A7dILQYlzOVNLIzkFJR04bx//jvWW/3LajNtl6FJcIajgTGX3TipwwsE+mNlQoQETXjr6zP
9kSW4f0zw4FYmjxoCEtzQ41QI1Vw0Tmwby9zNnMNGnw8PPKtKLHlTokW/KgMm5URYgLTaOrPUQFT
mboBjRwY2b70WegGjDnuyeCJx4vQxxDB7yWrDtu/GFc7zVayZg3D6soQDIssTcw7hXq7WmqKNCpD
Fl8ejpNDcPH5bFOlkI1Jt/c/amGww9ZxXCZf+B+fp5CdsfLhFHGFPRkaq54X4Bgz+oIiTyMD9pYt
9xHUPEYj9xKKSd/JY7D79bHHXC4b6fMoqpUxpuH/F4gBjnSiM4XKTDCCkOW1sNxBeEULcsX48apu
gC5meurDVuIPH9uyQRm3BVzayAbIW2ZJrW2xuLIeoZssCox9vhbCaWvdS+d2MJKjdbFFo7tJbM7e
kbbs5JCrLoAvCQkRtLd5jNH5rek7Ph1PYuUAIp/FoRzmJl328H1nfOvC7uYM0WLFLnYUmhbtTs2d
lpQcwrx+U4OAGLbex5I9M2Tondprv7+VJoIOkLXxwJJz2CXp7pzi32udauhUOFjCxD3L4Yy3JygI
btvgTQYlxtVdBNXYnw2OiA1vvvIgX9IgXvh3u7yvv6v4wcWe/Xfda+e3t5x4upYxZjDu0+uK+leN
D9Y3DX+B9hFR6d8DEADaX2Rd+RED7SWGZCGnu8JaHX3c6LrP0WF5DoTHsy6Cyj8/RGkPAR8S2lLm
Y5zFSUaquJK38/GCryJThIKKVb6ynhK75U/P+zdmJSzRzGof9XhbtryMjlv6flNl0H8L9Yw2wFl3
FHp024+6YBnB9llPrvV+VCOAi7HRFZg395wEaWP1JYCk2mOIhmpH1dI8j00FP5TlOelGcxmliHq2
mBe9ysliouqPgfUrxk33R9NgkQvfjT1NGfullduiNt2613Dchj8itpAc0D1RQGPCqzCiFG1HtRmk
3GAxjWAgDf/lSWF2ai/lKRpC10DhP8XD2cn/x9aUB1UTiz0RjVgqu2y/1rTkQP+8EBPkPgreBaQQ
weM5kBb52vgIfAfxJIhzyOvonfn/NovCHyzWrYf/GDZ9xMhbBhtOYsNay9iTGrM6ouHruKoZ3jFb
LcekAUMiQQqZ/kjD6UELpqaFVFt08XS3NyfF7WYt73heuu5Ath29bEXRVzZapOhU4mhA2WkwazaG
8IVIaJyaKXGFwtEiO9o+EWN6EG34ZoVpvDNrACkF+5ZdlbhZEDtmq0uNoGvv6mjC3e7E5zQm3kuH
Vkrlq20DCxb2a0jBXi6xbGkShU3zOa3XMJW6Lj6STORQRZdPcL3qMHp+PG9hpE050cSsC6z2NMNP
qo8yjJiM4Tbmg6Xo/3r12bKyf9PVVQm0wsuIGbCeK717WxZWTNlgBi3pPWyaFxlmyQXpVdXxwkgh
F58djcCJ+UtfFDpB7bbOKFT+yO84scuA9jfy6zHSjiEHANV3CsRaW8QkUoqIfFP5hEUkl15BJZe/
srINw5dxm/X9fotkXrQEfdm8NJdsciQKA5nLxQYLXS6+JeRpNxzc8h+9BW0lMjEy67PEwJtXFk+i
ckN7hgs30/rW8I7XIu5/ywnbR3R+dUj6sDrdrp81vB/WphxsBoHPpdqbDSvHnDZ9G71+I0SDKx6j
zmvZpxBMoR7+wtii58CgfH+mwbG2SM3c2E/4Z61Ph1t9qwOjVlXfBcQ1Oy8dc68AiScnTC/O2pjl
fnpdO9i3IPc6oSPzxz4SPwi5ti8KSMEajD9rq4Svli5HpJErx51zuAxXd6OAsaqCevDSplW+Hg3R
rCmnuMiRYyPC+xx+Pz/whTj4rNlKUvYhYTwY1fuglnCzlnpXrseLX/WHJ/xcz+9GkFxARoPZtSfZ
/ufh4lhJQ3PsQmsw3DNrb2JrXZ4DJ8LR2w/nCnMG11Yo8cWVAUw4xGhnMnKmieqFoo0mu7AIusoi
Or6S3Pcam26QYsT12BCjn5WpF+mF/CsqVuGek06c3vZed+hYYhTxG6bHoMBWO0MFIhr3UDe2Ovja
JUNnthDaoiS34qIw4L3zYzzyz4HQkrZkSIvqgbuj/LFRU1RY1Rj8W8v8mgED8txppVsd0JjDKGoC
kiidQRitqKgxLvgm0BTgkFsIDP52owiyW/Bk/SlTxyjH2ShDLP2Ms4+HqBmjHZzuTmI6qwwjeGLW
mFR3/j735915JuM8JezjIKubfe5ugAnMLQ0MWLeePuUQaY+WTro/R49Xm5iCzmkcf/wj9WVgEds2
fqSH3GO1SCJRVm2xsDAGb4hjB0z58gvB9ztnKDwEgm9nFfOXrZ1MH8Z0MY4q4vngrocQNv0yNDib
g14NTre+vLKZm5XQloicLLW5hYeDIp/MBUG2zF3B4r30ulRo9VwjDTqW1fcbfQEho59VdXUyALdf
+c4/eto62VKOlNHGisDIiwKjenR+yfSi1zpclXjUQ3LUXw0QkbYLBjcF3bR8Vdl9YMb4lIjiiHig
wrarn6wS7Pivl0TrXYLWh6/lfzkdtS2uyVOmiC+ln8KY4zqV+iq6Cg5KbVGH4A6RUdlkl6ldTH2D
nQCr+DAk5JBwwL9NfVZmIUFxQ2nshrjjKFVbtBkfBIYd3Z6KT0bm0T+TUAawtfx1o+0uvjD0qyG0
0bRdJaMMAmTgbgVhj2ZzUGs75Nzt42qSRRqXpr3Z5ibPqflFGbvkCcC0q70lHoUKmMoo78qMBFGH
OdmA3hZeavS3fzy79YwN3MQ5iJQhKcmW3/aV1dorxanVMHmGjW1sVvwCqa6GDZ+8/RzZZjQztQw6
IQQ4/hx06o0FpJJzn6v92jlygqB33p9ryKMNGZw6zCqj3q7fX1IaVd7h6Dr3Gn5EXs7nkK7UeiKL
U8KxvwVtHtA41epw3ZgmU8xvgC4qPbKqFPPUhlkbM+Hf3343SQjxoENWW/wzQXMsyTpcWy9eCeki
zktDzizvdno5lrw64W2Q2+Sh7oLW0dMNsw+8XLJr4yfKsY6KuVUkzwXx4OopW6/aL3lxPFkJw31g
IU/78fodUbA2RwsPDm1GzfwlsZEPsF5QZY0tEn/BQfB7awc0O4DEFqILex8R17y9ltWcfEUcPYtt
5sJbKD3OL8uMOz9+pVWq28beUZQBrPFYu0MbDN/pHRWIKBBNYk9kc7pJlY92dbKBC5wX/5J57/VG
i0SId6LaV/8O8BAy5OjSS4akG8WeOwGffizz4klS3pDGjazAqG1oV4k01H0l3+fw8grvK8YVzN5U
C1vuNP4Dm1r0fVyajL0w8Y295AWlSPbHDxWKGrryj3Gws3MOi5M0K0A9pWMP46YwKWr74bTouBxU
gUOj0v9OpyYZ3KRIcTEQo2FQtmjJl/0P0J/Da+Ug5V2nwS4WVCc6iQ813k55WgZxu/IrX8OToQGr
H0aGc8fkD8UeZNiz6N05o10hPjnqtrDQNhVHE+Z3bkYA7pfeFvGB3GMws6ZGSZk7VR37lPYeX5NL
E/WR38kWUh3tuOSmiZA+OVLQ/58iRVkic2BhjTKRsrqg8EyeJUuP5JaM+1R1HveDQgjch7/Dzpup
i1imy5JkaNCKV28Y33WY+ua/U62W1X2Rlfj6AhLEXAYdnMUPO+sJMG8VlMShCXOMg5NdYyHxc7C5
HKqz2t6fsPw4DmsMsKgqibxHYmHCtRzdUfFbiOzVghB9YJkAEotfHjBBeSWeEgFcyS7NH7GZfe6F
IGevkfeJoClyZ4NwAqaUUZLFhRY2tFSqSXjcAYQfzWsIA2uSNlg62mVVo0vJG+UFWa9wRrgL4XcG
bYbF4U6EG144yFvWyvn3Bt9AdR7EAd5mQy6fezHUJZl47NvMaL6kdf6e+ec7DGy91bW5JpLqPKVu
0WsoZ9813iD9iuYj5J+7bIWJCxasBKK7xiI4NHVrPSSLMXZjJ+8OyDSAsi6vgBsgGC4J+nOKtPrT
ZLXN8OBsgbyOU2tG4jgL69w4fKugeu++C73gr8/4N9zUSxQsOxonKUqNxyGavAolqn/Exih8OBEp
6Xh7wPodl+rmD2e4FUTmYdVjSw29hfJKC4hnS6uIynwOcWradWZmV8Dh50ExLMJFh15gY1f6M6iK
dRpgUl9gVvoWxIl4HBAEX4ix3FHcrVpDQhOndyKEUzF1Fopy7PAr1azpRLyJRfmbdNKC0reH4/qt
Xt7W63ZWOHpXtwZIVNpeUeQGhgHcoiqZPXjHBXZ7A3GRzqw6UNLkbnKObLXAhS5gruOTBH83dMzy
C5VwiFw5zmNUXsEF7Qry6+Cj1iU/LcEngUB1IW8VuMmB0BPKefAOGwQxXuDctcOonte8vZBsAVeu
beyAIxdB+4cpF0/w0TLtYIwpAbH2lzITC8kAssba1qHVI4tlTrW57AyOAnUMGHCEIx0c6meGZvvm
bw7b+s8E668YVyZpOiymCxtKhGQY2/VF9I5uE2TjBDpIuedaQVGGsrFnpUxSE8Ow9omI2pA9ALW2
s+S34/GLGABeYsFbhPmVJnZmlyrGCcO6hgYWzP75JaXCtqtKnfgcMA7ujCsDNcvWsJ9J9d370nbH
SwxoVBE1t2GgWzGRQCMQgmggwQWlA4yHinMIjnyjAF/JowZ8f9lVcz3RdYFc2kKIT6RO2fPP6lFB
q6IQbH8n+Idtya9AsYmwhAv27axAhS9xukNzv6V8PNMi6+KjlRcR9DylI1fvP3BZ/HLFpXvd6VmV
X56cxmROD4hj/YGFNWIOjXKY8ABesTXCFVoRvangKs9C8T7oinRqO+sNZNCoU+LC7j58RZkK/ID4
fHOHsqxW0SWYH9WS9LGqDDL/J/SNgufDOnMoc/eaZSfjh6shCllmhe/hSsjcdxh+N/buiql3f8zD
bA8Ah/xYd2zK2wPz5cTcxItsENzN4Lj0zbBwFkaE0hlwYhHrQMnPp0wjSXnM3p8aXKilIGWqhsnD
nY55BZkfXJFTHF5ZXfqB4sjsUr6AZcVE3ppdPeBLvZqRaSKCcsBfnyFX3qsYzTFrs/gtkTpGzNnB
WUSAyVmnWtwh1Em6BGHv037rCw3Y1lxKIVCpNiWWQ4xr3Pe23NweiItGdbpRaT78sWz1tjpfhZy/
U8w3+0Mm6fj3T6a2qjwlHulRcXs3TJzVLhRc2XMGwaOLjDwmLpvHjT39611y4Y7QhG6x+9j5HZNj
Q4/gjkcmE67Tlx5O/hpC0IU83SnC662WHJbOcGMFPI7qi38MQvoZNuBFTw7d4f6HnOuXB3L28K5L
a1WdQdEuswAF9Ii98KcTT3wjE6asEuPFMWhpTLJxFH5vdlFEhMruNNkCmP87gPAG1clGMyjyw9U2
R6GOyUfMH7B1qTeohNFxXLQo1k5GyFq8Jym6ype3d+Hp07+28XCN9iyRsyrhwHvUo8SPqZgeOwov
srPP38RplU+alpbFsGgHh7YRpOmM1ghpNdxRbCBcYhL3bDIe0U6FM0tKpCHY7h0j6GMXuUFL5uzl
qG9raq2+aivBdwg656JD6RoD/nSQa34mhHvqBTqfdrQyhRnt06RiDkSOsRVnyloCcG76ysNxpyny
5vq0z/W+Qwy42H6E3Qx8N9+q44uHyYJz31Kpcf6IXIvfpdkO8S97IpRZGdZNHn+CECnbwxD3gj42
PhyBBsYaVkiL9C2Epjo5EI0U8a1mGKQkz8l49oBC9BkJzL1tUfa1LZp8PvLNLBVlhiIm/c4moo9x
/r9p9Rs1w3JUOK1dgz0/jEW7BeDaCD2gagBthorQ7SP01d8s1i0x0FAvfCjqwMHfYxLL3vty26Xq
Axg+lpAOhfzfPXEV17HnYU8wVP70aun1N5OyZbFuR46c1+dECMjHUN8QmD8btVvpxuC2uAc18i7p
kOvBgJaSzq1EhJt0rOuS9msr1avwGshvHNEtZinDPMdOoBV275OXrXi/CA8bzPD1S9E40fBUJcFt
tfYGKFXZmx+rrJ2XSFg7uFRgx0RcjJNuLHsj8zBZAAHzdKPR07rXw/v66Fdkm8TyLUqnrjXL3zzO
9d8/cecskhJ1AylWG5vxa5uDp4AVsY7MdPkWlpMdIcVv8mC4O15teyJ3v0RZoFJMATdfVW9HbJlK
GycL1Qe7QorMot3JrB5edQGrlC1o0njZxGEZIWfUnFtTnV8xhNjBDlX2k1wFKu30npYc0/fimIND
X6Fft5bGdLPX36fMVmuvug0pPL4AQgTzn/5yLuqPpbFfIf2tqgkWbCNdh7L93t4tE741lvQCRarG
UqU+DqYyGlBlfIbFAaiyfgs2SXumOhw1p/Tgz0ZTcmRVwT1g7VmwUL6LfRwtfkPdAbuX/R0s5xNf
AgvQyioOtbd4HGDUY++eK6Mm0ion3pAIGfhH1yOlEWbhRZFRtc39Sf+xQQrLolv0+9KB10mFP2dV
VZlkRZuWWn5JBFBYyGF3JimNCkfwfjTGJCGR3aN82hsLT+iYREKXeYXN68MvkLf9BjZ3bjgN1vXd
6uPsQVuEWImR4h0oHDEWkqucy86THUBTuuKuvd420f3RAFmRYrLj4pqpxhzw/BX5+19kplbHVtfp
48hX748qJnwLBhP9ANObEWVhAQHUip4X+TkAgSKoHpk4Xua5ZIB7kDqkryIIHp5jvDNPx/ycmG7z
aj3A5g18Qiq6tHj0Q8rp1gg2M1QQL+J2m4zErStIo63g/isJnrwLG3BsoLqOOxyv3MaaROPknoZX
+IZCgjJv9XKlynedTRrUCQ0jn3NuVvSWdLc0SJE1TvWKHvSfFAovufO5i7ohsH3cRq50NJfEgVTm
fJguXewlPBRz7iubHCxNDEue9FrYOztuYRjRGg8RYay2hMGHCBitSu+j7zaoRUZ8TfdSzNdoXzEo
m4dcWa2HMQqI4Q/pMTqLcppRs7fjjJCy+ZarCMHTuSggolTNGxlVfLnR5mE0u5PPluYthpsbqFI/
hit4tqjwxU/olDPFGu5UhzoP0MI9giZsKcaZ0HH0CvcHRwGBZYWwseyc/JwgJ0M7uisXgDkL3NCH
lb7/29VrOSRaZROeKezMnjbTWr2t5Vw1us7HsbGittdNFIdR1jULhvWdwjOOnDuz6/zd9Zu4wz4K
SZ9RuBTW570q0QOVJhhpu2iMl5In33KXGw1FXJeBQW/IvhTRN5vPojssq2hnbIVjzCgaEhcwOgbP
oQlYYJPegEvPCrfRAmXiAievPqy0uk0EqOicIYy8BqkCJU1L2xfnejiSOOrGKPxZfJxlvsp5/QWk
UW7WyGfXv0d6PdgjOIElgSFT8+jWETvTwCJ5i5M+LUZJ6efeVPdhElmhTHh7PmdkRscjt8MN1duO
57lvlj+SeafsriptQvdiHKNYyu8pUwpf7u8Ec0gNBQK4ll/fjrkIUmJ4v9c7kuW6SqJsSVeCVG7O
iD0YtWAZPQxNOdibkWlLEPVzvg1DYEtq5axtsnd3kNJums2nx+NUAJVajGBVukXx6xTkKHl3ND0C
NH/Nau5+u4IWL7/ZqRwSvArkI3hHBWF8R3AQWQFGkgmWf14+7BTQvAqH/R3/4ZkMz/aN6o0uA2bF
FdEaYrp3dU2hhh8dBOqWXI28tAuxSMHGhy7bKCVhXSIidY9jY6NsDypLiLisrp5dR0Arrxw29jGW
r15cBoM92qeqPWXzhiMivNk8nqGyl0FnLSFeVQNU0Q6CXb1gmX7cv1TTRGDPNu6Lndaj9HRVam89
Embo8sJTMP9ow4J9Akd+WhISUQM62zokGQfreS8Fx0Wn/Q85W71XEsuYKWxqj6TDa4FVP9IqCueM
UOPGZgX4iyCTLtXwk7k6vAWto6YfCt+ha1acBH/kXrubCp6FdK0/njr/0t4DGeN2T98i03CYVKF0
xnPkua7I8IF3Amvp/IO4U9N6+B4RhxxtUXTcQZ+DgHKUyCUcsTZXdUS7yghUFd6Emg7928HlWtu0
zljq+snqd6MYehh2TM2Ev0z93bm4Adetth6aJ4xzwY+rwHXibTCoHtGUrgSj04SV2cSapgVadoFl
x50H0U9TEdLzwYKZZi7LzNNUsUlGh1PaVzNQWpvpqaXGdtfRvERDn0h6gkhGrOwMchnLxuNhl1+m
aY2xDv2mbwr9hta6qOxgUl99CY4gDMfTtrVcIdwznChBCXPKy25vErvokx/Fvx0fm9kQxItP56pV
oNCcWvMEby9jKPAI7j9KB/UaYfIOCF+nEjbgCdBtgth4JglhKpUE7X+1CMoud18WXBd2egqIS9N4
UIbtGQV/GR4MD1Ukb1Gp77YvbZuUhPGnkeUXRJ0rw+KUVOKCK5m0K2ZOYt+uXRH3UTfbF8K7RVxm
+MWtlvZse7rOsFYSPWNLDUhfsJynR9XFwQ3D+OgK0zx2cp3ludL3xVnTazhAFSnKGjfDheRbrTx7
pFdhgX5/cvMSLePp4d/A8bA/ZLjzev0aVj+q0FUvO13u1o6vXk+r8dr4lIwqjZhxcGbaxpLT3vFg
NSqc/pK6HQ3EWuKgTsW2prbLiVwxiiF30uicNq1NxA5HPx1iZqVVxUekH6Bz0tofBbr+wyqPQBZn
VWUmETQQ8FWVvRgki4s6c+gbf/Ei7OgZ0axVior8Hv9c9PHtbeQqH64mrS7BEdOqfhlkfV3ke2cg
t6IVt89frtYfJNSCzM3xeyf/VV2cwOztVhZVB1Vp7JgRDo0VA2e6dTK4ruUXiQdILUooG2JZWchO
jyV0lTTQzKv0u2MdmlSw7f/GgNDkknyBEd8ZugDYMxhIiwdV2WoF6epjjp32KU5Eg//dn4UkQSOv
zJw4webzDzSHwkkj9YJ/4aDbB2NMKsgSZGG6g5de+C7MlK1O3WyucfX+M/J+Lvmn0lvrPJpG8y5I
Y/3raSYxDksLmxbdjwTugV8TpMaGki37WxR1KlpNnQkNAM8aCeGQtpG5Z7Gprv7c+NIO//K7KlfS
zaPJFb/iGkfR1wl+rDqzduiytUEtVSAubyhJ2LU4CfvvnSG+O3tuOx6EJVyVhtHQwth4N661rQD9
mrSGh6Hy0Y/Rx1xNJnXr5lA7RJ+zVRIRKbaebWbpdeJLZZaaIPsJ9wWukKU6NZ10F8PEL85/cq1T
DNTiuckJtiCayv9KgtwDyc4vZBh4tDKVRLuAktFYG8259nhnqj4eO0Sun+JxPIpeW9isX4bUGhqo
ll1+WbO9lHokCmE3v7E2nwlDPmLLy8F6s5t/aI/m5il+dyFgCIHHkYXM+mCnicCoSg9gID6gDlck
6sq2ZvpISK5TzyYGZ/JPKjQqiWXMjoLrLxEF/OxqeEPWmy3fKevZwUkD/3CGoMcIRAx9s8LMvFyV
tRKE8AHTmqc3YaIGj9O9bP2fz7SObn1Rcx0QrayZU7rR2ckQaibvOdmlvNiSe/hLhpuiiQP9s5WM
7EYOxi6FPi5PEfj0gDlajYQ9A0RndINt6CiqP29L2px1472q/waatxeKyVrknrYnif8MmfBF6rmH
rUL81LVMkD/PjtH13KOprJletEs6qgGTD6ZXSv6fw/NnrIxBd0tCW67LCDcbLHNW+P6oGHn2OOKr
ybJhDeOTRR3AGj3ndC+59LfTVfILN6g8cy5FyCKCAWEVQ6UnR4yFcxcbJ7gDL70aPLpRIRMin00L
Yy09+GwfDt86Wrsg8w12ytU58X6x3yrnH2fLXaTMWyKw5LC85ESYDVVeZp8DiJ2nQQLOT+4XZ8Fc
+ca2BT6Wzslbbpt4IvW8w6LFwdnmkvnojMabl1o+lY/lq6GA3hwGbyh7Psq6WU8CPfS16FewlZoK
bd4C1WHbOehdyQFURsYXWLVfWNQJejwkM++KYC1YyjjoyQgqc5axe2sfOfYNOFA433tstyDV1yMl
QebIsSctMOZZiUc5jHpbWtQGj1cZLrk5TRqpCGBfWyrL4uMMMGDf9LCt6xfYPWj/RUSkv+nbBwbB
o45/3EGzMypJfLZhQL6Yrm/UDa1/32/cgCGJ5tZ2oRrnN1LfqMWX8OdqFpdG8sGZxETilhfxdK3o
TSYqlrdOLONrXxJEaJUuoPGGoutYKQH/LxOAn9VMC9krG2zHDJFMu9P2Df5KzEhzRU7FxhNu3i7O
R2Ja3GmQtrytDMN/54znQ7nYk3nFkc8nqPqDaNGou+SJlqs9s6+Mj2utarlhBexSTpqb0sXao4n3
/vKDy7RtIee3CUjb3V+L1jjWgT71U+UCHdfKiIN1+CdU1gAAD8mp10l1kauKCwhN21alRv3kmP1B
tgo0FMYSS3nqsOQjZ2xNK+CVB0IjbEIFyTGxVQBmoRqP0ixmPvJYBuIKwU3nJek58+gr/HOp4RKZ
uBtaYn+L/LYvEnKDEghq0BjIOx9Z65PWe+5lUMQzvg8Jwj2m16aHaKEII9KT864VvnJ3knfx5yLh
YAzizy/qomk2Ek2dAnbjVinTfFRa4htrarM+0rh7o+dhxDfKBmzmYLFqvdfgTkfm2tQqFrYpc4Ua
BmEEeiSbAmd0S7oO9AbSXOpbgBK3lfXGG4CRtQxDjS+kWb56aXr0XFHTQIgdxXpecoehPcaOE/iS
K+AODxd3RooLdNzYBAri4FHFXAqXTDIGDH9v0s8qWCzBTeXkbBnGU35eyUXtxF1uyOYrDkVlAlIM
DAUSQlv6c2Iqoe0wbeJ7wvagfBt8HK8YICTLUTeFXhcOJLmayoCRaovvKfBkDhHueezzBSz7DiHf
+T0j3KjfoEOBsqZcP8d49PQCe6OOuL0FrNZcyo7NnblGfxCFQNva8IWOByf3YeV3CtfYnwjeVK14
YutFYZ+W1/DDRsf0tr040+IXVGbJEKJmil18CqJGX7V9kai59BYr4XoLGocCgxsVdgCQr63NK+23
rP47OtxpJpmJMHipUCGV8YaGkk7267Qbll3YfUJAoVwDPRC8CLB5AjyJgMMRJLERuu5Zc5ebD+5J
bqpzJATXQUbMyc0KQ3bQbtGYWVozqXt81iRznoZI0+qnkLoLWxKWOQD8sbDCgZ0kx6q3eL3hfbQZ
wSGi5mbB2EuCeZKas7lOewObT/9fqTnmMlCbz1Vhm85QMPliz3YImPeHqlzg+SevTfW1f6g6o+4/
/8nfe870Ka+Q9lxCjEJVMFBF/7gWsNVFJkUAu1RgoU92e9AGmAGQE1dxFfPYAiCMHN+C0zGvXEHs
qtHt9b0nD//PPNE6Hlo+SGnCbhVkk8La/Q0F7BtKsFgSYJiFZ8dJEt7wT29jX7qPd4X2O30fGADS
JgLXH4uyxVgbQDckmhWrSaAoieZxeDhbnPjnLp+SrMY64pRnsLUf71/xBDZHLoRrXQFSPbBzfPOl
yBUER/rhxRV18z2+l8alFQ9MgwFlwpA5klyoqTV64gIkXV4X8zaKcfab4JucL4kHS6fbi5HWS1kJ
ZWQ8AdhW6+Xcg94+cJc5vKkkZQs0b9GTKhyZX8MSvBnCVnAfbKRsTA+jy0NWFGXol1RrR0vHpr6/
C+dER+xgJkaCiWHZMGIbmRF0e9MsfYYObXBAxsuI8mjqp/QjQYMeYhNU/l2fh0qNL7qWcGomPGnC
4Y9TdG6UDbPzV0ZF9t6tAcgJ8nycIRTrS+yDsd8bwY23uPxfuWGA8N8y337VQXfw6Fp1CWWk4WiT
zrG/to/7yK4KxEcnDfAQqDXvNN1T2TWALVEmAY8q9hFFcYgMT+0VA9V/TR7HBoFZ4ReUY9BTL5tF
1UcL2FyIjDJ4z7iHdfvtPPIad8ZiY0JcSyK/pTGUptw1WWPlcjZjfDpApX7K48yR222/heOBmLAy
APbqW16DtCBCJWvU3txOlzEzosjBHwIrI3s/SKDaYbwtK+QiKZsSactG3ZCAUShNG/5Dwd/q4typ
7cAc+FyY+YsIp8Ovfi8D8YTZzAIaPz/AmB9RLGxJ+OrQsryRd/UbwBZ8ypY/eQa1qMqk7sqv3xGS
WKdWbdpw2d81XuA8RJoVzLKpzdgnxzSgkx3uht7WbaZuSjx9hl3PSIHK83tNq8SctzZsb6lgqyiD
jTmejRrHmq/GP3gJv9yg1ikf2qNXNb5bciGf85RSdjc9F+ixajsZ9M/H6+gDetayg3BOYL8xFwuY
jsaQFJXa7vxGGrUD+g//IZKbdHeQutoRopbZmiMxFApPgzVDt2aBqkCvHn3KAlDmUNm7dElYEx5h
umGwslb6m6GVPcL9vkfCb6FHXtjPL5s6hWnL5uFCY/O2S3L3KkBLOUzSI9aEIxkc/zp43rTMcpp3
0wJYwN8BCV6W/IKaD2WIA4XaWMWFHJjB6vYKCOe1o9NqAdOX1AFLLb8yjJj0etfyvV+Cylv6bJvb
GDHoRBYUqHbNV3Ujj9F52RaJu3hTiz3V3GDrHIv8dBUkt2elaeu421WRHe/mtTqeHnJN6+HvUiur
CsYdQ5G/9nj7QB0wEzW8OWRjF9WZyyDokenswjs0b8P/IK8X6DUFq+TfJdTUxCZXGxab3m2yXGrc
eb+Tgeg5Uz5qSoso6UPu0PEZ+OUYoQH5fNIqI5oZzG6Sgmd00Hs2Vu8sG/7X1qitCEIzGQBudVjx
IoU1sDrjiRQvceiVFGIlgouHeYeIIbRi4vIJZhXMt+zQCMKk1eUxCiYOmDZG6JWrxDLhncEKso4Y
mjTIJTmE9tG6rzI7jDbvIKXzekE8LG2ql5G0G6mg9dTEp5AWT1vOho1k8wqnaIrMYxCBJIYxcqB6
bypsOfRRuUFLTtu6mAyaNIJRcCagBHBxnZq1bfURuZl8YP3mLhX7K+rIs66oe6UseeQzqZPyJ2Lu
k1SkEwZD+rW9GKyrTyuvUHbiHkQAcRVJMdbCpwLWhSIdauk8Uc1WtfVan1dTUd7hor7XCr7KGoBT
WLd2W5IAkKjBq3hHESfXkAF37i6DLQAyhLRvWfWWwr7/wcygzX/m0mD1GC9DfqtuhKc6ieotxWfY
voHAC1xr6dIQKXjhznx3WvbGkUDNWE7yAQbm46bK/Luvp3XCkF8bnmusH98VVCQP6NKlof/MQpdl
8ukqNQWIwZkqf2xPT3g/5OwwKVVniuiudMYoPReiftFjEYkE9R3mHTnfiVlp6vN0F3pV+cuETYhU
MFXu+Ud8Z1jqJV9LzAH4hdhKn6fxV7r4+lWEz1hGup6otgcwq+4P+trQidVaajr1/vvfz8Z1V4ck
K+SRf6dqxCLWacNqWfkFdaYCo71t2Rj0XBwPxUhMkfY7qRcnwv58CvXDBE1F4LmcTqi/VH/RJdNW
190Eai+La+15bQt/6IlrlOOcshjGCouBcKSL+6JO0MHD7sSFcLow5G2LyVHZOX+H0IYyCF9SpTJP
xGsWjccM0g2QJfcBPtBUKk1ON1dxDRUyplZPpDRlO6unkyFNMbjHQHIskoO2R2CbhPb0Ow+rMNB3
ThrkoG37NONB7VibSFe4/y5NmIBVXy6G8zDwZ27MHSzPi3rRNgqd0dM7vkv2i+D/SiFLOt2r9z0E
8gp2QTp4bfRvTifk6a+xg0eQLENJ0rnv+0XqU3krF5O6Rble4yMYgDhCzr42XHuJ00Cj4xr1MrmW
V2NgtNiZVaSpERST5vExASswDgxq1y7lMR0+d1Rx/m6KMu1rCp5DaHZo/z/oHdQbBj469KUUOylt
JnmMcbjHviJV/zaht8+JEaQ9KJpyUEdgwrIFuUqPhNvCy/qWRCou9x/VUh+9PPTOSsAdh72xg/VX
fWenCJoE4vCByhngJPalP382CXdQCUeeHHkpWFhwcnEL0NhhxzLrnjpX6IkuCeaxzKwEJ3tURMwu
K/gsYOpZA/6NixNrMXh82onlrQGe2h/Qo6YHUScTiuCMxnCB5OEGQSdDkTsLoKUUZDwg8kXznVjT
ke8hsixF7DjvW+GDLwv7kqAGxbB244k3Noe0B0u3k7rxWkvgCF8swpj9HuFVFXKcpEXb5Jqc2q7b
CNzBh9e03j20SbuxpK4/PIzrYqPeedQsZgMokqHmqgDj8wHBfQnzCIxSiffvB7W37oemX+H1ZMK/
ovgLTwzyZaWSYu2RRjdyaPATTda2i6K91Vrt5kMmb3zmqfVZ8lMZkG5CeaexUO9yt+atEisu+Iiu
rRm7VhdoSyW8nkWfzdO84fmEJUleJj+NQtXdPw48psvLIQpHvQ5hbWn11ICkfaul1sFnDA6VXTlk
oI6VGfOK//ba6WyBojln4rN6qY5LT7Et+P11naNJaAuy5gFvOSMkYb/rKD5fYP4Ir8WykA4sz0/I
83ofoS3IatU7q4X3labisz6xTBBvP9OMJ9/BT9yjnSeEvqNeM2R6c+4EE+PZhgEahRF9PsPy6HEF
m1ltVLOk5KTiiuu6U7bHZIS+Gu2erprv0Cp28swT1vlQcjiFWeUhW365wr+EFAamnpNnxq0vIjWJ
dnc3AXF22dtTlABucKvgcd+vsMX8WocE13M9OpU7RL+S/ebTFxsC0SRUb2sjTRRSkU9zBmW8zkQy
qazrB2xlY1VuMQCjEMkCizBc+YgNXRTojHsQZGwfsKiln64zzN094GUoFcAMKVR5xkcLwJLRRfP7
/hDjK4wOieaT7AtRT7WgQMZYx4fKWXXQsq9veEBQOgOUms1TUeeTWF3b1JV9iu23XGWqVeUw3zMF
l/aS2mS7+OWazEJiwYTm+cvYoWaywXSycKsfNGQnA+GmNzRb6ZZndrBDXRpmS5D2ajhWSWhXXX2z
FUoOrTxEvC7Wm1YfL2ldmFdxvPBb8bCIjHtBTNfeHTUd6A66SSkIqvL11Np/2/RoS11Sn8/EdHZ2
u9eToTHNaLjRtUq0POTYM9wAF/wTroALNMxbbvm/jGylI8x4W3jB9TPj6KqYaH8nbFZvNsKqIfwG
SxthAeN3rFX7frkwog75WeZdWFAKo0MI5rn7r6v9aC0gXQUc3z8UBCDRf3NFrlE++PQwG1V3m//u
dkbAT667t3U23ikh5a3pYIah1nFVGvK+i/0JtBx9jOQECJ+cs3t0soL0/e9aOMfCDwDFie5gct1U
xKK/g5TwgthEH7K1yNujFqjb9W9GDGPp/IRyK+Mz/pcY5QmSoKUha6taAGBG8m2Ax/AwPq+no8di
D4HUDLgGbInZmk4F8dp8HSl76avEcWJSP5Y+zKcAjCTLcM5cA85T+v1UFvRUGfg1RK4X1IU8tJnT
kQQKwCG5u1QtcU6uN/pAyynPrhTMkrJ0zBR7VoNv8UO+e0yEZk4dCzhG8qvDSOqVEgtjv78z3cT3
3bGg8mPMxtsgmxttgpFDVjsFQxmjxqBMtBUzyf4Bv3MuAdvlP0516eSqUafmHoF9j4aSq6VBW1No
biBmL/SJ/8OcGhVmt1qYewvnhsbZ5kPEUR9upvuDTPkS07NRjWmkq2zKUmFwd1xFjLHUd3UK2Y3G
UnuatiUhDQ2qNNuCHD+FXM9h+lzTHrBus+bjb0bRDw+4duxFyRFq3um9WFios9f6r2KmigdnWBkB
1IDAt8sua/0HkLXZjdMUW7CQgmnLooDgARF2eDoKD8s1HQoRTRHx+S+QO/5BKd63/Z56aqMzOmFz
yUZYhMhlDxhNxstraCoErUEvA9xAEd11GGh3z5DBoBJRNiCYqvjMyak9toxZjI/vYeDigY3lmGVp
9No24BvI8q5jmoXPPc5vnO7zlMPuBNHHX5OjfKDKuNbSeuHGL6tzzGUu5F3HHs5llLW6xhjtH573
f8+AGP8BY4exbx+uP2CAgaD++D40+1zzCgCbKnsWSDhd8tDwGWBRQZY+g++UoBvkb/1GCbtDZWQ3
90WIQ1q4PrWxWMTEj4TLt/U2QpbhX6ZuB/XsUe5t44RiihzxaeicOuN61PpnoI8GIwuvvtRJN1FA
AGQDy8w8cO4yZeTE3ZmBNTqC/yv7T0fFjHOVRm9B2eJf+pvO4z2trQb0wY2N9SlgM3HOPw0jxwgK
piQRfq/oTljwKl0t/sPlS7rW0KEI/+K3oXSMwEyjLCnd8ACMxL0seQ0jMMBt0wHL8HTQVewAvkRy
xrfxjvkyfyvkSf/e5zePz+8PxKSAkzNoUKQM4+jcr01qGkU850DHnIfRfmRKrmLBbDEvwmft9diZ
eP8q/BTWmOrVjlUbyeVzkO8hJFLuC9FQrLpU+vLXFmZMDLJXpUuf5+GLq4GiOU04fQmOZsVELx8j
ttQttDQovAVMcnaucQrXMe11dVSEkLt+v26pn8YhUiLvkS2iMIXIxK8fztpNzglNHZLNsVo1Db2c
USZdiPVKnihYAnVg2ICcsZHIigdhBVv1Rkdn+SYslSfvfd53k3YdZgF+PttAMFCYsLQV2F6ivSfj
jSqag2jgiMACPql37ViR2ultNAX2OAIYcMQXupZqlWkVozc1mtgKjyKavx+bnDL0xrw8Hd8kAJj6
9sb9LqQFA9aDyo220Gt24xivE5rCXAnJ03Ujo+wHPkHYQRg2VO/P88UdloRPTK0XtDMcPACYcyhD
vqpF1SuAd4pxQZOpDZoMN74AgsSN1/y+KvVswIQKHvpyUI0R/iZW1/kB19h0IeoiJv+ynMSHDfgM
bR79fHOVg6uuZwNi4XhNgFqPeltZUxmUJts9gemRWY00MZD+WoEwxCQ/kF6lOB2oEwyjcG/id7VW
+8ogETD/5B+f0uBJz0pfA/jNkRVmRq48Ze5jwerQzxHqTHRfblHe4ek84unQaUe2PX4sXffunyMB
5G9M5pjJ8ETCBmZRa3OwcMccrzVNvg0bnRYCZ+yxA47VevAk/rTFc9sgf/HLDuGkS9L/UCqyMFUr
37tNziYvu18DTtbnfqpUSv2Rt4YEcU5+gwoSr8diPJgMR+l3QmnOANb53qzbWPjm1mdmqXVcxY4g
sfT3XQA8iom5WwkNrScINm2WQcGJsMTwtxU41WeRQfMzzls75iUd15/b+xHR0WifId7vqmPBWMdI
Dk7JFUkA5aFVZvskgBKZs9yFep7O8ZBUkZdjKb/0CDgeSdswT5uBhP3x+pDxVf4OYO+xY6KrQtwH
IURT+u1hngdBwgfIyzhl53s/FF6j4xbA4OI7s+VtmtZga8T5PGkAJ/kGSZ+r/n2cQOpP8BcMa8I0
IF36Bi8cpyVlDJDDdI6vozH9IC0L1xmoI8ZRniAZRLXjT77AxkghTY/n+sw30EfLSVylJWUeqKjl
Fxqb8vVoUA9EbFLRk7BQB51cr7RkFOXyMg0bf+4zcnaGizeGDBGFcZ07rB31W87mY6+AXz6F4qah
J+Qq9rOGwNQX1BbihksY+z6e+T/IwqLr2I6VoOYYuDz3lr9TO9b6rUqUFBd9j7DuqUBXw4+HmZPf
G2JiTjZp2MUhFvnon28aLK/jhX/s0q2lYFOpLpQeIsjHajuKTtB1nYHB2aO16+DNDqw1MSVvjr/Q
Elj72hP2X3BNZ10gKZFkFaO7OZEFs5ACVXnXW/fOT7dpc3JovPIbdhEiTZm9ZPUKYQwdXzIp8m2Q
IMXwZnlzjeXk4m0eP9+SGkpuaAYceQN5fCWM3LbHZ8TNoP2Rt9scV94cvuYGcCdfvs3zSXY7b8Nb
W2UBOtFD0qa/1v6fveplgajj1K1N5uWw0tyuKJ5MUFf5wqeb4HUi4hb3oUiRIFiVLmBSy/HMDrPN
RB+i/IPhAZrsr6EULDUFM0B9pcmW8FSCSpe+yjH4szFMys9HfF60xt1O+smfxkt/9CDpFAOuggET
JuKd9aU99x4eLZkCcEtWOY0/6P4WIKKL+iWCaUfQSG+7WV22DD4h255vtrYVekCTird3gf2VbuMi
5JT4VpZnTck5kPeyKijI/SA2cO+sWCzb76wxQR6d0mSmZakKaVBIzo1d+idtL55H7tHIUzNG9S5J
aOUZk/91YBPxRd6etFUnafsLq1+LmJkA40RQgZpJkV96gcK/rOCxBcG6ZYMk77ktGZ9YnjIDT1Gj
SnYiby4l58Q3GyGrHdqT00KRhvXSTl9Pp527ikVADhCs7T6pK7dJ92RkqX92SEn1pPMSHdZWwBVk
Ovr/jd9AGllCyYtreiwCp0wRJtvprxqdxStjwsM/mSqozsrZVFG2lWNkNPjQnl+HDMw826c+ekl4
gYQZltLzrdqqatkVU/Qa6/eWRfKd/mkWSp3I+P8UXZ1moFRBVyrDbFA7rNY7MLV1fPsHioTxOs3k
fOvnZvrqcYoI1lSMb0D5ocVvFrzKgLoaF8urv0h+HSireU9yAIHe1rQGG7yGeH3SHdXdh2g5lWHS
jC/82xdEaRMqaY7b/6pTpPU/7gb4vIFlcHd9pz0Jyu1QcZgp9gO11RDkSWPoAO3ZkEbmG1lNCr+m
W5l+Mg0kYzHcKHcUvyVKSHIFsPHaDpm3WZOjkKf3mKVFyuR4Jifjc6SPnxMsrS/A6659d0YOlJRb
JcxA9ux2PKyRwnUzkMmWsyCgt4+2TFYZuUTjCFg3efZfMEkvnEfbraDtK56NziAU9GlV+6342Uwo
ALlF7t4nsuircbD1jU8WSQbd49y8We9Q1XG29YWwHMIxLZOvjYyp10F+HqAdzSsmP0oNzfBU6EtJ
QJMU7Q9X+bMs0bQhdpk3Ef3PFauZboj3Nz0ozIDiG0t6q+rgqpMIHAOWkHgOI20RLbuXhCZOVeOr
Jh2meZ9d2+PY4mNYHsqko8d+22tVH+I6ZIBMOeUgSK1ndEijMoEJXg+Vwh6N0MaaZBsp8hjGooo5
ebQi4pZ5Jyyi5YhszXNlkmWxsuK+uRQqm9JIFamBb+/Jm9CqkuwhRv5YxTBnfvlwpYA6WbCvPmqc
X7B9sok7zNNJSpt0dVA/cHn/OTpATQk9quzH4qFejbI7Az4zR9dporU/jH6gbC5xNQF+baRsKMx2
2GYtUMUfDFoa8K/NOEyl6BNW5UB21J3Zyvh0d7uIcUOPs0r41yOXeh0HUWiyndmuDeJ0mKDVZYCx
KsgPDSsC4PlcRpug7ooT/6oxNMdD5XlEYX7ZnMf1IgfGh8DbdddrMpu4Tj4R37Aujz7XJJpHrgD+
RCuJBVWpLRdpEW9aNfK1sir+tWgac+z6a+nXd5vpffJ3Bp5it8RQ2fsB99OYCGta9kfsy8TFypE/
6niVvVTCHl9ozalxwRnQ5aG+8QYpJ483KI6wv7hICbXehmGYx2CodSOtJufHPz/2yzzet1vN05Hd
IMrhv3/2f0S9t813hNDijZfAj094RfkFqh/U22slDDsKCcVgfe/26rICJAIx4eHHkIkTwxE8c182
XlDfYzjdsQE7hsi3DbgrYr5bbRDZxLpPe429uRnhMW0vDE0bE5p7Q+r/escGZa4Fq9k/534zD+kr
WbNUzk8iCrWZmbw7oAZ5/IQzqRK4aKFzS2ouTvAuFs91qEd1Lyr0tnYT1BPgPuicvVjLuKiAdEBu
XF9JQxlF6oiaNii42N8A/drUgYho24QfeInrjX1RdLvIbPANL6uMxegYp670ZZTjcqnZ5n9xSTDz
zeuaC9r6JVVjMzseIAYeh0Wp62TIsd6vEz7QBDloIQg48vHPXIyfP7KuZKB2+P416hqYmvXKlPdA
giCXZjiwzkKQqVLRPv69X4mTZXahDUrpxyb5yktdyMwUeaylsv4m+HmG23WoFnJLFMXlBUI83J0S
SVdVIFvrXlAF2Tp+x/WgfYEu6hrKpRMlpaRp3Oet4u7+RnWh4snrDA/zMqOpI5oBsN5ho9W23G3H
9kDZnsC61PF8lLcgQppsDJPXoiym0BTuN01smTc2C6MXO6NTozkd2cFWHdQp1W45kDhtq4Gag3nm
0SYZIpz+yGZAW1NxSUJs9STi48XaPE3OvjvisGGIe/YUvrAibrrgCkOi80rWsdJ86rswS+i7NDT4
DVK5sa1Nqa7XC2gQ+ymKEGpJ5pvl880axroj6kI6j6orf+YOA5En3qzGQ21Nlo6F2vgT12zIE9xd
SBgvYGemUwloVc4+IFQEJP+2O11L567Tw3FxD0b0fcU1SiM6Ne0HdbyOp0EfhgjeuJEp76kJOANa
lomxAZtQk69f/RgJHamKDtPVZ4xev8ddxrEKk2hY8B/5yJswBzqqlYTJbV8l+5FrIqDxPx73oFCG
ysWRW+OTOOZ0Zu7IJsQAclsxtJlHlsJglhhdHyNL343UBF4CDthR3+pF5x+cryMjIflmbwOuZWoL
5dwumiJDYLIn9z1Fg/uQkOJ8MWALemhucVcGHFhl7xH2JhacT90W/shkPl965CMIIpSaTNCJKOOy
UzDL/wc5mN2Q7BkDw5O9/d3QsP1kxD8Rj5CUG2REW9GegantoblmhQxExltHsY5xuSBb2CE9gnnE
AV33p7SZSDlHncxoVoqGGPIkHr1H4AlLllcNsUxviWhRxDcAZiNJvgn+I+Ii3PzteTL5sLU2lFkH
IVUW24rkf/CAx/0dkzsSNp6QiSsRbEa3IMRCDjY7ixO1UkrEbrICIaLT0SH5XYmBcQjcj+ThJbAd
K6zKluRKxQeq+CAmuRnIDcNsjhHfnyFWfO/G8beXsh8AbY8HxNBs4nROUB/PWIGni8ktlD69HmBg
7ntWJir8vWkJ3A4T0KSXLXoESwQXRi2KUGJi0dUROTEXgHyTUo4+78yXvDpqbdRvfedCDSn/ha9G
SmTmuOSMqEP9uNzpOnvtP8g2FUN6ZwiX5H2w+1oMLhibypXGieBDnDusGzq42ay9v3uqwfEx/TQ8
hlmNjGUE1OTd+35T02mGMo0LtUn5r/eUoWXw+PLdRSx4fwdNOoOg7eBpfOA8qTuzEYhNQmZ7iQhQ
rDjs0X58/DTbb8gtx5hYH1DMTY13ukk6wAdtiN3aXzQH+VD8yZAzwBNxPa5BJ1WCI8Vy/qBB/Fuy
ZjfHBPZpjypaWxOcNWh4S/TVfEv5Q+8ITs9Y2PPWDAGhcEEUpqHJgYc5VpGCZhqHEvlYCYUh75WP
qksRPu68yUULRrjF2/6NXejgWC0YM7qiCDVb4HR9iAPobcmJ5xBbvXiUTuPOybgStQArbYdjiIrk
+Y7m3xS2qgll7akuQRXobI9dV5MDwO1Jb/mhxZjvKiE9qm6J01ul8UeHS0jsHHVXOmGIZ4MwTb7a
ejeoY3LW6xA/OmHVSho6cvPA5MknxYEm/Y4rXB5d5amFLY0kOQPbzsZjWsSoEbDjJxfIJQIEjs9o
1yxcXBnUmW6gpS+tWbWgc2T7+ofCfihfra57ffraCCOYKnMWn0N6bLBwQRo8UwIPY03z0d6j9K9k
HfQ52Dhu/JxPBuhOat6Wr9Cg9vOZb/yrNq7REgozzq03xo7AsEElHdgyvHxFHwrrMOBMWx0mOird
Ok0jSDbUvuv4Ul3Jw8PseqyaiMs2EBHIvSksT+CwOJ0XOdECQoJxfxcFgWUHoHCxbilD1mfhUmJd
QNTmzM8ROEPp2IhtXVi+0DSWpNj2F9z+alPb70p9kX8xXEhiNlP7T8C8qTUpLkf0nFME4TyS/jDy
oP4HsgGlyfiTncNGO2ICIkNqyp72In4SkoBBO5lzaa3crppRagBw8SbSlafzlxW1YA+5RrRN/56H
7gVjjCvLWPI51xbPvti00d/ikEnlK9EGq4+hofwG0XSB8rXj0oQMFSO2oRM3ZeHWcG8+DsLiZDbd
s4+oU5p7G7ltDSGGFrH9YPU8HNHswgH+wKqi8UJ004aJE722ZRGMi5TdSDMeFGblG6XWoohzvbRo
BZOBP0ZGbPtznVjxpUoYNwT7FtUtCfIK9n6ZWvk=
`pragma protect end_protected
