// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
K3jK2OS4RT2A/EwTswrse6Qsh5Tn37vUHQFQsvhvA3P97dfgItqmBZK5PRM/voNS
qNc8G2hPsNefhUjA1d0pXTdJVXzlqZprc7RUXnnNfG1O2bIAYASZNBBnDmFU3bEc
T85ziwIK6+o7cj+40I5d3tjKsGXOkHG3+3bgIcwe6KA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 42576)
2iPkkiXBDShxjnWaFWaXLIbBA1JBonAlgWhbdlVqWBsnFOn/yp4DxQps8bBnWmRq
US4qtzn6m8pz/F/TZEYXtFIiUP7HAgGUjmEynlIs62wSWZCAkGouws004CWuIF5Q
Tv/Ny9DYKhsPMwE+y+o/RT0FN/VygeRTePLE89tNLsuuYbTNbh7oGyUDq7SNqadJ
/KNErUsCqyq/UMSHbyizbuvLy0vV/IV06MEbG/CEJS+rqVsKcFthg9mhm7qFAcJm
CgmM5dZmYjsPrQD6wyDJWuR4MA8tvRhWOq4SQ61tC8gBj4x0Kdn+tYjjDVa1FPlt
R7zTbxGSZysYOiISTZsS8lloU2o76rtFoUSwG1RImki/0GTbEEa16vLPuWuR4Q8V
/evwOX9Zq+FZBqMNJ6bnrXebD77gZOZPD7Yw/X/gr/V7ip8LyXQ2XXRuuq7XXRYa
cwtH4NjYvW7jmSCN9XVeWGyg37aZN5Eus8VAZXiPjjaY4AhP/KXx7xFlfN3X4K1I
/jxQzhEKcOL2/+86yxIpRORwN+yVLlK4mvzNZaQf63W+PopNCtFso07FIK5c/59a
xgNqalX9PAEjyHWazHLkB/w3SRzw4Ii+IMokmFvGPzsdSbU/arn3U2s37fS7LuM4
HaUHhgSCPodGPrtRit7Ji5jqm1hqwT6zd+U/G2bYkAHWL28RvZTg9ZvV7AwgrhV9
InkcFikdR9Luim9GV5qRRctBc6BmiVxAhBmzc5z5gTQFhxe2eYK3eSbsFeQaqNIK
hV0ldy2aMgCHySNHAr3VJhk9Uou/syS4k8lBkdpGs4VVXMW1zXTYz7Z1Z3veVHe+
7LpK1VbQTR+QjHomIBE5DpwlHsZOwbVw4Sivt0w4Pc+BO/v0FfHDPJrSbNXlzVMP
pZOlKHVKIQ9yiqLw8WhKAfqyPDxIbWrZUcRkeY5QZGnk+agj1cIX+PhG4Wa+QUsd
qDkcEseBGjUvtvJ+sjTS1V50v3X1ObFNUNLVLS3l8fZo0YfBHuccBkjCqpbx0HHs
TfmtJkcjypHakqrL5xOonBIJn+f6RYgjL21ZJ5kh6MIAYXiqphOojyuAKTDEFe5L
lmOm5r6d1WQtQSGmqBYqxDnqiWU3wSAnupGmMHMvUl6uUyzhxKz0Na9DnUkGsfOu
dbMmaydUNFyqFtIKeEKxZ+7M3dmG6NMEwgsFc6WVHzdFvtW0UjDKQ+kzuALpAmw8
wgezv4zIvUbHlxY9r6Qkfkx19dfrEouq++4HZpEMf2jUdKCWQGnJD7kZCfGoofgl
MzGWejwFzl3Ju8PigyRox9dUTi/CDtEw41PQRk+PxSeJpzXKoTAScM3rFDJb8NFZ
Xv+S8Z646xImzP78VEl2nJQ4Y1r5w/rw6Z8zGqam6uilKBK1tqsNwkOOELGWKdg8
eCv0hghi4pGTiB8o5gnNAGGR6wnE4ax5dQKK4b5uw552GVWcpx2IaY0IRi1IABd2
lEzEyNaErZaq/clC+cltuL1szgMTVXo6oh/daxc0R4lkPKSAIOwnTMvWxGpkk9JI
ireHs8a1JzYPOmmd9C8kPVjZf7i0pytUBJQvFSHvIsgYoVNQt8ZoqJt4cZuDcAo5
SyYix+hIvS10fvK7cmezag+GLlhqGJlAfCSqVdBtTC8BCXLt/K6mXPAszy9GzNHZ
mKj7VMlTzWbS8yO8+JRBTL5Eo+T21MWm5Z8OpZu+cS+Foi1UMqwrJToa5/rAUowC
jUagr7zGD6iY75MYvK9JgheDz1t0y8R7ZgRzHy08vfowz6Sq+COKIDs11ceQs+DO
gEP7Ce2CJEK+jNqHPwtfZ7XJMiNQM721XJeAKDrmBnctmSX4gCUwks4MV1L5TPlp
MfIERn1ZondlwsPrlLnHQE4Ka62aowCrraxSjF7iMzAKafkvFX2K+ebVQuuvmSG7
3zu/TOmRfGy9IkcWhI32uhOhHEge/I6STnfwb7GVxtnTGs9lgftC/CU8dd1mUH8R
/qyOo5aEx3BUSr0VEvV0GhIS57WLy8OFQEk9kXdS5/UCplgDxU9Yz7xK1Cef2Jn3
y+3piXT0o1FFf8AABdRaxIIOZoUPe83YjcfkJQMldJjwBeG4azC4Ixffi00q3d86
bRdtwjjso0h90vCRzNmCPlOgCqsnoG1QNu8VU2Q+cI+kjMpc8X7y8eW7fZuXQEp1
/WArdPSLAN/RFS3tiVlRrYLM9GHhwiWBq2/XBjnql9/a4nVofrihE8FuCM3hA47m
cUo72roEZaKV9rkaj3A1IU+iIWxcO36Fo6sUa0GyzTDZYSo5QAG1HbhSfcHn/Qdd
njLyWKBPa2Gx45pG8EO8Kn+qyx2WpH7VJT4qXtRA8eqJoRoGz7sZlAJoUqFUzTOh
yeloLfqnjXDKq7+aWlhsOzZJ4sEuhx5i6dTA6TUqJZSvpwwyKHco2SpWnurfwjzC
AJIa2lrJc6kjtzVsEthP+4+32D+gG6kHBxj0OOFGNI+yovMMvlJEcXiMmw2Im1f6
URz5k2voEt1ne3eehZiPLQjkwnp35cPxuv+3D1uxIm2jUPkIUTJx/jLT1+LZ4eTs
mBCTsHuDxlK5NnIlKwhZXOFVC4vhJ93+oRTVnuk2R2gPXBHccTRZIQukbIP7ssg9
W78SLIkHhD9F2FxO94SPYc4Z6fmKTw1U19JEiBJjWgA9vBs4KA4/nboJz9o1a74C
C3S7Rsl5+hfPwufb2KjGE2WRX1YpuRRvWdpYXb4tZsWjEdTvl0+dw8YmGb4DTru9
Pblh6uTUJCin4AvG0EpQcUr+SMH5k0aekgyjnEWvv8vfFnUgb7xNDi6IoLxkgJ7i
hYa8NGmRPhCuxXoFMBqAZyE3obKtzKgJRPdl6hnzrUnDxX6KcbCJe4f+HKHgqVXM
1ouOKommBC/fPdTd2xsX4Epjko307gWeShYB1zUcIOJ+pF2NBv91SeB4TmvxAdrX
BVhAKqni/KhQvQ3Lhr27b6YGJcQPYgYZBRwvkd0J33BzOmihB7ZD1dd/L7F9DegX
KyI2e7ZfeXjPCTOD5d/bzmpO7CHcCXB/rox0kvwX2yuIKDeiLQureT8jIJPbwIdI
wpJ4Oelrli7HU9t+aaffxH7VSpvKS6rx6/aUUkuTWy/AezQ0G1Qws0JSNJt/URGD
YxBRLIL97v8HH43JE3/7RJrX+clzqpOWvP0iYNkqyMgtbNly/MGd0ox1YeYnmmCr
hIdnXjKq87CL/eUN4zxZWKJRkAc97tRQm4kNDfA5yJpDX1z7YEOhmQkHolWxkq8Q
mpTVSHJkmYlfij2D/JL/CMzodd8g1SxgECZUl1t8wU5MBJpdgSbDO5Ql9imz64cT
Z5XIZqU+/LJIDXbQj+jAPdqlXtEltv4bxwU7bBfv3UAPeFQIiPU2ZVeHDJtE1m6H
3j1E4rFN6aUsiFz8/ewhyaw93gLohdLDD8E7kHf+u+Tb4LLFg4oynbC727HhIOOa
SYYCvC9TMkEYQeqftnvaaVCp4+8px+69KFvEgAqOyg4HvoDajL1eYp636NJhwtdC
6S/cMbHWzm205azIDWCwBdZS9B1oA7YpdN5gSbhhYSFFwsTRdW4iTsZ0+p4b4CDE
12sSRsmFNx7uKySJAxzoTmEsk2VmlB6TvV3rfLgc91NcpGxXdaW4H9/JN7LRyXln
p/OKtScuxoQ2RVu/sjCayEky805RDhj1KSh3wM4xZdE/KVgBWj5pmw+UUFrevVhX
3vlRUEhTPcwHtmvCdTSNTUVDNMZXFk/DDt+JEAI68etHBXVrc0Xlxd15YtOiSP9W
Q6MhX63dYoINgAH5lLpIQzImLj5JR8p4MpLAYLBOHPUaaTUpLtxopz3bow/8We0U
KSP4NxhZRFo9fyKHAIstRi9x24y0kNAnk+yzMIoM5veV0z852h/xrO/LRXh7Jnmt
HHgOtWblGsnlMDJUHG5wCt6PKObGp1IgoUxJnR8xT7HLKYV2YyTfmEnUDtNHXeAo
kZ+YJEBN5Q6GkV4FDUMaAyggJQc2VFEwX6nnaC3XziXd4NyQ9u4EfVc1XeLKUr2R
ci38nNc3r7eGh3XDj85VA9ETLaEjw/TQHZQ6v3R/umzfq7XZ8r5vCmH95HHpWmgN
7z703/WlHtq1hAGfoY+XJCrBFDQhcV4gsLOsxeQAnwxu8aWTyWdYrYcMn9u8t8i/
AdliBCoZTstgFDaX4Hkiz1Nvkd3aRKTSmqOLfzxx+sU9WlBnmsJmMdHNgBtBrqeo
FyhRUx4FRikqQ9XGVOsLbJShRnAKi8vPmyCIHkrKcb4SscrkxUnoBFsz7/ZHwg2s
YX3hJZVw4/xY0cJCgfFcmQAUj1qMQkEB2baly6Bt4d5nrocAkLYA8WHlnUPz2ubs
5v7BeHbRzCl1dfk73OYKUPKsiQg3BJ39bihUHxDGsWx4wfXx4F/zRzvdSinIYPAd
GVWm7ViIigNBiCDkG7DEgpNYUPHsOZB0ORm0agw4/RjvLtR8zuvdJCAHtpOLFl3+
j2fPJ4DnXJzhm9zmvVJuKjNC4dhTEdYA8Of4oWy4TOe1QL2sZO7iLImzY+INlyrJ
X0h4y0kzH34RmQ8UmZR5KnB4beVSQBZm+teobwFxSD8rPZ7Wy1vPhZkQiQfDbVPh
4ugGKSAXd7IorOITBO4k44S+l7802xOI9NGxFOH2/nFeHaDS2O7MewzOyhl13auO
hfg69Kk1nvi+zDRTh72U5qoHw+yIA6iE6xbKMiKXRMPkQ1JX/BWFATTyelIc7cLI
6q+7bzpg4H3qUBtcHtLP90c700wNYuDKgHBrRcuPzohNOWlJxNezjfuffVDOQz6+
BzJDz23RZbAnXOF7lpruTdI7xQbcftyI2sgzsaM6qc9vknEfjuzACtOYVTtkAT5J
49VOAz+2CPCtMpK9H/rZaeMz/n19ud0i8RMr8vlWKSiad7fbaTInpB1atL7V1NMs
+sNwwdQlNkGwJrEFGVVKy3czPisSvaWnTM3CLtwuvRngWMlS4Dkg+GzRNnWvfkqC
WeqXfd0XBoFBHYAi0m53uw5vVm2kTf48tNWndiF9h0s7zguHUaAlzMijsClluXz8
eRAHd4fWgsSvewq2J8SaoC9wmi0NYV031kVoITMc0p4htQFtKNcMo1T3ptr+uZSC
/l14jkqFuhPOrvwLoFuQluCmH7GHAUTd+X1+0gjVWZ4Bq25RH1GQwFupeHE/Dpve
PKzB61GxJsii3uijCBKNCbpI3pR0JMitRwgt2Jj4MG07QL76qtmcwNR26TzBW7ar
lp2lKFqEmBYn+EHl+GqGGRFGju4gXU9RUujmAcHewu48uxeQYWfl3fLuDmVbasnj
Um1bAhyzc4uHsFf3KO61dCE1XwiI5vWSy8Npz0EeQaiWr7CbdA5KP7Z+zEp+fZUO
MEtrshYczNKsR2ev3MG+RYqBYoQ21Sw1UP2ITMEs8knhWz3Oim5NVitTWRkDjfC6
iOkguW3kxDJ+mIxmPzweE+jHw/P2pTDCTnjfNpnppYDsWJT2nuxfdvFwRi7a3rWF
9Li922y5zc1wLNQ6IKFNOAZTZFCdRWgOvqRNH3Cc85K61WnW0j6OpBqt+GB89IDv
JoZ+Xibi1UeomYQGYt/ZEHS8pROASz4La5iIvIC5TN3EuL1OF0+oL1XQnURtQuOy
mw17V6zeQJSIjaEJShm076hlXE2ag3K3vmws6wJk3uPSpPBlbW8nxNI9XPdE5GsD
e7xZG1Yx8x/bXoJaK8gHD4vDrPrqcBAXeTR9FldDpi7/2k531O4tJIn9cCBFka6m
sJSubtNcrS4cNobnMw6dO0hzwiCRn7Bcqtd9eI1GrHpg8cd0+nL9gkyfNL1Gr/B8
AmXjvDR2ReoV5mX9AyGtBpL7UJRifrFkLePf2GD8rXdeKU/2A2iZnntZ7kNSlVoZ
0MYPxCK9eR7yDrcSqW7IMwdfQiDcE+/RAJthTeyQbudN6Q3MoxpE9mkOo20B5CVr
UCwK9Ma33bigiL8LAMBkMuua9XZpd4hYoG018QwcTSP11SZYoL//qBSCSM7F4McO
CJdrjJVSoIGP9CM0XXox+YwB2P/Am7/ZGFyj4pOJ1TWVD1pJTfvDQ50TRng5rL5g
pOXsrU25Lo1X2scYuwIhmhXKGoB71waVSzsDTLeYCYtWqRp2LP4WwDobjsRy/tMu
yMxUxyntx1AFUqpMkY/x99Xj35XJTu++Cm9UZOsq8LSGckcIF09RFcqZ/KnpW+Yq
HLGmBCftCGRyE5qO9iRoZiMSwdhBwcniNk7ULk9lqH+/6vW6cYdKBazwVpnEq7jc
WLXNYVbYzGNR8eq/H3Vn+8QQ+C7p09hJDHYzcKpeeDREuAVsIeAWao6XV+NgHgl1
a3ZmDzK72xq3CsTK69FUdyQfXR/4t07YkKbEcGvfFwSTyVULJwddeaa6iUpd6L+W
bYlDagF6OyClrDyZgyP1EIUXh/tMRJsRb4e9dv3tvsAq3lGK5jeh9EJ66do8HJb4
HpftHJFgZxqr/9JzvZrDVRqaalqx7UNFfmjAr/OfToHVPX3lW3D+YsmaaMRFGsaj
aJS1U/nxSpcl1VEyUzDYSMicgV/MulGlXTQMVfJMtrwxJXkJyELkXIA2Ds5FyPN1
uNQnkkO+qZpENCH7RJ0gmsRt8Pr/rqEzatDDGQyoDZPt7C0fDRIWHfrWPHVnFnEY
gbo6VTf0JIv/szDLtXUIJOErf7GRGUgxrEiWdaHEkpzOXQBlwZOnM34mGICctc50
z+GQEMBMSnXVaCHTnEXSDE3aCjyTetZZtLyGMNbF1/dOMybMNEx5AeRD64mRKEWO
5UdCp2AVrnB+qZL+FelqTZ9gZyewBgDUOOpC1vnNqk33AEgl0miDZ+772ESp4eo2
O2rt2hyL1+h2ajPUsYmKMjbVR0PlbPYhT/EAkzUalKwhZBTjLrbIltXHE9iQd1oz
lHp1BTZJSx7x14zZ6EGYNrFQzVjYLexluJNtpPhRU7BSJp3skoS5whiJXWEgCaaz
DwoUc0blIeuWKcwecYEsKjWrucAk949VzKj4EYvLdarwfhFTutxjyLIEIAHyQEjP
ZYSz16KBrb7ZzXGL35khKFVljwG5+7iiit2WGpMwDsUoccQ7AEUS3E5MDVKWyv55
Ap7iB8sOdG8Z+GABZ0dxiBO4amaVYJkAPMAbjhqbR+29Iw5Jxnv6o3VlgJgpUrzC
NklHedqyk3B2igSwMcGZeq0tNLnkKgcCn0bprE/behX/wgTxWxxkt5npR1+Wihl3
GV/hQhPk81DXmyGd/64TYpYlrqEU0jVl1qzew7LJcawmG1xA+gHwBskSdihxUqAe
Xd9CFy/ZLWeMF6fro55tKPro0UthZzwcnDAQthW490q7YlBP21eYNvcRQwEI69bb
KndVvRyrVIyRUQ+Rle7vQBEodIpefvArU/Uj6pjrKVRrF27k32LGSyUZT5hrRJSI
UQ+QyG3o4uJfslH3sqTk/f5HbBaxDVYLQ2R4w9HZiY6ET+BHzRgSfNNcbY/Jn/PD
0c2/4Kc09MT0Cfb2/uoGcf4RWGJXZ0QSNp6/a/eqrDZMju+6La0LUkRpMsI7MJ00
GznzPG9l6pMiONtkhClmBn04FZZ7rY5KdeaGpX3NPXntnO5cq63mTydn9rTRNUmC
PTWwYFxubAqjQLNOwIh95/MNFACWLTH0gE38E34JxbapblCRi+LRW/pVBMPuAUWs
u0i5T9yDLRUuDcr5ADYAM8T8v/7uHxtnBr7UCUrmTnlx4xGVIC41Li9JPWieoMYT
Ux7gHwLcR3uiR5UIAgVCZJzWqn6Mx8WBevVfQDEA6DmTicaXpL7ftircVi+r86d3
GjfwB5WWwKodzWh91qYQ2QNuAZMMbBxkaAr9E9C+/RoswrdpjWGTqpAwV6Aj9CvM
4Emu33xdp1kfqTroHBroTVYDUfqspNyiOpZQCQ1cRPHgtJ9+GsXz/DuDyD/L6R3G
3A59LrmShZvrtWKWMy78MuGFi/gMHdesQiMtUuF0mjbkG9B90hp1tZ1qJZ0SUV22
ApFsmwcJKZ9r8XSXN1HFf4hfxwBWVWEipsPqgqfp86spKtU9RwkyKac5cDO9brOJ
sUL/wcia0G273AzpwmoJT3k1LCsvGbJEGzhXPjV+6ml21U6kC9j3vXhy1P6tWBhJ
HSO1p3QPom8ESch4VyIxVZ4G0chhETv3+er4x2D5SE36kReYH7kuERe4pb68iPbl
KgUH8HCPdcIi+9+IM3vOVilEK2Xe713e7SyQW0XxNDv04lGBz02YNr9Q1bkA+CMK
XOmUTeCSrFPSKIJpHtEQLdlGirqhOCBVRDug5dCKwyiGgtTS3QdMWgd2kvTTMpRv
sj8/1Aq6ErbdKL0tZv/41GJEA+h5MRkc1iszzwm56BactLdse3iMb1eK7IYqjuJq
Umh3KKifZExwlE0eu3HcE5DkG24clL29IVrxl/11i4MAF1SkVbN0PAXeOofWb6mv
YAhvDvcxX7n+NHsqI6RO/IsgL8sjUuwPXisj/oXIVKfhlpAUbux3NztkUCEFnSSG
CFbDAwhGYhGbWaVLKxjdNJtfP7iixw9OqFYJ1lTeTss/H8ucEq8+DV7Eb5awIJzH
iq23UHqcykRVlcnK9z423AXSkvY4gJ+Yo8iT9mWwDe/Z8ziIu0+Bu9oM78kbKTYH
9CK5AkdRGRQlu8cJjQ+0oc9lvx/Ca1Oc8iul+Nw39cGG4vD9gOmS+1OxcN7eOsfR
QhsYqErJk2TuYAuq/wxcjpIESPQ1Dnf6WZhxC2/p8QFu+6jjidjoiczRdwDi3YId
hndv6UosESahrTaUR+nMQMOHxkUvyi08sX3P9UTvYvdjeI1Z/gPst3x4Cv7QSgVM
8kB20OFUv9IOK6iIj/UfTArjvMsgXakjyJWAL/eC2wxF19ssRk9crVHyHpfbUxmp
fBBPVWv6y2/l7OL4gCI9fqakDjnR1VrfS1O1cMiqkxFXC8x5MTwJ7jgVToZwVJHW
jK2Xwl4CaCdzw+EP1B3Bkd9xe08NbUJwgxmhkYzwLxRVSJICvPPdsbj/i2dRJRCT
mYgFQAqDtHQFywxWg6UpUhtpKs1+TgaMmH4Uq/vyFvrLw+wtt2kiHRZi402qe6ns
d31Gi/g3DpAkUJlEGAGPSbbZXsdWk2/DC3Lt1mveh0+IyJAL21WlBi4RHoVYVQ/l
0/ISOpPJuU9ASQM+BEemRUKseFt2V2LdZRz4xy8PxDZ40ZVgTEoQstoU48Okh8aZ
lNx/qjksODNXnpmbqUyMEoJOdCjeAtgaPfjkQE02HBhhP51gaTbIZLUIQOj6C/mr
1x19O8HDuu+g9Q3SjBtpxjbDAmTEXq15SgeAYJCY2QNlsfmUmICoYT8uHgBBbhuA
rWZcKwGv45hnl5Gr0nk1UObNjdWrxpDeUkoJto+4u7+i35O6W+KiL+NGUiq6KSwE
fzzu6368uAtYCOK71c7Zs+ywMw4Ksx3Xz9rIh1fScNLChneJx41TXqmX1/s0hTBO
Kul5B/g+S1VlHER6Z69pulOqv/CYtG6HA3I+iw1qJlYstDifhZzXVX0hcSHHROxt
8aDW8nivuAYZ1E6n5gqnDF3asCL/ykA6NJY8EF29uwmdNUi9N52fB87er1OCCDY1
UiBu09hMt69QQLPbn6LXi1Yp0Y+6PyxwVo2CnivxQmWIubgHxcaHO/1mFRZEMxLZ
0Tcjl0x5MdiJ2ZRME+c5k76ZEywhIZtr5tyHg+GGFz9HN7JGPNyEFBoe1dNFArHP
LtHqIVAe9rpcDf8opfv5bR5EfrDYDM6K9cHvSjIMfBSZ+hUaL81uSG0J5m3rzy92
51pTmRy20Vg2dUBWv5uQmXVafkSXR3RMBeVCtEBV/Sq3bxnHz83kLL1NS0sMxusW
+fHVE88sRPZU5LVzsSrmAtg4VcmyaUMp6xiCZgOkMf3aVuK5xZX01Q2B0knBgCLG
UIpDRQTmHChAgNZkUxLkLmhoFe3pxoj0HobpfY4za2algi/DHDyfgEwBP07TUaTn
1KopPaVfAaFIqgTcxlmKamydJFmTZAdASaHQTwzRX8O4fI7Ek1XF6p16w8/IZAfz
XrJy99lxmj185G5dnofYmTCnR1MK5XBq743QRFcte4jMFyvGGDZe5GQLRzlF1/IC
0f+Fps7HWg5t4fatiZTlF3jOQUWmccRV7S88Qe+yLbKxeAWMbZWXW5ef4WeAZGms
whnaf3wrvUGP/4W2q7/o/XcnRkpGOewrhmFXoHAKfuzqsHQ3NGPJl7O+I4AXbKim
rgMVi5i/dKWkrsBVj2aRVOKHK9I2qgK7lKIQICQgRmNxleT/hVlmOHgG4HyXSo2r
xPaSmc6eEvub0EnbrXeC8+bDv9fvpw7jLYfiuW2Yd1yskC4I6n923wPDu2zoNfvH
p4l/thqK6hqlCLtRsIBM6jciEIERA0sQGRLiPGif7tRPs7vold9BroJ42UKtTjq2
M/YXW7fMiK6h66Mjg72we20FMABRYPrGQLh+1AcnPY/M2EXOfWCDThv+8RXW1/ti
U2nE3RoQ5e3qVRAcYY2hlQIcM/jHmoPdiMR6MRa+InKmPct062oMiHJnX6PBBMj9
mZoj32U7TYRBRFO/Q1cSr5dCbLY8jcfDFtSJPl0G5Wi+SgoFHolzv2Xp5aW+8Dhn
hYSvYTGYchy8Ii4nFlPMmW+YhMJJDCGlg10AaUNfRNXC3oWolkwFiHYF4AwykNun
2MyWDhf1/fZaxSaXnAYoRKSoiBTYLYp89NHJTT0jSNLMj9Alh3IYcMUMZvUYV3AL
IVCyadnKDfaSlfvQBHZJQyGOr6hCgGakLbNuw3syNMIUNJ7FWO9C8RzswJffpMXO
HJuZzzzu+vrBIil3Z3uYPGYRPuy8/zqWyJsXswxDHRFKRdNLFjuvBHbbPt/HCgxj
sI/zy0dHRKHtJz6ZDw2lfqoxTfj5KBYboOtGrOSmikaNmfUaG9l8Q9YD5uGTiM2w
dLjAgvs1TkwqCmwQrTAJ33+Csehp1UfXGN5ACNUwPtRSpMu+nENCyKxMwQnXPyXN
8z9gn2zwmLWu7Yx1MozO8tNRO+vohw1TCNDe/RW94Qcm/o2BfzNEgI0GstiwRybH
crjd2IVSRUmkS1LezUZA7JUSjSU8xlbu5D3StWbC2R+QU0wGJxGbZMGk6dyvCQ3Q
RVeJ435jHFY8qKFZ5F+GCsc3CyQtElNMnCyfGEyq6Q4H/hzwTtvrxetaYcfPzQ+T
ejVDsvLUvP3XVM0+XRUJuuOw6EcfzcQDd715hZOOx1cnpVfgp0rbl3MLSFOH4nEM
ldPLGnJZ1Elih975nFGHuFp0KhnMIVl0/TYqiU2PP9WmC4ZgmuDYI+23v4XpjfPp
8EiK1c+j75SH91tWbuwD+o8ytPx/kTKpuJpjNJ2Qssl4yaIbZyIRwNwK0EB8jiJw
LczoFq/o55cKPl7/YVYNG9adpcw3UKTC8bGTR9ZjYMdOkg29kpRN+S8BWCm9xaeC
+2N/N0BLZr6Mlzp2wVEcGuylkCIcWLGbKlRJdz7+uI+aw/cHO3+sHThGD35WN9LX
NbBYiHcr7GJDF232TfNJ+tRdFq9RczcgTkr0yHRFYVS8BC/H3AlFbGalahecH/LZ
LEUxYqD/IT70HJlzvyYBQRZQUGhufB+c5VJX/7tGMZYNW10sCHDX+HKXmia+W88A
/BWPPmo2oTxy1EONMbrqpL3RDJEOskpqnWjQtxxUGyB6Cuu+JF65LjwjDCVWu79P
XR1oSrso7P8MD7cZU8maDhub3wtW1pNEPyLZxq4Wp62rHxkNFBne9cTPurPCskBv
0qN2AB+DcI7ZCeh/+FnJFJYmKqzmVXrWmh40GYcnOyqLoT6Po52vDsC6aulkpVE0
O0rlX9A/Gp1JLhR1wX/8wXvfVeRnmmcFio7FBagRyY9wWG0AqcJK/PJYSjbtd4Ol
5K/e0IHJmS7PPzoicP4GOwqAXrGo4mgR+nhnPf1DcUrOywbhDBWKS3mgh1mBoyom
zWLIIQ5PGZ1VhiVMUAhARbydnk9MSMHsjNfzNhf9/kYug66pQaBQN9t1YWm6at3n
+hQUi2JmG6FTfR29fE6eOZDx4SwoXEpTL9KbwTloSRZJMrQkdcIvMHN6y2aylm+c
AlaaMsGDIvury2zXLFVL/kYnKus5SNIl6iAo5QTrcYONs0F9vp5/viRkZpcjcxka
Yn3HV2il6BeV3mZYJUQxfLyRlNemMa8krd9UI4Gtc368ebzYGzgWIv/+DldUEVZR
ko96una0JOp7yTty15tMt6AZqs5v+VcAkEiEp8llWqt55rjCl1pL91gjHx2zp96I
ijp22Mw0pZDU4uV9G1ChO5CwQJ+CY/r42Dh32wBmmSHFOzG8BnDAoDvL6QBktYWe
59iJ4M5g5CGb3RLkSF+0qIgv4fUzL0L+694YXCsvHtWR/9kG0cPWg5u3m2be7jNE
QokOZsVBGdCRWZfyzKI/wm4Yu5RSfwPnwMRBwqGOAmaY7WAAuF68opsX9f5j59kd
rHJUerSWbuvLHKQbNMQoHUIvnsAY6CAbe2R8DKUEjxV+8xmtrELUI8k3PUD9VKpx
Sz10mPLsj1YkQN/XqNffkFjXo2hh9LU0zxRVe8qfLFYNtvfEKa9pW7FoL/mrDyQQ
GQXjdFJqisEQse0DjgU6LGG4IragtMu/AylMK6qv+2AuHbScaxzKRu9zbFaMZKT/
ReNF9koKA3gs+d44D8A2I5NZrTrb1RE0JAUGwBOv8Hc94pNwXgtXsBOkzJnJZoL/
oqH+PxSiA1gNkheMcq218vTfulxUULo4DWWV03aRRt68fV/SPehi+7OT9qY/VG39
TFcUCrU7KgEnYxIIZ6+Vx75cbyX7R51zs1YeyKdlSs7Zt0R0RPDQjc29CMSkx7ad
Xl16SYA3T2iRjz7981Ooy5aDatQvbIWXIvJfnUkK20MV9PzDwuPAsgKcv5eguHMa
e0j3RMJGcwZ4B1Xbp8TtUDiG7puEIICewprgUjdKQumWi2hZRBRphp+EJ7kwLdZj
0nhUZACfPXXZWoX2/pQft1dmFpvhBfUkg/hsgOGXiJZ3HAAlGqQ5U667sI1r+8cn
go6S2mwNFDcdKw2aV1K2wuy3JPRcqQPSkOVAxmlRnEx91XQfdz5MegyuF7/Q1NpW
TZxYDsFFlwlxAnDJuhH9b0WX6H3GIVs/X6YrkR3cD35xvwP45b5VcjlHy9F4RGxI
xp7yhuOjvi7o9KFupnm+kW2tZcZZ/6S4pgYPtOiLinqeUTp/SvJOQZG/PK69usez
KGrnbMkM4CCoCrH/KUDh6MJ79FrrkoH7Hpo9pjuJdG+FepEW3WUW/IBbc9X9BWD5
4lPwTZIbp6GVbMezd/1cRCkV59GM/VVA0Fn9d8tKdSvtYxzUyXkKgl2HO+uyi74o
wnf+ndSycMwMZuwiMQ86TBTSUvyHkGq8DqvOHAN+gYwaetDqSZcIAVfbFeHMOben
DuAtoGU5XZAy72aKOMNYy2FEcSY/kQN9+70jSGkEEecB0WZ2xR+rpswUq8kB8izX
XtuTZxZqSQ3LjzmV+WufTe78ZNl9bb52xvLuT9VoTl0Fm9ne6qemV2EozDw4VDT0
nNpi0PrRCwoZMEtcRj2t5kFRTHFtuTCI6Qpuz+7QtfgsHIIuHgJOX8box392nw4t
Vo2u/kWJyyLScwZ0HPdsKN45Knwjy1jb54C1oyDYN3B11/tMcj2O6x3LQpDDf08X
fJLRmVco+4wFfG9Lrg6dUVzTVSh1QfkUr9rKW+11iLvX0f+z+qH3MBu/sgavgOKF
ZefB9BQk1g8/+VR6PTpa3Du0UmcSeSxIIc2j2LCrWkukZ9lagzSlZgHuVMOZPomR
LBmL5X2SIX/H13QiVRVORNSJ2JxDPZyhtjPXQWsegkpzOszHO9asuZyqK4h/Qj3s
lFp5/RXJ3XFGaJZ+mv9YmjYAP5W8iXqN7sSgyWCI56RNbH5pc0S6I72kIPRdSLC2
aVsxoig7U8OeZ0hKfAaI4gXeLYllWYbyFFTKhiVrDiiwcRSvQ1tqQtNNiEi5Imk1
OFgZw1O5xDXmepXqKkGOyEMYOPLSXqRVPoeduc4uro2fOuFVJjQsI+XNJvmtgc29
HOdjg4PVQVvZPq1syxVCUY54reW4CFoDl8HuHPJZGTlmk2aaRrelFLJW91eBTTze
yAP6rPpBRNmMpKdfZZCid0OEdo+WogbD0DcH3FjYuoIeaqPa3em9XnLRpVhYw6um
nWlS7Ne9+Rae0JHx9Nwy4pZQyeHboRxlr+FPfMQZlNppPqMWsj4G1iAgpRnbMcKt
k0kCZajX3Y0pLFKNRGfjnFUFU5w9BS/Mp1dGnH5MsI5PyPA6u7yYpti5LG7RCZXn
LwHCW1VHOUhu+SmXxEtXD7gHH9RYcjA+BUlHl/3ELWOGsPdkMh2lC3Bsac4+ijA3
vhQaetKqf7hfZaEE9PP8OI1NDqU3gDwIrbGO/Eka7moC2JdEVwR3FTj0sTKXjsix
CCT+c390QBa0wtJoH5eSWRwC+HU8r8HiKjGbidGOOpiNPrCgXM2C1Q7HRXC6JV+g
PLSHw9f9uHPmRjRT2dwq9171sEV1Bb5B1n1Ulojvyr/JPhDyLOVfWxKGQb3veXMb
2RpCrfIx0kOQGLY9BId/BQq8Zyd8gY164GMhpOSMTXORvKne+lgHcCo4xdqBjVDJ
q4ESxH7OEy/uHoxYDtUaRaqlZSpCVuWesgv3Tot8IY8tH0RP6d/INoSCABhtOtZl
CWuhEPbjebT5ML/eZr4orHOiIfsr+VaZMgXH56b/8TRqXUlIsau/Pn+ACUuilq4x
UsmdVa7R1bxTYywlcHRMGjX5Qk3pepDJYXt7y+iS8DW2OpGKH22mVrivdKSe6GGf
Izae8YC+Q93QDpk5yH39ULkOWrmGxZmPbc+Fs1yyzjdwP+AhPC2QtGpkxM3gUDvu
7c0M9zfLkmrUJWs1Od5QVYL1NXXC8g4SwiBxQAg/gWTchTJHbPtpBALLX/m7wxi4
VEOKoZ8mgwhyTZyjT5scMVlGGXJ7IM5185/Nt3uSwigxMdIAKsmrTIApfEe+IVyr
DgwOMhDOlNaEv/lGc1K/fFOvTofk9mpQycSJ3qqY9CCF3NaZzGIDTkLpbdknnSw0
hyLu+NzvKrqn4NbtK0/WGnpOToTIzL7RMJUTUeMS8jtNIk9O5RDVz5ljF0H18H3I
Samp2CSuiVSercatwFJXbaSmsIp1QA7ry4d2mKEtI/Ytd5QdTfB0tXaXlE8oP54x
MXXypWtxujlJquDPFmrup6eAVI5pFYSkNRSi2470MPB0HYPesp8UQ6s3X+C+tPxb
DjtR3eNiW0su1PtX8xGuLmNHVXyyO4xE+QS6LwbpVlyDlUu+eWq8Th1JnuAmGzfs
AXV5NIbP9nVpwAFVOwQ8w/egsGujbuuU5RNKxaj32UYqol+DlJd8b0ImEs/ic1Oo
Ac24YGtfdKr7J/TQV9QFFg/G1h5fqD/Ji3RaucsgfTJqvx/1TsCwI/UUo2nRsZB5
WXiuluH/3a3h7QiAdAFYJVDmRlV4RO8iq/YJWUMkZtsJ7iC5qlTbr6lscXDTHrmu
rrWGIuLYBd+QPiwk9KMsaVKjDgAUzDcSLHldLOoFt51p9ddFEM5jPDPt+N3AicXr
jY5+sv2xWRqFO95cRXQzTzyOiUiWMnAJETcr8MMdHfRwjh+9/ccaF/yYmD85uCWe
yFHMcEUGuYI5hY6rdMp8aQxb14PQGzm0nPss8n96ikWKB9hsxxsROf0b5JUbvef9
Pprw8S5aDhckl4uXjlhYI4E9gcF2MzIR556f2Cq0u0dmn/Dlenf0qT06h336DFBk
6jpPJebxSe/EAIlAiTdl4UgYCWz7AhHzk/JlZpE+IxC0Cb2jq4Upe9KapU94cNDc
RZGtRSO80FUUqi4BQWDZNGZvAPI2V2y/9WgPzAkcmYIH8yGs8OAwBJsh3E/qURk1
AT86KoTtK4/PgMhMW6Sr+3Jj32iR3PodefG4/lwnP3zge9KcJk5xKSIoTRi6nQVB
+aL741TXvou02DmX8mOotSxmNMGjMbh/t25mbSFV/HM+dYCmoGmVPOb+eQx/f17j
OmblwT+KUKREz97WS6K0JSmQiS/8GMy/5F3JO/E4It6HLEznhsd+27Nm1N1RWQqg
pTY6UmkYuJywLET4MRPZ5QEIRKNKmRRTe7/qv9CYgfg3BbYXtVrzCDNpuY1jxhEI
/Ld0/KZYQnUALK2YdhkQKyGVUr8vXEA7IUp5M2H6u/mr8qlXvvkXXrVg95PA4KiU
XTD6VCWjdHk1q49RTSZnDmGWvoLY8oQbCuyMVySo6T88etfVgSqDWwsHoSfAVbUi
mKsjfqC21OFNqePVki/pANoIJgi2iLCyqoW7MQdr8TQ8Ch825hLsUurI6Ap7Q5G/
5a63/RvZwNNLGYdKAahA23P8Z2T4/pyP4kU+RJuJ9/jx+ul9nSwRsRGFQW/lGeKv
RavenPF7hI7EklKHa0S1JXk7FY6NBlV211wWaCTq0VBXKIord5UQZ72+d2r72HjT
9PGXkLmHFuG0ScwE47KKOQ5gHDe6h8dH/xzgLrTv4xv8ezSRimlph9t+Aa+TefKm
flWzT8SpBJzhI2GTN392AMl8RlH+t4NJezrSv7vbzmCJARbPZu33T26GuGj1prdC
HMnQWhhHICk+eiU0YPxiMDBGfwEDAYBz88MgX9uox4katIa5rXouycL0wZ6T9s5R
bJU2RdFThsFHZAW7RliMb1R2jKVUy4B0T4Jc87koViTD3MMwhEabWlh5Q9bRNJk6
58PHbZocad/hUa/v0Qthap8QYT2SQXKqHtxmTkZboiZuaJRFozotIj9T6gVPkZmm
zMdRUSQ8NAGuObH0EEL+JiPrmcaBo7bSu9l8GOTa5tocoC2CnM2KAHAL98sR5XOt
3d+tyKmQjlKiqBwE1i4uGGNfyEFY8Sm5Zh4LKYnTLQNiAmE7KBOvxFUKI7M5yIO/
iEelOR/iUxJurI3D9piu1rTUDP2HMFzx/m3x+4T0UUXV/3rkRHUp7HVeolkYIurX
Y2QDIh9CdrKwYzzZrHDKNwcsMNNxzCCqCmduRvfGv74CbmLABRTPuzVyxZCwVw8X
9wV9YJimXWyyAXMmP/EFrUQRVk5X4TIXp5muiIi3zE6q2p3FzwGDWslI0EgHpW87
66p/yHApBq+50gD0XaJlyxifyyOeVeaPPU2GzGlpziisPSULYaRnzoXNw3AO4KWc
VIOWYpeLGXFYYzKh1lIYcfUdnduCfZm+WHd4rpw/rDtBTVqBGJNhzOke+d/LfzZ6
txqcn3X5OMbGZ4ae/rEzb0lxoHP5jF/aBSltVIlTtlE1nDVOXHCxEjCuRyTfFfQR
3db6necEXw2vEjyRSkSEMbKWTR/K49hxXeFiqhhuFQ52v2Cxw0R76RuWb+79lewX
9TLZd3vb7fTcO1oohbNDWJbwTXFNBKLdZUw4eT9ov7juc3KTT50EpC7c7sC+LRqW
qkdZCJxAyzY6npqjRxZ5Zie1E0S/QMav0tZlMzm22QMc+eFJYslBi6CFihIFG1AX
2kMnh4uG+wkYOkxi1WJ6wW5es+qHvU5Qkno4sT2LtXnYiGC5LCKUu4gaHW+9OnGU
nzedTiLLrCE/JP77zEYq6kZxsWyOKa/Ngivt2xRYMtYIqdmk647I/R4PCPCg4ssl
n6NxKPisIrZDRG0JGqdzJcAYEyDeixuwNGuB7s76kExUu3XSJm1sl7OVHNt4AMMe
BS4vzURQ4Jlyldll4v4CXusaNBEaj5vsW3a0yOWaEVoF1o8hL+P2lMPWsmkCu018
U2id2eq9Wah1/LeR4Ca/efb3/PE46loDvvaMAZ1JaGP0cuNMLvUcJoWTIK0UAjlN
ya/gnI9A0mQ+p3O71HFyKYxZlEtYUcH7Dd0gey0rEWMS6DxOpCRP1H0nAytHm7il
W8iMfkeWKlPPOHJZVp2UqWqx7Ile4IqnGpSZgxjf/URRuY4EbzwYvmxFvERN2IEW
Zz78Ds3UgZbrqI5I56lyg2r7b3oj5nGwj2M7+F6qe8xDP3KKQHIvZ57eEaIzwEA1
RHdwAVxGDcvyEs3t7X2gxtgDgbZVxIa4TAOytY1q2I0BzvX45xtniCcnZvygtSEg
oTP8uzsYxyoHCLogYSPA8vTkffjAR29G+pqQEDO4LHI4utb6fhaE29+v85Hiu6ii
miBBFdrIOmWxwcOcKrlRovznIw5qOP9SMA589a+HmK3w6lrbKtyMYOMUNMuX++zW
0SdimLOFGIRNRhM3/4xS7Bux3eA92qphYdMi/bdNIMWos+ioSHGDnmM1FFARbS7X
5h0do7OALMwjkwOoBdQkj8APE7u1ca2ikCgCC4fbibfIk2601lie/THxB/cKHzsl
euRijDbAJKEmaJkjYFmMOUuieH/gv05W4jzusc47y5dzSSMJ6NXxr4gfwvbZiXRd
Twu72M3dfr/0oxGW0Wit7ekXQMEd4bHS55RsuNKtnT+L7hpGMmvfkNUt5tPom9ui
Oh3HU5Me4/xmLQmiMHePISrfCBgIIFrMrfwaS5XPNbohkIE96I11b/rRlJEm2Ao1
a2fgoxGepRg5auhJ9SCmtPlyEFA7gMbmCLwvyLfK0KoffbdxkCng80GfYhOVgCDI
Rvg6rlhEMhg6eN5f1O4rVNQjQ/6iUZBVhAfRzhFF1+tb1S9p57ao030vrDAzoYx5
zjw4bvObDDgDxaiBNy5XbKzzYxIH5ukxwAz+hTllBtdc7iAWfJW2sbHVaojQmDSB
J1Munct5teGoIcMHQsoJJANJ9b2Mu321fdxN9+fU8Au9S63N/AvRW0iqf5fNUjxt
5JAGd7aCknfeUxvLjGTaV2zJVLpA8paTlTrg6ST7FV9LM79Lae09SE4udyncg21i
bAqABbfuHB3s+/DWZ0u4+jbwl5bGYccbhs0Sqrp1LnX8AdR8wgVCSOMNf0d1utn+
I2Vvjb4QRpyBNU4pxe4TFKlmo4vnsqijtmUMv2/xI1j62GYaHFUxEDK9LY5gyptQ
BawL9lR731BIZ5dnNv8L0Vb05yxfDcTB5roTuYDhgqDA+vrp3CmuWd1rkecbETUk
DWJn7rPDKLKGbUNwFgp2DExFnMrbeF3Uluil4j0EnEZ9YjPye3zWQe8sk+0DLNEg
Bp1zz/hGPuli8R72oDMwL57xLklnOJocaaHd5n9cVlLuDWUKt2fv2gyjK16RxJKz
Dbs9O+3l02UEkLXeidRMITUYwKY4lNixcQSJ+2M5C5ToxPdhF4sG4ZoZiefjnJCr
LJWdU7lMcoIrde6jkHX9lpYVUyFhiwRhLomaR8fV4q+xZcbHJXoDBRigNJjJG3m5
uhfxydP0TNYJXBRNfKysbBDS355B/OlY+XtZVGANtfQes9lgiB74cwndlgr5AmAe
iO6sSmhvVB3X4ldm0C849vrcJ6xIqhN+xU6R3BYNZXwcyV1Fsn7VGeShvNN0/9jn
8XywQnMjvjRAPfIxy+AlgFJVUnJFuUm2guNrHCcRTIrD2SC9xQ9MKcwnjTE62t1S
TReQ8ez5EUxp342x42doCk0w6bXuIFyoGp9G5fj23xVNXa3ElOkByyyys1RJTsLI
UKUWiOZGv5p18x2H/i0W+h7cyna3zL08HL81UZBd+8n8udZ9jj5UXw4R9Tpo/JJ+
Q5pA6CdFy5oIE/2+TsX7SfSp8XYJ3vUx3u5YUoB0XcOYpTinPmrUPi5NlWmt/6jV
Omm8A0FbhVOHSbEr6FvSQWEbLjpGdPjWPQOFEkqd+J7IH0K7+TUvbZjhs61n+G7v
/6n8ryDJ6uvTTotL5cZpPB0HoASs4UpvsLBsNffDRam0T1+PANRSFD/yYG/o6uqJ
nDruHAjIOpatCG6gmfcolrn9mYKVrpRLv225pLmDRKpqNoomkYkNAWjJvg+PH8I4
pBuAnWhuLka+Do29x3VHHPHrFbXeaRgVKiz5FwiKNJZpB31ullxWHEE8PRyxWdm6
3B4oJtiEI1nVcTM3JOjSD9fCU0PpRtZ4SkT58KqRUk1TTnijvi1fUOEhM0HcBxmJ
TTe+a+zseqk3HzS1TRlHFsac/mQ+xdIZm8HHnYGr9IAmZ2j5vUwzg4eeR92lNzL8
IeURrCSF6mJxAFiE+el3I4UKb+iaLWpTlPh08whpTX0ep3PdM5rLkNQIA5vaHnz5
1tYeeNXKnIvy5JMFBjk77P5LflAfv90IXzd1o7fwn1zS+64d9Zw4gYsxw6xI6L53
fkd3j6tnfdqS8tlKN9+MbW8E3+qWnvHTTIZFOes/f7Ys78jAkSOYbYDtOWezcUZJ
BeyLbg04bZLVjBmKLdvouoIR3KAZ8DpSweSXWUnG9w9YX0+ZKXz9XTjiUqJMlYOh
6YRbz8m5bmXrpGIoaWQm3kCeRZJrzuGfwlKQgdO+aQls9F/kZClcfZ2iw5fiui9d
+vMHo7S9hm8axuvj7vKgOOm7qUSavhpSJT7ySqW3WcIw2oaLKf2TxUse1o1EMIrW
jfYM92Y8pd7UIvBolNby1OkCnbY1V2+SluUUljusIKP5WTxPScgRavxKo85lvhVy
MK6663PWvQafpJnGprW+r36nYGWiLej+JH8ZOqo2I/oszR1QZZntcoVOMcoQGTAQ
7fDSrWjdFNt3ItH+ORZRbtnPh115yO0Wac24tFd0wMXbn5VSivDjP9PNI1TuMqSm
ZjipGu1O06ASn+zPDOMDoqTmlK6z+nU+Mg560n/AvZ6GvBNckuFMwVK1/0V/xn87
zXH0YbVndAkPfahHL0qcy30bzoG8WUIxRnXVAFVXG0uwgKHVwdHiKiP9b7oCfmuX
Dc8UbDFyfQqOXA7kEr9JN/L9AdIsgCxppJNBFB8L4hI5uyDt5upLX9NzE/Fsn5pW
/Qn5NilY2fyp6aDq+lNvZKdTRLTe18Ne8e4ueVGa5utwfWM4MTS/65W6UDGsUZcp
IYnDa95bhXP83rrYqT1gWOy5bSzIpP+8Obq2+WzpSDXR/BezsTi8L6tgG98bt0Qw
VzR7L3PLG6lbIp6KiyNZWqXqOvvDXCHBLg64+P/npjG0TxEj9nY3hB0fp5GHnto6
oERj9n+DFp0EKZAEo9GdoxwP0D97lJl7F49kVohQU+DpdJfixpW08KwNnzn7bHQM
17CYeZ9JAXgq9oFloooexJ9U8vVDf7TrwO4qCIv4faFZkSG6T/GAD7QoxclV5c4Z
Bpe+w5qNYO87MMCqNfPBZ2VK+q26ldfb3I4PEsh7RdrrE1g5yVQ+6Oi+DX1GxbrY
WHCKLjjX5ODcfq4IXvTg4DUwpDrTWcBEYZZz6MdnqIL8VyuzR/KZG8Rhr7BiZfyh
YAYjel/WHhwROscpQ1VRgLrcsF3H8WGLzLKFrVprnS2fcmJAtTEw9azczpzMzD8e
c7t+c9uQRJSXGArxB5p7uXj/TCdX93QkDfTKhCTw0OgKwQddKRE8BO1vaHAqapVl
tSebJSo3LoPKYaGn5fGEZGOxkyLF3TG1bJ+LWVnS2kvIv93XVnjiZBWRpTtUFgVX
VKaRwHd7uA8IWyGhiT/vdluTRWCOfQjfztIxEiKXZFhO0Hd68riKrPx2QRX/ebUp
dfqrSmKkDL9RD/zt5ynCgdK/CFe0v/kKK1364+FVik25bIZJIHqVP3gw7tKZ9O0I
qyIk+daRbfj/MYqb8FFGkY4vHSzP7P8CLCzFOCN/xwFq0WccWfWVgyu9tAE566dd
L7UzKSP18l6NM9Ja1JvcNVnFuirXLs3gqYdUaPUaRT+JvoZgBg01Z7hKtk07+3Kn
n2xCgiy6MGoq/2xmVf5rLwBvheGy+IhVEqxuRitFOT/LNqpp+9M3bxaKWSONBXNY
SKaPV8haQvo37/V6JgD7gzzJvSNza0TDfG2ESEZrCxHwIeZ/7ujhPYZNifh1DN8K
GEYh8b0v9/rtJd5chOzlFVyzva16zsSUyMHTsSGFGBeYPofCqsMFDwrbWXSXy0I/
OnwsI/kM7mJBHRL9DRUdqkbGilkryJ5MZhlqutyjFzqeXr/aA6GweX+4J+4cts9r
jzdgu/1OnjvfrE+HzjiiR8KUZX+xCZqpf6gAqy9Vr0Oa3MBsW4dNV/HOG0pU1cFj
srkjnWHY5V2z2mhCpxGMCXLnD3wW7LoOx3htz2Ww9Aqc7VmoVeAY6tZLPwcpmACN
6e5kF+ftKSdVZh/OcNvYAg/XGMraB3o2Ia8iEiOrY6/ofoshjoBIz/ARfExocNa9
s4Y13fMnRycjnMci69bnzjgVIVZMlg3TOf6o9+VXOU14Vf8yHLu/TssJzNw7irs+
siYR04Qx/wj7T6DP40Rpe9LF/paaePo3W3QYk3itWEpjleVdS8KrogcHx9jTqHTo
5YySzAeUdZMwWiKxRs7DgSt4gKNdNtrseCj/khQR+RfKoa27VdgFU/u6Dn1p93+y
31xkmbDKVx0xpAmNzVg7Y5fI9Gn8WCBU5JDP1bvnaYd8VqlLG2JkRQ8aJZSZcQck
fIFFRBqhdueQi4My61H5Jp+taKNsh3CLeAHIr6cr5yDXXQX9g4txqUzROvZToamj
qriIEA25gANQ9RXfTe35P5zEqls2jEY7syncnM0p+bgZ2LvNOkxPc4IDkA68t6w9
17VOAd6zXBwNqpmfxm8u4058FbyFklkTR36lC5ammKZ67NUfK7CpWS+ngMruQsum
7K44GrlPr3BIlL0lLIaAGye7KoEgOqfoSMvliB70UjWd7k8Ot8Q2XOK3PWmE/v9M
Ub1bXhAFBF1BRNTQD8znTj1Gt/9CzxvwBGGsTXQEc6OUtyW5oUgqpF7KejysRJiE
v9hv1RYHJXuRuGDiM1LAxrmc4TnctZE+OKW5HJbklJGzqR0JD3+H9qdw2dArwMTf
kuruzljl/4azwWt03m/ei35732zFzFokHQMneqcjeAo7imeZhWUAPTtlBFkrrRcu
exF2TjKuncqd7eXtT8I2b71YRe3Zkao5hE5ce6ZJJcjhvzHFHI1v8I1yWfJHrErW
BjqodehdVUk6LAfTp3zmwhAEtNHUx9bb4wwbY7S2s56mMaiVKqVbur26UTJhQFGJ
mFl5tyRPZnczwr7vEa58pFqqPDBPh8uSVbfY75W4kyItNs/+tuSTDH/jk+m+0XaP
E4D7eNB6Eht6qI2laonAhLhJneInWuzHeJSWK66BdALAdqR1HTb6q91Rxcdm7Jne
Ne3ygfMxNdApBJTkXIAoSQ6uQhhqG6S4l9aegmMMlvsf/I9XhUeHpC7+PppgLxlW
iMPrQjAWCpei54sMbYHXYfrOmMqHUZIfE3uYpaz/KWcC0BB3HHBIrDxDryb5n0rA
No19zYq6wTT9AmbXbWIl0zYc1pd/iFn0QBwIAIrai+LNPiV5GE8a2bZgfPtbSfTN
5ImtMbjkHSMlvqrKIErVq16mvx5NaTpcdUZnulHz0fWzyfXLOPaZpRVTkt45urIs
I9auDu6VvNTfC8CUNjlakQZYcggvD6ws5v5nWkQocwMEX2Y66Lmwb4MAXKlXdAc+
uEiNPQlGvmOZJg2YWfgHiJ1wF0hg7luq1tPbzOFmi/cRD0qM5J5kKn3+2dfUvzLT
dAIK8LGy2CtD/LzwfoyljPFcSeu+n5Ow0NgPK/msP6Hz9YUr81t+QRjG6j+vN+Tr
vJMjJdOdIBdKiqrGL0FxtYapuXqqNgnZV2ewFo4KIWS8PObQJ3CQOZ5R/kaktzVA
sFu5ConphWKKqSiYap9bM0246PcSrGwND8iK5+EArKL0X9Dsl0P8YTg4XGZBRInC
zjMkR19YQVbpURrDwP3pj0vpP9RKGcjAomyjY/JZYvcZW+dqC8RPzjhvTp2wwc+1
518Y3WVKmgM/8kaPXzd0iU8ghRiD7BMnwugxoH/wLorZw7vIy2g7EmPOkJWGfkbk
zE78ZYZZQcKVZ6e2DKRgMuTlbD7z460Yc0ib2qioqQJEXe92neZsqezWH6i9c0zT
pVlJtYTwF60QMj8xIeprnt5tTTEdq8W0MgdWgjLuiPMwOqSWs/dmWxozZEt9JtPe
Xmw8f8Xq5rhv1zNUuG1y8M9UlBeQ9BcYXPsoyBwH/oOAqjRMGp39UqTbyj3r71ic
yC62qcD/o95BIDBBo9T4AfVBF4nrVCj9T0y4148X7f37zdybtMdV8RYF8JHasweL
hlAPwvqy4k892/Tm9YKAFf6igtfoloCg1v1wNK77SYne/ysg5a9q1PYReE6qjBj2
pYGVZP7Tb9pTJ5UkBzSFseNAp4u0+Zi5nDdaBvxG5AOf9dyPevG/R3sgFa+LDXNy
X4EM13XuNgj+38feT5kT/O60rbRTfARV1/COClkOBv+JY2Ows6kccN/ltYn04THr
+Me98dTNpl3jatRcUWOjWNRzxuHK0i3RScA5cE9MMDPmorGfjjcpSbPFONFThipV
Yu9BD6+jCUh98a705e85+cEpvhHmITGD/W88DuVml9NxYY0igmCFpJN0wU4D7kny
xbIGqCvQipfYiJfs7S1rKQo2N3wTLa1EzcskrMRdsGPMf4gSLqYhB/HPwPP2mxu/
sPDNnIODkTWxg1sXzS/pZVaAC7atuzcY0Mr5dnvAyLcMf59bFxxj7jbdoFpXDVaN
f6Xyv96arivNmVb2MJTogBOwpAucnFm5+zupey06I+DYJggsw7FvBd/BJHGU2FGz
QX4sxhQzdc/TYH37df/shcAGmBejBpn1qfI1ut6SBl0l/J/T318LC0n12D7BNABq
fEQyHP3KMLiDWkhnJlahpUgnA5fkrzOIkWLfXdBc4Lx3J1djlmiSYqvOx4tj3+8s
k+V3EsyjyZfGHumh1f79F0WYDU4J1gRPumRYgVs9gnVNbjE7LjdUujMsG64EKrJc
XtD61199ek/QUjniqoYLc8FzAjFVSZ9RfVNPh9UOG/fde5IP0sUeGJobGTw2FA0v
+eQ/mjIT2JNDvc/ZGZMzB0h8bEjzUrBFwnURR1qL11+KdPmCoz/Lv9aJ3JUEaMBG
T/5+cnyAmXDVIAgWA3nYWpArIDlV/2Nvig1m0YLR8YzfKDfY0axSfDQl8EgAY8aD
NYr70IuwJPF6fH/KXsNY2NDLjOkODJtAH9gaGTxQPFNrl6r1/0UD67bf3HRl0Rh7
I3oFlKR+MiXmZRjV0MWi0+0yM+H+EtLrsCFriA6r89MQjuYf6MqYa4RGfOIvrtGN
vKIOBKiX1bAvdvBB/AUY5OVG6/jl7H+z12bd0TaUXtR1zLqol4ozQigk91AYPrhA
aSwFdMagJln96wAOdmIXMt/zew3cNcQb0ovX2uWkGQaRAF3rTcMTKIRrrK1RkeKW
qA6UdXjBYCtheUYpki/qo3f4RpwYoZVEfidF6XLjXbCoO9G3uTbq25y7lyHRVYzo
9Guo9BQ+WjdAfhbxpFlMAH7ZX0FTQvBOhq/Naue1LHLZgZhW/nLrbJfz5gvbqwvX
G105sn49VlynxR9q+mx+bx/BsrbNIKD04u+nuoFvTIF/nu8xEO+ubRzDnkc1JILs
eRAiHFeFBh+3YxNybOdLEG5fsRiNaZiv0c/ktYUXvBtEx9JdIlrrBbN4unb/o9UO
EqlZae58wWDUHnAbA5YvQT3ojsiF9EKAw1rY1wz/l5pOiJ/h/GPPNyU7eubXcMVJ
PIOxSvp6MpKgKr3T9v483vt27+PBOLd0biAtYSx2PP2+Iny5UAbHdNxJFHTFpo8G
E9oPG0gPBM1BU42xpB+4LHRcq5a2xTOo8llAiB8Z1+gh5KLkSsOoxoYEC9Q4Hnxo
9Zzu2n4Y7Y0QzvklxHVK38IZTgpB5fz7UwA49SO25WCFiUBE/u+RJ0sCauh2fzgZ
vYH/LQxoCMhXwIs9ppNtZmRdRrLBsOXE39OKueOyB9pTa38yJiOaHXOkEsAFo/xE
KVf98vMmBdZzYg2jc5vNBC1TN6xdcQi46UovRdcsHHvgXhwIIpz3rm/IRpUrVX6h
wmb/D8p4zFHjPZhtkUUAWPc7/i2NjhIbz/0znfBnyN5I4SkociMhDjLxWbFJ9Hm2
haljkCZgCKBSccHvVFm9GionhOHNyzQwNuuA0tjnjLIptdzxIc+eAIswsKZ97C9g
ghDhvwW0sLFlkcxFWNZqXdcqh+2w9eMGevg4oFnEQEO7iM1ybXwvKPmBAahwkXL2
w3evRKC2AHNQkXsCCUAlpXdOCFHgcjkHIKmJAAsVsbV2cru0MjrewQ2JvKHYntrs
6VeIs6kuag3Bn7FqeNpR7t+2/RI03JSSKm5jEUuDml5AfjfCkTWtpX/ofxujSAs4
YdI9WKhSRQ3afvmQv2eVXAug+WUp0znjwBoKz0SzL4FfdWmlGlVYHZtnssGZSA94
5uhqYPo/PqVIWKKNAjdgpmXc5LNJzgekRHhoN4emAr+D/ctDHBdThD0RdHiCxpko
FtfAaVnWcbgRFkkwk4HEmlfsFGjExK8zgm1SGnhc7S/zrXLb/G6J0J/HhVJSA99W
adFaANJGKGydtLnRSDH2G/7VmUUud2U17MEXZoMiASILFuT1sP0LGEwpMS4z8kP7
+h+YlIvL+IPX/nzPjNiCxBWAhrS+2UxvhO6iv+mW4FXU3Q0+SzGV5uZs8x/0UaQl
7i1is9QAl1US39d2AmMoTELkU2j/Lg8RYRmxa8mR5wavBOQQRURjwI3rP56lrXq0
ddeTphypCBAunjQTDH8pRlZfU+8RTxpBGi5kRS3ODs5ujnTZDfiWI/pZl+FLeZ1D
nCpavgcuobuTaLl1xJtjJOKU8x1P+OlUWfSOuZ91ZxAgPQZ0C9MiY5/GT3d5G53H
/npcfjLV1mcBnDH+b+Y4BBukn6GCDjsxbOAW/ohxPwW2OSZDlz0kDU1V1ruHLRjU
7YanKf1PSmoGkYkQOL1wqUbZhPZwvE2h886VKrqD9KftUeYD1VUtYrbbDtuO0Vnz
sZIK7THJ4+dkkfNfcxso5/jXFRtLpr8YZoNXAwyB5Ez7TNMvLPTU9YOKlYegj6Xj
g5dWxhBNKN1u3/q0Br0aMcsGEfhLKV0Ag9m5X5Qw9MRjPsH29MAORaOUxYgeMy9J
8rnPwc0lO0+o00K1q9YbSk7S8rXrlNqyAz7b2t45zg4h2QgpUW1fFYi5aFZgggmo
o5uBxagpknnBs4FZzYOSBQlKCXAkl+yhIQjH0gPR12VmmlbcB80MerwYIn2O8HWa
0xXLjgnJHFn7BdPp0NMPUEh5HNQ1T7+V1VAwQv/knDt/P1hbhgGG2Qg0PJAn6pGo
ne5l2fBX3MIROLEQHRTSpiVizjSBJNSf2FlaQUYecC2K9uqUrk8VuGfnolpp6Lqw
Gov/b6vUiEFmF0J3jcZhf+R0RlBUf+PNghrdJsR1Jl5F4qg76f2o8b8oITlwiaiL
3Xddo0iwA08qS/TaBr9DHkovgw4oZ36ZNgc37HuxJKYkh8SFuFFsxD7YW84zCzB7
2VlZsFk8hXkObzGL/q7kKCVL9BqGc2MXMzcHwl+7brJCXigbk8jkglrMpoua416D
0gyy1NmMONNGkoceZgv+7iBm7iYUsJ8wIbuXNzi2SlPCT18CYMcgHUFWtSyiXpYM
fK+iePCOuV209Q2JQkDbyDZX19Z1yPAiM1LPziX3JyJvG9DwaaZOoHyJm9b/Gc3D
PIOAcstDG3/wiYeAPEc2UXr/xUpIU8NWUW3gm2Gswx4EQWh/s4XmVOtk5+Dvevlv
XuLAz6FKvmsaSc+ead6uyE5+BcVw+cn6oeTK2d3366lzV6Z8TzUjGTBTDx8C30Bu
z0eQLsZ7ob+FVqVj4WLGsSfJUZCoP4hiGEZWaY5l3cInGh67HUfnABzOUCT6+ncQ
trBB1wxuARextrTEMVNatN4uumHvuZEvrr7V09A03mf5MgsXjgbZgVInfRZO0oUR
rNytywnTPY4/rabl2E+bG+9A1KvfLgjB+dko+BcTS8swQ0+3liPD1163ybIHgsia
TfzEcnNO97bWfzb07w7u3AHscYKxxwmLW51dlDOCVDazY0bPc6xdb8/CviwGGkeG
DYom8qsjYLeiy2rjRM4Z/E132gVDIvrXrXA/VoHO1t+A5jozM14nlEM/AXS3YhqA
GsNDLJli1NDbjSy/1VSPBC8qsrN0tnx/kTvVONuzKFMA4ed9kJoyDMUjEMNyGdyK
pi6TjwMK/O7JJULDmpsCYdqe6X9GUQi0pRSm9XpzGjMIOmuBpnI87e+pvCn0hDIB
/1t0p8o++zCxtwbDSWK7X+NVgcbDQD6klldK4Tn/wnlksqG/bJTLrVwpCsmXsfGj
y3Et5iyqaM7573UNmpD4YWl27G7IB/WdtxaLT1+3XUeaM6BdnAnj3QLG6CrQkhn5
uF/Zdy2vJ64kl6G+Xb9Go63pqYAy1phy5U/n0A8+dtV1WX1aogrELvGLGgacgqSs
A23h9H8IvMJsozKW4S9iXMVZQjOCKykdlECXqr3IurYXF8dlz63/X0DhMwBgHzgU
T30HEOyxI08d1msYo69QCc/SgyTZ3GZ6o7Unvd8JzEZ1/jSJ3dMSDDgrhBd6vvgV
al+bsK84JkjNIABxwDFY0g3L8NeY1yRyhC40Pm99Vuhbr/YaUSsTTN3YipbdTtiM
61TkLw1WxK3xe6KVsV9ghC3SnVH8D0iqDkqBtbaKcFvLTkKXdUM6/5OTxXfyMORS
gY3yq4Pkw2bf0t4sv3PhP6KIw9hbTmdBAe90j7sqywXUmkAntg5OaxXEWKA1CE2w
+hwYih64Wwi7+R+WC4XyW+gTLCOCxAqwHstp2X9VgIb3OosR7zRRn4u8KE/ziqcf
gapdFildTI4R7hxbT/TNUMRi37Fk541PdYsXAX9263bKJrsNzIip+Nnfmkf9R8xr
PEjc6MTctbSWCrZz2lp7KakkimcyI1e3K1leEvXxLW2JRJRMK80eH29ThueIt/ve
cAwAaNWZNpZlOIv21X4u85+g6KmkHiXlTxSrDoHnTQtKhC+CGXmv8AmRquaJSE5m
1p7fuppZvR3gdcPEwTL7oKPhGn+2g5slR0krFWBcaRU4LypbxHWyNHkpb8Jeo2lz
hpL2BfH4hDXo7CwtG52USzZXhu98H/JoIFeJei7sXwWTHf/nq6DF4BGA9MEGP6rk
Dzr+CZFC1UQArmbhH6OP9Kybr3/2od2b8GKCk26nHuYs7YpwzX57BLjbdgN03y6L
BY+wxtkUTNC/4i6XzBovz33Yj3TwuyYJS1rItUjgBYsdTiP/1SElmMVXRZC6E4aL
eaaEFw/U+1OSIRilFg35Y5vc46DIIXN22XevE6+g+noF75f2jVVgBzsXxX2S6T2l
Qw7MyAgF63fimEUeaNJ2nPIqtJdoTlV/Qef/QXeKYsLo9jxyTXm3luX8NZrxsi8y
qZKbeRlXlH/JSUMEfk908q6b2XIO2Y/NnAJyJj79s0PwWXiHBlTTw4iH0GUA+yQj
Q0l9unK083zg5V28qa9papmcjg/1Ltj5FMOvsQLUWNeYF9VYw9xY7pFsY06O2p2O
suiysVE0YSC8QSAA9MQ6/wAsVWWw7s1uns53bOO/iJy7v6my6yrXqLfHXJkqhvxa
nsSjwhQ0siTYCtqwDmtP/QAN3ylEtDBlVemO2J41qyLnRPASLFA32IsslRQnIIK5
ph1Dw7IXz1wofcBo8WJPmVpD0V7ZQXDPFrOXszRI0zJwgE/BK0Gg5yF9GrM/fAaj
E0EP7ZPPuc4ReuNOm61B+jAwiIYSB6APbTWof39F2ARVfw2iwdU0fE3DVITDP+B5
ELoluI3hPI0hD71iKCJTMSpkPyBI74LxJhq5prqBLN9ScIGt5LqUG9YqfoFbQbjo
WAWP3pqGokrtjrkjabJbvsO2dNuyBf3ZfASta1656LOwQPDgiZvZFe0pp6QkOVmK
xmBUsm0U8ob1s7jxnE7poG2K2vXcMEtaMMAEAEuSWNW2W34DoDPtic0ifg99K4mv
xw52xvQuR3p4FoiODXvvUaeuh4L3zf3uWE6DRAS/NYHfICdF0cBfkmLyTifqfyOW
P+wG4cRx2dsm7KUgryNN7QsWFGc8v81v3l6WV4zLNnWV0rdJcDxlMJfVs4YnfLly
BfQtqpJrqG6CnKkKqZHSoWvNvl9jqtRrtA7lTLa25aT5x6uR1p25iz3yvwqXeAzy
i566sGhj/0FZnmIPKC1I+aJH9Y0dndnXvQER3K1X5tnDx60JY97AoS6vApq55mim
yp1Yh6tQJ7pSGyrNTKjM6gfkPbB5fXmG2XIpZMuPTsj3OyVH6JyUZIRY4+h7i4tv
EarpC0k7cLZZ4BA4X0KIEu8zIXtO2Mnnoefb7aD4qvsef1+SM6wLWjRnckevCv66
RU7rT4LlkDf9TlkyfPwLV/pzntYBEpaTROb3HlUPjX9g8wXK1oIDzIvWZ4ZrvdIi
QypbvFZ6uwdYoCst7dBxLT4ziJdByrCfBMNPjcanUjrj3351bC5jLh7jqMJHO7nf
ixrQ5YBIk8X+XxQj+eugMBJUnZ+GpKpApb1LOeziKX27yCpb05yQlrkqePPdOkUC
Co19Yl4vVq2rad0p42oEw8WGQnTNeVbWsrkG2d67YGH050kOo1coKLjJQvtGd4Oi
EAACFkVNeD7/NeGZY9lh2vUbnsPeFZwicxgN+bKximyVZWUKtfReD69o5NfkGdbQ
pGy/dt03/8VxSloqCyilv718DIFtOJoY7+UP4qbZ3yjGlK1AKVVBzmKzPXGT6tHt
sxArSNV+ii0iYscU+TJEZYhGYtQrl1C5hPuh3/Durti8LXqYs6IUWIa5IvaUYd3q
rl/wXPKuobtKEvfWetNGUWnZEU04qi7HbuCO7/elTE5qJhU1RqpxWINOwKn9WBHJ
bpvBMYfJHsyQNQyW5V1Ady0KXcYJpCy6K6j5dP1ZYYzmN6gzynRZePas1+oDByKa
B+1vgfZHC6UPv5wBSCJNF/OsumnEaF/0r92U+0mjFvDb5XblNl2kktGTxZYef8FL
OZpKhbuFRdNR3kRB9FsNvkFgg2jW+SVAlPXVgNAiMBq1n4XE7L8xCPMfqEzfWIMe
I4iAW5vlD+7DzyEFqPPZmwOjpBmtjogTrrDmg69k3fwMdQzay2hfKORof4BMgnsa
AK3k7KaNel63k3dSNzVjSa1TCIYjjHe0Fv35jHHgo98Mb3q4YJo+Jda31M/Hjsn1
J1Vl5qdWHolG4DBGm+FHatghFrZrw/vhQVqOqwMZb47sxaQklQTgfOqpu/lor4rt
paeh0I8khx9FlQ6gWKfyTs36jzFHibgQKtc+ps0gEJ7Ps1dAO9Knhz42lgylVNE7
7+5mXMhs+Rl/dFFYddHnjfFiEVUwN0RHUYa4hwNtGkVUWpA2lL7AVKJFobjqxjg3
MAfTJvQ0zYVL3e35ZNaaesLflgPvLsB/NkHFY/fxEed2+nEzwmag7klQEPmvVRL+
y6cg7t46J/L+EK2Ha6eHUzpEYxAoWUMwh0/dQEbTGdX+zjiRMmAeahKRAujBuqrq
Rk4eP1HMKYlx8oC5opDMvwShwOzT7xsnImsP2qTGbfLS5sQuON11DLWdwpf/Hawt
DhVbMgT6DWJ/0dM7csdew/OoPd/kPGz9VRq9WL3jfkOowyTo/IiaMPB+v9N87qD8
aWAbx30ydXaCl7qaOd36pfooJZQ6k/buD5RyUp2vID2RdVXUmBNcEu0/VJJigB+g
BhLqH1TDeOuZRPh6RNuQ+Kez1TNHoCPtdfuvK333YzHQ3fKoMsHaYj97ofEpfuYu
26Z9Ec/O90Bhz14DH8v45E163zhZRoi2Sldal7dbVXbGwiNBvAxFtDfNkrB09DZZ
CR4WwALNdhOLevePqnV3Aoz+z3mGIQ3FinCImakiK0W6I4MrJXeRNl0yuQ9LqpYj
+QT+LsudUIhKLTT+3b9dBogQTI7RdeQppEHwZrV1ChsTyGWR8sjeh42yuL25T8TJ
UTJwpar9Ke0+uRuv3U3j7QrnndZnaMPwOTQpt9c+2t4W6gVhJLl97cJYk1PUTP2B
H9J6DtyBmeeAUr+MJB8oNzIHR1Kf6VpsiVWRaju0CvKS/sSsrfCchoDE6Bd9WF4U
vM+gCEkbfhVvJcSU+pAO/GisJ3nYMHW5pfOnngUKUzK9NgzC0NAs8HzVavEhsNcW
QxWskxatjA33mpe//bo7aT2KXJARs1Nh+LFgGWTYzCrhfS0jgf5+GOiP2RNPkRDA
a66Di7V4rYunBNyCxuN2hfeJ4dhCkBIkXECfUE1grgKPJkBcll5eVedf+BDRtOVa
p/OQcdBJoeTHak3HkXEmWpILnt7fXdPHu+PjnV3vnQ3D4fp33wxFjIwLTbN+m0ok
fCmoMmIY4Hh2EEP6JYuNErGEKv5r/c/LHBw2rpU7oE+ay8PhpoVDtoxw+hsKQ2L8
AsBTRooouxPRnxOHt0rZ+emTVWMCHsOdNCJmCu5DIOBvWX24wXfcfigNI0O3G35e
dsj+WwY2RYdSn979gTdtTjB012YqIhpOXCG2os/5fXtT4hTmGC1ZPOU2P2rODI6e
F0i6g1wr77ZLtETwrEvfQ6qZ3VLOpz9xzv+jHdobcWPI31hgv6A2Uct5DTKwoQyZ
wARicGNxXX7OJ1w176tgRwA19PA/WUEECBCW9Y+9Q8eewMf1c/ZOzBCPRIkgDU9b
HY749j4Mb6i7AR68yYn1IOaVoXg83DxkpoJ4aOpY+eItQpnRPnFPh9yLFfsbLWIW
+yPTHzDymrma6NPNEEA0zt4NWoFhzybyTOPopBs/grNFbCe5o8KLqKCwXyGBvsbt
RhZCtFB42WI+uzOYGvUVPbN++tORWdQt0xcule3nohV/rhF2DkxzkHNbsbmMjKE3
2Nt6QsOpRmliM2KR8Vfrki5Has1J7hRQE03EZ0JkvKGvZa7qjDtHwvqG4b1NYukW
lLGUzgXvU8/sLENbF4Mi66PpKaaEQu+nqS4s907l+CkVkCEY1/1QqJSQ3ht0dwAP
rn16ux3iC0loDK+CGQMSLcWH6eqROZCr60sToNN5uuq7ZuCrscj0MZmSZqC0TOMp
5mna3lj2B8Obrp5tv60D7cav5x+/SPU3iztyXDrMFl1UpJK/anV+Mp0/7fwtQbEi
+6fjcjSh9lZuZRkqcg9Gonm8PFWcaEj1niAnP8zQ3Csb7xPaF04pE4zhPg6HmJiE
2SPb3w4fyq0gMe1wacP6s01B/TJ6HBau2TOCvERZmeLJIyr4J5XzryDcYHuYQaEt
DkcfnaK/KGT8brkBfZ37qKdQMhHhfQdVI40SIBlyoOkFuP0k7Sr9nvk7KwW0vNqt
r9Hdelq51wT/N0BCnvHHFC1aWM8667zUdNVoeADSLx65POJh59kP9VLihQ2qH+kv
kuWyNVIJhv7WmYuoNVycFvHiv51w8YkOORj0ApDfUTsL7k4NhUTGIGwM5AZUa0Rn
ajh4hNVex824bCHusRcNbc5eHOTJ1e9lgGZlBaHJXEJQJ810rov05+YjuNoHshmT
PiWYSlXCp0gAVsxFUhFNWK2TORpb1Z2S17RDs870EwctV74ELTD8VI7huGNUgaqC
k0I4uo0zjuMBecW6fIOUyh3KK52EgPS6j5Hh1UAWGHgYCzpTjVeSSSQ0C6MwNU7c
9MdFa/lKvUrfTj+aIvnSO+/FwtGwQRTQH/QvlETZuaP2tGRLdeRwtBlZFLfjNWPP
28o6ZIWjiyIM44fPtJZHzoDQ9PurcKkHt4cSFJ4+uAYS68F2mUUUNMVpDXMNvUub
KU96xb674Ak69/mY6YH5u6/faJslFYml1Fa+zeKSs/xMhG1Z+hi2h6+X5wq2MgCu
Pc90i3SmZqbgr6ycKJKz5dI7CSpiUUlITX4i+1Eeipv1X9I1RMQg5W55n88+Fo3B
MGmIFXq2niyoqmvr982T22Ybi7FEkiver3vfEJdhooZj089QYwua4ztDjQuYLk4U
DPNCaIAoIzmraH84Xyff06oc/G3tcXDk7gVzAf20fgbriHZqfkZoel3JgvCblXV/
H3FOXsmxxtsRGA2F7pRB+LkMxBsTWD5QpmD6qPFMDpeWEIdhbxtsuYyFKbegVX+U
47+9FlmmTZ98yMjYHN8QIVd1KTrfjHXkifmNIWPcGwrr13XkWPvkIb6oQGx7anX8
gTqfR/mrxWNNE9n0Yqt9Q//vuMwAtTCS+6WyKXowF485L/BS+P/LnFZXiKSZ3O+b
4xJd7DWY9OzqhVpnpLj4v655rpbu/20qLIPsWPzhHtXu4N1RNU3PXOfwOxRxtf2J
DbDIQv5cl0VVeg2wgMKCkcIM+ms4ungwAeTI6qkJnVdLu2sHKea6COY/NzMDLyMH
fmLPT0U2Nvdzh7c6ipCSrSsuWBX+2L2WGQTK9Tg2pwChdSzLaB6i1wEbbT7KoI+R
bnh9I/EEGHRFaZZnfy7V5h3NDD/fCZSgEBCfBnTy7iJxyxRAYaWZmUSFyrfo/dRw
RZftDxwXTMCpssN7wK7T47N1ifBhqlA0pOFZIYj+aHjjkzHJCuwMFP1iRFV7fPwg
ZnErN7a3kcRJXpJ25D4/fBOALs01AL+Alims4UkjXJjvkwO+carS4dPETAdI265C
E1JC/mzIF1OAWfzYCPmkbHMqGYY8MoQIDt4/7A6U8hChRxOh0b3rJSXjXb0/SbRx
YDblMTdxWduAjDwaCGtxReFtZ/NZf+ChunwDYNSHYDJ0O4BR7j5cRXYErPDOtNna
ajWzdku57BN1a1SV2uHA7GYDQo/VA3ul+GwKl+9KbqgDbqTebsHFDJGKnIC+WiwO
7dSJ808cDptlE99M28T55ge0x3QVTKu7bUdESBLb9mVggKwmeNPDXbH7qMqLpDuI
lYtrTqaHd3A2gFbZ4F9ENM57ZdCpXBODi4m18F/aRMqzyyW96xfkxfL/fkRDLZSN
0WttJIp9WeI/Z+5ihQhaepF85WcdsRBCF0b6k4hd7Uy6+HZeNmCtJKHKmKfi9/Ah
4CxU7EJula72HBFmSFK4jjU+zIAo2cZmhlkukrS2Mff6qyqUs+OEEciGwq1nVAcn
2K62VBjB27SkFStCSR9zqIWrcw6B2zaOQiM7BEWpT9sRzS3Q/3xxERtLrcWjvwWN
kD17/8Pf2rcPGbn1+hlpSLpInNjP1aWABeZN+jSIKAv3Qkz+GjhTVgwB2JsjCznQ
2FgHtlbSrhgy1hHJ6Jx6haOX00bNiiTHtvsJs6dujmkgrHIy6/aDrYWXfXNoKWtW
5QKaiczhQeltZgKvXUgL6601q8Ctt1v2ePwzW/2OD87iuex9ZQIMoJOWNN9zCEBN
i4KCg1FVbU9PjAIHMUlpxWr4IVj8nZF2DUrnULzALYeNAUVVvq9E/lD0jDTw6grE
sZA5VBLPWQMCvp429An+onosnQ2ow/hL263stuURr78sAsTTxMj2GwbvPDGI3QPl
wNl2xrWqCkxtInx+BRMMS+Rveqk3zjhZ8PBIhbvjBCBm/F0gUvpMTSWXd1ysqe98
YcqETMK7wKojR6eKI+b+DPJju9uJI1r9CRdqPHQ0syJ8sLi+5A32ZribjHuzxQo9
z7ujDdQ7KC/stm0IZi1rKuW5AIqecGpnaiqTMnfGOMifpYwiXterPdE2jl/xGKTX
ZP7qeoYvkD3cMD2GDZuTmcjQw+K0YAoHaSVqe8wgmD330OBcKjy4paocwBNUDlmA
HK7FnMkKPekkVlbmj6jiKaKfqHTLGyUbMhNZUG6TUS4YMaWEQ7mHqclsEgSed4y8
+tTfoLTNhNl55fhnG8hrqyUhRcZoHrx15Bpe/GpuN99RpbIOZsYQnxjbADxHCxlE
Q1Muo4Ps4rIDNIc2V9ohwOPgV0gR6CM18YxW8I3suPcG8WYWlktssORLehqQQcSM
Ni4p7nVBs0QDPOZCithIL3TJoqPVkwQCOttyQ2POMpQaN8ToOEBP1F/5udPXQncX
gPu1lsl1t/nnE9q/G1ZcJuMbqcfwwby7sBsc/xy1xDSKvaExn8IiKOUu13J+MWdH
70P7Wy/IsOpO4p5n7ynDPrTKfm8hxh6bHWJKAT+1vbKv+l61KlEEj13xX6AxlAvH
L4DXUI/944DMak47c+LH8QOWPcWmhDUZAIjeQQ8gxECuL+b6Lzxc97KA1UxjsMWq
6XV7Wbr7639m35MRWMIbUC8xEdLDLcaP6tZnjteD3NkvODZMzwx8dgKcthGfahSA
tCRK9irEhs79c+bWsvCH06RLKwGtTjI9Ug3YUknn4uCShxizaXGs0GGU9hZoeLT+
k9dMGh/2lRA/6vj+n5DTLgTQDPOSSuTL2C7kFqNdjfPwhXU/usmXX4CP09Rt/XPH
MR5KdRd4eDSEtkCFtA8G1wUCLsPRZM5ePmGXzPaZz1ClhRr68S/PCT5v6yl0FcI5
eGYy6B2fF1dOpELdmfy4FmrML7DetnjxwtbfV8y9tpk6j/WFj2UcdbrUva9/uMcF
o7Wp4ZfwSiFP5GVjd881nVXk/jucIrdcYdYOnE2X+5ZDMb6VYbkN9QK+GHi9epTC
la2RLOmv5rxNlaPQ3JSLIapL0dp1lNd5XR9xkT3XVGA5pKVYsgyl9V4jbZ35WDjJ
yiqWwBSkw2ZFHViINPiBPlzJ1PI+EfC73wxDQxWuDxf+LaP0Fx3wWTuU87Ih2/sF
W2tIsDKZW1gigE16KHnCLyCB/0eMSXCHR2D4QOODerWbkDuB8QaWFBX5O0P4IV2f
5fC70zaaxuiUVgzHzcFZ/nyhw+UPIJn+2vQYJ3EcaRAk7vw7WRomwW9BOmKcl50w
HchZvEhGU3rdZukWOh/kIar4tNxIYd5TCp/UmDw+LxlkkiaymqZXvquXqncwyx6E
dUMhzm3Z/e30c9d1YW7BOfXaHN11JYVwNbaprRWJgod3vAY4iy8qodeXekOY8tz8
IeTgdUQHBC6vd+w/TJYzMbGLhIjdkJAfn5JkWh6GeVsFaXdeP/eOzdB2mn+Qgn+u
/fcQuz3G29+O8mJaVVWwXmgv2u8HkIs2DyA9fAfocp5lZWtPM6JtNJLD8I3FMNZ4
h21oCgFaWgLQTGvuAwA9pElIWtQ2LEuIYOe17P0qr5vF6Ir3odR6k3ZwSkWdyyYD
CxEbACbHxCL27qu85x6yAo4DbHjfcatVuGbiAjdLGbST/bc5/QQIVm0+HikTB3Wl
ymbzlDa1IbOE8DD+CMZ+A6KahUfp13Uky23LcBWlX4mgSNRsuhGl4TQI33HSRgb9
0S7d2NhgFkE+w7UdaS4yT3CWxJINT+z20zMx17GMTsHyfAz27kHdiY0GfcZfg8z8
R5qLaMn0qh9iChbuZ8ZXf2z2uAHzz2xJPoFpq8fUXTlQfdFsfZ6Uh+t79uP6gD6I
ZPK7eENHHFfeE2HcjpnvlAZ2GfTrd2JBbRWp5Wrq+sJnixKhuTxxy/AFXXB+8Hr+
rKOM6wMiaEUqoWY2gsR8p8UmSjycMNj1c9giPiK2rhPSbKm4AY/XzmR+vUFt2Hhm
Yj88LFrVehOq9PLIFi9g90QzmdvWTZfpgyGqaZhsOzp65LlQJ76/z8JfMDfmnVvJ
NS3epid6LF8un5YgdkRhTrsFouEXLtVUZcK6JWGbVhLlWjtwM2JIIY4FuywJQDug
INUAjrzbYKoHQgwsnKxa67ya4+Lj9imKhzVTj1bF3u8BHLW8arIc3zPthUArmuoN
r7ca5p62HMBZ+kZ2KabNWZoZxSddjlPmp7Se5qZhB8W6QZ/7n8cBT7yktkU/ZCKo
shMSPJqsx6lL4aVgNLjIYgJlkGbFd82V7dRZ599CF64/vGMVnpCvc7JQYb+oeiJc
8SXLJ+5uF9KwZ5eQnbU2SbqzRuFlWYCgog3SatEBLqNlOYI06QfypzOR+rM1KkWe
gOL28CqORl2tzaA3O6OOTanCVG5H+RooF/DiJ5lfyPSrBm7/eBdAJ5foHHyRJfuH
27jUY7OdjALQ+VIOvaebCmHTN+T+Ga2rqcR7TzsyJVVsBEIhYUsYC/7ZnMaIY8Bo
ViCcd5QXhMVbvbU1mqRtcecvYtjGwAInYEqRdBzrKnYZmNCD/QgW6mjkbW9qgjjy
MiOL9EJVvSSUcaVQxiX2XWxGRGR2ozMzC2u0YCpAtGDtMygIZAslQA6pEcsUh48B
qS9cAfXR0ilTnScZ+ZxpZtBqTen39LQfJ3J60T5LF5aXF29/G1RnBrnATmWXsVpU
UBlQiTZwNMosEAlnZVRTGq4AaQUxe+sddhuTSGTGB2vvy5F6BMQf+zoaDZY0yyv3
r7Z/iFtayxPm1Pl2Rx44MeTcNHQRKcF3DnkM7fr1XUvDGypwvZDvDK3cz7+nSpob
l4hwynD6EKSGZBnT4VswkvJypTQopOmHdK2fCCAMuCgzq7E8vkcmECR60+yFojUN
cQVGpVOtHhae2ssJ9zNLPQVCZ2Bca4uPwOL8jF8sDywKU/6ikFztKBNzh4yRcW3E
Xm9k8sh/6hu/5o45Uip1fcykpjGFl2mte0Snps4uC35uLi4OXsUzC2LRvQXidtbb
A4NMn3RtkYJeICWLXwHHsJqxAwDjEFwXaz2Iac5t+bDQGdIE/jXj67i+6DwprUB5
1oxvdc2VOFg8p2v/REhvDd1RCw1xwdARgsbSI2/Q4Xn0gRa8bmrtdVLcn5gqJfT0
Mw7LVkI2Jpr5/XS3A+tke9ogQxeJvhNga2mTWWLDfXzf0gvCb1L4Z4k1soCM+oXB
AHSmnQ46a8aSlyVRVWvzz+uutcwM7BhQIMn8KUCwcHOJuGTQ+OQzUVdhIR8mkeN1
8ogb1heS1yZKCc93UoOkosgYSc397DAjedifZ0S+a/EL3i/YIHecFuUfPcizjHGc
/mnfRji5KrRIH/bjMWqgeSL1eSBhI94u/gmY5o5Wr2CogTKM0U6HEyNWfcU7i2jr
BdM/RHDgL7rrR+5on+dgOvhwX+/WRw8hp8y9P61ZUyaF8y0O2vLGU24V1yxtHJlX
AQqufZTNO0wgY+ZS59Sviy+kmkLM/vEUhEk7HzqdA4hO3Su3g87iolZRz01QKsdV
fPwTRPt3+4GO15vYAYMJbgeJRzIs3pn2JKROnmgFKy05yTbWtosx37Kj5IotbmzW
m5xI1Br0CqicfhbAhfkpZrIV9/g3XW6t+Q+XmE/ynqJ44yH/gObCkS8gE86vB+2S
QirhL2WN1is65fU2/In8vUNCx+IhXo+V+QhqFtd1XunjlnuFb/BVfSY0BXVYFdt8
/aevOQuSf+RPO2d8iOTwt9y3qEx6a0shaI8vcQ7TQh0oRVDJ3dk231d2alh6YmSI
oHPk5hx/NDkOINuSRFJLtmNJvxpIoXizDKd+UEJ3aTXSqjW0LBwVa2618VjZJjJG
4Gxy0bxXxdKbBloNVMDbjjP0UImGq/mjhh6MFyWK61F90mokw4cpR0pWNz9dLVFb
lWPdzL8F6zsYxB8Giebh5V8t04arqmW4K7gT1JC8vO+VocidTzvx4JSra+J6oj0W
HdGSQkvTW8nfZKxQnq0q0NZrYsJsRZ7dP/k2LkS5ow3TXXuB9KndKnc1C3qM0dAP
iw+Ni2GH/AETa/lMsJPykl4sYHjtmpw0Myf7JinPrVVeIWnMxblIMqtrMgGrQmlz
Lf9Bw87NS7jq+AW6zzeP1+jo3xh90Lt5BF9mrN5et/B4bbNW26xBA4jqpB8yiu4Q
a47+xjYL8l/qTXHS6eyqR6YGvVw/u3rd9/VP1khINEWDe0WE4HTOlYvdC74PRAfK
Pi8wMUNTWbW7VZS34fehz12Zs2kc1JOkoql8PEJyJfYsnqXEpOOq+X9lQ2WaCjbi
Z/Dh8CfkhIOuEOzrpufvXEmVe+tDxr0sDaW1kZrJh9SWrS/3MgcAU/SoWJoqCfmM
lC/EBRo2qbQWt54giFShg/ojNBjYTWBC8ozWrRwlOXP/rHbhJaNv2J6NCHKOJJCV
OuXUxEwM2Cg0/gjnle7ApEzCRt95D7uhkiUYLRiMQ69Vw2+MMYSDewe55qsoLyyQ
PZ+3NIXgaWGAVYXQQIuQln6ieWWNUICOJdrFE2p+F7Kh7kzIp0gvPjaPSFyyEDPl
rJFBkJ55sibkyuQZLLXHseci4/QhX/rLM7K/Wh/T3l40yZKvNW/8qHLO4xl/PWpa
J+uAIyx6DSmM/V/sNrDDnaleil8jrxStlC7UCif0m2NJ5A8n2oniAuX8MtTBNOZX
EWUpoS47wwcN4jTOgNLzCkLcyodMVACnzzQpKMRZC9KknzYrnspYICrtEoSpImDo
rRGDhHC9OhQO92AYHNtkgLEWQFnC16HLIj6frzuMn/PF/xiotJ45NPT2ZX3U7BiG
nR8DL7muoFREmK47PGN4j6YoTPfdxVppeStY9qVLTYpKivHgPyhamnw3nBFVgsRT
rhHQ5iGI4yK2kBYV34BwTrYW4bg1dlTjA8PtLen1fLnPqQTDInmHqaUsIqZKurlV
uP1rIkWWmbKpzeYFz1kPKXZwuJV1U7YS4zFO2khGYM7yLs174KYgIahOOG4UmDSJ
GTG0GE5TItG6780G3a+vZ9p96ENAI7Omf+VX8x2NQ4YllRz/eo0aOQrkpzgl9FZN
3Eh5fonwbPmF+OkEd4EZ9W+NZjRsFvHNBEXq26oquCHfo9YfZNESnBDoxpqN208N
pgeLOJwrAmer3X8begtTv+zia6Zh92txscWZAJlRAkiKTX6Xcd79oN+XmCU7+YQZ
3JyfQLgLqAoHofKSenWaF7LQNxqQRVBaczDH4w6RjkTzE7orvPB5hKfmTxoLnCN5
PFzSOE37n29etF8TTDuYmhaIYI0gqbXT8PDs08GNd1vBzeLgrpLE+kDqrEDOFLyn
4nn5MV5a+NKAHewAJB9KAnbzd98A/EfpFR/IvAyBEAschn4ymBVs1ghyW+CQEIDG
HSpikfBjous0j50jugBWcHEoC2Os/UtBIx1G9qCB8T21BH4exAer0ksPFxsUitub
ViedrgC8Szi/llpCJpNRHSxNrx9VxceKtOSzQrkLNCJSV9LUoG8NsR0m1CZaStoz
xN8DlQ1aiCuT8MD/34Ja0EzBgw/CYqHKXNLSjAGg/bsN/Og/Om8ix4XshaJ5ujGx
F/Kum4I+d/RgznRlf2VhgkaIdztA+VTI2wdOXq3nXmy53U6rXVTL4aXcr4gusvSQ
mVgHWpMigSYooX4F4RZyKCzCy9MMv9KZ0kGey9IUXxSVbTCjBl37QEMGDbW6TR9f
9wzctq9c5qROApJXDKArDe/YZej3h1bJ6avxXJ4qLBzTrV208mSHvfkxSwPb8lon
ljSmCbyIEu1bssfJsdCm+GeR1EBA7dVreZa0ZaiP3HpvWqSpwnaK1QAWGyR/BWy4
N50wp3ITuyJgADf6bASB0/d82Z63ys6U5MAQ29T1LHZWNuoohBq+2MiFW+ljXVp5
OL8qrFvG/9BYBN/wiOcK2gPAEbaf/iDtyLEBtp/Z08toIYf4L5HKpWdhYV8JNziV
tFSqDADQ++yI6YNZCf150pllOJtidZD/Yc3cHa++xUuAFvjFQuv9GQFxugy38hBH
UhwM7MW9jP7k5mexNfkL8um5I9tqnXj/bz+a8XmUstzznUF+ktQeEajW/nAWf9j3
QWtDITaRISftjzu7O2swq3G7haa5T5EhNBHVCoHx5rQKonGnQkANh1EMC83yLPWI
dPtrLqKPKJmxx97z8AAyr3t+iyDYKChHlB1cu1fL/vlC33DAF5sh0d6dP95qptMB
tn0hLOEznj5uD5jTscFbh3MCiimbJLg65tIf+ZxxLpv32rVyzdKRl2a/VnMSaWk4
11m6qkjNKPRj5QXu8H1dsbPt9k0793RqjYvWdeeArYN21610SKd/IOvmiMFlVYTA
ZdGv6jcS8+LHpwgy54nVHpkASRv6bIxh9n+TKLDZ5GwPaibUQcaW6V4mT7HSgNPF
tbAfw8Ret57dQtsQmqoJkUK7BtOq88H9Z2pYVIZSfCM01j5cNCtSt9e0ZSfOAnt6
wzbMuHQ66hsz6S6qb2hiQ3ABlLNMbfArGe7FAmfkfWveaDKdpikv0jqsYZ+UfxHp
ABlHJS6/s+KLhKuvv2LGpEVP4qMza0wtqfbVxoZ0wnNs093VIoi5+m/BAvrIuGD/
LsyepNiHWn4XCd/YqP32Ii7jbyH5ZadTlQpvEriEQuNLnKoSjIPoKqiigDQUW7Ww
BrdkMFNXUX30B/Gdm4Crleis0J2XwRyWdbgtqAhyqNLUg0kThqtmm6hwD30h+qRK
jQmHYhK/ask4nYK0IR7M92bC7laPmxqzqTraFAFFq+PUl9Ho4K3n0CaXL/705eg+
xS9ITDnlXYySvin83v+t/m75Y1+0Z+CUFWRS/CAucy3GZgOPCg6cpdf8QQqRvb/A
3ExUeX0Z6LDZSqObGe5VwfikzMXbucmCDEWCIazbBrmUigCeOUwNiMvzyu8h8Lvt
xflp/3JlIHx2KkKrj0beywdUg32JMC48StlFjMqnbZqflknWQhmTCyLGHBbwiXQ+
M5gxFdMRxnWMLjZv8j4PsHHnNp9akinK6bI8LUsVvaIU7w5XUh3HLdJrK3X2R5qA
VqdR5QzWYt5bFP2kVEcDBCc1gXhaW2yUl6hWyzfR4MckcFGKnjUlMF7aQkLEA0Ug
WbWMxTZKcQ/4RcIUPcbpmKUIr6VxhBGOJYx2J1boSng9dxf2RrH4neeNApx+SWeI
DWG3LEPLi4gTVyn4K1BushK6F83CeUF06Yg9681UduLgTRtALGCqO6LqDbMp7V7g
gNl/nf8smrjI2Wsk3HJvHTz0Tp1heSB9uxKpaWK/yF7YEYzrCuI1YD1u2diEO8eD
/9drmpHqQJRN98olL+Onsv4Y4AHNKeRHuwR4bPHPZFuU9T8dba2SfgIvL0ak36u9
AhBgtDfOBfhjuSbzBNXOFhkik2bXCnZvEbqfHD7HGXDeiH4mMinvNu/9XlFPwMyQ
czZR2HMW9kzUSiFyaE3wqB1Ub9xDBef6LMi3sova6UyYkE0Ms2PlnRqmEmANyDhh
3zjj7zex9Im62HRiVrWuHFrIaU4v9rvV+zeZGq0Bn4caZBEEqQGQ1dJjZo+XX8Hb
JGFELbhoHlRLRm7o8R+wRqj56rGOwJL8+sqYSe0ut3S+HWhbUgGA9XFG96h2h35V
ZKbuMLX/Ta+HkE8enYI7nGNcU5LvyEGACd6ofpckvRXAq0PUopEZAbs9GhvT0q0V
uZw9ZEcqoc5/k+pccibPGI6E+2urC7yklOi0sYIVG5ElCf4kAsWX5ZUvLGmZwiPE
2uNUIy9P7jDNXV0Eho4yzzKJTCZkjI3+jyyplv9S/QYpq4EdOGbseSYNBw9wd+QR
2RNABuA59mu5kLopblrK6WOWTNknPF7WUA+GZaw6x72hizWyL83gMqcaJFS1GLaN
Yely+8U+AAAMSZ6RKOIRi4YtX8BrAaMH3dHR4Jmc4ZsF44PCk1+QFo+0Lv6rinWu
LPi1yqe4mtpq9Bfvfi/5IC+QAm/AdJjgOSfjWapXfb8SRgq3xdxRBXayVgDkuEyR
FrZisVqNdTE6ieqaIlFvv26bKPDyNZY3beGqmeqlyKEzqwFT/rK+UyOKUX8S3aO1
5IYOY24GCeAI12dGvyEgk6ArezeE8ZhgLshBXabuj0i4+lDvanjA7CnKiYvRDq3N
49veB5bk72OHbCPKAx4gOQUtrEX6KfDgUfJtTKNP7TVcf/wb+VzFbAtf7m0AS2NC
NaEoObKV03kinjxhEL0RS9da45MUF5xhuzM4uGAEQQIN1/VJiwPIkWgvE/yDOArP
AAB6e7AjT3/xJI3F4LCM/qXn4rVhKx9cJnVfraITlEGE228yk2RN0Y07Jqq8yz1i
htr2pb3Nmqc8k3l3BKoKR1i6kHA2YGhSDP/w6R7f/7vutADvquvNwE04aiqbaLLH
GB9Hjo2WpJZGvaK48bPluRxRDeWyUSgmc5JMb45QBMNshhNK/NQJ+nDy+lUJNswK
9RaglWa9z2w+HK66jfKfdDvjEob82DQLmvfa/U8ExCqpUZcI1xKp6Y5Ti+B7e21U
YwZM4EAZ69tnRWhTXEF8yUOyNneJhq26hbfLTJz2FFmHRRlqgKrjNlVpvObgKphy
K3/RxLrl4XW30tUO7WUOPw3+f3CkedCwIpc1nUtIEPoGH/LoucXQ6hURKi3w7Uq0
c95L8Gzc5sF9iIuypgQaw69g4ryvC9+eCeYbj/Ly91SN80HfN7r73OUxt1r+qqyF
fJvcFnb5AU0Gu81ZRMy3jeXNxUD33Mkc5NL4CoSZF8xzWyU/3IzYjg0HwtNb8/Ac
cJU/7sKCrOpyIWY2x4GYxUBt5VrDIel867gmNixSNif9Xy+yqzAadpMOIyS7cG7s
8Hq8Gw+j1ZwVaRhVXPxzXSwyuykEfvEiKH8881rWCy7LXzCkdOcXcdGccU2cMmLj
LdEK6sVfqWlBFSdoUZY8SJUHz3gWVeRjXSkuCTllXBaUGF8e5UpwcAGpRiJzn/nH
A21BoHFVrjlCHz45D4rpHdhRLJrGqLjQeWPry5YuqHFqpxnoN8xDxgYKE2auC+lG
IBGq4uHdJ3XUE65dBCHiOcJky3jsso/kuRBQC3ihRNJd4V2di5w7m/AjpgYfF39a
geAf6byVLnCuutHLF/6sLKlu8kaFrWTCDLKKnW+0fFI0j5fZRqTAOikxddFjfKIo
0IVpxvTk27qKz5/CLaCvOBFprOnN/Z1AJeLoEKbX74pg+leKcTBNh48B9/v1xTb1
pAfX7hfRYm+P5Rui7Rai/EMZvrGWQeDDBL1/EfXmLHt/aNGCpFEEZHQcAIaVhC9S
tpMF8j7qm0AG0jTxuHduRJHkqvZD/OrxHlp8nGo1fid24TASQG3lce8pISCZlzsb
fI2bC7J0WbeLxPeFJ8+Ssew9O+pa4acD9/qpx0inyqLx00Luw2sUsBFn0J1E5iHe
nXZVsN6FvSW3gEIABDSN9FC+IJAH/SsioBETcQCmCKZiSfPUy2r1lx+WrTUOeC3s
ugmAHMIvNoR8Tcs6He4+Qm9rJovpFWvq5COloZyG9nCOoAJB5zMEegke5asoVlWB
QEtNsNJGmv8evuO8sDe4zHtMq6THCfCQ6uesnYNhP0lTPQfMiEL6aUZFhL2zHgWL
xP/fvD3mmTKlL65wgJEYkRY2zv9x5VSDeJ3zpZztGFKNI04NQ28ikUKCfvNw4+GP
JypS3E8T7HogrJMB7FxUuaD3ltwwSrQ9AsDTLw2yy8gG+5kP8VYm5iAIVWXanWor
QGqWKo26RLxUAqPk8BqRBd3+3UyEuq12OEx9IlfckCaEjqsfE1IWDurAWRmzJdLq
USD7ZkKUQOKiWvsxLa/lDdmWXcRprZDxfAgAQEQaqYuVgXupxmDDDZ+IzcEVlLng
2+Fa3azDb90GLDmM+jyHuYT6e97zIvik+Gwjm+fBVjWeBV8Eb8qsmILSE7WbVBIL
9ZfCaQz8tyFGQWbQ9EKg6Dm76Y5kM/jRodcjCNCEyJP9Qcv9ZZhG2XyC9dauwoAy
ioCT9qC8SeKldbuhOOQrd9+1dqclpzJTJ/ajON96h2MV5C9Z/+iYRxt98kVSmI2o
VkUvXQOEn7R7165ypIJIH7JDuKSeU3B68IG38gS/nYQXTIDtTr5y4S/JOqF4m3ro
Pfa1wXfvL5x35SFYe+AmCjHfLiR9sNPv4oNBneMp39oN89cQe9kEuTGItURBkcUQ
Yvzy/hMrIp5fsUKMeup0lkBCdQOeBMRKkiP2X3brr+3EuUs06g5LnHAi4X9Onrt+
PdkYFAL8Rpsn7P8VHKmrwX5HkkP/f+XvzQpkK4LvQaFfsc5uFSPmuiY95tPz/V9t
jXFmN6iR1E2jbGUa0PVB1UPYPtlca3qOeezQk6IoyJr/4JUMDm45lcdZvxozgUHp
fsvBCJJU6H0EegE9eXypRjvZe2hxK9QVY7zg0uHqJqiQYJBK5f43MaaQeEfev/1q
C0drYEj79siyArSWpskhutiPd7U4QjUvvS1SySgMjJuRW95p5uyHWZDukRs8sD8E
sGPDCaUPgMk8om2F+E3OqoCp54tUdZ44xm+OEXRufwCJ2CsgUXwGgUramq9gqXm/
WGUVmLuQY74YnoJ8uJzLqTDUSI8bTY6oq77k/QRO0VM8FfWIS9tdK7iUprXhrZQZ
SbjGFCXTl0bIEAxiJ3vQ+MmEd4fA7dgm9HNPEzpJtWvqVabdebSDlcyY63sHIr00
wpCPfRczbA2qIMrpuTZqDGaZeio8pIImiuBg8Ukz3jcFzz4OScXFt17sZl8sZfQP
M3XZsyextvlzjIKy3O/4suZAieY/dRlfuWWCGYx+/xUHfU2SiPg/KRb7ZQzEB5df
ODV6TeWVrusodtvhY/3a4gRhQuE6iqfL0KSHWcMzW1HDil2VhdNuLNl7y/0RaPuf
YDddCXJDKc7Urh89xl0mBVPHuaJ4BhvnV4ZIWLYPnQHGMaSxDNfR+37baeUMiCz5
58PUA5wtDYaSX5Mm5cUj+/24407yxQQyJ8QN7VIuv6sIaNPWNfbDSChwDpGVsFtb
igdy/49E/0TdKV6C+XTFgTSF9EjFfrlHaPkX6GUirBK7k/W7eZGG468a0DeGx8Dd
tSjFqxsRkmWWnhNMPxc1YAOh8sd5yma2PMWEEsWJAG+yT3n61BuAr8b34qsmBp7o
XbNzGK61NiUIgRHRZhmAzOyhal20bcFXpTq+wY6z/TkzIvet4g27xdIBV9pe0gHb
BqHjkBHOtCzEEm/258Wr9gfc3mFrMzRcuXKzs+Bcvv4UsRGWBCsZHzyWnPiuj4yu
t+VnxBV6ppzl1fHxdOs1ynyejgyoPQYFTJdTXT9mzq6LzYZe4L5O7ZcCI3kItNAO
PYd0hOuuaNGdJTk0zoTca8ueEmVCVwOTrl5TlH/CzWhNcoIyWE0oOle7JAbUSwNO
zQuDB4iW8ZJ6OPnmP0j68wLov4XI0/OuxRjENJ7RnQX0aMgCMlECBxXFRs8eer4i
Oj9zncKAL5K2V0GHSkR8kYgHmITHrmSN3XvLCVs3YDY0JMvxjoyaGfDO/YGnWTUF
Jgjj+1CIaElTqGbcjbwJo6TtuaSkMG8oSl/OKXgwM4CFDvsA3R26Jzvxg1tIBxij
3ruigNLJeq4WmUAws9vjPUjRGu7OkZpEEEiKwGfQ2p56uuubDsqPd+JDRujmz2iJ
8nGcw9gaopv1+H/9npPGirWIEP2fjomiYBXcMDtcsqmyK3qFxRmesgG9bTauflqn
lb/ZGMFFFF4dEJGiVauNpNKakihZBjcsERKhsxBJH9yBdZFCDBEad5W/tEWLsW0k
yE9p2eDE1L/j+ZDg4vfANw+xh0oZT2sjrWazTXze2AsKxJokRetG3qOlu2WBZrTw
ESOZJDuu6jUtFfd7+V2AkWRKiZRJu35yooqt8kM/nEU6J0jPzpYSR5fjGOOAGZzw
By3UmsJ6hUHqLdn2Nmcgnrc8gESQpAtjym35MfMPLumsybdoj+5ZNT1bDa6M3SIQ
OtTwbiUAK8vtbC3PEQG86VgJzZgkzrIF190l1ttLrG8EL4IONbx4HBT3I/KYNh6G
GmTiitBVejyU3/ALg2zn0riMPjtTACrfMG56j+3cNdFVoJbTXO09HiYEhjTN/TAS
c0sTUrL1ncQtJs16pIzJYDBI/QPMilaWEAkOC3CjSE7vvXcLh8fHmBF9r3z7i6x9
DP4uA7YQ1gq64xUNbEj9Ohk3YqnBvM3J8a5aYCQ22H1ObwTj4dKt3WohELeq93Yo
Ywtuxm9s1fXc9SAncpcLoH6X3vpsIybhOo+zrVoltpcyO8bOPnoEWrlnmtERmkVS
Jjogcgs4m3wGRog2OK8eQN534UFQjp5ZigHFaCQZKxuiLsWDBEUZijG83nbw4+t+
Npo8RkHO1SHOXDVDSE0PAvQUCuxAD6WO/FHb2CnvKflcVPaJtKreUzV35uq+BlBE
pUYAtnQcIyIfgkY3loD9tjbznIf5mOMAiyKjlcbI6tf20vOQaXQvOc7s8nG/xWSu
9m7ZyG4Wc5c3tfiZjj2HxG66oX1R03AHyuwfzajn/mEd+sq8E1Vfq/UTW18FtnM9
0qAZ9Ow0j3O6DS1l17J9aUkwzYIGanlyHPxL5bzrgoThv6SUWO5/u9hs/PsujZRP
mlOM2czB9OIuev7/MHDL98Bei4ukbZrEU+jUi1LUPRpvB/onxLkS524Y/6Uk/PKy
9iE5d5u2e7GEjnF9MKEgIQWC3AkKAMcR58XjwLt0nHOY3OTnVXSId9KaR2NpgLxX
tQxQX7ogZ9wMVmVtduPHjcAlcpLOq6i1dUmhQKEHYrCVk9dKwoj5lG0v09EbWmmT
KJA0eOB8Z3T9LMV8Ly6IHbMqEhfJQHL+jAqK+kqWx6r0HZBIO3cKfAjTYg9IMeN3
NFZKzTWoi7Q1MPrzpWUubRyzbql7umx8WHtVSEHMTJsSlPKvpeobcn2QnRZiBjXj
M4C/nNHUxEsfcRA7XWk/2klMjLNMXn0P05dCuqJJuaoVJ4r6zqJeCLdK2gcSC0zE
7xlJrJ2OxajZ9ApY2F5WzofTzJtq8xbclMtlaCfZNW1D1OumdmTq9Sa/Hu12c44S
h5Gm3YuUp5cExnxKUXcDldoPdBlByEHIDhJFXTLTnnkA01j95OZGChbCMTQxlWpc
QcOU6zUh1cQYaNyCOK8QWPdaJEuhG3RSruDAaxtLjt3mGTdNd/MST0le5P17cWxo
puTFoPKaS272od06aWo57+qfBeIUnEhMstG7nkkN/xStBvkXrITBRP0etBKJy66w
vQXwOWYy9eiS6GTiNwDvdVFcZJhN8N9J8uf1/OiokeR5p3PsZ1idqUqUuMfMWsUR
dpUfpss49yBZLHb+n8f+jYNIvrx8Mi4xbcNrn5Efami+leHeW/sjmf3Ty96Nvb6j
Tt5QMneQsAJPqlrfELqDFOYp29lu+tt8/rSKHOGdriR0Czy3NOmwLahQ1aCpngH4
E3VnJznQXh4OVKdZAFGDfYq9itZQq04+eDY+GTHwBFU1NXuerIE5xOgsjyX0wJSr
4j4iRyrJ9k0t1hHJnc0ZxQlyCrQAtEFTL2fBddQIwFBjgBV/L7or74J+OftjFE50
oftqBKeVI6KGFECFF54/cDNozp0uTo3qWPlIQMxc97kdPiGTQAZ0fPjt/f3+R144
nSzu1/CWciWSr9qg33mBbQxezZyOc630NEXuZ0L/jrc7PFx8QvRD5vKnoWKx8jZF
1HrSi51yme9b/SIVjWlzOqmJTS1CJ4ns/KqqliH73CVu2mEZKkyuULKkmWE2CTLs
Xw3UsZLyzJuy/VjpsdDmyS2AeKGcMxgBu4Zz7bReRRPy9n+eoimkWqxe2xiMUa4J
DKtYNq4rwTpB3yIyUEV0NmAb210OB4N1sMRdgh631ddwlrYAhft5L2TmyRxWP0Ab
Z4twthqNvUdHe7kPX3g1PQi9fJeCnzDT87qVDqjlDo7XkeH4ycE0zRjJV+Dlc5+U
aTwe4S7b9qGaTRhSb7XlOLRvfE9jXvNxH11F7eFvRLVriEzlRdiHc9vZnAqwGiKs
aTS/URQ2Xy2o5fTtQSirKE6FX2xnR5hr0flciu/STwKTINBuZJijYriyoJX48fk1
0/FhNtz4XG3SNDXHSBQdDXFgMyDZWDsnfxBQEaFIddchwco9U1mfU1P6KHJntR68
dnDC2e6CbCG7SWi49tN21hpUtM62AG0oaAHMv9G42F+o/ZsmQ8nGrOqeJ+uKY9pg
QPhsYIitlcZ3Oo5Fq6czrpAwfIVsrBwQ1FKRndPHUKJTx1DZNwki0FKURCgt0pC4
zJp0NyRdESB8Hde5Ka0BzK0ZytvuSflD7qNYXKQrG5PtAIUC6VuT/3K+OgJ1sPKM
ZDf8KdXaRJC+GzHP1i+Yz9ZunsIrOzjq9H49ua2iqIlfzRAuYerFuI1NypSmTiAM
drERqFHieIfieUDRjgMtV24fPHnY4cWHxFWCpiaWrTcxqN1wzTkUvMRtXmKvTsC/
5+QXK5wEmkCTed1rNtAaZD3CZe5X9I9+DFQOZ8XC62ZnYoYJObeugwc8WNeOeT6e
urYjg83k3dYcNR6d7j3RE5WrP1RK+nBQ+XAk7iI/XtzUHPRkI+hKQOIjwnQCxp30
eABv4K56G8r2tEJvKNFXCsFVEp7bSUXjaOQu0PiSMgmVjMOtoBOqgRpTSMBK4Rpc
Su5cg14VV5/xzMdRD/jrS7d8wjGY8wiQ5XrxsDebTnAIWsYCKwrWW1mUKgjf8mYz
RAtScDtGMe4tPjGG3/H/GqAyUFyeMtAUaz3Av0dMamC0lKA3Tw5X2p8e/Z1dOiIx
7MVYfOLTZDRzSV2sjKSW4ZRfqAgR5aN+LNAPHLkUtsq+DHDC0h9DKMM7+jHh2NZs
ilQfIp/iDinlwoSCcd4CtaYCL1l0Heujr0T+3sxHjRmFmpkKd2l1BxtPqrWaSLxA
7c/Z0RuzY/MiFRp06wUIcdnP3PGPGn3QbH3Nwmi/ZLPiOGEQ4ESHH8wU9mX2T5TX
Sf6xzmi7QRJ4ndrqKiId6W5TxzU8xEJUElXLyIOsNopPqBotqiIXzFx7sRbobDSp
wRSeR/309lNCnlO9Tt0Geypa/2/9c6dHtcDPG65NTCH/dOTEJhm2KITqCJ+VXH5r
E7ERld1dSPWnMvi6aaOVuv8utGmrV2zRvD32STIHLhX4HSJR+Y3R9qH0Q6WQomvW
f4/omgotvcb/xPLG/pzS6nQ9mJKyz2nuzZ+EiBv/ZVXgmQ8Dblj5S+qUMn3ebkVN
eiVAm5tfertESOU0v04j00xr2dfwkR3aFcxGKeWo6ktYsVnQQZT4lhCnrj1NCanD
mmbVxJ48vY9eDOCr+0jB4znX1UWmAu2CI8Xthc1/b0Q8xybt+6NEJHGKa92GJ0Ih
oaVRByQLl+5OKYNJcMz566vGESgHV4FpISoIoJaWBY2ZPbjXMe6tSCUmmc5koXLu
g3ZL9bw0dIL9/naE5J3h/Hv/E26b9Ra9zzWHXYHW5L19dou/ETkEBNghswl3WqW1
WCU0QOSz3cRHa3VCxCws0cSsa5RgmR1KrMWXs0iO02ZiHvoqo21rom4VO5Iy17HJ
ottgO9Yxg+M5UJ+kCIsJhVvtvgd4nR0SY/sELJRBehOnoMCm1M2kWGsj9iVgX6dL
E9ELY6Txrs6ZD0DKS9KYg8xmKc+Yg9SbCdM73wUgEHzZ3vvasWAnfqk/PkpzxLXj
82ySvh/5QYGygEp4aUkdzvXWiV0bc/lKwvX+nGBZqoyBOcH89w0I4gTl+/baPboH
h6Y3M7PYUkVGeYCFSVOScdDexwAF49am2/N7xF0+TIQR9ujtd8QrjG48f+uDQi7Z
eEcTsXciNpQqbcN9AaE1bJILXLHN891ftbF7g6YtwcTTG2tjxHhvigCD57JMUVig
J4pq6fnkajUhLy1GO86UFEXfD2yFC8M2Ga+mbyj1/2nx+ksqZJ43EAgPpcu94DRE
1O2jibKk2fs+cUv/vPYR/jQ4TV011LE7ikAk4Q6tVYjtz/dWsG0cFflqeVGFBOzb
znqonPdwIu9I+a3/HiXzgoki0ej09pcpl3RkvCIOQ5kMn/3zAUKhKGAfC0e50w33
XdQdKygDmPudQ2epVdqD6aSqbuRVUP84U/DiLqSiF5GdU7z5XH7u5zu6GMGWN7GP
6pwB96LZErPK1BD0PLRk7V7ulFN149C9OtvzoTIEqRi6VzZLAPCONXhsfS4yhjMU
ZFdehM+1HzevFFYgFtZsFaMah4BUiHm5g8/qC0GowxMVXyzG9LPGX3o8Uggvz5i4
uvzl2gFGKqOXhKFhTtx+Xs5lJk9KZb0G+XrlrUU8wS5gAyF8+3a6w9AiXMerTscu
dAtuLyA4lvEOXCuCLRBuhj+spE8GXjMNzA+dbDBwOMC46Ci6zWGgSBjujHNJh97m
EDRsPmAOXzRtLUxzPj1ZJSUuqOEB2tt/mCl3zXxOjhGOkkdDFEOic2Ecn08ZGYZc
XuBQ18YJI5CIg6e68cbxjgJP9cYr3n/rfdMOa3ufBviuzUNRziG9o0R3Vr9XeHID
FrDZlfMw9aUS7LxiG4GK8VI25ULUgVG4w+ypeg3rmCeZ9LyPIKafCnm6i2Q03vAe
inz0vaxpeSQKsNpRGjOwsU8GHjm1Pv1kfbBM/RyobjIjfhaCgu4J8D252nJhz2No
R8wKzLgPAUrRZanwyTEc+Q3UIVKkQ+TNKZrv1RVcRKf6MAjQ3re7t0piF4l7rHUb
YAOJIksQF2eQMprzd08ZccGfwq232s0S65NffjM3VJltUH7UR/At2wdvPIjPgKpA
zDCxJfBCiV91g3580YfhQedG1tjTDYduqNvwmACaiiavAeukwLjKI+NYxkg5a4AI
7bI5n/6C3zmEaOgVhrHJrUQtGIxYraDgbNnJSN2idRXtFzJzKqMAd84TzGDneQs5
AbuTYs2r95kIDChdH/LfgNuNXgkxbD2t+OpwHFKkSKqxxkI0LJLAkXLa2FYBzFWA
NlPmASenmJ6D/rmdTnE6XX2vyKOcnFbL824578zPQxDigwlMlRX9HgYMsXkppAe7
TNiE5ns8sh8QwFiaUwIDI/lfa5CKToK3gV6yrIzbUigH5UyGnyozjh0YaHlfiWnS
6jjMDwFc7A1MBhS5ghbKzHGZ42VQXmduE7LJYTHNTB/xwKpbqG0aSxzlJnxQiTTi
ZjQoFy5Nuq4aDfhqusMI+rK+pl8ME6NK+cyfA5Kber2HMFPPG5VZPBVDnqoFywrv
vjCOAjdsHbKCeKoa2TNu61Cqd0tjk30DnOKI1gJhnWmir1NHXNDkdztvMAFFXCpV
Nlp32hUIjT5ntN1gOoEuN1sI/rVKJXYTG56X2DXvdplXqZW7kO+KDFfrcz3DwbBV
bmnNw7t+g1O9y/++lbtlTcJzpJLeBNIdr1nEBk9sAqJUrU0L82iIl9HnIJKJ7ftO
0mdrHSkrtGGDoKcOJma2QfUpQNtefSA7CI2+vVbIIRBPzzIKjAJlWFNC6ulYMZYb
Sl7dzr/QS4j6ntxSGwiG7fIOIqjg0+EfbN920M7/4qRCvBDoavVzf79eotq8e8kA
RYGvqtzpsSBZ2jZcToMSW29QHn5kwP4epY1Z4LMlS414o8D3DJP1VkKAyV+csgsO
nxXDDoJ192VW7iTB13zMu7G6AbA8nBoaYt0Z2jxH+wu6ktCrAUMuM/Krpk8QH2hE
wrZUgdquVcY0xwoULi+EzNGrv9mKYMTd+4zUZAaQslV1RUxB/vZJGuKiktCJErgM
vP/4JE5qx+KxiuFZ5nwa4f8k35/CPGrAKaIZNKhjYPYRDCSM0rODBTC/r6mtZN0Z
vXum5gMc1cb7TWzhyg7Z/mxWgWF0wnVg41YLKjCl/nGNOqhru6vhRLIxWJzmrQb+
9OFe0/L2EMUzV3DX841yzfr27eXeFKS8n3OuCEJSeacpnZePBtW+woLROLUQwrVa
oGQJ0GbeGKqA1YlAwE2UhWdFKXfK2JW07J840lg7WbP6iNlxW9QtRnZC4RDvzIwV
OqUe1aQwAr61HNihPb3RZsYnLLpSRddU969iX9MtP1dizGNywgmXmQ/2N6pfV2zo
AzLCGeDO3Q6uIwHRRNinN395SUHTAoKVIle9BtJyH4BCiJ7tX7v6wnqZvzbk9AOZ
Tg6+mDELCgA4ByS/N5vV3Clx+6nUyfYy4MWDx5LHbMx5nffYxBK2BQAPgElH3aEP
MqIrwYS44CnBRAa1D+nkXUB7T7JJMfMuO1qW99j9cSEkeKpsxsS3CpDVhy5q85x1
AdRILBMA95rLQHujdPKMVRjd0mOos69Sh4HvgGVuW02LyTfs/p13JXq+RPxQ2dHk
sUuVIYi15KZQY5HhGy8LveCDip9SeAutunkm4BSa4YI5ZJaTV6gwQ/HyAN9gknkI
V+1PXBTknRyde0I5O3BwZF7sFyHOOnKu1gZomHGQg+ap1e5rR2+/s/SH0IH/uTaO
sHUUFAu03CILBYkJOax4PHEoY3NWliUATUc0nalhkeC44IU9IspWHlocVlWvU+ZE
Te+JNkrxBTk1jRRcajDosfiFtqXN5Pwxx3ASwNvB1JlHPearVWkqP/SVTobqpfWp
j7svkKtWYOB6HZw3P3ZSpI5w7YWuqCdBOQcnWkQKKdAbOgHe29GvfUtiIWx9edjE
fn3wULjN8ppLlMmU6gvlV4v5587SOrTYlkbtfx3lpyhDzN6OfKnNbPyV4EioaxHm
0ucuSsKz/l/fug9mS2UthGa+/njAn2JLRxYrzsgGYz0rs2YDzdotxl5XnI6vzrmT
4P39DBLK1GX/bjQbjpWdnXMLvZt8ZVkIqJdseqPdWDoSdMKVS2Uhc2fipcgoPmn8
wiPQKHCAZEH2PDUG4JSYltITnVDBWsYcpg0ilfwQuvzyNmZ+u1nWkEqdkLQhhpz0
qschKamRx+qjQtqyPSLWrLulnsadWXk8Q+M71nL3bqEH0M5wfDSSDV8m3Jw7ySvD
Ij0QaVGwq6Hi6Fq17bpP6UeGbQzXqZ5us2m0dp/ufNYb3TCKYyA6Sxc7h7MRWoks
zib7E1hUgPKD9MCj94zEBwY20GhSuy4wvwFsbDw1mF878Iw9czji7d1eDi5BCMqu
3J0vidsWkerZ9sz3IttNSZA+nzUoWFRuny2RUAIl+uUNpj/3ea1y2+OphbTfeNZ0
NK0H2NK/v7sRjpSdgZhm/m1hsoP/azAe17tgY3CyDKktsT9+l8QPprVysFjJLSQ2
P1GeruwceuaUd7CAZqTUzwiaffCf5diMihKHZsXjv15L0GaINjsY+cowA1HLG8uS
EHHiSB6jQ9+F00tt5z6ERk8x/aIurgpqybg4D5ZA0vNiwRd0eRgkxJCCWlQUCCsv
5UmmF+Snd1kcoNIO7DVE1wwLTMhV3ODC2vtk5vgo5DIdQ2VQikLJDIVIXh94lbcD
HbLWhI55qnuM2uafA02crLlIqsCN4IJBznaifq5knAVcbOq2VSzwxqF5fZXAr69b
M/ChVQRss0CqkdLsHDBDl/9priEer9SUrhnlJp1JD1jR5CRRHgFlpUjkFk38t3b3
7AVUyPM/JcZPV6PLVqWkRZeyLuGX+ZztGlouiPS4zHiTYWVDVPBn+znm7bHfm3TL
236CggPgU5juFRMrZPKYlwlX+Dj6w/lsx1FtFFdqAGlIV++nwIRiAFZz5N4QWurb
6cPvAd70Buy+NWo9y22AXjyUMLgfJUg3aJF7kILM8c9GajAexY98IsjBF+M8jpRM
Zx37DBYTO7fo0cnrU+sXS1bQxRBfB89WAm/KDVvenNB2FYGg/LYFKFElYyKJqV1D
PBnMdijH762n75uQQR7iq7Gjn3OLL9WFFXDMvrgdF7Oh+yKBePW9SkjC71hSuqwM
jSFIT9kSxo0h4ynNPKL2r9PNi3PRn0Bv0cvrwVDCnukqdSEvEsgZciUp1pVvENvi
NcPMJnlsVKFScHYaJO2tgnwhXnbKUxGf9nSI2ub6/RVmCfeIrJRTXsJsEn6T5UTo
m4SMA7o8sGoQsLXfVIOJJp+sBTHpPctfyelVRCbn5S5zG1KofQWlkrPkoYUfspNT
DxF/Az/5exo33Jrb0r2/9ZJIo3F8ZFeWcwtE7kgoxWhXnay88Nh6r3Xakh7DiSKV
DRsWkOrWMBMAwJGXAVdRXTNBgr1K25f+u/Z3ibSbWg9ef3nsQsQMHopAB0rDcrBl
FLWnje95pay/ZUc7FmjCt4ZATr2/4G/7wNWNas2RGq0XLiaJ19eXnyq13UsnWrCc
SEMuZs0ey3vZXRCycEJWFRg+11Ie58dq+oA5+xDj7meVUiv7gNcE2scwUvbipMh5
ERmQADpAsAUlY8OYX0TDV0on0Z44C9nLRhTmijdbKRB+RZ2oCBHu+gTEuJQ1efta
U4W3Bx3kxH6n3Dsn9OiM9KsnYWdsrptSSbq4w5KhfwVk+OCf210SNBnEzfGN9sSL
zN7rJRuJcphDNDqxUA7EunjFAzZJsqPwW9Rd1+qFqlrl3gfVsY8wW33qqVHe0wlA
H5ha0xjZA4ZYHQKbATmpO76uASpJMxY2/mNpLCc5CYAEc0lUylqw1B3j9OLnoz5d
iSKAxRZs2ffeemOD623ssHG3GDZvnKQ7Ct5O0LJS86tbys1ZwcJhwxz4lv55fhAZ
/TOwfgdexq3xpZDlv65nRa398YIKO6zGlyXuo8yHoefiomcObg+Gd573uM8IpnUD
4miWEFFFLMGU3CIfwdA9AfR82+Bc9XFrhlRsVJo6quEqrU2DOhQ/C85/TF5gu7Fv
VNtKx1+lYUr/hXSMutUx4gXtIFKObNF7tCedNhTMnIV9sQ7QGmxeylx/39omNIWT
JchUIdkA3AuoGPMbnNmqNcy/VPOy1IYPFniqoUMcysXZeJIZrqVRK+7/u4N93W4D
omNHpiaGbzdZeXsVBrb6H6EelghGfAcoBjqHOPx2WQlBk2WCVuITg+41zNYQfmkd
tcReQXNdd6d+/o+2C7VZfhpIMxrZlUSq5PCgWMj/pkCZiTOYGzLwR258w08ojUK9
5vjoW0madX48aCvFm1tvKhDtn2wwT5Lpx6a32YV/90hEzhQgiOQzeqn+hGtZgPcT
Vg1OzLf1bQmpYeSMjRpViYFf0+deQlNlAEovJnE4qVpKh1Qkxkl3Anc4TaSwyV5O
S4ZcY6JUNTc9MJs04Zih70Kgb+XlEXGe7uR9NGbJwU4dgfIxyH7tex7Y+hJqxI8o
nh+FmfcOvR/nqjZ/5XuKGjoWis9HRW85DtQ8K1e7S7Hp781Agq4YkXVKuF6eDQlH
ekz8nRZW2JMKoFsh17DLHiWt7tpqmRyu7e52yLLWBWsxEdxetbTREEsJi20DBC/y
UbW+z6WPOX6W+KUr3YIDdupxhUGx21UupnlG/IwN6m4EGzQF0TRFgPHvU0/+GJFA
`pragma protect end_protected
