// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:25 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CvVP9HYJYxj9gMVaU84L+1FJzJnOsGKwp58Mb+RY0p+MO8ViPC7zDUOILhuMz/YC
3EIWp92mBYz/1oRYQ0abTbKQo+wvL5xXh4UeoYw8n7FlYeCWogQFu+7N8z+OHOjM
gjZGHWEwxnXNnWdFj17w2sP+nXzs/SYpZnSLv5c/wgE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12432)
DmiPrAtKEUEGsqrfGDn42gfcG9I1uKkk/oL1vyUY+uByEhBFaT+2fToaK8NPYMCw
xJUOrAC919r8c2oSbjndwMaIMpGdT5WzAIQkNse3j6mwimUlScisxQnvJ1veE2Fa
75Mfhz1G9NLymaDld9C1znz39Mei9t082mPEkcmP0Hw/cBlaadE3V/4Q4voTUm0J
aEFWFwEVSZISjvAdPuaGVvS6Sz27pV27038h3rOikI/f7kiCsHlyLGmv0zAoubJG
84C7fqaJqjUrVCU9qIF/NN+3LzsObqu71zaiQXYQE9m66hY2SUVDpasfhpBHerkg
MdiyR7sYPTjq+YAUh1AjF8MyfuD44SSisLJ8da+x3hTtXakc0fjs4lDvrkpSc+Jl
EpGhSCsupUATiCLiMiJVseKoD2bmJ9jU2XmDBU4nbTQhNuZX3Ppr1rpWmoVrwtRo
DL/Or1SMcoiSV74viV/2XA2dF1Wfdw5RgTEKTnqS3Dw6A+HsxVGjljIZsHhQNX0A
1L8f9srwDuJRgVkxKUJq9HVqxl10guOxYYc9RHJaazAGVnF89O1JC1z8OSszSx7D
fFDu8+dculb+2wUOsW8FFjg7UMGQ1NGgetKuNqcw2/7756vhbZQnVc1Un2N4QvgU
i8+t4nzr8unpmTkajcUMNT744AQ6g7UjsQQnPdaaOP39GbcNzuCqE9Y9/7i6AvIU
5CJQ3LwqZqA7FD2/5TFoMOVKjFsOHdcSGTbbQelAQ44x7eJX5KT0OkfP+HqTYTml
ZfZdjFB7LIZEXyzQaXmSL0m5M74chOHgxhvHcKG7rLIRQ80j/eW/epOOVTPY1Iji
I756ZxmhHuKr06Zs5dkPZchfDgK8imQZqEFD2VDf4gD5S+FDHb+21tSyGspyKBT8
Suk08ZBErxTl7sD98/hvG7cHyJAgrmqxfMuFFcjc5R/Fpvg/lKRTLGp8jzqvWG1c
AF0c9Jz3pNlUM4AHFZS0tO05VivD++pkvAajUjk67lNTp++1fK86RVqxYQZ03mOS
7ZE4c3wn7/zIv09nW4tl3i37JSD0zd7tt/rY467jiwjsGqDLXDRl1XQyEVpX4+Pn
2d9RmIbR2okO49xqp1wUtdpDwYcP75qtLrKogE8it5fJQ8FDtjbB+3ZZfClL5fCC
1L2WAVqM/pOftIiupSpzsmOadlJcAc+z8o+m96dnKd4/sAc4ToEj1Qm65nuyop4i
6tFhJGQoPzYV0QWrbtX3qOiCkcEKzji7Pw5hAeJmCTEjB7V4Fw/9uJFV1ROIH4Od
x2bFMIwGL/BD/2JIWOGStml/69LOMPPqb0KTKA+0k60/JxgbBLlYfBnnWgkhawjh
cUJk89lWAu0vzoqHnB+F4P1kSKcezRRKojxp0eNiP48j9xYNGhjODOT1H/JcwvoT
g3cnKxSDEP8lbbIlRLHLRj2V/NJyj6rS1Nf1BAzbwizb82AnFy416W9ExotsC7PX
7vGQFgxKdidtSHvu4tFj6N9qiTljpSjvpOdHhXEAtZwPlsM0Hpz2C8WmqpA5v/Qt
e4w1EqI89NhJEhwWNgyA+5He94UGBc71B/rqakwhUWh6c3UBSmIn1WkCgt5HHZTE
wNuek5W5ZrNgRGlZia3I0943a01ym0YUpN7ozT4qpaRab5hIMYJh3e0lAaXelZEG
i2nT+yu2hM9CU7Wkt//GLH7cwfZkSIjc1Bdcwibj2JVjqmFCMRVO65kN8BCoxI8V
PKEq2Jnp32snZUTSjChNCA4cMjmbVg+K0iaaYTP4kcarMGRBjSdz+e8BxEwEykaF
ABwFcgJyyhG+zAJhwLPs5X7+lQYqanb6TRvSqf2690H9HMcsNccVXGGsPykCnUiv
v7is2EWswIdcdHBqpyil3T2nS7yXjqu3TBfcZZBZW49xo4xUpnJuECVipzEuCZTa
M4N3MqchB8gLoSO2vmazcMG4EFSMUL+Lmiva303HPvmAVbS1PPFVu9TqOD6OBjPX
9QY2hJKjnZWel2zZJZRAeZEFWo9ylHiTbUXVL4yGcTbYxAODM6k/AcyYebcT1Xvj
ZRiqPizXYpEWzguEA0ba1KSHq6tJRdkxXjaCtTQxPwZrHe8wWXQW5wtvJom+ns+t
D1x6C1CuyHqbDqapyUOe3VJ6bLn8EsDqnjbH+n9HIf4NQ9kM9rWgjexp6SaCzdS/
1PFco9Ds/jUDLXKvCt0liVENgaqniW+8bW1MPrSp80RIanlMZNhg5E1CRDrvkLLB
qlkvHGja2wQLkwcfLsDLfbDkZjYE4kxBdqMuB/whMjsOg999tOGgaBOlaIZF6YhW
B+GvdreuZPVhZ0RbswD7YigAoP6uE29Vn0wdFFoGt18YBaY+wx6ybwEHTqXKzusH
oCGuJc8cZAtE5vmQc+1/kHYrFXjH57my+Ynndl80ZgVPr1lFcM49ennCR8fhLdqJ
aDpewsY1JbEYxulkqX5Bc1N0C5IbhJVpTU8ZNGu8J12o0woJNmOgBCorLT3PfwO/
6xGbTzpCZdtJ/8NjdEbA5OxfaAIc+nzGCpzLF4UklbxF4tXWXXOR4E9CSRdjBCf5
AnOymMW0p2HtghJ0XT8orITbiOa6VNcVjbT4LUYTOzZINMAL7EAasYuQQ5T9L1zK
vAs5p3SFZ/AiljqOEKUSxIT1dPMSBCvvQVDAwYUKmREHcXhe+DTB5XB42B8zBswF
WzA5+KAQ0v93xeMEwo/MpJ9HcYFc0WpRXUeWC0D6eZnqvnyFkIAhEbMWAMmGHuRa
d1miqPIHe9BXDSahaWiRkPuDvVl85fcvrdP6/m7pnmw4umoM2vK3wel80TTY8wUo
k99lDGpMmlfzjXpWF2OJXZO9zac10p1VPOWEEMgKCTh5XbtL3mVI9nlxNVnwX6sE
jJP038D/pWnKoqg21mjse3GEuxFvz3NyQOOQoZxx12BVcdpEdBIccCmr6UCZVmfi
mIq9n2LHz1naFAFS/Z5boD05Nw2jMkTIIdb44khMFqNhdwRO8vzginoGiY56kYhE
SLElJwfc2CyxEjY6W6MxEyAnAOJ92M93vpwFlR2vPvCiIMIhl1TeYYy4XLmVYZzu
tk0lNlbgmTIcyteXH6qLPOpH2u8pOCVt0uskx9W8Lq5ifi4iXOjK694RAv2o+Rc0
bK2Eo7+I/2H7poC7Ze0AziZ+8QbbOS0K8YZpu2w9nvhQAVWUE3cBPOQgIgX4I3y7
atdVQD9XGJIBBEiVbVfY+AbPOYjhqEF44RZzP3oRA4+FLv5b/fEXvsnkQcbW95BU
JXFtJc3DFiGEzIxxB31mQQfYcVYMuI944pZrquG5lWHeNkCHUVP9vAezQjaY0iaM
b8NYgAsjOOKQvcnXHoQ8hSlxbXidb8YzF0+cxR+B4MwwP08Gqvxi08FO1PlcN75Y
OxersgTT2pIejENYwjmtaTdYuiOgMQhuL6v5LpD39fxAsMuAWbKbaBfVDSyULpWL
XfGUFLOGjbdC4PXDVZxnqi9PV2pG/cc0x/oEe99Ce9J89ZyT5man9DKmnKk3pmkt
4TAw8nwra7olV5QysQ4BRUXErdLlZmaE41+b+incS+rGccSOoFfw94T5oug34N/L
wggmNhhAUzh1X4yr1D2b/nbgXQfPFnNHu8Clbupx64SV8UPfPFXz9/Sc7p3RC4+4
mMnnZpH1S+/l9hIStEcxzK3gyZpI7BZUQ54qERv1z+gHHsGqBKA9GjD4SujE2wUs
td2B+QImoNNMckonbzXvcDmvf7U7zP+eDVS+QWNRzzfI7gL5+84toeHhgoGgciOB
scAlykM5L/PMhPmfSJkqm57grWOWkzvtkQIzrwNzYRz7pZ2SpW/dlQUrpdh1pUhg
t8PF66Td+W0Vztm8a3b1fvhbPvEEQIni7CNJSvy2MzBCM1xlP9qDXwcFie4saRKj
tr/ocKcTicopbTfGCaLKA+XoPfLH/mqZ5bfSHYnn0kqT5QqCxJY/W3SJEi84yTry
YFC13hLK/iCUtTXouxBEuU8R8F+a5FedDDQDSOH/qvXcscNTeGnjJKBXZjH6jPAl
Ywexe3K9GJTZFoiMuXFEfGTWxs4TmHn6UaXrG76AwU9zcuDzoFbi6J1dIVKemR8K
w7iklufJaW98E9KONH71dErAn+LqA2MvOUi98nn2+IdWtLvel1b0Rwqd049hsGzR
PpDTNRReSD/SGwPJzTmoEVXghXzwrfhp273cwKkSxqiIgR3M+A48UfL0SzIT61qd
jTJUUy8BxJJOUgtNo466WKGvGSm6X6R8c2GVrYyHOjxarELcEI0gcnDAXxYoH7Nv
TPl80gLYS5VQdnisO1F6eRFrSo10WkIsySTheNPt/yOF/4akAR9HQs8LGJymEVSW
DC21AWa4vlmOTt3O+SxV8x469AWdocFOIGFPZqin3NJtVCi2yfE5mUjbcORBEbcn
BxNAYiOScl8y06nSrtsMaPzCkSn76c4mdKngkt+HoNlvFcrY6zSJs1RaT7ZG6ZlP
hbtpf7r7Jt+p07WodtnW6up6LCT8PDAeobAiTGghvNT0KiSG2w78iic9UvR7AL0o
8eYyQyM2qj1KJELwKrziqNKNFNLYo2uvP0QfkCC3g77ASzgR7hCt2c/1NAji84wQ
Wi8ubLcyGWMUP4PdEk3KgBYl56iKhp38YDev57yAlhtJIh5BFKId6eUp2+Kck46t
Q84XDRJv+Ie4JYzhLeEjgxkEHDkMWD4VR+hpvF683I6R4vM2SrMRrXelHaLQ2Nxl
aa0R5yhMQ0tJMV701ehl+c0LTc2fLK2trDSoLKB5FAaiDiz78oaAmaijutj4WoQX
SSx/y+s51hH3spvDZZFEBsStqKlLnk2b/0QsZQ/PLRYT+hqCLHB8AsTb7a5UYqYL
+y+X+6HgUJ+hUY1lVxLyb4peIp4Yb2I83ENwaABPLVIwXRFXoD4Mq4TEjI1Hlc/v
7qBplpeeOoCxU4xzqGH4+HhGJ+tM2zVipK2qjOBEwp4GDqNKlLL3oSLnPFOBHrxO
W5VsmRM9JVtH+Lq+6uMFN5O5Hbem+WQ00DuwXZLFuawVtQ7FBU+zyXW3lEUUoFST
s/KV4Ix4hzNahaWjoEaB+S3girrqLjDyhAHsl8ZuyB1bC0HWjpw5bmIPVPuKjqL7
Tv7CVfUyg/Dz3ZxXhsmikqst0IJAH0sX6L/2sekCDfDUHP6THwzY0GW8htyWycxx
18EwcCOS6u+pY0A82ggU9aFCYNqNejXoqLjcqCZPJVJZPDqx6sLQ5cPo0xDdHItl
9X8mkIDBQg/LqMZznIB6SuV7cyZi2UxVlIHfGqOSnQWXu0wpnTtzNEMEn4tXmdS7
7D3UOtQ5dAEbe4+zE8aL54mk9CIjY+G0OnMIKqPFY1af/4Pg7tRSWBRN1KeygQTE
Zu+ddD49HQl9QX6FUniBwdlC/E+E+chO1VwudAikAjpza2Jza90Zw5XGVt5A7828
EPOVtHGRIwFe1URVi9Q6zDIPH3Bph5pVf/eJC2DyAaE32feYATqIqZqD/U//ofaO
eZ9bdGeJrAIGTzPlk4ersmdR9uzLm7BeqWvV1zPQbSFPBEaUDi4Arno22rz8kKKB
/yvWQGilISUe/fZtudN6YJlZbwY3DTreHlLkEv6PSNdyYjV8bldz3B9M8Lzt6eDh
9BkDgoYBAEbiI1TS5QXN2fZvOymzMUljCHbfthjvDLciPK/Pt9AKJktldrNHn2Dh
jfFQL1UAxTECTxHk+ZGgYrDXMfWYh0MrtPQuaWKFjfGJ5JJKB00AzV/+w6nRbi4/
NGxKs4dKlMZyGWPzNFjk6tQCEUag1O//cOnw3VAVCtp0WJWuP1F3HVsGOxoM2W1d
9vXkn4UnfvdUNq5RDLy7Kan+uIXLF5Pf/ZcL3n+H+5oZx1fDUdrtcY72FhrzSXkG
qlEINyN6dpUG7hoosmFh5U28+eeghNXmODMFGqUfDZI3qW2MS7/dzMEAJvQpWJhx
A2ff8tHXyJpP6u71UPDTkDK60q33cUvP1oXtbsWQ37Wg/Jeff5E5qSX7Yquxvnjq
IFwTL15aEH9Vvmif2MU3c/yaCVr9O43/Kpb2rnZSqKT/JA8fopDVukTH5YiwWPQR
+ZjLFuND2LWlspZ7c0sOaDwl8G72+Q2FNPXtLULFMXt7w3M+CtExFgdQbKYN+ZpC
YS/IsU/SR/fGOVmiqXdtrHm0kQmcF9DyZn/W/1YCHbNfs8KqMiUBg67WJYY4CQjy
FCC05namk8gW8n8+GVUSWsUc7MfQTuMq0xuW2ku4Cqn4JZ+nqw4tc8ngavVdRug+
uDJZ1MzpQ+BwF8sV0G7QJUzW/6d373uv4hxTBR/iH0I+qbOdgCDL+raIvqzuuYNB
tpS1g8O7xGRJ9iyiboRHhj5/SypF7w2Kt6siPg6VBuUyrXuzivpUgSIRRVPz767w
Ww8HAdAQpVnrdimFqjQj/3/6IVu4bn7wBj7w4kVDZbYt2sQLTf7efwYXFxT3IYj+
JEaJfU4Ks2OvcwnDjjNulfcXwlw8uOHNmxHiFM5Ml9HEvts70khSaTa7I3qgrPqh
/bs+IB6a257BtqG/wWqTb99/qLNyHlJzPl7c1LZEZxvdaxDgwyxGe6AgMZQBOlNA
uFA92wnaVJWdIDVy6gRcTnVAUlP5BoQsfxWeAMwDhBIzUZq02y0DmPX+2joTplYf
99piVR8CF/NRudlNY5z40diCMe0yLRySCsnWWv1uLvs968T/mlc7rokbuXGRYJON
Exr16X7B0+vtNW/eonu464O6KHJwGa/s7w95l+2yrmGJwSexqVelZIwZ8Sg0NwyH
9FzxpbeIqI/CKJRqhqEjBY7ZeHakvYafJXgrXg55zvLkVYbL4kyqbkHQ1d+5REa5
jJ4eOsdXjT9H+I4em426QNsHdug6vQJL8RoxVQr5rvMaKR+Q39qOubPhmiwwzDtc
PXnOoo+B7A7x4GfJwSmN0uQgbd4Xut9l5xENHdy4ynUfwqCSWuhUiY0euq9xXa6w
A8YBuPWdlM312lghMagGjyksKfKymRxg2KOS/OWdslniUCkbuwp6Z3e7s0jI+W/9
EkR6DCGxXffsKRk4bKSoUy+2WsFh2RxkA9+LsHXuE2gUaAqfbwf1EhZ3TiPQc69m
8MqjiQHKE6AzpAzipPTl09Px9sBRPGWIcbs/gLCBjvFdeeZzdssLn3dRzgHrojCL
OJSZpz1yO5N1Ui3KK8KQaZ2+r5f3g/1HMmDmc95845VQhilIhZgT26I3E1/4kxn4
czo5Ma85ObqnyVSdFReuFpLmIqfxd9cPl8WefxFvnFVEmfL+r5hMVl80FgRZC7+G
6BURmYcKTuuF70Lktpb9xRO+RScEH4yrZ9v9aLFJCLO/JG6O+ngVrt9dfk/s3lqs
GTmY+/utSaqed1eCGs9K0BX3UcOXVAMA3CHDOxP5ar+nn34LYynaXh0t4zyW9K1m
BDiRsq39lAYk0NYrM6bb6zZlZ1ieBl+aE3kv2qOQz8h91LXhVLfPoSBPR98Z5Slx
VjZn6mfU585VnEw4Y0pYeem1Z7Uhu4QyN6q38YTFCYDyXnTFXpNN/44YOTId9IjN
qMBt0d/KIZCrTRGgTWOA0+CA5hO5QJ+tNhxCfoLwgeWTjLOMXeHyA40UrVVfXMNx
TIvMAEzpcJqXmpQKJWzJHEp9hAsufydN8+/co1Yip0kJ/5ewIAy5WFZQvFkXhWuM
CCht4+hxnG/5KMb/vEZTU/TIy5CWbuDBM3ZYY3AosiSh4CKKnvWAYBQQDQ6Zltpt
guszlimjnk/gH2RQtCkqOnllnbxgySF6dPI+RXyuqo9EZNflXkUMa4cxSwd3I3rd
dKE71neETnGjkrXuIIFTfRxxo8geF68C5FfxMpZ3K0wy6G8p6bHzSacSGEDB87tU
oQ5OF+OWJKMGRbhjkSJTffzeteIDnofFQUABUPoUk9ppU33Zjr6UUDY0OnsCTQgr
6MWec+/0j726eR1hMPz4oxA9dgLiSPNH8qvErTMwzZWYD3eiaeV1AImkfI56cHEV
YLm5k4Cvc2bW1uXJJZt3tevSkp9oY8x6a+WCURhzPCZCUSXPpzV5uZOVSS1lbxeA
cHQOD4CBSxQtD92zrFbChzEU7wWQehqC1MBoeHh24l1KlxZDrRGfw7tYHg+Mde/x
mnxMmhlh2C2ew5hCP7J5JUzBsMsUJ1p4yRV3bKudXP1TqisHENatpS4vDgX+MFvP
TEzxgI+blbrE3B/DXIxNkAQD1Wv01YeXtFi2uAx/tF7Ldu9aOesS6/JS/4FwQDL3
5qn0x77O2ZUkAge70l00/VDF/2BM/T8pqsPTa4Vpd/zh0NWKli1KN+lPDmRtVz+h
JnwS8fKKqg2ktUaD2HU5/6H6JIxtirthzyl8KDNzI9/EcNyIXLgT8XXGXOEyYK/2
CVfVbNTEKlQaiKyioHPwV3W/AiJOSDMacEBRHYCR4Np71MGTfHbN2o1DWaP5Sf66
VEwXvQTUw3Jw+RmWXRSvZg8lNvgDvIXhTIOozm3mbqV1Zxc22LId28vuThsGf1dl
ShNH4VKFstfrJRmjI8ROZa3EhBM6UezTt9fKKLKNOE3y3LkEewO88+UNEaJzSJba
tdgGfwD57WEAkvHOgWWIG//GQWRRCUqsoYVPZfUU2wumFFUHl39QRZzUqCSkcxNi
PTSaHQ51iebBAKI+JfS+6TaLE+gNiJW7k+K3+5K3hugmaIwWEGmXk4Uw8lxgPLpp
SYkOjr1YWHR0iRCYljhAcjtso68ASbAN2evbVQ91Jnb7krPVUBJNiCpXPIP3W0D+
SSXdoa1WqcoJLGM0ifZKEl6NwPkv+nyO3o8zDYpO7GSRpNaJfIHHeVLgy1r/LJuW
1IUOT5TJvklhTgQBKB0eUTI/U7IuWufn+6DYwyEtoQsKX5ZFXvuRVOhEdpt+nHeO
FJbDLkyCGECxooL+WnLiywp64wmctt6dfYzNO8jcszVjrfWDTwDSVkQLbAwF/Sbs
whrJo39Dbpyb+P8oh5vXyayvhoErD4uFKSDWj8vxU9TbQSy+OjnLStdWcq6cVpjO
Hd/DENAaOqzoPyJdPZAwmgS9IFXRoUzXZjaSfq8qHVOUzU1QSiiwkmMx3bR2NmiY
w67chp7DLHQwcebmPRAyRvcz5CoVnW21lu7WNxI8KspPF51AA2qWo/X4+MpK1B3D
KaTOBzJ5n/+V5aNZakkAjVS/ESEnTDBm6i4cE4pbikPertKz9WUtsz2NZhyuSIi3
1ntOHL4WA91c6F2l6jHoaEeug33/P0XC5GXdR9frlvkPQ9CNtJzUer9uqSOv+m0O
kyLEXctsmPtt7IoWJX7/fuzDFgBqHEzk3CRbU1pvrsdCXSPYoZelokei2Eo2Rkdn
KL0e972MFLAMCLuNzh1QyRRzkG7OJFT0jm1mBUx+fJaMh61YYfxYpZeIsP+9iKRs
o62hdKeOgtacW99Xydv991yp6CoEhBuGICYz3B+Lgn94o723hmWt4F4KXlxHk8qG
jcazKJLB+OxsFw/3YA8g5o+S2FK/4Eu3/vsYb8sFYq5Rlpe4qqBi7upKVxS4IQJN
mHvHCWy2bLRpYfUpJ/J6Bi26jNmE74Ke2LPBNzGzJgI71sy5FPZVeZ69UZf894ek
1YvPh6A3VqaWmww+VrhvdcQqQIMyIJwZ4ftxArPNOBvmiKR2HxijUynSnYRbYNfF
wgHrYaJK98by8Zoujm+VcJ/dl54PQcjWnR8XLCOFWmJ9xe/7HMTuOn5eE+7CiAzH
RnQwXhbMZ5LjcUuv2pRNn4QhKwAZiYcaSihEXpXqQYOl0CyVf9/kY82fUVGB84eQ
3sDi8Kx2W+6aEbtc75kN+VQodWUhLkpYHcSFSN7sk94TIYpzz/VfQKNe/YFGOhFd
Pmm/g49ESINcXeM8OOdC5sUeWgkyc6hjWJSp8t5ZfuJzDClmOLrP+Jj2eS5MYiDB
n0sC91A3LycmlQJAZrK93AIveitJP0L+IbApoWfV083Qo0fzL0xENDJMKRWcHGuH
QI00TidtDJgR7DrtQphohmfGtusjp1ov2AiObTvYFjDMDapMnd2BZXH0P0arwJ+2
pES4B4FXx5Vnc178DOdncDHk40PzwlpF0YBuqisjY/5wg6M1drb/WNQF+YtgSws/
mwrxd2KGJp+zgf53Od5le3bNldvzT4LOxgF+Ob6xVEFQvmdke/grEmlum4E1M6Fm
Nsm9KXWm3ra30tmWa3Pawf0PjMGeZq868Lh0KJcmHI3z9N5mowOTdJIleJPfKsR0
W59FiKYyKCNKHWvNr6RXAlKM+UzEr2d+1fiY7GGXcSMcyWzKIvvmQJzniXLBkSdG
CcxL6l/NRL67MOVNM/ZMZMPr+pp+vlz74bBPTE5+jmcD3b7YtZySaExokAvpRl7n
SFQlqrob4Zsj3nhdpd/1m8fbZa7K+F8fKTfPzytbweoASRRsbAgpnRh/dKfCOEyJ
bphtTbJB3cQmLQ8ia2hPWvI4i0fzi16SloqwkwVeJjvogiKX/MAmK3cmb8vavb+d
EdBeheh6iNwLbXn+8GQdLeouL306vRSLRDXo6CN9wbPUJLsxGDm95/hxeeMksind
nWfqAq1zRotm5yplPT3DbCI89U1+VV8455IDhbYGZlhsMEpOLnpmub3hxxZxuixa
4SSfjHBnZTQ3NPb4KiQnuMAIReqmSXpuE1jQBpoq+3CcjafDw7VWUEqbMnfo9uqo
3ZZu5LEWs0OHv/JYaIlz7Ja3jm3ey3Zcm7AR50FRjqAKr2GVAMfgco/PzTt9Rh2N
3uRg2cC9842jDxCRF0Vb37uaVrBbduaPMr25jZWfePUQkqKe8gnogdn0J0bVJk2/
17BkIkVnsOZvO8bZmogXs9szQIk8n6Puhx3XCSTxB1QD1oHA32g4KCYhKEKB7TWO
CHMW6hY95OtqLAfinwXyHAO77/YGsry3kUsxPNfuFnwhKrsJqfcqPrkptkcNS1g2
NwHsbH4x2yX/cn4dfRcTZG91w9BxltrzNsNfhfAnjMStvcwuNx82FvVctPjUlQFo
1UHTaA1khC41v7HlRgvJDpOujRR0dw8ewH1JlW5cp/jif+OfuNxpa40JM/ykrX+m
+KAFWkEZcHXkjrG5EwNpwer7Gc5fi5BUadH7J+1S/gt3US1xc+YYYBCgUqLRpCfo
DE8ErWJVNaPKnaDyiQaygi4wvnB3VAEt517p6+VCIgpFBJaLkxmEner+9cm8ubhM
X1ESWR1dPIQx4QB4bamUcp37El5q06DGbrOILfQRldbzaTdWzZQGpPnh8gHa4wjZ
qkiIu+Bk7bBwkSXX/EsNucWeO6MydPw1ORCaIuaMReaZtJYDH3+j0AeImyfXJq6v
/D+sXP6soNI1GA9phj0JS1cEaBEH15oV2UkRzo9iz4u7Q44wncM8zJagJIZ9iOUU
2sLJFHiFFNQJFYVeyufD4jfC9K1N6NZQ0OTa+Q5GZMp8P8hp0pzEGPX/SF4dpL59
9E3ii6nd8zaivnLiBI1/cTYpIbpk1+En5G2q66+xE3xLydQXFsrpxLUE6ezXyMXL
a5ggrOdOQSmi7DUCPH+rdUi7us15EjXRM918tBtAKDf0OU22xTsLyFWw1H3Y1TUR
KdCiX6t1o0v718H3PJI0T6WFktZfHmGP3WvGKe0k58bHaFcbqu91D6PjR1k3NDWe
HHvituY+VL1v/GKV5xCCd20BuzNEjQdBkHvvf/JE44iFTmvWOF3PR+IoSdEevfCW
Db7DH3ByUqdl4/xKlgbPUGRY1ZALe0jF9SnJiQEGuGBDKNxyXiBn1MbNW+45BKqW
3QxuFs5bjXfrzmTBQfih+OvuGdOM4kbAlSkBMjFZlmVvOojE4OlR3Li2lAzMbP8U
RsRtV1PIV3PWACj/bFoAyqifhBmJzziK3prmasT6ME334vZDwjKCy7CHUx1Bl42N
5Y/xL2x8xTGivNOiFAy+LXi5xctWBq9+BYn8hGYK2fNVOdxjdsgPvlfIwIsZEaJV
iyfNW+bp5x69igQWFUm8ilnsNDGBovH5X4hOdKd37jYVzCmzyvL3gzMVxkPVb8Vj
YthSj5eHUEQ4yIEacPPIYeKLblmlFiI98hI7RzujVckNswkYQZjnBfJK0w6gGb+o
gctOayKq0CUWNots9G7hY1ex2dhR6ixTk+wyrXU34r8tBVazspE9Io8XSl4yl3U/
va/wRR6LYYo46x9PxKXUaapo8tMZms9EmysB3b5JdCAGl7/a2Gz5WlobZ1Eeq6/M
mWgEeHiML+A/01CZfp7UR0ExriJKjM5SoSlG1CjdgFflzZbijYizLmD7VkZZ417A
a9o+6vs3l34m/1bYTCo5/ZJFQrYLwRgvtj7ZUfsdXnFNAvZ3jKvr1pvyrqRrAqHo
auHzpOT7VoNYrVGAxKpTZB/K5Hdv0fjRBykw2mpq0h02qMwVquNzwa223buq6cmc
xxIpu9WJvaxhpCo+xaJfgfiutNzNjiP0ymzE4qlFdIXN04l9Y7Qh3xcesUXrtP/r
zPsltqkPgN+1OjAXkyPxyKU3492+RiQzY+QVifwnGlrP5rxy5t27Fhk5cTn2SjIk
ThsKV0dC04BNUFwrgppCRGzRNoQeWVOya8CD0BAPxA4F/Kj4FpD3+270ISRMgZRT
VQNI4S2Q/MT6/M+3PbfRjdfyNtSdKJZUAwtxgJ6a/RcGVmiTTbE3qgb8GQxPJLtx
ShKwTe2iqbgB1QlYJvrlyJ3rOrzEtiE6p+SmG3DeENpEEy14BdRt6tLj6FxtXJjD
m4fNKA4cCo7KczpdmP2aK8lXinOk5vcLcybdIh9EGP8D4MI5NrKmi8VWCmoDrUDF
NPFCk+hkbpr2P7e8Sp/L05/wHvknSnpEF+jKO9xfo0zZkbUTWAMEDKRBZz9tOCrM
rWx8VwFGy7O2HTmxZLhD5VtYBKDeHtgQ9BgUPJABGpr7qm0Qb13Bay/dO6xkpuXa
+sDAwa1Fo3KkIA3xwtxGw2KLymWAW1Y3AvGMHLyD2+nZ6EbdmtTaYB00exTZn6Db
D3B8zUNw4AyBWOTCU+X/MsUHWW7Of80wxWryrYDKHGJr2Qwg0KUd4fwI4IHCN+Ap
cwBEfX/7KcZlVqA4tvPhPZ0IBN5b4QfReUTjrilKXIIHcAaPx8qam9VdBL1US4I8
XusjxrPLaukTdDegE8GrBqtUqgBZsZDJKYkzhyWBIVXpXBJlSvO2F3FTKswyCNjf
Xfh9mLBKkUEx58G6OjuFqcmgkBNL0COWnTzzWHWyLWIZHbdM8DVgpAk1ep/MMYMm
OEnah/sPi13F/e0Ocmdq43MBNksw3Di0uR7zNomIu+R44YyaP+MGsbERWvO/LbQ3
FWmISDAWNEl//KToi2srw5AK45xEplVZaklorV8SdBZhIW7EnfPokMlY0BmW08MM
oMSHnA5YBJAUkr3FcUMLZs2hSws6NpxTxwAMRiFYaJpViYQvb22mGUsvphs2Qvj6
mOo/OTHaVh3GgpkAxicQghVhHGUDSiabNIJAFmEu6xBgMr9vvv7n2oI4iZu2Ds5B
mghIufdU44b2vBhW0NdgMd9BpS4tIXXzcOSO79SKje824GLebCg0bkcRks7uoAxR
kHFbJcKzdgvydJo89YniQISRlbGBEkpgR4L2Wy07soq43UO1391eleHrcx+zZm1Z
Yy2/9qHwT6ec0yQTkOiUCn69IdQRhpuieCym8nIZ5LIq+/hb1/7XyjZgH5i4F9/0
VtUeCTyOdMnWvQuy0aHPPkFNhXC31hu/iRaV0p2MmQu/05jojgZiFvhw6vpz0Udm
de0Ds1X+7PUZI9AY7mqhZ9wA0ONEMwNOSFaa3+VzHnr276yN45WJx3TjkIWHflbo
YOPsrpOg9guCA1yG0BfJl2iaxvWBof9YIH0D6cRG56aIAbG0yFKL61FCSyzh7YBx
Jk4VzhJ6kw+ek7kpyZHjltAiaGZXUo951YPRe32aOYWpLhzJ45gshWQ7e11FZNaW
xXyxAzWmPAWi0ew6EoKdxymKRsyNxqh67eZE0o5T0/4XBUbz1rby8AKKqOZ1Vx+W
XNUoZt0yyADzk4nOT382Cqf0p2ZUsMSkqvtpqo89dMj1z8IJk8u0OEQ7XFap0Ks4
KXSlSD1ceHPWq+LvlpSKE80TASA4fOHnxE1d/NApZ4VxOgHvJnnXE5xgJauO8C7m
JJEb4OTBP7lYZjL8LG2TFf0eTIs+zrqy45TDkAjzXgfzX9h/kiKEKnhq8jmo/xd9
W0bDUbibkYGgTOYWnAi8ray7JSxEysa4/gCXraNBiIWeqB2KlOFuy12VS0qZWumJ
IDc5GIha3L1QZoYjRoJLy0Ny2PL9JddF00A7z4pHzXLy3bCBOarl4pCtqSq2EuWT
2WYJ3WXR2aKyMhu3H/wFvV9EYvNu5Ibx4nqkwuycnohyxmT4Uhyj9KSDyiw4h9WJ
AlW7SWun8zkx3F1JDeh0/KcT6hSrJrBEF6vhi5bXluQMtKJd/XvvKZreRsRt2iAQ
v8yDFWR9FBHYb7oMMo35zviyeXB1mDCaYi8UhyFKaHoBp7IC/QbihgBUaI2ch7BG
zJZy2zh3RSG8AG3OiHBbAoarPmbjB2WSTPBIzgfcrErAzTysddhBgpk/uJ+a0YSK
AdxP7mx5yLgOeloyVQo6ZVb47UbJ0PfC9tAjkPb98EcN7V6tyD16vlbl/IcDadSX
hvfPSJztRybdGrS1eOpPwXz+fNZCrKN5ZaIrf5u1d5c/O4GCOgUMjKXoNcfKSX5D
ZnbsLK93qXgWvIsRr0ueaQ1h6DZQI6q23da3GikPxVnHW9P3ToCFpbWvW0/iCb7B
mjvm5aVlEFjJ5iw+e8YnFs93pCsxW5777Kr2At3c/v9v3fqFRE528NkEP++6ddzB
+tol8j8GaRMCLZXGL6dLMJNZKJ5NtPEKH1sdnkx+S3Ym3mVEDfaFswxY8XF4AFUo
J9fhVr69tDU/xslnBXhsoOzplCROort956jDyCmB4KERaUhHYY3rFqeWo5ECtAgF
KR+yOSbF4cnjYjBXZxlBT0SIUMvhXHjr4lWNc4f/RAqWJFopjkexoL7sdq1pVMF3
bTpbksLnaU7PasaSkEkSOgKAh24Q45SsDw3peNcZlqTBdjpsmlEPCcfg5pbTGxvC
Kfv1EMDsmxDPyi2rtuEQPKYXUUmdIJROnRY8bwiHgosxck/5f6J5SwFfqcShA2Av
9sTMhzCFz8qW1/o+fqxXeuxZJi/ahTa7sRBRwCNFvvCt2NFg7SLvb4AXGmZL/p6F
f52TTVuxVi2bv3xeRdxzvyFQWK7gJoElqW+uMGUw9SiF/lECmMkn4JS9eDDxG89k
xh3xVuo+nAvHfnYKsPxZs5PniQa1t+p8qTLPvQMw3CNifg0rnfAZwfhbAOm7SBfO
MeK6GdG0ZZqNrefwwgMEsQsGriiWlZTXS4p1hgaQv98CN/sRakM0G8rGNpM6AjPC
jIFMV2O+CKKwWNzizdc+4LIcvE0rxNUX94ZkJejCyamR7Qd4EvlE6twm0j6aWqI5
GZkwsQltsF7S7MpqMAM+GQJ5i67hxkjpWLZ537HyL1yK7r/Cw3Ct03Vlk+8qqw/T
1NOpn/nOFgGvFydM+5mA6ysanEHp1Lu63tv5hCv7aM3/Yc066X200gZXhAQwldRM
ZZFpqMGMhz4C7K1N3tZBH/WLD69/9b4fzcrV7oviDfSg2KgXeD2DGvTCcS5qz0Uc
Ng7wjgh0Q0sU9TFl8jnA6cqHtoY1jtojE2vod3V48BHIxwyBe91HhKxjeWh3kTLD
8XKS6VQZrcp1if0JKCN/10v87OO1YbLb3iIhBpdp8mnkzilS+BbQSgcnb6MoS9ni
Ey2t/nz5YqsZAlceWi+BWG77YtyBAZSolGwTL3Q3OvnBwbntHzPaiRdER+Fuakpk
jeG3oOwBmNV2fUvIXoKRNOov58yHh9nkQiv4RmqJ+Yj9Fba0s2YEeEzNRKW1Lz98
3Zqf4rc0Vgd3S0xXaBzwb3WipSuXZZ2LkhvMlZxEV5C3b153BtWgXeyB82B9V8tc
GTtwBHRcssqAjUFsw5hwmGv1K6ZkArKRuO9wxv85TqbSE7A19omAg8bR2MJErPk3
mXKs+VepLDCXzQ32934lYRTOECDLlPseRa6kjdiIEeRewGFVkcKaIh4zLK1IIjjV
S3Ahp0GCLCYMuIWPL5lAX1kXLpyU+I2lA3JsKliqn2Jj+4zwHO55Ks7IMHUwL7lz
ecZADzJWu2z/mk6v9SKsCeC+W3J+4Inz3BpWoOVWmKKI24LaRjAtHtPjbIq7K+TD
ABcGa1mjGz0JXDGfbVN9/beekfSu8DGIst+aiF9bHE/tpe7To1YdEU5X0EuctnFp
jmZDHLa4fN+y9JOvyp8BaxzXFdESPI7ThAehjNnST+193o89Jpcn4WQ6kZT8cp8L
5vokZfXk+hNtSgPKkp0xQjE+ZjS+Il7lGNqBlb78f5tYGR0lxfqDxfL1UQCIzbFo
PodCbbl8K61HLphuqZ2w/VhVG1yu3RG9dVswjLlUIBo1GhVBLpbZy5Q/gawekKwh
cVQD8EVo2OHRy5jg0cgyTSVckfmYhS31YfVinBXxWeHOu6oY7gSL6DDU6xWlS/8S
`pragma protect end_protected
