// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
D9v6O1xwFHn8zuUlY/NdLwQwFDm7ZfwdRP+AqqtomDd8yN8ZKNUI7jGeL9kbnDAV
ElHhty6dWy6dgt4SxQP8hmC5cxM76IasHneRmYEAZuysf2b3GTuitY+dd/X8azVO
8xbagSz1o2LTrd1EwmJgCuxDsBr9maXpTMSRsMzX0eU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19152)
+vaz8qu7e0Mdm0EsNpz1lFLBzO+YGruOdBlKTR9icLfBNNakzcGNS6iXQd0vd2JY
p6O+E2AAoK7bD8CvaA6so5QaiJPBzb443crSR//Ln3TZXNsvKFhvgjvEDwDd3CGI
sl7Xmxls/MDxRWNgIcGAdYm2Z8wyV3z9VjhHvrUn0dXSn8gHqF/RkIWXwb/pMyk/
Zcnf6sOf1YobMKTSOnedXeSRy3mInq4vjyyZRw/tYg5AJOG6Q2ORHFeaZExvihg/
mmJWSDWafyhJ4l6czl5x755+W1mfAoQ1OOg8/Z2AuKBhZgqGt3X9kLv+AnH0TNBX
NU5w12DwiIhQ//NF3N70hc6EXFGte6LFm/nOfHmIJ3lDQYsYLKEAPychkLbZ+Uoo
99mUTJeeJ1/Eybx6cECRnea/2LNEHNe4LO8YQoE+idn1uNocnS/cRd0qlC3JjiFj
BlpTcdwFk6dbzZBpFErV1n8W9qB/2QmA9zb6n54ChperFFw9p8Feo43DLxB+e/mf
vgHQoWnuTzkxffN8DNJBT38J57UIfVj8ABmCmmtVT8bV0mggI+dWyRXP6SbxGkuo
9nC0EglNekhZkIpzKDPHzA6kk9JjRoVxQGJD653OBSa+YzkGlEjUoBab/m1FV2VO
Mbj3KadIjXo1s4ZzWxSbZt2pGIBMsOTF2AhYQa/5MoWyDkbS86QkiBHeZnJ7mVo3
wk0c5YL3kzAtFBxWtaDngaveauoJB2rItNPiPcbkBEZ4EFZA+hF24OMoVuVIA7TL
kbnXRR5eWF86UtDmRSh71SicwdQmfVMJvl1RBxRBJsA2zl1/V9RhpR0dZCWkt248
csfdxVfJjRyjUmEZWDtl3mxtptH0kooPWBBi2H0v9hQKct7SWgKf+piLq/u4IhgA
gMI3DYDqBG+MXQktGao3NXAymStkIhiLdx3vSlUo94jFlqgtlX9Q9MQBtyreKus/
q2WDY6ron77R/ea3xespbcLOYDZ1941rnY/IOktlzyimsi/L/lkrmo2YYvePyK9c
21rzJ6IPAIkn7itqgI/CrBy4Np/mcggGlth8+FX28UgwfJ5Qx287R58f0bmH0im3
zy28wzBWFqQHsyKK3XFuMHDyvWGjY7ojINdhw9WdEMaUu5o3y5bTpGEnfNQxJLvl
6gHdYavjnxmAlbyTpBDyJJPzLu4sw/GO8YlzrqOQiFFRX1zSpUgtMvGqa9z/QJky
6uKbkltMzzmdNR7qevG4d2cwX0LWvanET28ljSJW3EEpJjqv9b1mC/2gKh8zhGd1
59+5RhnMltfop+5d5HC49L9QoOfEOktFI1f/2DO4XxDlTzioi2md9B5D+lZ0jvkj
IMD2qZfV5+1BUK9mPghmZpMI3/yn5eIHwTSij8LsvSzB9kZin91iunuHhSwsu6si
9e123Fwkzg/p6SxMR5SmGugNYsD3R2nWsieduvkI1Nr/GkyBGBzB8BVyeJV7pDD6
CAsGzjVb9Bt+G2h/npL+0uAZmiOUPRs6sAOdpDXqoOp59kfQoYB2o1VOnw6uLK69
sX/AhHFBS5K8yFhoDTQ62Tb28+wrnQ2/UiYRtG/2xcBCXIV3L4WVMibPygJrsIZV
uBYTdwS5DW+vF1IjxtP6kt2eqiTZJ5B61T4hMRdBJL5Bo3EE6njvauf96KkTafu1
/0iWHCrStEiOhD3sN1CKVR4UEhjgG5O2GhbEk8O+pbMz3fbsYbNtlyf7fo4DhhfU
5k6OZlpW7bdxiPsefIBF94x2SdLoUXrwqgVI8V6nC03AUuh5PkOzD59W1iuGJAvA
8m+iYmm2kkeQomw3EmkPEeCOr52Y0/FiiSViYJ5Wa5M3wqviqhz6fbuejXFKl4dX
V5uFBNCNU5mLv0nYRo4JmElBVLPMxpwTrBo3ETuhRVHTxOpqH0g0EiXfQyQdSbG0
DQwhfDdSfiHAQrEay/tJzrtYdRs1mT3q16vF92UxNcFaEd8MjYaqR+x11yYjRSW6
yIk1DzQDV1OyISjGX1ayeAhmt969E6eSjGeYcdETqMLk6AwX1xcEvUpylzyNJgbU
IWuIXlzjuUhkdPQ4dH5TwAXHGqZRSiAfgGdvi7yBF481NX4BVedosPu/8ADKqLo9
phfFYTeLZNCkmZ4QjJ0oiOaBmJk56uP+EkA6Pq9Tm+MKF2G9NHP5YDHVpGCw13bo
6Q+uTV9GXG7N7swS/nZKuOKYfl+wrY5yafZigs7oFTLGCsmoYMz6xvj7vMpaNF8w
AchuE3SYnD2gl9bxRL2wxGHTM//DyJ2d0X4IFmbspX8nHNF9Z2zUi0VhWfGFB/QU
Ver+hoIV9snQxPz/I7tZa8bQ7gUkw00wxNb91YQhFJGcF84qmkCkx2Z6+VvVT0UN
dGTgt4NECqxG1MisNKwGoEX0BA5+2ZN/OcOey7wzDBsiXv2bZv8tnoGGuDlljAnd
iP2fGMaN1tPr8w6c82Vi+82WtzFaYchCASiIEn2iPtgKfhfw5tbiS69g1QPwbE8a
CH8XN3hS0fgYwwLOEoNGn1ZZIUq4hFpsB2GcsIOrj1dxC6flLz6Eqpvge/zL0Qsc
afqI9DLC6YRLhv9W7Ze9spr8tcjGcibMCp/0D97XHYEcl8Y7CQIZ4gK6k8bow3Vt
7YIDGU3SZcm0A5uM8ZUG9iUmnI5C9hdtefk70MYUGaGNgTFK5V3/6RfW5ekDv83f
IwQdzEKGQRaJlBvamiOhfB3NeY1W8+Atn7kooswMcjPhMXgIjIe6C4ZdUC7JK+8Z
+mv/o63qIXe02/XRsNpS1CdWFyGvAGH4XIEtigpJbjVn3Jo0AR394mQiWaRQlkI+
xpDv049IS2Gz2opVOh8LCbhHU4WJzLzaUY1G6ynwWcZWc6nzZJdLRtyAHht5SJ7U
6rA5hCkxvxYAOcAvnTeEWUEyKM37ksM+njAfk4XPnzNJJUcBmbsz0I3HrpXfHHQ8
lyUPfQ1n5Dx1UGrwEJmw0xiWb7KbkjDlbMAM5aNg4qTOeNihkjgQ3On8q0Cifr40
k6JeOi3LxDJ5C90xbUOSR+vUXxrFdsK0HaAbdA51AnTI+mFIPn9mBMAsIwng7OMQ
smBwyftC+1xWTDkt5k+OevcKUS49gDsb4mh2uAOi0HmjkGmdR/00ARYm5uSMTcFP
5RAw2E6xL8GuT2mGacghI5AzQ6HIjJ3wLeJQmuvGvoL/IkkqVcjquxrCgIsHD99V
uBJk9rJNbR/GcmQH3CWIEcJbzjdolQucC1YQQbL8FJ6kIXd88+Es2nxSolpLcT+8
7AbPoK64fc5+toKrByrthsCN4+YiiUUlHKV2/zUwF/wHqvmSW4QNilPJpP4GTEv6
JqjRY9pxBPwmCDENOU/iDwVQo4UuWT9Y4tA/MZ6uAP5L6AMFKS/f7oQa43OfxQMc
PVQDwrgXB+HnfJQ48dZw52MilcQXYnhgFg8dfwSBjzF805qSNlYIFjBsfpBihc+X
EuOqptU0bxUZhhN5dmRMBVW9/75x95AcJQnYLh9uYeIaLSMuDCipNLM+iKgb0Q6N
tVOQoXu3aUyjdGobfkLxgfVNxUEJNx/TIoygjwf1yuGDrHibXRUM+EqRJoLUAN0E
dmgOM4/pixRrWtPEmKxacEE88FKwyD+oJ4t8SNoa1dL/17ffeJnm1e19ff8LXBeK
jlwCHkkiOCItRsc3ESNGhkAF4Shx586bi17g9ETQgZzXST4/nmKZAMar62fsBZTe
wdfLHSH7E+Gxfm6wOnaH0mvOW+9dYysU2TdRVuJmYcwxQVmirV+c+fw1gshD4/F3
BB8/NiWdccnHY4hk9x26ihhPtJaTp6pHYQ6KHzvLXTTQzb6FMGw+3jTbq0XmAUDr
6GhMkfSJTwzwgJh3odU1AhsuOKq/oelCMkLQsd/J6vuh91YvIAGXvzUqeB5VqTIZ
bMhf8+VWr1pX2JKhu6eHiFWZNj42UjQ5ZtwrPATaPKUT6zB/S19mA0ssECLxUnKp
8zXCH++wPGZKkjwktQ03hpj4iAnptr3nQ2/kqE0Ab1bHVO2iIP2oqITptR8KrjPd
a4sQFLwNrDoj53/8sTdO5tz8cddtNAlr1UUuIrMbi315dFjvYjVzlwFl8o4NWVz3
WHcCfY2K63AMFzRtO7xZyUPfzAgnnQd2X6Nk3BRef4/lPtaeG/HdzBpqjCfi0/+b
Jj5tgkgCsyznQvDNE+tdrf8HmhopnUZpw6Tq2OLOVHtp2VHjNk5XlLhWfgxFcsy4
4EhWpDEK/nX6Orl647N1PAgwCD7V2KPbEO6QYHMV8Q10CkzK2Mji1pFGHvrPjeTf
g0JaRdDjsXNOtiLmM6iaNKGwgiBSZuQyQjWHjhB0kYFzBeLPtXoAnlKDnieVAVHl
vQM/pKeGphFFpguo9aICpeAvvVVyKsZN3ZOAK7ZePjpZSk6JdGtHfdT3ico7xwvy
6ibLv2w9f4nDIksGVuAxoCdzp47pStSMKfYIg4Jpvd4zSfCgAEvp5Zmly1yYIkLl
V3EnqUyQZsZ5ktZIy+3VtsW2QMzUe9ilBN/rYczNYkLuPnnFK4IV59czSUSiyKPD
TxXC2yUNXKShB39iOaiR3PP6XluavNXa2/ROst0eh56Eb3r5itq97wJPto1jlBrl
SUcHxUukbhCAP0AAEiTXLTZ2rrqL9RtvowMcjWCJKZXAT3tMslnw/dylyTautp4B
7UhYly0IWiQOS0ME+CjeSSF9znky1hO6HwH//H90JQjeA7ImAG4Nu/2kPL8szuve
XUmNgkuDwWUPkBMz/tovW0UTBSF67Z1QDEjGNBTgp0U5RDOPohnoZ8AQNE/724w6
9LvzKKveSL/gjnA8I8wUuXXDFa9eTwShUObG9dyGukEEbdy/8xsP1rRw5YYN5Q+B
SPfs/d2zNCgBQGo55nxpLhar82XMEdB293QPcMJJg3DjjcEHtOsOWBi4CWPi4uG6
RWAyk5rDWwzVagO8nZzQi3uvYI47hHdc02o42dixjSiDDBNd0blF6qScynXiXeQv
3zs2Hb/PHU794nW/K/q44+p61Jwu41FPeF+rkd4bak/RuDgzltegJru9ICJu4sbc
/gGNdqmRMxjcQps5k5NDKKlqIaRnA/LlJ3yx+sNI3WvNapKmqc/LfrK0en5MlsSm
5F1ZFeIwWTdH/MeWiv1quE0RMmJx+d0V/E/5aN3Cmes9Sifp/XZVcO0nG4j04eLA
yZLYeCF2l+PKg8qXCAsRu/1jwLfSTXDEaAMWwETdIcfFvsZdZcG5olRzUD9y/7RQ
e9XRo+sykmbT4vVSjWThsNFPyUXWKWHRBfu03+fsXOvuKGhs5CZWV6N9tQiFOPXl
WMxCzg8h+7BcBpapkbEHzOVDkQW85z14DE5AwISuBt6BOzer0+phntrvX34NYWMB
nHxdyw/MIAWjMGdS+FctmOtYEXoHKqE+vD6f83V1mWi9r6dwa/0YNxvetP6+dYUI
Jt8OX32jdl2Y3QXp35rTK9YTY92fAU+5V71/i9cPyHHU4IC3vUVDnDv1RNnFIw92
+Xpsrg4eldEaNijU/eckdZa7pGm4GxutkRvG2HnTOb4F6h8wtcKaXi4gAMf26I2f
5Bmsg7v8sBvSjvYIj9Xs+/KmKMX4VO1UWJaUykFpOSdbR1vYeEG5zE4f/tmz+uhN
O2iOg9iZkAmBJwppNBHimn0rkWOaSDAAvIu2ALHlMb9uzbUYANfBikqrJktXT/KI
bUpQpG3iVEC41lLr5UC3/Hac/7PQP9kqz1m9i3tg5h+aa+0m4tL1rIAuYSHPPPis
3BO1jWujZcg16EftPsk7EOntBylJwaHDgT3ce5QAaBrO5Z7fFTbrMhYS2yj7OK6D
QNssCcARnZUsNgI/RFIJFKxXlwQ6BvlaS4e2P7M+HULOWvFICmd25HVkdfibDwYI
tyJxvfn4YQUOTFyujfliky1rtsvJbk9ba8udQWw8aN6wBvaNjcPSpkiaYVfdjOTH
kWQw65jCyBZclkQdf8oqzCO7BxvqH7Jn9WmFWSK/vVgNspKzXYHF734N9j7JYcwV
xcPGgPAbz9gTe7vvR3arrq02hYUNgfdmr9lrF+wAmxZzSj9/BzeLHnsXhFsL/EqE
Fk3KxYnt6xBBVXKM0WFbivr802J+TqKxVjfM/Pivv7USOzlgO/WG00dD1y/JPgks
ARBkhw9pcg+RwU7msvok6mScrDqYWynsrzzxI9E+6PSJFKefJ3H6bxHdIxm0MAht
LUhMF5AuleSP9sBki1ffHEHZ4eteclmq4SjNvnNJQcpZJMweQeh2IVIln9lf7O5+
7YqIo+nCjKWexK0EV/5v/5nnjp4RnU69926oWmxR5JO2HtUnj/kG4kN5NJAI5xav
rJfnwp2Q1virEhAgqIO6UsKracM0OtT89Smb04DUTYUPUoGq6IotX7fUiSat2cx5
GEN2Tx17TzkY+opb1dddHIjCajDWGTyOkLtVNvGB785FWUknSyXH6TybS3kp1vhF
tky8faoYoZOD81LC0UM9y88hHYFuQv2dOPTx2Nxu2csQ20EGMZ63EqR66GjI3Hir
F4btEELcnRrugDlZFcaFSkWkU3/pZ1g4DYy9wXVqbp4/0PaJpmF6Bpjpsg3/k5eP
pHGeG7s98rHptB3JJzvvuz8wTvZ5+zpnfBgnC9U/Si9XhhFlvlSjFm9lGuZhnPuQ
JtkgD3onItP5HX/FXAHR/xLgP+XtMMgqKaJQxBEpk+yzqso4n3PGYt6zaGdfjhXi
nmHS4e0B1BWxfSt5Laq/3J2yLnVRqDz6C3CSAZQZWEwRRRBv/M2T3PaqJAGbKgj6
NcgpS3nUsdcEGCindd/odjyEExj/rV9P70jjJEjs2HjLU2euDTCt2zwEIFP5/Vp1
tgcqrNiohI3x9YwsVDo10r7pZuaVc9kaMNlI56AS48ttbKsGcmrpk7A8iCfcfqUG
derUorq2dBnXX6tWok2XeQnA3luI12vli6FcS0bHmRREKARBOI+QhFgveABuof0V
n9r2T7HBaPs5bAB5dmjGU+1xlEO889bVAcsNcKekahkgAZS4OhKfXOZeU2v1Ti4g
1ipnaD26LtsJOPYxTUSdFc4jmoiHClLPqEZ4zLl5zxA4kRzQtDYJ1sdfJSzoDCoQ
9VDpf0iJBraPwxcRQfC8BPXa0lmj3Iap5IGxmbutf0BkxPfdI35zoshB+JqfnYx+
4lZ5SNJhKeVtxMdMlnL5L1phJ0OX96WaAKgvWVQ0e/K9oJ4ihy2KqmT1AwkiClPr
ZWrPFugyXX+kLKdkyyb0KA6LPEMIbJVxmnZa2cszLs8fa0iKxpkbK8QiYMVxoOa+
DQ1G1ulUv+y+YpQnknwSYJGvWRD3KlI9hvruloLf1raalzGHbZzhFTOdsML5N7OC
+IbFFVV01DQQVMvHheuyZvhPTFoWkwmbzfZrpTbZDsPCFIflKiuDx2PowWgbyrOO
21w5uGI9armwz0QFKyqYgvqTnhTC4fwNOb6cv4ipEbVTvQdFQ+m68lNOEUJWIb/2
60RuTSTi87wMxgdPfdb5S0TFfgClvZ2Pki7D65wYoLER8nNW9MxPatNhtJmFAAOa
zE6vnIUxkE9poKgSpO0Ev+1SpQBL4Ef8r3OSARN2fanlo3heWL7nN0hcCnKXhyi/
7/FXjuZ50h4xXkyRqkUrRXE4FBzOlxvy2yItouvvKdU9UWuBk/qVq058cAJ+/pC8
l67oX2d4hPhQFKaPI7gvYzU/nyOMbZ1pVvPDICUMONf50MstiWlDh7o2S3hu+p4q
awwIYgaIfkAqZr4SPHLeuX1dEJ3o2Eqk7FRH0jgOOw7oa8isegs45dipqx0E5Eqr
6IC360MiHE8o9BA2Uobj/raNt0J6imyp1vl7qTVseFV4Bhs0yghYxs4S3qMhtXA5
zgwLHd4vu3y+1DrbKp5oB7jeZGSZPGk36cWafDJchef0HeI7S7CqDLcLL3PC2nVb
fbDoZBpG5mf8xwx95yYOWJigNO7eiOTNcZGaFWnoRdzg6UYISldFK6lqb79z+pxw
Xgf7462xG72jyrI4FNZ98MMbtHyVE1X1I1aMTnQWIDinB7ky7xV8s5fUCie+Rxzu
P8ZGJ3i2/iCR8Q49IDvSoVVjDxMAmkrQcBHbR2ZTmy56LxHQi6YakFwhLjt6dYgR
336hMX277TiJHjq4jZcyTbnWzUlJoo/NA7YsSMz4T0f9GB1ONkv4/l9c03l4X7vo
nFR2IosqsTlytXpEEPE+7kQE8+M7BKm9qdvv6dErdb9yBpCYTqNQ8OPP49qJ7teW
Xhrdaz4RkMRmpUD2pG6dcPd9Hcb+9Ax2aNhlCetZLr/NncdbXbegBPSU9yESyVnq
+xuJfvv3k8Ok8rbo/9Uj5J3pf1shriGinkg100mQqvllRi7Lhtss/pdjTav2gWFt
umDV1YrmSpP9Z9GzKRHLLarv6wBs59DJPbZeqkIyu2SEb7RHKjIB16jGa4CzENbf
9CzvsjKN5jKzLv1T2SPXcJos0Dx5SmmgarXMTFjM+l+uoexC2r+Zx00rJXJXxw//
EJzWXBzkVK2eYkRZa12EJT8rf6q2GWOVo7cLqRyS9YUTBZdRONLoc9/VakzXzf4b
Pvqf6UZc0jSTkz76IDU+fT4rdbMuiHiXH27JYiJIDHViYmxedLgadbY2F+EfiBBD
7Wngutcg6axmoeVDaKUwDLC1ac4Trewnmt2SyKD7pHPHNCSe/UcTUXhLkwrPShhn
xvd6H+24hKidG8vfIEpYu7oDiFcFDhS+dnS0WFef2/HK1Lr7u18e3vwn40kz4oEL
C/HtlOPwt9xlyfv2GS1n0I9erCQRl5FrFCHLbWI7PUN3zCpP9Ct5iazBYx6TUSC6
ERX5/OWbIooNW4C7EKs1oCVuJAB0g95OyVMr0HGZjbQqWFN64QGyUj/5F8599ZCn
/O7mM8rwVKKuiz13vOmhUiIG48Ivrt69hSZDfWbucyDQSe9PaOhB41ppBrK6yCsw
W/TkcrV1519a7Y8NlKUcRHyZw7ygE3a55WvjhVbyHo+7xIzNd0P7e+W/iDHKduIa
YdBxd0/n7RA7Dy5eqhoXe33pEon4TwcDOzOk0HvkK61WbTsP/zzBMBkvcdT+mX0U
YT2nugm9cLTQNo0KrHVSO7Xae8msQheVnhiSLA3ZkY7eKL4wpi25FTNkMIq879c/
xMqDoH5+RL49qxuPw9RzVWPx1zoyUkQxFP4ZzvbS33atYhUbbIW2y+oqOJjRd9Pg
9ZD4StxrtktH9gn10vWS/XIv1mtzUsqP69nyiSCBkQ8LDNd/dRLcr1xhQHDDv3wX
mL7K01sX5KGbexpniRIhBYKTF8c49X4k2bKcHvWxJxBij3fdt9AiXwCA0zDIs3Mi
TeQTUsbFYiIl10qYnWY+6bICixBnkrfIQ5QE9gj5dGRrGEGQHLXaexHOnVunsbaU
aBb7sIqjYUe+ldlDFVBimBPlwLMzL9GeZTdc2tyEukql/xacDjDUgXd4dYymBl/a
3+ZF7aO8BHmqDJGQlCJI7LaYn8Xn9TXNdgpUil89JGrXTJpFWdthTJUVSDoe89Q/
5yY8ETG+sYZh6b8J4p9K4ovffAkZ2Ynm74zTtGb0wKIEZUy1pXZ6dSOvZdKtWKZZ
Z40Zw0zuNVlBUlY7DMn07KUtkQzk20okxFLinTZuIKe4AJtMj2L43TI81WxXcPH3
rQG9rZhLOKGELwAa0+6hCKjEXGCu1roxl2JWxYxxL+enEnr9Bk8TP7yYp8GF+gCw
o5Kyx83456y+0yEbK4w4aOxNUjdXmb3Yj/3H02WZmv9hiLO+i/GaANcWhd5iFEZv
JPJ1o2xtVuJyT24uiT4LUp1yhHYw0b/XrfQU0jAtADT5FqKU+7tq65CUGOVVvFtt
R8dnILb8NgPUeFrCNf3ByEt3kYDlDKbwxSEEfHTsnnqaUcTH1xC5Q4//8qj5owUk
KLHT1KGSB5JMA/EtbpLF8MYS2/pCzF+AIbGu4ZUk8q6ahzqLrxhmWYmap3VPbB5F
TFmjquYjHXTY2myCZ9FxqCpU6HtLr8GG29D/9rXM5i9qirP+EnYRMCptXrYaIQwL
BO86l/3eB2uuAzFv5EmOcj61QfjZ2zF0pnjhdrDMf0Dm28OBDQ1za5zhpqz1D+vV
95g025PnJsCj9xQrnZOFyAavonsTvpeh9rBq6eB2UGMup8/licmDUIrKInFhhkWs
60Q7e9kYfhoBSF6S+O9Ul2LQlP3Lct/vR3Gc0tLhHd50Horm8sVyeuyRUv74z78Z
5btPJBOZmzyEty8djt++fcmM6AKLGQw0WKDbSB5EYzulKntELmzNHUeP/k7KCOaH
ury6pImq1eLwp0/1j2qWPK+YmPkAO3w3Wjmjdt2x69utb6MwM097x+lxhSFRw1Xn
s+fW8xcKCqtwM3jttwtQVhvBJ06J/lhLuwH08PBtCTmBVKhhIMPvysXK+k0r0BtL
tkIzlezeNv0ZMpSzSV+6jEKNVSPY4/lXYrELFnp6//9H2nhVYUP4pSnqhCsEdxK4
US6qVadqqESVcmxbBI70Gxm4nS8GcMKn9ku8BR8YWHXHJOcN9m60UIi1BkOxTr+L
Sfgemn4N8EPpmaITEsNtVD/n1uoz9MARzNNvkmXZqrrFOHHEiLkgzg3oMoDy7vb4
Ck6Qxaw3g4UTK0hJKr4OUcy9pFxog45ketaRuSThSOk8RJNcjTxJL0e+uctD5PHz
mIWGUI2ExOV1J+rHo15XKSGDlS2DMQ5eBmDXpG/x9iQ6B4tL8peJL5Wgttg7JLZE
7+P8sQ/+j0iMZqo7/f+8DJv5+7JUNVEcH9z4SoWMLa2oCrMT4yeWC7chil3uPbwN
wJ8Oq+mDE9xfOsOG55vaUFSFAfk0I4v1xJ4GO4FhI7RwQu6gVHC+HbRYJ4PZXNOl
P1CoY1bPJsg2IOGhQJnbG0u3SuVjXv/xr25LsoEb1uRwJxHLS/JBtl0N+iVjhySb
FQl7eQF9MB9ozt624xrJMzD97wEFVqa13YiiO2zeMOYM5FMr5U8N00W3DUyzca1N
i/AMKZdixnKEa6xJCqQMjmPad2HUY9QoxkzPKvcnPcbFI16ifRY+AmztVI1aYWSy
OT+//GlFPEq8FG4+BW9HOaM4kdqlJB5dZ93sPV9mDTAwLb6IYwzc7sok2cC/Sdnu
APoluf3Pq+l3OV5zkc3a0knGjBlBwbh5JObCSqiug6sTpmmETLdO5LNkI0QrjMvY
T62ohoRXY6Tn2oKIqG+TxpTH3cSCWV7qHLjRZgbMD+bwQF/46OFV7RYv2QhArKGl
XSJ/tuH46W9i8cas3VY3KCgUf0NBS+ndNC1HuJuDVTFoBRsdHWVrgF2rNZhlPlLx
+e7aqSMrGl0uHc/TAkZFoISN7UKH53TGQD7vEWiYgjzrCGEg4n2Dj6x4A7mskWpN
tDs0f+sd4Z1Ys379+vwVdrMLW7kVxWTrvLkhxQC8uMZ+AZgduum0JdJFlFP28kww
PTN8f0iZKiUYv98d84Z73HAoCgD2T4zLewUxZG7CNcE6z8MzGeMvkVULr0MimCSx
biKt7sFGMhzF/hO4zX/EJtf/LdTrpRr/aMPRdZCSyuOTY9NUi2gV0cNZ/zVISeE6
eY6sfxRFzIFRstiip0PHHcGH91bCU3PlDRvNpx8tkVhUvDqWPQSe+l3J8c1wxf8U
zLlXdrQuvCN1lMiAeH3E5CUPpZD+/BWz3XxSzxJ7ZOdAwH1uoPTedudSzxSFrklr
qdBqubYdlD/sHRm17Rl1bEZ12Be8HYlyrc9alNrqIvjEYaGpLVBSYHIaj8OwMiDd
RnNgLBD/Yai5AFnSL8e9aDXLQa9GBCF7qop+o8HiRRqDd3BHzcr178t9H4ou7lWQ
NCZaE2Ryll5vVsmiqI8smZiDwFs9SFTs6UgiWH8yzjNh9n0eDuqqi3LmxGL1Oyez
fkfQK/+ViJByGRMF9iKvl5JJoNlgE441zOXIqSbw+YN8zIOEUBm4rtvZf+cZ5Poo
3x2B6+wuzZcVPYrsWPCSjRhl/oPq0QRvGF9r4iSLS8oqvERI4TQ6ICbxb01iL8q4
EXCAl7zGIc7hD+NeFVD5LQqfokXjvlkscPu/fzfRXtV/MFvu2Zncp3gzFHoQW21C
3f2oUml+PUaOOx890XybUZpxfgPeaq0Twc0b+aYNfyAHyEDVrKEj16tfbJMsEpBD
SmPfFDxejQ59dUAUOeWrddtkROQhe8Tn6fX7BtRsdgsplYiz32PwN6QTYOzqBtXh
3s6oSYuVFkRl4HrU0Yfk9jUSh+6CasLDkEHaJzVCWJ01i8JE7heyEsyb7J/tpGNu
gFPxeNlru6D3H0Q6SyzdMuabCT2UwnTrz+In3f1mFDd6ik7BfmU95qW6Oq1eHpBx
WKVoECP+ihQ4Idrj8mDnlRCJJhoWktUHsLXwByNIbB8Ggj/CgzhsUP+DvM3c2pTG
DkFTFcBnbInsHzGikAczNT2dZqwLl600XnbTmxrsV3JFeAloYXe9GUHuwlcy9b83
uK5t9lZOhYBayj1HaFEca3zS70QKyC6Z3y1gfNYG6dVUSrnCKdqjzWi4Pd2u1WaA
N6mIioJu2r5VbZk9n28kSR52caNkXnmD/drWRQqs3/kzN96YgEpl4vGtGEyvBMbC
z6w83EW+sTj6zef7j81MRN9rOvW1IQJxpEvAZV0UbHh4CHzkiOz4/uTv881LHwCv
Va1cEcGb0Zh7P9rnTxOyR9h/j/Ji/28GB6iu8NSZB89JxnAdUCYkzy6Lda4W8FIo
xEHROmZ2mFZtgX865oswqMLeQA04cdouehdFMPKdvZ3cfKRVnWphc5T47Xp+IfJ4
zb3q7aHgU/QZ9RLp6UgOxrAzp6Fud2XmfomxTWn/xyuPxv/NYRrP8kJYHr+1e+Cx
kBCGeXm1ss1iVboI+MnWogO1+of3JikP/YIGzVSiDZDUO70qnLArOuRDTD4bsLZy
pE13dS6i2UXoDn8Nba3UXAldYKag/vWwfav6z3MwMecX6HhgC28gH5RmF+4Yn5mu
cvYqv06CNiURLk6uckrSYIUwnQBL8osElprOZWIIEUeriFJMkXRen/AwVOO1XIHS
lhLxFmiJDvc0DdUQ7VB7ELoIly2l2NSCUVH09BnSJFa5EYmqkxVPlJh0NAfs6xr0
2dgESO9qDdYzbXqWtqoCfX1j6YMX9hTYnWksq7O0pLUwl5kUGeYjHiy5306aoNHY
Tn17lF4OFy2wYDzlO/rhr0nRFwAANG3+i5qfehOAyKxb7UhL45xvi3iXQKW5Ev74
HJ0blM4gNgdT29ysrU+IhgdMqt4T3jqjwpV7UeGO+NlIzcvgBBXWLWv6vHjerPrR
TwT/6T/goqzZ/i+oRnxl5QP8GsiQZY/JRFUoMl28eLAcerL6OWr8vwAxTt/nj+BT
gChzNb52vXXB/MFUUlT719XkrZzN1VtGL7tJ86UxTzi0uhfx4Jcsj5E/cLfQyf0b
F4//NDo9X4iu7hwyXA9bgcwnfKEHgoEwHE2Mf5p8H9kQay9L4t9GCO6wG2BiXJMm
Ca2/nnpvHmN70C7bK3biqMxPw8p2ObTQ8ho5aSS61ms8D3h3wkLR/kuP2rlZpvaF
MnNjNuB5zxABW+NRU53aa8hSLLOtLnR7rtGM6LJkYAswoGWP33uwv806n8QdMZtf
0ScCMeeXOomWedv7tnlEIHdlkZG9nm3qKWNGBRLIlj+7Xi05NbVRrIMGTwWNcrP4
SEdtDRXIM6mDMYlTA4PNY8MFf5HymjgZH4mJ5JtyyZt4CcbpRTWueoxivo+bYJQS
PIAgi+OTYBpU/jx8i3wOazYz9GhP2kTHEn+2IqorkFlLXcgcnyMNzFKqsWb5oBCQ
GnruOAnmHEOJi7CWjpY6qu1wp6w4eD7CRda+ZTZHjKYRkdHUbmyLpNLKEB2qDPrZ
hiptClSt6/Ao0bpx5XTedpX0Jnk2oLpVRwLpxIb0GT/CciJb2ry9bxubG5jITSlb
3ZOdUBj5TrJXY1ZISWJImxffX0OcfjpE+mDR8RCbln9k7onnfkgDSfbXCgiE3Ff+
kqjLv6eMP44EzeZ/EIf0Gk9jq3qiUkDFpD3xDbspHwdkY3FRc0VFh8JbPG8L2XeN
bEWTn953IE2CNPovoZt1bwCpyUv9JYBUOHX694BCzfz93BN1wGRuEo/0zG7yi29t
eFKbqMAtuAu5sL9nDIqu26l6AbxZcg+BO/EPFInn2xBQv4Gj+N+d9EhnYeLsgxXq
TqKBHZBfuabYD43PV7nhAWTdHGSon/Kchpfu8oN6C4B70tTUPROJKy8OJi8EtDEW
CDcvDjUAQ7LzgxvgaExXNGGozGBbfGnyE7/37nFKoBfVkpVRAHR6aHJyQ/hImX0t
SSyQ8lzoGSOQ/G41AJwojrRvAJ+C7JQOcwSYLOPS0xd3iHB8fG1peTtvfizjlwP0
F9lY5dwAU8aS30hTk1rKc+2XycQ/j/lqQd9Yw5++3IXWT3MHIQREZ4n1NxhAvjbu
mRWD7iUWyudQE0zsI3nQonBqrFyRJn7SwPuPoTUDTWySzn8ALAdyZmn5uHpzi/D3
RoM1aLIRRMFjCsfT3rGz49SGJMQcDHbTZOMOrGQdNgxrxQ17/ck6c4wZq5zWW9ga
aGTERyoOXKV5RQ6zL/Q3Y74P/CuqL3fkl/60lp+vSNVT4gTcNP7tLhkigvwRf4hE
g7GU/rCc7/3OtVi2w9Gr3xRMgW0CntRP1dPKpsiMzX6lsaqEySkq/P4WlXY5Iw44
n3RpNZPMmFQgkVWBEm4f0TjjUHFGs0blCNFhJ59Z1oW7JH84C593PPhpWLtZYC6I
w9daWYkmbc2OYMhmSSFLTJgqd6T1H09XuB8vaM7tMhr7gp4vpTJPYLXss3Pdbd9K
3hZAZ9PAiMU80ng87FD6SCxGpiivjDCcKyULJcQztg4xEHmxcjY3Fi5TUlo0NPtQ
DZO9WS3htKdPoNSh2fv+AYB7PtduKg2urLhsR8702Bx21y1eGf8kCTLOigo+a6yw
8WOV9oBCUEdAu4ZLtXrnLZ2ssi0QZbD5eGvlBFmC4SqhJE+o3kzQy4AFPOpkGTPX
97LWbtYJgmogzAGatdR4X6IPfbqUjo52aHZhv4cxS6wXVoxYzI1SRjCzMgcZchMJ
mNanPQMYkq3m552gdt6nTWI1T+5PZKMaA+M/4R1O4+TI8w4PbkHA0r22/SrgsojC
VDDNOkB5sH6CSxvJZxoIDMevZAggqzImbif2dc2C62G9O4EY+qdqSYVC0LD05siU
LbKp0NMRHu10ToUqaHuWevzd+gRb3/X58tCMyJ0ggv/t6BZ8rSN9VTB6NqYVe9TQ
d6ucsIMsfD14EcSEUkTxrJYeI0XqV7BgEa4RisKmQD+mKrgp1WjeLpKymx866Y7q
288tX6IEuTK1wyXKNtZl1hnEfH08oVeTVNUr0jUBLxr6ofUyYJu04aMarGKPRmTL
mB0q4M3i39I6fTWBOF/P7m2hTs/Ve8lUfAnQGleY2ZMntUviBCjp+jsazfxb1PuX
uz4CW5VL/1DR8A0s0fUVeNUvVx/Qg7K1gQ2LeEytuMe1ZSp6ltThQU6TCQC8aLKo
WgOalOtWUrsmXKgMFlUCA3jYu3WofZWdBMcUWWku0zt8zO8XY90dhPthuP7oMtYm
+yEIpFxQSSKngEgfUKJiOae60r25uCb2feq28/m7uDBL75TJZiUb/pINpRtTATZ0
ZNj7Rpmq12IDbqZUWXgmDowCHomvDgiZTjktYnEZE4nL+6B+yEuCNvyFzWKPk5+9
3Kckj3pgB+5BILYMYN4d7XGN+9WP2C21VhcGxc9y4eLV1QH/nZE/7DYyJ3B5/uKX
RMZAfl/2/O29voedYxt5/yDxnNA6kTJLUXDcaSDvAoyiTT8di3//bFwmnRrkqp3d
NYMGEhDXcITlTE4qadiQrDs3H9DGTp+FsI0ksjEnO1XarAjgAZMatdYodPrNH6NS
RgAK1oHcAJOcWidCZM/5Tdsu8QRYf/S0mqxjAHG/I7BVczR2IWjNex49Exc2k1ts
KNtWD/SwskPSJyxrYlxGGSFFWamk1+2/46gD2XrfM+P3QFkqcpBlCnY4KEKJJCFI
JnkNY6Yc0X9iIsEEid3t9sEK+Ye6LP/0C1kVFYL+UzoxlpyMoW9I4E3C2eEdCLnQ
GxY5U959aQdrYFU11YZ4KhV4qRB7r8iwDERITTjdHYJL/XRAJhH+wxmy+p5UgGJ7
ueI6L6HKVcXzsFMkCMXaP/OAWDVNLlUdogfa6tpVw+qqOKwezg5hP20nTr++wVAk
mrvn0XKxi9xoOUlyArYye5KadvDd0RRU6b+YH5sFjW7nD5BWOU6is07T7I/GT677
J0VgQYJrk5XhGFInhpUE74A6Z7qHV7aPl3rGmphx4PIBEkmmXojTsGJ58BAFiPqW
RL2RDO41fu8gH6gPc4GNfcVJeVnAEzLec1ZI1y5w6QI68TyHA0J6qTh2kJsR02WF
r0CX+GXiI2BS2JfdzN/HsuL2L0P66GUqe9MktGu5hrAk7FP1JIrhZfxK9dKMVgo7
KBBQGyjq+rx/N6ryvZlg5bHPoS0sA2Kk0rEv0K4O7nWhEoU+UJ2/tSgNF2PafJE6
DTy6UX6nz1Gt1tpCsQwStHJweRyluOD2nOnY55wSNOLA7UX6Zqfpg90JhM9ilrU6
JatIQe0w2AP/ywiRdU4HqPWmsXxhgE4rPzEUvjmIwxmDKvjmeTnNr/JBzQDGh1A/
en+X2QeTEhEBy7m4H5nTzUdACtmcEyYIVlhgGeV65nDzArwFxdHt5K8ljzhTIWif
5nmAHXxIeQQFEVueBDVamAu4HGBBlmjJBoMnzF2cZRuMOJXCBiItU/foW8szjJN5
JFfk6edOReHq5JtVmD6zxdrOPbr6t0ymHvGyd/p25gRG7g4KyDt7h8Rn3KPpA+P9
vFUdK4YW4wqwC9hfh4tZkqPwrlaMG4mug80PzrJ13nCT70IdKe5d/GXI805aTTeG
XNFrW9292dTiI1lZ1r2LK+r69y1vcv3nMUNoewc4M6qOizFKxTitOUPjJubsbmqw
jZMh0c9+03jG9T5srvTA+wrwp9LNhzUISA1rJTMpzAvP5gUi8cYlS99sl4xflu/h
EPH6XIiKdPTshR4z2hRYnII4rfL/s2dTktiruk6bF9sSnIwhld8Y+aRMs7SumxIL
qpJ6g5cOeL2XsJa3fed4GhqjnFSmZHrlbeRzBcBr/Aj+KcacifGNE0YttPtg1jkE
bycoowRb5pLMlNqXMd4Ht4cKkbIpgB6XDfn/OF27vW0qkf/HRmWONfmd8p2ltGKg
7EAh8aX5rIXR7V/knRBznxXvd1lgCFovYPAJgYCA+NXPk6ysmnPFPRod0OCeeFIx
3jPVky/CV6YEWVd/e+42BLYVmnUVuhnL0fF2b4df2fVjjEBf4zYiEXyLYEpPIKcn
idUTQrNVHvq/yw4kyiCtgsAzHqlHlP84LYYWnNCdeHS5yAS7AIIGONI5FuKAjihm
pCGPBh9P/WLWoDUdtIJzWCqwS1aZ7G7gC9ac4eioGWInLS2VeIoaIu6/ns2VSYPL
ZV1I5iFGGrhzIx7q0TsLF0BIdNdeYpv/KyWf7TVf9Bo8lZZ3mfl3U9Po7rdJKSLe
2RQFK/Kx6gaCXrS7LlkLihPV1N61OMh/WHs9RAQHSTlAOK7rAYXPo+bB/Tmi7SYl
dQdrhuthZggt3BxfEZKQ6vu2sLcxp+ge2L1MpS+V+RoPHeoEpLfQ1NN5jgvwklrK
DlrTjOLErhdiiX5wDfP2AsJimyqxKmVaXLRnABpZYgaWy6TM2hQ1Xi2cXdqujVnV
0lnNDuZRET0vZ93zjRd9sFBb7OBjAwQF0v47GrFTA9/mLDvtVuJqGgSQqhOqCoxg
QIKKagGZ/7yu9Ps8eA045ULXsd8bT0wBfU21zDRYmLF2k5nqltCgZiDKQVkl/6rD
CELnv9WvYFC58ovSufZC3sv2tbBnOoDwKC3qQ0TcIfRa5iO39XJO6z3IeyBu/j6h
M+vaZXDkrterVxlUytJNibdKSXHYUnW+ftnFJbsp3sz5jEEGz83F1SHR/8OQlyx5
C22XyDQvH2vab2+cMt0pwYxJO8XJqJVb5RxJ0KZniDRyiPJi8S5XdoBg3jXqPdlh
Xz8sCSNKehtwDRWSk27TZXjM2wC8+Gd3/q0MDcUXHjLwO4178vrFQuT+P1NaO4Ww
KpXEOBiRGC/loK11CZSHAz86NJzgP2yUd2Q6DnYhh/m2Sm9RJ6pJQrZi9MYTeBrs
krJF88dSg/ptD5jcp/vs2oI6IHwUfXck0ybHux3B+8ZocvEn6MzcBUiLPJ1WTcH7
fLLqVx8usg2bMFdb6LfiQo4grturO7bOISP5rytkZZs5cPtTlIkitbQTN6pjQaO7
8WljJGUFHD7LzZQyCDLLNVDksd4t832/jX4dz8SwM3WcI9lh3Vy88+1IOv7Rh5wT
4Y2KM35iFhx6wexix/sZuAgeksgcS3hUEdmXbDCTbrdfbZGw1BBSV3eHnhO2eQ0S
9AmGaDrF1aHhwe37z39gSTYqXmoX/0VCfd9skQXyrpGBrO/0uv+2xuetYuTjyPDZ
LRQ9mB+tbF3bwRJaQ2J96zaLt8DT7t6Vpdb/ltVG0/hvKeBKvLRdytflpuG3Tji/
2Mgzyk6Mna6D9H1gxr9Ay99jtXqLWQynlddG1RLmmUmMiidVfdtOlpvJpeS7HM2y
spSxeb5mCNUDr/c0ViCjMbrqxNnH7hWXQzavLEZRC/vTCZR8wZpkCPqUvjuSM6A7
v0v+9TOPt4veNqyAOIYWcGqui2c3sDzg4ZF77sRCC89JNr46eMjCW7qehwjGnxxM
KlE9a7md81dgqtZpwTbkPvD/05ddUBs+yzE/USVMgolWLBAnKKHr98DGVuw5wFqh
M5PbGYBdMhUNC1i51qPLLt95doHa1JzcbgnuG7VCgVZ0Tj1dJRX6o/ed3h5WEn1C
smWQ+oFBYikO0Hi5emjCx1DVpyPHQeEE59AqH/KczVRqOcl44Sq3Ft8LVvQmx4d/
me+kuTde+WWRm+o1/hI8rdrYbhT5tcKqs+jYW/1xOhRLrxujTpP0c1wyN/4OIKDA
1ZjkrypeKgkY/E8bZ9j8Hywar1RqjfEgAwrWNW2AlY8Q9j7DfAgkzfrj2cKzPDMf
XVbbN0L3CLdS/EZOHQE2QyWU96yAW9I0/XmPaWaeLMTlXi0Nac4+NABlI31+qVpH
TS6TbQ9Uoo7Mh/B8PfZKrBaH0cT+MPPMX3jepAiX1VpmSbOkUPDS7gOaWfclrjqZ
3SEP0gE27ZdPHGhXMWRFTobscpE5ENpVKOXrcZqB5zI22kp98+lGiojpOxzDQPR+
J02H9v1so1NJEh3zFB5SjaJw5iGaI8ZaDQhBIAM5MGWFx+ut6fWkhxemJ+cWn8Ha
xK6aEd8wiJwox+DJxNC2FHbbVg1axFK7NUqyOKPSirtW7bIMhe8gMLmdYIIqxwXm
Hcn/c9/J6MjEFv1ofHXprB9PZ0/vhaKxSFYV4y/5UoF7r43cowgoKk9tDIK9UzN/
5yCGDoZgP8qNfuuIchakcKhdvh/xOB0bmNBSMDyHLcgGEykUE5/JcRONMC+b43wx
7Vizb6Kpur+/89Punf83hy46Itj1i4ssn4n4achFg4vqVztzCfU9kaLfyQdkuqrm
uNOMvUF/ldUGlc4SMYgka7sWpPKRh5B8hulxEOdqUuB/HvbWtujrLGqLXBydgdUQ
GHShr/Czmo8aTtdhDgXOjPAITe47WCnc3xIoKAhEC3bE2syQhn3QorhjuQvylJTK
uQM4Vum5uJVJXOLutSMOboPpb2ws4vTkNAhidAtvV0rnskYdEWZh1gULE8HQGbUN
RaW1y/ZyaJveBvGM6BPotOGrEGckQvqkPTzWznsIbEzIm0DcrLkUidlg70azOQ8F
JQeOMvNVWvRL7hLs6kxt7T0POiTOGMIT0VtyJsvSuvZs4M5j2ECrNKMdVDXAOatl
LKah/647qG9sxPvcRq8l5hLwAgVf4oFcztKGoEERVYdcBfdP0rF5m4HqytLs6aau
pt+XesOir/CtkWtFMzm3NS8CIohSf3jr6rzGCTgcMJLdDZmUlJIWTEzQQ+0GFaSz
kWMpJ13o208k+J1eXdmmXzRMNAPGPoveriHMr05c10X970EC+rhozfWwBkSWHNPf
81SdyVrj2/sfIsKUxhH8MV0CwZPwql9T5hrYytldDFJ7/7J60YAeBHAVWBgD5Prj
LAwhkJ/jSCuHjbMhs/Tz+VGascHiqvP5CANLhIvYvz48ebnthG/ZSLlDC7R06j4i
stx1q0V0fiMH/mpygtAyKI2oUWDL9Pt77HKTmRKToMjcCH1EL17Einx7iECGYu9k
ZgXv4zIflmj69mr3VmmYNeOgABfltEwlo9EKpNmhvTJaBYhFGJtzEo+vk+6xpNuo
epAwzMpqFne3Y2YtcYeSF0UW3gEhuhRcgGtRiigmymtYhBtBQ8mpXnJmgksPyoQi
JNG2qtjZRWCWvEETPgBvhzm/D5ciWzVzvLUaHQe9sNbRJO+HXCq6HJzDOTCZRRHs
HumDgQbdyK2zXcADp5h32M0QF065nT48i+2ynzjbhE7Cs2lIxCuAyX53X4dNLlM4
8BGbI42x3HNGPHZCcbdNZO1ewJDJP6AZOzZvkpUlalH2d+UFz0xo5Rr6ckOySzdw
FswtSRD4KBzU9xS2TPm+6iEEdew8RXJchPmvqCGz9Wu6mBQiALcI+WfPBynVXBBj
irMoBLZM1cdLROWX+HDRHW4ShebRxjXQKdKwPyo3/RJloIjdj6SZccpHz6Myvv81
CdecPkLUVSWzlOgJ4lD5H0alPCT0FGhFvH9iDCDbnY7iCCDnAeBdUj/m1nHMOH8A
xwIuL1Y1Zvi7cQtSvVAj13WIV8xxvu/iD9sTVzNyL5vtm1D+08xr8Sg1Q8hSMfdU
UuT9aUAekk9ULVMF4J4Xzgd4DAnaGvSCG2YGjjLInXdhGDOccYI8h9rT3Kl8eL3U
1FqzXzvHpYsmeYravghIXDqhLuxkAVq6a/zuKnHCLn4l5+QObmG+pQmwocFtKJpG
fSIIK46je07imwhP76rqbpcx4MYJxlvgDvmde0BvW0y6GD/rUxTSZfZMLgx/7rGR
kmY2z4V4v8LUGwA7hyWkQ1lZpQ7foup8kYyDs55OgJYrb0ermNmmldgeM6/b5rdN
/+xZIrxWB5uNInLGUQ28TgieSpYvkAEE4NZGZs85AsFCdH7jwW3MuPwEgS6fd2bK
t15bYEzGjaMazg1PJ/TFnuzBUmA4CT/CdGAdbNE3EA62ZWyEmfmx5H/IZPlfSBZC
OWb9DWCCUCDO+I0CfBz7W/fffECiKXHp3kXbsDLBrNTiiCO/yZboTm1Fao5p1xCO
DcVl/YXOss85ED4nqbn1q73WhXnY86FIMb01a//UmHzMGqLTwd97fhcbTq+zul5J
gkTugcgdzSzUne6DT7rSr0eZZT8Qf8B2k07cNy4RwL8g+3C0yLp72F+AdR3exg1/
eHDperluirvwilB82vugXfUZP6MtIhM+EG6mQ76STGhm8LDTKmHZ53RhJkHMiWum
BgfP1ty0+6Uh5qf2uiqxKjD85XPeU7tkb1YZs9NvIjMnOsABsF77kwXSiQNosJz7
L+WetzA4s52wrVPd0uG7VogkhVh9IrFGlibXwx3og8uhh0Rqu+4I5uo3oGSDwhuV
Z9+gHOHeasUhVBCgcuqX7zcI62idx40/RYlBGZfmoMEYvsUnFM5YNPf+JnZ/MAVl
RW1M4btzz8ljApJG4pg9SFM/9fu/gqkxL9PMD9fPutwuJai/oQ4Cs0bvQz0MInQ+
JO/2hvpbz92J9CzRH1J8dfWnogrioer6xU9Rr3cRbqYzp8aeVQ097BMxf60ZoVSz
0p9hGIF3iQ3/7osVQxTmKKKcOHyyTOP224vzGrIPmgHp0Y1g7t1FvSD4Yez1YEif
KHBBoZK60TGBC01zeZmAQ8coGwjRL3ZmmNtzHhbJ/4BKlIvoNYvMBctdbECdG0hw
8o0rDub0RX00i1JczOtF/yStvuUVIk4dByJBHSGjSnf8NgdSI5lN3oeRA75kexwy
2XA39f2S/6PYDJpPbYATGS2rD5U24hJVXcmURUX8yqs9OkhKv7/s7Xfo/ck78/83
/b7lV1kpaMlX9S0V0HaB1hrAp1gzgCQp32eq5rqF82a/ulwUDSUqwrmZ+js/fGnv
e1Ye+ZIbBube3EPhn5qk+9KpBp56VDAtaEb0dImjVjUZhqmtRUHxFA23XRci9zAR
w71uM8DqO2/hYjapmytQoKK/a9qBWCElpuKHYftShirzXQkBfInOq+VhSTWCAbv1
FTMDASsAdwROOn/8gpOSEn1z3dUiIJRTfOJJX8Ec8FFAajcPHCMNs39toI6F5uhn
a6DDGXHQjV7d2EAcV5hdkjMf/sBPpX1U0ZcdbdaTidh73ILV/ycq+7DPwfgu5SYv
JtglUJJlb3htZgzsY/SwKvw9P5styaGx+82TDjlUrTo6PGwbiqWiIuwdLUJEziQP
4i6tZGx0n7F64gjdhoN71um+2au/bU5m2Cwp0pdsymW1TY9RfMG2fc32agZiF9x9
JYZDQYjz78JIOSNLLousccdeD92tQwlsAF//inDFe0gDAP/vtTTe6yGLNxEfFBbJ
lUfzZcsa4679RFeUdIut3Na+P04OWuYBT1nb4ut2NSXoIvEG29Wx2c0C+9imzEtI
CDsSv1L01kiT80cICRBU196aOxt9pqShHBUz9aQ3vMmFo3qAQMX1r2vIVuGqJmAM
N2+rmLJsFSTTfGQKdr02ioKAJazTxc31g3utOBRSwB6nn2AhYc+mV5QywmESHDvh
bVtttgENOjZ63viUJXO5XFmT0JOnaJoMyipbhLvJDQ9BcSRFAVMY7A7ECBaPuIn3
zA6P/5y+/gImRmcAXfzbkWV9Kjg21JSG+bN3pN3Lye97lnXZAzsxwoR5XvBbz9RW
i+37CDE/1aP3HsC3BPgoTS3wMcXbqv5+SfqylX2Gfz8HUVL5/6oO8xQOO15wbJbn
Sm8rNwzJg1KZY0dqiWgGJE/WZz0xtZQUu27adKl8xhUpDhb0Pc8AwxfrJmDX84fh
jT10EXt0c8QpBb62P+7sMZMoXUOeq51AC45Ogg++gsDb2tGdIq2OhgXbXHVTAUCt
I1LK5/iuQ9drt6yBK1haidVxoX2Drn7qX2wBrm024hg8u3sEgOXqvacEh7s5Joew
vTqEDV0Xh4VoLzZ+viikP3OCAgha4fJNOzfKkD+o7qk3U7fEWUYv5GBb3RIErPdD
wn/6JSqflMknecB76VD2aDU+vGtPnEv61AixDBedFHr79RsOFIzxAt8eu+q2xId4
5+iq67bbK8BHseoIu5YGZ3Ev3/eukH9sOYlINfizKC1p9IzzZqKShbGzmeC2K8BG
0J1YDRDT59bmARVrX8J57u4j3V/oIxjYWWnNsyUuc1h1UhoBmo9XDbllGiIpHZiH
KwF4QISbB/btlui9j9iq/NhTaFW+M0IHftg7p50dCLQoL4hDJSbO/zt8ba8h+7un
wIaVa4BimX8nfOVDgGM9PeDgbB22pGeg78UucDHQa3z3y+n9g25NOfR1DBof0O4l
IZw5aRLCjSFw7Z26hVgHeGISXJKZBFfYWnfNaxAXYVasTDQ/e2dPwczvrctjgWj/
p1qorYFsiHzO8c3PH9w6StqMoEhuX1B3LfYeenoG58cLNiqoWp7WPLJhc21Ft22/
hEG88zASFuUqyhwXEzkilRPZPPgJprqajnbHKiTMDSAKSWvWQct1J2h7k4g367WM
0vsakeENPVIo3sFquTFEEwm9GC+RzmfxVX6rknjPHSA/8xvsvNWd2awknoHwUoQa
w7J/6t5+mz05MpkhOyjadTqNWDrKsOZO7u+EJdNo2C4j5EdLwT56tkIJVNUFn0rE
lpdvmplo1fjPtL5gt5IrCytm2PvFKrl+t0kWCdaliofLkh4copeV/GG5DTdL6dvF
NBv+7JYziff1onRlgodRZbuP3Z/mHTHz/44FzOdA1J9E0A+5MTE+5AmtgttExKWz
k/mgvyW2M9SrPJn2Z4xLOQEvD8hec0D2Bwl8VP91LMtVbs2Ur20i6M+ZIY+800Es
8zuJK2hwRK73EnMs/zsf+WkQ+c0+AwhxvFbG9FDHh3HI/Sad9ey4jZpAKnQJFMTA
2YVdKMrv6TY8bVxHai9MCXKybSXncY9iwhUaCo0KobPOthfQLVInGZ4J4ickW+HN
+LtVk1uzdIkz/p06985PPyrnb/7fP/ly6/8bQKYoTnpwUoByeynmRD83A3rNZ1u9
pfFWXdwa4Rf9KJWEjU6FDPEl/RwilvM6sldh+4bfHBBCkgE5FQelvZ8l3KM89xXU
1CEiW/vSh8rA7vokWXgkIfYFYEar1JVRrKeo2+oxVkowofk4S6OngXLNr2An5x5p
Esvk2EeXA+xA/meD2ahmHpepXdiUgkAQThGhiAJgNe4DHKW47ZCjPHBeiL1r1NcN
9vfJzsvhZ/fnoaOVaXS18yrRbvVQXuTWboOeQ1Dt+WjBwGnr03cPAQxKCNibq8rF
5XO/oDbfKzl0GpPONurxPw5HcNzlIHy0sMzf52qXgfb27EBOYJaAASGnJ/7dwoe0
seQs/jLvjy0+YlsNZV/A8uNfozTbyJ713bNJdcOaQ+cDAU5L5jQUM0ImtJ5xXmHC
JCQ6IGHZs4FdZRgIFxfYE2waQBBKZEieHfh8Uw7zaxBR7lLMYM0vbDNX0F7iJzYN
mMP4R9CgJzKvBnm+LS1kLoOas6FKvvP261dnxasqzcScT87jcMBBaLvYzl8XAQ9d
Je7JbPzirn1ygivPn4z7OUZJ+zYB81W3NmxmzOicyNhL1YA7g8fOjSRExth7mSVm
N0V+VQYtx8KOzBwhmAIhtQJeFex2tDNWTtj/PIg20SqATrhUW1IAAT3CktNrMEVn
y/DBKbbBFvGUVV/s9CF7f0A6UIEz4PXRRYwDPRzD84DWlUngaedieBX/2E8Je5oO
dPqo/axYzgaAl9S0q/b6SLn82TvfwWueM/9i8k/xgNJbfdjjWxoFZqMihWOL++jR
iX5ac0ei1a4+iGFy1ooDI3M0SCDtQKVKKpQ8IABj/fK/UYEsVb6s3sk+uTwA850T
34bPrCN63bmCCt2tCnDK78goY2Mcy8FIB24suD4R2g8aFsnyeAkcKAna4ErQiK7j
jtmmQFcp7OfoiQcG/xVyL0qdVrvwsrEpFVQjOcnk7BEXPlW1dQrNXbr0WTDyoC/I
opMTCZ9CzpAqhE8oN4XhH1mhC3PxDa6lV/x8dHRO/8HjKqxCpt97lMyzqqzIYd6Z
CTht6hW5GtC7LY87DHIic0JZs1VpmgETTuYSq8NwmRPXE45bD++KFxUut/rvd2l2
NYB7ZNrJzT1oWIk46NqZ3eN1DY+VzwoZVmUrHhBLYyBJZ2Q9rzsounJ5+Bcwqy4S
+TsWtawF8Q0qQ8tuMn1tuyh4l8WyB0sqS1P/ziUodr65qCIMiYJox5WpLLD0nwAz
`pragma protect end_protected
