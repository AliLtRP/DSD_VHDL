// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gOiDMjW5HYlYHVphdJhnj5j+jadpQ/URFUynIMZRxZ5lCrqlXeO38muhsZCOC7XG
ObVpPmDqo3KzpGWQGGmCni+RO33j32aIMgHI+hyHa6nCy8uX7tRNIaMYY0T4IVVh
JgBdO1hFIwM8OGSrbfRbXu9cR5hoYq49ooBaXxkYghg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22352)
Kv5V95bgiOYpbii2wqNgVCbiPQRNFD1kXjDyXl8eJOeoGDiJjvNvvSS7KmIjaJx5
ws77NU+ZVwOFjOqt16k+xipPBykZ8HMNCEt2NOQETDo40FOZJUUDkCyT+HIVgszK
JGLi+ZDoYix3O2hIUMr2L2L9GUOYbFAt7pH5bma59YjlvP/DjToZKK0vCnLoUFlp
rhLvmZun9AV8bhxOdBlu9BGxg5eadoTVQHW0pWChIGZLPtP24exIK7ZXp7cP/aN8
x+9LnwtMns/YOKIxh1PPs72s6yFpMQn7Vv8GyIC5ti3u4vEdDA5k1CtubAuWI+d4
L5ASeuTwl/jOrRsOyKfDCO6NWCYEhZKzRCeM2jkA7rZQoK/+dClA9tTVIlN/q81/
cXh2Lg2iX1JMpsyDp3u/peyhvznqnedxU0JTWAh6IMPaNM/vUBH637Mx7W0u1aBI
CS7Cr7kQR4l9Q402v4vCYGk5rfphEjcFtT/Yl+8yd9qoez0uvvbTPt+sikZAdRRl
bo9SaT+rE0LruzsTDK6t9syQltIRx89Ff7CXxEITcVOf0MrfwmG+LKH28mmDtWlF
fGVqDCm2F0kFSosvTY6eajOZrEEd734nk3v1FRYoBIyCvTzTsrGMkIWVcghPC/5A
WESWaeLHyjFAd3P+5VBBKw6tfx+SzLFbjGCd88p258ONvxtDWhzTJw7icSrzgVSu
bguHdJlv8rgzr3vr2yfInqxAIILhrXvEsv6TJvbbOwaN3O4OOfTtOn6zvMP/P1rH
aPnlMIaYJ+gQBxUJhRuqChfZTWAwofdZQJMxOaSMH7wixr9YIqIsYobdAGAhJjn8
fFGUae08wmI8VuI8TC06cc/WYR67IGoywWHPwVQodoBXHAdMtIBhL/gIOgpHc58U
05otnwbqv+SdbsEbOxZu6dWMdH3PMhMAx478HIC4CQKKy89WT9Iv0gF2SpLBBMR0
D7BB7n1S8lPZMNCcw8NWYzT2sjJYD3coEavOmtQtPX0lBVQPAHp1GkXSjx8a8zla
qXhUdf9TPnmYcVYPrTaq6zR+f7WrExB9OkEjzfYqKDh2fZqcBENowZvhDUcNlMgk
IkQ36Go7xPQuFSTXo6NrG+EVtGBtEavL4UxIzuNuipWs0y4iXQxN1XG3JVQGF9wx
nh5Dy/xzn4cOWT/LppBuvOKfmoXNTb/gdGhxbppWd7ZZjOFZ6e9W3mEVZ/ypnDMp
65H9jyTqMvkymY4xV/uq1VXAh+khD8jUiHFgX5VaCJknrFe1bdOK6TMPDFdjGSLI
+qxaI7RndXYExnQEf4+J+lcbn/TMrlR/Zh0feh9QNGQw1s+8JsmSSgBuGZHNCsdK
Ul4i7pJPPhxXRldFUC4ZHHjFap2g9Fc3CuoTwgrWMh5Dsz2chGhJpYRqves9FSWC
08MsS4p0h/UZ8OqwfJFvN+mByFjITe7dTxHS+zxMpyqRKLMMSkjRCj6vqfAiBQ2/
KCXjeym58Jm9TFz8ZkrhOAHbisaG3D0pnzpjNqVUX+6QUDudrsB3yVsGPg+MsaD9
zXc0ZZpdRWqpQlH9Wf9Gb6dLthXDNoRTHZ5cK618VBsmYTWAN36b1uGXQAW8Yteb
sDg/H4R7MD478d7733M2pfW58p928rz3UZDDlc+kxkhAEP/7qs9nvgJM71MQ0XMp
asQ7StQiJkt9iSL7WqUwgOSZjMYZ8mBNRfflEiFejfBsmMlwXGTdT2w42Z21apLT
wnkOUaDkQpjbbA71IIRzl3Acfb+fWSLFxzDRRE6eQVPhzgx2nDNsGoQrctgauNoy
Tb3EugleLOWUVC2iD9tI6Qips5jGjvczbg6a+JM7pMZXjNXSk+RXHukYSUHJ06H5
BybGkN4kkzHiYee4m9Zu04DC32OV8STsaJ0i7Gl+13dqu0oNUYutP2OwjC+DASFo
nS6PpNIXwdhCR/FhHbBQNHN7bkouEXb93xciKxfDROkp5AoeMbAGVd0oSLYcslKN
nSrOzJAO8asktMB79Sir1hNmS83+PNsEkrI0ZMhBb4zRrEEasS/Dy5gieB3PHZhP
yvj8/rFMH9A4rtFMpROM1e6eXlBk4D9nLbb5c070upRyzPcFp8nQJtYJf+HbBil5
Oegtjx0MtI8ZPAF9wmx5c3qs3P1kuNfoZfZ06wuGm00ZE/wNbORolrzJX4OW60V6
kxX4Ialn7HvlsmLULEHit+wDIlRpOC6pfL3wiHt5Cv0jvHB3IqHVy9t22AZUeJq+
UfSfb/+/G5GiHKpdvsGyObdvRpuaFkfBtNrpuJyEGTMiAsvnng+waeZKGda9DgBd
UPQ6vQMrG72Seesk0pIoAJw/kQSf9ttF9oihG/L4EBJM/dmZedwYTBc4iPJ8dNcb
OrR4ANjE1xYi1ONKMrrWn4ZZna01wk2spjl14tuqMyLLsrZFaHDFYKFXSErn2vVx
X0wYLAQKXB4NQWG+0nH4USumbpNcASvptSaz66UUZUg2SxwbAdVE3WNjs7JitaU8
6h91TwW/Y43iXrvnaL3VPvQJrS79Q2dpGfR2cA3oaO4ei3Z+ALkNi8cPKwD7ZflL
tHKgEBulveKdxICoedVNig4t5OMNPL15MMknAS+FCwLAWUndvbJ7/zwbdRlNqXMd
Z3s7/4zDtDhvLx5ufYKxH6un3G7RLuyMddKFtdi+aZbRf4ZqAhOjtFUSv/Vqn2Ft
878vd/r8qpAk1mTTtiK84B8lFG59X4ApCkcn/f2ljO5sJ+NP1ku1M6yHI139tseQ
M9606/ZvUGAAVfRaoX05tN5ixs0CZdsq9ig4/GNbhzMjQTFjEezNvN1sz9iD5FNj
cIHZKJcqebuh0PnSbre6XL0a8y9nobPM3AkL4SNDGVYWBc3iHWeNQ1oRTOAhYYrL
nDVNGcpGdZnqAugimgF4ZIWJ6+nf7XC5kVQXrjHHp0Us3rZ8sqATXn00geqami2r
gpalzv1j1S7v0T41ABNJlQaw7690o7qYsRUVP6O5XK3aB4A1ZA+wi5iVpBmUEzKo
n0wgLVsUfuOK/Ouv2yvlYhXaPO7OEz4c9l9FSwiZYRMPpbTBJx7e39gwNZLzJ0fL
4IBypdXrkS3Sc1m4HlBdGgmW6aR3vdJzj8l5MPva9fDM19O/hjUSOSkn75DON3aY
GBwTKv2lHlwgGmDkQGz/KypSeJEAtZEAw82lka/2cT3UeFh0NaeZXH5Zl9alYtsf
Di8L84zuqQDdLy4hILDbXv31SL0ikOVqvQdCyHD20SbZ/mYtbbkMOky9AjQvV0TL
AVm9k7ps8FmH3YbfqSoXKhHXmROKZpe+ekwas+pHcvOOqeKBUnO/u1B9QfZtM/SE
NiMDAQm07ooIvEr5C+dUE2SJlogGg+v8J5s3Rna3IkVNawvkKmkPrJrBQs8CiGbm
thHPBu70A/i6yE/2WzNX5e9P0FrAkAld8CYk7+hTJ06SuCIc8Vj1dX0BT7vqVhp+
RAnAvB6Y/hS3vzzZ1YvQRtBLAyjVhTlUCxv9UxacNrl9FaSgB+TtAVwph2U0nkiS
vNbpREV2Z+QoHTdFeav4O7FwR31oALQ22j8D4j6FnkxeCymHsG+AXKOEjNutfxi0
ANwcR8adsr5G4I65Tw3k+E6d5YdJC28AK0WOeAK68amR9HvMVdWF/TjVMPPIgln4
28hq5d5aaAYy7Z698oKgmvs5gCX/atVisQlq2/swQD2cIhWn0HYz1MCh1uYQLwFC
UFhUPapz0N7MFQgp60GltyY+OjmU1ao/Tgic0ZAxF6yfpKpoOrD/ka/1t3Q3ojyU
xhGldY/AeL5HV1lrYb1VXf1oNAwjNQCp135Y9opbcyHF1YK2Rac6ryrPCkEBK5oz
oIR9f6hNhkjA96GzP7AgcersUw9VC1Yc/v84D8ShCXjPisdiwbhLNS23IX4AQX3H
6AzoIyI/nKCZcfaNrLzel7Zte/YL6hxiRrwVlJOu9GcWbeFUWRt26dX0DQsUc38C
iamuFwG2dyE3UddlmxAk7wOb+KlKmYyq2F6raYIBRiIoTvRqygM2WKWRcL2gyqhd
B7s+2hLbhQYBOYABGQRa65Z3yUhwq4tUCxZL1b0PL60gjxEgBt2LRpY9kgzkQNun
1Gi/wPaJiaRK5CvbvJ8cCTtpfiAfONRvW1nbSbzVyJv+DpKNeYZRMcnU25tEYeQ6
KOSfBEn7fB9h2mzqBjtf7F6WwJJ9RourYuCm1bifq25xGQ+jkVhSskI98uC7gRJ1
BgzRNWUyWjJ2Rl1VThtiB7y0yg3lWRSsQkF7CsS4T0mG3UfF4AEThmfJjzK+FIOO
y42wT1F7CCU1urHCeo/sOlSE1KHh5GcFlshCX04UJIkiQOGzIbJq9YC2eQQtwyUT
QlJvQQd8yjb0O/EWi2Pk7esGpd7R1/U0RziEy3AeVFGA+2UjgXdBUQlUNLclV8OY
611VPq7ZrhqCzogZ++aJ/mNkTQtqmE/Uh3p12aRESEbAyr7pxxNpweD/DCNiY4P+
bd4ZeJih1rHL6QwZgNRojr25yeVtfQGwygFHCFDU/KhN1ADJ/CyYYxY/EggG4iut
V6uD5BFs96BjQwj6xDdJPI+rzFjdgrQrwVTEjyKVLCL0NVTRPMLBVGGAbksgExW7
DHKIz3+7Jq/yyzY/PFUnBTNtMSCAsAn8pmRajZ7AJBY9pCXYQwdvx0XZNotlj5Jp
KLcUDfbTqPw5AUwPpe5LXz8ELlTaK1Pgd5X+w3Lzb7kxh6/O9LkNng5AvxB/ZwGW
P1dpysH1XCdI7/QqY0kT7E6ePwRVeJopKucW0FQQGLV14ghCWR7+bTYzr123wMKU
udB76f7EdsgXyWuut+i+Ln/3xWD3i9JSB1ycsNNQP7GN/O0g9w5J6k6d9HCI5qsw
1THk7iNcLgFq9mKw/ogoyUvgXMFh8jDMZqyjLnFZABng82MVbtIRShfZL+Gvf7ex
LSNRsghe3X5kx57ovufWjd3vnvsAUEXywdCdOcoOGcjOLmvGr61ao7KCqntFkyKm
XmPBm5/A70IjHZ98yBf1XXuvitnS9QlA4US6JXMMLCAyn2Wzbl80qK14fzaAkMxu
YP4bIuiDJKB7x1wN8W2RvE6RJMWEZEyZKhQO/N3i6p3FYQnAKorCWgm/PltFom7e
k2lt8RJYNefRU4ihffOhRk0PMwjRvdeI+lIgtXZ5OCG6hOtR37lSCZxdvWohnfi1
iwh5DTFX/ITksu9zZPuSlho9ZYbhCDd4zxkwZBZDM3U8rY9D+uGl558KJVRsjIUe
pg+Pqr2OgrJg0tx1rRimcPcnemecuUy2vmyiN7liYpmcyUbypm1rGUmLC8heSNng
Y3VSqTI8dd9E57ZD2rsWZYMJ+GKXyIs4lXO+wLMMTJD0qSs/Dqaag0lSM9GCkOLI
W3iOEcDEeLDBuQ6Aa0Ot2BRYXRq7vDlt8VEin9xVmWXBPradvsSNLyFS60nnoizE
z2N96+/lGlKY4rxqlpuPTlptk2n34bhmNR4HeTGA9FXtc4d2AZ4bihv53w/SsWyy
Hbsh7BJ1hqHrrYsC6jj2uDp/VM2a+zPUxZGyP18OJY5LphsyUajPX6ipjyRfj4sQ
HAPBvhf1jpbuX03/Jm7XisXa3BfT4kyiSkUiTuf5LlsR+6H8hsp/6l8OPsBORFXW
1fURBUq/eYifa9qG+doon+zlwcvXFVFKTUJgVV1qNK8AeNUlhNZsmyoc1MmjwA+P
DZXOal6y4P7zVaotGR7XIP3zWfskyHiFmnWjpfqSmDlseS4F7hfpC7PiHd68CoqA
wXRF5HNyJqplISMvq2nN0yInhcem8gl+LLoKVEjh8lfA3RdhGJpX71S8MgXRUUxa
GQV8izY9sxt4jAz6dzErjDDri+xhERI4DIBumA05HTTttdDMijXuKhnQK2997nX0
VvhK2aVdLwVGupbclmQChdZIYaSfhMmk+0XeZRnJ7JErUOQF/nbSDqBhNr9pR/x9
KuMuBHVs/jwW93MknBjD8Gs0o3g8k+5+O97coxcZhiMuTvjH9qCqsumbiZhkmIi5
pbcLoI+tm8ttclECmdv6TFtQMUZdR8oN8HSkNP7az/QqxDhzKplXzp9uOoNJJgtw
m87Mq207h6NGXxh0w6jTRsgTVUTzbr9ASecOCcQ3rT0Ql9tq2IP9x7+ftvVb7SkD
hSiw16X73Aw/uNbkE1VM/AhN3s8BPaHQtZbKoht5pvvEcCA/gPCQQZcCgEw6aysE
LtLAObKAS7vc+sqpsAVRbuuPNEoeQFnXNDNwS+ZS9tveWZ1Tyowv1r27mYPShfLS
k3HhQzSYx7lCUyEIBt8BFEAUJGVSpjF8RS4gBYOoSi1EqLgeh2ZPNc6v34DadKck
MOmmiKoNX4eb2tsKqkUAt1b0fD/sNLHciQcTbIFQu1nfIuqLynIKYfcB4VSGSIS2
iXqbZZw3wAXwUUklV/ddi5KbMiwi7/QRndQvNDH7cDPJEU7UpzO5b5uyGbeIpSW8
AkHEbfJ1h9JwciQuevROrX1felwmpL7jdaZK8WuX74M00JuIRZJtEJbhTlSg6+Ge
HiBT4Pz2UG/LwiKFx62EZtRrL65cAT97OT6VXiplx1X10f0c9LTxdy6gAiKYi7Hz
XMznGJB9f4mQmf9Tj1FGizXWFDriC6C9HzcBYF5usUJAUv6gWJKxRf/Iepznm2yX
M6tMmsNnby9YrH9ld6J/bNTt+aEICHb+QNd4cELoEs3BRecpkqk5ZmW7oLH/9dkq
o1QAI0oWXpBYTgnugz3RICPynXn97OGKpkC2o1d6jOhHuGTY9XQ3SliN3SrHhVMG
l0KW2uOnviOg9HX+iO4/2Sx7ykJyeOVNgs5YwdIbmA8lT6jKuuxDaLgO0wnZmGLv
DHh8sHqYoGNdVlb+PXTY7N2eJzDTU4uTvhCe+UQm9XsOwYfo6bXGbYzFZqoKnSgY
RU96o+GU9zNy81qDU/OHf+7Cwvd5mFkl+iMh5bGkin+BibeiSh9gkl7arCPfIfUQ
AyQNtFog+mQUrh1by1PPnF48Ra3DuSvqWjb0pWqQlKgIF6F+jVBmfhYw+i3swizx
AuaGe5SvxdzgFQS4IFOTJzcv2NXCImNJHFKwshROipCSVvvbSlpoVCit/H+xUYT/
UntjL6tX957oD/shGQuaM9xcx3ET9nPa7FXVE724zttCtkMeWc9fKoeIDe62wPQj
Nq0UkoZSRDaRH8S39GIaD6GovwOJeUW75ocNQ3Kxz7a9veN7rvbWkLT5AN52F/aW
CgbURdFY6X1bOlHujI7tzaqwYWWV6u8tJYcoL3e7bqI1d6oziScvMuXTQb6aNlLo
ihBLsAwXVMOsI5BDbBPuiMrzLsTjGFcb4Ch8m4uvQ4/Mwq//0+OJZpcFb+Mdn4Uo
JfuaL946uufPa+sm4ZosTMwuZ66+xau3rjaAjydp3+N4c0a9wl6D7+r/4g6p5lkI
j7+O5eZ5sYIUGl+nBP5izKO1XdidkUfAPhuloEjKql4wdBPzuEZGXTLLTV0AgDNc
FMejHORUUYkwBsQ1z2bIUG9Qfgoo2DKEQq7zPLmPYXYLWAC3UDJzQKJiVAgp0q26
kBAQFKIqFKunBF6f5bfxPo8ZedDG0mNGpirp0JZdY0Lw/BxyzrIBXcpXEpYL0GDQ
6zQPqvkU5jmp+AR9oTXNlCjrVLTisyXCVNs/bmHnz2bXuPZzWGmW6kn0WvKv/rDm
v5QsdlJwn1jqS5rToUV96D1n/i0yTwHmGcFgvZMeEu5f1IHkW1wvhRKzdCG3gIMi
guGQqsRgp632ignb/Na4NHe+jzOzt1M8wJIM5tqv4db+CYZMco8pgKmt1upm6uPn
2ARc0uicGeFKmgCnZaDjY0g+b/187oztaNsJaAde7KcGIvTLS3ByzAZaEECkKMxs
25uQ66M/cAdo/PGrTy0B2/8ZllI6l6Kj+pBJ8kwTERrr0aimjiRWRS7ym/4ZBhwj
Z/gG5WrW1fZXY7hAMyGx4dzM8UOTh5PLN4bTB2W+Ih1Ld6j5ueRFPOasgDvPoVW2
aeHdNdAv8TOHSwyRCyNHQzJL7mHY7QP9cQMbxevFyki7+3L5TjehKq5zC/uQtJnd
TKqYvgnztrluKccJoIBrHNWtbuA74p0VOi5TNKThEkqTcSpy3/jyO33ob5VN3aSA
jrflx7+bQSHPEwi8M0/Bgd4sdeFl6lHKjNMDL5RZtowTJJQBtYEE9ENCnSlqhkmd
Qe9IaFf5mLeExuCONHF+SsCJYs03dnYYXCFXTJpCyODPZzQJHJIHjHa1cx11ZZor
ihopeOSXNuj1b6SR3MuJXnYQV1r4Gal6U32+aPIxBH7TFYVvFYCvMO9227Zvgt5Q
2+upr22VZrZaaFwvhvbemrALdwUYNSOXI4k1MSWIzWUnJGB+zc8cDlq6UOCK2f2G
esRliZucA7UulpcGRIS76BboXSE00qkE9cWKUy5wA1Y0u125J0zvjzT009Fp89iV
hPjBwLZ0cB8CefGDBxzVxEc5+z/mSzr3hS4FVLXzuza/MHdyK9Cx2O58tCwNlpod
WrTjYzm2f9ne5H1h+5kesi79FL5o+SkSEq7irKRPqk5VWHW4fSAeK8zzh8QKOcfO
yvlf0H7kE1TReQuj4eRFGf0H2yNx7hXE+r/D5Pz3z+M+3m6tSDfz+81LSkd8tBfW
GiXYF98cexXBjV6TfbfWh9g3RY+UIgDbWc7hU7JwgzPntlWd2my2InfLNOka98CK
SSbJZV2xpJ9fSg6Z3dzSOQtMM3jrb3+LMHiHAIMNuDoh4lEoEg1FDvNf0CTIKnVj
QOhLylHGDh3B9qHoR7EUUGKQkZbkIwvTy0VQiW6omMueT3oHz8s3xzv4P4T9GTb0
bzsEFVcR3yuUws/MnA56PXWx99RoR3Az/9YENwf/7fHK23LpJ/VDhwN+T2RYzPMq
mB8iO3kPxIEpvgtg61G7DSEFnDfQcgcpyxOq7fhoAd8O6rQukB3wVygMTq+W5Bea
F8+kL+Ge+b8ZRjx5mN6ea45H4pfO3k/vPbpRtUhhx+Hbx9HSr+67DCmUGnBEtzI8
e1ETVBF+vfAvucunElA3HRpcs0CdaFUWWUAqTyp33RMfnBi5kmAVjje6qeXyaG9p
IMjTuY8GNwBOZ+y8NT/sWBriAPOnTzvZw1+mQ1qRDyinxfvuFM411oxe4Oy9p0p3
YBvUeZztq36gSH6xrMoAG7NtD/jcwq2KMimRMJPl1ubpiwnDJurq3i2kyLqCwTFi
R7Jx+JBV04IyzXmzO5PhBLXoKz5vWI4OSsen+wiooLDVeEkynSJaawMgwu0D0u+w
lsQGNPmcT2QfMoYlldESoa/LisNfJTVj4zwR5mpW0b3BVXHyq9GeOaO2BH0ArJzK
uwO03dr2Kaittx4WM2dqqn0knmmulzSXmX/0t9lXAdJg6FyfFiun6LvhmkVbPMZy
la/3006EG9if2yygIf78ePKI92+HtpvXWHIiVmRjIrcN9ruEdZrstz/b8d4VfnKg
+A1lwSQkbVk9vJASiGUshtsh6XpWV6skVJW9F368NVUH179wXgck3tFcYQROJou+
/puAlHFHb5hl2hafnam4CGkUQlsedTT9IHDQuQ6KCI4WwqHhzswhx6j9nB0Kyszp
4hXZEhPsD8Vb0bHtFHw9Bp/KEaY1WSqKTH2bzynKVz4rHVsVatfleHdl5akyKm0H
9YMPcPQ7/FPAsu0LzAGxLKLU6AyLwQq2yFMnrFPD8cPT982VOX7IKA/yNQDqOo2h
XEMgWyG5DVq43dW5tV+1Slzz9TqeL9OgHTOVy2P6aPrZaOs2GIsHFUQugwrOfWp5
C32quZEvC8ICkV4jbnpcf5kxgg2UNQUV1MArsjhUWTzeG++s45X/+3X9efzyW88I
II50Pk43lCH8EpH+XZt/pYXergpkI7hE9DXhwhxH23aPirvOj97n4vDb8WSYWYc7
uRoZkQnY4uSIOLj6K5AFIja3/BPTAkloCD+TVaydwlNcoHLP4VbCimTHAaTMq6Ov
ArfMshMfI//vw72jhwSfHi3KkEaUbVX3YD4jr+/pGFdff+yYTWINLKgRPBGowk3a
nmiyK03y6QBMMBePUhpqHcIcUb9Qztet0SYjmbKFrRURldAdjffRtN00fJnUDENa
Mae5I7zw6Y5WJqAYAKOY62os6Tjh2WFI4rPkG/TUY6JSFRW76aXHGhLNHX8mD3sW
aJ5zh+r/9hslKPgb8dY7L7ttc4DmbHFL8adcNLcaGNb8PhSEjLdjLVfHxtnnJjD+
tdN9N6v6zqnZcqweiTh2LVFOnX95eoEUIm2z8nWWh1f5ftdBKuNMn1vLrkeNX0pd
4IBoeB35M3EnqpV+J/4DxngpI1g0gzvWAf+ffD4vR1U8WpUTA5WZrX3dOqgVH20R
HY9LCU5I0UaA2b49Zfl6vlpJKFXgObg/tHNqPOGf4OpT4m9A+2WnXQ0cY3PG7jwD
0DOslpTK8uCVu6O7KoEFCPAJyjkE5004pvHV1GNnoeGsmDHCH1UmwhSaowFk1/04
nR/fJpFnkR/guVgaKhld6hYgAC1l9icr/Cb9rbWs8o/NS+3bjxsIqJu3ijTxpfqp
+lRwsp6UnJ83Rim46DM7yVvIs3sRPqjM3AXYU/j4fCDMSePC0QSHlj035B006GhZ
fgkHNxcjOHgwWcmUuqtZEvuvpmuKieqW+faQ+DdZP5e+no5xP2ct84MK7fo2B47B
idS+rscQ46pBwDWpNP4VUvpA4iknhL4fXCfiDQPgfHTcfJuCSfoT8235KW2QDBzM
hL+Xl0i2aRZXeOuZDn6h2juRvuI3AmIZlDBuG4pWKB8JLIgz2ZDQa+cmSla51LpH
ccWk3XJki3k5gZ+t4epUiT4vaWNNgA5R1H1bxL9OZoFGkacQrWoO6XhnbP6sGMrp
7fFGx3nROTV3wL/N0vaimJEUCXUaD+MiXr1LLJP+T8G1qJi5Q/hm1Sfwg2D6YmAU
Xy+aTZMqaMTKHYxctuMKJCpUASXawK6caGhZwr5uGY5TOYS2KJhJAf9W5A+XfF+v
HVLLx9GzocxHw21vheDUGyXwfq3USFlCKz6RI3jTRb8HerN3iBjOQtLc/XUom2q+
+a9XL1DU/1S8qUBwXYvuf49zaty3pzY27JLkB+QHlJgvsA21JwIrEdzolNy8+ysW
jsPQysyXZnhQzSm+8q62ycDwCOi9VuClFdEz9NIBMlD7dvPAwTjzDKimZ04iC15A
JqOwAVnnrGz24OVPQbBIzH+cC84bVXJdmksZz6IX6OI1QUm2wvuroD8Hm7psYAmx
QwJ4kHrQpwVDutPgEWoKxQvXOJ2/kpyQMq4iRTrseBqLE1vvFlCeOFy0hCB2zWDA
P0MBfSmE0Hok6m12eVohSfzFUSWR/8XWkTp7/RmQ8+Ocoz3tx1VTZ26oPSOYKEAq
pty1FenPrYrJTLjigA0FlfDrivyiWKBu4RnqC7jG5XQKp0ctdPTMLj9EckbkxgHw
DjzppakBY44xiJ3VZrfR0csYXItd++uBA0cbXFAvdwZmJ8qTX3HOJ9s2YWcM3rxt
z9mssivNc+izmgTVY+OuX0U5VFuqyMwfzAx6VjQwZwSSvurmKBFpjVj2ZvzGJwRv
rvSjttB0K3jcaVRpAUezq6MuBVFNbCJ+5rdcZj/r3MTzWJpQcgcVO+8R+vUaBLHI
ha05SSkaACPjgQ2JcjxIuVjsdVek8szUN2RDhEpq7/hi0WUT7Zo/NMaq0I1qhVZs
G3SHxYRS2Mw6HgqXK2wERJeBLp1KG6UDWBFh5PLWBMkrgRu/sXd3dP8EX41HHwzR
pI0aNgFU0i6QD4WtwQbF+WRn5hsy4577crBNeU9rU/FXEjKrTfsESOjeYFlOm06x
TPVWrPgoWrrvkKFnwc6JBMl3KnftTPwAetqTC19MSB3uBFI6Z7OC5xBlS9w+inHU
fYfEZ9X4Gj1OwHJMQI+QJf/L4pjScQrXhzt33aC1a/6G1VaUTB3U2M4m/JBzcaJi
RLsUkiO9+8e0P+7g1tyIANZ+O91GLMOMwJ+3D7DeUXI/JCKkx9Y++YMkamDWYpxb
8q0vrAeJJqF0abX2sKkCwqHBeFfEJ6M+7V1YU896RWSFxSwR8M6KeSFJF/oMPUaJ
ijB1b4AjehJ6wv8ZGGhtnq07oxEJ5VD5dFbbu988VY4tRHsnpN3PjCbiGBcTh8+j
SkORewSp1gA4Ld9/QSh7QTJyhfiGIWJrSlaZNvT5HPCpaP6kL8gRIPFh9t4lMTiS
nkJM+82bpUhDMDXx5lf6PE1QBTAJYD5p3azYdgmQ96ADwPlkvjXy9jd8MK4/M8K2
SbQ8CxX8KnWoNt4/uewX/5yZEt5Etolu/fcFpQ55sasFM7r1Br3eW7Gv6HWHIuFA
5COo7VAGNluvil3IUa2C0dS/PPQe/AUDapTu/2hcDFODDr75M3zR4Y4wR5J8SyzN
Ofn2SLfZ2p6eIA4qDWevd36dsO9pu3evA1BqsBpq/MmanXKvWQ9FSWwHUGdjvVEW
DvXeDyshAds0AbOQ0U7twH6rqDeSsLX6pY5pffSrWPwiIua62D8A2RB1xI47yeKE
HUqBF1agJdGoch18Q/8AVCPupr4G8wQt0hJGa5uC6+xg5MiDgDuJZUY1gqJV7v/g
juUfdblVKthPLLmjOPORnsCJ5nO83TJw495/TDHq2MVSg3O6EAhF9fxe3EuIWyAP
llh7L0XfJpLqrzgroLKnDr7NBpUF7eJComJRQo/oSMlkINbpxNqSGGgxbFiNk1eP
j6pcfjUTejmKPY2QA5Y8QGCFAHk2SPL0kKDY37aQM6GEAE9yBIHDKuSuwlZBZwMj
r+PoIdCm2QaDYWGSTlMJkkYYQXrHSbb0JEqto4LQQF+EaqK+iY7+1tV0OIRuO9Cv
r9V+zRQlABrCwo4/tLrcMyjNR8e7nz53E0F301xaPzpGbmi3MaGzvdiZGNOQIEea
9XYxBzUN6duV8kHqIlNtl8Dm2tmfliu2kjncr4wT3lyZIOc9Tx9SEQP5EiApFnUH
h3ZGiOAZNahSEiMJ4xU2mH+Ruiy46JeMTKmc1iXserezkHx29+eHwlqC1HKAtoeY
WWGevLozkVLL3mTTj4dmAafD7JAq7Xfd6hfj5xTH8NQ8xZkS/ckAzHFW1M7czspa
6raQslpULAsLMwMaIGYrEcbwCF9Z/tIgsEYqfEUrS1CWF+dewNw6qQtNcPbxyz+h
ZRP1pqzFOg08l7QSumXsTzCBJSLluDO9eF5cUarrj1rqC2kSRg59X+D5rIz7ozm+
tQ5SKxRH+dneMr6X/1y8kQi5kE+7dL7S1VpLHWcOr18FKf6xWomdR7iBnYICFMG0
jzyqpqhmbkBx1X9Sl+U4KERzstq9ACgMaebxo/KODVpD6ZUYq5HrkpbluFRV0UFS
XbKUUfUHHQiL0qpxlont6+3kvWZ9DS24u0j2TUr94qmyfzsfmmOIEFLHdecu5n5+
kXXNMp+eyof5U4mFCNkZ0/h77U4sgCAUkCvrA0p5uxzyuJm4iamV/n7Psee+OgXn
MpXsaGoSNTaTm42Vne6lNT/fFPm4nDnE2sk0lLhvyS/QS9xjWJEuzV2skbsEZtB6
b9P0bxJtNu5ut1uafUkwhjRfYQuR/IEIznaOMorXLlZeXh5zmhX4Q+Q/GHUfy6Wx
9nHlnDwi4xUClw+bplTs/PdyxJUA2WTpi3ptXf3bKiBW4K6bJ2NKEAvoeuf7nVLh
OVO4NsgZnjjllAiAdEfD76R+dMO7kiOXMUyXGigozNGMic3xBCCMSMGz23lYlJ44
jaoCQu6x5t0c6+EkQgWhaBE7LgT8KWTmDnEqaofnh8wdSUspYaDZjWq0E/fFiqVc
jLPB729vQlmQcG+WeQSfFYl6XJXKlwpBMrU4RdI/jteu98eDITOn9XZ/Wbxc/Pvr
SDUEzPi63j+xwkcB8JWMH70jhm8ccK6/dayjGRlHOtyKpkz6yxUrfRl1Eu2ttaOJ
qS17gCCuD7Deb8ElG4MdZ3bnDrpWrqsEt0nGzt6+LL0yDr4svRyikA8Btus0YWDz
9Xtd/iB/pVsZHSH2N5QgK8s7+Jos4O8KWIhH824hpSZvUyIgYxAifN0zrmP9xchZ
HKXUsZSY/GSbAYtA4inJQ4YqmMv+zk1dPbd+19gW4CwqXOO3Mqi3p6gSWOdjDct5
4fJI+m1e5wpwM6MJsYe9PzENniQ+/g+NSCJmf6/ImsZbxuw8ZJBQPRneRrQ4Fyuf
xGMSft+OBTWPCI/3vYi/TOZ4uqqXKkg3yTn7ZQiLyhBl7G2vlTNR0X7WZMCFQQ3W
T7+uW45bmr2WfbCUBPDMEHaM682oQFgkVlw/gJOW82MMtbYT7a44GKmazALl3Jtr
MTek5hisamcVufpNO4UzxpGLJtovI16V5yFtSuJRCOE6hAusktX0Z+UU0ELGYFXB
6RnfBtXQy3Ch5hNC37T9uKx61jfSHottHhZE7X4ttuP9pi4TuigjIbYwbkYMcHD8
phuDD44sTL07IWyNSgauWa+w/IaWOSWLJfKuSYTYx+uMHSijF2BCpInh3KbX1tsW
v1jjevHuIv4mwLPztafOnkF8/HuqF5v9b9++sJm2PiPOF9iOWwvMa3VZT/537RR3
MSK8AQ63RMy8F2riN8cCIQqzp9QtFQogTbkUhmH6UPyhqNmNCmvpjcDwRZQw/wka
jCpNxcranLCnjVwY9HVrAeDsY5TfmuFnfbbuOSoxTe+/GAwjCiEChofkmM3PXZ7C
9YV+5cy6+OWmYokDVMOYea/R3KNPsXCWXtUzHfGyxZdfiFMUrpxSpnhJUKAS6yu4
dxw1mOc5a5chlGzY04EVzvFFWE7vKCucx5qPO1HTy9q8Lp5JpBIhSTex+SQ3fe9a
zseOzxZFxtfSRWAR1RfIeDek0ucJm4wTSP6IySLRzqz/VQPzgufG0SxXPZAxVZ2p
hJHzfwMyc/n/BcLxifqfsmoZCxMCl1ninfJ0tzRIAo0+LUkLXefNNGHUdnDKfwZm
cLQJP/PMn6XJde5zT0yZOp0KpK6zZp9C89YCpXGw0pDt1r67GElRGa82wRweCKO8
hOkn7lkrBoldttTG6JEfVpVk0HqSuYtj9xIr3qgjCrdKUaF+cXVO4TyvKxg2sZrM
L8tnys3/tTcjPg3CiIQZ2QzhCE29Fvg6PL1MQZ9aQtIuILRtreAvmxu3EmWKCJOu
J0Bi0CL2XGPycVrIPjk5sEmitYOrafgbHyO9po7bG0CpJ4KV39KP2HjhRGnIl+Gc
Y15xrjkdjedA7Md2iJ+Qwa5W/iq/KDRM/aNmmECELV3RNcr7wMoeu4V5gW82a3j+
umA/AdnnSHHIEoFmbKzI01N9ePPBwgTe4yv+9usNxk7PGZMg6puR/bAYWZhSXLr1
rEcslWYhaLLoDOHuZUqgYM8Kmysokw+PlBbxIlUQ5061dmAfwvKBLPNzgCXF2BHy
8tRAp45ItR2s2fr2J+ZuxGkwzWAxs5AjlfPxY1uwSvNvFSquu8nXajfyKW1pkmB+
XAGQ6d8qaQaVmafFe8q8Qa47v9PMwU9XomMV+eZp9WHpi6/ahRWvXz8IsHaKP755
Twj/DCRKZ/Yd7C/1p99te9zVUlhDCzgJEB1Nq+58j8JK6lKn5/ODj7V8OopJS25J
qPuuiu5H++6lKkxrCb6QLN0UjLpa92SB6wdxQkVHYuzUy30IdGQYfbQOktJjs6go
QtzVfTLOjg4VDtn1Xlj0SCpqgtaAMlrY+TmS3QNG6/vzBRqRKenf07AthCF6k/OV
gGyrruKiTgTG4XKZ+LhrFJu39q/L2rcXmCoLXzBzmSOzgvvXedwAxbuQipnn7nJQ
6j2LmC1IJupcKHnteUIr6l+Az1aFqR0D8JtJlfz5I0PoOTsOBt/J5SpENgA8xJrx
6NDy1dSvBgIM0hYr1IU95il2LW8iyoD9MN6zs1kVP8tQgmPuuU0Ubkco6L/qXPJY
Qs4YYkdFj9XOUtP+BiRHdpwlkx9O5WLHIoFU+WmybW12a+gVe3KOcT53gts7EpwH
9MybBniS/zXyKyHYvDt5nv3p1DsLcLmMYfz97euI5QrEGywNrp/p0oa0sTJFImyx
FKDHhWjtMT2AoWRaTp8cbTea4C1Y+h2ntVWrpPpv4MmNpHtfAPkejwCPXwgNV9MH
x1yrV7nraHOlOfADu9XJSB+AU475fi0H7uBbTzpC9m9bsrJDFyBayvBE/DYWedxr
IaFKHkdnAFeHI3Y4wmNFep5mlrs62El+sZolOWkGw9nNkEZ5H459pU7DMGgIiC2G
jbdqMmH6QsG4UPMXwqmLwZDm5CBKYhN/smOo76TGhKgiCufuSZmXJLjZrvXy6RDS
T3YESPI/QLcJWEvUsDO3KiHblji+1H/dZIesIi1pzrgqwjbtO4YngtqMz1B6Za0S
3vvBS3ZrOuCg8gZKHhQ0fPRlfXFOERAN06pKMYj/Fg6xLvwXQ/k2CGC1wycXwEG4
L4B9mw5d+lTrkThJ20mVZhZM+VdnzV3gzsd5YvZotu4nh/HsuVqbSh2MbtGaCPJt
FLr1QiD9lQJ/vig3UA8wRBdaSp61R5lTDSbKOaL5EwtwCWRoqmkQIQKbtMxrlHSz
8sXVYq3lKAPpdq9dyaPIVGeqdI2YnNEFMk/aeJPQrbAfzdL/EwY1p5/WNE+5+Tj1
N/9gGEg6Pmb3xg8v9dSA5cWF/2q/tcS8I4agIrDIu9f+cpSk7r0TaBUdvoag14Vn
BSuO+g1DRc1rQxsmKez78zEnzzrt0l4CBZOF8fqUbIlSdLObvU2fPMz6TXZZoTNj
1/vcKk3VeJcTAla9z+FFFFhZFxoSVNbHqzXn3YEHa1CcwtL3InmzUGxrbgkd5O66
NQ82Luv3jmmIrwW7zmK6DlG3nLqtIS9salPpIrN0g/9RtdgDQVvixaOGGkXYdNWR
TpTFJfcCt4eQ2jZ7ckIupFAcRIgWeRcFpD5yVSgknfOVtuADqYSXFCJcSltY/QgX
ehTau/BQoVbW3xiDxJaYkQ81qY6/nC6NWL0NqbgZJr/O1cflWlcIk4vyYO8rVXAN
mzbvbZsju2XaFNopXXwVvgLliXJO22t5moiXuoVkW8NO5t34ZSFNZm/uQF+hBbB9
t/76/gLw4UzKPb53Bagfynxe6VD4+dpahiybP2mCEkCLPRGIJttIfNMdwhB4hk4v
NhKgotJhJaxYszEmej+jsiq1v5UBqzQvLyQkyOkJ+NYcAWy5R7kMs9kJ6AotMI/L
JDBdXEgNCUqS4I43ng6PCkzukG8aPKSa7V8IOOQxzbdJzns1SfbeH5zi3bhng/cV
2DbnLkUCQTuFBH5xvKQF/rx9S3+ACRse2fPLN6i0NB1l/pBAEIvxAlw4g8p/ttdy
0jJq1v1m6bQtrZrY40prIUOI1PFIDvTeDcd8pb4Y20zwRV263F9di7+5Ep52S7qm
fqrmaGWy2+fFV52sFe5Y7yr0O9vjBMs3FMsQQdGPsTyt87+933Nkma4ag6XqxYKh
49ZcStmhtM5T4Rvgtcan837vTZPuJjDYklIaFvzTsKD4ut6fQov34EBY5DfpBto4
Mp8lg7bGR5SlxmpgLcmxkfaZDzlhLS15iZEKeRxEwH2O7Mzhb6IgLF5OZLJDxuBT
mpwm8WUgWXWdzblav2uL/ij8esNUkr6JyGoL8FsOHT5hXESJDYHMfIoKCqMRYpzq
I9IZRZ/bm2mzCNN6iDIDDFM628jbAn35BGo6nzSM8kAeoidtk9UySJ1FoXBfbrM/
oh99ZgOduSfa9OvFMW8IZOrfRvfJLn0iAlyTAuz6JTBnfLxoyDhYCV9tVRF6WfwE
joIK6NkmvSewQzpEusRhPbPXQxZARt45Dcw8fMdaBwutMBjwzXm7F4l3d97n+ErB
jZ4jlD3lkaQUFe8KLHjfU/I/OjNJNqUfDru5U1Qqko559t8fg6ozh6hRhM78MXIi
DA9KJ9QqPCo2VZ3KE5tcgm4d+PlzxoDsqf54MxbjQ4/IQDqZQ87QOZLRfXKEH6Kp
kXs5YETqsqYnn5fqVnJHHHymHtN2RHkL7Eu42FnWTJmsVaFHz4i9gqroFCSsZkZG
Iz7QqzUpScZPrHt3twyPxVRs+ynU6ADjfpA0Nj12j10YqfKoSsv+wM7FCUuUn0GI
YAf1quJVqfMDFsLm22Dfpuw2+4YdgXlEsgBgK6vk86KpqtVixwZ4wawDYVsX7qnC
2IA7ueKTkw/JK/FWgbjWxMM7/zgg7dMQdNvJlwmvEeTzuVN5jkbRVqjMpmEg4jLF
Iz1liunvXscXICxBrFYyXebFkoZmsLRg4StCMUqXgskRgROlxwNYqzPr4Ls42SKX
LmgvhR+28WGN7oYCzTuppwcvHsK9kSPou25ISxMlo9wOiHXQ105Ejx8OZ6h8KSTW
UFCZA52ulZRTusFUU32D9ReC5zviYN9+ZLPEM2Gzd/0tIxf9zZo7V1MSjP8j6OW9
PxAXOpHTqaPlbDE/R8hEM3i5hvgXj0PTj78pDj38AqLjdFUgfkgRMTQyqK1Zs2Ah
EoGpADyrSJdI9CSEcWg14J0AR8/jpVyh4StiMa507SHJy4UrJC1m7CXHrlNHu4mV
YygeFa6ZtoYQT66VGrSPPtHF0me1ilAVLP+Vitf5R4UQO5CZmgV/DoYCZlJJKuTu
CO/d/9p9lP5VgUo+8e9Fbu2jAjHu+uOGseTQWublB4UNY/1cVTNsaiYPp1PuJHR5
+h7eVCPufa0CSTE6oKwn6L9uEpyae7wY2jTV4BkrwGdomaNYwqorJK/Uuo+VOdun
rXp45UWiSHsf1G3Rwd5+CbC0nYgucsC1Tl8+Ev8u0PwG2uLAS2x/yIURrxZf3+DL
VWwAFoG1El40JylONFduPvfdOImK/fi8GyXb4AZwbDZJY556D8a0LOoJdVgVbSOH
rTJGKxOZdt3shwI89XxakkA7nGQe8nIPIdau8gocj3+vkBKrdyJoM2aMmQJjfEJs
yFEbeBFgstWD26wp1AYwWOtGNN6p0c7FWd3rJ/K8hgIAc5Kw92rt5VQUcYR7h+/U
6dgnUrvFDDdML302Pk7JwMPDw3G3sgDtNhk2DK2mCMm7BtudRbSBXA5rvkmuTkB1
lzX5C0ixzRY1g0isiYCyXf0bVTN/RD5eepQvcqt3dA+j+N8GU85eKHsYlhbzYU4T
D/4OG0NWo905WyFsiSTzknxl2IaIl8n1BYppRl9R/jIPeRCsVnx61ZHK+CmnmB/C
78GaabYFc9o7PnaI0nCbTZvIrNykheV2e5kiTAR1Hw+OmD0OYydVNTfcsQBeJ9Ge
FLpLGbGl6gCzNBdO2pKroLPKcCOlOQZxXTckAhlODgNLs/Oc96RArVEPBvIcpGS+
pGqqUoDqZMaoflUnyIn9QEIMMF0jG2I4Ep0PsmQyCzmtkIJTvIUdq3Gv+PnOLHor
p/2x1yy9Ae6enjfSY9crQZPOLhPQ4YglLzvp5InjJ6ObJJHl512mnA4NveA3+e7w
QxbsNCAy9r7RDNEwEiRUFr+PcISlXebIZ4d5J6A5jmK/1WkDjI1ydztjDmDRboVQ
yTLwbm2e3JnRk+TXotPyU7hKfxafgureB/qDUT8E/vfzsO9ZAchGEc92MRrBT2K8
UB0xbog/r9cNJKbE8VpnM/o18sE8y/hqCkpOlagC0BReQD9ZCArgJ5EpDak0t5Jv
hoUqh3LIyXwn/AE3GsmDbECY8MhOjKqaXCbUS74Sh7ZQEyQKgGq3tBTcfyz38VOa
5OZHfuFSDrndlDQUSpCc50/Eppy77zWcYZ/6ZZ1XphfoCZF2iLnLjmaAvkuYfs1m
B3LZl3j0lLK/PeiTJzYYOpb+k0XpFKFqzy0iJZbM3WSHO7cb5PgfAO7dRb1x7FCe
rFQlDbzqKaEjPAbVzGf7nNggK7YOxCP3Qx/+I0zPUY5H2pOjlcFNuNWT5clykSkS
fL5SPK0b1E8xGqlEg7JnVOpMZKs+rvabHid6Ci+AnrUBzl5CjxucxsNOxRsPuxPw
jUfWJJzv7984Xdtmmq436siAB2c0sm8wVvGqFheOLH0ueMgcJpGCot8VkqFXn5+m
7UGQ0Ztbs46EjTjM3xLnkWt92d38NcYxfRbDhZ6wrz5d7GoR98QgUx8yUl9esl7M
wYHoEA+iHMZloZ/CgNmLEcm0V1wtEQ0Jplh2TUH7DFES/kCV+t4LF0IC8omrxTA0
6l29v5VV6vfYwZxRcaBnh9118F3qFEsjz4162MtP+l+3tJ0ENOsvmOdYba/N0EMX
3eUUeMJ4fe7VkT3/Opl7T0685qQd4sL1N7jHYD91UDkrBqf/3GOzYIQg5Elv6E2i
Xr3MB4tvSmgtmiLozGcsp2H61MNjIKR2ZpWxJlREwBNe8P93c/Lr8XKVsou2X+9z
WHj/wGyqB4/aoatKVs7YdeYw++Ct2qdCI3hMEIMFj2NAexKK16z9W1e6f+GskpEx
9MQQ8Wzd3G5XFEmdGtej9m8SdCKq40N/jL/NzFi4F9DkOM6mRF6mKcw9y97inU1a
gJxuIe/6u72VkB96AmhFWmkKAdOeO8NGAI0B2ZvC1GiaNW1avEluOKvqdtKFQBtb
PR9MN+bqknJI3OgzkmUtkrgsSF9RgXOPf67GCVvrQSRYd0sL+3WDB8FztNkm3CVd
M1GpAIQkNf/6gXB64TuV4rM8VlSvXmMbTuV1oYkJyz5JqGxkZW6zJ8asmlzIQx3S
Ijo4FXs+W+xZ9WR+9iR/F5/o07UqBVh6HHT1a956ZTMEuWoz0UeBYrnFaA185UF7
Z/lidzKuiY6OJigznOx5JxHfqykUaLRG7eg5AQr5og31h/ivKjz7L8xYYMw/q+pf
Fierx5yrj7R40FEZYQndsn56dL8luWZGFIUJLUfzha8yFr0qmp+tSK1tIMVbEk1A
e3mTZFFngceBaXxpCCGaQqWXvp6FNxhGVZ58RhWVPiowssLbMKuCWGWL7xwwRv1n
fG+rzAycJPx15OF7n/pjdn97wgmmlV8mVazH6DpVAXpnwYNIg3JlbFzQoKSt10iU
P7oslTQpWDK6r2y0D8iCKOC74Zmefr8chHDX6l9gUc2BRsDmZ+wnlbUXdqenaPwA
k746uvj3E0TKBGWNwF006ZxOaVpFKrVCviTi9G5mgvmRDZeIIrlFc1kNFqGyOvdD
nJa27iaSFotZahMKngT80gVbfoy8k59VkbcrM8R/VqyXSXS7IN7Yc2Bv20092s4Y
psZ2SBTo69KaZPfvvN67DLXplI+khRVCec4vcHlk3vfWM/npE5twmkpJOPfK4kG3
6MhypTj6OCS6Ya3ILWV+XFOtJhW4gcck+fW65coNzJCJKC7Pes7aWW1i1K4gyYop
XedyAia3LBH5WeG+ryns7kyzfLk3QD0mqS4M7jcLW++jA5l82QeGRgfweBZGpj6P
cTm+/Ff2C5vB5dHbafOVCoOgYrtSFrVNphmoYtGSrsXRTSdm7bwBtxtYWjN+pCHY
x7xoJQja9tyw23RCysJOzDAiSku7jbkVXBPKRPJt6BcwduCpjUyi3oNQj7t4HS77
xM/2dXBemAsbOHyXW2GZD67TFKve3Cg8wrlviAJ6THGD2Ip4YZuiBQCXwwzf9Vii
nYteyIz5lIXnGW57uhUaa5DMcchHH9unDYhP0zvDRjiQ2NapxGfQlAE5z3mB1ZNj
NPVRSVHkS+HV2GRAQWkL3DI9FRCbkhEtXeWGzv4MLrL8uQzspGBq5ggSngoAbwGK
1maT18M/e0w9lnCx63doJhD2V5FF19uxDQJvDEAj+TPXXOzSw8Iye+GWOQJsvaoY
p5tNPBh9YCaW8jdqPdehO8bmHr+ipeFy+GiAwkLr7dZQwE6PgNIHvm1d7NytPVsl
0C946wqbecCHJyEnCdtnka1WWFikRWqj6JYhGCkYiSnURRETbBJaybasG/2ahoHf
IrT7LY+DgIutxJZwdeOHutSovzR5zmN8Naag/wyjY8lwO7SPJ4oa/lyC7rywzt3X
EpNHMze5TMGRSNgVLTu1lHCV83hPPINLR0h6bQz6r1wM5YjR70gqVD3+cHFM6o2O
E8VxKJZ4IoVjSV/9W6tG55EYPjlifAG1DswOrcVFsZsVoEksraCaxgm8CwmO5rdU
kslCTEwMjv0+w7nd20dTAovJkeKsefQzSFb4YNvVr6XAhTSzL3sdSbgXhvoPvf0W
uBuzaaBRiD5KZY2B7mX/3IHbtr6w55NPFlTBF2z+O/BZrjJmJRRMGORT2Z9q31zZ
XtvuWm3mzCHPFWtL2rDsw9upuAc7Ly58m0tk9e6fHoa9HSS64gqUED6hmf9jEQWf
JvfLdmThoZwDOqu7vAs7vrX3XX0YNc/63jftR9+zg1cJSBNWJBNa2MCoLfwmnBZm
t+/snomUk8Frw5eGvd9A2FNNy5z+DHbOZJAulTw/KMbC8DY0qFddm/luBUycZydV
4aGGr5Kz6p4y2P5fzJflT+0H6ikMUHlVgQkSazdjWxckjnapoSEbpPTUoRBHdoRx
t5xGS2Tr9hxxvusjHOIUtPFKpp563MHNm1pDTU2VHqm+BhheV5cPIlYt3Ka2MrtV
pX8hMkmi46vurMUsX273D8Z2vr7WrMlZej851jhPYkqoa/RDU7HAL3fHpc2+Q1C2
aqKzC90Cq0a0OwOSeY4qHS5HZbdYkVxkksbpwX9XTF6748HtLDnKg1eYUsaAzluX
1X3pHQ76x/Mzbvq5keetWHatGkRvbA/OA1v3WgGylP8PSju8NIv4hOYObA8/QF/0
/5XPaExTtgg63dkHlRZDidzvEQRTYEd7cc142nU+J+m+89rVpcrtkSVUaKWtAl99
HD1touKVeH0z95u98EnbEkodJYP1RqaHZEZ5bMmPzy9xlC/IbsGX4k0rdo+WNV2c
SuCfm57YMjEfiFFmR1VzxaQYZzgDu5qGXXTXQMlh8cSi1Z+NLtXg16gIu+CfA4q5
+ZFyW94ah36UT1fGjGR5R7ArdPBmqkS/TeNgtJgfEsd92jLVQg5vgytDzD5QloWg
+kwhTA4eM9BtHIA9lY9uIMBGPiqkio3/8X1V/o2GObkLL+T8P8fae2Rw8w4s5RfL
PuGLEM2/BMjzL8GcymwOiVpI2yXvwQaAZChQ2jzWAskQ8JfHrrr4xDv72pfJ7YGB
8RFsXIDOQ9TI/cV27U9QOjIy5Yjx3KOLlUpzlpFYQgQp3+D8q6oiRgONEgwRPjV9
C9YPBz4KQop2ehtjgOzgi3995JJ1J0XbWrs4uE4M8pEjHFocf4q6Q7pP607eTzlO
bICaoyQREnGpq5G3nvM3TWFuuyjwQzNIv4wlQHENd6JM88vwNCcRc5VVTCOvw7he
V5RZuZupO6vjoGOiiTKd0+K/irIi4RnD4YTRZTxl023pwhW9Kg2S74eA7rySmOxt
Fb2IP4T4OvK6X3DTOOXQlvV3obFvEUzwDnMBwxFNWjkylNXYSnKJIWMgqjTiyJ8c
5yZ7SCb0Y9S57vzdz7H1GtHszlfJ/r99vL0tzUt52ow5GddwDLW7ruXVLvwBixlN
d2o/YGJ2toNqgBSvLvYvHXTZtKlms88eBLezMfFmbPjSx4E+hxb9lOSCc5jSWw6s
KRsptk04FNK9uy9jAFpNZ+YaWuHbfZfllYg8QJul99HHUxMHvQgR7Kv4StSz09uv
13VDIBIofGr23kMwelSLFIsvMllvI7r2IS+A3ZkUlXX0r0cLDzQXXSx0dn+2t4oM
NLCQZrBPyotcWIxA4a6rvI7pp+xziPPPteYBlOs70yfDLZwrmLrAWbqDOlNI2RhU
jNzZFtRBUcOcjcmVGMwFWDyoYQExQrLc07U36UR8ZfGFFY0wk609M/+UIUSDqIvR
at2zrsYHX2EI2P8taJePxygTOLRCIpkuQOwQR1pDkKqY6KnbIt2SCFssm4A9a/4c
2RxvTyxtU7JnNifNLwSeAgEE1WkQdQkuxFGZFmS7vYVyZkknYrw4jA329HG6Iy9e
qwodK6B5FBW6JkZAEoryaqv0k8QcCUBEQKzZ1MteQJ3DT0r5li0j5GJaVRNPKlau
qtBD1EYm76ojBNEJZt4OYIDxbZcN4oQ/gKi0Bf3IT/7cnC0vZWmuzo4xH3Ydai4u
i/ea30mFQ5Mo0kAgSlWcqhnlgwCajidj2vYEXJBteGQTLZonwlmXZuxBdJQzs3Kj
cJijecQEFhoOpxUKSmwcOlEbXa5u+U0d9vibqaFfSQra8ZybtonqdYqM0/ubsA8T
CulzVIUQBszgU2w1FCRuOfnlc+DLRK4Vq6imCEfWYT7Dozdn+ByxGVmyGlCiJznA
48pDaG2ssYKW5SLhpWvFJ7/prLPAVuJljy60b7JOlKI6W3y9lR4mESpP0wQ1ye6F
DsnCJmZaceMpRCDzwnMkcF9fZs3EPpV+HBhBn49eEJS/tt2oh6TkSBYhdFgEIJQA
kJv3eLHRcA94sHUB+j2Hh+1i4Dv/PBBbAZm+gkGdIckHCTt5995iYju+0NVmarQY
Wa8iJl6tUiSz/C1RBw2GTjn28X/T0RMC/28PUEtesbibj/ZokF3MoeaGmTw0Ec+d
U/8iFpjZ0+mSgyPrYrg2vQ5YL8Gn+y6fF71Bs9iRgcvTb6n4+dBPQBSMhMydPhvK
1Op/DKNKE1v1hZvvdyWnPSFyk608ySN1eStXnz7Z/6FZq9MsdA/Y7VJf2iU3oy3g
hMOyp5Gs6wzDKvshLsW8taFhK6+t7Vr0QTVt3y3lGlTpWqHndsZt3A7H+l4UsmfW
ej2ruObb2rDQScF7dDnn9ZW93B2ivuPtRPQcjuJYOAwDGnxySu8TuqjHLbZ/qaPh
tqGd1fCVDjaIAul6TO3ZrcrXr6IbuoH5ZClevcQLgQ/hVGHtoZ4k+MT2N5rvBqs+
+V5IqMPxPFtGpM235GLgiHrPfyybFpRkOBNqedkrReJRNFATUve0EzKtXBVXzHbZ
8No6L26CjMbglUf3QTkRSQmiMeqNwrIY3wSBh/L2bCFigcoKo5iBS82YAONBWigO
hCLBTAqY5XZc6/O8IDdH9JjrlwezNmg0Sv48V4mRsQEGzjBr1kMsl51/DXNwJ3je
mtiIEc94MYX7C13BD4SBledz6OhzIeqZhvtnN6P3he4OBHEnGAVQh977OIZQ2oXV
JwIPYO1GHgszLPV6kPOpc0rXbeJklUZoYSvd/asCgAiLVbHgD0lVRHW3pxZ4Yyjg
REYi+TBcYhG4YVdBDKMX+O8FWs34mTDPUphmuytU1PzAODZYIle+Vn0OXGYxuReU
0bwPUuihiNr3/TBjj58E08m7AHs2kOKMdSohP7l/99821QN1bteFes/sIsY2F3EP
CFX67Xor3Th08TLYxfOGhhNbc3S95++icn9LJFjIYN6wOfouvEGAZRi+acXTZpFX
fLPxChM9POIYcWg4sy4hc2jnDEH9q7Z87lTOoqN6bVGtPdiwFhhZ3DStKE7qGKPk
SxQdYtJQ/OMock9n6b+sqr4M6DxiXP/OZNLETeVqNd7GcDtFYShcj0blfqCy+d2G
a5Fud4OnWg6VDK19/aOyYhfBKG0y5DDLosq127t2jBGDsmOMfmc1fUCm7SfDIamk
0YXdFVq3Q9h83EZKdr04cah9ciITJZL08Gep4jDTCkFUkzgXU0NaTI6n9CpWZwWy
KFQkGLyd3Otct5zktrDddoMvxB5Y/N6A0jDZqrqNXdLoLwCvjniFDnaS/SBCHJrC
+2flzrFd9XTlzmriMPJOz9Y3TckF1AYNiRbJztgQ92lKJ5xvedN72P99Ieodrrbp
Nql+bcQ8/yRnSfjoNMPxlhaSVJfV69mmT73+OTPrTUGUUv5or5HERoR081e4Bz0+
LCMu7RyGP3kMjPM9XA9IKCr5H6QitTf4VlLjOyvFHxGvANhdrfMgA0kmXLzFTycH
H3jOUSDcBHn1fzYY3SBrnTpVtqXJZrOK8dVcuc4QFnaWLCIpyJrqB3VF8JwxbyGX
PyzwHULhkMYY/xD6+qd77yPP0RzgCF9lSXrSiH3XPDrhsG5qtxnxi60RcSAX0Q92
XbrdsAJwlLJI9q2SFbY8r/wrysZJtQNtbA/TbmJwVIygtjKJK1Kuho7ycnCin9tG
uosOtWrKN9EZ1hWbNrtURY8Y7YEEOXOCiOiYXTAk0RNucm2bboRO5HOzA20y4ME+
XSKUvyPV86+iAP0XNinJ/3zE8N46j5+ZR2NO1qKcfGkP5UMH/oPTBNmkbnxeJON8
H79jr59HTpcqUDfwQxxN4gsGGl3hGuxeCE5zFawZqBRaKjiCbPaKbF8ioH0dx2md
ssBv/VxU4wyCPvn6xF+haZedrqUeZZH1z8IKKXOMBQYNi8mGtb9s3xpNgpKftazB
JjI+qKJwVOtZX0m7FXVnDQEhFwxNtKEBMIKIwZ3hWQ48Xtuiz9ps2YKI04pmWaTb
3Z2kdYwTkRWUnL8MJRuAGe3Q38sNulIh8K1+HjaDHBTxCImfRPhXjyLgt3PQRGwJ
KUAf9RCd4ALQqe0G4uNXzVUct7h/6SgWYMwIF4fCCJ6E6fqbMvR5K0enmUgUFjVe
5koa0O8ApmLACMMN/qkw+QQlxChmA4fRvFZ+b868OrhqhSZB2UshWbg0xANhBZF7
lIIhyRuRaDRtZ0MUHVKJJdIafG8c+7DHQM9w7ma/4cQno5DAnCQXoHcCp9ng52VE
bfSUfVSzqN0JZMo5jVo5toAQuOAcv6LH/dypcbFWAihINQnIosk+5xxAxyAwlBe3
abHrdS0wgoVLTnTtY1MJ8zhN8kqbbxgCJih0CX+JH9M4B3DPk6Kr9QSRaN0UqkdX
/pouw7YrpXWIV2DSaUMVWCcSmoY04P7i7EQE4+pPUfF5ekFrXZjER9GuTOaMXxxr
6KGUOsTqZ9Lrr2CzKAHO1KFik+yBBF9kn/vP7yy0vTsE1TUHclN0vjRrjn+Jmn8N
b9M4kU6jN9UNufNzuxsWC/Bnqh/PtKGwT7ubjhJEx7+0hppq6Aif5gyiLe5OuISe
vSGKgdNRvLsdXZmjqchIgWSGKFQxQ3GIBL0jA3I2M371faH6bwT2/Y1Yrv/cGc0U
tWr5rUyN7wGtekXrGRczRTq6UFCuTJHVN6fJ1sac8DCEWrGN6SrYwlnsRMKLDApu
vq1N2a2fIvaZ5BLII9RAJjJ9NuxyFmL5nW4+pCA32Ct8e3yqMdp8IrB7sQJk7AAk
oA4ugmuyeWArF183880+2HDZ01u/1PsRldPxMX1svu2TiIB9eQM4nIsr/Tqw4Obh
Ke87NmOLNHNUmp44SCYZWYvMF6XimK4wN8wyvx4GUuyHSVLOvx32EkcXUT8dHtM6
fcHwQioWnbDtsFZOdHF0C8dNPb2aLYv/zDB028ieX9yioQ05acalf2uK79tzn+Bn
pjoNA65Xt+3qFrvRfbWwczbIztw9lVc6hChwPDeDizO4eb/q6sUWNK/abv60qecF
RxA669zwz4y7B6GR7B/Kco8M1GaxB9CF8K34APQCWW0uLy04jB1MVwSdkrgqW0TQ
pfsbtFb56+EFpL06WWmeEjOMoietBCjrg+2F4eoj/6fmb5NC9Mac4WqDcA1h1QQt
Z4M8/nODH8669WUuhTt7Wd6hRdQk2yjlJzHKw0VTDVuqJrneEJ69TPPdX6BfETQP
2Pm07Gi5soaCN3+vt1xlIpBmswE/FEkW6AIMMbFcneQ1f+b0cK6U68vgFMoeJ5zq
tyiV6yvwXibHKxPyPbi2Twbp2Uc2CRHXvC/DPHJzNP4Sz0dMqvZACirJQ8Cf+ORh
3y1Ni6gG1uTAzS7y2rHwQMaRNrWdw+ycVViAALnR8gdQ+jlqkcuosMNUnbrAcEFd
IoVhFrzANjNdc6W73hwG/NhAHp6/ZFXoXQPO9faYfKL9LikGwYF65oiHoRe/lnXz
RSbSgDyN4X6dA2K1Ms4UaVhu/Ni62Nzo+SPyRVnVyfwE4zJfeeF636hfS9644YGy
7DNXOl0+VZk2uoGBFewX0xz9POSkbfhJSfQ7zhl8ybBqSzMDuMEmpEl0vze7sES6
/JnrTIAKwWs1JEdfE4LUk5bn7wmO3iqyZjg2PFAzu5vN9Fb41fvWxkA3ssPL0U2B
Tlvx+7VUBJTGYW/4ubOg+Ow+YYQ5OAS7BQw8KEeivrzNDkoJcPLuiVs3fvc3iEX0
mZSeTgYAahyoEBzyvHk5sN0zXr/O+ushseJ6vo5fGfZ/gGx+630L7T4590/m8jAv
iV+BUwPyTXBxNU08K11YHNQ9DUkWR5iyahiYxUk4RHJJFKDLeUzTm+Npxdji4Wg6
y7lxrgSQK+AWDioU2WMJW2B6A/XRroCh3wI66tmzlmlE/7p/B/z0UAtJiSqO76TX
MXas5BtfszoDlpQ2QcStjY1++nAT6E1UVgBp6/XHxJFaZ1vmR7oH2h60vhwC2HBx
CZYE77w8QyUWFHY8H5JVHklEEl9H13OHZ2ji0cKfBRR85cgdcsrPmmbm4xtzuVvC
no8gNwssMBRWy32Vzd6HUuITvja6kedBx+IwPJMO6d4R6NsliE1SifuElkg2fuau
w9tMZO09h8Rbed6B1k28bgvmYUIW8tHI+6VvUQCFw7MxuS+ZTKGziBrXWoLmtwXU
GQeRHOiKGAMxrNk7lgO/W4nw1W5lWh182vfTowiCYM8lS77By5lVn4bVMKgu9yY2
zTsK+x5T39mQ7D58QNa0swjn1G1dkGw1xzZ0na1v2Jieb42cQ8zAaYyOBzymSS5u
4hxPOL1VCL3HIjjgVuURY0nYxtLW9gBYgLgdSftpRy+O9PVG9ZCSUd6VU/iV9N1Y
EhZqs/BTj8Ynl99A3sDZLo/GmsRTvSQGavwx0F6aOIuro7DGbACvg2i1fy0fCQEd
ok0NMuoREYa9qLrEZ+8e4y5ccOlia5VWRIK59uNQ1eVA6N9nGeqjafTYImT7AONh
dv8MOdkKR9rGywkIk8i93ZWD3W7LsYgc0BKRfIksv2xia/Avux+xlMHFcmJphKFO
E3UHlCl2pwCGGX190xCT8sMkamcIQ4Mamt1765xWhIbh4hOh2Ci5GhOb0GUuyLXl
G/of+aeHbYnACfDgsyHi/8AtOjlpMJbQw7wbvStwPWbOjcBHrmpp77CwEjUiPDHk
Mi/GUhIYIQpCF9jrwNo2MRav9ngt/t6fjjSiqgOcfxr3wK8cOGNLFrLJC8c7K4jE
Dz9fRvMRk5uACT4bNM/4vRNryIaAkO+VJRUB8pfmOejviWHgNr8REkfyxJRO8k61
JEq1S2REWP0VmyduV1mjXDujuSkDP4uHEeamWM0yX3tKbNGFEMOdfCdWJ0xaHoMi
FJ909iGXep7oNP20FlJzn5J9+rF18VsZJ4iKz+Vq5/OD5cKq57cA6BzMj+ia2A4P
dfJFuQPuPe3H6OkgHHL5ylsHUo5cB7Pul45kT2qlXgbCCj94EeOLaO13q/QIWTqP
4s/eaStMcbayuk0KEDX5ad90IHLR2wb2KpWL56LQKujGo522/6iwO0MwJVh50nZd
4Di3ulif3mde/4h4OoFPx+MAdF/Runq9VqkqQw8ZL0Bmy5prU8mrm/pVFh68bZkE
ztHYuC5FT9D0WKpR8tWDlMtyaH2upys5t97aTN18qt/yUHQ5QajctKWnrvhYotkd
N+C7OuqyGPOaFFowfGJoh3SUkqmRowwKZHDK4XbQwLGsIat3xHXrx1b9s+73qvV3
hzEEvm1NxvDSBPNYvIkR5wOQJwreCy81lQHAshl8D8h/ctAfT86q7zzy4TZbdLdh
Y6FYt7x/KScO3QIHMkZlPI3f6ZOsRwQJcaLyEZUJJ1lLyYAegwzQlIulIuLXIyue
EQnAl2FGAt0YAbBKznpp8QI9w4Iy3fH8pmrepp0IFnA=
`pragma protect end_protected
