// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
B+ViirE2BqOG8TX/e5dOL3OjRgR8OLkXFjubeS2SNEj8FXKapSZptl3P3upR+vRZ
prI+fqSwD2HhFrE8ePa3y71ezCCj90rXmwblyUkcV6/Pz6oD7gd/l23PlK3wfF79
e+TNbrDicyuoo9HexWu44lN3CgFJaELpklw9+Yn/cBQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10368)
xusf+YgPod5xNkuI9dyq7cKvN9mEHFM8omFU/HHEbzAnUqBDz2z5rNzRjZuTutln
GF9VLHz9kS9gDjIECWxtTkbJklBpOr6lcXcSH8lVUr/WHcKPtYiJsq9hOytOjy+V
ynnGf80l7H92RZ5LaWKA9660w1vBW3NOfiKIPXiXxaqkWj7iTBCS+45TuyNDK7qQ
slQFZ4nb3KmmFhVNgMAiG7VOS6bNz9J4o0x/rRfubdmu4vnVzSNLPU850AVMBa7P
Qo5ZMl9nw4hXOjcAvJj86EKBcgTJEN47NVmZuAZo0RtwyfM4bln5BWMIqwRpku1/
nt98TiSPnhwc7062PbgmSVQXahHUV0WFTd1eNiAwM5KKJcjGZDrf2i6PIhe/q80Q
Rt+wWS+q8cxJzz73GiFJEqXUSuWVs4flRAqqwzdKzkRwAz7szMwrLzU0V19ij+1q
zUnbRmXfLeJSIVUIefzXrW7tV/VRN/pO0Danr77Hp+K1M21jRiSPPbUPXM/A4Rng
mnnJdpCcDmhfV9hCyL8uBrIY9v5HFHdyth3HHgP3ELXcUs4q5FVNdDIwGxQuPpL1
0gvj1iCWttBu2GW/kdJGfhkcTydAXCDcCe8imtIrEcQthSgJZqGoLE7KlJDYj7RK
zpzkJ2BR17fKq/Ih9i1i+pmLKeAoV1pvfkz2rE9EcgfBQu9H3IkLBFksg1MSDo9D
Xbhdud5kV4zlO1zCa26tw3gatQS6esVQxNBwz/oZW+n27/3W5xPpe8IpwHbqSxjA
y8mW5IMpZTqV8XaRRvw5V1CABMa4FCpWLTuxtv4ymgDkhS+Xe2zz5cfLyiAbzfzD
t1r1eMvfIZLLLux8RxBJBFiTklAC3zZ7YknwSzn1BESvZfb6VEShYQreRPKchjmO
hr2Va1722lEen4HBXy0l2hEx4qfH3+7MZo31ncesa7/ENBh9vwu7px0mXAYe+ASI
BXHEJNq8LK9cnGro28Oa2gy87PU6rrNsfndbF3FONWbpmeevtI2HP5x/HR2kLQ8j
knywisQtBAKIv9UxQUJzAlBrbPrF6D4mgdzw3sVnO8zkS4YRSr3nZ4U+IXjrZkB6
dZ7I9VqkOero5RCp3ujuFROXdl1FM7wbUHHUV4xkHK86Y3fzYGEayOuT1HpvKGt5
X/1jUb7x+1M+COUTvxK5Uoa30ZDyuy2iIhlo+WOdEG70vJSJgyDKPzJsvo6q8Aw5
Dm1RVW8NYjdTpK6mIOZQnymeSP1dJzsPp6I2b9KQkHaK6vCz5fRP4kCa3P8RtH61
FjJ2gXegd97i6+9G6mJEXoC5LQS73I5XUEbVgMvrLICLXlU09ul2BbkOAbJXrsvV
w26rxl+O87DBr831f/Sfgr49o28ffuPjnKVmksoVZ68YB8/H6W3cwnYNf5LPWfu4
YjAOMvoQqFSB+qN/2N87XqIBugIzNfu+2DIIVpYB9UZtR+EB4F1fUKrfOiV/5882
l8xnXZOWWv42qA921ZoRHW9FDncczQe4uHcX4MzLGraLukEkEwciXpiH9FW6FmXr
NeJ+Zsucth6NydhIdJzBJSQPHZh86tOgffFUE6O0R6croLQlF9LzqMFR1dRqH3PX
A8dZOAPL1rpME0Rajpw3325jBhMVLrKtjuR/7o+c1YN1mgIaMO9yiqKlQK04z4uB
kovyyIF6tIUVrq5uetCys5T39vbVqWa0+TaDTKI+HayvM0TwSv4RhZxrElCWxkTA
u9M+k3VCPbPGM9mLWNcE8CSOQtFQ4wjF9zfLO3AbkP1df+xRqorWnKYVfVvrpTvh
KtGAqPpf5hXdNooLGk8TemyrruPxkjw3wXNOmoHD0i3hgfSQCvEpKrMYE73kloBX
6JlVAncr8CeJyFevb6C8HzQJHbQLDqh3g4Gxlupez7M3sjKzDbKGWLHmcgSoeIIO
Fd+ARs0TkdGFkdYvIOP+Ml2GJRD+4UcB3YEivg2EZBPYbleGbsw9xGcnz+1BeZvM
IbIuQjrTCkCcqQI9lrDKGg+AFOGCdVOw3EycmA0xwhVwlTofU2+iuPVic+ko8OWh
/RWSk04gUA3HyHwibPey35701Cc7hq/qygFnZlQBpPyCGFGRne2pALellBpWtDDG
QdK0dbhP8SLtCxFNOGbmJQMFr2EuiUikNrZKz1qWwjbfje15hecbfBgXYFmum2Ke
YbMUX3N0fzPwVZZ+vXRukd61UvHsnTTqcy1fDuPdv1zVnbyyiKE2RgAyNB38QnL2
8sOW/pHudlAECPdu9498OgtBF7fCOGjxnxwVTvqRtWK9V92hwUjMYjFDidAJQCXk
J7BrvAbtKkLAD//76AksP34/lOUs8RudTKmvFqb1KTs2qstSROmpgqqc2deAJajj
YPJQl7D1em/uQSwIDi5VuwMPlT8J3svZPfVEiFL1Sf3AaAAfFjiIZA6fICE7HYVH
HW1zaHLAhNjlHdZpHlNccXK7v+vmA2osQVZ5KzN5sNvw5GZgQ0q81Ytw4tDb6b/7
gROYBFI2WZKA/KDXTtnC/GpbexhqMzAEQxapPvrpdd/wYva+U8eJRuOs/A0MyJsA
P06FPAZyPX8xRYDgirkfoNxw6LzgObHEGvlrmusmtuUcerJyyS0L4OxzIdjEMxLK
x4Bz+oPElZX7M770K6TfD6eobPRZAViXdm4tSWgDnU6cEEIGJPoddaVGe4+lM6Kn
oKzVNyWDhoirnAeeHONr2i/Q4Arowz4AcEMuK6301rQt6/Kv5QeGO+8Jl9UuXuwD
ouwEkNGz9O3CCeYilB38uPYlvBZGBaRDScif92tZrs/YlRK8SuyX4kb7nIvPqF8j
iv2WoYaXm0qiO2YprsTacAYwqI5FitVmoLv/ZEhfZ6m7rJEDMdO3fNNzchRobcRA
trxJbPxLAMKYUw0cAEOdnck2JA9SD61FofL2jazwqYMPIR9yyUVI8j9iDykSLGfr
4QJ/UCxLdfebC/w6T2zemsi8xMpGA4JTxsH9kE7nNB5+0gwKO3XFopew5ozQ/maF
uVbhmhLKNY+sWNA2ygLR2WQWzpyEwLn4Pt+FN3kNpLLJYOKDkhQGp+igVyVbPZqe
aNsCYYpACnxcWckXekkcZOPEd2Fk4BsPGy5CXcH16jpchXEp4NGTgFoVz9W/MBER
1Yh6i+QRe2qH/4iPVwaPmRRTbsZoR21ay5n8JoVDbxR1RObGmivRinSuPtet+T+E
JWD/PYR14z7zMaIdEaYXrgjfOXbcpBUfx8DFHCkD0KOAfoaZcNZDLyinh7vEdZh9
bfLLSwOJkWBVUUeUU1mTxFI0OOtu4mpO0n6307IztkAjxbd2JM60afplXlItc6Sd
wxbs+yQMbY5i9Mal3VhDwA1WvOGtGEPAJewbAcdHKaHkTUgJjBbK/4wtLK6L+qbn
CYoFGeNX4HHhxVqiQ0oZwjb6Ds+BaaGxjn+IeW4G7nIRuuR/hNOVCqtE9PJUzHs4
j50R0OFzYiN5p51rL87r9Ji9xTFr7WQUBUrzTFKlLgJbrGyvuTIf9RHSle/uOHtF
KXDrzPHqG+WFYXHNEeHCUUYGHWTvpjyflUSr5UxoS7SIxj7tFriAYKqO+U/DbXqV
U8ClDqo9FLJt/pKCkDmidslvbvOnLLwzJiIJC7tV34UVLtGFgMI9mjI07hi4mDHa
LaYDmeW4XMnKQMabp8l4SOEsz0csSgqv4+vdn8DRuiKaqIfNAWOxRMUBN3nS/vw0
MkVJrqMudkM6zzc8Cr3KyzNWLEPCdPxydBpLGNrhHGKDBjSr+L5BKVZGT6H+Wzeq
PqzCFXNOxYW/qmVTI3VM1gAD3uWGXQoeBqgDqmNou0kRxE0RYj8F95UAKS8TBz1M
aI+ENWxOXsK/UyQrm1oLXdV1MyBC6Fu2w3yxIKHaOFt41lv0EfYBiYABqa8g0cln
xt7u1UsuCMcf+gQ4nh5kkmko9zHBU4D8q3E7Ec301GL3Uw1Hhuxx7P7P2tg0Cjk6
Qifbu/z3ze8t26x38k8y8IOriQjOHZ9xeSRPCYY8vTCiJCewbQwFQrcPw/84ljh9
ZNayser7R4jKfN24yg7PZU4h5ne6DxGlmNB6WEqWEXX3auaGQLo67fz0oq2LDXtG
9AezYI5eF7EZlIfZPvv1+feGhdA0YG/HIAN18htPbPlK3byoxzR3bcYeG5B6ZYkm
FfPwdwXrqsvcGbhl/qPGT74gSGLem+GeeXBPmOy1qTIThH3r45yOcXpSm2NscPnw
JP9XdQ2GaHCSBoMJW1dSlqejZLpoKBiicdogwplX7ebuTYPu+vXYfFkHPqS5l6B+
IhEjN/YYQYRM46u2HZt/Qvgd4tLFm6w4nmeJyCKTQSN+MV7MlEbC7xBjk2FEYl7h
avnMl5/48QUca7oUKqO/wVdrhkf4R1AxwZb3kfT+Z8obso2WK1I8TUKRT7HpD/9Y
eUGdh4UNsU+4LmLfFq37d+k3A1McPNfAhbteUB5JGixJr7rKjI5yHWi1YpoJgUuO
m50Qje7CvALUhlKyYD3SYsw9w/8rw9+ADwrVSLLormv+8bBhdqZ6RAQwtwVNokb/
EeaTI1Kunf+Me0GF7MNfawQlRWz4zQoDuK1c3XZJBxvEJ80ZRTKWF4Y0IWMaReNC
cW4nKazZ95mWoGmXfRB0HCo9Zt+87DUGnk4hoH1LOtWbls7dxO76n1NPkz+R5diJ
wgyMuYRFYb51jAUlAiuZ+3Bmw666bIJ0VDEo2M39odIqoHwPpejLoVnK659MquJz
96cfBQ3H9gP5lSjEr20iw8fkQkjURHVseeiw/8weeWJ8y5C7wojhzjmHzUqCOuYf
xfQUDhvmxkZ5keNqWtK5/ny9j6Pf/e4xpz+gHbzBVt33rpVxoLQ3g1bOYUhAR74O
9mJJrFM+kPAgoaGsbJMjKFb03kb60rTq5vysed2q5qpz4LVh54bIcwwl5YCE0yQr
MkhEEkOmilo/e48bjRp3R0ARgOSYnOV9h2Wr0YkTBCbHOC/LkHxYcGjyl+jrV+IN
KOh3eLokTDyEXXbDT62LjbB0my+SIRfgOUZMPud/cC+w4wCozNVF5nggy/Xx6mss
vQid8jaQaWMKJAiVX9DI9rbI70+hKnG9OHGdEZxFILEqb7oUijqYOWSOaIiMaEYl
sDUD0bR8HQlV4ixKgRnCTSM9XoXzGtT1WT7PBaPZsdMSMBdS9aOjCDKRLcIBWAVU
wLQfljO/0MyfI101MDSz0dhEp1zs0SpeMQ8VweowWvB9vLzJOX2IlOpjf9dplM8X
aTpeDdtnGfsrMOueg8gdxwgwXe/Ifg5Z/Fduqvn6sJB1T0+nlIYTLCxaEl1S4N1f
oOpzHy0ikZrzRob45RvfiMUeDA2nkYu0N+/NQL7jwdnxiZPiu3mCRcWlKhrNxXwz
4Qc8vi0caUrXuOM+8wxWInc/tOpBeUM28yWZe2tE94eVqwSGdhllO1NB74YtH2gt
+hLNnC+ehVnWu/xG7IxEb5hqRcc069mGXCxhW1F+IpZBKedL19lHO6/KTyYS8ad3
XLtgiputz1Ea1nLPkuxMmfZ406VfPztmobRUC6fApp6Mf5CBxb7z9615zBLHntr/
isYcd8dvid2lwsl74UZ0ziRr8OHsiv0ephq7MqxuygE46w+vdefcn1WYWbaP/5LL
yNoHqGX9yvx+iq3rvvXHP9h7ku76Kr+0kGQpieqxImKG7rSOsXM3Bjt7A/zcIK5G
JA0UFOuA9+gcuHFbm47JnVYxf9jKYukqPDgW/LI+knOqv21L4UUTFmQRurx7egqF
SHh7e3kymOGRheWSWLZXmgNRyaHBWx25AYJEnQHxBFuBF5eTVqzBmw1Mt52W7CgH
xCj6hkYpj7b2zhV046fKriGWmMU3Z8qnqEThw8Tdi0+2845vCw2ylbdACXfrQIKV
WLYY1HN9jnkxxRlbhfhV1c6Rq6xpewLKcGwZj7Yzllu7l/BoJF5qtQlMuEZoeoeP
vSHtKPNOdGumjbUKRZIUcZQnAoGBBLfTihal4KZO+ea+MlkegDX9m1Qe0BdzTajc
qEAGpH8OYVk2zIqBjLU+M/epuerBMAgD7sNvckONESx+su1KkLpH7hCTd6nzoaog
Xgku6wdESSrQ8UpUHm2MmjuxbFGxeari5QlEZ0G5bpgHqFSpJbe5Bap2d8bum8gC
E/tuoehEwwBcKL9rBDG4IhzGZXe1afvZAmB+CMkjW220ky36QIcMapFxM5axY6kE
wCyFmkOK7YweHqUZTTzLkSqeOcCo1UEKCFJ3rQeVhJuJw9pbv17weC30GGq2ZsgH
g39btFeYtbrSEyn/945VH6vQS3dzmIuIEZPOzzVSyxqQW/xm+w0ztr9D60yLNOCL
lmTx64Obduyr2bGm+yPpPCk2kmeSKwsStYpmg/mCOYDfzs7IbMRvmygPXcdDXdmx
0UFMloFk+VP3Q9UTIvjGPzm6kOkR0zE4NP6HyoLgkyNcfx7XmHSuaojJM1maHFcf
ir7PLzWD7u/s/ZV4C2eOmWYdqXuGY7MAiBGq48pl2Xuizbl+0oc3J9NF1MTZtLzt
y0Tb39M/nRmay+i6T4evTQF9ffvw2ayQZdZCnH2HnNWij2AwlkH6F6XI5e/9p/ea
NEIOsbmvuVz6V33yPCRdNVHXm7lSDglu5EZJU5NFryfLCCiLiTAsZTZKMvOei0IL
xm+WEaqQXeZ3Si7yCuicV+jfb8jVJp0t6xYjbnasinMKS65vymE6/mbu2ngUHvTU
XM87sjH0ZnS/+5vh8igQcpIZ1a72vccB2QqWInGu3ZPthVE3mxiRXqkn7/BKZnWG
Grb4O7Qpzgv7C2ISNCTXfYo/SG2rqphU2FHI1K105ihBqEDwuvNo4EMOIIBuHUAg
ZrGsAoGYdhK4WXxiexu49niXG2iDGjHFR8spxOhmtA5ZnpyHirBxBJwPTpH7SHeQ
wVOPSAFgkEM6cfG+no7iuZnEM9YQq7XwVAQT9YCCFHkqheynNVicRzQ8uiOTXsH+
qEIt+kX7i5ohLmyuIE14DODjXCrLo2ujNCDuS+X3UTkyPfiwJ6b6T4Fu8g2McIG6
r+ZGgWc0PK3KqZ0VxSxd3gBC84veDmzR96B3LqzQA8zxvefGR7MSFumzreWQbiTq
Sh603iuu4CGJs2EjdrZvuoxvxvv9kLgodgDFUL2LgLNaryO0iHI55YCVvBmr9VIv
a5iCxeydSTO+bgpLghlse/nF/8RlrISiW9vOVuVTE1PijybKHII/NtJ1twlAcVCw
7DdmN0jwWHoRKArWO7azclawkgy2v+EBn+Qvg3k2NJZXA9CTqhXQAwZdfW/2Gs1j
OspCiNNv3tk/QAhkEaiG+F8mzUI1aSMhmB27+UabqbsZIauMwlMBxud4MCUU6NAZ
I40MGHSNs0FZFAn8A8ZFGeBzDi+AGkNRkVa7EixqAEO3YbVz5xWwoKNeGxjd9K1K
iXLgEb682NA3glb6lyXBUhPH3zUQRrsbCNxJP5sgLIIVwGo9jer/EqfJ7eGXIZkc
wOPSjbH+qfs+z5Os0282CLBUAuAGFzZwENVopuoaNV+N35i9ZtmhYHud0TPZpa9u
KOigrqzH1fwa4IjazevZaY8r/eBEAIO4d/GNV2owLEMPe4hSNOvSNBPVGQTqqTy1
QhSnvA/XzglzhZMqgNCN/QyMtyOTdGBgJombwS/6rl203FJPNxD78Q6rr7k9kY6L
5PoKbq9aJPiin9X9AnwK31SwtXGI0QhUMokUBtNbZEBAzzExJujDkUAYOHg2ZAp4
RH3Zw9YSnnc2NRH//ZimjIyqaDMQC5HBLgP5V+CQxWSZ9NPXY8J8mqp2wW/MKDHs
IFRXc1v9+bKLxpoTbFFnuQDXhUavzW+75r7xvisyeoj7n9GaOJDu2kly7xmKSw3Z
qponib8UA1GJQeU2taKxkdEG9+wkvCUOM92i+yfNkj11sLrGMHkslR7ZweioLLQ/
lvstC+b5X223JIJ9KNevMFJco+h1Kol3bIrBDu5WGVOJNxdXst36iccUSbafkWRc
4EOPRQUr6W3U0MHjAN+/cxOJ2eAs3SpPOlH+5FSehRCUeKRBXDB8E8o/XQNTOAdM
NK70/wwgX0oGBsE/GcP5DdpapolczZ7/A+6VjXghy0AdiyIhRBm/+gnFfC5ZHsGN
PlFqpTyBjcMQOsST6MUOLnjS/pVgzemu/LzaAethG/wyYTxMx3/aZnx+askTSQog
zFMaJ1xPolUlZiamVmLd/ZT7WK/9n9ORp9T9iBhjubQpz4113ndAhFtNCbjGBQ1u
zpIpzQAP3G2MISbFvjwLqCtW9to/623N3RVZ1j8M3JC93vSbmggQ6mVjMu5lSvIp
zOsBd7esT69vEZ6XQOlXJV1IBvFYx4WKvPk1eDSyQp2QwSXIGcgY03PVjXa/Q4/x
dMPKKw0ZpgWENgJl7m3vKZwMjFJueZELW+iJW0CR3i6ACIY1NxR7UVHP0C/cn//c
p8ZZq3AiwQhO5sCsGT+DDQLc7F3+NCg9MsbhlFANpvmrd4WhDl7Qc0lgJVydYNuv
DXmo2HkesLzCeGZJP53Rxz27stXrW88GGyn8WQoZTqyMU6S74DFUYGmEzuN07bZY
+NjDAUXDn9dOCpadCmU6SZx4m26lKi5fy4nJ8QAki8PvHyAnZaBiHNgIBVrfY+BL
tT3Cx3FoyoEI1udWSE9OZVYN83Kf3ch+u4C1rTMEVQkpjAEGRteZRR9N/PLSxbSv
RSKpUVSwq7D/H6BiyVYeVioL6Pr4X7lNN+5IXDfML0PxWidllpvsrEtnfVHVultx
POWZmQCbh6/5+mCIdHtFO6vUGZKgbjSVZFWBctIdGCxh5uuj7UOBqm5ki1kjGwNb
+pnZqBwkVg91ZaQQfLragx+e+hKcj3Aq3mQDF3HzEU3MGAs8bWq4dVBV9EiKeTKj
pYrxFtnIi6fpbzGzsRzqYr0z36TGwqkT8PPkzHDKfzm0qtjZRAHMGvNhMYvMrPyM
K0IJ8XyI14axi35VNxH0kuk/XYYKf3uSkcKbIPPMc5InCSbLCDFqDTimYDViy3gp
mGGA/ONYN8fW83jYmGfjccNHGPTmEnXiTM1I7+zTKidU5VkobLCzRnGP6zUBb/lw
hh+F4Q8XQAGcoVRdglJpmMI8tCE7JUAMNr6aZX/IMDlpp8QYhXYwImrK/mh31b55
G2orYZzCx38YAGdU5fFFbLUsxMM6lfhuB4C8O5dfcDLv0FGPaw831559czGPXf+G
HwxYKbJ23VbusMH08YWAZ7S0wsHqQWt4IpRXQhFhwzhiGB2eN9GbU4K8JKjMlQfz
6602a4BSQo3JWJtmlRS33UZ4Rk8GEoaeZ3XOizj2ytsenakfqB2S2vyu29pXjmoo
skXxXqG9gTMyQIOVGoE2lDbBa2XVi3AadwpMAVj5XMZDw4zlQ9zq++oSdDFTYk6w
Idz/SRsQwR2c2srBO/MjOOKFZ43P0dFkPbLZD+x/OazMDsqTVKzYH1Q/wQ1ZWtQw
SMc+OG/OGiGAOfmLiG9DVfjLVIR4pKVnbmqApyVzgEfhqT/MwUFh7+2E9qRcwWEH
nzu/5wYi4fHmrDWHCmcMY4iCFlmVMQEByOMu6rFe5qQF6WI9sZWVOvoORBSV1HPp
zl0AgKGP5msP3NZsY1x5IrCN33Eq5PnGNILY8ZkS6fq1lao7+QCGcLlXsyQbUwoR
TWXj5W43fr84WC4PgAUfcB4m4TL6FTLIEWbaGTUYXkq6AKCJkxBVjmYZFSDTLNR2
22EJ8eZdj/mDjKc9zFUjJ5lXE4emQsnRWWFTi8YB9JOIkpO7cBTW2oEdU5jvU8OU
kmMP2aZQ5spf8P/P+CTY+Er42A2u5N/C0gOu0QmJgsaTekVUX0QETJ5DR6JGnYVH
L68j/m46qo/AQSTDAa7TVwhuN3XPZHAnEP885bNil6nbUEkQ0GLM9X3B8sDaRsRa
VYKc5/S1QyicjboxVwSYa9sDW7rF8JYlBGxoQWPvQRV/aksqDifiV5QLQO0iASUv
GslpaD+K6WzYEZCVm6/b5yNAWeWnzuGJV8hD+cSO1JFxt4daIVoVWXXcZAjV0XKM
QlNzqKausaZMZVr3Uo7KlZMcV6S7Uhs6R+CRADaYIIxKB12NpVWOPqN8VlCzZ1qe
Sx04a8AZW5cFEHQeV1owyHXg2XfZotxfcuwDYA2a6MzCswcJmpdnVdkNVW2Ud6iX
XouOvtrVy/viT3fUccNmY3Bs1KSxRm0WoR0QOFCLhQQK79+KAQMysRI84XMtlErC
oU7D8FKIGKdAfs53/bHC7uFGINcwInSa3oOQt6btzjOxE+WwtOTeAqHSbzrizSgt
0nZ9oLpdvp7QGxgiE3HPvMSFw88N85WJohf5JLL9+nejGwYh6/9ZlXTgV+5z6xC7
92nEKF8pSopAhVEDq/8TizZb+Vq//g3rjLgE4ns10nghLIEqppi7dWb/MfxPd/Zf
SeZaV80TUSRX42k4nRmG+04q1y74Nch57VW2r2uMusu4iv2vJ91EPkrZ2taXD8Gw
IxBCZ/RfDZNqFrkuwOjFSc7o6YdFF6yG/BVoXf0NonmQYKPWttBzFn++UW2mgFtJ
KEZndJxqM6+VU3FO5qdrH/eSt/btCSGKGg2C04y7Vnf6E/UgoilUnBb0j7OI0Jac
qbfkkRAxgg7At/ZDrz9SXik8MgtRKLTfI3g56DbvXCOFBQkMgRi1CSHKwX0qSAD8
67vsn6gp6aotmf2UZq8TBvFSoIsQbEFlYHB09TR/idT7Ei3EB9J7ZB5l6UuPN1yB
BZIt6yT0Log9XYwWll4pD5a0d9zojrS/lOCkxmyaEkUraIqczlQz2HIxKZKatjDs
BAtNvxJL9xYpuYl/CoaauD7BqklMEWCqXU3E2nJ49CQKApbYgAV6zErYOXvvrLQk
uOVr9j7c1qvPR2mqSW/5RQPNTuMZGTPae1g7sRFA+RJcryqyPaAif0PI45aus8SK
wKSaLxxVA+/mIXqzfN5VweJcfribP60U6f6jl7+L4pdsolj1zOw3pC/Mkl/W1GuJ
wnyF2UFoeBuDDXPjHdcE7QuTCT6sJTNnfuPes+gSAXz3/A8R0rCCtzYaUJEh/d//
YaNiqzVyTFasyHTZT722iPO/gHPDLkqbTlq7RVKJxKDZMlaRyCA1rUqw6JEOTaUy
n8BBLJB+ctvyh3CzrWdBmpux95BnXRhcugNRSgomOGJWKHj39BYO7HzzySIs7s8S
iQxq6/GisY2lfyMEPKNiRJN0kBvcFoNWm7/nqNUxhoyaYfRqsrQADSIW3fBSjHsP
McAjn0Hd9iT4pa6Zgso5jhH9imMUjhDUxFVXcQO/YbNMN5sR2zoR+zL9shynx8gF
9+gKfioK1RlcwpWNPbjhC2GNqfFTjSNbODdnqOnv4bxCHovER+e8jV4VDeiSA2Cn
I6UrSjauRL8QLmTG3LF4qOYPsn+AnQ8seA/tiy/XCFvGMn14hvf8g1iEzjueJziK
Norrt/Ui7wrWfbGsX1cKY8WeaGjzkmQKuKPEPkPathxyj489egkzzLWbWpMm1++o
LFORKvWRVBC/5DYKSgFIXMcTwOl8JbpEHUXtxtShI2RZ0QfnLFmM+3zG0SidI+rU
OBx6U3gES5NTDz0D2LhnKjHIyBZvrmnfJncXSHCDSsKvBlIC4NjxctkFdZjisMRz
igTKwrcQoFaomsGvYEtEB7EFodtysK+Sc5D3Eq84Jlme3ddy3F/M2u+D6mSrl/5E
Jc4mKnJFgjUY89X0HgyLGue8/kmIJjiMvd8fDbMqRdBbL6o5Eb/SqzftgtaRpxQD
LbUN1mvsMtsahnSFkA8MNKerxmdbUO0Ot4SwCDeP4MxHPcbTe+8ZA5qtOlU0lBfg
3kzDuQXMi2WLxPiEBumdvfkZTErZfxZF8LJpVrxCh3ZLrgylOkxUfGtmmwz0sONS
ehaQcwYyYOCkmXVnaBO/ZlsTtWu1T5cjvVJpKCTYjTAV1n9ah976k/jOv67um2EU
geZmwL3vCX0Qc4Nl5jhnEU7NBEmZJIBMoUwpOMybLxFKO2K28U10qqli54Ri34XI
MF++DuTVBylTPz+4MHdFHV6cCCyZ5Z5ZXdQilhBRbjX6rPxXszze612S3PEoP7hP
ti2VLEcQsd4pjYavDqCQ1EVLdBzWhB942CpUswU5T/WMJq6SyKk7ukWjxUtRhVEY
j14tnqBPTIminy9Yp00pghwIW+kRD1AhGfkzFbGJY4AN6vthKw3w+DcbTes6WESH
NsDBPQX8qiqPLKUu4VbwFvM7eVA6FBBpQyezKN3nKSKBdkaNpZKjp+5nr1LwnzAf
PNjM16XQaXikLuXSC1Gx6CcTgHeFqIwHsqNdKBWviyszqDxWpyZMG3vKpYClLioa
W+jjxUcwf70BgBBkV0a4YzoKEn8ke6TDqVQYN6pfL7BztqPF4K5wy+zNzRR0YIxq
dqC5rqPgceV3WxTvNodiOqhVdJ4jHDrwRG1ju8MKV0Y7JScV/4o4uuzdY1CBihXh
AXRtZjpYkr4jty1yjoeMYk7FHk+1AnM5tLKv7YTyNKgWJCPxX63QN9648gieGWFE
3d70i7dQ+LiEQDzAk6R6No8AESvpT1e5VhQYu/2nibipU8eHRm6f8+9g0RlPBOTw
zIIITRU/xJoHEigGrw74mRNWkt9VOVIWR7QKh3XKIiC7s+KWG3drwMPRww/bECxw
JR2j0B0g9I9xcqslkNjyKJhUYdSuP/mEKOgwxVqjH3sQnTYCaSx7uVrJqa+nuijA
kDFS/QMdVYt48a+yhhppxAFSa2FAKvG+BO/qlXkAimfj9GiAM9uVvk3iGYRkzpZ2
8Ovnylx1ETzB1WTYb2WBjvoNlv/Bc2J/FxS94R8Zg7RjUe1du6bEFXi37lrMctWj
Gw5Hi7AzyaX+IV8WuiKMHkGfsKE+wS5ewNPpgVA5oE6U0mL9w6iT3sjwYx+OG+Nd
R9zblkIM3BdD1otaXXa3ZSyEYE1/rEV0VQVrZP9Qgxnh3wtddYv4aI5ydb7PluPX
iCp/6gl54oJ8seo9DzeDnZY1cwAr4/MGKM/siPPF2F7wXrbdb1vBGBu1cgdRFICL
Vfo7Eat6cXwloIqPko2AKMtP5n456WGzjZa2pkmejTccv9rF9q9g3XHU8viZi6Gr
k4yKiB4vdsrZSvi3W/78VdSS4Wr3+1agiOR85Y2oKbZMup1uEjiPS8w9PfMZcoFq
vs8qe7PuH5jbqyQCBa7AUet+S4vRqMvZ2K2ZV4PqyT2dHbvNsVquoIGKfyNAsLg1
wg3KJrDk9meKNybZ0QscEviGqkO+t+cPcp+8nW1Eo3VCw+wR6NPiZQkTSPh92RzV
G+fEdg2ELOG4yLw4ySutrriu2+cLgNNewUDa1FqHw1Iu84Hx9S6C+9569HRY3fNO
TIaKFHhdG8XPm4UsIxXsc7PGIhfzgBTVTa42U98p3zq5bmgNdhZBSufcY0m2hxoB
6DKCH6733lhxhhLU1tOr0to27bktlXWyV0IwpQPwUyzOdBRQGeLUSDkxRgAS41/6
04D1iwqAV9DMEYgyASblW0I/QgfEKsmrkFD8KSsRNHTPWQwAnJG3UuEomVyibH0P
PumgjXg4sscOc1ATXfxbBcbiVICS7qBNlxB0FNg/nsf8pybV4uhnUjgzvh6bAGm3
P8lkTC9p6Y3kQSw78OWMphFpV+mM+d2ji0WchHHLf/gPVy5/JDLoecdIKVrSp37D
e03s8envM+Ppg+yg+kcoDhG05pit7askqdUdgDvKntZT2q8f6KqJ3xbFmd+hgyzM
fdXow80wlsiLiGrJnK1YPl5qUi0aYNOuLgVXIWsNbwbDOhP6yiTk7AnE0h+n3lUD
`pragma protect end_protected
