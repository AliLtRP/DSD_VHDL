// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
AnVxVRYm6f/vMknUJO4hjGRiVmm5A1gW6NfIHcK4ZPUAneXBNKZ4ffVig40msgGQATg+e+7AzbqZ
AFEhF0W+5EfshG4b7E4BaXnY0VAjOPTkkVbSiG9By2e5Sb8T6FQWKOitFDCi6JerCJ/i7xthHA6S
x28qJ8JkDoxju4qkU94H3EVQOh62REgH7ehGjMj1THlhqBZslDlWuW7Q3mbWLwPfKapVG4fX+cZh
C2JQ2gk9TzHrvcF+qAFkAWFD5z0QqXC8cZfNmBax+qxZ7rXjDqzFvQ90J1TIiObGEMBIJXK1g65t
LGzyjRXHL2+KBs/w542lMrn+P7elKZEAfsrxPw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
vEyigyFcpc0M720PDLi+bAAsV/EdYIm/o99hdXkWBMxcV6tIMpJwsFrrSQYX5aBBI2hH9w6JOQgT
amwU8ScdM28R06QW/bYW5R1udNZahlNHOH5FoNE8fwdZSrvG5waomdKwosb/OAF72P71zTvcsSaw
LOMNTv1rq8oUaQDpY+azScXeN3TuixrhF5DP6NUN40TmeiKyZuDhz5689GqS+avaJ2F7StJ2t1K2
fE8YgpgC7eyRKNEl6J0W26wK/KfB097S2gx9vG+1wD87BrHaeOxMu3wzwviqOvchtZ7X8R8oFI46
c6D4eAC3NBG4BMY9v3ATtTa3k3sLKv5uCxQ2EOazaNx2G2YyekNbc7VfwDyqH2P6doRYqst93+V3
AYsF8sno3owQNZw22zQyArKOsRhWXu4WvZrSdqlVfbCCF8LJz6VTgXOHaUKhqPBwu3eM4b7XFGL1
3Yku701ykXil+iqBAQUaCivcgaThd295RSzBHKrTL7kWGTrbiCtDZre6RAEsMxP0LwVx3yG0pi+j
lo0yZoJ5AZUXSV5VdJS/ezjXk1js70u4QJpHBJmKXAzEdGaUFUWW12UmKRs6oK/QRU/p92OUVozx
/HG/nATRFrjzEfAHd4UzAqX2zXnI74wYpwjS07rYO3BYhvPqWnEduSgeH1JkEtgUbsd1JoSv/NIb
orYoQoCUEFI9MloCyF9q2sSJXcNVGUb2bPROXFi/Yfwxo8xxC/gJhqalaGeYz67qEzUc6LNzvNTI
kvq6H7vGj8HyXSGPEZ3DethPjsiIW/CNsj2DCNm4lg6qCLfb41ojF5gTXdesXXr7nYJn4LsVsJ4+
0vl1np9NH29XmX0n3pSXXKMRWHA5B2L9fU5hmwy6R+PbZG+uMvaXevXpqxYfLCysy31UrH40Qceh
mSgTeJ7uaDQ6tTgqFdIKqcE7cdNDmQVMUeYbuwJRZYJ8zcXAri7G2IRWcn9moZ1qhfiJs8t6aCX8
Tyt1/fiNQpDcgNmbvzVCIX2SF9IhRuL3Ein2402UXrkZrnl3RG3ON1/i+aO4BGjsddH455u3JsNe
I8L1yi75EOA14dvXu+9o5qP8g6uLesW9lrZIfI18E3ltnzjJLtClOQS/57yex/J5u9LuE/wFl5wd
cI+n2qYknQz5SB0YTpyb7b+5jVHBFQx64WbHpbr2fqm0FmIDyu+K82ycq5d/Avoql4u6JcEyw/fa
ukCR3NrUjqx/nBHw4TZDlxZA96jtjiys3atYgexKtlDLYznBLIR7tqgMis/Vr6P6M2A2TzmU1sLS
6/HR1Zjv8R3HfE2s+LJkMxfmr45VyCU6R6R+Qpf/CQeRGU0ofk2midO/WnPAER9kHAppba3luNGM
t3gmqVFXyegat+ElZcZDV3Z80B72/01z6u0H4lGrWGZXY5bILjLdE+W7RYBODLos7ZxtW92/GNZ9
HY8DhN7SgHSiMzMiiRni3O+DZ+2HsYiRq4989mXF1/tRpJcYOrbe7Q5rzS1hf1TscP6oB43lyXUz
WziS5b9t64T8GNIGsaGvX6aQ20Cjx4JFa5pfxW9jvPvulrmvbBx7ZpUnBWUB3u9uki9R3be00cvf
cZO4AnxXFdOwZ/wdQJpMrYxwlrUz85iCiePV9enfDIzLmlQwJe0HaRdo05CixoaSOTO+D1iQjpZB
wvVN3K7lT51QsFB7fJbOWuqkVIwazPo5ZrRMDQcFoaSI8iI44ilPtr3IiGQ2r1dRnJaKHUz1Ihej
qDJKpxBgJal3znvxyF2wod5OdN4PE0fWcpbAni7U0bjOr6/3+nZezFVIULPjb3a1Jk2SHoSGbi89
JkhwUQqxEbQxelqHekysb8UZCZtdoV+id4pnp7z4MZBd72an7n2ILmHRe4XxGWlBV5KzgJeuOixR
l+os14f3sErfaiW/hnz1982x4rADBrcD6+q31HlFWafsbJkWfXMAlLVromEUF7GIXhbJX/lIUlRP
A1N6Hd46lfVXW3KdI5ZUZpfQd4Kv+QhR8YjX61dFpr+evPlp6/BszHXAMrCHkvhdpzJwMsEvCKAa
Bb/P0GZooUVLW7TrGQOcJsOVtg6wGTWNsMpopxLjUOEr8AQXhKS1V8zDFCPc5h0ZqUzobisE+lqB
cmKvszvqGaJsVeQ0tF+CiIYcAk2RLUtC+aMfItt3LSlgT2gcc40vDjocZJ8r+NjIKWbD9xUN/MH2
ABUXuz7NfDPqu73pQCxCyS3zjk82zDnblJXRubr2LvrXovSM/FCcle8JEBBVQbm4RRj5qElaEl6y
lFqLl87kIWb3fOfMyjqzcGb1P/cSuuClykBAn1Va/BtPsd2DkocHdbOa+ORF41KkhUTYJDL8UWrC
WBXKXpz1oqcgVdAlR91CzjluYBApfybaSMuEGtPKWqy0Ab2XkDQIARnV4f9er9/duZlXzYa04/N0
+NpQP3y91NmSveoZ4iWUhzbYYwJE8sENQVzqaeyTw4RSiAvhHfF45OH7Cv2vnvayZNKvuz2EVXg8
3hIEU4xu78NQvf5XUekDEpf3JFtjOmbbRRo9e+0iDrJZ4/sGQeqNmnpiCun3lX8NWM0R+IoqDPcj
aFDJcr2D3fLedYyrVsKqb3G2yy1hwzsJHgJ82SqYUd92Xslx2ZGoZtHO5T7O2Fl5wYx/Ee8J92EG
Xn3m9W98q4APQlQusvuvpPibPB6L/xM7xq0iKC8E87LQEH/oBlVdxGP5n1ochpKVAV2OPkGpYews
uCUFLi5XEtkPLsaUm5HwmMXEYjg5Zi0iDDF02kGDJCjCgMZbm6h47WFyiF/mM//f/bOwoC7iMSIy
XKEwRC32Y6TqzOol07EJzY2kQAu4ZgpkUzCzxm4emKNjmZOASDwd7jrGYfM4GK1RZz1k8t7iy3Zi
Bejtr8lE8qjc1MSIiubBPlHt4YSVBBkIZI1lbUkiNG0fdpkMlM6cE2DaVsB0Jy8zSooQmSaMy5Nm
8hENnBdO2sQBHRKcoVaZZM+WDJANuCs5A1KmvkHyNhqD6/YycZdY8ZdNAeRZeUOVUBMReKPBk0TT
SWDabj6D9VGuSTyPj/fUec/+cllWNub0y0TLkYm6qUZnqYrRoxYmoBLfAJUmvXd9qCOU6Nm8ssWe
9cBA7x5tV4ArxClpVy8WDtgshaaceLOjVwSwyS9tETJuSks09B6UyTN4JMwLte5utqDyiCmNBFsT
bk7IwGDIVNSeZGg4L8hp74iX5ySFBFjZA9grq2IkicEHeGeGHnELkIVcvsCPsfPuKOi1FgLuTR56
Gq6MfQIpEcl9waUlderqoHvmdiHqF0I914oobEgqHdD07j0Q+KciCzYP7AWiHlkyXqIfVda6FURE
b7NoLM6QA9NywcSq2z+5xUfXTFWGKa9QM5oO8ccX3i7q3LgpP2uFojyvPCf13FYaWahnz7kcMc1Y
c90Nklpag1z30R9RH8z9wZD+uwGbgdS4b4s8gKi2Y+L4uZLFzSawUsW1nfM5Tj/EZUXxn1BuRMVx
fxRLf0gtxDHvQb/1zlEW8MhxtFc7rVcgrUH/VNzp1JEvrllMPUhESDvX6eZ7xzTKp6hgYn/Bg/WK
jSW3nVEdCWdHnF6tLsFmjNjIhfghqItCu1f7kri6Q/j/B2PdHVByi1nwE7kvB1JHH3vbFN73TruP
msaz+irniybhBWDZBCuDbqjBa224HoMIrwwBxH/M7xdvZ6fGSAIiaTi+LGd4Hhky/D/PMIYSKaSa
KWlQ8Y9g3OaO28qQTY+CpAFRRKzdG3NXjvg9uUW4l3vpukRA2mZy8S2LG8B74vULzPaidKL8lcOV
Huehi6+xOpht8UDDHcAy+4lI2gbUcNtM0cFtCs3yr3EylN/wMih9GcE6PPkbYM2Z/NseoUxg66QR
2VW8OZLH4E9OusJGjjGgUzYxjxc1XPcvFgr9lGXtIml5qk0sgin09c447BiOoaasHJkuR0+3AXw5
2VVKLOyakGh0JXSFWyowlOFpGsHKiz1hSBRL6GJa9nd4t5uCjcAeA2mfUY+dAXwaj9bUGzXaAz5i
tPwwVuba5mYeL1hpFCbTGN4A5Bjg5l+tf8njrP+9Tkl09MmsRMisHBs9sMjy9W5ckWwPabe7jcOD
gVRrJDT7M6+LPCk1Oimx+xUus0t0DyL2ZkDwlgdTqHZT83ar8xvBTONeB3+EjmxtEdvwtsp7vxAV
St/1//L22FSrxBbEE7cxSF+rK4fWjjQsbpHWjk4unXKCXeOOXK2PN83BfjrKPXvWJHhPhXXvAcul
+YYlsl4YPDz2tqpfCpyK1WX+DAffC1b7LZITZkDghwf4mOv4Sijo8mUG65RID+eBrjWnv092+Qh2
68WUon+00uhSGfjD1LUt9sPRtHhPH9131IB8qgVzEEjF4LafdO/BZOroAtf2NwFZBRZknzXWWKAY
LTnfC5K8qEdrBEWGBCZ09O5qaVw4Ce8meYaYHX8Gfl7kOXz5QyVl2bBf7HqGom/6kczB3BZuIv+N
o+s4nfyVGjl1nj2uVLvmTZTJAsEKZ7FA2U4kGhoVpQVwMNMW9FpUyTI6P3HWdznU+FvxYKSNjjp7
IUzZT8TfchGw/lSRpp/9F8EdbQ1rsRrQovu/ntRsK0Y1Yd7BU9oBWR+1R52VjRYtGF5RCYHvjVCS
pi5EMrntcHVMQdkBv3MfJ9fKav9xdcFWrvZlbFyU6cEXWirrdgq1XxrW1P1jSDd+inEaHYLGWcwL
1zgU0Ew5pyUOHy2U1kiUZ3BHnM8a5Ap0ejh7cOciKMiD6ML14yYlWAu0WL/9c4+qSAdnrUcr9d1Y
Xz04LRk+wIVtxNB84/HZP7eUJV3wGOleRxIbKNciwPbEcMAaCjWaBaeGEChkTUAfmOVfEX1UgrGH
pP2SL2DEsvfCd6pRKyxRMAgWj0HQw86uzIn8Em2YF0xbQIPbKYFke5p1NI4oiETfT5ekSQFKlVc0
/i2kAUyrM3UcwSl/XKsU88PvNJXjI3bRLGkAFSYjNfw1aXJR44MKcaBOsxdCZxjuEQPSNZZsqkIW
4HZ5+zuwYEal2KJHT4h2FWzPuXC2XKlo+YRkXOy5ykC/s/Pr8eMQvrzoN3hlgMAHW5qyxJx2Qsgp
YmpXgJtcoP3AcICrWcyakma5d9QTL7biEI+4s4cwB7dBpsYeIa8N7fRlysvZi5Tkq6CnhSjnzjZg
FFoTwymyQ7bbRFCYTCt1iOWI522Awxugc2Us2xbbMOguSUFWQTtgc1dKwssyMyV9IOIEVcM7T/Wx
InJZ8CDiVYROAmj7lOyPR0oR+qS/1YPU1vbPKazEUMk4VecKnNvHsAybNm9Otav9CA9muXbltW3M
useFMt6//ecUCG8suyhbBCNKChXHRfC99PuVGQSPPuHYh6ch/kkVsiUjVVaz+UHZrPeuFy4c5JSP
JFcnjJOKGVYi44LoyUn/OyzzRuKPo7S7d72cxpJSLRTzlz0VxO1W22dWRgfg2H3jTWmnl4ocd2f1
saAUq1SlDZVtr4begZ2tc4+7s2zfgQAfOTJ7CotHztzon6MU/I/Ml3ZXBbMR8nS8DCO7XCU2tgFM
Fu0jdGpWD+wVB12NdfsDjNb+V7whKcVpx+icszt9d9R8Tov8YuPpjVORJF5JnMxdpkQphIG8ZQEW
WIwZqNVEyrGk2WyLNVESgwHdH1Z9hRWYo+eQqKczpupa4aUFLz7qAdfeoMtqPpQBydpFewmbJzgo
Z615hIpmNy87SUeLhKtP4z6FJ8MirFBe4cZQyOUIvr0+v5j3TFycOtF7vkSpcJ7k6MRFNsiKxuxg
lbstyGpU/kB9aglDS9Ip5HGu8Mu6Vu5lkEsSXNuBorlQ8ka3wjgjX2ZCx08OTb+L2Ml4BaL4l91Y
oerOyH8E6b25yMIREsQZP29jcz/louHQp5VmXsVv+JobgNI3uTltJp8t1E8J5ngzrHHzzqgczGLL
Z/A8qicIgIW2XW987Pi+ecKwYIrm+7/AE+DskqIqjnyQD1jrGR25JH92mgt35dAq3Fz0TG7v2svj
e6KfYL00/gaOoAFFqL0cJgZsGJyv7vYC0DYj/n47Iy/oXbq19TlD9ywJwEAUPa+E20rCmwUw4GuW
z7yAbPOnIbK8h/dsEbIOYVSXdoflKoXhoeqY1XQ35LtcsQjwoq7glOcFp14ZMFP+/OacE85kVVoN
cjW5fEgZbiGTDvr1uRAm5sk1zZWVHmj81CYCNn2KM91B3vxD2SUsRnziqMOVQmxT7PxSJ67edfFY
XtY0IriDMI4E+vUWt9HfGuS+2vsQ0Ysqkh0WYR8xostCpc9yzJ+TVcGCMAHH5DplVgHK8NOu7WVI
brzXwxHoQd9GENyx/sIPDtV0fed3isSUZbVAwSW9/MJHYtomofm1nrukhuZR+y61yIG/081vYX/T
2igRSbNUjB0R7TxIGIIszjcik2VkUGaG9iSVrRc9b68cLxknQybDyeTvYrIPZR0YWHAKarqcYHTE
Qn6+4UvOvQqKycgOkraY+zHFfLJPuIbu07D1V18+05OzEIVM/bCJBdZt2B3L+nBcU7jydmUyGVFC
tTZdlkUsKOQe1Gexf95X3uXq7nv3CCZMhw2egKAMtctAETy/SsyvH2+VLtUwgwgd9diEwwFpCRov
RJKCYS6VZS3dlNae5e7KZRL+w9x81bHbBT+cPUZ9d3hLtpvEsMYb52nwLke5dX9Ca7bTkBwJ7hfJ
Y/LyTtOUAEMGrYHGSUmC07Iob+C35QAfkBc9QLN8p6kY/GPygBGliT/HNzoZVg3eB95aymdTOxI9
vEKuRhfUWMwOtr5c5XC0hQrEsayQbNP/xQsdaR/pmd0PdM0Uco4cunoa4NtDIKM+jsEqRwBIg1Ng
RZUaOWMCu91GgZ88fZxZCOW1GbBCJw/s9noKvEphqI5QvEb3WujUcoYLRiMfMI0VrFhSW8dtOaLp
gZoReEGR42Kiuq4fG6GvppQdFW6RBjP1UwH3A8OZtYPz38uvKA9dVRnr4WGXO8X+hBywha6Gkv35
P2oNmu9Kg7yghS2rdfS5M1KGkX0=
`pragma protect end_protected
