// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
UXJrgKJRB15R3BT2NOPnsapL4sM5HlPrG78zvMivGwTFmbnATsKRji3aod+noJzpKADfjvrpXEPt
D22tOnDCnrpsJM1zhxY8EI3JTCAFkSiFmLVTSG/lM+hjGI9+RIxEfCLU/K+6bnJFhsIAq6TAcjBZ
3qlI1qcHauPr6x9bauX490d8IZJj1y4mN/poEjB2q2I81k0Y8otgo8dRsEqxj1CJBngiwleaGBBm
bJ3nR+5fVC4s6F5bNpfEKi0Y2KnXUyOgOthHVVMlCyXgBvayK1ZQzwgC9CnKhBXQpJoZNLvowgEW
xCUoUihDYvaC3bRCSs9gBVD4gUTshIzjXUGwZQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
j3/whhF1Gl+Cp0WqviWXTnetcI+07UrycCqCy+yt75RnnT+TP/F13a/PxgR5ANJd7s0+QeeEftVS
AOI3ZcYHoMbgaNjd6eG7edmnaRxHpyE/oq1GHN9HdWpSqA/bome+Tyfv+ifovJuXHn9tT8912aL/
EdFFKLFFVjm3hXXfdCkC1UVumj/rvkN5A7acMEdS43ExMXFyjuWMo78i//nlZrzI8WZd3TzSfYZo
mekjDwKgNV6ZS3i9egWNmfVRo2m0eSQoQcjzjOcWOIKSK2rGN0EwyZnNJQ8qw463sADjzrJw8Htb
wnB1ahp7u82P5DDs+XbYDkxL2Daw2JWkmNbauimCMF64fe87VF19Ty3PqapvqJdzmGT5iEDObWl/
Lg4rJflSLtlqZm1Ti5wGWSofVSTK1F4nIXKCPZ3RvSWH72UQ9TSqAcFlado6KGsZ9RKew5mASqIt
F8WoBTznNYFNcVMH52JVuz8+HkoCAzvDUtOIKvVe1KrC8qDZU5iMdpx9qnu2ph/6Bskk0y03a2H4
1X9d+QxagwLm4N/B7dRU6MSNbtUNulC6LoaOyZtoJHJwZVvfPjZJVIKiCP80D7fnqajSCNn1KAxd
m4RxGEjSdX5Kb0hNF5BGwE7LiK6SjgBVPeLRZE70k5pS/UmY6UTh+7f+uSNI88yCZw+lkJnlZKfG
fu5W/K6IDhFZFnNpJ5rEa9yXVA8AVz7J3rE4CXUdtlmFohdSI8Zt1GzHi+bjywE0SCptKb+TT/4w
Z+9AKpMRo3wXAMilH4xQM7kX1bdgGJFp23GFsbC2pL0qKDsYFTMOdio6kENamVw8h08XWJdvtNWd
LwIh2AvCNAUwtS5oW9vEPkYvCyc3iLjRLEkmFswEfqfOeOrgek1fAaFRC9jMGVfGiApi0LNQFJwE
clb3LvWnADNpKojP8VL7mackfQ9C2eruMod9ZOEIH7rqFveymIk5UzqoYWUBygzJqEGyIfnxprOm
b1HOzA4PVovWUj2QR097e0EZBfbl8XnYilSAl8CMRMHbgtQoX9OvMDVSC70l/vhGaa4dQ+EqTHsq
JHfchpJsISFryMbyIew7IbzTf9F0OFy5kILYVz+yapObStiF9ZrJXjd4BpteUr2Rsv6pU43aK71T
5oPxqdCvF/uafd0ug4ahhsudU5isV3SUacyXOqoPnHh5u82MId07tq92OP2zaQtIXTLDC3CkNBiE
ITafPYO7xlYoN3SHguUO8i+PZRZWa27PAOJ4zBoe6IzWBK5sZbpQcDUGorImGjNX7E68/2eA2G+e
8vZ8+brIx312lE307E1OakMmsHUSJcpHITKsCa06rQWs7A97MJGL8vNF4d3z+TDmLZhXxADwG9ks
0ulL8k1WwKUdXpQEn6KVtFOu9b5OIAqwED8hBnfah618Hf+PHwdaf64umOD5BUZNE7FzGqMd3yEI
0FKnple+OKxUZYwRuwo4FkmrbuNog5zF0qkobgwjPOo0EPk+KQ3s+q25tPndnQWmx/dJJhK8Di4W
6nat6gZ2KWaBqU2W61AM2UaXHvO6sYkc4Cv0E65L/+Bf+PWePyQE9IzHYks6Roi71hWzh++gseK1
pNU9MMcltdhcWAp1R6Kq6bvTMNgYFCKYKyxmNWQEq4BmAyrVPOzuG0dYfKuymxhZYCKFFfAXSuB6
/Tv5bgChTo1IsrNS7JvqG4L1OLMBv/wRfs0DZJe0hgrSd+mr8F+/Iqb2piykvU93I0n2QFXxp58L
LyZTZvEwyER+0en1JFWFXxgjL++mcEfZu9Z05CPOZCG2sc69K0/GSVo7de7CciHsu+6LdUrWU76S
QHtq1d7p/q5T5qTU75Ms3aB06aK3OdIeSemBCr0KN8/i1rzqZVHQ9tHTjQ97AxkdWQ+BgZrqLDrx
K4GzS8Nvedg7FMS0dLKfgNID2Y1poanWdl1J18wtXP05VIpM/kBTCl9tjW701rmXvNYHNVo+OeNX
vCIVUjdF/eEKj9QbazrUd7lHcJTzFuSJUS57aXJB9vQkSM51KZUB5myO4D1TF322FL9kyYdYEW+j
GLAFuprQTuJ4LTL5UVsP7bOVzbkAIptnl7ux8KgIgUzy+Fkig0vFWn+0bj6cMa16CPf9N286IyU9
GctLdpqn1sDsyuiNXe2eeJpRKFkv7FWqq0UZy2CFxx7B1m+rmtCdSoGn6ddC4HRMWdqiQrObGcRn
ZyAjZQj/yxlxW5QeyAbb/vQh4ukWrmo9u9TP17h8fwM9Fug9Kwj2eOQGs2i2SXFiPghfRJH3ZYDE
/wDHEWJgCh/8KtSI8qyqtFuQ98N2HFYtRwUvuSUxEW24YmFcE1t/zZz0Y7Ue9Al5oLkapD1Ad1p8
2MduIO/CTXrC5bvF0Yn95KZrG4JwHArBelPU+8WHqe4XtObMu6nFhMwjoHms07TkZqwgvHJMiZxN
5x9ENrTluOpOMQQ8kFv10VH8Fd6KRH/Scj87+V8jEbRWSjT3YnyABlclRdXxSlYM0deO1tkfIC9q
FIA8xERimpta/42/PPvr5H4l/9G4mQhCgcuYSxPz7DNMKPYD7Vf/nt3tj2mO2Q8Os2riSa8i9Don
gWPEObdyRj1OIDW6ND36/CYmUGO2U9jr77yzULRGgUKoYp56pN60dyZoR0g2eGU/AXZiPsVsZfWL
MmkNlpzIwLr4duNZAiyt1bb2K5wHhLofZIJ5CaHVJr3gpWBKfswbqGcx/hMMI7sZD+EJZHNQgvOZ
fsFHLfBWSbuugV7+RT255FSHo3y9xUWeAr1KS+0SYZzKaBw9IAYeCIjTmM/mWpxnoxrDIX82/BsH
hKyIUTmds+EU9xwbTtF9BwTf0b4Vym6Ty0mvhj9P9rUgxZ692yIQP0tewmaJgs7vqceLgTEKlpaT
19KRKnAEMdI8RURbISlzY7iKkcS+av7JYjbzVF6RDjcW6stErfqY0OaCdltplL3QWgW2R7EMHynP
XsvgyeNQlfq7loosDX7D7/Y5qWXzS1xL2X/HOjL45NYQPGdnwAcfY2IwKAb8WuUgp1KwfMW9NxIk
iVNxR4YY/JRlD1dtydSvG9lGD6Chv5pBnL1C2aIRblHcJLwMdGePRFZv5lbEUAhX1gMUKfcQP6kn
+7t1CFHLOZkdwqKTtgXzPKMb4uB4WFqi7kyVTAgpPlsxv9HTOXyuYyTPqCgZzE8Ci0H6C+AplSvR
sYRBUv3fg566hXrXlHqvf+URxe231ywFIoMeLSeL61iz1zqvaXUWGLO7KKhut/3W0zXYms7Lxrxs
sexCI74dsmb+AZQWwlrY3mucb2a2Inu0Qh6VobJtyWushqo3bB/fUkf3S4Aqs0+sQmLjpCIX1+MA
tzlNs90W5SEmoofkvQ9/godZrbibypYD1rxisn/Yg1ScJYXSklnnlX7VuCDJI3PZDjz8G1ntlZEw
QvCSxK/xsYrjvTMjotiDPYGv98J+dE5dcTJpirg91gjPhig5AhaP4B82mwCJ+uiKmiThGH9R9mgU
Gd2kKcr/QRhNn705CoN2fXjCWEsKzaj6m4zHZPL7gMXVXtAXzJy1UkQ/nvj/fBPk3qnjIlMt8KkE
m9HOw0YWSzm/dxyF0hIVRZ780U2hqCjkBwolajyQYCL1+pUCATEd4bBD/+65ZiJWG7zVazf/cJOq
tZbosqqxAdwnKCUGkIuyejiEUvgsbelOxmN8DIoF5oW94OmOYiOmMd4F4zVOfgzfDP2YB1HzS2yd
DMOhDCP486byVYP8knplCMDuIK2U3hPIzKFlLpoxau/N85OQW0UGIUhMGBnhyix/ubFXZkiiVZ13
wrWENW3QxF0r58mCCcSU6N9Y6F4wYwNa8YXNCWQ8QZRltzfiBqoNjqR/OFu1vVTL/dSPmDuDDF0W
m82Gt16KrnQKlAd+y8N6rh8YTjXhCK07tZPI0mQgja2WaAXHkqjbJeCeGp8vS0ooC8m++RdYgt5g
70Ba+Q6+EZj6iH6HYp+WM+qdYh2DFUrkjOcauE1b6s+WLKiiiPqrI0LaypiMNvQrSDZoNiFvPqDw
T8STYje1acQE24jam9Z24ZsLKUsT6NOugGLjNKCIx8Up0pDCOszytAOPtBrdJfTn8B/ZQa4nimRI
lFg9nqOP2Sy0bG/03uk423lFcfbrJuAyi3VG7CP9GEPkVXjyMeOf3aLJcojvEUbLgpnaiR9CVu1k
O02bOk0W3Tl9ruL3cqJLZQK2FzYSKm/sp/vHj4IX+B4kUzEboimq53uKhV/oSwfj6wHUp3RwvQjp
X0sV6qJaQJFzKHAf2jH+JlcSvRiYe5qplmZvwYIvHxv46vgqFH8vI4Bi/y0l7nOJ8mDf279gEKzJ
etlpuLs8L9KSnaFt6fu4rOsYdHdDJD801qRBGc5HiXItPtBDMkvHnhpmcjLEtDtmMTQan0ql8nwx
mQWP1a+IBTIIYnl/2ERRgyLnTTHJr/YuiKVV6iR39caGbveGsRtjEQoc6Wa7pDzZtOIDroiWmHgl
+I7UUE5B8cMHsGCdY9H5LdYNl2TVJfz4G/sddF/3PGmqriWxjMf3aPu+/YM2eFncN6XG+uAIva41
ICkgSuFIlyDLDgU3RlruP8W+xM6kR39ex1quUOSGv30M3zoWcJS988yzZNjiPL1a+9UImSOXHr4n
MOrCuS5FO6df8s1TTNBi35l6c40kIwFj04j+F1gCr9u5VhtQh+Lnvkwvj3CIi+sF3EaaNSytk7Jl
YIm0kbpU5E19iGK4mjoo9QToD0QqE2aJRIEyzM+K6+kQo68bvvgD+zjbLKWdpb9l9QhD8hUQHR8C
ts9C2Ce2m+7tYY0KGIK+NuPlUSazYiETWgoqvg48tJU/Yfu294onmIiTNKH0XY2d5ghTb/izYYcM
Fksc1Lheqx/h0j4197ADgLNUBs1MVyPP/xk6I6WVoF8KwErbpswahol1Haxcli5D+2gB7YZJ1NfA
Y0EI41gT9KyQME+LOB+xXYrb9N99BehYpBZNMkIPQV5k+OYXnV90QxX+0yw7UUCE2t0hIcnttJYp
KIm2kyuRiHpFZ9XiGa6ZV5gNayn62swUXhtoLWQxn6/Ee2RzMz6ADqTYgZsTEsLosvHGhN/MDUxC
Go2AOISYOFbO/tSR6J01TvCam04hUkGo0Y6t1lg0yYmt7PDuXMF/wGA0rCS2m63UKTzlFixIucyV
ho1OpBJMT7wdLz2WudJ4sCKv/FjdQjceL5xuv92+G0ZqV4pHauKwaLAw5FEqWZmBEqcFmrdt0VzV
3M8rMvpMUu9JjkaiHP86eQjB69WSKvD4H7ouM9gV+gEbPZ5GL5MOEmtvtNeHkQrSAOvYHZsTfwjy
4sCY6/GSmbXVP0odWsQjTm2hUcxlCGgRVZ/GiQq5s/vlGxOCkK+E1jMIHwlid4Yb62sVJTDxHuzY
+5rBufy3IGvXO5H9vt8rhR3eehcOjo3mRCAiGhnRn984qOsD6ittdYtNjXlfI+IvfNHS3aUFShQe
NeyDNEegKOQVy/zqcEbfkNn+Zw5jircdWn7bga36d/dY0hRKCHM2Zl9yi6swIHQ/sH/9dVMIk8m2
kn248ZPsDoT24l/pTs61bC5JBwwAtN5CjZGMPP3tVMepr7aQLguU0b38h9ErsM1U9UFiG7YsIswK
q3m8t3qaX6D5a0mZLPHfbPJFoNc9b98cTJ5Zc9E5XDTho5C4VAJpH7AKcPe7ygPMfzJZ+NcERr0H
FH8sKseeg++vM+5NvMIfNc40b1xDdiIpni5ZUIPeM28RekeGxQzVL5erMYvkh13vhxFZhY57nmXS
fHiS/S0LJIfq57vyDR0z1P/sKmB7qz48zvAv4pnLWrTXfXLhNta84dG063gEuuhCENLqXgWl+5AT
hK4wjZm6HMsjMXjOXcfW03Fb9PY/RASm1EFGop7RekA4LbAg3g112TytowDoEwKPcsXrxvCCDXXQ
hXI85EduWRQbvc1m5konPZsEyqFIueG8JU73jC2fhuYRDLpdf/g+bi5HUT70kXKUb6vgPD/3/2wO
s442684m/cYgutyR6LzB/+H9ktiEaU/iW3sFTVP3xCM5YpOmvCecreR2IsdokWpvlyPzOa2uVcax
X2Tc7FtqZVpL9QycU3F0TYlnG+gXo5cAv6uSGlmzFPWoXLa/HvNPe4E+QZJntqsd0hNVUqyQy53k
WiG5z+LHwmTLOaH3er8A7jU2eeABopYjbhZ8CMmd2b82ilBsQXotk2OjV9wdKDHaw3Wy/MzdIKBY
tyAWR85fhUZreYtNJDeFOjFNZiiH4RgNmaA5q8nhcNFmEOPwVDkq1g13K5UhiT6Znll1z5g+0jZY
5AJUiXaE9QhetkSo4i05kzN7aBoc+P4t79MjMa4vG+n5EagRlIcJ/3vl2nhDU8xB/Cn6xW53P6Fb
k4LG/MAXVGp6ZRtbzOsVo9jnRp1m/EsywW9OFjKo3Dqh//PjlXA9Y0DhrVfDpGVgpxuWs/B3M1bu
iF5Kh3yjAhalVIenV2UU9LoHskylzrEz7nJx5K7wCqlb7a2MgnV1tbPa/kwi6RTyKkiHf+FEK3fh
Pje2uXx942F2nAdVQtM7AAR6WCMc2Ij51zE92Z3JLFmzHfgnvf2bOKQuJuvAF6XSPuHd0qUE0wwj
Ghnfuyo1wgwbzd31Fbn4mQeqD6TxscIBDxRC9xsaCx2i+d4OeXcoUoM5W2uSRptzGsDaCo9sl2Se
8mzKSdTFZ3DaQTpjk/dIyAcOGTuC+MWOBPxaKbbiwJJqiT4Dr6wP8UhQ+wxBlWwLH5WvwSmXAP1O
NcsbFm3i9ErslUexM1Wk8FEY0ja/I9RVIXu+vjODwOMAqPcXbRgYq4pPvn6yQJkUqnX5bVRxOpad
4Z2RZBONUPAn1DzTdZt5/XjEe3m62snFU/UZoezU8mMlZmILbi7PfpOQSScB1JLtTwRdRMh1b1J7
kvOqF6MjKZA4fnbmVqMARAkPd8Vls+9LSZ1qr2e/WAUEbEkz31DUwP3e5Mfp5d562u0GMfETazTI
ED+F7jK+3VczvDGSKefHrfq6VFIcLpcOkHtgxaDDVM9CxHqLXZpaajyXw9hvmWq/oSqp0SrQDT48
/QIiHJsEjMG50bvSYxXduUpkqsuyGcGh/wuKOeoFaJgdDvtWD/pE1O38/e+zHzxkvDozSuJzkymM
NTUuTsUVJgWgi1+JmI1k0xPRpPTPnDYzGvlSq+vKc20y5cXXleClAhyA2lSOhOdCrtv3o5Lwu1Fh
/Jq7sGTLlCgxoTWtPQ/XbNOya6lDx1kA1Ln46Ydl7w5TQfqK+HI/wDIt4XfRUpFObrpEIgS7LhGm
Or6MW+YAZdil+i552SdImm5vaIl1w+GuoeZ2/TEYNYGWoIZBKIc0a89mT6xQP/oQtmPWfqQJNQbS
WdlxCJLwwtSwlrYPkY/T4uMXk/+PGwdUjPNjJ3a2VLOsOCUq0j7km7Jx4c+E8xZ9pX/CAl7MR8nS
j0Ujy1JSTtxvWjxsNLZnfIXnB/5QcqsxwqeyKtbL7UtI8HB+Brr4ApPbJU0F+0AmZEC+HkRapaWL
rQtVWBg9L1xg7lowrxWwrv7rXo+d3HC96MI/j5H8KZMZb8euRtOtr23H6rroYGEvz5FCyYfItL4e
sa+01ecS/u8BZeqipBWoyH/YHUuouAcWnswJm8GqqLl1MC9CMNwULYi9u3jZko4yKrMs45Mz4Oh5
s80M/xwWCA+6GhkoprvSGkjCZF2+0RtOuVNbjH9ncrVVRu2jRx0YaJeMPgbrTGEgBusdKwWNufh4
cxISVoVPzGtKTz/acpzVZ4sqw+ByVtzIL/aHxxKFAgHrOv4kZ/RjL2QRxuMKRbE/kK6864CtbPOA
igimX5BrM2MqoveoUnJMEvXFszPIE5PRnHX7rLLLGhpHObH/xqO66f/1QA8SQ1P1VHLGQ8baKF0I
MilebeWdtgC3rjEXvHx0WBUb+1zxYJMcjvdJ2O4+GkyPiItHLZFGoZqS2hq822Ldn2jEElLTDn+F
f86awvLgKRwPIJD9OZEsmDEO7RKzKZvDjswRbJ1xz5rvOGEJOYHogdrlRSJnRv8IYZU9yLVFmDdF
Z4GFivyhA1UQGuyOpXhQY8+VEuq3iMhjfj/QnqzbPavG1udC6HzxrJ3xXHYv7WRrYVSZMWTpQaTY
vDD6LW9g0zfOO3G/oLJAYZZXQuyuS7Z9405Pxt5bDio3MbGQe3ZGMHu5UxrO1RwAXehFITUJNKd7
yGbr1qhGhlOUWAqizGAWRDKyX/nPDAt7J1x/l4QIQjh5pZ4nLCEygu91dACPK/GX8W2egZLB1pwo
qOPdMC1ZJS6k+wBhaeGdq3mt42hhXtLYXYLWVxxl57YkjHx2D+TfU2cYMEC6h3xdSA9mD/0BIe2W
mu2D6ZPYIn2Jo5I1DCV+IvEM9dt2+4l2ixKuCz1NpLPrniwzQgIDr0KIJpuSsb4/lQHHzshpRl3J
cpQ8wjokUhuyGAZdYi414KLyEyWw4YnPNNIuRLn8UtZDU1TBpQaCzDkFJrKhdc1rl1XXUTe0MlIE
vMHp1nXP6RxsV/rhJkwB+YI/NS+H+B2TOrWePyCu2JH+L9MiDNompWSjSYEEBSS6gjyzciFcEH4r
JOJ7w+WpGlBftE31RiL+ZQ6UxOGT+VDWCje1SbL8IO53UeAZhHP8yZJ5NfypTAaLoU6QrPnr7l+h
PS0DYdaQyOzqPsA67aQz4mu+dlvM9uxjmwGQ7bv3Axiut1jmpRVc9xSoZXNcGJiOvlqXfaAxcdnV
jN8h1maUV+kxHxErsytOzzKbZMBMrfKSslBrYkphh1Cck/kpiT/fRVrFMKRRstt9S137POuz3fnI
CTK/qaR4fPzPNf1pdNxh7NYFTDe36v/tlUGKrBJRX+uRd7/WK1v2Q67UokoblUPDJDqi186WWS2A
lg76/+clw+xJkL70oj5zm2NXUzK4Jkmec9EH70yh6+OxylRPLzXKTbDhWOU0rXq8QJ+83DM7NtpK
oKUXsswrB9sdXWO8kQRsez2ZWJ/rkshIJvc7ISsYZHog4UP/2caCCUkTasdG9ZnWnfkjjktS7WG+
HUTliM8+xCnG6LBcPBAWdtSm1kSrF1mZXsmbLDiRbdBa00zmRzCkfhLWNngK9qKWM8PowxyB2yAU
jdtcFGJxUQQNRfeYrOavWL5A//uw/zeFCKUUvJyphRZa6kQwiLc5CC2olmL6Labq0+w0Jmfc+oZr
8Qw832qtVJOymodISZPl0IMOP8w2h8KxzvvAopaJjEwOGjGtphkWwAQWSon1MJyzpUFuL/lPzpLF
l9Xa4Qmy3tedINoqWYe6m/v8E4SNOT+FtYof+HIbgvFkOJa01FxMBf62ak1ytAR106kc1fFcUVI9
jTs31gpuw2iX4+kb5ljdYJHHepYsnuLEPeGchQ+qFdokMCL5ogGTrx5yG/FxObW3GPIuPDdvI40X
yy3CLGmTKF/2Bf559ICtcOP8Ht88iuEnKy0PFygg7xfb6JnR6fDldKMmGFoUOfF9dzQU0h/UgSzc
iXvO99s0uNvL8xspIavCdXsBq6ViOV9/rewtebQD05r/UKVXeBhhHnYV3/JOwiY2a17KBeBC4AJz
TBJe3EZxui+b/qO2cLA8rKOlBo1SFP48Z1a2hmDH/2YVjpLBe9wgnYY5OZWOjlOp+4Cn0ADF4PHk
MkscCqa0H7UH6sdG0gY4RRT+OP4pPs3aIe7XjLycIK56BErP2OogmI2CZh5Ae68F+xhvU+XTaMjh
S//Ck8yBv73zE4+ZYY0ldoAAIFFSKOwyA1hVv7b3wMjPm0JvFhDe757GVdGa2IgyXsZPHjz6T8dl
7LH4LgTQhdsNsPu41hjFqUW2BmAKWFDJUI4dKCW11QbUfxOb+qZqM6r+4y4LPe4Ms9pI95WiAT2V
+gnkwE0sG49KBcU7fAzrdf7YdH5HNdOCgJUp9vsQNVhuKN/a9RaKzo/pT6gOMnZNF+00EJxMa8+u
zBNGBeGuZGbOUdZu5IUcybwHzKD5wiPd98g5Liun7sXuXDn2h3ZVCL9eABk9/9obgmp2hv84phsQ
W6frp7jOOqz+fQ3XbbKgkE+8VXEmgDo5Qza4/AIwkOBVeHC5stInNOA0vE0mGT29KXiD0F0x7b1c
NGvX+1jtyaobpq2H5Heio3fd5COO+AwPLzWX2q6yffkdRu5OMc2LWZwtf6nimhLjm1nrJnDsqdJ3
rknSQNTM/xlAIGjWYSZ+F3pAG1ZKGGHAoVW9yWeNSccPEkP5fJ/QxqFK2mUAu6/lAiRN8bQxETld
yCd+KEY0I0culNN4a9e5OQ9soVHmrL4C2KAXWjqMsYKsRfOk8Yxd4HdpD1Me85xgxYU0bOLQ7NGW
UozNUOi0n2gDvyMfZFkp7bN4NI8lqxamNpJNBeYQJjlNjkmrDcwaWKNMm5LWGIcZuOvZz1ERk2We
ZmW94b5HZg69CMAjSOtlrOIKUEA5yasWoOa8z+IUaJvuAHYBtpbcg0S75wdgiqExWH/sv8iAhuYD
lEXGCaFtdBWZrNJ9kGgrusf3QfB+wNmoBLIqFpWYU59dMdl27u4KTslLMMX3klZRKUkQxeL2DgLo
LYxQi+mdku6J9U10MP9UxsKZm/EjTq+IrpjogWLhfTiaDkCixMADAqrULKXEamY8nfndHyHklD1P
cm1nLA9dmL6UjhMUZequw2ONtSutgZJ/qSMr2wO6lGX8EBq1iSIIkxkKEoKbNYQlqRWuDuscb1Ny
8qT7ZDqYWDnBvGK4Nch1XudNbupsFT35P1Ym7LV3zI/WIIBhCh6nr3cTR19V1zejHQbumZuHtYKo
VqiCP4tRL35LmGf+fsx2lYKVSxiamAOyt9wdF/fFRjOyjoZhBE4t27EJuGTkVCbpIMUEqRIqlCs+
3w6I5pIKdrf7g4X9kODBZfY3gwEJy9SO9i3Xi2UXCVkxeTb/O7gTBI20Eyej1NOyeprCvnVGP46L
Ak1nw/I1i7OKhJPgFcl1MOJf9ka1Es3Pzwx8YsG54brKu464nli3NA4zzZos6vWmrwL9wMgWHCgx
J+m9JQUWpyKyLvmz4HK+WPax/mWZEone67pWRJUpzTBh6AK8H4rrF5O0dMAf0/z2E+yE0mdSdXy6
4vOD9/g6j/PCok9sXHF5qW+w7zY5qO/2hXYwW595/HWJqm4t95HdE6dPsLRg4vaPYYb+uYaqhWmr
+60veoTvrGrnsbVDnixVFah6b5tlYk/bnZY4wYyYFTilpv48G/LH3SEMPa8GcicB0YH7VO49uBpr
zF5aSP4Acz+hOnPYNn0ien0YxrNphwTt0gjmoT+U9jYwAB9Xj7YOmKKGS9e/in1oHdmtWd/FsZF/
dU7Pz0llENBwHAhwKNgTsdnw8dQGTSkJNRZ/r/aksa6uZys+0rkArxuCQ7QoKFMISNysZQ2dNDPU
Fu9Lduy+9cYeiFIrCoBbCrx5vzhVdcUcDSa5n0B9yKK7c1dRcyrXxscm7Y8PrtsLE9ygooXIW3Nh
a9kJh6RALiHlfnXCTF3dzSowlLJiLHfxe6+UnOGHOXdVy9DjSI94MnjRO0G0nJofe9q+ghUN6Jw8
n+uhQYaMY5fI0NulHuB8i+aQICY+VgmDFkqpwU66XUtzvhFR6LcjBQISmy8U6BAlVRyHVe0VcVj8
5qu6TUNfG+fgsy7Ka9MIPTUaTGVuoKDoL6euXarEyXfVvtleGA67nuJBdPcsYnVtgaPoR0vJqrWv
9NFyeK5F0Mze06lCMrGj+opVxdI/uPo67ZDGivnxm40CbfKHuyEdgFFfDRuLwOX4IxTJpQOoikdp
IzRsr3NpF/pmgZkvWPJ5s8IocloYuBmF3mg1H/i4FbshwtY8IPHKee64FrRKrnICYqKVkSB8ywUJ
ialllDP9mUstTKKrn5tkI3cUt6/ut9oACXw7UVvjJgZ6on3E3Y9JJoRB5fymWD3urPEDJUvQl6Sp
wokV3W2S3Sa62rBjzDLsS5r+0hh4gQsRZ1V+Xs105GyZzE5ZAYRD5Ok6ApLrKG4n1q6SYhrmfacn
EtEIzT4Hm4OmFAysrreBDb1jkfzg2S5YcM61QvfPaEh/QPnd5ndx8cWYR0VUUXwkUdOv6YthoPT2
1e4mQRv1xzg/MNOAFVZ4ZXQ8KCJt24tGJSFobhqO5cnHtgaNO5eYRx8OQwb1fRmyczjXKil2V/YN
oSPVdIg2L1GCWXZ0ANZ5rkzjtnqB1Ox3d62bLJELf+BaLoDdcoFxiCexTM58Xr8acT/PG7/LwwPo
WQG2+YUkEGD7ukwTRoERTcPl/95OxvOFJJHYwNNuPft6EOU9vmx9l/NnFse++mgC+CHMxH2RKvEN
0vGCrKM/cURpYNsk3LYoAAeNDeDfN7UWJKkhY2OPzU9TMLtAg0CM776XER+Nd6CCSxgPqMlyHl6X
n1+1BFhPfBpi02doJFfSdsvEylHiuqvOmvYrMFiTuMy9SLqDbnfmzfbUOhypb4ei7lP57INtkIZc
/i6SgPjpPm5M1wVN0J1sm4k1kpvroKvdAYvzbuwxe2Gq0YXTdJtZbQSObPN7E0YaZ2/9pKUA4kq9
niUetqydIlVJjT6Qe0t2JfKofUh2pB+BG8Y0Zbaawqr5Mr1Twin6EgSsUnHxeHsaY3l8bTVwaw4B
7t3moQ+NQt8O8pPl9UyfHJz+8iunsu0Fe3+64evKcJiQT2GxT5/9vgnVpI7iciBndu9DR0SCJ/rq
HGPO9AvWxX3HhTAKrTSsIAb2ous3K9SteleVf4eAXE0gDrRw9HVDxZBV3bid9JYsqXJROVUhl+th
6KFGUNSddSt4blajOvWsrer+xEDJ/hP21amR9PyEqytsZ9pcL/6GVrnqy6dGICD4+CzkQqTWb+VT
R4aaRiQwI/H48910F83T3mZaJK4DOExzS3nN8VcMz2DXBhoLCYn7bi8Jy7RgkCboEtIru9dFHXhv
S4pJ0zZsLowcqiT4WdP9h+ttsRSUr71k+22TmYOMXHlqkWO+ubcoVv9qHlYQETiV2bQ6Y8A1g62K
G7DPNzeYyFtoU4PMOqZCwGXdU2YyOD93rI9g7hKU+ujgNej/MM9CBM4gXY0kb7iVoID3ykiGKgjd
tOgqbLN/Pf+4xoJcRWt8DTBovh11HXTZ54OtTtkAZ94F1BVzi7mPQZqb2ZKhydIqCvzanOZaAioD
dYaOM2j/6iaz+giENLoUAAJX5a5RFiPSXYrwmGsy0JsnB71HMvgEEKWfY0zPg/jAwNOCszpFAXjH
fgANWxmSGLBMyMmf54hHiekm7ht5CzjbH/WEZiZYEJkXzvOOF4ECJD9zlatHhINKYH+PRx1m90AH
f3+mfmILK/7ztxd4S1UymlWzJPD4tYhg2RaVo7kLldfc+Li00h7CuKJZzhwYACLRmaVWlyrkvS1j
D3PVj+nnhpm+sSS/e+4e4ZkZPFVPT9Om995lsLP9fEPdseoBuHO7+o2DLy5pyah738cImvar/k8F
ElzGVS4iZL//2FgugaE5ucJ1RhMsZYml+L63Qk1MfUqI6ivvgaDXvPU72I/isy0cVR6+wHNVJaj6
fvJ65fyWhAVSNEiEiO9VXHzS8rfv/7TPJgIB1cl57d59MNexYJiVUDh900T+dLiwGKszLOJu1dL2
Eh00jjU5wKP72ftS6hNQUnlzBiUSZP5tK0H3GzA6AC8rsWRDz7v2bVbciOeKLxXLUJRBkmhfKiOZ
FxQs1rpMzTv8/AdjBa0LM/7MTjxmzzJT83J33SSp2QX3x+ZI/aCFFouC9wod6Hr90k5M7ZogmkhZ
XU9j/YxH3qU4nAT6rpZS2L1N2ZoGsELQsM/yc5qiXDPgmdd+jgS1HArYSIUUt3rqhpFLF4I7WRxO
lKywWGWoY1aECwU7oOYfcVf1sKUCojDfRMgDgKh3R0BZuZpi2FEtY1FYJTieHIuK4w9B/gKflx39
oSja3I0o22FXIbIODTsSr50IDeQQH+KlG1s8we7GqXXA2TRgPkdVx1AsASRZ5KywpdMQm8uf6Mmy
/z6KXo+EOLOjSssGXRTLVTeTmjs9sh00siHlQRg8oAVfOc70051gXDFpD+eC/m8VWvo3Qf8It2JE
V0+KxsXcEwhJZ1R7CQ/XxJWpMF4jSn/IdIcxrKszdEuSw6xmLer08itZqH1hdALOWHubKGbOnTWD
hMfdWUzjBpQiT8odCY3m+5+uXzyF3tBjjjDTV7hx4qqDYeeYLcugJIhigwgS2PSXxYY0jJ9x15Jk
0FonnGtOyW0ukKa5TqHq1Ga4fNoXVXqt1tksIc2eUqOlu6HFbWuAv0Bs+qMa0u/HZKqZWbYsesrP
trP911qZPPEvGRI4Z4efoS3qP7kRFzDbUVu4ChhMsSxRiKUWDfdKVyOALXx/RLSFmaezl/HgnyGi
OuynNu4kkArg3kE6TgTuZcgz9ei+muWbId5ZifFfn40JX3SINimsbMvsWlGDVvGsbS/dX17LMLTY
AFCgawny5FNLtk3no+Vh/1KDmNEmWN1D+z+7GzO8OoRM2ht0IVL+wAiZkwpQHru4D8sNLEyCm+y8
BpboPLO+UJWvFkHKTBK24icK13CuoPF84bjX9IAoaxQC63pJr5l+IKNFOE3lZ3oo62P+neij+3ym
GQ9kkw8vdZxd7PR9DkTXLN4g21g3qpUVVjdxVm9AzDNVo4G44c0MFBb3dYHs/7JLviNe8XRakeVX
OLK/VSPezGmztL4LmfRmVrRVpYrp9Qaq1luu+xCVRJjDOjYDhorZAz0HNJ2+3zxr2hyb1Fxq7KQD
dOs360uAQA+KeC5DUpqJ02RQ3kZVOrf0af9WpbROMW6plhkkthwinPd62BC8HiQRkfN84MIg0f8Q
1l7yz8cth6haRCNEOnQn8j+CEaEkxJs90+dEmjRp454AWBonoXRh7k68OpeSsM8OtLT63NcGD1xJ
My6say5gxx29ocGmc5GHzPmPFbEu8T9mahjbeQ5f1qroB9eji1Ug49Zyossq+UdPLQRi2R6yv0v/
BIjO2AlqOzvMB8+BBQFpREj1CyhwOB1EV2f/hx7otEFpuAqZHxIS3irf2onVf/9Gr1SBztQaBNOc
nYJtMTYHunPJStW4QlrRkpGiu//3F2oJxOi9CGxX5CYK4/Tgv6CV9UuYDznbx5yus2jAVCuR7yIG
u08vGapHirRU3sQ1eoUSILKeF6MfGS3DYGQ7UyU0BQBQwMtDSp74hXuYO3ORf6CPhwpAx1a5DMpX
iDcUCk1EUck4vudUXTXAj0WSg2rympZaj8rs3sKbblhvwkB1NBjH9y8UgHgwI4TJCATMlBhaoO/I
N6lkDXqhIzh7Rqzjf1EkVXElFL7VeLggxKM9dQ8dJmsdXs/zO2+Sziw+9N3fXgUNaoC/7OjnP08D
7sx7OObhOA5HQ9ndAeWvqoPDTSYEJGGQuGZoqKkw9IQvSM5XPPDr8NL5sA6IfhyuuNdhIwufxcQ/
BEM0P9N8AYyPyuM/AhyA+ZuZE0dncWGu4UbjrMa79KdcjnlDFclzRRldsC4C1HqvLZ48SxCejKJi
DUq9KVLGc2ELnNLLWnIPc1RD1lAuprIzNTBsVfNqdzK/Shk8jjrLqh5RVd+fGLyCv7vHQQZK2M3C
6S/p2RGf2d6HKP8L1f1GIb84cfGZ5weBo8Wx1oVHb4bFTcwQE4MdI+kenenIviJk3erjgfk9mhZe
oRNYYE3Q8KdbG6XrOZeT9mk1evaUyPDPfRzkGQvCFbl3qD4A4pyFC0/96UloogdHFtkrM0c52sLF
A7EMFu7nNG2Lz8Z7ZmFng12utwarFnJSIcX0IrqsgrMP3D0zXleLtQoOPd1Py8FLwOSFk73CdBf+
qYTRqigX5WoNkyXbN9mjfSHQNgImbKPMdkaCVIHuMezkvLv6ZoGMP1aahEaEol9jGze0OAyEnGAE
YRIsoTwzoLSt9xN6Go4U+q82lWe7ovYZ+Qnx78jpQmbZNV9mToUNJkIpo2rfxhfK4JPNj75JM96E
SzZ7NXGHXI52DwIeT5Burz8x9Xz8tmecSPUwBiek13xHOctdpUdJDjMq00Xn+By0GCcqgS4yXqif
VU1iYk/KBcKdkp95gDbpbni8898JKGWSv5eyRfSdcJXh0ne7+weZZQ6O/wJXMPLWf05vRvKSuB34
/0u3++652/fneRC/KTu6QkHI40PmpmYwQJynyvo472lgtoslS+i6VYAmVXfqDPsNlJ93ahscEQZq
m5FcoXTtkAAclwuJ/SS/5fTjqj3Q1Ww5sgaYcWCi0YHV/S/RtlSiIwVB4dhXqmSPhudgDPcG1jh3
3BffZrvww63YsnV0+GIcBRfUrhFo5d1V8ZKqguRqbn/jUbY4iDfkvYqSGFSVgbY+kIFtpoal7boK
LtxP00T2WHo2krlKyqUzqKYv/llGH4WVJELsP48BmNeVr0FBaNK7BlOE+DfUpmn71zjIiUICPoRy
b/3CZW4hl0ORL9ZKM5kTVaOfIZVFkQBgb3Az9bCGta5A1qcehEV1ToHOZcL5Uqw4R4fNHSiBgXVm
TdlB4Owme3QPczhpoRSg/6u1Agmr8qCRLNJ8cxF76xcsuRYUScEljn8LfRIFioVmDw0+D2qGiOSL
X33RYvNo/Jnf5WVUU4ok5Nbhx0gHA6AM+bEgG0W5m65wXhoW0KmRHtrGr7/IzRf8rSuNFi4SJkmJ
BF1cS4hS9uxDinjPtW1kJDAg1A+NSVZPSU0Xu939xe/+UtOVF1tBMSG9z8NuqqkD5UaAUPgEILEL
9s7fXqskr60Ewp/Nb0kSOyh9y8IiE0ie0rtk6vBSHePKZwJXCxZHuetwUGtM9yf3+yTOoheGZRvF
rvwxmvh/l3dwwmulcrFH3AxLOribIzhH3zhZTmdyE89JgGwurKomfXRHssiad0nRVnHOBwCARCVU
alH+eekRmAaJOBAVvEc7nl+bsphE3GnYwUQDlPJ4Ruds5ondckGL6IY39i0ZdMI5xbptGfdHHNb+
cEl5u1ep/RcShvGhsfklYEhJBD8OrGVXFyZ7Lhpiz7xwKrRiHQxBLSUk8whVuSf2ovgQ5glTPoXc
PZ4Zr0asObbFW9J16D6USzyFpg75M+7bk6KLgYft+Z38BnYIyDaa/aZOxfIPfZadZwUfm1oowTHz
qw2NjkpSE80got6lZwtyE3U/B2LZNZEfDIPoHAfOJmzgTYMRwKT/s9gH7UWZG0e9tQhJSsOqGV8E
VAvmE2GGnWveTxhvwRjvLq1ujsQFVruO8dHs1X8/XQP1wgrDhs4bUGhNGDXXWzscGE73vkEVtzYx
1t8OXl4j+kHvoRttOi0W7Yp9KdczWcYZ71y24H6lGrpjWxGpmEfgjItT630Rw1rTCgLHSLHnAliT
95JjI1wuZxEeI5qeDHkZ7Fmwq609jaIIokOv1zmbILjIFZgZimdRhLcnfrn/06OP7P0Q7nGsblGc
hp58KVfXYnW7YpBpXNMQnH9F0TmBXhVRvxjacrN8aP8yRT5gatjDrbBp6JV1itM4WJ3ABACmxTA+
C+vUA43t4g3UVe4CXlF+xP1jReZexRzTATTPzil6ZjEGUWNRGNDt4sGi011Iwub4BZHAcNwUS4yq
75sKSWtU0jQGhd1US5CZAkS1Nkkntc0kNBwTCRHPE21ipfA9JHlIsyYvSY+7eCKus2MIzDeGVJxH
DzsXMw4vpKXagT+44k0Byt6btJv6ZfoX+PLlu9CbC34eduzTjJBDecePXXIVUm0cxL5zq3MQHUC2
SzRuK28sBnVv8ugDYk+Booe4fvuGhBPUOENLJusOe1U1JHMHsCqPPduqeCLarSd0OfK+w8QyOPbF
6M4Yv5B/OhiLt2pLwXSQtXx3JEWSInqPkPi0m24bzTp/AbCl+pVk9r55Slp4aUL7R3rS+oo8zcxY
KNvEuaKtgRwhnEgnWhpQcI4NmxRYsAvnL3Gql1hN51xD1tI/qM+vIoCPtkCTQlWyU+nfthU8OTGS
P9X0V1ydkZkAprlLhN6o9bGz23m63FL/gBnUXBgovRFpocRVJUBeUtrTsj+OwTiIXobjcweJM4pU
cNMA4Zkmn6hsRx4lMrwhWYfU7VSkcORl0Wr2BPPR6YZwXRxKjUg7RBi055qJXMGNMKQG9hvtH3BJ
oKtisa/Ik25yC+GhuNsjp2odjFfHBaDN0Smwt6mk6D4n5CxJFwrxnzz3ivdmqKNSjUNPdKYNCQqI
lJfeD61R0OqKCxVcdexJx932ZyIdD5DGVPHn+z49PZQe5actW+M9MiKCWmVHK/IHqB9r/wYUuV0n
Iw1v8vk4sUspm77XDGLk1G8PpiHhXOXwwYh54EqnaWMmPsW0ty8LrVotgxRC/hi9DEM1yU0ByvEh
A0VGgVdjFDni8ivDrZ+TbmbUPfZaibjqC1DfIrAvwBKvUMzhaRwKxyGidYmNGC3DME61QsJqt8L0
eKFaa1eh51cL9bLVv5937eI/B71kLxVxyo2m8e0hVz2qDErK6IjstMetBro64rC9rSr9PLjlAcLU
DYn+gupMTOJtKoPL4FdWZ9Ol1JT2rkIsqSwlUqvvbTnwYd88ALtS5d3c+cSHk/YckaUOgUDuQH0p
J3DvtfVA/a7OaOlRr0MKsZzaBBQ7kYKCyVdQCeLdHvy3TvnD+pvHMJruZr58LujtLoK1Al3/HfsC
ehR9IddAmscFAHi/VFSHhi2kOa67qByncrgHoPXz2CifEaMBj8+HFiiEt9PdzS+LAaXvKeZoW2Yj
xN+TWs/wCwNBwWeg6R9q0kxmOmsJuztlB1D4DAwqrV9Fa4FS7xDX8mhuNIDvjmRq1LKXyVadmfc+
QY7TVpaJCTN6g7ZK8ctO8yEd9gKP6HuY1nYXbJkj8nabhDxpCUEcrmlN5rcVy9mzbokoTYv7AUCG
FJnMQNXY89QwwxBukGVhBwi0FU29CtpajmcTxpkZ4udGOV0yKUoumREYDPmA/0T9lZ4eSjO1qx/b
maJT6Z8+8xJ3vOhmmZpHCeW7CArtVDhb2ZFgPGI1DNnZc56xidSeQTAHxiCclWOZChzcKl7r5iiP
gxmifMPRrQLAY74LdTXxm+W8/m/uRNRZEBb0Frk3dk0xuKKY/OeAph4G6nITKYAY4hsaWH5QdI49
Fr1vHcNNcYznNYXu4yK08lnvM+fqkEQOU9+OcUQPlpenUeWT24sUgCEhaby12lx4IoWsEiRgeO4H
BCzbALg8QsJOfJS1O0U7OJYjLn3IeZgs7PYI+S7HaBh2oukctlV6G5otTwLlLeStovuKhqjXnvn7
ruAtLTwYLYrFKO9lP8y6GCfbuGW1akapb45s1Kh1TUCjPFqj5YixBYHilia9ZLZJtzW1fMBzlZ/u
x/UnebCkL9q5nOknkoKZX1YukC9q7xPxFk//tIIw/jwO/bW5/nDL0iyPwtkv5TB5zeHhla2NYor/
R9pqAjO8eIOHcPRnYqe/DVZ9phE5/jhbwb5fqc8c5Qbg7o+mC6aksRWpSzn26zjNxstgWb6MacQG
0ToIDgvKNg/BHZljMpwoy43mq8PM2j2PZuByzdWnUz2znAVR/7X0mAZuzYytw8lIrqaZ+54bAMtA
YH/7Sd7QKJ4SIM0a6413SFVdYG9RXpWyE9k0X5Sg5yGjfwfizP/GHggnxozG6CCX9j2tH4Mss7+3
vG/4yZPHRDD1+S8lA2kkRt0QkeQOXQvMqQI5S0a5iZoz9WPZoSZGxQXk/uUQntVbMlCok1/EaqkN
I5omAX8A97ZUCm5OOKq0v9L76JC8y+SfThfjSnTBy6ByuHl467orx6y80IMA4qKWdPQ2GyQnVD6y
XN/0gECZis82/mwZ3ZHleI9W1/e8ydgbfH4KXHCqqwbLvglzxBMBqT/PkPhd6nvcLpYydHFAOQGO
awV31/C13ypNV+SMNfzRM7xsLKZZ7N2KclcDDn7ZvGTKxjpsiC0Tu+ZnByZWNxBJWuy6nJYViDV/
aOnZz1BrpDharYwU0gLrX6TeNU0h6m7bOZECJm8Q+PRseVYKFE93oRmO7lt4RVTxuOuJirRCqY5q
ReOh92w5V1P7BB36gSz1RlI4RDkjiNWvvmL7NKLiGFd/Ykts1uWQ6DsP6yMHHIUdevuelw8NN77z
qZm5abI05IlNz5RWJmDaB7DHLV1WL97WAJh+HoxT06VSKjb99INGHS3/YMrUNkjP+9ENuFOJXPFh
ZsZ5DNgxWsy41ADGWTRIU0B5ndbgOt16O0ofes+3+Yix5m0KFnAHaXnJAQGKF+jH5W1tRKPRu8du
nkUi75SdQ9r8JEK43V8xRREbNZD6Mww46CulVfs7jJLR2S9+Q3FWqM/1ACtN8c9UG9tIefvTyjrL
WkUwjAr3+E/FJDf8sKJKPEOYflxGnN9/WmixaJqyFRNo1f35dhHMyFFnlK6kbnrc7gcOMY3P0ekU
lQk6QqLJu7JK4IkS4xSO/865+qEUkJwUbITNIKGNZGrRl5fGfqZE3SBfPwYZnnmdFcUKtCYUUtf0
R6TCNpMkqbQmKcq4Fw9iTOu9NcIW3+28OAe7f3QF8jnTQXDWgg9agTng9z0uSQwdycE6wzPW/qt0
VmrU7PW3xXu5SGn8G/e34EJ5pQQcKXMw2O12XwqIuAL8y2zVTpAZcH/fAO5B63BpUAiT3aFA3j/w
9+n0EkROnJO0A8ccBjvIaNfkTCv2zjhPxxRb5S63/Dx/AwKlYaJDcoSv4JFuLpCBSJUuiRN6pr/b
7xXsQDpkZivhuRJ4ZidanLeRyv30e8HY5wZwtE4LkTL5lU2Fv1hapvoyCXjk8AncpjXsIyiXZL+1
BC7qSg9t+UfNXJ2ZCPUm1FbNSZ+IvPRlMoMVxkef1JbRYHi/JqU1byQPdQJlHmAUY+b4Z5n0ebUW
2YyygHTAKqaedyt40kDDr2uXgkihHWgO2Lf1fVHNZaXClGofh+ET8YjbILgnXjxxqfOYzwrmU5rS
HyFSvSUJBPV0HgZL97sMW4reb19pWlL/gzWd9EbKH5rCzp51VboWfUjTBxGeWhZK7WCpIHpbeTOw
wHVCNm2JhXPOXx6QOs1m1n5vrodpBScAeOu/r3OE6FQVxTECaHI/2UgJ3SdQZZOfu0cM2qbgYp7Y
VqY6D70vbSLOAubZFtQexR067wAAL61utu+FHa04TWXSht1vrizvsMp78HzqoAbSALzxe46MOL2E
oH561BZkiUjym01fs7/Vz7Dr4dTCJ8AQ+GwDuW5PtlcX9MQtUnGUuy1qs8Xpj/FDL5VDw7TvTTgL
HKF2nSZfJv58rlqmFlCLtt+MY/px4vIjILmGBOo/P2ohiGYhze1qX68FIIOUYZ675bVp1jE1R0dT
0AO16/0LB76SMYNpAcgLQmmCWJjcnQIPIXrSrUUh66SQOQJNMmxRWoCjwb0UC38vQisJ5DiKoXrs
EOU9FFRCz0G5R0mX3J5Sf/7zmZgTD1Zw9WTamelJ9kWee2ce98oaHWk/0dDjYH/WTIidiax/H7it
IDJ5PYM7sOmYwxkamsv08cGu5hNy3VwP4Ff1/y/AyGVSAPxrjfmEWRAC5PgmJbFtGjbRZlGfuyUn
jCqT63j2rvBU2bKIzKK3O351ZOvGGwx7EaMay9O1g2EWZ/Y/jrf4e5Mj/Ug+vh50n2MUGP7C5RhJ
CQrR3MNtQ9ynAR89dg1NnLxi3KJjhbjOjrYmtS+yTDN8Y/qBhtWyJV/vnce9opwfBg6eXc54E3Xk
ghS9iv+BrJEz+IbJdzYRoFUqCGC7zzsrGnVOZcN1XVKXujefw373H6aDnAq0dq1Q9cHZFSFQnjM0
f9cEBnqDwhSZdwjnQLWnkkFUguJxNvQmIa8V0yT7TqDQGzQqX7bwOu36KV8OqFCqnY5GtQerL39d
emC07h/Rbwb8Y1U1+jDr9dVHA7bfu4M0RJ9+fWIrrmB6jvNYpXZXRYsS9vyYP6BJp9wLgKo9LCp8
0uekrUtUgOJXswKtezJ3UgINTIoOiv37BPJH/TpH489chaVdAJKk4CM971pBJHKH+6PAxc1VVxd7
1MijlztejF12ZNfHoEa3V3ANFmBf7ICUiPg/IcfQDk1xqU8unrGclep2lEr0SLOXQQl9T05u5n4F
VlHPpgksohbkTOM47YLS1hcZIIJzXQ3NCZPHfR8+le6UBixpxa9dZX4Rwg6ELWFFHvhiJ31aYefq
bOAI0c1x0JgNLsx2Hp7fzXJZyDX2+vve1e1S+hgKVDLpTe54LuXOZLUA1AT2GNhndSg82l0wiajz
SnP3ZzZE2jhj1nXQLFXgkhL5X65R1sIexr7l3UTlshckFTIQqtSChHejq3ug2Wd/pQRssb4C90sP
MJJTqg7AJET0H4irmmT80Vgee3vG/hHZxF+wnNueNm6NzZORi7pJULpFQYFgRkL6u6cmCcEhxOmX
igfaLKIhFXJf2zdKryvxuDDfO4uDw2MD1uzBAVXZ2DEOW0Kj0Hz4PTv215PCrCzUp6pLFSZy6gBa
FLQ+Yz6PjLoNrc5V7vrXXaeZM8goijYuPoSLt9I5R53T+IMhSkSEiO4qNSYoUUddLaZws42dFN6M
bMAVgPcOwHwG+uUhiIZsATs3Qoxut4d1iZAaG2Fi9fWrzMKDbaCow4AuwBXmiBbQCzyUIeWMkQ2I
0wwHOfdqNYwrfftqRuPS7yYydJLNi+hkuEjRHXtDKatj/YsiqirowfoeI+QFKGhgGbGQGgZ5V8J4
1QwMXyaW9NiIxfheJzLQb/bjDyWNKs3kgn7FxYnmTj5c0+tvafZaOdQiTOLURgr8/gNt2uc74VeO
mYZj6FMEz7zhqdm1G5gPilNrWHvyDUL8tjLq9AX/Xt5NOiu1JBkFE/uvZaUqq9TXSgMftbLXsjbz
1jljGgYra2KU2AitooFHGslazzWxhS7eGeGqREf/1Q8/sDbJXuQqhLttCxBiAUOB41UlHOcyCqni
CqPPcKij07RL2Q2+xJjtFmDeGhTav51hAKLvtYFNYezudEAcvUNLAJ/N+G/wagi13GpOPE5+yHET
+8Rauj+qWnUmqgskn2HJIlvAX5ZXuP5rvQcUrsulECx8fO3FdGoZzuuICEQ6c2ls+TD1F8XOVEJ5
K5/v1n8niDbd2pjUW6pe2Z2dKtsajsESU5jjH5nbnHvWpdG6DZOo9aWGwGT6g8mvbJLk+yNs1fRg
crAHZ4wJntDGZTyimXYBoh6zWlpOIT2kHDd54s6R/4/wdgREjS5YRKNayQ/E2r5MuaaKHOzT/AK4
E3KbzM4G5xA6ASPjAmwVPHocZCFcSrWaorj6nFf3pBw0AkOYgnhp7vKpizs19LuvAC2hFR//DtNp
f4USFJqiQw34FS4JvD+elcsnSo81jkn9dKcNs7It/iwztw2nKVMirHU7zUx2GXTvG86K7/erG+7U
L3ibwPYOUA1o7fBZ/7oA8H39STVKTnrvORJQIVocS6t++tA8WezBqDuZr+ao5H8REGH/GGO3mqSS
UNxW99ooIxfmaiYVlDk1esaPwjrEC/9Ry+km5Egl5MeWdOl63qWqAxUZeI2LO1VXQlaUGH4+Z8bP
rXni4XiyfS18BnGjwhXvwSkJpcjef6y7yGDiMrcmKJXYeoS16H0KsuqUrRf8xwbGls8leWShTb74
cANZXIAYkQivBKm6PAen+4LSYpO78XDV7TLJDlXNQltreDYGo3Cu/5DcGCb/3mu/O5Noi8JSzuGy
7pAhxRomnV2WALSmrWXupB37a4rp19lTFCM1e4nBsivK1vD7trDfTx5E1zB+KzzDQwJ/pL+6zMP2
OxARZETTL0dhLpGsjUFGWeyq+90EKZHlEw4S8djuBdzsyV1WwXzG8jI0O9Bsj1Sm/8v20NYo2j5w
YDCfcM3VSMuHDR0d/vizxH7Kq6LFRS+diT49nx1ex+2hoDiCIVZ871Sdeaqb3vpBqOszgZSBBWB7
KjumcuUfk+2sPKh1IJlZ7XpLRMGZ5eDYpkW3blBZ4CDOajvq6BrfAETzbtuM56Uk1c8/xt+h7i1Z
NlsSy2Vg2dRaRva6JwdMx+LXbOWxZh3h8uqMqLCqOUioA1bO+84dlQMkjOqdEbYMcJZOXuAibySN
7WaVCkpCh83CP5EWm3znayYwb6rUWB1Yv3+9soSjUFhZFOXJy8nZwFM1hNshmKmGqtY9DLl6FPqq
v0OwycDfXeuDIIUx04mtT5tev2QNTTeQZJBq4Bk2YAj0hQXPKQbXMG0pNjOGqMESgy9MBok3jlYM
R4CizPx+vgeDzmAQoMPDwYoGqLIowkR2ZaEFStriCkzLYXCY9BArNAdmNhIghrTAPMmTK2VTxCLM
Df6cdWmxUxr7vooS9OFiAbV4uZ1DH5ZCjJBDJxOfJDJjM1wb0ku2iF7lGxt5ABSfk2oeJDKWhiXq
buYVKrvUz5xpWW4t6gDfFT131A5tjJ8C003cx9fifujhGCg+iMWCFoNrBJRgVqwQ9UYFZI5WU3Cd
HvVTdtYsMuVh/Imcg/vfDkVa4Ed0Qs4iUTcfef5cgN+6n4GvT8+p+z6n/OIKl/0hqP7yDjxjAs1C
4z8aIzOcz8xurfqMiqMuUk65Wp8P51fvxpzdfGy4QhHfZn0way8jKYuK8y+a+Ln1rEG8xAE4Wlir
cCcD3uBzoC+u1FXMBsjGXzNUjBsuR1MP1oQ029n5Se7pPlu5fqm0AgZ9WKLwkvabFJXLuELvO3LI
Oxtcd4jdzytXGBtSLxSGt8CnPKdJvcZaytQq7BPEn3+yXoRC88CYT1TYzmVH9Co455d2o5Nfb2Nb
tUUDL7+km8R5peroQaXxQBNEp7HHE/GpUPccWBvaoi6yGGrVDROGzSgT1h0wE+wwIQi+UZExetJA
uUzahm3TYkePSolJa0lOe79fg1UCCVboxJvkpcHEC6Fc78YyhUn6Y7a3NgAYpyG5p3HfznDWArNy
tL9KljepL0T4G7EM96D0MM5dFbmiB23k4bzjLi5mFbQvLUmHxYTUOd6NYdIxzH+Pfjrml2KtLySY
kAp9zrO6lcOWumO2zt5rSI7W9QaWU+FpMDHBvHZjAX+hFtGxWkIK+ZJq6nCWdWoxVg4Q8dk2KynJ
OGyP+RRE2jW86E0zceDPjc/NdYeVs3yy11j01iWfpqCVJ6JZdnFYgqVfCVSMrTawjRp3f42jyxfO
L1TcfyeqprlePzX1uOor4aw/tMJAlRkwP7BwBZBYsazoT8ObT7vFoQ6LbC/w+W0sNIQwbP0SwScC
OJqBbE9kziMM05xkxozze5YbCkQtgrR/DwdILpHoyaMCODOvvXvWT9edTkRy+8QwW3seWGeOviqR
7+upW1sWDPr1PCL0wItc7vyKYQS6m460hdUDZzag2WtiVKhRnaT+7sEKyEe+zOvruXHzkFlojA+z
la4f3BtSyoeZwWuo67xNm8UcSIG99UJPecDpjO5NXRIq+I+fQ3eQevw1NFVYmEOg/SHvcd0nrCPR
SabSRxgB3tR30FjiChEB7UzfMiZhG5UQDv1y67gKytmUNWvOPv4If7T/yEJ82oPi6igu5pTAUYwY
219CfcaC2TUER7VF2kEl3hNpKnL/VK0uyWKy5aw8v24jeS6OCC8W0xYmDYIc4Qqzp6k28gNtZl59
41osSptBA11/moYhg7oJIhbq7gMnvSJ6bdNJUuYpYLwcwn6QPM6A9Hpq6JCXwMWw4ui0Ln321edg
CbOdenpJNKTQpRjRpt0xUd3W4P4L84B25upaFvDPj6f2V/EH9AwmyQNPopuva9FzMmc3iVfPJBEd
7jNoG4h4U8Xmf1iG4ZxB73fNo+LlkEgCo4rxEj72YLNgvnwkWzveNYSr37kj/6GWH5J/iY3BEtRO
QeBwevv74Bt+28N0zpV3e8Sn5YHXNPBueEIiXEBJr22C3xbE/FZVrVEO4rhUMbxQ4bvXfu9d5SaY
0OtG5i9mIVU2JxyUoQW+AiUFtde7XOEZAKbXQTI6C5EAGHhACV3sSV4/HDi9nnDKrIyqMsxKJxTU
Ctg6p/v4k2eWuj+/hKFr4GdE2Vh/rYnUDv/7mqq4InloPWWBibVi4Wk5XkEt4MPGDdoSoF7DqFlv
zIHh5Gp5q7iRRscX4Pii9fpmkAaRJcjZiLpAS0So1XFr4PQBiqqRyp00yzqsHSXwtHe8ZaeXcW0L
MpnBergzhePTiAcoQrjT8WDXHYzYTfl7nW2LDVPG43teFUgBTvnNbY2F0XpSZDGvkxblQXpyi4dl
BZSdgKi77UePYf36Dt5T2vyXwNK8da6TgspDDldS40dapjTssPQ0cOXcvGXhrq84bIJnfCZBD5AJ
KZE4Ylc14jUJ5/YT03uQXnPcO8JgHBF/A6E3NaM+dnpWGqZJg14YtqWW9sW0gDDOuElzVbp+XBHa
h+Ydnhmwu/z3uZYTjMgrbvKtEydU5GU6UAJJyVZjvVNDJNkgcjQQLLHLOzq8EaPFG3QihgzKETUT
aLJ7yHrHs5Mx3qlSrwrhNOhlVigq3p8wFci+Y/q6NPjl5FdRQHAyA5pemnQGl4aGbf0r8t09yyp2
n+wDLo+NxxzqcnbI3IKfH+QSI/hDljWumED+DWj2/zw6TgbLy4aAUCP4iV32q06b/RE+9xhiCPbi
mpSsaYf0VzvatJk3xCz4PwYLv43kZTo1hjkwWnsjR+QcsGa+iEiYPf9gm/T5N0vqTxlZ31THPaed
yCiv6lWygte2AHMHzLj+k887HK144/NVo57Am0fn1za2fqW1zjqOZNYx+Wo4Xo18B1SYEkJUxDij
N5PML6wI+gH6pUj+UlzRZk8oWCZInyIqGBEGeNqSgQBKcr9Hz2hhhdfzCPSRQ2/ucuJQrBB8qfFb
ZF8ziZqAGvHicLav7tQDekEJr4yx7k6VwyNQzG3nCP2gDTDF6qV1sAw+r6QZehaoloCLon5bMVfg
kPFLu7byCRkaiATJErFBJ8hhe2OAf1FyH8PhOM2vRwfHpD1p14c4CSS6SltBBp/OVDnlURLJWXs+
wzm/XsgY6vo5i09i/RpT2kjSLH6brtNxe+ytR90V/PxsPkwDjoeys9NRIdkKz3x2kLEElxZgSj6H
5kNYHtwQsQXhYQBs5g6a7To9vs0BmYz3qVIpuQom596hxH2Kn9Rz/xEt6MoCdzvWvwM8YzFgFtmc
9mYbDY8rFEGtvVuEtMOahXFiV3Nmwx3eQo/K+I+zuAwcLlqDg4X1i/8YPRo0wP9Kd+AsAyiHuPkU
WewGLKVBrW0HuqOPwH6Zf8VaLaxRGZOpp61znvBQYXeJ3MV0MP6a0chsMLjCN9FfeOGzsdptWvvo
jXISJiZwVN9UOY0m71ngo5gEnianw3eGG0FhnCsoBYVLPtxjF2cL313hnDDWnOb5DXwgmPkdEoU9
9bX9YFjAdjuIcxIqO4nQM8arDgA+l79qR95gO+hYQGvpVw9gYvAZBDw5m8XPulW8ajHAU0Wjnv0o
vzmCUj3ke501UrBRYbzUhJmFHc/RIDd9MkB5Ry0pAOH/6b4gCXgoRDNJ3TtrCR9NChCmiQmNSCG3
a5ATXi+s+r9Bg5L6d4sxrb0E+sronZSGH0+hk7MtGwmTCcCDBRzqD4jM2S6SjLsfzIqe7FuDTOCF
Akb8JJKNwFhGAAYcRssGKr/5i+4uVX6X1Mj9DEzO2cUQIkXB27cx6ATFj26sA9/xLKZi3YiEY2Js
Ago0m02dV5uIu3yJenzbCn+rKIuDER7r5iMrKi0KUm1ksMQhbo3hu6uFVJDJmNx3gYFiyQzHl7Du
FPy4BE/tAx0+kA5PWUQEgAg0F13+/67k9Wi8qQoJYqkqkuBsXsxDEsCUsYyQYyEqBHaMtw89ZMhi
h17zDGTN6nTBPpBEDb1yefG7MoPa26WDGQQs4A2JNnDP+h4JtgpmQurVUB9ZMF6IaeFSn387m9+Q
c2rxCo9yxe73qxqyghPpgNJaWXBZ0nsa1WXyT3Xv9U4FJgSDy2ZFLnHFOCNVhA8NaS/eoP2bFyma
Q0U20VjYu4I0yFwtt+E9wfW9e/N2E9mc+o1jc9vYJ8+V6oPbeJfZKrByiwbRfQOlcej5etW5q3JQ
q6M574k7n1iSf0+hZ40aWwZBJ0efkBPRr56LwKQOUjErqDrlsHsDcw4zx1TebZcfi0D3fDA9sFiP
ik+cnlxaz988Gh/WTxemGGDxjhh9hLKvctgIDKdY3qLK8Gmp5hf8W7qBFvtTh23z+/lvS4XKdqXy
suEhGA/BFZH4F8yEOKdm4+lawFCze1SXW7BnW4jJomiH4QykhoLX2LLJHwwnu6sY0t90uCkc0qVi
a3ftb1pCPxRsAF8Omotc1I+1y2ovMhJ7/CZ5pzuKf/Y8b3M/8DBAnajfODC7vm3XpIqjOegZca1S
k6ZPd8qjfv/1D6/kXF7wGTZ+SC2AZbuqEBEKyqIhQnlW4jyyCfb0nC/yphG5ei4NmjZROga6fZno
AFyIUCznOauOdivAnhhZJKMoRoQMsx9Lm54gaO5UKlTMj12ccXkeo+syseJ08fKMtUD96Y2TQFLS
N47JW9ofsabvLvBetlFnoh2XFB17/8ggzoDWNqeJ+ztYZsOnfTvsbnsB/1idnXh/bbNuH2VlRki8
i3ZZwRwoaJfWi6DVRmD9NitbPKl1lcGg3Eg5JkmOM5PJ6vOxqug0AWEN6f/tgYZ0Y95iAK1BtWn6
jL9fm2/a5/LgM+wkYVduFA00YIJv8SLwc3jcq52GndrJxs9fj4QETp61lYi/tN8XWFvsD6RxAU6Q
a8hRmpBn6QX2kUziwxbAl+BicXY1U8ac8QAdHS1hzzdU0s5u5nW/H4G8S24XnnoYXmM49GNClD8K
1P2Lwm3ZA0hLrDvtbGl7B15PfNIQ5wcteUXft3pWLzrXVRlU4AjLxMnimAQyIRVx3+rPc+MzD7Gz
o/UeRyRP8essU5ka6m8aijXiBx7B5sF2hL0kZV4swQUrXstLpEg0q159Z6zHJY5B4Vl2kJ331dcK
oT+8p8nLVFofiii5nOo0o5dh1Sv2j6FogdEGz0m2wllgRc/yCcvy3tYzi1tRvXbjqylnWdQ/oBMN
38MEh5xUgKwsAnwWytYUv4gCc3jtUllUEwk4iGt2KtFQ7ps72woQMZz3TDt+dLymrURwE+Cb+by5
P+LiX5fxDjiklAeQEx1eigvwHFXmQ1NP1aAz617sNsEUT+xePVon1NP5vCwlsC0uwh68ByDOwr+y
szGdDnON1wABjXkRn09uubrpRjvfRnJe/f98yGInIuB4c1X1Q7Ibx4xQB1OXiSgcYB/9yQ5C1luk
iLCaRBecNx903PbKJBYPNa53nRZr1Sko27BOKw6MAITby4yU5ZW7WXDuRzY5CnlYGGFgQIO2NKvv
9JeDZ7/M7r0PFa+lSxQqC3Us1M9J/i8QFnO5+RvhwFtplL1650E0IvRzpaNy1yD4vazWeIluDBQs
9yG4GGPfa8snb1sjH61/thKV4xp18njvmedb6S/NnQj3Jhi1gOLNcDG7kpUZQlrVXAL0MBKbLxkE
ueSWgDC/tkIL+gjtKZut07YTtG7dmbYsN4OB/OmrNmH+q5wUbwSpvJk8nvyRbz+/v5pWf43J5bt9
EEhrSZTKBcwNLlEZPBiu/fwYL/Y49yLNCTWt/D5AffvU+Bkekl94gcUnubGio5G+T/OBFpqDCEna
lOcBDZP7OknURHPJEnAIAijDOPsMnmlmgv60h/JE47wl0oTSOHXlIYZQdkrUvJXHTdsbBFNbSFRu
ULPbxGY36un7MlGzJGroDqywIW1wgktxHOy48DaokNne/4X3J01tc+T17tKCoZ0WXfy785q0Fcoe
FN647EON0cdrr8kyiCo9dSi/kccQthnksKqsLFNTthTYISPasmp39Y6I2VAw0AcXetVZu7etOxuZ
StNRB2wm4xbgu3yN2TV9fmz81eEoZhQDmvU/E2KxsoS0SchtzRgOWpNWRtrxgW3xEQVrnrPKI6lC
1wgXudzFiGUOEjmKwdQKTOA56xDym6Keg4xIr3T8PPSQfKQrs6usYfLI5V174zLuxqy6dtNNws/P
VMyMezqFrP7eRYSnsoDGGrpuC1dV1gXctatiGvE8OyPTc3DhYw3qpkJ4MktIknbnkuZauSUi1rQ7
qwZDYIkVGHA3JzF0go2hr6JveL56GtYFtUQlmCXk55BGsZPCiyVjzOi49abj7LckQmdHW8ppUoFO
IDjJHCPAqcI8BDb0oPZW5XKQpiHNiT5UoSx6zExB/mFDQM0D/8CTHpNdd6eCyXDpzRlX31qm6wrA
8/DvED3QmCZ07KVkWX2kXCK44kZRpmQxi6QcCMz7tn2iEDbMJlrPVGMAB/IvCJ35KL/a2+aX1yKE
c0kGwLrDEd7MUTkLqs//FqnQltsvXv7wAC5oi/CO174/JGVSNDbPUnsyQ9f/nrZ4j0ecVjz7dfMV
/hvNaTp4gmaKP2sBXymlQHuabteHEe2nwmaQDg4QnnPRvmEPy0yY7h1ViHMB6uTdw+W0ibmOfNBg
kvSkk/JZkBvmW4FDp9byZmzoz+j4npMSNxsWWv9WvwRe9Sk8zs29RNdDmBGGKrNVKhlMA8cvWhbA
C0S9mxMe4vRD/s50eAqervlOii+mzJ2Tenrvd/zs/+rGdFmFQwbnDqFITBMGtwZuoZV91nnTihvg
0iHtuwbSSkMnarYo+6+nsa/JabfeCD3Z7WDlRCOqk78x6H53scOXA3uXmFRgwFA2NNXOobmJFPB9
+J8iBeFPhGg/3sPWmvw/Y0G+ngGrR3D8gKdAm3Ar1gJSIELEpE3yNLawS1VefuX8PgrrVT7U+N8M
BEapApJ1EOqKJuA8n4xudsyLVCPs88MLFD8Qlin9bmbkBtYlobhiulFcgPhUZDMqOWHNCOLZCK8N
iWu0NQEX3pmpx1YaoDKcR5XohABl+0oiG6ldBzfIuqYFgPzbPDr/KvX5ESe/Iys1SxuOILvmb+Pi
ZkddIAbQuw2aoP1r1U/oX+CvlzakejwEWfLz5WBZXfcywmsDtA7gC26HLdzsqlcy5HFxV4orAiC0
tSpKb6/yXFuoOIJNgAdP+720/XhIZO0MapD+CPuwlXPwtCVCi8Gg6ePeJUA7sscB1FMbXow1h4d2
ViGtAVQFhcoHL7ellTOe1eeAXdExA9vGqJTkYYYQfsxepiH6IhLNPSkTj8hERPnrHnivailjmRP0
F61KmuZi7/HXyf5bkUPHx9xG2RvolmPbnMj52KMQxsC+scX/RhYQyYR0NU2MMSzuZkTY/p3jpNGD
9D7/+xGlEgAAjT4W1N+4+EbPUBRI7HfjG3cQxKm8eSDu9DYDs7eW7/XBpsZ3FmBJPMx76uOx+8P+
WUXo7d5vWFqIN9Ng86SIOCMQjN9jIEh5oMvVHvC2Bgx75jLF8BEbhOoEWBkkHVAgeQ9icOsm+gfT
h9Evp4MNtZpFAc3T0MSsUnzsekh8+KKa4eTXM4rl07825/XUP5zX0OpLdziRoUq4K/cgBBBGkW3v
f8iXX73eHNqfPoQnGgVpLJ3pCLv54b2+MeHcrczHL+YdEqKj5htAcoqY/9l6ibxQDJqC3QCfeWHi
Dwe1MZ+oyBj0IlaB02IX2h0Xdrt5wzEC9pIOdnKSgY6b5JVoAOhY05tbqE4v7cL+8iiGKtPiCxGn
LbcCgGMDpa4Am4b2WLSiH/eM8YHZSNCIlFGpLyBRLIw7qS1TKPIuryJ2Drfrl7YR5SbgBg34kbVQ
pQ/LauVj98cwilyImjFZwRGy37OIuO5vbNEq7QGKQu6K5xud15MFeJp75PJhsFI4MUnNxeVtYJGm
LCKY68HW5lcYqcR76XTHdsNGfSlmIoYVtRR3m9MlaOnfFKkIm1rD8opS9n0gU9zGHH9sdgbreOci
xPGbI9AC/as7c9igOggJsKOgG70U/qEC2lL9ncDLE3kREP3604p9iVVY33dH21rPkvzWjvidgISJ
y/C/ztL+fC/vPB5rynDjFopFetL9dbplEwJ1TP8eoUj96pIpRlaAhplke07y3xZlp1P+5sHvr8Gj
0k77Mgl51KuYK2A/eEeLpThXECbDbjS0YFQ98Vk5nIEc/O0VjSongeIbg4uoVTI/yF8DAwEawjDz
XsI/soQIQPv0LTL0w8tsGA1AiAOKSNuF4C1oxXQd5ctyCkFRjIi4l5B5DslBxKfV4jOshCkZnrhi
GGK9Ot0f0Mn43ah8Quy2gjxhSYh9Z2EeYzVa/ZSgtZqXMdP3F2iEuBcm+tl9xizuZdMLFbNYYVhl
BE3OVaG4hoh3eW51b5ScMjEp/lGSswNNwAJkkll8m0ZC4a3Y9+BZQQ4HpWEmeLvV+IfQj5LTJMZF
nPshd4Do1U0qhielkR9b2DgJZdhAbSNPB9ZlgQr3XiwRXnBZ9FF2vzZ7zqHFTJ+G5WkKN3xwnqJ0
78Rpbpp47CYvNhehx8IvLZLtRO2UdzUk7Nh26WXXsL30AEX0Fc9t8lqpgvw0z2g/gQ3IfDAaNhGn
4OCOzzyyLKazFq0cWOsDrME+mRUyB8KfOWgGuKHGmkKcFMOreQA+WX17dBzcn3S/l49lSr2tuK95
s5p1JBXb9xRNSzFO9VzC6qyOlFBpU0oNMo7ck+mqs9YIZFV7FkFqR2+fc5RjfJnb8P6odN8qsDbi
E+P4B4NqmWkoBDTSQ4RStsT+IBN7OyMpuw5wHAj1S0PCB+7qcW45C0qzrnfkuzrM1TgS2sSRchYY
KpqPQZdek/RxF+5W2oThWEryyElm0VJu6eXrA9fMtlPt9JkEvdwqRGFsFDkE14hkKZ/QbzIDOGqT
VPhkRpdFlZHjzu+6DWdzabw4bHVXl/V2lBs0OLOjElvJTN3ARcREO8pXa7AU46XCdX1c604ie3sb
2NpQIg1BC8Y2XDc25J9sDJU+Qi+3GFvbuYLW0qm3kDjpNsWglWb/J/J/+nL4xR/sJKAbHygDz6au
9pAh1NjvCD1rxPuHUZrAYUBWUJJMCsmYmOgUr0sC7nDym5c802gydJ3F5s+komG0W0IvxCsC0mbF
qmhToUUfZcPepu/76dNH3IaxBThOPSD7B6pXtWLWoxeh3IkRuEj3ikisjmNyIUHLr3d/s2mlukfb
t5rj52G6nUFvGBsOQmr7sUE4Gb95CEhMDjshZiLH7GH+pAvCZ1pSw+uwzmwC6zc4oPPpERHW09SJ
kYuLFiirb+D8MT04LZpXOapVmRIa4WxLre5Mg4GI+cua0QVTJwl8ItdML994a0xS7043TZJqy87N
Eg1RLlxABSXkLbAY/htUtil0yGHruJIaOljpvTf84CoGFHubTOonZoymaqyYOPvBtFyZ7rSOXkul
7uo+hYpuvKzb8rYYSoN6Xc2ZA0PJRGIrnfH45FLzjtEw0pWOvBKsWGFpd6BuLqZezJu7QpdAPXzV
xhNRtHFDBSspgsn5FDq4ws3HaOzERTgaCkMAzDXG0F00Nare6LoA5qxQUy39diOKCimd8juJj1j+
fHs2R2J9chvw7r9Yh7FtT7d5wfk7Mddg96u/fZ9wQcavqYMcGhDzUXrUHeNOpS1j68BaInik0+nX
VF3hrP5WN+akAVT6JUyI6TeMXTVUxWfq8Yal9L5wRqe7xI9gsqSfnYAbYYLkDDRVbrSVTbMv9Eaa
U0c8chAPYs3TQ1On+vbNMdM6yUQI+VA1LLFZn5O7bU6uw/26+oSoPpDcnD1OMKwNBODehpJ7uKIi
81rBrk8Ux3ftaxtGUvfuknMFKxbEaAXwX6EWvbvMM3vScb5jDfRqoTQs0jkObtHg2p2htcamP822
goUhPDcGoX6tuWQUgyqzLvZPG9qd4UJqRr2iyysqS5vpCF5vam3+Vv3SknO2wR7Osbiey/HNRA7J
6iABH5D62+BXjSimmqOaPFB7Wb7/U2/cEqclb3f6oGsNf/qjADVFXOoks2WGXRl0Ru5PrFdWHZ87
gvGEudLA05kly9o/Yxqsy/cJw2/BnGU20tTk2KJ7j2kNUYTGP9MhRV6h0MijF1YKUVC9tbNqwV+C
zrERDODAlSzesL7c90TxiykZdKQ77YnrlBDCRI+CoAG8McSIUazn1FdLSmRCyIHiQi08Cd0HN2e/
UyVu6+TquELJRzXCdX0GuPDeQCUeE6YCInPN0rAtrBTyaMc3BVYtR+e7w5yWBwiUa7uriA912VF0
xcFvE4q8K4dUMn2mbVMB4tt0rjqnLYrLLEbY/Z45y9DFoWTX+RhePMk5mQT/aA7pUrsT9EzpV3Hj
y4/l+yZQlKf4xbmP3O1tfSuFa9eT9AHlIo17ZXBs574x94MXeCC99pbjDponsQn6YX/6+PQZdnHn
XS08eEVajyMd5xD85UzDvqqqNTfYP6k+en7QN+hrHnASnrkGIsVN0/5Obms2BDAAeGaA+LQ0YE0R
tGIXnI6RnFqg0pjYtoS4dJeaBgtbo77L2UePsqIvSkX1bnOIhWBWvuoVUwZY4yb5x4wcUX1aCl7q
bhCtxN5+Qqw78a5b+8J7AqlZLvaGZvmGSGZtNl2n1W4BwrwHhpP5Z/J2bVQXWtaE4knOj0fioQTT
4wYJdiA6sL3zD0iQvsxTP3i6f4S9d0lALf9obZDeaIgiqQCL4U6W4mCSp0tQnMFit6JgjkKIU5+J
fw1vkGY+ryUjMl/2pEOHbMXKHUVSDoI13T1o/0K69aHc6Fsn23HuD04Z3PDBTlqGodPLi7rBw+4E
LeHEtOcud0lxZVFtTMUImZ+Q6rdX9rAyJ+nvga8isTXHcyNFQoXjAFIoa9Y7i+sv57XE/CwPyT54
JqTydaRjYis6SVWKdjpssI8Ic7OmKPRh6ntlXMOQCYw+W7p/eCRTFVCBeQCCSeDn/SHv7oWj8lgB
YqS+JG/9ljhGf4GcghtBdwFVs1BQRLsMDazLNVOmG1lwlNUWkMsMxrvXtWglnHjridpgf8p8ES3U
3E09B0L7cyAytGtnBt3VJf0r9VspV2/Tbjs8G5QDRFEqrkKGKqpDpPmzS/iLlpoO9XvRguhxKzRY
1TPgUWUfbSJttniUkId8fq1FDRjR/vciqLkH+Pv+O2WTMmZKP7rYypkGKT+4qHNV9rtPICyPz0vX
Nq0ikRIe+4e7NhJ0MKqEJTwFxWsgC0FU+YNYM6nMNtWS3wmFIvWzT/3VVbHnpq9IcAGoKNKIcr5U
6I3k7F18+6bUSdF4Wrz5Zyhi6NfLxiFPRcfX3xQis5hgpJhyleb0J3Tn3SbDCEiWmTBbLOKhHwwF
591zgJY+UX1EO/IrmL+OatEdSUJf7tPWSuYwFXMD+/tgbvssHpdsmmwbE7+E+mQlw27YeuZsbCQz
ETAVv/y+ggrHpJK15FKkjZ4av6QGQLcMTbWrjGpOwDWnJzUEMjKpMT12YIiSG2jRKdgojABVRVTz
aZOKOu38MEO6nKtOgDb5qNiUhfhZ/cLRCaIT9ai00Ih9TQreD3RlgegN09ZuDBMtORgZ3OlKpWtT
jlz6a/mLgEp7xpbHw66YfmDqe45JvD1H7NZ3cOGFJF3e/J68dNILcbg2+qeei/ttX4yZv2y3cAdj
j4Sl1okgIDds4Yg6BZ0uu3n7tQdjbt0FWP+QThCTNweir63a7jEL/slGBDT2VwWP3gfDpp/NPQkc
KE+Prbvi+R/wUK6ZxrncTI1Nlt4a+SZcpAHL7H37z1odz4l2+tJBhj9cGkj2q9RLOQ24ANqrW9lh
r3AMQSQrLcWPCplGGgoI3d/ARwI8KaevPZ1NRZYYlAxGtTQQb8zbWH6ibkHF06Im/CEwSz3BlPXu
i1v7G8j8tuPtiI521YN+xbEy1nu5KjHET8/8e8NXpwf13NfL6xm1ew3N0H6vlZ9XK1y09cAe2mfz
klyBo6+pIz69YQkN2HSoMa9mTYefzLdqDw0Pfojtm82m98upqP3qaXT/RifzWkvVVhz6jyKI3L3+
omglBt+xoHD4ZE+7B8RatLVINonXH7tZD/qkS5ShEVOprITPBot7bjZbCjJka8oNuEeMb1FPtf/y
5rRaGi5+kQEsaGLagv4kyEEeehu4fOozgmgxxl+581ddpLvdpdEgXbASkkSfwsdEcm9T+LMF20RR
90Ey6C3c8WhCZanjtUP1nHm8fr0K7tMuWFBdTLtMtJSEc+zjxIVDizJnIx625drRYSA3g0b1n7Rj
R7E7LKhTCRBFadntcLSq7VA7hVzYD41j6Rkuq1u1OmlzZ5C6FMw2QRguhIL0Yy/RM9Fw/9q6O+zx
V+pxnTVgKFKBGLFGKwqg5KwTPSw/qICiLq9GXpYRWY+pSnNVF6pNyGD5ejtNmPwlJjvF9pjdCywJ
cwkQ+YOVEgB04LUeCtz3hI1D5YeAKhHjvvcn+WZLZbk4MIh1ko7dhD2lam5tYXeAHlkZ0ehOL9WL
q3BbGTDWM0GLaUDtzd9I6iwbUPu4cnGsu5TyOQLR3GYdjYkcdBz5NAOBKNg27o2XTs7ynw58Ezqr
X+Xq4IHM5nTPxwSasOmzfspLQ2M1EjbaIzFng130UWqWLFk2QGFUhBt6XAI0MQOmXOlYi74/HN4M
bQIPHKKhYH6dKbPW3Wf7d0ZzLGO5774iI4KZ2aXGN6Fj2vxZOw8TbLgM+UblC2fUSnR2h0NMAyQ0
bobcGmQv06XI4UBFLRS+UpK7DuadYMVnga0jD4T5/reU2e0lhSyOfyjv7pZs30c0n/qcPJy+P5/S
BrBHMxHcmZJTS56y6/NUIZJf7TJ+U6QU86EpplAqmFksdesLtEYLeWm+MkAY6qut4sj96ueYiLwV
655EMuOG0vPHbryKNRwhz9yX2ptgSCGGZvQekRiQnnwqdO5M9P7UTfl9jsw35/kVi7XAYQfbunTU
/OVktO9W2cwz3BjHqO0FZ2KB7MC27g+HlOyb3jujHgpNwO7T675aTo7hEWnp7YZp7WIhewZrdTVX
hW++CnHZO+E37aJy6R8dUIoQ6p7ahH0QOG6U/0+RnqBu+DvCTuYxbv3311Qvn6SFg7qmCx28pJH3
lMF+m4tXtdJZrviwwgMkg/VnlkUPkfGteTtjlGFjcynWayOKgYtEuBpcyY8DOdQ1YK2V5raWKFKz
2e7IqzwZ41LgnjDOO91ZFtCYNXe+VkSRdx+3Fy2g2phBpx40i4n+rR9vV0rBnDXt3PHpXAuIs6zo
Xar+cuwzX/i3+DudnKeABr93T0er4aBCe07AmsDe10h96Xrwm4fy4xySoylEVbI2KK0FY3y+tuwe
BktGlwH2yku9v2gL9ryGO+taZwxqNiL7MF431MpWok45EN+9lhn39kL59vkZADXhiNiCCYkXJYAC
/oRUDR1umnFHirSbpehF0Vc9WujQ9HknO0njsHYu5TivHnHM+dv2DRtvMlDzFnoQmC6rVcQPKPro
0MQ5nYXVqfmlWteIMfSmIo/vlDqhwhbBLy4IsYnPD7aHvwJtiCCb9wXjK86AF4Q+854q0urulWdC
j/1EBoV2cDFygGGY+0O6AP8pFzV+iU4nxbQYqZsNZ7N15RSbPhqKMjlWS1968RD1TF7mPip0316B
qhabaOyjvZavDMidxu/dakPiWziRJjAye3DbFdl9vgYwh/fXSrWR6Ho1aziUN4VILvxqSEV5Q2f8
CoSnUGi9h8pOuyNhpCPN+RECXgwgoXz+gSS5F82lMhLSVtqpqQJ7IpWth4TZwGXx84lpDhu0I+FJ
4uLJ8OrdguuEcanGfZNsXQaiHCyPTZqDC9YeifExfTQuYxYO27+aEFatKchDIkNJf655SO0GM7dF
CcIyIWvwVlGFwJ5X2ML4AM+9B0fz8x4q//Vhn2u1xWo3UxKPMEket+NMX6QiOW07wDYshI3Gw6fC
ejbHN+6sBRbUR434e5SATMOTgWVJBjlS2DXV0bpkOujdulf7TEQJ4DN+hb/W+T7l1GZKFw6DnDNT
YA+O/yC9ieVLXLkhqgNtuRP39Ksmh6OBUthbuiE91rwMNomr7SlvZFR1X68B8l3qdZwlLaRiW86m
AQinFsEDaWKZnO8Qjt09s6mP/ncwinxhTVYZLMbca/2zcMzvShVT9YmQBMFL8qJglucNowSsaU+e
IUaa4UduEMrZV1TSJ2/UO5q2xlsuW+KE9O+WM+vE8yLn9TR0zla6ubJ3zvj8/FeKmm3JgDga/D0L
K4UzFeZiQpSSIUf84rKvCbfVrkGLgRNuTCc6pQT1guaY3KSuCVBspxGEHF7KwI886ygjRkbv/DJT
e4kjiob170qlje+Z2wda+8PX+nXtpD1Ozui1bJxCv0arsYynLtJVSvkvNefk4QpREHSWiMbR83XB
AXpJK+Yy8sedW/1+XOEv+q3NY42GTmq5hwwo8F478MJ22sJXaWdl/xspjcJPqbuC3RrMOMi+3mn2
hsq3M+dcV+invPoZYu420n5YAwceP5WuG4n5iN0jgTLdHK+VlnMWO7gxdO6SSSXWcIGZlhWJgCxP
uYrGr9xUXjmtv7R/C3kK319bP+oGE2mDxetLkhCm9z2kXB0v/KbK3Fmc/4x+E2aztle6g1W7BwHS
HCrvAY8DXQUHyx1zxXHnjcRJaR7VNF31vjyOjtPLDgpo3q/ZdgVEcUSk2lLnxTtaTcNliZRRf694
Ia3eVpbGzFf109r/2vPg4EsBnIhO7asc8TKmSKY56aqWoBlCpUCi15r18UwgolnjMd6xIDLGIn7z
cIW18ObFkMYk2VGNyYeSuGlbmgN1x4vV4D8zkU4kRoDq6ySNJMRwbIoR6HVuAKbQc5VqNWs1OvDo
VXL0EZlROhoGjcJl/LGXHkYyQLS0UdTkz06fBvYYuHkLSt/qjsw+qu0zahGgcLtzgvbb/Q==
`pragma protect end_protected
