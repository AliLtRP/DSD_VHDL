// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:31 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QRhhHkjV5p9nNOVu1cROSEdZSOpRW2XPOgSPIWOK7djFmMUTjR3YZzrr6GRKPM56
Aj6he8sVlbDOizxd/AQbvjz8plLg/vFpIOlNV4vOvQo67azAGNTvEq5Sn89zccdg
dKJOg/xqTNA3ACnJ3P8s+sd75sTRwDnAMne76e/I+Kk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6384)
lpdEqczcZV59xCqhVtkZpFarbTCii2kNbDwBAO57vmKRJAzsEiMywCw90nNhydUu
gSFTcbJ01K9g/zceG5vqCnwKLwudcSmcl7t1vyCUTHZCJgNbcXTcqtv9W16OFtn5
IFX9gSpmbcuP5pDxEuAz7ckA2nYRwXVFFz5k0gHqxIUDDIFDYkzjghJ9kWOKNXXD
/WEIqG+FeVgvqmgJnsluwLKBO8FvbKIOojqcuX4nwoKi46BRvgAa1B+nn2bPdX89
NbBvMl375hGEw1VZqGZvRfU5m2I7Zj0kukN1x5pzgpepnZAsN4UkjJGzPaN5fFjP
oKHGSerfLKlSGVliXVYf2zDUu++5t2BXznYvznQ/zdcvhWm/q7PQYbm8VDysZeJf
dZ3LcAiA507R9K4vBEOqFWiOfYOAWAqDLyNbIKK/HwwTmhoy0ME3xXemefqzWgpr
euB5eCPIUyAoBej8bXO8t0qTSTj2pTLr9sdPxMIgsVZ6OO9cZMFOL4k6F3VWYZ1X
etC9F8zec/cZLGOknNg1clEVIrsgQv4vmPCOH93UWHyEwyE7ISaTPl8LccqtTCIv
35mijnyptsUUjQkkR4EvtaaJlvpi+UCPiDdYIjbJM9yQiiXGbeRde1JNKJa636ib
N4OLfiOuD3y9B87UHxxWO4rkJ/K5rA9miPt2uY9WofN7BQAWC+zsZlT3UTu9F8xy
s+8HHCn2ccwJ8weOlzNTsqR9lccc5P5JwbKVTFJR6NczpuQY6B923zNpiFEqtQFL
foee23yw7MIB86Zjtxj0RNOU44tsedry9BL4luGz/1rXWsCCAY10+SJ3jw5wze2W
WPkg54Qb7Op1cWbDoT9g3i8yB64vE7KkkzKXWbhgIwjBHCpCQZkr2hBep7eMSVIi
4A0Fe+gF7JU0RHh2XnuzCn6OzTm5my+jgLvF3tjGeynWOMGcCk1FYxmqPY3tmYYW
CvsJExiD5KWrmP3kJGhpWQy7DhwM/TPbPWcPTpuRDLunH8i0z36X7DUmBTxCcL5v
+b6CA491wHFukIHyC96HC7LwbbieUEbaZWgvQBYzFtYVYhlM+IhzPA+VkU7gd1pN
Brqcwd5RE01cZzdW2Bpy2nWQKLIMKZSGV3dh18GVnSvmnpPtoVjW3eU6vytJfiV8
VDdyyNcBxkWsybPapx2gNoiIFkzTqbyV3NeraqSKz548s55TKM6Zsu2Kjs0FsKWN
DWG+uZsvOhBFnGqjIS9AzLLuI2wzkJPd4RI/ZzxF0WDdv99Ytj8UCIyXXuuOJm6+
yh37UOuRReUu5HfpmdbFDxADT00pIHH9roPNPBIVno9e5aIJXKVUgM/NhC0PP19r
PHwnMz8WfkLr1LRLZUzsYNQEMJbDj/KG5NbPDNhL9zkHfx9dplgXPXMn2gQcnv4Y
vJrx0K3l2ST+U5Lo7qdvXhDoWQ6m9Xe0DfH+WjQRpE4IJSF5WFZVFOtcNTi+bJy0
3WdAtcH1MHo/Wd0MBy5JTCEY4rkGA1DlFz9PNxmqT6B4b+MAHc35L9WK1qodgoZ4
AdRudU+hd8pRaMgWNZbMcOeOAxKoAZpjLMF/JcdvFMfqzUFEwHKr9TuzaAWq75N+
Q6PRPbdKVjYum2+7MrT3QiTjXy3mjENpJULEgKRwiLPUHpeVPO5KIFWlUi53ERiA
LLcfBsA0HXNfHcYscQCJOgFyMX1mlzln2FEf4J/WSWYCyqoJkhZtrPB8jf1bGKmq
08qJeq1h6eJrWFO3EPut4TcFn/a9Be0osikwbk8Ej6jgkTLAGu60FbMIYi/CQcbY
jVKQ0mSpnCaW5pNQ3916VxBovOxBdMkW0YcEW89oROBbGLbMW34gT5+5yb2l5BU6
jXqWslLE7kD6quxrP0ryO9wz4OG0n7eiP9aW6WbKAqBNhpjiOM8SGxClTz9AxXpl
aojcjEEzSgCE0/ZVoWOaMOfc9se6m5cVrIte+Rv8yACygtkuYMEU1ecIODHV4P24
eHq0HVHA9L5lz0IYZZPNkIow3kmNCT7bA4ZTWomcIwePBYR9PmFQIP2lRN+/YMft
8uk7gw5jASMOlndsy+rgNXa8KlS0UVBZMF32KEe0Oody3uF5bubv6WYKr9QMoAz4
q1BOor9Gkh6poT/EaDYM2/rjS68Oxs+UVXMFfgN3m+03Ki+/76GTwOHDJJAeVrYL
Et42XWpmbon9sdEFRxpUjqdCPA5jzJhUnA8IKq54TRIZKDHpzsUrIIiQ+HUF/Qvq
oZGd/wcqiQHQ4L8KN0z7hLyW7PJWL7TIkIuvUn78BoCPJiQYcvSaY8g4GwUwC65s
TkjQRHWe4l5BOarCmgl/lnEwRNuU5VxMY7zXVWBKwpMGck261baB+r2iQ9PqLfXJ
XK69mVCa3CTW0WDXV7Jl6X+HOgS8zP2PQI5tGg2s7lx3zlXVzJyd7Wzr/aVeEprj
4UszKx2IonYKnG3AXub5CalE7ys+hnspi231mRekkN/0F4DyJuEmGyTiRppZ8k3S
bKHa+p6KtV3r/d3RIwg2vZ4z75rwtgl2WVo5gGJKb+1YfF9nZkhT2OcR/5afgMKc
107lVfEnhpvFp3awR8qEV1MEAERfcUIxgY/28CPOGD/fFRcYgkwiKHn11NtUl6Ta
xLy1zig8bS4XlzHjGCIRFEoinDhxs7YrgwHPLed3MMVlvP++ok+XDsw9MpMqNDJy
l7D+YYSUEZIkRGmTE+oQplQoZ097s6zUqMlx39zpfxSaLwehXU0We6xKsSbFCu/e
DtRtZf2YE1wdEqospfhmGPTPtJhubCm31uYnDxnNIysMUNPqHtT3yAjngABYTtKK
oWC1j3eRFVqhqzor8vXYh7E1pm49ljQmpNL52fyPCIRW6N6vh7Omu3+OKH7X5iA9
4/KGjwFZM7PV3O81ieiVIPUVPmBbd2qBbW39xHuYrH/JRBNO+dpBhypXKdYEnMX+
w9QIOo06tkVsssKcUuSnbyMdETOP6LE6IN6Up5vuK+GAWM4Og1en7iJW+3wNWXIo
k1X1Vbkl1VI28c9gDs+eNXlJIJnfn/xsRb0aC6jFmjJShjHCIblqSukZMUsQsHqx
ZuIgCuwm1y9PvXGMAkkQWJgzOc++xvk4S7SjChFmx/syFzVd5LleiYNbSjFLPSmG
npuqMWKF8pTue5iXJYZHIiZyznDXbrhGw+IoddmpXpmDhHVJeXJO9JylmBuHW/Jd
nUXhSzDeO6OTbun3I8kD+gCCEEWfq5vIF2nvFrGGJ7hd9e9rGC2Qc8+kWSUwgC8J
Kewayck5fVaBhaXmi7DWMaK0eVQ3O9AhVXnbRijZ4jTNvzkTV1BkHYvXhIaBuJp0
kdn98US/MEmNo9JWXaKnu7c3dPY/Q/40n4IM8tIg9mI9O+UtKclYXHncSAzE3xVB
Foe/ChXkx0qT/H76G4wYWVrdp1bh935BBDB4MkG+ZsJ0fJJ5QnY5fvm5yrcs3NTt
s3s45hWQ62pHFr5pfuu3ml1CgvQtwIxF9WTCri8lPeB7/8+YEhzf1qbpNNHnxkEc
mEUcaNUe8XTpOIedIc7zDMHnSpZcdhIECi1HSGggepsaokBbps+G/ZHnzUoe/Hfx
kWZm6vmz4G66XgdxytS2ZFOWXts8KDORZqJ+qSZjZxuEMAJmTCCK6cg1hAzCwYRS
DRtWyghhstLws/eoRQs6NFtD6gy+jU7YmD/h7L1Wrjge1A+22zY6QuD888f4ykUa
jX7JPaCEwlKR9HpoOVdmO3nSLypnafEF5M34yY58S1s/Dz7K9wIbvJkhr6923rAt
mHZyBnQc9ctFRIy3oVaqRSVS8RfiaUsBR+tFj1IywGTYb3nmXEcgsdF/Evhykw/W
zOwpgv4aNQySf8D9SYER4Z/30zH9bz/NtV4GSkHnO9ENtHQAoCpMWnpnX2Ceizw0
/xzSREieMEiezkg25hNiomtjxmVcl91b2tTIJks9eWBJG1k1ngVC1QVCZI0WsLkO
Y8zy+VQZ2Qr0g59pvtlI3sD8X+FM6F1I2lpdDtnWJjUCcoSNS4xChaNXeNyTIBmz
TUMAtLsU2IOsPMwDuvz6TNvH597F6CaKgF4Lq6BeZPAwXCsqWaTog4c4SET0X9iv
Ajvk8Z1P+41TRBSWB5gJvlMJ/khb/kgjS61DrYpPEAVsWRK0T4Iy/RK9YBvyxvbX
5TKt/pGlJqGxhwB/5KKufKMZv8VuxEGpbv7Xpf62QZ/LYmLdoL2Uyw2W64n8t0Ba
SOJR7E61ru6HiHZsL9aQ5OT+jTI+opQn6uv5aANbmGZaxbxIpK1aqo2LjtmiFshU
HZTN5JsSX/+GzWmJa7tXu3+B59aTU2Km6AyOYrDcglSW6w5Y2zmsLuadrglmhBRD
4TkRu49fBs0hNJl7C9wZ4w/Z3hPIJsbF/dOXN/KGVotpFGiNIEMsHlZx6ZxD+6Zc
9WlfVeoc0cuI8ZDxOlIHl0cw5fZP4JMNNd2Vy0siKa1Fnz3CP69Wi+h8e1PvFqrj
MfDG5lOukIEa+8VosfLqYIdXgomBifWhOi18pG8VnYafOofYJ2of/QehmD8xhqAD
QzbaQMNPWX7Qs3SDNMdrY355V1JJ0/RUegz+7lXvyrvTofjxaUEmtmQjeS9nnEuH
wPvgeiJlcxxrtoKLnsxivmQ7cPjaATR6pCwZjveCo+VBhxp3rb8P1Kt5VehrrRUE
YLtr0aT7S/PvXaaTatlQDTkhF9V3PO6qF3Elulibw75tRwoIVkT8eOgo3n4u0VfP
KJGW8uGHJR7/7IwkcZB4WLgL5Aysg7SGT4+oM8VT5JqtsPMBpjHLdzXsefUAE4IP
xyJTlrgk4uqEGGaObhCCE7giJHBc6t4zgMe/vzEFjNqiAVd/pqSHFsAwYl0DmXvC
7ZML+4jTbCjLvoNyq5J2yMP1FGOB//eXI8/y6h7GxHIkkKx8rh+C139oBw+n1Kod
Rv8uZqdyqnLDXvJYSv2xIKFAIGWhA0LBtSrFg0nKCBqoUXwDkBFtb8ZvaxoVdW9m
xu26IvG4hkatlIOpgOetknN8yRKAjUC4oMBJTK9dYxwKF6dNlIDZ28Wqn6HzvJhG
ypr1LMzr9P4hWp/UE4GwKQ4VV0rCvPhg8i1WvfkMlfRwMfOVHNPC4dV0hYTVWtxX
i3HKFRdwfELTUgT6RM/qs2vHBcezKEhdviUEJee5mn8QK5lGFe9B8iGTM6HqMyw7
3gzbp5TYRIbnCB7nny+oH1WoZdYbpxt1RTWswnmLquum3i5tx/JzAgCDYl8nXfbj
2ggEkEqF6nFhxGDq9vtSLhNEZTXHq+la5Yj2jcnTOENE4kB0DqKCXFyzCa+migZT
a7AuCkuqp2RuupEd6nZ9vUYKkQrh2O85ZsKIDlMHOG5FtKJB/GY97l/CV+vo1CBD
ve+Rcm4b30mWrn/AdYQsU3FeJlyH24zNgC6TCnf94n0MPh889wtOipuMW7pkUAkr
9/f8TW5jb+8Uz8NRMCQXFhXTBhBEVbr+wb+V+Wp/QoBOJw8fminLReFRSYJ+yrYE
x/BPD13kv9n5N6hHF6AytYaXSVnuDDG+FwxTSNyP7MUBv49txrfLkfVRNiGZYyUP
bDqobRJFgCaIKwde/UTFI0oDhv2L/VfJYzinBSwaBbp6P9XVtf745KdkBioOWaB3
wu+U18wgFc4DrZ+8OyahV/eeBirf4EaF+P0LgyM1yo3dXtsig2lcPyzaJ5tPP2tA
c4qiBDHvWm9yo/kBatDLMz71gOVJYG0Wv3c1eN6XOaU8hts0PdVR8dw693leIwYc
pq5qk6gI6ywsnrnVgjtHsX50N4EfviCLemErkmx6oZYMUH2jhesTPoG3/gBFIkor
flxO2Kk6+X/byGUV4/tmL0B8Azk8EsXyMGmn/RmlpKMGqwFOCjVReq/ZYeoh7Ftr
GjLQjt1D2GnJ7rgbDpzcjsnfezbDyUpAKi572xzDzZ0pS39h+IUSu0KrkPkPq1Zc
7thBenGEJqiJtx7HuqC8DPXA615v+CrrITmCRGK7U7jk/oEdzQYx/2Pnr0WODsYW
h61G2yd3N36kymjYsGwRvNvbF2duZx8Qoy5FpMgpTDPbgUcUmt2p3EQNtA+BbQsl
X4RRg68unuQPlqWmwV7aV4K3QCE/FsBsCw0nRnOKN+lzkzFziEp0Yaa4CqxmsYmk
wzh26Y8e8RjL+4BXj55jeV8VCcUllfjKxxSGzM+rP9EdK6IB8pPIz2fR2qpszENS
fp3JG4bBRcDMKWqfegUKzk7EF0Bye9WSuJ9ljNdo8Qz2hKvgIR5sqoFGaTCutzUH
vn4NRZoPycNJgGO290g5XMI+FBaAzblCUM+q4azoIDElapSoOoa6mtJKrlpY6VQS
8vT6IS+hUN+zxxyn6VZdRnoQ4rj3PKNCuzkVq0Oh6WA9cFmM7ihgjWU8XlOgK5k8
Popigwta+9O3IRpgGI0tGn/+d/hNVpC8NAIJ+sGVGaFcwTrPqXAc7YOdATIS2vbn
rjeyPxCpcXAy/NVnvVKHiTKbfaSfy9SyTGMlOO9DwYJjmOEohQ12GRgWJIVvP4V7
e1RrQOiMtqA/llOwntYUWEvUAqj9XYhlijKp0sLw8+zHQFK/ETk+rf4CdO/o2lyt
wUn7bskZ/jqZN7Sj47WKAfskIahpNejBPH1J4LTgEEw9X9RHpHgJms2pVn+xEZ2H
30nk8EakNg9QTNRQOtS875vSB5uZwDDjGXGCTVbcsANLrCbCJaI5RoIUzfdOOKlR
I94QN9kQjZSBzrpuNfHIUh7YB19ZHWD6zem9/A5JacjsNhknaVtJshAaIOTdxpp1
siPqpns+BOfPbaWpB9FXVRrqMNVGYYMkbLTKF733Ihc6WgFgOYZNtr8jpZa7QT2c
hxKInsJSosRGEyLre8fTPNvVoMP0WiQxgBdCcBZwaxk29ylle03U7Z7zIoZk3S/O
TlYqWBt2Ekcww/4IbLCtKyaI7T5Dta8MWytCQfy4BBP0ZUsdGW/2j4xgscnzTiqu
a0uyeDRfQeugXfrhSRW+618bbG3kGk8sitjPEOhHMvQUXNB/vqHWMPdIxW1skJ3p
fXtrtB0i/Yp7livFJLqkCXa3VQ3CJJYePeWUHXor72h6reejNUZ1PsP1eKN9Fxwy
/MRQasMx2Co23mZPEV4SWksMKfeq1NknLbPnWBoE3SrP2D/xl9VzDRXo+7V65vQ1
0H1pfoqSHP5hlr/O9Ul6Xo7iRA+boLfwFYNNsTHPiYZZlvjNspp8SF2RcLyyz4JJ
Ok6wixRyjYTTu6zGTXy1G8ATXpDOnueuEDW5OETC1BNGvDR+y7sVdWHPDMRF5He0
RlO47uBsTxmgC1/iBeUb8/kC4aLImqRrf15bSdwFKlchV2N1zAu4MraSbQazYNFO
KlKBNdqD862bnwawY+AqhVKbux3M/ttP+yTlPCArYUPsENeO2n+qJMUWy3gG6jxW
xyTpPPQEicDFFna+qGdFQqGrUNTPN061J7V0y2bUCWHZ5Vd84lvlUZ081ht1iFyN
kWU2M1uQVX1dtObGDVJy0pg+InH2zGvY/++se6c/Duci/Pj7YHTYQGCsO94YlzD8
/WsxB45g0AqrjnHowJm+6l3CO1LdU+VBCy3Pi4V1F21XVvoJ/F2tHQgUP/fbiuSA
1GNsXH06xcphKANdYR5EfoPr0UCWKuY6gn/fmwd2a6tGdBx+seNu0uWvpjJhkCmb
QfQKeZlOb63pPRMHcAv4LANy1L2fwOmMsnNoDEQG3QY7Z8BaMXBYm9nrMymHkPvZ
ii9vwYK0J2hYfDUeSa2FwqsAgsMIUFbBWt8YrY24x11c4NdwjBG5+/t/hylMK3jd
1jOqQjFva4R0/VV75iXTD53H5KxhAX1HmMAvJHjZg5IWN9MARqF/8mdJt/XW5P/F
86t2GNoK7ggvrVb4GzPxLqXx/NjVQt2D1knMVMygCtBQ6l7mu493HTE/F93jOt2w
JLFMrhvYcIaxIiwKKxBK3MQXI7a6/cTzHzB+KjwnR6XrY8fmw3v3rqKYIRAzzOzl
x4vtKsdE9peeb+CPGr1tL3sqN7F/9qS2xkiLuzcVtXC3WiTtsCTxTm5ipnv2OXLk
esaBGgYdV3O2MJFUXmNdM6n19pdF2EdnV+8ZhNHMuCwivptTfn4tQ+i3kISbFklC
Z8ATF9iVHgBlke/3Js2c44xTtAWM/mVpAN4s2P2IJHCiKit3UVVToE5xpWSmOeGV
KnRIHj691tYtsJ3V4/l4Gi+AjPbxvv5OmZLCeXy/2vtMSv4HDAXao6i6fizOy3fB
3M+bFRojpsanUoR23xkWBgtk2gBGhzM6F3NQDwSv85SXbYMN4g2XAEm0S/wHzSdR
lPhIfQnUgB8T30J+Uv1tdb2E6rWe+DwXAG6lNFfzEBTSkWXa50laiEKuLi1WqC8q
9wRrCY9DLdd2ZSrZHTOoXcB8OYp0T2UY4lK/RIp9K2BQ09j3M0YQHP9DLrDtqhGy
Vm3Ke+XjDyElzJuVEXCGy5AwAnBcc3Mx8f1ThEGw+H+7uTWCp9IUeTLoBC8I42hA
`pragma protect end_protected
