// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:18 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Bo8k/NGPX0qZwXnUeXjh6qhTCswVhJ7FWgsivMuYIggVSOmwn6JNBjgiv2S3jIa8
MmzE3kxp6UMV9aMzLxNuoB45Ph1fFm9kHyqb5uSxt/c9K3Y5JSA83jSr9PcQYeUK
GkY4WN0UVEqEzSBFPCNqBiy8y6FaDIB0U4F7hLI83yU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12480)
eAm7tvrf/KWhawJBqULFAv7t2yJJunaneryIr4ccTjW3FqfikQfskE+3iEQWt3NW
DrG5FZhph0lXyzpordh1t9qLRm8+3NVG+reEswAb1FBPhl6+xTzGk5MS1Q7BZS4j
HgBlIHa5WJR5NmAL+HT6fkOuvwe+TG2VHmzAGCx/DFyAgRzSr+6zx7nHjQZQNVj9
AXs7seF5ZVKEJxokdh7dflujoj71av49aLj/LSp7MRWhN7F3di0e4hLA8Mr8UIWK
1ab7onBK7hPCSHw+SU84tLIIyvLTRb+FZsDgWYdPdOjE84qhO26UQZrYBf0yLMJu
5nwve1X2desHV5Zx7+Rh8HAkCbxlD+Bvnyd0Yk4cPykvn4os7pZietKYycKRZIUt
kWvWIB1Dkw0uECYUqEbPPxwSrq2NyI3kJ4/AeepiMQMJSa/+mAFKsiukR+c9M3Dt
0K5VyqF6qh4GcvWUXhpbOCKwmTYrdVleXsBaVHW6IfcJqK+gFw71XVCHURCEjvYw
iA4yo/V30RbbcZZSn0uv0WgGb59E5BNSkUx01SJKGyPlh62Uwbf+GeECPHF9LLBi
IbJ52Nok3NYO/cP4Mz3bP+ZHki0cyo1mYJZlvaMOHwn24gi333ceEgny0noEEdQc
pg1pRHjJDMUnMCd5c2rLT60g/SiSo+NlDuhfSS6VuiAtFgfbZaawqNhYGoRvrO21
V/j4qn/y74tTwwi6FXVfjqGIvFp5aKNhl7xA1nshM4fWE43H+WIsD3TIFXcuyPCp
PY/G/5EMV/qDtlcnecZ+Q21XFaFqB8EzqDIX/WGnd3DdgH0Ap0yWpwfNYyShUjw1
jrV6isK/7qxhnpot7+NewhO25CMb+tciAL4cEZ/wHrW5/B3A3QFWxrsodpToPjJX
YZZyH9FXYq1oB4Zl268chRxK/uxVT9J89Sqq0GIRfzgXHB7ujlihCIwfbo+IOvoM
ey31pT2/fnHArvXGNxcSjnd/4u9nXOtylQGTxe5DmGvDM7yNQc6fGNllkSka98fb
Etzy3zJEuNTmOvZnsjaiJXPOg9CT11kUptf/OzO+BpHud2aR7clVtg/HwzcyT/OV
YPJPNbQ+nTuNaxpc2zIc87+ZgTcxn3kzyD2Yz/DCNK3ptTKlHKaQ6VUI+0hr3mEF
69OQpvJmBQb7IvhWJkFUanrZuUiZ1z+b+Rc0M1/gbI+5/wBwUnI6hdNhsmBNrg75
xzYkqODhGryKzpSS+V/u31boFFvTXf2Vcje/o+lTxqrpXHKUMxg2+a7Mmn0FMDCg
m3huh7r2Z8qVz2L4pDL3LhOakxQmlPqU0lDnutmHAebsD1mHacqEewddmx6KZOrt
EqAC5BxL64FQKeFSPfiSrtwfPIDDAeqypEzqKh0kIun+B8Mmyey53VjeiBK8zz4i
BZPJRlTNwvu+0Lzr1XoNprPbcKO7wMtgAqdO5B/8oOErK59jPwORXdT2cUnx0WXU
9S1ex7PPpTy9/HcKZCHsHtfduZOn7d/mgjAUTKRVTjOL0Ac6eNoabx5QoATLkpVg
2jwav/PZapr/8x8NIRHTq1JILJb9TTiq4JvZSQuySQ3nacbjVtc+VUiHu3d8xzaw
ykmBMOW+KCWXVW+J4WfEmDAucPYnqzS7lBMUuUcnYJE/dtmXWEu6QZL+ZRGl+zw0
aaTUM2XWMR2SgUD7GhvJNc9+PtArbfS8/WXCRETjZNYzSKqoV8OewsBHr+PpQCQ8
+5ZoGrCfVee6zcougLL+kGnjBCtyq/ymlpbW6D0EF04jHvhQJXLcHkQzcBOUwZJs
rOTjM0eCMN4HPXg0WZB7KXGR0V0eMQSyxCfmUBTpSV+ZKPoz9PhBOvM82Ro8XcJH
LIAFjw5+0HkrlcmAe7NVo/MJyi1bYCRNJnXOVrzsr93BhQSjWp1znALI6LfwRjJ0
vG9U9QruiUEZEz7HG6pm5u6rm3Zw3aKdWUCTsnHPE04qoK8wGV1x/GJgiLn24nSI
weKMsqFTRcoWqmUMNuegtaUkSeWqA79V0ZtfgYHJM94NWq/+7PQtN1Z+fSon/uIv
WCQjx4BO7d1gXkezJq/KIlZU717f3lo0GpQpU7bDJztWZaFnt4boWskKcCX5oa85
cIco7PuJ2cDySKF+0O8BXbMIK9L0bHc2Rr9M9tIr3e6rVIJFWYfBKDSIQSwmJcoP
uw8OM2xAwlJWBbhEN+GTZJElxO9ZYI2S0e/g3JBpXeVz94LmLZnr56maUZhO1mJE
1cllBKF1wTkYRz5efWXwLfsOm7MP2/oVOi/DJ7qOimllX2P3g+tcg76bFhewnY/j
DZHHx/rKp3I2W6sF89CHzTILi2GtvyIivoFXM+kqxxO0dvk6SZ2wi9x4zcx89DF+
AkNpjC/+ctTAWBVHjpf5RFzJWk7oHnJdLIA5YP9PAarSFvTnbRGZXHAknfgjBG0+
GT6evfqMb0stRvwpxfVMn2OsZbnj7g7/KzaLBCzggOgDzLXagrj9dT6sfApQ3qTq
E/QPFwbcXKBMEbDBGu5qzmjcqml0po95ZHmWBpRNKG5xLS3v0b982jDvkblCnQyP
PsOQ6apxqCLdma4caZ7rQNVLUzLSFpMOYXk1NUTuw+p4E3MjGKtN3nlo8IBAFhCW
pNBWPUBmswybTsH9gEm2XnCf0FQq/PjKLdPj+JdRzcH2VCuZaQrJvYgQcAgJQB5C
m3CsbvHWQ4ajlA9jnOr2jqQt4B5rVlIcJ2Pfbt99HYoebdTUMdx7Q6T6Qg/1+QWa
2vR0LVQR4eVeT5WD+spJ5qIm3JtKa1uInzqr7isoaeNwODSr2ofnuiODmuZCPEBU
9UbHQq6oiL75jhKRW1bzUdxSk+QVgFz4Y8k37vlP0rU3TTDrAFAfFsyU92F7jQ4C
WrtRt8HIaXkiOutLxkrtSKi6hyPrZvwX6FrrpN/AGv8cOPwYZjs3PgjOEHg3yIDf
XbC2eWdcBpyBnjE1EXzSQbG4QKiRz022R3P8LGKAIvt3Ffxkl2sWuXzeJ4lL1jho
tG0E/VXjts1h2CM0N833ON7sQP1/2wIt6Vzw8JdT/VCIBPom3vkoL1N0dJssxN2i
kW326DgztwclPErKxx/CEQ7AkhR9eL5dMo3uQ3LsWWgH3q3r3FgcMlTHffa/2iTn
bdOfgRrtLiL7VsWqRKcAS63m3I1moL+VAr7vgfv4SUyLk/PJMHheeHt0IFRmViER
uaYj7Soom6an02bLX3CtBs6U/QmCZHJJf/EmxpYfko1AxNvxT628g7vyXVgodld2
U9LzkqKA3czfztxCFfza/Oc+9b8lxG25Ur3Zbmza9+fQ1p0MzSvIBvSUiQyTpx/Z
+wMvFSDODiVlNKMZjlFONTTGy8WiWTt+fQYXDwJ1l26HDBIT7pY5ny4qC70gXeby
Lg4u1cySXc0PzCLzOPI+JIEXwrpqijIVNP6IMVpkZISk1Cvl4ZM7jTioMAYsB2Ji
c1kXwSY2cebqx6YmSyKqYjy4z75m+7/5fNi8Ax9jTS+lslv071o09yQXQW096B64
CfeBeaov7z0xa5rgAxlXcaNWYHjMLOvdlgw6Ze81kmU46ucG7cTjFjmL1YGU+D17
RZxP6J7Yl3BgeSrM++kuzTbupa/w8piN3WXQQu4Z3tH6vffQ77vCWwiU2uNkpBxD
P6wA//CnKv8ReBxyud0rIHb9B97YNRDhfBb6piGD02miXHiq+hxWdG0TW93c5Yzy
pHdta3u/nql9T3XwmPcHNNjgmY2XBgAdWr0pdSnOUqa8yNJnHPShqDqH7RqiHoXc
2h4999g1yP6RqREXMjTjO9gDK44qWSNC93e0mUbgxZrmtFjSV1kT8dvsRsrtBIki
M0ObwXGAY1ax0RrvAlcs9qsdKaG4Z7Cq5aAiv/3HvUt4ZqbXvW3hdt1NeF3N40KR
r1eTTTzCqO47Jv9GA1XoWizCs4I/d7EqufoYonr3L9syudDSJ5/0r9mbE1iD6hG3
Ki4v7MT7lWVzcUK+o7u7xyRVRi393BixA7m9eALol+UkiKMowEV7aYQsGNVGco8a
EeRPheP4La+L9Sb4g8OHpDNiNK+eCxiVs59WgO+iZbYEpNSGDXgQLs+FZo2TATII
8zxgXtEPsEHGeHFtZlTg3HG4fBLTCTYcsj7rZ7khtAl4EWEiDo6I2Cg32Fralz88
+PpWEh4y4AsS0uv6grw7TyGqGq2Av4pQmLnHOgZ7gNPU1VlzHM6FoG4AXaPV6AJT
r1AfmsMhHxr1y8fgj9w8kZOJtSL0s3onlRou6iJQRuEoUpZhpyNou7LpQ62FKRuF
HK0Pco0k4W0mA660KjvmTQrrxr9F1775Ctmz07YJx+okvMTYevNJBS+Hjzfu9CuX
hv5jwsW5wTQWtDcdzt8bgEVH69vS8pKuHWCQf7qfMj+EE2a5M/K8IRSbiHMlZTzU
HYqVecs9JlcfbEYafsEidKUKtEXjamrAVkTzkDYUqsyIxjOrcfRdUHgWj3gnS4f7
RwbtOf1rA4Y5Z9hNa03pgJSEMpE9JUNc5wQbB5LbD/3zoUP/3ga7DncYaQoGPdz2
s5+yC5AS5kWa95fIXBcTgTNKqQMplJ9VVkFGYl2fl0zBtNTorgsop6P7KzvNr3b8
KoFAbPLl1AkoxVNQCi28fPbVN3MrnT5uqGEBpIHrg2jrYpPY+HttFySTEfNnDcCA
Qbtxcyd4b65zv+0MohY9iq9ZI3xt1iX9FXjQzjpoL5cghHWtRqd6t2tcvdT02c/X
1B/gy60e+sp3C2w9gLv1Hj6JydwhIzB9pEFY3rtrxycDiagwlVYyIECcE9y0el1m
JBP6txziAIzsN8FvWs/riBN6SAzwF/2vcWYJWckQxZw9M8iek/pWN093Gw5xuljn
hWeWiDaUPb45NhiQPtOdbS6Xq8QbmzrMLVKyUltsePp6ldN7QPau5z4+mWNOrfGZ
fbXiDn5iTUX1y3rc3vW4ApUy6DR7p3wNNbDYjy4MOEZHW9hiZ6Z7vFv8crWfKgRQ
DMgjeEOXklN+fcdiYUyMfvbkCdi8x48RtM7cdCj2nV58YQrvCbcaZB30zC77j1BX
geE0a0Oz8khgegkJ5e81uxO+3i1Lod7bjwLKKEZSJhpUG4/spVQ2vYYvIrlMczow
XvR2xlkXfysPWrUjvq4R1jP2F9ZaE3Cx7zVhPx9BgJKi+i5i6tzPER6rH41Y524R
VZq5JUmgGlG2ERqLO5ceY8+EApEZbp7AtxOsK8d+Ur45gMFFp9H79pHsEMGT0WaA
3ujMHnjkTDb22B89zLLwVcZjMlS5JhrUVN2UjNTRPVPsUut1/iSJTixV8AwsdWJS
aklbUGRt6LosRjj9vaR6AxcBvu1Dar2W4yE/qMXQLjms9C/XCcuShPDevj1NFE4s
5cseBpKTgrQPJ8CqYxY0hJ4JmK+wXoR4LhSoNamruvOdQtzitowaObf6lu6u6ABc
mTEgbdhnliKRRNVVbfB1dxzwtcpZGmGrrGP6wPIF2B0SDrB4mchjGWtFg4qO1VEy
EL6609LJtZqna5qjWl4Bg/GPefumimfg+gc+xh+CEkb0tjhNj1wQU9yk1u9LIQqJ
b8c6oDnb7U4wAEkCeKnlD/SooHZn565X1v42M/7/ptrcGa3qd7z+hZ1AvhxWbhlg
Lfh0a/DMT/ZUwaEdam1Lk8SKO8JRN3/y6wAWMfFuAaPPSGUv3g3Hk4Ks56An5klk
LcLRQ95UFIU6gE9J2Xxrv04Pr0fSd8C3bbxOgCSH9AG7C8ZCQVIQgXh3Agb+NKwo
wGgJKnfSSsu6YLBgUn/yic+Z1h9fGXc4Vr5YYSyH95L3mUk0daPBk+aQiP0kJ4HG
SM58206Uhj2OhDY0KTUzG1RG0yRoogmj6PTSnt+KZZxJujWL+bGU0fmWYZiQa7wA
jd9iTplyLFLhNuMgaV7PPjq3BNjm3YpUo0NfZ9QGk71qu9ftlHD3Xi0Va9tUX4vw
lQ3XkLDv0UOmNQfiGtpoxgNrLeblBhniQmgO25LaW7MVUF00ngODwxGlUTySJY1Q
afIj88ygdOD/0qxa7N1jfsaqNvqV9z1yIVogIf2NC3hN6IRTfip3/mjxpJHUen5C
FQLDUD17DF17KOKNlce7vJjDErhbgDPWjVE2vIrhn3LgcZp/SPQ7KVQHygXOF0As
cmzMnqAQsrxiFW9o3sjTVOYxC+lRHQ3IA63Gxe2dd48cnTCAGM1R/UPla3QMi3cI
O59bJwmjpMJBcJHeVIR2px2KpeuBU7AE/RxNNuptfIwmyJNAv7zQ1QYsje+d4hnn
jmRiQQi/k4dqbjr1seS6+LXulKmXwg1B0RGXMGzFtX9IMzPxFNx8pa1IKPTBDsA3
HH1xs/SRd5vwXNZ/9xdqkKPqSXFFCfiUkJVyxTRNWGZVdAN0dmRphn0jDIeEcq98
c3WKi9QfJ0znkMY8+fpfR5B8P+hueduxT6tja1bdCKXdzl7bhb5+TBmMloS1hmnZ
vDFApYLSD+UxcOx99Ymt1QVihXNyAcvBHacECkgFbwiPi9yWZlnOSbXzrpSLV78D
dMhrkppw6jqwf1uO9QKzgmYRhDxAl5/TFYS/9Vnmx4+GqodbIco4+weD3yD426oN
5omsz4kJTfjFY1tDfk7YzXSE73IlpXlDBT2nrTGIhJFjVW1tMc8MVRrF8we3BIMb
RNpWFZ/TuCU0meKyQUuVnaSAZQjj+3bhs62L6sPrjqp+RbyHbVX1dA8Lp8/47WLe
MN4x3l5D41AZzsFFpt0uNOXNhGKNvijA+n2NwOFDsr65o+FoM4ALFuUuFQZHmuP1
EoVYp5S/NW1h+psvmjL/lYPQhPEHU8zpZiqbX1JrGzC2WIoSz2VALucB4tGESlkV
bwSQqGu1KDGAnPJV/JQopTmvBQU24cnf0lzao4Np0qrN5QxaQVz/T2rW/M3eGAiF
VgSLuehhQHyjs7+74UMnAP/X7BAAjONsGyd403w/nwzhqtLO482+APflB1knSUyI
mi2a1poG0ePru757Juu5W4diTw2AEZQT5dIqEsKHXEVC1A4VENdZai1DN+hIpMna
4v07F6bUT2daOGt7KzwyAUJC8TDBnx0qmp5/GA+01mbZJHH61QIcqj7OA4viCIcE
c+4EhuZ6HN/k5mjmsYDiDH7Uj8tT1v4qshDOal+V/0heQskKsW6QMftcThgi+ZTj
/PT53TojPHtBHvQ3nejQoYCMjkOKTugs4TEJ8wUBQYfOlcihd74Nv895sJd6ZCGa
96cfcBUIrXgzxUQfwA443tbAG7h0onPrZ0YOq2IVaeA4U+bERDSfs9wNiF1IlAbY
ZQCbskyJDo8bF41amIG/PAe4LHy7pQpHSO4xGkRJYoDDixvFePMiDsfpV6N+KS8r
8fJBKbWIHf1bOnpu9EwnXQSk9er1VEcEpaEvk4O6KQrz06VfNS+xjCs+R3REbZ+M
tCSf8sF0hO8RlOhesg5gHI7n90Kk+cmz8SIqFwskgfVA/sXi+G9SReH2TvICdsLO
GaF5pbDdWxodt/Ocw5xqsrYJEKW0K/oI8gGUzsevRAYDhvciH4PoAX/j67NVbkOx
tc5aBVxVCdia5PBafagiFazhUati+WDSY6wQoBjQFxvSdTPxrfuDxijXFUsbtgit
pinsCUnGkvEqm/dVJ6E2oVBHJDm5ZZ/g8BDALJxrbcVpfmgFnBvrnwY7Bz+jvbna
ZdGHEYn6N1y3Smf3Jd6dV4eTbVnUiZsxZdSLqt9YmkINlIsIyFqxpFCjFVXxhxLI
HhhvbBbbzT4G/ij6Gvqa+nJZVQi7J6068kktz5mF3s6yO5Mgk9eUsx/d9laZG/4W
FO18cn8SCJGMT9htEOXBVscFtyAg64+3yBlTNTYgi5QDpxtLOyAwo7CppdRzIYRM
EuG0oHfBFH8Sd8vxwDAdvUMsrzUPQfEkOqqKxfHno6VMObqMEF2Z1PVQrj1GlHPC
15DmRxienkdMOmNnbqeEY9InD4W1wkHBJxdOv4SEsIMQEloKf8GMg0pJJ8Ts5h98
ehZIKkntIcbizjy6dpTCFrj39HX8/YLOMEo/iK5RHHB+3LRWDBXVFr3ma5SD7ZhU
6FH2DH8AcFx0YskGYCTba+Jb4+szMSJCT9K5I7OWR7hVI631mFV3WSUUxFt/4rNQ
Q1RHnKVj4lCmbIM1/u5V+0qvDNP41RrraJ9mAX3dBQ6QbPu9+qJflVBENw5biaBN
FoOXr0CDf0E8GNC9HqJm5cDmakerQqKKZrDVNSqGzE9b1ki2Bp7uZFZZIOIRsQxT
NxfxiXODbhYjALrl1JXeYk8W3U2rsP6m1tTX9kycCT5ypAF8y2oExf47d5Y+Unz1
m6JK6uNFBFTpVm8t79mSv7GtSgLARh5yoJyOUvektnf4kq0cU2otHAUuUMbVL43c
Az7rg1cDSR+E4m1yqE2gz7730xMv0Mxof9Y6Hf4g7M8QDPBxIkzVi91qWjIgN3ai
xvl27INiwWyeQX302YISuJ5xLN+rEaI7h0RjLm7JJ44WLIsGw/TIXbr5HUpkhRmw
i7Fdj1xFXINB0VAjlbL5yWIsfRgOevg9AnPAh6k/AX1Dtsk+Xg8t/2RHhJEZLQXm
7UwPH+rkm3p7bNHQXSPaWUSJIMgjhjS1eUJzzilj98py7inWrtlcq4JTbT2/MxHN
yD9VkAPXPyXMccgLNR7tXGi+bEH1AC4/AII505PASUmHl0Xjxiq2P8UXQ1Ql0JlV
7k332oP5f5/rNpr7yNzVUdUwDo2YTzuN1TTYMYfQGo6EI0PthNpau8H3ks47BFVi
WoKPWRuj/oG7Nsdce7Jyc9feVZ9g1lXu1P+6D7gzXUUjlVi/ApLaj5bwMfjy3XBf
8bbRhwnblfEsJeaRv2xbGFLPuENTxUokC1RQWlDRG0zXemg910q0uReboUf5G9mK
uxrjJnlLqW+cGp9DyBSC0OhLNs8MEO7gPbhbPtQPS6E0U0ddkb+BKAJMmZmxAsSX
IdWKr4I09eIAVNULue9VLdimQHrNbt4tf4ey4A4H6OT+si8n0Trt9nxrquwBa2bA
AG2Cnp0wMOJkG6PVTaMfbtQ3XTDhmHa/NKp4cc38jGRWeVfS5qFTYbK7pkHrIGWW
Q62H7r/oNmJo1DVZkXhh7R8eZr/NazJsPiDCRwta84GzzHD3dIzGpCBPd3KRs+8L
pnyRCl8vNwCZg/J7NZnh2Ky5+5/6XYT892YX2mqi3qGQdropJag4fBggJcOJMFmD
rOBq3hsmLDbM6RceSGu/7Na6FZSrbRZuXJ2yOrrzBcyPFb7vRpbemXMabxsEjOhd
tVtPd/46TmkgE4VaafYtaRnT7WWM1IX2uc+egsxeJqJE6SSEj7I7dmalEEuB5thE
fIxPi3fgSOK/OqTOkf6wWVqgNwgHxQjA918vzeEf/RPkX3Et0GPgkuW0a6mKHqS1
dJQdHHkIujskvF4W8t90CdMOkNX9jz24hp1wwTpm2HhOaxPezdP2PkVZiZC1bj9b
A1pF4g+tPIN0SQtZ0ml3rBT6z+Hqz3eoItq2+zi2gdkRPTZNQWvg5QogAczH6QGg
T6QI4gWmNoSSvNaylSxxGh4+Dy0E9y6ara/z+1MhIK676Af0hGXfMkTnj41ryetY
kfdHJoHHWBwzSTG0eC/wLTOvc7JI9gTKhdBB48gBF0GT4HfI2cFthNrQ2jvq1141
q9tREXBEFzSGiseHdKGqZ0MHUqMZ4UGNjWtFZ71ZMd+1WPiJc+nlgY85gO+HJsCN
EYcDT+fdgKnD8wIWhc9Th5Elf4/qCfdqS7P3xI3Fup7cHUBy76DRMz1eC6o0iqkJ
k4CGK/09XnMU3EcFFhC84VCS3SkyQnGzqyzaMST57qkjBO9VsgmUkZZfnrexbkQ6
o0UXuZV1xu7zODW63ByK35Gbe4EXEGp9jzxZ0WT7NMSEgkgaadK6TW8R5tVAm2gh
7fjNpD18bv8mjBfGSVhzq0d8LsTElFEdvJ9tU3Wx9PqFxzcYvg/HxtkP625lBp/B
smBHzXUVod7V3OpIMyFpBQGg7zeNh9oTD0Kp3l5mqdb2SDyjOogGX+HVZkejuCPQ
rLk5mCYOEvI9i+HaP1jb5h/WZvnIU0NBY/OiuMSpI5LWPf22oJV+VXz00ahHIAdQ
tH+win1+tHhkZst5f8MA9eDqILfA941J2rS8KmyCysQMg+llS8jTML+lx9xE2qSf
bOa5HsTjUUnO4gAsmRUJunA2uDgv08HD501OGosVwVXkJCMrNBltl/13idqqsjhc
NB1e1PTIbkp6LCBO1gnaOFwbd9NHTnIS3YK0fBdpST/QNkEag729rk5AjlEFI0Z2
aWrnNpdsLHyeK+1vLbfZusROeqHpgaI473479+XE150wZDLaqjhshUyn6TAtR3Oy
8REkW7j37DpzAQCedocY7SitORceyVP1yfNjXPBYyKXH6PmjMozo79xzCFO7o4IL
3m0wMeTNC4Vwo+iEQkDt73gAluAGUTAiVNO/8In0zO/cXgyVeP701jXjUL6kt/il
ugSzb8F8Ff2gCqoEmw42P0rwuRi6ljmuhLzO00zjIlwUnsYCQhraZo7y7PIhsMx+
vUbhe1lL/XSCQq3IT20wHluOeqVLE/Si14Tx1mEzdqt2SO97tQgDEPH43OFwF8d5
S5Q8MT/draOK85zxEo4z3svi7ek9OvEFvXuVIFDJNH9c/3J00RXfhq8N16ARdCiG
bXDFfDijplQf1ZCV+0EBOrLXT6A9b9ucBpabRuCdmUy7cMA08ArEd+pkkOjdBWTK
g5Qw2rzPXg/RqY8r274WLM42inq1bYo7hTjKbd4uEFIkMi4L1XwOynoL2fDoOfij
SQuZay4Y9gR8hmx5SL8ueBs4TOjMhRVWW8+wvgn5pU3XDPyUUDsbSp/dFHexT+ZX
4ovkJzbOlxPCq1cHFMDtuvxG+nwLW3H5F4pQb4493UQ+y84uO3cWSaBT3/b1/t64
1/5VihcpbQ+AxG9CGn3S7zUrmN+PRPF2idrlCtGsA5KPzHloRr5Vm+WzBC5YaxXZ
EdIQOQz1RYA9qaQVDjMHtADxlOMJ4DLMXvYDlLYzYVwdzaT5gpHncedzJhnx6e/c
PN20edtf1xEf+e8kvbDsDfkfvI2qLYHfRwlIJcOtSWhdqeNL/r75+FbSfRR919dZ
8i1SJUzztwI+xPc3j96G0viHVjc27wv1jzSlfcY+19alJig3nUv+SX5d6dBXvatj
fOOHt6wVJDJ1I2miJ3l8d5Vz2qM5DK4hNu7ubW48d/0YER4YYwk5cdVel2bUK0j3
TvxEP2iK6/sUXDRMIW6wOlo0ES3Qba4x2mN8wUh9JL9XfR8JXCK+QxaWXFVAiYfE
/575XspMuReXGuduff0v0tZHKapFsduSsh2GC9/+B+7hXBrEs/z6btuJLM7uajB2
nHwOw8Wdp5V8r5H02EmSrX2bKe44CXlnozsNcSP0zHikvgk4SiYm9igxubxtT0aP
2ZP7tduwqMJT7TLbXPT5akgwh+mHPNJY7Pp/DdH+Xn3ER/2KIVjY5sEth1X+vLqa
3sC2Ug5WCVBblGg/A0QJxltvhDn1EoVvCFHlTajnJkih0s4ls9jfSAmBfBasRoM/
fWNh0/q6tyqxEpxEcoBMLjml3VfkRf1iqcayJifi52CpbEOR5qVToCGyK9BXPS2y
rCNNEhhojPSQyaWvfAAmxngDFW8whnqG3WvwAk9gpsFwRun5Ya1AKN4JlLGT9Hec
wCwZE+PNiTT3OTzGTLqZX+TyIpq4oCWBDSLvPMFNTLjJMLPhazihV3FO+A3CYHAQ
TV8aba+pVLnZpX8iXZHDGae8f5zXyaiTz4yQFUGDDaSof2S2BDuXddjnyaVOLktY
vR8zbb2jHoonDhmur+BF+46XvQSN7upLUQnqad87kkw2gBizpYL8nV0Gh9O4ZCAZ
M8UYJY0LFdOlZC83569BnS0AQOlJ6BfbWEOvNgx6XEA3J9zrbgBOfiP40SofCwmZ
YPP6IiKo2FAu56ryAOZxbqjYwXYgl+Rva4A2wMoq1hC8l0lg0y4I+6OuYuKdPUQj
oG17fXWmUCiiO3uroPM7/nfGMqnbLc8lpKZIHdm5tZmhnRub8b0Z04EJE0mr4Kvb
A7buQ9dYjXtmwkJRMddY6VSi9kfctbYBxVIsSau+QpiwxfeyyzE8gtpX6ntMD+8L
GViwKr2fR4tJdRId868rGod2c4KYBsaYJ6ssBVAPlHJz7AI8lPM1+TDU0lAZardT
WRrPnFq+WJUIwU6kzYr9yJnMD+LWM91pZgJjG8fpz06WC9ZEvRBeMUFftZLI+2Y3
1xfs8XQ4AOmhjvnJnLSzsVPcDo/CufaSulIpHXhTWuQX19HoXcyhPua3wQGR1aeS
1sd8RraZvbSH7uS4qpiVUN5g1Ny+HXie8iXKwmzJzSXGByZ4u6X2TFI1lZ16VYaV
lo9oEx4Nsmgi8UXpqNJWZmEyhjyh83xfy++ibODzXk6rN0R2UrOMp2CsAVjeqSj7
agLsGPSMgKrBJmKgFkXAvQ6jxQnA4z6NSitTd8Td9vULiHevjAwc+LWaeExUNdG6
d9QdqLEXiFn4xLYwnCM2N8tJxvbVu3+48ZGbFwFL4Jd2cLSPfqIUHAB9TyqZfBvg
wdb1ihGmb5MAV7j6mWQ0MOPZQ1Hokjfbu3Qo1Zb7rLuQ5C5K5bFKtd7fWM0APsyq
zdp3CidM9wtmW/OxVbjPqAEZELb8pDqjtfESbL/w2kvdrfxUaqFYCyFITS8/FI73
LoUSjR/USyTDkNvt3MdrwKOZib3cbDQKJ1/2eIWXt8AZ5MIhKg2hFTMM9R8VzZjV
MjkqPbfRB5t+1Ia/LHA13hWXs/o6+WtJXIeA3ydO4tmsshrtrH1t4Gcr38Psu24k
yepRPAd3F8TD53pXdQYx4/rOq8Rn2OrfZpaJmXwS1786NmBzHj2xo36Une2D1bqB
eFuCu9ziuGNBo+YC4D90Pjx4NQ5JAFKogVyvj/eL0IGphv9mXyL7PoK77IP7G61S
CIf9qiRZY+p9d8lqJ/m3JdGAWQgLvfJiLHFxjcBIDEIreclf1zycOnX2lMJtjdJk
guYiMy75k/MKqzuYCi9yqhm4uUiw02ls0ElFVJAHvd0u/eE3jVbzeMM/mSivAJ2r
rzebtIlE1QoC1gWQJeTc74fdaLmhhImPdMwY1X8Yp98jb/dwDYqn/woF6Bfv+9V8
aajLVBrzSUaDKy4yVL5jd0BbyPlpFv1uoKDSSZTJD2rf8EwatVI8sUxdEiweVBQM
weW3imSX5v8JyqYt9aWsbrQFHOJuFcSGV/dTPQ7Dxs2degifC1Y+SHR8uJbH9u/r
V3NlObRzM0jn9Czv3SYQwUC1Uwu1ofsTq7lT/9S4LAIokXPKtpeI17UyefBrWKZ0
DDvm+TuaOfLds+l5olj6AMusFOxw+fzOzPKOW/V+J0XXqK4rzd3OfiZkpFZercN5
43cZKGuY9pk2N3qPLyPJ9XBI18zKKPiyBD9iiHKxAZYDtgdBbxLTyOlBUKVa3W1r
0JucspVDxs3qFN1+GFBX1/YlkyK0o8H1xAJMvDOrq5q5gYijGRoRhgYCNR5WpG0S
/YMog+yOWlfTUe9Yb9M4AAIN+QU+zqU8Yb/dsrh2JYKZG8JjS//jjEsQv7rcTrXR
8iaY2M+ecM6CmfCL1sZaXdrLhdNlB5mF2GilAhyb9tX8d0krEHtAIljmnVSETQWg
1+oSt4XXukNKvNBtoPMR2VITLWRoxrY/EsG7f3+Cmo4uKmAhBwTPtck28LfgLj1r
iIvjJAScHiYrRDq7aYHxUGfyhaoel4miYUaY+7Io4d7nP6VRohQRB2/ZS2xHzfVg
u7K0mHY4kEv1D/MtST+Ziq8Nbe1xJNYK9vciR/3YhWhtDIXwZQldCP0EyYDl31Fo
VAm9drGoTYbzPibhQLFEf5XSa31k6WuXV/Tt275lpSHG9x3PghYULpi3hLE+FALx
M7+bEjU8xCNQICgUQL2KSzNgomz/tsFjmqiC2q0MZFnyZg/HCI08wS9koHMYzvkk
swlD9/o0igYzAkaD7t2jVSG9hFv7+0mV/Yhy05+0/48s5AW9/rgxYUTQ7zPAG+IH
CRZVJWBzDu0NMPpt9zCK0j63MypUod02j4EJs0XrgmVDFpM128dia/rFh5njE0BD
xvJK9MlB1VoQsEjIQac0L6EDbrl/4mSp0X5ycrvsYlJz19bly+f3M/5BrgFQDNxC
rx+vpFAwAiRPV6NsG5b0ae87AF12Pyo12s2UBlM4NH9K92dseForj6zaamIZhHU8
mJoT3ES9cNxgH01MVVOWU2EmT5wFSHgCebXi9ha5BU3mWoDmzPhwHY/pFQFDe87a
3UjeEN/WnAUhyYHxb7Hou+RUhHkWxAPtiBj7WdyQMISKfRVjgEmEoK+cvYW5QkYf
mkTKq+6I3MXzt0P/wOuxnNiZvBMfqrCjLgaiIe1F8qlqS6JA2TzZtvQ3iBivQTKy
5m4W1fFJ72nzXzRXxteTL1pQS6sItx/4hpj+Z2ZN7pv6p258GON4S4mKkk3K/Ovh
Nd/NQyiCFabp1/BgYxFDlJ7i3KolJeImUqaOcfD0dpbDp/UEA7PODYQnp7ZZU0ew
ihycMHOKtTGo8q0QEotXoVeEoObUe3DGFCFnKPnE2nNGyawRRRp4RAAHNmJ9v9cv
bV4caha8phE9p4kOG32b2ha7ZfvsAi5TM9naklb5muT8luRj9Ga0DdoutZA7QGys
CQaRVuv7aSefadUNu9193BboE4NhmPuFSN1MaiExFeNZ3Dm+CUXVUppOxHmLcRoU
kZldx79Ej7hngnOcInkhNXLEMsHO/ZftFmKYwq9L7tSJQLkIPFJaWZ0xAg595/xz
4wUJBXnxfseP9MHvcT/toDw/akKiPJdqa6Gr3Su8BBfTAOwaEITM7ZdqY1Obu8TB
rVBsELWEe7X3/5/KrMlYTjBqqqKI1zf7spQ1TwNKb829Mz60BRPlJdsqXkgCmdDm
15pI0J15SjxhEJKdOu5jKrruy3/QoY1Ck/KkDU1usH5ZZ1vzvJxIak930j3fE82I
Vk4S0Nrgjn2AP9VX1HZQCq9otIt6MXCaLAE8odnQnXEJ3/SHwQuFiqnF0a7wj1gT
n/+Cciamms0pIBJhkTg7P0vNyHa93iinrkIWrQ7N7QvUWNteh9PnqiSyn9SDGWN4
vXXV6TYPhn0tuq9fVbSiJT+G1MNXoX1IIC7HV/kRcjtSIb2nS6azLuJrCzEc59s5
WYwVBEBxYbljgADkQi/i3TL/8o7SGa3bWEtq92ZunmkMLwgtPYne8b/RdebjIaE6
gVUaKMcz7avZzkWtcSc1ceKrOlgmEojJEpYG2DooiXKr6awMBB2vl833xz2uhjQs
KQZWR6HIpz9dbTlrF/S3rX12SJQbMz/fTUSg0E8ndPtpWbBGTUTVXFtEA92U4lBv
5l87s5uUOOQJQVnFl0DdZgX6zT0rbNIahKqO/gWnqpdrtPjEvmprc5vdsaXdl0KZ
lHGHaM12s8wYj4rQCI8rsErODSkZeiRRqFxh8xBm1+Vrm7jNd/g/kVSiaDbF2W9U
KV+hBWaUFFmdeAi9ZqFSd/vP55hQNJ0mpea8y1eY2dIhBpi2G+Kk8ofqZScxfOXJ
QKik6GPZMXsnSYcdAaPCe3fSBTb+uwKeeKuaMfKcARuZSQdlkyDOwvMXXYbuQFxV
irnW66VqoevXnrwAlRlws56zggFCjDmjAJKADjukHXRJEkeAp8/E0xMHEH8LYuqr
o9jdoFPbNvsNb30bau+lWthEwmKLcEZXCMpODdqZKOrvnmdadezay+E31uCjv0+d
jRrE9UcrWae8O0DMldBUyPy3kWNTquOKMpZbZjLrpecJARo6642Jg5080le78drc
BtJxMEiUY/oy4A08dV2jDw/0fpMRsio80narCKb8GVpKphQp7kOYfixpvgo5vC7G
JJSum13VM3ODvXQM5WiOoVWd+ubkPL3oiDmPtIi1HCFzbWIkkkC4Oqmk7UeOcBkw
STHdjqXM5s64p3A7LukuIIXzkj3gdfCvLhzQxT1cq+N3qdXjvv7JKHG5bb9ZbVOf
zcWUM9+LN6mvvSC/F1bk/mud4zwRfWCcjzbKxmiEabIG4IfUpUCJ1hFVsftKoK4u
pXr1GdzUbw4XvbxPB+518ajO451jtR8mRSmNPWeVGYnxtjo/+VQDSw3PQWJF8E9V
96Mcf/ZYm9sF6BTxEDBN/WDzkRYlKFJSP1OBdDLjNsBrz/Q+9CuvYRf7ZtOELtJ3
PhLmZ1TV5+CE1zqXBPNHcc/QXfUEo5RRG5M/BxXR03UNTXJc4FjkyZiLF4DEk5Dx
p7+5WoOXA/oSCFMV5o0TIf7xZuSNT8qSJDFlyRNcF5lkK0rySOPi0pYmpM5rJnLW
++A2kn9/MyDcmrvjZnWU5ui/3hMRslTHJiUh0Ach2Fcd3vdbE/Wq3VRwzHmUrFkP
hwqgSjWnJR7srRLD0CsMnLMiEBX62bTVu7p6vbhSh/gI5bs98GfpsU42c5Z0kx9G
9XBOKh2wHtbofjnH9QyohLrpYE+6+w/iCANZl4BBMcX4ihiU1DcwLvyEpt453BGf
wuSbZdGOaj5lTLS6BzRPpVrIlGW8qK+Ypabh0vmf70Td331lCVyFl5oN4SV7NYZ0
`pragma protect end_protected
