// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Et4kbHcF6iVTS61kcmTd8sNwGZf+/uEkmZhiJJIkCRyNgdMYGm5N36c7Trcf0EFb
2iH6N+g7U2ApPVkUfumTE+mkA4eeXf7XwHZ9HhwnzGxExPVkbeoUjC6b3BFaRvPA
7NzJmVl0uFBLdYgvA+Z8u8ef78upMSpB7Xe1CS47WBE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10736)
pWxwF3us4nsddQlhtBAvGuT3regtLvVffXeFsfPPf+eEpBGDi7yvaDGEw6KDK6Wo
LU8RymZ87HSFmxIM0ZsqXmVdC5k9/Br6l+3I4JVZi52WyHloBDCTc+RRzYFLAuLj
u+ZXC/6DTOjXQ56mvEf4iXIsBzwypF2xYNrlYExD2XAn2qyd3d6rmplwki3y4h5T
Kh0j/qVJUQTLeHAg7Paoox8xpwXspMyWP+Pdx97yCCBibgzVSujQGtmKoqsj5zSc
C0tMTcqqcaXUwNCNztG2E0PfDgwdXS6STUjGTrivxuSy6eZIWmzcDjXz+P7LhLss
/jTNEW1B2tZQMkYEjiQEMipvJNe3VEFAd3RxQY6fofo6o2oQUrKvabGBuN0WlnO/
aVRfXu+IbwpkQvz8YbzBj5oWrbP4Er/b/57ZWh6FjN/E1tIyNlCqCwuB+l/Wqp03
3t8nAXUaXpkoylSYMMudzwtZfgAdMeIhZJ05vq/r18NGyT56gErtMDyOzXvZrThW
diyr6OODOwvzIPEAAfZHLQvc7eCKNJn7WKgGyNex7V/oTobK/7hQ4KBcaCvDUzCn
MwriXy3XWV1an3StOW1mVnQT32Nm8a0GA1eHiM/fjEhI0BN+bXETWJ4WwwNGFTen
xBlzRQYsW2RjQChuu4Ayit/Xz734AmB0e3J70AA3142a3+8iuBTrtKtmIwCAUGWh
lRsEhLXkSfSX8zRCFAMb2NlU7+HyUy7Kx1AjM//JLSWiWIf57iUae4yqmZFc76Mt
AGE8rqFlk3mVbwLjHIS/a7TtVC8egJPzWqT18WuZe+Leot2kAtKosVyq8VVHL6l6
2eFWWqMW8+wr1VrREttaxWVpaJk/BQLa6EmAJ71p8IIA6BFxhNmIXI5kt5k9hbmR
/yDB2uOv1I+joj459D3lBPMQcARaboqRufBzNK6Ah0dWRG6QSv1ldEEmZGI6YWmH
uuRB6RIPOgermssQJ2KyQRivmK8SPoQiisz3M5l4r22oKGbPq/gyHFeqT24ShpfT
sEBucrze4u3m4tuweFnUJ7w0enby9GKyXCivTMdcKl1fyITZVQpoz6eRCKsv/8XY
5kxYfp+fqtZlemCNbe8suH7XHlJVjS8tHKB+Hs+/MoyChbBuwO9NuBWF6S8/oR4d
fTYciJSgjIyRO3aXRTAmCydyJxXGeqIA/UDKcQfVxpsyvIhFVmQVZfnY0WTMDnYp
p3AIsZQdQRZBMhzpnUFQ0LUmwVKE4F9L20xQD4JMTYhbXkxD2k5JCkQeCgG7Eyu9
C2HE50r05coz2IhmQqRdgQvwal9kxH9JuRjNazX4NfUOXKujyhGVGxfj3NJTe6rw
dbO3XtS87woqRsk5j6yDwyp99KYHoxs0C6ZGwKntVPwAWg8d0s588Ka/6ha/ypER
xW0XgfiEn9MvYwU4xxxJV7Byv+tpDClzRxvPeEnWEIbmbA7LA1yGrTiYnRLmlxbB
eeYG9JXOtzKNRBxp/A4gLpMbMNatjf43bAEEXDT/02ESK9thCJdt3AZ//cRIkijn
6rtmiLOKkoKeVJjuSOBSAvgfWF98BfrIQFfJWtQA5P2NmayvSc96E459EfOmAQth
Ip6sdhDm8NvtCa8IDOC/PrjyT4iNkSYbbabQvmW209cFW+VwMKeB8NYquJnlS17z
uoSgpfzZPyFWm4r40ebK/4VO1KaWtYD3k/YnMBqAPJcOvj5ptCpYbks6yKqWAAOg
bSs/oiGBDw958uifKrDF2hYJMJXGdiP9JgTq3KcrlYt1sbAwPLjweAa+pU1chigq
Js1M9frpT0oneHNJIyefDwrQfrstfap7eOEDGa8asgxfCAdsBsOu862n4ZJ0+vHW
8RQNpvPotKxE0RHXOuyc6y6MhREurr0/XuchV529h0fBsBghJc3EqaenFM+Vu1O+
r1FSiv0w6l7xFxu3PDmukDDU1scbekYGxue0o7QWPpa8LniVxhDb/AvitHdF3YQC
P/iHMgrSVrvDqVw3TBnQwCVTIRasRbCOn37c5OhLqQurZjlmY456l66K565IwU3i
VYRxg4CWbCEe/RwaYv+3zQfUXAy2zIPoVMFj+5pkTIyCOZDEU5szqdXFpLA/x0cD
eGEe0ewQFyDJtCehF5vcZr0D9Pvl02hsvvtWOtjjeXORbLzPxn6j0TbOSvuw1PQb
o4tBbzJcqz6EULFPLc3lfRkF4tRwHdCT1rucA5BTpcrXphRlMTxWcCCaV6vITL8s
PJHywq6SFE2TgKiV1PYejvGL7nsr+Ntu18VqdPMI/huD9yqL+0jmihIM+6HAQLLw
hPLvHRuSf2xRWcslHQoBNIiKScw3Y06jf/2kC1A6nuntgHDBim9t8syImE54AKZa
PyEe4ftDb4c38jET9tCtf/iDa5nZMoqhiL38eLN+6IY74FOtZIOIaN+i+FeIVdXW
aQsnei+VbmeT22ULCHol6LNs4cWq0w0UtQn5KqdWLqCHkOB8r2oUdY2DopAcrBUT
2bU8yPdvp2ZsOCb+dzrjEN3OJUesAn0xnblGufyrWEzX1ha5qZ6gh6aEszbEUzYp
B7xcJ9YlV/jdzmRpRxbXCKhtln7VldfJlg3VMT5f/7JB4ORA1aAqrk1WIydDIllL
Fdl4uUEPEJ371c3O5Kcw5F88yC1DgnYg86uTQFkaPnyzbCGjNlmpts1Okj1JO8eA
2fFBguq4ElBob0TUEWImJqvAWBtrEzVzIwvStS0iIYnOZPiTOYCD0niU9IykndCV
n1rvbp0s1fQacezGYCsjKCzfPiB/2t4mV11GEjF4ZCM1mnkcom8mX+HTeeZ/eWiW
TX8mlcB1dgnUq/n25JqGHMaDPXbla22mq7Sgoph3kbZiqVL1+27ZaA7Ftvrp33Ry
vIjd44JRqA4qe0JMLhpn4zp7BPkIGWVXbcjeB8CPalkva6atPwiRiL95V6rEFWcY
JH+48gB7iuWpf4nWjax0kFjAFbuYiIawEmyjKkVnAawLTuiaxV2QOjrmTF7Um59J
UFc0v1KK4QNSUofMYOlPdv+pR7Rv0qc7U/ldatvci8591zmUPRwdUpvDjrxT00yv
9Z8MW7BLUNYqLJJ3HOUYU4PdVvnQilx7omciYiQRt0S771viu5oxA09X3dQeN+TX
4JwYNqkMKNOr+LCMjzBQKb0XpPF6Elo8AGxYQKsXICWjAD8ah4/RI0C0KGnLKdWl
B/szK4IUI4ZuQO3PM6CIvfym09E/RXfKaHyFkxOJTzi1mzAD5um7CgOBOp9Ycvfy
pK6HFsK4u0lIUgnSMgUMlTl84sj337MPrewC4InKOL3gnogWufQBmGammpASTQo0
r54uhSsFLeEPtYZ8z1eRnuOzRAgKkavZOcElXl7YO6tV0YnYe86jDLONyKkQzQmP
/HgpmgObejkjA1hUV6ucLu/HsJkeAeRr9qWB0Hj8CyW43VXZ7d1jcaqywxYLBxRC
3qZGlCoscXJhsKY33sPcLHOzFaI8PprjbKjzKdchEsxwFDw1AmTXGCtq7NTfAYHx
hgqoS3thv96MfcVKv6ADb7+XIxx7/ooW5j1kHj/AkKvsV07DJUp14JCApD4zqryI
Zse7A8mWiZduLmXeLZmaJ6YJBZpkiX84wdzSAj3ZNsDXZKRdpoSMZGitk7uCpCWu
djojd+Ga5i18IUS+7jM0rbVzHcWP5Nard8sGqXcqPONe69xawPhhSmrs/t2hU/fX
umKxRjFBfg/HCDea43j5ZQtXJre/sK9wRNMXnttvlvbQIk+YNp0m2l3pGyOIbHiW
XvApASzthFTAfYn6zxuJS7EH0oyBsbrko1bffbdH+dIDpzsKcQp44mRaeY10klz5
YONOi693CKtx1x9I94tPZq7lQWBHDRrLgbh3CXl/5dnC6sdqWeOjxx0U0eQyqAM/
XTrpYeMSzadexhbh15iVLqRHXK436rErj6Uz0XKGzD7b1CdHODjZ4CBTNXTIBcTs
YWqWEOKDj0I0iloCYXpMuyV7YswTT4n+IbzjcXwU9Yp6FZqYnOPVPFND2o7J93Gk
sBax+SwP/vhLzIGdHm39FUz0aBewAVtjmZOcUqFfdSnW2g+6hBOb+y8vvFMy5oOp
DZj+1x6CeFabNrm1etJ+uu7mKkEXqgSef/ukKHo9QjzlF2utYojfvuTUxer4Mktv
bvTY1SYvZN5cMgfpIqnKY7PW6D6IN5UOU/GSwcCzgSbsKsWci6t12WkCpS5IT1EN
DG9DbcsiJuKeqF5V3We0AB348NWP7Lunxu1bu/b/nbCVDgRV+9jMTUxXS7ukqhEd
uwTB+qirxsL/fy+pcQERxunRJ2jqCqf4kdRNxDYs3l7AtJxgjm5sdI6/s5lwv9YD
sfd9ghzDwNqad3Jm2T+VSIVZ6AQupVTuG1XWwBYZIpY3BVT7nSuaOqwAEBZko4d7
qUy9s65FTtgqXQv4J6UJcX3DCtA8o0W6lHITicqWDbic5QhipPeaMj8WfmC56nzf
BRIh/RWbH5MRKeWuTN1WsdfAfNnsoNMVQMo/Rz2yuL8GrJQn+rUwExnIujHum298
YXPmlsA2J9kcqOomTopTyCam0N+Zrkp1hJH6Z4EILsCMg8IVED2pSJ/hDIJES/l9
Zba5BvUYWgKo6VPVldVHNeqxEmGtpcPMF0sxDpJBQEaBvwb010a9qcSkFSlOinlZ
CiZ5yFw+5yD8c7BKPiEjCEvNQZgX9ybRSNJ712OhmCcMLvJqmpjvAM7uCMBcBdMP
U1PUFoK0bQoqb0ETgdD22NvUHaKmyABY7F+wNrpmy1CThKLjAdJCkij+x1xsIKBm
RP55fzpVoiH0Cs1psbRiXn3KEEa8jY0uI3C28IVMBFcXvmH/K3cMSonhmp8zDLO4
7hsQDymcHB1GBs0kB8JK//BtBpqZhbn4wSIzsPNUTF7YKkats8ek+7y4ckIfaEMb
9SfAC00qOeejx6zbVLhSgZ6xbO6HA8QzaFxRvXju+MmAPAQK2Cm4Hz7YYmOemNlC
a4SiTlC80dykzaQRD97eW/7v7NwVpVAvQtw8YJjTCnwnBps2dKUmAB0HdqkmS7CM
fmUHt1/LVX42NJliihqJWE1DnN5HR9uLkanKX4qcg/pdYB47irynn6NDLdyOHXoF
oJFiksdHaq2EY5Q1H+w4mAPBoRL3Fb7BdmTYbfzAwavmEwm1NAPcsNs3zbjh0moW
HA7KKQ5k55HDfLpNkjncZ33DD2fdLcjiPQ43K6mEmeza8msrkUd9rCgsqEorOteL
hEwEzbrl/jJJZ/0nqPUj4mO8w4WYnKKQxzPNm61NNw/yHiYePHqS9vLBzOJ2kvY7
/lNuPpQaXdKAZMQaLjlzbNvfH+anpzowiLvW5SW22j7921xWPDWpgVIi/eqi8xAe
p5KGy5bmEMuBeYQyvhafLS1+QV0fc0uAtYmFE8WBLH+AxksjWUKweK1K2SdLY3qy
07HA4OAwWarXCxlwSxa2POkc0FR5kjcrhxj0zu9FEI5JC0sU2Qm/u1cmi5PFI2+r
hlY0ZdAqTmddWBq3rPMe98jPA8LCaJ+u9BgVGtX4bwD/FjCp8LePdBFQPA9MeDyv
pACgnqowOevGHAD6HY1XK9eWC2/lvbVC99WAwQCeCgbcjVKtxOnUVMhAidG430Mt
/IhqlKqNaW0K58nEK3IEPV7BdV0oEbQZk4uNmTgJx79TeyRjHFJK9KTRQ9TY9mDB
2q2qkX5JT8MG+0iRYNjKBthJViSlmpdVlV1KpeY134q2emi1njiYICA8lj0V98+h
kryfXEHliqUYa/mB+rP0kjT+F+b/tauSrl2IzMskMVgTbcErmSr+K9BSj2KCvzrf
RTQvG5kOUUrRmACtetZhWTTIU99VrK5nVc77+1wiqgUKuvwv4WwcZHJAqJ/N/e3J
afljgv8eqoaKDKsFgdxQDv7611YrhZi0ZnaCD+311Gs5GvEHSNZNyAa3sDNYE35n
7TOEZ5bD43L45Zo2A2sq7DkYRSzpi5A8kMOLGabs3vcgcxVmVs4VGSIz9e5FBZbO
jYQC2qat1N39FbbO/qPdM2l3SsXAIol5PIMQ7Rbuv+JUZUKwKe196h5GrwKIJJv8
ltOiW0BqUiHALaBX0r8m/fcIwniDaFSOMrkB2oDCxvtVVV9t/bPC4oCwyyrp7MXE
VXxG/tg8QwIk/oMMcAlBjC65LknVb7ooWmK88XCjIzm7ZjN6JTqFjYZQTNEQYUjz
0Yx285SJ7vgXCCGUbk/EZh3xpk6Ycf4i4qqE5CLbWvraOb2tjENZXlQbb+wRMWSE
qxxtSw9NuSFgbKtrIHaG9XJEozKFoloUoeUAY7c+5NSd7ZjD1jjB4k7HUM0wFPL0
9o7ttBPW64lTuvEEMFGPJFs9Oem8Cb3j8FHTHhBYUOsgkHvxZgBG4ylgEfei5wjJ
2go4AvL82jMHVP0T0t86C53Ix5bRsc2P/9x5fXLLd/6mUuiWLUA7fgG5smDAQXiz
OuhWlGPZ4zfe9o5zVWGlShFD5laiZbqi82nKKwxRHILap5HkUZkOX715OudUiplM
drdWicIEP66My9uUH3KQeRmlcmIGCGR+JlpQTgrJCKtnTayppg6xmyIkac6Mxy1z
FKBiGcvErgwA0v3YigO6bmfbhqd2HdUEuG//p+Kd3+7dTepzZLSx9R0aXKlqRSkA
WdTeOGTLDWh9FULJ9RUKXwJSuxI7KwHFnBdYip4MRC0hm4oi3ZiQcoEbCQbkhyAo
5AMMS0ekCq0gFjvcO07dyTvho3vsMOxlP2R5sSYgjJFNd/E/nK33wcHzm5lruEGd
oyRaK6lDKzoGHw50aE1KhAz4l+ykw7aqiEXI4Fx4p3HSd71toG1f0+ZFkFEC78rB
+beyo3P4VjQiu++hYBr2MH0O0ucDlMt9FDZ/T5T6qZP4Fh8PVjNjPWomD0gpBupW
N2O3MdgByW00TNzo5J9A5LZfDE2H7R+Pm1zVhsh8qp9/9TrYyUNy6bqZHUbZ31O9
Xv6LmH58PQQLbyJ81UNsmaXPqtxXFdqDigGIgerC4xzSd1I63a0ubSLJQynahdjb
RqWronDPKDr2R+Af5aaINDMQtWO+5kbypk5VjSOJDNVDsR78eIYyuEP54KzOfpDq
L+7iiS5DmYFEdSdORdLPSvMPQzeAeSVXnG4NJM7qqOtdMdCll5aHw6pg77SZ5B+e
vbxovnqBNZt7so6EzJyRpLnEWNfQG9FvOXCa96IAJrUxw5RZsrVCcuLl0ZhNCFvL
MjLGxOJr2ZNgyl3UtbaQd9VrC+tMMW7mVkvRvHGyZDM+GXD2HuSjfyTeqkaMvqRL
qfmjzSZCUKby53gwGsznbYmRh6cCQEZk+51QHecT1Yffc+wVk9FTMAAVCBYpXq/c
nTk8fOy0ktUvuOcuuei27keSD2hNNqGFqnd+tpJp6HyQhJOEnsti1mqMWQT4LqS/
WmDBFMiBBWRfELk8WGB7iOeCkyzacABIDIPiDRmmfKPH/xv0dx13meWZj+xq54qF
S5ta9eex4UVE3ZLz9ohSraOxMGAtA3EMbTjv6G+3LAyv3BlJC7xzMzUyvFWLzqH9
YYa8x+slJcjRarM6IRgEFJsU7/3VvGC4VsKRZsKKfinLMXJj0V8SNmOkzDWjm/HK
GKCeBOMdr47uocysQVFBYnHCH7j3W16mpqFJNxNgx7ZhjO9Ia4ixhovOq366ivN/
ANDOI7uqPefKUBN8RSiHJXRte8UylimBp6ib0oU3EQ5VpbhYUIlNIwXpiyO992Il
lJd4UUGe0uFLbieI5H028RF7O7xRSW12BkICZGwXUMdhuAiWWmt2WzDHs+27XTgn
5YChPFt+4b/il4CIPMWevxH/q0O/1XDeGiD66Wmt1rcOfqVeePtWHC1PuMwVqsIv
zqF5SsWij9aEDUwxkOlQSunzwOr+zHoYITih5DbRy1F5s95CeACTwV3Ta5E91zvu
8leRLN1mtHUEC9Y+mMjZMnT6eMz8bsu2mc8uB3r5VgqPSACXlnHkJ99/Mo+kURWq
evtsO+QI7LZosZhQJB2g5yLJ8SK4lrogcTt3oSlAuZJKUfA/aqEA6uaD/GtRDk48
OdV26EDEUwnBaWLAKVSZlYNfTx+gcMSiaRCuTEoLXXZ43e9RUFhyafrcTwLiN83c
UQwcn4bKGhDzn6jQ4+zbsyiemayYDsswvptX8ZJhx/olRKLuk83yILYwea+3/5q/
sNIlHQAs+1+UhAgxc6p0yQmn5FhN25edsKZLNWdtXH98IYiNkbIcysPEYQz4PSwe
6ZHo1cfomauR9ryZyuVvyCDU80iyoFWCrAZKTKXAA3HehCaXEb+mSVFmTmItRc4p
+a/wuInomlDRRqbCiljIZkQsGUb6KkGLGjfhMrc92XJFdqmBwxPsdhat5uP6t7Op
NdnFP5bJQV55IBAFejPi48H9Ye4VC3cLnFDc74bV9uEqy8e1taZa9liyh2G2tTuE
HgfpQsvdVDh/24S4f5FcNHLLf7jsgiJ9FzOoFWtc0h7B76QoJOtTbCiMv05h8QBj
qudXucRz0pyHJzG6V+FyNB4vNkM7oXn6huI2uD/5AAGJWGDgWE45/RHpi9f325ci
n4okGiDxM1JqHygyKEobUWjA2CO7In1Fh4SISO4mynmvY9/dD5d/F5sVpUmKBb/S
YxqIERmkOIdQ5oYmAARcdFIukx0CFx34pO54fCkqpA1cKnh47Z1BOhNdJx8iaOgD
OfUyveaM9PnR04XVqdGqsDaAx3H/oxWk7f7YPvZguPcbm829BOKutBGJ7CguKqQb
9b3L2Kn3kxNw2bmYok7ih/72SypWhn6oiieaZJ92Zob8ZNLGQn8rdic6E7OKv6nx
eZ6iBdA4QveoPZcur7QCMtw3yXyGx7czLTAGrO2w82YzjR4hO4zFw/y7l6eYyCk7
f12c95ipNJI3N0WCPOsa9KSTX9QdQQe1Vt+m+JbjlZL/iO6n61FtyYtTyO+z4Ija
1PP5akAk2sukfS5yXiJZCAn89JbbDzpAMGNkhikX3x73+MGf5uJacv15nzdxSOW4
uYmQHX2rbVAdQ0YH82xk1+IDEDtr6/hSr9h2QbzQoKi34988VRRKzysV1h4MnN0a
zeb5xB8CNhxSc1foXhY8Vbm0V+HCcmWzp+4rcD938z0GPgFIMFb5knjfR3shiz4S
jWDlGnLALXINA61qQ8x7fyHkd/hffK8aPJFWLSeA5IOV2mX1iCy3Bpr7O8BQfrqE
wJ0a2OhJp64JmV/gpN25mfHaEFcToEHRhfj7RbDwGHt3QNTYOXj3/85ACDmZRrzM
qWB2OvOyzf3oDkk6NWTz51I39hGGVDQQnw8+SLPGQRJhWWm+rpx0wkueAl+Gwn06
C0eURCxZ6uVEGAv4Ly5I3kn2IpwE8iuEjC0MryDHj2ay/beaM2CkDLxNwNkRqY6X
riC06vEeIqht6r43L9K/bvqitsazKWSOgavb4cLHitCm0BCI+M+HueE8RTdYfhgK
b2fXzuJ6y0SNBiEdvY8pfuq1RdwnumOoVGsiICG+kx2ja1/qxO92/OYI754xLduj
DEu/vjmeLDc2w/ke6J8Sxa+9cKqMaQRhWfpa114q0vBwftLTcGBr+rueIedSUox3
jRadIsNKL3tdNrxq12oJd6mUKHZkwr5dT/yj5TnbcMl0NlROkySxe4Vmfa7PrIqF
c8csDrBYlVP/a5IUB0D8sFmhq0y2scmVUI2hY+4yxtfVGFPemJPsGCeynAjoXFjP
lze5HjY/umAzArj4TYfTCyjo9tUauVf7+yPJs1gr1bUEH4Q57zSzqG1xxCCbhYOO
tYikwFlqAzvFJmHkjmxDcnNQk5yUkCNRK3WwzYyy/W1mhAWmcPb07XcjIX3jTnJY
InEDomHWiuVAql5NeZt0KWE1RmKM5MyB5fVhavpGbSFvNoKprlJhMYxE35QbXANR
3VDF2ik9UIekQnoWYd0FZuQbtWuKV5HT9FLc3kQX+s29pWatIfujKEpOTZl8jMMx
L0rACzV2mBU27H1NzSpA0QsJmUft/WA71dI8o/2N/XuJSEevOeKrI2vIHWJGwdHT
ZsbubxJts/ahrZcEReZGKgkuwy2vgSek1e9b1AgpcMFtGzVjdtK0VXAKytWAHTPT
NAZMO7QuFrwolunGefxJAxhKKvMQWBSo6Avot7W8/cykmShBGJZ3RSqSG0rJBblM
CSx1bvBICnw1n1rSjpnqjWC1va0Dlyb12i+NZ0g4cdPg/yw3F4e/hjKuhS8yzDXd
xiXzuCkI0ob4RhSWeQ+x1ftPoEI61XS8Qqfc9cWb9niHPepiJZFRo78Y9L67yocJ
+rUsdiV3KJSqMSh9AbjLvs5MymP4/kUpZ1MfVrt1fmYU95ShRPLlRpzUZmmo5fJV
spXUwxTBNeEEZQmIbK5kLeIHiAxW/26B8SskheO8yLpFgiyP6UjhTvMM8vxRYNaR
pvsjrvHesMoq76MsBTxqNBH0iu5c6WcSmRKIe1ZPfX1t+DB5FJZr7FqyZm0WsFAI
3M2Eu+EfvQuzRfazu308XV5XTYpZv+y435VJPbTCk4V3vd29XL6HK5asynRQTPZF
89OS/elo/GJaJanr5n4NtlJHo4V7PR2R8CdbJTLtA4M30xdM45zPaX9+Sja33FFV
IiPV1qTFxzqfKOxl5vixEOKmWiJnd3V9URFO4vYVWfF7vYS8fEGH1VOow+JMQx0X
ownFpjE+TE2Rzql5dn2Ai5d4RgGBdHDbMAlRMhYPg0lr34Pu1wnS6ynSkox9GUMl
lN6XsIFanBxL60LIyuEasLeodYYyXtsn2iXobyOHh91zfA0eCGWKkA4hYgjhtulb
qBEBuoSWvDmyG1DYQakkgjypX/zgqXHwjoFX2DnYyjG0iBgRChDuLV1AtEjVZNke
RhiuoDuvTvQX0adS2Ru8S0wyhQxauzXauCEelnLBdv4fGYzi3neuHOL9wpISwxIG
kON/frH+PqGS4O9S0os3peVPLtUQbTjZXxND1QBbpVxnFHBqPIV7HLN7hRG7qoCk
BeBb8qwZYIG+QPJmtvp8RoNgk6BE4ddjYpM9Vqlz39gklRoV95rjVcJNXRrxSs1Z
0Q2v7KHVgJEmsoQfSU9PizWTb4xJbQ/NXRaWw1Olmmp53oalrBn0gEHuZ7TkTPwb
P9bA4zQggPa8fBX9w0YY3ioAiv5KkW91fBCc9RWXulei+Y2GlggL0kjwkRCu4aXs
SFwp2ACG178HBwO6p+e3VR4+Fub2BAyR58zt6LTf+TU8OrvqnnjgjqC+fbnvdmOp
Cv3llAh1w45Ndd5QfQn/GaCKaSFdd0N0hErzlzaBU3tBeC5GBYYG9iyLP/QxKHSb
KNwWTZaUljH+/XKFuYxGdrs4ziF7EmDvRy6wqh5kkqzZmKoEeyxB98qUcQUp/Vnr
8mbrMPxufKGQib4kZ1jt2jkO+xJGoid1qU8X/gS1h+565Vooa7wwCO0D3bSsH96v
0uWDovz61BX+w1ruhsh4+CjKZQpYw+4O9MamDol8gBvbSpoJBQmbrr53X/q5imIA
hfewBkHPhoMM9u6BhZCAT2FJU4Cvhy9Veh8zXURE/BJz3P0nZzFB/oBMg2RZcKFe
aEYLj4OfAT9Aym+mfTp5U/aUbWrRd+63KgWZsBez9wmbB2OiwaVuZgheMBtl6mgY
x/wSOzqXHx34ktc6RNKi/qsT1Zd9gfWjln+VPFkZ05hHUg5MairO8gc1pSMm/xqM
Z3CDBKUI9hyuP9KKxoGcwtz181gxavuNchjFnh/sYyIf/1Agyx0qjSNqVu19EzK7
6QPU6xPcSiUUTqEv4HQI3t2m11cT5l5X1jS0Uvx+wfk5XVVrRwLjwozFozakr3dR
jPKvxUtMqv3egW29x9ciFXZ2HcZlXsOkYpLYMdVt8mPyx75EFwkV0R3AEUwbBwR2
a0psydTyBsrwEaEiEM+9eVrplp5DhNAW7wrAWAS3K6WZ2nDEG1YKMsft+oM/4aQL
Q7L9r3Z3nhgwBDWEfCIpexR4rtVPorcDeVMU1Q5xO0jLC4bDoVBCnfogWzNm8d7E
Viza/338kwJYZTjnwyWq+iHuKWkRKFFi+MHoX4mzB7OHsxdMnC3odbMMOExTQdFC
yJtcfBlBobY3S8EPhUux04p2uD5KcJIujby99SiGE8BM2wdk6t0WNbYUJMEHeJq4
uq8izbzADEdTWO21E0VCJNuA1n1cRfdDcLt8jaSDiONhrC7btsVJuxNF63mK5rPw
d19Vo8c/cmO7LjJ/SFZYLJ6KqXOI3igkjDFXarfZf/b4o9WAueXcZ3/MXK+qhGsa
wdwYsGKUfOEa/aCkAdy1zXv2VlEJIkOeTS6Gked+Fyw+k1v5NwYxj6NVcPPdpHUL
yg+OMNb+G1JBcW/leETWpFEHO7RKCbYegngMfxr8L0Ex/gME9GeoPcRACVvFSkpe
Su9Yg9wy1dxXBROlsWsY2JIWTH6IQeFZoJtKMURMYTU2tgQbdN2V44Qq5q81AaDY
SRhmBthRRLW0xxF1sXmyUAO9OPfwEJCExCwNiJ9wrQJS8Y68wtOQIAwUc5ZCsRfI
z8rNyKH9fmXzDqUzImCFI3AoBkAvSqoWmJ/diJuyzsTd3s9GeTye1unKv1ruoq7I
oLqa6IdTeK+5N8VHTkmC7Gw5XiRIJHkQDFiSIHXtmx73CurSlJFbwzGVXcjcikDB
jNuW3b13BHloGwMebFTjITadLgW9iz519nE90wWdT3Kojma74t60wwsAvhKdst+N
F9aaassiiRkJoDg4KmCS6OYdt0+A8OmlBRvpy/aZo3YPQ0CeBzPuC4xWnoEnPi6d
elN8N6H910gpir1MdbMEOlT8DIZrS664A9OCjXUGNXMWejzpOK+OK+91Gpbi/53K
eGDo0j4SLeFSHX2I/iZtjii3Bk3DhCz3+g1MbJgR4JLrgnOkEONbHOs0YGMQryGT
dVVVTZFZsN4uAqDKbfySgdojXoyIBdISGtRCvaeMFPHll67Re59WQB/6yaCnED4L
15eTWxHSp9pPZcpJ9VeUGmHVfIzgwIbwP+zJzu2yEOR2C/NtbW6PwNUsnC+9BF00
EfUx2sjTA/DCHhhTigEFSWeGnreQniclEnNqOjCMS5wxQfSf3BHfknd4GWcz6uNw
HY78Ch/aSGh92Dg+mIxZ9YDYtmeeCbeDf3CZJ9K5bg7PeQsQhEblqQrEaYAoCTaH
LLVdOUcJa91osdAxMG6IKCi4icTyYtEY6AmaTt7LFWpH+crQUkDTsw4slMJDB5in
oPi2lf+K+I7L90UQyc9vE0o6yv3uFBWUnVL/SeQ+NFQJstTMWC1zaAr10K5f9y05
H9PWrSDD/ZRHJagO8GfwkZmEr7F9iu9QcZA0TLizczTZqEQr7yKqM/jQF5uMGb9A
+V7kayLS6i9juEsNI3YbgCJxZ7RBQACNEdsPFAMu4OqIKAVuwwgBKFZsybmpTCjO
O3YOX8Dz30dJGC7LFx12TKLNAWlppuy/9ejRGv+rd1tWZ3BUAefozaZ6qIv80X5v
vEaSp+7P4ntgc3+ZgTH9wAzbVq6trmpTPnDr2JQRJ70SFIpF+Rq59j9TdxRfVZHN
xROYd/B5hRkBUd9rjEb102f3Kc2K8FyTMnvhlgH86YEpVWYkwGGgbx8ieUHCJduD
zB31pKEuZbIWbua/ShlBFoi1xQfxpgXr2WL5Hf3zfL+RwD4KD/Pjk1fj39fMubqW
KA++rNYFdIfsw7+xYFoWNwPHO4ume3kg5oifGlN6Byq8DL0GmSB16BopKgo5UEU+
VQbRUhsL/QoS13yjVR1ZKvAqFhbELFsP8F4HF0kv6RKM71GbAXyr3S+vcsGOjQpx
/qeKwcRadpdTj1A7z+gQJcSqdNUxZnoZpbuKPoAxsR9PtpLPqsBj6zd4YaQeVMPa
EgmN1HvSpLJUkAfk/ySw3nn/JnodJWFxIh3gUwb3ca+GiydHWtG9RKAtz9cVGvy9
SbrB9Rass2XOmfriJQPQWl1bYWk5gusywFeLtYZXYgJPPtLYOaFGvZ2YOtC8RSuI
jpFKdIpOhMIoVoXM7GxFeGMPccKT9A4+BnWh042ANvtLYk3lupTQfchUOyRXb+Rl
TxVK4NYd65lLGuzXMoKRmWn/qKffTseL7eYqEA3A/8u4DNyA697+AncM6fP9gVMq
5NpoFVCAq+v1nFCdbw4L57v+Pj50sZMtL40EUHLyF7odC28+E9O6Qk0rhT0YbbFo
JE0N+bN5jhZ088/cNc4Vj0EKgp9jeKcx3XyG1h8ZjLkPKvLtPzlaPO90/Ocu7wBh
XNP8imH/EP2wgznfx3V/395CP2elqK/ayM8Ok0RZ3b0=
`pragma protect end_protected
