// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:54 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PDmakMaATwgZYW/trkQ2ciTwpA7dmpPxS/t7OqLTJJ7Q9xFg4dh5eJW0hqHjJEwh
/+XY7TKcq3dsnvAcZNxW5oEPqQ6DrZItEINMBipHwk5attD75qgl7qifBYjEeLcf
EotIB0EDvy2AZUCbHey6GET0eDVxw6IFxURo3wHGnJo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4240)
asim6eipCRmDXwPcPa2t/6N4+9Q5lNeSbL7iHSS/QOSrwFb48MgYRiIX23vDN9Rc
8IdifZSyeQNxP316Iiib/PtR/Ome1yuR93bLBgm5T1xt05pJpxDZYlugQREHjYpo
pGJ6qsp35tlto6O//5iS44oQlHvquA5vURAEu6NUMM4iYqIe6xFcOgEE+lANo51u
LXF3aKxHnO/nq2HspHVUcmRr+0jp92gD/gmv3RX/XjegR/rps6HFLtBl1EQQZAOQ
bSB++Doc036DRY8qDy2SfGwAj2Lgan63pzoJWYvbx4W/ZCY4d03yziMMqeKIdPMc
S5ICvphXX8iuS2BGkIVmlXe7MiioFuzVl+MO6mDntKMXv1OBAGyyC6bS+7k5UvbH
K1XUIllwkD6VDlmHAUcQc4QTct4F0eYB3mta56A167lbAZoSf54X5vwkvIxdxa5Y
qLzZIeS4y36pZYKmznVCHVm0tAuSxFkZ6zQ74ksQVPuI2vDIFVcOf2X5TN68bHrR
kU044ZovteIwF2v1oTFV0ZVNDG80v4trHiGpHs9gD0PLKpsfkxgF5jIvQxROuwOH
R/YDtvPBSw/P0HFmEabxB83KP2QkpylfvHyNuhJ80COC68NjaD9HDEOEr6xo2vcC
XvR1aF3dKHx0TR4FvZ4SUKyLqnxnXhkZ4fR97aE6oAi+daZ5m3NymQvUCIdxeg1R
o4Cmz9S56U/Xzih3LnS43KSWGcgG9jXBwzOVQfXUIDnEyo5eiTluoysBZpHtx3Tj
RLPg4XIGPgzJTVf4EHbO3qjK/QLRPFQw9xCAS4agWwTIaJYvodtwJenEpBloGvK9
oGloERDq+/pAhmPMDxEcWEwdwvqOuOCSIgy0y4ICLdo6u+wcw/PVR+fotYnKV39s
SLS8schVGBciCx0Z81c8mXKqgpmaZmot+zbzz594wlkGxIAuCA+1RxePcaACrNek
oFIpOBnhHOorqM+fiXTTAIN2tfKj32dWviZM2T0xzVGr3Qk2yD6E7k82AD2/qLQp
s04Q1xCLgyzp15Gppgxqqikd5ASKg+mMCAVk8/qb98dHMLbL+0gm+K8FpsrM5led
9ybUctTYVeIXiryB/DTfw73Ij8xXZ1w+VersBI4bGumap8fub/F8eryqhHONQ/pi
KFTnu+0f3CmgRcYdX/upKODox5BrncTYwlrNEf/HGKnH/kJPKO0mqArjzDsOVfjI
Svc52DEOevXJDSeorjut0eWiMwchtW2IIzl6n5BbjXFGVxzXtTFMJvZOOwmTPwRN
GU0q4JAvi95kpCX/V0EMWyB41xn344A9ytuk/WoBnwXfrY9XsSR9zGiGk/0G4D50
9gvU9IuqZ96w2EhvwtWrWDt1I3FfFab6gvQ/+BJ2qKd+tQwkQD8O0R0kvcNFlBkJ
IyfpeuXOAFKMY5k7Sf2acALmsqdWZ+QuuAUdqTCwLjhKuHr2xt2hNj8che4qe5le
mk9Sg0/m7Q+GDgvEqEqTFjRBTJ4XL/W7zCDrdqcNGoQQ8FeAf6wiDhl53CuT3ZL+
tcv9u2N7QzrxrbESsx18y2HixD8VKBX9ewZpRocx15KtuVoUeYA5rNmz40MKh9qp
DM5r8nHX09J0JMsWdX1gFN9/tSeawHco3BX01kvIgWeJeZFNnwmP2FKpvkMIWvwl
bqDs3YD7Oczu4TM1v49CPKPGJoQQ/xaoLbByuhqosTjSpLtFRzxuiyyMJ6t0M9/0
AiVXYASEFNRV7hpN+GWRIkq+g24hTgl5Nn0bD+QWclrKigAuywyQAKtU4dVc/IbJ
EpwIhAtsUSIJMDjtPajYUSsmq6VcuJa4UdqOYFOAI46uUFSEBV8KIdn1KAZDs+Xu
rHwFOC4fCHVG4TGxYo/GxNBAkZ75alo0HuFDGXDLHeL37iNj/NVWiuhka+bHYh5B
Qb6WfCzJpKuxnmQGiQZ4zzvJtsW4spbZY2JUq6JcoR9aCjHntYKMNcxllXDuQ07w
LSzfmsKsl4h7qa3ZmVHItBpgNtA7L4TQv4mAD4o7IOU/ruDTGjtBCDLayLuiGoNP
HwOTGhBa6AdqJX8A5SnUdEVQjg44mQzLYxs4Nx53r6rUVDzNCBxF7M9oFjT519ka
hfBEqNc6F1WHofHSER3GaXhuf545HpyhKOkSGKgDbsEC3zwSJUkxD/jUlWzSx/aF
9xp+mEFljF/fZKyIa+XIRtx/ZEyCvy1R5Da2UekCDiph5OX1kPOROdxE6twr8ENk
iegyEGpkh01dAKs0vPTfk4Jt/m8FNZfvzKlIr+SS3595bcm0O6JjtvQHd6SyG51n
DnvpH7JJXX36lkqiZBd8E6uu3KuN+t8nKc7yyDAOfrpsoUBwjE79s8KxotBhzpqW
LjvlWKnaglF/h5fRZTqHL4Ypa/OIrnz+FlhAd5dxXEJeDTZY3is1VanDyF6Ne/9Z
A74AiS9FhMXSYey56QuqXrK7/Tu61SnYmaz1GcMz/0ExFmq4+lyQz+eZgf3iaxyo
lzxg8ZZBOGYHZE/Qxs2hVwZuUu4K1UBUtL6QIH+ap9DPoNOoKp9EZ8FRVUEKY657
o6ZNvJrFrHsPUhZCGKZsCaJz4P5kyiCJgHAdwu9cjfh6dTVzsBP5oVL/lk4FFrPK
Yu8VHGLl4rZgKHqgIbmaxPEYnwXFEkcupNnWBRWZLzXN4f2/RCiliCjNee/UCpLG
GW8oFgYWPzH7HnAXDcYXj1k2SxXOPOs60SYHH+2Njj1i6AtctNfdh8kqgR4jTMsv
wHdxYKEcP51yY0YNDykM7v1CD+LaCMYxOkq8G5cJfSVKOFx3pT+/9iBrDVT23HNg
wUThe0hIixW7DcCg2XRaaPS2qTsaqi+KEEmRJoCTPx0mYzNLq4hhH4o3MpigyRhK
+JVXcjoiCDR378VPkEeNgOEAqPq2QAZFidBz7Ef3FIHSNMEKXZmbHUbjTPDv6uiK
LK4t2bAFsTrAk2Wn/desm98SbeHtSN+dEiiTyxbjPxVKBHFMF6ge0zovwNo00mBp
ZGV0ni7nXNuCqz89Jo4TYSVlW9H88uzJEOH65lF3dMvTQfC+KQKWTk4AkrXZLjwi
BYfXe1Y8vZpQsforyciyEVpuJEi4UcK/md8xMa5MctRSZ9ynbC3J+NyNj+gZHMIC
eZRsdhzc+EVf6Gfxx7O2LyzDQbyHtWiRV1uM2kkLItyEZQyh5TEKQN7OugCkm78J
yCLPjRAcUR2rW3s86GzlUg/D5x/t1PzfGl2z2znipgJ1Ravu1mOxTYGpxwrXxvD3
QxJAL3dJdywcw9ocp3zAvUU901m5eQ+BWek39Q7+uZ2UlrvI11H+We0ImybLj6yx
JbVLGONk/DZmL/lfHuu1n+Dt48cMDVGtKcWQKqgZPLsxMtHrp3sxOqgxYuUvjejf
zkdCBSaPcTEtlOzw2qUWxwzauuUidv+j46rBmvjUVA1ArjzbwdlsU+SPSqNsZw25
D1e8qsD4XCLasDfKxuRIVBx+E6X8WwJsiEAEw8+qz2AU96NgSRDI0t1hv2X7Mdif
WkMqUyoJs63qI7XwNGAK4TlTS8z6SFaoZgqcqsZIRSozW0yq7gomEXtV7T7bdy5s
tLN/pxyawE2Nd2KGotjfdx86991jcMLeKqkJCDOgG9Y/BJHX27HiGP6UHxqYoXgi
jPimif1D+KN3NuVDnRXAFboyarsXVOnidnrs0+lvHc2RjIsOBzFiZ5WRILnc3PS5
tzfvWCYE0NvvK0D3Fm6c8S0oCx1TNPpgz0UaDx6hp+yywwz6OSXGg64W7cIun1kn
O/d51MkWlXf6Jqb1H5pAYADjAr7jhbvMFDnOIh7OAFT8fzjhFQUKml2cqSq8Gnaa
bf5ye1EZyMpVD9rFfgS92M2r0F1hfqof4Xah1HCpgROZscQE4XSKKfxxWQ44YHCJ
wRQXkFt5EgHK/gPB6dWBORo3iFc7Z+pWkaDGL1VJXxCal7G95uLCgAGnrJNBXp2l
qIR94o6YB5bzh/Y2HtOQraZb0+mcj2zf46XdO5u0w85gmIgNpZ0W2CpZUpHy7lKZ
QgSOwUe0NeRg4WELO8NDAV2sOmjOp6YzpmB8g1YbRvfGrntvxON0zbfbfvkzLaf4
qcitVXVUpNmsJlvlo2+iCHZ2M7tGgQ+1TUh4/1tyflGHAs4L4cp0LgcWeflHG8oN
QTGGDRPbmzUM2J4XLddR20EOm490lnFsa2ii8ZSY53WcGsQUbWBygVzid0pJJ8RV
+Rtw2/HX5Q+iJibuUj89TGOuMq0khfeQ6Lo08BLUwkCff6hzKjTpaE6Ki3SM2HFE
4riwn7KWNF0DXSqNbSpRNfe81JytH2vPMqf5uMnHw8HUpxIYeq332WUw5szgQkqc
VOlsg1Lcis1jaNAmaquJ9J7td8VhiuIjHU1r8eIDs8bSwnortM71mmyhIkaizoD4
T72OrYGXrwro8Knis7+xLoU96LRfoFehnsTRQfjUHO2eWQ3ZhkajIjPduE6tHOY1
O6IFaKbpKU1G8nneXQuWdIVJZ2A7PUmn9bFoqAf/lwX0bBhNJtkKyMA+UV5yapdT
yCiinS+0nm0XM0RrpjNSvfRFHB47PQmCjoK7WzFsoBgQXwRK0jZlpzXs37oCdE1J
F9qziZnNS2NoBvTMX2WwnoE2IR+RbIEmL1jUBKzcZOa7dY4hioeApNPDeGRI0Gvk
KnxTrfBf8LUYP9HixkrikeJOhVmeoY24Z7IVXjVtKmdaEkTjRxF92D+QISj7NxJn
cKGYbV0AP7046jRDwpr7HSMRGU9zRprb82F99bd8nz/WIBFWMS+Hnr7ttg9YeQvI
1JGcbWJ2x2HyOUf093mRAsxiiwO41uPxWpGbyiDMHJHNMQBrLk13zlr0GcrVVRec
BONyRyGOPtWoJOiuiH5hwCpgUIc6lE777vogDJv0C5kTp0ZP0JGZaqWlyrurUIN5
4wDbceRWji4Pp4cvppdu/bYLci8CBDpdWV9zODdDaNKNlWwEf/lDZiUV9CWe0phW
7Axulsqapr3m5rRqgSO3xI9NDf3ONNIr7tH5InLVrXxb4/0wIGZzL2SHEkzsV7g2
U0roVIFZtRFKagU2vynFVDJ2XCaPHwc4tw6dFi0o0N8wwNkFNTPCFAIREkMfPDSq
taL1ajhaOFYBqDwhERHj1CoBqlWbnXOZyhZHY3eQclLGH5ot77XOJly3rxRSr3jz
gjqQ9VfDRGy4AriqvjlaE4MQljrFZTxJdzDUMYehy/pWO9Tn1vqTyR5vuRr8+gmr
AVttIG2MA0toT2qfeT90HwAhco/x4VvBwZ+dzmJQd5soQbmwDv4zPL/dNMJBRWAC
hD0VHI86zN4NsxisIaIyxdzzNBV/zzqwfEuEVQYfY0DE7Ko0eK4Yt9Heas3e2tac
VgJN0taZ8Vw5k/eI8Wh15kZxxoZS1qSKTKfZcVe4bYVBZ/7Zx33+QJI9Q1aBVAg3
lcyq/TrpIgYdfKJT5QBIhWSZs4aSqB99JAEWC14sXwL+A8YgDoxC756awZlFW3DX
uS/+Nkur5XA+qmKvAxEuFKipz7+mafTBpnNMx8O4HtZPYaaEzCY8rsvugD0QLJ1o
h7bRv+MfgfqgB+wdq2cgW/jDHNy9rhs93J1Huzozc9rNAOK7cmUylPpguXQ3nzeq
+eOQMvV3aH5f7NFllaXHOQ==
`pragma protect end_protected
