// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:02 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
klFZikRvFLj8oEJyu6CcNyf/bPj9QN2saK0hEdppSo3WpcQ0ZkixUw0NHXmJDAOH
13sKobPrjgHvB+kPuQ/mXu4855pfozCRnjPtDx4ptd3yWVIZ/xIocxGptG21XvzW
xD1V5s1+y06QwdUKu55QYMGdW2+m702JKJPDffNXK8U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 82048)
ZZpl27bfQJl6Bs/YRkgTwtp2GQr1Zu7SqeIJzMne5g6ExvZEd/T6LLFRbIWNBIyE
SKardlZToTksJk4Vxsonqxd1o8vtqZ3CZpO7OLmaEteUcZD7ShPgHBYkD7igQ0a0
IzgiG9iVkeK7RH7u+vru7GSTzHzfdh2D1aQZQZif+xeMwutq06Vfpw+lFZHPN/Et
Dli7ZDK+uwQ10/HlTgPNXh/1H9ecXzCweaynm7ebtldXfjBeCQYYBKL10V/ZWrGp
/4oCG0gQ1xf32p8G71QvAHy9WMf2Premkhisy4Q66Sh7DpaiKkYv+0DJ8si7EjY4
vD563swA35GWgVcGCqhttsDtC69GTtbEs13DJWPMkCOwzVZsjVteOhS+VatuyYNI
G7moKl0kYgco+AK8g21/Yh8QJfpN7CILQ1BeTEVaNS7+WdHX2nP9qUNsaDOaDazW
QCn0U04s48MZGSAgAnQ+CeJmz3WzMYtrrtNtCHv4HszMEEu8/k8SKGo1I57bB/K/
QB6ne+24WYtZxvCSYn+BHRzhz5VFdQrLYXcLCu409geXZvH71fzpKIr9IYsXPBBp
Lp43WfPMVfUxrvKPRamT3AO7Gwku04xD0sfZDysTmAJsCnz+B9BBrm19c6K8rIDX
jnIKzSr35n/St3bk5nGcWvnXhUK1LbDIi2kmBIhkMnxGwPuz+4QioauFIKvWhHvP
6x33ZMku25cCHocxpPpEbmXLAlkwTRrn2Hkajg/VJn+taAB4dT4uOpdQotItEoUm
/TYJUquHUDNBQJQIquqxu5WEqKpZy+frbhMBYn3iRx20CklkImNPtCGgXppBqtwD
mfptT6iVtab0jgng8ECODStIpi7e/T6GE0nmXGA8xuHUyeCsLqMTm7/KrzEdU267
Rv57qY4JjLnOp/yphh9wdFEjYZcMOKdhqzqdSkYooUMYBe1uLS0k2BypUhAZRli/
k+HrkPYDKEM9gojwzP8qmk4z1RJn9+jD5FWN/QToAgf+Q9YiCnd8LEg8xJ4Ab3gI
1HVZ4BECEZwpJ7/titdQAr74a3M2pJcZr31bRMYws6c2R/57zSnYYCdc2hMCIWP1
ifzsotbI/jCEwvoZdeUcNShabFZcpgdF2kZvUQl8HHRQOWLDBQas0yGtE1JW76F/
WcC/zkW/9Xv4OcI1Nxs03Xdkz6r8A8YgWCV6MTZoyQOjaAs/sDzTRdcmGh/3eR8t
0O7xWvGrLD1ktcOmiqKRzgguEZ/7/oWcWdrGzvui/MNZhsV9jJfXKsx8AwWF51ty
9KZE+t7YAaDljsNsXsIEBBGIhSo198t2a2vzjR+ChPOlEP3moxaJw8W54SSf3qA+
6WkFjf0rePup/oefqkzFMd13gaKsbhjwoCR9ushCi8et27wMCLJSZy9LM1+6rhM5
Iz/TDK5pQn5lU6073TzglzpV2lVaOtqBbHJsJ8t6PiiUp5sk0uLoOBbXvCGDteQQ
9QPot5aotwy17+10IKaGjgcYtlVQt9ro03Mw7Fb9l6PJH32cUPHGUC7dB2sdAuyb
/YlgiExEjskOaJdra/BJ8OCzE/dv8FUPkJxYxM34fWAWR3gne48GEDwJNBYzXuTx
bZ2e0yZ+5R8iAuRlos6WECqG9vkvd3jhuexYGsFrC8qvsXakvJ5iiV7In1c9Y/AV
074DXMrPlexZKDZWyVRirpogBfYaDAqImJqyqVj188m3kBdlRaXxKhW8blzVuIcf
qGWxFsonTQTTR6GKGyFIloJaFuF/8MHj23ZNq80CDCpeBtpuljGg9g5n4TCbmJmZ
0ovxYHWzzQ2clrwu8km2p7by+pbUbvXUk1fZ6ENbc7aAHV8sWbJyxfskGOgWD8mn
d3OLVvvxX3Fn7WhRmx1Sn2Bgbjt72/5dPnxRCEyOWI1qDRxlDsz/J+Fk7fevc+0X
gHxRz7Vj9Wr63y1qLjUsIrFisvl8/Vw9TMzp7rC5iGNH5oQ+OuRwYF0h8yQYCSkZ
KXzJ4YmqqWiicxz3PzAzMdDFDM5pB9ycDb5I932vGNEm+b8QOb6aXJ1c4SCsKJbV
6gNdFqLP+PIVU8eqNgRKrv1o8ZontDkUoIK856TE3Wj5ToFLk8qZAwKVZkOHrMQR
g/wb13QZ66DQ3w733OPL6FOnkniFFbLf7B6MywmLZUyFgx556x5kMnQcQ4Yh0iJV
As71zIBRB84+NhrLqJHGCP5QxkmHU5/SwRkp66boVNpq/Do7aEI0I8ApMOA3CktB
XGNOPyBlUwxZqIcm0V2Np7btRyp+NJyqUeYaWFAVW9YzBr7BFjYu3ZiGrFufrKhr
AMBXHLB7fAt16xsSiUKCSWWVUUXW0VEMv4raNpH0uj0o7yQHtImQsULE+Gv7u4G9
DnQ+YaDa1g1MCKEl/CnO9EceYSKYgJlhypzNMcnIvdItZQNRX/LgpLuCw2eIpQra
64VgoNaa4THXoDod5bqYpFEXnllnkvO7vsqzfe6VoKPcXiSUrqFU09kJnHvqnZGE
EVCD/WbByogByah0MU5hVYyAJolyV3MHhcFsRBoUFqfZhCMy9k7qOZAdKgSdj7MT
LB2FR9d/TOlfuUi05gluc/EnHTawDWMRWSAkrwR9ydM2K0pT8UC7BEfvTf+bcyFx
Siltyyh6jvqEg7Qegjhi6QsXOSV6qqEk+DSBttUE7unYF/8I3JCodCCR/L1Lsjs3
a1Mt6/3cUsmk5bKctbS/dHvrrmyI/0dsmk7JEN29NcnuYKYH1TP0Ium4J11MvX5h
BDvs0GlHShzRUlj946KEMhC5gTYHXr3Yc4b1tzfDjvt3LAppoLiejmlt9umVEovk
GTauHwWTZGwmtEgV583LK8PFhII5NWhggIesyp8OrtOC2kb9Fmsp/p2IjBig3RJq
TW6WeBJxeISJ6kAd3VcbPWGnusauTQ3P9turrdD0UlnHAIOy1XEw13+GuhJ/m03O
28/9JSP14/0PbntvfSOmS9SwIXP/DgtANW4nPOp5YHI96+ut2w4iGH5VuHnqKFwX
/qg3cwhb+lFBOdMFz5qapPI/nysmlUBjpvt8wKxVBINvnnjb0kTWvncv502RzVD8
Uanv8Rm6Qq1ol3Ul51gJ6S/UQt97OUmLT5F4aRG7QES6KZqxoKXqQQABPPlZO/xi
rO/0s22PkSnPrsU7snAF7KYqtZbN7ii7ZF2bzQteBIDH7xI//5GlDmbFrkg2xWCR
+p+aw/slFxnoNN2fno5IPwDQCdxx7HUOgqYXwG7ch6Vq9WNtnQu5CDniHtYtttcR
E2uIlwnedXzojl3rjxT2br64oUkQrkOjz+UXCuLPTpRL57U0EMTV+ZupocJa+c6M
yPUiSJ0ap/9c+y4utknYe/J0GtQclBR0/lf7uF1nfWZxU3cyxB8LnWMm0HCuel3H
4f3JfVnHwzj7yi3UMT24810Y6Ov0YqDTRQ/56N5/W0MtWFHUMCVdwc6E/cB0I34N
kBjl4VW03rqEFo/lvbZmWFkDn3gXDk3rxqLL0opMWkvhS4Kqy21L9QspmGN0nyyH
lh8kKpGoeatgmUINegO2tsfdHPa7nx9sxAJiPHOWB5y5x9iGifSAPlWg0rJo4LYa
Lvg+f7oNfJrv0ACqwhJTgxoL6FmtaIGmzMpaKDmbzeA1+uTlvpYuHqMeswQc58wb
AOkju46zMlTmgPGWtQBahHdYh7cw4lgFPsQxRX7HjI18XrftLsOftJ0Yk9J/tvl2
CwNV22zC4MbZBFa7WTr8xS8hN3ZTgxahln1ziNPwUe8/QG44jJj3lo7rFRvYCiFB
O+x88mRQbrRQGFfaAngNIKDXGN8WGBhtfYQwh/WZTG8zHqFaUR5PtkScBGA8axXk
E3dyiU3a27JDh5mJez02svQtlL4w1gGIxO4jvczgzPaWv+WPgMfW7GZPivtEwcoI
+/O+N7CuJHoMLqv1BO+3vw4pJC83qIQ0EEMAXYmjV2HMYh5VCa4hS886J0PvUSYS
OqEQiD3mHHB+kPqcvFi3uURdw+y3N/FN8K/oHCz6+yT2kN9xCKrkrDRC1SsniP99
lacx52IJfaYDrmS4WLcBXHOeZdDixpW6o5zYmeD0V+ZUXi1ApiuM+u11OS2ieu+u
uvKyEGLthslf6QzAE58CMOlkm/DrW1IvteBkG+lCxim7/RHcR7rt3vVS37MqLVuD
7fyo+FVSILgJF0YFNrlLwBXgfZeAjIG5p2jDbRHJM+U6bQ+bn9xNRDWydLLbAbGw
54g6Dxy7BfRIh/ALvzF9paOHYXi53Bh75XJhMk8qCeKhW31FydBCqT7dax8XVSx9
/3qfcXmO28zLHPmjcsjhRlsm/XF59ynoekhvvN2zSWxWdUKHc0SYfR6xbKRRhlhX
KEXJCTTVQebUlyrYMOFre7rK4+LCKF5MAW6dH0d8mrmSa85xcWGBXXwacxAJH9k+
CphYL0UvQpszMHxByh6hXqmoHPLtxhla7jenhENzkiXFqDcoSInIfwUNzDo5kdBf
agzDC5AjnIo/EWZnkfxzRKJv93oiejQeVkhqdf3tmetpiWeY6t3b22KmEcvO1OXi
aI8Zr47ZfwKBqVp5FpLA/0r7gy/moLs3VRGx9aOpGHD1fUNPIVR2rOtUZ18oXrsT
NrdA7S+l0GDDIH5yelQQ7Z0anV/TrJcy8+kRj0fMyGGnCtcs1ppVO2tKq6LGGk+D
qi29cGNl/KP1xdQ/07XzgAyroNc7u3qh6M8FA7pKouQH5DYqdyAGLp+ZdA15CkAB
jcksYHhhb9Kryqj7AUatFwS/7H7oDcz/phJSl+tumKe9wim1MPfP7F8AZ3mOxwXS
ce2zC6NX70E5zwRqqv1nQZxgPkoddl0JoxD6ncDySDqd7qRW/xOa3OPEU/oPxO4A
11vqvcJUwX0ZwIkzQkqgVaXI/PIwLHh5gmlOZfkD8ftw6cb8+Vsg5PHvam5xdWwo
klAy2B/6ooA61HRrHdH5t/BPUK6EBaVfQ9jU2HUczB3+N6Oo2AD6M08suPFa6eo8
U7lTsRAp8HfZMWjmx6v/8iqwcfe501zeAE1nxBj6NDe/BjkvxDeqk2Ij9DYnutt6
RSyshIf+jOrL6I79qOsC27C2hNIGWWMBYuNVVdwhijdXy0FH32JBZXR76WEwJ7qx
5VLvHX0d3+n8/Nh8BRQqaqZBxC1XRVgQCBb8ezjuhYmmIsZYhWQpN2TZjquamvqD
/zdoa6g9eFgOSkJhIeGqrYmB/drvVzXlDNCyQnauHYLTUsZtbunbSf1X7DpqbZy3
pVjhvju+EPS03bN16C08n1ZaZnQlIFrUt1qpWdENkIWaDtM3c306sLwP6p1p29sG
mwWu+DhUvTr7DGbpdv2BZwL4ePw6fS8EhVzle8LzojlVTRP49aIBzAKX+78gdkG7
CpJnHvL/+t7HN8I9ccuQxHED/C/920jauXu0IgXMj1okp0cfWYe5OkoNSST8LJx9
KvXT6zHUcvI+UTZHJ74LUMdn4D30DyTwXm2ftrY6Rx0haBJAgtHPByn7KvrTR1k/
qsqMEYdCnhY4d/h2/HKkXPwdXWYgzon+jYxrox1iuEN4wSyIX5tddFph9VsjoNza
c8TxGQ77o1u3oIC/k0v4kpic4fASGHcAnClOWssRMKqH+FLUX9iSNL4SygBnXtge
RyQPFbfaNRFxKNOW67OUllZCcwbXW9Zt1CPIIEF5xYJsmDFteDVq73J/2EqyYFEm
Cs9yHl70hLD0/HZSifXPBdQuJMM0KfgBMnqtmULxuZk/MPyIEZYkr3fpYoUewgq6
vOSDvlyR8jxzQgwvzvt516pZNNvwS80a7hUwHJPFaBR40wsvA8KAmzByd/2U/XGC
J0hEy3p/RldVadjayJHqJxRTkZM+b4tsDCO+5BjlJcK6pWytkeanJQ719dzUpoSI
XsmARqzKthtpKE9lyZ/zKF1xxmbYN/XP7giadlvYmsUi2lv4AdO0GphodYCDCtMc
f+3RxO0+rcWkoLvpCqe1YeN1FUoYFKX4bmor5VY4Z6hZx4wPyDU9yKYWPAdp0AKS
mMxO8vkpy75zSI8wdLc37AmYPqKbfj1uJLoIp6eCFH427phz4JdnC9zgDME3uD0w
kJQvtM6o0NWMRP1vpGpLGBW9pA2uu27EtTqgqf9jNcfsdwyKB8kl2POK3QWPKZfc
agAHuMIvdooaOfdtzJpP4CkhpXgl4d8LrCXGXAVaGWEOla/M5gMdXkWl6bDHr/vl
HxpMQBoxVThYLh83iM21jxTF9yo6zRMxqnIf6bFus1bDvIXsGeiHOBLAwLdva4H+
KpdIgDzZJ2u4Q7u9LkqUihtOvpVHC0JcA/3f9sArJTUamjkD0rNT1Gs/G6pUWbTb
eO0ZC56Bzem1HYlKBbx8BAoEfA6hwHhLPxbpAWekKB/g88x3VR8JhvjT0wFP+AYO
eNXxKPFZLHZT339DipxsWe5X/EgcMZOJh9MlitZcim7OhJNKixY+QLRUBRGzwjjS
B12IhzmYMn+zgJDBavBjqQWIxOhNRM/Tm4DxqTk+nLfHAeS3ErqDRV2zzJdR1J72
rfq0NesaeQ/0YLX1CK70iIV5c+mH7aNXAxataoR80OKSAps0m878YJroQlwt/0HR
ZL6C76BE0PQOYLVivIvQXNfK19U5buEoqMQt4lld8cMEp+B2mt2yEyWCInMRjNqv
q56HWgCgy1BX1wPgEENnuwUqcoUWFjZdKR6JDZYd75muaE3Gh4PqFVqtTMq7k8kg
nbvn4HW5uqYxXB/F5ylVFqgtXRP+8TVNPu2afhmmQuCtWo8Q9wcybgCSnFGsvPui
VDTtPmcL7XeFRM4auijPpIv199oyaHwwhy98Z8h86bu9PRZIo6miXKWaNf627J7X
rTSGZn8pQ0UkwllAV1SWS1PHaIiEl/Icx39YVPU4lPAVuyY5Ahu6l8c2+1rePRZE
vI8CTteYU0Ng4okHX0pRypGbHHqfkrT0Gwnj3rAnpgFz+eN6n538c3eFrr/rewLC
JvT89jhZP36mJu8ugZVSnsKPHYjt6+wkNmxJmZ/ZncVe0lWA6o9bECJtXZxD8EGb
2FGhbRMnP/Y5rw+vVzgXu5Dcypfr08qxwup4/oa166E+LG/IW9fg13oaXTL/QgBZ
zezJ8EItKKVJdEcZyoazr/E0BmxnmPSEjSFVx6pZIBpdQaUNqW2r85XgCNA5OBWE
22I9zbFr37czH418eebDen2zerI6PyYQ/WAW/qiXfMiWUD/QcAmH6ZRS5ZhQEVbu
4kAqdApyMlf9Bgqq4dBmiRuOFBSQg9BBXwib1Qow48EHwbz7HCqBqiL0omzfLJTg
EXqSN7tAMiJPelHKvazIIJErw9o9lf357Pxg+83ztt+aYw98Spuscw8NTP3lv/R3
a4Og9KgtSVU6RB1Cc/wDzS4VqIqUqyo2FWqXuh+CPDdMesmWrWTfQwY93iL+Gp7E
4jVyVEyEBmMMZ7KtwQ4Fu4zT13PbZS0y+Va8/WNPv02DW/RnDoOqGT1jsTS0Uop1
mfhg71w3xR9xve92daBP6KnoLynS76wpcbffbZ/VUFF+OSGNlp7FwqvNN1AOMz/X
2zo9AaiSrhDojQ1nv5vK0ef9aX7r2gQ//6O1u45SQB2nbpMDuXeN7FCTAKocGvKl
UCLthj6r/z9R8pzyZh+IaNCEYhUpxb0dmrnmCd7Zqx6/2P5/IpsrVsMcrykhmbmb
BCidTR/lLroy/RqcLbrooCOQ/WbUE2Rgl52pn2HezuH2pkcH1vdLvpwPxWqNyYtA
UW+4lM8VT39jtqlV6ksY1/lPeCejfeNUEuR2/ie7KJQz7x9cT6dD4K/oaPmmV4Ls
9BsMQhqHPD3BXI1CSPvE7unb4hhGeVQueHEXBOI9yMHW4Okq53/0KnkQQcJYW7If
Rb4Nt9lTw2G7sOGtNEJQVrV8JUYFucLQVerz7s5y5NakBwdwba3htpZsWy2R70Gg
6XyhC5g0/pUJOEj1hQfBpB7VAM6DxKlQDO9r0blKhb75A6slnQP+LeEJcgZBKo/T
WMW4HveK+WiZsxgQ9q45facD5c2v0IfMWYdLHCDEg+9QK5R2lylpM3BAHoLQC9uR
ucpoSzk3xZszJo2usdsaDcz5skZ0TrLsNob1zpV9Tr7eX8LNMqaPBBCgZyV97H2H
rXHS99FikfUVe3vFBAtmT5EmBXgfwMoGnZmrNQyYhfzezW5FCsQCBvBYYp3lAQ06
7bCNsk1cym/62ePTO4StiLveo96LGjCv4uKb06vIjl8OnmMd/pvqPIGXQkq5Qi20
9FW27NbmV5LZiYsTISmcAu2kOLWRc8rb+WR0BxH5MC+SP/Gb8ITAmpNxYUHWxXPa
1gLleMsMrN0auS+X7m3v1LmoQbifelfhe+eIfr89P2lbBX8x2r0cQkeNuRhfs5jZ
JyFoyOH8y4m94GvPt4xJSQltNPyw6z90QBhXwNZX4Zo8zuvlLUY4btNvXzMLuJ1I
8OEiAyg5b6cXnH6kRkK4/de4ZC1/zfZ7cMcg/nD24epZLEf3DrIrKeWSuahh78xW
gXy9myX3sqeVXkiv4uS0BayDlt3Hn4ce1YZ91Yr+T6kVfxjuXbWEZv+29ydrQqhH
tBnXKz6zCiruCoymfoNMJfyX5FOd8m63Zd3gX+mZazFpa4a2+J1Hp7L0x/7wZCZG
myC5ULWdK8VyqrOGHa/JL86OtwkfZdE8VU1pjZpKFTNuWv9txoCRdQ0Zlexhxf32
QlXo0KnyoTLi1A/Dggf4Uf1yO5EX6N2v+EbHJIHA8hqqtcmpld7ENSDuzTpGVrbW
H2BOXHmBkmtVODAgn4gyG1CI0pzlyUJiV34UBz0T9FvV3TsWPa2zqYIMCRQdIq5G
fg0rOkqHqwGhK9foHzsHdmKPrXCeXmjNBCQIzOhwsrxzfU35kmrmjLpgfHBXDoCu
W/2Kstfxm2T6tg9403OfV53x0aWy8fLbtjPiZTnQWC2lAXWGq8k+IaemfuavL6UR
zcZOxgkSiQzck6e04hRsymHuB6QcxnqDepcxCNNdY35CEACGvbUCZhgrvIF0ygrj
/geh1JOSvPU8FLSYR3MR4MEj8a822tg6ih3GMxJYje40V6zoOc5pEaggOWZ7PNzy
CqLYQb0E9OR6K4xhvRqhPeBwdqqS/NcNfRUGqYp6NnlRhL4Qjqn1s5iRxHdCVtIX
WodbI3Agn4gX7Ewka8b/UQbUtkCoEARbjS0xSl7b/+YiCtP47+vsTyKvx7MRcGuZ
F4myTZBkhLAeltiPh3xhY1EavugaS+BoP2RYbmaqvTekmje0R5L/KTQ0CEyglp/q
DDz0S2Wl6NElEEOqVQ69SyRU5K9o9D3ZX5LUoCZKZiBlAm4B3XZA7wDyTwMMc8cI
ZkbpZDmGvqiSKckfDNhRsZyS+Ih4/CmTA7UQ3M5F+InlXPsG0Iqct+GRQuc0AY9a
WeW2RoUQEppMNHIXXiRg9KCzUtooxccoQlO0T/TmLb61C8uOMxz4gHcKrAy8muM0
cAfDWMAUADdshrz0ff1EJBOZSE9MVspSyG1UpiO3fzLe0Yl/SYvAX7ttuJgynJju
DjPFB8pW151InDr37aNl/DOcGar4N3eCGkokrOhOXmomGsp66QRVk/0xxbnp5pql
xAW1+HpsGs/SNPUJn5fnKnl9khHLIpHO2Bc1X1Ar6qpaR2g/iU5Ru+Nd/MTqbAJY
NZb6z3RjoZb5nNdznVlkKi2d+Dmobghb6+p980Z9DQAQ7+yHbU5Dini0ESk3IuWg
K64isiS3u8i9rWdjWenS5Sah+O/X4RJh4cV74BW4CgrVENpCF2fszMqeq9iSrMjy
WuQoMIf1YP02vlSA9mde3leyn6+9K+ATtOENlF1kuuf6wVagMiKUTtPpjgMopeYl
OuMe8ubBTsSBaf8+nkYc/HKdq9ZPaN8+pt1X+SIcflSrl7zBY3klGVwHs8jkfYiN
2ig4PBdruMEFX9MdneeTL6DwXKJ/CHbLSH8OzBkbCFDfomg/69bIZVhsZnCdyAOz
tgF0YGsn7HOqO9z+sXkq10q4E4/qYNFt1f6uIPTdZlwhYyYFLlHQbA3k9fu8oajS
z7ASHbQ0TVrWFovDfnSsiu+j28L6HhNAgzFJImSxry3KevSIdIxLpwXo6ezjIgyG
65wuREV+YRtdpmDvoU6AlS+mDAlbixlvYBFb3is0fh54zgRnOgHONiz/d3cl8VpC
aFDk5mXZjU/MffWvoQkfLWy6GKdV6cPQ0it5mU4b235mGmzdyM5btgHGJ/z4C1z8
upvqZAOP6NQaWKPX8mZGDbqKiLd9xLUKut64KqEmxBCFQ/MwER2x/ACg5u+yi9Ug
HAO5+zHbtk3x2UXBdWQJj1cR60zu+VfFYXfsiQBbeR90azMSbn/ZV2kmkKPQyF3k
Epir3sTzlCJtgSziSDfn+7u+xiq7ls9ndHskFXj1Skyg90z9773w04KrJuqJ9ruN
5RQCg1o+4BJdvfPBcuPZDVOkWCkD3G2dZkdKoj7a46NrVcCyCk9LkbITHRMFDcqA
j3ilmROPL5m3DC/0iXRqs3w1/fB03JCW+mfe6IXXTwodexzff3bJxZY2nlYUdRna
B1dmYVgTgcpd2hphwQyxUQrjLzPQaU36D9bMACZTzCAb6USmdnZ/AEPQhnk5CnW3
azED4nJxB7LAL4ThdK0Yiy7f/Px+X6Onx8U3W+j1juVPcgLbQE6fAar4z97t2szH
f1eNIN+KqBahPfEfB8Vms+TIh7ntQ60dC639wItXhIe4oRif5P5xKShVE1n71ueK
WX+bpEh1BA4NHwiSsFefsGYcOytzGGgzJ7m7UYhUC/LjO/oaNxGq1h8c0J41ff/I
Alci0YHFqXjksaGcvV6JLbsbS5PJJpIzOANiG/yyWYhTvGJo9FpsjoO0qe8rL4JE
vdWTBVaILZm9cYvyeE1QVl/Oke9Z6pMR72lAMmQNj2Hw0zAc+ZTODHpWF1D44O6C
TSxhgNMwJvZkux9rc51zbUiajv56e3lzjRYEHWkKtM391Eclgp4Y1S2fDpdZiOFW
bTvGIcQtIklttDZNHgsmy+jVTSctY0ZTF7AmV4CQSUpxLAgam5BggWFjQXBJyA1w
vAxsjW69F0niuPdWRhldFh2zS2pEVUivfCeotmt02H3oCSQm5slNpPTH+2/tIfVm
Ddb4Gg0eMPJOFpCaS01QhldiOjDHE+QCPCMYAX9mUPEET9UQnweNt5KlZhoTNB6Q
BDXrmNrQKkqcDSXPrcekD4YEtlohk7FP1gJLDmYlc5tR4dfhOrEAimPTUFrB523O
clFRjNjQNZLPi3qBLxyhD46K7aaZzFJ2tui3RvfwfO2CzlhH7eWvxLW+8jQSBu6Z
P3LGbIq+i8MiiwFSFl7/jG2kCiL7ZX1k0T6OoGFWPvnQ338ikMWk6K/mN9+StaEn
PTFf4aqoDUCDZJI+VY9bl3YCw9TN+mnL98x0IYevhy92IJv1bSU15WariMYrjH+i
iX4UDbaev9NFAHm5bJCXrjUnA80NVBVawUq9gaPz0N80ENoirglDZsZDxwdB6NlX
XUeJPM0NwoDXouZj770l3W2KYN95sON/f73+yfW9cnO7yVeJYzCJoWn6Sxxljp1I
5dh2C8RmCoWIexSuwS4hlPrUHZUi3lWJMJRxB7egLSsWVVJHub+mYvMt0BHVoStD
txiuygU+En+muk5dGkUYXhfUGsN8fKJpdEO9fH/c5yldxxn7dbha2b4pgwn0uVH1
fQtSUM7sk9tLKmZ8yvUrfDqO6RNO2Xql0pW/T7735op3ifTyd2MIze3aVx5mDdSA
+1f5aNO7P2JhsOVh6yWZFsn7ZmhFimgQDJpVxAsNoOhOF1Wo/p4roGiMxwLVhHe4
X75SRVw0UMUH5MtdoRJBdZsbtuKFCY+PthIIWGdcBnsSKQzuDt3pfG9fjSAC3MqY
Tt1ZRAblRaEug78ejYAcVD1VAyUyOC4plBR4oAyoup98cznKKUqCKi4iM0+nKU9j
yZnedzX8Rn7Pm0azkORNdhOG9CN+GYJcMQXL/g15UG+0HjFs0X32YOloxdNDuv26
zmIuYK2KZRbn56iFvukuZ6EDi73fRpIQJrTXJgf46MhMpjpdbG5dkpX/Jspq9luj
caFdVb3o8SK/X2v/DYkS7ei1dOsJ2ItpRjPLDy3hd/3ijWUn0AlnXJASn//jQvTf
1zII6H+cqSUpj1iETsdlAtnOcPdDIz5XsAd+/FfU2PMEckRNwbZQku/tQPFXiGbP
wzX8eCKAb9dAQ8LZoeLfXCSyKC7vFzp4GkIGZuHG0ynogpVSJhLqi0WO8SLv5TAz
CkUxa3emcROAXjhqwvz+nHt5MY1m8pQpVJiwl1MbmARWXbKD07pK9dMgOseaLFex
2CU6OwYuwRhsttEje7ek/VmYjcVA9ZfM2R0Og1yq6tvLLC51ephLIfmAuGKDDsk4
6161i5TSMyMwYUF7wO0CktmnReHsh6pOjZr8pwMfJ7Yt1PDAH29J6wTdScgtkg+O
BeYZIGxTnuT+VYFn5CjUk18VKPduh6tLz2ouEDX57m5k7BnYdhsSMSw+YxHVPWH4
xLubCe5XvEKdQ3VE+CsPy7wXSi8y7KCWxwWm22RZasUm9CsRXNCATpK5viUJY5+3
iwrHtxP/ISqfIg10TEa0Pug2cfANyXkaVbL4QHPWk6cK3hOcc6Bo0tzaxkMNAhuj
n2chuSJzgOpxBlqhexpdvutihAgmqXUSkKOeomyBBUcWlsOeFRcOAD4YpXFRR0et
ADz0TQfqc40yNl4f+ZC7fqDJ0cM78f0I+lFvuqnBqxIZirnW6kXZlMP92KLJZ5bG
5+65v0getxR0wRKHSlZALHrTlrgTCNyUDo1zdUldpCedmrZmRnntXMQThVYJ3xy1
Ha11qgCMmDNndFJG4KqxAYgr3+cysYXJ2SG2+l3JdJE7QUPmKLMgU3J+x2x4978j
2t53hK1pe98k54s0UyF0Blpm8VfydNOoLlNFrwW/GQeKmcqk4SAGAvL3ziv2hp3o
/AcOSaK3Ct2I9bb10HM7MWP/gZhr9MgP+rdGRBEYDqnITpV6EWVIWpZ8/v++Yjtc
M3AyH6vViKpuZlLRmIY7ZXSkTejbXcmOfl6r4hsC5GTSYqVWWRAK6uzB/FsLBAYn
HQM9ej28zuFmagDAVvOYSBobJtJ1hCunQA1+gY7nLGc0qMZXH8cxg/l/aip1KfZp
Tj0KlZg5nDsGuTpnhoaLAZb6yboQubda/qqQ9utEOhXtYo5kq2uslUlvJ4W31AJZ
1pIYQBSd10Ebjd3rmSjWwVtfOjg8D5ET1b9bE0KBntJnJuxIIsGLRTi/yMMTxULc
nU2Gbt3j0F2sRgP8AzA9iFaXdqpqrAKB34EseYyRWGQ97BUdtj/9UFjElu1Esj5m
DLESzux5vHafLpUFl7bcDoz7GA1PcDLhr86EY7hKCeUYid6Ut3w8bq3hNCnZwokY
FVRO85lzS2jf5AUgc8+Pr/5MOaYkgqH3qXHTvFkKKQsB2lhVs9GPY921BASxApXv
XeviSI6dn2Hyu2NPWQiUtFTOxePuvy+SSpZlYz8aOg0CLnLe2G2SQaaZUMn8nhVJ
QvVn3SNs+3X98EDLGPz7qqChuNx82zW80CTfe2FMifzXAZYn3HzN8I3AtVt926Ub
cu04DeqF1nxI68itCJYH8+DNqnxHHX/AhrC5AXwmLNPP0ssSvNsAQzDw3TLDwNdU
2Q5La243Jeub3Pk7tW0xUIsijC8SsNV9SxwTeXy8dniaB+Vu/YKJ3RuKt+iaKFKr
n4b1HJ63NCXFfl07bsR0O/Y8Ku4yzge26SRDUAhWVAm3b/F86a8pauqiLyOAVxOe
a0B5NC4L33HVyUhXDuZ0Az1onCmbcH7ZfdFTVQuqza2Xyb1aVo5+ZIdKW+x42aoh
MfzVFovvgKT1b/bULpSbavoSQzBzfTkScOM+OTcthTe6JGuMeZTDD2bAj2JOu7yW
0fmmoxZnyTDRR5LpW0uLnpjRDgY+l0arc1B22TXVXc5Er8LBtMwM7IKF6dBBg9/r
eZzpbjg8RQLLjYDln5Tn3Nnthnl9isWDCJkAzN/HV3YXZXWhvmBnXveuG9W8+8Lm
9mo87RolYhp04sX0Q7CiRqNd/RXk0ul9IaKGRgWzSt+yggQPVwr+LI++mmDkVOLb
deIawlrU+FL+KkE73fdCjrZuBMnYlxqKzvtn5EaSMlVHNKNgLk2O3IfJ0ZZ9sRCF
oWifZKcXoRp0OkmfgytQcuk+IOjHlSEWk0Nc5DwRqZeSyqQmEL2wTPJQqDi75Pez
pnQLaqQUokTe/DX/c8rQZNP+TqVsrbpFMLCcnTrnIDXQBJDa9bAcHBGr1uCnZiIb
MnjiDjciSWj6NjZtI1Uc856lGNAlRT8fj3itbmuVZ/gXLFkji6urOzbBrSKneTrP
RCy4gA0fcf7TJYi+5fYGSKmefz4n93G5m7dfVAyaUoG+kSuUv5QXOLpoQyugfdJ2
B4J61jsMb0zbdrJqMhpQHUu8sXw39eb267XRycp79WtbVZvU8q01DRxkKJD3hZBI
xLh3/pGbQK2lj90RKwifZTL7P3weoUitpHdoNqv5D1LdebwCdkooglF6eL5MJSrS
c0O6nSHakLeIN7nAtkvnRfLgT4iVjef6QUl+xWAgIrJSLldtoewW1Gxn4ClGgRQ9
ERka1olVIf2IGXcYjmpRtYKV+dmrnsYYGYGtlFgFa4j+XJ+Su++Csb1Co19Oclux
w2mvDwrRj9VRbUCrTHmDQdgsu2SPIoFGR3M+yYsPKvMpQtD0TjR4KR6XqE8YlZmZ
DdnUSYDrRTOCmC2IQwy0cWk9KLmWT5duq2p912O2sCjH2pHab2oOIX44eGoyxIcr
YqPq7VGwyZuoz94dUGraOsrJan3lLFutIF4c065d099YI6GUuLn0VHIJaFms1Fj/
/aSbjO8NwDGzrcTvAxbg26BT1HE2xCnaZ9i2prszHNDc6lIECE+Hwxcy1Rp2G69R
5yR57y+hjE9xTRN4clux9Uwlw8O5+87w7y7dJgUCaUTMGZNb5KHy42zgWOVHa4lo
fDQ10w/3yLgftX/gbgHHGTux3rui8rhvvGVMZ+od6kXQOLo8XyCOUdTViSYyq2OD
aPYHCDqcvX+f2k64jaDyBkaGqHAEMmlKo6BunlJGuHBFWLcCdhXS9V45N00VoL+l
TEVIc5DdPo62BXfHS99QjH86AfRpzI0xea2PfzVHHiV7CzAWFdVYH5R3987V/u58
65SAwuYB5D7v/cRU+W74CnVf7QxJXLYamFVdZKf/8xatJlf8o+Dx/h+lQwKu/bT5
yn3H1t90hkLQcer8d1jIEaNpwuzRdHx0sOTWwm6zCWjl+2vb+i+IfsHPd1IG0jj4
NzyPk+ZD8mWCtdBmBsGDupORazA6lWi6fY8y9N2DZnzR5JnMuANaPHAQ3U8pxfiG
ML0EdwTwbLhPCkOCkevlwP/DbQ6H5qxqiOj+f22b6ghuLT9+nhnh38Ot0tAxuPs9
zyYYcvNEirRNdgcfC5apDN2d7BQaM8w5ylhaq1jnSKfWEfPOCx0piZWKpZFwxsKR
rVP1f6720Is7op5ggzADBLuzIqnhTck5vw5lgc1ug65OX0pDMhY5g36Jv711aL94
Q5I718L/D/0cM7H8bqA0TN69XtoSKD2U0SQ7FAvKomx3oEuVT66xJZoIsflOjgr/
7MHkLnHv5iX9UwgixEsgGBZ7GtYhhIuJCULy0r4NsNGkHSTpx1UaXxtU91cnnPhY
M+2n9it7b2DDtKYPMN6yTYJ670zKb385MMMyFipSkYFOI+a+jQivVq6yme7LGSYb
s+GOiMGe2wg1VLxNmHJCZKL5VrDOkZXHKkIpqIaMxmu21U5W8+inLwQqoajHVNoa
UCIxt2PHZ2/Y4REJmVdEDe/jSFvBaY4Lm5Yy2sMzKPbSinHpEzivKLPJvrq1CvHy
Hv0deCpdKzcWlyMTfbRe258JBjOt/jl/4+ontbylwv5SnoXzVwv/c/fxgZPk1wBg
CcK5i7tECuOt1BuC2/OmocyzidfzeefOKiwN/xvjxk/i21gGFfgCKQp/2v24a/1o
SiHviFkZOJzT3dD8E9itwwJ8F5ucVsolgPWI2bVfw1GZuiiXVHD6CQwfmXzWuQJG
7/H0Lm8siYkl9vgR2dQ0stbVDmH9oMAi4NnNTRdS962HTaVRRVuAL0Uv+BzsYCwH
ceQWDVsBuhXMfNvQ+JhD89dRNrwZOuvgz4P5UVdTodKKA4kxObk3YGoRM8RLjyFY
U390lwFC5AHeyxP1vSKNpIVLRnt8IjKNVpSeKhMsuUeCcjSCCxne8gB6vS0mna7e
DK1GjTtDul9NRR95fhlYGLKQklySmiyvEi2qBw3TTsoEiEqshkoHqGIzimnqSHsK
ne4PUueVXctgW+mG3QEw7ko1GlNMNe+vkpO+tSJqs/5JKmus/B10XG25AjGAoR0B
qUMGLlfAzEdmZCL6n7MuL/8i2PpzDF7Ymy5c+fc7e7kMdN3pioX8I8csP76UlktM
TQJBWVXIgO2i4eaC82Abu04pihQxMs/3NMiB0yahg52gJlUEWFDLb3tBzzgA1Fuq
sO7H4nPOLdcGN7QJx5NKuLlHxIVy/EcpMht+8RnhxspKyQXOTuD4z1iM36wAomqJ
RvUbu7sxQbR+Y21mEPNDtIMIrNpAotjdAfUxjWA3hrqz5ym75j/rgPpoyI6QHn43
wEMSH2zOqqdVT+LhVVCzUrbNAgLE5r3+RHP0h45P/WOCG6KKmf5t059UTOHxDh+Z
ySviVcAb7h8NCaENRVKh4M/NXYH1Z9PNjIxdNhFbUXc3xc/mm1HX9PumNigWaQFA
Iq+6bR/7WJEcauRIcWo/FuLfUHfPaiKGtTMWUK0Anq9SamWmebi2iyraypQT7qBq
M/fgbgVFw7JziM2IKbpATNupuAyDsR4PSMZIDbVZyYfgIuAqGwmSjLRBtSmPuHxG
dCcPaMVbDFssm+/1iDCW0w3Z+NvwsJee1TPb/JfmoBJAmJCpLYRyRbEirY2Wh/z+
dzBnnIPzxRaE4xrI+WEHeBWXJyfw/9p72u1xKhz1sXLJwvLL1bDIzie6r+whCq5r
FFXLum1AqQ4sVg20P1D5k6zmdN8/hrjYubWoNFfs468sYoT+yi25K8kY/7MInpwH
fdej3F5wPt1quG+phqT7kQuUErAIyBj68FFnSh9Bf9LO2VSVgO5UwmBMMOTZHyGu
S2dTTlspsK2Kva9Q48lR02ZsGemVH2utFfnKkki6s54Pkq4TwoezdFlYcVwAmc0V
8BEcenHGAUD1CAFarYHQU68QeyVnjhe23QyW4YXdPM9qsxRS8HMtGoNj5Amti0Wo
IIm7KpwYt9LzRw/G3NqxFrj1SNgYYXSRlw8UyNfjWaWsyxUVdCDBkz2cOJ+Bkokh
kum1IVYUrDTexNgnXIWlDkLHbBrHqfHzfwaOpI3kEjWzV3XiFya2EOquBFcaV2g+
/pZa1m9Fy3M14bIpAVpL9tHNHVlwoT18JLECcNyEyUkAq8zgHtJSRT4pdMmW9RDX
Ar9lNI9cOXu4kpWwmWYpamHx/ojU107MRQkdmcNB5RmHpES7LmSk6IkSu5WI2b6q
UJ5lYzbI/1J8lk8YZ/nFcp/RHv0B2S8NTQZAFlZWbGI3RZQwx+S3gM/HUa4zeh0S
QLsr7Az3CJo2JwZEoq3hv1wjWvuco3uH3AWqGyPpC1/qrZlA3YzsVPeeVCQQhlt9
DxYdxD5rfqO3J7ieQKZivAzi0NDZorcWb9kCoEUW23zNgt2pYfg62pSfcZsV/Dgd
avKdhw66dKJ77SMTbZHYYmD5O1GoEeabU/z1PMgP2LAEKfrRqAcbVc7vxCpilZUL
VlFcY6PT2GkqmMZ+aBbXFd9zDqCGWofdgcikZ7N2fCsiEwG98CYd0n0p054iVVKE
08zVHVhlkTZzaoz8jyS1gbnectPhhkIHa7URv5mFdvHXOgBw2c8n7cGMZ3TZ5RWb
p7FuN71mwJqlqI0CYy/2zr5xdP4Sm6YP8RoZ5ZcoImtNUFd1PEQ1Mml9iBbzWdJv
QXFl/s4I+MwI57lSsJ4YJc0kmXgnAk3RFYcz1hKE0IyDhNt2gkwBAA7+O/HymdXx
bqg0sNVBZ0csYgR8+2kr1ZNqB5fHfymDnI1PwLhSodbzrcMC1jwrNTVnY76TPwF+
xYeMotrNKebtN0wcHIrcy1LSWhLYhu8qgSSDqjGN3vZK+IqpsUzaEJAxj7XJCcty
5a5sPgoVPuL7NzGLj4/HamTC4awJFNw9IB6ADIFKEuFUoU8AnvoLJKXVwl28HSme
BYE5N74IndJ7M05xSilaQQi4nlfM7sQ4gA81dkL0Rkp5hhL5TmD4ofUMklScyphf
mRJNmsrOi8rN54fYxxGpeEaQHieP4EPs8l6vRprtdxaz7n6hRhfXDAxBjgFwX609
v4jGnhJFomicMKKymFxqExcMi9OmdaVOHyUbV62WzbAzba/8IDlAp7wf5Vw9bsIp
NVukALBbXcngcJrKgblyY5iZt9WYhY3BxaUAYSiGTYByhDYF35SK8bE8gmTGeJQR
/t4nvqhk1tkz3RZLCNVnJiPRQvjsPhGqY+5tLoOy+d9n0hk17TuEAkp3DACJQ/ru
Vn2QvU3oOkCMb/1sckm/qGzLWCQqQytWPkO1jN4hmRSdaCD7ainAzuZcr4db2mGn
VRVPnk/DuzpHdjJwB/0gFoPUQXaApGIPU50ILq/6xItrd902tAhczkINBiENyWDL
XipSq1nnGm56kgDoKES8HSb/j9LPcj2jaAcjAMbXsPoLmrqkBgaNHTZGMU+IVSNB
bLfhz3Dwq8MAPcmxr+VtZ+HiboP8/ry6cqnhXaN0lpopfMY6Qz4lhTWvOFPX96dl
jcn1j8KEviM7xg3DaYd63uq6JlNB/6kVIuChxIYDH6UC5focgdGWX9XIW7UAwp/Z
XJiX3XkkfT7QSwBOckKctH83KMoSshOa+Ql1rhhv0OT7nhAZ+aiVjCXOJnINQRgG
aun+3vgmb38Eemd4PTmCGsLaNYEW9dUNWFXVSiyhM+DqzqjRXMwXNZNn0fKHp1I+
rc+DALdq2zk/0YL0cP/VaKQEgLiPryemlwhAilGMLbsll9k8pSNNHp7tZEOfYSDI
LtGqrzeXVQ0IoX7YgmFcfuI2SP+N+zAtnQVrE0nWIOSxL1Uq40Aczv/BwKJvu94v
xB0QFD5c2UDLizCHTRy3/hR74anB1l5I1DzrUHB/wyDSUJH12uZcN2FFW/22t3+F
ewH3LLP4r1M8HeU5NHOqJoujWQBOeiKBndN0CPSgsFq4NtWyDLBOmdOEYSK1hwmj
++QZggl00fN+yOvALJ7NUW0EozrqLMW6umJiGqhuoVwj7XjFOtNbKzaQGB/5kXUB
fKys/k3E0QymyO5LP8VUnClwCBFtMhcM6ieREMX1uy1Q8vpVUcy8m0kDenQpDMwf
rC3s2Vdm0mKz+C5vbQAxm1kdDTzsfiDPjbMP34S2TktetGljNAGg7VoqTKVMMGjy
FCTV1uTbiggdeMpVWA1H1PuJHdwmswJfXWjHwE93gVNDTHADdG/z5tAxoJBDY0qj
3V1Y1ky69g6hEW6UY+c8wrqVEJlKjui5PF7VVc2fFDlHA3gejlW0kAN0vCHlpHvt
+ac63pe2wkQkcwBQoAqnGUjL0ECAA5vlbrNaibLEz+Speuq3W5oMhpgHVoAgQIUE
fwg/Lk+LVGjgAucHqW4as5xBwXE/+12sePGqanUHpuXg+kJI/KoCrQ50GxqHjNHY
HzidI6wTQCAQnMI3emmDjZ/QPp73JjZwvyzbHVq36AfsH1aCDuvLTfvr4BZt/iRs
7VPIhvgZ+Up7t+7VIzLZvVEmVqJQuH5hfcfXM/Ue+eB5CyggDdiUnOPvHe2qcT92
ruxEs5mXhUlclYDK4dgfNr9/TX9qcChRTrToMsH1icfT6Nx8HsmWg6GAKS+wLu+M
8omTGvCB/ViAnaL6gM3aUfZ3Iu5O08sXK3tSWKtJdB1LzoBfp1fMdznjcz2LfBcW
RQMkntV2R3i7HkOWQDRPiXPJDEcuG395/ZCtamBMzTZDsJitWxoZOSrxj7ZN6+aw
7R8PC1IwJQSgpdAEyllWff2UyXO7lJWkNB6dg7YZbQ/Jy11Q2TdcVdlT4XtZNGG1
x8d/po2ShyctJq/3VSGdtjmrXtdxA4Fhv4xuOAULz8EEglUqZnpBabu15xXC0c9O
VAtcPMDYK+4Xl64kNGoQhTSnvOPNGgaRII66XD69few323m1XPvKJOi+xN0tiGxk
yi08FiZgzjQoZI1T3VmoWw6MWtW2hME8PZgVP3Ep+SowRtUjGusSHlL/MxD3m7+5
A3vcpVlAYSkA9I6xFsO3/VVTKBbD+/umMDr1I3gbh/MDxZr5mAJ+pfLsIvMpKZ/k
gBw7LN4v//fMgRFIsj7aYL+ecsZous0F8Nb3YbOQIwLlhp3sXhiLS5/TIxpcXY4i
Ie//EghzdEJnfcTuH9MVWezcxH8rsElKO/Rtt3nnkKCIqkAsYAcoqpW1TprA6bZ3
6s63OCG9E1bTfjab/R0HotsXNh4zPiXbhMPDvIs8M1BE7xUrbZcKBDgfhHfzMguM
2rpKMOFuLmjA/aso8JAjQenGximZmzJcacqBxbqflsEyow8g6b7/zrH2WcvQLwNx
83qBZ0XpQS4UPG9JrINTlVSDiJQQfb9aR8PnXJdbstmgkpSjjiJcOy74lNNUh8UL
msYqqOmywOKHlSuklcJaw5Drl0J7EnkrLeHxMSJspGeLQBnxnpXGjv/IC7RwECyC
WdrcWpjdz4yvMNMknpdurA2MYuYHp/R8SiCBUil/ZSANmH/Oym6kmfcBnt2xV3hl
tCcYLQ+3EQv3Hr9abG3utyU+qnOZZjGrfYgPtk/AiSlOaftUyOytvCXdpsYEwdn1
09CwGOJEVSbXPltSdg1TmJbNTSW9CGdla8fMpwpkCinJM2aRfY/DgPOLYowdj6Dm
KPS6HF373R8hFBY5sw/MhJJZdYScOkr2bO2nbi6jW5OzA/d8uT/BTOX8hRnGwDGa
XywamB+BgnGWJiyvyJu3XLscvhJN/t3WjXtmn+cfeVS5CvOzDuOctzsxyHI2y6HB
45E2FngsuBj4id4QJ5xJNeKO9UnKNXQBqnVMaiY6P/9kJaLEE88V6vvGKLeL74Xt
WJS0n15iHyy7rxJjsNtBWEBqxBqCgft8uf0/TmYpPNPLJNeHVI1KgmzXtdnei0Vj
7dTJxigD8Fb++1iO96VtvW5p94jDzK19IGtrLVQ19mQABRHOg4IkGW/0xJFbaSCO
i+8EM6RFav4G3G81tnRkJr7tG45WW8tfiCJyWdeAmg8DKVFdvc/ny7r12F9ue7oN
MVuSKg3dpmyB5WClIotW9u+Dv/vRolAByQVXCfr1jc+HyhbTcCl/2jSJoM2iP1Tz
fQM3IiwAJmI3nguM0jFa7j91k9WoiL2g+SCuHN18SGmk6pmIZGtPdR0aEflnFUdc
DdGxrklLSr49an082W5bdKSE4rB8gP7T8WQUCf2kmZIWx3MpiTe/DyaaVyzYSTf6
g7BhpS6SyYddAQAHBYForICQpRZVPjEw0qTbyoIczOfY9x4ZJt6+FDinEG8oQBwB
FMMDVyyNw6lQgEv7+W0tRBQSfdypn03LZTfaqbLFdS1TleWd5fzeUPcrapXG1d9e
DCDum4wTA5eOVbzCEbDzRip3f15FLrEAwZ77DUUAGZOEqZhSXixNNm/WcWdBPLw5
igg7n1tSutsKwYd2ZT+n1qguQgssQatkSHic37VSiIU0EIq/pLaFZRi81XyDcip0
dxI0W0/MCqV5+//se3c4Bc4aJDRoTV2BQC8eJ4W0MFLAK5CECeuRRhHgGWLqp96C
r03/q5geTcSIDxbPFwUmH50sRTdmltEGcKeXwqyQ8oQOZKIGdEx8w9nwIQpqwo/d
VYsLeN5fnM4apANHs2Vlbr4866IF6BIwpPfxOJ6II+OH5Ho8Asc9Oa8V+i0Q36Sq
MaJlypOO4RkH/JuK46bwpOBuCFsrsL9u4APJS+VpuGWQfWlTPuEEvMzss2Msha83
m/qGio9cdXxgBv1kJOrnhbdL0YWfXibWooTVTnMbciRT2/Or3WTvFTOJnef8ly8B
nrIO9A2D3Y2YQ/KoZXGWD7aSoz5lFjsCWcvwccCaW7lsPibFdNLh/ACA8MDSceJt
2UsTn3K/b6aQRUp4uLqEjQaZJLofuKn4ctSxLUk41u/p/Wp8s6ZKEmSWQvKuG5uX
9HnX5zc8wlnHv2Zzux/wFqM0HxdVQgwokQjyXam/h2hNjh1BzATJ4/d6wcBPEO6x
0UJwachliNWqo6ubbwnZS03bK3W2qJUsfve9p1f+k8NIxP2zw2rltenUX7OZSleW
L8AczkqhqcOI3/mP600nFAZWXi/RXWzYJPKzGhbSjoYyRk+gAWeicpegWH22x81s
X2VPQuCKyuJnWw3wngYYA24yiFvqE23sWuDbKpZlJxqJzTrQv6snRJHesHqoAZrn
pmFrXK4A5qxqaJlcSv7BWDwfHadqaWCxSRniZr9uMR271KsyKiogHVbopBMCVpEV
2LdL3nQDUMQ0DeXUoBLOVssGNa7YcKLPuVVSQ92XBrRIl6cvcg30C8HHSh23Phr7
VX6aYEFB0FObowWUCgaM8gZQ8i6xqHn5yHY1i7pZ27QJmRDhJskpiWNU5BubL0fa
q1myacycEmZJ69viPb/sG9iA1sLH7VcQexsGVdCWytjmD7Q9cbdZsNXTBUm2hjEr
0udj9bSN3ausRFbpA+su/wvDyR8vQxqH/b+SmX4plpPk6LJ14ummqx1YMV0FPNHI
gupPLty+xlJ79fxVKEYEzbRhE90DpbNM7+JmDdM79ZfkIfSz8jwFt0NlbHH4McO5
2zL/FCkQzQ3HdVyhFl5GP/4nwKky2HCeG0/cX5p7/7erJIMm88g4msuk+nMLBUPL
+8vAz4RoPg07EFqaMWpZecob+mTEy6cUrspdu3iEVDUxKeamyVHvnBOsbESEYt2H
Tzs9hPm7rL475y3V7dJJHNgHmk+aEqcHgSdpiqr33UvFVZJAk1I983CtZD3jWkum
8umh1LxbgtzciK9O8mEID9uMcK7DZt8j2GcSbkRxt86lOKFk/TBSdh135ounmsNL
68Ltnq9DphH9fGTzWF0FJfv0ADA1Z4psKLle9RjTlzxGYSHM+c5tAhmstZUey1ZK
C4HO/VAmn5MKNxtXzsa0gPk/dBWAaqUlrZrwo2w6H3u0XbNmRpRd1ObIIcAC74ZF
rV+EO0dbN0mCjRCe9HL81aElUuGaGKU0GxBr/iklsoUfrdO69CMNhVMJMKDEYboK
ltGi/1ytAuGZ5shPGcHsQk6MihwsBIG01IoHPqZhXf9Wni6jDmkrOXugnD3n9Jcy
+gPV1QEEt1Z6hzrNtNvL0hrx4cibhocnECPTUGy4P32su26YjilmcZfKRD7bKGGK
YjgGFGD2xP+rvItR8RmEdDVvhlCoXAcxb0myT2WYs+XFFQEQwI1trz+L2ZIxc+5m
U1U4ojc7g0eEPK0NRmp0mL9wbJ1Xq1fHkc/p1MgZUlAM94PJMj0XlHxUjIYt6AGU
mdpInhrlH05vmr0ydi5fqrUNvX2yHziXpyaZLAcjtvm5k2IuZRO1xIzitgmNSSZs
uPF5wvH51th+8AX8hyKtXMlTgGcKIvslIrZ0jq4yyWb110bQQBRufixrm2FaF6NM
dhYHntVe06CoI9kbZDeA+LZIqDypK8KY+4aXc7MTJWV/rn6OLN9Mbm8M294dQQ+v
FSQh2QsZvJ2yNoNq0PGdkw6GtcWh3fwBjWbBaRXrwI1ERX0ov11E8czDed7lm1Pk
87wZMYe1bqMWALbqYi0rjzL/gmCrLpaiEc599GlUUceQx51QvG0L8FrdwZ2Wn2wr
QYuBdeOATHHtDow0TLXVUK9ATSlyG2J+cl97HYGgl695v+BpE7pCJxxNV/unTsL7
268dvH1Jpeh0f8+dIm1cl0c5/tYkRjoyU340oWZXU4v9NZlg9ROTJVksRj8h0uNd
obIgFSv3sUm/wU3mVbyq7p0jAq1Xvx12ObDm8k0K205U1on5RJEmN6ejti6VM+pX
eeriCYh05GzTkekKUVggDDKWy157WeW4SJtZjRBePZvuRM2m8A2M+rIlaPfpF5wB
lCcoD8AwzVA0K5KCG7ix6WF2OiztyFfQISW9rDhPIF4ZMsJbqxJnzuE2kccy6yVs
8QGqf2M14qK71eTzGYIpzY13+UXbxG5eI8iqYSRk4I9nD21R5USo/RtQMNPTX05U
Se/vh6H7YMVMZ4JSjtq+EL6pbaOzfLG9Vfw5fvZMY18bNwUuikHfzjhDlgEPRptn
V2d56e4uSQ4lB4KfpvuvJZLKggxYrqh2Ik91sboedxuRhk90WFpc1jislX5fD/v2
c3AfjtJqFwd949IZvwWFtIKYUyo/DcUrT8pOBwwwg0LoSc1k5WZ66ETiB13QhY+R
6HMXMNm8dDoZV72yf2VAQq0GVSBm5Io3KTa4uTNVsn0lFbwoKFdkb7xVrOa5q+nI
xQgxLCAuDZrHKAgIfVAxOVo/nMLMlBOaWHQNkefRt8fV6XmsjcAWohKPbr5h/r6A
70cCzxBUp516b2xFTAfIo7kXLEognAdhEiOgbCalCebdh+piPfSL9c2iuz22tcIR
SwQd9aemwwfCOaXunySXg+1PWXpCzfXJNpPHa05c061ZlNo8+rcwVh2e5aGPW64N
auBZWXzqsZXatMYP/I9laLTDTH/z0bqPTXHAvvXqIwQhT+qIXrP9H7mzk4g1cOhr
IaLsp690H910a/qbPlUNxH9Y65ksBQeCeO6Rn4SMpnrTiVYg7szQkrq1jCWLASMI
tX3IH4tAka6jpPiJ6hZdxskqkW38hKwy+hhafuIgZ2RvnOUZWLgLFxA1v3NCRBPp
56VXJx4XAbpJj9drvbPhQPAhmiWbsDM/66r9vDI96n9ODpYIVo2YWlG3K3uXjg3J
h4vAX46XpQvl16yktBtvpbsvM5/CGvOUi323TdaMmM5vWSYZjWbJq56Lu9t2A0jf
RZrEuKx7DdUn9Rh4r8ZR/M/NcJzRzLcTS7VU6sTdkTZzlA4CMWFU3DEhkALqVW2/
RVjpQwQQ0r/y2ZQUp0IU4sIhKdE29wt55V95qyUMo8zKf+aryZRZpmqBNSy0eCRq
LHGrUk9Y9bfYi0G35lPLpCQoaJDFT2i3yzObXf5ZmtLKySut6w1KVy60cIknMkSY
jDbEx7jRp4w3HGLJFMbBgiwfB505hfIdaLimD1mj6nSWHdrpzxqAhkyL9FopD5ty
xccDh74pVNJyBpq/4TxqQ3HYmfQIaWxZEZv6MWo9yQBBmjb67wg3W4HCwmOXvUQ8
eijohdQbO38q2ehrKNEa3mYH66tPD6a3sRQzeUOQwuRMH9nninmwbnu41LZ2LipP
l+9i6Z3aZilgcvNJBbSzPMW2Gvv/rxjnRQ7wDmRqGWZsDagNZACf3SEhbcMUTzkq
RnIocrd5pFyF0OBh/HBWDAxS+FcF4ScZCZY2BR5TL9yPfofY8m/S+4ypPFZ1LJXG
CpHUQxYEbRyntOIyQAdIgp+M43pO0c6+wvznvNPQmPuwN9piDU9QjFdUCsvq6qBR
BN8Rw7Mwwp/4NJCUqR0QebIM9wM3oc0AgFPQifdwD6Ic2ruAz23MLQq3jv/5c9R/
9owcXwT/uVuwwxL6ilIX/rvK5W+WGT1JcKTkWBjIaUU8eL9iyXHMVtwkX2jQykFk
Yv1O9zWvoH8SvlNe1+73ZhhFT58u7+bzIi+67k00+3Em2h3siDCzRjE8LIS4VDQL
YXYtHv8AwGscE9kWW//QNKGMraC20KaK/JPcnEsXk297yWVRM7v0zC+zPsxY3Yb2
oJI9pWBkGK9Cz0DOlXQfsO01ztOBxVWPGHnzLmCSi6KvWWzJtD5w0Te1BuHGGlIe
YOAZT/auG41IGSxB/XBeRMwIlCeGuocUU8LaRJpTIKRYJgcLsVxUmVDAWL6C+zxU
JoW6i6wwZi5XrCpDbfVotGK+OtjiL9LPkWRYp8yXOEZm8u+k9Xc//RrhvDhfo2FC
g9o/yHCIa7ZTA7yb1wIe40LKUrb7/O2WyRaYw/1glLzos3pGm3jYrbyX2Yt0WR44
EKeG4U9QTWnD+bm68NndLwEZxy57EpFFO6n5KCmFOATm00PBc5VVi9xIvOYwsDeG
pCPsjXeNmT98AoGUp9qb4eMe+lbHhgACHUSFtY8j2kHAuy0PyUgzKykxakMqO4HA
tCNZGuj9p1dcubh1c8jtut+l8Sf71CEbBG1KomM5suBiCiengAvi1ncjXc2RkSDr
QpeKDy5Fy/Vqn7tmpneZNo9FsMLhUqGzRNaqSe9w6VxxZG2JmzX+viWB2PtJGbOS
6yFz374kTB+X/ZAEOi6dfM9fSsZAE6ZwIiRfYv3/h2LwdFVB5oiM8Zd+st1BLzkY
/a0Dyxdzuv918Lay6X/rBUJW42kY5f1lrlIsnl7z9KDCQyTnF7R4+dhFMBKpikjE
nWC5hcS8GkYkosLTcF8X5nnxCV3Fbyk/pyG78j/hPMgSwQPV3k/7GzbgmqzO9n8h
Q4QssZon/bHPT82/v/xsZv/ArARF3WYiroXByUwLDhW+gdhj2QKq+pDOSpm1CxDw
XIpWg1sDY5SIXE2aS4A9Lb9JclrQJiby6iNIiD+qBoU9t8slpPkIwmbElyqHZ8GB
hTeAgUwbKKjKtuK8vrDlnuGKyiwp6Fqx0UKQ9gljWXcjfhTgGeu1u/xj+xhqmNBn
qc2rV9R5elEfLHHZAMAI+98k7GvEmrZl9QMtaj1N+PhmgrEDHW37f6kE/hDshEeW
4o7y41KX9eaM+jY1od3cX6D5uwpI9OVlC8GwnLZgllIiRWlMhlJw4D8Bd6rMDTQk
m5K775hcKgM9slJeWHTtk/JjQrK6WryAPxVjKpoN1wBpPojAFjlecrogVspFdxRD
GO/5//kyV1KZ9/NFQ8rU7zDVEDUcn6tHHEKCKWjxJEUDpRQkeAre9g8ydXiTHMXd
16EnBZ3W3E/LbqkZjfnxL0wkA4j+y++3EGavsuUVwysFwuVSrZLQ7ILlpWQ/2pUf
IPCsaJGwUz9+iDrR9uKEmYMVjuZMWM1yGQf2l558eS5DXl7Gh/UC/QEKkRy8yscS
XQ6IbqOcqIHMLYC0QxUvHwCixUnOI8SJt1qTTvUeDi19/FFF/HC5mXqTqPWXumJ+
ZExZvUuL3hcqwweMt4xZ0cpB4ponxgQHqXwADPWJMRKlULXdSXEmeEZ5rIuNsOh6
pxaU79c9Zlr7JWtjnaBqYznlGO4O8HvLXQZkwJPxQX33mNvdX9R3yZhzMXcqyB89
E2G5zzps7/IwGU9WRP+UwCjxfxM02IkGxDNLr/LoSRRenBAybOVVYqgn68++n869
e+YrIQA7eEjRN3RCWEtafQHjU+wba2PYm9+PAXpiWs4pvkKKIe3xDAtBCB4Ww9l4
gir4xrxCxzafIX4+7e+l5RHCSPvfMGzIIE+w19xQ2hWhvLxFntC0g+t7qm3pk4gG
wpwXjZh/1MTo7nTkEiFu4qfF0ZBCAYHFQuD6P9nzgrqQZB9RFSbe39NGfuJuMlOy
YEdrDbGM2nnKJnVR1QeJ3MAKpKWLAcIfW0CtMGpGj80iMa89C28ieewRFrrwiyTk
DHdP63izfLo0dlpsILv8iZcK9Q8/mvZb81/Av8UyRDBSS7YyNfVafDVYcaxeumcW
+xJGpc3uWogW+iZ3BHq1Svf5QXIiaxS3E0mq3hidNfIukKbM1xa2hj9vA6+jto79
zywUyhFOnJdL/MPndYD1iwqnEIl+C1PN5p/Yx34ncPbN8ezC5zF/FnCCCECn/MPm
qm+mhcy0Y6tjI1HyBZJ5sv9tWJ/mXEr+E/6edAlFYoUWrEpIoW0onoMOVgb1gE32
kL2BSs2xVMgfChRssvpvU5vDdivSqTEOG8Ms/SOXfPrf0oFlVkL4tSFH0m5UXNFh
2ysL8VE190o1M3/5+x99CsP0cWXZ9EjLFxrRzCgiIj1Nct0dV1gOJTGeDOF2vvg0
kRHjNa8c76s0DEvf4idRgTSLq+4NaMgoCsRS1M/crF3B92myFEVMCy9pikABZZSL
B8pXznKPjFfyP4RHxIonoorm7f46/yN4Jlz8OeqnG98SiO03fW8652d7DQWZgPTg
C2P1aAO1VDl/sIEp8XepAsxpK9R+2647iuSdK4txP2aNfHEk99jnAuglT83F2/q9
JgutyJ4rxmsws5rybSQ0I6aHjVZI4mNx9wG6sWtLPCUrdCjs9STbc0rj395tCz9i
v1d6jNwOWK3CWdZL8Wz8qAEWmDC/CHz3EZuJDMKlTFkfgban+nayHpv3GFF1lvN6
NHTyrzyI4tyLyZijAcXVfAtssS3995r7Dk6QtnFK0IOKddEUML3oYTTwJets9kY1
+a/mITXSNkQtaJwHmn2QmWrP9Izlo4wXydgIwkeOElhf6Yg1PPyoLOeaVBHXeopc
VYc44NOK8PAoogAQ2JtblyMvNco0ucHhwcSMM7bDS6JJ2r+15dl+FjnHlJL+Eut8
ey2/yWszR3lcfsrvpwqo/zKdGs81H38iVhxse9apEBx5KO1rY0nbaP5XDjK+xO8P
hJftNsoAJSUyjd/auRhjd5A8rpY8U6D8Mbmq5C+28mCQ+6IFapEDYWF8qkYNdJBf
m8lXy3eC45SSosoDSyoJLg8kuYXJzPgwUzocRxewbgeRfosRpvmdHXuoWzdwyLju
3aBY8r/wt0aJm32F/ByimnvY53iMtSf8mXDGDxJ+u/CkBhoUWlO4mwaM/z2VZjPu
AA1w8TyCZeNnndEfniqUs/pXC6kDHfsWoRISaYKm6utuNlIEH13iRIm0+m7RMEpB
6XId+REkg7Aw7AysH/uS79N+iTgEdww79BU0VTbbbrN0c667dUsvPlNeF4GM3ke+
lt2U0w7jMBTiM/W3QTBc86ymbtITf8ZWLHlCvQiHrbgGbVlyY2E55zGYgfFyUu0N
FXtX0Msp21yUNL6REXqpHfCfGuNTvnWz4FtdKd1PIzbL2/QbETAZvXl5UfC8Xj+o
e7GmFfiOzC3/9JjmOmFK4I8ftpW7Wel4BdkpvWNq/K6ExVHNYHEW6/BV5l4CwuPD
ZxBJlyQgvqKQhzVSw6Eans53h451K+2o4AQ5yNhaZ4izKutmnXrMj/+DjghLpbqy
aSmuc5IoM63UoDdHifilraGw1xWhlJik2gmLks0WUavbozzWm0NHraV4yMCbvwUq
37SpNo8bngh4sa4wc8k7RxKILRnZqZ6x2S+X+nSYTu7Mk5u38i2DvWxVRKwYJAa1
iQNrYA/617+pxI8O1qU0ex95yobzwnd2P1B0cF7llI0/Ujw6HykoXlysG0dIz8QY
Guc5GGZ4BF0HD+robLUcLrS/VkxeWRTKsAooxgamA6tukhv7V0Ix4b/IeKIc00u6
fFMJGk6eL+gE5KegDUFAeFtYv+LdI33TkD09RV/8ya8B/Ayh18QYiundpLcdc+d6
nsO/pI+8MpRmzhc4nGqfkErDBX8btidTdNlDDpw/aYnOY3AvGbxItPvTcg6WARId
ywIAmML25XkwE2aQPt1nbpEYo7VOXRSRiq7HQMcBLktgQEi7V3vpxB0E3YIKA+Ig
j46kjbpbI7t/96fphHCvMtFVN/8FbQeTCDaYTV1ayKREUnYueJ/WXSvvmaq0GJJq
CRLYhnepoiuD9LWEtTVB8XaA7UruTjrfD3DNvZDo97KBrTdghgtEzUxpHndfJVkX
wBD02Ne65d6WVJrqI4SKSclN6GfiBN4alPs1rwHR0mf85iXEUaC+9qaOci8kBesN
a+b+yK2TvcH8LYhsKI7i7BVFlI9wrKBeYnh4Xt4r6zdRS8b4MJ9JiS4Y3opatxWp
+8908FbykwQWt3d7GTsiFOlzHXQISjzYhOP9WSZFiL7jOwHIi+dyWrJRjyRwZYN8
1Zgi2gO9VmI/IWKco3qzkTCHtBjN5mZjsyd6Zijtaa5Xv5/aXoXsw9rw+LoaRc+j
NIHahc/hzIibDKoUa5x/QPTOi3R4C3X7J4fWloFJ8PQlKBTe8pKaB8AsZGYWhOrR
8Bjk7i7+Me12jGFzC8ZpJyN+ct46tI58qrgEixX1WxZf1Gd21ze/ElDt54z2MeD6
zDkdQ/up/NzQBEUr4keH/DBgm2XQi3+L40HFgOpeQMKOnhtCj8SLQvx62cB9OUP/
+LgkkBhFds2AwR8cdTVerSPjGKQ6ZlWFbEindNDuovRl8y0Q+9sYeVje6YCbRaDN
xBqMVcNp7yC5fJzXkgTnNHr2D16UfUb8EGgxsPbfQv3oPYUdabvryCVA+GJRWCzH
UeN5zvqhRX1IDAWs7eKVRF66KUhgENyT+bKuY1wJWaKGy+neNKhy6Fwwekwn5VW2
Nm9kf1gwRJ7KAQRbFoVAsGcOozV7hruTo39khO60jImmH8atbnaKgMN1YXOIl+PD
y4Gg7y/cYhhNxtWQQC5/TVZE3E/uWOIMa0Ss8t2eJSEjVR2rvVuMDtw7Dtysdz1/
N/sLYUVPNLvFeXjo6Y+jtkiQroL7r7m25qMDgblqx+KYo+fBTXSrf4llBWOFQ0AH
+WokKkzb9N+Ik70nTnSx5fXL5RV6Z6bgN4ZmJWsAQp/VGYjxJvrfTznjKs7brw/l
3HWcP+aNyIe50koKz2UvU1AQrbi7GgRwFVZsH6LZftNrj50VFY9C3JAcoxVz5tym
WZSuql1PtjOOMMNdX+WjPCq0oyfCrS4IOqx9e2gffNIfMWOslJhUl3uvVoXM4txN
/M8qCQy7Ypsx265cCF6bh+WP49YjLInHGYAUK3yKiBp4y3Jg3LZgbkUajwoRa6ST
KHEob7VkUkkh4HENw7BkQf3Z8S8vCBKS/dQw3Z7IfZSH9NppNL64p472xqHe331B
ZcTbAqZBfCoY3mdsI7hG5EI6f4KnyYBxX4b96Oj2MK+Q3pIAyfdwXH6lO9GzmbB4
zkb7IugceYp1tC1va6HZmhvu+l9Zh/R/DKTotAFdWNgjf0TdNflBMy8b/DVdYvM1
rtuz6LJzLfFf4cX21hpcFUl9GKyNoClqwky1oGFPNtkN2ARyVl1IRKl7lWF7ArC8
o+mLDRKzqEOb6zAdGn+mIGhllXDp+wF8FcHbWOcQTeyySviX/QQVo4qi5HJb0ACk
96vq8zxq9KcOPCZKOKGgD3dZrrmLup34OlZoL3uJjL0JsHv+N9zfqF+OllU3jFyx
s/2eua5EajE9feFCK6bPmKuk0IFR3abVhFuapZuJbjc3UlCxtr3Oh6Sek2eU/PtA
9GYpuui9h1efQMeIzD90yrka2GBbTY9CR4VtGwSuYXs5N88RPFTnU0P+wHYp+EJR
vz1I8pnQi+H3NvFUCBdW/L0WIfTSNZxnXWtAyMnW666WAF4ufZKgU+MLyEqWdmXf
UHUYi8FZ+igtyxAJkbYpcJ/tHvnv3SjOAgbBkhDauXiDCyZ0V5G5pMFHG0x1MeC+
efBxbfyF2NWdfzvZJyyb68RVL1a/KRQ3OSyF04gkxmDli62LgKQapCmt4nowE9t4
sA6sxfNARM3NXDXNRyKkMRZy6GeJnpy20K5xokpQMIGbZ7kR+xshFo9FtZ04GWva
hBVLVPKA1wPfM2mJtisjreuk9xdrfS7KN5tPmP/dquxdAgwLXXN40ys53+3uMNKp
tiQbise/+BN6QFWRxDLIs81JcfdZ+kEISJHRIPjSM3CtppET+hrTymKKasX2zSuX
CinghrOoQJk0/oVdzqerUsQ+EdhiZiLdbYKm+DmkGV2CT5tMjGBaGJkZ86IJur5S
AwgqtD+IFmiwd9ToRw/E3HHbeXR5pysgWON2cfhGwTW4nS/7atSeSsisY4vWHDq/
3pL4N1iyivw/hllThqCM4fmx6KpfXQXzGxiiJ2giSfmxOYh4Cy1ixHnK3SAkbVAw
rRozvCIcnP75pymvur7fHXqkN70qokuWhSrIdNwjv/3s3kBV027S3b9YMybXAo1m
JCvUw4xomCajeal7/tt+7L4b/4+KFn3yUNmHzs3rBNySxZUg0JT47ZaQ41jclDL/
eMwNgykTBZs2o4wb2/KXTdm09t77IcTP7ABJi7rrPJT9UoTgc/KrKdkWMKR4hdbk
mOMbh2cGET9iKj8fgp2e7NV5qo+lvU1IS073LnTlKYPvOSRrQCgoJXV3x7EtnJ/w
E2f4BJO7dRPr0VBHsRGmaQ7j3zFxiGswspJMmrZOhcfdfkwkCkmOd2y80MNyXZYj
c3T0yzY1UejFfXE0/33OGxkfgti/GAW5iEEyh1SGqvojdIEUenn4s4ir/n3aIp3Z
vVIg5ss8tYoiVNHu6eyfbez3bs+FbNQhLPBWUmIfRiRpqPnVikmwssMxmoP2WXqV
TqIS7kKUo1/H3kdG7n8t7Zw31SYyd6PW40ciOInvbJjfbILC/5hnshtusswKWn49
QC0YneZ708f3UbzftV3S0+0aQLhqyG7I6LD0B5STItfbeQENVlwHisQD/2JFXmBv
urcsP27s2UWd6uVep1A74C2xH3i9YmynT4naoHbmR5RU8wTMJEKorwG4v8u5ZjJX
ToVnKDf70TMsAjqfteQlBG9CajpAjzXnXmgKr3ySzMKSdaTwdnj75IroTKyY7H1J
zYb3uv1qvyy16NGnd5aRUn5WDt0ItIyiBzwvqqFwtOVebwCdpXxSiy3qS/KVwABo
H/8m2Re+b3yEi4MzBP3VRFJ9qcNLm1i9m65MkZmlnR0g7m+sdaci1pSs/qC5jtrC
GQw+TwvrN7sc5ErUf/gh1BRSOKI3EOi9oKO6vqK6I6rc+HeftEmWdUciOH/I3rj3
w15UU2+c1I3Cq6J63TgdClgWgjWPfmAFQRuX3S6DheP/6Wh1SQZn+KxaIjoflW/x
55I6RNI4J3DcWnavi0Dm1G/4BAAmQj+OrKbP6V0CCzCCNt+6GhJkX23x88AxWaWr
o9a2c+utlZQ2cNVbdkxjABxliCAOxQ7jL4gZUlosWkeWZ8r56QYD9J+iik6LFvwY
AMzVrALymGJK9938wBlrqM+B1+vtR8gtyC+7n5oAFJpGXdPJZeJgdngNiZEV2rIh
GExcCWKvE+HpHzN+1z6FxPPZpY0kTAtME+1qsYfPu3N4t1OGV0ALrNAogp+Qm1YO
d4Jr7ZehaLC3RSmYnGjJFV/kw46Xq29vDySngz0b10j8RdDnqFBKyOmw6p+GdwfO
Y7HzfzzgiRthE4oosDQdhqaO+R1e9hJ6HHhzCSP/+5k3rguTsz9G5GEKqI9DxyHQ
BCoevi1l4H7lD0gt2UGlQ4i99nQy5I4R8hhtvmqMofqhbaDxdUapF7FoxMNPLGnP
dVChhGrnWi694kBBKubQd0TGemZPzP0KT/W031xbg+Z9dQuC4StgVxjfaxewBlTb
5xvBu60lAX51sO/G4gxJn3f8WUBFX4tet8a2V9+efpPrkZwjrpfzFeCUjdyNV/SA
UsMRZNPvNPlMrnu5lfFzcI85ZSJzuBKiidWAAaacxhjNCnI6MdPF12cFUwjanq8F
DZbWB8LAcarPcoYiR4Mr4EC2oJ0YlCdVef/bCDVKdXlVobc96V9pQp9MjA5aFrTy
i+kgKVjGjYkEZdkYxMqZMSr5JnonOtcWNlwc0u8kmAZ7wC+hTegxq7HukWSFUE2C
8hnupKaAPUBf1YB1Vw4AiZKiN/5Zbochxgg4DZs06bM4BXO/QoHZQgGo0krULPWV
lrVDAHRJnc803+N7jFSvzQ6zVUzVlnw+Vxiy7Ht54dSxfY2gbWXurs8gpY+cHXcV
AwUU0F5JstjtbmlcxqTmgo7tEPPIcqbIJjlBwVMe5OzLw+cpJXwOCdJQ5Sb5GN6s
t5Tw0LTHq5l0LNQarXOWPigxJcYhs8Zj9J7IoFdmEWuGJt1CxIzSvk9lRcoSSC0v
+r0EbJPbEFX8L//4IkN+27bUAXLoR0HJgk60az519rRh6zgm3fEEYuq+6/QLrEqC
TQwWHiLQVjLjceCbVRsNwFTZP5M++t680ulEh4FZQ61+9zF9CUiT7OBAApDxQnXm
iB4DOIxSGD3Cy7E3KaChZIjwiqOVxWJL3XRr6dyMbpkgdY4P4uTZbXRruNrYmYcq
UcGZr2m8xvZWIR0+LvLD/kPxhf6rMLc9ch2DT3ryL9b+aWAuVcljy3E207qfOsjm
OyoichYTo6T97Itor7/Zth9O08HYdK1894JRAKmTL07IdB2PafMxtL7wrdOyHDnM
dywLNLnDra09AHjwa6BiXIQs5TTUGMO3ZS1s31OwRegJ+2Mn37LHgiKXbmdIDBxE
mYm3neEGM9oKGS618xFi6USkR+PMYMZlwYjZ8MLxOkl/ec/7TfmpO4G7379saosn
gLxvbe9MYBnnJP7aGqpBtixyZcqFzoNCQ6rV657KV9RlOQQSMCSv/9w6SqcKUpiO
m7nFfXSqsGZvaLaRs+Qd9ux4zwfvl2d+QeiivtkAQUPWi536Tf+8tScP5S3CnX2H
xmVvGlYGOcYnSSS3M42g2TTrPDcEDqa3VT4wusTI4XUuBw1Rf1E2MYb20y632QNj
PQpHIhH7MFoPad1cR/Lxl95tADuj1cVXUc7pPdBpsqbdr+AsXqfjoNX9vsx8V8Yw
Wdt+3WxB9Q9hjMHiuMIs8WV7pUYhl0hbv3kx7PLoFU/eFIVkzjs6pXFnQV4Tv/BL
jf/Ad/znsXexN8Req7zNo9eM/hxGbLGSF6uf+A+0y60EE4CYVzKGR3MYCl/ZWm6m
A0a00gXWOxK+MW8ELUFG1EzU6oicp+WTReLGW2bGkxba8qia1tl7DpLl16KmvT7z
T0m0uEJh8qQ+YYTdePN2OYKmSr+zyhl/2uh/40vrApAXpquCrfOkdiCKJ7mPprEt
v3PKvMyHeCgOtiL5L1wKDDUmwpD9WBIJlNkihOodtxvt6pJ2y0bGzagrhKuR3Mwa
gyGSqdzBcCWTxYq/AcW5vvihcEB77bGFBGrDnD+wRLPpKvHhC7VSguhLEUxMkSpW
zPHwmtFoG3Yum1SH55Fil1bIgAXVDOilR+YULTFsFIiQcITWJev5+42yRmxJv9dc
WfedWPqvjoPo2GbyvG3iukgaIgkzEUQ7zKbPx5Y5xjPNyhc4+TZN1SSwCwJeAVCa
MST0gu5Hwmz13XuGI/Mek0DZwm/9W34YVS5ha2N17LqHRkfw+PSyr+GdS2lkdCvW
ol0NSCK7GdLnanaho9LW3fshQIhmLtiMlsDDMXA5X5/UWpUhFeoFOSzfauQq8Ugu
v+oinJ+pobX47akt1LGjb80v6hJhgdpf66uj0TvQ5gu67nwmSFEBp6DZ3YyxvCR4
Br09C19/wDTJmS/SisYD1KL9SYLqe9piHYm5/6/AurLWXurdt06nxZ7pEtMZQ6d3
OqybZpb6k6CgYhFUpUjuVhrRXS2mNaVbWwQUGXnmWncH2BfuYtZTjYzjl7VOprGC
utHf7B4xZSorR0JvrOO5K4tCA9kU3C0re5r+n2/z8CPe/WWmIQTtbpf3uJqIHWKC
zxUqQB7F1R4ADiFKhx+6N2yyc/uqLeqpGlmW0Ns7parEY7K0bdvY0L3lEqkFo9Nq
7W44jbemN+Rs1A77C5e39ojLul3osEHCYV7qsYKRmYQd84hLJCG2DFYBIbPBjRzC
VpwcdsuSyX5EmMQxrveyJ/R6FHR+d7GAgutXlriEmALgJ0XvagXEH12B0+2CTXGa
1JCM4TSflB6YFJJlrUS5xHW9Je/Z/RD3EU2bJ/0KFyH18xHtlsun/MhdjvTCxBSG
uTtmINKKIK7EV7whzJfixAvs95xb9XO01v5MZdQV4HBxVZyfCCQrQQ0hIaDXHAYp
DP1wu68Q1sAnA1iFx859RTu9h1WkArSCkH8wB29qixHmJmLCMrV/c41D5++lCS6G
dKELq/7d19YxQePCqcRRUjcVqXlmc925NyXeshoPfYzg5tVnokfv4Klfj0MUwheI
ZA4y5n2rfFt2RsA5sugAFrp45yFI8uNFu1U1zSeY9VN/IDx10XzXmSu1GCDK17cp
LtwDgixWXtDA6NIVXIR5bVP9qFMFk1+VabS/qwaLSsBlAt2naJP76bV+cXcYfzvr
pAOtarXk42+9U0POLObPSKQ1/Wf7/uAgWo3ytpalJUjNnQcZdACsof+Hau9qFTa9
iOWLnaWJTWFf/palxc4Mr4+Qo95eUPfZCyxDyGJEFv5fc+IxMUdPbxq/VLXyqaCG
lIcBDekjhxWXucP/ldfRYvfI59h1bPwJCMYvsuZe6AEIkGBXzgtiikCz6EE5kght
vxKWflUeiNd+haL1+Gc66RI7kN8jpEeU97TfkT/SQ3z2sDTrYqx6UXeqcrrwZ2Hu
oFw3jHjTUBdfc6JXhX14CpRxwNtGwb/e1Lflalt9o9cLD6FBLBzGaYgG54+5ZROZ
Ij8kYMJ/kh/0+WCl02mgpKjhUEQuAS4elLjKS2e0xbG3/2L8s0yuIk/k9Y37U0h2
QU/ENHdfXpOUFuJqBplNfHGrBq7n25HrPzplzpQ17fWBPDjGaNETSB9VOIQTH6jq
7tHjWil6okpM2S925ADajOlhvcMCIij96tyhHNDr7Hm3m8AzMfYYcTwdmv7dHCmR
RGBiQQcdh4L25K4UnRTl/4zArSMApoz3Ezy0IjTjSkqsQ8BiFGC14d9+70NfgGqd
gYM2Fw1dUlAh3DyMxpnXtvu6jEqim2Au2sdUn5G5GIUx4Ooj2i0X6kA37u7VdWCZ
rz+zT8nT9pZKREHd+lFOZGeFZa2CtJOApMy6z7k3TJWBHzmhvfscqnciX05AzAEX
tdWrNxqsffCOuzQOfWCzUpRvJpKqBU2qyknIApZ5cUQFsuFA9Q3rKG010VnWazH/
NAj0Bn+HoDU14gHhlhi3Xp4NR8YjqV1Gqon/ad55UXf/FuA4qmWCo+mkCk3K4jmc
wpkbkYPTggxg61teBB553/5FEqBwK7xWQe04H3eZ9eyofFKUB0NoXnT1CNRmAWfH
ZzhWZwGFGfONyuY5fNg1QZFwgCCJkJHGpMjblQFBsdDN4MUR+9akd6xck9FEzcUh
SOn+rbKXA5ujozRttJw5ouo9piPyL1376HX5xZamL+p5vPZp5ILalAtliKODWvYO
YTdJaxJ30eWGvxagC5S5OHeU4Flx9E6CouqYoHgurlAourmYr9kgEsmxb6BO5ZHG
AioTXYaDIP8nwOsyv79YwwiVv5egq/Vwup+l2WGluM9VXz1BQWYfw0KLJdHDP6M/
bgK51FFHrC39UTPPYucpVKqpDSG174Oa41T+3BGyBqjnqqPuwap1YRkYa84ZuXEO
3M2b/yn5qCiyQTv8RL55KfrwDxcP6qtZhY58xn4Nrv/l41vQcEDQGli0xZ3m+jj4
+QX0VW7pjU35fwqtSmyqebEX0Ayi0HbEeSXMyE9bQXWFKvv25vT6Gk+5SZUmiHyq
GUe4Wd8FWAzTbktMhFmaVw9xe7tiZVGltBwJpsI2KWHm2iU5/ij/xXgw2+NVczPc
SdmOSzchiAsLI+tTjOGJkpVVGvEi/NzTpW/KdJd4uE5m165u2xr0PFqh0qdGStce
A4/7V8mDZRcjyNUo83t9prh9mdu8a8kagRZHHH9wppAdzaieVo8sCnTt5YCz0OON
AKsZZVK4c2BKA1aDdPMZ9qePdfjgngONy/cU9qwTVMosVv3c9L8mwOzTgiRZzgxs
H1EjZjIUnL0aVyyE01qjtIV6PXPk4oS5/Ajuz337QK8Xe7Bc4A+iOzxtRdvN8Wz/
C6dWTtk0NKl2YIhAlo1993ZCK+/Rqq806JTBVJkfSEqm4uhLI2rDTN+4LRUJU/L8
zcszJLJ/XSSIsLanvgjVBRyOo/vTLEqzVApkt1TJisqUF2vjsshsFukeWggLk2Bi
Eq8M1feQAE48TDLNDENi/4UlvZ9qp7Z1HU/feZZLhMRLZFtx+pQvcbhKtthk80su
sJub5ZTBYNXe1S7qT1Eh43xO9L4r2GwYhqlrlvfblbuI5ojQ/KvW6y9EzQs01j9V
4KEDTGuyi8RLoACH+JLPnwjnLRZwJliWZLGhqLfx8S7zqwmxpTqiHOWyEky8/gO0
qeCa7DjdUw9ZyAh0/oESIOabTLyng6Dj/0pVmI1t+xkJUHjfBu1JNEz8HTN+4Gj4
/U05RHFGBtPXGV6EpbVQE+u1mnSDeKkd8KN14ackSbaHyTgCUbkHJpx8J/A/ulDU
Qe3jUcnv6NJ7eDMkPcmuDInwrBxP5H5HxpOTeu5goZFsE3G/xhxvJ9eLmS5eWue/
aHqX6z1kR8IwVNZoVrpgiLx6SPgx4QcaV8Tj9yemZVRKKIwJpo/KvoeEYsUhw5Kq
VLX4mtRmCFOmHCBZ3fhv93rgqqQIxprXi/5IC6Vjnmttva1hPchVWnA44ZXOlkn1
OUkijTGlobtHlEFyrpD6GG0lDC0Fz7t5VN8fHuCRbUVcVnWMbKKIfzyUlz7QTmeE
BrXO+3RynQbZHeWsz3O+9sSlvOUPp/VcaWvvph6S84CR25rtkHrkLnm4gPLdntZS
3xtG5o3h0XeGDLvWr9DWqINPAmYldj8AGcaoRd71oIYVSfe/35+HiYf3vni+PSFj
Y1wLUtHxpf5ufhPvt6y8E+pjt/bCy3MAxMY7AtvNhiPROpgSB6SI4NdeYTlI6KIP
HYEhY3sZNSYIr1VBVUZOJnQ+r9g9OxIe79AUbCe9AzZQyYzRxs7HUTtEyma8VaDt
FEgwlr5Jy00yTCSzCsgBmt2Tr3QqdunhLKiihufh6cPQMTJl1nkC5s/NEYYGOH4j
Y2SZylrqAS8zu0U2FCRxxoTYnWOSYVyxQzPiweEzMFhwigbHkZZavW/SEFX5rkvR
ZCDHJQVprre2Cj52Zm6dyS/OCYXBuI+gwOiihuuWlZf8kvBWl/Js7QxWq2C0gkuY
RSo31uxu8CeV9sV264TxNH1jaBQ1jk8OXtNs3Q2t4GE1ZC5+vFmcTX/1+HlU29c3
eNrN9ltUOJ5yp7x4AzXhc8UGCpxpQ0yI3/k7CN6CRkuFcRNunsQoZri69q9KuUZy
rUzVgeKveQecFFP9YaRLGjybeSsCeLDP8KXfFcoFcHddlj7GuQjK7+3VXjxyzhun
P1JwnnVOfQeAAuQRL5JY8bA8ij7LnZrb/c6tbAr0opxjnNHp2DjM9ooGBNk9ZyIQ
NODC01hbLi+UeJFxS/MgPC0McFfHW5BhAs2YtphjsCTFDbtV2pCu2b/uauwUw3yl
aFoVlaO0VbT/I8F9Bt/l8mMs9MpqEYy4bRfLINs4C1/IzhuKVLk+aPmlnlt6zeWx
OAx8B22m9GfGbaH13TCZmaxA11+cBKacVRTXtQJjdrvlFByhadzX/7BfoonpE411
eVcZqRvMVa19bvB1no+nxPzyCVD5VJIpOMdBWGmwryrapzOGqFwqt1Ipxe912x1R
VN0qjp7XGF8eN8hYmkcMmTiCClZHCADXpe6Wj14TOHvaBsKU3essS8BB4uP+I7yR
LGzpTiPV1bqknEvf3tNgrMkPIwfJH8EkgAumcCLCx5wnaMeqdOMzyIQuh+UAloqs
h36CWRWFVoOYoL+De/jrR/DZE+etpLgMuukk+h2bqoIxIWLZ7q7wwVDiB43u7Lm+
ex2+uEZj62RAqI5RTM7gIbDHAB5EmdWYaVXkQSdxlReJuwz7IS6quq3WZ7LEbM2e
eDHMB6NXXZuVSI1xt3CwJT/quz4f8hHE7N1xIxkr2t+kZBNEDQpK6OVOdJsCLW0k
OCFz7/o0i3Jmiam5ciIV6BrcJ8+BasfhlSicIW6IwsvGyZl2ibm7p5fJumRKgvzE
6napZgo8VPJ2W18wF3heXVe0S4KUwqGd8aihZAgvdwi5B3bj+GiWW8cegqrosjD4
GVCRzdZsrQLBGNIfVfX2rx4P1Aef7iTTHFf4BH+hGRigtAWcS5HW++gWprW6YS3s
jswZniK/VnRFUYrKLwFxqL3Ba++uAZmfNxU2LjgfPADS4InsjhQbT7uBPa4uER9V
qeSFRJifnzuYEfO1MLjl/crIiur1GiKQs/2x/oZOybTQN1k8JTZtajduIumGLW+O
yglNQ6kVOn94tWd6+hL4bDENH7/bGjOE1Xd7a7GhBfFnDCX2NTmmV65j2sWDa4Ra
mPSwS34TbmgNtP0QnM5U6m9UIYNUKO8fx3wBkXoZExvTUK775l4fay6SqG5xLT+h
bmcms1Fc9YGyjPs6soPdXpCSGr2dL/rF8Np4rZRPBoILd96ymAUQNqeFBT8Scmnb
L/CcvzEKiAphlmUuI8p0c1yIZDsOkA46Fqw9Od5bzhblPJcjQ9d4dPYBHx94RuzX
N9eihvz48axtwVlxvtxcaPwil14R0pbgg2evcJX2JprOHLzgDi31WChVvDFhaMzJ
GJN8OwgAnu343iuGduHD76Z6xhhVh7PlH4R4vKuL8GxrORO36JyV8Dd8f1+RYYcM
I+r4t0jgrSEHx9+MUyN9QFAnwXAZv8HxcXxNO6G2vPUBrOq9qwYYhRKsC/Hw7W+Z
UUvgLHjpjc2YPSbrufarmkhGGkrvUAo4uZwHtYpRXyBjKKDKtXXOo13In9IuqKUN
5/pu8C/vWnTK17MikPe0tpqBYdQKUE21UwHITtP6ZRD7DY65i8vOo2O4N099cr5t
wl0+bBsAZhvbzxeWpPpl/AKskYRlw5gQBByyLkOYeg3vuuURF9Nv408s+c6twkPx
yz69HX5ugX5n/TWf3L++zb2UDcJzqLOvtyWJ7yzxg7CYwR9dcdLRu7do8GcDv1pS
4fnQwfuPeJOEyVc2f2MRNko2D2O1CdTNA0RgDsbLkfaIZG/yx/hZFkPJsQbrqMI4
frkW4iHOCEdk1VEw//s+5qyjf1z/StDx5vi7EzyqeGREQ4FXe+x27mRMNEo1VXNZ
01B5ayBxraxpHb0Vxnf5rfdvjvM3H/YgiIFQF7EiPmgH32A3TXLMaT3CiESkLGN7
4A9k54bJ1AkpaXDzeYfSBlNvOHWyU1XWPkNrc8lWLVcYjUloiAPr5UYeInc1zXGJ
SDF+MQMM2ujyLTVkwe60T+mgJ3hrRNPRvjdFHeO2LmRat/bv/ZLOsqySvNTdelFp
nFBYK0bfnFSEKLxduWMjZXAr88iDowYo82y4mPtuix8mSnMUmntzqPIKH3AlUVmj
XYbXE8ynIn4KblX9ffvEgqPdYSEHtd0+FdqrR0Az0zjQcSZCtuLjfu4vqvUD4Q4K
RXFoSaFIHcs7+YPTUppfULJXJ1bVdQljFTHfzIewI7/AMXWokvcp5YG3fnU/LVVB
orh43yMACBUuOqsqECkBrwZCtAOwCeo1/neTzfB3vDWedHgtCLBpPeO7lN4P8mXV
Y4XBVVTfCY5jnpSks3WqaKrmpY7YyC8A2gcpvvQEV7Jpe6LeMIU8M9/zT2VjMjct
Ni8aIzHhFIDvsH+FpOOwOXxseXyHUtH9zsNOQ/9My82Fa2PYkvAAUtO3TWKZXbay
XjiIvNVDzXEwgWd1XPoc7JxOWNse4eXa731U5eoW0GECJPG6t8Scz2eBdTpqzTsw
5HYmZgO7f8kw4ynHimmYXceHGrbIWfMUA4k8zyaLIOcQhyFN6H5u+SEbRQmbTv0b
E51qUoyXPCTsQsHxiFD1FMy+2KNODcGjZQzQjE/0fvfKpvEmSy3ozygtcuKPVue0
6PPdpvSVQwat+hnFx4uETm7C753sXnzuO/5FyUR2ff+XRjru9kWmXnbpvGoT4tIZ
C18PU1WLchCg7VqituAFgbGuoSb9pwl1fdqH67M++I4ENG1Y8F3pmo5doFiHXz86
v/OZh5ftmNGKQIpxhJJ+8sMQuhFT69LHy/3PalFlRmqz1Unx5wmern54USz2Hmmc
BqvUvnDIzlKe0jQ9unjcKSlHfe5/vZIAQgZiJgVaVcG0HTYvTS3L6tVtE6SfsBKH
4cO90DemzZ8TfjM4CkOI8y7qMZghag09XMiCKGvEGNsfXBbA5i/84EODU6tuDKub
Fwl8hTUem2IoktlkcLNdxlDljCkZIt9/hoc9801PRkHZXzVVVhLQvdYolEj+UwZP
B6qyfcg7Gy+4hU5DMyhQqh3EfL+faOp2wN0bFBUK8+ohBclW9Ab8Eu47NhhRgS4i
5cdHXjwiCPPca1xt/msycFWhoDhJFQbf04p2k3nc6M2XCNsQ0Jb7Vpj/FVIvirO0
5crSqZt0AF+5jErdhQ2Q098pCi5GV4nUC3Rad4Iao3zVvOqp87kEn1BhJymYiN8P
ijvpKTvwSgDFcKQtDOfCBPnJ0bHK08+8QRr2aWejzNVOKz/+vdKDLHQUzWBejYBt
qy+hsWs6gC4mKMqoDzrEIwVS/JMnpNExC8LjZ46DAt5yJADxNT4sX/w4PB08YksK
IP7c8LZ+J+lbEova+GL7kakkYHGF8q+dMRVHL3p/wBFveixXy1FPhglnVWi1FZfu
iI+UW/r7S85YKFiC3JDy19D94haZ0FTfWWLigpF5fZituNIkv/XkJzXsUWkvXscB
KV90Vf61ZS4sVEEjyG0+C5jKQkM+5NYG39fratl/iDxuwAbOi3/3zeAz5pJIbh7E
jL3lSNCfGpUf9Ry6OPoHSsnnij83hPJGNrz5UvgSovI5Qreh26C+uthprzOMarD2
a4NYf3dT829EUGDQk9UQcD4uW5d2ZHuA5kGxsEDIusyQ0LzSs3m9Rm+c6xTAbsjv
y05fwzYrg85ATtcEFnJzZDhmsxFlDA0lQ711TkJ7gjotZavf83w5dQ7hpE9a5/Nh
A50z7HsaW8+JisZxPPJrNwbWF1VlG193ma2JgZWdjyzJ6RamVhr86eZQYEe24oH/
vLWqDJTrIu3TrOY1POEkEx0YO4W6ZRau0NN+TM8b0JU7mPUhLtse68kUQBQvppsK
q/BedOFRDQDb25PnYyz4uuzJuZHBj8Q3LRPvMMt1+M5wqPv+Qw04qErnGaDdYn/f
KEgrEaZWH/IF20wQmhV5/wXyBFjW73GRVAou68fd2+xYMtOaPkhbZ4OQ26xCdYGy
3xl7zPkkWi6TpPD7tbH+0a1mUiwF7RnlroQ0dmCV6h46HLQarLIbHsnUf82Nneib
16X7Or/hUA/2muGWDJVuOED1ZWbxcS5fv2dNx/99o5NFyqU0gink3JIKrNpS+7ID
dllAXVc0CRZ7ceQwLF1kJz0Qgup6mUKsiZP8atdmTDF3XhZ+W4ACFyt1GD2mkMmk
7PEmIyEKRuca97qMaBMUhNJPvP7orwo6ELLP3CwN3c+w7Hq0dyM/yl12yF7DsRI+
IYRcZ+hO9aMkYwWcUy3qddXzJG96/AuHLHAoyTkeuySGX3HF30q0QRDha5UB79Nr
2Ba+hBxymeP+vwixBsaSIApzsL6EpqITeyRXVYo6Ut8gSbtndkP5+1Qxhm0tRXlN
yTRWD9EXajpG7Qbj86o6W65SDhTQV51PfUFZAKsl0bTjrq4sBwxJWbqY+e7oBm0j
TtV1ia2tk8Y1+Tu8ThCJSqL1FYR2aUHUDEMbwG1FGRI8nOHMwVrprnB3EHG1+dsI
Srb5qzidrVBWFgDYXEwtBfqD7wShOPs7Eq5m8EnDwX2fUh5sj317pN7Kr8x8pGhm
GKzsRrhxs34LShXNLIuO0J9NB3sEnRi81eDgEkQPBIoSl91ruH6/orOFhNClDXXg
iYm4kkjKoPGzIEdzI3nlhYDiaFv6UMBuNvSMMeEIdBapPDT4gbfrxva6ZG8WKXnI
FAz5k1gmDAeZhYJ4SEXZf+pVrRSbuL4mZvnQAbGpOmTdU3mBiiLhxHrmA93+JE7l
ereH7yW3AuQzzKXbGXF8r9fQtSx6Uu82UJ1GUoCTdtqyV2op1iuf9ypLzZKpIKsL
RFo5wNFKq/VDAFrADN8HZ8QLgRVwMMTzpm3Rgko5BzwcAKb/SpfASzu+WjBl16qZ
IL9T5IohXnYWzlvTtb7+bWrYuCfGJesv3sGctNic8PSFcMXKCMVAJpWexy9px95U
zUHMWZGtwr62JtRWPU51LQ4Ll65X2/sp43DSmLzN9aiVWwR+0WbK0QkCQGtNyxyO
FzCZbtRGizo7VB6zTSbt2MhudrSK3mMVrYnkvNbqkP+ofMbVFjSbQf6vsGnA599s
bMy/Aj/QLdrxqv2/VCetnjMI08q/MmL5S8aa4yUh0HNcxZw4oXLIrC79AHzCVMVz
+rbIeWf8xTHR/aPMs7N3aa47uI4TPHng4yefahSNaNu56cdwJbLl7R9kZvr5esEc
ar206itZ0QmUMmKhIlqwja5POdBxC0HTJ59H3ycG29QDWLJjcXhzitHFNhYXD1vw
5+g3iGxyGXAFy0sUrIKaSzPuBtI73eEtf7GOFOgvQn5WgIKtO2n5gIbO/jvaXCov
WMnp5XVaeTsSj+Cf7m6rZ8EnWKo8xrEg48fvQlGTWYLj2UyBaOl/zCDMYAaTijQ9
RaHbjuBTWmwFff9bhAmwLA6HLD8HpRGwGpv29HpPol6n6yjTexvrquuYcUWcBfsQ
BMbjt75NiPMUNCx9GZphob7e79UJI/uE9Nlg0N7XC26aYkg1ySMgDBUFgB1fPNbE
Omo51Jdq2yUPG39ah80uCl88CTQ/Ed3EfT7MAa3gAHgybq+YCqJLgBD6+H5J6/4t
FU5CEi3vvzMPsz9PvnKyNTaqxPMcZOT8d/DHJBMCELlDmopScH87AJBITcgql/CW
Q3vzigWMMjO2lVtvDuYJsGiFnFGNXb5wV1iV8cEr7UstTIfSixZWCP1J4IOPKjqP
fiaO/iQT4tvMl74bm7afPJzzwmgrJKBJYShQROmaKRa3BevCZZpnRVkFOsPkR5IU
RNUjmjvRiCccnyKpRi3VnMMvPG95r1dNBolUtjw5jnoEqQgFNFq4vCPlIzQ+uqnc
VjVaP3AeBDciQjsGO6/xAiF4or93TjSlHsEYW05HTZ4IISSOjpkM0yMmTHFxBkkg
7wQLdITkKta92h4uR1uoJ044G1ZOzReEUI2qhckqrjH8oV53AtVegtKz5wGBdJuY
L26odK9Q0eMdaEFi6IQUrgCuHUs8hvK1Sx7aMnwmjaz6G8dE1vZnPnfShIr4kFjw
TTfX02RILVnQruv7ROqlJnQ/THQXPh5oKTAx8oYNGgRWLiUwbXk3QO2KRmtZRzjr
o168z4DGj5FHpiY3DXXOepXOVweKZsc4Ptba1GthsEKkrN+YRnlQNfSgdFaBS0MD
PJnoJM5otQtf6pl3CLCeeEmSAd3KDbe/Bp8qKuk9OuUdhQI5ngScUPtIHf22nf7O
uMO71zUjtmfYbThvILv37fZTXo6QIX3kVJgl3+yBBbX0S3OlL5Xg1jeH6uBSW/su
5aoRqLWBpoFrvXCogs/cyYTwcX/o0azYJcHi7mMTXA7+xjeS/b6RqVD8595L3tih
CO8xfy4L11hactoJzYYQsGZMQEfCEsVjgDpn4l5mftYvEzYGWlJglbMoWo+mSWFL
A4oYiHU7Cj+1PBdM/Xsshmcspxk/ducBMx3bruK7m5bX08efi9y9/Pto1VMlxsAo
ScZKcQOxVOp/zzOZScEQkyvm+RbTqBmrTydRRm3wtbhzZABAjQKvtfcRF8N4mahk
YFSkLQv+8eGab+Kn2MoUyEq+GjpywFach5i68dhq2J5/atwTaUi/rYk6A11HNdpg
LWjmRq2RQU72J0bsgLKSVLPbjE0W48xOr4d9ZhtKukXCEbyxsjzW7XMqBfGy+vnQ
z2QmnmNg+zrBCRbL8x3yF6kIO9LzIgjYX4yb2NHjrBDTbIgRaeAKJk2NZFYY5QsG
uOlPPw08GVGWBuFyP5/VbXgkqajJtcLRLDxEW9PO+u10Q4/tBXO3EKRjjxunRgSR
HfPP6RQTw8iLIE9m1FU25vAie86FUb27i5JfPV5YaLe4jJnomGtXc/jqoRzJcN6C
le9Wd42ipS+fOqLGsz7RmzQIFBfu6FMsGc+wurYhlyH4dfUhMU0DYOkDC3ni+yG2
YIB8wILvEdZ+qmM6pGC7O0l+6Js+3MpJ+HIj0HHG6iwqVx+hnm5CfbmQQWoL1c7c
FYrZuCPTHZQOZrlsv52immpX1XwswlKsGkCZo4vRSNzSvarMIaOqp+m4BNBjkZCn
fAwvrUVC3oE8ZZvwZLMyI4gsUwPPSihmFS7I77QKq7BdWl0cmpcbDD6jNmXiVScz
Pe7Nku52jzyUeJGYNVxtrR4M0ZzTTqeYZTR4I/UWK1e/hYP4k0rR+nl3YFzOixWb
mQWpqF/gXSfa++PJHHJk3o9QXt4taJIjN9MbNCMIKlIegAyEnPv3Cw6IwZZCQyBz
5Sh4xGYeNLYOkM9h6px5rVMK6+YuwnCmKiH/xOKx9d4XExKCeBydQ2SBLtT+aUvP
htKDXyWTFKOWuYraILK/ty2VgopT5kz6ann4XqIt6K0s4fGi0vfzYNwcdg/ur5Ro
fRWqvxp+ROZfK1Ms2tE1nOjW7GTZgFRiy/aYkqInfqNTU5IeGqbfd9NOWHqg2/XZ
tcXmCUFhzh7gJOzuaC79UE0MlvsBWu8JmiqusPU/BGY1KstG0+DGTMW7arIYMkUN
ki/4N+su/NjlTfY23OuSoNPL2BrbUZxQYpe76rv6N+XEraoN0v0tx7ZB9Vhsad1m
0bXeKiamMzXp63WZBRTJzy4n+p7Zbdn5c9ZyzfW2tdCClMmigTF6BadoIL4GTPZ4
NtTx+m3wqV/J50QBsH611vKSUdOpfdgGU/6h3PDaeg4J/cHOWRxmGyn7WdiTSEOF
dCQEicrvxqgznBi7whsQli6PQWdhi2ssjwD/La4xuN7m9ZuR/+ZaDUi9+4iQ3nCE
IS9KV5j4d1OmsXDLFoiBOGljvc4d5kYZUZ0kRPtSn9ZovZSueH/cgXUKo+J81JiB
R3dcC9flV00puwE1uAGWlADc0WZakOJbUEE8/kkV4kRppoWQ8ZFpVghaZ/0vOjVS
NGEORK23NIDRFOWtFnhChUcvNGFjcdEIYlaQ/3AbdyTk0pcCXbt86kCphTsbMFfq
krNTVH3YtkzoMucUjcSCC2wHbIXUmEHNU/gV7936hZ6S9FQcRYQ5jTE3+VljrgAV
yj4t+eVnTTuoaPjGQX8H1mV/do4r5D24JiWjtpjmY/k2Ko71kQFVlWD7blKjyD48
MK+NSUXss2kanpU0TBLGmRajhQR+geI/h5CDzCXhVMF/qqdVIO0zYTa169TUtV8K
EDXP1Lk/DkMF2CpakIGd/DZLMvOfpMuxi0KYdlABqSSCIJi9GEzPOTkfQ3ux7fWQ
lnTzrSirNM+Bl5V/yS9nzooDkYMHoJQm0pcqqh664BpjYHS55xysjpIIh6pC49ye
PgPCS3hKCATvP+md0XJDuuhO4EFi+Z8WRkPr15PQG1G3BEz705jY6QL/rEWyNY1k
jx6huEvJ3yqQknKF7IqAP8NQn4MEAa5DXjYONBi2nX4akuJ5SxjyLlkeelDrTx/b
suTdHnxw8AXLRsSzDjPXqMhLuDgzE5AoatpzKZp9d1VRsQ07lJ9JzAyxBhADSSzi
uZQ5yIRBg5LedvUX+98GVC/2t4/ri7sNzyJvTBfmIzNaRvBEgMnuC9LdM0jxWBxM
hQDBgPUe5cu2Mt9cJPhMm/BFQ9iVJmTITa94b3kP+A9PAq+S1Hk2xNQN4A+zBr8t
gk+JWUEzqOxE3BCdVt1pujJRf+TVKbBxHEdlAkF5kdLwaezQaryDpscE6AjuaLu2
zNGuWANlRVTudFlSG4SFAXe3eQh/UvHzIVlq6wFrc8c5rYyZ0wTd6PqboLABO5yY
Ojxh2c9L74nalwrGJroxMxSnjpD+IzrE6hHX1TuRultzxvR6fI5rhDrmsy6tMdZF
j3broDObYdgTg0u9tyVaHqVKRWkiTvI/iwecgZpyJb3vq+tRS5zKElpXypj0BDZH
Q94huwoBmXWZuNNRgJYOOA0S1JbM062vy8w4cl01si7i9PrKiwhBx+98SY90HYAm
9jQTU3QPAMpXX8otPc4aiKySntnHlwR0ZqJteL61j1hod9t1+9toQkxap6Fu6VwC
eCEgSxihMjkmnwBQ7/o/BFhLlWmD20x8I/QY465kPGIZy2EqDePFO6jl5Y5tO4wN
OBra/Aty6NETdcNryysSNAs23xQGmDjB3t1AzPd2ZXB0GOEpxxZKeSNVmgdtP1F+
F3c6+nv4dUvLOrgu4IgzeeXe7YjL5CVL5bhLWXJ1VMgjFnKCB6ZZrSh2tCpJjgKY
BuqdoFjo6mzHSsII+JV1R3TOiZbvF7YwHWats4cCoyxZCHccfd+5P1kYOGCJpdtb
W5+HtLoWXTMnCxlaBb3DCoCivHPWTdD0DqSBv6DIrJXV1vTQ+M4ywnWeJPI9FCnS
OUDAr+OQ9zNK+t4hOIaHNfH7he7+7rHw6LPBD2Ctq7T6H7mKamdkgazTOjjRAACl
1KmhZrsBSy5Hxnfd4QTrWkGyskxwFcO/HQP+qMp8GrtYhaNsoxiLMUyh281Wxhqi
/YmtwsokD9JFcFT+K3QtjSHkz2dfll+q3E+2G+h5LDlFON0AvQqT86Bfa9yc9A3t
9Yge7wNueHtY1rP43I6R1yP0k2UjUh0yogbq0A9FRSFPzYegIiPofFodS4F4Z0z6
qL+broxV6gD2OuZvClHz1emlczhCBa5j6CjB+TcQET+tV4z+W6F7fqCoFvJv9c/h
UlsM/Ewz0i6ZveVFcI2dBLIs7j060poIAP27tfUJU2SD1XbXakVMYTutG+pyrLAm
2yJyGEkuAPfnetw5A86ineFl3NEAbf449/r5FgqTyWjAQi7KhmchGjK7/Nt2PcIQ
Qw0fQz3yHiD61DE37uZx++61x80DoLjQSs4vMoS4cmv2TAC2V+V7u1K8uiQDtIw0
8DzUF3i4kK7CjUv+JomNYABiUNOQdeLKNED80+IqQt/4dGV5dQvSq4HrqI4RVLa0
AVm1X7Yg3IpPJDrXDenQLNHekudGRXbkMJg1ccWQEHXleszy9b/JRzTmyesF6G1+
J58MpaY5AZkf0XXCIjYcAhV0dd1F9I50/FygC4gyuYsrYDWrbyQaBiEtmv86Ruq4
FDpls4bKEsojYggX05OZL9cs7an60sX2wn0JvKurW9WDiIrwJUuYtrYxw+XGaXPi
5qs115nDXreuW4WTE4yGpiUAjplp2aHYmYN2NoLkAY+LfezIO4r7t9r8pRDZDuDf
cMOj8KijW3nhddw9uHTBukVzgmpTbPS5wPkBenIwejQO5AlS8NdAjV0zBTnEL+Ty
FDW5w78VNopidUI2629I74iKs7ft0x8Nx7cR4IBf8RfC3WyvS+kGyatJPRnIyAhm
FezKW+L2JBcfnrvsNtTDqVV5txrqH5P/HA7dO9A+J6ABQPhCzdgDPDynDSU6w8P3
dobY7EhBPZY33x0kPXIyuXIQk0I0bzY9trn6o5dPtDvOUuFZi/QuD0ew/eum+u2n
aUpDUJLerzwytUZbsLHOQl1R9O5qP5NMvOooi3n8KL1Q2yLvSwe1vwCx7A2mLoGV
puKRr9XcQesKhUsyfRQqKhFwKo18fjSxD6WBacRYIWitVwvH8gQX10Mnlnu2O14w
4aIU2fzGkLnuhQG5E135SS4nC8rdemflEjEUY0Kh5v0+OwZbREntmxpuGcUnsWkk
33ML5cQTGFWwQIcp9SdvUMbrTTe6T291bAf66jPftGXO2WoJGdX2y6ZbNcIPBbRW
IMd0EkUrlMkkKzEzeBlgQuL/bR29EA1MQaCpDisXWPlgs9lHQMVTsb/lT9/wdsmB
pK8omGOt2Lju3DGVh3hoDchcHls6QgIdLBBc3HKMQ77n/uQ90e14X+PGiotNhcPw
nb3nhJtkfCWlYdOSE6pQgPShQ0aZUYVlaxxxscU6cLgDJH6K9uXNSWbgjaF9o38k
DKgbcLx04FohSYIpynxjRxjdSBCdSuAg0cM4ShnpdBiML6pmiQ1TO1AmOanJUmNm
czseQyUL0Aay9chYrwWQsbb7O9kZizo+o8yLyVp70ytp7Qu6GOX9VPgfJYMh4ywk
8ZOnQjMK3zxgTvxZh7WVLWZsNzUH3+MMDYkLhJW/89AIQJGWXAjS6UU+F3ZdDZ0s
MsWod6NSfKAG1XZTChSyJorG/8HRgbR43uMB2RTmUGtMM+v+TH+FuN0fUfIumsGs
yhVbIZrHlImMxsk0kWnrdKJ08U99rNcK8LfL7mJVoNm9vQh7mrfIWoBtresR8a6L
sbwUYq9rAUkK8K6iGfy7eoNiBjiMluJuNlCYaQBehSG0YI6bVOmUxP5puMX3c/LA
aiFIEsqEYOtXutbelXUjJ531m0AI86dN2u0OUCo1hJNyuGn3u+ybf8bjKwgm2W/C
5QpBdSo0/iFOw3LfoC05XgBE2+lejB4CIxP/yArUuQwY4+BLiXtBl3hmK8UfzA8A
jgDXF63pbjPOW14YG1LHbdOUHBkOcYLMsltKHkk1sD8lrEludGpkYhlDNQ+t4uz8
WUuYdy7+LAZ44VepDDlq+PWuzXfULdYpgcpn1D9OBSab1ZDYle5vDPJ7MaEE14mb
/1hHCNAk30YAC7f5gHMljnTpnShcIUB6Bdrz4/Fplj4XGoyK5R4MbwgCilrlRTyH
L2eehrSwrdvMcVl3B6ELLl8B58Ed/scqtRKrHEz7dqWJLunXaxtE0IF8pcTmzAx9
Tcf2gA+hDvabXNySBTNL6letsxeK0PaTrJhH2PnP32NGR7PiSb2QhN7VJ2xdThfi
EzPQhdsUSfq6Kpf76mGJz8rF+TYxTrIIgXtFoL13Siw5ptvShhW3kBscmQhEdqx8
bOj+INZQpzVSqWbuCzIBMJQ264vuOLJd/ikMmCK0XqeWrP7Sdx3kRJd5njNdAYb/
EO4ITJFtHjXMtOEnEOSH62tpivfA+MkiC96XV/qmnQwpwEHVSDMsM1yi5Vpux7mW
7BAaZrAOTLNvLIM5dGSOBOuOLzHu8Kxenxj8nNRVaJ1wm7CHeNUOs/YhHT+rTkMw
yJx6AjG8lQnwN+6CcmLSWxwc9y+LPpnx46l4GlSU8MWiWoS2wJqNqwdIBqfewCgf
dqUIErDxki0ijeGTX+h38N0vpuxtDY+EK793cb9fRKRN2UgGjDT+mhnHeKY98jma
dluMEyD2AyRqSkTS5DLO5ZQ7w/0rwmbprH6HXZ9td+Lj9NrpFdPRvQda81lkfydp
EDpbc53W53wOn5VZ3fR9daxp7OyOf14wOiR3beAVBdd6Ds2TE0sMc0Zg+S5WVQCf
NykeGuKQ2Rbbb5ZeP6IffJ7R52FBzFvuZQGywWzukIEqdqOtBzCMyCR1oyH2Qbyj
r7vWN4cA5Juxm9m/QXXkDtBT6LbMSCsGiqB85ubSce9Hi6Nh+zTPEeoOlqSbkYFQ
STrVBidlGZIpICvLvzn4w36dyn8cpuyt0zLvPbyl17ReGWbQDQR/cqjYlwztEmJX
ltPXzsyOz5FM1UEOWWOmkPqfz7zRx+NMS2hZwa3mtB7yvVL/7KfGcopkx98Z7+2u
IiUqEJ7nLA4cSq4EUIiUTJu0u73Qd4AZC8qGQWezJuktEC08Dq20krNHrO+KO8G0
Mebo1AAxeMjP8zYNpBId1/GtftdG+k+CbavBGq44o+TABNJbYVOgabfvwhwSjUbc
xIJBQyGy8oFGumBOPnw5MkWEFes3Pgrg7kXdB9u65S5EZOBSe18AHtPvp9surT/0
XEfCLACWtnUd5b8AXOADBZ4ffd8L2YTaRatxeHe5rPRDidOfodnP/MbLjK17RfNN
YwaBzFs4Gf4AYGbT02y6szFL8DeUkH4En3rxFtFIh98jPNpLSZIJNBEQ1doMQePp
D8uOjckyA5i4Abdq/OYCabT+a4H08975KVqO2OKWbVG5pmp/L1cu97+fqI8YW79o
0YR9i4PESawQmUX+kgFIiKYzD6Thnz+2Cs7ztHKA3au3Rp6l7AImjqx93ZBgTMOY
ED0sCjBvGKsyQCzWsTOFDgRGIQIuAop2NsdbD08VOZO2OBlLO7LZsSB0/yM/2FXs
I8nlMpuZNaV6F6jVi1ttiuWVd6w4mmrkPnF7dfjSFkw4Bj/ImtuFreOi7oRKNA51
0Go4tEmHW50jxpT7bdEA2xd+8GxUmvCWP38EjS8R5Ayw7u26UHqROEOGV9P8xKuQ
xeCOHJL4FQQ7FeJnDLJX8vX1AloulFhOgxXhGEAO0QeYb5qTy5QBcLA/ObLT8bQ4
HAORaB5Q5RSuLLLei1xeDTjBOJYUBNHkS/GCFPXz519EGgoEXSq3euMckBMqbGGU
tlj1py7zFtw3oNM1AqFr3LKSZMgSCX+iGTVq0lTxmb4KolBHLfDKqpg3Dj9fzphF
9w2SrMGC+8zZO5CV7adkpCd7MfXOCcbrKT/ED1KJmhWhhoZywe76BED9tyV+6p8h
LmcS0qM8lOZ5ZQVT1L3gBIMRu63qYf948yObZskCP+4RBGzJ7bO5meJIK2Sc8INs
cxTIt35Zs1DjO1A7pDuYxWddqSZOAQGWZrb4qYvXytadKzJvAmdYONUjxkc+krbI
JmZ5bv4H8TAYXHP9m5B9B/pkgCX5GSVARDG1oGovYuNx3yBcW0PJ2rt3i+OYX79N
TrAs/sFT7O2MV3ZOBXF2qgvpA/Mz6+LmMI+u14QzQAV9Z79vw3L6576YaoCzJvRS
K0Tba/+QXTO/y4qxdnNn1XXgwZV7AI9OpRa8npFoYpGrSWf9+dfOUiJCKbPqjyu4
P7oZb8WIlMIpwng5gGgZMzVipfJCxvAMRK/5tQ7DHTdlUg7IAHVg/LXn+4dWtBzK
HtkCegaOI3qGhh0jEa6S0pbbm+JPlVK9bmONUGvUhiV4U6wvd3Fvq5mpPke8Rw3F
FsV+ZsFh5csgV/QBMO1CGoVmm0wEXHs/49tOpyMuLnnK8/+9MuudbC1VqmJK7/oC
eDJ8rnc/gfvUNIAXJt3ojYjMEeI1Nalo0hP+dbZLWeam+U+gEb5ZgeYJnZwzO6aM
QGGnq2C0bstm8NntUOT0tV+W2UHlOmlfXMCU8cs6X7wmwYfU6EuXbanmVqnBuzZv
FSwI59eexANrtJ2lw/zi+s1MReDA8QwZ7prFVzeoJI22zHd4P4/8uxE6ecYkcYtC
BmRuMnuBNgvcDeW5PRg4g3K1lgNriI5ijwZ8RYbOn9VUB1+UrSmmnniCho6+rbe4
PCrfUOfO67FxBmMOKLHvwVkLDsTTyRy0pmWBvlWF4tez57+yHzM1uHxOzp34RgZk
PMX73K7sb9ErfbN2SAd6AI1qTCMx2gmLIVAGSBhS0mqEygtwMjJlbkQsTWmSLxVn
jTtHTh38L5czIPOtHkPOnwgxmN6i9AqQ0MAYOC3adbNvn5I425J3Sejag58VpW5V
lknTJHLXPNMUGeNqQs1bOlyPDURd5+kl12VYVlzCXOUIZ26m3L+nIqB0gzkTRfmD
p0Y2F+f93l18LPEpu/bfK49Y/JcwOfmsc2ff51W5d5plyGYH+/gKT0Nr736Jdu0M
v+iRcNNLJ3HQBBq7uWs3s9qlhsaylbOtsJ8Y1orsUo43lVrpaf9gOwNtEYIg6PEe
RyFwVT1+ptLiDjuGNjEgbjHYsoEwIhBbNSNQKG2TmxocFCWVH8DTxzOcDQ5gOKs/
b5ioA95TBnzyxadnqysPSr6daU2iJ1zwplw9EXB5TB9BjG07StzOioy4btBxILN4
PbN19ZZpKNO28v4bhVQ+6ch2KMfntUNZq4F4uGaZMkdto8oQicJYIaYL0beYoKoB
swEefY2dQYxqQ9U1Us4oHBJ1FVQOVwI2Mq137Z8/tf/+EZQn4nCNrt05qSAdNkp2
W7eabpM+KrziYOfoAIH5x4P8FbGoE5hmyeqDm4PLz3LKuu82qfctT0vaIN5d0Z+0
PnJUkJYfqcLcZi1ZwEi6BRf+aQfneou3xk4uU1i5apJuWH61CTkliB7ojINuTvrr
RpepLhu8KJ5pYGMRxJBgPGeJd/o/co0kc5+pfuVTcEdlPPk9oCxjyYSERt9THiaU
csX1XY9eMipL7nLoDxGukyelYG74PjCZiaLI6fx4P1WbGdO7snAR4P6aavKZU69M
HoB+6Rhsj9TpFyVb9KURMVBCOwxmiU6GYFkRmr0EDbq1XIaccjZeC1FxTrFXZ/uS
hEUognATK+eEdeytXDjzitmsieefMiR3MRBY3WQTR1FfXM4QIgk4lsAzmb9/MCEW
ETgMumqCQCvZJkNdAVkkVQrqWAxlPjSGJKuc8kZs8vOLY8x3vr1Ue+uG/pOARxTX
GzuU6SSkYSYzDrzBRQ1s0N+bKegav3LLG4r6zb7UHV6Eqtb74T57QfI6Gi5fZiX8
9J0ukpbl2fvRME46vwld8kHpShrx26+gmnR6G+TRtOw0JhZFh242fMpcmIKG+Thp
SzTlVfKwLKRrGmv9u1DFYRnnD9O//rdDIsMg8r1kpXKApwKAqi6THBVG7kvnmO0a
gxdhw4hCJcQdqBh5M4+12NQqx+uX8mml5zB1MookCnIOBESLH+cEsSg8IPBr2+0Q
psbBplhVUz1W7Pz3SRf6urt1YXtPn2styplEqGv2ztbU+hEoekZhmHBKhgUYZyKe
d0ZlagzXiUipNJvRFky3JPBX4+4r2Ww0X/D6eXmr/8mzwS4XbFFSAJY/7b3BkWvC
cREryoOxudQutsOz/H4wMi+FTj08CAuyKAG9weogA8mwnxR+3+T86YApITMRGPkD
t/G/Hmx/DOKkgP3C7vWDrNhyamyDz1dOoKLhBv77Wk3IlUcQo6s+zWqmWPg4J6R3
kLAN6HwKDNEVHdRv7tA8nbS003WOGGNNUlSR5Jfr0nIVZL3ovvd08mkLxy0ltRhh
PGDLIuE2nX1dpukNyWHi89M4fE1MOHru+FccH5zq7uW5qcdgLuFWrQP1K1l7PEeY
arKft1065eAt3bJTx+5gM+8DBQmwiiX7fDAyEjshOdbX7cKcfLcz297ptfZ8uNwv
3ytS57ORAVJZ3LWLMcnTaRQpVevRFi5tMMneObv+sO553IxnCCw6kTedhW4Cf7uf
hPLSBS/EeaCkh8xjjGSwqUV+gLl2t9Te4mrM17sg0iGPQDeZboT6R8EXE0kSpwXl
wPC1LvMysrLbrvywYJWWBK3vro3jNArfduuuHAkZ0iByhZGT0yYcUmE29AXyTAo2
Vu+F6AsHEBUKlgpNINfzKZHX9hRSfHcT7ECIMZYXDY1xpcenpb1qoLIdj6ZnzdSa
SYUi6XYaRIVYLTH0Q9gqQMgT1Uc5AxzrdfwcjtSmlw6OAvnxIVtSixq2LGSplAC8
svEl9T6qfUi9s92xuUS86IsXHyl3TwqtPpa2euIksLsuOoLVaI+bYEaeiPykcXCN
9wbDDrlyFfBJQQtl+38OqgdGuatHnj2kqooj3p1q856wArZVJDLtIibVHpTQpH1K
tCDixuQLdN4p1Oi73g1a3D6i+GOd5QrjRwlQjh1PqA9Kva2tNom3EEOQUeqAnZKy
Oj8DaAN6I5B9OSnbr3Pr3fM8/qlbgn7XXLfZ59psLOCnMCrmO1tGV0iVtmjfsV5C
GyouSttHAvxXIlaSxS546lm9rLuJHRaT2SJi1MwvY4GA0i1xfhTkqy63dNkujfNa
qkQIyThaGSvDrCmKv8vWCVph0LPTFxNMwHsM/2Cw8j/mhOnBjY7tzy9OBbJNTMRR
aW4uiYWB+JgyZZHY9rKseYhjQvskdxok6+82laoPes5frgpqO6l96mDpoEOw/jwO
I4IaDiIjkxiDNBwWF8EiyrQsJ+cMjvH/IMnGKgsHeiVvuYCTEzH/hBRxVj2/O96J
mpoeAUZNv74GbJynH/EP4zfsMo70b0Bn8qfhgPEm0tTYAut3TcfQMYozEXcAjdhI
wQgEc6A/bHe6SlqTjW2aRdlUL/Lwkf32SD483LXbMo6JN7upbCb7Boz3R0ERX+cS
FjPFtYN0FKh3DWKsJeqMN8M6M4IZ4f2wIpFgkKb+fTjxz/GF9s/32jBRQSMTzxjk
HJIUDpcto8BvLaYeKry7Lw2h7itNuyKJNhtRVUvfJoWiF9oM/KJgcdwZH2+8rZtT
6IhzxmbkA9pJ/C43biTog1oZEG0AUxhH8W/IvLdRQ+7wrhGxfX4JnnGMR4pseVOS
QQgobjznsSQFSo26Bhf0w0BzOZiPv6JT8YCMCZDcumR958/cV2pdQ53WY8PkeUUF
szItDcRG2FlhS1CzfDBYQeY+f4obDir2vcrPJitVQK+YnDXwym9v3hzKOgF8+0Jc
IFcvayEr9LLkzzWH4JvQLuU0jQpj4MMWVZr+j4mJTpl/sJyTnWVamoECHv+v0Wid
vxfAWGdbQ/2UIXQg0jMKHUa17Z2KllrHW8ySWa35kIYklQAmK+wLTnn6EwUZzuKq
s5APNUbZA0BuAZ+HTNf5/1ixIsp126sQqKNQ304j4rRJe2uMJ+jscSVqhINeA45K
I5QVo6eJkJ7K7+El6fKHCJxXxU0Y5an8a5asmEHfV1kguDNwFTUQ9oZZj/sEiNk/
6McR7ld0QpP/HYF+2QYw2wWnS9FUxDdtp+mVr6iZuPiVdqQvUEjsAdpu2VsrF+0y
LWSX4ivhXwjvyL4zfLLSEwtQVq2MPf8qq5Ie3k9RhybBMXMr2S5iTKxqfB6U0uxu
yH6VMhLJXtgF4QS7ECopfRnuYQjFoiHvfZQiY7Y2YZ0tAJq+8graeP1l6Z5gpiWU
7Lh7zOX/TwdeB+kaT0DwSX4Zl61uWB3J+OWX+l8wc2lt/tw9tvdHkISXM/iuekKZ
YZaCboxFoHC5yCwjY8kvnlil3blIfEdp7xwR6ZZM/zA/VAgNKnIA68LIGgnrT96s
q4rDTJJzuzsEkhC/vuVNVdBdYY+YMFGV8eSmxKZ6hwJ05Nj8gLUUhkN9tB1J4BS0
ZHb6FN3+QwMVhcYZ0P/+a9b9KkG35QPLNNm+Wv2ded0KY+YYtp1DqK9xlw83jO8A
4lv/7EvJRXUnAQFJQfu5l8gMeRpcN4zAgoy6PyBHphwkzPHr8WekMtkQCU6Tmbjy
gTJ45ey7UpujEd07Qi5EbbIhOP8duaKi/A6TeXf27N0TuGytmb5bo773nubIMrQ3
ZSJczNknzFk4TBDMnvMl+Y/Csykiq2k1z/6oBThzOx/G1KMjtU+t/huRF344eWDm
9bUVNeo0INXoSms6Cn602iO3yeTmtxnYZJIjOMCrKnR4jKuLVS/x+PVpBsaDFMMd
inXsDyWGu9FlCuJw5tNrmLpI2zAxo5cl4I+a8GT/8Gs1aN0oJUOLrFy+lsYo/qtC
NOj0X2q72kY0aO1nWF0jaVfq7bihcZSnWR2c3iRvmRMi0Vm/DJAkBIEAjxkq5NVj
/Pg+dKqnPva+ZoEYc51CJ/QSg2TbJJZLm2cVfjQnbln5tYx5gnti9yiD9TYrtrnT
rArdj29v5MB+am6dl5fcRZoYpmWmBqb6lI2cRValrNoewvqyHEMp4JiZPG3FZoYy
DgUUss7PWa2oFBpCxI5ZOiFUH64Tc22saQcb7YnUXBoJnaPq92N26MK+aInAaJrl
XYXsrrygneuaYaJgBNstbylD+QFm0Pb9N9XSWY55luuOqfYxpgfVyehwHSgTYQ0U
fLviSuMf4GgEgrTj+IO1u10735VJoOujauERamp/Zzca8KNdn/AsNrXVDpc7Cxa/
cvqjYJroN3JFepqHoH2AeSHB9YcV5uG0ibXhnLbveVENtLcLye1e4Qp+z6cmjmQP
GsU69PDB/q15Wb7vZ/r/nUdHVElqlRt992kXiKj5OSAv5erPo1xsp/CTDESiO+Gr
BfCOTFl02GeVhnWPfwpgfZjaN+19/GJTvuSrVPMOkwi9dHjT4FqsgrDuWI+15C18
dwMIbXRclgHY4wyUBv1wt07lW1oZdQhLU651puFXbhI/UaYfwyZun/4YqnI6j54q
5sacFRY1pfrsCAQmGr/105/iVCH6d+PX1Fg3TgGuWiH5u2JuOekfp5XJSKeK0IPU
STvsxJp4kumBaptPl3OEGP+ZYSz3IxGRR1TYowJeFZBvIWm8l+g/dpt2HpCIuREu
lUc2oblZ1dBFOcITGgkEAQgXfL/dtQbfSg5fgGTzovm8p5JN42c+LNQMkoreR1Y2
U0LO+agkFnMKycB+G0ue6x8GZ3H5BalOqkuSoKOGbYa4kKSM6IwkAkWuBbQQqs5M
p+8Xgacej2yo+n2Jgpyc5ZN0ivGn6G4zyf7HRz1VBfJ6JIVix/gilbVSpX+Bo3JP
OUxFKfHeXIhxZKwX4nKWVST+SZuS5GWXnmw0GgTEyZQXO7Zsjv9Hah7rsfGgd7WM
P4aIM3EqqTbJG0XNr/k959KzH31ZBf0E7waZshpWn51l1ehHBWMV6ReLrUpzTn2e
kdPS1J1xeCXV/nlhAh4iObzvTUf2ErY7G/u1yqS6M3sBiwbFxw4JAq0PlUFQ73jv
lJISBPSlHpj8NNhVdFlbBnRQdALImSN3Z8aXyTn/y4d0xc5bqawS+i8P0idfIAWD
HkT7NbH5d08Gabc6LHLOIORI6r/vhQkedhZ9bJu8HlZoWBvDaNNP2tr0laCsxWpE
Zc4pTgT220LpjcPIehpPzz5S/BTctr6QKfH6eCwLZB9Xbar+cCdMB/YT+YwvRaNK
tIro+nBV3iKTUT6FEDCiHCtZz4gd0gcQrsK3pnO0dlHghyMhhSB3/22V6kC8dBNf
KEiqwXlNOZLnu+Eux8s9TTasew/SrRep+/0jJs2nEKYPf8d0YrHgFTwnbHak6PLr
tL7fY6c+pn+f+z7tNSZyPvO4VQCy0XV/NPb5n2Q0usr/RFsBVV7dqqP4MFWmpPSd
XmZxT9vOlNHFSFkN1GI10HLDyeqgEKqovH/Vrih8M72FexBNktGGtE9xBDD/3KFZ
VuaUFMcN8qdtLVgFvXN2hzK8z9Rw/QA2OWjJ3yfEY1GibwCyY/bamSshqXJZ+qtU
BitPQxo2x6N1F9JjVyZk0e0jbVRhofPfzcrXJ271vSaRRTJUtsKKMntfauMTY5uH
+Zxend4RWrpokFMwN015YdxruTqYQeiQAhkMVKpngvQetXtRaxIc1fQmklqKo/Fj
eSnRBXBYOi5kOfgQDPoaZlTxgQZ2U4DxuSeIBcmsXrc1Q5fv4AKbo4l+2rrrp4kA
RKlynPnaWoYhpZFRNRAgxE2EFLxdU2c98c6r7ZGbY0L2S+KEqIP5Hs8xEmUT3ldi
ZxmOguzHMeDZHUfor5KsjbSNhph9tMPmj11Tl9uZn5duseGBYWYuPlSp5h6+BlIF
VcJ3csI7QhVKQNM1/0HuHEKmIQ4aFagc6kvKHN08bZLHgHF5PbBgl0Kyei3/FvZz
TALFGfKbaKrhNB9/PF6CD7Ry9/eaMFvq8duof74Tx3aG/NszKi33M5t101L8WvgZ
dIQp7nD16fAwiN69eFjklluYeIOhvVpOrsIsiL60TIigjzy7JG4ZInq7ixi4Ce9F
kvUaej+C1c37443EZMo0RaWwWszhmr5XY7z29wCElegP/TKL1yAhKj3ouv2K/53W
eVEjGLBPK8c+6FrHM8UYmQiew4Z8y5ieHi3Rx8BrGL3w+/JPuweV94jNZ75kciCG
if8C8UY9NIYZFT4PYxnhHnJbLHZ3kg/zroMPhYrAYQFQQefG6UhihHN3tKepLSq9
jwaUYXGEpuKTn8IS8VEv2Ry75Up/79nQvxBEJIRF7WFWEeWRWZGiMV6anr21AzCP
gXEngWdLhdNlJbNlP9xk7G2z0ODROCsBg4dhY6BnBRYPXF27jyP1Tdl958S5XR+r
joo7gF1r6avzsur61oXA6c328tD5rWRzFFSxwIHOschtx7yYP/3c4Mhrn0S7TLyK
HS7ZmHbzXTs5sCh9OGf+l2NwbxVVzJIuPl7JWKCyIcySjQTAzK9RPRRh406bZpLY
L9cRV4KsywHNv4UNhExUVuvcbAJwAR1qjNlghCu1h1uRrFOCmGRGdAKXpIFoilEx
wy9NSVfcHgI4dN5tP8JzQ+iKS46UCi0FQXBezJE5SJRnoe18SntZmr7NhH5c1pMH
v5JNb+ukK1EFMNu1/ewvjHQDBtu/Qi0x/kj4Js95Z+DNCgGEwy1B6mbKUgRbb7pB
BzUME6nz96ety7m/ywMV1j+RROZ+nY6kDyn/mWpMWjujrh1Y6wW7Vtht+XflfGRm
3ySmjWb0UybLuKhHAH50Gy+4BRH3yGsbffBHBeCudycrmSdIoZzrLDaakYhglLwB
d8pd7n/n+a5cyohBDpKk0EWQNb32tR/gGP4CXg+WrKtcV+mok4HIELNhj/l2LtjD
HHjDhGiQM74H+6nXGMkOAMI+aYWrqZYlNvert7M593lJizVln2L/2U64cbaknQcs
/qgqXhrGtV4sb0NVVIp3Ib6hEDhR3IKcb6jXv49K2eOxw6canBKBtvkT/vxTtEOg
gjuMS1ktudF4GW7pI+Tape7Qykh40Y8hhAC43j7pyVI1otA4KbcpomKPDN8W4zOQ
JCyRf/8gN11xGUCJH0/w+RxJCpxTBGvtq7OycQ9LMByxTnxF8xaLmfO/dor6frl4
ldJ/viiF8AjZysxq8zsaMcakdWQfOHSIa0RejNG3sCx+BCwuX+kcbvTX7iU24jpo
9cNIFkdhwWZtnhVP5zDPU/oB40TgtCzf7L+O56uCy2EMSbydTcrVQDEqa2QW1h1a
j0x1YUNL6XNnG8ElE3DzYO1/Q5k2BKgrXmtG9Uo1n3m/Xs+Ptl7yIKG+/2ztRdAm
K92S7eD1KMns0RA3talMJ2A36J+pqtAM7lTrhALnpDlI+bM/LsGkzX0bdJESAHWP
sfHvbwewSeRaaIH/ri7euLs9m23v0w58wikbOYKknuIMrSRKq7YEV82KWkVGDaxq
HmPPyV3yR66YaKpZkg7L0ntqmHKiXz/ric/txxraApkV1VZjonuPS9G8Ffrc8638
NK7TFFEXid5SYqC6grUUhsBPkePCSN5shHTwD/ifLyjV4v+8kyJaPMlFJ2Xmk/+8
nVIHEpg5WtVElB+AmzRV2T0yIakGmiwXoIOQ91dNZOT6m0vtTistTmeLHIUENJP7
Qjp9FnSa4KVKVV/n9gPahYwS7R0Dpx1HgXWO6pDd8LlFmP6R4RqzCSkOsSWdq39C
JzrstzgVbth+yI/gRkCN1KmypBxDqc3wI6nrGvl19HoHnHFeQ842RGn7RrxRq/HF
3zy8KzL7gico7PwIDukMjGhMzn415csuueOQqadzPOdIn7SwyLZ+O/k02zyCP53u
M+iZX+Awm2JG0t61L4/f5cgYPEWqhU42In+qGxe2MfyzVtpE9hdGg7pcDtkGSSGb
LVIBZsgR/vGlDogmCN2nG07C4E+QhjNDUC3G4zTmMJNuIJ61DJMoTTqGVhO8REJ4
oFo0Hm1qy51r6UfflF7g8qKjTS5HmOr3ELKekNxKgLuQLAUf9HHZFbbjBlLCFrPO
j5+R7ircVg55oC6nebX9b12RKoGT9j4HatCe7qv/Hrmr96DOdX9tT3LcJHRHWnWC
EsJUZilg43VC1KgXS5b/qapv56jehRZz8lIvhjdwy/LFfhRumU0YHJJSvBHvgiXr
ZJlq4QVX3xD2lSE3/V/57ljV0Kzvf/mnNKO8r7rM4dHlvZTz++FEjhMlK4qOlWZ8
cWpB1tdCvh3AJPumk5gBcutYmV8XKmKM7o78xbOwaAVd+voxM9O/xvBVCch9cJhG
OoMDZC0ux2Q2f0FbxmSg+5dcrd6iVQ1EGXbhm8tHsFLes3RhSM7NV68yAL9B2vQP
2JPi6qIqozaMhmaXt1akdWuajSeRPJ9R1xngnBmHox0PxsTV6B8LyajJlEwmBOSh
JOJwLnoG9190IvaGWpTK6QvSRRtLmxypob0rXFVoxcKS0fnYUHK3RzctQ6XcPNnd
4xQN6JGkSmidjefomKIWB6UYOmuyjUmhChi2QjtLI+8hlc0EoxaD8vDIB/ckYzHl
0IWBuogwqjh+Bh3Yh7U+By4LcD3ZHbLAUKb0Orq7xp4kd3zWkIDb+oBo5oXVjw3l
sUnkfnWPE27M2EMSmKQjaS7m+H9Yl13LiidqijbmDQYvZKR1xmKc6FzBTvRyMDeY
1Bzx9GNVuCNCpBeB9CRQqO4BD+03NKMOqKAlcwBVlcq7r5FDelFHxb0y7L3Bvog/
gNgt6RAauHHKCIt1izl8UJIoZtRrMy3Iy10WeW2xlcgwnOCZZfSlBiITHmzS4rzF
p8WKlBFqOYA3MTdouLwlC7X8H4NTdbH1ZJ6NjRQLaC2CDcgQ37bnTnd6rd6234m9
O/+M7Rs/7wBHhWaY94LQsS2PzvKxJsYlikQ1/dxxmiDB19QsMFr8rdAUfbpu8tVq
RxClekzo4RCaWksNuosYVa4h2iz3hku5xP43j1EPXdpU2H7wvF1rSPtkTR7a6Fx8
W7Nchw9w7t9+eDgjtKxSIlzu+zamnp+oBD17+TSo4ycFRIUd5v9siyQunqxLUHrN
ttBw6i6vHWvgu7wjmYF8MNS+eSQpaaBnTwL6jOMYxD0zYZtPfQzF2gMr/mKFJnMZ
cSmkLuDBwc7fBWPOnThCvU8sJTYF64NMHpKYqVuqo7jywyp6+4DvukAXJvGLAFxf
ZGaYm4uyvbcHT8THc5Fj+ekFb7CgHrMQrH1nsd0s5ZafWo+gy5njbY5NRsScaNDZ
M6oDqzaLVl6z8jz9J4xmkhA+LNb+XBqCVRJFnpJbPJljnLe5PLH3yL+Lj84Y740/
ytbz5Mo/ncaMeTWvgfmWc77eRQdWgq0p+7FVZTT/gIqA95epaLIfWPqffiSNlzLb
lXgvMknrYDlkyp3B9s97fS5qZ92TLwb9Y/CxTedTuA1cxoHn3aHLKabM3oTpdrgG
kLDGryYFK1ruqS3H5+IunDv4ZQ0sshbLqvdZ0oWMb2SYLGmAxQYpjmqWJuHZ0MK/
lgCOCgsNJOp7ylCk0PeLs73pkU01tY1bB0OoRgnhu8soLc0XJ27U2g0GqGd8R0Y/
mMQRt54gapFBw0ChhsRg+/DfbAI59Xc7+YGbXIiRVI4g9UKGhPrRaQXGovaHJ6HH
jzXdx4x+l9Gh13LPTsOpIt97RB8QDWYjiupgz+nODE3TlVLf2p83AOuBTasxRJ8z
jhBs8JP7qr7P5z2BcSy3+wIVFX/dHvHxElzdV1MxFnzZTunJnwGR2NcKa9k/Wm3P
B7IvheJCzYh0707L847Z3vwoy/iUWu7MfDGUACwe8SDOh7K+pVMdVtw2ffOKYV3y
CH5Nc4s6JdOoR40di9kJb4skATjsJ4Gylze/LvY9wPEv2O7WqTxrPjAbu/yrLe4m
6ISup0fnCDqR1YvXwJHezqO7Fni/UlzAQTaIeVGfscdRROmGjr3lzQfOCNKGRcf3
cBVoGszh324m5XxwEZNjmO3t+1uiT6b0/G/VNzBW3GvyWunWY5qC/OFHu0S4nD8v
yxps8wKQImRuvzZv4hgFfgRYL309dfZQpHVFIUWqzI7hQCz8SJX66rtfDoFiP8Hk
oMku8LpQ6fTib78CD1wNnE0+aBH6PtELXNk5wIXDf/nUL6oYvE6pY7UYkrYfTnKa
RkR0vqp6vVZDz9aS9V7xIB47B2vLu6fdJCXex0w74vKgDT032K24pkCQolxaq61h
e9bZXvzaLLg2voff7TA7tF+xH4rOz5Ay/cd8K8rjFP/0cGxIyUbmRwoOXwWxtSF7
OhNh5qTUh63poYucPgPO1CELYiheC1OnIDipaa0klIUwLLpOyMjctx1w+Xg2on3a
IAudKWQ6ddMpPsccvN0w5U6B9vQ7sVeJGtUTRhJ/rDLRCIxkeUIYqmYM4jp/1EOM
J4KKepD6Ev2d0YDyHAu27FHmYEYrz/PEgSLlpacb+G7UN1WyqdNkJRlnzvXGQULa
g/8hhX3nWzqtOMkEI1WWbiuvd9cbdub60j+MZergdvuahjHrUK9PfBvAQp77p3vk
QgOujJSkffzV6kdnvBNLpcS8XouaEcP1rKK5CQpfkl0vG2JSY8T/dEOeCjStZiDy
CKNSZlewC8Kl0vF3A7arlOeI0vq/nylvDkHfK4+DfPuLPhyURYa0/m7zwlk/Uk8j
4C1lVxGigCwYCIn5ejFV/hfHJzD5yrLLZiljaHF9AL+CP8ZQnmyaTCcaJuKNtBx7
TpkgHi5QywCKdVCpcgd/kis5lCyDCe1gVPcsMgAbbGhz25JpnsrNYWJSudWeHvm3
dbEhObiZJhvn5ag3uZhzWGuHt5R6EpJlys8nnBgO2EVfbmUOK0DFwpweBXeTykpX
3xopKift+b+v6u/e21sofhqRu0P20MpdqCzxRlF2WPaE284eu7g+f6Tb4d1waKaF
qRImdSofgNlDTsuS3FPoQ/c8CT4MHY2aWG7YHuj8IEFLhvFyHizO3OTFGsppiY5N
RXnNhJHuXkTtcOJGh/a5zw98pRvsWkJLnm7GSEKHSNBD/93SjB5rLvHSIf8VeTNs
VGTKu7fRjcMI9ZH0VgqffbqhEgJSYGxvjjE9fyUL/Qkx+80EqA9j2cvK4yyfyvCD
8qzoueEPDmz3V883nxiLgBELm+B4qx2M486gS3P2nyqBypmlSX+6gLJv1vBki4EY
GFeKbEcan3DFO1kdDS+Rgt/DXU2iYk+tklH4/umhZYPRz+Nv68wmwaWLYOUhvjHf
Q9o28pGMbeC/cktDLK7BhbEEn8Y3xKAjGzz128G+HF6CBt53cFbSZ7ITH6vRUSYr
mDeL2l8raTjaevNmB9bBE9xhQ41JLxipZwkYk1UodeC1vu383u3Gkf3zVpCB4Xdm
Uv7WUlWtP8YnyTUZ9VcKuCJZnuiE0KfQQA0KwY+j4H/OwriQTEdo7QN6HT6iIx6h
gcZwDiYHjNCgsxVRpE/0EwwVhP/Ab4r7MzYc3fJGcBMyngiA+rvs7P8YFki7lWMR
o/SqFn9bBuVu4xjAKrPAVaJdbYDzXs1ylshRwq7ZzzU3zwEuo8Af7QpHwtOzBkur
At5MoGIJOlmOjhGwAtL15CLYvoL5K5JPg2jgPUehBC4I5yqpzKu44AYrsdQcFtsg
mxth/TMOam2OmOsSM8+zjrHPo7NrkNhXAUjAw/ym3AeQTnpWHQ8DUrZs/LOr9biz
2cQwVY1mdEPrW9XHh2FiwtlDKjzbNN6fvhf3f809hojNGybwWKn+LBXJNagzpnvX
3xzrvpjy5P7neZRHFrPJH8K+i8rXLawm9D6AVPnD0Lf6Aq2B78X503ax0Z+DlIOp
LMaL1dv3uGP2gZzQlK6FMwxzWlkirj5zWJgP++KcHJLd/HN/nVD4xClJl0QRyGMk
fziCARoDdgV+DKA68RDiU6M9BNwb0NkYSnhL1UYA1uIuioFD6Id8FZg9IT/v2I5t
RW4owHAA0EjIejciBjbYfZpOoC7az5JYWBs5YYSD2bTmA5e5bASvDed4/J2aJMbu
FlzZlVkJVmb4tPoNql6sX+u/LtPeF7wJaXJwqz6efN4/Q/RTCZ/QTSqOv3II1zeI
C/KM7r25Vs5cEkqMFDIbuW8FpZvwDxqkVsOaM5CEDFkatBSDdgfw+tlUntD/VyQL
lG6WSgm0tVBt8VAjqdPxVjv8c0LSolHCiAAbaGKPR1DgHyRTxytkF5QbW/L0Trow
SpxZ1OF/chIhfbiJYLHsaKPy1ExC0E6UqQ1mOw+lHj28Rr/LW13VueUpqoqafAL3
ITsPrRx5zyl6OZqpoej0PRd5V7s6DBzopcaY4yiynrEjf7MoZF1RgI1X5Ac9PLxN
n8/7g+XilhWMRybh5gyXjFIM4J8ZQJ7SsbBEOLw2LdT1bTfwS4UnHaRFIb+Scr0U
6XHnw1/B3UGf7mQvOqONpq1QX65ZgQGsqbvSDqEZg5ErVDmkKEaT8eHDNEkf3uxh
9KP/0ohZ/zt0BV6iQlDM9FC7zVwd+hmHVKkkXMUx76imt1VHiqdlqVqvRxJasIt/
NqiRx0FukA9UQtrZEBJMIS3swEyNQB2/pcs0XZSdv1EhHDPMPnxJiV/cSPRnvwWY
MMEgzEAoGU9CGKlS6OkhLEjzwVgIE/dZ67LaOBbxBY9Ffhtf0PjRl3UUi9k9GSjz
EqmAZwLb/hWlCEkbYkGjMEiS/ReqxcJAEKwoWLbIawhLieyDO1a0px8E5+EU/FKh
7JQH1UP3S0H1qNxShLtJQVRI2DTEPFKStZI9rPumzldnPU35Pgru32Cls3BUrAGc
sqZxUfHrEZUWHH5USU1zwSRxI0D9Ndttz7kYRGbm6ylIlBRq9FL5eNrYnEDpVsB7
x+dPVHooZxzhtYEzTnYJu5knzYpiR4UIfkJ0aCuVmBUBVTBCxbttg5F5uyseNAjQ
scPYBAEmCgsyRbXtPlI1ECDD9eH4+z+x6QZGYCzvCSs/tiHvY+HAL4sZNXnPlclx
EeqzqE/LgjCiPxgn6MjkBzTUQUodXVstP9g8CinXW+80YtR5FWlAGDxu0yOI07Fk
rmLN9qwx0nUIFpvyDs+14KVGjFQvWvCekSPT/FUfsuiRCdWipOg/DFFaclj9vqTG
OUkHg56fefK/IGq10Jg8UPSFY0pUT2qwM33qmjwnPyovSxuhxAvFey75bbVDJJRC
/N0tou6wNWdRIkh2rKjmdy6YDQu2tWBcDcsu75oZy5vYAaCFlMsRHvV5LRSJQ2lF
9CBe3Ixz5IM3ipJym4C1tW7xeXd3kXYemyPl+w4JgjmhAGmym+L6806B8JGJDk1G
7U0rbXPDIwZ53pX1R5mkGocY7neJefmCTVzThrbVkFnrNqjXTrH7Lx4vy2GMhCS+
iNSOsw6KxjrhjkSUkDYn9Jv6OVvTCZxqfsA3sr2scgjj5Cw2zBcyMVRS+xdquvsa
FA2o0itIO05s99SZ85goC3o0+45Cr7X4TbkkCf0+H9+pTTIEEXARjbamvebQF6pU
oyQA6Ku9WScTRfypq/KXTBaobLaiV/VnKzDf8UerSZm4np6HxRz74ysp7LZEsKbK
Rbns2cx2xEQvrXK0KjPfHDeCPgK9jZXip300yo7sMwbf5WmFZuSy6L42H4VPhxAA
sfBGEzCkF/AN4ZNovqfCsPV5YYcErzbVS0nx2DeAlTTpjveTw7+8Moiu9cyMrljW
OCw3X8QS7IhDHiWg1yyDx/qsfaMV4CVcqaWKDG5fmUYWXFoy214ncVgILOMNjMj6
tXSIbE/uBmgE/DpBtkFQ/fmh0lNmiK3v45HLNXAoAkSvqEWS9A2nUeMenWJ1htxL
nWyHKCaYsHVBbhdPS2oftc996G4vNAgjkDOM7MKTnjYopL4/oUyfzITZdyhif24s
rjReTq8HzHylzHX1IVsktg7nQUlUPq28BSjGnvN5Bd7POqS/+P1jhuM8s7b5ywlJ
3k/h+W8Mzz6WWMZ3KXyK/HCse3lU+qHGWgWQ1U56UQ8luF9RnpDP7o4zmlC3Tu0c
pAjymLI+c3FKYTxBH6efPZ6io6fMD+ytgyjNxugt2lXpZJYKmXDL9Ldh/0tfOAOv
lkz9Y8X/5wNxh/J0VDx6ayM/t/w4uxBxthInbsODckeJKshThgtK+ydNK2e6toVq
UHUEgO/qTNrhzloNpAPOiTpMoGpCroMixA0jibGCB4ZmsdsNh+kYx8Gds/VsA3k+
+rvbIkhWtAZHbZ+2nsR8UB7VnTM4m4PpZENDzuy02msLjt5UlLq5lgXAY+IRpqSW
S+u3Loi8oESvZEBXs53avYz0lZ74wv6QmB9uC4hM9nQSyCobRwUCATxUH3QG0iuy
0uzwg1yYvoNyLveZtQyRGQLT50vIBido6FgiRovou6Lf6vZqMlJaDmaMOcZup9NZ
y83/BFVOTaHZokFtM0ThV+xscAdLLP5j5XJD0Goxawfkd06MpzknHcRW0zqkgbfj
VmgA5XHufywKmykUpegN1PuMUeoAfMYcTdGDuSQqUtd91KYaqb/B5ARuO5xAn0m+
WVAEZftNHaLWcVd8dWJzvbzkjtPjsu8O058K/ZqCEHi/QAL9vBFBdEx09QwewPPo
D6VojpTQOr5xyQTpbje+WAMa+Bqbi6EqVgNrdqGjcbpPXTWbGYZi9HsPUUcNrmll
4jX1oyPPKGMYs8WFGeXR7ftZ2UIWdGF1PN+P+7Ahkdi5TgvySMRLVNz9EpejAjCq
ToUAatxP4otNnZqQqTCfJny4UkcGL4qtTGY6FIZQB+euwQZEUhMq34HJjhKJMm2X
LyWOwkf0Ps0FQUtG3iclRqc+V9Gs8A5kN89cjS5+OPePhz1IVIgQIDg4K5bXz9ia
QHUldLkcB227DpqFuihrpOTv9ZxrlgaCaAvibuEUIv6cin63hSW2tMLnpUKulkK3
8Ch0Epdt9uJhn1EgnNONhOn7H8k1Iwqq4/kCAZP98eg05LWNYBSHLup58i3uGfeU
vtMpdq/PSAob5hVy7V/JkGNj6gPauY4Q/Bj+zTG4EMGF95bq0e+jfA2eoyxLvECN
ygb4Til0vyJw1uD5cyYZ+iKfV2QYKVDDJZx601H9Z6RXngO3JJVSQJRz9AUr4+i/
JHAFgZ14UiWV2TBfFLXOgr1Nepf2sMegKa5lYhn209RHwfgc/3A33keEfbY+YZWi
7s0n7DMTQUfqoyDhyWVgtqn9ElARD2NoVnsXg4Jzy8e8YSGBb+rIfnjmia0yPK8F
5xMBXDXle97NhiYk3TuWzh76tH3gQKcFbXRhapMZEe3rSqe8GL3rQDI+6RFQYbOM
eBX63Jq8HV9IHvqyol9kokOzi8xi0mnE2k1WVBxUzSpVX/X8J3ECKd9+9ZaBkYOh
oWdlXDEI3SU6HlHEIAQo2pR2UynCyF9kyljm7r8v3+zpUXgTVBHoOCmPfr4/KJCn
wT4lOtbBA5ovzRK7PmJnhiuafJDfKk0qNoiZV6+umkzde8oZ8TRuL/x2gUNLtarr
ZgRi9cm0lhBek9I6r8p9MZ7iqrUbh4Prwc/BJfZ9hm5AKPmRzefgGEpF+24OBqKv
8JL5fdqDoS1+4iruUoP8qS775wiyrrDfHy9sy1ou7v2WdSCRZCKmfhCsyvYYDaVf
Z3yxH9mW+IjDtoEfdG5ucI50tiiizj4pkCyqVfz0b9PdK3HQthTCcZ1gEsXhjfwa
g+jOAztkT3yMRoZWfkTtSyam9S8+GtBN9/jxh4KaC1XuNOnhFD1cFgjv+LqF69oJ
Wbc4ZC3vGaKGFpFzgEXCdiDfyPJ2Jitvgz6uDe50mze7i9ImYVCrBOPsHSWWJGDl
4e5zfMhnMxEqC9g4MvTrwLxI5y8CPFgZHxrzIUYfctKUU/SvBdKaLMX8zbDp2zVT
4wyU/+JqKNud5RRA7vRx0wQI0PtaI2QOWdCqaLbATPBdeqq1/Fe9xTon8Y3qrnGg
I/touV3xYq/u6qlTZ+7wtddiNm3GQ7OSrjpXt1SrmW5JenJ9eIn9u9iiX4+1KCKo
YwIr1tZyRBFSVfAOfk5cm3G5i+ql/37IvB96bq+93MElB1/Q1GfLlBlTjVfOJkKy
eRF3LHVV+dighTvK4Wok8owkz11E0c3W6z4QStlH0TYljBM+Hoq7XaeJ+Aug+jux
dSqDrT1aUro11Zv89MJv+4MC4RQnb03Owh5PdjDMrC0tbiXshBNXYoYIU1K7ya5y
m3wsJTjVbeID1TRJU+7rap2yFX7tCWZl9/nCqM03d+1EYaYC8kyHJ9ToU6OcYiFL
kmrSHuTqHdrPlKmxSk/02p15r+lDSAXtdsneQqHedsTA1XiDWmCYRo6N4yIPpIBq
7GPcM04BMOGIav8L+z+BbgEJpp2L778B90FA9bI6MfdDIIioYTVKuZVSrqXZay/V
cu4YnrsD1FPcs5a5z6EpwY6LQLQwgxEgWtC8WJ5l8Fnk7IdzPZLifo/dIm4tH6tX
Xe10dLgaYxCxY5nYUH6RPp4lE0+6NS4Xa6l8pVVa0QwZHSOqXeG83rXiuw41BxN9
opv4roqfVyuTzYmb1ORjjV9CGuwXCNjnfxUVU6zbunriilcBvbCBuawE9Dnld+lT
PiYvCFsXPf5GDa4iPxLFfvWPGS8N31G/SawLW9O1F8AJKkG01I+C/NhKFvGuBNvh
ehWIGMdJRXjHgT4Cdv/84+cDtablJPnU9eBmzhmb9NCEdX4MYWuBRgyMFHLF3t6g
viX23phcK62wMYToCDUJh3lpv+Y73Wy6CLRnOZkEhmjzP4HrRGmDtWBYFwbx8MDb
OMNCBT08slQzudZOSn8w+1qqV4EYLLK6BuoiPg344epnF23iuwwgpI79UZhjtSjt
SHvyw2FxxOaTgemlUzxgAWiuAPKnrB/tysTdBopcLtBu8x3YGwwdux++sWTROLFx
9qQr3np8y/S/CYYbgieNI7nuoIVcDigAfDpzhx4O/TvaGVL8RAifx1Lu6U5rBs/e
6ScHeXI3LXJJdnsnFJBzXTL24waffqPm09d/AMRRNyph1lHCW+1MJl2T8MvosJhC
8PAStUd+UpYObhXeFdSGJVB6LbZLoTbp4l2pVW1+fCFXjcryvayUoF8u7Vo0h1fg
QfGYF/WelNEmE+PlGxvntvRBGIjWJi5MVyp26qsvg9j7M2AAaLYssdWj6b6Bl02S
VUbGWeSDHKhOahDoCEmwd7uiQD9jv5PEAOvbuzSbyfEWqPMAap+y49ynO7APHFtn
YwujpxUx3dQkfDjsBJCSkM39YbEf9b59UZGkAukEZNWTAgSjNroFfijU4XzulsaB
XqV/LBLhhml8f9+7l1YHS2qjy2itfz4JcW/IyyPZMQGU8sYGa4jSK7UTTDgrjDIN
gzJB7QucQVcPksR/pSg5IkCtQ666LPYfBZYQkCDvg2lMTJkOQt5bDm9+oJNwEeK1
NidSFHDaQMrJiPv+7bKi6er56t8cwczcXRjh2Kr76+uM8TUo7hdeAJMoapOmy+mC
3ml5xsHuldbOdEZ1Q4u/im3y3VhIUsAYWSjtDDhg/dZZPLWGId762NnHh5fSjQJP
r2vvIXdJ9rLmYLwv6vACmirmAg4Ndq/3TgBF3Y224xh7iMSP5L3Inc3UtbO123o9
Ln/o8o5OKBxZJOxjxE2ml7M1kQtz51YkRFZdLRYG0/bQsQaSJ7tPrkynxZBB6CBX
xcFfSmFme/OLnXlI7XxS8CWSHccx9V5WgQZeCjRWJp/IaE8i5e8u2s23x5jHxaOZ
eD2wl1OQMh+KDBdRDOHbM3zkNeILUkL/tUqiWKif4ckmI2miM4oMd/C4SXYrWx8R
FAc5aszux/ycAhI8yiilMqhxA6ucWWfN+2Qu4PZS9Qycui66Detfg7glHSCn4HSL
tmQqiCWArpDvQ1iDdARmJQ4Pfdr5nb+lbR1NLf4wVLefK/UWxpSkDk5CFPrIOwwi
4bhvjotGko/VcCUcGUHC/5sG9XXq6P54ZatYNIb1QtWDkopvk047F30aUaZV3/uk
a19ILVyCfAcRDte5cdkwcJTPxUW8AOiBSGu8TfOwhUb6Ri3rxVvILOf/n0pCLnad
UJPVI5lZrEpakw5hBqNNU6gyFZlK6jJywVNuHzCNNGsIWDJcDJcHIJcedTB9Dnhk
n7QMaRdJ/Th4YvYuIV1s1myMRvRo2+hP0EKMtAOBuiaWU+ssvjtSf9rOjXNo4EkJ
rubSzVQJVv1uL+epesCIMiz7ue1seE1tx2nY7+Sr9SQlM6Qdhx5Es7qfDoup4oiK
lmG93/PBWQnRd0X57rax/Uot8eI2Ag9eSgDl38BCKHd86EmWomLSU1I62R1ZKB+l
ay0ktbOagQQEjceQp60EzbdxCKLh5JAhhTXXR/jCzV+AxFM8BaeK80YzxNrrXLZ2
j5Q7Rznaaoo97naMz61dhClkqSwiVPUz6KWqs6jpPmDQXrxIo5reCtfsIFdWYMEk
MlVsRXWayOJZyjyJiQsEBmWePRN3HVlLMR1L0Oq7aYlZOCYQCiBnn6p4CbSk5waf
qFlu5VQp4nRhAqROGMoLVHqTlSPtPGnO3oEZ4ssgR6liDpI8nNxCwGUem/5o6IaT
m5yagIYkeGbdenDYPg0Tf+M4B7ZIpYwcbDPe3EIaox6jHaYPefMZm9YxftajmIDM
8hD7PPoUMXEI3kk2tHCRcZvUu/qA5x0joS1Dl1moR/sLpBLvtX+/2cIJ+J8Ihh6W
SBo59/umiu5RBSabG1Vi2kAsQK+4vw2Zxl/Mf06Wc7TBma/pqDirDRyoqnn4t4CT
zUGgMmo0kxCn0PP6K+XVGtivImisgy93NiVgcfYbqDc7GoDSvjdhstquqPlTvTLs
8Xb6VtSgN8jjZz/VmBwI5LOIBPMuDzEzJubR8FmHY4EFcnDb/V006LcNI64mPMc7
XZjffa9/hZxBelfFxRzXb+lXOUHJZBYimEQuTro0DpnLXhgzmjfih8JNjDK1EYkO
XWUtlWZTJGY+svnL0GvhPRkHydZ+UTKbV219Pp/1Kq5MyAkzX1fPWwi15fm0TWAq
766xGbi8KwNHUWbBo0zt00/jOxlLU2Y8DCMLKy1G/9n+4F9Duj9DxlDbimqqIXOT
WFk0tJhbRKSLC6Hc6OutBwyVYCEarL9zTIyeggEiZWp7iXLFFbAsytH2tOTP5uTH
Vq8LnmcZ9Mw9FSvcuHdicrkyxfDdH1ajph33p0c+ZEvZim9UCWT4Rk6bTuvJ3b6G
boBGeGND+a9DNTpdGGItOSOmfqX3IDW+Rp8Xm6NcoQpgBhMd48v9Aoe/kEv8NTkX
OxVEYB3yFmF9lq1DFo0f+6i9nHeAkbkYUd+03PTxm8mj+RUMNCscPNy44YzFJbOt
2EKdJ1Y/eMtmqmkeF9Gg4YC1jALeXoQBzhg/QSEIpBElpv5jbeXiWomjfahfz65I
xxgmwECoaZlWBqApv6sjaO7Rym3MrF4o7kQYwSjYLOVBvs3Z7IGQue1RrGqodZHV
M3Scw/4ADqAZcAvx+xkKmkuBs7ZtgiuCEMD/m6DpFFTiT6gZrTVl4h6WUzXIe97H
W2eNjzPZVZWlyvvIqKkrlpvB11YUJIqo9x5s0J/EX+X4xCTMZc2UpO4SEX8Buysw
nmfGUl0ERDifT06m/e5DxvCuForINV7jtCk1XKG1OQtPGdcZjigOnJnSsuJpGWuA
2JtNrYa+X/3G5vl78X0UQ8DsI66xJv/zF9yWGRX6mMXyfUI9tkobkKHtDa1EzQea
gFDOjWy6hrStCE0GUWtkgW5ebYxjVtVr3y34uk9HXFiehxFVi5NefOYSznrDRuLH
gjO2c/89ffn9ORSrrTZrd/CiWX5ZX8It70tN6QvO34BknRv3I8V4sg1WaFZ1HSUV
J1NeAX+J7Cd35nD8FNiwEYgMVmRh4MUV9u5/FB8y2FW1LoaYSg/Jth6fsR0g0GFO
IFLRgy+rl8KvlYG5m8lCx9RTQ/I8C6iRyMTHDeZJwsjUw5UJumKznZ9eLfkt5mo6
BQvpaHihLxevD5ppqun8q8itMadHxsJtDzeuHElEoYgKVUwuJVup3nqNZ9KSk41O
loAv0QQ80YI5+2oQc33mKEj2KWe2ZffNLJ/osVxeIEw6FB1/gu1TCrbWsblYeiQK
7LRLM7db98RDL+KF0Jv14rfEuO14H8Hnj+Ven9jvX71pnk9NzkOQrCIOpimGieix
+2SOHHVZCVMdbeI9A/rcxR206hyp7lyF8NyoN4VI7Vq1k4AmKWJ/lfD15Adrc6g/
iWn+TipBzDWGJjccwdhbHnRKqnUuYxOEpXi/KbgSyL1o/XcArW2VeYazQUfk4+n6
1TOdKvY6gJOu0Mh4j8rQ8gvH6KpMe3e0pEptUq9EFAkMYvihZgXmcdbC2uIr8ovB
5gwZiz6gjxalIv8mpe7PUamCRL/vX9s/KsQcq4esavB8Jy13ovsC/tRG2MqiKhMt
SECAedSranWoOgJKodMZXFZQwYzL2ujNeCkdAuSt3pJqS+rfQgAFuZPHTJOuQFH4
F3Z34rKrSln3dUBPdNQUE5mNo8N55PAS9wu77l+DZqrW9neMQT0gjPO+XOJGVeLS
6KEKRE/R5L7hIM1Xh29zEz1RtCDjFxU51oYyRKI9xTS7g0i2scTxqLV/SrpuvkPW
WYz8n4YSxph6CrGSIzVTj2MW39XQOCJRx3J4qXkFqsWVqjh2eiaThXwtH2Sdzu0t
2bZVN/D3ZpNGvkgY4SljYsBJ1ko0vLQLbykcKVQzCJRVirdZ20Sum+3ET6LmWEXy
5N8utRMCNVgwG3ZcLUw/N0+rTz3hfZvsI7CMDbaa3sgPGwmU4bXoOeKY5oC5lYjf
711tZ+TIx8fMb9mOML52FvNfHKlT23WhoJJMadyHGbEM8qO5W+IDBW4kVsLdeBte
Y4U03l1Sv6LAMDNeXi8w49491btSzlLA94YQXK+W3j0XHr8JExz5bP9rctMRI43f
zHojQXzbcn2gat92i/uoye5qFZz/9Swqe3dVOVx/QhTdbVeVhrp9zR3sBsE2mK7e
DfBJCHk9WJKXeT1LrY2+VC4IbXz7bV1CA+m46SfSFSGZrzNZZ3jWAq8jq0vAw07D
Oh3rlwGxkz/Xok4hneajdkuuq5xKodRL1JWywuA2BezoMB4TfzBEY7d47W3HFMt+
YI48oH3N+4ZE0kcluxpZnxQTB/IQJhdIYhgWPwDv3KU4/SkNH1Z6h8L9KS8b527f
VpgfmoYNf/0zu9ej9eaxlKr0q2pKqSIDiEm2fVPRk1cF/DvRvy/b9pQWK76KfacZ
qOc++hRtAETrgG+qqeapckBJ0rdkKfqnoqp/h85lXTw1spzIwd8wzok9LSqKzvKJ
GbKXiUAQpUj0kKnSw1FHCQ7hBJdxZbLlc3gtZvkAaSOwpwf7XoJcbhv06KtkM7dU
1aP2NujqKNaG+ORr7Z9BXckZRYJZwSmR6k+1xkeKbRdP1/ubZLoE3DvlKsc6ROJv
t2j6fmbKqCzSzR6OWSp9cuy/MFt98Todg3ehVRsHwd+VnUm81/tu6GJSAI95Ecp/
Gn3OzG5FHdeBXeQWCsYQjcjzT3cCtb9BdDxBif06ZITwUmu4HEoBvQ2Lnd4HFZvg
nibe84n5UOShrJitNUqr2yHlHoEuaNgMU5F/wrSbbWgjnxnAO/k9v36b5frWU27u
OnzQizwZqxwIXV3e2Wjf/0CxQcAM6IDisDVHYjown3UaEEAEev6JLYx6FORcN85L
UtOeN1HKijq11DLzGQBWkzL51g7+6Rbna5cdm+IUFZ6LUFJC3AewRKBsiHcfJvKK
FiF7zEBeZhaU+NByzdZEHHEWLtzWvPJRwlvQN9Kfupad8RW0G94SCanbeWqMXlPK
5cRoownimSH7Ty+k9TC+KY1OtD/UZZwexzwxBgUNxGbC9GUl+3z/hYCJM/D1z+Ez
3e4r1h8HLVOz9IGE0AEEnvx/m44Ti3Pzwca9UVKhQyjZtEELS5EnBWEPjUpinsTs
n6UWizL2tLLyvlyxRZ4E7Fe11xEHi6atgZo1bKj80pSQht3++8YskJXVlnlf+G4H
5RIYJya6lUAxUTWlYw6dMui9ortpUG9uurcCK2YOn8c1yXuQ3KRnsMgo/3K137Sv
2UTYkO52tpljm0qy19N5qIwaqaceyxOo88B3wBbPF/HTPtavuYhACEnb4iWFvdls
jct93YC5P0EQm/HajxchXzo0+oI4xugIr+8jpl139WXpE2NHfLYIWPYlerua+U51
QvvnTV2Dqmzap+umSxu4IJHgBHDW2GVBMZoSbDSzkuj2GxZwCitIbwq+ZculsVEU
1lYP5LHnLU9vU8t+2GU0tjL2LpipPFxRHtlryxkhqKTwrtaSNjhMlFg/ZXDY2yLe
3Dj3Ky7Y5zu51LYtCjCiXOsaJt8yICDFD+pw6HmetnC2JU95hoEgyHFQgO9dRlEg
H6SYvPJnMZ3CVI0jrbLnbSHm6ezxRdzE70qdLAZxFhdoQWVJ7WFsABf/k1KVpW39
ANm4XG4MOk4SWA7eIPc2ZARPfvgf0YbLMdkYAey2iMsSz3j3GnwtkLsyZwt4q7/+
r7ErdkBOnU29CDQHjF7hQy4tqXNMkzBWe6iiQR7Ptf6mHb7ZV0/8VVV4uzOTED8+
4y9TXxd8dRw2CxxR7jUEs5TjF8K4FwuMPYwNJ+U9JEebV01dQqFE8BhWDrQNEWd1
Dv3XATq/kJZboIS0C5gLBlLpnnceRDmCdvocs0FnTSyHn+cESZPLBhRYTmxDVg1r
wOcsZrTTHG6dKelCmA5776eK1RTdq/NK8jkqbvkEkzMBdAELhSH/2P6E9uZicSZJ
4MsMKuH8tTx7xxM1Jp6hoj1Ip9aEaYvdyxOXd3e5BUeRDjcygOI+kKs06mX9Xtpg
SNsiy87DF0h9s/5BbG0ifeyVxS0jPrWBE9Xiflnv74bWVgaDoUDNy8ZyT9h4dQWG
q9mlpPOd4bbOmvk3qWghWncvMhqMIS/BrjHDrvx9FmsDP8InykQBiMvS/cFGzbK+
bQGezaixbtgxYAhG8Jh+yoxBqBpWAbsyi4UDdKdO70Z5k4WY8khG5ykdbOCETCrr
peclQ2oVAIorfc1qhQ3n1QLa+UcfGQXsvWh/I/L5Ih6//PpVZDXRlQ/kQ0SsqJYW
YaxKiPnTc1SUilgDJHGH/8KmrDDb9Wqa0fm2q2yE/hDMuiKlscIuGfXWPU4HMXR2
8WPsnQEMRa1Cirf6FUv46DCI+mOAxYQtC1ig0n5UmhSlFJs/JAg9zE0e6w6PVl2Z
FqEB+P+kTOfTGGabqXfL+1yNAUNajMPig0jnQ4S6pE0x82HgYtElTaUszUZ8w+PE
T5dTqHvUO2NPvAGfNnrKlbQpXWkH6eoV4jSg+YnAt3y9hi3E11OYuAFECLch+jMU
In3We8RGBKsF5mT9vmTiElaKsb05kHK4JOrytBNkbXE17wJ2gNJWcNYMj99raVrm
GzpmWpIrGzU1nTE50K6VZyvnhBeE0Ei2QoD3J8PSpbcutJcPrXDvwYP7PG2OUX5X
n6acP1jAhPzN34YRX8gx2W1C56R+glKmmn7EQKnASrm3p6YTlkaVZC58up3vd4wF
h8TR58u0oe9FjEmXxf7xiuxW+x0mIT9T/vLirEFAkaOWXSJoXZbhgul58TeBIpTq
/D33BtAR/GDeIAatktwG6SpBu6A+S9MnI8YOi95FFDxVW73xfPgZi40vY9jLa1Rb
DPd+eGFfq6QZL3Wz0S0YFly61A689rHq6/ugiXLDt3S33VS6ke1ttFzU5TylXp/u
nXMBX9hvpdRRiU6Hqk4Zhc2fogIisHW0vsVmEPubdHyddc9ZgsjjGEsj4fTw+Hpz
butUyvTRnAcPQot06v2VqeINAb4vc9Ej13CVVmNxD19UO5EiysYw1viy7jAo3cOq
T4ttzcsf4JK/3dGzgaCX+jPYc7sxvOWZ+ND67pu1rrfWFr7fJ9yIgH0wrPrZm/zB
caK1WUVSzvruJi6xhugsPDNDTBKAZ2TB5y2HVOREE0uhs6+g9D30uqWYGySg77M2
T95T6utQIf9M1epkK9AatHajgg+JCS67NqAeS2f891U6HJeucUqbXTZAsCexg8QD
SBiJWwdoDn9aFwtp2shQap2Iq6+NCrjkX7oB9pm7rcoOwHlR0wFx0hE2evvVhB4c
IpRG0jX2IeziVekOf5koGHm9XEY9gjVMaAgJfzW2Z+TIEzn4g4UKrnAdsxj8+tSc
3ckgq6AYihDFir7IVMRb3fZOWw/8HWKKuO6ndUMCv9uyaWObM7DBK/kse7TrWsfG
0ynmmuEGMHivfLY2t+1r0h3WYi4EmmAvSG2KoPcax2gzKfEgmqYcGbgQMDCsApq+
JHwvFvfXPytkznUYTDbfu+cWlNdQzKB6HNZTue+ECkjQgFlFjGWjjBxfA8B4u/ov
ekUmFYrVHCvSjBzVdAOL43ng9iR8kTJDnz73YQ7v5DbjYtY8+qGzlKTFz8NFYU89
dkpFWNQXCyS7lPWiXZvD2P6PNdH6sQZtp9+NzY/UK4/HlwWHAHmoH3pVf/JQ3BXx
BxLEQVIEFzaPE9R8L0wHScVWKRwFMZX3tpgd3i0Z3qVoQBRy7mUBbMRMZOxSz/Cb
NEjGXuUP2aMWbgRxKttmw2eIzNlIAD/CHJiTauy91395Mjrmk/ZLdflbGzggBcOo
3O3CsDw42mAmuZCqzxmSA8mL5JFlkxQTe+tqIyqTGQiV5XoKQWHCmz6dGAiED4Nn
thRVA26EJQz+Vv7kqXKjC2Jt6leDbaUEmv26OqEqMfXGdDILZR27RsjXsJdHJCil
p/M+m7o9RUekJpuPUcj1fmLONkZbr587DJvMQKLTRJ9cgrTHcf8eLqZ029zkZ1VS
rrFJo3y36DFe21kWoGtBX+1LA2twzXN9GaG1IbLJup1jeTc02If6hsmuN3jOUAwD
b4q6ZLFfEqpewFLKeFP/hpLZOjrcMRzgOMZDYDPJr2+cE/3r+V3PAh1GFebqZGXW
STMtoOt0RN4NOmDTsuagA5jXSw1l+YYahl4Se27iOHHuqRTW7qtd+mXzibZZRmoO
kNG2zMuLf8K1KYR75yEOLyA0EgUz4616sltJvrWnOyxMRKo1IDtymRA+FBnzgQAT
4jNRd2k28fUmI1LIpri7KFLj/jqHbVLmEIo/E1i7+wTjVlICgssqdxiB4+KLcdI4
2kiD7zaGdVpCVGEqjA0ioFANu2gdRugZRUk2eA+eQRt7mez6gDndwdLyR69GiZNk
F6jajhx7QLdCJQSAhELUARea0FkCwLH4zqCiLI5kIO9BHxaOjnM3ZaRSoQO4dwAJ
KsEQhoypmRIca4PvSCchV3STvcKC0BHrzEx7ysQPRcvi2xpon4y1rEahMlJZ44fT
SGeZBumetkfzqh41dAP/K8xL9esf0cweKPwUsmGqz4ke2I2mC+KNH67VL87Z3iWS
NYqN5q6Una8U370FA+OqGDYv12QMZO9FkCZdfEVWn0p+o1gmiK9REIUzXOrxlfgJ
W39N3GH4Gbq2eYWe4KlITzrNPWayhd+OR8H5BbKCnOOHqlf7NbZA16AaguDM3eMz
76OKc2ati1dq+vee8EiWrLwzqr19O9lg4A1SHcZvO+n7Rp/1bB875oO+lotU62Os
czwn8yybK2Shk/DoN+iyZcMyonETTjuB4BjyFuJLWIdd3CtDb+9y/TdEtRcfVcSX
Xh+hdPmgX7e5VEtfFKC3lvah3W9ItQdBX3gHhJ20npCrqQs5FO6c6mWryztSGkKe
3HUeLNQxtqIkjQarcgsiojCW4AwAQDQpJmlhlFbtMW+2JHYiLcXZJj39YFi648VO
a8im2lZNv9ROBZWvNA9B8hd9wq1IMtC11KxVfXOVpBFZbAdb7a6gfHhBKCr8Qh49
P08UplTxIm+q3gZvrxR40PswJgP+ldR69ajHWrVqHtCnR2bbhke54ojkUbvEIKz3
+O719OiP5z704S5OFBeDZzys0DYVgA8xZI7cX7G4g8+14oaM4VV9PA91ChUElGNA
80gprUv4YvvWQP9no3JIZQ8qJ2InXFkoHER4tjnXuhP6P2YZjsi9LJIG8z7mMwXG
rqG6WHdrJPkKwn/liUt2HorJrXwU4cscmkLM5s5k8qJCy5cZYQUi0hpv6GnXrusW
OxUWXWq+3PGLhjHOUudyQ6QjNVpA7mLwn/xdvk7uKLsds/x6FR6jZI+lNHg+dI7p
+tMmZQ+cHR0nP3xGkHV7tEMzBGcI5oWsuor3AbYSJ7FljuFkT1+/BwjSLmE1KLHk
xH3zy5FHlzT5D9kebjcHjJ3BXhBS8V/ByyN9lPcinrXEPTVIWU8errf9Oo1NJ6lX
KpXod7W6lA49BG/VrhNPt0JYzyqIqTMSKGdvMBaEnw7MF713m+U71u0FZgk482uf
L/+6hvEzkGwzoUBnbW8crSTKybttHEq2m93GjO+H+a6Vub0I/u0sI7lFrv12O5rV
EsyrsksSyVkyjw1vEUDqFUnYkX5t8vq9mPHx6XiWYE50UUZd4vU+qq/fGZwkcrol
ffp+4ExOh1W805V+69ziw4EsdNrbsYcngvWxJKBw24uF1ZAP0HmE2FTNXpx3E3n1
8yI7uiVFPeX7UgAvB7xvVFOHIWvV0UMyka5Kf0tH3MkxjFtSO/wfRfDC31wAQkrZ
CI9P46VE5uODX7/hd4+KXutIaTLt6ZIVIn5d/DmaHn3FkrUHic8dOvuJetSC/x0y
JFnqJcJ0O3f3U4CE6dAzlp3px0Z6VRZ8EPjiyZmY3143DtBNsu5IAs8U4mWThlkV
y5Cawq/AIwfhzpi0J6dXUYkLEmEoFR1zIdiXYjmOq+EeQ/I2WpkV0cFe9j4jXQfV
UQ2Bhl7SokJPZMLI8IX4C/2kp+ySMaeEqB0s9sahbdJ6wmfgOA7oZycvwVbSUge9
q3fP+K0xq/Ir+O7m9qohYxzB0x8Gt2gNoOMOUsssg8CgNYUjdf1npjlw2UEpg7JN
KAgb491Y8EqDKa0pR6kTGentleeDacbeWotj877et8/Ln4qgmtMOoFO8b1tgg3mT
2j/+LhKDlh9bOq9X2vZueuCLtqr3hqctqSL59yQecbUoxURkE/L8NGtHOwqv1TRk
1x6vm08mhcgaIW5OSmaiUf8pc79AyFfCDNPSKG0JcZnZBuLWjcW/xI+B8WNGg97r
GIK5wcADJ9UwGdVW6+LUu/Pj4Mi5LLiigj8hkwgDGgvf3ZQJsHhuyZKW6LmyKZ7o
bPNKT35qmjKmRB0EkD4T/Wwr1B3MLoowm8ebaT0JeLBiw3AbMqH+SRZBXC+U8JHn
OS0HBtO2WleHFeI7/CSuNwQ2Jf/djFSu7QNduxzk+TF8k8WbMbW3gH8lT9HZRf41
FKoUFzGZxyOpeAMaQkpIxLcS6qJ0kjwhyPhjx6Vw1hFxb67P1wu0RS7vA88939YP
7WityvF5qXktL16+0/AUdDb9+kCnf7LwkK4085ye45FMZAazjl/5yiAbuNGMoFrf
g6rA/wZeNi951mNwuwDw8OY/K7yozJbL5tuS6JQ3AMT3RAHb5Vd6/QmOjUhnF2IS
DFPYxPuoFPJMCEBPJBrhBPWAhWs3XAtP7eLGuFM3+PhdeYljueGBqsdUDjnw/v2V
89jYWI3MuGFWujx2Hom9+B5tMXPtXCVxQgNljwligOWNQLazAVArL5S9Ja2PzoP8
YxKMA76aHNUGK3N/MhG7hPxicGhFugRR5UPinSpFplJj6o/7DH9szgi4iUTjJ87i
c7rEomNg1nPNr7n+Zq/c345kL2NBL8uQe2p+9wm1r1MOvMRq2xcTXE25XWI07fdR
lJVbvqg1cAtIJBLMg7fwU3KMsscP5QbmRGW8sho8QRcU3YfTuxID0cEbdD8sOB8R
PWBDELVvpZaPVpsyJZp41C1BEl4LCi6BmCicSqpSLRuHfEvPLlSop294oys5zdix
iIXNHqwqxi5ALFdrPIWUZefcJT6wjbJvaUL/DtkNDd5EqgJ62EuDupa5Cdypgrjo
nNrCbqOivBX88biFQ6/92LgWUMyLLTWalY1yjowknZ19N0FV7+URv7wTC1YGwkwK
3+R3kf1/dD5nz2caMD7X0/5l/dpfCa21n0e+c5GBK1esSXnMvomjdbbJSUNfdDCY
j9uXZyqTL0Gp0nTkKTqFwftLD/ASSYzsQ/wdxTefnKPHuAgvbgeShM2IHYTDCW+T
24HO/UpNgkaSUl9xPrXRH3UqsRc2YfDL6pZUaxyfemiZdgMCgUgtEmw2rW1a8M56
HOqMcU/Sm1HElsdU6qiF+0xlefQjZbyRh57cEVUC3wZpRJqy7cCjWwH0TROzQdPf
7DzRAbc5Z+0Kh9u9IcaT6uPb9YPiAyXQgo76K+LJGQVl0NigO8Bj5Ggx5cTEsTba
+G211pg3eugsFnO5owI//tRWYsvJAGzT5movmeOFs6TWJgDgpPvv6DAtF0A32Ieq
RERKqap4Ld8f7EZsCgHY1HCPP84p9tgSOggD7GHNw6Z0pKW4E7F3uCC57ct2M+MH
xLjUSj5nDe+YaQ0NBljJ+rZ6Qp3heOidd9gsZjgFtmpl8ssbvfW547ONVFdy8Fna
xADaZywzxWPmiX0Y3LJ0cD66xMtO4CIFBvNUa66sswGFKbfttbsDtztpzBaNViBv
kanUlHRt2OXn1FWKQbEibAZK1XKnjq2qA8ujiWl01TL/FORQYBZGZW+pW/lAb8IR
9UlTmV7JhmT+AmuruZRmhIYJhMScjCNI+NnAl5LMLeUS4+YiB5rmN77zhOWS+aLK
LNf1P11EyA30p2XmZlfcrxxCK66+5gQz7mb3TiQddXZ45n/W9rG4RxFQe2vhEe0C
xjaVK0aNQcN0bwzJD6p3qW1DYuFDcAJ3flXqmHnHTdUMlzEgyc74C280ECThNDKf
xDZDwjIBVY9gJ5bh5k9a0zAtyq9KB4Gk6dNirqrr2Px0nX/bb+hPWiXYHUre3rfM
xg9zJYhHsJty/zw+Eh7UGXsNxmaoljxV7EqHzDZ0JXZfrYGYMXEEm7sq3bUezxyi
/ch9M9+Rd9mn6eAq2pCF7cpAO292p6mIYvdjYWOyHAr1wBYJINFoxqHxbXfcXM7O
18L9VxsdF5AyjULM1rQHb3NQqPF5wlrgA8Dz6Jyr2CGlD8KszIG4kml1DGCpcX52
1sGFd+ir8zW1+8bh7xZi0nBSlBCEpGnx+a2bxyuKgVCdYJ2Kk/zdKEOFkSdlAI7D
X8/j9RjYxnqgbcoT+Nh1PxdcAHqnrYpFc0lx6oQ6hhCJ5JMSjtmsp+tV9ww8eOn/
hIuaG0YMEDzWR1DMOQnQjJwvuey3gTJSgZSCnPtR5IwpiwjUjP/xhHFNANRwx/po
BWKqabhK54qB5ATbq9ysQ2LOTh6p64hjQCPPyc+3a/S1l7VSz1GDRMZAPhNHxPM/
LI0CVmB27WllROzGtdTpdBrt1d8iD4nry14cZdoY6EP7K70k5JGpfkB9DcC1rI5x
lPV/BGo2+5ifcdlx7tY2Ln0vSqD0d6JQuNc6mk72NcR88XN9b6mJiCGOk1DfZl7K
XVh/KekNoyozpG06H/mIY/q59jLKLX2v41vZpVVm1JiMuZLAQPkVM+jsrKTWWvfi
Ns/2be1z12GhhQoiDg+uvIo6rZlvzwRAyZpxgbeWjr5+CRagovTwLsV2d97vUzHI
YM0P6f4uA1EqbJNgHmX40WOhzCQfMX/xWYbkUit9jaw3SmoYMbVG8pQx4aBYQM4v
kk9PmIokVgGFRCMEWVLbjNkaxPAHvTBZvm15RFcrrKjdtKQ0cU3RO/u/64UtexKb
WCxKuIdkejnycGFcD/c9HXSm+b9I+UHbl3PXbhV93FM+piqHIUZg2pXDTuc/SNiG
sFi50gIPIt+ZZsF2SS6Jbs1Ur2Axgm+9l3HJ/JYb+Y6yMp5mJY8quEnk2X9uT0Gb
VuM2/YPZxx8DLavlAW0S26s5dy/CHwrhdSzGL4Er1Oy+E+R8WDC0dbdSEsw5wzXH
sEt9gAQ1IAR5MMc+SAvWg03THv7/PNCl/y5eke03j6W9uhc20opQZ0SgUQYzuABc
op6GuRoaB7mFCCO+pjuxzfuszMeCDEV1y4XLAyw+YYKgBdi43Tvot4XVjCCNv3Xi
ETqI99vwansfR6xInxslaItoaSpExkCEHufnAH3f/dMQNGtt81l1QFebccfJI25+
Bg/FyaZATWZgBXOqHfCNzfRARKOKKT5wLkSpnswtUOro+CWbsMToBF5pPctBOtFs
L3yP7/wWIkIXxjfXIOIgVAhSkGiA8ZQzjNZoxPY+ZUZKbhpfmMmDFIAdK+LnojAj
Tms8oPACsS+xqSuzPE3AjWfRkkEZ2aRyWxa9YXf84CaiLlznkseBJwdmKiMrkbQp
yi+kVQcXUxW5KqBczLp8hq9wg5ks2ZM/DHhBiFnhTfbSRppODNWOXCYtQkVg0BAn
za7zPPCSwkq6pnffaPUXrHy2UrhP84CfeOnnrJqySdHVXg2GRQAbM0LG+j6NK2ki
54JgxlpUp2gT5Mii5WRZWPlZwbqvwv8e0Xa9sugkfHe2w0iBFbkExX+96C0xrruX
jup1rkA+8z6v0eoYfTkxABnzG9NqBgfqZvyshXCnSVsvG046cwBf6+aIp3DKTiFL
CggNiEtwvZArZIaDdZNCnR4TH3bhRSw9vACKkTDvW/Y9D5Ey6epaUKddSxVdrJr1
E0tCDVzNypeB9N0GF4UYjyBnkK4hsjMyZDuiEttQ052A9fG/VBkZUk2jBfBHXyKQ
t8MLAccf6J+cMMAiOuo3OgpkuAd816xdB/RZwkbEffCOqSjsV99so+8f2cVeuGSQ
Y1Sdht77kyQH9K3hu1B4cd73GrvEXkY7QiWrQwa3YTtIL2ICeB/ewbhnRCbng9Qv
fsbWVmteNtwu6zPM6libsNEhNdI8u91hdoYg6v29V0AIopEwO7ROgJC1dt+Ivq18
sHuXjS2gUGZwCjcyQ204PG0bkEB4SDG5WbbCIvJD/wruodcrO1o7s47SuTzPT6tB
SHndmrmk0mVykEgco1JUvG75KSPcG5SkWOjpVd59V8N06w2lLM27pgfjOghWH+uh
wEAL7bA4rIxH0b+lj5lWCMUcf9z3Jb4CH/Q0I5is0zOoP0vdoZMfLr0vtczJ74zs
+d031tCHkrLMIVu4xnKCZSWN7Mp3g1+bbqgPPcYZsYuDek1OWR1UIpOAb6sn0zeM
EsCtUpQ5TETPfmoXdwV5Z9gmB2fHMg1JV+n+HWizwFHsNBC6zaMSVezf3g0X2JrL
Xwy1ginrOZhYJPkLVf1OUwGhp9tDuZTzyJShN5Rzk5HWyGgo3VoD582lARnnd9Mj
DJjIc/j4PcOp1vTKvLu3GtusiicVTWVQoPsPfzB3DBZDCZgTeJfea43YOrfg7Zht
A03bK8z7Wg+cnlJrFCayFfCZfSs2l/gDcaTQd3VbRZ6QY8B911DFjNqsTjCg4cZV
n7owJX/wqn8dltKdYU8nPpzE/YNKQLMoVWYqJCsEqqw007N0dzuqQjlDkMgVUhJa
Jc1qLQbfrc/OUZkXcyQugdl1hZyUanwpm5gSxPnt5XvTmKHSsoSOSlxkJuvcWJNX
gXiKFMC2Ywp0nf0b9INi2sFBIhTBWA0yUdn11d9PInLSWkojv/NR3ojYQrFwkBV8
PbBesTSsWnw/SLxA+5BwcKg/s0XhhOTmxw01HPgAYGtsYk+hQYMLp8+eq1uMOf0X
ozrsApdipHiXLE4W0Cea0LlURrQ1AbZgNIZCWQ1sVdhV1SkZBTgNJfpZmmUqomsR
1v5hV/RnC5XYGiN3WSl/37NWq4Fi0Qlqc7WfpCh6vB/3sg2+gmrgBhzl9MpMs86l
RP5i5zrhnfRpR2GQAB9MLtuLonMto4fmG+Td/fojkt5IYJ0EHsEKL6H1maAidhry
h7u02Avgv9h61tLI3grdWkDwuDGNDUCV6CzmyEHlkuMOtuZXKZXxC/8ofk0/oiBk
tEVRaYyqLAUIvfhWsZMnYbNQ4emm2aP8JR/nzqxTUa5esTGJEqpghDnK4si65KuX
7h5tNoMFSaLVC0LDLQPnZGVswPZR4PcO63w8dzEyLq/f/+aUvIz1ZKzs75VGA8zQ
/rQwAB/6CidX1wtppWQlPIn7Ur9+h2bYuB5y2SgkCIsxPjRCFa3/VjQnSA4f8P2H
xMduG/9b8htlxd8/5bUgdQqLGfLQ8z6XgMTXSnF7M0CcK9in7TSYprIRS57CWOnj
ukH9qDnSy/9tFrQQSSrdePekRnLfR3v2K+aVXSn/Z8RvgEJulKmS+DY6wLfJUARY
NmpSMSFHYtsvDg6OxL8dRyh5CL0Q5DWesZoBXbCnM+6TLWdX44syk/YW6siIVDDF
AlAMO/vpf7wQy/h8tiWoXBE279WVnqj0KDsxFa5JKih/mqiEiFhrlHbOk1HMtQcN
mGudc75aVi+QSYpF8XQhmvHYWfTdKEoi64EcHhPlvXvWti7rKxt4XPBKuTzJgBuK
1KX0bJfye0dws60ONXOLHIjf1dDbvAtzPck0o4ZkAqwRzpxD5qWiGmLd9PZP1ifb
88kPTLXyy1a09uuCHlI16HzBUlVoY6O+YttS6/Uf0xbJGT/kOF7fGPVC7UXWuJfQ
l7JJ11tQPfPJ3kC9B1FzqFqOFNDQDr/Ky4cpNQ/FGMbtqIvPpJovo64a0FqM0I/m
XQ3f69xs/mp6Svu4h505WZDg0fMsCNF+qN/4bT1z3ZsRC5vpaaZyFukc+4d4nelK
HsnaOnRCY9ydVySI5pWHqFpWhp0Aa2rkwsh2zBQjg3AR5xXejB/zI8qWDuRdtG62
5/i2Y8jwf0N64ltZjQ1EA4F74+NgIcS9SzZaL2tlO6IEZcR5jFQtXpJvQtyXXqG5
x3wVtaYiNg+bgE1Eey5c+AXSXkNbp1hsbzpOyMju+jupMOEoqNmeYLT+YZ13N2zU
0d+gl1mU71R9VpfoNr1gX5Gc7scrvhMHpQ5wYNc9AKDyHBK+8f8XQguX1bRI9jt7
1UQR/2NGEhN27dFkiTFFCRlS/TikTyF/A+C0pwEshJaXM25dTeLVERtiEandFW7c
O0CiE8UTxO6r/0dW9F9gfiWjG1n2Eos1slTo1hMwFXUsoENG281pUuRoo0Qde+gu
eIVvVy270ic//8mZJPNAOutnZkAdgtVzkKmK55on+eIFZV73nF9YRc8Q/PP5TyRt
Xi/ojA/gOyQJ/6i9hu+bUpKTVRQTKwnLcqfbY10mUOWBNFTowfVVeQIDh5bKy/po
5vpHyvoOEsPT/z0AC5AMg8TTTfVze+8m70gM1nvhUb0FTIfmWu5/Fh5yWu4CaBXM
bGcHoYmybDGmeijxs5V8Z7urTuRlixOzT7/F8inRCygjDFO0bZmoxTX3TJplKq+U
WykXScvJldEe+FQV80WfywlcroBxwvaFHfwdP2yrYaxM1cPSH8nPD+S8jb9ssDjY
Re6WhibHo6uQ60DsqK6+hXGb27U78iORBsQZlqg/J+4WG37jO310BaDA+qZc4wJd
rGcAFDfbJIORT1pmDY+vuakOqKshRpeQwGdX97vVULsZYmcFZ+GtLpEqbvFwB7k1
XYDLJX++GAQ88GYu/xrQTRr9R0ACODTZKyuuECdUgPYgQnjEpA0/lNr90pUFIlro
4F0eXwMB6a2vbYGocsTsd2w42e/M9OmFOCOxKcGbiYz6WwvIjdm6fswWkoQmrehV
dAOvXMsKjtXKPiMYNu1tbHiRo5NT5lJUh0HkSfD+Q5BCJUA7nlmyvMwhi5fXl8Vk
HeTYZD/hkmrcPS7UUZJ//pNHWDqF40D762OjR+ShA3DIIK22u/HkznzYUE0f7GDI
+FQEyO1t/8r8Ne95+WVHor4pjlOmMvy+uFoO4G9H6T17IPGEZ2W/7L/ODF8bqtsc
cHkAg70b5rDPqRgrUVGpiJXcQMqIseKxylTvQW9bE+DST62L/ZxiuHVMIXh9byqN
9Ys6wURzBnN4sfqRxQoGa+oSX4TUt1bvcSpn3oeHXB3rY4IdRp/GNmbCDmqsU+AT
Zt0BSNH7Ksn6PP1qZ5yTstEYeuj/FqsS/z16LudGoN0bDBy3UfQpOnzxY7+XbiuA
VcAMuOAp8d111JRPGavmr1hTaq8QKaIo5hULyjeY8ReEDZHcg92V9t+lgbAZFQ59
E6kyLf7qTt3Ns3h+mqlPOGu7yi+dm1M6qjx9nPJV2YmHtlheRlg5Yks8Ndmomcg3
Sv02baBYf7NmGRswa+3hlVZjRDJXtHGqqCE4fUUq+06Bw4Zqsa+jNQc1ykwd2Uqe
zTTrEmS+vpqPcmTVNgPWP21nGzWNlfCAfWkyyIAIf+bHKt5BLM/yP7Dwe1XYpAWJ
CKtsT69ADFg0JsZzxxY3Ue201CeOG9jl1DwOD7kSXFFzQhJ0FLQmohrKVFt3iePH
+DUE9rUmoaV/chf0oeRlQCUVWwmWfzYv+RoEriNOWWTAy8XqhcRAUBCSIzaBbO9e
owEXFiy3V8/cpCkQ6UDVBgjcFikWiuWzs41CPZlge/johs8ZUEbLTPZFsIR4LkEG
JvPWSL8RI0+VZZzcmG3UlMFdWonMPVsbd2WLdLbFUpv8bsdVFVUigUax3BlD2klZ
MwIdZvCRMglSnhbonEQWL2yvTFv5gsIJD3ICHoVB7QotC8/kPgL39erXtUYnfFoq
y2ZSwnwBAsjI55kvOAFja9ZJdgXZV8kZ416DVYddNoL2+IaL2Eh2AWtZ88QEq8TE
BZEYEYMDNxpo92DPnGXMIcorRExcQB8z6L7hp9dBF9nxWaA0kRDauoEVoGx0dCvI
Ukk973IqLQHNbfivXG0191kKKTL/6ZszTn29GLDzKj6wF0gs7XZDZiwBa1kG2UDo
oC5The9kqWYKygikqv53/ee2zsAEmsPJjOt7F7FGQilQPJd/pfi1rb0TS9MQFg95
kGlb5s6byVs5aiV5pISPF+L9xwSnROvD5ebWnv9UC7lkQRmSVjw1GtEFwqJi0+v1
QSi98aiRzHV5Ua8ikrDUP1Z+yAk2ypTKo1kr8hEYlmMrrbfa1l5ehJ9vSWwCEEr5
sKKbK2xs5JsEGRuBZfx82WrQ52v3fHrTmw8zczYLK/e7FpfewUYLp0KdKPHB128E
0lf1QkXNuLk+WN3NhwOkG6IC7wLfPX6Aqh0vZf6/awwDQ6Q9ZWbDBk5mO5QA1P6s
uOIX4RB8BIoWUutmPAeB5cKx4GDJfrSZx1ns+himhd+Yh4ipig5iuoQtKfWaTbRX
qEglbpcPSHF/QW3WFvb66vVwM3ZgAMKt4UDTuiOz89xgSSHTW8qyZ4ETocLo6nOX
8uSKQYlEHphvUYukMj94QRdyLhrR2zFIxUOvSdQ/61z9XodEO1u9qmijkL0iVi6B
2dbrhhs12ptp2ZPx2S4qoGR+Z0Rv2HN3oOaKSkeZFFRboVWpMoj7/kBcP6s58IG0
tu7fo5aeOK9yQo75mTmtrQu84xndCMm6mkIF+vs0snGnpSubBPX5rUFF9bieDeak
gVZWkxeI75eeMtKUENAwIHBh2ytckl9HenkMyTDSGChterYqjfeIyMos/8WPrQ2U
8+Tp09Sg/hQIgH8KV3ICZuvn+P0E0wXfqoNkWH3TxL8Qby/uj5ANJYFzbe68v+U1
vqoVWQ0cHPiWBbSStpfkfGcuv5OpuTh4jDRiG5F4dDKcVse/5rLjVoRFXm895OPA
dNlQfjilnv+ha1tA4naJmqvs34KpRFRyPTw9Pr7C9DVFPxlJ5ONv35nQAXSfQOUW
GYH7/iIZc+EUmzGHrO1PU1kj727RgkzzopjeYf2yX+cWpMw++6nUoB0s384UfDqH
mRHL3WIo5DS2G+Jt54290HRIUoFvne249zdyS/r+PPfrTwE/szPmALCFFfuuU1cm
LABJH1HJqZMUiwEpPkP6/pp/nM2Ms6+hojqRULoLKG10Xb1lbP0gYS/Y5bifCKHo
/EH+Qz5PQtBwJ8n3wPr2KbrzTHzSH+yubb7xZI5FO+0dm9neafwx8Jq3o7Ap4z/C
bSY0EkAvgDjmksZ4eMpocKWiyLWgJI2RwjqRbHtlq68IlSC7b00hQZ1rRoDjgzqb
+xh5yiwa8r+9DfxgcU/eE/x1g+W/daPQcaXKI9DB96a+O8jhAsaTcqqYMZE5TaBO
duhxjQM1XJfwdgOMUm6f6aEAYsNp1EEOMlRfLXGE03dTNL5kQkcUbCWw1yFyFaHe
eMacSy8rSCudpgSTMIzjNa3zvbhMnpLZvLiP+Jyw7aMfURKzZS5gGcU222pkQkY8
dRxGrgsbzFry0yNAL+5vEGkzpBj5iQp0dHlPVFcYg8xO/BQ22F+UOHxvoizI6OrG
w8ycUfgiOIHoBVRsiKsZHsoBLsJUuI4BOxQQsJEdJQWnY7jKsHYC9L35VOYMJcsm
hNM8k+gdr6vO/1QDirO1DunmSQuw7pT9ygZRfE47x/D+mSGiKBzTJx3Pm7Mbyb3d
JcYimlF9cpR473eQ5LEj6beCgySWE/OYTaNd4qUN7y+V1Z2Y/6r8mKWzkqgJ5mLK
rCnXroDtfM6x9MlriBJ5vTMVttjNyzKZmqhKthXwvo2XooE4t+Nqye4T7SG8fJaW
k6pBFkqU+f+1GIUKr+NnPiCdfcD5+OGmGRiSgBrHJgWrQp6L50Fh78g6lg/cPHek
npMO+7p4UTYY6QxRTMjWAJSBgiK5IO1glGGX6mZ6b/G2+uy+PZcGGhxCVOtb2doy
3kfF6cnVxZSseh2qUe7JTwglhQxCW2KHzCENw/pi+/UerKhQtidY+niGPuTkDGNZ
oGhtS9I87qHUVikIhjWsaA/Yc9DRSkxEw3Y7myaE6m6bALnTa+Hz6Xfc7RU+EktB
8avj0PegePFa4RTzXezsh27UQI0uPh6ffKfYlUeq+m7TKhl6qyk3dNF8+3hCEVde
p3jOOswmTREHw8WwB/McAYq9FZ2ShZdHgXNfuY284oGlIGiWYI2D+i27sGOsa+CC
bVg9N+jCpRIdGvuIZ936SdcqXrdkcKojNTjSFIzNGnlCzvoPMcIhQqxgKjSzVXC6
mvAn7gCnbGWmUz3G5SE75q+xO4JU1Z8cUUGDn5OGHFFDgbpO7Z3vgGzc+VXG7fDH
Ms75uO5JzCbWlJrgTTTOVcyDMyVO1FJDDfPR7JVTGJzkgAe+mnLoMAHUXz0ZYvBZ
+ESQl7t2QzNdrPQg6IQDYlNtv/r2C1pTTiVH/1N/DW4I+iCsOAD6j7Hmc6hHhtaF
KrjpXwoMm6+9Rn4nxevWHhdHrdteUyAWMkSjjRzqxZpZ+jCbruMA3EBAzHxOiIe0
2SWoer+3j/VmKsttM6qbllhyYH4DWxH4lS94x8L4nkipSPFRFMCalVtIyuWDSuZ1
mkfPYt6kjDFPfa5IRI1OYocXNh5JJOgRMz4o4vhWh3ksExJBam+9N0fRF4JNccf5
KQoD1PYQsHXUHWPAOHyu2pbims+HRB3d8/ImZBQeLDLPTr2bPfzOSPJy5BOTBAw6
jEzsV0mV4NFTU3OnswtflyQ7hP8lCh4wUE96x0afIL4n+LhwPJwdWl9bJGuhdNcD
Sg2zV9Dx5ChhTdH1p6NWvDDjp9MKzRceQRD2A8jJY5pgGJh8n+ED7p5+N1NuS0Vq
pKel3f4MclqJ0PAIKz38eMSV/A5k8lCxlpRcOnPOtarYK0ljyb7Y6nEYE+hGmFLl
qj4yoP+27nQ/e1Mif4BnzY6O/Ca61cdj9t3/EM7SU2owlOTqo+eQR3go1xdvhp+D
x0SNKneIZ9ahVm4kw2T0oGIb1gnbn5vn4D7M46KMpNT+QQEjl/a1iO/qQ1TI61bw
bYAaMyTcdT3Ls8vxXjz4nsl3DCZ69JSdfeVAfY1m2oV4kRKRt8a84tmbjT6uvHVT
ZDa31Hp+W4+nwi5C7tD2jqvmcN6Y8Uo70YXE4iJsZIb6yaaS0z001NcLio+3A9Xg
+4yJltM/DANUTH+57FPuiIbUAy6X11dGYcdoC/aBpEk2pEpu19ZB67BpCcrC/oxJ
r7RJmr8iJMk0RIZ1gTtKMoNsM7pvguTMte8cyaA1YxKxlOCAyMuhOfkbq7T2IJbr
F7oT0nvBvvKkv/U0qLTki6GyhEyIiJ3AJ5ckHpUF2NvQVID2MM1DuM/vjLBVReUB
IouA3XoK2rOnh2FYRv76BBRnznXSTLEF2ou0EYo4ruDgInQ0Vt9L+j1AooSr1nNC
+6zRVwPfNm3WDNCJbWxRn0zlHToVd/s78JTJ5b9LGzy4gcP12OWi8z4UkgS04oI/
pfynioVL5ybr1WsxOTwQVg/mGDLLStgjbr05k7FJXzKIweo51d6VvT04O+5JeaQu
keJfZoMRHML2fVlutufaVn9IYZZ+YP/dTlbqCc81daPy9vurlJXpaPLYG9XhjoUb
AlCjHAWIvpnP0GvN/CkLwSlPbRbJsdlDxfwZWuw2sw3OIBSQJZARaKO+0NH6o6ZK
jNSOXbBEW1ILlvFlOoPGkH+GWgwGm2NCaXeo/XIDxqAOJ/ZQtqQ4iAhyFcSCGqW3
kLyN7cjjoubNHSg4p7LjiqjBzvYZilaeyoRIZsWzEH2qhNeUF8Q1qOCZGNbBu4SH
FCzf5XDJEoLIS+6egxcpmeESRKagtnBAzn5jqYHuSX0vaNZuSoQ34cbtcUiykLUo
tB7032zWWLr9VDUgcLOBidnazoQXdqWY5BIbitGdlifpmUKjypNDOM8PHO8NPrX2
h0TidUZ8EORYHwJ1dmBnzF0gl4kQivWRRQ+gUiMY38uVEMSq+6erLpIFB4jcGmJm
U1k0V8ANCj8Dp53a2lVk4KXA9Vw2vF9CGsImuhkRwa6S0jlemWU3PS2AI5j92HEU
+eH/oWx6fduCmId9KXUvFUYBjoN5bUQwtXeMXTdOGsQnJiVVzklBZfdeH5+NzGp7
CF2HQsuqgj27Kv9XkJLbvZPORalKnTTGAFtgQLgSlgbCAj/BctvQPYCEFayX2EpB
HsvlJDumCkNP2wB9G7T1FMWmacL9bcI2Ayd5ai2tFxJxC6BuCRZAJzRcGck8xITq
IFhZatlNqlLAB+PGly4TPVnDR4Z/Wec4lgu7spfTiXdNWByO2eg+/uNnCFXRxaSV
7q5PWLzTz4a9S0JoE2DSfEIMQxLXeStPE2T3nRfFVcqlaxXiYK0It9Y69/W5HJh5
bnizrvYDBYEj0gBKzl9BQ/9j8k/h3++QmlH7wr1/TyGDjKdGA8MgtBNC/4hib8ad
HS9aZHBPKnnVWKr9ZrgDpgZtK27Ugg10Y6+YFztxaVTCNnzSydz8mtCfMVabuiAU
9thROSuqsIJl0T7an8CRFMaeWb8eiJ9gBckQc0/KpA5Xfvji35lfvJfaM/g+FnZs
/6dsvmqB1WAG80HfCZqer4+iMeSE3K0FF/bnxHZCqLecE3Z1TQK6mhkM/NVWO5aG
2gmBAl1+G9n8VhRMJ/BnAoJguGW00AdBrbNS/XXkvcURWQNZ7Pb8PNothAus+R/B
m73ZC3TYUKOZFiqyF4n+447/Hvfy7aaQnF8PJ5ieYRovXdUHeIIL6feHZaxzprT6
PKKJslQs7AGWbCxdj/hNPfb1Hb/PMlHk66lECUswuDte93lrsoWlmY+IAJUXnEFa
BbhWvwuWksEVno5wyjyxhflEaLwokAcBg5CN4kJVOga7mMP7nP87txi8AsCDL8+N
UTETyo7N+IYltXSK0/v2cACA8s9WPSKYnjmck0tvCaSq+v+u9aGoKttjSGgf7hr5
TVPSxrRbAX1K8wh1OQTTTEzRU31KMjlpjQuMWl95OcKlP0SOEhh+fLPFrgDK9ZLR
Fkv5minyYGNQGTfJN+epra9sxdbLDFQLtxUmKXHiejddywP9SnMLa2xjQzf3Qb7G
Ascx4NyOqy69uvXqiExwkTuPTNF/50W7VSJHKX6uN5kdqlIsGYD3ccGkSjAKIkBu
HutX0fLpjH7K3Qj7d+jWWd9ZLxvXEyspHaEjjtNK9lWq9zEDOWs9d/ZbwuGQyvJw
qQ/cg44w5TDw8OjhwcNWomkHJoXykPVsYrYCH71rfSOKrk9sfzJGhc30qXx8Z0mA
FHuXaorqhVxMf6Fi0z6ABVn2LUYiEG5g8+dcLH3hYp2iAVTKWWnO6KEtzuoDN4BQ
AA1xK+ynbDp0jBcnoHvDzAdM3BZNyF95rKp0VfjKVKq02JM1Wl7bycthSCe2JjEP
syeO8gx/+3A1hhuKi1syAgyPUGe6lC54jF48GDWC64pM8uVwFS8Y/T0p+uTveuh0
pMpQmnBI5DRxCwJ61kGAaBQXkUrwJSVu7m7ImlRft39sSS4m+OAPvdQP+nsDd55+
rluYx1Zhe578ktHYMSwUuYi6dBe1CFAQybENJOcH62RY8ARjzY7bcEbCvgLBGt9f
el4gl7GFpe7SkfZPg1BmRVn56rEe26pIv/D+/0zEzHKXEmmJ72/SBaKAoC5dF33+
MqYssu4hkleC9yj8Lm0+aGotVQ7MzMY9ll4AWe3/zXnQqIlaNOY8iPmBisC8POSn
652GhMGHqOkPD+4p+JrGhzAVqY0Vak0rDbkmE1LH38a3vOwywny+wO1HWNeEnFyO
kCZ0cMEHb5te5ddBBkKpXyb7nk5kySq6SBiGxtWega84F0mq3hbkQKelbvCYiwqu
60oMVy//jFtKiNDDqK6QDqHuxOBvxeb8se+JfQ09uRAAQQ3/0gyY6SpLIh+36bbv
sJwnXGDcX6KN2/b0RoS/S0ZzD/t1XiQb4KxVNngdDM5lmz4PSVPp8EYsB7LoRwk8
RqPJ8JRrdrvVv2yVKb+pRNUdXQolz6AW63wgzZgeTgBchs2wGxT8neEl3gGYHH6G
o/uW/cJckWycMdW0ow0W0NuVYkzG/PzwRAJme9Jj7JOGDv5l3tuJmXeA74nP67MW
nowjp/Xo03DQ1wn3osikSXhd3OTSUtMblo8GOm4FJYzDH5N8/7kq6i4jiwFWtJw6
UexmRV09CQYSahwb7lqJhG1aK04x7Su5NIYNBA/Xxx/KSdDQwk1+chveiws2jX+l
rh8gp5/2os6kvc2GWdBUChd+OALDxMpWg97SZ9K9EftUwcOeJ+323P5eV423IUto
HVzKulPEvhJ5OuEsMHMH8kZ0h+GpJ5K2d1Dpg4FRXHUYVMy5di7r0TYt8MiDMH+h
KFjf+JWlIdH0UNEYd7ihbQnc7QnT9YRED/Ls8X4iqar6LATgWvJEB+LYqwPs5eQ7
koYaT3xezIoAUFwxlN3isZNL6oToof1grD9CnCSP7rIBRnmkFKL8H/nQ3tUnUChy
CUpOFeSKTDxoHpBuH01lK5VWJ4ZARCVvKXPDgpqUoOC1z9kpdp4MZq9Yz1Ou6oBC
WYBDQHtEn58XNwbrK8J5XL2FLb0LMWjSpIhgh+yTLipoeg//lSohvz1DYaZIAOLj
aWUjJJyAN2UaxXy6FCf8oqz91a3/cqEAw+XnYYZbVVG39/pxt21eu7WHPJjL3TYP
yYpUGY3z3YuOndhv/mjf1ueOOA8XGYXlRqpNcQyvO3/z6pkqiSxhL/uBVnXmnbHQ
GppGsyKoChyGfEyw/M05hITlvAfVcG3lrKEJEY5qovwHrJYenfpKiGNIURXee+ZC
fOnhkilUEeIKZFEi3S+ZuC99/c6hKG4u3dyhL8eUHPXXVsc90P5FKqVFo8fK9GPi
ZfYNxyRC2nQ0xtagaq469ZnL0Kdn3oUySOiijVDjYVH/InJhDFGi2kvqHbHWldHS
kSELJWISv4iSMddRfFeGv6scuDs9h0egxX6TqcJr5OsFyoTzqbYsaSGssPMvABv4
h9nVjnAl6V+GqK0Qs9EmsRDQPhu0ugjtP5oG6kr68J3iX3LoX0LlnOOMIqWpR19P
A68nVm/doYOLc+NJZkjHzT4QKIaz04Q5vN23p/fvsB4XR8bo9LNRc1f4mvFxjM9n
mxusSWf1bHKxnIz+/2bOLK6YNQp15c47xKOyC5fRiJTdnRzmY6pDmaCfq6G4bfiu
rqGsHhsdf4UhS83EBA4hBqd5MQbaGIsMYuskfVXIkIdzLReMTMlfbbTPPY+dR0rv
XEHkkBoCxtgVHlrUatftNJlrNp1DObO0SYBMrz08RkZESIO6BskWLh9YvMYPx8MW
FOdSMefwutiI35/atjuTcQp+G7rX7zSMs6FqyafBljlYXwvkxEPQqWChLPSOCosD
uuImOraZ2JG4z5xFQunBUPxqHo1DjfAhSIv6UBNzOlcauyKCMeOy8Luib/7al9s6
pZxyFVMUhxRjU73XomoE5UMZtqPsYoI4bHjwn01PN+qlFnAPgiPDhAsEl7NmDuoA
NR3RniziPbL/8eqaERIc+fJGdKVuo6B5iXuYpvglc8oC6B24Zr4eIy9d2hlcleuM
e5lEhr0mNoauk2ouxU9nc1fbglT2MyioIIR7sxDFJ6CygZjllCQ1Lu0EejTGFzIw
z+gJ0m4OzjCyfMGorVrxkqhS13RSagwy+nxscxt2FNVPYZNkOvQ4qjDRZ+fN3/2i
I2FuXPlytICq+ULtkWQ5KVa8w/shUAJgD18tV3uDeX+Q/nkTlaJM8iw00uVnv5gt
/tU8+JsjFiMk4dJGRvnAnqSvHi4CzuflS27mNKcnOaWDOlsCIvwfx+WqErgfIKlQ
gGqOfigIRWhbJdD+LvKi9LmxEugxTCgcm0zUAI3zk2v/BKtxI85g4I3HxdX6o1QR
m527alDbdqzqacvqfD0hRxrVBEMOMMiz0bRZSEQIzpS/iVQ+FzRKnHrO9XLEolU9
zd15V7Bonb5TTVT2WJotdyVAoIBqKCjbBNxmvaLtjSyE67sybiBpEp0teCBr6zKd
zG1po85bbA2hZK/am9tCzjBtR6yM6+UFEDKmD/y94pnk8I5C0WVYce2ZRmsjBA1E
VvB3B5nxzUhy2XCBcmonCaHjV3ZIplXh5kjW7GQzJqPpKoKKF+e7gfanogP63CtJ
o0cIg7rV8BVfloNE1aVrgu0detWIPRIY7SVfkZYq2jO7JPrUiDfbmRs7UsN6xtzV
v9cgjqQ4wh8SRq0/rNt5CqvgvoMrEa3u5bVKm+9s+Tv4sxRZXJKwCku353GDaLeL
EfpUsMYeepH6Xju53dFIdl7SUpe5aQNX/UvdCVjogWU7Gbm6/xCspQ0p6feehRWl
+pMnCMsyzwG78v46kbUiI/Qa8sXY+MKn40gbxbIFlwcQrTLUSKoxG0eHSe5XFJ5h
k+k2JXh6stsaqYB4JLLfQcvtkp8q++8uTm0eGI9UP9mhCSPlLOt43exhSyCOVDjX
VOIj5gIKxggZLpAEEJ/aeC6U9z41eNs25zxAvKtiYF4zF1oxF9QB3ELNDHuSRuiu
LDkwHbKsX/mB+cfy7gWOUekXmAw+KTA5Mq69fX5dK1JylHVriX8cRDgIfiph+8Bz
niVdALOd+tQHNdo8mieTVrcNeakKXMMGFifXhAIf4vPR5TGBr94lPcxTo0nFQSUZ
7HcR3+ynFQPdkGGHjyY1QqPqHNsOw+iO746/YfXR9ZFszXyk/9WI5IWXeIbs1vn8
YKZQIiP87xoMnMXLXaiWwCS1NmnW87nX7psPNgWs62BQda+RREAfUnukQcRrU4Fs
AvXX2Ssr6teUjslyZCwvUmOMSyBLpjAXnZ/3c9ucO2Dvp/0pcFQKmSXnZ6oqI5RG
1TFr+56cssEwQnUIiejkB453txHL+PcZuRDUqIXe1khrH5NTHG+cFmFKSpqzf1h4
K0XH03HmsxYvdq5SUlJbv602Qz7ul8rCd7x9+i/UCaZKqkLOuVFi7D7DX69sVGif
rtcw4Jh0UF2W1lrfUB6jKFE/ydVOKuAY0MNOkEa4EV749cGEIw0JLQX/eAZ9pFeV
bLpxzO9FiJuFGFHOwPRLXbfGlOLahUkqS3A/tKXqLL43a7DC7DaZDQIPLRe2KFJx
RCzPH/9lncGjnhOsDS5WFbg/pRx1VeQej8M+nPXwsK8LtOv6ch3850o+sENRZJO/
70BFk1tkn64iWTB06h1XpzB6eTzjdh/I1TXmmaO8Xq9qGJO6F96T1Nl8NrBzeAaq
6PdtDxgbMVsh28KvAtumLr3Fmd00SFW6JKRIUkFv+qdpXFGiju7slAg56FAHaxqo
cDOC5N/66XpuYBXNOhV7T1KUK/4jvpwlg7apGPwDobhmoKCque810SG8kxkSXX+T
MK24M796tgvs2tRSW1Ea1dQjofQ7zcGLEs1I3h/a/2Gl2MIUS9l4zK9wuuZN0P57
2Ht1fZ49OQtZUR4jVcyepkDnKwquX/Q8oRJlCUj7viWEiVOM2veIJgOb/O8w1Sxv
SS1op99gle+RFhHVgpsuF2wG6BVmJXmA9o4Br13g7ank9APPGeuSyZpzdLgnlfJB
srToVQPws9/jN/R7LHXFJVFRP6ZLn+7O0ZZ/3LkZigVPj7GbISqjTtHuNKqxUHCM
DQk+IjnV1UY9lwDPGyAW320ixKhwHaj4NOx5kcKPdd0kLjRxGX7DKpsmFse29nSn
wNIWhK/0tPYvnAQSqYl2sduwuGoPKXykdXUru+5qxIGLb1hidIehrrAobJhz3lzk
9f52Fedpsxl7siXJRe0lAEXZ5F5TR8VpsXh17A7XiZfOxqf0TZzHWmTrUFHFIpKu
qs6owJEZbTP4caXug9W4Q0cEniv0kD5YJ8YADaBf8M26f9/TXHHR86/h/rDT1w1y
M4359aZXNDrBzh5VQGKGQJhyGLrsw+XeB2YJiBKkOhG4u4vednQF57/bJirRKTQI
/pTBnhwepikmPyQDj1Ek7EYV0qj7MxGbIm/8dz/j1/vyFoyEb7HcwZGNjXcmJmPi
PLB+n7ooGQJuW/gNNJCvYsgzJClV0EjDgRl+DXCoM6xII79JN7jhTcmEQPtF3IP3
GanctdL1prmGKgrLl/4Q5xFqKa8DOabGe8d4DsOI35fjq8k4clKIQkyNn3MuGmOx
o3dCLQCuWlPWt30iHPb4zC3C5f7rDZo1KjLQLfsgCZnzrV7R/U+9xz3ECSu0Y9w2
W0eivkcnPkbnPSCXRmR1bmIbfg/A2NfKkebk1EGlk6HTB++vDLbAumRTq5V2gpao
rjn9MvkHZW2isxk3tRWKTJXTVZLdMkgTZOpq+gYRNGRce94NtnEur/a/tDMG3mOI
/WfAU5XPCXIrC9OsCiDqLVxTHKdgbuXYy5zHOHoCc7ipsaU6jxNcAM79y2xJDZ4Y
M0pilxRBPfVGA4bvWGa0i1qWFjRB9X7zJ9B6x4hX4YgBDdEuWs2rz0yngAnBXwp/
lEHdLKvgxMSg6EZlPWNK0HKRdY8/U63fmPxfQOO9nsPkfQj+LmIv1lFFpYZ4ODEH
+UUNylZ9ghH2/eZ9lc5qgRSCUgkn+TVmPBXqfTTbbTL4VLf2NluWIDZLQqjf52BW
hAxLZdCeW05oiJKLguisUOFk6h5Q7fFef0+BKM2Djql/trbJi8LLui8akZXkNAii
lXZh+p1cVxUbTT5whY2htPs3h0FyMmfqlVwrIWq6hIGIwd3R9RZ3KCwR70mMqGo1
nrdUF2zPD8EMmyQhUbImhvVpRRBkGZCjLGnzTEAG2chVKJYVuMrguH9KIPuUUJAK
H54ulp3gIfmqKzKNrXjciReN0v6CTewA1MPHnmJNyrTiSRYUbU3OUz99jViaL6TE
oJduePFw8wmpG17E6eoegZ5e9YqWlrtWQc3FOENIby8s9goBhYqqOakE/bTDMAy/
KMlZN81eXSlLVdCuxq0GSww/3q8EQqDLudrPceNIHr6WjcFZwaa4BlsU3YQb267u
mQIrhue4Nu84KkW6KqHIZ99ND1g7tWuRHLey+cmOfqgLEjdxTrTgJEtI4t1P+zUY
HX+SIR8o24/EbOhNcOYn+mXLmQzD6m5kqGYgNY3bFVP0oo+bFavix/Er7e1D+U+V
FADb8VeLCIEIIFarqDrZ46/gOXQMfEVY/DO1dfqMGvWnronj8nS3dcyiuTUPKtAW
0jSspJvLhY2IM4SxmW9SJuv7iJY30sDvFuTEmOdmWBZwM1mIX+k+aLfESxo+peT5
i97a3a5XRoKkJrd2eitP5c26o1LsPcUsoKuQAtdkakkS7JKCqkum2MBDEsYoPAIN
mQm48cV0V6IDcduHPwpxck2v7RSlm/DKO9vDaHeUEeIZ2XDxGtcC2GYqJm4+Ctt+
gDdWwQFr4pXODHlTPGJb1zwVbLd/B14AR9XZFkxjy1jfMD+vJUxRt6w95Fnm6D1T
h/j3sW/bos81ddsnqblVV7f/6q31qwjgYCFKEI4dE0hV3srdndB/FV6wKOLFAf3k
3iud6Z0FHIKGWCZGQyBIvypYmaw+c4ElOHtKlLNGFAXg3heluCM9nFpgX814zIpT
H5oHY9wezr3Y4WZS4xffd9ZzgnT1/Ixva45qUefyo3qBNhh9002dtK6Ta6YAlBsL
7EgSoTqrDhEe16eve96heB/PYvo0BP7mq/OVoAnV+MVXwwWFjFfBWEpw6INpmw3x
k7wNUW0qbAMlB4p51nF1AHloHyo8CQqu/UzKWKhyHxaiP4rRcBechrbiiAK47y82
qvtyelO3Yq8C0aUDr5kPrjs1S6uXHUIbmOyq4PB36GclSdqwG/q986RGWISRCGlz
mhpdcrZ0Ks8TBZob6TrMPqzfsdPduAqrFKNDupZi7FpT7NecyOYxQdzwCE5oNX+W
mEv5IQyL1H2rClRLznu4UYzr2xgHZjSq0Jetu9zXlnTHr4iF1OEN2L91p8kcTo3W
s6G+bwVwpyotOYfSqcskeaWytWGqOF0z9kWOC4A5KN2O2JJrUw1q+H/EriSjAOhg
d8WI9LEJAC1P9ssztzwVWHdo1z07NRwWTO913griaZ7RBqRMk3owRJ1qLAiXffqh
rDuzHrJSnfEsxqw0RRy5fIyygghwxygJLrDJSjBx3nXarPSzmLuZxpeMYZkN6veI
UkRfowBOI7Khq5X6P/QQMYWySY4gnYmpTG+fE7Smj7dHzRY+zx9fDJpjz6zxQj7i
Rwp7dbDMHd2GE5H79N2w8G7pbAqtIh5l7m0Vt0CKjWyYvN88jQWOU9JHtOWZ/se9
dn5RlJ1k4rVMPYj8Ewp5AkLfmaR5+hbr7y5nQ+zBlXyi2Wx45ny/+dcgQK4LljpQ
qN1omdDz18T8Q6gDO6kywGjG94bNnpTcnMewudauVHIwqmWHQrSfRZEJbffG4GyH
94mAwEm6DNjVHkYI/bsqqPL81tzD6ZZo0Zgn88xJcV4/iipahp+GHI7qjWM/2mW7
MVYFA0y1LfM9/UFgCJWF6JCgmAAKJZAhkxnQF1d8HojKbuUv46BhlbFa4CqcUs7v
6IAf7m042SFpQjXvVuY8DLFRv+U9et6wsIe7rWGt3BC40z/Y/pveYp9VhzAA7+BN
/qGLNAQ3oVVDRnKxu+82x+9LG/Ndx82spYIAsxE/PK7i5iOy2y1nbmT1g1R6VtCR
fD729//wzR5fNNPanas5ydVbEGgSfnqj/dYg4fc54Hn6Pk9iQYmxavp7OUsF6WfN
KLsJ9GtO+SIwcaSChCwXQQZZj+hdNv+tzL3FgfODnL987rDGo5MBuEbKD7TbsQS1
9KGyLHpgdb0HCu93MPx8lxBltgMCWYuXRcntJkKtbNZbAnBe40v8REKPKPHdbF8g
r+tbTINq2aG+czVsMzr0zVYaFXcOJQbAZ7IaWzqh5klzbZoELE51t7+okFVKIrkN
ldp5OOF+jFuCFS+flsK3IlPvV5BYqflUFFj+WDh7hQxFjMaTAq93CYajb/crwHL3
0fMSfIgdrSkIidaACFhv40+mpsEbzny4syJvzZuy5rVxy64EXr2WFrAs2TTnHDYh
difMqDixUizKs9Iethuo6x8KVXigcaws8z9m3fzpCK6bSZ3cGzwka/o9WrVWsW40
HthZK67UaG6c0CapuEhd9vcAl5/9mtarqZwKd45WYfFJoNyEVo4SHlzp1d88tUuK
z2GxLMLk20hswQG+Cl5mmwET3S+sR03lrKFetIixGvQl76R6EIWuoZlxsap4pQ5l
/oCd2TWL//jn0S5gz+5o5zAYSrQ1Hsk40O/qeKJ0bHo2Zg8d/q9EktTuX/4EhVGM
t6k8ha6ZUo6AxM0Z9gpxE0DNTf2uCsAOI1BsPMae5dbh/p0yFg1Pqbc6sge8Xbqs
m3tjgNZw9aiuZBQJDEySgkoW8mK8yWD4fNtlKt45bxG4xiBcExDgg8RNBNtONy6z
pNFTNfMGNNpkAJkHiqGUv3nFI0/GyF0inTZ1RvJbnaWf1hI3i/VV/FqF40Ksutc7
PyukmNW7b9zHZU/b366HvH62bsawi68BjIkfxO8QByz+wb3lKJxxll2L/com7k0y
htx/b8bV+Itoupvx6d9ckyXI1PcFaCCkTij47IaGDQx+7HGCa2K1lEp39rTNfmab
EbERBOQyoIcRS/FFAS15op2BjlJCLQnzm6aJ0Iff9WOyAz+mYvL+5dye1HeptJu9
m+E5H/KKno51gUXpvwiSEWno1oYwOPDIAeZZTzqKtrjeGEU0mFjP9k8wcVAoPD1I
83jeKm52Zorc0eNRWrGK0DW0976/w5gChVNlJDk4iZ3YwnhCQXdxocxX1SzX0yHI
e0oh58bIFOvW+Nb8UZnFF7p5Y/ILlUPWFGpkdPhZ5TOn24iRjMw9pjhLcNc6cjWB
G3RuhXn6dPqq7lXi75lBBy2Z8ZDm7lHQnSoRp9AJpJurPYHtjT8bCzyQI/i3D9Rm
diF7ftVwm3XlnjsvXRGui3rxTeV+smzcbf5u589rhVenYtIMBfFUzMH6ZMvNtc/D
pd85V0dMZY2cnEXS7h7xsR2yXYQlnAOo/6anOqzT+1p77Jaq7JTAShPlxqkm5c4t
mWfeZRu7QKakj+Q1I4TFHZ6wzK7Imjyj9GLA00raMXBXyQg7ef12fyBTPaI6VGQ5
Vyod0Iu5w54NU2jOQfS/j96SkTOglyNDwczeq4gW/SsirxYQB7LojyjRyeGlCmcY
qRNb9+alxn6D42/0YZVlF4Ews85VmBCGSM2FhZDvknf1eAh4yftvuGpRffuVIsRc
ybXsBqKMmFR554TXHuYWwPC+GRkSGXpT6UWeSerbGS01Ty7CDyVCoYNSoapfXgf6
Z4c1P2VmXfmmhkk/hrzuE8R172ZCzCkhLOUE4cSp0bRUWcTmY07U98rgAYPvckbc
4kaZ2EcyWtmxG4kkCHMGN8548KEVyznVd7tvYe+vyOkXQnOjNolJXC6lr0zWESLw
gxKjQKy4IIgtaQToW/lpTFCCb5B/zVHsvV9J1sjdSvdAzZbqp1TxIEKdS1Yw9Osk
5yXRTHnN2rrtU2Ic4GFCsH8MWkIwOn5SHClbGpHO6pbY/vQcocw/2ftx8VJJiMST
EFWBldWm6XToqokz2sHmKQZmyCdTNZkgclfLw7EVWHeBnjXqV/sjf/qIzRaV6ku/
Bx0VOYLIFZ+lcEUR36PMf7Sz+ne/u0bpZ82pCk8jj7HVwcMnboaLcSnxs8hOJ3eV
LS7UjYF6iPyh3B4WD/ead4usgY+9gS7tXXOaV96TNt3vMHyuGUlKY7RmXS8UaV82
L79E3Y5q9NdS8rN86dHYDEWAis/bTdz4BS9O74YiCILFKrYtE2WzZnNl37zvFa8K
CCEn7RbRMGeaadVvWft40wm3NlubJcr6A+2oBVp/StQGdS4bRTj2rfJdQD2hKOhw
NWE6DTGlg3OSy1q7UGzGmQzgeqAtRjkp93MAztp3HZUn8tG6tnyiiiIt+hb6Czqe
Vx4qvtPtZVFrsndmkkderN5PNbaS35twBoagi/fxkEpcez2DgLnH0/yQCHdWj6FF
Q/hE+SIjZCrmRXsb5y0RaAxt8AQ9Z7sqeK7dofEkSjJdmToVjby8vG86d/p+Pc/K
BDqRNIXRSfG6f5glXJdA+IJYKf3smYgkDacsVM+UtcoAjKD77mSkBrUMPaOAItZS
cA9hpZwunIgXJaa5Sl4gBFqlZt+HVUg8KSwS9xvpJujubi4m1G7c26S1D4Jvsia2
1J9wtOGMI+avOZie6X0Qbfm2PcDQtQP71rCIzPnm0mk5Zm+eQxEsOEtgMSf0P0S9
dqPexA+2TFvrJFHgp33fHQgh7bEvnySQTVPnFFACDxNzP1EQQC5lzRFOPbomwS3u
bYEEBSb4QgRxikM3+36zDVa5SYmCLDAsp3Fi25Di4Y0XkOiZWOqBv2Ot/iXkEnie
LBUTR94EjuHCc/Pr0MnyjD/K53uTYLsTw3gJtCOmzOufStE9Nqv0QSMP6boNZOUJ
5jL51H19pytURBMrVky4/8gPquPgcqrhFle8ssHDkIaj204WdZeGrbMN3FrJCkMH
eglIFP+bbJsSXoZjCT1BjvJy5qxA3+47LZz5Byw+VcaPYgN3tXNyF/MrWeOVsm5e
8PHa1eCrBvNFuXXfu72quvGweAhPVia4nVBXvIeATUQ4DwFTo6qEJteetqwlSseg
MsU2Fa9F/ySe2QLmQfwLNP20I39tINle15297hSa+8uxvdnPFIBnuWWsgAXeeLGE
PxYvfahiu8jHYIZCRCORmNDsEe7/UEmeSbgOa10Ibm7h0hXdurNT1xwocw40qM/u
4w2Yim9X+qenaEEzVIT6SzuL4gawnh9+b4SRYDnmtpkNKdSY2tiKKhmD95EVemgI
RyYFlbYIcTcXGbKjIL29wT+2sBZN+G0WoFbjp5lt0m7559GHbMukAst1udit0evG
ewzXqGvD9WbCYCJHzyyMFt5TLhgjipS2P9HP6J7R4UtnlxPeGDgleKN4vgS/84ok
AXfYEqBuLZMqRh81QjJFJCyaQBakced/9tB1kNfHvXb8rbH6H66hTCVZ7xb3wKVY
5OIIuIXA7K2eMXBSiCuSBGaJLKX12nTHP6Vp32GWkPIYL4fQ3AT8qXux0P9fapB4
X11Bas8j5T8XpOUz3YyF4iqNRIZ8qbP7u8N6E+2c0vx0OEsZSCX3ZzJRY1s2j6Fb
J7tHFi5ESenNH61MbUHMCPm7yDj+wO3xzrZ5qaCtrapkQmOFAMSoCRY4w3vP/eXj
jkLbILMqoEjAuO6OIyr+3DELyA7W17GRk/PAH2eFQxgYv1K871lgL6Z/cfWqzXKO
GCWBbX59Cbs/4EqoNJRABOI/bhmewMe8nRB2U90OjIQlvOzMODcA58eNO57MeC3B
DPoXnLDSpaONjlyMk0IVQSfFGJlln0E33cu18Gj7utq2WdSOYXijUw69l6nctWgK
Yq2w0ujkX/wD9ThQTpCXU8tK/9AkZkEf6hC481WCz9p8zNxM/HYUl044l20mnMDW
63B/WkOi4XXFz4jMFrI2F25h9+Q9cWj86xveRY9l6x6YmbFsCM1fsHfaxAAjTbUg
9hOclfR4bOZ8i2Dfg8QbdECNkXmH9VOsueFYTqeUCXuYio3xJwSed2VMiyZNMacw
AlDyfejR+iOswCKEHlDZ0wyWsIvDwK9Gk410CHvgxMKZSVjWhAIQL4+aKDEZS91s
1h1hj9g/OtQsW3PmsEOC2kJ1P8KW//gZebtle+DMOJO+TtDnBi5iedwScc8L/c9G
UFLHsg0JF5t2K2V4tf1cKE/UxNZuJtUkzSGU5w1zKgS/MZgM+x3c75cq8goK6Iqk
kM+PSJVwm+YJlKk/G3+EIAlwqRNYY1afeNgylgSOI3DsnJWfwVMfEuxY/lKvVz+R
9x3E99qoEwia/SZZMntn9NkXrup+PzFm/oXJv4tzguaL8n49yd0XwBuG/MQt1fSh
xYNNOBy1yKUt0z7KN/pfoSOX7wdgAULMXG3hNBXNYOAdP/mjZGJKVw8bGX+cjagO
m1YYDIEIaDPK2/FGYYe3uUySZyNSaTSArgGJhFfEPsWQkwxU18FDGqxPUBV3K01o
ss0TLQ2TFKuX9d4TOyPT7lUy7sPhGJP4lvUHfnKl1RVOgIRqAl8F4ZxYPU5j5Ebh
OrV7Ceb7oc5Umj1L+/AH+I5ZWN5hlyxDfffxbYgc0uJd9sX4eIIEjU7wccZbKdfC
++Q34ApXg6fvlzvo1bXveDqpi8Ze06iq7f7V3D91mfpoLqaJSi55+eU+840DN51a
pqBYMWPIiT9njXUtMbspQCHacOzQ9TWQ74SY/8bOba6I4hOrelRQ83zaHM3W6f0f
oe6gcVHSjD0NVSq0S7AFNGtkWLaImnQULvtrGgSbAS42UgTIEkKqGNG5aApdw3HC
hyjjAOJOkYdLD7IKu+idorcSMqlB04t+kMDmRbXTaiqGUMHh5hTGiwnbr7CgLCkX
ZteWIYpFszxUlLPTTW0j1r8WYZtgF28LjpvfOigjvGX64yE+0R5wu1CR31XcCEJR
CJxsbgVTK12oJBkl/1xVXF/54P+Pyk2iDBSgTer6Qf5XN03TP8vBWtAn6tsPjOlH
AxRuG57DcidiJFodSveBCTkOHSC4q1WHeZtR4oEFpl6mlyneoJzhPF9QByXAGaY9
6ZhSsyW+ZWz1KFiPxKy/pCgbltcq5QuSBwz8GPZ6DqXj6bO2zvA13kM3It8sQ+HO
fDMOKgVd9XyrMeUvol/Iyx/HigOu2GJRmLoY0dWRqYhspm/AwEbF74ZXwhaBYGGQ
9GwBVSwnFSJMAoYSlfwUJrbg4cPs1aC6UDDcL6cmWWu8HXbsHvuU/fkhqQ9QNtfY
611zQUcTDb78f3qI7yHBVi+IDCgJxaibXf4EzDCp1c/8R0gt1hlH0sIign2XkmPx
l5ifLdJLRDH+A4mKXJAPZ7uSfuFi/gdX5Lj2055W61nSiHnRT3WB0T39NpBGh5C7
4SaQLtwuRSpt1i5M++CQrXn4JQtu8O/wgfsCPu8Yym5VeKRoU2MbJYAi+JIZ4Rr0
KCnaPEIvyq17ZrhM9+q4PlmLJFA4+Dm9ADO6WdLAsdKxNsxEGphc1x0x1iLgOvQL
O/2BXBXLMX50EG7Fw1l2zE34ntY3HllnISkmx3LUxCxeJhAvdaQCJ/UnVjNqjwpd
bqfD5Pa8TUTMNeyKcz1lhPYEhCDxWNAfxe32t+qM/X4PEAL26sQAh5pKiDRh0aP/
MTbB1PNPDHuT0DbWA66fmWl+Lp+99qA2CQlcE4TKFzu/MDaLaXWs8blfDkkgvIh7
q5ssjm8pvU0U/cTUuXquCx06NGfbIJss35asPIjFprn8ZjnAA7JbuPA9ZOD4lZw9
Lo9VsKM4NDhYdodbQMcpKwdpHWrpKNk9oB0Oj6GzR35D7+WvsUGuOyH5fGnrilx7
VSUQnNFtntU3uOhDMOU20xiA3NotWymVnA8yzWaFNtAHr5aoElTyWZdFHo2+SEG2
SXBr1admAfChgXsMMemjA66PU+nMcWvFziFt9xLpFrNBEaZYU0vzuKzj9rRLHXBr
2fR+NjaAWpW33P3YgReYgjsLn1Yh9UbyphteQz9Lod/QmcxGNsMKZJLceMI93ChL
LvOdPCArHNEaaqgE8/d+95RmoGb6OSfsHkIB0jwenEZLDcY4oxjWkgv6Ec2EA5bD
ibLlalXyDKqyr4IqcosfVk+Xc+PsNG1zx7ATGQtCDQyn2XxUpXBirCk4mRuDZzj1
2frowmLsQ5WkF5I+cF/IWuGrgoql+w8gW34EbT/iYBMhYAH6w1SVlmg9iy9Xwdt+
rQXAMCZyVEn4hcXwn5OvQc8UpUYO/7TY59jAnFl4dMLY3yPwoldxqwuG/xBbuOPs
MaEfMu4/czj/FvlTCCvWS372HfDrbYL6137GTI/Jbd+Nod10JXEbNbv6V2p4mMpR
i1JMttXNs+x4nQTeqJIyCFJLwE975ylMYz4/6rCmh0muCMQKJy1dgg/iSuwfo48Y
v3tt1xXmiem9vi0zm/AQcgsxGbNylk0iwY1gfeqYwvxV1Vi+zHxvakdFh57oxKeH
0x3RnNgXC8RtwaRf+yXXgxIU8TbDVW+8aSilCgXnqbCGe61zY0p8Fgu7rICD+NXj
PLHILBq6tcH/EWRzPKZEMBNLtnRsyWtBRoRhVz738fNxpEs6QFkswIxQrzj8WFH3
AEgwNX1RKsVT+R5NaeUHQ7mkhKzw+o6llG6rNAoRivc1wkaiPhxI5rKiPGw3O8/G
UkvJtJrsSEf/wjauUChCLfG27czOQmSVROh6U83blytOC6lJltHCOx4pDnanRZl0
p138l+vXP86b0WwfBYmJn0ivQncIgJRE+WyfHdViMRdnri7q7VUVtBtsXcg2EEbx
CVnf7dtgDNg/AXfdD3rvTTgEZSEj7Dp/BnmW+xhFmEY11gSbCEp1LK/fzGBIAwHS
bmi9fR9sdoghGl3f4Sqs+zsN0tlCQvxS29zMtdz7g3yVPGOnPVNA/B6gL0K2rhh+
llfxor0Yup+Yh3Z9xW6GOXzAwArqHopgVh9yXvvGcW/LXtmqfcHoHB31LzczI5ys
3bXZKhoMjno2vZQ6TuxVdd+XSnK6mPGV6qvmjUnOKCZGkafaMq91asZ8OrzhEt6F
aiMPVNj4XxP0FcpqX2fvrFme0GvN4xwO1YsXDe8SdPbZGiEokp3YRQGoWEZHLk21
S9N7FH9cOUALmQ0oCpvDgeNDqUzNpYYRsbOZdPbxUDQJnqckIURIs28gQRZ7LrnA
DFvJrAkGWz8uKRzJumy1P1OjjmmhjRilygBoO38VKYQwCzt+JvUYEVbAPRmuU1PK
BPyi5K5uhToPn6o95AAVqPCm2TW9M51/QbLzojF0rFuIfq6x8RQED7IU2BMy8ubJ
WfPk5XXpxc2m2BTA7cCNNc9soIsss8XYudM672eRQpMSy6GMPusZfhidkOVTHvvO
wyJmHW7ZXVurvcKgqLuiE0gADSgbrws9v4GqQO8rYeNXucAeAX6Y3HMRL0rcC9k/
cg2OW8DQFxYmDUzm+2eUDc1dN78yA0D0pGZpPzO0HD8j3iKc0pCH7p4YyOiyA+HO
8vvlEEWovhObw0dmhW4Pa9xOOtVr+YyiqeCdboP4h4ZIs1aHMv2kmuH4VJ093FNQ
1gKgU4kkGjfkKm+K6XBiKFz6PqBF/kgNkAlJfERAPGuOOaLWRUrITI+GcjspX9Bq
Sehf/qaaPrJsG9/MmehnXQ8PWy4QHzjhdVShbYCijbMQHC+IlhUMIJydOdPKMyeS
uVzHR2dqSkbe9iy4HxtHOPQZb30lvC79DKFPnrBqN3SrpAB+v8H9JTHFx4f6TKMl
Tk7k2pgBS3+wwDtLZZwdJMr76dYQ01xFSe83zdCVaRCHxR4dZYJB2QqGrHyva1zm
eIhFPqWu8RYOro5QekB0bxlVnyJym5NqyE74ZzQV2/WJQeDW/LGY72xG6YCevjLM
iwyTz4r54YJ/FEQErF8sz7Yc/XsAJWhYwPqIUYJUWzCW0vXxp0Jh5oZzLitrdnke
aj8Wm7iQ1Y5Sj6bkAhn/GWvaX3UES8CX1LaTuUcTQbjVOnNh1WPozXJSs1Njsa1T
WJCjoEnKncDozj+PvTtilxD9lu3m2h7tVTXPEEW+AFkbbDiVDmAYv1JuG/k8XGmE
IufZtWLNrUMACehk6HBlbhI6xzcRytyS472SkelLD3H/JJkDGBEmPAP/pfyQA1Ix
24/AhwlWQ9iyjuK1oMlnwkqKcEkUuHMlD8DBA7VKibLMzuabg5YfV4Q6WJqo10cR
6QMk8dVfORzYMdCO7FGD01YL5RyDy2Vdsi12oVp37pCy8XOLE69eDm77IlddVEjN
aZ+cp59H1cXegzMtZit81+2dOG3uLjXniXJBvu46kA5BP69o9HZ88SktgCtIGjov
I3mS2mbIk2aMnoF5SYq/4Vsc9otF5NlVIy7QN+mar2y428vrekb9/pDuHooHoZX7
kJtmWm5+n/DUxxa1okl8ZfmpgpqpNMkEflz0Tvs69XSEjFs7NscFDY6fkjk+H3ML
/ei1/7CtzMkRh+fW6JxQLKFYenREtOVQ/tlNEw7s5zp4gOyH3vwZgkKK8MX4IlqP
e4LSaz6AT5RKu2G98ZzRQNSaO1GwQkhvDeF/1AOyEe2zgBESbFymy0W4K5gGKA7r
Xn5FUvObsUqwHCB6IAKIuHWGICfYzi8O1+Iajz6w6zdchGPayeTF7e2kaEHSy3rg
Ien1oobj6/X3RJpYBKWWl9DkojTpz9LlkMozNShoPbTByY3k1OSpo8VKESMIAGVD
8guXt2/yUpAkIdzHcuViwg==
`pragma protect end_protected
