// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:17 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
N7T/MPPsVfHU8QO+t0h7NEuYO2oWpLOVT8T8a9xJNtakUlxEku6l/WaLVKdRphfx
r1OUxuQ3w88Q9Sj5t1koCQczammO1RErXr0TR+ZatgEf9DhskwOIHze9k/cdpa1z
3wX2lALbNf446bu1MBgGTrOkeIN19ah9Jn4gZvyDc7M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18752)
lRwO+vvT3IGoirecdKeoDL03Y+He3TrEtYeJ5cbrSCKC7SexRUmRkSX4UcOsT/Wu
BBpCvZU7/oj2n5Psso+kiE3Hln1Pfp7T2mpxhFWvziL4d/Oe41CWJ2iMf77KvERS
ME2GXAumzXun5CT5zIw2A/Xdml94z/K7cJfDn26fp3/FPc5CHqxxQEEqat6Ay6PI
PORW9nuSZAg8IDBdBsBRGvgeEYAJ6GulUqNj1WWDTOSVYL0feskSq9nOlRKPg8y5
MyR8guaSUzjzj3Pgm/0C/bs7p3p7EHI75v2vS45j8ybslQiQaTJRGFsLg3MkhOJS
zRCZXr9BMGl9oXScA/0L3/Uw+DfYTsVcK1j5IGckzdhWShRoiu4roPB4L8/uVL8r
fgP5/gBKxXStzIthkC97+92QYOa5EotTPd1jzgRn4PNpfouX+H/I9CAguW7YrGtP
1MTFYNTQ+6CMS1Kut1izcz7OabDjJyE1X0jyoGU2htmChN5D+qMF/rvrpw273TQJ
qJyvIwrVjm65TObnp9vA/l/7eJUvXTBLR/Og1S7Q5Aso6uXh2XfaIVivGfyfGAi9
lWUTkKc7QEv5uzvqu44GgpsmEkYDVlhXDuPZivPwVRN723q4Mc9zUX944Yc9uD/S
GhYDRwB1qlrX6oD7T4XV4OSzxhuqEQ9alYk0OF9oAm9eYvYLfDoV78ndKBPNVEGx
pmwHgrIA3NAQ/fSryenIDHJk8WwCkjME2wkIWp6m+LqnLB1kzvdUr1J7+kGp3wZt
scqAxxb9jHSbULmIpCWmwO+TGd1XgQCZtqQvsgNZUXJIO+ICDZX9WT49rXsdWOW7
/Pq/AtAJbSpucjIdRtOnerO5sY/p6ZAHkgXUNxJMAg5yltD2c5h2jejhH8982cTi
ob+oCWJ89Gsh/wZqd6zDLf1mq0DQNBnreo1UFqtq9HpPA97BUxVM8PPK5j+ac4pn
CtqmbElRsuMbjaNDbapRpDvq/601MpOd/jsVb2oWUadMUmhdUDwOkbKESD29tBEQ
onn9qpDByzeZ3NUv25CouGTFOguPSOwk203pRv2LjbHqy5AnIezhC6LhnmjFl6N2
O0O32hgQF+/rO5obovXgViNQjguaV8rAMUxn8yV+wU/pJxBUM75k45nxk4M1Azpy
z0mq2tcJdAMz/clRw7q1q7T2ciEuDgnE75UYu9CvqH1OTg35YkFpniIOtAx+1ixb
btPYAWP7LiCHyXoAO/hhfq3tmlIauUId5iLJqpzK0j1nU0b+PELGLRxQxUex9Ipy
6zizpT7QyCnoyOri0BEzw2QuCi5fcUCXSkgEX33ux+Ia3NR82YyKhLYLJnbw0oPf
c6AtP456qJ5/KnX8pFt56xrPOgq9PjRx/6rNhMyEQazp9vZmM/NC5Dom25ERo4wC
gXOphEmrkhuETkPJvwUgkFMLQUuXpdy5l7R0iNrTo1DRbiq4S19UO8+1et1EJtah
LXd6++fj/kEyx+hLBDOJy8pSpOSOcpbTl7MWrW2lS1X7cbN+5OLxPuTKvb6cabYx
ra4+BvZs83EDjWi/2JYy3kwX7jSrzpvzEzaT+pr+UW7Fclj4Jd46o+JI2I82XJFg
wfCTQ4WfYqIIqxOZ2WcYD+ExEAjRE/wMSbJ04xLN32ExjrsFrknUkYcdLBrdetBe
fvK8RkfXayZlLvKurq2QOCj2I3i/YIHv/3i+J8agCihBo34Xtq0+TT2bb7Yh5wYt
BMfH2p0vnpL5gL6pkpFbgAthHretAfsEBGZsyveyqx9AAPntDMrwzdwfkEdUBkui
zZnfzKew0A2FNQCqdahgpz2mdT1Qc1CpIB+6KOD+Nnhf8L3K/Jv82KaIjPQctYLn
AdcVeSE6I5pN3IsXHT1fLXF3W79I0WDfotXNWvrKjyjZfUt5huX9hq+L0mJtpPn1
J6fmEVv7M9MaHWXIZxP4QExLSq+4Zt/NEIYj/PFh8IGN4Kx1T87WYVCZJbSW6Dke
Jej9950rJ0U5CMY/T+TuUmM5xgqHUfR4IrnLco7SJDpNnRpFDgSXiPBYf+gzy2t5
sE+CY8X7dI7ky8TRVt2trgHF40hPi57S6mOeUYmtllXxaYO7E8nkCy11mNdbPoQF
jJAe/JzWasyBPARFcr87xYVy2NAekXfHKaECQ/GZ6uk/97HFUlOl7+u/1TSr8TPs
i6OcJMVR1kXEyS8B7bhwKrZK9D+zl0CcombbpyA5YVqAXDEqYQfkXPftD8IVQQo4
Ficb6KCCqxV6ImX/PoDCuIIN51eiPUbMwm3P5rXfaZ5u496UbhqH2bR0oUL5PoYX
sk0Yfjc35srgMDy0bbbjAWY/V38LZBlxKw1c3jKB+EIwDLBQfNIhE4Y0Ln7Aa6GT
qRILKfTj0yhXukmK7EKR9CPpaQkylnvlRmeD7EWqNXKweST5CEx6mQOwaG5qBUAI
VN8cHVxpUNBbQfRzDZdBfLBnV/B3fqXAjSEE+RnMCnMD++vB0gCNrAa2NwLLHnSs
W/ChswQ5Cxr4F/3rzxf/fWtqTq8WJaEPaT344pfH4Y3w0aBgZmR4/Qn3XNpZY+2h
wRHcmGPgn3sFLEqJ7A6yd15FAvBpXIWUI9hzE9KCk3W2IQP/IRgcQoe6SV4Bycj2
F/gzrIlojjzItlWfjg6xdHPXMY67T8taCws8CYwwpkc76n2iYLDYxnrlfM8cFx7j
0JXeQCfTrgcW/T7xGHm6et/MUAxJ9SINbpDEHY0JBkEiy8UTKfWciogfMmfhZnq3
TGfAiByzvXnPsZxF5DPKaNmCJVPyt5resDfCoBhT/vivyG5jwuJYFisfxRLxJvM/
J83W2W9cuQ2zgkq+XmdtilUF0LQH8TE5P5yWrZ33Ot5VwMEIhNZMlRwwCDTwc0M2
pAepATaq2nUD56BSK+t9eOzkqC1ZJxf/obSz0/ZhblVbVU2iio1Ci0qSR2jPuaLp
tc6DqAIK1UYwBuuzu7ffGgPGn28KdP2TxYndHH4eFAgYuZGRbTAAzzMWt+EE1Kc7
TGn4m/4yHpL1ByNXzmVnk+tegwcndeYCxKDfJAv7Imnq7pooNm0KTBNmf40lx5PD
U4kVw/ZMrR7EW8oIhidd4q1sXZ4IDHVROEbNHopXB9dQwaxZicSVH9AyB7gM4hIG
ZKvWkxySk0TLYpaK7GqWorXL9w/SdjPs03vgQfrgq9o7Fj2cyXy5jVRr/SBdzIza
LiaGDLsk7v3GPe3PueinYBXVK9V5O0hGecz/gPalSopYuQISk8B8OnIKfNtNonxF
utxz5YqsNoTnRpjCYl4xnXI3Mlv5ihwC1AlJX4hrF8iLoeSNYHn+IWMoZSPnJMXG
G+3vgA7E7Tk+W7zeOHUW1l11n5xU6qGOUk7vDAB3d6HLk1HteMoyDpd2ae57xc1V
vI1BZP8941spSSOFm6jOD0qduNnd340gAYot33VT9RYQrCcxUjl0mZHjhgWZRHg0
oB5/T1E721uy53OJLNueBTjsvE1dQUrnzdzSfCX/9rHaOVzwrfUG2q3gM5rNWIDY
KTkjlCW4O461A1wHX/+nzLbtJ1nD8cIpfel8gIoLmC0BierbJuuxq+kSM2GksiNz
wRwRK3miSK7XwdRXrf2P6JDZpS4tNNbV7qo2RlSf0kwq6Z6cUVnRS4zsrdK3HXWs
FeOqKuU9Ut9UHjjDi2+MWYe04zv7jrXiOXzBHiFtAYW25dvfpcpwZ553xzCDSDzE
rGrd8JIdxcjbuGNcnk1N9JgsoqCWCB2va7VErRazpsyqDNhAJB0tCPL2EWG7yKVr
HQaDF7uhYbPeFWdVoy6FKQg1iIrpCxzJRAtVTCk80BCiZeodxzvaJ1XBmkNk9qqC
8xScKDQ6IERL9YO+S655Fl5pzFJ9x1B4+629XrPAoc2oTRHduOsvNqEcuPNNn8c0
LaMadxNa9KFB24mg7E8epSRJRVDeLAF3haQDX7OatCjsq0TsZE72XvIFTi+hzusg
ORULxwi1/hxnMPmLzIbh4tHusOl4mwzN8fw3wAL6QEBvrcUUks/73ofBAxs9L6gu
Tr/YTgRNQgo+ABFzX9aWYx1ZW5JFoGfbfnMU0dYDYy+DwANGk6GlNZk0+uEzSx22
uBITIsffw2Xy/UfPAQk/V0/Oqkccp0dGI7jyJfeq3gBeOpWtmeVTWxJmVOKMKN1L
Rn4Nxg6hPgDR5VB9un6ic4ziLRQYatY39OBZxhVUouykmxgBJij4jaQXp0o5EclN
VGG7oPzr6lRVe1bAdVRcKcEg3De265lRtDM/ALdmLpPFnXlVFq3oo3npeHjjE1qU
eT5UAN5BC7ZJvBjfDENP2J34mI+GPkgfb1BlDauDQmcvOturSfm29dIjbY3qL6WA
oSvQJfPBv50Lj+4gr7j8Rtm9hsVAlIhgFLOSbXmtaVw3KzzFssNhUlBVYqEZhM4h
IRaqa0nR/Q7Q+h9KtUyYvCv5eaXFO6QotJgaZW2Ip+GiczvYWK+2sBrJvVmjTnJl
WyKCx9946NlZAZdiC/Or0bY/ildwuRBu6skGHEqYo/m1pr0d3RgxYn5xaqHsBCyl
QOjikURocCIhq/DPvWdO810wlO1x8R1fT2fr9ApEM/3wknL0U0UhF89ClxuIV/zr
eeCr9MVXdfdX9NsECVR47Okdqwe3UbBl5e+fJdAIb7ac3entVTcBjikDMY/8NdFe
iOa1WwJucR/wJCfrFa9gpoE79tY8sLfSYFUNlz3qUx1Fh0+OZZgvPENEoKQoWRZg
Wi+X2nRvDUE1zIiQAp+I5sOn6f5gpfNeOZTalNUTnxPBSaXgKzkv9MaLbIyJXZp9
ASwr36t28B4+epSL0FXBuai4vPCCACaxOI/VXyzFizA/XH6d61S6eSxrqvxLoy7J
0/Bg++OO4X1+BklaGO/+tmmSlNAudOeF2n8AjdEKSjRtsWP4yK/sdoVls9j2SJEf
YJTAnDwPyuMCmCnI7AlA4GU7O/5JGyzTHv4nw9yu8i9g89laSlNRUlUTZKfl3iNX
GZMWyurHMUVbdN7XTIA09heaXQsykENfpXao6FWi2UgZLrSyjAZVZkBDd3davaBZ
9s3XfVSvOenPc/127jjQ6a0nhbQ9cUH83TwsaHJPuPBDLlAGVkYeGWhxdcgOAsxi
eIQJkWhlvZi9dkPyWL3csSVfZ0VP0Z17a4MRlSN+xRF4L5+aRRlpjRVr+B5peyxU
HGbGOMxsJyWRBcvF3VfdijgGZh1n/AGoOG+IEiGhaWTVxOZj3TAPP2G8/83amVl/
1NwhBfREBqEiKeEXXOk7dynvjd4qYczBhG3xuIfvpRDfnFPWz9t1+AkSkcfMejBW
fevEQGkBnq8HqOXNnfK+jmguhT4BO9iRboRrrbUV5ZMmqHLFAYrR4HdT7n0bfVkr
wbpnKW9Xv6aCMJnwUs/2dbZM453YBpZv9gJ6EYguYn/nmMNKM0JHdPldqJlrWSDE
pmP/A1MN4D6O7wE5CrX+bFIQTd6EMlKtrQkM4F2qS3k77DmvuUK0WXDw1yN+1Lyi
bS7l866cfC07r8+XpxZVwYR2afPX27j6myGViZMnnUD/AK6IlQ40XiP6qiJadMAd
jiZiv0uRL36cIsa0Fw9GbXHYjdPIAfvYgmG2Rr/nevf/wTk9bKGIb/qEGoE0pIKu
EIf0/c2Jy5sGzHzP1LIoO7Y6a39nPk91ypuIvdsACq3lxFzUufFGGoe607LWwZHv
Ico2bn2kNvPanzmsb4NGwHzL8CdqaC0Z356sB/s68JqYNmDxkKQGEsYcmwdXi/CH
ldHbYSdsG8zgJVWEL6wHktX744Ouf5QZmEcaQjEiCLOVYOBGL1yS57Ip7BYxzHvj
UUlnvHVvXMmWMGX4NYyOGWrcvwnGQcEcoOOB19Y0gRWueBUnO6znnkPJaDB4Wopb
f204ekrVs1B2CC71OZjeCHHVOO4GjYqBKwj8lTbfUw3119z8Zd005Aiw8K96YIEk
5izQ/ZKb3AKLDnk5BxfYf2g2T8tO4QC8RJOWEHXebg5qdfHTT88A8WZSmWKOKVoF
0VvtLcKwBKVFgUgOW4PMEjvivjkDLNFNS/xgxf08VMeeOG2XVsHxKieP00ZXac46
WnjO9eKtqz2EHoYuIigXDeH7+9lJvhAGx8mDj51TMvgldGE1fDabwQXX2qkzmwFe
mD+j0eCPaZQojoxitlXvZPDxEJ+2QmZbxWvzIggo0QElRH4BoxGqwzHPBZ7PGiHt
ZDZaWl9/9TKlInby6YECsGN4HRz/o1lfXxrXtsOIZ7YmPiFbm0QaanGLgkJdjKFN
reqtKqexy4DBuk4escmSNLS6Hdi5WzQBYQAkDQZpDNsJ5/mjza1p7t1h5Crwti6F
UZDNx98TPHh8eNzk7bv72dH0Grp1FMejMWchjX1fEZnle59+1VZrS0vfSVqtpjnJ
jM7XplKYYZI6wB4S5ac5YTq+BXvD0qOI5jeC5nZdX0rO2Y6pU4boKCYEtEsdBRFk
vUBkP6B2y1QHJZvtoeOMszQONqFEEyjtzS6JIHSQ5QD4oy9EMecuV/+8JwjVU6EK
6348JfnTYGopXE3/u+TJVmZ+CVf07MTmzjy3V1m/4O66fB7Ijgb0xFS5UxaG3u6m
BXgoRpO/rXEAOOsLqhKxCz4A7sYkZ/03XD6j1sG5zo4t8BOxUCSLQoZRU8o7HOh0
sJJspZPMRcCUps63TAbc8n+aE/RwCW4kBnqAkI2ydqjOZj9XrjeGD2ubq2w/gB8A
goYmx4BNUE2WEbBuw7wlu3Q2xXv6ocbEzJvil8IBlZXW+nV8Oyd/zvQ+QAB0xOMV
DCjGQfMyCc1XS7VQn1ZRA9XsGmsc6nFYxuDojnt43fXxSkcWqQ4IUv7JTmR0oQkO
iK9gGUt0BMX/V9PLLeJJasr8pDHA+otD84ipe0Ue/mmTLnKvDhvR3VX07IfBI9jI
vcLImKbfy2JXxatfLosidJj0jUS1xoReKc1v8ZFw5SjJ16bfJZQATiNf+UeD+pUC
p0kvQgCdtrOmMs32NXE5PMchuqf9AjrKJAj0S5Ug2W+JfX4r3KrjQc0GSLAwTMD7
2YhB77ZsS8OEPkH6lgyPGpRVxXEdpbeO+xnibYr+1f1AcQLsc5ZRjCo7qhrKXvJL
rf/5M+mCi5kJ9my2U4WCg92NYQ6KgcM9Dsp0khT6qFx71QKGKyeMDPiLTfGMbMG/
gEhlAW6LnIfImOS/XuoxSFGyFbTh4TN4zh9DYJXEM4JgvAupoP0BVT7BtAD+mbKO
ks4HsbJdVe4zZIDCtdmlVlgyUcF6BdIfFAPzmxnNn8h0BnvTAAs09pMpCS8nCKjJ
mILriRHMH269+BxG3HYaZXUZhjQ5Um3QovZnlbUUjQxpDqUf4EboAcfWjP76cPBF
G2A54YvxaG9DqXva25XbYiOxEDYXdLmUsrMaElZ0MtH2qUvVTOsrxoQcCDelGQ/z
WbwGwWEZziHHNNbys1QPyuiINN35tUFCv7Q9Rcwf8c7POyPrvi/PZP3nJm9G4j7+
+hbBjr6nQ7LQo46NiwwbVUfRp34pjbVLTDJ+h0wYBfg6qmxNt1X1qe5LJFPnbole
X1YbAFDc0I1HybWYwO1H7HPvId2ukcG/kTmPHl4DbsdiluwBPAnWUcvOV0Ihn6cM
4qwuqOY6iJRIXF0UjzQDdXPScKM9GK6+na0IsrPRaJ9X6A5q+3901tFJ2tMJnqh5
bkLKg5Nuc6CDWDiZJcajnksGAvdzogagrLYzhM0qgNwqelQiQutwRMVtcgU4w4qQ
ImAozhJ/Aj+yU1vKnJ0j1pYOIZe5Rfat2mpc36DbrlTZOdZYDYxnyXAFOGBSaMXc
aO9vbJO+khOcJLMXSjzZlP9JhId+KhaHdB51622rDevw1drahGK5YOSa4NbcFMmG
K9PVd88U0YdWE5ncqqyRt/w18MnVin5DWtubm4WJXfhjA61Y8gjQaksv7WRb+DiP
motfEvnqmpVRckIfTMyqjRCnyX6RGIOXJ5bdwm14MotGzJWKUZhuGvsTGqmaxanh
2BPboBhUqbrtJKtNbA/YaflPZ/GA6BDunSMuJxSgZFjwyyXRvR6mINqsMLQpznMp
FYs74P4B4FSubkK4pwvXdxseS6r/kkehUZIJqdEKPyaBJKX78VIwycTjUo1Y1BwQ
ysfUV6Ejs0jhIQ1WcTvzskrmSB2QBnwmKwnwcgkHYidtW0LPlXK2oeG6V6CD/EKU
n1MJ0PYQtnutv/+Lvg/CI3i9Go4QgZF/cHVMOKSNJhnBhLESktBPDCgmA2l/R43s
GrWt1U2QSRz7VmPZo0A0gw0xmK5isHkVkXpHybuTB929Sjxhjir2UB1Gpmbt+rZE
d9L1j5KXuzNlLnP0M3Ie8PIC4tEEScJYnr/t6Wjtrq9nPKvL147fT9TeZwXt5mvM
/PIiRzTNrJM4aR82Cu+uHze4sRzxkKbS781drsI7grBJeVqYa1RZviUXdRwGpARY
lOF2SxuBSBNLzYKoY/RvHI5SdpchNDxEiDT6k2LFJ+EtCFr/doYeILBPXPIHkZn5
zNMYD6xbd/S8lcBC0Xe8B9nYP6dFOpSBPzz1uQSN3kNh9/A0yetAOtS5Ow6/Ssxr
bG7YhvTCYGkyi1MCnWNh2/0K+n5hmudDtvcunxuJGsLuC3Lnb2L/GWWL/0dQcII2
ZTndgSCB5POsv0FB3ZtitQ/VSQEJyowf6gX2ON/2IRYtFzgXBw2Wpn3E13R8UyUo
asx21x0LSq77cmdVWyuycyETMh0uZR9PYhEi2cngIO/VJ236eG1dwqeLGw9Bv9De
uZxrgFz6USndIktI7wTXUCnrIViyYiQAKgRqqYvWPogG9oY/hQSx0+Xu9anBmkQG
JrmfYW8cSIc3QTE1XQoQqIbhWrL8esxtdg/t2QspbBqs6oNaWwbF/TGcmjM6HyjV
7R3y2NsUIJQi0YoNVIhYzPDNxV1cLJBf83S61skI5Yj/GuxGs2QGWj9sSgZq+Pzu
WPo9XM5ZP+0XZd8Jf+VbXCZuD/+yhGufD25aZIwmZoD7ViDlQrxFzsqPhk1hwrlY
OzLpBJ83SuNAMLE5w9adxXUJfPDyVjhv7dR1JOBwp1nfd3VLepxCsosFrQ4DUkbk
nnJ6E98JE112HQi0r5vSEM3CZjmf0ansB9srbY3LVRu8CLt+70rsCUj/KKFJaj+x
kjWrYCfcCu2IncLRSy/d6Ni8VpVE5CMXKz3GGVemkEA69ko4AmIcni8R0VA1pYKc
GElVSxf0ohNMcdlzMDPwwpwl95EDj7OEeg65TOVUwP9IN+EOz2EwHel4dWFWZzWV
nhP19v+US2DIFGhMAFcBIJhgnG9dwJxmZBNFm4M1vhddFPE5nvot3Jj2IvS5XSSi
Yj/3h2svqhNlQNBkTH1hGusDDmuHbfmTy5tlf37sugFStoWViWK91q5BtHp02Wrx
aPz9/SpBHkR7786eF8maXwPsYb0vd0aTfBh6+gBegzCdzppjJSBHZoNVvzoADNPf
yO1z1NkBrIqnjaR3ZJVl8RIpvNUB6/aDp9KVan2prWEpHTroh/FOU3UPhW5zhj2I
IDDYiKmWGCai2xkPOxUnOk+GNpS7F9mw1Afyzx20y4rRcMLoUwIeo52N9QTmnn9U
cOsR1ce/mpaXeBt9sz2Y9b9M1gJWwKpxORQ60e9h2RXaPrdWkppnYAJpET/kCWjp
HMglvgjYbFC0fPKjcw2H/Fislvg1I0qMO4X1QHbNgaboWs2CgtR7WE8Z9eYbcwOZ
fjzTGFOiQ4p0FhdU5Yvx/tI7NUuxqWeBInICvJlduvmU0W8R1uA9rxjc2Tvjqo46
NnqXKpuHqLFn0yC25/xKqE8qKW34d5mY054NABCCNc6V3o5Uq0Jjuq5x/2EaYBlO
aP09Qtg1Vd7t9RByqPde4fNTNXHSvDeifelUoo+1dI1LCameX5vnGb5w515pvVt0
07NNA5ce+jlGMnDESy5cfDq70i2vewW7cT0Kux8JzHCv/o2EWWEeoHD5OoyM15tp
JsRa5lPwNdLoA20GSfiX5csa69EJvKXvZMN1ZCP6tpGS409yvExNvkhmk9PZ2TwX
nAS/jE2iodSZEvfsqqxR4ujf4E8N97UR97fRmg+a198Rj+WQIvtcuTSK32e8iOJG
aFoKK+eQM6DVrARybhiDx2Phi+wICmpWIyRcjXXADeiKvrqpvyy8/bjmgPlWUzUK
mKAy+BB7X87TTcRCAEPjLz1nceB2JiOw+sHJwePn7kepQeCs5pse12LogDicW5m6
+hGDEuQrINIMJh6YjYHcBlqc3C6ovNTMHC0vPlN1r2sNTnAUAZTSR6tm6GkdgeUp
xVxgXT1nIVygJeJb3duF2XqaR6SQkYrrNVC0q7WsX1GD00AN+DGSaSqgtIwSltyt
lErORMK1tOFfksDR1mgaHBmbeaGjlBRcdOe/zFi906+HGurZQTKlEGUaiL48dmwr
Fd+N7Iv970AhSoQ3rav4dn7qUhPaEpH1H1NwPlocKYSIlqT9MwypzmT5iJBmnc/q
rfXaNxHiwuILapbsSlSICC4GfTHgOdKcm96pnzUpVMfkRr2OLXN8sR1ZhwTwvTPm
JvOTIAU/7gpmErAxRjHwGC5y99UxUPsVS2EaIWvXKM0ImxbkwGKhMFLus41u5QwY
70k+PObDVI0nW1Ea+nwwKdHUtqcACax1S8VjRecMLipkZXcfXHalP2NPDyDLDaI1
krczAosdrTucNnVcWVH8TN3WwOcDysoQR4PfFK9ohHkDORmEoz6b+N9ZxfdweE1m
i4fRaAtnGpHTfTWir7g8/XRbuTeS/YdHTVPP+iKMAZor+qWUEUuJmHzXLYvNn1uL
18sF2lE4GUxsEf2EHC8RztHiBkhtFg4Ke+S16o4w2kumoL22eLyDqTf+rEmMSk6Q
PnYjoU1rVLwPrX9Sx+9hdM8CFoZndZfIu52qH0lKTZi7JWO87WG8U6F7IbPbY9bg
5kfmwz/pNRd30gfJsmdV2WrhQun27aMvG92sUQHFQ+6/NKv0MVZsLjAEvd+jryYs
Tk27ktViBYcC9qvP0HcoiDtcWW+xLWsNHsKkBdwiQuFJF9RNNSfq6Xr72Z05Y1Wq
zdtB0TAPWYIL8nJfQnhy1u6/fZv1d8wb2ILwXCsGhszZ5p7YT0m/RbGi6NZWgW+A
4aW9I2AfJ9lO6d0yRrQpitg6oDsaeagjAIG3VS7EKcB/6LHEyDXhFz5xJ/3drarO
dukmnW0QSppxPjR+9a2Fo8aTqJ5yAnnzldAEOALL+JnSkG/hUSPcRviGxChinnhp
uPIeF7u+bonz9UIbZbpurigbY5U3iPVFz3lGVcJI0dPnXOJya/BVXmybFW7oiWgu
LajMLwI3P1Cd8l6me+aQtKMnUE36BzihUhjp+3/sLrVGRzJC3Z14Nc8Qgnrh4yvM
/O5TL8EEGEs8gU0OvwRU5Cbk1tyIfiWD3bRW3+iesjDmMUgFUwtOtPyCnNRpbmEM
Z/nImDCRXGEJA1Y8z/HbfZjbUFrbGav0ZxHybCFm0sJ9fdZz2w+NhSt29ysmLv1g
tpvySv+XMDIY7mXRfET/2o24cxGSxTw81lmPn37aAHxdwqHsfhqt/aMUIbTbqprv
+vtCWWlslRJdjKw7V24CNdzMdUsSennv/Ji84whCzOmbCcEEis8H3EHIWKP4PjeT
undGyUWPRaJgo2jPeSNfAC3l9Q5IFZ5aSE53uzrsp6NzSFnyHL6TL23k0xDro4XO
OfaxG2372ZpQ9O9m1ICq6sZa/cfxMGOwminyz9xx8KgNUt2jKCho4MqCO7Xlrgmd
hN7k9WgJDBJY4aPGmNj7hxOg78HWjQqzx5alaq9iC36CnhR380wOPIehd7Pzj4p7
A//p53KGytgUKlgIEgVsStbYOmlCeCd+hLRun8/R+4hqgSkrwxy6mFmvVwv34LCt
nJkCl9mp9wIyrwrFYIQwLozo4vnVIenAlA+IRwv6opya4ufqdzveV4IHutjvu4tM
o5vBYVYv2ZNF4EsSS+Yx6kiUz5OUY4XRLE320r1Olrd/+GBTAXmoiudY4VZI+PFT
mkTYlJhhCv7SHr5F/3ZvWHU3NnpikAUhCL7fACzppKD+wtRa3/QG3HlGFUqTW8au
pzkwavKNik65oe/n3uK9tSg1RfJsDn4KeW1dlJ0LF+Tlyaveu5bj99Llac23wZza
sKd1NB0+fofpI9XBtvmPteA8O91Qjv5CG6vXjCCK+s8VQk30tWJFreH0zwGIxdVq
BDkRD2yWfQt192Y9JRK4OPVeBSwWLxBFbVd8PA8XSB5JUeIcnH1f+5oa4W24G601
vPWisg7ptngOsPl289sB3VYpfND7dFWzHZTMZ+slPlrf0lox5OANpukMplez9viM
0FslQ0grK4W/K/7fxfjQ+5B4H+sB7hHbH1IEpX6Qv+dyFAW09Z+AKAj6YjtzF1ec
iKqRS/nfJYFVTycfAg/Ee8u0anJOyi7IZaRjk2c4+xNqvWtvwvE+D2xno4883OKQ
RM5ZK7ENOae2veI4EK8HSpoJgra4pmi3+C2oTq7uK71ZJEJ60nmbRCf1EwXKbYov
pHASxjRMYuzvHDqK5X+NL7FUELrFWeOAMWL6X/kD13t8i5iqykmf2aYQwKmRxak2
qTdJ4H8wUcvrXHMcAPfZQMGzvfHkH/db7fEJEz+IjhUFACTWPp2D1ivtFYSsTvhn
Oupn7FO0qum/h3pQeLaq2PGV/KBD5w0Q2A9DyIG/TMVZEG1M8QLLE6zF4vjdzprU
lzUYA6wn3ZNrw0BMt+ZYwX+8BhvfmJ+/+GlArvxsVDnokCTMbxTbX+vrqRWgRlr2
MFF6eMG/DILp6ltmgAKh5F2SyDGN+IOKbBbwcx7VcWFAabob3boESX1NE0iwY0YE
fLML+19/QyznrL292bBcVReyhki0XH+v780Okmvnw/uMaC0f1K12vnEoR93eI+y7
QjY0vC6S3pB979x93M/C0daV5bjgr9aebUeQ37EeQAoY0o4/mhH2Vi9B37sRfBcv
73UgsEP+kFLYixsty4ARBM2SznWQ1HVUxXD6pQFe7hvDDXhqtv4YOu36iCvfkhfw
FtSLZ0l3dWRVdhbqmi3zD8bd/X7lqqp8yN11dj9gfjgDB7WmBfsj6djqF48IBkOP
MttpWWGoE15OOL46w1GQfH63z9RejXh9/qw+tYWCFY0Khi1nseaw8Q88aw4bVIrx
YPMwWmOWvoGRK1qTthY6TxKd7qqvydn6150xT0vfAho+uu7mg33jisFwSF6bDl9w
59aBUT2BxmWOPv6BGY/F1sPXggCOcrgI7P4zP/uwwcLHOIAV6PDn7l3BmHho+pkv
opRSwXKNpoUaBSKC+FA1yqPtO08eUJkmYO/XhSqJOb75wkmZgseeQuzboESQrXZ3
fUTKHJDhTC6qcQC57rFDgYbx1pMgTQf76VQ6VmvsjLUufBUzfEVTjPZSdT4CgTX8
/zRiDQNbGZ27k29FbaYP6LdOIQUe2C3idEyou889Ah2ixbCVQ3Gy2deQN/fKD7vE
8C6G0EEDO3Q46J+zKth6NNvx+jvK2UvlAH3OY6ZOzVN+Vas5NhTXEsX2m3VK0pfK
/wQegs0k83u93vhv5MFEdT6p8kXW1E+BJLCPHwA2zFXb5n61lxo5UkiT3RbfHhiM
2eYSVsZ3dZUH2hksodkAsfvPoYUA2PwmY64vl7Ys/W6LmcBrsgT5pchXD8y4a/z5
YDLSIE2i4vuFRRySeG+xW+srnjbRYtjszZkQMfPW8t5Te4cBmNBlb+YVzPTedE7v
gE5L/8v4Z6snHs6G214Rfs9PylYxBSSVjsQ2Mu+W9ua1/5J3kTJhyRVIKloGl+EJ
Q4Zhe5PgTeLrluxoFiof8+tLIx/HwlfBPOwc4WHbB3Ih3CdTJrJa2wecobKGXclX
s++AjtgjLINQcVQYY98ZhJ8umgnLwOUkdwfjMFiqnVpjjlL1UJaV3trqWapstM71
5PHODwd+jScQMIyvrctGXcwM8zPLjXp+AUkB+UuLROspXrAJldLyrwRjVwiT23zx
8srsxlJV4jxtoDLvASzWt3t6/NiQ4W8K+MLi0gMciCXZkUHqbOJsf8n9MOqVFwEB
Dqgj83e96SHI4x0spdEVwQBtc+X+rwLwdKghlOKB9SlWo4ccBng/3LFkC69pleoc
wVbxliyfnZOyCU7pdgul6thZihURQCjd1q4gD7zmYEMg0HXuawLPt1o22adLUjTX
oKH+bUiKW8YPEolbWPhF94QKNds//N2SNRzeNVlmsGO8J9EqP/SoWv156dkWLA42
sVhycNCfSJUi05cjgQc+4EN4bUU5OyYA054w0UP4dP9Aa6vbTUYv13XcyvKLp0Ps
8J2DEv0Mv4AdkTRJ9Y4vIXAgcYPd4x3RSgOvVYDuD1Y8+8d3Ww568T513A+kenMN
bDeYeDgkqUuxfPeUSdC6YqHxewcGphretA7RF+ftkbLjZPmBNf2uwAljc9jMp/Y6
kOqJ2ZJAr+Ig2IqhJPVMXFMEWB/FN8O+1rVaHGj7rXaFEvqIIiLno5PnyRofLVSs
mlHVrmwUkWSmuHzNH2y4sHGvbiT9kBujeER4LMiv80A27JA4PTVi/oJOxfZHe59W
anorRCkzCbv8Z0XC2+o5qBq2zo7raixR0GrZ5sA9Sg6vnGch4wKE+bB0/jzGkqKT
dm/fFAEGi9IPdYLMiDkaG9GrVxp3c6i2Q5gFLTuE0a0suH9zvJYlmIDhEey/xae2
cMKXMwhS1kcYtnp/98E5YLUFzE1w1v/r6oeQyjNHsEbaHBvbpxwlyVqTM2q5ofdT
mmqAIm4/YqbBYZauKAnumVPbbUQisjc0kFZtr9OqtAV7JBsiDZ4LWtsnHo2LkjAW
dJtb29Yz/TuPhjr0ArE2wa+WYp+qHqJOM7H2Orb8vY3NcA9eCIhQ7vVqphmBtIW6
yytilJlKjf+jaNQVb3vpUCBTUOCtPw2D9Og//IxsqN4e9EwJ5VhZPziXWPZv3HB0
0aL9H09NssqRXhujEbl387CCzEAOxgNmSQQZ5l42ifDiE4pEa5TUfoS3ZqwfbOS/
McD1aUu6nxkElhchtO5P5nSIT6fPKtArBnahFD4iZI4HvCirfeZHmYYojJ91M3fU
5JfK8i9X/QJxv/+2e7Qof06ytQdS/NPxFe/fGqjD3Go9oaqf8Ua6bvg+yiTorhx7
Z0Z5cK3nfUz32b++Q1IthWsi08rftn0frqtcHADZ+etexNLu7qzVJ66SsJnQC9ZE
Ydgr4duK/bTTE1XzCoW8AdwPJ7cNmzUvQVtDd5F+QhORkIrHQ94bgg3QQpH7rNgr
54M+CuB2baLzRlOQK0LgZHQS8M4rccDMfZl9WBJtgdGOAcVSw1ZPJD3OoPHEcBAN
SdRvaUu/k1RB48kZDm1GzP+DEIwZNm1+AptunzoPYZUuw7ZYj6O7KYhQWvuQ8qJj
bIpbCspNq9aYh0obAi9jLCUgQJSc5bkjIp0HVzmcTHOYy3TS+cd+oubqMu7sqWiB
tez1Jyiq2btyyGhbPg07JvcktTGHoXRAMr+9FdEx2eD/RiSyL+/T/nR6MciVjtGr
ZRuVialU6iLqgJQQJfyhliy01mP/cfr6dh0Tlw4Bqpn5vEx9uNy4CK9OCRm/W5/Y
t0bVsAyBhhFP37Z6fk3Hxkz3amQILnwhmc4ImgOIbxGJ6gZUEdr8AvNzgwTNz2Hg
9s1RN7UvoWhU/Ndvf9Dr/ZN7GceIjKwuWoOKZMzshkmlJ3jv67IQyE5ckjTitUGS
RVjZhTkL3/pDOfM8IULXt04PvTXXBCm7QPqt/1qJICYrh74awS1OhJWmfwrGQc0r
o5MejoWGeL/vRMHk/yxsezp6wGpENPJidLXsEtO9V+oNZit35fOgparHeSF0XKTu
zRrXCS5Z1cWaHUBPLZY/Bz7KvWrQtVjWh023hZb5u1TUWfHX+JJfaeOozZkJ13/+
/7GeF/FgjRpeLUVgVElodDdyJrTFNwKwK9VjV8Z3SqercTvGq96ZWww1IRn2u9mZ
MO/LjrrfN3A8SSDR1C9RgPhntDUkPX0FD9sPoHJa8FdmG9eZXTte5WYXvNf2Svxk
BO/diiyK89rowBU6cVwUNoCMPHzjrDG73RbpNjUyIfSRWYrNYuJsVGrC7pf1Pe0y
DYlBizvs0/jMPnBKtt2t/+ukxDPnJ6G8wUOaTjsPlpWM5KBQvi4zWkgyPvua2X+y
Oo1A0VmyLlz5R19/Pj5JTKEwCLFt2uYhtO1ytgB/6Hx+6qqYnWMz5ruNXAUyjrPP
482DsIqMHO5IGtSRoUZn+PMDr2iM6GQ+hth+omQqjfyq+XmnPYsLq0sdVTCS3qlP
A/oE+w4g1NWaJTcysJ/ATn4xfX19lMVrtGEZnw1pbyZBAkrqWPAI3ZKj5i2K5MYJ
onfECDUI1QWtokwOBtDIHQMOMMUDOuptP7A8rPDfptetCER5oqAkKTkOcT9eToIt
u/RjxHrl+XYHOXHh6ckSriBhL6ECUCR+cfJGEo4DtQj74kJSk4VQSzKFff2gDU2N
RqJuosmiZD8uC5KMIYcoRPzJTqTnSC8Uzz0N9/s7iGM0dJZ0ngJYc1xQpQXIUqmh
YYmM5KTbFBZEI4hjeBAcHN/U3PU77UA89yW4phShSBMuwuUbe2x8FiQW6eMqDLGP
6Pk5w2U9euGynbomY3pSKzQcMXELH6HU7BibPKwfx8EmI5+5gx7RkGSA1S9Gmhny
QIkJHbHHzhBuzdU6aK/dgz3ROdyN7ncTI5p5CI2lBbCV9Gvjs0Ygj5ceYguT6gNh
RP6icL1Ni53bzfePckdncIcr11DuzHNtEC5yBAXohYn+U/u00cyL80DCV9dFaC6z
DiuoCZc0Kmzqf/S1jSySmqSwPMAefKY2FePxG6Xty1+12GjNefCjJTPh5YGJnX8J
yydzfewpSLmJGR/4/HHN5in+pUG55lG3rRarkA6OYAQ6hgzmRDSRJWUd5FQqjEDc
OGc6dCibiDcgbcqfl6SI1XbdmL8+SChdHokVwU1rjznIZrLxlNLhuj+7GsBvTtZm
G/+thIlW2jTYw6uoyr0SiAMvzSep+mIVNfMlTCPCFq8ijy5uomkD9b52Gzn+0KOb
d/QwrM58y78NROOxCLNlSDSsQYkp4VKbnIwS40vSRFpSmtdV3ndDaIsuZKYEAPS/
P7Kjchfkthz9A4jZkZiGkKWumRVSU8QZ5NbSNKOoz93R4BGnJ7SB6ZRZE6fnlr2w
kwt/lR4cUsJz45p1Ah+39rLxhUU372DaaNahfNcQ8NUCV/+X+p0/xGfqRN1e4eXY
5477Qp07GlUHVE2W4LCaxvKnQKQJygnvm/M6/imrqEEbG4XJqQzbJorWK8+ZtSNh
kVkFAEtDDdQyoO0DOSJPi5jIWq0y5e4CJhTf8vo6cp4xU8fXdb5E/pedpC3x7VSg
ZyQvqihmWaCk+7SQzkhDewP6K6yf4HKqL2yfVd1JPOOEbhBz1xoUrXKZsaNsFJsp
KYbytTDNqk2V9rWr4X0LVR1z9vAN33xS+N/wQ50STQNHRmZauj7Ipr3M1F3sQzNd
H63uPiUPNzq7YM1zRAA2whyR52PVRvi7G/4wWfr5WrLb1NSpXiODNFc+4RuOQGu4
Ecq0ACJoOLdMr8/iVE6BWaU2oslxNhgIxzwLHaNLX6rsD86PlK5lchpzO44ZcZHc
NWja+0iZRhDjwFWogZD81L+Tvn/evobmdCWO75z52KmU+h9+pc8rExgTwDIKcAWs
jXO12cXY1EPQJca6ZxtIkqzcBkY4iCE1Ft82pcAcZCVP+XqdF4r9lxYekYI8Rm69
bTfFFEFJf/Boqma7mJQNUqopCXTdLslibBAGGAD2wmgWWjJKnkY0hPJEQf+YMPEH
7Pt7g8yPNpTf17bYUYB5C9nQjqlRLZDH5BMaKg1cO+FRuny5FhZYnsQEajMrbBOv
9q2xeFPLv+nMQ9cYG8sBhmSDDsQp0FCWs4k7ZwhAFBJ06cx/NQM631GMRIv/BUHx
yqFKT5apVDW8V2NH4fynLP6lNQQMhrygVSqIRedHa+k6GcEaD3tuZMd82rpApObu
PkW7fkYVojDCFAnV4gMbmpjLzLVNYsHcGOqNUj+48fFMlIQMK7+ASy/TyBH4H1LV
WTQPuEx5Ch2tiV7z/Um9iGfwHBkN08r+h9ubZPqd4/fkdHuDXG2/BQfzKrz890Oa
Dg6jJsai1e1f8KBeBEEt6hnEGFcUoddv7nZgYH4Er+LjgABuWtYSmA2xSdr0To2u
y9sDz6vtEEaE4LpifKkzq03tS8NQOZ9/xmu6zsS5BC40B1Gy6jqfPxNfHLQpcbc+
SutGmFZhUJpK9Sic8ph9nCFCzzpDsjW/D9oS+G1ZBclX1+7A7fuMPBSRl74Fkqja
vYnzRTErvXXuEjPtoIAtfuNvcFFdR9gLokbFto2i/WOpT3T3CWL/NwL3qD0x/2Dp
3hGyruY8ieKOuHnC3lcIr1wNyR/z/ZsCWm7YV+wj0dqxPY+97xe8sSTU+zKTbXpM
+tPS+41kAQfd220C+14gGL7wgPXuF7Qa5rfmmZe4HyGdbnkACXP3T5mfy4L0ATcl
vN+VeR3uw/mR3ESPxG/vj7Ba8yYJg2tFasbgrrJ3cljBG8asRqnGS8RsTxUXhljO
XtfWcugV1U8dGmB+lVeU17RgW8nr2SvEPF3KHW0fKnlYWcGVU8aBa0txwEuRsMRB
yDJTKUmxw0VPxSXnWa/GHEMv0sFlYY4efPAxqSq2ZuEuSnMBCJvA7Oc3IMvzRxfI
R5mq2xiLUrkjbFwH1A1BKYlMiOczhkMNcLhYTGueozFdvW9Af8TZroBsiX3d0ytA
1qTct+wM/nv7M4GU+9XuV3Cue8lmg+8zrQL0mjG0Ab3ahBzScfh76WP+/zLJk1Q/
Be+4tNW/MfgrGAqzPh7BLELTelEP4QO2MUlKMjooCnPM0g3WnVX6UvfWPBTgW+Lh
QJNKjGJP954Xi7XNO89n8MlRCZGm/07SMVyBExYWfzcF7VgZBPLKflnfPMRfhMk3
nK6IgmptDFb9FUOf4Fmciqy97eLBkReF3gaAzTrbxoh4432+Tr2fC0MRRH5qMz69
Qbd6z4LwkwlQzsybZlszrGUDG0y7PNSwWWv1qZFCDKhmJxpv5a7P3YgxLFAP6sUJ
qRCWzqfoqpF3T41cvKKRi0DnHCkK9na96FILqKxvyrMlQAEeFULlN2fivsYC+ir8
10oNzjPc1Cc49fdhqdVzQxtFCFqf0WAsD0q33HQvO7wJMqIVCDBXDH52YcXmMa80
/XJwMsdII5RSoyM6vUGKDyEYFbo9XzKlf6z0zgRdrTapmL61AjvUh2aq1r39TcWo
YizTsPfO2uc4n21Q6dLGpgFT+T3SiQxGF0XSvr9M5Kxf2M4BycusO68ASe/s9Oh1
jRpzlMZzdYPUf3M0ifj4C1HB2rhvJ+95vLmyy0mHGSKnB09fnanwd5M5aAZWs16e
Bbtt7tzWol0bQ1Bmw2deF1n06KNt1oVk1WR89ngxbZJmyYCDKcNMSY2AK+JqaG01
Bi6dq3CZryzEeF3b1U/XHgLrF/FRreLfO1CuQBdA5mNgVwJ3KkQNqtJmUDAZSuZy
HtXqRD3J40ij4cJHU1+hYhdF2Nvf0g/Ff5+aDVsFyuW8LNMAcolJvu3NNSSWUFDR
3Cs95Ba8cuQRZlfsMF6hbtT7zb4yttQYLtUQ9HO9BB0ge/Go8YwJILTNBEHU8Fd4
wjMh7ht4fkhEB3gsHWmcfkLQVCdHFim6Mgh5a+p6cP6aq6krpPHLj+PS5ugg4pyX
7i1+QVoguI7V6FNDr/+yTd2LIJpy2LNUXkkux02y34X/UG6YUvARGkfO+DU8tlZn
rBgt/k3n3eh11BwUDG5ebNu43wPGAL6UkWXKgEGnwJJ8PVJ+HhiBIYo5YP2T4Ywe
cUu7WfpM2peG6yx7a+/wINOtpAJkOmERGG6WgXQEQxxk0V8tQcEiVX5zmKZSsGHr
6Zb8pHJOkPAhLH4dGNGbZdzmhxMbM0/my59dpjcJqYEewseSsiDNUTV+Nt+7YBfF
WVgSH1G9kxSVgsrFkHX3ZgAw/O28y8fbHMp2hatVHZHThHpqTderaa/xAJa6BCAY
yC6DxfpHfQ46pHmpTsXG/dQOD/ZHjg0zlDO6KTLDDLkn1DXlXB3tmWCqT+BZtL0V
1D6myJqhBw7cxK+2nPlZ6aI57Y2BvvJ00Xs3SqVwZ13B9GRfBB3JMRzdeZKVr/UV
UTYLMIsJoMM/LMv29NM8u6BX9uzyyH6v3Ho4b4sf7XhjMUPnSsUbkvMjBsjiy2tp
qhfNE/MWVD6tn42y0sYZYfucAi1LLXgYBXOlhOcPJhGIziU4yajJN4Q60SeM/+ZQ
EaC8a9btQ++2T3DIE7NQMI3acDhT8Z9iRDwO4vKAm/k7xtoAr5yWAC3bgT+gXn5D
BpbxVZG1YRfxVE48NAWK+fXXCMA2CJEuTrzo1MP4ePLgewxek8qW473rY5nbcL+Q
FE64fDYsYoUm8E3zF9IrTIZMgLsT8Tnpjn7YFLXXSdIJI9ReWhg28z7zn9e2VzEC
XlrUhRaLQ2VJlgj9t5eBYe68xgGCLf7+gFmawzkFTXfoCH1heAGk6/V+TtWWRP4+
qh5EgXAWEh5a1TIpKGgk7lmOFUh2Y5ym/8nGgqW3dKXP8LEjrkVOjAv9WinTfax3
4TGCpFOAMeMyaE8+Ygq1NZqqCDNjbQM1JyG3zVNjaqahqq8aXRQlAQZfKqqrfONS
qZ/ljNs1rs5kvo0Wq5U8Y8jS3orX7a7fjK2E+lL94EkeAlgjekIkUpyDCn2lrAoR
5eu1XPr8BJED7cuYR2BSfwo4RKQNL2p0vhKq2u1eOIVOIwdLQMTb/1eVLbU8mlVl
E2FA4QJ7JS5DDPJlyLlQlAuMZaS8eqhjUFmS7uzAZndDY0AijDqVoWan9cN+UTvU
N8iE9TJ47AKu0/h6Y4FlMaZmyYxSwz5JDZbNI1Vjf2KMtR8BlXlMuGrkiTGjb4yT
Q1dgDd2x9QMFgq0/WHSpy2FCJ/UntvG6qLhNUtf1ev+8aY2mS1mPZo+cK32cj1vd
TlKlWr746pJgy1eoR0UwoExSwk9Cc1AlXhgfgrvTmI/HhQbxhh4an5xrr8Aq37Xr
CjPVfQMrc1e7JgGkTKi0Sb50x0kc01U8p3/NEUw3HItfdb7oIRRbP4nMgd4+Q4sg
zsaczvpX000sl/BOQyWPVQ4s9HZlhUsxjn2kTa65/9mZ9xc+RDIPT52nq1eZ/WtW
70758Kvhu6RmgzZ6zOCQQlDmdDTJvrPJcz1Zh2Xrs+LzQlGPdG0o46DTWZaf6xov
954EQ/S6IzjDGxEFx9KfsLdtcXrNrxZw1B53f9UL9DRy8/0E1ps/Q6qxtz3jewIc
x82Gc58v61mteaXSHJax//QBxvpZrIw+mX9GzSOEP0V1iIDVf4YR34DNdlHWXUAh
4C/sCvMyvMBUorb5IuTu4u8JNuoZICJam5Sj9nWGmeT55m2OBH/UEy5GpkswRPDH
d+LSiPMfmLyi1JTyJGbLQ0XvhfFd0WxjCl+bPXyqqa2FSE7g2bKSoy61/XeouNMR
LWUP9mHiajNakE9HzmEhiLk8ZN1qKTzCm9Oo/45LiztP5EbxH4FPEmH1LcS2sly2
jemZZWoYjqr/elcNVJuslBhOCK9b9WeRzoSO7bh0eDT9yYZTH+N8WkyYtyXQnrtQ
kg3Ow719PL0qIe827ANk0ujd08i7SrDhVkVEEScKyD1OubGJ4IrTSVt7nbu0PEke
jUjLrMSvDQl0Z6oGkELCqz2fVO8hgpRzJelmROFZVNE57dfMt470dpp+lJ65Iudz
EL9tbA6h4OcEjNCDq09cQm2E4MnFgyvScmc/iDGPj2NE8FLHyIJsiNzmzqTtu6zo
uLK7UEKLcrrlsHc5iQ3HbJYC0C/3CeJcpfOUQ19ODJPZZWxEC5pO8hm7GG9sVJPt
WG+ym2V+8WeNqGHQAhkrXpFLA1fDbvm1h6Z/OdyiRyTf47L4QHYv/pv3D501xY48
83/Kc9qH1fr/WhKIuUz23ZeX22jHYE36QeB9ZBmmU07S/qcz2KJFsSkJArL3Ku8+
z86ZTyPg32tDP0E+Pzvyz0mhOCPCZSQWVJhSzdlwRBAD4APjcnWhsSAMHqmufbmR
5haLn85XceMtnfz6wXy42F+aUP/gOtysE4a2jwZzQDjNpJvsAqzDMvSHZZonke5z
34afSKv2FvuNCJWjt7TMIGo4gTxHaJI7CRsJ+AKppkYgVHwWNvHUy4jNJ6gNIVCC
Pwq/nphfQQEUsr9l3EIR/S1bZ6gyGB6UxwuwJil/+dQrirxUWIyT5YrDgab2EmdT
n3RC4Kd28nnJDWtQBo63P8U2jv8oPsr3KuOxYqFRfOCqg2ZIpQ+HH13T64mfaMt7
+9LlvaflFumsH5laQPA7LppRMWUrEoAxPdm4JwiaFbKi13tbYoFY4otvM6bwIcYu
Ukqd7jfJdKEwPQzPO/2YEod3K4Y2khpL2hUiZR0Jp7EsbFoGs2yx+CjpAZg+cVAt
5IkNmnekY5Xy7n0bQm8NC1IQYSbtRGrub/77pN5Yi3RNVbdW9Y8A2QVwRuUlycoo
r2OqzfqxHbfbhgFhX0QUC+Wj95Qjiy6ZnU7BAZuVPujWwPcADwOECA5eVSEVCNG/
tCD1tWPm1E57hlIKhRYoJTyPo49HzbRRPg2yalDNU2Ouwylmq5vNq+D/28UAgXe5
MLJdm9RSBfE6kXnYPatpzlz5VCEkcOwdqEE91mdGnxce1xPf8AJEFFDJSqNOL3Q4
Eryh1Cc3tA3eVbeddr/LA0WuN+XbrBldmzxN5ryMQG3L34h+Q0qXJv/NgMNw1KHh
RZ+hunuMZmM1345cZN+hZnmjs5zOrlU403SdxDueX0iOwC8XIWkdpFhlou72IZlR
zD8D2wrltPILiq9DNcwc1iuW8ZjL/oxnas4ITWhcWnF3q/J+JWgFHcOKo9LUR8AB
WPHcuf6gKpTPtgm9tuXukhnyuRtMF0BcoMo7PrEhw7JO2l3HFAqjM76t0iEWKczm
Ar5NPzyGnbgJp0q4tdvEKqrXubbfqDzDIa2Ix2cmZmxtdtzJDVEhvVTUWCOcoJl/
xcIp+oI9wNZj9p3ZzGoHtr+GNQhvHHGLh6PVssyrhKRM3+TeoNG9texYwC+eK2AX
YYCq5T97aKDh/QpuXPgEMc63P9/uulmgbXWMvp4+/mApplBrwCipJ0vt1qxQ1g22
KVW/eK2iTPWEyJvb6488UkstM8FCRD4EWatfO41vgavCvEudbzq/CpDmJcn07YQx
HTxPB6kpa+I+2y4jz247SMYQtOwFfWYIdcT2uyUHzI82rqi5biCCbigVVFP2LEI2
FLhvg11ne0moQ5qT7rGlUeY8Bv2GW+TvgqHjfMq1jW6XPoxfgJifXXjlRBMNxyJ4
7eLoJ5RrXGFLEoyFSZfKa2wYQ40x0ORo0zevQUj0kB3C2SBByIC6uX/MMHEZfB02
ULD3TgWMvmftN6NFGBAFfUZLTWhjhE5EGhXNDOzeP7Lc2DlYH174GUptFg1eUgyZ
l3BiDGnyZnb6vSB6VSRNOu62VREcHOzkYXREAzLLktfcJFQCO2v0nyhXfbrBrPIR
AHiprnlmnOUWAHD8f6/OPDDVfXcIUsE9DWwjgH1ycYLpZZfZWmW0/FbyFAdC4TQT
rI9YOGPr6bsZDRr9v340tP55YsGeITVGyw+DXeEWLYs4zaKHXJXd5TgsTN9P0Dcd
RN6+qFTeelWiy3EC1jYSXCsUWzF+EamtP/hfK1QWB+CChX0ae5PGxBUnpM2Dk+lC
Ms6l5u5A66R6U/6TtGkcNA9mUg78Pe6RZZiJp0wT4OqXvPeVIwvbauDQQYz7alRJ
k9P9DVC399nbZOezRGAjhdNr9Vx1FlXgABdX/XPe1/WohcFJSAcpsYOd1cS/WJGB
8U0FTt8RLHbU+qekJVIUYXV0PH7+fQj8iOfNexUm96QduwAxpysP6vYI3lFTDmbl
+691xGlgQwAWgQCb1Lg+IMsW5O25u7XDqE49xopuiaeo7rSOpRyH7H2mFlf/igI2
752+exTaraNg/wRDStRA/5PROabHXaKuMYWyxpzKh6+ouszEYmZlboeY6wOwpipN
ss4XbPQyzvemWhGY7xVwcFDZuSx8ZHSSNZYu7V/nrZ/90/agY/hHggevArKK1QfX
YDqE3nmAbzx4qTFidAkpIyfh8UOKLZ6xJqsnRzfq/IZAwtuMsivUvyVlh0ieACIC
kCUj4RaoR+ADQ7usxtVCzv6mLVyxsIoItGIyMx4D2pPqU1CsNZTn9uCstt/eTR1t
EtaBExAJfM05EZeEzXQ7eQrexUGW3mXS340uNygKT+2O978/YOIiAEhe7vKFtJjd
1K2Hh0wYi/4LwnWD4ek6U3Ie3ZeO8HfAl+hlIBAPqm6q6SVQ6VN2rvfoskTVX2bI
Igm+YqWlerigtd2kRSSRntN/nb9t6qUxzfdzdDyt/2Kluxd7FJ60erOZU/YQkZ3r
yqMwb5JMoenN8cuy/yb8HfSrP6lQPqw+Tfxlut2zFWaowVecpOL+6N52pp721Xv3
quPnjg/C5QS/IEhxKoXVLrxqt5L8GPuhe5QZbSaaRkf85+vUQVNiGXn55tYtyuHW
hPA8nw7PL+Mt8j3UKPGWI3eAsdId/L+NzbzTBuA7T5rr0FBqvJ8jdKARQ7Q0vAxm
8uwnv7iDNrizS+3MnmFmhs5CyP2Ush6kF/UY/+sC5bj1r3S7C4MlNy7teKwB3kuK
v+cqptup2OVCX7mXPqhYCQ/kB2/blbEESs8y7/01QMPrxpvzEtd4MFTmCBm81bxq
RCmnHIyE2my9wHmNklyzyXXEIWliyzBT14Eoypwd/ueldewuWOuJs8oCTP/jTA50
bMw0TJ+EPaO3JDV/6ZW3UmCzV27ljPO6M1IKUfgNwKZWycoNiF12K8ar1ryeBj+1
aq+npFA6cj/XG17+k+yjZaK83oWz42Ggm0bILj5GjK4=
`pragma protect end_protected
