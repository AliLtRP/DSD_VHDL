// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:15 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qp5nqM5H1WRJlRzJacagRnouB3+ho9KC4ixM0gQfkMmBNSYqh3ycNX4jSNA23amX
euYtqYwon/mY7RGK7rOgjxQ+X05dxrxl0WoL92dqqU/acbgU1e1ZzwvmgM+hG7ND
nzb/ysRZIy4MZreBzMvqRTIa1CGDZU9LEEF63besSg4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11120)
i1rMQIJ7RTuYSJO/Fs1lYo5ziDj+KfGwMD5kIRqbi67hOR3S+me68FcmoMfQDL+L
Kouy6cqkYU7Fi8xdON8jZmlAudCPa7Fsr/GN1sa0E1lvYGL6Hk3sHbE4Wry2IZBm
gLoWhxW1QakJjbymkoM+JTVHziK7qICSWdoTz8TSE7tBXclqvyR5HDgv+A6KUrN3
IYThJqpJtG+HW710mCV3hC3THsL2iw4+4fMoqGEAP8RwdI7xnPOcrhQSYai083MU
NQCAaGL5nafy9cl5sDvHXPaNS7VkiLYuFQwh42cbvBNOywsDRRi58zjuYKWYr/Uu
djUKVrNG2ZZdpEcAxfH/h7/gpUEEyd3ny9oJY3IvsxFUMX8qU+MmppqSquJLO74v
XMLmVvt2ZoZWNryfrosRhe7vc666fproN8cEAL4JdZ50YOt7LyQlGQmn/sR0MLeo
E9Mw9HwMb0LRPk8RzxuGpiTt6Zhf+MuFHvJZfVwtShL13lfMh6bM89hMiagef6Yd
qsngES3bf73Zmt39ye5Y7azrjkkrsjbmeOiT8g8a+67iWff3xC31Kupt6s623Ca1
JCHVmI92L/MpLOY/Pd9JGqSJUN/jzYHUR0giMGgsY3MumViiE6w3PVNQn9cu2vRX
AjkGy2LaUncIpPnIQPDP7dnkS5LGU8evpKRi67mAh8DDZTrEXKIGYkyQR8SzS2pR
bTwFWfDbDWJB/iTksCFy8eIzLUwb4UpnAE2toBYv4STwWzmIuXCu1FpyzuITUMtF
cR0jSrTLV1V9GyYiZvx0yHiUWROz814bT0EjUm/40bDn8JHrHqzyQ8MxsFi8Ggnj
6QxSj/fyA6bSsjB89P5d6g1aluQoGw1/Ji8bDQ1zZyEM6HtVvdxc8Hro4Q7vmvzo
zWsgwjlGCpxTuTXn8WzZDSSD80FT301xaLVaY8vnzluB6uoYSfbRcH932GwPQsE6
r9QASb2RlC1NIfIfCkNraa3S9kkx0ck78bt8YJ3xQNZY0pExWjWAvV0ZvUQFvOsE
+ybQ7nyKk8SZlj9IoGgVIJ0b+qcqNW61V7daGkscM0Iss3oA4+IMSgloNqRP+5Wt
nKPynJkfCuewKL+2UL48RacktV2IqCwSGrZAa09Ax4pidMNiei40zmTTaHzcNFBS
aVAOTfOqudw4qG9SFo9aIMkZ1F+0wYKes3hLdMLY65zfEzMijVBmRULam8f19rER
5nxWOL2QbN0eKLOIEU8wm8UEAqWGqxvZup9pYWP54ur/aIIhSkk3UjYkvi34aqon
tzt19nvF5jNeYzJJXDPfYXKBLCULNltfK9NIMUBzuBLuGMFJX6IGwiH7f2P2vXaz
z3K3FuA2tyTKv8OAyfwk+hyOG99PbjuYTWoBTuJMVdWTQL7b/aMudlCCkqdn2nUW
JcxrK6GlbCJ+LtGVdAZTJRUA647bDabpqA6ujthkRh54qMU2rh4yQD0Wc1FnkJkk
FIvKquPatUHfbemf90oKi96d4q1rcRY70LzhHoSFhRI494YuvcBUmN+02+PYynUv
k7OHtnJtI6LYrjOWf7nghJEfGQBw2FYyO/DpwySfD1NwMTTcn6DhWg/nm98U/dRD
chsK1EUaBXZt0+Rqt2S9ouUYFM6V6s0tV/CdqOfRlIYoTW6hPyjJnQYmZ9nP5mG2
7wmbPBHVYNU1xOemMzMfl0OOdPzKjzULWLLW79GKxl7lAt8JuqV3hpMCrwfeouow
yTUKgLBi/jrvfgqtOAdATQqCkC7K7Q/hafnjzgePut6rr8+br8/+zRVviQEoWloq
Zm4oIJIaeOj6EncO6rGm5+6BcCDu1Zsez8OhI51/TTawrKkaGY8LbDTice2k3y0u
cJH+xE63S1NNPo2serH0fvPC3e6EKbJn7fPtjTgMXpMqLBmx1YzJHHaHMY14js5v
eN2V7eBy3fxNOlXAt12iI2/f5UHY4gESmGMD4lNJJbBvKrr1llAGMxNyG1+SRE0W
st7PtxF0lVnBppW6mBWJmEg236zfxNInP9J31S07wfV/5g2OBZ3xpWYSGysQZyhr
cKd8s/yNBTfSjQ5kIWwfkV6z0PJ09K7MO8pjtAa3iAj+CpF95XADnmwpGny2NzzF
U8LgrDEQU/Y8kpdxjPUZIJ67O6cuKmsWxrbew8X2QNAY3zplPPHb246qZ5cNfeyq
PKy9rpwekBhP5F+ZjQc/qRbxL5jknDmQfYDDDJ2u9tgZ4Apfv43gAIK/2wWY4LUZ
+Yk+6rtkQLqKmOzkgY/OSCyYIRh2/Z90e4AoZEVTkl5C4EL20O77MWCRR9LrKcvr
TcikJr5n/BgjeW263vmyMtcQAI2o69hMRZSGjFzouuntSawnbOojBwvT51rudyJs
BhSSPwvmSdLiC/x+6t7LO7ID/TYQNLwkGmYTpoNSPUDdOQw33dxVbqx9WZlaK4gY
TO3u7rGyLfhSXM7b7b24CudZjJ0LH0KGR3MziaTj75Z/3KSo4xgA1FBGIefdlz9T
b2vpS5wX2T+Nd+b8MHXhdua6QahoBitsLYAq7RQ+7FKp+uYNmVlz/+gnc4DM694y
2fQvikOHfbjdPjdY3bi/yBUroYCwkQLLo67M3kPTSrFY05A0x1DAyrPL/gQ4wd2b
7Kostb7nXgLJAflfRQYwcg1jjT0tKhWgljcriFMsEc/f766Ca7QXiWK68iyWyF05
8JDMYzEO2prp1kpvZImESjf9Edu9+RgU/iOAsprmN4MSA0W65hAA5lqeUN6QKMwp
AreEW0fI6Yb78+Gi8Hg+SF1VQtcMdP5X/23IHW5OMyyvYzdQMunlsf/20k6xCjfL
nOGcIbBgQdaYvxw2ImoK0alavKN85rjQYLVCEtFasJ8ugHjWbyKpdlTbrXk0jfoQ
7jbK/svf6684BPaxvddHNLDazmuF74H34sQBYy9G1JUQ+gwBxjFqGVU6Tu8oAeX+
ffu0I3XHepp5daXgjGXcmTZi7UHFqE3teXSnZ1KeRfz+sO/YFgrX+8Rnj0e+tzQh
b4A0BgSvAVWhpfS+PrZoA6YaSa6gLuZHymqNAdQZfDtHD4RRZe9PNds2PsFD0+ff
H1rupAtQR+FaeFQfEwzl6k3NuQ9Betmt4qcdV3PkEDCPozu5Wlq5DJpNAvGB3reJ
rtdYE5MhhntOmbZLuTeScTDC+RZWk6OVVWDnfRo8i2QH+Ra3KWPTu9wYyzxSygzS
0h66baxhbxUJexhNqqi/l18+GrEk41Fn593ixKvVPreJy6rVmFotyACbARsnrHe3
OEBs6TIXxvpe9Q80ia6QOYEZjriZ6L8EhwIyGgjjB8iQbsUfWoUGJSn6cILrVI0K
VDpoiI4pEK2HAePnAfYQAbJxLiOgI1TbUBlJ7qem+OKRrVQp46/+0w7utgMQDYaT
iUh1mDSFZCrN3pvAgb+Wx9JVgrK6XwlpERuFz8blsDdAubQQDDZebwNcA8y73Zl6
+PFgEGD2wcmhxDS74JQ1CpKSnXBgsIhVQNE5jmahNmTJD/qWEfqT5nvsDXuKsrNT
CdkYb3OKSge+jsxrKnnSkFJOJoQVv3G5HT/XF+/Rz+wnLmtOq77lTpu7L01MVKqr
im2L+WiJc0T9Rc+nqUsSTlglyncXT72mkUAOi4HOkef+eVGmCgmF85JiRSmDcxI9
wdsOVuz5lHBFqAnYi70jciyMBLn4tW3nYk75GOIqMyFCMvAWV+sB+bymM6QyTQVl
cwUbrT3abeZiQwGH/CUx6qw6RA+KnQS4hDpCmiEPUhyTOvCv1xadoYOqHqUIDoTI
6bFtO8droACTqF2ap5DothIupeYjyqRqMd6xx8g1m7LeWWFSWcYAXsWEt+NXgqDI
jBE+LrmQ++UsWB5yn5eWQRW1UD7LzV0hYOGh3EZ4KhWV7oxzuqQN6bfleUPCEPSg
Me8+gQvRym/0/nlFwJjOrRAyXnNKJ65G3tiajhpKAyzgvUzHlBMKLQdEkexEHuae
NkxaUHecZll0bnk6z7FHwkHVvrA9QsqvhGs++MWRR2e3xl+Zijj2k6OMo3oBmRkE
mifzr/2qraBBRf6PNbmxOZBpAngvYhLz8dyCkM7QYN0sTaFjbisxmUTMKTpZbOCj
Wc23tNEH5oJgvvzcDlFzOKriPu4mRq0YYdjipiMa9Ulz93lld0aH5FVdx/LauYi8
ReSXBPCdhvGXaTVGKqeFUWWXJsfKTEdZbT5/5y1BaU8HMFZjO+JvBgZ/2PhqSC/q
NkeBYX8FmDHH2iWw9NyBYJOXO3xBQVKKPJ53DduOjhxVmYz260lkrDGqQjrcptS1
6mo67W2DCyZ6nRdurF7Q+22jeGX3Na1L6wXbjaVt2b1q9wLoLn8GMkx3epZW8W9n
4iCIf94Zcv2z0NJ1Tfw4KtKCfI3GmDxUKJ2snMNBnrldOkQUxxOH+s4sROMDqwNl
C0snTEixzrHLHP9TsAeYK6PZi5dMXF1fRe6Ly1wKk48BXpYeo7t7NyLVSxB+EDyH
jwdoGcC6xzNCwfcfdVZ4SjCzItIKrnQKoww3n2/90hxhRC5nB7SInVQAUR9AuegT
Jk2Pa1wDbsdeU0Ga5bdYinnXtpZoefIBfJe+JGJYrxuQiZDNvCOII5Ah50e+WQUx
Bbp0BxstDgUSTHkMXSonjNhDM1hp2LJcl4loHcHMVySP9Ope5XKihdCZn14TELYi
jN8GEoqKwl8quP0M17WtRzX2c2fESdZJ4CO2dT9aK0UnKfPdn5Gpo7wurPmyffNP
SHMlPSeJXaM0WQZJS5nkJcv14u0vL3a1Db12KbuA208qryvQZxHHLO9brGE1CzhU
j5R4IXRYBcu4F7P4ZK5qe5Jebr8XxIHVHlzErzqyR/pEglZIx1ONzsvzAaNgWIUt
XiGKI1r57yjCwp0yaA0GPFe3ZeEYpDcFMg4Db85vlsb8n5MASf0JRgCabz2FIY8Y
cn3u5J3tfgjexIC9qqXwCYBq8KscQLTT3dZWaeR1XsIaI34IZyTzS/hkxKKiyXEO
KUoaiqVQxUVYDuH6gJtptLMqobf2EcPWhTP6feUD/oQrQULRof3oMciEW6ZczEQQ
vIh16HQcR+orObEztbWIndc0EU08D9iIERSDFwLrmpb7UxePAPPkhX816SRccFPa
PqSXu1hqyYgvxR1xUwWCwb/4mfaJP1+7PjtzFCKhzbu7orICnJyY7NlgOBzjKYI5
+ZqJsdcXWnw16J2royQ8I1ePN5qhw3gwSy4IOA9elkVv1OOHHSAUbSFX7fWOK2K2
4eYCoPGfw5QXqDrGWHjqlL3e24c7cZ3F1XI9onN2cHX27mXd0su73MiLdRSZaPRA
l7pN+MD8xeUpkzleb1JtDO80bb2uD9Y/JB3VqB0lBucGPPXZNY/8zj6Oj8MXYATP
HSKz3LR+ah1cCmwwFNrhjVYLheIytYvzbutb6r54sNay0N3C3l0pJAJFOtCSqZTV
s9ccyWFXcPfTHvxTqW/3KV3zCT8gLajzdMlD044aovcJ/D5/BI4ZjmzopO6pF2fX
soRXgk5TlBOMMWj4yokl04iViDC/ChRJPXpQLSew2Iblq4qt5SOKYQv012qRXveq
PgazQcZYoLJWdwQUd6zCZa6GpEizrzFVv0FwfC+lZF3rHY34vkM5dZbaiGvfPTHb
P03Ydk+Uo3gR7SMsIe6n0sC8ZWkCJpRFLGivY8tU5w6eeoS5VIQo3OrRhrmZlnWG
cUGRdJnRfKzWQNhK/K/HpDTUuoi7T+OM0KuZLNJkAbl0wl9olCkHrr72X8lKu0H/
7EFJv7mqtqEEczJE/al7zX+IQ3ScjRdzDfbbeH+wrSFU6KwX+/Wejh/OkRpoCV0L
OJ0NpzLqzDhM5IjhKJYRgU8HIebLblJ47ZzLUgYrYtq5cHhl7/q8/iBlHYmtzjpN
JFfzroGPdLEsvKmCAgzAXij21ESYrMs52CEJ6+zxSYM/3O4tixHHtxZp9Fq8DfBv
l5J7JOpYp9i4JqCn1s2pbwJZ/s0AwQdnsbguJYLO6yfjKI6GuJZ36rQKzRX9PpCC
VMUYsPxWQ0wACQx3bxDMtpLTZymY4Mkbnj3BUOKtKwff+DPbXXapdx7/ESjEtKvW
yNJTnCib0tPRt5Vd/y2owscChpNb6cnESB9aJgh90GIOPWteTv5YAn0Gxe1xwiu+
LlmcdqzH0BX25PGfVet7dU8eT617LBZZKDdqIc+JjH4XCYwJt+97pTEben9rUn0P
sNGtCqJPatMRSuq2v+bhocTS6ePnlykDoYKNLr2pzzcXSR1+uAU05yCiiVaOQQVB
+xv+VpmdXNlcc0tH6S7P0bh7opohIGV6nAe340EzGxe0Dv+tB+uEUuYYpWAOQg1J
iXgiXTVTwcNaGuKfHi4WdRySmDa1oVTDXmsFkxGM1g0twDb9SgxMj++XHhx7KqMO
2EWscdDhES6curWQCxBBjFLlj6dd4y2AbF6FIoaKhXEwEbufEPN0j9MQpSSwgX4h
G0TbuwESFvTyACIDNE5Vp68oIdw0mLnWI2oJi9OEEgxSGYXaTHKNuiKocJpHF7kh
kSVjaSOO5m/PHWI8TtpMV5OofxUvb897Ob22YBUaSfDCxDTLVTrbd2cv9SQtzpVF
rOmbnciEi3CxCVhXK7CBoLQ4I5KRyJB9Eq3FSz91N4yTVBuKbB45l4u5w4thj2hz
7BhvPj7/UYmISRDE8YFPTxeOdBut5rXjvJnYu+HYU1XovjJ354KoHY/1dUww/nAu
HoDKgrkVneeE6Kk/adZ7lqBDdgV6Qa9Zs65Oxv26LL9/gk7Z5gp6HBATQcHUq2Yj
mjD5rEPbaUd2eSf46E68oy78qMsxAQU7eayq5sS1IrTqJ7wjOeqekITXTU5YwYtb
Tksf/OaOX9TUF/g42JQkc8AWwqj7EOZ4m/PSsS5qvtM877OD2+d0rnz3+LjtG1Xk
DstKFT6O8TwVOO/AhougvGQ3eP9ldYHqCjfmbaISpT8qzaorluCR0oryqrygY41X
oiI77Wv+gz5OryVnjmjicJFGWejqoWlZgX8ZwF8nUd3AdjA5hXan6Wo/k9ne+aMo
Vq0QHOJ8/hm94JrwmUyNN+i9woq4xK1PSfF1bWGQ+ahDmjZwG8D4byk2pezFgtjp
qKlmeLi4swlU+IZo8sayhwEqQZ7VyeHbfcwFulorjlJhhY6uUVy4mQ5n7mvc/zZF
RIn0gAVB1joHYTqAQdfYX8m5VwBic+dFfZG9DCd/bedKJpRuFDCBZW50GF9kzio/
Nd2nnZok7mgD8GGGNyMVjyReLoS4F4IuTC6BK8nK46+hLf37xdIz8IgBz8Eai7rk
xQVkrbx+Vj6FECUJt9hhMNM2L7QNyrlew2yhesXOQYcupc5tGmwzKVfGyzicW9kB
TKnmxHv8yX8u7/E0K4Ln3jMe+xp6orozIt8ObNF21uvriLicc4WkPlXG6GdC3urw
DhkqC5U5W/VW8z2ixGU02bVPfpu/yzCX0EgtJdEAX8hR6hX6GEDXhRn+mN7TRxXG
gonU0s8WTfwvdefSz4dCLcym6n5b//9jT42dWI+KY185GHXrerY5V0XTmYhH/gki
I+b5gvTMHBk6HtWVBeLq0Zx/hjgekG216y6NeFvt1HxyXk4vmZnB3aFQd8s2Kz3f
dNhxG32GKec+irnfxE1LSzsaJ04Q6NXarC7eo1eNNRK3XlEJ5hMsk26dmidSZmRL
/FzV3SP8aKJ3CCpcpG2VSpVSwuYyMvriytPTkEDju4wh+AFwabT7s4anBW/eoPVC
MCPXS0shjlaI+AxzJLL1Q+pxxFkgw8qsWbGi5ZY+S4yA9/W7cWGw/LegW4E2Oxl6
r4HeI1kgyjP3pS8sd2yyl6C2pcP41tohypByLlARh8D46uU5BNKhH/6x9eDpnF4D
BRJunlCiXTPenMBMaSlZuW3WezL//QzQg4tSMI4XtmsV/vqrPvfgCidAXk3caQK+
H/0Z+TdJaPiA1DQGQCJRDyRqlnk099WR5ztvXW6uf/mF8Pz6ey4yTzJ1ocA55olT
pTkEjO9cD1bOmy0VodHJ+l0oAAeqoaB7GHxF3u9okvJveO0FgOyyLeZpoJZSppFw
kHDj356GtUjjRU88Yig/3K5QfTLhEwrWEB947nZsuHUyJmQjpQLjnvh1tkYKn9OK
KyeYWtoNETjFMPbsCrNoHmKeqXH3r7hCP6U/bS9lQBouMV3Z+mXBMXncq3iZUtWC
7zrz1n/6Y8f8WZFdRVDAFJ7J2Oc+H//DsKMvbylxsp7v2AvcrIxglyz3/eJCdp1e
NhUA4yq+ATloftjBp1+fs6BJNtxT2zStl+iia0rCnokc7SxoGv26eaXj4G2oG75G
XrsmoHFG1kkuBT2mkqo53TUJ/J58p+xgagAVSGqurUs0rwoG0vVK0TC25FSxkisc
3LRIgUwbSYX2GBokphJgtgKgDfAwTbGkDz8+SoTgEjnZBKsNGUtEeq5Uqg8maqcn
HxbKOAYAKTsZ9EkdFDJHIkuY5OZCpfOmBeKBfEyOEgXxtcp5uJ+V9dDkrAy8yRUh
1a4EOUmWljfkdS+e3IA48SqI0N2VmuhJyaU1ExH5MTnpiwsjl4TfW/DxBd93QZpx
jf1D0qiNmnnPPDxqBzvGHTI6adrffvRxkrTWI9F8x6NLcTlMnGCd/mvODFN2AtgZ
1xbWbTxvxOCqNLDlpvRHDIeSt7RZx4LD87MIWKD+NZZwy3N+nGZKFGZSHHGk3s64
h2mdBmi7eh+b8mLUYQL9wcrx47OCRGwpUD87E6xz/9Y/8+5ixHDtXBUQQ1BqhmQb
Nh6M+Ba726F6pkpwSrW1wWnwImTFRiWtzzEFqqb9iJ0Jwjse2jPn2V++nWGSkQgS
A5O0VXVs7ttoMlHRxPeDbA/XKvoDMXA8WVidaK9VSoj1R3ywKy+blATccbFhlMbN
c3fieR+yIdvP0hnU1RPV1qB+Gr59X42rTQd/Louf59Bu0SJMml6rk+FhvD9LmucN
1pjX5tnsZjRUwOjrYkmfCBtGjhpD2EgY7d/mBlbetZwpDXi5ZGDOKdJ43A/4OIVv
15ywPjaSEcaMMLYMX9zEhrp6WCCes8ZRWBR6FrPPTs1cQJc5LKpbFlOOYUSPQl72
n5cc3epgNAg3ZlEw/qk3Cqxyja95sRsCdjhkuIgfqEXhYDlnl11YZG+GNBOLtD9p
Xg4ia4MNr+ZSrdRsz5+3tpgq+J+wHWTv+MU/HwvKIlZ3fUeFvRjMjd6HUn/WlRaa
A5mXkY8utepxns9f2tS1RM6cFDXJJ/G0SFg3+omTJEl4Q2+1saapc+E9nB8BNd/M
vOKPHygF9ZtjpyZaZChUOpE8PHrai5VNHAzU0iLrjoFt4stcHVAAU/a7ZfwJz2WU
ysM29GAJ7I6f3j9QWnrkwlbO6uk+pcp3IpVpgIoCSkVzHFK04VL6pEBZ4nM4Gmw8
YBhWMCcFTWtxM02jM+Y3HDCBox+E4FNUplwzXWuAIgCoY+4WguCqBKUqVu+mUKK1
sUL/XkKYglY/PSFR6b4KNoAZGBmqwDkLsBnfGH2Poog4nOayUtvHTnUYdGoM6Wmj
t8MRUC0A3Sz752+kGYznY2QGcM+NxrULL49TxxyrpF67dxKhF06a7WcuVQKmydri
sw4c4YOWAG6Qou/O3gVMYaDoiJzGL7Vr6yUaykPuZ5Xp7H42GgS8nZkBebLPwXBW
cJYC2U4tqsbaJPZBCM7zLcNlPHxKvtNPkoSh/eNtNs10UTv4VkjbvPFxZmmiRUil
Q79ih4xdbbZrOWJ9B/h9bWQKgHrFSBtoQkSSI8UIBppdfn22OZsylJQwYYwALZHI
QoQ9tP0bgmIjeSSw6gLVo7ADNVfpHrJJ017dYzICv5mgWHzOj9fntn/i1mIwiIss
Z4xbOFHnDOZjASFmZ0J39ZSKN4gHcJ48UpAM3nip4/x9ZRaYPHVo3ez1dcx9yYG8
dWBndd+J+4CWOUgubHjGMD++PkR4MXuR5eJoGhxXj5uTl28YM89hPQIe7rggAQRw
GK7tCnxtnzjv0C+8E74XiHJ5UPW10m5TU6yDN35wM34ez/TmWgdHmCv/YGSTT/w6
u/BjOkTLiSBvgqfvdFL4wqTs23lWv25ZNNGdd50CZAo/kTYy5bdH9vTT+0GuV5q0
haXZ55leaEO4XGMg4xiS6TKahK/PZiIy7TlceFTqBRLcmGFQ1d7J0B72Bx2Bqk4C
wB7hPhZtga0rJ8oUvK9RSAgX9JZz3Rb4ZTRZnzahvgwmVehxrXoNwhiesyLAfxAL
pfMPXoEVSYsSQDBlX7B6C1X6cUhHtBNu23tMfXdNCpPkpc+/WeCsW3gmUKZyXEi1
pWd9GDk/QKfHO7rMBb3mkmR7zOjbMI92mnsW+y3CrVMwu/F5cRFOVY1quKhFEEUD
2BGZ3cDuTvJUSmPGGSh70KstmnGoq2m/Z5tio2W8HsV25KZLmQ+fpBH2KIb9fucN
INJW0gIjpSNi1ZNXThWunto5ehk4G1AkFa1RCBPxqo9qfnqBeqiieFQRrzMp22ju
PPSQ6u36kYdpAFMIuMV9pDrBKeLC+3Gl2f3WZMn4I8jEJUsXomS8C1bnnDl1A/H0
nwj+MT5XXFQ1bEWVx8dKSL6x/5l0XMwWJxU0uoSEyZyZwcUpzfuTsrD4ra8gMesC
5ccdFUb3lLHHLvjgWUX7XcN4obsxiJ3pX0/I3yVPy7QSPvACX/WjNygzfQQMyMu5
rWInfAtmL0WtudiRVNx1bY8e/h4Ghqq77QWeTISiJAQ3iadX0E75cL04unsW1cyO
db8STgRPhVBHfcPqYVVaXO4GkdopI1LZnZyGgD8VWsOONQf7z8hHti/aTFkHs4sT
alGTbzKVhdYWKx4osFXw9y519rhVBp0TpyunSniI+oAAUSxeuv4d95JmUEruC42D
PpKNB3a/2nKIEslJUmZrjCnTwhiS1rdQNwfjHBf4tsGYDujkgtmEJpA9/0/2gIZ1
D31PY0J20sSXN9jKoGL/iU1n8HZtadPzLvOi1DnYwgpIXafBXH9SGYcAH22pvcmF
40TKNAcRfFq4p0t5LVFy/DS0+6bnPclIsasLvjmzT2bksmIwX7NnimjaG2q8mplS
jS0Dz9YSw/0FSW2bIwmDE02qLHifwQ8QEWwofd6mBrHn15CjYIC8tHTwI0vASDMr
aVv6MFe6hEZeDys/O7DeoCAWMqbmcgLYNUcqpyz7o3CjPTe5IRfZfkFvOG6ph0f2
xGTF27oieLu0U6lt4XhomR6j29coe8UNigaSVfNk+ZmAfLJFJnWA3eTkORZH68EF
x9nUx6X9RIZAXq/U45I9nsgTeQA7vv/4fbUYfR58d3C56gubS1DsrZjrgadorH71
JtSDZ63CQ1dYcPv5vldRQshTj/cnKe4m6SA5qNFXYPA5fJbcevI2pEEXtrrX+hoa
5XZqTH09giKI+s+3UwocTulUlfO/oda41tszTKOn4S2IXBzL2er+UH7yFsIg5yMs
keyZQKkkO1co/71J0e+Ypbfq4slVzxcBwv2uyf+/D6lLVIw3RIUNNz6Hs84eJevu
pjTIKTTlz0aERAuN63yRVQyk5sl1y/aYAb4ZoJfPXMeXNpOxSH7MEn0WStmtMU6r
pcYQn7yJDtF9Gmg0KcnqdNgGfWorEorIKlhWkenFxkzPixVVWNkjDz48UhIJ0QLz
abItqKEaQAjeJK9U3yHRY37mzUadKzb9wHpglOpWNRjX/M6ASQpvNlGY2x1Tj7Ei
kpXLZUEDLB0uFHYb++2dn2ebm9kMcX3xoFHRBbfzlcM0t1YL8ZmRK80wKVM4P7+a
XO88mdrMUmu49z5+zQDqsidB6oAVU1o/gicR/yWOH5Rc2RA3b87Zdpri9lAbOjXI
vcW7vneFvOCtlg7Bk+EKMCVpFkH7pulkkv7KVerIXEo5Ny2zwUGptpp7WdZ8/gj4
blh8ecG5lqqvW8t9L39Z4ijPG/NTHpREYrgGzGSDcHQ+JcqkAXglYMtua6W8wPRP
nvnCE5HtVYGvx1mW20lkU+4rjGojTkQyUO7sTepuwZFuAgRxv25kO3o7oj4UeCXU
kD/saFMMmoIXecnE2QHO3EU9++0V8rUpk3Vhos16koTKz4YI/slu46N4BxNeQaD2
6OmIzO12huEvZbViReaSEkKSv8ucdKPDjng1M9gi6mHcQD90N/Rip5NFKvuuVbcP
TSOUt7BqHjCwXjfHUaHAnS0+d0Jdmsh4sqJAlCtEHBmaGlKz5qhqcAoyIWAkNJCc
soYAJNXRFjOKslJ0vjjbbCQ3hIOcec0XcgSZc7VKw2Onjg8XjD4XvSCkU66KAWyU
I7y0nWU4pCnLWRxOWQ6rzVBe/8fupRvx44Tkbb8Bdk22KQ+bG58Jt+wotoP4QWFu
ExSfWHEA9Poo19bxM40avdGH8k5roTGrornxZq3N9O3B+bdGGFkjapKQAzCh6e1H
r2t9ZVg2QANNc7osPazx4SMnYwk58hzzzpphk2jlYitlbIJu+Mn+bflIWNtlO+IF
AtKvp+CHQxmptnYDrdoF3amQK4hLtLv8VBmVGYIQuyYyum/bz/ciIZ1GWom+sPsR
I3ZzSiHVC8eY00NmGP9K3QbROh9MQPi3Z2WMorf6HgYjANGXnwqWXVFck0oySqez
UK74yqhvg9nOVZcYFbQ31HaV3mSQ5277HIBH9CXT+Vrmr5XI7G4u2qoDA0VTVDrL
g2yqG/NRKs3P8Q9oXn2TK8camNSa/rLMS88D8BFcn8PLk0nDXl+rf/jd4gHHi5z7
bzG43ymMEz5OgO/x5aCCls/TlCqAu0jAoEy7W9xJg4hc4K4WoXhIeN6vKanQ3iLA
4EFY9zoCooyiilWRPAqv1TGAMfL3gxOgYsgEh7EiJ3uy5WWC+xaWhyDCQuCKBhcH
sTgv4e+vwFX9Tj9NaZpjmltFsbxpz53eJbmQrToYYjBItaViUe60kJJnKrjHW7k+
ViWj7Z0Ptk1DIeBazp/jaEtMz4v3p/T5Rjh4mNA+oK37M2CS14qfW64Unr3RLpk9
k98TF4YDq5YZnfuQ14+yiUl3y8eve5pid9ksb9RAQ1TKJmmnHReZEOBMfAZASsg5
mSdDS9qKpKqb1RKdcucLJ68r44+ZBbg8otkttioh6D4y/6YQisBBS3BjC7gG7Px+
x57Awg1zGF1LRgNwCUKV1uren3rA1TiFNFxYGuttQmeLfsaZcH8sNPc80yd/jK8O
Sq2rl++fI5C67Mqiz+X45z8ycoWZO3kIc1NKPB8Z++Bc8BZ32Ma4y039KgClZRUp
rHhwjXhF5kx6+4pA2Yj5H34pPjL1SFE0IyIQuHv1pRzkAInXC7yXyIRq3VjN46N5
bZgH167YFuhpP/Yy8X72lU41n6XGtS27WPrWdmuBVxXMHMfkhTSWgBOjnWZk2kuV
7P8N20xQxkGteX1ggBqSdA82lVYdzTrBanFXk6vG7nk4TQhZiU8A+v6mYv6sEQAB
MCfQ8DDlcv03fFQTWq7sdZS2toQg8zjYy2lJepufHiGhSCiRSUGWyHJjN+Xgwm3K
n91WsDFHOVE9QKH+rpuSBEO+oqBAPFLzp3r4b0KGHV+MPTxxJKe+mAmG5Pe2GJMF
0MViZHlAsSV1lSo7pwrH27MlGzFAFMXGt0U5nPos/GM9wHzyHRo5wTrJu8d3neXh
pqGqnh/Ecn6GYRTyZhb8px+k7Q1S+tJJXZ2Mqv0EvVPQCh+ludpw4+YxOCh77rEm
drP04L+4cEWLobLIt//mGT2DAh1H6YhU07lUngPMOqsGncIfieMCrzfCRr/JYqnf
7nbQs9T41mltlSBuzOwUWUwTYovuYXWdygf+e/YwFfYODQu9CL0j5C/819uX+U4Y
CPIc12afrRgIqtKwY/yh7iyvT2S+CsPd+osKitcYvFZ1lXgNmQP4+cx7hOMWmYrB
j/fpBd290c3Ggh1x0p9XytU9Zm/YgnxF+NQdxxYgMMlaUSh3dSlo3DcXOGy5o+3K
aALNUkKVf4xrQjCdVeOB67Q+b9MmF7VXQjlB2vZtoJyGUSU/aF593CNzdeFtn3nm
a5/6p+GR8+XVBkprkQwDzYyQw0yLClbCeMVwIU0HBOX6ZJVk9jmu38K7QjK+k89W
Z0TzkJ4A+0Uhx1aSBHgu3Sf0GwinSKCHr59cR1YhZ3Ic0yNYpbJNEpQOXHE176Dg
TzAg582ledZA8ABth6x0/8KmP1ZblWgE9CN7PLF13S51ZoO7LWUqUwNczK6R3/2V
XZDpqQrqPhbz10fOczc/mEC3a0gJHMVv1UY2N14IMIrDmWWqfDfWHi5+fSs+gFXI
pSlXk1H7bmKxl3OGA7wSzr+s6+DVI0NyK09M+6UYS2kn2HeoJyBrcf3UIW8gsnQz
Wf+cs/nk7o02is+QRlqAum9OfiEGBCssDOEOLM5wCyH77UQ+2f3mltMjrhRz86Gl
gweZNo43nNF1A8afE0QiRoqsP1kXSpnGPkO5ydHrgsMjy/kPqjoe/3OQDcnf1QX9
fBgrvrF+V7pTstJeVecr/1lvIG8IpCnlnaP+RS6/jS00B/+1cSiIgL6CohFQmpKQ
/jvOyfKhl37ljfNoXlmAC1oxAj3F5NqVx4FRvsao23HXKwuhudaYic4kWM94wwCR
1/KHb9At8O8k2mxTgm4kNJ+FbwEPyvPJReeCXjdBWOVbW/4kUPIUojGHJWOyM2Si
qnRpRlqd5WDUU+dX+1SzAdneQGfCcE7OYpBRuq+a7Zetfo6HGAfzlxqepyEYa1/u
b1xhjgi/qXjchdxmjDpLEfPVxmUaPGagcvBO24Mt8b+przLa9EZWEalG+Dhk6bTK
iXzk1onyjTp/jzfvwmZw3igwnlek4F1rUk/mnu73/Vk=
`pragma protect end_protected
