// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nlUPmX2gk52A1LDVn3iNHGqUL7wV5Q43+4R3bbuRJoisIqtRBqN7I6NZ05EfTNyv
nm8XWqc1TyIx8MXBBNaZDtvKPBqdTR5//Yw3xKEQRhmUSN+GOYnIDxaj/PpqSmoN
rL1plg1aAIf+C3tkX4ocPhP3pjywInN3L2sLIWbDkYA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4032)
YXp3tStoAIC5PxM2qrWRG1e/2APToNedaaQWFkJ98Cv/fDQ1798wEi8xXNIaw3u8
uKUyzUoVD8x9/CDJIDyFxJ7SOv3mCbQ1d3hf5Ce9tOpu2bkv4ex1jXCjVxstfhu4
P8dqyPj4RQxMOy1PSHufqe+l5fDkeAQESj44Ryx9KwZU2q57or330JyNVF2Nrvbj
N8AJ8s9nzRCUG43McmQ3dYGxi2DkSXUy367W/iS9DCHqdylJNJ072xQ+AR2jfXIt
B2WH+0/CrYWXDqHX4X+q0U8sGp3va6llqJWDxEnHL474vVU5BqJpSmd9DS6JnAj0
DS3z8aNuc+EkiC9R2DF7DfrSFPc5TFrBZWpyX9XavvElH5HC4LKrPLZU1HmcOPqY
90iVaUi0ctHxaFxtS7MSKaCfsoyBKrQ28r7FHLO0VIu2hK87o1LjMdxrsE2QQ493
V903HYidN0Lb9E7jDUKDeK3XXSOOtHJlR2LQCa2z3UyDLRp2fT4QMmePtBs6KAE5
bWbWbjYlAw52x46ZkokGL7Wk+3y/nC6zOotd+rtrqN0syX7f6OGKOfLrcauYSfzK
YRhEE1SQTNyFKra7TyqAAVe3L1qeFOTQ+OYx0ilh8di/a0nWWn1opkl9wlI8f5Vk
iOeOQqlqesCjWdgVW/iOayh9wp8UhTpBuxbMh6O+NELiUf+13AZsze+IhCO2yZLG
0yO2GuGrcVeTp5xJvn4Wn+ZLRTYTzBIsSYLW4B1++i2WCcZ4O/CN8vznAQSdkGXN
l1BMptWOKEWyonQvhW3gfRdPavTLYzujYy8FGaGwDPehn1SWy9ArcuquSZJFhEll
4CuzcqTi1wJtjmZDgAz49pAP/9WNi/v/2erm12q/AluqHqUUkQllNn2AJuIlYmz1
X/OD2VnW8ojD7IujUGBiZNSHeEY5sjyMCCnIpCINEWrgZQXqSyVbpVYYMmfGI7Kv
N41iRrTp3/JsprNW+c1aMD8XuSXQMM319PkkKhFg70soMbZFeSHk5+82d4Djwmm3
TYr9CqjaU/kLknwusuURpkTNDbYQr+nBYJt/jkMv298HJrrUgDfiJ0+zU9KHc708
hvBsOILJpsfE0FmUQjnf4yAe7snIuFj1Wi1wVDyND30APLC0ovVZrtMoAkNOJSHb
Fw3+NWkJBQurkE8b4OfC7iIkznn2gSE0o5fiB5ph3zOC6R98ODkTO7vyhBjHtG50
iU+bm7SBdA7QIQcGa2bg0O4xIZQ4pBm3zbWBGIXZworyBywn2mgc5lMVB58WOiQw
RpOarOUJtKNDNLDs/nQubPioyq2CjHM1i/7S3rh5+OYBfGd2p4Dn2vMlE/jIPW9L
YDC7yRfOWd/7+i1LKx5B6IMT39z3vw4RcvfW9DG3nZf0GxgNAZ1SeTDWBXg1yXK4
/6MFItUQdseQw5e2ulV+b3MvjycGV+Yg9LF6XF8Scju2JRtehznz2RmSaWEuILek
EwVaIExu9CnLJWNib3XdNSpAO0WixkwjeJv1ZLkwlbI44eWTw3HMTrgurr1ICkp0
cyBp3AA7xFXeZBrMBr9aQGMi9wwhkPUYxpDtYs4LalExOMg9CDIOX2j8bVCreQZO
pX3nGEXI6UJtNN18vdISiMYAnkpSaXi8hZC+B44wOIvwtZGDDwREjTFNyBFMqnRj
EScalhklz9VB/fCXGLncXyZLVuxPgW6fFd4EdFdv6iEFvQ3JTxMNlQv+uKXYyBjO
igZr1NZ/jwJGuEvWq9z8yC6jjzp48UKl10YiLnn+ANuk8vTw+72/hd+N3llkW99y
sY26p0UZi60MqRTKXz3kGWhSIqZMfunAj3em+kHB7xHgv5LBuRwYUvGpdaioHmJa
+vKwqqEpi9QHXgRoKQOEH7ittqdyq2JjYaOg7zJTy+aV9TGWacde3yCQSpb1OV0o
6mUv0C5S3jHMOlaChl+6V26lRM7fYsCuZedBxVNhvSTVg+Rxx3reADOhPw6svBE0
HlgkxTO8rqLOdDAXvT3+E4T7yIRsCzWT3TwddPu3nZ2+IPz/BjLFrqAQ46h7IiKy
ODP1Zkif1z21QKO2yXdxIuAOl8HsRblZmfxMysLKIY/ecFISxObr+XJLXV8XIUfn
LFnmECVLJp6hj37Ncraz9c3D1RNd9kDUWD9CuwJhG8zVFwisINNNO8/2VIUv/dv3
IomKeADRzfa9bYkqpKp40puAuNyTZpQSd8rPi8/wT41TxZySVjn1VpX0Ef52hKlI
o7v6MeBHA0y1aX91hG7KKGZfdBHwihmuDX/L0vlaZM6RPyYxuOLq6GouAWJ1zWOd
D1mj8gfhoM7XSzjgc6/cbkuwoyrbgk7+CkSKEiv2ohdE2p8aBPaLQkh/jJjKqJV2
DvWSAq8EA6Arx5W4p9Yhtqv/YwBHLWK9i9ubaCqAHixSU0iTlwtECPfJxcmXBsDr
iNAS8QVGfWrnJeEeLz5+oybd0g0yTgpKiZTWsBRBYez6LEbljSDprPhaekhPm+VG
MEDYiBcHaLJZ/6xug4kPxE2fzqzV50nKkuMSAbveJcoAxn7hGxYCRazXad/5PBAk
ifutmMCzFTMBbu557z7bOQndbMej9p9W2jMaPRhajzQADaAkvVPlITitjVIKRj8z
fDLItyCNcfol9fpeIgRukHIiF3hxs01vlU3xXe/KFVgtOOgsn00oivqun2A+f8bn
b/VByacNZGZcLMQW2TEIxbiyJ2b2wq7P0SowgyC3Wfl24YwvnctGiOmpTOFZbF4U
C1bJqHbsVNcGgU2wQJofcI9TqALL0guSQYLCfo7tcQ4CMbPa/5TdTk8+pmu3RRWL
vulDhPJPbOikgwKwFXUz7OOmTgmKizsS5d3sNsHxYOGeo3oOSH7cFNM/qVA8NLjX
w6F9oK4SZC8Q0i8fjHXq6cLPahykkjIPDaMD5vrP38EU5w/MpDkUgFGHBVr8vMa2
4N54acCuqahtX9ffUBXKl3NdrxlZ2CWdF3c1FdnZ5rynluymWSTdPVv3d0L0ciBM
VFDc/wHo31zTogALZxy1NBvMub5MADj98ODEeKe9cw1FCYwZ01AZupP7iJ7RGpAG
3zxmUHqzfM0a54TwYbDXrILIrsyW0ntT01elz/D5n97MAvjs7wWn0SEAChvQCHY9
ttV+5/CNOpfdiF9A1K68fPEJbd6udLt+bzGdQgl+16u00I3NWxjGlgLGlbMMYzK2
y0UImSoqpwbSLWdiiLnqJ4/UhdLnZqWrORWUIj9fLI2cReuKvGrjJTQ6MqgELv20
EAP1pDafuO+Egw+EnH4iniQ6S4r7z6qId3HohPYKnfLjy27QmWqnOwRnbC9Ng4qq
/kW8B4sdYjKKqf7dM47M3kGRZuNTNIC/Ek5j3WcWr5oQSdMro26aLNvXnEgDv8g3
SN0yg/Q2phUleqEN2KtrMdXrv5F3LUghY3E2P0FmtU6mP4xCgTNwZaVbiJJk9EhT
dlG/Ya4eAI7oiJ1KpqePwmF6Z+c/o1efYmAi5PDHxdc1iIPqrubqmoOnG7XAtm90
2OJTSh6XXR3V1gKgr/UATKGYgtKMsMqQf4PJgNW54H1qVsqPo50704Ixfxk2+tPN
iyjoIrM2pGeK3kbSO9yjkpdr+T2ikuRUp25lewuczyi4JPGAqEuleLxcngsKLBjH
+NL54MpwsHE16C3SxCVukr6wSh5ZO4gb0KiiWs7ydsXIAR9wz/NHmomhGVEPU2K8
fjuLEW5/+it/9AwvOkYFFgjMcO4cDfSHqny/jgbotx0jjFUomWEHR6492BIT2pyY
mGtrXHFWdtVgGT1NIKryLA+xwm6wr0YQ5gtKx2WwwMUnRinvh/dr4MkDav8B1ov4
mWz5C1cWTegPoOfgi+B9CwabU4CUmptLWjuBHe0DctUj+zPsQPxActpWN98J/ofc
8Lscop7ZpDeIFW4TxHeJJdbOiEYFmHjcV0OunXVJEa8/ifhmVZ4vbJuMdJ/hBG0J
HLGB/pFsmkbuoj94SiIyV6+H2KjoHjSvMlRloNlvMT1vObpGqwgDxVZBAlU5MsSC
lHsj+xNzFG18aIRu0srZKibRwv8ciS0ZRq0HiOMTJNIIrF7YGQal+EGBa8vMNayP
CqykTQtnYNjMzUizygjNot2ofE2rvQpNCNQ45BJsCZifp24M16orX4Wl/tSAICA3
gBl6g9BTUy1fWCeWBU/kPFDdpTzN/jQsD/nIzslug2ZPlxgo3XpNeJ4m+zbgqPJ0
Y08CmlKoXFbVGiC30z5vvKwfd8/ozeqtYOyNENQhLiQNKYUhTtluc4QfjcfiT0qf
VKvP9SuFAx2mvkp+vZ5SYZJjiH92puA9JI9JPYkNY+mvY70Gm1R82utLKGCVEDxL
BDjk3mxVk4sKNChW321M+OteBGf11LrODD2ljL8tPc+mzv5hoUh3igXQMw4ky3IK
kBnV/Luun0KyJETaSJOS8UJ4pg6LGhYJh2ngR9mwcZqkguG/7AGonA870k2rdmRL
huRbS9TJxQ5LG7CMpdNLGEfLQe1VHgcMyr88e9PUcw0dw3DnTWaL8XR94E6R0wyi
X2n1+9CyvKIacQASOmqg2xF01ExnaK/8QohK8RRAun8G30PQ55OAC1olxyr8BpA1
sTaLZ9/xBU9Y9FAROrozEram6yLAMmAy3GIm/u/akPh/fRXF2N7Q72AX9SmVunRA
8DWIn1qRoF4hQzCgLRS0SEHtl+nvKG0iavvqw1rY5YMp8MWrizbt9IommWhdxzxY
1bqQdoiog2j8nb4W1igVrNaC/NdI7TgvSAncvbj6ihs0pyPdDZY6DX6dVgkrqoEz
d+0fcfwr+V4a7h2QEJJ+Uv134eqDCIZQgxXP7esuMHQJMKaxsXkMibOE0vng3mmL
6UjG5xR3PZiZMXdCoTbrFIruqOnYuYJuKFLvnjTfjpVmPgmc4+Fw2NZfCctGDaIU
Q8wYXonC5+yT0DoXSodgqqfctoQWA6Y7pdM5PAREAlQVFpnidNP68kEMEU+A4iQc
FHXQ0XMgJLBvmxwzspXrcCZlWYlRFg8kXWs8TcWplcx+w3+9NT57nrkV4+JPektQ
djI+NEyTMaIfOmpggsdhqpgrKqFSr1y5NzFxjXP4TjKWpH4Crj7G1d/N8oDt88iF
wu6outZg6U2OiAmkqyJe7VxTh8rxepmStuiMx4drRKmJa1pUg0Mhzb+7Mg1LJtMV
+SzKjJT9Kv5TDt+LWQvxf7Phfg8FIbmRokAuuyWXmSqdRyFydh+yZMG+B9lJaFvV
8uisuREdHuzWAjwcLfqRvJFLbpzKTVPKlZq4TUxpqypKZ72Qo8ldMAKPQxbOhG0D
vKeQ91VNqgOdFFKyucHFcbRhFY2cihytkcYru7CynULZYPRhs6k4Zi0rM6QsXo+P
`pragma protect end_protected
