// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XCKcw3Nt42qKQKNJuto6y6yX9KQpAyq0VDaFkHPhrIkaqDuDGsd67rFI3j8e0ICi
YFZHhiCwE0hE4bO2sz9Kk72YEfuxBVVvMRRg/YSbOzHrv+UBzovh1BW6od59c2nZ
xq7ooxdMs6iyuM1ln/5DONeNU9ssh//23uzPtJ/C3Po=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18736)
aTYB4qal0801pagf9Vz6wKD4ipiZgkEYwtWnWrjpr3SN3bQ/LUbAfEXOZBUMjyYF
yu2Qke2TGWpTLm9FKpDxIYHi8ULad5iXFYVC6C3XuAzA+Gy4jgk2AnwiQpJR7E5p
uv8r+vQy0nirggGCkCH96hhPmPx+Z7/F10OnCYNVnUWPWjZWV47CHhwKrBtpVge8
vk/dUfU7CoKD9f3lGzn3cKXY9T/UXjdfbfPxXD3Bjn15h3CicLoE1StRwjxFkS2L
Y0jgoQxUB6f0Sn2A+PZTfbVtn6TCvRnVINZgvPzqaGxvr2gF/CpyoalyrbG3E9XL
t5gHvWvgGVNRxEyjLFlBut2e760YmlM4S2gyi4tZQQ7Hlec5w9Lq06ZttEgBQ0Xm
7PwgMx8MjJTDl4POm5nGIqHRsBGWZL7aIkqXm3gI+2n46CUdrhG5E304yAVBuGQp
sAxQOvIExJEsTDyPt81GLUlCNTT/bE0bh0RneSv7q1YBwjx/cnFlD8vJqfXHte25
AHXlMI1XSxWcOp4gYbh4VwwEXI36fEaYnJbLeez83Wovq5xvECie8bMaCSoJwayn
mol0I/bu9JMgbgxNFtqN06OOIQY/Su8k5z4ySrWl0yzu07hk8EpY7TPECeosox72
Qx9PwSLGN0u6z8MJWN7yD3EfSK0607xU4ZXQEmt0G4m7vFZbUO+DDxepXJfbFzmf
yC5VnnrOqIzg9SM+ffNh9q7GtiiUBETxhpCc1cFrrjHWAHRD+LeThCpnDHV+R6jb
57U+uwGQkBXGu0jpf7/XjNbdX5Ohds3I6z5mD3xRA63YQWdqWjd9QhjrQjvdIL3E
tOjJCQTUbbnEQlz1EOuD+2qo9PRPkNkDdHDt76HJIJxJjLVW9kLjMw6rrV6nm/rb
THuNMCBnig6z/3b8EkdpKwNTI19rjA3rsm1UrQa2K1c7yuKGrC48IlXCpdS5OHZo
zlYLVcBqJ6Ui5DGcfVk/XspXf2zK7KZ0wKIOOopxG0pIR3nhjtGyyE6RChpQkTJd
e14JS42cJ44/QjREwMYnXzzlDTV2L9pvqUWvqI1gESSApPednWgN4QTbhbyHnQ1Z
lsMhSLDnK5a4ceQxM+Aj5+PMY2nTYyDv4VzwMO0I7lQXkiMjRGCy0MrSRcH5qUFz
jpzwvwOOqfzs1y0JqTwSp6lkwq8eiee4yRBWkaRM/Lr3MutFzJTUEQK9DgFyjIxh
+hPJaMbfATgE/k5/S1TXlTjHDL5Jbh050MjHujpbprGNkRJIHfmlVWIM9IrPmJjn
o7liIFM2U3t8IMEw20aHwfwDmQyev4zG+NSVHgiyv0SrwOQhFkaYcXhLXW405Nep
I/Y9EAADzap5s28bOfrtw+/LPI+eJ0dIIFZtIfc2PLBlDeT1jkYasv0bTl4tEBHL
no8kliWgjce1v05hj/d/QFqHtLhXbrsOJ/lfxTIS1ZmNHPb7zZShFPr4ViMMAFW4
vkiqp5LFLBCJdhlacVeVudnt07iEKgrB496bnPzj6dzTDwHuG9e3rkIOzA7R4tt9
n+DbIlhW0QJdL81/lkP8s+ZO58O8/KolnoHXSbwuciohyJXHgSTA14FW9Ru8H7Cb
pudx2w/qdrmW5kQkelmgEsoBd0SPOqyhKBwd2O9jY8AkuqNhCsAIXYekJf1WcKMn
MLiRQ7TEtdjYJD6Tl4PytsZU+pAHdRJC3AJ+mMYiowk5psiWIYDPwakkDj2d/OA8
/DD+sKCre86KsxLgLDLfqDBGrwVmIQdm0i6f4IdyaLmyIBA/FZ7dvbjh5qmxkCrx
Y+dGJP5j22DbGw5Eb9Ngl8mWxdsnZknwL83s9pvLnruUMfXOpYiszg9j8aUUonOp
lAFpfDrJr5DUwmFqXnHojExv5z21GYobxADdSvnIDBi5PyQkUxBPqzLGgMlkUzMD
xkHEoK4jvf5KaLKNvtzK2hVV8WPX1TZRxsFev5SHHnUyqByAb0Hz3jKagME51KsA
+rNE+l/vS5aBPCXDLxE+fRafOHv1XCkLAgVSTqUUx3WU0baEFWLgh7IQEo0+E4aY
m1dO4uZbDwJtQDsw1e28F8t4Lt0ZIiEuTMRU9dn17FC1Hy01duj8WIdLKySOZTLe
sa0G0ml2jeFPbP/jr0MHqMJEGDh9RKzpwP7M4qs54cds0wbpvSdM5ads0xDtWA86
nEHtwJqKaR8+Qj1XBlwsFUT4WG4MOzwJvQDSxdGRR/kefbqBLyvtPUe5bwRRBZcc
XElBq5BxJun5ry63VovItYjXKwJdax9B9Gb7iKuiwMSLYdiE+AqyxZRcZy20n8Yv
f/xOw72GD1BhuwZvN/qxxbHDncTtXcATAgzLZLDfilcum115xvFOmM/ERY9EQy91
lCErA0q7mc/9y/y3jNIYlsCXEqJOL1LbZspb6Av3FXh1vujIBk4SVJDAC7Fd7rFF
PvOovxefXswE4i8FgPo6nsPB33AqhZuGSe8ly39qkRFFSq8EIgY/RVLTzMry43pn
5zRAwLitPMBlBoif7zP2DS9HqHkhTfBubH8Dchrt4h4HwI2XzMQ3BXwM4cLKvx7f
DGUTXQ+RhmrGJXlfzAj4GLA+D3d8AALznV/+McCtiVozZodT9QWKBlJvF6hEx5G/
LXyrQORl6Y2N9orABY3/kdK7HWNP82w+N5PSfF/mnbp/jCnk3qaNxdYHagcE97pm
a3BmCN2eP5ZR5OUcxu3iOjNVx3X50oKBr+zdpZ0CUgeADqFfOsRkjYyZzvwwCCZm
JTKqKZ1kJ+jQ/ijcCQVcwNGE7IiVhA8RRLeb5Ii2tnd/OJkG5dsXi97ICU0InAyP
Ihp0bdLieAGAmHDSXSRpYQk6MEdcv3JGGbxdknB0VtDXKVyouggh77yU5wFdjiYL
hMgJwqSBz4V+mYEuQgdFrU2+VrS+FA06Hs4bEe7+cAD76wHrg4ZyXEvQLp9drb8c
61d9HCExq4iMxW8/3Fzr0FxgsJq+yOWQAK0eTgzgipuFkB+LpZMCs6p8RvT+RZsq
CsnaKAAtalVQojMxSlgObVhbrFngcbE8pYJFB4YQWIcBZvX6+hOE7E04gqh5I7eR
ScyaadeZZDhhamo/ILIuWJ86mhCS0f9uH7SI8o4OsWaNmSCxfCHc+p8+b/wR7q9W
Ny24EnYgR1ULtQGDZV2OVkeNd9eERZDsEwztvNPSbBsjXmh3OUbbO0lcBcPkn72q
77GzXE4fCvUkPIJjxpi7aBdDmiLtMTPK80IuENTGwGMLBEYqK8o1N5/5HZojK49Z
hLam5ZF6/GHU0Pov04KwRuCeQCASlDBKNQBRFh+tYhOZhcjLwEl/PZPWQvuWgIlI
tncl8SLe1VLNjgK9ABD65JwX95qzE+s4IrcyItT8FamyzRwQU7y7pgjv3tg1yAYD
3WADk9RuhSVibUU3BWwLmThNBFKj1thTssgwAO2Hgh0xP/PPfddANui18+kB+08J
Lwyd7Ldpa+BIwio/LrdziJw0cHTsVDhkf4zvEipb4yCjLt9t/oXUCouJY1S7n/E4
+6p02u4tmEKR9ygBH/+RmIdnz4/w4g3gto+OGONiyUM9PuWEPXWP8mcmUqBnE76u
X9tmhzlPSSClOrA+fOBLZ7ncDGw97p8gKMrAtGy70NXABaanbec0xLxqqIx9Ddxp
LDM46tZA0aTIz++0Q7AYTMjiDYJC3n15wBnJX82rZMo9+oew0jZ248V9RhTU9fAQ
N1xd7urTSOXE4M1NMWrJSPz6ROkMWiF48BmbGePEcodLbod/FDKbL1m0rewyCJ4S
OlVWIyQZN6vmxtYUBnyfZCQvu1SjvnGM3hHoIbrvXVI7u5I4VQpNSlik3ntl85pl
ijhuyGHw984e0r4k+q+cXs9oBjgFS1ZpSFhz3ic/X9TO4Wf/l3XIvPzYVjiMB+Fn
lW0f/MFMzOyAjP/v344GZkENG3RSlK1J0aepndjj8q6tplD4J6LZ6tFIf4MKqnnd
54rQmySUHFyvqr6QYy80VyOvV4v9+J4WIhXTArIJBZ82pr3d+zIRZDlT93rgb9cP
+Ue2Mh+0DIXsyT3Ui8e+NRnXnEy6eSAWt/SdNmURmD7rhJU4eykV/acXINRGiq01
/nwxySYlbz1fX22ERExgrw4Q2FUruIHwB0Ue2ZBjjpAmzCU/q83t7jwgkZDfAyk6
/coxcYqkilPGIhnTyKDUAB5GLXEo+XJX8ikeGXm7M2u0cOqAg3BPK+vH1FtPCaw+
AbJQc41BdijrcmF65NFv7md5yw4GWfhHPv5/+rkqrncDfuHMdLfREHdmyGG6A869
nzcnvyMgPnPBqe3KCRsZoLH+7XBVE59qBRrHwaZCNTph+Dz4m1gktpl9iM99Ua4u
jucMQJTrwN8H6T5Ti/tPiGthPYnfoZ3f4I0coHjwpbtmKk7AcVzy0ilcRtsE54SS
aWfLPLY0EXFC311RpKshJ6Q8FQ7aGeI3zDvdNSQNBlg2WEeBsHZ7jTEL+E+T6I+j
np3pmhVO2A9QogEgFUEderR6CnAvs/nsVzlgHJOeG3w4gF8wBJ82aM/Oq/HIUXrp
URLufRsnrd1qu19UXw+ihGnoC12iv1KzAqBEVHxI3++z33CnkrMhCxpD3IMCQ+G5
5mS9A5zq3DV0ANmYGydmDLf+rQ8FkYgLWHa8CfiYaxSWsLz9IBzy0rOVWGgslBL9
/R/31j5eVxAXV9Jk72zDyYrZGMU9vfj1VxuYOuuf5nKsnskhUvQfm3L0i7pFvxUS
nlQRkNRnxXAtXA0xBzq/0hdOOO9KJAL1B25tIBVAXoIWo+APuLf3wZg3Tv7TTGMm
Z923YIfXn2exKmhZ+JwDMPmgGsfTZ9lodR8k9GErWxZByXgVKUnFRp2Nb5jcVVE7
Bd0dAntiJAZ52jw5ta+znyICX/SlkokEsQ7mDLMnrz3CeINGb1jDNYk8DKm5p23j
qF2ucx2fzJ4HKsmDruv6REEsUZvXV+/nlTfvNKc9dGZ/IXV8baEW4Gftq8TzcOFs
aAwatts7ApauoQCww4Zga0wmpyIdLA3SVs+bc0iI7IXK78U1nI4jaR3vI8I/fpF6
d120VOCSsfhn2eOIXZaicGpuFta+iFLT78zScw9MiIOelUcm3q+1ejj3L/dMdf/A
NvIu+NVRgpd1u0P+iaK/y5vI2PfgrUg1XQmJ4c1/Dk0ncdAjCLr+ddTDEAFCrx7e
KGiUMQ+QV6g3+5pa7gP8ssjweEf8922qU5Zpl4t2h5N2l4rh9AgMhNm0KE85Imfk
KSFc+I3+/O+CZTw3W66+OH1adVixuA75K362Ec4dbGjWf6ToFGtzaKhgX1G/I/0p
WsSiErovwMKMjb/Zdfl6/ke79OqZ5AO46uLR2TI2ihKi15+ACnJUew7OO5q1gWAZ
+pZwpuVs0sxhbHKogvF/xarBBBCVlAaGsDSWaunYJSB0gp+lmWUeGpD0kmPj0z9W
677Y0Ly12VkNpWYx+KVKlUDeDrE1EdvUodsHRSozyq6ONsI1oZd5gHMNy7a2HpYr
fLPo/PGxKD5RnISpgWY4GpCeid/g4L9xoGFITK9u4pqgyA9iL8SyILVirdk/at8C
A/XoLwitzb9gD1Npm9cYP3ZDMqGXLOVbrlIQdKy9KmYulyphcedrru0M+l4N8DeS
DcRONHzK0BOmb6zY3+VFduPexU3g97vAFTN+B9OOIIRUrXxRbQGybWK1HluDI99z
ubRrpZCUpVPbNSy1dO+Hd1ZH6xmvuJ+lCmcMN3X7gpch/e+r+MYQK3Gi1as6WKnb
DNM9T6uovmdH+6JU/NLmuKbdhGolfYaucIwAJvGc1jXUSBWOVrfXwoueAJk3U3EQ
oJNk8X3Bp25agpGeBtznrqU2ScgQAErTtWyHTHTXenFbPOMjmyXM1sVLXy9nP9sE
e1wLDoY4saf5joqW0xUJlh2gnnEarLzdTmcOOIs8sIRMBVS6IH4bhr5IMnN7y6BD
J8mnC2nQP8ZmiItCp9GEuZIq2c4yuD/2af//Ly7l/PnPC1/miYK73k5NiYhedn+d
wipFJFB1s6tmVUyNPz7cU+v3+123epID2PXPaUpPsO+bii8YEIj6uB41wq59U3sX
OCNvJKdUX1hs4BfvIqQvGAmje2onK3EJmAArxheqiPyHSS7TF1SUB0/wQS4NMz5H
DkcWjNY/vozLEwu6yc1RDCZlq36vNi3EYZHV0nDofO2+NoH+HDahMvXB3gBZYr/g
wZCjSiz2FZPwEVm9QW5keW0RwJsaw2cQnOoSnl/2SOdkM65Iy1N0q5MzI/kQpWSk
ymW2WndQSU1mqnZ4n6j7ZgjBdeG39ffIqaRTLy17iyFPs77d+ej8cn25Njx+g5Np
RibQYyILam0R66+4ZJ5f5/cYa478c6OBodt23YoyyUcHt3Byvp9Fi/ehYUvlJDHq
+FCYPPgmzWizJ25/sDHwB4sJ5OplGZAByvQXY1Yt3moEzljGwvaJ/B8ZeGsiM2KF
u6K12eovEvqwDskS+Q611El/A+nh6UsjcYIqU47fj6Ahh2vfLBjPJrJfck5RRbYX
9YLjA1RK9i0wW+RQwbnLcmh9s9y27OOXPR6ZRbYeW0UZd5RPtV0ArpsB79sOeJ/e
NwAjBT4jyXqHIUqikLoTtwN1sWXQNFOF33fX7DFJ0dwnOuTbVP7EBw8qBN3ia5SD
YDWzt79iHuXbAkN584RFPXltnhhT4N4A8lMyNq9IU9W8Ol9oqwZ8xN64L6V7h3SK
g7l/O88qlOEhvRz8t+587qLsI8G6uSeC463Tsm8AhaxgRrz2RhH1orgUgAvo27di
jpA0B43SaBlckesL7gHL962HonSfDobqY77mYnlex8Di6RCnMY8tEtOK25Ya6p1n
nuZmqKUTmVbGIjVpjgKf7EcJi2At5r1Wgn89Xgh+jn9sxfrsD2JTdNn1ChPRwGsR
wRBNuaKtuq+2bW+18TQt+zz2X1L3oZNMWxXAtkwetzZJyrsG5lzzR1Y+rCfu43c7
zl1Nu0FkhMjgn2nnBmWj3QcYN9NfYghLhphlO8g/GCLx86R4t3+7l5taLgJwMTYT
DV9G/avzGYHLOXn3/StSkJvqkFq9D7JA/swO/bx6U/k2odE5a8/e7x+y+d6R6tsj
wQfV10J7tfvUKNu2hSaURkTbF1AL9fOq7kRSd4MMCpd80W3CYR0OuG12Egeb5t8k
kbdkXB+jxWrwBCHRA6r3UXm+AMhigvBMMKqh0pbDQ692Vq+uJ8yON+nvn0KIE3Z8
SOQEUQ69J/oNW1nnipIEi8aU13igCB4V6n8PlH/yMTAUSwaGP0ikYzWxINHK+u98
oYg6gmhLBoUPNhKA9J3LRbJ+Q0b4ZzJGD6UcZ6yCOkDT17kceQvQWgiRRjk/53WW
q+alR/KcBMXEJudERuUzqZXMdwnE2NPJjtH98s1tjNQN1OJumbTmvt0jb1yFxHsG
bFLPiEBXvZp8r5MIBYTt18GJlJsML0d5ljA5X99yUfZHDSwIF8B9dwRzs2Ksh2Z1
d5GJV96GOV2uwzbb/Lar9zTgFISUHGzETXp4CUuJcijJs3igzQ8gPfnHMdeGy+Sz
lcSVPPFP0d48UaN6d78FJfTDuLZou7RYythEplrrle9m/aq+XQoHvumlIFNXWJYL
Ke8C/9YrVzjK+1k5c3itOa5NoxOgG6Ebup3J7ElpQoGIohiJcjKIG4COC/FE5lax
ZP1/3pifDln+AWeeUuqnbHJz9k2lLEiP/jd2Fnxa8SBcRekjrRLQztY4PAhSlwBE
AH641DtLKw8NA3KENHb9ILJG4bxtNRAJPUrk0GND/5AjWIyz3lAyAGbUJob+6QOb
i/tKeYPKmAI2IiCCCiI0NS0xwG6oipfBSpwAld+oE06IhGfs/PEV6ybMAKlysLn5
p0XFaIfdHi9CSxD5JyOt1n8imKqVWKDlNhOZNx4TppcGfpAIKysSXACYZSLS7VU2
raYd6SmoeDuZCOJbsGCdQai80xjHvaSWegS8CdCZGjznj3S+wvK03STlL6VQOH2+
qjZgRKx80WurK0/M75j9BMyDaXVL5xSA8GlORgAolzwqdU17l8T+xjnAkkYVZFP8
3jSxVqgyQubbN6+4oZVlpWXVICU7V+JEoLTflWszKwy+XKKg/UmLg4VhqfnN2F96
iTX7BWzLpM51+ImU88/da0mRTFXmnYGfMIMbfvE7SmZ0N82w3VKuyy/c+b9QLnwQ
J65+7IlBNXj99bBpSKOkfk7sZJ4jNW1WmBH1NKSDHYbuaZA5SVb+QzftVixFUYUw
thZLjpHfujTUdBekhP/MuoZcOixGucTN5rwdkvNuOn4b3l/13vKTqJtRrEyPVvNO
cBguYCI1LvPSyKHhDppciBf4xotc0uRZKA5d+3Q8zmzy+7CoJOKUmOO86jSEeN6Z
oq2P8HSU88Yj3nUVxTLsrucAYoxykHQa4v/B/u04Kq9osNjuULzE10rpO+swj5JC
tKWQgC8ja9E3x4DrCbh95W4Aip5IguQkp/iDORUIiKM4ifvRiE2L3hVX6V+QsZJg
JP7pc7kWQ7/wwdggjjDeb9TwtBCMTrtsJEJk5JDkkWw5vsqG7GX5lg/Qf8irg7xY
h2LrovulB4GXlQSlhHkx/b9kLrN5MGPPJpARVybFX4TIvR++xTqPhacF74901moS
yGkeVAEXsM+JUJMqKYmM2uivHP9QpgEho+1n7wD56oKEHqscItQYOw5zWEj9gstg
RIuHE6C8OpU8sfkpT//Y6KBdZ7XVFEnVqMevzm6vIEZ+lAk29bGLvUCuN0vW4hN0
ZMDS2U6M7/7ky/TXmT18y6fPJLu3JyB6qMKyWE8PwVQcnBL+IQxttGqtEJV6CZPL
negSl8ZzDJAFSxLA/w6CpUNDAANoDgtuZXMIZF8XkSv5/HjTE+R41ggkudv305Mo
lO0k03UiSzr/pCSfwTGTtXUGbOBFjUd2iVaItUgGqghT/cxnrTeD8NAyhWcz1Og1
a35yUZmtCdmgCg6nFHnFJtLTp3E2NZsD6DvqM6dYGvaGCuOGsSWMlsiRQKx/17o4
eF2Qvg31vv1i65Ge5GQ5pWyhQ55DU4AlaB9kpyGuc7WbFxoC5/VsvSjTWkyCShSX
7eB6bM551XiOWkxjDibcSanehS+MhqtxUTJUlgEZxidX1sv0Ua1aqnl5kOILE6li
BzeCLlOVdAhRE/D2mAOA/wOWGJ8IGf/j8At06nFe9oVfDULy8Jlk2YxGnfg2ObLR
PAacQltKZ5wrNilFY72VjLFrGm/O9Mh8WZA7agARmeR7oJORfBMSwfr2pVO9zmBU
4FEljdndTqwNeFqzK8HPSixIskkqXLUbV+AzUFaTk6f/CRFaChwLB7ybkjwzoaBg
UqMh0MOKJDTFAE1iOhTCz4SIeZB6+yUT/iB0EDrfSdaCQvAEdFgcuA6LeGYB1LED
BOE1ZST3QdzLu1ixoRNy0GbY9/K+ewCJcgibEtx2ybQyA9Hf5KmAyuvrEvasZYxp
kg37Lfjtt+ouaTIb1GTUVq3hlwpyY6CPO32icqCpKWmPhF4WRZ+43hAEb0jMrChX
7Z7FhM0djrtn2Z5SxXJp0LI/oLClQz8N7HzrXB5A/WTEUBUPulvV+moCgh6dWglU
hp8fEIMee98JN7Z29IkVumZTjy9FuSJvAYAzcbc4pBeADSdM/U733/E40HVnYra9
mJUvMlNb/hJ3rwX0m62G7zO9QkLQzq8GTisXIFgXfehnhKJgHYDNGHwd/8XjTVHh
8uxV57N1eqMgyyVwLU7IOvYOq7W/XHC9rXjBZ4mCBgIv71ZjtQFbN7ylNGV5pSfT
JVRJfVrA8FXo4WRGX5hKd0zcAJas+jRKkF0IoEdaOaa70KjuN2GLuMrUp4k+iXOJ
yVbVM3Pe8hC/XwQmp6A0ozer91OHtqQGd8tqyQtbVQ0dBy8t0/HAqjKWOP2mcaIl
wu/nBviZbmGU1u+kcIopEwFRnUaudPPtZmwoebUAKTNqD25+ybuVk675LJQvuTZb
c18RlJwwxSBJoVKc+JpR7SB7mIV1dyCE+VnNgTzSXCecG+laskcDddoWqrlF+gr0
ErarhKUaoFrBobz1dPcI/G7PpOy1VubYMJw+A2knS9w/uzbpDFeaOSEse+VsJfwW
FS5dddtS0MR4QXx6wHBrEbC2Q+eIG+OZ7wNlUMT++qjp208nIaGETQJ1+UvXxsgN
4xpf85AhLresMeKrG6kvVt4vGjhMcz3VlAGxHi+0Q3THh7c1IvC3sfiw0ivSQvU1
S5bUu/mlLLRmkhF/HifASTOdXGfy9j7nYXztMB+WQOmeqnvuYLGL0u5ahvDugr7e
7yX2qFQ9zPBL0lKMcvUXAX7cmLlbDQdDj/0r+XhaxyoCflDACX3JbjyvX0baIZ8q
fyF8qhzERBY4b0VOIE800IEOOCClGpko9f/Qqv8MGv2hsRITgXq7KEiCrhhot/0b
FAVz2+Gu4Fc8/yIhHtifVUrMQLaYdcV+tJe4IoBWFaB8HZIT6fnd3Xqz114UU3YX
hPlykxwtfGf/7Zaerf6BQGYUll1EBs/T3UyHQoZEzlrQeo5z/er3rdTlEjJb7rTg
N3stKHoMco2seNWmOZoVTpyAYMZ23NyZb5DVxTCRjDKwodujVm8nNSJtMrB9MYhZ
Ed+1hopfH6N4UTz36qrPY26np0gu63K8I4OOGiO3SPBGs4KiUDHqI6HtuH0Etqkd
1N2lW7ZH2w80ZlQeKhFDIzFFvWa7bwpoaI7Wx1NHEW/Gtakys89JfHZyJKOh1o9Y
ArZG6S7xRhSRBVUpPgZxMxKQukLmD3CQBRqeNgYyxKwj6E/V3we80VIq7OTec4mD
jyN0G2yaIOE8cGexfgt9BzurEyyLef6KoaZW7t4N03jIhcyIE/uB02hAcklfxTPY
vtakvOrxv9mSlnf0WmYe9+Y3iorW3uV1tiWjjYHofh9msyKmU5KzqpQdXlIzKZXg
WuMHkugcuf8a+v4Jv0ULp47rikr+uwXiBNbyhY/yy2bllXg5PVgo/LZIO83zHr7t
xF5gq7tD/jlsgRWqrx2Ffs8gDSfhmV2YMM3MvciS91SFIToatCoG7v2X4IgyODU0
wFayyJqTRWsKf3S1SfgClpC5nQVkdeSk5ZH0FR9dNbXpEMz6msApum8RQqeMk5Tw
L2xU79q17I6qJD/Sy6zhGKPElPgzcMqko4vxsF/vUPgIp2PRkk7OcI+guVXEfLwU
a+wbt1qsCKpPskIi5aC8VQ1mScppnMrfon34cvtfPh3E/ABjShKOmKRrtBPVNTUf
BxJ1lS5T2LAzaLrW9peoBgT3aEu2LE1guPfoSceIMoEcAGisMhPfJ+FCiHIQ0v54
O0LWySqktaQU+0CnmtC1cm3FLzdApsxa9w3CgJ70bsn0wOZC67yjCC/4ugc/QdoJ
BLkd2rYCAMmFir16gLyrq3bfgdNyt5psyIoj0hTaytqbXHQrSTDQWAPirGzNEHtC
IujhhztywCLU1UyUXAMZddt+HatNidgPat58IGZe3DF5xs//VA5lLHTSzh8Z31iE
y2256AlZ2rskuR1Carmvv1L49+WgX+Ylwm9LsqcKs+BYU3CW1YYmsgEcSVILxYh5
JobTdalWuOWh5eqA0EtwiN8pKhwRT3lzc9ML79EuQxWKYwOriwSw+P/rt2QtvaC7
GU5iAMPqyXyBJgOTpNk9Zfy90skjKLDuMxEWuHqerhJDpO4Sok+hVhVOkFjZ+ADJ
NALDuw6Yzj6MTq9fqQR5xZtLT7YdGqwIDqpaxA3GOOP7pYgNyy2nRmnSr4IrWveI
HlDSdLzr5eMNGmfSrpRHUS9Kde1NDje+eKKk4rSzqJ6rechNZvgKbYiXKSljkrnC
HC3B09eU29etKRmh4OoExH4U+NXyYjaLGm1YGRg8m11W7FTdrBdONlbSR1qhKIPj
z4C+2pNf0eirOEWWRucCOUcOGUCPuqR88gZoWU4ph2rB+duXFae3LUDoZQRHX8yi
by8lkbFvixH/cuTBUDmuj4dySErURMTQWyGMBK7iDoVKUDq8DlDekMWaCaCu2f8n
ySxGhFUCxdgiLKaNrxxn3iyFXjZ5rsXvus6KcKRv/7YdV4Sk0JRFppShjUkmiWhS
dTKCcShs4yEg6aVxxv3JxsPtcD+I1k7teiU+vlUHVmGKq6HHZLBLHAL/LBT/200s
VNdApyC/j84KiG+yr9Q4Yhp6Zj7jTnnFZkXjTTKZQVaUPRSgGwZ/ukpEkzNRO2Dk
PnWQQZSoY96/MRq6g4JhM6EXc8yzr15GD+O0T9NDjG9uk9lfJp1vi+bfrKt7iFSe
2l4poG9hhrsHj8VI88Bo9Da9judMFnZN4rZHj1DrAeyKnGpBBkPVhfJ3XbwRC4y/
x71iZn+FyZhn2PJs0MwE69RtYOYAmdiAMVtWr5QlYuZbzAfW35B/V6f8f8fwjIqZ
MLAOz9RQJQTm9/TUNb0SFVbgg64NWzReCgv0raCDr5tiUqLspxWTzIbvsg0pczH8
sgZtDP1KqdwIPRgPpW7Av7U/Kq+olQfgY2kbDWWBBB0ZHo2Il6EzAK9uWlACNVZt
z/vp3OtTEFPHwJ6f+VZhsDsgCj+QqXDa/G/xh6bKeA/1a6Tqz38kqwZ9XaeSyXtx
aqVXzJTvJfMVyqWXiVEQ+6613qVZjHrSTw/5/09u6Suuol38RUIB3N6zGMzgttM0
j/I8CrGUAfF7sLk+x6EXSeOwjICLrekIvIYWSKdYg5eV8DdmcfPH6/XafW/mckNB
6YYKMUlKToEOIqKSCu7GZOcS4oUd9w0OIvyhFCPuH9DzCWAKFZs2jd/Yn1ZjLN2F
3KvqDov/Om4cOLbCz/H+aZ8wvWEappCg06lmMHcdpL/kexZXFPLWmkmuQXz5oINL
jqIAOuhgD88R2fBXIi3xFgyBDpltjT7SdyZqpHS0cfKD2j1uqPtUuZfI4pXjKXkY
7C9fm1+Ge0t+sSyKyY4+/IKEddOdItiLXQdbgSgjPZ2N5B+H8ir4bd9pXLbZib6M
ABH0/yJXHrrsS6e31AagEaVDczLelO3nxnwwPJ9HPYc2OzJ67JYb+nswn9R6Pxp8
WsjV10a7nLg8H3zjvI4YtIS0yVYo/yeX2fGPktnEt1lcY7isUfRtbP42KqaDU87W
FT1jzgmkGiGwT5qek28iSHazJcS6k6oFu9N2IhTSinEDWRbO4z4r5drrnB36RuYd
Tu6btmEx2wZxOs2N7oZvWRYQFI0vWTclfymS0euoiJ5Qr88dXCOgJGYb4MDlLwKz
n7H+Z3kf+Vq7cxhNMFPNpvEG50BFMyXMi1tkmUrMZM726eBQLADUenRv+hwEpOd+
63aoTyXbF1eZP9UHKTWQY64o+IuEXOkKNQ7QKloBaiClPLLKdsNcCD1h9cCWtq6+
yWk0efc0vA71b+MTNMPkdP7PQf/v74DE2PHIFHgeWVJhAs1+P+Ejp7DjL0E1Rqyw
QLZY/uAEt4s786UFI6XAE0GoRk4aaQpPii9rIitbk9I4EaT2ErwkHTuLp3LZRzDj
iF2fFCBij8IF3WU2W3duJ5Kopb6C9g9FpQzf+kU0b2rNcdGt7DoC+l5CUXlTFfZL
I+wJxudoPMM3qXIYDddd93BGzbnLjdAiyYR5f7nPFjAuve/YwVfRW7JFW72wowDy
T3/FDjA2X1s05kGimRka4u9iaLOmEx/n82XQXhYvjGl82uIau66SwwH76ugyBHc+
PQILNf9jej3wwk5itoblbuFaJnefpo7t656oeMgt8jxERdSXOb4DGCmP2W7zHimd
ODgesl3wpW0P8WO3uHy7AfciZzaXec3jmwAjkbf3IL7zNiOiuFdV3749F02gvANr
Lw+irWTPmYpQpwcSnIJ7JIp2SkaGOA4dbxWefv2AFqrG7SFYbKxloCwZzwFnt+Xq
LmEE9WNATeHBb4gLnmaIwVjAzvx7ejRMdjJEs38gt99RnEr8s4XJnGuhZ5rF9K6P
Q5wGyjzzHL7b0bElwiV0QsDNFTRt0SefUfPog0wpLEo/lPEyORk5L3zouZQ48qkN
gsfidh0HhN+9ax2wLZVpKrJjeVT2JAAOC0F98e9KvFNMbuBkBaXCXfsIALO4pV8g
8ESRH3JHR+3Qut+uJjeBtTFbaZKOEkbxixOXDgZWDzHVcpTIarldiclfMkLW6sPP
6Igf2daEUl7/fXX5t/kq/Wxw99okjCoaX2HDdJr/M9VrD/j9BDSBEw0zqVmYGxqp
+y/NH0+RkFz2xHO/Z9xnsYLYSJToowxzZ5bunVD4AIdalCTxcwjTmG/gU8C0zz7R
/Vz+7k2WfFCSfBTc2nAxtJEGlhX/wRhMR5Ec3sNUTevq2qX8FJucRQAytlKQulDn
7PF8ZOsFQfjxVq0hVWxBqjhsisSvpiYTSE2VKf8quDervO6cjq1n+Lnf9kiWAmz1
rY5OvPEkS4Sn5GkUdg4q/4q/CqsvekKPaKFDqgWSGrl2fnPX45g55Lt4FZPNhkFB
qESdqxuy1S4I4xO/Q/v33S4MQbon6oTibuSqvkTPHACEM4qLQpiN9V8RVdltruI9
BakdbJmH4lxqv9fZYhMCtja3J+NheQQoNwzazWs34XWAwj9DPNh9VgNKqk/TbRYl
CdP8EJybnPVlL1rAFN1/v9QPCoGBEBq94WbjPDdVlxxGdjMcZpaUc5+aexy9g3af
45UbqNIf+1cs4ohGvHwf/ulAPstxTZHPDET1Yu9YF6FmFgFUErkJ2s1bqux/j3qu
dfiW4JS9JLGIK0bUpHK6auwKscayXE6cJ3i1PZGV3aGLAjgSUy4R7XXQIYHk/lZS
id7AfqR2x2LDNLL2WtZWrRgvquXrnnWdxmn4hdlM+/cuUtQ8/lq/hys0/0jIzRcq
emWJNHFiCORTyDjXehc4pTNkNmBQkhdjVrF5EZ4aIZ9EQ39ku2/H1Y1DRg2U9WXd
3MZ711nuKgk2vhY7fXPoL12H0sg474fJRt3My861NRy+cBeQ5iv+tc9iktgII25u
+rbpJy0WGPy9tH9x96UE9BeX8fhplTOuso5kkrkbGujOmISEngGAB6SV3d3njR9q
n3bvlNEyYT4q9GgI50k9QtiDDUBrI+NxKvcZCS/g7WgKkqNvyu4oZ+Ta/lCnnSeD
yxCOxLj/23hRd51BtPnhDc2DL9KaR34yKrhTvv+4L0pi4ReJ+PEwtF9bF+o/n+dB
CH/vPrA6ltalVTSG2EYHclHeyIr7C3MNSvuAY93prQvv8D+kwOhfnV/ajP6eu7nq
BLLHaT45FxpkYqHmBgGoI1aL9XFtC/1QTVP1TY6RO0SOBOEZ8hZAGHSO3ETjBg2A
j5nhUIBg/qC9yHeimTP2W9O+bfTFexPW8N5zJbE3d/uPzg7bRwnWwzQJPd6E3+Vr
ncXLQ8FhJ2Kjv2QndbrKKNzwDVPba3qrEkrlwUZ420Ax/z7wZ/+Hgg3iYz1veQqD
rEwmTjaB1sFCeQJkjjd/wlg3JoA5A73wd1C0iVfxuELXlWz/AthUyrz9zqsTcpib
f9mZSj8La+ChBZYui60hlNkxrVZJMcQnNLA6PIwxguUV83cQfbz0ARaR+MhLH8Gw
7FATMyuXvXpFkNxax25u2N4TBhf3x+XrWo45OXEH7gYqXAD2R4LHNclKm9n2OI88
a+NLQssPO3p4fw3SRSXxzDYJXIhb41cf2JtsoFwcmdz6XJzha16OzSdfZTKKwqdM
mu+IxYjqb/3JcFUZx4FhgJ3NywXmTZ9ZdqjaUJ44AbSMV9UNNCyJ5m+0XcR7mra6
TMlwDFwT13cAXDQ8dSlg+XlPH2uC9jo5xKLmfju6WtvLB7yIqN9nz/PSNMAxwYFt
AyhEDWsOv5rvZMpUeKKOEvMCS9DMxbaiEI5XUWz/a18e2uqxd44BqaeKoBkOlJsj
t60koF9POpqNFWa9fyXQxddzSYhsQK4y2srHDEuE3wgFakPw1z42+1f/2s2Ti1Lg
deSJ25ZYqIQzJHNWJ4Z/z3zC+JXs9eJ9HeGqVg5ecZSVlqprodEFvgly77GVs+0I
SRZHzJ4IkSL8/lTctGhwke3jkLqrBZ7AXfGysR/fAZ5k1jL3DPZNar35+/5KBrIl
ZhYF672zEgUYJ4UtGMVNRHbFM2bcZ0O1y5b2JqQkB6WJte7ZHT1a6oZd8kuqy53H
jKH781sTAXSrlYAmYmqu0nfJK7UnkKmKUc48v7lsLIZ7lIMp7GkmT5g0hBGnZDmY
tKr1CUsHLQbh5pjc5ucNK4DmksOVaYHC61DjF5PDhUkftPdj4/NR3Yif2N1CBTzt
i8iaoKBdL5if03THQ/pYC6fquhxU+Dd1TNizHT0YnVQKSjaiJjl72H7/cj6U9yqB
pXS5Ma/x8T3Kf7fik6CJYiyi/WNhr1gfW5btZNDTVlKHCtK0o+OuGn6X074yqXwC
qrYNDVxzFGfXl/mW9pDAYS0+m4N7GRbnKCKnx/K5zfLxnQ3lsbYDN3d1nR81R2cZ
8LRBHzU6ufkdihv0TiJTt9WALMzGgEceNryosnjEaj3l++8LrXnetXaQmXqe9HNM
Sxip+Vz/ACrpQcfwq8Av13r01emEZckdxpPzwDDbegkfvc4lYVgZorH0rW47bBPh
eZpUjEd9okHhaqs5OEBuru8cHdp2Kd9NsvK97xnxfBc3jAU7HZmf4yCYhOang6FH
N6U6PwQrNnpP4kwyYP4joHYcHhQOe3ay13+iQE5QST8X1LGzLpK8SkTaqbKtT168
mig1uHxVsLj9fXAh9IDfp+wZLjuO5CNJMkfrqWZ9NwLXrNX+aA05njzAD5Cf1t33
di+AnkLvJGqMI4ASPmf61kNqAVkYan4nfqRuZld0lvBolpz1WfNMHnkefH2u2SZW
GFi24ef6upo2SJDK7XO464qikD7WsRDDZqc+iIB9OoQo9/+KisvtDjCCQ80YIAk4
GCHhw0C0XUEz+gYI/Tjz1zAdIyuch0W+OEtrPXc5i39CEP514BORB7j8Xy0UFp7E
+8UIyF4ds6MVoOulrd9sHBX7ry9rEzwZnK7y3+K4CaP+WsVZGm7cO/rR/UAyX9Ki
sHfxJa7rByz9Tyfsj9+PWsFnbSvjO29/LjNEfz9P9biIIKr3xxdCKCcZ0eISugJW
1JuEcWuHZxcnJOds2pMmWTkWxqVynCP11pxQjlsidvKo1GptwI8xfCXOFiJ8S8B/
XrzusKstn2NW/+Hhs18N74Ac3RulYPH/1UC722Hrl/1YaeYrtRRCOfo6I6wpBjC/
wSY0N9AQci6bLmDYkRoa1u12oREFPvTqz8HjB2TeS4E7HXMDGKJkKNfVkNoIouVL
qDiGqJNtvMo30G4Asm/HcLxsf0vjX+9dkCyJloPGnhbgf85ohJOs5hWOByI5pxu4
y6mSNYMRXp9DIsVRfZjtF2tdvXOC+UoCf4vfAOZuZBzUzDXdKALinnZl9pP6u8hb
B1JH/UPR/bA8upl91tBX/Bdi6WNdY7W6W6XMS8VgTCbvbkUKFTG0M+A6zkEhTQGZ
y5HPPIfnb6TNgzcV+Dt7QSESQKd7VMtfNtet6OVUtmG+PlcsRcWcXnYL5WmTbDFM
Zf5CXRkRvKnutNTa4v4PL+DYXVVdzTR9XIRKaMmU17uENLRRLD0woSYgcujCe+8z
3RfWagIQnc8Xtmgrkn8382e+krT1RsDeN5Hx0hMUhIIPcDx7Ca3IwlYuMC6ltClF
BFAQSOl5FZZR6BazqLKcgm9PVmnLuX/02RioSseWc88weqQ1Cnb1rSfx1HtQ0uVE
520jZWPDOVFRcIS2hkGs6csIOaL8enXD/nFn7TMwCjh9B+GRDRJEaRk9yozjlI9Q
T1LZOR9XAPw4AuN+w6SNhW5hK1/+918gbSWZYb6Zie0kGZaru31kQyy+vbNzbAiz
PnfbV8i8jXKhN7JdtFVOsnCBLRA4sSZ96vkvUbg41SKVeyQrXDJ3jbtsqPR8Tne2
zGOe4lfAPCiV5jVvEw1slAMNdkQPfJIK8F124pR7jip16JAW7NmhqJcBMDkWYtaq
YTivZFfGgDLVeRBBvOjQEuCaYIWxkE2e828o6W0m4fEQyVNTkIe1KVyAciHDwg2g
vsHt5bwzdl2qcctEh+ddcWQm75h2BkHh7X9KsgVktiv8iD2RJ57ytjD8o5Aa8yhB
OpEKfyPg1fITsaQDKiftlDfGEdSdj56w6GVx3bTWxovnqvuAOa2Z57+9qtYUHyg1
OitiJWKiUxxjXo3RprjFN0ajpixeNn/HpfZYDyT0HnS4OacnheC6mdi3DwoSm6eF
7zB3lz1GPiF6RgvXP3BsoCTtygtRSb6fz3b3Q+eWP3iegO3FH7O8Za4g5u6ccRnL
+PJmdfY0y50A9VU5y9kV1k2KtrCC2j9g1sjcH9cc04bco4f+B6Cy9ObUzVG9Eotb
HyGyJ9m3krmWb65fzUt8xTmk9ilvfmnH9gaqBBuq973iG4yKw7kIGVkUQEO7NUiq
EJqz/6xyQKkaEvrLpjS0CG4mCK0M1tIq1thhL2fNIIyc3bOz3DvnCB2xL7bE1d4z
BYFmVHUWjgZ15zfkbgHfDip2Ftj0LsfJWzyBXEYgCVaX7Dg5pPEejF23UotMgl/q
5d+5giYdGeU9D7l3k34XKDuUMLZXp/zzsnxJtfHbCyMuD5HAf6okRT+KSKlCu2No
nPqIYJVVRnFMhKaWGNCWR6SeCr3gCU4/w8Ayph48yHKDxNDOLB7IrIdEmTaQ/KTu
wyP58CSjJCi+11YgXSCpwCeVPR2teKqN9NseDscS9+TLzbfzn+LbC6Bx80bUWzvD
Z5xS1gwheRIxk7rf0c9yyEVVSAU6PN7QDo0YxDDxeVVP+WDvdP4XBrAfNIzADBG7
GrtL9GLxEw3zKJzdVpjRj5E30UL2OoUmLMrwpbSUg+Lv2etaL5Ki/sWHbyYbjqYC
E/hPPuXDvLSTPFGZ29TSwDacacltvt81AXnsoZZEPkljzlpy7EOmP1PXvoeuPFIg
ttySQA4KDJmCAd2oqkpHXK9eZ5aK4ZDQ8005wHuRRJoZJmjR3rXMWjg9LvqjPSML
NPvc5CZODFNbeB/wNJsa3qG1KYun3zU1AWw4X8lPoIDT6lZ1IpHPAlkLo6sStdr1
xcL0E3cYSbRQZRBQlll/OcpmMB6emPmgRp4bAsKv62MLHuO1flKMXeiBCKRdsPJT
Y+qBVzyb4Z//oFzB43eVE6iNEJKKV/r7uvKzJESInoBghxdz/CM911XwBZXqJlEo
VU1dJLpMGUoqoK2zptlgVOt9Z9o7K6ho+jLmnAyreqAe8RMsaOZWx4IFKP2utNEe
XMd2BfOlrv30FYIdln8f9YV2zjIyE9OWP8mzm9ebpxaTB2aJ2Zl0msmzR4mbiIHb
GSrCyHxtJOmr0BmRs3kgzur53FNyhx2kvhEeVjVfqWMLvrJT52QTfO88X9zDQO2k
JrrIsy8qJG1bnfoFj1Viic7mVXLK/HQivHB1/Vw4ZulNrVLOdN9dC3TVmUfPwfEP
RBMsiSn/amzZB46VJxVwbKTXO4IA7j9RmN+ywXKYOT8JPOq+436/OimdKlM315D8
Kmdh3s4tuwYEtCDCXkxhwJYScD8FwFVYhEPG2GF/9e/zQ8+RzaACbp5kJN2YZ/5p
R7HS+xdy4WZjmvZcDDa0b2OJAJ0U1A0GmiImYuDKJSWGj/HRWwCVJ4W/hNdkNoIm
C7QiXL8z4ZrqmsGjnChrTfNmmnzaduu7zwGMpQnbrxPNLQ7xB3oHb224Fe9EPkli
NJkbzErkagiVDREInbQ/6pZbsJf1Y0L8di+s4s5K1bIsbMYVDo/vkFAgHBpFehCA
fDTXuC1Rdh9qGrauGtJxYdtqtNj+ex1+/r85cWL7y3WtJm0NLkCYfM7K+MZQKung
MjXduXftBhbS/8AfhA8UU69YR0VuajdyAxCWa08/kY2AVdVU4mO5S0j6um13OGsL
GNU/90TL8fVnvBBnz4L1NIMQfL/PGehFruuMs4jr33fQBvXp3ahOMSUPcmfVHagA
n9zelWixuYlRCrIjemTcuesLGpBQ3IkgueanZVIwXKiDOmAchYNxsTKBXXosi45i
8GlS+SCNVL0T240O4iYtVKZszmARs+xfeoCpmstZnHYn+pbKHxSwPvZkFhoQyuYa
wd2tjS5stJh6FfduRbOcHMOZhL8AnQEaXoIPTCBQH3yp1A/4VcsDeE4OQr6+sIkv
9Pr9BCCOktbrB8Mq/C0MOwV66f/4oHyLs53ugSH3SUUJ2zY5cBotFLTGesvEMIjT
uhMfLU65vZJheBoaqSih4qQqju0i5XC1hGPbh3RXvUOROQYubutPRrMJQnNAsBHF
7wge1I/Gx5XWPDiPdMGjQnTGg+ysWQn9UDiVugxJ8KnlOKJQ6XS47tOqOtPT7LtQ
mUHsciirqiy6vJekgoNpu/Stt/Zoqz4HTS7dODi6qfBcEcA7y9XkKeuEtAWvBvcS
sI03x7QTV9rKVIMXU8ViSsWypIchMvCHMfvvaXzBUfn1wvPF0n4hkVoXjCyg47XO
PQwzhd4Cm0Gh92hyMSbD8durlX5tuzCMeKAGRB2dQQkVWip9coHMAm1VSoD/LVVc
r4oQdpLkRFSWeDoIp4KXwnw71TFI4I0u8zvSl6QPKxJjbuWRMP2IrvjiOevQ/FcJ
EFU0mubjEH2Xz+ChnptNTYjpxaGwxAt9PNtpm0Qc0T8UHz2bOGiYvHmdTASGwXkJ
7c2m3lbYE2D3Kfmtk7XUXB/IVxlXpQhp0cM3aQe7Pdm3Mc/Q6zPzWS7SSW/x/YoY
IXF1zTXwBrZLfQQ+JbKWDNbaVlZ+aDa/ybh3aFZ/zVcFJ+VFCYcV/nRukAQ49Guj
+C0C+NJrbp+h1shUU1vMlmf8u69j0Z4jbQkDwXwo2TMXhaSNvq94bocb/Wv2RPP5
HA/nfnURaad1NfaBZke2XpnVTtBxIPo3Oaz/zW0JuN5lqwiaSlqTaefnnKdWDXaX
UwkIaddVQfc3UHfpXDwZrupGdue3AuQYw9vdOhguRwj/ifcP7LZOG3QOSvkO1zJ6
LwxCmVp+OCNAtsY/RWp36eBW8hl5qVxcqMelX2s5P2gb6x6peCm2CUuaX6rvSh3L
eJYde8qtwzjq0Crti9DVm5VgZIOJx5aGlMJeTIrSvkFJRgaqu2bVuqs8H315UcM9
tk3oRB/37AqzmhNtE23X6Ki8vDCRuYMYfkGSw+LlH3BK7GSnud1kCIu5MQKsIZsS
03dAOJcKY1Da5jVDDmQdiuqLLlY8u83N3W01HMn8R+gOyzNyOyRTYgqhOpqwCSnP
fM2OepdwjD5mDUxCfeP6FJqeZXxyfQecYg6rdXKd19T486izgsjDVG4Ixr7W5uCy
GQFIahWIJLu4WRYQacWZgw1O6gRtK1uV4p0orsl4NRumi+bjy0XBiFufiz5TDQts
gh6e3hsEYyfkSKFSU/siz8bMb641LEqou27FxyeMxrdFxy5jOiO6eDh/DxRQK6N3
wZAs3TDEI0COezAzxHRPxVpQ440CRUPGaZddZaHA41wXP2cjLNvMtrb3tL+W7t7n
Ctf8etmVP6braf3l/7wbAWTkiN0Kc9zAnMrQ/iup7nWX5KChMruY1qWTDKAkmlXE
Ami8vBOEl6z+Mkuo9w1p9fX3DVo11un833bOjG1ILujIhSv7d6JVG+2bnrAwS+Ku
JhqCQGbb+FF/u3CrRR0NpgxxPlUW75DlL+2/YPr84zScsimrhNpcMcstV3W54CsR
BiCvjJxUIHHEK5lNN/w3R4SR1AgDnAu9fpLRk9p5HDlIdAMlcDB2ZVWA13UpVAnA
8MieOz7upEw0FmL+ohqdTNaDirmuyToy7pTqMJgbDcss5ghQVFgam8DNawxOiBIO
dbJi/Zj5jmKy2yGXE8NeYdhXd53+nZuRfjbk6IFxjE+hzopoPFbe9Rs4o0EP2PnX
J1N/6UNv78ghcwqAPuGbR4UuLJP7+LnceHTtrbTguOX+1YzqpWIuNkRK/1kE7mIv
YP7weapECwvKNMGIl1F03HRj/WiETqzOb7xpXdRjCuI9o55GraQjhb5YFcdGK/+T
cksp90uZiilpzourpdTpP2OJoY7p1QKLdAHvoszg7hYBNdUyLl0DGZ9OAhCKtiUD
cBIXJPTvMmBSTnNMBLdA+uT+4vN3TyIHAMagNG7tvDKNyUEC9aFHtPcZcucimqf8
PVpvRJpuMq9yxGlTJiBmAorf3Vp5XUKocm6zhroSuWWrRAFLUGq5t+FkIDLHCeo3
lNy98Ytip9F5W6W1KI+vjZN8S+dCGD9B5f/IiDkNh23GFpDxknphj5Hk8Bjrmkcg
3aJl+4wj8ecxk/Th/iponW/d1/W/ziHbDZjseJwcFvvtDj72vVXvsiTx0+li/pYG
H1qSub5VmOZZnFrY72riZizJetyP0iqKDnw0x8AgAhtuzRoXFgODyw+VbW7n4RIh
wS6kG4oDD+AW0aPw8wFo+5rFMV4SaM0sXqdTJ9XXCgQylD5fqfTxhBXDcsP2lJ0y
wz8niC9KNU9RC+yVRGoVXbhsbjyhTxhPxnmPa4/b37lOERvzojunuP0icq4z1HW0
YSqUWO7XfrWMYh6haeerLGvDL+WxFTo+j5dj/NIUAWP3w9i8vT0rfhCOintVDzMD
4PDYSHeYKa0L4TCeORx8Umv4jTKwLyyEdp1yVzst85UaIPej4t0ghSZZ7sOTXWwN
f4xm5h2OZlPCJSp39781i3fA8CML7yuAkvR87B93TDTMpd6B40/hTrNcgFh2BMVi
FyCmZ3G3hhIVeKoBZkvQbvfpP594q6QLN1ixShGu2cZCalmIT2182z7rNXRrekHQ
NDgcFszsvwDepQ6azoVMCpEj8E/QldfcAzG7a3jQqnpADCXeK/x5B849B+HHAwN6
Fgv8VUuyFwNduwgaVVNJhjlhXb7FUU1c5TMR/SEtUZGb6Vc1lNHqOqmVVs3wP7zv
VevwGcEHP1yxdcljajdZtLRVoYfYG3ewvM45BAOjQP4VK4UgjmoH+uzqWA/LqitR
1/KlHAk/I1YR5U24H6DJjTHjfybu/TEiIR+v/eBu1XTr8s7vaPvOwl0vHduU8aNR
RftvO394JCuUxrtI3BQUYSRvjoOFQjdmtbIqxfknrzFwFo5L65fSR2kZAB2KYVqo
BdDlhMWrikQmt2jg2cJSneRnDwoFrdK/gVUtLwOZVpujPAUTXvL4IJsqtzbHYeo2
yHwCbF2chmmikTQeYIZe+pG+CSYPxwgnAvGScNCMAT+0kGjaoVVFA999obmWwwio
gmySy4JxeOBsQ0meuZaR/jnDTmOmXEr27s2bEwBSeS67r9WI6Hk2GjOuqv8KdkwB
fABvxhFvd7upSHCxtqmb3jNslPutWnb+pX3UvddZEdAmbxsYVDOLM6vNBotuTnpz
AvvwQh6KROn/nJTxKJ5h1cPO2fb3LkZL5jRNEDwazcPkzaVAmN4lDB0Y22riZMyw
gB5/43hrWumMfHAkJEmzZbHi4NAaXmFYhHYfC2RfcGfJBnuir3aYnXgkFUtP4oI0
hDvl6cv2jiBSTeRX936xQp55h4OLM9wgg72oRdxjjZT5Co/XUZXm3PnhSi+p5O8Z
PZVFRKcDwj+iuICw08isl8Tj44t3WeNDqWsnMPTsh1DNaZgEF4koAUE+do5R1dsN
370giSzLRkeP8LXuRTqcyNFbwgbWH8gQt+glzHr/yq8JT/IIUDO9+k4LeYSFdNsW
8WgmL1J7EXnPvfEyi+th1bECilaVHrM1mZ7j+ye+DRPuJr/3C60ciQVtGqUv7lJF
wjsNksnsd2MjewRUAn7IfWEhaCOgZH2nY6m5Hy4/tnjq63xw45Egb6ZmrgrbgMdl
nq+yPDnBbdAxAkwg+eORh6oxuFVFJyRK9t7rWPxWdMPioMbpiXvW9Ir3o1Zruy6z
iVhluP3pmDCmAbT6yFSGefm5EfRuC1C+Zkts+c69NkGzAs4cS9jhrYKDpfg/hsTk
YbSWFq3x6loTr+bKQyZwHrwXcA20q1rKWi6TNeb8oUBHoVHZ57HBWe/ywAU3STYR
GW+iylnctiGEOV4eibp6c+ZbaKBCCrwteltAzh3/dkPmYz699+RDeoNWAT0T/gh3
uDSvg9ydk05dtph8mqi01rfiMsWFjhHLSkMfrzW1gZBDsWMwD3TTljuChXte8NV9
6wpmDPrP4moMgPbi8ykXET60A5jEly2ri1m4esp2GgX8hMrwnSZ2NxV57prBOzW1
d1W06JMXQNCX/4XhWs6F5WZxIP6mL7j8G3aM5RJyO6tRVulL+EX6VOd95E5zEin+
2ngD6JOx/5/jVLGnFR7i/wF/vVkLueQINSuZPr9Mx8tnGbpXvd26EwUrcFQh0Hbm
81uhGwHmOBnEQdBl5kdLQB6ZEhDXxWCwsVA7iSRUMpkTYIXlVWMkKkIN7OvlsMyz
7ACLUXHUyer20vvynMWpHe9WNlAJ8sKzGZkslZSRzyhPXOtLyGCj5RQ8oOubwUWL
1KofXp8BKa1PImqd9CjFvy3KnqoTmcAD2vYobn5Z4u+AGiHEC0scHa7fnbi3lc3c
O+hz58X761CUhu7cTWUhl/zqGgh+bEsfAhg5GnP55h/TPUEGsZSsZ355TaGVDy3M
Dvwh90U+uTBeIARfIbgp3ZgKyQNphath6vUYMlLVQBHNUL3uolpA0Q+MH9VJuVR9
oBL5e6NuY0YKeEFs2UmgaxzhumS9M388Sf/lRGDtS6ubopdCIii4bh6vMhiAs/Hu
YstRptbJUrIWXwnKJ70IoyNVPLYDZvnendNIIfJ7xJe1vCeqAEIGwGz/HKg38zXg
wPyqx6FKHmecwpueR40FGqRDdR+1Ubdb/ZgFkPkemttSqCWUwK48nObMUhyO/xAS
4Dwd3Zj9jtop7maM0IsShs9bpX/O1BWkL0Joz+xC1oeoMftKYTFFp7JjQUCXyIW9
q1VKQ/SGzgaN5Z7zA26Qv8/GYrhj3XkX/QUYFD52y70LaSWbxXDI2xqMscE8j+WH
DVpbosMmrEaOsrwybi/QuQ==
`pragma protect end_protected
