// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:17 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
svXqU4JfEU4yLPF+agNwgOGGspBdMlC7FHtlY1cS9h5hYzhxKnFyQ2dncAx4ctCk
BmKv+nBAsmmKVEca+CfPFVPGBFheRCNjChvKwnNTnAUAbfIsosLoZ30Yc+R0a50n
FGmM1J1cbVKw3VM9ncm6S0Y/FNOMqix+lcPJ3maVF3M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28640)
XyZXl6X+qBCzWMwGEtPjFoyC+CZ99djf1U6bKcEjh81jkv2/NP4FNIV+gnaUNDdw
TmI9PKaLjdDtEQpxIO/TktWE2bgZFqkOnFEmI9x6pZpDvcCMU2oxaZyf5Ramm/0p
bws7z2XxURw/xcbZmfonVrt5uYSWh9Xht5i5xsWPMM5RitJvSKUCpQlHhSCMWbpu
ZrpfPF9vSwUjY7v2A9KxJlxQfYXSWPqLwBG1FiPjQyBcabw6eJIcdah6c0p365Ud
oZkJ9/55syoDHrFGE9QPrgerrIRX52XOr48jGzcx5O6O3H9kt48FUCeG9JmMSq88
GX/ajQiPxsPw1QD7uFbRdGLjYI5ldTsju1QxCPeq12rEtgPihuGkkH7VTDZ3whRh
oy3PaDCbmroMA5HurpPJ2cNJDgT2T6PxJgezJiuGkmvmi8/t9/xdkYAsNyUgtG/g
8v4WL3phFbPNnCHRQUS+L6c8DNnERZc/4Nh1uA8Oe9hWzbulZqGjuFUW99cuptqr
OIzqdr+SZQdGzmjrI15ZoS6wX6gk7hqdV7cIqX80g4idYaQC5p1sNY8TfeSV3uNa
KgTDsVK7eR/C2eoIlfSyvPaqPES8AIaeNa/QDVX6IFRmeI16YBcVyiwPYXznycCm
/ByH0rLF5H6rqymGT+FpR+PXDMRxiAVeCSUpiDCmNyF3cd9AtYAfkflIfzsahmd6
wtoCsNUfc3i8eDe/4VFJtdbZdX8K20T3OqfSP9rFF1Qn5Z44CsTtKZzMppQcTiQu
TUHrcn3Kp/1elnNn2SgSsCZ7Bgq+EY5/8RorCROcV+wnIzg8x1tzf1lNm7Dj9a+8
BUtSY5YIrrYV57yVeja5R2UALhm/C1zvXeelGOuaFKEW3pIBjp6QPzI0sYIItAYK
ghXtHCtYNJD7cDgIEx+Dat2dQEfC3CvWSzWmkQV47xAFNN537FuGtDH9+TIHZOMD
ul78VGrkXW1jzFQtn8/ah3HM0ZGuxPTQy0Yp7ulIiGbU/ryOYwyoi1LQAzWLmq7Q
khEEmxEBDJU6TWEgdVUdJuOl++tUhDwSC1pLhgYsoa4SuSyzl68RXi27Go5ysPSC
m03QK68boSSJAE8nTui1JJtpN3zi+Dg3jElscxvPItYMpPz2azWqN8APJ5RuyGKE
JHWYWSiOLhe7Xw/zNoG4BjGvvsUUgk3p3UTVyeg1NTt0/ISfMDKbCISwi+NHiOjR
AtviQ57CY3yksYO9gGbBT2+4/GrWFWjrYC3XvBxfRDwQ/iuZ4VjpMNdAS7vf1GTd
gs5CyfcIAjLBTZsu6Wy5OWVbzhj7ndnqSbd9gANrhlC+WH4x3XFuV54N6EwJHStI
aCWoKu83FwDd0djjTN7u5Wm4TGcc08QTWgvZVfjkpEnYdxDtS77p+Mn2KhCWXZEn
oMDZtjbj3ljh2UWRvloUbFklwwrODcy84CNiiotSZ6/+x84d/6opoAg/xf3wHBBX
f1FwP0ddn93e5yrGsHrfeIAymRg3H9VTSnxpU+zo2/gyLsRxIpQc0FqVnyMWdHbe
pZk+OoWdmHpeN3Swx2cUkaG8BeNfQXmEWxDPd3Q3YicgAcmO4THaTLSvpAn7KnAp
Yd92J084bY7ij1Xeg80TrdMK0SOnwxVtNnhZGq8ndUvcUrEfF3pW1YDMDj5vaO09
c+grEmN/+crTOzbEocCSfK8Uy90rdLV+6d3r/BdI4Q6lKbJ+xgsZ/2oMT8BjeErt
Wq1WSHEylLOtd1Xhc98wxZeCBK4jaFByxtATTE4q5JE0bPiEe8G2bcfNpZ0cj2wP
FQZT2V3F5wdTZUIaNeQ/YGBkl7JHEjAk8LEL7OfzvfroDRqkEU281uWDN7MEUTdw
2X8KpSlMD58j1jGvGO4qyNo+72hoczGintDDBM8c+2jUezALmMSioLAJ80I/0eh4
RUlJk0UZ9FIj7/aWPH+5Sk7GY03WLfOKXYmVg99p4SS1OZXVoWnw4pk7By6V0bS6
Uo+/F4C2x1VxhfOrulHrAfNJOmiOdSWtb0XRztO/cwYp2lrD+o62xXYQuYcClMNL
6U7JAyKCYrf1moKsPTbGhtjDQ7yQW+exOmZ1eKMeAAVAlghR3ZUF0HQnd4q7O0WL
Tj27O8yQsuVve/dVNyJUzk2jy916jDaX7Q0rdANMFV6+gxE2ynd5KGMECngwnWp/
tYmBSxyOpYVUKhgaA9NOALF/C1oOXCO3Kb6ZBYu6RnAI/OihOHVNOBb+WG6RqXfv
a0xgQje3F2spqU1Ohsdb5Jcy+pEggcHt2hxzfCklcWVf5f21z5EkUchf/v8tu/e6
AEdqZou+o3d4GVQA4ou3vVCfqG5vNsZjHAmfA6m/8CtrrZkv8RmGgBkJdFweym8v
8hkwGYAtkXQ6ihrDUljjQOjeBOcI08fvU+WC6LsYj1fHoxdOexUPj8pCxeGNQxmu
gqC4tu/yDVQ9/oMVim/PK7oHM/OqY6PhWJlodbi61GraX5HskVWinafupXcaVl5K
EJoqLDzSwENNO7uqRqASAD0rsYWOXoNoGobd/DXk3ayA5WPuikQ25Oet6RW6mtbF
zwoEkzAwZ9dK/O0+7DjfbqLFu4C9332zDoFWJJbe8wJArDfsvTGCHK6srXTPro7q
JIH91uIMlS1yJPhbmzpcnmi4HAYSrc4696DXrDRXCKc9i/nK/tOryVVWAYICdrP2
3tMzbweURF7Pa50VRPVMho0XZXAKmzIZOggiwLxX0Rt/+AYtXEEaSpY1YWnORRkC
RiefamYIl2NzHvxvYh2GnJIgNBYxubqsQBMoAqSFIYZIWdjlbhNMxrFK5YWymyxk
8nnM0hLdg4asLypssCtchGar4O3kC3POVQH6bmhXmNarMBQH3vVw9if3XitcyHjU
ma8zQ8BTvNl8iAJ4ANTOXzM7h9zj/uLQ1edSlyUVY4MfKK7zd08Dn7y9DzmKJpzP
ZJnFOxi+hBch7EpqRhYV46XhjwUqOX7VdjJDd48FChBMrPj0l9LVJn6wI6y1VtjD
hmonUf2K9LDKww4xiqC6lPaGtWiT9SMai2tDSN7nR9U7Yv1iSgCQ/IWVPpbJNo2N
zwbkwONhalkc8genCUdskGjc1ul2RJb/XdDC2B5fGH73hxKsSjdd0U2XXzyS4H6+
boMYSAR0ER/ir/rX36DnebIV0r+GP0ZOor9EFhSJgCKM3b0Sx1QT36BFTO+eCGri
R1ZI7Y7vmSZwu8gDplqcyZceOlw/ptARa0Zp6dZVwdMJQ1hZL9j64Y8e4kvzdgnF
JHNhSnapCaOAHludmjE6Yajq2V8ljym+VoJPy8N3UY2vscPJgQscaqVabzXkhHOf
Dtt+dvfXOzrxxvbqr5FoGmXXZvzHvc45J52eYFNCcMVlMECXebiVbz2ZzOc+0pTV
ZeiEasz61YB5Ypv+lIANFX1ETL7FIdt9MFcYSD9s9Cb7OIOpFny7BuVftJRz2tQb
GJnViGo3C8uBFnkTuSXFxOxkzSAHd/WZj1jOP/QnozXiVIKqxFm6CJfUiPzKzQFu
XArWq54W8SU9iSeRSbyeBBR8i2FIJWo4tb825HkHhqk4FAyQvpa3/MuMMP7LcbFB
Sc8ectqJcG7Tbmg1Ie4hfGDtpuhnIHZNOWXb3bUDUrZQecAVG40p/UipGNUYSc3t
cpdp/LhLqMtIMB3PGb98jK5ySPDrhUVpDCXdqDaascasUJxT1/pton+tSH/Cqp6U
rO8JBDHizWpviWBTOsmOEMl0/rM3auDn7sqdFJ2c4DCFlwWruh+6O/98MXNnKjiE
Kr84xDGNhCYALyrorg7HeKSvj5oLzvi5+VuOZp8Yd0AD/6SLIJaYySQYdeVujnEy
tzWFtAMeeY7uSm/PdFqN1sav56vFRW7m3sl2vbtM671EtEOj1Vz/1bNf777ruJtI
WpDzQd03hzRjdiDx0Vi0W34na8WUkFNoIDTvhLiyTTBesfpZslr6YGgCzY+oipQO
9UY2jT329WPTuAYDlT0MMc53a4K8j/Cqw6sGEF4SBykqoFNY4PX4DGL60AD388Oj
Jk5YrvuwwugH5tgnMwQtr0zI8n6O3k0ADBkW/N/TgN3lIo9w0ekQnbYi3zxg6Z9o
xe1vCM2y9jwgiKn0MXpoxEHe4CkxaaLKuO+z8hqbhCE547NahzKDFUANQWjZNYNq
KmdInZZsQGv5vwYD+XYedjoadkBNoKeIZhkMkhtSBQEyFNp5h3qb3c57U1wy9QHM
DS04xaRZX/xHFmb0hllAx3Jr4FijiKMQng2yiYEshziXfdC7RsNjBaqMYkVV9Ty3
Ot78MGq9fggF7NHylfXuW8LOLtbsBkPO0O0oOObwFDpzQtfU2RaApC6wQiC3ZS18
8cw5ECgItdaJ8BQApc1k5CCbKuEIXcRzed21zw2puRAJzPqBP3jZ2RF0HpjfxguP
5dbyFDOY3Kl5vcb4e2pg/rg1+3XFlUsB8OV0tOS0/w0bdHzbhietivojGabZyA5D
QBxI0YNp56BRZ3bHKtz1M+iu4YGgUre56AWjUO1P25rGBUSCXt5WT1RofXwiRdfc
YOt858Re4GsjPlE/pdeowyL775ch70jq8/Iewgvy+kEUhqL3EjWtqIw1ApwtwhPJ
iCH3GJIkhOFXuW9P7ce4CkqeHdk916f5JrYCy32YopHhHxoCeGNjj+DQN5sKyYoq
04/s+0at+gG0CTsv9FxsNS3TFM5OdW9PhdU/UE05mmnu1XqiJjrSkZU/OfwmUyEh
fHthmZeYOj6avy8IVy8p142qisi6cWQ41RBIaeoNnom2a0DbyMOquQTiZMp4hshg
IGVruxRBbfLuGCizwFapKbYVtsOchJ98DMUXm5uJj0YUQLAZ1g4EVpg5IvzPXHPF
6jgxGcAI9uJc3ENyWeano6aQh3Vx8QAK8SQTsPJDTFDSLjsCaxFuppqKPXNdftO4
L5bsSq0B0zGHitM3Sl285/S6eoPeEhSXhMxqShkdBU88M7KWoNjjap5VLxGGnxSu
bVt0NvfwhWd0WFL0k+v454UCdakMMtGn8gqpUoZyha58XGykyZuQ22Wmfv6tqYvP
p7e3Sci8y71bayPpTd0+yR3GA8QVFX+l0RYBnmMMHFvFDxKcGZ47PjkF/F44C+kr
bKDNHY3i5vFgnLKnVxRXWHPoAsDJT5waNqvTlCElqUT3NKNg01K6BLXNBtn8ztVq
VOkS4ftgG0RktKkkMxK/R+R+aOzKsReHWcMgAGkiI2kpx7Ovnz8Io82cNJTZBT/K
DalDSPJcrd5VsxcGnHioCpipokX8abchGP4gNrd1PdPBKAdvbh4iS6lA6l+ut5An
EDfQa5fHJr1XMIdWkUTCVfSbBsjaov+Ggpf8/ZeHKZ8KEcQADCBZVQ13lvDbGRkL
01zz5aFWQBgwFI8JAjR1Z1GiqPukmBLbHGIoIchhMzRXzByyuiYZV6TMVTV9lJOr
GABxceGb/cCVWWEGchokd7qR01Bfgkp54ebZ2K4CaTG+uor8UEHiUjj2oDVI7Lnw
HsxBE4+0oK/BmanfVAx3XBNXMyYftH+dtn1CPmp2uzUXyTvC+1T20wvt9BFwA/xX
/1YyYEGR0y9c+iVCbsPcx3wbT5qVNzOTfijFy7Z5p2bsKMT7gyWNPJClB5LIcaIb
oy9aKURZ42IsUxCeS2VcNTrQTxtt1qf0TvQxPG2kpzMoc74LVfkHy3RlAEAecFgo
8r+1H+VhHp7PPFqRVzw8r88DFnNB+d6PuyIeIPBxbwyN3Zn/cazvvTa1zZrHa9xK
906q9W/qmxLvK3xV4qplFYv3TJ8F5XU2WPyJHbmFytimAZCk7MI65HrzqI8cwNFc
gf7AS5+8xb0Gc8P7XnHFsEt2s4KUKjBZxxhG2u65YIAwnPfoUfQt2pt/b8huFqeS
u86j/EbVA+yrP/xesU5LJ8WM798bM7a2+YJaUs0OfJj6IApmKN1SkF3+nTelhw+M
8Ubm4fYiZtj4b/i9nt52crBeH2ukNHAG5c8/39/iMoqdjjuAAA146njEniUPx4uN
zdWiZlQBvSqs2YonkNi/zWC1j1CsEnmEU7A5uJ3YARoOJAgdhsROjWYPrJurRv4L
Z5p1j4MYFxOry7ENPAcA9MvFeK+Lgbhxu7V16ER85zyv8LlcxJL1hYy/cXFuY3CF
vK6Z2lg6zDUj0yfsH2q8VygkSn0bnYYp20a6mX1WVW6bHQKYuMPjZRFNQjdIzotz
gAfHJGqMKf+yasQqYsOH33ok6A6+RF18qre8jhewJ6WQ+zko2SZ1CPaQY2A8z9NH
zt7cL1LNpTkugIaWAlzyB7w5B+fLK54L1MmF9Zg0wV7SGF5+/92H+iVIu7aGSauF
uIvUZHXMPPGpfidZeWStS7ovqbc6m79NM8X+33lbfUuJKEsvvD9BBjp7+0V3hlsU
E7AlzRc1aibNAHFNb4R2QTsuR2JW4+v3bmmgcIy60+c6m4YEfMTxAQ168wyNDlug
7zHYPSskVtAZW9cQd57PX72tRCgXruQacUxl+akxca5XNxp4mXaeK9v+tWXxfXXD
whWmYazB0a1NZcRhmDfM4ANP6K0MgT/U5PLfyux+7MsQcLc9svbgCqKrZuM2fhGa
wKEnWQ/fPuX75P59yGMQspO8T1yxIcS3w2/nNzafFLS45J3pW/6jElLH25s2Vv+5
iizyI3a5X4JOZf/tLbDnu3K4JrBiMzc7xTBSWyBmNtR5xkXqlT3MaKzALB3OIPxh
HzsQenNUyNaCSp7vclU+N5fy/kSj3zO5xcryW+qAaPi/IVOiAW0TQkmlCZ26jicv
JGJP+Tz6YmB6n0sugL0cz6+AIt74V4SjfPccBERbVeUSGaZzwlCG4ZRjGskEvnNE
uJ1WOUQspcNIvYAaCEic7Arf27FlT0IZYqfAQ5SgY67DjF73kdwsyuyRbOshgZgz
DbO75eaKVDTSzjWXX1ztQOU3o4LDTjKOrPCN4qkfQzkF/wCEBumIQWxP58t6ypqK
B4xmPnj6NhqzfatP+T5dfmSg3wP8Y5SYyBhFZ/dAOErT2OXg/4xucqMsaQyQsHiX
iwqdbsRTcHNF+Zi3LtptwARb2xWY2EhOLE9OksW4towdbSavFHps/nso4HNuoLzP
F4LsgvzfwUawamMT1rayholRmP179HoqqY42T97Ct5hzePc/opXTGQ7tm3IKhiFr
EhtkPaEPzJG1XkwxZKuUjw/R0gzSsxkxoilnckVKvRFqY9vdbR6E6dZuxWkNkixZ
CzdaH9j5acFGX6u1Ry+onREZk91STdf1wfpJIhyCoRIYYhhJoL1U5Tq6xJ/oo3Eg
6G76e2WWOcE2G2YggHrVUXyKu7Y1k8QOxtcv1g/AYHmFJuxQhRYV7AtuFJ9Fka2r
X1Cq1kF6KnYZ7FMVl2BidZgaFlhEDGI+Y4Ke5HXOxrnPh06I6ChhxrK9pCpvLXv9
xs7pe4/myxI6BLs+2OO60GFDPwRJSpaYDPKHyIMUDFfbtG8B4g9FdRdFFKKdxBr8
TLYgYeiZH49T5baRW/DD3A+rm5RugQgcZRTJr/lDpZlfybx6688Ap17kjqnuOsqX
84nabakt941oHfrOaZoI8vohq9TQfRE+g+6cYVdNlmZ5jhh255JSPnxPIFsWi0O6
QWOr3Y80oYEDkkSbp3DbkVgz9IDCc+BUGBiBKgowE2HVr7EYPF9Xg1E4Xx9H51ti
lGFqd+v4UqAx+6Ftn4dKvyMBTEGBBazOg9tAgnz+Fcu+z4GrL3l1B+HjZ7NqURLx
bATjEbXLQHeuYbKGRJ74qiXQXAbEHwus7raKg/QR+xdt5PKOFe11AUcIKxMUow+8
hQxXXj4fVIKM9P1gP18NyWj3xt81G0bZ1DQyLOCIxBmM6MA4uJveI4Ohz7d8p/DJ
H2J5SdBl9M3KUldgIbhPaq2kjueBoW4fiT0lMrbzTORb+950UfX5TuZuS0IynOnI
+yvndzl4i6PkVCYS3oNcQh79XZLnqQqCVJEMqqMHVa1Zid+eA4f83oTzl2NUa11M
iN0FAFQp/m4yuG0syGK4PAJoZcJA1Yjyz73b0PMq+lU2YuSUMtZZelTUgaY7syQR
gXbWJCCbEAvQ5qEbC7zYLV9hV3CShXl49wOCTwtDzrnlFr1Lz1FGDRI0WnakVm65
vIxo6stIuhwwED1vRQzRqUZXjI1IdO5syB+L2oOEMi9vjAfJHB74JmMoPi0cnlE+
EU/0xKhwdbE2nRgpnz2QA5x9znEn4odKdV3yR28HztKfspKVCeDYB8Jiiabt1+0y
QmYpr9RXyQPUPBG+WysGh0QQrsejMvIr6OFAvja8ESvZW25P//qR9ndo+b3NxzeI
eur/o6YwcReFUso1dEWKpvlsVbao2GFAorB4Ef9/+r9KfPCgJjALE/BNha6F+9hc
5ESziYSz2yHbQeSpGHby5WXrFWAycl+CeyZdo2NojgGuebfyo3h+Hh8r7KrVVvga
vdZ8/YfPStGqh3kpwk7LLIxo2LWxLoB5MRIqyij7bbdo+XE4szgVPg+N+d5g7gEE
4sXdEqO+BV3jfdn0SnGYuSZMKhI1qanxEnTWBxCGdG2G0Slv9uznpjOGIn1XI/Kt
3V7CcOumVx96fqJHPln9hiNyLxgNywHQ19WkchXoW9cYox4/QTYQZkyWJR8lNsRi
jun/hmX1aZamBIttA3R3EihDAuCilqQows9674c4IrgHmEI+kskNIvivIb9Eemwa
gmQEeEPx7q2RsSUJWHirDm1Yc+9P0+fcDydLqvzlmomVUF0GdAg3y/3oGNRFshDr
NwskT+U5mCp84lRKxnp47FYiUGERs8biT236x2ziwLoZ2XIDyrTO+THk8bJcFXEp
5yrSJQTQ+69llqhBKlj+fIjd0Ikxobd2M/okPmS9/x5s0zfAbAm8+imbdQ2niW9P
vIdCar/pFNtUp8D/sb3ZDp60l0bMW81AntZXnWMlrYtvhsWV8opezniRIJ6hh7x7
u/k0BNCAP7KSYd94XeAZ1AAznn4rDSjmzw53rdJoJAHKWanZoQxN373uLy3DJx5j
Rgjs9BRS+dJClLv7gQsQeik3b07c2NqYhQJqohPHwH6lyGy20nDi7ocKQRwevBq9
QT761TIPUsvLb8OZ3unVT0bZ+xdqvKmzvYFhO4q0hd1BEOuoIsQFnBjcN2GnZIJY
p3HRvpR8+rz5ODXFknRqOlFjne+64bOVJxE+rFlhZqdVjjhiKKbl/ysejoSiopjb
5EXzVpMf8gS0VatHlDq1nzJGELpYJj7haUyfUPZ+zuD4ktexJx69D0vO2ztd0y5k
94lRzS80tIYhn6cHVEj31B7XfS7Wpb2wfR/EFiE55+9WC9jCNw4K3sIHbq+lx8S3
f5B36PwUH2RMxXDOfeN71XQp2lwBRHj2vJmCPApjmEtWkrZ558+HeBvEgtsmdD3b
m//3ZSI86wuOLMon8UAa0k/gcGSeT8jnMImDD2ZLzFBNuRkoGkWKKo0U48sPO1ki
G9Wt/V+m2cKTVPxcA6KJsZML+kNqH11Xgp6AcmG8eoC8lwVWmTxOOLx0CNGJzzjI
OFfWhn7WsKzbIyPuSnu5ScGLqjQw2qYrcDh0ILFY5UaC4xpo9n+E4jTdbUEgPpMt
pFw5HLwKUZsJoqDHVc2BMQynh/Pzc1x+bxXiMKYwlWKrag04VKaItpQ2/GxQ8QWI
t7CUFXOk+gWpN3bbHlMJQb6MpdZBb2EkV1l9MIs6q74RVXXSsJCVVxaCHZ34o2kb
UJaGspHSZ4lZrNZEWoV9y9pZvW4S32VmMxNUGOmNZeskTo+XwkfWC6O4959Oe/q3
FxhcXrSZ21QGxETZCNybPFk0m6aEKdJ/yoJVLhy7SEy7+BxEibsxNxDbfq7LLKzM
pefVgM6sYuEdrP2t7p+XvmWu+0DtjFSee6SooSIiwdGBLUl3PvEo94ZmIYnpwoR1
Jyd9N78rN57TxMCk1loVrU87aQ4udmeM2JvdTTyHg6X9YrcRcZqXQPCjG6BAlLyq
cNAo25xxXpzby3jF7Qc7qmp8978jII0lHWDvYv6joQd555WCdBuohwS1XWqinZ+j
podotjh4xgLA6YlOaj0KpjQDvFFfCEt/87YZG9xxUyqZxEgz/T7P20iMudecmUNL
RB5roPzVzkgZT/jXrutU1Xww2aCc3tBULvAaybIHpv4u+T4/DWR7CTC0ccYnDJBC
5Lq5uOC5TEg1uOeinKwWron8PtrqUE7iOT+BqstDZ4V8fOMaduzpcXy75ySRdNEF
RYpLyowBUH6qc/yhtFKJMrBVScOBBUT1uY5FII4X0kQtURG7XhcUqTxtgeziS9cQ
YO/QfnDEihT7NdX7K+8YhUlkLxRBY7viW6foJ/mqes44lFXe+3a5UoAzQQGymkNa
alEc9DHRt71K46M2zI0OJ4hW2kwXZ8YhRh6xwMgoX/rkObnkqmRXUeGfpw4hZVwn
qUmJ0XW35PvUK4b2RxfmF1vk7mioVscMYQnakcCOFfWq5LqgfADZ4ED0WA0b1zsr
4uJre07Dtj84/Tq6REq6/O55p0yZveauqXjnEOhUWGXIo6wdFJyZon1KON+CgXLH
2/tEhevyLLtepuAcXZCZbvtblsQa1/aM5BvKlN+NTWf06BdbSljyVnWVwRz9BCrC
UsmPAb2o0vqHCsXaFeyHfzqaQSHD8iPnEVrtTtb7NJKChN+ZQxGPb/rsDQhpv014
zEau+UueZubMycFnv1zQaf0FsZrDGzcipvc9YLSUn0rk0ixRc+2xXyv2F0Cwx8b5
GxrSXLBLmVcy1MdCbREmZYvmTqOb7Ja+mV86BBluqkSsfCE+ckFllRl3bQzIQZZ0
TicxFLzkYawUnUatjKxJz0ro7gQhntRVYHFtaBH/0XfI98o/v2LUnGtLVQ/bLPu3
mLapJt+7Kg6RUe9Ts4PPXqdvCtJ227iHLP38gEqgnUHHsWI2k7gUO7vjlTpsvn7F
t8yiWG8U1ZP2pFEeY52nv01pexpotgQ4yWc/w3zWGKFNOT3q7l+wWEoqmbMfh6h5
4mz+HMVM2aWk0Kvl3kk9iuNrbxe1Eaw/Q+o5iWV4ER0QingPQjwuq04KkNi5ywJI
nPzxzGpkb3VAZn5mEK6cYG8/+xD/X/CQHS27eQBOWRhlfc8sfMg5to9bnUcHawg4
1imW4295sqhjZLm0yhD2fZb0GakuzqT3Re3GOgE0ocmKl7DyYJ0oDHAI9tvmWgBW
rc7YIEP/DntBg012b5MOI7waaQ1OOSXJM81GeXKknu7fQfT33wJY0JjpYKwepT5P
GNXh5ubQEcnRUuqlzM18tmUeemJSN9UlrLy+HUj5vY0Hzm4zhzYAonUXDwQat/fo
kETX49NOuTRWyMl2CgNY7ZLsALrg1/rlt2SOwfbFfugsLKWKffUWpabTJCc/F6Q6
WhAvRFMbkMABSrAz1VMWDRGb03+EAKL2cIP7LN5aPYs1VqNSRc/a2hFJKIxu8hZu
h2QnkW9QnIFeg8b122Xm5mY4qZnNPfryiLaJ8X8gkhDLUN+5XQIahyT4lzSBw+TA
ycX7N3SUhWnGE/2NwGosLstmV6EmJq/14Fc1BEDhYNUEDZVuS/TwMVqS5ZmxbB6i
7gnwIjzYK77K5NJWJS1YM3YdjFrZv/j5lYedaPmU3npnvLo1GXfGHeeZrPA90kkF
BYoWl9ia14mVOx/6yC1vlATybZKUFIkhXDZkGZizxfXyfFsA09sClDha5ZI6W9pm
hUD3okaV2vdC0GS+iAUUmyi9lZ3v7NegV0KXpJGTWRigoQuRa5tmD1Jnp+q9+Dgl
pXTVpmAOm7N2XLGLXVw1TKLBO5FLNNX6v1dmgiXo1wkQoiZDk97+Dxm0k3TH5mdK
0LwvnN7PcCaN671ZcfjKJmddWOrdKzc8ElsRyeoLQYe79ctxjB5EFvPGDDreix4m
QIu2jHoqRYTIPkiTmTAga3VLjSKYeKs5hK0pUfXm2fl8anSexUg8XJsAIwbXgx2e
svd6nez+juneEh+4RGDIdG/87CmFNS140yYcObrCPG54NzX3oz8nzDUzEXkb4aPj
zYh+fgEjS/lsINjLXlb6fMVWoGrDTR9462Dx/hFZYfJyJTnbOhlnH0yYtmNgrwyW
fxHeGczSdmm0LSsqTPLYqW2nInwydMlNaF9THoMbtGNgmS0/JJ44VLJSJW8zRsQM
LgHWy0KpsWUBbi42qcSmBjAp12MEOGqRpKVxR4GiAHNQcGn0rv/cLkNmWVqYx9a6
+ImcHdM8Q151quL8Yb8/9BQUGLg1+3cFmu60Bcvw3m9iIaFBGS+A5ZJlnl7xNRsS
/q7AL6j9Qb4ZyuzaWdwfxJB7K9nO6jQzzAuZypmLcYTJGnlXLAXRSeJRBfXkIb6G
bfhLdvwMX3E8UoPZGVaRz8lb2myINIlOJoL40ioFzTUAxzPofOs7oibaKDmj2MF1
GiffRyRBdZYBNi5HkrRCTdKfadB7DmDZbjwVuL+2h1navNW+R9SHD/LrT1N5m4xJ
qcvRM9BJNoEBcl+DBUwqlmd/VY98seQyfUmzsngURfaAsWVkOb7muxDc54+sWcBq
io6ZFEPL1uhq937f6I6/nxn2Fs0+1A8CZFNdZFhI54RcvmlMO648K6+Q86F9xAun
KmMUjZ429oN9MT2C0f13UfmDO+Ml/wSHXEGgyxL4jg3xS+g2RtOao/AoaALsiO9D
nLXQGRYZxS9SCyNL74zZ/JqB7ElFZWBpPNnZJANAJ1Qcq3aW1KCuXfO+T7+ciejT
9iQyAn3dFZZ32hhP8OJqFD1PXXmMlzu8EpQHSU7f2GHZ5FsiYFcWbOFN9gCiF8It
r+aQKPSZzIjD2eclDZbvZKMtfb5Y2w1xbeFPrXKcfB6X6ZBLn4K2+ISk4lrmNyAc
2WAEW7OAl/DyPCpyZvQ38AMtfbzgsWcbbh0MoaOWlRt8ahriRx25OrNEHmYJM906
Nz8aATqjeQdZI7EjWAjaySqZ3Dtdil2M3vG8iEa70oO+Vq2+83AtEjewWqG5Zzvn
ueWFjHWkW2HX/pBiZvsE4HGlcd7JrgnNfAOuXcFXy31KinWP2PrHRL58B3QRNLJ5
OQ6zDo/CluY5BHM3gmvlQZKsFcWMpy8hdfeerdThHF2uNPGBYbMPW71+PiYRsfw1
nIwIkrj+b9Ot08LCDvODLe747T1k1zE4F106nOHG+gdduyuEJh/kpWvOT1T0SIYZ
OqpH9KoHgK1OEDDjiI6dMzylIXYTpUnKbWM48094wQg8hORuKd3/lnmnB+kQ3hQ4
3KlgFpe+4VxUdMhRVhZ7f2+mvQLVKkUxqDN0fkrojnjgyA/GxFRf5oM1Hc5V3Y0O
TaUOmOkjlIziCvSIUV/mcCuInrcONJAtGUaES41IzedC3A7RDB8rhr6QzNbOiLYf
E5eUwpua9IAUp+9qp/2T26ivL4qHj2jBYjVBIrkMdk1x3CZMOELUaCVsJjiGykjL
ClESPfrWHTrxUpcHzmTRTNH/x5HS9vm8/4EpSijXWacCYYcoCgawRsJn/RB669L+
LgI7sDCdyniYuqQsigsybQosEdJ3xG0E3usr+P936eor57/Nd3leH2DgyjEhb5fw
jjmBSglJLWebbR/BZrtXwUQY/QqJcdZbM5juXj9ljIryBA+d/9C4zpF1zjiUYqr2
HknN4IF5bHpMnviGXjlaJqeKp99wDmVGue+eHpbRB8GJFkQ+Uikbe8WLsiea810h
RuJrmNGtGFkMy8L19Ya3KiX5u2HRP+/wcQdp4Pvdcr5EI3tPWklrYvbXjDjVt6vg
qwG+POvWWDK5wEGBoaN/6WrzNo8q2kmXyNzVAW/nvPWPCyb/mDP4fd51HFNlS6N8
2k4AT1EgEgIkKLbHfp6564rnyXwcLy1Hx5uIuSYaCfU5Ka5brlmk68WgtfdQ79Do
piLBTXzlDMKLo8lHKsr7eTFb3sjr0+sS9VJ9ksjTWWkK1JSJQoYk+M70PSh3TvDF
YfrrQGus/N01vUacHNTDxfGcp9Jb+x6m9sqCIoW0CuE6ZNgB1T4+8B3+nwZmQs7N
LsQdF0SFpkwXsDJy9FG16VKYeQK9827IlOabSzEiMYPPtC6cP16ROug6BH+TwkLR
LCUzb0k78X/iUbWMtZOhZ/csaG14MTwxYje0rPguYZBJt3Uzhw2FsyjJIplsGIGw
6guzNQ/0jLUVN4LUw0FuW+t3ui3ST/8wkB8ciLirf4AuIUyEcbZjonHuSRmzaa5r
h1J4l4vn6NsH3+ttXPdmrg0rx79UgmRdOnrZEpueUXT0HLRY82vbOV1RfYq3zQ9g
sa45Dc5h5IPIhID9HKTECPZqYoTm1JrVOKjACFg2zNbmT2ZmuGJSPT9pZuLjCEUO
BCNbKftVewKm/C9F2LAHWcY5fr2YqzqhRblqPBmO7DKOe+jtQbE/cGyywXSAdlPZ
5EEILb4KHBu9pArIpCcBI9VZav/jNWJhCwGetPrdeurOiM8OXQX3pnxz06gXtrAl
1NO0nrRhaQwYrs811tTf558Cr+qey3ojWi5dwenSa/onW/iTHuF2i1sYsc63aPKD
/GK9Fj07AwizA5moP10gWuQIAuCQxcQqG53LDIxAMcpOdLPyakOfppaRUPHre1bg
MoRIpVf42aoVUYLivOEcYxdqju56UbTVqkcNipLQG5t6FE8/oyYYAC+5AB9Twywr
V2OFtPI4ERZ+ZydlxJ2U8rwzXQ+lH/7B2xjOWVAILDe2AHS/VMvqjGnq1McFFaH3
Yl+ZkP2XtokM+T7bmFYJiHPGEGxYM5rU2qywIzGfDGnnRoOy1jJDXci7DePsdE/g
BCdWP28ZcB95W5apQXGlnVdLqZ07CR+pJswv6P4cSdp4aNId+0pc3bRzGbMwVNCR
+YQguRI6tAtAxYxRf6VBR/VojriiCai1hbTyIE8gokPa4QSMY4DJo59qtY4URsbU
OJhvpI21blI/njFRnhIhtNiXwN5lC9cKS4/NiJDpOFCrOHZcfWA7mRbD7ezQtBfE
dHJC48uDdFTW4wuNlKxjtZIkzbWW5k7WmwAE7e3Q2qEKEbFGGZbJPlE2/YRQ3FwP
UZ8BFp5zTccIF5qRUKEbE//SAycPN2nZ6yln0Oc52PSSdKSXbTLyvz3m0N9TQExl
oOqq5mxKQZAzIXdISr8UwOdRFAG4GPGFBzC1ffQVoyXXT2FOpyx53MdlvxQztERZ
GUkkKQACEYXUgp0xXtKM7qeRgzMYga670x4Nd+RMZomXjtSjqrokASTM84L/ZW8q
D2C6qsOL0nckDZeEyV9+4+xPV9dzSfGWZo6MPE39MtqEUSypd1nq2smofF8xckOW
kOeudV0Q2tqoGZyKt15zDZngPKju1XETtKA8hQY37LIO39VPIqpxMN5qvhqpPbAS
pfUrw3YOzDgdc8wcZmKEl58CVRBbrqIgH4VPx0or/5qDbmxoyHs3mU27jv8z6h93
sYxmzvYqXDOpH4mKue58E03OHEXrm0nX0ipu/uMYkYoIAwbzWtxWDo0MvkO0oz1b
sv85V+B/r9oKfDw9fem3bFD7Hd5UHMKazW0+7YUeUWzGCKHt0kKHAAuxeu6cEYzO
GenvectfhPWbWTTywxgashiXpZBKcXuQOnjpVq5MNT4f8Ga9+o82D7nWybT1t857
lQ6VmRTwEFmFgZG0ISojQW0fWMA6/cTguTZSSQqvlZ+3b0bS+rdO0sp6268mvO17
hvxJM2yIQk4IjB6L6as+5RIJ5soxSLZ2oRZCC4yss1MBLZrStPhXTE9FjjQI2hA0
DtU3WVmZuCJi9cy0jLy9iWoPZsgCO8SrcEEWEQBUv9JuWhMIMmIrM4aUQ5whDGg1
ZceJdzLJGN46ahvvTQL01mdMebEtXwwd5uzFfOw3rJHG7Born2jG1wIOeLmBJha1
NGcJNOfgrQJa8eb2hogz7GMiJ87IbJ69HI+G+OQ16It+YFr+hvc4VDz62QuKqn5n
pX2wBgVdNsC2/C0Ph6mUA0DrtjjraU4AXMavTgvaMFgfNFeisI0iLU7R+qihbDtx
d0XyPr167TLg0/teKLQJqZBZheAd3xZ4Ai9V2+3BZuKayhOrgOnAmamh/ACi1trv
rMF7x8E8CjP20Ryd0gxT9jdRlL/Q7C9043fPBamlBdAT0JvEGwm94mAdMk3tj7kA
jToNm8J3QSa19YARpCwGNOReEODqdtu7LLcQdZHnnO1noHfvImSlY0oYvr0ssE8u
iKmZJ8Sng8AGNaJbRsv5J6yx1xIuWWCBkFQnRp1L/KxovBiros7eJhf7Hgo9Ho9G
NPR99AgnXvGA3JUsVaCEUY3xH5qSRrNDDCvkwbLdLkTw57Ke0D1GgVsvATws7EXZ
36AjjNJxFd0Ij2Dhf13/1APUmNkWfhrOVjR2jf1qvmbs4HJlgjtT4mCny9QnEAGa
f25MTgN9Z8UiwQtdXA+irrN/NmBadKgjLzG3L2oQFbiiA7eG/1FHtLTJBrCLZvWx
HY5GWS8nlTgH/1sg/OKUpGV3w7Xz2CUb42YIwQCFQ3zXOtsHh2E/43w42W8Y8tRg
xwdzd41+3Zt2JpWJi4DOp9m78/NVnMWbedbkAYKAw14HEXN/bNru5IOarGk2tTks
QoO7qznbNcu+S9+KkzTgd4SJ8kVuXwJVB1FxsO2Hq54j3ZWbpyId/KSRKbMdvYAq
PkABDJUJXryvdhrP80KET8ZQ8abs2o3sv2JwIlfPO9Dsm/JhhRyW+oo87v5Fh9xy
wjGDWsqdip9jioVzG2W0Cvko/oyAF0G1b5qYU/cwY3an1qV53XLZf38jIMaTiMsp
WQtL+G+PBk1J4gH9M7EgxKWhZsoPAnM5lBRmMKe8oJK5MdNpbhwEW/mBkTDrG0ZB
eAjigbV7I3Ih7e4PFPVLSnh47Ca8vptTTbZRl/TBDXSJBFobQgqMYcCNLqEbMkOd
pIVwB7o6rctxzLU+7IYOl0IngxSxm4IC5FWE6iVDjptrUAWEwC5+XiEqMbBkzqZl
SR0JQCRC36JxHuctOSIPE+FlNHdTlGCe/rTveMFwblmhcE4eL6LZukeb2jUiNeuf
kM2WgpnR978Q9tZrY/RbbSDtZW537nS26oX8VB0sVvHPO3ZVejPQhjhE0ltEAoU6
nKjiCzugDgKHRjM3ge0RY4nF8yWn1BBLnnYsAzMngjc7DJT7T3VYis+eMxK4aNr6
usVvjzgTu4lajCTERr9qr9zSe5Eme7SUy3tUSJbRINWpWkcesj/HPb5uF6CXlrD6
iMKd0+ekaWf+aRnacRZFt+GCHtnTQuK2ucMiKFUs6JOjawqJC2kgz1DpiALER5VM
jtdCHf7YuCr8w/LQGMaQP9z5xvlQTjUOuN8GR3e73J5zFwNF05YonMQPT9w+3PW7
8eG1MfQwbziJzYpDkbje0GjaFTf7UXJwvg0/YgSYKhb1BOduC/HnwECTEehpxVDl
hh71gvK6iB5HYeJ83lxDix3oCHtlzuB6ZS8ufG1yUNMZKflKCIi9wr2pw5lnhwvB
EQydAJvI+hILTceMW0zIO16ACTifpDSl15rQt4eJ3ocHfeMkvpPSogi5s+hsd6mw
HILiYW4aacqruFXYSmeORwjW/KLcgsGzXDDh9ySpHoQ1J0R/LlCitkuzw+Y22CDF
nLXPZvAd16NJdNzOA4M/kJ/2CKzy5Qb21WJmu/XTh5fKlkMSYxyUbPVMEIBQXWa8
GbxZ/Vv9M0nGp5tso2e64HoVGuuxcDsPKd9wqvBL7JfKRMLfBKl1kDvYHU/N2s7M
Jw1x5odNY0JH2R22hE9T7CPp1Jdj0fJAk891HTqdYh8EPPJw+vCIbAgZhQ/0W/T/
jq9e3TR5m1wMyiJNy0C1hXBsK8Jo3CqV8HxArwRstpBe+sXQ8er1YpuVLq2sNpqh
gHambjF4tMXLAGKQCRtLU50rt9Dv2l4DvIgddQx1JYgjWbFT4yXEYEICUZh+B5uC
r3jtFUsDv6yN+HmQXi+e/+urnBC3zhRsZTmJGO/M5IntCctzgKeqUJ5HI3GhoBv+
zUS/9OhOyB52b9DixATSWQlFcEGjas9mJQgtovxuUNlpoB+AALpsFp5kt8niZgNT
STqqMwFXbNnjasNUJ48nnWNDuupkmknSVL9tWEKUxlJ1FK0bZzy4TmmgQ/pz7VMZ
L3C42zM63CfhKjWZaqoh6mKQ5GUqG5B7xagmVpwctTRdv6YRMfOTwHIwxdafyrLy
r0vaRclGh3GhbFprkY2MQZwGujgiBUFqpyvJ+lDiygzwzUqxjIvx2CXSY55ybrqI
5sDmVN/IXUR+cwH6YQixfYKRcxjIC41w/JjhwDNpis4w2nb81ti7Zg0zmUVuNIC0
G9714Fyw8+0IGrFVx9BsfoQkX3s4XFaUMf9iPMvc8odSZ7vZTHg5GhnORRtBUX9V
7UzK5bAiEIemze3BM/xttDvPWkJJFdkKGPPb9yr30OgVTPrg2Vm2oKCIIe6qPJW8
Od0EkIqs6at1kCBSC/15Vax9By4VUvddhtMouIXOp1P7gL0NKwVolXt8gbX9utKL
CkrkBY/QdMhuE/I/N+fGNf2CsjaeVwPr0ZXFcM7NHQrJ7uAmpezD4Vr06D229XNu
la2z4zTCaHRBn2mOZQAmtUbo/8rtkprATuxgfVzwj92rkGf3lyGf5sbcpnYaOsBg
PTlTr6Wuyd8FWRBIus5tcQFqsRfazKKaoI0wd2xLCwUVj+WHckWv8AMlBF4oVtxk
++p/k9z3BXyP5/oHzXemS+RllfW50mu/AW614frzA8mQra3R7rz7vt4tV7TVBgGE
iL/TSjC10FRqCAeVDWAESYTNS60520Z84xR5AH5oqP+15nuLhLZ9GBqsNRroMRo4
FVMg8Hx4e5AbjbUleg1VwIrIPSHqFnSOeNiw66qWtgE5h0tMx5q4JR8cJVpjiFpN
gR3OOrn6oPXAaDrRRRKU5iyKc3SVkqSyLJdkWuD9NJ8hvEktdZV8GWTfDQUi4KRK
vrjT7eiMCc205WExxw7naVj6lhswGhkiuinEuph5H3eJLeOx2J/QZFynmXiI6ENt
C3YldKQTeGgMOoB9oqGWNoZPyyy58APTZ4FHoZEpcGhnywxszY2exl/LyuhHfQmc
GL4IbjEVu8onDd7+m8DZfK8O6IeUGNkNxq+DTPlRUZSdmyQRAIWOxjbqoyzIMd0O
D886R3pQ/KyIUygADcz9/9Gowja+Olsl35gxTluW9MOlZ/VqvXeAjFkqpDWBUiwt
HxhpqZJDyyNDMdIQX82XD3Fcm9YviGroU1MDWxMcZrdMWv5FNlGps12QxQOYyGP7
BtkKQXx4XVcgXyhBTQmXKBXm1QM/qFAB0lmQBpo6n47VoTSUvkYuXXWfGisAhodH
gDPiJeg9YEVVUOmvPBKZA1hHts3dYf2fWE+gwncrN8lI7heYugMsTuWIDjSzr7G3
tMeVn+8Ck7vg+9dyoVpq5Lh8+0UjknJ7SN3PR9zSyBOeAgboT9ttQ+pUHXLFIytd
a9MvWRmJHKrfljxdzesteKa2IH8m+TbAd7/DwYUraIXiUqo6rFZ660WqsjfyUXZ4
Q/bxQFCR0E2tC5gqcVRYb4jJYKM2DB9XQ1SuIrD1SFrS/3wYM2uzZUahPP6SoBAH
ShNC5wRavq2zot6PVpNur0WJrTIPiqV0IJ9QHMGXKafov1kLJBaYYa6hoyqkDCIe
UP0G4AsQJgR+R/YisrMMfB4jG8mgHje0CtTksKoHPLgioG9u3QzdSCoGl7F4fajj
oscdUedf1Of9Eazm1lnc5Sax1gAcCFCm+hMC045LRtrLiKdKIpq32avbv+RdBz/F
q7rWeX/j2ukQ6YtuaKjd0O8WTgQJ69gq/C8zEIz7F7AjSf/i1oA9rD0NLfWzX1zz
ra3yAMaKaO8KJKLSvKSoHWqjLqq6eESnZo5tjGSQvObSYS4JT5VRP/bqB37ZP9uE
GT6DvGyvZ7DeUXLLbNzaYLyOOo0mPTxlF4JQZQJB77EXE/tJnQgYMnNyLQKMkKJB
zJYTsVEvoEqfLWrK4gAr4+hcjnGBqufhmrDk1F0Uvn3afopOGFj5U47JX+hrJdJi
JP6uUlbqau4X8RtHK9dSX2OHbXwZmB8aOsKvEEAG3NGc6dW0uO8g8yz5i0EkdOQn
feKiMFPRAmxLVfzW4Ai013qamC0Yp8JkSxGX85cfIyG2/WZlKseKJrD8yIdUl/08
sxZ1fjPIcDXZoNS0hNohyo7QdyN3Us5wplBeEt7RzsBjE4jw12RguqhdcW86Mpdr
/bOT31OVzl7hzVSn9Bo8mDqf9aqY+M7YJB0kapR5OEDx7JVDQIWlbFc57kNO6XPF
G6zdoPHfCct3P4XHKKt3W4x/Sgfl6u0/Q50psHciZatctib3vYp+TT7qxTppXzkn
T0VHO7iWr424wy4AaerIpX5Lygtb4Hufk5HGvJK7nPwh7n5eCG71x1CLx8sO19Bc
cLZkOY8KkvHeD1ElE4iWdYN9BBWkYnEvxYDhWd0S6dAZ+iOMVHiU6CV60eIaJ4LC
QnuknIOrTYIrdVnnMY3uCHM0Qk1ecYK0o7OoLC1LB01sxxohOG5XhTX+Rl3wBoYy
3Wib3VMYvdoLEEjzjTRVdLjA8EqK5+N+1zTDdXbL0RVeshK10r8W1ypBFRabtNKB
8aUiiSbB8sbwF8KZOIlPa/GQhk2G5SP4SDfaKByUB3A0fLf5Ndt+JVT62+zyYwuL
b4kPEbACIDVcoWn4lwBXI0xeKCGz1ihDziXDFrvf8by/zddkPg6v8z7qwTBOSPfJ
ePgv571IVJh5tgY18kGU+swvoFfy4dr9gt6JOAym3ytNu5SxF8RGvx+yO+Rlmu9l
/azYK3iIRN7IVVOTaIDhZw6yZ4T5bj7jCQu7QHJMntXyxpF5+CfNAmnK+PCGW4bB
nVmqUl/sr/Fc/jLW9pjjr3C/vgZkhfTtc6sndIZA/5ksC/Bo50v+0meX34UetSvd
kH61e2koA6Bp9nNxPtwYcJUH5IoWxfWPJLEvAn8JKUE/gwSKpUoTsjbXdcx5R2J/
M3abY7HgnrXvyAeQv1Cm1MYyB43Si/snNpr+o/UE7vi7AX5LIi6H0iKb+cX9Kjz5
xP1Y9o5T0r1lT8KWWCFfIo9vLBLMOhQHDFsXzgywyTJmgmdL34q4kiJVJhjcVmNf
tgCVGzN6L2bl+nxUSSpRQLyxO751SrkPyLFyB93hL8Jo0vHeuV/31pDrPaY+BfWa
I+B9N6MHSa4sLicPn6lqYpij13+n/YamQ5nShUKLBmkklSKaeCdl2dE/7t2mE7lF
747cNhFSLh6W3U5mBoZi6CwxKBfDm+62/KpfNkmU23tZ7o9cNR4rNayu3Fg/KelW
pPZllXcnMC09+cOnojfQB62qDviL04TVrPNJbLLiY/gOLx9ge4SInwO6FvaXQTs2
KjMaRvPRSbrz2mXHnHTgBXv2QcI7lnmjSzH2WqnNqJvN1ZIOyXFURkHpPuOAEK9p
j2/PG7uhXk5nrGraDGybPGdESYFgs1yONAff2LFFOVfpoZNYyMnh2+rXjZxGbWVn
27AQq+tDG6d8XeY5OGZaXT+07CLU/SFQ1FnmMtGtjYCkUb/bYZZAkdPDGjFAZZZv
nWwWjcMhjqSGlRLp2o/VbS1LCPMfq+keHM2baI4UusBclH95HYJjgSJl/dlpv/3+
XmduSDNRby8TMkn0x0bR3+rwk8yTgGiCQ5rUcPjhe2NPgDtFLIsTDdxh6fiUZ0yQ
+UuTPcwR/RdRtF3d4wLA5XIiB47DWxe8J4GO5QhHSx0QTLbr7ZFIDz8aR4htcglH
C9hwpel2mgcqSM9c/Ce3ccrlb4wJaJs8jICuZ/cKGqGsur1eQNyw9mQs3kSvp3PE
QTfVeyj4E/r/U5MglnQE0xU+78hNoX0AkeVPgOEysgQ3GWXwI76ND5fKkdR05woM
B0WssmH9W6E8JMAAnk2UriXTqoxF06TGTxQaNexOtITCanNqdvH0vbAKec+EbAdg
QbSDXIfInwXObGDHWGasEFIjEFizPPjNzFbs+t9ybUho2/UZe7PT6uFShDeZcnfv
3Dl0ZdwEHMZpNjtYTnTJ76EZ7pW9fVUw1qiW/ATuzNUAZHoxaTdr6B3ffzkLP8JF
p3HfLt3Z2Tsd08mOUopM96rLk0/Gh9tEslC1ERTeuzFNM6jc8PLh6PJ3mUEop2eg
GCprcG+yicm9p4Aj++MJoRyHlgxkpguUxwwvNNytw2JNXhuecl2LScdUl2gXJKyH
/JGoAngl5T6JNU0vzAhyHxKOWvX50f4ZXyHoy82z7kHNpa7itWHQwJ6eFlTXkQfh
0uYzg/N1it2iToXb+Ze9T8kBAe0n91hcMvXBtC/6xMnI7rOFflmJiyiXLHosHsX3
7wf8nS+6fvRUdnoaFs32Imh4b9UKnLgEHM84Xa1hoEHj7tpUrfKvsj2qYXqoWQ3e
BPFVDiLdfVR9Bkb8MC3SnKgekRPaN+ZXdZKP/qWwJgEYvhrYMBFjZbpqF8rtdMHB
ormVrOJ66TAwI9SrvwzHDNvIsnJWcqqQ92tVDa6NOyNhBlc4NAkuxwtGTLD2crOr
mp7A4je/4S9A6FB7wodFXrkI0If7TdgVjTkV3Ll9e7C9N0+k3NIOfd57sJQcKbew
8EvN/DEp1AxrCoDDlGw0HbGWhpWRR5LO4Dn8AZ9Jy/33igR8xM9NQMpTTT4bR5rX
ZyJPlhRoC6rmP+lnOKmW8oJckDjFvu2AvhU9g/1f1F8z6rzKH28lzg9yr2jt5UPL
fQvddxs8ZtQkBDKh6cAgdfMgWPbZz+X2oD5XzDZRVwB0JJillGJwwlae+sXQlik+
UD0pqbZRq720TN27yU582S7Q7LcI8JkM8JvVw5hfxSgAp5XXI4JLLUUwRcmXWBeB
9zEOBQlFd6vXhrqT8RZ2F9+YIWS3y20fRmizEcqZpTVjYt1mdKiJ4MtjRx5VpaSp
IDf4IzUJOI+9TV4NIZgx4ssA3T1lV06NlpI084M6k6rcuFtT6ZEHdtatWVO6xLbx
s3cLQYjc6SL+IpCKOmVSJk0zC0ykYA0C7t1SzxcduULst1fZItjUvIOK9E3T/zgr
71hjt+/8QvKfARzHQQPssj9D/XPTzzRlGZWefMXh0+XTuNnYKID73Hd6ExdTReSN
u1YJaEmH8j8aQF/2oZICONNKaTpJkjrfJgifpEuw59sSy7FfCSZCsD3oZLA8rcQe
mK9GGyKTMLQn1AIMwqSCGhu8N2A3rrPA6DGgYW8gqXBoa7Ad26cyRwvTuhWd1+mq
5cBx5DKj+55Tng8Ic1S0a3o4TbQPnATTTR8kiNAxleForJ+XDSQmennRb/4zJd4Q
FJbWYg8tqtDGZfpCK0rPqPPy7ii5o8gphG1V8iF7Yurqvuih6tpfdrAxNGiPUfik
0HWR41ZlLsievZTJ5ga6RRwysFt+TBo4uzQKXmStxUb1EdDgk57Ja1fSW5ew5zIx
kJotT1qFNrDVkZPr3uwMVl5nGJKPIguKT82sNLlbyVL1qewuBawppoWtPG99MPLH
qH+VSJsR3zACXxvxZyPq/Em1El2illkxhEKK+sbwXKaGm67M+Bzs3P2YCOeZkui9
+61KUkn4DhDgr6ujq+lG27SXGGFRVP4IOx34d0IYK6QemvDX8c5/6lhQIIgiambR
q7rJt9ozJxLXMrOSun5ml4VlYCvRBckZiPikJr4AZygJvnvPPPrCuz2czAXBRdBM
Z0q7NTYQU0Ha38NoUCxwPQuC7kUvbF7vJBp4OZbfCf7KXCRnd7cSR+4ODOlLrrYk
shYVRteHSIqbTHyGV19bTW+QV0wn8Ue4qa7AfcnimQceLwMBMxgqmsbPhNoth5pb
YqXNFxK8swjnIZzM8keT8zwqRyUGej8p2a3igeR568hYo210lagLWxQ7u5xHndR6
pn6yhqKkFOsawHwA4zu+5ntDuwfhqZJa03VsjIeNWxf4gcylZUjGS0EexenBRVCC
SmyzDxtcafbb8jnh2fpqJHZD6nCuHW/GR541kJRLUUN3iDcoitwk9riYGOVvjF2W
xx7B7vgmgH3rhgJcrO1SvVp16yW/cXdyRO51DpoV1WKLaUIsu6DloRZ4ujSNdS9A
RNMbL4lIF9+6M/PENS3RmMNAITzOtrhHikz2wwEDvfiIMCLZDILdUI9N6D+wtIW4
6Ga08Wu3jaDyop6nOSJ8tJukvi6in9PL8Ywmkv1LK5z7tk/Dxuph4lNgYC+CVdKU
tHKXlwk27mZ0aMET0uRe03YJEbG+WDiKYQoKGaUegBeHAb2ja+Afrls1Mn+W5d07
/EZUpxawKBQD2cZYQXifc+GGqm3qldXFtl6Oe1IGdKd+h5wimyYXwr9MsDI/MOQr
1T27uBfWYcCczL+uDcwe56syvjROjTVrxDkticyhrYpR/iM2prV6bb8iZswz8Qft
cgGRMbRlghvp9dlgTwzx+Uhhxo9hWizvs4TJeU6b4uKuzpWmI+y9EnH6erCeGmav
Q1ESO1xwCnHZAvqV++4Su3p0n13g0A4rYnitMJlmHRhBPv7iQlLKsaV4q1gKpyEP
FgEmmyEPjcYSot5RDhod2oUi8qnoVCiPMn7V9gqrWyPnvJ+gYP+SaTs7Yv9YWWyf
F7VTWAUIT0Ubmsw9p8+RcvsEriiX1DFKymWboGawyMwrT5IWlXbR+XwszlPM6uc7
7vqTiCk856lW9J2eGeapADe5NdmnherDE0mHwHkpClGMKa+U9ScZqWkf++z2esGC
CDI1x0xA4+km7UrCc8/6AVleorXwjNUs7jPIPlGEBrl9YMgLlhrt2sDYWhw//zna
YUPH+9VPNwNfsyhtrm9YHLmHNqYk4MROTWhNIJ0ytq+7c2aNJGYhKRvaHplU9yx0
sNufTXifJCdlJdKn8V0pNnsKcgQPrmyhpYuVlOMLPzjk3bcgKOoNfXCO2rcPao7P
hWXr//KA4l4+bhnqML8WssrzbsCDvRMJyL24UaRF6qj19rmXcdLYemBM1Xylho/S
t+h4XJ46EVyZHTQvpn8jf/HGFQ/dIVywZ4Fuje4lS30EVB6IOJHDYz7We3AdLLDK
L10yMz3ng4RrAU2BLhTm4fTWmPZvOGT36+UsjL8wnN0hNB12li1Iw2HyoSdSXEUw
+O59G6D5rJTKwacmXUfhpFrMe/gbbSy+09lXn3i09AvliGO/BCo8rvzUOaJ+ibBs
6bArT+9i/joAy10UZdxVVddxwZMsiE32nxaPzvq1Uwkfa0F5MsxYFm+YFDjsrIZT
ogBx7nCtg8hbu3HIPf0RfzmDpClW5zDdmV02fWPVY5CKlAm4fhTC7ua1PeRln5RT
RPEhRzlYZO0NPba6DMj2PGGsE7hZ+3wziHTjIjLGc2PGloqzl/K5SICdgAg+1nFN
FHFEUF/Ez+vsyGrUybq7MieBCy6vRPJq1vPzP9/0Mp0gJd3LClK+dx2xlDjc9zYp
axgNRdk3tu1RN9R5Tt+TaumBCMC7r+rCf+KeaCFGIq9XYiH/2zkQohq3BmpPqIFt
WcF365eCmuErc4+XPwK2rOljibcv7ATj440u3jNvxJNaVm5SgfFLHyTxizEKWecq
vGjnXgwf82zbOyBQQzr8AwXj3W0sKSwo0riFHH2PmX7gfpP6sNGRGToUzpAQ1UJ8
kVXOGFm1fYAUUZVLSVJtRD1od17TSvxJ3hAYGmJaBA4GcjPcbvilM+s1I65qUu0y
o3w9ZtLgGax/Ne64K2gsxcE9PJ5gMe1nYiE57PvsquzxeR5kSmllV3Y58EXLFrjK
CD5gfhpAp+gnEsrf1WwJtss4UvcovxKIqzsE+QKqP3PMF7TslLiFzPC4vNb+lmSx
gkc35WCP1iZxOjKtIw9I5FRyD9w/ZW2QWkNv0BdUu3cjdptoEUR5xOKaLfqnGnuN
iwJOyj4wZPESGwulpPlHhzuy5tbFW8mCy0c2K6oKuXHzjRqad8p3xuOgdGGdlfXu
rYdEt2PQqxlJwL5ajKESQfmj7mF2QAkINtawAYLUQYQliQuSB3ZfNgTJElKJCnPh
uybOEzsngHBX5CPGdU+dPqJ9Tvy+S7IvjRnIpcXW0RJo/nmn5zCn8h4wbi+kHmRx
kyAsDwvvI4rl53LJhaB7aj/Z3ig95OSJTO+3TggWrFGMIvJ/+rxAEa4DmcPMdpTq
OU2/Jv5VrH2kMOk+Cl13gqlt2EtZFS0p4dfjHnzJVQaVkJv/GQ3GZNPOHsFgA9Ey
zKmeAYz2YRYM6RIR9MvUcN0NnXayobGUTlNcvNjq+XUcvKL9eVvOW3uiGvRYxupy
ldChHHXj4AeNgbcvEz77rmjKdhntIN4pWik65TqBEPoNc36RrADLU9pUzWC4yTkJ
QPxJ2h4iMoep8o/ptqYfTh6yFiw/IvNaEa+zMnhvy+0dEWbx/BPc4tJ0mhqw/pMd
x4COXynSzVgELg7Hklz5MLOs2QqofVRU9IHiUdHlM9nKbtqL6UJ7rtMKZtPDae2V
DjSJCSB/OL/HeiUvFLdHutiRn9PUfk8QL1d7s3boXjISnwoCVxmT8NF4DFFxi4qv
tas03bwLgHeRpDyXfbCxiVCHJ6JpwPldMx7mqqxciCtgJfvzMxt0XuMbrk0Tr/T2
2Vw1oZtASOT1+fPlSgweeXZ4uGVF5AAAv0R2S6ScsAxSqGn6qIWTwhIcz2DGWSY/
jS+09iXo6vNalwMzPAB04fFKZMNOKLCjr7Q6UltsAvStsRtCLTpI8fABuuMa1UvG
u+44E5lpGzye4sRUf89gY9xXPUs+XVvA0SLf6LnsVKrObk9s9pIbhZz66SXg9YNG
PHaU88Qfz3rJohJJVm0QnBNECQQyVIAfQ/8prEmT9CE8+pGYlkMPgqDThUTpwj+Z
AipST/cilYcG6zG95u+4sbwWRc1ys2nnUVVxi6QIwhxxpUMKbA+Afbt7tNXXy7Sh
ODawGLBK0VTUYOTs9hCYvh9u6H63I9+K65U4SuZflC1cnEU2VqK2yWizOuwwvhnA
+zcXid14L1ReKL+x1De+tTBW6sS/1ltXIldYrRh34RZoL4GkIG2vaVrBWEA762T5
k6cOsygypOfw7xq2tpSgPvgaYBhTuybWCkPYBAMPZ0ZCYYlhVV+Rr7JAUz+PAqUu
0RgCav1332Woju5aqXI7aflkyBcmvz2b261uRY4Mmy0Ctl1NQxxtE70CPjBmCqXA
MYzZC7ryDs5y9cu3sJVdbQNGaKZTYcEtiAmz0vyNTnx7c6Q50Po3L7fx7VvojIsY
ehMBqCl9yDlNjyMI0q2rNoV9n5neGV/TO7GNUtP/0xhxRMHigk10YJbbPpX/I0Qt
B6H2SyMKlgi/zwt4esgomZpuBXwldIVoYGgkDF6CcX3TUYnVbQOuGDIHp4ow/AwR
8B7pp44O2CCLPnZ+7L0nCYUhRqRypxGdU50THq6UnBS1jeZpz+Vrf92zfILYWmlX
XOpHM3KcgjdlV+5JlUHYVpK5stX2Aj4yuf+9zIpBsFk9mcrJwDCtKyOKC0jJ2CMT
LAmqs1yl8Ou0bTfJ7xxMKN3aqNL2cGhZuKI9Z00Q5R4gP6ImEhIdNCeYD/ZCeXj0
1lmPpmltrq+2AqOzrVZwGk3MVcceAa3iLvuo4EFLOrDbvLJ4ZRjtsbNRfow77MSr
zBF015gfwjCPs15eTKb7tDLiorbtOICc/5veGj5iZfhOJk3Qzrf7gBeqKml03UlQ
oyXgUD7SzKQ6UYTWgqiLqlN1mzPmqJ8Z6bu7mu2Uh00ZiK4emZgsTOFWJxr2MUYS
+85gVnuCSix9DFkymyxSh8l+qrQQ7l+vePFQyx0H0wR5JNxq+tNTlZMk4YqbVYdV
RRdCLdwdVJuuMphu5Fy6ZKwmCZQxe33bk48zO9Oz9t/fTDmNFmy3cm2zicCIkXPS
bDDCAy0ATYxqFo911hqTZL1ku+qeNObqTGfqnxfw2xI4uedxX225DLCpqNe3frKK
AaU1Cvw8lJ9HSEcJ0EFrK84ql9NYKVWfE6/bvwNvAvTULbKyueWH0LqoNTJibEp1
IhPpHCiD4vJnOx30tPegq2BE9pS1pCHNe/Attf9NVLhb1iytqyUX74iojAqjp32K
1lHKX1INUPP6wpZGAiEq4zh6Jfncc2lyWDsdJp+zzePKpE8MUu2cNLT+k2OJFOnO
TAX29E1bGtK6By/Vp9AhW+DyPSKDzcsq0BwSZCvS0fVQeaFp7+8ifwdInc4xBHQL
dJTFqy65k1z5xhy1v88pSZJ7FwAswmeZSIKR2WALdbkuV60N69XcDTq7TFjdLcuh
y3ErbHE1S8QwtrOIq6gFyWSzOhwgb/4UqLLz3p3HpxjVAmD2uqI39kVd378pKhGR
vo3MNGXO2Vil3hK3KXdix/4mHOisCZ1wpy6TP+e1mfALTJPcNxSTuEqysQY9xYf0
FAo0RLHWC3+HMmIdQPQuGVKh9O8ps9scfakASy3wRF4sU+8i/SBnBzSpvmYFOc4Y
RsnFW7LrPeM5fabNuSQl8+ra7Bn7Z6X2qpt+VHvAaIgQu1yN0HNLKHsPkxKbXQYs
HCntuYAg0YM2+sXlHX+MECC2oD+KcPuB7o+KS6X1/y0wLYSfHJ9vOvIwtTGTs7iR
SyXR2lxoPFf4ouSn3zRNnNii9WDUuNv9nkTsoSLYwQDzHA44RuhFtxur70JfEx+B
o/UkNOn6i+ohcWdLe3HbukAWBAxVzvB/BQleshwX8opx68VmnLQfsKEUXaDcWEc0
jtIgkiSrKcpdiNj/xQWdsOCnfp0089Em8ClWWTN7p70aQdS6Iwuy/VwbEPOe4J7S
fJy4yC6UrBVBYBCrcw9HyXgwZIW3vMjfRM8ESpwZ/ohsAVmzLpJtw+Au4gWBRltW
vyFonxgb9SUcPcGdwfXuVaNeW2vmnU2/62axlx1nIl7KKVgQQyi7mWsbdyDNdDXm
GM7lUswYbWz11EVzOTceCh5tjfeRQmjkTO3TRhTf2PtcjdwH9I489S88Koe3tRzz
fIth3+U7bTGzhmKh8IOMeElC2u5Xy/6W016hWrxOlixeRFl70AHNHWs+DnHVEjjm
XrBP3X4D7xkLm2SMXqS7bkUGcv97M9xYraa0S4AzjtKc/MHj9y5r3pqFRVSs1uxZ
Y0PF6NodGPGonHcN/2KTtys+pThkoyQMiA5g5BIQsnU4OuwjGvNgCRzWZZJJ/O1/
mxnsqAHBasgBeycEQ4ndnvvoAGeGJKnJ5mDkVqBaMSVR5aYSpMnpuCU+GhmRa1xU
DqLUK+nnaqAP6viOyqShrRTlLI/c8beldk+iiS3Pw9WYWfLMXiOQVS0aeOJxcrEl
Gvhyo3bkL7wTHyF52RN94Nv7RNJIx2dcgyt5bdZmHeytFZwihDuCcYAZe/jfKLzP
GIVDRbu+XjdTlrBWUGyMfJPegbelR2LKZvW4S5ekTRx6lljJcf8R10OFPdt86yfa
eOflKxgBqE1edAAtZrqWkPGl2LmBc7Upmgv7RGdE/xQNT3cohfD3ncsw39PPrzUH
hXY34l1ZNV74dHU+2uX7d/mriO8onv28qJig+WbHGpQ6Bg8rJJap9OgmQtdpg7uj
W4cFssRh5OTjw3Wxtb6PwbKqYxX0rLX5Tk9W2+KjP9/vnscI8lYmyWr+mNiy9xHS
Ug6q+mwyPKHyGKjedPVuEckpU0QueaAb+22FbfxuVT6RCGQMmQY6cVnE2MyAnHgt
ERef/CB4le5lj6gv64Q232sIFFEglSzh09UmKNeoHnmDOH3e/INxBqrjtk+qMLRC
qhEGY9IwA1CIzuMWZPh1URomH6/QPLYl6uxtxVI0LDiYbKW1u6jwN6UcLcmNlOO1
KcW1gTvUIGLqbdfH0zDwENJIohlgunG6pmwoYuXgdVK5h6/+8iq+g3IX48Oyeqaf
/H4IT12xUjO7mJxU7o+EKAzkyKIr6MFSu/ihGSieYdChvFAUg29TUqlgaB9NJ6wG
oflTH3zB2aeWJ5oKAUkAqbQUUeYa1vTNecw7zxFk2Y4RqOMWE2MUOr5aqOTCkcgn
eXAItk1WgpJ4jXPdy72sl/PMxnZlkk9HrB/tKmTg+MsJgFcYscm6TwyJdSRFnE35
dgmxA8oXADv3pzbfJJhuz8ZatJaKLPU15PaU/DYlb0HJEezclZ+v+uYiIIyQ66vH
fCMaMipAbqnzZQu3snF7qXw93SY3QKaEBClI07cGfnfIbAxJ9YIY1hVihivXdX8W
x6+DNz9MCBAdr/vc7q+SOJXTI/TgfLwrRffDWSq9o7zSEihbFDOysWN/Wzx7b2DH
zhxF7yy3+1cpKQ4Api2WOC6WDjZ3CdnfB58TdhfQ4ghYGn78DIAD/W89eZRSnRhq
cl2U6lMIzZhSEfbgflu97Jg2KkksEZZSCexfFK8jR0LSitBUOzcuLVPwpa/OdStM
fyCXP1XSbw4TB8pgOG9APXubvdW72Fmeh69lggVDtkJubSg8Cs+bh3f/Tk/ApvWZ
WfqSqwq5woex8WW6W9AYOnrbdnlBJj6pgDKdCof9HGIP9zCyTAbX+kW1bmicgfqD
n977xol9nZEXdRtpGlUKVTUdo1tRHJMbmFPHnAHbB9Vsf+48vWt1dUkigQjpQHAK
83VSNi0micYlqOYuXElykNp4QntnlBY1F7PzyrAbFOkU11tROjTwqjPzIiuVGO7v
5sOEweWr//9xlgjegT9O8XnwDkOJIxYhVzXO/U8fXXXfhzQ1tWk4g0r/JY7AW8pH
oWaWWUxgDTnFt2MgrgMFDzJWAzvOr8xsrbJ5NociRmZbNZa2B5THNb6hhZAN6PTP
bTgnYbhGBwr2DVmN9yHHxUv3bvqPU7GBEXQGhZxY+HHc6QOqbiPO4foPQYYrvzQv
KTZCqJKItCMkPNqO8QErTjUMkY0OwdSSEfP3DokVbzwHnjf3tOkxIo/qLJg9Ia7W
AgKTX44dZm5325t62kl64AqtjnleRYtikcfpj3hdI4BCUf3EF4HtUd7u9Qk7hlqh
ubom96R9sTtptl5hrKAIFpAPsJr/kkPGW8+glJCnHySJEuYJbYyXsJ8bhA9s8cal
H3CK+QicOH9k5a85MhF1qPHaKSfP2FM79PDXxVcX4KCMYSJ27NxOZ3tHHWTAwALs
Z7/rZv9uYpOh9+NjQmBdYBaOw5KyktaqPHYdmqxAT1MgO//hSj9sBW+Bf5a76+8e
USL4hoyOLj/surXfkgelCmnVlDOJc/JcZajWjgOcWJddUJA7FwJGoPu/xyGcsPaN
BXwxZWH2hgt1C+m/bvY9ehO5tzRrQUgysdBsWYq3Wzu1k72sjouC0XAzKdWmGE6K
VufuKD1yKV0Ma4XM2E6nNDk9S+NNfu4SIPJyxnimDYYXKRFFNNBMXziha6dvZ/5g
pDFbSKBJpCrv1m0q1n4/0+WxQW28z91J6Yv30NkcaNCy9mRr7O2dQ9iC5LQ4vVy8
YKSFkopRjaAnsBrfzYSzkJMqchqnqPuXVgBuoQFrgrYnm6SXuJ9wt6MJqGqQcVMR
J6XQt4gDyCtdm2uIAviPalVpUJH3ou7eOUpNfzMSLePUDLNsuC7yL0WM/LtZKCSJ
7cGgm4V+DBB01u59eW/WqbCYc80cP2yMxea1hHQ+ia+S5tWVOU5EtWXOv3CRs/Rc
htQ42rYNdPVczuFVf4aeNYWD5Eq1AfwGJdR7ErF4U0PfEppPLcp436NlsHFXzXot
KihGOz1BmzWKD3QYBTBAX9nUIHqgwm1p4J9XqrAcJPnYchDnBb1H/dRl5gSL/axb
Y81pJsNVoWDLm/UbL6OVe709iY2yZvGnTl25hKkXR5RRoZjEvs76t6eFcbbdaFoC
fE5cohC+yeYlpKBNBUkKOUURWWLZDhV8NW5PKkj25cb0W+l4VvrqntX8MquiRn7o
hkA6QzFkTOTLV+dp13jKEI+eIi63AAcYoN867sQ563TqTsUuKkVmjhM3zInoT7Ih
eGkC4MG66LvoZ5RdqzMomnkTVTW5c+AVO2Whu/dY9E3RlcwWhf6K7Pr+QJJMXa9a
BtpewL+LpNmLQBv6SoEfdAsUpxI0ycI2V26KOlbLeJ+YEDbSpb7Q/sbGh9eSyYaa
RKPNrFbEI1ee/4arosKjnACARDw19Ad7yQfSpLaWV4Qol31u9RewP+SywSsA70yQ
tC01cY/8eiTUZQo2O8KB9FlGk6grTzPJns+MgLeG7R7XcoeyIXmZefp47P4g++if
8u2RR/55tpkp+HylfpYoihYTScb/35JywGVG4Yw6kTzzwI3wVjCQbOZTKXMfpalb
goZeBglk2c4OmmlqKpcMeljKP3BxrvJKmcwuakI2kbaYmrmDkks1qYSu5uvQEpcF
Dd1+bxYhyrJHfSsaOVm4NWeK2ycjUSsQavU+/t+qGUsxkBGZlFo5VWM50bXoiyBX
80pu6Pyr6iLR7ORf6egAMLg0rrhBTlxEHWAyJbmzcx53Pz+G9sQ8qIkrK46Cuju7
XMKYbPVVLuTfplFpdvYcF7qYjzq+Qpwv4ZyjRCjJ2Ufw7+DkABPkH9tEb9uVOXQT
jfHCE6MrHliwSDnyyUT6fA0SXUh1Qkm9gIuncugA+Ymhmhe5oVJAwXSRJHnTk3h4
nzddb1gLxC5wsdOG8syblITZiE8PKLYmH+/EuksIN7sbuioafIBPJ1tqig4D8rhB
ecRXLX7Kqxi/tFQntPFqvIpYYegnInnUGxR/EdTOCsxU046zVftxaYiSaNfGLW4v
SboQ6+fb+29puSQqp4SKVwV1h0IIJWYCxhLpO7e2eOQAdMpoRb344jb2ZYz2llGg
nlCKEIeEOB1TKlx9UiS5QidSbBRj2JQtDaDcut2ei2kb0hK8wkJI/ayIQVOm+H1/
djgS9onIOIy6oEynHKR4DBboA8GAFfZNf220YCBbyyrj3ex6ANxP9xJLS53WoB9t
W/prFo5WSX9OIrZahNpGK112FujA0B2SsNTZMcqRZym84xO7djHrstSdICFKANCl
+6xYjSGexMCOkTPaJg9waEq6LLBbgLYOtG4mw0Wwu2EtyACH7O22UlmCuj5k6tfV
cghjeeT1aWzsAVoZwLkufj45j+wO6IzkFmL5U6iv0pQtyAXKhPnN5Vdcgmaw1Yqu
Ys9RrE3pU6eylMSkkO61gSEKUVIIfxroAxNGJEQJmd1b4t1NMql0fe4unWNW3inF
V9nXnIspZ+YukWQKSStHNUI3U+f43Qbo4uYM7o7LicUXe5TjVZFZmBY+ZIcy1xLo
5dJCesxeTlIf2CbTJnohgFR6tGrSffNH8ynb5wz2Jd1F8H6kwOKVWcKMx4fNxfq/
E1Wb4QmuiCxohYgWWaQYW5xjGUaZbkqwzYH6scfDRhbLMcPdykH9+gQ+Orbe+1yN
PNkliXFptFc36GYqaBDCoD4BaEBMNLTSSPFXpNJWAeMaB2TrDEgTbTgf5veAPdlo
fVPKYOFcdCyaVjX75Ossv664whBBJApzUVrzSuLDwF9Asb5uw4aFJYmk0f3qiXHo
NRcIIkrNKtHW3q6pKc200ENnIwVsnQunULxdMXOApXl+k6bHomq5At8JzkDPoHyy
8V3hwXUEi6eAsEGegcfzlpicerJsbnGv0xfgZ8xZHH42j10Ngyxp65it/ETD91Xy
jmMEYSqQsA/CLdZ1kJWWZPHcsYzbGI4D/JZO1z/I98TDmhjajFde3fXbiBfFSqEk
CJeH22/zZCrHxm7NcsMR0yT04UnWTw1oN5V6XcddILlhR+pbNJibswxv2uuGN1Z8
BKJKYoj2sKyQYM67gKgoNKz+kZF5tkQBAiynYLFK2gYj8rDHUirwlXVHuW6NVU3K
TBA1Hw9lC6O9Hb0gAIpDuCK20ozL2QHipuRG8TSjjAEHEenIFtoVA+pDQ5paaYue
eycIMK8CV2ERhoMy2OHxemoYu6vyt77Ti1tr5QI81tSjWiWS/N5OvalwuwEWMPdo
oehnixKwG6MASf/zuopvLjFPDsD83S/StV/C+mpMNlKbc446LPXa9J1pdYsABirs
e0iDBrM3G49iVURic79Uf6a1YRKhoJiHyTa8/+Ut+Dm2JYqR+mK8H9eDtdQPpXrc
4JhEA2YaX3M6Cw4+2OQTEYgq4yZ7pTGK5UTxBci9gaXGBIZJTXa+nblZ48y3MRa/
AKUmFysi5WrTjIhhIAlypS5U2FAkg9b2ODYe35YmSsYlwhbgIh1+qwWZUMYwukzy
QoqERRPuNOtTufg2fzJUbGEDyt+wLjDBhP9lpjarhJavD6x0tk4xsUUA29iMjBVO
s+Nvf/e35p0In7kuYzPC1SESS6xGuUrw8r4vodfv+jCrej3cVkxavrXaMrWBKFTh
jbcUBg6XIiTE1cdAEE2RlkX57nE34qu8TT9U40hewWZBfa+FycGMQh8NeRyIKNWA
Aw8aHvtKG8ck6fOdZB7QySu8aEt7bjREk2IqGXtj78Xj/kYjj3Tgq+/+urj0nxin
XuFy8OvkjeCwTHqJeW2p78vdxndDG9+wkNlAFU8qIkzkyq77a/UpIS3v9XxSl6V7
DplV0gjtiy7E8HE74z8qt5ksJgaD0/GwrL7AiAMURRX0P1Azl79jwc9PtMV6qn99
9ETrbTP0PMFyLV2D1rF7xaeZF+DoXN/WisdKqxeDUGM19bjDBn1SNt2zmiRbEI20
iE3DWAPhRimaEkMZvj5bjcbfmc8JERz5jQdYG6QxI7ko4VlwRRC4NpEZ3WkW8P16
8Ml1IrFNKLZHbS0bja90MVWudFoC0CDeFrm/Qd196T2CTyObreR99rZBj7kW0RU8
K+8rddgv+12hk6lX72a6R3eui4684bhBhploEGyxae8AoMUsrJpxhQn4AYAKsu6H
C6IXZ8c0sUXTWsdn9yvJf24v4icyb1IjIAwbXSY/ec3igo0gDj/FhA7RKSizIyR7
Wu7YOE8R+xiWFVhr5YUowYK/+YJg9IIJOBuTQcQ7Q6peSSKqk/h7+hllU0HAUwxj
qSCSD413E+lUeyesTEOA/Vm+7qU2yawFhVVxh6+rd4pRc9a5qZXy6fFtJLUMJOuq
ABJnYpnLKUxglhAaSOj0l916qdVsWYTcUerkZpTHlNl/ukGAZsNF3z3H7HJko6a5
KYjIQBPtmnVJk/CdUcD2Kf/VSBinkyorVTeyymWYkySPcYN0QKXuUdqcvMDtXHoz
cWwSUiLhQ5vAfxmG+Dw4j/YD/hTeUZy9ODdFixaQVJoRfX9J+pn2gy81/m6j+A6S
4ZztsKABu2oYz1luNipob/Q4mnEb3KIQCig777tRyMgVOgsXbVoFbMUUhSeOF85J
2s4Ha70dnDAKm7ucPKUQmPKLxKoTwfJUVzncX/IvKGb9fQUD/SMeyLUuimscraR9
3weBTQy+nDz1EmIHzf5l1xFJJQ/WcNsyeJoS9WhqS9cdqKxP7Meo+mmKRAbr+c4T
ie0BBYPLlynhkBplOdm+N7W7h6ro6R73JIpDxctRLGjl7AwYhvs11KeX/XK+EQpN
s8/P2O9Tzg6h6LvrhIRKaek4hhv5asupRq5rnOLIkricdop5JkPUPPd7s1hzRmR3
BxyEgXNUG8Zy+BsjasxJ8YmduWwUchL8vly1IkCPM//4vfuhHKRsUmfZZp1nQUyh
+bbbRBFi/SPJkggquxhGoaVxQOhJA60obmQUg2dTCPIQzzBLYqlsBSLBAZWqmYrj
jExL9KvIWFNAM4fxrAvsx6KywVf/QNWixb6dM0skZV7S4nKGjMUbMevcEj17E6vS
MRve2VHf3p9AM6InrX3cYi0BEL9YhVoo4uZp9M8Eygc5o0+RS0PGOYIy588/blCv
gkqlBcc0HadnS8lcTTs7//7Lb2kYvE/0zEZcpGaUg/sIXOBVfTHn8rFqb7gOmeun
LVbmTo1DTu4nML32dRIdmcTt2fJLGWPCKObzJIPpvaA16wpA10C0yXxGmUU+MEXo
cQXjZ6R/vK2z1SPQbysYSVJZN7Sv1OqibxsTbhTBngA8ZqoOcpfOt9fu10h6R8/G
ThHU5E4XL54AAJQ43onE+ftyrU9BjETsF4uMQ6Zac/AWhxNk6ctn5IZftplojGKx
knJQH/yXppXCHwhLkmNLCSoLTcINIsIfrEsFO1vzGe8oa+m5vGw4K+OQuBz8CITH
1MTAm/jSuWLsFISuApqu/zVqEh2QMLlNF2WFw3r/ZfnfT3fb7rh/D4TWUoh0Hs2K
4e9S8bxVKxL506gMDAlLkQYmvy+CV8n3JFde+ZtNkiFjLdwcGJz+wWxJANu18Qei
uE9Rrvi22BsAeQo1qZzkRFuYDix2z3dlGlFB1hvRk80CgaiI82jCwFcgkYtAEzKf
YawhQqO4mr0hc8C6udDLjaoQCwQOgxPN+Zwg5NICBDTPd6VgIpuyEXLhOOETgTJU
c+NuJRw7x5qsegKrY/skMCUT1NSbIGA04wT857lTw2blfvh1nf+vt+xlxM9xPSsD
FD83z5AdH9TFTCEigjhEa1Rw1PAnEwwPoRhWF9CuC8uwUo7PI7XquIRzO9r+wzjs
/aT5bHsse6Ct7kcqF88oBvX6vImva6DEO5y+Zj9jfvVY3PM/4t1gtktKedfswQjh
uquWjg5g6l4IzDVkBO7mT8q4MbKvmFDtKvapGGBqHiHmU0VmyokrYpKTWLBP+44s
M2z3BoD2e0OfHS9OgM8THraOFXFiHirK5OX0s2Ntrb80Xj0afqKNJrW5GeWjB0sW
5qjf9jpRX23U4KJvCl419l31WNSfGk8X4CdFPxc8y0/UlEAtaY5QXqsJWTF+IvPW
1JagGN8jbrw+Vih3OOhZ9rwyOSFupwY0yS1x9GYMaSqNBKBAv/iBxRJ4TVWBh5az
Sgv8vCdNLSZ+DebWopofBvm58cVNJ34olDbGGKP7t/YNE1zCZvTmLlJrCrrjOUrs
/FKtqSaXmXdttA7MRQA1gt8xk24gTZ26js8YKlCRLLTkQiVP7SZcTE734kUzZJcP
WSTZ17V1/hOMdvV1ItKHw4rHm1a0HLsfGSDSuYZm/9xGY2uTpLJQLkJY1h3zDTDn
aLgoVyhPl2mr0R4wESGayqxEkRN/PmdrBqAjIO4MiEdJhFw8zluDscN2bX/MEWxU
60SJFiqF7/pamXaBS4hBEEZXmL7p6P5fy8dy5NROGowzcu4B6NRoLrLignQjK7h8
8FHtEbjlGoFgY1hkvTP3WGFqRs676YAWmz/BVuRKkjde2I2Yv19wvGT/cpJVs1oG
YqsMGZY4vRdhXFAlNYEGwComv9SP1Slc+hr/nF8ycdk2VGexKRvHcqyGut5qXphk
Aasr0kGwITCCG7OisbaXCbh4uwKIsbKubHQanNLkM3B2POo7efJdBqsNaCsRr8nW
WYhER5HSRYYnnC76R3HkOrdOQr7qbugZBvLi4NMoYEKmpQkqUpcQj2VFs5ojp2NN
q5Kpm2XDCohwCx/uih5Q/X5JE/+xaqeuK77ukw4FsPddFjOsBtYTFnC1qKx/Yq/a
0NKslun4GEugzVj8357/39Ft0B3Zuv5xZaXc4g9DqX7idR+8erBbS/kn9nE5kD+5
kos3ZOycCRKfrd3qg9+DX0KcelVMnpz3JFVx/gZckZl913kE+ftEEpmlFph7H+0Q
cPdwiDHkU8N9zfDx/1HsRamOS5uAPJh4DgTE/ca+Et1iiHidaQXT3diW3tj8seVp
ZnjgSR+io93DMuMNpJ3qN3lBXMv+Ykgrby4wYQpAHsV/xQlMFNFXjcHmRdg7XUQw
sWb13T1zYdRJPUAqNMk5Woh1BMShqjWyvYXcRUveWtqIp3iWOzcYlPMGkDychOJK
WfxlTBDPaEtDTC/hIz/ARGMtYdZtfP+C2yAGaSJvkH2YqqIim3dyi0QFauRumr4x
iQmOYFVgpuV00ql2iUgW+Lt0hhmdC7mjU14PktG0jRZeDbz/65Y83oHBHkUFk5RB
JQWjrIFaVuOJdIJmzaQf0jzdfs/0ZQlTMN14G2fmW8BKXXTC8VBNOgouTdgL8Uxi
IFC6XIG6WJX/fWbv9w+YZvQY0/THdGAWEqVgctYEU8d/iBMsE4hXFbtNNdJNqFZa
BYcHV1lCjcGj/k9ZpAWcEtZs1D5y74OJTfXLuGkO70LRPJ1M+awTz3mmUEQEMlIh
i4dAXy0212p2APLmVrbrLnateheWjq6ttgbQrN1t+mjhlgO9kWRq7JwXfNyK43Ax
/QF2otGCOT+vCRvi3DTlIExX1vSMTewU7HeANDuEI5KT9HiwQv0L0vGyPocGYi4+
14PO2Zgv49SK0HHnFxbI4lYYiLvhZjw4Y4F/k1wZ0gg=
`pragma protect end_protected
