// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
rwZkwplnFg+lECULw2fy3PcAPhf603c9AIjHZHylcb+SQDBamb6rnerar+FfCPxeE3KfhfmS/RPX
CHXV2HNxbnxbL2JZo9jXx/uwehK93Q1cQcD4iqXmyHpn2FMQu9jyWHW8XffaM+vi8N1KU6Z1WwJU
yNuK69kZE02n4oP8eM+vSvzzDLm1T9EgiXj8Vh9ASvvWD2GB3DLtFU4qd+WpULSmPeFJfCD8LQDZ
gPA/MV9MmJBLmbQJn7D8iO8Zw+u5KlBump9ZDIHmKtihIG2iZmWWSr3zLTiqP44CtFmBXGUmh2PF
DewQQGKI/hjbELJLcrQQyNI1ZwTlHWASatZK/A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
I02mqvQQY521YSZa8NkYQqb8QSYFK2QaBkkqDuIHktl11Zx8kPCa4dKW62xX5VVLVZJg4q9ruew3
GuR4+dZj8uXMop3gRlFfwhU0BDlpSMdG4bWTfijl/sUiGk5+ob+2ZO2FVRNsqu9PW1AwppHvphyt
/E9b/d97+ypTskRXb6kJLEeVFRE5PAuFy5pPqHcQ7vyZagTff17HhyGvFFbyxH50Lk2IttYmw9FU
8Tn9+UCqcwLrAzbbBsFab7ijkSSrYmXmiJkqGvP103UK2h1kFcatfK/g9RcAMhlTb/2Uvl/MbBBH
rf42sFh4lx4dhP06KencZEX1afXdXSKH/23idmTQh7atYMp6lTYPJRHQegz/XusrrYLDYmiPMv/G
Es5qmYVp/sits9SzYY6zYTE2LlmZ4b9X16AhY/V+TYIzQZJsRuxt/5pRQwcDXV5ABI1oYlcSWvL8
PKDocTiA0fPhDiAZDlIHycDMlurfrmeqzJRxfYgqx/LcRIJGfA5IahKK4ZcHs6MhxoN7+0W34DHm
7syFJ42NXZr2pCFkYc5+Gu0rnT0RZwiKEUQlI8QaL6E88L731NRk9rqs0926Y3OD2pm4Wfxkv6a2
zTie5SB4IiQ+DnivPwGO74+52skUyU7ai1Eq0u5AkndDTixPcs+ggKESHn69Tsl0d6UI2jGbG48R
jjXDHNMSXvFgp8MMk+5WxpRtlFRWXp6aNkXUvI2TJeDTfDPJTQCxW8xclj1aV72cwVrQG3T0MVIe
o2giFrWkl4QKADxJX8Cx+UhREN0lerd9B1RakThsX1QHDspgbW8W1XTo69NMqV7qSGl07kFYRk4N
syZ8nhs4JsyuT5vqlrOTlWXLKbU+S+B1+yf75TTwEzgK6nBxEKHYrCGFWXQxgaTje9XvuFL6n2ui
+szyUvbs01X0SBkymzc1A+q3YF+Lx0nTiWxm8prFrjcnbKZnJfX7bEydt/DMjvDUY1uIiWLh5/07
QpN7VmNNWeI27hKnaLiqM8TS8pSzgocNawTrXEZ0tDkSftBbUGpMKouJH36SgvqSIxX9jN46NEf8
4y3SS54DtMaCneDgMO+UxhvdoARl2fiPgU5PXbbqB/Z/GVrliiumq3TJkgxTu3jsJqsr2SRvGn0S
EOeLz/ZEa8CVXmMVxbZcYN6ucvyHLLxrrwZNZvg2VZpRmGwfyBfh9/f4P4/WCN4RjqCO/ebN/fTn
47UaL618jEXJq3rbkOc/049dda3zasyKWcZxJadSVvP+I7rYa07l/g0tQ1dOSuHwvFkgtBj53Ohd
SkWtKYcdgbnPhgG5G2NbQKFbM68LG5DXlb1Ligd0M4syW4fTWEgZNuBL30AdtxOJ0SLX833PErm1
nQEFgyWi7q4f/9SJ1xMyibZPKb6+3PTnmPo3VLd6hllWEmJOtqvRrpXFpqL8jXAzMLiKJAtldrBE
gIcW/nj8wOg/H153feSa39H+SCDZAHBLL6FeKZyPiLpv1TUKaksKKaCWNgc9NFw/L3TmG1z0lbj+
dBhURAFkTTBuFuAV3q1HnKUOoT/OF4DWRSVs+xsA0lIiA8QeF+OoLWstmxCKj9KAYosirgPSfuLg
YcbAwgFJxk0wBNJuccuif7PNVpFkwemCuZ1/lE574aoO4qbPWYFhqj74inrmtZxILc2D6DhU41zt
r7MMR3eMnPkUZIYXzjbOf9vOU+MGqONNNBgLojB1WdmcnmGAVjgjyQvmBlCcaCaW6nWwCQPhbMDB
1pvIMvewNPiGZPonUqPrEYsamQ/VIqKY0ee1GTIcNgR8UA+1qurze43f4bJ8rpPP6Tot0a8Iz72T
Mzc1zCvwrlYp5cQu30so1I/FLczQyE4GeS17nZfa/7w43oexe5d6mKl5iH0aEwyumtnCMweb5Y2L
9R4Xor5JAZ8OhUOH+VaGzTuOFFHkJ215TPO2cJ7MqacRwrKsA/L5PjIdWkGcLxAx6mCGLwMl3ShX
ZN9ac33DkEo5WJdAzP+iF7OhR1I2OFQlJkZ13CavzJEwxa6VB4uxYeUbiOdbR+TYgASwug5Pj400
4/ZyHb4eeiyGwZ+F5b+2HiKEw4CLAbQ0L8kkkFbkrMfmeMGf+sIUwMvt3ROXzgoFWIKdXBO3CKDV
R/Gq8OxawifsHV9+kZYTfItvfKBLRtH6jpSqvvnVdlixFNYPvcsjffSgXpto3hwT0/3fzO8G2V3p
TPuhVYrVcirBob+CDlfiXgmAKuI9P639/O9U7YHoNfb6tMJTqHJfflu+2uyID6zlh/s7eU+24m1L
uBgQS3yg26kUrKnF/GyNrd4YPHwqiN04hqEk56XSlN44PCDg5WNSsmNP+zFQMYC3DPwj42iVkuKN
VaTnqD1Gh1Xz+poXxIJQNrxSte+h9ZHd7OczRMQdqnzs4AefRzrivaswbhrrFVjZQtOkhZwJYS2o
ZMfEsitJArmq7qXhA8CUe98P86Yy+Vy8IXsrT3/KNgBegQHJe2T7ak2+1BSAPnHlUzfEQ8SbCBhm
O3B6ltw6JcPLeZmSe/DTui4BwdmeHziGYDV9NieHahQwYUE2N0jsz4+THN1EdnIc+Mz/K1yOZPSm
4vvjlChm7z6l/pcaVaWFRW6yX/31Ok4nvQx2JSQ0Jru9KW2NHwRBpkT9MJgCPL6KJrrIF1MFWjjt
xpo1oGRAxWA3qg2QrYaG2Gu7AFwMQ+FVBmhK3ZxoNzW+gxzlHxk3HbsMJJmJ019QbRXr61DZdUqv
dyzKM3bZpmXTXn3gO1SnkYhwBUD5Lo39Pu0iVexHbP9Y3PobTl0ueEJnrXTsfsGNKDbIgYr/w7wB
Q8b0TdWY76i4oYGaUW0y7/W5uy8f1I5EvWJ1zYNG+4YhjEmRJanCBZSJynKWrIJI96pCvMWJXuH3
G2mF3SJ9Ox9HOzfaBjT/THiVctgQxQF1olQX5ofddITM/H/NPY3Pa9Pnn8xN+HkDNfuEuLsyh2Hw
QQuwYgqM+eBi8jAsT2kE/q2eqC/nulSFtggtujxekHaYQb3SsHAQcrNN9oMIzOth7d/JnLVOOIQo
Kh+snF+SsvzWFoTVInnTHpypE+o3/vYOgSR92unS8X9FsRJPvrTJtaDQ4I3FJb2jMP1IqZi/QUWw
y1Rf4olDFXbSHMupFPKa+Nlnaps4KB84XMNAIJh9z/sByz2q80zdDOqFaNT2kETRwoOyTVX8IGPf
nCaLF4qGqDlHgozqm7fHklxfVnkNEeSvhqW1pkjygB6Ra9yRf5A3122RJLonV9vLaWHqBGyKfItA
ngAEGzPg5q0xBY1DDoUy3aH5qzy1GP5kRVzLTT18XR7T2Bgbta4MKt5kkNkXzoWpDssxkBOUT+Zc
01R5X1jRjb9QczDy+HE+Er+zESxipdJwnBUaj1pRdQGkfSSWF30h+7Rfc4VlUruss+KMDFdLINx0
fdmeQINodbs+xDDs/XgduXqG1xJ8yWXzyPsRvq+YHa3qr6vySGblQmBKSP7KZ7bPWkjKuguQF71F
o1i08Kjp9RFgEChDN+k+cXWufHeGKFQk/YSNq7qoGYuWACvMFdHYRywLSw3HV/EccvwPjJgXNYt1
rGTQTpmn6z/zpz0Bm15dDv5VyqgTynmXzPxbSC/nyxoz3EVwxr8sIUJCHsbIQRQTV2sYEaH1FMBm
ugRaW7vENMu1TBT3loQGSiFWWa1aBBB6ilIKaxAqSKXVMfnKSKDMxWn+n42VWyysnW2c8CdfixE9
K3SBAWWEKF9U4mWJ61m/vOOzQmlkDNMe2+2aVWWYzzlaVxyOdb8crpP70eAMHUqjsHYNT7nkh+F/
BQgAL/uxaXCoZfHm0om6+HD5Nh3NQoeFCmVoe0JLjSMOyMspX9qsZFb9eK/Mf+yL2c1RhEllfmqK
U1RxgV0mmoQcWiWIs9s/G/bwzCN/ROnO+Cvyp3HMpykaOzvnaTnnnWD4fcY7OWPcaX50Bk9KAMK7
efgkmMx4CUOwMVMEydtO7ChzRDeCS6feuRQ0Zr5eRI7ohhYBWWwFzHNTDJFjVwD+cDhfpky9LO99
a2kgP3iDuDKAjB7roIqQaXUpgJ/RS0+oF3SDKzhKnirfM4d44MN7sT5S4rkTQ8tbkLB+GF8k/GQM
XNfRM77KjJoLLV/v0wUH6A++1LzXtm7L8ZJV7jLUiybPJ30wUxhAdjsEwHbnjdI9BsWCTffqwkdZ
4R6YozDm/5wPQV06u0RoDsJA3JePwTlYhHFx1LgYHwm73BvrPxVpHnIYERrr6i/+5Lwmi3w/tqTU
/9pJrVDqxK3LsqtpMOILIaTDb6Q5vWAwcbdoLy/6ETDAo2X0GSFhn8l9VKjehMd3ykOiEZjZumkX
IehgHmOlgJZFyGD6G7c1NWA6wSTzyEiJ5vgSdFwTUw7jcFqQRAcKsEM2ZmJtU39khU9oi0bRDJdI
IavM8Qp++LD9dYBetvivdwQJPM+Ij9cB7i0JMWyOr4iuVYJ+uSyH678h0uogT9MuBh1/uiGAE/h/
oy7sI9CpLwJLqLkpYFWQCw2wXg/9xDfTKDO8dzpA50vhzyBTHHHs60WzbFQMWiOYmpMyuXqlOZmG
wnpJIwBNmXgOgr3PXC3cvXItUm/2FqYSKov5An85FhkcoUhfucXn2CGyeDnzCA+wAZdQ+ZI0j4+F
JyBfb8y4ThpDC8XJrb2Erckipr+HC+Mc69kzAeNFocS9ynA2EnPmwbf2bEjzknLr+DyD2cw40kIc
QgT022non19pgY5tlRLj6i9V7egAE3wFk077Cl2QvJo6QGGBO4gxf5cV58O2ze7WlDnS7VS1eY5P
yc/PkxfmOAfOOBDjExdah4b8tZGLU1LMgVHi4eGtkEhBzJmxIuNzNdu90X2JNDP5QLW/DOoFTRpA
ih0gus+6Yeoob3VGUmZJzPwcaz98y2XXuD3lHRhazRfvAqxjZEuK5XT4GzLGecPJ1uXuVcetfE5N
bBeCU5FkF7q2S3pmfmsB7XwvIt0uNThR+BRpzx8G8ICKrxmaDgXp5wSr6NyVmxPOU9vO3aXdGFOV
vVvp35vF2ZPNq/KY9SSqAq/RAi8AQni+a82G8DTq3gr1MsR1kYaFc5JDwxus01m3NtYDgTV0dHth
DHXv1SMkQNzOPh/eR7U5qIIphYeOnRFXiNYyAA/ZtIKwVeoGag01ysdwOnX/wm0x5KHL2+nr/taF
Yvvhw+3sqY0FzGFmhaJEzI5HErbZSAukM3Sb3/tYwaQf6Grf9101om6h+YFcw5mvVoYSgXIx+CeE
4IQEtKEx+XcHxXPodlUZYin9O5pjnDZEnUnIinyQ/MpkL483FwkpnF4MYNBnOb9lmZKwcYbz8EsC
tIKudFz35ZMOZXgb9v0uWRHwqUafTTXuZt3APApqx5vDWtdORL2aoHSEWKuAnXlFtAAmDOMbxxxP
MYETZMAjr5889NSyhnOVIYrSTKxe7qTIN4Nk7r65m2SXcYRXxSfMQVlavj3vVF2MZBtuOwStqKt6
7Twutej81M3sqpoKD7Uy9wZBEgEOHnWMO0l5xxOyrhSmZx52p7EFc+RFyrgeGS2fze7XkVcc7KH5
VJZWKh08VRqeP09DmYGq+2qT+F/bwnZT7LB0Hky1gQ9QTvskzwmv1uPVL1fBTQpWBvSibXxevVvr
JGjSHS4Tsa7iQuoIs/St+CPke+dhnaDQG/CaQgLqJ50ovK4DxMxFCG32oa5+JCRRQXnBpEC6vge9
S3tTM6YdUhB9n3u6XAoSYYj6BRYRCgrfHuC1fJKRWnJMo4OPy4IzSz8Rs47Wrhs6VYlPjY0O9vMw
1iHRXxDfzzcfkoqkSO9UHAVqkV+7e4zMNg04Vd9iqH6Rbnpzrkb/seuVyWmPS3jndjtK+8qDiFHi
G2AxGlCCsILHrxuCHmcCfPh84uvD8bCosOXpThLO1P8gSAgZZl00pACjJdz6LbP1bX0yUKrY4FkN
bNfd2J/95jaU2OYxwuPM9jSeq7+7cjIUSdnvwtEnk39dqvwSecNis3QKOEz1Hbb/sqbhAomGYxhv
ZSHzSA6TVuJpkWNH04MyirJ9logXwmyi/pEK9Hbw/+Z+ufQhjBWflb3/ih4/t6+tsyVdHC3JK2Nh
jicQdhVBUFrw+xdKD+hZTQSyvyn9B9cGDqUBFWlOwff/tPoAWvt9RRZpEKnIon4YcrWuStxKp420
SKpir5LwEpikzmZVg+JiukiANAgEQviGkV6bKEzsn6CZxMCplQ5oxPgk3JEN9e6Wui/Z1J7ZMtLE
rcT+fUHLML+vPR2Slk7RLdorNB7bx2igXBBnxp9TAlCLdKJUMoJoZL/6Ert4cFNC2VxXbg37Of6o
ax9X8Wb7K0FMiRaXPA40srW0sFxsg+mwiura+nPYeyuUw15pYe94VBtGXgUNDXLnKSdtL49DVGUK
eOvSgmPtSGveBzOGyZhJT4crHrs6XQ6ExRNX+txBUVz6JHFH8yy+LmFY/bklkFcOHQK3nNrPiPH0
pqe7YS8Q/IpQzsVjALDhgv/Ncl13cAw8m/GR4OuAtxpJx/niHwYSfd4atpem7b8zw5LxRL2URqji
p2Sg13H7BcaTiM2pczH9P4sfsjij9yHHlefowC+BxExtK23S/63G0fVs7AjSVGaPu96D46WkduM2
9pQQVBDNqj4ak3ni9QLMm83vVihQEHrMZsB2XxVRBQ5cNhmuLj5lbfnnTGXmmfJrpXi5IysiijUN
X6vYPWXlHUdLmDsPzyyT8OsZlk1ncyBQJzBOAn4CdxDjZZr2BBO29rSVog6btGyVVfPJYytP+F49
6WHhW61zQBEu11b/mRxZIqfryE8ZlpuEcV1epK/pTAGl6VldI8FmP/Puo5CGQAGTaxTDNBZ1wj1y
q2pgm2kXXWGe97USBENFq+ryltaZ6M0sNUZhT9ohHDBiGR7pxrs3VBhEal2B2eVJVRI8at/3M7MA
yIDRk634UPDIOYTU+9g8Q/DD3Pbz/HbmE0vn1wy1SI1guGBk0vfWgH+3hJqQIIgsU4ZP4ij9F9EO
Cs5D3ZlzhvAjHCO5FYBy1h3KVo98nzYsWjVKsar1gi0WBuVterDyjc+x1lCsQDyuDQsVpY1W2GzD
6PK2XVpwqovdexHVhjUCKh8KsZcDFm9jJlpgbq3kw0PJAlWoLacMTlEZ0nywKrigtLmGkZylI8Kn
SjS6FxV7DL7sIEtvR1QnWwhm4RCJ/tGS6AjbnRxNPZaQsKFxwsNFYUY1VuijeuG3XEz0rkv4uveX
H36VlxlUkxJs/LEJ8w7iMHga42PndzG556ykiwFz5iSAo75Dpgz0JMFIiqiTZSmMWtwmlpXiGlAJ
0LXL26qhlIetuM+u7jh66Z4OLBZt4DG/H7GvY2E98LzVd6jS48ZFi8zqSAAxnTJttnrh0Yeag0rz
ygn3ceArpfR5OBrCIrLfFufLVGXMaS4dQG/MHfXIEEpB9qELJHgGVi5/B8+fAXvR09gC9vc+K4gD
VNdOkySplCgcNVR6GQbTA+lGOtTGWj8JCTPpRGKz9eZjzOm+eTEBJampFedmAhgTD7ukG2l3wOkR
foXAg+p/kzbq54ruJztlyZoo9E8xP7YFu+1sLh6rhrHxqBeIGxtkNY9ETLDf6FwXhEzZ2eDRAond
ibWANA+xdazzJE6Nq126SB6HmT1zGD+qeMTYpISTiwLX3WqQnpiY6JMfsqOmnftASOq3dTIyJl9m
BdUipf0L3Ab618o0w7aIj/h/PlAkK9OtuikGg6KjcW+SNY+tSw0ppiaWwr9E7z2QvaNrTGojWL0l
iTbeY42kf2aEV/xATU3zMoguVBxU/rXBL4H+TsBHFWYYE+QYA94mTC+rApXaz/VvGKe5bf+EksOL
cuwkL7Ky5U0kWioqSURiM8p4Lg4WtHHwAcTEmDkoc9RXVaKfqxO+W+5tjYt9if/DrGfLBI6hljpG
igTrjB4pRL5VV1GuCkuQJvRjS10fziIPlaw9NDIz2TC7jiCxfGCTevJLlQsKItD5B2sbHV1vTPC7
tNbP90ReGV2PKyXLudBrH/kePidmyvBUQBxvx/HCx9ll/AmyuFG69I8h0kDIX7d3m2zDUMrTddO5
y3TxyJ+hINZ7F8gtLOSBbtrOjgvl8UIO+HwvdpUhBFl9EAKuFkRBK/z0y5xxFwXR7Dgl4kiNFZnE
pRQF+cMNgibj00RL0A==
`pragma protect end_protected
