// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LRefxzyt7kmqF6y5PFZbN81Y4Gf0Wv2QFqX3AuzBGFoe6IOWTYT6sVSfeqX0PjhQ
eKuJWA6Ov0ZS2IpOOqe8oaZnipGUfwk0Q+j6ovT86Hu5r0UpwJ2BV7ZBfFkJP2xh
MsjCcg/azxGXtP1kOt2AlyFsCfrY4o9kRRb3op6Mlk8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7392)
cMcnnHHxTk1P//7fA6jWWOhgEscZIAPQxog08IKlngw1nw2mROnq/ZEzL/W+l8Oj
JFkd9vXC0oiLLIt6mdIsEvhJSZXQL6h1RwAq9Z0NPfBXbfW6KlmfzguTlNY6K3HC
UU6KOyB+3rp1MMAMjGXNHQ+PUnqr2YXDOpihbkZfFqeUEA+hgV5TlIOoV8Hue6dB
Ks8mJjxH/DBaXe/Vnw3yZIoiOkB1LjRrR6GaTJ4du8bhlQlIm6WjpDt1jCcn1iBT
PsVHCSn7roluQcFm/6vrZiLHG1Y8QLwRR/Fk7LzVs3hUI2gfwLKrekkfqy4cQd9Y
KBLxCR7UCoDgxxDS3ICm7nipBN+W7gcs984kN6FtRrO02leAqt3gl9QJCOaopGFT
ICRkES0RyMgt+qixnwUAZbUHFHA4cs1UvHa8GojhcJs2/XOfaMarDoLVu+EhuHa8
+n4G95XFohLsh3iVLAFKwyqjBqDmdd46aIPVwziEGq26/P6e6TfOEZ/21G5O+eQq
5+xAzVhNi9/EG2d71Y/ixCtB7/OhAGFFxiWst8zO6zdL0dd0jZygXIJm7Vr3pc4U
Ij+SHJ5cs25z2/UYHqZcYQi52iVb0coMRQCApywBokDutlhNrqW6IcTzdcCBAqsh
aS4DAY3PAAN+tjQE3T9i27GpopxLIoAqbHvduYaF6rhFg1HWXOooF5bb6ahGNdqX
u19bht/xfHW3dRNmYZ2pRWIjw7fIXz53NpVraFfyNajGlJNNXlS353HCrUVAdV/i
heAa6tW4Hpp0zW84lCYFSLD62CnlwCDbUnrBKM9paolBa4EInJ6Q78o/tSkhrnzN
bPQAr4+6cNRBycZ1g35GH7s7ODqT+pVwsY1y7aKlWDbT8pIsMYb7ezjVk8LmVIWI
sXTzyTdX77AllQ2mVNzzKvVJHVtpLECp7YYVX5DZyYmxVvrHjUgbfXNSpFQGYLYM
gAgZuV4zpXaDZXemXnJ42vF4+20AOBBPds4pWKkh1LaII3GgnDBGgQbzuE4XYRBs
guUslsURuPJC0Hy67KpuMslsvuSUmGKAbRxKch+lb0XEB7Dz9jo3EMCtuBry6dQH
CNRzd5CFP8zfcWE8bZzFpGpsEtkPzdQ6JGdgAeU4i0b6SEMwrlk0MDGlgi6M4WUj
TXmdo9th/tj/vcdz7UOoeW/82EobbvNvMQPHFjEgeWM/4Enp3FdxVwSPUfME+vfU
gX7g1Uo5USMpyDUdIyDEZ90w04mt6BKnXkx7+ScofJfFYDVfC2Qg+dfDnoIN28kp
dyKwDtqvZRaaQ2VTrwwoHshVwJjnHO0/KFwjK8kUlMlHyVMh2sXfHyLuyIKOVQZ1
MqSU81qgpVVq3CmcA5zllGK2Lrpz9YCnlrXajSZz/tA/gHNI7oodbS9+i9Ma2aHu
6vLDDeieOVvNdS8PMiab5MnVp82tY7BabVDLOcb8ehk86q/zUqPO2a6yUFheW1NT
2OyzqqxQr872uezbt0oV19/Z10jItDSiCsFu1ZILdqaBbMVpfj3+3QAFaYwbnfh7
VIY9YFQ20uslQvI/aduTmfXuVStCxNev+NNPOeeeCknyWL6HwFuD8rYEvYfivmSW
fex3Qx2UgPIDCrJVHPMNjewHVymRRg07uZPLcBHYCU/lc5vZwJblGiyQXS9Hv6CQ
kz8pSt6uJTJk+tZqh3bsZzVJz+UAv4EUdIN0nsNctSUvg2f8Acr1Mpn0xOqZrHgj
9tge5Rkf7deWyO/GlUf6Z+lMeYWGtEawfCQ+OI3OOmX9r7hZ1FQIDA11oesKpjZQ
1m0RKSHFlIE0i4zRa04MwO+p7cC6TXheIilDEkSwvC8PZX2LL0wFfMxskwA+jIzp
uW//Srt0CgLwtWcNKcfY9nLjqL4vz8Awq3UmtsbW+PPxLehFPt4B7qK769uDc/Cy
OS6EPy3kBaOTitWQfkoXsoC9XuNUfJ8xcLAM235UFtOoIKXP7n6z+tAKZEYI+xTV
nWGnMFMrhVYPlVBRp0BlX7w+FcJ1rznpvYF23f83HL2M32v8uZL2zm3U9GQ0B4u6
UN0ZTXoRQw0U/4CPSEL33BGJFPuZIT8gUbw1WUZhNA3uF28PIzCikPjfpxJjs86p
6OGO/zoF5o0NKeOFcnR8QBhvJkWGgSQdUMkajnu1/tlcZLPOC/0hQMPPRo/IDA9H
GFgcxdR8/1W6hLlB+ODM1sIA9aCLWPLkBwcBMm3YLVMw3ByK9NAOIhYiGN4BNUL6
bEbhiUV99Gy1H8/CKRVXthgOPJ+bsTdLDh25mwZxSM+xbjZz1ixzAR9mikIO3xvJ
e5t1JIRCjX4iBuVpTxsMpvDPwF5zaEDKNbYQMBjfpjaUczWA7Q5buPcufvLd+xsJ
GzsjI/CoblwvXOCIFHiYZOQL2JIB4qKHm7FxGry/a6HEDMtyKu0gOd3rvNGlKuvk
D6SM5bCz86w0YgUsG+embZR+dHNtNCoMDgWR6hE5oRAd6hKjKJ35kdjWSnkHYK53
d2o7Q8JpdzPvCqkvJprKX5NFrCTZsj+1tVez6R9kK12q9TiE15POX4XKiUEHalRe
mAGd8yyldxHsXxlBi7u/P0jXpp2RUOUycullWnbuZQ63g2t79rc15jvJw9Ts5NGs
YIbGo5i88x3g49X2yzkaHALSbnvcDzXvFnW4imSRByAC0iFGwVQGda2AXjccb66g
04jjBjES1QLkfWxnBxc+zc1mWP7ap2IkOpN+4xGMtvle/MB5PspXNrskMOAFBXtZ
5AWM+1BO8HO6dK6MjnfkZ+zZEeFRp8EXJlS/4yg6W+kde8BFPicuXyQXVDkoyzq0
OzPg4xGJeWxlea6/smbff1ZbMzyxbSGsHyyFyQphHg9nz+WYz00nV1ym7NZyHlHD
ZgZp6Y+Cb3nmiuV0quVtnqitJcFjOQTyuuhgspGlXllXNMNCI9bRcvYMP0XJVE3w
kRbXiOpSHIkPe0vRSgt98Kp/+QFUVTToS9Ba5gO6WFti8aL2beRMqW/eJdsPbRdB
Str4Qfa2v1Ak36P5K9+KOXvmBeoPpVN1xvz3fXdW0vSnXSEmOM6KrOAZPgEcOXmE
YuzdRYczgXlz31fgegrA1S/Z5Ib2PgYNzNNknjHb/0+KsnRgAzLRf+eiLpG0EZLC
mE9GvkcWl+yo9P3dYW7sKMbsuHy6hdSMjw/ZY5Z70ounSnj36i24LcO1TPwHN9X0
e8T3dTxIp/eF2oSGhQpWOvGFgymPzc4aYT5nHzp7Wc8a8LKZbigpO7fNoZHhY7VY
okCcYAM0epjRjQuWdxnUJDSmvw9ZxXW5iyCL+u6vijSUInt+ENCu1hzX9vCgV4TU
Hry4CPDdYJzjCvW8tGJQYe2nmKVUZhF/j5SL3gzld1hlanOfuZiA7ZTC9xSpLyLP
WSAg0pbABElbf46OmeYy0ut/UK0Z5KgAIF43d04Lyf7ABsF2fOHrbTtVfOTHnjJ+
QEx6p/uzj0Ht3DLcutuQred4IoscVPMpckd+FXs5/N2kEZpDZ27JVfV8OcLYQK8L
l58fLhfEc7wErqvKaf0Lk3nHMCEpJWcJJq1n/01k6w+7u9+nb8jS1EvZ6a7JIuFC
lKR+DFqew2c5DCdMFjXQJNpD62tnWg+BqJH3NC/NvhuobpzD9sZn3bOgZ/bwYwGC
nDceaAG+Aytzkb7QReB8YOOmefaT/RH47Y/AUngpzlMgDGznp2yTA2k9tiYfAS6t
GvlJjHKu6yNNpTPd125nM6uPoNK+3fGj5h/tg6Squ11Ld+M+WVtoPqWtEi5cBJQe
KOIQBrc+waihHPBJlkMdM1PcfZGpfHjzdR7/5rcXW77QF5hatEXrxROJyMPK3Vbq
t5obo88bYjrzy1f4oTKfsOlTzq1Wis38qqabuhTHPezoz7iIhdkekY0qP9TKdyYm
oZ2w/O+3xCa2u40lgAIyBgDlTMfa4zDDtiFKanLZTsckqOj0QhL6mAmJommlEb6i
Zl+ZOTI7P/05ukJwXas8uKmO6eVvFHG6ETGI0Q+n8GRNE1nM6lmwYugj0cNAbBdu
3ag2NjaM45UEWwS07vBN+aqieygqK8rJOjhGFUMxEF5zztjuO+R27/yR/oXKjfpL
/xTLPi3lc8Rac5LQz70SLBJjd+u5P38zJSAUv+xVWuB3XAocKuzv/8o6ato7x9e3
Uc7xyx91b8mXZIdIVAAkNv8gLphWFphGZ00NwDRnRi28/n19wpx/bZzk3gT0ytwa
yjoCKqNlHrQcjhmyp1N+80CWVrXHWICmy7Uh9CTKdw1p05Pj0sqsMAk/SKBqBC4l
DLYtj+egJ1kELeTK/itcbIle73jz2hM74xlrtrp3YTs3vB8khr1HLmHr5w7ja7li
Dg+oeX3r51lar6/XuNzngHRwEg2dMz4Ca0F9dWxpMbPq/SAXYrZobWt/QwBm0cLo
+bWNriiag3sZuCcrQMnMLTYM0pWYikWRecIKXRkDhfflBu4C58OoN05pYABacILL
yk7k596GMcOTiYvRDWjeJXsDVbEWMwpWxXHl2pIEzLA/QMZOvigCdxWZc1WpyyAq
VRxqaTDxI+w8JgxUM+ENKHyc8bbNuYTxU4bMeQa0R6ZZd/xL7EpoVzaiD/rGc7cc
+iiAKlVJsvR2z3RgdUQH0/S8/m3ifNH0jis5VxrjTmN3wBoBMv49cRr0tcBRUTQ1
TWtDu39Mm3dZKfX0lEQmxMugERp5bVMzKIs58x/iiIZtG+FSlLt/VbLUm2T/S8QP
jIr5YT2APowJE1cZn3D5vBuyX+2U4ivawdQLUkb4yuhgcKhnD4kPVcbxAVQIzGu4
vOKbJa13WQvWIHwsDihbjw2mrw7kxOiIB0KnczMWr5J1vCNbU7YFSMY/lL+uSlX0
Bs8pKwWczNQDw6lmOFFNxrG9X13EAqUWymcDPwTBV2vJYFDW3Dqt6pCaSnCZ3849
Ob2Ugrn//+NI118hAu23MPD2Hkf6pBd4yJ/bQyKg3cFaNl8USsV28XIMbEP3hAM0
fo/kzGWKIfgYntvkeqEpPESYxH4bMzfXFBlvVAlwgd1bkPrLbw8OdgiK8TFhaNg0
MAqXZZSgbv4AQyAPWDBCaFUntVOtzTePzL5j7FZGUI0IhpEaLjnCNlVfwVs+Zqiu
/AiKyojjo8P7p8dSsGGDm7suF7CX3GCMGyTPmBb5gy2f4rIA2+PiFJIP5ojyDKRV
5VXsvUfnxUxeN3CAxu+un6oZKgMjQIFvTGrkxxnGmpH6d4797tQzDg7MoH0dg1Rh
GGD4uRXQQLfHVmEhC/nWh0xqrbHFhSctGBn4LmwbjzUQRtnvZOXL4rXivVWkkmnN
4LBZBFJnP9PAaYN6zPVezvRLJlknM3vTzbr7bYj8F4Om8XdSPM2rx77+lfh9QYW5
DD8qgrSnimKAZHaR1gn57iXVkg0gC4n8LMpbDlTclvwgM+E5YqyCZrgOvjBh/WXh
DOSs38uStHKzbXrDxq77a4Zo3GTRX/KUdFFrum5j/yPfFjDkXUxVGNC4OT6eRJpV
KGFfNb+WB3IfpdYtk6z+nGTDaqGz+L42Fe9kgmJJ9mYahfsXw61ByxSliZNmAgFt
wh99vvDKSezBAWCcV+o315BSLzFJj5FouFnqjN/CpTJtVaf4PU4FUI2CG5x/aYj/
cM9n7h7Fj6t5a4xqzt79XSazuo1QSGAv75IfEvcT1ma1r1aNmg31ffoLK2U1L9eC
vKAKufYuRV0nPHwuQvUfphrEXQ3V5LtTt0LCVZthbjB4rDr7GwDkucU0AHmmYmmp
F893406AwRddUpg7Ny1dXFtLrnWLt23bFQQhJQQKSygvDQAeeP7V3fEJsA8OOflf
0+dzlNu2TvwX1DA6alRMpU4JX2iOahWfQBdrbAa8ZGuMukaE5eHaK1/b2cT8lI4E
qKTYfutlft6pI6GQaKHQ02ep/VPFGvQJ586vDdukhvp3SKNwEG0CSqyYmbwOaDKE
YMo8OxuLq/0OXcFZpqB2CdMRge741E0YS5wAuFifArrgtNLOd0qXtUWouM9ge0mF
CjWjGznTMgalJ3Eqe3dq6OVYoLG2bchTWbkC0kUZ3OhaSooJW2xk8eqCmHgfCWr/
qT+qQT6RzpDPBjyL3LSeN2lDcZWfscWqaN2bNMvTXCW2yxyyctyac4GfqwLPWtk3
O5UHW5XCeySaIWDTgmJ1wYqi1Qcfl5+Wkz8H/9Lqcn/bX8YAYB/RwS3NKzawaae9
etpgtBApMbrUVMWFe4TBKIKzXVDSpL6CZm1EufbnGxLR3XVRTHSDfQSJ1W7GF/lJ
0cGP4PAQ8lPoJO3qmAgetoWCRsUjG6DKnQkyF6LDrEYGZcoNYtWcEILfgVCqtcbo
v61nG+OG5dgcCqbAz/XPeJGRspsrIpN/FwwK5nTpqye+u33RZ0LheS0HdJY5L+IO
naiSBbSskiwCR76O/GN4GEWczXDHxm4+TCEcINlhL+1XTx+MG93hFRh8+GCdtxHJ
xCBMv++gKflHehFq4TvpBnMamtJQ0R7nyiN/Mo2wbRGcuhm1iT50sN8osKxK9bTb
3Hfw1iobIsErHMHGA9VGwW2ofNU7PyYXlzz7ggDV2UB1sl8Qa8gHgZPAWfAM9yTn
zgoHznbyTtB82EqX9hAG3eD0mMGzWTXOpt1zYgZNI2Fjnh2IBFO7UyyGVpPveSuA
8nQpfS+FU2VeyyksAxsL8VmN4idnDQD1j3hdN+brq9sa5qt2lBI/cHY4Vs/15fVa
tQJf1XwJYtCEvqfcqZYlZrBBBihwWVpzjNeHJDqSUtSgmJyIP0DSJZOnhd+++T2M
1fevVw28+da5ABMHS5kTsuSx2L87cBlBl+YbI5QCVN2VsyYJnnW8K64Cbeb82EAb
At7i20bcO5qcgpCLMwhFQUh1sgTKNbHz5O9/jyAa1dw2lOnn9lKcRdyQrRQ/XD1b
BEpyUAne8trjh/RUaMhgFMDKRpyNKFu7ExCaDypGcXD76C2s6SBaGgSNAo4jl4Dm
TDsfcEP6fOGXKQM7ac4iWLWaQm0qNQVGEWrIzjeueviCG9cNOAT/qEylqO/vNySn
l7oivhVKiEc7lKEfOu21uzEE8bP7aAPl8y4VlykWdDavNmbbpsy3QxdpoQ0njBDD
dBQcQ7ic7jnE6H6vmRGaSBmHEf2lccRzRgDTovSLw7bR7+Do/Kw8RNAuRl8sDmCE
ubPtqXU2edNaLjTU60hn45zCcRu1e7hEiQbfls8BivPEAsP++hfOjR1JZkL4aZ01
3+J1DGwyeK88Winuj5Mu2SMbx/94G5bFnr4KWh4er4OHX9cJkif4X4pdXPts3g/l
CCgub2R3iHWHweTOwGSS19TxRm/wJBrhWvmOdKmAzXTkA0lNzemPD47TkY11GsQL
KrcZzAQc5RzPChMgfCtHMNtvV6e7U/WWSmORz5djs29vis5PCo4bcWGSG1/639cw
4h2Vw09ermlTTNA6zRmWsVyy4E483iHIvk7SHsfTniKlspV94zjoCqlF+XwWyJYl
DqyToGhY0mfrZFQCcvA8d6s3l6i0ld9VIg3yE/U2o2xZntgMV8jxQUMHlvsIXQrA
zGmx2H1RUfka3FPt8jSOacxH1t3GPETloGh5ONDmFi7PwmUm0P8LqqcESoWn4epR
NdSgo0lCgxTi8/qfKKHOG3CndHdwMceopAdhHVlJotp0XGNeXoNbCVRGFvHwXLwL
/GmThoXf9zOZUDRQjAFftSsRfreclMqNCr4s6hLnIXIEWZuTlOyum4Y0KqCCpvBt
mboZSyc2yQwAPEevLG6V48tPj7+CsW7MPFPFwB2phCkiVo+WARDXRfalRTt5Q6Vh
VStitUd6LULOOJWfIuvZWOKkK6Y1S5SPvVg40aPYZxRsT5y072VI331/oiCduXiN
B2uUhKNiX0YrIrtlGy3j+yTHoOKtaL7MVa1D4sy0Zak8xzwwZtoYIgL0BT5kVKpr
SEcabWSiOwjT9cVbJUG9I41mIMLnTMxXtEL15yE545fc11tS9KWtzS2saYXqhO2P
VTxSzvLl3yfbNOiS8c6g26/Suum4pIQalPRNTVFjY8gmY9d55f3yA3v2YtBOyUI5
iFkSQiWHZndR6Idq01vGkNFTpr8rz6Hq65H9AGKSND3AZ2jgc5MzEmCqaeutC/OZ
+ItPE4EoChywvybu6UFaGgqT5DLj+k4sr9tgX+c0QsTzL/i9JHR35gSH1v1Akgi4
oseSWY+BcTkennANk+HjgtCmlM2gxnLr1VSpucpuByJs+uhKg71ByXm8WeL5B5s8
app6rmbXsp9X7LwkFpAzAW8/rgUytRH8pwdwr9H3jmBDvPZnpfUtJoD0Yp66Tile
L+EJCrNtnf3ipFH3/7z71XyNVcUxFdHU/iH/7DgkEe1WnVvKtf1gR459YdcBJeOt
gmBPK7EW5T3u7SKbRM/LxoMgHRb8EmHxDnJhmUaXgelBagX8moP/QT0omCnKbo6W
n9EpTlldjfMO+bxpKEnlHznV7muYrzpjOw6Tdc7v199jvk3gYfw8Ivai93Gssi50
QTa61KHiKzg+nMBvL7iLoGNcKpTGyT0+34BCwuWPYhQLzpKqaYWjzZBMmFBu72tG
RH7ucitadOwrjDP29rn0GhE2kjZ8emDN+d4PXp7v9hNJVJAei9Ht2lUVsTLLTZxY
TPCbsJphR5Qla8t7E/5641nlUNYz8AESl6v+UHPbXtPCl2jgKv0X8poaJq0+cfeM
k9H1KuPCNHvNNuQMgmeB3JGbJZiPrRMMy8r5PVZHcGVDrsUed1AW9pvMyOVpImUD
llQ3nlKnYp/8qKH8NCrR3D/6rrBI45EHDZeiYjsRVvHiAnIQYHnVG0tbHGU/KfEg
RSTRRkkeyrbG8Kxpfc6qBNq4G2HUFLiNImrTclhEIkRw4eZG2KGHWpS26xj0ogZg
XAeBQ8i+3/wU60guaTzlqSYrYdsYhO+QQYWyUypWA8jhI0Tzcbop4Xya0lQYJ1eq
Mv+pnFhKf4iYC0bAi5uJlxiSG0kbyGvE1UEli7BpACQYNqfW1Z+AZSW2IQL4yZ15
AkrlFkejVGhdOeiKJj4sGSFC9SdO8trn2P818KLat6bHXCGqysPMa8hBia1JF091
qnCkfyJ2EQAjaMK2Z36kOeTuho8M8NTAouxWZuLWcxbsDbSzV/5m9yrQIgu81yHr
UJniVlRk8zUMrPFpQzs9SXj5IAHOC+o29lebDPpyq9MOYSm/2yM3w/t7iFjEh4na
y0aBbnUeuGMyYjbp1I5qYfHPDqw/+o+1t007NXVbQXIBsgLhBj1ckoKyjW3yUS+2
zMxSWcGdXZIH2bQsufhbjEvGOKMTq54xt+8Q4f/SGvjpSGpdgg3HI21a2XgTmg6u
ta5+94ltSdQXq5Q+BrTcPFuq4rb+F72dvPQ2BtjWpQ6JQO35RWilR++oCSlfNCFL
vz+61PbGVKrgrpDoFkGqaoqpxxLuEP2X+XsxcfiXQ70jA2nzbXuy5lrbJi3U8fUN
6JlzEUmF6v7QKKIQ0lEhi7aW09685e0d4UoQnes2ANqXS4T3nt4uS6wpmbzOMJTj
5rPpeTmn4RvUdrxW9vtpIazoCjOWM22xxAmwcfUHRj5nEP4GhJys8zOGMYIL9yMa
qfPPrXn8UCo1SQj3csnZnNAsecOkQzZ4BPcehH4/ixu3w2XW40gOounQEskjs502
UnDerar8dEEOT7RLjoyX26eA5X+UNaB4v6gabcs4JOM/KIu+WNb0ZPe8M2vxVVh+
7YeeKA54HF6TCyyUqxnKgCZgJaahIoC1S2vT6DiHYl5emDZEb2hfjHbcOApjPoHa
1oEiUCWQN80BGKkuv7tmMOgnb0K0prdnrC+ujsK5dY21Q6T459cK942nFbo1YXRz
`pragma protect end_protected
