// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:42 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dJ45GmiDaJ0BA0QbBLPhkr/LEH7QD1MHSTF53ubzgSqlnB46kUbAV5GuRkoZYru3
Nmeynix3+MTBXyr4x9j/wSQvseDsJRYv07UXtrhb5nddJvv6PGY6+H/LDDqL8JM9
JmyPa0+7Ld634yAiz2WVxjlkf4rUtsQa5hn+pd6+0fg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10768)
3CT0NeCGDwnImN52onR3ihfn/7lOoEB/kbbwVgNUizKqLApyudEzAB685hbVrvyj
mw9NK8PH4j4dpINGEuTjVUWVR9087CL650iy5P8KZBGJevJiVzcvmNatw3y6FO7P
dKDPtwqAHJxMEX+l3G7CFlpoHmV0ld41JeieGgg+k0d99f5hs2/Mf0CqgApHk3G2
ZUBJzDrMq3oorpOVS6usg3zfLzivIBvwTJmaJUkupRML4SoZQXfXNvod/6H1iYQN
qEGgWKYjFKvNrrhWWH1ulUVqt01JttpeJS/V3Uo8qXouIVMSV4XvLxHkt/5+uxLD
tlU+yOTrDRUcOXEAd7cMwfbwiFrPNdlMM+mCO3eIJCrRkT6jpHDQvDxPzX+I1Ix6
RuG8nyDI7Qlsf92NTYOhrCG8yL3vPN2bQUtujL2JBmsF0raBQKTnmf2gs0/BoO3R
BYM7J2qimGC1m+N86UVqNgQYjcCu4nA+29tzwL7BZBmpRIWz+vNgnB8bdfIwbgN/
trBdVd5HzJzhU20dqE2oR+joxeuqXL8abDAkklyOIA30xaUF4mDpUpRY6i0pGRh6
D0ujZR1XpAFyl+fugFa5RB1Ne1wu/Hr+N5IUN2OQrP/UiAfYcUwtiD4rLvuVb7zK
OXhmFFfLbnI0DaiRWvOCAYXnPMYml74zDS6CBvbrbRYv+RF19/M9wpETtHpbHTpX
0desV+qD3G25rO4AkI+tm/t7zv35/VTcTZC/1ed4QCxp492FVaN9ZmMgIECQaGS+
HUpUBj68HfSqKEwMkWANP/NdXSn0yZcAttFUsc20UtHUnXIqOVpqK3odilK8YOll
/Zk/TFc59LQBD7+RGse6gRbI642XuJDMlMPxpUENjXZTQvlGuMK00KgSfmoyVQpI
6vxIVYMBdw1VsDU02aiVGS0H+cwS+ao09dimq8UBsYsBvdT0E4AQLl2+MJ/sDPPt
NOs+RYXDadzyha6tWqTtLUB1Nw/OIDm47qWgtESAgQmY2Q+hW17cjD8kb2VCa5rf
9EtKMf0xpO1PioQ2xjg7uW4XCqBBBQxcnHQJ6D9NYrxHhOZW0iCXrb4PdOtaO0gj
mLABcshyRw1eq7vdyQ7YduMkoYYN7dV449UoLTPhxxCJF26MNKM2h50a3qP+FZYd
hHDyHjfkJSGULsu9QvtcYB5YqYahKATYKlkAd14s9ZwY3SbbYGlqA5vgR7z9aT77
1wHaiEpnCPatx8ISFnxBl8zlqLoEAHcgt8UlTSSd9wmt4Em3gomcJbkU90cqHXfK
V+ONsSikkcaj2Npi2HrpdgBYEhlDylIAPSN1FZSMMymxarwp8AqrP46zLTzZmx/T
mZTNTa5jgD0d/cwY7nLrUJAXUrmm43fTx8MwuWd0CuPWv1g2i0OGz37x312LTURG
BAOl3hdkuO+lFJTyHM+j7VcDSnMNmC12scSh+EJ2SCJWKq+l3W4v23/iXS6HD7nl
DZdJAR1PJxr2ver2ZHjY74QUDygKZ2Lzld51jdni9C7Ddv2i64rV78JIib3Sg7lX
sND/7qltJY+R6XPzQdW+FM8kfWv8kcF9tzxN/Uv0TdBJ2SgLGiT89m8Ml51cvk1I
i4hwChDxPfo2HkAHXi6CsogCrai2byjQHqiWRTXachEU/d7vOawcgf04ZKVPlHNz
qv9v83o2vxS2sKgJO129egFG2TAdtV4s5/w0vg8MhF87yWiPDKXIEov2+7xc+OiY
ABUJMCDP6qdDzpN+S8nGUcu16Xpz5LC+u8BfOUXAXPp1gv6G2m5K6PU4+HrzCaC6
PW07ljSAB81khpS+BP4iBLEOKTERH8M5uhU7H6rxiT6RTEEE1bpkwQa58DDJb5Xt
LtUy0Wzh0PKtMMCC9yhTru0m0BumT2nYER8f4xfQITAEAN7UemRWQUG0soyp26KJ
8nHfiO7k6Dcw7H2bKQexpqiudbgnkLJwC5aCKs9lixzfaxqOP1dAchM8fpjNB7DX
3JAtJM6kllRMPYILAGYHMQPUiTDU1OCNgJPojn1Jz6nOYGNWDZR97W8ew28MBHTC
bhkecl1ME6GQQpZaPRXPiEzcVqMsBYL/asIzUh2fMIXuZMuTbrjudu6dm0n0fGjV
UPlBEwzqfd/NK6xr25GNh3UPlIaHYsqsXkIeuNsPE6srUFQpacIBppcW39IFS9Hl
vIsjuiiCA0cu+DvEkxFeGYNQyzRCKYgd/lGOA+2GmY7U3Y/dHfGCAZfLpIVftcZj
KvpPPsXTim9wxgWAX1VWVykLuHLv5JioU4ujuY97aM15gRLOQQLCvmBHtXFcpOZq
19CjzdqxrWXci0ss8R4NUeYcmzwgKnD6sUIVTHUHnze5l9FRiihfy4VHGVxASsb0
HtV7hOplMF9vanjQVecF6Kst66M5cg2lJHt29IiPHF7UbSbQIl4l1r6xgU9CPqEq
MEJetqo1I4Ie+PQu1UmDw/An4VjzI18l6YKNM/g82sKlaT45c0SI5tOWQzcksLZH
35vrioTOn8pVbmDYiFQ16kN4vdHRh742rZLansffeTL7EHktLUpBdW3CALtaA5h1
ATxFg8zwsXxmgFKk2hra1GszRaYTl0gdmXS/Y0wwdwkpYiDMNP3evr2O+7uONY3p
6aKKsGIe91hU8YCisstS56BTUjmy+hyL9RnIjtnp994nKdwJWxgNwpwIqDrXs2vq
FP2JcyVOwimSWS/gYZDesdxW4RCtLl/8zAeVbRkQ3dkE6oYm+UuSY3e5Z6vQrtgP
a8MDCnUeK/xH2TCKWXic7wfwdN08TWmJ8+Ru+KUqBRIkaBiREIAI9a3+Wu05wBDo
tscI76YbIBQyIT+GuWV2u2ne6B+5yIPJNtx/Qb29XG8iDkkfQSIaCQerqbwR2FhG
zKZkT4JNm5S2YlvqAvkTdk5Iw340UL8eCaNlQpUpfuyHGx2C0U0HGoeCqq2IY5/h
6Avx8He7UwOEWsAE0LKjxD8msAlLy7A7lCjJSVXUwbF9qUXTGZAyp0Nn0weWBT98
slA2aCUNqlsyup+UeHsc27nhlKpFH4yVXkZzddB65HrNiW8LgbcYqkx6QrkbHpUU
T3vr3fteoaJnmZ6ZWnmaVXFCngXv8VJdjCL9aMbBL1VKhHvt2Dr+0ygQdnF/lSSo
VHCAQDxEDr1raU2jbhlZU9fk2oz7SbCeQQ2CTlH4Jon1BTM6VPWRvLuXY/Uw/Y8V
it7NWWACEE80SmDb8IOBQVPCWs01He15r3YFzqBAG5CnY7V7OOGvAF5XriWcbqLS
c99Vsp5ozsVxKBy1tX4cbm0qLo5Yr9AkAYk7PfB1RT+p30H3Ztl3s7/KgVFjOeEk
AoR2KxQIKWxjmh1arbOJpbI1IR1kazTu08YTYtJA5YPd5XaYMctP/spZv9Ne2Fh3
XV+U+lhAfAGcGc/ces5IZb7d9nt/thdDkPSH/LNRKXG7n3IoKiftNrHp4H/S+LU/
3bpKqP5+WFJL+1ToszAIHyGCIKjwD8YZKadFELo/N9peDWKt+StDkE3wiE26loNV
1/SnLly/b6pZRmO8WVlxQL3nMimwMvjxk8Xnvxaoa2XkJyOEHOWFNkg4V5L/9KSg
yRgKjvU5lTmJibpUlWV9AOhvz+GViNfhzAflAuGMxCbP+AhFnCie+7LpZfzviXhx
53qUiGZAv/+haqo6uUX6hrHbqD+tjNQ7pUAh0cC9vPPif0wmn0c0lLb9A30brjWS
xpnNUVoWH5Nx0urtTxIf+SWpHm6lSwU60Ke1OHAmHMpVa/8co+b5cA2QDyR/Gc5Q
iO82ff5VZLLCALKXaYm82K1YLMCH9vrAUe5cxfdoQzG0XGHCY4iOlDndeSYojt/+
34iE3YGodUvklg//Ce2HGtzdisEXdcn3F3BT2QbJlPC2/0IFPm0J7yVkrV2PPb/n
1eLLJRhse9/ZQG1rs2Soawn5V7+bORjj9rR+dwnzB7RpWLQJslcr2kJXVwbkyQ9+
+ASfH9+75wFJBnqy9mTvKqJCkwCGqmGsBSK+aI8GKLv5I8LK+K0OckK4AHg/hF90
RYCRDYZLtaww8F5xFHDgQhvrJoh7ZODGxxUMgVNiTfrIvUC6Nrjh5T9rPPQsxql5
qDtbAEFM78hz24caZ9ZE99ynNGbIvMm3h3I3quKMEpl3KlPrNiZrPwGvk1YkDJfr
kC9pOJiD9zonuCzJ7CKQ+jvxwLDrytjyIPPCayhwt44z+xUv0xnrqLr6wWDlw9RN
C6lz+9ssyhcK1bUa8agL7N2wqVvr5pzEkC7SWuzaQVWQdVvnWSaIpYMIGeu1Q7P4
/edBprxRvycn7IyI6uhvfK1ggqfRch2eLj8V2R+Mf9wSkt5G8a8QkS8/EKQMBvLu
XgsVbMIUyPLtoBPaG9aIhqjK+who/kmX/bnXJl7+H0xSd4Wo98tSAqBZAqS8wbXr
mrYJbXriyeo3PWorp5XhJcDaZ6G6u4LKE8JtJQ8TF8RVWp7Z9NufOLLUaJfLkqUs
1cj2xFT6MOU+oek47ZCRxBbhfhMfGeMnkRytx2brYCJwcQgn1mEfinEoj/nteEjE
h9muSViQNlYzKMQXZyAnyOv4d9xmBOjWreccfyj2VbHXx5iQbWyKBkKB2VG8UWYs
B6Ha1WhZ6+Cg6l3Pa149nRAphmtglwk8MrjCeRA5kz9BnnWsaxvvlSpr0C3sWU2h
h1af6EtzPjfW2u4x50rpvpRbiLdjaiWu5f6Javuv/aVkHtSTHy9xn5FJSDYbuQbC
EdyLJWKmWivlXTQYQiO0qJVH3at8SlcVY+PkELVB1Gu3sa+iKWJVcEuHzsPwaRuj
lHL9dpJ3bIBciCvdJzDsI0V+o4o6kbiLpdstTEgvNfs3hKBjv0uDDzVh1iqj492E
n+sol6sg4Ee9534kk09S3TztqcoSstc/HSJq5jnaG7LL9J65lgiMtInpCcE6j9zK
0FkPwUhAXOL0WvfVRgUrlGgp2oZj98CZY42+5bScp+EluIVcutBa2Xct7kb4C9yd
qdBjiNuZ3XSQsrjuYAC/5hq3n9pr9olmTteD6TU4ztJjJSKOjfSvZjY53hdtpQrU
ssD4YRsDCSGAVTLfAR5OEuMm85ZwhefcPIroH+uPNZ5V6BRGKhgOQXRyCZsj8RsO
BwYsefQ4Vxhr2e5EAvCbeoZPssOkqt1+4hQ71ENvELThAz1jgzUF+5xaKbyBMjal
bhROW7/GZBp0ZD12It+3WImArRS0sAtMP4UQRL75He/ZfnXctEmR9NM+9mvxqbmy
7buwC1hM+rc4df8sGmdVc5sJ2Eq9Lv3IFKDvH0rkRIarEqZjRwNhrq31+J/EOdkO
FsZGyzMDZI25LNRDBksoPQU+MTFOkPDn1b2u0UpJtCpbFQzH4HjEU+vBICK27ic7
yybZh/NkaEtrz/zZcNX77CaTnqZiyyU8Fbi1wSNUpVcnTdmuwPEjh6w4KDVXglb2
XD7JNmX+5YFZ0jV1mDEHaI0ZxuvV1KJPRggDb+tNPJqjT4bz5PmwNfjs+ykT6Yku
/nJ58nDy0PNk0x/THP0i/xYshI0xGy3Ddy32ZZcMIKXFuFfvb3LkoaZP5BhyKIrY
ijvFPJusf5qDhB6g7FxknzJ3QRvdo1wbLcbbzsXwVIjDmyRgd6zAILDhU6NusipX
JoEE3d4xiZDm7NHRCvGbSES1cmuxpomAEBrDHEsV1jMdoUaOR9TYzZW1i+fckz4r
jnt70NPKww7YSyMB1EsG6RwSKOeh3m+7fE3LDVqrg7TnBTiyHbuiHUMAOYn4MNld
PiYeRYxvaXFECe4CiHN0LkKpvCoSAaSzyKw7Pwtt+bXd5JH5zOkwPRP6IKNZggK8
dSEI9iEVDNcVPG4dTfqbQUVPfQZ+q6VHtM09wD2GPoJvxaLlGRMouFtNNtgc16mW
XjIEyxIKl8HQaeQyMxoJ3B7rGmp/XrLJ8aP+SvQgv2wEb5He7z0mzp0L0+Bd1U+K
SwtTm3GNhDGntOAjI3GlANnjOLo71s3eL6jr3u7SpB6/jtiLRlbPdUzZfeyUg5jz
UqnAMSGyB610dNRSflwAxNJOIz6mIR1ALAW2jXMdvae6lOsmPOwIWDndBLK3+9x9
fy/XDAk3ZqPfAYkZDf5bj86FdG4usJkyuWL4aiEnwCU8I2sKR+BN0RYmpNJZ4IsQ
9rqQHOoMAw84r1pfBbzUf7G2WOOObFIBL5F9CAXIWp6NfQ/d5p8bCOwdFdAVTMA+
+4plcuzhVIrqI/cvqimWsCPvxv+3wVtvxXmZbTKrCAbDjWt08Swk+mu8MQc5SY5k
bPO1COp5ZRhADpgELwJk6RPcm1ZRCkLR3slXc7lgvIV4f0smtGkpB4df4Hlvh+pk
pEkEoB4VJl8UH/NNV6UNaIWDrN390h5YQHC4egSoMD4FVkvt6m6nlr5eNOo+ebCc
auEdzel0Rhvp5lTysq9ggj4J8m+mthYpPkMyZsQi04SRQe2WMdsRzjjv657+DVgV
4Ocm/uuXzGlbBQgqSydg8BtvpKsh4/2ijl6YXDOH6j1pjCPqmKvIFfS0Z+TIIiRr
12XGs/k0ULUCQTjTJol4HHVkhF57x4Dh0+IXM5phDqeVXMGlkZEgWfqEx/wNdbuN
FkNxawLdrZiY6VEAOizdKLGQywyUB3qe6utUnZmLwC7siDSsexkK+uReNhsIkpPK
Vi38i7yCF6hlLLOqeFzR9lThH5+WnHahyAHCgEUznWhPbDKQMBxZej0VxHoKGZbG
+Nd/VNDw1FQzPRtZs77UCtpxJpnHdr4/tjCE1AQxC+Ld/zdvi+GU1mo72x1x1DWQ
mpblzLXcOxXH4Qn5W3kHC+nYIwJvtWjiiccxd08IJPJXxWmULNMy/3YZam/k3/bq
zorVhmzL39miIC3UlBvhx/qezu/kGYGTq/YVMJ9hsFuKuM26pmfXmc5Wwzg2LJ71
ACpg2Q0DnTXZ7ZeNMAsgBJqdN4NbNDsZsU+BzdQmjrAS1vPnkQUR0198vPgh8y4g
kPuKgIJaPtPciwZrY9FbuPTSxv9Wa8pCNXdOrLAqJV9hFXr7eD71Ai89k0kLsxWd
l/ssUJU/PYsJJHdL9KP7g35X0UfvNnhTZUxtPCLL1y0uAcre8/mjEkFtksSVNfdp
Vfk8yWlVyPAw9ourWZgNSl0CnkdBm9IK0yWZzG4+AGoPngDMjpj3dp8FmWbJgJ5M
oswBuqeeUsLjMBvc6owSwJ/nWVnItZbnnSqaYHTBqEeNIdGPwy3+htYjdoz4n2/q
bhMOLppxaZJ5Ew0It7gPkVTLGlPAA48R5Rn4zblaDlHvmpdhPoUli5eX4WbAHM53
8gfgUIdyIhvkzHMnIeekpVB2cG4LnNiRW31EIryPm3Gtw4PivgcMJKQek+K4LesP
N2XORoUkQIZiCg0GDdwy4ak97+CaSxEEUh5TIL53sHHZGRy1J0QwBOugPI/UnGcU
UDtvIWyrSLKFyi9zqPCPYeRhjn/E/A/aym8Lc81NhQdg2CDDcBHGyCRnIlwhKuEM
kUXqd5iewty7iOnUOPmxOsCSaaPBzNjlgzUdndi0MKYevuvBfTTfJtyVp/m3t7Dk
VDere4vllBkUFAPZLk/RBEynydx5IeYQeVWaPClWuwOms6t7D6JHnyyS+4WGbhxi
Cr7/gFT7yI/cvW/eNsNjGhEWlETMymVbHVSlhXl8F+ENMVBxPm+DEveAtKYPPuZN
4agrMNhNZXEhxWOYvtgOsHSGj/wA2nfSzGS6NP314ltHJ+rIfhSw/apd7u4TrP0q
gU3i/JMRChV+s57hkuE6eXMw5cXCOENDfV+JNbpK7t8f8QTqd4ye3SlZp8AzNOYZ
ilWayxr4B66iSjvJCQBbNgcfCyVMqhfj9p0nsEysHJrPbtQit92kxXkelR65IKi4
DLIRuPb8/S+sYIcPuFJ4AvK2MrYmg9SgyFYrK3YkkRwoedKMgPC9OCxL3JNndcz0
Iwiyl00Jm3LoxpmjnUr5KmKMIhqxpUhXHIsFC4sXO5I5M26/zMsKhI6Z5I0DCK0P
78xOej4V8JEG5Kb6dYh+WUYOLkL5QMUwXJifOcr+L6afwbIOIPG9FnJFY1fxqL2c
apmr9pxa4sRljMCJuS6kpxcChPcDu/grhEiRpDFuDSqETtLjK+bYPS/CYf20ZMMQ
iQyixE+/FQ6H8jD5KJ4p2qibLiw5pmSp6lJ2m0GODnkiSOuYyH7AyZ5mbjJWgE9s
puQapBKZtfbgEYSbX3qSrZ+GZDdCwD+tRgJELJtFr0M1HI6KTbNZ+wazUUYWD7iU
IWNcA9UgPJQf+JFfeMeK87G/yiZ4HhmlTXvSW8ln7gZfcf3BPJS8QiTP2qKadPxI
MyL/iusBBoe+mNtyPywIW0ROxhuZSIN72P3m5yWPQWExYa1r4i4NhBfkqzaRq+Rg
ArB4u+mf5wl9YHfFziz56hGB0+iqhZ7rGUnYhbURv3vFUQayCXLWGZV6nNswYPWW
wWXUnjIktW3nJYGiG85ctsKLZliEcsqyKBlaqVpok2DS01yJ7zXvcR8V1CzD8LWO
+Sqlbkblh9B7Fo3YGWvEZGs+1jUAtFEuV5GGS1/JPW5q6jodXMhY+PPYvTHFAnKg
yE2ahFP6RRG7mLPUmIhjUTRvBFVjxfWnHjOjpdo2iGRB8ajAzmonsh0CHds93W05
yXTISleVgReIYdQBFDsYTmpQDmxqIXNjOh2iRBEMD8njf0fVCPJd66NtITsd0mV+
E201q+Ve/R06AMTE6HRQC1qJEJaeuaQp1yHZvI/7U8tumo301NrhINBWlwFztaSU
Xx/UrLZ1pzUtDFZIkE1LDIOmqouGgwg3h+idP1Lh8VIYXTOIbA3ZeMMcNbwI4/nq
R+DQ7jDVLbOcEc4aziYed4PAAv+1/i3Jz5cSvOaK9bHf7OO6jM/kRzdrWRfPmvv1
oE8zuw3RylmHtC2nFq7XA5a7+6r3UtPE7six+Kc27gfWQDaSu9Gol7J7uJUPS2nx
FaxT+Ep8JnHxGN7mlvj2/MYw67MEwofl6VkGOX5Qw5qI9FUM4fovsMlWwpzvLht1
5lwlJOsvMTp9EAUDt3o4w7KNM8UexgJJU/U2jvoKVg1VhOu1aR7OnCL4qZAiMAw6
DVo963Fi8AK7E4EUKdi1RypJDWu2Cpbx2pMOdByEzgAsP8cBZKw6DmYUrHjtdQEr
a4Fg5AW7yrNCPnNnpLkYqfIX/LDDLequaVWyJr2yaiUtDAiU5sdpNLAUSoCefEbf
pGsMri0AOQhJYT/HJyuMNfyhyrb/xvuA7wAxP0or4GqL2bHqMbwCRxyvk2jEfC2p
2YypWXdVEBm2qMbnO0egYr2K6pGXSFLxI3Q76+HqsJH1hMCGpGJxqbvlFDLVJzoo
Wa1+cV6SLMDDFBE+rcNYjT9xnb7cZlYuUkIfjyrBEPg9e/cj8U/8cBIaC4MrcM+j
YKC60lh6TIgnxUBoz/QIGQZ95I3lm3+EhCOnJ7hcnMLwebvQG0AuuBoqelk8zWZ9
de+b2hmYQEt+JsHmgbyxg2IWvlIvxDtqBNRkI1c4yotNNbFNzc1klIrunnGBYgfG
KM+cgVYubeAnzj6hzq27rJ0f7+yaVTOtHHX3eL9OSyaC4qYkfr/BD4Whh0RJHkK+
qvvQsJ11WaiHzNLhY9fJsIQBLlL9itvv7Zby7Ge3IWXMeKSTrJ0JG7fD9Zw89aNW
3flMTHRty5xiS/R3ftbGT9FLn0a/oFW/Mj79Osj5JqmddbRTCktaSpzaX2x3iiHl
uQLQOxh3mw8ClvxbAZMkf8LzcEygmmTvskq83gFef/FORQCZu4VYs/Ere39evyO7
ua+8iR8GnTK2od6Z8FpTkprGA7+kzgbBnw0vgTawLhzyqyiPL/Jg+xFekPN8D6oE
dDiZTCBywE2KkX9CnS7cX6M33hrio3Lor6jxOPlwL3OlHSoZ7baSuR4ovpJdsOFN
6CBKoh3n2lhG8solYK13upKUNe5+abQObbEgc8RVW2xwEQ/ImqWmGqpgUS/qmAa5
/gEH3Ewmx670P+2DLie0TSU8HcBv+yBBzmxGsFk+C9XjnFN4f6m5Q2b8O3A2fmy3
3AI71gxueu1f2E2bV0UWRFHREvy3b+5MDXjiLNNxodlu+fShf4QBBb0mxTKaQDyw
P/rUhFVkdHRYqgxp5BdlzZxIypFT8rn0XMDOJ82wdRYeA8pe3YAafsoLjfRrOW2/
oKIgScAA7qRRMOq7/kiR7uMCwp7CBkcZpKhl3NfcXaFDPOf1xltwOWbuMUDnO/5y
JoMlm32SG3Pae1o2iR2dnJoZCIRjyNscvbODL+TTR+bmbMVrTVad7ewGF+qCoPsy
/1AJ8Z9iklBUZcNdh45xEiiYTv7ustG72KkNaluvTZc4p7sOaLcVM7L2vCHvhTTC
xGq4m/NXesqzsZtnmvozJQIrdPzFq0Wn83wBwupA5aqRY4AIqzmGgoBTmXX83XB3
TKMDgAcP5ZjSeC3Tp9wY4Adpo54TpCe183ToIH0hdLK8tLm8LOfVcpyBl+2Bihc8
7RkrULCx//AFLykbFuOrvKaIrQlT0BYMcjHzJ6MMs9GQFG9bFRzInrnE4fP7do3I
WpfanQU7OiIcY7e+OsOfPE8VZYSAGOLT7/mAYQAi0FpsG65dXdL14g61IEtrQiG+
qR+xR1Xyg742XHhkhZhU9qeIyAg+I+YrHE1m4etWys1hg0T+TX54OE3YHWNvaXhN
Xokr8kQjHQNeeB8HMUAvRh11eNt2/pKjHQ4voEuy2fFFCOYpDK9oTvo3QKpW27SV
ZhGSqGa8q0rv1KTe3c1d460pYAO6pLCtjCyKXDNUFfkwt9laTd9P5Clboe+gS4TL
8TLnJP9iLrqq/7aZPhMyFqzFTzOpr02/MfVvUaRNG9Kb7GsfTNndQhmzn6atwmvb
9N/i3AzgYV83hi8GQ0USr1VSOBp5osBTGXXlRFoYmCOQD0TTHvdcNW4E7TpaDzSo
iiaYMH8Mq1eUDTqF2px8+hrheMga9ekX0Bu2uopTzjcoYy9/Qf2vWw1hIdtespIw
t8im1+jCs7Z7jzywfDWL5ldV5gUs5aJlv8rbXwoJsWO9rZN29mh7f4AndYOytb4v
6GOpyuv1CB5JNLDthUzTJpBbLwzs5Siec5zfmeUGOI7s5kfuuN64AzmLyMufdHlL
VXaKeuV4rKR8nLKmSJCEsLuSjfpHjRS7OKMm8bU+e4/vcFmcm5QmQaXBb8xUQpsV
QmRlytAR9oISbG6exbjGrXMi4txw1WxE92Zsmu0GHqXmA47mz9zVoLb1iu91o3WJ
yPdLGzrZbdgZ3ODDRVvPcBcqzShLhcHSlpyiOlT37WgWbpNwQJbGSHe9+orDOxkV
SVkySnKjY+kTJ/SDAqeBar5aAbY6JbFYAU8282fGV4qqIHA9Xk7pC2a6oxFD3Bss
bCdRBDFuOhadCvlVcpdmT4xf8argyej9vdxC7mBC8LLLQJQoxmaeMq947R3kvsNc
zD48o5LsOvB6GKvCxlR2iMYgZxj9seRYUfwdVMBpTaXcZ3hjL8HCJDhn5GZ5DgO5
r40iZZaV6I9OsNBXk4jnQ76YOFEy/4kq/CE+3Y09iHiV7Gi0j0LAHDDRX1w8Scp3
hCqITe3+ZB7cCsjKmk3mVovrcqkAQjYGTg+bIs6pdOtgEXIkNoSw6IPc5+TIea+f
BRWxlgkioNLNHM3s8jWGhHJ59oYSXXVptRk+EdGnW2khlIiIZMy4kjoIY8BUJAUC
j5QJ5s/tnPDXvluYvqLdtNMYShnPOuCWf5JV348mW0WLmG06rPWI65jrhFj+XeEa
Xq2RA+iboD1y9W/QcngbJT9+uEDQRCVun4a7nnguXv/hUoi82oPvrq7w70GBsLAd
RS2lJ/lt9rYyU/ggaAUx2UJOT2qeGKSkkTc7RqJ7ReGOQaFvbxS/EvdUQF9HdXLO
gL3K/TEzgEbvwWP9+ErFDIr8djpBxJI3KwuvQdHBKrm9yQbk0gskDKtMNeQI+UZ1
oOd7M/bqwrGb3+oVYPfHQMEVeEZA4oywr8KTqafoztYeEm/VaLa/3uM34tETLHp6
frEgIt21YaHjdolik/4Mi3sa98BMeaA8IurJqGix2TCcgaBecYgpD3M8uG7oEyqc
Iz8B5ZfH/wxBb69Rlq7j3IjReII1vTJ4p0pTT16bSot6UVkzGRNjCDhTYuXFjX28
HvHTfl5+ZO+uMPfhgLjcHd/jjWfwEwgP0Eb/reQTA6QXQJU5PTcXH8Qwk8ZJuhG0
qLRdv4NCDgb92XrLGkbdi9/PjH/vfqE1GzjT9Sdnkzi+fRfujAf6bv1yQC/fIpce
DMHwHQm1E82eBicKBjErWfkO6OuxUf3fYDfChhS3ZSpzSTnl3IS+/KzlMVnxfyHO
XQjBcDnoz04Tlm3el7jI68NZ6JPo4xU8Rx60cmGLnwqVyTFXnc7+/1GchZ7yv0rS
DfD0ZXcBFwCuHbt1Yz/bJRCv/E0t5qsZU9Y0kOGoBPiK6W2SmzLCaTP3sHlMQbOI
KmTeUZRUAb1mvYpbRqKs1xoublPMqigvKvfBIM4tUJlpOH+Kt5p4TzBll3WNmOFO
WRIm3+0qK+rIO2JDPRFofIo5EAoSMvHhHQp8P5PRVhoAjGCr19XdeP12sszKt2Zs
zB4UbFZABV1cJxKG3TjPM7XHZyZWy3PVu6EyN3kbAA/PKpEKnz+XN98Wb28gDvXm
YU5bH4iA53qJXVhlhragOwLIda2cMXcoqvhJcgsJpDly/HEBjlOoTKD6cv88G16w
zuvLJfR4TKcL2UGq5iS9H8kKgTTKhbLz1V2/5WkebKyPBN1KXbsPKTA4ynuyIB9P
xn4Nxak83YG3/YCrDFDxnA8QMNA4mKTsdrGrVPX0S8DRAYIh8wq4F3nlxD6Sk8Dk
cAAb7rPHZ66ahHm1DiBgCpQDkBE2XRpHgFvPT46f+i/S7rlx5104A8lYMJ8iwOBO
ZOa2aM/zzLGB8NzFY1F94E67vva/+6gvjGK1/8VDtCUy0xe/JJx4IrbvP1PWa8ac
SEbg4KcrVelqIXjYZGgrnxXAz+vCMOHLLx29OfI1f2+ooUwzaD9jbPnuiSmwvUr8
84N/+EaYVJDa65B3Isd75qLcb23MG9W/K763pIRIapfiTRRJpUf+AUsY3O6ih0Dm
kYmiI5jv2FKCZwhKXYF6cR1KOz9Cj5p7lc+GEP9KG4MhG6qj4yql1rwl7yrJqwC5
a2V68T9nDb8B0XKQyYQoPo0bc+3oIKNogqqsn8yLM0Sv86pxvKKGMZ+/GOqTH7fv
njuQWQokNBJ17SlOBmqsik9BqvlOgwKqR5BDjkZiK8p3pCzfAeiagcnutalMXqBI
or/UuT1Nn2+12DsCjncL1aLtjhCBYiPYK2nB1npOEhuwxpxBAbOH7PdO5o53Mjom
m5L2vq6BRQLCW9f/K3t0HtIjItvQlLkCl/WAQbC1/cH1tRUpJjKcpFwJQqgoIJnr
H2nbC6zL9SHe7vVDfrAtZx5tjfhGYEwRYTQSFNAVQzX8EqeMMyRjZYN/PA9l+W4O
x9xelpALGi/04hDziHA5RbswpP6YpStHijAcWbfzmkNYi+NvLE15msvVz87n2eDU
MtHH7eJ5MF+T8gX07E5m8KP1Zr3+BDJZMiyb7fmcRgD4qCG+HAyHRjtM3TJc/sM6
0kBNEBCkVPaVwC94ccbYRZ/Ml8zO4p/yRSwc1lBmdcsuv3NGx4jQFrAa9Y9wTr+X
Kuxa1snzE/9H+PJ5dzWMa23lTddI3T2iO8rCX2N/jhff3xcUg2InNf6fSUfSNuF+
TO0BH58mXHLk9pi+tqXR5VAwnJwab+j4KesW8TZ8y2XhwtoCLXrkF7XOq9N/F1dU
INopywzigtWLkBbX8OodhydX0ecbM4Blvi9ZhuOKFBcSsR8K+zPA3Kd9LIGWj8/J
/EoyjWfiwwP3N1YkmxOuFnn+WQMOVYgKoNT+1Gowy6Z2/u8i8u4ZF2bkQwunsSdC
pNqyW+G4zpLX9oHrqAG8kf3oJfCgVqhwKtW9+RgAZWW4p5zvMgjrICFkg/5LXmll
PNDMxSo4b8oSut2CPty1AqthyJOkimY9lAqk6Q1YyUQ6o0hnL0r7Ltm1aOwYOwIp
rOY466BIlAzuIqewXY5UGT+5O+LSJ9STobkwyakjeoUmoWLH/OENeWkogLOaFxyx
n94Ly1jtk2VPerG0gn8onCcjxGnAKsI7+9BVMF89ygwie9tqgmz0h/0tSSxVWwL4
DS8gR5eHcc7jIfwb2omfx0vtaRYLdS6pyUun/lCHdKipSEXwIdI6oOY5Vdq0OUy6
qYlhrzbTihStKinRe4/HIl031Ik5NujOuIRNOdJ+pIajp4eaQ1sz9ovoUKfL43iu
4XDlfQP5YuoyjUoDb5tuFw==
`pragma protect end_protected
