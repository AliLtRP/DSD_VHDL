// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:15 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
P9mufEZu16D11gUHzADDUSEwPWbQ9I5w1EOApVUxT++gNFCtIY9V3ocRoUHQRYOL
dynV1CxSoAK88EjP3ix8tpNnSoWzrduoeECMmsm5yX4An0wcSRftMsfAjHTrUCff
bfjzYnLPqJpb1QxCTAFweBIFWGwuN9J9GkxFVQhFIy8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28864)
txo7zbXbUBqbI+0ZlJOqZYq0gM3jqnv/xS+T8TWmkC5gSA1atF6uTFVkHHQbCJwi
pR9DZ0j8cPJHwU6HGtQe1OSw1RSzdAA2J19FcsNJd1P40eI+dww3nWOd64GHasCh
KZ1NzrNDBbGz9LMIZEjQB95phtS9M3g7R19QHixoVW9A4ICDlBJJbfqZEvwFN+Rp
TKl9ICz9peLLZxsaA7LRZ5QYJRR2gZSTGsI+XX3FD6eJMt5fesbsC7G3WhQ7pbsC
5BfkPt8mPr4fKHt83AOfUzsUN4ensa6lWU8gbrYjFAv5zJ+bawVIiWBdFK11X1wE
3fHMqZxMakm2wboOA83gmQid3loSZHXrSwQnftHgphVY5MZ7cuwOd8NNzIpoeGpS
8VG3xMvaxR15Zn1To0twdHVnYQhiaftFWRwCvCzqRRL1Ctlc7ksyEtdqRNF11b9/
pkKD0LDtoEJ6JdZIve+QF0zff+wPre0F0BX3buFhYGOZVPC6rZ90+MVWDqsqB4Yo
FOxZP6JBDdwHQqUgzPAG9YxQeLgq51iDv6MdEvEFOgXuGeOeuRX3+EM2/vYymyHP
n7u78vTwiDqEJ0YQulreQ0i5FSwyU0A+RGRjiKvK9+jFOTdi9hwbvPDsPegyjhqW
MZvn6daf5hme4fy7q+Ah9W92cYJux+m5TNruk58tX0MJlFzHVPtCTkFdsESB0Dub
t99KL84UoSuIyI3r7wN9cqoxCWBElqtufUmy7zDiRayxZ9hfWtmkBvkUolNqKplF
a/iYLdPrOwKZJcw3UNGBnbeOZVCCjHiZwgjuN3TkBHCP7DOvKXEziaeyGJO9XESH
SqXWyiGBistHDJl/HytRxSGZH6GnNPFOb1JJxU6S7rQW0RGNve6pYKEXNjdFBWzH
BM9sYirzLsva+FQ5UAIghG2I/IysXeXD+iPhUEQjzJCHQ463L0+iYXszh3DYI6+1
Veocev1kUhqjc6BJX0MtZU7Ghd0noGjQuQGn/BjJIiM9JsPJRIPJBckWgB8iA1gm
+JvEHWM+CEBRh8eYmKcN6YidIzZYNFnsNqTxR97JArK9khxgkoGeWFi1vor7vyUd
Pei/Yoco9WvjNM7Sac/gvrzytUW1lOPwUOVmDwkyh8lb41Kcp8vWDfLm0JcXWa1I
xzMRz10n7WtD3rIqvz6EFys+L8QD6H2VrYWcK+/u5bPjUa3qqKubMZf96DTNdwia
eoQ+fHd/L9ryO1+sE2mHaPjM2TaYk7goRhFYlKEvpiilNcVFR5LqAp8GJm9J9YLO
dYYSNlyinOpkC3vXVVHqbgZwPWp1Tbb8UhFd/1eFkzMgFa/fV03VNkFpKt4Swf04
Ls27arFmsKJtbx4dkQTIBJW6IZeH0OWRP27S8Hm80g1pNkzwHyW0DofaQOQm5d9E
U18zsdaU+gd3BOeTjoePtVTFM28tkTfbXRXz8gjkQYB8f3b4SfuipLdONIEnP0Ik
0uYPwFLuJpKN2/kn5t3RG0oCW6rt/2mul7BrJ85blZcz4pATZvqJkKGkKAy3Z6QT
c8s2ZeIRYFCItNRz1Fqr0Q2CE5EK/izgDI5q5sC8ho4oP6XURiSddbprl/j5gUks
PTWWeyTtaFBGlS38hnx9iVNBk0I01Jy0FzmofnrZrwylzhpUFzqXGIjFyJSC4Evx
Xjx5Err5qx4JZAH7ns6uLTWCgXouAYXBCBTUUqCVkq5geJcaU3LbRi+zpAJ8CItf
yCSPs/0NOvf5GECo7lXZiOYQNKGfeMO903V+Up6d/T5bLwyP7AgBHdJWXlMQQdR+
LfhpZ7NPaGYg/F1+gkbbUXBV0trAm8SWV785XYXBAtu1EMHyxZIU8HUIBaRg80BJ
VpxLTZZCRKNSVvKGMCVs5QiWdMQHEfMiy31v1TbkDooVNANMIzvSUE9cz2M2n1Rn
gqbOiHF/dEc8s5bxJ1pKHPYzBQx7GGXDOs7O+FSxYFAgtN0fgg0r76xhgOcjFYAv
fty2N70Tgy4og5beD4Vyj7oWxY33OoiwmEmsBAPQYmdBDDUrALpIkGJGMsdSQDs2
7wrKR1BgCgjtsesC7ol6TdYeMZJjsSbR+Uu0fqoGzfr9fImQbS/CbXeB1awP/DF7
KUQaTAWqx73xUP2nfHiVXypxqrbGISH2ZC+EgYPBMX47G1GXVUO7fLKd92/DSUVP
/VrFWXbJHtLTR/GzQ5nveUucC9K4kLx7pgBiki3Xxpv1gnQayvE3Ot3XKoHVcQR+
7uQC9+qiPNYBYjJQ0es/Qoo0jAhGStE5HyxpjgFTwU+MD+w6IIAI0o7VQRRVWpiX
uA8E8vhR6ehPGbVSPyv6DflRA4AnPNAzzurbAgZrSyDKcWDeRO0/W8tKa6fZmDbW
eo3F5laEaoNKYfc82mTI1hCKq7m1kfgH2shXw0PAADvhzbtv7ccrKfP9zzQ2m0EJ
hhN03S3H5ILKhu9lxwhMgGUQqDJL85BGk8WTu8Flk6ymF8R6ohftBgmVqbGjL4iM
WEycI2Bm7ujGbhAmWSqDEsBB2T6z/99CMWUAYYeRKGgguBTwa9SgowYG7+JJFlOe
9PB+tQpm3lhRs8HS+16RDkbRBhbq/PSpOjwtZJWhtlZNa2f8YqIHj6HlnXBxjYtw
r76cudWpBiBXXuSBrx2e+Ra0c2PpFTmi7zqZmVGGgSxnhTGegXW4WVHn+z3dIcpY
9jaPn/yKMucjE0gSEtf/BxsQui8rzmyxEme14hLOtAX530CM4qo50U7d6rt1QMtq
x8f+HGWERgOhnIvRZojRHSIKrU2lBNy/oHuvWcGrwunAA9EkYO/1Cue3pYKyixZJ
n8vbiKX5sgYCyDReNjGKZJkyVrBYDjMb06hKzs7kQU3R6U6+wSmbuRYYkLzCE42e
l+Ds+5X1uDTUquW4O+FJHj4ViR1G4HrPnCdw8NOx7p4aTEj24shEoUM0NJl0pCLs
W0VrB38i6J1pCOD60c9D2QxX9U4XVp+7QneZR3Ju9Gm/LlCmLqE9KAqK9pTGo1ko
oMZUjFTNMqaFIiGSDU4clwGR6YivLIp6bY79QoGjVy7VMIzld3K92hRW106w8bQg
+SGVY1QdKil/UMsM++5IWRja50bDfgYb8Y09xEfGik47VZ+HPrBr+NFXdtBH4Ws4
WhtOdphaPehgurAEMlZYIuIR7R81TREnMdLGfwd9qBK/h9NVpBBT6gB7rtRtjkzk
xnKiYqRiCCUdm22aLjNk4CzBHbelYzCUe3vWkzqxxZ7eWuyIJ7mlwgfQhwZ5Shup
lUqgosPBWR41it6yoKqJ8ciYt8QUqYtvOSA8L7L8O0fSK/wzah5aoPpd26BGUUIj
y5vjcZ4LFhhf9w6kGwqstJIAQLoREf/GRL815APW2EwtDTI8eXgxfuBkl4HhJGKH
oycJHOTlv5krHNcaaesAM5ruZLr/OjwIL8s8Tm3hNqiN812RVyl7M9R9lhQZX8BB
bRjApUgxNBR2gAb/EoqYK1Q+DwTUv2lZ+FCPHK0lNW4fvcpyspk05QFezGfP96li
eav5r7sE3Et1yJ/aQ2iVDvSdF4ttsHZnpRReE1+BBpIwQvS1n9dkWd5/RFLJ3iFg
szyQRQMPASNLUfnU7JTWUifV3mGFWrFKhwl1X23SdR0JxHKs0HiqV9RU0VH6aXRp
+ba5ZFy2XRzWGwV+C4bJvun1+t3qa0mBO7+7ggWVqzlsPu8f8F6N/Be6ginnjb4z
UltTCxSiuSRDnRClF0QlrJSLceHWwhEcPnioKldu4AR/daLsQRum1yMhNLtLAT+v
WbzI7b6Xdek/FzKQeEvBooCr4sLtWjCv3iZ7Yfpv8tfVlL62GgQ/wWP+6jB4DGcD
fRcmSd1fYSMlJP2/7DLlJV9UU+tTZQiqDNhY65Vg/ijF5NY/MWMbLLa1G7BQw2f2
GKhAUzlFUso/RzUSHnULm6bxNsWg+8T4MpThUUZ/MQvPcg1iV6oD7jxlr4hwHk06
hgK+WV8AjxB/Oq+lqyoJeOEgFEK9GYzoiKAGDD3l8JqCF+MLQZe8ZW3E/laUpFSB
lx0uUUbSUccI3ZO3eKVnWgomTOsH8E79wyEBWEkcaaHeCwrMGgyKeebC67LcX4jD
ljHrMhusxtOl8RbcjdBE9aCQSkAlVSV7sFxDOWPQgfdYKPyBEvZ6z+iLZC2t63qk
yZhnyL9mNAFHSYhh+qVLmm9ck+P7+cOOEBtEsPnKL9UGwGx77pSrT04sfiUq2n76
gMZn2xHkoWQqetv/+0LA8tYqQdR44w4HQo49rI5uIdWGV/Jav2Ehx9Q9FdfKtgoC
eLRabM09dbrsRlXSl1XyKbCDaB4xNu6l4s0Ykt+IcUJegILI2ncG+YUA35qkAUcZ
8ufI2kEiIldlId4O9LaZAwyJp6l3FmfDz+aluu+IYuI5jcRnS6wcBNcBO7mt9ivW
YBRhmIRHqgX0oqfxepECj2M7lJvU1x0Jtw1PIEtwZyTxBtAFnQ7EAFog6mZMbmLK
ElpQauDHSwmb+SGNSBy9qR7ILEwMGjENrkxKzci3cSsaeIKEsI/LPF9KIon2Sq+Q
l2bAaOnS87fY4AV3eR5/q4frfIbNeu3IXk/B+U/ooEhAQCjhhoTOculQTF+2+9Qq
0PLXBSUB+ekXSr3wEWHAh5OaR3FTq+B8sYeyqpzlKMAIaq4GvO1y1SSZnlhRroS0
FjEoDSbzPJm3Oy1d2SdQIVR/h6TjQTTG+AwX3g5O3uaO06SSPXxggoR0t/O3f4k4
ayKFER1oSC1YJ/+0gMOkrV0FON/ybuBpLsy76Hi+CG0nSm1s0K7NrpdjJNMybDUC
UOoDueNcA1nf7tvlmOVqHWTSIUH2l90VCoRrCTntR3A44wt4xJ2Dg/LyHNdcVRX7
IzXgpdaghRGfXcSmGA29JVp5NDW7LN/vSg9JdJE/idPcX5nFBrU/QJwIkoF3hmZF
UP2PR0rKYBC9auztNOGSKXLG1+mY3sy78ttf6tnh9NShCfhLMY3elIKSkFiPEVSk
3FNbpAwpa5tt/e5bosGrGbM8P5e7POPxeM+pq3GAppuMKdP/vM5uX/MJ876ZHROq
YJZOfIxNAoR+Wql+NdK4eBrDE8VTnu+Jcp0CaVs8Kvv+l94a/6fUYO9fWq38Y3j3
/TNZyrDCco3CyiNMqyEBlUJHDrCdj84AkqKyiEZSA56OINoXxm2dbT8dP7ZaSa+s
jKEeTonvkGecj5gD3hMOMbPp3v+ky4EQJ0vVdhk4hgdF1URt92Rr27ZlQ/y3R7J7
GsgnAmcDrczYsfD4cPvSK2aK/EtZ1bIqytRgXGSrYgs0oaiSQzcvqVcrwGJE6+2y
WPZs2EhjqfdzSqaL95zXUjM/ING1wQQHMxB9VGer+KTC5+yS3UEp17/i7wpVvGGu
EYPFgV0XPmWavcYoASFxtAeNwap6cXwcErFbzdkvcIPWFj7Nh+EoHovZwfRuhWDB
ygkTK7AphEgXVIGBH+8Ba7E5YJrvBgnouw74nnrWQf/qQh45Sl11Gd2W18gynzM+
Sa0RyzVGBWj/9qFWWx34+xp7VB3Q3JDWnyg2o3GN1ou+Yyyz1aKKFQB+AGjXwP+d
lGNuiDdYNcq2Nq6IPwCRIzwLJUBYkrPhEIHve5UJzdL2MiEWi6pJbTF5HMW3A4hS
VCtgW2nrN2DDeFwBCjzkFAYV+0hsdY520h+V58X6P3kRrd3NUZRCkvF3piKcCz43
kpwJYB104T5DUr3/eNR6XKGy0lbE+sgKffMyBbGFSRHWkZ3xIaGS36nlNB4u0IcS
o529rTgLiaf6epUDRIj/sXDcogtLiwkjP0zNRd2BWOv4+jOBMYmNFxYbBcGGvv/A
JI09SqnG2XuCoB0NS5A3eF+UZ2hhVBfAMoHDAc/TAT3P+JB0KlUvKCEkI4N9zxpe
BLNNdDyX7JckIXsbBSGrX6oLY7ST8mSj2NNtGGkQu7JdjH/cm9lm1vlpZapgREVv
qmIlufcaBdhhvi+4IFmoMZWea//ypbzFFdKZtkszZHYzb0vj33+HJ/1r+Yp+PV4h
013XFHGthEakEfMqZ1X3MGPRx1O954gC1PxgUF4gUZDUNgQU8mQ5CHUsbxCdcApK
8rM+MbUBxWI+eq02DtBKD7H20XdW7cNwcVcQajwMRlPNLbdMpiWfZRpD4hvkHTDm
lIiUTM9xid8o0oW6bDf8NQkxz2/32S+w2GkYYWRND+qLiaMmYzH1zBoMcn+uZMtI
gNXe+dH37xV4XjaF7iGUxyz2qBX2k9CeGoZ3keOiHr25CTCh7+sS8cYiEYJ2/6eB
NpwcwjjdaKb9iLMsJu31OIf6coNVGFBCkMq3BjzqkoDUhKSRfXw1dsuFncoV8976
z+Z4GQb3anyamil+WnmjwfCrWFfaFbPQ7m6qYAsYU2U/j4guoutKW8X2XP1x9CUJ
dzUkMsgBVOoCJFZH0qc5ULbrZP6AuaYyXiy+oqIY3PmsHmRro1h9z8PPq56EXE+k
LM91uo/LrsjGAsuAQN6/ZT272ZjzdDumGqq2eMkyrBU59NTVTExLRgEFt+7O1sxC
lgZGdPMDOlSBYge3RJLUnFXUuPJmu85FtYs//Qc2wyNLOI4+hBu2KRVJ6RRxRyWc
tLMlpabU1DveFBU+lugosPsPLOy7NQjbWOMSI5Od9VoZDzdqfZlRngTIQKYN1JdK
ghHl5dFeBtB9CJw4k/8IJOBneGE9B36pEch3hCuZ3fQaRHsAE28vWX71hccnr82P
7cNO86CKiuPK/QgPJUTWwEEcGrUE9Y+s5ea0OgvtXqGiMI1JLM5/fmYjYWBAWM5V
8+1NvRobAVdblgWSbS2aYXnZBwArbGyh9aXJJb2V5+ovt5c48mhJ47ynw+rGtX7w
1jqyxFolLdwNrC+aVUNxZUxdS8v/wsmpAG0L0Xj/yMwYPfy2q//xsPho4bumCjVc
7BKfOfIXPk87xuTZ2fAOZ2uUlQSTFPK0bgbLujgE4a4vIzPR/TtUtq4n9L1JY0R8
V+lFVTx6LFoDNM7W4FRlJNU8VjT2otPSIgcvF0hx5l6YEy+hrC7Tvrp962qj09Mh
LbWOVrDeEx780gOZELJVXc2nRHYJbV69JTgEoZZDUAAIK6b8hfWYswQaOcyRQeBA
Ziou6vE7X/LnmwLd4VoTGAmYPwGbJTD+kEiMXx9N7PiD2Tq5WnIdxBtsYlo5gkJU
fYuaPK+dpB6+cau9hR5EnH4t3v6b9SRkqxsMu26WHKAsMajyRbCT92IxrPbZGZF7
h5NpW4c9VnoFx9Wt6DRHL9RtTX/59IwcD65bog6U4xRFll2VVUCqnogK8fhxFjdB
LGblS02+Psm54HjvWzrSOT6tvRTZj0VqnsHcHAcOAI02Vtk48B0bAmH29n79mDKf
Kx3L3DRbasVf8VJ3SJSuMjp486UbdZ22YbBxgjfSkR7K4OFAmr6Z/rfeUCYRk8mI
5pcKiyvTX8yCD6ttuLDbCCYk+FeNhuyiX3YhOW0lhaZqf4sUTfVJbly6/azkEDla
GJwZEAv50gnPROZCsHKVeNdsc1J4Mfz+cXii+p7Q9gUYOy9o3uIHgNphaEyEBYWj
9fgM4DthhCDcnWLMGQoqfOlvfYewlWbbAlHnONwxCREpfnxxglRlFuA6k3rivPIp
LsV1v+aoKKRS9o0F2pNJZMpi6kEZUtUIevD189wieFtGjIc3IzpZkG1Vu030/1Lm
l6wMgFZXlRM7Oo193qxBSknoRNIkGyintQ1pXisw8dnzmSx2NmupwJzBKG0BF0IK
kK62SC+C6vlV08kOZoxh/rVPbTV5dCyqSyK9iKNRoizjFcgu7qZ0VaSYyoBgR5DL
i4tFc5rPa/ba5Hb34y87tWBQI0GYKxhoYdPLoCXuyulxIX99DqbcMT+OZ3wvjo60
oCv4R8xkZvOjplbBiJSRFmqwsZUcG2hcE3T1ch2Skq8UhMi1rnI8eIB4n/AYdd1D
vLcF2kXMU38laIwDQbnG3cEZ733GCae3HCs6WI98S1YPDKWt5A3eho3bjeBvKHEG
MnUq8ncFp53jOmilzNrJ+6b+Wp03BHN/uSM7vnElBORHFquVC6NihVZtpppm9oo/
EiAnlL1VMXPOHqYApdWPlbgzmblo0FBjUH5A9lZjXHFA9iSurWi2rSKj5QnjQks6
FC6TYaG19qG9qhEJ5nbF246dd4GQYEhL7JhGr4IM08aWKYg0KL3ywq44Hj0vbYYq
VZAaRbB/oBDygSdFWlx4UK+1O5xg5/6Qsy10J4HiQQyA2wwtJ/SR9O+v3o4YinDy
E0QTw0LmiM8gxcv2Iv9Z9/+8I6YH4yKdw8ANVKKkSVMsDL+yqwvFUrK7pKZF01ov
hflHT9Sod7xsiBYBm6XKlUl5MzIXYSIbqMCHoixe8Z0+l4BMTfnOEhpLKTqrfZEL
DNkBCcKTkCS/g1SkadZSDaV6KL+7SQo7f/8kGNaAGN7lez2PI+yYct3VSvh+MwND
PC1Xid82hZdxjErt0SpwtEmyyEqHcBq6xJNYsJ+3lBO5T0xuCAoWebpANlfMnD4D
WDbKZDCfSxq0J+qj/HY1AMFfualuUq7ZU7scy1zOmjCyrA4UHADRWX9zBv9o3cWI
qW4a8t63FA9y+O5tRDyBeAG895fLSTLUUBGaaXjvjA2hIIv9xOTiA4+u0PC/9ies
c+nq6E/KP+xx0S2VXaOGbd13CIFvy1j5B2SMTouvI1Hy2PBU+H8aBPBEbU5Ztx+V
klgbLSEwqSjn3yJPXWtCvnZuTP1YO1KgOmwe+AGKgrQ8IM1azOpWYKnZKPI1CkUk
9wq1s38XFxNSgpR6DSTBmmd6y2qO/ofw58y+B//HTQS/LPuVvMyVsX9kkLiBVZwl
XRGHl46I6aqgtpN+O91Ad/xmsrtHGhPRdTOIXQWsm5uPdMf7/QqId8iygNi7FKhX
rsAEz8uYFPR9DikgWCjRQTTBmSE2pV4QckJMsTEi3XxsQsypz5RPBhPMww3Je12t
YNf/q4l59FAodZfvTXEsSL+z4ApMLs4T/bdvUGm8pbrEuXijcbFoRKApmLTcTQT3
UF6EhIHN2HhDSm8P57cH0AUS25Jj+lU7oHOon1JEsKVZNgTKW0EgDoR8ruXAZCAG
ONG6McEJg7X35KJYvrz+ZGXr7NC1q8Fl+nPFjHIYTwgDUNlHk/6FszCy5wjyKUm5
xXAbfUsZn0VteUIgP8owmtAddP6ibge9EHgmRriCouYZo/2GDCg35XN/NVTtmDvB
8/PFGzrACK6dixOHJ62+QIRBIxflSB/euVw+g4XZFlb7dVnV+DMITYbY5YrMDS7g
CM7jnP56k/9vQXhRCPl1QDaW/zUWGkgEPOFPXosdsZdol09Ev6LoUQGS5SmdHpBp
gcFAjgYpgdD9UrfARn71A1QD9Bo00OYLs44lH3l/2rpB94ZQ2jgKc3zTBTfT1GyT
CpOI6Z2hkCOD9G7ecyyycOl9Vf3xaTrcsVDMwKuiqRBrVa00fu89Jl2vpW9qPWmo
ebrOTaw6Wm5l/6nVbPBTIRYYDNAxxgytl8UAHJRYqlQ3bY7wub/7IfY5R+qIevdF
COStGYtdsmfmXJYxSmnPTNRSmb8iCxN9LqbiYVbw4YTZ9o+pC/g9LUSAbX9Uq1g0
+nIGlz32GGAonbN1dhk+RUQ4cVtoXam9EuskMwzqdxNtrlNc+M4SeoQNqILCJmt3
mE1VuyJWk187K+S7gN0M+iAWIWPWB1dWZOjzi5s869wOeag8ueRaShjzveHG19zj
pwiXHSE/wK4HlKtVBvGVYbmnjSXfWdWLKSUtmQA+hi887kgSCS56MKkRL1RbP1eI
kNf0KZJtp4YC53Oph9ETBOW3VHVJr7RffKnxKo5rxybA66xE8x5UamoQeGhRgm5i
bjx6FCNJhG+dOWubwxXfaiJmhxAw4f0lyFu+gsD+wYzr5gDxqK/7J+kPXq0KNXKC
I2xnDHbD0fn4KyEZxSumrfle+9pQffD6v+gLoqdgEDrvMdbiAe89R1eFk8xQlfr7
Vjoc8pKdIWwyw3pUHCF/yTBZhSnPiJR788WjTb+xXSQ7LLcXMCC8Bj1SUhgYz1fF
cY/uKmgJp9BU5iIU3CftPxM91atWSO8t04QWTM3A1vGvARu0y62+LFV1PazIlbXi
+Wlrdlsq+wYDy3v8ph/xTqSY7e1iP6gnDIEh6sKsbs9V3RlJ/dDv/zX/kxNRnO0p
6BBvrWkUvcfTRY/vpotegwAaPNClGeM/Yn6tJBIRZhCvmZWUUPonn+lZSRGuPFfE
sqvplIK/I8AN68kWq9f/HaXl+pQswsvDfcnMmFpZFlWz6pH6XE0V/6DeqmpofLBN
vyXyUWbJvO+WUkTwADIjoBUT2s9Avi4JToxl3B//dE6cC11FoZJJt2OE2Atqb/fT
tccKfFp3A7MC6ylb1W1wZVOlJp0M8rvHR4/TW2KlW4eK1UuBbGewywysEPY/L+DB
4Km2UnDcQxfcLEC4RAN/ni+FD/mVbVmea/s03tYA/MPPzUV1elI5ty3k5oIDOayn
TTuy1PMgXMUM7Ya6+UjSrDX2IXmanwGHjlK2+U1/pRguqD/OgZfzO6pNsyJ5QxIS
ipo2vrz0BOSXWJ//AJvYyR2FKveUZQJkTEUk7TZ243DaQfrrOpwfO/PBXjsmXrwI
Lz/Hk10gDysDtNeFWupoOPDy8cU05mUVZvpeX86KdXwKcBT3pHTmvxhBwn1O17LO
NB8xvpxTzpirvLUM6Uf9KMw1Hs44yoFK1t0q0DQLJe+nG8O+8o3qSeSm5hzvT/qM
2yA2YEXFd/h2dP91vu01VHIZsrA/+7aMo1JrS/vv0E3SE1pnY3eTTCvw+xPBKt1p
QRQ5uR9rpHqaQrLELQ31GmdzSqK9VklKDia8hM6F4pKR4lYmWDQtNPOtz/7Vhhsh
T0nuHIwZvu6EVHdbHxolx70dUkQSHOr6h/AL14cgQi8g4q1nAqwYpRHAoI99+Ywe
tybFg0FpUfZFGk7GU2XrnvMrr1/LP9GpNdbg2t+oNKII4Fk1+1aAS9DOfQhCcBDA
RVikjhUUj+zYCIlGBEtCFCu/iWa0O+oiTUes6sEKcaMqHCHXNZbfX2AfkKc7GqP3
w9ZqBKwrlg5HYNi6BIlteBFL5UIixMrgxdl6gxvKCRw3FPvQAk7tpA2u9guR5NFy
5dR5ozgBSEpN7Y/wkNUL1DElafJtvc3m7SpjWMc4FzuUqPXxlRSO/5CbiTKutQ3n
pEA7qHoBQDYeuereLwvKdIk0jdZWj4hQstU6FtkKA4cvrH1wTj6WGQnBZRjPkcBy
HeAo5+rPjr7q/u2388IHbtqG+AO4OLZSYEPsII22AcI2z3bcPkKtsenLjGXHkSxD
GCmxExTUbkS/uz3eYUlEoFRvIePr9NYnkwm/7TWtV+IY1VZZ10QwsWQEjZW99sQd
OBNaxRXtF3Ecy1QG7Pp3q3sfw6Re7x4ucV2EPTuJHueMkhiNaVcqQFbPre4O9Mqh
e9vg8Ssto22Bxw8f/M/2IKJuQNGN0mVmpKETnMBLcn1HoE0qYivlhrRH7TmpnHAr
OtEnpYAZNFZl6oLkGoLagTMBe6Zr7vnZjfqL6mIUK93MF7/SJomCBOru6ivwy5dE
cNvRoRJz7BQEQQM88+F3CGkw+8yl8qc25wzOjeClF24+gvXmJHSENOtApL8Nt8MM
slm5e/rm5TfJFLBXTCWbOidRem5PJDkYmO2i3unEhOzdRbF7RPyt8YiCyn0ry4qf
WDQkLgkaivl5HouHYkLlytpC7U44xPpc0RGuazEbFT04atg4k5xEP45M9nT64wDr
kF1b0D0FpMxH5jvMryG0EGoeQlUH2tAHDiwQqLPblSdONow+Xbr3PlQvYg75Hb4T
Jsfglwi1G6uJIC7jDGt48ywB2/532xKfCujwCQ4Qq+3kkmAAzlEtszn+zxu0dgZT
GykGqCWCm7cyeWex3bcXnTf8x0qHbUqbqDT/DJyVpp5Ap36clxo3zCH03XrbtLeH
G4vgGmZx+keP9gd54Xu8SxNbUMoY3Mn5GwN+pwu02uIPOAmMbpwUzaGcVCLZeZwD
cw7UVHwJaM8mS1MvZmPKhbJ4WIKVsGp8m4j5E2CxPhnH+pvRopbKj5xzdIa1znJ9
iexSqoxMJ3bLuSM4dNgpZDz9SVDH/B8Lbh5ww/6zPlXpWzRHa/cfOYJDasEhQxEn
cLHadycGlJ86OXo8e6jsmFjS5MtG0w+uvLd5wp08+ylUzmm3GgJG6LPHrx6J2avP
s3jJC4UMVEBv9QAb1No8TVoJGX+MN7uIuN6mZGzeU4AgnpA7fiWyXppplvjnPB5r
B3icFZvQy4cUPFS8vr2Q3RW7XlV7iwZBX2H/MPpfdb8SibueDhab+NhuEKOyMryA
rC9kd4xnB1TPkHB8fPPD9AcHOoOXJNYb8xSaP58Az8EvTGLpN+QV990gAwFDGuTa
RfLxi+vCngoK3QFV7UKoda47cqi/wTzVp3IvZRIH/l7uErHtDLzJu5botvlbEOwQ
kKG2t9E+C7bkiWr9IDsGX7TECdl9s+Wl3K393vruwCiINryEWTpcpXaQJr5JC/O0
5VMTj0Rigm6ixiGPT8CrlsQQg9vjiBmFV6mg/WN0IndbvXdURMK6vK4OqxME/y3W
y99N2LJjfctQxU0Z68qgMIuKBCcSAkeIT38hZh20LGkWrAvt+HYPPsrYq0EKL+Un
CrW53+96K/T8IF15b727P4ILovSldCc3q45Vq5tXq9szuDk54l0sMnQDp6oi8Kcv
MZnm4NooyPbDRF4zm47SV3sTYCeu4kxF8pP0VNTEIIM5K0UzGFGtHe3t61Fbm6Ub
bpqBBljU9uvz6jLCqjryJ+JHi+zrfil+4V3/5woG6ho7/77p3J/8arJgIgJK9JHy
MEy1oGwiiH3NQUWbqTkJqN2SuiDgWjDUvXjgWUvSBaf/0Sl8WWaUU9S1plfzVejn
3x7LHCHVykE64uYII9CXuXkcpkvKJ+/DWf0iAyZtvQPJoe8Wd6yVQ++WyBlUOJiN
QVCHot/VnKmxVcekjRCPmnDcY8+V5KpzBF0pXsUIl3ZQS49wrjbPfMYahkWzpJl8
zRtEinkFImRvalTNkeXa9wT7BbnVYitSaq2nfbTLPBBGljHbBwmzyh1qCIgrwL3B
8P+O70bz1lNvyWw9qo2bHWN0VA0IbguoHbN6mK8OInvY3ja5duc+q8trYqKXS5ig
SNxbScvxY2D1+SxmltjW3T5/qMv2JPNKLfdtJgY52In3XfCGMoRAWwa8n4geRTtH
WeZ8yCq0Wz+58zXTEJJX5RGkqnOKx4e1Zm90RRwGgrge1THBgfvQnusRe13DD52/
BvB6sGIzlYuk4aEM6eGK1owlO8C0icXeG7HugykWbJypDyLvmYvs+RpPhxc5nCTj
rI51czce72QfitAO7rTx4smVkXh3jG9xRnjdULQMbQpNXlNvNwQszCzEi+zpY+A4
9tnCucDSdzoN2rFyGYi59NAfTAiGKWT1x6Rihn/aGv/RdnnjHg6oEEsXhscM7FtI
K9M2tqgP+OX8VT3zFMs1cgTTKGmLv9wdi1dNFChvoecE6MNVOrAC/clpzSNodoiY
Kk0SynfqAmsJsaRiJ4zPlnE7zSWndTlNmgz0pW9Ghi6xcMBQ/Pysmfmqhj0h0dla
7qSzkYHpE9IfaYJeLXgVzXCraFK3Je3Bgcu9Pvs6jnbTQ+xDrQrNWFG7Li4rAhLL
xaf0f06S5Pumh2wtKuupenrY/Kpn9Qqo+Z5nZwh23NT8DW5sJgdgay3J68abpKpv
W/I9c79IZLrE/85Xks7mTBfkTEEW3Ik6T1yRbfr0O+zmzb20ezjg+nCF3T9LzERf
SpN7mTTZO4X3ShIqWX5xVCWDAW/sAWHFD3cqi3eppKgS/Xw9IIpy5HefFBPmJ6Ro
lsP4fxM6hGSBW1iTdGjjQCrKXV6FfSbEIB4ft74iPHIuqVNHmnNz4NqV0i4kyeaC
knuUCkXFqYFeJun17IpXv88bGuwP6sj85psbz+OH8lNO/hlBcU9ELmE124dRcn9m
QNBzuypfmd3g0h6xetU81/Hh8HgfWBWGR3XRsuH3LoJ8yUYwbxJYO9MemLF0NZ8z
jhUjMbP1lQqGMCDkhVvgzGbL9AfxbQXQSXSbxyfSfseh0j4qu51cWQ2lxeRyN3sJ
2mePIjYK3Dh7ynogJ+uICl5coPWN5WUD0RG725/hATasBNYTEWmIugUv9SbfNlB2
ms2S8UzCSCQHc8fozVHhv0THRHwyOhnOk1x24Otr3sHuo3F1K/xVTKPlLURHoPwj
eJ0dL6TxVY39WZGhMopvYqSNp7C663FSqf9O1uHbF31lYisoBomksTLp0F5TQ77U
DKlAvjf4WYO+4DY1bvQurIMYLOHPLet5FpRJaPHP23jfHIpyo8UlByX/1yTdDVQA
pKnZxM1Mh860MLTYN8PgsXFJyCUuoi514bGqMPDXn5c1l0ZOA+xBmAgh+rKqxV/H
dQs8jnXmYqn4/5vmucwlGLjaad2uPq3fHQs51N6uUtaCrBwOcmuZ0oznhr5pFT6d
VKptVQDevS1n+768FyjQGRQqzEKj5QV9X7AP+OkU7KgYZSGlTCPBU2v1MMSatDG7
IZZCXkRJarjv4Y6JVix7ZdgYuqEeLYBMn2LImzZfaY2gMTbXyBmOry3Q5FiaUVx8
R8cF9u7GrYA2zEpIMgwqYo0CE6Hqbb8XoguVoZjHGjBkJLvp1g5/Qs0vELXKgeS4
OcZGXpR1MV40hJuZMZYdDa+oLttrkj9hQuFcxpnEMTIQGZLOGT9kKxUfagxTpHoD
Ow6BR/KLnd3QNJthZXic4KS7FNLe9mhNfiYdmcJ2Eu+a72pO32otcw3mrxdT06Tw
AEY84YO4PSzt01LUrC6tGI9KG+KptFNGWE/JfU2rsgHc8mwlHRLmsFsD2DYqg1hE
nVTcx9lco0p1WnF+vMsP1jYvrnBOO6KKbwpKSh5CyY8C2aqdpX8bRQ69oyc50wiZ
ogH56lBgXpvlll13FB9bj1UtzLn6/TnuUNI90aQPJtstVMIqt0YedzJgSTEgztzC
X6m9uMRthZuFqLzsPZN7g93PRp/OtXkguvid7VzFwKLdS3NNMAfl7BCP9zXYEXRi
H13gbhBBxUsSsxnlj8RYjKdOVpJxm9NaF+56golzcf+s0MV+RL6dpylsZWTFLlaX
fkNm77ofG4eZ2phSfKAWiqM3jr8HkJ9rYeZbyrfb+gFDR5T3BIUJyCPIx5ghgR0y
2NNhA/KB1B8xw6Chz3OpcvSU5fIIDgKqJk1kQ0AtKHT1mPLP4w6it0YdGrMvkELu
NMBqzbE0Fjk7EdR+1RS2y9xpcn8bAYQTo7ckxn8yllmFcNFh0BzwfPTIdfba6BrL
nHUJQL5Wml6XUwyAktF+v9Z0ZbX74RVlLGDP2YuiJMfx7Qo55hGBtYleOkqxsJ1a
pA6YkhYQpbdn6D0JbXShE7if2yrEtswnCump407Dzsh231Fr8DZHSmnyvuchiMDJ
1XVv0/aWqrIWwlHg4+pmqFYOqZlV7i97hPXwJSVYWMsnFzA+b6uWJJUvd0zt0qDt
N7RRdpCyo96AHFe4U1vMV6AF58eVvpZOlrWCBgo86LtmDoX5SSLByZXd5aaX4dMc
8jhA5T234SpJK2f/hUM857d+lCm86QCGgmogMzh6FJOYVQ+MhWHDCFO3k7Jpl3Dh
mlo50PXM18poX0ubC45QrEIxb0MgXhAssh2hLF92j0GpVmDM4qAB8G4jQ03D5znk
DLg5EDOJ23Npvj3hu2xEcyxyLD4Kh7kckKiPbKZb0oXKvmcVUwr0ICTPVLyRJ9sM
l5IyWfyNr+yGUfukTXk660ZFG0jpb1jqB7LJv4PBZpiQuxWDDe3cm4ciKlVfiBfm
jFvVgycBZ8SA85WcWyhHgaLE5/jwSYuE3lmMqH1bO0pwt0bsfZFszN2NmRnTr5ai
KQ2qpCKdbeHz8PK++hXv1o+DOO1UVVrwahkH4Rdldv7BqZazOwN23lGWrSjVoKH8
rXFRXEO5RDGdXUtu8BeFf+usc2JCinj5aIhJygcsQ3j9AsLPgV5T0qvqyqakePow
wjwNeAQ3IZ97sw1kLKTNOjGfF5VzSWCulkH31FtpzkQqEN6+gnM0V8I/uz887MMm
fq2S7cgCFxvsp5Fzx45ICE4rbNfFrGAjiX5qO6qMhfPV9ByDWOCh2iCr9f+ihmvy
TTqcl/yAhtLZHOmy29hCoNU91hqatQSLMZaPqQxm2qYDh9v0+HxUljnl7tJEAnVG
NpetHaw4KVqzzzc6tOY364n8BXT1+8kYis0YwpT9knUBhydmWFqNXb+KyUPW6na1
6Npwa8lNY4kSdJ8m3reR4M9/Ld+VdhZGsK7bAXjloF0NtCecndiew/Z6AeetuMVf
6zCupEpZ9+gmrY37EKuo1R2+FKDSBVVyvxLrrib3RfjRt2vlXo/dKgRBx9UvZFWA
dfyXvPzAJ8IKVyc8OJ0BxlCnjgH7dvkTGEbbdi13fg4F6btH1tc8nAX2n5CBGHyX
EdFbHC00xcXgQIjzkJyqVRYjLIcXwwdDOz+oR/4wNJO1yRknelLgCoNV3QnAMOJe
IdFZGqqIZpOVxtBuzA67zcgfFMOApEYMbArsPZYffZJ6ZwJRUXwTFtoQYQSDmFVl
qnlblXswzUAq7DZmVeeDJ2oNdsjv1OXw0munXtVnW9IRt7cR2TQT7GY8Mtfwoxd8
Nm2LnxHgAc7BhjnOJy71u4KpkQgSrn65+Vdq8/Ot5kXWSNAPzwsIbQa8YVYUhtDT
FhkSfRg//k+Ig+TJgiK5giBPIv+wfpYiMc0zK5/FtQako0i0cshbbNUWaslzNQ4S
fYtQvgLlJxsihNdGy6h750kWZ/TnQUVyptO9EbvNRSAVfzRyYglljHQhfFMMR3VR
se/EEOEW7ALcS24aVahFKgBWRxY0Jo4Cr6lhsIvIffPeShJ468GY6Vr5OzP6qPtT
GMG9g7PiSEbvDaPm0MRRG/orpIypQARDNbbTpOVjhsceAW0/lvqqIKQNLQuyt+PM
ukv0XHe3vUC58JiWR2BcCEzadAck2P7oy+AE3izh/Gh9oeJSt9NxzdH7ugsu7LUc
M97iIBtZ0nIZCtpV4tLEJpIW07nQa0d3n7Zwcnqr+Sf5ISGL0VdLGqeSHw1NyhpR
MNNqCaAMUeoNdLsSOjuIZmUcvsP4vP+xWUEq8dsPNn5w66o0vR4m+FGMZ+JRxi/8
/EHd/2C8wOLC51o2Cj//TsLpQQE/38pEWZRg9eAbhQvb10ln1Z7lyZSndcRoNZF2
74qsgD2n2G6C/j7KL6XFEfxYYw4jz3BKTtX4UKIUBEPzBdJIqybfDEh+4wuQdlHB
WIyL2HfPGatQVN4zA8SO7R/xcc85Bq4AY2iDPjyE3+LkkYj2fA8HeGbvsw3DBLWb
EgfIR7mETR7O/N4/s7t2lmYF8rm4gzdC2mLgjiUvw3DkECGNHU9H/6WnLqkdZ3mC
MJepbKiyWdd+NLmp5gqrVBKuHh4iYWOrxd9E5iUUhXFEBIQwCA2KrCxSsUd8Fpne
ZTB5cHbpSnNYDGSz0zech2jAB/XSr1HSMGcraRUcXK2Gq+hjq0JZxijUKEZdhhWN
lhRo99GfBVVb9jwo2u35U6aAAwZURkGKYflY8PveS5EtfSnQyOKZJfAd8xiajANC
BeJvN6qwqaBqVhKw2wGQlEK6hpfziIWKdEtMazSQkd1ytolaiDkkvWxwgIC5Ytj7
KrT8sOTrfRR6nzaUswIU81fFnVkeoM8H0+5v/txg/zqfoH/WXXAto9ib3o2SpuhD
CH9TVzp7CTuuBHyGk8Uof0jcn93mvGh0IZWg4J0VwYkd60cfH6GXFcNa40RfMn4u
bNy7vh3sDKIvODrozy/kFlxNW3mw5YHbgXMm0DDpWUrBWi1LXiWMwGeZDszsZlac
PB3CXmmfMZ6yDIXEbqnFQvjLCMgUfbQHgRsbk2ngVOieWZxZWlgYEdyaTVSMAQlC
2xzV54voXRBY7o8DxDc82sZm3QglsboiGnOxyCQYH2XXd/t+bl50O9rMWB0Jw7OF
pY+iiiBAIRYOn9Vr+OdDTutpqDL/uBDjk6u5pM+EV/VOax/4eKzKg+szoqu9Y6gN
EZNMSQlNAO6/j/lLEv2m7K7TN43K2ZiGHUXmXgN0YjYNS9M5vJV3pIm3lBOyuS9U
Nwi5hzCbuzXcD6lmNPQWxbRvewGxukLKH+1/cHqaIOn3zrM9jRU6iMMKBJlC1Xwh
rpur9L1o7/prQufob+ZexNn3PmkqXw0+vaTyfsDPDawqBafG8UMrX6qCfgKXSySB
9/orhcAx/FdF1j8drtq3vnWqCEr/EAaNFt7xd8fecMGRbGXcy0q9+6evSEf00kIH
oHJTJXnA3j6W0fTymaS01NNYt80q7cRyBjYQoPjzWCzdJn+g9GTOPzt+Gs4F9KV3
FOu3VB9lzEpAVwRa3G4IjWy2uMgh9NhJ0jq2OARXtD8Vt8zEzVKRRpKd6abz9F9V
9iDCmO6MAyL/J79nIOdlT+agsFyE+2wrorbzmR+/nf6fYFiD9aP9hHHG3zfM0beg
lm1BSvuHpdpLjMuLvbKuQ7JmohmsaGcmFVW5zMF7mJ8IKLKVnK2aErCmQxavpY3/
pbdGOBqPrZ3pS/y8PkMgh19Z461m1VwDQ2smvQoUan7BSbxeZdilaEyBlQgGsQE1
ghwhZgsXMVwHVy2Li3tblZkRxedH4H6biqdE0+E7utZDg7MPpsuMS5LQBzCipp4u
u1nqxvKsEs6wHdtLOC0ZzY7swZlid3YLh0yXGV02hp6SU02V/1IuMjDdjuLBiIvp
mtJJmjlKLmvG11uehxx/ezCp5rtNA1jXFCSeyYO2TbTZD1PUJ4s4+uxM1O8xxJgq
41Nyaprc4NdFO3UUZsYcOE+n6TTOfWv3rS7G5ECZGavVK9+TUHkdKkYin0hhb693
RmMw42jnV4IOFC213H8J0hkvBgllLBYxdYShtF7Cd1EtCgtyU4n8YZHAmK0tT3UF
O/h1hmJCTTWScNNq/XV6h3V0cXk6Gsm9mYMzcy5B60R6NttdstLwGbK0klAzCLzK
FpGMu2pKH7beU40hxvnMVpZMG0lc/vS6dolxkGV2T1x+MhY/Gv+lF8Wroo9NDh7I
blOFjk4iKHlzzKCDt/RCQSaHIeWXNiS94LFlMwXh9pe7MzrqMHHxghkaWstT7Gt4
CAZZkez8B6vDYPud6EHCXV+h8DpXpusW0iEu7WsJa1wEovp4/IaSWSCvY/VQXinb
vN6Ok/jI/TxNT69am1X9vlamC2CvZGxpxrdXFzbZNDoRsZJbnZ8IOZjZwgWPHUeA
rg3WTKcqxX0bmOLCIG2Jyadk75RUslKnubXmenZeUfUx1yDOgwBLK8+G+Uru4WrB
MufruE+dx6W+ZmFGuxGaWLtqtWSKWIobYx1eFgJdenNz6okRZzUG2/LLzuYemDLA
j8qKFQ+rtT3qFayxckWuMaeEsxpNshZkr2cr7Tmfqkksl/DSJktgc/jXETCEgNqR
YbWil92JBcH+gc2fGeANUK1xxUaBsC79Qap1rG9wCyJl3BSD7BfR7+EUHCVqutfS
U+q1qVGffZEYaV4EVjcewAG4OyCegTLgwCOTWzkQq43gQe02IQQ0eWQbbQ8BeXBi
3CC9AYHL9gztWmvD93ONBVucH16X7t2AUvsGuSWqihFytcSkjhBdGHZc+RdPHOuG
vRCM7ndpwr88ek5h0OWkU1o2IdtsCSy3ZwXYJxSgtY9K6CaIQdAZ2A1BVJ2lZYPL
6Y/BniwGuI+m+fEfbPIZLFjQwfw13MgSpQi8WPvehdC/06tX535CI1jm8M7im+YI
DPkf6SE5aEdslHxG13wcPQWTjJ6IvrBF5xWQ8G/u8jgiwsAMZHmKUI9dB2a/Lqs2
Km/1RScXC29s2nk3Bd0ZJG4PJ+4la0HHc6AdYs5CxZxNyxnEgPgUFaW4oNllUYVS
EviqfT7WFkIbzM9LXz61Fa7qNCWypQVyOblnQcHuJJiAqKNt0jFRsUyS1+ITsilr
iMmEbPaFJ+/LvKJUPBnbgPiGHr6ZkYCPKPuP4qgMjYA0ojZ09646jR5oiUsj24eS
vOZ4h8zGTLn6tFhC9YFOinbYCWfMv4097E8PTdPrPGOV6oo26fUFBMCaQWkPFhVQ
6DgmKIXZD2/69gAyFDOvfrgXkT3S9VeIz8A1YwwC2jU3RACWr5B/W0iQFIhF7Zzh
XMCYRwufipo1jyY3d8kZM7I9oas2Yja3TCWBCM46Fc2CBM9KciOb68cohh5tQsW1
2KheJli/zrtlwrchibYIarYmJH9dqQPNvbsFRPdeaHS2BnnV616eUS+p1DpFE00Y
zE7bdk4kCFPRbLNdkwiLW/u5+Gx1LF7B8vkgQ7ifOPNYULngx9PugMHSqLiEE1iH
M3phdUvD8/ograBmKec/++lB9xG9TmAn/h9/GN8d5sImrjDfdT6ZlbkNlJeZvNJk
sM5+ox826sCT5x+EhrLU3hPaN6BIWQtTkEtniAskRTpGsH1vQyEXStdi7JIZ6NEC
hRhckvfTOuGgu9XHd4pM/fEIpp8ur2AfF6u4VEbxuk77ErU4FNbg5qpvxYbTqNXt
dO/j7vcAJDv0SujE8j+38fK2fDqtNL+vC4tfCbLjJzUEHSWQ4QdEnorU+qy+19Xn
2Qd/Gv06sWkbrGTj3JwwN8J4rHGvKUVGk6jpMfWyB0USmkf3SSoGggOVYS1wyHz8
0o93elmLZjb5RuqFd2/nWtf+Jvxg5Z+X4+vp4jwQg5YjR4JbTcl5M02sIOYuOa0N
boI57dOrXlLkxlv5YMkEZjyvfyiPV2L6RiIbV2BM+nCGSyna61Tt6Pk3i+3P5uND
qXBVaedCGj0xOc4L2KEaot+NtSYMsjMraFFKLNj1Q6FZ4YMJglMnQ0oVHInv4dJu
GNgVrGaeJIQwM0toORcEWxstO4TbTRevyJz7v7dhXY0SYUok1/gNgGhv21rtxYr+
IuF9v/Eeof41JElsSM7s5cCCG+6F8WDQg6oz5QvCJlHZVN+GHY1SHVEDIPPNWNjD
y7uclKpcNZea+cMTP4PoisN3ejKa76Q2fh3lgHnVbmwygUX1nsJGs8hrQ7kM/V6L
PlHScNfZStyJz+QjfBH4Rn7S5etN3UlsOAsDHA/snixEIab0Ws9FEOyRwB9sJRNV
iteCEZhHkZ7AuXJz+rxpA11msBs8zrolMl0ofopWQQ9/30yPu5j/YKez8wQpHrj2
h9mHuJSH+wwAu4kE4EhpCtPG7QpPQZtoC7jNpheH1bWBH+o9FTRmG4mu44aSfa9S
RiGwMP/KEVKFZliU4P62NJxY4/QeyvHaOeY1CtsLZpyoZbpak8VBAsm7TXzn4fBs
7VCWywSWPnW5lsZSQaKFfeZ7KlYVvL5o0ap2sxtfBYJL7Wnhmomi9cCQkt4M9TM5
X3ydmrk7dWO7qXrsTbA0yPXEEnA7ayTPsFo8Z6yHYerybr0u10wqK/LMjwgEfwXy
8z+SPqSCLhfZPDg9oPZZswFSQgf5iacZhYYHGM3335XYCZlz06LiXz8L447XxocD
JdaCHc1S0ZFvUtp67GcJpQpA/oujI1SnwsXTsIjwVlSsxzbSKvdW3YmrxRWE5ngS
S4Ov4vmz1hcG5gyEnH+UMGh9fkkFQgGEavQTrxl/jW7SvdN6dzuWRoW8UOdh7z4n
y3gRfrKijqyyOg4deAXtL5qRUSL3cUgjIabAgFax9ijBv7+32vrpIs0ncWkm9N6t
4M/4Wcc91AMZG9fwb7/D35SCiP8dHlOY+V7rYf4+ABAkeJuAmHu93oaDJLvFgYod
hDOea7gO9uTJYVz8mSRMtPYe5+0HKXriMPTrUdhUieWX3kKXDSBwJQZkQ7J4jY7Z
7LN4VEfSBpO27QHVlw8CeXnEBqrGHWVAxaxcFeH3qF6ffRzdNe8+s3mV7VtuanZN
CWDyClNAammLZqvHwzikFmOnm4c1o24D4pr2N4wtDibdZOhDSM59J+mfDcpLOW3F
Sn32R2Xl/YiZzFeZLc5DP1r2uhd0uICgmYQSGI6ae8pz7BasrZC9L6HRasOSz+bl
IIDHem2jb8Cne8l65HS7z/JsBnuUOg3CXMcvX5Ii1S1A7Ju/dCBQqSh9Atxbbp5P
Cy3tqlaVDopzbFaOpxuo4SLnQClwmAeAib4l1RqTlIRKtTPyYxY1OYQSn76ZKlfk
O070dPHsPZzzBzTa8KzgdvIsVW4Ot0Y5rAJg2ni1Z8eiNOqP2pY8wyboIdDizvxC
LqvkeiscybUkEZ8QxLVDsPPoNFQCIWzTD9l+IbdVMBep+UQADk5H5iHeqSoUDJSr
QMKOvrnr9RtYq0d7NFSeNtfo37upPJ6z3aBDBZWGEEsy5Dkt+GZtmuZoUHD4X0XK
pd1xDJZXWTjnBahgB9d/vK+nBKA1WprGFgpTH6RXaqAz1fR4ESzxtBCrcQ8jJ0Wh
qWdqvfs8oTfXqcx4cUPji8pn7iamI+4NntGDCPDawYKr/OcqS4c2aQG/txHgKSHa
yKayGFJ78fPAWHGr5V5B+07akTs+A+deO5HTuVE0DAVh9hog+aQPErdBQC/AvVGv
9W1iKjXRncMnLLU9dmG6Go+gg3oHnc7Sj8Na4BvNoMFJ/36kngw9vlehjooq2Zrh
b8F6NZ4cVeMetsjLiRF5QhxNhpq2971ii2XC0DKAW5d8M9FCBznDQAgCdANzLFAa
vMyx02yPxEuekjJMAOS7nMPUKX7ITROj6pVu+78FSeMCbBLwRY2LHB+OH+TvKnzs
Vps0Pb+yQz9ShaLa5SHwrKUkoi1RBxt+AUr4DiecELK67vIpdPn7L3cmmYE8ioUQ
GWTVd+pYLMk50LQfH/85LzcJ9XPtHsbkUZmK+XfZwHJZ7FAVsBaPDXnAhLoXWtt/
RC+bDuH9LnTSkfUfdRINBK5iv9SfRAVPKhcqZyJiXViNegGwODpAGjbwRa/kV95a
QanRw8/nVqxZo1h0D4bKazkCLVVbN+fzdqvcTK8AKKWYCtrJcsuzoSUrAE9Z1kNP
qG2X/mL0yvbXR0ks7BlPAlu9BEv7JSN5+mqFxPhbG6UBUCfj/z0gswrjC8EhuM5F
wkGdQj73Phl+WXNnyedcsZPbcZ/SElfrGU5y4si1E76Jio91f9Etn4coSzX3eEBR
tKGW6SP//U+3wkmerl3CkAfcZpI1FACOIeppQXoe5W+yQs37DG2SUAJ/P7Kimki3
tXosXdA00WRo9M75O9O5a4WQNHuuNLMd0nt6SBxmc6k/gB8vwjwFB2POwx0LZXbP
jSOyZLHxmYcIbpo3gf2JWImf9Qw4i4OI0fvkiVBxrt6FIcNlIF39V5/BnEqUGwkg
K5Kbadm5TdK4S8ghv1NrDzHuB08z89mNu8ttSu45GHg2cf7iA7wt8uZULh7KxKCe
c9UdVIrtFdr1Hf82x0MwLtNHzO9MJRi/Z8NmMIDBzIV7ACCkNiHMV0rn7cRuLI8X
F2uEdGLE+wGvF7KqwvPB9JIABb+Xr1KEp8VXWoCb0IqRczAWuNTwP4z8c8y/8qZE
x0hN87FHvNdd9yT88h1dwxNC9Wjg3qu6DKRdLxqrBsJKtBqGgxgnilcii1gqhmCA
uEeyR0fs3CgpKPUlrXKvjN0K5aKxj9muBF2hfHfBTJuvRyElRavDtodHW5VndWFK
jFJ/RnkE+6cO6RaC1eHGQ4fu6IuwKFRBym7cHXynyFaFum5urxabUa3veGU2ZyL1
EPLhjveixH8EvZzNvLMTbzraUasdWMBuxV+YnHA28A4aKQqRhoXDd7HDa71V+NIS
SINe7j0aFkL6/fYe0OLZjXr+fRJjk9H6/0Ly8SLvAY+krpPNXfvRKqcMzBug0fNN
58NURpptdPuQyZZMb46g04wOGWwNtS54N2bR9aSR2q2SMHKRqfqXLyyF+pATx1Uv
nzM6HdIzE+g3jbcrQEWBY0QY1Euu/l+xyifk+vuc1xcwD2RUjWjzEt3hXqBn4IEi
XOKNhHHLj7t4j/tnPqWcqmGj3w248Xh6miIXB3KwL+j2UCKwPkHgr/LUVr6/ib/e
ZVHaDtz3jFLRrJ4TZr0YCzdvhmsNYc9/EbB+R2BMxbIjJ4SctGNhF679mx/DSffE
/xfhksp+FCWUfdeDiDiRpqkhj3/LdKGU5KrbBAjRyrKq2czwZt1vkIiRSUo8zyjj
xOMdZWYe/cI9zh0zZWmsjPnhdQR1WOfLwu8V4rdg+HBo+F98zQj5we/N8ME1tRG1
FModfF7xnga5JrFlwWB8jbsWN/kBe/F30mDsy86juoNGnB88ZaHblzxCefdFvqpa
GwBaQffvQuFv+Wjzp3wvwpi7+QOAAbbFjjTT0iIrpg/rvuZ0EDFf58050QEahYYN
H0KIaOOzxzBuSiuObGkrhc39Thcq3tvm3WuMsIjuQU3uvF4pi0xtzuEWBWRhvh4k
TJiL1JHMjdtu/IxKjIErJTl0ZRFsATErDiQbXOQhzTR6GcquM+qpBYu25sdgyuUQ
8sP148tB3huvRjHuejhzSjpeAn/EmDe4CyTgPqyB2gkiXhkwTITHonim6Bydlsos
1oUaqPjnC9s3eSFWAL23jG5vEIJgc/JlLvZZlS9r8IuFNvx/BaHOBIWIN58Fx6/v
Jepy+fD3Lli4/HOHaPlsvHQ19hZYpxtSZAPDI4kQvqvjQOMbu/s02oUiP95gkNj0
kAAP1FzrBL7uCz32zKahrTh4DQO6WJMZ52dT1AxCGqhxzpNWdagCH+1ZsbpJ9P9O
8DWxc4A0dZMC97bfKOYZeUyjjwdqMqfRudUeGf2+CftrBeLfEjd+p2uk18LXpQ7r
Ha8BfOovhCdZyHQDRWj056oLaN7ZXImCGytOZvWqM+E/qcGYIc+weDFkW9tU630j
3M8T1xHdPuVKNAmOXYAweqNw83gsSb9uw1ki7rd/UK1GEtjsrPSTUu5Gxa8jlQNH
qO9+5WY5iQYLmUocZ56O2GSeGMGva7vhFZy3dociiau123ekJP/OVZSdHKgOnSw+
MtofJ3fusvdQ3pAxYrKcsVvxer9EbI31UxFfWpKl+OFYc4hTBzJLPDJvXqEplVNq
XWdM7X0LEhaqTQfwbZvIfVd8GxoV07eZsLeB1DCOaFtdbnCtJLXMdbYlpaGoK7Eg
Qk4Y/qm7bFgh2NVo5gzD2yw1r4SO08jxpdATyNaRSMBw2BTl80HKIU2DFXys+vzr
BzmQbgDtMKU5sGx/EPNIVDvHelPwlydcxVWd0ozQClWxayOJP5F5teB2Q7c8ShWc
FyZpxFIjFfu8x/nzcpZ71ylhTGjG1ukEt98wDNYh1ZyB/ktJ72QmzJD+5RnfvrxQ
Dlq2GT8qdVTvTneAx2FDxnKb/4EMnuaVd7czcd4EZEDzvixAgtZfPHWoxkzITuHz
KOrt7i9yjlwfVWF+/AhLSjfYtkj7pp42dXExiKofkwB2mRpOFx+j54JGMs++tKTc
f8o3FoJ+j9i8lmJ2wa4iAaHVNad9IQ2HTN3cV4xtGJuz/eixKiAd9sQCOgW47mfk
yocjM2iTChcs034VqhhHxlKdmWcCh6oD8FeckVB6Srn4CkfDZ66D4LA2UaFKq+0W
jgpOOHdc8G+TLOdwGP+1/8ok1eZD27MnLbnkDQ0IgQXzzu1cCQhPT6aV0newQ1fF
SV5JGJsMkwdoMSsUENx+AlynBGz0sUFEusd+TZhuKlJrcQmAWDInix9qtE/iZ5ir
r9YIWR0q5JJZ0NoK8zlsM6Oxj8YBED70O40H2p4U3LnIq8AuhTZx2xXBXyG7gglE
tTuQNV7vwzj7NM7T+ikPp7inXBnek/jhTVD1MhWaZWVJtYO9Gn+d/i67KAb52ioi
nOBXuJkh/4HK3ccIG7qFgu/6+FMsfa2PTrSJ9HvnQHVnrJqLVK+EX0fq3HfNH8BZ
sQAv+hdYVNr6ACoMdsiHECupxVyEYBFWTmy0+vFXyLJmLVXRkSZq4ChEei5ahxGF
iC7GiaK299LVIK52y0NkyjadBlj3MVDWHDTzkpUc+fqq09Xvw8yNWx6+XAU+AJhW
En/eLTWOO4Gj+QQSlFH+wfhBjhWkAujfh/zVa3P2oIpk5jjAZd3mkDjdOw8zqGLm
P/CzX3Y209e1A7+jOS5tdvznzoMbArWZFekc1Hi0lsmfY5sr++eyEJZkSQUDSd1X
bMJM8Ho8oY0G+jX/UQJUHk67hz3dJS9YOyrN628r/qHUDMwklfaXT2IOEdot6D1j
jwK34sluGXUo4bO04jB3VS5j3GtNPSJBLWghicLfyM/Chjv9DGu9Ya507DNN0aQl
RBQe21qiRAskKqqCqKfy1z7BRNegfu2k1Nc/iBQhKlIQoXeqKo3z9yZjaWdu730Q
UofUkc6EetpU7DEt5jRs6pItSHhoHLVVdVCpcyO2MCgMuUEOqDRBYaGirWMKGSyc
wI/sZVSAdqx0Gg3nvkSBPFdFp6jbYV9MLJQrl6kQ+U/GYckxnUez6/X8oquZnJ5t
zK8YCX+qASX6wsqClvYsllaWVQUuINTteGREwHWprrRcxyhgMn28v6i4R6LYgc3a
CM3qdyGRqbfxPm1L+xCDjaztoDIiIESduo3HTISIv7LqYJzsEoqpbmomixVND1vg
ohJvLYkzb/svReDM+NTnPNlsD2Q1pCN9G5SS/ipsDARn+gN4Efp6XCBQh++BiuV5
hT1BrY0bP15qCsld1R7A6W75XJDyUjvIecPZR1qIUVe5DTa/wJ3HACz+Glehw13o
pQdaezyd7rOGz6oQJmh2JWRXHbVqBoexxdsaJqIlrez+Z2ZPNF/sdBysz0WJXhDI
Id38F4SXzIz+4r11a69/Uk4Bc50zaNAuYKE6UItRESAXECVLfvPJgGa89B6irivc
yTgT6XZFhTJvL7JVBMKmN7Hg1TY/0J3QsNDP76IMoSN3I7Xy7ULT4bU1acczgasK
/5E3ow1dZN7DbwuhPxjBJGmMRkINmPxsok9HfIhmsn6h2e86C/OMoH4v81Bm3nbU
QMMqKBq5VbcDVaB2NzhtDbEhqMJuW2v3FgjaEenTKtR0KIXBWRDeB8iEHmC+0c+T
0Sgp9Z1T685NOnSKzDsl8t6WhdNoZVVCsa7Uqkcfmj2BNYpGB25qFgG/b10Xds+9
EQAvg75+mfm/CDemXGkdvSZlJfj2T0y7t0usteO+sgiL1+IReoH3Wld7HQ91lGyB
OUox8M9wL0NTK7SfeBw6ZueCe9McrUtWPDfHxOFhO7HrQys5+0tIjeIWBI1wP70j
6KY0iaUoI3R1EWEIB2HIcIb7hzW7ZXm49jletDgoyFDvNr2OKQf0QAi3RKbl2uEV
nXBTMPYIDVfIz453uz8sGopfFWFvQMt89x0DsglpqWDjKakZnRSxKg4jNnsyHcnK
ftvmY0DhuAdvZaSLQ+vz/u8+fNALFQlWzDLIpZq9GugeHV5Jg+a62/Q3O5VpX8P5
JrQrvM+Km+Le0vrY+K9+b757sAUORjH+ykF8zunSt9GKHbdPKi+f9b3frBewYwqs
y99T/BatTABPFz5KMbAqNWGdMIKgOXfrn4Cn9SrI3EehrUQZpEb7SricBArX/I0O
tpszijsG3d6bkxrjebkGZl8tDop3dhOWLdIHd02f7oCQ5VOOTCP1PEEvFJkdX7K0
wyzIpLKoXSzX3btXIKFlGSK0f0Q4Iith7H+zvYUKPlB+lp+Y1stpHwr4hW0JeUVM
j/D2bP3zG8YeLpHbBS8efocAXjMD7r+wpoymhUcnASaNDW9g9NGlWMqaH/YaPUOi
zM7+vYw5nbpqZC8cZzMuPsB1nEiNzC1IjiDW+/Hubsk8zRZhhwB58HJks3s7xsEf
Y67HTZ0ZrOpxt+MvpeMTc6F8dMPpMRwu3xi/elbWO5J1IO1CeIbwoY2te9UohQay
Sx59WgNvQYq/ebAaPhT42BKFuS/2bw2tePN1PlljM+EuK8kOZbShyJC67L+RSl2Q
mD9GXy6TdI5SXTKg8bnwDaXD1Qoo+aaSCApOi7DNcW5HlgzasQzEhi1/ZL6Qjlil
H0UXk8CErizR6iUVEOlji1pFtdcXTpLEhCisJpN254ASuDaqlqzlcTGmkO86KOm8
zhpJc9jyYZcyohujGPIHvbhyupXlasYoDEU8TCG/2gkRpFEjPrtQd7TpV/9+fcJ+
SKikzw5kM/bsjBxpkMNeviblu2yAM9iWyGpNg4dEMl58NLBCX3PdW1LivsdiBTU3
sb2QqGQHtL/TyGHHJ4ymdRFcuBTSZwI9VHTddCWxHa09MqYnwiOlrefZ1u+wxjL6
1HlrmSgnndW6gA+nn8Jt+k+EqKPBkA+iVIUNiSGuhRbvcXuME4TMrP/DpBwhqrMn
3khXzsE6cUsAgZ7dEDrZbneKEa1PBejx8O9G8504yTQVi8YE+HthZORbfqhS7kTJ
qjlQP69TBIGSh+Z+rqk5a0VU59Y2mhF99aNMAe4H8aFbLIltpW6ryLFx/ayMPcYp
HsmWjEb57WP8DCp4mZLQ/LIufTsJ9YYJNG7S95CUflx2EbKUJBAHstkfnLpAYEGC
SdiV78Fek5stx3gu2dDoUe+U2s7CTJYS0vL2o38wLuh8i6+gjyHYQL3Elft5froX
L+/MHkJSEpGkDmfBKON8D/ihR/g54mvzVcYtv4v5/3goX5aNPvcfVFEkO+dOLcBr
i4qmnjkMuw587T2kVeaVJSkxtV340ESPL+f8xABdJ3bKwapoH3JNUJboh7iLaQ10
ZnkSU/ERDExZq5lUKdwh+kfetc2ichYFIfob5qulY7mWqG9zkFpEwkuvmZvsw0nz
2zATKuPguVoxxZ22+KrENERsLnfoDeC1GP/ol54CJpQ3rWerU2NsJj4VdhUKGmoX
l/onco+AaeQ+sWI1y1BNeqpEfzhfACJNfcamN+B5RvUJui/UrZQZ8O+zg3Xe7l1s
dJHsFFQncZxKx4XOWfm0pAjCO6PQAmF2UoQ90Sd4ph/eyuKDOrewoVs/8MSnQzmg
jb8vtMqGMIoVWOR122GkA2yhrqCX/2LlFCOolpv/e27Ul7LZY5KK6BmBrrG+tXkS
2kb0uuOKsTCQXaGjkrkUWr/C5UZQDt3lPhqVN3DXTLhr2XffC7YRRtUeJg84dW0b
J2P1Op85cCPtNVnjvJn8cwhyQDBC1h0UAYio/L86c6NQf6rIB7dGB+VX9nEphVRE
k5nHG+vNNgFJymFlV+l7kF4ns7Yw9zOVZBlZXwYgOQnAEod8GNiujR7h99+YEv7/
FRUBiJADAXNDbIVtq3oo2GtazBgv8w8ivzKQAjw5Km1S6w3h9QyvcbExXBwsHPkM
1RD2ZB1ffd7plsNRF7GrUrOYq6CRhrWmQ0ys/HjK9MCOE37Ys1rs7VEbHPsmGVQb
on/MtG9ljEDPUaFkyaWjlz8VpUScCVCAXiPyHZItgP5BfsJwBo4gLD4doXsckwuJ
TXh99ywX0Kzie+ujtMOorzFhQLpGJ7q+Stlh8MG2YEuGISbmwog+oi1JmnMJ4eU4
V02QjHjvT3sc0vVV+3rhtXWLKlPEJs5kBJQ/2/b6maeixLVGKA8n+tijSXyXhAPl
bZN41v7OvIKB+YI97skoxx7jfHDFOdL9o6j6+mw45fDTQ16u9511hcWWZX+OXHhf
sK3KE2RjkqHNo1c/kYmb/IWevQEDEiM4WHiXVhkjvL2ERLyOAqxooHFbIP9GwmX6
WJSq7KXTpfwIJdqJTY5qiWYNP7n0RNer9Q0ZbFtJcXXHv7XRkjisHlTjomH7WZDD
Ymd8Z+FDZIMR0qZukPLWzo4NJL0PH9tNK28DZUrFqyHXu8nCKFKVUf1I/OC2Xkac
T2V3n0GusrNwabHjPVkeqfjA9YCYiyZ+i9Z3qOhhBUiPLDK9voCdqrQYeUOEnfOA
QwxYVtE4AFvaS/IIUTws8/C8HLXPiK52qi81h5alDsj/gKreuHrlh7enkkaqXQpF
1Dc3VY+M+zc5dBkrTGMmy/61oDGcSCzkc6jHt2mTYE0RB6Cmplv/SxHl6e7ZwVu3
ERdRzvlsHTiXTDqWjrOeHe68xKalBDtn8WUhKLm1SKbYr0BrnENdxHuVun7XRzBS
T/43okH5JCUVeuAmQrAlVG/ajXb1BrrPo3qEoxsiMw9LPjahQN2E1+Fn1WKyB1GM
XWdb/DXtlX4p5tAewimYCcGULlUS4ZneML0ENyvTnPP39VD/Z15ZJzvrMNQUrGcL
5QD4md0JWSe+hOwIJgk0cIOpsA8qJ9qFWEL3f8lxN6HUc/jGWns/WMAJdpFJ7EfX
auXbJDEH7MHzrmVFDVPs+MUvItK4J99w5qrqUI72iAOzpemzrDQ9jdZ74yYbhVbX
vVLrt41Bdcqm0ScFHFC/+0i3Z9GNTj9WhPYSUZuFJngCux2LV+xgoK1o0wSoV+xh
kNe55fQRmVYo0wGPzscKO7AKjeiVq1/+arjFteOMuuWXbsBMtNDepvlAZkM3vOGT
7PW7EmO973ptlwoTqFvmspi/oPrvmzd00htYq5s5i1Dmse7o/fpcW6UzwHrtsGus
UL2pK6qtdH2+Fl7qvmhxAH2XF3/HfJ0djKcR8OMsxd4jN37/6cy1Ir/0JvWe9Qrc
tbq1O8lKSjOiVu7pJjXyLAZw7CujQ6cZ2vrUt35/w8NDiPJN6xJLzk0ZT+sD7rAt
8mNeNEh/uQpVAqMjPPXB2i63BTXYpE5Mfd4hIgZUTJDs+w8jULPd/F/QpPNbtzw/
EpQRAsW2pcqxbtTdDU+upvtIJfnjqlqX8nbwhyq7RJqKAUq2Sbwe0WaxmTx4b+n7
qYuJv5VXEGNwZZP1Ec2uYXk06Isd+eRjxlGsHV1uO2cFQEL3mHUmrjbcpHgnxxaq
gS5wvjPyJP69vQR34J0mITJBPRYoH+afuUsI0VPht6UtEqIxBgOFFwEj+Czs939k
+slecVB9KF0bfyMkVL3CLDckjIs1gAD5SUW8m2Tbqhzvbsi5xCLzweJMeXXPVOs/
AIl/m7HoXIoqq8iO+tze+uEHq+ONmbMg1MSxKmPGX7sw9mUNICmb9fH8yZqkcRY4
m85EWNQqdT3+gpbO6K5DjZiXGnly9vQMhDXz2kvDxY1i8Donqh5woJo7SIbpZb3R
fKWipb/3wMw84N3MTH9OB5d3d84u3T0+14obVjJeo1xP+OWdoLL3IOh/yfXwFzu1
3hZTK+OzzJ7c58k5PJLu38kJKIUtk1+4x8SUkm4f9wHq+zl73J6UBGgVQgv1ZyKV
U0Ar1uwEv/ZvAQxhkcJkR4xX/d1Ct9fY339PwM+LLsrMxkLeb6QEXUfjgQhrP9Wr
GxmV2kQTeHznstz3A821Ua0Ve/BgeFSh+0qSqlHmrmRC8P7WSeisEDLGg7pxqv4b
zGs4/YBkSv7x0Yt367gUeQ539TnIG47XIZBsfxUUkRrhZAnlj1jai+tt1ABCWRlU
nGiUJf32w3JzjBDL4TVDWGe+n2Y2wKeArxPky/tiehyL7h+IjIFilyunBTxNVSam
ZDPYMAL4wfR8jwxgkO/VlHK6cSioyU5r3BsXTNuV46R9Mcyey0aayCX4jEijttsW
FY+3AqEde6VJZL+2jRupdqf3E7h7gKZ71aVC8xQVxRqtswlyjrY+Hcuky/nyLg7+
mMxRXsc6WrVgSmaYncXkXv9TkamIUuseoI7AO5jshB8+RmmpjALV3KIaE3ol73gB
awq9/6ZQswtTwCKu925KnA81Gg/ZdiHk22b0pHZEH5+GtUcNWuDAFDn63oTKwAg3
bPVW65YAq8oOP4mxQ90ZvrlQaz7TpKSei5fDZ5BeJopgfxCwYnEjTXl/96SzxXHW
BmEYUoU66z6kq0wq9QcatGmEOo+vp0yz9l213Ws5nFVtZAfPlxks9/XdtiL8e8eu
2bbQ0hiRMH4BujP+mSD832jxdsoQkqK6FwgAbecEAuQbZ3DFTteDCvB84QJIMd3q
R5seMmuR07sY96yc0r5jjanczAKNRZR7mpwp4RwJV1ObXA/SUrIf/mAL2KhCGZre
j7VAuSPMmCJvMeYy7SI87zMDjfgS9uk/bDOY10g6o0tPBN5gY6qT4TeDrqKgtltz
NZdRaBNL/V1zS9z5s615+pn2I6AZRR4a9PUlz8bpOFRhhnfCrr9opV22XkeoLahg
1z2Urug8P0PWAbqKPDcwFe0RbYVmEv8UvBnEeINFkz6SA3ADJc70r53Y1QUA1uTh
svn9ZkmtW/HE3AFIQfymzcGGPgjpYqh6pPOQnryVQQNDYvPgRSRNB9NH/PxJnb51
+02UBdhjEr3i6Ow2aJMZEHuWbQ7WgXN8NpxUDsn/uzAJkPHCbB3VXc1Kkfia+Ipo
wwvt/GcMOK6Ciivi0JRYR+IPMajKkHPozF+tz9vLXLQkK7ysW4/ULpKyza/xkZz3
qhq58Xzh5mxa+CXQ0n5C5AfcRznDYMzrYvHRHmtLRLvRidI8TgXq0xVBO19PNCUa
OdYqwSBBsylN/2e5FU716hdUVKbbQcrQ6TDMV5wnmGyna+pksBLhEqSphr9FVP+k
772m75Notn+7rUBL9Wxz3Y7OpExTR4mZpI4BBrCgJbw2W9mVV7SR+1JvzEMk2Arg
jjcTRJ9b8m+a82Mpt52ooDTPysMDGhLJN6nnSlbGjuyagfmEewxKCX7cu0jNHM69
ppuB4VUeP5Dcw+c51sE+ZBNdLr2vEV3+IznOrvj9ynGbNWLE533SL6h2C9BCf+am
CZI5JC2oj1BjWwhJm4g2K2x8+PyanDdtKOhb8oE3gqhiW7CC852h2XpzDTJc1Xzf
yPkSo//s8wW/t0DjkJV8+S3CqI7d36/l6kYKZiUbPdRd7Npb4g6WEkHZGMuVCMIY
eZZ1lDo3G+WDIin2AC2iO7wlH/ikcTsHuQDYsCGm2Ca35obCaeyCxzFaS/Ii+fQp
v7t5NpSOTBll0a4zEaxpU7Mqhal1fLSoNJQbTNYW3z0t5nEINACta3P/ip82sDj9
e6dT4yy+vS9bg3cGxIvolzA4kxU4uafv6QTXpV17dAZpQ3sXCabT2gEwUsCNZVFy
qouMig4Tp+RhiRgeuAYEhkqxGNj+f/vFxkRWBeZghgvkiaHCcDlxRgA1yevsYf9R
pWxc8B6PHNIoU83F5p6cB/K6mxyx8V+ceRWuoMmiyCjozoCubNzCKsNOEc3uhZjS
DklpO7jWeqCmVwWWDtvWySafKWq1h6kwkNphgYLXN4rpzBwdeQG8XCcCCpQQwmxb
Xqzwx+jPk+q+BXnSBxqCi4d0hsrYWERO4W7ocXSeC+QCMZ3/z2Qs8UpdHBdnG2j5
VIzyz/hnt5q2ki7Qn0mS60aALYi9GCNiXLtV27bRDBrrH6RI07y0ZFQaczMpxe+L
hKvNbBv4zCKN9+1DKze1OBCp6B0ZvKoulX9YEeiDwhsJA+JpmgiFH6+T7ALqn5bz
CENbDdkt0pan+7xW+ncrGDncBmE5NDJsX1LFtJanPeqlOFvhA/NIJv5lwzt55tv5
02/6wTa/U9IU7kKSVoyizlSsGsppHLvfFG6Vc8+8Qd2xelvREOwBj84ifwHJME6h
VjPt19aRuwxtBzG+SQyNooQiNEqmcZkeG0KPXU0fMVmN1FhsRMg6Tl37KOhpmeun
OpllHI9K2dgPUxzpZTIusLyOzXkW1xXCIsudBZ3bAnIKcFvdDNpEvm6lVDsmktqm
oH8KQh5lfEg1KyYcbYmF159R5U3J0YkULhiZKWHVATE1MPoHpSfo2zycsdqidjBV
YMgWjA8siomA4UEaQ7j9F+5yE6lFgsfUVaH/vo9yEAACelgomDxp45uSw5oaMiG4
QOc8TuwqsvvLIQCMwEr1vm9vZtsHDx4l3ML0G7ue+7AuYe8LBaeEuL8blZH2n5rs
9cvbKGYVIEQKOsePx30MHFsaLlcLrh/z6QaLc3UYNc3ofVAffNRqUuaRmxXt/INM
0RJpfLcGpiOtOWI4nco5P2X6sTbDxI3demxHbJqT9zdwnPRA6FzhN8QoEChLRb4Q
L5vFnI+Gf0fssDePwRNJJIgAwGLoRjcvwY3bqquTSWlRvXAWEgH6TnhXuWmd0HQY
qu3dMXEoRJA4R6jldVlgpLu1tadzdlNUEnDtDW0/4Q4FGQy3+VaaE4a4Ax9lihYK
cWMoaHML3NnWKUID4Pa6xXtqDqdOJVkeVTmoZ0PLb58P2nXacWcxqUfNVHvxkIof
m4aFZfzIaBAdxfAJkAptvhDvguHw0/TagOEg/z0mKvU4TespOgPOJAebxmqv674n
wxBeDHWMcVf0Mif3lnOXIEu3hhDiRM+rYKi/CsEhIS+kbFkeJmSVyg9X34m+dS2f
QqSBDZ02RXr9aGkQ6iMRbVd6kAkzh64QWel56elmaEpNMIo5NKt723wLLI6B5kdk
JKnYIOQukWUrHExzYIc14DEvwnWfqHuVu/K80GdbY89sn6TaHsSD8stfdDydCbfl
DVMyKIPtwqZg17qsNZ8jKuO2q8hTIJEhAJaaEcSATEkJWTlJAtQaTS8mV8+KjsH/
uaeeavjR/PPHfUTMXYdO+E7uRu3KWDy8YnvDDpN9MlXLE1kcf7bmhP8MWLfPpMgI
UFHu6ueAMsHIE8eSTZZxqNO6osskmuj2DdLWh91BmL9pGZFXQa+0t3KMdPurrmAp
xlW2wbX9eVkCpPXqwbXr9tW/CwHoxeLfO3VM4XUBc3t2ZUfMM3qK3b5dkXZIPQpH
Hn/VSEYoV/UsIN1JMhbm4xAq3rMuq0wo2oLQe9Hr/RSn1AD4F/edMLwOAs2+5yLY
eQmnCY421iL9Uxmcb9Uv6dvnTkopqs6UZu4T/ym3zLSj/Fmotz3ZkU+fGSR7LhQS
qBVfUO/jOK70lJXStQQUBkY3M7qrp1SDzGg6qVPRGP+U3Q1aGv5fWLsboR29cXeS
0BXOi3ynvgHT5wtuUkGZ/kc3Q3ssay7OZcQn8JGOhuRIRXmnMSFg9EQnRYyNkiYk
89rn2DRo8xeSci/Yrk3mPvKHmhCaqjwHzBoU/vDKDyugJaGCJeyZC+ZmI6o/FD/P
cVm9bst8sC6HI3LzoDddJjOc+iaY88m1Uc2+bLDo2Jgfy/H8RxgnVFO4riL7ex83
+QgJM+4lA+1Q35HX4XmWjLXRT1W0bd/+JXPN0BB8r/uLrF2Vao23QAzSkIDtL1nT
cY0kB7HY7429LuTyLULCwML12l1TskmULF1EM3qL/H7LeAGp0xldKiWh3KVSHUJp
KOcrcSrePOnVmFjIjA1m7Ob/CQ5neIF9FhwPHttU+7yZjprLSiRKBVfj425ZZoT8
pj4nUnITOEnyBegWNsWHKOOxnMfDVZIH5xRYpLbQX0WwV9kX+iSfXd71WaNdfMqy
VPV6icF239e5jlhA5L1n4nEQewr562+HW47cZ5BznUcrCX6bcQF62enJ2Pb2I4hA
Ln16tQR6YggOyJ89mfknjnf4uKHKg1W8JMzGjxLPCVnH/N662+qyfDX33OcrhkSN
8zldr7sK7vIUW2bxJBkAcrBGjk9Mt1WqgdNk5EDS1Pn93sA1mB3iUH1rZ+7Eyy1Y
YRizqw161fIwQq5knQY9XQfvb+EhdZYUinqOlW/mms09sktvW2CrQOvMjCHd/iMh
IlCdfGHPCSo6JZXGPgMy4SVrOwmSBOAV+CG5F02nNuEpCF7uJV6byaihMl50Xlcr
SKktSGMdOomSZldCXOLGeHYdx6tSE4595e48f3FNy2ry7CZCeUitGvZGz28iOSUY
24OfI+UoqRxnLeaGxC7O99tKQvm3XVn4dsdE9SYvCDgxaH71N6MC6Wtx4DiiE0hs
Hl+IE/AwBseK7ImaclGrhmjYvxWz1ytZMRgqZpMCszBoHsb3usK39yRV6vWIDfg0
btHa0fci7DRyPlth5zgm4TkVTJBJJqVZId5z1UA0+xPLXusmwa5V1S6WYtLGvXol
+l1IsFBt1EioJ3vW1bc95dJZ+XirodO1gEQQHmLAkbV0+g7nKBshwkpakY0YQcaE
Rce2iOI3B2EggENH1FUbFZcvgO7EmDbHem397P3N0lDQq0mOJxjOiEBbMGhoHso7
wIDOy+1SBkscCDg4q1ZCr1dWGiEdxJgyVuxcVTsm+6wVPME8L+KCUHrq50xVZTJg
fNy25b6Ljw7YYNuyhLaI/S9hJTLtnbHeXK948ZAvLTpBznijCNFatAt8aYBJtcLq
iyHdSPJ4F6bKeJY5oc2MIYrAwuwGb5UL9U/71gDBMj+Lf9fT+EpqKFxZP/nIRz7r
T4S2zP1a+5KdKY6MF4Ybx50KNbLspuJGioz1j9hsuDrcmzPdRzypOASUTxdQidNm
/FxlWumay9E+uXnYF34jZo8s71JE9bYE/GMZbMCDVMkZyE+iNs0AtTLM73DkeTwy
PEkvvN30CdlIBr0WcC7zGnQwvTJCE59BnX2V8Kw/oNpfa3ChqZgzxeNBajES4ngY
bDSQndcSiCU1cRQR9kAeP3kK3xe4bIRGmLoUPsdKHA3eNGFsdpQxI5lu0yzb0nHN
awgMVNfvJRN9WJB1C6caM3TwEZ1XyyHN85zOO6ByCK5vcUfgQxas1PNfgnRZuZgz
t0GPnSSOIHOqHRsCaG7CR6m1UqypGt7/fLZfC8noiOOA3v434SOX7GIDxhSNra5o
S5g2OTT5VWzdbTQ90tM5j3XInnoYwviCeLswFTOsQhRznKDR/xSzNiFs3m4H1kjC
32Xwim7FpK9yRd99A/6sFGKq/lkK4zlSvX0crGU+HnkJb3OuS81II1+aQcIJjG5B
6n0gjOTjl4pDIeNSqk8SgUKKZ1+yRaDSutNY4ywsZB3nnq3nKTCL4MEA+UqBsTMv
2E32g/T+vuyzxbCNfo5W2J2dX/usrRGmLmktBiveZF1lKPcKf0gusAdcxBGalxZ5
ehMmlfNMvzGOwV+50myl2pEiEwTLUxQ4JFXSYU8bhr+zWTMMH9OjEr86MLPMzWpa
0dZEYVtmNlSmm/1+NFS5UvFS1Ri5exGuvZHHFaYkOLX/wZDODy+GfYC5A3noPdCe
Y7ZOnmbBmlkH6F2HZ95re+7qNy5Nnfftka+iLJFEOFWLzVZMhR8BC9ZBBu9zJ7eE
JhnXlhgK2x1XJ3sMoJsePYVhA58ZbTwZPGLMm3HQ9HUlNOAOa+kccDi9j868jOMC
9VvIWjv6EwQFjmw1cr5PvSw1UkQkBLWwDCQWfwhPMWIM//gtN1Lbapz7vSHLLkPw
XvwXJ+ND6zOvUHcE/nuiAbdZ8act6r0+qpENvI8SgD0PdKLffzKp+2wLIB8qnvoG
p77Fj1qdSjR/WNxMHnNJ6ilVKVwdUm2+BW8+hTI4cdqu6SblrpKhtCpf/wpRCGOH
o/uif6/XdfjtUZcVY21HIDrRIg8sGneHOAvtGLa2hgjPwIwn35toPRjYA0uJMO9D
wh7e9SBd9+WIgJPXuAZLBtp0WDmSyWq0IfL1wKbzg8ywq3RcYw5t/tAXAu2EHXqY
f/jACcgVjAPv1ikoGvIYk9us1s6cWSlQxZyGzj8sSZB7DYanBtFxN7pZp7azQGGC
2D/v3QW7EE0xKr0NTHRdk7OQao5jbfpH3oLv6sRW/zKeahjbGYwiUhrZefl/BbR6
ToTnWBBCcP/H01AKI1kwdtSj4NFPoAU4MbKoSb85iYjraeIqOjaTpvw0xGxAWSca
pMQAXgOfS8gZ6GTsfV+J99rO29wM0NHuE/GUKuWej7+OHxqMFi40NH6A1chy+MYI
z28/+0kMf5VJVCNuWnZHUqvUv3e5OO9vsn6z+GChyBwGvoQvpfw1mFdnfHO9bya/
xD8nkZTrUH4AiIvlDlc26F3DmZ6KAKd23dWFdJMoQcAKv+CvJRcO97libX8Fkb/Z
hhyaGKqLkz/TIkKut4tyHBTCF9WeN9j7gDeXH68oTlDQL1SGBNoihhhOj29DTL9i
Du2p6ERT2eV2U9cPmQVAMd4rJGUoCZVN6LkUPVV14/UHpaQkT9pir6EdKIoKpE8f
SEo5w6b2J57C6mlnLmhk/Aiq6Up0geUjEnj/X7LD6k7IHTw4MGNq5Cr98Cp3s5es
Z3apKYv1fl36Yqj1pw4YkkQ+aJ563t4HJM43G8dfX0qSAZAwkgXcrQLTyt0vQDBe
4q9rO+sYamDHozcSfPkmjFnVwQC1kTU+KXSJy7sP24WknVAASH3k8jgpRNkJ4LOO
EQu/cUX6Ke+tkdYyR++ov03AAUC38Q24wKd89TKmcWvhg3huSQSdwNjc00CScO8i
SxB8YQ+6NnWRG5IV/98V061e13iERWfvj9u2BgcoQ5Oe0Lv4zc5pv3RamsQz8I3U
cpLM+c6FnzfjXiWvqGEIYTq3uw0E9tA/KahdBhzqpCu9BoenCxHcp1sxMWQ1P+JT
4rj71NpnW+MP2drhHhASgBwnuOzrDn8SCdZPsKWcaCOH3EyXzmyw3kiyNEg/aLaY
8HjvQ1Ne+6AGaygCG9HAboaz/jjaaprepmds42CPXrFPKRdNWZJJGOtBa1cdz9sh
ZNMcLBqTAIN9AFQphDppfg==
`pragma protect end_protected
