// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:27 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JMYL7/H/ssAezXJRX/P1Qmb//imsiaasUwgSCN7I7lsPVjWq/WxS79MNzlL87omM
D4DBIElhv/+liqQRGUSkE1D9G/otkvS8azpyTU9AIct0dQjvi7rkKyf0fyoePi0j
HeO86mSGmYwsLCJBSuisNn9lP80Ocq79WrUy+ncioMM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7376)
he1jDlrgSVaDdPQQr2xuFDuKjFi8vDTdQHr7RU29f+JLBzmQRoZsRRZAdem/eVdC
4Lkr93rJA7Jr2s76g25B3iPi+AZRlOIPGQtcCoc9bs4jUrqDkAtrQS41hHgheW/I
V2bcj0LQMLun97BN8vhst80ZTjP7Hj1VpVSHqMlb70gcxW1Qix+qn4+X1h1zgUeK
0MltR+TqVT9rfBrwR4f9uyUwVCiCF88OxMfmDzh7m5QU6a13gPIGx3y2Xu/5qSdD
MyDmQpRrZfm0HAoDFUZaAeXX23QYJFxr7YV/e0yv2tYN2HnFAY3puOlVugmdiwe2
PyQ0MLGG6BdkpkyDrudfEOLc9Bl+bRNnccR4Y9HxDIW9bTPq0dwfuJL5FcnyLhNe
A4Na4h+yDBGkuKH0N8W7udk30wlplojGll3iBi5cSKOE1en6x95x/VBKYrGYuG75
INwEIMOmhwdOF0EPUC8EFmwtkyoMKba44/BMiGQFPggV8+RZEjJ5/UklLqSBKqVL
sCvd8WMC1bUivesMtbWUiFC3GDjD+RHUPlkbCHMrwl1W1v1FL7iP3EyjSD3g3hGz
tvFqD4tdDZ38mcBz/qT2xInUeXzy43Eoa3xGbRfbNyZUemVI/X2fGK4SBmUFLJxK
CXP10w1bWwv8gfARnnyjWAjr1GLPHDGDTMK7SucRhZDW9x9+QVKSITDInVQ36w/j
nVKDMhQUMSY+0A37B38KVLFE9uzQZRhKAhM/Hck/lMojkXDX6uqUhDejsUhN7JAY
kxv0A6eLjNTrfrpwckkQJFBCLdJ4ug1+lWCDjpdgiMvBSEjNqVBFmV4xqNBRKmr3
0IKt9wTWvOvHl1K1Jd4wbitbP1cXMrlMzNS+yK7spCVHikjZm8C1RpY/hqZ7g5KM
LbB/AV2kN314rtil6qc3UX98usGxdloqTlqIV6zxpOwjuVUkIVS9kE6OeduRB/iZ
LZ9qOLSWYsi7O2KBqL9k+rftzHWopqcvs72r3Qj2M62e6R2IrtHJnqp8eOeiw1xi
ROIF1bVC+Cwvaxr78ThlZJTydt+Cea9DQHPIY1T55CPEIrI0Mn14aCJg3kPaLmcb
OxmGjw/Zi55vEIzgTQV2vASzJcbYCxJzMH/Umd+AcjZPueFVuP0xw5WWMWFsxFGB
iS5jEYeRswH3NFIA+vYYndj+IR8YcHOSd7rUc4atrPvGvcg19ngxBJdHgJxJX5GY
2BUow0HrEq2ZyMvhNRnZD/adiYM9d+64vHPnv5KU4P5vBrhdR3R8y16HoGRFw4/D
WuoivTjF5Npw2H0eKs1A7gX76emi7jAG5w0zal1Ps36y2JrFiDR9sJuadXwvBd5w
UPJnV9FVRm+0IvL6n/I3rZdSf8bAVuVAU8ezuz7HVwIJieQmbFemLj/tsDAr4/tb
ROLy/cbMzZo3dBGoBX7Kv29MwR7nqw3pSAo1WoFVRYxAOwncqrd0Gfgj4HHJxn+K
JdPxuwZo4u7dEhFcRNnZ5q7RVI/yDgOfvQNsrjspwG/peHIky9MHwh1DqEI1fR4Q
nCuqrU5hMP8hVpIRdzlvamN4ma+i/CG0+SDntRJZ/aJu6QCbtjHygebhNZlEnM7r
RHS8dlgXtiMsUAWhkY+pDMHKIlZT0zy/CwAd1rWz6A1kPNm3zHgCn5hCgXEQlBc4
iClKVp2G+tSbVSjaWB4mzgbIN/dM3Op4HdEe0k2U1iJyInDCnL905WFgTOFfc6Z3
dbVO7DZG+p6bCRcws974uWr+dAZyRYfKerPrig7Z4hZ1B8BQiv98V80YiUCRJ3Sb
gu4Q4TfTQWNZIEQm8jRV1hbo4+3DpOpOwiJlOmoqyMpUS8bZkyrRi1hVrfDsmt3V
5ZCBi/fd0+6p6xs9XgAH9fPWVo4HbetP5Q3qgFUabyV0iA8eJLh5/luJT1NHWPZA
2rebUGv1hyqDYaxDg1sEo/q69rJSc/pexWULAzl5QWpFlJlmdgcusVfwiEzAH0nT
Cju4c4ngrGndABMZzBYxfMMPBYyAcq/hjzW72a3wqsy/JT4G5d4kGp/FtxddzGHp
HB/iUTJmP2kAlKm8EnU5w8MW7Myf5mAbE60ZryskxNpg7UlxW2+a1P9MS7PS+xb0
rqxIbf8O1Zpu35g/6H3TrkZf0y48AujofTBue0OJpx9eMiJx3Dc1okjKWQmSgb0y
0DL9hMi/QnQyHbiSrsIS8OJFwINR8kHEuLIUZ6b9LQ+FKB9IY2tpxI0o46z8EQ+1
0zCHTdyikS+xFPUTG8jnQlTn1IOUF7nVI2f6wANzNvZC0OL/j0uHYQIwW0G1DwES
YqjmIPSok+e+yNPhXFleK7FEx4ntrot7dWfcZ2qZzuWdDXgNG7lCa8WqF9SoUsgK
cQjOk2HA+M6gAlvBVpzC6zYlYCZeFFtajjAuqRmVJMK9I+Y8srdZgZnk/mSK8ZvE
CgZtiu1S7ipAqJobEcsgozTZADSLFAbYO83n9/HqEzxv4fK1jvi3Eu6BoSh2LemN
cXMOn1+iwIfKlIMu4HXt4LIONRktnZ8k2abgca28XDbX4ptwutSyzeNyFn1X9FIU
GlCOwsuZC6WmHzUOA2piG9w246lUBOk20TFZwSIQhQ6eS0Nz4Ui9DYSU3wDBqH8y
4eDIqqOyrQtE40613kWue0JaK+tjamBfmG7kHoTjnpa4Qf0zy40ijAGdwIHS4Nv2
tmWzJI2/BMXs4CiLhy6v/B+1neQVrR7y30BkcVnWqFgPRijKVla5iiisQhOscAgP
crYWnBASfjEAif7zHF65v3ov9S8be7F4WRHwXqsHVtrhhaV761RXdlPEbkxFQbm6
oqRQ9Wyn2sLtndwzdg18vw9qcacCNMpXiLMUDh7xmyR1VOhly/K+d82PVNAspyYG
w5VA8TUycb+UOlaul+S4n4An95+Sgl6bDe4PgoylnJjRmIm8Yp8vjaZo/R8g2700
4k+bA2HZunUhMMKBLpVxpltSxOlIIKoyN4h3HDqMUld0M0NnvnaTSifVg1CDhC9E
MkaAWXNZ4QN0ojL7qK0C//BMxflvNJM3/nK3unYddXeasxysjskLJK91djqRhu7m
YS6lEjWsAh/RQTvQjGi3PWZm/zzP4pBI83V4U0VfQaBtzcGSa4sHfBwxFW3AD/sq
KN7EM4pOh57Sg0zhT2+Xa0kWzQ7lmwDztPG96XUVkvIUp8VRikw85hUwntC9lood
mnbI3mHAwyNduji6tKYptbSstXet3VRqEtjeCSvy8iVwj2tBxSfWcVyKBpu3/6GH
B2YURnwyrOTDy+i0IKLMS0x3+JefEqKQ66kg9oFeNrvzJ9LB3LGd/vWQrsOzJUcV
nKR+kzkTghfHeQyWYhRK3ZMcWopU7eR8HYEB3IZuUPNc86r4tI7LNCfMC8k0FFit
x4uppYqzXdM+Ld9n/Nmq6VRu5m0ZtHUJGmFUtDtia9bHQf5NrvIz4OQPINr0SEVU
C3t0P92xZ2gWjPrYV0SMuOEzks+PaBun6/RchMoSpWbQQEJ2Q+Q0Kzfozuc3NFpq
sznX1fWYmNiGmo2gkdV5cLqBjyoPbTsUVO+uRh5Az/nAuAu6wV9abGpuVxZKkd23
daxFc0ssLtk+8NyWnww/VAxLTLRPgAQSfq6SPio1YEFsWQI6RYVnKddmBX20Nfd9
OZ8Do5d8Hb3ZEdygAd2XFcTIpJtva98fpgd2fTZwRh4F9Y5rLLmErkJyZ7g6JdKF
scq+6IwJAL/xGgxB0KoMwymkUHWB8WD1cSnNDikQO+upcgztgGBXITibPbhLWQVO
Nf0qEwNO8cx95yIcPiGafx2DNcLFwcx8MfagQrf1sAydnZF3JHi0777UQ0irCZJC
AlWEeco+A4KGo9lUvW0sWMawFFk2LzorgF0m4HT8Hy08ssUDKiyFkAFf8kJo049X
4r4aJJ6UIH1U2TgW9p1mk/bOeht9b3bhDvE5ybpi488V1FhQ0n+KcWCIGvBXMeVJ
UJNblijXf34kCSrdqDSifsqhCGo4sMS/R4BW1YFG0odO01XZ5fbIdq+aGy7Fu931
v/I8BWYgDj6rKj43tyQ1G8Px+s82JBT7zo0DV3Uh+8OfPQVriwc9hZSv5SM+VbLI
FC9PznllbYjjNiWeCnfDPE8Prm0/J7CYoanQxu7KDKxbQpZTkAcFaaanpu8Stdwi
dpIfpTzlBb40y8aM3BXxhvCMnLpYwb1G2FD80OEfHEKTJaCHVSXBatqSOsLhZcMu
rVPbBGKLTkbOOiW2fmFz6EzqjZCtoyYhNUzQSIESt4GdjAPosUU6SRM53oD6JE9D
aiq63YRtNulHF7qqlypGjsHoKUitBoeBCpta6rSti6Yf5CUSaajs5pgkIlIeoSCi
qM3WshnWCZlAB6ZCpnR7vWhpmURm65nEo/5if1rcSrgzP3UoMouIPb8mt84Sx642
oiseAU+OWSdNXcAvO/Kqo11Q9xJpE5bywAzR+MkRlciILQmc95SfffH8CywjZWSD
3PRQYuh1CTp8/WqVnFVCAl4r1gFPdypNRGhmH4lvASpKQf3mYDHtByRba9jfT64G
HA3RcUFrYtI70nP2y2ZaE81j1zJQfhISmeK0C1gy+MHFuUifi44MMI1erNKhlFGw
ohayLdoMMP504iAM45d6hkvYiXN8koJfI9XIi+/9Z0cjSAEBtayhUBrFzfytuiz7
lXyUpyl7R5jELekbgJIVAfEqtFubRJ4pLMW954kivFCevLMrci/ILWDptwpRu2DU
MDAv0CzOuQ6P2m6YGf914qxilR//mct911KFfpN8H2zs8ZxgKw0DIiie/mfEDG9i
+MsJh5U5GOyjQl5/OI/LHV4Vo3YnCjCyH1wZs+FMS3p0ERlseZ6VpkXEuPrLavd/
wMaggnKBqRpwpubdJSen9OYydayHqTyagi2c/9yA7uXgdwobDus8udqWtz0BPrYr
8Bso76ZqFggLPHGAFIBVWLF6cT6mfgPcDmv2ifOlTccUgHMtiR7NCJjx86rgR61s
BIpNoLiqV/8FNMp5InEgpCydifgyq9LT8sasLjjtpNKOyr5gZfQKzeY5BEVpWx4y
hCycx1myM9RufLXvreImQXRF/0COxWgVy2jmySggkB2EqIXAarzyqJxYSKqdtp/F
TX7VARVxxX7itpsDlrELtI9PvWpyrbIQCuQh8JYWLGDKGSg33OyxNGPhW8iIru3e
4IDgovqxhPFkVO/7NmfAz0Z0Op7FHx/sPEFdzzVH2HtwqGaJSUKvBKYeKgN95NP5
wS2nnsq6GacU5tLFDDYK6ye5N5t3qi0gna7yvRACNVfat68nfEeXjwmHjwo/QSqB
RLFo5EMCU8vAb0oef71L/OiH3KGUTeVaOGH6nCIe8c5jREhcKzm7QiJpycEv/cnu
zaTZE4aJbUy8vpkD5bnEjkmzhGjSUbTBc0vh9N8ZKO/dmuSjxefkwF4z7wd1ZgPW
S80du6sTR1wqGHNsKP7hnAalsVz2lIUu2dAVn/gqlIqB4mS2nAhkcTz8ONbsYb8j
YLTN+8PZKl2P1JpeU653Wi5FbDoUaM0n1mg7HMq7xRvzg550gYAilKCGM55fOjRZ
7TrJk1xhBs+F2JGgpcwWpqeGg0xw6EPbTf2u79Iku3AX9Owy06nzZCxgxkVykKZI
jnTqSarstLLD1AdARX3OxHWwXGflQWqTV6qkOScKOdJnN2fFxdRR5/LALCKVN/GJ
1mI6bMrHwRkoGU6+3eF8L7vFbMO3K+S/VIpEfjgqMvEy6GYh+8yhccQNrPFqdUVh
7B2LTQ5ski97rjKJH//YSJ/GWg70pR+Sl+wsonARNOG+4l292ai9eNbCWJOW6r/D
HzUpRAMr2avDB5Ixg23/5HGY6zIrrM208QHu3c5JWyiivdSTn9ifMZPoRb1tbDlO
fxqKrxL3djneZ6X1iIhnU/rhYLz08dhIH2CttvT8QJ1zjLYJV9udWVmRbItjViVX
I6NCIqHzivZIBuoIB4jslAgWdBtgo+oogxNcRtEjzVSU1L5Z9JbewNBVhD1DxK7R
CPk/jQS6uJ5V7hDYmC0sqnhU1LmRL0Qw8qWlYEgMwjatzf8TgnGQ4EnqnwYpq33a
Pl7xCB+3Y513iLtLUnw8AjOoxT1yJH0DqNrfbkLUhpbcLtZKLRIeVbf6jwxH5hjg
iOUAKwHifGXONhqHrf+YMw5Nzo/oOCF+Ne9YyuzuOHftM3rRMup19QgrkWo5pnsU
OlRujh3bYcAKDDd0Y3qem2NtOwUvtnqB+8OAo15oJnamj1bzsWyxJyhP0zh6P7s4
osnfSbMgrfc2YWv6kyfiaVlg0roUjZMzf25WxO0Os+2mpDqpmRbbcKms9vZUGIH4
hmUPeP4AM001hBxz1gv9KMO4Mx3iXIPIWNdsZM2u+XhNF3d8aSLLOmiAT8nKApwV
GXDRKDDe+lmiulO3FLGURyh7LvPAC1TOWYS31W+FhPITlK2FmxG/bJANYyZvQbg7
m90YYtwMLfyYT0CM0yh5RtmaBa16n9S4VaAyF8VFOafh01Pc0DvxqJJBu0+xKZI0
b6g2oQsMkts+rDI9iImfbbnCMn2DvRXJgjwg2rE5s+gech5LhHLQXI/aeh9i0P0N
RagV3ac+wvR9Ark7iefkx+feYu8pVYJxt1miz9kw33chnYeJ/du/db4xn42UO+Eb
4hwcTBiWZd0kB1fMywofKrCT2hgN1QDJN6H7+Dr8C9grUIgE4tw7cyAl4f7fl382
UJk3RL7rSvqat5d9XZA6PX4b0skHIx5VQkzoCU4RktSsCXXZtmK2e0BwIgb4V9eq
jmTrIgUNaybPvoPgbkwSiQNsZmh+zwcLjffClPLLvTMmtsbjZ2943dJPJpqC5H23
SYAne7hbYaJ7ohTVDtbItQH2iiJHGx4uhAsY4AyS21qp/aAcBQQGKJLGnvB/Beea
agtYeaKS0k8U97ztdssWqHMxWC027PYMnAfvLF8oWRxElmb40M3kP1ZPySXZFJ4C
Q8rOVHtcwfepe88e89YmrDwZ+4LWLm7wbzJPIT93XAIbnroBv6yGw5IeZT0x+Y9J
ZcN+EdAwhyp4E5pXPF1oTornyH7Z7zipLP7AzviqYe9BO5U/s+JTe6CeiqoDfbt2
GGoURfXePmuqo7tjbPwEeDNEST1m3HiLkLlk1M5KUwAaCtCE+ASSb5dMTkDeOJsl
auygG6qORf2BRvkqqcGqe/5j5ld8C93zfao9wbSggx1gqa36PwtTaVLpkz75k0KL
JjS7sHs4wRElIaC9UVYTKczFzi2MzGtD5dSdERq5+DiIaTjraovS5wbyzarq5BWD
brwaPPQejsurBAAuHzhpk4A6VYCwYH3gUoFPiaAhV1+5/3exWhAkzu7T24HWaA6E
+nFdQBE3P16W7ijS5esG0J/gUDKYAGKnxD1dkOXKHkgdMDYnUsxI+oylkO6jJK1K
zm0Vt/i+ZCtQfApp5wSNcgj0+986SKYOe1V1UQXS4qPuZO0WOcgOVHYW+N6sZgpo
i1zrH//71riizEFzk2RQWAufu48Z+yNtxfazSs/0gIHurcE9i/QKQxEtFoVX4Usn
vRjyTiWfq1FGq+vnTugnmBqn7g3cVUDowt8IPGx9CTj3qUfAabIp/WpQA6oUzzzG
RbrEO8Oc4ak7J/oC54oYKd3ivlFbGAOT7gdRRGN6yeuXSNgNsvxkcYDQUARb3Hoy
yfdxiohx8sGSOpfzsYTclrx/VqNUo1utGae3j5adAJ8f0HqoGHxheUzUwetslmnp
zdk6yLBU19HzRLZALgE9zRKbvxtcMsBkh6u8uOuhvAEYDPopbZ+pGE7iB3AzSUQA
XI/rN2qI6TXRXjlYOYgQIBMxUXrgPyHPrj01UOQycEVuZE6ZWVxBKuGrdI5yGpxo
Yujop9/Pguq8B5AK5+ovICkGSKAPKu9c8FWbb3w0dr6JmKal18mF6RKoD4wmtZUi
uH93GciTzzV1E4vCFQds9ZOsUNEyQYGsvpFPgW7Nv4n9HxPsZgjo2vQqQD3GSvAZ
zgiNMEjNgbwXbYsK9nzTX3I1NMB1OtNCP7LQWCduI4uycaklcOpkfM5l/cdO3dnQ
qHIeuaKcp55QEXzUXSiE+JuWvAoqWmtsvcYQ0WbGKZ1XFEvv8JMU57+kM7dz6MQg
sWvBHARms68z/yWaiby+kckfBsLP+8tZDD5wkKh5G6GwdMnnh3RrLzwOGW5I7+07
G4HQaHRuBFuoG/SuiQvUR+mzpG37KYiDXE9wqvnPxMNx9+eBCgeqYHCmtUZgsQpl
adhHNguohiSBz/LYxVCpNZc47A9haA14aq/78ce7RJZo0UWBBnJvS+9G38YscyC9
mix4+csD9leJgvyWkebVpOjZQLlniKdjdQY6vW1oqxTt8Cuhg6ZeU+WzXcXT3stc
EIuFmK7ZBAIEnG6w/Hn5TyjoQFFZMmH6DYCGiZpOrhyMUNsYwU7+eGCmOR+32se/
oatM3ntks8oSa9r81a8XAGYZon2yigKJ1RooGvsVEqIF+xQjWfsMMgxRPn9kSeON
2gxXn74NmS1YHJ5EOvNeccAsMpfjXn5RfjDsyRb41u1D7Hrj1/N8b8Ebuqjl5pCQ
fnko8HDCMJYM6WM+soncWIi8T8tUpkxJ9cYKFMfD0yRbSnmijkvkhd3PqA7KQ9E6
4L8MpTbU8/VqfCta3TJxG5eSxPJY4SHU/4fgKwVNL7IZyzZMJA7dPtPT8n9ECE1N
QyiAV9eaJ2dNpyRT7DvGG4ncUOlEn9iIs0830/ZLVGtpOECYaUejlrKw2q3VbxMU
dXwzCH6FmCeWbK/xtEBOMw30gUK/nl5GZps04mZf5Wg9xDO4sBenTXAERVmxOdhz
d8qD83wUaJlMZFoq2GqMUcwty9THdEeOqsSqfs2XGznCu/K9rYYsOtk5P5RGeHIL
+DOeyeUMQSlzSUlIDuw4kt9AvzWpW+/3ooymJaTU2qilaK/9tY+pynmHrjgoSV8/
yPVkFcSijufakamyucC9s8fLWROWx22jArhBqK/qd1Qi56c5DF5veYIrWHEWjedM
Hht0TZbDMfOYMuwGPCVBLJWKkhdM6UoSReul7DCXKv0MIajaO4KBMGSdDNl9kHLz
+xh8tQR8YtHF7wzo0d2TUkqQXniJv7TpN5TaRS9iJTv36FvC6+GD7Q9Sqo5hMf/n
sa0LoxmfzpmRDl2NolkMH+XvtgYOH0e2hAQhn/67sPzt8TIcSNBOc9lPFAcOSxRH
9YLbfu4wpK0QqCqcwo/hjPmfB7oOVQJ9ySbqndEvy219oA6Se4dpdlxnamwFjP/U
4rFo6ty8LGqU0AqYaigYXjIHyh+tn1yG1alrrFbtZtdugqwpYVNUUYmugo//PDbh
Ctf18ovps79pmVHmwpNH3edW6fRP++lP++00a8WWE8SkVzbvQg9yX8lHa/g9/efA
vI+SXsChdcez7lVSCa5F1qMlRhmOLCfB/wob/z45EDmgdE4wjRrrMh2N1CMYQdtu
zB6RvL55MazCQHmUNDfGHqbCGry2BYi16SE/5TXs+7tO+07SmB6ZeNv0lFq6rB/c
cxF2cTSY2pkw24ZUNof95Hc19mrz6bL6hkyuOtIJD1nSg2yZvgLYY47b8ZprizB+
6JdFAWYvCyxB/HoFKZ8FNw+kSvvHbwjv4+Nzed6F0SRBGwb/NkpmDSBvguI0kk8x
IGeqgDXRez4dyy2e06/T5rtflEMkfq05BwlrLB4oWz2G3UI0lIkZTSMVHIpTY2iJ
dYEPFp1Tydnx8/sizo8OXEOr7Iv8sS+IU2fDi91q/YEPX230I5A+aGBGffTGb4B7
JGPTRnKYhfNbQbf9LzgWKcty1ntIybYmseJP9VkxZ+A=
`pragma protect end_protected
