// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Prt0pZzggPe6Q+UW3wPLgliKehS7nKYm/fSyCqvrGdg0HABPE+mok/3ydDSVJD5rSUy9GN/ZQQuU
ZkdEDv499AdcxvcdVWy1Y9lGvgwh+z0vnYwOCMRCiTDaw8AUJHnz+VYB2xm3D0R6rutVDbD9bLXA
jpmvrHJOaKX5oKpuAjRrLJ7g7fO6rZM81XEtR+ioTsvWWsT4k1tgmeIcraJtrCPAm0A4GdV2KurS
v9q40o8xcsaKz431v9j5V0U8LiZZ37LLsGTH0p5/ZnHTdAe99GmAoVP3VFJdyUhIPpSGaISGpaEk
XjTpKHq3lYXLgcMHpOAl5OyhWnplTOC/v+3p7A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
M9cmpvD+wk2t7w5AoB16Fq1bcpYt3JrRWL/njeJ6ztg15ea65l8FTv6htVNvc6o4h9I8Kv8OM4BB
5kOfdhpE9kl9gB3d8ZPV89PNcBn88OXCRHGoUa2cCnVKVslIECBUtZxblHwMRvSKPXUUR/E/cXMO
bZ9buhew7JTZ1YXYZ/z+2R0dDcK+ilXGZqam8SsYbmYno6xp1smd0te8UguJQZzQyJIQd0TZmmYk
9oKG8rAe6GvmHGBkY3fdvY5BNY0RUNRJGGcSc3puN0ZgIKwOiVdaE/KJrjdmiOr0n31XKu/QumKt
Y2Tax9PMG7FwI7WVnTUGJX+/wXOGHDVGVxuhq37je5dwit52vFI1n9OackdwnP2dV5WjdF3Zsog/
X9GFOB6XANS3xw8kDdhEqIvN5XWQSF93Xqod1F2sPCiLu8Rb/8xuuuYnvGxRIn57+q+IhpGWGmwD
xb/cKDsMd8xT6lSq97I7ErmIhsj4+pkJ0efQd7/Ma9wpbQRx08h2PeqVwrOqMK1gSA13Xp0y9sYq
+Xd7XGGXNOFuk7k1+0Xl6n7916XCT53sQq2q2+rhJCMjXC+Ovh8BdgixYB8VyU6rUMIj33MubVdC
rspwwNbNGCgqRxqUEDewo8szcz+kTrg/w5wAXq3oLfzBiIqh7nrsYdQpmEJovDCmnhEsJzAECZeR
3/fWeNzf+ux7REhnhCJb4CTwKdYddFgpiNzuIVAaPDPbc3JYJAoHMbKTBY7W9OuijMVEDfFD8eaB
F4wiw/6yQiNpgrt+IrShkyO4u2Yw12LOozG//6Ca1RRKbFchzEkf+XXAc5l98TUOusJ7T+AK4OWu
OFzdimmcrwHBx3ccLLEIQ4I/ffNKeb81whOqYs48Fuujbid1uaoZpICgoGGcI/yb3gaa9Uoddkkq
/r3jkrJcTqd5K2T4GKG9nTRQu+RQf9VKQKR/9JbtJbW2k5dHzt2ECo1Yy1Ak7LXphho9peVzqVE3
7Js0jwdeEDlnDWiQVoLtfCRznSKMLydz70Cisz5FUa2y/AwyPe8Vs9X6JtoUxNoL1ZKgXv5HCDsj
5mEYtrBFGMxcUlAn4kCgxEX6GDdoEwFzSrIQzNyuEffQUPRZfMRAr9P8p4uugpPEHgIYv4ymrYvA
gyyhpgSarKGaDqx6xiNTqoYl56WU6APU+CVQsKglJ3cx1EC9l1AEmPbQElNojPvUHfm5mGa77Boj
1Kg87JNrEM/8+RDm+M11+T+Y/YYz5QZuRRe25RYwJcG51FzyFYiW7SSuZileJkbCNl6t/tpaNugy
TxK41s5F70YflJvd2qexQw9wBM6L2soEFDiYRHhClrzkXITgfXUz48pQ7TqC01YKTmbWRbCKwT2q
0TvnzqNGOpM7h0ehEhc+bRVoW7kT8g/bhM36UISC23wiZvDKi1/1L/MvL3t8Z25Az+R92b0zBVaa
oPKcz14BVoDw1mAFpAIQJ7Xcv+08jqGJu3Sen7wr/NA2kd8X/keCYXZjaZUx5CoIfaZQxyDRPMUS
Q4xDicvW9JjEWKEACGI0N3n+J3sMNp5nM+dc3XHP+HJLZvDUdL2KO6whqKdlUkZJPIYxRoR7Yndq
wLAs027xYDPTmHmeAvEBpbRd5mZZUJODclPUn9JBNLm9pt9tk7qRoMwwtvsKR5cpbjDqacbzqfUK
+IosITgSM7DPWST5T1WdLri8HCWFc4gm7s+pSh+F2PPeSe0be7sj9URIW6/F4Ws3Cfm4lV7ziD7G
5M01w8RrxW0Nn6bE1QsmyahVnBeX24T95idZTOV8KdO2OeYT1LarCWqTF+S2jH7qHyvAU1JIfC+j
2CpLGcSqAxIbAT+zIRLEd4dJPMR2GOnE8HTeljQChzEpnSb9wrQjr9ForwKDYBo6VGA9vHw59GMS
tGtbfgucvTggo4kPTRcT5yyt3enjhkmneIGTj9ejJZF4lG+xnjD9vXBPQ+64Xttqczk9veDoky0U
wDGm4vvUO6qXhwfbfUQbQ3oWUUb7LF5J1kWRRwaKTC5sUGJGsH6o9dO+tcQGClk3sFg0MPHd5/vM
hh+46CLx0CGHDJIz4aFtpDbZ8cP6hJW/O9TnyxIjbrYnwJ+rSm0ZEzIiT1g2t1GJhMhczp32dpHH
KL85rm1xmR21Nez5nNpbAixI86ZLoAZRRqd10sEm6WuRUzWSiI3mogAwimt9iiHzwK8KdNRqhVXH
ynF2CV2bA1lWyhzIL6uPhFib4Km80+hCwRdKiJVZvOLDTuMUJaMHoHxuDoHflmjWEZSuVHAljeU8
Tf897F2tc8tOKEbfb4X1qhScfqyZTf1X4K+FpPPbkbm4Kw2tDSJo2P20VedYzcvmxKoMA3rDgnck
pqQHqVe5r+tRNwNKub23kYGjsgHpJpI0EkfZsDKHVqbWxC/bDxS7Q07UE++YdU3/xUT1uVeByiDw
N3yHKOxcdWirBzQgUr2u1lVjUMnmgHL1RRR4/x4ZJEzGDDYepmVKHWh4qBIZIglQyjC69InXthKW
iLLZOUI8vOipZdTOAiYwXGNRTCjOA+8eh4lEvTJbtsg2qrs8MYmbcXOZfk5+eN8JJHfRB6DiJhlo
n4rP9UEZ5G1PxSbBx8pBT/TYn/q0uNLHHL2D9CRZKNjcEYZjKiuBUi6GQLVZntPr4UmsBLXBsaCD
UIFdEH/5NjHdLpTGXih6c60YCkhfZ0cBdMUORpd/r8u+ErAtdDa/DDAlqSXhVgkdrFySeziVFUim
xfG2ArFqtJz8eZQyyusPcjtAMMo67aSzvG6NtVT0Df0TI0cxLYnLaMQJhYv4o5H1+WZt9cakeoNe
ECoLiCN0ZjwESlKxKGL557X1Rf8WxUJwzDh6Q3I06TKHJsIEs7JwPs6SzHZ6GnTsSR0AIftTJfz0
oY5Q7BViYjsWltK1y2xx+I/3indk5Qv+uQhNtqqxEsOuTYfCn57jCfZpURQphBiL0pUAJvm+x0f2
S+cZAgFvlkjc301uzisZilrGvm90jKm5PaVS8Lz6qO0r/8qXTQNDZHYvRZMPnUqhyy4DoFXabnFs
UbulgJWfzJpc/t37+1+k5m9NcQDtymo5Q1qAR9trNYEKcSjyeUuuVfnHvw1YObfPpB59aRx58Rv7
VJ7Erq7vQVIRwnll+R4//kODG1ja/iU+CW2Oe1mPwkBfo2BOb98vliy77TCeB8I/zjaKN+omLBPv
YTklQ4cIB3akq6mvJHYdJ8OHG0SmfvkFWZK0OKbxlJoXfcNK+7Wjb7j3AF6zhzia/TfiAKvoKWZD
t+lD8Zbguj5XmJFj6lwa+IA0PfKClaZMdenDjpfjXAz44HcZxSIcOKTtWMGulj4sDUIie4eiFh5u
cj138VeCS6ZwpFW4WsouL2PFmZ1MhYS2Hel1qqIm6o8fYADUS1+dWJ9/6t96ie8Ru57LXOXVxDrx
5RufAc3TA1Qa6NNpcNffbS/KmV73nBEx0Q+cJO8URho75tKd/eUtpWREwvAy+URWoq10EHD9X/3b
5AWE4ON0kbHn6RtNwMJX/uTpw+zRk7l1Qs134VkK6dfHilLMg6qF1HrsUlE1kMhZI9zeamxD7AWQ
fFDzB2waKNXZJrgE5DuQ9l+myikuSp4eQulL9jhPRdoH0QuYNbbGcQJRpCDdbKinAdqYTqKa0nfd
z13DP/gBU9xxfdTNbJiqPPiI98s8Wr1UUSXDZQMZ8FOhmOu3qf+muBqz3+WvrbvPAbr1QPMJVjKl
zx3/+kDc/WQFPlOGbjTLGSlQdjFcTaTPbl+eK9olBqIzSzJfOqMipWi1wax/E84LBZwOpDx3v5zt
C/Ti6Mak6PYCNSOGETe62Kg1xNGPXF7BUHdXNJEEUwUwAGHuDEn0jV1jq+66n5+N2t8WaHDsb8LP
iB2IokwOewmdBWQdIIzK5UKdFoI96PnsFqo6BqSnhHmKezXtBCGLucN34kNalKVT0Wzn/FI3ANcN
CmybcOPRnojoQaVgzoxJzl2iIUSe5Noghamh5PE2GgDhQMKXPNYuaoo8KBKfmru/WKAA4UfcXtRJ
rskl5lBWWBn1MApQd/ribR4TOj5h8rdLhbr4k+rcksAtcIlJtUmHPIYNXsvjJXALqFaBn1edlpJu
lJPCgvf60jDl4G27jJCdjB8ZI/yFGVmHVyChDCHM+915I5ZuBW61eahuWnCmYyqg8O2N0XwaSKqS
cEeF+dNC8kttzkBfDnOeRZfW+E0jZoxb3gFGtN1YxabvTdCO6GU+CC9O4E2fW08pwCYNeB2y6YFd
tBmZsBva7jMAalmfNYgrxIumNUXvfkRlecbLcHYQC7uDlciGLNPu4b+HoE01NUPIJCE/KOq8c5wU
DrMGtfimAA4O+emTFRINIMiXHKN58lY3YkW2amOik/wFHU3c3OAoNS2iPAP5hbmjhmWV5v3cRHUk
0NY+v/St8qYITRn2l1SRQOZzm3DxuQk4m7UPMYUWQcMFAsh4EaGC4QMBzPL2lwQwKfYlsrxkbCGj
sIw9FIdZliRemAXkEiqbWsEv0Z3UFrafBC4w1lqBAGQtg+HigTwRBOL+HDGQuajD2qdKqeiSuqbB
8UBsmXdLbmn4qD/H30Xl2NxrgwhPrTOwQfv4VM7U/NvPALyyU/oMe04lgxjpMKr+g1FF5D8AJQ0m
MwQuKwIdYLg9dttmbzoPhek9av0PfipC66NENo1l+mrH0qVKenJEssOesQzZqhQtnxCJsNBM+PL7
DsPHX6ExjRfb/96//Y5BlsKPCTqf8HiOmip8tlZRQfrEgi2mmFRK4c7+t4LTq3oEbnX30DNl1Vvz
gGqv8PeRLxtvzpdxE4lyVdqQnR7aCzNvyvnqf3+XOcPOSUo0WZ3WfT6H1sUtTIjDe2GFgT8tJpQE
vK5DxrG6HQWQr2lkkimrTUgwof5VL154TuRS9XN9iLhmUSWjitIxjtrgZFBe7IiIp2SQRlfMkuYp
j2r4mJ754bn4Qu+oRL4GPQctkZ97TnVPaCPj9WtX7naTixgxGOOGTCr27baqNgaBtxrDsG1CAE7Z
lJS7I/W/ki+pCOxo25a6LNoXkKhE8Y8hLso0gZCuswhm6pYkLZsMSdmRlTvJAUxZgznx7Dcl48kB
FCT1zbxKYppm/J5JgWySn6sPfl5q+AKfH1quNdOcq9gN9AteyrLtTg8dq0lCcIb7Ox39s+wEPJHX
cGtqvX4etO0IEcttZTxTODoExYz0FaTIzZAEfwOSREyi6JujLdM+o50gwKqK8Zi1AV2g7tdkmmYL
8G+MaWeIwYNYrE7EDQweMCOne8LLXjFA/DTm4SWGKb1ulzo8HCkZuT8NiVwzY0vC3a/1dX/cnLna
NuJpFfvdqkhOR3K41JknKiLtFyQZkTTb3+0t1FZOaaAYEI59q6ngDDrRga9V9dlz8CL2XBJ4fJ2o
pA1LAI9UGl93jh92rrsa1czEE9MaKnlb/QnoWryFBWinCm680d7YUVgAiLV/dW3tsoLpF1eBRwry
NeHI1ORDeRVi12J37L38X1tLldD5UazNi2JslfuSoh7Y3Vgq5JG5kXufHULlfNu/4ODTb4Ao3RwR
KUKqDs2c4aWevBB6SL4XIeIWSGBorZfaEa7sOhvTlojKrLPgTR++e8v2nmnf2oV4LyyQBzQQkJ78
yys1dq1zKRmqPYavod9hJHoc1hl2ZsT8xtj8ZNgQr8uJQjWMRx8qM1/6kT2tmZXbyzF1CKvgfLGJ
tSTasm9TLPa2lAk0RV2xuBKXIuUJZFE89iRSPfCcxtr4RmW4OREIhSy/rqoWyxs2955ZLYkEQbTg
m4UiRxu+yTnRZncu1uXLUaMj6mU45SnVh+48D67pPxZ7YImXezD4MLFGkCHGumKiGmSvQEb1XBOD
hd/+Giwd/BgGaRj/fVEvuG2l617rkNDU1vzW+nK5wSgbBW4+oi8omR5qBFp8+53oodpcEtwwlFPA
85d+VelUDrAozL4bVAr3/ldtQ1e6HUx6j4bfgvyowQtENqDT9jvEOXt5uQtyfNLeds5b+WKdO1Zx
P98OVg9JxeKoPBHRwbiR2+JWxnbyOEW3vOymKLjC3V4G7TqFlzl2g1dguc+RQdslmu2a31ImYQzh
LcWPU7jFevNTIOU1tTIqYzZgxa+Y1+geKxlXg4X+tcxOjaG2rHeckX1xpCuCYNJNFKFJfMaCrjno
R/Bae+bP+kOnW9Ov757n0Ps4/bDdqYeTRl9Ugpgn3Q5q7ug4fqvH57d4fgCUdy2TdGIgSwNNKDdJ
PHH9mP/AuIAk3M3UKt0v6NhmfXYkR55PXy6dOpPPxzK/MtqfhRQen5DmCt2ZRl3EiCeLXyzPgMcZ
Sa9xNTrlNBuXAHH6rioSjlNqg/so7hLC9EvyN+HX8NRpksUs3zIzyRrg/g4QV3/fk0HBP3rKxmO/
KNbUYYpQXcjVsUBB+U8VF1FIwox4SPmoefCd8ZdfQqVyHAsOrE1Vv+6mINQ9grC119eVVmMFCndG
Kh+QNUumMw2sH0IH4Mg50mIRz92qeXiGgKfVmCcJTwZJhXzKGxXn8OSxHMzB558KFB8KQSJATx3N
IlgXRTC75/I8qAgK4yq/RDPnc+lF30oVKByjV4Ud3p+FoGP864cBjJKz7L1KUobwsHrPGSHXRZ1m
2GdZkOxgcpzmkruwTZstiMVbFV9ESq0C17gtipfhPGDjNVFQbn091ApSWpfnOaWvISkwhxpMcqe1
Tx+ZYdpk9E5YCocFeKNk2WBv7qMT7tFioZJ/kzch9/DQk0afmkpV/n6owkLkconbQy/gOLWv0BY4
JcscxVN1zlBdcHPKJFZTsyH5w0Q8dRCXcSBwXO6yMAB3jB1I/5E5nJc+1uU2sMVBbn+dXuZXL587
BX6ysJSWyMcidSnnuEMkYk+8ZfnRaeYdA1qv73CXW5PECvTZCOpilZKO7tVXz8cF7gpBPyk8HrdG
xa73gAA5eEXHHnMbKGlJx0cExqOL9/K22Yl0IFr9nVMnjWL4W8tpBFR1/E3r/PTzaCUMndce5JRH
XhtYo9t5nuoKj7+BjqLGtF6Vv8gQ/0I+LxeKZGnzgWuqc3NM75IXRNW4nAZL3uDMMLpK6yCSSyk2
L2hXliXOcLJNCA4BRMo1c9aj/Bb8GjdRE9woZVafOKI6cfgd/wEQdwCBYqaBjlw1c8aG7Ggm+81c
otn4YuIycBthfNbwNXA+4lp7/mLxLWG6f4P9Cp89hRF1wTlluZBfZkoFVgHSUwaZ/a+jVKws48lS
htVRTPUNaQPp0SRdK3Lsbhc810OHPoBMbnPo6/EYOmbAv4+PPsHczsIcvia5JKfSrk8OZ2f+ptl3
JADsLu0/bOQz62b0sAhotn75o5PddqWBewGqsQ+QvKD0/KIco5Ma/JOXuXKCw9dH+7VAb4hoMWno
K3k/srxbeq6W1sn4UHtKDWDqQ9SlpJ8MfSL7P3EjaT2GyKPN4tKgulOAz0RWxBcRvQ+9vXi+51pj
5L9Notok6fIzZcP6ElFx+Ozdsn/xsxpmACVxuvTtU2B8tloQnTNzSSeqX0lChRtgSo7CHt7EZzO4
vz6nLuVdynvQtaQqQ8OYCDIF1gLGSL1H/yJmKrG+iCY1lbjXgd+ymujbmqRuf4fAApwSC+KluGru
Y2cQtqTGAkVDAiam1CG3yM/RHn+Lt19hl2LsNn9flxbRcwsqJji1L4cIxVa11sCn46Me1wgOt36P
qJx7ocuz5vQcwv005GI/KO2FlgqgSsVHKAptWCmhMgjmS6VUDT6AQ8dGNsTvHkd5QYpJWnvFN9fi
hu1t2mnr+7ZjNrRQRQ2fPX7liXaf5DbdAm0TOEmjXodFOQXMuuX+Em83PZLxxRpH98rgHLnGvGar
rsxiKao6XGks5g61X3ZeUil9hl4BrNjEC98VIJyR93C0xz8k7GVxrdTxVTiN7C7KXZvXvDZSHiUz
ZjCi51zLEfF+WJazXyWsO7qfBCOHe9MTA3iVakyXXHzUMMopzQocOJBQSA5g6Ue0hVn5wXvbWmKr
UGYkqWMup+apn4JHzzsH9SnKEnQyZI5veodXKJth5g8ePE2VeGGmUwKkFuwlLg4l7wY6Ak1keJWn
9xvfng0zCspty0yb+DR2n7wb9n50HxeKwN+vKETPifD2jUTfPND6XHZus2nG7n3Ld1zKtccIn/6m
jlQUkN0W/fmq6R+5Y/GJY5+mOBiS/IMuQZL7BIHac6a/AwrltL/Xa/tFYnfZ/UxRXyJA+9vwjvel
qOqSS2daTuww2+LniBas0ScNAQpHL7v2j3J5KN2L90bIZWg6AEnTZIjs1Y3lcP5PsOmqIcyHU5a1
LK+mbOdnrQCnD2a+NUDZ+FvDXLNAXbu7Ask/AVEUTGxwQFfDS35bnRQ1+3AOi+iAH0rqitVJq6KC
pa+eGvt8WEAqa/2w2FFHHf93pGzKPIefwE+gyhTpGuLZrH1Ufotx/oeph/q/m+6wr5hgIsL/JD4w
+H34GzF4SPTcXf4QVFhPGRTSYX4NE9BE/YmYEJi+zPWY3eWbxXr7wjPv9Py3Ol0ZQk/SaXYg2SLp
mXeRHyAJnwTmxCpozla+Bhmk4/tHmYk5RDO97c/g0DLK37+bXNN6EBNThKiAUfJ+xZmkpHYpvMv2
KFesgmPeLLNPDXWZF/uw5+9lStOjUODy7rURQ82UiYRZRAFJLhjLlXZ+e+hnUYqWskH9NTZhEm7j
evFeo1hi22zogZWKBn06wipm95MRbq7bqXZOfgZH5+8BV+EMvISP76pFwnalpHFc2WmTkzpfE8mW
r12cKTq3SbdJ10laSoEqqaZ4Wvy7qAubP8T8xbVEaMcGGTZe0Y6ZWAuWtPeDpkiAAO5JoYvWeBmj
sE9PO0hp36G2hA4pbHTsmzYOwVLXub6IsV/ziSNBnvHGrLQMUy4msXNW/1y5Y0Z88RZOg5/NebOO
05cjWsnjL/9rm8nrlt+rxV/xa4RdJnPX0QYs5kuIK3gBqZG4yAzNLwfNnnjJUY18sUoDyVy6HCjU
n9UvdPW86/yMpyOR72SdD1S6gtS75QKQitS7MZjHhocl4SX6Gvto3S3chmM0O0T+4kHsE36TcZfx
A9uzeWoryzk5YUo/f/IxXMmHEpGQzu05UpeV2kRzivenCZtqfrBM6U3LWP6/a/AficQ6ojkMYs6+
z5UNQ7cgW3N9+hBLb+PN91BShIzjGzYjc5DXU9bofmw7IE4vIQYAliPW4lkNQN+E3FYz9R+qVNQo
qwqpcrwhxXGdZ9LZzY7ErmImfoZB4JA/dxrrasjBqU9zu5KhCdljvflUiSK0QD5hyIKi9k1pch9C
GD/gjAXSQsL0m5tBLvyJA9/wP37a3gBne8m602yBhKMHznY156hq2VHNL26+dMU7ln3xX4TPrnk1
+wiuoMuWtqkRc4SomSq0ZqH4gyEqjX4jJOMXn6RoSVmJQ3j04nMCEqGsFlikadYzpIB2e1W0kGNG
+wwalohoSryoi5kjN57OSozPjZpq2PkKH/6VSVOk+h+PzAv6mUCYak4O30h9mjhKB1Y51QUyxyu8
lL7TAAnVHI5W92lVfKcKIu3yZUOAi8/xwqQLi42TQiKY+PB31UlwBNRttK26kTzGtQ7r1wIV0WEm
D5Mql+5Vtyik0KxzSKBHwrJV/cL2NKAesH+0Ck42KvG5tOIfENSHkWLaBT2Low61CxqW8s+94OZj
FX6Q9i85aThhd+YO4yfUTjTYQRlmSwJdiIUMpUkbYqbB5icsZ1E11vfSHoZiBEgJbfxvU7zfBOcM
TlRVo5+Sa7ITurTAKGt94gxuV95Cgd9X/4spWxeKWQ84W+vrgyQ5jJ7BN6kktOZ0jnbSykB0KYz2
SwX7FbyglpF1tQt0DDiaD8qfC5/mpVugd5jH0lkwvfgkXrPcIADqoKcNnZkt60d+fpg8UrdrpLB2
kxV8HvpQe9bi5BmHpIdfmG/7ho0yC2LJoSboSSecZ9iMJm9pq+Q99fghSdKpbj6r041xqYuiEOCB
KphCLfy0dOMG2Q4UB75Am0HFGu1ktafRumJ4ZmA6Aihc1iR1dg==
`pragma protect end_protected
