// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:31 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ndtEubPKjb09JinUA0oIKEPgUJFxEDOQAvx4hsuvRGJncyHPJSMg3+5ocGVHDHVC
XYWZON8OaN0kq/8QHQ/e5hlSqzRX+mnxmEfp5qmy959HBm1Kq9ZulJepHdxngmo5
mvNqrlHItEu52kb/w1Bqrv4WlY5774V5lQ6FR3qFlh4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19184)
OpuZNcgAH5C00wp9Az4b2ehRK+f/g6FQepV37QGolvM9qfhW29GHfSTw6svHZwX+
usOK8S0CVA/ldRhHFPKxzc2pF6Xqvx6PzbR8B0avxnY6Xdy9Hd+al8INq7z8P9Zz
54OJuEt5aGJbQmdrTPNnAl416oaTLs0pnsv6NyOAFkq3jF5nOdMFxOlsvPr1ESGm
5J+/6sDLbXo8SYiitTXLMFgf8w7NaewXCW1m21fUMRKv4N18ISWwV5ewIEUha3LC
7DvazPf7YoLPglMyth7grY+eZJgfOakveqKbp95mgQ4L/7HnYrzsdE1Y8SrygzSy
7twc+dwUjAca92hA09LKpAAnJQiezW0uEJ7wp9opRPGPgNFm3UfrvQiT/e/YoxmY
bbiJINhWi1zTVsues7XMr7VyIH4H4dwtvRBBO6IslN9bdu2BADCl+UscbrnhWBBQ
hwIiOtmwWZS+JptCZRI2vXhp2gnK+LqvJBQcRq3aL5vuplm3Q2WirwmZLDv8A+Q1
586HoYAqf7WW/RoyR/GS1nch53mrQ/XrcZRR/CfDFD6a3JnIbcOalmLgUvRGAQAf
TCiA44+/SyQbezuMl+IwyF8GBLDvZendxRfg//+xLPDWPXzPwc+T0dHjbGzxBLBl
8HNNXSPyDlkGSunAN+03UxNOdwthddS1Tfffz2hZNdnYVKdoym9eR6psBFi5GfW/
TpvTCmCxsH9981nN5zXZtDdA/Dd/KFmIJGsjqpLzStO1E0QaqHL2i++newl12tI1
HHzvgmoC3uZV3pgf3yVStYxsUNtS+Tw7XDvTRUwFz0U0ZnVrpVWNLGdQkqICcEhm
dM1MGlEbvaRBfO7CNKH+3r69N4TwhswxFFCgH7z4wv8Lx1GsspkOZzsgYXFBgXG6
sAuM4xLPQ9c6TGypxM8PKAF7Wd/ekquuXwaZXRGDh6O74S7JBpgIJk1CAur2H8Mi
0DrrMLbt98qZ10CAWqikTdUoMtzIljQsM46G7D0zYDcOB2guPTPC3nCGe+mUadOs
RT1cOeMP+hCl2DWLq/gDXFj8BHxGCvtS+QpEYoLFphZnMmO+aZIvjJ7zqjzBNI6F
Xo2F/j0LBoG6kHILbcefpBBHeJvDBWs4qdfm8+pxvV6G03hjlA0lUSZzjzyei7oF
0kRepXDRFzGbPlExmPvRWetMqEtoP+Ajqt0GF8LRzBkFvEgPlv+ujjZfACUogEA+
1H7UcRiNDyDh/cdyFercukAndmrQQ0Ot+82TsHwCoFoIgBhz568Z+Y6+0A7/5BtA
iu1a0j+IvGNHP0HH1rWfGLuc2h5O9Wd/RDdlCmO9cwfnYH4OVn9blDFC0xJIK0x5
ihrPuwDc1zodPbN4231RQvHgmAf8fvGn5u/oXJrMLcGz/8VoccKDr2x/gyW0dWbP
VsOLlQt8fSA2AP+9uRbnyRzjedT81YaVUUNYW+3vN8TIhGYToaaSGfpr2UporN5b
hkPgsVsjcW8qWCc8EJwL3nYK1ukZBzrqFwLfGXvqsr+NB/ls5QPvbcf4b8VT5i+0
bgYWiz9ipy6RoAHQ727I+aWmwcuKpyECEhYS7ejqfkbLz1WjtI+LkA1j4CMd09Sx
UIN2vlGPs+0ReI3J30KUG2d4WKv5gXZhu9wGUwHDQpRnmh1YbDfil2BTQ+IXEG9v
87EkLZ8gze1BfRbC32f07Sxm6bqPW8AocZKfTYp8ftpXxjv27MtcRRXE2unFrwvm
H/7Ktkl4voIhVYk9OJRs3mCu2BH8Vx271wmMSfuspkCHqZIVfY+7iOqjKY5aauJl
e104kPy/dCiQ72yb+xwJybTbrWzWNkOeeU8u85olbhO9DYVhn7x1NYpw5lYAN5/X
J0IvXoOgpOwJo1Iy8dJfFy5VASYX5zfe0bHagChCNYUGhqk9WtAzZlSWKyy/n2ol
5WjvV6tY+IqoksemmiHEKPMQAIthCoX/IqrmX8B3L3/N0D0l2hDGxj0vSZ8vZBgf
cvo1TAlsrTPvisYanR5UwNaKgHyGY04I0w6bPP3YPSW8MRPH1GowVReOnHkISRLD
wrgS7CP52KfLDKr4/doPdEaMHWaIuBM1Ppl5NZuncR3Qr6blZQpkb0APmyj7aYwb
wcSNg7GXj4khHDPB3kMTDOix3TBfbmPnbM7wJb6CIjUNO+LnviCLKj1JKHp1IfX+
Q/+zNfr189Kjjx3VmMC4RjqZHgUGc2JHhfrMA6ciSHItC+kyYT4EgLUVXzEhsYmS
BY+9BcuaE1zdc3+DKDhaKDzLmpSd+yv5LDMPW4Q9xJ/9RY2YutwSDJeldsQhLLbU
NfnV736dsVeoLmdkQ0n+s3u+ltQ8qghXOi3u4Kzk2ueh8JfmPDDQ/q+VQE8uIbs8
sNh+xmFzFuHekXApSNylEf+I+EAnGdCd+tPsWtoj6kJsRdsCNrhJTP39Zos4G0ER
Fa4eASMk0MCDpteTZ5RpynZbfBR582NrHtV+lKvCTHO9V6PzId6bp760/Ot3bFZp
3nWkQ33MYXlIahT5Kb1+df9+pk4SZyxGYegjXDcMONaxC90OnFLENubiA1eWjZnV
79zD818DQoV9rYevlamM1Oq5qq5h9eUHWz887mCOcdKo9/p65kcdvAi6iZPayGea
DJ/aTo6FK0w2i7N/XBawZjJGRLKk9JBKTYBsqrlas31l/7qkJU6SVvKF+VZeTwpC
5u++vtwYIFI2LTTC9Pf1Q9CXxjYHF9V5v/2jGbr4kG/DwT/tWtvRn6CnyvHmlAGQ
8FNqiK6FPTFsqTh4SmBzaDdwEihQDB9J6jtynzPrOPtuUY10+GcL+fsYTW2zTBsv
8IDD55V6XOcLAthMoa9uWRkZSYSGjqBu3hj7Ff6SQIzl4giZ9M+anYAsGqefQsyh
fwof6zqss1/QZGhHOinXStUu0bnAXS5cM9MP487Ud0779BBshacQuHFVvdVdKnaY
YDcC73lUaDeEkCrN6dudUkJpTIH3sy+1HgtkKIH6FHOsUFvGsZ4Bv8SL9XRDrxVJ
EILrRY27yu6KpdUBwoL2uUxb8nQFFJ2aV8ML9ejgQv7DZN0M0iEuaS693mhOw5Qa
S/zhElQ7eVWeqm3Fros8Q+50NrQGTPDcRcJpPeEzBiZPyyJN7XBnkFc5zFoN0W1I
NTb5NyXxZIve6UOkVrphsWj2/Rq5gwoC+uSqeRx57Z8zcLnSX0DqG90t7Fbcu6ZT
2F/joKTskKaGGyJSaHwrvFO25B7guR3uzloroe7eOBtqOYLJFscomB//CPsOl3xi
Nx6HZV0vEPfuqP92Xj3FLfBo6gWijjnTs7/sT1PDVLMVan3sl5YV9SsYAcWsKsz2
GG4RKRPgy+yzGhkvBwOQSCHP9KV4NSoSnq1+OUPIX2EDJoT5LKbyOEX/eT6oT+tz
hqdkHs7TwUqBwu3BLHjOAu8ellYRe+G57lrvABbb2iVI2OMgY5PfASPLsETgdCTy
R1Npi3mM5k2t0sE8yzKdK3P7y2lqvJBJFPa95JKeVTl4if8SByj5DNcIT0HhOeOy
5q0kZ8QT25dq3G+TobazCH7tzkegaa68A36hWiEqI9VFD5OCIu2TK/kwU5AL1LQC
fM7FkUDGQB+o1t7KCI0pfW2f9ND6tiopO7O2EAgtbFwNikGG/AMsYM23ejVs+7Dq
ZSr6Y8qbfzzCdCTyRr1NkN+D9zoP020uTgct7AzLzxkwwqkUchVZdiAXNgz9gRyF
ctVl2/NTl0tFjqPmICHRqVZObR+2zdv1kPPq3YD8Ws/wuZOIihxvL6TFkymcRSqe
3agWwf1s+h93o2m5T7hvaC9gKCMcYImQBIqtJTNHWquc6KV8WGUVGRt9DUmb1aQ0
dxr54h9xl5rDRWk5NAZVPWCKU7Tc/ThUxlAxMKj+4WXQY7KJ9PPTIPeMzznACU+R
VmTacOqR33TClC962r4yrw2U/7umeTC9BPe90VeFhL8OFdbUxDUsbbYimU0dmMh5
z3OUrpoVnRK/tgBsGeMM1gz/4QnFkJJ4bfLLDUdl0xYaQsQYvU4O4n3x/FhnkHjO
B7O+uLBOxPJwcdUMWVmw8mqd7COvB2aK9QLz7a6ieBs2ruDNo+eCV5wtqpPOTKag
CUiNJ5zQonRP82YQeeliAJIh4cxHA5c9NQOLhxVf8SYdOPlbdchyBz7ymTT4E7PW
blfFuVLJzJ6ffxdpS78oWKruL4agfZpyfhLKjj3spti37VwCU+4HLGz+D6vtGfdu
wFaYybX+/Yom1tJOJIXmlapkGyMmOC1lZXhioPjrcEqqo7x03I1ZU5i4XJlJOsHb
ZSiIpeO4c9d9o2tXowwGryG0VLzABGbkL8Dx6108qTjt6aqS7RRLRy6ZDiNPV1xE
Gk8BVjqF3RXRRalHxdcrurtDA7iN7IefrffXZzUbtXS4bj4zkV7nxXbZLAGv+xGB
tNRTvpBFrOVmAr4Ze2HVOkixN+Vc9pfbeVgYH0jlipP/i+uX+jYCEUMH/qlLMkKD
jFOgLwQISj2gzussGVC4/kX9hJwJicbaVdtxiAyluRAsyTEYjbI2RO2SzScg0Pob
Dn7oD+XpVKBvCOffWRs/ud3MFmtIHoayRV74lpJkSd5tm71wmYyNdE7UPIalbFm5
Ya7b75e4k7RJ6rwdqEOSgFy3D602/zY5+EIc8lIbk9BdXQknL+U8hPhP/GdDi8hG
DDWkq5OLi/bKrwWXojN0Y4by8NuRJh9kROktI3T5Mf4LlUWViA7BT91G6xXld7ih
XY3R5fuzf4DKK5VDFXEXwvhSG9F6BcSQGKSjMrZYLFDnd3iqje7qS/bu7FJMFxFY
HPYCAffodyNcPszY4l6ra9ntEXNkzfCVJxu2WfCQ+z0FCXN85wgLJCd+udcd5DWC
H8zeDh7EdGcT3bNSUMeDXW+kW2u8qizCFm+zKbOeWBl3vsNv95yZPFNfZBjPnJuM
cxMwp6LlpLD+eKEnMGBt8d/ZDulNXY56UOFcg63GXHKEDUgJMBnAMp2k77lNdDOo
z1GXerUYuqkz0jecjcJM0ZzDQJ7O2aEo4xSvhZcqZ1EiiTc6zx02fQmvxbfrUktJ
Az46o4HHJEC+tRk7kqucBQ66eyKcumZYOMKR+Rl6wvJbTgvdkwzvXcHWWJxkey5o
kN8x3xyr3oHmiFkwqAwCFH4MxlaJJ4px2D08jlBzIJU0EVdAJM1jSCESkTCyZ4SY
C4ffzviAR/i5tW6Yf8A5U6PA0eUEp3cNQkkst7a2OVze9YZz/yl7Wykc25g2TMlO
aJQZ1uZVueRTNLStC+f8DZq9+Wh5GslPdyj5I+zTStQjFyUbY7fCQobwgklp6RN0
VMGl3vWyJkuTBHNum6PgdDObvYCMq0GdFvnFLSuB0KwYDO2n0LPds083B5+B604R
So0lJrc2Idz1Opc2X3sHHTKtCVSxP52ZzhwgG6CNo4BnV5EDQL+4Q5slYLVqapYg
zVmNjYMgmh7b2pBTJi+PsIcTEz3ATZK0PMInDo5mB1FlXnzA7ZD5pCXNOHZzuSHb
ONzTGyJvHHJVXCv6NL2P3+KFSZ4dh/ZMOyn4W1wQ8W4KGIyA2TMQVYUuy8FT7Yf9
Ponp7VLoBkUSn33gyeKP+mx2coK0Tonyv8abvPbLm6+mmPvTC7boS1zSNdY7gPHR
5qn7vy5PvBg64T0HzQjEu+Sa2+6Ir83h2WCDdd3/fmJhpv35rHF2kqySYh928SFy
YT0PrBq5E3ZCqs+kow6NuCFMjh4ZsDatUVhoiPl4nNlJRGlXU0ZrQsEJhMvL+vaA
wz/H+aNhbwRF7CVBalKq84zW7TdS+hg4t8p3rTDjmDrRV3f0FReKhJ68gcN/Ad0S
y6kvB+HhgSdH/1Z+dVgJ6tKjn+Tt24n9s41yf7TiKjQGQSRZCg1lJQ/9BiR9R9ak
DDe6eHS5aDi2XikfPD7L9bhXmPn4IXjqgp/t24zdX0zjRvND435u7zfKAN7MmfTS
Tq68GW+Z3NXZQ7iEfYkU0nSG8TtfLe7UPOAKIH4xulpJ9h83+YBMKtlSZu5a0KRM
/eoZZJZ4VTkq1yEH4ULfDHycLetYrrPSfdMHGPy9VRjQxPjZv3+UnpTChd9FSrh4
qLJlhj9ziecnZo2ziQOCtjeeKxnI724lB2kf3GPkWhRTM5ojFJZdhPK1Dd8qj2+g
A6M9EB1xZpNcPxkjrSY269mWyYxBI1DA4C6cs+GXXuBAkBZ8WT1kC8hI0ZwWwRgc
nyO1II7itnKX6T1YM/cefWLTcnyAHSv6DbHZHNy0ux0aXUFxf9NRLBlAgC70SI6B
QEjh1e2BG7j+2pyJq3uSQrfAdb8r7Aos2VOwezNb8C7h1JGgR6WCse9wCXhdZ/B6
dtJuTEoiAQlkFkPU43FuAr+i3h/CYo7zyiP8pLHkfDcH+JxZ/yuI4S/590qrNPyV
x9nmuQNjwjdFw1NmL8hLkZV1RFtVNnRy5so8VOWvb6EbgPHKlvpnkq+lobgXyAgU
s8cEiojius5WUY0jZ6tM8Y6H/rre2UWTHblKZGwudmpZXmXd5R9V4iKNzIJwCs/j
N4Wd/HjWzDtqzAyp+S9AIy/8cIyzgNyNjPIyin98jMzG5BOXRJfc+ITTe5Ba1aVf
Apbo5zEOZyh9sJTlWDGt18XLRAt/+jChmbTzJbtpaFfjE+72PrjqHi2vk6BzSJiN
bmwlPMzLF17rz22fC/sVn3SVd+l7wyQ294FhDb5TjgWHNwvAXUlX61y5wpKD4j9Q
GRSIEdz2SELc9dPbz5aUsYP3pLipqLQsuhV74jL9TfDzMpcbszY55vA63uXyAwVs
SMytCgfU6VimByW8obDL/dpSxx4I4vPQbg6jL5VsT1d2fLHDbnK6e119JK/cOjnf
DeNNo5uNszqFSs5yJaL0zjn6qJ1yS3QjzetWH/MFMb78V765in8ckg0HUmyWXNkN
sA0qDJa5falEkG3aIShqPniLJOVWrAScqQ5XGz34YStsRLNi9GBmMtyqsaVJCmxF
dbPbKKVLj0i9RyMJJjZZH5XRd5M8x+jDt0UZqVX4QF0708I0p2APOWomic8aLDbM
ZgWPTiFymx4SP5/VmeUyPaGolrbFUXSBH7RfIGQs1JAnoXecXh9rAOdhbFZVA0Fb
N4/9CYxZSU405Dw8JnDDmRYXiK304NcYMtT9d0Hdf5UskkASXBvcBzIQzhxxt8UX
TMXVHDYmZr4nYbmot8k/+PL5L/nhmjt2+Rvo72prrtJ2VRwA1TcMoSUndm4j2tLV
IqlbdahlKxVQokGVdIhKaZ6hhEZ8HcAVusMXuPOlNeFSgZX4BOVWmoMH/nzVFhTI
J2uFdiSf209klCVcVdPMvQaqgM2o+bvzDfbYBquXrxYSZa41mlQKNHaQY+7y08F8
LN7G4o5a8EYEBS6k3UAN5hPjxJKAXX9pE1D3EP3tyRP6kxduww5BmsJD8Dt5Lsde
8MESET0veb/oUWyqIx4A84c3l7P/4moghqv29MuxXEk6Uiu576IYwGiawkj0qxR3
WGiXbXdKJyMK3cYlGffglgqAQkR9ZQf3MqCWWej/bisIVEvXTd80HBt7+b8iFc53
JgGc6tCZknlNM2MYKvapMueDDA+SIWNmYVQvvGjcUD+5P7Rj2vAmNcWoZQ6rI2s1
8ugYOMmAQs/1WXxOlLCllF5rbinPWN1iWbELXovtZmv2+SoDeUoI5LfmW0TwNPfM
49fPA/bKU6TrVtmXYZvkgVpP0jlYtGVcmE40tVFPSXTm/A3lVJW/ttTuhE8SeQ9F
ZS9jmCKWbv7lsQm4p7UC7tlXQpm9HezNli/l85j0l5w+VMo4uDSWXU7QZOufiXgY
EGMwctVUhGAOEz1ATbWSBoNTPNypRfgZ0eceOH3tvq3XFybn4yGcknp7Btb5b3ip
7b2qsBKpGLU/P2XoqCS3hUkYHegrxGLrpjue5vRtgzDsv/zEMlzRFr/NhugkYGvb
D4+JMvvLbCRfpU+UyCsHLVNi0V+nJfPKIW8vKbU61zg8Q3uF7zr+PeXzb34FNCC+
J/ZMY4GTeAEI/+qITxk+zAc+wJRtJokH+KROSStIJyQQhbEKLRsCY8ckaxKxpjwH
eKYtDaX/tKfdtHF+H+Xi1sBZohCjBv6rZ+qUvMTeu5C8/L47/zfwO8qH7RCui+3G
Uk1Luadm4GiTnCgb7hD06BqWaM1UwZr0vMDdgML3zu0rbq/+GhsUMS5bW7GNvUv/
7blK/gIG2D58sCWeYkxOABsWUfjhdt5HgvPbIqpwdFivbtdVB5+Rs7ll3olYFh8u
7Fa8aJljP7NIcRFlTcB2sNiOoOW9KadJ3tL9bsbr8adrgSLONMcnK2nvHUQM12e2
o9ahWNGFlPHeoojcHniAdedGfbeM1yqfLInPzZi40FJb3tYg9YSopBDURcuo0YuE
t+aBe/G0Ck+BcgOetU5qfo8B2iHL0Exdrc0p9+OLAboTBxt/Wn50+tQFP0gV84md
Umq/3ia7u39MwBIemdTi+qgIRlqtCfng85z2DcIF3zraGDWFIVFRS42crROSBwif
RfDbX5kRGSHp7891UlcH3+SHp21B0dyLlJEs0/2hxhYLTEyloaAr+nalFrqnWlxy
AmIqoplyT8ElTIMaBjNdMSOAKoXFZEOQe7ioeZADnq8MLXdPrybE6x4IxWWFJa0c
fTuSjDBcexGzE2YdTVzOfbaJGRTaU4oqesqzPOJSBjJ6GhIx29q0zfo9EHNsuZRU
w83XpzO8LX8wnPsiv0eYcy28xJVBZb0ZuxV/JwygF3ap/pFXeUUGgNp/yONeZPub
RuqsJ3ZRsMN5/s+qRtOahfQHWGsgo/z9AIwBBMtRwRQEMZ4fLN5In7sii0cpKrpR
5hOqUAgLt2atM/dWpldmhb38q3G4aNlhmewqfaokoVUl9XKruSzXCupgTrJFHote
M9oBId2xl3UFpOiwH4DEKRfdAphai43f4xSVCoHkH4TYZ6qVkG45Ca5Ge1CCIIUu
Xhykz3QK+4fNv0gMYLsMCVY10oD9gjXNFyjlrTRok/E499ckZWo4I9wuG97TBg0g
Z5zSCMcYF/ZIZDXtf0DUaLWyvRyuJ45lvyk35IB/QtJWTXLfEyAUCEdK0SK2nj8t
rOemytIuKyC7g8hgtwx1Rdhz3//k1TY/eWO10TkhK86Pj0eq6errOLOuDd/qaXbr
cwGFHIxFqnKgIO1PLF3pGRZyPOi06hF4pCrX0kfW6PW2uOMpIerveeRRwi+QTEHi
I9SXE5IYuMwBs9on5CdJRW1r3gFP6ZohLxIaTVXFCTtBd9RsdlMH+Sq+bIGGyBxy
hUPdqRASnPM+zRDThEiskxk86gb0bcHjfoFqO0VZq1y9lx7882MpKdivWelkxFZi
EzjHBU3pcSrYE2IbhjNotT4fGoedj2uBG3IH2Y9S/L2mQlQZGeUXXXPRM5uqzRh2
V1teXZCMyy+/3fUWOOoIHChgOKfSmp6lBSD5larjgpvAbGGKZRGcwywQPxrcq6Sw
dnOGlEcfbQGVqDV4i6yicIiPAwWKX9W4gfndZJlBGnC+329EHPI/6kn9j73CVr31
iZsvjrDYvYF+DtrZIhU+laW5u/fh7t1lebfxaUEcTdSgqKdizVAXfR+FirUKEUCj
m1bDp8E/7wxH9LwXPIrPvdfxzTy9p9fDOYhawBrSDqUvrDcTuxNYB+ZRZIoOFec5
8Ufxmn/X2pspYPG81zmUv8vH9T7E1vk60N1o6A9R3RX8ZoVXnczjQe7oqd9oeqtM
07sISYytTSD6WU/9IakI88gaixu06FmzyC5khXbgFzpJOB8c2lb0InMKQSfwkn69
cekpOJ3CjKoPX97YdUldw0Y/dG0ljiuI3IDb5CKtZfHzoWBRUqfIt45zs4bvW4sc
yNIyZ9D7i2pTEPg7wWb0dCHfEguJOS0z8G3BL2UGOY6Kxu7Ft4hx9g+/tkJ9dxYb
JPPRXDnc3DyvbLJDajpfVeZGFZhg4I1ToMgmwMIXcoFBX5ufu3UJzA+PMNKr4raC
xmyPqGniPuY5kbBjhD+xNyh5jrUeaxrwwu7+QgiGrxwCDBlqTZ/lPMiX4w8QeuTe
FAqym/4anmcpx9vKgY7I/SdXAVdauCafQwGVD7zVMofmVV6f2GQ9QWZR95h6iA0S
ToKyqB6luJaKLyhMNJODCtIXttf0iqAZEIvx5lpWh//oq9CJyM7lbvLDd8sSXKg2
B/m3O6K3KMEmsC2uZ9k8jmVjIKmtb5M43yarJ5aBxjnHdgXP16PNC9z7i9qMsEEp
ArW4JW+UmP6/hV3VuFDquc/A8ZVYRNt6wqINoWCXo62QGCVjeuKCTNkpHuac8Q67
XxmdGhPmctr2EyGAenvoXbZWRrjHp48qpsmDgUgrOdaW3lxQ1FbWtEFEM3DuYK/a
qGvD90Mt+dah295t71csCVPTIoDLj1TvJeoKD2nymWczERz69ARNqCW3buI8nHe3
hKVNMJACQoXvPStnB2rr+J2NS+F/9kOQKQR/Gh48TEUP+nACk1Ia3tHMCDf5IkR7
VpZC4gQkjrpXXbj0kWd4Bi2UqQ/jKvwJtXQCvGACV57lKRhtUNL7eE6rPloPTWcV
ehrTrQOQ8SQa1C4G09elNbt69AtpcOyYt6npQDwaOo8DEnVAzhBPW7BuRqHQemXy
BDpkQuZWvke+8dzBXV2iadZHcITngPjDMAdA3pft42DUPGNyDeSSVVfbFVP0TvKC
0Oz8lvFMOCamQFx4jS+m8H1BrPZBiUrmX7F86GFNJji8K70y+OUN4jhhAGhis922
OzAt8Hi2Som1CSKUdtZz/Xg1LoFQl2mj31DcdxYI1tml0PwBAualDQ9WCIrU3VdS
jJT+pCogUoZXUoc0+5u4BFEPk/P8HNRBAP9bd66C1FSlJHrkl7/p3ZFtGkEYwlwK
LVCtlx7HvE2H7UF8JxOHDG4qL9pg/yCR9Z4PGXZKjcTPNFlcbO/JDDE36IT+L2fN
Es8Bvs2QhvdbpG3u0UCJDPo42qdZmeitOZt/yyrJQlTpsblsklRCfQIn2HWlpVAv
/uLF7osL8qafECSshPeWjzHxMzyhPLWCxVSieKty2cwwhwwShoVGz+MndDyK0703
cs2R1ZMO+xD5U2guCpDx9vg86aYbDQiVmc6q3hFa6T9TvN5wVuN16jGApfl8BEN0
cR2TKLyLT7yJr4tBIMnXmFnDs/mkuK0gJtYhOauvHhyWpwCwmnMWTo9ZCtgHITcY
yucAimT9umfu5sn7RhuNhJcMSc/KBvhvVUrXkOWyjHLVRGTzPIOyHkSSvPo9VfXc
F0FfDDpXIB+zUcPs+8ZcPCixhERHnfeM4QUUhAKVAM8VQPV6LiPjSIbx/6q5XAYP
JUVTm8yOU5RDBMwc8os9/rbXyuvq5RwSnvfNQwcvIBXkNWMt0h6IsrhL2WWOA/t8
zhe3sGXEN2qSsDlwgQ88OmiFyZ++uVvOylo7nIB6K0ObHOWAR5+dHSst9I3X+0UX
YImAqhHS/t8W8w8AO7aOAuOsqEPyIO2erLCxYukcnqc8kRlTotkJAU1W1rTA2oRR
NiJ3994ZW9s9e12JyAHWh9MKsc0bR4tdXECbXyZ0HJoE0RbCO3RsRcba8c9o9JIa
zrYdIfeMf0oLFFCkdYGWcyVyXTSggQJYprzZ3NDpH5kmBkudfVZYJ0p90mFi7Moy
EUFmaUgQWoHgIAnVkMd7lNXSPkNDWabLIIpCqDhDTXznTPxGoR0iE4yeIlaHuHUU
KvzkGe5Wk6wPcfE8UQpIliJHgU3CPtnQoAbHY66YaB1uTCZoLqZ8LJ9zvNKUKcw2
1Z1iJ7wqzMwcDhGoWmiAKtt4l1ubFGzDu0BRS9uKV43UxfUFO9uWVJVDogmxluc+
75Xr4l5+agq8HeEVxmoSoZG2D7XHueC1gDym1BoOHydk7aZbHUYy3egTLU8gZtQK
Bo9Pr2hzgZ1AYios3Xc3UppXSTam4koGrkMchlNajK/d2GlGHaJQasS9uJwLL2OH
VcnKr0pJZ3xaRTfmqxjQhkSCwEh2Q3LzsS/9BGHk2UxWAgmHboCGdhd2ui5evcWt
Efpqb2Fxxb/bIh88EADcJKjFPjW7PXV/0GvfoeV3nubia6VltTh94OKmSFTnlRwi
O3JG0jfKZyODjPLtJyoNSiJ/wkQq3FHQu+CLQT1UTNZgdfUPZj5x6V73KcjgijZb
vOoijSKD+S0IR+cG9Mr1LA4CAas10GKvwGUUWm0fe4XwQZGrvjkNfsl5Z8kI8YCl
qy4B8qJa9N4SG0t1l/JZdticeT2CQgHJd7Nr/+lAexCxkylEPuOuo+2wIVJ1pOIN
aITjHRkv0nnk9Kfz428Ipzjc7NBpbY5Hj+mPgVbUH7QG8E+D+O7z70+rx2cRvTBZ
wz0/yj4Hv8cP4MqM83Xf6A0kZZy9iEcvBq7VjyP8JurOmnhqhv5qNR4g2Nqhr4jx
1zJ0ztVx97JYhjNFfTWthhyGiw/S+VsV7ClxrWQKSMd5qMpsDVABQRQbDRURy8tq
ViDOhTAnJBvLPiFQaG1uTxsUmRZrcDwz/GQZir3nQEiNgdrmTr6pG8CrL9Q774MK
sJ74QkOkQ96xq7lCuPsswRXMSKrlxBN4CDxpdFXctykdq8pbjNFI6SgTyTT58ViY
dC7eE55TLNUpF4tcjEXI0461B56q/db1PIA5G5xxobbugGnUfB35Jd6PQwdjIKBW
EO4Jvpw9MWmtBKH+qwM7XRl3Hefl7kPavlF300BhAeVBw1SmqixerfKpBWQUsPSb
3rxDhJn7tg0SAFh7wFqZaIbRuIzZ8y2yURE9vnfTbyfYyd/Epi0JlNZrxwkCym7U
L5j5UDiD+jG84rgN/hxzKiyWtZ+Qv5nVGB31OLLk5gouBokQrbzAQqEXlsd0bEec
I6MWa0DMPalmH6iXMasbD5wEBSTBVx473DYPi090gEtYXIV34P9/sQ6opBFyeiFZ
Kol1RAN92Bash0mjtkIDtHSKPn1TE7sXXQ0dEg6jE93HCQTvrJY/h0sPO59rPXys
/7gf1jJM8ocTfN/GgQI78vKgNx+e6hMd/ez6oE3fxqzwliHTex5zb5dtXjiEKkW5
dJgqeFe7+I1alz1HtTx7CvQYlrcVhH67yj4+gEb0gFX60pP0smSdAslB5N5MQFyl
Nzt2La+50utBQ9ZhO2cjVJUONzL2Jz/9P6LNAERGqQNliC3aUK5TDuHnjt++6Z6i
Mw4hzjpzDFMJu5ef9R1Go7xl0kDKX3e8OklXaM0v/nZ9o+l8Qdmu41yznGVIvdki
PahppN/hrzPtDZUOkeuibE6sshB6Bz5zn8ufGFr1QiXl0/VcFIK0ORiEftGVVGd6
RkoS11M6S99TduAfscXUpNz9INeeg1ofJJSyf9/oTkAbw+/OfPege3seE1aTiCCo
GHiinzTSTfBNSgg/PnRWbprNAKkaEc6fK8nrKHfYjMXOsCRnxVtogrxkUWdULeDr
PYjXqY25ORnMu7hZiOn8EoK3UXocIC9nvbFUtlJ+xanetBmAo8NwKiDsJubgsihQ
VdPHQMJ3+2647Auu/7u5l241Bc7edWvoTDAcAYdQAJyq4sUb2n/MID1N2rqK7z9L
1CpfdnQGnKVbaoOgU5G0Nt94Uljg35XmQaTgm7Hhsq2Tem/4/znp8f6KXSdmOfUJ
vhU91OEX062YohTAUFiJIL6Iz5hRfp1qfgEnkppFHYfgcTvwun3Qq7SiheZ16Vgo
eSNFuwJEwg8jzsEig2cg/rCt1YF1WzoenvxLGtiG19wGnM4CJS66IkqSYyg9po0C
T58w396vP73TpoWvNsKJK/NENG5I78PYqYlGntNrBbrjzKGVRrT5Cx3JUCV9HtoB
sKUDaL7Ul7n8eeym1j6jA2XnfXfcyy8ThckOJX3SdqzVyglEeBfa+7s3Tn2gGJkp
fqoQoV8ECZV7yvlYhqRT3Q2V5whfiTAiHQUTkka/syvmsVlj0YPENQm1zG2CR/08
D5ycSL4Z/q6PXUSKbWCTpYh5HzScUCWPc9KZ8yNGvTgLkjFn1p95AEcgKZdozdex
Fgi/98DnINr3NpSQ5GoVgKYLwOutXieNDoBZZXyVyr/vAcuh9mff2Mp0HWzFUre7
wsz7Wrll1rAo2cpTB6igng5ensIRX/YCx2zqTVjrB8SfzrJBpoagVutR6WaFIElY
x1wBH0kwjt/pnRoq30JO4yWmHHpfMuT5z1pZYIeN3EwOWajSILXeQFGPepbYh68d
34q4FDgF83RSDD+TO0Wz2aa7NhtaeNJFVacAFJMaYwp90al+Wy7GbQCWW1WIJzU3
aOCLNAtG+ovDdOF+aLsttEL+09iuBRLPHN/xJESZCYVnkYeWJw3uTSL0U4kijsay
vV3zJNUxz1sD1fHN120e9VYTaQxUAwiQq9pDYlJjjDAq2FusWoLkSgUUu8QZpTi3
2EFZYDya3VJTC6qn1i4BG2HhoOLYcX/6sANR/vcmPckcIMcNQ1SGbwcxxRwKW4MC
2GimTK91eIUlvF3Zoa5LUePzU2bPjeukHtd7TVyKynahe+jbcHgem/Idb1c21BD6
/Apdp2vrKwS3vlzZk/jTjPChaz3bZZyYPaka9YNi6cm9lGaq25K82JwteDmRUPfG
b6NB7x55BYPjbWwv6wcdDpsJ5ro/tt/OJZz4VKPVdexUljMniIB5pnxg/Q10/5Ex
I3dwT6KoG/yHzvccIy4kflNnVJhIlrO3SMSNiQ+ZWrLwhZ5l59z9dqanESslH9dx
dh3nYil999jIn/0Vl2sv/wzCnEm/XY23rU9fQoft1QeFE5Wqb+uQlpj5514Rq1A6
C86ryK4YFbFTo/72dThIF07SSyidsEq+Sgb8HeQqlVkzZyUIT1Ly2kPTJgRcfzUl
iRJLQPhkRZITBa+RirNMj0ugd1O7XltnWj8Ttk64H/Oxi9j/syydSaeKdJibYQAY
+2xcytENtiYBUMgIJSwYhkC6A8B7E7XooSx+EaQ6jixWmVVmGe/28MSy4Ggd8QH1
RTFiqJZJRRxfJcpjiX4y9ER5fpIWrbm30joHsqIsGEw7QJGGe/3xCxxT8wASjzIm
Hq8I75PeuZYKJaSEbfOcpsfgvFRSXSYSY/J8OmfeOR02D63A4ggEn4XDgLX3Zt3l
ISixShqdD8Sfaiqc6cAMMKBwUiMlIBceTDM+HIFZ/8i93rbWcfFpzji0xalrhXTt
iDkC38kYUjHu8YttExonqIuLYXTkNKZOmWHwu7sp2adPmlSxZdAcMSBpXm+jGyfh
efQMi0RPVzCKumd7cYmhBePLnnT9fUs8aOFgz9Iieeid6kxRgOTUp7kZVK8xFGfi
udfJoRvHKIRNcuK6cvBh3qRe1scHwAQcm5COgL9HJT03xsxWuCzat+eVRJFDA2lZ
icogHaqQtY4uk0fdZzVMiwOEzAYP52KM5/g/fvKuCeZ3fk2H/vLByvjaH2WXnhlB
ZVQanlW4XXJE9m+2oyT5Nb4SAw2LyZvOEM7wIdKQDuJ9M0EU8d6oWGm0necCH6Li
0hx/0xm4SFPWi2s25I2Cs6EqEL+1autW9uq2Kd/yxYxcHwGVcHcibPCs2e4wVG3r
87/XcX37po8eX09BFLXGA+npMpHP0HZV9Or0bbvqpHGLIFnnx15mq6LZCxa4QPgu
A2adwQyLas1lXLxh/on+wy6wCENp3uEOV69ZLA6CpaCPPCRB4Uxf799KA03gxNe+
OH5YI7cKm8wT2q0QetlMxsSQ4HO59ue/NijLYEN5k6ciiylzGktfyj4QbGlKALxb
pd+hyUyA1xvfnC4462zLsS9Cff+GI7+sVcFYbjPD+03kdRqAtMXJmKyaAIBBAFwW
GcBwmocPd5nY3ud46MRV9TQqwzB6t3bMHIQHR2Vx9yDTZIQioDG4RauPKWMC+2eo
l44Fg+PHnxaQhZbrHg6/h+YoAIvKIyjQ7nDs0W7xqW4o8JH/zPjhlC7/Qyp2ZAKW
QHQ2ChrsYHrKiOlpqy6qj7FPdabzY60nU6ta59/qT78KNgNLRGNcO3UjckSrrpKW
+/JYRS9VYPwx1Kb18gKrg30LPeGPD8U1rwjwP1DIIAW3c8s/Ow+mj8V9QtYd9qJw
0GexoDMP19pKY31ltoiBOKXvslkiuJEBcuMcG3n70BvfoiR7YwNdkrmlYVrgLF9c
CQIahT+F8DpxDjRd9uj0kv6/ipuod+ml84+onAgt/V18qbON7l9l9JyP/tuOGoLg
bkftClx2ZuH9oTqUIDQvpzNHN5RXClphpwuC4LECAtYxyFL0aZnI8BhKyG1exOtU
wXp5b8N8pOz/HGgTGv+K7WIOTBVLtrV1I6lTX4Z3ModtK1PoLMHO9tXYtb51e+XR
Gat4EQwwHOsa0yU1wVIKnluXKg1HaIA8SpxevdoTJkS/iTrFOsRomcT0TWM2TAUR
evCUhaS0JQpFMnNFoRhd81Vir1kxg9GmU0iUgx773BCjjQzGXGlP2qizHRdkQmKn
g8jq99JiVbVyEKhLi+BiuJPXjR9Idld8X1wLWwL9UCFABAXwfs0eYlCBN7qHpofe
atvTeQj2hF670rPExopfDcUKY0oKlkGOjj9CYYWV5S0rHmpiexJ/p4huJmRFzgVY
W+XRFcedcD2CQfZl1bn8InAGDNgZQ+2rLm0od5D9w7UuoAKsvsg/NT6XzQ0XH+Nx
/dC2D2woM568VUnhR760ogxvAx6t5yjqlSZp1lOh9oDuA/BB5ZfdDKQuLZYlkNBY
4EyHT+TEWE9GSMeoYEoaXEKdj65npP6J2jCXEKSIfZ2pgRdG1Baii9vE9IEL2e6e
J13kf9fngdY9hfrlY2QGyMmzL3/xvl5SGRzeL1Il8tQvS9H6QnaEAzRvN8e7tg7q
BBB2KNkKtIpx4LrM6tQCGUI9T7dxGE3kjUMut4TychF5CGZk/4jso2SKw/8JsUQg
++EyZLG2RdZbcONc87YQmYcVBD1xnM1ECrgqU2Y+DxZw7oLTQ+1pAJZa7MCWDzla
T/Qf5TznXn/yNOj+7zh3vbApGXST9eNNNouk7cOyPznoVKIb0zkQXBlrj3imm7j/
HMd7rnDDXY5QaxB74DB3/y09JeR/omqwvPrTG17p4hzfW55IegdeVwSjSfNhFEEK
0t1CL8kiIbsUYYfGDBgU/U4etlsQ/AyDZFP2ujxLXRxqeVEY3tR2Yb8iA1POphX0
o2L+3i75XcsSg567o4QSqp0nHJTfBM7Cn3ElT5biLa2ELmHNAwazSsrEvMmXss8P
b0XePE/G9vQJ19gUlhaqtH3ikaBnMVxgtxivHaoyKaaIiwKFAiaCs7bhASrBG687
iyXyEAPulImsgsPShhhXzgZDuQ8iO1ApGGp/wz3VL0swuOX+6lc4YdtNDDC5QoAp
uHA8bk7kDiSVUYuzuVwG6uyHp/y/iGZBViQKy2mGbK6xxU0H63m7gqte3Kwp0glm
Dtc8yOGKurDi14Fk7vQ8oSIe4riNBnQmynAQtg2I5eCF3t1Eeio0zFYHg+OJo880
uy45jL51tMuARPwWWJ2EpyamL0qW3xc8G3+QhfDYKnAZu/vErHCDIAaSVPKlEQEf
efs+Ja3C5137fWkAB7xsSLFvvKJO1PHWWjvYJpMZsgvoYcFgzGfftnx/AW4PMmmO
O5cbRpmX24d5rwgjWqOAOqdU9mu3WpPSzUPIm+U4v5nRkzz3bK8uVpWACCLY4eKZ
HItX+NeEeM3c2UMYQ7/+igPN8jInbiI6Rm7oSLkRZ4R97mtWhGm2t7X4+Sm8bhnW
iiut+pTcjRSn+WkqU/ERBTL4j1zE7C/Dz3WIlyQGK684M9fNIGgMUlXQcLZTHwLG
5AaSbcOqstFVcZ08QrsA8Ai7eVt8HxBXOmBLKCQSmNpCHTuVmpjvTwn/6rjs8QlP
37Qf6JDm8JqFvRWDcmNTtWHdVYbZZ6D7Uaa6GNWiqArYLtGABZuTcYs6D/x/J4EG
J465yqjCNNQ4QVtHj3M3nI0rc+pDi19Ft6mL8auO3DViqo5ubgEPUwsjfyblCXJ1
tjCQ7d4fl/1JCNI+VnJiXvTM3n6IRGLQBPIfCfKqgMGLeaa+8+nRfuE0Vz73Mvid
E6wmEqc8RRUCxAzhFmnc4s/4BdkM1sSbj6Kx5Shbb85rx9wSnA2TatG6mFbaEDC3
SKcoKMG5JqLat3NgAJVdKcubvcOJbRxfqa1vkfxvFfk1Ppe1ueKTDeeT9FuzpkYh
1A3nyAa6Rn1/NnVniXHCAMJU2Cs85AYXjeFl0iirrp3XCfLDk4cT3qncpie888cz
J+WBTB2LT5EZduSoA69/zNronafHcZrsHwmbpfHQX5nrXMwhKzjmsqtHwWn2wigs
16F4P72aV3HHllABe4vkMHdLbnHM7AUOFfMK6nelFsK3dNR/slugHwrSzMMZEfKH
eA7Eh/wfRgZ9QvDtE58xPphPYfcHhBqVn008xuAZEKjzsbKSAE/OrXJvHt2AMXJ/
IoC14Eapm+wtPQmP5ey6XGBBrZ6UCvOwXWuzStsGbS5Vd8nn928fW2ff6hrkcOCf
egcATjdkEcWtXoxN1kUzc3vxZZfaEuoYEOFQV3b7gX6uEiYTI2DEsajFrT3w7wjQ
eZyRltAeXuBn4z9NVVneculI8QJNRoba6qjLL0sdUdynT8uIrxiOG9XyrE/J71/h
df2qygPkGk7gwKNfGHBSOBH8elFN17TrgXseY9DzFrPqfgOS+34eOqLi6KGnKQds
jSNR2TlH1c5nvddCNOp8AAdD9/1y7raROHQX2LsilKDdbB5p6A6Z2pvYhIN/zxkY
NoStsZuNJerNFnUP0Gfm60lXZIVoWqtul1gT/PKNhZiCt21kLMaXS+1GbPPXkttN
Cb0PL7SR25WnPIEQe4DS5SvVr2Vf1FXZpssXMLVrLvqAHYExMPbhLnpwLYNOkNCG
LjTChVUbG4IaDIaoLtxoUUtbYHMBaNE/BOoZ8IonQBbGfxUvjx3dCch7K68hRQ+u
lBJYNDalsiSDOJL62cCsvhrauNlO24wDKUSHlMi0tFNFc00VJv6Xa4rJhrMW7JKO
a+uZwgqKxO1STsi5NLQWra3vKoGPUnBbDjn9hNUTRKxnRGNxdPl37nBJNKeJ8/AW
fsbuMR0Dr2F8Os+tAIWoi1nUrGcERy7DuqG2UjBL5bTjpPlvZMJzvnwTu30zzGHF
+bxvDNs8UOxk9XCEEAmmjwHAxFA6IPfUPCLak+D2Z0YYoOfcIxVkSY+HWoQERwso
RjWGCgmW0q7jK1EURndoTdES97NZZa6maBo9Hen5q/j0XSdU7J+F8EE9rhFQg+aU
1RrhKFSG9pZgJffUAnnDOZHlOzWobZ8vihnGIjIu+ZphaOoa0Y7wueY4xVV6xJHK
2KUTNm43DrHXcJj2T2+1cGJZuoqaBAEtqLMReLVrKJbY2GX0iPrL4iRZMluJvGKr
rr6pfCqJGBLV2rnd6qoFpsS5wV6hdkS0+Hf5uBNuEEqtjfG9TD+KB0P12eJyEgsx
+m7ry4R9+JB5HJNpImX/vqb3DZ+ub9STXM3Jeoja7sBaCTXuAk7CgWhXLXdAR3/8
y2t/fBIf05AZHwSTeuQFcCFNuSJJON9IithH+GsidVzJ3WRk8MFf81pSQ47ZNRO/
Nsbf5n1dozboiUpYcXl8uO6pHMa+Gk+HSWODdJI/+KifQcXL/vmFUfMXtV5Syj9Y
VHBhz+E6YT9rQj0F9KIE/Akp0qZIgcI2ZPcZ3ONm4UFs1UwrYnWGH9++U5azlcUP
oluDPVLNOu3plHNExWqZLdjj2ALBxDeo1B+TvQF7iKo6mJW79l4dkrsEGKDnw8De
s6n0LKdCL9EJcwGNOZJZYI7PMXM+i56HmQf2GrvxrObcEAWDIPetYufpD9MH7fC6
siMCLaedNzIqJvHg7NbrIvgmiGq53YFNc3zqqwxMIWFSq3gxrJtfouU+Afa4UyP0
pXLw18ymrPGkI3IZTYfJSkwB1fMZsGRhsudryQa7RMyIR9gi1VqTQBYbHm8ulL/w
8gfbkYd69J0/ynw4eqEpxYE3G1sPn9//zOcU87LW307wDfcDe4jMAI5CvfoInSQ6
49DBV9PkOJvnVx0As32m+zrJzgPb+Fo5DreklGnoZCqqkkL7JEkxGpOXK7svD0hS
Szqk3Es1DDuKdxYRmVs1gnKuO4ztvKRSXuWGCdsQHWPy1DUA5mE0we+5Jt/UvoIQ
Vf7ZdB/J/JCj389RYnb/G3RwN6h7Yo8v9Jxmw0MwckBdgkwKh2z5qBrUpr5gXpHq
YVwxjBlHtPFF6nTgRs4UjHzGdI0Ai1mEA3uBtGJn6HHsrWiuGpQhUCndmnHwb7+R
1q47PgU/fhCFLNBo4mdgdPYlG5WvYqKxDSEZZXLe/FZdNc64mGZitEJ8NnDntYcg
nHxwW6uaBmVWHPkbQ7CVHMdQM5Y9OW6CSr6tWQif8RBDdwjXrRK2qFkykeK1JTVn
YckQeAokVdw02CJvPYfe/8nVGeyCi9HNHayHEdmBARs3ozeRg06xSyr/ZBBxL0HG
DXOIq3VGcsWv7bPizt10pIs1szoRNNnHmoTTFR2HtIs12AXDwwCiTFDy2MvvabmQ
/Smlip/DYwY2hHfztdVowRr6ieQfAPz++c1wpxSnapRNurWrpUmV0gT90tdJPRdF
tMJRuxWGWQNgUwUydM+oN25F/kQpteMbQ28jcm2YSZNtE74QVI6pNbatsJb6JGQY
pXlRR2yqwL7nq0KSOAymGBJnMmXDS8vlr7tFjVt59FcsSB/5mf1wFkmQH6ucXJ7n
cv4cDsLUYbpoDBSjLpFli9WVgG7/nt/bRIcIPYL8iLHQN6v18c8h78NSFumejpO+
Cfy/TOsfLk8PX3yCU2Z3WHfex46osz+bYVp1cUWnBbsRn5FA6avpHIcTRSnarEAc
HV6HHsxmzRXJ7f0F8V6PQKfwD15jY9it13ZW4EyYagyGITihRbZbqm2UtxF/abzJ
JnraB7rTHWIBiI4Y4tmRZab1N7JwB2NMcZ87d6vKgrZpe7JUaKmwA8DZR/1rcJ7f
U57dyQVMGlnA7ltKXD2z+fU5LEKWD9OBIsbgSwWAQqckxy9hhq4XQP5Y52VeGiZc
t4nrey9i5D0D7WjRQMZREznYP6RiHYdsU8lpdmfrsmNxNCWlDhYbEQkJnf56Z9fk
9ED9USZnLo9Gs2t1V/yyT8AHI2qPj904XK/Zzmi9vfRq6ubTnqDv1R3b3H99gW9u
Tc8tG8nKuAMeMPmoY4wGyEC7wnfiFk5PmFNqO4crcqhsOBLgaGpR2sr5Caogt2sW
Os3I8rMlpeOe7p7KUYcWqu6EaCox5fUTNv5gSAFzq2BZf9YTLFSr5Q/qZDp8d17+
oPP+O8hcHiBflZ2Au7O1x52hSNAMD13iFuDfxrW1gU1WBuQYv+6WEk/7zdMY2LPN
dIy8R6Zjb1ZDOlrczgk3aXrfPsioqeW6xc74KQqNH/WesW4eMprOml22U7B06Ki4
06uz3e2TPIR+E6H1EsooSwl/RHZCB4+VqGGXoewlapK5yHGz9eAuspHmFrmL2xMJ
iKoGJ3yfuoMlWH1bUFqQ84794M0t0f3gak3GQBSjOkAjBGro214BuoDyzt4NSuwf
K93Ism/l0NG6shULF/GNriMsI8F1MpNClH+0kYJyFxWh+81rooEwwnpbTvJNzNiW
Y2gWJKLqYmYztPqHSCXk7Kxp5iWGAkCDg0MVjAKRO2c6x7TrcwszFhGsQ18Fcs+B
cq2FmaQxROPPoaxRx0Oz6cEwLrM1kA2dsyQsIqZ5/ty4gLLk4wCF1fTdo87A5i+l
4dVikqy6rzTfVrMWLa7afWppA3338jXJlVQb39mXliis72NnbYZo4PXZepbDVuLd
fDQP/Z6AX0+Dnpy/D1d+BPk1RQ0gBQ7E23nBWPR7iavYdtuLGgyEj113JPpxYf4C
FVuGVTfVRoNIOzwcyT2iagIMJg/rlzZhQHfz0WP1mzhRlVdyUF2YmFyBViaKuqcf
/wsDiBmQ2fXbziU8MJRe5B8NyqsGrf3eP853XX2YqkveYsb46Qg6aBuoX7WOD2J1
d6e56uIuXdJjrl/MmjDynOlMwTEDVi/xNNzMjgMp+NNkKhkwc5g8feL7+TzvF+CO
FOyeFehlPv6BdUoCXoa7aSt//oTFoasJQz8VFjfjHLrwx9AvbM+gbJkVDkwrlEN6
Fn6aHp+B6I903gbPgEqtXsUs0GLM7T/Yjymi4NDB3SWtdKEgLXij6Wy2LhHFpoOt
yaHIy4ni2bSp3LeFjpP859/vLO0MkNwfuOeigXqrtqRRS8xGaO2yBAMnBMo3L+Rc
8Gr3nwLZTXt5GmYwBHA2bXOj0oKbGtbfG+fRet+6WyYOt43LJAocI9w+bjCKi0cP
sOmMEubx7Wjlk5yUmX4HS2zn/0b63+MrNi6mBaPebF4Nb+beQLh56mwAoD/N3LJD
N9Xvqjx+IJYuum1Fo0KCy6SFX8Kb/DwfBL2v7nBdM9OCPfmvB014u1Si82enz3Pn
5PkDRwQ97hh82cFP00Er7H1c2S4iPJyXtkkcPxGU9R6LY4ITSXUIGh1UF8dIQ+sm
Yx+WMxyqpIuZJdLjugRsZITj/koK+ud027Fg1PVSwFJ5aF3wYi6o6/ulC9wx+Pzg
Dov2a9bhaN+TxXoJuPAcYgWTPMAqOryx3XDSsuFkabRo37H5WPrHMRdJFliiHb/e
SM1jYm0krhqAFoksQDGQeSUPCij1WiIayHwPkkwA5vB4AOy2vUwe7MVHjxMo1Iij
PTMW6HYH1M9sbzB0f+I6sq13uCcppex4oH7jDp5PoXiOPIIciMChv+yC8Bc81g8u
9aRbyy/vIgN0jvsLVxMOz0nTsCUy7OkKp+VfznL5N7oDevbjeClinfOORTw8ofMF
meXsn8SPly6xMn4WEqbiM7QCLIUXjtLx1jqnrLLzWdQSwQivx0vwFASNL5Cl6CRY
JlEkIdkOfmr1nQy1yZpeNoWuFosrEUVVUaJq/rm5N/rH+6eX/EK67rzeEzD6APLP
HlZ4KdyAe7032bXpTQ3C0oFM5MygzCT2+tggzXDEqrwN9iv4R4u2Q/eZGR/CNqNZ
pOJ3HwHNAKPOO6Be1welLpZIaxpkSFzXhw6QSR6wMyb4wEotUs+E4Y7B6yAhDtHz
ecjpBaWB941+xabmrs2j9wDLy57pUWbkRnK7B1nc+rhu6dzku9jJyEBqAj9h8Lw2
+Gv4+7RPflyF5lBctGiYy3i3W4j4uQa8zDvdoxPLV+xOYsxDo9eUuklezWMo6i/g
i6vBoAQMagYt7WIii9xlktVV4CeX62v1ulg8weqb2jM48krEMNAjYxK06N5f+fcE
MCOm7zh+X0XgzQbzaKWkQV28n4MuA0U6VpnXH8Ku5k9Mja2ZoW10pY3vIxXDOrPk
7v0BUesN7bpHCBFI3G8yPsG4ic0K9HLOlNsrK7JLuHH7zu98TeR7UrMYrx31VCNS
hw8ABe3ASR0fAovizBSHkp/VyAZ+e2kLG4+IZ1DwVBCyDs3aBeqkEwACkXq7Vt+o
botboVYt1x1PzJ1uJeIhxrtCrsUUpJRCSLlkH1g3s6gZ3T0z/CAGNSY3rTQ8cCT3
1HYc+0YxI692NQud94UZp60xZCmcjKx6kTIHeve9Bf9Z63Hkq6slmev/HKEbTJ86
eriviD6HYxvByreSdn6GdiWRqRr9kIasB9ZpX3Vm6XNSyNBrJZDpAeOfgeRvU/ld
fRamgHXUyobxhGXp9S1cJoic48FELdVwLZzdE49Lo6gJiuw/x1KA8nLyFLYuXHb+
auYhcmzWMDfmA7Ne9ReeK06qd1WXVgvqDcwdApTmpPTd85sBSWKBzSH3zc5VS3K8
W1iCYQKfi+sVclLEx2lpE6433U4LWUTc23pZUSqcAxPQ+K4DFEoZXIzEqiRycyC9
DQRNWK8QkQUwPi/RSbRuAPMBizftuXkK63ofBf9htLl9q7eWrO6BygfcipvEWFGM
XGCgDVLf0ae1EiaefibMvurN2nBtDS6tojtv9cab1NCZSQbkcapJugEGNy3kVpNN
/rg7OOY0VrQaOFJiLOEiQyNhIPRGRfOb27RdLaOcrpLhBtBaAlR07IjOCDDv1PP9
0NN/YScSTJJLUauGUwgQZZ5HEnAcsuHFK8DjwsZ0gGRyf2c75eAnL6cP+HP/TNHl
Id1lHa6VzBienXOYfD0IXXZxtf90pu/iXC6NrwZbdeNolcPYmFFYPwgwM6dD547E
k811Q1QPP+od73srV6J1knTdcedWXIBwcwb/2ygHIJkts7nkIzUyXzXDRLuNH7KJ
fxE/1O/8JgafKQmmAj+r9l+Jl0sZ4wTFK+q8eNlp1CespgBQF+xFFaaAG+9XjPpT
ahLuNjLxq1r89ZizRIY+NWoGEbYZPzoL/6tWBxfWPdtG9ujbvEsYS+kJHfAdyg1V
VXEBGLUSkvOClq5W63/IVyF2KAqwLW3ZWhkM57Dyv7GeJzAbawsgCi8hLwBw6MPy
AxIiQD5FX4o9tMIa9siGpi/IMNmLdT/h3ZsYopNOcd0+IQpeo3OuAbEPChUd4Sxe
jgDmNLEADnpM3OWYRLLUA33FUZhC3ZhXsFVgrIt/xS0NffGX30IZLt6lCt/84dLE
KwiSuvPNIwK2GqKenZqWTa1hPnOJUZs5t+6JKMvNo/qwwp8lSgwMd86Cw9HCnGdQ
2TR4p7l8rGsYI8MxkG2R+Hl7v1bWhYVwKHdtd1wx7FxpwJh5tZipJSl8PTZcQqPk
wyqWq3GdJzaYec8QGB1nFhegNrgZ9pQXHzHDACWV5q4cU+Ki+VB1pR3A2UGWggUu
Alz557FIkEjNaIBaPjL4hRwsI+/RBUfn3uLYbPgKhgURZy13ZF5VMHOsJ8xh3l/G
o6u03nNSmNJgkQ5H7YuM+/6aweocv7o3NQduo+zY/Wu7exFjA007aAw1E+BG22Ty
RGoQNlgGGEcqjOzxALhRV6H6u+7vxzQKwXSsc6BYOmc7Yc7rrJ3XjpQ1VinynkWb
wI6EzvO6LrgV3g+dq1Ipq+Sv0svZnlnrZ7obuQNJhcxq14hJ00Gq+aaMCoLZVRGv
mu0/YdXGBD2Z6Z+6xT7Azx6GJaLO27K+1z2krRGrwUXZIHgGVlCXhd1k2aO0olU0
J8E3YTVmgVb4Su1jZDMepumoOQQ7Pc+ucRkIlgadRAXP7SnhoGiGVk2WvYMS43lL
EuuoGg9GgVzNOA0vQCTVeB2eqag2Ll2hqB5B5deM3Gnp+mxAp390+QmP6Nc4BwXf
AtfHWO4PR2YH9SpWGffnBSQWsCNl45PzjYvRexiTBY0KKD80a7D3lSbB1Kyykxd+
Er5pMKs/dRmDXctxQsaHJGn6Kv25FZdmvU9r4UJkqpHiheRWhLkzQsIJLeY7TdrA
w77XcBLj9d90PqpRG2llGNSll5jMiQQEo3K6M56D0fFPj0cXpG3DlXLgekNXYfK7
6Ik/+PjWoPAmR3wx78N/c5IULpkuv4kcjY8uSmQcbVhK8RF4DXy/PeTTfaP5rrsL
5uXRi+qLk10OZChnMyuI4R92qziqnBG8tLbqMsMwSXAfijLAEvMeG3agyQFqfipK
7ZGnaH1rWBSa+kyfr4NYsrkI9SFBRcDKyf7w/ObP+NQ=
`pragma protect end_protected
