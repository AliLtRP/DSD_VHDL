// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TMEKceFVh6pniyv2lGUcfrbp/fO1LZhedNhAmZYWVgZ63fJdfSK7kU7SJ1vvXRAG
hJUSH/Q/qlqg0hFfGmlKTike0f6ONqiyclxqj895eLdbGSDLfPvFq6Gt2fMXNIAV
gFYTi7FJa5UKreik6J3Vek6Rs9yD/2ansSI26Fa2Sps=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19872)
Pc7Y1YLZ79xeFWwyJwtsgTq8RZbON5027LW8rRgVNTQRced84Pe7p+SNrHctZ5Ky
w0xO4fA5dNTk84FFu64PyZMVup+GOWCYGb6lpwSN9CLafv4WS72bEhErhxa7XpsK
p0MfZ/cRVa7keS2UnDYmibi+MzWOGI+fcGW4iquAdsV3Eu9TkwSusfV9opq0ElVK
pfuGnAKs2hLdB8DQJ0CzKXq9ixIBZHp9yy1f8TT1wZmRHpyE08W9cRvYcSkDWz4c
tC0cjqJBpLZQD5MyzThnuhjHVjIOgFfI3Gk27Qx3wJtP8jmqhcPnuik4aj+x1ftZ
/jvlCHMT5+BhUkyWbB1zL5cpAFEOz8G+sTzXz5/iX/wFEk6NLufpjF+kbmLKHrrl
PT/CssmyCBYwgiiidYwqIVgB5FxkW2HiYYkShi46Uad3Va3M2i2PgpywOhfOqAna
sh3vVsP7odWPADkWhg/bs1D/94pbo6KCc6s7A69m+WqLK7nQCY5R4Q3QdeUChK7k
uE/TUKpKiYktuCFxonBiDSqyCCXsubB94LJdjSUdXye36qYFUwO/vWeizcjo8fbF
/GaFPjZkloFrlWA4VQVyIkjPgvWTy3uoaJGfvQh8BcPrNBMjU/cY15eGV+T8ssrL
L9/WRc3VJAQJJd70zmfVWU+umrQR90ZNql2yP2Mw+ORWOtzki3IA5jEPu55DTsj9
5Z0A7ufQieMAx4VVLxcT53jcBPkXNhqhSR5tZPppMGDOoQcu2JZeBi0GrUD/XOyu
4sGhEUA1T85oNLMrPLwKi0Hs4WTAAFnVRqbZubHGx0+Qzm6ArZKTvQbbfcevk4Ys
BkwWBlQrtxykuPwZoCYqYxgTZX7cVu8WRlRf/tFVrX0bH2slsaoAoB5gj0yFDjSK
gY6ykKJSkQvlwPvCAYzoHj7SuEX7IZmK12zKyg9RWOJR7HMSToItBEyNApZbm/h+
1ERk8UHoS7RaC/XZxeIVuTepp8hQ8rQQhBtQIQasJHV6gDgIPXRMgKAxDwUKmKTL
mvdwiUskIcNrGjcrNykC0dHnjZIznyeXLSOkFmzeG2m7i2i3UMRqbqhbsSNyX0Ne
puuiH84fr1vSXWv7zemf+/23v8T+5fH9KvQedCKKoGMBhQWBl8HMG4w5fRsj74LN
rYyafUeIo5SjON9xljQErfvlewO2w3UOq9nsqS6GTBcXffmfuJKPQe5c6PAlMyjG
ttaP8k309lru059LaA1QBwTZ3MJJynRfTHcYAcP2V3xibTcaIvqMRuiaal7lFF1z
3DSxN1BfOUAz1nawBgPfm0hi1CzOEZsc/6IIyUKuaN+JQfBc46cTgYVl44d5G0Hi
fpeRKfpaiTz+q6fsQjTkG2x3rYrp2Kpb3AhRKPJhLx1xWsx9OwIl1kdXN3FiHuUr
IKZz2qY180v8gmU2Q6X+fO2x1ChKsNR+XAudljXhsN9Ec6JSzwVeAhA1OEQebBhW
ERwsuq48lZ3jyD7pEdtfW2U5s3EKrQ+CGCksOLI4ihWSIM9SUEFcPZPjyxE1dMTd
SqeMpjtfIx0Db9qCqdAcqyUVumQkzyaQf+auEI2JXIHO5P54EZ+ObRs77KDavxVu
pmA1QmAq/2jtzIoMkJ1MZ2r8/6lMZPw1f9fQXWaBlR+7m9aIcFGwF7X+12X9s4cI
/sbyegat2Okzzmk/iiH1qRNauf8reB/4hyQ2Wih0to0tDk3P0snhXxkfN4gYr6LV
Ix6yRegidx51RYjMUpL3bFGLiu7szZeh5Q9lT7rIi+9xkB7qbJD+XOd+Q5P6x+lX
6qtgU9dNxKjfSXZnMZ/UIOmqS4Crl0KDIvB0upVcmtHjDu5teKoB3yzRhpgAy/4b
cAlYHn4ibvr3rU3nF7/9C2j87tK30fyNDUgQN/PytksCRUU9BWoAhI/24yptL6oy
bAjqZ8qYYcyNPwiBh4GjK6ROGAm07Agq5+AFxc9tuN2DtrgRSG7CGNnjCR81f4us
bKrQ8w4jmrRC3VlSf7SfEB6nydI/27QhD10nsqKSHbHkbbZHvGaMj6xHx3qZZAz3
0AKxKu4aDX4HIvTop7e2zpCLPqygBXhJuB89vdmjdRT3+fg2o0rSstyCT4lT2f/4
bOmds2PRRmpnIYtcJgNWKmS3BUXbtK/IMOqJQdAwABYqvsPBIrbf3esbEch+dha6
O+K6JuW7FGoH5dZmGaE3DL2rL+EezPjtyVZAgZBDL5lDQbKpnq7EIxwpehWpNznb
vQYU5D7CjssozI2LS38cBfSsjj1501okKOdCP06Ozhu8y5Wlrd1rrhoqrCljFKYg
FDo1kl77tZL1+K+MOzFlxk2QDfoLd2QICv7Bc9h1l0JsBwflGK8aZeAvkCH+/roM
il9zOQVcmnGR3fJ4sph8SndJdYaI7u14NZAxxQAJ3Ag2TCRU3a2iugjciSC3Y1+O
V8igfjtbwRGjcf+0VuO53D5qWP+5YMy6s7hkGO6cnWdfOGyCuo3C06mw6vXQHEZ8
Opini8PORrnBmY+b52AHiPO1XkCltFsknzwkbfxPRhbg6EdDgPp20BIRKhFRMh06
RaN5gZws6lBY+ChpQBXM47Rix35JyD5Vo7reCWjHrbIDBjhKfD8ymKBToQ9yTAgN
vr5IPpNTcT2EdxZPeMbZZDwmdj3sb7ewagGD1Aw4uWbWdd1PRFbKmyOTWYMoxj5r
rK3VE3bqkUtdxo1b6Qb+1VjQf9Yfr8892ADidLHK6QECzqTgSqunZO+mFbMFy9Wd
y/7VFuZ2e064VpvE0nQMHMwgePkBBdg3QWnGNhzeoO2gOW9K2qLDTpeOff8Bjatx
5GmqhTCDVig0k/IzltfqyKvsFTu8ChMZCAyR4HLl6MDqfHtqR8kHIHyY8D6wq48D
QamntvXyxQ/uqnzjUSpy2/ayDLaCEGfJ1yOCq4PdBYFFSySuzaj9xp4Y7hQuOCpF
TpTq6ayTYkLe2FjFFlObFEsz3ssMg5e2VeT9WRDmGksqTCZQg9Hm3KflvewUStOk
gtLa6Ohrx/12xElZ2kmvwcKeJuFI66LzhDm7hM4Rz1F0hdi96Ty+o6JYf6mN0Fu4
tHdOUhuPNCrBQ8956XWN6XeSlZIvC9AmmRuUllazE6JRV5Wq4eqBcNdUzpvZ6Wg1
3SI+o/p/wf8kflsB1jj3fL4TqcLZzo6gg0D+EYbcLvLbqB5ZhRHN5M0+DHCiWBip
ZhvK33WS2w1fulHjcghjJ4ErByQ4wo3wEji1sqrN27vv67nDf3rJvyhwhFMktjAC
GKL83LR66pZjdgFt/MVVlCOFERCfTnaBzpIvQpkD7LicSVBRa6mofiKZQFgAmb2I
itPCU+OjdtU7Upq+c61UNss0nMIwL641gtck4NVldef6nLhdtJrtUSglZI1a6OVs
tyo5mtntQKYQkwsSK9T0MHfal2GE2tT+xb4WhuTeKanbET8yvd3Bo1ttnMmA26I3
dkKOIHsJyaJPICBTBBm/gCxpXi1r9Pqo/NL66us+Sp+/AUIoyKhOoA/jmjxkaKN3
36v0pB1bWbfbkToiEUo0xJ+JugDNyHv2Ou/y8UI8Iq6Z6Enjbe63tk56GiwPQ5WZ
4GsX0ypzvkjT+Dlj628G2QY3BZPtBvxfPfTcSZGM7CqO8Aua5E5Wj2CYlxtaJxt1
NxMveql+fUPBmhjqS8RugZELDmRq7u39Ux3n4M2DNvHJAzFlDrBj0WH9bJtH5EUQ
PyAEmCOkCLNDQb7w3e9co8qkTGpJveJxBH8dS6wi3NwfraMDVt6bOMdi+3cZuvJI
6Fj/rxCWYj5LQsYeoJFyJnuBKlmgFmBqHfa0ZsEC3k/7B2adSwfycPIVor8UM3CE
gR4ZFoDJu3TuRLQO12FZnbGFHgmenOG2aX4/SfQpbYPHNDUIpyd3jN3QwJVsaYFm
XirLW8ICS6Y7A768ff+1oRCvLxOdlibZdTM93meXa0ZHelxVfGNFuRTfQTA6Xvea
gxMK7saFVNjOqOsUYxe3Pf/+UaheP4ltEnmj5N94Ah7hr45LCkBwUzJCHOf3tsdy
7JvOJe9jbfAqHMSxzvDL/qDavWIGQ6c0mGc1K11nOued+eWwhKpSeeWagiMWN6fg
/7YlUv8W7jSzM1G3gymj9s1oGg4dDMozQO3Tih5hCOUHEoXDkHQEBrZAsI1Vw80U
XInHCaVGoyCa7Svf1pdR103qTGxp3bfUV/fG6d2AlZQvLgGQaHVt8VYBER6OH0FR
cPJAGnbGUEAJnupTOIPfQw750IUZJLsOtqcXikVRAsUNFFkpin9e4Mm1JY9CovsL
Vqg+2mKZ8IeGBn/z/bsBrwmbH+CiUuXS1nXCtjOGGXoVxK361cR4xcjp7YN7ji+2
UiyA6/x0hI20YZ5dIGusiIU9te8wWBdF9UqwghRBm2XIblPpS3miJOGaJx2BmazF
KpUw2lMfW8q+e2BpyE4JNtRR3bbBApxp9HMDKGHmwhH6tvt+vZDpPqzdM53nVgcX
Tu60K/YNb3s6Mt5VKxNIqf7JqNG+FBvarAXQvgfzR3Z1xtHb96glfVPHOv1tPzoZ
J9kVa5ELc0iBtdR7myAM5lTkw2H1LDYkmfjbq2pXVlUt6tZnGKmWGoCEbE6ntb+1
+sp8y0rn/8nEh2wQr/Jsk4r5+LLtmSFiXRkCAes5ZV+02rBtYB7eIXEspUms8b+b
a07RUHkN6bvmNvTdzXG33yCLk1/IDBUq1mukjwB+niiyBb2SIHzBpDStkeFP8dF9
lcGcZSKPTyhhWJeu3omvUOvgQS9qh96DVpT5YVg2o51f1OP2gJUrOI0D7XRHjDaK
WhvsGw9U2sszcR1WKLrxZxvnWM1x/2Sd1nS0eDY7Gbn8p8Ms+kqcwPTFHUOKtGmC
cHXqV9WSWH/U+67MPfxTqKoYgQVHzbfHishKlKYLcx5Fi7uax69h3yT4i+ZkEaEI
GM7R78fOHbElM4hM8cuPP79eEMz659+jgXDQAAs33rblvUA32BdHGEwqaEyjtp4y
2SiaKnf9n8kzZExews1uP1qMeCChOcD9bhECARcyaIWTtuGt0GlRNkfUm3dDMEPu
mUSDXC8DIKBmNXbzpiKLnZcaY5wgHgSEc56QfdwuT+ZCxrhufMX8S/EYzDyCJ+HP
Yk5o+1Qm6l5LrsUQGmygmrzAGbZCnn5v7zNeaqwiPmZmfrOpHXj3+PBDLTWPKd9B
2zilykMlIKN1ut2drEihSeDexRq091M0rlfnuPC10p1xl/iNu30TVvk48+SQTNr/
KxVRXA66bDT5sSA5AmKE/rRo/rwEeQ72K+/R7XV0jqV7+V5kNIfMLumXplSOCk8H
oHAEkH5jogV7B7IWFKnazcJrKOUN9BB38KUMphVXA9EUqb1zuAeXTd+0AckXSuTn
Rd6bVDEqQmxtzdrdAV55KZkmd7g2QNU+iSKbGBVhuwOSPWsWsj3s814r5QLbr3iV
e24phM1Yu+/M6qPjsUxLp9gXA0R4/Caol3tgNG9/liSUBPihWg46gixSKN30Cgbh
OFtJ1aJ7c/tGqB7tIxOghj2Hqx0FwWV3Vpfvzi6siepQFZSERj6VFkcmLNfu/Afo
/4mnpfN1zb1YlmpV703+/kVl1YkeDyYKbKb9jTg77e/Y1hbCTwP1NGlL1xpxJGlh
a8hZka+xsLKsE/b3xCO4AI10nI65DtrFc31e1Ei1xCzZ4kwVFPPCW1tecw4w+w3u
mOdqxemh9mcB3+/geWoX2CgFpNK3b5haEF8DIMjJkLAW3A2FgYXs7PmrSpy6liHt
GVUtByCDoHPkCjHOBjsI+/gdwwPAmAbrDA8MFz5Xuz0VS7LdT9S4cpTnZ/jIlBmu
ny0RAyzRgvGoPFleFs7jx35OSDnK9uGaDLjsh5TZbGuhxGWIddif9zDjPt1z2J/t
RJf1G/tMAdUIcMQ3du0pvirkSsY6SZN3LwHzBGlpe9Q+qxQPeqUSY6wOPNI8tq4S
+G72afb6NM8vd+Y/cKlYblwEWbHy4fnjwzWWf3hRh+m3eFWk0EfMLoIZax7cJUAZ
H7nTSnBE9foDVsio38qVmD6aZNhUO5JiEnPaS2d8Pnsh2u6jjSKtXHNap8O46fvs
7c2/Fp0L5DYod87Nbf/ecEYO/TenW8irp0WlHedzbWNcXza78tRnJpBT/k2b9lgI
wJ6sTWOHFMwwwGOZyXdTO+PnYhCcyyContDYiATd1S0o/ukHtlZtRe23NFd0SfN0
n0xIj3u3T0/AqyWS11JElbHTaQWnBPh4vmsY/OwNKx+pYTyHYh32ALjhppgdTOJF
u7NwzT5DlCHR0Pqo/zmgpw6uPEfsX+bEkdswBEtc+mnsqggT0W/xLkSjrtMV3pZ3
DQX0sI4Y+kofEJfhTg0ZvqG+8K54me9gGC4oLiu8wT+IqRSByhPMnKZ418jnCjOn
2NQ9BZzuis6BN6wsnQtni4rI0SFtyPaLAucJ77Y7vsNdOmve2tqbh1CzsH9LpYsx
pkfwZ82asd85wxvXbc9grEEN7yLTxLzfwGo4iZm0LzqeTB2QG3jPyJU4m3pF6qvQ
rqZJfJpndCimWhVBsCIMxizr4SI/131c2LwXWV1ScbRLp91j1LMjwCa2MIHL3AEa
LHFPIe/y3Uge2Q1DlMFz9qVEKhj3F3K/0kUaglSzTPgwtWRGQJMrQNrFeECH2mSC
sqiSX1VjeiOZ7prPsuZ6zG9lITqQLH3dETZtHbKq65SUGkyXAefhEK1QpsYbg93X
ENXz+dZZ7c4si8M6Dgc3nwtCJpd/M4cAle8KJsvwEkw47lO9XoXVMYrYnEPky0TX
MC7uUE9sfDbN7qgwrHZFPveHIBJF0+CtKm837eNYgXWBx645UuufkPxFJPD86EpP
M5Ax8dEAMgGF1v4CuEO9koOLjWSc7nglvqq1u6xTu/Z+BMk6ZoICf6IvCIAWufk+
JteMJEteG0kqKV2bVwHWDAKW6x23mYe3B1biTduQqZL/0/b2lGYntHniLCeBD0JH
+3XcHmYfAqfBIEecQejhOLawWNF4jjldtdpd5pONrV8lsnQJO+zyw6XcDvfc4w0B
qq0ITkAzrqtweDj4+NMMMsWWtxK2XMoIIfoflmgAf4oETRvtg5JkIP4MD0XG3GsR
wzns5b0syvl7uNFTL7tfOMdK7OAcmGAbkzm/So9xg8oN/PC+DNTdxrMp3e6ApgDV
e7tKtzA3WAvq9wyHU3jk0pl/nXEvK10QpLD1ZS7atP0d6kkdED3cV/bSiOcsUMmM
fum4b4f6xDLgpvVXjN4szuM8c3bfl9+mjZVOvz1BIUJBEJ7eyuQoz9Pe2y6y1/Zw
5h6G3l4BryAJgo7z2BFArPVeiJ0s1hVdoLsbBudLb+8jTpyOMKxDtHPevB0i8Q88
bRk2dCsa03CqF5yA8heiuG6AdQyE6gqWRhazYl6IdPtdcSdFreUWk/t5kXjj5hvI
gQSh6B0jW/8F07OTp2kYgVvfqfcfAaTfhRD2BrkFawMa3ixRKDme9QWvNzj8QGWS
gzmGBsV15Kz9M6Ce/H/ppr8r/bObSJuZzRAzgZWUwMSqSyh+zW/R7cD35b8AFyiX
U2FHYsQ4ay7iZoAwCx+Ci9CFXDRrJf5aXg1QDX1ltJgKNxQcYJFYKiauibqOyHkU
FHmZRp3thfh46p2Pk81odq9iV61Entof5KqLFBTh/p72+faYzQvokGWY0EZNoKiU
+Q7zzq2RSd+cgw5vr5blXCb7iRswVafxHoJ+Ym1GsLhMIo8l1bNJFbKBKOU0BP+1
kPmgUGEC8lJY6uAIc56j7PK6iYgQLIogV+k0md1RugZp/+uU7xiuXqdnztGIHnH0
5575Gh+gp+tkd40YkFpfzyjuxjsbOIvME0qWO9ezSLd2U3+NyCRsjcUemdPI454P
ngI6zBUdUON+nC+SPRrbHIUB095d78wsIo54k81KlUnK1mED2Cav/BhC9MxkRR+4
MvWxRulwS3ul6Ty8lMOk06Myy2m3y5CozIMe8Ws6bZfwBGZZgJ8nY74XBmuwGLze
K7NQwmZoPyGQEGnmO50He9bKAsbA2epHpJLZTaZvOOkoq5Nnjj9+JcTLL5d87YHR
yXed9RJPx+DF9le3hoK2IcSMMcB98AqIDNSLBvcZXPk43twAjBHcMmYU1GlFv59z
KiwOmkDz7SVb82wtEQLg89CMPB98KiyzoDMsfKn1NrSC009LbGEKBU0eZYuT44YL
v3x29mXOeiKev0C3vQwgnTcBqJ+jOWFVwQ6ncnOe8M0U/17qKDkObUcX7Huh1awJ
k2l5CizXsMeBS/C1gHvGcoWUMC0mfT/rwi3xcpStRJ/8Nl5Gd3luovS5u/irwMo7
m1n0XFz4S6ly0u6x35LxgWDHUOhVbloV0Ncp/q3acQS0ACmLi2iiRyZr2Cy2D2Js
hjrLUtQDu8fJL7lQcD4OU6bITTxgm5blVBRQWThqf9b9icAUyUg6qQOwzQCIRArz
aSPsoB7mPvQCHN3gbDGafpjOgqWtPybGEqWIimiHAs2t8hilF4ERduDZcYbA2g4t
ZoG71DEdObZiwBBE4BqaBB00bIlaPtdFOZ5cBuJvl736qlbXU59DS96H+nB/KiyM
zUWiLr8Mo3z/89B1uiI/xIBI/mLKVTYwggSGtyYdbPiQHCAb4KE/PCD7gixsASHL
2l2Qb4e5W0dhPmUL5i3cQDtDRY6604s4+dlT5TMe8W9nX16DAzZMHY4axx/+vJA6
NPFLofX8pQFtSrXMpWFTRRW0P3OVRaLwedzitOO6CSYUHjJDT/8+m0XEH+kzS+wu
8OZOsbl8jK+1YYWBp3kPJJI84neP0u2GpCs+RsQHJ/i0w3R2feCVTAhutRr2w1Ag
oR2hSZQpZbsfIiFpQkdYcosM31iWvkMKFMNuipmQZIpVJI3YSE/iBh5SNVCEKpPI
R1gCG9AtYG11FYE5W+hvs3zvl5uuJoOL0IovhTbJhD6/qZkEU3oHEUpmDojns2pY
i052RDZBTswLx4czMgKtTTwug7YYFZkyoCamjt1+cdMf0/qThmd3vVGTB+Nda02F
iE1Y3xY9RouWMz+Ab8yAmsYwX88V90yoC2uLI++arL6Q7gj17c6di+fqlN0dc0o1
7MCO7HqS4dWPjPalb+md28JzmWgI47AOprTUnR/cWeSyOQDZ/mrOQMyf7z7I1uNL
FEJeP/cgr9+/SzS6lMcnFJB6fPeMgPO0+67ufmuVYT27/13NNQATSHu2O6xlqQ/e
/PR8Gy1dDb7et2TD08STa+6DaY1jOGaivEzphi1qfLFhmgrvUYHlte3kCUuWdYmg
gxmyp3C6+/7WYk1rGDU8lXOfY//6wZg2vC+E8H/ZD/5A3shOMQd2JO4/X+9QsMIL
IPJ8r01wyamj8KF74LOzZ3r/K2yEOtvHoPxI9IykY1MrCbLk7BKfiUfQb2rMu5/c
cAQALE4keH5Mc8idaQLSG0KSu5Hl/7/23wapz66yNjeaXXgDaTvpC4v72JtNyAFf
HK1NFHaEVhvCrB5jFS4HroqBo/ZKdGdMZDCN0MZWA0iOzo8e+qaO2ATg69flOdDM
53vvPBj+xiVwqqsgCnkcgt1PJw4TLdnmUzhsyEDRXD//FpLmz9+u2elyw6suc68P
77pRikID60q5jWEiXP5kJXv2UjVeUF9wscrLAjTUfUybEggFrdo8xeHQGgKOgFaY
GU5r1pKhiZzFwjJvn71uKzvXRdQw2HgBUQ7xJ/eWdMxd5hD8tlM69Sv3mJ3pWqTk
cylZfI1jb6px0MaSKC838wPLSum7FCLAc9d1NnfUeB/wP9hnubgdNSYY/Us4OLYt
rg2L22LgSSheWd5XaeeU9TWIYMz6CIOjLOFpl8r12dGUDj9oqjSXEFAULh6WiDcb
4O0Ptk8Pf1jHcY9ynMNRW13lVosskDiGXEjwUfNAN/WeJ/GM2dpebFyruzA6XaXn
UtIVRaDAtvvhJRkaNs/eUO+FbtKf9fwwG5TbKVlD0vm+HzW8HhdkpMFiTBQyyy90
GGV1o/HpUxnrWjRxhlJWACPWLwoCFwwuKjVvCv1zk32PAFvXqQecoMWm5wYnPPz/
AI00eJ2EmepTmwKt6hdlz/eEPAfncEjGSfffMIutUiMY0Pm/RtIQWKc94aU9nx+a
77GkeV8rKMmpNj1I+L9BHnvEackYHjC8WBG8fQ25knI/S3c+XHIiglOTSM9wDJGD
QtBk5XFTejfw0X0CQPhkUMUQS6muNS8KjWor0qAJhC6qnH1Xv0VqxpbqRndTnVVv
kwxCFzLuX3usxWnqOpvKRfml3hBMJeWMPsrXw6CMlLUprcbQCL1ji3zp4sjz+4Cl
DIeyf0GM8/W6NwHfJJLr1rUBmod39RVrXiQtRYZ+Z9HJ9UutOOPrIJ7jEps5YJsO
jJxhZDp/VWwB/fkd55l/I3HEnQ1d9dTa8+0mZtYYKAJ3R1SQcil/S9jrlWDl5YO0
x4Boe39fUjAmjvAfzL2Ck5VqX3I4vr/CaQeCpSgfExOyVUDh+orAvzLTOxKpS5ZR
YFFLBcHDnB3fNJNenLM+KHa4TDNza2NqV3YkNDDTGZkGpI0zRQ9yZx6LUBhRYsBR
sdGcefXbiwRBmkHU30+o5tYT3wes1uT/Z3JFQqIbWBdH9VjR85tYjTocWzm9fN4Y
iYGN/SqkuRlno0k2XF+cMsnyiqONHJO7PZi6vtXnzaykXmO9DAe2TG+WucYj3P+u
ZEkKeTevNtby5KqRSMGCZHN15aWUMzgNgB1r2KGI1GAgiCy2ViFgISaCX3nEICPW
wlnl1dkMT4tNPXGzRagef+sqUU8EGqIF8aKFJCPafMnX4f5RT5S7VjX8iXq1+ufc
lQYciQC2IG6qXNfzjc946XaiyCjPIuofXMVQyB1zmxWPSNnI1Wq/fuYusu19n7yM
82gzR6LqxgMK0oSQ5iPDXNSftpmoXWrFZtPdMp2HMkp/wB5yTHHkN5gzc1wBxVnt
JcuBO/3IIV7NzhqcJKF9/usFFTiTZZIw4YcKzZAeRTtS7oqJQYx6pmL5Xrmd5XVj
yCE/zmA4pkCTxoFzeeOUccAHLuF9T29HXAuMNl4yd9HyVvptnZcY40P4Td1QF4Od
8MLcaRubp8U1LdoIVDRTx0BAoDOM4iHxtqXp5EkwnLABXbW13Qsh42s1yhApln8J
a9us6fdKH9raZYPD8APPTuKGgaV/bQVcuWdIy8z1LvgaP1+/vOc55vX1OxOpm9a8
niSKH589w63fFG3eEPoBfoIdkRMfryzxTpoIax2Y2WN9tuPaAJ6Wx3Ld44hFjLD2
CX1H98cqrxkZ15PgGpGn2ngW8k4kDPMwyO2O6BKjjcvy8fWfS+Atg+iTsESqMmVr
GVhNHXY+EiqAfEL5Zc7b3bdCFEQnFIcZ3jlHh/T6OoHq41FLpYeXn/poawPyo7hc
04o7FwxfZkrGhjqHMJrML8MJg6AGgZeSE+6d1c27W28cSVyu5U3DGwGpOLietPal
YiOFk7pFfZkRgqw4ZQg127XZEpxqaDgQMJb+hbQCnJAxl0vCFE9N9XqENAzP0MwG
xxVkVOO8Go+YQ7cb6nys8mMNhoBNL5kVwYm/oOAd+7mm+tqk8o6jh+hjEEaa4PWQ
DhEruvT4L0f3JNwHLp19OUQ60h2uLmtRmV9Iu9NY7x1GM4+EZtQ2hvQGmNUeVdgi
CKTR6ZRgfz3HvfJynMTxSaNx1x6ngxk/jDzAo/I9yferYoEe9A1wsjk82N4FcWNh
1dgB71ZC/nbZE5xZwnLfi03eKj1p4rzfvv6E0bZ7Uf+uPEDRdLUjQkjA0Ma73Nin
LKm9SRH3vlwf2fNK5da6upryJ0bjVd0buekcn+CCtuAsBVh4tT51XU3zo6ZbM7ce
/3uTBy5gynfudsDznF2bDhqyxEDwKLSRGKmpSF19Tc8syUR4N0CCiapDgtGpyL4U
x4Yu5ZLrK1Y0SrALujtl9rNYD3u3vPHajViQWZ+UHeiBdU8/IUemVBHkTynSsmWj
fotIcBgeHSAKAUsOmF2fwrJi6hggN3r93EjYWoqW1hUyQE5u+ra0AK2JyZbtHjL5
NVAnvSc1a5frdTOK76VydXZXSoe9lQPXGmMuoaMIetPtJG4LSSuseh5NZBhhQ94e
y7Rd+TCyS99fUiAotZF59YCMpvJmic8IrzY4K6fj0hl+mRM1D05ogy2E7ocXn6KC
8S/lwCkBe06X/8Q/IqIVNMFJK9Rw8r9Z1Qk4DMdRXY3G0ZxbGASAOMtAThvSqzI2
cuKLuABcuoe3Axs1GSFJfMSFMKjNTg32TSFgxI7ZPFVUA9GyxjK4TMTQBr9nYQSI
7PIHSw+cjmgDpan6SBhMot4h1uPYg1gaZ/Orn2zdThete7yQLfOdyp5yNcCFJ+Gx
9V0uHL/RxDCWiXgl30vKWfcnqHxypDdgHNK4Y80hoCkvs+rr++sAQQvWNd1wonl5
YqZ2RDHOhCT6NeelAUTEmcpgr8BJoI4QAgL79a06S6ddLkEgha4q+TtLqVARhw41
pi3m0gpCWTWCaZeYB5Ganq9W3pUIU7ZZGh1ifT1OpWKpDBZ0W7NlkesVI3bfE0Jm
yJ/t+4wpO1sPhkecmY2xckhrlytCjTOwYwsF4eacwK6ucAken0rWHX47AUq9EQ4A
QqAfZ4qmEkQlncaG4gcaadHbdTsrwWkLYIuKPq8FrrbeC8nTmIDjC/cexFnc91n7
CPvzmLVZ0InMDyeVVeJ1/sZq/BaEPn5YzTuN3u4Ikr0qism5hwNkOKUI0ZJ0orj9
qV6z11vsiJCBGL5CKPvFJeWBiPDAJpuJTg/xtfrgpWcTyl0fNxrC1CbCr+C6ZivA
21ykXzk3jtx/SFg1zMEg09tSKDZykLZQA+HUXGen7L9wFgxFfTK7ARbHkFL7e1Pa
QIfziebLLivIC2NqwI07Qptojvp0uIxWu06KvFk1+/r7yNMvzJxRUVpjT6YucNWe
jzafMzLC+2+DJSZVwPpDP7fErn2+/AR3NKmM5AK9VzUOplWD1uncxu9d/u0LGYpf
dEj0x8I0lK0uBzGz6PkNdqRfgFV4Mt0t84Vb+YGGs8BsEvRjErpvf8oJUtxFy5jI
8c/FlhUJ/TCe5hMD5Jid5JZv+mzBbCqocEAsJ5pDNAO37suNgbH41lxTzGnZ8tL8
nYG41IpLhNpAidRIG5fwK+zs3kQl8vPSw6pKQNx/2jIpXCfUV1+hS0swX3XRn0+4
uih6rZUfuaYQJd/nkDtOSNUOa6zx0jsNfu7npzunh7TH7PS4YJJANYuOliloS2Mj
7LvVJwjlrvd89j7cmH8KbwuPizLsdh0AEMMMoIvcL9mrzboxknRhvLQa6Lquika+
MbaylvJZlSK3+qqW5E74hCqKSfIS14CB1NJKQZZvHWyVxHo5DRenA8wYhvWigWbE
gWzgi9RuaeUMnd2qRR5VGIYzJqvz7DMXYztV4ONRKplNTTfueJR31MSD9WC1q8mx
IDgi5iLwwBuKShVShraYAMUVtqMEtWQ+Md20vbJHuYJChbguNQ2m4M893EhH8gls
EyGZiviYCdsBhemlvXNI0KjyWyCU2jAfJg1LtMSiMitoUJqk8dgAzk1FZ0YTaK+L
siM2ibinneovK2PxmGZgKCsmbAr6CAX0rmLDcz95lWszucrsCdLMCkd2nutYMfRB
kdN6cLeS5SZ4pyQcvGqxKcHjiXjzRUlXyZd8Dtmah6ne4CxRfKaMENFmET7ZdXY8
S2TG5fR6WwWhBBpD1TsVTh1+H3Zy1tearOMNy0w08WibSmITCDTShQ95zloKz63K
VqsULswCqbC31XpUyLrPEXE2kKznqtf3VN1QK/UF8aSXRyexWtJH0fFiLqzZKdyz
mdkb2efKMBgquYPPd6MtT/rhcVAO22tmYte3UNaypfKxUQm4nktp1AXK0JhdoU02
eiFbpsrvMjeR1rulOvHnJRvTwr22RqzksMmILumiV8hg1+lvLmTXf/dSqV20T6P8
szSYanE4OEGlOR5O+kzw+Id1w9pwKgBci6RTXe7o6flgv952Y5lQm01Zr7I+sITT
5eXpZ8wqiHYGlRtisnuZoEVcn5IHHMF3UviDgDdOOfCrtbWL77xjcucYYmiQTsb4
is/FVv6I/sCNZWOo7XbGDRyMyYPLqA5JPyJWISuu+NI+pPfweBpsaR/n6xHg4jGH
0uiWJD5Al/DAyNujzzu0X5H/Tm1SSGpmM4yFcpJbLFMKml6b9ZyZoowS21PrPJMN
Vzam08OADOAExL5pm9zsv1MzGCt6R3W0M/IokO6ezQk23nzuphDLWwufNHmoAjr/
liqAckQvd8tvO0cYLH8kGANBarUYyq6AoKo3aOeJsaeMuGKfC9d5mFGpqaqrXP9o
VO/iwCUSFqxi+ibx3kaLT/E3mv97cFVW40Zo9udxVdGJ1kNAhVeApJlqiLFnYx0F
+9dnFHAeRH+KFOj9munlGHCzpdE/gV3VhA7GwwgH3X3XIKAW/oLfzG5yVwXzuaeu
LAB5HVq4zdPs4CW2GBmJbuXARQ3F5KOaJYUaIBzaB0AWBlbCn4SHlVc9uH5I4JgZ
E1svcE9iPioeWzehhNunNk416rJuUm7pjPJEJ+bJMqaG8wqacV7iOHR9mswwE9Te
49XYO92xAZRoMvP5qhY1+3ffFrV31J2gQR9nJvcc1I2NCciGfNHZyUUYbpwbLj4Z
hvqccFcr5MRA1/eHeY4/En+f136ucuQDJfWSs0iKjZ/NvaKOoFUA1DH8/QZ1AShB
eCWRwiieUM8A7s9GEMlufXQnuJZmiAt0ct6m0oWcPgGrHb508mcWhB+0lDHC6of6
7voU+NbxoOsub6MDQOxUH7xhV5aF0dp/HLepF2A+NTvkeKQejNEEdi7bQiuX1Aj0
eXIDqbzj2tAZUcOoFyfqAGMu1OJlC6V5vVqXtIPwwEaTTPgB946CvZZazk5SYB0G
Z/xJSb5gpQzn1NpIp/X1lX51Sj5+jytpXrKRePPY02BOztqr81blyhdxFwlOGFnS
OhKhknMNeCjDID2DIhSrgzpBhtOAMPTgpktohPMC76R4ob4SyctAF7sVvKJ7/AcZ
pWgDe3Lzo9z/GWhDBtx2lZlKVD1kliDeIaw03HcuPINS4HejVk0IBsDqIjRr5+1P
VZxBZlmrzHafAQITWMbPl+tJERYYp+uPzsobR1/yBkXLIMJw0rPXBVYNFs0L0ZbK
Zb3Kdn7I/zv0bg80zoLWOm4iqWFM2W2ET3qwTgNvvvWuflFls4ygtYU8UTx/HRhM
Ajn58VWmHn6zoS9u46rvJMA5YI5tSjiz9gfpUVmvAsOyC88TTaN+M6aCkGNIyMH6
oKLJwH64dNSeQ2n1cpzxUhqf682ytd3BPQ+jgNUIV+YSKzaY8FBu8eGcieyqkJ6i
YfN4o9SKgIhXgMWNJeQcChpDuQpie4WSVFatkERu6T/8hsIk9K+PgP/g7Jzb6kzl
AiEhKbZ4XfE1q1naOKu1ySCpuZaMgBLI4ctqXXNDg4iwNfbLg2XLdKucpQBQek/L
ezmDAGAdfZHh9Uk/gIBJJLK2Uuwl1dpeb5/SnpNsgkL/dPwJeNYryY3oiFRojhuT
Ogdg4D2AAPMXw7A8fU8ASLAUI9aog7aGvZCWTknH1z1Kw31O4dE1UPK+HKJcJvLm
naangqBAR0DXQzm4UyxzTHKGsvAjYgY4pYKe+VCvK++pNDp22Dx8u+JVqNjVhXOw
BwIMXO0ru79x3RuT0aw377cWz77zz8pqFBW93Gjt2QXZdqhTbPCI0xIH8kDarMJ7
FSUzDh8iTq2R7sPL5vzHqb/+Q+Nbp7nchCT6nKJrSO1VqMPTRBipXJkxAp5/ob1R
BnObAlIUSIdOyjP7m2TXyXlLlJ9QSDFh3k/HdzLHZC/SvG1NQxNHw57sjCRvYZ0a
myQYCulPUGoOutd15aIhG3Z87vgQiL0d1nG4GSFyhm5h53HDNt+pPcctBXHk5AnH
3io8lhzJWnLlnCl7yejEufwxAdMkLrpFwVfm/F7tFpE3dtV63DDbdqYGcj1hisRy
z2VddFW+mZQ+/lX68xN1Q75g/riNTQZQT3yCeva2h58My5j/yq9QY/bs49M6gszS
/yYOpkVn+Bzhipv7Acnj8CSB8a2GNWqARoFYL5aNdYcdATMQdegHgfZoZb0R6sCs
u9KopyK3dyFHsyIeB6sKwVb9MW9I8i0SAhXHCuWTeFbtFBk46MtvB0esIT0OMQ43
X7qfJ/r+dZtQ5EOrwzXVNF3cs3cfhQbVCyJe4QpifQ0DIooQtStq6S6ot275ghUj
Nw196BeHG7/BseNd/326hwshMkGJVl7csd+rV2CXIealjqy/WsKPVypoKuVfOWxr
vF+smRyn0nOdzHaCblGa+qX9wiL36OgQZlpl5gPQE4FXMVLlsmUgwHNck2xVMBTo
jY6LRQvN/5jq+ndgk89mqOXexzZx3LLnoAWdbgUHvxetZ3+WMaWHG+4FehOELoU8
/WmV35X81Jb26lrhdEA7NUHSTHf/RTbaK7zrroI1R6cdHE7P9HY0Fe8DEWpdw+2L
0a0I13Pws09/wn2AA+BK2X8BbuMbljsxy9iEj2qnXSLD9WGj+ksUKxsQFbwC6rFH
XeVnV77j0irPpwNwpKwWKe+nad0x6l7+U7prWYXK2VEsjDWOHN73jVytD99tIzxU
aRCfsjW1E+X/HmNuBaS+9sU6aYVaBrcJZfNH7ZfvK9TmSBHWvj+93vh7QOUOeMrI
+yLLle4aqQvSYoTu3ypqVWzwUeh3Mw4nvZlR8lBy+oIPyMcRwWSf9/RbKcnbR54q
6DeCB4TbOMEqhibGc6bgwDsckmYvRkLk2I2kwBtyPjsAvQ8qplRrTVZuGcBoV+FC
E7GdwqoJdCvwWMbWy6vezHiu/KgKEEhoXyfnQ8o4NeimwWlDMxMBPBNfsI/LaYsu
V8yu6gb3xGJYGzIoyypqBp/S+b1qGH1thMGURaqcbkCDvuGlT70CjbpVAjJFp1Ub
p80XE7kxtGp20UGoaMZRfIAF53PQPUWkGRMNMo1OvT9p6b8H6dc7RmwtbRC103Z1
AKbYHHXE0nnwC+1cLZigMyujLJ7w+ZDY7wa3mn0BLc+7J7AusT/96bQjBmpzobz7
R4SlhKVEn1rKBmWHSos/2g7E9TzVTCsz48sxnxLR1dgi2u5E/1GXb2eCPTPO34m1
G5vrVu74/83XJTXzLnIuzUxoxOHKRhVTLDauwIAPdKjvwGEK5LkjQX28i1ackULp
mJvvnMjZcIb0AejwfSvz+RKh55kRHfd45cVCgYaRRs/Hhvw3uPxLYnpBbhUj2orN
yMdwkzOCf2GtyMEku/ozNIvXg2I7KjOW+OZOfjidoQVQ6O+8nyf/skXrM+Mk8kpG
HGB6SM4IJp9Z2kYU+mrZme82Uaq8BkCSc/bQL61z35pEgdkCPl5fh0RstmxR5+9l
EusRKDNJrKsVDyaX4JXbLd/nhYnOq15Vosz0wP4KyC7wJny8q7ewsWY3ZyKMNfTy
YJp8EbVBnajhm+3m6b6DwTMDEWj6stcCLFVfkUR2j7jlJQDNRWcciXKZF0ZP5QMX
zNPfSRySHcPi4n6nCGIcsEyfdz49WRrRnUYs+u/e9zSWILMgJrJ57dU+KBo1Va0I
/Y2NH0C+4w4jWlafoU3XgmWmDUjm/qz+mogP5LWOkFhAYs3vVTdOIcfnsp3M6leK
qvZug6hEDtjcqRXQxpTpe/Yi02wOV32DCH64waOGQde8p3X1VP5/vMjQvWRO5BvV
fhEnS6eAfgKzdA4GLeUprU9xfoi7oZJklVU6w3TozQ7TQo/E9XhaC38lFUpXKmO2
44kpyPr87fNsG7fsAgsPA1iIEubiFejS/pkuSDHhmyMhOFPwv+65s7X96MsPLcAw
7iuyo5KBUXuWd+1iG90m04wvNaNSSR/7/Bpm7Ajj8e4o1FuxgrYdC06HsGHXqPzK
P8eizbVXdltex16JA7KBoba5TGakVzyru2cTrW1+QLRUETltNgkckyoS8TDAMzJq
3NHftzwcMZ4M72iT3HdkDHuIo12cXWwFht8yu6+SuWdEAlhPbDclMP5bOPjmIrjj
3y7KBNSdOBuu/X4nSTdnQRrn1mMAYdJinTcCv1fGvwZQrDOshyfkfFWJMj0LKg9e
BmrHTx/uIyjtqEeQgUlY++bhTmPT2kcGmAYVA07yI11AIx/Io+TF1JDcI5G/0Pii
UVIIImb8BXQF1hBpSfBoLZVu4Smtr7p6besnzlqcg68cf8F1iHpGUyk39q221VM6
YBV2/r2q3vudvDh5PFdUbWAPV/SngFwycUKlxdmmtZvIoUStYd6SXhF3PfmyUcsW
h0VXUx+NGvweni8muGpM8Hv+OTcPcs9aR7QyLSSBpmfefT+jKIclElzzEn93tK2L
4/1VGG5iTDjiPA4XcECbBZrV5q8WvlcJk5kFBpQ8cfipKVsEr/3moIAD22FxOlfD
gf7QEc4YGhtEKq9wPVrAyyt+YsQwGUrxOG9YLmNX5wGVte02B4rMS2tXEjFnVUTt
MKvndzE9yP56zxKuG/bQkQxPkrSe/8tJ4AqujHBW/p9mLyketNg30q4Lz7WCSq8Z
h+FNx5jH8pSCj1fAUsizddrm/zLqB1xRviWovaUmsaG9X9WLsPOxHdQkqwbBELD6
5v9zI89+oUFrl9TPYg7CSqSzBLy03UWmw8K2hawGMnAcjnZ2JpM4mLOB308n6slc
lksShJ1F2dyN6h1C6dybPbBUB/Ne7WbkCpDPIunit2ax0E/SYiPrN3E4wpVMp4X3
QbYFy89gtM7l66GZnamRyvLXfrt3AeaQxH8kEsyetIU8ckDnP0faqdqUnmqN83sB
+UPHRUIFtUDdIQNNUrBsdK5olwTu4iCu36i/+va1R2T0TYa9OBw+mGyWpH0rQW3W
pHn+moX/+NQJZuH8fWvXhCY0iRoYA9SiFvYGxoUtunVJGwxSia0jzGxpgKxsceWm
4Y+W6JNPiYjleCRVJU2wOP0ujl9erYt1V5zz7j30SRzPEgUWkv6RwfAxAAB9ISy6
BvdJ5MOqJSc748S6EwIxD2Zct180P6//IS70ZtkwRcIz7m+gYImjMN5WXKhAO+1S
LzkVsicNjbX5evUj9fkHVQ5ZIgp28HF82onhV549uUPOunrYGtij+ccoJUuKZKYb
am/ZNhLEtp2LVE8cE+PVQI9V6Be6UmiadfnDYt0dW+Z3ReZFs5dGKYIP/8gVYDfP
0ME+qoq51iBCLrcKn/TcvSszE5vaUg7EP4Js1MxTciZe6j4kfdVnds08m86p2elt
plTebJTHw3GGJtrA0Bk6Sa+b+iIUY2/16NN9/RTS9EXIYsfcnP0nk8LzEcHKf9di
mK7m7K34bp9ltvK2pPlOS/OA9iaIrMZvnRF/FYwMo7RFmBMhZH9ankErb2Q6XhWb
abdylDoPGM5Em20J6db6PhoEO46PEzxwAiaengd6nOVIxRW9qUSlJ5stXX96pVGd
nZkqqXIcoOkHeGLDd+7r53SoFHoFZFa7KYArEHnSH1MllPlYHVKrtDwr5fxWTWfq
NR7PCr+wl2moUgRqmNn8C2cw2gW5UK2kVBVmrOlEjR980gTaZNRX9q5Ha8PNHFw2
j0jXs49j4IHXlRmYxUoFy6bYah9hbp5G5G/4q0aQiGf6XZonznS9NQlwKgPed51s
92aZ9s2rwxR4ga/1c2ljdzgudrvvfUWhLe072+RHddARYdHwuaWB55sVk9l/Fga+
k5V24jfR2uwmTuo+jFztKhHYjN63D6TeaOhVrFfU0dKreMmRnB1Q1UJeSpCS2+7r
BEMy1NfcFiAhDdc33kAOzE8IuIRJGAYObZ8A2wMb9Bb0d7jBBzbWm50cUcs8WWTG
M9pMUsS5DBZmanoaNWtRYmaJT6Cc4YWUJSTahVgDJXdE29spQjOMCHGQPWh5oAy3
Niu5ksm6W03B+xhPeONKfGTB5Vp/vXCDRMo1pVDOaUieZfwNib6GC2uLk+3kYrYm
AVxO3C4cur0Lg+c05rEzannWZT+5QmcbUUYTfIxasXeFj7ZZXO6q1h7gTNreQ5/Q
ZjEVhLWFiP2d21+gCndoCLpyWqWXmdEdRQ8qCdVPK6XPPou6wU9I+kVIeq7Lev1X
zmh5S4jXvwbrLgm28mGl7vfruLcdQLauFiNPSL0vJo224lVPFyFihnZIM2z5BIEO
eL2whWlQ1LBeq+M4Xuv7wxHjTTLDoC3TSsGB0wEjqzS4ci0DSSK9+atpBZsKyQ43
icsTVUfDab+vMS/w2ogtWO1o104PmeTAK65wtihc/sHUtcKm+JiSm5Nn+CGRBnv1
Hwe9mRkKpp+dkthYll37Qty6G4zsWabCuSxjLK6oFQOnT5lNgnfh0Kel56iucNj9
9mA11U4SWMIea/i2Am+aSY+RB+/mY7WPo4amP9HqkgmJNpat+6z3df1Lx+5vy+4c
+6DSfcArsLHf7Jyg3MvExWPT9+td8pRghmjV7Temk1Gp7t8pBFJ3UHbnvqUcaBeb
4ifBVhdaPofN060anD+scDqft10MXAB391WS8AHf/xhbTLwnD/6wehxR8geKl+6W
945aaO7p1UJJWmE+njwG/3Gul9iYc8w/Z4c/+i0TG1QAbaPdqdAyUlAtF4GUHR3L
SMbeW+1PKHZi5gthQPSMCtD//BYDvB5Rz8zgu1rR9V2c3IT6/txks3l7Rjj493kb
OsAPsh3a0LusEmNzHQR2Dqzskg/DPRpuF3urvSisqzH/P+Sw/0uUkhK8dFBS1eM/
ebca1q6TszH/vCkK+Ismh5u2eV9D+tte4HTVPj9j+nM3aw3nHrdlvht4fMUzkpS7
SdsxUlfWo7wcHJs2UyUViPWBt+Xk4EmzKYl9MDPPcgCLv3V+z4FttF+4Pix4Zrru
7hPSATGzVDDdySjvSF61F6U0P/Ml3HeN9pexFG6gpmkteTSTZQTOaqq7CItVrxBi
evG8CTGm9QbaJCSK98V6/wG39tW8hulMhHOIdJLY+4R2vJxbWe0HqLAxJqBc/ORh
y/UjMgDWnpYz5/mpx+m1hekAdkxtldJCXGxzo2ci7bHdSRlaiGX/aeZYakeeQTfC
wEGTVJfKtE1Cbpm9UEYZ+Yf5/kIhNNAxGA9dVejU8D8oFomBS3uN0SkSQD7c+2mR
bGGfGj/G9jzI0WJiUIX2ex5aqLdN8zWmKjZt47KggevwitNe9n8QLJMRLOzAuJJA
6treqzs2eroAX3tn8qbPkxwaX5qd8VElSqJsIw4ghBtbHn3F90amWV+5C6lAOrtO
KBP9mAM+oJyUWda7X8xQ+yNfCDgZ+pn6enKXTV6nta+yA0vjO82cVU9nQr9ReoRa
0Uyiwu7DxU/1wlwwrl9RqNFlcgi+5g7eA2u6ugIRgVg7EnN/7kmUuScYHdzW1AAV
CtM10xBbJE7QbmXf4RUtrozqOtDfpv/gBKFgVn0+RPM6Ks/7IJ7y2Mo8x7AlQmRQ
upnt8K2mxklXfMo3UCiy8PcBI1TeCtrLD+Js19rwOArrXTCZFEk7znDyo/K2i35q
Ybjh27Q2fd3/hA1w4YXiG4G6GRGnh2uYRwA0L9xkUrmVHze4svNCBR6bveh18p+P
06zoDJMT3RKszYSSDZoYL7DRt7noceb9b3955jyJsPGqtZZKs/vJbrSn5eSTxNQk
QdxshuE86rz4juL18SrgV9mRx8qfjZSZyA5JAMCfxCkXNsFbOUKb5uodStsdSMsC
KiAZCmcSxYH1kE/ft6vK+uezoZsvBgh3H7pLK1wSGCJ9e4DZ8WYyxlDbyKksknps
DfGFlFh8u5pHbbcDZRnkZP9vQ74M9tdMVUe/AGIzcLxbSfXkHW929RMSVoIjcVPk
OwMG0++F+b+esR/eCXTK4JEgt1JbiaGeYqw6+Ojb452r1PjGlJXI4CWVNnk4Z3sB
S0bR1KJWrYq/H5NgsuqM6Dfj8ELLZ5kBmTovtCo8cddJGLEA2HWVtJw+XumHQjSI
qCJqjWWoaBMS6WnPtvJKXYCRqNO2W0DhBrMcYvtD1FAQrMWhPeWHYSGj1z8lMFm2
xG2hCmpP7J6rtyetH541u7TyoTP4FjBXINuzrIgC19JRuhdEYmJSpoPUq4BYfaXf
TXtjHcJmXyAqoCdQ9dQUvYF6CN2dqDEB5+r1Icjh93UK/nU11eY2HCUknG6gcQpG
qQneFyrPpkjkZQ+ZBBbTXzJK49JZE9LwHVRfhENkk52si53CPuAaTVQv7KQG/WcP
aEao1pqJjYNO48drFE8X6lNRlD3eKsElq74OWnfuAzdHsHLqU2Pgy7jivlku/PcW
UZt3BFY+G9e70NKRYDR+bz2tSq2RfW1ih3d/1TDOwH+lKdWrnJLnOHmjaJt//ao3
WlbgtuiXwkdMyRRPbPT7RsgdFBwqgcROP4XiICsAiP/Ko2NFbxAml4fMgo/CfqFY
IOsDwcYVxkyRlf3OxOSROSOrebkl5gOJgK5HsCeGSVqDYD5WKaLqdkupPsAgQOWl
MiHa6iSUA7MsHkx/YpAT03mKAwPEAuCTtd5eaxDclq/Cy43UzRyIhwjCQczhcY1w
3Hgh0EQtgHOZM0uZPhGgw40YuZ7bZkajHuJPttJQdhOkSsX+DkA+gVrkCZojxcDz
SNnwMC0Styng0yEQZX5EYTo5SImzKilWFkTX5+OIGoaeh1YGQk+I92OAiEButdev
cay0KHNUkZy9d0G7C+kkvVJWsbgNwbJYyr3kEclbV9p9FpKUALD7X7ktt1sz3AB3
Sw/DlYsSQlnKlBgJcm+Q38hvrka+eR1+XA7SlKpzP0KoRQJS6CiHF06esDCDPaDa
lmDN19h4nCqDdQpSmbFDBw2zZfXeoJqYtk7gfki7hVTh53FDJ81961OCmQA5qDb2
62AI0OBgCNXUsO96eAcAGVZFdKLI/MzaM3O4R3y8KjV4jlA7JMkZBjI1URMJIAAa
sEnBRQapBRy2T6dHW4sDfAvWTQDqqR9JaXuwt35Q3siFloAtUNp6gu46lZK8RDpe
QFiizogPToeX0X4K7BsluoKJvCT5tmDG0x4IST8XmaAPwc+wszEQWoKGHhAOiCSt
bZR6LzuSoVwssT9XuNfL95Ks2QT5GQioGK+Z7mbr96ttQTED1+4y5WnSUacbSYUf
j/J3V10lczzImVpkpNZN+UrsLGxIg0Q8HH+nelMX3t/v2acGzqOPr1gkzqERcEam
QE3smpYixXClu0B31ISc5/ZSAJGJ46sgtf1x/WQBhpQF1V9vPnutLE3JmgJt/mlg
oeZscLioez4kRPiXuyPqN1fzgePJ0RVrgJoTcxztg8t3wTVLcDkjsOGbIr65SmPy
4JNYM4ML4G1jvQiMZCrMbu434XUEu/zaeu+rytrtg/+ZpLhGoqCULKQorDH3DkA0
8fHP9Cgc+p9TrM1jMIoo8OClzpsemcw/u3/qXAhP7Qp7xnXzoqxWD6HR/tQjBtOU
UF8xjQShOqJcycKPlTfc6yTRsmrFNyxHGZUIr1NoJphklCmel/6LYVhkOihOzho4
TA/uWrR5u2aCPG67Hzf5O4lSb5zTteUbcO2TEl84xmfS2mCOH0wTrB4s+OIP6XSL
t8VnQbwnnu0ydsLzDM3qlNWP3zPP8LCT2+KCLhvWIYv3s4MTdZDXMMzHqDiX7R1p
dELRVhvxjmcmzLA9E41RQxFk3kpdZstHyIVSXK/QnICyOuq7lC6u6xyrRI+FU2QV
EU9nibeIYYjdGQv4rwfow/nqWkRaj/ptfKvws+acoVdvXcAqqEMvPJZ6ovTrET92
gYRSnDOwIdxmexHLhaKDExodqBW7QWXoOcBWhgC+t3VeTEOV/APfRAs1xCGtVhgx
EhLp+Z9uF+PHpOB4PnPH6kqU/dhLmqJPsp/6Q2Ca6XrmEGXVQtvwS6nrCmEqIqrg
6+nga5z9KgHcGUNKOHfT3uteIwbYHD6qU6i/8L+kXY4OotDRzajnZpPqTXjfjgPJ
UqdoQ/jXnOJ2Kr5rIjgHdQmLQI1fJ22QiykTD6V2FpJ0+ueYmDBbta6Ds48ybIh1
gNEIb1bqRwWYcjM/FR2fjP+flLoavKbS8LyEVXlyyCge6G7Tj2xmee25A/8dsySA
Fez8a3Ddo4DalV1d/FzwiJJpZVQzL8MXbygOPqy9HV0NdLHc6h2hSRjZuiWKUUty
+YSb64lVMQrmH6jvvFfa4mFxjCYfnVE4OMmKtG6y0+XN0Wj40FNgAfUWC5/wKShd
KGdno/0Pn7ffYsG8IhUV7lzWkgLXi6Te945QPQLF0AgSt8OAiBeyXV4Ncj9AmFx9
0lNXtNgogoNIAgyABnkxTEt/F0L7Ehy2JwUNmh0Y2QygA65lv3H4qAiQnG3gC2no
3t5Xx8JdLkY3oOgZCPAwR6ULQhmfzluGMjr5hAcjokpKVoIh0MJ7qo8fyda+VEdi
R8MuZNOkpPzBsw5hD8/fQ5LnfXcSVQs2nhGBsMICXAbkcH7GnYTztaQ+igAbldg7
/YqWl+0qivYXEyNlJrRIUV5Y8/N+s22sjzoZVdS0L4tR9YK+vheJGjYe4t0hWNut
nW3NUnNDvdp4N5x/xRSmIaVN1dJ1n/n3RDdOcFDayVaAewqLq8IT+hep0KE763xK
vsBcR5gxTDxGdRGe3aT5jbZlvLixuANt/WTcfMe4b6Yxolt1CxD/DFok/1zNkGOF
RiXGW+6GSqC56l7tLkiCQsTetRCjyBuX1Kp924D2wm8kla8ew0A0ywcbHN3m1pjT
z9tblpR7ynhzNCbkI8/XRjXJWHacrGqOwHAvbCRqe/SusIi7Mn4EDNRwErmlQrbr
RJQlrmv4KfJcduZkVu5yWFgEunYXreX5sO9H0uLW3PxNVZj+9yvk9JLWtp6F4Brd
+CBpi+8inBIr8WtxXlZBvwdxsHWUk+PW79KeS1HgGqwDtA3dyU33SplHWQ2Uv/fy
IvOWc5fG3tk+OhGgtHDOSON1NaS+lG8AJwcEWjI2+5irWtkSNNixRq6I9B5saWLS
+niruV7ehom8iaat0SUUVF3uQOoqcCBUhLHFj1ISlC6f1AdOFUwy2Oaoe/wuv4Ou
tRZxt4WEkuPESMvDrvGPQqgG3XBGl58iol+YDk+vssb+r76+R+36nTsrcgkxpYam
9UZ7lpcw+WOMjKO4uFhHVrP/qfbTQ5fV4oyIL585cFZ/HStdvGYyhPpTckYF8f3p
ztFT8724gwzvOLAg+5FQQ6I8XpD2AgkP/q2TsOhZaeKLN5ppXM76puEl5Fv8bUGD
0lzPR8vveRv/V4OS1SehBfYVJwT10zXjZs7S54mJDK08f/ZLYxCX9RIO3F0z+2Fl
3dUT5238AcMMp8QFq1LyhktL9bIdzqUxFIfoMmdhAOoLNbKT95eLVtIc1yRD6k54
lAdHOub1gVop/flRmNvuPf0k0WJkIDWbvHrq91vZykTnvtZnD5SIZQEz9FLBK7MW
Z/2A+iJjIajZHO6v5HdJAysZ2xSSM6lWABgAoNxisenKdoC3U9mHUzMoS1QJkQol
wMQCn9FAlMbraEoNbdLhot0kh+ugmyj1+cc3pBqVmGj0qZhIrrZZOeLxjId8mvZd
kG8IVtCFRqifLYkFX0Z8e0FLw5CGvjoHmHopCdQRHgO5Tz5bZFGjAEBSV3FJkVth
ZzHVOKIa70XH3T7ZtO+BOPm/7nKJB/u0vGSM4Q7KLjXvJVC24Nn/i5cRHZFZafcJ
ZDhuBx6k6CK3HF40JKN2Aa+xAVPbbQA6jzQ0WXQ7gH6S/KaAKDXVaiePxgT1BTy/
zC2uh7d6IiUWN+yr41G+ymR0djq10XBNQLKoabzgZEd8Yy9eIlvFlhpm4/81o5J/
t2BywRhFepqM7alwtiReqffP8RZT/CCFa2FAugfGJuV5Vyr18SesQ6kajwPF8wSj
LT5olnUex432GDtEkxM30rwyTIKWaI2jmM1x5NCIi8VcSbr4vJRUwpNV9vpco3l8
mU76yocyU+k1/uI7vqu30lMhUd9WPsurGXKrxEaqi3hA314A4qSOPLwVegDXmTed
G1jbPsdTi6xDFhCJwUzIFtEX7vfRZabexYMNycpkJJgNlT1DrrMnCsbwbdDF2D2T
PWJE+h5WkG1g8w7XxTLk3IrT0fUybn+KjPLx4xGXa9d7ckg6cKj23dqvnJzzRtmH
GvKl0F71FrCNDoRjCf/bKCFaWx6TuTE73cy7rdySu5Is5vvRlV1PFXjNrqTuePLV
Rrex1CqoQll0J9PnbcsJBcp8HsLIgiN2igyhrIImARuJNXk7B1kp5Py2/taTH5Dz
ybQk9wWDLkHN9VXqWrJ7/Vp75iFWf1rrUV0YPkyoIlMOD+TgzD0LqVEZ4LPw9F+n
SzLE4YuxvcXW5Kt90NAg9s714S2a+7G0WK+Gy4HX0gKW2jMK2mPgmos++vNHoYgg
TeWjzizHxnfAfeqbBWI0dBP+Y02ptEhkODYhAf221l+T0/j4ek6HP5+f1KrMhwEw
tazWd43CwGT3fN91Mahrtx/ug+gy1Zj9+qMM6skJa27fYgrEvECVgmb317+r+g+C
`pragma protect end_protected
