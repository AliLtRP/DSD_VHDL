// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GR3DJQu5aTKNp+P7BRXRhUIt7aF3YwbnRrEtB+fCDOjaTgGIB6sxMvqRUGdFc3tY
+9euo0ZxuaJzr2p453J2zQVt7WSdVpeEUAh+uHzsEm5IyjQVl77QrAQOq0V1BchS
zflLZW13d6p+gG7lvC3NgfeR2tNjvJsgSVIthR1Fwko=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
j8hEN1dLptZaA9H54poidWHcb1iGeoXpjdJDwvLc5rTjX9PdjrgYzCziTEbqe6dG
nbL8WZPE3XxmBEbIr1l/Wuu4e03WVLWuF8uSCBc6iHKFfUUuT1c5xc2M1hrTp7f/
1XQDOyFRZkunJ81hsRGoaUym5fmCW3aMHthvmKQY3XQSSfmdiOZ/fb+AYGpw4tul
bm0YUvO40ANsOuEd1K46Bk6UaZRTTI4jPGspoGuI+Hz1ytjEu4EYdje11nCJjZWt
lJFXzLIYznwNYBIgWjRAhOig8pbpLITOMIIohGHFCI1iMebtKYltYD3nk2oDNZna
TQYpUNzg39BFvcDZg6ClePqxwc46XlUmGzPJyo4zNskfWHoswRk0GPePVt3rZvv1
liThKMCxbhGsYn2vXEHrqfc16o6Vwr0Y4iUK905rS8h0Y3FzWxWD5xt16KGLqDbj
yCnlXOuA/1pb/0R4D2YhZVroegnML4HUMp2If+df9qGLoAHCNUdYRCNiP9m6RZAc
sGzaQiftbbhis1OPGb6eVcudtwRTISY6E/zIeGe3vBuL6ZKaFacilqePCfLS8aLV
iJQLk2IreiE/mCvpfkhHDY5uzu8ej90k3yofTb/8xHKtWTjl1MQL1uEOAzlx0ymf
BmKZx3Q5XY4V5rrBvwgBuNf7sksJsnjHrVgqU3t86C2venqj4BiNhXS+kHfmy8dq
XGDgLBfAimbKTjKSGra38AqQaXf776gugNSAhKOvYEocsU32xPmbm5/1d/gjYtSA
1NEsQLXvFaZA+xsbwDL+PpYovXvSVyd1cuHtXCVNS+DXGZM+8MICtCfUNTLDjqEv
knyAwSzaR2x3NKYREt+oacOqAjJs30vRwRYQwL+bjBgvBVufGlOzBPB47JY+Z26K
nMEML8rzg+lHQIR5Yql33+foUw0EX8a5DxcebH27tGw09hpvXEBt2TToHnH+E3UU
iFuNQA/fBIYUa0C8HOGHz1+Zkab+rP1TQVUeYREwF3JMELUQSpbERh4p1RvQTB5k
o18tI8eVTjpfT9I2dU0O4gT/a0INl83mg5NI7SiaLaSglsoT+Slt0UkenGBJfK91
W5z+ScJ3GOZvFYfFvrzonal4DiKYw6+MdyaRhTKAfWucWSuDzME6VcUW8lgTQOzf
xUSAzLglm2yehtVO3jkQMxclqNEblZyz21znySQmmlfNzNuvV2fNSv0YXrqMeeGa
r/HgDCcibqYdeE7HIhZKyiP9CnPTrrB2+347RI4dYvU3oWGV+S9Ld08En122cPkz
9924ggUqkQWhXQV9ucnOL4kfXB0FrcRieZ2YxjHfzxs36u7ca3JPSlFtNt8rCgZT
8eFDSjp0lXxycAq1QHmrieHhvuWqjd77hY/HiDejeECrG+Xh17z5mUO/WzrQq21c
CmOFBlgEOfDijgikbQP309gOLpsU22DoGcmTKXJnmdeTXyPivSrEx/zkFD7zhyRs
nFHjpiPDo187NNLPK8MKh8vdOqIgrmsiPgb686iW1LUzbQs2m8DNbiZ640gtFEYA
rk9yyz+340BhSfPYhigiX8dgn0mDfk0rmj9TVv+C6MVdh157lojhCEK+KS8XzZ2N
Yb4hp2BzuE5hedyceG7qOJhA3ExBu6e233pRuQxtjb7l1p36XrX8rYBhu4/073xp
YXhRRagM91ZXKhC7ak8BqX5kljKamc4CwMFNeKkSsRAEVZStGMuOSR2KPCv03lvm
8cYpLmoJJGSkdmnaTgA3NVKXbowS/9MWgN0X8J+1kO15QnD4yU8iYd6hKgxG/B1p
ylJM9XIBU+UCEKMQrOI/4+CBm1lnN+kUTL4CyypLmGAzsYAsSy1bA2pIEQN+LKlU
L5yTV7uInlM2vXrvE7V9mp2Folvd+ZzuGGYumY4e5bkRW3QRpZ8Ddsq5guwE3i3O
7YdP4HWe7wJVudSo22Y0tf53DJXGJRCcHMdZ56iWZ2RDh2Wm2tE/kF/2OAFx+yyQ
A7lkfaB97JR5d874gMLXe1CqEPhPC+2FJ+55bf1aX96mnbv32x9+UGklX2TgSYa1
EMWigbej6W1KaHyDs0pVUcZjuRSNT79jR1RM9Cs53LXeYBzOhb4jxesje1iFAV/x
A4js5jxd5chDiQCZszluMWrSVR2lldQxxuDvIWXK6UfLH8nTMDOnuHP4I6WHxLxf
KOre2UghacuXr2nMO7ibQ2P6WkRzfLOKRHxxS0AERR6kPYHIiIjjutiyLaFRu8k1
vh3EWrra4L2mKzFGzl4Ws+TE2gNDyTkOW6sijB21S6dEmjOBddnGsNxuTfCdoLon
7ewutxHQ3ssvlZ1/R6PEv5MKxSbGOloTfr2FB0krFLsdImwiM4THxBhW2UYoumlM
K7xcPSv8liJFMI1V3LfHN8qFJ4Y/6iL1jurAJTpoW7APizfCbfuJhpmRQgeq91KL
WL/F5F7SWQeacdrS0qnjQhvH6eXyUrKmXCJZhQRJ61LZc48VbZvVkH6eAUH1OXpe
5H+6rtehz/1NFAbLdCSZO9JiIRsbrL2dMuplSF7gatnfTLkKPyMEGxs+umIvXY0I
qmHwKAG1KCSTs7q8nFSWPiZeLpWsIoX42ZWq3NYUJ/YmUBTWHOC8UQLdIsA+K6Xi
mAnrybbcVBIJMDKOjMetT7erQWp97PVsLmP/Q5ujOSZWjfA7fWqis0OqxgVa/tW0
1vtP1OdBOkSNNUSiaZhbH1AgndiZj29xnC2aY2qm4np/ozf3OSvKUuiVW97F9Yad
8yoyijOVnjNct7e3J0/yya2F0CvbInQ+S7mw8WoQF2fE2nUxeJnl/znY2TuccocV
UDW05dN1q7he1nS+sleyqTHG7u8jrLFPWKVusbgvyHrLXakg6sE97sepu1885USI
hpVXaKjwr1P+3CbJYK3mN1kqirDFv3cANfz3B+2sUN9Rt+x1VYkRBXXqP6ppB+oP
DVmX78Vx/ws2dECD1QrFLPCpZfCYL7BRN7DSFvr6mk1TP/6MN8SZhwnEgYAL9c/u
yfI1HSo8mj7shj/LBxr+To3rEd12t6Icjt+Qz0fOwP3+akF8lZipnXhEsW5xGRC8
sCpE10qipeTbv9KyjV2Rp/T7g2QsjYSSguE2K2h3WUjLNzFjXNE+JUM0mPXZo58M
55tHp6nBpdvjTujXZ6xXYURW0aSsQfcOk/gNabbqQOtIVWwx+cAh9ZKCpLRZP55l
yI8NT2NdpNy+pAMKEoWGO6qvyjLMyrkHJ6Qtb/b8EOzZWC6/aEDty1w6lLp1WlJK
MJ8ch7r5nzXBoQSrw0f1PETYE4naLDeRdOQg2XNCKf9tByubto2CcYeGS163hFRD
b5YoPWdXZhFVgawAHi8i1CGPgAFk2aHBIglvBs93jrv45eIMnl6LL620JF5GeuzZ
kZBouSuuM4t39Hq/eMHRTX4I4iEDPWDi8+ZOyF9bA5rSZ+KThpob/tm1c4UmFaaI
RoIZ/5yWutfpt9eSr5hTNuMTGcZLtSiJgAl3V2fDV1rQQQAlHx32mS/yac7b1LDg
0RtyZzF62VaJ0au+USve+VnX+I+XXy//2qauvit0oQ4uTKhmniZytQdMZ7534Tck
DJGnBKfBfpDl3UCYb63AUw3doY4rbsNqGwLhs5Ih4RpQ+IyNlTqqhsTeyl1MweJZ
ERMzgq6dJM27z3Rr6NrTfZL1ssQhXsD3O2WuvzXVdgtcfgv1SYonHhE/PzJ5lts8
VqNmnbcJQ9Oud1jqIz0GI7mItlHtM5WHmGX2E/Fo+/ArXE8FhasOq7ZRs4gXwThD
n41yvHSb66s5AzKRJIBjlO+mxPR7c9qeC+CLxB1UYKpIvrCcaVjVROieg3ETOE83
VTi8j3mMlMBWu3CWCwfJgY7kw9fn03i4vBGlAGO/6RdfwjStlv9PeQPQcAKdCJHi
e/T2bs/qSoAzg8cWpFPPRSpJiwcpapZIiiTS/RQIwxs/IeTVT22Ln4snXRCnE4P5
sXp9ehj2i1jmVRybhvuAKEmW8jdXYtS63N/PaFDmx6hsI+7dWGR0YG8qorkq15A8
6QESC8ESZY1YGKrD2oPFUg==
`pragma protect end_protected
