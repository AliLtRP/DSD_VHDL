// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Ll2KRpB1io3VUpJ7IQxdPsPDotCHK5rE949JpVr7jey3n5rKiJX04HDLuehxdANUnLykUzBc0VRU
CyNwIpxzrON1CDyzu/KfP4R7pkQC6c+FsyM3TIo0UXvjRNMgAyvdv+mQTG7lUO+is3WDWSBeiDXf
KATEsj+lhJqPgCQP7Xfxd8vMRcfdQd7Oyq93Hym0ci7VV2droJQ0y+jmtm0gn+HEz+sgt/daCxn8
huczjvrMayDNb3PtSIiJxfgzu4elAtzJh0gnC2YFIpp0iuANUHlxtQk/tJke0N08VmN7pxZH+mor
uUWHSDsUL6p8Egla7X8ExGvpQMR/idMi7gdmWA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
u2Lowe4ifEt8QJ+ZGoPj6P3afq5B8US/+bv5DfRzHc5gfTtHv5q6G/FAf3vHzZsrpMg4W/Q951Sq
3R2+U9sJ34qw2EULjCAwUL2C4Y5uqO3u3EQgJNBVMtsBplsxoM9StwYF8FWwI2tc6A2kvuGPYFtb
B+3QqJgTc4TOSCI7f7V1WxRrMzS7PqRs82BrbHdbKr2cbL73H0E6U5a+QfKgVdCJW6f99T2IOn/h
4wBnIhXFAP6/OWt6Qtl0xNUDYCNsARydj1aB8q21MCwO+NtM8kntQPW/7tJq6FxWfiN1JPis0v3J
UyDUGFGUzPc+nquSpd/IsphLw2KNKZrsPt4QXAdWTgcoDaY7eg9XME5VqKtic+k290s4OmbxyvLU
X19h7yjHH4KzpRLZ9HaU2yMkhVS49eUimmR3LEr60Sbc0mk3OYe5bMANQAUXfxf1mNWp2IEASkbX
yF+3+rQ6u4YEhVQ8FNMqAycQGiMwGf9mmzCQXXMKwvxO5bHP41a60peO/bodDn2mYrDOJm6ec3AY
+zjTfGA+PcneMqARWeB7ivt70+GDF0wf5H7JsHgeRJ6gMXzoamWAHwEfLAjJCtQqCr/mdk7pkkgl
aUlqZckuJ8I2Yo6zlTLX97XpaXEYAWgCHmO4EB36pPi8IkX9xze7I+ynoJ1gTXwk8+cTCcKS0fMW
40SStElPFF6KX2QEi16FiTAqcBzZcO1ss8Ljg+T0O50wMeUg2kAJ4EEssV/XwIfr5BFszhlaLZqm
2AUMMhX4wUmMP/1P3X8YMchdz5r53DskH6cN/oaNYavmGVZo5E7jyxYAXidJRAkZ7eXdbcutsYBK
TD3Ww+vBVXvK6ukqtB0j3fQfl6AjLpk1T+xPAO+qV1LihTLb1/0K/aG549a7IATW16sPcIyPVaSe
oESHjIHceIm8zb/u40fFiLxGMCuZiJKOnjHYEbqBfJMAieoaFKaCBo1tV7c35lQCIzM8ETJ7MgzD
2nPBrE5bKCFlI/6c2uOJGvQRzASaW6zIYPp6QQtW4m7LaBP+1YyQ/BwpqX6DjRSiBva4502buJkc
PKNiex3vGaujAZdlj5Sa7/dNUsdD8xIWGsuRo/4ARLxWSREInmuxp0u6g7RoHWDkkKfvhyrp+Nfv
R9a0T8OcbnfXhsfhSdlsVWPZeBUkM4YPBukiITTQ/ZuIpWD3f/pYoWGZX5zJo87C9xXyY8FNDWEw
JwrnmAsGEVpI0h/ZyDJUk+FLLP0lPDzHASw9NiF/bQhf+j24PGUCUPWFvOq2eq0Jd50WUFUCbfTN
Ivtyer2NHVVMP5OGfT0DMD/2GP14t8fCTVinpxL3mbQ5GtnVI2UNiU+FRFOIOW8TqHB4tDpAafK4
b4TNs/sI7IbglGD1D8+DTOHFXuNUtXFizKvaTxqtjBzY4uOJHG4xvYGtGg+lZLV3bj5zBbgXuszs
gfR5bQ8/kklbhzHkqgr0xcAJx1fOJd8X0eFjvOVvvZepS/EMQYWkRGIu6tiv5qhVxmStZZDY2Pyb
MJSDMktbTWpDQhtqPCzkJYlvpY4WNkfXYCvibNghuw8YeTuzPWhiCCCkPxvY6fQaYyF3KAhhkn+H
OMQpfaII+stOxj/ORrK/0AHexFP0nfunuAY9NC+n2nxGgWI23sA1fpCgxw9EW2RGedc9rohrnh9Z
NzbWhLpnPiW98+xMcf2tsKeLtQtt2rO6xmRDPiyMETD49bzIUJ29NiIIl9kjTKnJBdCBJEfaW4do
CCJPqTrf520QKOUj9A5aYb8oUQdTkBVuQUgm5buiWoVrMqUUsZapgh1v4YcUDpF8dJx9L8laOFrj
DGukCP4WEewuP9YNR+ZOlRLRc2LpzGBiBdZDTRBNiqtv9Y628IoLp65xXpW4nHVqoJ3JUB2pdS5n
GKbzj94EIQrdKc1TwTdRYq5LTlS1uC90GrHMKNNgJD2FrmX7M5dq0fqkMFmMmcR4lqRmdpJNmwbs
9ZJ3sFnxwNRCYpwaxr+WM4SKbeAel2IBi250/TJO2By56LUvJcUBm4xN0j208AqtVb920q7CTJnT
DDc3divIbAps2kwrukoAWqEs0CsCahHR9NNRu7LOzvq86bRWhH0wdYoNzOS7qDOvaIhD08LchXGw
LLK0tVOp3Jr1+T75KUjC8ocoeJP8ljp+5EMAl9IE2tVvCUdB501XcVbrDipiebqkQeU5hSVg9cEa
lipUfTfumfigYHBtOe8fSa1m0P1oIl5TVjBQDqi7XUshLZBaUM1fJ33xQlBpFhIsJqSEYKKNHXMT
66qgV4hN2+uXg7uM+HqTb/50PJTP9osxsBpdDeRFeQkDENQzIBIXsx6qheOJobQhhZ7wJQWxF+AD
2sk3dnMaO+YdYt/2xeX5JjaHS+x/VBWjeVIuLvayfxL5PCkQO19XelUM6SN0er0a0cYJe3LY3e7p
A0J0Rbv63nWR5UkxZzCHjZ28vqL8SSnZimIlocOFdaBkxdMk791OGQ8ZLMs6VN0li5C/af1ATi81
a6wMGzzjsCz7l0FVr78CDW6NsCEb3bdBD/olC2132tC6lndpB0VlAHY6mGwXUCQiigPo3HBTpJ3Z
TCerMC6GcuKE/kLovW2a5yybSTeJFgLwRucsIcQVjIIjmjiE8PZM5kbLWD6QoxNUVAKW7SXjTwko
aV/ShXhkBqaAVSpEjyxYkucvy4fA3NgTk2mQjE7aDHy83J+HX4Rq1pcQ9DPCVAmvhV4Z16vQjJJX
fXxsvp3jyD2Ln1+BaZYN7CObmGNZFpvovLwppzdI8mYaV8HU2juJCcjvHh8vyoPdrGFH0/YWVcqW
tYU8q5a72hhOEIylivFNNmVjwC3Jwa3D7f8bhuwlDvOGFLi8b/MMF/YwTvJaaoc11Z3JW6NGa6/u
WTGK+ZbzxZYCvssKsuToKK4FYoMjnTiC3ubZmSIRGB06YsFctlQlOKAgRkONmo0h1GjwnRpsUxuq
Q2d4DtjCDgl6IrTUmHnRqOT4EKHOa2/dyS7OOLoLMUnRyuqNM/2F5xLimEANFnlvjKSzNBqPvUdq
LaOCfWYD4UWLEM+LEzTihBknszlGDCf9HQCIRSKTPZDIomGUk9OMhS6L0U6OGmGGxtYwosgtatjK
rVt7SSrWBXrwtRZWdpfwS0DvGzK/Z7jME49hQq3qZuoa1Fb+nY05jPFNL2rRgnPB9zpFUaaeMz55
UXOW7QYsTgcfqD151qDsL4bXrpw8hgIsNEbfdyye0bWSallrE2PgVN23JuvDw3e/a64Or2O1sMVf
INU/qaQ/g3kIbxtO4OqwpF8zlxyXq4XAi9wsayY4NZRqE03/iddUIpCilQzHk4LnOx2WgtbzJzp6
LHndc5PuBfTwMPD+WtVhSB1iSljjq8kHaLRwDSCJoccwYndUWcfYYi5/8g8yEjJfZx6N/ehBOrAt
12VLVQEQ/DKwPl0rDbmwPFN5u9RnVyKH+9aMcEB74UI+uakK6PmszB42YuOGEOLtQGeDqYpD0Mwk
tgtctk/7UhFPBnT6amisP+SAB39eDfw7fj+NPS/4agUIbk9Nyl9BNzWr7VXJueB3wquOvxZDaZ1d
r4947IW77peacVeFOQ8j8oD9UhWx8o7lci8xpaC/LLqWW89veAjYkm+fU217lQWLAEAg+jFPRpXo
QK7WsTnchOYdDkmcBDPijxMBA+b67XTfY9pev31Qu+reNrjYugSbI3ot/iwh2IiWeJQzdZyiywWE
8JCBP8fjylampZ7+huE21W4j+soanVmB/urQvZRk3Hq3QNx37VKa8SKA41yU81ZLDdiSgFgQk3sG
gnuvTovp7FLXUhtioF/9q45cMQPV1s0fafNIMkXNOppo68MWcbrL5Y6XeKI5CyYOHF9P2V3CZJGk
j7fz0ZcW4rIHxXkyb3+BVu0rX+1V3HH/p0dmrNuWzT3CNl0aLkvi98r3VYGZceYvm/aOiAO9KTgW
/bUsZ3MEMtzYjw4YBVidEJcWaOvFMoUYqdQ07TfsOa6NWLxjOiArQMsflS+53N2vQA2BjQUlZz9W
GxrzeK+F2zkgit8QzDgTKOT/Hb7jn6T4RWG4iR1kR0mTsFRlJSlUBNFdrLndseYYdabmHUi1BDrz
syQ1mZXKuxEEG6KrZfRB9s9EUoyqpgNQu1Fidy99dcPiNbn/0O525ExX4ZhBzFzyo037MbCrvTSh
xPbRuely+AsrXd6csgsPbrdezuvwwPCD9wFCLOOEELLFN2JDzwvIvUU9UxjZpDAuvhZkadm2bujx
jcsW0q/9BFP26zJ1OKlUve+c4co/BYzyfLor5CVP+AHqJkE+YK3Q1GsBu7n58ky8o+1h1zLRNurD
WEgP9wDCtgr5t/aDK/Ywh7ZClZcWkgyFLjV1zEM9+tToWgz2g1QQtU+s3+tzRbmIzkL2maRP8S+2
1aClg+3Mify91ofpiFLAhIPeRkxpIV2e9A2vcl/o/Qpgcvt4yXakMG+77BMB1rMSKxGOiw34Og4Q
06hx/t6Asp1Olfq9juYgXQUHehCRvF7x/KpzU3udX44qmS+whqqboWxoUV9IAHd8geruNgmS18mH
il50p9b2n4b76WAmNaKBFB/rQ/G9sobO9CZcFlsfzI/CygcUnbn/oX7baxrDqGeB+a8E/5LWidQi
J/42aKhUGBmcsqzBigyeK6Z/d021yVmqdLjq32cBQI2BG14vt4AWaPIAiZYagJGQw7kTt9tnb+UV
R+ZYfqS6hSXvSPmzZEZOv5abIi/T1UCHHAdO7VBm9pC9cAnS6cpYoDkjT/6AtnVyEpgWBr8KxaSb
KghUNsi90byjGCvKSbttzqTLaQbbpQKWbD/cwgO/Vja4yhL5137+1aTjkNaUb11edmWrdkuCRZiP
OyYB9CVzsnHIlyFupre+H2+2DQq/w6zF/iElc0iWYz7SWSj+z6kglnkIgpOvsUZ2qt3v25P0SlYN
7L/H0puz7Asm6rpiSSYTqEMzOuAa+oUxGQYm+04MYNnH81jRA1mwk29Ub1k1DOS2XXnehkro2ZrF
FCKCQLWXkQiFzLKgnwBuXDTfFAcW17lnSe4EtAAV3fO4ebu2PUg81kt4EYfkA/61zxMWiMcArlU3
kgKNC+5vu8XZqOoBlnjgFf8VLO4mypSmaLN7KI6YDDoLaoegkmZVHczcnNto3eWyvWc0xGLxTE6y
m32IvtPcDMpMIO+rS5Hzgy6zPrHomKEotY8uSH0g7iS9HxpSw/6nCI00z56czO+Oo2YEnWkdJ3Z4
PVjulHN7XsPXZWY1BuxmGD5y//SyrIHktY3B2Dl+/v34sz/Zf9AXUVbLjGZEAuRkSUCMvIWiuyZS
GFXW9DluJUg3JOEvR2RbQSGTL0mr6r05zdWHFeml39mACuDHcsE/hcXvE3a+YCRqxP2PTlk+VjZx
D8EB4BnGitPvgX2EpZ4Eq2dUz2OeyawR9DxNyQGdzQKmoFytJb7i4WKTGNB1ks+Kyj7g858gkRqv
ZnZGOTUCmsiwdZElznN/mQdjlN3+V+SjLWggO6DFMq34N1BB7KjkBiAR44z7CPjSwNfTk0LuxsqQ
pKrHP2egD+ooQkm9J10l08qr9FHBynG8cz0cmNdfre1ZngEIAL/FjE3R83mU326ROjZEOIeaEuC7
oXO/JCBHBWr0y8E+UWhoIypzpsAN/fErH/cfvsw+fho/lcg5FvNrDvA1bsAx6Xr5GPYTDeuQ3RmK
/cn159FuABulYJ51Eq2p3sAXdURRF2vvBNHjpL4v+xcIl1ua9sswVKfOBMIW5VRuOjRvVHa6x2jw
W5eMetiNkLUBIaDzVFm/GtqZdFI/n37uDL2It0seI8C4g2A/O/5UGDohCL+spNGuxuGN7OFPxS0V
0WAYiCxOda3QAgLliUq+v+DjCb3aw/EVSPRn50lQWl9SL5jB2xc2YS2vUwEd28P3IbytZqEW45XI
WN3TyWSJFAqHa/toYPXG61kF/JBSqsJVmFO35BE16JtYF9Y48W0SRZuyH1xCGELmZN/87Pyk4lS7
ZH7/8YTB7UG+lQJGJXP+hQGQsXwUvYTanDaZ7uJ2xgcNMfgtt2JJxsaWrxYrP5D7UmkvL0Iq5vsM
gjDzTFMd4nys+SzDZoi7uthjSqB9DWExMDgRn1AtL6+ouNiO01XOtfOPRof6kcEeCHDnzTqCmx6F
ChCy8z128ii7ZrgPnE7v6VXmhFr7FVRQk2UUaXAOPh84+hiGU/WQYoDPplTq30HwkfFVmnIMwPpX
3tUmZnUJKxG8f0yEJFAa/iqi8YuPmGqBoSPzzx6P+gU/8SWJlEA/3VuHVXfLwUZ+3j3t9d2sUSGx
3Oky/mb9UrCnSlzElgQA3Lco/uXyKXeaoeU40E4R/8Jl7v7xnu6JWWZpR78h4XPrcwmI9a+qWdRP
5cRskYY3WMmyAsxtiBww8DqLjvw12fGPDurikCDqnvcamJU7a7DMJI5ggF9UEUjmzhSq6Yp8/ge9
Noai/9nPfqntNl0ZdRfgl6DUDCZjXLrnDYO/j31atnkrKTq0eDPqMCe14B4Hq/fFbHbsWpDXtLco
k932gR9qzkucjsEWN1LWdAlUin0NLTWavnajTF4adw6+KKqNOvYGKMeVL33W/sCoVv1lvURFPRIq
X0gouZeFeWuqBfTWJ5P84ErUvMQ10Ci1ArGchG3cappwy/UvcC9puByc50k7QKPISR2x3IlNxTz0
e/LAVY3jXQy2UMVUUqiHWtNZJwkqdJFq4FbyIxx5ZROi1mYtVJOVBVI7JafKchZN4L4bzW0lEQem
N3TN+0sWhDu7+IlFmAPIN343OtMg1aAmZifYuit9r1vM/BJIWFe1kUOJvZpa8ri00elB4vRRflpH
pcLEj3GsOCC4j2ffOMd/R3ckFzMSU2NUaOe7iwnI/uxN9UpSRwkJcCRjIv7Mbx7pudCKfUsEfFTZ
lp3I1/tm6OWK3mC3qSHsSQnwKzud8maTwxGRWAE5R+STW1ol0DVvZ+D4CmAWtJOMQBchMoEahOoI
b902FHiRpo+NsVsGmxXd5R7Ume3pc9EHa10MywO9WrltEroQLkHAVhjBIq0OrF6fYp7KSp4eGEFL
7qucr56gsUZfUYCD4B/fAuHaAaMnSMSfVHU0pdoNx3VW8phLbtN45KH5dWbAr8wHhw10CxFM6bml
l8MTCeoGDehsm9AaBfPYd9NpxfzQOo6neqYUVoDO+7B36fBa2S3+D2j3JJ3D7l9u69jh8XuQmTMH
LZUoz8GEC/LLk4kNBLB+ZoS6FdashgFDciN3nea/iOZiKADqpI78Aq+H1fsRjO0X+taYPPjwDKx0
KX+ragCmVXGvwMfFqd6eSJEgrHC3+eIbQAgt6q2KgA2ReImX4InUDU06mbLwNmYVq0x3uK0DUv+x
7ctmLaUpf+HcOKEOzDK9llwDXnlfqUh7ytSJhGMHqSwN/Kd7uvDVHuBQ3B9PAPX3HtjuH3gUInag
I6BB5CX0F/KjSQF3ijdYrsqDxSRUUncX8bf4chcQR8GqSa4XrlD7oGO1KaIR6s6mRS1v/3j0d/+i
k+ME5+IoHLkDmHC1SSEmTDouuP6EiGbuOkfVj+9XzElU+HskFdxTV+ge/Wl6pdbQrSEFUcCgAL8U
TR9VYW/7xJC9zn2MJDsiYlHCsj1hgDezaf33td0aXNY7EvslK7/6x0foDCUw5cWo93Tjvane3TXY
APls++fliqc56L1Uocwey8DsLFaTImTBD2/H4PNEBKEeWWnQt9x/H5YBK8oWWCEBgP7UGdnMG6MH
irLlOeayP8jMPRn1FYoN1UvQb4+RZ1/DtSBm64ffgtallYxRNrDRVvmYBxQO88f9yDz16FW/Rh7x
HMptZxRtP02ZW7TG/00EInGu+oW0hXPMI4CprqAxtwsDnP5UgZv6moaCt+Fu1i8edoK42MSK4i/R
pOQuJ3mic/KUk5vOIj1JyRo3HRBu+3pD8TqyzywL5jfhBIiDbE3NYvf6SLNZiEucgUN3ThJy38X0
eKbdJf9SkucRnSVnN4MfUUEs8OQxA5dEHZks3GWRPpkA0LBK33LRpHvDSADXERjdIx/IdMArh2ww
0ZC9ezkd6OrJcUuRy5zBOfPlolTrfiEkq8/aFkl5S4iDrUR2WjbT6BeElXZq7e7P3sQY1eE1Ymy7
uVCwFsqWXNqYg3Z/Q8u55SCysR4370ozpQgHeJEa2Yy5G7FZd/p4BJPITUJlXjhIOjfJh4fIXmuD
IRTWQCU8QffkX400A3+oQq/7PK7sV1WY7fkihWyyms2Cb9JvwbGZ+Ilv4nc72xEeJGx1NjFYBXgL
pqPoGLkGotgRxZ8Z10RZ1IrFEA1YW6KBRDsu1/F9h/D37t6OuOm6nGUNpI2n4GwP7LeWzw6tBPHT
/AfO+bWXsxyDPpHTqXQ6DUNqKntvuFqYk3QZGk/f37o4rD2ANZ9ITCaAgoTwiIX8ps7CAWUCbunJ
Cf5CbsReZTBua5UP1L9daqizIsvMSn0HIKEwl0ILqEu87gwyfJ5S3DsVnwAMgLqDpVamUoQU60va
Oqb/7EYG/PpxRtK/IVXsKSymw1WRMs5fhCTS/dVkQ1LyvG5D/yUaQ4W2h3QJgepJT7rmQY153+jC
eKgw0BnFaEt026wG3WJI+eZGNnSTFl9SeQhWPeMBHp085bGvPiu3RlabbdHO3A7e/N9r6wOh+KnJ
3pFnBx0k11x3PwRAGQ5dHum4tQzuHfrKyEANWraqMgw/gAhHpXuOQd1W/ZaHsKBSQLsDhYYo24X0
Ql+6uiB38o0JZ60CYwaQb2gaKZLKT4ORTig75nd7uwhBPpQWJlQtrR/WbIePtY6s0L0dl0t9WNVP
YvMkWWEWwJJ7nV/ndfRC1K8bsroMmkEUAvnco17txlJGTESjlG6i8vuRGc7rd+0D9x0jhOG5+etu
Gu7IU9IvZE+QBtqzvU9XPh8Mwy6sPY3MwXQXR/U7UwlQBJQCN722EZ8DgkX1THkloqpfALdt7s6j
jSVVMJkN2fhFwXKRCsoZ5mmt/j7/A/KqrLi2Y0olYMmX+lV9gQIfpi4LdaSovpHrII77eE9W5BSO
cqzA2n/bwCupphsbSwruJvkoakrf9Y578/5tTFJeZjZnqV6XQtMIM/DDkAuA31fEDFYOfBaDYt9T
iGhDpyDEaYRWqSW5KskAnarNefGjpRQ5MwlqVSSEas9NkppQWTUVFtiy4u39yxmLB6SETJ5eP/dH
ECOOhSAnhnQz86Ibw+l3ZOPPRdrIkEtus8t+ZBQugdTTruKqzSDq3+urvwhknspw0Zl2DziXkyLO
GGeqg1qhuSAYVGsEEojUoYU92T0B80i90EaA5TC6rCcaEgZnGxPrzWMZgg4/YOsMOKuZxL1WI9+U
/HINTiJCOuC7X1pzEbW//1e6RiGc+nQgCssNL0T6drULGWIswZXIwQssZgkkU2+VsU8LHhphrce+
Zm3ryUHXPhMFs/qC6ISZghVP04z4X80dz8X9E7/xiF2oV/khF9Gg1jU+ifKM4uFwtkUAWoK8rZkH
yYpFcMHOsTllhK72ngdeahlHn6bRrxWuqBq2ifEvgt1u8NATswPsDavOkZCE2mf1SxiTWCUzEnzY
vExMpMZvmguAQSXVzmGpu+DymQzwjpDAX0WFnDBAEdeoAQcvZf4kQhrai/tTscIK9feR/1umR8q2
NmTHEREfT/e+CslkU/9uqMQaLRbgZ6ts6BHzPjrbM/kNJiGkZE0GvqU/uEiAE1IQdMXLjBE3lYqO
7QeukXtpgn4yoDIQVL+nX9h4fM6w1HuVwAhkqtxjWXOLo2C2rj57wDxsU5kIIxRp8aYVV+yxh2+S
iG75Lvpsny23KdqV885MRYEQ91fCY4zIbiVJv7VnRgWJb3nJoh094zWRamdvJzUvhta1PrTRMTfu
uOuB0rkzxJ8ctj7TzKXDIagB/1HSsh1B03y3hL8q8aibzyADOnI1Otzrj3gYLHbmkk3DhDGxPKHO
JulPQx6w9OrlmeTnBQ8hzFbO107mCgaP7kUmEr6BaF/61NfVN9qejWQfpjjnAAAAUHviQmZaCHJ+
n8CEaDH2ar1JBr+vc1Xf95jtONYwozpCO/JBgrgL/UPeHCQktYJrNXthquLCu7Mj3MibuG6J4jZ6
EqAB+xKkSv1xWcjBU1l1bxoq1VxvZhZcJPiqKpModEebiUOxwQ+lw2Ic9jdBNaYt955z7bo7e14L
JfvcLAdmrah7k/MXrse4c0Hjtt4xZqvNKtRaenFGQB0nsVs9NtE+DPlr3QJF/JtqrRnN4uU21F0m
S5Irs+B8+K/J6FQ2LTq0sjuYnHeUrJ9OaVqMNwOZ30S4x+kOm8VfHwyJwQ1vG+uDNCD/EfAYn6lE
m7TALMVgCe+qzuvjgNCag8hzhmQs4ARjwRurbrg4K8ygxb04CQkcOIRmFJF29x6gIKXMVD0RR7CS
H8uJGTlfgxmDCIfFDB21RK9YvKgAaVzxTNBsY6v/v3/6OL+rNfUKo7JBI38sl5Rjf8J6FhttlYvr
Zb+FrLGaVSoPmzC8DsawBCqiMhwpUpnGPzpGjBE58Bp557y3pEhGdLpZSYpEawXV0lHKlcztbewC
P3Ay1Y7Zn2Etfd9U/+Zj0IgxZw218qxUNVQobUO4yA2eMwFlCZ6VBtEd50wvwLf0b4N7ESIBDvSQ
cWBgMadk+mZjQ++JZ2ooTBrqroHWyY7j+qsRp8vo/SPoQ6LPo6To0jpNaM44CZCcduMwVeeu8F5G
xs3ZiBAFvvUbVUq55hgxJUPLj+y784yzZDZHklR7T7KTrwxBXS8ZVFQSpBcAxlRPM0sgL41onajQ
/jAU9a5v27HHcOZ1bZqzgDtMf/mLh1sMRASsCYWOkCG98TMaoqmJMOu8XLDCl/Qc7MSL8MX9JDj8
62KPcjbi2R1JMStCsB6cRix8v6rYn++rYTmSPE+oUWgwm2xSgPHYDi5ZKOdQ0PnioVWsdymzFPZS
5+CkF2EkSFnvEM0snwdIq/CxfrLcf8dJRROQQXov5UGcebjsth1QqdGFlmEuYbviZGF8N09pEE7u
f817r7OXiObfEgk4knuljhmbGJVE4dwJZMm1hXB/EDxrcAnjjtq6S7abg0c/yOAdOQ6IjfIrLNn2
MD22rQ404URvkwygHa1jlj6bYJj4arG4pR6sqAgJGDjSGVDrzusMoMl3Sa6cB/nr4CgfGXKwtNF2
BRJvDyMiUjKkmubowIrrCff33AzJpqsM8OjCaEhiSM2XajKznpj3n4r1nq9DY4NclAPdqos1HkGa
pVsJZKlK/LXyJ3yantbumzXNrSVaijjJ9LD4weIJKh9zcBgZ0fV/dH/9UWdSCFOJeUZwM3IgxXZ2
nE5n2pHsL7ExuNQbf3TVbG8B53cKKnwIRq7zUFhZ86WSykDfJvn5mGVKdIR3IutnZFsjJ1CVDTtp
WeQ6BqHF/8lMqyelp5HlRZoX/+S3k9Me/03VJwqu6x1opUWOfPm1KTQqO9gIYGPLk/bNj9O4diXk
bS7v8y47ovD4bzfMP8dEThNCLq2QGdEXs6FXn3wWA5GMP8vZdM9et/KTUTfGoPaAA73P/f/Ys3B0
7uVT4q5TN/2NhCxhOL/0tDKTZMsQOaX636AdAOrfnfeDR5ZFVLZ2KYlaNusEhBVIaPmsRpgWsta6
RBaOWB0+BO6QD25zV5MinHEVinfLhbcMo3Vra13A8sDdMI+V0uq76W+Cp08pGMGaGpQBbC4CKWEN
sLtw8xwMSLDc3xeN+hAxjngtSTpjsjecW33NlMOx0PiJ5128sQNc2F0VCsnDe8gwk13uvpeql36q
E3QE5XS1Ez4c0xcp88NkE2Y8sdcx+tJJi4n3Yq7vz9LZBlCBBA/sGBwBr5qB+6FZ54gbrbpPw6HW
YenyUAAdLSCs2UYt1XidyXfRYSQsBW1VzD8Oms+h/5HePmBzHrRk/ZudFkO0Ztv4kRug2kaZmJZK
EKHT0X9HaB3yfv6fjAwC6O28z8eMrFPwtwFB8n6A3+jkEF1+w5k4PaAqUpsbWbOhkDNKolUTLnZ9
YALkaJVq4D7BNqMT2NWYIfuA/z1p5J5ZfueGttuAu36k44UTyzw+WcxgJTsT8wrTQJAXfIGD341/
IA2IAcv4ytKE8tCaqGvlF3YFMgsO3SHH239duqkcc9P032q44jebataCTvhNmRFhGE0F7T8xYDCu
YCUo+rfjPWz2Xj5Vz44Vk9ef5wkpr47qd6d6hjiD8jlU41kYfCbXmOpuRlFVQ+Yh29JvQMQjhyCj
IH3Gub0nHmMFHEDwOheba5TR7HQRJbQvVTXgrldLcjveCt1g1dCapqMpLDpBdnMZqOeop9K4ooSe
2mKn1eHybJsXfxuF3vIyxjSe+cnPVHjee1d5SwIjUsx+T4QisPjGAM9b2G96LR8F+/RkS4sYR3zB
fq9hGnSF0AmfBq4zRk7cZOCqZI4V8U5fQLIK+2AsQ9Cic9lvHKcHg1/NeVmlb58rcgGm6VMfWvRb
GEIuhrB4rIVa2ALRm6z52NZZx6xiIA7pYaw0o7JwB9Lubg+q5hHasVkMGbGt5nYjh50nZrdfhV0m
yFCFkRXVf+r6vyW86bxYFvGrKcOolzUUjPxW35U5dD0iP7AP4A4G3lJFT725nVwDY9KkHYPVBpt7
zICtb9i0n5Wct1G+9ZSu/54bDx6in1t0mYguD2ot4tYW371Dy9eeedTE54HhFVXf1ZIg/66VOchM
mK87E2FITKrlV0yMe1oZkCsuIu1EFAsV5kOxcsEfV+MPUWkx7ZskxkSDrFoyOGzAuZFY47LFY5Ph
DrY66t5oDOz/PS9hCzTMQuyS2s06q+7fbwiU0XxR6zV++vuWMP3z4ToKuwOOluSy8f4S185/ywXR
AhS9KIJPXjSb/uyE4tywuuEd+nWgNuBJnR6gvNJrMBiolbGaIr509V6pmY8e0r8LZVeckPgT3tS/
qX+edAybwdgvXtrS1sQfrKgyPf0VrYORFoo0ELIg/UjbNvUa/+lisU49VoSdyPQXOyqtZgUbtOmu
OYXMLMtcHK2P9AkTBpUosKBvuEY1CY9LOeh2D0JKpB0jpFiG1o168RHaQ3LBz6aOLQbqfOTvl2jj
vBWnmHxzuyFvwbwxLlUzPbivOs3MSR7a+qR+nCusjfudL3wLYiGoGfPOyLTeEvjVJS6ADD551PtI
WrNkC+ZImJsIJu5lhV7/2irM01l4IVgOzWt26atU4ZHVEmCD1ClpLih59RiZVU0SmYbBfVtZgtOV
2mmKlMgfHmQtH+RkFnxze6U4TwBYk60oOGQXwZgr82XcUpgBk3lO7e+wYK35FdgqeGJO812+EAny
a3pSQ3zlddMVPICkvMituY5dk3I5eGbnm+naThLNIIrPCHuITkA7/GvFFSAxedJKexUv+eZcpEY8
jYPvbfU+cHWW5OtUE7PP6D/aAOKVvAxEUQtu05d7wSW0DDq8Em34fiUfy1jk/sAIhAPPI6KGLavq
vJmDdpwYFCPCvB6DJagJje+GWfhzn5ykRmny/pGTx+FKFPkorONP+n6R9J6afcO2OAClycvlFnlv
zPCrQd3OVZo9SAbh8Ou2R6jMMu+S/TMvVdSgCxu0+RicP//uL/D/H24oeh9K+W65dGhuDX6DGGuN
KaUK0Oxt5BY24k15pq0mC3K5CJ6JfmysepjhpOBs95ZnfWHscYxF+abY3YtuyqQtCbjfWURlOCLR
89u6OzAABy7Jmi1hX0XeHDOsALWQaXlCSUM0osdVMAKgAPOXFcFYD8netCE6L819HUTghQ3K4aXT
fMwetDVpbgqR5GUxB9Y7WmSox6lo5xUOP9fioj5THhAZFYE55qFPEDLNSd6yj077amAvSzI0e8Dn
UmGfV5cQhhuTISXZPDGXq6h70706R40ZSICqskv07okH36gRVnTG//1KxLsVm7Law15hKSDMyzEL
kyTwLA128teeKQY6DRpQ/3UN6Wd3D2QCyyOIdaa5UZQ2bOVGXoFTjm4ShUlnz2ENa58JGT5MYf6Y
humHbN7dNHK4OIe0m/g9WbOsuJlBhzFkTfYtu55Q02r1HijUdRC7pcr7j9+lYvC8/T7EgBzvh4Rl
wxpkCReQDCR8BG2OJ6BMw4y997iF9SzchgnErnQO71hjSC7owohRUmh1TsQnb74CNi+xscKCuZqF
mgxtM1FiUJ4xYQvhgcuF9NLwOR67Lh823f0UXLebRzowm6rTeeWp0QO3VWPpzZQQ9abdRBETcDwe
8Or6ECeYmEWd0f9Pyc55MWYWNN2y/evQJcKdtFY9WbXdWf59URANxzui/NgRDkXbeRVQCbDbHlTn
CYl8IcSnnV2oJg3Lm7s+uFH6eL5SaDLJMU6d2bq8Y7DGKTQqES57JdBO5gA/2hhqBGG2F5JiddKD
LbdKRByGTeHyx6Ye/6MEuHvHK7piP5id5Kfto0r55W/ZrASvEy55fwnKbIerPE2NL7H7Kw+DfGmw
sElQcpQXw6ryaN7iMoxiE5nCLozJvjssd/YIVkBdNpMtrPfbY23ouliAcjLmBi6p6zMZwpUypZXT
tpnMh1rASZJnFE4DCH3aCnF72x2pPz2EwssFzDqKFbjaMTvo97vRYM1Gy2a9GfMjhCvbruNAHqz4
ZejeMc1IQwJTRVQ2oHVcbzsFF4EiQGlG6Ws4vxY/mDX94+fuwwHXUggJrP4zhM/M3LxYxFZKuAsk
MayGm6UVjgwmTxzgqUw6k2NfcnCa+EFBfNs2q4sz4EwcnyUTY7aM7PhoRcJPs1UXKxJcF+Cd27hK
F+KAc4ZfMJuvVk0R5cyFexOV3AyECmmUp3/xmeQxwiunvxd4BjKhu4YOsz84B1+8N4Uj7TEmin5K
9sI56zU7Dij5+mEpOYCUcJoryA7jwdnY6w076P+Zj6+1NP/sL79S1zbRyjLyL78Ie2bqVY1V5pMF
MHdOoFmGwAJM6+XHbVp+fiEyiRSUPsYko8YOSQWuKRfUwuwGawzi6N7kkPk0YBoRjOB9K36MSf1D
GUOdi7+Z+8GsBSBUL3IesBOpaICwUTyQJBFf2dlziEyFyoPiagB6OuwcgpxueB1z5LbvI+H68OVV
rgh5hcUDsZmgB+9S6KdnUBrjN89rnd0+S1p1XWDDxO4AsINcbklNZoB9YWeqJuVCzuRbcOO3akWP
I5kyLECrIT8R4G9IijqbdkPdS6bASLXSlWDbiLFta08D8cDwfKbL61mqxc0vjAXy8JluoRxGlLkV
Ucx7mOjvvqcO2T/ygxVLAF+ouD+mWq1qfx7i2DV6awXKyMbm0HP9b64bmyq+hX7u6yyxq7GUsVMx
x2yw1Yal+eDsrM6vd5J3OkSnFhL8iMfKcbTgza61G+GRwhOoFBi6ljUHpaRjlQbu1mn91SI45lrd
XVn8RlahcL8jvRycMITVIVGdmepRZKPNLzaumQrmJojv+EMVtinz5lnPRX6IqLH/4ohdda+0DeYA
p7tPcaYpY+lIgvxPOwJmirxz27+RM0bO4+pxPzC3cMBBl93wd7CQJyVbv19XiofO783zHcjLYgg4
BnUdGOIvHmOeCEUyROct0O/UnjxxXfRoJfAR9x92PbMFAHHJp3f9U52btxtGoJm7KiTyRlo6kBDL
Stlnsx5T5smsBlMnY65J6Md6j6pSiOsj36uAlPY/nQ6XUmoVtXpp7gLT0ks/G9Vp+b9cH0QtZelN
LPu2g+zsI5WF4d2t4Gt/JIwxh30pofJb4b2L48t2VWVx7t95wMIMORI2DZI1h8koQifvTC2eWydq
qU+5Hsi2WhhLvk0kfmuKR6wPvY5Kvj7eyeulLUfe3it5opRM1iPhm+1LRggiL/NCcYd9bgf/6diY
R9rnmGIqvob65hudcgBd9omZQP+IaSfWW1EbeJZoRSUUyybXQ6X3NsB/Blm/JlFJdKj+jpHXQXjJ
SmDoPdhxUMfa7RsttdMIgyX0A+UumvC5l+qeQtg1Q7s4XYfaqjSk12sSs3zLCheYKaEEGg4pH2NH
19O3gtGh7I2Eq6PAyU8yAKnjNkT0aEQHPPbZGYT2ZO53od6KOA5FvuCypCPUFUOaJQsS8+x+InHC
TipmtvZSX/Wjr61XYk15nJmkZ57qn4KlxgePp5WXtjjLQaJSFC92oyXDE49nSITs+qqmO1iCY2xe
O51JZf+Uy0UvtPR69g51uQyZ4gn5A0miYCVc3T40cElKoqJawo1xnIWuoBmTkgT7sGj5UDIRpXZX
GKB6oQ2dwaunk2CkhWCeuMoJdGevxC09GaqeSVpPGkfy+gNwkPARubRXEElZwrPG/rkRYf1iNgAX
+XVBZkwFESP6Lystix2DbFauwpiTE0tElD87aNvYobnP1G9x2DddmHUkfraGJtepp5yEVPr8DpJP
OhYMQUg0p5K5v4lUqZ4kamGSXKJApX5GfqK+o/st79jW0NOZbObkk7NBv50+MyEGNJ1K64Gpjrt8
xNDyIEpYXBgn4N4XVV0f4zUIClGxUMI5kdAPVl4JsMhPcqfURJug3KnVG0fXEV/LnfpRvbJFcf8g
5j1NJIZLtGcGSBYoYJlv4MefevNkWB9DYTWbM8kH761FY/M+Q8TBxR1pDDvnFmXHeqy1uZmlc3QT
lo8WwkVV1frAuDSMu1qsirITizrupJi2QPtYnFGFakCmD2mQ6oWL0mPa8HQUELvGm0QvfU2Fa9jU
EK66bWtVGKmhG+J1JqdWYM4ua9z+/XtgU/rCKd+Taobkk+tqYhAK8wpPIdCyxT/0YgnkIVnnondw
njWwlzMXJXCMVJIjJXdLwdxDLH7QHb27NP/CMbzY0vnHyAkTt/vAjBO5xqjGtr/Ihdr/eB50Lh40
DhwLhCaW/dZM2uN1svGp2dkH0BwhuK7pZu3i0Yb10tvk6+yePHMfQkgyHu38HRt2bqr1uf4wZpTJ
wR6Kff1cJTyr3oUdckgy4t+HCNGwq8pJOopPY2ldvUovgGLNttWukj1gvz9x6ghREJ9sjm3BaAL4
kvuYGOK+0DgU2pgNHMR2ObMfQ4G8WbqjoAbJKc/8BD4l+b0GPd1cI3PhEXloOLQkEZtZOozYPOLZ
Hw1BL3af57a6L+z6bWEm+2rLO+lTepgvXoccrQeq3vLHl+ovj+gc86g89pMtW4Ldxh66JrZrjBcU
tg0Az50mPmS4wwiEV58pWn/EBTi6LHCdtBN2NqAgPITPWgeKAAlER7zB5hiHxbKvuOt306JtM73f
o9R1HYom6bimV+fLaHl47qxdplZWZfnw09IK+3OUfHnEczDgZvyojheXvwf0YBRTEcdxFiqofJnB
lysV74fKOJacPWxiv6vOoJO72lUmPVcPAkntexh4cayd68gAkzZOhe0hmHhbSFo3jSewPPb1ap6E
KWWmKBkyjGqbH3JIQIWcmz6C2YLDW/NWibzK3nbeMWzEtIIzRUPxogLa4xiBbYf5zdfTMJKXtCXu
Moj+bfubTgEvHw6Yr54A+VzbG0uHfkKiSk5O8zTC2MqSHiUj3r60Nq51yCD3LggYNiAynd5zNehw
D+wmSIbQr4iCyiGNPMNv7pUVFLigwv0DRL+i+23Ovind2S7Ql/WiX2XOybx+n26uiF4uDFzLqGw3
0qhc+ScoEs/+3DHIU9T+/cvEeWR5DrgjzIho9zZ3Khu3AXgkBnWfI2g9hC3EFKpUBlnY7ehepurw
Qf/9Dvz0vCuLG57amDyLBhNDAllSbhGDmWuYLHqF8f6uErLQ3daAD74YmIeCeNyoqIhg7UTgpY0c
uC34KEZkAPvjHUCIJZmu6Rz3miE24AQd3bCIHWUd9UrsRYMLB7+bgwiaaeZ4sVIXQWMPuXH3wLr5
yTjVbN/KZ/slS0NsrHaWwX4jeXnwJ2a3kWSSXm5IMED3JqnD4B/t16S2WSTkZAlg25OOxouQlKSc
uqQMFzEZCzGSdDtJ2K0l7YvYfFSqOr3Srz0sIS+4wAplqMvsq/0zjmQkfaQe9vfe9Jw75UWOC3x7
EgG4YArlhdWTFOA+sXAm+TwTd+rcI33QYd7Rcw1QFQ2GKHT1W4MeOOvHuD771PNvJjLih+odiI9R
/xaDwDoIVO821b2ghMTXlZEvQEq2muwKrAv13ODSkmC2g/a9b5IaXOjqgREKjawkyD5acstpm1Nk
IRHjJaJy7dsE1YUai27DyQ+BFwLKk9m9YpmTwYdgVdFVSfE3E/08mEr+LFjB+xxc+KnhoCqNyNfo
wd8ujiwa6WarhbjywX80HU6Db87a4P+KxZxOF2wmuRr/08O59T5+NBZefQ+eGYxWEwP0cBzs7m+Y
nISDs0E3PHamMy0qoThqowXcP5HznF6ihf50n9BzawWAEfXCj0V/se8qPt3FQmlEKl/GLHtStXlp
wBVXbCLa2XOSIKAkZSEtteETPSL9UPBQMLT0gw+GA5Kn8zsvW3431wNSV4pR70CJtGax25ipHeFP
MtwaB35rU50YZz91H1SruvzmHoqXIwK992W6Agql7eTVmri1EnniM0V2uQWSq7OHs+lb2x4FQLbT
PzPy2NMO/dx4P3zFQbCL8jftwGLGwZsdhrkywVc5EJVFWWKAAYiHtXH4l6tjFJVEy0DXLrJPUUyo
J4rRO8on+z/vSk8reOfo8cgT+kzcknD6pb40VEkBZw0HfFFTcY+ntUn9t71PvtwOurTiX4sOUJRN
Oc7MQ1F45Byp7gehoMZTJMtHQNbbNW4iPbNKxMe5e55fGNVVvD3CSPJa886Og+snVZ3Au8xcwDS+
RkvTmULc/3S0J/VxCKF+gOVp5rz3v+CTu8JbAVWYH5IRJgEXtUSXlYKGVCoqxcGEkYb8cgqc5scw
veR/TA2NlZ31jJvJOFYKzbKCU7Q7XnIn0IPJysUYJxCvFiTEG3nogDdCjnUfuaVt9ig/dpiXrHF7
IP+lD40oSDjAxxDslwzIy385gRsCmGlg2ksOPqFHPkQXV3cKNpb4ie05OPyJ3ocRVrMk1iZFXwy8
79zF0RG5bny2GUO1Kv6u+CIuuyLAvQU4gTWp2RtrjDBechlkOptH00JX66O+7Curm+gmKg4jkJkN
udJcPAzbxpoq0phcKy6TUmRX9dalPqZB360+ZLNSY1wMylGE8OIvyNbRdYZ7j59aIYjeC1ihGdjk
qo6CcXzsZN35909iiOG693KD9RdUNaprZiwE0yt5+2f/y+nO7yJIHlOEXyn4q/vtvXJdFUDCGupf
eY7BXYd5TQLc3ZWh/kgWyJo2UpVw9HkhRIkQCk2YWDzxv4tDmq3oMPaXsSSPQ+RVwOQCkN3uCfoH
+2oeTRYqh4A3CJmagmSrPW2WhEjZcgWdny9j3g8kooqu9A42Ur6z0PQpAy6BPrOiPMSStJddB26K
is4npsgPntOd3TFK6jkGGBMeY1Rh9YXhkXHW09L96jpiPeeAm8xKMvq2sJ34hZkjc0rf0B0xOfN3
hTIPbsUalffReyM76y73MtJtyZz54NaiFLItpR8VWgMcRQ0uqxI/wYqRc1c8BLjsfUjqaM/ubA86
VKaDQPlUjH2CMKl3GhF/UcrIqJ6VAxrg4jgFBvYCj85QKyt/De5Sj+IRk2TMQqGGg0Dtt0aa8fQP
zyUpjoVmyULFWkwAAeM7zwyjF/5FvN9nT16c0hv4grqE7t9CEM96zO2A/+uGAjqKxwB7XQkKxCQ2
P+sW7ARP8NkMRPUjgzVTTz66UtDvF39VUvimUk98NEogF8UlkhmFDzqmiv9+yaH/Fv94q2felDmd
hZCQcKg1QNgGHhmdaoIk3CgkrCI1v/Nt3Dbfj3ib9LQulaoXw/zt70lpS+5WtT6f14rAmQKC9iqX
lyIYEe+NtpGsNDCc9Kxlp7F+VedP7v7I7ooAtdLh5UjbY9HFDonCQE+VIAy+ruB5bUHkhvulyVHD
cYIAaviOeJ7G7njS+BYMGLzd38nNTDxje7wE2yt767uIQsUolDbtblacd0lhjcbGlV8a4CKxL16b
8WzpexZeNL4+RGsr4xxyNNOq8vtYm8hUd9hxwiIjGsZvQRpNnY92E4PuLTKW3ebuuvT7WtlOqRFH
VRMLjVR2kb26fBMkWTdRCLKh1TIX/6kp0sCoy4SMGjRw31ABhudMbqzC+RsVJFyJuw0qqh443yGX
Sk/U9otAu0RQ6MmXzGgnPKcI7u/UUcH5P7zzF8apA9Lm3af+HCKi9GLfrX/yVhx2x13yBNwGkJ1b
IvJYeF2AeaXb1wfMMpcebwA9OuDweMUw8llB2DQXioPo7mr2Al/hRXd0PBdfadQ74ETtud/xcVbi
kNSMCEQSmD/zVrJVY7nHMEmzx6iwoD4aBfkMYfPZI9ubVKNYRp99pzPqLepDeHdVL6TEvytHxzmL
6XTjipuxdeVjEz6m1VlAo78zjhsnN94xljOmjwL7B8sgqbw+0P0jfBUNHdyrq0Ozipr2zCQ5W+SF
NJqi/dema2RB5oaKitMacEkvFOg0pO+135qU2HqlKyY9QL+by/QA/rFTvVXyy00ooWp+YQpx5Eh2
D4GnFFEs8KugOMOVZ4Wc+52SXiM+jyLGtGquwmtQEzuaBqThq+73nLSqbomF1jJuSGA60bsTk41T
rh8hA/4NBrHFMW3yWR19ytdZRqlc991mGCZUwRM1cAtozHYr4CZTrg3GCOLtWpk+tucVcaipYaVa
o8atfQjBKPUK+1LbJObs9K7mITymKm3Pj2UJzGBPDw9N2c6t8MeLIAw/gtGAJaPEDW93vAXfdtOx
Nxt/FPgdziBI4XBlQNmE99ibVwtoutMagigaWWytGResh29VD+KGVLg5N9Qi143X0sIAxsgxXT+4
CrdMQZ5bzGGEFLHjC159CoyLWMF2uq8XRoJ0qDCI/dnSsKcfMZEB3bb8ONV9I75Z6PnA2Y2N37jY
zZFmCjSAUt91sOGk5aE+nPWEz7PClu60WecBKNKnVvgGQgW9Mh3covsnqo82EiuyE95jGluaINru
yGfaP5ypQtlmOgv/pdb0YMfmtMLikKVEKBpF0+PSAaE3TVjjwZjB90nVkphP6uoEDDmeJUVlClai
fP5yv6Hq0WvlqbQMuGIs7nWwJhZw2Gy/kZ0HqkmsZrDSRk82GalQpSuQPlMIHFdBhn3fp2GqkvHS
zHvEuDNnfXOfxX4nyeXTSRvSYifuYUvppZFUvWWsCoVAza+eu1S3Vtp5rGXOJqSc7U5pKwoWSROl
3ZkshsuFepGirAUmZNZx+L3Vrn6Q2a7XGFvj+UQoyiIolgDTwAMftYHIBhDVcZxm+jo/fr1pCOjC
Zm4P+icGTkQ8pCF81pIkgTYYI3pQKgbWOulKMKqxVUL8VQjrXiqhwRrP1jzPWhTuT+k7xVlDPiYH
OTWq+EawaVxP9mC5CsYlqv3mOfgubPeHGN1MS3TTNS6rkFoNYFvLQqAf3DE56iGKLDgs0hTis9v7
eoRcsoc8Flhh4ngGyXuhZfp3KiKIbuPuWPMALwXowsbWWJsEvQ9KLTbHkCT3L2EYpNAwMNILwnpg
/DMw4tbv04mYmnw5/OBwSYGNfw9/eDDcWp6xUEM2FBAuRV4jNGAMGvqr0hsCrjlSoEfMKFCzGoiz
rK0jZnMFeVuVuoY4HyvX/HFZK/mXu5aAMlb2Gy4xEeRDCpnDF2CmgMZfnnkUsDtVtXSkNUnEOY6V
RGFtjbAkdmtBRdRxjXX+dVeGNWFI7zXUVHhHrmbyqqnS/CiIBOJFa7AiC0U3/RYXZthqW8hTY5La
0tT8pkap+Iz1BCOZ0MnmnEEpAAk7ATxdmUgSElogAZoBRX7OBqEqWHiXfJQCTI6uP8IvVIrrQVMd
iUzsQfK9dgSk+/2YP690eKolEZguL6Qp8VHBD9eeXS/+SHKGd9PF9+euVGFe+CdDT5+O7RsF26Uh
s1AW6UCkKPpdA/kxWAdLZ9Vlas+PI311WVMBq7LzP0H4TCvRl2OnMVt3st+D7boNr4dLJDT2xD9v
vBxOvdDlmFN4C8AKK+5ZJu0ik3UelPm6H6OfjCfzMoZI+k8eDkc7MQCT2JmvLdHiCy/m/vNW/krE
lFe2i7Tx7q/8KmjDA0jiHa2hwsZhpj/0yV34ZCLDSTmNw7wPuc4E5dRAnpdXWHLzxxEgkCCx/ZFu
zh1614D2bgrn3Wgjpll1xJ58sAu3kZJEuvUxAYhscyD9AD2HHWghYslAo/F7ePu4BCKjf+5pQtVp
yCty4k6GZpAzcNTG2UoIkBqvr0FMTRIzHO18cGi2/hm7cvz0BOt4qw7x1jbE8x7qgl7MQfIkG0WL
fVYkw+j8TXJMAqfxzpy8JMq2UTFv0pFibKL4Wig6ZEkUJe23QoW/ReL0g63rRZc0iLyp0gNVHIhh
che7sRfkpb66BVxBkGPsgAu8Hu4T1SRB+bdr7+FXK4lzQxeAqU6COwyw6yLY/94lSuWZcaMKG9hj
Fbxn1Vdm32EWqx9YLJMtvWDgLCTCpb5IAkc1TPIspO37tcMYQV2pZjuKVh6UCto13T8cLWmZyaZv
eCU6PjjaWGM9Q6qrLIOkWlvaCcwUjrz/JJoZsZrDdvK8vlaN1w1SuXnLW1EWoZUOAdScPl8v640O
WtiSZKKpL/DoyPamQKSn6g1vXwLqa1HgygeT1qLK6QkB+1d6sAXLf+CeqVST0sC1iwf+RrZ33RXl
QvLeJEIpvrFRfUPM0eKPX4kUy3vEQt1RuStdE0rNyfQjYblyInybRTZPNus28okCjNBinYMNzgdq
xF58ZMSypCkpzpfRwESN2C2H+Tx8ONa2sSLyeqMG1ghkSTYNi9mwBnSCPk0prLjMB7lIy87vfnk4
T8Hvg13Ap/MX1g2csdV/PCpee8AMixO1ojau673KWz0whsnpdbqs1ZoSrCyX8vk45UHcy3dObk/v
jX4jMGRKu8fg2uwA0im6BJBkoVubl6R3Hak+sA6YNKBHTVwm7FcxegAjnciY7/pTNfEhfydXmrlp
jhbI0gm+l/7TzDIGwjdISeN2DfH73BhKu738gd10smxlqTkrcPu0vSsbl94zjBqTDihIFwZGBT2+
IBjr4DBMGYCFBcmXH4+ZlarxmSn/mAyYLt/KFK3we1BKzWkWbCB1luCagXEpqwqeTwGs2ldjVlX3
Vor54vy+imDiexR8LI/AZJ1U05XBOFrNiI3XncrBbOXMem8wMKqh6yenHSZzrcZnNQOypR9WT4ql
NebWqA9njIiEVAmBWQcjCozCh4nx+jqhDnavuS4yXcF/kJm481Hv+Yra8GJ7lumJxdSFKrMCp391
yg69l2vLI2moU5hcBUL/l+vohdfRKs5+1SZzuLyABULzuWC9BqxjxamZMSMwfsAl4dLmebtZj0BB
U9Lg5lO2qCReoxL+AtOfEWCL9zY6osYZd+A3g4FpUZ8nhcpYN0WCQnaO5c17H3OT0g+AHaxy3gn9
a9FJ5ZcBGq4FgUzb2cdR+GK6p81nAJosNL0FtqEieEXYFtHs31ZWuCAtqKPulL07NA5Nfb55jS3d
zixoLDHt9cszZHtio6CC+PtxPbBIrkzeET8ylU4DvzIDhAwopheYOLLHV2cbYcvk7XBkiJmqE8Xq
iS1P4QC3NxEr/31/ENFzSaY7cTrr5WNv0OdyrKMaUXd0rTVGqKgn4tqR+pUwHgdQTIrKd3xSHDnt
4Px//ozk/LXx2wVsX/S8OUbUCPKTjUv9MJW5jFo5SvB2crTpBn0jkhBPRTn+PCRHNABgnQd3kdW2
09n77mnW3B+HUEDeRxZKS4KA2/GyeKgBtpt02UNDKakG9lV90GBpwb7DCuh7txv/RmvZpf75H7hS
mvhMogLJ2UcUfvnCh5gfNpKH24mzPW8K+cEJuq111yLUUD+PVMT6pMaXv3Ed8xa2GF/nJ0yhQB6x
ygjooS/FNlXgFLQFjtWIcV3lEgAzRkyf3FUsx8WPERRdw9m6w+sEwCBPaC7KhvaREfbzbxa3mZKZ
OJE1JBScibIaNsIoOW+Ob4h744vESUyeSQe04chu2bdG8I+ijL56wbPIXRqJZ0V6e4LUulZVtc2l
Kfs9+SoWyaSXM7qg/gquTnpkMS+bfQF/lVdQuNHwCiixxPFzrY+lrAEF4JKjvcKK+MKokJSiSqA3
YpchKbORa9i+LbxaI3JKbisRtlVepsRMhUWbDp8+pHu3bj4ctfnF78dZdurvXZIFfbK37/KM3Tem
Pws1pZ+sMw1blmbdQGOKWtD64GdcdmanvwFFlFt9rRAUKgQQ0DfOSmB25zerLzqxxM0aK5q2fsh3
3uX2H6dsIO/u3fg9NOTYYcBlwgZH/9L9Mtf5VQOMKU8nCQ3gmu3n1GZyVgeNMMAuuEexABVMv1Pn
br3yKTm/3a+EQQ98xjWQZJcTPw+C2TQYiFQVSJ1XczsBViP/N4VE6AlHTc1+URLmWBJtzqGCWVVC
MNXT071v23P3kqRs+mQS9IVOr6DTfOabTXR1IRGF7voE+SpkKU+43QMYyUTlIUWbPDoJbbu5RYnm
WinyNdEeQdmmg7qsKz9TQerteXJRnb8m8tERnVv//0PBQboHKOBOjCkWQX56twgqhnZxE9zNDrQL
adXVbH7KOxKOLVKmGBEcBKQSYTs/SpxV/MiUK+6JxUXZ153SB2y3uUc6tygOsaHu5Am1ULF36qio
1NApI60hIxXCmPyLH+DO/ohts10fLektn+jPtE+omXifYPO6Z5DUgppiUyJLrEHwXnm7k9sNOpqw
rR/c1kDHUIloPBYjhC0GegRG0GG9UiAZi+upQVqSis7hSrDOg9paE8FQEnuqu5uG7Ds/PwTPb8FD
JNyDZFAFRMgf6dfOA6aXNBgMas9xADGAdHJGzK9KPvJMdiGfY/tLY8+loZUgx638PNE+MLP31NxW
C1PCt6uaHOnyi6O6S8bBZQwWeBimb2aNfWXFlREYqok3/D5rH5ISOHGDrCEwUk0JGWPhbRsm+sHQ
wg8r6lDXsFQzR/mWgUYh7tZk4UfTA1LWDDINVwktm/KFiAT9vb3mi1ATp5hDsElkk6RB15ZX0JNy
xuPx5sH4/fwOL1ndgiUpkNCPe/VilE0efDoYmesRyi3SNCI2swSwRIJp9agJ8IUY8Y11daFUlnMe
MqIaKV3eCSYoBfL8y0V65v7jHJ+m/J/FrgU6Jhs8bj9zCcC14Vzp3zZQUwrz/SxQimmZoyv2l3I7
JvJBwgxpO996pOkfWnodPS1e7EJhR2NlIalFY3gC8XTkukIKV78xxQxvjfSvyWAsegXsjg0lZ1dz
VfVfLIUwVXSWUeiGZqYxacrTQJGvK/7qxC570qOPn5Pxie21s3/HElfgzZVtwdRQgyeWKvhNNvl6
LU+GornMPmIBL2jpTnWkuFMYYIdzUu5Jom9EfWjZ4sKNgKXQtGtXKqs1XEn11SW+pEzgaSetcre6
uC/3BNQjalbRcbGXaHnrYmHjBsSSBYUsj+Z1DReXFg3hOc3YtdmeV76vTIEUWc43kIwjcZSHqW4D
UIO6IG0fX0r2j/LoWD7Qn41sujmHGZ6D+2jhrCaYF9beXcw6LYk+75uGz/+FdbFuoUrUgxxPvzSv
v7riInnpHhMC5YytRLVlrkV9WNoZFgXmZaRO6riRJfBhSeM1rmm9cEUQcviWGnu7KeIC/kzK2xD4
z/eXdYOUgPORgKJwaTKHGRY2IpuU5Uq+pOWMysA1tycTIxLkj+9tPnrJfBVK+PzW9bm0VTNoMvRO
xTvBSfXIUiyI4uguTW0Ttr4STbKCZ8dSpxgDvbUA6GjH3PAsy06UObXQyA/nQfeOYy6zzqws3m4R
in67+58MJSIHccNFGhdDRovLrzV8au5fnzrU+pTsRPHAwhbPhLi2TV606b7hzRdRwBZOuM0BKAFN
pYfRP30mDyBcisG0Hr4Vsv3g3sh5ZPO1Qfd8R2zOgiPAVO3bBg==
`pragma protect end_protected
