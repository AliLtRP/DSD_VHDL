// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:27 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SqH8bhLXUavdlBJTevkcolMqtj49FgaKRD+GFGfzUai44BJFZW1iwPR9WKi7/xLQ
T6RFUOQsgoEtn9FP3yosOH+MTCIfpJJFEVjUgzzvkLL41fasPBvz207931MOJVUu
zOntuCmXxa2/Jg8+9awJPmCCAEfnZNf2SeX818vx+lI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6736)
FYo0w1D5L78d/R+oRRyJ8V8MtQ2/qLFjhjgARrbUHRNVJA51oR0tQV9SsMdSPvxN
OkcgJRRQsitf/KJWB30pdOgIwRiBs0mGhzH0Y2OkQsNiR5BQOSJS1lxe03ocheGZ
3kxBKu2r2ZSV93oAzoSd80nze8vZIIt/QLa18tZAUbNNYNGKHFN6BHeuHo7mU9SF
DE7xPXoQYWTyj5X3bDwHqsr3BM27f/H2v9nNHe5+jB5UcDkafhdPzhW0/lV8p9/Q
CLA87zjrh9PeXO9mzltVtkUSjPqglqCdvN4BN7YzrrNARI9pnui5N3QP+z1QYCB9
Yz4A2cGNUKGsGFGaL1XqVmvUrUug1V7GEBI0rHSKPFm+KMKoUTfZm0qsk1k1KSdo
3gBJZusZYKVKwkUx/+z3p1ago5+IpQzHmo3aFxxtXrmpUy8yv3abOIEIAPwkD51v
W0ag8U3ExKPD7Uu4+oZLSPsDqPSjxGHRWGlOuFvQ3FAOIldKAYAc9srjxBQmFxWe
mHSdom72MZrga4u6wn/JrB8kFWxUgc0hHJcFB1ALco/8Zp5f37ADx7QP6Y6+7Y+A
q1a88MbtAdRRYbgAydgVMsy+I06bbo7CRNjcCrkuVvRVSljBLhEW8GHzBF14MnIs
CZITDp1e07fh0YHukIKOX0HVQdUY22UPtqfcaRJweDMpWpxNXirLwS01wY11CAPX
NusB4TqfCZ/WurCbImQHEsKcsVVi4wO4NZNOIrPANlKJeOOyOLxcwqtR2WHMDiOF
Ftv9OQwzEhZxeFO6hSCpmF7ty1O2/BNNsm/v5uXQ1em6hSe8lM01R3b6A0GNUoie
gLPDZ0hY+GoHj/VKJJTpGpvBAWaCKCtFS7/TDjjDqDfmPMxSYb/Mgq/cP6Jz7vGx
8TRNNgEwejkR1NXHj8K7nKPwFL95goZfFcEKmT/TdpNLhQq0P/CeEUOherVtAk11
NLwa57iu91psdEcxwLeNItDAkrn6P/l3nGMHsmr4aWURpsYlGxLrRAl5+12Kq7T0
/XA+tngiljcL0TiVy4ibXeAH0VCqT11LskNRy/boEdMjGtJNwvMIJP2WuTiOtKoR
1p7lfmF5duUWrlC9umEearvV9AFriNX+x/AgcgDshAgwwduqdQo1pbdc5PHdXVht
SiR+swdYs1TeC8crRcEaMjTFBfTIm7lpQkPhqXxJKKog2gYZe8z4StGFJnMX+veS
SfUIgRU5AhLgbVklh3TjxFFiTM/U6t/1toCcMQZmZAXvhaKnGfnT6eat//sY9tmf
Itpl/CXb967KQQj5GaQ16CJXZkScbxuEKx/wC0y4K3K38gWMHcLte2mUYm1PsHMy
GnayOQ5FE3lNZngpMKZYw+gb2gvD2KfpQ8f6pBumL3tJArG9fB/V7lATCkVJyFFi
6XFLgw3MYJea8VTaQwF48EJej6q/kuYCiZvHzgkhcEoi32tyf5kWdm1DsiJlDEQl
ceDJihJo6KT13ITWTf8qq/nW0uNp7aKpRnVl6xU+0iTK+xMrwUKT19nyQtk30o9K
wW9+sJJsY9JmualtZzvN8CCJMC5HRWYPdfnCMkjLtUl7XCQ0AxHmzB07ehAr9a6H
J1Y9mPWvSOD9YschaKTynPCY89KCh03wHtiZugf/u5ECcX5I8pmVSOlsil95PzH7
6sW8iCfg3+EVf6Qt7UTl2gbpPkSfnOvWh0lJrOmQAku9H6iXfUCBSbPSFk390lkU
NhzrDLNpyBXx8RgnHY7ACDpSpkuI7VQOtRo6Bhc9F/RMmtzXiLVcwjebEnWK16nu
LCiyTe+9kio4gadB7RjRLIX3pLoilWXAj+KHSQxSpfZshwfDDGI7XFWkoX1Rth/V
Vy7Zl872O/PXXtKxb3cPqFGU3KZ26M3FTqI3NC33i+D3Dt7Hqg2d/0JHMLUY5ZRf
y+oZE6Jxg+Xl7zYWOqF5WEozSkGVOLhnH9GzsqtrF5Uzbcvdh9dfT6JUk323aiKK
88lzuHTX2lpjWX1bmadgdI2Av2ardJet+V4ffF80NDuAQELIcQ+jAVOmiApbWpjI
iPQKlHUnkc8g7qMOBFAfKEth+o0y7BfjbT7CIJI13kS2IYDdBDp39GDQVc3U2TS9
1tcd1u4ZsLtRAiK0nY01aQBlQX48gw2SOhZy4oSj2GXgR6yI+/uISwFnkxRNpQC3
VEDrSseUkApuzDfWHQj6sFhlFMvBdDXWLqlFqubvkHCJlJrRwXihooA2PYDuyRu3
MBlkIPuXUD2tBaPJfSJXwS9or5msx3adepvOFebjWaeuhZ5aHRYhZkpsNcIVwOI3
3WeLcWXKP2N9Anih3lBFllmsJDTN/qh+ZFuppxFgtslKrR70ziqdP5SeOgS/EyL8
5IoUFl+X0FK/T17K5+EI286YkgJfOrKOj1qALBzmq6B/3tRTBrXh9HcAwBZMTJao
8yF0kbspfpU45dVKEc4FBDKBJ34j5hQNwRgkYMzT89OvcwmFWeaA7suUjTx4xHrj
vYsPFLBgz4qBzgr7dWsddDnIAgfHjZAw2Ely7XaDH7izSilt7DaQWZqu+00mwY/x
on1gDRKAvsyBgy7IwRYqQ5QQdaU+im2Kdv//5b5Def5mVqix3ow0umM9gcd4SYf4
kv1hZUYPqP5UfuP3rTZi3Dz6Gdxn/yLBHgAzdCp4VXuuKe/vC4I1Uf1FelHueghB
r9o5ZsrFLNCzEUVhEis3fBPKtmAT+iooKAN+WmAXTybMc9e9bGeNYB26vO9SmWws
m4+b5eXs6JIyJ5XJLcOlj3Nc7yHio3JFBBFZoGytqOSzI1YhHjx53oAhBhWV4kiN
kDCP0lp9cjuZYcstgJsm/V5QpH306/fqUx3GyWKS+P3hM/QUPH96mx4ul4iUj8y6
t2w27/g8dzg658bmX3NpgFRLsYpPbLHnZvgpBDpPrazJH5fNpZjti23G1I2fNmQp
IBCCf+szDAJBDHNSVqZy2unqPHoIbB1Fe9l86aYrLR9If20hM6PeB4+upFGbNYUx
ZonFjLVd+GhtXMLFNKENUmI74Z4tQ4stdpOC1UP62IzdjQjMhraCy/hXV8c9rXIk
3R+1cV+Uvwpy8ugjxxCG99DtA8tMlKRu6EaIXsEjy6qrPf1SORUKWpezjLM9ZQq4
ApsRm3krnUZS/leUF3hjqbdmzf5b5NtZAcfx583TYE2iseTDXdg5kJH1DB6LgDqQ
lHcAFX+v3VqsSgfTyV6QQrWZLIBzYu3geJxgLPZN7Gp0UtCgjsiHoy+t5RtOQA7y
dD8MweJTfx3g34kEyXSF78njvWIvmLZUXHhhPHEN1ubSecVDt+QPU36AEjy7qXfT
ijMeBwj/LrSeVSnOYjKayRNIODpxkT3rFqnbTQRpHfbxODiDEomiUhN+dmlcDYnv
0UwikH761YcjNsDIeA2nukVhiv3Reh2J+pi5WgaC4ZDMxpX4B+XTiEefMjB3CCS0
NXtpqMIF2Jx/9S4LMZsli/kidnt7Xq5iuo6eYfaiPS8+i8k5aRvBFdPgT/7AgQva
rWtM5nHQWKbPaAFBdBK9H3abG3R9+ltqGcaKEOO9Nk9LDIhDh8IQyMbhwUNJ/BA6
Vy/i/DGsFJJGvT0DcDUaiRan6J9WVlh5sLKPbZ2kbp4WWGpVtjDJnY/WyKicX6sc
HfowoWbz2N4jV5pfFjZS2BuMTlkdkPUqUHGKv4P+tyJ5tAaROSHtDXHFnIMtuMps
H05TRhjsEnK5eOlV/liJd/2nHyC2atItiRwd+LBSDCQ9MDrzJT17Bqlc19Bm1U4a
PcDHYzC8EIO1pb2j0V1z17gFBt/pNP4FOEjI0MkINOXH8Cxx6Y2OiSAPXXbHT4rh
Wv3leKfIxShGY6IHulTtmWyV8SFJHgqio/vB3gu1oXZjnWENTvkIH8gK2R99fr0N
HupdUUct4YgiE+QT0hzMextrY2AD2qfL6a5y2vz2Ib9fatHB36DMcI+dLHUcnNkW
t8QDO2FEA7O6Pd9JOV9qJ167fy2cFHQocAA4FaVAzFkPcri31JNtBiTmV3/L4O5w
AckUeTGJGoSrZOYEcJr105cM7CUs0pAAHEMg2s1C4o7Yr+VYlMZvysQMdSQzUUtK
99fTWi8AnAFC7Sj8l0gMBCtbAZk0groh6vNxlzNITJtc3o80BL0KFa1Ye5U+BF6E
vUtxPZlbGqLuFGvsKb7aII3lx/HmuVnYB+PgDQiY0dhc1S3dod0gG5ZchyUeFCTG
JI2DkGQwg59XdsAgMmBQgu2a/3rwWBGAya9jBDl9V4PGW08A30U3A0bwdwDudsm4
E21W3DPd9UzHBEeyAeKUIzeqRET61QtJML9HLAAvuXp1aGQXIck4sDf4yZBRnAkC
CLrHk7nMURkjUOGezzgL5uiztDv8HVTt22ejT4U5sygpk3mkicCo8fLOFd7+vCTB
mcBSkYH7HW9FJPnRoKWXCZrQY1HsFlV0oFZ9kAuYqr77Z7DBrs73OQbwpnXotJ8m
j1QW3moGS0b/ksM3rPkbScTz2fEpuIeuPD4igddrsgxUIXcW85OxyLhqV8gwJnOq
Xsz6wAbSnhWQHY9MwrLOwDQPwvKvVZ+CSsDbTkIdurHSZFhN2fWLpieNv3bZ+QD8
SxfrR7+mvRtbj3zSJ19NBoIyrGopm25PDva65VfDZnZoyMS3xPl3yT+R2H1aEBWi
ms53AcUbeuqyCB0mvBrtc//a90Nf4541rhcO0cgvSgsNKBFvi4+3hiB6AW7cUyRQ
y1nyOcl89fjtJqMunDzcjg1uGoFern8rElDjBFbLnwizEdCQchBhz4OBQLiJkxWq
xpllOoUlkmGnYX9W9bB3S/72eBJKEnR/ckbkbwms40S5L49dyX4CkcDbLobMqtEz
r0XPGT0Lh5683T2E5X/V1qcvWETGr37T5/WxbXWypyrRm5y6Ymnin9gI/iSK+nw8
Lk2Bkz8XUaKtSCsoAak/9IInPH+Me4wFp2ApG/ZsowBq3Hzm8o1+iBjURylkZQz5
xyKKK6r2IRc893vROgjau05Fb5PLxGwSnDBfVJ0ztPEI3gznKeSQZJrawq8Al/MB
iGwAsA1DMBNR62r9kTJMEVP1jhFsYyEOBqf245cWMDBtd4gPkleai4O/nw2G1dAG
GoomVLCYqNjzZwrMH7zHkZJ3KQ31RvQFTfKOcLGSfAxU4GsOZMNqxiCUmlMmm+42
dpP/KbbruCBHBRsFpIX4HB8y4D3FZ6zBJ6bH7385w3fC6Mmzd+JzHb5NJDlyft98
c1awpW2tTFRLdjHgHD1m2gdev3U6O1CzBsrVXd4cdfn3luSq2FvNah876wgpnXTN
dxYAdb9BiBVP36I4bACMR8fOBH/I+Zg64gIJZ6c7PK7W/bGnVb7XiyxMJXUAGdoC
sWTNEiX+OsHW8P0x/1DebjpogG1FsNW82JmrpWXDWPCfv7WkHFvwcGpQLyulRmUT
l0JGl83dY8WU5iS63aocHyXt2MiMmHqeYi3j/WrCvfa/W+cgrIHovYzxJ1tDvSMO
wRaNT8LvfDQInKZIwHM0K/oS9GeOD5t93tARYCEsLto/Q1Ad6as1QEeJQ8jzgOOg
DP0BkBbd6Nz7S4LlRmE5R0BiEXFRj9A93iGk43xuOLBOnkl/hcAmW9hK+H+o9p9C
EvnA9wAtexDD6cEeno5g8tdwyiBzUyLC5HVp2tmAFR6ynJYM/VbeMRV09bSwLn/f
Y2dqBo9rV7/Pj0ek9sEAOi2VMEJHKOHND7qMkirTPcTXRtLWluxzqiiekFiQfLDJ
3R0w9eiq0KogANhVQZrw+H+mndF5vdC4FtgAdCEf03KG0MMDQYAMHuwSE48cYZ2z
z5goGML/paSjSbmY2Yh8RTl6n5aLHNGFpkzs1QnpZQApcONUlcAuLCGcy4rey/wk
AYLL+kenUc0m44JSIIEXBeeI2lGQM4S+OmTa/FJ7SpzVjaeYVQVOK0LklBw72pPF
MJX04mGpJscRrX88NE/M9SO3gsQBkdALU0SBc2TbdPAEsWG6FbgxnAMINwxAC5Hc
/NcIMcBLbG4jbmDr9oKb8PtScmXFLzljvhVycGHWXvEqqyBSucqq/ob6EFspf8nh
eJnZ+4eH/fRYyLnOf216IpOiQF3gnnPAeOx/ZWzZyTcnmBUwcnDcbEp1nhubetU1
tIgofm/Zyv3j8envJNcbghjBHiS0y0niHtRVaNo8PshgfLicyoL36vjrtmHEHknJ
JVHF7RUE0x2rsVW6gFfitM5Ht3PFsKvv3x+y6qL3GT2GfB6FtT797+PBkGNTVOFk
B2iGNf+k4rnZSEtJNHiA44qlpyKr1f9s+Nj5CcZaBGsP20RAFVlnwOHHF1gzh3Mn
3Mk1o0pH3nfjW/lbOqqz0C2QWk9Z0pUpG0bnYbz4zGj3+yFo1ZsrU3gW93yjvpWJ
JuJBGcal0hQTdIZszmjUSZVOSHMfDTafqVPrE/j9JDLaZg3XU6u7EyL47VwkReQY
lKeZ1WM+9fZDa4I9B0ExetQV3qAOgvuqjgfQKd1p3aYokx8Iiay39Ly80zB3rs5X
Ce4aCwSHPAFw4djDVk08NMssJJk2H07Y+CT2d3T2wV7WmYVSAl7wHJUqSILvEPOs
xeTO9HHWlaP6TxwPHCq6QirHsZfBFshyi8A/wkJLlzdFXp1dL1FQ5wditgC2BveP
e5ui3dAGHff4+ktx5evNiuQ102U1yFiBqmGMiZnhdhe6AEVEKC0pqtu60Pr3a1Sy
3sJuebTUmZeLevz2eCI5QJjc43taBENq+FbyH6HpeuGGoS77mY2/81+cqQg14mNK
V19WjZds8ZjLMCm3LCpUWh8HmLonQOZCB1oj5zGsLahg7UCmD9fioiyAPhOGGEth
EI+e0FzfT1S1zCvPO1UCGfwzEAEVRhTQSb33TajA2U67Gx1afwy21pd6K2598mdp
ca1/GRkqzcbNsAG7udRUkSLdKirzEtRnEJHpYdIPrWUYdcDeXcXTPrBS5b9Kj2wI
QcweHXuUeh3Qh58cNvZbefGnuiE8SN1cqNoE111g7MvJOUNxvIfmCqHKe618rn2y
UYgvGEAYeFYIk5F+nakcjY20L0mTximnLsNxvK8Ic2wvVoSzTq9eXr6GbCRg6gvr
8fNR0cq+jIZ6jfH3EVHtISqnOs1PcFKShqMXR4SQ8ThbvqgxIe5XIvy+6nnaLkFw
Tyf5RDHHZUsr7XLB2rGuPmJrum39ubqdgcZEmvbjl5N4xaCPglIXpP7SPNv9FdUL
brarGSxXaE1E3lTi/YashmXv5Fqt0ANT+8NDe5lcqyri1r/nia5f/r0yEcFrcsL0
HsWBtfQUzLk/QrNuxtfsqbF/GS3W3C68NSC3sfyIptsfyq5cBa018pqRg5iqKyrK
4m4ExOPReMFwPicMDXEeOjTeDmzZJJ6h5JUk+9Uz3wU49MwEmo6uiXkTEyX3KmC0
dz7/SR5B/kSwDqGrOEnzTqA+a08JcUG7gOjLB7eyT8xGRV9/zORmgIo2UufrHXHX
+jnYPXYS13GFSyGcCPIjViK3/21fO3gVj5cUUvJt6iHG1HqBx6KizuHYt3eqt+hA
QmQCjss9S7WMu+0sWVfgQfcvaAMtviLHVILx5Hkmnb7DmHIWrEFG2KudtS2wbxUi
EXUTrKBZzixNtzDFDIqMlhuJkQdSHn2eAFaRYJaGahAuBPNYKyA6YHT5iTxpKFJv
m/y5lnqNGmWN6BWAMryh8LDV/Es4CJZ4YrCxzlDoFNU4f9XE0vNDnXVwM1D7T101
6AOQsB9x2Zt4x3ysZ2pzJjTbEqViGUrkC1kG3Px85tyivlv2AGaxOc3Z+0JfFXrl
g1L1ikzy3nLGZ7atkdArK219VG96fGQV49R+lcVk18hoLD7zdeLhlswHgA+qKzXr
ROE6zvtZ9kUKBTXuuUeMs7szlDmY0D2Z0+FqnkawU1KZMjPfobxdenOL0N7op/P1
OvRsADctFu4kIZOwCg/TDCwrtnmRMEFgB0h3jEmHOhkyj8QFLTTvGzvry+T8jIS0
lzF/bjEM04h0/6XEiQvpLIApyOJS+n6X6loVw2zb0H6rI131PVDK4ElIZmEcb0aT
1NrBOq862kR2ddYDyhJTp0PMmG42jo2DmnnjRmuNHmoZ12VxsmbwtVBaMV78uy60
e7dxUaobzr1tGUoDt1cgL3SsBDWM2OL0nG53bEphZpZ8c5RoTFpV/PsiLUeGzPeb
sglsnZI7ZUFGCFE1yW90O+rD92v03rGXGewDm3MTOTtxlkQvs8/IZ0MnOf+9ej96
dUgfQEzidm/tASYS7ugddTdccha1ID6f3XSdLUlN2jEnG/zYcFZZPTz2+++s6NFB
ZC47886R1r9uSWXHr/aqW6VtpoLsytvEDkYLIoA7zEVtAwCenvFbc+XOn2AAYaCW
ffeXCEB7PpsQ+4w1Jl5sKLuS5N64U6uA+/GSy4dwdL10iUpXBVbl/ohtbtrze5Qb
la16s/IMgylVzp4ODVY9XKSzq5wAl7YhAMQ0xcVwvqv1xKgk5YbSYvF3m7GP23Ps
3fEWstvmj+JOppj7ceJZ8+L4DEwZZWT8+7qDqLoS4TAzG7p2TL24BOMF0ZmBhc3l
grVyrICIJzUrprD9dhL/SEFCAfG0SEZRuZRKyECxJxZV1oh+Jr9SRJdyB9p+YT/e
pJ8AghtB6kFwJ2HpUafVTALMOXL1CVjfJXKG65Wh/Ntf5QJzV06rATDYwgkeYkJe
ZHAnvFMqQMXqirQwjBLOfrWhahHysPqzm+Wh/w1rdCnQOoOuIrURSZItNDtKZCfw
WKddA6/djxg74UCq2D5kPLRUxbeAGviIls/EviWRRAT8kj73kfz7/pAvr+WOhdLO
Yf2emRC4/NqxodXPKDXq12xMngAvO9GpoyCeKU1O2vjaEaxUy7jHXCJ6rWprJhZw
uEkpPbOYLwqG1BSgBMAzZ8BaEAKaoeIH56igfOGcm3VT+LBaXJKf7cBDQJ5hVJTT
mZwHAra1YrfzOVBX67o9sQ==
`pragma protect end_protected
