// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
o3ML8w69o5jnjeDcAEof5rvX1RpFNDPmxa998yj5SXfOzh70Q9kuQmTNP6Sd1m07
9riNQ5XMVDGHP2fSUZPCET9yZm7u6SPY43oUc2laPBlsY6B3seUmsIrH+Q+VqKq4
IIMSX9JyF6nvAqZhYgOsj0pdfiGlQKuH04NQZIP48Ww=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7872)
xqwdT6hHPg6Lb/Y7KUL4cTiDaDd+DcOHemHZXBDW8eHqIt6lQbSjVOtuLOj1ThAO
/7vt5ImPVqctaoyGiDGNvoJNZXli/+Mw+tTOP51cRjxFN4cJ8tz3+OZcW/MVrqHr
q4/ZcURiA4MGd+HWwsA2F7a2PFNNd90kb3y1EAcPAMBBcsvUunKv6/kVUL0CVNJP
zW4uhV6ozLVRQG24G64QQ5THspxZARro4cdtBfr6Tt2hkMYX5+GWbsW2x8LiiQep
hvDHBk6gJg39Wex8/ChfStIc955KkDMpNIA2ImekznoWaMuDWdcsUQBBR/9YxrdT
oPUf0lU7BHhSNjep6ZKBFmOy57PFRHx0WnWCbhhP0bII+ibvoeodSfjXMuZkffnT
xOwJjDc/OJkQgUB8lrZghfgSPSDCRaQnLXgkR36x8bVeb8y2hICLZmdeiME0W2nP
Uq6lHNYNanNIVoNMf2ppECKeM9aaJxq6IPrZKp/P54xF77J15ouOI/8cR5XILEfJ
WJ19kyt8ndhzQpPnX43wAmZDTSCGS1BIqR5cKaHMc4upkbziFFW0iYjVdBVkR/MZ
KB7UsEZjAdNey53kN0HqD7pUzwQnEzzJI69PjXwyLEIFyyO52BeYamRr0gexxQQK
VKyn8+z7d51BFCG02jL6mMC0pgOLLwG8/bagdYx3jHhZLvg8X6JE7UPQgAyN6bA/
If+rTbYhfM2wGfcG1EaZj0B2s6jNS5fi5P6V6TW2yDlK7idnl1YBK0iMEt5tjpDT
QJLbZM33hdkcI12EhZ5hlZngmiw8TaaOjZ/O6Z8rr7XvmfWGmzbm9MBL6z+TmYtb
VWXJNSfj7q+6+g8f2IOw/+lVCNdFNTy6/wko015yANj7pL/ZNcZyvlVJPpdX8h2u
s11G2vm1+10IqjrR23r4csfC1RmA2eRS9EivBYkr9yuk9BpELhnloWKZj/dUD934
mpK6i71HudCZgpNE7ePCu5J0vPTTjvLZkC/QgGWw5P9hl9WEOc3e2hHVGhsLPXyb
ygDCRdGQJH4avke8xIbRl/j0zUEHUWidQhimAOmOWj0d7e9acVp31gdgYHq9vhUU
BYyoADfdP2HCYAt8vzoGx9PKo8a133mtNrKc1pWqmssbleNkRy0BM9sTIG8ERD9e
B+Fz49oW7RlXeuzfcb8O3u92CD099xTldefAxfmh2MTXm79jOd5CSLdeHrxB3shD
VCEA57AqbzuPQ/UFWrFHuohJvOwLtFVHNyZDyDlnesERB/2IAGG3LO7ctsVz6C8W
Y58as2akVRxHl+IO5BxN+kiUVZAAZoP0qAAIQKnbVKN2FIf7ejUivlPbmF2j3TYP
WgvA900PMReVD5GDblipF4t973w7Nioj5FjBZIibJagZFh1ruj8yIw3vy7a1qXVg
ae7XVFCQyuq8bHwI3HgUSN/cSEbkQRvNeFqf1Wzsa42AaX6yPpJIhBshPU/JNZUo
+9MHJNOdcX/rRRl289tRga76puSdCYPCc4sbq+Nly5KjavOKslrNEYSQ40gEA62Z
pRrN4/TIYik4U2QHFP9fscaTX9MUOD1bKAhRrwBUDq4vj9xvPOLlsDFWBzL0fq7V
NSGLO/Gup3N28cuh3+5C0rPNYTOTMaqee2h8p3rwcnlrAVr4Fg0P1FXtJ7556V0v
G9tU2jYj6uPcNIQkyPKbmHwvhtKpzqsOUt9rHzLw4WEi31wRVEcpazD/iEKiox13
9xg9arFuV0974P6n+0r3Pk9NSZVzIjHyo/aRY2srhFRc1f67B79vy5ceVFJccBRG
Z+7x2m05n3VcxwmZQQfZYG/6grh2lvfo52sBspeO+8xoHLy1vNDJYhTH738JY75h
d/HHcCk+E2iQYXRXLe2khgY9nKyCvaa/wLX4rmWgpE8eZN/XSqIhW1n0SW0kXIzq
LNW18JdWUxKO4cGlbqjAGFUEG+QdZMbodRdv1tAigqBb4/ncxeN52VB3ydozYMn6
wfp0chuOFRn+0yus+HkErBoRi9/OEwFCQ+zEARvzf6kCaTqfPO3pXy78luKlsFU4
np0z27ap84s4zLITiPWuXupoSjZT7PDZkA4jbBUu3z3Mkwi1S3Sq4su3GhfisqCx
c7K7qRsMQk5KeUpXwzm+zuFLJJRF3qruWdhcgUJVYmOZipr4Jy956NiXZOsr9bxs
24PZ6Taq9xEX8AePScId0tMc5/ZrlwkF0diUFW5GvhaJj1EhTxoUVtYbJpIrYe2c
zE3+Xlbw1id5bpB7frHRL1VCcBePri9a3IA8aocC/gRtDBw451DgktqFplSMRq+e
hHcI7IbVHgXrdntg6FQZkZE5kslyRiQntE8v4hSc1JVwLZjwKtrSOANak3Y6Qh6D
Gib8d7OvLS5bAPFWbNOpYC418m6ch1n1WykgrNSBksWb8YfcFEEOSkoeGle+4Vp+
lXia1DH20R8xya3PNBXC4cbsXMi7rdSGHBxQru9eocn3eupjSAk+3ejq08e4sq7i
D2JM24gqCZ9Z8jnaLb+pMcPw7UcUxQmPU+RJu49oxxPlgW0BvFPwDrSxg4kb1itn
FKX71fUk/D8INnGJgsi7J7nEhD9CSdedMeh12GfUoH0n36z2We7otxnpwweZrAQF
Kln/Touh0OvNRGQW8S3mNwdf3nI0lcMKFHRYefKlOaXet/LdYTXbvkBQ6R1M4qIJ
WeuFNLzh9rDDiKtxXdd+97Dlv4byNR61js99yqFfpc3tMWcPuavg/1vPwW3u1F0v
tLgSQniQMljpnpNgNFiCONBuB5LKhbg+a5MX5SZvKeA4/bqtAZfsH0Cs+WVGWCGf
PKGmMBeQssvgO27WokCJXBvdDBJBRTVl0QchIUKLQ8qyW6+qWZOTn/od292uauQe
DVWis5UdhUsYr44n8Kl+R0oO0MrYZM1WQQWrzrnJkVA2MCbVPb+GxzCzs27d4f1x
BtEcTilbwP6RUQhcRfhy5tOCAipV6LRyCpQuScqZLVJBizBemqMqLbjIbAs68nvU
d2wsI6fpbMjBd6LG+D2Nue/69nwurXVzlZtV024KkdLGbC5MnMrWGMlLoTZP4y5K
qBdefpZXN9LLtNTP+McJeh4nKSBpxuDpYvy80orHUEEgGrdmKcG8JDcBF05dfFHS
PKc166BP/mrU4kQyiLN3YZXv9g0eBW8OQr1FJcajkUvDPqMF9zJnP2jqCd0jFXxy
qtinZwpSYsztQrUUQGyLBzOdwrxk4TH6IMszoY1jqbihuYw5CHrPfGiGzKG1zhf7
tgkgL5TJRifDSmi/DZm84fNRTRJnKGVcBhxMLswWTRcW2OnOLMf58YzfSl35vHqi
/nElECeUXoc6bK33x2QlrJUe335Yq6+A04rzgwsaovzJF1gMfQu02bAyUYTblhBV
QO+wNh4OEGUxkjDuSvgVPXPkAbV7tKnr2G/93hvKH57WDw973iTy0Kjm/jrqdrvF
sM+u8sk2PCUMW9RwHTUg9YXB6gxOUQpQN293vK3utZoUP00P3SteNpCe+vJ05wce
egwFdk55ZA9tXLKmGcMvvHkNMKYKPxNLJTsqzsJskgM+0vemixmQqoymAUPByslC
ST9PecDwXF/bGDVFCyDUGhH7H6K2nKpK42Uq1BOIGUJBQqaS15aInYi6LkThtu3J
rSept/F4Sv0d6hXvmk2b17YpR4JblfEXaeQJQLwuS4VuwxPvGqGyRtz8JTDu9gEp
xhgYYumkB/MHdq1wzx33FYlQUrHyfd2Gx2NK3c+k57QH9bsLNDW+RtUJHcEboaXV
zvzl8X+ECwB1T6gbaHRS4wGhUoJoR+vvCSDzEP73AxBxZpF6TYXJZ94GhWascSFj
9YXfPk8CsZpRGYwSQ/nDWcoOqZVXKGTVrULUklQVRbThoRTr1+3CVpeXIMgcupcS
xEZHwcmtcT6kDcPt5PFdOqMkAbHLlnoXiY4A/HyXZHxw8dL7MJLFpZhARTlyfP4b
G+RH5VIp6GRlcU0V98rUc41jQ4KAIK80SsqNxAu83rxglg1QwM4EpWUB6wMzJTf6
u/OnEb7wlPVy4uKS5E7gR/2VAAMBXATXCIv1ZI5prePTKKAgN+OYHQssNexC/Uxz
Jff0JhSXk+1QVNiRIwqrftK1cUy0vAKTfj6QFnUovrHl2NkhLxKDwSPMwCkgUJSz
fIbzEDEDgwdxwLL2x7rX6sYeo8Wu6nvFygetVYc58xl20q8frTZ6PWNk6+19HVFg
SK3J5xpsyIMbkE4GtckplXYvss0oRjkd9vbvu7Ci2kn8NQ3+G8MlxBWC+dqKHUTI
aAld0F5+XcYup3E+Aey4sdWQhVtGrs3E7hhNMTn//XWMSROyOcvFUkwQFA95d0Kl
zMARfxJq+YSnGgX6TNs4fUIhaX/ga9Na0F3NEMvXP3AilZrQsV32khlPTe1CdOzg
IDliXvsnVkr4lxpfnJnHFxn+BMx8wE6GAgxuiQcoOEfXFyTExCdWf3K3zObzfKGX
Fds8oqZuOPb+4OIAN1yUZK0BtL6/qJUCBkax+dJImUiyHEdHCP50CZp+A1wwPtG3
DOc9bywH5To7A7e6nmnBe+R2OyXUHm3/4CCwt5rUdWTFc2L/IssNOoLl7P+c11wX
F0UM3C7bEZgZA6eCAJdoipxP4fa5M+bnGS2zLkVvAoBWa3nKYRDIXY8WSfjyjYin
BugfjRW2H3un02+hTyNEP7HGzS8pB3vTgqqnKRNV+hVRHvr7X0pleX1d9npgnTZt
OIeIFXKWWPGwCgGcGFrzoqhg9vpcAxfMp4ptwQ3/gAoOw2l8KAZzIxHB/MHLVOTC
ght6TiD12xU3tktOe4hIrTCex1fZALd6Y1RWKFm6wvZxBv/Z2WDZHYr6sg5YKcXz
zwR7MT257ZQMCHQkWNRWTQOFyE7fOG4Rfg7LqhlZoihOI04HyAcemTpRfkPZKnZM
sQ3afNzx9/TvlOuPWtSNV36YKCveUXsaa+NNLQgBvm05iMzCsmQVQgYpPrbi+bMp
6uwdCVo4wZ5jz4RIRoijNA3n0ej3tbLP1wkEo+bL5fd5dBNc0h+BJ/jqM45eN0eq
RmYrtZtiJSOYQ3GhA7tsFx08tYN6uvHvJv9VMRbXZZfwRAbaEm/32q8zu3qGQ3qp
ZlruOsVunbNQBQJsprXUbFieVbaiy0QlfG91mOO6naSd7ZSfA72yfhSXPig0W6UC
9bbSXS/w56FV94X/AHd7j1e8fMul9N8dKdRQa4ngSZ0GPSSdwraCMs5NnRWboTqr
xlrQzWwMN/DIYawrirqpeQh4jckhsdWc30WoQr1oPjuCqKS57HZ+iRU6nXNSYtv1
B/1s0/FDqyngAhCA9FtldWba3CboVnd6wYodp5ur5Jq4HALfODfyZHUxr0qqmzI0
8F/YFTEd9Nqu05zj9r0wEedO+JIIvXHShwAF79hUyv/9xasHN06ssT96i3tl8lkx
un1H1wc3CdVch5Xsw4mCgILQTfH1HXSoDU5eSOwzpou/vxTQx0r6favIREvPeZlQ
OvAev6VUaZfWOcKe/7Kth91lg2Egi74vvDxWsVmF/Pjcc29ZbHMWnP41HQBwUDQ6
EiYxh/LViT4ZkJcrHLIigzSS7P0qa1o2q3FHaV/JXJkqW1wQpvSLRijfh5qa3+BC
MBLTrIblyHwOBhPf1iU1OX8UyJERe0Z3YlB+56M4e38+UeAeH2+5iMRB8j+uPXJ/
Cz9AeEzl17B5riVoz38OKBfQBjDImUam9Kt/Tk9Lc9DdN3uQsW33L+3aL0CDZBPK
QTjnL8f41De7dRm1zdkMlCH0unczZuMWWXPvecjVBr4c6WdGO1c34ShdmmBIelFm
Eq5/QRuRfZxYhQe37EoZozh/76cXnfxaYp5YNsGs6rYXWYYBiJCkUx3WK5P42qha
GXW90AgNKnY20GkMPFOPq6V9tYV9mPnEO85s4AUGHyGTJ4b9x2YgctpNZI5VtcF0
PrKDN9yD1q9Y8mK7JlqPdpJv6EXEezrEuBjzQqSGsS5Cg4Vfndg/5N79vtBx/HmS
cEQ8oJJZEnEo77g1KNqPZiBLuvJwcjYaZZ8TgoFRezEzPRz0CtTdPX0o8dki6SlC
3IDRQiGrkOSu8N18pwkW4z6tHxPHfufKB4B8eNHxayC0rk1UFBmxAuMo1T+154jY
72h5QCKyCiI4FqraaM3XYqacPaLE0FTClKzKbo986Cv1SPq3J6Lo/JnlhKMurhsY
BkB9TsfT0fwXWzPKmpx6hXouT8a/thhGhmHtO9oDPuHcpnJH1FMeJKJJ8m/f5E2m
fRjcvcwqDl4A/nvmhxNXmfL1xOQrmE77adlK1KVFDR5oTlQvzKkaEKMHCdXmlBD1
VG7UksKMnPnC94rDJ+Kvq1tp2pR/7UmgUiH6XG8E6KTY15qkZ6/yukkVmJuqD7ZB
jYu+oXCsvU5ctyJU9l94DRnKRTGT98dxdfdynRSFlGy2Sc813tKXhYMgrzKV2NiL
LCU08BlLrZmiWut6MwbwJGEuooPHaMtUf4XviwdmJ8zSsAn8cyXv/xuFlqyDTPdy
7kYZJjsT9DLG6m1rv5ubMlHM1IfPgVsYrlII24hzyoxTyfwfknmZR8J8IkAS83x2
3XqgGpUWUPCuOGvEN2mv5mi989FQou6LUVHDGzuxNIltMo6gpNpvkpSevR1HQEJE
D0ZuitDNQ/fdLbT5DKn04jm+p8J5bDqvpKHW7ArXFU9bWOq7kSQmKMMO+n9CTlp6
h4kJDDJUKZ6EmJbZaC4bKfpE6vCbb9upXNyon3wnOws7qqNeCGkLbKwXOIUynVep
lOeY85xqWiCAVsvE9npkwVWT7A0WjAS8lCMsCha/aBiSvhM74zk3jXE2pZFktsZA
C1U2ppdhpU854qZrJXAn5e9Bd0z6llkW+uT1U18xXJVOnBYNruznbVXNFQirCFSM
W0/MUFf2RI/PURdbQaGBC3p9T8YbT/SxnrOWtgsmnus8gWmeQY+ArRmahEVn1K5B
2QD1KTYpNK3arIuL5eZCzvK/s6BELrUyxlbylb7Bk/F1Bgaj0d/c207jjzp3mh+t
XTGaSYTscBgg3uN0Va6E8+xIKKWGCP+Fe4LXg5tmmL27odvuSDf1/7foyycYeMS4
0NDwfsWIUuCFhceliIKpH+2K0IFhJFqlvjOiC/ygNozHzgxnsBJ+sX13nnmoyb+r
++DGnX2DbXHozOcDcY2DLAiSTLmrulFGpGpaWBWUe955NjgsAewexRSiRJ/bkodg
9+CoO9Wt58huYMI/8Fhs3YNbPkPuP+xxb1X3PQRnBJcbQWz9mvdzYv3GaiwKhaXx
MFgLyb1deqSZU+iLM1frcqBN/RRPLy7YwU21CSyATV11wpjFIYWEYX9HhHIJxgTl
v7QfAJDV9T4yWe1NmHKS3lpkmB6dbrRV7Hj7kfPMRS8mhXEf3q2M4xqqL0aZzGA6
j7LqYG8z8w+f3F4ysEgxep2qtQoSpfRTGLQBlKjtEGRMPKoft0UjrkDqgDHtYLDt
6mAV4wMzhwggqDF+rn5RBj0/3fJpJzB949dXRjx2LYFhI/iFKxsX81sDRWCXjljt
egxIkZILI/u2vMszua6qXx/wtMU/YOOFCATfYrKpfn6U4oJZSJozbaPJP0a5Xgoz
W0GvDHnA1j8JHe1tFjPzHQyPcs9Lbt4OJSVIHmOSDaMVmJG07UIxVeuuxQrTI2c+
EJP0tvh22gfg0F4ykek00uyWZjawPIa+vQLhYVJEh/CFZ09iLVsqemuBL/C30549
uSttz1/BkxATNWtN9g9D9CuQecB6gOKtT7/sxjC1/Fb/KWgr0Y1r4hASvrpD6x1P
j1G/S7kNPhczmdjjVbwhCeN4n0FzSBAc/Er/7c4524lFSE1rfCpRG2DQJmLI2JtH
FiU0OeyRD3gIVDA+kKCb6xD5LCAZZjiQzmyxYwC90loQ4SdypCB8pI2rrjAsjDS1
RTSsjDV4+wCo1xQqRr+6XtMqMq3v92GRUWMFcyCzrxFubQQ6XOQMx4BllP0wBeFA
IiBTjeo7lNddITc4tfOUX/ktWu+Z9WTY/ERdct1iJp2ZFYgefEcV/uvGZzup5VG+
yA7o4c0LR4Oiwsq9/VZv02bqJ+227oalcXT0+PyaiouuaWt1b+ImsE9Itjzbzs/S
TSQ526X5zM5+oOv8/4DYOo74dPHIcNdbM5LDPX9hOFnNJeUoLB20VdMjTh2+biJV
7jnk03ol42ReC9lJf7QHbYt1vL6+qe6vWDcYj1QNQ4ueoaP+71dfmV1mJjbGfXK/
T1NNhRCnKeBzjkEFCviv7wRTT2mztFrvBS+xBQxWk5dcm5ynksgIya1czxrTNAsK
zuPhWkoGwl3xViEEHta0NavNio2nfwreGWfVyHqhyc1S9bUl1Y/e1XWNMgs0lEPU
DCcc5mqCvLcOgFR+2dyVeGtEfi4MHw1Cs0swdTmNHyn36WC2XEUeYrNHZ6sMkuKm
VGzXAn5qzszbqcG5kGAbL9OtZkqEz2QI+Kl+homsZ1aNlQdMrUmupAwEus8kjm7/
/3xd3W94S5J0Cgp8Bp1PA8dLgvvyaDZjOyJKA8aD6PeFg2tB3H4X+6Eeosqm/5Yc
EKbSg3ohg0/VeWivXJP/GVplnLF05kGxkV+uI0+3o/18l7fz8Lh7+wh4SiD2Lxtz
t3IDFLbGn3gIPzHlyaycsPmT0qqAR9FR+U0sSSkXMs3Cls7kbnv0XZ/+K+Xam2o3
N936Pcc6quMz7J/ixvWl7oCjYqtlzTn9r09Yu8ROJJA+qUrvg5YsNBDaNBjQSOkC
v/r30HcXQgOW+/2SE790RAIJa/6lTPIA530YUknJmw3OAShxAWT26Q5nwyUljKP0
4HDhsNzYlvFw0Wo5ZrbSA/alXTv8N9ZaXbvff/tYA4fuWO+icJrwuCsdiYiZMxfZ
tkcxL+68tukURul/0GStxKFO+54/EWnHdLRH0o365LakvG3+BtWtxJNVJQ9dkORQ
QCXGp1D15SFfF0OUx9XWtf5ZWqNboQctq24D1bnMbB79xn165XMrvBIadifSnndX
wiIKQo5vmoIvVB6pIKhIO3xV2s5xEjllVN2Zw12/oPHUZ4XDIsaei0wKKOsoVgbM
PkVFGjPKdmbTVg9K01D3mi258q2fgD7+WnGdug89dVj/N3JGRt2UirB3q4FnUVe4
VXjMqprgWHPU74HZMOD9QpFCb9o1EclVlxhtx9fn8yAy/PYHphwZ+IKEe6Go1FKD
FAZqxd03jMKRzDFuoDSuHiYGrfvJiZ6IRFwpl1A1hM+2V3H7sRRyqIpM5EFrhk3G
v4+q1+MKyvRKZrJblw5EXxp0gszrlC8Z3GJrUK41qv2DX7ABgIgVe6b7oWnLCm7Q
WbaqhTAU8yfIyBw7Ud0ESd2Z+0ZL8pWoMTBFWv3MhiRXJsxhDLxS7BfPM1tWKhti
zApRhpT3aZXhMCRaKzn4BxJWh1B0PmlMHJ9x42B/47GSJM+opcjgxcn150WsYsNk
vhO7sCzuTwWzy8EXogg4+/XAf8+HnoUt1CG/SzuZ/O7zIqwyjVXNuUhr1AXxGg+S
73ZrxNwThPBIO+SefnLARvPQvoNMBjqa7xfD+FOGPekhP4ew6tAV/Kbbsc0sfvXh
iweuxw83j+7W/1irUMHVqgs90SxAqgk1ZRNPB8ZO/pgB3KW/33td4mQojJw8Nl4H
2Grr20xRx/BJCrTYgN2Fpv1tDGHs7SD8CqGUJ93f3O3Js/fD27ABAciSVk1+rFV0
Kqj/uwq+x7LEnI930XFFkepsryeCdVTLmeE6zqttuALZSSUiWuaFsXRFl4kMF1rk
Mk9uPl8FSPvIL8BqJMZzHmIc7A+41aUo08Eepg+IFBGv7+FPQPzL8RtYgWtOIn+Z
3VvLZwUyfRBdSznCkQtiILy+9FFX/gd+IZQoQ8ysg7iQ+XtiqSJzlhW86buoY7tv
3cWZLs0/Gl7R0OECXOdJOmuimbpxTg/E2x9elHXhO55RwQQfJttejzoBELujritV
NbKQ0L5bLkxDWtZynsIcGJuixU4fkRTLEllOQbuDg0Qp+7LxCRMQJ6TpIUmboqxi
asPUghqso4MBiW+syI+ObuAOLRrD2noI8E1NU+Q028galJF1y73hGWd/bDj/tD/6
hv2oSYI0yyKB60zbI5bNbSBiDyfPvYrDz49ZKb15aJxxmGMgo1hro8j8KzcxVCI0
nCPuKq2MoxXDIolDldqbW6InC1vgEADwvi2zeYEO6A88bhFo1b5KXUUF46v//lcp
l3/ZEOLd9B+2mvP5KhO0vImDIdwLhQDCvKK32egH6ne82bG0BxeN4sj5isanJSQk
y7TSpEcaRLPiZ0/zG5nKCLlG1SmKqiwuc2qRtk8BZ0t0XQhjHKJ55PKKqHtDfirM
sXcS9ypveJ41/NfNk1PVgVGi0WRPiz2sj+eI6DFQPr2Il7bRhdjrSA0McGhZlgi+
BjMK4WofnkqRl8iBg20GcK5KmBmCBb+e8GX76iT3R6O2WBPMzLk8PuvHJ1yZUeBE
`pragma protect end_protected
