// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
moSQA9wTMq9axZXALqBs/YD3Z58tmVZ0//B4rPELBX1BxakNa6Hl2o0L1CZFUKTb
POcUZlfbGMiRQY7UucFgqJWT1Mmz1CP74wwEmLpoWAAPV7b604w+z7kdCuyVzXov
TUy9JFt0vfu6GioXBZm/5ktRxQiF6ogxbBH9rl8BAU0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10096)
7DhYXbQxxmKjmBAbz27CpcB1ZxPQC5jsU1rLDE/mazsQgEiAHV9QrDfdzU59jjt6
TQ/bBbdmFcOXQQRy54Ltw/GM4ZGcX3ir3BoSHKEbKtSuC3hnSqt6MtwVuS8wf/Nh
J0siSenoZJOTXnaWYMxc77dnVyYQHBOarDk23UiB+4ij8mLyi/k6Lr7rf7nfKS0u
OH4jwbgezuOmaeiP235Xa7aGn0CTFp2qwYcIq8aSdPBD8E9Qtt7FCygoTrthDPSD
VaFO0ekLnr+fVp1fWpQO5IbLTrBG+7AS7Z/cxxuYhOK5JkHRuA3CviOPhBNJF664
im5mnk6QgQBckswOvu9yJZwqoRNm7yytmMj9IPg9Se5ohf0mgQlqM5nu7A7j8ZJl
UZCqXFOIsw9O9aM0O0WxYMSRZxqhw6i/izoyhVQMnAXoAKsfTvxnUl7NsrFYYLBO
QdmrwdSDupjeWJTW2i/m+vxMciMu/YYYwbsgBcPE+HhOUn+k3pAj6lpgSofjsEii
4vy4JGVJ4AFpv39viliHFaBVa3eoFnpX5qq4z++e3uc6rWHwPCKKBNjczILaVGCT
PYRkVet6qW0ChtRgg/kpCvu7RlqpW1XrwQ2S5Egd73CPbs/jgDus7E1M5eJtkrAl
l13AZwFcrx6mZl09MVtIDcbG52EpjmVNlOnpypvqVAtdXmUEPkH4zXoUn04zFxUI
2A0f4BAbrTjhf3CRlVxZjrww4J/2vb+XllxeNqvcWTVRug18+O87LfIUyO1/IA0F
d+ihm9nJruf6nj+HiPfrgJLxOKwFxtFmPj0JrDn5GSV4WV7L2+tLcwJt/Yx7BSja
GnkWEcb44Cjux8Y3BIz2n6ZjWaIe8m++OdA8aINnJf2AGyqkZBHLLjNmcRaEPN7w
Y8k3Ps+S1Qp41armot3N3n/NCmPNHiVN12ETbshevvznMb9QgMlDGgjZyLK7sjNZ
+zfcPktmbWVAzwZ6SOZEEgNraqEj13nYxslh7UjYbMHg4OXghDNte9h5ptJPXqTe
a2CKL6NOaMC5NveiX+7+IiHYTXH+Y26Bedvceoqjapr9+ujQKa7ORcv2Bnbn66c3
pStdYJ0wQM7mlmmRb1trAOHpDJQYh90NrB7S03/zz5lAX+0/oirnxuRh8qHyFGZR
GSUUojW7zhidtcLmeF4s8HSwL/QvuiYTsMAKPnSbHzNXRyKar8vzdQzlDBqU/7Aj
c3Y+cwof3bJ2YHadqMmWq94Q9wXVG4LtLY6xxQCPUolCHndLHpqYA9Vp5vLhtj1R
nG5hZB+RyWzUruTvzl2KnDxz2hgLfUShZmSqWKy22OQisKaENSs0+K7kTR6a+ltw
zCt4AgeJKmSZxuQAp9osuBy84UKGEPKZwHEZfyb8OhmLCgSn5BJh8yNFIMBy3RQh
sCMzKJxF+53rg9sf+xCJkresS93OBlIJ7AqK0KBN764zlL1uxTaXEsQoHKKgxPIV
0pscGaL4mLoxxWfWSYHi2Ez3kPxBzE+fxOOjI69yVua61nqZHlPm9YQoWbANqRn8
ExyQUjv+hwlE8ZeL7RV3uN5O5WdyWwUe+EiU6A+5a/nX2D+k2dvwLlVfevXW7vAZ
92Y3Hr6sa5OsmL8iqwNSCHOh5DQG4HOZLRPM+/M3nVObSioBywsvtcqsaGdTa3Un
pBJ8dadqbMXOYANiKCMKmZwjbz7SR8eOfxJLQmtnS47HxxM5DHhLloxfE+9mMBN5
Wp1Bf/kaS9mVBEDLacpEXxQta8LQp4AzZEwJucITRNuaas4EvWp8cB44mD8u0y88
lnopHNAcXMnj8Id5hYPRNa4PAXTIR2oMLHiUlrtzkoqbARDS+OvIKJxnIx+iZHfz
/SokfsJKnYJgNQITTqWk2FALkNlZe9w7rWiXenhYR6pk8dmgAMt5E+MSNtQw9B7q
NkPNV7okQ3acnUe2SMvsC2Mho6yyElJK9df0tDsehdvAu6Bg8Yv+mpZOS6VHsZPX
nGn8oZzahgOXzpTobstTBGkEmJusIO+wdvcelyTwybQe+Poq7ZdMZzCE8rVzIvvh
2VERYOcq8sHs89dxbnDdm8UYfGVlPHZrDCacuQgJPhlYtN+XRjsICiXokTKt6pwF
E2NrktfSW8gaLCJKRUShWckRErf2geYk7ChQzMI12yClB7Tue7wOhMVi/UbdHkt0
xrfD9/CDCXPPu/91i3vzWtyhL8xWbxrNzjpEgtbM2omkHKqHGdoA9yoGFr6n+LIG
z7PeBWwbed6HOrjpyfrWK7LhLBxF67d97CRo4JCeIS7L0niBKhlO6D9p/DCwRHxY
qXEzjajkO3IEI8OjYBu5IBQtmsDOTFsVq9V9HBOpokPgFbsIIlVgLIgxH4/TAVBH
m83t2mj3qp/zNPUL7BFhqAmJ0hCm5pmx4REDgFd3IP3rP9KhrQr40BpfOI2wbOGQ
s1ubZvvUxYSUvQuLlzt27q3qy8n9B5R6W2EshpaP4E/dAUuNkJqMHL3YTs+LQtLC
g2TrkoW1e00M6ccGjxP0DkxotvxVnPGhlmqXZInQzXrmVPB1QWN4WCfvVYegSa1X
g7VjeGCSFzD0n1TRcQiwhqG4cvxTBHs7Ht5WBoPMZExF1BfZcBwwu99v62mtznTm
PIBGtsVvXj3DGduwFl6zoTNFftrIBs6QTftnvh3y1usabs2fNyqOKo55TgXsMiUj
D0sO0tgSEbqeLX7Mpxqx2sSAhrDFDszCZgtBfJ44E38B4km7Sm1TUwpJaGld7K7i
uKi/83Dw5MdFgjPeNUHByURvuSCXe7rSIMzACo3J4aGG+E2sQ3k0MC+YrH/PzqUE
xwj95s2zXh9kO6otljUpgdxdmUqjn+YiZpUmKFEvG+gdqQ9djad4UhsQ2wAfl2fR
2AtBSBTWZ/X+ZBCcBlfcb6fXiPX4Fusa3SVG6WOlvgl3tfFjdTBlk7iKONTmtmn4
a7nCejqAsA5/HAnLu5xv4Vox4S8vfGxreb936qkpMdmFbGZmuz44HoMwb6M3nyD8
TaRb4TrH0jgOz1qcEd6/m9Un9pkODcvMOqwL6643qMETaOOwLW09Els+GDEkwEqx
fp3RoR+wRPPDB7fwmL4mELVhgWwVPUr/XIqMMO1j8DA3CIF1VYTMC8RMYng13hTY
Dg7UrnI2MhBqHwheSfKijClYIXZsOZFS33m2eRUfoka+4+CtNix+/XYYJFF6JqDL
vNZYehDof7VvqgbUWYqixzBSdJExjSAMqE9AqEPwQc06icNRq+H4qcnX682lPxq8
xuLAcOy2CV5oVbbiblrSaF5NTdN+4NoX9V11BHUv/DD9OkqFAgIZJeL9P5dNrZK/
peSu9SACIBK5dr69w0EIX/eIBUORzuEM2ai/Eef4FUR6UN+3hIv1xiIN5KZOdaRI
+MHDWcsQS8JJP0ZF0DPFSmbI8hQ3t2luPyHtlFbEOUt2+ndlGBcAqxT7CjA2mg7u
1qLP/Fh3N1KhBVfu4pudhuuqQ97BGaomZZKnZ4T8sxOgut/vD5DvmVybjIq3+O8E
Lk5slgD4HUvUMqC1u0sAJJFE8ZxbG64jDAPfpjJO3Xq4GQ03JBj9lOMB8LRpokpw
0O4+IFD24Wh1OP1Kl7eQnZoSsXHgL8/g+bXjkbszrutCKghz/dx4WTxd8aHGsXPe
naAfAdpYxo3ymd+wxt09z9RFj8onPiSP7Il8bJ2VOETm2wjXicHFouzE+Rb7be2o
Cf0jf9AB+XcaJlWEx4eWycg7212PU410b8O3BJAbD0sXc7K8bTDBWCryJqVya1Xg
R12W9gF5PlbQKnxqxtSd3k8F8DDXBt72W8Bmu0ihYnSzQN8sNa9kdOOdvld7+Gok
gn8QvEqowCMskDWt/CZLFpZevjPPgbVnqJb0JRlmR57gBLXRmgtIsiWgjFf2VbO5
nLyINfBG0i/zh2vGSCkGQD5y1y0hnsfB8DC8jZiGebzmj+FTL7ZuNuPk3f7MSEV3
H6L8XsU/0H+xJUaKOYYNrcZJVoh2EvSP5DF7jp5vO7XyfaQsR+aPUCrLUH1Sz47A
WiwzlmGgeP0uNgAYDplX1+Fnf6kC0oRbkCpELsvVVHg2BQ70/tEaRkw5BVc2Xt6/
osguZX9/Uh3E61rgZiO04wSuQ7rGu9TNc0TjLHHr4c/PFOjK8dRTsNxmuS3g9rSD
938TGIsityby+Hg4E5N1rSsOlmlSv9M4stpKchN8HzRA/l85hROfKsM4FibGVVHW
lcb16FQznVasRXi/TmPV8IaIkXZOstrr6y2tCALTiHb/kXs3qBMqGRAwy/L+0m9P
HewYilMmfwZGNjSaJiP1i62uByb6Xmc66+NMtvo6HHIQ5DDcQKetgP5V6k5Uj+/f
jmx4jXS5DIruzou4ddD81gRvb4v3D1npqoLyMK3ecEyFsr4E1TuBBrDkiAjYIcEv
XdgC9PpNF04u54lNWahdQeWg4vRJl3w0/AjNY2iNIArucqdqqLvhDtef29kTXllI
F7OW1teJX2f+2wNemBMzKtTN3Poj2t1YUkgKmn2GopprSV9pH6jfzT5M+I5VayBW
WR7YkSbI8l1c6YgqbXQycti/uYt1v5K1OHyyjMkrYoOv8BW6ZO6tTUNcgqmsmn+I
NWo3+B5EkWqRjKJwpqHuBc0ioHQyuyS0QGKkC0/onBtbFNGQMsdVh3Fu5sVZV7X/
ZnIaYyY5a+JSw3AYUBoULW9yjmtICOhOD7kVY02Pw/uKCoNGxealkH1v7+FYayR/
I2/frdZyjVAeHjrgkgx2D4iSXQ9s0YtEQveGDpHKQzRLBB91NSluM69J8PQRPUmS
JVbMVJP2nNg0xuY+nNng1BlU0KvtcAwgK3pOeBsHhtJJ/kE0RhuBfMEKCyjpYtYX
haYZTalzzbCssnzf/d5uzAKvl6On9wPF8ZUvTTUvATTII83CD09By4tqPTvP9dxl
4ge0CiQ8EH7o2H9Rcrg+8gqeLhSAIjn5OMf1ND65bdAqWP7DmI+RNTtn793KSXo+
BNSyu1n279zg6euQ+TdGYQoFQE0LCWvFMlPNglMTcoxAWZSJFkJ6g1IEoMAvYaiO
+01gIJIovKmERq7YZn7FZ4YRvPfxQSLSQm0dUgLpXufNEJlZQ4QJywl/yBUddFCL
2qqL/9Y+ArodqTZo3Ktp7y/9BTUcuUvl7Db01I5LGin0tfvo9YLkvaJCDesoM9SE
LMGq/0Qb2peloecyULJ4GHzpIU5mkU5aigZ5EQ1YbIeEKXbj8HuwRR/QZ6PKkwQb
69DMM7SFY4m0Z2+dn68U20lZLxg+9Z+W6U1MS+HWyQDVA0AXwEwIvgeoCHlB8oaT
l+2hl7R0RtV9W3yVWFZS2514ugClATK1AN7FL+kfNmMN1Ey4s4MsC7ABO9/CLG0r
49hA3PAAsLMJGBrKvP7u8v5NAmH1hS3/eIxQS+RcM+GfljBuO3Xq86heEOEEtB44
FtFQENQAq6tRwAJrmO+ycCyynAUHKH2JW1yau7lk44JsxSH4MNKhrFv13uP5Tu/b
BadwjvkkTNlf9/nMpyhgO2lh6gwbUUpmJ4H0mZaadUcd9Ly36hILaez7iC4H1q4P
ogEVs8+VfPXe/grzqj08L2pY0KbOBxpr73M1JevLV43gACEHjQMllhMxkmTOFX82
EBMfyJeJqF/zZi2EyHKd7vJMEVSeLPmMch09UlNfeQT6r2rm6EK2aV3YHvvGTi9h
AxtLzn9ql0/QpAUPREfzRCObOO8cRx+H1aQf4BIlZ+qupubo0JyVdB9OKXjhLW7g
UVZ5X/FmJ7QpBpju1OcNDZ2O6NkibHP5DyWGhlgn4GNY6G+XxJsYKf+tc61BpHhS
s3w1PUH2TcImA/h8oyh5k7rHsfiBozEr/9PHfcWANkqSmt1SEncHHCVnSWfWxAPl
n7cCjPqt03jDUKETH4x9IGm5Pr/aFuzPE3cCY6eNrshewQQ0dZqMVo+w4P+Li+1w
JuByqb5k3nodFxXyG5vThbtzdn5OD0aSf44sQtQMu+gTmASft208KVKcvrgB6AsC
Nt9zXGViJfJB8JaFVp8YyuuGyT3zBhVeLOx64Q9VgG5RuAUhbpSpYitHN2dGsY5Z
2suqoYRjG40+uyelISfL40ezRPNCNY0DgNl8tos/60Bw4O/EiqZkrCWbTCigAcC5
UmVQmvvQzIEYi2UYWDlH1wUUlDqWj32SdlCCXau9M6q0Jhp+fI4LJ1Hci/BeLxtq
gLuVAc2xeY99838IGEkwdG9+8RuMg36ktEZtSVEmO7kSaRC1qth22CsQEvSYHKmz
EfQrAy2kJ0I+ABWo8U1cMzEA3vn7b7Ct1JQGJLxJy0vfdJmHUanu+6aMAsVRG1ld
MyXCyWPDhKk6fMCaH3RiGQU6Avl6ZBYgYCIFjRXPh6nRYjVb6I7Tptb2JS3rfsqj
iBKwIwVpo1XMK+XPZ7ttrA16gyE3wFEzUnnP8HGLp6wgqQxOWxYomSPR1ATl6ZNe
AAdmSylkU/T7aLvh5KaLEUpX5Bo6rCNqbnRV93wat5xC2BU/resjyj57krTXsBNu
gISGIcN79Fdo9VEHc4NlsF9fMNnaxqlxC8UAd2/ySDh4jQClau5t2PthJeWMS79W
Rz3ofLcJm0HCNu7PdlmXrA6r7t15o+UBhxfn/WS+BOv3no3T3ykIXs3+uSNSHqJc
Z0BR2MhuWfPPcE/oyqK15fgHJi8poEnRb7jbh4E7RCVeTbhO2G6bPzO2YaQ6io9A
X9rYhRmVWKfDYrJAbwid6EBsktEBGFDtPA+y75/78Db8yFMMRuuQ95W86vocIcyW
h+34ERn4BkJQUBh2ca7lTnUQMuZljdPt0VKfIfNK1shLtgBedYtJMY3xqn1kRC/w
4qRgiIoPKAq8aTPzmTfJSg0fLFDQsfxxSioXuKvgV5H1TDbHMy/I8nv7jCXZ+AmI
HGxW6WvgjyOWjS6y8WGYiLyAH8YgnEwPfLV1sgvTiGynERfzVOlws/Ltsgj2n8zJ
ovmYX1ujk1WDdFPOI0zAqH6PLh7Wm1xdqZFVe/M5glypMICbwW6rkhGpmvQY0212
6cArnU4BAwU5n+mmvJbw+J7KhQ0L+BsrJOWuCpIEoqbwbwYFlLMKwLPJY+PpADH0
VgdCM2pSauNZ3VybH4LNfVLpt6iOMESn8MYQCBG2JdzKV49cJ4xucnMGBbYV4zBM
C3mw0vGca6YB4MDRXJtKp9SNFURaDlWBHz9nfzOYuIOeIOXG5gmFZ1IhF2rpi4ac
ZmgXv1syFOn67rc7vTjCWNLEU6jqjc3SuqKJk8AQx6ltOkVFv6Y0F9WNA2JeIn4q
LHcPGFCk/pEDc3Dsr/1ERRYuL7SEMGIAyMZmVDNuYyprunFjsbVupjvap8B5sySp
IGRpsd6amvgHmYsjkynQCIaUGf1v8pU3yUVHEAyLPdXW8U/p7k2RUhSIRY4S8MUb
HbF1l4ySnzWUcpkpQnAN/M5hQrN++6HgpS832vMyFn5sp06sWbEH3Va6kmu/41JU
VNMAi9Vx8Egu/ijdyStlPMSlKlo5qOxrema/Vispg7lUw7RpzkMNxmAuETyqstt4
RRNrg/hTbSVuOGXMqCn1kWOEvBJDPEZ5ba3tLj99ZVmJctF6nEuA9FCzEUiXtqMK
OWv0RtujHTkIvHC3EwFizBrB16AX6T/oUVT6Jq/hJ4OzBd/kcTwyssVrF5fm747N
yb2m/5/z4DIg1xPQZFmnFu64XCqBQ3+IIiKrSOkVkkLP1k435G9ia/vFR8yle3Q8
6ncDApYhB0z3JZKbwh/9vLjGVjFcLVGhd7hWA4XBtomaouAxXvZd8oe5dET8uVVN
DIwBZ+91KCvXaIO2yBAulQtKDLC9xSyG20rAHQcZVCV7uduSY8WIlfpENo8bB1Fj
2DMI/WT2PSXhqpLEbznNzQwECHTYm9M3vLviD2RlLf0wpYqVFrAarsnY6G3VA2vl
SsMYUTJ5rqAdmOr38yvGvzq8TN9FciCr2hyeQJROEe5X60ZIWpKRKYB0J5s7Cz7I
gHZ6zJ4igmsSdVYVFg9Pjb6lbHWezNSq6rIF+yLWRJ0SZLMLKcgmlkay2fXXY1nh
VTIVOprNlOG6kXWsJin49eZE1jseLNUM0sOLaHoeN75SZNq2pcQVmYTt9fXn7tJ+
T4hJNeFTwVFOzmM5+gjQdZOpVBOzZnTfxJXw9SreGINvIwG9ItJLm8HqNE0st7+S
sOQTjuIB3JfZK53MdgshnvhPxH/mYPlahRf8YkubSB+ocQ+55sl/RZ7gzRQ22bAD
MbWUqnvPAMH4oTqYEzBi3BPFFzPsjB+oYH4QMPxukuAVNLwU6f/W+FkWIyAzTUsu
RTOvjD58RohWiaFRfDXD6ZmTQsWz6vca8wKbyQKl4DvqESiKVUn0UcngpnnWz1ZX
UWpz/nCH+Ss3mJQl2twDojpy+Q8eBnSJ82lbs5FQxxAnYNKrhz7NVVGAWs9jtJ/4
wcGDYZPNkuzYL3Pt1h6a940ZVgRKyB8GYGMx8kuTsq8C+jogaZdPH/3ud0aJlltp
YdLCZ8Vt+AjE6V46uEZZVLwJVgJxMqXq8LylenwJIkf/tMJ9ugHh2GAaDKa5EIbB
ZjPfJqn8EJMMx3SM/KDRudHkq7Qmw5Yay+RJfCs7Wtwvx9iWdQt/9QyZC3aRvpXe
JtetFd8EnuS4LeUtf6KCmBZwxn1Y8/gKAneT6Q3cR5fzN+Zv/IKmiAksTah68iat
G7zwQGxAW15xyuOdHdo4ZJrztFvuQz5kPXy2wYk6fWhUCgyhb0nSrBFWDEihdGYQ
TFvBdDh25RKTmdJt/5h5622OI/CIUB0aIR/luI/w+wV67BYR1KgRh1cfdpT0baWu
jkL5YQcquBn1FckT2wp/bAiAtXLJDkITmiZABd/OeSTVSfl6ly4+8ZDBysl8o60B
idXjlJjxhHf3wuNrA5JfsWjMRMzSlTOHh1Lvl12PSgkcQ3lgURLgmda2WuDfxDj3
3I2DSqfI9jQl3UZHCf/u/xZBaELf3AOsLW+b/u5IHVupSkIWCKKWVMjhJoEPrn5T
Wvb+g+d57imEpuotnjtJ40AIqdVOuJ8/hpGoJVPZJ3NurZHcf59sMiw0/hTCs18/
TXpWq9qA6xEU5SipTJde62zUKG8q66I6IXABfEu90P6/H8VuKlqPw/wuIpqFvie+
7z30OVt5Di6vrkG0eRXOBDEb3hx852aqXBoU/E49OvlBSyMpStuCt8CbT9Jv7Crg
j2U2iQ4dD8wwvkQ6wdKc08QH/iWhyWmksjNaPl6Gvkr1Fmv/UFqFQrn5u0aEOAYL
aYm+rReg3H/CpcwBfzOK5ax741tP1+lCfdZUNM2dHCX1CAr/m+bl5o56apW7nXKk
tzfcgbYERd3gprqflqER3B5D8+taXBEf03VojVgLpC8pkijo7zHccITld6q7Mg4V
uI9DpJC6BpLQrmAfIxcu6a1kCeNxaD4/Ly33/JnrYpcbKVbSS5mwAE1ICuA6q/Jb
3wI1Sz7q2L9Z8AnH2Ftsl3qbJnI7hecQfdxUKNFIfET/XvgK+u9vY2yNlIF7zPxs
ZwbFXkaUaju5kD8RGcHnjmHN/oq/W6A8BxsxZg8E/w3OvDRk4jf4aQEjK4XBlIf1
H5fsC8CkAwnRFtfhALDrVdLs0HsnAOvuEjgnEnCsCjjldwwUzR+Y/96QQ3LoL0Xo
bQaMcNiTIuDcc6so1nqsCymjz9eAC1MyMrEL+Qn8eMAyZsTYz6oQ/tGGk3Xnto66
pX3j6Wbc/D/I887MkMqihPwmFOlZZhed9hQ9kDR9+BbEi3IgrjyT1no5V5BF0SP5
zIA8wCeLL2HJ5V0VNEtAO7mdXM3ZQaEeKwwbGy/d1VVrXhc1Cv4xPLBCNn3qkK7y
Brf1pZnpRllW9HNk+GikZrZPuHlWq0y9ofJikVKihqJPc8PxbQBHxiMF1VxxYNc4
NnSIIeloowAa4G1FBiCfSGfpLZ1lErqUvCQq7dZpnNCHd1Xt9Gi46jkHolGAaDCA
VLA65osAZsyc9C+PDqJ/JhzmWusotTwrdmF5Km/0lWGmp/23gKvzR8tMsjngwzqJ
XyuMIZWkzm9p6qPJ8v/r4nC7vouFlZfu89OdRBGPOpwo3rFo/7YvM1KQtum8YN9O
/NNMv2uFIOzSwyDbQNERb40mHFNZjnBy6wG3579lf9RlU7ySiM3FBRfIweLyL71M
2FHM0ZDt/uCjqSnoqMXjSu6iN+POXcznojC0RtZbaMs9IMhhyHy47AgGuWwKf1ut
tTB0YwoPD2LitQDT74EfMt3ooDom8H5e1OXHqPFSVfEl8iaYDoP3wn3rM/6l0/vD
b74ZPPUi21BCyy/XSQdwJqX7oSbszb3p8ep3/FamYkzo2pKaBfU0pv8GZCMnifuI
gxJ37YZof0xnw5S3lnHzPVinj7cEBoZcWKIycUOyaEzrkLK9je1NV6z5L695Xv7G
k5U2rS0GscwgbcLiiKU4gE1Rh9W4gcw7qGfbvpeWjBfa5P1yhi74fWH/1uVyQLK3
pVoHeAGI7YHlpTopZCD1qGf7JphY9xfpDECfDnzcROnhOZNP59XASeILM3MZtGCJ
jWLVMRWYyoIW/rr8B4bk6R13EyARSdecM4r1doAkHendCB+JO4zptJhP20I9zhWg
qij66d1CYwpFdTdawBtYKhPrFF/dZl3bTPmBhkJvmwKAQRGUFfrk9A/N9/m/xuTo
8THBtRTFPYDWgSz6rTcWm9dOKWqvcNvWpPYPh5xiQeyMIvbq8khqqbYWXdnb8JSL
lr/QqChb3D90GEMI3PnfCjR+BSnubaL1M88vVlRrfjM1qAvZ9RvOYoMEaLNweVP8
y79Mn53EFc8j/I5gz23l7h3M+c8VfaYOigtHBgwPrFVYMzK1X0tO1cc11C5lW8+6
SCShWAbWV0/4ASeN1rAZz/PJrwesI+8zVhICP4JjSBakJvcOVHSUeNs1CZ3r6mRW
rh1iKw9HeSlDVkWC1uML4/g57i0GQjw1VHrskfrQ+m3lm8+/4E6dF1o/x7XTA/7C
ChjhrOjrGuFvl5z7TQT96UIghz/UaJXa5xr/mfl1M08PJLF3TxzHHHwuDNct16T/
85CjoESRLkqn7RH4i5H9+N2xg2CxRLx5sUhVC/UKii89b0AUWrwloiM50K5gO9p7
nsP2sQ7Ph0Q/TlUwZGrg/PXWW/xH8p5G50T9dqZE4s7yJCTDscS7KVYQz61nxuTj
VUtXdPeVCAI/1x1oEA0BpdgauYHQB716BvG0u4ugVhqoHx7ORh53GiUPVMZP/O7v
eSeGCrmtYnmYUADypMzRbzphD3KT9iSLYbNzZh7oFHrWFl9mqS7IT11FCotCTrQn
ShO2VHOfYlV9OezbVkNpKNgs6DWLlHJDpIxkJx/J+2xcW/iMWrUrzKcXykKo/I3F
m8U6BqkJjhyRB/3lhoxt12+GGyTO8KLP//H2mSaNBWBPZYTAVGnlFXQS1y6V+P6C
Oc+2fdNZRlPEcayQV2QUQnckl1yM+5nH7jQBY2YTaUGFQwRa6BcFDmatVCWLziZh
KxLVcYG6q7gYms6snySMYBbUha6FDajoXF7edT4BJQ6fpOYlRikkAGwKT6Tp7gtY
PYTXuNFJ5yQ2yM7l0Vg1broTaDuusvhaDLlF3FNxpUayn0ppZHEmrg10d3qQanwi
/85mKXG9nQeqbhEoJe5ArFs0ObBLJRtB07TXDhPvkc5+bUZ5i5/e9rC5HTl0NoIg
q5rAKw6Oi9PbN3bk1UeGUOdFviZ3eNc1YPwbLWoQ6tgNaEfi9voOagWnMGJ8jqyY
2sbjsuBuI68UOdW8Xx8q8YhZ6XXJN8GlcKqyBvsgFDK23Jy5I0GvFZ37Pc8v4tXs
8oPf1byuE9HHcOXS3UC+cXK0iMSU5FF8OB+Ff3A36XkAJdxbc0Oxab18vcxfMrGL
MQABbyturHSnmLbkpX1IAtqr1p5WAl1aEpN+FlgKpNRlWy1WOCpG0C6h0t3w2Oib
vUX5HrSbIudby5VoRxvvDwyEiezhpwNNDWM5xfow3itWdw1d8jeKHn4eQrfyosAn
BcV2+BQeWxfV9KtNHLTgUhyQhteSyDTRnj0T70J4LVLzg1Whqx9Ez5+8d8g2f3+9
URKyRKeptm3mbI9XxTmClY+K6rB3d30dmTNaVXSfHuRe11uPaqGcI1KkmyacbUNK
KmiveUNRhwmxAuDvyRFwBPCkrOf0S8a9ootGXIeUtJC8Z1TyEstc1pLabp/X1B+a
shXvDU1J/y2rmb7WWIe4pVuWxOJjSanWfpgcXNqxbpX0Wr/85k62p6nuGG5TYJjl
rCMxjobcmDgLCik6eMJuxK7acnSjUkzEZVUy1yoUQKqt9jCGRDh7xQ+2hkgYGmcZ
iyjblujIjTWCr52gB3mx1lMnO5Qgs943pX297eiH3tklBuMxuALZ0Ipu1GkF//Sr
FpSTIct+2Ey0uuI1JqFlzi8a0/dSSMt5P5baqTG8ZDy6mhDANhtm3plG7TjyAco9
qmZuwBPnW4aiRg7s+Wi+2UrFgGBbbBghKtMFD2P9o4Mm+Se6WNqinRMgKSdR1usR
StbFDArp+BYg5SBkTneWUwONX7rFUTiPxpyv5TKPXSRFiUxeY9SJqCP8PuWt0o7Q
Mn8IV1pyulNEwEB0Vra47OXvgVcOPB4mM0Cod+UKouKOQEy8fN6D91KnMLg4KmlG
ZcVEFWida0o3LWlqzXsexeP88lp4DdDHtJjB62i3lqidUnIdocnFco+PjDRo3rcL
KoerM/Fb14AwAq/QKuGgN3L7Ab+mghvD4J1r6vBW5aWTyyN/o1n176y3D+fC+S1+
1aLEkxA89yxIPCujq22n24H1wt7K9w+guSxtZqBLNdzKla0hztG4/0PKrY9I25Xb
/YGPf+27bX1mXJZ5TZ3CNyLPnwDRc6oO1dY0N5AowKJooQXCstYBhOhHT8zLlIVJ
aMEL331NBiW3F6YyryXMehQCOk7jcLj/bjrElGWiuqMnSjOpFdy2oEFaWeG/Dond
6+mOQhTVafGa6yZ0ylBEPY76/aKBvl2/YH3u+Gn/WT3TDU/KLvbFJDKYLsuv6Pvr
tOWGdmx+vOcEPGYcNbwelGQ9rYD4mkmg0Beltzw15j6ZeDeSaNviGm+mbiz/6SoV
wBJKVhudrMjWs4CSBIyuP0DmjRq4Apzfx4jjDWBlQ4nUyV5jk7yNbZUiEbwrMw+h
qmwOEaF8fA2gETWiQbXbMwhxGgoF67ERnJauI23lKWXiP15/DumRDGtctALDlhgS
DoLMNaiLxoP/GOfF8Jjhssl8i9S3BZJaR5TJJRmjy/IRjZ7V8Ehy+URfB9OgWbVN
hzD7l4V52JhWrYDOzCDAdc4cYzWXeo0bC7MaWNpnVBPvBQqpYuvbls+tsmjcOZ3J
TB9se71vbvtZyN+Fng8GsOiVuRCDoZhTDMr3p/khsE3BvHr7iygq58U8ci57JHnV
UtscGeer9tRISjesaJPHLg==
`pragma protect end_protected
