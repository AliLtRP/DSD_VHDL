// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:46 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YQfSUYfiIQ9pwlNAs/yhJWHIXefQOBUnWmZZvuCjDYSve9fc0sSpnTKDqHBn3cRQ
J4pxYVyxQvw6gCBz6MzS/34tcuei5TP9AukvV1njXYZ96Y8MtHRjNKgY8o39SIwK
PLyF2qpXg7XOTX+7k+hOEjSexgrNOq2OwjoDpSqvQuY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6448)
iepkSyrmLsMFawcW5OPQQ6FynfH9YfTj34WMF5nUMw4wICcOSl8zAdNGtuUVAT9i
M+KHUri6269FJg/QT3xHpV85CRNfhKscPdN6Rk6QqzMubzsMaUO1VFw+fyPYZHy1
8IW18S1zbac8RZL636XkwMGiOh2kuKIfXIZPHMcisGgV+8KhT6c8RhB+0Riyq/An
scAS2Rxl/XSj2QbZvztpDPi2rmWuMOaKNB6tONY3JmltA37yIQTHUG0M8U7QZTsn
X1/aqlaH2rv4GGYyn6RqA7tGZQGaQmj04R/hwNi7SAnqoRheMTfJIM/47wya7vBV
31E6M1LajUL8dMXtX3Xtn7qPqucPctqxXNXkul9asEAv6HS9jvLjaEJh/AmJrqYz
+xLsDtDkEJAbViZZyV4KjMUKqx3gw08DKkQafdL3Yvh16T1ju1V7HizcLQElzaom
lyQvM+rzekKhhelMTZFxKILGNODwKwQbundECfSE/u8OL1Rcxb+qg4SQZbQT4/FV
dGLj4VVYnTEzYW4MLSkFzmFbxqECEM/oRqrop/XPJoaCwBzyPdLb26hmIqMHdK7O
x9Na9O43oHeU9rjRTs5Bhd6FolhvwWYHwdwkhsM1ie0j4B2I3TC5BNGAJrclXz74
md+gw8rUq7f+Uo1mtfl/UYIhYZ62DYtATVl8tBH75TJ8szftrNpegG+la9mw3bSi
eAqnMXIrZinWj/B5gResG80THRG/g64pE1utSc/t15AH5E/FSMIiyOIKN3JTATWW
ErB3ys7m0rAWnMetVYld+cb5uVeRRwvibq1OZOYylx3ykhXAZqncIGS02C6RqCPH
05AUvjE4BjW/Oaj6yvIp8pDEKkm9kjw1/Ni/74v7gg2bosmETAPaMgZrQvNzOmcA
MeLM7fCXo9Viqki/9DMm7Q/x89bKqYaFZiKvfMxLC8w13OYiTmStrLzyJ1ICjX2x
AafODgtKqR7k3s87o97WRds/U7wZuGTT5dZOwXhHgM7OypZSuYu1zS+EKhRfyRvP
fCIuPlgMBSoMsBK2TqE7joITgh8vnWFAAw2BR6TV+GK1EbjXBSFX8nKygFGIQXKv
e118FjNjcouhpoE6qirYWzyCaZZ9y7uoLauOV7hV3dDX3AeDIMUWBaK6lEuZqKYN
uDh3zRCgQ1li1q8gJItdqCwdiT7hZ2I2TTqL46mlUw1SZfWg8ua7S/urJtJ1hHLh
CuzYIaeiHzRDaI+jdLgEAhErjMr6m10SkvtRud5vgbhZx1emYI43yzqnAtZBbT7L
frals+VwV00OruJni91CFgcUV4sFy4zmashex5dRuhuPnon1uLYKEES4VNk2j3Pr
hevxrhTbsVhuK34TKb7FaO06NCcn90BT7I95Uex8MUbsW6XfHttIc0qRlNYylCCM
bpmXVddxa/WlnkZ8/Ho+ftTPUpkp3s0yO5spEKwhcRijExV5MZYzJE7cqtAfQHA4
MDzs8JqtZxcgKyBqIqzTJjv26igK/yJc9rQRgW6+1wEcs/181QaIm4hjVvFCrY+S
lxyF3ax+IcQASBg/fdS64zbeDh95GRBelpyhuQlc9Q3CDy0KAFA/FmHYcChAXv2Y
2Lc/1FMOdxjF+61hih8qS3PmLoSI/JPKGs4lW3RhCp1d5P0iH09cneP7So5vr0Vf
oPJgIG/9IA3uRTZjIfxGWCp1QqmWHFXexJ1r7pQOjMaMHoNS+7D5S9jC3jkSeHDc
ALgNdpcZBF1pe1GGFNgDkUAMJ5j1r1QMW4ROPd+dkTIVsmpDnzHHbXEtFKlr8ard
D3RyJcePpo5RGGGz0aH6gpiSiQz7EUaveGAJfnT+Zwjf8R7nQ/AHI+oWrPuOvzo4
Agi/jptuy/zJ0M+A0jNDW2kl1yXT/Hz+FKzKd5MFfCLX1SZmjz17+KfnADHVZDfB
XppwZlVzOJWkuo+NJWQpEZ1TwjJ8I0+BYbPaDmHvUakykQzv2Wo/bvB0l6J/PYqb
BZJMBS6AjMUSym83NZei3napMHrYBjgz6x4r9tzzEPQxLaVInsRN7LSLjka+JtHp
iQ7ZG4NX5oA+mIqrnYv4aOQlqO5+pAObZAyDTOQm+QNuF829FXF+S/1wWx3aJgPa
RvUJEjhhLcnGddIdgYRzg/ivHrfGc1RLKCt8AAiHdqEQ8xY8lR6YEZYWubTcCQrq
akGIYTPKXEJgU3uPzi6fCrilIhOH43dKwzYFcMzN+tk7PsTeE2cQ85LvAsFL7h4d
mOII0LMlHbZd8qiN9MJutQHYeQ/6UDq1pGea82TTUNQQ+BbR8jlw5jcI4qvU5X6g
vFR0xyK5mzqN5ogB1VSbHLx9Kv6Y8cIBqtT5xHUTWE3NbAF/S81OkU4M3Ax0/Or9
6xn9PhDx7m6j6rltdiGw+cV2J7inqMfyPmjuXx98tCu5EnXYjKhRffjCbRK3+rIx
yAwqrhw8i+U/cpaWOazqGh9UJ3R5bLIMhtBdf41s1TLYV64Defj9T0suaEVYFci3
qSRhuxPZOV2bL5vjEgmPm+B14D6SoOB6+Vbi/VZC0wBUQTVRi5ESq9vjv9USoQw8
GS8Fn+EhT6jBvqZBWuXoRDL+0u8OCJk7uNKTaBwHBQhwPYXGGFtkTzptzFi6cSI7
QP7pLnNU60VX1/uigk8yQS7S5pFute8cRtvvwdYFxKEcMmQp5kEqgGKMS1X72rY7
Lg/tG0mprq1P4XZ/uDd9+PX+1omrMr/UGjVQ0ww/mxi1gwl1z7vvRZYrN1L1tddu
rUWFrTx+D1WMTHMYd9NU0uLLBzYtN9qtUK/gnzWIb13k1vY1g9tvJ/JIDcHEDX6i
hx3G4yNxANv39DBiPlNDE97iuTkijxINGyeq1GisSAhUWZ/0+UNdMtHNKjdmCrWO
xkdIrg6BoC2AFCGg4fAPKeDa87nOQP/XJDhz4OVkHlXDxoWCZViqHS8+6o3Hfmuj
grh4n+iOhFSQhh0HpdfCk0pp/lHvzePwsfs/TSWaqFaQP87QO4i2ednNfziZ0y6f
dOY9hM+i79lZQcutpBEclubYw6kSGGHj5OyHTFby7SsoBFUNY0Uw7waui1nWm5/n
sonQy5il64QdWSS/z0iL0nlNCub+HIE8lqzO+G5qoucpwPwr/GAhuvroWe5mGl5D
gY6F1xOBETC01EuPfptTsuGYPVRTrO/n4EINjCkSkpaMVtnofX/vQXZCH2aSuwoX
LInqzJm8YgiPyxwFSWmDRAnSu83JfEcDHRVaIv0fBPKh4NmotpPToyrnVrIpPcM0
eVa+5I1fsuLySxl3tyalhb+Dv63w+nDO0XtNk7OUkhOFKsGbyr2LybxWPojawjHi
vJ/ki8mLrvvsLV/TWxoqUGlZDFgCCp8LGLDcjbYHzrPtP1y02OkyLyfeeG2/76Tv
1OlVih6a+So1jitoHE5eJe9X9frxJ8s6fPf359oNAyzFpdDAla88ME61lEPiELvA
4pKKP1zvOmyFuPlqq9qySldSKNaMRLNXCWodbuG7HTIiiv2viHL8sSAjkaOa+G5J
sgUvitHp/WFTIVSi5BW2xDRKzcPBnH5hK93aAIjlv14gZsPOmI5c0FdaWM2V1vWb
KgSsJxSDuLcU/nI9/Awfr89EMuT6uzfsNgUQYiKjvivChLPbd56kaq/3MFDEGOg2
IxnW8pRSRd1WCccY2CDZWnLXxRKjg+HhJe5Xt2rYG8IrYuPOor8v8SsumyE7zHAM
B0isP79rnIWMBYySIMd1v1Y2CumC4IA3bzN2DBG6ttmuXIfSFoYEV+24zPmJ9ni0
EeJUD+Nhl4NEqhWew/S9sLAIQYlTi0lb9G8ewXnZrO8iqPl9do/BZhaw45hbTkAw
zBasYBCwAncIDNPMGmG2FPzeZ0p1u5LtUhJ5PwZ/htnOKpfFz54KoLmjC4Fo8OAC
DQBSCYFC/qrXMuHTBtfvn/WiMP7IjhJe3EcNDvwo+fPtyLCVqJ4jTLWfUPZlJFwd
sGRaq5Ql/juqgq+s7RV9YDb6DLXkvYv0SkwrriHOoO+i9ExIbEd1QFJI0+Vxe7Yg
XF7R5RLuyMl34AXxOKNv+WQYMIojzlLMcppnDLBPlBbITk3owRnFKmDwelH8akG5
nQAHS3xwz1FssLHyJdIxetb4WkqVQbCEmMGfjMcGyc234DZfzZesEvUzlXSe4Ehe
n6LYxLa7Z/MWZqbWNlGibhhck1t5JWRzctAuRyNj/hIyKOpbnxuu1AT4+CGiH9pH
/vk8IDL7ePxq9qUaN5Je0qaeT+FBOpyUBfqt3IfCFThzX+2mdu7ilmYl1Xon0l62
NN98uYkhN9y/XxAEFavoaw5h3ssoplHieR/hMmGsYvwrbKDLNBqF4RiETMi0m/dD
MO1aVV1T9BACdOhih2rkv0LasCB2s2ii2AkCRNbKCj8JP+wvRVDa/W3j7Hme7Jrb
xp/JNriQegNHM6+Inqe5SSgWku+Vg56prBzVnz/t+pOudt88C+ZAr/ctMPhJOADV
8fRFC2InmDgjAX0qQFVF1dBxhUuAT8TNuO5wGbGtoWGtaIz+n/xu3GORzMWkCaQt
XipeyTeJJUSvFtCCKbWbJtJoKu7T8xraBEU9TMK4VZ9d7uufHMVa7TA7F87/YO9E
p4iruqM9qYBl/Q9G5DTK43X2X351D5X0vby+W1YPVVh5fpQP4AKsHx6NKNOt5FF5
+TPU1mATnH0yHET6yxEuJ2Ud7dAUcW2CaHKGdCVtM4+jcb0wb9AdLFZzRyjVXJzL
U+vJMJ2Tv3eGx8S2kdQ+5rYVRUAGt9O9fxakNsat8W75QGKc3+VkH2W/Fv33bhGZ
dtgshryVWTKKa9P44OaJe5TvWjOYKi6j0SFx//nyaNqoppaNnmxIsqrYfavNJxUD
+pQbRhZ6/ejJ9ca0QcqqgucylMCHa0nQMigLnX4RfnS43S1Sr1QRYhMZAcdmWac3
tWv+7g59h86gsRfvVgpsQkc1C55tBKSIq2eK0vPoWnh6D38Esmud7ccZUdEVMMPk
E0KvaCCD5EZB7psP6tjwU1JBd5QBtpJcYysSaM4N5WSbRpbYGAy7uRs5sKtEmHuX
YXl+yPZR54q4/jsEcMjy+aQYM2IuYzdiGQrI4CoIh1etkX78uqLKo+38zrcm6G6V
cn/nEBZBUr6xMx3uAU032wqqwol+H/PefYLtX1c2jeDUYOqwO3L2FEYH4qie7dZb
Qn+bhPxJ+m7t23kI0nbtkt4HiyAT5G4+18vCBJGMWVE9qUuJw8lQ/g0ER2aE9GwP
lP5Nh2CDFl2G3Z8gIs+HK/vzYhaluIOULzPA2oYYbNISKVM6fnV+iQJL3AAeyrod
a4V+6SfSsxaHMMwjcMz4eCWHI1wkXG2VRROUJ4u5yu6ALUfP7qsuB3h3/K2K9Qrr
AkZGwdGoKHfdywYWm/jELEargHzR8awJdSei+Dh3Lc5F4TcyNDcZBH6HZDhzK0ZK
aa3xIZXhsnSRcZ89GSg4hOcID70uc7eS3PstSPfN1wUom2nDVI6qb23eKPfIVFoN
YQmTp/xwcLmLpf4VhKJh5uhRc9qgXOG63EImWc625a5EEmDgibkJ2XH8Jwj+OtCG
L80DT/coFRCy3J+rHSDwla7kahizVrcLUOV9yZVcOqsFDLTcUSblgBIp7mfgE7sr
NxW4n5ObsXLBwgmKX87XOe/eNWLuRK0xDdKcY3M6qHj0klgLRaUv3gXwDGEJ97qq
RYjx4EXbiIuYFR6xbJRpgLfaQBJSvLs0VVJpdK/xrI6jaWen8NwynPw2R7AnJYj7
4m3MnPEK1n8C9mbjqgyTHW3daW7VKbV3QRAwY11J5Jhlebk5P3/PueUR88AIW4J8
mqiLgCEstifwp5kDj96j5IW5fi+ZUmXVXKm7Gz2jAmuxQpTzzk5OBDisJNypahKt
yo65axT9q9hezdLUDgMTE85SRL169pNOSxX2A/SMVggJ7O4NuQNaAwbakwoLsjc3
6wm9aVooHiXdtqOCKFH2RuA6k0iwzZ4SAqltVcsFGheVzFunisZyMTQA2XK8U2Zh
i/qiIocOATvB0gY3KIcBfL7NwsBbxIgpOn1isy1Sj7AzmvSVoidx0IrVvSHwQPJv
1csQwLmAn9ff55PmlDn9YbFFp0yJcZFNxkUtzo4RO/FFKK3rtkUrk1ISi29G9ssg
cNtiC9wU8+QrNu+ad4yLHvD+ldLVo4JUqOWCG/87WE6+GoOCFzzcr3QMborqd2nH
oStRAKB98COR965TwlCgkuQW6dzwX264psL7iHF6iW+6e3hqAJ35SoaHPwZ8EGqz
9q/PgAmKoG1OkRQquHplwnEbHQiT9a8Iv/Xk9NKaU0GuZivqSM0t5egrXHHIcHl9
bwqWTBmJjEWamm630qrAjDxidPgrh7GVgMgDbTwbZKdbishI23KmpHYU2KW/A6po
lomGmW5s5Lp4D7O6/Wxu9aBZMA90MW1GA5pyqU8feZmqFP4rLzV+N21owQyOVZD0
aKxNE6vkR+Uk6cZPc4pGSn50ou9CLaLqX6MBMagwHBLa64K6op84rLhbp+2TBUsd
yap+/cARuZfJPRmvWeStdKgIT9RpGLV17rOt/6qagA1PhC3zb09hmAxMLLfYw5JU
/Gd4JAPOs/eeZU3hjEXZ79efx5y4MDnsWWnsOjZCZ8Curr/PRfNvKXcE+UzHlZ8N
unJ/kCw7cf5AhS0LFzQ8lrF4OkJZPB4ktSxCG16EH7K8zoD5n7H1966lxbMrQ1RD
lyadq+hU98sSyoxLCbP3hce/SwHJmre0tPpp8czBI686/eTJHgHt/HC9/tEVZGxJ
0vF//OstVv/o+MaR4ajbRzg5Dwyym9OToOaiJzTWNs7NvvotGf/T8iCJxhnxG8HG
2tU7BfIVcV7x0bxeerFawNWenw6AI+p81TpQj7gZLHib3YIJvpyIoOKOqfeLrK5a
ZwJLXqKCi3g8uc1BBfYuWLxAeZ3+PEuOr1dmZkPk1C3kBZxmdE13F6THvD/6fcPT
VH+WsXxgUN4pt5OuTsrahJgijIic+K3pfyNb/nRYJQlYyhMOXIvzdrol3WV0yRrz
Mu/qZCEt0S0lSp+BMtsV412Fq++P+sh7Y9bMwzUY+z5cwVj5bTJiBw+Sn9FlcZW1
sYyyymhL1DWj6JSm/pusgECSh9+znBhFNCP6yLF/T59zhXBPu53NVNZMaHN0cIfZ
UWXr8j7+3jH14rqgATB+PH/m35vYEN7hmcUCVM3ri3C0Njyti7DL2vzu8S5+FhNY
li/HN2qRB906AWzx5pV/9Jc5GX83Y3FOIBDHwEyRfFBxTifi7VRBDJq37ofS9SyJ
/u+C6HpavUZl1qYA3+MDqYDCAmLbXSXjwC+pj1n5Vw/g8nAZIMo7TF6WZMzTUeNc
EDGKEW9tAhxVRVXvk4ynLIJMeLEhggYAXtjHk4fT2rQTpXNj8mXQ0iwNMH+/0ke1
xWTDqQbvBcSApnIfnwXXk4nMVRikpBgAeWuPnWWSXd6PVJ6eAjzwcbE1U6rI6BJ9
viFagYh6vZLfGw24BtGEbEdCoaqgjoJtEuhSI8ab6rYNMknnepv+8rqMGmavHybX
/6ZKsKcfTfdb6xUYSJV3Y2RhA7pWE5/rwkzUx1rQ+75RxolD0NuwVm8BbpCr61S7
wYYeZ7bBABGNRAPceEhor5bue0XPRdnFkAvKTbwOnAlN0hoTpvUhTP+obRMko2by
wl6m2/Zxxgo7yHvhD8pe+BehFrp3mF4rRxGNoHY5W5tpiF+Z6MH/qMidPc+fQfQV
lGCakB1PBey3HZpHb8+FoasgovYm6y41ug99KZ9tZojJjNw0/INU74xHnzSOiIWD
GClDxMCsn2g0BUIW4/ktooxw+5AhhP/Ma6LF1FUI7fmXVC+bfIFKD4wpoQ5FhSmR
NSBYBK/eIWOpwlBXQ0e8lnnB1RAGfxwRLT2xzK3z0QMU6QKtQlh/zodQy6RFGmJE
1TRQIQrpgp7y4vToxZegicnjyqKWMOrLrntCfl+7ZqrlU3Dgp+U/61dJkrj/aXIT
U8dgQ1j6EWgqqtT6Ci7iNtu3q09H8BkGDoC+sEwrXWy0wnEiHqHOJzgdPEU02D2+
zQposmIBnW09+ULTrH2uRacO8bKuWFNEzSdka71HxdbKc0kfBy8+Dl2ierasN4PI
+Sc9xbPJWxF9+cPxS4a+FFMI4OzCl5XP6S0BPrMgBoR55mOlnoo5R5TqoGK8omMe
mbBmJn8HaGaAeZlb/UQS/9HEJCorzmNnwyi9ySEY9VvMhtXpaBUdnCRXcnvKOYtD
g4hZbWAp876BelCVArebAe2wmCrJKXKZNcNEWnym9ZnWoVPOot5GTr62e/LRu8PY
EMaxNxuTBq5vfotnQVAHSmM8yK569ogm8UmCi5iTzVKuLE9o9gVXuzzQE42G9Hw0
Vp4iAHmHg47EspRN5G8eKgQAu1VDb0ncjvn9HmG3jAx5dzqqm8Kec+NHN1e8z+2t
L/QyaKTvra6ztxw0a9sghNl35mXPnruLONwNtT9Ol8E2EWWA2l2yxhQ8F4n5QKur
uRzA8jdNq0raOdGLqJzdEnGh5UbsxF2GU7ocukgYYuqRd6d4qiTz23pmNQK2pHm3
P87yyTGRT1owoQEnfTZ/tg==
`pragma protect end_protected
