// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
m8y84QvAb9pxOjMqCLDWUlezWVqAzVWBSAsW7qV8uPwkHznucVAeh9Z/y9nlYdTTzy74045s+R/3
KlxO5ZLP6wVDbW91MATC/z18Fkzy+XwII2zVi4u1ymbkNuQS+RfAgy1A+4eHnn2hOkDhEa6zEcw0
7uOS/bVvcsAZE5lU8i7eSDyHdr6kIjkSwLweBozyJWs+pkhY8qRmwGNd2e6vzQJ0w4bKg0d9ZUUY
vAfMvsIXmE2g0gN9LGhXLgSNkA2XMcknKcuBt5t6o3iEzWtX87j5Qi4AEttdsqTZhz3P0urpTnfX
ndJZCzXYzF0aAjTND6vvR7Wt022BVovB3AgzpQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
z1KAIV5Zj/l4yxpfv0A6F7zVNXY33MrBGyOYZuL5pt1Ob4/uT37A3w2wAVpVRSGf5xRrJ/0s6GZ+
fJlSLTjQbf2XAb3MmJDIkzAKtaDDqKgE4AbV3Xdw6i3nKicyJ5spzREqd4sWckEUuJG/piIDN+VX
KSmv16UqX+8Yw9jcbfNux8Ei0jzV8IC+Nmq3STzvXB94M72/ul71JlWHIHs/V5O3qK08qzcteTHw
ClLXhzbryLIpgGb/4ZNFKRF5q2Ys9lUQyHP0GMxvRedKxI/U2FsmbJ0s0HQ24cmKs9Zob4WjUhCJ
q8NJ+DahlG81nrQZNpkYH8R7iogxXIJ/K+3m/PwcZDe76cm+VplxISiSclMxsiOHZRiolAUmVMTJ
+4YxmMXRebS0fJM7WmMcK+k967iXjsMTpYFZ23YjHAh3TeY+1z/zjdRg+Vm4OehBTiOLQMND9I+P
yf6DxfarfSucSG3wjB7xtWNdYrNVg0PwqP7zZdtNBaRs0GYWkFXiuToO7G7tw3mP51Toi+5L7MtW
05nVX02Rsax0xzapD14b12s03MpuwFm+WLPZZ7tZNDq5j//rnRZl3+snRgsoUs0GE6uevWBNP5eU
XrhUhH8QqJDQfjt3TYf9o6bvSlOw16hgzrEahbShhng5uj3Z0gnf3/Gt4eqRrpiECj3cl5oBDG0v
UwieZ0I37MaWtk+qYE7q1K3rTN4w0Y1UbazsFQ5q3eREEshizosedi1ITeEKOspwE32CZ+1q1KuK
gd9Yei35hVIRZ4CmygddDAqeopfd08Gp7i31l1JnqfAiqBdRvVLRAIY+eHrDu74dciN5mk4GXF/M
qD8AOADHP0wyDRwvz/6+kEPuFixkkyHLyek+/66RT8ruMOQ9Ye0L6z2z1QHrAFeTK4QUwxQCAqcb
F/6wnDBPBp/MNCsFPorj1GmqngquxTLROSeJfpRQrMmmanOJHd3mVoQTYq8LDRgiy8zJXU7R/aTX
GiPOTz4xSiF0BcTSDOa/Wzc7JUhFUoTf0xl8yBZ33DChvwQt/gxsXxR65zYt78zfZjce5MR4Kxxd
HLPHtR62Yv9TCCqPRQGChUzobHqZvWToZVBR+AGaCTJeHl6Xx0Mr2ciXT1dVe4piL28mKBbbc7Dw
grX/ilKQOThYK9cdyT/iHoK93CZyQapu4YZI4zxx+bMs+JkCNfUC9Q4JSnl1vE7WESpKMfrzoDUb
qb93mJKRzupAyiOH5P5nw7XQOJy2eUBrasPaZTf5uJRNLTYwkshSlMY1CVJFH8Alz1hy2R+2Yijy
71TCZH45ZhUKTESihA2Hv3XXIfFoPVhh7SfRNUhiHzR3kHIwQv+GIAnUY0rRgHk8s3oRfeOx1CLv
7VlflcyFpBhHIoiXr/8R/8igXriuf5EWHUaQhs/fH1SxnGSVPRDEjsZbebRomzDLvVlHyp3Idb4l
PAzCXRlwHSuViigAQoIdbFKAm0ZnWpwHSmdryxzy+EYBKhCdBNnc+fg/Bb69g5oPJ2AB841T8rIZ
1ok0hEX9g2dZnfkGPJaeFM+NbUSZLSLnngdk1j8Oo1uD6iDL/+rr7aQIyA7l13QUocIGWF/HIbMg
7AcGhlSpLsV/koKkgZxv8Q9PPVwWkLzXeQ/4x0minEARLrfewGF7LCpZdBfIYRVsA0UkGImGXqiS
WDTjs0L8wlTYNGQEs1Gy0uVZgNY+dSOg0S89s6SdPK5rjTZ//snVK44y7s5s1uE2EBgvqdwIydsl
VTO+5borPHt8b+4ek7/mLHtVKb+hsDf4CSIgVocyqu6kz/SlDQ0afsFetZwJf9iY6L/8KuTzcxpS
5IdbKltHga1V82kljVdN8KZ0pBlR356ccdbXUMFENERpWn+2rQggDPQWpBXC38sJ6PV8finow+7L
tmhTVi9Wpa1EYYcZZCQa2dGiIztpNNsjhQJ2NLuHjnjHOkh+/7WjoTeRhXE1XUvLO/9qoZS2hSB2
BQn4AOmkpX4DDJdxz+tr/tZ32ZeNpKiB6v0DAB5sFqyMm21BpnFnIX7j0HZXAA+l2t7pPLwKf3yr
cwYpJeB4ieIkQRA7mREIwnHk3WudE37XW0ACHZTvjj7+HOgyAvEpxj+3bRz/FjB20VbNI1Yzc/zi
A0EbNfqEJYcWrbGFM0fbIshot9uap6ilV4vk8G7zi74hnyZx9NefnU4R91qSDQFe4CvjvqnDZPoF
h6OGGjCDQOuFrw75pziQs08a7kNkBm4eZcAyPBDTUlFakKwFiUqdLSPJH0QxVxBDM3jZG3+YawtR
6LUY4RJu/Sk/LVkLW1MKYdVA064C0tcaI5Inl+kOtjXDZrhd4LdnEWqPUXMbsneDfyB33jUWr06F
IdwL+l8hd0F5iqhGdO9Fxf+nk1Q6TfZPI8NW+2CHVfh9kge9lcITcvkda/8oSbLuVpCnBZpeAea5
xOph/Atc4N1Aa+0604ZY1xEV+qZlEE9HX/nCdETTUKubrSmtK2Gn0+0+tE+1Oh5VOmr+4Ewg/N6c
zJXlyBSVt4z+E+D3A9F11mZjiuVeHceKFoV0ZRyAUXSG0Xsh+Ic6KOoNY9MT25zIpaAW5ZE0uixu
wq39Hqyp0OYIgJPN7Q4aJZiRuQmI1g4MmEGG4EwDQGVnhxij5IXDjBLXqfVeVEcTa8rR01qvqME/
N97RqpN6XvJhb4cwe8VIEF2bo4AWV+7lRxHNAnuf68I/Tj93jypVjU0mhGBE1bFp/Q+Av1w81rjH
KkcxB6NH7meLOMrTB1Gc4PwDIWKjad1pWMh1FtkBIB6kCod0lUwXZpy+MIPH72k670rKnr6LZHL9
J8FbNGZJRQQOH17FdRkMJiHWirQgAbxH+fZtBgDcfz1lSrVznd0CumdNRnAp8wo6wEMh3zS6GSb6
CK9CgTQ6StlvswSFqPNl7UxCXTTchH3JWkukFzV+/XvCWZxvjrGhCNWCOOTaAFtonTYfH2ii6yPQ
+kqMwiax1qCRT8pcThE11PQG+ziadRo6jHHUxZ0Hd/YOa8kyxC6vrVmVsEn1NQW7qTfGWwmWU0pr
KAhEFjU3eK7Qm0EM68KWm9k2OSlogYX17pvow1nM3O0HMYmf83suNH+Ugj/g+UHeZVyAxSMnxk0Y
gkV0BF/9SnsQiGilK7kAyVxKosf+wyOViD8jV0HC5d9LWaB5Ze6VJTjRjFzawqHSMT5yNijKNGQU
Ad3mp64htls3lN+5scMkiFMF6GFMnYCCtInai3FJESjIGP2sCx86UBIZT2gRSWseIYDakbmI7iQb
2NXDBshHqmgKo3SzTX/dCbO663zBvDgSyCoMrsUjIn+RL3F7zHESJCW4eJgC/RExEkJjK1zmVgyH
PCu70BTykm27AR9fwW9C+V9dOSyL58nJi72RW/wCBrc7f/2IgUoK6YOG9kKK6FWKo9hxPAQulox4
8lPCOl+j7cb405gCGW6WwlzbUR/OIzAybh9nwY7enS8fpiAzh0ua20uU6jsNiZUrZEzBHU2eWCro
uyY6uJ7rRxo9epAtx6I3wMmoILD3WyeAt4xK9n+9KwWwTfIcm7A6NVcARZ186OBhgL3qPWg0Wt0I
STJy7yuqEreBSfHBbNcqhJ/VFw/BAUplL46a6EateB5veC9R2jJJjjGsiz/ZKtgjXUQqpXtfGGTe
PEoSbU391p/KBAK34e2Y1jv5QFyVyvZBoUBqvZo+c3yXZ6KytaOTjritDLU0nvBfKGllDkTEItwW
stf5no5ecv61Tdu2a1+UihZU8CPjPZEZYZF/lW8Yshrk8X720uN25oYQy3BvcQBgjWr8VeD+G5nF
VQcaghURYJPyYbGlRcb9VXi2Dl8XTeE0idkaSNblAbPq8jwoCa0jq5G5h1ofsWr9+gphRGxFidFx
QRonmucOecXqUwuq8AOXK4WVMIzNFbCAx3iO7s+wKc1n50MPgpLHBkKf/tNw4DDOi/G+PaCd3gIF
U4fp/I96o3Qw8agB8V89uRUmblyDkqgJE4wCZJyCvcmJuxSWlZ/bzNX4zzifwnfY92GP/c6uvBzv
WXpGW2vr48KfUiFHkmnUZp10NilG9SgjrBoxNF2AsOpSYifORC3oi/L/I1/jfPk4pRquz5CF9Q4/
yFMh6aqZ9A7nmOgRSfeScpar2cV5SRWWfDkP3DyLmTj+DWXU9BTlowR5WqcvuHLLiWtcrcbVZz33
bz12tHPl23xdfuv+ODwM/78vx2rFf1v4RrFM1Nw4G0Dsme/Ehy+p2HLHSb//JXqeqTW1w0jB5mq8
bDuXTC90z6wwdp9q2SuZVt5hFY1HeLK5EnvlD4s/h6JB61z9Gi0c7FJo1/0kFW1u2A8K6FwBnodT
t+SmPLiyhzWE8crZO9WWf0F/y/IiB08VRR7LDEDmPoiV8l6Lyn8kl0hfX5x1pJ1NHbtcufRPWL10
XSg6Tmcn719i1klyALmUuGURtHWpuvTsh7yltOmRiVpfJSAAR2obkvuObDpYOmabv4VBeBrhVu0n
j7Axbh/+2aVfIHXHm8C0H9KInGqEUkmkvZGnNWzxseOxvYex0XdytvxdyLRymebMwndCvgP5mRp/
F823cqzyWJw/t3DTyEvwl1zQnJcugHH6q2oDkdce/wgNGHStaXu11i5KKNjypT9OFA97nYC/Kgff
nkuyvWFFa0OytVcTEI4Lcuroh1q12BE/RbR/jmPxACvS9vJYDsKnVmcIEtwsVCzTTaTfbM6aUImY
0MdL8/BmOQsBgIF7L1FAKOSrAMChGr/YX8TaUEPB4WWWdy0GbGHwCvK4aWo7n4tFEVp6S2Euiss5
HBom4zj3wgoWJgSs3UWaXdqTirNZlaBDDMhpfVRlq8sqIKPaX3Fb61mXpUebzO8leGCLbMSOvsQp
+d5oVOZCUFlDa2UKC507hbx0E+1wRbO1QrOzpirF83si4JjAh2pRGA7QQNaJMrdJKgWz6jhgjGQ4
ot0yfRYwhQHSWocsPitq7XD3H502Ps9Ci61nLyefgh3iulkVEEIB5n20sqjqcSyNJT21kackq2oC
7WjZWJTWcRPIbaf3Vh7Bl28oGnNlaUJnSkh5cL+r8iT6nFvwu9qCjnjRi1IRGKiNCLi+jvVx5xJD
oe5+/6kuX1RGTUfTwe+rJAEpzUSc9mfSerPinxL4NTQij/lCjdGP5hUVJ5sp4rMFjVFrDIY0sCxI
O8zF4zNmh1pthiIpPRsFMOx/ut5IBkDmmOYVG0n0wA1bxrx8tbLXY6NYxyVVHaipBw2FmEYPOrG0
fk+yQ6nzwDJVJkUPTObM3hrZYkbTAxCbEpuvgE0DTKU4v0QEF6uq5M+N385AQtll7Ls0dAK784Fp
ZQuComkeK2LRZU3FD1JSEiVuQ4bYQiIYrGMXCBUsTkWAX7xNLv9Na0z/hvFBxVi1rktL0QjDpMO3
A6uiuXCVy0TfkzVJWj0uDz7w2pLfhtfBkv0OFQ+FyQIu1mJ/tooeJp1yRpKhAzp7CJPzRSBxZPGZ
bej9+e9srvPLuZlqSL81O/T4sTGqpasXjUtdgA32jNryFlLB4uzUyvjHxcykE4jWHx5AnYMsvcNX
A6hN6VE0NbPKB8Qi3Mb3fbIN17zkvTAlGwHqJ8y8OwvGr73j2wiE9eEfQfmFpcpk4qJvOxRq5B6v
wAjgQ/fAKwKmnUxGbr9xGSb4UVndWm3nANL5aaMf0yQbvPj7DkWUxVqp4uMNybLmy0VoOtR0ZKyc
8oGMiZlesqBooA14ly0l3Dq+yOcTQgq8FLVnP2JFm/UcfBvSNSjnWLwuOFA0y6t2EkNe80p/KT23
BPVwBXob2WAFaFyxbe/WgpCHU9GjicniYTiY318kc3lGTcwBOPPBpo3YVbZdVMJq96gxPI1tWE+D
ep9qHsycIvmbxVM3OQxw29QxWfMdP/eKCZAK27AZ8um9qDet+hENxO7P7j1zURCxzPLfoH4geYrf
1TdB2D4qqTy5ho75PdgPL6yigeqQWuyXJ15bKFaP+VqxlNAMI0KP+cC2HEiKyAKUatL9+6ikOAun
o1b0CCgw3Mj3WS3f1DrzY3uRMuO3txXPG77hfqNMQ7FHvw9lYop+H//jlV2Eet0psaNDh8cQLSzG
drn1lAPQ09hHMNuVQnAL7kkPAT0nxSMAgf0GrAVQYP/QP9xNP5Fd84m44gIsU7JSXcIUDFS7uPe5
x6nkQ/BS/qhbNlbvJiByx6wYTGk2m9bWwypTID7eud/UTEYYkDOEaILwGXNIoppRAM3ZqtBbwuaU
CxNUIC3kYRsYWdsangwTnpaRF22lr7ZfWuiFICUSGE6rD1GH7G1LIbK49J7hbZn2oPZ00AmWr0DU
ZFtQD/RTRq0LLPXZBa6Oj43FIERScJ3ZkOziRAorFYsR1py+moaJ9hK0isWMq2uFpPuoCnfK3qT3
9qf7CpNrS2jStD2xHgBj6zfswyjlYKFJEm71W7MGeu9U3WYOaxlAMuxRT3ieIo2qQDLFjAiWLx4z
LQbn6JSydcZZfYtmen/o09iLAghO5i5LvKWj6Uf9hmmea7Cjf3zCPAqbRVxfPRKympEjEgWFqajL
jDqJxPOeXyaX7jnMSeopDvDxoL6+IH4GdPutrnxg4qIdG7HK6ZWO6p+vYHIrzb3MmNyiVVuD+zKM
FZYM6wiZy0Jd0IYs6LipKKSN1+M4qehxBcoJ2gMxRC+wL0doVrxz1LlM9poLBic7dh0TcLfADfNE
gDYVCyRr1AomIB/b3HYSf8afLYDbV0XHdH+l8pylCEUlX7Jv5692dtwkp9jLBhnZSwsmG7VptOWt
UFwR/r/z8pq01QmSzAvvnPAJJqIiSgPBGTG68z7D3vN8HM0WJlfOj4Cgq4NZMqvVvLheFF4nyml4
gASHtxkkV+lN5K1RFjnueJKc+1aYmXSaS6/fPsgF6U3f7nL5vPkAcsKCjON5dok7YYKu/r71WUvh
SZxXaO6k2/5aQr/SJUau92sXZrEptIiu0oatN9xY/gRIB5zF5eUUoRWFl+fMURtEmUeKyLc/k1/s
Kro/9SxGqg8jF8lncbs1Ys7NE2YXyXdqm660Mht3XoTLqenodWLrThIFnX3wEufgwgWaeLEdwIj6
Z5+Ktxxk4xY+K3WDnx5zTWzJFohPau1jOOrcp//cvSxK7TAD22Kf5NWJpvk4PCl6dL2HzGgbZAG4
1PEfP18qnGRuN/Uy44QYTl+ie7GfZM34VqX88adSLo3hILoY3u8QLh1Y7C/Blb+alGpzU8PAKngE
xzOj8IwyNkip8jwzQ0+mBOlk7GxNRxLnUbv8zkzU42uaidGP/vWMNvV0H3/FCxNlKFFhb/i9qQot
wcRtEXBS084fIKS8+tdDxmpYFAuFDVK0BCQrZ+7gFNzhsHZSA7PMsWb+CRhvU2XHBxXy0CKks8eb
Nb7mR9yZk8cXRkZal8UPkB7GAwqLnCCHxn99Kos7gk1U6HL+ibVSG00UiG1KNfwyeZ429xjDas+c
MddPJdsAGLyeYMkytnZebNV5uqVuHEQ/oMK5mdyWTF1fWDuUHPYO4XusEqdwnlwtzNFHSmwp6LcD
hJC9OeX2imvZurU5ML5EYlJEC1tsJabA1yXTcs+T342WEZjXJE+daEaZqwuXyTkyC1PNGI6ZKh3v
QtBQ3VjN6moEB2rgrqBTtD7q9uARXIHhT+puee79p/zMCBiI/Tx7h9YPO1veVYvkjPjbkw+x/eSg
dJxxPL5aryD0yr9vHHB4GwEVRic+vmeSUz+PXkSCtRfRJM6bF2EWY9c2j4Y5YGSZaYIbtiQo+Cba
uKgYF1Aw6BtdGGvn5MKbg0r1U0izUnOliCoaxtXzzoknwN5jp8FuXdQG9Y/MIhs6yOLrGhuQXybA
ec9zQPZyafjaZtHFT3lU2cGRd6i4EYfR339Dm5RaqJKftwxoleAmdwSHz/F1GU0iscwFypqu55k8
hrtrDI6rYBD4hBq6646F1nLf7WJIED4WcILSyNSLOuPzxz6+pFFIVEONFa7fcxq/20rHZZ7OuRd2
V/NIEoF54qyMzOob0vBR15qZOjIz/jFC6jdXMKLvjb2w+vTsw/vsv5RRorn/uit0wDWS68EErWvO
mj2dIPKmvq/t2eal8TDClceZuVnUeyr5qm3NMhZ/g8X9nsbGUtVsHoXkEZP2Pyu1/b9r7c8RMeYP
rI8/mSmnIFWkbFF0IJMSjaItepy0/yTZ0BhyNot78Zr8o4Y/i0SvO12C6/qnYwcbziA04dpzw95t
KegdaPWWAK/COLTSRryEkwsT4hxBi1cGb5J9ct/NiGhDLD0ScGb9LiDldAPRFKuXtFLYtakSFr31
/GSEkq1AG814ba49YhForqi16o6YLI9OT4vQp2AnPpWhQicP9IcW72xApNhB0ejF7XpePvmWPay7
AiOB9biomwQJAeL/SYbnVck+v6+uCGlMy2yZU9quWLIwTUukjXIg6i3eqKkeUuiE/s6hPztFGI44
OWIJbHLznBzA1LAssorI/mRgMHil3FD4c5kcrcZn+jo4iOyoVsQk0q2infPbh9d71vTlVd+baYxq
+aTWDV7PK92B9rBzbjb9+nlupZsHyExEocJknCqZURUJmYgmEt8OLHOItyJhNabyyqO5yTZgBePy
LdgkbS1Jp2NEDiEWIjLNWUWcyv+2O9oAtEQGGpC0Xcf1f1m6yOBvQ4qdJJPUK0iIGsMeO2CMs/2Z
swaq/UdqMyWz2TtubUKWYZ9+4OJz1B+yl9d769EeS0xwbdNDdVNnoegdZ6XQUUM4ABK1UQlNhegs
SxilJFCkOXfNqih0s6SkL9yPAX0VBFzvVQ5UpEvv2Xtrw2DB6Diqx0pr/ivH6H49xJMVqLZrbI9v
fekdOrdapMyf4oUYV69I1qiJMd5OHc78bbC7KVRgF0uQCRjLfC2AAz6+hPMQ3w3gtegL3fU/XvEm
xiAR3y0464+njzm/IxJ9MHIpBfmBGJyzVSYYfotKuyEUSR9Tb+QfdbpxF2DvNGpH3TEPci8AW2M1
RrTbznnB2D9GsSXWtSeVyuECzawOwrvolbyEOnWkCJHxCjZQQ/aajxMON58J1Hp9pZtLiQ4iceRZ
rGYfivqf/PoPPVMEEvVrxtaWQ9or+JJ75GsFivQhBDPyA1oujkzoFzzRDgxMp6iV5gxZCibqjBKl
yObqjD1wYM6u3sQ3A2HfzTaind36RDWOrTvZMuqwnu1h/pySP1q+dLbpVw6Hl1dXf3Do7r6wgjJ4
rDgxUQD5BmBRYNgRnMrim/4Maeq2Wjb0NQxmgEEcYvzlb/uxcXNl7pLT6+f7/f93+K/7gVMjR4EC
UNfI0N8X2pDn6xGTvV9XUykE/vdRQdZS1yO7ubo4eQ1TYGosUFP8wKUfEe/aeVvq0WxojfmiKl1r
jzn3rS+Cr/AC5WVHID4H0FRxso/rUMFC5UEEM/eb93veuvikXlJrUdTGolscIOGu5VT56oqevWQG
XwY5kEf8EG9GjDiNIcBS2Pz9vO5buZuU1jGhkEyoB84JTvE9Asu0p03Sqkr3buI7j/jTLcgNUlpc
UoFRZ6o447y5hixIg3WcJ4lJcAUo/h107XEh9BaaZvtnYN1k/ON/9S+drMDJ2pST2W62pzH8CP9A
9jZhMTw5zAE2YAgfzONpigQuJpQMLwHh0R8NaULVLa7I+GRrVtiPXltwtcRhZrzrJAc/v0+nOD9T
dK53f9IKtaZPO80F7NafcGqQ1KBRGHw32Sp5RfDhgO+zMmk5wTRYCGkKBHBfTnG6Gq94IwO6JqhM
EC74HHM0b2HQKhktnYrHHc8k6i1CFjLWecfu1PvBTtqYqvnHTm74pA7moq5FgBQN/pZfDNTvTtnb
NALbvF5L9TdXyyeAqMQVn4gffytrjMIonfEWoNEjXGf706vQNvKE1VnMqti2Lx+Kkb+wwfFLmpR5
UV3UR3jFu5HtPVYXh7LsqsQf3RJFr1Ajlm7nAfEApYtgP7maFMcCe+zIPvBAHCIipJvNxIMIU2pf
BOI/bSAp6IoxiRDVxM83PEaT8vjME7lzLPpWBdZcdxC9f5mg5nar1yM5qB2zKR+SvX9DAq4BSm/R
4SlvAFpWboXHhIFr17igSQjLuw5xdeyYO73D9w/Yu7hTFFIPyiRgolvjYAKubUQQXjN87RboW6Zs
HmWn+SOKSk5is3qZXBrnNhN47Azpl71jUcbJo7tQhJako7r1kI5vsIYA7Xy/ssoofE39FcrVwQ8x
i0qDsX6mzY7fB0nI1Vy/ZlR1GUd4yM5q3nTKxdoG/uXKhq3mji1sxjeIOhyBqM/83Rjmv/wUJzde
/2D+ay5wibi754sAiQh/9V2+3CMGOERlpl3D/0omNASQi4wzSqfaAAqbIVxRQ/+OK+hx1+ipBi6R
Wo6DHhbQvbXAuAuVtLkl++ZrTKyxXRW1KCkP/veF472aAwlh0ythfAP+Q1d7q7ARyE6dWI73BGlr
uiKUgDwkIZxjYVYdhcG+tJEJ0OXoeDbWhJ5y7H4/NzUvJ6IFperi0aCwHvuBt9E5eOL+ZOJ+gTeZ
S0zpUNdIyU3b94R6lbql/00b6IHAkSmnnacmzo83673J+BRFF8u6AO9L8o9vq1LrkS0mtIVnm3Lp
0sNjNpZpTv+GGMDd0su6uWpBZWPKq0wLku6gpQJkulREkPhXaZHEoCLpxCN1M7ik1Hr6HgOJ5y8k
3c16CVpjqQRXlQ1/1hb6sVuaGJRhPw5RaRCiA9FEwjyCbg9DMfNjax8A7xc8udz6jLAwqpf9QOVz
IeDTV46FSXhJazKNk9wnVBXjIKlXTgLSl8Rp4ys6LJzq1cSC5LulX0Vgcd0mXCpGZZdFfrizE6CU
sdVNyMM/1MNAhUC0ADBpHusHpMXjjQ3HKepPX9BX2CjPdfftRxdGwMc3GgI7tLdiK2+NNTzONX5B
JeFv+8PLZ1W9RYPwaHgI5imtQbRy8lW/4KLBs1onJN7cAgZFgHhXUrGEz7g5IqTT8vidcJ4VlPiJ
kmcZ01VDpYYHfW9LavguTjVe597PMygp6frLSW0myGguznQi3g/7SOoeNfpr79vowYgbEtFRd1d/
iAOQLNUUG/A3iG8X06bazrih2deAtaDngwOPJc1JQGjwlxrI7oDDTkF8ilLN7vg4oqJpU1sXaqKQ
LBhLqJrgzcrhP8ClZcfEUkU74OH7zqZbjrs/MmR7VeOKeA1AiLJ4eyVRFySpNEmBmEmdPQ2ojHnC
TTSCU95lESjPaWmem+NAZF6hSqxrjMDCv/6yrvpd7P39Xx0dYK5PNjBykDwRPU1ozA4WwfZeOebr
6OeBxBqNikn8dO440BOXS9tfplGGvRJOMfOirI17bQZB75XW/jus4dkzBhjgdqm2iAoQDpoZmkLY
WE6Suax530Rg8zjLHFy4i24TGV0puypjjt8JC1p7WeKhpHi3udpyQJITHMF8GoQz9fp8W4TnssW1
3PHD1igUhzGthOINGe7LEdcxtCO547nxuVoT8D5BhSsFxKuConc6RXVAZimdwogrn7HpoyVdZ+si
ATXYCmlzrOUV9nCliSLg7OYKoOasudJBqWUL5+B6o/d3VOUFIoIhgUdraEzjSH93Pv4W4XsyuC9j
2U7tdT2RRPG/KZOrvQ2h8ouV7EIu/snglCKBp/B9Q5+ZRKBUG/18ORaumMvTPy2jUo3jPcxTwkCT
Tc+JrHs34RkzJxHeh8EURraQXDAZsbZ/RfPzyV2CeV1edF9mcJf1aB/stBtB0g1MhERe3L2a/MZv
yPF23FS8x49sEUpLemCVLyG8d1OtLJgPOHT7VfIylbKKoKWbIKe2A5lj27uRzHnl7CEgrDrjN8Od
vKGZ7c7OTl6VBY/StUURPnyvF5b4rL9YqMbwZH95OjvfKZkMVbWO4+YPJbJTCmBQWugOrtf0o9pE
OYe/+26tosMa0bW08pJt7bXHWbNIx8CGrO5Mf/F9jF2RsCs+mmUDfDAQuCV4j/ot9qjXdjYHX22P
VqXkfG6rP95Br5c8ly0Ko4elYdHH12GahqeX31tjGrVsKEpEVsSS8QR7QV5wTrY2dAMihNs2eOlO
v1h+354G1yEvEm4TvQ0kWOjwBmmR6ZGxkH6o/wwf9mv3//ea3IavUTQ9uGNNv+2P7569AOFuoagy
+L1fdLkW52U+mAhwyoR+kVkz2N05015HLhOPHax7cWlzqhXEfqYrTjPTjqqLI3HYm4D2phTX6OYz
IuM8BWMIA24IpQSyZgBwVlcFVpHuCD4KlxEHvY1xUJCUBPPQhp1jlDzYz87g2rrrdz9ze5rrL/4d
I/VxV2Oq7Z+Ys6beWe0oa+7dnzYnbuvGr54FDPQl/v6ofbqjGNSW8weZXR28O18WeNAxkoEPB9Sv
PP1LwoeTySh11U+KsE0mAQoUDtfNAvsIclLWRJpj4+4smNtfbLwytjyezBazjD1KAGgroAuDVPvQ
mdblBUqNJ9K2m5OWwgNmciPioVt5ky3wMFR98fDgzq04KEGWKd4u7crRGKdDVU9z/FZXv9MK4+Vw
mXV1+Y4YybhOoE5t28i5JcgRwrSUqpdfW76alFt0nXA+KYm3MdOABspKAmF0c9s4rlmxsXJegPE6
WUpg52kimCWBypKmUpFfbFJHDgHwwsAWEPMdNFItQY4dErfojkCQPEPtd1/Lw8Vtc1Tqm1hhXbVV
Ho8CjIwRuwrmCqrD52IhLGsZ5tC7yp/5g1jBITJ6rKabFQ0t1vPrdC6e4H0G9C6OnRD8qJV8KD67
fgAvmozIhC8wzs9r8orZIavWh3kXpICuusjOP2GsaVAWYTD2/mYVaJBlCyOB9KSuo8HGcGtbUVfX
hCiVW+zNReMo+SNU0x5bMbNet00kFzPh6jnEwlhRhIVQMt88/nOpOlUcxKoPbEld+UZpsSr2gSRp
UjWtQGBbg6r+ddf7g9+dcKyr6k2jx+c4hRnxxrzQh6KnNrs1yLBpQzh1IakeCzk+jWbL6MwU4cDG
mj4AwZoh1JWdNAiWQFmRF1XQLk0NPcNZWfu7WTMQDaH2Qwm5negrrsj45jBhinTuRPyal3GhgAe5
qFoJZuhLLPsYC5IgaZjaAXAtMLxkWJD9iy9nSfElyMsJyyy0PcMm3M30mKEuH3TW/1q6RXl05CM+
fzLuQyhAlAdY/4OCW3aRJjKX5n1M7/+HZRQJm30beGQKt26hVbAS8Q/zOiergBO9nn2S/2OqKSwT
dOMx90jmhnrtydACLdNrrHrxPLJszHpEwQ6CU2lguMMIUoPBSUISeLYgf8J4DLZ6vX9APchOgKEe
RPRGJureuiAYYmiIihJ6/xDC6+JOJrS8EIWXd1dMwh/BjLijFIs1vvFdHyEvWVGIHTf5BuNdYfTP
/qvfFAzUoxfkATn6xqtNIrVxIOOUDbsIRlQ/NeDcIFa5WOYSTgKpPZbFpC/KzEZQXe1oPgGCwgqC
XXrTiiDO7ZExPIFoDBdarDnY56jb4h4b1TVKXD0ZrtpLYpajaPCHJ/T5ruUajwpKhm8UAHZhSoOI
9EsN5/BJRLuSpMOpjeOup9SMYacCHdzPgPgJmWW5Spt6O2nkbDdsIustXO8TMDqY4YN9/YZmzGpH
2Z9a3MbObdKeTXcvc4MJzBJKbEkGFZ9/pBB+PV7NPDcbpiy9YYfhQMkzakiz52ZN2QXMPBW3Y5Pn
9VM+HCXf1rTNrQLkG8Say5et7hTsOc8PF6WqlZ+tcJfuq6B3WL5XGuJdiHdDisWtCDXGzgVqzX0o
35gaknyE6seBH0cF0h2x84bjnI5lcyXzBDH7uTgDhKcq0Y4YhqV71JZ4kmwB9QtgmQH/5cnJI0+z
qFA8flJgSydfmhMulQag59BIWEsK+/J8nYpwTpOFFupi5tKm0I7Xhxr7HiRkl056uMMDWz9msUT2
EVzqH7MNA14d8a/Ilk7FNd73eahVE3UUnDy741fdkZLky6JAwxv1usvDUcNuv9k5AyHkFjYapTo1
rw/WCFkzHQ6joehX1e+8knXXAoBcSuC0lQ7bCf3zsIDn4UFMvpRgKhsHqQTKPkpqiZJ7BaAsBwUe
OAjiabDLSRKPh3czJQw+5dmcb5XJLviLX07W04EC01DxLItxc8higVlQxlb9fsPKYu/X1riWJRYm
ei+uerWiYAozUCDp/bZsfWd/sMT7zx/188nDkn4QVGfZ/+eunP87jokT6YAZQ0RNMrJOz6RX/3YH
iEamhWrcrX2lJpXL/DMwI7KFEl4jwWegfN4Qi/0L01ZmjMEnXFKkH+/5y67pxu85HrmDrrtIGdvk
PzK9bYv+JB+ay9nmavhsT6nNEEP4UEKxBfvWgzlpg702xxwB8JdbC0dU4izUj0bEdmgSBlb8GW79
17fBP8GAnw8ypxTsi9YgxpEHrx5LMpRADKBcKVXbFKthQMSsf4pupElKPqd2UNdsGb+LrqDQk/rP
2JJGgziQ9/szsOPBo9pw10kyCQTkJ03t63sFDfpnRmatZs4+qYBIUqmF+YjJQFCb68zzsMy1azd4
XAkQkDiYwrxHU36am0HWYMQUFYqCeyhO14rSRJ81+2wKN8mmn7v1rVPqgZ0bKNAnLeFan+8RkWFE
A5eFhU604REVp3+lAw30B30VWdEvI3OUEgHtotqtvHaIPaqxD/wR0b9gXtDuIZVTacqbVUaFBxN0
aNgbodykp6AiPRMlWCiS2T3d6vbHUaWyK2lpwzGL41GrxS9P8n2ss6YlPh19lNRU01hs11YegmiC
L35usWpwSBQg34rh0xKZSLL4Cy7sT3e1xUTUlUO+XGRcr0TUuqEaUWS0kmsEEqNQ00GlHwm9PFFI
yFr1q5iqsUHBL2UjudDT2DYnmq8rD4KcE+L66vXXlCFrvEiyYZXC3658vM/h7qeQtkMyTNca6S3c
rlVSnXnQOXsAUPBF+Iej3w2hewSul6XA8l5EiiVJL2zzU4A6Et1AIEtuh35OUseHYvDYmR9A5otY
/nNNyQMUuxdcurbPA6yYf6CD5ZRXrvnfzQfNtBbsazdRSdHbuRaFU8HhoNpb3InS6MnVxOtTarvp
A4UUVzQFXWZ5HV9TjK0f/dp/09PrMMQDzHYoQVi5jJy+kIHsrf3ynl7ToDyY7mGD72ui+NVrb0JO
y7uzXlbHMOGZDTonwF4FWdmiBIEXlJ5iHyxiU1eBmRAe1hX4Zyw8+tr0m8QlR8VBecZX9Blq08zF
K7Q+hAkQoxq7O2fO6UPEqEawzvWEgV+Z+0fQitumWo0bgVeFQ/Y4qOpQkmRfO1K2yfTHtw4t2GaS
yP2sgQEMXuNF8Yph8rOUAfGLi7HjCWyizF+f9OtkBjX+x1LT42UN/oQkRe98yk2kV1piF6HsAgLF
CpJIRFdwP2VaHxO19RwfHvdMMapfq6kPO4q5Wtz+uLLq+2MskXUnNkZM4rd++JAJP07EWbkijJ/z
RGiTkRsLxddRRs8ciu5elYEjsbA3HYerKFs7SZ6UNP0V23/2MeR1+PDm8lbPABgI3L/4uR9qD9PT
WNJFN5XIgmh7i9QfOI2o1/QCt5YTtq1kWO5B1D5giyrhV0cxqx0OH+UzzM48fT48lilEcbWPKRkw
HlBQnE39Fsm2nZ+F/nqpc7iNrigJK+Mai9RpYGcDAK6MUtD7Fiu3pGzuQHKx1eRt8Ey/pSAoO7Tl
YdK2Keo/esGvWXF5Jcmc9FQ6B3tgV0cfR+mjCh8IOCbc/wCjoW5kXfBTvj2wEv06shuAD40n1kSt
N40fWfKi/9kNkJP/KgfVRHzI01AtKbmGf7heYQzxPAS1fe8q5yTsXo5jRDu/jaTeVOQsVPUOpS/3
ixB8ArxwSUQZfzyHItagVhJ34MZsqp7yhn4neqScyFokkIO5XNqMNNdIgiAORoFCefth1g8FojbQ
YVAluBrNAlirWpCdU9U2O4rOvHLbGlFPQqurAVXyTGRAiI7LOpffqG4JnftVurEjfYbxu5TFOlGn
pyeFJNwL9O6r0SHdxQAc4e1LVILsBn+1lXNXQg4Zk4Iyi1gYeQqqFTAn+Oq3lQtwUynXzZTEmYZx
KaofPsaEP8tWhUuigwbrMgfKBdNgR7+vEXcW8coq09HiLNrvc/i2TR/hQ9RjHq30kckAuNBiiZdG
eqjlrt8ZgviyhL2EtLZkFKOEgIHy7sVpZMOjPItY1YSaPOMj/4q+kkjzfd/6YXyuQtRf2j9rGoiZ
+i+vBwjVuRVf2kugs8BXN9NolZgEEPwuVF17jFGckClioFy5+C6xQvCIi1Qyqw6IsHlrl9TNw4v0
HQNwNfiVefeXak7FIgYo48Ia71hRzmdYKtsj6ZZ7vqIgBt5EpGcMY9h6Y7LIcrqgAYgId2a3+RpL
QqgG4S7vI4w05nnIQRSrY4E7fNMvaG52Bf/6FB1fuOsDXLXWXCrzKHeya0oSSi1AUi2ywuP4/AfC
KJQGxj8Tus/x69eanfVwn7g07wIOFwTn1XgWLp4Hs4TLI8UN1hYxkQnVMB+38LnSQceiuCkR+icn
hbyLUfwBl1mEL2+h+CN6+n7OUNRoQaCNB6rAqbE2FOiT8xN4uP6LMOXaHkfUY4SMjk9m9UZiPJe0
47NyTyuzp/ScdLkbUGb5oxh6qYrONAXd00Nt3mAdJoC9Bhq684OvFJZE8az1dqbjaAZYI7CFZyQ3
FQsbIuQNgYUPdpSH+w0KPC4znssMP6y9RukGN34Y1oFRPHNBTAkv8KurB/XXs8wN7etD4qfJdDTG
I2V0GjpnTB+nQdu/vFKdmnQKIIE13YgpVF5q1XanLTxe5CVojMLuSeMOWjNbZh/k9F93xMurFE+u
7cVydvdnU49lXdHQvsTLq3yHpYZIlAPZgPjVbl6cWZlWq97eS7tMp9oo8OKcH/IXCnNhKWQYJHfj
6n/mY2PoW3qH0eU8j87YrYkzZxa/awI8KRptyDuls17SXdfeMOuVFtrB7v2P1QNmJD9E4KYvp5bu
H56EAYc2ejrrSxGax5yGkTF5zxFUFOnpj0o2tPSjhp6XWEdi9PumV/RuwSGBOyn2RE30ET5bOp67
R1Nq+Zvni2HX7XlSHWHTWPfrLNzMwBPDcdQXj4JHp0XsbAGudCtluyKo89CYAJqSLHdsPLLEdR70
GOyEOQbegWgLIt/4FyN0XhqqspGh5wvOiN0xSjLrA0YsXepFi6GpLkqC72g/rL4JygzFUFPsXmYN
68A5bualkPnlTA2+P8JzCHRcdgzgGucG+MIQTonQSr1swnLAIedaNEJBpZ5fpPdmTkh76geJJQ5M
+/a4AegwtYWFW2Jx7thjK5uONxiLpxq78HWlNU2X+mYNlQjAmlTCG6kPdorBNouAM/84xLfbQ3Ky
71gxc4hc3YfXfnSduD9xcTpGBcwMkoKuByYHmrPRkFEvkd6ODZgWs5LEpgoLvmz8ZifSdFM/j0rb
OjMDazYVFf5LkOoDNOVEdf5uh3TDhUD6unKVMg==
`pragma protect end_protected
