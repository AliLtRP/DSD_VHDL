// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
P1hGK3pNNq1x6dUqmIvACfoOQbrJbBKHYYjfGePdSOswIdLxU/b8rFTHzRan62dl
buXCFtIDodfyBughS9OaQD1WOnBOEKoEqhYi7xjLym22BdVGJJyHYInCx1KMli6f
Nk4xziD1hhpikD4cZa8zvteAE0IS2i6G0l8F4WOLnac=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9808)
ZIy7q+X/2PhgWtLs9kAuFKGlojFnaTiltEI7vFvzXJum8wOq6W11RMwLyRZZAPht
JsZbtJIVMCV4SXGwKsh0ge+2NMsmRePwOxaOyxBEfeuV2KVLdN6kvZJptZSqvish
WHvV9Svbd9BX+aujTlWEf1YRoswmVTs8pnvFM4yQLUnvwPiaE4mi0n1W48VXlldg
8wenFcTZYS7J5uBJEBWeP8ZW6QNl91bMPXf7IeySTKmYQZfTT/amzYa1y9GzL+lL
yS/SrkoI3UPiIPPXGJVE3I/0IRaLZqB5Hul1Q0PpdoSfmm8Oz9S7NqIDsC/kERgs
hDOQf5eTs54XBlm3gEHShkoeSSkCR+xPShTfDuHzfxpOxZ22leviOXvPiRgNU8HV
A669BS76F/pGkXLiWn6Dxgj3QGYev3tFjctIjQcFsAo7PYfUDWEW4HS7djdSv5oq
HnBgLhbNtzjRmyA/mW0UUYBUBdGnFqnT+DlGTolbdqDlOUA1DH8N6L1eXVoGYANg
WbDol8E/9lTwPp7Nsm19uFVQaEPCoObnxfHHTnRylc2mayUz2lu10gewN7gq3h8D
8uNlWPcPrrG+ikXBFtBlObVk97c/TD+5IZUzC/4cqj8JbpYDcVwy+/VBHMgWjBVL
gMCfU4zHSse9lJvTDnM6yDNe4WJS4E+nidAF+MFWmXKys253eGCziPrfH7FaRpkO
VSNYKJpj5aqN2/xYiC/ILTM9VndulwfdcvIHgnOfSFhorZJyDmCEjzWjfk6eiKWA
8LhlcbRJSBr8+qlz4KyejwdOqUvI+uwJ/j47NVlkFEBKpkFFXLmhhPOYTxr3x214
yTX7sDN9mpFGh/7gQew3U0SUQSNqNXYg9A1bE4NM7hVUsdHFBPjJtKxuqfrHBXET
aYqU9mJb4NgHd3RKirM2UQ6bBTccI8NkmjzaPTUJcOi8tmLlBvQXotVnLmJogsp+
JMr+EfUF0RqVauYzwyAi0CrutTYj1VrvVRurEkLmJGPNH2YPJ7HNbk/MkKXZHnLn
G/O+DauYyVbKwcsmjsMF74eGpzksFzgOgRbhhlOvMlx19NpzlfQ/5wvHT9KMAqbm
YA6cK8gcNXk9368c8ocFFfzv7QnQIbkJyHrfP5T+3617aAlFE57Ysy3ldYp35o5x
eHIsmf/zwOdi8mM+S+dUqweumvGYprX5k/zaGirmdAgfh+epZH2aQPCBxII9sxyD
A/HSkJ2dMCdRNk/fanQQML5BiadCaoufJ8y7D5rZsuRbcC58zlcU74BvYEkpyYTA
nSuZEtdUMHxxQuEsTf5/6LFcBoXq2+G0mLBTldKKcawNpq7YiQkNYil/JiP+h7ZW
ikZ7VDHr0Yq3ia4UwMCGziPL/f1vk6M6CqE0bHmt137aS1rc27CDW6kleaGqlWJP
AJp4Xc8ID7aN5EZCZSOF3pphO4EKDUZy1zB1x5i2KUfJHiI0OJXxmDv7CjSu/46P
1hDnE2U9bg2jqsNQZjxxEdi9Kgl7wenh5UK4azMcaFDTjVT4rNnlKKDTwiKPPVG+
HjOW7SgmKWmPO1vM82yzTbZvVdxY0OgJuvnxykqG0/zT2z8cwr7vPIAquaVsIbLm
eSAeMfiKAR8i2l2WoLd3mWkrbXPMx65pYeHYfj2fm9c7Z47404m9GAImLVjOBIta
quO4VjlTe8L4rCvUV461FJ43sYs4Xb6MJd/fwRFgywuCREz1x1DIjkvjJyDCvWn0
TMswjIE/uDn8A4eEqDr8iK2dulANI3/lt2hszBPHXaOmaXbPYw0jLm5NriNzxN1K
sq6r3BVtcP4lNiyRs0a4YCVa/cPwR/eIn+98ri/S2qElGYuzCg9nNXNpEolJlrhZ
nMKfX2dBmsf3iRSEZRqhjTJNjS3yso1MoL5ojOIYDQPgaeK2K2Dr7Q9ux3fYI11/
s02Yci8q47m/6VnKg0pcZOHDCIhbfx7CpF5dujioF5sGBX8to/R3Jb9Mz2N7rRp3
sf0CUjgIYg0T+NyurA9+7tsK+Jv41q05xaI+Nvu8jJNLNP6YSksmRScY1qWMTCZj
4arheKxO3tNXOhcnOWInQedJAECM270TQUEZZnpxsukClnXobmi5HMun2AfYM1da
gK4rBwPbj+lGSM/EA8Lt5qRizswrERsxjJTB//Y+UIwxiidr5o+km2vvPO7d0MdB
vhlCMtQTNi/kxJNv+fppMdCX29iUVWhM0RKP9Be0+ZEsmMOT/mkYXPo1APE60V4V
wIMuMfGfTvyRLl3+uocb8K8CWW9CPvQ+Y4eTtfluFLMI8RZ+IGq92SeLXeBPlc1U
wQya5X2sh3brL1giNgBcoDfDuctYKYRtvKQ2thelJX9uzBri5HOubX9jL7TfkAop
/3aqBWwIdEBfKXN9CXpM+Vp4PoPACCT6QcEuohMIdS3OMcJpQBZ0nOtOj2yfojTs
HlvqCBGuv6gcmDqFi9NdEtzybRUfvjmGkOF1GIN7adeEN3gyZy/YwR38xpy2Ot1N
8QPax89/noSMEmW7g8zObijYNaXEt4AxRQ0V6oCG4ktxwiFqyEGQswxV8KWebkLE
VlhDPv87WUFj+OTH0fwIm6E4rD0PlhKYzdsl8zCI0upTQFlZXL6PNsvCjBnA/ZGv
KnpxpR3E9H742UQB5/HOMWc5BGKoQVwys+QmIbDcwc+80xSZhrTs07fF9KEn/WUW
QfgrSLd5878u++VIIwLvCPlmPFosqvzPEBK+To2OokpP8ZcCNpzCzOnHsWmTXgjb
cK26b/RLMDaoXAUVTSO5wWwMBx7TvwmpTQL/GXl6XG/uLvzr0U2KDP4h2wxZAPPP
B96uB+0Tkbv4mhw/G2xPHB8pCZ2LDZ1NFf3H+kxp+Vda6dTGKfxYPVGr1+EqBnu8
jWWy+kI98rp/V8tA+lVGF+bsDCNBlaJowovgmQWzd4BkpJXtIXo/XYPf8O4nkwNM
YGIGJCGmiA2P+2cGZdLLhluJ0nrpBqq4K5XAPZGY5Lhnf6PPqYBGRBI7KUMMK8WJ
FAwcQI4qbqjReoduCAwpXn/C4z/sQUIVKZ+wCu9E2blZnORlmKR9ydnDFP9BzoTf
uAXE7ri5b+IbwQ6PRXbYMMzfgh8RJ3KeMFS5jIT0Ep0R+FW732Wwdxc4AENJo5V5
uGnCSg0dwDcBWgcF2XV6bYRThc/COHFBEvRs9C2asyKCzWBLQPKv4LqK0FbKYWFX
MGTUL4qG1Y+npXbftVaXL4ojTOzNJ/p2ju3UBLnbCFqpzF/BXpOfrC6tSCGrpq/d
QlNUGocC7LCPOMqemLK6K7CNgRyTWFGT/dQeIp42HBe95BALWb0NM1zyGqAWLjYA
MWfzCPikXdYOj/SeupEmdei6X134ggJJbb5+gx0aUWC0+PmjZXh4PdssBsfUar9l
awDK03pevrO67MWzqi3K4nFkDYPWibDib+iTRZE5jLiiCFLJrEYeDBK+aPIAwqKi
8dmBnTRndl6TFkLKKFFPDajsjPhsVbecB467rgGjlO4Bxq+NJE3AyUWNqDBGL4fH
OAlUuxe9Kt/tPRPaQs+ZQ5W+dS2dRHuLUOBs90L9ljjHKOUi52PIBmxkUovzMxqt
5U/2ihe6aYdb91y/Uy6T7RQ+WJa17p942gRmgL9gSBwq2H2wHMUJwQVDBexuFZWR
o/fI9ShdL2HtYtF3/uYzBl9xGhY2p5EsEFVFLC6irrmS+HVNlLLpSZzTCDD5Nrak
OBUJAopnbYxPbYazHYB2tgBqTCMQSiy92v+OgYS2FGmJh9ItSvB5Gfzln5XXrUrw
9cusfhV55sgQPiEW8qF84pGy5zfmcB/JWu7ltTks6Zfkvp/XO4mI3JrUZNth4CR4
oor0y+m+SKTYMLysnAHihHax/AfDdTQRF0J3q3deA4Ohx64FRhMG3eqraM7Xopcs
OdKlFM1bQrg6t/3u8A8MmhFvMeC+4oF+i/c6inmPvB56CxogvSEy4ZW/xjAAVPlP
lsDG2AWzO3qHtcaJAoZdoSWW6x+9nkpd0b7N5GVGFSpzR6UDauG/eCy7CHUoKAKe
on6gtpLXU1k2pRvsVwnpHnzWDmXb/81PbG/kK/ynn2Q7LrelRdQL8si39sFOeWcK
5O+JO7qu/jevoRx4VcUEGgTmizZZwsiYsyj+sd571TVH+uQzP45ceN3KjEGYdS2X
tQ9MtA2dTQvHIzAtsp4lpSUECigN0bjYuP9cCPNU3yefGkVhPc+YNmxOaXhsOPxB
xP2pXWeA+Cq8e5BWUj2sRoxNcwT+jIfAjYr7e0Eq+bWyhhceJZHiE0jKrmiT8ICb
OURobhQPoMOjk64fnAS1cjsiGUyYRQkKB0ZdyZAIsGGJIK2G7mQ6zDyNwHUAuFvG
Wn4NGiSApP88jkGl0tVHWAEP4hXXtsF45FrhgPp6x8I8NJ3Kmh9W0iZLZDviuI1y
AFJwX+x1xLzjWsyY8VHl/0Ou3MzDXPaHUA6tzOHMsQ67vm1HQKpaEiQLF9US6/a3
i6xrzQjHoQu0eSDgZKQOFoNxYQLXrlkZ+i/2nDQGySbrDtoWTyWvfg2tsCdhG1cF
n/vd9QfG/ICk+CzLEMSgNI6fzqq5dsokp56pWv8+r8i/EEQJMZ5/AAJDSWuFLQDI
3IXjUPVIfgtBbt4q30T9lXRLirUYytP8kRml94eLLouR0csOGUaCgEjZJJOBySiD
w+Ve1vO/vSc4Ygkzz1BZpvlQf70GioYWJ/DTNYt/6gnIx0NiSmO0Gh4oyYDmyYjq
55v1wKARIkYTwhafUjRyp2o86b3gwQdL5IPoer9mGJgY44j15uvd6plPv51DZV0/
hbR+erQl8MxqZgdHKRVsmYnxP3fbCyqL9rvhrM1vNaI4v8LGKJvL1gH+KW66IwHR
uC1haQkubwFPT7X+I1zKB9m2ogqQL/Q4j1A0GvhvEogmmxEE/mj9KZ2KXKOlzCEm
L8AF61UrljQC0gw+UGZcatTVKmJUlKX4rjDxjwN/lDIWNuZ1Zs17smJEijG16r46
CGbWVU0GQsoW9QzL//Eu8MFOjhGtAWliixxNTbQ11UZT0qwBKrz3jvUjE4wfuEW/
skm69ADqsDnbzbQFTBQ9e2RV8ryjgffewHcgqL4CSfTBZihjGInz0FMS6E0W1y/B
A/Ri1LdYFBoFvQukqiWfMblR6XUAj/qhNkkWdhrCJxNjBcLMoGJ3ylhM72r8CYgv
3if0UsxzEYERJmpKfGeC8Fz4rffN09cK0ErHY804/+7W5IO7INcnELajNR0alOWp
Nl2LhSyqaa0Z5fMEHAmIMAvu9NcPsx7RGY904aJqqpyoLtFAzTiQQjFLalNgZttZ
jxHHh2xHFFTFK15vnDETBm7jX3fVELk8y6g5NQ5eQqUo9mqhU+EtCKSR4nEms+dB
EDyTkLqgdw40xGfWxz6ki9rtCgAD59Vx2YmG58fTk7Xte8CpPYEw5HVMApBBY03a
yAMTrv03ICHAwKCWFgKk++MaYHf/ka/xk4cwOXwJXHv+++iIjflXywKLq8D83Qeh
vJoftfCUSo+Ehfrm6O6cQLe+zWveG7KAiBSIMq7/iWBiBGylAxsLQeKaN6UGNPLt
QtKqEavty4m4a3T6tYLBzpC6y+zSMe92xd+b37udZMbbvqSdf082LAdIdSiDlNZb
4PubJzs2TiJFykweMP9l64GA4wnf7omuucQvp+cx8y8euWWHTR+vR2gSKdaSvve8
B4Ah3uHyF+PvrF4ESHL8dCdGZtB3uA6nWenxryzjmMUs1LtgskJpooGGfPfNC27U
g0Sohyn6l3W5cgz9KLg2RHJc+RXfYoAzdU3S1vzQtveYAOH2QhWal1fswT/0B5Zh
nsseI6RhTAE4IyAiwJi7/OncsYz+fLVzSzgfHkPMlYVRPGTx1REGAqQc3dh8MxJp
GroT83rn1ASMtk6lA3z44ILDV7xtYZ2UZc36F53KmnBf1CHic4DS29141HyxqvM7
k6rTEHnZ2CdLEYES3OyLHw+EQ4OVbLM5JRcgs93j8BpjjR26qrzvmCfoqoO4uNsE
DPSrJFELvrV4YzarShx6hJgQP17awhliuZLRY9V/sHwZh2INpkhVI0vv/YQPZYQc
OLKvWFkJ7dVF5/oQIPyHo0tyFisdCpecTq/BsSKsjBwLp52z2EgqsSwGBsfi4CYu
DFrErYMe51LbH5wy/kD62WJInRif2ODnZCg3sV3kcCwy4PeZcb2vWEQpgvklMzIZ
egbuxlxGsZwcbP8RX5T0hTtwrIPH+SbL0OcOkCewffbE1wQ0Ia8rEotPFtW/gPaS
u3m4W8tBRBlBPo1b6zDK0MTh8VxusZrABa4v7R+dLb34ScxibEb+r6muDhChDZq4
yyLW+N4bfq9vH1pyDCnalPSK+DielFQJ5b73g30+9rgQApqbkOxzLUQRBlE+p94R
5kgwccugDl36Kqsfv6vFxAR9zA7QkK4D/xuJryLZq48XzBR698/Uy3mjbeo0wmga
eEjZF4/syOaRo+HQ2odUD87Kv5qSnY99AxBpdB/KsO0l5M/M7qgoomaqyw7bqiZa
Rstd0/MvbCGGoG7GG3VLu/yH/AzbZE8IH8xOcLTt89q5VvlGz2wMkQujTgDr9btk
v2qSwl+OXSYJnNnung1s9Ffb+oxzVHBJ5XF4pdqEWkx5hO9S007BmwL+p26YMk30
8ovTBKu2z8VoKvps/WFNm1GjjffPkqv2BeLYdAXs4pKUPnrzjN8b1/RfKOidz7Ir
Dh++VOQpthzGTomaCa5w1px1/SRPkeu/rwDTh3llTvNd5S1bZ4Tz5av7yLQtUgkG
eA19nmts+f12/RuDSsbV8GkSKWR0BCcWv076NUne9KBuMO4NqGFxW2sI4wOnxTjb
C5uglIbpfG3plPadaqNEDGjU1mBP4rpOHTjmYKVNGjZVKu2LLw5cWF/EyGAXv36r
1QWgGlnN4/B211HqkGfAmudc2FsyyFWsj85/99bvWqbAKhIP8ORFPJvxV81uREfv
9dGW4E1e+YrEaf7GdRkjr7505ZGlbNSijJq6O+FIEuvc6LnOEdHrG7cDhMjLp/+y
DAe7D1VFZEJqE5jG136PHE0szgN/3+zZUB+/wzd6S1xLC+VK6PhSIfAhV+x+LZns
7hSP5tJ5svIUCS5B0w0AoWNsB9ehFSix9h9bRMsDAqXm93LSaZBUGfVteCpQSx6i
DCSkUzKaNmazbhvVQ4txQqEsInAJh6itY3wmIzFngMYHF3eTSvXJ2wuWAOGTi1B5
FNTlL3KTm7QSV9GAGwuXiwMh0GaRvxNlA5Eqz+a+akL7oQfAXcvZdNa53fQck3iK
GSZVPkOv0dcq55MvzZf/ffbll+bAWvSPrw8kbNrBTCL6CKbNnfbaoFUWB3paPTrf
vSHGrDl3qrNOo1x5gjVAi3CdLF8QbLaryM/jHTzLeIo3uWOSk4hCCE6qbiYHovRb
2da6UAsNA3vB+PCbTAIqcSm6/OHW97JgW3rAUp1UzsBcF/riZXz73qH+V6hqxIdP
FHBSTexhl2p6EAMF8tByQj62J9WPl6N3A/MWju7Xit95/N1IM23nIkkEv7v4ig/v
F+tVHlhjfumgtIvDe8o4Ig4VPWuEuhvw3vF5T2Kk3dynuWin2EeGsqGtF2+hZLcO
x6FLy/6DbMIEaL1BxQXZWPDjaM1LvRvZMeW9eUnCyrBxbkSmtWCrMWpEG79a2zpS
k4BnzwP2BDaL/l6xh0FXoGTyRP+l04zB8qjhFZPMcPRQukr0RhSt5DLjyCmgpx3c
zuIALy5INmkpkN7f1d8Zz2Yla0F11HnCC8VYZQP9suIKEia6QiikdS+8qBe5h2tJ
dWhZCIRUKciD6GjoA9yD26dIR7GPuz3CLQfQ6iEAxRs4CbZHA/O+1SWUQCNEUTlA
+1RQzzpEiTSHzvMqLP1sYwWS+xBxFPIIoeuhjFc76NBiyz2fXH7LVs943JrxK8xC
IeUSMQyMefcV04ACXltTQnc+yuK0++Ub3BSertwOzfygtpQv8AynMvcI7LDNTEz0
bOa5kEe5342+WIdgTliy6uksT26T2Dqsac83KKHiOJ7le8Z/iharnJ76XnQ5Ix88
C5x+6qnfgdIMJ6HoJ02rnpVizsBYg1GFgXUB7mlqa9nPpPLvkLV/SsB61DLVqO6z
WNA913uKEN7M4KEb9oxXljmekNp5B0klqW5dF83UiJPYlX5faBkHHUeQYMRcKI28
r6f3IZSLr6geiZU2WK4f8X6eV7ri2OIQZKq6V8M5GAGjLiNPWe8GpqxCCtWwLWvf
Yr9A3Kr+ILOcHtdgS+VGwidg4qKGbHxpvrI28SGn329OBajLdlpZFtkXHxBa6Mut
ciO/Y5t6lH7l1BfNxFERmNXUIdV/4Kb4wlFLiJ8a9lRV0wjEdMAYi4IkmhuX7oU0
4ygI/fLr3gWriOW++4YJbhwtu6co28kS0xDr2Nq3ajVwIKO4r6xCsR2yVIKVDS+b
wy8ZK0ynyA3ger/MsIq/tSfD+Cmsv5qcoj0D8/Hd0/ctyxD9HUQelQjN0ebOmWid
Pkpj7/+ixCc5k8qkjQPTuV+wIl+P6o/iq/xf97gnGT7QUhN+T2qllNo1xLnztlcU
83zMPWqC3GKI4TFYuEpskp5bw8zyW08pa8c+7QkjpAznlJ1txekTeVNo3vYqJwBq
fp9NLRpieSpD2IQFK/Nn/ujsFWMZ22hGMgqV8em1AH55i1gjmDqzwcStj60658Q8
l7z6ttdgSS3tCf6voikZfC1LF8N4K9yupBcdmUIKwdnegdehMj0qbKz9ByhR4bS3
71dg8eqrpARbHjLNqDGXmGtDpt31GIqcBnZ8pmSPZJmIjh0WAl+cnHuUlUBYoDxs
rx+UrZnBwc9r2OyulIo4SI+wb0mshYJ4I6H2EEXnXAsukBDnrhvacqSdg89ijd3I
r06HqcRJWC/AeNZGLFtWDskJF98DvCYc7VZFPuqwyK+RK5t3M8z1HZlyjCoGYN5k
vPVVIkKmowh2/9A2YvpZ3ofDcSYjTRzeL5Mwc9OJQkRXQJa9C0UAFmspc1dOhPPR
Bx4PMjt9za0JjjqjRscFwAjws9R9wjPMgw8tPOlDJ4RHV+2VY+EbIs1o1YASEegF
y0HbxnS5+UntoTw1g1xpx4/BIkKDRqjQdChVpNQpOygGkeaQdVPfF1gzP/ofbiZl
IcFmnprnNjORN2ZHUzcHrba1SZQKFHYmpu3g2WyjX+8EuPMgNg8BuVYT6R5EBMvn
A09L6yiwA9VIidg1HFjWSTaSzISyKjlM2qw1AQOKR9FBqNg42MJmjGGeXlIe1MNA
u+3HpqyPl5ZjjE+q3Wydv4UZn1ioMpPUfFGw1GFhMbb65nKxrleueHNKRgZF5mkO
Hg3g02b8DVEYNOkgL2QnuI1xmVQUEQQ1ylNTlDF3IHmljADkBnJ3hzUWb2rsO1xn
y7lMj8JqHZcECYuft9mTqkOpwSHG5GxsvQLZQZTOURGHtL8ciYEiDMX+woJLKUUt
dOivuevek48xiIjYQU8WMUALpivamfNTnADreFWTdN3mmR4Zg/twxX0dIqGfA9XK
3zO99kgkYANhlCJCdqd8RPPUCjnb/rTfFeOFnMy+U305cT0+vbVZO4jExS+I7jaf
+YokV/84h+DZvq7/OP5YqtO+m6jNklPYvB2ysMnkBYvQ+XVKo5DRZoiALlkgNkIH
3DWHk8Iqa/U1p4CzeIcRVmqSJOku8L+F0rjQzUuEJ+40ZCyrxyCoPpkY7+7eWgF7
kTtOj1u0i+eDdlBnc7OXrYg/eSCmKkWiGNDNPZHnplZuP/fnoyhlrVmwndNBcTG+
NQaj0DFFjSNr56lcBGuNZdVpC4uw6aFF0eqeAzhvh/d0qNopM8iJ01LZM8RhX6U0
3YQ96JsZo4IHuFLjNnBaj+8Z4Tj57Y1JqYl7zAnJGsSWQDZTM3HhGxNweyIna6Ht
e7gh0E72/HsDff51d2nlKo/sigNi2L1kHmBLIwjKWUvU+6aJ96qK9khKxBskRXIq
D5B7L7E3M2AS3eFaslCk1usO5PaSucvPFLNk8+4v9oTFyyAksDWP2Syl5P9wRFdD
0VhUFOqywO1wb6af1qKhJtpn0GrqabRLFeJEf7Jte+cBoCwIlAzetVm4agOlYG4G
KtMnIkEYvMzIeviKODT7VMPl9BB5jvYkC9lVs52tE/9g7vX2pvDxQTqUjdVD+pFv
UOEI/72V53ywfmUQ6+04aSnUg+zwkNoJ/vXKSh/9MMNOl2zxgYeRGI5ViylXVY6I
8QCO+c1CMr3jrN16ngGSLulwECLFOiQ6xfDGtS0Tn8FrQojvzuVVZ16XyJN20cQb
Dj5uwJLDctumKF3afUkZt+gRUk4XEUfgTld4vC63lfyNK7bfxEn6y78sA4TvQKkX
/cuYb/3W1WbyjAM4gHGepoyDI+dyh8SXtZNCaURQLLTPTpaIe5U8ipHZxsYgXknd
remPcAZR5OmJFffw0PxvXbJ4Cul3c+StRqqysvLZpVyznqbOeyFRFce470kf2zD8
Z9SjaM3MUawJdrsONoUlG+uj8XeaqFE8zL1TOrPRrTCaWoNaBX5nrsP5+yDZmMRc
7fQkJIxDu1QcLv93DikyjtA/mTpRoVtWJlduzzIMfXVGckjjE+b55Wxw0JzivEq7
EZH1jPXdOD9pYFl488VLhFj1xXe4AUZG3iX7S6yWN08PWXrkAc+GZN/N2ymPJMCA
5lFpK3KZHvcGVPzyUmgmRFByZjkpm0xgOUpA2lmOxGaMK9EV0mxp1CJ7+hjivVL0
nsWb6UHbCdLnsB1YZnA2vuil0k+/KDGu2l1kZz2bnC7T+8cCI5cJ294YIfcBVEd7
tXACYUwc1fll4LOj6vSfT35erVWAPoJ5nJEWYcZjH68MlEOusY/5zZjWg82gn0nv
hDVAciYiZhcLn0EzMppRCG4Wl/+f/d0U2BOm/MFKnQnuHUywBpTcmdpWJm6Sp32s
aRrbP3K7WSYFm4a8/+Ye6L26tqCjM9kCLwussSM+Qg8nUW/x9UkU6L8KlNZ8vGRw
TkJivtPf5EGto5le3McONFaxf/MsNTFU48F1JgTgGHZ63u9XMyzh8BxXKVbU7JyA
rTUsT4EvdZdmw9Fr4jT8mLTZJVVlnVgtG3SPYNl2w2EtI/eYNlQXxbV+1DRsgRXM
NaRpdC5vqwM/RL+Rko1jCc4nwmeeLBDTGJKgNAmYWQy74gilMeBO6Z4bClsidJVi
sldgVM6gfRAiX6WnYjtJz45Y4iVJozihG9SW9/D7yBwZYgyhlX7ksxNJ+CMJw0xt
cMVW4EgUjIATchPR5qXNBQVLbQ5FvJGIdT3Zfd3A4nEdLcy9m3qoZ34qiFLUZI4G
Ydwj9gtstxMkRWS0SP6yaVzf+xFmVQkJtx2yayFg7SekshcQuxxAZd9LkGaDp2lQ
l9foVm0OyVdTWEh3Yh2/K3LQdnLUmmiyTPf/Gb3+VVH6E10Xbg5mNRuzRV+8hBET
kLvRGHYZ1Nq8jiJx813loADqMG5rPq39i4eH6Y8JNmNMh7Du0kSHUjJ52dAREVlo
pPSmG4vQk+0+aMSk3yBhl+/J74UzkcaprSEBcLU1HUjy0jt4mtJo+gYNKYc8h6KS
458vYx2Tt0nxYd1J06jhQ3kVPC93O++I2VtpL/r3oqsbMcyo6ZMrCsqeA04Nu5pX
/2egwD6nvznTaZUTIAqjxYCIoANXXw2Mya+Kvv1d/vdMJ+MQOoakAtGONtXJULw2
ujYoLRoieCZNfXKc88w03x+DKZkwrVUGurDGw18CLWesRJYsh9+d7PKIpY5UXZIM
jl90N5DhnlS/SNqdKdFQPmk8D3JSoA/uH8a3MW14WY8TEVa3rQTAENLOzQZ7/HY8
56S6xUpuwZ+rf8wGgjnbAwswp8sQvYSO48lshjy/2+HIU4gidBpXE/PZnQ6kEwyk
kprtam1T8tVoz3gsx6uvxcWt3Emdk4ZLo3fVHwWCdxyBkZJdZh3F+UCbyCkKn3m+
QZeB5zSiVuxu6HcYc8CUeOe4qjH4abnjcUvoHyv3TxROCxJtx4IThycZjWvStJ38
AFPmXxa9SNje4rR7YZo8UJksdHEJ60dYFLZmEvlR3Z0QrzA0ycXZedH9X9mTSS7b
Hb5BeMR2K992btg0vg2CjGrVUhZgmCoavhxl2zt2wuWcidWQKRZ04X6uckD7YFU/
QOS4x1gYqByyvc/UYoeGeIjhlE3EmiglErCUhcF9jsRTaPjDd9aQ1lBQUqS9yX9s
J1rCnHVlA3S7FSFrMJWxfU+SENL0h2H5mbFks+S5T1LmNx/yKB9o2t2aiYNgTgYr
AVGQoJpHwGDsUvRPV1JUXQXDSsrn3GuzpJUccMWf2nFncP7bBQzQLaU4bbAyed3R
mxM1VKGv6Jm1AnmgPWb+8qozaj5GxOhc8i0gNCX/St+ej92zoFKM0SRpEnUDapTe
+AgpXcsxNXaa362Zl4GrKLtSLW12QiwHbPJHvAm5Pc3aRLLt6nV+YvOEAS7zWLMB
bsxSkMOF3N74qU+gGqhd3X71rN1G/BMRxuuXFBvjEncRFM6Tgji715l7Fwu4Ji/V
fqDt26bEbxC56IPi1eIEwOD3/UP6cr0JqbNq4PJS8a1c+f+KLgQ5He6fPX8VvD87
OQsziYcmUSH8sEUE1OusvscVF6j2vRNOlA/Sw/BybO1koidU7iY3AieBQmZvnXyc
Ad7ru7j1wsEoh9qM4dmqio6xvBxPyAURCLPEeElTXKG3JNs2444k5UDi2jknWHXa
opON9ySdPkdlnDIGPdVcNKH6AFg4dvoawqsalpTq5DNPE1yXFlasRpEQP12sYcC/
e5BBOwFeDZbQjWjv+2G/GFeTTNxpxH5RH7mkvcJDV3JIyjTwjcpkVZhf/b8vLsTC
aNwvY+68YZnsXamH9o1345vGNkCaaAeBJYQOYxxS87JDeYL16Y0fvg8A9af/yQuE
iQdUvjUn8yzz1XSyZrWFXpEH6lK4KJp/YyTWFcD6ScVMFkSniMCfp+mpOaJZNyAd
qg6MDYTITeXrMMVqmpPmG62Y32/2+RFCbzNIYcuHNXI80KNHe59wavLqdqv8OQWL
QcY3nA6tp0jRr3LWXTnXhA==
`pragma protect end_protected
