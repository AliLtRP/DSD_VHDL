// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:31 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
l1N2gLuSPyl214v4/UInADXu2hq8y0Lyrfa80nuBZIiouJdrUhuLlrfUX65ViBl8
IWjBxEZMBsMNcBsYCHZwUX3d8mRHv2ZUmek7ZNqlYV9X6ap2CA5sTtHBNCCcaZdS
nateucZXYLsLTUZSfMczqbZrCUme85OxTjluR5y6KvM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19088)
sTa/G0sVp8tnUjqLBlmyqhXl7bKYvtBTZE+8ylVpntRrDox03+TiUULnILsCU5vQ
aO2/oXpTFR8sMuKFBMmYCuxiHbXhPtdwxvBCymnpCBgQX35W5Z657ujcs/MDLs/8
lAMeKHJ9cN0mXWq1SzeYqXebuKdt3Au3bCL3P+7YvCSdbl0LoWNq5lQyux634Whh
3oCw3w9XpH9Js+qpyUB4nuu4AnmqjTa93Zg9GTcVVZZvpp6K/PYQpep15j7hNqaW
yUufG3MDgdCSL4LKDUKok4yIpMF3D9oSo/7oCwjVTNNkRzIfRAhXS2maKiSIv2+u
gKwtvDAaRXfzA51z4OWMVm5HIL1AGWaewmmg7OjmPdcP/xPKfKtPHvyIEvAExe6Q
c9gpa20ya4jzXvIWvWjWLJK4k8btZvV/7TfOZxWZtFH1kxzw8M9/ctPE66bJIYZu
AjRY7HASa+HH5Q+E4IzEDx1ldDLLbtFhJRG2QhMPAcPFTsVstJfdLpe5cW2XuwCK
r+pyHNPBbZEZjsF5vxBM9QTZ/q34hxakHZgSZNN3ibSSjVudoLFY3qhLJ2UZkg4G
NaCqFiIRFLGe0voa9QF3H2Q8DFsBkYVc4WaYAK9ciZYFr2Q2J6JL1PqelUAuJRiX
cOCtgTmx+yLs9pMj5fNVn3C5UhjrrcXIAYxCLRyvtBTQeOY2Kpb7oDDvVVZ74VFt
g9IkrX6nV1NSL3OO6sGRQ+5Qdp1qRB9nDuaTsYQeGfAO7GHhWiUsymsk764Xvdbo
HJZDC2sLq3KMHIfwrHn5/4HIsfRNz07194XtkrlfPPxaJgvlVkr28a824RyhBT8g
Yv1AoUXar73sOWHUMKR4lMPOgncZE/vttbEjDEHZ1cYIHaqsndyR/M8c+mQSQ6sx
mve0uQ+4cQihjh6jqjMJW9TJRW7EY5FLfTQKK/LfIKaaN4eXzJQ8M/trhDoqvWna
9s+uGSiJYFXAeBvVh9W88neXudLDguHS7XhlCVP0tGUON3gm5ynS9zZd8xDLFJWZ
9x4Umo8c8s06ifarhk+RVKavVyB1B4mfAO2F/rpHq+RI1tM05PUTe0BgpKSC2HNQ
GlWlYjNXL8Ima+4oopCZwb2kbpflXqhJmfzilsX5NY9/nMovXSefy5kXBOLVxXrC
BI95cQDbDvrZkqkspDTdRclk9Ps48a6Z47GI2ZgFPOR2/eIcN5Hxx112T6GpRkQn
jh+bu7JOgK3fe4kQ6hhQOlgw2L/ICmU1bLIke+otrAi8Y+wKXN2MeCFw9sNsgBvs
Jg3hHRFQcnMd9BMzUHEhqxS0d+UwyZxIzNS2Sx4czktmVXW3CICb5iZNYda3XFvN
/ceZhXhJoaY5kucoQgyKkyNvmnYuvbS8JGkyRJ/3gAXpv9hxPFXQB7W12ngHuerg
8QT5NZnNc6BR+z5n9Mg4GqnkM9jVgWyDBiqG1D0S2/ChHgLcurkK8s3DwVYNmPu9
109A/EI4pFqn9aP6Hm/uVstjO/d6LVSpAMPHTda+06kevu9MzKcOci9Dr6RY7u5L
KEg/FqdzHgxJx+bXGbMCHfQpFI8b1Vmzfz/syooJywdNfYjOMxMrYra3/L6ruMbD
Tu30c4vZmBUsoJcrcanlBAh43loWCwdY6NkZVYSROEFIBZhtXY6xCsxTSlMxDry2
Ju3mckBvIiTs7Vcn+eS/R6Vcdf6/bcp96uqzVqGqYu1Kw7ti+cEH49XJ7bhV3Fuj
Zk4yg9T7B2iVfU/5sIn5Pqmb785lfC00E8s08QDMIBTrS3WuQy2k8zL052K2d3eH
FZlQGvF0LUJxvVp0ciMO+251s1Xx+yIkJL9unYLA2bViuiVW4wJqQhQ60FPVGTZd
MbilRkGy9t57euPDo7eqejw/gdiMMfmzG097Eb+pvJReLARjanRYgpgFF7NDfYTh
0/78yUnDpnn9Neg0iDVnGU7ve0OhRW8bEwJmwRy3ZlFfM9wZNTgK9/apLloCNScS
0QJH5Fn1QITdGeZZOowMTsYT8X6c9Qb30OIm5VPnDFC4nEcY33C65rlxsXTZWA6y
SA3jkhQF+203u4h5WGndynIfEQlyC43wPvLIVsB/n7TFYlOqSBJo9KicJgZtQCOK
Fho+fu963bh5qWxMXF/CbRYcUuy4Lo4NMqrIoKq978MdVlXFLAxkf6q4v8FhHVAZ
Q/h2+MxtIQrloIjCROz/Q4NBtP0ZOaTDxAnQ4i9bDM6thIBdtCmLSGbbZSU2Zdj4
Jy9XdkVVC+Ynd09q3UjaFxCj96EIMEbzzxTAI4hrdm0xfsk5KY8u3BT3Qjk877gK
LehQFcO2URNcZFnhNocQIxnaU2FjwSCkr+Z3uE4++ntcPpRo9M/u3p+NCC7QEgba
gdSyDFgsXwITYmP66ucklsNemHacPWF9el/qvid6gBgI8+NKf3jTnMcvFHwVQIKQ
RHfJY8uPyRfIeUNdqAgwWiYbW0zzMAsNvpEBda1gmyYgKZrCS54QWXYJ2En0P706
nzjelasmMF3WEXHkXyQKPvB2uhqH3h1VzP4AczGPb/IBjFFMH+mosQvMDUyWpFzm
GPlMoZQZUHZ2ek7HM0w/DGSDYXFlERabTI08MjolZetXYieWwyXa+Lo1GhMeQCiP
x+mcnNXKDU6bG2ZnGxUUfCmyB73Tb1zkOVtxHPTQzkJO7ihmiTvtP9vK/6QVFI7r
jwv3/gJeQBpzPBlSahn9T41hZhCrrlKOUmTIiZwg8TmHX68xj5eCVCNGyQ542CPf
+tCt1hQkuGoSEawJcX8uRDJhF8Hfdu587sMA2FFTZLysNE93nKsvOBc4Br9kAVde
3zPl/rOLTuDiPUwfYmQ5YmQUVK0NQ2I99Sz31xaa2ApDEHSWGeIRSbKMRRWox3My
ikA4wqujvM+G7OYPOHo13bGiULmtv+qHbsNvlLaqspjksDW/G6d3haZ5LeIALvV4
h8SbrLuf9lockMlQhjaqwQFV/zg/qt0IDpXcBElFMOkfg3Qgj8wz541VBC0jdgLG
rEWx+5RFO/oiNdRMcfTpHBjEucoh18IJ7DsfiJs0TgHXwssAyIiGYrqQItC6Tc7E
hTMLRKGiwMwCTLNPhUTOKD4HIbetOGw4kP1SGSHRAmFpl4rZ0aKQz6Fhebw0w0/R
KSKq5PpJChS11O5y9R0jZNlDo1c2cVfJcMAofc64hMXoFQpRTIr+vqk4QIv5uv1m
2NC9mg5M+K2hnrzwAprt0ZWpNPaKMIwJ+8w1BcPIBVSPudNfNDA1+KVzAVU06aJM
qLdXIqiQz1+bJ9IWAQ1NzYjvshWj5Eid42MyEaa+QZ3Di54HnQcrL95PN4VDh8bq
WvoUVROCcDXq6QZYaKVfkSW6V5/x4TlxCkZjuiGDklx1LDqHz7Yf51CZtCY4j1U9
ee0HAwy6yfIwluu7TappocEXi1KJeCPwwSdOCbqR2K+DukXSlVz8sSp1H+j/KeiA
ZXShpJlc06HMVakuurh29g6nNdezcnQ6XnbVRDzAM427CCqtllSMpbfLKRBTcIYR
OD+De6bDnLcMccTT6qTiYZivser6X7TLsEXGoLE0RBTRvNuNFFPRt3Cg0qxLRfFu
Pbd/gwE4+3e2aGha64mqJEewxN8/oyGiyWiD+Xc5Xfa0t3Cmzoqk/FudLTIByiBv
M5i3V+ebrOnTeOLTKdlgouT8sHjBxVlY5jy9o9M6ESt8j93zhfLMZp4CZamCEMW5
x6axDorc9J2OV6qUxLIsC1uqeM5a7XlYOTHHmh0aaz0nYOs4+Le4Vv/2rloap0Cg
4G9NKL5/SBDhP1RYtwF0z+YMJwQ3nrMmefd1n3V88LK7LoAK/Oeyi2jEH2FsLgOU
Qa+ss0+aehH7Jo2CyazruBgeHp3YTZ+6KaB2HTZ00jxxs1xrpwbtrmB27TGWpCuJ
ctBbar8zj6eOhyMYuAhc4pIWLZAM0QF1BIJwDwv+bJWU+v73WHUJGzTaTWQgprwM
V+abD2fsJDg2JQ4gcrT7hF5kYxIj0sJEoyaIyaaD2pbGxUvsnGhZVrNf/FPL7pTZ
9u9dNoeZ9q6bviZtwvPBlS9Ba3UIYai7LQ+Qc9Q1pLvbflX+Ep6fvse1mqqeQSmP
pcaqwup6elGXS/DjGrdDg5Z8spvIIrhvoEgGXoMCAMXVgNe9il2N3tbKFFz1/ZuN
w1/Y9K+coo4zF/90QA+SCzvGWi1SdSw8BiQP5U3a7QAfY8H5Xfz6lF3aymRIddwR
sXLuIbCvz+vO501ty7NtJf0YkWu+eVowesTS4Vx6WEWpRV9dDhMc1/LGMjzCKPsA
LGoOlwyQ+G21DDOQORsXjM3jegVjdvYnMg6F2B7feU5MS8ZTtCgzYg/SIhQ9a76a
BBIAu3YezoDOkyFt1ixj5mcc/UlZNQUKvfqocHgJYWr6YOleD55WY5o90vvn8hno
Jq32MoSDcgFf4QGWBdrtJ2SG4w5tZ6VVSV9j3AndBigCICID2orfQjA7wCRsPg37
NGgVtvVtnBz+iUPwNktokY0dcZ6KyXk3CUuXEvGJEhnyUgO5toxgV859vxHM0Bqy
B8K7NDPMjdb3WdY/s5XfFJzX1TnhgZb5Ttz3euucjD6d2ZxVCHdsCjFj5CMCfqRD
KI0+j9nVHNbZFrJk7fDoyH7UKrAmBFvPI3rRzPL6X1+qn4eyXhXI3bMEvqEoNeZT
awK6zGCHnmgwZK+klgHXZYGn5vy5JqWYmSbnAei72fqRbOcgMpSiHGR6phdIAzNe
HYCsQ4hB6NNwjFMKIJauIaFl/Zz8tWYNjAerS4yZmFvivq54QPHIYFqMeNEwNk9x
biA53+G8X9ndOeLJ0pN8zsGk1h0cDhVeSgQGB2QLJBagy6OvW1hIuK/XFWYU0GAg
1+CzU8Z4Cf544IZKY15s9QSgxWQoxOSvAzgnnMVtFyHbf4Qq2pu7c0FiE7vzE8LD
CfGMHPd58so06KvHl6oRss1h4y/MsnPmLTLEmbiaAVrUqOVvm8X8il3DU+/v2yq8
6DMp8UnKNlgCGNTfOxnUXwccKlvQ94NfnN4+iDqm0XDML467Nrqo5Se+hNtiuX5K
k1yE1isGv0laJ1LsgZEvRITFBjaITB91q0ZC1O80cshd4DH6DlsxFGD5chClQtUk
E1myuRY8Ae0YUZ3XoDYEWTpxK3OaDQgNqEekq9gOp1VUoMrYNFs2ULmm5ILIPUtU
MtwrFjQLy31BtbIBiq9LLnnzbu4MzDS3HS4D+s0n1gkYmGSgBPTxztyn0kKulhaI
jJXnGT3H7BOy/7CGnPx3fkz3jQRktARiwppiizJe1sRlALcpzYJkvr1q5be6HjRx
sH2YdvnyvKgt5jDdCe0djIj2qogIuxbmZk4PLnVxb0sR2lY5tVQNk/YAwIconH/N
5FWJ4e3gekkOoYIEBHXsrBmOiCW9k7wtR27n2LCnGvXwOIQzkH6uoId0iTiTdCUB
aolLHuEh9jf40wj1tbAt7gPsSphcl2qr6cazOfoAu3EYDPFQjyxnsEejpjjc9qjG
7DuNmmJgE1ZUiUSRgBGbxU1uEXFDpGu4fkGyehRfsbHyQxFhXqbc0gSn0g6JlpUt
2xGWmqMTIFj26xU+HXCiuCNksu77oJ7qJWEQr8sNCypmMUm4Bkj3v9RapsxQ02KL
4cETy17Va7oGhpSqUaQHlix9yw8TIhj2ZvPTeZy6oBM3zpVJENzXMsz1ywq3x+XO
y6Ryk7npSIiiAFy1oAS/oNrsvlNPdul8KNtWOe9Es3tSXUAnddHwGHHaSN9KLU3u
wveNn4dxBymGdq94oAWWWsOtr1hEse6m9x+VQsgz59uu8QimNpeKnEZdc5Sfy7Tp
xeIVSVjfuBjV1ng3hbdyttDQMbjs+plrev6E7vuO7Reig3VwFdLeYToCr8rPNGsZ
t6QSMupuYRXduYgGcBbDwIbjc4quEoWA3ZZkd/h84JC7QPD0SjjVLW9NF4L8ZeV0
oVujLDUxqDOQq3vyVQJ2DAB3X4+VBjlslXd2HThimquYTTfUG/UgQCx42T2PRzo8
rnLG3Pf5IJw1Mz3vI+bKPUZTKTAXgyfPK9t6WEBmtjX/qpiOP+Aw5J+YQgpzalWK
cLnDJ4DCiChU44hKG06fxESOjNvqoVH6EPu1Rs2brZCBA0FqtHCx+KAieY7aDUAp
eZDDi9+VaklOg910FE7191bPdhUyE6P6PMnnHkCjKDpHVkQIe6QL4GVBPrG8Fxcl
gaG2PuDAZfyM/XXyEg8vBh+LbTC+l/1Dz8vWT9RNV6ginQPAwAGJGSLAQCDm5Zb5
nUwTT9zpIRzi8WrQ43viCZgzt8FqxG+agadYSJAR2HYKNXgkJKf37SNqIGEdHHRa
6FkrkDaw/wl42WXYHeLfLPjnHbaZkOvoBPbf2V6CSWwjsizmZ1RkCScKb2cQqR4z
byWNsg8/ucTJd+WQWPpOP9WAAf4wAkheH5+03CcyHc7yc8wHs45xqTaU1VaKZuso
VyhMZ4ESb+3xbRM86ca0b2UwW7Yce7ZoeImrL024HTDIu+oaUu1HI0+n0UjIqAA1
z61fNbev38uDvjVbDtkEaBsotP1oyly8kBQVb+9OaFMi8PeE8h3l9CSNbfUCTjwO
zpoePTs5lUrmQ6kpcemwHCj5zOD1s3V8a/RwdDvrNDjqQ/m4k+Lkhz7zBTbDGeEc
BJC2ESRQUYK+EmFaqecMhCZ1JfZoKcBKBQNTELW8jVBtiWsfOd6NhNWxd0mSWYU2
aQZ+lNma9Az42LMqBdh61IjxHev+4R5rgQKXWml5RtEijz3BUrERU2arwEbryMlJ
6LjY7B7ehm+MLGz2sEsTeZWVDJs5qIMgVG+ZFB2RAJlbQyMKmuEeCEi3XVWB3wAl
1qODZUIiK1K3wrUe8UCayGs4kOrDcuTDGsHiu4//Ndi6N7+kmLBUPMOOc6HrcxtN
dfHznQJra9LvI0oGdOBcg4oo5/7d2lsC1Yh8JrPjhG4Lyb7h9WUbR+RE1Ja1br2Z
2WWzFEvGouUEyJZJdM3hiWbcKR18kzx1lWWTX5qwJeE65LWgIMMpONoXsw2qZ+DC
2dkFkGJagc545Cg87GsTWXqsaTRx1AeRkUijbvN5mr1r45peLyhTfO2KwCqigFOx
LMGQMusKrap5PebKKN8DpyHgGgzo4wwjO1KlHR3JkX5L9t+zWJFAnqCOpOvYuPc+
AHIjLsMtjVGXQwmepa1c7ZWt4s2bm2VXJtasbmy8ZwotE6T0HGVaICEsx0YrbtzZ
jTIAQcKkmto5sS1jLlnesmTfeZ5LEBOvH2+NwTJCIXmZ/Y2rfTgIbhdh3cWe1d1u
u330uZ7RqST49EkYCdp67a4N/xQkGW1fA8QXExDfZD8F+nZrIdcK55CLvFuvM3Ea
3YgUzupGwAo8eyi1AH+8q53uGD5LxAunwXODTwg43nyvEe3J9Uzq/feDH25bN7Q5
Ag6N25PxAFw0wNyyeJ10UmyGPmK3GpyotzN93xqwdf7RnSXB+bZpbQGH97uGrrXX
xEqUmRBgI0j2LEk625YiyQKztY6pjuGp3fwNnxeaGerOYcrM+IdB73vpwOGYGPVP
vmW3BWxuZet8xn/SegfemdGJZbMOBk3U3B+x+sF0/SPfjFU2iH3Wpz5jYN9G1+0e
GoPhAfCmzjduptyEa2m1J5jlmIdh0uid3sFOh2Oz/GR97eBK3drb2rp591wSfHP4
gwTZxHJZNZ/k/kEWoxGyNCTl6rKdzkXuKjjUyeo/NbzJy3FpQjvrHJYA8Xy5H54c
WPFmHrP9wqq60mn0DBBTI55A2mak+b4dq1i3BrM7vF3SkeGhUZ7EzrVfX/NrRr4t
CAczrMFL1zWTJrS2354HUgKMDx6smnHCzJIX1bnhtX6CdAH5PDCWNQyNONNBIa55
/d4UUb5HqQ+4BYybB6Sccc+rg9BvMynBC5E7jXCbq1+6V6K1iUTZDxOKyuexHteG
629MFUXavFh6Gn0LCeDqzuRLi7D6GL7+kRiKI6sw4kEo4PBohm9syfu9q48CQqob
G5o5mZN5Bt/cxplHJnvEleJgOSobLi7r0yCIeDdpuPR2MlM5YDk93IyikQboWW7Y
CH/FldPcTM1mIAFk793Wmjo8WuavH5LiRgcoH+lg1sJjB678wCosMOvsulqeMUJS
0qkfbEE9uNVK9j8PVS6imChh4qwsR67J9WlTSgPeGp0r18UqPBpddLVximY+mH7x
OB7jsPmTcsl86NjMWhoRuGcYNnFha+HdYT5fhwdZFfOhxVujM6pfCMQuewiZZvwB
xPRXuep5USXbZzAiqyEoGV1Nz4V3CWHsYkLEwvVqRqWBuQwEtg2/Hy727pmO2f7S
DF4xGfPNQB8X00Q1ZThBcvj8QABKCcG1Qe6K2GNtbGHHdf/qrGsXBJZ9Jb7spR+r
tNwHHtzh/za09tMAxiZSXUZsWCrkXFb0Thf7VobtA4Tmo+gtv777Bw2qDV1+DkiQ
CmQyZjld1MiA9QyCQy5zG03/vrvK2fquQU9hA/NrmnAhmR+9WvmG/aSoZscHEt8F
zsbQqMbCmbV5vpR862Nb8N9Iit9r6MuefqVhjFuZv/wMKXkrEj5jBClyzOEgOiEe
Agi3LQUKNEc67EOyAPvHm7yxm2VHkVPgqBo5ZtJz46X90hPMqi6ZhL1PTITW4GW8
w1OufDHFMan/UB8cDpV6Uef1wjTxVHDn8N+N/1e0wrsUmgehvR9KdfILpEsMFkpP
jcy/sidRXX/B1Lgi+1txKPXdsOtQDvSqGQni2qcQ6X/ruWkrb0VPiLavBQt3DQ9V
KGYEy6wFg9FR/sofbUhM4Ie+nqfuMYngq5dFdJFCryPza3x2Ltp35TlVadT344ew
DCu+UhAM9W2pbb49RyiZd+L2dk8ivqc1mN1LNj6lxrhsSGI6oJXZLDWTATn0Nesk
ZAl1kVkUmR5bEliHokVaiR8aoroGjfIDxArd/4ImCnAFQsX25xdgfAfuP/ObkWkC
hc05CLyjqVXrXuuT9yETzA7/d0idTWvOyoDt2MGV661YRmXwUiKJSU/oAsC9qgnV
fqCDNOr93+Job9r4t0gNo7rokH4lT+H8zh7QAeAMx/iIq+Dt2vsIqeyGtfXmTYST
8nrQhLmTTuKOqLSQAa0ThOi7bOwParB3JsaFmqxcKP3P08tx7VMzgNzht5V4VCpb
f7PsWsLyWKHVU7mYWagygfa+xxF5zCbz5jlZswrPjYNAHbFk7iK2pDBNkipz2A9V
MSLN6VFXR1Avl0ujgS9erUQYW3dKXgG7XVwLRJXmiBwrt324/KUXLTpZomQZCwHS
tz7nw0/dNerH+WFzMPfVvJz6divRAA+jiHEBiLQ0VK2JHFYMh8RslYJGO+wIa/nE
DBNVWHv1SziRzXpNIAFgyoavfnIVm+sjBap+wuBi5isb1L5fr3UFW78EJp/S1ipE
TrjMZeXrqOb2JI9gnG+I3Z1UgYzLefk2iPUpJbFbfI64Q5pU++wzsmKM7OGyj//U
EKrQ324xERy5f8+VNhlSoNjHjRgJM8uqHNPXqNtZc8IGpUJpplsDVCjJ4DPqc9XY
wX4C06GIcglPb8DdAuds3x2VluEJ+vym/BvBo5bjeDQgPKO8RXpYyk3VRno0Yg+l
j6DTVc38VvoD3/xj6nFh0Rl+GUaS6cr9bqSDX9DUjwFsmJIvcdr7nWi7KG9CJXNZ
3Fv2amX33k8zltFc6M26VKUgZGEyaJhEn7pynBzNoBTVejbURkq/2ALAsEtICgyC
oAzKTcHopsedBEfqb2KYOPCNvUfXHM4zwEQQ+qXgmsd+QvasA62HPYra9rCwgrR/
Ju7l0eANFJms9+LJaNTWPx+SbnIFhuYB9/0MSl0AVQHhNS7i9gS/1YDlVbOfp1uH
V75TMUyVO/DS2Flm9EzsAq55EKX9T0khZPR2tfNtyjnUQgScMvjvyhEl+dLP23qx
O2HMHLdLf11UKdB0Be1fod+tFjrGMe0XZZoQna0gg/kj0RkPXv+qiT2EWu25vrTy
boSohfjM43Elrowcuutg0zB7efIojml+J1+rZNcabTlsjziToInLgwI5Reg7R9dK
d7f4QE6Yze01mD7lDCGWF9rhgqu9HfV4zU3eFyXxdpAk+5v8JGazU13Clu8dKnNf
ZLEZREW3vFVBXPWDE7MY8FW4Y70CuRcAvW+cIlgs7U0MJ2+GBGJSe3IZyNanpcd0
YKKh+V+HUb+qBDCfhG4mRJPa/q2Cup+hDlx0VymeeiShI4bj833pUpebbG8820Lp
R0k0Nshajqx5YkQgVUFNOkLow4P0AGgDMC8adEjI/UVANMPjKNR4D9Tv8KYATMFZ
CHEz5tBByGSrT92Q7lE776h0SSECasc3f2O7upCPyhsg3yrKdu9flF4ZuBfaI2q+
HONAHiGeVTR8zqC5wD/pXvp4g8EVH8nS0efPxcYaYeNY1DDYoNYEvbwlgoGqgWrY
Vs7mO8LmQZ/ohyZaYIxg58iTSpf5wJdyy9C5ZrMc0Irw0j4oMRBrOxzZyV6xTgfl
H+2G/E2ybNksILgkNIVO6TfUaGLWuRmusuX7vWGesQJgBmBS3xO1PSLUA0axX5M+
Mq6p2VtJRUwWZrkK67YDjeWbd0LGRkPkSnDi8Q4Q+0aVA0rIrm1BdIBk/meV6/fB
n4ef+CRL1dTlwFwJI+d1HMrYQjTrys8kUpUFWh+XkTQsoWft+JLtuOKmK3rwdTY1
tTRDIWxfallUMBV9DI5C6aZUgQuy2Lz9kIPnJXwJ7mEBZ5GnpZHYtt/tyOh/UmHM
70eMsQensJHvUr3DDkdExDi/vvxi1PZRRJ5Zt0yllD7VaWNFweQAInDdYvy14brr
d+EH4BaZaut0PXG/WAUU9Ir3M2grG2uuLXcXPkAYjVqPd9RJmqWf1I32Q/ScyErg
cr+zokuOiTntRLPnK/ulhDRLU4R4KT2WD1qhkkyaEq9ER8fzAHPOmMHF79fTZGah
hd7Tlsh9U99cie6JLkzNzTZumHIbSdrTfpiAndv9yxyWd4LcQg64YN+4jmwNHl4p
5l3B4nbPVbwTh21YHhEB9YmT8tnPv2E2VzD47BkBPfW6pCCFbJwVYQLb1vhZseu2
rJtU7awjzMqHtf71y/TEeFzifU13w+fh3QS9oNDqJfHkgffFz9vNXRri72cLS+uT
SOjsADVK4afyW9ANkHNNSWO3kGoatks912XsKaBH1Pp2fR3PpHin9vOxQ2jJhawW
E/wKS5tgBsYSY3ExoPJ6gpgv0jjisXqfwT8LgF2kBvxYoVUq+vnZv4MqNoDLgi2d
GrqVQMaT+/XxkU4ui5PAaLjm2yCHMX9qAjYLy0cGPEGW235b2Laqe8ub7tIbsemY
NxRLBwa6+oJDWAPJOexKaO5/uxTceT3E/i85e/8LjabvSJnEqVQQrvKIgdRfNK/B
9drPr+khgWXr9+OHRFyRj1AAgBXEUx5oIRH4hqPORRlmdzVzSmwilRn2RzG69D3c
gIzQQdm2AVoto6PPY1Y+XYj+Vxnm3NHexyoJdVhf8BoIcOHfyErqwT+MjsafjWZP
x5rAYKmndFtEM5cWuDyT5Yn4hcrT2OOq7wenRKh84j4imqepy4dcFUzKOad12X7V
rlkgUB+uplaz3XpKaoCMCqWp/Ef5aDVhDipIvboNOoP//b7E7XSISq3ZzwOnpLHD
DeAL028fHo/3AtFdGZGpOPSdRbTdLbqeTooyyi0Bxt63STeHgZ+wzYs2hc6/zL+Y
+RQsjYysl+tQhOCV92h3bMcyPcK8MMMMQu2Hzf5nRj142vAMTLvh19ui2gb+SoLP
M7q8cksDoO4wiYOxRyfIl9YnOFo8Pkj5Zq/MKxlLd7yZG3ghYCGjgp7nktcTcMPU
d34+lUX0cCaC69ntI1QIoC5z9pvX8cQumYOw5P2yUKaeECBq7OgruqFSwWNNK/b4
zTn+ZUCEVrFSXnL1U35kO4ofM+niEWVwRTLQt//dKdzm8Ny4FCaijcimCMstiLSU
02VxeJ9tsQ8eEslZLoQ4/uTCtuSfJ1Mb1B5Lz4YMMQRy01DGAQcqZEjiyG4T6OyF
C8KIcUIBSORB6yRu24KxrGbzY7qzNFBKxjIy4Q41cK4E/VuEMW1ayaZndzgWkb9X
Kop2ovLFxwfw211ekLbkWhOHcl2FjqPRn77KziL4LguUP3dt3ncMUB+0qeOGQXw2
K1eE1KKa8aVRBZ9XyhlkzZcg3MFhHI6EYFKSfzN5CZYQ4cirrNOcfVfYMWL/BPMn
0nB6fBdcj6gL3a3Rc9TpSysURx1fHO/bwq+pXK2g89zamkKqbd2NC+iZJy8Khff/
p1EPZPfM0ZRdcZ0/p5t5Y41XURkNO8cBUJnQaFGy1LqgUedp6H4AuSeo+AIFzTa4
FIi+CwQDV66F2ipGuEdr5FwIhvW2Dpnn+Nlg67ZSMUZcfTVukw+WcS4iIm0LVzXy
T9CjOsl1g2tOeJ3NjMkNyV0DvxskKfpHUwMhzcPjM9IcwzhXP/WDuGS/7Nfb8CdN
ipikryT8YHvf0Kxg+/4MT9Jdi9sSeerNjwfd4egapE+RG3kHSr4AXWl8KyZgHj8h
O1j66ChojtEx77Q+5WNn0U68uDXfOmsbc/Q009yzNJBL+10yOHSb/aNHg3K0RH2y
zfQJRw9+25WjRDOYmu1sROiBcTf2rZxhP8hiy1UG9OOlaZFI2BK1r+e+3LVT8LKS
Z+3wX/YY/dDSH2Rb5iaIV20B/2Yc83u+3BssCsrNNfR65QEQevWC2sWUvKZWaOz7
UIGMAOgicCLrDIDbEILIXhxUNnVfaobHQslacZCabyrG7hRSq89ULZ7CmA08sFwL
CRHRL9hWvJGh2lrXEx4BTW+hNLz0cx2QuVsMnc5ozIU5IyP1wd+5R7Awk8EQ3Va0
kDees++siOf2tNplYtWHUi1eqylAc0LuNWD1PeMAdNaIhOzEINLMu1Sb3D5P1ukQ
AzhWjuBdFfmrt8bw9nXJnJQA5mHjK5mLkY7mgqen5Pd9UFtF81LW8w5Pg7+JviVG
XpmWVU8FiUf445OKqf26uYgcaf1rKMyEp4JL9UgJ8GOwowa2d0DTvY0v4lnyoWs7
/Z5IqOFbm3W1lfd9441F0YRUQMlxGmL7uXncFTKDL/deQCZCzSee+VYpoM0DeEzl
9cDIq3UAXBZy+rWsiHvoAkpjjFgyzNqwcjcB/c0m1gAMXKrfrgQlWDU00rdRFWL/
j52fN0YYYQ8A+cBlSCOK1/bQ/Zpj5zAGRAEJQmv7AF/oBHxo8VZzuhvVSa1+vlNe
H8rda9BRevoaFyXaC2jquSd7NZxx24tOBOL7XxORGL9xKYampl5vZH93LMAX0dWg
Fuun310a2InxQLS1hwxyYmP3S12oiGVBTZ6j/OjGPINnxTi10/tGU6pNHRy0r1XM
MIN9sMn5uGEsiDi2HYXn2N5UCdLW/17Fa47ClpcJvcnNKMqJduSnv+8T1Dn9tEgj
VRVqRGeF+Kg3XGuEvoCpN0pXJYi3Xu4RWMQM9gfEjc4Ze8JzlE9jSAu3qHfrEttX
GBCFRCKFo7c/9g3W5iRbQlmoyObjwIa3XPUDXL2uGdVyzH9BhTo2lDI+7vpDR1Qs
MOsfftei2u1kqsx3V+EbJBKfjFgK3j5hfkywWThKBeF2hy55zDgC0py3PoHmqKPM
AjsWjxBU8QsSckciJffviYnNfBtIklnIiaZMJX/MA6K31nMhwDMOso7eUETR8Erd
+8T6FmBLFA2b2x4TWX4oTLJE6AIdVJ/GY58xiQgRgUIzTFsNWc/YYuiXfEbUXXhJ
HjVrbXVr1u5ltKZg1FVbQAzu59eszS+6S/ynQ0KYfFrBR6k3yN0PsnKw/fjkZ53g
druFTL2OdTcdmMSIXuh1HW0dNBtMknsTcE6oW6Iaf1TyU6I2x8MuV7K6jMNAOYBh
qrN9jmj1Xzz5bgE9qrs0j85heu2UQvYjSqocSHXSHbDCh2oHjQWWd2X7CYs8pbdL
3iiqTL7/QmEfVV0GUmWMcxwtOTtc+xAOEk01w14/0B8cT9qcP+W34j2c8wptA8kk
aw2d/CD06+cCTAybSge9/n67mb05fjcZ0eNAnwA2mR/xbGsg7cyISQGFib6rdP2I
swX3OyQ0HkxiwEg4Gkx/GV2z1o2GIq5dUWJjvXYHNxZGma9V1UrgljTTF04hDaiZ
mqM9Xw1kiK2CXrxA8d6ZcrAX2Va/GlkCBmhzTrafnsxcj6tscJY4V2P0JiffrmE7
WHPGE27H1FP2NACGQuxf5tiXPpaPCxQClVdtQhJ39RY0yDAJMJRP8qG6K4YrylEi
K9nG6cpppEv/Ge7fbzmIiGk0oiqMlZOvia463QlOFywVlvZVpPALJmiusAsvXIS+
C/auE3TXo8PpbsmXF+UGl6xeHfKAEkzy2LczQwiv125wDpDTkcX3YUpdmgkkWiCa
pq1+hxRCS/9BVBEPU4YBTMD748yaWdrR97fVoaeYmvRfBtkeyP32DjXxkgVFZfA6
ufYzWVaY2prM0GUHaUsc2AncR5RnGyvn4nPimsWYODr3N3nCKgOBCb8HUd8kqpbi
O/SgtiMGMQRMQVAlM8JG0DMjcuUrHvZ4XVEeUkuvQk8oLByDfrY1Zf5BwhI13GRX
BB/Ay8CKWmxCtnyEutkDG4FEeEy12NIRKT61uy1cAoTKx3/7davBaOae2InxkYlh
q3QD7sk70iFhVHy6OdTJmfwN+k2gss24MEwqJnDRG1VKXxpuFdQxQCRQl//E5vaU
i3/lx8DbKv+Wa+/ytG1g0/lMZP+s2eBKLvG2KtmjMvZDNgy+87iZJoSIlzE4u74D
h+8uFDEaUEY2r0C51p9jh1GzrP7P0BLXZgeaKblvAWWTyqVOHE2tkWs+yEXxFv9g
WdL9s/kNsPEvEFEJ5e0qKsAi9cN5EWMX00U+kGane8MD1i3giEkXvh6A4SD1RO+x
7lEZRllSBfAvksUIAd1skZFXUf5rq7OkklDoLfIHC/GyRr9jWg0nEZUAmmLV6Y35
7vuRdwnNzsk+YFUSpnkELilGfGTCz+0518ER1kF+MTFPFdVhG/1ramgb6LEOo/yH
2IhnajPvk7zGli7VXI09y22/hcA6o98PaVs7eSbXZU29nrHWTvgafNQETCFTMYIY
rz9Vc6vOQpoHnR4I8XaFQ7Y48Ya+PdLfcGbelIPIKUaHnsypkKws5C7YfI0amp4r
XCVDVUbIc+VnZl0wkjtoalvUptB9eANIS/3sIIdrADZz/OFPB23APf0Si7zLujf/
LlmVcWsEGPxzTxflgPsIRodj4YeSGneObhag6lGroAIjKQQHRm7o8D3Pb9QXCDD6
gWVZksQHyv7hzv6640bXABVdDgI7HQO50rtfI7LQ//tRUPw1AiZV8JZobpNbZm9i
rIsmPmpZbOqvQJsKrbXYCO5uEAc15udJKexVpdIdGXgFvNI6c1qHSWg1JOgxQJyG
/J/tOku1PmOXYaoGkjUEBEuoDEfSs63pK1AsfMaZ+EekRczP0jydn3q5rwHOa33W
VbwljmgQ6uS0v1QYIko1sBI0llweBNfYRWU55n9bv92F5tg5xTf1eysc9U5fts/8
ZkTFnzxO/Gqty48Swa/BaKwvEAz8ampkMyA0+mEta/FOK2efzqSgRAdRdIG2+qgJ
XPCjmH+Zc4ftgY9PTGYlQo8L2ei8wy69dPt0l2F2O05Ka8CqNBtwuk1/YIs/uVgX
z/q7ks5jiZE3SF3zq6be3PDVxrUqgmsUdXf14bxq6A6se+YPnkqcvq4D7IkJIAsQ
R5EeRWNmH8l+I1KnIX+vXKid2xrcYMhW1kwGyQjJyjMkeZq/Xc+US+dRgT56+ASQ
lj1iOxST37/ZLdrvB9wlxv/jWtNfUbJqOnyMbpcLw5DAvnbU9IlXTkTO+BsTUdzj
Lxy2G5GhF8TUKHbLoQqNNAI7BMWgs0O2WBN/XssR434aifN5BpaWoJ3ZiHI1fFHY
kLQdGcbvq5vkc+Ps1NNtYh2pnsCZc7zXEPfx76wgEshqxZOrVVQYt05hfKX55VHw
jwQJGhzCUuwR7zsFPaKgJ4kViOrQrsvIsedxOQDxZptUW8CoX8nnhSA3OVbw3toB
Q5ZTpLxsZ9UsPIo4C5Bggh/CnSizKARmQ14gKXoi3kQn5PuYtdcV0c+PEt/WtDQp
N2v3JD5XDyd9Ty4BL9bYE0ea1u0urTQilQYHnXvoJhhphDqXbsA0YmOFs3XYlpAh
bnszH4AwLs3EkMDglqLGsdamucTcFURNmT/T1Uw/qVa2LpMirsc6ECZshXNaPSz9
IOpEonkHeu9Btd0+Q0VQlx2csuy39VkRZkA8w6WUPRYKvpFK8aVWcakAvXsEVtLJ
C/oGMshawEStk1WZsuhjR6SG8VH02gwgPBmXjJloL5T3OSGsGGJPJCMRiPtbDgbI
milTdsXvrlNpZdrUnzeznzpZuN4aUlEJsvkHWb84lpi81Eie/DsbcZLrxMEOCrjF
iIoZZQolkk4Syog3SYdfKfAWx45Zrm5QVv/KHVbKMZLD9zFNY/aJu4FqaTsey+X4
1iUWXciKFs/ZZ2fVooGWpQPZ0y1cyTPGmV8ZvhCx3Bkx7EmLYA3lZLZaVFZKHpeT
6n7Oo8vd10WPBsk59F5+Q7j8+T4SnSeNZUZvRZz0MXM4+K/4ZLQAdMdpiB1MuNgh
rXwgKfi9vLKiwbuQ6CuIr62GGJzTTGfHbD2chFoXHnujyUyviU7Yr4k/TsLdO2GR
iqx0mgmWjb0Xa2gUZT3LON4fn5kXj5hmZPAZ8yPYZCE3bna2D9pocolTmdT49MY6
/vcrLpnMLPHiYRPbilCpGhrlJyKB43neISL6BQiOGxYkATQh//YkCpJBaMtBvlkx
JjCmYR6U7dhUJzRTlZ+bTn8II/5MUOieklvRScb63psHwpLCxlQ0QTbcHdu0RWRv
qNmJazXhWffbGgPkaDChCSN+w1sPrmRc0Ww9Cqxb3fCmOUOc0M4bWbI7R7Hjy7ZB
MZvDkpSsyx1ET1dKGqDrzvzROlmKHj//3ok10HV9Hjmfzp6LVxTzdsAqaP12W2iB
aK8Ozf0ITswQC5j9K4oK2C76n/nu8nF4kHmxjb3yz3HEi3bfHemNoj/9HT3ZP3xz
M5EhURidyql4pu7ef37DsjFlQLZqVWGwjPfb2rOVWBZjIqX/le8zjsGJ/r3t548h
sve4maJ8tbfCRkw+0qFMVKXk/QrrO45nsPN2J+cTzbcSN63tF45M5y34nJSKo8Uq
F9lDPsHS2VyJdXP0yLbdf3+puTfH0HUisgl0bs3vyQGWZDtivaiH75/IdimOmjFN
U2fg3DLyT1Be0kOV8elLiaSToJwgNjbKSHIZ5FFWJ0y6y3j00RNcPblDoIkw3RgG
rUbWsZ45hVJXd7gZfdxtww77SKdt088DBcgxi3DBXRgrxh5l8/YQewgRXi3+mYf3
FCN3fiFLZcNy28NIzsKD3r516L94OO6cuLATkVAdtfS2yKpxMlfa7FRDkqV2lBZh
naKM+p3eueeQ5H2wpJCZitu49IY2X+rq0gLoCJeDax4bGGkpJDe9MgXH47ybwEDD
JiMwII+sBIChFEMDB++XM1i+xLzwyRxFuKwIbfmFnJRS3CmC62yDudhr2BnJIvnL
BW2OwiG7sMPKhn3oZ7q+MKkgc+P49CH6ckVDTgpUzUYOcCEqgeIThJn6EqTuIw9c
LxPJkouo0AuLQQaf3mE24EJe6w7HhTUOHPspnZ9bTbh6tnJMmeHsict123DcAMhN
aS09RQ3BOF5v+/vGFU4wD7edDiZYvw3jkmwt9Hu8moVedHdCy+55JONsuMFzVTls
tEVlkxUfCUl7e0ZYvsYq5CMFfkDqA08Z7pMNNnwpS6+n+akv7UeEfelB/KF/BOiz
ioTnz9ZNufXeVCI7VCLv+e2no667/4ENTPG83NtrYJRP4Aw8WqXcVFW+IPWdBCkF
I91a5e/OYVr0jtDT2F2KkQ8kU5JY2jdbW4ZhYbUy/PG7mBRwKZu3aHYH+YAHPFbI
2S9ilISIdb0TO7t31SzvfPWNQOZ510+hgaUAp4LJztxT0sD1J5bBXAvOOAOUkwMP
Der3dk/bMmzvqc4nzOEsoR6qc1jL8aFqWlCCDexLobWaLUDrhKrHU0wrTmUTYlBc
iZHT18qyIfwpLLpHhnqJKtzyUi0SG/tcp9zWlysJc2Dzgg5s/JWWXDu1ylMrHo3u
KM2vPnUXeMMIVAH+yjO5WRh6nOsN+0qdev0GwV9dSrJdHxqLvc6l0iUKqOw4MVgM
mFezbOv4w72mz3UvHfHsal2zNY3gGZfv0g/iYhPC0I+eAN2DmF+Jr9caFX87Rb8l
g17KydKcrCbgBapUKjTVg+xW+idN54ntiTnc7a8XW4icLbLTJGMOQuIzkhydx9oQ
N49GutGR7OwqptgVyoZ0nPo6HB//Ws402/4e0wRAmqwYTQXq1rrPckdjMBZH2yBV
z8kHNnRibEn3bAQ93ZCkKC9zUVpAPskqwcj3pKqmx+/BxEJTO29Zebf+BnkB6/uS
qZkWH6NoRJ1b2LXu6BJl5brDz+qM2LwcYDgQ7HDGnQXGGTlSmFZCdHhcZMzvYTYN
Pa7y6iwnjIl17ghrKE50aqVUcI97ZGrlXH8n39TXwufyuqlb73LjZ4TZ7VwDaGDA
YCEuSVZwo0LFjOUDfkR4VHpyvl/1q+z33kJOdWwVcqnDrzuT2brhiROVIlBHloEn
QN6VFYbtneR/q4gDvmVDYYika6LxrzAAi5LJJ0FWTqcQ1rJoC1ZOksJWZZu1YK41
SouQrPZN/zrKKsO0JiU/+pmGh0JHTGA/2s+1B2+PcRU388HJIgv/+NicUKLlcMNH
DD3i34/eUsQhXJteGKemYNPrG88yFjBia+c2s6eRZRrggtj6ZKU6yntExOu4jD18
1M/qNY4ETkQbklJmGPfVMd/fqGZLEiQthq3tYVrLjv7kxyjw1w3U9vyqlq/YkBbC
glokTFH+5KoeHATGQLhYyTcNrlE6XK8ImQFt91myUnKTe6danv2dH4G0LbgbDMl3
Zhcum9o2u/W85h2biQF7UkeNL9eXiyQG95YVAWNkjK8PiN5sXLBN7fyvnkaPIdvy
sL/H6tiduZu9csOWBs9Y2FKdjgPkXBOOiYKsV6lKQFQagG9XwXm1fmqPzeAvS5Fb
PuZ0qoC79gU7lThFyiUfRkd+nHze7+Q7lYcT7wbyYAs+TEy33CsqHIoNf1yADpw8
2SMC9NPlBSUcZMcxqyVHl20kCo5I53MEbb1CwJ+U5/9w+Ead11KaO3MnCayrZRnw
mSP5Ud25a5wHXYm/Uqwrn0//mt56XJ1Jsln3u0AstLlSWI7g21WTxkzRL949u2Fg
ZoDP+t9/HX83zLDV0kBiQm6sISAS+tQlhqJy4Q0jjuD7+awRrN/tER2QEtmYHqKy
QpHhGvTDypi5drJMVwj/BdaOAKq6yyTjiI8FqLWCiG+DTmT4kmBv9r6uUhtSLlu9
HFBBb3EC1+WHNtu6ciUj2YvxoVYldD2JURh4d29ZpKRWIL7RoK+hcdA++5MWtGyK
FUoVitJnsJIhgaXOJbaOVHS6/GNP4mbrIEI6Rd64LjW3YobnVNpPdfIHftHNhPdB
c3swQQJF9ktqo2YaJhIciATxPDncr+snsl56c5GyBJUC0AME6PPcVfMQgZuLncVS
hPXd7Gx4dc8Jd2w1NmQTlUOIrQYJLaUmu+K4SBFfFPwGu2tML20j2jeCZyGBDfpg
x1clilOElwYbx9UMiD72xNNhBAkD5BzEkdgzAORIqBOkRR6ZeYJy/RXEcVrk0vTN
Cn7Yjj7291uFQTVoZX0yeN2na1rbG1fftR2i4T6bhWAcn177OekZ+DuE5QEYVPXL
l9jUmQ4Skd/khGoF3ExXnyj0k988wQU2P+DFcsX/of4yuLbIL2DZj6572UcUMok/
vE932xaJPvke4kYk0zfZt4zyQ7vBtuDFI6h3NxHztPedkgku4qeIthhVr6fJMnG8
mwc/XaaMi0BfBobhWc9anyzYlrVPsha/HlKR54lpRPPvPolOjzwaT3tB5RZCeaUN
wZz8RMv12lG0Uf85rebkcPOZS4rdXQGvpo4RAe4XP8dO3mCsy88FDnF3WaeOMfcz
aK4bV6mUb89hzSYkkbxIFM9TbSms1blVTFz2ZKUjwG2hz8CCINnJzFmyDPWom/c0
wlPFpLZE9Ud6Nc63C0a+1PLu0269Gy5oSILKbe1p6+N1qQKETW1Ml6tel33UmPIQ
+HFZ+HSAn9mHI0it5uQ3C2W7L2Xi6c81EXC993X3dRvNUxGAbl2Sv2Hq3wWaw3Qd
qHKYNso2HrLYgkeQci5tEJHLhmzXb2/SEV+yCo5DQdTon5lpaaTJ71oKiwBQWJQl
Q3STI/9jCKm1hTm3MyHrocPaBUHgRoVC5aNFPncNT+Qj/rOq3sY+k677wKZEn+MF
TWxus6Jyq2/RPqlVmNizBj9xe0fZ475r6MSvjUzLXqW1qmTvgddSwrF8GKjbogul
m1tifSR0gbUOSaeTYfggRScXSOatw2g+IuQPUh7lMJRs9UdYD5zT7FhOV3HahNS5
CTCjNCm2IwXsuq6fL0RrBN100pYY+v5MIp6fU0+6wGmKfOu1I3ydg7+OIeEOwaWU
uqIi5dI1OyeYXZofFb/cDhEJjzPRi6s61sjdOm1FZWKL0tO+PjpvdXSNyLefK4Pb
nyyfo9HUUqrxjga4K3kWN2EmMkxRix3+ovwDJvQkHIczKtySHrHcNGqLfYQq6huK
FEX8KLK0PhljIcuE/S3sDDZp9VjfoSwqVmSMt7XMCClaDKMnFdz2ae8UKCwCwmL+
SFEujtB/EN4Z2Dhr6l6oq0C+PmZ1b/0xzTukH6dwIz1ava2k5CBjnJg7EXFsUfH/
ZPq33Vh5IRgmWHz5ikyx+a4GSgqokZNa8lOLNGxnX/dNL+I8mT4NxoBGhmt4qn2k
Jfc+kcCBkitS7gaTghGnU6wH1P4y6SOTefsW2ixArFFdSpA4xq5AnmIvcM/DRweI
pbLt9RepfA/eGp5swgXHZfuKojjOsrnmrQw58iTaGxc9L1Vj/srilBpVoxNihyUI
oq67KW/aYpC9Qq7KtnLyLeqNCW8L9MdP9zDP5zCTDslc5JouRKt7jLaiNa46l+lV
CusNV1YfQnlrPIOHPAKkvKh4ocjX9KLgcjcv8L8DpvA0OpsRuZiNIuf77uVNRFc4
1ovK++RHnf6sEA76/+KKQ1U36swpK3C/6s7hNbhW4IbWoh4GKXL+KnFymh38mTdz
ndvfSBQY8LqJqcNY52dESVjetLap8edWV0Q44jibSf0piMV6ZJuU0r/9uyoLfe5v
9FZixdUoGLamjuPJtO73B5qWG/yuLA86aY4u46D/sV6uSW3bHgtwY/whYYDWF8an
6DNGSfBBgrlhGPxtAup+4rVT7HmI7tRtNuyl1VN7L1tpm9i7tWjTZxqmJT+Hq8Qr
bepa2IuEosTfa3ruG6pf8UU4hCJO6SC9c65yNFUZMeia+87+o/go1njSZ2s2nYUc
u8zABG0vr4Dq5AJoWt3S/u2VNGjaTu3eUWxgp1eLAq9BQRHYgBmpMXU58dcx1U/G
QUYSrAputJk1cGzsrBqajV6/Cx018QC6XIDQO5J8vUjuZPYcL7v7XC6FMy1Ssqzx
U5BrzLroVADCqnfNtnG4cUBwWlniqwf4bmhNYACPckW/8EIkPNMly/0LuN1Y+Asz
yWTQ+dD6FRE9jPQY0rSIY6XtYBheKlLFpeiiitk1ErUGx1mnuO+lKXkQAxBAMyj3
9uJ/Pnx6rtt3LbkH2aArOxLFH1HUUSfhjuBNjPDUFIrywj3BX6wF870fsDJmLZpg
IwET/2DIWtn/ZrkV2hQMX0OSLIYIvY2lrm6j6ZmNgRCG7lctbchA1AMGZkTDFdGU
BUlHhL6hw4cAMsMJuVUXAtGf+tPHlET7iBlyIV+4opIlOcBBRj2vwJCj6o7skbtv
xuRCKgMpjuynn6KMc5X+OlRRl78gWXLBml+Tard806zIIBSpAO7xmt5sPSMK0Trx
p56CG7IkxTi2tIGahhjHdlSYmWaPqP5K62UWuUHk6kV//JerrsridEGcY7eiFBmT
l3w1hsQtMkJ4IHoeRBj7Yd+6r5QrJkZKjoS4B26cgUQMalryvfYJMKTl4Zv4vokL
oClk3rBBpXri5Csd82ZF6IHjkzVMmzuCBU3lv1vI5Qxngkfm+Z3BK5mTOCRhrZab
EWdYhWxoch+Chrl3z1TorYNJOh8FkRsuMs2EOIf68XstEQfK/tUE5UgkJV5Emxy9
79hH5O/yc13CRwF8ylV3Zi8L9TAt7da7APgH816PI9L4uKG1xkSdmitdeJqQXHKv
fXDoO85KIKDdte0KxQIyLdwy1LQJMHBJj32CnHepYXFQnXlHYpwIFfQYp3g8vS70
20kZjmS5EgykY8dVkiosz6Ndnq8CdVeTQLflQWIA9yPF7wechHs/8MNjThdy8DoO
RY62Esa2fMV2C9EmZrPWrY5zPK+VPIRS+CqoqzvV+WumAHjRFNfZGCbT58uw3DOJ
xfDPYIJjJhNuCsUQZJDGema3uKAjCBmSAjx1hBttqZjg//hy2XszVS6NSIQvGkOi
qHt85crFXdQEaFMU3MZZcFT8Odh/W9ZtMHpr9dfSqvxeOflH0Ees6B46KIuGfX2m
smT8fwgo1MTUBRhgcV9w336JJRw4ailG+csL0IrPPqbZcuU6qlCPoerMOeVVrWwv
9YRIFSF9qITNnjCSLwGxXwloA8GUXh84Kri3Vsyajzb32q51G8xMDj/OPuabVgvd
rijGuPNDhva4+S/36ljrU1OPvfOvWov/BCXyzBAiqvh4FVpt+dzQsG1BQ5qsMvDg
3bmYx1AtMzkQr3BjEZ/I0ADA4ag1Dp7HtnAzxr7pb8Y68g9ada86X7YWN9lpP6cI
N7oxiDLRjC6TZsbFmn6p3JafB4YbHdL91pSEIrGL1cdXHsmhaCILz7VtMipeHJwF
/h0h2MGwMKYhNpKkGla2ynqz/tOKoxkWumtc3+wcdV3UvgZDzle1kO0n4Dg+870j
4cRN5Jlfi3WfkErIzwFaJWurpiO22M9wInLtpXKh6glrZfHNgoAcaPgOMglskbkQ
y3fz4tpWLbV7d1P6l6y1E34/zhETnRSneesuc1k9BB+vUyqRTIC2Z9kUQ3eageDn
0R2L5t98r5DUH3LsonRtUquaElszNrfUmueyQJInyz+FUxROj/cwTJHa/pDZYQWm
iYsCmrCQZGxobeHIXKEzVEP6+3rLeLDhbS+h2QG33KUI//i9VVzJOmF0iDjBnZQw
7NoW2ivGn8bMqJ3n1piwkLYp1eqbnLXL24JjV9VTi3CX6J00IWIeJnprOuZ3qdeg
VN4+YpDKW9rgyiZVJV/K6b9SJV0eZB2hSRtTQAQ54pcUHLz2xeg/GSTXMNulWigO
q/G6qyVCXVGMnrx2lt1JR4VbrldmEGjke/njzm/5wyM0f3mrdXY5cKh/1eHC+FpR
6VYAsyXs86THgZki1SqMeppzqjj/bPtcqWLyiIXh8EAaTs4ihaYPYFj5PHTcArPN
sUaaR+kMTS7/rAR+nvl78/MK6Y1JGmCzBho6Hk07/liQd45V0eZ61mG6OpkzlPHT
8K1YBSeJaKmAt3uE/0CD3J7M2O1VwU1Z6qXME1203QCuP/o/TMZuECODliW2tsif
Sr2LC0ihw/2TK4itwFlQeWZXjG311jhA9SaGOPoWUkkp8UI2+Skig6nGtQiJTchx
tEgi8vFS+vvBLnHk+d0LF39ZdgjinsHCQOlnJnjnO7Yjb/pnzR/NhUo3ownezthi
WFstlcCJu9mW5d9Tr0uu7KB2VchSmvATXLD0zP+qkMdQwEGV5hrM6PsT/LRkzt7X
13esvXheR/1z9F4QE3dX1K97tc1+1My18ZFzMMp6oUO+PLd29u+qewbwFkVF9xCL
tJgG1IinyYN4JWW4ttnWJEci77HGvpMNlkCt2CXE/mjEQf3t7mylMXb4n5oXCcVr
k2/ia/dFsVWPPA3/iFkHe7lyd5B5T61n0VvO/rAWe6HgzDPi00PiXENt2/KBA46r
wtOkaQFLfziC8Pfkeb4CLykTqEerXOY4aHs9I85/4C8bLob1x3wB0YTB6OAkUuX5
6/Jh66hN4jwhppAIh7oF/wrYo4t5fpayHzQHocx0jR53uYU5avP9jIBlqA2BxlAZ
wJmMmMWl1Q2r/Dt6yt7VBD0ReUEUjWpMKtm8xf/5c5yAnenoANB0yMWhOP6cQJaJ
BDku/9oqjnARFEKjEC5db4NgyyYorTCjhGB+N9dBYzEiby9xYBlZU6UMa4Vu1ljH
y2NYni8v6+3X7WXIz9pIdCUGIexY8RcUF6illyPDQW35eKm7rWmbWllecqgYvLEj
5huk2kzbegH3nsC/ou+wwnsTyPoHmg/cNXElIZTWMRUF55VraKmS+ouEnjSN2KO5
prrKgLyjT+y9h1aYDj508ChNfeC7bc171ZVri3p9aRlrdN8vo1uAZTcD+hYqVYsU
dm7w9/dSisAz9/YFaxvo05tu1j7JUfusYS/4ct0vBeiIY/tgu3UYA98vokIjW+F+
nb0JGMlb/o1Y68G5gtxRpzuHOmurMrj0ifMk/lFlsLlqJP1ZrGK7ALjCrYoo7SNo
xMJvHn9lHtUBxaBJncRFFq6pZkAHOcO9hZ9eRQcf35Sh1Z8JQs+/Fo/YXjXwH1J5
sDPVxpVM6z06XArSeA6ahw9Kx6lHhqCYjo1RRVywcIN029aCYL7oTtZjBmzG5MRK
Vr7xAqOAExDZX79ew32pvb7wJeKlmCUZd/XTfAzKiVD2QahbPOzQ1A7rPRR5nUJ/
AdNIptjxX29NTOnAIT8Y9htvFhzufu2Gq7uY0rqL2lsqWzUTYfdTBpPMda+cjXEt
HQv+xOI3N0jznR6exhKnUI7y5yHGD8gwJnfmh0KDI1TNduQPwWuo/uXe3IYLl4eZ
KeDLf2IKeIFOW3Kv/8Kd9CaiePvf3ZWg6ynPUCBZlWs9loFN8Igq8xmUJQnq4NXh
rlW+fHhm5xqushCQDG7CuurLUsFNvu7CbURVz/OB20Ql1WSP5exhijX6h/Kzcpx+
HSWjYDRmBck5TAql4oMTXTLoDMAtuePXODdgCHSV56MqhzZjOHrJ3NOyBulsAZge
YrqdQH/GzPj5FCw+PDRFgb+7VTzK+IvH0U9BqjKu2aZx2xUtVnByv6cIZ4w/EW2I
e2znHitXANRInchHXd2j9L5skRHOM3u/PEyZoUiUaMSCdodDljGbjORZbRTEdrMc
/DKZsj8V2ssQ+UL5CwtE3eEgd7xOBpbzUQZmTesmc7ioiYpoHIyQ5VQd5Re9rFem
j3NYREJedSWfBWmYtb5F6jWzQUYrpmfG0YrREgvmSSHp9BVeH5fvOm8plF7xOXWl
G7cTvFdpfoL0njhEIL83u91uXVsf+SAJNABa3AViB9A=
`pragma protect end_protected
