// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QFEOBz5YiKdDZ4WqIMaU60GR8ecla+/q+LK19qoPwOV4S0Uj19x/U3T2qDBkgI1o
LY56KQFF4WgT+1EdBpgX6+9Mlf8RJt9kEjjkrSdCNSk5hRYDjPNX5SBhBbD++v4L
tVpwn/9JA6EiM95XNQMz689XatofL8Mv1c3HhTtEETs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19008)
GhrOAwnCQ2LrUJB+ARJ1I2az78NHyMTpJ48DpfbOGgR9qV4QWMmPVbOTuIpPpfxG
arrrU1a5+3DZL24ZQb/UB3qKK4u7AoHzaQyMoXZElWJTrf488i/Efrp/WFbcHlCT
RflIuoo6/8zurPi+Gyt+pWzf/bWgfTOSc0VuOgJ2DD3LMuigsdUgxtgCxNmD7LeZ
XymaKYOAcSNMgl0yaK5rPZFSJ7p+NWaYY5uTIAyGaqCy0Ipk4Uv5u3ZiIPs1ErwE
M2FyUmYXFxGvvJNNCAMx7nc2xdwlkm7Zn0gCXfiezTo6P1eON/5ZMeNStuUmoP26
pGYkMZB/ChCBO4LMIjthLeM9qErP5qXkSCXss0sTjA0KFa/dWFFqla4Lz1vlcRQN
kDqOg+CTinBVFwf8iPLr035blYVSTl4QKlghmvnWcQiSQfPrgGM/ahE0c9LjymHu
UmRYDVXEemiXPJIZ6sB1jqE4/5IORwt9aU8I5RnGt6IH7b4uLCL1mfFz0zrUrVy9
ZhgMJHGHlYu4CdYNduiql53+VAARlPYDIiIxEDNNanhk8DnkbWMy4ijjxArU6RCt
k8aAPOb1fLYsPwsEEcGgQC5IxAXTwUrBrvqxfhMDi43ROqu4MtiXys6S65bVU1UJ
nJEW19Jn/Go0dYrnj3rsa8IJgeLRMhM8/drX5hHQr2OOyBlQyb+l5hktu2KrfjUo
kBc50SRjvWTEMu7Dv6J70OB9pSIKKAxIBxKhAdYUrB0yhpMlGjr7Aqri/MupFmYr
4CRQA4IULCAqgmR+x69ZCksaiB4kEXVZYg8vcqV4P42NWRyk50zYQfvgfcwQN6tn
eHz9DHQTqOnzGuFB7E/XNnHDQYv+OAxEmI2w4JWX6Cb5eGccMza046XJ9286MBfb
Yemmkx8/9tudUaoiXtyX29ZfJpQIcTpAkcZuqxY5vhK09bJogbTMbQUk22PlFYzB
PZdfBwd9MeAzo55OzdLbIKXSWkRt6I+GWGJSaz2sgX5oeY/PmrWDrwqTNuiVCQ1U
aUJEwWHUOrMc604lUGPDd2q41/WzNgv2oBSwEGrJ5dpZJbxMxiVtt449Viy041cS
tQuywrUAoFOOY9E0LRbbYsaisLL9RY4ZXq+jKyjS05k/SAI5mDZerrlEXffBeanJ
te7/mihCX8KllD7OgtodgPdQFBPdWBgFc5MJGDF44aWI6LFUqAAfaYXlNMxNN8pr
DqrXKmtRMSNUMRt/lLctGY3THgSjTYi7JbFB0FULX5/sWOYnMGLgwey05Mjy8A+Q
gffcPo5XfOSgHstNn2yNKt0Ypbhr4yYr9lXwzx90D64ljhisDoYRat7tJ65SgtrZ
YcWXabbqXid/NopQQzEibr7DbF2Rg6K3xyphHfbwL/1VyOYwr7LgAFqddTk38wTW
k5lWpzUoSb7OBuWuiJhKxyw5rH8BWlA8VwcoMvOOoDGVNznT6xTyu880GV1CNCzd
Y0ORIdH8G7qh5AjF3kHYhuW901KjsKtBleoaqwOvsLoxTz3UUHP58A+ju74uBXTW
ym+mUxmO//aN8vVVUJSgHOGRonIgqHhL8FnDS646Z7i4u9J2EI0xVYkG8fCDlKNw
e/zBdxbhx2LqUMEl5y5ywLQuIhTrTfrKDxY2+fJ6xUIVD2vKF59ns8UTDmRPjCpr
ISo+ZqhZ+i3al4XxNecSNH501uYPHBH5Ujb5d2h/Hj7+/n884tbix1Zq20rZ9vSY
YDjSHp2RQBNYK58CWWxV0pcZEK5eM5FVZwoq16GuPj+dTLhkWyWJoQ3AQfdKc83X
6Mt3zTUJgVhf+sX0GByzQyvGufUS2GwUWcLDZq43lkGTBXV4lDHsmgzL4WEa7+Bf
G3r1JbrTr/yqFsgWbGzOChJU8HJs80hWWe3gn0/X0uB6BlPqgQLFheL1daXRCMsM
C7DgobANrfil97EEJ/mclQck02V/3SHsMkmWac+fR6pQl9A0q1HeJOubBTlQBHLO
/LsVwtAiQzWZ3y9gQYuvV4JbiORl3dlc8QQX8ei+waH453Xzo1IQMptnaNF4E9CZ
zw8qiP3JTSlaUvSBIlf0ac0mhEFgGIp3Rh8sOiBpRKNFLaqRb39T7hAy/wDGinG1
LFBZv1iWRfOEUiR3NwmYasgpQY/dwuQiWlDNLx+xuzzpMUDuR/vxTnYP1u/UrGLG
mMFnBD+QVDi+exx/uKOOPi2TgxHE5+52B9vlmdAQjEUuLNbLGgj68Z1php9074ho
8eXikTMfDbf4eJujGwn5pOfuwQEQWJDDLfwEH2qbz5BC/Vya/Yg8wykzx/1kPqmj
qcIsgNRXD/HfiI5SKsLpPa4A3780UxTvgHKVLudKsQ7rCe1u1wT+LgL5ZIpBnETM
cjcRdEDXz+ze8ItWgk/QjkUHoTJl3+T9oxyAP2cqsZFGJ7xLbmgfJXgSqJ+5LGyd
qXSPONbhiQI0us8bf1cZpfvrOOkynZhhw03AkOHUtMYXGB4M0C5VK7r72aS+73P6
uzoJC6oH0uohhesNb2y/xZSqTJ5gSkNBL2UEF6JA5zVQWBdT3JfVSKq6Vx4suYCN
xq3DLpvSrRnsIMfOV5bJ3jvs9bXTmgIylrv1/CX9Ogo5JSyIMNhHMT1GX3W0Sh5q
ZI6QS3TV7QdXvfupLrbXpGvhji2+cIXw5ISjEiau9r9yztmulbstcS7s2rg4P1Sw
1DaixSpPbG7pTs+eGyZdEn9+EPVksRF/+9d/wDPVW9/FaRJgMGJ+EjDWGyiB9Wbj
jLraptPaYc7jwvwGAIu3i4zM5bUzKVXBEDcWLuDmqspPegve1RFPKDWSnPLK0+L9
57aozX8f2iTXGQJUzNySR6WEIwDkpEbNSJzy5E4qQn+0DTrsUSFb4yJj9o2Kt2/7
beBty+2eC6oIcqzkIQxK/5yVVniiLAahbhDyP8CekzdGriHgnzzh2cwIUTkvwCuq
NM4gI+YXVx4GqfBB9yIJuh8R1WT412M+6w0Nil06WxFq7F7pbZiPyUb3fCUuOSFg
0M7wMKC2V/A06ez8j7pBUaeTDHNIYDfdIE95EU3yCJRWhyubspIzcHiSKOhkkqAe
6IZoGg1/b6UjXoOVqvktGKqKVs0rqgpQRg5M96RhozKBjPCa/YEKE+WeHTdtbkiw
DamjnfGJMWRh4xYcy2kn/ILDpu7M7HeByu/LnLgkwhqaMCxLA9DS0+5P2TXTpgit
bY+Cx63d+QOlYxE185NTzWAYksEBLc1pLh39x9fupeMyENc48c1oHU/B7i1xoUzP
wenjiuGE8+3tKAEj68ASYuPBbXkcdbd9Ag7TVmMRafm42eCthOPSCh/c6qjy8v0m
uAUp3Fi4KI1KTLG0FVlyzirZ1AY8IFq3pM2ScfFSUIhMWEJzMVGDsOJMMzgmYzP1
5Ra+YOCpBQLIMoTFWG2uXds2SbZfTf6rDxPcnVkUI0/T4oqcZCyKuS77KxNMii21
b4433ksAhuQwcLkBdD0kViazMmODi/j2utsrely8H2yhjLP3+48jS4qwYW/ZBZWD
JGpsOlWR30p9VQmXU9xbB4nSIGv3Lwe6ymoy/SomhG7IMa29MbzxmxtqB/AMucVF
//6TrV3OyxR+G9aZ3Jfb/MTMUSUz/hxKTKao4wI1jYUeWswGf7n1TyLNptkD3ug6
o0nrt8Ys2CyaAuIp0Ltv0/3mHUf3TK6pcUtVl3pmngP8UWSkXZGhaFvbx39MUyDu
1UjyvrDDNFJuXBZrRgO2wgtpCkK1FVC0yoW0y2TniCaO4FaUncF82UOdcZL66b10
z9yDEGPEA6OGiYqNiNdk4NuEFzhn+NfBaDClUOXIwn/gVeqx5H8qi+omRSnQ9I0F
zX94bIrzZXK02j8hyUHqpdD51lIEv8oTysZ9K5AiPuLzOcL41T5TpHZurg4ppRH3
bZ0uUDpve6kfHAnYWSc3sxTpRTahopYtzMntsRs8FA70ngHehLkrVD1qxuBP5uyl
yKeOBdtuABuLvywEinwtYueJ1W3ARJdENpjLuRQb90YUxZTES1ACMg3vp5q94Tk5
0uFW+roMx1cXnbJe3wKEQsgg2Hs7pdcdZ4LHaLglAxYMbYwG8rZxQhfsfJ0YSP70
uwjW6PntSMmBP5AvlAnE1LRioK8/H35dQdYr68PbR5jKy1qrMRWGVFRRRLuxrsTC
7++rkyzGGbzePqg4kWNTQiPP0h/Gd8Fy26inc8El4uPxAlA/4/2L2kdV1NUowz5W
+dUBxka9ZDqgrkKqpcX+f4X2TZkjocX9NF5JInz+1s8XLho39uLCNJhqncBeQkao
ESSKG2DPbMgzk8gmukxwGHldZBYQelNTLS9e7RfAWRETXWZkWQ50lIXBf0snkWja
eCsadFqPp2eRQMzS6ZFRkPxHSZ7bHqoqZuBdp/ISdN5ml8KJ4LQapp12SPzWbfk0
7QuTRxUjIeiXi5MdGK07XhaFZlllEUJnxleuISkmEDlUV25z7k5FH+KeLvzkPFpO
K0ImPlomvk8AnFAEyGtJQlLuxXB6ac69QA7yfpaMElnQ9jQ+Zlx8NsGjOfg2oImo
Fq6rgwvjiYuadxGSmuURKrn/kO632X9ZUKPkCXygSOCBgBHaM0L4W8pBOEzlXEgD
2hrcVOLOF2JjRbT6GnU+aI6rMbTT5ioerGCLV7jDWZXUwPGG2B1tLeKCmazryeN/
wVpuQspX8hN7YwPElXdMvuGY8ZJwpYjk/59tXYtkPCxPsYC1uf1kJxUfeZmlBbRn
H1Bi18qXO1mE/wyIzZmnpmOj1+p8D4ZOlrlJokCfIm4F4+6A26pb7SEXDVjj9Qfw
2B4IGtGntN0dZBvckfFbnMHjq7ChzqVVf+Yy/8Gxrwvee8/NHFhuFPM614QSM68h
jUi9gRx9Ira3UwdqDHPe7Cu+YCpLL5odlB5Rq/V0xAjHjbzVsQMGmdoIfhW5xM50
UM57UCWd6vL3FoGjIkBYZbZvx9xalFOGsgUtO3tvQcnvmvqjUrYpZ8l8+x+acEAS
yW4WQ31GgGifoh7wbLtA52/43z6ixiLz1yg7YRnX8opfDmEqg33yQpiSShTp3R+K
8gyzOL81WQ1HIsMSOIgGTG4aqQS7A7gNQVzvA8PckAM69DBl2hqiwIwVwu7QAAQC
OeI57lBe6MDLU6cQN8V3K9mVbW5X6HgG0nP8jImD/qKxGAPYUTu67E6m8z332eit
JYo6FgGJ5Gz+D2MMOQOtMAV3hhpE3VWJfQUsmy+Ke7F5jiKPlhpZLZjvRbFGtPCw
BRN74cxguJKjrnm70OxtKIyug1WlU//C3GOFR/ehwFZHGrVnSO1LDTp7FdkeyNu7
iW+ymwOcqKxCYRV15TWzZuMICK8Q1RcNZuJQI+TEnuZ9/X8SvVKsmtdeCqU8t0S0
QIAbXrQma0f3ouczGcjpvtHWV9+tuWaT5gbc1x6OMxaBoh2drav2sULIWvlQAJl3
q7uF/0neqYDhYayM5zimF+Oj9dgwkM4SyJ0lz6NtVZaPjwT2XlWShmg+bYw4iiEg
Wx3GoW+ZmlYnWRe26Icd+KFayv8GLKtP5WePQRUGKKJ/DnZECi9NXlQuiWCCI+ui
CIe+X4NEOEgdW9RwY96vhW1Ui9rCwUrl4B+DnCggYLUVf6DNB3tXDMqPLDyyxdfj
ETogvfUA/N9Q8dVw9QvcCOGg0VYMt7VrVR47KK4zRUufFxWY+ek7yISHh6HltlSz
8gfRwW8MKj8mdX11XPYuBBEwHgdUJ4qBNFFK5eUpl3FuD2I0OeThg7EszcL9YQud
rxQzLg+YgFwgLGlUXOyBIDj3jsnYXZqeH/6OKAPUC2gss6Ni7sIhspM3+uM9aHar
LgabbL3abzKjW796mQlgWGeTtV/m5aubOwoMk5oqfn8oHx9qVqf4eY6nAj7uGfgW
LITEjEAIqwpca9MSkbsJQAL0jDUOTJ5crNBiGukLqKwwb83U/W8DU4VGl0YLDi7T
VvyDlhkZs8DNHkliQ3ZxQjxXzzb1Nkhvs9/tNUNTbWYgYItblCdUAiK3KtVG2HEO
lWfletlhGJLt2p4qFxEnRAUlDQvZlRV58ZSPEinjCn3Q5qFJp+WKGzr94Cbqb9IQ
70OV5Q8RNrr84KcQsx7rqlKFcCX5S5AMk5+gKdJGAdOZTqry2ZLHvvECJDrFkWbn
70TdBLmf2/vUeZuwJuemrEVcbPr2TVfkSKCtplgIOL6Y08U1XeONR6NlsUz7XUr2
5bM4nxOEw2bEEfyWLxiWhhZP4U5AcwQbDzp4r+S1fcH+frCganlNBUmxC1TYyPB9
yYj8iuzTPqiqitO+N5erZJkL39Mun9Aip8zBhARtk/P3lZMavcBLOej7vGYCBw01
FQQWvo8MAgAGbXIKpwybqd6G5kXRb+ygu2vgOIncRWTKi3gthq9zaVebEGlRn+7q
6V9F4ESaxkXGaPERX5z1w3eUX0UkJTAm8nTmthPRut3nMEEZ3kCxEsYkPvL7wMab
XMJLNP2EVq5Bbg98r8o8dhM1aqoIvNEkvQpQ/4Wyu32p1M8Wp4kNuDgI4WKes4eD
m0PiUlz8g0OIlFqm1K2fCn0aH7s6eyugZ9XGrTDUr+Tky2ZwZVBT8VtIeyUrBIA7
s8PX3Qq2g1NqgeMafO99xo5rOP96cO8ujxzobhR4uuVB3nXWsbVa9FcEkuE8C/FM
ZMHiNpQqiLZeOd3yo+WOhehEd1Oceaj6UFF/r7Zumo+uXh4RChdxFpg8fG5DFyiE
rCx4/9TEiST2slaxsU1mk3hmFOGENlceg2DAV3CI4w/vju3WYYFt2ykGp7kIIO2e
d8tp3w/+5SRBcRPIwtTHaxdHDfze2nTF9tcbX1KBalryFPo8doukuOfyPE2+CTku
GOVQTdi6I0q8dtIvx83Lb42EWBIMWasGcn0MNHMJBYULLmzpuo2efcmULMZG3uWp
Nl9gLiMUPQQSkbsc6dc7S5VmCjGpX2kFhYcnU1i2QI5sj71rwfYVWYzyOd/9KIfK
H+YdGMJcLqFQimk60bLnHsk3jNU/W6DUI5pv/ooBUFvIjAnr4pFZXZouw489crmg
Mi94UNnIW10a00sjIQXSsWFBLKJQ2Sbp+tnae+F1ONfpEr50e5k9E/qKqUwvx0xV
BGUyas2ztLUilt5IINdw+9RusSyRwpdA/w8FFZ2xOd+r2s4CQ2tZjKnaFrOW+Fgd
s7eLlYHYU2zM26olXjGjrYwKF1VKtmjq4KUwLuim2BzUqorKMb4eEErIscYO/WOs
pXrg62MotQQvlKQhUGPo5nIZcnHzWhwDQxF58evsjcEbhHP5hkqZjl4UlYxBu0fT
pHKqCk0xX9v7YIJyTWzk5L5Gsv2Qgt0Ho1+ZytGbiq1QaVFNBYPMzm6sPvCLglQ3
qj/gnsvlOjoruleF65M5I9GRiq/AMey9ZHRLteumzhW5fXjdYhYYqE8+w0iI0xcd
B/e4Obot447d2D88UdcAzXWf5n33Panc9yF1ybJzqNUpZWD+iuvKE6LCpBiU4Prc
pZhm2oMaTpw4id22gNIUZKMLDzh6nkvkav41YeoPX/VTWfKwv/OJe++zdjsW1jju
Q+ffApcT25zr1H4A+qmv39jmmi7EG5Ayuw+g0OtBu+bXzBXyDypoPKWWG+KWsu12
Vu4iToHNgMAEBHUBo5RB/XruqBMYGgV+LYLYZR1JpUtsR3TFgeM3CZKLoLKeLRZa
d9v9mpP6dgup6sFPb4Q+M3ViMBNQmvO+TuSnsL3v6zYia/h4rB5qF8I9j7OJChFV
z0aZ4QxXRNwD1rQHpwdobG0EiQ1npSi76SqXDQzBX5oF8VXHqfJxV9vFyUisw3jn
dK86C2TFtJu/3nJXXg/zK0ARWJ/5gg1zVbG/GU8Lhv+naxhRZMnS81BNGHIe0HWb
9Kwka1dg6lMpFUm80i8X8UzfBktG8m7t81e0gFXz3ZYsuAz3+XLNgwgmZnZ2uaso
VpMH5M1LC78QFFtgTRw2DRGTV+Esb87MMdn5KaJsWIAuI33mU2E7XWJ3b1h5nUJv
4YGgn2lRaFQqhb0RTwK7vvr+GFsTuRcuxCGq2L5qKe77KJ+7bQZxJGqzUIJJUkHL
P0LB9LP0R5+4Bk6KLuZe/ncbKEf429uAyfJJS2/ED4+Hwweo36VHA74GvM5ANlrU
jDwQKUpiSdtEjIyCL00Y5ubg0fqtz9F0ZfhLNmstKQDb+U4t+/JUsYeI4gAdduQ3
JVNT4OHbA3ukgFfaWc3uDVefQkyoDNpotmUwv6QCsx2YxYWh33niFbuLVLHWAViC
bpXPuFPPmtoGUdQtLRJWtYJ6cA4IWZf4yoErsdbJcSzX3/vfCjklzNDgJIR5rrKk
h0Ih7KiJ3/s+Jbyk/cVOtdXipR4mZau/+y/m3q/pykvW7EF0yhBzlH12ZClyCLd5
+jnRpqu6waWMGJMhty3sCJz9ZbybmGhELmuqhwguwgTJDjM61BSqBnCNELFKE1eo
XiA9cV3QXCFi4JHK0KCDwcC9lnt3NoZZ/i9zWZDkSzq4UWJW2XZKwA4KZa902Cqe
qD8FfRTRBYTeQnZWfGt+7ZXrlQAKQWR926BPwlNU79BNCNN6Ka7XGgtcrVrmRgkU
ZxeB4e/QMTVd3mmqBK4QaQp3pmWchLNBc6hvC9fDhCDIdYc2o2D+jR8b8+nDUnMQ
ja0RYq/EH6VwTikempHzM03U4UfmzPb0D8tMGgI61qE+rJQCINAtiXVlk3NS6V5w
AkQ+SGEVkRXn+W0bbpVvTDYdt118eNToJbO/rUG7seIe1lnkzl3A8cLGRFUtR5q/
kwFbI9Ra8vxq0NYcMs4E6tkwWd9ypD8tuLH2gRoIqynkPEVlySX89kIvO1MwHK45
Vq9g1+b7UATzM7l+hUUQjLRf8UJI2FPGEBlTnMZOwm9UVgaG2L75IsTGkTKHD/Hq
P28rwVEZcjFe9YeEAfPmSRRqdPwQ62CDRgHWWzU59QkG+6sXB/so/uvCBT1KPn6G
C+nixjY29dSzBpEJOF4U6DyNa6amK+2hCdRfs2IBsKt0nVC5/Iowd/VPOfvNEagJ
fPwMOMfsq7He0trWRnwnF3GWcfnOKqZM+zyHyvmI+nFQ2YT+XPzj+bzpGmXnv4CB
0KQR1++gl0gcwcuqc4x7+gZvWHO45eH9AyE8IcvKoQJRZVkzFaIa9XJyVUSwM7Lc
B6v0hu+5nRDz75YNAGYebePuFydN9PUHXDcd3Vg+8voLuPUMzGLkap0jfoyP3WES
KMH2KntEKp0Txje3QuudI/5hFgN0U2gOAh+hZZaAHJ57fqRRp4gbDW/L6Ka5hPiq
99cDLE1oa9jKCxv4kP+pANEwHR24wQ20WGtcgMsbZcm1XqAAoPKuXB36cHmJq2N1
c54YQqYBZzjHCB0nqZtEWja0WdnOAhuLLYXr/G5ikd8jV+P1NV2DnQPNxeEr7CmY
8CBqfftWEooRb7J9sPECTs/TJtEpXyOFtIkolVf2X9YWylB1nR0kN8VO7K/38/Pq
KDzIrBl79kWtOn9+HnEtHjHQLTHtmi62HtdX5pni3fXnui8OGLZT1KtdHu+bE8Ni
tL5beyEk4JvYkwXxnnX/V/1odBUGJ5c3NevxDqwA4sjh3XzTvlAlDpXB39NiUT8X
YVOhJcTUq4JVdWleHU79pceDcy1fQKV8sn77+YHR5sd8l2NOtFLezT7Wno9TwCgo
JhI6PoA9BWpAi3Ctl1tcXo0JQSttY5p6eWfdm4sZSYuufZiOxFBiJ9TlRhIleMF2
PMtcwetWgHNSXa9g/SMyO/iCrbJpFQo0vyFmoBajxowlQeK1epUKDnBBX39xSh17
lgBmw+ldmfX04mC+NxYelYCqGI6irP1pM0yWmrCKrAG7GB4KKSl6WFOTAmgf4EwU
Sc8TbDzyrTQ6X5wx4xc3gT9h17sbL94vmP1GMdEKZSV0AeU3EwXQP/ObDJU0ByRS
6ntB+/NEr3t1U6mtJV4HlRWvlW8dsIwgfBq+p3IyT12n5NN36C3qiMXFqZtWHoE9
YJl9lY43bs3df0h7pcN6g9ati9hAG3CKplAhjxdHP/mTgIPDRWw85c8rvw44eocP
TSWfPHr8a1OBAYqt66iFFxe1TEX2Cpik92dVlI4VZqKlp7+0suzA3IcC+WitREXZ
UqqIVAyiwGezSS2WmTHKqJUJFLx1aVwLTrzJRz5NS9/MA9f3x7//flv0w69lXWXI
sVfuYm3mz/gaNH07kkJoDnSN5VHsLlFMZ6y1fRffJkBif5n+MhabIyzkFEHACHpp
3Y6qBZqJ1/wxLMGAwXCY98UHCfS02jURvIa64mXb0BmTozev0WjOj4h1Zy/bI+0y
y1fjF+MvvVm46qvwckn/5GjWeGrit1kJGQHfF5Xzj/mpl0tKBAMnyYjxGbSbo0+9
RwP/ziPkOb2v39OOPLNZbvphXor9NR9F+P7/kgl49klfs+sy4bCQGYF4ckY+K0Kp
/OmNqaZD9smc+bEJe/WddXXMvzGpBcS7YeVC0nHpTJvsxRyK/xaYvJiriKLwei9P
4MX9Lx1f8F6FbiiKdh5IRm58IEx/VP/Ud81VrcD3bNBcSfJ/pNc7UpKYSyBuuyaP
0Ct8vBdAEeV7c3oZp6WYQK0t6WUAL87cOMeUjU0DWz4uEUvh6EfalX4GBa7a17/L
0cBuKdJ7R5GyA9d71/cWH6W84fJ31K7zTiubN01F1izI5OP1G3sVyBgRyAOc7ymJ
ftBCsjuSkR0GeybixXMb0elg9RKM+WN0c29wGNDTzmg42EmPlHw1ZEDeZ0x3/IhB
Wi/RyOKC1voehq1Mfh2vG2iycMRwwLGIzySPmaYzTLjsOVVpICahqdJJLCOHeWs/
DAFy2009qXrDUs8cihEe/Mrlld1CT9unVbGNrFDdYCLE5WIg5J3+PCB7IP64rRb8
1ZJWVcTPh8vQtmbG4jEvY8EGGA5k/+SbmX4qN4kKhpeCJKLPKlvLFFb3RPbPhSVd
xbaAXDkX3RC3WT2RJ5kGS9AOkeRS4MHgiDG9QnueUP1ay/TT6RdofDIinwWTCm8w
eJbTWhW7jOFJBLJHa+diD49L4UqnKTa/l87JqwdhfM61LLN5AG75aa4AmBHt2OLU
ES6wHNDKs5G+xvZlAWMXK7FBwF0WphkcNqgcDE1vQ/2/kRXGiUecL21N21Lc9NSK
JIPXOQXz+wbmpXh9mVbRYMBkVkIXAZ7CNhZ6QXwHOL9rdBMs6KIEqsrKHtE3l8xq
8BbRf64bGQRj3yuGHB4ROE1BUXHZypVgvNaZjebSrBInanedgdu4WajSPzVi4kNY
N6pv5E0R2t7nRAaYrUJytaUoPHY+Tl7y2mfwIa+4sj47mQwZkJGqtr7J+UWCJ6/U
6ysTjkIHp+MfOIiV7+wOgjUBFMA2AsvZFyBwWbZd56/Bv/LVYO9vlSJS662gc/5m
jwjeVIikFbpNINdlEGIn5RX1nspLwevlUrPDpPTgBKi+q+Hy+B5aYRzER8+bDR+I
C6jRwEy9l15LRetbVbLiNSdwSuhwFxpMw8WO0bdEvzVjRHLs2pfP8omfX27ql50V
NYbEywSOqmSlT8vVzJu87MGw2cN583dNKfs1yzh1JX2SG1d7SBcMS1a6HM1ffViE
1aReC4+L/g5H71Img0Wjf13MXuSm/kAPGEBPHPPs+V1AyFmQ78UzS38Nyr2EdVZF
GEKfOxJujjdM0ypfVEB56M52r3ZYdilYNDnBi34z+1AhNxgtVtnsoErGVDiMcatg
Xmn25RaQzR2liKe3T+iTETXZw6knMHNsAM2VJe91NesMWMbGUj3sAp1rM2vPWY+z
Z+PQ17J/+I7OrJWL7PsqC0cJjDaLKWbTMNC57kUvJvwBSKbpa8rI9LSUOC+MRZqi
0slZju9ySBuCe1aA0Auw7UrRhprTQN+HX2PpkVt7I6UwW1+aHaQQcJ0XiTr9f1AC
EuAGH2Mj3rIS3xn8t+LVAcRIDgbSe1ukHX0yReDKvYNGSmnQsDhkZEfQimSc4HKt
PxKSg/0XTXxH8nyyMHUodOcgqX8nPEXDWz0+umRi7FSyjfhHf9I6ijWOG0mGFTS2
sYR27Btvmdj+QE01nzh+F9qGRebtM9UaxWaM76Pa0oB34YXfioUme5RZUCPp/OBh
tYFM26vKX46IcaPoOw4A8LRt4Hpc3ftwmVpIq1kKTRHoZf4nJRho2y8n3PlQd4TV
BTxK4qfuE13nK0ExrkMFPsGIIs25ccIKA7YulD4EZ+8YEzsCRqmkGAUUjad2+REZ
t8DEMfq/SPp0NKrBNMfC8ryO5bSifG3P1AyL9ovgXm+AZztHsa8rYlLsYajleW7c
arfkqmYpilf82SfirsTb1501l8DeFr2gD155VaV0lP3ZT1U+2rPlgvNjKFeNNUMo
HuGxUKAowVjCIyU6cZ3g/CFueYL6Q/PT4i/UxvYf5GB18TtGIipLwLPmkxsJi1ZD
+Qn3I6Bb2Kz3onu/lEm0QvxbS+Mu9ao6Pgv+MkEFJ+Nld4BGiNvGBZa1fvDdgteV
rDOq6/5pZGEFNskMfeLn9r1+BmTwQXJsF7YKGicMkRhdRfgd5H2nJ0ahHac73WDu
0KDFc+pGP7IKsJqd3z0hmlQGd+lZVdMm4ZdxMv9iEMtzdYBKsda81MeEG3bZoN/6
mELQm2tYker/aNQIw3MyhuoEaRToKrrqdRX05RSkkucYIvWzM5Aj3MlYjlWY9bTu
3XVzJmtFn8IYSo/AAkBbSmlAOkHFhw6+XWeY29QWrVvQ7fzffWS07aHqyA8SapBt
cmDbJcUkM1Y63obLC2h6oi3g9TK2eELcIGbq2dNvY/RU+otzVlLVeJ3I1FsW32pf
32hnT9AjHXko17TyCfpUdBcWiDKNi0ddGkf/wZ2HhJm22amBF/eywSbN83/z7J2R
SW8K5OFwDNF3sjY/pF8s/AXHPAamUEn7edaicIMmaCayO1cJwLr0fw+e8vPY/T3Q
hOuC3HdFfr8SI3S4urZdtqSXaRC6zBqfbvMcegDizp62xiYbjeziZaL7cNZJMbJr
YT7ywspj3ejdoL1GfnkTGD7aAWwGF8MhgYIDv7bCUpKNtNJhn2TGATGzTSE4lTcw
za73OaPq/TgYkkMuMiNr0JPQPbAqPkhCEy375Jh7n5j5JnsT4S7+uDZGjAIYxwDw
vUuS73FPF0BFE/4eEYhmMLjxFtYEHr9zrgT9GFQuBbp2fF5U2wACnI0dazHspz0d
ZuHh41MyTUfHKuUHMJJCJJpVqhyhduu91hQeTkpk5hWrBPl9ZQjgE8kGa7RIBdU5
awMHc3JaTuwYyjW0pvElv7IWMNgHgWqEM0aAuSJMcfLYlShEH/EnwKdLczSG+hu7
LlvGotFcLXaNC+yXnqfunbP43K2BJY4YbanAsFFBEi9qg87JXqT7lOVr4AoHH12m
in83RZB89WUPHdeASNKB6qZm7LJqvhDv2eqDQBl2LQvVeEYadJvaEv2OCi0bE+5+
j/vX940SWXr4+qYCPSb0JZ9dnkePQfFDJlLhO/YypdryRfJpeLnQia9DOM/M8xmZ
kHKq2KKakkUXwHmFwVHJ6HcpQU764D4FA83bqPLYJa8H9E79BbeHbdls1l3bVTKa
OrY1gmPouZxSex8zQ0QW6V4PJlJKEbKqv1N5UbkBxcwhAPrEN8wjGKSPfexhCTuw
+FIEh8r8YiMCf16drhfBzebWLAAqzUbqGk4RFMHgv6CQvebbp8SJKgr7XSiYePhz
2Av+bvNlhhecBQ6WxU77vE2R5uMnCOmnyeSFSuWJAXY7o+bnOgZJoQfTSoq4kYKq
06+jYVxgrCEBTSQEdKS0UZ1RiqF5fdpRdvdkNAzBkCwt6F6wOm+mtx9JP5FAtjXt
cdQXTfidV8hTcesS4qYk15xj90FBvuTztPjUNYkNnPx+Gy/Mi3Ls3/1AycHzrt41
u4dVOxX8VRzFHSTHx/dL3/mTlSog4u2aUqg7Xe7wyLF7sBn2EWhhOz7EnBxeviIn
O/7qf6nfLPPG1rUC0MrlrAePeffNrL3Dk5aYEQObhE6mB1KFXFKUuUyCP8qL5XVi
MeCU2O6S6w1zG6FTg9kHgTpFriPDTA7fJtZn5pVM2/MG0S5DScPh9dd3KNF/kA2c
IE7pSvPnXghxdh+x3+uzaJGii7cjKjPzHfyTyYx55Ns5TLN+acvVl9YCSal8yzZm
vKcQ8PZEf6gSw2GSt3fyY0lr6Womp5f7+PgqNoTv0tdwWSH/uy6ujwe4GKeFhNWz
KTqxttVjny/7IqZLbWWbhKNzndRSXCtn9A4sbhD3GB/PLIknlxq91lwiUF/GQ3sJ
C98k19FacHVIhMJnHrRhJ3jPQ8iiccNzLXF3Yh1r1FG3dMx8iQ+8DDFuOej6Djqs
j9qczVMZt1uJlFtDyYwHFtb29WlW9bd6DJ7jf582k35RLbr52LhOl2gWRM3y/S4i
6F+dWRaStuTE8iCKPSDqBJj0Gu7hhMIO3oNapru4SH/GoIb33c6n4oaUiAD2qv+R
JU8KxN10n7buz/EdG9VW20U7Yk59gBjCOSiHXWeOeX8EpRuA7HVsQY2EHh5yeMgv
CveP/6QVzE4k4UI3MAwgTbar3tUvsMRin14wqBLA5YVzXpz7PKCfApEOWcXr3com
XjFyzy/VAKcxHEuWVTk1xetO9xeU15uANymjFrhqT7c575tV6/Zrvzn6YAHkEnJy
Um+qGGsx+iWz+KZzPYhQ6h9j+MZzK9/jiCK6aOJPYpxhnX4Nztw/pRfYAJJoIpCg
ARnXVVIEgOR5ta4XRyxvnha0O3001Kujibv8T2NvenIbQinEuxe1jiODxoGpOQRX
vscHddJnEve1rBEcCJkMqkdjKO85UbkgjVs4j78d4feIO5vY0KqBiDSpRFgaz4ML
SoSBb5QZc/a9V1sCmYBlumvcOXpNFd+xrqc+ZlVLwH2t1rIwJU8jUQpBZyW/QH5u
TIKUp9AjVIO1RoQTq6YFF89SozB62KSND54DY98C91FAHwF9ftmYayHl2G36dUui
m1tdKQ9+1nYERrBV49aOYbxiakyrLq7cjX0v6orNMB+MPe3h3gqfPGJ73dN43+0B
ZnnYpQflhZdKuuqENnHQN+Oz774Rs5lWDsIvOisZHjuA4rnJgkTm3RlFUoipVp/w
SDaq3Su+Jq4HLnzo5NdwA6C8vzbNSRW6DX2Lxx5Wj7c2UrbpV0CHMrK4Q2Gqpg7P
6HRgXcOwkmFLC9eXSLTKWvKwmV5v15dyLJ4r8KFAJeqRReFFz4QYYGcLIpBZQXDO
p9lIBGfzPcJfzZ6yA3PX2R9Xl498qsae1VtHzU7+2O+6V/NxDuTyAl7MV6b/qmnh
R8fo68H91uLLY5LNft/aUUbFF7R26n9IjB2ay6tFFlSEcv4z7FGJdZWKzM37Ts9p
PM4p13vf8Fzs7YH0WZCLBzLaIibj3AS+i1k00L3FKFP5QC0ihoEZ+kzI/DtdVcY+
OefoIz9+Xvk7mOHQ8EqlOeHsbfPZGNQMYuNcgACI6BqaEK0r5Tlk9hfx1jMSrJpb
PZfO+HTfjx3HLV3rmpI989zAmw6yep/UMuI8pgQRpZGou4CnOmhK5TeB9lAkDk8u
/OfVpLW0M+EDztheL7BfL4SBq3xzQoeBSh4N2TpzoKyc0h0OUEQBqK2g2bnytLWM
6q+TmHRpk1jN2eXax1ejbHsRj1WTrY6sKkHqCAXQNP5KblU9jHXnVOB2v6sdXycH
IssNkZf02ZHEBhX14Q6GkvlJVrQkDIyUSEQaOXHKZwBKv8XTaz0aW9kEeHA+qw+U
2W+f65zYcnc+s0GgmNnWCNymJ28SmGwOIWEF4R/uPvgAYc/aX4ynGiCaS3QrmEXT
PSKP/ag8rdFORn+FYWUZtZyECOWZASV3aW0QQ/ZWTODhg2qvvBsoDln/yvrOWfdi
Az9F9/nxByBTDgSigErdMW94w3q2zxbbJrfeGeRJb5Hz9gQ6vdPJiJ78p5YnRAdT
V9K12FEX2KKS3f6Ewvm4atak0rUCDdR07q470/TlWzcFOsWC96aLugfLPrC5acRo
YjQRhYNiu2mKRqGpfl3h2ZgbY2hqrypd2PtezUONTGRPElLVCqd8JBPx831vhojg
LJAp498vREvGx+M9DQXy9EUKCH32TaMNahT0phedgx1xz7smNw4N7RBKTFq+11GE
4Q3pl83blhFiQqPmhbFXqAK+5hXcvqxt8fb9tCCgkU9dwjcMDBhU5TnSK8Olqrgb
MqXXEJipeTK49LDxzNqH6NlkERVNssEBHoNu4rW2MjDAulAsKn3WWYhjLvbigENg
NJiV1wcoqYehReoVRrYJVKMnbPiG3CfVnFMj6/VAXzAL/jf3SEVx+m8iNHj3aQw4
BTyQsH7AhOhIwOEAKvVmYx5nV74R4dqAmUMx44rY1aft9TtLROpJgz5ntCHbHoQZ
xamRKMBRMmz5MWU681ajIIeLQhU7voe92rTLMoYNmf07SMpVNEDmwVtxPL/+vD1U
BRN75FPL2XTQFVn+Y4Z8SpavtXoJ1ggegnn08jEyYgp23Gsr7dpgARb79gxXic+g
Ryw6XYFD62s7mYM2Zq7eMsTYlKcTEvFCESuFMLTEumPkCInhjQMRNTMhdBZsx8R9
cZ4izXeY1V6ADinWVHbUCYtaNXDh1VB9skcJPh0g8EvEHKSYT8VLZmB98IPCCzT/
ixCsCInHSQDkiHyCe7K4jhwFKdb9m0xwm+IDWpaJWDD0knlaWhRvXsDDOI+72+LO
ZX1LP9kfhEovBtikXHh888NdqOQ9DR7iJIvWW/eipJv/XTm2yi/FxrvBBhvDTdCv
LMACa7Pz3z9h8xRgEE89IGliGDcHk9hHwKk2lTwMus8dgaw4Fo2x6EdC+kwnCOgQ
MuXL85H9ra3LvLYIrC8oqGk3Adc1ESTIpDaXmF+m6u91KMjWJ6ci4alr3JbL9bid
y/+QWnk5iKduZRP2Q2y73c3FDzR+VEUu7hoJG7XYu18y0blfT7OvFf+dvk5t/bPa
UHPjOi8f3o8LtdYanT+wZheFBt6UwuuiMs9O8jQROLAMl45WXUmNMSNY1OQDWs2v
Vf6jr3530TB5QOYbUR+4wey1etxa5l7Yz1rRdyJt6SlrjVP6Bb4xmBpEBGvVIOTN
U8Ro6SqTytxtCyFnhuhmESXFjyGwMfiaJ3GSLcO2PboLpXdOoZztk1HW5AfZbViz
kFqZ6Qi915ue1AGn6ajJLTQFLpo+GRluKKjUKF70RE9UqFlkBY7BP6j2zoYiz+kY
w/jgz6VwJqbvtbL7x4Y8IFHlB9rg1JNKlDLI3Epo97T8JCqIk5xawvcZY+b72r3z
e58yKOSvgPuPF5apULyahoCdAQtXFA963bgUASuJvtqkxsLYWWadfpDizqvUdfhg
DrvEum/OKbEbFlIwFwOBKjyWYbHf2VH+5BsPpJY/G6Tt2E5RjoiVxPfSAxV6mmm4
xd4JEjXazcR2bamxBl+OTFFLBdRYjFt3g+I4dalMVPEz8G7loDEbPdH9WiHIDExr
B+nHM5I61vo7Q6jNBQozIEdgfM3KJY7nb6Pw6aO/M9TO/rAGjX9ZHk7SOGK7rzNB
a6aOGC5iYOZGPOO9i0C5+TVM9brbLJhsgzKszxe6HSn+Kc/ykpH56t2jtZGrBskv
cY9kfnMDmxPvQai8rOPYEKqbR0Vz1Z6h9N4m6z0L21OBztXt+X9OlcvQfJjO23e6
hhtpyIDmfxkJt44kWGMZbO8tdywhS1yQj2vAByGAdaunj5MfkEiWnbTBlTuRhsfC
zjCFWXblQbWXgOpxdJ4zQasLTxCvc8ylHE9QT7QQHI3rbGwbbHKgFt67gD/AqlNM
44L65ABX+Mz+Qd8iEHN3ezwUislWpCNgHsdSf9Qa4e2kMTIi2PGwwQJY1Xz6b9IB
3ahOgd3WPwLluoEkpw5/ps0c49KnLISX1WQO72Z4Fw2IuFtKA0xWzEsCkqgKrXF6
sRXkWQ63RqaN8ftlPgWYqk493IuRXafOIjKb3GS6LdvbYDzrMIkP7oogsoCtI1rg
q6NVfcoX+aXT+IMWQiFLybWCvLLGEL4hqDbvTxlYwuv0oaF1h7jPVDvcJRJhitlj
amdlG3QV0yz2wwQtRPK8qqgPs0cd61RmKW5kR1pFSrP0zCgqNAzoY4ci9tj/iy5V
5BIlUgxzZMc1vShsAv59EeCoL2oY2DTbB06BoyXmYFvAmfAxOmWiNqEYo7vtqxMw
7C5n8n2dECD1as0fFj0q6xmLuF8UJ7CtqcSjUONDvSTY11pFeoiGMrMIYadP5UHl
EPGXYpilNjKO0ankr40RTRBdogrJUCFfNSnBI1bj4tA6YdsheMwh1zfrJousvA8H
v42uiCIM1L2xgLtlSoFBTA5hnTNxCMqtZaNVQfCPlajvfxkC0wS2Lv1jNPogv2tH
nOz827jWDFEhLAaN/rPTQbIuU7ZYcYk6TA01wjVzSxZkyiNpSyW7k1z5DucUfY1D
oVAyBJ+Nv9oUK1f5IJiiqYR5vgWS8qzf3kntG7pOqrTQLfkrkBVPa5x0z0fAOWLN
Rm+fhFqrqjF42+7nUQRLVu1bhxZUyRSuZ5NiW+2ycFogk9cERLi4Z2xKufq1sGIW
LwbPOyV6I3EwQPdhOwWCR5b7yww+vIuriULAmf3C2myf+FR219j/TMXDelvebAWp
YfI3LgKojMEZSA7tuuFc924vkVyYEzMdseKQA2wGJcGcKy+4qqkCE2EpWvEPiUu9
jOi7X6MjXB9pMi4IlPxt3srOkjWpRoqxfEZDJKukeT2Qs68hXIQGeDlYXnvHNm2k
w8Uf1OY2t2+LkZJT/vihMnH5XxwQTRFRxPhnGtChx0H7qHLwgu27vwJ899PtbWBq
dASQhuAHluQ+mKrFaLgBaOIJ97IMmeN29wQdBNsEy2Taco3h/tTaTZakafnsvVZi
HfXhoZlnUB5sOKQ6sW1LqOdF4mV7th2cf899JJGGSA2yjeGuO1FJunasI4INXz5P
/x9WBEZCnnYigZHIAn5Li7XLq4Q3KPTwXeTshHIldQ1xxo4ItpnBjkYOKuR4YLBg
B4xTx1wnehud5d7xU82iRXCARYt4pIwUOEAp31ewGjo1+JjVr4G0hHJxTaNN6/Sz
CH9oy2308/xGf7O0lQylRfH1RYl+74d7Yd5ylvx/u7r4OiqJldww83KjlCRMv/0k
9xgHW4xQQOmuewZcvnPmQSYXWp54CwLP2W0oHKRUv3VKHlKO4I4EGTf+pnVIrfOE
gewY3UviLjY88diTCg6jcLOhVLa44yGdXsQu0ymxLzN6tbPYPsz6mBqhX/pkGsXZ
x7G/EypElBzJJdfErQaMDKoMHjNF78c0NdeWMIcLx7HzzA9LYhq0FII2Lx2iZ2Ao
EQWcfQBm8KOewVWcKuLgTULWbZVjf2r8ENT4B3eurm5cJT7fKgZ03pGskoOvUR3m
wWq1z/ow+o2idyjFTUVukcsTmhfjsHlV09Mg0YTLds8d6FJfn92EFgLjl9m3ESgS
Yyg5cnl7qAX5hBOxgFV0XHNnIw5YmyTcVRU2o5eDyVOOoQeASNIKc2GZGDh0aC3n
gS1bdMaj/zxxD3zJaVqChsANz7CM9rvN6ym+nr22ab999H9i3FDYmoxKsjw38xFx
d8NfcHAi13fQU41asHb+CYDho2MsFccL1ASiNt+1Lh6m5cQV5q0me3Q5gbxPQao7
7XD7eyCS1N1T/GXJKdYegApKP/yi8Ule1UOFQuqOAYd89XUkb4ZuMs31d86v9rVf
B16T1L5jVnDy10MkGdrciDhuP+bW3P6yBP78zZUtlkmaaviUlnn4Dc0BglPCnJ6s
RJr2PgXKkoGBOvLLWkw8xacwUWh8l08gThwwvVxRs/qYv0JwGZfjyoV6EIAIOtW2
ZhtIqg49Z+Xt4y/op77ztdr2V0bp4sc9tAHK3npQRuHZ3mee3h+Np25CXzqJAzwH
d5eRPSc4nw+9/d3gi06IRKhwIUI4eaJgS5w3U2zw4YGKLHGJ4com6A8WP84hF6GZ
8oDkcbd+y46OYPGrXSwGamqCr2M/2FPVNhDygVAGLHr2mtz+AjcitUE1kneJrq3O
HuML1TtU9dAYkjX0fcIr1qt4ffJvJ1lIOMtOdmEmdp4bGnHmCFGLz0jKhLmcUadT
QvfI33couQ1kkCHIjS5iXZxzJYc9V27SRhFFGnbB+fwim/rzyI8B8tq2oaDXJTEN
oSFK2XtBLErRBoWi1W5cAla7k+dhm0Wjnf2BjAAYWuYZlRPfsZAP56Ua+pB0xnud
OJHL9u1v+gXjFJxmk2FTFgII4f+3r3lcLGBgBtKIYEWaPHyhEILR8aEM0Wp/C/9+
Mk798fnIoRqPGV66XwCImPR+7iIflmdsahoMuLaWGNqdPdAc2NWmG/lfys15DRVA
nD5KU1/XNFpIycKJ/jmIQ6xWt78muwahxTKvSb3+rTt57Jh+Sz6Www4n+5eR1ZNg
d4r+cN3B8CE9M0LQN+bGjKYDEthrXi9/30OtrhQ7qFSYvVrixNhCfY0sQDIuMr+2
05AvpsaMnHj/k0zfqbwBUCBJ9b9wvljvUuoaSoVIoW+cqxvqVwyF4N7ql4imBRGB
j62l1oDVGFRX86vbJ23z3SPsodwfrssz+uUak9bCXEHFW52NhPw9+TPQqvRD3L9e
UIfcqzsZnyxQ0QNchwkTzwWsuvp+TSgCSYJiwS72okdXohn/XVM2D7cc7MGDKYU1
0PbmsK97eYSolHCQQnIc3n4F/0s8ozEcAwniAHFyY8IC2pfCihfPxdJRlawu/5QG
n5crUrHzc92hcFwS/GsWuO0W/dbJx4CPweJGqT402WYTMcOhCFVVwcLdMCaM3eiu
sjfaMLu0MH/G9ov6RHMZZMztuaXciNxxBfDFehSQrfETlDbucv0shg9Kv+OVvevu
wuwjnhIDD3yM7Fg/78zbiD4pfnj7sD55cfka3pw9Tk4r8oBr3gqOglfNc5TdjknM
iNGiuSVmMpVaDpsNiPn0BhpPwi0Opk5T6ZSspzHNUyjAEtGRtocgF6tLeZJ1YiOO
CoMIeuYy3She9jbuCx5sCvfA9Eo8MQsrpZSpkhAz7Waenbxjf2wPsMo9dnYL80lD
f0DXc8g0RgSlYEhs4yawnjNEGQRBIYql+Mu4cvYn1aWonehNt46j7em4Q7DgFPPo
KO3aBEI3lJwOPlEgqkjgiMdtzgBvx46Anl9HRO+yVyBSo9Zj13wGjC1sLC8OEGnw
kJDTdTQKPd2M1s3prAK7VWyJfaV2VgwLcTHtED8qU1801igCSre0ZchCQ+y0NX6q
P1i4KvE7PWlQESfxAdDpfXs9Y0Guts0KnEAjoeqc3VA2/j+EykRABeM7dABDgYFe
vo7fyiugIorwHssYKCARHtwmTUz6M9BVIaR+Iy2bsR1riRMFHsif+N2JF+xu7ASq
k95WvrbkFv6yuA3dT3bSxUwKONt3ZSfx27pUhHnEn3JHAxYes5b78WHUcJKUGcbP
TDEzVGL9YFyxeR8OzjnBrbFE75oZR+//1heyZID/TcPdq2ERV445N8aJFd1GCe+7
CxLIiPsOXgFxqp9gF/2RV6Y/axTygQOo/Zhw0FiEwf8DTPq9mJYLF8CRLrEtUPnk
5BjA95jFnk+fCJFCjKDIi7KV6GundGgCUtkUUj27XGXK1P/6hqwR7hiNHE831ilr
UZxWFTNEn3iR3kWolYrAi5Z1Km3y6opfE/1QgbB0X8I7S9ybcUqzTriaoVWl+Km+
uXxjT8SJfoHMwWUK3oz6dSfmIHBRmgF5usNi35lNl4efoDhIk5/wMlwkj7Qo+Urd
ILPXgxRh0kW4pBsKMaf5FmulcZkTHsV9aLZflEtGa9UJvJD9nmzxkPDjqthAAUpu
CNX6AhvZLKOI7tGdvn3RKf2kUc4FdDhrvkD/yd1TZ2UV6Jq4zqCgfTN81kJD/voQ
PfCuHc5JyOlcWJyVtvYx3k/MSIPZinVgecRZDYARutz2MzSxdGNDlIVPwFq64I2X
uezbY0IRmxooI1r712MwZT9cRCKo7pypy2R5wCuGrxg9x78vYoI7NjEG0Ob2OKt0
hHL0fIWhv/JIAhfP4kx5mq21S5B1FOJN068SoVRAy5YnDC7dKuuEgE1DriiCFche
2q/mFISm6UXNDQBaxHkP/u8SsiBUaLAXEuE39B1PdhbYdyOpKFzHcRd8pNE36MDW
f3y5KeG4MbfiHVbo3YklV/itCFVFA7U25YB+tsXogsMcuBW0+hp+bLESKyH22htb
wg3nRDhQIWDVZCTfAKeGgo9LXFIZKLB6WuikjtKHvvgoy2Sr1+4RmXfGMMCQqjkY
F6hOeJ5AQa4n7P6FIWc1SPJ/X1p9u3baF7h5E0BTCwcTCUioRJyrZnG1Jm8aTpLm
MfdSQQYhR04vSyrq1tvfEYE7kTqlVS67I8zODNi6px3pKugEpRh7Ra4a3eldS5bh
oJ8jgfVRG8zcKpjjonF9PEWRPIU8n0DwzvPOrIJAQHRt3oezSN26jV9c10QYD6dV
AxyVxSTHtNhTz/K9jRQOemsjaLRKaBIB47LsHSD9ENSua91djuZeucUNbdTrHs+T
uX1l8B6JdT3vFdaZ9SJ8nPo5BLHCJo57SM+5dKQ8ISsgjeJRQXj6nuZ4PyQxUi25
Tdw5lruFZzd1EdgUMmlu3X0U6zYYtra6iSK6qXOfXf/sFd4O5mSCF7YQaiyOnZLx
LaY0Zt6BsoZzDYtTJ/Tc2y7tyQ0QN5yynXBAiTGKD+QKSfiiuvTQ93gcK50tubN3
tE9MDAXGPi4c9hKIsbOahEvwfu48Od1OFyy6NJGelAWi7SUZw1LnjmM9xCcZu8Xh
vQ9q+dCcmpzFF7KZjszr3445DDFUyhvV+z/h88YzNQ+IarcP7dVM9G3CZLfVS5rM
Tim+hZuOQ11AhNb7oolsCr55RKT50jNSEcGeRWBZ02u82QKuVFYnlrtSVoz44A2f
fH2YmXf6oJiygbbwMdv3kZnEA6Y9E+yzEyFLi+7NxET+sGElz7AuJVFPQjWvbjN8
MIN+OobV5ZbFomnmMoAUS7ufjv6NihFaMpRQ5rmSrHAUXA3S6YLpYm5gt0CLjldP
YIvkpIZqIsC6wIo+J42JISoYAWMd3yZEyR6OAGdCDgO8ne0R34jN4Uc3Q7Ns1OTS
l//aBJqUTmAwBGC5Ik2MPecSYp1m4Kdpx8Mydudcz4/cfHCxH1/oCRfOdDc6xn8s
Er+BlOv3Gojv2fVZL24Jn4lO9ufT1HFeK+RvArApEEbTdhGVgBiuVIugQ5mQ8Tyf
VV9+9Qd5SZM2+UkV+kqWTZClxOtJ9LE/TiV1oJcuvZkNKIaTB72RV/kTccbG1aFS
MhkfkvZCx22SGkmHATBPTqa+g1uHz4G+yySk+M5csAu2MJ2AoFRZ1W7F51nSqa9N
V5UqtsCb2lhSTh9UwpbyhQQ1xqIeXLaRDY5NmDqIr1WZoSTGQ2mezdLVBs8hX28D
fTgPjjngUquNHPttqnL+zl1wlL44+U1YeNzM9qlhESvkD8miq29Wlqpxt8XaGIUz
0GhmGZ4ieYCpy1FmFsNfeavKYcjVN/jYE0AHjzNGhFdBtA7h8q+9gSWGzmBaK0Fb
xoRxY8Cmb83fQCAZ78POGlINFgxv5lXFoArREqAih72erYsfkpIY7tYcicgZydcj
KnW/sEpmE5o94uSL3tTZ6tIjqoQDLHxjfEbtFZ2iNE/rbhYj2hVD5+YN1BGfVGg7
s+B44SY7nj/nJDnbrbRY2Nd5VcbnBriVZE7Yc4DDfl+O94nTSbBgoRyT6nfwTeru
qyUB39zUGOJzeoLWf8AA8AVppJVZ00matt7v7H7/SJJqMMlq1LKHegmdlz4MKgak
kB/wDeuuxLMgHhvvoH5icTPEpW4QRZ1SrsuHHec3HMC7eq63Tz7i9EvviVT42eCJ
SBAhvs6buEKRF2zkl1ZHiWJsxERTXTh2VjZHQZA1yL/YSxhJ/nBHzR7pqMMyQkfe
0WF91s8x17K7UDh4Ee91ONjAWyLBdRdUo6KeG1fkdz7wstd1+/JPX9Ii2g8rF/oe
alteCMz1FsErAfDzfetU+pjZj00cQu36pxTFxKTFW7V8Y4ZtbqeOO0SIXdoOFrMf
h3m/aHLKzJnv7Xx9WiOckxUzXGk+2GESjK55X5NB4rV0CfzDLLrhfus8b1gTVTAD
kNF0Tf06mXbHSNA6Fk7cGknwneFLBnQFXPDS5sV2yN842hOZ1ceKfUF9yXXZinrL
Bt0IWNyxAot/y1T6NZKdmUUk+azBHGs65W8pGVH+1kS8bsXgXiPKLzGbf7GjObM0
vt6fdPG8mQ5LZUOSSUYtFGPH36/f2p1tL7USGG6FkWFNJK3nPqEU1+oZ6xThSuEB
A8U4uUe2KPZMJdx55BPI0upjevexa31bpsR8ixft5LwuRwt7nCm9/+6AC4OvvCSR
1umNKc/uS7ePj3kV6a4blR/vcdvpGqwhSQdtzeZ/MM5raMDBX6IqtojnXf4DtAPD
OQniS9JIy5antyDYm9myCpsiC8F3PMtpX+eSudePBrlZkcVd49MbL9CkUYozDGsr
ROJsxV19OtkIEP8DYYs0hSZPEQCCsyxOvAL17fwEAs6WByGMGwDLlqCoATPOB+Ho
IKqdZ6T1GfyDcsayi13Ee78uJ6iVR+PM+PIgO7D3HaT++kYD2RPdrBChZnkHftRt
lmO/2g6sjQFpdFEjES9XdvYnBR3NO5qOnmpg2W1eBJH14+QDXYTnh+bGrahiTxUu
lh0ZynqWoFBmY1h9GQgC5IcKZPJ2WP55IcClGm8WU/aWXCq7m0brAiCabBBQn3bD
9q3TIMRbglpFYwkEcvPnNu1FzKiGUf4tF+gf8bUPEZB4e15Zx9ZcsTnChOPulDv2
pMmnBImZ0mpSmg5p7tTfbcRh74zot0kVfapsCG9r3EccZRMCJVzaBXntXzVvTSYV
ikuVG5UC+mYA2QP5apc0bbEA1/3hKaAYVa1IwQ76YaU17JRQGE0FHiVf7PvJfw72
DFbwdLk/7eqWStZp9CFW2PauyXo1Dz8uNWF87+5uYaOJ7jfv0oBcGq0g9MQiOvGd
xVu4fxs0rm/0ZV7mPCyMH5D7T8lWTQOQNVRy13fa1CIAqrxwoxGCMeRL6qupV6Kz
3Ntby6k8e2QEHvRLeZBcn7PAYpAExaPUFQ45/9MwcJK+ahi4Y0CAq9i0HGueGRcy
b1+0BXozYxPqm7eyw0X8fbQR3kOyHV0oFKUBm4HgoaiW2FD4pOIh/U9Vr4xJN+u1
k1EM+EgnHfWv7Li2N2ZjqOyoprrZ4VRPwR8G0Y2GMT5LzSKv5yr0XIBj0EGhpefN
PCAgxjnU4zyyrRSjYgfXXF0gBE9pB18x36mNW1fBMQIJBuBeFuHVRTLM3p3YYhde
`pragma protect end_protected
