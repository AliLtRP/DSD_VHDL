// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bJdSkkEDNm5JO+xwJ+0A5VBqdXFGdGIm6efJEHylve9aFefsCrDdGwIGm0v7mm4D
Bc4vGT2vnaMPq0s5UJR9Ql2F+xHsR3wHqdXOUmT42ClAYtnar53LNnk0He+rgHOM
DNWz20ELwwUgzKB6FkOK4rKSAh5eTQmM6DS314i48wQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 33808)
ER2nmuF43a9rV4uTOxE/f6VnpLuyitEt2Znlx1ii8knNu7OD8s0YQWA2fBMva5Y+
fvKYg/OcCjY2ADYLY9Vk93x8a3I65bffAIB2tYJjKryVHPxd/6fyqU4yHiZxM1yk
2B+0+QhbS51XbMLPrXmRzmkL6TEcj3zYDPMJ9tFb0GI2PI7CCw8sCyB+1uF3IFdX
Q/pjt7VAGw6bgbsCSQ5ptyGNO4Z6+0RYzTkZ4n6iPnvOOtyTzUHxe6QuUkIkf1bR
8bfb7yrIkeVZ7tR9ya1fk7mPcON4GHWdlxhR/TRopLejbCnzq7cnF7A29WudaVZt
GxZ3BQl6dlwVlpkjfA8pPLyShp1PyVHTrCIhf3a3HOvb61lk+EomnTHiuvUbXMoU
9S9O78fGJGNyBCqJnOKFjTXZ+4pLNzFMWV8K5zcZVON/1zvh0rlKleSdy9bg661a
lfbKF9IDYL0XG9H08mMYN1CN0OYww/ayzswBFyISEmFyXh3pK5WoSzq3ac7xz8Zq
Asjvkw+Q1B8TkupdYMHeUgqBvnVUBVMM2rlsUOCJw1nIlTZuDadU23J+CqcsdiVo
ksp6fGlgqCo8TjZs/mYznctWTam055A3tVB4HoWHAXkGjp1q3rsEE+iGzNARyr3v
RATIOQr/DGZ05AwrV7XNJYTcx66GirEpRFrr4Mmh45bl+LjbNv2uJtTt/203IAwU
8kAtjbCxg0HjY6wdkmu2x2kJeFA/uWwYLTyguDPE777ixYXdIs4+gA7NpJ+l+rMG
nYeknrp60IbRocLlUSuG9Scm0uokGxgIjcyt54IomvIgC5ac0ZhM/E5OF6Ebit7r
SrHeJVxtr0ycyOlXFFIjineVz9lvdNddBth4LyRpWUw6o/8QoJ9IejEZxkmlnv+O
6AVPCjaw0oxOCEAZOSDWVV9colLAvnKMth87MFOIDYKn6su+Sg4TKeD8WoduwdpA
0bJxm27o641g6qt1TqQ9Xl8oR4q3jWpS4M6SrQXJFzb6e2uttHdosRflZX0TTebv
4K1eFYxcfgL1w0/aL012wtw5KhP3StsW4ReSdcI4Tgs/APk6BhP5kXV7X5Qh1D7b
gZVrWhZjn3AWTzG2KijYMYcjGeNhD5zczzW4yn3ETn0kFNO8uknvAp0AYyUvFR6c
OsxDxEIdT7kqe3YpGYkXF87roagFPKEABp5dOLsu35/m1GNujuECci0ublD+KzYm
UHY1K/M8WiyxkTjH5lY8GJ89VCnKLCwz/Tknh2XNSvkZCJv+IhYc0J0w/NzbJyby
rkpeeqJaeFpscDgamGsdjRwVaVUz5JI9ArCtifmHQ3dZHbpvBg7lIf/j9r+RlVIG
oPA9zCNf/yXAS5+R+w/cd7ft2LD4pU+Ge7d2fd63SHiYj2BlUKaWLUuB89HqLCAe
XgHozw+UaF+E5QJ9l1PctRnDgHi5xfBbZjNUwCZ01fTG7qX5CJsKQaVr1fJ5mLZ8
zpWJheD5v2nJsAYBOIiGu5+HLsffYVHIt4Yll0iho9r/48CKzKj3WdDu7YRq/rBl
uFSF/RKU3NyE4WQjoWqaNd5BL2F75pqHYX5Fu3hvzyS1vy+G+JhKI0hjglT2QNyc
S4zwsHFrtP/HVAvzKYkA/sNMDnUWcybTEoysIcHT+GAOvTnxQprrQKQcF7exSryW
lqbL6jnR/eWgVdH6j9wWg3uIK2n+kpCi+KfgLvd1fDAWa3J5PIW2yl/ebeZ5rbFZ
IKtubXgTvE23OfPJB4wl4wXzm0Wz8JSO1AtxTPBY258vlbgOgxlQlZ/QZENpnm/d
ukmBO6FEd9sZNRRp0HnlzO+LvGUyspooRlzcC0yi2pSNTZvyWnY8U6ScpgrcjUig
LdyoOsnzvxqnA7Q06bBENzbArYFTrl1eEuyhXTUG3QJoT42tiJyoeZYNZiDeh0cY
byGpFXfufeDvsnt9oCRygLnj+FICZPUec2X8182qBmSFAaTmSu2rL5InVoF9qfwm
lqALx4VyieDFIQPNFNWpS0gpgSceQouuZ28XqX9Re+E/zLJH1omc0FCv+p/t2yUR
j3TWQGQpWlaAuZYnLjFRRdqlyRuTfopgkxwXLcjhzeQFMTqUa8ywefTuT2r6DdK1
+APEffRK4wE5fjlI4/d3vp/6IOqCKti6ip4x2ilxrGfPVDXRiKOZgBL09SMb5v6y
nNRnclHSgRT04+vUnB8B9teletcogb2JPxzUxIhWRI4UnyYgkHHeeRWlVuEx6NQ+
smSYh5gi83oleUz2qhJk/VZ+7Fa8fKAJxy6T9JHWrtktS5tU30JNeXG+IVVGa9z4
sFwQtd30xII1h7XLkhS37jZl+cKxBlj4l7cxhoFfnX7YsqH5eWmWLl4HVy5MjWgx
R+eF7BFeDAekB7WxIVDJFaRS4IF1jyd7lT2+TFDytMQoIZGwyWE2RR1CfSgBwBy6
nOVt0thrEKbpd2lvzFAbmkrMUEq6URWjELIlgnrHU3cOYQetw2ALTkZl7lpbKCq/
+tM+d6OwWE6I9p/U+p5/FWLPwGfZlJrm1j1gynHGCDttIM4bbHVPUbRfZycXnBhf
RlDbKba35Xmfnfz0QaPg14fWudwzMt1NyUFueuds4JgG+6kY3nhPLZg9YAoCQa6o
jJWsSVl+iAUvY+2ZowD1BXubVqzPtJhL4EdS4VmvHPGA6dj+rzsulPcjlENNmF61
kZsmEyzga1fj7LGl0dFbTXmmvUF0kbrhTBqQW0F6FAvTILHD/WPuzetJoZVmGgVQ
pVVKkczVvT8cHOlrrV5LW8JmVopPz3sjXnxBt2vhOyTCsJ8LTXRqx9Ebh3GntIHv
dbVSL6B5bsvCev6zFLTRwod4w2ETHXJFOwdGFmc2Jb163Y1a21A3DaEhKMWj6GJ9
TlnzUc773j4/dNYBS3j8Pm/f9MDgPonSoCpKitojwgSsRZsnHyHJS6zU6MW2qSrh
fIMjd97CsRyLRmbYl1LyOmU3BnOtQPF3Nz0VsH/OYd9Pu+kjIrof7+sF1OETKOrV
b+1btOwFR/VMTkvmlmRel6KvIvjMQcD2LKEzb6RHuIU/WIbbeGP6cL4dMysHYtjX
DZVYKtagHld0CKl3nDhg+yfCr8xT6bTqY7e7jEJ0Ek0gkMARn69apK3m1EOFkjIr
i7yG2satJGynV10L6qN4zvzA8qIKVr6Mrnr8m4terX01f0R5eBMxapk0nskOSZuq
ydCV5LYt6rxB1D/6LLO2Bd2FOblNpWc+az6CB4dxutW8556TaY99uM62b+JgQbgk
eV9BvJ6uXoq1XecjvcvS0MaeQShrZvn9nuHRm880MSmIOdgWufSXJo7J5/qYLYxd
X7Fjth3wayUXtYFWicpZ8BOsaptm81OVS24wtLVIg6KefnsfCg773sfWoRysMgCY
nW7OjYH1jTVSrEs6+eBUQwPgHF5uywGi43SCbgnUWRmaQVc+YbC3OgAFm/yoriHx
h7JMA00N4s0bhlibA7GIYqhurhlJCMi7Kj6i9+NiDfnwQ2gn2HwvddZ71huCp5nY
+7ODn3gJ4zjVAxF4ptkEjMpw69ATpXd/XANYBDh/aoPjs4wZrzgkB8zEyO0Sicmf
cZOWDeh4770i/jUU03ddMxXp/w0ZqMLYPSkMbU3FAFphqTWTEg8jGPAHsCsgZd+b
k8fDgAgtCBHxrANHC3f/54LwXyHEewVHMopuSXZL0mCm+Of1Uki35D1r30NXrDtS
8L+7MwvEbKmshha2GhT1n83YDix9j5mlmU9nfBnlSSinV74hvDjSUcaqkK9kgPrK
b6PY3Hgw7s+EWCKwrc99f8qQ43BWWkw7Y4qP/awyMXv1Rd30EHV4y19B5TlbJpzu
b21eF/dmtcEW+Spvuv8G6YQ2cXXTT+Eg5rco5vY//FJf2QOMyuxOOiA7i36L5UeD
7DdgWEwP8T5irwKKqeIr5NNWmR0jbj2I8Kw/LHCaHFoPb1VATV98m9/9y/B14T57
UeHOtX+M5qV2OMVBAn/namSprAx6iKyNE2o+5bFhx9Pmq4XSNDmC7bM2Zq7IMB8i
YXEijLF2v4eZoxP9/y1+yaC3BQGm8sf0EohKCCr9C026F/KpQYsh+EesSyYD52HQ
dxKxJESpQb8Vlt/4bm6ldE3t2OB8tP9HzrDF4uWnFMZ9caZeZxE0C9fE/sssmcsq
A1380vCkBOaxjK/gDjDwwxFJQyyrq9GD94YDsIxF76wczQJ3qLv+jIYr8KCO8bN9
zQ3XlWrJlq2A9EPbE4CXiXC+dFgmvRZfGb7wBiEeqIxMipCT8AHLey9StAgYz5i5
QYFjjCJgsr/F8Td0h5IcUJggO05QBMRIGT3fDVRl/S/S2TdvGZyp8+VpJiz7kqVC
O/gpu3wu3k5qlf6n24ioEOE2Wx3rMoktrKHo4c3uAaJ02gFH9RLhuE4TfkkGJZw7
k0mkd0dlUTudkapI4RfolE3oW+OBFQphmZpYOvSwGCrcvR463Vqxib7xbHTAz5IP
cGld7F+w2aSkxU0jqdgTjjC7pvz546GwcU2nUSkYTcUiuulWh+tpTMf8qlslDxFA
+NjksUfYTahYNfkTkN145Gy/QOVGftf5c2hjRTWDVzqzwfSy02XBjQE3r2RoCmxK
jkl/hCfQ4LxI1yGtJdYnmTrE4+RybupXB2aVt1xB3IfGPAInc2u/G/V+ZNicxE8O
Aaeezkvb4kpPux2+xV06crA6NlcvjmIc7ud0uYBdjPZtGjXq8KGsgiHEWuF172Fz
1362lC4OzHVQfW3dSAb34O9/w/+n7CjV8aCkgn+Lj++3uOORv73OCxXoVcE7pUFx
0+UcwKLaLyXM3VtCdl18QMebT5emVO9c04FN6+e62i8eNAyN2RnB4GXTTg5jXsnh
UpvANYysCmhffRinQvZf1GbGRb5pZ3nrtnuoC7S0AjQuITbWVfzlqGVCiAhCjbSi
Rm86NeFLeY7eCF/kFy/6cmkKTifR6Yjaidj53eFcIUKw322ZENglOIgGECgPwP+C
roP+L82/2ALSB7WN8MdgpuPJoeLBev3R31UMD2tK9DZRWaUA5kC5VAdS+LdmrrUo
B3+rL7+NdCJSIhYGRhrOFECYnySmpDWYOApKp4bW3BFtreCsE72DPiCE7qQT8ZSc
Qh4NoQdjrhVD5m3rRdfQNm3czKnpDJqklAegI1oQ2coUNu14p6QTR5pPC6n7Cqu/
+U0+H7DSsCGiQOrCuw8sXvhuClJnbfAJL0a/gU2N2BAc24+pQitEjI6bLGWiAgwH
LHj6T7+IugvUaj8VjHzDfRpRId+zOX2HhFlmn+jLpJDG+YBO3C2ibrKcAht2Zrkm
Kx49+caEk89jV118V3XaTaFfUE10qihjRxIpPw9nfVZrwVNmnwFov684OPcrOQDD
mw82dLOm9+mQItb4j3+B94HlYeOKASd29VqB4h08l6dN2RAVOlCNTsruPfIdSTaI
ANN79ssN5BxZRece7VLTlJbNTzWSkqcS5qd7SNNeFWPAaInus/hflH6TmNVucXYa
h9b9WM6DYigFydH8HGTebFYYrM0iH6+sA7UTdy57TkR25fL0qtbiREvS0A3Tqkxi
ZpHFuxLtun1Buq72/COgPi37v/EfwpEX+a99BYiNRQEkjcSFzMxDhbslc4WdJ4I6
Tms7iIoyIfHQfGuibk8tMQT/hRoJEMVchv3POpqBzwvwWWy9LKrr1oGJGjU2904N
RYeLPx3hEtH3wPW1fXWvIbl1D2JrT9oYBC+LuSr7nLOBoYa0jmqY0J52wiHVx4wA
NEhgKqWfFdvKCfXvqA1x9/5scIGFwygYjmLWsjo3eXg7woIpNmkiQNn8j8b5heIw
pBEhPqBhs43w4Hi4pAVu0XsyYRt1kEsb01aeldBz53b/RtYcvG/Lvw90KtpwxqCu
Yt4Pw+sp9KW397b0b+XKyux+HKlZDE3iZo5XXr/hzqYtiCy8Lzwmr5tPKav5Fnfw
j+rg35pDzK1cdiTg37GbTLXgnYPUde/nbns2VpvjjaEZC8DdhKimMc96Yv6Wh9U4
wqvKtxE5NbToh9kUADpwdyREJK819KsvIFEbA4kDxfsXcfMIslRPArWRJKcTD39Z
Qr8THZ9seUYpcojxwjLfnHNCwsaa0+eDYHjMLIUNYjGxAYvkpcXvFuUXaw9tBB1S
D3i9Qwadeh0B/CCFvz4u5ublHgGztJ4NE6NmpbtBFii56D2m6uunWhmqlhEzyT3Q
wR2xKeEFIiCvXq/emH+HAi7okbCJCmYu/Bmm+E60alzN2abNKP5PiEQx9zl1HNsd
JlIJ2AKOXgg4lYFtK9Ui77mLTGgnQw6fXPc4flXef/PokJkx0VeuOvkq2Au3CwBr
YgyISXVncjHeiDZ0Xl8YoTGHrJ7wp8LlZmLBP4wZxKNB5jQjDvpLy0gi/1ZPHFSn
7CcHPUlEXAdtv71tEmQLPUvs4cVu7gIERrYuh/nUWzDp9OsJ/jaE5r9P87p9Bgkn
fZiAXmTCjBM1ddOutxZ3ZCq5K+SX4uxPr9uWmWANUgtAJXyTKz0SKtHKX2BugXUD
qBEE/t9aJ8UkDI5baZhlMfHaO0s0Nlt8qF0EL+F3qGJgB+oVWAN0IuTxs2FodiS1
XPYWva783ZjYKD6WCnLQ9rLI/gb+ID66Di3SyhagyrKNk5x/I4ocVs4yUzBTz6ke
KKeQZZ0p3VT8hwqc15ZEF5tKEXWJDj8sJGZ6kdKr2czi2CyFOuszXPcOwkJmAiwn
W78yyhMzxrso0trTXfDY1XaWY5G2D2nr98UYYri/I7tP4H/tRGNOjFI+ZoyEQbJ3
B6SPTV6XfDxQTEyDGPp+UUQhJlXW9NIRpjcRakF1z7yFtkyN6lxW27yoe2dnopgL
98kZfMTOkUoK/7IkmXeisvCOtsmLunnldjr5KN6eRN7PZ9JaSzsTU0taApmGrhoD
WsFqz3VjaN2mVTv0vKPv6Uv4psEaDsQdZyUaWZkKZb+Asjp+Xojr1jG9mdGkfsjG
hYtk40ZxpOGTKKNKRqT29W0X0A8u53K5BXk+lPF1urgtvoMkkfyDwWn6eJUIZ2ec
zQ3EN504kz5sd5UJOuOVTG4MC45pFAb/GwUp46MKkNsr8on1oFRi3TZeoeVfY2Zv
7X9+lFAwZN4MneMSK9j3oQLmB3Glnlf2FTwI38hN/kiVvnMiWICT69LpKur30Z0u
zEJ3EZIHBpC9aXj/KR2+/FJiKfIiyWvtxYVMmQZB704SfShucjyuMZlYAAirkMBT
v5ratUyA/oUSXc6czfWkGzBQfN5EQcOrKmvvmBQnP2x7TPuwJgjRHQSPq6FTfgre
oUejFwRzTIsqH31k8xwj2TRtvbFrntb6XOSs8jTqU4MitCJr0PePpykCEmp6u6cd
6Q6Akr4Jxtp0eISi1RdZJnCgfm/jL8JXuhQsE4AztOGojay+48wO3mj6T1mRIifi
1qve4lzjlXpwdrZLvZHCOsr6S3uSHmEmzmbGyG0pJWwo3jOiRTNQYYJNwGA1Bcbm
vhp/w9sjGcBJtRB9MJmnIaGe/ai1pb6EMbPxx9WBe+T6GhTN5ygq3lNQXL3dUldi
dV3HOOSg/ew6EUulhgbNBAVMTQdoHe09VeTe5UJ3DSm9F8a+wgwI7M2NLJ/HwoU4
P+h6WzNy1vDAuGl1uUFiYoSkllqRZujUOqLixu4jDTZFrj/2t5htHB6gQSaumeU8
iLso9fOBBu5S2YRzUT5ZJMm2r+4IDYjPQ5VqDCbiywHl21yEcU3D2TxlKCPU2x9x
aAzTy1EO6Hs3B8DrsG+46nO8siBUuToiRsCNW7pbUpN7aXs53r3iipX/lK21vaDv
cx+LwjL+bzi/dDSq3gO78PQ5dUhNxBWpVj5JFSv1PylcbmPWlgDGaczQ6T+toq0j
ZxV2DbFjNqxVdxMwEU9VdABcqt9L4TStr2BAnMIkV8+snJxpbVvBbWrNAhYyjmPf
z0bm7AMiTN//K0LxHJ3sGIiE3jz8GJ5rklbjjpTuxTh9Y/4nqd3masLXp2nOMtrn
mAknRsf2UzkW2L/Gsu1AkCh2V9HMnWaZ7qFSmFPa2MSSkWg6rHcK0pqw/fHQpYfF
o4DUaEDlSOAq0UG2W5Sy7nmCU6+J8Zrnr+POqVYAWh+IrO+QM1eFckEwKIywtYwt
nsNmo0LCSG99vcu11PPepPUbhIMjoEqnyeESMFYOKsDAFtQ4cQUH//LPqEqbkUB6
Ppq3ECEe34v1kpKXmwpBaSed++ah46DEP6sS27yZ7DsHdSoHgVKAnOZojg8CRSp6
XONVHakQM1IaScOWI6qCil66qrijLyWjz41vPf/GGeFzhFNhmPdBD+4J3XDHghKA
zJZdraClHMjGxkVbzNjta63TJbHQtFaPEg4D1fCg0o1q2xu9bUEATOPON2ya89UL
RDURKtmP/Eg4fFi5YgIffJp6t9Hn6ZIP2WMW/94bpmo+LabU1CMTtScYR6piUOnb
tIMkDx8cE10aqSCzpEXMTdDmKUgcCRtwHRHRSaquMFl4qM2CM4kEa4Pkt2gWW700
0d8nOs+/OcpU+CCBPY7ewge3qF0W4QC+UhvdMRjLYmkzntzzI23/orV/uaNGj2Nw
UewezHUlXAsGycId058392sXpa+QzYd4P5dh8IKGRhHP7ioqc5s0MRagcMM967+v
rRpkwJ02AO2BAU0JWwPah6rNk4S5oenVhzRFNwxx+PghyebXxbJAxhu36vZ5mXdF
cVZ2tTCHhY1gHNqvbQSN5OrSDbgdQ3U4NqKhZipSN+QHX4rkwyL4iBYjgqdDZ7Xl
neJZ8IimItizYT/nJZBJnE3/ltXoLOkQsoc0EbyzxAY5FFjNnni4625o6CkeBlAA
Oie7Tu+XeEdXM8ZWpKSo70WnS5ZbK8p4PJRGpmVeRWLeaX/5nKwOLHluIrfNeQc1
EMYqtdyrkZJ+wvJXpF0DPWlQ6S3237fYpSuMqNFTnhpNNzYfQvfpHzMEchEKoPCd
81dmsInA22vlyVL2HnrMgzr7DLRxieJsO9qhRu7PHAr2lGIGOxJ3gP1m8oUdVnGB
xX4Glv2ieIe6uNuBBeWG5B0L/XDD/qAgfAPf4N3SV/S7LK8GVd0x5GAmc9GtKI89
2amYsAwSLrHEblglK0GygbNW1mbYAb56gXF6ZcZtDXGq+8ib+uj5c9L9cjXGSmzZ
GMjQpS/tZDVJcdCfcrWAkxdvIWHD/jVPVUJL0yNokRLUK2MEluBPRbMAEljKH/wp
05qtSSJaGy3DeFrphaaClk8VuPWMjJNx1eaqr/vXG6UL+0bgdrwXwiWShKEBBynV
fq+1BqPlsgp6Yj9Yt3IK6BQyoKg589kdbq+T8KQ1VRp2FBS6BX/P8D6Szzp1CfGF
K5Jt7wnq5GnDUCJN6pWVspx4OLFr1MIe2QQosY2/NxzIhYklbsH0bIGomJt7N9q5
g9AUnKgLxfdC/2Ag7a6noHmR57tERSC7agxaHCWMa9TXhHTSjqbge3aXZ9UsLWuu
VmHF8b7i7VrTzoFZZ7eQGoV+VwnN36xNf8It4odJ6dfqDmhg5MxUJqa6G8IMQR+X
5r+YhqQxT81nY5CEj+V1p8pQCVNX9QFO+DiL0jYAe2niTTvV5OKIEWopBWq0NtPz
O0wpoVX+dc95Q2hjuQiaa6mAUeJ/ncrrPvEv2q80PWOWZwZN7/Q0C6cnDEl2EnMa
kbRlCB1Poq9I4BnsehYk1t2NaIbbJJqrrqQSsTFuPpL2yDwHU9M7nfkiDUJZ1gcM
Q4CMAlGBPv/iV2R4o3gXVyF5Nuc3nQKJPN0VjShsBa7hmcOCRUenuGIGYmvlnnqQ
vZq16T9j/Xds64YPZiOgLQeh0K3SxnLmtKnE+3hntQxDiuMtk5VQylpO4YyGo9CP
TrdNltB6wQqr+Lnlasn2ft3HJEKvg7mKg6XvBUnyKyMPKHkAEOAdo2Wq3A9zeL8z
9qaz+/H63Gm761oUzkzXny/DtCuwUAk2g+g0FH4/LSEAOd3Q8ybTRaXIDSo9R0Pg
/jS/rwLKBgczz+0tpsFv/bDMjNTWmuuKSzfveLUFkA5rO4GWTspQ16sfnu6E6pYu
9WViF9r1FmtrWK2jaUQWzY+eAumdXetfyR1yeJVYoWW/VvG4CnuyeKIdNCx+OaFd
YfURlVAeeIc3dy/xS6T2mX2SXDgnkeoCw1KqUzlo7mm1uAw8cS8z+dmXJzkPR3hL
r+c6pfUoW6w3TtgMqfvm33M0zBAxg/y+F8xzrXgYfFeHGEUcdwnfmjMbg9HtZVL0
xFokFXWa0A+pKZaVDDJrzEASQ6QGK1bFO1P+R60cZfajyyAuIKPVu62ugm4fdxdn
pn+HxYTyKWl3n1A/p0en5gq8e8E6dKroF765hvcOjiANF/djsDAQOe/DtT2WzXXY
Ql1M6IYm+FES0kSJ4O/AvLqw84yGDl3lUq46pFWbZXa24zw/AtZEBDCKKMguKjbo
qHryNFItx8lZmXwHdtNEOGrVieAR8c6cA61ztGPzcJBLXBB5cZ9WfRyqLy6NYRAN
hh25MNpqD69rMDjVHbOFfelUt33H8HnofoaWjVGNgnM5hvb6rdn6xp10/SlAVGfI
plSLf31K7zUPiaGPvr5a1Qp7OCen3+LlIIcePUWd0VlLa6Gl5uC3f4xOdcDExKYf
uY8ITOyghoefjf35LDFp8z9zhP1yAJs2wVCZ8K8G0853EiAkK6SXPQzE+XrQWzxf
FkGsdBKy78LePcc2J8sYj/bOVZ5LcqQkmqLD2hmrMw4uzTghYYfmmYYBgXDbJWiM
aSjlOUdU+CSCYwmd9rA9v03k4uXcV/o+byLsoUuH+ZDkmdbTV6kNSEeFBGFZbdF0
x7wgbdi0CRxEfmklvTjO/a4E33uqAQlRbdm3+GUzfaQfTN2GAlgj1rPvLz1VRijd
YTw++QgtLj0nDF7CDCgp3Al6+cp+/jLjKlBAZ8XXltb/noW9reYyQE3RTNWvAGni
8KVwI8WWZ6/7y8VNkDCiSwf9I2LeenZJASoH0M0vaRRwFlOlQF3bToVO6zqsDz8h
/T4hae6/5tfETIohpzsLX+Gr6MliV3XrATm1LPIH6w0LSpYxZM+ymzCbJ5Qm7e6C
qccIiYpJPOtOxHSaGo+gZeV7qIZt368fPkeg28R13dyMPt/S9oiyPJKVtU2gE4nU
7mBvKhFIBie2slSdnsfpEWvpitR94ASxVgpkWQBMQQZ2ANLX25ZYY3f1Yz406R1y
HV26TrymfVGuk3wfDVL8jnLlasulqnkTRgdC2/2NtlIFZjDtlgwuXA4g5ahFQgat
Htb/8s4qeIuBBfpbrNPaG/5JqozaPXHzf+GGlma0/Zfj/YyhJMh3rhD0EZraQ+BV
lToABgcdFhayHk0huzWVHKvB5r4JPc5Ufag/WsR41M5sdFm2Joh5hzIgCFRsnJUl
P1WmAaE4XQi09UPJZWQnF3kfFd4p6/J1pT4EG9Kg49D0uxiG6+l2JpYR5iL0Cq4l
KPxL1s2FPzOHsXhDJJ5HGA8mN5lL19TGwmvB78Dv8yLh8z50eZ2ai0SF2TEatr+b
3KHXaxtS+9r+Vz4Awn5yOSwm4TuP4wrbfaMflvYhRYuZRy7NkEPUQ5Ah5W3FiwSj
gPSZCf/EGOKKDqNxdE04lVEZg8y1g1kL5fRBwRwzga+ZMLv3xkDCKMmKPK3nAcWm
KnZ4N3SB+ezRBigcsyiSWF0hOS+R6mqH0cVYI48F1+u46E774RysIgb36aJQX0iI
AaohEF9vu2KMJtCoON8Mdjo2DhFQxh4qFSqKIwbQDCmVKqN1Tt4bhEj/4aNtlt14
zMnqGWBsLiup0GhQ0esGJKOog6iPQ4VJlVTh/xlKduwX07Ieb8csrBA7Vb51ttbt
Mu0xplg0UD6MBUKfQi49Ym/zWyoJESI1SX0tAeN9249toZuOq4Rc3J5soAbCBuzX
qIIsnwLV104e7pshYQH0lsC4IhF59cLm+58u8i16OBAo4oxkYVIAicjjCj0RnbXk
Qmz/jsqg6zEcndkXSppZ0dMEEV2rvv6bp3Gw1QR31jMioxo/EqhfAlgPRPHwjQ/l
24yivRGNKZYIZ6FXLvtQreHj8j2ShFiYHjOHshRyWIMHb3baYAWTjSNxwafUL11x
FAxi/clvntegi0dUZiDyNlcgapYxw68SUm6VBzuub6j9qeP067LLGeI5psYvh8nc
k2GhRzcVezU/VZVeor5mtg3c9QP7MZu4ejspfUP9SvE+R0uRmoD5sLczpesWH0+O
E4dyGEvUEmWGcgC0JjXuOCYEiaeGwNf1b0zYHVi4aHgJmeHbGkAxsaME/dlb/h8K
IDIDMJuoZ9iGnnnU9SQPPkC8oIIP1ubLRdCm6XDO5t7kD0TkD2lvCkiF9M7DyxmQ
Q+U7BkSPvH6N392zfc1bU48CCFNh5wcgeY0cybiGmOEkD2WvhoHGtlehzZPkmkJA
qlqaIab97CmojbIcT9DZ3wB+MrveQAz2UtEe3MNNxPb34SqoBmjF6PuJjfCZmE8L
jfXQnLqCGQfiHZLL21vSLtqlUvrGqET0DErbTDSvzL1tSoo2uh+sbCLz9mXsVPCa
/diBRTP1Pw6Egy4YB6+bRc++gW7IQH0UBTZPCbADbrBv+yQJ7M0au1iWh7qGjQOG
Tg5uKJz4tHF7u6ArA5XkQGg3kyn/tYztMTms1cLWIKwjFeHOjzy15hpeo7hiHTPK
wJjqen0knFDYRFULY1M9U13uKeL1v4eIz99lxdk3lE0wvynBAZU0SlFzNc5Kyu1R
6lyRkyFLEmYansk1hmb2iQKe3SKBgAGMvgettJNODk6i2WuKBQvrTNesmGNHnMaB
t3qAhjt7iUHNASDCypS0nNNFRms11N9LnZCQ6ZeKNvxpQHwZlOTY7Jk7UHD/3VhM
3amhd/HwtKmbZQkcjAJJjn1KVOj0s3/EqyGu3nEc7rbtZJtFOP8KHGWPrPyry4wh
t1b3XKPBVXTCasVp+yQcyAP0PVya1S3F8XmJsLdt6GUlCPxe4m5r+V6Ft1zXeWqQ
IRKCcs1+OejRX1sxbeZTNpgIssL3u0ZNIMLmwR6sIAjMM8SRtmxQXLlrV4esHRzb
zPxpUiBofV/79FHPKY5UpAfBBoLQlzPHl46joHx+wYLxycHyk3XtQ48V4HgfWVYt
3mOejGHI4jPsYfIzTZi8V/0T5bpquAERgsZC7/eFIGSGMOYM3FBm0HKjvjtUka7X
AsDhJ9H5ewW/zl+cxMny5vwMa8K9KyQNdMfoURLt+uN7mAeLhM6Sa1oMCofWDieR
iUd/oooEJ6YGlapyyB29a+dgJTNRerLRa73/91zeRDmzfuw5+wtlRLanZNLEYnWz
nNlFSZ8WyzF4XIcM8RqH7lGaCydpsFGLu3drs8LfYq4TlUSh14p/Orw23GrqQEKS
QjJXwkyYDqjEU4hksAHoptMhtKSFlOnRBuPSUAuIWjLqjFjUwPmm6ybh3FkH/2YO
xmHHQPJL55qdZ5MyUz90voIwdDgzj8P2aS4Hvo2N+UjcmDQaD2GI0s6uejPyE3wv
ZnV+ZTy02f7uykAl45RhYTfHeTSFYKS/ntrFNIrZ94HIcXrwILWjxelPD4w/wqSz
t++tvIbn+9aHA+DRY0lbIddn7za51e7iA8Ri6jAtQU79uYDXpXTWVaYOp4xdenaO
bCgAWgKEWdsJHXJOtSxJlm2FereCmxQ7R4A5WJVpBD9PZHnIxyzpfv4Rok/9IPCm
/R/m2Oa/lqcMCQK5LwMoLDxEgcA6/uEublkgDl6NiqJy8OiVecejelgKaYkSHSeW
++4qBp+lWDfoF3xBz3Y2RjFgk20VLfXgp7ggUH4heLqirbqJ+G9ObshRdpjE7aXC
4ETVVblweE8elpC5a+aW240w3lNwq1bTOYG7UD0ms38VYsRD8Oh5N0Q5YpvOlYri
i8nOjzB3xTBRY9gORv+GvQE3SFrqF+0QTjIsz4GcVW6KP+ztYYiRMqzv8rEr9tfz
9f2N/lxJXCrgPDzMFcCjAtrPJgeF2EpLJN+COEHz/dpE9ILGgnFY2hlhc46JHTz7
0wU0/3il6T0k0SCK+avfiWtalvCC1UEXAozYlnNGzvvhYOcGiMBRbJNXpqpbFmjD
XoJj+Ct2px/vqQOl9f2+EoeIk3ERv0jFB4ZUIKJg7LDGdcdd929uXXjOtqpG7s5S
9jPBsQH6pQEJWhlqWAaNc9Tztx2uw/r8/EXU0co8MAah7xUJfSdClE4fTXZ04HjJ
73fO2R1mIqRze8NdvNJ6QfvOQTK7zW5F0hMbs3SeSeG1XS5Y8bh7OH7LxNgtP2gT
g2nkXyu1zyaniiCFqrQ2XbNn69K15tZcWpqh6SyhYa/HesP7dGgNH0WhCUuQVVur
UpEDZkLrClKzxMK+pUJ+gymKNbxqiYlzlrGhqO7hraPNCr3w2D1udGjz7RyGpLND
bMjlIXGgGvl2CO8sKig2H3zrK0KIK/cWlSFGutBVuywUkMz63jR8bsgrpiyfGhma
ttaDHS+u6o898TFAAGjaxThsmbF+hchkTd8vB0ISo08NHYRzHOuf25doMeUda4xS
aLzUnTx6LchltFkr4xP24haO6wejnMM/HHOf62vifuH9YPSFrL3Q+VSrTBw9RC5o
cb37ItEE0TRQepvfPjEzi2ay+e2+Y0ywRxD2y4Cd0EXLWBaIYQtR6rOE+UJ3K7tI
2+cvMXu+SrpjEuedg0D1bF+2ojDDNpSPHNMTewFHAoesbODKMa5kxbz8MKVvka8h
DZx7OXtr775HFv4iWwVmBrinfvo7ntVOMkAg8l10p9+mfgLSivfcObQglzkkpFND
ilrD6p+oQmwZnXgSwGP2hhToyIlopCF7v93Tn/zSq9gtHNEoRAR4eXTQRBNk71Mk
Qfn2BEb1gX+xIeIt7fnNaCHN4/saFBI72x7j+3JAuXRrfFbM877pInO85d89JRNB
oTuN5IYV8d6Ipz61ei8djtSLmwtnyXZu87ag2u+eA3+wjiDRlikEqXJZxFvWN+KP
R0IeiZVNbC5BvZYB/mGPsnEzYQfjVdae9JtquAQwGjFs97qUa021OQPY8iQFCl8R
TR2f8I89UqKU+sQEfZyeQlRcTKLN+fjbmPpRzYxvBPIYAgRFGyghiGqw4kLR1btD
TaWn6Aq7k29bFDq3O1DivrVb43b8ZEJS1cqR/abwkv7ihr3wlFZyJA5nCPkH6jvl
9R+YVM0pyV4ZR+zbNVwQ7uCmXBINiVXnOTzUF5am9e/sLx+Hai13ut4OTxvNmr2Q
LObriKm28pZ/XLh6o5JrOZg5QXPMJ/vGSnA5iHzyexX7vbnRxReZYFVDlyIWcWyA
D2Q9rqdq5r+KER8ippDpf9p1nAYoEm4dG6jwEZXTy9DtE7VP/vmmaipbOnLzg7fg
ywALHqVBha2MLPPza3k8E5ZBbB13+lv0wOQWhvr2mcY2f6V8oOX5mdy8M6YOttHl
w72sAvbrZiERcU674uqie8Fp1cuZ8sCVq4QXgUUrmlUlqiE8BPAhJINMvIF86tYT
eW0lESVEZWY1s/fq2o6k9xxx8XHaUNvBmrZW76w8It5gBSpvril8XbcXMzqVRZXf
zrNGHmUE4+kcRPqFYV/ZVgoI6+1gNsKZPuPYBqNjB+G29nDeQMwTx5jZ2jlf2Oko
Jf1w7a0Wz837A+Gci5jxgJROZ9jEwu49hDRT+4qnfnG5WfR4x5ezwGIjtNHBumAg
YpozrpgmN//0OutHIqHwgtI2bGgkT01QLedWGZN3yWJ7g+DAPFtn3ub3sCPIHVYK
hewVqjjJApcf42kLCLDURJTqw4uMJvpdcDhulAnqnqp22+3bBj86bz4gFFBsrlj2
Yz+Riw8DsF7qm1WSjzPIo4j2BCBOlWNbbwmBQmkKdH28QE0GZcfO3tYoIgyu9CeM
DCmm+IPAY4w7BFTwiSi2s22L06gLMwMT/Wh1WHUHz2yMnTBLZj9OZJrVH7HPKvxx
h+Fc9T2QI1w2xzR5c/GdVaOnexIQiR1IKfo/PzAyLWOrt4FVig/0naU4dMc2SW71
Bqigo212T2soSgA2lAS2JSpmpDxorngUOmRnK9i3WlsBhbnuR59aPJsba9sSHNcc
nk7Dg9dfv4/JgCbwHJinX+SeBx9OAKV/obVcNKlfP7TbZ47mnGXbstKgTIIlV/j9
ynFh2RsrE6Cusb9d4jt5mo1b9me9yVyruSC1lYmBQcgEp8KjTV2cewKxGxeNdhC9
pq5TexYzn3UobEBvRC/9qp/ytvj+HKJRfWG8CSOef+2RpmRK/a57RVrJ4qHyFGd6
cCk1R56lIni7uuw/q7I9ylIIdbZYNJuuYWTgWgQTyoxUnX2i2JAGQIQn++na/QB5
5wDSIUrTdUSGFlZxjCA0vNISCWRs8W+MnoPHlItAZ6U+/dWTEpl53h3h66eD6fV/
etSDShY9Xg1/JYqH6q8ZcYJcCr1Z0JCt8od3xLlhlhxtHsECo/LtohNubZBg7WTt
xZLlcEi86Z+GZaxm/D6MbrJg34Hr1GlzPryMVpQIuf20OuP9BjZGecyj9hB5sWa/
tTph3mz3blIKHYywjlTYevvP/1ctabxhI9YFytJ73ncYzry/+2SSri8repyKk64v
hxiH1svDgukVflnJt5/gLDgfI0aMaXDkl5dulfTmZAmx8eHGkveodF/4CKxMKI8A
drhderrR7arL6Plr1B5XgIIM6wkEXwSpCePVwxzlAn2IdNP/QlrBXZt/xUfiELha
1DRveATWxa7CJDJSuIZp3YYNhLKrijuYhHVyHF180FOSGrY3dHLQrvLtYI9JHz4+
cyMCYUY7k7jheuTNZiXvmg6cKNwK5ohtpjOLcTfxcfMKeXxbk6hu4o9qAR5uEmn2
UgHMaM1yGjIV7Ysg8gH/ls9LNWDQviLZkMSglN9bqk67vSIcPHMunbzaSfTocevK
ip/TNW6k+HKk3by5uShhrPiITqB669AWCw2Msj3sLGxeqtofDqb0WjS79mHb5QBn
5Q5quQttLDw0PTxsy9vGrYn/RoYia2U5SnkR5FZ/C/aI8ryr0Ry8uTLKJ3oWFvUd
Oz1AJua7EDChO91pnvwSDfDQuMXFS8T5wToAyA9hsXc33OwoPtBiXdHZKO5NS0Vu
kBIUsUN4zf+c5CpwKYeZwgZqPa6ka2ryB6rInyT65sEWzXLpmYGX788xD6hD5coE
jWG9Jpo7b4eRv/r7J8uYC+jOzL+5034fI/ewoV0FKeffxnhH2t3mJTPUjvdxUUeI
HOTwo1CUtAFNF/K34MHgy/w/VAoxHNb8V9xO+1NAfjEP/cEePzYWkar5Obsdrsu/
O7K/VsF802dJoHeVfaxjetVzHZ8EQDrWXsnRA2ahRDrRrNma/FwO5IGv/Eg+Kd0x
qshLtH8CYS7NEOinLrlWXljE8vF4mw+wLPF1eeusGqBLg7Q8gdK5iLMpsefA2r3p
rVE9rvifgJR7Q6QxUVW+LZUG6s7EAcoPzBAuCwg9bquN2V07QwBTndebubo97U/0
+o1/uY2JADSHO6fbrAMpVb94+Js9x496OmngDp9Uw+toZGj3SBtYrwt0iawJWYuy
+ayU3eir6qHDwLhPvihCzN87aOtpqJWcPNzrcRgsDYRhRik3ajLZ26NjvoJ32a0+
To6BZ3wLwZ74l7S9zEt1vH44cfWmjIpjyn0plzqewAMZqtsE9tRrHPcWh+n/xkrL
1qc/YnhWcjxc0/dm30RG2YaF8X7cikTZVGuN+xn0I3JqXu/cK/NZ13OPL1NuMaN9
woxsSdJ5azuYd7YCBPRtyn/bCXsJQ76ZmPq1EW0ugUnCNgelAzufxsoQaVQE5SqO
DEKFdYh4uiOR6BwD89RcakzWzE3h1Gx0dEdkXcrGa9F9npLCHNMgsZE4yQqwzdr4
DSifIFQojRywkKdpyr5vHusOBk8LclY8xGRioywD5RShCQqO12NaVn1tp28+lU7e
Mqyt8cr8IWe4o7WYjMxtCm4tXp0oPO4lNz7KMFiPzolKlV4lklr1F+YxwBDczwtQ
mQtywLIi9SuUkJofzuo/8LfeJwtDPfNwUIHqQzFkxjyCPUpyIf0YAu1L8WVgY1FL
XqOdIj8HEU7LP1Rp6PqpMyfJ58d+VjMW9/vsxM127x0IZ5At09JHeRl8RkuH4UYy
2IOPPzMDTBgay2ONVsjP7HNttofzjGykmTBRptAoPWwR4lfIFEfL9HdCJvHa4C3K
frXkN5mN6ygvdQl/soxtHKTOdJww19RJuvJvJuWVEA8t5VrzHuJIO+bXZT7OOfXN
pd0PpmHP+VsM/j6gOUGKj9Ji+2TBTOKo4oO8gtPZfSRafVmcEnjtglpYqbtuzR9g
OBlr8u1aMYzsrSceg240SbTx9Ux3N3Ph9l268XczHgJNSlkGF7tqQCCfCPPD7SzU
R6+BIJ26/RIVBSc4gX2/eSJcSOfSMYD0ZlSGDSNtMHjUXCuhi5q73Gsz5YfK2XAW
Y9XS5ISIuZV83JLGFLYC78S9bOGUdtvtqkDN2REyre7BK2HHKLdZi+HQIOEgZhcf
maaVhzJsWzpejHn4QQwt+IHxJVQxauSFzVAQknS1s/kN35wa91RnOg32NCZwjHJ7
Ryzpe7Kp0lPe9AXrZ4fBdK/IzXwtcVbl2OAUnlZenOtCNsdb6wJ/U3WKRGHa3YF8
Cv+5xB/ZPSaVDsYM8rTHEIsE/9zPalyNrsjYG+rQqs0EIOqnvgGJullKve7ihz9j
2lv/vJtcZj1hlpKuzMTIAUD/kqiLgclOnZLXu9mooKdfmY4NCG0Q1/r0cruVb9wv
cDhinfy7Bd38CrwXS5Ss0IRnbPtbd1BsRMFwVqLa9b+OrSUJYCigVKsCESvkjBuu
5jkIU26nBn7ZFA8AKGNkl8QBotZ5L5VBXjPkm5h3EB30nsynl8Af8Saj6qbjVtC5
YQ1JLt8hFZ8SZ6GLOPeWkUkC8KAc6vDFrxJqUGd/FFbH4ZqIvC0ruo6j1raiQ7c5
ehmcUi55LlCPJkLcb9SqQo5PXdK4q/vV49VHRB30LwgXu5jcltFn/LrPIwBrSPHb
LAVg4XM2s8CJKtsaoXKOwfTT3G4pk385DNmCUcq77Sw+RrAQByMwW27CrXQ5R6z6
IAeF6ywLDCWmZjrfBCoB4RDlB1KkHEUlLDZAxODB3NRw9Rl/BGVGqWH/ri3afa71
LgrxTepBioHklGog3MkRKcW4ASH7xqbTtQ7ukhCL5i876l5OS3Gp1hLlUi+I9sA/
KpCVot9ENEYb/ngappPNkSp4wrslsfaVggmY4QG0Ilx2BR4+BoFOg9MY+dyvEukm
a0infMl9bRrNP/slIygmtkJNItLjzFiACBkRyjAS1gLNr7IyZZG9xuQaDO1c8cSW
Y1ZguecZHhwAYPUD7vM+yN5tGTfH9CYxNqilUaBILjC1MRSxaTCBmaAIh3A/DQUG
gIUSd5jk33L3vPdv+aHH+LAu6ae7QubDViB7QKfq4dFC9bItummesi6GqZgEGrXO
TP5uGuZqKw8SkvIkpYZ6L/gjBxKK5FvKKM6mOfsapZAPj4ZeYcHQEm09iXoVyTNe
w/Eh5Ila8I1fl3QmsN0sIGHlrnFNAtypHjchTIfVuNoDVWVAWc5SNOP5qQ2nnC06
Kw+kXT9EhX1PbIZAWwpLKq15HxhYb/CFRVA8KT6ZOdsldU3DmgK2yjZ5axBvM0V2
+77H/10iRP+egj2L6+GMTkvBFoajQtOIzSDsC0vdREihQsAksLm+ibTeuY0rK2NA
6jMTM3qvzuvd87UxdgLrFjWazSBFs91AjWtB6Y9en4pQuW0096JFt+a4vWV2Snfr
QKxcOFt7xWCq2iGb/reCp7IvNJywxFIocKRGkE6d6lm01Ew/lBbL7mlDbHHA2De9
Mxlk5YhkTCz2y6rRpuRZev5kTGTuvgOwV9HJz1Qpztu1PfkQPidmCKMK+PtnAjvy
S4XP7E2rpMIgyKT5LZsXfMkNDta88sgHS/NnSWItAqmkV85jWo55k5shUZmyCnLT
pPNctgUzC+JtXWrSdpyykXW+WToCjKtRFb5hblGYDZAx3D/gmDb7HlVGKHoZCt2q
KBhnMtEvltbFJPcrqYqBw4eNUalw7UCEOGYqNXSJChNSps9giXYjR96DT3135uYt
CY3mhFz8D4WbFtaANpPzqxsK+bLj7iIkZTLqoE+9Xjrei6/OdPo2wSFAuqSnmfon
OskKv1hTcuv9L1W1fB1r/U4MVn7abxZkTHBpw/cg2JsQSG8xvndwuu529fc4mapW
HAYzsBOv/ys0qPES5CH4RUPlQ7lQzd5t4Z4YLAgdP3aq7RS/grHC28N4zZuCYA4K
NF2uBm/17s4dm59MPNxu0/uuCRchfZ+yvhuvCz/t6FhOKUsvoxQ4wPqbTL5ouuti
UfPkL8O/cmK1zxmYc11btcrSZexTnBacqAKf2cec1moVwx79iFYHP1TzSqrmU92E
YM9zuQNFPzPcCWl9Nzcoe6LBAaGtoEFk7WerK9fz8TDnmTzeTYCkzl/M/2mLdSP/
e9fnJFMrE1/BP3Em9u6i3pCndOH5jRQd5+/8h/ETuKZsImprumgqfHNYUeiw1Uvs
13N5ezM4xHmmZOsbfNetQNwWX09AcpO2GCYjJTJaeM3ggw7Y7JMoJo5li4NeO6eR
hb2ypdYUofIYZw8hRhjFVIORmHN3ao4s/SjLqz9OhbVDhQZS17A+hReNtCNGuL/o
kHmfnRK8/2quFsy/aBLbKEr0Ddm+v4pdckBqAXz/B6uxVg8T+oOdk7OgJaDezMyw
uyMH0Gd6AXpjAP6KMcvvI+h0eBFmRSZ3aM4AWFCpBmXPqNeq5GZpvfcO2VUcEKlf
gPaiMBnvVPyapVfzHJ1iqWQgXMIJooqu7zOsJdUisFVprT7cdJmV19ue0nqITn1n
HR4Q0ZFVP07frAdQuY4orC3b56Iwk/mL5PprJrhPJc0BK3n/5ziRWeU83WqoyTIm
S/LZf3kl2ZJi2JX4H3n6+5bpkhlBTf5pXlGjbnSVkKoRrKWkWD5rpWKXXHHqzkMz
OeRfOZxptfz57Zh9HVF94P+so4edCthqVMWYTkCeSJ5TKFrysbF++XaVISivHPtP
nRo3/DWmmnTFdUQ1GFPQKOqlvdeNCaTruhvnlhzM3fTUL94Cy4KqyC0GOoMnK+nD
Ep9uZZz1cjdSAf9YaDV5Ex1xKqTAPHkgKbsTet+U46TsLMNIHnaUmmrG7iHvVX+J
FHULnJFvseUi8nX8bjNNQExagyD/fbQbKnVut+D4XwpZ5BPdTZGsoqrWJ3/iieY+
cHgpOfCxZ5JeB0497D4Z3JJrtn1wWe74Kr0Wn0vhXVZmdFltMmH5OiB/iUfqbaY6
oKu0eKLcoqzojMwcm/qpaPveBHigEqZpSo+SMI3uX++m3TVNOB4/VjMClkxjpmGr
DizaXV0dVYeiCG9d/BdMS0kF2WNb+waZI6Oj1RxjqmiT+7mqHd/eqwbMcQL9kE81
ZRVVYi5TtJPW2Ma76hkhhSlGz7r8TMi8OpWe5CEQkUfzBhIRlVcQ38m+Roukq3fo
oCzSKoXkUS8Tu/crjtc2dCAYqDtcBYuotNjUfLd2Nhf+wD0MSG6UkjJFC8tcDnn9
i11WYPzeW89oMKtdY0KO2I/XkLuUJYGjjWouNMZuIfs4rElddgYMeUVJ+MJInBOE
QSAEHLYEBZ5kZw0DtGpHz4yHCYNF4/j1eY6bb8yUNnkHBDbezxjzgBVxogvX75UX
VgBsibhtmHGiz/SLC227iR1sTmrQG7mSbqgKVO/oRVhaDFvJ6TxKa2neILxNSuSk
qHl8QP//oKmtI200r22/Yui20pV+6Y89bM+7RC+uK3XEEaDKTs0osh94z3dkSVKv
xyFI4IsL76+1ZZboYf24xwanBDHV7TjP18D+JlRhFL+H6RpenEPQ2bd2toAKFt1b
Gn5S8HRFc8B6IGnqDyc+ymLoKjudwafyefFM6MSUXjyljDOLJpzq1pOomj3cjRDg
9zn4YDIlwsK487R2Fz7xqSNVdjSS6Mo2tUnSBXsIYixXfooDWkPEHTCwhwAwYA8z
dkCQ4KbNT9nzwJ25dgRKZ6yJEGlmOFZcwTWN2NxgqoU0SPEuGl4Ol9CPqcxLiZiR
MvkWJIp46+EhyjhwgFrTNrQcf1zB/dJFHyF9z94vAht3NAwD5j0jxIR9LYDoQS5U
TAT1/cS5YZpPqsAplKHLJBART/dtcywUhDbmzfUlJX2NaEZaNJMq+RUoC4t4GDjE
H+5q8edhmrk7olNG1R5nvjdKXjMc6+KWTvMReEyn2fgg6Qkl/olTCoKvl8m/kc44
hqu/taFD+X/zp1qEDQWwoj/bUeqGjnGjZ/2Sm2Qa1LkzopQiOjoDIN7XQxJv5tOF
Vs/XsvAwqs1kNDiK9VNfpUGGvbUf7Vdf/Fgh8wIxZEsSsMJ/nBiMVljKO90u7yKG
L6jrbS4SvbUj3yIHwSfu+pKK3VwSllF7AZPWEixn7hNFxmI+vaxWS68F8kQSAjqo
Ys4twIw9Fihg595T6LTfT7E5r1uHNRh5n/+sU7eaypfR1tHFzZ/Ldb+aQ4XqnzJJ
Gzbyl7rUwn//Op0ymQriTLZjHZWGP/ersSLvuQaxpp8mm1LtvbLw+oNOHL31U2VC
MBFR8H53rOwBH+SXgx1I44OA6ozFZqsUGlfBCnEKAhEU7v9dEzVpx1fVoOtbACr8
vdmU7kf6f23GdqioNWiaJR8MrrPBZ0xR9cFP1sP7Gq9euOBkmqc3hOlrX8Ysr80S
igVxmn0zMHWp7kEFrBnFwQbkFowMxhh867Tr103IucJJZ6jO4DM3NNhDfQOJQo1s
GUOj/ZaLVZ5JsLOtECZIZ+cnQ/R27dsctXqXDDVc5UMJJyO/Cxt8M5yIMoQkYDB3
TCm1TmWQL7LV2Gvw1ReDX6/pm8qVD07Tg4XrjoStp9TjpJYR6g437vCYFQfcQmU8
g/H56Rhft8aNFAqwrqZKXkfOSubkm+PclmsCsJJEe8F9f/CGWUxJfE4VqsFyc4U5
cTmTq/QAuvV8bpcKlZGULcFzgwRcTY+S1aVa9vV7iiu3dlRxz9y8OwF5iICNxhQs
DJkiYMLgpYw1VwW3sYYdhuvHHn7HotK0ysJPSVs6ve1V3WqRrZTyBtxIf9Vkk81K
97javAoFVA6ImQyaH/40rdPCtQNtCPUChuwAzTy9vIN0fvZXTDXRJ1TxsqFCizuI
F7ASD9rvXVFrEC0ErH8Isl7AvVu3POONl5YmLyNhwyo8f7TFP28Lgj45Rm+fpuqO
N7ud2y4WHdCZMy6vu1kLW1k0pI9MgizY2PALUy5Cww2CZhLlHgOSxdfHjA7vrfgl
ywmravFIW5WBDpRL2l533X+6hEDoHyicrmKSo3pp9+td2M+ONgsTvouU6azHUknu
eHPR51Y1lBqLtaTVWvGdgMyvOdgWcRyPevMfMFHDDZjy8n5y1GU1UJA5IPrfT4pP
+Gsd3POpq6tup7eXy1pFPkDLrsrztHI/76Pbc344mzpsmOwPvjMvVLczI93Vkpzr
jSoVcGZNMi9OpH2R90rqgamRSlgPHT5+ix9KUmTGCHCOHys7tBy3JsVUgGaiyMhH
Cx+wc7UMXLLV4dlt9VgnkmedLL8ZRaSeG67LV64DijzU2TsNXLh91Qg81H21271F
AyMWBCGDs+aPwyvvf+XjqYo//dontXjSCkfra7CEKq+j95Ey+KEUO6Cyxspa6dEw
cBm+DgdsfJfgz23c2NE4oaBJlXSRzH20Ar2LY0EnCWH+PqSkklKGmRh+OJdPeHzJ
UcyMqousDQxTIlhUcy5wK0htu1yhrTD/MgcXh2ImSe/Zzfac60j5Awev0RGj+LDQ
bM/D+tMWmcbiTgJCnLJIqHu+zOk/PtV6VgMb89TwpaU80xTxQHFg2Pneg18hNbUH
FL+a374Q8N/orEGhO93sStaKcpQwDYK2VMQy7N0wXvm4NbyZDIw+FueiiB9wS+Lq
iuG4aqhFxkpmoYb4wSaC+dAb5RBLvORD8RU1DNpLtEFZGrMIFlYg2ubgy9Ck31Ae
7muDphSJ7KV81ljIUhymOF+hGe9jCX1UHA8THLTfbQkgJeXKBvqcYSmKXeUzs+ew
pL7l1hY+JTwHBk+TY4EU1hb13HX6kmuCzpnc5nFyCS9ttRBYD01CaiVa5hbp35Af
AWM1iwOplYlVmwXkamQhj8SPjRpqRoRfxzOWXhXQ5gTuquH41V9U32RmIAgGz3ie
YfDSkBX71mODge1fkHL3GxD9MTzex1nY7tIp6MjXSGdsYwOt4mwGwgvO5JbDDgTf
Vx0BKR2QT4UJoRPgoNOIWO7G0xB249yj9vCK6Ki5nBfDsJNFs4F4uuhxiPspLKRI
DYiABpEGui7uIEoWplfjhMAnQhjNacfO0L7tQ3HdD6jTwqdiqjcQCG/8Y5kg2p5S
M4gPT2VQoptj2F16hq42mR4JxlbJ4BWzJ2UIGOpWnFSycqCt49QtgM3kA9jbMlCY
21yvxymjVDfkmfKrS/ezpeTdca3p1pQPQMNBxeqrr97imlb7xMV0QXf+tL/FKMDE
0R6+ZQViHxTXOJtwZjgmfD3CA7CXakKxqTbF+p7IhAZkhji3+twuZ+xCd0g+lSto
Fqg9nYlABU5fVbRexXH3YR/jwRtE2sHIfjhZ8X/WuAF1f5JmQVcLECGCz25svPVU
Yn7NnHX00LCUMjPM0lrLEu1JEISizXM7yl+O55P2xqSIhhNmbY4wTxIHbtYY6KYI
uYKX6t//YzCW7GD/NCi+JaOlbPV7OySdNjhDbeBJb+HQmfFvwFiB4+eXBprhXEif
SUwPy+gZgEkiQHyp3/2j/Uj9tuKMoLT2NtiSSES9pNJSEcPic9UeMH2mE3hknYJu
adxewK8ldAgMRAJ+Tu9oJ2Ws9LdIvBDRcYvdn8lvBJwr4u9Hizrr8B7sOrIj5A2h
PSURaTpQD7tiMuTlTHfAs+mRMXpEMrr8RCKn8WW1Ca26RR1f97JYjUlDDJDr8bbj
zYbsk+zi8C1Ka8/KzFflZSn84w888Hz2MgaW7ZmWxwnvKeomgn3kktHdjLoN/tOi
2XVVRtSO78o7W/Cow7hG+MfWQUX7DEKQVdGEwYDrfGR+fXAh2pdEY8FQucECV5Le
MAwQP7S5Jr+qFaxbyQWYAOsWp8JBOs72tdYTc607Zu7/NChffkZG7SfDrqqCKLS1
w88jR0UesAiVyTQSD9eHPZgB8ZIelwPqyHSnrUCI0g75kf3ru9uYu9st7l/L24QO
S5UNTseQ+VQW4deUnT6o3+Na788KWE2Tt1OviyjmMMU/UJi60eQE5+24FmPzN97Y
wp+fjFoAHlgpg99TEiZSvz3o26Eg1elZTqvqWBbUefMYxBcpdNpPjWZ4d2cwzm2I
fHfy90pBA8zDoHZ8peyVxJhuERMhc7C5nelNklhW8f5H1g7fZK+DJ3rg6N5ctdrw
vaNx6YBxPbNZkSQUIhx1LsfzH/sJI/gxI2PNMB33TzSReiGfzkxDJLPBAcvcfHp4
DQ8FAhhISr5HCPR8XdXXQHoM+UX4IURjgdVfhIz4EfEQhz13J4qU7cxGAm7vvbDK
xYLiPHGkSJ8X5ABGgG53eR7FZoC83U6JtrBUSl57iKuSpg+vLJq7jEjO8w3mQUsA
yr5eJ1QYSkJqik91AiTet16qp/86TKxgXfT0RbaNlhd7LCH3nNj97x+2McjqBFpq
tSpzx5PBKfSSAw0OLvtYd893ZbZN1f0WD/18OKXS7XmPLp0JbYMAC1FdR+LTqc1N
XVn3Xd4GR+97cNKVxX5UefzO+zfGIZF3ahmBrqjqU9znwwXmPdOz1cVmk13daNu8
gGgMnGPGPQfFagV9KkzSbEYVPNVaMjVWJWqC3YH6n+0hhp7sZerkSJYYgccdbwF0
rjoPCYFtAQs3J6eXab8vEPqgNvyIbI+lkzB3DcorvYZreK3igW4wQnnv0SEQWbxN
WQu7BrenhCNKZ2IE/mNjtCzPlxT2JVqWKLXbGnfjjoFizKEq7lUXT1NQydIafc2N
H3IVjDTqrBL9yyXO/35eUxB+KDNu0DreMZ3AhuydhByosSdUAwfOJrhgTff4v8IV
I1oPtxjV5BkTrdQKiKUlmMnkSoBneA7B9kP5HY67i4VOX8bZtj5hTLT9Iiiieh3X
unu/yYplVk12fChh9xY0AnQMH8xj1qRXEHU3A2aNjyEU4P/OFMnbvbxFdOd2lQjl
yk32xqt7mpKlFVP4ezOABegbWCXq42ESMc7FENQGWVNx5Nk1NNVxkpuMP6Y8UKgt
S9z+d7LLgWgAvr3rJGyKuvVcpi47rYDDpq6WBdAnm3H44IRwMh5hufNVL+uVkKgi
4wo5JY0EnFRVLUvUpWc4Sozp/RZj9RrCCsL4uFBcvuwflKHXGzNpq6bN198y5dNm
4+kCiUO2EUYs6pgJmBK9p3cTr/ZjgwfoAdl33K09PrKDOUvV+sRjdrBfrUeaHHV3
4hpIMV6hu81HG8prmfPEtryVEIo/SJ3FE95LtcncnypVuta/zyiA8LtoZvjDnNBJ
Sgb86H+DpH8TPHZlffCedE3+G2N6Gys2UTA525tlkIDgsGyBHwBN0oYPNK8h2rcw
f9cgyDIZXXxiWhPeWYAdtbL86rsHHBaGB7hwk0EwePgQRBXgxAX4YmxNhxAR1Zhp
Ei8amNfpG4WfMiaMCtXW/ceEXlcnaxiDxRim+lsd+9qnNxyEi5jtvhcsnktqFwQq
W5IURN7owDhIVRHPAjbTKPVeZC2lRDRL1aOSyh3RNHqeVlNakQGmOuw98Vdx6bXT
CRTi03m+dLiCTN77iZiRzjGGJjYJXD30N+JWpt6RbcKO4ePlbJbAZkXT9I+JbPRR
UVrOcPxITQgdfqcBibbkfcG8Sz+8PvWrXMXKX8JvyMj1iM8ZS75XKXsQS8S1gtgX
nCjIEZFB5gCFYOjjwjGClx7aGJ8YU09jJ4SFpIHIMd1CocZlxAJ5/4cavsztzXGd
0q4HkA8pgbZJ1o4wCp9fBUwL3dG5bwIAEKQ2afxVGXgbZFMaS9yWvqWINRhfRVMC
xZbH+Si7S2B67R2n8X3oI8Kg0l6KAn1dIcLorjqwqJEQ5CqosKgY4LJ8j2n+B4de
nls4paXMuJAKNXHOliReiBPwyHqYvNTuaMLBax+fAkD3rstGa4pb0O7NP1e2uKnN
X4O2KZWX7ZP6WJ+IqBddih+AO2c8eVM5w9aTMJadiVHqP8JePmaeSidOtseT00fH
8rKiJIkqJFg/kKhRirt8H0hvGSl+r2qM9pbdD9KbtDcZlS/MsgAwmaa0oUgc7O+q
24cjmqfVnsitYZOU3ejbUL+uDUbTdB7cADGt5ASPPpqKMsoSarbpfxE8+K65Ou0R
H0kWLWCTfF8XLVeVVsMQ1WX3vZJZaNuyuW73EPg5KpwEonyWgFO8H3189Ru/iRH0
h0+qpQCLL0SjkPAdqGRdTCrz40u41InwWtgAr74Kk37dQqvUczs3zoo+M0PRLPcB
naF+Y/2CmU7bvzycZEollMWAz+FK8hPcAZU4TD+1HlfgLKzOC09gWkRKv6vyAmny
yANF6ItPPE1P5kH7p0IppEnQUKU15RzruFiPvyv3qb6ZmtjWkna/deonm2o4UA3l
NDzta8yiw+SNQl9I+t4LA2HQdUQ8ga5TE4IzLHzCPM8G7kqVKM/eK4HXekLFkg4H
5RPiG4PXGgxgmeTOOnpY7/9eCsW+s5y3Mxo8ANBGCIrJXjwWG65/r2w9KODosBTA
1Twf+TB+QLvHZjWR3b2cMEzYdHLeo8jfczVJna9AN2PO1frCErew2TU3V7iPRXi/
gSGGPtDWnI6NCLdcmSV/G3kLKqSmUUb1KfTeP5Vrv+zWMJ6Ck3+FXW9gR3oCx0rU
XrX0tQMj+KEVXFdLdnBqb7txAl2q0cA3mULKB0IceuDoSCWqxcffCPqz0OIAXcq9
3egHXGvJ+WDZBlmkwBj8OZW2N9zKSl+dDDzWlDFFDvmRWOqhfsbcv4IzDjFpTeh9
1O/Jz/oX0gxzbl1oEZ7iDx0dERZP6h+j5qGiQmQyRCgYuz5QP9zVoOdQyEGKWbqQ
S223A9zcQCCI0hdp5tLNVmgy4MTcS9FPSFVFIZ6sPKPxOPOXo+NaMfNgzgqiKXSB
JmichKyAgQOwgl22VbEkz+dtIin/nTS8ukt/cm4EvShBcMe+IwU+W5OOAikbk1v/
SLggZBbA465DRnQlMF/ja3S/RCurhCwmGtmvaYdWl8ehlwJtYSHH4rYCB+NbO8Jx
LiOy18ztl4Gs7ElUrBdSB67aG1Y8ZNHkc4DgwlUE+HrxJsUpdlAvCcMubCA5DMCH
xxL7K9MP0aSyEdXIQQB3zCIVyy/4gtjgFsVF0B/Giv8EQQkaBCEfzE4OQfjx8ld6
+VwmwPrGBraq0R9CyunC8zI8ynbMc/jRauj/iUXm2hrt7zshRfyu2x/GNoExibBZ
Ymhcem1RX8UCq03XHku3eYLUD12ujpcqmaqFerGgNAVj5EV4iFDyDtmIBjJkHWIa
+3DOprkszUtwh12Dkk/9SrPnfPQFWIfHjZoZ/AOHhTDN/vtMkhzpAAjOkn2fnt+J
iZiYMyvM0y7zcSbpkRczdVsHVYTtLl011Of/q8ZOmaaYqroMMaC8Ae3pF2qUkgOd
rn91nDn0VsMK5lupMkO4Y7fG00zJ5jsDxja/AY0mVS+fW3IkBfNWJcCDBm4pUA1Z
tlgtibxDS+0hRzd1RvMJdNfzwKwoISDFN+PO2aQtwTO+zwappqtKl5kNhl2Gox+F
w9wcvSulDgfPa7vOINDdwDyHdXRPP1HlM3qqvANJqeo6OPiKL30fPFU3WP1L5aZJ
4je2QJY4vsl4rrGwlSjD1ihYInrWXu5Tfs11aNGjP+3SDFKtbIQmDgXxNq2Ej3ty
rrrtb9WsGtDQxKFGkYkEihE59Woku9xXBLG8BEx9D4YwlBBL/vXCyvZIFRXn8In6
3ggVR5vVsb8ZTfS/8Gw7OYBT7PfOnrB92Vwy0lr4GBDK5BA+XNGr2BZ5BgQ5PfAt
Uju+IRQma1aELwJmJ/+J+OJN6vk+6YJE8FkxTjcs/QNAJcV4ogYBWkR0FkXd1u5Z
M5eBef6LSAd1YAb1Uc55w9zdoXw6jxbtpm0ir/Cl1AhwI+tATr67ptZ5/gfPgVqe
cqXmiUJGGdCoBaWiguDUhF2c5LZrYB8L1hTOeU3m37224RmmgeRvNi5j2b0LIQFA
+BcdYkMpdl84vC3OVSwFlCPzZ9ZPwy8H8HIOFB8LbYJLTZKj+LduxXPylsytJHgU
S9cLtzPUpYDqBcKu09JaMEzPT83aiuhqKRyuH86uK5wmMepagzrVT0ry/hbXNZxx
58V6/wvpbYI7yZOEZrhgpCuijqce1Yi1BNo1bV6JCxF/iEIl3BCQyFMao4AdSUw1
/9pEl8N6KQDaiDm5/pBJhcu4CX8am7vhzkRORBQGSy0AJjNv+nPI77aFHYb0QqQX
0RIogoKlv0jcoqYmqbD2CkLDrIaNQ3EM/i0G5GPizjCpCeCX6ZglovJdGXh/b7wX
apc6N5REsW334pY9p9h5zp1QHTgRqdWG+xzEcIfV1/UOT7Ys6AF82JNEdSM6MZjj
91d/FAQGbL5Ksj4NmRQk++o5neRcW1OVbJeqXy2C4TApl2WRHvcnrCa5iRsnfJmw
dVxo7VBf9sihP1m1+9IdQYJA9ULnocXh8T+fY1ynaihatGvV3l7+SHK8+5Q1GFTT
RG6Bn9pxq3/GRXTUyZBER1Ox+NWnAgwiN41aLzZSMivY5In9Jo8o5md5FReKvVrN
xSr0l/QGr5B+yqJtfeLC5YI7qSL4MfSaXwxdXCykycnuANCC7JA0W8ALgQYDa8B+
Nj9RPxHHW/147OQox9b0eDpAnPTtLMuQT7XfmmtL7WA8GfhYUaGr0V7N18NR12SF
ZPT2xGrbm/HouvR3JjDB4NqEWQuLvZacaH9su+XRAtVCO+KPvn3XE9LBY4DstFT7
9k2sgE4ZcjogCKYUiXKOS4pdc3tQHZjpq2aKVPBghHWvwsAQwiy3WjcWGbvyLuZ7
tFQzIUpDq+15kq24MMtFe8A1im0GYMBSKvVUbczTMAfe0f5/rVP4u24fJ92c6H2L
CtykOJNg5fZSs1HbRVur7KM/AOfvyN7Pue5UGBFdHI/3fW+Hgj6iWBaO8G9VmNfY
RLy3BbZyMjGL7na7MWf0e6XiHOO5Wx++HbxStC9/wwMPvAUXoQKiQFDfr2TRpqSa
o9dri2D+hXwynVvGXnNlPLzyfESLCfT3BTBL9PNCtdw6qfMxz/baioqQ0nio/Cfw
NR5387x+JwH4fOFsyV5O/K+s5rjl9Ulcc+AQ8zlnWegbIrItBTvVxvKsosp9Cicq
qow7aikOM9dmTi049WDZYt8IZgCsdJZUZ4Vni1stQXoUSLWMLUal1bOlrvrkQGCJ
W7MoX3e3k2Qla/9KRFbv80A90pYB2DTeFP2JhSzo1/AFEdsgqsNek3GHIWjta6vW
pBDMIuZeVyrKNsrOG4mZTB2Uqp+62F2E+usUL7mv5gnN7yBZHNTjU7F9KCygWhZd
uIAKghEPxGZgn07aph8DBmn1DsouDZ6a3jZEklh1/Glpb2+afLehadPC8W4g//yk
P10ywdw4xOx2w0bGbuKwFFghca2ZxQbHb+W21oPKknB5Xf3z7MpSIaAs0CALZduZ
v+ojviLGelf3TwbxJOFRKJa7D17Rro8SL48SFwfKbqcUA1cgPeqygihni5rZ2gW3
GNmGAQk3HVNzTn6qaD1zjbv69Zw3P33BO4KWHw3GZisS0d761b6tCpszcGlcOjHU
h4gmHb+FIsJAZWMBhSz5zc/t816S+fxyRrsHKbS50Ibi5g/8crY2kXjKgabIQV6a
s+PkPzPWKy8FyNqlBVu8z3V3rQwPRm5Bhb7u/nK/tad3oMMOictaUbOSPji5J3MA
eFEowXPH1du1sR61fE1iFUfRudr/9NE9S4jZO1EX4RV7DVnp5w3qPDM4JhOt2XDs
3aW7Kls0UxB2ghm2shnHnCxtlm8tvayglBJGVB1QjPfGVAc++k0VZSnAfNvsVS+P
I9z927fChCVgGyhjTRCc3kwS7dCioK+goJDe5zJHhMGW+llDmeyINQ2rEAqA/USo
N3JvaJ/j7E0xNcb2/NB9e/9KD3BAgt/vp//yDbPQqSF71epuCKpC0k2nU8BbtJu6
upHeA9SZjCWjJ1QXZAmwEc2Njj5po4Esx0/rinHxF+QK0fzmposEbddXVY2EqGom
FEEDtK254pIeiKciR2+hu3qCngyfE86GxPfanku3lRkSRibnoMGd344pD5CiBGsx
Xxxhgoeji0Oa1kbyeKu3wWu/aMXHw5E8+CWQkVJNGsvGpQFYo+Cgrm4YfYOh0+5X
5zpAaXiq8RsO90PC9Ga3SEzKTsubdCkAhkfIW65s3JDHFWhEQCveXMzEwg/EVnN+
yC7PHaVwxfVaiKF43bi1Yyoprq5kbk4ekyMdH3NfxS057bQG3A2D8scCln+o6GRp
RSEf80VKAyPHktV+oUvRllExMmJX4LDfBZTMU2dbHvMC8PAF7Zdpf0yH+sxsvRki
gVyrmRBbLzFJidJ1d/a0qy5fzitVznNY9rXEL8+88NS/yQkoAvHUm4oTV4bI56/b
sJ1jEhPPeDaGeexO25MipcqXb/vkgbBUasdOoiE8+Yfdg52hoW81WL62oBnhwZg9
vt1EPI8WB1F4rIcNHKN8qiZOCPESHT7r+ZZr8AWnR/GaavwTWYdy9KyvPXi73wtD
DFLepzBBwx4KBgkx4xJhXw3AQ2liFCiXKALVhlmN427SVNa9LjZYCfoW8clk7ZYr
vOzWhtTOfeF4go3J8HYYdH0XzIIDDPTLVp6nyv1WYsDjtDUzo0NceX57iGx1bu06
Rgen3P1Y7D0rAmMxyT1DTdzE8vWXMSNriGWhbmcE0z6scHxl5oRuYJzEQo4TmeHf
jtzI1fUPhp3CyBkrUjrhcSk8J43aB6E5R/7TfhiP6/4Y5fbwqxxJxN8zyvs5mzD0
B0l879At+KMLfrgpHz818Wsi8G0PvT1WtAFKRn6Oee/9cknSyK+VVvn2mbtN9BCQ
P//HQ0EGtA8475v01hcoxM+jKyE6qX93rdFlp5nI07prAVCqxJaxsIYIDwB586j9
1CXgY+D3d3bkAvZ4mGKDjYz7bz5LKqCHE++ZmFgJkekRVRYE7pMmxKB7r4SXHNFl
3xF/P/N4DV5neIyhs+RI0Xwat7TvNhJuqRWzrN8eIFCfRe+3yh57USsxWDa+Z9Vk
eunpCFkZ1sBaBIf9r0G/1D1u66HUq0btZqNdWnmy2+yjKCjQfDslg2Z+nfo7Pp0c
bm0rLmusMj/w7gV1Sx6gEXqbAhXeXwMSoHUjwjhpSvNhpks1sTT8+/x56kOjbWfl
hgQJpSechiEcPJeY6ZAJz88L837fnoiuUZ3zssF0v6lA8WJGUqsMvhGnslIrTbAb
yA99puBImNDh1tZLzqElifp3V25jLERKiJmdkVWXT5dXxftJRqN2AMjKQAoxrX1X
cESbeEr30mE4oAkka78wiMqfG6ZF51MC47lX7S7y1gtB8l9dhAY/KkeE1rUAXQLZ
bKu40/MGzmdVdJkvkzVkt4i10gLVoiMkpIG91SjVbysN5ASd5/lTA+ZL1nioS2db
YffBy3KR92+h+K7rkMm5h0//k3Ca/wXOHYEiTzFN6cr+sm7hiacpDmr8jcJJ5qiB
oKn8r6YDzz+kQy/OdU/+P5fHdRHWqT1qf+mFlDmpsfOtdRcMJigPLBvGbOprHw6z
qwR5wj7fTXdCdYynxe63NF6M6fvuxXmOPK7jRRubpBgDnc8pmj6zn4oMefgrXpWZ
lEHPpGoKzoWBSC/+HMlb7OSI9bAISE4Ajar65vVJ7mfKOq6d/O0QeGi+36RGhC/X
sOlm9QQZ+l/ZxFH1VZzBmqhAAv44g2oL04Duamq097KC83AFB4I+eKCLC5XKC06J
r4eYDBkSZVhO550E626nXgZKwGsSO6Nppb4OVvi8gCqRkZTHZo9QHTTDgiPxBpo5
gSJw3Jg2pzPxfv7RRJOkR2HuqJvcyihxUerFX07z936WCvMWKwJZS5UW9P2RLjlQ
EOQre1fSbg+BM7KrRinzYPLt2ZaAVrkwr7aWnqaC5Q9PVwv3z8pbL1ba9clT55FR
G3Mt/J+eW+ixqZNl/QoifwStVANmJvua2KjNpNj5/2R96jFntQQ0umyEVuQy6XFh
DU2+rar/iuHQ3hCsKlsF6kvq7OccsX0LD+vDv90lFC4bRwL9Wd4sRGUjDvQ6A3iH
/OP0HbYuv2ucA2SMF+SoVDvTvPIVKSr/OmJx4osnltJao2ysXhLPste7UrCftQy1
dV8jU71KFiMTaMDnVUjrwkjR3fES48aralXjyxn7LZdsuenujSAkgG9tACeW4UH+
Sw3gXtcjBu3Xvw7Mlk443FzgVf1RmMYbQd9LGbPwSr3H9obhAhjRIcn8QWpwcliV
y4ZHmINQWaUFntvLmTT6LhJhadDLxC0Z1r9w2I6qKdkQiV/U8piW6+7t0J+X67iH
fOHy1qlmD7GHQ1s3VjkWlnlmbMWjDS+VjycJWOJ97oAJM1MGJjCeDUouDo8KiUnL
BRyDzdnnwG7rQFlQkTl1LYKM3WIcybLv8s1LVwpmIfGN8d3DWQsTi0SLyyc9BdLz
SgwVOp92Z7XDHq+rSKnLYRHAzQjNvx3/rdTaw58Tev2AyMsnGHLQ5kIs7dJC5/RA
ckZY9dtJrabigW6Mme6/WqRGW1QPbMuxqpYNuiD572z4imzd/BzBLGGZuQ8Asq06
S90lYfpi3sCNhPx48/Bxg7x5+KvUnQxIzx2ad+3Qb/pBd6kOLrUzYS8lCJ0Ndy5E
1WbXYVOg+nTvuNXTcfgqEnZFBM5xavzHdgwMamk8LXwPnm92vgIFtK25h9lWjh8Q
OdUE7R8vBI6ERZQchmuUf2gEQr+qHLTxczvBVMbMrsHpIFMuu/NXsUj9zCLYYssR
LLfcm6rEdg5It3rKiaucxWo0q6F2fE/uMBDAWFrvixmn+ITQzT+Tuzg4zjl8ilzP
S0HSO9EBymy+y7OBpLNbnEDZ+VHEbrewPZmNoauQwnN08JhM/OggOkWulTVkFhrA
VzNMYn2w1W2Kfp6hzdVcWzQHKECk/ZndxB7iZ0jbqDqKNxleODgf3WU9ChRHi2dW
MK8ySMz5IIl21G9PD3LyvfENoAJRvi1x0PaH2rU0yTzo6eDg5s8tICGKGG1qVsg9
RvVpQkvyppZdd6nyxIuD7DtcUzRlITCvjXn8wBa8EWzCHCMbAi2C+GbHsvHAOh0H
EiafF6PyinwF7g3sh7lclO4ywx5EixVbCoiCgoQUtmUoMm/ew7bdatorjvwqquHC
JKDKPuwHMFCj51ZUrFQY5X7Uxlr03pcWUdKknRvly6D7NhTKxadsc0dWlWDdXkQ+
U22HGUiQ90dT7A9zEfHNd+qmkXXY42fgebK/004hMSnndYoXsR87kOt7OypC02g8
uskD3DrQH2Sxe4l67UN/BrRmuB+w+K35DicjxFEIXMxinp7BUsI+6pXFkpZb4N5s
1RrDC33gtMhxeoykudiESx8X8jfshjKbv6zofG+AkKZdfyQ9O2g9JHypGiJgtMYx
4qdeN66ejOLRc0CSK1GbnvEIMOqAC7RtAOdVGf1Mtaf9ceokTKSbwzdOX0jg6gnS
Vb0YMnwJTfKw+6aO6c0W46PmzOQR+u3kKtxD7swCpTAGQ1yDmaO3pcBj5T+cC/L6
8qUui8QayL3QUrr2s/sqIdy8CwjWsMB2LaFyXf3WvY1+kUdTfcIIKnFYVKEQPT0C
a22ApAAsYTWWlInosKyegjBaoz6w1I1qlKuC5TsklfZwmkH89NAzjXowUSt5xnsn
4qOOPGqQ1kq/22MbNBWM5RbClhTD6H/S7gX2KPbcOTeNtEDyNFv9/DgHZZOPVYjW
7/znPyvfN8t7IhBUEJAHwI9E5+GIFz7rd/x8GhuIPNl20GPbruEBOZ6WRs44MpT3
v2pK66Wk3KCAVyn05j3oSbWO0MtXBhNVM8s5vDxz+4RyHkekWmjJsAIfIexxR1uP
9BGHlRMWgF6um8vCg5HUjY1sUPerhFrnYMbts8HM5ZmIAeTijURIvmwnh16rIFGg
VsbDH8P1ElOncdYU7d5PIq8iA/W8TPYi2cyWw6Hb2Snj8LTEdkR4g+Gbi28whm2a
V+cgW6B/k03+amqagDswDKduns/j4IcWT6GB70ELr7NxtTiM1+qOdpBtUKj0r/JV
jSjVpU8ic4vpGUsc54pxggb23B0AloC6T/cbijonR0pvhPtHm1HGmwl47Kht7Ap1
RHeeigrbOK25dPoelDIOPwvAwLi2fykA1kByPKR3c7bv7S7u6gNNRdHqO19bFIKX
DbLwZDn02jabv7aq3ibmtOcNA6Iz/Yqu5lmOotMnseZ02aUzGbnIDbOvFhK80Xk2
CZpWFvMSacPKHvwDC0dpm1oMyjXzd9laIYNCsOAsYgIPglTr6NMeEHBCxRRWKZsU
jqCltqfh4HMC1zZt0SHcgEVMcL7zFBWlVngeBUpbNnQnHD7P2/dMRIxWS2hTYiVy
DcxoIEvSn7fyyjhJNQM02wDxzcCIG27AdB5387KKeJxB4y0le0/NLHHscZ62auF/
znJjsCFQGOAuwDOE/25Lw2sPLs3ldDGbnnQS6DbWWCFgNrNyjr50wEKLebmD2mwY
hSM01IilV+1ZzbTE3/o0VXvltehx9L2XllBSc5Q5bh3RALIYCaPaDkj7ChFDIdjQ
Xb8Ib68/m1tjt9Tf5p0l/G579ULt08zh+7WZwd/HQb0+qzed2ZUGVhFwto2FczeM
OhHoFpvSXmxzlHZgZiSRu2LTqP5G5GqcLLSlw2//4RtRQ7ODHkACjKP0f9p3dHAQ
q0fctKyZUtBSYISdc0nhk8OQF46OoZ6Ouufcd8PNMkVe+qNN5lp4qko+p7Xsz1yR
4+2K/R1rp2KCt67OuaKDPYUWR3MH1X7zp0qhDgD99mVgQvoiofpyXRX47daos18i
NbzrzMNb+vSwBZkD5wHSdxGfBsTlL2HqpacOOa+BTl+AXmpMrWJLWdifK1BhctHU
S3e3bRIyS00LmcTfnQZDJ0tP7Z8NwJMIZUtMDxe/V7PxEnuNsyUSAM4BLt2FzV13
WhnmCScMiwbwp6BtkjHj/kzGxoLzJAWllOLcBLCrrdPkBOe3MGzIRrCRmvrWfDVJ
dvn2wzUtOFkzahnCtWMsakqfYAcBk1xIXNa+oOgg7q5OdcYsLgMxUielXlx/yI5d
qUjCiLqf+agSqnB0VviyZ5hDCpjHRpNDTzVgqZFNGlHY4NreG8cOEAcQzSr2otpS
q+piUEiF6v6wJy+mZAEW2/kCx1wb4/OA8n1fUCE+ns5KRihnMBqXC0dAwze/mfSG
9PV/qHZL/gSneNUkcXgztygsaPiIzYD9fR1jzdeM/S5u2+u01feRGM2c486kdK/V
/GxU7zgq+4Zs5tRmGOoqWdmgjXm4J8y0BAhU7ZcC3ljib8jjhuMw51UYl8a3FF1t
Ef//pwWPBjCot4YfLMyK+clhwpAQAMWBlDjIDi0LTUAGSfRoN+ShCqXGKcrOp7NF
DWaxJMH9IHBfGWtJfUoZjScC4VTjPAVuoobkk+Sp71OqvXt8hzBYpjSy5qZYxxv/
gapv67fUByN7gIVoxbOoN5ZnambuQcW15jle8C2xIHFMd47ZhUKtZnqzazMh3xCA
hxosNJILrqqI41Se980o7OyFiccipcDFM1b9H+pkcx6dEjqLIzaAKMdYeex68vZY
P+1OwJ3wpuoad6buam/YzApY/iYJX0yBeIXgmn5yJaV0IbkY1W7//EjzMpR/X9Xi
hXcMjrdbpP2MNUDDEK7oJcgqjAfIGb7zlQkdwFlUYfQDWMhhqxSsCZOzIjbsSPh6
uX5ZTyyA+452Ezmk0AG2aDd89Vrz+i9Tm2Q87kowjjV2eKVLd6erdUHt7jY75N/o
ztHI9e/qyI4nx7Yci3wd9oJOMR732yqdI0Ku1huTURHW7KzyIZ7xm+D+jK3PUSKU
EHu9/HXoOGUfYN4o0i9dirZC2eiQ1ibc/m5ShX7s1b9iesiZlUm0xttdK3tH6Vdz
b/ZCEur5mNIsifPLzYfvH98frNITmMrZgwJKcDOXL0L+rJHDDg3RAUtosrg4GchN
3zHM2lTH1qiJj+7Ck1Wlg76U3ekFNhD/2bXA37R7AWanOSjM9xKL+IDtMPzdhpJr
J6e9KplmFKCbsRU84Eqst0a6iSq4tWkNEExPBhFocMkwFAmQxp1YeOtlcHcGVsb0
aL0EiU0HgdULWEu28tN8qyriWNXLT2TapnrmGuyH0Lhr23/S0PRnTXVxNo2We4Rw
8EDfSMdv163CS9O6YB6CzPTnJNf2FK+CAXYSqu0c5m/Jaf1d/vbbEvGr1lhDZt7y
CEzNCEX3H7loKCQdDlC/Ez4FFXeBwc/n8imy0kVYv4WsK+QI+RGQ7Knq0G173018
HLqRfrX0j4lxTW7qbE//54VH9JGjqBb+9fcZGPMJDLlAR/MS3JIqIRCF4aCdLzTT
A6tY06jIp9lpUrHgaSsBLCjlab1Mwh/vOcoJqSwx8xinibdrU+WSJ5C5EuTmG5VZ
vIVzlwxa8EPlWtENxESoliIPmTiLmTSwDQNAzcSDkDMMIt7ZBfV6JyGSYzDW6a0h
OMBl8UuNsqT3teWwT3Ah93ssGRnZjWDSTH9OCg0VRkDenuOgqmlYmxyjMcWbXasw
7K96cYqojhdQpDpWC92FMUtNxs4KpVRiQjFAhrH7Yr7t9kkyAcY584VwlN+u1qOA
XW5dKwT8czFZiTTklPthgj+mnSq1L5BJSqP00jtOF7fW6MldFwIosqodMm9HAbmg
L6pHupIMHAcWRI9IZ++mdIvyea2RwrvfeQLUNzK12Z1AbRBqQIZ5NGvhZGCYxbac
TFqpXsuXSUtJBDbuWSHJl+Xj51gMOZvuQrwTFgku7NsM8dQYyt8iuez9w2ipJ8xj
uPZLexmNElc8LIgHXkFurmEyuHs/Bw94sH5gfjwmkaqTuZ4OJ4NF5L4BPGmYFhG6
KTstKkuC3Tx8J66S3ze0n8tTJYbHJBcQg9ETcOz+wAgzcX/KVKRdnEZaSufiwOHz
A+7X2PN6S4NfyNHJ9qzyelO3Zi7Y3KgtC54e6YRgOGhSM72QyXrK5WAQzHs8YNwT
YJxgiMCUN8S8Uon4CgDn/HUQpdOQE2EnynObKB1DnNuKNdgU2edovPvdvX6xIJqm
7T7kusMn3IpBrxUI4mBqHzGeYb+4G2cEkXqbXSpQznQSjDCivEsNeJfqj5mbJv7r
a4rKQZDCKCl5iW/XR5J9DJlW4j/fOo5xcCX3kIs28roja9A34EAj1TP4/CLgjg65
ZpnZtjUzvw0UQ4ncs1B+qO+DAOltSDt2cOY6FfS/AsvBtKXsfhCUKrcLiC6Q50Bo
CLPJ86NiYSw0NpgHNm8eLqoBlKG8EQB8d7gf+gGf58n7DyhCsanjQDbjl3poeowy
8Wqgb0E9ch/9hIsXoeCBP2CAKQd91yDNpB0t2hZfEJaaKb65TjB4KQAVTzDCfPpv
jaGZLeP2z7woBwSD+L0Ly5Wd7lSD89yLRa7kghL7lk+pLaFXrtwxKHm30fptO1oc
m2LFz4GNEtc7t8ri51pdxokhWK43yfNPSV1VysDTqb/DWkxfRJH5H5AoNtCuYoyM
5m4i93Dnxp3rJYAdpaUGcsuNVTNWf3e35DeEDNhLztf0kIeGMYwCeGw0lFspWuoD
XAgjksAf4YCkMPeOvKi3a6ah5i1NqN4CyxBocxEQ/UIk0zIjOW6l60VETJGgmArK
hhDxPbe2ombMhy/HWkGlbXEMNNIvmIsYv6fXqIUUkO29uD00SSL3tKoWCAfhHiRL
qgoJvRnbOgjkF0Jxn/za/AlIcZOjFcD7uVBHlZ2dmdxxgXNb5+QcLyYLgSFE+y0p
8JFB3raKjGQYG6NOa+fvKnovtMFx7ArHFEd30vN4yVg/rREhkxAyZ/FpOp9FJnDh
7UCdYHHQKCfbyszWNR7lY+YRz0sdFEwhDTADX8NuSVYIva9vPxmGMpMZe7dn1VWi
sa8b2Cw5ooNtOLjF/xcwqqmBdOp5v0PgE0sCYcz6lufwpaJi9H0pr4JbE8K0fjI8
X24QbaiC8sOhyT7uw6CzxD/QZEzB5hBDK+W/Su2JyCvty3Jdr78+CkHsrM+YPLaw
gzCmCJQhiqKi4ZvEDYsj3SnTszdN4T89/7rrAZTlXfwNKFAFdEbTBBB6W/wNLAV0
klvRLOvpHFRSEgv6wffbxVEK3YaKneKJhO+HGOENkpKoopJ08aCTnSd8QbeniZ0C
GyyTk9IHVkcjHoira+AZTduMfAQxA7OUd5wh+dskLFRGuQbG9ngvp6io9SFSSW8R
rwma5h24RtogkO7qEV/2WC61YqS3hzkxThH4uEHfHXq6gQ5X3jCIsI8gLxzBFDZ6
qaVe7caXQpK5mZRBxtQk1oDG7732DvbE2P67gwZL72ki8HLHxUWy86wn9SPVP+mP
05+SzDBlVjadCrYsjzSaue3eaYU/CnsuJNdOOCHP4fsldczBxGRDN/T6GFuzHQhi
nUhd0z1W52N2fMbDzKYENqLquY28GfeQCb40HRlbpBNhQ4Yp7tr2pSfQNrFp7i+h
Zvez4MLtux+S6Se39Ju+DxFn1zPqM2H33fhRXzQo4CvqdCyY0hhQlOZCoJT7tH6f
YoLQ6pnGUIHgKUCqPEz7buUgZavYoqGHde9Bmomev6QAaMeHQwC5zsQsnElAp86n
fgP9/bdWfNDbkHnosqbuRhNCEUOIqefph0joLrOEgvhR96jwws/ce4q6LBWuDKBU
GB7ByjXRDvkPTuppCauGNOKWq/5+fZ4XPcWaL5LIIRGDJN/9KtHBIEmH4O2zts/K
CqSfwnxEsRiirzmYJJ7NAQR/hl50M5oWUKqAtFA1tS52zTWbJiPpcczDh6zJu59X
5yY6XgxnxihDie/3YDdCl+Z/ZuksMc1yQoqQWqNfcGmsMvTy9l4LORSmx39PeR+b
TKCO0pTDWTdVW+28dswBInDXH4TYjCoLhMcnqFJwdTbPhiGi/u5L9GtYKyCymjBe
AbpCXdmGAA055KdpLwXlMb4LFp6juanLS3OtUPidTpnXlU1r7cmOnQf3b76mtYPt
8KGAhKgCiXMiIks9YWNnPK/hsNUwgsa8qnOytZKWYqjiiG0NZa0P8a1DxWI6g1LP
dbMW4tVdmvzdIbGy7Zgx0bXsx3HMIPERmMK6DexM1hPAOvh4Q47khQRoDn2hFobz
qsBrFNZsEaxExeJ+iCHaw+2wUITO5uDejA0CXKc0FCYl76/voBNZTJ1KppW7sH7z
fQsa8TnnHdVfSqI6xdEdJ9FKitsrGyrXQYasVaAuqsj8F+6dCH/jSWZvzTRiqOD7
eeGYlL6cCcweQoRx7gDOrQvaIkYesEpcU2NAzPCwoGjosENLAMsGZkKQQQEzWF13
qLGkWTFS9RiBcYjSfrEUE0ED04nzPcpJV3sZYBYIBYUgHoU2xbbu1sHELqJojoTp
sKJTzdzt5LO20jHdRJ33UTX1CH1C/NMgBaEQDS2sfZLX7vRHwjhOz28avUGFllip
ca/xB99TeaxEF4Wx2FAIK8UdrUyZz5uEksHjiEInvxesQRAprnv1yeRbJDF/yujm
PqKhxGiu1Y7l4Vi0xQGJx5Pll+ZsFVzMxvgytEndg90WIZXBrWRA7OgnNAVWqedI
YKOjajyHqXHSW8knl6YIYZeXKeZY8ElBewseriUWP30VKwT0IShQDQ6xutlyJgHl
sS8M4HLR4RURAyKWbsGHjdeoya4ncZnUq3WD/qxbtbT/bx20EmTZCcFzRNwzr91C
hoXG/4SOkE8lZSnTnaskwF13FqJoW5fyEw5EZGU51lw0aeNUNscpos25T4ZihBbx
usdo2RjGr/Hf4uDaZCyT6Y5m3pzRe0mDVCpQHd95fvyqTsPCYI0DN9AVK0Dx1YWl
W2YxRvVRJIrFqxLdahSayw2rziXz52ZAHr/WNNsaJ5RC4Px7xHBObB63G8Vp9gGj
k6R9tkkwFOHUO1ReXNRozFBFafhMFbPr5T9Nkhx32HszxRsoX9wteInohsL+2Haa
UxOjAIE2i71h46A9hjJEnic1lnvY+EGGJYhGZtYzdICcnrPx7gSY9u90rfOgHOZ0
a3tkDXOd6YdMqH0/nz2zj8tHFNapWBOoKdtojXbUxMdcfDmN3dmRUZuMkVpTmfKj
pvIbv4x4Zh7lCYvDOs2MFQmWqhDebwUrqXA5zbHF/v1X1j05gw/LR2oGnS+zICTf
HjUPkkIYLxMZ0k66XWU6DuFWcXeGVXe+lfPKRy5NZDvDAvTDoOYjFvvbNbLTJ8Se
PjO54pcyj6g9oRiIC/ZRYu/gLC80PT3St3CQN35aN3E6jh6patnIuja/ymdayQIH
zwJL5NxqCfQo4LlGRx2wU2/aEEb/BwlBWEmoQ6i6lUAKbXPCyE6Ic/s6qlnjyHM6
n0s5kOJnomHVikMTnHTzYLdqlGeYdSvYkf73M7vyOmurMJyMdi/JTUyCexVQumyL
GL02dUXgx7aIjOUJ8RKryDJw4IwwWTRK55Lvyqcb1U8obvCTva1Wk0xtRR7ggPFQ
ZKLZlTmZ3tob8RW9xbRbPUw19wtUx/6EroCjfKrQCaRBsY21fP4nyDVqpKPBZqb2
ytzp/nScNFLgYJwIaUIHo0EEpJ4Hkdu1GOpKDhUSpYvjKQB4WhBaJxHR/+2naLWQ
YrF6WFbXTzGQKej+zwzS6n+4AufFdOR+cj23TYndYBA3NhQ5KBaQPwr93T7meHWG
VP7BL0EPV++H8z5ZpyrViL1FwnLRMikdra29n4bqNWizz67Rx+WiIt8WlWM0t/6h
P7RVZVGeskhFn/6kSc2n4qNKIThwzhY9ffC1HYIY9zmPDRcToLRITzzAXoVI4dhz
E/SFtZ1obFGWM4gf9BlGPX8FCFw08/8RUsURiZLxDDuYGHIhy1lAOmM4tlLmlbUt
aMqHHR2n1FtCSO2p7cK1U9D5Q7h4PPgCRWzUZC6Z/+E6f+Btl/0jrpz/HtnSWeah
7O7kaR3n2MYuXag7mwHIT8xhFlbewJKA50kvvvcvFdCDj/zP+UAg/NM2eHH9pGrt
x+w8UTfoonc94Ql8+oq2LVxsDexYiH8rameEtl7iU0jD8tobwPH5GejW6DJZTUYz
qaWMbCNeLcMLQBDrEVxy2/+LqNay6qfYAUNhbkMwL0d/kktFqSiqrltdGZDu3OWo
7OT1dpkc7WPhyVW7ONz7KchgtynYuyasV3SJOevetoHGtnN1+vr6qQdgCrDCkxb5
sZMajv2SMIWS20gCamz64uC90i9tK/gEtTjCUaPxhcyXdwPwGbYwnEEfVXpbiaqT
WV8+/RJ2VZEACrSRfCTeVQiuDvqFxNH8kNgDTKq9GDEhi0PMj+OxPkWGGAqIkR4Y
sx3jJtZ2UUJF86iO3jVjyLEEG6O/IKD3rP/kNP39gZ6zSlW3tsv3Mq7jZMohGM/T
hgU5yvWfD7de0Z+hCeoAA+SMsOJfWnbGsc/LPje1uyNdxedXx6N7tFBhQ0kY46/q
s7r0GzmaShi9s5T7LKzuvhKw+B8uGqHEyPr0Vw3rn2qNA/3fTE1Em8/najVA4FBm
ZaTJHXTj8JhATlv6omnjjK2Jdy9muzv5M/rzO/0Expa67PrJIcvDBne4Wqq5aDkf
H6rkXFYWlTKJZoz3Mo0vDc6Qe1RfvMo0Aw4Hv2eZzq4ZHqBFWNokj78HqiPNH1Ax
knm/Kc+9OB/sLDoP5jo+Os+cmEr6sf1JqUR0SShrI0na9CTfX38ea0o/xRoYizdO
hOb/jC178TjjiJz1EkU29HEIbewohRCSFnlPX4U1cdJHU8Zxlmf1FYpBLwzaJwSq
rvic0juDjfNmdfoz6zcTSeyAJv8BBA3v6BGRTj5e0WwmhxiLzYhpOqZiKQ1rSozy
BOdfUDptNUWqcpC82iSa3f2stjjcnoC3i9PnzIcs+RZ/alsKccDXYEFw7sHmonq0
cdv8mgz05x0P/5gTeBBObpbzp/aaFI/ulDAKZ2vRK/2LvcXx8EqonY+4NM8Hs/zj
2U7S3wNWRWprHzE9owdpeqJPvrIW0YivCWGr+bhTDHLxTfZKSDuAbd/28xyng8uK
AfKsrs3bA7iX5jFWWEVSgAz3zHRjHDVQwU5eiWdR+pxGiZhaJ3aZOIX3whiOzzBC
2lTc9T/O5pZgme2l7q51+tcG/oW/7nXwwfJ3lasgj87707Gbna3IIKWg/7KdAzkQ
suOtCPYDfFsuilmelgjRa1qH0ecupQQVX68RJsb40cuYKZDT7Ly/FHUpKggJYex8
grY/wkss4UjDh4jJ9PieR2l+ptp9+aovbRF1ottVLbjoPTWplASyx/3aigjZ4OXI
ZhmLcUOvSgmm57p2edVxD3bHrmyCvLzPyhPOqbsNa+WV9o7On0N6h+7lmLUqHFCy
Xbl/BjTkpUFDXXO+hPxqZWN5orhiOjal9B021pT2tRaWvRHTieaZpf1fVicUN7Ez
7/Xw4FiKuqBa4lMG9sMPbCQEgaiJ2gS87X/zp6Oz4ktI7+BA9cv6DYuUQbfmpuBw
dQkilrcKiqOPkakPmGyMigRjEO9NQkOy5efw/YJqXshEhdBkYQJTLcA1ENdn1pHW
bRuAWvLqyFLsDmKd/lUycHNZCK2+ZN4eplclNfG686m6QjSYY1mGyLCGaRTK/jE5
cCHFrV7UTvJCTas9ROof1mxgEdHmqKowG4AOXdiYvGY1ax0bctQgsMNy+n0AcJ1o
R/w4IbyCtN77rDBxCC7IbQrnjmDCV0ESYA8Rb/DqsNsPjoGNAUW73EUvuqqch11X
aA/OxH02UNW24vNo1yy9BwnNqPc6rw4atnslPMd7ZvSgaeIMW7+jo0kiXOBUhprd
gr9ummdGmophI/Fv+MiBA7njHoFQh/yctpz6wM0A5kC2cdyYoxk39W6smsq5tPLZ
XZDioqks3Wap5+WhHOMmETzpdrLp7kDCSRBPiyj9E0z0LuR/MjDVpu+nGndI/RE/
Yt7KgHDgXAa+XU4OAMQBHjCWuF4KpVACu6MV+qlPNNUMzsTsp4QbUzoiit6Hq84P
STyJfD8gA9qWDa/cGjwyfG7uiZdwqtfwTIRYuv9/46QlaWShi8zxmdJd3XHCpZ+q
0hZk/hSY6r0sk1LW55ec/PVF4vVoK0yUcigiYMxNF/AIsBwcCZyeWN8GImax2AHO
+HvWBQSuZy5lV5AmJ8PkVhpj1bLmCbYbN+FcJ0zzSrBW0Wnw054PR5IVtbqKJlr+
pBbLcN14901QJU9lBVrIbFqEMo8TPOwskTXTXXweZwmJzlwlp0KhC3uZVUafW1HB
ynq2p3zqwXbQVw7GibUFFi6J6tCbZ8a+ZCpIY9y1HmBRh8IMCSsboZfiSzFnYK9j
69P836takByWuo3GePWLNMqNgmEB3rmIX7Ly9E2GRTZgdGwAUAlfGc9cDz6EPdBw
BcK22cIAeyx6jgwONhAcDxRnV1rEvIWN4jkKIVEkJlJng1Xx331rWtDNLqjRPYaR
Mzl8kT8M53mDjJp/BxUoc7LSWFLbJ0sdSzF7ERO5aqE36enR3vi8XOpNuOQOS1gj
oI+ypATuTJkxb/jNkLNxopTNSU+IOq859H6EQ8sRVTw9yzQ5lGSOItY7dF4rZa7H
5Ut7VM8OCNKsBHliouqPfULBb9gPRteLH+eabOygdljeBN88dks4mjfDycC+GXc+
GSkHY8JGklwaybGdI5nGrNpG+vPRDUD8ztqJc1N7f9OXeAVSmCg4qwcdOYKgWgTR
3grAKRJLtDZuPKAxSuL98gJVuIDivEsrmuqdD6eOQD1Hdd00mNsGNpoOZRc5xfJI
HlPZ4G3LE3u2HZigqaiR4X5NK/qbeALydqtGK6FbMgT8vToZe6yv8A6alxfD0Oix
xngBu3yELWCPLiFxiDAtP/GYwyh+e77QZJt+fmaxVLuqnmc5ALLFTfI6wXSQucld
KR2bxvj0d2NGdtoxpDs6Mw==
`pragma protect end_protected
