// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
N3vuFnRf0EbhDTG2WooUnvpY0L9K471Za9TYJfcdQf+TMcn/UYHRSnUl0Y2sySJO
WRj2ulGO3npfQQ+oUa/1pwcRwl29w52xO65x6lsy0gfcmYGIO9Hhu2ViamYFRdB4
PZ+WJWCSqG7z0d445TJztV1M7jz+gKsDx95HUXqddKI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6864)
eiUojBomGT6P1ODBxW2cMBlazBKKkNkyFl+6gZu4enRSwpcGqxINPf62ubyUjLU7
3FSftG+cFiefQx4vFzPPk91ZNA1d+N8ksUIFaXFxPxBKHV290xQa1fNOF/HJBiRE
C2ICzihlciYB489SyInNxv1wyqqV95XAokbV3LYh39w0ztNFKkZVC3K1QbTTZjqk
XsNDOvsDCMUYz6HJmTttymVtZ+XKZ3TC2QreWfdlL2zgVBa8kGvzryacDXybxhC4
/hVomX7vSSgdiozF/rn1LaBaskmbIVzXu9VofECevwQCXU9ZSvlTw/hQWvAu7zkV
NFM7G8r8Z2GAWHg9PtwqYz6fOwy3lG2iGivJa6uyOiLDreQ0yAQ8O6xzFhpmTe50
NqGhOE0i/Zs1gufbBkJjs2uL7jmdrOahfi5tpWpxkVLllCKbpBl3o2xCoIjOafJH
1w8oHv1zfhXjOotl6Y/put0VK7R12kewbWfsK8xeg5Se1x4HhYvk0x+XIRMZFyzK
wt9EBffXldSjJVUi3+TcCpdaS5SKzQMoR0HE2D3XcBzNN2wzwoj3iYfno7vocT9D
gREUX9657hgvM93VlCf8jf9I6DE4pKuIlcF7Cje8CqRRn9l5fUvoHDMt+i2DeW6g
r7GZ8vvygm8MjaVZrAIsbgYtd39pWtzxptOsXSzeKXpI9VJ0skFl7g7UZ2q+naGR
DlpPmxwbGAiA+3tiTg+dSF5ePL4u1QFUOxOVbhPHbYb8qNp+NNLYrlzi60X5PaO9
WQnjeRIeZQ9AlzghUpaIeYSyXo7SVr0sXuOG7vjRq2UwgW0ciLOFMxrt4fLnngmt
qczw2lukBr/RNO9HfTEjSScqAkjBxrES6e8hd63W1EAPALhoPHQa2103fPx0sCdV
B2LMMQBRs1Mjfpcbsb027VjEpxjEU0So2XpxTb3e2o9aSAhHKpKcPbCY2rSTs7/i
OYNgvFMlTRsU6gAY6yxyszARTTVP/R9dck60b/J9OS5IqLIVTBWZyoEr1UYewG/V
sXA7ZRPeTYmvXPKPphCO1H7rsoTB9Ez5u6yesnjHtgXLolM+I4q1RgdpmR3GAbwu
K5fGyxIg5Xn59q7c1O1dEkPSJ3QQf7b7gTDOME+/10Fu6J1h03B9pEcGiCETGB9Y
9rDwYvlEfNbwWIQi8rPp8sXqc5nokJRHqsLHOeTIoKa8yZatbMol/vxI5QKHRv5G
o6pJGDdd4DGIr1iaMCjLxEqxBMoQ/CC44ZHpAtIt/1NhRFQQAA6Ty4u9GH7W2Qb4
Xxwv4fR70ldTwSVhUApehYMFKP4fhwRTGurKLGTMuAw7tu3e2C1MkrpsoaFsrIXb
msGOPBZh9/xaL/pYW1KV4Kx//VGVH1Ac4Kue6vo6u6K5dmyIFDDcbuQRVQ8tfu3w
m/8onXUkxLkzonxxDnjY5O4QHyD6pSYxLqv2mEluIEQ2iMo7KdZ20/y+cEwEsYif
MJJ6AZtAbyqluUGja4Xj9yY2HzGOHDlmffChhVXEvxYlMACF2tEQlrtj3H7uVOQx
vNJUz/S5X6nv3zvcaxFxTy/UBJZAP0yfsxJvqb7meQXFGFuilTkaiH8vxvloeM6Q
d5q7+CicMTB1Swul/kpwlITAAYqPf50RC9wpW6pt7D7vvuc32tLTLbEtXDuFXIXk
d7YKKngmVFXRtd3hlUrdqpCprXPFVgvsjCnaTIbtybEBSgHCvO3s4g1/g1/TWuyL
ZSqEoB/F8zvBKEqnd8vQUmPe4CuzlPXoz1ofGhRH/7r4pNg1kOvTyQBCeBzj5tDs
d7QqtBjnKr2HDh5W/slcp4ux9CJA+mljtG0D9U023RUBjvnRVH1d3ug0qe2dw5Tj
SuwbqD6lbJfL9latfDnA8sHWqaj3Y0UZwgYg7ZXxaFNZfarGwdo49M4eOl2BPiRX
2Zuw5LNTvXSC2MFOsZz6nficeIX19pCgQiEJmDMhiY1+H4ID720evTABb2EQbM3A
LL5XM73GZ+WQP8Yl0JD/p+pYhG462kzYte1DXzD7tq/4UdjQ7y5bxMqcm9VEP8SO
4W1D5ObfNJ/K93ySYZyb02obQGkt6UYRdYWvzHsEQNhrQgIk4MwzmfLU8NqaPpBO
GXg/3iSh93qSkLryuhVShgjlpzqkr87FOYNsiVobqZNGp1q/n2c6sEVMAkmAEoBu
YsyWwASbrSeQ46JgP1s1FhJQ+lZemgYWNsnCJk/0YjFAuP/gI3LULcfCEX+rdDaw
M8kEEHUZ0ekgVFiBrtEYVz5PcdunlYJqTOmHxmPqoYBlcxH+oIqSiMJkNcewy1OI
j/n+3cP44YIe1tlUeNP//GswjY+Pib+ZM0f5KfsIIPMF3WnYLeDfnTqT4NfZJwLv
ZLnLAuzNg8tfIZKuDS1qOXjD+Ngngqb7myT8Tq+CxDhViaCi60htwNeZYHDNidrj
GTSY9c+ruGgClwl55bJdqVCuHhkZcJCRKMEFyBSLMtjtH4Pj+XbubyzAMOgsA8ct
l30I7R+C1Gsw9eie3ILJMWBAzs6S1y+P1Nf+qLYGa69XlerXUjssskbVAWxZdzoS
T8NCQiRiGcdvy/ttqN2H4W3h7fnA96KnHSLIzCFRupXq8dkiGvAzMsTN7S8Xof1O
C3pV2s07rwqmKHXVG7cfDLx24F8IUH3sp4hTGk0hQDgiRqKqpKYUAjs4l9Q0ASGI
kKw/8+fUG1/vnNyzOKSIvnDLzacrhoPaVHK/flSDMH3iobGza7v1np5i7tDMtyWE
mwm7XqocKu5pqotbSlFjeavzWH/EUbewLuTNx5VGxXYMLfFjaX6tYcuPUw/hSOlo
yJGP/Ex8CjIL8uQNkeQPSM/uHJnkBKlUp/Pm4Rt8Ma0ntwzF5hv6DZgNFK2CGOS0
LiSHqV8Rd7cdeZkCngJChJMkU2FHkFHTWcOXkFYuv48auLDYTCM9GT4xSddhEJxR
z3UcvGH6qoRucq/G2Nw7NdZ1CBJqTUi3F7NdSipSBVO3ASZMKoNngPz9x2CmmajF
uPj9yxdkreGE+JQu2uotKmMYCWb7cq8U4qJ90W9JVHQjIoD4pFlkpCon5fBdigLs
Z05h8pnlL0TizS4w2qnZTjY0FOwjCZ5Nu6Qlhrmc/z7KbYGBHiPjNFVHZJtE+UKb
EN867YpkPOEz+shi5tutxlQeybd9BzqByxCvBUGlGC4AVumGYs8oJvU2eqP7YL1z
6dk8vKZCaM+ZvzYiH65Ifh0O/7X8Fnoj7dwJ3SCKSEFlJ4Qwsl8lQuhjQr0jxmAz
7Y+6zs3WZmsiUUGX44eW4MT/cdhJBm3wjlqZBxKb5sJXw996XJAniok2qaqRKi7a
CQ5XmYtAVD11PeBvusdDfzUYxlvt3v4wraJ/sOuUN8gtstpYCTin/8gjiOlyXKDP
6JmQVyp14dzAXEG4uaPjabMpcJxKMCRNLn3qJOh3ufk+chQjkNWk6uG2i2jZSHot
27SKI4OO/4dXZ6Hbp80PM1bcefzSZnMbOA3iuGOnP6HLfIJhbrhLxJ/9zdwZJwip
Yf7qEdypMtKYHuKZFX4Os9n/nQzl9AVkoIKBbjYMl/ZK/zJ2yBCGq5J4stBX57jt
yacM0kGOVdiHa0hbWmIy7o43ahqUbdXv4KnPS5EvV5lk1jVtmXurCHGgLlmF3w6s
vya+DhA+Ps/oQgbAamXFSloVJBlCwU7zT5yZxsg3vXM1XzsbKNMPkqnQLLnMrEg+
joJIv/FXhoxLExesSfmDX5pzRDpr7y3AzGXQcnj6Se1r9jOg6HP8Y83dXvd+UP4r
G4a6ek03Vs87SB0eDUO6MuhB29GJfgO1QVWMHbYA3FIYYqw8R8MYmFLiI0r/Jvi6
s5QxIKQD6V4mtjlB95NShaBoiNcw1Ga3LAQPONZMWPZ/AlAfu+UouMfLvRXIxsbx
48l/7QmB45GAferi+IEltZHJKSJ+bd0PpAKo0nSnZMDBLjkHmUPulXKXP9tDKpwE
OvFyOm43avwIMIfCNdvl3cKu+gWWlRmdOco6HxcLk8E0yNUaArWablfdyGIF2pTg
OLSHFHnu7MujyfW+8O0PcdKAdIM3yHBUuiorVhIjXlokgeOt9hGguTccjtYcNgnQ
i2PW3Ac02mvcGfdI4RUQRZfNaE0QlW43OBzE0HDMQ88Sj+XTCebzbzXp04gXPc3W
ktxzw2QrtVrI2l9r4nABNTyxwrMOV4PoMjvVg7I0k0me2kKAO1rtn/558OTExPJv
X+rzKOWhzh5lxBf0OElIh/37WqTRhF8NfzFL6OO+Jw7vXgZPkWlwVfadSHuxoFDx
WoDk+FEZdkSpUxGOuXI9lvxXp7sclvJf/pGw1kdr/diifvCZKPmG/JickRdXNyyo
pArh9HXAvv8opPHhQIX9nZCPsn1vRXm/kbqur55EhWHOUJvAKbADlM6CnaU6rB7X
UQPHd6zK9LUuPrlM0Xo3jUKvzX+gfYVKm6ZyVEzCLm1Zcb1hlSNoydm7K85uADse
Ny0IBMWgGwidD6+Uh6nciP7Gp+5e5PLVzRGhrWMp5EtkBa1YZ9Gos+f4k2czPVhl
6TRUpT4su6SMRFKtuuX9AMATd3istZ7ew7cdJAjNITJ/yL7XTo94rNR+lRR0lPwo
Tek1rFLHfGwWsI4LTZlJgs7mcO2IACsBAfSa4Wg5b5AFgQfEnMLxdJou3vZCCAi5
Rfh3Stlyu6Cvlem2ml+CnFIU+hhwVn62jUe5Nr3Nppgl9knBEk+7cabxfjRdPFT4
i0T5lW5wEeD+D6MYoSy8XSaCpL/D6oAwi4EdkQ6ns90n2ZaI+Ng/4/cgO5DTE/LP
ui3MziQr6xzXK3devbZEUE8MAON2oiSSGTGtLFzaH7YFbZGcohlGlM3v6TwEoUgs
U1DDsyvcL9W4jw7n3fj+16ZBtDf9odfeqK4+j4jZxgmICU2Jj7RKXp9cUFMyyAJA
BgoPz23vJHXta5AQ4Q4teLjXgYCv783ypYb2lwupkIKVmggYvG5sbJahBSAYXARm
Jt6M/hGd8gERbKJgyAryucoS38J6T5j0ZIlBjijs3bDHoBESBp7uJJikB04WCi3f
r6DtqaqD9GEfOmUDJKJqno9IgmMhMB0gVxl1ZuR2J3j+i8HiawW7//b+qAsv3iop
L7Yz+jlmj7RY4WWn1DLUFY0czPte4vlpKX7itvOU24CdkFC9Y0emq7RAPfN4AzgV
pr/LJcoHuRYluZOCLjAMTadYOH5teBn9GcXiuKj7kHwN6ufhr56ST4zV7bnRpkmh
U3CQoJNGMexE5nSkaiyJHol22hUU9M3jKxihWD7JFiV58nO24pG1f73dkdCXpsB6
S9mb2lXTpyDPkkw33EJp/bdzOPqlw23JyUXp1dkaxhVAX7x9+U7PFY/q++KK6sAo
oYmlOSWzFhXC3k3q2O+CetL3DcDeglLlATTkYq3skAYxYbMWVRblo0tHhBa+mKRR
WXme3LewH8BTsn8Npq6rCVWOP0lyA1Nm0x1Cnaa67uULHh0CC+61Z375mcoDpJC0
jzS455T8PZ1/oKRJ+SSlJjz9j6hICZbwfWYCvWVY3l9zxayOt2peRaNRx+zqQrm1
jbEZAHLrEiR0AFcXp7U8vGeldNpz9yWd3LmkTejggrH2zT+dElxIoTD4+cqJTVtu
m0ZR4+75AQi7TSJpn7b/jDtVsjdm4sae9A/OV0glSzTkMfVsnYO+z+vpiB4udumB
CbtpKVpdNo4lQWFbt4MJI6E+dkpDbEgLksqrlOUSs8qkYtxMRhTTJ0BwilEb/CXB
aTKXZKJcVPvAHtzCC4Dg75eNqiDCFqWszT+/lw5t30dHcU2gHK8wAWaTC41z7E36
OfzfZlviAxHjfhcFFuDSANvFAKEyBMPlU8B0GAT4mSt6bjhXH3ubvPiU7eplwx97
y1YFW2nqwOSKH7MNveCrJoefKu/f59ZDu7eO6yoyzxZ5BOVLLt+a3EgF+3Me8jxV
KgYC8M+PG/ASJP0Xi81XoV7QKBlpgrrGWeN/zsZ4b2wtIMlfJ6Z2tuZzMJnPLiOo
zIvuTtkVGI9RRuYdqkqQ4WtMMmjL8nx2mXflgOKX/s4NdEySVDOTFhSDvbH7Cdfs
5z1AcGFeMmm63ambMTqCwHx2zvllf9SY5vwRBd8fP2CVRxJbb7bynR8OjnfskxBa
zvMVhBVH8Y/BwAcdJDCNk7elhfHay3LxxzPIz4Tehqe0lqQNLwa7Erxt7H5o+w40
PJCqXc6D/P9dRDtTofMhULvEcdVklmjCAStbs/puf/619JcazEMoppiTZoEDFxD4
opqpyL6BWvcxCLuRUrxl+JHfCYuQ/KJeCOUg2w2jDxw81w1YUVhuOMDgz3BIqsK2
/HPzR7f+6arUqm+RPoKgX0xqeAUXslldNY9cU9sbZhytvq6lnrZwqQksBsmPcpQn
gyMW89U38Qxh0VgDCLNbSwfEUl5+j3H3o48GaIcGQHgniFlVY+wJrwEz2enIyiun
V5lyyehQj/pHKTz9QBd8xA9W/o/LHv5fOhsLboyfAJlESCelqvHdqtcxh9DnVZE6
WdLg5IYNOO0osFTMrDY3zmgyKnl28c4ICR5hcToVaU++0SwOzl3AXhvEA1cra6pI
VrRU7gGS73EsFAgROmgSnzGucglDbT5QRL0YGeFjMdDtDnpfEJCTFFWxQDyRZzKg
82m3h92fEqvlHegKh7s7YL8Rfug3oNhxbG+YHpMxj0nOlFE6KEHhNHSFIP9pAfyg
V/2A5fteZVnU2cVp+FfIbgNm/LMRbOLWPaYWzitQAwjm2MTiRe9iGyNzo0uNrmjj
gv7fF98yOQBMvowtxI4fw3sjQSbWS8evkgmVBesq+sYNpQYORzCyOwefVFsQIH3i
JGxJsFGLrAt81oo9V08+BFbssRTqImXdBVRbXB+CZuLw3ejGC07QnppW+Jg4LmX8
41kudOWbR8xG/se5pa4VHigiaJ8//s6zjvlnKVInxGSxF/EiQyFaZcDdpyocsEJi
xs6iMo/b5DNf62QSerNY9XeMdo/YiVmZ12l7w8Ae9SwK+P7pu3NB2sFyf9a5eEZi
dzAihSYFMy+Zfay4uV1uwsaOKCPz6AvRpo3OwhL/57IQ/k8pQXMQ8W3O3iUlow4w
pKcKqScWDq8tRduoo3+oA/QV+g+BC9OM7Mpg5pXF7vAQP+oIjBgHkHpsNnM6LSmZ
ZHnlHwOE5pke30+DrKhoIAyFN9EwMKpSklZ4x3SC0iOStUdHypYntMDX+sskm7lT
cb4E2BlgodXwISMqLtaW4kYM5erOTcKDrEg+zg9ukh6rrqxXHTyJ8Bg5RlpwYZ9f
Trxgrfd7H8FHK1g/Yw8wtkQQQICAx8r9STcYy2Yxw7EDRH3FwbINZ3Qtpi6GYdsT
OG82vu87tteYgcw17bTubG0eUbT1j9L516YL9t5Rbn7hwpWw+n491skXJTtuIanO
YXAsikQdUDuT//k+UojWudLxb/j96De5V7DEs1mW/OnBM+9WAHP9tDFUVniqzGqq
NSdugWVwd6mvjlIZb9cR1HmJl7+QZx2Xo/c7r52qgOKnCeT9BxV6L+r0HwAURkN2
g34qRj/qCtwlFVns30FnUBBE/0hp3Qg2WeXwiWxfNpafsfhNWcXry2ajcn5GQkPD
9XfO4FXXHsMdcnUs9IMYcEqb6xk0UCXFm8VGAbaheLlqxpZT2LeBDe8CdkCvrRb9
Ch0+76DPISxSCloJBJ8B3iRw2/n7hJJQ9ligiVcX/Dd0sesy2SXCLcULYq+YfEb7
5qqRmrs44QEi6IIPeLPcHgXw9hK1Xm9GM5X9PBf/pdzuZHcBjgTXCQ89BamdwCuE
a6msT7I6CE0ae8ycx29Kf/BXjdokKjuf+b7gPfOD7ZzQ+HoSwaIZOS8Gq+ubtIjB
8rfcGXl/xkbU7u9z/CM01F2EiC0LLY+2d7B5nbBhim57uQ6esqmfQgEV29nN0k+b
+fE4ALqZeEzlsbeWWCLXZ3BSKiPvtbuuCLNr5k5HJY19ZWYQMYqZkB3tTss6WeNr
l+iI+LcCypQ5JUeE0OAWV8uSjohIMKa4sLQcehfGB32SksyTaLJeqzXP+o/S/SVW
t+lH7es/WKKIvtjlyJffiQknvuReGh6Bzx2LeNkwnnY8iwM69ne3Fw/eXO1KW3XV
pJTOhfFTPCEvm9HeWNFaH6pElj6z0JrLVWpcvP7WpVrmAYCAx2DDljG4dcLQoNMF
320ftwf2Nx+rC7HdBOplmR7aSCLUIJp40zyoR5zWMe2tnBuvom0ezivbyB4sJ2wr
DnR478NLvXatMV8rnp5cB/cI52gNhHkKn+koYJqzkX+3ABcXsrdS2+v9VfzM3B2c
WI7KviRecN6MQwFNFenm5WW6aNG2jNLa0fXfHLQ4t9+vKtBB2eGbwPQ/Rlyq6/7h
RR0ue/6v2MzZY+tBkXgDhO6Qgh0p5EAKEMqaIEq0A9MRDD10ZEyZeJ5antfwwd3I
IedOmSAKgP5P2fHUpX/S2aIy7hyktgCS02eula7D4Tcw6s/oIQ/ZbOYXvMAHStEb
veRecdCyq5n7q4N1cdZDOt9oIs5+PKyjB+hUzAz2+IU21vqhIZsHlxCHi+6iKil6
LFNY3SpQLbLtDnSo1eEPO3zSf6Da9I/gqhRQitJ5MIkTudsSlYBIgkLrzDddj9LD
ITsg51COZVzNUN2Dp9MeqjF6dP8xTWXScN0VHTpQAZJ3F1XJBHVJyd01rNYJXk3w
qs8GXp5OUS6gE+CAH6XMmduQNO1DwTzy5wI7m/H03dhrrRooshOMPGa8s8FJrEbU
7QuY6rZKEPDASjg1/JRZ5mno4Ofe5ITEvgAFaM+LJW1wIVo2adNCnH5sYUZ8UbDB
OE32mf59sOSUWX6cHvi3FG91XUdV3338X8cRfmVtDbLIydYcS/3+RIa9ih0/ITNh
gd1vYaDfpni5muOOX6r0Uz+7/iQP03JW4Y18weutvyhhTQYY8VUnPAgLz3DJvDoe
69lKcUZJvm3uYNUojhFYRA3bqgJy8/MMF7Vg6uLICLKljn/n+EV492bLb1G6ARo2
LDuDIC0PTWpKkvxTd/vSF8dGWgPw2wQZvWhtiT5ACKjINMouUhOINT7ylfxxDAbT
b7l9bQvCEnwn7LdIUd5Fas3Ma9gprlYxHXmzRK9hwf3AJ6BCMoYysa9uKM6bY2PH
`pragma protect end_protected
