// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZNciEPYPjHeNb6ghNbDGmXylShzgBGoD2Orw1BwfVo6JyYEu50Xe8Rb11nCSwkV6
q3IlYyLMM985K1EaWoXVEgI5y+QP17SGCSa9fXzZn+bN3nYoxe/RlWWmA2nnnHvR
Rz0dZ5D05xkr9lADmJgVkpvJGm8MCdXVMsv5Fiy1ZOM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13840)
N9cOeCnNdS3wGYJUjWqSmUflvOr+vJZz7q34h6pQ52D+TdbqrhvEs/V2ByxduRVe
rAvILNvwkFPzRDIIO0UsU8U1hnC69M+DbDlka0fAUVOw3HN2s28AZfgj7PQoFiNj
Y8bwrjyB1p+QpIHwjtcSKtdl+mbz9vctW8cUNkg6ejC3HqUCamhp330HS4CwjWY+
GYbBbUA0OpGmMvHEXTTj5tQmYJl9GuD/qr8B5DIbrEloOWXywzCtMRgf/pqPJ0c4
Rb63bzBr1UzQd8X5egwjgCoXTuT066S0sFLtaRtXJea8nRpOJJ+dqYsdnX7NcRyD
GB7y3kB9lyeMzCb2uoIxSeRLftqelHFzBcS4WTE78JK7ogDWncuFslsB20FkpW+P
tcOPSfC+gkODk7fdbU23xRQUsCMZUsd6wv2nep+GF6tubNHzJFclBBx/OUfCyVZI
qpfDX9XZ9eNlhwwTc8ggjF3lMEMKdU76exFSbkpB5jymJFb3MtwFrYlmfziiLb84
Zk5lUOQwZpvovuq6Ln0NdOHfr9dpuPEo5Fq9F4GJbHZhYwwGHvMGruwkXF/l4+8s
pLV0kdMcYjY1hVMGahlBjZxCR7CBtnHZLCAU1wKN7R9OqSsPgc+V+RXJ2ijT0+nJ
d1RmCqmrKGDfRbNR9E6ku7H2FKUn29nmG34CdRKrE0KhmfLKKy70zFwhAn7B2Wi0
ojgwsFyTMgmvcnG0cV5iaLasvfSkFjSSeQXJLe+Ou/OjmLYCCBbCyDAVPXEllBAy
9mxOJinc2pQu+MDiEl+BC1s3zsty0dK8XTsk38B8RlLBAbhSKKKgZplkzGuV5Mbz
n+v942OhZhc7ARun3WkxHZPYyu4lKhPwig85hNQh1i2dVKrdQe/QkBS66vKwxp0X
5g67/V3ZkG2jyo8ItMh4yI0fvt22J0r7jMKFyf5u3Jc+oNEZS+Y9DK4V7yE7rTK8
4J9vd8+nFyt95vwkagCm/4WqZS3xm5sc7Xh3aaG5e7e97ycBTZ99Y1vH/8lCXr9/
K1gzxj2rNg0i7DzBseQNJvc8ZPl3R5ojp5MO+W6BI/uGtd/CG4sEWDyENUBO2Nd0
NgB8JPrIyX3D3W5znvE4hGmmRahAj+HwP+ixktKKuD8dsaAmLfYUQdc5Ieu9Lgf0
is2x1UNHbqrUwwHQXeVriXlrlHMyXUrTr8Vf29WZ4qBoW0/qlfQj0zp6c1mKD5bE
TUywgAlHyvYnHhtYKO/Yr6gLNHc9VWIkLFEqquVBDDJuPZOSCdbyNAPqD95kO30H
hDGkXtFKd+SzVl8zczYzlfP1+EB3mjShYaPOn858KiRgC8DySggA3iSlA4gsd3GN
SNkkkFPQvzV1ZV2rhKvxEKCN/3nT7qzHuyUJl6nXuDXYk/aw7wg04IBxIIN0Se0c
qjoIEC7OFZinxncu44APvyZEIVctM5RHWol0+rSZC3j6MGrQ9Wfz7zv6w+p7382d
VuV2TchvEu7TI3H4UZS4eOVIByxnROEMzBl60dWDJDKII1IQ1/JdG6+gll48gv20
NTDbCjPJ07wv08qAPhf6tx4JJs8rOkcqCjRBm55box2mbb9zySMst2Z+MHsUTviF
KmsPorp9TFvOHGC+VqFMtr51U8hjZTkRYOcrPugN1aZCtrUj35AXpVlErJbtuM9o
z6KkNU2UMj75BKJ/cEzL8MCEfljZOL+Tq/SimcIZJ6LnSQwcWkTZdmSun4D97SYp
W/5xcJELC2LN++aEF4Ba9PBFDXfNGwPFlfupTzQvgz26ciSI3+HzvNEJJqOzXL9m
GE9s5NyrznHZn4A2wZ4UL0csHXgLUIEoggMWXC8vsSy/2xbESbn58M3nRD0CcPrh
blDML5gZhFaAe8fFwvpQoDRWZ50sYf+e6N4KNOm2wEwahNaECFz1Y51iXKsi4lqi
FUmj8uIUbO0jlZJxpH+RJcqXQTktolmDERfmnqLgH1wAJM2CCgin0t3yo/uionja
L9ecyq0b/Mg4f/mnPJJ0v/mj+WcEDQmiflW8d3Ru7KCcZ31CPqwBe1E1kKlwtXEr
Wnn+OG0u5Kgx5V9DIdt/YVlmWvb8lFnI8C9yltQ3+qK9Z7uEaJaQ2Txeggxq0kDD
ZaOuwWIYe95Kz1SXICdHG/g8ZIagezX2nQBNfIogZnL76tY+wKW/lLGuIeOebrtT
xjzG1XgxuKiZvunxIOHODFxF7iwnXeBzx2td0yzBHEIvbWgIjd5qOXo/57E8x2xZ
qLRosHsLWLYOOrN3GtUIhRkkbvnP3ZJ2KJRoZUGyoCikPLCWnSIu/7gNzrL1bO2e
NxbIb3/iI5h/xRIJlw8ujevPz5OjXb1D8Cl7bSpWnUvFM9RHM24U4DrvdamOZgDi
/guPjwf9hEDDCvGGeHcDaZYsujeq7iRvFwZE/LVfFqyXtUNtFXothhISiWBwRmuS
IQa1UkOssBGQqsBVYnteatvMDDPn0LscmV7H6Vt0pEtJLUwgm2vDSMZWh58AHlG0
LStuRg3jgbfqEOZVIXuzVuEXwAtYBrsXtJf3L8NV51ss9cCDx/ILiJoZf4lJsfUW
/VzFtg35kZt0nukWjCrtWL9LJrdHDmGTHtocHEHcPuNOt0PQ0ecCkNBJXOnAyCN+
3aSQTfBxhwiARLCSkAHz2IbHxyEAMHh3zPU7JGYmlxrKoXJ8EJVXoOvZgJLgUUBA
kEuflUBWuapTsnxfwLf0gCwE3QDWrMbHn/s9pS9wfTRypAEg45fP4fUCS1K9QM4o
KFf3e5mkcDqEkq1qmAxn227PQuMDAESGD8s9V6s/rh3poKHDR6338OqG1UZvVjhb
Y3X5aAJzjNg2UxrC4hOobic0uQqZYswvD0eI57sah+AJd8ABR50s7JkJ0TRPQOaP
BZLViuNLPyOxZz+jrsFnSfaLVqTNhfHqAY5tAIJCrdRJpvuXb/H+DlOiydd2GKYf
IYb3aCp7mwnOJoQf3CpVs0Zp1m7XXbmm9VH20ISZcDjjWTVTRcVILbD30xPsa6yo
rs3l8O6FU52FpQvzN8Z3G4+F0x8m3GVtzUPWFzzIh0728OJC88iWedOIxSqDZIGG
p+k1gUC42Ynz6W3maGR32gupRAxvzUv//MjLkIaOAMUMarSIbbYMb4iRofIrRmlr
DfbRbhvYtt6YY1/n74fnrDBTW5rvh1WMUo0Wg/JVXgfcY33SJO3BZ7RIIPj85xTx
2srGbjRXcT+yHa4EdXwUKnmVunBk0x9dlIv2jzFrmVa0QGW33oUaiEcdTYif/DdK
cUHmaI3Jjg5Iw4tboQNKinfsvFvUb+3Xi2iiIS8LtQ7Z2obyEXT1P8MklCvyDug5
UAMozsr6epG7eVzUKoe0MsJ9JEAYYsexDPx16dyb+pBb1IeG7b1LPGmnk69tL3uJ
+qwhQ7258MkDBAoKYT7l47GvTlnmK7Z4NZijE9fo7qSIKyHDWGmWgZCY47A0w4DU
yKYfoQHjA+q4VZoQOVBAkfrFoUHoYuhvau2C/JxFengMBnCqPjeMiiVZSNiFvmfB
3wvs3o8x06GnxuxMtdgDHzGDzNwNwLFVpr71VDW8WUpYCoFaqUTqttJVrqISl3qN
WrAQyHj5UYiZsCr7CsWYHHzT9WMAQKJq0CmhyK10/LTIbGCZhmcJNUVA5tZ5A5Ou
uqizFRk8V8Qt8ktuEZ2OCO+U5uHaLyY5+/CqFMjbpEeIXkwVwM0/E6tPycegpUU5
VIMt8hCd9Lkp28R8daoSuIfyeRnzlGuSzS14D9CeK8P+TEJfYQCu2EOvyAnREhmY
IOKbhobth6xalxvOfAdx4j9QES79229MsnEP+ZXEMyE5ML5lKOWqTzJVKT0+maNd
0RPsGgp/9RJKV93vXnLuJdoIh8W15U4wpo2TzOqc/ulST0+/sBIhFUs7k7l/yjM/
yqvH1ezMmCZyWbT6/EHPwFsfsqNzLh+IM0UH9QIoBULCSW4jGH4VoU5BylT7XNkx
rTwdCJalwz96y1Bv02oc32r6UnbdIzUDEOt/tnL2jQ7NRFBPzp1UA/ZrQ+GeuVG3
zZjkiHl4F+np5HGX7uzTMKEeGU1IsXF7UaJrI5UL02ufxmliWxxDAfClx0A/fuCS
IETwbvgzecmgB7SRJ/Rq/W6PWicLQvi0JrjTD8acjPgv2BHOHA/QRXv4QYRUpB/X
ZRVd6elIeZJ0ykgk5ZUm5d2I9lpsWqkw+gGwQ3VGoe7LSzn2IWaP2Aalg7KgYUxq
cb1x6nNMpnWODp2kYWsvxf6AtlEKRxGBf+bMGjvnLa+y1+CNn5ojHaDmy78+yBVr
1+vuXUL42yx/rUUW1D8u5eKQQtEJkeA0uLc7tHx/s214rwoSCPqQxKzQSbE/28SR
Fl5qBPwWk+GzgMAjelKPeDVqOP6QetR6HMmUx2NKoDr++X5m8LumqPmQg/hb9QnT
Z2D5E74Z/tLlJaYI383Ghi4nR3MbJM0lsFJrm9iOq2k7avnpc0zJ1fQPYL0X8MnX
vrdAC6VJD14QJeCz+H5vZSlIYdcnN1EoBF+L5Gdd38hPaWqxS1be8BSzp35WAllC
D4VuO/oLqzihrGOBsD4ZCqUEIFNUWQv62AgoQvONfDWmFQyHYTVBFKLt4W3ENBRf
a6cZ4bhddf4Tj6fjsZKXExSyPC7TGHbXTTB5TYg2X5zK6pB/Wbj95NyOA8xKQsUh
thpUGnH6qXpLP3zOIJhUxZYTiHR2es9mMTgLyFZdgH/eNSEKoCtmzV2qA2c4hmuA
iEEAlZxB4uNunt9MNg9D/PCF0Li0NcjWnRLRACjt5YuSz6M5rUqysUYQrNg4mKMV
XZTve+I6AWOelndxOd3ov6umVEhSXL6YMUzHB3mWyj2eNJcwSY2Js21zwOhyZNvM
rBN2GpqK1IH9FK0PB41S/ANWSxg38SlyZklngIRsjCBrUiGKS2DBrIFury6CQCtO
qu2U9gER5FTyeSJWJNzo6vhi6ZPiyR5mCsc1DiZtILF6767FQNkSZEV9W1i+cqkz
PMq7hhL0JxMNOkp0PpZQyHUAGhipuVfXPwti++7wlMNl1q9gXtcM4449Lon2sPAZ
5+vWUg/7hli5V40VpEzKwX0ec3v/124EUwp09q2WUFOsdHMN3R3LLmvRejIa0KFo
6WM+9B+rR+d06i64vg20YtyNLWPpGPRFoZgwCzZsdfrqBv9Vi1i7VJhmHY0gce9Y
T57O1yieDVnkDfe68agNCRcsDO4VqfsW8S/xPX+SaLDvBGxzm04uv9bpIOq0KnyG
/5uwX04/DbmgKD236y9pTbpSm3WcPS2X4nm8PtqfxJPmOdtbH5dCVwayApH19kR+
DExOY8xRJpx7o3hu4kbdyZnbtmlUHTTrEEDGhdOAX5rxUvXcgJyzUCBqIhPcVHL3
I6v/NTwZsvpRctfkDGDAKRQ99nK6nTIao4A/zjv1BHlgdA/kh5zKJnnq2nWu1BLd
37zro0Py2E8oQGhysWnHHuIy/z6+EBtmbZVffZ/3Hwtjn2xraUwoQBclNl3VdrXA
EOzjcbrhFSbO8zZO4NQOszrGCOXdupowd3zMU7LdWnZwgN2NsTAYIDnzNNocf5zS
2jnONn+G9iPDC3yvQ/JtKfvTPJ3ZgSiYi1eMHVmIOsjKoON9OfeuHVI6HcYP8d/N
+jXxHKKVpv5xrUB4j8NqHp1W6QogTgTKxlpNo13CU4bOOOEJxLYrwCs+SUgqjS+E
gIvzkFBsBO2eXzvt0DCSygwtTdHb20VfKBxEDFLBl2FYdt80Auwe6IEvtyNMcBS8
FY5Q82OeemkfHjc/7GmCB2plPk8G8ImWUsk6eKlhnZpWRSyieLdXy5Llbj8BDA/L
cNGtSXEz2SzNXUYFReSJJTpI61R/zHfQ//aTyW0Z8ISLTce0rg4qhk4O6ibx3ZDC
DhAsq5eaPxzTP6hKydAzcy55IxaTtClFAxbUdZNS+OllVqd4AsB7ZANV2dq15wvI
tPzqCZPMQTH9TvNk3/FcteWuKQ0BvEShWdxoayLPWDcuBEgJ1nljitQnsgWC4QXj
Lb4WfYrPVtWYcz3WxbV46DA5UyHiAaYcXc9JZoatKN2GRnl9hU8a73sQmFHhb6UX
01enVR6kIf4CqeGBPbJ2as7zleHVWgZIno/1LK5URPZq1dMDVGnOvm9hmGKCgSH9
kgpGDNEmT58ojq8NRhE8GZCE255exCXko6WycIMFyQS3RcAf1yGJ+rtwfjNko/Fr
NPvB3LkEzkDysslvsukprnYhIWO+8rl1tn3ndbUl869lF+s8U0mlleZswngYA6r2
vLspOpoxSvluDRwUa92iixhs4zHmeYyprk9ehYg+Cx695JW5L1qIhm/JWm8kEsOT
0mLPzC1uko4xri5uu6ppDhTQMExEm+3MfAv+h+FbYLwMOv1zUKagsRKEyNRMdj0w
UTFvqfmzCgHThSr2I9DUs3VzwFkvS5ZjCpExbvfEKQeDMwLBfK+LISUr134O3J+q
Ueak1xbb1aoGLMdpZDkMOXzl0J8nltVrP18ysn5W6cJDY0mq87qYsf4+PxWAzXfi
i+7sBTPjv/2sdbae8GJ3kjRR4aw/4ZkWEtejh/Fx2DW7dm9tTUOA6I2X4V5HyMVv
MUxcsNBHLPjNPrWqwJzvi8Mv7107mNzW7YNBbhKLG0UuDzbUlqMA+iAaCl3v2pSF
eP9Jg+57BdbcuDvYaU7HhamGcemMBm8a+yd/WqlioKcbMzP9TC+1FRtWJWn0GQUv
us2LxUy5QRbF/tUnx0N6gP+w7ROULXJKEKeplitwNxfhb4V/aeokbjK1DCMopbhe
E3DY1whdAuhDFISalbJJuKQJYM9G5wxeAtET4w3p5H1QVpNiv7OwtHn+HsVJYOWm
nnwuZIKwMgIlf7TgZA3HSsh/B6y7n/R79Bj2akyYExYfoHKfbcagrTWqceTi/Ip7
8XqfRZi69sU30Nz+SqYeM0goCT7cIXYeReKbntPWjZgOWL+5OWhgqydREGZpRxEn
f1jh2I4P5NBjSN0eLTHn4dTMkC8UjMJ8blnI+zzhW671kVxrz7uwj2h6td673ven
/TGDdQd2dCuBpFrPdDAylkRp3mqt1LObBoI/5AjLteVNoDVlJtRKd/zGc1jaBrTx
01mjOyghYKu7aY/bMkX/8R65Im8xId3b6tpfd7ITnlvB/8PQqp1TwjFejSEtzRJr
wsyBdEfvQrh/PGcqfHg5Eh4USyNlhxc65PakkYhMSBQ6Ven/f+J6pR61Q6D+i7Ca
EBJpnq+aTVe6oVvGTKLDGk2hl+RwvX+y8XXCoV/c2M2ns4fMh/+Zkk0f0vNPwnbA
Zzbu7/piV/dBi98bAlUctWjgjg7Mgfre8NmAB4j96HAhmZTDDcOjHXpeWwg+9aUA
lOb7gWqydPU9CS75s66PjL6BNmUsmHqHRP4wUvywTNnJeMoG67Z2QzTFetfW8SWB
SYOkqSaSKkPH0s59IfmXO2GQhMEzsPaBmg+omc/Cd0nmaF3j88HeNjm5zPKt4gpz
TgqqR5Fv2hAt1WFpV1Z6ColrwDoz/WQljON57sc2nzdRTYf2YfTfFT1ypJ8ou0xr
tD5scRRkNU1scbyRq2ZPxcFJGEP8UmC/9QvzOEnYyTmbUNDcsib5ZCeA8vc265WP
75YyBeDN9YRB8EPeikGIIcu53fQlWv75FqRi3lb1po84CF2snrWGFabDzoSTGGgV
rKNX1wZiHoewX3MlqTopiQ5ZQnROD/jJApFOc9sKyjqZP7twBPXWnpzAtSlbP4Po
cNjWs7PpU2ARvEYJqsxFPuFymVl+rvsK9Jexm6QsHyorconeBKQG84FW+90l1uBH
4CxC7sI3Qt9UbiCw66fIVFV6ORtdmPDtFzI+GO9aPS4GJgaTd56N+RANjOoQGKH+
NIpz+osRjxkf6XfDkDxM7YPm6oXRS6dJugPb3wZOq1ACS8ugstA64neqOMzznCX4
JhIUjmzybBXhbPjSpQNaEC3g702YYzLyeeb576/mtUXLgFMwLAO8/QEM7mdaRFH8
QrGlElYjaSFHFmsM9p1olAtbG6HrFJMiTRnR5rfiq/HKxmeMOjQQ8h914TeiVy0r
9C/UL5jC8dZiFKVrhw9ndFrKkn5KN/mvCXwl8kI/Smq8uq/cikqcwvjY6y2Egrfn
hvO4QBzFRzOMvzg8VZkA1f4lLgo+m3K7guVCnd5gJ81+4WzYUtPqtTKyuF7laYee
wXH5ibpv+GeH/G5o/76DBO+Prb2hFS1Px22VjedBIw0XmQXoNcoYTPpMx7o49Zge
bZxarH99FbBD381rwAb1XdqDeM4kVGCJabbDwcsQlsCEHWB9VHQmVExaSLLDlXVb
NGp7cjBEwLdOZYkIDAh5OB/ONz2ixuTpyOgeyEeIKKLXutJfcoA3hvCair5kdepC
QPwBj68LnSqxW+yUZdnoKPGdepPH0i96d0iBBRdRt7HucB8Fbb6WOuFnAgbqhWPU
zkgOHmIr8R5nYFTj37Z/MHTTYZvOQ5QadaUBzp1QZSLn2NpNDXWasNnHj3o9CdoK
BqTHB2DeXB/667pQFRgaVKJlQGOK0Dg1sTmCFVbR1uG2ZFFJSHf8VJY4ZB+B/sci
PqSHR2czCli3Zm7Q78TDfpMXZC05udiS8aJ4Fk3iAkeVLbpQunVR9lC/5TVzRJMb
xdDxqJMJEQqydHOau+ZCjoJavEXwe8O/CSlrd/ZzNzg1WQHh0HvJyyVtQ3A4TuTw
ydKqAQYb6CsvA6dqOlv8F8glXD6lIWsWnu3ztDtxDf2+HaNV2tB7100Xc5QfS1U8
d60ctj8VxoOjg7pzA6I+7fyJjTbFgSEj501TzD7Us9hdEzlfaWXmJeJpGMiNPu5C
uZ1YA23r6u6ni+72MFVCkK6UcqcAadtOjsCQTO8+JDIQz9wleAGnwViZUMF04SP9
9AuGX7+e4zgLn3OaCTFp3zMwqt+xuQfktwEuYCXHPcdPeqLAnQ/vwkgYtthlqafJ
rYfPD5dxvCBkojWVAL+M8HzH6UXZv+qsNl/H+ZBc0EiU7qEWT1HhGtqLmvR4Hpxx
nOMfVP7IDfrJbqgsqNC3RetN6IvMFiFlVjFOd09FGgLmRMSHalqPHmBn1EMYsVcY
h+KxNJu7D2MpfXNrTgPGQVeXMAzBwJKwfgR9JuRvqVo3OU5hrs2GMl3uE3gps+73
rlzkf4LSZjItYYStPPhBlBgFx8VDJy1Ci47xVypOl1I0bb+zA6kIHcuaHlqzbzNe
1tYoq2UANmMwkKkPsY0JrCHtoXpM6ZmXHxwxx+08rcSK7RPnU/HxLT5Nreoc0YFq
QrjVwGD9J7G18NBwjwA7sH+DW99MHtHXUHDUvjS81wxRcXxKAgSsCLhNEiN70YQc
XJrMagrxcvPsw7X8D8iWvxWOcZfIwqFwSyGur2vDPqFYg8zs3XlvTXU3qDfqv8g6
kLHDu3YpK3r7lGPoh68Q+OhGYqs16Ky1iBeRn9IN0HI+3FJhO5mVty7kunVRQTsq
zjxndBqBdrescIeIMQlHZ/NFG/0d93v23wj37IYYm6Tg5mXH5se5VCwGkbq7IDO1
17USeosdUchVwePICh7qQidZhoFKLGQh9toYirYmPlSpcyCbCajp2LxSINj859Xp
MF1+eQWN9tzoOdrA6hosFsuveUKxJt7dZ1uYJZEnMmy22hF1HqzEs6cztmsg11Ww
4hKG2C8ZgOTQCtSXREL5I855PxtNls5xddtGETo9Gj/xieILSVOO3EN7Wo031CCL
ooTH5zT8Xe8N/PSoRD13+oB5TDeQHl39+YHSIpmQ4+SvS8bByGqcYdjIWhJHb9k5
Iffjzmkuo1Svke0ZjBgd5Z58rUCd7ezyO+/iS/U9+UsWkZ37Q20AFNUzaOS88LDW
ZMg6V05EQxmofM3nsoIaKX1ajqlQxTVND8JM6bCyLhLjyLI7AAoRQvnjdmUEmCDp
HESaVXQa8bVBVUuRYcdwoyXafDpoQs6r0dMp0fWymg5JalXWKtwmaNBuIrpVk5Ol
EVbLkZb2gIofM3Fg9afs6u+NZRmEnZYzRgo8HtpWqT5w+VhI0qVJt1DCXUpg0n/L
ufY6NWv5ycIkI5qhmZQFg9EeeShnVSxLcuhlxsFAX87+TXftU3CW0qsgrW2H3HOf
GwF/M47MOLTbeAn/E7lJ/3vSyLenvnlnTr7kavbS/dwHBpasUUcWC0LGFnNHfiNK
HuwGXxC/ESglPf0wZbTr3zF4Pr3oFt1BcBJBaJHGGcUd/BYD2UVePZsgjuOUwe3S
iLDA278UAPRZSgfvFncWlyhArHBuHZFCwzQnLEH2UjYR664yzo9MHhNMNgD5S6KV
46JzmScFE/oA5M2uE3GJT2tZ96BjR9YI0Tr7qKZAViu5SpDoCb6uDvprhK3OG3Js
1vhHCLWeNORxIBVDbSK7MCn3dG5z1bfttD3ZztOCkWJ+vbtnAxR0sx3aXrFNdpIP
JmPkorVQ0XCPT0CLLAschm4+IXP5eRyViZMruTmswXnSiaJ6llweN/LBi4GRGLOJ
PlzM+B9FEmnXdK4ZxtqqjOLmjnClRUTlg9I2Noh2EWqTapJM1kqByS7wiHhY1qAS
idOBBDlsQ8Ax2QP7By6BZM6fT4/jnt8yF+QMHXqqC9jrAauRq7A4FL4v4ALGl3YW
vVc+HzQpnlLp/uqCQrCa66AgxYP1dbGbqf87RjGHYc6M6nAXDcA3Pk0a/JjI6/iU
lDbzUySqtuV/QeB6vn3TkEKWHg0WADzd/J15j7LDi1QiItB5gDDgYWIE3qPAVaks
EiTci4lNSiUSWfdQWhPGNDdehgpAwWeNsC51TfokdX/0lcTh9nB1dPaW0LPExFrw
0qLS9lZbyBjpA57CUnPdZLs+OGrZzvo4F1WD3HM4Jrv1eTf2lNRYCseu0x+OAHK1
d6oW8Fa/F1r7vAQu4LwjHiyL7zQkBmnB4eO0FdFjAm6jDI/0Vyj2wCc8dc1+sAR/
yB01R85Df9R0Pjph2udEjRcWoSrwYmE7KM35t3sHi/C35GnwNetD3nSRspYasgGR
uTYYiU8VlkneDGoDVTyfM/77RpfEZzhbrpa/5sQ+ZmSboEwrLVdJEK6kdRV51M1g
8oDor1khp5LfN8hUm1TWUjK1C2pEqnfUKHKL5aVbWoJVahs+dcMJGW3L2DBiqjOm
MaBTH8ObbZJrOLtEMDrzRPscQ46Imb1dyJcVkgyR4oyHnNC8G1yNFRE5kx19QePv
xNzONVfUkXvF//DahjPtyP5V1qrsw5tpy4cEDdivNE3d2MvchcftKBwjgKGQ4LmF
0Mo97saaVO83Bx4KQq0j9c8yAYIINnOiQ+4hBVsDgc+m7Hm8yvL4ljuO3uMpe4fB
jp3VjB9NwPB1yMdRpVWx+VpPY7Y5P2Azg78RZ3EaZIBfw9PSJtkQqt85z0KoQqqd
fZeio6T7OsbZjsooCRRW+mwMqfu8e4RIMcs9voFDeJPA3S3peHyMr3gPx72hrdMO
Rt7T9WygRtbDFc7lTgdG7dijaFfQDGkpDu7ttnAcwnZ4FFtyUz66JbQX+pqrPW2u
i6SnpN/dtR2HFS3o5ioi2tHv4lYBHN3tlfnu2hlwRJSGRJSuI1xofmB92lPvVpHj
pFuo94jgfBgz3A5ry7HHBz6aO9AalHa15lBDUU1zuun+Lmc2X+YKg/MZJIPXS9xu
m1hE7JknFm8Cpf/ARPUee76cKVCAxuoGRqakph99pjxPR/GysCss9nKU5k/d2PJi
qFftlDzjmM+B3yPazznwZ6B+oo1HMvzDEYMJeUAYzVVCYWOKlGBrHInRVRqxy7wm
iTDIoONholQu0T8QtYzxLhy16Yo9EppAgi6ZLqiH7Dhe8cncZFKOfd3p/1FXESw1
tr+eey7nIpyVr70/Y+4gYIOSvhDGebUE57u4WpeUpfS0jpWO3k9oYRUyv66Q0KhD
HFfNgrjg/zVDkWEluZg978JrTnLYtNFYnrwbRNxR0ptGHDdtsHNpduj0P5pStZPd
Llof1502LRsKtLdyaU+739TZNlZPPVKu1bRt9wzSR73605KsTuvN4U8H+mLBoL7g
tF5WLdq8PF0xoT+a7U3/WZ1/BksISXuELDTLcU3TmI/t9kiLOLbodgdjHhzd2BqW
k5q9HFcZLf5CNdlOhLlOJm0Qi6N/ounbJOdYCYqJpvQFb3AdRoFbUrPmoUX+QT1+
sAghmwl5NPIYBYViQVph37K5TPu65/LPsTmJ0hQCS6dyOKK/ARKf7rFm4rfw6z3I
ayYF/PcTwuf3coPNYyu60ma0LwkWAF73hFbHX9rrycY6hXlg2nbu+KlK/7b4FfDF
e+d/zJQyZP1kBkG88GhDXZVuudAWFu4hICyOgi2o/jYKhW1usE9LgMhhX2kGhL3O
ihqmPBncsTNz01422ONO00XOxoJYXTTpPt4NBo4GHDc8B6QI0BN8oY/gds30cHCd
TSz5HVAd3HsBXX+nNXgo/Qrks3qygruAeKLGL5WC6Tj1zYFPqog/uPt1dl/rafUJ
7USvFN8pWMF/lYzfT4SW92io4DJHpayS6DNJmJEYkTQ2YULL1feP1BGKwuema1Xo
dWOHgVFTA4hwQGq01oXhkNR1HAXYzpp0rnVL0RNSFu8+e3W2ZH9RKTVVtOBDfgFy
XX62s7cLAvHh/DCkv2IRsPxSdKtMrt0tkYJ/MjEMQSdECuUzn7jzIfExqN3PX5gz
4ORCO+nHYwyV+nXd2HTjcsLknsykGFExLyU/fbvsit5TAGm7CAYVPwn6RkWlsPog
dPtahvAa6fsPPSi9lkoW37RPAHW3mF3Ee5TRJdrb7WgEm55zwwBSabTmeaEW+trm
RfN0IxZ+6FliTBuyr/3d/uo30cBUCB+axvUp7rRdl/4+Cj4NrvKR1dyQvX9CeRde
l39ISRgCnHpJQliT6zoceUyUJ40pfHpqSsSx0cKeCyqeL9/rS/yHTBJqp+hKjqtZ
TkGNeZCBGxtQ4MXnkyhalsYdlGWY++Qk7oZVWE9Yosbe5glrwN61z0KhT2/3V+1Z
1CDh9S1BeHYIyL0B/zYTcI4Zfzm9De0WHNEB74hu5UG/WA0h20i/GpDIvdTA8BsH
2vAnftdzZCahxnQpwkkoD45yWpgtsksokNOzkuHiJodcyoqImUy6WcdRjAGauD5S
Pa126y/3bO4EUR6Co5D6ndjKJXobtNOBIhSIIr6L20Z/X8WDNctV3BICHNFuh9kg
/t5uk5+TxEGXgoulc1ksCS1ZdawS7hnfSiAf3GuZqWL03TUTg3N/T8fprtAE5XKn
O5kteY8v36hyYZ3kV2HOZ5wCjlKDBVjMBpELSK+TresTiWRaPdh57efh3jrsbJdQ
5bNaRntqoIcXVr6xA1nDcSzo427jvdOOQDbZeNjrF6Ibsj38i8WyrgvHjHNMb0MJ
DyZkeFkuAkeoRzurT++TGc2gSqFEBbgbU3bK9aDTU1iac8lYDQfmjCU7wbexU/1G
+FvpAPhTFaJBa6MJgEAFMMGMgKtDmvjKTSZ7105/TGa1LKaJ/Ay+Ulrt7IWa+zdr
jaAsXlKwOS4/3IoQRgix2sUPlKzmaTUssu/W7EX2Hp1YxO6nhg7aMCjyr5Xk/AVO
aJv+8mXpQuKNyaJe2GTxM3WxTXVPfOoC0QlfWosAznod7xTi2SDTwdVhpSBEH/D1
YNHAb66kDK1FSE/FwMH0ymUAPK6jSljLuc775NEIDmTm85nhNFKV4OeZAPVe/DBu
Y8foJmus/jjqvlTgzMRm33jgiFKx7iB1z3+RH/jE/YD4SAzuL9gvPYabu6RWqbn6
SEQvcI7Or61olZ+BffC8e++47RWJdhBOL156S3fyVtwTt4uj0NMg9E7EiuJbKVIO
ecxHftaBBafcWt+93BJ4+FSFLxRi5SfMFR4g5nuxWCwYAB0eg4u0/JgM1EweJ/SO
OwpTAZXQjuWNIxfWFe3AbXh4kqYlaxbdLRJWyuSiaJqA0ymArpf4n/YMTwIFNlUX
Tw/RiIwBkgvQ340p3vHWTs0MwoiU3UfPUXYtG08DT7MxBJqqJXuZDCs5rFCweDKb
NVyGj9029tpJpnh9ZzJrVG4lCL94VyWtHQrxLRrpFW9Yawd4lLHewN5X/9/+5mya
Zm4gdQCTJgBS7eFNQ8zo93CYKAyt4FxDe2CDJibT0P39txqXBvBxZb0bPjSJGOwL
UeCku5DyfdIO+A66OpDXBMBT8lQ/VIa1H0BlKZUEAWXP9DaU2i9NaLbZZ12d5Cse
fcfQ/eBUMvrPeeUa/Mon7YlusJJXDfQbB0Z0HuR1CubyRe8MsJJYnLhAl9X/JEKm
CL+uahpeCYUgOpDoVvT0AH91S72q8vwEg20pF10IElNI9ne90iLc6S1NlzAF5UjT
nvxZBTDGhrRrBiW+ICddOId0v+8zXF4VWTOjRBbnKjD+L8bZi0NWsXM4euaFOXDZ
SbpuN2RWPqyk45WE6FBlgfMaTSZHdW/RFFM6DirMR6LLIH7F68bWAdUB+9LiUayU
VYY4gH7CLC6o/UH66kvP8o00R0pllziKfsI1K/1c+g82M6pNOcxxTgpBhl5OfSlx
Q+VJ9M+ybkIMcnxm2Y7TKtKivLySR9+PQnW2LThPXWqhMKevJPITCba/PygjPv0/
2vTrrg3NURGNsCytD6bL3jTZVy2u/Wu6MIh4/KEaluSVN6XYRaSyydADbu7CT4fT
oiorIOWS2ep2XzenRDv4HfBXj1K/K9/55tR7MWfOcaM6zFyRzOZypCHSo8QE9biz
ODlCkCEa/T7DnGbnz3qITOWsYLzcKfckCTeOt6XHA9EvH0wujspg4l20Mdj4xENk
CFa3S/Ib8hiLGKU4JHazu9agAmmHo5Hzq9CGfG6m6M4UKiwqBxy9Uvtr5BE2z5vG
12R6ClljfacTMhZknyMmpB/xxWfbbRNv1oFOCONqD3qOVKVkfQ8HGoJ1AiF7iPmC
P1cc/vnrbrRftO8O0P1wbVRYuCHj/Cktvt40kRqY6aFe6Bu1H+7OkG5Aq8IEssTB
hDzao6reGPrpMNj6ZdAOKlH9BNB3J0J5C/Qb/6F6vI9qtmm3BfFIk+PpIG/aVOiv
SwI9Mubn89aYpBQqJy0MQt5Hdmbcu2/v136gHTEyIcnEuEvJ7ppji+Qzvvtzu3/M
i6UDLFyIC0WICG4Ky6G+g4ssto3/DRzxYGUmNxKvVElXnkECt4BZCnBhA89LF+wa
pCE2ipDAymrOT18U1SOTBzfr6Dd6tPyPDKKTKyfOONo4SjTkqbTeWo5tOLAnx37U
uPfjhPhsa7QWf2w7Tnb2oSTtRO4HkhENJ80mjIg7sODUTDvJgWkV/eJNUhzc7Pvy
yG9V5U9XVn+jLUkGNwaQVg5f/aRF4AF4XWC3At1hSpySEbG+orfV/8T8fkWGhsF9
BuIrgrVeNJR96p0s2crZNiuvpdMzhEcAkS9dTFkinWGmSDPxnHSXIJva2+U8jAIw
6CDludAeP/rT/W6zL1JVeAn1NLitQLXkKZRhSvwivhmQYOQ8z/U0bUmCHztYJusr
vIab5WuWa6ii9V/dd15ULVaOOnE2V0HltkxKm2Ik2Bg82Ye8RY/YoUB7iXjzGO26
Qvq5hFQBt7uxXGNulq7feVL2cV7vsnnRNpLgtUkNATSFPp0/b35DR6SlP1arjG9t
nkqohS9nrHzbS8IvDKnoIp1Nr4ovmmskfcmVbtMpzHSZx/Cn4FHp/1kMuJmmplgt
n8bXPpCm5YB/FBkEUls5hH+elTyXVmS2lEQH1yi+AFjvZmYbssAntsbwlA9sNGGD
bETHtd7JQPXJu+5G6HCWJEAspjAP674ICIti8BbH4yC+Ca/MbgvcnjaeXe+55L2C
DKH7wsTTccMZIKPsiWzBOl23KcJjGguKwjyqQPSU4AgxitUxs2ziQAbtSx3s8qE/
Mw0yYZL39sWqUTcNzyRwqogl3YfqE/lhciLdGQZxBj7bUJCFr06XesgPGCwwQtru
KVQf+nJAdf7Y5Q8hVK0+tQXwD6N91Ru4havda1LiCdZJ+WYMD5+k1Jkcto4w7kt1
uFFMXwKN97/4of4CR/3XlxfOaeaUcfpR68RUMaajVZTqLtcp9ybIaFrjzlhaPiV+
eBokL6G+ten/S9m4xerfF/sIKiGQAbfFNy0lJZye7EMNb4GU/HjcqddGlaB4zOPD
jTh387MDqdNttfrKeMKJIBuOjVwqo2QoG7u3yd6Pv1zJ0UFe2V1aChTDkFD4IWhj
1uynl2S0Mar/Ia/KbvMpZcmAr0IyUmwHmsZHk/TsdsGfCEgxAvQAcwJBnW/v6Pvx
aisAQ3tOM9+nhZDnT7CIcT4WZhXFKYLBHoUBs89ZX1+vLKU8gr6wYN9c+mhponLd
p2h1bXu5844aMjfCCRai1/ljpFFSClKZq5UVsFBksmZsEf9O1ldesJSG9t9awfQ4
g6mGtA6VMgtTDjK8xAfmsG4gSADo6qM4pIWVWVKHDSbAzBX9TNfc1Ts0iN5TAiy4
gNHjf/J5m3Z5781LjtepBtaqCxDWP3QSQ6YMKxQAxMXP2xdJrWGyPMJE+8NvYyBt
FpUGzsRBfiDADfi8fAN8JZ8Ih1wnzxh8mo6Dopp/+gpK60H1GMF3760vnqBsSyeJ
39M94zgHGr95auB2eAERBzkYj6keI4VuXk/6gmsPCdCtrZmDZb8IL1hcqorFKGZN
amjqZ6VC6NibhrhnDEWWm3QLrRiYQc2fKEQKumEKefYkygQ+Dw99MPBn9OS6I/Qg
iOmRvWltwesLUf4h2C1UosawkZuvVvMoOUT8MGpifg+QSizoyNMfT4NFwfIcB5h8
QEVVLuB3uSlBW44uS5QZDMKxVlR6qGD75XTM1zZkji3LtIIbwJW9VBWI0Pm2JIII
Xdebc4i6SmG6Itbbe4Yv6CGFwunuwyLSn0DBSzif+Q/4uZLj6igVGLJicxOGDjm4
kZBsUGA8Drh1o7fFKKNP60INZA7p8ZYFRX3oGpbo0pEb8inFzXE4au22/C6vFoXd
AjvYjpdZFBhk0MZwrl4+nN0/VCQ47gzWgk/ioK8WhKGILLDcU+PMhdxjtkLYSqiW
CalJe/orV4fJOj3fX3h0Nzw/TflMPKnF9hwRd6B0n2uTFXCYuBQfwpHvpU9gcdo6
tSRNoUprNZR6S8YJGW3otUbQsRma/PO4KZBKlOZAWlYGdoQkEPcBl3q4UUQHQFLz
Cw9RbaN+t6vr+m4IsQuWlj5kckIz931iTl36My4ij1MW9Gje5g4O+DRBw6heNq8a
tvhVtVlSmnI39eJIzdGh9I0xl4ZleacVvv+ffT+F+OelNm3VYBBRIfVcbc3puNwG
VUAqkouW/G2VHAEVamG9eZlu7Pv31zwGeeyx7LoXyBQ8y6PtDsoZ9IWNFDzZrv91
E28wAYTLGYALw9DpDtoEdDNUBbfOTmySNWjOKU+7auOLIDnqCVIpffL3gk8sSUBv
MubDnBGGIH9xRQST/ANfGK3OeoIGmAcqz1Mo8qBVU9K2ZcLWpy19MgXkL/id0m6j
Ms8fS8WMDRrZ/WEiFe5dUWR5kiRhydLoeqQiiI4iX5K573sr3gV42ZFHILvb6nYP
k38Uj5ANS1dFIf9gutro7Ndzh/Fn7NT813bBnpu9mo28bX8SoEQwXBmkm1OLcIbF
ok5OHsqamao98Lbhk3ArSC22YbtT/EnmXGmeg6wQ51yOeZomWSXZVMM2kEfxzyuI
kklA7T0poERA4AD2xf14uQcMAirq48FU1oUdB8fjBcDcDATauD1ksh18al1cgkX/
j+v4fCAr7q8RTUMj5fUnyJ8qXynpdRYhkF8dLHkxqp/T9uOV4EK11s0V5x7EHHjK
mhgz6BQKRyQlokoktFtZgBxJcWmtP+pQxiiKS5cWoy9EDWG1ODAFsCqGVLcGZBqm
0K6c3I1CMBahQQKIVLgrMROKV/DJAo/1+CijGLcITgx4VhJoxlkPeM533DeQTI9C
8Utwh74RXkDcKGC6Deh0rP6Op4Pkkg8wgHULO+z6h45dKzMmggL4yJLD/t5U9gJO
XJyVpmKkJ1TJFCXYSPnZtt1I7gq07uiIuPrAoCNiX61mCfgKUQFuVH3kdyOrnZ3r
2mDq7NkrDKFlkt32bAw0VK9k5VNfOYWLEDibKVbaUhHt+UJwGwzgDdwygiw/JRUH
2OlhjYcCDT8/oTvhhfgdKwt3XOq4bfRbT2OlwI8nicRwAVOqJwUfWRWd88fAh11H
HJ0HJ9K07ewN1MZ1jLyVA+JKzy0hhrE8xpyKvqZTlD/sZnp7tmQuJWsPUIXUolxL
bzXXEr4uKxqpaZpkQZxk5MnOW4gJXJplXfB+KOXRuR2hZBe8vgXxjMw031++sKur
FhAPMnBFcvcdSCXtaFHYKocd/9Ryc1ykvVqGZRDEe5jflXwdbgHCj1rs4c8GUtLf
grFpMUTzYewpoNcxDK+mk3yv8a2pNrhT1z/H5nTPhjDt2JYAX7fKkIFgBJMMCih5
u9LlnyBE+mH6qaQB07iV8A==
`pragma protect end_protected
