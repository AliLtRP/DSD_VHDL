// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
aXVcDce1/S52wM9p+DNbqLOlLdbyv8xjSMYdPq3LcAEAjk8AcSDOhRLY7QhvT/gu/ijmdNVe83zT
0w65sRBk3b9r5KeI3zZfnj81M5JkRA9qpcOEe5HH4QBPX/oSQW8R2Tt37IQ9o7aUpcNlhNxJuDeT
J9E5u1Kj3FqH/j/6enOCau5ZwlZlgLwKdxhCEPVUq4PnVKvwRRD8Ifjphsf/Bt3+uB2XR5XJUnpl
1tLgjj3IiR4IC/wqGJ2sw7GmuyVBMcFIKdw9EfCDOaiFEXrqTwvDLF1QaY9yzzQrG5alKHUM3gja
gmFxqHCcXLhRMPjBLq+z1N/la+onLwh6cQeJ6g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
8CIAzprl5iDhM//b7jfnAl69EQx1GCgzUa/WEkRVnOBXrI5+fUJRCO3a8WuQzOpUjWXH00jG1GrX
GZz6cXgoC+kkEO+7tGNyOHDpjYltDVxiCfSHfSryd4IcJrZEMNCAf3Yf8NHJ2KSY8buBDMgsZIC1
nvDtes23PNKe0DhpMxg0phZCoAwRF9ouNQ1w1lK/ua9HJyRURyCdIsEeMAWZHIAKX6Mus72zHhlm
iemZennEoGV793ufuMHFA3H8BqB4QPCBVyUv1kZ/oa2yuvCV9yrxe/LJiNZ5aEsR3eZhIzuydvQ3
x3gmAwXaaRsc7W8KR552/qGI+Fi+dMHojs1srT7GIx2mWWiRjSQ5gsblE4gKs5M6m39PTphNVYNy
KZIVyRqtuZxg0pz2SssKl/7kyAV3s9SLB6yLh6rAoNqKDe+M96v1hRzgSt/PupQv4y6wh0sKelBr
xxPats4BE4WWXWE5Ni36ed9GehJb089pa5BPD0zXTRnhFU0kL7qlI13bByD5i02FTOhZuZXGR+qz
yxrBCwF41zw1mKzh80DDL1TSj8ddNmzjuf24kZnKCbd4amsnuYb0el2CfcGemJS/h9/NtP1Rjwex
LL21tw/Da+dbzf0qL0C/UoPtHp6bbEPLF5SIyLOTerFShWZ4VkNiyAcRizDOrmadkTeIKCNH0U/g
fRgqkZIJCZmrC3ugh0xEveQ3tC/MbPCUDjG4KOQKPw4QlBxg3oSk1ypjUeIQivr3BBQ3pChRhhsp
XhqfOZBAakqisp35rmrgrVeKmWwqHjsBBWwU2BWx4a6gvBDmYxxOAFymarnTvUxSZRPHjlhtxqcG
CfDuqeP25/RGFrzAGjX6lHZStvePR3JvEnHqi6RfqBt9ns2LNOI9QKY+o+ZxJSSkCqxfv7+1qrNL
YGOvVVyRXvCr6SEhR6nFKl8hxJQP+hImvJLRcztVC92aiXakT6iGY6VdR2U5qtY8CZddfUYKbv+V
rLx4RAb8L2LNNvuTYilPLH0WdzN8Trn2io9PPBrDPKm4XfQUj2WKcCyK2J7PP+6i7bWZd6fpVgte
5m/MJXVykIrHhETqA6AgIOyEpBR3d888833pC1/GJGUA6HMHGYO3uaXAMN3h7mbzr6YxuygE3Kih
wd7YlMYpfY9Yuq7LlMJtrlIyPPuNF+Od+mPDM/6hIAGm+yg02VU2SuxtTpvJ+htVoMvNcr0RSTv4
1iuzffIhLZOFuOg5lY1owmQ4ufJYW4mua6EkAubapq0B8ppBljGl6DquQrJ3t3EZ59b9ocPgLnP+
i370ea/dG95yXTf2J+1ifRyXux+2rWQZFo7ZkLle2wrdqjtOGWh7ljGUg/bcNWR6WTwotUbypNSf
bvdyRtzw+AXbOLZQKcJZMz6smdQXgFQSBzunagXHn+526ecjA90SHDadK0xHR7RvJOxlDu4+f6u3
4DfxWhBier/GEGJzQnl+vzkuAW211JnrBxI5q0Sks6QaBlrM+g4OHCrQLsc5SkTEZt5W7LRGetQg
Mx6+BWtYx2JfES4KTE5Kt7kOwfsdRiK3AtfddDipqttPsUVuhE1b+WED6J91v8sw66PtXKW1lSAz
jDiIFNnuX53h4M4XUA1T6jZPH0ZBPArqcWdzqSrSJmEl2IwP0uw6rqcASdcgIBg9ngOIIy9R49sJ
ijHH+/t1SE0JL3PKLY0yag0lBFw7hh0uk0K/ev5+Ar1tKh2cCT//5yz3PrtIRgn4xyPrFPgTOYre
yW7F4wz7rAqRXBEwxS7eSbD+H4bAJY99GMLMrrJ42oSU68Ztn/kq4zEf7zEuzKOltxPXY9CVre57
CEbOCbcTH/0VG8t5CwVtGVjz2XyeMtFRSYw+fY4G/B2QWQ3AZJl8Cu46bQwFM0tv5R+2QYzGOYYj
dtLJRRDuv9P9Fs86auJSF67wsxlXGc34WaMthEyoo1q6RWTa/vdqsxhn8pA2IlTsH+1hib+YZdRO
y0xH1Yl4/PS1HQW4Y7cqB1D9PZY/D1/BiSGR5BOMPLbs4m7OSIw7ughXHLjCaZKdBmSgROoKcfiy
ZeOkDYwVdkDick+zQX7hC9+Ab3ueznZEeYYIYLStatKuJgvWqYTHJyfuyEsbktYSHBakq6aK7hKN
JPVFYOPLIWRkLNmcBC1kImQuEiPkAjHYj+HLl5q5x5bUgSuByAd0cVUDqcexeSSdadtmiF/wJ9ln
z1zDS/gid7pmi8mVX0/nUgwLKSq1YHAUcsWYmJE5fb/DxegevAQU8Ubl4l45izqYgtHUAUqlSnbH
/lwV9SYzQQ70as+x/OO7dsTdUrMz0cJhKBSebVlSVsVUMb/AGwXq/X5L2iQQUpdkoDqLnpbAMKnG
u4NUbRuRNBmZo9aDaC2a9DAVlXkMpyBa7N0/Zi2Y5Xvh89tdIi74m2HxS8elgL1QReRu0eho0Yz9
SDyhrYnYsuq8w4GLbB3UnW2FVgtkiELmHPmihHiHMP6ZpELu19gTqLZdzbnvIDqQ2NPdhkmhsA9+
GqY8X3+fwCosPYk4uzZsQ54YjR0Y2TMn4Z6Uwp8Rf8GLQojt687NLJJYXmNohWCt2wu9f1Nq5ZkZ
kT6zrJfeueckUKCv+tJTinYz4WK8DzEkK1dzynOGbx1KnkYrNhWhNMUG7nuSzUxyyGzYpOw3sVgX
V2vCYzC6mKi8OhduvKEPtcYUDH49vm0KFcBIzs45S190fIPYEpC4485uNpznI8Y5QUsniKTEvvdi
iEUv4M21vry6Zsg83u6VCCIIzzfk/NHcmiIaxgGKeRCEyo33IDEOoXnsvuT/qL6jpb8Fik8X8yIm
IS3I+8BellL5hh0e9u1uoLpXvaiU4DRqPnadMSvuwYNAhr3hnJ7lD5SlgP+XANZXTC3MKHmT6FrM
GL4Gxz3TZU5a+1uIcCBo+P1c6j3z/uaB2OMjAUVme13ihe9hopDK0jpnCGoRAPW6GcfWiqeXn8l+
EeM8HvLVN+pGEOfClMxx3D4MNcmr9l/1Do6AOoyP252iuESlXV9faUU4SUlDKYVvVmc2ejo1x2Cx
KcWY6z9I6cDhW7EL1VAVPsXhfoykv7qs1UzJ7aZQXrmzdV+AkMSVxRWkj30WDZQJh4+/RvrAs37d
aymaSQWszeay8f84+v14tWip1/s7190GBaRaaUCZHtUPKEXm3BLiF3RubgQ6zX5xHHt5ZpoGj4N+
sLfAfUEjk6jX7/ENXzlH7pLd2iy2xC6v8F8rVnWtAmy/NymNaMj/kHYljj+21wDH7STihZAv1FoR
gQZVTl2EnPHdKlQOyTWdZCOLjermyRea6jjQx9Ua4PySq4Egux3vbZPpZHFQrf1ID+BaNLG/qvpD
s+jAhfkfVYiCYOputtjlMTjy2AJf0WaCX6qj1iuxL9ztQT+KFQqdX0B93hLwBXKN9Y2JZBDqVIAY
QWk8xPNEmAOLjc3RS/9ye0CLyUmw5UbSZP0uHERkeqqPSb4Pp87VWvK156iOA7XbhQ6YNG3rzHCQ
FQC9y0pPTbECanDKWpLmgTmq6ILs/QtkDDL1OOhVWR4DR9migxQyrOcAm5/u83Mz8nEVnXY5TzIx
rdAASGwjH0fGAkY9c9lKF7aXiQGOn1oJXA2kqpJHVIBRrQdEBBW0jvmN+M760fRe6VI0vtGTrAUm
RY1Z0WrseahPxOI7AM/3oPWO2ac5ySOeBhBC3LQwqQtONgRnWo30IedcVkn3lV8jtXBoP7W+RUdz
jpYebdsVNq7a0xUZ16FBoIZ83/ugBs1FWJ/UBUACyArf9EjDxus31d5Pt5ZInUQgp9Q4xffR/ijZ
WigKrrmDN4nkarrm1GoULa19W1++0ZT6cDRiPp9rdAVF/i1317l8hGXWnTPhMY3zei5xf3nVAiqf
YUwJvxyh2VVTBpJws9pPlrhikXhYqzZSSS8poDj7YApqvZjsnbnKpKTEU/XYjW86WOCLv4tSSv6q
ds/qsQppRfcTqOpkoY9Fy3e+TjaV1LhO4UeIBrKcvhx50wlSGp8vKaGVaCEKU4GpZjve3QZYPS5m
4ZdCEjS07bsdd+lgMDBOjQYdZQzoz+JiC3TpWctfpfkdLd1NbGhS1pjyHCT22D0HQL6zciyGSkW0
ghCZKywq7cEWT0PuBc+yDAtINl6pzoFO+aYv+9prRF7bkImW9Gs2cOyjpqwuUAuNy2+UKiphYnXb
XFwUdo4d+M8L9mQL8UARMmk19yN7uQ5xIJsAn5Iz0iSIMT7HK1Zv9CccXTexZudTFVcx1IGKfYZX
kSJbmlyOOIvrAoKaXwHkqhcrwjNU7HNeoRvH/4K1Pw9a3DvewUvgSdljs7CJy5Iq0poVAFWV897e
TkOQsdVTxGbJvLR6U5e9gCMqK/zX/37+EryBmgDh7QMk+7XnDbL0mRfptQpo7hQy07ElIa3JHtlz
eQKTP5MbLI85WZoKiaqj1Gy0YbLPjGD1sKjY8xmfZTr+gIHvVGWeNLrpdB0a2qAXxvKs1c0i1izS
8e4KhmXn9OVbIwsLfKJLsXPlmp/HEG6JnAr3ccTRLXdx46gEtHtCw7KtY866ApEJCn/1we77oyVJ
Ws3bZZnkexJiZ2FiuOor++zEzmYEPgrEcD7la50TAMcd0DAUAPuCOMeyMl+Yg3GDsucULO2MYqaM
KupFUwVYCn7pu9x3OrPwRk3in6wCbiT8fR0FUSAQaad3w/+uRIzXXCNzDbP1MMYywuTcMyG5qzty
UB2J8cS7paPDvQ3EzfKjRMMJP3Kzg0ol2lqSq5SZ5ixsVFpYXfpSaaQnvodfdZfCxe96EwfK4VDF
p3HhHfrk26n6EAs/1BDepfjwyQ1wuZ9PLb7Avvs3En3p4kyNXAD6g4tzk4WwSnBleDyZgyLm+W1t
gKqZIz7Q0PnFlIsjsKeVYwcKcv+a3OoyLd/sutm+dIOXZwvVGtyvX08ZSth47eO7H3vo1equA9hF
a7QMziDPG+AvMkkvPFYTAzbIyvAFt+9FrHUSqGDDVouIxiNEyUlO+moXhUj7pBglaIQPLciUdcWO
iHCeNdyh7wNc9v40YIe90c0tA8Ks28vpJb8A0BOdTqeHNUg80sLZDzMHwIPp2T3CA4j8abXs/SvD
bebaTIrvA0OIeXRHPeqN8B5g2GLvVT98lBKrIvAmMuhrcNLzuj3resFe9yrgOu1enUbVnvFDvefR
VRQhO1zFKc03hYuGPYn80z8NrcRAqaRRgk8DccoVMsUktrJppdFSV03pW9AvXdwpugDDkIUeUrnu
s4rJ/1j95n660f4jHGhDlSZDiqXkpQydkk8SAc9BzIn308qZmyRrWNp0cwWU7G7y5D3a4uLW9nR7
Qe4zYcTEv92KMkKs6AoFSqBR/NkFoJaABO/FDDBt8/SdzJL8OylhncBMF6ViHu8yN26HLokuglkS
CTzIlI08dd8mrL4jxPV/cbBpSePGQENlHa19hSLUP7fohlPI6yxuJ1TtxeKFhBcS4kOlOmrr7K6i
/gpPtqPQCwL0HTb0XMpsaiSHndvZORT/b2Q7JuMdkMJF5et8IOgYQlY/a9bDS7kVEqa6uTEa4945
GrV+JNaZyHJ5DZFEg0Yfu9L8stDxku0U+ZHb/AjNRbsdxR1uP4e6ILrilGgmvV6mgxHD7dDS6vxE
9Wx5Sc/fujEDAevI22UEgDIc9ZmeKUg6SC43YCYgIbCVgRxw6CqP6cx5Aw2DNJR1yPgpU22PeJ6K
CMTWGM1vRBny2TWqebksLirVbzU64ccT0AcHO4Q3dj/i2XfVefDK8QKr+6pZWU6MOUcAR5o5zYsf
b+xOYUAsWXLT4CyGirtmD49BQP96QP7LyuMvU9nuCiBEamNZUG+WolGGIROHOkgHZlc8Q30EanYH
mBqmxvSTWVeSsAJtNKBfNWnq1Dze4vVf+XNVZWPVI0QfF2PQik3JB9aJzxpVGFg1Hp8PlZv3o1w2
cDI9rdWTuAwXCNmabkPU2V8mtTxb7ZtA1QfoUSsm+OzhMflC6HVetOUo+4LoAjI5Qh23+ZWtBhWB
HzFGET4C3dP1OsRb5C2CpWgbBpupI7EyC8F8781ZjhS8K9ut85GUpkQZ9wqg07ew8bP/gqF1+i+H
tWtTLbIczPNKGvqLU03XoKMvBST+h+zRjuVAhMv7POodJmpIJE2iMjHJCTQcHaJWvPrdFSpZAITz
R8+23NQN8GLA26CV/SbwVcFFPqHOUbvlZh8s49nA2ctmskYxbKLT4AFsmyOTWqbMy+saRDYBbnJz
ImtZca5MGaC4I1IO6SrYr51Cr1JiEi5jZipv6/6ZQ5EnHBqIJgzd1/CMBSt9vlZcf2erqvtuYdTv
bEBkYGRe8GnAleemVuY0+Uw0BD71YZUe9bZqE2sZpIAbY4TsRJDXm8VZcQssRb8ynLNNnvXjs6IE
nGMzAn2CP1BmwAMANZpqt5ImBlXFJZIlaQT4ufL2+NiCiGx/w9TxUW8HA6xxqXS0RQCF+ZA4cWpS
0t2nTiG2g9YV224bLTK/m8EIkToRai4+SrHJ4mp6IFRLGC4R4BAwbJ6m8uNJA9mbLK/Z27seXPDR
NHor34CRn3gUytm/OnsoY1g3yVNQ6CSiEmXOdPHgbk2dhOx2Y/34zymGkDUPbkKzKYxRS/rO2qTi
1ofsKEAXgBixtuKFvPKDOawb2ow9fI/v5A7JNvU4BoknRN6j9E508cbMx9BZwqk919poYgKj1jra
4CH9ugR+3NhnSf/mWIryWe6HjlBxRhuAuMS5EYM59jxILGx9MjyWJsEkJWST1WY6zREEwPBCsjjl
PXJrmPKajJhhADnyZuoAyit91xr7kVl1gQ2gT7yo6tLxVvsU70/qmuYnNbf/hs0yB0rQDi3LLaPO
3RqrbySVfxkGWoJbX31bavGbLYrnPLarKJXrAIDsjokQwiUn1CS03DKwFLA9mpOgyq2RNM40hbN6
d9OZno9BtcPZ3DTpvGudSV8c2sIzSOr8CRRCdtPvmRX+fmI8oTRmJ6HJFz1imGO57j39wLy9TtZL
cLb1h/yZTQZ35jiQg+IeVs/xX7/1eDfLfQkPdh9EAoeJ9+Fmqw/bzRi2LPzZFb57PQN9HF/L+hBk
KFrQVJoR/ewDT7RC2NsYphwQWCgeqNB/3+OcgiVRozCr66koGCGkM7vAlIsHpDEW/y3BK1XUXq2r
gHxALN/DcOf5FmusrqlDRYIC7t6vewYUdKFd09TNUNfeQ7W+GoK2So4fat6hOwSgUSiOJ7nF2HmN
WXTd2edUoACePBCeDYoIzc1L4WwdoJgZ68cK+07kYDfANtpwYTjcslXDHk0P98cXWFz2UAoXf7kD
4UzRuP4wLs3tKGFjvjV6XzXg6rRNTzXX91Dyy+0j+oWbOC47tSD97k/SSBosfM3XEPG2dQRfiI9+
IqD3Xbppxcpcc8WsfOpJB2YYBhroEBiKWnY7onxn8qxx3r7yeIJxXkcfI21VbGY+x+fICrj+kNMq
xdfru4/oT5aJRCL98XGOPmh8RQeaY1PkPUVCqJmeTUanxzPaGAuvbrWWAkkStbGDLChOYeWIWIzo
7aZZMBcpPbdQacFpY/wZ9ABuqhP4xNnctws3e8PnkZAAnd/TsEyHXk7K4Dr43g8Ou+nr+yIyH/RF
A+lyaM750n9gd/NcpN40s/Db8fJTCSbZ35MOi0Njt8ZzJK7Eovye7Fs6xvq3ihK+9FVWlJJW0N+4
0fNXTI2/jA0GFsnVKT0v3Tmatc03FPOEvoIyoCbC40iJqLd7mBOpVjcFhPC2MWjh9j17ksnbJ6aR
p1pUB40t8LY+nUW29m/rzAwOQJS4LjNDaYFlZqvr8EiL84xtVGohwEcceL593K/SzbYls/Mq0oVS
Ebq57lADJxZF+2yUWJ80yIqKSRVl8sEBdnfs+t0VSvkqqVgRhRscwtYNu1v1HSQ0qVynPX3EsR9C
RpTM92ogC+2hJsZUdSlABYAvAmRxdpm4n2jUkJ/12YfrdVM9Fx39H1KeEkFeipz5WroNacblnepb
93680Cms+gQisrM/TKYBxtlyKnIEDllCLq/CTw92coRIm8WVQ7vQCsAB9EAD9O9v932DGTJT0EN1
x86+I3+BmdvdPY7jUKKn2PsoOWqeGTAej1dfwR0nx32C9iAsrX89phg63+pTsdoIC+RBHFAIe6oX
fDRG9qfRTRrFt82GOJYND+3IMCAt3LYgazBh0CPUR1VVaGGRT1t/oxSL7R8amwAQ1DeFR2EcbYT/
i97zmNDqP4wrBQjRMb8HEDGVGWvIid9WFj9dqVlLx+h08FiAb53m63i2ND1fk91aDL04/CKCrWyC
D9gLr7wo9iOnMtk1Pl73A0M21Vl4XRPnz2lDA/761r/MaUDx8aR466NrYXkVFFALhoBBHXk4bS4t
NER8J+rKhb4q82tJVGNoRH93NnopDkOdy/i+aa9KG3ChcDnLPYtoS4niPDcbnnSWmmYPL4OjAfa6
//7lOhZEXkx0ofJKb73n5ARplP1WSwJ5Izos/iKiF06KQgpdYi70oTIxnMhTXQfSuO7vX6ixJH9O
g9ZBbpG69PG39cNlrPI3SIXy+pVtSMPY875hRaBK1gj5p0vNIKzDYGnl9AcnRftrmVL7CMwsL690
MKaoOxwDiUFD/D53cs8eH/+Vg5JaEa1C+Q5wtCQO48L1zYGy3oiS+b4IHBnSRkebpBBrSGKuwpWW
UigB4T1OSqc6Y4wAU5yQ0WT7sxQhKBuZfwVjBdft
`pragma protect end_protected
