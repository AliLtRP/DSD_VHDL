// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:17 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tMcZbmKNdfQH50oZWClOhEH2wYzAYGkVvkfvzoLXG46zKviPspVrzQ8V5F6QEPXi
ZehbBod+FbphtgoFzzaYRO7cqEs2vtiYDvujZzzOT0wPWorFzWlPhuiVGGJXgqZf
icmVPoIx6LWt0y0sYTy3+Do0SpCj2ofTQ/ZtSAcw3a4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3248)
vKaE94D8+ySu4LFVj640N6h5AY/7/3hwWcEthN4BvGxjqiwHo9LtcNEJjj2za/fk
c1hxh8I7g459a48YgoiceRZ8E1elnkJnQN1Qw7s8uSe5VhStT/PM4GLyLFPX8wag
F+qZv4cSWU22QxWr4XORzpdKG4rjFUG7bjkVzR08UjZjRWaarWdA4Dknv4A+4w3X
89FRdH80xDqMvTY74vnJ6JBpHRx4b7qc4ZKRpM+8PsMjL5MfkK95nWhDryFD6L7I
YzPXR6JcUumyxJcKKIB65C4hH4JhIcUnBT3UhI1F99VLgJOMwp26WKgDH7DXEBvE
edcAhOdcMgmWuQArwSOAu57bhfVtJYRpqI5pBxGq5uhx1NvHdKxjnOx37kamajQD
Um+8E6ikyRPjCXqkqiyG7C0UQxVStNQNGfXj5hVT4cJkKF1HQ/idIiezy/RyNizQ
pFF6DoVPhgu9oqU+T46kXPMqVDwKqcxJ7eA+wIB5B+kK9yrAmac+zX7i9e3A6dN4
NNw5+qoN5g3CPLbEHlFIBlcmijcDn0E2axu/uK2Wluk6xTzjA93KIrgwaboTjlck
0++5lzESnOoNRSVuo3shFi51utR3lRK+s6wvs21YRjOocqSP+t2oo+5x+4wijdyq
KKfJgP8Wvac4PNsExFAug3Zlwm7XB3FtRQ+PN5m1oXHTup3EgwXSjUTeQtPYhGEj
U43hHwg86ftz2kNqHB7mFAJcNe8+qBK7UrfQgCn0JJR9Nc/dJReNMM6j19gKBmb7
yt9sc1Xg9dyrfUrTWVNRPuUuBRWl7PGEmC8hdWBVPnFnL2v0p9Wuj+jbXNeW3ndP
3sdeAU5pIDfC4mn+2c8+OE+CWOaVTjL6yjbbxi+TVLx2UKLwyvfIaRZi2z43J6Ql
7ZUq9v/SgUkMUC+uKoWPwiDwXzsYJD1Co4eu+JCtM1sUNAMTFFRn8V+wRbvquHFy
jOclCctXTWVciqoxw2xX+/R1731tvPGnLJMCXioIJOFdsRd2yB1uEqy/fpNuVbtk
tYWkchH6Cif6LzzPXuweT1KywPAbH3rMm+zUfrS7BOJxsyX4R+Pw31ckzbrU32sb
SmV3r0lekENukgwe8GDMmosieNvyhEE3PvR0P319rwj8drMjDZ19tiLZDCYZQJRh
UmIJ6GlLT5XeQrO+PbNUefy3yY4Hl/o/qQ68Vk4pEMpEFmkFkvqPhPisAJX1xcsO
1XzIMD+XddK5dFR1BhUqIROGLlD81K7SQM3+gAQSTxYnO5iDIk6IXKOKH2bxnVpH
HKb9HrQcHwoUeHksXWOnsdjnD1GHZ7GBd5cHII9eWAtYTfPxbd4xF/JOW7wB/iTY
/osJDX8GrvT5x1Ya1Cb2x9kKWTBdARC024pKHvRJ5o+8FyvVNt3L68gIyiasZPJN
hEGKFOeNdEp/GKuErV0vC9xDE3mJUnHZj+FfLNC7s4QNMiqoB2BwzG49fKsHIkCv
yGI0msvvwwzYoFnhbjD3u5o6ymrL0XGrJk7fnQopJWTIJRnj2irSGeEMTmeJHxPB
MGMSnJSAXEpNlEc1RYACUI5oKeQtOQhxJrRtNV8gvg/BcRahhBqerVfUlAAkFdkE
0eP270rgAg+6z7HIVudhaf3cE9Uf1Z5p3giwmO9iv4C7sKfqZ4QJ+3jIFtbWsOSG
3ntzdrZP93pdRyEVLkOxcAM3LzDRcDtvufqfa8P23LRNHVMCgqyI2RCTg5dtJeUE
uLQYL/0vYZHDx1x2Z7JBRo/aCs/X/yrkdYuP1wQ4opNEXz8kZp4zl8zZIXLx4yCh
iCCfvspne1ywL8TbwbSiYV3Vl0zFhyDE7fh5TY7in+6eNbE2GSaHFI9tdHUDLSYi
IMaITPPpLwuqfuF2HxTdfK81MJlx1an3wFmcz/vlUiLO5hLTBvBOrPfYwsUNBAxJ
9I3sS75eyJOAnTop8K4HkuymoduWnkhJhtJrax57+EzvAgK/QDhrhoCKizrX9xa8
jwOtXUtRsbr833GAmhT4o6hakbHZnw96jUZrBOlkF+PGVHiE/ERd0QYlM+sSVnqx
3wBn5gZZIOCCkMDkwQ/IPZo0n83027tDQufYFC7uVghVnpu8ywEzqezEK8boh73H
iPfO+9L+JCCkJrak+X2hXZqyzTXxWSn0ZleiEVf/0UyrEcQFJHgzyG+iR7CqTd6s
mdalGksGtaUU4+fxVxMAs8e9aTc8njVHIIU79n88bWHVJnoQzSf7C9ZpeoCBCw2C
qridxiHDWgIECBEpb9/54hdXurbgwunpibAKahm2KSKicL7NEzAl4/uZIk4o0WFe
MGlEXiALqC5x1g7agTfY0ybI61LMAoCcpkdS3pIIKldkxqJaJz7P19RhFh9oKDzK
2lH4iDrM57DLDp0COYVvheTz/8/F7PVhaUB8CMbqqTFYgzIs70H+oCyOUuTGrkEW
HloxiMi/9Cia//XPC+9GQrYlEQuy9wqyDir4X1FMgZNH0OiSB3cbD5b/v59I7a4p
7D5lx/gtDazcJBHMkLKtYPCipE4RICkr+G5sgSjkgc6w9M3OIYmxlkCjxn/rmBAj
evPBP1HdXE507egjOKl6o1ST7BKJw7sQGIkczaLMupdYe2xtFXedS+QkKP6jYG9v
zK++j8IYXjb8vAXTYTObIzmYV5GtkF0pxkrg/wQOZN67cC7B6YTnRMZzwnrDHDXz
2NfryeqNZ/FAArkAEnUYY8OCE+0vJHQBFJQ6rZgmheoPtV7QNsUdwPJFeXIZB7mc
Gth4GYR9xtWG0Ra5JfzmK7bEeBMh4xTfD7m1hOM1TqZRQG4KRTH5s+sRfIdoHAEu
sboC8A+mYs+CSehZuSMqv/X7o8YyRth8Q7msh14ppx+UG+u8SW3ZoWAlJlyOky3q
clxqZn+LRe2HydonAREkA7gSmdhBTtJPtyfsuIMqHKTywBAaAV4wLlgd65DKpmNS
0g3nvf9tWjYsxy3Iana/YfQQixY2vdNF1RNCRTOYgBpbuUXCCjjh1Ax2fmrKDX6o
7OCQQLnyb6lbWTLRix7KyasQAU5gEsXGeOa5lzdHmyVR3z5Q91PR561jCCRe4zSN
MYzY0AKxpE1NNUNjyXrd3MVJ2ZFzC7hOkAPc8COij8EXgOFfiAD1/p3AcweSHbwk
FiIscFIb8KbkQnFK3wxkOf349oTktLutGcaw3OeXQEzVGD51zSHq0uLCHU7QrLRP
7o0YrrxudPOu0FE1Hb6VH1nMXX2fDgmABQc4X5U01YYjyN1m+K540N+CydyGn2mX
zS+EJrGVpfrbAZltVjHy5Hf6a0DpDJ328eIfA7HfC1ABhiWmI9zq+JrmibBL5gjx
Hs1t4K6+JmZwXx7UG2T6/drPyLC3Lhmtnrr27F90Hg4tQStyUCHcRFUiiHcr0d9t
Ysil7HyA6AbgEzpdakU/RzAdQadW3tXhb7x/lUXrOWcom4GFe1kQyJmvSDJLEsip
t7NNOcGOqCoVbv3768Pat3yZUWP8rYETcWVAjnb0gNx3byeA8eZNJGzWeywN/rEZ
pnRbeXTIP1+uEL+TQ/X3MgE4GrPxKYPp3QciWX4FVOdLHpWObbfKZx3iMfDk8PXX
z/J1WSikEltgy2IqAU9odevaDNWaouX8lfaqpUJdV/YF2Ppux+FJpUXw0k8k5Xqj
LlRcYpzGe9GGHbhnF0nKP7BKZ8o5agYiSJC3uL2XAljlXp2z75PjalyW42TZUSKj
9Pp+IDKE1c7/MhsQ9jZs/s2nKP5TksIszDA8CMNY7ZG6ziIJ/SYGUEYnkzI9jflE
VpRRYQn8NTExpZZw5j0HlLnQi3atDtvCGahpEHiApwYhjlWZzBNfEAsfprCbwgEH
XRREufqCXsqg2bxf6Tti7GvEOKIShWIoTSoK36u3nOcqDlF4+Ny3zwSXb8iRZ7YK
M1tDMU4lCYXLlGrA4rBjWLJFXg8L4bxeBlJBeNcfsTw9OpQbvaP/n8MPY6nGUlcq
f5R9oqQkqKpeIK70eAIPKXbDc8+GVWBQjqW9CoJR9rDpwf75078Y2XOB/PGJQkf8
z/mI/mYb9sgtCmsAq/BEacDE0ynduWO0KMKv/Af9RFBrf4pPi+FeqKMOXsuE5Ih3
yTmiGuZhVd0WGasBtfRTb+QkoBWuNbGuTGuwIBYXvHQUzU5QaVxrqzndP0tp4sGe
8P/MI1j96jc760gZSRAXWtGiyZEAAsr3E1Apd1f4g+G3qVZRzWPR1TBI3y2VPnqF
k8JtHd4fou4Ol+JP3LeiPHd6V+iHTscJf7cqKXGFoMqhLunedtFyCC38kTFUtsUb
SCX4XfxdH5k8rSnUnHguP3hWBq0dgT8w0JVVXScitGs=
`pragma protect end_protected
