// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
n+l6ahQJcQzW3X8UtbVKWSr9Y7cWJL68Vz1khNm10hla+t++NIkhTo2zwdyGcvUT
I9NcS2jHU5mqD3Jb39X3yoUULfUK0b4bzub5PIaNWLpodYTqWW5uICvmaXYNpXDj
wmq5ciGfITOa3jGIwRuywv5kJYQwC8nbfJD1xYnqQw4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3328)
oXdAztPUpVPa5cmYkuzdGM6pvjhM87k6AYmeg2VGu94tKSkb6uZ9zO+ffbcIIPIu
TiqhfJw5LT50HRh6kxzZ2LAguBZJapLNT6AskdBTRCN8W6wM9NNA1xouwVhx87zH
xPxzrmb5+r+ltQuCdzU6SowiJq8CXT5N9ZGVGtps8CXUrCcPVGKVikT1EURIOiyn
0rbTgl/ui1MGf9cfDy0jTGZeTIaYtB9nxR7EqpnMirlZEDJI3967zHAI8saWLSn/
q7Bn1b5nAR1UZlZskhDDH7Aah7yZZnD0a27duXJyLTpygIrvkBkUqS4XdwpIKtSm
3Qbe3gwzxLTgJrFNpRhY57csFEoT+IvrUdRTZosQ1NR4AMEP0rJIA6E2zfNut8Gr
FH8rQmezZ6/VIqVNA92dxv6rk1l6dOu0gpoCKDd1s0cLYsW1K/I9brMkwsrUd9u3
wBG6W0CxBkolaDdFI05fCZbF95dMrxmL2o+tjhmOJm1Epl8Vqx1+IHCNCyeyiQaF
w9BgMfZlqxcVKWa6YcxIfa555nn4w6lqhMeStZ4jAXxHERx9PdXzo8bh6UY4v6Kx
m0vRuLRlX0nWRK32IdW23MtwBajWubrwxgyU577d94kPWV1gUq7b+5VZMXePlCw2
WFcY1Jf6cJHoVqvKPQpLy2bjmZJHMETBEe5Or8oiwDS9ziO3231M/InRmQoyoSyu
K35+w1OTsbI6FAVhuSkhfNSMnZ/spWzMe0k0BQAerwqGCmGxP9CC187n0egKVedH
Eo/zRbbT0paReDIYqYCUVmFlsk2wAjbUn4djQ7rUKRM40Qd5PXfZ3Ihxubju0NPl
Rbl7ZCb4WL+B5qAMswekmxsCUSnZltmyKjz3BHHU+1y6Mw+82SXSHpktUBcKcA85
THioilF+k6fHxY1pzTDtz7NTRhfRkNAXTdnECau3AB9k4gIiVwB4IJJQv21AM2go
mjkP7skaQOpvhVxP+HQqpNfSorTkWpeyYCCovQUHL7eYlUA7RrIo2ETzierRHUWn
g/I606eqYj5PAYy4TDyfiGcTEaaiSHsiLQT6NV339uQs3WhnmrEMZlew4U9JK2G+
XWr+iDYRSE7BywBecBZ2aUSP6Ivd9zmKkuUQIBAvZoT/bF1Iicln5rQtmhvnHeVB
zmJpkDBvfCvFbgdKzhc4fRN/UjdgXbvSe9qfIUE7LPmpnd/aEX8qlt/yUuW/p30q
35rwjUx/xY+roQrHzab6cKrgPUICplMVpsC/k6S394gujdz29lK34Qk1LzRO+Qc3
Ze+1N1c8B1h+10CrKaI/lgoWYOvk7x/gHDETulSsKxM6waKfs3+es2DhdmkEaSHN
lMWU5Oejuog0+OdWNx1gN6Qld1Ox5W/lNpaOkKYIgUm4YwnFuzFxbayyzx0EpAub
OLCqiUM5qdZqBZnbIf2m6vi/z1Vl7iSvOjCL2/f1q+cTy/2v3pySlGlBikoKzytf
Gycn5kvtJDWlYoZfS1v9ib2t3kdbiKLeXjXOKUSj4tE3smETEG+6SMY4Gbnjo4if
S3gySMo3ff8I800IOux4VNKD/EUZrd2DLURM7MlXcSyUcTor0iZfxKbvhgH5OgmT
kvbPAUvVxzJeLsMxiDMIBaKh5sstfci4sM4v6h9yj+hxiRgzlRDsoJbZKNxv+G10
2sLpDnrwz6gYsz2KydCiTojZxozz1si60BSu9Y2VAkIP2TLAJTRS0Kcshd5b4lm8
L0IknMaPoZTUB/wlD+VT481VTu/jKX/drWuoIbkD7NqVWwv3gmjawiMgSpm6ZEx3
hU7VaemGLJprxrnj4JPlqVxVCRpOgjqWBW+q1QmRKljKJKPkdMLROlQUH9KK6/gD
jUUnfnX1NhHSQOmMspMG/kzKirf7GFgFvHe+rAaD8vZi6MvIdgTDviiRq96PisSe
xo3p/8DBcPZ6VCe4d+uwYLwoXkxSIlSco+Ta8KChzd0z/8v+9BneO7qkL6Ly5hVp
Cjv0GLsJo7tzLdxhj0ZZPsTKSeXH8fk88uCj+kz41r3LpverxCRSgp5TNWOYEJE3
3MMty99TBVoZqPNDvkNvpZV/Jy3UDHHbUyPUbkTLPALmxZdOK9jAdsDgse5oxM48
ZVU9tNIqj+2J+qpSu5cMHNTpY5xspjGWREmH9IByR8mLTsXrTGHw+eSfwXAxw0DV
7U8BD1mg+PNYmIFbIc602UYcpQaQqvok8WTE6QKn+zu70Kw+pAtvMuBybLgcuIP7
aUzqqYNBuToZif5+4T6/Ei9Sor1PNYdHoevRRCL9cNmCn9skBubXwSyJFX/UB6Dx
LkN0ealj+p2Jgb8DIUa9G6+9GXZ/gUqxcqKROHt3xT6lMR7bDbnOM/Ww74A4AqAI
6NtTHyfL4TF71EdPwozPIQ3OCD8ICG3kzjrJ5TfT+PhdQbJc/e8GplMu9b63q8VK
G776v5woLgslbGF2QDmZEX3Wmd0lt3G7fYj3V1fXp+cDzo+leI3Kc4A1l3cFOFyc
2bqVFaifVesiT2OBrVhIvKX7rn4L0+/NK0ao37KEupdWQ2ZjUwTYGwJDaDVguRMO
SMLEVUdDfJiQaN0zsy5pL937lbxkt3h6h+FH9PK8XH/JXbgR8Y0AAqDNlqXhyxd/
vimFH9LMrg6spPa5umjJmmAPWXKAG7Q3DPnWv02EJoeb4uysQNUG03h6oJFC/RSV
X/DtjGIvhWARcbrxsob0XPDf9LhjV/Mn6y/snflZNbL6BSRct0niEsmO68ALMVQg
GW0oEZ2rvGCAfMDKVZeG4pXuakaLlI8qWw6gB08sY80oDqYERVD7zVs3pQWiS9H3
jzdeiqYQtP1KW06OhJDVBXE8TNL2Mktsi+TQqwrHUTJDbvb+jkiZ8pSZ1ZZbZUgN
Kx8ZsUCJ+SITh7/yFXJcvSIZqkOO6brc4WIS4SCEDiB9FhAHY4it1+ueJsX7X5zL
eYKy2UlcdqRpQu7F8JSWbHdqqKLRgJ7Yi9CSKTJXYi4Ym3lrMfZAcGAPjo7UVfUq
dMCCs9pC2152dDr8VN33gQXGCJR+lBRjJk5I11lP9f8KmDyOC0zMzInhE0EF2tnt
bzXxzc9LZ/vxNjkWhT7ZE4PqZviAgqyY1C3QwfLMjjHy+xGYPS7s9xYSBkRY2qg7
gLc9QXAac5FnTEcjItMfhmlqhErCHI++JXkMAsj08w/EpAE3bJ/W6HScIBO3YTwP
kRPIGOmacRp8Gdq2YfUxTLNS3jhlm+NktJQhuaYQJQ6mGNgH70bta4E/ShfmIyyH
R1DvGWKKUpLi1IVm94GMzBDhP67380DOmHxfGyI+M43BG6KAo3bjU8eKhAx5FYkT
T2flMAZW9ID1bmb3zuMhpbvwwT2Vc/AQDp7Ua+wNOuC05C2FSK7ilVroWyR8l5fF
c1b+zMCWu/LlNHrqf4pPzC4JjLKauAjleitSc00NehfAvUjvooW970QpDBiYTQD/
YTGavbz9NHDONkRVg5cWUYgressstb3jvT+WPIAKiVM+b8f9vO2AFbv1U9jpgodr
oUGQ2wAdzEO5zA/8CnmLcnN+5h5iiE1Kx/pYXUzLd0R5SSX4eoVNfdP0z+nn0c+m
5ztazMfOE2ASDBneNS4Pu5iJhEK1RFJpeO4Dn0T/4ZMh72mBRu2EF1Li7cEqFNre
nCimyoG/IXPRYJ6aw+UnaRQuk+5DuvhsbhNvAFgE1MI4KOhWQUaAP79EZrZ01VIa
dhT4VLoIUrdQ5NJxarCoREuOzdwbklbR+nAB79NPrUaKnic5ECvESZsDuvtUocnj
FinQ4qX5sGo6UCipsoA5Bfzcq/e1HiiEbHsYs01DfMvTKuqWPQoUQ4fwqXhP9RJF
kP1QtDs2VhJDGmynLyIy6wPf+GiOk4QQ2z4L+QciTcu46giBWufLZNnDzfLIdQ9W
KUjcPJhpmm9pPwWoq4QHlcIf2S+LgAZ/2kfczPYh8sgxQJ+BlpHNLl6jwhq96wve
DReJdD50TrnEnvqd6B0oVjFlTvDyobulcOzxXy7MCY+bN3oU0m0A6C5mFhW4wyCW
BgMxvlx0R2cxkjqvD3js2nT8Fc6tUugnuX1wwCWZvLxJF2pv3ZyMQWeNHc+tho4o
fXdP//aSAajYK1t7NFx2ZL1XCFYL2G8Y8gosnmIf+a1ucfivKJUHxuDAkHXJCrf8
zW/PjmRQsAhf9efl4ZyfXD1mOCrjm/GOZDfXzuPFZFT0aG6xHKpxk3/eUrzv2tFV
c7jrfn2TEOGG7gQyNXHg1ot7ePGGca0T/X8T0hOfcXNFbpM/NbOX4HN5oHR6uYjy
AUkuWfl6SGPFy4ERRzLPO5ChVQmmcs17Dxe7P3TukTHc9FpbCplHrHIxmEr9Z4MD
PaEnWWzmw8Iigxqu2ovlgGmGfSjklGDAZ1O19FWwB+hYnwlaL4zgOEcMl8CwvOqJ
OMUgGMav1P/jl2O/BnvVig==
`pragma protect end_protected
