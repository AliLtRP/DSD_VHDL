// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:19 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Qvejcg5GLkQ30bDc0PbecIo4WhIlCRG62bhmkCgJz1D46F4UPZEuaHXLdQx32G/P
4igw7IfJMY4Zf2fqtXkchKuWPIGeB0FRaUmSG7CBeUebFfG9C0EMvfkQUYnCZuYU
4qbyrb4x365qhIaOaPYF1wI3yAg/Eg6sm4VG/0MdyMo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15552)
bxcQeFtI4vQMVprXinBl+MyPPkjqi42Qjbw3CkhnlJxLzyom8kvvNujSveW0slua
KE8TxqsRaXbvwSByJJErTYuMUQZhP1UjMkz341m7JSYpam5H7vplyJ0eGhVih60J
eJuv2HeltCvvvGlgNmtsJ2NOcR/0uceff1rJpFTqbcZZ8ih87irLZ71qZqLz1mRi
k7B+nCCjYHwtGowChUaDfiBfR+4NBMD154noib+99zYg6bb7NwSkNnAz0OK6Y6DY
s6exfcYMwNZQs3Qxyj1OXxy++VfJrv6RflK05FoSZanZ2D+K44csHgjRgmDAAz4G
H331X3vSZ55K1jzPJJdk5AT+K6qB9ks8ZlBwrKs8Ee6XgQqwGHEYN9VXYUNF0h59
bs/5ASppm6yLsWhStOshDjI4MHCAborpFTF02r67U9i535TqjD46kO3avmMWpY/F
9EC7iuiQJxovDbAXv0XUIFjIRg97kQOPcPLEvat64Via6FXYIELM2FecM34wIBCS
5GEg4EqsoEom6qWxGndwhp06u6YUtuG8WpAWiLs0mhwCNppKcpW+aarR7DI6M7/m
/fH4zYfE6pdMu3K1LOcCuDOoX4ad/sOqDdNhVjKtcwk4nPqp0FXmVHtPJpg6XZ4F
IqL/x/oKRE+Gu4NE6ooGQyeZ6cWc/THaq5A/tTvcfO8n8TkqU2mXosHdgMh2tGPR
A8Evql4b03upFuhlFLNAjbQRLH6mlHrRnAK6WyfYlCQU9Gha01NOM39N2aUQlFNV
yAZuhH27JdZQiE6xIxO4oEMSmM/re8UVzSC8D/ZkIJZy+B1r8hRcNwd7LsqIsFh/
UCr844IdAkCGtSLMVLwVvJhf5mAhggL8D+ZMQK5HdHLcGlGM2M/cRuaDhS0xw+Mr
QQFsztoauhvgoW58kyHtYZ49kTPCMb3gow/87fRJYQvhB7/XXFRh7zOmtVe0DKiL
YS7HgdR+kDo1powe0JjbYBgP5ypUorPzY/J/IJhZCj2qy+rl2bX64xBmaQUXwMa3
nYUiLtRvqFhqpxsrvE4mPeexjWEmz65p2VHhQTtWgMcafrC++yXZLxBxtzOTkKko
LVOCkRZDMMDkUbC8gTXLktwscQ+vHbIoTG3IcDNv+SKF11cCd+uXWtwm+0/io7LY
jEHrBqmtPbO3PvBBDNbHELhhWR75qWj9wYdy0U6d9Ebdq9J+MdqmGp6GjosIDVoo
8XnmgNmE/QtDhQ0opBYGiJNeCNFqcgTrTfhxpeAYlLQ/l1bDU+eez7kw1SIJq1NV
6cZd2S5yjg0rmtFypwsbcmODK2Sj3K1zfEkVDeqH9F3kfHTKhRyFclzVPpBwXQFz
oJMTvW5L+75oSCyzMZ1Q7u/Vs93Hng6POdzFneya2Ou1QZLujho+UO/mRWuEinU4
2qiSptbi4nZL2SOTq0R1VUvY7xTxxjoiGE57//b4TNfGDDXRWH+utQCkL5/vd3o9
HEu3GC+jwL8TYiOUGiwitdr0/GwMX9L9yxHyEvQXTxKFonNvvQ6Ylj82WXN+fLBl
t0nUW4TE1pVs4z4Kw0E2NnqdLMlS2qE87Ylco4d0Rehu5T2yzPS8qW7DTMK1bXIp
ZUYKU8Wc3aiUB3CP+1OUXnxziuBP0FjekXpk4QD3V/d8msQftZjM74ibEWhjM+7c
jZWGslQ1qBqIey4KeaBDgGPneqtElIsgxbZ06VWf/ZpQy4PXVk2gDcn3x5QeshdH
zFoXVNL4p9xFKYagurf2UzxjN4P5v46ZJp7LXQELv3Q/ipbYXCOPvGr/bQiClrOd
rKExev06uMf93UiXy37tXu3y79V1wPgXacKiEwkpnYd5dDmXXnYL+ibWZLYI+60O
DEfqGl1rqhnGafVuUAVVASYOYQ7UFq3IJUV6SNDUJu1uBgIwuz91rucXNYrcQQ03
tTN3iSGHgera0yACfGJ3X4JOJWLJ2rGWP81BrMALS7iwLCd/ELNY1jd52xbkWAJB
QmJadaxP/70tbXav6ZQVzuCdH7WpjEVWfrmeJsTgYKBMj5QG5TcYYiUZFLKP0Xji
6CXXRJsz1m9NI/OSffrzXud900g0WNxSYF2bqKwrEktAPJOUZpjVr7fHFDBdZwBK
Weh3fB8IO404cjJa+ErW7BEjZN/S3Qk4+yQYhRzRkq5N49f+qU5O9JKVHDsxumkE
64BUn1aP+Sbidb6/izmFll2fvoCtqs8u8lGuS5zw8ATtFEZHGdMxO6NvFSxqPZ9a
7alrWUuBNW1a2ZBamGyE/twJP6svcOZOPzGhwbKwkgC86ZyM8kpekTALsurragt7
lkDTQAWcJnVS5HJOwello3Vo8XrK2r0+WbYtYrKrjcBZOhImiBpxr5IvAVkdLPSb
Xey34VwAWJGXbJzSW6wiiRVzYT8J9E1XjAVlCiMsR5lNq1L3aij2L9lkpotI9zgT
f02j3VQHBB0i3QGymVipt8qeWTPNojual0x7/EX1a7Hl6xcqyCG8Fopuj2NQHAKx
ivcPrsRgJcEJL2ig9hzZZT3Fu+83Ua18iurYzJARKQnf6ObCdd8PS0YlqmWSo/Yq
SaTWMri3KngDUh7KJxh6QGKR1kW4497Snm7ncLvKgsjK63o1Oj2vGOu0Kw1tFZ13
4Z9W0YNYLtT5dBi6lBWiRHOk76EQi+T56JOP+K+eX/bm5i+AwZkk7C6LnDINCcsS
jsFOf/a5jAK1S6Hnc3qVYYGYL5CInq1n0zfUBSCaSBLhzx0fCgi/HcodPkWf5fyC
1RXDUdzz3ujLH18osRphJuvgdXl7ZxpvM226Wh5arbPyc71+KePRcnPV6Wp3Ia5j
DwTEDfm10NHxSoFvQW8Z5zH/3BDAxhnE1kfKns9RqyxMtLZJ/RF34FZjr7RcZLrT
Yf/p/gRLhJySntYUYxaUckrspEEwVQ4SEIPOg342NqcvHCtLj+08cN/SaePJikjZ
W/y9f8QWsiHUipZPH0ONuFQBT/N695fUCozY8rqn/0EjVolqHOwuGqyaWNTLwAqs
XUHKRjaiAQaxR6mPGzWE24sbz9NX0uFukDiCyaHJY89x8ofq/RzGf4Tnhtsj20eL
e6wQu0ftjKlF6TqTSTF7a/tLv1uN4Y7W1WHftWisUQpIbFOOGxTJ5OTxPuufz8zL
d5tooqEmDPcEwMhwanAIWYyOkUTBGF88UGCD56lVApH+tuy5QmANlDL30Gnkr8FI
eRESj3WgT9CsgJFM4j4r3U661Qqxrowfsd/g0q/QK8MuS6VGuM6PTS7CYezp17ac
tyySwW/Dni7QQuZuZT7KjTccGnGtEMpmEzUUNWKlJq0igPI5wORoqmtOKLfO7kCE
Lhu4KCa0oHbL+I9xfe70o4otLQxGVAvDJy9asjcqLxtxsToCKWB+6YkMKsXtAxW5
Bcg4XCkgtFV/kL5vFZ6pf9hVqnXOxzb3aPFZ7qX0t/yfSTE/XwCHkY6RAfkQxc2M
WCq5syg/lwB1a9zQTFIzyrdF45fEpCGLeHLFgJPpfX9w/QW+dgHO0TsFnQfhbmJE
DPPRAFKp/eAsyTYI8PPDLgQnIB/v8iBV295QbO0egGNu8KLVXOh5UuazQB1iCVAC
Hcn+ESfOlT43tIbHukxw/47XQgDFZ2tF3XFOq7cqLC28GKf6ooxotTk8BAWYAaHQ
z1J6crikKWTYKtwZsIUyvEANmXt1QEMzw5D73PtHP1AWEoYxrq4r5k5fjE379yVk
hZlkxDk4iu/w/X8bkzGxldjAD4VVFh0h3Qj5lKIIlsSwzmtX48HWL10FZ3dnv8Gn
eEs04dZgz8vyIooO85G8u45vsYYBgz/Z4eHp0uRz/FMVJCGBVsA746WEo+r8oE9u
WyynUC1ixXYa3IWtBBcH9be9tVNgtYDR0QLPInv3+So68yz39wkLCeH8IZYifK13
cf5ecXE1Jq3Y6QXtaUsizemPBaG/nwiVDLK93zRGB6Rg6dnl8wVqiapieHcKJa4O
BBjcUJ0xmaDznWC+iDmTnfVnSsMrcoVxDEW/rCuAEX8Il9h9iNu79Y9tJ8FjBy6e
Z8J0G/7MeDpG+n7pRkqCDaIELBrKeDWuVpdes60CvAejZcJMtaW15ZDiz+OmI4eE
Ks6BZnImXBhWbGW7kHamnMpjJYS9R8nrY3qZH096hQ6VEtv146N8Uf6K+Bl0OrRM
ejakYotaPCOOwpzkI8fZmLOyZi9BR5Xa78ssjCzkYFMblpEic9VCvqZYyh8OsOGE
eVR8wE7fdaLJQz3A8v1PQlRDKVAzIqDSovhl334qcYbvTypRxrZwQ+bHdXhqSAJ4
8Y8ZsxVh7kHwkUgNzzuguIlpPZzcVpYFt/4S/rA8QOrXAqROXIYoPYoCYyrBd1je
oKRDHa0ltKW1UjxHE/ArsjIMMGN7gGKICrVTYm1qTWpeWD6RcJL0ljr8SI/mK7Cm
19p34H8q0ON10fcHzPKW6EvmXwfCHQ+Zrv5KBRIXATaiNkoJ4I0l4oVifJkykotj
ZnFa1hajzT/JHlP6w39btRFORTqIZeCsAdykLqv08PM8m5CzavzfR4tXdQLqLGCF
RLgdg2vkmBGSyOTSdQHZEKsvJXw3S6SuplkQ0qJlHRsHpju8BD5HIHd2myCZYT9w
1B3RKkaF5heCEbD4zEa1TR2+qcmqknEnYqeyzmvQPHnV8goShS8ROIHqiFe7Pz+C
mpSpoKCmZ8pYxDIe7c2cjyCpMKs63yKXNB5e7lKG/CQ5ZrW0rcVcWOzTgwQExlrv
E0rEf6pYBgaHU8f2yV02Fr8zCj0lFmZYgQLVdiwQrjlXxOE34IxNzTE4gIiHzxVq
nszVk/jMq3JZqqLW3v+Kd7NQL83qcoUgK1eFRbA3UucIwexl53kxABWhm3s91OXK
AIEPEzOTFKggwkyDBnF4VHQx1GKw4dOB6cw/CNFbVmKUiISGZEmLyYqX002+dNDy
HbGCkvDLrxnoX/8cD77H1aX9U2tvWnQ3PqDrSueM9heZ4KVV2skdjxA+rtQ8Ky8y
RnoW2TwxMKPto9QRT8F7kmc8fYQFmi7hehQs7LmndplpzBjp8WFnbTuVjR5Xp4Gl
ZKGVWvHTPL+58SVvVbmKshKLsk81/uJ/n3PcDLf2L8cW+KoY7DQGlLcowr6rxE5P
Ak57ACU4dvpRkd2EpwndCG/XI1twKXnACG+EaE3U2JD3ISjMskbpMmN7adYAyMHP
zRemRDMsGlb+JxOb9A8yLgkMgbdn4GgES0SI0XpxUYjSMz3ShlN6HpjsogsEFI5+
Exqe/veWmGBa0KwZBPfxxtNZE2FzrFLQ7yrRqX9P6Q5Zfohw0CCA3jhYFWVwDAvy
DkrOO5/EuXXCoRYhnGn3M/nxtg/P8t7adnDhdn9r64c898ysys5Zvu+rVianmFQ9
F3hTjNFgihTh0Gd3VxOAPKlUirCT97pX7fuSaQPr6DIDN045S1eS4+mU8qYRFTFT
GsXCeR3eni51lh+6c3w1xgg3PH0eYSBPlSnn3D791QdXHg6/vITx19ZkLPNZ5TNy
PVC+RyMJ+VaFeOxN51pfMRnwMvzHryOnhOT7tqro6PZ5d6k3h8s695mmVsKYM9C8
hU1RnqXZxe1YDI/jAsNFe9cnJA9+dfwsqzlICHrOP7RWyaUyybtjpZabSPGd7aPs
sAXQA7siI+PWx+yG+Ar++j5VOj04LZYqFxauBNxNb3uimpC5cZPtJNT3Pq8gL3Fo
ALyOHN0nnWwwJZJPfV0O/cbMKQ/g0iKXO9x+js1j26BP18sR/+JDDWXJD+zrXZPt
b9ia6A3R+h6uy4s/3XNKT0VE35+okwHQHGtbwGdH3zMZ0DbR9uTe4Cpg0wF+7zQe
9bCocpEg0rSLdwH72hi7JR/4tpJYl8/RAVta38TaXXa94N/6O2uh58hKkkgyyf0a
8DQjWQMoweZM3jy8jf0dFYdkqj4G4og/3s5XNRTMMoxlxiVQajEVivc1BjOjSr1l
ePh9kOTrP9Gn/w2KhDsohBBGbDUMcTYjT378FllRBMN+cwx++u1HR7c0jE5f4y2g
FbGXkPu25TrFn9HXUl/jMpxj+FnT8k5zT44u96Qo9b4ANkYA54Y3UxcJZz1VxYH7
yJJTlP/tmtF/cy3IolRfRRCpIcjeHBWccX7T8yCF/+fmsWtIZWaHRfFoiH4uD3mE
wrNGQHDX/5PNFm2VV3wSw+eucVtjn5GeOStSxSaox9fFpE0l8dkg6+cReQP32uQu
z8wRozOpf/afVkEVnY7DrAyaLl1tAgJFfmqpnOATDRNw6UnqpduMoNhRpL6tAXXP
3mBwfdnxw/bDmzpDh38R1//L03MUXHNvm7Ro6hM3Eqdq4oSM+Kmmsqw14AQClavv
fdQ14tpFv69M6IHk7rdngw6NjVAerGPPNdBRk6+a2pGmNj9Xz1HOjtT0CytLqd5g
1YwFHGg4ZaSHOQR9MC6dPvUJ4fDjJCTRRxHp3KPgF221FRf8wGRvCj3bHXQlVPO2
7wSDKN5uqRRy25CiMSrmwsBphaTRCnfC9Xndk7VgTSRE3gf74vWB9piOvnsELJop
+IoIkzIpSvQGDB98RWLiIzLPDckvgJg+MbJQ2fttJUZdGPb07Q5fBd86qLlQffM+
ZNrQ32+0t+yTjAixgdXvkp00+01sgmLMCQV4vhNDy7mG93tDPTDv7WWDhkIS3xfx
9tn8AzOIpJzna0FPYu+SJ4eHlJ84p8iwKu7PoAnlMD4u7Pr5NhC+mwfwbBfC9myB
LzOKeBUMyTsQbzyf27r2WkWwLESlJR/WV3DSwqG9PU2eP1veiJozOtot2eawSBi4
45FldE0ARzK+8wTrYvrKXXVd3JLyj4SaUUdDKpR2OhaEOaEsnN8T/LlSaJWLrn4/
QENSHioVN/MIUs1zs3mSwSyM/MKInjdsGyusMWpOaUU6RTy0VByn8nkCBkHLYJn/
442G4WiQUedxPw3NNaJ86nb9GmXYaAoX3XWN8eI+nA2exlWWo1bfWST8pROcAASG
BahV5RmB8Fa4yDDoKzR7K2XH3nNaDTiOIGcVIK4h3pqk4K/BqMxNFAWDNnwXQaVU
seUGSs6ycwArHwKhvjJIqu1LHBRV8q0oonMNseL+695T22Ss1i9OPfuLShZ7RrJn
fvUKuj8gQh2S2skkAjNMUWkDeZ+mjgsSGH3cPlakDiyImzkuCPs/Prxv/+8gwDMt
mH9quco1xLm40ZfBrrMKhgHfG79A81PCQ8yYSIGPrXQ1FQ5PfNDamwNSjo2ME6Dz
sretT+MLrLAJHwXoqyyC1D3i/iD9mKs1ZgbqXg64oEyzxhN8ICzedRG+F2A5gX9U
ucrkMp6IsfhFJYHG/To35eIudDjpvQ7J33u4Hep/6JZeLHSJaAYInY3GptydgWZ/
T/U+w6FMXItqxMH+YCjOODVs4uE7HBlUrICG3fB8U3IC8cEzQYV3JReqcWehtf6Y
Jv00uifRsklI13EPNKDWyHmaZBQc0zbm9pazN85vNB4Vbshi/S5xPcDDwsoJXYGq
CkyPNoThnE5FOcmNiz4Ug7AqxZuINytRadpd4EytUAadhqHlgjeHFMxvzSJZQy2q
OVa0icokYsLs9jdadUEipmomiDjhdfMfN3mRDkj9IjOHyHCg4+MdyA6R4cGNuHV5
K7OP7caCUJkbn+qR8voL8JJ+dVDdO/6EXnneJMnqoY0wZpbCPI87MhngzsAEkLdM
mq3XPnr7kXiDlYNWGfkKG7Q8mJzIkhckiKISmYaH6Ze464LjzV1nWBF/eNU9jUu0
Jou6RgLu4R1O1eXCze+Nycc46RtODDrDSJn+Vi2fdnWSJB25g2NDqyR+IHK60D1F
68T2H7zbEg4s8vOBB7GmTGsmShMS6jVx7ttwQfP1MefIcWRk2+zqt2O//wDYTA37
ubE60gAkFl6TorQcUHgY2M+V4lDsPDd5oT8P0ZA2eYZoqdEsrTg5WCyxQ/FHgDWg
2bKIYhJ9T9VB1HheNI3AhkohXu+x4oQHHEg3Uc7GLjKc6M9utuafumTIL8v+R7kH
RX5r1aDetUers7bp4kMkokZ+2QRdpcjo+M0OOeYmaZowN+pbQ6zK6b0Exw4hQTdZ
wlBp5mpdYgw5GVYyl3MEORQJ1zBazXhdwQlXdYiunjednrfe4ypzSEuACrLw6fyQ
BwL5d28jI0Nho+TdN7t6Q4UUYfaQKXiP3Pz8lRYm05ZPWG3FFZ0mAGF32EIdZjom
Em8+4qg9v66Py78N06VtKyoA1aW6USskHWJ5EmATHsc+gMUWStAcyMvwJ7EGrIDz
SONglCdYAZQueDXfAqzU4TPonHJ3Mmo0MaqUW+0W5tHBJwj6PCPXSisIS666Z7Ml
xpTZrQGgPBzA+qis+eXIpVA9bO2XlHYRfNhsGTm1gHZUf2cRogNDANrVZDTgY5HB
4i6TjSAtb4S24Xzg8DHSdLtob0hFp4V351LV+6miY9CIT7HKHIuaxXDymYkJl8T8
bqaJvlI4dPqT8TXuW3Kxl8c7d46NxuBKcTbC7QZLadWR9YYxcSSUDShBETGvDG4h
FAmo2KE2v6K05BEPrEvecFwnr71D+GqWjBcAlWAiyVixtTeU6uMnrNVkVq2z7DN1
525WavuYU+wHHcQVWwuFB2irDDUxP6fGSOn5Db7RMtQL8i499sN9rB1TOxMgXcJs
jgmsRuT+sezrwdwiR67XkK17pUwVTwP9SMsoiNUHuM6sC2Wy5B3WpVxxwu2SdnF5
1KY43wY+N2TKBMT+RTCOSDSO8WMyoXU+V/+OuqC+cLqcnEoYKL5TCqBxFPSrLPdF
fCj82tEj3r2QR3Z5hwVToT6cquVmnD2HZq8nd9iQq+/YBe/WD+hPhW3TRVDVltua
iCKpbfAScGychWzGr/ww8hZRkrlxE7xUv4rsc/nHMTtrEuuAc8hHcCk1+cdjs2Td
/H8VeZIEv3RBxnjeM/Sm0mUntDisLf1XrgvEVJakdQcfCgqI8LwgFFcqGTnMPKnf
MFLi+XHpj1vipcD5PuqcgWSE2okhD6+uf9X64thtYImpS1SH/uyN71eO7oIKUUvR
Wcy7kaJEUO6xmpCxhBJVJq7Hmzw9lnPUD4uUIZZkICmSaZo4EcZxrcUo7Rtnkptg
3PHEZJ5EevHewocWkKNk4OPMKtHJinHR+rTgEBXUytrRPewkCvR1EKfaYkMQsVQR
3U4O8e4rKiqhZ6PxvH9iyWoIX8tT6BJeMWjgVS3GTcTqPQAtGRmH8+f83jdO2+Fx
NvkuTiBjU0FB5o/l5BP0hTOFcQQRhoE1EiFgp57pP+yGpMDF1OBme4PZGqXmeO/9
mBrJ9FYJFFaRom1EE7yzGgEt3+iQVlPJjtnDCVoCmC59r5lyiqEkjk7NjTTtESVO
yGctibE4XJFkuHT5xBnxWY+jGT00QurxQDht/W8zuL+IbQnQ9fU4AMTBrR04Oz0M
LqK+ZCUvrk8k8LG0pzpgbe1R+8D3j+mArxH33KD1p6ILmRZCIaGvPfQrSRkrxibG
eR+00DHiOUD7t5WzuLktVHIYGaQJCesyxaAWsQI1shpj/xAcoJzj6yr55MBP29/X
irQo1hCvIXkrt+nFUnpzmzTGmYgF4nnqlmXoYicgBrcddLm2E9Fz9TlAsB2LtcDc
GBtQ2HcPZ/n7NYO/ws4UgtYVgs/TrbzaLMWGfHKuOX0LEeKq5T2ME8hL8vfMvqNq
3JYsZxOddOD1iSpruzXVJA34syLbf3A1mcILmErc7Mk+S7usUASkIHybIOqi1S/U
vn9NCXbesrVzq7NsIkVwIWk3KsKcK6XmI9DF0QHZ8EUZ3o7epRDgBWXK8O74KtCL
z30CD0Ks1wwNBUwluEFBzrbwJDvpwLOP8vjyOz51LsMJI4XsDYyOpj7fYiBJEm1P
bHzyGn3xy4zAc360zp4rU1wbuioBddWmN/4uO6oMiDWNMUOupZRv62486pKz1AvS
UnZBlGIGpl2orEb9yRHAF3abF2+bBIqHVwr04nkv/kq0Zk0IhLoIrKg7gl/+bY1L
K3JuGPlm/0oxeoBGTxD9LcDLjnZgx/zc8Ho0BWngefTc/u2MGeMEDHVBtkoRF2hc
DFc6+knYPMTrurw/GN84lUARqzcdK0KBDOCtzrUfJGbWXquhcR7WdUn2N5GtDURU
n7Bwy5L5EtxV5xb2fknD1UYpSLIFja8UZHRsIGEjN18bmypYudvaGKVKzA3HJEJL
prQZ8IioKk6AXagtMP7OQKRsnT15czFkE8wJKYESlhdb4PoH7P5Zomz2D87Vlbn6
glkeYlavJrEWQMQDerxQht39n1I2QA8PigONNyvBLha3vnnrO9+KGcxC73o2yQZ7
P69Pn060m604vj924twRKSU63xcBGC3lFNFRh8s4KwSdU5PdYt+4WR/P5xp8y5xi
lf2IgPfkylhvm433exbrPtI9EaEBxDxaU1FtBdV5nzoK/h+t2oaikNy29R9PxGDB
I7U1GKuCMs+1NXrHRHDWXMQknkYFsDEj2e/uwrBHTW7JF+GaF7P9VFO7yHPzekYh
GmM+/U0o78UZWNfqNnj0YNnc6gfK2vghzOZtYjUZELR7IsINtlFsNtZJYKPrUEhC
3SWHYWKWDOLww0p3bpuJIOb7t4RWzNnCQFCGXUjFO+b/PxpAh/xIU7HZ54iBQq3H
GIxdtx9BYfkM92Gx4Saw+ZURL/wENbIbhupvx1XzMB8/170lXu6XCdO0Mk+0B1JG
cQxE+pSmXUkCyfIo+e40sylJzSiUe2vYmh9j089q9uKL/LErKUNS7vkopLgyS07q
bWdmSAD/xY/Kgah07+9g59x64g3+hBe60l1RgKLihRrtDQn2Jz+3bZC7kkjkajfc
x/jhGlZEULzlC3ftj1GSDAfnrJyK6S6pEZ44Aq+zWkj7h2DEW9UJ52eNxYC4VqVB
8w8CzMXxY7mN3vPASYCTUbMU1+QceVAAqXhpBsZQji/ynwRgTCQKE46lJ63a9j+M
nIRDwk3b6rk6unpy4j+zldK62DSqCM5pL9AC3GuLZSVenc31vtzfj+l4RAFHMil4
UjAmLCwLEF+faaRMhJCH+PHZe2uV+lIqT+aJbq4KKTdb9heAKWOKLUet0BJL7OQe
7bjywVtAwA75x8ZQ1lxD6QY1rG5tr6cl8skB5It4W+H/6QzGRZ+D8JFRdQmXwTo4
yNAVMtJaWG7WxIcsVGMT4y/PqeArXa/PMEBDfXX9ExcDbdzIU8vgtOzWOYPhelIm
ex3PkbVpipOSrG0gor4eA7f6AK9cDU0L6zoDP/ILP6EoSS7qy3TvP2QUqFuqI57G
8LAQ72uMxbS5SbXrk+QSjXTNhL0k6KhB/bDKzB10Ji37Ois5/85HDTjz8vjFvHEz
RmYC3Ez35K3zVfbuYgck31oaXLmmZu2Xb9INgekfT4auqIc3FBe1VV9VBHotyH4V
ScdotSP4RirE3pjoYu8FimZvqNyFEzj3YHur2+VT7MxPH7NLPysZs4IICuivmEWs
xNfux6hzBM3iY8/O7yr8e7J40aoFMZOI+LTi4NyPcrNXA6YevXInVOShda+Eyi2U
l06rNpVQW/YTS88F+4+1LUGKWEPIZLLIEmrvP/EmsUWtikAaVJDzY6T7TTOwYc8A
atyumCn8eJNPJ+8nq1/pCk8Z/U8LhQXUFUwnIgt9xNvnQIfkGuyYmftLcg1+YlPV
gzB0F7YMkPVPitTY0qkPqiYWv3g2lMgGPeCYospKzw5R5cyHEv/aeTuVIaL5yKg3
6b5a5ql82/8+L8lxikzowEluLmi0hlj/Brpd34ojoZx1MuT1z0mI0UR0PT0iR+NW
kmZ+18GB/Svy65AgTjsVWa1ej6lJxJVVeD5luil9PpKNJ4emgeXLjEI7Y0nEb8Fy
zHeBeA8a83YOIcHtTk5cbBQeeGJi0nLy5DogAbB9lFgeTRePpPDi6RvM65gNwOvZ
3AU1byVSwAs0BlUKQTxpZmulcT1iStrGJzraTuRWxpircKWAda6j7DffJvQTHHH2
+Rh3HD1K5I+ck4nyKlA83axqxqO95C71rVOpZOdUc8IRyVbDWwdTvxZgDUdELjwN
U2WdufhSznfviQ+KokBToym/W/y4X7yfPa5+syfnvPWEEMOGjuXH4AC1K97lXvRp
RvsXBnXDCUB61ZodGvgIC5E73HzGa+Kt22zcyqHd+ca7xIR8FLz8bN2ILDcwd03Z
yxbYOJiphO57JS3WGXfLlOixfoOzBzQA8L5vzodKbPzJsZd6NwOxWp9Rn87eL/RS
wxDydTR8mO5BWPTvtS8QAoN0giNJBOsHyRpnEq28im/wXphAYB5ZD9pwF0MBLvrA
j7ihmHF1SfRjcRPaW8IwP77QWwyxBx7xnvL+lVo3h4VZsBS8NkE62NWn+Nx9Hyxg
VO1byUin+5OQkptf2l3JmiPxTGkkNLfflFU0+BMwhRhpnYp1vMMBi/vkpqhH1tID
/oF/Iy8tEUiWFAuHSh/U641hWC+Z+KyPqX1dG2FHj4uYPrSnjjijiHfIsXQxFKwQ
UDUfYF66wxKuNPZIlwxdmoznIOPdSnnjVlC1OgEqYO2/R/xRo2XxH8xnPQvNSkCA
eloVbZ8NzIZg4ygwMyq0HZq3xGCohBWJ1Y/apR7PQIzRGJYC6FxfynzAIheqquGs
QGDBFktWbf1EakzyWHVLvsyFKGLlSRNtMU+XtnJx4IpAhB6QWqcU35/x/v3JktDt
OEaZ4y4Id+tYDkH1k5Fd/oC4jyI/jPOiaHtyyhGsvUZhsQKJsChxjL1W92oHJ8kJ
uIBghW1dtaHH0sKxKrX8UHYWbxUhDasyvgT7dyl1UEXWLVwkmOZ9fEcCFbgG1++J
HalJFDQ2+cd9QyNCl3N1dWnb5UdiAJWLJrNkEHfDKAJDRKtBpjvITok//ZvTfG1n
ssMLjlMd8zql1Ap8xGPx1wZQAXTT/6CTy6A+owgb35JPCVcleZdWkTt++GerxfAx
/Z5KBh2zRvYYh9PqXMegPPUGpyPKsKqGTemYirlxtLj4Wx+gZRXADdxMHcvbzrWJ
/X6N2qUYMdIsDejcbPbw6hQ3ycbWUzzTjvtM2hZS7ZQG4RjzOAWq8izAD0dgjhpK
9KIQbWc7VHsxywHwXXIPPKgd8ssLMgXXUJLcePoCYgxW9GmxEeoIxtduPyDp8O22
7uL6J9QR1xuCQTqTN7x4QDxrrHpr491uyvl4KHnFu0TzEFyF9hGeGh4F6Mo1tQcV
T1/u8OYX7YFEGK4Va5M1FS4XgfvNTXxeWuC0rb4ekSGiP0Wdrja68sn+Xyyf5npx
YJuKmohcGVlvPdr71M0CwQ+xECIB6DPLkI83jTvBfnNFdzW9DnKXEcaWaU5Py3lK
VaUbcajgXAJ/OxDR7AyznN/1/J/rDEA2I2ih1Xh+LYfhpY47faPi6k4MfoFAV20m
GcbXdsPxltPNJUHth2uNAoUlwINyeuOnWHcFKzeUHWb9jYBND/ZInQXBfdJbB8B8
WPzosHIyABERC/1kjqbja9O1ZbLJERYQUjirqUx6OheIaZk5OcfN38wEZe3kNIMJ
haLdvC46IblAZtcV32szPHTja1GfdG0/hSCYgS9jkBRNKwUJDqGtsj5tGx5MRvgp
wF+RpF1C2MDLt1nkqYTgGCqKZTIv1U9dfydZnHI0PmZiWKBeWp2oEA8mUP8ndRsy
oTXsSCJwy5vM6PPs+sgFWYiRqbHAezD92thVF74JzCNW2Z7Lmblxu4AeVT+YSj2J
/PfpF6b2kUEqquWUmZsd0dAZlsiGo/iI3wGET898QeaoierTS89lU8tZ6KV2b/4i
gT2ta4pwITAJN6+F5OWnHnSMF5QhVeVi7iL6t5/0hFcNtH8zeqc86+0IDeOcfNjz
SDhM1dUK2k0ZM7XSibSuq+TZYB/6B2jWmqCgxO7o3JbgkfCRC1j5B8oIt1Ov0nSa
gASxUzCRuW0uLSq9QCEsByxM7k1FOYpjJAAcK1WVsXGH/HE3FVoPgA0UG652V/4g
I/+9K0GaPvT/eMHRV1VTzyg1jG7Z7WX0KMheVO+oXcWj1BtvR/jPcfk9WPkeeNJf
200qK2usV5sSJQBNZ6guDF4KGtQjHFl80NW1WIMn1M6/aHLTCpCjP8raKmDwEk/H
JgpLzcSeHgx64wBT8I+qSAgt08azAVwrZzPWvDW25SVK0SoZTMYNYF8E4dMNv3yR
ETtXlSl9LJ/O4pwpUH4GZKzDijuvJraDTF9+wUtfLmaENBhISiSx15qznAGokJTv
YRnMilFOvAAcbVqy9RKFrBnnfXiV7BoSN+tXoOV4nm3sf12UFQFCqxQFPlVqtDNn
V3miDkhNXAB3LQldNWckSOfceo6iLTQqZLcaTM/ISEBIyuyonr4Y476tsO+Y0qF4
dW3F6SA/4dIBFGWjkWGCOHSZbrYhqud8VfJqtuawybEXk5NKqXMEI9BZ6vqz3LNy
OxoUtk67EXlxbAKelid9ynPNaRlpITKyOxJanS7iNIGIqgf8k7B69xk7WMoIXTGL
DoKCsU5fg6/ruxaRto8hPFnh47mbZT+sMblHb0z64hEtVyP/lNvCExIj/4SNcBFb
VwI4TkDcIkjwAM5oznPfAFX4FVybHV9TPNflBSvfavNUSqqI2ln1JmBmQZyQDA9K
ZMk+fqdXcCTPxak+7NQpjL7008Xx/5KswYuDumjQ9cgvpPro4GjWcq72fbID0job
KJqKxAdjERP2csgyVZIonmyKCzfoiHzZtkP4gQmaPs/pGVlOOqDK2Qm9DOuszawP
tkRzylfbUnZaVOz31Vr5R9UnxNHshSglshB5dpIh+5X8MO491o6Fexgt0wwkGgfG
29Bul8sOyRD2l4PfGiMoLHlXO5agSIeY7iIkiqm8KLIXMpY9U+3nvsq3A7e5mm8H
tFHvER+jVHWb5wYFZ+OGUOCxdCNqCEc4p9FkEZu3y0kZhDTyV0arn13B2smE3wZv
cmNZOXtZ46CiawwL6k8+n1TaYjq18QlHHw5egKD2IUGVo3yTadW6sQKqLQ0WjuPK
10v3xWGLf2sHUNi93lzH3xSRk/A+XHueDf9fNTlea8VlenzcjH7hWPFipPvY2WLZ
UDPHh+yjAg5yIC0XlxQvaQAV0Bc+XFxiFvMiekYXkOyTXeAQk5ulM4ZThgjSxZ7d
HOl+l2jNd7SJbglNmab67UfszEyWypdNkFqyCqWvS6DBt6lsx+t8mEop2kVXWzT+
E5jzncKJfMxJjX1vDqb1dzfd/lNzDj0dJLCnjF2mq467oLkznws9BFyUcI8guxqJ
eS+ONYbIDl4XZVFPpCZyzgqItlEAtkZG0wuUYRsMAeFdZVCeiFk9RdzRBJFGgMur
ZNx7AytdYqqQgbxAnfMHbhTkwtxBaxaXt2EGGBxd9KjjQ6eZ1pMXwxBM6e2NUneR
AhLIub8wipK/Aef8TJwkT1k93iQQOKK6+ZpiSzaQNhUpl3I2hww7uBQZNcc6HvWS
ds+AamKC0iYbzSzV66h6piXNQ1mLLddz+54xrkL2wMcAdndnfjEdODrpbqHBWcb3
XaKCg/wfK2b2mPzX8IeyjIii0efpGmAjb9/KoDYGUilt+fFK6SzbwMF+nwiWaS9H
YRbi0od1xTsVuueV1KHfpHz8jaeexPpkyvU8Q6LabJ5OCd2um/0YRtTQFrL6Ai4m
/yNinSKzUlldvJ46w7SEF+C1geIEWU/MI4bx0ZoNgym34N09AlnETDdY+4Usn8Bn
Z0ATmr4XuPj0Acevleaq5vPmn4DQuXbXlNJUaaHO1I1QLI2WRJUZ6RAgHYqEyJqK
n06dLOwH9yfkQ8wCORQHfEcNDyz4+/H7z6HDT4PlNpdmWCG7nQe71Ezq/a13u0w9
41lhv9YxtD0omSjxtFRt2zOnO/iOOWNFYYVwP7msUrNmbAxtCLJVHeAIndBU0dCh
BjXj0Dt8sWGag9wla0X2hIItj2GMNd2wozb1C6wZsVEC26Fzf95+9yj70+VbH6VV
zXntR04KQAzo5vFsYCDVjyXWV9oK/PdAvCDU0lDvw7JINRwy/1qvjn9xkbWxfWNH
miQHJJeEdNdwlNxybtjDFpmbzSbI9Rj3daWv0Rt3G7u6bDUI2H4LOy9PqUlwfLrz
f/aZNnpWigjISRIRx7Xnn8DhPwtvio3llxhccyTeXskY5BeWs1oZUU/Rd1Sl5a2l
GXROF6YGjTnQxRQ6ThAZLWsbgcPPNZdIf7XBcnbvhTvmCRczaUKqpAKPimTcaMgu
0l5vQqhow8rZ3AeMXMF+9vHZ1BWxcMlUVGzWxQ2DCLjHQRyafMQt4JtW2/2txR7F
SkzQLqYEXFqR2yt9GMnK+yvCsWZ2svcm7JCLK5K8cKzjYgIu8mAgjpopFHMdzG3R
IKjoikU+6EP9APJAc7h34ggFwcGXWppbzEeIaR/b5fR4yrYC8oD/gIZoYFQz9Alb
EzZYxLy8kJe5FcmL+TGq5ss7oS6OhDdY7/FF6iKJRPeYGhqUak8Qs3UT12zxIY7c
Epdp3NkAkuCm2e1bpZtx9hhyvN0kfa7kMQjvv8bLatunquBIpNB55KVl7Kq2FCCs
DZZa3jrHcflCvfHMoQIYY2vS/29tKPW4GBcM6xh62Fn7Cwfu1dxjLmyYiWSF/sLv
DSEPHNpBm/raiG2wkrlrrZ3juhmg59911Zg4F+q2AUpDTHUsdteZImjyxUcCBPkJ
clRBRYAdvABUiVGUD3ZCLYlr1wk9+lNj4emMsoc/vXw++NwvIOY6hQwWNCtk1FDv
XNE+kS6nbaYwAt95hXssXhWpo4T8/cl7fIpvvaSEmRQL22ISpA9zhwKFZR7S0DKS
c28iaPOTbUSVc3oEc1H55bSCAYJMCWdjW9NUIihaeSJ/jwTwE34soXxiTDCHM3yW
JeKmSTKRifxQVffY1tFYVeIEWDYEIk3k9xcbRrMkNZ8ApLkLDrbhFfZ6gb1+gp8e
4UEr5QiiG9AFvubxHMsLAEOHmFOuQEc8L7NaozR/96uZNW602k/QYgkD/4rAeBOS
/gXZVGTBMxkITO00waHxKucBQ9B9rwZv4fm30fS6JdJqv25b6xiJRCb5VXs3I3Yq
JqmRotQUtQSxDjozuTFoYsu2BFegIqA72igDSeI29sCcaBa7/NrGDBvlt6uxYyfA
/OtFIXOfV35OdOgxF6avlH78BADiNMEU6bMgGZpyL7u5u4N2YcuDAlU3n/Lpd/mv
Xjd4xtX9wSRTNgzSlfCnjxwkL0uWo4mod5YP1JGXe7tFQ/Fweo3v0zN9vuGvT6qG
aPug/VmykwCmSKthNS7be92qK9TUEE3hjUF3lkpCEWVJPiFUzgFnjxIw3DYBXS7S
MJMKVd0kP4tankFKitEBMahOKGoal7lbqFca3PUvg+OMM9Rz6krUZ2qgpsw2gbM3
vG6+jn8u+pFBeS+a7mthaNtYWu9rMTyq1EYfTpNGP1W0SxlLww4n4eJIvXBhyO0B
UTG2YkSGtnu7Ep4zUryvWA0CQobVV2Q7ZfQHXRHlRTCw/TWFa0GyEksGMosaRVVm
VzVCk3GUy8xdJhWnQEQPCoWwPIVfoRi+ELgaxv43Xf29CNuX/hRElzrjMhKWgzfA
ArtPOYTRCu2xKP7H3rB3ILjxioFj2klaBNya6cCL76lipvboLu3D0TZA533NIeOE
0ohWKGAd0bLo126dCfGcOmr5e1npKw4Iqastz78Qu8q/N7at+EMAj/5cxR+IqIho
Q8nU0QrBMJ41Z1oC7ReNbhfUw+MqC6SqdYqpRso4HOK38ZHaNX2AQP8c0oiXfZsg
cLXHeTTzndsZsUz6a5f+PaGfS+oMEWgdUmZplNh287qrzPK0LzyiEkTulXZ9M7dP
zoDaWWJcYWYUcZTyxchNQ0CX50uWbDfuG5wnlwGHePD37dSfKLCdaJAhnq5X3BzX
2tRQZu99IXAU8u3exBWhgFd3N7rjTZPBcZhrlYJIa47f2BPz+9CE/9rRhvd4FMHZ
QAfrdu2eaz/BNnO9D8789XN6spMxbv64u0g9GR0VUaZ9rBQGZFgKphkJxR2R0bkA
DaWXmQdqrank4qjQ6L6vRM97X+vsM5qFnkegCXKmcZXKNVxVWLK2xwPORPcCHEnw
ZhXfoRpbzaflzQ9MqM7G3kcR9l4kLezW3KObIUjBbarUnAA3xevI3qnHNeBvjnTD
VHvMmU5BEm2+9Y8Ny7UkfkP14o1YAIB0GCszVBlk8pvjPQYGJMdo5hcJZWxV89Ir
jSnC8vYzR4SgMEEyKYmPGEmRcWeg+rWfKBnY0f0gDQDlrurVmFn3d4CVQPIWoDKY
TPGnbbZX/POo3pDWRU5Pqz9CdpqrAuU/BJ/2JINZCyZPLvRoKIJnVY9JdlOICG7z
B+o7eI0PruwriQyxDHAS/ZfCWsBVp5+wdKDEJ+F15EQhrTPnqnk1h3Wcok369Slw
/5OAWse6+SdMJ4+DdbWSXcrPFnqNW+MLPlUPdehPBQlmxRlHhKd3LmTcGav9HEnx
uG2i2mCw/FP+hGJo7Oipc7/tyJW22BUOFnzKohm8lLxg3Uxrok8rcSZ4oZ6YcM4x
roaoPKKwotG/GpTPW6nmhkubF62+ZEltZ4GLq9IOv085i/ppKWszLuIU/Duwxfdz
GtjJbrChWBIHCC9jmMzsnWMPYI+IS9zLQs5UMV/A6xMbHzDurX0ilQezsZ4UN5vm
+6bjOa4/snl2jtkCfTFQoMH4pm4RkYEAMgli6MPZKcejYTfA4BU3VQY1o5wtTb4i
xwEt0MdfxsomXYosqfj898WvdQm9jMWrRctENviULnUmVHsl66lnTDj81PilhXK3
xXB8bl1vN9FtESQ6p0RSmSOsDW8BeW63DFY4kjwHRTktxBALqQDyF48zRSzV4kQl
y9eVt0MnJYNHmL4sSsMU/1mS4D/0GCU8+xQEt+Eg5e0VBUjSbewhTLIW4IT2lLBV
3uckJmO9ECIAxrfX67lRe36uPFs8ttqwPFPscLKqSqIf8xgGL9uGiyYzorvTbEjq
DOlXHGyNkaCDiH/w/0JJ3UFWGlBH3f6CqjkAgvPYk/+Kdoi4bM7gabrlxRei7Hsn
69Gx+poUphyjG9lLocx1Thf0nmnpz5KasMdggEtxuTUwRU9kMqezd4wAMjkUkWSC
kMBagrw5K1H2SE6pe50CWCSJ9J7t8VHTnO7TZfowgGAUKA50fIMYVls58uoyHDAg
kGZVAiGEjWBhO9vGXfBryg0DSH7kFHWNeoAi0ZOKMKxlpp04+ZeXNb9vc5z2ywi5
mb7Ch2EHIPVTxrcrGqbMVGwJInb8x6mvcyEQsFgjpwMPPiukMQ8FZtnxs8VAgu/t
6Y9hyYaGWMujMMLAyOexot+tGNfUMpIRyBIScGXC8VBJysGAVi2KWKnj7WEAZsSw
Gx2bCUg01LXrOQkr0GP4T14JitPUzi3ww09QT2dSLFgGg+R9aCuuzbrLY7J9MdgL
1boJruApMTRQr5Uwsok17jh/RWfZh4ike7beQi6SUvKIuuRx9YLsTUtyhcnClHXV
mxRq9yT5hBWDSSFB+8qWCGWLr2f76vH1EeOjfQfjiPp1EkP5V/6sFqgbRxlsVAHW
/wj1UF+hSuqdLaBSmvvwO1LABOZ9rt1jZ6U8h5tlu3gfQNh077SLIvSgHlfjxf8e
pcHLCA3VGu/LFhHVe1S/1AXYhl57prxRBlm4eoQ26VuHSfz5WCDKk+MYX9n2t5Hc
0amWIcJWtaU0t5jTbuczBi1ZV9k5nDjH0A7WMJEAR6YKOhaWJxRYqrC9bXD92oYy
6Z55yKG9+sn8x2p+hFVJgv5sGg3WaaQ5oH9bWGbnUL2/931MZL6EHTR/bZgYjuZ8
lNaf7KhZSybfnPTyzrJ+6H/MIehVyhSC+hJspBjrqiy3fNbXmgz8S2JNeEzlJSvS
ZW+GIaKZHjo+HsXsucj7fkk1aQAQIIPX6BXrdGUW7AzHOm7FmIiyH22OGXuPbGnL
tRVbuWvoZ3NMQ70U/SXPireEmY4zvPFV62MNV3VUyEESehAfGdZvzr9ENl3SzozL
7xy1xAYjrlPIKsbD99CpgmlE0j3FG1/gaRidjqvV1x02CIc+U0J4XUOziG64a8fT
PJG7NzCHVA9I0H/N5dJjxralEfpJIwiyGHw+XTQCRb25lV6jnHsmTXZp2S/l4PHy
q10rPi6QPiFy0cwWoCQj5Q528vvI+Yys9V4EKSJggL5yE4q5kaYRbpcQNl6c4+n6
95ZJ7nDidcR332yafQok3jHEu51keoPj4/jyJIhol5AKGkEylfuJ3aPdKi614oNH
gxcMFhFb903vRh8UKCN7aYuiqI1aEBUkmcLE5u8Edl9Fs0Qab5KpJZElb6PBt2As
gp9dKHyC72Gu2XV/FKBVAhzn9N6iRROybjGZ3ZKF0caX9fvDKuLJ17xeQMzckMX3
YOLdyZoXSsmpZPo9gf/arbkCmSOwbmN5OjFfaFNhQZMCg3CU3QhyJkOxQoDP0iIw
hihvVX0chgvScS2rYRJ/8+3V7UuIVva5fD3PxDSOE4cf7Uk+ntA6EFK0DqDuoKER
2H3xsIysyGUVLy/dWw1k+BOfaZBqVodzIlKR9GzM6Qi3gdhDsPd6i1N4omnbbtQN
QpWNBG8iw2kNcXLL3D22vBsH/JD2XaqIK/OiJo0KsmX0dPql/JHWBBH1jI7KGmvk
bWJ5jvO56JZr/AZcSGQ+yhaR0yBtyvu51fIQO95UMhtEoONOoDWYxuZZkMsjSVQn
Iwvg36ZIJW/jIc7N61OQg3dayZGbghpq3P+v3gL5YPZq4qLxDweSlkXTaaLCp+0n
`pragma protect end_protected
