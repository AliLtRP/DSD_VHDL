// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:17 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pcKFLC+uVANxABF6Bdllw2AfJJWTIxrWkRn5rOkzvw6GUTb+3W5feHVUEciPAeLN
s33oY+X8dsiTO+xGRw9C2zvXASQeRPN8rJ77Bsf10hF8kdbsPQyrSj2Axp8LjNRU
b5bEr/bgP+t1Hi3ibyXwsOmanOnqnvYzzcXFJ/K1+s0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25664)
FaiQ2RSrKq3M2aZFnU7jWa34uyzqSTJXkl0hPJUU/xdWyB4oz1JEO3AyT6Yp3/YS
NG5vweTmwny8A+xl2DHFT4ESev/E2c5uospsDnc+jYdXZoWhlezNg1q5bwPVtbfH
bqI87i4QvFMzQGEFHwxmy2ADnlBQhFa9CFOD0EFZLeIyIZLW/U3MVmyuL63Ihyaq
7l2DU6tCN1Idi4ZSsuR9bBxObgwm2Ne2YdJ0gKp24DY9HNEJo0UL823xBoe9zgss
KUfEivjNSbvv1N6pvCfekVer9jectvpEJtUTlHIkxaNKpYv0QiyRBLdKKewZYT1Q
hfeBfPjQz9JY5xMBwVVD8+G2uFJRH2J8EmRM8wscOthOx8PexcZ2bsMNvZTR1900
vUipi5BcB71IV4ZFdUlHJujweKhG59tkgIP9RsC0X9eP3S4P0jtfOwNd6JodWRB4
qRGxUGLSH1TMr3fMeyVg0hvW7QQDTMUjKszbOE8N9MlIr61RTuSBXtTWcqhSr8kc
oGnYqd31v8Bl4jjtgTCW1vz+/NNN36DMyOVbsNXVnqM4n9eFyHJOjoPodrln+l0C
Cw9y4HlXdXyIuK5WjofPOF9KJ3YYSzPfjeUuYgu8fRDfLh/K74e0gQivEDWgwsEb
/t9DgI0VqO7gwWmLLgcVV4lB8uVu9c3nxZMG6aZ03wLu4A+DOZRz04OXB1aYE366
PCYjLsvzJWG5LjKzz1a5rUIXXHFg1Tom1aL+Exnxy4rOtw673goDD2pwups3lHk9
270OanN+LzlCxNz1V1ePFHEAq999CLXaiUQCe8BTgStODxNeV8/qHS5DXE5kzF1G
Cc2OVa5/SxoHpKBow2rGxiFDi/kG2jbj7MwES10RqvYc3VAJDCvlKFS0zjV7Vkr+
o8LqCsYdl8lXZZIuXLBF3FMxltCFpby3WNiYWfce4+8B70fLhocyA5Hb0YEmCbfX
Q036/9U2IbBC7XQmxdeKxFM5sarwcMiBSM7CErhdNkSi2wITmr33t0IgYnzbjZAB
UJCyXdWgm4YH46113F+C19E579mmcjpOt7Pz3gHaQPhm9GqmBQuYArmca8FdIe+n
WM0cDP+IC63Qmls7VKwLQ3NsRSyUtJISH4eESFtT5h3tIJu4bod9sAb3jubkt0RQ
0lprnHfl0Qx+iTlVPYS4/UN6InlWi2FRCwmJCWC2yXDaPInw77W1zBjP27LZvlL5
NTRNd2AnvdhorF+u4NLp6rPH7OXiEkWuljULF74jpm/K0ZAoQE8EJ4F2xutp+/oM
cs8tnVlsIml791/I+vMFB6b2+tYeO6TN7qz9M2Y645EEjCnKE78i2bbziFKUX2dy
1HS4bsuHis5HE1xmixnM4DBO3BWUyYh1JPajb1xIG1uK6K3Oc9MbbHGcdX2ohcXW
Jw1kmut0/Ac4o2WDK1hgraVT7vBkl1M4JFeG3MdY0HzFMY2KG/6cGtbV7CruN1kF
prZS7M5V8gjOuvYC7X3ShtRNAjyxef6oLjD1Vqa2qaRxPi5RnrFVLrDNDHCxlr1Z
wrASfAK5YQ2r3XG7069pe+5QKnmLUwQjBFxmSiGygJZut+4GSnveLF2AqpbfL/Tv
S1fTiB3U1O0zAhddd/YgE9bbALGko5TsxuUw+NiC3d/Kd9Iba/tEKFYjIPhiOUwW
knV4BvFm4KobTyrLny7PAvud2efoDPPaciz0I5Ig415WLB3Dxqv8agpPpnm+yd8l
nQj7D92UJ5ETfhxjovuJqS5T8TTJPpcH3pTyU8wVbuhbu12Uhzg7a5Fjadh7CsWy
lQP/cqmlRcDfMRAhMk0X7g/T/cpTpC9bqzofu3T9Ktbvs23cGY4FzYyYpGgCtODY
9QlYcB0pK+YnaEfk5C1NBb2AEWcEg/KOpO9Za+Hc1qqSSkbIEtF5sDZ7HsTPL0Dy
zvl0BZmyBkZaiGHDdfKsGyveeMjLGQSy2qkq7VY183GL5CdI8wvZAdovYFhI48jL
4XkpR073fxPIx88L53GUCgVAAp+R5CgPIcBU+tNSBNA9eQJoqHbY/ZWZPgbiC/TV
07tMs1GDlezti6uOOY1oSUZ4lsVwEUEAqN17XdCMzrJJbCAiFc8syBxNxMTAYbaR
BIM5Z3wcmxp6qGuhaQeeeWoX0gJofOc2nuTjaIfvh5oxC5BpFbZAUOcK+qokwnk+
+hpqucLWTriDt+WJZttozc1KUJIZ/JeJpRmZJDFk++xLUxL2FwNMjw07qB+MxOoL
hYsrEUfVC8BH3Eo5bKcswp0I3XrskfcR4mL1sAqK0fvC+OjaqhSgR99OfNz4pzvf
BPP7vE2xK+j7h0wwVWpIz1bzauoO5cbXL9dyJTFJcaisAm4YKFwDNvEPQCQs5tBl
fTU6vgbcMEPiw0r7cD53w3Lt2hXzoaCZRkpcDR5HQfm7NPqRd8D8zOpujRyuMG9R
t2BBzUkmiEFghRU18635Yfk20rb6XXQpmKVRNdBbXuK40GiKXfkseIvNbVSIsTli
LSl+MwMvvDwSshp2rU9NSbQL36vaF+CMvzjeqWslZ4asIaynaJLFsfo7OQ8vXNE7
YBtLMHd/4y85F6uhBykIsQHynE2dt8M7/e8sxcl9Dd3dnrwR9lKzO9rijvChwfT4
cUeZRY0pWJ6gWJbXHcI1c2L7pz0LR9VPyufVWIR7rPCMfjNAUhINQWE+Bx0HVqN1
X78zYnnoAcEUkXzrlClk01KQ1Nknip/QrmMTMrGm+qoA//2+kXObbvHFEBGbboSH
1/DGsLidwTw+9vn/zO0oJR9ZrWmubg3wYcf+GOYD4znc1bqsJt1qMJsy/RRNqtjc
OrxAkp0O/SM2LbS4iVdarDDgo44879Ejz+Xj5/i4P2J8up/G5DL3lDZ3EwimLrUB
hipYjVD6h7ToGjURn5T1JDCIGQJQE2tcq0S3dv9AT5MfzU5plN1Sgre0eE7Lr2s9
zC0czXMqU8gO1pWuHDe0tUlPOBJQh+MzMAA4kFgFeqVf2Z8Oyxjnp5j3L5lNNedf
3EtMoA6C/DgESzl2Jtgj58p9gEeEe9W+9rTdNGql2aFVYxIfRVuPBAxlO3TLzkwr
1m77yaAc17sv+G7lCj5IJk3ml2fo7ntX7hl1yetL1lIWmjnPgYyhrZC1Ls9RxXUo
vKrbwlAI5DdBeOwwIvgHzTjUr78So4FoZmLefpz3TVpQIYSm0E3T6ZV9cStH4x5h
mKfSjHiwa2b5h/ShDRg80E7C6JZCqH8kmDkxtE0pSsu9vkwIvqWKLWYgkLDCE0a6
Dmu0PQk/HnTgYb0DqcyarwNCZOsMje593nmXb67G497vgUyyquQrZR7j7xEzpR3q
WeSYR0g1/KugKYhG6OUuFKDOK4ACflEfEUu+96z1SyCkcKTdecNgu4iL/e4IIRkR
/8Q6bGWOD7wMUXZTsZ7zH7T3dlofbCvtGHmsr14f1fTMQpk4vm3bo5gecn88hlV+
IyVithdbf4OYz4h+0EWn7bSuTlBDfROAHbSywHHZEHUC+nAxXXeuIHjUXEMAmtO0
Ok5+98XESL8iZT5NtFsLYONTBWkBGr6Cq0lctBQwc0seBzwhz3mmIefm0h63AB2o
jJLhn5z9Nz73gxpUOJyKnkY8rjwe4ni1oiFjktKlkA+pnvqajTT33eUuGQ3iIuJv
zOdfdk/xKj0G6DhLQZhDy4Ywc0KO4eEidcMul4vZq3ALaDcHGwut1GOIoPjEtTFg
cKy3o68yQgAgR9ZnXZswyncUAne9+o5rjvoZQ77ntN91gR0Lw1aIJbMab/T5lxIY
3mZkKDPrVqfjWl3DWc/9MrQlQaOqHWwT+06MIawdjViEucemGaiG9AYuZF4YG+KC
pANkvqMqGAnzh3e5StWMled9DjeV1DGV97AcQAw7JEu4J/2OAlSU2ZXRyA1IChd0
yoyG9217c1e4qBTWCiyXG2mc7Gdt1P/Heo9kalIK0/VV/dQvK9dpdhqijKHG5ZtQ
+ZrlmAS0VNjCaCbSPMjhWNRJ51qxAOzskixYBYLGYCqxGYOJxfV7VllXyqUcEQoY
dpQYN147aV7OYfeu4oBgrJSqJtLLV8/RWP67HS5f3HJdhvVD2qxRMxvINi0OQZno
O2pvivGA1KV7cgmx+17nN8uYJDekqiMUuX2qSpkwfl29PjmfVLBS+AaWnioI2PqO
WV84pY250oj3H7PedYcuBL24e7dByyjsymzwR7inpePn8pBq3TeMEnUuJ6dvNyk6
ZnRkMBPVpjt8FOEnaI5hi9TfRmfYDSy6LqeyMz52/HN6qLSxaUxg8K55xCJud6xH
Kb6t3nXLENsHfp7qakP6h+kAYFAsweYD2lr5DZM3b88Y6GDGAVh9Jfo2HFGLfQy+
Gl7AK9UFmkSW+Kqmjzmc7yVgPTIaGiMzL4qI4VyrZu3l8/YCiUDxaUbGK4dA9WkG
MBUdqtCrQPIaJ+NJ++ukC5CORsF5LA3m7kvgzID3Jh46l9r5kIXewhipKUkb4cCD
z7ugxnHoVUl+urJsOGAyM9lIexk+h+OoNcnefV7SC7VdH8h61aWhDzxkMg4CKc3d
79o/ARSDn4UHA14AexnnklBelLTwyC8thLA70eV+r24j5GjomLQ0rFbBy/wrwues
mLPWnhx8yXEBqDhscJ8U8pxPm9VuVxmv3tVtoyhO97V63WYprR8IqW/WnrNPzdbg
6qwyEFoVQfcdyQ0w7hAMjO8SNuZhAIEsG2BKiJZW/lrG2f9/N7e6MEaelDeD0VVK
S8+RF0jqxN2ZME0Ii3teqC/WVXJzqtKyckEEmHAHWAnbeQxBYpTHJ18ArL4MZY3w
gaNSA6+GDsPUNendSE/iEVt6ZBAV52rPBURyOxWvHXNh4s1IW49gc9kllUMU99ik
6Pmd4ppncodkKzwy+NwIZiQZ8oOi/0aI3YEePKLZ9btXklwXHljUVO9/DSyBZ+5/
eCcKClAorVOOdcyfIAZ7qFt580qPuqGKNsCIAeoanpflDBQxRtCSE9RCRmCvFJHC
JUq32jWhpC9nc2rbSekuYhDO8ZRgFqXnFi9HWJqzU1mKBqIXuY4rNdK9i7ZLDVNs
qgQaH4Ua7lKKzH/cxP+COPyM3xbORLFfIMmRWw9ZnvKnJhJHXR9eD3suBP0dA32z
HGVY9rD4F6arVN+VEVsdL4Uq3jgvDgJJLJwC0d7A+ZGOXr5RQ+PxPPbC0b+aW4zz
BnxKdb/0X4Ajh/P2bPGMinKM+UnHxNoH3dJgwIMsTGseONZm6x8xmuO39TDwbiY4
70C0848BrK4uoIENq4pT5slCQubx/payeYCqNwU+4spFy/FZBXiGtUF2oUvO+fCu
FHSIu5UT+12SdFIqGLeYNN/8ddeyRL/s6ov3q3OP99/BJcwMoI7LaM15k2Rp4TQo
cOpYoLFrsp2n8NUduTCfcYY6OI18bkDcXX6oGeLgzsvsCrSnqWNhsCab5h/rm8xT
nsUTsJUHi2VJeQHDhuxq7YcOWAK1RAkCr14RQmZwmGSR77O67SGLDhcbCndfID60
iNzEu9L5TURYSKRS1dI5LpXQrQ7Eq6V/i5y9JJxHdEjVa9pMUGOzXzxchZYwglQe
ez+0COjimOF3YJXMCP9Rc7nKYV4ihFt5oLUMHwMiCgxcY+QvhBCAqJ9Rjp+HynX3
PgGh+9/H2rYotIVPnXRye3GCOWXvUC5CRmGiDGOopPqxJrNxSOYpqH1+OQ3/gIjF
BwBVRZO9mLL/tYBgn4GPd3zhiry6KAmciPYJbri5vueUaEAysNF09Fy1VObg1CrS
baGoqoBVwOhoZvgaKnn+uuilRNOX63VHYNizu8XhoWL9L0cDmWnxxXJ4VinVeMCw
nOuyLzYXve+Sqi7u31lh47flTbUmKSTgoTwAWxDSaV/lq7fZGW7L+b7nBeFJDbft
+86P3f8q+mJpw/DLZ6ZXirNelHDq/Ohlv2StfVZEm8MMInw7ZVC+WZJvPBvGtP0/
zDfru0r4i4butaNYHzDk0QCg1TeiK1q1vFBTYKGyd6KCxa4VwPk8t209aVpmEr9b
SI0xNHOTblXX4cLoRNF2o5r79KklnGuacXoRFimMyuFmdA6PsBmqbTsyrglTSvzv
aFj+nL0Ecn2qPQ6UpsZUiupFzRCyVHxSBf3C2TIYo6Qd4VRmouZOF+vDSaOvtNB4
Fee2Ip569MYx35/39Uj8u6mP44saRg9RxBbxZBo6COBCBeVC5opJlA4+EQfcpoCQ
dhvxLKCb6aHf2zs4wgu2DGb/9oroFmhRQtFHfHcQ3SIbtt4oNRe6padA4uGCK7B1
YbbBZrmvRzdVYulopJ/7HSDkgcshZsRbG/bnT4UfaaU2ksZdZZFDeuQuukS+UG5o
mTEgKa+YC1hi18EXK9LufqP40UdTL18aVpLafRa58dx0y9kdLhBIXAuPkXt21dpD
VK5xehCt9tZS5xJMv8bBAZctCDNxn292zGVcqExH89+nQpKT2TFLkxvujDgPzvUM
vqRo/2czCLQvfp7O87bZdW+ql57MG8evwFvB0ZdVQKIwQE04RuGXnOR5ImT5gOOj
zUWLOc06cEByPXMO05wzgotZDzLrF+Vytq3W5GVUK/TPnDL0aPgUE70ulFFzNvUd
LFczXb0P5/7hVfh2fAjQXcs8IWaabdim9RGgCI+ALnOLdRdjB2mWrltTSiPdNBzQ
Sj2YSv3tov26ZipPSuOGzREEi8mcsfQ2yOg0t12FPeFtyZQSo70Q/hJPUdyusbnV
WpSHus3hSSQQIa7h+nF1FVIzgoGvHmbdixyUHpcHVzost1DttGNbgDlKn0zLjUtQ
gK3FIMH7UH/8SF8FBjAzb/cwS6/lF9o7tYzQCrPlSfuIZrhY6BezaSvt1unXoDe8
WUWRZKkccs8QRQ68z+H0GEy5nqOCfmN6Uk8aTcYIWpnh/AXyrK+tcdPdbXeepDd7
LECr0K7/aoU7sqgrsvnDsssMuejd+jdzQY1xmenqVvV9n+SFZlE2xNf5KMxNFZ4L
AKLs7tSnUu77oVH9tpXyx0pGCPO19gQvropgJEeDEbvyawEn8XBhYyjaUreUkv5h
jFlmED+bbCi6XRLaA81Y4978oZ9SBNQdWy30xKgpc/Og7ikDDNZJiiWBLhmAwts4
M8HrNVp+CQw7iZNFyj+ZHlROSGESq4b07t0e0f350zCa5XPtSYhMEkdJBn1Dnf04
2l7FNnS0fqfxnM54561UtV6Vt9djy3/6L+CCNZnbndHGkVr2DLzxT31YS3GpsD6r
t3WCkuQ9F61gZZDfLH5TETNZ5H5Tz+RJ4wS676CssiBrA7iRLRZJHcuot+8z7Wzi
DDS3GedmJMP51goIJjiVcljikNogSzf/W0gM5vgsITKwl+Vuxei5doDvvpbIB4ea
dxOa2NBq/UNIdFtHvvRSs0ngWs7LKDWQE6vxOB+OwfcUuxZoWaYVoEn6hSt90eWa
l9vdzS9PoklK25LZ+VexFN8fd83M9f6fcGuqlUtBabkhjuMkXsAVPz7b9JDkgaGV
pR14UORh84OqIhyIRXkVHPDTBiC62IcgJBygF1Ffv4gzPnUKQYjIPfd7GddeQuNM
nuNMBpf0PZuv3iuvApyrM3/7cOJYvx3ec4RLqNecavqMEJKaPJLSjin2afCJpT94
fv2aPzfbpJaigsBHKI4T54Zj2V8+gu4cqO4n1waLsYQpW2CdQvepDOqyuRXPK1+L
cg2HZTBXym+Vz8ePzM1TQ8JiUCaTZjOhIUBmyzUOLX5b3SaJCXUbEFF4BLup1XV1
Dl1n60daM5alw8VmafzpuwTPuCnf11Sde658oTCK2fPQHBs1QveTxGpXz8WVWDRS
4Pt8Qjb7x2z7K9At6hrDz4UDPKCN5cT7L2MLShSgAnLTaN3HVe2nHCJfq5g+tPgq
FKyBFa1uq5XQhyd6foGQrgHXyKwJU10OtksvzpKbC6I0EdTlod7nNIXgtQxfe1Xa
ZBIGV7lNJfwZbkEz9zIOX2+D7qq4A45UTjJn0rTt+ujgIpoQamSdG/p2NJ6XN5aY
O3WjpoaExuUQmAwPAWlgud5BvqWz+3zHemr/GX0QIQBzuoeakJOEgtKlUpPdQ+jF
AxIlKpUoLCKF39yFAJjfwOCxwq43wPFyFjwVSK+LdK4KaoY3KiM3u5Yi+t9ZKNiC
Mgl2krjvWvv/Wr1kpulXB5w4h5lRPIZOC+fGJ/17fjlTaUHgFY0frYeOdvK1czKi
jiKj/9PANuOquO1gjLbq6m3HlzS4556U5dz8m2JrXv27BBgAVPpWD2RaqfhcxkHx
sw+B1EyNMKi/nodIS8iqr6iWbeaSrNuZBAWssxEnRWzdU7wAjLewLMFfaLGiwZmv
W01iOrlgmDN2R84NS4NlxKHA2puyuQr+6PPuKa9K2SpHo9joGm4VTL3p2jUiBYJD
HPGkxKKg7d0icmzLXLS9ilSz/BqW/ssAMXlFfc3d3PYgODKpupZUTn9voxGWIt5f
cQfzQBcDjNvBST7RhY+VxyRVTbsBOU7Oa9xsrRXYY8u+xDW7+GXOmzuSrXlzaFjG
mpgsCmu/e3gwrNAAizXT4YRCY9uq+gHFh29OraMbS7APKsWYCTuNK4bJpjs1qbKT
DFE8ktD3zdTXtyG2K4r3zQmIQBvuj5kEdVjpgv1ZBdHrh7aZFafVkQERaR2vMqTz
Cap1v18h9YhRMIXxFogPZ3U1X+2Hk+patw9SsQi5u0Zbse988PnWshi6FbARWrwG
LGAyw+to/PaOjug8Prcmor/PvF+xVzdM0LfEYqbmWFrT9TC2kIbNem5SxUqZEMNB
pqk2hrU/nV9/1Q9IAZAf0nB1OPpl+AxjcA8DTRRyfMUxk+kqKANNINwAJT7jgwTV
KgKG+QcrI87WWaZ0dzXZ6sgvJW+R0qQ3UgmWFMqpkWYfokiYNF3q/7ftO41GqHsX
RZ3LrHjZ/D+CvpZwm7y+nK9H+06ifJ3mXMHmoTzSFVisf6xkc3RFyQHSsBIAOG3l
TgttevgMVIL3HjwlE9TmOXZ9ScbPF4PC9hDmE/hjfHWAraXTVk47OnMOKPy/pJA0
6+effBAgI3CqB9FhOrtmIuVKshmOdW9V4ztO1mjTdtW0gtyz1trxH6KXj+/T1ixW
ox4HKQtMqMJgj5fKfF1fVLzlM9bHLrM+g6xgcjuzFrV457JW1iQVfJrDr47VxFxF
u61qsC83pcO8505pBVIbnlDtidzwnqNMraHKIZZ9Rh9iNfm+CaRx0/0URHzrHq0+
LwauBwRfED8Oohy3qTzdJSRdlikQZTg1DFa3WQMla6DGeP4GjIC2/ycNLLTATWT0
mK3l855cHNAGMhKL3rrQH5AW5FIoYSVju2Ez3pVxkop7NSfWQEGmxal6t2Z0/a7D
fAoQl2bx/wa3d2pTIfac2S74remRfCI70uwmJ/xi0B2flvHThOvs7V6//rrLg+jm
u/WWPeT5rDkJvAkQA7v88/JWVaYaH6lziaLFSWrV7vzFZZ8XdiRp4eapP3kg4H2v
gLhpdx2L9mSygr1SwwhZpAE+Fsc4NvQnYIH07uoI4f4dF8AzgLi2p7P3LZ3QOrLQ
i96hebpYk6oC4Cm4j3MtpdwiWrWbzDn+6/n91APj3dr7iUAb8Nhzm3zePVwKrveS
RW01bDbwQLMVKhIkLY1gUn4WoZN1gXAKHBnGg6Kxuuj2RhDK0FM4RKt6CQljsQwm
KWSsja4xo9cfW/N+3nXUC9SvHT9o75JiTS0QulPzdJW/zJf4PHnvFVg00w5dGAxh
ZWt2wn+gy5J3kTbU0kcdzOYigjz0BFPipGDTC4nZhArA/w7yRTDiI6nizlV2imBH
b9uOA8acmi7piLKi2M0R/SguNT/7lJBkc5FVcDTtryjGHHNUFMJ8pkgfwtjpbZwW
TrLoN+v8Lk6ih2pvehkNTmL+9DMFY7OF5/UZDPEB60qyFh41p3u7J2Ir0Auv0iJ2
5KQUDKmdZ0PQFR/bNjD7Ei3eT/wewK/VimWPpGQzNeg655fywfFnhsUijScej5Yv
Tu1doLglH42HL2kyk3ezrYoWZPlXWX65jQQXqPQVapWF1x59JO6VjBCG1Uw30Cg6
9TmnSV1boKF5jmSCRmk+Mky1ttnVjwDWh+2ekqWuiR7Nj9f25DmBGgLIEPnikFvL
qFNnHI7IZvB9IY2a5uQi5XCGYZJYnPHW3XtHn0JVpBffpJGoaUlf1D1Q+zQeOsH3
tpLl3DBlHVFC50X7dPZklW72KdocIN3SbAVuhUn3CSOCRzqKJJKvfklWMEvO9ynF
Aiqg6KExZpddsl+OmwR63d6OFRPalFG0LBt4MrW0SRQS3hHIHb5tD7oxcHhO4hO9
CYK+mPlF5qyopJrEEVBsAUqENBcj68rYPq5q1gKnj3xPKUEK9fvunFWt0OH1Ylkx
15m5SztrqCFAFkDEafbJue+6SRsg0BcpaUHFE1wjUG0VnzD+E7jWtrexUOqiERtO
bN1/PmghZgBwD+xjoXTX5a4JOG9liBg3fGXFkZ6aC/uOjq6oJNz2/rmfxSd+LZQc
oAMqEKmxzhQHQh7n0LTLO6rawaWuC9laXTQvd4Q/G0jNojMtm8KdRJ/UF/bas/7C
EISRkerkkLOcjyzvGskpGYucQjeTEBl3MVabG5tcZznEwEVR6+aCDQkWPhP3R5SB
x1frKcwCUk9wWarFeRE6o+XYzMJOft+37sfmWCwrmNArV8eNIzVCaOCnEIZFqdIz
VRBjlFK7jku8okFJj1UC9I10CHyGaavnVAdEJPGLfjkaXUl+I4JjNTDfoujkdmm1
P1beeUfJqSuE4/D464s6TGxK8D0pbgfU7Cnxdes30kkRNAqCmzc0qrhi3kBl6XKs
4NN1paOyGjFr4mzj7fRoCXGG/SvNgCSr24fgUIPQsVSrESYdN2/USp21KGb+8dIm
tTIkEfYJqN4JgGAweUpi/YSTGXFiWNoAFzoUSiczK/sqHXpiBr4U7d7XnJrWGf5m
xSdu+sZBNCllrBoaqshqaLgSaiNQqNdrndw+iFk2GsT8LDHG/TFK65RXNAAbcEzD
/fcumCIbz4ac0cUMp4Hc5vLVMUpPtZJuIAg38gb2mLZbow3ikS0sh6z0XuUGWyjX
2rWC941VzDSqZfQBnJJgUHOea5epz16M8NyGpJ5jjaJP86WbRJzVGlHB7Fjp0nW9
fBj90wEddrGPz0SxJ5jWthHnHMXh7ZpL3QXV3HQW5iDivf7gx7n5Zka3X5jaylJI
6pdd3qizSqBjlP/BJIWtJrFv0/8IvOjZnu/71mjeb4FTf5s31lon9fHGNMHHLHpg
sbswzDpc6oh8GkJHVGz9GDs9w/4i+6/J9th6vpPzR93ZFkEjRTrAixWrMeQphN82
96anI5fWY0fXkmTjNxYcvb0somlpDrSHJNnRMqYpKT0U1ZteKxSY1GvLdmizLtuL
pmBDrgoYGzH8dRaFEOKJpx9ZdDYHWj30Zao8a27tyUQSrRS5kH9r9lT2oC4IbEk3
fTlkbOQ3HuOR4hvPHx7mbce/yS1FkOIi8gDDaBj+yE0xct+yqs8lxrLxZ5236M0c
tcoiO9lkWJGFUgMIRf5vlkWMYU6SIs9FkKc4kXyw4nwqbvXG0oZjDaFNEhLfdFVS
Fta3F363YMf9UPK1Vi576XGxoJBGNXzk5ifDv0OvIkG8YPpF2dPacArDZYANbTHr
eIzrv3zn6o/ZBiwh2yHb2shR5w3h1hjGQgR5vhL2aiV0Vh/3q99pc6pyJ3M1M3+V
U5dwyKjWvKWm2Aw9iuafjQwPTgDmOajb0i3b4O4dp0DRVSSLaWPlQNSVGyvTJncH
vkFDpJ2ZxqsBOUN7lxnK9+cybsdQmoqwcf+z+H5UM+gNK+puYOtGREePNDhXBuFa
xFbwz/VzLx8tTz65rECUmhdFBp/5OYpdSHVTwGblow0vASZauEg6mGtfA2whYT9H
hvbvNbwCOt5JMDTl9TGZR2tZjA6ga2eqik41Hli2XjWFLDp6g7aO8z0kId5q9SqK
O3/wbCBGYigsF8fsGTVNIuBRyPPn5itvMpgoUCn62UMh7rAOix2okdP4nlI/W1ya
1PV95l1T98/AEIKeTyhPA9FGmlyFc28aAT96Ie+ZjsFgRX4eqTbFu3mizUOY9H8b
Rw+RHKsDgH4+XF9zW/kpPm4XDDdr3c8vu/uHNp4yEDRm1PY/1P6EtoPj76AxwmuP
b/qutuW35i+Nn1JBMMaPDssOD+laB9md0jPe80aHa1EY4lJn8XucADqdwFWQWPeG
fVgOd7CEQo/v03yaanBvblhtIJrx/a/1jgZc3NiPQaicd3aolmaDAMOMu03eLF7G
iECL09unwGE1xZo6QHWdTK4OsDb7vMaZ6NUwwHLrTQyUhSGEg7Z9ECJdfnaS35hj
WeW7KzYFbmcEH+Z+6OSYtCI43h9aXJwl34iFgWHmeWu5rmvaHEzm97xTcipYh/fA
JRwzUt1ZUjjubBLrNvtPfQZy9swJS9g+XA8WaPYt2p8AXnuoyE3tvAx64wNYpyUl
glEubFI9HvLOA4klrsIfjO845h54W8pHCyqipEaVGlbd1UR/tcPtZcPL6pePwoMU
/eif8DNkNXlZdT6nnOSFsRrf+wo7t5HKc8ecplqmGJTfozCDMhWJxRs4uttjVILr
jGxxSQlMuvr8ABetDxMuS1ORRvGGWHOqImAzmNVUd+sPsfddX929Ecabcj3zfv8s
8U29AJAdiW/JRve3PG470SJVqS7IzQrIww587P8+CFFHza5+usfP0XgeCfLE67um
lc6H/gXy9RdtGOM5qs5gzK5OV0k6bPqlDSj6+m6uvJ2/CcNYGztdgCbYLh7su0e/
saTR15gcyUDmEUS83Tc45/3H97qB8gneSqwQ01K+OCgOIZDzMvyihvIk3v0YzEHA
0svNqfIZ3+PBUsnmn7S4NvwPQlSMI757t2fBKPEKNl816GRZvaatDflClcXtaO//
4UqAl4/kXuZxtqBZuXOYbxyltAfl7s7LfUeKWFY0NObJOO/+nbz1GYXhNVknChml
SwGGaU3r6v9wRmnnttbrTTYxwucDf/zkVWQ+YZfxOI+KXjib4Poq5PqXcCQ+U7yh
ZAOksu9c63Xikm4ILcEmiy+PsMWHngnACW6Q81mhKFpPrD3M8iAFkuCyFrFFTUwe
PIHcSbtgcBDydm5wUvDoyYTM6pCmj4HWWA/itrGi2ZxsVm4Hjw+N3+jJ5S5uixnl
giECMw1oVs7TbqD+9fCB5bAjWvjnAZz6hk2iBCbpadnJqNqjaFWSGve/3NSkzs7L
os1oQOq6COb6F8ChPL4UX4s8zGzRtoJhETc4Bxq8oVOlJjndK2CnxlestXEqJQ2F
10H3BZkbrhXZvTQgEsbkfFmlsmfvHMyo7kZfR1Ss9DtCZD0KyyUrTup7VFDr+wgU
1xKi05LdzcRogREcEO1l5x4dq4Y3rWBqw4iIx4uZGVk9dRh9nepjM3bJA6m6BhGS
dGpBOa+W2c5250+flAqSrQ1sn5Jt4Ww61vY/rwFDVM+DO1TwwlOjk+cIBd35uv+q
9E9VzZokIgioLNbqgTlFqjxo16YMr3+4cH4rsLqn+KBIFwt1lL8RILV6Wc61zRXg
WXc7MfTUu1OemOttll9hTM567i+K8pDjZoWCtoAGRcVfFVeRIWmr7S28HdeMSB+O
/HCfnOHTaLNv+lPozyhAubNjxx+rwmd7OgzQY133sd58CgXF9tT608V7oO5y1Alg
zr+NcjBsrKTuWR0uNTRBmX+QOf+gyr1J9rETFGp2JJ7WsfpZfhASkxUC0Q2OsR5A
dlRr88ODZgQpZp4H1AhE+jS0ze0a2tedjF8exDcu5ACA5safnLB7vB40c4GOojG/
y48YWlsPbDthDDiJB/1U70xI9hfqYAJac/XanrgqOvhpq1RumelIrNhQckKSsc9g
iSzC616tSvT6pI/O3BzUfBCpYhYMy2+gHNU1P3ae5YPw98gPnSzmEEnDpTjtcpnQ
15NxUnpv7QYh9B2F8fYV0JRdkJhxJwFr2AauKUfkf3Jk6As0lXwVPN+5g9HM/Ggz
3nzMnmVQAvs/HKDvKKoXECEo3vw5HK9IO0cF76OaytEsNZYoVpMWNUGyqKz1iMS3
Ep3y4f+n/5lOWoh5quUEV8z7cBorRDT2DCRXqqiDcej0oVWqMjtdVgZNM/jZKOr1
3WvuyrWP2sLUrvCkpCAmvNirgQgAhossZBr5ui2cEGJUYJxr66qBTtBO9IKsYLQE
PuD2R2BLr3yTgXjbZgeoRpHXSeWDGjUqgVD4BMZzdcPfpZl7z+WNirnX/dZKI9bA
bzB26+6k8qdeZCRHcZjfQiG4UP++s3QjuPg6Wnwp85DMVZv6FzZDrEP5rkbasGdk
ZNn0Tvw8E5JjHsolfLqNBh5SJuQWMPtQj4EjEllP7TNo7Fggt5lWLwVw1Ko0BKCJ
XKPQMzXj0rjm05vNLIO2g5DRw52HHdttZTqY7H64y99KFYVmwz1o8RFCq7bHWDkX
vZiFEgzGHoG1YVtJFrauS5qg9puWrYH1OCAm0n8WHQcF/Hg+Y1FxnyjfLdsBter3
dTB/4Qzk0rH5pgf1rCK4MkfVabcPZYGTJz1PdRJd3SQ0EgK0nx/Hkl9n3uaEaTp3
T/t3fgJjr7VnaDm1+nC921GnmYiXLyq911E0pjm9GjmBggRX4+A+PNUTRPR59kyW
pIPvCjBQ7AErzhWfAGsuRozkxGgBWwfkOUahzZ+vxkQ7LJdHp5hPi9FbzAdtUXpK
LirMgQd1EaxQQ8t2ZXCOY2lVDkZDapGcYrT9u1SA4RStJtUyXaa81ozN8MayJl4U
ZMa3suTCHGWusJaR5lJ2HtdcNPJWOTJRzkEhj/BgpCSAArGpfc7CsCz9kOV+wtjp
XNuCVWcM5z4E8potthM5hmGMDePu3LlpatKcugebpJuLFI4OStdlndSy64kO8vKw
srpD0znbXh4Atn92w8fmUL6onqpa9Y1cIwKLHB0er/W6iN411cfYY97yJBWQcaB3
RpkYXOWkGcVAqzOc3mmjhHz+0//37Am8vmYaC+JudwOulmivcrDepk+DyqAI+m6o
mXBqlwawO2hylr4qEinQ/FbGOn9ea57BszV9Etfes4aKgKjQr2tiByIaUo7vAb9P
RCuWU6v8Ze5v1MX6Y35kPfGT9qJu7AA5vzJFwrs/+O2z2YWVW8utWnEoLVsXabNL
RLR0HDDp5QuxKYp4k/oskeEUzdEsdzGyv8rEtzmYNzXHl7d/QvG+T40m2xVm9JhG
UINhf3XjTkSmj7LDfiYgVJ2YHX1gPfhcqhfO6kjxd2Q3nsqgcvxXXBanGIthGup0
3lrkwMdBijul3fiTXbJJOK8/UxxwsmSmnPSSO27iIaiqc6Fw1qnBi+UznJr3G3sH
8NjMpJy5vwku6Drl9nW/HFD4mbsl1waL1RuDi8slqvxcX0CGV+0iQNNgCsmiIuZU
G/GfvAKwEGvzgB5HQKj5OtPlu7mEtLvSwG1p4cru1hODeRYvsCp5kO1pBG9kzLoF
G64O+9p9HN9j5wdtIL7xNR/XucJ8gihNNdPwtQYUDn8rCtT+je8snFoKdlf6uwoy
hU0E7WnZh5a6pTNBb8uNanH7gmZx58LBIdBqZHL4cuZTfGoqus6qLm4ggMBRojJl
e6MPqZLojxyjV8KU2pzwn7zbYcD73UBG2D09lo6sd0VYYmwmUDEz4Ovp360U/ylY
k74XEZlIywpwAVae8mYLJ062kV940nEk1ECBNto8ccQsrpTu8rG3zcRURrDcLrdZ
qGrUr0RsaB2szhpBdlJQnXnxDBhiWHC2A4Ekh6AvaLpEBxohQtsBihNHdbctfZwm
b82wVLMTCpRVHE+59aWo/JoSaX7FWFQTMLaGkmVxvlFzMR77VkIBwxGclUklRis5
6arEA3uaL2WRDhFBTLdJFxJyIgUQca8u8fwlpDw/EG859txpNfm2ZlV4TvY45fki
fUnqxcjvqgxW3tbu551YfMUDG8VO1zlgye0IzQIkyEZFiAoFcH6BzuYKoKgrPKx3
y+D7ciNNgwCWfHKQLuibKMLASVF8H9F5VzdKOh53l4VMyYpwxAU9ukboKbiR2Fs3
FHClJQ931geiz4TNEIfS5Q4oVBYKPVAsxqas09bXBf2iGenpBEZzK8JJamM8kAxO
1BQDYaJxLGX7TMFfjKdK/9v312ahGSULTtStF9GNDGRhno+Xn7JLpiBgadjmmunj
i/eN9WxA4SaOWMTwpi2xFleuJ7/0B1LJ0UhJrGbmaZmvV2/3UOH62vbhgNrJNtkX
v1PHl5ZsskGp5S0BYtNava9zxQ2m9SCgB9shJQCfKq5CutTupOVIIEZXFcMGf6BQ
kmA4gHYbDEwcqbMWardt6e4I2y9yAsOfFfM7nQ1Y1tVuuXPQTqBcJI4Fpp87Fxrb
Aql5E7dw8jEPCZt2UPE4hUWoGUJSrHG9PKlOxYkGevQNvXPMpurf0BzcF/2A4XFL
fPBg9rfTComhryncwjbKe8mI26mO6AazQyWDaNIWbBRyfD+0CwsH5msDcEZ7UDOy
o3EM9yRCJqsE0LUBOpB6/lG4QgIEUV2JGyx5+FDvLDLSnc+ZAOeZUxv0wKDC9/jO
53GZJoC7R7iRhOpfTjO7sn47IvyZ260tYOMQHojubD5YSrHCBtjrR/y2LgUuvVw7
wSR3aKVDeAAlVgfmRn2QBRZyIFoPw2InyRTzTLdjUPxN92KxPnQzz4uPeWEWmVUc
I5jGzCFNuiraMbSBaWVxmljWjwoeS9dzLL5JiEL0vClEdPO+NVrwN3raO+OMAgEi
3ckAO2uyVzq/EYdRfAJ6RA3r3XmDI0b+flHwR91IcIUZhblefcIGcze2JXn9zrsP
OIf7Zzs5YUOtZMTwIBIDXADAOeMW4/RsmNgQkpWZt59OirGmoB5y8S9Bbmwlp2or
lVSMF08qqnZ6cbPdsZ+E6ia+I60Ub8J7RmhfUzIL/6+roVvxjpr0HqHNDQzYe5vJ
7BiMJb3Ye/yCTXPtrzkt+IrOTvfueqTIDmhbRaJr/+mzL3PpEMr6lezUnR3sDBke
FjKxv5rsAxa0wIU4sMpQ7m3xEMGdPO6g+rsaMwbBuzDofQVIVUhKdQT6YVwwSeeJ
4XzMBHxzqeVZtMO9cj3H9Jpm3u69/u+DH9p691ITk5ihL3sqZveU2KM/xIMn/DOi
XwLgWW7NRSRwdZpnoHVQu+l/gvVBFByzy2ngAKYBerxjwcJKIcLE1jr6qJk7Smxt
1kQkBTOE34CbG+88tAjH6TFi0r71M64nsRlBjW2NiyD1PuVryRzW06hrni8RbZQB
ZQTCCRG8PPvZ1ZZkr8dxDpiCJziiEAExCE1eZKV0jzhMIWNrG77EjGxXvlQP3ks+
gHFZsMIvTJAoELxHMAd+eTmftXNB9TAOmHrhIMieiYqXpFD0OcTFCt1uicn87O2H
Tks0So3vYVEAwOhBShRA8jIWqJFccP2gLqizZt7jKdu9YnGjKj9rKmiRJplJw7Dr
Q95TubaYVvk+2RVAC/5R6taQxxfCta4E6Ga3TToUu8q1wTN0ewUKEcZZT+9d8cOh
X0H4w9H0geoXQahIs4enUSu2gp/P02D3p9p0QOnphqk4CgPOT/2RIZioHMl5CxJb
O//e8CELU0L+PoAd7XS2yb4ICOT41rV9OATD2DQhPIXIqX3alC5TgaSjAoX63gKi
31RUw8JJ+TFii7kCrYKhnshUIfaN2EmcqGOQSGA7q2j4pwwAZz3JXRWhm0TjVGsD
IgqHbEg+0oQS7BNsdTbD03J38Ec7xuk/RtD4W6xleCs/mp8S0dHVJe3Z8LAMo2qb
hVxjRjHdYYUhEgrOkMyc8imgoj7ZQsfG/QH7Xk2X+TNsokFKfMdkP8kBfR+ygA+B
73BNDNB92Jv8p3Wr8BncGH5q6kG7hjBC+VOslgzgSkJQ1DDhca/IWtbxVHXKib3g
0kGF3pRWosaCECxmkf2C4wXRapf4ez5DJqnaR21UpcPWdQBkgpxwTHTIvjc1QpOl
lcZ29LGJloOhMnk0tjKv4MjkzFzMfVMcNgoH/JtGFnYp3C+Dcjg5qfcPta8RtiWt
fIawSvfEOPu5vumo3gFUbd+ZnwC3GUdVlCCpGU6SLCNLaSNYcoZCMIDQb5v6gWzA
htsSbaFnyYL1k4pidCMw1DvIvk/IsPa0hhUkj4m0XnEs2Odkko9FC4piCwnlQwaz
DyoItNKruUi7MQzGCGbiREC+HMVATqmcUHziHEo/7eXnIKtEbm8+HYxA58Zhbqpp
zgzWbQQ24Mj2I0hVKKyIU5b6brLbuxiauwCWpEb/Cipx/ZdYSuWA21YK7Ag4Vi+W
zsR/+HKWKRDT3htS8ZoaXKhKj9AOkbytjOj3XM83/KhKt6j5aaHMQAJIQRSA8HBg
VOp+1ebsCXxuh6RVQ7eoWyvwF6MdIdcaoC6pFT03NyQZNjwOFAGlerRJ7uT/VDIZ
FkcEOlXGzhZfKBFCwjCyDj9nubtcom4fPYhfMIMygVOhWmsmDJkasn4e2W6TVAkP
V0da1YsuAvji/MxvS2keHQZ6vpHJ1HVjC7UD0dymRDBo1TpwRhEOyQIfUeBv6KCr
D0lxklNkCXzuYsB9w8sFrZLgJ1OnKrIV+PzPoHzZ6Xhyx9duDmMlBXuysTGNwXzR
TXvUdtdBSOJdcYhzKb/E7DUxP+fjvupxzFrfOeQ7ExLsGDiPaQFBy43BnoJlY4f8
+equVe+IKoPu0YmieQj1y2HB9zK3GwGszi+2T8h4o9Vrm7mJbTXa2+7LDVTrZyel
x4GuwC6eTTr9vfjmOQ/zMLwBVgMFmW1iGsFQA5c5NT30FWvdKgB3GcO7o9ZF3MBQ
IaCYEohpjECtvHU68iOYLG+NkrSqgHMJniGkE0huujE1pEbb4Bo6F78ijB7XI3wL
qau8X/iFYmaMgituMbFLUBps1laRZp6usVLuZTrVCWvEFKHNG5/Zl4JIn8xmsxsr
1ZgTi098zLjgVHCZB+rNZmoaQw+q7ugUJPcPxJgpyhxYCvh3E/PvE9kZF1TFdhgL
BNT3kFlyba6axrGbu3l7svQGYCXcheRd4ZGfo+vjOM/9/CgrbOBN3bqUgJMQl7DL
tlMzlPGYetEKW8xDPZQkjhM7HB9noS0kQo5dCRTInxFI9rIAr0/cicUBIgWurJZl
l2ft7qcLfW9rUMfCwwLIq1pAeUGlevk3zqVXnjZlB9g94mX3cyZqvNyWdptX/ZqR
c43IFOPUl81sJ+FYx0xTqJ9+frJGiZODgoX9MlDCSPIaP1bkG/hSD36DL5XXlDFP
UcYVU9U62oT+1SGSBINl9zpQFbS/QBJzK2ALPFbTIE/U3UHTAwRqjbA2xzt9GHl5
WBrqp5ZWb1XXrdbEUtTzKrSDaUZrSmQg2n54mFHYFRcx05Y9yYkITJZtmKMH0Wwu
AggDo+UMru3HydIy5xZEks/exN+gMpADckGpOViCNNHdvMyKqgOUWxwogRaUwvR1
ZJm8JVNl0Ccq9BAfRezEGd9QYdVn7Yx7KZj0vKZ0Ah/1/LTw8LvwHMwPYo3WOTdU
KS1Q0dC8OTQoEgwKlVI+K+uV3KO1ngjf3gUvhRP93V3ggk5RUQ+4jJwecqQDPmlx
oqlZzZIbJuX8vDHOwZ04ParBiV06g8rSHrHHKSjYoH0jNw+qwSTzqSraprSgb19d
lrjiOKkyLZcwK76luSDotgv6+V9nzMUat5bru6um/DqzDr1x1TPmIR4ZVlRZKzv9
CYld76R2mO954gLLgtjUA1CT0ab7XxhmHqtqYAder/FSJWvwWRiyjOSyykEj2O/Y
pugCshc8UlwM0kg7kaHb9bGArxJN4DYorUhW5WsqdnDvAPh5gAIqOcN7g4bIAjY3
1p6nKJK+8+qLL9Viw/GrZQ1ij1bjBbGHn5pOx2kp0xON8exdqfkrUWKniniUG5bB
6PQvcbk+IbOMxUbpcIsPxyFWSN8SrDJLwaE7y0BRStTMYlS3HM/4PAu59eaHRQp5
lHE1wX5hpCbE3rmxkOuhPgjCb1wzKI0X7GR0MWf62RzcHg/IKS3LP5JIj+2IoCnL
8V6c8J6h1WIlNQ1QzYgF/xDlIAVTF2oUnFj32MZXitVpsriqR2u2S+mo6Uj9Yux1
MJhOn5UjLQ/dCQRq2VbGOmRyOGJrXQL4mEWT9vyG+T4QskLvOxg+QTcmQI9ISBhe
Xl6SkctF2Dm3GjyyyVy3XB6iyAbka0WScXgnH//Hp2HQoELKqOqvYAlF+7AR8PEx
6ik5xCZ8silnmv+Lck2z3HTNOPNTRrhbv3ISwHsTaUwuyp6tTDrp/0dfbV4hUPkL
n/h4gkmRkK10++J6l4N3Vt54ouk0IBRbCp2I7oNaaPZthzUDQqo3r3436tJXXJCj
tds/1ksw52MTTcSY/NewbTO1J2w3Bb+85yoVkV2SQYQ+unsQ4mTySYgEOFCrwxSC
uuectoo8SBrpmItspVcmAUPGsfGFQM7tf0IM7Zq0uPRdKo5oX+OppO8IcnNzNtkh
VK+jwqLm9VrpQuUNPigJz8R97U64M9Rk0UN7fqYBaDdQsthRhyx19gN6qlMofmrR
53touyDs4IKqKC48R5hzpD3Pumk1YMPgMiCe0ppPh45DfIOyophMgCfbngHWfa6L
6lAmIRN4dtCD/XVhCm3AVulKug+NFs4Z8yAR8KdfW3ERf53jtNAsO4tJUpaX/emW
yLYFawiBIrk3RGqogIE+82WEwcBsQDGfEKhKoXTRAlS4UpD0mO3lGcKnIEHTYnpp
k6PjTTE103VfO7CK8bK47dmOrDhJmB7CxJIkjYLKRSqOA2oBgV+DVE9OD6aN3QpO
gGj14qqBZNp4mllFyFsGKOqOm9dUkPs1Ejp94+sSjuyaTRK1U5KHp2FGUIZKpuTx
euHzx343pc/PeM26WX3S8z5aAxAuUnxFJ5NPZZ2gbw03vJ12/XbaS1WEHwEIavb8
MFTi8YyhGYBk+TSNg3LhFGLgdlFWqQvOKFQE2+2xGrEwOIOc+QUxvNqlVEfl5WkJ
V0p18goelTWwLPC5CsCu+w7Yl0GpAU6mv/UveVSx9zA7sBEIoQXkp0VzOPm1sAzi
dmGyRwBZmAd5it3ouwFg1fnMbmGnHFBU4KUSK6a9B8F6T3fS8s6H9K+pt66EDk3J
VvMsiVdcM1tbv0W/EjtIqzMy4i2CRBPNTJ4g6Lody+uzHDGxj2fJ/SIRdWGVTd90
dL11v+TXC8eg7h90bwWbXIFvcVBcGFb8aGFNFk0gwc14fvbq0/KXwXa8xoMGSICe
fZeLPf8/bxq/rWMn1EBgqEZSdVMDO3imAVpi59FopEDmEhT2t2eHBX0+0XGu1zQL
udBGiT01RzGPMsq6i8o9wsRj6maAgAv/BvmUQOZBWcJdGlaE8VlFaUD1mT5KSde8
f7p15jt117JKQt6jHFOs3vin0wTCnnnmvn7sibkKP8DaJodjiQnKt+8i/Amj/KZj
ngvmY1lbzWnB+Hd6pi5z/zTLPYLBO/kkZQyXzccEB58dQGHxjqKOhR1XcBFhEEOD
SaUP8KcuqxAaZIaDo2mfAgRFb0l89uXdcw96ZwmqTzL7TOW2LmBMpv3ed0vPNB9P
aPyWXTrCBQiUdSnTJ4Jb6V8EEBN6d4ZXT4RxViRGx3h9goVeoHhmsanA+CbpFKIJ
emcrqYYkuSw1llD+oqdrxf6udRJK4zxha+4ae9DopQHqxDKWPBZo+EWGassoGJ8F
6jcL1aFKQ/xyE7NZ7XT7gWFcTQAxSGSIIH4c7rjG7cAXGs3dBKTtPf9sRKnNky/X
N5OGoivdlcERbvmoXl8ckpDR03kqvHzqTzTJwPPzlzl14XHe7MOkljb1+sXX918n
d8UwYg3N0H8SgXquWR+ldegyJpkaiVITzGkNlzETkkxdckQeFb7O+eVSsQ32YQpE
EoLRz1SeQWJMfH1Yzpkdd40V0jGzglmxNR/LNbfyyYukCL3fndaJkGM/q1u45e74
8q2P8f06a5XjEWFvbe97/lob0K5lUpsT6gqkAiIm89a5yrdN5WEYz9v9636szCvR
kRZYNzq6n2vsSciGm47ganmQYBzToLny/5HyrcbhzXJCFk0gpWn151RSlN0a8RPf
gAf/OhDCYgztXUyjrvVwVtfGrX9e7WQDHxBmVW6JLS09t00aXE5J6nQnMQqN1dX5
qYiKcXq4c94y2eBz/Zj+1ELJCGGD+vvaNJNRyvZfafEbAvihcBP3WAKuae32ARD5
k90LgbYM3ZPFUbQD5kThTS8qPwZ/DJvcAWWFOUFex40xwQnpqrDEmgx2+JiHhQf4
nLmnWmI7GZ5ZwitC6zgIxcxJ2NtKOzfaWDfkxm48+BtuO1VUHFsOTz5LsDYEj3Ht
JkOpS3mxzgRmPe4UzB7I3ZWXOnN2JbGG+PjxuDSu2iLoABIZjgsMFTkMDT+khiwh
TGlWhL/FkPVkUR4A9VZcBQqo73MSrBJ8dEA7QbO8pHvEn/U8jTK9pPGhFBWuJrDT
tBK4Yi7kHTO1AxK1kZO1HAo5nAO0QOGijbOWF7Shlh2VwZJ6rXuLtsJQcibfULND
Ixp2yVm6mieA0eqtZYF4we3wKnAdFy2sLcDEnvQr4dDvqZFDl725D4Je1L9vO0Xr
GZRaGwF4RkpNn6hGCjszN1dYlHXZITD1m8ox451KOH+ZuZKVS8ovxDdqGGdh/230
aOt8/SBg+i5GW9E4HXsKeDGG4ofOC2+3UNPKxLKnKAl2zNIauL6k+BzyQNfW6za4
kgXJjeFHNrDoMTk16pcUnmNxk1JRruvWQLWH3yiQ2uuJQaASm4+SF9BQokCPx4yl
VIfOFkFekAgcPGhIW00gLM4LovWwnEMOCNTc4YNv9lA+wM6x7pIdbQbHQJSl8u2N
EwA+hTu4jwhDOLayrKbXBPwfePsKh1OuZnk9MUd8KKiWeRCbTxLITqMVHCQ8o0f+
kQEQQj/J9Lz7xVPM+S4OpBnlNxfK1thbDBNUFs/ARX7aPxTS6CgpzaDRSDwKncnj
rGKDoa3Rij1MEiUPoV9FMHTxQwkvjYK4Hay3IRZKrDo0h0Fh/1qEvSViytXnocA6
xxyb709cAdPc4swlT9gAQUxY1BmP/5lm1n9h9YWBao36mD0al/GHbobi3mEa/goO
UpO/Rr+Cnm+Z3ZbhctGX9yaim0/yJj+T5hhXgCrLbbRhZ2zzISk4JlhPTspYeUeX
uUiGss8pjQ+DSzn0/wxPKO98faHNPvHBV8fgI1AucBau951nbgMIZ+ab5zbDP6fM
cqyTPWlxLIrg0uWMr+JkoJXn0p0LgRjNmPPoc5P1/uSEuBbXym2CIxeQGq/ARKm/
MM02j9pw46ywyROinj1f4hDEzfrmhPEKjULCZkfiQZb71xuSPP3UrtGTIKIx5m3n
CTdxocW3YO1o5Bhqc7dnXjUh4YW52CzOIDgMrHnxukIn53FrwSIPgTUbJKPErYLT
mBYDzpjr789a+JcfZDoqKcFaHBrkYcxQoNoZTTr/M8mt6+xjCksKUkpDZD/lp4Av
kXt9bFREkWc9xHmucRRoMnaDGvT73xn2PMKia4vwI/DZnzhBnfCBkt29U8cRb9bK
ixkt7LLMohgo5Szp+mLCKZunE8LHvOx0783vjKEAfXIVbFUHzoaznD0exGpTeh04
rjh8pkfYAFt666lFwIWBs6VEB1Y0VBYD1EL+rS8tuu7l1z9Tuuv0xkIICBAMefS4
381r7Yj8nYWCKp8wZHPp1KRT3bPXQutfOKaHA+wZVJjZT9oi+5ZAygIUTJENuyYB
lr04G47bfv3j7SwvyXNZMYnrVxOZS0LnH0F9itQtLT7exCoEud/tSN0DwNj8wjnP
YlxFCy+liS7KiTM690F5JLhIJytnFcS8nPOPyG7FtzxBljl5owZkNMa1plYfX3HB
RMcj+agS7RD4DjBx4Lp0H3hUVTRJdB1C1jQMMfp3jxkIP2ah/yV4ng4NuW7I1ILN
0VW4baiimoI+aV0YndVagRLC/8rHOZY8i83SXiRIQBVxi7l0GDJ3kOMsyTCYTmCe
plc99nZcTrUb4bxwPH2bQIc3+GAddxpExkGfPGslFndZH0fgFXwE+CSrQw+6+ygA
Jo8wK9Bec5Tm5gjpSXSNVdA92wcwepwKrZ1RzfYTT3qsIpNAiHZyTyNXos3LLUg0
iCd/zjHgtkm1+CLo6Mg3wMaZCMAqTH/UFMEe2j03WPXw51dsgtLO4UaU3A8PvUR0
1Du/y35GkNBXmwARXIK+kz/ABpRuGO74nR6zINH8otvm2J5LvnoyfNDmtdye/WBN
0MMP1qb1tC/qZdX6nVW0mcTd7jhx6cHGhZxOEeXAK9O5Ks0LQLPKHvxbjzm9KeRF
6Bsh75/ggpaBAHCbRJd1363y/aMAG6jeMgRcOod3SKHoLuiNBbdKye9yAnjYalyy
/mHFKsdV5JMZCbtEBCQgMqHSxJalwp3KIMIdS1mCthX2VtsEIxVOz0ZoXTcGh5OM
rOtvcb45aLwVaiGv1sHqEMLqr3DU9VSir0FNwUqioGmEbL6B/FfoFKb8iEokYL+3
3WjFiNWvAE/GykjhlswA2WhZ21dOnxYiTVdcjXsnof6PV04tgUmpNGay9pZxWLqN
a7YI61UEwpnblU5txMjFQPnVcKHQryhV27Fena9+gmYCqUXmbnqEtja60qmFFSsr
p/m4EfslI1z4MbGGVi0WXmQv9HbUSOjiFT3KWAUj/mNTpuUw+I7BrIAt4CIlDeTE
jJGEWJcKQ94+mp+sidlNn1p+DoTEM3V2w1quOQ/BSX+2tia+9mpHgEHGwKS84sx0
LWC3NfvBBQfiYNoIHt6uyqMjTQfym4HYLpUmwbhncDh76wOIKzLOmLRGlZ5iFJ90
kky7zuQwHROPKrg2hUAGbqhAtU7ylucMSfsxCAx0lb4kFGKcr0ZjUoq7HWaqit+B
lEA3mrnJB4gbXvMEyzha0EgUgVYTNo7HzeKOjcClNXY1GCQqpnfa9GY/Xnx/raad
F5dy1zMBeo0oOTAsLe6sL5Rfbbb0IoizCh9zDKh76e6bENAlKE8D111zl/PANyG1
Ygzn2RkVlQil5zMCSXSl1sQwnpRmUooqfYySUUpfha/quQhYoHkobDI6NOCOY+0u
Q520Jn3RFRgsSdkTAP9D+PdAWKC3uNssPJJXyZNJucyjFpWLk88SYeWCwUtEZhek
m6YuGfNeaaw655gvUNL5J4zj+TMx6ATF7Kt4yE9NCPxSvENonyY3/6JaOjX4VhQr
DULjFs6dF14qAeZfCNlGiu4V5l+hgWc94JSghuFFbF00cN1Zr/wckA8gh8ZQhj/a
gRuN8PicPZgRmEcC67JIZTK3IMqxXAHQkPRhOP4Dja5S+5XdayrEWLQIc6Cgm0c6
bvREb1mC8aVvdlqTE+HDleeYWjH8D/o3gJed0+HCc5kLUOyQYDwswsQArzSffFl8
npqjt04OMcJQr+oHajEsbbHAhlBlqLnNMd3ziu+nW0q44NDNEowqgHJwvMdevQmr
SSDOCwDNOY54Hf+SQS0pPVdkfSfLNT3xV/2EBaz7tgcD2Yph2BBPGSpNU33LIJoC
a7+0oHVk/YTytq9lewStMwc1dgQtNPaXE5l2h4W6CXRuPbRjyO4+6btQQB/GUxvS
4+MAvAAPfavImPA8CAj0kEHiur92fSgilEQswKzj94FROSMC/WnLeI8N0E+w6O9e
A0JQVbQPh4ZF38fUy6IAGF+ploBjcLMkw61BGV0JyEBPNxvuili6+2zGgQJC3Gkb
YjQ0X8yHUjDETxC7Vrw8a8r0fRtrj5XXCnmYAt5lTlj4mHG0Uc+gPR2JaxUGP4vg
g8NcBgZEscsDnwpOpAAmF3bAZhKbeXYNWTSizwpsfki7YCDMmDTV5npchQX9FWGn
03G/1DzJyeSMjwz7j0k4D00VxD0iGUIc1yQiST8J2RpKUthzus39ZUAaLkK/X2Wu
LhE47BKCY3HlMxeDCmyAg/utL7uMIw6wlvH/4t9vpvVe+phaSovBzB4QUsoYz2l6
Kx2+iweVbWGCIW8+8IshB0QUuO6Gfc22rmW1ZYf4dWc+QAdOq2Qxn195X8God2Eh
Fg8RkygaK3kz4XIeyPEzu3XaL8ky6reelEqipPl5n/X356HdCBBPPRSR6PcOgZLK
fej4VsvZfiy2CnyLxe6aBQ+TAYqNwtdZS8blHbtt33AlwJ48+ysuBXXRKhiacWjQ
Mt6ZVq91KrhFPescQ6wPKiwf66sn78tFkovTFddCA/oTcnk67RiVQj2w9gWhxAss
Ro8MSSgjp5ZelLsR3nUtNQSBP0IEtkqV1fWYV8cG6VOjOQkONvYLBCtAvPPJJ+Ov
0Fr8m7eKzxsrR6ILA+SuKeeBE1wWsaijvXvED5KnPN4Yb3Lvkr9x6sEDEO+hUIqN
KX+MqWI/Fd0t5dsYbe/Rz+bx7V0UI7AQLz99t3nyamSOFv4Tci6YpLdxEcyWeQZ2
zim8/9nr+qMiW8cd+T7i5UAe6yGUnCQvUuw5t0jzzJXjfOdXJ4ZL7/RelDC7bQy6
dd1DPabGHv4CCSQ7bSzjRySsGwxxQd/54bP48OlbP4/slIbJAq/efDInZL8MyY5P
Uyo8dFQYLxMRuwgtf6XPD68vkPFS1oR5ufT3ILLWMkpT4Fc1DZwxlGWBgKPpNj3B
5q3fyvYdlZbB6hbwYZYUFpXh5m83eOFibu54fCHB9qcWXbM35UEtcYYjpqOgNXrU
WMbRiSDQ4SIl03VuluQ9Ndzj+RSH+zez9sO8IFugwOULNqoJh3e+1Hnw0hjyPhOT
c000Dwolmmvk8DqHy3jOFXZMW/QAeng3GvI/oZCG2r757L6J2eVMSpqzOLIKoPt9
Q30OphYjd7VA1X3OyFcBF8IdK5JbCQKU1pbY1tRoJtXltnVT2XJwraVOgMkfvQCV
Ul/BkMJPdo3quMPE+zWXE3Wl+mkoBC6FjLq9SQ5kV+QGttSLV35VZGP/fxmJlGkX
amFL29yMVZsAzNMA9+kf2u2ognMMpO/bbC4uSwtdZ3ibkRGQ8RIVmKrqc1hfp2+L
ITDRORebDSKQElU43cPvtduJyUw8SBxw628X34/QD788xSQjYamjYVjP/f0dTu5a
KEOUwhfgK/ULr5PFv3bV8u7n28P9rZj3/x47ZiRMZdoYUeanON3z/7KRqr6PRguj
bAsqsPYmp3+2TkC/7BjWkKwf65FtYFf8BLJC/A9Oh+Ma/6XGDwCSGlyy+YeZZxFv
0HX4c3ihqCLm9agp+EGS2Sw5A3Jengd8HILf+7Bd5/g8lVbqxnswMW+7nCPJpUYn
ybs2CSb1iqQhZ2iW9e3H0fiwgdyunTGFUepfMQOBbujqlZLC0yhNIEXWo0qaSR6b
Dq63wEsv073Tyg2vtROkOkQ9VXHxxBpB7eAqg/hY/BpWupFL7TLy4+zhtskrjKEd
tHyeeBFZjQQmx4xmTP1aNZl5A170iDyV6LgQ10UNufu9s4XhEWp0NkS2F36jmVAi
5s1dQ8sjgZXm2aoAz1tFkjqSpKMImrIIO/4zFyVN10Uw0KJyJIIKI2a/2PROwUWC
2pvlgY+AKJkfx8F50rJmM0LVglJCXdrqO15eMBBp9Hm0WI4B7bzPk07YOueVzagf
vaVYNqfVFZG6uLY6QqHEGk3UFAlb+Z1YuICIK71QFq/WjMHZi9ZWd9ARiUpR26sL
NkalDKnNR094WZsVf1fCTP5kAs45bM2ng36dGNhGFHMYusHGefTuA/Wvr+MkiWbr
tNzziqoq2U//ayoAE9kTANEdGdYCbJ9krDxTWbdbemigq1h1sftTXzsbb8JtMHZw
c3PpQWArnH0xncKuyxGORVtRnuB+tFF7YXu8b7gJtXSYzNImBYr6pD9kQmbVz809
G/59n24wYhiEC/4I0ZEz/RP9g2KcgiIHSFKmOrDLU5l2rlsD92iW7yws9fV0LBsO
vPxMG3D+qVBMUJC/eYfxMWOw6yma5EPlulA/bTfupoxPpAn8xJrJ6hdZxbcERTQo
9Gy2nfz+MwoqnbWiHwmscp6jkUXEcTmWzlEgaozBKqPG1AbCxYSqccLuXBZMREND
NuxixScODPySq6PTZMQ0266qxCJb+NZVYUbbc9/erUt8K4RNQqyJPDOjBWr8ybKE
/dziRo6b4HYNXQ/3SIIenoM/41DHfP79YNsL//KNW9qJwjMGMX2CRJgvdXYM93Dx
9HWWljR4BooUZBGotRnOeBSwwiIFXilW+oM1Ct3i3J1Emq10d783My2CaajlSKbc
s6mNSTlK4VgNCQDhty7flOwIDb5xq6H/6B5Ri/5jmc/m7C5e/sQ8Tz/IhX1FYLTW
QEnKTKX6nhmP69UqI/unZU3/0QX25uNEaICYcoWweZkpzXonsZKchZ6F2d+0h6aS
tMxwlwKPceSs5UuIrQpsowygAkZn0YJ/mVsQM1O9YtkUPjecmU/ee9Ptatrq+JDe
h9JrhLLkBncyDql90uYCK7H1ohW/9tn49JHR02MbsxGVAf3q7WvYRmrk3dsHSDrs
KXPizjsKwv9jlyM1UDF90zofzT3Bgtr0P4AkLH9NxZxJkUTcrAPF+ZUc7kd56r1Y
2+OrSvaKx/8NDWpv3zVaogcf8D6owtbgEA0nnF2ViSKaLR3OtF9hX2r3j7UnlVEn
SBo7qwx0bMRORVCXZ7ZeYujkQZHgBcqe6tw5scJExMT+jwbtKLSfjfc/Lyl85dzK
nD1cSFbQRbgGv3XFtp8/08+N5le34b3SfW0wOQMztlcj1nULbXN1OEha1n+OkKY8
IyRFDR9D/RzNgiiK6DpBJID422BAlUYV4j4UlU5mLiyl/edahABDzlEhfu+k4Sdq
HcXQcxkx9pk5WhNTN1b38VOiBOYe22dHdkZy5yUujGnvWaEs5bQh/z45mlqJH5Ed
HMWns0mV2YmomeJcN8NTuOo94gWvPzCT9ZQ+aGw7E53PziK03QrvTFEhGj7B/2Cj
4LvflB9oAj7E1c0xFL3jxCkN0iLrvaYDFoOHgqWQhNacz0Uk7XbGoC/cyg7XNBOr
oNT4l103QCHwWFZw7bwtpFIs8ao/La9vdK6qz+7MqmGI4J8yO96zHm0ALd5ZSNQn
snwRBh6X8EinC4Dip/DtCaobASj1SIo43JhrNR6lqo0AlRS8A/3u8AisI4l93FeU
vZga0OwOfuWhufvyjESho92RF2Le89/5IsZ30yqZLQKjtWscLOy7yEuHWxUD8qCZ
0J2qgYYwUkgZ7UV7qRjQ+F84paRUPeQT+2ZYOieNXa13VsmzR87ywlBb67iLm4aR
g0PaGg4IgpYhw73dL/dFlrT6oxMhyILF3C8TiL8kGy0V1+DVCRYXz4fVckRx6p/q
Vl5BWM8e19x4aRZnvpwtCzSzsBuIPZZA0uNv729wnBv7XvIS9bOxCQIvU8iw342+
c9cri9FnNBq+qfzHIIRW51YMbM7AF8aTtMUyf9D77Zn23Yas8EUUkitSM+uozxpp
+GphlcE2sok+uBHlZEpvVFHq7jdQA2YeMMpm1t0CoWZx2EVTixZL0R0e/n/Q8/7w
IlT14/WhvUCWkOWHApl/u/IVK9uUeBoI7FPWKjhdbcwdPuRLdDznI0kxrCf8JygU
XyO2MUzBfJHYlImxBJo059xhHzXub9P6BTcCeGeV2EMMjuPg0B659PQX9MKsJj7R
L0rRD4jUCI4kI3t/x6VOFhEIvDgWDPCrEAfWIXX4FglQnhIQcfQYuz06oGhOxPiX
WZPbe82yovaRDeMPhDTf38zWIv1ve8esNkv380Y4Y8gxDY9+7HrNJg3o77hj/a9N
XWYTQbj8YGpzNiCIJIvNuBuwB1Peqk/LuLzqY9SVZaPckUQJrwe5Ph33wiqvtB2U
Swio5aSBsfcqnjI9PqvmHrJIkF0EkaU9Jjz6wXzkjEDPqGMQnqJujpqqxsOORPQY
2KVMQujvPFOvk+6P5DWajyPWgCDweJ1fsPOQpgDKB+XLspav3hHbVd+8w9kywB6F
QLOrqUaJMJX+vh2/wo1JsDxiZkrFgNpu+BXzqskCWXhR67wlTjcwz8YTEZ/sHlDm
L31N9tYwkSbArrO/gvNMukBb0YCRjcH06MI4MsAjTqh4xJxQlKwuY/X3bbcLgftt
1wGYxJgdPyw+15ypb9FVS3E+vhYQ4OPk0diZlNBXhXuHPKK7CBofCFONmxwcy/Z5
Ck3Oz5q7fo13dfneyWLg95PPrTYnqXwIfT35Ll19MkDs7tzxxEhB6OIZmRP9BsQg
iwr5+lw8twsWhtfz8Q4y5WcdofgWc8MmM8In5yvjBvy5XJCHr6deJDqUeT0+rxhj
ghSOWTdkGjaWqjYCKfI3jYiKZxsYagPuJZBc43mV0UJm6aHpqpfrnDSa8wP3uozi
wmnT/QhPeDALEI10bLQhZ36TG1aAziOUNEb4trNF6yb7pFoPE4WnEl+pwS8GpL+v
eCVJUc/J7T2V2MkqGazGRBknh0Nmyl3lP6E/l1v6VgA1xEDhH90dpTleTF0TTsau
uRhPXs/gHwVKBOKCHddAN+ZRp4r8zJk6LpvMiklvtr72k/lzv3YZSHbAQF4yXn18
pRmT6lHVaWTEFI5uAo02n9geviCB1IM3CcrNtCR6HkEtT8E89Z6e2ZdYu6aqjbDE
2IdQxRPONUB6tpTNGgHn3/2sfv75AE1NUK5473A4TYLwZNu4uG0cAgtNtK0VOiaH
EEiyXYr/JQb2Wp3gLBNwZFJwg07silYVfluzpHpNLSvdn7BF7rHAjUDxxpkdNXgI
+MGRqsX8+Ide8MGq6iGu4K83uNcYCmdaQ1Yde31Zz8kFPzKtLMDHILgiAMYAV/8f
CDAZrvN4rPZ06qXO4vAsTI0j/tpST0w3KmXm2m2dPUjU0dvaJyWCzye72XNXEUr9
SJ3L7+3sfytNKw6Lml4TX1Ds24BFDI4wvojiryxW54DcAoGtnVDn467Oh6K4eWgs
1Qfyow3UqI9a6iIHmqjk7mmkEJoMKlTY7pjULhac8ayBa2CsKaYh+QcO/gYEwfCw
SwSERvvx6W9GrnSzfWHsw9gsmSKtauSCmcHYY0+0sZeu8qnZBUrnlEkNorFAfYXJ
wEr6n4myn5XsvEkogMqzk8u7PX8GSa+DaLQmgZK/PYJYdqAU+vw/x3//NWCBytnt
x0uFil4ZJ3vWAjlfLrU30dzBvSdEfZZEP2IP1yojrvx9JkvuLzO6yYZud1f+bTi2
OdAUtqAb/PchOmuRfMLVgeHXiAcHf6quMmZATcvM10pqmf6KOoGdD3/1140WcZMI
2U8qfeNcBo92stKXNHd3kCzsT8HpgIVIqhZhHBxK7QMNRwXo3iVaKtrvGO1PqEw1
UQVzICWEIrCFwk1zgIFZiTvxvqKA3g/P8GlcoO6ScAHYVWOcCrZqRKqJILx4/S1m
pULC4mdtc8Mf4HrbvYDXhwYFg0lNTFIM6pIz2uLXoT25apoWANQT5oxO5yt1lWJg
KD/shVL3mMD2VMV71ziIbaRzFpeiSoWO2+vHHGuQo/MVf8yqy3uRpADcJ0fwiobk
PjOm91MKI5jivFEXmJsgbR1NYlSNWkd4HKHO0MsHo/xf6gv4EezFx4LQrkNT6/Rj
8A6EboY3AcxX18tMYeKFTZnFx5pCEnZPKrz4coviv+g61Bj9OrON+aolol1iBWhR
bP/XTW6Kv7LcVwnaMjDUC/uBCJilaoCAkkIYgdhDPDBetjELborAr0HL/gc0h+Mp
jaIKmM1wczd08yHmxmmJ3/cpUwrqnn6sEhpA9OT9zxbz/JOfhKQkf9D/W8NOD5wQ
nzOXBnlsINR1vriJDjRriQQaHbYMKOSoUY635opZM5UrHonD0+2t+gf/uxuebyOl
JC/phr/nanyxnN6hNMiL76hPwarRnGHwHngzIbDcyEfjnYzjjnXCeTnBs9JpiT3m
asH8Txj+osP5RvJFmm5XG7/vXBMTNU+94nC/arCHQCZQLQSO/nnlN5D8AHJsMlqg
kyKJccSMqmul8RKT0C1nR06GEBPHFnN728twv8qNPW8MP8bEGC1O5DQbk7eqxR+8
cOAeKD4KSy1m0dy83uHBVvvwZKjyEGSDN5iOMXAvXdsFCbwGOG8dDbyPfVJZYol/
7z+b7YC8XDV+rTR7P+nlz+5SlBkY5rCyeiDFltparkFqdwdl3TBxAKhyCPGyyxdp
Xr9vVqk6FcsPg9WWFMnrDKRrhXqr2W1qFGIQIB/C5BWCZFe7XpoIY2PjWIyzaR6E
e93aR0R06DCRQGs1e8/VJvf63uHy+ZI7HmGgJ4Y4JSIOf+FYvEL1kxe3dVzW001I
BNJelqpubnQJengCfwa4UAiFl5IA4X266yomC+V+9Aca+JOdTYgRLHSGQekcvlCn
gJm1ODPGlu8n1B0UA1Y9bgRbX/j+bJRIM7u2oW0wEYt/I66ZNH5X4ALxs/Heqksc
ojivYgStGs0tIAzD7KUElgK3Oy9O/3pDYZqvJvcX6gCzBDIqahFNwoFpYYcByfnh
F8S5xPZ4eIE8ljyYN7adu9S8Y5+4DLqBwoYN4F2ZYh8p0LyVHVMBhPz8JS9OvD6p
5QJct+v5qWosBaNxHhQVUZzOepwkNo1PTHuMoB4MgIhXpPQjQDLRIRcriZ6hXhCR
VX8CO+6cu9VS4hdqliyyfEuE7vsKWSJ7RD7KJLQvC3wO7Y/QK4VDg4lOxHhhH5oW
J/meWabqfDAJ00f6VAJ/CTZB24SmmUsYRd5ERQ6Cbej+Xomxy34NYp0PSDTSTEbt
wrGpM5Sch4gyJ7ipQ5EW8/+4RfZ6jPwL3mEdv59SeL/2uRdVdw9+FwpFTf7v64U5
NYSyGthXQJX8pY+f/a5BpJE7BZLdAZgzJSzYFG2L59GMa2rqRRezMWJ6lOkVbJVT
AIj/mbGy72qre/6HOMASGai8HlOlkhYsnONEha6lT1RygRq+kDrcUeEt/KbZF8Vw
lKer4w2v/ho9VGGotMnvPlTrYJ5ubdyspNBZgRgxNjczBi4Tn8eZvb3GXimMorgY
Ho9sTDQb1NalisAYTv4vBebQaKSql19eBPgaV5KA1dsxrljQHYh2qdr1JNkLojFo
yThv4ZNwQZsthPgz86GDW89wJCTXQL5ts+fPeUNBSCtMIyABaLrQX11tcyK0eWtd
rWgFrzib7lm4cUixlvou8lTxyKbxdkqBht/xxTspNUNP8HEyobm59rRM8rrlION3
fpG+Uq4mD8woSwyCQmh1vKmkBkVO6Kt2zu9T/ML1hxuVUB1ASoUv6YOYuYUFmDTP
KL2XKhUydX2rzEfxI8la5FtOejP9v3D6gU/d6pLrE3HnaKl6de7zdt8JTZquv8Kl
HkC0JPQb6B0cmVvhIAnuayKPVvrPKNdx6gxYlvQh5hmNFjcJ/ne9Z10pct45QzIb
ayyUSe2ojBHKTHGohx/RlbzmB5u7cSY1GJtKv3a4YHMykPWFIDs+QpBOETKr6BYe
4KR5Zf0PTxgpci+KShorr6B6L5HsGP3QQbz5Vi7cQ1ZY57ukMc+lSubNnCth662o
9IKyLezxSXj0NCOKKwkC/fuBhpRmUyCS5xPx2lOqD0Y9aGmHlctj/+kZBhyupE1K
El1OGj/5/QKvvDFTYnq4j6htxkm1p12giRsqWYyxGkZbAFV+VKXwiliHSSWa4mfJ
9AqbPBZ+7JQc3cBuzBn57w8rpDW5UxGYYIIFm2nb/TKHAjvzZxV2WkT51lJTu5Nv
CAT2fT4edWDPZgcPqF16nOutkpB2p2LPmESwMQlRzkijpXo1yxcQfZg/RsaTWvHs
Gg/od3ctV81Iu8eFrYBEefFwcxI4URMKUHUF/QCGX2VdcCa1+uu+WRhtYkEV1dHU
M0QQzZK+gs96rTHzS++dHkxjTz7ahol1mZgj9OSggIx+kk0C6AhkN9Ws9txSfyl3
keHa1ukwky2xkJXwJQai1tN5j34q/uNJiC5B6P7knk+Vx3tTlPktlyqdEL6VMbJs
LXp5igGf8YlXqGbLPwowlyNf/dNvItVzQG6KRvjzCRzPpQk/SwuyU7exDKLC155E
80jWMttUJy4PKnCnhIVVHmVl5vsgdm7yyJgNs1nJXKIov3MQOWQr6kJfg9AUdGH6
BeB9DJxcAldP/86BycQZW4VQGPI0/3Hc7oax9etpmi7mAcEN8eibWEJnteujLU6C
/0KwW4+4f7z3YB9IbcQxwQifMSuvA3dbsXrKzBtsX2jzQIMH0wYfRY8GyqySBuCg
UpIPEAKWO+X30O2mbYdxHrIPeW8G2Af3dO3TGXMh1lo=
`pragma protect end_protected
