// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
d4vbuif+cJWin9eE7CHUwH0Q0rLYOod9qaztUOuMFW+GiOH1ty5SyQ22zxFk4qolxbuVm/V5opG2
Hao7ymnZOF4I/Wa78B5gFQEdVNjGmT2xyI7EW1txzGUf2EjEhQVgbqA7S11oC8bryAw2yCiw56WI
em/kKgnOyov1us4YcAxjAPvnSj5HJw7Q6XAZfuixWS0RNhYvZc9BnFlkrTfBP7vKpAbkTUTajkbQ
2DaC+hhSyCxDapjGqmCUbbrDjwcqNkAkYYUlkW1j1ICJoaH85JpZJbEAoTuFOTUMBAdYjbCEkuAk
mg0sW838o4R9MSmQVunjynSw9UDPHICNF8I3Xw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
bzO7okJPWDTIUoJ1ZkU37Db+db8P+LvEBiNy2AmRkaCZVV6uJ8BZXYrwGt5k3XLfSuRDpK+Nyr6+
jFce2QOgFdmA5c0z3TGg3bB3YLOlhwkoO/uNdsXitKxN0QxuoNQwwv94qYfDkYLvPZJm92B9HOmx
JCgojvkBPPHQOIxnDs/BoNW2lYE3dhUz9sQgP6LLmKhWFDaDbasox/w1myAjbjmEf2o/wwgIEaTi
JrWI/E0FJCVjH70Z2vXlNgvs0DGA7O0LEqJJk24DCLeys4DKIu0/tNSMm/3UNhBxhsJikf9Zs5HM
alCyEjWSUlAvEvHSA1RQeagXTZBGCePWrT/9+rTrMNqznmI8RpEEiQdfIgAFF2rk/qW/NoZIOL/3
otJsZoPGTayb4IpJTst3ZXfJ9ivaFA9C4KX6v6w04tm2NvPcm7pfFuf/KGqu9VyDUinKy9eFpNVN
VooQ9YbP/bR70xfVJsq2V6E7Z4pxOFBe5emErUU3uHRYWflAYc6xN+6XGRNPMaEi/LT8H3+0HLgz
eVowbP6yOBhWDJ3Rp0kLr9bVoB1BEOme1FK+c5Ffa/bu5SodDmbG9YA7UgwFJtkm5KpPawVTGiZ2
K+qmQ0HRbjRVXtxUy65wFi4ES7T07xp0cMgcN9rXUCC+2L+QgITbvfqq0H709ldwApihan9/BWPs
mIGLcQN5M/9T4l/DgcmDy4iKc+u2ZdFpL513dcrbarzdW5HHrgt4FniOrGqg5eUWo1j3d3Tupba6
uwiqUx+/28N8leTUSOVwfTHzMv6WT+F3/1euegBXenejcQeZiraO4EACPsdjcZjC0wiX+2PuYBKN
HTrU3MokrZG+fIlFfBQuR0GktkU6W5OA6Xx5wQbyrUksNlSgo9gBhSTJI4WQNxgRBjgrAd4rJIlU
YYU68B4nGsx2eA2hwQxwQoOHZb7jbqhRJn+UAqKA6W0SWN/DW2yG5cndyplhy1B6A+mSZicqy/D8
wmxLAdaTpEfHDd5Y4lgrGVubMeg+kiYfiw171xayFJ/bLEX9mYaHxgvj6EBpenl8ym+2TjvPIWsS
i9xQKV6VJcRhUQeV9LCNbWJbXYVSsKluWmS/wRiBziEwP7OjJC/INiKjprHcFJ1VE5lO/5XSen7Y
9YZWTe56CPogls1aInWF8uRLzZi43LBfdPXR6EeGxjZyJ5o4ZLs/5YkeolT2KfXybfDZMucv++FH
m8ZkUgHrmpmNbfEzDQrXAKnaejrcYX+wMTmHMNc65H9qJW9GhEVD6XKolUGk9QrWQi9/O3c5dNUe
wgFXaLOoEXgFhgSe8QOgCnckOqjrJrZ4zXGBjP6/4Lya0cIRUXVwriQBub40et1mCiIc5C3tP6EK
GSb8MeLRLSbrW1urSPqWbz9Du58nlh5Zh2beO0WBdU+mcuO3a8smWieltsThYr8llFRQOuh6gudN
vizcdnG18e+BVJqEFpkMR24y+MlZIQaysZXa52EuW9rhInNm86bvOSe/boCaBkDgZa4fKRrlQT7y
5Zycc81IGGw9NW50LUIlwAUQwWuEErvxalRczfmhLNTr4YQHusZw/yoVtD76kLn2+O7ng2gM3G8r
dQ2t1S16skbU491LTz9YbqSaiR8b5mQ//9c/VVDQf6nwtX7fiWEIxR/vItl/m0Vw2669M6LsDP+g
tGBoFFNIisRnGkzrpzwSAxdTxJNl3c6H6AE/p2+Rsc9/efNpSSAIXAhaSWtBL/Ngx1q++ReOeJvj
5D3EgJEE3FKB7Bn2fnsNaAcHjlmLO/hUUEfexXsSe2Qwu+FC9yh8O7j2T6YqiCtqMM7FobHjJ3pV
PDQLenr9QyAfrU6IP9+3pvkVQ+zrj0Lip7jxxAl3rof9VbQfb7cw1Api4fb3c7628zdwQllt05uu
68+iyGeB4DgUxfBvtXje8+a061fUDtw5CxedRWqvXlqc4hGcF/i8SMVUWK1Z4W5N+ZbRPg0yCh/l
qwsKNutOdJyIHr36VNr8LwjWu4b8yMtE6u6yrLkCPK3/TYxQ2QU/p9pjHPuKiSX57Hy5TCNUUWl9
JvQ231C+sSrlZd/mjiQQfhLHAp50Aya9zm/UCDYodQWo0fkIuTeYWA5RVf2d8DA5HL7NM2qO99OQ
OKPLNrMAl5UBP/eLE9Pit8/8DW+PPahLqam4MjFCwHp/1sOOZJx0WZNKYfufm21PGXCcUsPPgpyP
eSoRC7W3MnQsTpqXsJLNYJcPsrPxdS9ugDwBJqEuayknOqZ8a0D2WG5uBx4gKNIOSMSJgF+ZWmsY
aQUrmffGMmTZJGQdyXU0rkqY6B4j0bsoBpaL6FhXAeuMd6dz8TCSi2SxmmKebPg/8u+8DNCVg5s3
qSmo70aiVaEnItOVFeeCL79EjJqKAjkOM+kiu7Fy4RgAFvex+eLMJ+4rtyt+2SzBpE0x9cLpAgWY
EERrs/In4M2/LoqTvXaQyvh3ZPk+G9BIXL50abIG94iuPNlzScCdDiqUyNsdYTIlqLyKKXaf8iDs
RJHg8fKBxX3PSkmqa+cufH/fcBPVy8I9kgUemXbgyINbg+Y7P7OnQspgl8gblztTrMJ9UZw8zP1U
QlFmn0TsZ821twCyw2jutSJ6gYWOtSh2H4r5eeJ9v/YX6KNiZYLpvfxsd3l9j87dFCzF79jonUBj
1vgG7uKRXOM8sgnauR+241RTv9XxqE8tlTaPWruTaI+9eFQMHpmwIltrFZNl6RxXZywcTY0HYKjA
esr+tut940x5NXA+3LYTyvJ4kq8OEWoIT8qTVLqk+nLgcIy8Qg0n1WxOtC4uu2U7FX+1Nye75OhV
QTkcurcexG4kdNz3oAx93vWonYMA6PqjTLF6ybo77MrBp1vc0JP7iHL+6mAzTeTYF5jWvw2VgHmI
bgIG0l3m6HdmYVVTaWorHMVk8/37yq+recpn/b73a8tQI7HovmSRXvx9lclIiN4AvlwowyrdOPP/
BRCZUu7cZqnU5NFgVpH2pykTxcXe+P4AkXmICJJvpXnm0hHDEPHuTE0Z28CmN/8DMd2Fw471H8NU
TgEKzIe1NKTgbizCQSd9IUMEV/M7P7pVNgSgpZqa5h/kB/GVXFiuZs7FwD5NeFGFuspL6Drzf6n6
k2ymVWfy9pjWFDMEZgYFzx30grAr6AkO3t5+sm0oaw6AzMusV6GQK9gjIleEDnUey9cFi0a/fkop
OgzZm0LKmGtFDUBHPSfqE1fUk9td8J9+DV+lbB2LhFL2m4Quq5xjt7gtF07wyDLBb+0iwD1l9tsn
gqFQ21FPG2fmWMdcThwuSf+oxk8j00fVFYJ9yMDsSEOguj9DF/3sbuIVYqc4/UhC6QGFByd8nnYR
QCkoclDEnb0heWkfBqc1VsBbcANpMO7VbxhJopNoplZLQ8ue6Ye48TFnnFNIRYrrXQh9LWIua9sr
bIGt90JMMAGQnNTvmKRjJCxIo0oavqTeNiRZYTOoeQUdx4r1CEtefromEVz98KG6yueY7rqF49fg
ANZyalcquexge+A13YGS/uS+PeafPUiLWBRBvQnsJvaeztyJwjoqKz2kza7a7i9cvChb0Y2ZtVhk
9gsXEgCdrabkJIv56Rv/rMat9LxcPRxlIMaJlDOzv28KI15YxgozEwVAyhalmr9/ttE5uacNEGxg
lMpVtKLznKLlMm+I9cZ0sYfJsDCCHy/P8MZdyNRdhAxheqrbKkMGT67STRpfKtlO+tZiSvSBi1/y
rdX7OU41bP+kTdUSBDzt+PXqfmx8vxKyBJJAnL7C17FDGy8rZXiTu7zr95CHjQJRUyScKguzgCy6
NrBChcB57bGfLJGaSn5ZQxONHkKUbdoAgX1S5TPanMbY+lyuARZucBWofapaa6KaMaa/cqJuTH7d
8vC9tK1Z+4qvf4fuZQuRxRt9KNj0Llu/C3khiC9iRbvrXAcI/KiJkCF/1EEvWcRjBmPHeHnn1Wop
xgIWWW3+n+/4E8mmOubDgjA0Cqc9Gb/A8qIjkxb23ARqR+CgEby1yQPNYHGDl0Ksca80sGgJQlmJ
rkWdlhe4dpNIzU0FNJWcN5CC7GOgnz+OoqtU2XpGUjNgDbzFsgMJdhgAudk1jB+TXVAcitabwKjn
C9GBlSLHGnxWqqpd5rKoXBZiy2OmhLDZMJcokNowdh7NPUyOHAX4DCYsBerY/M/x9cXbeKBk+rIY
1T41N8mkx/6m1AllflQACfM14zd/zv6M2+D541amqBuwolGUpMoCuBgQ9n51wAYbKE/uFuOKwpN7
D3RuMiiyXPZQieB6kf4PNYP8CIwBg7dhbAWWYK7lxInq5wtujyAErurArJVl+291q73LanLV4nV3
dcXbh1jNexpFmvKOl/IueeMNs4ZthCag9ImK8ZYGzJ/8Rl1J5Ay1t+Vy+DnbI5W/9iM7T6FpkQMp
3V5e76f42FZsNiXDun+JI8n0DdEkNWgom2uVQGh5/F6qyNzKI+RWl36cI+Dr7K8OH4bYV8YDqg9N
u1BxfFNR9MUn88atpo3ST6DCTxLwMBwmurFwHVPcy1C4LiB4QXiGeEbFOCLUY/vyDHN0m7ljpoPO
tH2X9gr7XLEKJ6J1FCqS83EuHOHGrZxQ6cxm8B4Ygqmzg46znMb3xpJFcCUcG2riH1rKkNnQhHvY
MFD/CcMavuVhBLldz+GJDYHqRFvk4zWKhILbZ6aCi3XpfrJl8F1DAdTZ7XlloyfLribNiyZOyE3N
mOtmjDe0l0ZHoVPFwnnyegXgDPW7RAm/1Za5SC+a/8p76un/M9cUuBqQUzojkYkWH5oT/2Phfoy/
aQfRakFQkzI7YRkGXywIvDQSBk6Km9ulDEXWdgNWmVRQehpBfr3QiH4NjNpie+K14xpbzPdGLzz7
ymWmoZ1c4zKaD7YTw5J7fEpFxNMnNj4uUUKAo2vJQ6Sn6HH3eRM3hNyAqfue06Skvs1F4gMkpkFq
2rYxJ/xB75Q36qZKdV8cLZxMw9xF00xlX1AVy3Cc840DAbRTEOxOQMDFbe4GQN4qQinIJhYdm+KW
0y4DS7waH/ebxfYUko9guV5Zbn8M2uCcUsD/pjdnUSTkeO/jICQyAW4Fsbk+ReXBz3BKh+RjYQ0V
yf4L3HKFF9q1FK2RKcxXdO958TL16ApbDC5orrpQOsnlzt2bEoHXCJkuSR8V7llUrNNHJq0jboN+
jNPAa8YwlWEKD47lSoxWFEyn1idPvptjs28R/IZTRSi7BXkd2RaB8/ud/VPped7y6bsUGevIm3ER
ogAY84+iHRXS5YN5BAG7yGT9tAnaebxHG9DeWTieGuYh0ON9Y+JgwoM4N9vKXiO4i5oHN57CvElD
O8qcmFq0x0YtU151eMxmWYNkLMbG20C+bLpjuNOEolJR0eYbgDotiVl7ORX+6ZqRJMx1bDE7HTDl
b1VIeQdwHPqXVC+LZfgJ5cjCpWr3wX0E0vccaUqWELj+7NOKRJTB4MmJozjE7tacjxnn6UCebrd9
jTQ2rwEZ8ZlmkC8TFRPT7aMk7uMjNAdFPrPlYYWW0tLlmNLBsATeKrdxtnQq9xmvQmOejPzl7P9u
+ntsclygSjMIIxYDIPQ5OO1oE5oigKtNbehKWYr0HUsZqotRNIKRaI2LN/DxZue1LwUay7yUqk2K
qjIVWd6Xc1EVxtZnCJeoEZJkIZTFYHSnHv7ahXU4cNecxtoGihBD+mzZY3BqrU6y87j2xPhzW8RW
8XsHhMLBboenVB+nLnwGVdRefdr9tSdmEXUpdvohrxLYfQr2LFYDxKZ23MMZKDlNL9z4ha3Wo947
McOC/ept0xUQMS1mjByrhdTvoMlgOl/B+V49g0VPSh/gHVocJJJ52UsycD1wttXG6YTdJCtPqzaU
3EWsaQdflBxuDPm7VD8FGGO4UlKCbxy+mqjvkDX9kutP4NSpFhxAROou7CNe4reReOJ4n1I87zah
1fBz8GTRUKaMcliuzOjawR1CG+199S0YT1sad2XaQ/wt9EvVmAPqZP7UXlz0KWmJGIIDjf+/veSs
WApT0lOgYyCRV4J3vByZ+ZjzAib7SSRW+9OFqSWPscsmGUjXGrQKpPQZ2ov57lJvHGtxYPEq9873
eb9KIauiWrZnzAb4TfL0aDBMTtil+gmVkjjGBMPDjLu/QpJf0fLzMbKxZXUpmINyHpOnHNpm4hgH
Ntq7K9ZaIylFLS9cnwfiihFIRr0jXxf1wnSGDlgyPitw+hUV6vfHTy0FJfDdRgY7mTzewTJwYjbo
NJFobzP33qyn14fFJBujUauVjx2yC1aS7NmAvJzGkxm+Jx126FsqG7vxdKNcv7yJoOJuorCH9Ton
kZ9LCOxWU7umm55KwYbMtCglkhwU0FTg+qp+fKXTx1SHIqQfUx1L5qZvAuYRxu0CU4nzbPh7xQQO
RLSpZdwMAEKh2lyhqJlpgQB19ZjQyig6FqFDTwSDPpVxUtOGyMemfLmUmUON37S1JBFkuPDge/SE
AgR5ZVsdqQZP5vXMHDsUtjr7nwDu1dc1bvzCfyO7skKP/wEiiyNz9jAJ0NOwgRi1D2YmuDbeRaUV
5VoioFY+AFdqSszei7n4TQqSs/4lCmlosibGNPBd8FMlySnnf3pYR2gd8VCFkoSuMgnluJaI2Ikq
+OEQu6h0WdIB+r96dyQnyINWKFNk/dTqEBU8NWLNRWc8vZV3+FMM9Fxi+MFlQkXrmokQsUnGEzpq
7pw9YEnQcUs1IiCqnbcylb+CIEiFsHatarmRPeWMWqVDlM4OaMS5KJJhhDNPABG91HyihkgOMX8G
deyk2df8WfTQwkOyuhR0ltSKzoLh6shbLHP41IXa43o25z6gZvC82CbnM/bwrlGOqc1jGu6KKnAB
hgS5crUZOWEJdQCJpiZfXCBFOXZCaANl/vU0x9WaKNoQJe9ef2Wf02i93pfyWIuYLQ6NZwCop5Rg
kYsyz/qCyU4FkzuIUOk/W8czS8yqF0L3WaevquZpceVNH0UN7vnVW1KvJLEkFQ0OD/5eIfs5vwIn
388llTZSe+WRjuZDHL32FcNFD3TbKNMnwdlwHMrxpwr3tB3snA+PZA+g1vlYZYmBtNmtbSGV5ozI
FuC+P831Pi9B5o4qgEmJa0t1Mi0oZTvOlTBkYCw7iaIDyo64oJG4fCBlK4NysHPomYmQA7vkz0JX
6AA5O6L5CYSYMPod1vWcLsgVrK8C7qdApdAXjqhA5SUyepRP2Po/W/dMf7WIJjIXsZm0ZIyJuMfT
URPFJH22oZQmE0A+CB9+wjDZWMwkwe5jbeUNjyzkSVw+OTdq0DmiEvyqCTzY35SNIcnFKNmO3LOO
gG7k5iT/+3OjbuxVC1/CF8buzwd7BZVhNfs84wDjpXtHbmUeSHde6MCY2MnLgk8TstcUP0paTYVr
NVTXEByQgT2hb0WslMcvsX+vsDo4v91ZWGk1VkETQg4euFDxrYMV06wYJe6MNQjFx6B50Co02NjK
A2nBKqOzAJ49/BWMHL8A1D2JMnBBdd1hZ5TKfOYFSo0FQWpGj070uz2ixDAkfPy/kx5PSYavZlIZ
hcvr7a6TKYlXAWMhFFtl83KMOHDQd40gXN6YgqZG6NUWqf3XkWDfzyoUeSFrXuciq9K3d/3PrRCX
xApFhj7IvNeLW7eghGrLL3Rj2GdwbDqkCokIatlSsq5RHzWi9746m6dW7nM+SzNnHCDQmRLm6qAi
gm1O3vrbGKSu2nDDGEtW9+JsGvhIx/Sy9B5PubhcOrVUGhzigdwM6czrFzAeLjfZAjroH9jIoJkG
mxm++UM2BBdJzGEBBlcNuMYni0czs6iRECLqI/BR11cqn/n1j50jkwPNqzzuaQw2xBEouTpx8I8z
ttBGjBIW9UE4dRVoJGR4swnjlrN+AwYMmqX5ZYnm+yhbS/EXd2InMP6c6+x2uHWZYYEKTmkBjx4X
M5PVW+I+C4+hN7ueupiGxJlhUX56Y8JYjZ8c15NmzHfGGdGF1cvQ2K5yDuHN+PpsJzTZuZ8Ku1yZ
zMNSj+It4eiG6r2AqAQaNYE3axZiYbt9Q2+FtkmQKJpgl6rF8qZkWUmXaC2DGHLTWJSJFAvVMQ5s
IxAPxJCqSyTukJjtNbTSxT6dFn1Fhzo7YfXAXC80YRnhltsh7l03K+6nfLdVAWBtPlCwH0tFgqGm
/XmjCbtLm7LKzjCx9EtGu2hJyLutCCfEz7HSD7myyl+jbk8TFRJ06U8V7ce8fhFO1AkjD3Rr7noq
OePECtUiuUJEBG0wE75L9kGNwyjep2sdg7/xSwmA1afCHfHlZoQxR6nOns4A64xQxRdNK0rrxXYv
Ytqf7OuO9srQe6FSpXHGDb13tuZf2JMjxlgP0ADSeyPvxJPralq7ppGP1SdY5NAtNYyUeZQkQsfn
Hb5/6y98elog+hZC+9a+xvzbUE7OfZQ+d+DVlpCclZCmOleejr2lsvwAuj86nWs+Ergtfuqak8K5
Z3SsYxHZOGxkeJhxDDgdfgW4uBHvi2qI8eYO5NO6S/dUsyz5XOQ4C8m63P19yWhPsKB/LEa9Su1D
xrnkntjtBJ20I8Txec4jBt/HzmJfhS7bGoaii5x+UNBZzEnDYEzHDR7TxxkvGpQCN8lYBRCi2wQv
u/l/a2XHCE92Pnwh29hsiy8ycTWvnu2ihgTu0trpRBQteNnW55tnfTKymZBS+TbjQpAnjDgs31RB
O17wm/1RF6En3YoDHOO2XqQ7bzSr6iJ2L/Sb5o/6vpAKYO00B5IYN1/wI40r2J63bDfkvg2eiNau
sUlqJrWMoiG/cDdW5nG1VJEEfjkWsKPtLdXNrjI8Hu6ZQzDBG523Bo0hxwFaYI2/hEvabMoyJ/Hb
AHYnCspaugU3VqJKAxleOhycK+IVrSANJAl5Mf4rrPZHH2QROF/DZpUFqPKDSNU6gqbi6BV2fZd2
8V6XthMq/F3fr4YYdIS2EEf9SGBWwcUH8XY4MfhZxn+DxJQYpvX4u1xb4nba1lLu/3zYwMy/IYuD
wxBglcyK3+QGRODzYJuxGlliERddOfrqbpWa/T7ojefQdgrqRhZKtSd9Y9viDnU43cSCqKRjAKyq
fTBtoNmRPz7j9jp4rgsqz8cD+2+ZfZUR0pzaNqViJV4fEkZP7QA+byx278RPl5UjL52D++Xnr9cm
npWmsWsN6RrEF46dtu23A7z63s6ImkgyElCzeFa9duGTDznWsNzp8oLP8o+cbeXsGCJm22970kKw
DQUQc8qeOZ6L8g7ywN/pYdOwy+yjayl6pqxfLK9vUy3xijOBJPBkFIPDu+hmVFhmKX1OmNleua0q
NDm9n93CD+dCCuk4SSHiBvjmI/NPiaLsdVFXtvuUDg29FlTz0Q+DMXgud3KVvepTXvit9/Rr2UiE
CdqHMBP64ZRG4uNt+Zf8CGn6paogUyZdf+0L2EATngKGjExN2xD65nCug4DHDi8XUNIuqKIzGRfC
aPHKF1dVpL0T5COWX+pzdnaxE97ju0gdpGB2pyJobF70xh0CHh+iBmhCIhX7kd/nilSF6OcIi/wT
d9NkNOeRlv039b6YllKivCW0olJRlevrrqRLua/hGt/AEsap5JD2ZpGet0YR480zY84QYaFEj2em
Wtv0bboOhVeLKnqrWEDAPIaGlYy/MmJ/ziv2f6B2g1WreHPG3jw35nO2Of6SBdTuneNo8RNODp8n
tTvi6ATaycZZ23q8kZCJvQ4hxwFvNa1zOUFwpt6OQsEpHhMpmcJBPfSIb+P427Cm50Nm5VRGC56c
w0s/U3YSJmOIQ8YVZKfmp7YODkA/jgcLu/dHusWEsVgFJVlBdV/Yu1CAGIOygUyu8dNbw1KQCrnU
Xjw9G/v+L2fPUqHRU3Cbd/+SHVs3ITAh5mybnuZpZzCRT1Qtb8tddoJH8IkXZAqoyZX9+7t7kyfG
24BFfeIWEAUDVN1HuTSdWZ6pDUj8c64r61apXfBFi3fFKmd/xz71a47bNZ8a+R3yrC5aF2sJ7RIo
5L6EK4wQtrVYZDiOR3eLrTZwBy5fNJqMvOlU/+3xzCgj+CJj7irqJOK91vWYWegE/VH8UcLXWufC
kKbj0YTf2gN6vfFZQ3KLumqw5q6eY1hA96660pMMH3rCiqFYi//gOcXxdNwUSdlL4K7cHe9ijp8c
snU+Sd8esCAdPvAAsLWIYRuclGH8Bj104ghIvg9AHRx5JmEmIJiu82hjEwtvvbxxytoQoCgVG6tv
vmr8zprZr7cgnDjhgjybDQsorwD7M0IYYCBuyK12SmDDlJfEfn0nWc7Wncmwib8+sGlY36SEL6yG
YQO4STM9sTxFabApzkit3x1x9NWI0UDL227eDxqpnvLECYnjx1sB6rKIZ2SPMW/SObfwF954hMbe
7xuBgnfD6zOHKyuweXFWKt5ByZVJrNnCH3C1sHOzweDP6X5TmSUBexexm4RKyEp7TBgq+ZutP6I+
jNs9xEZjG/oaMwWWj5qzwKckvTRE2VVvSAtW3MrOtKfTXDx4SM/yjLn/5XoZFyDoW6ikBrdkc6sS
ROgr5ayRsYechACjyRcbIufDVQSxUfQe6TNp/Bm5YUKfDuET2fP8s3TQat2i44wSMZJ0mNGz9WIS
xDkVwlK6PqXKi1K9DotddVbDwne9NVwz07BVpRF6Qqh6crzH6Sq05yk6wLR8j7UbDG/ky0YAGUbp
d4xy8PmoZ1lb4WLAQe3dn0YF4+WEP4oc8wsLxpvBxhOor82Kgwn3DoXzuqEE2WkvdLu2s0MByhVi
KenM+dg9LHOYA1BcL1pP0lfukCCmsQg+i3rR1y4edZxVfyM+HxhKl5lYwVABeO9Po/zEqtQqL8LW
1Rj/qJFKbbuDFIlxG/XyEscAQ+a0mAuEMAOJvvbdbaZY7/5vr2djelD3becFH4YDXXKx/MXO3N9J
mAfKOSXFVPVcrykrygK+pRSTciUnl+LciHpHg0MWa4pOdw35A4OJYIP7RxHVQ4Br6NvpdcPGWZw4
65ium97ZEcVJtLPkJS5V5gp7iBGJZvxq5lxGjBtTdrot4KEAzYmsCdNaNi7MKqsaZ/XHRqu97IBu
twAeNvUbw0hBEI2cyjfad9Kat6zMtGHKwAAbhe5saaQY/pXzFvGcTXVU+qJUuUXhxeUvsGGC9C3t
sfkan6r1R+fPzD3nW+rGNwrfCAg8RzWkhWER4Jz7WhzdnQ0t2pmWwqfaW845XR8x9mfsf4z/22xE
ZdfYvVD+yTun9Z3vbwk9mfHYSMi9DZ4jGQ+P0ImhHmJpJdz3ZOIRdxGKKg90dja1VtbQ6E9aI2Pi
O2el/PUWJXHrsMuyxZkDzFPkVHHrjXzUAjqN9tgf+6T3b5Za/pb0GFYFuS0XGGCIE8lK7kDrEXgJ
bE5jQzroyd3zANI7gjZ4G/ATNZ/UD/INsI25QUcLy8/Y5Fd0XfVV2b5awC9VVQ3xFaoxwxsFhDih
FeexccXuSGvSzSnUR/9e/E3x15qMAaB3SQ8/bUSQeY8VBvI0mRKGhBdBaWQe5xE5KR+yCqMQeXZ9
IN8GqQYczwjQCylSf0rP65N3xF/hRlmUxUEZI7PgNp2Ud3CdI43BwlmNZpWZ6Y9DainG9claohH+
oUnEJsq3GJZmIUsNIorocAbQPMBLDIfVlI8DWhH5xgmMYe8mJR3ewxOSaJ6S9idOMgjjYdzpjzwq
b2Ral9zamkYXc4RNaSzlbEvM35VDKzi7RoRlxZ3hjUtIYX3OUp+W7vzTGPxtYNBPxltL5Sjqwf6q
wv0eu9Z/DI4RTjDViEqoV7JIZS+zHBB/YWfMJI8CfveKMyQazuvPXCbd5Iid8d+5PRvFPyRRv2PS
wihGnQuQBpZd1XYKa3Ott38ryPlRxa/HM2OZOt/byhibtdmJksod3ExWU7ysRRxg0u9pHI49oQ16
Rt259YVgCmvyzZhFLhqeoshV1fKCpcFwjzH42JVALr55PYjX9kyRdg0PPp9r2I8e3gadFEqC5dRT
HECNQReYyHVV3x1OWF6ii+osFleWkYkES3WukQASaIt92SamcDNCw4nUh4wgMMgFbMXnF1Xd8wps
XXql8gjHe+47A7cQqR27Yke3y1xxoXMoRoW7vFnGFTfIQ24gsvKwGTvLzwhxM5MoH4wNejP38r2O
tiit9PZjwEd0emp993Bt78TiLVNtOlsyDLoZNjuT8a4XyxdPlt3LOqAkmO+yZwLb3vVYQX+iEKc4
SSfD3AazHxhnnVvRpBpqEBRKgNRPj2obWUbDB7sR/vnYfhZ9Gb1wJfQNwbyoL9HCF2ZP5Dc94l8a
99tjSiQRu15bOU4nh9IH2zmvQXE1l/MFrefDKPYlXl0QFKWmFY4En5JqCKkwBwKO48W3FsUzkCky
n2eJADvpkTQUEPJKbqdtHvWHnDKEuhg79nd9MdKXkSDs+mi1/QML5HLocBIWZZjGU5bNVM6PlYrG
N9hCoRXIweJvONujZ8FU7MTRd2bzNencaMbpeDzMaxj0tZ7pt0ETUkj4HM1JQzudvEDXLhc2XI0r
tJxjolgibilnNaMgjiBRbveaX5hPUoACCZzoVvtyp0wwcv6BeujMiDTGlhrEXPr5BoJe30O3pmp0
rGzVgNezAJDALRp9tfZXgu1G2E2mOb5dKSjHNeZyhhdx1N5yCC+D7mo5d2I1oYQ6rn4T/TfrNdYt
dmcaXGURa/hDHSkyAKErwxGV96CwkEM0IsQF8pLq5eXNvqZiucPaVsmnyxezTs7nAx01u86OiXR6
+CRpTh7KdWWQtTC4lA/MMFfGRnA5bP9k1W/9nNtp/dk5LbKDMAJUQKWGRI26ixv1iK7edzey7zm/
VZ7bE5+kmCP0h/nFOpCwH7kZ6AZy3lxVLP7G9pY50A9TV+gD3EuAeV2dZSK3oXlRByqvoHT1P7mS
ZzN1cfwWmRBAQ0lOx9BBVesAZPd7md1rXjwt3zcofJEdx8dbKfOHTIUUWPYhbuRatRFLCunR1GQ0
jp9H/vJypmlK6/IslKA/mn2xu29YTXQKVX1/qKV1tPaSfePYck/3Kdobl/O7AMpM7XTPJhygeULd
zdXYs7iEoxzbphXJTkNx4MLXF3u5YhjE3eV1n73I/sHHiHm1d9shKlHMc1u7elCjCXfj+ARbknUS
DaAZyYIFJ8ybOAkWAxUIEBAUiuV74uYixKLdJeUsUEXO/eDAWOvgFbrLwTd6hFa2EOqxkg9QP90E
e3LJZRYcMDGQ1G+KZctfMgNx5w6x4zSLESgGforJ+uGxzEdEa/mv9lmZnadZVeX+zOOUvDfuzuLn
r9NebFRAPrtF0rrxbJ0CjZQ3Ptf11XvSuFX4rclK1HOcbksnPqfpppIcIS44oMqwMhVkpYg/ati7
v3FVfkDHRT0gFrr7FAMc/feNZ4p/62KwxmyEeO//Y2nsgIYo+1OsxTEaTU2OCNr8Vl/68LAOl0rb
1XNlqCVuA+BVo37fZATY63KpVVC0OrV9FaD/Fz/ZfMFbxDoqYpEkA5yLXwf5fpnEJbTcohFDNkpG
7Jfh1wEZkqCYH8dQYxT9JLuSE/nt1g12lo5r/tzJ1+Of75z5gWekvM32gcbZmlmVi0WebJZPySVj
YuyMqovy/0lUTOFdGDmuFpJ5abasM3XIpN4ED3Da9cLAoIQpx/2ADiWf5FUTo3ee4+MoK/zRwB3Y
vp09MsXk6fptaY2lLVLyDtfGM1knndEQ+RwUtH/a80KEUOx92H12nSnycXKQfK7QQKEpBeWVgYIc
3zCX9lIYW9Drbf5iEMnAZcbG9bTEo7b2e+Y4cFwza88hUZb6KXX9XJKOno93JZ/cyzixYy+wUoF4
6k120zkzp1o7EHd3gvkRP1QJvB/9fKMMkdwlYsoVfgHrMX+cc164eqgovShrnaBICkWD+YFGPxnx
uKMuwh7iSqtlPjtt7EIrPq6udSQKcsbs7VDDux9mZbwtQbXw6D6n1mQQ+e7s48/JB1HV+fQkmvy5
fuC29S916OZ9CLgq7/rStZ27kF2B1xHOV3ZPyx+ANYYivZdbDMlPHzk/qyZRNogDUeucvG/6haW7
HkbfR5mDdSygODGhseQZdWYU0oYgaIBLzPkzcqCbfsZhA7KlFyNui9qthZz8QOytwFb+y/f8PQs9
uzmSm9sXx0SlVO2Kw0/kEkvdyiHYfmYlRg19CPxLQ/j+aYsDTGA7EsJIvMAioLZS1hNbv8YhecNA
r2og8DqmOG9KqmN60E+XHvA3S9Fcpt+/oVqCSEHbecjJd3XRd1ix2dwArGO0NhTpTa2UHfUBSOTH
YM0Uur0nC/7K8urSBfJpzvHlya/TywzxNWgH8MNXWXjpCgftbIueUfHtC5l7v2p09hd/CgX/F23+
Mi7FXpBmX74v8H+kClTFegOhos22CCTOqPIqLc5xz4mSfKv7KeQrU/WooAwnH5RZ0cRN4nPvwpZq
M7N61fKnyKoD8kj2+qAkA1GL3nOh3Ajfc1fx8bjlD7dnN4wtD48sfUyB6pIRLAVfwL/XoHVKIh8C
PSwqOx3GhrpP4K4ozjqbDpgl/yVUaWYtbwl9DkNFI5vuTR0cZGIMma1G+vpTWF+evo5dqsiwUkQ3
xh8ANUrVtJhpQlHoQ3NG4t1BnzGDHYcVhdbF67LSOaA619JgkCLfXmhZGgh6VpRTnBx1irWf7/ON
MKIpbypjhettoXhaKassjwkkZCloF/Etuop7lzfDU2PWZuSMei9QI1oMsaYYbD4Ok2dN+ArzCbRr
xDBo1A+IkbC867XKRp5Ii6Xr9iJoYMoGphqd9ClumXMe381AuuDqaVAFDjJ/fDlAh1MQfUB6JmKx
okkkX1UyZ0ZNLyniGKXWMYEQ04qPE+gy5BMZOay57AMcobPoTjZU2u2nxFtyu0vY09gT/J78oQc4
4gkow8Jv+q0vsRJ/xYyQNv1NFLD52QLtzHWQCotDvURlHE7dwsX973+LVA1Cuk/kA/FqEy0sPzJs
G1t8F0ANTIyt7KeVRLCxYFa/cgOnbDRl/Il4ig0U/UELQln2V4i/Vd9Pj1UQHzHPVCSjKeD+JFcp
r4Xw8hcwPb3lkab+LJk+K7Fx0/NvwoHORIwfOQZ3kEQ/BbeH26xddgV8AkoDIHTARIcD4T2T8MAT
h09Yusb7xRuRR79XwX65Pj4jStH/63eF9rqqc3kcDvqsIrIef3UetihZjlWBtp/RXE84Ncct3MMz
nReuZXKAkidS85aFCKcwlYOKdbZEb7ORoq0oazNpeEAChba+SBNfzC8+OxaNvg4DWK7aWo7HIvS2
f4ItkVgGxPIhhPhb3ZRzUvURCbu5HOgzbVidyV45QoTF6wZn+wM6GG1aimsfx/7KvSL/ZlU9P2qt
7nLNN4W4Fu9hXAi4QJNnKTz/lWiVn8JE+qbDbzu9OK+mK3yeZ3BWiaFHSxip+ldygG1KW+UXkgPP
+mXCP3Wbsh/b5rrQ5Id+7TdwKH8XtUWQjRE3tm6Hyz1Mj4tjLgCI4YbkLG2StJssF/ZXJ7gmx2gU
GHW/KDF+wR34OoiEWvJJePH6nony2LPO+f8oO4sncE/ewRqevwaRbPgI8oI/Hp0spEKaUdHC4Awu
oBkjZ8/A4psfQygUDftnGOJWcL8zjQSbYP21PxEwi9V2qgiMmi+t+xGZ6RNbsGesn1mloxW5lzi5
2W6zf6evxZcVL//ZCiSWcMg/cJQaPiz752UmPRCF9k/oaXDbIeWHIpflNLFO9333vz19KIrWh7jj
ePLk53gJ6UTsIJlhI8VytuGxPKNYX/p9cvA9AH84AzJw8VXmmanhvM3mfIYQEsGJND07CTcLLbKM
DMZe6T7eMGmoiQWjR19un6Hgf2fCrSMLz1fsiFCyVxuBdu4bz0yc7EzSQ3ZxGg/OxTyKdxHx02O9
W19IF8N6K4SyLWW6jJ5CfagKhBl0GeWJI09SebMj06+fY0WYyUjqCeivRJaYRATehgAYzWahCjuG
zDmajUQlMvstDmU5muETu7mk3cgAX/fAa/tvMwraydQt02+z1zO0DkGJwjn0srlTd23SUaAsjE6J
BrVdCKjA/7OSfTuPrPBSehaag2h99VfI6jbdEYu+7Y85U2JiDssigN081V2xF5V5L7DQMTtVPPfD
o1qX3Jvk2rtNvU2bbGFhh99K9+ezaTKZD97dEBOFiunDuTu1188q0jf0+czbpbZzcmcXHsVT8OGh
iVtLCdrCxFLkjN9YLTvTroBc8cc7YTsswK+ZxuyzhVMCdIP7BxgjIfuZIXihY9DoyQ0/vBeyFMt/
lsH98Z6iCZ5/+h0YWlqu8tlH86bXBnCXAcpZAcf9XEYLLqhT5gEXWUl463hpJiKyCDRMnTZ3w2Rh
mNzk/f8x58canaHARcmwrU6m0JnXWHZ9GRP1ZkpOVzeDUCcJkkq6+4/DCgUrseBdOH6o8zJasNs1
rIwAg7vW/VYsweK9m9qB5f8pnD31QRtSck96xTzWDEUTIsOPgRBwcBylICoFK1tNzAshzyGPML0O
P6HzeaZoZSr5eOHicBxXo8gEnhe4wcmC2cH9sOm8ZZtGuorDvPAhs/Tlr9cylofidVaZOVwXBq51
PXo1om0E9Qs4yJFzkl5ohVESiRar+Taay+5tAiQv5Xq+UnRQhHmuGrBi3HuTJl/pfR5ReL/rErly
mRY3SzESq6VKhmjj6hpyL1pQeAqgY1ZiEnMVSaLyeuUSg3mbwvDPJVaeOIcn/Ojo8FW0BJtqb/63
ryAdxkNESPk6GkpW7AXwBro6+uM6ZrQp2hBEd6FfyrYAx8za2VBSecyr2FuSX/B+9ZS1RU8cFww6
NisQCHugOZUbjqD53ON1ph0+/9EHR1QE8UEqI35GekHniWTMiayORbRwWaTXuMQtxWvc355QOK/y
SKn3abVeG/4Vokd6QeGCndYNRKKURAN632GtgeY75Cy++Wt029dgDa62ek0eq/qTlnnvFvVhd70j
fRNa0zYDFKM1EJAlVn5rqLz8M/xTiWf2WCUqk5XIMnBX0ABScJrYi6lFAoZsL/c3diWsX+TyQcwy
4eHJu9p5E+WKg4cOKKcD7wqlYKjNUxQjaMTxS8HTbCy9NJtfvbhfZ6hs2MO6YisM2BbI+sYHDzj1
GcrADESEWltJQgbrlMXXXFMDLHpYa1DI9RJr19BJPjPzR1w3Lgkh4b7rRWSe7NatcgkU7JqsH1zt
5s97e8p6VKZYsKm+NDxn4vTUXEqlzOHmuz7OB9XBjEIlqOhi6ttjCwPY/pO4frZG7A896MmVf+nK
ttQXH7TPV1H1wFyH3x93R5jQPSMhQNKcyaLVayHpz76laZHLLnvNTVeqYORrEvbgDoHdNXDsNKHb
Rlsulsppm5CRQ3RNSjUnCJMCBHw1J1i/IyYM2kWcg4PtpXTV28DEUSqyBXCGmZxmRox4XF+aaCXA
eM4IVZKxyDgmMDFMnyJr/tO5NLGSwuqRvFZIXvG0DzvjbNRZsFHTxi4cXJXY213bNwkA1umTZST3
lz8VEpyN1/WfmvsajsjbTO3e3tVSjB0zQOhhmLWbldGhhCwxvO614kVJyd9X8PBLY+0/eOjzaiH4
1YMzM8+cKDkst3bY62NvtAoV6rSMIZy+4RdEw3oZOSCDHbarrFLqUdIESbUKfJeUrmgISujfXKKE
6JMjsnTX66/S+IFHlnQxWUN4cyur356I3s76Fe3MakgtsUKuRPP6E3VMq0VvM/Uj+I1EBt0KLON9
yl+1/PcBnmkNwAJnLVT5zWL9diOSrdNi8Q1ZazkZr/iq0PTtBG1D0tXLUMeUcNamEJ+29T0XUepz
0a4uD7enX8IUGKUJd4idDlb/63el0c7gH76gLBsWf5ly9T4yd94eWs/lMbiLXsjZsjH5Y9n+oC3/
+3BXC3njRnRgz9zGFN2JaDPdaOovIYRdYtIUb38JDzJHuuB963JGJ3Gp6AESl8IweWCpow7ApTwF
eTK1F9Cy2jO5tlk5b1CT4k9PmoeKIeecDi/FJuDXYZzUIMSM6mDK16TdS62C896aX8ml1QclrZ8W
0s3dq2sniTXhMvYLnU9k7tQ865BOc2KLwUMRYaDJl4H609N/H+jrYF/9bppCdqYGEt7UauOclXNu
XgmEbRJ41JWhzFrTN+63nkKvRJOvPTfmgSvbwMzDl8jXNmULLOO51KzD2qMRl5TAQq+uwmfH5wKe
vA9J2ViG8BYoYqTU+t86i8NT4mV5Uc41nc3pPlbxYrTc8K3p2WsKFh6Lpx5DFhn3P82vmhNp2ycg
ibZwhLyMqKV7lvup8G1wM+88n58OB4sdRlL9v1ZsZbhgNO1z8HkMO4+gLztnxdhDURND/cRsofqB
klApp8fsM2UviosO+I4f5wYxzjiV1kI71fxtN2rDQmpSJH1Kan3IYWEdr51WAVD1XezrZVKlkDTh
INOSFoFxxefAtpVKejr0veSdUkg0eqL4+wLexnVXA1yWTiZiFjazIMtRr2YcXU9oJHuvMMUBdWui
tNT/2SleNXFkrwb0fTskPrfKv1+gb137C/hUYv7x1IA8rysLbG4C3Oawb8ZFP61B/Z1XuPRtIXb8
7d+pb+TEQ/p43DAsClo93s3Lra3t1LgT3yjOBVOBRUbjt1iXDp+Wk1o4zrH6TAKum/6ZqwUvXlwm
yvFOq5w/WAyqte78qAULRDW5PkSYAUGfuGcO/FWKen/wnci9LA+Mbhe9rsJ7ZwwdsOEqGa/FY4qV
A8A9TvoNKCMDH8SJ8S8x1R8q+3YNMBiw76SAtgPmY3W+D9++lNnF5zmmaUnXpw6+lsPvG7c6Nc4e
FHS55UBJiSmfM5oz5l3hgiAIV6TKi9o6rPvu0xF2X1SFBnRKiohXYu0sXtBqY+Yw8JXHh3tsRygu
SHtfQ+E3K8yGKtUoQo/6kZy5STZRQKydlXfPjT79GZmHc2IbQPKt/lzzMrVapDAoS/1VoH0vCGNm
5GeL+yGqn3iaUI4wmE/ZOzmYwDMtcY2srOIFcRex4nJsk9hq0PnouHMLeKd6PJMKt60HbEpCMtLb
f/9edtao3pOsly6xzg9cTTQYu7o15vFmWcDfQo12VXiHVHDqAjAUsm+IjRYMy2IUgcFzwb7JOGKk
zh2OmmzeoezWhMz0UELOu96G+b03ybJNUeR6XcMYDXMeKUHFcoW9JIGWIuy1Yb6SO1vAeKS5Yvtp
NgXsCRTVlvb60FdirpifWqmgMEH2+RceSRW0T4zwv3GhhpxL8M7/Vr4EwgCZ9hOgj0djy7alRY0E
ogxO9n/ncSFDjdChraFr0fGiB69MIkDX0p22WrwhuXtt23nqBNccJUAQTxxyFxSIgLILHojaweIk
SA+SuaIFrqrqiJg25w6Sx44DaI2sLv695/s3ZNoxDGQMOlSbRgFKg/l7F6v7LKgeMtG9uE88rukR
c23yZJ7t6O60M+ZsZCn2YkbdwaZrj634d4Z0X/0eOvK0YUxAaPL8nrQOOXEOfWWMO4lsI05yzU5t
U+aEkQVpE6mMWZCoV7J4/NbrUn34A3gPgc9vzWgFgVPW4CpyWg4OtBnXAOBnCiv6h5xXlIXBsEp4
ee2j8UFPYmguKFOcES9F21vYQB11ztKpcJc9wxhafkcYMHBXmS/IavS3DHCBZ6FWTEwy7NLozFZl
FV8T8jPMMVEIqRHXeEfRJ66acU0Y2dULhaKvD1zvx0j2aU1PZezLYu/BKNoCBlMl63ZjsHFfs83s
o+uCYQxPvWLkIRNR2pXm0keCXrIsoJZnMYuPDZnIB9qnpVzoHk10Vzs7WzaNxpGd/C/B4xslve4w
FGt7relJVN0ctLTM1iTJJvDAT5wRCihpYdXwWH3x4QZ41NB9kdPoj23plzUcGRLzVpP31h8XuAyX
XSAaQhNZAHK1j2nLQch+jdhHTr62To2+ovkkt2K6nvjJhBg80ClKW5joYQ65nLhQeaF6uUC4C/xC
L04xdAbBMmmDlHQUsc8HE0nYZE7UZvksG3DCdSnDktvzSUUv9UmfZ8T0GWj9uRUg7olPBTn0wPrY
8HElVe+3tpf7FhQFZilp7OFagogLk+SyODO9fGw1U+juezktVoLr10lLd8+75+c7ZnC5covUxkNf
sasgA35xoPd7ZhnEAvVMCKWoD4+G+LeHNiLX6JDpl+/1jbNXEGwJslbCOla/Ei+0siNWjzj9RJWa
izFl4er6dyIDX3zf6yVpz7DRrr3Dlv+fmHw3iZCGbFfQd1U+KzXmB9POwqp7so6ouzSjDJ18Ho8S
OUUzr7chzilDWntTm8O9lt4HJsuAE36ELdrB52XTTJ4jMT441CD0mcr9HUGadxz7GAosYEi+IrT/
wjJcBt1qxKNusZBqWhv9vyIvCotu8DerA725v9Qa7zPBt6v5cWccyCi4nbPCU/9fWL3OrITr+zEX
yQh+9mpEXP4PM2e5l5vkoFFWON4IeqWQB9KCqy7vDNsBHkk7mLOgXE72seFLGZQ5/4ndzrF2WBhk
kBG8P4kO+7hjMHo8WRm2V+RPDnJDsDO1rEfQL15smgTv6FNibMF1XQT/ckSDHvhXAldaAJhXb0ZR
zvpk8jAjFfPGOmRJvN/An4ZDcWh6IVemIK8mHxBVM3SRhOy9ye9XfNihGHyl0h4+g9TL2npn/4i6
fH9TqEhhBKpT51LBTcR2T3jsOaWpvny5MATgjWhKOCO6uRG/okbIp8HhxR27gcGvmBP42Uo/bhW4
kwc3Tn1j+lYj/nRrYLM5h4vaIflMGvsLPzznKlSD+GC3a0rLM04MHwSg2pXE4WduL2lCcBrXVPC9
9n/jsnVccV7+cIjwJc/GK+aMlLyU7lD7C/ByHyH8CYDLDY6EjdMsG3Yyx4dpkbd9PZwt7opp5NoR
Xf0oQWnEy0jGowjyPRJ5NRTMeoLbsubYO68inxtSQoSMq+Bx3YUtnInKwKycQHFoV1TH/ja8jJ3f
AN2uMSx4Sj9Tr0L8giNXKixH2TjtBxd8WlT2Yhl2eyhi5tkZ84b4XsjUlOFg+j1qhzCnPU6I6Luz
FNvWjvYC0llBHJV19pdHlBaoOE1YbzpSA9iqcQoem3MHPWA1aiH++LFQPiKkBwOnZKu8AM5/QYxp
gmkekTIZqjFIawPdU0LvYnIcJs75Cw01aTkwMuPP61Tn0Pwo2g5kl6cE0Q2HUn0W2MbI3g6jvIqg
7mDsfpU13nzAIYJdeZJOrqIdSarHxrqcSTdhb681DL8pW7kGk6Sttb607IbNKkxKS8Re/StAHk1L
VaDT/y3vz7kSkwjE+HDGLmZ42jVkWoTlN9qa9VNWnBS/+EBG7lQ1ArSO2rOkugFwHNXWSFCJqNAB
XM7bxnbdoKHuUBNDsVWj+QVf/vIoNYgeHpRpLQULoy3v5csrzAWqhf/2NV6IqOkpvIcukUyXtsQN
s6u4sWhAhAzWPduuo6UUmq+8ylRtdW2Orop4bUMcuD6QW+t683nTWPlE9sXptRggmCPpgc4Fx9rr
SzhG5D7V+xmOjdn3WIS6ncf2uEv3ZMF4Sp3duixJmCF2VS7bUEu5kmVwsaD9lGAAHXaNeLymvttu
Tg9uGwn/cOBcH1qRIRs4nrakFjLhZfhjpSMFsGv8Ixh/05B9y4oAddnLXgPkIKhM8B32MexK2Z8a
NglE1rOyyt2ldOaIqUPlhSJj5L8fZnM94qX7CGkEmszsGbdeaJ4CJCq8l2BiSJfVGPF7uaWES/TW
3TqpX8KsxuP0rAUXuyi/mgw2CIdb3+JCypdWhFR9KD3Rt01vMR9oKr2NCbp1bSbUJNAwuJsX1IdS
mY7XHTPNOfhzp8ROU3yJREGNEz0JfUgxz7fN4WGRCzAZjBX0MsExmrIxFW2gUPwjnbgdEZTRNBWY
DJkQr9N9qr3coqPF4kT3F5Hcf8Gu/SdsRMUckTKCi0pJCdngZGjzdplTPc/jX6TqlodOeolnwiWj
tkp7VhoFX1xs9KKSutjFagIjSdztfxbgnvjOiu+cOXKBHUQTcoSz019AvlqZRzRhSSNo20WhUaWp
ifz35dNeL8fszXRDEkKmSCfydn+zM8BfEZvfMV/Tcg3pGW/fKF27+lH9jP2KDamHtAsQXt+X3HBi
llXZ3DJHjMvUk7WWy1izx0x6/DWbmRriQZZAuTYdvrYp+1m/LpXLqKSE5UbK+nTJqfiP4wagxj/Y
xC0zpd+ea7huXDpL5L0Z867rvSqBaCfkZZa04jeA6TE0EbNMdDGXFAhUqSPuW0GFRquh/TI9RfuV
4I4cG9+E2d8mbg17OSTM+4U927OUXBsNJdcN1zE89VXTEN2gSiS+N5BZx1dXqdPgraMWBmg6Iwl/
0aadljVhWP7YIH3XmKBEMDtMOZ4Rg+7Ory1R20LsFBoWcHcbPZzjz5rK0PO+CG/xmXpZDII++hkF
7xMfO/F2r6gqQCRbgoNPh1iROZWbhZd4XyHKQQv24dx0c5pUrdS2rODPi0ZTiz2cY6cnMPVfqQx/
VPYfP4n6wAdotK33tbJQ9620jmDnPIWLfOVz2rfc2uStccvtVqN+qzFoHcZglAOPmrHnlU96EJQF
irrHGU2hWlPEZsdwbWd89qukMn3u/aGh/Z8rlYw/RA19B/EPA7bV9c1b9JNIJzJ2NIjfvwqKz1H9
1b2k5pYkAMITC/uS2rz4B6JBdyhtWemAt5J2OL4BU46XNZ6imRwDZS8Oke5hqbj5GR4U7oF1DNh9
cFi2HYrhGlWOJngQa5nB1o0tv6YZWSK0gtX/FPy4bBEXLWbMdEQmtTp2IxJ/EhzrlxcLxJdMcaDd
lezOz8zc+tappeFHTLztDe2eGP+9tEH2gQokgx9oFmrEr0Pc8kJHDt2rGP8WzpVD2ZSS5m/zQ99u
4Lsv3e3zjKHcb+TIRC4L60kRENrs/0d/GaOwnrLYi1DwJwdiGBID5ZSNakvHkIGCl/i4BZhIsAO7
M/Q5VSIXrVL8Gcm5F9fpBOZUlSuLNL6MTKsulRP6/KCWZkNiXm4BU+DuhHw3/l13cQlydB5Iira6
4PS+0TP8qcQ9hFfhS4RwGesQGOyNkT66HwsJdv7E4hJRpZ/qohK1svDnoEXUGj4+4k03pw2aURfK
g0VdaZUjcxNUAmtvp1PL/kLANPwIQ+BYjAbvxuaiBPq08T7tZI4BrtysWe7l82jQZ13auq2NV7k8
O5nFS2t61fG/xXQAEJfPBH7ww6GrCAaNIyaoj+A1oNGwNH5iL48f6kM9ny70bagLY5Yjs7P7h5Ol
KSdDilmr75X67FJGG1YIjSxpSVEfTPVN/Zipdqb8qoknqcphrixeD9A8AdzyEkI4L7fa31S/7VcM
bObIWbslT8On91KbOSwrtjvKQx1jQCcRkqsGj0CJn0E1VkZLZgJAYEtuEUu3248pBkSsWkeovet9
xcZVZaYzEkKvtspmYlB0v7QzCvWsbUpPOtFY4WYhKLYT8WRmamNo6XLL4BBt+7wq6/0b7khwMAJ3
Wh9r4DnwBugSryvBUMyakf/7vz9NGGUmm0VarDh1aDDbolFSyuDv3TaqLaDIZ2ShrRWm6dbGHZvB
awTTEUqr0eo44L8vaRz4JaYpEd23NM+S3EesXtPKG4PUxxTTTQYnhVtUlgkSpxCSIL0VUMut4gcL
HjeP9eD1PfERX9fHX10rEGaI2N+An055kssh9YCWvputZlDOFZo4Hz0A77RazH9efTeVrDx63XG6
/tkP0J8JmNmcOcSpzkiXVCl1Oc2KeHgY+vuianijUG7ewLrd6HxpyioBwE3PSCoEmLLUovSU0mQO
WNx/r1Xon9bNMXCqtCrEhBBFJZqlIMBXTuetRCKXRj4VXcuNFCkcnzTVxY/FG8s++o0WHuDAbhls
vw9SEs/nma4WKG10LGy6K2w6V5ceSTGIOjsxNUjh4vPMuFbdiFDuNBVTAPTDjHnGRQmDImZeYZl7
E3pn9d6JPtWKjqhJ+vsT6hUYutT3Be2Ha8ZTicf0OwoTXUpxiKb9uqmyDFhP8/Y8Ya3MmRZ+z8SG
9XHHhp5zHbKa0WtW63Vn6EOKOMgAapS0wNYSFTsKCRmlUCfq92SpmgUJ1UvUIY/pC4GjZxzeiyiY
A84PxriAbJ7GHLfXVDC2Nzgs//ug+XXoAkAgacM06CjzAVyk2TGXzjTuc3A+exd/fD31Tgebnea8
UXT2Voo8C69E9P+6SJMAR+Sx81KWmXB/mjgV4Phm14XxTHfpPeBlT7M27u9Bk36smOPpd7GaLwFv
so7P8+87KFCWVPTrwOVLwRxqNUKb8M/4Go0dmXBkWo9za8t0BQ6ZCAV2usvlp2zeWUpe6WBOhieb
0bXJAYKDuy/KNnkqJcrrNc9y84YrHzUtPEizBexOuOx3/rv3Jc+Wn+J64fVXm7gI5Hy32eJQSoPK
Hu0gCsyK5amimS1si9RxJrw3ybwP+IBc3wswhSawjvvBXhRkU0lHt6BXWUmqCgwEM1LrOy8jW2jT
SEBxtznjIpqYO/ITqJTS7qN4w4NdQ5lRvuJGKtSkcYatcxhtaG64L/ooQ246y+rGXMvi5aE6OQVV
tpDvHqeoRCK7B8qRyMPmA3Saghp1QMFsVAtJr5AXyfqhIFky+6rHHiMRb4WFL+pxC7FdEiEXyp/3
pGoqTwYh9JFF5QAn1m+fpqfz04DvEmiilK43oFHau5ZY+txuakGpl3Ehdl909MYdNeVceFdQkhGx
C8ptaamzqwRXCk8NGw+1gGWUTqddy2a1zafUICHdBOqCOjee4pU/UyJmUoEFk7YkvhTc0lSKfs8d
RK/RuXlZZ8GOyXEG9uRh95owiL5Gq5HZ2O0Msrl0weblNIN81x5nFK4sBXrVTBY9NIX6UyCbVMdz
klb9JoEwEAKQbOdC5X3EShV3Yv6lvU8TvEIuR80SvI+DUdIpuzCe/R34QZ/KyDsryRUMhf1FzgMz
Ze9OBuTjCUzEx0pQpdZLUimGva+SDuu3A6h9biqY/NmZXpqVnOFAKaqZLrNYSjsVnElBAPyGqOAS
u59Irv2TVkjLl+rT5y/TeZ6a+upKOVmOFW18yR8CUin2eWVmy5lt65mQJQ0lEADjtFVkiYlX/x1J
9KHr5yIWi4GK3yPKuyC3vMkRhwiceVAapn/TIsm6dwmhuE+eD+03z/2mVeiRjEzn3FZKdG+bs2No
QRCdOc2ozLtrfyjksprtiEBxOkvrbp7Oukt2FQ8FnJla1pupzmfyy1d9PvcN1PriDvS8PqyzUKba
UjW7DWVuuQuIB+CWqV6TZ4t30jiMgmE1Hdee44ETGK1seFiSj4xe0qV/JV6lWSJ+Ap/kQIEuWEpY
SxsNs132zxJ/av4A7TKFgOx7AvMUxRa31y/Rn45kecBRJjiM1tw8naJEc7t7/1ej3Q4/nROZyBd0
NkRVX1GeOghoIxBqru49uq6IhgItAgPU2W9FsYs4HVpCa6z8U+5qmbJfCQhtuVrZ+VEvmP8AAFQv
VLjdCfeCLj7PwEZmuJ62bdWfhf+NTv66X6pZoJqHtXTaY7eylo18Yz6JnrCrScrx26/cOcMNAVUU
omr3N4xuccG0gRg5QVfenmKKdLtZD8DlU0YnQW1P89EiEYAP6zxH+mtbVc7agoQcoslvBTaDNCkB
nLgbwQHKxsgnuaI5zu5ieTAKyip/nJL89b6MYLRqHf3HZwfhF59Dz6c60wKAb3Jp4qdR2Zk6oEPp
dpWvIokZ/O69Nf802aYZ6LX7vXFVDNCOyIyxFJFa76815g/dcMd7K069vLe57C/i9KFXGsfiPfRg
mwAiSZ02jLR5eSyCb751ThQ6yNHLMV9mKaUbwzF7mHa6lGNw/0jnQWa4nAtinkBwfTQU+RjfJpme
m2T8YQKcVcSXBel9xc+1ZSyGlS8aq1cScXmv7di6ZJbHEfnhmxyErHYF6BwPq+/0mWa09AMthauH
pvGTRtU/4BXlUY+vTf4a1zhT0DDxqa0/gduWPSGN/n+bTe+X7/QlGH4x1zF5vP459hhYYgeaWBbh
BwLYfc2duatwZe5jpkMMhvrMuZ8RH9SgyiS32WdB6eBBuEEfH12rdVxf4u2JZzjR1uU1JMVCWCR5
K7dKrj+6kj70EjtPrbyM32BkYfF8OIl4Yrq+BAZstKNbdSPhB97e4wxj9jHPqZvVfnkWJx486uln
RozS/ZWqm7Tinm2X0hulqCN4geSzsp29rDRsAISSU/TpwbnRlUMOtSCD4yQqX2HpKyDfnQqtDbIG
FRYVZk+JJYfO2E8abTjQqSd8QJUrH48Tkvqsao8m11SlU5EDNAnZEy3nDkDt4oLFSXtbCxztAXyA
Q46lSUCMMAuWv9FGBK2JFRv7YAEwFT2Fx40H2KtFzEgcksnWV15LTzjTi+mvl5zrflbOvQU6Yimt
ladsLxp9vVImkqA87SFjR0lxwnmsAw/BiKl/A6kl4GfhSvC9lninjQFItMW/uiHiwxi7Tc9WNWXi
k3a1o8dufXdpEvyPUdcftXn/l0tx0KQY3v3gg0Nz5J7d6n5rfXocXjRcZvXgcSTQ8gxZz1h+Qbq/
nLIQKLpvUER1cmu0II96cJYA/gforPd2AyN6pV7KDjC8i+5qfosHrlkj+rtWnmlUi4mLqToKvfCf
Aq9TwK1vXTsg047+W6waXMYRH6tFt+q0yu+fbS3YrNDhu4cTxctUM6kY4Oe3p18/xnrzIT/2T+/x
T0jjsbMxCDKeApROUjlChguObEQCdnnk1rLLzEmMa/l9oyUOICMxFb96vA8WEeCpUrRHmWJ6jbbv
uto2S9pSJO0S5MUF+IutgslMi6lxydAfAOTe30ozNJpDvEc5pDLXX/xjmoFNutqOjsstn1emXtTZ
z8PjB6jagkfUG/mPO56cfkR8VxP7yrS7BPOZz0v97mXfV0+GP5Gdogomof6LRj5VBN8b/5PVrr/V
Cjrw2gKNKYnsX6XsWnU451sYiu0vb1Oe/D8zjkk2yoj8lJSwG1j857RB1ExLxbbVOAC/ANAmK1Qp
6jK68YXmqgqhI9JtXRgRF/6l0p8PX05m2yb88iYeZq3WUBZxx0r3gEHITE2UZb2k2pkfIWbrPX7W
hdK6f8zKVhmGycDbBa20ZnM2pbbUhEMUGOnpi8EVf77rzjy5VzsFSV8BAes/KRJ/vJdf8lNlUqyi
sGOBjZw60R0TWI7k+cBfYa7SQU6dQqZfmFBue3aPJROWrvCHuXGpavHzYGhGU/4T3Qdtb+7fh2BM
SUk0Js9i0iQbvj1dakp7Z1mGN+x4vTt2x59eJalMlJDUen2n4q31hSWbUU6qiGt5aboXiHWwqrUW
2fWtMVItyHu1FV0Nf7DYkxEIdViVb5GTPFi2LxIqX+w26Mb4t622wnlAchwS2aOEFYiojlb1bR+P
Q0roQyXQBLrQhTb30OCFBudyVfB/TORR/VFPLNVFCzfo9JKtiEromnNUHXJ0ZD0kuIciuYp/wXIA
qv9miQXfb1BbVGBqnFhaUd4H4Y9azyx57xBW3HB7s6mplxWmQbsqfpuLC5jIds0McZMU6bB2sgmN
TjJSa+rAvWZYl9/7KF3KP9ME6F5Jg7aZf5qJYBjHVk9q39AlKRcPszmZEJjvgo2f4WnUPJguTFb2
X/jxz5HDDckSvrQS7uZnNIjbShA3GpA60BdnYE/fuqzPakPBy3dfmfoUsxPE4cblRtYjYFFvYb4x
pIsjggRpFAxTmdmXGaHF5macau7jKhTBjeX1SqK/B+5mqWkrB35Jpmb4LzSZBDh1rwE0fXymp2hC
k7uPoohuIlD3xoHMnxUR+y8kb+9RlPTE96IgyaQGAztKYFdoprAqRPQ6QMhFjURPjFtx5QZ4YuBA
yfmhxzu8k9F41DfbvAdP+T/bU8ecusy1fwlpr3m/mWopWWSX/Gcw0Jz1HhulgvViBkHh8EthyJww
kY2YW7kAAn4itsbrHl6mPeDL6+wtdZsUdv52S2O7+4Y1k5SvKIwmNOLhaygzRX8Fj5sgswUEubql
8yYpVidPp/I3GNP3grdMM6ybsrVktFV5HV1q7JoVnRvBhQm8WH0RI66D5+/H2GzVG/mAKzfWF4MF
j2uy6lo1d2WFcfGQg+VvWhk14Iecw96lthaC28zQtIOjP6heXrL2y+QhjrOwaZs/23uIgT65VTsL
jHYvKOzaqj+zC3bj+TYnUNQOL9IfvWORN0avD2mKvxR9sQW5CLeD7uIxyIJl6e0r723UB3Wj8bap
ejg6/6gNbqqo061+jchjXJBcgp5f448iE5J3V3qlX4WrmbHAja9na2M/SkLejqmDmpnRZpbY6T82
fSD1+5/LeDN8DOdq2q7Nt8Y9vFmZQ5pRYPFqSwqZREAKy/DZFyMl36rzcxm7Y7xLabpm/kM5DOe4
BxxlmOk5C/3wbsdmpZTLrxXm8aXAtjG/lM4jaB02izjvh9aA1KO2WhM1gF3BCVcnYDTdBDgTBGzl
SiN2v4TXBNDHwzr5/PLf7xL+xiI5aMeFIAxB85RmqNbQvIItjnr7bs76Ge/toHWvmj99vwAH4WKm
JRXnZzQrQXmPBNsZiZGAzTZiYSoeBrYlWW/WDPPLCfVDwAdfXbbTh7Uzqq+hJcxkGS+ch4gH9Jgl
8Yu2azo3JYO8x83oeHrR6Fp66/r3lLa8/phHNRqxw7+yJSxU80EkTn3XBUntcSH8EbWVmwIS8jD8
cYJBIvTS/VSO3ndTJ1eVqi/b5SFvhKwC4hq4uj63b9o0ZuCy80aDQULwPab1Ou2TX0WVl3EX1TVS
Qh2+R+SwNK4g2yZpFFdjrtuNCzg2Xfdw9IA61ALk9PYxXMnHHWOAr+n2SIXXigc3dYy3u5lGcS7V
xgjdgV9D0pyZ8ok2xfYKrsj3PGWDZjjmmxiKZT2N0qayUU/6Cx/8y2R3Y/gZeXXWAbLYzIHieYgJ
IQHiOIPcyy35RHe4nDVw8A9/yEtLiB3MQN/CIpAC0IH5swShz4G444Ad861rbA/avsTvpnXtWarL
OxIQm2lp/mCzpzTHE4fPCej66Q7YQGVtAKZ+Qeacmmx/np5tlCahoOvcV31mqQjvns1wqts1p8kr
vZKfYLJqk0sU1BaQt3ql6Uc5ZqL10m2x1nio95ZrfRGoKsCkX7ZUBmSI4c780sBwecbBmE/hjDNK
4Kc265qB3dSeK2FhbC8hmqa0foH6iCQz9xkGdZGMsdAdknPH1BHjyMSqu2I1Ts26W9axjjaYmhO2
Bd9LMxkU1DaJ5Y5iUMhTfXkK8L9pKl6gOpyyonXvXb+Nwb1XAaVbzhhrxbXH4lymmUnrLAlBIQhB
04yB++kR9w08yRAC09mlFPkA00kZs6iwZJX8j4zI2R1KPRPyx3/F6J3O4m9wabvWfYXioLZJxzeT
whfIyqOaUaK8ogsvupJxpAf9WW30+TxvH6N2cneY+oNmwC0f25N/qo2PVGzT+mWb2B6rGcdKVIYE
aW/C+22SQEAFj6tgCbGxcVdelU3vLSGp8uv3mCOdIWn4sAo7gTILs5/cRkoFCWZfBTU7vSgW719V
xAcH/VvZzVqUg+5tOxfauBV3FY3qg1Ie1NnMS+iprs9/o1miNCfsNXQhq3Px2R47oV+Qu0aWyu91
XQ6uMifEqMwOOKeyn23ZCQn3ajL4KK0B8bet12iZmzYn69jb73tyXYQwNvTkDWRIgYlkd7KL1BtY
YGTAXpu3WUErgGLS2ojLJlbFWCj6ix9HRi1uJeEG4j9DKs05tVo24m+2dr+KCfNjQzjLRvHHB76I
udGywwNfILHML2CKUlYXhgPAKrZBObK0rNasoCACDwHcepxDDpxFqu0jHecJ2Aqomq38n+m8ODi4
jnwhADCeOJXaEElDrAxpnIgdCA2aAVz0vDiCmy+BPFu1tUAQzkPKTMsgh2mRlxsGLKVIot2fjNiY
dAQ1BkMnurolmjDok8VUiMLzJLCVDBGF1oMXJGoy88jgTUstyndQkvnOz64S+dj/LzmqipX7CoZ9
PUI3wx1YSlM02kxu4ydbIy1TvISWEWlrcwbE6J5A8TOi4USs4LuaXsULUORtT21MrGwT2H3+NJy+
0VXdGYwSSEZSOLRghWEVKYvmzhbNzGP4c5TykTH4SAa13j+oJQJXtWqqQTsu2SmzER/vwgypn1Je
ZW9x/E5bXAG1E7lsH4IQJGJeWPtpPQM6wMReliAJ/LSFhNyd1pBcRYiZQaEPwcqtiFQqpbulwRkd
Y008KOvZL5PurGel7ftgJzRCIMZaH3kAFwC1L9fXT/fEO6mD/+p0onkTWV3Ju9/MIG3m3XcEdaoc
o/nGIwKAhntpSjflxhx0nLi16KlmQ7DN1yVm/6Irs7x1cgaVHvpTnfsp61gnuPJMDFlYMpx+F9CZ
AIGF8ul5FVdrHMHgKQHzcVUTo0XG4oT/AEuoB/FFE+hJHAD87x1kXXFFb1ge+DNkNj9X8PZtBlNT
nEcm6WXbpvVwIEX3wWUKtczkYxmngDXdVy/NZcGW1wOI6tOiSQDrE11/JwGAMv0E950VGeWbra95
QqRenDNSKN/2TZ8d4v+70WKbJsz22ekHxKqlg4KRhkYHz+YEa75hUBRDdxY9/Xtn4EOAGOlHYrg+
50Iv0RdPlhJQRQSoePqqlY0aMmAzdxDY2JUY7eExfj1e7bb7tnWY3X3v4HB8o0bfhlOBH6Q5b8a2
ZXeWm4nDjI8faRirvpaEbCfjOVJeaVr39dmZ70J896S6eZ1hcU5EoTPDmFQchI+ouRfNds2EPliz
VbIF64QN1iQlToGsiqqLRbmvX0+D/8Mjbjq+JcxUnpPN0HoHFVbTUrzVsQDUcdmTulmtAUccWxhT
oC7u3rXS9YiqXrItJNCvLI9OdZSSvz15gM2nEVyaXfIq6Zyv2wY2MsjUN2JjBOblW5YNRd+FiPwl
aZcTlbmsP7OSqBuKa0dqsoQwoFZodxh7QPArX0dl0nqS4P8I1JObHswTR7crnIkuG9n0P6c7Q4ea
tJ7gJZQ6+gS+9jLe6K/EoU69Pvcr3dm+VImVjcm+M5Is5kyJaxWThBHi8b+YLWExhCwbAfSybiJx
IXHQ09EQaoBV7Z9nv/PW4Bgk0XMyfiu+q1YyWsIQ+X6QRYRV4Rg8pBhSgBql1RZDzJaO5yIhM64w
5mux6IoAhBLQ+bK3bT1uaOtml1LsannGF6/hXNXlAPRp8GcNjz0gGi+7a3r4bOIBbBZaqWwup38D
4qwjNuw+mudzf7i0IptmvinLIo/9gn7uaJF+xZSGhEU2rVAjONY9PoxIX/uSNWlbLaYyKPHfhuxB
cVUqEoLFHzRjQXhhOFPvZdAfElETdZ0kkdCfaKmjZqRo2svNfrkjvax8ZSVBGESDn49GRgaCF7ji
OrHccWx2wno3OtEJimkzrV6H8D4OLzECzcFgD17kX2LAnj4vdqlQVh0bOA3PJcm/aPxWGVPXZm3s
c+AxVYFPpSM16IH+kq2UMbJfZcER8ZlPbsonRVFZ5y5B+2sPP/Msxyl0m1vL9ecYJpwHosbwH9mD
/SRGXhIPQFwx3L7rvbUAq/Lakkqp9DjJpfHlyP1IwFuZLg0AYrmxIfxwwV2BWWyYYGPX0E4DbSZh
ZSml6vHGsNwBbaYoifRh02FvwjhaH3B2ePdXFT/qTZAtt2IdxSlsOEZpljJtTr+jR34z6cg8gIYd
46/T1xn9BXWf4XCjzYUIgVkZTsXbR36UNg9pB02FrO+jq01VWl45aTXZhGMpwd6kz8E6c3rBRfrh
xyxsAQVT1C8vpGqvlmVeXdb6cCfuYllT0kPLUOv552kQNQ/A4dB0S+6x96mP4AxJxM13XTRgvFfD
hGJhiFRWXzof+MyX721yb1Jrf8TaCzLJzze7Kj0HmN5eOkpLxyFURxeCekZq35wTQCSJQ4q3fcEW
9nObb7hiYuFWm7vqb2aLk5SEeNEPY33S8RI4lKbqOLfFyMjSnJCluvmjk86DROidYkqLYjQ84sxW
9IN97W1vgSoobzrvKQaF2Qf3c93YnWwA6MwvCbRd37BVInL8X/LZKKhdxBmk4dZXO91ZufBsjLe9
IkCii3FApiKJ4sveC3CeHin9zilUzABC5i3lYfNXggBB9oTtXNZQ5zJeanzVbbQRnnR0IZ2mXs7R
XXQRnOlJvaj4rstvFhRSRSf1ONg1Q+0W+MCgmjX6k3bHPxDWwRZjcwcoNqJRGSxebuFz7xUhH6j3
Tt7lXcr0EsAPofpBj9GH7qWKxbvsfGpmpp11BWBAMD0P5nDXge0ZiXzAGGLhr6KmLwH+EuxF+K8i
gYe0bFqOh4F90X0MiW9GLZP6bPxc6V5cQWkSC6HIEcIR8QMxBpYzfziblln5DkXZLBvEc10WmXG5
Zzc2pgnguJvACZatVgjdTaqhsrXhBZEvnLr8l3OWOg6MVlK1/YUlFfUE72lOQrFBf7U3nbj6yn9z
KaxtcylquzItAotRHzB5gx+lYIT/X+kaF05kYKHu/n4i4+asFHOdlYglUxfKwrorvULKYxS72Yx+
vj5eOkyjE41Va5iLfUVRKGPEKzVNxO0j98fJLfoUqx5P52do7CTrTphc5d8DnNovJGkdurgMpsWI
x/waeSlsFFI1nhzzjDG2PVn/HbBUh0HyafcTPWfJaVV45atyqP7pvLXV15BigfabBdGNPDjmJzGe
aBTno20+dKkMHiIQZk9W/Q5gWBpyhTRiDZ/BuXSD/NGUSQQgDNp2Zv8lj4+fF3H4/V0l6V3cOGp+
qlMMhAHrARnnXMVTADrPBuYS/1ETb9k6ifby8XOX3dE3+X2qX8IXBnm/bDKgEq4TQhJI7NVIIX5u
WmYMxvSTOOBL0QVSOsmIYbIC10dC6PEJdlOlWDWx4C9YCzfERQUOCZqKsjdQ+/ie1WXENGOyeKFq
+4l4UbJGlE8CGC+GNsrMwuWcO/zAaSYcvJqMEivzj1sWEEJKoBu589voF43dkaUaqZXia2tPQMv0
lBePrndu353tUUTAd8UXUk8kTp/aNkbYRp238kPidVFgP7CrEssr8pD+84YNdRrMkLocvmtqVhwB
qXKtXC+o1JjChTjE3KXKjTTk337b86fbJ5jtAWWa61pcmkOBEVg0Ke2I/YNgLorJJ4qjdU4Z2M3Q
U+duY4DKp5z0OQQiAXZPSG0PDIvu9b9Z3W9jZ2Y1SosSSVs6N4KdALvPd1GAo5qn/dzGqVXL3psc
zsCCTmXv46nziR8y0nQ/v9Rx2KEiriHFkOWGTcBkmzvPb0iJO4iL9oV+XIHr3xT0cvzMh8gX5jN8
Ggh5GiIQxt2rBj2B5clA6lnBxOMspFQKWYehpYN2s161Zy6NbvMxwxx+B3WpB/buSNICTQfOqYYh
MY7M7jsi+Vdl1oJajSpWvCehqmTcfUcLSeXEWRzJK7z2RiWzbmwY7FlT0rFu/atn0shLkOC2IZUB
RxE3a8lnnBnfzcQDxlAIKhYCA3XYBaLB1uXBGL4xEf6joNdy5JhHxndzN6kFtq+aQTDC9A4Z2A2A
hdxEvcny7cOse9e/oaQdFeirrBFKcXlSOWlAK7fwmsOPjqs+RScPjQooC6Nl+pVWEXhAK/qCbMJr
8WuOXgzbS1gfYuAj9hfl5RA44a4KinQBowTv6D6f3FGAMstJKVC0luZTJvtH5s9SGViqOL5zBzXX
TlWGj4PV1Xoqv6PGie+7JeSCCt4TKFUrMSagyT92MKdf6vF737S4FqqbM9uSB5+GPBfRKEpiYGAL
rwlV0GvWXwsnXiQBTkCm7A1S19Wkl5H1cVXF62pR1x2Tuhgk8zqS67e7cqYy6INH8x2glszo0ryl
UmWnmaqaVTek0jW6TUDbkAPQozo50p2D4DASnHkVpMJPOf1awzrbbLJ2nGXJwry8weo76oG0vJ6A
7cb2Ym29MRtmBCtVwppwuWOJaGE6nvxQHPyvra3+YeGapk7jigYrbXKPZyocaaBzG53aeVFiTV9J
+YW/nNLAZlb12cogiYQBD618IvYXUbdSFaAMES5zonnifzrPTp5kGFcjS/7Ck58I5+p8Z9iGB/h5
V8wbD9g/4ZmJyWawB83ea5M1b2qMsU74JloaMEmVKMWwXBNX4/cQOHUp13fCTW9D3njckJXnKQte
lus98/zgBZfR2CV3BI/20atc8J5PwFW9rJ3uht36F0CZSnV+VQbQ+AvnXdgDCTAgcRZRUcUeQfP7
HDc68zaReLkFikQtCx0coGxtgmwhMPeFb+vHGreEVdEz1TtmxszEfSAfIl2B0JBxcwxpwjHuK4Nx
DNLoCZAXBu95HcGE7swhwjjsdzjbhV46jxvzrDIcKa8xivMMyyODs9gn3J76mwquaUi6hyREQDnX
VyW9HtCCPPvbWvHjx5sn7PRmfpOm1lYNP/mN+mCAxmUooAmhQ3zlxuYqGYnpclZLJ9gQXHNQnemZ
0OZEpE3LnTFxFT2On4FBQqUweToeXCc/r5tqjcmzkqhTTcuhBRm2nGQj7PqkW3pce5KjoYl793x5
LxbsdGTHrJJ/P/mysoFUHacJxCqkpYr63kGtm9AWAG+HkGjpmWfIeQ2/kya4UCbAcjO2zRHPNWzF
3ArPreTHjZvOgE5cosl+5KOGpGXkyt7mErHV72V/q5IFEy2vkPGU19U6lilevQC4gfOFjJHJHHLm
CLa2iTRhKrCc9F/yqxlO2ZqwPuJDweEFCWvwofnDpW2IeJ+pQ+OuAobKXawJDdAKe0EefuH1REu3
TOz4Q9cKP+mLl4XLdYZKYkvUUjZKUwX1F1m+9H39aMHFTx3k6KNMY4SINxI6sDJJF8jhby2RIimJ
TYExrCMjKRY0GrpjznzceLv32jQhVRT7kpkW1LsFThZaDkXHcFX3ROmber8lZK3WPqtwbQeaMgSq
CveMHVo13c1lq6GyD8f1nblx37DNW0eYBHCyUBFK5ZR7Lo85CeXH/yGZ84PC/kW+k0z5/7k6RPSQ
1PG3L0pcex5J4YCFDnOwPnjc5RRk6NIYVN6rt1S/lyMqUCdZysFV4RMC+pAjFC4t09RalnmYATRJ
Ei9MLhHrasNWOKbFy8jYZrSVe9ayOFcNVGpZ6ZxLWfnPIZ9kbUHaU4AVKhNj3/2ZfeDa5E94eub/
zrD/B3h0p2jkfGnZ1mhkgp5TgEce82Yc+yZ0F4ZIzrVfHvEOcIpiUfqtJ/zdnaBMUCjmFJuYU/Fi
uuUK531RQHfMjHvz+yEYcu4uOSqq5AopPW814Ab1FQuNy+zOfZhcGGKsxA0afN3Ey2Hds9zG9jrU
jq3rgCXP7aYssEFPUVNw0N3/H6X7rf72My0kP4GJVC5XfeLsoohgnAGH26ADxzX/iCD1VRMOni2n
XKxGzmtqgiNspF2RMSGyblR6OWQQgs6QFTVYN4jT9j3hqvUiCsSmcnxWIUHRKksRLXlWhBTu5EG9
kbS9HJ7t4LxQi1xg50Wlp1Muj2KbeOggDgopJ/j0XSmJIa7pA4NLIrZkuLlopRFrKh1HDK3a9sK6
fUYoncfqA5jrxEUcLl98kdjOl12EV1suHsUVB1EYYoQkpgRAq6FoOjSZzMUNXckc3hNY5x2kK+pL
P5JdT2pSd9/8GAlEV6Zn5FKbyN9dJSOLYBLmbsKr8m3DR+Xse5rQzCV2PJTeSFZp1DHtAbQlVsHQ
Yn/M6MZXhrogW+pviT4OUXCnXtl9p3RZ1wPu3pF2+WrPqc3Y21W/Gx4bO0HBp055GwiC4UWzeqy6
6nT+cE6DEyLpRCVcay6W1TVmunYc9P8ZNB3GDZSLROheDWh5UkwS1J7iEkIxMLaIOmyPFu3tjbNr
0RSTAO59fEY6oQfdPdK423aCpEHZN0M1wuanxo7hH0KZ0e2NNWAYN5xa2Q+D0OlN3GBf2/UHzE4P
oJRdOHOE0lOtF/rPmsUFjxD9k01vim+noc3sb+umj9u7RHOx85P31b6cNP3wdz69au3grnbKobN+
jBuKOxYNqD25rVcDmUOQbvJjWwjmd5+8EOXe5JTITsfiy3LTsRumPtXnPKmFEWbRLcVy+BUipu0h
vyx+nlfTAO36MlIig6KJXnL5k+k9sdZr5rowrv44SopGvHQQF3ZDonApxluV0Cqz9n41/N3fC6yz
VAlj2OyoI3Qo76cSkZN5g0byldaXY+dri61GCvDszp9cZAKrorTEnEILHY5p7eXh3lAcFccp2Jq0
FYWPLWbOyviPbMnpbb9RHNQ66yANcqVMqym2KI6PB5I7vEnhNBrsy/wD3dThxM5R69TAHr4l73eW
gt3G9y1PjpyQvF02JcE8DqFeow4RNYUtOBS1YD2Kr2EKVXoBIl3IgCC7Hl98HZR4Df4xDFF+Srxx
UNAo8yKZ4ZlE9s20shOEnUfsnyDJVrvUCFRQSKNh4opCaU7LnCMJ1j/JIcpS3dSgWFtFx7UhGX1S
nHU5j/Uuge54n8AmFlzqiEBXDCRn29cVRtjOQjisJZ9TAZjLZNaOSaN5TToCoQ0FruZoG4356Zn2
/1Jovis9kTIscbsNM08g4hA6wC7xxbvzX7aQL1Sei+g3OdBwsn/Ex76EQMaNzXMjKCmePEMsF/eh
YdRrH4cMAjtNUiE73UbbOvMyvUtkg2O2DfL0Y6CNPLGz+OinYYygqGU/AzX4D/r8IHQJcCnoiNeZ
iMk2yDanX/HHok57PoLnwrHrpQ04zqA75pDqQRm2DOh/murbfzi7ELiQpCuk5ZmTSIkfLVjsM+Ag
JfMKNNsq7qkFoEg42shpVuMkM+s/Bspnw27/YpvX1OKjVCtysW91WkjNi54t7dzdJLxyXxKEyJU+
TLI5x3CBtu3+dcFhysd6PM9Hjpy+FmqIq4rCzQnbrtepZBUTL7YpnrhkbxZ3/n6JUgj3t5g6L5Cy
JWoWhmXZt0MLxiI1fBGvnTGHnSNTVqNvElC39jeeXe6wO4FM5cYKo0B2+V4CsjIRU2ul9zG8riXu
BgzUaF0sTp087QLkJ4NwP9SmPt2DkchdvqB/GK8Av99S8B14bfjYr+34bkQntN0wCs5iJttX/GLl
dCebKzyjJAEw0BLSuG/QNqk59bhqinehQRZ8p3cMKavSZypDuvWitbQ8KPB4ww7eO4ozyLPz117d
MsxU5fvQiH9w/ul1aEbZUbqkIvIA7RuhQLIzBOYEo+qChzGrPSMqCG9nnz+PennYo7SBVGONPzxZ
jh6NaIG09yBXG3AiwyDIhzYpeGuDpbX+F2TMRq2jNaD9J5PBDtk8r5BgwO8Dm9Hi64wHoUPSkGws
t03xGVYbQhf2tobBS51/ezv3T4B4LgG76D54/UXZY9WnJhVZBZwprh3K/cjR/M+UZt8mwqDdijsN
L8g0daXs2qwYibHIw81UflH11YSLt7faG2Yw58XzCGS0+yDxsA6FQ4ag0Q70sYJ4L2GBsmlStN65
IfDtGIHuuO/FjbVN8qhDNUfbxjl43Qab6+2H7w53Qi2gg85oDFH+Ouwb9o5SBY9DPNAAZhEKzDOc
rOz3bWEplwh2RyUaJzpJA/XUlMrwny0QeQ128g/BRSIYxahmVvXaMta/4bxyeAf4ZbcYRp8MaYUO
//RSOSul0oeQ7XIQaf+q3c6LdDZtETSsByVCbyo7w4cQZUb1LCgT+n1C+DpOdz5X2Sk6uXy8GesF
nqhdxQbKqHBBb1c2xIKiebEfO+zgEXQHmsMfxy7O9kUO/1nHxDkLIA2G6S6AbsmoU5c94mZ0P45I
nCJurndHDpRPvaxAO2EKHGPHopy+pmGD9csOKHQcONplskJgd0kQSV20BKPPgTgrXaADq2nw64Xz
ycQGFRsH6M5iqJFUCWh38PV5gTKF8CgdZ7v8FSrj8clErRX2SnIraOgr3mIif3wdmbE8eC+95Zc5
B6bdPycrRULQGIsKyyJruJoK+bjFIDV0peRt3PvpcMQK2FKQ3ujTB4Th/A4y8w0Q/QGNzRkuzwD0
9P5cvyo52NBW+t1x5kqswZXt9Q0oDwFl6mOhwfmHSa05dO2N/HfR8zfVi4/PSTo2kJh/LCypAeUI
gylAjGGXPqusN67LzXxkimZmnnkdMFforiyuyESdHfykfooJyd3b3Chtu9vr6o7AMceps5hWVLiU
vAInCwWEYPmuOVo4PgUuizS991kRlxvfr4R3KUTmiVpaGuULcqzMUJwWBb6BBa5z526PxRiF8pGo
NwzW8tiKYTQeYzsHpJIe2ptnTaE9ISAa6sASoBsTil8QHkp/KCFuMJc8SpJH/zosH2+axjghQB0q
XRFK6hlFmBE5CRE0Vs5JPL9NVhS46O4a/Ei94ZD9B7ZHkSyI0UKS4sXjKObOr4PJ1KklQ85mCN8A
dYTcaGkZWQOPcIvb5DTCUBQwG5g99GUTZ3y/IUaPOb3BfEy7PKaejs2HK1fdSQeMzvrRibOqytvz
kBizRpHNqbn0XI0/KZO5zHaXXdlRhk9+I/INaRy1Y5a3QuMHDt4NLAS+PN6swtibQaBTzzPh9NFB
KsL0JwkvQ9hrvQiS/FNZVVpS/A6ZKvp7hGY2TD/ZWZoQgk3NlbOdykdPFv3byf2KreL/cPhaPr8x
b1rw8EBcne15aQDBwHWK+We7YkaR1ulxwQbfyD1F/yHqvCzDB8GtPPZSbz31Sjwt/miuF8NzaJ2X
fboRkJcWLXjHUpZWRXaBCYvwfNFednEYh0l8B/6cCMF+gPkx93/BURyzi9jygE+PNakrmNMBkSmL
Wo3SUlNt3QgeYyvED58urajMrxrtdCEIGS832kb+GhzbakRLtTreSxooNwQRQK4lp9oxBsyxZccs
wO+ms8SEDfpPM6JpEOcvuvsgZUebSqZAVHdACATPjD74FO39jm5c7k0/jKiLUreAN2Pt7Vpi15CJ
0atEFWEXDygDCIqAuq2JNM+lmqc=
`pragma protect end_protected
