// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WkAVCaWAiQAmgO/BS0XpTsbMiMKV0+RpFi9y6ZMCXc5MfSWaPlEV90jhX3eUYlUR
0qeqdeRlldu6mAdBhyyEIqlfD9WdwYrobRPPNf3NPvwvReYQsXKfdFeYuvxDHYGY
xN9yCbvhTE8tE6GLNWHIANlbFLHiTT3OFfeXnGRf8DU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4352)
Q22rTxAdsL4+tR78QGApd39QwgvbrqEy7I3MCVSCs588/pKd9n5Jde+bG0jJKNGT
U+JZrLV8e0io/XcIYJWH7uLmL+rc/8a1mjlDCSzDD3ncFFyp9m6rG5r+tJRvwSXz
VTtHbf+uEB1MuCzqve7+rMzeW0LtoElrrmXjIQm+mMgjhSNTs0CsVBm2qKtrfDEc
abZ3//nDWHzFXfvz8i4rKCS/iC/lChU/h6SRgZm7Ag41agKhXVrs1dWcFqExI6Mg
z6FQbOI9sjNSw2kgjho/XLzxEaTr5vdCJ22UkLBEVSBWAnwcDuGRYIQyJETBPy8R
2nFKh3EyzeFTLEeLzTBcQSjfgH59aqnuV3L6K2XDWjKA47l4afqGiUbn1/qM75sB
IqwMjZFfOVcpYrxbOhIBG2QUA8GDyJB4yVuG7a+lS/NDJCdF9lazs10l5S7ZLqcn
1AT7ilKR6qd27x2zEtFpWiLykRBca6pF61m9IC9I6aH3ANOlq9mXegku+DunFBpk
7s2u2tUFR1UIH1iT5IxSCPmXccItB2G+BGgj2nUa45CXvUDIASLkBL6Lv5WPGxDl
Ict/LKlPo5oWEbdFCVvU9xhtWHCDxLiR34e2cANVFObEqs4O/luvDtq0fK3v88Us
N08ayNDfMxAbFu0+A9vH6+CbscSbmFJ7CnEDjU3KroyhBpedArrykBnPadPufqXj
EdDxYlblNwvDMrBmfWD/hUh2yWokos1wlBo5t/r+PP3Ktjg+qlf0RRWoLIxq/5pc
ibU1K2noigUNDBMYXXIqqhMR9ZpNxa8zpooFBkm9cqHUdzknJh3jNJyBgFgCUZCz
6SOLSwK5Uo/19F1Xrek8EBfb6jfwPNduoJxC84Z4dpW0DxSluAXYVE56nbhfoL6U
Cu2Er70v+r6rQE9gpGDOy+rUkBq3gQquwOoKLEleCmPdZTn0hWZh1YXl4Mnwxiws
ZSREqqXlQfINLHd4DaK7slBNodDc1rYX/SwDxsvwKqL/ZtLYOHYE4gnwVhkX5lJs
u5Rd90OCEQ2sYr1DTchVehCjw+HY26QpoJ8G7LXL3NlS7tG4jOVhjewZ9NIoD88r
cI+1p54AvcBR58t41swKltUL2B49F6C/J0ixyiCl6iXxPCbJbtaFe98r27x8SJSC
SN5Qac55PUGmj0MPh4XKh1l5i+Kw35JJzQx762p/4ofEQbJFDXlG0fyS9jZlG6a0
X9SRJqHq6CrX65cShuEIDwJP5gLMBM9ZjXPX3UNLCxA/MTQMKKHVlA2aBZ/AnJER
JzdQ9IywJY7DueZ25WvzYPRqL3CwewEeopMZE7NlQk9CgPMUkMeG/oJqeGFQYgs/
/R1X9I+8oYYGO1HGRwnkeqSAv7KKJ6OEzQvAgbhxxRe3vEH0CxwFhn0y7pSyovt3
KYm9/H9/RDmlZVV3CiYSPs9/kM4KoRvWxVkQtnNyOnOyz6+PczAGqmS/vejG0+ZV
0KRXibE7hxIE+9XZj8HAN5b8LYb5FeXoqXEUJ2BTJWindZPhhgXAhVp+y1Af4SJj
KJpD/9+yEu7natv2D1bs33XqS9vUALbW9RHZ8NZdjr0VFXpt1mSGB0q3GAgia756
W4eOuJxDm+24TANNxE+5sfJeeeozJNHbqDV2CXmbuewr0wfHK8W2A2dbtNve/B3G
X5m4NUyeOPaWTO7ln1z10ewCsoCeJsKkWaX3y3khPfHy85RmUgzruSHOZEqKjEPj
CsfBh9fkNwnHs4hZOtgCPMln8n4WTl12u+D00aKSNUa3DZW+EUJS8oz4scfWxb3a
Q+tukNK6jXjvBIy0+aqHue2mLfG356iLizcfpZFyVhlspHmvDMd+WSEVzgVi47Sn
oZnnb6aEH/HiSzfBYWo/TpUQWEiDahjNMVXGvw+uW0N1fJy4sIMldm74kLwCIYf0
Q4sSs6B8QsKsmkGNpYokPp/3HX2DcrsDDbrYIkjlWXXwgkb5BHetwBuN8sOt+cHn
ndhDjt51DiB8MaNMGmGuC+rYUi31HlikE07y5E8zVam9a+C0ueraLMfgoxsivUJa
VInt6lxAVE7qA5j0GBWnz2AwkVu4/MTqpn201W7Qgb/uL2WSz/gXSg25wh5FXg6M
Iea6U8aE/c+nAk6sJwuD7adG+eBrhmjzvkG4/v5F0Y1FJ1ebGcc5kAMKQVQyuJRM
+v4ohdGVG85AuJ/f/uzS8YZMjVXAoEMcmI4qg2nKUKY8iovrWyeZt/enDggYy+jf
vQDKlOhHYH/DZPWfuGhXNb5E1BVKiLakxyPBGfj/8SmopZizWAfpcqmp9GC+72R6
Q9KXuO6xG0s8VCRwHPT5vynObl9i6dP0mYXB7PZkHarBo8qnF2fBUzeWskzUk4vu
35C0x2gUCSRxDGnkt/rb5K0G8oYAtFD7YF4Dzqf2BaXEdhxUCiXXo0QmiGHljYp7
64yseDoT4D+ZeFmrZF2QsmErf8i/E1JmPhKK/K1jbnRbjs0r5Vj0VIbW1O97ENLv
BAU7RO4xorAEs7tCwNSbqhvAom/cMVcrCDcqxDS5xb9kmoJoWR0Fces4JeS+fzdP
1vci4wkfQavLJh0lI9RISyx+CN8LcW6bthFb2LlwNH3vC2QILt4xQMjgTmHJC0R0
9unq1kap9D7isZmP4O6lMbb/+XN0b2+BLaF/gcr2FDYZUrwvxofFdUwhDKqtIPn5
fQYSM+Gt47+z6wgQFvifwrR6fRm47js2k+0gg8+h/nk1eS5NgppGyv054VZ3S78d
GKgFnLhQ6Jq96YhCEbTmPMhn63ER6X/qGWso/nSCPQoT88p8I+bWt0GdY+A85UUS
LxqFm+zKFmo4HE1EQO1HMvemHXWz8fpn/OEdPoAgO5WDXPLMpwx94vuRIHOw8h/r
Yuzj/KzYKx1ZG09a+YVuYvIdteTKi8Bc0WBKljtwEZv7wuPvuR8OjLXLzIQc/r35
IHsXRZC27cGbWNzlVG1S/10KUstsIonG6g8FxHoj6DvRNh0kcvfABtO96RlHq55i
ZOB19V+lD0+bLQ5OvDfpmtIMW1DlyuupqP+kisfqf14ua/WE94ISAPmkMgz8/48p
XHCTVhOJfkGoL8quEuIu/Zbn/cO7yW7rtUAwAknKX/07uiFxYptN0DT+rjHyhf+X
4p4QlbUS7ttUXnCjuhbAap62ulkyfVbu61teQsx+rBCPDTO5dnAnB5Ys3uUkBDXQ
V9aPX74nwTQqAml6MAV9/dKaKW3Wbp5yPMJL01CkSRg2FuOR+f0hOsu78OqyHRUg
6RjLXYhcQLTppUnnP51oj45jsMG/Yll3i3zGcJUWdAW4dP/VcMzyxILefFgs6i9B
DbMedjqpSYG4Dl/VadxTGvT8xWu8qXGukL1rXJczn66DEth3dy+ji6eT98ngEu/k
LrHwLkOJxp6uSJS7LuZX5hVrhlky/S7iPqQYnN1Q05RhHdMIhT8BYY1ByJakq+lf
SBfBixHI35b59HtRWLiXg9qIZko/eZ7fikWEjRV+vv94Em17+zZGBdNwkzDgEt5c
bQq+iVOzhP53HN8jYm4Qyckwv5dWGyV0Xvsun15H9RFG8637UstyQ8MCSeNzQfWq
DcHR0LEN2IZgNbsukOyuEokgevb4fycBWTEGVJwx72brfmGik7zOLb7xG/rUrHJE
qi4zCqZQdMK6vGVGzvUEhmVCsGO3lPYLyc+saYbC5H78CNWW/UAgTe/eM6vRnfOp
WJOBU1Bg3e6H68d8wz4H9+iJkYZY1LMJQgsWnvc+HRc3CIc6p+SvlJPMj3/kgi9j
nA9bUyjPxypm9QvvpDYr+9syISquiZiUy7Cz/cs1LwiQN8yn0+BDRm25/AFhDB/F
Bmsz/cYPBCUNnqllej+u9t/IL9K9lDCIh5rETR6P9OXBsZjtjp+UImC08PbzvDes
31U5+iLAfce/DlG57wWvDayHzYlXAVz++fBDadzmsj0KPxT8E6ZUN2B77vEnhZCy
D12QlRb4NqrW/MfjffbC4zw0yDcWSL2SH2uhVf+SzBtmRJCt1M79O2tlR5kPKS9S
MA+qTSoLlJMmWapOaRPNRKAO+MOuWoP98lpeq5HYb4IMdRAttuv8iNjID9/ooday
I46FZuFtdLAciCmlleTH87OD/VmKJ5wnqZp0mZD6pdJWGbkcewOk/TT97wmaQsQn
cTvWk94kNd+vGO6mb0aQqY3ztXRvgqbjhPU8/2OTNe2vZubwf7PVdbqImyLQut/B
boWtFuLHKgdqRtyIDThoxPwa7g7gNpEqTtrro2M0+L7fNDB/0h1xIfVWmCLNOjC2
GCrARjXNpYTBm1n9y0rl3z6S8cydcE+QvWAudczefMlQWfoAyrfLhNMGR6OBD5sO
1DXTWwVQ9FH3SWyulXd81zMIjBzCVHYto+bsfpyUv63qvXCBfxeSBIGYV4cNvCcS
PcAwRQr2EM0sfNCLAOxPgqbDkIZZ5DcvvVIz6mG6UwRqynwCAdl8u8QQuKh9ZxoB
XWssWF4hpx7GiSfxU6sXBFJXrJfBIiPaq1Cw2lbnKWnHwvf4xRp7Is6Tcdje1kSG
LExGYhOZf1ZVup+9fXRx1z8jzmx25nCH3ZZ6J1cC5TCpXExy9mj/gL8NJmQPNNW9
df6xEtjyY+9VNVY0O78hRtnlEm3059lvHGK+mX/rZLk43XMiHS6AC7kUC6KliG7V
HIayQoWHR4mOlepGVOAqXq2m1yM+opIhQi3FzN4WzgxrkSsBJuhnp+9UxZpwwxND
XkIPBTOot/lXwn75aYYywgqQ38yEY/zyQlvoiXgokW9wphVr0ZLCkOOAvvktQ3pk
ERINqrtXC0709iI+2K2nZQPzRWGrA30zjjF3JxJ0iR0X65dX9UlV7XibfhmIuqIT
zD2qjtYK3cSulyiQ8aDr6it+13M1DvLTnKJcxTB5N542pXjiRzidAa6meopZtTA3
pmp6y+xqcdqqFYDtky88kLnWwgMgjxMTq2GlmNz+iNdgKmyzpmZo3JsmNuUc0RvX
n9b+4xR79rKnY08C9gxx0JgSjJk7qc0kLK39gPeimGU82kzLTtMnc5UiTItUEuNm
Dz6jPbo7xCqbQ00IgCaLjW9aFzjSdoEn7/cH6U/aTFve5tsZelI8MGk2LTvdaKvR
vW3RtLRXN9xrInRVO337jYzwp3KYC12/L5k8nl/UQDpUkNsxZdFRK4HmcqMTVkus
l5PFJC8FBF5e7BRFsFfGZubhKLLeGnyOrbInBb6pgfGPbhD1z78Terre6Mz6n+Xf
N+Z/WDdBodMeRWagwnVVPf0wWXWehcvUE0UhXWnlx61oP9+U0kgOlhIAgyNdWDWT
PND7vxWHrj2AS2Oe3Jr5iZhgeNwEPmtQsBEsxWoTgrJmljOkMjnuBr0uFe+2ntP4
iPeUVJH+YyaJ2peQjlLQ/F2v34i+x/svyeMQiS+VMIo7C1Sv9Z+Hoeg7yNt1hF69
gHZUfuY8Tqyh3hukwJeTpcKvK8XCoPVPViIG/XKaHVreQNDCqIhefiZWKnHQk3nX
LUkFQS1LcIHilm8G/vG1sN3CsfFUcG2n+j6mifght+bkhnE6dBN4DLCSgXfIFhUL
OEnLiPI/Ttm+vy0wU00oKdJ1O+I8JUZ01wDNpxjTZWVCUbvkKlEkA20Ul4ktFKUk
eBBpkCy8BeYYj5LCdvvAltGTHsG176g6+ZNixZSvzKI7wx2CkxzjXp02EtFwb3lT
krl2oEZcqdw22LN+DbPIMkFGq02+J7KmnqbvpEdIUVLkX4BaT2gdXBVxZjAKYe3o
cvCMaT0EnVBdooY8RKggBmDxIkyAdkufGSIF9hA9VPE=
`pragma protect end_protected
