// megafunction wizard: %ALTGX%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: alt4gxb 

// ============================================================
// File Name: rc_s4gxb_tx_2pll.v
// Megafunction Name(s):
// 			alt4gxb
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 11.0 Build 157 04/27/2011 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module rc_s4gxb_tx_2pll (
	cal_blk_clk,
	gxb_powerdown,
	pll_inclk_rx_cruclk,
	reconfig_clk,
	reconfig_togxb,
	tx_datain,
	tx_digitalreset,
	pll_locked,
	pll_locked_alt,
	reconfig_fromgxb,
	tx_clkout,
	tx_dataout);

	input	  cal_blk_clk;
	input	[0:0]  gxb_powerdown;
	input	[1:0]  pll_inclk_rx_cruclk;
	input	  reconfig_clk;
	input	[3:0]  reconfig_togxb;
	input	[19:0]  tx_datain;
	input	[0:0]  tx_digitalreset;
	output	[0:0]  pll_locked;
	output	[0:0]  pll_locked_alt;
	output	[16:0]  reconfig_fromgxb;
	output	[0:0]  tx_clkout;
	output	[0:0]  tx_dataout;

	parameter		starting_channel_number = 8;

		//added parameter
	//for MAIN PLL - 148.5MHz
	parameter		tx_pll_inclk0_period = 6734;
	parameter		tx_data_rate = 1485;
	parameter		effective_data_rate = "1485 Mbps";
	parameter		input_clock_frequency = "148.50MHz";
	
	//for second PLL - 148.35MHz
	parameter		tx_pll_inclk1_period = 6741;
	parameter		reconfig_data_rate = 1483;
	parameter		reconfig_effective_data_rate = "1483.5 Mbps";
	parameter		reconfig_input_clock_frequency = "148.35MHz";

	wire [0:0] sub_wire0;
	wire [0:0] sub_wire1;
	wire [16:0] sub_wire2;
	wire [0:0] sub_wire3;
	wire [0:0] sub_wire4;
	wire [0:0] pll_locked = sub_wire0[0:0];
	wire [0:0] pll_locked_alt = sub_wire1[0:0];
	wire [16:0] reconfig_fromgxb = sub_wire2[16:0];
	wire [0:0] tx_clkout = sub_wire3[0:0];
	wire [0:0] tx_dataout = sub_wire4[0:0];

	alt4gxb	alt4gxb_component (
				.pll_inclk_rx_cruclk (pll_inclk_rx_cruclk),
				.reconfig_togxb (reconfig_togxb),
				.tx_datain (tx_datain),
				.tx_digitalreset (tx_digitalreset),
				.cal_blk_clk (cal_blk_clk),
				.gxb_powerdown (gxb_powerdown),
				.reconfig_clk (reconfig_clk),
				.pll_locked (sub_wire0),
				.pll_locked_alt (sub_wire1),
				.reconfig_fromgxb (sub_wire2),
				.tx_clkout (sub_wire3),
				.tx_dataout (sub_wire4)
				// synopsys translate_off
				,
				.aeq_fromgxb (),
				.aeq_togxb (),
				.cal_blk_calibrationstatus (),
				.cal_blk_powerdown (),
				.cmu_rateswitchin (),
				.coreclkout (),
				.fixedclk (),
				.fixedclk_fast (),
				.hip_tx_clkout (),
				.pcie_sw (),
				.pipe8b10binvpolarity (),
				.pipedatavalid (),
				.pipeelecidle (),
				.pipephydonestatus (),
				.pipestatus (),
				.pll1_locked (),
				.pll1_powerdown (),
				.pll2_locked (),
				.pll2_powerdown (),
				.pll3_locked (),
				.pll3_powerdown (),
				.pll_inclk (),
				.pll_inclk_slave (),
				.pll_powerdown (),
				.pll_powerdown_alt (),
				.powerdn (),
				.rateswitch (),
				.rateswitchbaseclock (),
				.reconfig_fromgxb_oe (),
				.rx_a1a2size (),
				.rx_a1a2sizeout (),
				.rx_a1detect (),
				.rx_a2detect (),
				.rx_analogreset (),
				.rx_bistdone (),
				.rx_bisterr (),
				.rx_bitslip (),
				.rx_bitslipboundaryselectout (),
				.rx_byteorderalignstatus (),
				.rx_channelaligned (),
				.rx_clkout (),
				.rx_coreclk (),
				.rx_cruclk (),
				.rx_ctrldetect (),
				.rx_datain (),
				.rx_dataout (),
				.rx_dataoutfull (),
				.rx_digitalreset (),
				.rx_disperr (),
				.rx_elecidleinfersel (),
				.rx_enabyteord (),
				.rx_enapatternalign (),
				.rx_errdetect (),
				.rx_freqlocked (),
				.rx_invpolarity (),
				.rx_k1detect (),
				.rx_k2detect (),
				.rx_locktodata (),
				.rx_locktorefclk (),
				.rx_patterndetect (),
				.rx_phase_comp_fifo_error (),
				.rx_phfifooverflow (),
				.rx_phfifordenable (),
				.rx_phfiforeset (),
				.rx_phfifounderflow (),
				.rx_phfifowrdisable (),
				.rx_pipebufferstat (),
				.rx_pll_locked (),
				.rx_powerdown (),
				.rx_prbscidenable (),
				.rx_recovclkout (),
				.rx_revbitorderwa (),
				.rx_revbyteorderwa (),
				.rx_revseriallpbkout (),
				.rx_rlv (),
				.rx_rmfifoalmostempty (),
				.rx_rmfifoalmostfull (),
				.rx_rmfifodatadeleted (),
				.rx_rmfifodatainserted (),
				.rx_rmfifoempty (),
				.rx_rmfifofull (),
				.rx_rmfifordena (),
				.rx_rmfiforeset (),
				.rx_rmfifowrena (),
				.rx_runningdisp (),
				.rx_seriallpbken (),
				.rx_seriallpbkin (),
				.rx_signaldetect (),
				.rx_syncstatus (),
				.scanclk (),
				.scanin (),
				.scanmode (),
				.scanshift (),
				.testin (),
				.tx_bitslipboundaryselect (),
				.tx_coreclk (),
				.tx_ctrlenable (),
				.tx_datainfull (),
				.tx_detectrxloop (),
				.tx_dispval (),
				.tx_forcedisp (),
				.tx_forcedispcompliance (),
				.tx_forceelecidle (),
				.tx_invpolarity (),
				.tx_phase_comp_fifo_error (),
				.tx_phfifooverflow (),
				.tx_phfiforeset (),
				.tx_phfifounderflow (),
				.tx_pipedeemph (),
				.tx_pipemargin (),
				.tx_pipeswing (),
				.tx_pllreset (),
				.tx_revparallellpbken (),
				.tx_revseriallpbkin (),
				.tx_seriallpbkout ()
				// synopsys translate_on
				);
	defparam
		alt4gxb_component.starting_channel_number = starting_channel_number,
		alt4gxb_component.base_data_rate = effective_data_rate,
		alt4gxb_component.cmu_pll_inclk_log_index = 0,
		alt4gxb_component.cmu_pll_log_index = 0,
		alt4gxb_component.cmu_pll_reconfig_inclk_log_index = 1,
		alt4gxb_component.cmu_pll_reconfig_inclock_period = tx_pll_inclk1_period,
		alt4gxb_component.cmu_pll_reconfig_log_index = 1,
		alt4gxb_component.effective_data_rate = effective_data_rate,
		alt4gxb_component.enable_lc_tx_pll = "false",
		alt4gxb_component.enable_pll_inclk_drive_rx_cru = "true",
		alt4gxb_component.gen_reconfig_pll = "true",
		alt4gxb_component.gxb_analog_power = "AUTO",
		alt4gxb_component.gx_channel_type = "AUTO",
		alt4gxb_component.input_clock_frequency = input_clock_frequency,
		alt4gxb_component.intended_device_family = "Stratix IV",
		alt4gxb_component.intended_device_speed_grade = "3",
		alt4gxb_component.intended_device_variant = "GX",
		alt4gxb_component.loopback_mode = "none",
		alt4gxb_component.lpm_hint = "CBX_HDL_LANGUAGE=Verilog",
		alt4gxb_component.lpm_type = "alt4gxb",
		alt4gxb_component.number_of_channels = 1,
		alt4gxb_component.operation_mode = "tx",
		alt4gxb_component.pll_control_width = 1,
		alt4gxb_component.pll_pfd_fb_mode = "internal",
		alt4gxb_component.preemphasis_ctrl_1stposttap_setting = 0,
		alt4gxb_component.preemphasis_ctrl_2ndposttap_inv_setting = "false",
		alt4gxb_component.preemphasis_ctrl_2ndposttap_setting = 0,
		alt4gxb_component.preemphasis_ctrl_pretap_inv_setting = "false",
		alt4gxb_component.preemphasis_ctrl_pretap_setting = 0,
		alt4gxb_component.protocol = "basic",
		alt4gxb_component.reconfig_base_data_rate = reconfig_effective_data_rate,
		alt4gxb_component.reconfig_dprio_mode = 18,
		alt4gxb_component.reconfig_input_clock_frequency = reconfig_input_clock_frequency,
		alt4gxb_component.reconfig_pll_inclk_width = 2,
		alt4gxb_component.reconfig_protocol = "basic",
		alt4gxb_component.rx_cru_inclock0_period = tx_pll_inclk0_period,
		alt4gxb_component.rx_reconfig_clk_scheme = "indv_clk_source",
		alt4gxb_component.transmitter_termination = "oct_100_ohms",
		alt4gxb_component.tx_8b_10b_mode = "none",
		alt4gxb_component.tx_allow_polarity_inversion = "false",
		alt4gxb_component.tx_analog_power = "Auto",
		alt4gxb_component.tx_channel_width = 20,
		alt4gxb_component.tx_clkout_width = 1,
		alt4gxb_component.tx_common_mode = "0.65v",
		alt4gxb_component.tx_datapath_low_latency_mode = "false",
		alt4gxb_component.tx_data_rate = tx_data_rate,
		alt4gxb_component.tx_data_rate_remainder = 0,
		alt4gxb_component.tx_digitalreset_port_width = 1,
		alt4gxb_component.tx_enable_bit_reversal = "false",
		alt4gxb_component.tx_enable_self_test_mode = "false",
		alt4gxb_component.tx_flip_tx_in = "false",
		alt4gxb_component.tx_force_disparity_mode = "false",
		alt4gxb_component.tx_pll_bandwidth_type = "Auto",
		alt4gxb_component.tx_pll_inclk0_period = tx_pll_inclk0_period,
		alt4gxb_component.tx_pll_inclk1_period = tx_pll_inclk1_period,
		alt4gxb_component.tx_pll_type = "CMU",
		alt4gxb_component.tx_reconfig_clk_scheme = "tx_ch0_clk_source",
		alt4gxb_component.tx_reconfig_data_rate = reconfig_data_rate,
		alt4gxb_component.tx_reconfig_data_rate_remainder = 0,
		alt4gxb_component.tx_reconfig_pll_bandwidth_type = "Auto",
		alt4gxb_component.tx_slew_rate = "off",
		alt4gxb_component.tx_transmit_protocol = "basic",
		alt4gxb_component.tx_use_coreclk = "false",
		alt4gxb_component.tx_use_double_data_mode = "true",
		alt4gxb_component.tx_use_serializer_double_data_mode = "false",
		alt4gxb_component.use_calibration_block = "true",
		alt4gxb_component.vod_ctrl_setting = 1,
		alt4gxb_component.gxb_powerdown_width = 1,
		alt4gxb_component.number_of_quads = 1,
		alt4gxb_component.reconfig_calibration = "true",
		alt4gxb_component.reconfig_fromgxb_port_width = 17,
		alt4gxb_component.reconfig_togxb_port_width = 4,
		alt4gxb_component.rx_enable_local_divider = "false",
		alt4gxb_component.tx_dwidth_factor = 2,
		alt4gxb_component.tx_pll_clock_post_divider = 1,
		alt4gxb_component.tx_pll_m_divider = 10,
		alt4gxb_component.tx_pll_n_divider = 1,
		alt4gxb_component.tx_pll_vco_post_scale_divider = 2,
		alt4gxb_component.tx_reconfig_pll_m_divider = 10,
		alt4gxb_component.tx_reconfig_pll_n_divider = 1,
		alt4gxb_component.tx_reconfig_pll_vco_post_scale_divider = 2,
		alt4gxb_component.tx_use_external_termination = "false";


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
// Retrieval info: PRIVATE: NUM_KEYS NUMERIC "0"
// Retrieval info: PRIVATE: RECONFIG_PROTOCOL STRING "BASIC"
// Retrieval info: PRIVATE: RECONFIG_SUBPROTOCOL STRING "none"
// Retrieval info: PRIVATE: RX_ENABLE_DC_COUPLING STRING "false"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: WIZ_BASE_DATA_RATE STRING "2970.0"
// Retrieval info: PRIVATE: WIZ_BASE_DATA_RATE_ENABLE STRING "1"
// Retrieval info: PRIVATE: WIZ_DATA_RATE STRING "2970"
// Retrieval info: PRIVATE: WIZ_DPRIO_DATA_RATE STRING "2967"
// Retrieval info: PRIVATE: WIZ_DPRIO_INCLK_FREQ STRING "148.35"
// Retrieval info: PRIVATE: WIZ_DPRIO_INCLK_FREQ_ARRAY STRING "27.0                   "
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_A STRING "2967"
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_A_UNIT STRING "Mbps"
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_B STRING "148.35"
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_B_UNIT STRING "MHz"
// Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_SELECTION NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_DPRIO_PROTOCOL STRING "BASIC"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK0_FREQ STRING "59.4"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK0_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK1_FREQ STRING "250"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK1_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK2_FREQ STRING "250"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK2_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK3_FREQ STRING "250"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK3_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK4_FREQ STRING "250"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK4_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK5_FREQ STRING "250"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK5_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK6_FREQ STRING "250"
// Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK6_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_DPRIO_SUBPROTOCOL STRING "none"
// Retrieval info: PRIVATE: WIZ_ENABLE_EQUALIZER_CTRL NUMERIC "1"
// Retrieval info: PRIVATE: WIZ_EQUALIZER_CTRL_SETTING NUMERIC "15"
// Retrieval info: PRIVATE: WIZ_FORCE_DEFAULT_SETTINGS NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_INCLK_FREQ STRING "148.5"
// Retrieval info: PRIVATE: WIZ_INCLK_FREQ_ARRAY STRING "27.0                   "
// Retrieval info: PRIVATE: WIZ_INPUT_A STRING "2970"
// Retrieval info: PRIVATE: WIZ_INPUT_A_UNIT STRING "Mbps"
// Retrieval info: PRIVATE: WIZ_INPUT_B STRING "148.5"
// Retrieval info: PRIVATE: WIZ_INPUT_B_UNIT STRING "MHz"
// Retrieval info: PRIVATE: WIZ_INPUT_SELECTION NUMERIC "0"
// Retrieval info: PRIVATE: WIZ_PROTOCOL STRING "Basic"
// Retrieval info: PRIVATE: WIZ_SUBPROTOCOL STRING "None"
// Retrieval info: PRIVATE: WIZ_WORD_ALIGN_FLIP_PATTERN STRING "0"
// Retrieval info: PARAMETER: STARTING_CHANNEL_NUMBER NUMERIC "8"
// Retrieval info: CONSTANT: BASE_DATA_RATE STRING "2970.0 Mbps"
// Retrieval info: CONSTANT: CMU_PLL_INCLK_LOG_INDEX NUMERIC "0"
// Retrieval info: CONSTANT: CMU_PLL_LOG_INDEX NUMERIC "0"
// Retrieval info: CONSTANT: CMU_PLL_RECONFIG_INCLK_LOG_INDEX NUMERIC "1"
// Retrieval info: CONSTANT: CMU_PLL_RECONFIG_INCLOCK_PERIOD NUMERIC "6741"
// Retrieval info: CONSTANT: CMU_PLL_RECONFIG_LOG_INDEX NUMERIC "1"
// Retrieval info: CONSTANT: EFFECTIVE_DATA_RATE STRING "2970 Mbps"
// Retrieval info: CONSTANT: ENABLE_LC_TX_PLL STRING "false"
// Retrieval info: CONSTANT: ENABLE_PLL_INCLK_DRIVE_RX_CRU STRING "true"
// Retrieval info: CONSTANT: GEN_RECONFIG_PLL STRING "true"
// Retrieval info: CONSTANT: GXB_ANALOG_POWER STRING "AUTO"
// Retrieval info: CONSTANT: GX_CHANNEL_TYPE STRING "AUTO"
// Retrieval info: CONSTANT: INPUT_CLOCK_FREQUENCY STRING "148.5 MHz"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
// Retrieval info: CONSTANT: INTENDED_DEVICE_SPEED_GRADE STRING "3"
// Retrieval info: CONSTANT: INTENDED_DEVICE_VARIANT STRING "GX"
// Retrieval info: CONSTANT: LOOPBACK_MODE STRING "none"
// Retrieval info: CONSTANT: LPM_TYPE STRING "alt4gxb"
// Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "1"
// Retrieval info: CONSTANT: OPERATION_MODE STRING "tx"
// Retrieval info: CONSTANT: PLL_CONTROL_WIDTH NUMERIC "1"
// Retrieval info: CONSTANT: PLL_PFD_FB_MODE STRING "internal"
// Retrieval info: CONSTANT: PREEMPHASIS_CTRL_1STPOSTTAP_SETTING NUMERIC "0"
// Retrieval info: CONSTANT: PREEMPHASIS_CTRL_2NDPOSTTAP_INV_SETTING STRING "false"
// Retrieval info: CONSTANT: PREEMPHASIS_CTRL_2NDPOSTTAP_SETTING NUMERIC "0"
// Retrieval info: CONSTANT: PREEMPHASIS_CTRL_PRETAP_INV_SETTING STRING "false"
// Retrieval info: CONSTANT: PREEMPHASIS_CTRL_PRETAP_SETTING NUMERIC "0"
// Retrieval info: CONSTANT: PROTOCOL STRING "basic"
// Retrieval info: CONSTANT: RECONFIG_BASE_DATA_RATE STRING "2967 Mbps"
// Retrieval info: CONSTANT: RECONFIG_DPRIO_MODE NUMERIC "18"
// Retrieval info: CONSTANT: RECONFIG_INPUT_CLOCK_FREQUENCY STRING "148.35 MHz"
// Retrieval info: CONSTANT: RECONFIG_PLL_INCLK_WIDTH NUMERIC "2"
// Retrieval info: CONSTANT: RECONFIG_PROTOCOL STRING "basic"
// Retrieval info: CONSTANT: RX_CRU_INCLOCK0_PERIOD NUMERIC "6734"
// Retrieval info: CONSTANT: RX_RECONFIG_CLK_SCHEME STRING "indv_clk_source"
// Retrieval info: CONSTANT: TRANSMITTER_TERMINATION STRING "oct_100_ohms"
// Retrieval info: CONSTANT: TX_8B_10B_MODE STRING "none"
// Retrieval info: CONSTANT: TX_ALLOW_POLARITY_INVERSION STRING "false"
// Retrieval info: CONSTANT: TX_ANALOG_POWER STRING "AUTO"
// Retrieval info: CONSTANT: TX_CHANNEL_WIDTH NUMERIC "20"
// Retrieval info: CONSTANT: TX_CLKOUT_WIDTH NUMERIC "1"
// Retrieval info: CONSTANT: TX_COMMON_MODE STRING "0.65v"
// Retrieval info: CONSTANT: TX_DATAPATH_LOW_LATENCY_MODE STRING "false"
// Retrieval info: CONSTANT: TX_DATA_RATE NUMERIC "2970"
// Retrieval info: CONSTANT: TX_DATA_RATE_REMAINDER NUMERIC "0"
// Retrieval info: CONSTANT: TX_DIGITALRESET_PORT_WIDTH NUMERIC "1"
// Retrieval info: CONSTANT: TX_ENABLE_BIT_REVERSAL STRING "false"
// Retrieval info: CONSTANT: TX_ENABLE_SELF_TEST_MODE STRING "false"
// Retrieval info: CONSTANT: TX_FLIP_TX_IN STRING "false"
// Retrieval info: CONSTANT: TX_FORCE_DISPARITY_MODE STRING "false"
// Retrieval info: CONSTANT: TX_PLL_BANDWIDTH_TYPE STRING "Auto"
// Retrieval info: CONSTANT: TX_PLL_INCLK0_PERIOD NUMERIC "6734"
// Retrieval info: CONSTANT: TX_PLL_INCLK1_PERIOD NUMERIC "6741"
// Retrieval info: CONSTANT: TX_PLL_TYPE STRING "CMU"
// Retrieval info: CONSTANT: TX_RECONFIG_CLK_SCHEME STRING "tx_ch0_clk_source"
// Retrieval info: CONSTANT: TX_RECONFIG_DATA_RATE NUMERIC "2967"
// Retrieval info: CONSTANT: TX_RECONFIG_DATA_RATE_REMAINDER NUMERIC "0"
// Retrieval info: CONSTANT: TX_RECONFIG_PLL_BANDWIDTH_TYPE STRING "Auto"
// Retrieval info: CONSTANT: TX_SLEW_RATE STRING "off"
// Retrieval info: CONSTANT: TX_TRANSMIT_PROTOCOL STRING "basic"
// Retrieval info: CONSTANT: TX_USE_CORECLK STRING "false"
// Retrieval info: CONSTANT: TX_USE_DOUBLE_DATA_MODE STRING "true"
// Retrieval info: CONSTANT: TX_USE_SERIALIZER_DOUBLE_DATA_MODE STRING "false"
// Retrieval info: CONSTANT: USE_CALIBRATION_BLOCK STRING "true"
// Retrieval info: CONSTANT: VOD_CTRL_SETTING NUMERIC "1"
// Retrieval info: CONSTANT: gxb_powerdown_width NUMERIC "1"
// Retrieval info: CONSTANT: number_of_quads NUMERIC "1"
// Retrieval info: CONSTANT: reconfig_calibration STRING "true"
// Retrieval info: CONSTANT: reconfig_fromgxb_port_width NUMERIC "17"
// Retrieval info: CONSTANT: reconfig_togxb_port_width NUMERIC "4"
// Retrieval info: CONSTANT: rx_enable_local_divider STRING "false"
// Retrieval info: CONSTANT: tx_dwidth_factor NUMERIC "2"
// Retrieval info: CONSTANT: tx_pll_clock_post_divider NUMERIC "1"
// Retrieval info: CONSTANT: tx_pll_m_divider NUMERIC "10"
// Retrieval info: CONSTANT: tx_pll_n_divider NUMERIC "1"
// Retrieval info: CONSTANT: tx_pll_vco_post_scale_divider NUMERIC "2"
// Retrieval info: CONSTANT: tx_reconfig_pll_m_divider NUMERIC "10"
// Retrieval info: CONSTANT: tx_reconfig_pll_n_divider NUMERIC "1"
// Retrieval info: CONSTANT: tx_reconfig_pll_vco_post_scale_divider NUMERIC "2"
// Retrieval info: CONSTANT: tx_use_external_termination STRING "false"
// Retrieval info: USED_PORT: cal_blk_clk 0 0 0 0 INPUT NODEFVAL "cal_blk_clk"
// Retrieval info: USED_PORT: gxb_powerdown 0 0 1 0 INPUT NODEFVAL "gxb_powerdown[0..0]"
// Retrieval info: USED_PORT: pll_inclk_rx_cruclk 0 0 2 0 INPUT NODEFVAL "pll_inclk_rx_cruclk[1..0]"
// Retrieval info: USED_PORT: pll_locked 0 0 1 0 OUTPUT NODEFVAL "pll_locked[0..0]"
// Retrieval info: USED_PORT: pll_locked_alt 0 0 1 0 OUTPUT NODEFVAL "pll_locked_alt[0..0]"
// Retrieval info: USED_PORT: reconfig_clk 0 0 0 0 INPUT NODEFVAL "reconfig_clk"
// Retrieval info: USED_PORT: reconfig_fromgxb 0 0 17 0 OUTPUT NODEFVAL "reconfig_fromgxb[16..0]"
// Retrieval info: USED_PORT: reconfig_togxb 0 0 4 0 INPUT NODEFVAL "reconfig_togxb[3..0]"
// Retrieval info: USED_PORT: tx_clkout 0 0 1 0 OUTPUT NODEFVAL "tx_clkout[0..0]"
// Retrieval info: USED_PORT: tx_datain 0 0 20 0 INPUT NODEFVAL "tx_datain[19..0]"
// Retrieval info: USED_PORT: tx_dataout 0 0 1 0 OUTPUT NODEFVAL "tx_dataout[0..0]"
// Retrieval info: USED_PORT: tx_digitalreset 0 0 1 0 INPUT NODEFVAL "tx_digitalreset[0..0]"
// Retrieval info: CONNECT: @cal_blk_clk 0 0 0 0 cal_blk_clk 0 0 0 0
// Retrieval info: CONNECT: @gxb_powerdown 0 0 1 0 gxb_powerdown 0 0 1 0
// Retrieval info: CONNECT: @pll_inclk_rx_cruclk 0 0 2 0 pll_inclk_rx_cruclk 0 0 2 0
// Retrieval info: CONNECT: @reconfig_clk 0 0 0 0 reconfig_clk 0 0 0 0
// Retrieval info: CONNECT: @reconfig_togxb 0 0 4 0 reconfig_togxb 0 0 4 0
// Retrieval info: CONNECT: @tx_datain 0 0 20 0 tx_datain 0 0 20 0
// Retrieval info: CONNECT: @tx_digitalreset 0 0 1 0 tx_digitalreset 0 0 1 0
// Retrieval info: CONNECT: pll_locked 0 0 1 0 @pll_locked 0 0 1 0
// Retrieval info: CONNECT: pll_locked_alt 0 0 1 0 @pll_locked_alt 0 0 1 0
// Retrieval info: CONNECT: reconfig_fromgxb 0 0 17 0 @reconfig_fromgxb 0 0 17 0
// Retrieval info: CONNECT: tx_clkout 0 0 1 0 @tx_clkout 0 0 1 0
// Retrieval info: CONNECT: tx_dataout 0 0 1 0 @tx_dataout 0 0 1 0
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_s4gxb_tx_2pll.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_s4gxb_tx_2pll.ppf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_s4gxb_tx_2pll.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_s4gxb_tx_2pll.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_s4gxb_tx_2pll.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_s4gxb_tx_2pll_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL rc_s4gxb_tx_2pll_bb.v TRUE
// Retrieval info: CBX_MODULE_PREFIX: ON
