// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OCWUFBH6w1UiVQBjgQNGNAusUMp5AFmlWsHLUqOmUFve0xWljZcIvbljUITWC2u1
pVGObC/0igiisVZ7kfP4DPczdbD+WyFpmnhUtvJR7N07v+t56WMfxK+jKUYXDGZZ
zqGbKBA2rcNQDeseLWzS+xv7srs3xRjM1Q026jicJ+Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10736)
u0jDP8EHG8yN7S3zTk6S45ntwBSw2XwNeH6RRf4aCvq0Mt6AJOazHljEj1ItXD/i
sKm1CL+gCtuFk3KivF+mCIu6HPWjP/mpNfIFwiNOnzgkc96eyS7oHo/NETM6t3wg
mBQzV/rQshWdNYCxyBVkSQp4MSvdEN+QOkLo2UYJnZE4f5mvf++q8462Ly6nw1VA
rFHXVwc5P3k9qifkHXOTz0pAVYkvqmbHKg5Le7Cc3gOelhFLxD4Xntk38FWgvXxV
QKcyei7im9G4ElSq1O/e5dkh+U5EC2cf0b2lkZZlU2oycBl1OOCdFkusqZm8dwgC
tHRZUlDMk9KMabiTbLRFv2QOU/Kv9TJJvUCXg0C+0MgQlNWkcAvB5GTtzkjdhZyH
0Kz54btMsXyTbGwEQUHUQZd+nRm3dHfOZfNub5YG+HFi/TX699dN4XgR/qQ/3JZQ
lAwuLxKXpPMjjeT+ysIV5u/cn8zogTluCiBA9m+cwA4viyp2VqUpTRH4OBnb8dUr
tu3IfdZrIlgBXILgZbYFweKARTk8s8WDWj+Cvf9EIS6iwy5GagWg6G5v3by4lp5i
QzLZ4RAcdj0ckfpz+0mKi/FLmYYDS1jaRNiQSmit+QFo94DR6/tEoQjx5xr9NqW0
jBCXehRPIq1b5Mpp86IFxSnvs4Mo4xsaNn6Qi1pqZMH3MaJcp1+hqUAIle/FqbZm
SjrX9RJBZDhQEtuDAeGFTkMq6lSMZNiB18Ch24dQggAmZE0jP3nZu6Nhd8RHkIFm
CONoze7T/obthamlmnrZm1SHd+EIQrm3zQg6sYnV5qz26S14f2VxO+DbORjDAsQr
w+XszbLoT6mUh6/W6sY6Ysl7vHCzX45mxD6I+PBMe8l2E1BqKxKh0KWL4OVAc5io
Kk61BkhE0bofg7Nzu254suLBNUQ+DCO+9mfkuFyREIcxDpPHGrRMPEbICmUpNoKT
q+I/I5B99xwNFc9sc6y5xBj25DPp4EVTIetfDj8J6NoRuigb3SpvjogXua/n1VIA
AtSyyItIShGFajRbK1zaBP6eeIjiEeyt9sahVXcJ8tVC7LZ5A4cLJUX997HuVSnJ
fe8oFMuIjBxSiZrYSvEG5WlBHcrk/xDbCsOFCblandqR6RWimcVmYXKZAHxU6kbT
74crkR53kfKne2A0mzOoXuQE53chKrFqrfwl5X+tb8s2Kc+QZKUwCRNlXd/++vpp
4CrqWa05FGfQBLAy8yi7GAYXiwM+48kIHDjUnyrhlxLGLUzSt86hOI8Mx63yl7Uw
LWdiLCzNxl+ktiWqJbFksEnlO+NPJSeOX1U+bDeb4ZB6ZurcYSMU554alOsp+b+K
KAp7eiNBPVo0OOs73MzwSMWZI87lsPO2aq9c/y6rcFpKHhnDbgflwddMrOAfLGql
IoUnsxswtwPr/xOn8W3gFuDTWAcrW/1f0nSXs4YPM+EPxzRJgxM5FQjq/JzmS6fJ
jDchtmbk3ixIy+m99DAHlHJkpHkeGPTwG3+V9qw/ChuOSCHpiYOCHBE/H1ZeuLAL
aBaDGZipkbMb00HyTP51Ac2NZd+B7BOsbVrl9kFrWM4dKFVR+nuH0aUOIJ/JdRC7
uShIzOaXsCK2xv7CNkfukFoFxaEQcbsalr5BwYoSAPCeHqaIIxZ8OPIQWXTsHtLn
3ZjY3tX9mc3PAS5vddM4XEbu+xTGwhS4ogvoPmsTpw//sUrJaY6Wwy23eDi0Nj3q
L72/xwwWr2V/JJP7EPSvS/KoFat6LUVT4WVvdDZZ9lKUqCN2VvxWS5ARHJC8mZfA
SNy4VrTVk5nr1jmKyk8ebM6D6Zl9r+wMwjS75VAcQUOmDBtMySGoUjhHuGuPVjqX
BxMin9xHjmVtsE6aXu1a4WEHPb1L7uVvoEnW2LWMUDn2h4a1PnugQlvrfXzK9Jcr
AsNxsaoIDGsCyJQjlNriOCRTUtK+ACXvjsRCqhhy84M52Nl31Aku7YCkgvDX5OE9
+CckvHrmZXObicgW++vpIrA2fFxXmnE8s2g3Hg5us7Nt94Q84TeiOKutItP1LWFm
A+cCDZQ0H00RQR5oY8zVhPm7UgBUXVVaRqaPoX9xIqbDXFsV8g/uvHWiU6VtD3ij
J0w0TE/TwTGJ9hFyN+/3yc1nTEfLfUvJlWdsQVsi9ry7i+De2+LIXurC2b2h/3kX
FGj79UE2n3otTPXCoJFbyaDfRIuo7+XRRxDr4tvcSdUIg9eFBaQUmyxBqKt0G0bc
7O2T4CIW0p9taR7NYmeGGOfEgQTnuDc66A0Qmd/bHbCg1YIbZDwxYuXIvYN2wTRz
JViSVpgSpQtfGc3LBRUs5/1vIBVaeqcWyCFGbveEl8aOg3g97dl2FPCMic0x0V3H
jCmKCuZiEhcVkvBaxLvjdruVXQHS4QdfKNO7n3M0d6Ke3npimIK2sS+aZdroonrH
DOBca5rDhYCU+b2rBsTsfvlOS0nj698SpmQeF5OmOvFqltXWYSDsoN4pJWVGxEsk
OHlWT37j1bcz7FaKfsmuYTjsc5/7TQFX66/gjjVwee8o7HmqpRnLl0jOxxTeYstF
oKXsoHJBjxi8JBz+2gLc9zmfx0x5AvzZd2bod50/wBBdrkyh6Lc0FtLbhTBkvFSx
eMgtiVrai4FfuM0WN2LhD3nHbrGt1oIBCznAOeybTcP4sMGSw1wjoV6vwAsrH5s+
8qVpZaNLjYmUMyOHBcK0L9KvMR5dlSStL/EIXw2hQd9arz75phlwGdS/FojIqzxe
xYaaVXV63bofqisaQdppWsk+95LHan/7qUjIcesUwGJ/IlFfeZ2nECU8ofYTbqhA
KFBtTQ6Ux5otbGgI03hoy6C6hyvAWmWHSXcBKeL1wIhPbfOvgdZ1EpIedOZBNWqs
gQWWED2d/nRZRlFfSlj3fQa5Z45K82y+i0DTKv6IBI+QAbHhfZ92/Nctkxmsdr1S
n6gcwYj1ZlJNBF4idBcExefAKTAmsRmpnExBfmmrRYdWNwKJZfyN59f2aWHh6GZF
qLnMyV1BmUFn6eTTDoItaIojlcTHNmW/XvvsDR5Esqeqclufe/dJZ9XHN1oDfApe
ubg4v2oKa4CTZoPa+CGDmWIbSUBSA2ttV+vfci9ShZPWQMkJMuTo/T9cTH4axFxo
ibHPq4ULqBcDXaCdAEVg7hsTxJHaGwGXHBTil/fmDjcrcbSLwZ1oHlkRSFZ7x0lE
BUh+e6/eXYamAwwaQSsV0aJWuNrZaXmyJbi/bbi+on+G/BDDiuoa+ZBhCXgpjJin
xO4C+8nDAOuVIs77hm6nUVAFwXUZR7JWN9Sgj8D9xVvyUoYuAIZ2IJtcYsw8zCc2
HXVa9Vn/WwlAUb/zrdB0VqZ/GC5v6uFqY3tpJze9FsgUEzwjMHH+7hrmiswDVp46
QTjFrkb5In3KpE2WCPYjZboYszyCJq5ao1OV5lz2/Dl0JnL6eB7wm3o6sPgoXjtS
mBR8/x1ddlhEa7LTGuBUfmygf0j9Wi6cUYYDyWHiAtEzI+Qpy5RrrfkbNJpmy6yq
HcTCdQKNn5vL3Lpuyr/IlhAIZ6hNfLby7HyRBxUXCiJGXdx6t7T6yDL7w+FVbl6L
5zZjzGpMEjQzJtA7S/Y1gigWcq5E1IIPW+DKBGiccTUDkSWgCbFAPSCrfHWvifkM
mzO4p6tLEal8gE3ZZmLmqR50xZybbsclIiJA6dR1U0BgRcp/oJwuVoFIFTHChqtD
sJ/YcllpdPkDoJ0gxIZtnOl2JU/bILfIJODdrFo0MlWv+94QlwbCh7jxG+yNbu+/
p7BbAGRNrR77if6i0stbJtFJNO+tF/QWLHcgEjPQbYAIWGjN4bdxP0C4bBh74Bv0
yyHpc81Sk/jiOYMTlChq4yJV2OuMt1NKgw26tlCh4frqMhl0GQuAV2ppzPspczxA
fs8b1ZaLvb/O0bThtEYNF8p9dOXrWz2teg94XqPhkD09cRggJ6s2y2bZrLsWE42Z
NFZWOA2c2MdB/vuagtr9iAh6o2wg55Rifuy60deuE0D8nXyywcT/Zo6lzuymBSI/
lBEv1gLYkB3z29d9D1imkIgCVCaJQQ80wgBvBCH+l1aq0bImVsqJjhPN7Jittdvt
2h6fv0yI2CzuJQGoT/RDlceM/LMrohr4YzTGgVJwCJaqySQUSTxWxVNBmsX6jT85
D8N0WjkOYvHWycMlTuGSYTlWDWQDAHSY7mjOtbYXYqg04KJRoC1kcdhWf6LOFldm
j6RbmP7drz4sf9cFZUU3Z9mvVsCr6dh+aziIgVupAqYd3OwaQvi/mcFxd7Q8IOEC
81EqKXBION8UZiihOHlDDbcHJ3XdyYoV6l0SGX4rXDhFiitV0uhxX5BwObB0k1JJ
JrjRM05WbkoX0CFUPQp5/VHQK5IkAvLqxVPeWOHGGviUDMQMUVi2lzxRrQBGybqs
px/f4cAKkXYZ+49IAhRSvfi5cGDuWrsofNAtV6zASc/kb7FcUEnELQIC38dzriUZ
TvGbFN7W8iTTha6UuVONU6GaF9F3W0ogpTd2zpCHGPh+kfxgg4fPS7epqUY0+Be8
M4aqfClbCxw6I4qEgqQddAjfoxIH6KV+d/6k/+eqe7EiHwupYF1lNtau7N21W25+
7hEmHnrBCkaS0TEUtCoe/IYiayavqX9hBw4FDtaxIibWcZ5H8MhmufxIq/LVGNPg
k7maeXDk0C1lY8nXqvKfqT3kSsyKzjZO8GPWup0Bbkvz1oKFKk8njweIiyyoJxeJ
A9mOCNvoOa3LynAFThEBruaYr4HFpHBjMCXOlhp26clrU6ayIn7q/rTeMakC91WM
6o/dadpKff+rtIOqRn0QgmeNMiSQaAdZEtQ4pjuuz8EOZwcSlV7c9iPEZOIP3/1w
H25Fn3rY95fgFyQ6Ek+B+WWs+N/GzeSiD7qXuqR/jWq6+lTp7oSbTEsClYloK/fn
fo5EpZ80JG0xPm8jNt55fcnJRHASJD9UKcXDmhaRrLLfdETKM+d0dOzOtieANxwQ
dqWuw4EBEEmFvS/R/yAlzv0+P5Ornp46bXjlOpMi+ef//dHMlhm1kiLeozV8LrUt
Bj9aH4qriBkbyNo4OKfW6IM4K/zJvX5rY8cCZZIVXWOB8pvyRUth9rjYjr5ygMrm
1yLLsYXEQH6KV4RXph7Pr4CbhfijTkvO71kuSGkzz+bQf3zeDPFmpNay/F+Gz9e3
ddKGjXB41JQVHxmsLFFbcHDuZA0fng7Ka1tO5eXQIk2MSgUVsrkUVishuptn3cHn
Okx6B1dwB381UJIT/ay6vhLuRAFowwGMiebsTFDKD48G1w8N1jHdk0yn8HPiMbYb
inIRONvZUsC+WvZWzNrHT0lt2gFiNJEYfPSJGY4H+DSOIB1X/+0N3vvJHIs1FUDx
3vXuBJ6wptSrF9oxHsa8OjTzovi0PmYmLn6S6EL/R/yGSCMgtxJ7smWNii8Ozqb7
/daSbijDhpupSKu9qOpkSrju9LGV+DAGY+ninAswoQcjqJgvPIjPsoX+hLh2WK6P
AWJprWxcBoDuDzncwOZJjKZhzYMYY6nCPY58anctX8b1DI4rPec9xKCCqy3AIU8b
PPHE4RasepJmMKElBPDLS4/yZXpjN2BqECmu4ofcigUi92luXVyQBI5cC8KHJutJ
LzlHECgKdBB1jGfdgQyDGlWwcAeCJj/02uNUGuZYMcwBW3+t+b4M38UzChBLFKvI
Y/aWgi3PSyTg0mJc8c+iL4mwrrU9RX9RxKAmyA9sQPSK1N6KHW6IjXKnqw4sXAIh
zG3f6BDJgqVaRh7q20Q446sKqzaRSM6kl5+084tC3ohe5PTdsecCOQXOShJPDfs1
1jlYwTSioMMibNByrsIB8QJI0tgo6E5njut76jNE+d4UxhtD9psCBqK2oiXMA2Cn
yzpRZ5yS6OyCmSPxa63AOPIebJG7ZoxhiRqQ5mPYiZwhMSidWoc9Q9/25wY8gKy3
ALtdUnko5Rbb8wSa2B5GyTWEGENp19ipT7txh05kt4iOIbLPxFC0tbSQ+XeK+h+S
V6fhmf0DnOFdehf/nXZSAPATAPz7RQ6bYVx0QnNjCTkWYveKakzIkQE9/128bhXn
GXZ6v/j5aalNqNI8lRdrHxdqGxhd7XQhfc6IDmXD8M2jjhh9XYeSylWrVU+dDfBe
5FNNxdpxyNC10s4hkQ9may3UK4lPblt9rkcsM6ejHKqA3it0Rp6BEYYVgdFYdeeD
V0was2Z/zUgeuQo8tvKIzFXU35CW9cAqDgyvq0g5J/dg4NoTibNDXERQF2DzxHM9
gc1FDjDasoejdc0q0wm1imEVY7TplZ5jTsiFbU7ruozE2ZPS85ZzC4+s6K7CT4rv
qt/QW20WWlb5g2QwX1+vXavnStKxQQ8I2OO9mbJWx8h+TegVDhED1oRujvkezB84
rxNJdCwrMh1FrKBMKJ1KjoevvpUgPoa6fisUYK+6BMOpletTyOYgVq8HeiwEJxJd
RQWewzUihsLpA+z9jSJwQZUc7gws7xfuEpKHg3ShGM0Z+1xcjI/shX3IP9wHwFz9
ba/3AJV7D6HcSkJZstmebHNQShhSEMZFXiTI1SzXM6bRyPKhOr4XsWcD1euhtYqe
fS3aH3BaXv9pSLNiwbbre73NicrsbC5mVwg5/9NdfCuekIoqjkcqpIJ30g61apt/
oIgoYwSp0IGT+era6ygUk3mMyoKLMy1G5lOQwCXVST6NLhqI9jY0576I0XV3cFoH
DK+Cr9KEW7vVXD6ceLasMVnOInhfg7HeeYv49g56NbLBczxIKpd1OtxsviDmYiuq
MPGMGV3Cg7XSjDTkZ5a8l2EZGbRs1m7JgS2Gc4EGhQ1P0Hf/qeaORFGE9rKwc0Tw
fl8RwusAKTrwejcnZNwsHihzLn8WEwWNrsadJTjicipb9g/GrBicOLwS5zX9GWoj
FrwJ6tAxlLRv5BcLbewDIWJSebFfmI2GoCQEZeZPt3DJATuzvnRQZA27kDzHBrBH
I0TO+MQj+2HMop1mQlMQwyz0wJwC6xIjvIh4IB/nquLoDNxayWtiIkLEtO5M5Wgx
wqhebxNhml4wmgle5SMVzwtJa2YxP13dtDHYiKuHbur4Fwl5dnP7wpTFb8Uv10g8
CpxlAueMpdSo/wzxLGW1HTFcy7H4KLiD0nW5ESWPFqzWtdJa0sYaFrD33a5sIAG8
XNUZZgcwlGBFmEZJsed8dA6VbGIPSvNa7Av/280CI3WoreK5SGIQ8Us/j1j0rWAa
RJEV5ntxCSuCSjWTYYlC6W6qDjJJEig6XgRSPEkWRnPQOIF3nJWiNr31WmdfWkV6
354bN8z+xUBKf2i8fsuyRILVodLbsosU8mLPsRS7H3uYtxT5eKPiOp7+Hy8CJ6cf
24OHFbC00j33HRgqKNIIWW83Uqv09NuEWxqiHcGvcc1RNd/5G/SXkfJZY2vfA1Nv
GLbfPTgONs+5WApldlpMe6kApxw4TFeqckTeqEfk9wWnSznaRsf3OYXeAanvFmPl
bcBbxG7jTAryC0OjZfxBcJL8gp8+VcAbXZSil6YPeXQnkx2Q502yeqlIYt8JafKD
YV1u7vHe2GNDJ6ca51hORsV0Q/d/tz9lRUeqWyGzxL3OWb0Ay8h2cTTEhw1yaDTh
KcqZH9pQn4bLN7NBT+ql74g2AfjNlt7WuP5Ww5DvFglbG73iwg4xbXuN7ue+6wfM
b5dj/gUdk8943Wzh5sR/lZy3CPtPRDjdQ5YQBi6OaNPCqYkqH99tPKBiJTeWo0Ev
lJRQSKTWym1PmI6YbKJZNXdmbBxjXCjYldcIEKFhuSSHICNCWDrnI+mZfyk6EIAp
AE2gkSsccRdbImGj/yZL4wpjpgnF8+/3rqm6J04+lD6DGNERjZSugvbW7Aowi3zi
awre6SfmBxjxdzVC9dtpGw9d11L8891SxNv8tiOIYzY4bcId4ZJJXrFuH8VXdH7U
xsT99vI2fcJW0hqmDtvKytJwoUiVZdFv+aQo20/G8WPotgEqwdCvQ5g3/FlYmhrK
z/HKLfTZPuTYQKJrkZF/WCFZKCFyc+4KUCUWv9zPR7Q9InheH7NxB7KoMdaiziMo
gUpmirQaUZblpUf5TlB7qTjYt/fBx7825mLEpqGL6AIJqCEHP8TODTnZdn1d+JKD
7G4WqT3V9pS4O/OmabX03Dodug7Hvn90dE1jHEqhENDmJL3G714NjmMRJCgMlL0J
kJOTMwdRU0jRGMYXb5d4KJw7GV/NENvq54PbfIHYW3LuinWjjdtyy9Jj4J/29T7I
Y4pf7CTFPt+c2NxJKA7tERloTXT0re37cgZliLOb6xH0sEr7TxPo+dG6nf10iRGz
zOlFcvZ6/TwM4VHcxo2fJWc9dTtaqsrMKDlisTf3dDuJN6sQxbHoGzZLJevfrR3p
1BoqbMvExP6+7EQWDDv8+wkiXJi757CIwcYfP+2L39dlKPI4SevYDxsaC0nq5EaG
Qnu9UgYOdPSQXZJh7EMzmU1lxcdP26lV5hfm3M+ixLahN98mFd67QlVigu9YvG8J
1gw6cEJrKjGb6EBSejVBv3mD/NVYYAT81wbSrzFF0GuuJveoxIDUUK4Emd1OOpD/
Zk8DeMRlBr7Az16sJjYsR3tcNxh36bXDTM9oxlaKAq3jZTFvraQCf7gLMK0NIVMX
vRy95/ar6pwNfZcC5tTRvqKU0KdiDRVh432ZtdmNZiLyXkWYxR93jEPlBijbd5Au
L9REEHXc+/p+ro33gT2IXvtvedJFLhimN8HupznOAd26ZUOkM/bcxOsgbVk0avoI
wdgsRiy2U92iSWa4Kcdgc/c38FK4bojFyuJBUgihx2O2dJ9Y5TmzNd1JJ5dIipKk
lwfk6FdbPlamq3zZeMMP4yX0L5eO3HRzf6Kuh2DVo5eJzDZgVFsDZFs2kBHBPWUO
kGQwjd49jLTIkdr84RPMsJdQ0DQYSsYS0vWF5WsoZUGilgILlJx15K1cQA0fm4EQ
YLR4WhXboUMaZj//E3EXKw8zhRBfSjLZazYEOd8hx08NeFrzcq1uPjtxS1C6tV1E
+nbAkbV/CayNWjCIpzpDuFWUA3mi0Fu4KHxuYDA4rRP/pH2czMfQd+GaiY2WIIR/
/7lI3VKATK/cLpQrFReDjCpIPqq8NkCfCEfkiVjFx93epCYe9KZPFmfCP7zRFnuY
kwdJuC2ZDJtq4D38TnBaKjpaYiCfbE6rFP5Tdy9BVj0KCGbYNHiHMX46S9YdDu+h
wqgIr0aRX/Zc5iiZ3z3rTIPfu/Z6A1NBJbuz/Q84yDEXfOt/HK/xDMKjkr8vFWJA
DMekEzBfSOCC2djIC1sZVEppvp1a5ORVGHWSLUiZrmxsnNLxipu+/+kvb1P4aHau
Iwxw4In1dr/+rw9DNKpR4xiA+Q2VNOC8nmdSeV9IBv+efT4fpA2vd4wOAiC59hEj
wWbF1BthM4PmFvtIG+n7v8emlFVZEIYiD9HDWAo4xeMBot1scMEvByDIaoLU2XET
mfD8HGQTar8EhP223Z1u52MAvD5xH2Z2r6slwKrSP9Hc5g2P25TLRnYveaQrUjfo
q0FZpy1QaYIYjDor6EnLdBFgJXVWAy31lcewnxHTBdZ7mf4itD3oNKyE5O3jcpzh
0e5u7g00mcKq7gRsBB7pFt4Dye6qsSeSZnsGXXHycBV1E0CY7J2eq58NzVtVTegW
wwWWs0xsZdHJ/Pd1t2Lvu4PpsKGsD2xyXyn2opg+xt2cDhRNXLOc3I+5pg9rAWAA
xSFSt8pgsoPj4POEmgkG4XUZ4D1Z+qzSvDAlkA4RvbO9pZhXYmVXyUGpPvU/7Aoh
T7/6oj25b8jIiuJ//JugEI4G2XPJcDYWNMbWyWy2k6DncrJvfWLG0VyQo7VjY9Xr
CiCWTp0f6XIetgH6zZihBBNMKEzA4f3h2cbZgRosR4SWRu1RZ+qFYFLSY/iK6Dh+
nNOxILZFJ80DeV1y3ZXUsYexoBqtArUDTBdK3xikEnuY+3L4ScMqOJclOrFyKo+3
WU3PQVVU+xwloic2OAhIE6LSimbgHDBE0k7CXDa2eY5r4Wdz/BEqpjDZ5K/IDbdE
RY+5o96L/bxt+NCyB2lVxyz644slxBuvBmviWkXOikU7qLD4W+lVkcJ7e+Zo69u0
fR6eqE8MpsybRTQ8tWEhoWSiKNH0YvPSEeF5hBat5JdOm9N2Tis1yzTNSRk0x+OJ
6Y7J6W3mC4g+fNxSrwLP6llrVqAOVIzzL+lKi3x/FJKR/17nVL4xM8NxXMwTp8La
8HgBs9+a22cxgkgIG38E3k9+wWMFfn0mtOGDTjLoR+NkSBhTahmaB3cTykxW0jn4
g/XKp7rbrCEIg580GwEKVQy4KH1O7W7mvuTCAEERJ573PFQmwl374tvJ7851P0cd
aRXbFczc48u2Awxg4rfbou7bWm9F14Qzch5VM+PdI7Ui5b3qTZBETwIzQ+xqVn36
tjx9FiIDU1wfxnmQCHjMtKlqJBE8yCDYN8tLL3JLwuggKJHHWF8vRO3XUhRdg4p2
/5+TqbxjoKuSJ5JLW9/qtssw4AQYbg2KGq/4UPhjE5UdD5nEjx3sDLpLZKVtsCC2
e24QqmGqgi3UNYjUnKkcY8HvEiw4g7k5deGseFC9G1B0opW7cQyvHnpqQl4InfDW
itklafClYLiftFd3wRoijmlCoU1RI+24Y7nwSlxKeXnye+woWrJcsVIB4hQDfcWh
2mEvIqa0ghR9NnLk6vk8FjBAPTeCnS0h3EeOSmB0FTYmmBEiXWifRRD00xK1qSXv
ht3CpgZrzSLAdNjDjy5K7+q67Eyj5SuogPGDNtpUXRT2bUGbxmLLg+0VoElI17UR
RsofgOiF0S66rpiaFtYvg6fFtU8y92WvzCvuKjhSHPKTqaKK28pGT3LmQCkn2HEf
jDXNbWUfgNdEFft6Be+xhWKyjxlUVrN7w2+xIabKHmCEZViSrRnI3dROQ4fE8COd
HP6simzB7bTMjl8LBS8BwgtuUcjh8DmULuOH4dHan8MVuXbQNWkaQd8w/0eIxmj7
MJ9BdPilHTg6Sfc9nUwQ+orIBG79Rz7H6vMvS919NYbRTJM/D1HIw9TjHc4Dle6c
uGeojLHihFzVeBY1TkFfkRbiTHYW2Pxnl+2MwoE5/z6Ti52gfmZy8zk+tFCkNivS
8pZXQv6eHEFU5BrP9oGt/i6JAX89/cKwbM61DhbLnI0v2tnb9IxgR+TMCcgqRA11
vGDknT3+zaRBUWQam/MfXquQPSQmqL9ruh7+8j+OZF2iBf37xIxRrt8qn11wq+AD
/GtV1X17PVGyPb5m2sLlTmQJoOnomsi1e5KfbAYcVyMFlVMWxZ5VZBBwtlIujPpV
ne1YzrxA5gRuR0rFGK02IvAsN3HAfDyrV8SBSwWPOubmjewzpXt0fyYG0Qlzc0Ao
ywaSnjbOgA8O+8DrMvopyBZ/yoXHVzFZTYroVrfiUYDA9p3MH2YXte19QfxWNGHd
T7tpUrVBXh1zLn6l23Yagd/IOUCm1/i/g1zaHowhqKzjgEdbE0C3MvdayedQHsfD
56jWKS4aIOYdQVBXD+KLt8zmshv6dDUtX6nzTWABDqV886QAEeZBZNkbXdjcRj60
uEKaqY8QnzBWAOY2TqFgH19tGnGM8g5lJobDUMtodWYaRApLPgXFK/VzoAwkp0or
MxLVtVsYwklfTfSqtiS4SvLmz9hhFNrXVdD7jLZ/+aQytmo+665x0CGYpw0Y5ufM
p3XXaPXd0A6jQASbJXa7J6irJJA16jg3ZU+6rtFV58JD+SOC2YXkidG5RpFeNbO/
kNkkCJfv9ctrWTSQam5tHh7o2PRxaYjTxVjd9P1dr62nDZtYLYLbBRk/N+DmYAgP
yhIkbtYGiU6oh3zj+8QT/zDuVJ7j9HBBbtqnq6Yz2y94QIuwWMq2cYw9OMIRTEQa
u10uU5XSpeaale9F/wbXC5fn5OIHtQuAEZU4aU+y2cgdUzzrnjNWyEQU6OZNlvgt
c5oQY5rsScsUgag09/aaTRUqjVOj0CV2UM0oDHzFLde9MllFG/LlsqNsdC9g0C7d
9qxFibxPDzATXoQUPuGNUUGkHV0yZwd6Eu0acdpP/n9eWeTjsymo0LF4z4dbFgTF
Jo11Psp+hcQwE3TZuMDouxNR3f8OXSJ5YAhtc8QAVr9k/XWRGPIg42RCLz0w1Fn8
hStgrqkmhkBUY4aK7rHq76YPaZFroxzdk14Lhfxj8WPEerWOmlA3YfVMh2MsBFVK
SZAP3awK7nkzMMyiYaRnxqPPoAA1vOR9Ctxk6luR40cs6ssYlgQUU+YN8ZnvEddj
C5uMjvC8/4oASHYi5tDLEOaoW9UflyprdMwvXBTG8wFnFVthw3b6yhr08DDet1Bb
Jb8pFNs/gSX2CrI2yoUMeYp6kH8awekWJSKQjuUeL0hP+ja/iWsusJoUD8cIVRNU
cL1EDvNJqLaSVPWCp51iZDfNIyKjNecBHPmoOAC85ypZTrr/iSFgKEUckH9lIecH
ZAu5WGjyQsjD9JNMaBYR8jJ+TQcDM+uA1rD1733fkcEQgxN+SBgTmYmCXXfokm07
GEfakxOg/ELpSOFtKnNtoCNi+KgLc+YLBmAKRbDO9EqLAO52BV6Fw0wCzdEMKl+/
tDhEbC6RlRuMvA+mJaL/6rWx6SssfX+6JnjfK9Xhyzfbp7aVBnvXx1zOE5bKWScB
CNzw4GeW6id29PwwU00JYhRazOUNLDoCWafkZ38KeW3GUFjQ4PnoRs23u+82bgwk
dSXMhA3pvA/orPVIkUzk1j2GIYIkvyUcJj2n9l/2VpoXW63unjEsKIE2clnu4Gij
SrK40iEISZwA4xufT8YS/ACL0xABu4cLxVnnxHhZYRxelkXPZc8wzA/C6c/SsIJM
1KaJEvdr+LztCucZAPfTR3dlDSN8TDjBQTObERtY/1+LdFoMbsxY6dSHSb0Zgg2A
9L6BaIkmn0RvN+MeLMf2dk1MOFqO1XGRxpAjEZwqa4ivl43nB310M9exx+2+zUrc
5twi4jsXY2lW17xQZDWjA3tsnoxeOc/5ZeanqJl6YD8QsWpR/Jn2f6eRcACCwWUM
l6T9+Ehfh+2+/OLxImA0VJXnUi/6uZs94juVLFhIni+UW833YLzM8rKOpvqHHBMR
mljCdSkPzPLV3A7KLehpcLkzd4OSrSwSJokRXkoRhJnwx3ER07xl2ivyfqvzUCIA
oiZe3gtvogS9Ee3Fu1i4EzOCxD7rngnvxU7lVl/sRzgLqUZyhj5HBIJN+5jUTlqV
s/41K0DOcqsLPr7sIQ51x6j6gcVRGD0R7iFJ0DU0yL5Y7XgPD66rn2Ng5EeqElhX
zGcQSl5b5i0XZRLVeEHcOAjvBrgB53scyGfL4XM8Q26myO8y48zlnZN2zdUSA89o
5wBJMo2fbQ1jxyZ7riJqovnZwH7yb3hIJEXGAKwhlBW0UixWzsi13WXsijwcK/AY
CD12yjDtWOpEczfLsy5fTDyWYjVHwljH3H7hVbYA/l5XBwL8ZXCyguaep6j1wCc3
jMS2dH9jaJLQBCfa9PRKE37eaqzjcWSW7jVh+dNZGSEZkKpnhNOxN801DvdsaEWp
0iUJ0AU3XSFfS94kbTp5+papAmI2NlbfafNgkAkjl7071FU/vSM9J0hL0hUbvN5q
dXquSh2+PfsFMsM3/txLHw2aJw7Qztfg3e7XmEpcXVfIVZL0LaUlD17m9Vi3E5FS
QG+DUYOxJSeG0BKLgOXRo8Fft1bXwy/rUEVMyH4nOzWGEOdQ8yzorua0EcjpenZE
3OsnmqTyekX+NuZV6FZJ/JyqTxYsgbnqA3BK9+7s4FNsdBGMxjbnPlbTJObLH4fN
lwYUZ1jxFaAeCSe/7X3ItQ62s+m87yWNWGAuvYJgHTinasWh8cQq+ZV0gBTf5xx4
Ysj0wJf56PSI65B/H8I/t+cdUeAwfOez3jCJbf8BWbGlNFykZwsUoVrrK+aP8Qyc
VDCk/nNljMMAkKwDF7vj3I3ya0CNGpiKyqLt2rNT0Qqoe170/nTRRqdq42EC8fgd
tJQQ6bpgos7XCa0OCqT8/d9JIKSzr+mFg9uIxJP6AiH9KuuJV2ZZEL56rGENdLaQ
/JpebG+xUtHcA5hQHp4TRc41vsE0ZAx6ZMElcAUGSOGNe/IlGFaJ5edDEnIx5e7q
ZdZuEZtydGNALiDtnouz1XCihkxeYM+JZck9LiQYFrIzyDPlyhgUdqz+9GXO/fRW
exXkzlWvlxOw8Wxr8fXmE+7kTQmWGTNQzHavBdAlfmMiUGY4rvUTwsbOUHRCdOae
ZG/s07ewgIk4Q0Rwq3jcgfsyMJD9jhLO6nXPsZKjytE=
`pragma protect end_protected
