// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JjDT1JFWSUrxGqdHK36iB2Y72lGeNhfarq2v+b3XPgYLvfVnuzY8jVD0TzsR5kVu
vDVq/VU5Hk6PAEf+uZIVgpnlF/pi3O9SInPWK3UaSNMgTfKZaSlkhNniH0994Vc9
yLWWOWaQ8+G0hixdCnn9mw3qC6gfdS3F1jygONfavoQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10544)
exnAjHXty5bcQyDY3DNGmW30TsmHHI01ld10ycyiMk82pRAqLQd60xDmhtWB/8UX
igOOWOhpZW2tkogvwfV/bfmIRac+MWiC4m9P4zOCaT/AIqN95+es1Mu3xZiMJD0E
x5wDGNrsjLu0uAPRbnSmoicUq19mOSZssEktEddkRGtYVT993dKrYqmr3F9OsGZU
D0ZWVcqKZ7LDivEH2qnQz4UhrUYjsh08wwkSOAh4IJ7g5cweh8OYRDWiKuwppksP
pRirjYABKlEpU6uiIRcy4dprWAczjTD8+QXOfp6DfTt27fr6f8b1iqOBL1tDD3yB
bqTJcYTfCbF/4Qb5vlaN2m2MTtb+QrlnbdrWCD5ITmQyqw7Z/dDzPde/XDvM+s9o
Wappvvdw0q22/I/lQ9/454+cloCBcRF7xJXbSqqLeTsNd9yNecy14gPs4ZSTMa4U
Ekj+GSZ9U64t6WbQQ4V9vnMsVPEl6HNAUwK3baSen97BpmMx/60c1tBuEbavrXrG
Pg8wvzM12ESX+9z+J18bXBttxGDwp8zylykhmaLZKD7zYbeUnBOziCKrhGzB0Kun
6WWRCphPwhKsAhXpHoswgCQyYojwmO9lKrU5cWrhpW2T8u2cGwhezYoz1SuKKNzV
7gUYen9sOHpChnSV91E7XyWoq3VraOj/6XD+zWzL/k/jDAm6lK+GnS9xv9+ZMj2n
Rtzi/CmfHO2aUvp1NZsCnJpcGVekEEL+2TEYsHYCZXinEk/V5KNHUH31DVPLvgKO
3NEZAoTZAN++iVqqoUby8Hu1JsbK4VCTwkP4usOho02pIgLYWwhBMsgXVXf1X0tU
MeoLMZbxX05fxDrJe08MaFdQBcMe7zFykJszGefQV0Vjnu6dKYohHph861RMcRhV
HKRTfLzTMbvMiRnEoa7PgtaBZ6jcgs5Gb8H/1etOOote7Aiz1a0SjxZ1lbvKjuaZ
WNV0/SJStYD6V0UDlP4TunoTxNRfsA8EhJDYUQRM/FG7oRBJMmeaDMvvigDF7Dj7
nKPL5Tj7pJuZh3P1vqyPubPoHZoxmsxhTJ369Ixz+FMjxzl+Nh1wAeku/5MgQRPJ
7lxV/Om4avB0tJ7jSo8aHJ8l9IzMELnkdjXx6VYXcucbvwd8EjFyjW5MghIt9WNZ
vEpspLGNcqpu7qzz/wpRNQvroHL2kuM+QVXyrRKSlqUjQJeNRuOMcTKciyu+7epl
P9AZ8cgWVt2Vxdfz3zEFLCcbTmqXLIujmSdD/TbLMrxYZgNzrLyGLxWmrIPwGssT
OUldDJ7iIFbgQl23frYiROxu7Fy5AVCb8YqmZ0NwppwjCQFO3kJAYUhk1oTk6Kwu
VcDpOKyrFkDmLvLSuCf7onsAO8zProimP5Tj+SgIaPYl2ihvPOYH1NLNCoVxWaGy
JAdOpFfTOJFjU0ynYZJ/jfFzuGxhc/luH/d0UH2w+8STfLyXWYYUt0je4n6ea0+N
qdCDmWjjWAGTdcXdnQ+f3QlD7v94af4ur04Ihe53tY/o0Xe4mY2DGvg4jH54QLB0
/JQZIxfjyg9vLNkN+aeyeqTQMtfrozjyJltJDxHpMrKaNvmiUNBHnO4JqQ1aST43
Cj9MMQZ5gyck7Zhp308hjB3vFWYLd5OxndSnkkP0j1a6p+zR5Yw6MXKeawdKZ+1S
kvOrFo6RtP/HNqUFvplBqBCS+D26jVsLh55LTb8HbRw0RmKmUaZxNjLaJdZm93CG
5AYlJneEkLDOFcbSMpVdZBD0v6M9FWfz3rUxpfk/WWTbzLVoCPZixvWGmPeUj0eb
BCZ7OwaYmHAtm2o5cGwuJJt4Ku6HPM52XAKIJUVDOOctY1WGDb/e3YflfQ38UecJ
X1a0MSVSvt+iTjzDZ4OncNW/h+v0ZaV0NjCb1qF3K57OIP0xp58M/2OEtlVk8rVw
0P5O6DawiDb+DPyhTjpmSesHQ65gkiLPpyD7nwcphVVEcd2ad89BK6B/gMFb5hF/
rbdqfD4otYYLW+3sT/C3ZwzD9hwxzGvNe9/Onam6VnG5NsXbhQRW7yP1JawtED41
Fn2AHj9VSIE27BVe0sBW4ELf37YATcVowkaszt7xdOKkzLogli4vwbc7b96vnRlx
BuiwrGyS00/JGrJ4RZHnC8cPyUWnWV1T2GH2ONVTKqWOi/ZFHiYBWoEbLq6Q2f/O
n2+8ylVyNwS50vZKijY5JC9CIKpU+a86HYgl79AiM5GR2IW3Of4dGERrNowiyO0n
8BYrmMzxk51fEjMYC/r5ZkInnntinlpVbz9Pt706klVUqFc8gEEIeHYjdo9uD8Wg
CurGS8B78YN1YwjlhZKMANgHVs2grWw1WWBEIVYaaAhNoYicuYSz6IrZ7L/Hshla
yJuNvO5NARl9Cl9Wf1k24Ds5EvEMvHf9Sk7VFFKUQgY7drggUU/3lZcoM7/Mi1Tn
VlzZqw/WWxLYvtpn0K4jE3BjXHgaeS67KlXsEq9MjoCNuN9aST2YlS/TXRlAQJ0S
RZC24U29FTyuAUWuC6jSlvs9eeM+DhYOqUFsky7560NMpolUlaPgBI+5uBPOqSbs
jFJk/GPFOU++sr7hKhG2cgamZ1Kf324plg6PSHTqSWC8jpYovrWGeWcylgjvGR6O
axCpG6gIeFqcI1HCkd/XjGJt18kGrqpLzkw3ykIOJ5RWSG9OoCHOg5qff0ww5751
qSb7eybNU5RN8WJk4MrQ6tvmLxCLHkYyF+VZG4jhSnuRDjiR1eG6CsZbBiAMu96j
SKoCoPr3BNefuTbTMBWiFhYstgLCe89GsHVP5gNpNui4cQes+kZmd+YuStTRpStl
eLnpo4rj+ps2zoZdLl3BDcwjL4pD86wDLp5ppE/9M8XwcFX9HElaCdMyLkkIoxMp
cecbqVtbsq+Swt7dBuugylMhkZMKev5D46F/Qp8mh48l7YzWo7eSIv0r8Y8IvC0u
EnXiyRMYVE5f9enZSH1kuRGgRqt4wtwUKCs+BkTNryy91F/7EN5ETsBzY4G+vhEM
HmGQkKuQmXrqY6C2dA/E8zT4ryYJ387pQ6HXKYqPlvhARvPwsQ161yYktdvaaL9H
9PsWZbfLPLmg9GfbEIbmkUd5WUriPQTHZxDPuhL7PBHO+sIr7CK7nI2Crcn4Hhsl
su/UPoJECswfL58W1SHiV9x3BvzQMuY6+A9epAc973B/2oR1Q2DmqrwaBtVlNtAO
3QG1ms0I4OzkVpJc6IF02Ofl9u6JuOZArQa4UXSX4945k4BRjebhYSfulGeS2nXN
5Sz50VQrVTfUGT/7S2KivjG7i4YOn5+2ewIPZq1SYkdqlZeu08vWKcNv751hpyTo
fAg01LjDWB+jW4JW2DhbACi/NBqBbChoGS3cyT5EU7y/p6/kDmFogd7CIVLZ07+D
sIocq1FsmUXpX5QdK9zQHcu96tOeO/0vGSN7ZFk/rSxoOx7lRcN6vY58m7jpcOZF
rnIEAfvlSCBAbpDUml/290ZcXg88JIvkHBhI26FjLtMXKFOPLZcxvaB8k4vAiMRu
/m/4LyQMUziMQgHAOOjOAio+xUXnwx7b2Vgky82AcUzHPsPVK6F3R/Rg21IDXdAB
6vKOE528k6Ur2RgwfvhEPG/8h7jsbvgeN6xPX8uwYSwo3pNUvFegkKsqspxe10S8
nX21vBdxHe7cpOQvu5MQdUclGdYiXbDWagZoIISeKbb1cb1srh0Va42pKnPA+DlW
D4/vdXax8H3v0w+27t9+sxfKtU9C/rNXTEMRcRYxRZ4wtDFwRbqg5EGgJfmyWGp9
5xE6XHivDvKDwQBWSpBUuptZ6oPLwHs4e3nnzuKso97FWC48D/MqruX4/vc0JeKj
6GQPehU4Vlktt+5ANm3W0NZgL9Ps6wquOtC5ybwmYMA7ZwDaLjJXn/ADbSkxxxsE
FTBtz5wREH5Usf1WoOcKS6gC+9dDP4FeHziQwXJnpAvL3zVJResbnYAkktMvKK/F
EAS+T85qIWCgcjy7gLLsBGJNMOzRd+wcBzBo4tOxYJa+66WlYfi8dJRoBiWaXZp9
cQcuc4fdqxNvpLfE6i6T5YKkfwww4cZu6ZHUWEHPRa+jUl8wAk1FJVp9tifwLUZ5
br3v22zNcQK8CiPWp2DybHITaYTMQ/4oAr+zf2AO3UelnTxnxC5nyCLfKbyNgnxt
JnD8ub9EYDJWCCfGDV3zpBtQfydBjpIyKkNYeE9Gfn4ZAW8TGK8rPRjyadbx6Yyx
kCwebBWaQtkLwH2AHmblG1IpZIbZuaIUCk7k1gzlRbXql7R2SAnWHWTayayZBtm8
TkJGqmN9ciTLPxYP8gYrPj/Ky9y6b6dS2Bfam2/v0nfN5oBOrg8Wkbt9DkcOUmPj
fD5X6t4pJr+vHoKE6CWZoblp2j8w7t1yIYr6Zw2MJUTGdzF6E5eYz4NHlmt/8uKL
s45fy1WSE/8HdLM2Q14Fc/f/1z4OzARNBhRLVhd2UlWUO0nJpnzW7bokiuyv0i2N
RC/9w0NCc+4dtP9IHUZxKT3O89Zus8fcXm76c8zviGZfVHqeOC7R3Ioeg7NEbYKq
czCxU3PAg51d6LzYD0XjNXoBGbwx636eUQ9W1CyLAD6yG+ycLyQtLppm0HZDgWTF
1fZGXsXBCj7JaNWapn5/RfmN0q19SgLRuYzuzFaaTXH5tJlGbWXKhcMOgyeUHNcM
w24/cZirYuD9kGgWODJb0o6fhsCOFF4DSgDs7Od8vVstM7Ojt4G7UWbyf6ezxtvY
mJnKEq4AWf/uhPvG69E/O1yJSgt1JxdWK8kns29Ax8Q/J0RikGDj+2+b9zrCBw7S
PuTTmsZWH5TeDwXdOd7TOqlqiSfbyg7V/yR1o8HT0HK+lXd5l8mvHXl6SZfpj1Hr
sq6xb31/laOe2a/V8qLuHF86QPQcPLrrfkAGANBJKb6a7S9i9cdtaUveWss2d8FB
xA91SYoS3ufaofjYZWIUF0NiGodGyTngqi1D3/4pKqG0gzHeUY14Ld+fIBzeJ5zB
RbpdSFhG/MqqXUBpH/q43Ttv7TBB+ave8t1o2MiD3PFl7ZLpbY7FhQc+z/B3MQ2Y
vRJqy2NgDVXt7igc1jjUNtix18EaWVBXCuK1BuJ+ct/cdbIcSfVEpEUr6ThvV+et
KT3hqVg2rwQUeyG3OItaT/ZQmG7TWCK88PquJvptUPJkWBrnHzpBmR6ALrlnTurl
V4epNLkZhQXNxXPvcWWak2qwzR16eVRVlJ8rrZ/6L4A3LnUz7FpBJUUlj6viaD6f
MK7bHIdnC9yT15/i1RXdlnV0aS3dPHadTXDlMSJImvIm+WmzTGLzaGZxivd1hteW
0UASoAxQUtKKrjR0iMW5Zfg+bSN4cDFBp2DtH5Tr6O0kj/6uw9gumKpYXespb543
WiPhF7RVEY/JzgSADBX8H+TzTonSTzApYh1CdC1rp2o2+jT06bP+ejxAtcCkAWF3
GWPhYAGn30zRYgHBxGAYCwJYqUnQ1fXBeyxVmoU+SU+/SMGdBeAH/gPzI6vrEJd8
7nkI177QcbVWkhxGRI0Am1rk8XPPmEqz3rPe212c+hNnxNYAVblOD+2MI7zhjPVP
7ap6LcqzTrUTYrD0vztXW/PFBHt+5BafbTiP040utWEKJQIyO7ZY16c8+ZzzHYrM
3l3lZaTP5RKssaUrZnQKR0bMDe0qJQoxIswBGMOsNecV4fFsPthwPRq7uPmr3U8q
mFKcOpwLJX5jztwB/uqa2JYneYMqICbM4VJijUs+irpuD9ED4R+eMirteL0sG7lp
p7hI8HZev7zdJfZgl0SYKuCiIKvm3sqeg1FkebCwS+hAuYZeVoZ+8QJ9MP6tZZeg
GeLfg/CGoeeEqg/CuWPJjAqoGRcILqWTWdE1Q5zd9ih3eD4X930uhY8OY+UGUqrk
2BwToSw1FLCmcXItztiQ95HnXB/lHzu5MKXWH4D2SlNt66f0zMgm+Nth/Zu0yeJQ
rgGPV5ttNPyvQNnxLB3Ku+W7rIB9FpRCGhmuqcqmeZ5JXVo/Bc1BoMsRI7n1nJ+k
1U/Z5SSdAYOx0v0Yme4v8tjP0fdZ4Ukn8s5ufOgDNg+Aq5rErhp+UCuuI8YvfH2X
r9bPisL/udYH8EK8ZmMSUx0MzZF6y5GAp6Ka/gtdsymWTrFz1pEsGpWbD2hnFOuR
JevEOjQQt6TocFvdI0Dpp+OSkaZnnPaRR/uL3+N/7wYJ4dbRwSP5ahD1fwnCbvSK
k2KO7Z4QGRvetOU5nXIKFQdM7x6LTA4v1XQQrF2Kjmr1RzXQ8NCy4e63+mNIsqYY
ST0EAFqauyXxfjxWm3jhAdVJJA5Mt4qQQdjTA50quLBlBQ8YuTwSu7rQaGFwnVii
wG3piNRSVWQqobdIl0grg62A0NSPFQeT6R30QRYlU915llkeGAV75ec5EmaQv+6w
0+yS0V+NBw94iaDCRUcFglXoCDA63HMzmz25dAZRpWtREJoq/5LIqKOW8FMUAWaG
379D/OlKE2VOwz1iOfzQQxvOElKWVM7GVNTj9Dr3UZCmurG42k9f4rr3odoiOUP0
0Mz4IlkiN2HZ/02eHYlmUSzDfNRdjc3OrPZc95xsTU+x512SwgpoPTF8oGlX5/U6
lywFh8lMmXXprm3g9l7ScrriXwfGzqVuGgqQtN05LKS62Y4rlcx87KKMZM8LT84E
RuP6mmXZt/wYk1R0uikAESNGqDVCgzsn8HxHpF0aInyiUbkWOj8dmhzQfP/+LdoE
Qp2aWP19WMTnCGMwXldw51VdNF48PeF738WSaKuHjiXHRfRNkPZyHZerTMIYuiQg
UGI6wbeig9Eg5iqmoF7GJLuNHXi2BsKLOWB1F3EKqth3rMoHHU82X9y6a+hIR+6d
IwXqqaLskcPNv92UHf6QWfa7udPg26dkPjx5QLYzHvd8jsHuKKa0rvMqpqHM1WKw
MDlHw6LVVsN0vki/gcokfsVMGoCH0P6q0J3/giWJC8alx42/cv2GwXqGoFu4ghCc
6+lUZtoFCihThKxo4yGaDTmt0njGFHGr5uR4ruQuzoJZSNt3l0jMg/AvxHUoL0CX
PzbenVwvoDAU2B8bU/WfYhhO9g6WpldX947f0Vdug1fEv7dsRi5vUdoi+Wx4CYcg
GrTjT50JD2QmiwAYpxsV4l0ZZl99Z0sS+E1vx8RrjjjpRtPZ8jT49Te/slY+1kDg
YCu9upp55DJMrZqi9eCI+ZOKIXIFnGylxq12OOxY8pEfuUGoveOBPxhQx3ZAsbSP
Tgf7Fs7/0sSBLFtSKQl+YUwV/O3YkW0et4um1qVMjYJUMb9mSsMpgM8l82psveSF
PqZF972c0d4tnH4JfvQ+Vk5PoWEo81xZyQ9sgCOMvzBUvWFT/YWcs3HpQHz0TPV1
kYQoSUbeH20kVO2BkoFqv6wWccIu44QPux485YaQmbYwQiobsScFfBrzBCA0po70
HaZVD2RggiqybMWTW6/rn9UT0qxKv9zUty77KYqESdkpbezXyFqOO7EuVW3lWekV
/Avu1u9XEFZJH9HWxkuBfuIcGW3fUx1w7DJglMKlUW7xQUP2yi1pMAWOefF7vxvI
phq4PzPDvc3D3UYAZksE6qUJ4hxprXz96TGjmNWDeGy7wb/Ep0kPMAiLHIcoPuei
JmyMPZRcsiw132SMRr6Z2YF1LG3vTJcJTltrYtsdCYs1r2+vim9RmxARFUruig4r
xvSMgt2TixNYUXDYuRTiFKNhHIOUDZnF/QT7d5PO0LdV/YClkKtCU4F9COejJQIa
HOHoffS4V+jtlox5vSrUi3aViMZj4oAb8FQJ5w2nyS7VXh5qRXfGE6GdfQUlnUdt
ncyDZvuu1gCOw4HsMU/n3FTfzpqFfsh9XJVWBXtXqnp9JMBuUgBlLiZdcJvreeVC
12rLgtlA/2lQyQqIMbW2f9n2Lhr9BzdeANY3eO5YnGpwzDUUV2MghG/MAqk5H26U
WnxeSezQH/G0K0qlwPi233zljoaxsL0lOBTaxyRPrEob3dPqOGXvZtx/3OlGWDIr
nre0UMZkELYKIPX89TQO+B9NMuLj1Y1CwW3khR2JIn4Fp75MtZ9KoAv3HwH2yzyu
jJsY7jkBKyAFzyjq8OezQsg/YTsP4DM0s8JSi62hMycqdBK2oUz/CNVuQKElRUkG
MYzgfXUajwF02OSKzqCdU+C38eXXhUeuruHkJAze/LRUFfrR24UH4lxSiI2nFkcr
l4/YiLdqtozPjsLzdRDdosp9EY/O8tWuP9m70DD9DbwOwD1Yw7HJ7y0hFTDQwxHa
Bcl9YsyKC8HY9g1pul8lnYXIkC0Xp6n1w1/olAucrhDBmOBmXDJmFg9Rvowy1Ljj
V2X0a5aYLxAA0vzyD0Ji/cWSsVfkM1kiXw30DCKB6eS97xFNVB146Z3q5MasJ/Q4
Xthq0boKzoldE5xojtSnCZJ8bxTPQ2QhBSsog4zxKtVbSSF+FJXGDT2en+lbobz4
30RcBELy1chbkoslGbMneRukgm29PHrUX3CzeUDh0w2UoSWiMRtiosS0eoMAjLKW
IrQHGMSmYU7e6Bs7+0HSTuH78Y+GuhbHkbEZj8QenCPbYISDIRb3DiohenbNR3GE
E9Ur3OshEsyWrHxxGMlScsUhHN+BzVs4T1170qcKl43R+OEw8j0v26esNRlwMDAw
++zg/3AHGfVof0TRLRrlIvrCM+VpbIYkaUSnTZvc9LUTd+szJUb/q3SpPLBkrTzm
sDlj0T7CE5XEFE+ny4W56ntfN/YMRrEteZPYgOYNaDeEVxbRgMmIrD6iw8gOcynk
jfevtEbw95NKkSOhNjAgmfWc8FGQ07T+dQPjkF4tUlENvCK9NqCkKVRnNXlSqswg
bNf8PPqShvPqwZdPV7iKqgnnp3vqGeuudRXJhwiAkRme9NFyNncrhJl90JXaWM3h
RAKxLWbbyTK1/ik/aNHNdbtOjORbNR2rFRlSOkk73xTOK/3XVa6NKjKyUUpRHgks
n/7XCxACTQdz4F/cncqdskdd2rQyfU7fq9T5N91mIYcDmJx/2TkyGk6pKQypBno+
6/zIXv3XCgNYj8xTtCjSvdTAN9Z/KoTdgNSvKUpsgbFm/BOvAlv7DuCgeH2qCjun
TCx+zzx1trYEQ42FtQeJ3MCjf1YvRLZwSAkBzewDQY350U0GdzCJhmzGXPq+NRUs
8qjpyYxzRl0ptQmo4wIz0rEkOtRd3EbM72feVfzDCPChIEnHICHuZc9sQ+XfDtMP
BFn8WUN+jrkdk52uElXHAPtiDMbNQDu0LQt5OCtcQH2wyYPV417fAxUnm5bpJlva
6+N8/+E2UFqd1gwCeKclEeQpO5+B3A1PJMoFkYX0xb/ZVB/oA9f+cNG61EClCVVe
WTc8v3l+FoOmYR5DrN1oH4vlFzrbDgs3d15+3AyVJ6lE7o588fejV6SHdx6/UmSp
DHjAplGik1pbZMf9yL3WiQvR46bA3v1p1TxuL3pMDKl0XsvQ6qiWiGPOPPVevTr1
7+QfP16MT+VPH0GF5Tg7SRkBCwmbpNCz4+wJw1485LYSrjc/V2eqbNlpu7qV0WiW
mZpdjdZStvTEaug3IgVTDPAArkWbVrEMJnSMD7+iuOn4mSh1DJmJrQwbDWeqVyz0
hn7tJ0P4XXJFR1FyaAaS3abFFNgQEUitwma8nvChDEAqbiALjX29Y+qOXVcxhZk4
kKqUIokETO2tp6KQyDV8/NMoW7FBZYmGwJsqzWehP6gKjX8mCdJ8QHo8zv8Uv/8m
pBp8U8jFdLf/zHdkIKwR8IKE3+gd2tYN8iHi7QpowAi0cdm/pQVnSQ+elArimCbe
OhpXHtI40H93WTHw4K7nr0knNful7UJ1GG+2nPZjjsm7hmvTbpQpKWpRk0AfqVJe
v/6G8xqGmtl4GzteJzEBKOAziVg55fu0CDPKIA9fIPDAWHJ0VlJbuzzZUrx9nuvc
lzBChXy8wAWEHtILIEGUe9Stuk4kqp7spXPsusxHuTUFG4tef5gcNdzxsDwaLI6I
GjioccSsEYkvXG8oy8XVT6pjX4rd/5/uXVxK7TOTrjLvTUe+j+93ADe9Z7fu8GcE
Oc87BcgLZi8wGUviVG8ckcVIu8kMA1jNT3aii55cystJwtbST9kRRvngJ1/2ra4d
hDCHkcosveeEvxR3i5SVjO+QfLg4AsdLvwXOUw7MdSU3kdgeuN3uTai++HZJrnW2
XqHhk5UtTSv7gAmkFu4plXREPLtnKEjRfVpkUcknTRLIBio/9IpV25Oy7PIBXCtx
ubkfydvJXx+4hbNsI70voHkD+kDuJ12PfqVgsR1MERVRHkE0PaKEl7PreN7xS+fk
Jfp8337m9UlBf7KF0z4ds6+7UQx2uZzZwweOJ6JvonrytvRmo3EMa5+es/rCRCRo
OsKQTINFHeUNvK5nfNiafAh4RpC8mlZCL+hdzvT6QZ/+16PYKONXbY6FVOV7whyy
BApsTeAoYZ6D7vTiSMGi6Y3CM4flhIlRZ5BkCWRXQCUHmenOWciL05OcFF/hV302
xZguUN7kdbIXz2lCkr1NICTkpuk01tVSG7ilH5kFZpoc3KsDCuUVTT19Zlqm3FKe
CDxEWOTx0kabqHJA52WlBwmZ7yFTlC2mV0sS7ecrc4E76gWEvqAKrO+iWYz4MXPF
hI0XNEzPEQ3ASKlh3CHIrmRCfR5G9cPnkk0hDYFEf5S2w6Z1Fsu/mNN7DFhd1SSx
JHPsclW7Zp3lmdycCrpJUoe38DrrfqiD0IxVqOmoH0pExR3wJAej8Ot9snzC/uto
kQuPVk4ElbVlMgaZO/1ypCkS+uUQEK9djjkG3XzfzKn2jUwhwX0iHiuH939mVCGr
CX7XPuOdnIST6DJ3MExh6NZs+Im6rdRUHPMgsIkOUH6o1eVPv7ggSY1L0zZbyfHz
GsEKDtDaHC5AZXhUnk0RWYJmeGiRS6a4xzEEdGpeT2QA96atfrP1ijCe0rtq+8Kv
pZwzDSTDHRex4vwZX9AkPP3Ks6txCH9dXXVSG9ofFyWi0fEvQJOgjRJVETH9WDmO
MTpnhssvp3yBC6aT8H96Ors3Ich7xdlV/xaXmN1q7MECbhaI3bZihSijqMzrTDRf
TXJSddtID1/0BbMMo/wvPkuZL7b2YM5QIvGvu1c1qLpLwDy6B1p03xEb9ZL/rZM5
icLDvOZE/mAyk8+7n5v2QuNtden0pAw64flcNyYGx3MbHy89YCsJIorVevjSznsJ
DW0vHLlvboI4OQhEBJcEDWB8YFyPSthX1vgCJRKROM+ZQzu/f8ye9Jn9MHkxChV+
mfXdvIfFz0JTeRi0NSqZXo4+vVJdG77UN3iNMgiVyZwQ44ia6ge1sUJrZyysr5pw
fBaeBYKRCBEbgcs+7Fir4vjs6KmkAHn4KZ/z+ti/qtUjMdKUg3x8+2WBOJq+9L3T
HujsFMT0N57yhSEFgvIxtSiF2eZxbP2U2GpWhwz7CwYlnnJxRGhfzx5MfQhuR9/H
UGyUVgIhSr3PSfyEaXh4QRhMBc67PaPLPJlTuld6aC/KKZnZom9owi9I6WSXKQ0F
LBRGGlcXLiOsu76aSaRVzfhxYCYw3JikXrHEZ9jo2RUT+gBMciHueJ/8r+j6kFM+
3hMxumLRjzaf3ZFoB6Q/c/pqgiuyX6PazqAZsnA7BOG8XXIR0xEeb++DvbHrPKBQ
8aQMnaPowqtTnr78XkFI6IZRDCKzeGFfvE8B6AOmMXpI0pBYbKaI6tdXzwIbvH+i
FFHlFgOxfS8POijF5ywdWd+f8CA+FzAykgh7E+SAokARFwtD8xvffvchdTYb2Eo7
+iu/G3gX3CjLrsjpQpUCzUoXrAJWEmx1bTNxx//HjeO4ma3lfBXjgi6K9s8KSUlX
ZWt75p5i2sYAWx+JoQcRQ7pmXkhpwnIeytw45m/P+riAMSXSlThjDXSQF+skUE4p
dY6rnwZhQTjg0u1TjX7CnPhEm4kitJd1ZyklIwWmLw2sX0xiE3TlEZlo1tD9lMEO
QYF8BYwZ5TU6YjgrUjeoq+NFWXDZ1OCjMXo731KsYNi8pxfGRbaLLPJLK6WfgXBQ
YSWeKLtZ8u0F3NXEMj6uHophWIFzOnBk16eBiAIELfl3jyu1q4O9mK+i1dSImqf8
jZsXm5MMxHIS1riQP3rM5cI4hcXKU79NtRbFHa2Xwii9mQtc8TFQ/ycC41nVJsU2
aEQ+I/Hk4ZC4DioZK4XISXBhU7oL+AOU8o2l7BCc8prTozL9AOcEgZCLyIxSUUfl
gzucdxeuCRxlpJ3eAbZfwbzLS9lVi2FuUury/q7G2nqy+CJEGdkJQ4pGk/70l1A0
FTHzJFYqCM2z9gkZ2U9fhJGt2cc8vIWv3/fSODtvFzUUSul9fj701oP3UXP67RA6
E0c9Hvhh4rw8KOWLWbqWowYbYATtFCFVI58wEtaAthj8Dw9XmQTMkrxHjaluxbCy
4vgI2XhCDtdkeJW6m/TRMsT4x8pSeP51weg7/dhHB0moaopKpeWL1lcxKnveBe3s
ggYkQn6uNMNHeSn6eSUKEkF6YsMklIXbFP52g1NSnCeVQJ/CujHgy8qEADBytTvw
TBiErFYIjIsM0ryUfNcsAZOs9w+0kHuTXbcyIvrUZJlr2WA9Css/077UiNV17OB5
gsVykJrU2rbc+B4Q3X8JWzRPE6ZEhrZhTGAxpsKNxQrQzvlsfEd4CbpZJuoR7NZL
5XAfo7XsYYjJdrEm5U7civEzZvt7bFmy6ZhCPvphwRmhHtCoN9yth1tIAlMl5UbI
NY9j8qcxHR0OhKFP8GzeU60mwAIWjek8ZwnO6M7uCRc0MKJQVsQIzREWHN6rjWkn
mWAy4OjItjxS0LOSXzsZbcb+BfIxjAOpDamC7jGKXYrMANvY+QPLF7N2nB5F6BUU
jPLpqaBzDp6NuYf52RpHP+584KqsJpT5k9btFw6kk+A68jbPLR/OJyt5Nt0El7Zu
fHs1UTufTU7nac+QLn3DQOziT4uIP98uAkjaqX3OQPTePd7b9r4MK3/1EEZ+3xET
YjL2hjz6YYqYkX68D+e4eCQGaxy8uaa0EtGK0B7zD1f4UFzZwsZPpwz3RrsaE7cf
TKcicqVm9mXhJdBkkFW9S8CMu31dQP1+jnEypeeMihBBZyWaMBJ0KeDTUKcoBIS3
gmz2BO1gyV8ftBDkokpMLgN7sKMModRCjLxTR80pUryav4gORaQEpF7oMqw2ztAP
KkHO9gvfnV6ZGwI7coegQBEKLqsImATu6ymur7NolzZLtryia/hICDQo0e5KHiGh
vM2CpLwN6rbi1VbvDRUW5yWPQSK5hcC4SUwWz/fxC1WlkHStGWekFI7nNPa+ERuz
v5JXFDzwkdNhH32yrFPIiHnhLd4BXELERH99rvD6LkcPuHUXI8PVVyszurqT40uk
0+fmx8ZsbHkihyooSETb4Ul4HJ2KsuGyfTQa0w0utC5UKOA5FTEuNInKHU3AHh2z
DvlaveavNCgSEraLNANfDEd7UEgdUCnFydBH2FPQiOdizcGLYAaWSkMvV412g6wE
ZWuFXomoyYwNSH67a6sQnosJFxHw4miiWwcO8Yv0uMOV65dF3hxOVQOLy72+N+hk
GDyETMkAN/Vy8dcedr0cbl4wgV4znBZ4sB35zeAmykfRS6xSk2TxsX3OzKqmayRj
N9s0kB3vNz7AjI4CBQirTvamIsltygVe9CEE7PvsnZJJ+F1mwDDA0QN+MwSdKM6f
wnvR9gDBTLSnWpRIuCPxE9rOOyDprtNFBpSpPzcDgese62N253KnzFGq38xFoIxR
wYwns1HS1NQaY7yFw/aQLd3do+5HnhnG6i349ONb1UbizHoJ7gZ1WRKq6/SA7Jry
jlJ0vqfvoM3sle8EUZD+v789m+SDaG8YQPtK/w3q+NF+9+MLkNYPGZ6qpvNLdYV/
4sIla3ywDhOCipdFoaCf4ShU3c8FC4nbNEv71pjJBtpNwMjaAxBC6GOHSPFG1aVB
Jm1yVlMqDldkoekjdJw1tX+oTwgMPDOtAJgQpEAt8M6WTFUebCN1cPwu6x2Lafs+
pXVG8rrdXuuwbrOB7fit+BjMJgBczh26pCCg348cphg=
`pragma protect end_protected
