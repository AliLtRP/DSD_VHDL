// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:13 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZdboEX8Ftid/qqlrzClY5XoFpUhCzT1soF6gK4ydsamVR3IKLvWvb1kf8K1rJrcx
CNPPwoCFry2KDp41GTgfS53CBc8VE3N4UwIslJ8SGZezVNvYfVLXO0NvTv1dSeDC
djpsjh7jOUP9elsP1/QpXhEfhAM7z8TjAQlCXCGISB4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15536)
HJaf3PREceKsxvFMi29OR3IeTPKRA79/EYVyS/SUi+HrlCKOCoWQ/1zW0XuGBeBQ
MMfM5cU5UkdfOHqzhJPJqsiEHisRjTYoQFQb5JBJWwRgqu8xJERxNhi9ceiVJO94
seW5ruNqLXltqDeGvk11+VMkVBEIuq0BSezno6qtKy9gdvmn7/4pFUo9ppm2Nsrr
nwcmS2Dy9dx0z8zM+7/G+3CrXEVO/RrkAOdn//fEhIszzGACbIZAMK6tvoxnPfuS
aETx12fUMr0uWfn7W6EPoF1dSRZleBSrF1TEnqOu2XJyW06w5gKTK/TEEg3o77SD
fwIQ5Bg53ettmOC0XAxvBrQtYKxrGHqPESgjk0/7jphK94LXIbuyy9PxBvvfG+ZX
h76xjD7mZppdS7lz1T8eRTd7hYlk3hfnOWI+/fo/cT612VH3KxACY05zBavUjblt
P+TxlTYFup9oLfnPhtGOrFcARzyfSjoJPO+HAOQOjmzJlNH0PsgqMlor17VozQig
Ri5fiFiVI6lYuDAmfK5wfUux4qAbziew+nzAUI9NBxgaAEA6ezqUrQBivM+EHNwA
3/WE4pFAinhqyMjjaA6JTGwKTQy+B4VWqhZj38zEMfHGyounKyZzxz7265PK4GZu
impjlpFrOM4qDeDRbAjfBwTw4qsdbWcdGzK766UEe6S4wpjBYI9Bloc3uIRQB7HL
HayVFxV4Z8qsthDDaPeuv0cS2q3VfylOsaFnZKBpoTtsanPKuBL0+0tKcK0zjhxU
FoS+DAzzBggikEHIlNQWQ54gAnQxBK0ugyVLpT29WsilaDn8B4MLIL7iY03leQXZ
WMxE7M9VdKc1NZOeQ4D3r+ErrUOYpqfTq4IpGvsu0Q9eoJ8VQ9Ls+MDyamGap2hi
yb3N1mM0TkeLpUI+WSxnLQox8xD9nwjvHi7y5PtKJcSxQNWs8QqDniIQQaFdogst
YFuz23iqQrTIrypeRYGlFoM+h4aGbbRq6qH42ysMG6L0YVjuNK7LiLhT3mU3kdex
IUmVxjxwecvQ1RID9/r/UxflGydvSBHD/sx6F/ofmWhTsr/RaR2e1unfNhddNBGw
Q/Kvx06zeqTp3jE6fl3o2bERokPBQVCOIGubY7sGhCde2zkJrlyFGABYXWB48s4m
GQkWlLGmlcBMMOdGnrF5B5NidUuAPSvDfNcfacpvbVDILNHCFD08RNB0Uu8Il+Z5
kZM7Fc6jHE+YwNNmp0z3XfbeGksKoxOeJo3+FY1Li1TnqVEygcTIYEDYOY6GgGTg
Nx2rU2hKFFdXhF02bD+9LNVW9bj/qVnutL65dkQNaP9Onb72OrTw3A8aNFI+x9ZK
w5zfyJbp6USQVBL3pvSLqGumf4XML/kmYA5aycD61cflF5upUlBLAcnbVIcy1wAb
ktb82UKwTpQ63oJy5Xv9DZB/0rMCR3/hEH+bOpsEJWHgIDO4e5FCJlv+4ivF4ZlM
dOetGen3SyInfENxQBMSjmTvvno7D4fey4v9Xr8yenMCAcPKMeScQFclJWF2R0rk
5YZ0uQ6bTTUazUP+JRXQFhx9JdXEOz3aK5BpWkC17GPzsnohVjbPmkt275NJ7D32
mqvg0xdnInVwpseBowyzfXRcG3wRDmJX6CDurarF8SVNxEhMPAPWj1/H6kasNKj2
h1Re14iCcsbIDZWgARS18vUO9F+eFi0ZZbp8D/a4uZil2v2j8Y2sdKy7yScpT201
vOgu3ENgx9TO96TCYDvNhICtb1KivIlYpK8YYqFnjekclMx8CwzDlnp/ZbYEhMXp
PQjpN7Hxaw/vUAArs2sYo9wLFKkMN7EhMZBnSckNWnoZvdonn9Rz4rWf8ozZfTvt
yVYP2eMyyo6Djcfdo5cL/M/ztGOzjEuAUbfAE7esutTsqFiLIT9UPO1GW6lXJjgT
WJZokgv1Y6OVi8jpOor/ApJdZmhK/uHEZOQYVCr7RZ4TBclbE2rrKEMiuO3e7tJN
IEmY2NrfEZSpPtdGqNnCY97ri+AeEpRT+vxo07I5xr//3VnHjiLJL4LET7VZeC+c
vCPG7+Jdw3K4R+myybAscrY6FA0+jbz1S3zRy7wMVzq4sUzk5mxKjlsBVv90E1Kc
mVy2uvaiPXGH6s8Z0pL7kaIt4Pcutw2rxTeuWJwLXi73XWHZwjdd6ujBi9QE/qk9
DqRC8VvJPy5QWqavmX47H5HEMm6uhjUQPEJ2O3LTIJJpET45Yx3ihglY7SDW5RuE
gO2RP3SpTV5zDkomhdVrj0vHxRmuRWra16jdOGb84eLlZLuQWSK+x5LCAfHoXNWQ
4aoWHqxEjzN8BlKksBK5rOj6Lb1uCDvbY2A3Sjm4tebOQcsEwaFx+0mpDiIQe7vo
+Uk/M73gnzRco8NXrqjwjDmI9lBvGVUh38WVuHZ1rP8JeMYXAgtRD9/d7e2PDNEQ
Gi99k/gOlLDgTLOxtk/0D/lr2kt7vcvkq25j9JC/2mdKCeNbDQxyY0mjJzHm/qEW
Ls1kaqGJ0xgdTDOBl949IqvyT47f9oEVz+TIPXNwbYKzj+JFNOT0PQeAU1c3x9IY
FFp0RBLx6hRTPmT3PS3QyUrvyp9uhU49VNhYJ0NelLXlVjmDCYwq1RCxy/sQ4YEd
qbXfzSDhE6xuAlbAzq3ddnuLo4Pt0fvAMTZbToNmlG0eyibNn6GLZCFHNSFB0an9
I023JNuUZG9AChnreWFz5S+PVqrbhE0wVs+gUBZDuSKJiJYZrKZuQPehn35X+A8i
/FdCVW4rky8rng/iV1gSBW/Iwx7P4/ykeJYdWqBkX9bvP7HpFrw4/qGdsjLN4BWx
fAoQLnrxhMuJAJp5B3SU0RphBlF251AI3Fjhmn6vQa7cwOSYLBIX72QOPWtAdV82
gl0wKnpuoIHHxFFvHllOIOufKbM6hunu5unPQR2S5chJLUDQUsujETzuouhjHzwX
3hA/4PRUfsugcd+ZfIJJqqkft/+L+0FORT7nVJSDOjEBgZGAWI7nlGLyBOgNspgK
5hgMiVyAmhFW1y9zlYcyKesmG9jqmXpzxJpWi/RZZwgu30gq7ATHiBtrvRU5U8HJ
0mgFRkp2zRS3dknmREyxFy5bTFu6XAeNwoGYCu7gm2RzDG5/HYPrT4VQ7T3gG9ni
QSMDVQgbWkDS42+DscAk7Z73Pfm3rgyOjwxGP8/OdMinaZVA0gj4nA45bl5gxVQf
d21e2sF4UzDSEvzQPeo+HW4AIHxfhhWylCo95RTPa63YrUYGe1aCflTai5xB31JE
hkKie5k13vQZ2ej5STAbNXMqFfNjINO/T59pn8iKJpMsSXpx9Rc0ZklldKplb+lm
Qas7dx9/BpcZt1+dmhnsG0vG2XJNOWgwbZbDx9yHPw2V9xpFS6liXSKgImuYjDbh
UZAPL56u9AtLgWnBTtrNWcXSoCXXF/5oPFL3ACUA8vMDrJ/OePvR7NZdlKBUiduV
SZRcRfYalvoY1q0IDPDH+aCkyfdb2XSgCbyzY5n5NCQ9Di1DjB7yHm/ukMIBv1kn
mpi1mGYMRmZVzObpunrWCbWOjL5ycP/bkwuqXcsrg1Fgap01dtD/soZZrJEa2nx/
CYtbFEHT59vz0tours7Wuu6+ys3DPLol+uvbAVHe3lDyFRGp63qwum0EiADB/Hv9
oadqWr45Za+GhLkSe75CTMqdE2x7zXnvMKyWJhwOaq8vO5x3Hd1WJU5iurCh5dsE
qNVkPgBN9UO9wi1BnHgyY/2gzOJKSRWO7r/ZIYWtRNcsKBK1EGzOaF1kqaSIxg6X
iQ1clgGL2SdgZbgBvh8+C03ynSHGo3F0bWcNgDl6UWpaw5wPexwDm1UZadqcmgl4
gHSudfe8/4xysg0O34skNgWn1UEnWu+3mi7UwF0cDvCVFXiwIKY1AnhaXOpSmxzG
nJbWIZs3C60uOrsE2Bun+CvpLx+71eCp9/ahT2rwq+O1VLlpvteCcZEdS5KyFXCx
CcBZI92EW/eeSzRMfO4B9idulvoLoMO8H+c93loBXpc9iwAtCPqyXkKgWlMfhguz
X61JWmrcfE6wXjBfcoGzAXHkh7g3pWkh4oZYns1Dcdiz2+5L/4DqJ5nlHJXjDWhd
8/CLkdodmCntz6o/zq27WdudJfIrLZPkWrC4Bc7dHJ6CPp2S9kCqjaat8QejiUeo
zesA52l4GOpMtxy5dU/V2257FQJ8GOeMfnK05LywgQUP8qG//tEeTCXrhBr7C0DP
wB0nD7nFS1aqc1IvtNGy7d3L0n9n3yrQlUMDBCSazNOsOZGwIuB26+J0KXMGNCeD
tY3LnXsubwW1xxvqpuEH/bBXzk0T1P+EMjPzNBbJBpAfRt/dd3hVx30DDZNChHL1
k6UY5o+RiC3rg4e8eirVZ7dzTvdJxiDTzgGy+UdoQujfnGs4qD763aWfeZLsNFe0
OfOm0oRV59U+ULbTbys5toq+9AfnctFtt+s2RONro766LfdwGLdrKyk8IKFM28Ay
0SKm86xoLlK0cC9vsB+OoBoB6v4eK0Oincy+OccjgSgh3mc6gHPadLEGkh2vyX9/
h5bY09IihZDhx50QuedfvQScGUVJPTSJPzScseiF3gYhFd+oxLb3eJn+Dez5butO
PdwmMYqRsda5oz7dIm4bHmzqM+3fIwsPbVHHRFXGdHWPuvgCq54tmqG7SEXPUX8G
hccGUmA+Z33azSv+S0Sn3vBZDk3bvELXp/Y9dwoGqmicd52scDm/ZH/rcDUS5yal
JvJ00q05wGGY762k87mW6VpDt+5UDMZm/bXoOCQ2+0VCGzRQ2Rzm2h7UwRMAX4iu
CHz/Z60VEJIMOPaRscx4V3dlALZygAeaTFelIEfxP8Cb4vS4LuyFAwY+SQZUrT8Y
HU2jXKPSA/rTRXuCK9sQL5KmWqsGvSkmKmSpa6BQ5lcXKW+icmJjk2iCorXQV/xI
S5nC6JAF4fEo1MF2u/n3cnJQsE8RrmH3DAjbEVI+DUFQvunnIGNEWgrSlyuhgPKQ
rjCLtMgSRfpbwdxPh4HMNMlV5FLePNw7AJgi2WT0pjGbhFSrC38tgAs6dAA+D7fL
GFqDp8SVD2uuqaQhs3XiJCXCtPMuzoBtPEGjmQzNlNoCOeB+1QzW/YlgH58Wefdi
Vf39y28RBx/oG7KoTzWKcsIC8Q7a6x8tPplUKG7zxeQvPmNyZe5i6vrEnKkyNoO/
YS//0tmHNO384BeMksM6o7nc1i168pNWHWQPhfqxwH77Q8FTSGXjsNIQA2o+FaHn
INrzTirwacXSzTwfiZC0lQSgdLB56SMJ5PebfsLicMcfQz+TCSuyOngVefl7x0+O
PsvbIQdJDL7NS4yWCy7dfP70tg+3MHP6xJFnaKus6Iwx0gZU1IJoqTPAqyjgaMpS
eIPVwFLUT3TiLmuB8lj/wI+9ZB0zGon9/B1kVcOaAYaY+nbp745Ei/0aNqV5tBIk
op03AhDjppNWgU7baZX4kuF9C8sApdXM+Kh4PeMruIgv/moy80iBHpOD26tUbVCw
xmggDhE8lXJqRxTt8ai9huufISJxjQxFuCRTBVl7ws7cuFg8aNXwnAjOs4P0KYzL
jSFmiikxLf6FAk+cjffv6Qqns4ZV25ar3ReP6tDcVBkCMI2SRCWD5pWx7r8YIlSC
lokJ5ePijzCmEDT/leqE5kDrVgUOaLs3Z2TwrrfKAek5FKdg3bZCrkZfmLgzcNT4
roOISeZmVYFY0luWVpzrXFN9Q0qw3g/JdEtxvUVTPcuWi3+l/prMJZzMc5Cb8WQW
n/ElJ6yPgFik2fUQZ+/0fnhuf8NYdC00gwZr96hI0X8eUgFXH+emKozPKZ/6gWG2
MXO46FzkGEF6ltjF8EblBiRqiNBj+GKJKvKxWr4XHQjItkOxinmDUWf08gpzPIXO
BrYMCFDNvNA5HFsLusTuAx4su1TkTj59kH63FdPMWlX2kZnEpyQumM4aC8l6MYSx
v0K3Xj8GCsRaLzQUsDXRI2NK0QAdf5JPwfho5yS9QJslZvMc1rRQYJDSreWi1lst
Zpj9Vhe/XOGG/Yuy30VAUV+TnZ7UbSNSYZl+gzeFiWAYXQsh+4boRUNGXb0D2rWe
f3gtasOtrLUu8AxwdSYc/qcXnsDWRjEZamCYwdJqUPn9OuQBAXHKQaBBtwOBhEFb
blOsN4eHmecFANil+DCG+DxqDlB2XjkYXyWpA2JsISS7q9zWIGxdzK9KU6r2FneA
6SOzhDYOYSyR4LVGRMe1GgojvTQbl+pby7MVSByMiBfFHspw83b64D1/XskWXkr5
0T5q0Q6fLP7TblqFVfrF+vcRTiRgSHx4BRWDynKLHX9cYNIcj3VMnIaW6hxLL3Gm
DL/AaQr/fWtNvuJVnKQzcj1E/ahW2QDvPsTXI6lRfgaBfo83g6/BK2aTz6SFzlNa
BDEtqP8H4s1rWjFUA43MX6Q5XSBNLHG4LJNYL5dWOLlnWmfLw2k3U0RxbccaO+mI
zKTHPA0hjf1Yg3CgCB2fHeVdb30PF2Y2iUEc5Fc/f5p6px7IlzYpxbJDAv1e977Z
gWsSPYRl3fGWWNajLwMHjJ269JDq4t7y1Z8rApVDTktGYlo13HbyCXeKHoFBQ5Mj
JQLb2q4pgekm53Y5T1Uf0LjT8R1xR2fzbnSdMo5ZuSVkDXCE87rh4RSJtoxFHZ7Q
kU6pveW7tA2NaXnSDeN0qE3/7oFaiA+4E+YYJRu/Hf7x9kL4BwwJ/CdsF72ee6j3
nXJrFzFUuVNc+6SZtrVd70yjoAXl8QH7Izn37rhsVN1QiFsLjMQefXuqb+fffuZr
N8YuxV28rd1fNlb395JpqnksCdFKh6Wdd77VLbO3+fVIlS7/udcFgSRSOMoGPEs8
GdO/abKneDId8hIApliVJURCA/+fPSkGHmebYIjvLxlHwSk8sW/6hdZ7JVDRgoqq
DMFE20qFS++XdHn5RtE9CQuaIQPu+YM17lHIvIgvObVHyPF2BNZ2Or3TfGoRo3fi
3tIEcNGwXmunR8iPWJMt8ZNODAaGKYGFfEq8GloOqIF1K74Bc4XUX45lC1jClqVl
iiM8xBdNEsoArK1PfM9TmjzKIbzWFANdNRyKoBFigduf7Tn6PXe2F21/eJF7S2uu
no+Mm6C+aBYR+OUTwcUiWH00JRd2r36NQmrjatkxerpvR7ml4Ymi9F1gpA31t/gz
9Wb5f3o5rTro5cvmcsiU4eQ9HiN3kWhpc/iAR2kv23z/ppcqDuJ3adUdSM1Rq/BB
R/+SaEquCtZ3N4Hd4+TpL2t0AwliH07TZ++dybdgflM7QxvhX8SqpajNsstEEqtA
D4J3q+767siwQKdVwMLb2c6LSXzK9GhSZCpNd00rH0sMJI6B4cxSAxqovEKN3Lhg
ofCjIuiJhQKGNmDxVPzNWzGQRylieksYIPwpvYTKMr6pF6ABRlLOBLYxOThbH0oj
LC3kwaILmwJq890JjhdSjmUnZce2J2mz8j2qgxSg3ecG05TZ8uf6im5HG2nOfusP
HP3L/EWalfZYQ0DNdDRbYqFtbD2yT0ulD6FdjQWLIrYcKDJdbFP3eVdVoWHsqYXC
ozPvHcxcsMQRvGKkRu5xsvhTGsazJbgpLFXJ32jKPA+pU6hBtIyAamwV81K37WCB
Y2CoswKkpqIPgalJwsGRMwNEhYAnJBy5aB8b8jxXtqHN0OZBxnX/0gR47eDwivo/
HNdJeRZq2tA3dQFCCyG0Yo66PXuJ5UfcTtCgGcYHEDRmd2srqYwzM2a3Lwd0z0yo
6vRCr9SJk/TluTVhX/YogdwbDWzqo+0gYj4tIgQtxcpUZMzwK1N2RlXE/3K8vK0y
zewpnnQFz2S2Zn1yjv/u5MO6BTrT3ahVSQSDrx4pwudT6y5xKa3UmL2V5EzmqZbb
8g8Xes9GcqNGwcEIYP7Mp9Bb7zGOUuOAjUiCZshgoruti+FwONyU2BGMvMmvmXbo
Ti+UF2v1zLWUz4zqlw0m6oF5qnumpSVmfssnN9K2dVIA3dsPvJggxk/PPUkusZyK
MvJn2Q+oV8z+1MGC2RvgGbTWCsAzZYg6Ebezzxw/B+uUMYYHQQWk5yStyxChVqIo
NnRfzYdrh+uFvcofHnfYssUteTJ8YTKGsmmeIB+3RbosGqmpj+3ag2ye7/ifyZjg
H+N4a2hykViOvyY1rROeMdUW8vURzxf6SLUlEGz7lFtYE7NssEJ/e7/BCtJ4ii2J
mNOJJ3ythDkRlUc14uzW7NcEpHo5w+ULPian4sXI51mDMAkXdPwDt6Hf+z8dMsgd
5f6oZdHFuSB4x4QZ07UAg1TI9jMrYY5r90Tmk11Q7ck3fIT+3b+E75Zb/Z5Ny14i
yEkbtZDlGq+funOgtNXhmTh4v6SMGarmIcWplaw6hkZGl/ghELOb7NXS0k7t6Pym
9P42quH3oW7lLXqHD6Uh+8kpLWfr4px13TMppd7a00SyUkkgZc5ZJAFY0EAjupOb
ES3cpXnf3lE9t9cwEu2ZLd9+Kqn+sQA8HvQb+PImmzYfqMOsVBbzDeMC2iGsoJIn
5fyJuZ60vRmxcN7CtU7yQ1DEtaPSzLUapFQYbcQzXKUbZcNxRXyo4+713GH32Ahb
8a4nTVLJNamwFmWDVAeNZQTyyyeRdXBzhccHjeIc0Q3dr+x8vutyj5snhBRJhXck
3Zx2B7QFms9NUvLQT/oPShNwoJeii5HW11YE1ckvhkJ8VBaTdMmntwrUQxvn8Pnc
l0W1IVOltVKe0k6lexTKYUn9EBuZs1pkmy4vkl2STp0GMf4dVyQV3TWWe+/Ihh6P
pUFM+58g9HqxKVllocJGxRyeUWevar6TDMt8qg4AHAQ6lQ64LKebAYLCjv6O445G
2WXQg5psZmbtL3jNvL2O/KfDrh8wRCQhYbDYPyk13b8Bml3bCe/leGGZiVvbovDI
EKPfGUG13H8aUGhnIok/B9FLctJ5+3lMbnx9JrSDWKCnAWaYFHiRdzIuXQ3z5uc1
gxQgNWa9+x+gxBeooqDVovMTDLTKZelT5nJCrdI5ig0l9No0NuBH417zdLqVqvB9
XH3GIKyQlyJ6E5IPPx1azPX/JE5z8ILh+TDmZFw4QwrHbZ7A/PWQvO/+tBJToWJy
IDfUw2O0kBE6dQu5k3E9OeoH4Y07XOrEnIbPLIz39aPFfOVSBY22tmXw4XNpQXdQ
x1/R0Gz8mu1YiGHhrc+shczsQwU42yF3GcMTtjT//Ra1zImwKOJLTUhJYiT7mnnl
BvrxZGpsJhANjFO/G1VhYgV/gTIoVc77jTgljSFKXJPhlH5IosbrAF4NsH214PPC
yJIXEwgYn1DgK+h8TgMT2GVL7sMlh3YuitQyNVTEra7Mb7s9SH35EzMCbx+Wf76u
rEWY7/tv/xJ74KPnOT16S4VzPcms0fNrghZQc8P3xtbQo5rwdN2QjGi8c4QCR9qu
4tCZku+p6e+P8PLlTPzQxnHbKlWvRi15L8S9aJFUdry6LJGUlcboHB7whl4eCRKe
+zLNw+6kYAwBhYKf6q08QOLzkC8XulHrVdxffvB3Jg4M3jvvJdr5jTnosm6dRzo0
ZscGM2BaOT03QGBUOkvv0jtiKcRuTSmagZmWqLTZCpMEycm0rJO0vLsCupvkSEq4
bSx+zox66eLYzpB53ZdtnK4ZWc4DqZ9pLjsPzSc7RVM2ZIYhsVoR+rZTp6nYl26z
1c8dVlqqRsxknx3HQO+z5DzSsWMisbdDjPLpXxlJdm7qSqismHiIsPdaoM69Scyu
KFm9K1eMBA/5OfA0Ci5mlkFpYCj35vaUC7zRWRCfU1cbMo1N5BTqJjbG8eXBNTtS
NDdwKIRtarlR+PzmgZcscU1gdqNeTH5RCjckkNCpatQ0n/8M4Pe8Ga1d7bjnfcxr
JFNQkxKlCmJOxXUzBqj9PhYXLW1v0Mdo6wE6QRkTx9wjpg1o/TlAn2wsmvXnh+im
jmCqPJdJmv4ud643IJb867kSiKI7hE3/s5ZgWY8+6+a0DTb66teYPK8gFk81LijE
juLuyCtWF2bHs7Q5Th25u7Ibwcj0KaP4CdgUI+PKMiEttBjRHeqLGsoSt8dUAE8V
xPCrvO//sFXu25yFHx0QfsHeHmHBhc40uam0+lGlizkXXfb/vH2IhiJJGOV+rKDH
VCu1w+DZsxYlZI6GzGw80L6JNyqjfd9j/Ou088VZHiiK06FLhRx6qBf9maGJWYWF
+qhGoz3nwxj0AYw9FUHA83jmxv6OFnEGPb7vUsfNNk87V9ggyJq8GS6cvZMxYYlK
00DXzQIMSCGGQM2/0/35FYZfMppUSvfiVKdcyCX4pOIgfhqXkkbi1x4hRdQUrVSK
X2TTUBAFV1U4pG/myBQ4LdRpbkJggP/PL68XPwp/Tjar1b1Y514JX9BwiqO2nUXo
z5flt3Od8lDu/Jdvqoogz3zZpzzacf8g+BuBDMLaUnoywDuBtm+sn1FGw2s4j9uc
qzHGbkXZiWQJpd/Ez/UhZkLTOff5upAlGly3P5/UjTTSytAxCydUDnuSeT1JSkyg
/dQTBogdDS82NyADJuQBKCfAhP+Aw/YsZjpsBNd3WNfEibW+fTaoTD3yTgV5oOfp
scKJuZNlIl0TduNKjdbgPUk4lFmFXAuYfj1f+MzOrb+xoYldXr190mbgcLMhAL5d
i91KgqC6GVHPpbMx4DKE8i1e7uZz9mRvyDBz+4WePHWL3k5884QSSMgnz5WbGcAY
6Bzwo33ASiArbZWofyPRhE/oloMe0xmSokjU/iXL9ftf8YCe1E0LmhNrDVfHQ0hT
lKHoGN7m/5zJP7fCBG0on85FyEvsrVmSzsfnSQ34Jjyv0tA/zDE4qerZuSjxrexW
FjkRb0lYmAQCRXufutHBCnr3kvrLbTW/GAclfSl4Dju2/yiuR3Uk52YMYe99V79/
BwwYh4W6IvSxc9/9XLOGF42OEf4LOK4ZO/wg/OQb6PQFPbDuOb2CqHsM6K4/xOUr
GaGkTErVT0uogWJqYwrfIHf2vfvBsKBgAnhHG6Obbk4Zr3XBllj4OYWpmKmyWhq+
t6sCir5U7+wBiOJAefhvNUcsJR3NIohU6/YKxo7T4PNS1QjWi8IeSzcqXCwVzF8G
5NBEkkBPJLvU37qDyC9lsbxr3MF2R5/NL6vUOYSOIGd6ndtLYusDer0oHpO4QOYq
9RUlGVFBuSaWkkr/KMc+zIYD6YB5yKAHIR82Mq5G+gKYGeoCf61n9zuVuAsHuMp5
w32PUv7B13XpyjVmVrX6xEYLukLR/IjDYrWdYJvjtrWdxKRvbRJyQtann7FQEXbx
CR5NeWzLGtIFVNJJ8VKfL/PPLGQXLarVUkQ+L38PlDYnVLYJfv86EBwaOdD1rllU
zrbukpLpPq3naPwu8Xb/JyqB7e8xz1aogV2BZQwiABb1lh8e+xAkJeeHyWRC9MA0
HB2DBdpU4NAttUKOz0wHmEfwPjam+fxzO2la/Chaj8bsxC/BxC/73fMgx1g+o/m1
+kgF/XsqcetlIUcB2GeL+4hw/eD052NKa7UyQZO1nOJE6/KZAnDHIiaWi6RkO1vW
5hhtEZZsgvsglXBqitw2pmQuC9NxGaxTxk0S7HMIHxoeyX1WctKd3LgfkTSbqV86
WGs06sZYJDlUxDH92KcnR/gwS8ilnjvjw4235wu4e5/optPwZUOLdRXvmBMHhLSG
6VfcqPSSXymxhkoazt689RdmICjFMFbYsDWEM4ShojpY/qqEbFFhwWcpwoOBeziv
py3tcP22E7zDD0sTkXVMPKos875tp53d7KZjrI65Epv067WJQOv1m4qNm2KRO7Zd
vydeblGfhWRXdiDXgbMy9FNUhMgYdl0HMiBu0U4hbA13MZ2lVR7R5K/N/HSf8EX1
7S1sA+R84duecINRzeJLpm1cnRdrOII80ZIGabmgQRR09qPY+MPJPqY81roHhQZe
45e1iSykrqm8HLfwhRX7rjV8mqxVcu0X+NO6wiOs3Gan3os4WdVDdjsC0tKVGsfR
kSccSZHrqo0HL8VGGJ6nsssVNfvKFiGNXNnoo/uTzhYQO5cncAi9NTolE9FNLqrG
N7p6nSgPc8HyI8eVsk0sKmnDZxDsmOPEKflRaqkHjtnnwRqHUaDoTqjzp+2MrTSK
EbO5LPXe/KWF2zy8+sODJQZ+tXxLGW17FOkF+1V7DJn+UTp5MfDTAqd4tIpU0PXW
yx3OkiOxjfPBiuaqxkdmeLcrPtMSuPtTyzd26rDXLY5Toz8Tx0LwqqGr/Ot2pLf9
ExVbiKVzaSAXgj9Va4rge3OxSEM6sZGAwmGjDH7P2J0VISUgwGHafErHcyfC0u5d
ALPvxBOSV75NdV12dwWdVjBlc5XRJ+qqa6SmLKr1qPP1p6/W/uU9o7zHvSjh/ovI
ocICS9b1u+1ELsCtV52vPZqpByIwfJGY651t6ZHDmMVQlAA2y209TIF8pK9AddBT
LqVTq9Q1GNZH0ny/O9DXe374zCvirvmaJKbS5ldncs936WR3ZeYOQKP3rsbXeG2A
m2oQQ6jmc69YpCIXFCEt7B5bpQ88O66FV8WjxblUzevoL9LdFcmOPX3frGYyPwlK
euvAs3m+fbdwy+7fozJfsXNZZi7dqCqSNO74Ts0YdkLPGTvW77wG3EbSEk39dGxr
xrtlATdtojY4xHy/062b5inyD7k40unulS+cIM9i+32/wNHt3J/oIXzbm9Pd3pWh
nT0DSU8gt54QVBRGf+qLk8kXxOYqfSPJGLnJP8TQX+o6G1WM+rRAO19YBSrcidtJ
X/T12EbRJN++bMnfrI0FIIeN2triDlbCgytwIEbKUK61C7LgRMIVA58QtSsGgJ94
ifWBFaonCbG9Ed+1e8kuQE3WPe2fOfUZJGuuE9y9Sats21du3Jm0jvAtHrY/rEIW
mKaxVVarFpJACqdJbTmJS+g51LrL8T5Fg0KwQl5rH9ViiYEh7ayE/8HLVSmhBQiE
UkWqcsYkQjmaniM/k7ikxZo6G6eyka0zyomVQ36DRCU9ULjLUnDx/ByESoAwAEUw
M+d63bHWSH0oQ8v3siqm71YsXWPRGSE7SCI0sSco0ia1BYF0oTRiLbrkkHfvDMRi
sf5Pf4ahmHJOAOG+Ec/22earmc7Z5zu68N7JHmDfH16GUnqui826zqkqZjP2EVWR
Ha1ZxyBGSlvbss7fFr5vSMpBwfyc+iALASWzUETJATexURlJH9cooKXcLngLIPIu
F/so9JIivBKhd58LZ1vsosHQv4D0cz0IkPHta6nqXTD+unu+4BmxyTvl9jAVQDPI
FyeeNgHRHrg/Rj2zMO9GN9ulKiEvES8KiKfHXvpxPfOrncblry0GnpgO/aEY1qxp
P48fzsnP3Qw+B6CQI8zbmKUSsxePe89fFMJeo8JhRuWhke1wJtYc4GUlh1ZY8Zh3
loe9eTfYQl4XhFxQqOEnSF4Xqtl3b4euNmJikQLXgDfdW58/n+yD6nP2gSwgqep3
OF0oHcMcw+yMNHrWJZ+O2wDEGY2dSMQE5bbDv7+puT8bcplf2Ek9v3s/wU1Z5oXX
dXW6Kd7DVHp0V7xoadalYoH5yzrQfi3mJwpr3zGrPbS3xWn3Azpav1xjTEULVGzl
rLzv6gTfASrTXVtUVsMehD4tX+koBwonz3KTr3G/BX0LR8dKrHR2GEyZmnJcO0j5
g67lIznpq5NW13m+Rv2v7kjsiNZ3z2CFL5eEzohsTy/s4djxtntJkVxn97Ke72S0
U08R1evRwzFAxOqNBBftgfJC+YBQaHd/o96YdSfHV77qJ9r5csGwu29T3BJ8Kp2c
mjnMXp7JoJUux6A2Q1cTivsPliJMZ20NGNd7Dl1Ooxp3KUp2iZDYfcSPuSbjfAcz
gMpt/4cpTdHcL/cDkbaUb6yCpuJcc+DRyGImKukhRd6FCTV5rop0owqc8xgYEg7j
37OZ+SojWOfhYmvUjFZONtS0iwWzUx4qmwV1RRIukBzaHFPhjpeeZXDUUPwcCojH
UxLiyCAmMBnnzVCmz2pj7Jsq/Bw8w8RVL5hML0vonZmIs0T4/XbD1qLNJ8kRMqDY
QDMTephzZPgWtFuqMgX2Br+QoaslzEz77aTsdcW9X/1tEnz3t15TuvKAk2zKSmE/
U+QyXf/feQvdSrU+iP26cUemQ4azK4KGXc6Wc8tGRhwDV4i1FCgu0RWOYd52Q/Lx
JVNbldPC82lY+nzYgW3KgAOO604Woq5TTOCsE9U1Xi7T/XuaIke9+VVC4kTT1H+Y
sYEc0oRapMyWjBV10FDh90o/vNOS/hH/CW5Z2DAqGDeOyQLh9tbGC9mjHdmo+59U
K1mW5HfuqPGT4aQ2X6fFsEqfRi2iQs6IBGezZ2Jso4IOJtyua6aOr4545q0ppWEf
KUsrcpYWu/MrXGYaFg1kbWxVXtmp9O5p7ZzbleqQPQ3DNsdLkGjLmVGL9gvpZD0x
c+Kefv6pncqFdNR7n/lLTq0BNHqtNVoGQmSaZFreNw1WzaUmBpgL+OwxqNyR4pru
38M+27dMf7/77wRDvUUXbKuCCvbWs/G2z47Al6Yu/5MdxdNSpgG0A/ljLz5BYfHa
0Ty/T7mqjNVX7e8OTWy8cVjgPBS924BKVWljp5nPJ3NGchZ+hpcDBA1XquIWGNu6
l6pyQ3Hha6k0RCPYGsFzy7SvAuzTcno7FyXlHvD8R5A1ENkfxXWk4dCMK2Ryo1Yg
60dMj/2nFRkJRYUW6za7FSyU3hfkdeU1+RDxPqR61fhkaHGf7z9pY7c/Z2MJsNRE
Vie6V7qSX3ouz1Vo0DBIuLzuwydwmXJuOq/MrO2lCCkImTrOg75QBmz6tQ6Ml1Rq
FfPE+s9Fkj+Uj28CAak4Ekv3FteTfpciqaLacrpfvNAhi7s17wQGoJVbjg8Q1bhJ
xlAWoNQ+EM7QUl0tPpD/+kJWSeIo/P/vSRA1IS4BxdqyIKUYq9g4AqIkrZV6o+Hw
jhEVREHTQE4ITg9G2WvjPrLdbqBST6vo2faqDDGWoWqmx6Dr1Pz7HZAmA9nTh2OZ
435ma+ruik17172SNDvIMm2jaft39ZSsLIcB6LBeriQVkuae5aPrjNWKHXqMdvs5
osvluwgaOSy6mFj/IVbna1WsgiP0vAKibM+F7J4NaXSGBRSQ3IPLD+A1pJnfEKd5
9vH/5PmqJo57f7ttDsBsRb5rRGZ2bQ/W54QtNyr0I19U9DsUOCTTfEprfahD9NjG
WPmFGkXzcIqyzQDgkQbodfW8kvNoS7+JGfyREs3leRUhmk3+LK6nyYvAiMFfMwIm
2y1maEWmM4lYuaum8SshfDcfP3aA5WAG92+glCf+kRrl5ybjbDsVmntWLS3EZQ6W
VCQ67pWt6W8ljHK66HFIOFL1KBPYNBuBSQb3oCK5biFx0wKdikS8vq9Mw0YPQOv5
5e5Xe2bAtVu+SWJo4ekmXQ/jbXHj6qkZmAsPSFGcDxOg76T1RdagoXRe2Ve6mCyz
+WpfYVGQeMBEGeJwGObid0hEvfKu2tm6h2fsmhbJ/28wG16EfSlEfme9pqmRxgl4
SIOK34naHgLULrIUUnl8qT51dVY3BjdlumwJoA30X4/uCQXzirNxnKlTZ27Rb/qO
qW0FGqgalGxrj1Xf0F8KJEc1vVK8xT/h7WbBXBPrU7g/BRrqhROSRZK2Q1H02di1
ZmkdRsc7piiM0BDhBARja/3Yd1UiS0DAPx/M08v8CK6jYUqQkZJwR7gtV5dA1GQ+
eAiim1/6emxab8cEKAYX029o8iKvSgWdIqp3+3cE93J/379ZpNL2PArGUe+Juaun
8SQ2O9LBFlDOcf1xJKG23Ux+XO3EPKz1F0E3UbBwvX14JuGTQdp6qlWAj1NBr1hY
yFNZRKkRPXyva8sfEs68gVHYlq3S3tEf6RdtdAOQNbeOgEXM5eV4Qg1OuZyUO6Rx
3MSzr0HYzHk5kJtGmz2i63te/i9hT41a+8B/QJZ+NuDoEcY+sSw/ufD/OLl/mMc9
MUTI4sOob0iNGfvPPGsKerF84i9swk7zAc29kITInZMXZCrPsm6b6TziN+/iN7Jm
ZlCLWdS+eCojXDppl8TGN7znsol80T2Q7lTBOwAFS6G2crvFqML6kPvkwZ7AMkpz
fvIwi/X2GWIA6ITgjvHALQBKjpxwibIIVbwJgWYv9/Gik5C0iilyvsCCgTXIaOat
0/230LMUQyMaZ/Kamz6CGx2bsQm3KBDdYcJhzMsYfOYZ4A6z/VQJekdCVhwPONXG
pwaiexgfv1A0Xa4QmPpjLeCk7QBtJkHGFL6Q6q0uyrLt4WxGKh6HdmeW3rf7P883
eHI8AA4BoP1t5IPyRXFKGRxamFwToXkwmPqyHPiuY6zd8Npneo2sIqur4lB6ePjN
NYx73qnHI+KasJOVGVsR9mmM2UWtYftmqLSVnomZkaMO/a4eUf/HNksQ4LKfi/ep
Bm2Xqy8UFQ8Yi/Xby8dyz1/qa++Jh3b8BvcrYdf3dzg3alUdpYDqmdzXkM7UXu+s
MmunUm9qKsemtT7MFaDn751Oh0VwRAGIUGUl3KWZe0uPa78H4cCBudN1y30doEdD
R9ObaVvwrah8goM9mj1TT3R9Ob3rgiht50YXVNQS8br+3HWG/fTou4XEwBrgc7HD
DB/qtP+NTVUJMb3NG5XEMGBbzr1Y2FacGvEv9U7mxkjPHcRN+WXbA1evHdCIliAC
2maKX1qusNATPXMDt9J9jRPywQ1RccL1VjPeTltsTc3HL7KsCr02Nw8M6q5RFHlG
wEJrC6DPFTIwGbQH5USWXI4adDjsxBtiBKTRas4mcM+yP4r2T45x39GqJN6RP81b
618U6sDyac3Zk5ShloMF6iHG0/1Lsg7U4yMCBAxti2Jcu3EEwybHzaAoFMW6NXCw
7onpzhlSA/LXUH9H6siWmUPHF0zkE4RSPiVeB3GdwtG+CUuDOABh05cFHwPh30wb
Azrh4Eq9XVHBqTR9Di9P+gIoZRad5/bmBJgXBOy5LMtHTfVh1pw7k2IQxWLZffgR
I/r2abmbs/JCJUyxheyQHSKoslSfGCBt59sRcYtEM27WK7ekZEOKmDKQ5aRPX+/i
vq+nVDvAHpfUAlgQi1fBacmp21s5q59YE8Sahcw0BKERlQ3x8fulOjMCrA2gqwWS
L3IYaWYW36+56BFnHMQKNRLaGErf6eRFt/kq+/tPrpYhj+FEPZG5L4xu4zgsVswm
I5weGFGEZ27Llx0xeEhPmioALg4IqvDUY/+J8g7sEg/KaEaY1aGOzp+GXxXVwU/N
BVe4haQKcGtEQTa/A0knDj9JLcDEFjEZxFIrYrnBOv/gO6ItAksCyBYed8kkd0h6
ZMSvXGGVZSkYSWfP0WrtA4+rWXenUk2HusGQ04698YYqpJnEKa76MM2wTgYgLclN
ySYTfXDhR8N6hk5QbWwVUA5CXQuVD+7/IK3X/+sOzCMCYS9dNPuzKK96njICUiqh
s3b0rReR/keDAUgOYokwoj8oaBqWAJr+xG+a60LL8q2jjk2cZzvfYe5StyzGwkx8
OMvJTXvODg8kQC9Z+VmoctWyzBn79Yn8ax1BrXxqXiVrhGcvzT6RXA+bcdPVOUWr
oMWzDhhs51xrqj/5zzyhTk6YE2tJ30Q8dIbI6WMkmCYaRLuNjy/w0Hu62fnIwhjs
NiQqxH3D/3KF28vEcQ/XK23j1yBH6IyVcqe2l+NeQKZ3JeHSYnZAuwd4ev/rT9xr
wO7pDEU2SYQPq75SXaIaJcU9SACyvln4TH6Na/20kIMSMebAEDGd2W7b/bcIu/Wp
Cw9QBEryFBZ7C/bAl52XF2ZPS7vWIQIbyRB8i9g/+70A0vKq7jUbAhARHLNT08e9
B7UuBDzSAYLn3eL5Ykt86MfojCFSiAa1hZW8Cav0m50/NEkqwjXCkEv7Hn5jEvqA
JIM7XCM8DLzHFOYiZkArDe5neFdAGTDA+Qb6bBjF43yHxr9Ts87jjROhAmCPZfRr
YwGOtdWhnvNRT24XbMeHwV0EJpRetftCX8TCkzDyiVoa02tnGHqWtGDXrtjWiLs/
eagKqF80Fxs3i+O1azuZ0dtPTuxu/fPgxw+oEjwH6Ep+JqqWUYE1b1vIiiZGG4oa
IPJA3d5WHfm+Qbvor4b0yFVFi/FEF7M9UsjzSR8rigptB2lwHFcF7pEWe2grwxPd
oob1BzTwtHXH+8JHA0clMPoUJZLUuDRbLDakoJ9mhgah9BweH6SZ+Ed16bSvL4ns
huXdvygms+asvKrP0oY/vIJFRK3E00fxRoRd6KkX7F0L3G+ms5KUXhqkvQTa9QL3
E0dWSnwrvkzzzcdVTHpbWVAfhiBc3vzp4bBgNbmYlEiubU/eTtIUEhaw1mlMSb21
R+vfbmW5LbFkhIi3xZX3ormNzF9QGKUCJY8UJa96y0end0fmByWLUYMd2KiM0QJb
CyIYzUmunfY3ehZ9Hng8pMilmRLswFf7BZVUJSydlfCHtp3fwsAe7gjsJwq2PVJM
6XyqvrpJ4dKqvA9brcitp4O/mt8PCJEeNVHY2QqAawGg2X21CAtYmVw4tNUjiHtV
V9KpQ6oV9VcVaB0rbsoP0RWRrMXTp54w5H2a9v3XmMP24A8Sv8LAllZz7L8w+J7+
n4CBZWkTRVUzwbH6lrxKaoBg/uv3/pms0k4K1CJgMo9XjeI3p+50qjsa7/D691Ay
wyjPTT2SYO0XgDT9H5YfZpr6+f9MM12uFyiG8TnhTDHV6cYLj0o1oHji/C+VEdpX
aCXUsZ8gSyjab/X+VFUMIl0aPd7X7sJkWu3KIKh4/JygFn/CgH2abqQbS5XM0h5X
6je9eQhMimwxQvWx4UC24NXbp19IhMuUvrNea+UhT2P/6kkOBmwlv5BPwxw06Yq+
AN7pYMfcfn9e6Jw/te+A4q7BNjRLD+inN7Q9KAIEWN6dtP1zpji36Ogs1aE9zTPB
YMozxuiv5bbmOSQGQX2Rt8zBKov7QDJ3Rk2bPmZxegzhJnqMm64ezxtjQR00b7Wp
aG/wDVMkyUpC+0tmSyKn4cCw2bZrkz6cQb2sSgfUAv7F16ZA+lTOqWNl6XxM5X6N
zVSz2tpEe2tauOsiP49JCfyU42sTzXbnNuTX3MJcwmweSKQuXMKluChF3guiozL8
EB25MTeoqg4KpFVM6NVrDdILJw7X385sy3uD6UoLMcYbc716vneSfhnhGl5YnOtU
HUgf5syOflfky7krD9ho2dEnDCgJTFId0SWeEyn/FF8c9w3O/TVi/0R9Aqc1BwFd
VmnyUAJ8FBtHt8hRSyNvBCigeMFhytSLFBiHeBc1w75zc+X3EeXzaH2LijeHEPyN
eJB4M06voDnPGXo7Wsq14IeZcygYPOmj6a3JGJMM1MEAZoKkjhg2WR+P9MmV5BdB
YUHmxPnpcUD/aG4Tae9jQaxUVTHNoujZjYBrQT1ow9jx/PAUBwFniQ3hNO78zbXq
uaFPDRzcY9xsAp/G2K+aYuarGvqBDygMc6Fcr1e06wJExDaMAGEEk3SVkh621LnW
Tif+FafRKDNbJxtVKqQ7KQ4nSL5h0zDT0a6azLlJrxb47XNjLbMJrGzKA2Ak2CFt
SLcPBKbMPpAAZMDq+ryXqvdy9BazuzFvTHFQ56XEt5DDowiEixNF/jJu65nSFUqW
FKAzcCJmqCkY4y69GDfFiToChw7vdNwZ3Vm8l+JRiAUzKO3eelJ6l4EjYqWUU5Ad
dsKwdA6oCJcH0ZDoGBvUCFtP2Z53f1nrn2bMQXPpR3FMR62bBjDGdogJar9CBprT
zziiwCyafJDoIIlOffUdz6ewoNXZNevr2L3DX7p+3ssAbR55p51c2bwT0LwT1+8B
c0xGPwnnqbyui+s8C/iNrQuIr4Rzvblx6wjiERbfV1blPKxv47xhTZ6SoCGSuLdf
ecDSTiGRXrVxRmXD3Y/mvOTNjLOfGOQKhNJReNCTLw/mj9s4PdPWxZpDDH1slIDt
Av4ntmdgDhqxjVkQvymyQeqKwldJNsP1oMvN4wdhy7vnwkAKzC48SsIcxcxSaA0z
pAE9JejeHke2znMOTBjDD4Axj23qLaAK6K2lalw0YLaOtXG8x9GSR+4Hc8cBSIvZ
7exEwqwR8KosVDE7TxeNV6YcOjfUI6jYQvUOlyoGSBS2kjlPiXKIZfPtXk88PmkF
Rla7w+yE3ATrMMYvtwvMsQqnaPss66iQh/od6Hh7/Fh5++gKIPFuxobe+r9Phpiz
wvMZAQKGOAlZBwz1zBuo2dX8OgwgLx6KHo5vE0NQu6jyZykDPkZ/8AQ3Dz5/JlMg
ODb2ryHywVhTCJha5VYI48UALxhFCyC+ZQpOGZHgJvHkLroK+GXLf3HO/J0KvkVJ
8FtsWKpmptv7pkKhK9xKMlIdDMC+sioFppxmsLz7Ur6QEm/vTQvzb/ne0U4YOQw2
X0fpY+meAOQ5/5xPk0au2/n4jXkY9I6v+QL6knQahRVLn5aNJuU1hcSbSO87zK7A
aR+MxGaS5B7JfxUKOJ+NQuOloT+igZCdSyHvP24XL+sW1YnEMwHLr7sZ1iZqwD1u
aes1bsnq0udGvCke/g30omz4xOrO1eIqbJqGi4dOUyShP4v0HJtaMtbE/qyltOFE
Ji1Dpw4RvJttEwqDMBkuW0HNm0mPXgz79+EgT0tZMLEj1o7/RfbWqZl+A63eVNti
IoYJq8nrCFXZErKxbKPnjyhi0oNp+aCcxIfymcsldMNPZSGGhS9MkPaBJUzQzevH
oTu4qnFpqjzFxDmay1fjHFe6DBbF7khJjXR8pW7/Flg=
`pragma protect end_protected
