// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
GaUHZphXsbc1yBNYUD+oD1eJdcJdv7NoUS6W192jzXcdlS+BR9vXYFlqqxSKYLWCmbqHKRSF+MR9
291dwMSOBKitrlNN5tpKkJ2GdUvUlP3wqrneRsZi5rqivCX2y4Knihqjxvjm5+PioIBI8KPH8Kuh
e0xt6Iyquyvr2U4RZg7OM6bNEhDcWFdbdQC7tka9BxcZQbBI9MM9gYPaW3JaSqrV6FCsGx91skzN
Xjh04pnGxRmbCRPea76I91NiUPV605r7qkd5K7vgWmxgl1PfSVeD/sL+NWZ0p7PH98Ls8/Dmz7Rf
B8Y5KVmXG+HAULIzQX+yT/FOJX3gbH31dfjRdA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
C94CLzqVDTZSsdu9L4nUqrUTfSpKUjqDziRCdI4WAFWpWa3NPaoKW1ZW6TamZxgVDZhwbTCo3ufi
dHOqMkrkvYpV1eER21d5OG1elIedNWG6hw+CNLOjFZVdbA3cOFhkfbZOf4A4evm+T2X76TqBpubU
7GK0ZCvUT9sXIbmF0K716KuYtRmuh3UM4OkWyoyQ3xHEm6FURwR9Pk/Sq+nxuow9zdAwRlvvCQ9B
WN8jOdMebolcSonYbsqfWkVDHRaIr2LTMfyJuhCplObu9+0HXLUQNKJWJzIqMQk9YqGv75/Ye+Fw
Sm9moWYw9s5UAkhNS3nVOZpXP+5wDFbbt8x1MYH+I7WxjBvVuV5UZlpheR2prIa1j3VgoGyzNMlh
n2tHG6yrntQrcIjkoTvwTZaJaOrIHwLGM1QJV2JwIPXOIJ/anZamikU2rRdHk2BbC/oIZItYJS+0
H2SrkSOq7vAopNFOiFLEQzNg3441ZEJNDA9SpwTZu7RNiE0CxQJ0+uP/9zzNIBUSVlm2Z5x9Ux+C
kkTr53Kaw5n2dLWpRH0Q4dNvEn+/rOqbcKt2fUAACrOZzAfD/+kNHkOCYQFLnvj29GZWxIl4ezWX
5/N3pAkevoUiEqb+iNKx3rWl5TlWGhVZbRMfiqhRXKzop/vbO7/Ioh3hL6p3AIy0tUV/53/Tq7L2
LA6hwh1C7zn6yxSdJJkkxoNOKXBjieCjlHx39mr6nXrhSmv6zZlxQGZyvEZiJWDEe33HFNIT0RBw
RNDYejNS4kls3tRYVDNATDGV5glu3BF9D6ZG/+ePrhgBek0juENRDTZzuA2KkScieHqIGe+Q25RS
0ywO1LbBnJGUy94Pw3ykQRPBTxzMYKkMk/GEzH0Y3p5rHoZPd0DWX5heITBinkvZOVBP4l6vGWcT
c0y9EcvMm/eJvNuIVqU8qEaQ8sd4cmEPk3sgM2baw3l4iofFzwI9js1IYGwp+nUDvGhwFRmabNuz
lNzVXn/GGWmUCnAlXGWgzlAVqMnsdCHu5cyWwYdx8oT9riGql9IX350sedkv8FB9bcsxuNMpP6uT
/hJszIbCdgvtJuNyZXVQwiuiKTRt0MHxGq0qpp7qFg5no4r8357fNb1aQE0j4RHTJlUjwWJwbFHA
1IHJArUi1Y+OSMREVoVxPxxJMdvtot03yaVZ0eyTnSpPTG7U6MDOn5Xrixml7rOlLjff9RVFwHiV
Szw0SEhWXvoR/SNatadjej6wsE09TXVrZLgbz+D0C3MAi9Z8IAFPAuQrY1zcL2iifRCJwd/cbXto
2kLlgiqbJ1P39YOFJzaEJqfb4Cnw5uVDu3kqPAURmqLvrnIBmVFoEvxtFOoTolcyPUNMSH/pExk1
Pd1SR6hmZhTZgC9veuQiTw+zEGmcPAcZyd3tpEtP1EQmcAiy7vloGrvtGqojRSXNsX1bGia852Pj
uwu/pkJ6ZB6KTKXZjhzAnJQX1cwX03hXUuWnnPDe+itNZS4FqCmdJtOwx3lK2ACTWJA8mr5qEza9
Slf8HvxP3ZgQ209JuCxEccEiyjiZu8/xyRY5i/w0IBF4V+4PtY7APFSQI5GJ4quvnBy/ay+fXu/S
uT8u2P+qSCIN10+JgLuY1QqkSY0pVdKt3wvTc6D+43vlKlhbQhsA3tT9udSg7T39jKkFXPoqgyEw
DnYI7MVSuLWqNU2J+/8OpNwa2OCzk2VqCuj7SxX719sE4xCu72+sdS4VRzYQQOSs611cJ/spHisX
1dI8f2034nkKmPQtAujmlnUI1AR4PijDIY4HaycEr5KLmV5cADPsa5ODdHixuvyV9YICz7SxYuTW
vZMOjl3p9kI/W/9icrie0pq6v4hviQp53/RE376JAqMpyrNutfqCBU8oymDplsriOG96RV9qJ85R
JtZ+Q+vK8S+NDyZ9Q2j0Wog8k6mj39e/RdmGUEJhnFwBPsoarezIQsjv93fNm1gXDar8diCcThuk
LULBni+2zWt92WDtDQsUh/WxcKnQyNh05D3yNHxSVtzQ5vpKyqW37S71OITMKqoUBHUtP3+umaN5
7wTeZ+btPmAXAO9vQSOZ9BSHrjB8bcAAdFF14LTrHerRVOTXSzCCm2C6CAItCLSJZP5UhxvSfuG6
vhj4olkGqZT4bV6FtSv4bJ/v6wQKdP/QUHEmPGejccg9cBylZmeE+bP1yZCzvnMKagd8OKAdnNH7
AoZSWpduxg64SBhssy5aQ56+zv3LQUkZq3BVkoYBPtASLjP+g5sSro2wH4MIru1yJztfUSdTy0vb
b0NORs8DOIO+ho2DyaoucWV/ASQCayNnWH5t+ZWdWriXVL2+2WQLSPsa278n8MMDJd3t0qgu7iU7
i0dowKDDdDcb1DZBlX3yTmnLeRpjTOQxYGHu72k8b6y41NSmAglN2DURbaF9FssGwOXoVxSr1gdM
qUqSA4prLvBLVhIv5MNVtn85ybjgLVY79HlRl74N8dj3jz/LO92DlDbgno5AdZr6VNuOjRm6yBca
nobwc0cel1HkC4SGxbr4ym7+haVysPClWGjHKrP5eox74mNmIguf4cbF2mclX/igl9LulwAqma1O
EEUEtY1C38tzDQ4l0ktTF4V3sgIEFB4Z5Ct28y2pmPkHI0scAXC5FnZKgbjYt5ES5ns0lXgBOTZG
0edis535cGLUxUZ/xkZQ3bdLYMdM89hmABbo9s0+fn45tqvwiMfuhb+A5/iUgpi9xtkovqWdmHgK
9N3QkllDGoBDE+0EBGSIlpRTOg+M5RdQD8RNKff6cMkNGN2yRcnzgtyjcORQuNafEIQQ1Vpgrofd
2MkWDKrBkZQDjjQD6rTwVtr5heO6YZuKK45ST7xliNeD8RBciR+umOOaay8XDOwrx0e8bnOfNpuE
fz8CiNNcvCWA/WlWW8qgvO/YZs/XO8fbku4v2T9IvY5rd66rrNYH4peyo+fLHvql+UO3TGGxgU27
YjrqGxkep0TmzejM61MBoI93y++vbr1TndHjSLi2/BUQfhwJvN3aNodCraWuNqsEAb5+oUGyGBPG
VjV3rKG1Bpi19bR+1Z03AhSiQMuzCi2BCPROnPjGPp4KVY2U9BzsVLdxecFdiuiLFtlneXt5fZ7P
UprvUpSLWEuHHzY0KEFQKwid+7K74XyGmEQF4C+ZoYx0H1dxe8f3h1ZMaH7J8zepGhPcyvZRUzIw
eGZen02SEspZRxKOySnBdkeOJjWct/ISwVuvrWb8B3YBNVvZJmCUqgbalYz3YlXp9k38VymTfPsn
jBmKGIeRQ7CQ9LW23rYEVdqsapOUDRD0tKmH3StP23UDefEXU3kK+4cQSs7d8Do6Tc6crK0cRcpM
F0zDsBiI8m9h52oEzzSj/htli55cwARr1XP8g/Oy4A5SMPRpL7vCePO/q1zjTibsDRZCkkZ2LLmt
Mf+gSm2CLeRRSGMf+UungMVKEMj3sUWf7eA58Y5pmW0EqErVggWcyZJN+zGvrkGwZyMPc6fXBEbz
e33+qq0C1gYh/apQIrhn2M5Hkapz4HjskgL+ZBUB70DqMlc1pYNhGKx6CZuxNH68fmfIHJsHYhct
DYFxCMWHA+aVevsPZApLJavozbMFIqHdI+DOxQcAg505xxvFnpP6XxTl9FKzQuJdJ5XGEJ1q5oZh
8I6rdyMiW3bmQhkgD64FaFifdUW3Lx8Cg09qQ/Zs5bAKmxTACScJ4JCo8ZwU1b7m2nc64IsKBvHE
uIsCdYd8C/hRGgwVmh896IGkytg2N7Jk4jAXo3N1SocBqNb0pyqdTklVmtg/2FJWTR41WRvoqXur
6aLQ54lji9CUpfAcv7TwEB+PvfijV+n21yEwZ/y5kbVAgZz3U9D00vmxqkvhZkf9x8nGXqdQAa5d
GQ4CPbld7HbwZvZF4lb9JxRxwalBE4PhVEh41RTlmODdA7eY+I1bedpyN5eL5HosXjm7vx6d5XTf
A/YfpUb2ej7gxEF6NydgKGckw3jyhm1XT0zMYTFMPPO/DbSmS6r/iv3pfrIY5ImnlAYUOE1wkQIi
TcBcCmsAz0aWfF5VYE5nfMyXphwFakK5e1f3we74WwHca2hH5Bm6aPMhT98T3A6cU/OoBBHgAnFK
zix51D+hq12lHaU8zlyLGxice08+BjloT89dAe6/deakeEj6EC1znPEGm1M+2Iaiiev7Y+HY6Sf+
IrY2BANXFltF6FTgmtGMkzgt6VizLd6Vv5qvRS1KcfC8m+yhvZ9Sjbv/EGwIyYgRYPALVNGRVr6t
crOkTFIkOAkZx/v0shMbbanrKKXPidwfuj3F4ec41dtsrsCNsKYTRuvI+3tB6sRMj3+QxyOwEyD3
VgNiLg/+0dJbwMtzIvxdAhNJjH+4x4cTmiwdeChJ8UHfllg//dkuvpIuCJgBqBmNIopraGdei1qg
MODhRNkzTKxo21w9BdwztOwrus96xwwKjToHhPgwzvhZ0cQSAJb1pmvo8+pLZ6PQVcDINIojEMAv
bAr7cuTXnS8HW5YFqVA4+xWsNdmZRUkZ2vwRhpRr093/1Q6Z9QTWA9PClUC1uOwLYEvU+SwT8QcG
Fw2WKAGfOyzxfsIucT6X3wkGHcjzM8m/ZXG6NAqDrnjqXH5lEEWj6tyDLfl3VoNTLTIoPnnkSftc
BavWlzJV3hg0m+hzfemrmA4pZA0iJ0fYPWr1wDFi0y7bPJtnMQpbSCm/mYBMgk/yROlCP/2Pa8Qd
iUFknEOkEKEMrEcYoSrPG3/tqbWMHuDuj0HggfBcu30bQ7cIAXPeWd6XJfieQPhXwSLpEyH9l4j5
/Z6KXtD69aQIhnTPvVSxHO+sAhbJ4zyXvB7pGYfqgsLdOe7+UQ3QyJQbDNVQfG7idBM7juX2gLt0
T9LJTIRMHYI/h56LY1w5lgK0NYamczDg3qC8J2HcOdhDCsgLrkZo4U98Ob8wW56xuf5AbI7Lt6lS
BwPCrXoDqbNXz7Css882OV9xpXsoSrWDMV56nN2RQO4716zQ2De925xj/ox3EgRf1F3alaC/e5gU
T89cxDTpo+NWUjBsB8dwYhLULOrfvPqnXYOkjHb0HJBxOyDKNJFyxptl7utT1qRRMiD4IbHqhUjk
IZ/IqqYYDesZ75JiRw9gHPpsl8hs0imyN42lgBWaTI3e4ahVI+RMdZddX70L/ntgJ3PXfkgzaafn
RTqRmmUNaw1oLxS4A3ZLp45xfJWYi3RltPrV0o0v+4XEwdjnZHBFMLw6A2o6BIMghMIRfxe31xok
zlRvB3Y9t7VvmN2oInAmchigmIydJ/KbyoQDC5qupszub1L/jwWnS3JLRsDOU9xXh3FHiPIcAIV3
1wXzZVZMOOUp2FijnJiw6Kz/76JiAt2M/S+ctVdrIe/kmspJEtjncZXJKLx81mVQivGVm4E8Qne2
3w56/vup9Lr3X+sg0pAlctx6neT2THmmCDk7JCH2WmuXI1J+vExsfB4FTd+ENNvw14IWqq2gB594
6U5H8yLhrqU7edQ5lkkqk6SeP8kCgTNGwTLICiCSLRq6lPDXVclaCdeCL6/NT4IBDZgWI4URKW3u
0V2z94iTszSkwRZD7cq90R6nC2vmJROUdVLJ0fsP7PYMbKagFEqeYbwd/DRfYdEJo8rDV7KQXvEk
3qyrYmNK2oW4rjOgd+vYXOmjKfSzknDtmaTdtkTc0EPPTEStp2frgMIQ0i3XDmaenRlqC2uC3GFR
Cy7e1NWUYACgUeyKBEdMGmLKW1yMEY/1BF3QJ+ng0j+/eLtWNCLlDF3m9dLorqFqWxq2wR2lyBuM
q3MP+n2YldK0kvj7zVa1Sa1Ifyy29v/toBjJCj3MKHQhuz9OG4fJBbJJ8TLdjI9cU75z8R0ByHrQ
318ZQpDnEbg1w6DgSl9Rn4GiH4HKJrACjnplwTHLFGuTPlrSjvYtZvPaJ0r/huiUrmF571pYtxZF
tnSARsHQuRomhDC9L8mEWJWiEcEOMY7uVut3LLXtjuzexSg1RHdEaHuUwUzpSsD9eb3zf3MstQF8
mYishTQjscL4U4VIimhQABu/WzP4nzbH/OdEfd9pHAIttB/3RmYcW4xVJIRFIT1cnODdweOrMgv+
BL0rYWyMX24+OJB2mTUHwDdm3tGM1FfTkarzKPy+vXu8PGn57banIsETcsulbhbvIlbE9hkdmcu+
CiQv4hh1E5MekcHR/gy6qIfsCV0AmaKI7P46d1fEVoT4KrC4V8sgNdMsLQNYSzd6/IXTVwoYJA8+
svO2K/NFtYlbWFs+zvWO5A96vOmzSTXIca+zBIFkb+C4vdC4eceO4kJoH2Jk7LU5xb4Xp05jANEl
FRMnpH1gip/QOHPybx1kdJ3DdO329lkPC0QWTGFLt0RgRLZI51fH7dk8S6lI28dq4FX9t/Oda162
HLEWhVjAIQwOna38vrc2XS+PPncGTtB0wjZ90QrWXKlqn6nduqHPZ5JLkf7gG79bZaAD0qShbfNm
y7FjhvXMdn0q4S3sAyI4a0DmH5hfmQWtFQx4YrB7yx4EmPjv/Uch1V49hp8YXZGLKynOIY2CoSU8
M2LEdWMDf1msOZeoY0a/D7F00c43D3nMYIe9dsaEFggu9eydbjmNwlS9MjEe/i5YNStEcv4E0BDx
ssLrsUhhJ9FutiF0U4OmzNKCRcU/ka4lLZqtg4JDY4hCKSjiyQmxF4KRtwjfxKcnhN2dCmErA2FT
nIMbBQZMDhNaIfPg/I0GOOyJJN8Vt/mVH+hJGWC/qNo69mQ47L3t7knnWNf13Ccd0JS1CsJqLxlR
yxHCn6fpCBCNf8GBjF8t4MI2/Z6zxfGW3apkQ6eEytmAQBfKv7Y+dtpJmVjyPU+yFyGIPTDHIFEB
q/jg04wjcIJY+pPOlcrs0J+b3DUYreaosi5ckXW27VbOSjYAELdkbJNn1U/fMEfn7Jon9h8fpVYz
3zjHuh/YimjuuSWYiThJrQrYzwTHcEQkPR8F4+DscwOCg+IVnfUBflD5QD0tHJmfQevB+RCpL8sg
soFDDRpYMNSiZCnkMtz/O+Nt/OHyjqjkjlFILJcXrYrZZgEpbtCtPxfLqHCcFICfNGI3j++W8ynp
Z8xxFRLGf5hXN3546OR184azCXZYuwbTMNephUBCfbiLDBPRb/cIKrd9g5lDQa/5XhZq+GXC62Rp
eTUsgXxqCXwBvks8GZ38wylhnnkBEQ55hSGxgHIQE4WjDq0+DpW8+Ny18jCKM1pUjc84rdmpzDeP
eKeq7NvnKtAt9f4BN42XbbnkoCdVXvW7T33YPKM5DjB1bhqrp59STVeYA4Tdh0pVLWU6GqWu+Me9
8OoE0XQggwdDIHRDtOASmDtIgxI+xh6hnsCuVsQ9Lb5j/I9RmPngkydQ8ijaUYiYpfb6a4jMd8Ph
yeEPjJs7A0G4EcBYu+OvNswkFMa/KHlKlAH/WbS96F1GS3erC1Zq31e+ri6Gh4Mc7s9JSnPuqFJ0
fzBz/swiY7+8z05VSuSL0EVb0Irlt7aZcbDB3EtJ0JG3N9lRHfwMzfv1nYzOfbJn3xmGW/C1oZ7i
CFmBgTLuRp+XHCs6O9hoKxbotikY21M6r5K2n2NlSNoKUf0Xe0vpd5jQStAxB163q3L5/kjswIDj
ZE3pquWtIga0OUv/lJAavxFvykhtgMvdMhA7ch8g8XeQ0Mf3zn56G0BmsuJgD1WNXL90dVqgPb9O
D7m2qyfKYVvgpxLQD+zRKS2VIEIs4X1P6d+ikwxnuYzuv8w2mN+NDwp3yP7ypjFfbPHkqWE7C0l6
5ICEED94G5rdsxQx2zHbj3d8+NeiIiOcOpA09BE+0ssjfLjPxIB56QPJtgOq4Fdq6L2zn2LUcbyQ
mbNwR9G2LQZFFa9Wz5OKzKnKEca7IEHOLa9L1MHGig8yWGz9H4zsxKThYmyVCVRbZpMG5IvDxvPU
U81UALSN0xnaPfZhL5iF7YqyJtvVPs2RXRmzVrx+XVlnolpcWSvmMZNnWXU2TQGTUnj2lz+m9KmG
2xYqyTUMkmDApbwy15DtQsBf7zBpK+bVFyHM0KGvQaDYVjQ1htmlnt0lZGn1kt5p8WVCL9tfCCnJ
bivLkotFHfovc2hwcim19UAJRBtxk6qH5uCoQpt7D0VXWbf91fwqxmcmv8q/BzIPBYIfR1Iro0NE
SBHBh/WhEU2ACLBdvwW+B8ArEMvL7K9CBqLnf/q8hGAXY7H1nbQhj8I0FgmXgMucDTATr6/j1DVU
sPljs+XsvhSNENG8/IUc+xUZTvbi/SR9x+pUdhPL5zvAbCyutNjpQAb/WXY1YqXgrQg7CBSi90lK
M4mb/eZFtqSWeBuXV4EUfpQTtaVy/lauUGUTg05Kdh5x/Tpzl5BrHDRF7NdqHpWzFOQOnnmoP1ZR
G4SQyV9/1AVzZPBkyuGMawawToUVoRKotyCpP4yRNZkieZRfqnK8Bfj71e0CjcwUCjHgNdMpapx3
0aZpdoKe9U3xOqpHuLehvqR+tSXZ4rTM7MxJNyOzP66NNTEErKOB+SdQLAGFbIk3kkGgII+jPxEY
PsAHKtOJmdK9fRzIgS3uT68qZ8QD8JTh06Xk6aRtkoS42atF43JH/LV1nk9PjnppoZFwhoAi/XrD
BEr/Uw6VF0Lriv/3WubVvpBeVheFeZL0VIBPVAhVvV1JGnGzw+m/qx9/AjLB1uPjafyXAjJb1vM7
8ZUeWTVxijPl0S3WGzvwDWd+gGeD8+ZUHL07I7dAF7WIG1KDJHvAl2vDZ5+sYI37GY6d1elK/JS7
87ReSPy0k+O7tKDber0Vl3mBcPyX1poXrVGtiGPQqPXtx/zUpbXsQi8ONkFKGiMgb4vjMCfACMs4
U41qPWu1FO/sJT2talGuZAXn4j1j2ugbzFR6dIvsSfEee7MjrxlKBWX2pHWXxfmUVcy37lBZqAcM
V+fETinlg3d9YqEjjAItY6YqWBQJA1whymZU9+5ASHO1U9WAnQJyt1yFpwFDV6ORTg1BIxzz2ZmL
k9Q7nN5/UIX786X2WazNLvDrq80G1II/VTEgfuALYzLjc8lZ1WFpuCecCaEx6Ygs6NoFFvznh1pD
1XFKq7rPqSFT29Ftzl77atdEZV7yjMkASQFIOhT7VsxvKDQGRPa4e6cxFIqZ46c0/tNy4BZC5rel
O8eo1AjDDhp3n/l0YNBSYx4k0nyFbGljffMOtiNT3ZP9gllLUfeGNLBL1PChKrTN/xX3w0Ab2U2u
9uA6bIR5FFXDEYHguzwEWonp5HNzFR1NpHhRtkgW8HgaRfeaQkfD1PDxZ53lt+FllKhSjS5VGAB5
vuXfqSa4jFClU1ynUgrqcPOkrAkWQrTV4zYGIp4UJuHVOL812qCf4Cn8zTN6vR7WCdtFWk2RiP21
4bU+Dstxy7kD50lWnPWJY7sV8+Cl1L+TwSe5V1IfBViuJyP51KqkQdHs7mV17I3TJdnA46Jvvq2B
htPoogxBq/uEWN5SLooxBToMWiLkLptrn7fbGBFW4Smm3yLHRv06v1U+o3vgGhkNACRX99iEnG0l
I/EENjAgNBcElAwoxCmAZgHDa/BZRRibgqWhMtJ/Ga5RQeEWXGp1NQG70AKz7nUsdnlCNP0+Nnbj
4xxvCsFtLyEMr0njV+ScGkwWRSoaCSI1OU7ekU4TwYPyAVGrk2QRyhPpWf/+VbyXny62dztcmU/V
3HADV6GMOp9cn0KPadO7sAbIg0VqIiRFSx9ajNmq/Vt6CGpH7b9x2Rj2/iX228j3a2mNjG1jFtMr
ARuEQ9DYBD/e8a7s9cCVPXGNQq/hao/XM10lok+JiJUoJbwspdfDqZLqHUkTTAgc7CojORiPvW51
MP5JCiQuHu9PxfaBhwyF6BVRbPmRDhYrPbN4G6kCGEMXxe94nGiLDbCkTm6zrQl0ALqhX9733pfq
ptMrrJA+aLFeKZQZ08Ol6EeJe0hu5xcL69zktqEJUGj4NRpQS60zCtPs+zrjQL00vvINxAO+/YI2
YlXTQvX8pOVvtg+Ks/qOFBxT0ZA0ciabbzmAhgVV/AgT6nkNrnmDnZtL/qJ2cAdPQiJQnVeLzsUM
E2noZEto0ancTxtFDG8GPQN9sqfcPii1xkc/uxz12yLveL2M6LnTLeZxdGHnXc9SATuw5w5qX5VE
xGm9i1x4989hWsl5OM5Kvq7c1n3k1YziWNH0J0YR9gNKRG0KkLHq/rUzKxDUDDwJPDK/Ce6+ejl6
ji77xyxnf4pE8W5AAkplwBSyvUOSl0gfCIJ9CxOKvM9xTGBmZtUeeOUdTSp+BA9ShAhMgXl2CnI7
dcoXWOzu3APqa2XyHZ0yCD0qg5PoPt+lHk7ddcvCiWmmKOSQyD+TYTzG2i5taYG6SQeGlKykqLRT
4GLPwOKd2ZxQu7pQ8wVAWxEGFoDH8YmZgQW1DwrH0hSrzyW7xxcZ9To2nxhYOtsHNXO616Gy6a7j
11b4Nmx27nq1GI+oSiHULaPpaEAdsgk8xaV9Z341wMAn805D3kDzR9nG/fDQkQu2r5dq0ZXkDzQR
nfteHKeWr0pFbkxXDmblUcSBOxzm5oW2iggjqSQR0juYJDkRIWIyriLK66ZIJgi5cCrj7zDdP051
Fa6IbUniLk+L4LeUnll47Tc87FjkCSvdTJh+vHCJZU63zyf+TkEgIKSpqbg4KJB0/Lf35vP6ByOB
pPh0a/+VpXV/pfZ3sQ63vWKLU6TAXBXQq+kCONmqsy9S7KrbOyJgmCGHgRKCoaEBABCR2324GRpr
xZGP9E0bkMB0b0w/+JJ31AUfDDl8U8QlCB8gUr4YnPv6fUE8T4VSG/K8P+a68zOuQ2bNZ7B4bZHw
R37QLEjpC1BH0TojklA1XGDtO0t0zURka58s8ShYH9krf03wjnr6YwmQ52SeHSuOBFB61aBNO6Xd
SDI+Uhjb5LhDoSqtPo0MxbA9vQPWD2Onb47oNZ90kJ7Wu63UI6KIVccTeyY9TFij3M7ncGLfHcb0
sqfZChmMxUkU2MZJybUvc40LZ4PZIkIHXLK8twPIzlBPC+kEwMVmh7/G9f0QKUvyHD76/50VVBG/
vym4k4Y8y06LJz+S0gbPdCbCgtUUyfTF+LegwbfG/62jDHsNy7iO53mbxt8LHA+67OLUOoMM3gO3
gJFL6SyAHj+gkhm02eDWSvmublTdrFJb97uQ5V8dApF0vaiD62X9oxJVQ2bBj06KZgNboupNRsaI
dKDxZMXgKkNyl25Rz3a5897RBZQQRR0VLrkDUABtrW6QC/RIfN6G1Y4otBmoJhfprKxD567e3JXf
WhN39uPm8bxDoVHPJRkIMwwj/7Gt+3AQlEkDmb8aA5CRROLPcnbMRHJjCi+Od6g+7N4ydc4umSWA
UI+YqTyfrApvzwTaNL6hZerdm31vQk2LJ+g9H4rWZK1+bY3NxIDcteHOo6USfpT9vFMovrv6xjL9
oY3kWzs3hA3NgqHyhzUeDpJugyMCvv4OyNfJdk2tPBlI7mLdTiFJVrVOY93KHy85lsWPwfmyvIYS
HfgE0KKxlkfaOjGvthj+lI/spfARPvsBQxSxvX4XTKajLI+Ix4GK5uZxqkpSiOzN0/Kntz7dzf4T
QmQ4+kRr+59JV6RTRC8mBR170yAJff+yRqUb9wDR2siYOHEBwuAFCHSNJArpn6TNud0DXjCtdF67
L5YYj4BaccUGjx6jTFiucKCb45kCSmxwttiAswDcECSOwQZAiyE5XNBntZ81p1hNTqnl0C0fhc/m
gAzxM2nGMRC71hOr07oxVM58sYixaOMOfKny3gflaR266jcG/HH+1WoLGoW8zrMtqSJ2Y4rupd8p
gpErWF7AQavdU2xRdPmgufrYmpCQRgLHm33Y1jg2bLcjBbVvvaCDi77uZ2E13ouPcVu8gZ6llbt1
L6wb33fzNiq1quS+W5Sg+jrO2HKuLHBxV3X5QjKdwmPI4+sLDo+hIrsTsVVUrMk536tTZ1dVrgv9
54/KOyvUtSfUxojxew3jWoHrr310LHc6LqzMB6L9r6Z78noRsONpChptZi20nxzAtGLJmfYkXdCh
8iwwtgsidxlRep6VDt1S16DpS95myREt+eYf93KBlQr/m+cq7lL0ivJ0SsiWOH+5ODGkgoV19gzV
k0Hn+0Al6ufgzSFHUaEjUhdR2lJ+OqdYDczMs/k9HisgdDdYQZk8pLr7wZLmcyYLXnwyR5v79FcX
2JUOe8H/e/pVJ0l7r8rZRhLmeh3XjhfrqiOKTn5U/IpJ4KoPc0Lk8Rgf2oJ1c23hlAJxFNvdlMlL
Ay5/NauHe1og1DW+evA1kAQ79Es4nD8vb79ks3Hqof/HtzgH/MtTAWVHyfUerMz+izq6ZOfNPF5C
Pbww00LpGQWzortPlnLgpPeJCfmxl6FkBEXhGzhGtys6drOYDUNUG0moB6VetukP+v9dIy6wJm09
lckAhENpz2OT5JVuhloSFgjMenyk9NZEgPZzfT1SFFkb7lY41z5WAtM8yx/okTt7qSR388z5iINF
x5khqfoNb8djHhDLBLbOPlO7SOjq7aLtPHVbKoeTZwAb2nI1TtQ+SqFTxq6oi3VuSkOrw8qIGBIp
ilWihSlpcxK+tMmGQhuprHYA3/jhDp62EcZhEZNt63YgTrrQBDpxbKXRcKo1awP9HRKtdHVCKxbb
1sVnLoVztQJIAmWeoEwMycMJxbqX8D+bm+0ecVfKl1UEvjGNWfBkwKm37rhsHqq65j2meyNR1uLO
Drx8h7AaLqf30XcpelIVjgB9VQk/C6CZy/d6rbDdcFGSzdZ/qW49FVXFVO0yGbz6s7rvE59uNjl4
Urec6ReUHhtETRWwQ9OTQ2lNMx0E+tNzt063SX7GbuDbmGS3/FlAJsecTwj4D/ncsf9ZDtWnHCqf
BrqPoKlBEqYuNjnFn6h9idKP7nhcf8lU2TSTkRLKX7YZDLd3IJBEiKzvp8qW+obSuzungz+b2J5a
D6LYVQkD5BcWO3fTMwyqY8P/qATzv8AYYFjwNSOYn32qopS39XsbNi+aJR0GB/hpJ//o9MfTvVlR
OWjCl47Y1EqbzR0hUOJ0FIeHJW0LU7O+kVud/gTd7aGSyeMAr+H0mcnJQMNjLeWJ9Vf8FlLxsQYV
xtfM8XMVlc4zDvLFFl9cYHD8y4V32PjMcEqXTUBJf/QqN5fYN19U7K6pCScnquIAx8QT2j0NJO1q
sl3Is15qOOPttuk0/UAWXllps7I8VRHUjm/eCEopHrO00LbDSU4+d3HaOIRTiatYKf1I+d+WInRC
UNJJtd9ycphikVCPUJESwrXeiBA2oSb39q9xzbqrO8VA5hhJK/zOIfHG2Octo0KwzRe9rAYEr5/h
IaBfN6okSfKAkW2pCXEnxbLhNHPxR7nq20k35Wm9qNg/AttDhYPAhFnz/0KnnvPbrf7haiSmWD57
rvi62EASRjprI3y+c+cRgjdb4W+fyXAQ0IKbccCGP1biTTCrz/LBSb4E7KGvnV2Vib6uRqLP4Hi6
TtuMwLWqNIqDdnyEU9oF/AdXkdGnNSJhaeUAmiwyPxmhLy+AV+A0iMvQOJTkGUaTo8RP63lQ6Q1t
fHs56tdr61c4etXu/k4lhdYd8G1+zb9ieZOW5RQpX/w78++41pE+pB1PK9TM7WbS518zBt7xLYyV
Hy/riyjf66Vb/0la+JpzkDJyxfbd8vz67h65hhFKXanpZ4AroBlVOWoNZhat1bCA5c5gDzwLkTdC
7BbOCbYdU43o0A+N3nTr0W22xH1PrmfY7DR/0lhQtU3Tzmz1bOtZ91yYNUlEmLXA4KqHb8EaCW8m
H69cRj+hVgJGCdfq6hHJi3o+rK40jsWpt9sIxkTOGme1vbiwsonjp8zhwW96G/HJDTFBvZGz8+xK
B3Rhbp4kdoco0Ul3cj6g38k3mduQwBFd6aeNLndFZ75WSv7gfzzpcPQMHjGVciY5rrHPHKyvnpRo
2CMo8rmMt07uWtMukbZ04QUFKpbjo0Q3cmrqS1ul5Y2khF+luqSVwwuFpJkBDTYZqo6QG6xNd8D8
4iAJQrtzV9z/vgefIvCUYLrGeRvKkDvG5dn0U4X8CDx94w7HY1fxLlnhNbKUzdjY6q9bD2rhwhzB
9XLsy9e04O1p0OBPSlfIk1ghORNmnMGDr5gkVUl1kg6RXUUz1Qm0TQxI6bLcFVUWxr0qS9YLntbd
d/7rpdWhJFJFpakPURbJkK/1uDujJy45dsfMMXOwWI0y0hd2C47AoHG/7BBtoChG7xPfuLOrjX1/
mfqnPsw/eoycXF/ry+zTZpn2SR2zvgRgO53NPQG01wTGSV4XyLnedR/iqYdOpVN8f3nhNGAVWk63
v4JtybIKMdd6IYA2WmLaQ7oHdKwtSn4xEQZ39qaPVaK3xpBZ2LWRb5EFbq//+/bVeUHLnxkbPENp
tGena9QBex48Jgf9kNMdIQQjkld2rJeSng5bYUjQIEHm0wpIlf/O4KwNzlp9S2GXt7ozBkHza4CP
fjpLb+72hYo2DKZ+xqBBPoAzXltKtiNxCGgGqtcTcCMEyoGD1n4LpBSUZPuR7V0a8eT96RlR8RYL
z5eVNdc3NAz4ModbvDPEifyO248x4+yWtQlUt0IzpgpfLuvXW82JNHhx2o7V95qC7zF5t/pD8LQB
TJnd9kavDhZI84mQvP31pNkpDSPoDshf7mNeTpD9sT+5ecXfnBWBdYmcbV6YyFXfwPA/0DCmA6Ej
Zp1aPNkNrryUl84Uk+lw8Vf+HkoZSj0U99xqW0O9ejoID+ei/Ns5LWqBMdS6cN+BwzHfeGBFvlrk
TC6rXSwVn2HDxKPMAUmUaZikewss6HgltNM79UfZE63Q3v28ZwF/3IceV/lK2hPxrMpKjY5+k8Pv
ffJpa1MpQ+zWu1lE1d5cGbW9kQLqhLJS/taHY7bFzdkraU0TaP+7PWqdWW7q/cEJPKb2PSzzd5RX
BZiXhDTfEzSDWsdaw6nz5VDntXS/i4n4IVCBlYreUi0S1X4wdMDCaMexU38dzccmsRFKfP3RAupc
tq/AphAnNrdiric45eQaUjR56leEPkan+YiRjftVIKQmB4QITLkrGC6dgn/NrzylIKJZjYVQL/Bg
SrMcRp3XxZBueISf6O/z12CGOorpYf2pGfcmWc3KTiRqSbpuNvv2BCbwR+l4O6f2iYEhzf9iE/MP
fBTGnUxbO7jgXl5QG647xLQ6JyHYa7o1evQWhxghAfUg9oOL2Zs0M57J4EsN6Tl7RzYWDNCAupWE
vKmcVA+DOR1bpThHeOk2JQmD2/DbFvsp/ZYkYDtHULH5FpipV5dycNJ/j+Gj4mmPD572baoVSsvM
Rm/D1zyNFaFrPBY2qC/vE9s77gQg6su9z9UDp2AdlzZw08MFNvs+x1ZCQxEIcukQVQtfPLgcdoBU
zqp+OnUgfmEtSwFWSMjj7CEv48H9s3Qv+9nCo2kDdf8v1MoXvPpCX+BQBsdJiGvgAofbfogc0r9Q
t+fPR/7hjy5KswucTCX0yZHDhOjiLRcEuHfZ7VJqtzxolIVmh4OOp/DIxy1GWDVGTXAA0alcOUkN
u8f6HbJyFKkvDBGuAn3bdIAD/mpUMpy/cFmaqKzMKnwkWMd8bYguaHbVGGsaj/SQ6Z0RV1EuCs/c
Zu+I6n5zyUK3Gwp1hmrJeQ3t2jafuWQUlYVF/ZG8gptZ94ssy1SX8/nKGL1lPjYSRuNg7P5/06kP
/x5hCjNP+awvbjjhFrTn4Yx5wwabB72WEIq1sI2kzdHLNes4pqL/2v4taobN6+inSmr4pa18E8LV
zxH58WxK5gxmCUdEvsHygWYsjcuZvBYFVYz8wTCJiAZo+9geHDoqNdjPZPN7BuUmP2tsD23wMbUU
lnfsHPIJYtR8SEcCHZvRKl+TghXLb5HaeL+B9vLqHAw+RtD8Lqwgwb0cAQX1cvzu6/MVL1FnpydA
TacFMec0tVXekv0QmT51EPX024F4ERvFu3KAx5B1fQN+LPYgK6KNWkQOo/VVpbuUVY2vKBYz0LLc
bKdENID1Wb1oFcLga8cuGrHY2a7d+3kqetrhYxzVtc77Mqa9Rvj5pCnUZCTiDdL8r7vCIgwdJPy0
8yb1N3VZ0Rfh5Ev1d+PhczI7q/dRpjwRT/i+vW5gq0sNHoT3KjhD9TlBrwoanDfu8SthyxGA35Hi
qgLyNN8SkqepHlTKtZ4Z9FJ4BxCGr/8gVK3qkoAzfxZeWxJhTo3W8uJk/dUywIPPqnIQKO28lxFb
e1+kcib/xB6/6dFvj0p4PsmsdpQIz2i/LAl8VCAnRL1mdTfjuzaPhd8WyE9nAML2UnZ6/oaEDwBu
ke55qIrSDUOa7IiP8kc1upALCWeeXq5oib8CzV3Dd3SKbOqTeRn8g/8qj1oEFlqc8j3Kuwat+SXY
ZCC8cXTEBfaxBILwxubjEwc+PnzzykE5D731pGxc6oACEAGGAHex8Qk0sOqf+h6hwAoDup8WfWLh
EhIodyrBtpEjpkdI7r+ujtC+mTOoIcRTPZdJ63EvsXGrLCEy+8PBm8oR9yGhRpyO0L56IkdyD3bm
mW1BWCLwxkaAkiAp2ZJUsVLd9dnHy7OnpEl/gfzEJsRdRs9kT76Qv8vAbORTyMXGB5SbH2+VVHmQ
BmvWX3/2I+21inXVxjHLK2w8knNG9SJN8U1txbb4JrXsDNGeDtrEOhGYJUf1ZK5k9rkZc47ixjti
scNWL0sNUewZURaLZScD4849Ct0uBZu6iI5Jxcn4twjUxV9U4uals2AMTCkMO2FfTg7K1hgciJEe
rKz7DIsYtk+PMKJPhZN/0W9BflMAXRWMF6c6RZr6+PBheU/pjSO4bLcwdfMNxHqNBlHw8ikMGswT
uox6nyidvSVRXe32fncdQpETagssbhax84kymMDzm/K8AG9G6GHFvTai07mDik+gTPJaXF08Rnxv
D+WYkXtJgT6OYNya2QksDalrWHjmH9yZ/SXXaH0c4t5Ja6cC2W+vj40zB5+uwEa4S8GA4Aq4tbgW
Xk3fIwujbUAiMP6z7zh9k5HloC9U/J82b1+WzraMcwovIB/7MB3Twc+dcwLbe5UmWDwb/MC9KD6C
jRxB4cG1uT8A1Jw4iz1sBG9yCVqn6qyxXwwnMTgZPx97RK9B017fvGQLVo8W2qNwwxeYO+lJViXk
e8HZ3WSA7d3iKkiS4sKkqP9fabOT1QxAIZDrwJIphhR7+sTN/mBsLsQzu9XuWJIXn3F8jv1EKpbE
BUzOGE1beJtZZzAESWe9THWu8nFtqNEDL8Njrli6f+3hEekMU/h5G0Dd7wzYeeP6Sl6B5qCf/bD2
/Y7ZbLLmRH+cu0PA6rfSL1LDmsAzSHIpAj8U7YGciaiXULN32wctLL1/2i28f9HF/E1fcXB4B72O
lEldUAqxkWBf//RsF+J114jkogBh1bTqOR1ERmW5PRXR+usToJYKWL19WaPeqWL5SH7XbXHz7S+R
9KBWj+U+8N5jfccEq0Ea6mj47mqYIjuAXkerKUDXNcjnBcWZi6A1Rmqy/tMPHD4wqLLfG6nKBa0Q
lFtufl7eeVadmrPLUTRuIvJmCN8CzzR1afPb60nZEUA9/gropvyyuqrBidyUpfZe0Zv++9U4gOte
lDLnnf5b2qrJou0kR+08m1ABGbJdO/8qqNUp4IvAvDsnw59C7zr10pcus/HUCLxxpJeQOvtm+DHr
OcVYTkquS05Smssr3d0q41bCu0Xt5BxVCquyfFOT4Aqt37WCTB2rHBzpFm/+AOcKpJCx2YRPrIqX
wYKia0UtKfwFeMURpPp7r5IvtOT5Sziixv078nJ8zStFEiTVeBw9IgLv/JHnlZTPd5WsmoyGqkmc
9FUVU3vrXar1N+dzsHi2omxnk7lPPEfkVvbr2F9KzDKx713SbGjhTgmG3rRvqBCYECFi/r5cwLHs
GOjkqCykyZaGjBgF8oQ+yGnkHnby/S8Ngq/98NFrHTwYU1ynCGVmOn/sg5PMuxtmUWLMo/jNpcCH
eoMBBHzCRWwJm+uXfmw5aI86/YsZOlh3ma+z2rHr/ScMoowKPKmU/hr/TM2U81AZfgRRm1dp/WHD
g42QKqqLF3lmyuwIv1Q1tsVAxRjLSUVuTrsqF6jlG4RfhaNC/Bzt9ncop96RtInv4Ni3uYPTylck
KMEI/gxWjeB0qcSOV97N2yUs4/zzptsB0q4jzyewW/YXSt85jApAUqMrOZlwq156aCSITeEQ3SBJ
vbUzqHb/BMj4M4sUlEEXLdUV6xOdEyBSqAMEAt/DK+B/JDDl+F4Ai37kds0/d32sKFyV9jNkh6x/
F5lyeqhz2fFB+Df/P3A2MrKruGxqGDKs18DCaAS05qleN/Xe9oVy3mJfWCioOYETpzcYVhu8TDNK
1WEM1cdY+INi/i203pVaV+aEMn6G/oN47jHLLk39mOEFDY8D7II1+cg+RpV5cEkAY8AcfeTsCqPL
S0pNihsAJ8VgxiAcD1I6nWxFuFeFeddROlX7PgdMG6g9WsOLHMRzZKOVQ8iburrSTLVYphni6866
y8YxONSAATQs7zaiAkdmzZRFzkxcabMqaUpDGlXtlrsvUjad6wUKlBKU2q+fY6Cc6VtO+4zKn5fl
OOvekZmg5kqQfJ5HD3wSFRGQBqXMJE+fWDlEQYiOYsJEQeMWXuRblWjKzwBlAgNufLFUfivwqVNq
vY8HLllR6+g/BymXNY0aZoHRlcvUi/kowUHb6y6Iiy2qV1LzJzvMxtxbQYIbTKx/bLzstbIAFX0N
6plLxI4aPwke2AiFNfDvc3XyvoEoyCzZj8dGAP3XHHl3Fod/2ElGjditdYLGd0U7jitt7i/3tk1j
ZXcSLRg1BX9/hH9ErpGiXC8qAGasZuIF7331WsMd2P7GtJAqaj45CJJGF8Rzz8R3Z8bycPBG21uF
VjI+tYtNwUDnIkFEvxOR1lJUobaDppqSDHlAX499n0JILzGd/+vljWqcj1bC0g1fYMcbalaBpXSn
FJANu+s1vuTTKTdCZ6+eo+rrAMuNJwYyjI3wVvU8eJUrevHN8921lrvMN7B3QSC+y38aVU54M3O3
ifounool0xogU1cmCsuk26UizSkjiK/h3wQwIIXNdUAZnzbHwIICHDjBANVN/KNUd0opyrzNorgN
a3+Ln40OQ9t/aQ8buqsx9hRIogVkUMnv6W2Q8WDzEq9fTlk0fD+5h7XpvJb71nR4vtYVPCPMjnZB
nPQj6OoSPHYDNphnL06ty39zIi/FHjPw+tW8Ehu6DZTMlaefTBC6zBcUSMj9ySsIARuHV3uo8Xtc
LzC661Rl0+P1VLdNhrbyOa34S8IOoVFgzewW8vG2Wb2LmraFh5GLtwbB1cz8yNnbQQW/qPYT+OI9
ExaFZH4wT7GDkB2I4xAnlmNLQeaXZzjFVEj+yPeBul1nx6uhIyU+wBVH+AJJm1isF8JWT+ij8YH2
U2ChFEFB8zA/QqPg7q3ca46IgFNceIvGIPpcWUm0a2aOFmnbep4YLHLjRt8II3olGBxOvwiXOT1V
H65HXaTKofKLoNMQa0+khaMiIQ+XrhChfc3BkPsRIccE9EcmLep95890LneMsWLNDR50byREOdGL
ieSfmJ9b7JQVXgIYWYhjZbK8CM/YZs2kyEHTzfPybf2WJN247ert0BtqrxzVDWYqYvk7q8E8/FHe
Ocxew+inAi7hjuqi7+GeMEEm3soP6VBbhmgMo4kb3R2TTr8bxxF6M3KTcVwAFyDjfKZw9zMdR+hC
xji24YzZ9s6DLPDgL59UtZtq5wD6y1GlJg8zuqNp42zkXHhjz/y22mP7CiGRL8AQ5O6HzJ80iA5O
y+TNwESJzMQFFt9rH0XmjesD6jQ2n9JO3AZEmANcGtsiUlxnmViEeuSGaXP3KZuhtjIQeltNWgRc
JFYZiN9znS6ixAWgvfMI8NAYW7KXsDchJcRCIFfHnXude5rK1H865KZUlbla1bzg5RbqA/T1EC/Z
vBRThhv+LeNRQ7xFiHVK//b17nFMaeCJxbvkE07odKsPaRpFQA7IeEMj7WUidJxI72Mnwy8wsNx9
IH7ZqEppUyoE1lcfaj1hlHD1u+DvDy15r8cAHZck987G1ECnMLSivsrcdrz0RX5oDqh9NELGFtpw
E7USolwKffEazpDxvZLQRX/sPly4NrJ9SVevp1tWUVyu1BYRN7KnM32WpcVKbsYCQlkAUYvp7Bqy
nK1AUv1VM0O42oXTSTcYRp6Wut5Hiu3Enzw0CSyq/Al/o1IT62dxsIJ/tF+N10Ay8WnjodoZ9N+P
MZ8Hsm3R6RlUahvydvDQtDaiT59QUTTiTzhIEm2V2SgH4nKMIRgpzPyWIbZhAgIewfWaIOcGk8uS
Mo4qYJ9m6akr7U5OdGEFcCY0+9Vtdo5ELDcZhYaROFpBcSaaCeYacwpEa+eZxHllbkWRKGwn6nl3
m0h3eXTSnEMnp8cLPQz8zYY7UBgY7WMLZObLlv8Qcwvn7aCL5YX97UEPw7YKdAQrYpp7Gm8erwhf
23gt14VbwJ0lGGLL1WUHUu5QugAvloHBBCdPCfKeKreA2Pg+oHnf6SXppAjZTgm54sC4/ktTCaao
5YFQnD/EG0CSMsSwcKVI+n/s15HJistyh+L842g3rugHdsQLSh/PJ6ioNBPW2n2+ezCuwK8fXNtJ
j9TKsqKVYjZCKvAF0cCvkPazTqkI76keMWm91vUXe83uES4Z78ih+qnUpTXXcONK6kJDYHEAqPak
8dnZUW8AkacU2jpFfqSOblGKVg159Wd0g3VK8mceHAO1jPVJQoQKb1HzXp/N6nrbTkONHeHOq4PM
g6nv1DlYCiVf2CYJefBbft/Ijx0+TGwDu7uTgqp+DehrGBensCNaEukjVM6DseYFM86W5L54CC14
n3ebiN3FQ4Tl5wv1aXV6ZeeHA4PiGFAGEDpiIIYXAqwB7yRAiCdBeZ+oG//Wvmqtsq8WjnGs6k7d
AucndXCMMggelu54mkBjabAzqhx9EBlEadLQ4I/kJL7/+1W7Du9b1d3FaXnuJL/ffO6aaMsNBK/D
GL64l03HCPavbOap9Z6XL0LbTiYTGXYk9/lJdrevqCTXCtjODPKi5EAIEoxXY0kh/6Lz2xKVDEQN
AlLvSEFETrnJYusOqQl2u/22o2sFPbaZi7PdGQD+SUbRCYF2pR2TI8eFvaMn8yr5QngjgtUBaPfl
kMqUpbuZJcSSkWKwoAiarnOVpPscLyimjCUhH/YcKlEhZLyYFXF4abfCiJSu6q0okCZ+zIVUhop2
zw4DgyO4J7FsPmu7LEwaDjYydkTSgFssxhVTsUp2eKsGibnmMLg7KrLOQN63P3EyPskvcAyzrsro
ItVHPhZEWlne8Wr8rMhZi+/WpqFQHx49AgekVOalPHJoJoNtsk0aIVJOctuBcMPVr6JHpv9h5rHm
lvTrpmwjeCwaJ86EDTJNPaDFG/kLc9QCYouq3T3KvHz/gg7P/NGP9GhZ1vOuvmX2FdlajbX2q1y7
qlMk4FU3so1HgK9K3W33iXBiAa2W/3dENOIbpQZLC0YBpUPIjDKh6SsPixVJLjqAIqwtstqGzkEt
zPPtQwo43898KjdDDNFvLFm5Op8y4fOM6k7Wd2oNtKgGUgZnKsIE0j36tr5RZcQEU90gKmbCZ2Cd
rcxspEvKJDGqdSU52xfDxrNaGNTOMhVsJ0LoF0O5rYbx0Ua/xHX17ceJ8F7sL16g5lF9leUAyrK/
F99n3/lJ63UTATCkCT4dwQuVTi/LCFhjMIM57DsBjohimZcO6HPtroCCGXm4QqX1N5mjxWJ+jhhI
DFGPy9+8/grhZrTc2kWCAn4HQP7KFFGD5MpcITHNkwIKdaLkyoQr7eO8SDFvshIV1AFQmPJQoPkG
tg3E//zwkZcKnU7EKmO2hmdDkL26zapQRZec8BwkrH1nsFsaVjB7Y3z9NbQ+XZtMYplVdMjeAmJV
r7U1umHfj6w8UVLAo9zMj3mRYSn8YjZuhM5RuQuIjBUNvrxbYdI50iOt8Cn0WKMXP2/AwI/2pysF
Y7bVnN/chMeKEp3+F6CTyc9yPhpiCaDyH1577aMCZdt9e8zqUSMLmuaypy4i1zZaHzpU7DVAz0+N
armh0CvXCSbsBCdlbm7dqnv4Vkd6iytoFhQsbSmti7edNh54YmXZvhhJX6LPKN8x3BVHIEngFswS
WWVlgz9/1+vNFKLQFbveiMJ9mSH3A8KwFieznKmaSqbaK/kTf6vG23bzsoRBPfnwqUnjRy+wcuNE
ROeQwfZY6nuo/lT5k5u8wVwz+TpTmc/GQpyXDy/4QjGA0x6TsfpJhUI993xNvKcxjK5m9fIHeUed
7u8HaztTL4bEA3/ijbhobGMfKkugKJQKjlkLUhvo6qE3IkyLAtAL59Ml9QfQpNXOQGil8b7SJN5p
aeM5IBQUNfV6+NkhISKmiqHl0TwsKY7OjvlrNFsDpfnjWhfAW1fz44FeK8iP905vfYH45VsczD9W
xEi0qL8UkniqlxdhLIFWweJ3g/gXgMsi+8yeKtDdXSVzGjepzhoZHpNatDAir9EP1L+yzMSUi9kP
M9SiYWVaJ9Zf0dk7NjvMTj5O8FAkO3Hm4ToeOdP/qT3fXXtz18OQNh/+g+r+JoXVRMeb4ybetg9j
htEQ0cWo+luVcyCzvXzQfo0Vf+JCY0MkwKiKP6gZ6qOD0zOzxD78V0T4ao7JD0X1dYg68SY6BhKl
Fl0uVZlt0GmKRLB7iiXT5wnJFWmacjFDI1Ovo4BMs9tVVxoFSHLn7XOzJlYKO6Xzlsg0RrINFP6i
jEr6Cyi5bgopXLQEDlE2gWL8Jf/ViK4FAWfmNKpYSqGeG5/P3PpdXocFON1lmZhGY3+2Z5ELcNqZ
SWntUbFX4uqB7xmCUwsUDU99lp/9QRzF1A7OpLwrXo/yMrU+t+5srjBz366lvw7snDkREowYRFde
NfEDxBBKdB/wDp4S0WJH3wTbyVQb8oFHwBNc05CuSnE8CkvHhJkIvcLnmhLbM0/N75BKkpU0uh35
Cj3VEsNaULd+vkJk+swLyttKag5D/NRoGNc5zqK5uS5cEwBGf32Ya7JVLPIwGT21qnqBxIgNK0ev
RBUujfutOqBGgaycxLRnT/Sgpjkd27CXl9bvZ0esD1BDs986Yp9T1/gZlquGXMf7+6Askq2Wua3j
dPSFajTuRh2dj8r3p8sbokHPa8QOZ9JANVAzzA9KwcEf2+D+ejTtGDMygaZ1H5sm7RY1t3aVwYUX
9vx2REnfiT0Bd80xtX2Ga/it2oCIkvLgRUoX25xmnh3Gvv9skBwtJ2QHWC5QukfSn+5jjAsBrJAR
NR6IRw0cOrm9h3sTfi9lW0ZQY6OOeOhNFQtmcgdkhkY72S9w7DyAmDf5n0KeZpgIUfKHWrPKfezR
JiTCjRc6cMlKifQHUoxGNHgskJXR4RjasAv3I6HWKQ4scix3XkXOf3L/igOirZgrIMC0mO8wKwms
WPJ8Stuq0K1jjyUxEyI9zR/GHJQAcDABFZUY6JAjEYD378tQ7iORHIVEYrrk/m02buXKPjqtmRtS
R4E0Tg1I53thMfmpdeonF/JNkHukJoRczEF/UVI7w+7PLh3kTMSiG2s+Ibp6+XVElk4N3H8DpmhC
ANmeUPrLz/zr4pKwXL4kk02oqNibk9e2Z+/E1XuskvG9xmse0LwmUOCvbLRhRqN8OzSqtMP6+dht
Pf7eakBp7yp8Lo/BBFvtrc7JFQQazTPnm75jh3dCUW67XhBFnNqtSfFILG1Lx1W4Q7I9enisox1P
OrtwonvjxcLEQGmdgdVHV782vm3fEJvxFeI3o0fuyG9r1wSRHZGL8loG3AykucNYTtEWDc0Pzk5p
BOUabgciQePPUjlZDbXonc/c/FA55iyDid/7x22xf0IPS8voBgJOUs0M8fdPmt6LJivFuutwtksu
acqa0+cnIta1JP8BQFIcOQzJcyb6iW0fo6P9MSFKxBNdhwbqVy7WOzzg68wUmk5RGeOiTKM2Nkp3
16b8BmPZtswPUMpIqqo5/lMJg3tnEVW0RrRMpavxYwddbXwVDjhD3PRl95j0O3UVDYZmtbzW8Wdf
D0GiL5VOlpV00jdd+Winn7Jjr3x2it473r8Twmhr4Q5kY8IYUU+X3fiWPzx/CVhNwi5Dw4KoRMRU
6R2iudnydl8JbwAht+/vqONzMGgm3k9mIEgRAgo3mQ9eSLpUHoHnPWmUjd66NTXzG8SMor6xuQyA
Okw42AFoOdEubKEYvP2h27M+BznHO9k3OVms8EumNWBEjg==
`pragma protect end_protected
