// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iKzPRSBGVWKz95LQ6s8JuP2RRKtGyP+gR/ZVEwJnVjrUyN44hgHSalub/IbwfpmN
BkeSmd23Rujf/NitPX8cL0G1RW96yi/fR1UaDWkcsWcy4YgjW2PLwTGjDCwuyY/9
TIvganqE97PaBs8NuGoirA5TjCU/6zNAat7YCKpAbwE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18160)
xL+JTCy9JGGHxOx/BOXaWnnJDxUxyn4/U+7jguLVY75j/I7usiqHkf8kN14fTJG7
WMSEf7eKQe2W3ygWOdO/rpETcAz8RBtGUu2w8X7SM6QYdBuwlaD3odrP46/9kE+8
gUlso8leF/nHidM+tO5CBPwIsQu+SK1Xadn11Izmx+u7CDXEMSyhs/9HOXKTv2vG
/pQ98y/rTFTPS4UlktyIrn8xdVmVosD90jTpaf1q++iq/4W6H4AyFRk80X6h/+TM
s9xSU0h+vNkxhOPNEUETeyUiq3uUT4caDXdGrNNLoLK8jZI00v6Jj70XUlwQHpSl
fonizQbClVnrNjOEV7HIZ8gL9miPOqmDm0Ad85w/aYasiH/j+Zs68SF8bNuKLmeo
1+uHdJl57UGjpRhYXtMrlnCVF7jX9l5lbk5VbQQfX0KT+HZkD8OotDOPHtXwXXMv
HH6Ifc8Cwf6Sg+i/FjXR0FUaugE+X+7H1x5uVnW+yAARVcsaCnbI/f3qUAGR0LQp
QpIQT2MqnBljCNhg0BVITsu7qB5VlYWsc/30+d9yCpUaNzkuS7UMw9LR0FAhPW5r
GfaHGMc5fEMSnKuf43MVtU2iWuStqqMaTARUOWHCci1sdERXCtLROM8qsbcqT569
z74AShC33aMDe9YxOPKxe8IB+Xvw0QUQ0lQoUancp/Tm/cqjok3kUvElv9Cg1VAd
eArvk3Xp0bhyEQL5u4nfgJcsCg9vkqMjffKSbxcChDzhAAkMrR84yJWjOapUKsYz
DHjW0xUDlsTGYceL97V68vEhovRjAePBlmBwKOMPCstMVj6f0GiaLFXBV/yH8SyQ
iMdLDfzIFWw9GNlCjMFlMNVa7/J+xy/rt0fUaP9HEy82oXTXoHeKrhEZjBMbB7e7
tktz6NtR/bzdEy7JGfrqQ1/nZQ/qNTdj6BS3v7QrTpa0j4dNgHtcRRM75OLKd3l8
6rhOOxu7Ae9vNUZlXLwMxG04sbR6v7RP1bw+KK7tmerDZdYfbnjsSstAGbt84OEh
wQmqJ7wSUOm6HTUUMo7RSfohRKmg4IMLX72UicvEm/e7CjjMIIFJn+c5mgs+WbXj
pRfdf/ItIiAQOBE0D4EVKFvkfBEb6DHP0FVJ3xW60sKov3p3ojWetxUm5p7upJI2
L4v8QeuvA/yKl9UFdxggYUvkaPJip0mbt4vJ1IIFJZIPuZC+Pvt0mSmkmeK8zTiY
wWoeoEQLBAkeLbjuDc/hUDWeRPrrrb+phZmQZ19HIY5j9L+t26Ck86Z7lCPgAfNV
lwE9hSPpgJiOqxDNZxU3MBwPIibKMSDMw3px5d8xdv6Ytmpo64q5JuxaLZFzJnNG
erY+1dCHNLDGMfviKRUw6SuTPf0TXv9c0XYlM6BLK9igI1i3pj6Aba94a7a4IJbj
7AVf9V1hLs84gxosBQIKNZCgorg7Ld3fsnmcciG3u5zThDjS5gBkL0YFOXmLS1kB
4T4594k+Gei+PVrJXhc7QM4weNYGN74z/LU16OR/0fucnkW2E0qdlGhgTM2WURDv
0pSDoef1mIhcxebIis18Mn90S7+OlZ2Ztc/13xs5h4uAPkMQHOnvFEQzZ2IHTIYu
WViJrYUl/WhGZLOXYJhJjoraPv5Zjv/nTmrz3JNZgE+yRuKnTTsY2N0BXIawSrMQ
DUkUqjuJhVoKFmi0S2UIJhZch9V9TBLUd0EOVUEocTnvWVwFXzNwlT3xH6YNaqbB
a9SPXWbdZ8kkZWlREi2v8yIoXOZmRvWIgFR8rqOpwNZSSJZOkRHun31YNJB3c0P2
XfSMku8WTdfFQTUqCqa9xaR+RtadyZAINUVKCsFZZ9Rux5z1o1ws9bWn3r7sPQU1
QZ/5F0T97ocne/dMxs0kq3e+5Y4/uzL4o1Iz1mNe0qPlS+C0xcXBF22FCHgyqGwo
x+bGbb1mgQ2SQl1Uq2FgWOujEDq7RDjivZn4eECaq5LByg+MfCckwrArF++V1imy
aFlQzaG/bIu5JpjTIu+oFrfIXqlVeZDEY+eqyr89hDWjSCNaFszJMJVxKYC8NQif
VgQBP6k7ekST3LRZVS2BXhjaqUaq1WrRbyrqPkid5Y0iHIDKu74bdgyiemIjU4M3
0EELE2XBr+Fvnjb3v+xixFhcLVxSJwPkE9nIpmHO053bZRvKkxWF28aZ3VeMmaYw
7Qg4nQyrNdFRXh4S7x6WQXlyb9/VBRHHSmFDzx0apXd1p3Pq8pIp2l4shk/ZaNds
1CqYqFdceKQGPHvQvJzf+6QJ4jHlGRK+mCnjgRVypMeepdUgQZNC9UDXtLHFsvAa
+jstCWoN52lMjSKC6WbYQGugTir7LmfEkNrvwDECasIs5KlCwJ7mvDod7aGx6FRj
0RBLnVPUFFrKs7narm+k3XgM51SCg4nTHTu6RF55Um9CBsPqXkMANdih3twi8/r6
sIulF5vZWA3X6TIlTTcAP5byuhWAy21xn4NeZcKoatAwKgNcekkqz4IgucWZZEeG
pOOk+nTk2zna9Vk3wxpGvoBb3A6b85q/4asPxXrbF/bTAIRD0SHM55bQnhuM91po
2WEpc+zbrbsorjPt2EwLcqy8UOTIEFnzS4ehfWOGTAWccCkC9bvWLNCmAXWpXLDr
fa3uDl+z+oVGY5GQPeOT4oYPnUXUFfc5i9Oj0yZbMwE6jcZ/sBX4rZtmX2qekIwQ
iSwV0JZZE4sriUXiQI7728fgk0k5EExvImV/czlFJk5k98EQv/L8barVbzZ/cWng
ZMXcpiLt/UensXcrVHz7MPuHhoVUIrRSuTef/86dVE6KyV+d5BKhV6G7FpOxxvwt
7166O8b6xx/CkL8bQe2IkHpgOgfgOXxbfRK+D0Y/p0Ty4GN3hWOvXFbZhTv2sf/y
TaXdhIJXJt5a6pTj/6Jimdg1cuViKd+dliMZfVMaICCTtyG1Au484GCVuq9Hn78r
Ova2MY80IDV/EQKENbVlQoR/WJnXG0gjhLXE7uS8xC1A6rPEapKXD761vYnqlFXe
Fg3JpwNdy/7x4jtwp/Z5jvqqlu8eR4tDBNiq1IHzqZN1l6x/t7Cb1PXKsB8qS9o0
eS2gDz+HASFvc3fS7fWaGirpEGfX3eMJgRvUw3XVVN7ei0yePyR/UG5R5qysPBBm
bQYQCeAwesEnImh0OojwLcQ345d/pOWP+jU1C7Rh+gb2YN/fMYCBu0Vmz64ef4yt
tmxEYh6+X6U3c5VpaIDB26Ix17uG4nR+R+Tr2/XdMxdh9IZ/yCnajcnmLHKn0adv
dg0hToGiab7eEIlGF2otGit/XL81WI9l5cQUR/NC6iRi4hv2yzkWJUkBaGvAMSRv
8hI4kGfgTPiO/Ztt4jsUUfMTbd+7Nv8mvkL96grMR2CYJO/O+ZWpGluawxNedAnu
bnd8VDHKAOD4UN7/crQDT7cimyhp2CuXOrn2O6jb4tMzyBfmgNDHVLgArPAhy0Un
BbdMbet5l+07RfSKxK/Jn6mbSSTJUhguzj8lfats27kpXAOxoJ3YNOsibRE+9+jH
TpFG3OcR4/Jh19wvwrEQ0DYLt7R4w16AkKAoD6HzM9niS+UgGaIW7Br2Y/NiSxvB
tmbsRF+Wny/aFg2XvsmkbLNYwEP9AOZgSO3XCG0wyPKTk94SPYtxZtNJnhrJ/5vr
q+uWSXq707Q/lUXIP+2FuNDmtPOXM/SAP9gx/kN/7Xyxvp/7GgBopKzK1jW9vy4M
nAoPZLjX1iEozm0kBEaGn7FTWAN1hC26N1eFhzv2L7eolaDcKynO4V425+t2wmwy
/gPxYgY7BycCtNV2n24pIPk6Ka0zWdXgPp4UKR5p5O1FR/t79bUA1lzPaFK3kxe7
HypuJZjkWNBNl+AFZ/cu2tpDdH72tO9Gzr+TDYyVfT/YzaSeKYH6fU0qmNpP3O/I
cENA2SpzgzrAnC0clhGy0WGhmagQJgx+YtHi/X5SJw8F2WV8/0yDSNEWGYsj1gb2
7S4rC5OAF27u+qsGL+h504o3GsS8rnmjZefuQ526q+02gLuoFpEsE6ASCmM9dSm2
P6Oxau+OKrXk6o6zNW3vLlLyWtgZr9WvGh7CAtjdmwOp6I0ZRaJvSDnlj0LqddS8
OjAqjvxnapT+HOn04C7ggAs5qgiJ9uTjrxXqWpYjXPgOUUx6608AEOEX3quBmaWl
piJTBKyblVQLJv7Lyo31KH5Y2gYkw8xMftaTV3NeGnDWSwpTWprcZFQp7xRzF8EM
rjsPlYSjfXksXHYPoAMrFDAP4UzwkJSoqGn+xY+ga9s1Updv0PlFP1XhRQKi/qlV
3r94DWQoqUEKIo3zB4hmpuZaYW5qEU/cKNeZUaUK97awQi29zZBhvOxHXkJxL7ye
FDdo1tealv8+iaKCnY3V1AWA+u1DMNG5e5MQRNGpgByKLQwqRI+hIYWKNhxvm7P6
erhfw4YeHk78Ufu+ICFy0zh25qFc9OLWIVl9Mmnd1YLZN6LpaHkPDbHGW/JNpZGz
nsJybTECKWKu17eND0unDODpn0PYZMJUwnL7829TFX3gfOPqJpW2SEQAgzXZlaxx
JVhhefkYTfepSaY6vb8CMgXAK25o1G638lu8SBMoFe8suwQXN7t5dtzPI4A9Lin6
E7Tq325FNSgoXBV4OtmEMGaOhWv9+IVt6f4Pb0+w/3gwvk+bUpBBgC438CjzMY4m
Oo8K+l93dippuP4FdzuuJv/Nd2P8IfmsaKprYrbZ5FMs+7JreUUKTatJeM0JlMg2
jCdB2UILT7I+V1p4vSdYHRlDkHdaLCi04xXZYNh217mhk7Z55kaHfrAnTbHEd+LX
UI5fpzo4q62PyT3br3HXJL8vwPmNAAXGbdW2n99RYBb3XV2CPYZwMMuEYSBEkPOb
QRhOlIt5TIn+bcpECwgt8lJCY5OVx+1tkagwreXL/5MVH2LJcrX1GDMp1dOL7qLG
Whk8j5WFQxl04JMMEXT7OTagDwEFE/1p/QOIfXb/eU+A5OIaV3Ifvw6u5tTyE+1G
L1NiiguxscuaU86+DeWu9hrpXSTDoOKKp5vzFMZ1jr2aaUl/cQZzNy6cI9uj9Zas
ZK6ojhwSgXt0wv1QQZjMPNfZ964aZT8PYK8OWUePI7RUgy37IC6mqamEuhH93b7K
zAcoZ/EUqaA4n61fjvIHw+PfdJxWevV8xXlmCVX95cfO/nEHRmtIIPva7vq1Qumo
RLCsoe/M/7ub28fOHh4bbriG2ilbqz7iVwoZ7q9BvmyDh+5v2DsAEkxT9qujujgZ
pjmACg2mMfqW2dc2AFE0hMSFPjU9tPte6BZBLwMNRKrWv7WQYHI+yTDFKsukbyD4
xZaDTMenh/iYOW+bNNcZBiaYX7axYuxkTdeTHVwdB8LycBztCRck+i/Oxr6j/FPQ
/PMlFrLUOuQRLLLHndYTjB9J0VjJZLtTX/+34D6BG6MTQgMGyKyOhDSCsUkxvvvs
BB/ey4iMuX8p4Qb/UM2hX12Jpzh4MavUjcfuOxi3chruq9Wb1p+3GoDTCl6lNZhx
NAoNjvnTgh+UMlwv8Eqf5EZVhro2fMdSgZqW3uMCvQkHNaLe8FxHZyDeRz147AMg
TO8sfdnf+TT4ui042IRy7rEcATiz/fZDDw4ndCukeeAYXs/kb9kz3vywqjCVA4o0
KhljjkXRklNozTIqvnu+N8OF133RTbgyHnSfFL3IegC9tDus7sXarZZaTgUIg4Yk
8t0HIjNDmrTMCuTzfZKMf/vyWMEMu4wcuJMIHCMbGD/a6AeQE9HkMZnm+QuJ/XfV
emphznPiDk9fZj+SYMqpEVTeba4ICDfcjdZ2FvA9BZ2+TwILLxJ0bZhdZtG4EwER
ltnmLmTeSnM3ylclCcxu2y9a/SdWDjAxQx0H5NARWWNQWhxu/sJ0e3OCudnV/aBN
QXLs0ghaF229E+sWOkXVzFtHyyVpqkcOfm6UtZHw3JxJZ+lARMmlfkW8V2eb+8IS
HHCPbluyYhPjh0OV2zRb+vJnrsokxrI/7Zt4KFJNSJuB1hSonIklNLnulLKB85FY
p/1aLVYPT6/OE0loj7dWoVlFuO73QpWlNQH2FGUVAARIIwMyMF3JcE3oPON2TWSA
AVH7OQoVletN+YNvUU1eLCcOPjKacuzj27oQykKeIExmoC0rWbq0TjH04UOSlsbY
fMAVHXMKaNSWhW5VHdBRao92n/yQSNhnHP7HYdJ6AJz7RZOImRY0w8I8UKlPB9Cn
gkSLYJIWIsDwvt/GWHkm1/1zszzPAnD7NmA7ESRRUddxEpzf6Nwhv+U+CS9tBwkf
S5ldYB8jgATppbBMwKTXtCHBu+lx8bmtddMRy4oX8CS3qpukAuldlU35EV5+nP4W
6e8T0hABaMwU801FXbr0gevG0Zd3NC0kUrK936RBnZpEsYrE/0YTzu9gzBk9MdRY
JWg0tABdTVMIG6eWDRbSCBT4LE4/QJx3qpYDzoylAsaYnYFfv54X7Nnr+vLtEawA
zJXIrml17bz02uRC1jIaXts49oAZMTaP6GJnPaWPeVYfbPV31cltKw22J4mSuHON
a5Kmn4xl95GnUaF4SNDsMPwwFiaEf5UgnXOFXSsuwre8Dl3ohy6Qf7KXD7eJ5GH6
JJzZ6UbYEyeb2uApTR3NNf94Fwim0aoMTRm0I6hou4lpqbcYNoDRhn+FfEi5CGAf
y0ceETP7GmJhpy6/AMe+v6XsJw9TO6lQlYFiX9RMojUOs3x22/tPmsnInZ8ZLarG
j5q6+30tje7iKuhRAHKaGI9wf3GSiPTaQkpRmnan3ZXOhVhlluo5zpm4gMU3EzKU
VsNKMm1L8lcimIc+WXyP8jz5+pZp4aHGo0U4SQJPiLlUG8kduUykuRB/ISDKB+e8
NaUNSQMhu2xW8QvVSVL6bnj9TFov5LVbBe8+e9HgbHNF5uciQKZY9J+f9+Gv/GFc
EyUeBQYoExt0ybi0PQ8xEbCAYYqIcrPELC7AhekK1B0ccWbEtzN5wJlAHcimgo+q
P69MKcmfXtze1i+2IW16Q6bRFmiLDvlU+w8IdjfNBqFetBI87cgP57VwlgRc9zPn
PmyBQ+sQvb578UMgR0VsCaljJveVjPmKvfPC3amsrHZXCXx2jM961RwUCcZVQxnN
K1Ij7e4GKLoA4WSMRLYRTPb2dcWHc3SagGqZGW994B1vbTsnZ5zuNVwFLONB3SdY
f6sg2AfBWs8pcWu3o4HZwisWdQS0eilE3RS4IKe+C4EkAXXnZg6S3mJjVzvcdOZD
BSSAEteUyIrUF2zMQwhVsHbQCtig2iNtf4OrgFWtZU9JinSmPIANmHXVJzIqGsHk
IOyqdafBD8tV0clH39EhLE+32yAMxkEIMyBp/KFjl3b0Eq5FbcSeYYvjJTq+FEyN
eN9dZtmDS+8tzYEL9V6jcCQqGrIC0vbc7A7IMPXLBv9etuvEI5GnAXqvUOlEzHm6
n1zLzFaKPIYwmqtgttgZdcFxdKrpWWDtSxp/GNDJR6j2fR3Fxvl38ppKD1CSmhYH
1BTl4BXvNZkHcQchjdEPtOg2M7YWnHE7js9fE7dZLQDI8hWAo0ORcHPDsLrKywKE
7ELWIxvpCWjI8wtuhKOLJbuIEC8qJihdIGFjPcXHFniq2jxPAPaRZAh1CkqXxrO/
y7Ui1J+XJYzVIrjjkaiYoJQOLGbOZ+ale6z24Z2t3b4+YMob1+Ca5+/UNCxbylNu
ijhhu0wXluQvOGXAi+WpvJ2kaWIU1rufBx4gGjJrGc1aLpuir2caJSofFWlQeF13
LH4zK57yCLIQgx5wgoF+WnuI0n8S805oXnbw956OhOqu1JYJT6l5NB49ZxqPQJNN
nBMqwL4wVFBAGw+fcDa/iC0dwQxYYCPvSdVJ6CBSCUxXlDKN6D3DjKg0Sti6A0A5
ckA1B2xLC0MkBLxTymvzuvCChNvMvOM191wi2LauoEOmYi9jUGGhBXnT5fFYhqbh
6SzNZjlgXKORuO/libbm/07e7tDF+OTadPhXa/lHiWssTD5KjwmXHU32k3BuUyPm
9mKyI3N/pYw+JXA6wtNIM3TvegEjy9ur8WthxAjxrf3h3z02WJM0AjmCPmou4dB3
IPR7GGLAfvjlwiCetwVSRoSEYSJPGza5m/r+uxA6CYw7Tr1VamS89orwCWICrWik
Q70udZE0e6pmTUCu3U0jWFa78NWgpTwySAa9q2vomsCGIr9abgLNU2Xyeyutyr/5
/SZGh4hXGZ8l0kxjAK+nVB3LL88mv8IbGottzZBuQ6cLwZqIfv+cIYfLYEJoM2l1
6bDOG6bY7t1n4Dgre2kqr52yceGjyzkuUdKeelUR2W33e4MopqzqIi8P1yHBGbbr
mGPzdQ0DFj0INtHD7+NMxOsW4aYqUwnu8sGcm0LSYKMfjX5y1w1Wecc+LuOz+iLb
3k3twXKu2veNyrGZ9qyW658+1CtYN3HtDwgLb7qBwaDEYIkZqFMiq9KGAKtAvJ9o
F72N02ueg2sQxfUCfRYbIUd6zmHYrw94CHlEHHdKqwH7OpfSHDKPxIKWEeWQoPRF
8L4qMyjoyqIdH6Ishh17dceRSEAXsLfNx0snlC0aZ/3RV4TQM+oooe95yrv46hsz
u5ri4VSotlUaiVJLZaGI/BqS5ni8FkjW7d9D8dLuPTsr++McGgwwDvjcomztN/C+
+sE7WWLQNB0hYv+kkpTZss0Pou3n8wgCWfu2QdM5Tvfn9Zf+67cKiaoYrqwWBvpL
lT86T4ka30M4yyY3LgT+Hl0YX19Fxet+YZMz6HG1C7+56zwfqT30EHEFpoi7XsXv
GgYKzsxCkB2WMkvbyiFIsBSiLf9MkSqUG+PI3Q1kB87DiNQhhOsy4I9EmY9TtcoJ
fOpUgeBNHEN4xPktbRMLRETde86NVhbkFluqRtLi1KWAcGLH3/zZoNLP2KBh5u+y
1dRsWdT5O7+Ze1dPsfMgEvI2rXqq7IwisEDw1cZjcMZPmfvi9sv838pw5K7NKH56
B3Ig86jKFc+NzRlY892/ud5+C8Jl9orDY6QIiP/2HgtJFsLlYvteUDQG0IrXdW9r
flgeQuC+q9RfowuWjgHXK/C9h1UjwhLqvBS51c08rKFrHEQl9RON1Yo/pV7kY82A
BrZu8XzuIiA+KpAG9eE2q9NdEKyxXLNdjbqp6PIhrvp1YcQolMjp0+4qZbT5tJ+d
dB12d4sz4JW6bt+WPFo6m8v9XMqnooZBATFS2k2VpHDxMz2QRcnUzoUE9bj6agfS
MpwmCx0pwChUgraCuvgCbpf6vyBgmjuaXhGh1VEVlrLa+99vAng3J8/uEYTfPjft
tKN3kjgHuqfUp3f4mLCv3YEuk3v7rbjq68wVPg23CgsfzzDmPcJ3cBGV7w5/mDbe
a58pY7+ndSEKsU8sf3nw5lj5fWEbUlmlDF0Ko2pEE5glrvtIlai+ZKho8p+1dwfX
Q2SmnndqFs69pZxnH7DlbFyipPA8S7vmQkAT1z5jG6o3WCUXzJZtRDS9PfGWA+9R
w8YZAglI77iFIYjPRheZ6oGbJ7MQ00ctANjWJ6/TSK4PH84yiKnxZD6VF9bwEA37
qoaFAyRtoxwZVJ/MCYPwj1DtTIvn3Gelgj22N2/YAwIhK2cVFVTeqCsGew94dmAy
BnK9XGDra5KObBHarDOoy6I3ZWLsbpJYWKSIYS/8IzqWPUZZor5yGP0mnDzPkYcZ
9NJ3AOlyLz9qVj5zj2t8vhge5HA6S6OxMpJekb2Gx4UuM+pAGFABdCJy7gHcGL3W
upgbZ73kmG2yoUd5IU6JyZ9XPoS7K5DsptaxxadBh3eOI6hksOg2Me68SyI3tcxz
hjqemTNfkGKK4ink8V/QvD9CTRgaNbDpWMsXzNj9+KsDi9v14c3OJ4NMqkhtxv7M
ZWgWl5w2dw3hZlimk4lLPNV5GLdBJGID4kLN/Mj3OuvNdqAxNZdw6aKiyyqJl14A
E3u8wdGEwqbsyolceKCX8Y/vHVOTZbjSY6JWXZcV0B9PtzOfeOWUxn8kwHg3nqjO
yzQSv/Gxlm/PGICnUCMdqXRoP5ZqjbLy8ZDqwSfQCQqP9/K795NJt6+ZoqSZgQyr
33P/ZS2yamxLEEpkZOvMIY/36jYJPsq4WVDuqx8Mkg1pNYzTZYIaEMDsKAg8z35c
M1A4toyTA24xcZGz3tb34Ld8WXfMJAXEYMMVxYwNDdkLqjaypmq3A+PSKmTTrHvM
BS/+reyHJpwwhb6AguTbz6qHUUVBfwn4mdA1oLcB9P3bk+wtEANY/x6V+D71UjwY
KqMV5SwDtib35ukHgiWJDA6o6zIgB53TEM6EAATr1TMPSDk9jZdDESKEHuDXhwfs
Z8JkoxGQIi7nnP89o5hd4GD9vAFE+mXN3FDtjSmiDommq3CmgQa92Z18EDV25O49
6PB0cLVh34/tiAsLWEnNeVPi9Mcr6qqIPrOtZt9MzUSYw07P8ZP7tASGWxf8aVAT
1/TTByQPnuYqrqdLQFG55MmuvgJEM9MI81HkCvFG7VC5p3cVsKQDB6nOWwuDVdln
T3FbqxdVokhqlx0NRCMrRku1nRil1m5FZXRfUWJ1DsvMRA7MjNYerUmWkTuxi5Cf
L2Ta19Vd2jdNeOnhhR+7ho9CqBtUZx3lzccPd01iF2wUOQxjqIINStKe7eLVD8BC
tBicWTd4DgG+97nHRFCf/Wdtiht67jxMLcv6clYtdxp6MWGZxWMlbogOl8bq+ecn
FnO873ls0q4PbZapqIqJvw98RLlrbiTH38l9JPEMl5YZhtFDTUMiXurctGWXhQPY
AxUvsDa2jK09RHWLHK8lp/LEYykC6p6aYdIwaikQCbymb/DZviSEUdbex6UPjH5B
WU81C4nxY9AmuL1/zZdDROCCX3lQsNvJtCi53ncXFbGSPiWAG8Kg0DyC2J+SMcQi
Clwxe4ukeD7/10Grs8NVZWtIn4oAtmj8GsngMEwN3l6V5LnXb5Ddrx+YgENyutJM
srLo6Fk52X6cxQy5ZcjzW6kNejc0jLO2VTGS83SAkUDX3aiISyTEiirGZ6Mzg8PT
YrAwrM3nbM9qJ1qz7suLpDiURzMxq480bM2T2YYlQrnuT/FGOH6i2itoL1EPdDVZ
3wwkTakSI2e34PYgnxvBL0H+ucq8IdKPqu9ofDNePqCCCJaoTskGElMxlEGnSH+D
3mIVDTlW6ukV2jXouFkkGnZJFYC9O3/z/eNv7YCr1ok187BqQTnw6AI3QgRmqYy5
VB4bglLScBlVXfxr8PRQ+gI+S97QIJ/Zv3MiBNoPORnTA/AumS31AKkKiRat4QKo
3z4HvhYabftUMPj1PKixrpB5lG4wA7YSk3wUIiZmita2lo+b+GTAKeMhYwtuzpXI
oZkeeFYUITDGrJCLrBmsjFpoc4OsGD5aA3RYif2lEgyc9pTgd2ALJEkblilqxt75
xucVgvV614Uf9dQI1vm4j8hHSnnjTWPiDT/hOP3FMvN2spF2UNrD4ZXVWq3EU5R5
m/CQGv7fYk2uYbaX2QYOcphf4foFhPbHk4hJ07Wz9j5M51QA5Xobtq9Gfh8rnhvc
/3HTQK3y4ggkloRoT3HiF/Z4DyoTxPjXfrzUss93qGT7VjL+UTl28RByrAy2lHFh
kECiRc6vwuczqu0FJI/ojS1o95K2lNMwtAGB3fPpUAQ+JOSHK0FtbZ87RCqHJXZ3
OvOzUomuTERoALe42YQvSFI81TmuhkqbswB0neBtLmWGMLUxFnvacCh/qZTIYEBI
3hamX1lBCtiwyFzEHuOhOcNyvY+Iab4x+2gP040nY6NN0sY88Z6NVlaPPlCS8Lne
H7QgJafCo8arkUVk4kS9X0wZfuDSJtoTP08YLOBhWzgSICWLHokH0mlq6J4ia4Hy
3B3WsH0MqhJ31lNHiKO6nZ8GimRYOzhjzqYLyhZaip3tzsDC16/EnaeY+D3HQYVB
/cHRcqmH6ChfuruE8wfH+VUR5XcyLP0bGEsMMi0iIFge1o+YxHDGKfIRRdeOZo1d
LK2N75pZtlPeQqcXTfNhVsdI9PlMuBR/860/ifr+hYbEiLCojnCPO9xdVRYZn0OY
z8pTnBRYFK4qM+rJbCi1Db+3lriI3WJFKBUpEjirFGnoBaty9Oh45SVwhXhGc2Ap
6uygyQmFi5/1jOp+b7yilvLeZhfU/sC04CYbS02oLWsyLAWA2y+4iLp/D+gpeLfk
EgSkw8mcSTs5/mOD4Z30B114LyGSL3a2vEB8GhOarHfJ5jmT2WQjkhjuyBj96/QM
zzfx/ykW8vo9+aFaQQmWjMDp83PO5ymwTKF2kq/2juS9oFOjiqdtjA3TwXIAnNFS
qBgvcCuHb6n+j+JmllGxZVvAIgEc7O4WATOWhw3K6FQ86NPPSlMvYM9ho+6kQEPD
BZgMKLGc4dyKMIBuSQ3mtLSysKBTrm7KGIh8lgnWvgdp2y3yKDx5+rWkzxS9Uo1Z
2FzUGPfFmaQwn2vve82p0C8Gr9TPinhP+hiZls8vHIAm/BjU5FsmXMqT3nncNyhG
59fZN2bzzqC25W6q1FugQzs1sU88V5fx96tXfpVeBHQLF69SKdrF4j7ymUcRHBCz
5zFgdeQsuEjdjBQtTM7Mq7HOAW3pVigE1LJmihQJ9sWKCigiOjXZvB6xKtsokeUU
AjqB+bo0nLeXq10P/4kB4w0W+UVYrmk4q1u0a4ZAxU6D/6VVI6hm9C9sqxkEp3EB
U8NlKkveR3BOPbZoucO/8pYGgCQoEnTzDRbFloaat3z/ztVB1oLe98wg6+1gFpZI
mPriwyt7yLkUop7YlKs5Ao3cypbRoJa7Xs9rTubQUHX08N2J/R7gy3+BA4o4pKBf
CcCx0p4XJeK8wUqffNVZ9UGcZaieT56oDgjUfCPaAFfTVPXSbcGX3H3/yyOsdkyP
cfwhCXqvyyfRJgIA3WBuMGYgvTA9ZlfAyBGRO0fZ8YhPAnByfCPbequoUqAwnqFk
A/KMIShtZSC7UfsM2/MJcj6d1KjgX27dS1mMoPtyhmg+Dv8oRoCGVFEuIBzyDiFi
KlvvwS7fJPoCmjpPtDHXEwtD8aq/9tp1dCiNfM4j8tz4LKvD2WbxmrxIYScTDgK0
pJD7f86AM84Ee2RBuC2GUsK2BWJhbhnRjfpZq+DE4dvHZXKh3GkKn0q0m0RO9xnt
xZGsASL8SBzwhEpEcitm7jZLTeIRJiTGzit7PNv2RDbYP7L3z5pf/Yw5MzBT90O0
oOXNujO2Q5JEukRwCWE1DW4+hkT/dU4x+vWmPmVBTRW2zT+zZ57dl2NVIgS+RPmZ
5onRNl/wwDZtlEJW9oKq5IvuKF38MfoF0WimlpeNRvhzYeH/9DhYQGfbJT8QOcMf
CxTlnmwigRvH6o6lVGFOeeXzla2i+TunVn8u0l8//kh0m/W8yHnl4YLQ4R4/zTjv
d3rOoTu+ceACI/VlQLgmHWAkcN3qj/Yfz5NRnfNcTID7gLZd/VwnIy2IEBr1+CvK
luTTKqPKXQVGftaeitJRUsLpCa4XhJ/exNDG1jeaCKI/LJKRIdDHO4eIDNUMlzy+
fqwmLy2OgdTrsYJ5eeusDwmWGMhzNPa5sgulKVO8VWuRdhlxo8sw/PN/5/50457M
avHLq7/RtNT8c0kt4WG+/iqj2GMir7sPLvUcz7OeSY2YJ+StzOvUob7IuzeRAyKa
0l5wk2LKAYmIt77xPj6NZ8GsR41E6gKPETvP1qzYcE/H6h0/J3DtQA5TAuydeSHg
jLBgQ5vObqBgrJELRYbTTKXlwrim6xsqUe7QDwksjskCtOFgCBjv97j2uHPYhm6y
Jguw/2tCcfJuGOgyCz65EjysNSSK3lUEZmaumnPfv0Yq0NAwcmEhNIa3KhN9eeqB
ld1Xe70yibLfIYG4IQT/tdjg3baEwMn5iOooviQblicaEGBeF4JhmmZBbPBLEpoq
VlBpu6VYwLPP6EUPcWQRnQVrLyhfNd+6+mRNGDeqJFpdqFj9afR4HEsSK9jhMtSx
/KiDEYD9MeUaiVd5PtMyOUpH/WV72R2XPzs+MwwZ+1rflGai2KLteazsNrkIaeI5
GRfSKa649E1FLEk3ImPythnGO5BC9bQyVRN8eIPpcZqJpNZUi7ezWayTN9c/3f5j
0GarBEjxa8HsmWhqzfxXM+G4Rw25MCI8gGA1rE4mKEINHpDl0mFKTFHnBMmC1Xpr
/JKiuCOR2q2LgBPJ/X2/GLxTnT/Da7y6rW8Ma5jQsPLs1cJmGYjiz9Tdu/WFFDYU
swElbxN4gmFlSjcpJSPpmepnp79zZxamQS/RhNlWLjU5LS5A7tfYJ/DFMtq64kzt
Cu2Odaur1z/fkgl+POSNhfNgQwMmbDVn6aK+J8mNvziyJXhXba3/P+XkIqBbFGvo
eV5hjElt/7M3qIZfu1CSXFqkIgqs37S2FD+1fZrjuo/WGpPtYqxeEWoZrFUWLxZm
gLNhjQgaE69GcEbnMe06yhoVt6gfNYUY6/HsDXpaqiN56NVbj3DaiuBzRePsJ1NN
8BIO4Ig5+ahHDzHKHLIKMeR24Pvrau7E8L6WB1CHtjY9z+rFiUSlN6HhcjLgtUEk
w4CiR+fbRWJ5XGNBHQpO+jveUDC5BijYv1BimC/kyXpEQtKz+r/C2u2LICRrOKsE
mc+M9c4OQRMF8p+qzcgQWcvwJf4aVw1C3j5W12Ub8VS8N2STpDlPmkSXq4QCgCIF
kSsVpGE4/5T2puCqCzmfwdZE7u4JHKxogyEjMY7CZXJs1ZvvanAwkbaeGmXrhXwn
pIyq99XKG5qoxSIUWPIXm1GBVJ2xPKtWBdGZS9dbvbC664Jjst2wmckYODEOxuDu
qYKxxap9DU8nC9xJfa0HPkUi2+THDxLwmwon/Getx/eqlISraB+qrg67sX+dqtrT
ARM4Lovvw5JUUkOBifU4uvzl3MSJrP2LaWlJNM6lDqzV/izvszpWTgINkd3JnHIO
AW7/7+S4aU6+JZi8c8+IInbZhBlOaffRmvaACi0tEGKen8Q97eNYdv0+kNYlkOUL
gU8eFBkFMPEfwbmqPl6tNDWpP3IKF5RQIqq+7075m0vv1YJ/WDn9BCJyzakz/v1R
HzoYigFsJtwRvM65Gfkw4A17jdaoy7u1tgBzvNQeXTvKh7/EVqxwTeI0/FADW9Pp
rkR4YxaQoP5yWeYUdz4pUXhvVDGsa8FnVOSy7F1IzAwbgt67dAvq+fq4tJ1UDIHT
eHdxTIkR8eqvdzUmLV2V24TZtePf55rA9KtLX0yC/lPFInt5M0a9k5dWxohqFMff
L71e9pmJcT/abeKD5xrEUBFPbR4xzZf91HfaZZD8NYDW+1GtnhaoO0LEXCYzr1r3
A3JwrOJtLEJTrrUxlEi08ZYxHIC6K3LHMtwR06FaPIydDS9S37yMycMMGG45vrpp
5QMOSjlPobASj3RRQMd6ZIK+KcGiWWlg0KAO7CzfdvIaTrc7geFUUEYhcemh2L0b
+25m6sZfMbpEWswf76bcPwGMuVkCBWRJReHFZboI2L4ER1QmZkcpw8uXLMVTjvEd
PL3ZPnnKw4VH3Z0CBXhWbrYOk4cFV94rfHccsLiHoxV1Paw+ExTS6W1BTC175yq3
wsI+0PDUd0lQDykB3mmoEWyDpBwCqpyW+Ubz4JdxidWKACTFLzI4YIBDUBbj7L8Q
kjpPx6LUfjLuRVfP9M3SDofuOsocinOgDuiYOaW8a3bX8Wv9yHqpSXqqwTHsdxii
VPV3wTfq6yd7Y9MXVJDe6GShx2TpLiqZh0UJYLPB0iNstdkTCrh/bqoBZGWv7APS
StACwjkSEZA+Zy0wZmdp/Gm4+Og8non8D1zwihcTMbZscIpYoDG0/Kpdt/rDnK48
K7VhpaBoNhXqCBpLNBACd6Lps33oxJrapveAz9vNJEENzuji98ZcVw3aCjs3qVrI
noUvDNMD61OCRNDMknH9912NYh+8oObgVLzLhQPtA3aVCbxx6Ppot5BmpojiZQon
SiYRL3wZyt5vtGvHQfzbI93pL3Go7fPVFvzVeyIe2oGKwmvwLOsYhClO+S81rWST
IJzwyx442YNu9NxjbIdA9WRWmCu5Kvt/DCOefe/x8KxBplVYQ/nPNa9TcSE7FfyO
kY1hcq6IaSVf9WKEMaWI4bElREukFLT810yjTm51J0Cq0DA9Sktg3PdHPDPw4UOZ
Ydzg006rwcBfWuGVeRiH+zN7uazEB9KtyYTOyLzkCMOd7EmGq70HmO6xyJfODW/n
xz8Y2MdnwVaR0SfTapaqsFo0Uf5ZtjKHTrBTZrK9Zwt9tyYWxlVMxuTzuW5F97aK
J9WOt4b+/Lt7OVX9d0GGE+yksJ05pZb29WpCJQuBBN6PNejxsMgyV6BW7Ug+TaQC
nQZGH3S7UXxTBCEp1AGmxuWLnvGdwrLFFYHtZ/JCHsuOiLKCD9fHkx0cA50MDcz5
ksmD1dqMErLEejQT9kkfR/Z4DSLg6wtPViuTlLpgU2XWGS1Jf7CH61Sd8SDZrWh7
D1Md/G4w9KCV8BgJQHHttED4zMUjKz892ZY4V7UYbaeC57PDfqAbX1jAKe3oIksZ
JN1jK/S6Wa+7If5uN81WAGJYP42OsYzC/N/VjBJX+gVSllzzLTIclS0nfyPgTvad
I8e89Ey7TouYsCNiT/++qo5/EbPrzoPM54RV1256famGZH926FA503uTByleSQzK
NFZMCcNuT3wkgPjktl/zTDIAq1BwAyO1WOdE+XWfAVwqpX1Wj4/iCCbvoWbY4N5O
LX5dCcS7Tc6uIhqxQvArBZe9aQPwb6xo0Ic+6UXXwTvYcz83sZTrJRNbw+JWar6q
kO3V6QO1Mx+EGmXl8FVP5lnLm+d/94qdzTbkPOsIoUd5kjGBsHmm6ZHI+sZ/USwF
dSSIvebkabocXwOecQUcVkWSUV3JSjrydU29RAGx+zC0U8MxhyHpOXdaEOGHVH3i
5V+pinnXX8fpYgCPbtF2SuKMSh/wyWSlBBHcjXXVKy7Iw4tyaGyNhedkGQTqAUEa
If6WQzEsOVQpygLtw600V9qCp5CgaOGURlIywb13+gYML2UoHtwZJaTZ1/LrWNqa
eUIWJrHjnWpNqmXX5CR/rlFwJsZIrPhPF7gD05w5s1TQ9ZrxetiLU1I0+fjlYlRs
zT95FzReogDU+RiIww9OJp+LxbFZLQqZFH98cfmdXPl0Gaxlaq1/qSXZD7TLqoET
0al49Bnd9RMnNuvidy1dsDvYqiCx374uSyFfW9Vvf03rObnXwRW81lx8IxBtkBsk
m9SyzFSQmk95GHJsV82gjJCGfdQQD0K5OFOkMjp3yjYPjNufjDsYZwNAXa2ffsnD
kM1ErkZk5KZRZrvjjlzLGn86yi/g+Sn5/lAGLLZ1rs3jwzyShuj2SYifWeV6t1Pp
b9SAHPxdpdUqNk1JdOLsMJ6S+gPE4DZNBATHhxloDHOdZfVQe5p6X+mRRrykLddn
qEz3R0WoWOADe/7lMGDLoqIusRxD3Vf1jskGNiAAyO0Y9l34gppXSTwd6m6UmZG0
PmmTpZgw4KHznYtOiVrR7Ze4QqQwV/UK5evy8WHhTtweWIOks3pwcUQQlNxYFP8H
JLcLLG+72smbwfl5ltYab2/L4HAUqvQweG5wi9Nqa8LKPs7Z0qzXTQeh9fYafS6n
+ZUPUXgED2CnMp+iZLKvmNVqIcfn3/tM9fuWlNsB+YrVzDasQozL5BY3zMfmj91R
VQTuS5KYkrmwVO1ntNdqGyExGHAH0cAB7M4tP9O1fuJf//kYXuTl91nzu9bH3ot+
EDs+ohsv2Q1/YT/aKPRjVmUuYsJpv3kNs7ov2hB+LsqXcwkD3JjBh2SbvON+gxWw
1G55lRcCvuyTCx5znHc9YjxTpwHiCfb6TEqWXxuTq0FmTOTWxFq2XwZ+dLS3ucFt
HZjdAQPL0Q9w55WhqRpNR93n+TNFOyxCXY61tk6O7V+Mf8GH2842Gy7FRP9g5hfc
qDhc1eQ6/3KFM7+uij2SzEaWFNLHK2GoOjLhrUyEDbdNx9wEohSaQef1tl19PJCA
D+pjvgsZyK0QWggDxucXjZJwFX2gboj0XJNUo9eezWnAGT3AVBcqnOs9knnJn7ri
Nq826Qfat9SRP5zRuY4y8YiGYMTHnBvtuRANDMBaknUGli5gePro5GBIXgyqZwnh
Wge2EOtCapK4gfWzC8n746XNLiWx7p3OWZQFeb9MpECHcI6umOnjr/KuBZaSJJaO
q0cJDUzXWllXnVBXAVYkHQHxQg1z+fHAby++J6Mf/QbjHCkw6H5GYofj3DAcTJgM
Aichh4JbYMal7KQNBNqE8nh0aP/oKozoVDInqF5IrgbwwxswX5CX83sMnC2iNbrS
asfV7PNax5hFgGKgvjU19NsDH9Q990WAJDtsdY4+orFXm3rFNYzPWdSUdSf2FH43
P3IliLyjEjGLT9vYveoU/e6Pu/cWsSt0HfIoRFiS1W2KfpTf8YSuA0Fq+9kQzpwF
faPjD5mRqc+N2V+Ey52aT+73nNyX8rxYRW/VI36OSKCxrsg/C937N4A9PFxmFvql
4qTMSOh4dIAqZ7aJnHbTfXe7iN/ON9Ck1Pg1tzbhREFnO1qMg60kagjcsHFXyPuC
/edlBHY5avURWHPbmx/GJfmCX7Fe5RcmBCM6SbKSdoqFfU+5MwvgZs4HQAvNodFx
7s6oRIoFGC0hcIUej5uor/h64U+MkU2lipaMVYUQ/qOXZ4g9mIuGOZAvL+wuDFSW
fqwms4Q7SzsmuXD/Bq+xavpG4V4nRatndVqM++mW/nQeSn7U+kgLXFGmER+Tgmnx
TzavcbB4RmmYNHE8H0JMlp93zQy4d4no7wc+JVO2r0xGpkVqlkz9+v5paRkJ46pq
QEapCw+dPzYlRheMHQYzov6r31ZftstmMqmWzkODqdXQiv59Jf2wutvoUJuTQ1l2
BAr1o6BmsG797VZiDEOYOnVpAvAXnXAgXaDAVrNdMl4JMzu+BFkEcsRSIlsiFdV/
sgqIftze+p+j0sLjOc7KBTghJryysKlXQa6Tf5xOPCmnxoUfx+YcRKC1w5oNLwPh
TWFaBGuZvfZMQvODdWNTcqPfaLywQ0Alko0iw0ZlJz5z9tVGZxuCBx2cJ/Ca16Es
Cv2u4/ZIGjdZ0s3E7/nccVFxostXZ5m+brzzU5FWbltbRvdxox71EiNT6eVgUmOh
kFw0E9dT81F2IgEW8tDsdmAhd/tWDz274oI6MMFQqi1AOI1mN2IYZYVnGxT2bPrl
o04pwaI9tHl7sH8kZld7FyRHDos+I38evCxMmN+k7h/SfdksHlAHP1T/4/yBAKcR
RLFH9Yp0nFfjia8T16HnxrUWA4wvB9LSW2d5vnp6vIaNebuyLClc17U0euoN3GOU
oR5i05D7cof1VyurTf1nCTZmLg79Ge8hf2O3J3oqAuHvat0PVJ62HI90WgniZ5Li
qFVYeYNRtBYPqawkb6eZ+10nP5m8xQEdUbO6WtThQOnodrrXfWsQTsI5ajsaFaOB
ko+Uszn9Cgbn8bl5uyAas21Q4xx05y699QSAP9jyfjDTYSuponEQhdqJaCjOt4UX
luffPAo4yXhxKK4LAto4k0BZJl2FBgXoyp3LbMlVrhb7jCG53U3a8Rtlcpl2u2NR
x/3D1cY+GAOsiKLlDSrorbNkiuj9WkMKWh+I8fOqS5GAR+OAEU+diTsmj8+nh2s/
AhFFTUxyR0L6p/9UAMS2iI7AdCynvBRj4/B+5LvHmJ0uMMyjuaOuoYsLe/epHoX2
xMwQ7X0/vpm4yMJADHk8guJJtBJuaEvD8TFFEPJHmqWFEDB+1DCRJyUq0EFWLVlO
DzePEvSTmEamEYN6A3yZIxAtMzAw9Zbf7Xj/4DKwFcZWm2fsHlvNnmsHH8Uz55x3
Zfk0lijwyFPBReoM1shkidMdyGVnVhyRX43Q8CeutXyBITOChR8CSkTXPl07EyEN
INkrqqIxuZFMK/DG8fOCxg3cwEjo9OVa0u22knbEHMu/L0DmzbCPlpsZGowoQIsZ
mjrqi7/o0VpXzqy/wJ/ikoBEaM7Mu+VKnhl0zngv/019qEB80bY+nrt3NaXxDqNY
rBy1umV8Q8XQIHak2Uww2oTdcP/eKb2l2fxLEJ5p+XWKgKs3oUp85o09hLCmVjec
/mfcu4SygcWWi+S0r+uB4bXbcVUI2srUt8J3qBXc/cJTgPT57m19adub1b07pIUG
VL7udGjMM9cF0hMz3bDmLLFPoLg5/B5sACaGUe+fac4b/uepZcAvKA7GtP4nKK5p
RmDKjtEOLKpknNkmb9luSl+ZMZSbuMeQ3NaA8xbA6CQyJVhXuN9ZVTClGSuqpdhH
f30ifRaN0gyWjx5djxGy7z9HhuZFUAIJjdxs3GRVB5KVibCjFt6c1TO2OdT7n+D9
JDVVeyzqwyb5x0eirqUBVW+8HwWZd80ODy2ZVdD7l8UrlIW1Wx6y0owWUCdkK8M0
5CooRefhSOnmeKzujH0+AlkXx8cg1wpaFG114Y4Abyb2APia1/EKqcUrqGxB5AMQ
SOOKGI3IogK6dSBcq1YGwgk4L/xchKOVpS0qFoBon6q41atHCHC+wr9hlyJaUYxK
rGrzPeYqELwSp9+obtfFq4cFWLglhkGdE00acGFzlG7Ot3dUnROsDT8AxMoLAygq
y9TY1NWDM08GwraT7x9vHs8W86lwiaa8dRdRICQcqM859L5oqYj4wWFf1ymYYDsw
nk+DYMigaZotmMEfC8DMyVRZw7zAsuWvnFarnYN0kPTtdKxTKqfNtb3KHQq1ef4o
b9ZXLPktRboxnBsar8o6L9JFitJQX+XLvdqNmEt4m5FaB9N5UNhv1q3Z/C7fM4Si
UV3nJ3u/x+AkCLFMCGvJC8hS6V6xKR8mcercR7ZAeJpb7M7oBXeUuyk0of3Lwr7Z
t3bjn90pImKRTcMsr9+rIqYj/AZ5QftGyBPMh6IxmRkf0Jjx9mD1IT6jFMQqeNPm
S2JEwLXX8YnC6BShXG3ShfAfD57EbDKvPWbOrHMqKmTKeoQO/2HvVE4LLav444ik
8h3f3MnzqJytq2oXiYbtGH5FuFRT5YS/RZCNFu21t6TtKD+tyHM2ot/Jm2CBog/F
lcsZnwPBkVcuRJefMNz73jROYgRPaOC/pacFn4jxreFyr5C9W34XGYqb55PZ5ihz
CgjZLiinzbraMNXjCmhr6PJD9seT+IV+I9mdagK5siv7fenzrijSpvGKm4UbVCIg
kBLP9lcWZU0OTUNt3cu7mGciQk5H8wIS0UAsJ7/EgEZO9P9g+BWdSdk3vQUvuppF
E0ncOWuw9JAWCTxGVl1T1w9/iSjObP4vn57NyQhjnhz86Zp18KtZJ30mNTIRx/WQ
KQLQm+yDTKcas26C2AKC63VOTd9xYA9w5gG1HynfB2COCkeo59Ps/jrOjr59UFh4
05naig9fIhqh66hHy8fMjruui4TRR64/XwbUmNevovkFQomtKRJQWKmow9HBVBW/
qSEHaA4vnZUH5Rv5f5ON5EPi6t1gn2IMMU50ajexdQ23aXx5Li0fQoxWsCt5s8TI
FPMLoQBh5UrJ8nZlbDiOzIKwWEbrbHI03mNn1A+SZrZMQOIFrt6v/fe+rwbSqAsd
GROWdpbTZ22QaxX7eMT98oUJ+8Lf3iz7S1DytguJiTOHamtQkA7pGmWoPJnJlDw7
R3MjTNCAHP4Eey4/dzRkm+Qp36qmhikkTLMnGAEB2AsojXwATlS7wyT575H7E28M
5cwd0Zvcdoqb+Zfdbr8gAGl+u3yDRuAP37y2e/V62+dC+Jtvgqzdn3/6yCCsl+FO
7HFiwJO1OndpXXqBXpvuTSGxhxy+RTHyaey06Ll6fRN0H2zPDyOy79V9SJnr+Ycu
2stsDI5KP/NlhOLLjKkv57uBOjRqY3THxw9wvIlvHK30SkCcNgFanRMMWEqLPbzO
+zb1ZSYswUvBPcWG/eW60iFTkxwDFY2Z+vrY8d8ZrRpMBUFsyBk6HVjnk3oJ+LWK
1XMhq+cn4nFoYnqBmLZmboPaNpjNlmHJWFw1zbjVYX9zDtenoWHP1CDZojCoB6PH
srW8vkMVq/gGxB+0sUNYPshhaCbZ6G1d+2nHFsB/RbWxZjELdmtOJZNDOKrLi4nJ
iLKHemWkExrKf6eauu1Crb5L4fniUN59KX6rFEKZxzVlOuwGD7v1vE7iS7XM/A/D
PENY0FRcXSVH4NdjvMiBgQPU0+nNtfCUqBxl0616t9MVCL00zpmfLQZi4hlur3EZ
ivpPTAhtgT1O8qdZlK0BfpCeHSItmWhFD8ImPoc/1Ak0Z2RUXqWYlkR+1K56hzpG
UXV4o6x2gdf5E7pBD9G0ewedy+e2gCBCZS6SaL9i2CQjSHVcEf9/85OaJgmV0q3I
wMe3a7UMXzf8O+7/GsVPe6qi3wxP3wRTe2Y7DfSd2UDIk7YTwlTZ5geS45kCwC8e
ltEuBcfygDqzeahbXvf5ba0Sr+k08CMznAJW8fqcAn+2+YqAc3YRuTXEI/YQpToU
CdlCWvYm4d3596FTd7iyX6t2f9yRMoWomgqxmFFSwMnKJVJK8RRpiu1a15554b4f
rjddFyD2NSJoQOPWf0h/hgqOVH5V+3yYdwN5Qw71cEUtq34qTgYRCM/4y1iyopgF
bjmGiwWB387E2+xy+/iv4FOvbpnZOEjnqv3p8NARKcgBNhXVabIidpeN5KgmQhSK
D7/b/KqU97iTecEwQsYSyhYPEdQUkcAyZEOU8/PAFNdf081nzxBVk1kJA7KmOY/Q
yz8BsJDXwTtmjUuhG8b9vAQ7luRjj9yuTiNE61azPbSmRTptKiNJGH5H4BNuwQVm
Si6CwGDZsL659qfqLF7AmFjO4Qigf2vuP7vXsuSxGPnjl2izVPxA2zxgvG9vKtnh
PSUVHjK0gjDb/4pykEzMyICBFcGEfN0SXeamQIKo8T02A9I7HsIgWByLYaxSg4q9
8WTV7MZNDx0BrnukYeRRnoD0StY9NHvSEdABg3WlD7gkp3mF8t6GtCVR7IGCGioI
64HjudVof4YZt4ge0A1TKffyzneY2AVvF0fhyI+WfzUHxJqLccCC2E34+QyJBz/0
UGTB2a0h3/tpIcBvPp7UBY2JCCYRF15SSqxDN7qGIuzWFH6nWD7SkpzZhIk2dRmG
ZLeHwkPbFz3IleZvqXxoIXGF76Qq7TVfxAePMF3A/e210fsjk60DEyqfu8UbwAAx
OUEkgNzuj/nl789rRakm76kH3ddPH+VB4rzoRDwKAxug7CUphRBcQsys6nRlq/ku
+mPmYiGdGh/Az2VW1qrVZpPopSuzyHQ212aI2q6y0dyQJQRzlJn9LTpyawPkMnN1
xlExExnzr//iAOtJ9aq7EVY5m13A+dWZyYeAW6Aet8ugySHXsKZTbWja2dHvTETY
p8SDggj1YXI3gORp8NsQs4S62nEcKGKm99CnCTbMyng5nUo1I1Qc/Y4MFcaQ/69q
Aiwde3SusWqxIIbS+mMRWCO5h7moSRQ54Kc0/yDcTM24f5fG4JrVRhXftkDPpvtP
7Wme6VOVxumhpGy1kTbErFKdXvazr4E8hfOy2s+yPmOAm2AnMkChGlZPm8juASod
T1RqhKTv0kyGSLE7RPAQIYceXTwKAE4Ij22eYZE29DCOnp5IE3jG8MpMplmMJCso
BQxu9RsGlItt6dXfX3Dffe9q/suS92Zn95IB6KQY14pWkzyzFkF6DV7kzp3khrKx
NnRWZ8D8u1hVvoXye4CvLy6UeZtgakA3PiZnMMw49EuOrLfuuksa8ezwgOkftCKc
CwdaCa48MPRCb7N5JezUCpiu1z7iV3sJqfR22LU3Sq4120Z0BkuQjVhvem0BN0Q1
fDeSxtg6T9HGoVbYOmmjtvXhKG3C8KlineUKkQVgQwWzUhCcBwB45/Bjw2HOqKxQ
vPh/pbb+DE4vHFbb50Vbedho9hvWC5DjCCTghii7e719enfLJmK2GH3Z1aeCRPbZ
NmMvHgLuABD8rgRSvAg4FTHFdV2LRJ5L852ZXzuWFi9gBbTOlObHDuBv+I8tz/sI
aJircbLrHospdwW+M3k2438pLQl3gESEygypFSpNk32zlH/ZRodZKs/nqb6qYY6A
7E9AwKiT/kA60BhFnLYiReX29gukqQUmQCa3qR5aTk722IJ/0wx6uwU7qg7nw8kR
kh/RNJ0U0h8nf2aEpG+J3DtQ9gcTJ6wckAHIy55Twy3Ddaqw3y8kdJlU7ZNSSn/Z
/CpPISpRR7cGWNskYnLbXg==
`pragma protect end_protected
