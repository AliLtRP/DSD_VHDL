// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
BghYLvFsuk3W4WdNBYETRqRjTMMLGY0a0SVL4HTdsM6ILpIL6MYTeHibb0i3XgNwJrP7daC+c2HX
RQKpy6Z6+Hh9Ls97bjnYetGTQk5nhfpG12kCvVZmnerBTAxrcQrLoQsaskgd5rlNP/AQkd7586LG
d3ovKXFCFPOxpWqAMqXBPawpZiqeBzBa0FQ4UgAjWaW+lQe4Olba/IYUD3WV8SUHmx1KEhiXiQ+3
7xmU7wo5bv4YB3XCrXHWkcxiyDULLQYSq2nrn6Q3Uv8/dSoPLTJw3lygtcAffLILSFq4wAYh2zwS
dUZuDpzuvFwJ3RtWMknNxgWempBQO+dO8uiDVA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
UYiwL4dRYPNw3aQwtoyKIr+JVCgbKyr0uPnES1hjmPCCDgNaUjzlcRhX2kPcFUqB2ONFFsF00TPg
GRuw90J/QDHBQIg3o+R/4qMA3K4F74aWwdMqHhCKPC9furO161R23ZxdhSWqqlSQsWIwzoiAKeCd
eXefINH3ha1G3Aq8dWYJ5UbbZSixwyYw87ermSvoC9P/D0fmSmn3lfIrHcyww9yJeupNemqCwYeK
KEkG/S11bwKG+HFZ9TdDw4NlqtVs3m9YrB5KD8yoqcJj257gSZtEOg3kLCX0sYwBYMeNrAf6iFqF
P7I39STrN5enGlEJs7+qeKDi0QbYY8EHbZVpEicFH2jSN3Wbck/gJ5X9SI9r5H035Zq4V//JymtZ
jkoKHpUVxPC4TA5FSbzROJy/eZP4bwjw5uanLo8Bc2+cuJ6ieYoB98ZX6pEuSAt6EstFdk3DAOYo
v6c5yZDNUMivESM11T17AhUpLRvo7uqSPaYs58CoV9DelendMWM3jaPpBbe7iEXDB4BhV2hyBzfr
oExDbzNHGKAogBvgDj+/Nj1YpJlMNVyMK24B67FFHjbATNy2eOLoEu5xw561lKAb3JMnxD7hmhFl
N47CXoa48evCBE1iTJaF4grfIYq4IIzPYtlOSNPqd95nEjaFRlQyHTXogAfoN5GSrm3gItS5GhHi
5jHRjWOvRBiKmyVgDb/zBC5kQWBUzimF3HY4KrCtAnGnPsmaPdDfoqIU4SOWxrbvScGCnU1RgBPl
K2CwxCX4l3J4MwV97MQg/41cywJ7AmXzBGX7B3BJmztfxHiu5mbztdNkrxumEnTQ/yuh0tTedAZa
W+Gbdu4cVZZq0Y46lsfhwmsx53Ghw1gupCKIBem+5i/9cXNTKCJzMg3kf1Mp/vtMXF0fXCIpEmw9
f2z467dZJN+1SxSAMGrG/WSEe4TrblQiSrVsQuEFmXt5aFmfvMClarUbMCcKfeNgCPni4VxzLom0
ncZJowzzWkshA+qK0f48cgOgoi5WVNgxhCP6CMjSE8TTiuiNOa3UlR5nhOHbfViv7aSjEoTynHNb
4fCWOEcDUHc0GmwGOsshgB1WVxutmukY++QwhpXLMeJ7LtGOm/TUj6gi9jiYDnMkiFopULNo4kfg
ua+A9ySnWZF0LC0f+R4+Iy1Opa9nyh9tDiexAgmtwxXV3/Y24FkBQ0GgqAOSNI/k3xZ0wLvOY4AI
/4fjdju999EncBVZRExORQdpDb8KhU8KZ1+YUQ9vBXpoSUP4uDpyEhcKY0gvucnk6bTRuky3wyBs
R3NFEln+ofMHhxMsUS6IhToOTsqSh5wqru8VsbQh34NDJ656QwzPVYcghlRaUc5jcY/m0/ZJHWid
Hfentsu4UYArwln/0wy7lwzcklhL5IvdZDwZ/9r8/4rDOSMyh6p0D/CEy8p3eDQNHH7yHvL6+wvn
aE3li5+eZBFynwvBqet7SQZvTxKIsty4+QJgBU26UctesuZkQFTIbezzIwtESK1dmouRwtJ248Y7
lBu6AG+dDB62k0tUVHDwF0EvYxy0+/8UwXA1DEAurgH0D7/qXxe/aZKNaEABls7Zug1UOjhqfqr/
DpJNMm8VZONXEeIAiIxSh7M1qFp3LSgoOj6pPt9V9m7h5lotWzXyOH4cW1vhd9FBinInAqtyPTLG
2E863WCY/9Fy8R6hHmFxWFgXHjPe7OeYW+f+TuU10ABcSB4xwfoMI9/Bn8wY8hwT92P/JHcNbdkc
455whZ1R9NkJzuI3q3Mr6pHRj9h9X9ua4OsQlME2WCD3/OZmqd8IeQvlfvrY4siLWkFWLvsokNpX
v1jB5/yxb7Kqqq9i6lxRjtJWHE1/ZjAPV9Xy/TVzZhA5eUvfKNgUuSOcO2YJvDdclU48W3/teS/f
hgCU69V6DyjonuJm+9UoDG3g6NoC95H81atv8HTS38pVR+p16njUdDELFhEQg0hxiYyaRBsLMWp6
MdBXvsRnVFSf2uDqbY30Ge7RFLXrVeRm0MCU0py99Rz6xjnnOPxoA7JmSP3cTqFqa5VhDCDkPQ/N
mxHdjuZSaH+qgYzIUFvoYjfJXud0DU0qkKlNFrVs0ZRArgNrSkGha8hEHDF5j1EmrlHlxtSBMb2C
pvvOKnMRdfT6wuffWSpHZTJCj1kuYh+6QQBdhB0bUOdWCaPQJGHHd3GtzYPDULKx6DbPkIXP+n3J
IZdbyehFd6+UCBHo7xCq0mqxgbFljUReeubeb7tNnCBCxppygFYm8qm+kv85bb8VPq7VdoSv9gG8
0/4L/fNJfT2oPcg4kp5n9XjAK/qQAZhcbTi6o055aC7pUWigcoP39jKp1jSP8XQUokhRBAPBi8cg
2pGsqzNbQDQhNTm0C/JbEaeefaiF59XAAY4yn4ZwRyGvfafjhca5TllXWAHmVPYWVGtj1tBx/fMB
20ot/luXDSqjEdasBrXZz7bj59hIGKUMMqc5ZZQ25lerOGqjImfPdyuHLIAf7dPUUkEVU1Erpajs
AmONC65o6IQhFNsf/knhiPGn+x1DBPiDVCXLOnAY24QCNY+4BWKgdzCs9yx4HvRzIEyjEi0hrKPo
8FkYdIrgP+odc5Q4z0NI+m3WwVe9plSMWeMBE5v+E3v/kd0B1RsVygOwrLBwwHTymH/A3Lt0Q734
XZZqD5+5dlVKp2fQWRpwdfGlE4xGqFQ3A6auZ6Mh9jt441mkG3RwP2XGZh3N5AxrrArYq5pHVLUr
0eXMmbBPiBbt/Dxi0SnxFC4Yz0D1tdhdEmBEx2OT9VEHZLawtg9erxUJn+m01zHDJhuhHONslrvv
532dtcL2iH8zfEHUtVFo0berBQd2WX9Q22iF4nIPaQ7hn9nC2qgfDS0YwBRRHdxfVqHNXtwjWsoj
3AFlPODiiknvwdCHqMx7eNCp3/qAb+WTu2mjbRv2Z8wOBok92VhkaOY3EYGIed4Dmkxl2JqaM2GQ
h9JQGl62YFFt3k86qEnW+M1lYLCikU4GTtAn59qHnpJ95g1f6ZGt6319WhNPK+vv8TTKAnlynbt8
+BZFYMM1sMBO9NamvMjG5SOCAZrmSwc0ozIg8JReTq8EaDG2cxHgCqFQ/ZwpyRr4TgOX1jqgrhcO
LWnBuDNE0wcYgnUYpXk+H8nTlUn/vJwmcdZNNcRFlzpy1yqxdSw6fdBZvzbDyxIOoWShpuJpVX5+
LiIjl28f88X59jw23tKInR2D1RMYMUOGLTRUvzFUTThOJoxDLCX7VeUUbg2mXUEZqdO67lkqHpmG
XG4Tuxmv24ctAXS6V9u3SyTyD7CHNKk9gaHhWy4j4ZQbvX+eC/sSrsB4haNqKf3qiIUhg4wX7sbh
yzJEBIK/YOFnbnelphD8dO0xIkgGrx8YOs8npXMVSC5p4QqmOeeJkmA0MiWkhwgpGrKIC4Z59MB0
W+iBa75tVHY4QattErREOZZWpeDAZF2OiCvI0WZoUfz2D43msnEc2Moy+dji2LSE/kNhGnunq9l3
wRp4fwmyD9XOxg1f0Yb0EEr+DVEPzo01zK8GYoebS/Q8Jq2IC5txBchlRo+TZJuukt/JJPPUgqzg
fXlWFPcGX1HtUY0e/qjiSRNH8sJoCByKJMlD6OvJcPBmxq+A6Z47fWF547Kuz5SAeVx/vbFgnG7+
rNFP/G+NCPEC2IvxEi5UhgCBUDuMGdGwJB4u3oOtm2MUYR/Ck90ls3ZM619SIFaaAz+auc1fwNpy
UqYNr297xqMroFteyNSpSoeEtKJ6TpJ+EuJ7MumRzrm2tcuupcSAr/JBdMMR2jGm8NKoP5mRli/S
7gYibNLrLb3e8wuX+HUvqnHd/vqt6jq513IxIveGn51+lK4zRHH7/bvWTz5DlyBL3NF0SqWuVXDV
XPPn4REk9/YV2vTPUEf9/fSO5IGX1seCy/07biNyfctWvNinXuZxWM+qicSDZAw3Iy6+uqla1B9z
FM56qLSvDYEoF2kVGVdKqgIbC0Hswr8izSEonKARLsIjg9YL6UbApciVIGZ5vAKixQ+8pwXP1jRZ
sUg/nYfe42hJW+6aNKtAdADFcDKBwtyVcq42iQ5V+lmYa5Di/02Dvg+ubc1hFfQt28qzRZhTNU7S
1Dx0DQkxISToMDfCNCj4ct5ustw6HyS6Ff7sc1AMtocE6G3ytl16CE0NiGUKa/YRIoQ85bGz/sJQ
0deTGBNZ5j+lSYBM2tvA48gcdRrsD6S++QyXWyEyTs/4r1DvVQCeqwJZFklIoqrp1qQr/mkYf5NU
rUF07MOJLuuGyqeF2CUkJg70PkoY46r03kdHo+ILPUXtF4KWmohBxpIQWwsQpc59HGnjRuSVIREB
TY9yPInhX/eZVXGgRs9XZrd0Zo/+9qmyQGxV/8vqOZjXODjnHAwUFGUz71EiJ7EG12jBTcttVuvJ
yZgKxFG1a+s7I66q4iyNSNCN+YzKEtc/kduhqKsZGM9Yiz9dXGPsxSoGKL+iTKFotSkvTxGh0mve
e18SLS89u48wfpD3YvjwmWZddWaEUvirw9viDB0X61IaQUQBxBW4xBpNjkr6UFTLw4jndYt+d6wM
ZRFw3cINRlZDyrU2zO0FzmSDo1XHpvPR2Lhf80fmgpHAJwkIPdtRnwV8erSNTFD+ve8PUhL9uRIS
avM+8dtuQfGyuvvHAuZAHywWUAIyCeqyu614D8qghIs42Zig4aHuFqi5e+HY6re4PrLG04+KwUS5
KghchHQD51QsKKe7DTcNr1568KSx2EgbyNWqsz5ZU1YNibD42uvPwuWhLwECfJD8D3eY+RDJupJ0
dCA2RFv8jlYo+hTaRb6HrfFg1q7hkoA7GEUbU7bkZmENgNN1d8xIfh44Onr27msiNlhAvQeMKyF6
mVMp1afxrRW4C6jQgI7/d4pUbls6bN+ASpp5UDekBbpF9leaYJf+z51FAVEgzojBtb0VGS7492MB
Rcb48Ps0wEp+85nS58jv57fXh+WcEmyRwmhSdmpdDAHS6WzqwO8O1glRo07kwGrsMXfuWWaCYNjg
NXBfN+Sg25wKFBv9Hw73rquA9XCu3I2+KXaX3Vzn5HICa1GncR4umkzk40itkmUz9GB3JZJ/cg4W
xnYF0RTEvt25pSVbSOuUtAaTeb0ePeyC/w0CwwbOjd7Tgq/hdjhN0wWtMx6qJIe2wZGpOPG88e2u
9UVgEtwWFmRK2WxtFll4RHYqQ92N8Y3IrpHe6yW2h8m9doeYkqN77rgpG2FeYt8vx8FViAnezlwX
xOYjXl86l/d0pYiOSIIxyudPJ1XYIVsph3jqkl45IG8BodXkRKB9mBbTdnwyCe+BRL6UMuu8kbR6
dyC0vBpVMq+MkuvFXumqzVlmcMYg33XXBRogpfDr1NpTCeJhtgb2L62fkREWhlsP3uAmcVUZ/uiS
TEUnx6KuVJjF1p66760JP4g2iiNqvTFx2AcVhL27oLEArTV+KhvKeQCAbhEkO7PBRgK/yaReCDdA
XqLGRqy5aiVjXjAv73GnqIhr1F+3L0Xiha3D20AgdP/GK/jQfwAEWxgHOrBTJQNJYJyz7J7+OW/f
Tz92/9A78YjG0HJNHqpSc5TCYueScYqtkNa0z46eSn0MVt8lhbsDYkUpSOBwtZ/x0Um1D/b24+do
pQAyy9+7iqXHyq3tgR/YCpHuPNsGBzTM01+04JX6Dk7enDfbM0j44VpYXSFfCsGaMx8lLD/a+sUP
WoQZxtkyMCF2cN5nsW4gc7xQd1kQGJeOEGcLrRMDYlYwZiGLB7Ad6NBYt8Qh5tmtEY+yKzaWZyRb
s1AY19tAJBq3ESMiAwB7N8+jzYUDxr5lTgHc/dgrvpAIJEMvIvw9biar1ncamANZ9GtUEHs2JBcM
MGyWvQ9s7e6hRqEz1nkIRPyGBCrcdly4Mwn33MeWu9ako4SHPH+RRkKFoPp7n7H8635mA51o9Ref
zcfBbr0ON9dL/i/c08lKB1o4fO182Neq75ECDm5T5x+ThlSp0A1Oog7Fxzs6hAjnc6xznPL7MhbS
9z4MBK4Nbq8jSQG02A1nSYgW7a6RxC1wLt/9l9Ei1tzIMSOl8mxRu8LtFdq/sPecmaMlV3B96Ngi
hLHTgPBE7GYDlk6MF49gfUxbLcNNKY2PLZRnrtGnxEZjMg53TijCqI8rBynKaS3e1etqLilft3bS
8R3VammW4naoGySfCUXkcCYetLv0aSTDCMiBEXJWXH5jh2CUNFS15VQzxDldmcZ9DeTnVfDXKIF2
lrHrsuLnS4totKQEaixbCRyZuN6+T6+QqV60ArGG9eTGAaAzszOPrqhNzFJY0nIkCNWq1oIw4pD4
F2YXfV57fwH70KYEH4xLpaYuehhaHnb2WRSdINMdAQ47FMgyX73L+SSqKtOQN9NPkrbJFZp3VcJ8
IiYQcmb0vrkEdsQfD89lPTvuAV6lha2fihtCBMhJ4S5Su0m33H0oUgQr8yGF9oCqRG3PkN+1Zmtt
y2aC6HujhxdRMq/ItxhAZgrKOjph/sgQOmtEro8mxAYzIl2vfncivcz4a7Z+WRtihp7ixSDe3fSZ
Ew+Z2IvbL7mOX7xPEhW0uHqdMn5MPo9fpbqyViYOec0UYPHLodKC/5rv/bM0GyFXtz/+QMlCj8n2
+kDcx4ORr4kQsz7MbN3sgZproKDpKVs7nfVp0u0a4O1vpsjbviwPQgDLhAY4JiAgQr8eT8ld2GKK
F4nlHJRbZc3v/KrsqQxBlI5oVvAt2zgJ7PAR4N7uNkfl+0+JixHpGs26SR1qB5L49UvdJEtgZ+X8
uZI4fr8127NmW56GKvGlEIFmgubM/t6SRNVS4g03BoOOv1cYR7KLgmJnxYD6Rb+KH08kB7y1ZCEC
Ub2ssxtVy0S8zZqhQGFRw6PkX/knETPAmzU7eb6+LRywAugVVaKkDCZsPiKBQ98uc9efI3QRbqdK
uLyzhuUJEYNxC3o5I11RUflv/WbpyKaaVRRK2u5QMkxeTXmIuTLKZmQnJHD0o2VXL2PUzsoIkemE
3zPPThzyhLI6vLcoL44ZADOSowFcktgMDsvhTNsyuJBZDSAa9HWOiVj0xf2GkNPNQUBDgIMkYKt1
d9uAj2gPWaTKGlwrRd9GNp8IWV33cjlqko5j4KOPs6NtHoWngyWKoyqn0gTi1uNmDHNEJe8VUJ5H
Pgig26oNwnBowy6Y6yN9wCNr7wrSmhccVZSjuHxfwh0mHiGAQHPeLpLQOYVtLwQi8dJlqRiZOkJz
O1iDcB1FhZS0WI4c8hb1uY5ymCTNwIFhgqkscEEz3WSgz2bOT4lj8uyvCPIr5UYf8hL+heLNgl7d
kmsXyw5Zd50TYbmDBWWzROn/HgP9O9NwWXdfIqCx10d2TumKHV6KRZDpqvbk3SaOvfzGIZLChsOl
kOSx6UuOOQzwmF9ByttrqVk09grgwyeL5eAKOgirMQBbhHCjYcT3zuWuxcCbLcAVDNO32s9MCPw0
PR3Y05izLIBsyJmx2oj36YCRQHtKDgADytUJcDS8lkIaRnm507X+0vF43nE/QF6kG9VMw0gCCKE+
QIF1NrebfHdtSL8Gvv7mte1JfFbZLZmWYIv16tQDj6QJcjaB9UWJyEJDDa0PXLvbg/PZuz9wj7rd
lhbeazRdgRKetCcXYEyRhW7bFbV6mwLhMTfsNQgcjR2wQkA3bQL9nUg/Nv/alBVEw+4cngShr4OM
CVK3uuJM+bjw1cqVOEJpWNKeP/2D15sJ+kCSACPXDx0J8RJNp/uh5Nne6XN1iU/Kx5FtgTKmF1m5
JfDkTYn5qU5nz/jXIEhD2K4mRw3+e8X76NK50pdSF6Bo2TDxdmD9NXVHjoZb/ca2qRIhvo53ov7Y
svZf2d6pMx4nTqBC0LBo9xchRapHZyddjUocOzK95RDZkR56bOuNety4N5cLLd0VomJvt+bsTaTf
HVI4uk+OZwRdCpIa9cOaaikIeCeWR07/+pPZ7i3JzuxOa3L0a4B/PO3jRCwwloCvQt1WC8ZtuwAk
yvOaPR9Yw0An9k6A7J4i4hd8xsZwnzvrABzWzkBdFTjGB5uBdnKhvPIXDiaMeCjKstpMrRFiAjBi
Y4DBYLRArRn7WafmYm8EGAwO3DS+ZlM6/sXauiZxhCgsRD+Ed7Fq2k0qj8UbHXj/f+GRzJoWmaKa
+gpBDDYu7Rpk1+tAlCZW6LGdw8lEXL0DADdXKmsCY4SbpJewmobk0He2M2gyGdxRu20o8RwcC3o7
bphi6+sW9flXExku+GLffX0AJ76ALs8j9esm2xSexLsjqm6J94IaRcEOs70N+HP2cYWfr5toQ6h9
/b58OrWXQod4b4fuxrZj6g4H/hUk7KtDy/WhxRljtXOamFV6OlJmfIG80Jj80A4dS0zZm0YySZw/
mUBY/tG8O8plMn0ZqCGAa8aPa9wDYtms6ng9q2cMuFaMi4OugRpdVObuCPVZSjm/0LFNVGOq5C/K
FRTNoJQQPlMdUkn0tkuHgCvjuhJT1aRxKBKY41fEci2y6LepMYyTvoyv3KMJr+IDW7/FRszgmjTT
k4fg7TsgPF7v0vKISCRLAaHWx3KtdRJ31of1RxEV+1DEVcU4cR6wI1yXm67CtbqmwF+iMQ+9/CBB
/8I5IcSWoTITaIYTI2yX3j03/ladZsrHbYDyHu00/u5xbxTt+Uv0//6JVEV3Xj8mtIDZNK5v9o4+
XQfnnXqrGm9jSyGnuxjwdJEwBCK6WxrlL1E9j+b3zJFcKcg/9yh6R6Zx1xzhmcT3bMxmadc3Uga6
8Q37bajx00vjql4980ziSKyAR1jmqmtHIzugDh4PGznOxfIOiLXPUMUQopTFr3+lVzilpyZ9cier
5u0+QfGpcKWtTdtlAADy5cuyMvJ5ywLpTrGDemaaF43P0wHOKI1gArKCTiD2/UtvBfg253CfWoGg
rtsxCnHm9JRcjmHRG8ev17RQMK9ITJOuqAbUoTt9KyoOKpG7BEWoX30TvDSU9DIXXWIPwobDHfGa
LcQwO6EM3g/1mu+ifQ9cvxKlYexaU5Sy4TbcSWRz7nDtyK5p4+6ygZiUS+MfmoYjIewJAGnAvGFd
sBi+6vQEq9Qxnh1NM5Qu87fCzJWnUhiTuo3zbghLk49b15qKgrUrtK1R3Ylyq0dPsR+9Mf3WDTK3
XPhikNF66rcAduV9W0/tdmuuStk3eHjmu+TlbUIQRpF7uqvApE0Jdj8BzHkQ9f2SO7mpH2N3YIrR
7Wa8rFC2Dn2psk/MUioceclBrwNPG3s6HGoJAH5jDcjPfro1Ulw+M4RL188oJWqTRORqd68ibHXF
3ZojvXxB52RJWI2ABmJYtNjL+ytWOSjs48aTtxsBrvTFELuCgp8PY8RCHbxdz8rJvbX5Lk7j5XxJ
Zm0uPsETo1VBoerdBG7f+ijPSvB7dVlLad+ZM55hRD5ATQjQ4lE3muphyqif7fbD4Pwwk9t/5Xut
IAIhiHENhGywqiDkJARAsstfkbvTPwTCgyfhKfS82JUgzb97wvMIjaZe9jawnQAhLpDew1rnuo4W
4D+433338XVqnZwCwyO9TbM6YVTPJBV0nxRT1bGkn6Wydd1a2nXtAdT54xz2/P+2LzZ1iktLnzDf
9UQ25LbBN1g3LqJnPdmbhOoNm8Gve4RFCUhRJE/jLaBy9wr4aIaq9C3kne4lVX0dvCqR0gAtznMJ
+g3VXyGBqzlarVBJGIyQF129eqTsyDOKBbVEZDanR3IxVFviS0XVqnIfDXPWO/ue9dtcmcwjCPJL
lfQ3mBXjQAxk+uzjUQMGMYzMsW6/G+ZPu0w2E5lijkt1fPwfgsYMgGjbzAo5hnUdgd6R+yGrXIK0
8mZG8jQrqXmTjIsHvnow/+tKJlng9zKymRImfQN4uO/BMbEWCozGJtgG6OPL5YwVj3XlW+0izBP8
bSQrwml0ci1eJK9lL6VlGBxjPyXECbv3LCSY7Uz7knKFpJDzS0RqnCyM+jmJeSjY9dREUwO6q6KJ
QhjqE5xINLaht6FGcnyTB43skYT30IUjfXfeaxmWP3umDfnji/wnZjtN1XPF7ivsDIjQuP/ENQ99
JHD7Zv+F+9hbkoutXdoHNj7u5qKLqoL9c3ctRATZ2He7BIXbH7TPVkwB4pmkSIPDp4oqIveePq83
qa2Yyh/e2rohkHziP+aKSGw2Q6kANtBqBtB1hTICpsIH4j0yENnXUYFHm/UP4pYPII2fObfyqDh8
Vd0w0pGpKxml+x6hkwiGH8xBh/K8rzTcl6Q/rSQDXWc9oYCA2TbLg9THKpaMKKnzCfrpw/8EDGie
VAHn5l/ClK2nbS9fB+OEwbhzvT9zjvnLJNHii0jTLmUHPzPM33lxH73NZg2zaXiRzO3LokwCRAqA
+ogua0WseydR+6oDEGW1KYOec54sENrgfbsVze8ey1YNB8YUxqh+Tp9W+g2d7JkVBf9GdbCMUAVC
7Qefj0pBBYBSYToL4Id7Hf8LbtByDijglj8F2e8wfn7z2X2mj3+mHgBICgp/CMhKhyS0Jlyv6mJx
3MnW4QNHBxcFYs+h3OpDjH052nW5plpFe7003XAGxczyx8rolt8CXN3bMOzhXZhoaN0qZemZs0MX
CKEVQULfyaFhVI7njPO1X32eaqxwtpcUqlsbHLZ0bJV33LKTu85bLG5I+P244amW9hxl8+QC8mwU
qcHbLtvRYDZRfB/E6bwUd9elSaA7vtPnSQoQ352N0V/J8ol12S7pK+vniYC4ZKbI6Eyr8ZLfY1U/
1d3c/a6qXJEXMfAT033KIyBhD5Kiio952mQRbFSc5BtfwUTnVCYFpu0CFdRpzwl1hL214A1BxIXS
neC0F3YcDWHhlC41cs9bBP0IhBid0+KA4mbC5zySGtOIj+uRYSRhWCsr4QGq3UaRB+4TKvcC/+1u
gp+LSGLGCeSVYqOaCUVj2454we3LCH/IgcHuCWScfbgIQ0kY7JKde7aNstysaCn651Nr6ox7PrjF
x+hcN8216O23A+ScLZnqkdjrN1cP/vPam8FJz6ubarnbyiqrp1pBNCjK7QXVJsMVxHOn149SPawL
n0H09W3us5pIu3TlMCZX7Kx3Mn7Zm587Eh/vuzzPkVXenSRyaBZBTsQuQ5sNB5YHdKAE1lWHljx+
A2aBUiTh0P88hNECvVHdU58zSotkOIDWIHALaPQSvX/9GrEXQkfNOT8Q9ziQh5CuxKmthAlYvyBR
iLbs/V1o6b3wK566Dm5ouEWuu8mvDVajxRgC9pW6R/XKCJd8Emt297kcEsTILTW0O4K65iBJrO72
Zj078dHZzIkwRZZqVZdqqls8kwbkX68T4nA8Vmc/4XukMVTmghHur89yz9xmKtwAeDpLYtwUZjla
+l9EUxz1FtfFkPe3BgE8NBQa6M7eI8ko4jYwip09aTGBQoNdefA+nSlEysGEctWvQTJGAUhmWpGU
GBNyx4HkmlQEmIIzgLyX1s1GByOzE03eYA54vwVL3NLbcyq5d4c5zvKTmgZhBuTKyEx1GVJ2mY/v
0Usd7wyhqvkfpPgQlSyB1ByqPAWjJf7coNaJlMDq5b0QnpjLFXMGxj7B1hIx17vd4/Vmpgbnx62j
Ck781+1PL+d3XIYpnVa6i93guzzN58b97idb74NJ03haC4Fpk08lQfQUVu9i6XNhIOM4H7WxG+Mf
ExqA3QhAOSjaPWXWopFOn/SRTLJ0CdY+LlT8jcOz/4z6vCOuq/L+dZck1C0+nyKCLHsVHEvLCn5s
CM3EoBtZ8zOTZaCJOhQ3LJTZVkmN2DhphUVSXk8DBTfETfs2eZyWibl/MzVkp9WnJNhnnPneQUMg
fRPlUUJzN8iWDh2OL9+pmGtUvhylVfajlLB+j5cfFhiQ7eJk9K/QYPpvF5Nchi10vR4o7rEwwzYn
Ne17bEFkM8naLB3yUsfgJpVqooCbhocIgr8ZbBKFTRFYZtFlvQPqRt6lIYj+jUDLslYYwR8h4Jrn
XN2FCVrbbVHewttqXb/jT3ef4KhkK7BbIgS9t7c6iuFOb7z4v+hoq3Cs10CJri/5ZRCWflkqE922
Svjse1UEDh6siHk5wo6Zj6y4SjGgZSDrj7nfRX2OX2rE+f27Dnyit+n5rtnnb6YKrwSlKTJ8CTt2
DsINqoVeaUK9Bqztnp3ETVQpOy3jpWVyTRNuKVWPccqcQybQrVDNJP4Ee0gUyl+qeZSlmE7/pDuA
rtZwkQSPdrx5B9x3VJARPQTWc0uTmVRNQNeQUZEUjL1scCsG59HTOYPl54D9UtnTg7sXLCX2Zqtk
phBINP33rgnzrfvi/1W6RLVY64oJhKB0D2kxTBbf4OtIYbgxgXEQudC5S3s4igIhtAfug2yAeLy4
Aqm+hjSLI7SsKNbRodTZY7V/f+DKUJWnWJqZmAPQGnaSOP2KyQx1H49Yclv39GqGWWres/7sn8Z1
yK7GoRb4ArzxnMGBFoaWN7tLwq9YDr3PILborp8AE6wLEOnFHnZJlhVKxcR1hvVYJtuer4M=
`pragma protect end_protected
