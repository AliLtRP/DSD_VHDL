// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:28 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ub6i9bv5PByciHO08F8D8ZiWxIPvQfjH+Sg+BlWxU7fRdkNjaegxHgFD4vrlJhFY
inWC5e1CxbTuR60IDQpyrr2Nsl5XzPjo+2Yvl5mUJ/lbicxTK+xFA+FTQK4lLxPB
rpLRYm9x0ixMOcFF8bh/tJ01XnH0GBUky3RkK8/TjcE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5808)
t2wjY66p7Z3UH9oqP3opt8N1ZzDKsBcKlrHx1zH4xqNX06KReNbsLv/j6ZqP+t6I
Cl0AvTbkk12JCYRGQFr07ARfe2HUU1N9BBR1CO3Flr02/hreAjA3iZWou6Fn1ENK
ToJZu+bKDu0oNXUpT0DFiD5s2nSfgJUYgbeV8VnO8Mb+Qssw/g3Wq739MuFOb9mH
ocxEpmlf1bTqRKPUt2k7B5JMB3doMd+AXth7rxFv9WcTF90jKJL0+br9PKEW1Fcj
r9sOb7emhV5KO4CYGlcEtuaN70kKjqg0pYV0AiWHVoudeuyzqjaD8Mz7O0kZ7bsI
SlEhBxDZU/K+OevNQmsDbJxWhs+0guVG93cFUF1Igr9jwjVSKf8BRBEg3UJJI8BY
/f/aAitl6+797vrVWHx1Coui4hoyF6LOEv9dn2zDhzHemaKBnbwpO3Md7qs1DsWr
7O2O2w7Gv9zMFHUvI8q4X8vO2+dz07pI1OLSvIi6Bv3OIOrgq3lpKPGCvwQi0+VP
GQ3+ap48Y8WBTPECvH+QCcXDCsITYHoPesBAf1XNRDc721lCA/qdq2TtkSofmQtt
iiMOpUKDH6ROhQVNloqOCnW0NuQDDm6c7hVkPsZdSi+Orxv1oHVTvhRRpFmVA3L2
OEYOW8m3ysR0E+FDvvzNsTXIt4UPfwtBjaCTR7itJh0FcIxNh+B71ChkHJlPItZz
DLYV04hsZ+qtkzj5on/wjRs3yikjNsqrEW7y4iujUsB/FKhWFGc2ssFkeS0GdkpM
wZVvwQrhPx/XP4EJCGNnJQOTltdwj3D4e9yKXXCJEeZc94rmLKRVynjAtqu71aQH
2q8z/y1JeSIMxRWVyqOfKnLKOOdtHCT49kOktkEI5H9oRjXs5h32eUt0aNt2R3ww
LVZfElEPuXAf20ViS3r7vLSJQPMJK0PbwO+PGB2EkbZRwxGesi/UbYKGk+uqOkuz
AvLSfL4dhlfsAfgQXpvIDz2m5Bt/2UsCbeAdZCUO2Ri5fD2nfjAlABdRs/b3qWnc
5Q5H4NgeguvoXa5h7SV5Iy7QX4i6KK6+9j0b0mf0iKgU/u+Kb8jDYyLlD422bBk6
QDAezTlOq2oNNPT0T5UtpY+T73Iy/NcXq/wm9YsQdfCjv9dFC5OH2S/+cyml5BE+
p0X3Irft8JcY8NNwRkqhWLhzBlfJgCK44muKmvu1nqwCjmDOTVCtvl7qxgcj7MRX
fH5EOGMwWZ5ewJ8tl3guWqDOWBndaL1Wdnvdr2Wx8YF98K8TcZ7mvgaMQzBoxtcC
r1h9ng7hvEb2PZWtqJTqCHD+/xuKxfT9xyv/rHDnkNamWSwDaRXtfpaWyMJJVbbv
REj4yk/J2e2IyxsEhk5P3wU87WoHpWHEfIGPSb6Ob2GY8BmfIhJ4DA3q98ynV/MF
KvWiENe4RFjbONxDMmbt999n3+q5hsgVh3BhXWC0qY9kqpVrJHNEfEst/rg3H3oX
H73c5GpUYLhPxQPLTGO9QzKxSpMM3w08C/gjTd70tLEg0qLRCqXD+nlTx4sp2k8g
GSSNIdx3prdh0H2i0HYcwqrlzOyRYQ14EAxva6DHLZ+5svRJ5JcFqAwgdLKSksy+
r9i2Y6hwt39a9r9OWl/TOLV29umFO3AaUwoBdLqALGUsV4lO4M5b9Cfurlz9yL8P
KFuEEIjnUWRN5SaUsVQinvrAfyL5jgZg5lljbmoBsup0VbRiOmOd3nuWbJeQ9aDx
P4uf/R/2yPAOOVkqAtBuwoEAjn5UGgmNw/D+xZxO+HINUara5ih+9UnBHTxRKm8K
36lcvT32Z4tmQXdOo7B66aNqJ0Uv63RGkVO2zXkYte3sVVRwpiIWuMRztPEol+v6
2O7nqIfSsSt/BNo53C121gXLK76h5JezVWKUqPbAAYJnf+Q1+VtP1+NaEmd4SFO5
T346nB7ZMTCw8V7EvIz4Hq/7Phi6MySY0z4o+GaDHz0Vpcu9DjGkbgiWLbarxWx8
PLJaccAMAQArrcbO5TNUMjICVBZWVYh6A3azSSJXl3+bDhlQdIo8lMCs745W3k5m
NQPRURkidIFyxfX2ffWSbikB4LHWj14UnqVsjXC0XYCh82QrLUIYd82eyiq1Gfq8
Ev8cmPneb1LLc+V7hVuuQzQjFPNQmFrJ47j8HAx0TBOWIx4w0gbgA1GxaFSav1nj
EZbUjC/5tPrjPCVwwXoZx5lc9scPCTuk6jcs59iNFxGe5JEk6O/L6LDSPj26JUMH
BOAS9/YZEC2PVSD9d4NvOjnljr2yRUbwX/eK/Y3IMxkp2Se6jyolgXD3EthAf9PB
N+pyGwTDDMvGEWSg0dbg0wOi4v246KqrVqz+Uj4JuYDrxG3X681jxtThF2PeNTOa
IlJFON0yj7swyaVePNqvHbYJrRBTGBe64nnCTJ66sOi1JiU2Bt1DQdrmznKMu8Jw
KfZsimvUNxaDDJYNuEZoGPA+y0q5CrGfUbmODR5Hqnf9DFzYsqxL6Ny42abeWIOQ
OpYCG6MxvxRO9vWUfpfKNbS4X9Aqznq6aRzc24SV3qzsU1JhrhOpkW9W+Dckdj59
XouP7D5+CTr9fZoqCq2Dt3i2UIag7zw2gk2YMfAajwxXQMeXS4MQObrJEPstC5D8
/XsaFqQb2TwcmH2o/B/lDI4QLJ5rP4qOFZytcBv/BhGWoJadQed8QekibuqFmMMc
i3RmtfZOJ+5JcgCV1tsBF7MqBbcGRALFjQ4JRWbcIB9sr+p1aSZxkVu4/oVGe/mu
9s8SvHS2glKXojlr39fOUxF461KDjjD4FnCG/Bhqj3VysbFM4fgvSA7xH1U1wJ7A
Gaib7qGCYV973Q4vUM0iXWELK8ayoytS+1VBQK5m4iiFAFZ/K/+3Fj7nLr1fmlKe
x7iWLY/G53vzorJ61swhs9lj9cCBTy/XrAu0hg+YyWzDWWY+o7+YaTK9MGhkG+WX
zqZ0RNLbgNRSXEa4JjdsZ+O8sZIxOXPwZGjC8J6I8ZDfNvThcGEH2i1gi7LoZBPf
mDz1G4mNEp0mqK3V33jvuujpEZZbizNfrXt+Dguu5SLvQ5G6d2pkOxC5FKvMZnLW
jYadCBmIIoR56RioZkLHmE0nDA3+DQ+NkB+qecglqVjvjIiGnc0ZZW9BYm7rM0TC
VaXab9XEGSbvukgeHdlpINErigO+JE/bXpP4Yad+Rzc5e4Wlufse3qD+zQJhg3vn
lIo4tX+AIX381tWfYFViIAZhcBHQ5Ewrt85f3y3SNDxJ73l3hn7KVC1/7Ehg8Rya
xG3YtMPgZPmBmmL52si6y22vmNpSFX/trCLsjF8hUBdmFULqFG7MQwbLBdZcrFDg
xVcFnVTF+ryI2Qudz+E27rg6HY3Th8bE9iVXeg9u1sk/lfr9BNjORL7vqqe+BbVR
0u2IWtAPVilvgJQ2uihSym5BcdlT6T5JUvZJgqa/2h1uvlqldKJb/3GMYBnwZ2Bm
l1t1gXD9Y+Nnxta/8f9LerJKgMQ46Y2s0f/J1U7WmUw4MOjuaBNcj9LNkO3+CD0P
AgUr6mDfEhUI+4PBveJCNFfEOaJun172j4iGG7SXPzhzN48NDT76+TFk8Rp0ibV+
f4dMX2Cx8R94r3v1V3u/nQlw+uK4nBew8rA7iUVc0YAJUTEUGzJsmaI5QPOo5DEK
GX8hAwRMb6try6ErOwtn2DTC0fsIIVFXCdKhJMZpm+JnO1SM9yhOpOMPWh7WLT3s
0dA8y48D1xDel9q+VUb7d6cZJ1rnzJL0aD18UWFYif/KjPuU9duMm1IYG/e49NQm
lGYJJ+7XspXkY5gV8niLysA748YRR8D9VNKqbKPj46KOeQNJJdnOQ77J3VZY2YYm
7MzRQbcmWDJp1kHxXqUKQJz3b53EkWAZKg1lbe+Dd/YPOR9oR1xnZaN4cIl3PTvg
4EVMhk+8N3Mxl5mC6UtAXISiVkh3AzMaVHwmOOsqXy3aEZgq97xPpyQPWJZdtT1T
UvYMAKMweQbW13nDoSJ/01aCXGauz+MHB0SYR6uy1Y3TuNRBlbYkvhE2LkG+/pj9
wp4bZixMG76WnBd36VuDBUn2nt56XD9JUbBCOKEBuALaIGMXuMbUh9YySx5GieY+
oX1zcIKldoa3kEOSVFAUR3vYDAbM/e/O6Hmqda3UTp3AQFu01wUDHWrUWmvmZT2t
mW+pH4GxCgpakzJbTPUt4XSrfaG6HHPs+XkHdw/XkLTFiOcWiHTUAcP8XOMN3mzB
Hxkluxg0/jXyvWLmZ3tVhKaRmQ0lwbxLuIkhbemOEtBwRjNRyyL3VulQEJnizFbi
FyJ1MGxKD0Xinc4JqxeZ/GjJ2Im0uIcEzxKGzNsxjaOq8OPPFwsrPp8uBZXVzrQB
UHVfOXZAANcGmLnK1R/3SWV/v5NYt3VOmQAmXtMhX1Ch+PpgS7GTvwdRuQtpLMD7
DBtdbMA3juN+m/jaf4uCitgqgM+bpNq09NGeDj27cqfWoj3rLHrAC5wXIsyWzBS4
r0nbbShdBXwbIToqqwAC3koTHTwDQy3dsDWqwFrfoFPbLwfQAnmI2sELXE0BM94+
p32PRcbk/9PsWK/Nx3wr4phOhc491IjWBSYuCUEc8cAMS0GRRzWwNeFTyddC522J
YUCRaDefojENAY2r0h3dML1Py0yVB/ZVchUfMIrB0tsafrEjDLke2AXFcXLNx/1x
4OJN5aaxa6BT6hKXm8g3Tw3bjRZ9V5OvJoMsXxc/S6zSo206s/uwAnlnJnPg46VE
Y+oMMGE/cbBubFIhNaNysUuF1x6d8FvYk4T0LO66ITP7yqDR6xQnnIyHQkq/UrEa
gT8bHmzIMshvrwliW/0EXVpb1nLkQqsjuwMiDi9f+a0LYDUlHi4RClhrjY1UtgYJ
9U3Nw8zlkL3XMwF6dNWa9EwcZ7R2Iy4YTAI0y0RLXBnyxbCn+S/3htVS2XGzkXwz
edzzRN4SwBIkoPIJA3zQ/QMgaOIDpefHRXKqSKRo9UNjux2UoSe4lXurBnUJJ+IT
4x6IV+l3W/fYKf7qh6vN3mP84lBbVngNaT7D+lkwa/12V6CH7YBycSgPaol965SQ
r6ZrIP6si/EQkHGaRe8HKbi6tu1VU684aYQESfMx+WlRCgiTrM9P6Aa8jt5uu4sr
6mDpfCguacTRs6Bynf3igtgQgZUa6PNvRcURdquhqyZCMI4nSRKDi3VTtYmKuSYH
r9ujBmePMN4w+tIucoLOOxyBJXIRrQwhp4D7GN3jDScB30RBOO6WyZFa162HG8ee
GKEGnZYNDi1ZExh97iLAZgQWI+YPDwEyTRW2CVH+Wj5FNkbn/JtgWL1wH/i8/OQK
Xh1g3f6HxU6aac47mHOdq/IqF3oKTBergRzEnQ7kIJ1mHivHAD6BeTbbt2iqBd02
FtktznbRgttHu5bySioFfpjXZfe0KR0wMivNXIH9q3g5V8tRC98P9x0gGgCBRlg7
JWzAneDv7RcQQyvIeHSCeeaamu6GdatUbedDlSUUN/3zb6g+a9Hd7fhhzdBkBOtr
Up2fxn4gIR7J55xeOipFF/p0a66F7MaFk9eFeJcT0UCIqgw7IOvo2rrMNwkZNUY8
B1Y8PMln2SNufpwNgj7PkJdDBI8ejZlRp195FGYiZZUC6g49fFna7FkKSnxvKqP4
VC4iO4HKElU8v664i5pmEZNAMdM5aW5/31lTsyqIB2bTxqvmtVz1hmsZqP73QQWg
GUEzprzZ83YlPFeoIyJ30UhVRJCjkx1FJ2LmozwZ0aTDEkTba58UZ1wACG+e7lmF
eKPhhhjIK4CmEyBWHWHyFtBm5SGPaIjP6qgjGVKmG31p5EjS7yGVJTBNLk+El3Q8
v7t1nr1S0yERzePq0d5uPuApOx5NvYl1zLhLSSUNyPmrVWz3yCyfzP+82dZuLBCo
JrufQcDZpu9W/xxa0tFjz47VhE9vecqNgnauyxLJ/gMMgn5llKcJ3lLaXhOgco0m
cFplAtoR6SXIyB/3OmmvdnkUMp0N0Gn83GgSwKEyzxU3F/j+fUfUwhS4V8ct2QEO
zV35w0v6Ks4jZBMcpE60oyptCr0Kj6HXS6a9z86pYU6vSayPxlTXJ1fRXhCAzMrj
VhbIPdcEuXz7hFzmYsI9fu+k4ntbJiLHzi7WyEVytRgVEpmCS95QKDJFkG92KYbE
5ceI8utJBXTquHmuOkdyqLfAu5MQqoLgXMCEtXwQ18AXChG2EzcaPfLOF26UyQDP
lk+6OZvoCOT0vBXQIF6hVwXkylda5mPkfO48l8t9UKqqpyhSDcY946ZvkFdrfyCT
7FLfoorGm6WXefmHG98fPSfyYwRk2p8aQ+17yeXJif2P4TN3/i0YyOSjka025c36
P8A7srxpnIUk6NwMxoiGT0WQ3RDppaSzPQjQoV0S23bJPoZYXHotdkkQuad18soX
OFVCxXzEfcRiPdISRt3zGCDfDfrJrWejRPN5f0J17xdj2enIkOYPjgSoZIsFuob0
JU5mA8bjtzWl8nKv3nuyklYQ0S+Xo7rLf6rH4fHKQMDLkdizpZBpE6eYvGhBoAmT
fuI2QWItA2NBjv2tXTVroiHOpDvh9PLYOS/c6cYddFYs87ljcAXWIFJd4ycgYYe+
bfhY0i+e/jmDHVu3U6KdXzD8ZtEUQ7URgc2PR8d1pJJ4EjDEjZOxv8b0vDdpKQ0L
PA1ejcVhOOY6oDAtpXcqH9hmsph1HZOFsn2pILe1Kx/l6cxQDyaG9C3447NUv+DT
xHVMMbp0pafAmYKKsFaC2agO0m/ZWv4h4bBSdlmFvhIku8RFis/wwXs1UxiN4kuX
v0qrHif4cMqwuRR08xULHX1Q2HEzEMl1B+3sjzhxhhoeaHuvN8hiqaz7OMxrifj3
DKXwhhaRoPHpi6oBmKpMWomnj6GnoPNeUueMd4xplZWcqjerUJAYC59rHXTQ7Rs0
pqDZ7H9LI22RhqrZIvCGTBgiJZaP0Ff7Xn0UjaSegzE3G96RKhoqo4tlqL31LSzY
tRtpuIyUgprduHIl8wRthfHGifcp95EihWf2+nQ4X/Ng73X4f6ZgpeGxLkFGGUxR
9qOsN2DKN+MNcvk4ypnfU0TcY+HGOc0hKyT05fJEOZcR2nFjp5LmQi5YizBm4wWK
4+u7Aj6L0JXBrG36gbyUmwZIqmdlWOWDhneZfyq8Ftx0ZF1UcE1f29R+GTRVg9VE
4aYIBaOFbzVDcr1zvMJqbNeIKoCYEBRkhlZOqTeI+sRxfjsZMYyvCiCESQPazG7D
G6CLwuGtE7g/YtNwIb2JxenD4xyb4GPly8QfIUggpqdDRs8dBf9u4Zrt6JpGcICK
ETL8kboOnqkBuUu+Y3wTTqj/jRhXcRmVNrZWEBWcvAwnI7PdEMca0bYVUg4zhiHd
p4T4cnpEDPnnJsh9NGz9b1DDcBEuNYPxL1ZVcolYJreYugsHdU2gORfZONfn5/Kk
5Q+o/NKTNmZ32XrCl4tLnSz8oKwSKuxOiEe/7ROpEeqfd+tyNPBv2wlViG4+XtYK
HWxcyARMbKGrC4oMInkLBsSvrq9geOMoqwwPrk2IFhbjvnoJW92lKsWBxei9QSEc
k8+5qSenNKshg12vFOeNMG2vgmBzKg3Fkaggpb/+zIWSLfWq9LQ+r7tNnnj2Jela
9UuRN7umGSvfFszZKe1HgO8q2mPK5V+MAfTLRSe9Egael1hbdxr/ldyaKU9dqp+j
56d+dR7EeA0ysp2FrQKixeHq2e8qCx7nmin9k2/IzKzqEXhYWmokJU6ehKxm+Dxb
`pragma protect end_protected
