// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QHa4PQiD3S4cLXs2CYp3KSVcIAnAV8ilUPSjdGd9jDhD7YxNP2cZoMaIUk6ibcJt
uNXI/f15RqV5PQaP9OSlGjhe6VaX/OcXBGnzEHnN03lqA9N8p/VoSoI87Kqae+c5
s1B8o4i0E4KguxUIfiWfaqvAAy4wkdj2D4GaURwTKYA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10320)
bhdZfTbMHx8jd+VyQNkYpsRak1IDTxRk06VR2dG8LLym49Cif62ezNVS/9R8tAbJ
JSTOd4pZrGAqbvRedSaM7JImEiz/eDnzajXAyZTJe6OXcfrutGngNfJ1ABlIq41i
z/yMe6Z/7ONUf/cW5Bkx/k69eSNt6fR7S5PpW7PdzwsABfJv3qNuQhAkZXkLZgW0
SUHaXaitd7pgiw4/KM5SEWVe5kWT4/lQb4VnjqQIkubR1pP1h3H2QZ9fkGK7axYp
Jcwm0GqzvCp3zF2Y3aNl+CJz8rSJKMlpnB5CU7UAfRWfxMRFkIuQLOkb0Eh4fnMg
BKHMxXAREsIRRy7PBuukM/xMkDjcFESiXqEEDqqKijfczEE3gLyCr0cTQvhO78eX
8wQwPXtsY4zbkfKSS/vMoAdBs/GuaPMBX+yA2D72QuUwoilhtCM2Vj7mnDKEy8EG
vTPwrEM6rxEAteVqqsmhwL2e8KsnVLRzKZSIziZkXoCABbeIaKh+tRMOKa5Bj43b
eQDQsJxThe2GbKN5jDg2QuT+En4mjdgTmDhlRG9p5ZltUVBMblJGOCsuChIW4qJb
qTfteyNjkxXh3unWE/n3nfoRCdO8JsdN2aCPDV7kc6PiuroFpUzbvZuQvPzLkX8o
pAmThkNAfUZ+vDt9+LhjPMMxa5EkbXD25xgn56Lk2Bux/nSUD//4lFBwwnZ8bXxW
T/HgOrUtDY0j6kUKD+en9noF8Kw+LAGMEaDD4l4SDK5jKwa3rwJPzEBYrpaio6Xh
/q2uaa35C5rULI4cfiOo4ezK/dGLrfyBdhcPsRCe6jkQEl/uoW5x2P3c6/kDB90j
gAYA7vgUah1YbADOdFnnKxFlbqM2H/EM5z1yDiy+6nPwaugBSkU9yBzt5PoZBpqx
hV1KxqUnM8Hnn1XFpuPqjMo6YXCdGGVVLzPGh/+gZQDC7XI+AlKqSLQvfPNXIFLA
p0Ng83NGjC2IIM4h/zgldIRvPMiwzcBTO99f2yaFNtkXDwij3cS5ohlcyU63BGLR
yuiYqqj4hW+kqQOilgQ9m2Qkp1uaBzK5/HYObQLAk1ULmFJV8iO0T9gVYsC37MF2
wDZyUkX+qZcGmyHdYCKAPQM87P+o4U9vgnkxfxCPZKeGbbHdzR0efLAB67CenCUd
35g6xB4OFD1KdOHeSWQfF1e71ffLc+g0L3XKiRyRG8s9fo15lclH94jpellkin7r
jzDioIiEexzG2TTBH9LlCjEUL/jZodbY0h+UcrbSdIJvI5xL4qR0MKA4/ZeO1etr
WE/a+HR+Ii6ZMQPBKvwfV1WbMrHSK8MeuSqqCcmUtPalh8Unx47FZ3YlIdqlj2yh
3mXwzQgxZcW1PGDGnxZdPMsZL3wpEO8b8itpi1+0vxBjCvYE1MM6Ju2C1keOw0Tp
JmPEz02A7vf5eTiFTHmJwvADvut1k2cssfrQJukTjWthIJmHdY0skdM0a1JwEMzP
r/3uX4hMoXYmDajGW8vNyG6nq8sKgm44oCAu7CM9Yt61LkZIQs0KbYa9PelqkDYV
74WjpbmSM9mdKV/1XcKscJuaDRyRsxTGZ+U4Yp9Ykiz1ibm5Nsj8LOZmPESInbz3
OsNqY6QWsp5DG70vEJfUraFoHQ+69KCguioERqK5isotJ3XJ5kUx6tBK3fvNBLcD
msM05g/jNTcjJEpHXcZjmlS3naThZbvgPtK9DiSTLa8NiigE3OH+jtxPzAdOYDzU
tl8zHTJP/TC3zVFstzPkfNd1XcQ4i9R/yjuwnU9nlAnvpGNtz9T+0GuhwqEtYF9B
77oRSu3ybO5RsT/4CP8mZxy7n+HE4lGDUG6AgRcfc07L9XU+v5yvnD9+45FEl05s
gkfRN96DvJZKg+bkhB/N3PaNfkqCWgiPra6OqwYXdrW/NJ66FLbUL9uAWJk0EQNO
0UJJT0BArdgYQlmxA4q84I+Hwdn8C5w0zhY59RsElIrzA+nAIuRv8HQ+u09RUdAT
wV5lv4ZEE4LklP80x1UFYD8dXqyO6NWwzoTfN3C6ADedSjUn3085QciJ7yD7jWZQ
ziv7jT6EXjZm27H3B81QBClwo5qNLTjSSnXNQhOdixvXM0rO1ssgymDt7V/3pUZ6
MOa9EaanWg33pTmd11wb39koZ25998jE9koMr+KvMYRh+Gnv8hLLbLLzWwJcw2hq
SvaLxs0nRtRhT2Qez6/WF7uzl8k1N3dNNgIONUoO2JhP5YFcZFzwzluTnvWwoS9p
qO1lQwPQ9IuTg5LV80/Fdi6DcQdn4zGLhCJG/kIxhpqOPnLBnbrINXo86KeKyBYZ
fyoR37AsW3LjJ1Qk2+U/Xs4NQGHwgpFpAVHP5XRTbuuLthRLnrMSOYElFeK+LeOx
PEw8gWV4svC4YJERN0bbYGijujzKtH5FSSMdXD0Vv0SvKVUvMdABk8DT5SJL9BAc
d8z/DeKihcGZWNKck+IImHP12HyDbmWAbddpB6PfdkgvlKGWQH46i1eyOScKE+Hw
3mQqfpVqTp10Wz1cZ2+DrKp033SX3HLcneH5wtkxVyxKNg68tA1Kbppj1U+BLFyE
OOsi2jt9vwu8jS420iPrQOLsJ4+Y62ul0YBgcBAu/PXvpmvlml+DGFwcwaQBrp7u
EJUZnuLey/7kIyZgpAn38F77pOHVoNZL8Nq1Bn7zZQCe4YL7PZv6W7/fYcnOxfWa
A/lP9/xnFmiQSz9hGnJ/HE/5lSAVtmzGBrcSvgnPfUP/acONaEfQ2BpnqKonEBR+
Vq3KdS+9pPUZ7/8sUPLzC4X087a+8xtZxKmcyXKx23g+RdsWrJOWpBw37qRgFx1/
oAdmJYR/hl9nmRk2hsIQxAKDK7afT98vm1//a3W0J1HQ6gvRLjfscIAttQ+TaAm3
HwVGI6kyM9k/2QIO+lKq9S6zaTZzEbKp0wj/gTnwpx1Fs/FnkGrj5GpWyr8+xu1V
mj+Ri0Yz2IWtKo+0b6ohp674AOxY5RT7O2FaD8m7qp1oQs30oKZ6aOOGIJ8V1Tjq
TE8oEVv/wC3dM0xA2G3p3hPKmw/eqnrIy6mXDboguo9Wi9mTrqy2Kz9L1JV9g358
0v8UmkGYF5c8WPRqzSJYu8mGgWZJ405GjnfOsJIOd9tYfj76hFRdPL4FUfrechNq
CmiXfk29eAoaZwyrby2Milg0RK/Hr8noBnvG7zmCFsCe16ZA4AWi2by5NTp1cy8H
ElnWRWvHBHH5Vy31KBvROtJsFFQZOC2siKwm+cre+11yd5VdV2Ih2Qo015CQCdDc
3IUrV6Rb+Bzg0P7BMiRL57NXo4FJQVhaPUiXfGsh/eKbUfPk3xAlEPVGDduu5hZ6
Srjy7dKSDHKaUglpuL9Rxap6JIS267VrA5+WplHTNJt7l1Zn17jLhX3crRSnNL7H
SooQHyptFfkfXXUo/hvW8E+zCvPshmMjZ/AXXXuAAec+WQ/H+N5/20cuBqFyChy9
fDvvGj1KM6bUsao1h47HCXTsX6/ce7TKJMk3L/UkLz0AOVJSyhNdmBG5B3zHkmY1
9Y20001AP+V06Wm/gQsybtgFDKDV4hJFgSY+U/BknfFQvsRBXzjtyZB0krEVHEqe
nCLikHYBLQsjNdD3THxy2ZM6KSY2EB5pHRpsYr6q/1W/6hZYsVMpDJgu1ttbrSE7
mM7Yr71mL2ZaG9o/HLCAylF0bUuuXjeq2bGZf27lV14diZZ3BjVl387j6VYOEBeB
I4J5CI+oE/wCINZ0Tx6K/Rb8wTEATVVK9uIQbV76x7i9CKVK+eITGB3ZtbApM65k
8Fwm2Q9xZ8cemM7sbuob9uHob+MXIjMb4SlN0f9TRn//NFsV1YubTZvDeqHqdk1r
JNSHGMID+NnW1RJ0Qg78NjkkjzCQtlc8gLSa8NYd/j1iJ7X3FWIhwb25PNojgIFQ
Pm5jepN3XJ7DgqhCyA/azs29hX7Fbjb3MB9hF0+TVMG5v7DauevRPKzpNNNhSDjZ
ed+zCSH/r9NScRWhuhJ1VVK1jl+3ocYIAkMsA9pR4DYok2vUrrTmBC+JDjhcstW1
qoVnaaLhxBv/TxjE/L8dRLf1Zkw0beIAiMnypkIzA0WwXUKEBQH/v44aSlA4qATq
FiZ8jKF08G+4YmePqCT2ucOkfUz3qvw05VEy0gXhrkk+WKjA1ESp/4ZPVjUypjBV
q41bQ80wXVQpyoYaT6XysycNGbfmMbUTR8Zaz6v9kdsdqz7qviJVkNzNXJCvqCr7
CYIBV34aKDm4lomeciu9c4aeASor24zq7klBrj6uymDV35cvVwinXajMRziLreG/
a8QyAFO38wJ77POX8Ggp7964zviKPHpVOToJiaTPfbqah5zZwPXsrqztEB7w+W65
+P7UsIUA5GwsAVQa6ZCH7v6QKh3eOlq3Gmk9XM+51H7MdniSPRquEwR1IgigAtLH
Mkitfh0xwWRC9X1dqSS/LtnECwj5iprIuVGbjjZAFVwOZ9Ljz7cncYoZwKW+YN3O
QhHTMAp/UaV2Y0r96xYIRHODmJotlLb5k2LbWLXlRTQqwMtZQxrCIws9DQniLGP6
0MELheWFEQAtwTM+1O564O065IYldR/4q/FKkDa3XQ2KLgLa54TsIVSaVZsyurfS
fBpDsj6eu8AWraOZPbkl3oDZoKK7WL6pLj0EuoHK/84EAmvwmSJhk0jAqO44mkgh
dzWHpwIHvRUHEi81qojvAi/7fc9yKs6yoyicYB5UmOXsIV3uwVeFOqGWoSNvEmzA
HOuic05HC3u6LXFYiOHH3bkfnQOyHba3VKa7ZazMfM6sBvRgNTw5N3fvKHk6gfCT
7mIQ5LPfpP5hz/hgzI/CNpJNZ2EHcVzts6qDM+tUBt7J+X6ybin6TQ8uhkM1/20a
uKL5fu11lKh/s0++VA8Mdk9Qhzd0J+xC9Wl4qo+H5WLWZ8qdfNZhDFeXSiRJE72/
vaHe/of9Vmx+v2hbxHRAMDViqb/pU0WNJYeV8TNlYbaiAMVQrSobPxSZGeWL+Qsy
0qyqniOiwrh6X7+YG+dIrrz/OZztiBIv+Ihv/F7N7ltyR7P/wS59yi3QDrq/tBi/
CGU70GXuOpH7Lqo/Ac5PQrPN491RoNafO5nAXn3C6gck0ekf7WlXK0OshiC7v5gM
2Nm8QdwrdQg2jvoH5RSkV/eWlyGYuYqoDkzjHd+6R1WSsIe4Ui5u5ubI0g9f5rYU
Arg4ULOcI/aTqLkU/sGE0DWRl1EUmr9noIq/0fzT/qyfmScUWOMaSeTq8n7Tapm2
2oYm16Ksk+he29xDzd9j/yltGq3DJOIBVyG3lP2ddICEOZwiKKepnyGod3xEJrdy
1B5EeNKhh0qQpE9x8BvnB4tH0T01h3y7FyfisGJKK5uWx+7XQBv5U3A5FjX24kld
11rLDwy5EVWSCtiuLDXGie01MaB88cQt9QDZThHziHiB6huXrtwGKSb3zkhoX+im
H2p+MJ8IVXtWhocLM6APnh+mTTid88u0CGeSWUJJKVdxsmuhd5HKhRI4ciReIOPF
41c6vBq7R0+wgWK4iEGNqzMRk8jQQHWyuICNGqrKNz8zVJALHO7QYLk9xOlZXz5A
pX0L1ByFP1qn5QOV1sCnDt2bwVnW2jRO0qeySqQE81CVB2IhAySDRncZtTXWLFwU
hyHpUT0S6tf6YxRFqEkbY0Zh27wEG2he8rguFN3qE1bCIgzvr8sUymGzVLMP5CU6
VvQCW2BMeBuaVAz1sqdY+pM6iWhNbu+lPQA8U3AbE+sN0x1RL/86XHnVjVdwsVm9
REHWFruf2Q4AhnXKkU3zNrQUaA0GsCYAd0jC+ogc2bpxOY1bs3y9k8Rlm1jtaOu4
ZFMIf1sKydQKfeNANwjziDvBzi3j1Ay96+B0mCuNDWSN+0RjUs8VnTa8AG/xL6wJ
GRC/mAKXH5GEkhqd4npiCeyj1BjU0I1XeULCTjPQTXa15Zhd+42/a5fg2dq9fTwC
K9vZo79pXZoSb9FTnzv/1W6XFzvp37cDFiqBtRwSnBEB67adIoKokpUUdwd2dTYD
QHk+Nxes2qOh1gnD1b/+94FHEHLX5ILHSayzpf3hYsZuhySX9OwIZ4aNk4mh4oc9
Z979hHZLhjG9u9I+G8EzHzR39J2/v+/TwekY+su0sq6xg3yCuvXntxvStWzsXwO5
jUBOHrm6NYTqXNkSmXcf6MzYsV5rGcV6yJNyhYsLtWwOspDIqfYd8hytCZn3b6Sg
CgfZNT7hcwkYQKPMBdTUZhQdk075NWGW6LdaAYCaD0ZBuR2aTqqVSBAbyPwYz10N
VS1yce9plfk0tz8VGZwDEqc/O4PiZqwg50aJiOFSKes52mLubvndOy0v/U6Mr9Mc
Jv2EGL4MEP2ZGcVo+uVU1SPCO/CyKaxBREVY954jlbII7mI0qNp/mXYCafb6Dq7m
ISiUTyEYXFam8gJbbcodE6zRb8nfJbtQ8yhjEo5DlPTtBPLvXuVKwWpWU3J2yTIt
DAo1m/gdybcYdr/b3Y0LwVME9gvKcZddKj1qyDjeIURO/SPnWiEdEf9YfjOaEXHO
jUoY0I5ttp/2kpatsxODS7C4K3NT0b0k0WuS62cOuORgk+pw73i7e7UGx40Bo6Fe
dgjddSGLvB9JBFbEtTBL9EvCiSSjFO4pMZFDQEe1XZuF/nKdvV2BIeDC6qres8ta
lzYm1N+cBTPVMBx/R85H3FUwLOrJpWyPL8K5OyhzyfhbNYzP8eys+GMgvV2amdpb
D7yWNOdP6Dd708Oh/oHiLnlPEYG2V+e2WTySvSB4+COxWujufcPWW49vhaP66KdW
72rYu5g69KnyWsfYoX4Kaoio3+9CJO/LrmL2bHxdg9BAhoMAiLQY0tU7UYBDiuJ7
/ElqTP8/wnCHOYxxCn+sTnMCIjPJMNNl0kabezguhGz5dfjN+1qUx4asHL/y2/8K
gA2hJQN5GYDiGu/daEziRyocEmW8tCMukUW4ZtKwsrC4IECad35tWQ7cqQ5aU0tj
M85ehVVHqyDOTdhCO2rhj8JvfCP82aasZyHs3b6fAgEb2lfwnNo+86ERr7o7clr7
bLERPmWOLWu29yr7gTLwXgm3K98WEFN+G+z23uu0pgEMmbb6sqBmlOsr4CMGDlXO
zqetyWVGVS7RfpW6SO6c7rCHPwk3Rl0VkZqw40JeAYQrTdQ0c9MSDsTSVpz8XcQa
P8rffk4fDqHnTvi3zwNPeWKGeFleUtjwA5PImUnc25a3Rt/Vb+eL2Li1k66gousA
6umOVLdmYEEcjQ8b0jP6Xs0JnOFFypYzg3cvAq3Src8TYRIxqlfRix8NiHvy9mig
WupwRr8owOJjXhslox6vANyDV7XOSXP6W5940vdZUnG81OKH7NCeHqRFmup4I/oQ
oMdqh2u+eacY6tNljHDvRu2tmivP8rZvhf6IL8vo84rrGeeSv/h+C9CWSWtq4gYT
Pqqf33ZYYNmdBBnB9w5RqiFJEvkqLrfWSQnamzO563eJmXbvVh9xXA2o+5do4Cnr
Mqy9wCBaUCAIPzvXpaNtZolf/0CZauQBCs8PiKy5QxmgqvCkWTW7fCRhtAXaNVpd
GYFqlGl0DGvFXNkxf+C25MjnlW7Y9VzAt4Y9AsFtAwcbg9yJYYLjtzQBBYwT0EO6
ASHaYZEZ/rk1x+QacitLI0wNyUKk2cafhkp3sBaHFrrz08aM41+UF13QIAYFUfwk
EwiTeHR53VM6+DnDAoGxMM35bmk/WZCpnFqpM6SaX8Os+8XJGviyvJS0gQQAZGe3
ETaZVBOUJNlJ6offJML8CQevPeCHrhDIMruoWD4c0EpiN6/ZijbXTPWBDgkx7vcZ
4JRj+hthz5+HRsM66sL7lyc+lVBNh9TaEwJAByajJDAzbb7YUp8EnepJGuGnAzyO
oDOgWz+TsRkyjGSX/c3iBcyWyCv/POYuQ70lzoDywPGL7+GSFAoS4lFVmSYG2Z3o
ZIJnsrsqbOwUyf+AdMwn4eofNX1jxdD8YP4biLYdkZ9YPT9BMAlS/HNE1Usp7XPO
F9SYiV9NHa/j7rPYAeRabyw3xZ1dihwRNbx0MOpwV70lwuaxHs7VkAOWgeJi6l3P
tk5iu9oVqSFzHbkD5cvZLq/Kfef7v/x2M/kRxh3E5fwnN6HVOc6v6WnXaNqKyZGK
MlO5hY0I7xDiSsd6lr0v0VQCmcYg3tXMqrNIFmGgeHgFXGd7IGVDVbRvWe0izvo7
oW45rTG3wLUToi+AkHS4r/lbQ7TWydq0V+8DofMINY1I/3AgxvHvMXfJ3q4sITQm
YAeiBw2A4MoEeKf9r2TWjTdLbm0VbLh2FBtGKICHRaC+5Yl+QzOGyS3vAGZ8LQ//
u5PNVb8UhS5MOBYrnhWQqvDlHbm8YYfytKtNbY+BSWvKyKeijuhAhzqwZSRAqaRU
xUU2pnB3eWchNL82jHmsAsg31E8KH4S/tFYydX0fR/7aIpWdIa5vDZwQIVI8xqLU
HqR1yUhUuGxUFDklk1uJgCdp0GehxLz4bsSqXIyb926euKjX/WpH938xrssY2yG3
Md4agK723Qh5ll3ZxHQGOWaAof+vFmzSEo+Uw2cERhX4fslWx7cdOy/xjZhdKTJl
6CN8gl1VXLD8ihgjjC1vN7eottqpx3KS9V3l10cZAwPqV7vvvxzcuUmRfXYweTYX
nbMk7gcaLCEY3EhfyZcVyfRfC881dq39CnaPT5ihuWzLdswARn79ybr7zW0nh4NV
+u2Iy+sRlI8sbkZpZE5OMa0qwuKfk9PnOUwRTtZyiBzZWYn2g3YtSk1pzbnWNu7T
bSGJm0u2WvI6mDvrN92Zl9jMsq1qQT8lG0k32opL6s9pKdoWwUhcJfhMBfHqf0lC
5cpFrztitBd756yHSpoWRXRWAOjSmApxLMLsocsIAIDHO2sI///jRsJWAOKFVp5p
uHMYr+gvWatI/Dl46rjnVToP4x1sFH9PUAU7Xa/9X39DFpMta0n2UDGINWVD0dG/
1PSlS2VDkE/ujAucg0hZJMSR8FJZw/QExlEl+X6y7m/wW+HpQVIoJ20NIzYL9Iwj
ea/3d6vjeJRyKGTTp830Csbc8z+wxKbAoxq0LWMKKvaWnvaV0cpb+CuAh7AMvJjT
Ks/kH9m8Whtf4Y+2QY3/VzI+1HgHk/wiHlIOjkchDwpgVarkrmcKjm3dQW2QCOYz
yEzJ58Ouprhs+itcdNw01XlnSvRgyLw6mLbJBIwaPuHIOZkYDu7DkMa2xA6rxYnr
eyuqaEEsrIoK60TGBxAjpzAVK5vcVJ3IsyaCTkYUMb7fjp6BHFck6QpSakmuRy8V
gJTyPtfOSysX/yW6IFA1hbvD+urYp1Xbyq2Eiy8RIvFsSdkigtYsX2NgUIL/PLpY
x2edhaH+0fUZ9RqaSbrFd9Mt/0/SISYmbh3c0HHGwlcNin39YwDCmEGYqShsZggx
qKrU8VPgMa/FNQj3e3ELgTk/mJN1js9EyeG0f4gCSPHCxSCWePgkJqCLNhqJpztr
artxt7vubNcUpXTTvZnuWvC6/oy4UwJsfiEGgDS46VklurJXNaG/JpiXHMHzQwDf
6BuqAueMoYWNICR9AwYHYYhzzySJ6lQYWg+MeEawJpfCUWVBi2RH2Z+rIHTaCZlq
tn0Mr1T9w6kgclhyH8V999rEHmoWlaGN6trQzynUdJCw4N6K6/YrQ3JNWJzQkFCK
3WH2DT+dS8NNpO3Tcp7UACXVOkAes86z1gESLWXg9A5t8WL+maxsdrDIzWPZDTLr
yyJubwPEjd3InLku0Pv7AqJLK9EkVd1tVYeuuTuEVL/5F1vbOj9SGtm1qhLbZx91
tBA+vFzkjaMrJejbrZK7cvItIjaSTAgCwQyEICAirSa49qC4jFTSB4gxZvfAOB6J
YX7lM8FEJKfvOVXbxutqzYLrC1s1NpA0Uxd7zRADcpAge47Wi0NLmEyeO74l8WmM
XkG12ey0MHxNvM5sgDHKXAg384jDiT9cKP1c/4tCna4gCgEjYbv4Zs8LKZFla4UV
SggI2bCiksCBupCb2knjeAgenwACHV1xqu1gp8WrYNfswYSLKNs+rBiI2cSwC9jF
xCY65Q4xN6PP6MZijSxAcY8ffzBLja6an5lUX7O76pmc4u6G1OEYgqE/jnfY9sQe
8IeODSHxn1TPLt9lKRoV/cubEiK5kl5ztXyhX3M09LusUN+oPu2gMtGbtq9/9Ux6
sZpnGmABaYzwZY4ADo8wzR2m8boKcIV3OYq21SBxK/ex9LJq3GWOe4nSExbN0tPy
hGe7y9kWulL8tZ9WU/SQs8qZCK96S/7Zjkpuv+xjetGx0+WIPfnV1lJ4ULte1N1n
3cZ8Ikrgs5cuxA3b3JmBAYPsgi2/nDad5jQ/Ez0DLE+ydzPTJ3A43ApcO9ECoXeI
eKwuiG13doh+nm9nmD9AQzzgcvW3eoRZGGSqus3GywQKorL17tbey2tNZftqA2CC
g87WMVe3jQlXzokLxyCvjG0yWeYyZInw6I+j4Bu/Am2GqNATR2gdhVhJ5o30x2TP
3hdLfP6uMatpUvyufW35ieg0NLSKGi/UJKCef6/guzPdy94wgi92/Ciuj1Yx9ZLK
XdsmBUpz42Ewz1VrZS5Pg63dxw00rnHagt2JsXJ/WnlGA/cwi8UGrFt89CXexT6L
vl7+JvxkqbjL3EAO3fcypDpbvYVcpsrW+WH7p/1POz8lw3JDS/euhyxFfnNaZHLI
p9i83fukCw35SCAG/r2VNvX400M9FNQ22GKYuZXExwvXJaTRQi1yv3y/9rfU5Igv
8W4z4xzfweT/xPt8ppgTrUyGZr5oJmgKWgydd8scsnCiLk5AtJTc5YyuQVDf2qsY
MckUqADwAUG7zM2ly0g+CIt8Nyx6dUV93F8lk2cVF1eTYCL9zghQU5WtGz55d1fn
wSGtcvzkz+MOwaSIKYkFJRY6Kks9YyBUt/bTNAdTJu6BEZj1TeYZsNtnd7zZXp0q
dfrXlSmn5HtoOa/clHzw71QWzcC3LcCr1LQrHMMWBIiAtV6MkyAbk1aRS6QWlUdU
DQJKE5/1dN6Q9EU39wX1jYF0u81JCOgsrD+lrkewvSuKlhd/3pxqxlorFX9KN/z/
xwYjVyZTzkRytN/iXSGajuG1EYPqrKrI9aSRBOsv8r7yQLpXpRrw5os9D9jb/7K6
P5ZHVzylG9pvji5LWf24AIjnf5PMKsGDcO3sbqmWhx5941egkVIrfIMTUaBSm3qG
LOhgrj9oxY+Ae8f+FPimT0BXi65GGOysQnUN97GenVlhM+d9+veSC1g+aNc4BZJW
UCcEzC2GWKOU691m671P7c7zgiX2uhlEeqBVrTO4FsEwqPZyS1dieAtYZczlnIcB
n3tzZ+kcD2v/umnKeSvrFVklBqEmL53r3UzOkuIb2FgUNeogBitFR01ohUeytRva
PqhkveN3kJBqy+D0xmUzT5DbWu2QHZ8PmZaVu9zagqvzFvn9ImnAkpgyEntuiSFe
DvTpfYiZ0cusJmjSSjaAfEdprI3leZomtdMr9KkUGyRSvni6FTgeAJdzXs4Ep0tw
aritt1LGdhVCgTqbJ+p2lNaB7UkFzLlOY+bddZUxoINl28WnWA/+0wf3DiDXnvnJ
M/XLf5pbFVJatq/zqICckf0LWa0yqc9EE6TPoXyOs/NKFw4MPwc0NRXCMRumXpN/
BaJ27SvAkH7fnHR79kQ0Vg08+2x3/yzcXQFsDvpMv+yF1ixrPtT6AkeLbMRKj1O/
WxdBDuTt4AUpP0um1KZncU0HPPtbidgYcY96wXmis9ZLcU3xl75tLHfLBBHbD4ZR
EXQZuge+tucViphHeqYP64euhFg4xpr+EEN2nAvLCODkDBlfgZrIzZKRSQ8mQD3C
3T/mUgcsufObFxVvIRs4kM44HYm4c+z03ZA1geqFw6gos6bbKzX/4pWp+oXjqIwX
6ffsAa8BjWKuVuvZaHsr4NxKkCOSozA/bzJIFVp4ncJqGo8w3UbU9s4SpbbD0kmJ
POFG7gRVKX9SeBhKV0Vc7EdUkukUGycWBHiawkRS1usGjjU7i96NjQ/0Jq2ECLzo
TIB1zSG6CVz712wt10vKGpg0imKR4wZjG1QGpux7f+XqhbB+KEFYRdy09y2UUoW0
t4byqNFZ2EfAsNkrZ3Bn9+3XQdyTlBhw/BOmT8Cre5j1pUnxGFTOKTIQeSBCs2y/
j42veqPAvLAFOz+/uPZKIdiyi98IoWMUYv9vMGTYNATzwcNWMdkTTOuAYFNsceLX
1NMprS5G9mqY2kbg+kyaBOI9hjfJGUIYocps+JpAFNqj6YzV2yuVlPKGp0rgBtEb
vqv4A9fXq1WR0y3FrbFUYbm8f8hRKXXWwziEHRnsZ4TWgilQRGv6JTpv30HXSl/v
vm04baV3p16zY6i+lknhQlo5PPCyqBIc4iZDWMK+nd27Rvd12tDIDT/yATNjTcOe
+oou/dHqE91pP6HpTdw6kMg4hicQm+u8g3eETyXycQb62n6gu6vckZx30tRPsE0G
nSbsQ25+JlSF1OiUnhx3gjnzyZBlhkp6c4zCiWoz8WMUg3qV5emqUIuKdHCFZzMx
x5YQ8zvvx3d38iOEafiW7DkQ0QWyb2vdtza49uk3VnAY7/NK1e6d5R7K9IYNobgI
3clzEcYSEbjE4b/8fAnXaHFuK6Bcppmbe33HtjrokVHqw4Yii2PvP2vFbvsdLSXi
oCcFbAWAENkTPdJ1TtzaxOpYAKM6l2DDoEGw+R82ChZcwjI+clH43bOYqCtDaVLN
WqJZrxA94hbljqdu9TbZnWEpWKgeASJVDAdiTz2l+1TEvS66qH6imddmG+pSKUri
7WNVQy5IiPgtOsx46RwIvFD/7pMQGAcGj5bYt5L6EXLotHTHMxgcX9wx+AsgqE5j
IC87MYCu5HJkW9lwBB3R1qUNI9nfry/eBStAIn2ltdGEcFoBjqH1thhDm6nD8HR5
nckk9VbsGVJ5YrOcNEkSRXEq1kHQxdgrSkHhJ18Aaq3BSf1D/BKudP3YWgV07iFr
AwyXhE0mSjbjbuS88ro1NQUMaWrQE1v2BUFENom5gOrB2ibmCGW9OFWZTGFE6zKB
TBgbt/tCaZb4PsV+AkyWg8Vicm1oRUYnZ+YgPyEv8n99UZ29rYZA9G84hc78hCAb
dh2p0eoT5tSlqW7Vns4n9CXJK7goQX/gBc8+6HvyeCAyeDiBtO5QTnVApyVHELfY
42TTQDMHfqsoEW8uPKeRDvbpvhLAyfRNo6XgoBlv9AqsyI+xhanXBOsGcXeHHiug
eO33WKtGAsyUG3hI1+fyqaIXpko1IiPR2Pxu7iebiugVwC/NvDAOcJRw0g045Ib5
0wT/+FjNOco/eDujOBW2Jl7nxAPKDlcpT8U5SaNCFzzLnlQm/qEzCwwbP5scj4q8
hBGFpBhI3TOgGUbIxZd38AmatQlJSL9mLECqcJP0mZOClc3lXMPr9Om+O/Zu1O5h
m6xNXAYEPhmrdgDq/4Rx63IM8jNQmqTOJUAKJLSuXOvnFxK33+Wuop4ESkIk459e
S5QO6Ow7I9/6xxtAVKpmLfoEdOpybPK+et2Nhzw8lSHvkS8YkYimq36TaZsmo1nj
KPMjUyYjl0HqISSmw6F4sfhuqvmrQp+FzYCVF5xYy/nyZ/fWxIOutO65d3ECswSb
UjBULSJaLzDJ964uQMngFRBDXpGcKpEo6RIn27GHT6f06ixuNWexMCn+iehoNqEL
vbD92f2E+bHKmtZgrv2lZJgSTK6Og2cf9jNqIOKcpo0NP2wpoNUR019ZhyUx97o8
`pragma protect end_protected
