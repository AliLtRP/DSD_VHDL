// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
iJgN2OyQvltW5eC/e6uIX2VtbPMxGLLnJyugS6tfRUqKbZA1UBDUIpMacHACOGyhMF3/OGNsWZmb
gIvLrAYvm6l4ZyGD91RpN7O9+B+U7ffvdvmxGg0rs7CPTDsh0VrQGh8ChsNFQ9iF2t8dlNVzyWsT
ZJeqM3n8pkbq/48h5L7AQaOSws1fhm7FxsIaQHBpHInIaTCQpBJUOrFiFFuOSdwM35zbQyb3Uy5b
uT6dz5wSgybKaFQZjE9UyUmiFAsFjBWD3IHvXH70ETUwDLEVo3sp/NZ//wRdHoOHzmtmq8HHfHx+
+q0ZC4ctuaEJj8nvar6//UlZ3EtTtAjbL3MNbA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
dV9sd+XtjuA7a/C8nMC4kmdx14J8KLX+ineLCPWA8N48kXHJR7YHPjLB0uLrDUKbJvPD3JaPNarA
Vith0T6Elk6MdbjjMxIgahtYgI5UZhFDkKM74j/+mBEHQSMvz/t/24rcYnZMI6cUPzgQpIZRQuOm
PMpc3FSZJlKOTM3BgGC//IWZ/Cr9+663IbK7jNhpRjxJ46jDFLaBn8DtkUpypkgLXx7F05gFjXDh
mdx6tfGYLXmEedFdklw4MQqx+0PSClDJ0SslEptgkKC2i3i/7NYYeEMAokvbC5zLA3Ukm/SVup3E
51V0vXpf0H0YoZtOdyODIBD2Aa29khysox54tylzkgfqgjwSZOxXGxLxSjCvFuQp3HxE5QkXMDm3
6/51l0Tfr/LSKh0vc9ewHdHB4rvr3BzQnXoZQ91AfCZIv8MWTHr0p5fuTZetuBZC38z+VXBZ08kO
tycHjoQwpsuh9KqcIit6rGfH4KV/0EyZ8PRXMDpRBBl6TrLcBtZfZQO/Y8dHsRY7T8R4wjfqIkS1
rPcv0ofxGza/PBFnbXW2/GrfnN6x5kmuv7RO/QiFkzJIyoCpdooM7HVo1qyCorfaUBJBZ4J/CK1x
AAm/dqJ2u9rns/7BX9I4rMF3aMA/OyuN+2vz3vCvFuyyzjOyaF485bXGPv3kShFVOmo9r65Et8Wc
HLaWtq4+7ygf1BicRONbQh3yI0rZxRy8PbMOt4kIDccgNyWhSHfsOihaXT6GYG23ka2BNq/hqQfM
irpve+iFNJmlvfzcWrM1EQrfdxEdaAkdnGNO/qLJIuMO+ewW/NaGMqxtS/tqd8fNqu0fM4D/KUji
3YWCzuikYwGIbedzBonptcNKptTWB6p08ubavjxxg4x9jbRdRSi+o2Y2unlzPxA4/wWRITxmC+X4
mBtVe4qz+8cZuy6lPRNG4rHjed1Sqy/D4d5qZPewotjbGIrkz8QAax4W63XX5Ksb1EHRx/wbIisc
FIANJBJuFqysl1TAnuz6fGH5lYJBLdcgtqVD9vsRrQO5kmIhWerX0I7Es5ldx3lXUFYPlpbba9d3
6hKcTQxM5QmO/L1Jg70JlKkbE2901jbHiGpPBh5SpGxmciLxSccYRaJW1GTAIaCGISFRFRcVGVdU
0+o5vNCYOesjkJdbJsr69u94t8tyqwFeqvs1/TyLGxY3yoDZsS0Iax8Kt6wPNMSLmxdG5b6rgIrC
16wR33hg7WXktdxi1EQ7uBm6sn0qPwRwK7Cf6Y4bk2+8x7WzEy6XFWccU7vZGnwXlIzmUsBiQfZa
7nb8vtkDZblPRdAjzFfq6ZMyXXb1au59xkhikkJD0CBiiBnc7FBEUjbcHNIQupXl+CJpBMVAeg4t
x/gBNaH2skxRrCv+2No+TAiYuYOr+fU7VedGMDxnO6YUpWK5cChbXa5OpG/HspMyTkVDqYSOEEg6
Peho8N+ruLq3TFTnFtCXmUeSYqfIWi8GGddfeIxJYEr74fJGj5ehawxSpoXfkmoCGopnfqNp9LdG
sinA81ZzEwKo25n/DV7FKBJ9kAe6Znp90D0iqw/x2biLkXuyyXB3RlQVfMDr3TVUaoyz1Zn/OMUm
rKYfqubyVlezXviedKt57+eZwrm/QF+XQEiWdH+lBsXbV8yhUMx4IAHmspyPXU1m/8JwurYZB7wV
RNUn+et/mZuLrDp8OdntYiTHnPr+RIgGTSVviboqZFvJpP4wNqOz3n+m0W16PlyIIt5wP5/pponO
yVgAKLjlh5S1Huvvz8d57kTmCvI9uIs93qwJVl0Bp2sI4yNvdN+G0P8RS5py9ia9phgkSTneZ1JW
q8GB/FKxX9pGs/8bVXMVHjo8pvBrrtXzeLhfRhtTF4jUvStGS2peL3JZ12wPL0rdfONYNsyBNZoi
agosBlxzJFARiSk13qgmxkpbagm+LjyEfuQh8yVafNJrKFluR8w3BPF9EBc0iJZ4U2lYN6mjEpmv
8L6E6VyH/U9OYn+PZWsHcw2YTNMFSgUAB1b2xUxZ14H+oqd1Qtvx7FdOyKd8TvHWBJF0OYcCY7w6
LSwiA1MrGzC+6BAlnriC2bjRTM7XSdAhm/Z8nOFhrdomTfvTE5wxy6zHtOAumlnmyv9LDqxI7YnF
PVw7SZiotmF9bgVrp0FOqQLa82bMIArWSZlNPRP7DH1F9BpcS/ixVvd3iExtxcUDFdXXSnFH7CMH
OgJi8IecoKh9DOIDo3oHmaisSCIPAzTEyJOMkSqWdvK1i9NDaoZpXjhDOiGw5U8UeIPVhBkYyECB
0/qCaWYkksoSguJf/e7/4hm9Iw0WaKkykK9zE6e2zh7AvVbad4P5At5raGpLilrqIEAZecOqS0bq
X43mjYb1omYwNyOpyX8E2FOAzIjeQ+PHVNJQJ9s5m40qAiGgOUYgsIE6JRTZ/LHqeBkw0LXq1s/T
UQNQPK266/hJW9B9g3mzxSSX3BUzsymQ15IKgMiAkoWwCFsGYvLS0AYnwP9IfDe1ZzTlk9KF9ATg
9VP0WvwwiGh/rEyL/PtXRbta2sub3AeE3gWi3QrsHr7SnvGYPEv9O13JPfm8crUeZW1ZBQTm96cB
dIKLdJkI9TXrOMWF0YgTJ38TFR0N/MWtTbu5sg1zNSQyeAXC051kow91RrjlzRuoAma3Vudd16OF
Dmk+i6gm2QAtxBCS6Fdgz8JJysZRILkJ3QltasTkuy22ycuJInKQmbocOrYur34PABJBFFpPui0v
UtMo9vL9Epg2VwLrOs0KEslIlcnIOgV29Nli7vJoRoJSLpm7ffyZwQ6W4FXlliVGrRVhL+UpJMZz
/x81WbuGKn5WybL+yYOzFDJ6qjV5MkN9OCV2HhQzxAwNNBfNeMrngvS/M4ZH83GggQhXzsPA+FXS
A6gH79LOiy3VhFLOcYOjn/9uqdULvU8I/uKHiGLAT/aYVabumy3bS5Q6Ht9SDbtsKFcWwAHgzDkN
7PVb16MJ2P27oeQgmx2Y/qdo424mU/QknHIXtS9nyJPFUKHVBjdtkcdV7wQqONZAMgiMrnTfhxpE
xSknpqLDnZJwfaF0Y54rCMAXAyns2WG6qfFTQj6T8lKqzDOQ+bCf/pYhyzgTfgWprFsduX0b0D9w
Q0c5iw830KJE85KJ72XehjDRp0jg+0Szm/ppQdrt6s6MkUrr7yOkDBvcstgnvpDDMaRCbvJ05RrL
1KkrkJ804tHLbwCqym6mpbN+CGCwQe0O/ahr3zA0OpmDLVBSqIiklKSdM/qREBQHn1UwqXT+stj5
M0WUc0opiDX+WiTlegtUvt0dKrjX28GIUq7Etaxu9FRDRB8kjGghQpxSH1O4wzd14172cyW8drxi
Wts2QOmgQQ44kD31BitKhTeFSCYz4zK869Dy6cS24+Ug1f5FZhvz/7FG5ASPojz2BywdoZi0QjW5
FWJG3ba2DaM32FYyo5QXaHdpLve3RRNNSKkY6a9kD20jN7gloE9t6J/OarZG+y7JIO2adnmMPXw4
vFVhRLutP/lSjLNoIHfpUqukIYqKEde7jqcjyM5HbKWwokVFd+QdbUAfywq8Yt4Ae384J3RAXiur
UZ+QBBCUSdh5lhE8QzetsdDmeMQNkxL7j6/QQ9ZNNApajb/zi7sKmBORywjUBhIihEKpkjzgFASf
kof/TIv7CDTXpqyCaIVIcSFNQpqRJ7wjtp9cQk4BUn7HBEHH6IoUAzB7+ojcpGM5H45N3W+aul75
WpyDBxrB2lusX6yYPV3NVZdTOjPevWJ0jHHYb+CX8yB2oUELqOJp34F1VD0fSuPCKnERjmhpwAsq
ScY7RpVc9zkncycwQWX5DjOIT2LN+Y+X+PZUWtD0natlw//WrwNf3VXD2UOxsVIjL/MSpODcTCK6
ww9Tks2pxBDkmG8URzWsZUjClZKt7pZi4OevmB0q8Mh9EvPjGSlKeuYEm1ArGKF+L2PSAoTbitd9
Yz6VrsZUBXBXOFs4UTmMy3Lm4wRb0tGwZ94vObXpzGmmLTkClEzStpOiPP73C+wZul988GyKcR1k
7amYw/5IkjubgYJESxbpg87KJC5QKw5Atqq3i6ejCI/fUIqP/5/FJoU417C5eFRTBEKg0vfKCm9m
3M4dzxn3O4JNlm7H609GUv1Z6oPAaE8t2n3sJFupNr1EW8VcMhkVxlQWDifNbrSl85XdcvOHLp/9
jZS8Zohbd814mzEERNHNRxBQurZ277ejbmJCmBbmFjmFL2f8zEiZetYfBr61WBsHvP/zMHgLHK6q
1LxLQZPXIHSDmwuv2SXYJQ5P6OxybWdcct1Gi9g9pme8HFVDHHwMVF1nKq+tVwnmpXs88AElzq8F
1QOvU3qpi0UHs9QC9um1Uk6toH+s1Iva6jXgMctXTvNUfQ9LjuTlCjuzmsheZLZr/u89+zyQsEGW
BY2wkUh7q7dFtMThsPN0l+bpm/u9IN0fGprrloAO+Z8acrF4z80aEdFeKGjjyAi06m06cSnM6+e3
Pt7JBhpajGo50AsM7pVyxmTeAqGDWynVAjB+Kp2mMNA2qW/iXx1zxOHIrgTzACH4HFtc9XfNuqfn
vcpiI3HE6oqHmCAbd9kWbzu+vjbKF0EO0KmEkUlHfujCcT69BxZD8sVBrHqGch/g6wKs2yUA+TUj
mY7jSxsRrU3dCs1++YamlpbwYNuHvN0+MtowNyhzhBDU0hKCMATaaEsQ4pKsnvqqJl+M4YEmEdhi
7BLu4+tPkHbYwC/FQ1+I88LMsFf1Vfud2Z8RZRYoM+YrNEINUHGTrQAvnsqOs32G2+RfYM546T0z
Ku0uCOJvspwop0r6lQwegDjwi4b5kk2reWBW4zPqmanTWnZhZcixf01vvkCoHsNg6fdPV0x/UEKX
2g1Pq8EQQJ7uo2BmJ+Z1q9hhDmy8T5023vyRVKmMJN4g8rE8sCz+t3vlw4mlRKlR5N2WyEZHvDs1
SN4GtXfxZva0dFo1WPpv7vHIvCVmBpGK8yFeu5HsQWfJjLpTcH49JafQ9rC/WhDwIWYisaY2vrU5
duNQSNrHcn9sHPQeyUH4d9XTOLZqfw2MEEsSqIdMUWbodydBiT+TTv4fAUUw1COavAIHHvOiJrsH
yUstwPrt0aGOvlBV7a6SLhbcTxbigQWyBRZ83DgGOkpeRO6mxwdbgXFoAWb0d2XJbA7paXGApK37
r1HY+ASSUmmjgby1nKIiSoxwG1nS45pw8tNxqw==
`pragma protect end_protected
