// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
n71ijifR+XyBHIoruYwYfpVjH0Sgyr49bhZatmHS/l61LjAmkKa6TCT0XxhqM078
+S6/i+w/cnxgIO/g1vnGBSJ54tPNkeR+fXXSEqVIwSFwhda90dCVFQ1AgjHHpuRe
Cb4OI2VDCEq9IK/NkuYViKNyPk678vNjMGV/6L+xaO0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7632)
qpn4yVnPwMm6DqqBwuywL2V5A8nT8qkFxYYs5LVL+jQi1HVQ5PmTNGh2m9mjPTe9
RPNRz2eIkL+f8TzQLJvnttnd65QRBme0qEB2TKX+9aUpr60lNmrl86rAFP6sKy9T
MSGi+fYvfvIr91sRqlGo5JhvnGfp80QfAclGXXnffTPaAo0zg8V9Ky+txYjAQPom
EJSDSegMSCZrnxSNUCxHu6RCbR2w1D+5Wp2NHwf5hE7S/RAXh+qjT2qO1EAMtdQN
d8GirU/0iZE8T9l4Dmyhg+SgJuiK+JAZnrakIjBR5cEDUYXRU2vxMXN++hdRA+/q
FaXKMwMTOYvarsXZFolmmORSxNZPDz/odr0c1G8Kzqh0bY+6umKwkfsgoZHtsNte
IW+JGszNB5uS2FpisXTZwe6icY3oHBS98uJ9H1RsLnqLQTXyCgFEzc2RnAuU0jGC
/MhOJS4HKeM09ftJpUDOo1O4wxHDDXTiy6ZM9v1iShJyUt+KHAI7ZCCYPuLiYaSc
/9gemwt3HRDEzFIpa9wOGcY2Kd1bk6OHJXm8+MeaHfwDxq7NwOBKz5SriX68gDb0
Ji2c43wuMxSA1yASnVKLHDwpobJr9c4X+6Kj5tYVoj8qLVA5TgdVnLdxkJynAV/9
E1VYG/32ywsc6NBfvPXFyYPP0mPpmpkQFQFCkA68EKEH3kpJ958T+7W2jhRghkcl
of1/+75A6eRlJdsTphl0DtnMlLbHx74Y6h5qwJZ3aOUgpoCTz91PWxS13aeRqRj2
q8g4KQRHQOhgkZUDugo8P2mgapb4nrc1Tp1yj2gn/Q6GYwPUt2oyeMuVe+2kG3nH
ilqkMaI3/6t69ux7MK8hKqwYnFZaAct4FHtl9XslvObJC0gSo/Vs9dicnq5IUUBa
+x++qjSyYyWyUT6RjulREpup+6gtrOTl0/MhgJRcGlbORQSinRUuIn3INSURqazJ
IRt4lPqPcc1N50VQSIuSc6Ks6yo0/0g+Uqwkh0hOMkbpw2BQiS3Q6fjCivh5qa7P
WTvFyNrAYaRNk7GDJSf0WIU/bnc1asBVR0x94SmRCBV/pgWoXs/NfRXdR978dDXB
LANuXihkgdXl07oywb1cxhoMpH9DMkW7MiDSfjQq0urK+SxbKvBYlfyoQx+yrlHI
Oy6HDLE9snZRK7y/IXtIAsOBv2jFQ7xnGxUvozFCu9kKP3C2jTmG2NW6bFslDrkm
CnOvk1coYLwBjsYq17enoLuGausgRhHCPN+8GknoSiDuUmbKCaZSEYR/8RB5TIlg
xf0bPqd4vAy7CJnQULvVFPqxnbz1Qr39eEGGzOFDrkf+B3arKfGwyqoI2fUBhqcD
gcJNFmNRpuNVqcH81KOeP7MCqE8N8R48Znpfhw7nPNJOR2OJlIpuOiiRbxTNuORa
FEb+Kx+zVDwzubdMsIbt1kFzBd5B587qKzoDD9sUSqxp4WOAUwKoVdijM8H0/+S4
2PlUsDfr1BfbcvHFWMHeRFQ/omAd9BQtIR0KzSVIqkfdBTXQK6qwpNsmVC6Dlyjz
cd/zpvwvV66tP8ad2LT6Ds5OjgqeXjDXXlLs2zeuuEfaL7Hwel5Y6dbJuRbHrJN2
hxwQX5IUtFBpUy3yVGVIfu+7jL5wYND0wkOXcZgqEwNXR/7vZ0fyY1nN24lF3JjN
yu8+rfhv5Yv2hGp07bv2msc+85DajmPZoAv2kJyhgNDCSVDl4Tb5gl6cRB5gDZ/w
VcsPlD4Bkh5rzr0otWXJyKmF7/x9olS7M3aQyiP7d/19OHPCvcGz609AsbaUoRj0
zpBh8ydHsdyoci9GTVttOtXiQPJrsFrNzTRHc9uaHBJ/3pr+Vg95xwOluE21cUzs
84oyeZB6IimxNIVNU0Y4F/k5FU/MT4uBJwOqu9cddR/boqcgoQKcvAW/srgTsuhL
U0yNaE4GZJc3N+DZZCanlWYmNycAcisSKoD2CHj1KciTDh9BM9YYlDPo1nknqycN
FzeqxKnW3rtd1OBfSNcPQwyA8ArMWujPKuHrBL6x4Qow74sStnyi7mZ9i4+uiAWU
of1BGlUSpL/A9ebBMCeDVPvaDdgu5MlgMwCP+tNoCnRfD1PiFS8oh9w7qu4wsqGc
It34wSf/GeCGXIbHZmG+wdxSPD6LhY0mQCrnyBGFWk2FPLf2+uUx4SyDJUMWLByc
rTynQEogdjLG0etU08J0ZsMUUzU5YyyrfQPVz85OlL/9w6gt50UWoLqtyyX2vZuk
LhiHS8ljopeA7TCtFLXkkQTzAItxnnt/TvDaoZ1BTuWSCwmLoHFQzuhR6WKTWL1c
o5qtd+AeIxNoV9X5LEPyTs/Onc4KH11UUcl1+X2HnRSx76/K4ShD+xQAFbhJ7P9Q
fJGWM0rZ3TWhPWRJjGnFHxifrBgA1cZJSgx1GhzEbNl+N7Ssv+itmkPjR6kPiM33
2VQle7q21jg64btReoxPjcY1rkhgGfC/zGQlgwiD7lCv8Amqau6Ve4Dsu+hbKGBd
tuEQP0ptV0tMccPmB93X9h4CJZa3QytVnqWEbjoi6q+/uGkJ1Vlp2A3IKsARpJtk
BS3UVLluR77XIfoSJTR1dhwd024wcmFaN/Unt7WlN9Wdus10wRTqPC1VNDGQ6Szw
OQ00Kp71Lr/SkGqdiK+FZaC8ywA78I98VjnvQdJFSF8Wm4vnXNfueXTTU1FhguWZ
M9yrbGPomG1NEBcJqVLHtcUSM0nPQY++nFXFYGRvDpYyoYqmWirxsAMXhkPAX3yc
Y6sbt9uOS0+nfPXupf2xgyYzKxh/f+Lbp+nB8iZBZsAmmZWDq6ZzXPHwXkquzmg5
/q4+o4l+5XEk2GiMwT7q8tjvswTTNJGxJqGw+6Hw2tAdWSIMEEcGMUNEw5af97AP
uOXjDzBp5hyypeLnLB+Cppdr++pn0BXohlDP+pLAhkhJ7+UVzRbJooXBKvCIphvm
5A7WNUya1ebfk5VYdIbQJ2d+hJoFJq91mwzlFu/mRi38H7fQtHnZQCdpwQpVMWKp
XU+IJZqYvACq6hXFSSXrv8aAcASveDfwC+RdddEVEBEvDUP7ltG+jvQBvJO5c4G2
w6nxXd11CTUR0WawA9BpQb8UySc/iT18157KcHDNdfZ1S0lzUJWQUtM9+mSHHVKX
y4OlJ8Vh2IrTubHEOCj/2FvJlfThjs1dX5bBNxiX2a/9WlDL5HLCNRU4j0PIAf0R
1dIIyHqF5D/n1eFMjMTg8zLvwO/ABzlY0k+9lROLpdRILxq3nL1OFU6mgt2kUYIy
K13ruk8Qv1Dv23Je3rp0DWD24giQ2eLGxVDyOLVP60tfXI59wXlLKyrm2Xkj8ICV
A1HfLpQwvdyVV8Da2H14pzQ0sHF6vVBYKLeaw5Cw+dxPOjOSVv2L91vBvJOtYDI3
ZEM0Op71xZ6RDDj4laQ1KiLWToEnpHCIT+7oqZyydy7cnCZPmaz5TaX7U08zqqOQ
a2eTzQ1ke3/wcY3iHyYz6SrQmdc46EUYrz7djdpLYja4W3h4vscnAymfzeG3uUZY
jqpBQsIpHN9aiMZcoKFZkaIRkNLG/RSU+JQqrmc5F0WGvWuQpsnA/JUOHjeS/xKg
myDgpOILCg2qPPyIsIQ6z7x8Pb3MAK9k8FDfoZ3ZdrJ5Oki5pWHI4IM3AG+w0jBz
onSnNKuTvP/A+CPqvD0OEJRIvsNTqCWDAKURiNnSWsnKLarXGnd2sRhwTfW+xDL3
kyyeLz1E54dbc+4/gj2qL+IQg1sY4XkiBv7hMiHGPjL7f0wR4cPx9YfcZwk/ieoS
qbVL33xTCAPRZ1cqiATC1rlbEWrNIoay8AzJZD31wCp+b7TP0wa6UMAInetsYVjO
zySChBeznlNluzfw+RhjSouosr+jLNO/k9OJlx5Il3mO50pKLZyxCfa/m8D9BiEf
fthevh/0Ju8wkNs+mJMBBwejmDvOTnmSZotaDstsV+f2e6jZS7LdOjv430OoDUVQ
SWymGFsFKhTc0lvXga8QWVlLss/u5pWH06Z9Jwm4ldaa4X90NmzMGcUhcmSi1O8Q
4QGs7zWWwtJyAAIg7ze/3Djzo7dgBFs/Rqs5g38L9raZdUOv+QtdIIDZDNCD5mXL
xTedmL1b/gYetqGOly2/Cg7TNId9KBv6IFQVOHNdJF3sKd17a1BB/SAKAfh5F4l0
/FMJ3v8sCjQz25IjeFtaXKQ/Fe4rwAVayKbpdAhCIbDEvvfBcR02zo7VpqmGrYvk
fK7ceqX5vSFyBk3QrTXWe3vgY/lwzG6ULCSagHCA1/HRHSy40XvyRxzzjob9ojD+
bXkWIjLoV1N8W+nvvgNvwbEp580Y3YbPQw/ubrOGzLfc1RR0Tw8EbaRgWxgnZmoG
GFOMGv1pdXyvrEVz/sw4TA0yr/KPLtKtEcquM6tmwlASwSwbpeR8fpzaG1BCj8th
SMO34zsLKPcoY8PYgJZMlrDZ/swY4P4+adhlNJWEKap/SfSLn7N+XI1QEEup/L2K
N71V4YTY+mFsS9mm/NEFl7IgV5XhQMBytBXbxpoXeXDOOtkyVBURZlpZ1w/EjCiq
LXctLDR2lzDYUfwFTKzpVjNy5zRcK63PXMByEKmxJ01b6q5uQp/SeSKe7a+uXzGA
boPE75koTpn9IeDkgEWy1Yj6c0o3gOnv8GHvvJPI6x26XpWxVafi2UJ/0vyU0lLn
kb0sjyCND2xPHOnow2q4Nq0Zf6TlBpn4K3NLpmlBvjFQMTUXq43waUKsTX1Th9ck
Ua7lP50bCY3rYEifld1CkoxU+QGiVWcRrneoOeUdf9gfAsyWWgBq13Fh/Riykv5j
yFisLeqQqKLN/oYKZEpWuBTBmuWNe5IUMK33By3noNXOoKnWiHR0q83d1pSi+UJG
C8iy6+thyq4fN+pogwQZA3+0vURmsofel631BlYhIygLrLzNwbbyNm9nb4UUprMz
lx+rcFq0wVxJOSxsCiMqDz/+t+gTHJk0228wjKWcO8AfxzjBOHRr1qgfQTW+yXLU
Am0ISa2KwBDiOygjBMVe+k3Cd2+Jb35UA6MR22fEvDCf1AdVmCuOmM1x57H0+Ef4
K9f6qWwv3uayMeG/AhuDzsmunoC35/xdcPhmT6XBVIav/ERzhgSmW2hSnybDLJ0h
PT3hNXf/xStRy9c1m/iv/yvx3xNI8lX4jNQvrKynoCFth6o/S79SfgzbsZVnX7av
fFcJoE5iullkoUpQqJfYcXpjtQNyIru2ays6BJxZHtm+G3dFphtn0ofcpw4iiJeZ
Nx3Aypg3X1OhcGvYA1Q7h5u4qBF65VJeD0uWKNXEqiPjBGXYEu9slU+gl7bbYD33
7ETogAc7molix1DqIpoy52aI7Sug/vSUOphi35FPCw2TrfKM/uxavBJydnZd2HrV
w5H8vzoq6ALfM5ISgxzcB/4L112Xu+Kqph479tgfLofIwUQMBJmWUOyeE4I23wVr
be3WoGYk1ZT1JpRKnz1aj7BTLjX84L1xfXizekSMXrIGFtd18YQIK7P2792Gi3er
DTrEw+G/fc6/iS5/mTO9vbWBGjU5yZZ2HPsLv0nw/IhLuZ8x4KefpsuRw2icjkLa
iOqDz0VLDCX9Q7/d7USqzRobRaHllVb4A4ppW2aSdJxbovHVTj49neZw6gxg5MLY
fvNRf6xiClzk57SmEFrT1Yz81cquZZUtvB11K98rSLKRehAev5VwLMWnP5AfIokn
OGOILrMiiTGWG8MmFcGRFtu7gFAMCzPKcg1l1u8MBgv71iZLfeAfpG0k/L/rqH8V
zan6sR35QVPK/V+/Mf/y+1Wq7yT5apBTnCOT9Kkiv+Zg4A3cXoAdDmk2/rVTICie
+6WD9333VaDUKmXxYY0EJJzyNu8sFZjjbYuuVEyaiJgM6OTg3FZWauigUVq6axJQ
+8Alju+8bFj1g5AedEAeKfOLwXMGPmmJK43uNiZhgCO0LiIMLwU+EU6bOtNZcQCa
v78tdaaDKQ7x3eqsedMrXNPq0pEW2QPYB7FHw4f7NoOZ3yj92wPNuW9lvQ6Ggn7X
HWArJmr/9ygAph/pjKUJDhWM+eSCNrc6BH+1TRqmjBWvZ3N3ZeMIeF2xM10wstW9
qcRbwulBCRH1VWic892UxwC19auMUtuShoBbNzI4wDc3TfqRDJ2fsEI1TLr3iPM7
4MyK+q6rLkw1K7otzfdifY6XgEXU6FR3Tc5mk6QKCBJFQEYJ4CXoXMRiLm48+Z+t
gcnGXyNLZ3OKjXCn+UC+e/6iiSXPdUkT6waGUR9j/0GnVR+p7xGop8D9vK459mpv
sZw7bQ1KbK1niDtuvNRGymdeJ8H5hzhfMDRsAk7ka0sr30MRuDFpTgYX4DrJdTtC
r1gItSKBVZwHXgLdf+e4inLg7eFKm2rw6ZbPXqyM0TKblm0JfN7bK522km2zC65x
VDFthq2AP8uSTSfdUN9eMChpCq2WglJtQpAyvHt0VL6LUQcp2H/FL9gGyUm/4YXQ
wXCBFLTABHIFlj5HuZfJDI2mBjszLTBEt569vNQ6xEwop0qxAtPVI1FlwKepiWdV
snwo/6/aDv5NW5zFANcPSigxP24UYhN9KHXfmMMKBgs09mVz5YFGd1M8usOmKPLW
YDJ6lz1yuG4Vq3udFlRM2sbgsNiptmZwYoipxqGcHEqPmPx/NZXjfolisFx9kX64
H6hu4SDaAeS3YNdNoMyyzcnAZvZDYTrNgm2Rum8kiN3D72yH2pa4TfJ2MLQFeFx1
AplqbN8KQtRLSXwpOPxvjBzbEN84NpxYQe8HVAWaPOMWJKZ+EiPeI4FtvWh/Nu9N
yhtXTv3g0EnyOvCk64LvLcv6+43ImIaChg/SGpI618ECiavgNY9qZstM1TNPKm8z
mX0wCmmh/BVsYhcOOgL86mORlVq/LShmvUHpKPms9o3H0ykrDkymJg5z7iUELmtE
nQ4B0L4grVXeDVjXIGlgQbVSDipuoOPOUQMX2ML2XNYjNm8DBimBOgOsgpX81l5f
uxx0AVZIp5e5OEBkfWkHIt4PgtFCglfl+joQxRCym1Ve6Ml9p8JSAVZ1oeG7W6e2
wdqcfBbdjK+C0wd6fdcaAxM27xdhbQKb6zwsxTWaQhiwRX3VzSXonvp8nk9IeYUe
WgYPRHa2g2ZGZmIQxe5UByUeMsZRumBtWCPKGpzxuuf9UZAMastI4K5NIw7QcmI6
NoUeMIkEn1P9rbmLBO268PUMsIUaPJuHi0HMIWsKat7CMY/AwqrislxjkmWJPw14
U7hNi433Ug45bN8wMzkYrS11TeoMS9tv89b5hML6MHEDqC/rwR5CFBVogkyt6Ndx
mPONX5xPZ2lKdysVVVtNSQ3WFPaEHNBlOVWJDR+ZGEYKZuFfRoQ8Y7B+1IrcNtiu
NXvfWOFAm/g/1INz7xtbcJIFBPHj9+jZrMjzVJoxzbk78I9V5358co5+l5ytzpgB
g75QsLb934XHoqnYE68Mna2Pw4g7P3lNJfWXSxzVbllh1PaegHj/4MtYvq3uXxux
jBi2Rr7OEF42N18sjwnxFoNYRG+rgjzujFMXQ+OkbPmRWhSx+RAm94ku/HQBLNA2
HiEj9Uv0LBklPhyxEBjtFgmKaPdOUwD1zSUHTTUFY+yLKo0rSAOFyONz2Wm8VWCs
/eDw9inIMZ5b7tVTn3wIWHFpNdGWsBrEHNdO8G9BDbzzdABn4DVo5wLT4KpHkPxL
EmOW5bqa4HyHx7wfm/M5AQLOI48k6lNlCHAiv+OhYP695vsQkP6v34GQKsyH1lVu
nwlabLgn040DfHy5bYbb696EXUx9zKMTJQ1t5uExzgNgg7BgEmqYjSUEKoTcSkmQ
Lngow+UwkFCG2sluuvQY1sXQ637I80sx1g3Vs+L+BkZj2ChdkJZHkBMvlmhGLQky
UNYZ5x07ioci3DCUVop9zpQV0wzx/wbOBWo3a3k2E3HiNWr/8O6eR/yc1I9R/rAR
Wiz8ryPqqj3sldCipaOlQnRKZWzVBXDCtENfH+pahD6H8QiB4Hfn6AkJOVnv5FMV
/t0+0ipsC4dw5ji3NCn2QNK74WhWNO/j+UlmZszPJfd5da3DLknz5JHEIYoJ0Hai
X5dceeHq0Bn+qbAlVAkc/Kw3ligXnC2X2dtvoojaJk4h9BZrOlPgBSEOIA04fHIp
auwFFJtSOTSqcCZYF7Am9lINNBX4FY6KLjor3gGWtovZraIVK0H9lAX0Iv+6TNb4
XnysBOiuVfT6DAPmQImEkaQXm8w20SOvCGahixTL1RBBcIHrFJ90MMHunCZAFvdi
XTzgtM7Sk/T8eR3Ku8OHijQBOWbLB5U60CN18kfHIXSkDfhIBCnP1sEjR5Tv08hf
OTGTnFJgn9zIZAe33G/ypVdN7/GSm3dcUm08xb04RktYr8Q3lmAJdDyXArWgZp55
u0ua97NNVD+7t5NlSZv+eFWk7Is1YHKJ5QuzVcwg0ZHAxBDbmjw7ZrI+sMb5OwsF
meVIlxUCvsZkI+HtcP/khclEgmdxf/9Sy60q8m9JdIeNsHU5GrHsZjBF3G4hijzX
YqbOnRfC1dcEOe5qHBvM9OM9p1nuPJdf4Hx3VmNsUnO9569xXuWu1ctRT1m/v/mL
c+GdyYSIfWY6OpgQbS6rjyL+GKAX7FnJ1VG/KaWvsP7koFV5/Hf0mkqPKbIkxLd0
i7BrL+m40fKWtGqLyF07VXPtHeG61JaLWXqDfLQh6ddo6wB9RO8RuaNu5AagFDeK
xW6flZyN51Nr/HweCIYj+rcyUCnLcoLKuolNt5WJ9rzapudi/qtk1dOnOWvxsTRg
/99+5UWQsSQqIPLe5VrH509QVgZ52zkj/Vy5ZtwfTOeNgEqTIy1pvOqq3Xxd7qWr
dpN8tSenmcSc39c9G6uIe6mKzH6QGPXJN1TrblCoYnGX7iQLWzgrHhuMk7qEVBKW
tdFms5xN6vq3/WysT//PwTzkLetvSEqcXj7SVpjGCoCcqOTeWIuBq51PPYptXxmq
Q3lK6B2CFpcL26WPGfx7zW+V7zi2S1wNj9xwqpBp1b5WsF6KUnzTugweZQUTUMBA
TW1Rd1af4uSXfuetYsb9I/ZkAeyCHemdtaJ9RQ1ae4yuMY9AQHDcd2Ls7VAwu7HT
uUPC/BhcDaWVZwjSchWiQNW4HBRFWKuSFCeW5N5dh9Y1C/5IU0KDHcm6ZzCG/vnR
Ou0PQlsvcwx3XOWm8DxRyZPNeeT1fOaQlN47RhVguGb48ZiEgFn/akOKecYb24JS
FqpFQDPdJ0l4E6FKxERXlNSPC2onjOuP/hkCukqHygB6E2S0sqht7slXAZe0+Djj
YQc9U9qTNttICY1b5yIJopkAUTdtgfyWupf64sWjV522F4kXGmy6Qc7KOKOpuODv
E3IS5HY60C82nvognQ+iveDd+yInSVlOdU0L0VmX7kenvM9RVAHn5ko/FJTtSLz6
kNNeafzKQAYS/IctQ0i5ylDNAW5wa/NMA34G6OmjW9wicOZxdrzf5paaERh7XqtV
z4pVXPOAqn7x4wwFc6ba1i7yr24BBf2A/Bop/Fj0biK2eAtaX7sp+jh/yUHKIfdm
gp6JHF/WFcDsrLen658ZtXeOWEDs/wzcNvnwTeKQdKeHogyHwAwdB8TqFBNaboXd
n847mCwAKLhd+TwrQcXBgNCZVLSuZfD01STMjmGISWpEEFiXSIiZm6oifMkLQs9r
Fi1uBith2E76ujCqyNuTzlBYf1BLGfTGLBrvAD6cEqnUQ9txvflFMXDgzhZIoDe5
3NWkvIN6uK1NFgRVrKh+QYPqN2KAevVA4uROiG9LdWT5rCat/z8uCx9NAOHy0BZ7
TUT9aNgjjn2+SX3NBmgcmqHXRgI4V1mkP0JHiuMvAa1yjy8p68wcF1eK62gwo7HB
r6muqSuYkPVnEVe1zKW3Ki7rsC3Nq4sb+1JBoGwtUO2gwzhmQ9wCfynEQ+9M8YXG
OWKlQAgpPShBBWwV0sQks5VkalBLM/Ev6vIGVlfa8i/ZEWDPsnS83MhdvAt3hp0N
aToILA9YkH5b90ki+PJoYCrQLJBvC7MRi6nQEtaZiR3m0lapZrAfjxAj7l/zm5Bz
YCpEz3iRo07r+KRdJoIbxn1IzI8lZxBJc966fVJc1TljL57Vx6+EjgR1unQ6Edh0
xuAvswJvlDy1hkMPQ/xQEmT/jLwlzNZgyaSFh/UKtyYIi6JL2LRvF4/HSfbs5+qb
`pragma protect end_protected
