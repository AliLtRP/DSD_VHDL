// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:47 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
isEguRW63jWtsxh41pU9tOvlwz5bw5oUeM94rgSy3IMCtxpNBDpF2f+PTzQvQngY
jyaK2ioLlzg1OAMZ/BbgZHLC9Ctd0N5bjVZAaY80q0dyJmM1H09V9mBDfc8AlDVR
7+DTDEnFpaLjwVwiCSrRw9IO593/u0vXVTA6/0jGe20=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24192)
KJUvNbY346oGlE5UriKUtlp3tHXKB4mpScWiJmzyJsEP09DHnPftd0xdglIayA9Q
g+6843o1zz/Mgd1dnWuHtDOT0YLF/8mmTlw15eMS4pAwWsxRWJDLg3KfN61Omaij
TpnJFqRh8hj1+kpPsWNBU2IRP224A6VC6dMPfu56qDSoepxKObWBMjHO+BceBlLk
gn47cvn0NX8f61VgxONn6T4+rEUYw8oZCGFFcqN9vx8IwvwhmS02lHxLj1dJgTnU
IhHRC7prwsZGnoyyjMRPOG8KHksDXdQPgaqqUOq9fpDtknnfysh7U1GNNpmkTrvc
ud2bLytu3xMZZj0HG4avF54m4tnlHK1akOci6TVFZ8Qwx6nbdWvumzQQUKGssMhr
Bf43epd45BaZ8+Lcu37muiuGpW3Wj8UtX5R8Whcy/KiKaM2k/iAU3ZGLH1Xf1yAb
tNqh6BP71poqe24fAFIp8yOZ7iBr6lgfv/EMoAXE6kFKoLRLNR/dkKIlFiCUjlTB
mHKcpcH+KZtOZ8jPo4j5wiBL4YkM6b5TgGr3rrWCfFnd1y4f9CRVr5isk8BKaBTN
IQVdo9GA20f+scyebn9mrxJ3SpzrM54CenS0huK18W1w298jg6UEfgc/6foh9c40
BQoHt0d8AbR2xPMgCEnX1TUzPaEOd7J7X8LeJGG3RhVyOS503wo2vqpCRUPBDSqU
uk21D/LRk5ecYz48lVSl9vBuh5Fnh4d5LZGXex4y6EAaFCzr5to/fP8AhR1RamAw
8BtrkAZ3z28qletSS6uK+i9w0UDk4UL7ubWapjac54B7ololQbNxPaMvpNoMWZAb
8I239mgc0OGzyUYmZQn8XZc9+AIMk0Ld9LZNFTfGGx4Wi52Rcarkh09F/0fYiDEK
IjFG4PA6tAUp0nCih7OZakqQcXLExifI9Azk47xwQmkvKB1vsR7+LGJUEy6ltMOA
cE4slMU762r3737CkRfbfdYprYVR36ZEkNSVOmQJgnt1mQoNzDW3b2KxHVUSXKMy
KE6aFustIvUrwIhm+0KuS9PAHdgyQe5Uqj4GhXPx4mBx8b/hR8Ls7hoBvR3xHkEM
S0bhIWCzdo3YKkZU8S8Y8KMByCc9zy7r2kkyNOs1BDvjn5aTUGFCUiJ79y43u7Zl
ieYn85bVqN7OVzowrVFx1zVaMZdtQ1w9OET1ZonOf8ibbf4H2jnX/EPlsEko6QPI
jOPuxltBp4VQcIIUkFp5GVN43JoqJHIwkE+AXDTG3St8rdZ5ASLVM0M+ios0Zr9B
7b2HgSNGYkLlwpvraHyRdwZyhlr5p4Hkbk99GMMY0VEvWP5e3UFW85MpXzjtYZGP
fzi0j/Pu91wM9E91bHv3/r11rL5hStZnmwrYZKLxRiTzjspcT04BKsGomOD8Hctu
vUmC0YahQ2NZKEOOgVk3NBJX7OPCJDHxwOY4cVzKLE7BHTm4aPHWSWMf9Neh5x/f
SpzStol2dSWnptKGOClQYEB2w0b1D0y7mezlS9ABKZu26M/zQ5+lycx/Ja3+op5p
VyaoKitW48kFF5JYhTHCI6LTGz2jIqzoHrMoGK6cfxPvXyyCqyEGadHRQzaPI4RS
r/Y9OY1S0P08rr0xKPzWN/jMYXkiLCrd9MGVnIm3k+36EUqctMssrQ93G1pXFJjr
BRSmbYHguZIRar35LDTUK336xE6QQCoeI/wzyC7gJqu5K7Bvxp1ffhaXrUOd6iE+
0sQwRAkVsTrIROIvpD93cXJDe1TyF9I8Ex02jZjXPRE0+tkuR+/GRYqjkeSbo/5W
VWeioBzGpwChW/qov8zuYer12hBtM39BjJpvIMVfbkyunHM6emXC4tfXEWiNmFta
qSoX0uMAkYNgE+UGuYdF1OAyqcJuYgiJVAsTu/6d2R1pJuCcIvpedMtnGX7/QQyz
HHTKU2m/JMhIteAEMkU5JJvum5T43sGzokQr7ViL+DTJ+iPQhkwD3BRZ4l3nlUAp
+JRh5BnIeJ5Lv0daG3tzDDJamMjOIQ6oLohNfHkbK+dpya10sJjhFve/2l7BniQZ
M3KKJYhB5o2/V8XxCpKi3ji1/iByFt4GSLljlVsrzyirYRKZwlQl8c09DIL+qX41
zYlceofzE4X5JMMSPxGXzA8D7cfsL8yam8QnQWqbWYCwDlK17RpQt8BIpcn/rRNj
H01GUhVOjntmbJIwN9ohajGTcFUBZxiw5JPPPatHXHmwyZ9NtBTI+OQI8ExQYAfK
K5fh7gLRU6KfEmdRyFq1vJjnKyL3qI2GTa0yuewbYEn727/bsb8idZdBMEp6089d
fSiCvALeJwLuHucU97aGWo9pRPZFnxVmIah7uW6QMTK1OXX7S0DphrQhhHn1Dqof
TOjmYYIFkCZzefL1DDdy7gqHQqo0hhGhJ2baSRjh/mIiEN4CHySqV6oTBipObXAB
tk3efA9P+AaUTrlqefzUbUyC0K8tvBL4cy10EVs+936Radlpk9nR2HhaYE6HMgW9
VKwZHTZWrG/ppww+uASZAuF6eAcDDeuBTK2CZIDA57oXwFa5SwYjh8jqlLxYlfdk
BhYmNtBXgT7bV7ZzIbGQFmcLXHW3HLUOVhRlj5JZ+yR14gEVi6vCxCrPJzesMpqo
khypWJ7mjoD55oPIllG+KigKJXrb1pzza0OA6LFDEeyeYkD+zFLNV5uHJaKaSs9N
4uXYN0QWJm2TAG5SVaq8d3QDSsOXzPDqJaBgpzgHmvKdWodgITrWcaG4jqV0dUCL
UnD/41IrY4dgpjDVZhrt5IBWxI1zSL1pvNoED+aI3knwFp0FTNMwN2WAs5Ngl3fG
VhP4aZGLcMspk1sm+3TPJn/4sUrV3QIkBio8pkb8jrc9Dy76zKG4Vk1Rwv1n5PTN
6a8gFKt08v1cJaA452EQkiq+XEAoUB8Lz9E25hArw5Q4OyjspPRUq/Wz4uiDfNPw
Bar1sqb/jkAV/bJWYUMf00RFlTvh4idwHM0TVWpgVTrWR1zECuiMUcoDk8AsiEC8
nqlVrBAP33VE5DSqNMbR1O5HcfCSBVrHIpMKZKLpRzDhjehtjyg6zMJPsDOB9W0+
6NlYorIDDsoo9LtSoJzxMq9gYkZDS5WqwbqCL8KK6455cNqjMm8ABTkSTwfyEoOI
fCysrxVlnpaO0wFZEr+3ZDGb7Cnth3S7Wmg2IpWOnR8IhOMG0x8JM0cWDx2Ruq1P
+Xgezi5+/R5HYClrKGEVfLKma6WZ9yT5nM787asULgR7d1dxrd6J2mG2T5rTIDjp
QkP5SG+ribcwXu0b4RXA1a923q5oB6XOO7DUzmy3cNuXBK7Dd4CuKdCrnhwNKjos
dLSUxVnX2gcDW3aAVp9V9WLTGIEFMidU2sW9vQqAZ77gSwhvG+1/3bxK0MtyEfhu
a4rq+hty2ZIkbGFnwnUTUcEdeEUxBYpq//au/kusi0Qnvdshm/gNYiU19XKvmNeZ
kdFGk6Hsb/FdALWJZuZ5UEst0aQoWar2cc7tEo/dy3g1w3TWElapQmKdVew0OTuh
Ke4H11+OCwsil9xJ5X1x6CCT47SXHR4kkF3EfecElc21Ts6RwmjgcY0UHXSWxCPv
URdMzF1eXdZRzicHrSqFfJGMU3MhPr8CTK359OGmNmhesg+wPRTj22jeuAEFblJf
EZy3DOWDuueo5sI3yKN0IgRQ5wjiyVNODezITR2c/ccl7CflVpE+4PoTwUpibiIY
5OFi6rm2YPJgjLYvAWiHhsVt7l9f8Sb77dO2UX25YwhkeYbW/XMf/41e4VYnW/06
I5HmddXkAJNYutr0MwN9tK4uVhtzFQarYytJUkZZfzCgz/Nwdoo9zk+6wbBH8iTO
dWcf3siEZ/ByWu8htB6vZkZHypLtPvb99N/GOPY7Mg1He0OQXA3Z+Y4nLy22/tnJ
GtWYGMANdkcqwQu3BUw2HOIlIPiH36t25zPCRHLdM2D2fqetRWZShkdrEw+7oZWi
n3spcXNI3EmEixicmtzimMOqZ7pNPpctVVxzbnqpbuV2obytPO3NtLlZw2KgENVN
YPRy+HvnC58BOzYDh6ld8TSqdGMO0qIx+nJ8B8v5UaHPVOGziva83yWiprjomajy
km7vPLg7yP745kSA0SnMbVUlyFwWIMLikHcdc/KcXhlxdSHoI3kOXhgeidjdeI/h
pQDW/UT3vJirC3a4Rr5tkLzhHa4er8QqN+ofK/iDEifCgbdMc1fnrb4f+i+7mXeM
c7+DAN7CcTOZHPQgTq89jT7Te9nYo4AH8RhPXKRka6erO4qJWNJ/Kg0SzuUJsl33
I2vuSVqRdSdIZHdsqdsIP0FCOPav8uYL2TqJvLzXvawN0WnQikmx7o2DqYADTGc3
Blb2g4tMi/G7ixaJIUy3P2FcwdYo633dMuP4dODcqILOgVmrkxgQe+yfsQ75yu5i
xexxl9W5CEUHkp+cGnKFk3XXc2u8rL5Q6/A6G4ByiDBphF1S3g64M+ka324sA4nE
7ICvhgjBnrBI/lxU+JHyD5MFGta+Ix/fv76ZhglvbpkJfQajQLs4fblfHNHiLLKr
Icja4ic/uB667ZOWjLT+3f9L1dzqAHV7HCrbT7rEJwLL62UiW5S1mqIqWMUMBuS7
K+AKCsCEn6GGOeVNH6Jf5wy4OpAl2Sv7hq5XxgddIrFUoN3lEzFEtN9huZ6b8UTb
BDDqIrliHkeWUPOVBL7jP0SNbJagKDEHh3q1GB1IJTwEk7uRO9rQor5vc+YawNO/
NRajpNaTh3RdH8SjAjFiLzVNbcIcLSC+lEyQu3VHaVxn2wl0bJp+XZU156QoShaZ
HCgtG/rKQt61u0itw3u3Jp+yGCMD+gs8YXrKdBo8pNnBQ/dASHi7M+YGh+3ku5uI
kKEIjW6mdmgL8ys0zqeumQ7jdj3I6R53QoPcRCkFrVeEn3Wb/RAkm9jTLQBN0Evn
ybRzwwHxMyHesK3GfPOcehAg73FYWgJIRBQU+PXT0zHSGmErE/06Yr9jNje3qyjl
cyQOg4woeHyS16+Ykc/RkXOs2PKle1DQtQfiOS85ceYqyvE0b8986ovsoTcqiXT+
+vKuF7NPnHEhUge/3cNkYTgUo1ULjnyi+99Xran4Ygzbw1sa0v+4UtHe6LW192YG
FPT539F7XaFs+ofxQKCSY87rhBzOKEpq/m5mnfETDY3fqGaqjJwgkwaGcAR7nqSW
ZFx6UvnGH+Nszj3q+WzCd3xZmsLUfIMqYrKQXe+Y0oh/L/eWaKIpmiWezgJf8gDu
9QDDBztReA+07BS8GmVbKYJ9Tpr3VhoS8qTDjQTiv6GKJHvLqqeIgcH3wnhriK/f
bve4X2aXINbFm9y05PJdHzaLJNwKVQAeBkAo2rEQBHvbrImRKQKocQEU6HxaQ0u1
WhVVb36fHQCMuCpnKhyTB0SMy6/RFTF5JvLzaw5iAazw1A4Lq8R2wnpv5Xm8d67/
UyY9ZC6jmbvZfNkHf7aO3meKqU4qCmDPrgs+y3grBNNDyTO01ednpTnc/nGok4BG
HRpefTzqoDOvsN7yl4XcfpnXqrNhtjPQePjtwRq3mOq/TK87lPCmeQisnowbUAdw
R/VVutoAirJUevPWQ6qZtoIqv1BbeWGkTqsAJQASsPbNc7DRYlBdEeffttD3uPMn
6jWWYikKyDdHTbIOetyROq663yw6X6nn1aUUytDEURQJuyjk8whpFcIZJ5fhIw93
iqFoDT7UCHrcrXXAzzqB7NQSLrkanVs3WXO+C8kRk74Luy3WGdSSAe8CiHJJLjDq
6HtAAad1X1TDT9901jXl+E7fKqL/YA4ZgR9s0YB6uAj4yEEBad/uo/mKp11m2YHJ
iaq5yFUAOQQ8vZlFEWGZ0NgaleFmQgr9Ph7l1aI9zl/Spt0UliHreF/MjRebdU8P
Zungb5t8dlPiEwP4ZQnrM3tWeUFXzqDcn6VlOO0TgEKbz4nFM+zsREDi1BRH9VRh
GTmJC0PyiBbTGENMTs28HjcAtLtd2nHWYBW583lzL8dN+pAsUibyD20nHzvDehYa
ZaJuPFjWf48nUeSn07r6JnnGa9LUKtWjMyYU+PlpxMDpVGCUqXeILo9TKl8DNVJ1
QwP96Y0axfypPI+MWPfUA6454Yz2mMvdOX1Pm5XE8NPRDUzOCESR0D1sCXF030AG
qD5sD1ODwLUCyX2QtSowYuV34SFb10m4kkpEHJhlFG3qxJqVK77d9e6W1yQkBaHq
Gd0D5g0cU1Bk1HWH91bDTq10ykYmXYxrI0Vv0G+9nqDPrsJ5diijZXKeeAfnSJr+
26tcePqpwjeLx4IvDWbGgh+KsixPsClAVrFv+IMEMvU1KkapRkayLahk23EVordJ
2eaMKVrqK7YuY5R21pAfPcL9jaFNmAf5XINHBCF979ZAHssxajV8rA5JaPTl20mP
67nQHUYPNquLbu3k6yRFdsjsnBH5cSfJzrZdxWfeRQmcHDpX7O9eTvpDReokv/tg
cf1h7CDbC2yU1FBK0S3qA49enXkN8Ztv0gsq5lH46Iutfomyp5BKLltr5aeGNw+6
D0zgA7A6i966vkUmYnZ06LKr1FGgjzdGIkeUxDnaBP2d+qaaKUAPwE/iMWEjtOJ8
74JdoXemTN9nFEyULuTKbYkJHvzxZbFPypko+LUGTWYhjpCJ0m0XCSb6h/s6CIkG
aLAioBB4etUh3cpqdIr8nji7nr4aFBKqvuXEAglA/RdSHDtJV+KFsvTmIq600Duo
Snh5NtVvAd2M0IOknNzn+lu5gqOK7seDfXHbmFInYBBdMmC4b57D3tKnWjlLCI5L
WeOPDTCvQ+DCgspm1Lp6rypfaAocYx1zLCb3WI14V19fJeiX9VvflGEwqNzlJdtd
6AW811xEpooZZLE9fpUzRx+qdOwPFotVrDMRN1y9v55xv5VG5TS6gpKyzTrIHVth
yL5PSEd7144za+wVsEunDL7BMDcaUlxxdqFgbrsGjUYe4ZMgYP7IWr3Z33eiMhqT
UOKneVYox5jW+eQmXIh1ovp1KbsHIFv1r4ie9UynHngn6tBiR6hkCVx+8f7nWlvs
gCi2NEcF2k4ODBc/YfoAyHfzFFdnuuuVkE0paRH4EYPQftMPyKn1u9o690pj4OXV
0z0GdleMDKelJ0UUA3lUsIjqCI3XontP8e0j6cCrCQep2OvLnVL2kcH13ZDtejC9
dEkAD+qSE0O2LnK42RI+R8pUX8P2PCdTSYQV+726RLgqffI8d6JJBwqp8HvBdIvz
5d6e2QxOFbL7sLCqD8e6qAFuw0oHOuYKJgwXiltwgOupNHoY1dLILXQx1pVhDOs3
8fQTNZ7ItK5gRA5Xm9xfxd323zd9bTbGAPWy9TneWOxdS728RxkCJ3H6ECdMFlvE
g4gahl7UfJRFQy/bqDl091pIW4wmJOKS0XY1PG4KJEmpZfwjh+O9B8JHPfNmMwNS
t9VTfJl4NZQ6fnvGicHyvYVNVaylPAtpc6zSMGbCLDGEu8AcItIRIj0gXumPOIjs
7wQsOhdukpc+FkHCSouuOwpq80NqCdOen+Vg/zYPjmTwZ107XngJhTj8GvdSvwjD
lV/a2dq2veu5C5GXnT5dxh4AQ9OF4XqUFD173EjA1g77k5TyyD+NjKqMK4j1nZg3
TiHheaAAKBBHkLIw+cXNuG6rTVcIt1eEIHobCu9RXhV8tpwEjanNXu3zg6a9Y7yp
ZYH+BZmSe6McE2kKa+yXMzoF/zk0G244oXCBtRKtONAgGYLraMks6AlrgdVQKTbO
cQ4n/AQ77LWSTmRVrFK8hOSlR2W1WUoJ+2UahOGUbERmaMWpS/P5PsOZV8C/+jXN
+U8HAQjCfXlhluIpfWJi0phI9pd7+VU9OFu2AcxjyjzImJURekDk0yaz/yUePLkw
Z1SKxmnhT0maMey1u3DdP5+Xrc0BxSRFwQYDkw4aN9XfTxKPv+LEXo1s28yfr1jv
VVzrZGQ92gRJakR+kzXYmUWm84McMlMZaEkJhHQrZ9mYjXz1BMRlJ2gb6cHvj+V1
mpZEjtcLdFuPOcBWHgOP3ZwXAAfDDjlXxdlCxhh21GZaNADbBmj9eWrGJyA4mei8
aHCK+7IVz143ZvpUd/Kx3lWizJV29dZYkzuh9jjQU3Q8NJt6HEd+Dx1/gABfsVyD
sA6jRh8mGaU334iONmopSqPKz8CXUjleQhBE4XhhR3+f99QMKs6BcQhnKQkANgZ4
DOSaIX9OK9sV9OSYxleCWRomrgQ+/n9S7xlONswOQL1Tf4ntW2N5y/cEia7J7HZL
2eQmavat+pvAIbUyX98IvOuuh+8I2Gv85q19fX7QY04r0AIjb2zuoCVms93/ssFS
jIap7tAucj1JXzMvojdskHn2GvjNMwLVdvIL51pWPg77AEM0g81SwdG2S62viaEf
onA5rzcnS4I/xbJ4SC26bsJQ6k5moTNR8r8Sgs7xEugkqHuDNKQbwyXeQwKkse7d
bPo//qTsx38suoAmgOQNsljksLImwwDDWeJHuf5nCOJV8EJvva+UvoYaXzh/3CVS
jSFZBRCGSH8tpae2G1TpAgWiHQ1uYaOXvsxl1DzE78qARYo5ppSL+fUpybfgUJRp
SdAVXnkyaZ9ffg+6M/wsbh8cWc69Gs57XtA2MHx0ks36S5pB7WVHBn3F///LPvlf
Acmgjvos56hcvMn5pUs1ts4zXHJl7FI77JhyZ1B+IbOFg+4GQttRRTLrh2O786SC
9G2EX7mJnbPIzpYGBrCV1iBOXuywRWynKJ1w2M5fgQpEJ7JDwlOv3v/x/QAr5nrt
+v009I37wUBjQWS3N2+Cv+PM8J57LiQ03QBqDQn+XSZV+hlV61Gd5glFzc9FVncC
V/jsSoEgjEOJ8LFGyc9oR5w5/41lp23XZxmoIDbwT2XNl8/q6KCfxPdyGatW16t8
Niz3/ZnLHqR17igy9JJ9Ss7DFKz4sHxW3dlH/uCNtzxlbPuPZqqstS+lEZC2Qwn3
KHRYQ2YfkjxxIA/UxYgZQYWGol3EPEgMKq1hSiATtriOHHNHUf8oT/HjaFPu/7P+
1fAUALb0bTdWfS58zlUDmppX5lekqzvtoRzeJ+qnf1TJNBUzYuU9wBRt349wBQX6
AghfPkoy9NlHeV5N8m67vA4byG2zK7mee1J0XswOkHXLvck4bYSPet4/Jam5MEvT
B1ox9S5OzFidZ6dVcgGuL+DEpH3PiC1yTxi+2YExIO4cAXE8LB3Z+tGbtG8M/lg8
t2ENnqE/ACrXyiwbpQx5WtvBVHVGNJPdTjN9+yNzUBudBtaFqdCbf/PvlaUivisx
cgmBOsa6rLrMbkntGYg3a9WMCasc21eR32UA7Gwwi58Dp4COJsJ5qB7b+4Q+O0Un
cHkH8plRoGk9ErlUr1wOAjZJmCshWKrARA/uKjHjngRU95r3vPCcE7oKf7sYuJsA
4zmtivCJzlzDveQJU29y20s8jD1fwCD2Zqx2KyOIc0gGmZLsCPTS40pmlenFwtzs
05HQsGfSTz4rSAM8yt4NpJ/8A26H5pW9fSvNCtYKv1KU7zrLKhl3cCEjD1vBJJso
CpmHK+43D7tL2ugULI3UrU2ZuLFTZ3C3UiqflDPxwGLeXwNlipyGVSc+EvDRf+ai
O1b6oSXeqpR7Kfdg8Zv9UG/UKTKxAmVi5qPAJLQG/4IzZ0ouWaN989rju1AFmL0Y
MqimE1Y+HtMBDkdha+y+QGxcblONwZRPMuFAwDzrYAi8RkfY0CjQ03aol+u38oHa
MLflLx0kJgQicezZScXEzqWd4ACJXCiaWgP6DdiRxFWSlyQzWoxDMa4sZyqQ0kA+
R5Hd3C3HhVTR/x31L3fOK8gNwMynzIVnA2OHJ2W9YMF6En6QeNcE4rI3LwBOjCzr
XqWnvf5zj/qC3iaobbw34ZRRx4VWElGDuyGRVj0f+JRocdQaJNUTgADT2p1sdVsK
6OiI6hJWeNEt/21DuI15ny+0Z9oZhY7iibvQkWKO4vce3tqSp2QyXr/s4pgpq80j
Df9EE+R4Ud4+OwvtTsvR8mzbLB52QqSiGkl/5XscDvQYepkTQXdz8A/pOSdOAEI+
dBiAqQNuLtiEDDcwQVe12sf62Wp+WIwiNWnISWVoCLMk9Cv9ofU0JaulLVZbCntf
WH/uWPAYuGaBWBI8rcLq1paHc/UJJW5VVXaabpWQ2swWLzL+YKoBemuOrsC7yyDG
SJL4pcjOPdiyHjRYADh7NEyXD5c3jJ9lh8X998KX9HAsyFJ/n15taehEdM7NvXZU
2WkEFqZ2QrBp2jOMjIyUCoJKjiYPookZtN4duJykYYq9zfxfLxBTu/+v2WvdgqvM
HlEeSxFm5JNq4dcVT4XFA68N46WfVn69h3pq/9iI1lTsPu1UpFhW41NCgL6C4E8w
l7q4zjbJlc2ScR2VAfBkWCzk69KrqcIpmMfaqew8KKLhV9/BvMEXrtXtOBMxLSo0
rO7xdF06YdU8/C77a11RQgKmuym24/pIJZl24At13OUudz8HgElolHAeJGX2aHdJ
8S0jJbXKWrni0WtpvbpvAIcTDf+h+vGMykZcZbOTY9m5D18l8v5z1cLXSnTr9Rwj
kQVKCgqDF+CoG53vj0ybDWj7qcdtJu6k3n55cyH/lSVx74EBR50pPv3UJRzBFm0a
MSHPWu1TOiX1xCZAi83NgRInR/vMUSvEgKHcFXmpwf9/c7SQq177t/y9cJh33GYT
9rsCEvr/P0yw3iJRTdlL0fx3hq2CYk+L+b/BDdILtCYYLMON2Jy1Q7ruosDJKUzH
eVhPRED0dPVwX12bsyEBm3o2jL757J+fcTIGctvPvG9W4YI/lEaZFyOyKP0A+xYr
wpVXv6jFSineLddx5vVH+uO5KZfZ4Ai3xgkAa+4pQAZZy0uRhLuSyW3bYwO3gYaC
CRStQMSCQHKwuiizfmgONth/8cAfTyEpcEn+2kssftj2LAEiHiUKkqqLy2wav0tH
QBy0LyhD/WplKLnk/Ts/9usBtbRRVdPJHWbSonQMFowskhRiWd0durJuTIRW0z9H
7BugP6zMoldDP6XVF3urtt5pn+g9T7MWV6cq0j3/U0Eu71aqDrto2yezeIh/5c8d
zIFUn3rMawyuOVctGfsbJZF5LqeoYTlj50NWgOQy362YzLhIo57yFFNgftDdH8HB
Jf2rTJ+1/WhvTV0AMgl8GjhEUt49IHX1NA4bsDLu3DXGtz83PA4beY9NhyyhECy7
oJ8A/GxSd6sBJ9ld3iJANu67CNOPiSCiVTIa6LFWqrsj9vdKLcZgB1Slag5dgZ6Y
XL1jZVhQXqPM4An6NgkBES3imHEFY0hdOyhPn7eEKqm9OJLrWRlRDo5NWLE6h8JO
lU7FSL+0cuIAQKghI9uXj816sQyhLoyRJhOl3Ddsq1tkkuQa5GnWEDDXt4E3JydH
WgBgmvj71rXs4DC/IbIaPRdCp3WTpsTP7O/j65Kq5thAkIzOOAJBALzU2EIfhMY5
EEcND+6DI1IxUILHvuOYsX36Ko8nhTXjepvLodkt8QnGdEV3BYEOKOqP5M3uGZy8
jnkHdCXzmLLdhVC39fjv8A+EnTjWI20DUeai4et97lTswU07hNrE3i+QNu0BYE5j
BEchUmbbMIVEEr87bwVv48PqXcqAr82v06X4yYr6HaqtvjC/ueJ8Wm/2YASem6Ln
1y4y46+9zjNOUIkAO1uTTe+2DIOUBSBlZwxNclJY48h+GeEsBlyMgqFt85dcMb1W
esSYDz4l3AOXBK4R9tVa42IfwXR+DLFbPDFun8Mf5oI2nVwMduLElCFV1YM/kOQ5
ZfSYUnaZJYG5RN2ORCQet89qUUeuVXPtGwbx2qqn2VhQUEiFT3Jx3OmsADhHoTTu
c9nHJUCa+fOR/LxISWwfA5NFzMyy27a62scDQoDBwMEwMvBuCWJXRyVCdl/q6xbf
LFPPCossklUfy8RNu8qRASqu9Vc3Gijxk6dfovwVc4ZzIMYRXh1yK2bLNXGHtnIg
Z5N0LuR3dIXhZV7fvWhBL9WDowjiP+y8Ajdf8Ee86ep3T+qt8Zm5/q6zcLxXa9XB
O5RO5C3VJDIgrAfGzjnQSo4Ef/LNO1EBzPrIM1UARtBtyZuyg0LoPMBN3czSbQKf
WfDQ/pu3hxA7H/6m6RzL+3YIWlbP0gQne+01uHUu11r1VwUPNl1i3P4wsM34bokX
rGSv2zZmsNACWQdxh8/CEW6ZyEnOaG4H9m9cQOrUhAmh3RGD8rXPkOQBUvyilwIB
3wAR+9aFBaV6p2dRT6WjwrkwiiGwkhru5Ni/qltAifbJ1g085mAMgp1lpj3gaRh0
r81JdBHJZSKRerYJgAWVTayy5kPiXAMOw3sPU+jAjhND3jwzuqeyJpM/mRa87vao
NNwlnCQS8xSV8gA58G0WvzBnPA4r0a3OZKfIyFlBet4LjNwDtWRD6/8tBfi9x5Xm
t4wLcyuIMNLqDd1apjw5YM0eci6TQUA+hJ4ZMqoSkUcG7orRQ5VFn65LdWk+S0ec
N494f3wO+GREgWF1JXNpXdDkQeqWQrYGlxRBgepLO0svNhT9UQLssqJBjKkf1WVW
5yKpoU9y74cFe5cF7EJRzGHrY5UtL+llaQ89JVuvCuR1NasgEnl+GGH9H4MAVs+F
1KAK9081bWgs8TVnI7MgahhMuxk6BgO+Bji9MlLbuf1wCu7B1X81K9u0yb5DjFPg
grCLTgWiLNrERB/kY+9OIhZ1bhKwNs8m7pMUMH9AC7NHEd1HMQ1v44FusxJ/A3/q
xvpvzcOQv/QxOCLUPJSHc33kdjHqLgfwpE9fMYQLX05yA1/iaytj9HXRLNJZhnQS
SQpkA34Kz4KjErhyMi31W/6AsLiV0pPfa24FAZCGYalFCxghPw1gb8LUoR2YQVv0
kMWvMWjwBmJjDDr9INV4BOvjtLS5pg3wwtQGVTJC3iljtHQDOtJyY93QfudfJOFR
M1VowCCezem1Ic44p65WxsNK6HTrnXelPFl854x00RB4j2zWMilHsA/w3Ma8desq
H7UJKpomGGg4ib3lDM//GZzBh2G64tN65/udEJv44I1FzZ4qFTP+Rcpk1WWNEfCU
OXk+cL7GLgZnQ4SjW7NiVAWF4Hir2xcaL4IQjNHD6R+KlZLGPOgq2/Bete2hY1Js
1fufmFz7sJ8OUXO4PDmMxEvCQex9f1+HomYs+rqvKPss9EQaOtY2fNZsaeCIzX0B
hMJWfamWXNkMVdShPwD0BX3voAp25vrhTUxTer748h5waa931vBg+kxG89YhTtb3
8Byj+sMfX82gl9WeT37xeMcvFcNX4bWFP1chF+STxDkBfuZd3dPQF4kPNICiceMd
jIImXPIUpDPonqaIdSXn9BkOJKcOwEYQmqbJLmVAzm/SABy6AaUdRy0nQI35a0Ld
3Kc6PeD6hTE1oixeC7cfGALHdHljMYQwJaoQCbwnRR7d7a5R4E67D5wwTCeRpnap
R89G6XJdMDJEiLb+Z3f0ZJKo279+eneAhdsTTod41xbPkx0BC1mPdPclp3amz3Wp
PVJ6F1VCmC1qfe/7NnNJbH3MyBtzZzKUSSDOxuhN1DpzcA0l0WWjnadrMY8JGpHy
E5rQ6hOQqDX8svjeQPoWq6YoEdNdfwKTECip8MYS6wl2Z9UJJdPvJ2Z/d5uvx3Cw
uV2oWnL3A+BzRQu5p+K48PakGZdpZb6oabW2Tv3+HmmvtG6jw3H+CA80mUH3XyVq
cNSJ66Ay8D3tbNtbATzjlaVHigfmB/xYCHkLfUy/gL7atR/j3d1n04DkMAyPNa0C
L6gX5w48jMi5NYa/yxaec3bWpACxe8Lo3lTHF4ItCh3E8i9ZsR/cWGhJIWWtb1tJ
cDbfRa3clVgdHEPPe0DbrhIsW3HKPshLtxMR3foBKjHYBOisL5w7TDO/vNFAmxiJ
1/LoMaOlQBTYESMRRKxjz6Bpqrif8exOsTfhO0wAcbQLsUiNVbo704IL/3i1tEPD
deFbWdgXta5p/2la+QZTjq5qGR/mUGlgdcHA7UVwQIv3vn6Q8c0/WXC22lp96ml3
8qb160biY9KC+MIbDEe53t56rabb3insdl00G0NBRm97IW2hamHmL3AkJ8rYrJS1
OxjACJ9nNeOCBHOMU3aS/o4iqfYWs533w/dlnMq3UgQjbXcQBL0Q549+3KVBRVNi
Tnir8rxtiAT6GGwJn+qTcov5Qxr4hIVDFrLPqkbH5fdNInnoM2vMOL+uQHNY1Axq
9bvcevFC2/34P/EuaHnEkqmAqUoX2dwwFmE8yvFtAa80bZ6wBOM5ALWbB3ToHxLs
LUyE9weOxEiGFpyDiW+qu6tofJKgwnTDNrw6zRu7L8ooGshRCZnRSpbOLlQS/CFw
ZbB/bjGo8TJ06ggD02whz6voCfKzYJD2xUo7eDRrly/sQwVUfMAGv960UV81Po+C
WxE3fOj+olMUjz6F3QN0y0+gQ9V8SVTkzPeiNfLegCwplaLQo5RbClgPvTbkQ4VG
VbedbK86oqiQ1DlJSaVzKiiLdo1mqbtEgQy2r40lahFasMBbD8bfPVnXpasSmb9w
hTC2F0mOq26mxor8/90sGFZHE/q/Q8E1PX2A2+GrJ03DYDem07aetBmFKbWWN9ar
dlmQQTj3x5YpHU3A7RiBYG+XW1bR6HAoeaoYlWByVjJMNbm2lGBK+NCLLBket20v
v63ReDwo5wCDcLKkIC3fevlMlFsyD1gtweTShTO3MJXGl6xc9jNkRKeTHZXr/pa4
BqBKHxsb89XjlzLtpFYn+RQST442sKZ29f/fLxkhmwGAbkxzbVvftBn9bf0VhdHO
3wLSSeMxoSK7X5Rdo0pBn2rv43L5QTPk+4IredpoONDPJa80wSyBPC9zLk+gv57B
50p7B5n+P6roC3or80o56yzXUtye0+lcxUPFwfQaIsvNRv0ufmahTT100xNrbiiS
UATO/uLNvIt7OwGr/5FC0SVm713ETJpi5eJI25tTTjEinatP2YqxzLVa38aEPS0p
oHyij+6km7hNeN4W9dvCWYdFBxm650PWCNd7OD9KKOa0WIVZyT2+sE+qZxabLl8i
EH6+YGi/SUMewDgLrFQg682Lpw0n/PD9EAUqZAYa2FvwB5uq19gw+L8g5nWs8pza
QWOwTsjufRO+HA3nBqm2vxgqHboMz+NaJnz/AhsaHMRW2XKPR54gxplDp82OGgk4
zKx7On7+a0PBFEEBflTkhbCT1S24Q0CbBEc75zlsZ7Wd+LFSQOeiZTSw19Kl2F+8
Z5RjLhi13rvWivLnXCWHGe+fuc9UWAveVAWI2qjpw0dBpzdZDPWF82xvPllu/Z44
4FPT48TPfVkixbQaH25fk3jplV4M/628IAPGwkh/RuHjkU1nDlweeQRe/ZTkKjoi
LdEBF2ts32z23NpuEMyQ5By7rzLUuFK58Y9s7Wu1cX61ljFnBoiM2eSpDS+d6zU0
JsQUCygbw3G+yQMG0NmX9RN/BrShl2bxHEJNGuWo2dUVin522Id0yIpsNdeKiMYs
F/UfKXevE8660U9rDklQTbfnNu0NpXTjtKBCqlgEAypyn+jk11p0iYnrqBbR9COS
zLzSIdC3QtMl6IJZactQIdzl6FJmITg9chOnXkkcGr1l5jMo889gv8FfPsvs60Uf
OEreudZGO0pbrlYu+M+0CMtSyLWcmjQHwVILUvKMBAC1y/LZMx2pFPDgQTFztgTB
eqkFt5DeSCeYPxE7CX7FeIVBe90krly6DXFgWpM95KvfsB54PzQnfOTXH2oOvzcI
tN4Y+2SStuL6ju2rSr4/bjCQVPPmjurSgTUt/Ldpc3p5+p9cwI9z4V/53PzmTRvM
jUEN32qznsMs+PbmYE5hOz565sNdnEsfRaLXbXAqA+axu6X7ZH1zojq1K+aorbAr
+3yoYt3fbOc2Csh4kfpSvsCGOXAfgXtxIOE3ktc/cxd6tezj7efu8EbDAmJuUpRw
r8c5hIirCkvx6WbaxHOjGj9+QpSMdFc5SvN/N1vVcAvzkUXv4TBolOfivyb/GgyP
tmezxOdBfJUVj1unl3L+dkt8aWZNr2vsoIOlW9BbgzUHrnbNPEC9EEE02BlzAy9b
mfaYA2QUB8SbmEEjn0HyNEErdgsno+bdqIXGrFX9uozQHmSNhOU2VyMhwTwq8rMF
beWgn0d0tGHYGT2QL+4MEnGauHbOuZDQZfbbwM+j/aQwgDIbfAw1Zpjk4KBFWbG1
awC4k58OAo7lsUmXt+iypdQemqyF4z6yDVfQS2vLnfScFvAfd2nL/uzUpgTaEiL6
l8fWe7GDqK6FRYFdSPD/aXH+SBjKe6zIYx5oMp1ENXvFD7TYyfLqIvFOjX0y2pst
pNhJwbvJ0TSTodbVHEe2o7u92gKtEf+Kk9qWfRbMzLmbMrfIpaut+1q3mqMoJzA6
vxLEQMFarYH9xHFbV52OSEaE7hv+PzjSW763Hziq7LyTCzLT2LgQwgQi/kEDNZTK
Z7xhlJuTWGzHX4K+roBl5+VEHjmUa1v+J+nY4lDcaWoNt1hWSmHiEbdTJ5knER+r
x/thLVI5uK/dXnfDoDQ5GiSgBCwgR9ey0AI1T6UA7yyWL6IdxUGDlsBiOmDAQ//l
q3C4onGtDoS7HDk7nQ7u5BOU7rlpNh4bkwhmt2/Ve9V70bvMcs+7YLf2N/Q6rWlp
e+Iyg9GPRHNOCWbHAkPgryBUbEnOymg7yKUGj3mW5RBzDE3kDDarUGcqfq1vlfOH
ICarGJZY59mCDBp4mgM8nucJxom/q0D8OO+I/o6brZ+qvs63KCgjCFbANWKIF1pD
PzuyxNNK3VJ7z2/9aLkx3FZZ2LYLaQxshRDWDcdLl77sbCddbbtDQm2IDWegjcbl
0z7jpsI+Qp7ZpilrF/cOJ/eKYdUvllMtsnBuPHOVl7Brubz41rFluYlaf5qJQ049
2FofX3mf6LVUdwjHMjK0eZyEw5kk9kwnPR3yFMXfsTH2GLGsL7fDIVtTCp3HKbaQ
E6MrTPdHWLb2y+KkSrSSauo2ET/HWaqO5HOvgigC2WwolCTvSe1IQ6H6WzZr53Wn
Ggn1g1eIf/bN4OpYi6Sah+/6HWYG7iXoeI0wmA335hNM1DcwR64WCBmACdsWJy3q
tpcfO8OSK70hzqFibIj8UsxqximCyfDUd8Vs1VUXdmyIg1GMRIP1nTYWDwuS3mlx
WVFo4/NfdKKUjMelACt77yomatKwDoZQYCjJFbiAzdh6+G552kflYYRVjK3zp9J0
9oE8c0OJUQUkDBDrOBXt1xDAd+aTpdepoUAa7IJOWS4ZBjIFatX1oDmfZvciCgIw
l6nQh9bpXisgM8jIWZYK7dGHUVfeo0wra+hHZeeLN9e2nav/XtjYtDELTliiinEA
sUwUBpcc0sfXfETmmFM24u7iveOUpfsbKBBXXsXLscR78tesMzYhTIRFjSgtjNan
BIXK4kZ/Jaoby8K7LyEa/eaNfjugIUXr8FZYbuu3hBIG+vsBbUk6ZvX7ak1BDTWW
EKc58yYvtCwlJSYkdXIB6Ucfojw0nu4R7lBR0ko3AUVekrQdxEEwdnhkVOIOPjSI
v20moFkYK3rLZVv2oH4lm7QB2x9hcvcpCpHRT3O1RnFUMtVI6tZfHMKQNOaOlzTC
vH+4NsnM7lCvjePs9U4vgDQl+WYNcrJm2ifZ8DEUvyMTqKX3xumpdFH7px8XFMJZ
tZS5n8VY47OrJKg0AuCBiqJif/N7htfD8P90DEfaGyIvYlEmPJMhTQeDXCmIZSDB
xfmw59CzOIXnMvgU/hRAxpqvGi6D7/qjYkB7YdW2laDV/L+MoU03NUGSemn/djkH
SFZVgxlbQMZS3Qv+i9jtqidHxbRXFws+KlZN3FujbTlSCDKsrD9oa3mi4QLGo8Ht
hhL0xqjNYyTJDGczsm/q7b2pxzuA9XVTx2956LgiWCPaC4fzV922W54dsU0zh7GI
bQtxBcxqaq0Xxcl5Ocn6hVPmHy7+Bn/vA3yBicx53eUH9Z63EAT0mF8JE08gbMmN
wNZ6DbZpigSH5+Beme8Iec1XBAUvg7fPOXW0PWBtbHHHuXk9iKgCgLwaV/hNl7Hf
D8HEphzM6PwJdCZGA3qa1mM0QlAftgM1i3Y/08XUCEKUj4H3FuMlZngVWhGdyWDz
8eWfNa5AeTdoPSXMwzRyGUlTJhk/Iz0mTDjp02RSIJs27enil3SCuF+WDLvAvKgi
WQHXIW9Uxt10WwauZEBddVSzoo7XkXvhmrAu5N2wJk89V4sL+qxk81vyEzPXS4a0
e8sVUH7zhYWUJCuuZI2qk26zCj2f0zC98tVaMCPIoVyPMxAa1UUlzcc5exKvzvmi
/BfXlg+5pRWgQ520JIFkSZfvA3tJANB0w7t5zEjdgJRUEnBCXlWF7vGplECXX4M7
BPMPxixG/aLSud0rw0Dj3E9Bb7VH5fKb+319jcryDXCgDOJBw8Dy5IuFa31kraFi
mZoXORZfo1fdIqNSFbYPMm+7/BLrUoCKRJjt+zafcgK1T02ucSa6eqQZNxST4HrG
PQ26FchWmEqgGi804CHtJCB4dlY7RYV52dV3bVpDCrGtT1mI+8+JFZsOr0nXDbjr
Ru2WLLZXqqOLOq+FA4P2ALC3YIFrHcXqLhq3fHZw5bfeY7u4RDALn2jFFb8RsN/J
jEDMc07vcNweCmDHB1s5oHPYs3hrxGqpAImwofF774Cr4mz2R0dXd2MWlLhSh2ko
yGnozzNYSlIrYj/bwgW69I1AeKOS6w5qQOCI0GXShhpVFFzckcFJSAwwgyzLUmuR
TP1ZQBXo9HmclZ/uJKRH1Qeflz8B4x6+76U18hqK2INiAegATwq21z4coxzl0QgH
Tv0yVnkmxzXL1D273whKy6JN7+o5xxjIYbtKNMKQvq22TnyXHiZhSIt3FiTh0AFg
mIhMhkTRzmQzG6zCJLxRaHSVhPMuEIkJv6/d24uHDyK3S7/ScCJEdxeyOwZtmqor
WcKjlWBqWOjvPo02GpMr2zrB3T6XBwfQjaaXDK5yl9aHUHuGStbdBWBIo4X1t+Zk
ZNJ/P27fx6C5UYiprnltwd9I6NiE8XlB44tctdq5s3qJi9Y4C9wqSzYAXuOw1U5Y
DShKpz+F7H+ukBIKcMujCHW1aG6jUohOQj76WusgOf94hAT6XhkUhJj3QQhso/ST
V0McLCd/bnqn3AKZw9fMtQ5KB//1jMkcsSM/HFKkX4GKzKheUnTO7/+S5zNUbus/
qjDxQB62CRnHw2SVLo1m1q7Q+kZ2XcvUPNkfD4SDUxuNzy6v4LPHDpE8rtP8kdal
vOXyKlo5AmqETJpsZpO3+24HmyB1DzI7zzMgyKhHyjloRhy95f7gy3AJMSLAIUiC
fBqZ55bMxBEXrqw8HvEKvnpaa4tdI9rR2xiW4IEqz5Zmy/PjGP3x2VPXGi4X8m2F
nHPyA4qtF/7k0R1OM05FFImbXqTG8wvEcX40D7+rany1J0He4wY9ts/ponTTc2NY
3amMjVejA/3C0vcPjX8zTPxEwwSFGTW28alternzARe0qfbnkBfvQqCRlcef86Co
qOzF6H0n/HqjGA7JOgayF6t/YPPme68BZ7cAzqfJ8AmDxR0sFWLQw3C2bE/xSBvH
XMPb28wT1pm5Tt1jAnuIKw/RZ2WK9M/uiXo7BSyg+G+gV2koJOw6+aSEPSI8OS6x
tGEirMrSHNBZ1iY94oaq9+cBtflR8PprWM1mJC7CKK7h1rz7YjPcxObNr5g36UFN
SeaLeX1KO82y+45tSENMz2jJVqaxqvObg+XcCTpufeWR0cF0bY2yeC16risDeLKU
KaJQp8Oezc3x8dvreV1HC4lhVeRkG0WMCYutN1ugSsPSDOuzEWMGFSsUdLVlrx+L
6lnFDtYuta5hgxOvWs8zSyhfJjRLimNx5mJcKg08jjRiqsf5mLg8wNwJGeFALvL+
+gxnlMW/hWzoahFSSA5uW+fDW3PknQmfE0zAVf8Dza+6YSJbwBVEXKy6b73zBUbH
CIpWe4SoU9JbE3LIhPsxc3qMjB6IsXM+XnyvgOYAtOVQIpBzNyG9YscFozwS/Vau
1cT36WbSCcK8cw4RJ86cnDxQ1D+PtCt8DvELkUT1DWu86TW+YkYAF0xRXirScfiu
UmCDS8vZOKQyPJbYpA3oqvModdGG+2UtP97n7MlDMndD/zAryi2oPmZRidjB6l3O
7HwN8sd7tBXsBj3oGsUoE2YaBWLJvV9TsMSUFAU3jwjM/DmmgPS7MXUwSW9R1MUn
xT9y7cOr4m9YqG5HuPJtFTSCdB4YCfWh20w+AYWF7vLNDoLSUZ85JJmDipTAmdg3
Oh19UXI6U/Ad9Q1AzPV176ECN/lUpAv1tsHd1i+M5dTyly+jRBUxlk9W2Gm9G440
FaX2ZoVLPl11pm1b1SFEm2jxklFz9cJkRj/tHlEaUssbtjskpqH/1VWNRvIpd1re
rZS68My4nSWKxYuf3OO+fpk9W9vHEeglE/6wIaOvDk95VY0qzSjxKpQe2pkg/NP6
mxQLHO82o3mLMJvBOpgpD3Hf7mkjBOHtbDq4rdO4QWBfjbFFohPpbNSw8YT9wrYJ
JEpUBJwnrqgSCESRoFk9IwPYoFRhf1A6bY/mBnm32GpA3V8qqHR8/cZaI+lOtqYN
dyHl3S8wla5YAPlyDVDnKcSx2J/enVEossyUcfSdjkKmAZAVBVEKr95aVX5jZ4Bx
NsZLslHySS41HZg8qAKibC703Y9grW5RXkau5PDk5rWDRpIggElYMx+JIA1yLN05
p1gBQRByHErzFaR43KDiE1Aqa9D5fUSFU4XsANGlofXCEkwqC9Ts19nZGoszlT9L
OeN7hfaVV77r6F8lhd+arLDOZjROgdADgHjUG1Jz80GPROnswSj6vmtL6wNa9g8/
pp0xwgXvJeGq+1se5r+QuEYFFodES9C08zVU15llSA3DVtHKOho2z0GFVvWn+16y
0wyxiTLA+1GSI0JCF00H9RvX2giR+YDYz8++Zv7y2Ax2MmmnzUWEE+US2gT2zoR1
StgxmRouwx6dAqa8wczesQQKXOkFOLP+TxIgQk3iee1BjjxMVJb1m6ic3jXqsPCh
0QeaVN8kg0KlwzaUKeYZA99qkSjxY8p1Y/cuMku4LuDkM+qauybLOAMjMdfEMKoz
kWsuUslf1VESQ6fI5jbFFcsweivHRZlIQhBdimQhmxNYtdgz9JJPzBNBJgJuWiSi
MC4LsHifEyBj0jXHcb3iAN3VmcavmsI7H6LcM09QDQl8BjzM4Lu6M9f+oFX0uKBN
I88KS0LJ/QqaRTPHBFnoryoVYUxNJ7fMVUFRRLWazcYIOcNjyd32nu83dNq7ohws
ZrB4npYg/LW7cxhPos/wXTO0g5gXG96iZzL6sAn+Hg8srxFQcNsSiI+Ga4BWaR1y
AJgNbMV2WA3pdGOxYhspgKVmvIozNTlk2QiwuO4x1eRNH3PDs4sItXxsZPLud+kG
R4oxHUhIR+PWeziOK0as610WybhoY7BtOqa4w+WnMJdIj4oxrMDolStlcnqyQkrA
e9+Zkj7LlXWI8XUc3ChsISlPxcCaPPHitr0HQ2WrPBVEoBZFsi/GHGWZ+7tHcUD5
q4egkYXJtxqLBoWNLV+zAlMkWtZh/wkMgigZ0LOusPu/Bwcx9DKXintM2PqPsOQE
o4yiIfoBcAY/KetdUtUVMJnPNeW+2D5oXZ1TSaYM7uHUX1sgZszJshsYF2Q/T4/V
YwWUw5Be/j/2Z5EI8fOOn6Ib7INN+jQXVTrB5ezkxSczXzNn046eog3NYHxWmzxs
27SHtMMeMQEQzSytSrIeUcY1/xav8lacwP2I7GKMuSB112wqBxbWm2uRS6vdnrPP
AixrekTmcI3SevRLIZsbIRf+nVv8zUDRdAFsMlIr8hCCtkI514UQl8LrzFPa75D0
HeafnwbqcAzY5n3FcJw6xiWkl64g3v1mMbDLLCxp1KqjRGKVmRCCEb21zayyAcdB
/KitnisCw27YPt8BsuYeaR/mBU4Bja2YqWK+U7wb+t4EWKVH2+eWSIS4hj5/R+B8
ewQ4xDpYlY0xej9EXMhcHFr3opd341IEC+hBYUnpv0PDVDX0dabWNCTdroVIyJpX
Ea8F5V3HhqXpjwvbx9KM9steacABmBCAFMxp25uQepzXtiGdIL6rUqmaWk9SfWxr
9u8lAKEmxnvGC8Vol/FqeIgy/Qasd5tFWH5WVn2Q66+q5n+kfDZFMQiWokS+hGEz
9FnZnnB1Ly9pEasJIFaTPVZry8H1+HKRjNd3a6HjxL+/GhKu29aTWYKJF2b9Dyfl
yYjM24Y7VX0wOXTuKkUgQxb8MYi1rfnhK7ZfT0N/B/JQcpMfMEUH0zlklZOJF0FV
GsAeZwDv634rmhwBX0fOys5sIb2o9psd7Xege8LAoX3PBHBh3s9QZNjQ2Se7g87x
vQZT4dlnttYco6TXGhcR1qZYF0Q1NFNO4TRFV921wj1qahMdneJI3Z0qJlyx/2P7
o2T/AbOu9cX3cBWwtwGg0MT6sgUc35VDNHc+a19WH59SrdMYMwSzUCdIfm6LAB2i
FVUKWzPy0+zRs4EIn5HxkTkBSeybtKMXtDguQmbSTtxYnWasnaiYky+WZyU8Tyy2
4xWTcNLTnHAYM7R8SLWds4lk3VYGAqE11qxBmKMME/GrQqovCIRbpzBu9G6ILJjS
72um8A7p2/KO+cm1IKNP2gndKX3jnBrj/+J5P9wscSmkeMRyXQUlOaqcLRUm4zwx
9WWlVLdPwWBHbnREviQDL7pvOrCSQCw2gm+W7n/p2cmyAxJHZKhAgGd4d2YSftUB
E38RpOTJ8sOa2cPUcGhXp0t52dNuxq02pOw11ZoJgMVDmY/09ZSU6/SE4/R2eJ65
kCOIq1TfoICEkPWKiS38hleLWyqqIqpSy5O5US+lE5ewANiVtvfBXAmbDsM0M1Bh
Z4JzGdcwo2IQrtrCUKBmQSnRkDGDmJnq16gna1VuTI4VoDoWT3mnrPlpby7W7ua3
lElrFiFtB/zrly6X56uhKB04YLD8qaFJbYXRJy0LZivgGA7YpGOQkx2woJV/LQG3
XWSGNsjgQKsHyMnIdQLpka0hz8n/P4Q62JABxg/7qYUNWpoTpW6jyrhaUjJijPhl
hQc3KAPGhw2Hg+5Dgo0fJKcFLsVs9SRfQkAZcKWNh5RRSOdgLVNuxVQA9FLvDFLc
Nkj20VTOzoCqNBWgI1078//16b7FdtuUZKkcH9Xs+M1sXuI/uGjG/I0G0JjUpr2/
uS131qvpcwf9W+6giz6uKpMEO6IOwc8KXR1ISoneefUK+o6jO0WvlomsuNdrgwGo
BNZ705k+0JwnYFinqcSjBdEPgc3telPo4xpGtgXgVFQzgmyCnKcgL334hyi78uDL
RR3M2e+EO5eau81N+CwPBzFS6sQUJLeIdb3sR0PsOyqRn7cJydXW0nyEWBGf+Ink
9oQoaR/3tmiJnskKqKF78zbtemKgU0Pz47Xtr2OeZ8Kyv+QRI76lHq1Jx/0f5y3f
4STWGdxS0V3l1Jgjkmg7C4fE11toiROezHKqisRSgT4EKtVdnsgiG8IykaH7ghI5
ZWsbZ6AknRgWEcx9Basgw+t5BTGXxt2AtdjnW3hJZArN5xiqwORymxBsiQgvODf0
io0fJYFs943NIf28gsycGje0zGAMLMENN67ES6moRC3kC5j01ZwKPkJaxuvw+/fY
6iLFKM6b/ZAsnEQx+PDY+ol9h2mnz6CX2HAkehMZZEa0Ykf6/bSsXNhqjvtrLyr2
QPDuhTNKUyQvyBltQFH6t0F+m5zuv7oMy4x+uadxt7U+XCG+qJhx/o49GAUs//jF
g+Xn6KiKci2H3Ex/6l2qdKVO6R6SCo8WvNRw92ahW7e62weGS5xgYpXTV7i3G8gs
WMhGYQCY49oFHwu/3731aOi/h2mbakPaEgDzOTjgil2O8mPxcNp9yYHJz5MajXt+
2/qdHJ6o61xaLUsZiICwDfFN3FdIAdv1V/RGDI1Xqa7Os9fjgkFgNiPGJDbRoOE0
osFP9J0VxzdP60AHBwzLUKZGmIAS+cQrpLgMDFhy5ewtAGkSm77Puwty1ta4x3CL
mswMq2krZXM30P3UuOpfdyDvPk6/RLFoWvSAr6Fw+oG+uFZ1NLZIhXGvgSkk2ohV
kyx3I/HV4tpLhZs8mTK3vcNiYGphCQZ6CB2odBJyfS28NgM1DAFooW0S95ZR5Uxw
+9MKq5gW720GHj6sYWa4zinIttbjjlNXlZC5UYumn9RXqYx7nTmBe8rfF8c6yrBV
s73jDQ3CGakJTqDZLMswXgZtcmdRasDS8Ya+zMxfDJ8bUUBcinNe/Mxabdy+RyeK
BRRgM6GEoTC/OczXDxIwmYSB9Q1SSQXvuidK/P27s2g8O8x47uwpOnFI0HUcG+e6
oK1ZNt1wb/7kJdth/KInnsXPn+vVzk76lCYJd9m/9lPmhLfOYojDS4pZbB1IoP/c
/rCf5lq7AUUtRzuAt5254Fdb8T715IakkPwkkPFegmnnpCSnPbE0GN4Zn+H1uO3T
TxsuFQV3GVp0vYsd29CkLjonnIG5p/7hegUAC/EaQvJNOLMM2Ck0lBWAghWLoqpr
fNUXNOTHBaU4BBML0poLGAxUsPOwfwAeYXXC/MJcT35F8Kk91+m/9JMnp+zhyREK
/zhNxe4l0VLJbmyI+k1wrjvp39NOndryKz56DVyEW7VDaJfzSZ6+7y3aEsRlbdpD
W3VDCIIf+42TjXAJo6EAvtuydw5jrIIxmrrbygOFMAsl1/AmbjUDoi7opfA/k2jJ
Ju0g51mvugGGPIJbqqXqy/n/hP/DE4otgCPn3Woap4dqo/0t0cON3k/2JlGnRj6S
dU7SMjxixtvQ1R7kFuAItJxbpw/Ow/4DhdgyoJomN9dDu7VuEWIgKmoSsMfiPXfj
vRw2Hx2uRpb2tsPHae+CL57uuIF7lRKkLIlzH5qyUncrJruV+H3QhAP8Z0xTwqgf
h5H5KMjJixn4yR4G8dX1rWKy4Xwj7SyUiDCbBv1Kh9JA428MtXUR9OACp1Gtv0CT
FMPXhzAvGTZ6OgQT/qfBi6Ut+qqqS5rWHhUoKCtwsk/HTNTHG1et81v6KJo4N4ck
ONTfRsvgsd/bPcGDEB0mp0L8+KjvUCL1fYUdyVKEwRQnSz1UB0e9Zz4Mx2hojyIy
lSG1FfO4qNFH7KlKd8kFQpkpv1S9d11X7zY/LEjxfr+fYJXYNV8t1s7tWwPVcgx4
bHYrnCSB3zkXQEiXd3fJHn0wZW023cOMmEUgaRAK/dT8ajoBgAtFYv/P4dRRoC9s
DhuW9Y6nwaXVL9keNKpiVrL63QQyk25Vx0ddCgZG2B9L9Ox+Y391jOMRRuFPMeUf
odM7Fg10kYGMFlmbDJlNWKKIL9SyJUJ9eV3XPStGbdiTGBk/YNWoe7lM0ZG4wKEI
GnTv9LzrHKuBeF3lM+c9DetFUKleHDwr9GQXeq6vkATEL/1y4KTpY8+Aspx2a2Wt
AMXrX/bTGqDvJUWGzVmWzYANnNH0KBOETNkkBed9pAtqUHiXtN2ievS1MYUVdvDZ
5KTZN7/CDW1rahxvyEuLpyoUy7fNRWsEBmhiFQRZ5VIIwUQb8gYGs8SQ5CTK8x73
Gt3rQoS5C6bF1iF+UCCiNlzxMGxLtgvIsyO7UeEnEYoTpqylnAJo3VedEqtn/BnE
6I1nkrLUt23h/aA6fymKzBKXqcN7tusF7wt/YQyJeNOVL1s+xw/QdFXCAUxQpSrR
w1b4jcZkhgSTbevZ0LzyvcXdElXvzozvYUQlCjlGbcXCCdcB36eK49Cx11D/FUl4
eqd51ENr2aZwCK4AUrsv/2m72olTwVzXqotZ4mFXJAbY/pbVAhFzcIaPein9530N
kZdtHcVFIdneIn8zvXbCDVojFci+TAovbhFpVPMgT8CihMuLPr64ULI1r+ZqnUuY
7f4yec1uHVssOuYLYCewZzzCoQjR0HzQ6lqT5CRZ/cct4K8v9KQWqPPfz18roFCX
LdSuPYrAVwT1s5K9zfakDPTF2XcTMktYmHlIeDAUiK4e5dAGYWNvTvdQ87gd1r/D
udQ8pKRrkMXLWoOGST9V/qHO5hKHe7z1Coj7FOqpu4P8IotP55hRBZ8/75em1Wv3
afn9xKhrSy0VbOCtZzMkO82ghGzSWmkQgc/N/Y3hcmu9CpJCsGNcuQeD05ccCmAT
3j97nxPFE8XxsDPxiIS5smjIR7+0T7SGnivsMO+2lf1xs1F053Lw5YJu3dPRyGZg
EPdyWCYffD9UwwULk9pvJ8mGDvavmsOm6aWH+x342JT9mWQm6wiUkAIk45Fpt+GU
NPJu+vKzBqT3LPNAH9bjttNBQegnx14ChmRl/itvMwGJqIIFcQzIcExisUfzVVix
5dyMomTWwXzuMQ7emlYZI8tADzInMs7h4jAY2yZpWczrRljoLQ82F2kkSeODoSq9
z5U/havoYZPwlnOCqwR3nLf3L+yQTIemMfpSP2mmz9Y/YExPgfVqpWHEpBOh0KJ3
zMma8LYWQ7YSRQiE+fG7zzIINnZlM+y4t335r1xs5lNCqwkrP342qvIneoLKgJZo
M22pTA1KZqemiN8utF84yDekhwzIn5+Od8U/WnIH0jjSryy6gqMjQ1kXX2Mf1I+b
UAHq4blZ07bIGJseBebbiQ8XtqXkIuVl9SZDmI6mAMrNtdzOm0gbcb6cqq7JMMfL
g8N7+jRRUI7unv5QMVUcDwDd8+a7ZyGDGUP6aoYK1Xx2s/bdGBJjuc9Z8XEEP4BA
QpwAr8FwBXmE4Q3gZ4Z/H75yDyuVht6fxMzNyltSeViF0FJ7sF6UDwAutBQ24+nY
z0BXgIqlBaPxzD9vlMqzwbJNewGWT/Y3UY4wDzbUQZdTm7eVXAW/rgJ2Oa3gePtN
dgg2iT6fkhpRqbXMecwnmknpUnhfVxh8XwkkQD3mpBPuyGRmjsRx1tffLrwWS7bD
HcA+FD0WHUZ28EoZ4s4yFjls6Gqve7QevasSnF0Lnhcit9WcaQ8YjxOtBaqHMRyU
F4W+u/pZWH0or2mWmv00wQE0pkKbBQyDIcsm+wYWvLnunp1SzdmaKDAeIvse5jSC
yWOs/Sy37c181mVxxsAEhWbZb7a4EbsxY/mNfTIiA0NRnhv9SZahs+XiCADhTe/n
/z7P1XeZWBchPSjsIVbediCoEVirqgG/4LttckmRQWjN3tdDsYe+3G+ghXoUMMWi
bhxvbaX0M28yaaLRTk2ijS5fpDgqdpUhaMFViDBob9rfIPkOHeliK3A18mDSxDfb
7wV7RWX35Z2Tsp4bsXh8NOiOzAt18jhEeZWDhiu11q8PMKWk3mdT1ykdTZ8fDoJK
SqIKOiFPTnTRws2GatIcTuZQ9MiAb8ckMskSzryvtcpR6bD/vhDCvm5haehZ83Si
hFRUh4MYJCSuZkTBdtn+MD7pOFpgqVuFDEh7Cg8Wa2nqdJOpQx+Wj6XSmnKdxdGH
gHvDYOuK9D7d0Fb2Wtp2eExsRgSebhFO8/3YAdTpdAt6A+2I2pkRTVbjB3Bio11F
snEvRG0O2i7spJQVwW7XHZOiLhX6/3qWfIpfl/lllyf9s12oYiNqKj/h4DXAizaM
VYeXdmJ8z9bGiN9ScTKcx+kCgpRY/xya3sakjZbZ1slpI7ympt+lTxXBLQXsrMf+
s5filV6pxGk3qR8r8yalBakwvc6IH9LzFLE7S6zE++8U0KMP/NdzAtUPTHazpu79
cFE1J4PbKZXcWwGY+m/303RzZ+afGXOpzoLQoo8JTfZIdWwHnaJeP/6QMhxo77Al
R3C/j/mUb0pCv4dRZPYgwg8xW3A7cv1HtHP4jF7dABWkatSxIFBMy9ZCzAq6x4pW
odVGN/9Sh/SQ7X4qBcZS/X369gd4juskmhmnoVS+mQaVy9ZcEhxlPymNDYjTOvr3
Bx0Y0Tt5nIZmI+91fyBRhu+fOTD3HZGWT1DE6imREEzDs2JxqBS8PE2aEa5igI8S
kW2XWfb3Jy7GAOJ646GkF95Pq+teRZUwc4FFmT8VNi9fvItAMj1KWYojVcigTX//
t9E5xjFf0cYHfN7QL+bIRCCZCShhKPf36vsUWnWORO4OlGjlPqTqCC3WR6zhxnH0
bh9N5mp1NinHF1/8V5v3xzGbC58fyqRrWWbi+cNMlaoKbPZx0+qsdInmioED9a+C
9K8JCg+ZJ0PgtBTRHWhSzHaQ8wx4bq6TEnfb+zqcKPdn81uDn8oCJMxCPGc97Wi8
OrSQXKFCsVZsIALOOOYm4DrJQTyL9H6prGHK1E6KyySBaD89cVlcc/fDUOnHjCft
mMXsf6RrZKs/ZGFEsV/B46eOjWSC3r8sEDqVJ1VdKdvIwRsHmtp5HfyK3CmQTD8m
J7ZXfk/eK8L/LO7MtFwLN2w3k4wJLn+iWkyCwofVNi6BTMjlVHcttsV83MsKu5hd
peENnnlF4z4HHKI7ajNB42ds0QLh5JCeMG+VRHvRcsOlieZkNtrxbzj+74Y2wuF7
8+IuwCKJTTBfsmL7EjCWn4KJ8c2JItT1XtNlSSlvmb7QXY7SQ3V8OScWZHGkD7ZB
y1+UEL9U5vqiVGV74/3rlRsneAkcuoNnkxPUvJenPrn1MQMhAUbKidSTHwTwpY89
EbeeApg2Qkow28lyDA8LCH5XE/sPXao2OpSqMLLXrdwjtV2q5QVh3UXNlgGpVJpV
plNezASwPI4oSH8lGTjTtIVcMSsYyzhXrDaJN4LDKr3Ej80A+ce8tEUzI2TJTzVR
fao82UPecpGpWS1m2CDsPu5D9ehfHynLi5Toh6eG2jS6v2UCe0eK4F8WN03FOSdl
0EhrqmK9c5CskY9aZLrOaTdGrnaNoMe7C45TgEri7G9hHuAlr7kCyZegDgFfaPdV
XchuPb4WtOBzQ1Mh8HuzXzvFP8ho+e3ZGuVTMULPgI+R5MPTgUoaUqCoAIGn+qHo
aUTSRru4LXVrIVmsuVZuv1qPUzz7/zk4ATFHtfHGjZxJvyR0UeU2tkGK8TWMUUTE
50Adih9d3OqmEFoIVEpY14y7iSEPjj/QgVV4s7NmWWYc9VpQIWFJoblYJp13Pmpr
BR+fGtyd+4EhhYLJW5drMACXFR7eqZ3RqW+LvRELdKcHY5TulM8KOx5QgDTlfZ+Z
4LuvjJfR1NqLVOYQBm8OujWKg72UzBu0i1wykeNu+BfZ4alnF0721dzFRn6DXgZ7
DVl0FfjgHa2lcnQQR+ARUpfsxSVHdJ+/9Ml0hbprTc7h4M1hpM9iFuwDY3xhiAAC
e0mnktK13zogeTLBesZLYAsvPEr54mDPJfW7jbERwPkouuRUsbDzyMrZTxVVEm5j
beN5fn7haf27RQM5A/72Hw4KIWw0ekqGDv4qwEq1pji0D6alF2MG781qABF8J7Na
BSygsztYfEey/q82wY9MuXe8AdKcJhmUviumyB1GKlk36UvV0zFWtB10zDCDTGkZ
qyP+oJtJvFqr1wo6vWoFvS41Jv13VYdb4X/upCxfVhcfIFPhInoOT0CAfn/qBihn
eEb7mWyNkW0nqHWCbl3IDpVJsSSaTmYaua0t5QFaFRZuRxdxQ2R/etvw0y47C1tD
wFVxQl2h9eGiQnr8VA1v/WixqJbC/M3gNmF8Vh3h3lVrgWdQ+8WJt934389HORT6
4hkrz1WOc5MSrN5MtXCp3JCC8pR+bGW7VQAtn7EUNjyC1Al04EletqO9vIhScng8
90sIjSK0I9dHBbIRv26tJb4/Ry4npTzEXz5dopCPKO8D7Bm/dYcRyGF0Obdyrv+0
pfRQEbm2eRdPKC1fdUBPPX84XEN1HLx69I/+nLlpWsYIGqsqzCL95JAvYxT992hf
jsZHr6UNHJbBSH5fywsJylLz9jNjxMMloRy4b8aXgt6u1Mda6kihWLAqUXxFHzJ9
Pmb8wzzht9Y2XbTYCuPZiRVCEIne2JZ10V5Dkv0go5ViX0zCF/2e+prdJPGMAtKV
HcTXWaIkT6u4SLeZzNmZ9oQyrTCezuilMjf9Ans8ZbzKUM1RumrIdu9Rp/vfIfDD
+3u35Be4o8Hjb+MNukN3U/aO+WhWmzVxerU+FxPPjiEKnXycbibYzpGBBdd89MkN
rq7ibyCWBLLxUBPtFegsCLasDSCdFn4wTzUJO9zKPSmCyzclevwNx404nr3CDPO/
v27vqIzLe45cypaUkZjsXxcOVq07N1COSSovz0EzstSoNnAZn1y1RPzgKkfuakzC
ss0KZDxpCBTHtPKYj4+1hcDXu7B4nIddJF4KORyjh1ayFA737iQCsIMhkG1ZKWfL
F0vWCD8JiqR8CX21VZY0iscf4/DJowjBFfWiKsEH+KWqs4O9sFsSzcQRiFVFDuPY
A57GwoBNatpCqcDRGidbWDV2yrX7m289tBum+9OaGbTZrqzVQ+hhDCalbf7tOZ8s
+26YL5+PV5QrjDyBXli9UiWgTuwbeQeq+Lk046TIGfgmb6CSuVheuUbc4pxaLdU0
cjNzzkcDe5Ev8fYYDbw//FkMqOaoxUv+ma7TlkKrL9z7Co3686WliGw5sK5fM1kj
zfRcApKUr5T/tnlSQJgdE7BHEjQLaZjVgfuYnBNToThPWgCATBjkbfRtjwaCDxcf
YqVWVNInlMA644XV8druC+F9igGhoZWDJ8ZgXSMctY/9k5l3/pz/aofTVwEda46U
0T8b/yRpjkoidRpkPt19WgBKS6HRnRPVJJnMpYUisNqDYNSO2TClV/DbIlsyYExC
H7P/wijNpvmKZHOWNWYlhnT5+ZbSXiwuD5/w2qXk7iX3M/OuRgpm+k+kTmJprBxy
Lj442S9WpYXMy6rw6FTOFFirrM3Yhd0tgReX+cX35oBQPJnboXWkxSeosOWHSupp
4PQ4NFrnAeQyP6+UD+3A7z7a65ssN/J9Xp+l5SVxKjt0p/DlOZ8y/+dp6Av/ELh6
8lVB0m6bKOoBk1uBEPrIWE7J9R4oN8VGO7T6Dda22JB0Tte2P7vKOh9mLESM8ii7
uw91wTTc4/6xpBlW4gaeHgHwKT01oZzxwzFdOltkusQ88GFIGl/p+pFLUqS7wNWo
9EuUR75fN/JVo4AV7eXoXaixYvVeCL2RbggpQLeDAU1U945EwWUT97o9xHhT0fkk
fjD3DBLF7igxBcmQGyHmmJj+IKK0yh3fnA/XBzs14w57iFKC2vlUEUFgwyYFHGya
7nXBog1IcXNKo2fbDFHHhO/fuiCivjUDNfBiW0Kd7LxDqg/CYZSauPtDyu162IJP
BIMDy4LAdnpFSw3dmh4J/pDQs76+70S0ZbuGR4OFkqsVs6+tY0jCF8Z7vhPeJF/p
qVD5araEcSVtT2sVziadPQ4NCO6iBOdFDUjEaA68cSwaZwMj9lUDpm4DqQ1QB8km
wvLBpjekqU6Pie753RmUJEyO6wRIcUCAeBk3OrefihHGre7rJUzxFhGkzLGzjWRK
HA/mP9tzboychJ8ts59reqfX6hkolSi4YXnZuOC5XuK0qUkWI7K8CHOljuMQkp2n
XMXLt01k+hXlPMyXdyotB/KGRaxZI0nndicDYsWm7A9h+ua+AK1VfHPmh+LwA6Hr
xU3MMEx//kYwF8yjr83uaxp09zo7WgIdU5U5t2eCbgmACGNj+dvUDIYs2R84S7n2
rLEbNkfd8nQdwtVC+42RB91X/n+KcI1vnbThRnQX3eBOTF6SB4qtPbmZ5kDi1LEa
xnZ9r9pCkMxfS3AKiG+kbZ9/DcDyIQUEmZS4Q72ghjzs5gJNk5lTZRus44EB4Ft+
hx0OUfLoE8nVmZUy6g/VtXlg2YkJn7Z+g1WE9GiqYEXOtlB56qQGsfj3q8fYzzX5
8Qg/dh5Z2MWyLPiRShH6kRq7m6LRNzpa4zLBdVy3rhplwUFq/Y31ez8VFx0/JT2f
KsINwHS6tTHw+B7kTJMfP/WUoQnIBXUKoj9qqTzPg7Z0G9vQjeseRvGl9eD4e7x3
qCJEQEDaHFaPM+KN6m1AFUqKtcT3+niKbqiGTR0cMkJkgg+YPKOxbLxnDtrC9tg4
gbA43iXb1C+ZzdItWiAspfaOyyyunrOzg9sV2YHDJH+3dSjRPd5rBs8YMOcJozWE
YGPzVzC4yUQdzXACjztWGozClEjeN83WPMYNWPrVP+GMk3xkLGTq6ebSVYjJfFc9
qyY6GOjzNK4gzuLAO85Mep7fL+fL/6jWJSCddRqlu97rui473YSbTXgUTVln8c0B
lnL1wRt44eVHqflzLE/5Rg5WOB468wlHMpQjeMoauKWruKpI0TANpMfZ3KK/gZeK
`pragma protect end_protected
