// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EAz17TAMFH2Lc3ZD8PHZQVIV/UWxlFy0NrEgvWAqSzyeUl6W4ohAJldGdNyBo7sr
5JQ3LgJzI1Wft/Jkn3lchRX61G/WAFl4SxJftaK4Y/PzgjrDgGQsvJ1SI6v9LcF0
41NGrCwiaX/p73v/4cdlWuM/EJfWKwpdQnN87lJn+As=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 23072)
LW77bYcHfVuCtEf693kgSTyM5L8Xehnq3lN3VDzSRYrrIDh2g6nJkEtd+OOI0o3B
ax6nc3yURdKgCqBhdAWU3aYYSs1cwpgqdoXSucDX6ymwpOu55/JBxZxISUsHl8u+
axCt5cJZYgbnfpjcLF7CvqG9Wg+YkTFnS3E5033qiz26EDhoizvliJbEeSPFsjDW
PacWrNH2XXKGykuq3sGEKy5lDzNQpDvzcS42FjXI8RvNa4HblsI92nxCT+l6G8Ip
ShAXHYWWnFus8amXuIg+voeqIOtORrSpL8g609c6TIxV1vUaxASRgTAxLv867uez
Z01br0B1A3gJ7PYPmtWkw5iYfbtsxBviraqu6bg0Ap6vicwKzpZXFsEvIWlkWqYp
LV797e/S1wu3JjgnJltotlNpTvUlWhfrezWZhszEw1kUXIgyXKpcgg+CGQZLeTCA
lX+pKKir3/U8csj2d7i+0ttvi1LI54bUqK9xQx53toU2aVP8d6gzFDX4cQoi+WDK
xSAibpvyAzFJspRcejIP8vAKO1yNf1zh9L5eOVPmZBMleZqkZ0EUIY8SEbBXC6p8
9glqY0gTTstmZGWtsFMlje4knshtztunr0SZtFoRToenndug3cPwW9i/fvGteJIV
OhZ4JXTHo+uIFR6yQiicwalKoaXHPVcR4VGFnauE0OMRhmmjk12uAp1m/ya2hIjD
zNxyBTTmLDvTmYZDsRhAd45ZsJ8sfF7JK3tsC3CbYuWM/27aU8bTfL5DNhyxQz0G
Utc4HsFjtc5V0RIdJFY2Euo2RJGp464v3nyH+VXVOUxjKRJEHZftru62+NGsTOg5
Z1JabrvbbzN2BF4Ulj9hF3lUTLPuCLGAT6IENuHsTybKu1ECbCNKE1PhEjV5vYfT
H71YBl/Li4K8vrNdlrx6V73mGVdfpi3vJucZ7EjsbI92mcSocVhvaTNomIvnQHSj
ymMaB3bxmD6jzDVf7zhefe4v3ZezlDof+x4CwDJsaVLaqYxFYhYTux9s4dnco4gi
/+CnQRCenQuV4HV9GY/RZV4Hw6bipTguqvRbZ7/S9+dl5YiQxeZtOo9i9bQhQgJh
Ik4Nsl47AUqMV9hgkMu+9e2Yz2hA9pJMqDjIvM+M2EZZ3IJz62y1+J86xGgNFTG6
mMJuhWN211LylH3KC6DtjXHhcSFazWns/BbuCgo0JKDweAhrZiee9snv3y2F0zlv
0NrJ6Z2IiKk7fHE49Xx2/mT8lSA11BKhD8YeP9WGSrbyY93htbI919NkrDu7jgR4
b11yLWvazgfJwLQte8jWb/NnbV0Xlu4h0DzVh5yB2t1RuWJS9A+IozFUYQtcu4Wv
1gl95Ab9w6ITSxqHOHNN1RqV9JDvM+EXPeWlL7Ol/BfPJWfJlOZTaV1mjUF8Hz6U
jNy3/fhLIGXsrKNXtOSOBzFPy5uhirMOZqcJljini/cclYd1vCJLhuVN1xk35Idg
rn0ZQ0g+RMZ3Ii6WqNhOZGNJ/pG9a8vy1ASMSnhTX4cfLFEX/dMkOXGtFfCUgQ+/
TdvNj30txterqfhsVPgAtLZUUt9fAtrg2CUTr51/4IHyXg0iQaaztO29eYWczh8D
Z4zFGt+qrXxu77b2sRndc6WQqU+bNft0Tq7T87X1HVK8v/+f8m4gUdo1jnHgHHZK
42hX4K6vVQ5oOZ+cnlztOF/qWLQ3eR5tL39SKXVXw22VJKW4wPPAQTiNIoxqEJBJ
Q4/ATfxrfn9vhYynaDsYMs6IGGGbrpv8IwKjwyxezpgJjH/4UCMCf3c0yr0nLfWj
NRg6cuJfbknuLC4NooEB7gmcHI27AGid71adZa+ZOeoJaiUFOU2ccu0y8zTTzULW
Oj5Nxsj1+r36OqB8lP/OJjy9dh/5SOief4HrcFWwDhlSeLSqrw7Fu1AR7cygRhkM
Df8DNUDo4n+zJWYgwvs6XnE+YW7lOgrKtNpVY0dh9mb68pp9F+rhLOZKzq44rDVm
Rw+xlpjCDI3nk84otSXmqrGWKoKD/pG0uBkF+qAwpRc4o4pMbAK/wtnX+aQZXK1c
1lTHu6+zsypnVX5p5BaEfhxV+CvcF+Zd6c5D/YRUII6s87BL015CHeR7TDAZZhpL
LeNHmUWybFjKQwW/dLO8W8GJhdlVmU0WfOpBChY9NAQieggtJnDOHCy6C/XbosUx
gb80MwsChw8MmtUJ75ljLj2CA9sM7EOEUhfu1e1GVHs6MQWek7Ivl6CTn0iScqUd
/agHfl7fORlOW1SnejYaJuLf/zRehqjIUVLnwBn9ymgE8tIB9IHNi6Biao80xaYF
mBW6yfqPQ0P6rz+QIX/DTaWVkr/t3kM4u88jbHXImbkeq2dk/2ZT5cwWyi0Q2oPJ
fU6f7rOsKQ7RvvGKMZY9B++mnwZ9YXgF36yNWIAdFFt2+5Z17K7u43pyko3M88SF
6zI4JTDv4Wlv9bmZJ/cqYp3AOLvCm7OW4J9Ft0gOKRlqj/uNfGA+iZ2q47WuCg0U
vtmUSJDqAPPEeEqdppefWJ7b2yhIqf0WnAK5iTUVLMD3ZsjC52uJzpPjFJGaHMhn
Fx5w9csMHBsJsC+AtazofjnFkB+ON8U4FlRVdoedcT4WIG0goYZhrYDfQA1hJjwp
tWY5evV7sBe0SOE2xUNmDWyWPx0NzWoAU43fkWJ4Maw/lepEDoVlD1rZYIHBbwXm
KDKMQk9WDnMEScgSK+W64v2GKz9eALdRmu7fnV5JDjygmH48uywGG5+20ibOTLZU
a+2Oz9OaQujmXa9PpC2n1njI5GLkWkp3GMElu77iGZ5jrX+ulocoFtT4NRTKo6hB
OUNamzm5ecOSmH8iRsr4GbmKNFx2ovN79pHRbpcaYaT9bRA2XxfFqURPFpFrW9nG
Qp1xhqpGjzsR/cCP7b2G6OwHpD5yNgDC/JBkaJ2dP/nU2PjFEX6IVQVWvESGR1LH
dFtVMDL+IL9mOP48mFK2e5Zjhv7LSaj3iymnb9/4YIltj70n7Vqa1hN2f+CXiCyS
2dczDhTnS8gXmyr5khGkt9a0cdrBstxqwzIYfM6vvi5vD0167V/YpDYAmMQ1Vn4u
2K5QWRwA9hEOjXPq4BC2K4x2fsvBdhl0Nl80JJX+m0tE9t+xgFs4HsLP3VnXU8st
jto8erfku16JrylsH1fRV+LV3i0AoRkPHnf0TjI28Fkt0FuhdXuxvMScaxvwNyhw
2SrmNHoNeVaoLYkyk2WtSXpVfy9DctZhOH6I4lN9UGd8oyxNOq0ZTk/sqquXtjkZ
303sZ/j3xOP8SMt0P2r5UWstXbHfR4UJk+HF8u9PcmaQS0a65584I6Bp2YqRybi6
yYxC06FSysYaylDdcxU4KOgThUqOzq1Hw9pkbwPWipwwl5HVzpH8WGl4HBNWBV61
2cmZjBHObfm7RC6iQQ9hLcpD6jz/uoXNYjWoBj/1dSxzBpiBR3DMngqHg86t9iNc
+HohrW7u3njd2ZymsVFKEZ0r9U2ShJPg7r4s9Tdqbg27/kj04cp63I48MChL0Grd
aI87SER5zjWdfXO1SM77TqMbBTQQ3ke+A0m1YYwMvH+r79JHYLBmUh2URQC+AIMB
mcuO8umH4WN1LOwkgZPEU0SkfR5AKbFXnlqO/dJcC1fEgh/KiZUvpz2qHX7zJVI+
rDDadKHzbZ3Lutd1VsNUqA74NglqITzNNlBGBmyxMLjbajeJl/p3wTdGHxFAobem
2xg11xi0eQjm2EQkSAid6AnUQhiAfkMjpK2pjth8DIM69fn1m44RnoVSRPJOEAcF
PJ7UutaTdPFHV1g6YkmBc9aTVlsUEcQf2bDjJZpkqqFcu4dQGfQuwtjPDzOQwP+Z
JCoBG1WQfOPwJSOIktI77fb72p9zaylxMbBTVGBVAAYyY5tzN1I6KWdVBFb8fmgq
MV2j5a6asWXLJaDZB8MvUbD2jL6xBaMyzNkUUVv/w+5FXgcmDFuGrxoMqh2Pp8Ik
P4a+ttt+b89mqHXKsc5+ya4GDq31bYMQjadwTRQvtuJZGvBkoYXxpGryD2GeYqT5
GBic9j5wm8UQvtHPq0ucbWwsdbjf852CMrO/L3PiyiCeA4mrQtAtc23kBLEG1GmM
dqJeBU9FkJ8zXMKTZYKl2sc6pa6Hq9HBPGxFoch8hAYUAZoqbre3avO86od/0XzZ
hHueTA2xneLMpRLgII3EgDt4YQIliTAIPevmnQuhoQpuGFcEWqdXqwa3atIG9eYU
lJUSdrYCjH1mLZ8XHmiA0lDl6oV4XnDQfYlrh2WsmwC3OIFmLdBJ0l0wyx2Hg8Ye
HxIU+w2bGQI7WBymWyDSLMY8UJmOsHMKv1EQWkCootx7cmk4bmcet5QyQpYe7FPC
/n0uIL+MNjrBcJr7Ds/gzMOM9RxCl9h8P9MC6Fg27oBkCbdgqcIRBHvLSAu/oJje
V/Nrj5TONbJSuIHzrNseDTxYABCTVLY54ruaimZitrXXDDxapzUVfKr5LoKkWqB7
PxJxTdefp8YZZDuqssdmML1jMDFq0xfZdTXghNupQG63123m/rgkDReBo9SQ1n2A
bksr4N0xe4MA+pNsY93ymjYzVJU/wJBV7s/RYai+zVTka2ArWV1K4JlPwZKAbnDf
yETV1kLDTl1Vp3f7QIYVA/Pf72Xt86P5rLDgd+re4b7+lsdqrSe5aGNkCNYx6ZFD
caWXzPPtTbMWPoiJOD+8OUVvPWIrArK5s3oJpNwwC4jsboLt3tmscYrI1S7dhszQ
1LREt+WMAqpAH2UvCA/AilPqnB8sR2LVgy11n2Hi1RflpCIMA/kTfbg7gkcD5y+N
lsEb+IYnEpt2bd+6vRstM58XTOBKEDbzUUJu0ZeF5sqnqE64ci5W1s3U8F22JQZh
HyzzShy6InWgsp3sHjl1r8GDg0eGl7Tfkhh8SugGAT6xc15/6CggAgPsztWOcDcF
sdAOnMkFYjh86LnURLynoIOaiHL6sXyvYa5YRcRoHZ6VXybh4WAd/YR6l8GTrP/Z
osbZhlsRwsvnuDvYqf2JQyL+1c2V6r8zHYsZBp1s4bse1s5rtOMU6SZbJs0rMMve
7Uytobyn7iWOPTTIvczjX4/raO+23zKM0lDVaHPnHYuHDebqswuI1EPYE1Bi3D6q
FA3GiNwYDH0VEQaX3mEejiseXqu4C19KBj7jD+nOSwy1/ue8EKfPF1/md9dU3cOk
+2pgpafTy/1IBDUORZl5ChfFH6jAEAr8zbOSsbHEO5+w+7KdF3Uqx9pOdZcqjeOX
8sjnc/wX9W0C+qay/VGEKu71GDTMrIuyZh3K1/2trC8YbNRHSPa9dAzuV/qjI+nR
zTgaZJ3eZnbvAqDPHTXvE9117Jx/DX5qlognQy7twDv1l16vBST7UjXfgeuFFWRh
lBHYUmKaC+l3Xkmwz8wi+2EkJ2X+s/pfspq2Hpt0GWRYbD/sNJGkD76XyvjYqeDS
Wf9tqzS5LDy1JG1FefkSVEoProNHREPTrfNLrqnZ5obmaDhRBJv35gyeH4UJfUgA
7dcc7yoK4P2D7PkTG8R2AgfFaGodbEAFLiqqquwrp/rEiUYrrFTD0e5SSIiJgBtH
m0BDvajCyh4BJ5buBKXCQE0Y6x+huLOfMGuGZi1AFxBr9yDt3M9MAhqD6du087Jr
gupy/4oDVSVcGmyZN7qp6CsjkjOaMVjpuzdtKb+aIaYgONpU0bIa7ZAiIDATYhYX
dL02ox3pA5JfIhfdZIedOsC3jdvpPTr5FIEvilSv9Ezn5ngNifduknS6sEV2Ctol
UrLg4Tm1501K4+W5x6iaebHrVbh4SCnxHxpkYfVx8/nXetcRIDEyjBJ8bdAWhU8g
fo1qxiU4bL8HpzsANNd3DN9NACj9qaCj9kJc6XhStdGDFd4IjBHAo9qoXJHAGJMw
/HAmiuuDAl8TezkdPwd4mURaKaOrIjc+tAHpLaZjk+TFxzt/8NlihJrGgq8yTpks
BcTWA1Wys3Dp04A3OUElaILpLdGYMRQP05cW1VxXn4aaUedw9+DTL6jYoPL1K9mB
NYg7Yl7x5HcZrhH22vlxGEsXTDiiYqug5LPsxgVkBweOdxFQu9dla/UAligKMJ/I
isLAcHasnjkpHNw6/+D60DrBzsu3Oc/Hd54Zpibhc7W/c0gnuyodvHI3KLKXXIJi
hjSmiehOItA8gU/ZACJhY6bIp/bXbvQRWqRwOU3Dar3MDnbQ1j0A5l55vNkO0RZD
mw6MkBkCf+1OwPY83WCU3pqtNzRIo5Syiw7eSZJLQV1l0W/V8zZxSiT4qMg1lZ5r
gGJcv+SIbwFEaj/zhc0sUiWCT+rad8khMhr8fn83Bt/LSByeB0NNLbeFRR+E5ywc
gK3zatu1xhYH2iF5lkdD0Qic8Hrz0flQFeZW0ALgcNimct6v4i8Byrt1TbanvBBr
JiI/3e72bOAU+qKTzjhA0Ber+mceSktsHLqAl11wK3kPcaBM0mrbdGckp0FwJ6pE
ZmQx5e6DVUKjxDtBNISE496GKNa8rfl+O+KzBlPzCjTOy63PX1GyKJjGB7gp4pCE
rjcU/kj3XE5UhaXGvQBtOjBfd0xnfVMAXZ/wWpl7qjobgW30w4kp+bV6NCd0OpOU
8I1gNSqAeARcuuWVF02vuzrEKceeU43MNe5D49tofn4pDQkgKwtVCByB3U4m502a
UGaGNVbbDCgWnEmP45MddQlfBd7I+WlIiE0IBGU4Cxnum5qOD1lOYinNQUhnRLGj
uQ6JdONOkIShy9PWffaz1/lV5UCh6LMBRM73Qarjq54yJ2SvyQZXm11lneSo5oeN
yJlBHufOYhXPTRjOanCYkV5cIeDZLpI4CBTrlQhHa6tqaDXm6zC2PVXIHxXfNKFc
VRy407boj2cxQ1HzGq/2zHqLkIGwq7R5EAziIQrmKbBiiwU1YnrpJUN9NDMQcIex
iEDioz8RaaTXjQkoCqBJ4wFZqXupiNaooZfK3VAeUK8/oUXTFchMhXwNAF9jyGv3
6g4hxvlPC27EFZ6JLnbzm+uiGmNG4X58QYQ1tWrJn0K0DJlAzxuDAvKZ2iZhIXpF
jO29rmAa3BIpp+sQxvRXUAfuXRpY0Ycsi1FlHCTRMngKAf4jNiE2b65o9vTYa+h/
S3I8DcIUm8YVkPusK8Gl4uM5ZBTTTJAKFv7S8iz3131ki7cA+MdBZ6+h3bEUHCkG
wfnOjB8hM8dRDdTIgYI1cO7iHMqQIpu5xNTi/8PEZ9vR51iJYhkWjxT9sXtDPGV9
H51Q7zMzrx8wsfgak4ryWExkRKGB+IU7oQ6cyz/dy9wDYXb+PQJS1b8E7k38iV1W
XmhD6DMiAtFRmLBVY5oxyRhxIetGpx9BRL4+gLgunZn8rLsuFC7XhLn+8ZYA1Q1+
bESZ/He+rxEe5F6G0up4SBqhONapPkWYkIkT8fqGRpIyZNpLWJ9iBcHMYSiPyMLW
ae2TdCVKL9+IM08YNPGiKmpymrRzXBaacKRf2OaMnl1XwIX5h2QZQzO38G0pZByW
g31mxUn9dVier9PcTWh7+3HQo1Nb12aRqdt2B48M3ny+iYZnabFL0LTgDnuHwn4O
4sTyuYJv1VR6oJ9hb5eVSDhaaI042Cszaz7IrkI2KdxBEFXzx2J7QgK5hCoWd0Ud
xS5lOIk10lJR6WQgYwSYkK5ehTL38qnqECuMNEjT7/IQeuA3/PyQ5GFid4HWdUKt
SMMdTBW2bGlNT43/cWHwWlGgwqoxXEvT4Y2iOtM7TFsopfTxYtAYpwsu4sFSXoxl
wO2z56Ns9cMod7IJtV9h0vMP1sAbGGt81bFkt0c357cjxOtwr4IZT+Bi/mMudm7e
pI+T7pOCdZMrqA5A7n6DdfF7wacaQgZkc8xkzyc+vuJZmyQT7Mvg8xO+QJSq9I96
/4K3S+9s/9oHKJwD8wq+uYbW2KUd494yZdRzKSOAaOCAaw2s0mSvBtEfv3NC0y9C
RoTb8Ta+WyptbZmMniJCITuBXKGFZJ4reri+zdJjZg7OQn0EMNdgcq9jDfrig/r7
WfM6sxSIDOQmVeshIF2lKfbZBcIGd1vYZSkKj/LVW+YiWV6pmsRdbG/6Mxhb/thG
EGs3vYV452OeJxTGk7PxZz2d3MAC9f2YgdRkxi2LLLxvp9IQP1zlyUyqB4Duaadz
SeLfNdec+MNo3HhNSe/Lpxrw+uc/aNymWBobPSu11PtDLZxPOytcUa96pbtEV6AT
4xU7vhLYyVFZU6d4qp2X4WRc2u/18rNFQgZ7Mx6C/I9oTzX/s7/EzvscFfd+C7ic
FLCvU1mCyaYITVJsWfiVKo0EeFdaj9SsZK4XsBweJmLJpxhaZ6d3KBkYcFbv6iYy
YxXX1GKQwUXiGQ1qmX4Bhm+G8i9lyi9OHShEMJ1vcRMYGHYGkjaE9Rg16bdf4SMa
x4Ea1ZiODUIC08/fRPPzPThzZrfbgST5dlYZ0OT2rGW52B1um0nHPmLI9YhkP29w
fd5NpOlYgS83p316HfgQ1WcCgcCD1hs79iFRTlvh9Y35+HdJ+12sj3Ec1WmIQuUC
Ox8r9qRCjsWg/Kj3wFSGeW5HjK6pD+nV7X/gP2o35YgqtYMPvVfQypN/6uao+K0H
CZh7nW73fUColHJNYm4ZgElxoW+Ofwj1fnpkmTHiNUGlZ9Iw5XQUcBxFSpWoCUze
p7iQsN3p2zJrGm05ChCbrWSrDYpgSN/kev+bMEkSJHNPA5OWaq8vJvbit/mD/Q5U
MiorxU/44k0oiUNyE64cTtiJVs90UFDnnnI70sITEsN/o8B/+OP58yQDDpQdsTY0
cIJPTydVkns160AlaKHO/WxKHgTkWGRXmlobeZ9OwXt6t5BPt9CVOzCD3pqb3aoF
0lBvAg7jU8qbrh/uXtVFn/j+dArbONm39ORfKwB/kvO/ZC7Z+GcpO+1y/O58QkGK
G+g3sHaatL8ZBInIkvOdBt96HaTcbObhnug/EDEAmN9A2W+5dNdSEikYqT04yt2f
cJPPzBddlZU44fAcfMIaiO65prlK+kBzqr3NsFNHpJXl1hMhrF2snI7E6q/DrTHU
TlLnDQL2r5h700WmR4eTX5/Ckraj2bUAiL7BNpt/yplUw3t9Mrl8Of040HI5Eefg
zMM5VkpYgJVz81Mge7uKK1ENTepgQ9fdPANrPwi+n0WGtTBSvCiGMA8J/KogdxWa
AZrT2vwxf2Z7BYxcqfUJnWtgCeSKtJJKDSN4qK2EJwCxFJnsNZRYviO0dNQnvI5d
+Gu2UjgqPFVnSkI5nr4LkE3xdxzg5BumxcaqQ6pb8znz5vxZgDoF0289CPbCg+es
p7/Uqt3zeAwqjger4JLueQSJB4+5X2ionNCGjITajKAMRCkd+igycGAF7c4N1E45
iuI7IzoFTxM5BeKkVUk4ZHZmDcWRA6k1uBeYEREnjTzcYYCWQAh/WBBkYwAe3UBR
8+fEk4Y4fpCZPqjRtC8Owd6eUyW7Iay7nov34t3oI6xZu1XQ00aNL9E0pIlWBGQA
yt8URKGQsg02GZ3MxP773D0n8DnwImGrFi5AY+RqhOK5/wnOuEmgE1gZGKjEuWbO
Ay0zWOwgMWAwYGPlGcKnFmOF/mzKcmi8eV1veDjvBu2r0PQQ16xGmkoV7ke3Jk3I
vjYpJCiNtLtVMEJqgnAK19vdMwOPuGMNXJZQZGr+zMNYbA5YxEAsOKIeTCv1Y27f
TRg2t/86E8ff34YGsKOFcPyWPvF6l1w/oZCK2w0Z9F0GNch/deGxc2hisBynnkDO
eef5j43yDP/MrgcTCxb6vAEPIqH5Hp1/goyKM8+tjKR5QSW7Rb5yEA2D0fOg0o2d
q3+dY9Fni2TWMSLwLCFiBj6UpvIIB2vkG+1X6XwQ7eeZGo7ZiaP9K/LCrKYCCF5C
6trY8wOhrN55iQofl3gQYIZuus2fxg5nG0f59UmY93BkcvWP0BJRi6IjKlC+EpFl
IY+8paM50HMJ9g3dUa6WcG+dQZSkJLtqtRMVu5L47NEaFVCsqtRhyosoENzhPonS
HlnbbXUUtoBam0/IeA6m3WyNy7LI7/RJY4uhXXuMEItGXfE7zhgYvUSajO+ONknj
wRnXw8sYu22YdM6NvGVkOSwq2Yn1MFbEGr95EA5lFTM45N6FTOEDAg+nbqVS/64s
Q4VX8GmQ3r4Olkuc/iE7N17Ygcbp7b0BeSEkKBre+tZPEuKCh/NSRZR6hye/ygCb
U5MLtbXSRuLgwPSkFlSXD/PfxtI/QiPQ9R4DqIoUJC+2bjklUoGWmEBCZVFK5/Ny
vFRZdl3usxn/3QsBKaaZIl/1XEPNu+RVJjXrlqk0jD6hfuQFwi0H5CfyzPdHn+WF
zXh6spWi4EURmG02zBfilsNw77aIm7wgwYBiAeQ9irPs75QVp91RyASm/eWM7nmy
4huMCLtolsJr08RlQ4LaIxXG6x/C5JWcUdTGlPI2JO6SR4bqE+Bs9kah9ZX219uO
lnDfRjpxnV8fvKzW+Tsocvj/TuZmnvpDb/8qHDVswpDCMFRPg7uGMdfgOzb8LnZe
gcehoTUs1RAQwVI6DDGr+qAH1GQQeSmm/zMpfA+kv9Ow9KF0pcQJMaA1KFomLLvw
RLFCOoPNML5D8Q39D/5RMbZYTLvqASmnSbc7ZlpJOjdaj87D+/Qec0mV3kYoECfZ
JDb0+4ttJG7Oq9VIFxIxUTF1G+fcIlyxmyQs8opDtAjk9vDJlD2Fh61FG5a7NGA1
LtXmxnXV/cjyvxx0ZJov//zV2W5EGSYdL7UIXuAQFl6TTb9vSt0V/LGgw7/5pLV7
/cJiPhCWhn+BkzVwpDTlJVIJI5qa+erJqGXCdspj8UJna1ZBfA3mmPZrXcIphdtH
Il6J0uUxDbT1uMt22Ls3lcwSaVW+wDpw+t9BI/rqA/Lkp5R3DYmyGwmkvfD5PY9W
Cpk8hb3oZrFW2bA8q2eIl/Ux+PE4HW8mUS6O8FEMS5Ik+OKlBo8JSpCPRRnGx/WF
D5fYVrm3pZy7WRCnOGnLDArOoAsBrL8uLRnrYnEDYaEERp6wCCbcEeaGJPBd4z3m
CEnn0Xsk6p5QupE++RdVQ7amox0mMYY37WOswezcF02t906wfkIB16TwuQvHV/UO
rc4Q3QyMN6EFn9Z/u4zTxk2KDTJbo5vV8TWzzTBbj0eQzP7nPkZHHIO2hgBFF2xb
kO39fCRiWCozaasPmnIMhskKu0SJgpsxdK8PK22ZKe4fbspAG/5QdSEcs6K+gpGK
Z0DQlPgs312EaMR7VYEzghZk+JgkJ1Pirnjo+5PVOEwkuuzmh/NEMdPmi11kiJCE
xFPKh9HLqdenA2nU4osQ8BnZ2BrGiRHheTemOyqaEfrt7p1/32DyArrF+Xzsk776
Cuo6yDRqmEiMP+WdcVaJD3KeJPUa+K6RWNOBix2XSpGf4HpRYf3lVHT77/PE8rVH
nwEjfTmVKY8dEadeIt76xDIkaTUBt8MoQQMubXKbB44ciL8gmRZVigFx86vcKnl2
7+HUhYGFemChALsoXwk17ZJI8r/P+B7E2e3x7lX0dUBw09KXrkJkXeGiW+PDScpx
e7RDKamVzqBX0nQayTOY41vc0o5h2/PrH1imuQcAWveTkPjIRSJ1ZeAg38FkP8rL
Ez0VzFT1rIBcpKW9subW6rxWX3jhH7+TWNZuNMt7wz/9ZxmCumD5LiHeoT5zA114
JotsSUZbq2PtsOb+GcP40av5pvX+20wW4dzytGf18wIYhCOywng1nJkuKe4bPxhs
/coZsGuaDT7h3zMal8wpcjnujshKsy9ERMa/3EFjoQGrurWTAFIuH2jxQWQzoTyx
vnmMe5YH1gI8txpom0UlgFerxVnsE2jZXXCdu/BG9Iy1HbU2JSuARqGDNrG8QiFq
mz8w2bll765FA5NXuHmQGqMFsTDTyhtsc9LdYG+oY5OkITsETh7GsqsWlk4jqtUD
pihVbbrWgmydh/6vMo8vBi+RkScizh/Hu1jbS2TYOntyI+n9cwjIm6T0WUNZ0SLu
eWdJPGjCg8DFUzVryu6d0RluFBVM1ASbmmFsgd1SJDBpilpSQG9iyvnvXtwfp8EB
6jrypJDDv6sPr/YSCzHHZIXZUnoeh2sU/RFAyvzIiDOYQfrW6wgg78TByIRT3rz6
bNHZW1IaeT9vMu8ROHnxkyqmD4eeomgd7DPXy7mXfJRdU7WfBoi8ntj+O7mz3yNz
o0fdt3zfS9bd1lkkus5mJFe2w1qTWwWqw24gAO/FQX1B0JZDqss76DAVyH8M/DJU
X0LyVdTSAUEN6nU1nZampG6qm5EARnQcieLpJ/et1oGbp+pq84eUTOShYz0ZqSGK
Y7Q7hXLBaTSPt5Y3CvXugoPCsMFBodXOF3kC+lUn47+G6zBFRL4ckbO3J87ysJKf
4qwdKAZzUzbBDI/zgLrHcWq7DALhTCKyKi/1JaJ5OIU4nYW7G3qBkpeU/R8YiEgM
fGzHd1Cr90fvVOmrYMYuqWQhjoOG6DhA8m2ZdK7STz8gggDAKqItliZGpVxZe8T3
du0qdMYl3kZl2dwES6mybO2/uNdLMavjAbFxD4Bw9PC4WJpZkWARhaoYh3LfqOck
6n13Ko9RrEHCYgWMbbNCxujSagRZti0x8pVXq4SBqDR6AiM3mJ0GpqtrT21BMJje
PTRhHMB0uJPDKZoGTwCxy+eTjPOj7QtBHr0nKh3uV2HUv37FSNj8TC4Wgp5nC/ia
ZiXWEBDSePKz7dSBMUyyGDjyK2d03XynwwS76o9qNx8oSPTTLXgrECP2uRB7zztg
77EbLV/so85RNQMuZj2e/MQhDjtKFKTe3+dToVogH3vBp4vBYxA96+SqbwvotBoA
eZqIoadMR9KQUrHfxohe6p+l/MeXg6E1vRw1fV8C9um+O6zHToW9RaK6PGdZuW6L
FeIm06gXUPTKVPqfkw8jfc178VCn3Ab8a4HdrQnTL4xNkMSCVS2XeYStK9vjoJ1d
EysxZKa8HZU+mlRmCvFouubMC3j5TQwktMvGArEVZ9jM5eqKoruo7BsWNY5zQmA1
qCCUdxveqjlERRgUtpVgUghy8/l3NFQHzbYJU1mFufKUNqmKmdAKcc6+4TNSAanV
lZHUcpkvOPuMXSghGKKZCyiU49D+Qu4QiymkEIBF+bzt4zAPwZiOG1BriVdUgTmN
7GCXYREYSlNCnNGXI7KKmsdP8ykOSMBn5vcp/nzvGCuHAFNFeWA6mgj2Elizoq+g
v8/n6b7qZQfkxjvJrmCuNXYVK3i9VTECs9FjEVZLnmVDfp3jwtl0lt4vfqZzIyyn
+q4Kn+9c29wJBef0/uqQ1o3asSLAUx04R0egfhFU1M9Fk/r3l4/GHDaa9mQ7kors
mtrrxFKUR05aOTprNOOGfSc5sRL2IxtglfJulUCRcsavicl1Fw/b7U4So/OfaaDi
G50DupbEyIHCbKe6q+1ORxRkH/AOphrqFX67fyvuv16csTgc6Yb/q/JILl07Sx6m
74AuvnuY2YAEAS4J9JQ0Gsdpz0CfL4C4uHEAfkfoqy+WPUlCLgviG2yMKUVxxBry
joX2gqNP1eZVyl5bEHa/w30wwAhgBWjLDgyyhfM6JCeFFSn+qdUxohR85ubUUOCv
MtCvFrItKavTA2JryK3SU75wFoLfpl1c4D1Kk8qiUO3sFbrm385Nz4GMAsU/HMYr
nRQ4BFL0cjGdHHwgUHcDNZl673QIaG1kw/g+s7HS+i8FshpX7BlKcX+hqN35Gf/e
1eYu02SWhteQ+XwgSmIH4NkHelNLxVhwBWTKBakoUTj98n+19Il+OQSBYu/v3B1i
gby/VF+wj7yg6b3YrvmeL43afTaE8kXU8w+T5VfVQMvvlMSaQpsufFdZReTPcuva
/L+zQ/6rSAbxEgBofbTBzTbMtAvsf6CZWbc4x2jgG3P4SbzDorWrx++0PVuiC4Ij
dABcGyDDHvbWYCJUr6xS2CejPWZ1/RxBMZYLUuIY7wEVFk7an2OOHznK9Srr/9or
2KIahKRa+jgV7r52MHEccQZagakr0xrTjTmDv1NaYGakw3VpN4YEzcJsScoPZYzH
wLsfhpicGvXSAy9zmPosPSTX34KtaTgB5yhVO2opok9PaDkCNHiJDxBH8QwQ+BT3
r5OqvdPdGoRvwhAtCOQk9kzEOKp6Fckf9qwuxWxW5rSJsbFOLwKDWSBG8idrigur
N4zOpjYLkf9meAI7VtE76ZC6Be4VxPJjiS1ESYHf425XpNW0df2+LaIMh7rZYVMc
b5Q7++ECUo9C/wK1vpj4YdbGhyjM5briK/j+/MMtMlpb4xK5VzW5nA7dCbpC1ajY
twQyJMiM+5Ph6/2eDScPeLSYORJnQcZhmKv3THp0SrbM9bZ5S4wJzumS19Kp1nef
zRQQAJvXNlrge7Q/G1lm3TWqUFQUcDArcxB/v1x1vszmlKi+ssCEj+Hb7fnGKinW
GRF1rSTvwTBm3THkInouc6XrOYKUmLjlBAFHZxLqotn2owtjgbkGOgfBbPd5z5Fi
bngxyH1yCSWysGeOpaF7XyeGiHL8OqS86YC2E9FJsIPkjdQhZvribOd7Lc32ESgS
wAI5ggFaMZbErz5CPwSWF/CO0biNNf4OhEXpHQpj4aiF/cHyCYlJJfjIpt3q8mnN
0FVGb4nuL7SsyGygk+UV6KbqwC/jzlz7JtZEysUNbCChnE9S5fJ3OXDe7MdUtrGD
sliEEcXGBBRe9kBcW3Rep3EY1UkF/+5k8I7vvk0kQIpi2Q6+uxdMg9i1yqvuHrFe
xqeqHAcQYxYCqTctAHUoF9Z7ubpIz+2yZ+IcB3nJtLTUbiRqY5TV5+StPE9gdBDV
0bzQg7aE44Zkmf5yZ++2SyGKWrUvrHxJHcJ/GIEB3jszAaGGDnPkiawJHtw23rIV
DrZBWco5rXQIZqFrh/xrqvGGTgia9RWavvK9KgmqS6GqvgCG7KOWfPDa3NrK7RNS
5+/CgAYDRXnCZEn49gKuIvYJA5NK+npGrei3M6c9hO5ju0d9a5Z3ME7mpOsI9pBF
xNXZT9k8ofmoE+yDDD9Wn7eOoAwHlHAkup2DzSSiVFr6lk6nhbQqGnaz70+RTo8V
fWZfkVHurpvq714ThZ1XIXGb0PwgCtGsQGrAh8cWgITwv87cN2++XppM82KoYAe4
CoqTvo6m1tEbPQQJVJji0SDcIX+fj/AHJGii2uaR658ja8b2YVd6eZYA5XAxVC0M
3G0Ru38yrYEdR+r+kGzBm15jLWTk7FkrUQQpLURACaglI2FsqigxEp+PBqWRK+b6
GmPVCeq2x/rjrE2ulMCZ0DzB4XmTOF+/9MOr4yAn0ZC7PpssHDM2MFhrbdgNYUk6
AWpUpQP7Ojo6B4qqwcUvyWK/RiVnWvh/rxc7wIZHwXYXyM2ciQH0qwcxR3VwZKfR
4iKtuocVWt5yop68SGulgQMrITbEAu5FY68OqhX308WyNxcH8h7+D94IEzLRHyLR
VyJ0R19ceEB4GrJzUi/Ik9UfvxbFBGTAcESBRCIJd2Vn2hAQ9QVHTvQdntNXEDS8
fKmIQqv0fyxvMwBkM6W18avVOd/OWiJ2m1fxgChucl6HlhVa/7lGWe4VT5ehXvBu
VzOgMcTaG4Hpr6rpC2x5Oaa7xPAk0KeW7AtlCGp3lUVixP0GGmvV/kD7LO9gt6tF
UfqCeqSpLO1+qSYpNPRs1wm/uLmggyUNMAyE2Bm3JNxrZsLn7ULkKUvV8+pSO+oM
grkQOUbG2KpPEytzye2xloAJ7fPPH0mKmaIDn2uvkXVYLOJ7EBaLtSmqFjwrBwBW
X66fKi1EJpt/2BKABs+mbv5iv+rhWbOML3m/q/VYaXfPbDW08hdkm9u6rh9SJpa6
T4QHjXMJ0qOS7LnN0KhVvmkb/9+1/ZXfZ9zGwrQXtzagCeDVtmiTx+vgdayd9upr
Pjnjuui7gn3pAZ3gDdV1qs6CUwzTf02c1HcRfHCDj+Laym3Bwif2OC+q8f8ilfIe
5NtNaKKoPIdmWc9twcMM/OkRPT7kv64NfwrZccgDoiTxkvv29AODG5X5UF3HRKuy
J0lLKz1FWQF4kN+4Q5uozi0XBXFRjTvYkhlA2Hxu5tgCvQnD9ysJ3EEXrj/JC7pW
EBWC6RybqK1t5gGxidzNCmt+DjB7ByVUh8Vkx9Ftzk6h0riEH76k1iaXOy2O5nvv
OauDmW5mPPsNinl42h5/zc8R1L2c0OpAMANtq48K9+JaudnSu3RyWSsF+E6WV1C2
RtKBLZ4FeU04fst/QGVRHWn12njUHDAIIBwN5/4tsnAiU/R0FliO10xBn47vuDMS
RoIrGathmNaWJxqHGQZSsTlX3jd2aXcXF3YibavVUPwUTN81J9X3xnF+kTG9WrpG
ontpdhwbAHl3Q2cHaflFLZsAmgyW+r6F+cQlerILz7kzE2iNYWObKy7mtnp7XXQ9
GhIchwTGcYYfIXV4Y/RT0/6zX3tuH4hzNZNhBrWo8MAwj/IxXFoIXI9NPU8+326C
JlaD7hDS4ur+VgnblrWZxzsULVDO525lE1VeOWhbJDicj11wiTsWNl1ivsKqHcjH
jPmCsFYog8tav7fnJ3te1zi5x8PCaoNNDxxgC408bFp7nsQJBO/3pL0HEoDsqpQb
Ouf2Ni9NCcmjjyjsDzCB/hwmGwcYNyVMSvpUwlQqSx4Pzg2PovgYUdovzC0sNrnt
ZHAhTiJyWrbD27df+uXcJ1h2Q28ZAQfRTjVwbBI6oB9LnCuIF5zaGkTcvqjgx642
Sd3JtdOvsZvJXt+n89fff0bTShXASlUMfpTdS4OFVNqwChlb1IXbNupEfgR3SbVq
aCbyclZ9MIbmQRhrOQOoboONMuAXy8NHPhdHZOFIvrAGXeGCoLke5seBdUAkf9KH
HltFJSJZ48OBTprBLYQZJ9Mki789YdxzDhEhAxNx/BzWxPtN0wpf7DBRaX+X7oP0
GEV7d+SAoVoohvYVGKSd9SQS96aHPYqoonH7Wa+mo1D8LPzVIRERQuA8Sm/PrfQj
KCQS/fgmfHc7MT49HSMDVF23Idgu7vcycoHJqugYsLNwwYj49keZpwA3W3D+obAz
3lPzN+eSVz52X+oUhnAYXGmn9sqokfTFNADwtjNQMyYfck7TONU4bzACDB/RAOXU
kyEwhcsa0BxsTVscBCh1D9jEAhUkRl33aDrRgtDJ6ctENgaUVJ5dki39JVfkSd19
Rk/ztUf2hAlxKrxH41kaIsCx+01CZjSCQ9Pu4LzAo71ngDO9il+W2Pdr0j9viQJ9
kF2EJj2P5VH2jhbCvTM5z534VzorwlNKIm4BHnn5fmAHAd+irTZu4MqJzqqaJyTD
2JIh1Gv0mNl+GriyZ/yeeRXg2x25AFCwHsrJo/AQUcxx3rJTFV9m5ylzkHkFHmbQ
+RZ9YYj9dhf3TVsDCoWOBS5WCw/RI4UIt9K/cxycQXJneRhKp15gVmt8g1o2rk6w
94CPUY6buLmfVqTjy/oMZDCVKolSxEnZ6W6bv77iqulHlLfZs4tKIO8nSqwiiqqE
0COG2NpIl0s7WwLc4CxAQfKRpWOVY2cXu9XgfkANvrA9XK/A/eP4jlApWZDdIIob
1vZrvs+W7/qqgzDrtoqN607eNo9n494RZsME1Ld4zJgZRqXy6a9uugkTYumyUjSX
GNVUrCXYfna7U+IFsRlILC4XMEY3v9aC8QUYZ+D7Ho3HNfeody0y/ujAT6cIbwPn
Weo+M7Ze/vIpzWQ3cLZpY787m3pZL+6e1Urwbj/FD8Olb2XorU3wo53XBRQK4G9T
b4XsUaVd23cIKVRC8sLXf75gSzYbbDXHFMr+DbG/5/oYfQc5UGkxZy8qZEFXmE6b
3smjTEwqv5oLie1wfJLCSjuSq05supmpmlwqFwP8jJJcwrcbN4HOgEMWDjUrLB5W
HCs0l+K6GMJPbX5Hdnn6r8BHs3vwNqTnBS/yA8Vjf8gAj74TWzYXL6E7c0PqLG/L
Y4ui0uGlYS9ToYpu2Nr0mANK0Wpx6mQ+/sqXUNYzJS6EpU0cRkjx+TWMHskLtGXF
3Ve+XgNOv0Q8RjJfliZMkr7iZgvWMn4SNajFdhmWAHr91MMIal+dDrYTK9QpNHfk
vxC0cTnPN6CeYJ6yIgA8OfAt8oMe2Jogiwj+BRJkRvKLDuEJTFczn9HLsJHDCuIj
BmU8ujgzBrW50OkmNZnkN+G8ZY7YwdKyB8IspvTtxeYSIsWLWOCm+kAZoOX4+Xfc
55kVa4VjZs9yyCDe0hxwloi4nC4Lj5cjQzP2z2Ddn5gCoCSYhKCVjOu7QRFtELpI
+ppIG97+KOQen0iZGl4mkGU+GoefS3pHxg0NAZiSl+IDiEBloU8TPZ/l/VkN9r2e
KZgMW/T4VU+U9qo2s+Qfl0JYptffN16Yp/PpgItDA1prJim+dhLvtjU2QQkW1ZK+
6tBf5dsMtD1PBGD1NQnFCzaqRCq+su1CSPCYUfF2WM9f50OcOywx6x2ooSX0+tyI
yu+XLd5jFUyMNRO/IlT36SDYkC+SweSgpsDlN2h4F2LhiVS5Y+BOfqTUAncYlnN+
+mIfTZPn1nDAkFK7huQdwaT6evH1+DmFC8MR7PDUBIPwep/mRqzSDdELmAUvVDGK
iZbgQmN1kgVZtq8n0kQUhgSnPbTtdiICiIqEylSGNvTi9LroQIP5CM+UjJ7aGIFc
VMD/MgXzh+/G6UI0Ez5RwZf5JLsk75TbXWBG/pxL39IK8sP6G4ByuxJ+xocQ2Rom
LpNJpYIs2j/qEmvOJLLsqCVJiRcW662XfHvB64f277ZuEP97kPoh5pc1z6RpudUO
wrOk+Wj6uIXi/0SuSEvgC1ducdbghUHkvjCqjQfs6co/cbXU/asGfXHcxD9BlQhF
UbjJXjMAo1Tigropdf/y7+kijkQPGL/d4+SZRLYtc/kWaxnrcqHJAYLDZgCrqf/b
TQaygeCTqK8t6yr0s/DrxI+vQMyZGRgNl7m5aAShYz1ltt2baRr1pe3VsG9xIM94
AdiJqrDTk4F9cIRwzssLmzHeoDn1PlBU/rRL5+Sv5opJxvnx2OoJ7kYJa6FVibgk
0Q6Wgh1+rOYIqU18cGoi5yimhB091WG6mXmDkR//2fMX3+1WR+O0E72G/zYEDIQb
Itj8P1ZezwBA7y31mD2NMDI2pzKkDoLHKkl0WRZqPPe0eE7SNagPSxhlVQPdykdC
KdysyVYEnJfLqvJJ/ZgCanSRv0BchF/aOjYI9X5BaciYI/f0bAiB7Qx8VJdxiM0Y
VGX8+SuiwP7VZIwDQZntJsSksXDR9ES6vbuhTzeXZcyWScD3apfMMgkbWcikxLXA
9oCw3awdpyPacjLXzdMU/S1ffWv6NpDvaMtx2Dlxe/NvIOzP0GNjr5UyvObDUdpz
Or9L4ZucnT5IEZkn00aIbjfRwnF3i95Wy03nEwXqKVGBSo/oY1cK/Mxi1L3F8HBD
GtUhqnFBn7TEEuHlkppL7yt4RegZ5Lgdh1Froi27oukrVK4kexgkObtQI7juRvHC
n3xEJV+hiC1SZ4CZe7FUe6G22G0D4YDq9D2K6JPvYF8o2MlMyeGBGWfcfuLeGCaE
mz1Kiezi1xFCvFa5EYXjGJWQmj3W0F4qu6utl2SkVZrK3LznNgtgg4P786NN3fuA
30YP9X0fc5sKE+mvOmBvXj6nN1zlFHTpG6lURmub9Ca7QG2nS7EF4TWJ/nQFBvZX
x9dufYvNkF/1EH/qFByLxlYcf7vJ4EXMVYJp7Yi/WuZUilG85/eqVWa9bY2qyFmS
ZpqVdODqFFqy6ZNu9QHyEFlc17Lk75nCYfU4kwOtfiARfkl0iZh5Q7nyEHUQ6JMd
uoFjXofx/FT3ag6HKo58S+7CFcwyeuK4dfjZI1MDTXLn4Rl+UtvzhrDPcyA1ywro
yyLoarB3YmI+QwuoyKcFWrsFUW8OtW4n6zfXNN+bS3PY0kp4RvIBFAYm2LGzPaAm
41UzbOfnRCT/NkdPHEMH49+KqKyH0jFeMUzvhaPVa5L151grxGAO26KbpLjJ1ZpN
w/86avr9EVCsei+o3GuhGzavnz9h2a1Ko5gaoqVHbRMwToP6DID8SE5LNf7gRHEJ
tUP8XacUOOL43F/dhSo16duhu6ybdvVGIn1/cpKS4Zf1dji04de4rhITfN62QSQJ
IjmlU3p503YrK3zn7JMJphbnpJI9ESskNbeYHeATsfNwVyNyrKF9rD4oFX4aesrl
EhPtWqMTtf0sbZPBenoNQmbC9i0NKCdsti55JxM7sawy9ROevucTNT6pkCE6C5h5
CEAseIBgSyfSpbPNK5i19FLunHIq6DqaaUCpTRSNT8iUhbQhZJtiLpyaf4OrI+gX
1AHYJw5Qww0CA6jSANSb9I3UpPPgtbo35et/GPrmplZc0GBYKq5wC2INA1vmmTyo
cVgl8UF9sER0d4YuuifiKBMFjL5/97J87WIO4bCyqN2wl3ZihaO6oL9C47Q+gQk7
CAE4c5YzBDuf/H9Ag3sn05CVy9Tvyx9HHbAewkMWq9TNkb/gPvUqCiQIys7CiEbc
vRNkOGP5KX3kv0moWlgXGoQEPw+xfeTDOP2tXBJjtcvdqSBvTdcNNcCzs8ZJQkV/
hRsaAzrfjyqeKBmGVaim4wtgzXaAjgkdu3MojZSU3fNiSNVakPFUS70fj9QHIcsV
btbkYAQFRophqUrnPwo80AHutottUTv8rAAcki5Ccf1U12wcInE7A0is8waqtAhC
VW5mLWpoyJcWhfiH7Wt+UT/YuDDMY5USAzqCXtBQyQvMwFnzVpe6FwMl9dIH7aa2
YrRcl4smgIXzTUCXyewSKMJYAX6XCNPsqSxH3EVnj8nP+Oxaign2QF/wnT1cgdzW
zdZNSusWk+qD56Tj73a3X1g8SvByGTQMVTwUJ9Yb/xXxeCkf5/NpHRxQY1VuYI0t
d8HzogbH2h77HQ0ijEH6aGgpJ8gdYwpGwXg2bSW7HVaPjGNiMnB2XeetiolB0HAy
ds8srDT2nkwD3KDgNAN5u44ieS/pAsF8oO+L1TaPy8ARaKR6j9vCh5Yp21R6n6A+
Zmsb5+ikLvlMBaf9grY8XxsTxQdJkbjzVRVOj5OvuSIUrZTuHrrQdGh6ElY76Ew9
jJZWzW/s3ki5LufWC//XiS9vV1noLSj0RfvcQIgdZWthBL/X4dstFh1BONTCHmf+
tZdX+j4GVlG/qMBH+v5KlqRWcSsgcbZ6vL9BUo+lw/utnT2RfrcHvK/q2SzCNkAv
stQZP/dO3B5XAu/lCaMDrOlOIAiH9Q74hWpt7BnpVG4w0wKIiWim/Q06LelJSggC
o6KiZMRetHdKL3END3Z3H5qpeTa5tnLsBN2KzhyyVTaNTLmRK6AdD+Uj7PhxsY0t
MgUhxspcfVX9cNjk5Za1ZtXTYJpFXn3nn6N+FDfjO7H82ehHSK2Zbs2y1YVjqeNG
+o81Tb2fXuD2lZSsCm8scgPaLFl1P1xSIyZI0zps3fir+C4cqbMMT8C3CsV5C0nC
V5yKr4rywSqP9nSxP2QkzxtoUk7yvBIVBcUiv1pONUH/CqH6/Gfa71+yf1TvbCP5
Vg3jYvnCTJR6KGEvGS89JIbiLsVWN0Ms02B+NC3AQE+KtfPupB0KlNKNxurcwSKJ
0O4hu8L93zjm0fMs4KX9+Zvo3ZQhVZ0AlJZit3Gx5hW54Kof3KcuG84Zn4hRGYUG
cb77C/8pppVhGw9/UDGloxBzIL3TIIlKGTIDptP8SOSpz8gzV1xXVqbfK527o3DZ
IuOFiySIIr7WWzrhF+9KZQ+6DIqVi/9/JvMaXxNVtFAp51GL+KKa8LH55TelGq1Y
ihP/fIhRbm0VjWNVS5WNGgI+kDUfKUozkE7jSV11JFKrBcf1S3HIJpfrhG3BHuiO
DP4aROBC0D6LhuWmjLUzaTDSmaIMMjg0HVprgqf9TQE/uO3/3dZDqrFwbPxVWDRe
rvomPI2NiR+/AXs/Asfup4amlh13WST5ryrxr6E6LYByHb8pGBiCGXb9LJ4rbH1R
WODgPSBxP7OFcC/7faTYTrLLuLsF2jerX84CkxP9yLhuQ4Cd+OC/6GJYEa8tczle
MFozEUEmcaO5IsKeX210LkVd95ymcVOiO4q25Exbhy6G8Me69Zt41MPcXzm9yeSk
9bu7bPYnV+bHloUqRRS654ZRNgZIruLJ22IrKfc4GZB7DFZmrWfbp7nn1q3xdIU6
LmngzBaLA6w1sizTdPYevGXWFZbqXy1lHWJBByqUGEXiUK8p3hkrDxuzmSpVMXIi
lEZY3Nfq8HOandRefikPKpbz2q0omy5INFggRBbqUlcaCXwgFoBmO4zn+DrqpZps
NqJodi8MT/LgzjG2nrRBNYP7vikuGxzjZAQzGt8cIXdx7mki9bzX6JShDcM0Ut8y
frIpmLeuKdFS5vkibNBsQQrqz9t9ExOnT+R+E5G0xp6/QgEynF/qRxzxBqiGg++u
/4t8Yry/Kog/VM4ShcmbgZS0DMdcVksj30pClkPBnkw4IZDd/xMIr4X2lqOP2peM
Vmo4y5IubB4YKcgSKZewKXYv1nuHKdL1QUfR3O6D4HohyQLG6Wgbft8/fj4e7q6r
HrRZ4zburCNyhnkz7DMaJ7AeZFHKRNgfTfEWlTp3Rg2CUnYtKq/yMI2yji8LhadU
+qcXeKRPI/WQrSRuUVy4u2ykqcYntEINDJ/nGa7l9sOgxk5cWVwkP3ewXmK6C9Nb
DmxapoGYbbm8BqVyq6Nl3OQYfIpezE7Az7Q6hk9h/XSQuf3snpduSp2qAeF2Bt6d
37ZZ+qQ6ETx5UaNLPxzAamIRRut3Pu8Hoy0b3tPr6BJMXOf01EuoNSzIqz4BSrtr
9L8Oa4p6Z+p+u/Gry4Qvo80NFpJAe1EJ7PN+VdHe4LyldkxKbM3YqxwLn7oO7hZ1
WBA1ZJh8c70wt3jEvPt37o9K+j/paO6FpF+GeJejr6F4Bhmx65dWcAMMI5wvdsm2
fF42ExE6dYrXzdAaGiQOK33lvhVEx2DcTbT6P86VAUw6Z8ywgEz8qyrooNu8q48N
rHraOzfQIxhBYsM8zmnUNAsK2YxYXdPQ8s7uEa9Pzmn60iaGH/9Z9f0b4jkZfYFx
TUn8zX932n8UJ34DeEw7L0CLyHMlf8spP8G5IMkMgb92QaTyld0+hWbO+EHAT5JV
albS9HI5lvGP34mwdbrKAXQMRZQuBLFPcoO95BW/j2S+h7wjNerG0j3Ri/+7YYxD
SnJiuh0JNeJk2+AppFLvuFVMLC8nSCnufrHZz74SgYc1QMOnq87dFAbL711CdAZI
nJHT78jKft1ZCYtVrFCfSHJF2+pafvIcJ7oSYGaUdPQVUImjS54gpDZqXPYHkpY+
GeArXu1IOf+p0V6fTWtZP1wL0LpsIEi2X0ZtwQ3hbotni0Y0eDUAmPl1IqIuM1y3
Sqzn+FrybZOi1muVv3xW9ArXeOyguEWMJGJBIuuVBOWOKDqEyXMxp8IfQPS0bpW0
AST2I8Brd2E+NsU7Q6OMGR4rvMX2JSiw1KlODyodvy+NvJu+C4zegRVVQCnVMYcs
6fREA3UVC5ZpPnHVzQocbgcLfAfsL67hMkRclmAZoE3IAjYDlmDKGzz54f8NkaIw
odACGkJ2uSyaaGycfympmL8z6AqiquNct6cl4nVxDHZeAh9sBR5BD2DyIpxXgaZR
FOok+0js5WGGA5IRt7YNBpeZjRStPuMuK96oI9nPTKV7nlcmBgsgv1RmNBOjRhGX
oR1csYfTKPQgq8ulyWviCUZ1U5xnMy12jVpnDVsjhc9P2rk8Kt5i4hay57kXKrE7
RqOfWmWFI9NAaEBwv4HJaVaFeF/y6b0MazQCZU6s4R7LHypnGfsKL4BspeJfSvd8
EZQkBZR7GtMILpJeNLmcVWSbwZPZk/o9PDrAtX9ok4AVsQEPkoh3Telz8NbAmJSh
rzo6k+3zr7tSBYDKN4XJCyHGgibd+7sD9vN4yc2dw89ZQW5NzfYgfbrHT2LLfI1M
EBHub4RJn8huUebyz4FWNHwwX6XwM4VEOZQAOmrSiqxftP1R/yN+PiTq16X/+F+Y
/xiwmNgo8HW0RCnT0Rq20Pu30xJ22pFhYSlIQcc73CI3FLrEM5JNYutNkViANaA+
1D39tT1m8L4VxPbIRYF+nMyGkquZZqPDP8POwompi2/Kw2tgDnzHUMdffAirW7Rm
qAPuX31hzfoGzbK81d1rmZ/i+pgVjvfKGKRUm711iaXnUBDLlAYQEowWoN3jMQn3
k4q1+FRXzBtyQBPYYtr37gB3sRBt87XEX87z2l54EfH+2ueFqQ/M033Lwr2FwcDo
YCUYeFZ6nA+AEvIOnSA+lztOx20bWb//FL24xBNur9dEX16SrkHFmRrZWadX/9WM
Ik5l6CkKaZrCjloFC+5jXRD9PGd26aBk5cmJvdKdhZK839LfDCDViOF7JZf9EiV5
Rwniydt9bwTTCEmUGF3Ayz/DQDHPI3pPtTsTpASlXvEx10xxRWBirOQdlWI1RTEu
H+tbQXF6ZrI3GkeZQHHntUUqpKLOunFL+ZkAiR88ehb1Lt+ikKo6cPdrP31I92rK
/ES4UKEEkv+gSkTAYn9+k0Linq2fXbQo/BQAhuBPpeR4UVjwvJLwKDSobnhVbVxn
N9FZiLmgEhq/GdUhS5cvtOZQvPMR0rJZVdVH2awX1ksqfZd+m6xzRWVy5nbvfye8
FT3ZoVPcGdPqV1pcuOnwDYzv4ENgwRFLaZWel9LAVeiHzt3+Frlh6kb/Cq+CPzcQ
j0EcVNTBg46vP8iB87k4bNWwuN15AkKYVKX32ldrlWMNtyC6WLTYcWSGfJVDnyTM
EWH8WLr1SkdNjRmGWfsKsgjWsOa/vIFalWFS1b/X7WOA3qjwP5K5btgo5OrF5Cs6
/hD7joEcFRIlI2xCp8kjxZNs08bBr3+zoE+TQGw7qMtFe6p0ubLOX5oR1ug5rw0p
KdWg5IhSVDjA20e8c9pUNQreTj7xo5bh/il0ohTXmLGMX5XFuJR0as/uTW6lrr+0
ha64mX2X2jrb0y8CTgaZDUQfOtGtl53C0BSC7gDZ9Ng8O5kAr6jT0DjzOti5BbQM
UTlmcEzWmcdRbTs66rSuG/1mm0vwUM6PNfDk2NOCmy15+N6LeqRheApYHEZCBsLo
kOMnK6Z7KF4UxTCmJl53RmuOjU2JmG7HVQtGJyspyeKvUNKfPbpKUtk1MnnR4pMz
fAZcySXTbdjIp8rDMvPY00DfghkbXIBm2Vzt9gmIIS1Pu2qtw1Y8EUQvpBYyBGZD
3fLiTkqu6HNwX02tIFv0Q3iNSwFdLuvKtNZBGSuUdZZm7E2+zLtwx/mRUgxABXnH
wuvJ4Ngq8gBvTDGM+JrCdJ7IJnjnMAlOhu41WgfQKIBtGMVk4T/r5mVAjvJOSBrI
o4LsPF5KJTZpUD8AbCt2cvD5KOCkyJzE/QGl7528zTv7NKGtNaIFK62d/zCJ3AUx
APE6mLrgf+Zi7QDZ6e6f/xu3F9aQk8fFkB2SY+e2CngCDZsB5DiBq+2s4rBPBhkx
QjuYziSRHc5DLDtc1hkrPhVzjRnpzh6A/mebyVVBtX/QgzLTIb62x+kCyFjJtJkp
HZ80WNaWKSC04KUkUTXiiEQ0+OTcWs+284IXtuVmeQawsql2JVGpUfDDbdvToVCK
ieRhQ695XmRPrRD+7xuCEZsOyJDoOwekYS+Tv0F4UqJK6djJPz6FeLOrE4wNaU9s
Q2J/dGL3H/1ORlAPhYsOwBu5D9vPrpHnZmQmiqtqOkjxioA+7rqpoHricqyeYY/H
Pw3qDVgNo2p2vxOAgVyRAN7LT+fGbxP78GKimTpVyyC0jbsKMD1BpCG2DUWA3XxL
OircAyl9g9w2Mg/N079mr0dCw9nVzgxXs6BFHXuYSWl++z8IyVuu0bhWLBUKdHU2
OX13x/NoqYppMUFYftUAQSw8rLepNSg2P6OdvIWtjiwqK65pPsei1f3PFt9LKBQr
WgWQ/IS0yYPu4CEqLidF6Cen+rUkjeiyOxBYwnivr5hqeoQgs4i8WQL1rZUSO8MK
8oaBvbb7Qwb5EuDQN2QqPBa7FH40yARTg+uKB2+TAcg9VXZmj9NZgZ7EzqN8IOeg
RMGJfRnBc6WnK4Sio9l7jQr/krikkQfhe6KlG8LiKbnxubRHcFmNJUKumY2SNaFZ
2zkR/RRHsLaNxM1MzaWDJUDK2oZUOMOeqfDjbUAPkl2mLjhWKAS3RdWs0fS3jROR
W6Ho34nlBJX1ENr7vXCSPfEnaXaSC3QwouuMSWwjx0H11p6Ve9OpWjf0ux186xWJ
9PYD2QeZzYVnnu1Pe8/YojxqHZ0A2YXxBrqAMPTim5OVjlBkxoN70iC0FesMfYdu
9hWlZ172MBoZBNVLyy2oZFCA/0j/8vhnzCCTPuUC794+OVUL4sVQRf27MfEnivsR
psElSUYbPrXZXmd0uI6DM88fLdpgGFs4WNow8tq6cn7SqnWRQZ62+26vgFCiB6xu
S22RPQnc86QkIvylAJ/six92h6wRYEgRN4LZBpRKrczkCUDLNoe6cKXbjJgkZ+OV
2Rz685FZm9e9ehRZlvfuLE7vFd/NCgSyfl1AolCea1pc66xhzLA4R1Ji+5roFukl
di4jaLS2wxHIU5E9gREkPYQw97QFx4FQgH9bUFM8lQ9+RoEJ7K2pA8vVmNiorkjV
d18yDfpLcEymMZcP1mWxlwlB5v0PiCP+Du2cylXbAlog9KeNa/OiEwja4DfZo7G/
dtg610pPYV+3KYlgSrPCeutm5INw+yHOYlzSLYSVqr2jfhrcFizZi5GGe7RZFsAn
9wxA6uOeY8Z+b4leyfFs63N24mDPcMOrGONY/YoMwLhQJm9nR6tFPJT5GRu6/6Nt
gFN6Tr0pJlPyMGrULtkJwvlZUt/PSvqCOwciCWtPazMy8brQJi6VRBUCu9UVbMWH
DrOuk+CeJmpKge2WrA0v5uwQrxbNsuMPgEu1spUmvvBrrccMs5LcNlFdR2Q582Kn
3UcvPm/jb4k9QI92N/pV6p+FS5e50s7YgfimQqazxFukUtDqeKgQiQg2tJMxaTal
5Olwkaw9BVWrns9o2G/hovNbAWyrBg7af4uLnSUoaHqoXyl/xHSwGYe1uRKSNEYs
Jdusk6iWO4zzI8XdZOV2vl2SwMljCWm7xbJ313GRN6NOTPPx29KfAk3jIqRpAqne
NqF4oy8tMauU36+Aa1nCzL2pDINbZZHtJv3vzA0Z7vOj/GdCvq0l6S/joMYhvU9C
UCjtHDqQ5WLteaw7e0yAmh4TWHEfYL4bKHlXExEQ4UucWLcE5r8k2FAp21veY/K+
8iPIzUO3u67VWrVXypDOHzzIcHGoVZ0PVZXMGa/Bivf8KGMVk4ICwMT3Z8Dn+Iru
sCiApcyV5UHHgHzWjJNjROWTod7ZdXfGqkuOoGMT6r2FvWviFl1MI8L+xabjFyEN
5eVDBpYfTaM4KtnOJuQr9mlppZtpVRpljYdI7CHPynh5ZiURv1YhV+4gZTZK6836
CL6u/iBVYw+oZaJ0iY+n4I403QG1fH06pvNF3eO1eACHrD/wWA5uig3XW2ej+ZtN
/pk3noBaaLyY4cZtjzejDJnNLjmfXX+pxnn44AYBt7yfumosW2KTFckQCXUdxrQ8
EcjqKcZ6cTTQRolvmfI4jIya1+i7I0rLSkX8lcuKAspWOQ8ENLuHCX0Rbod34FMS
gCaM1UWYQ+UNX4PqryIf8sS5xL8n1G9pWISrwuc+tRZC+d2851GCv7y+eKS4l3/R
wVfD6prGE380xAVo0foKBArL4zulwKc6rueq7PpZ1nW67KEagwir4WUzuP7dsGyI
TaNqewVP4akq9WeztULjEmmHoTyk2JKrPwbGvXQv0UzycIPqKbYidmBlFluVioX9
bRK43VYI79uVNLY5WPTC61ZS0kYWNUq0j6gp7EWkE3T5TN0YygkhoquOqoiI7suX
tuRgSMZKJgzROcM/QkYxBYA2/mO9/JJn9tL/7hrYStHdD9kg//92kbtEsfTJ8OLi
iogGV7KnBE/nJ4P7r7tCiHn/fkO2DapSL8ub1IqrOSBDbTrnSdO6mAv6c97GfRL0
oXYbGyS4iE6kgQLooFxplCU2wi0Z0kffe/pgjzbxWKN+q9VUiK/VuJbWKBu4zoYE
JIhQ1ip5u8XMAa4YGqdXr0j4RD/FasqGQS8ij9tVgANBFQwTI3ccKz6+Itaslarc
RYmuk4LXJyf7/vJQYmdNclaPE8ljMOD53sR3dbt0UX0Qwn3eTVuCsNUVk9Iz4sw8
fCEC/NXe1r5VxzPn097UwpZ/pfQK/WEN8KhfyNFhHx9YvNQjzbCAu4hfkQOJVfWu
6SL0PSO5OHxtv1c28gicbXG1Ofcq4RXRBt0tt9oGWCPa5lIpXR8jxh9npdgHZT26
pyvYe4PuAA9ua4aLXOnLg4aHwRITu/9mDM2Df6h2SaqccgrU2kCrqx+AMQUZYCQA
vVIf4hRDcRHXE2mng1eHs2aYdPkYAF/JM3ayJ/Rp6+TY5e5t5zG8OFJkM562nood
Aj00+Jn43AWJZ0+WrXbWbPfIoPqodcQIYbPqX5OdVYjfUgU0Jbh6mh+YrGaLflFk
p+EirZyAX/jfFPR8m7PPD1EYTx5hVYI/JjJKBa0NUMEstmei8RmFVJ8Q+f2/BD9W
A1zaKg8boOCJKfgTorWWA/0xy1iet7tnP6NjtzsgzCkmGfQcKIAesCcVdFo2tvtm
xV98BuDzGZFiYuGG0T8D3THwBWCSDsS0+2hsHLzKq6iQKfqJG98vGJ3Vud/CBGa0
XT5R6oRlYjz6tGddenYqvBBMBuVH8g3d4B3tIXYzdu0KtCFs4Uw86uZatoG5vXCP
3LuLucSrVwhqczgviQTRPYGpGru/xWYgR6PpfZtHLntJCTPfKjS+VHjnI/ZuJiit
/XPwFyZFdTiyS3oiEYzoc/0owus0AoPxu27z/c86RGWAr9n1T3VwCj6WIYoSTvh3
sWGvJ4DMLmSkOA9cyZ4lCQp65OAPVwZtJ1oXKQoT+1OWVfmOTSDbxvJE+fz644wO
dmMLRKEaNFU0UDbmk8pcrmdPcnUYAvoiCmb51rFQsdrQxdkkpmksTm7TARntbNV0
XJd0J/Lrlp/kIeWve/6etEYWNvtPFEI9zekfPyjGUiypFr6ycCdkUw8eAIlzrvY6
9xBQsj7/RgCRCZ3cMUzXft1WhSFWdl5BGFRr91oNQwlkmQsB97yVVfUGEUV72+eP
blgj28jho/yhuFyDGfmYGA5dxh4WEboJGdlIoCaLlvbdhHsqWd+je64lMIHT3k0y
GKQLhmgK8D0OmPBJaqUP3pYjyU/LjVNLUDZ1prZ3mtUKghawx5XtfPZ4hKIvKhUL
qfWUNZR0w8yQMUIYAIaBUTKFiQnw4u0RdVD+W9oWC/G/emahJVVdInqH4SQdg3N2
MXFkLDle9QwrE5IJ2ukyl4xSVRXTowcscVL4XxbhSpkuTY+iuySDMsjUSLmdTRl+
Jdv5SpkmMSzUoYMBzOZrfs9XqmBIroZ3mkNSlFbIla/X+r5kWLTsVl7JVVbhGGgB
sWovwMbxvPi03ItCADOt6bo/f86XZzxFEhOhmB2L6AGW1LDI7Wp8sXgxorgK6ztr
zmN6/0Ge4LAXntWF1Y0jpMtwIuQfqjFAOVHBT1rSv5NDrMq2ZuLPGqRpLDNdwO0K
Xl5SN0PtzEhuLvxMj2dtT5VWqnnsCIAv5t1Vi0vZKdyF534J0sd/enwiE8cHGG72
ZAC7GKVdMWqQ3tUKBe0dZCNWGXzF6KZyqEUrGmwAZ7Kqr2tRpKc069MFOknWqqBy
a9qmrnN3rVpnKRx0E0aj/8BxxjO/GnNguYFZLgBcJA/Gnb87G2tsBERLKuq55gBK
8ZTz0tc728t6zlkYWFWOPuhr2I4wXkZGNAhLQa3cRbb5jC0Cvy9rZN1uIQEoTPOI
2ZMCLFVcJOmpQuSITS/08i72hxwJW+cAvvWciSknYjgrEB66dA4Lm7SdVjr/JMf1
Y5chOzeWlUMuFUdf0cW/knTdMo//aHQnBV4nYBLzmzUD+cMZPPJIXE5heRTMEDCK
O7CWPnUltKgZ21phu+tiAF1Z4enzY44Vu4kLdeKQlRoX4/9kZvDyjC+J6g6ivwjI
IVPEd5K9aoGpAKXIU+9clm1kbl0DQ1IURboI5knqiRkOmtQbYRdK8TuKzO2+u8ko
Kx3vs8/QLmO26pVZZI8aA75V9OIxOQNosr1iuI67nlL1wcyF+wgamVQNhYUnGIVL
OoxSSBuDUEPrpd/Ik9j/ylq/V6xKDr9MXpaO5qHYrYmQh/a0Q4LPLO3qf9ruTCfn
iUzlDplJyOd38gMxv0qPylF1wo8ClXnz/xpG0KB9zZk49auhJ6xQo6O7OJpbuFYi
OsdEvO9SGriFyi469N3Jc0Gs1A+yl1zeeRB8vzmwSWgqeSO0kD8NVtXp9EV/Rkgy
XCvzQRgDkYedASwZBAulwMNeoX278/9zk7dzeAAv7k8tv/NPgc3GWjJo0WaXKCmM
Rrr3LkAvTSdqI0Sw0AXHNrRB0tOXnNJkuiGtLNqz8LQlJBCPNa1m0LhiIt5i0ZyK
lKnQP/DDFDQyTi1Dwut1kz4C8T4T+AO+iNsf57P3L4bFWHlvURKKxcRsY5jI/L4h
SyKaxEDLxWukXUcTv2QkATVJSLIqGWVkcr3HAIxNVPJGuaoUSl3qvgOJdGFTV9WA
LI8WFmV48VIwpGJStRDc+bk9k1AasGjwtBkEOfbsqVUYSz6qAdTr31hFljgDz2E4
+fvmq1GgU/5QdHL7IQ3aNdPy7KqV6JnoqhbGL2DvbM0=
`pragma protect end_protected
