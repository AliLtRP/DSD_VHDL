// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:03 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YAs9vPuf9MaDcPxOUhGQuK5CvuNipKfx09NOJHcLBe7utxnTrGq+KJ/PkTbjuouY
eJABsHMJDRED/+5ep939Cd4KBv4231QeJ8F+rIpCHKcw4Md6WHZeesIdhla/FNPG
YWmA4XiEfRlQ7VS37DP6++PV9XHxWdqY8eddq77xtrk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3984)
SWKR5vyG8zqj54/GKsYwXOCFsm7z6diw85Tj7IpFbzmi+sBuQNTn6hBBZvRu5iOm
35JNfoTGgJYugjLV4xx0gr+mxjSppYstWaxrleglCrnR7Y3Lh8YnI09s3P0KT/C0
SVKmFET0yd840SFzInuP+XOsSXUa8lgLc1PanVSSIWQq/o/MYCPeUpT0098T9d1L
hv+VaZpll/0D9GsZ5DwpCM4U3hrxz8rLDFXpWBIJ4tyTpwvpqDoa5DUR8Mez/0ze
7kIZSFVgd+GwDtY4tudsnc3rQJK4rQQ52kLnOArXygRIXXSJQXCQx9gw5GGM8l7u
VtFL8xu89zMuhdaLYjBoukr5iZTs0J81xSZVMYUB2ZnzDvMkUQyY/wvB0kPwxHGS
nNkGV8dRWErs8QZt3uZe748O6iC0EbCS4XLY6TBLHuyDhqifiKsAr8YcdGIBkkqr
wEHp5QSFxBWNHTzUWvLJxNCg2qS7X+hSYGZVU6eoTKBbYjHHOqftJtLhbiRUWDMG
nGxk6GfLQ7kjRbw9WKLFpa+zmFEnlAlyTRGfIIbzVfMs0tsUvIzl25LqIRVJlAVQ
WUOuRE5ZZrDjbUMzN2HhR+z6/FXUHlC0tj9fas4Ryb9O5mTuKACr+XxcZf5bdeQm
VE0J0+LdPTPjuEzfoQWJ4qNN24Na2kggzQ0p4IDEeM9MdyYNDrZD7FQxZQGRnlFD
vasaiIG2qZh7bURM7+JNl0+EiXx9cK6i/7cjtSUBrlk++w/MHnuzMA1ixWzRtHRx
qUoJDIDRIt1jkyQNMHn7nfb2Ha3b+K0fHg9tbMWmslt6gigzjucEZoxaIp+yzZN6
uQzUwLAEOo2oawtBnH+5NvWD6N8T+rqxCsgsziLzgIWwEapr1oH0lYOmLi2qZin6
of9mNJqAkImvTBLW9YA/PBemHFZOdllWHmalWL0iCwVHDdKzDHND1ZFUaLhS2mNG
eDKo6aOwPtQmCEB+hkOaHLCrQFNCllxS4dglg2oEk03kfkH98kWtCW1fTIZKBKyP
K/6JqmQsDPz72SM3TrqJtUMYkY3XSqMsh5q4CzEN6hPvir9OhqIL8ivqN31bOQP7
BpSRM01wG9u7CaiB6IEe0Iw8789ZK2Fm9qWpJrrQDEOYPDaATMDukyoXesf2OOnd
52WwT+Id3igctNcDBfhBNhYIN0bqkmMSwJzcq7goptfhtqlfefHs/jZJ5i43COdp
2oJRpEKGF0Ghq109vWEdRlAZob0lUjFtyEyWhZqFJtan7x8nN7oHQ+tgW8xDKuAZ
8bhyJt41SvVrSxXkNa4IRNAg2dj+ShM1+qvCpeq4m6LIpqEFyGgHqCL8APv41Kqi
LwSgbHqe8GeVAKAl3pxGz6OXQbiTaw7CXcnk/3ueRdgvbyDQfVfoicM4brisR9e/
+g9f2/m3SSsnewunCYn74WtYAXOCKDa7dv9Hv3+gd7yRAlo/ABoQfb4z2Kyxv6Kf
Jjfe8WKrkIaOKouUS5zRQM9gHjxlMFE0BjpRWsTcQTWK9uucv/ceBxEKS0UOQvdl
Rt7KBr93baP8zeP9ZHT28FllRZOlHJVZqYyjtjUwWnDvBzP9hWl2QyEGTVxvSI2s
54KFDZxpvrDvgK4uG0l/RQWsix809UNIMOypvIve0aCEjka38ieK6pjqF2shd1+Q
qTmNBkfl6ZMUMcUoUQS7+Jw555LFS5vqfVFQGowloRAsEH3/mvZj9H9g0Fes38XG
UayiobCqGoFVcNsstFjodrV9gcMtD3MIpee+su0cBQujg+gqnii0SH9ZITfOW1R7
TX/CQyH13Yb1EaJo6mHqFaHu9BdJlNXLT8iTvX+Ipi4qHT9rHVtSHIm70xlMEtQZ
fWRPDYJc3oWzdDlG2pmLNSYnDnkdatg70BNioiUNtUGluU4Ywyrr4wfj0k9HR9S6
sr/uQRqg8o4M/ContFbux0w3b7GMGHCPWiHKbBJBziw4DIsCURs+CdNx0fWGmPQ8
XjMYZm4oqYj71uGzbnNB987gdbKAgKr9SW+l9o6QoviY6jTWPrHpBH4ZYX6aeovq
++BRII3i4s0RFEMEqTMsbqEzcwkyDEPTDeaNPrcm2wlY2mZFKIGTS2pa21Ztlc5T
/wVRqjzobtibIi5taYpMqH28g+UNiZ6/yWiZkVKMXbKU46IWL5iMtLFn8T2cIQjY
RXGopSIE3Rm2oWetQfmH2SJkFE9T4KaIbx7M1Gt2zN081oBlF0Xl6JyVb2vo7ZjK
fAIgwWRIcyUvH2YxP0JsKcCTpRS4mfnkbOezo1h8rrKviY+2OmtIDIQmS/5mQYM8
+O0tKyXV5bqg8W4lP7E7ZlunTZWEIpMgnJZTYNYjs6XM9r305QvXCVHmpCkfNq0x
sShtneQ9mlTwBFMJBoq/M9AY8N2zs8mb3l4iYZMHwpp2rJOAmkjtITxYL5gdnOqt
o3EcI7//Jpc7UAD/yH/pUepHPJdRdDheS9PZuZgxlSxfXx4syiHM6SRuEyUlhwGh
Fz8g2sh898a7hyZipRKjvJkkqLt6vW3doaTVElBmBZS+5dAoMsL3+6Ls3fjIw5Bu
s6/YLJdFnQCzsoxt79spEyLSBrQ9prVDJW33mCL3FUjJs9071TyIxg0BZtZL9hoP
JA1Xw5rWjLvTLK6YXltT4oaOsjvt7KxRDUTEb833PHzZ8vEBaV04d+W3iwO2JiRg
p80+XpfwSmVi3xviH6d7RnRMeP4BgDEdWcnmZw/13IT2BPRJ/YAOmccE3wQSpP34
tCprzGsXxofqQx/wZ9O28vmjlAWDMM2oTLkpP2/cWOEDPBjNk/GUglC7xycnDQgK
j+Otqri+VH6YwfMMX9De/M05c9o4Gpn41EyFAMtxPadQrQZKvHAwxZ1/y+hr9wPC
Qy0road5ouqsbJ67iF03oKLVdHni3qpCUTUSrP1fc0YiLENxX4gnOlrGc6SOHzYE
s9UA6+def5LgfmAXnsi/Zt3MPwn+FfeGcb8OFbtZXaZt2VXr3yTwrfqbyCi6jJyS
SastziKsURoC4AdGkvGXgKU7j4zvU8ZAQwCecEcTkICR2Y7b7sdgoRvqysYa1owI
FtdHVAXjPJWZ04cSWNlBD/U+Vx5Yn+Ao0Nw2VNiODmxyHPZjkXscTIW3zg7g1u0b
XZLW30fImmjEWUo+XIiR7Q6+76bTptJk62A4h3eeuJGI6v3BV2LEADZhiqiM70Qd
hNg4h58DyVr4AezKBuNpLD6/MHe9ePX2PL4tR03QSm3QeOPqseB9JsdS71KjD9A9
FSaEM+bQoLhrZZp+wCi2stUh87DVfrhpuQQ8cZGB+DQvT7xGeZLxS3KoAcRLEhIK
pG8szFgS/vy6M3Kg1YLAFTLb/t2GvFWF4yb+F9ElA1gbeFs7E/qNxtGsxv2Vxx/C
KAc81Q5xgGFCknb/7hx63jcVjZMtT0g7eUT1rCck9Ddv6q2i/1UuDWydlQDSz8QM
pkk4rhUQXMNoyzLsgr6xUhX3hzTriOqdMUEOUx4q+7FK58itq/1scLxim4cVZpAg
sBTSPQaoeBxCDUfbfyXi0lif/ft+6P+hxfWWxp3m6tlHbC7TTtjNb4e2tCJbeTHz
HBXGawv2OrjFO9hZLPqRw1uOUgeJM+DUE3P6i1Atm3Sjf4NWOVba5ikCRJdW65hE
cpC0YjVAzthf+MH/22lBbZxJu15AgNvZFjyVrqU5Mb2UlxE6WDqwOdjPEam1Iy5F
fLbHluQAu9dQfHOq/c6NM1oaNmR5MhV0A+IkMfBomz8uCMZ5CEInJnqCfBeO7/2R
tAjf9mmkqsO5AM8gUT8hr2Ky8nmAz4lUmj6iVUsj7QROkiOW5NquCnlI8pbkStu1
5iF7zIQmOi0wxnxSE1F4sm8EmXFZQaIez6+cCAMD0q7gMGSW6IGhXOqvnUByi+rb
AZff1QiO+QedXUXHIPDAm+sFWTwyNGb0lyR8ljWtglXQ+FstpvMw5qzskWcmC2/y
B20Sa3YOUpw/XkesjNQy5dzNS7c63ssx3rOX7w7ic6ZfFfqP9102l6Ge+yYylecz
p1tVmiRuf38ZQ/9NX3n7sVMimv/6gCbLam1COwNEPj9uEpW+6xsVsvDvvMjoUHLn
YUUDNnMvZwUBvyZZT4FEgJ5j3OsKb8gOTMpdg9bqCpg7fOMN9uF6QutZdQZSePSv
MqnyLfaHwPOHDwvk6a1F6BRoSar16BTO+TpdkSDkxRytgUywkYqvtGwGbSwvIuUY
gqqb+NCue4PZnD9bulwBc6/ZAVXWO9DDPLm40jJrVaJWL5c1Pz4njvkcqsfQLVda
KH+ZTzvCgY+gPL96uvsFv+hNukUl+u1p51DI/4B/0FnzOYRlTN2nK5En1gaeVHFi
Im/fPt7R4v29C6XHCt8YpYQzGEUlYs7636q8ADnjPBHc8bCsN1GxURkG4qqx8bh5
bu5Siu8/pleuwkl3PDQl0U+3/2jZjWtQqPiWt00/gdzfHHBNUSDFkJgT+4vzGQr9
Mq9lFhqzWKqih6/ivVE9VWgzAyV7gKpC5/mn4eJlI89qs61rGaq3cOr7EU1MRxgn
WGslRwneO87/zJJGaQFeShX+tgJUH3lgQ2/Yh8IyGIgFXXaNO/Tg9gj1rAdMw3GX
311G68ckt8dvWmLgFd2EtEsoSSYJ+q+7vifM8Uo8sXAmzm6qlocjczg9VHB5bX8m
t7Bh9kOKmX912jxR7Dnzgv9ltO7xg/ky2opn8ZF6krxnOdOMEYK/krfUBM87WY9s
Dt+fXV0VdTJwzazLJtCVQ9yqYX6g8Q2OmjV2tHUsCpS+N8p4+gnDlYtjIm3fKeFX
ZaMBrrB+Htf+S4jeQnmbR5+CCgIC/14lA7OVXSt8El1gi/19kJy5u2Vb9y/bVXYE
CZrzyJBkhQQ8MIFfIopyJR72lWUG+7RUwFdbv7l6tjC/N8UQcFY0anTVCFRvZIsa
bwXI9L4hgJe3xC5dDGn0a1hRIOtB9NnOHPzF9dks/KxRrxqMNYzv1dHzbEdGiPLX
TNGyNrNwkwEwHKnVWhlMZrhqpCl20IUuQn9Bj28Mb4SNg1c+ggIgrrSok6lmN6tA
MVGWans6kQstqTD83wLYabC9W3srtjCL7QemsZ7YLRpkYMB9v5fsQR+wXghhiHFk
z/K6WD3UBP5St5MC4PXu24T6ZF/q6Bu6QqqfEuGO5VfDNqG36zD6yJXorWz05rSV
l4RQSmun/G81U5nUXc5QH2/XymDlqPhrBV3IenZhFWARXY8kVndFAP10rQL+xYGc
Rgg1Dci2IhZE/83sj0ItDP5qXFQGePmwQVooBi6AqN7xiftFIgauQz+UrPYR2WXc
`pragma protect end_protected
