// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:30 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TYMLg/tZ79V1/ubHH/mrnjacfAAhDVn5txXLvDEvSdOH+r94U9zEU6wmacI71My8
uYl33wSTPoBXQ4xZejLyNSWhvpSPus2xKsrV+Hv3Y0YIdl1IVJ9x/hJRskt1KmCA
PRtor6v99drnQCgvx8BZ0gJJLf2tl1d5ukCKhrkMWDk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 63392)
tCXhWsanneoKePM+Cuqw0dfOHFguVZ30mGT/jCmACVUw3/P9cOIzIe//Bakpqyxz
t16HUeJPmCUGn12yWLBsEGIq4bCo9VoTx2KqsiH5QUcuofy1T0SvQoqE8ZOlhfX5
7tDpi+2vcmyPdeadsgonCYbzSMZ8bRZGfNlMOKs27nZ+yDQ/iINZK4c/gcvSS2xO
2WvQRCJn04PbgdJGihigurvMxYBsIIb72gfhfMVTZ7CEkvJgOct6HObQGYEPDvOk
qVpa1hDi+6eZyueL6UbPrBdtAZTwG9NVGlYV4zGkEN04a8IanyRRq1DdifEuUjeI
Oq3A0+EWdqIoQOVWGzDxz7+MQm/42u6274kTzbCqZ3kLsCoPlFOAUi24ik4+RYNs
4niqEzctbjPJOzPJXUyYPksJ3+yRGvhy0MisnlMwaiECMlTiQRqFRBmoUlQnrRgd
/PXkfXqUbmVwqlItLun3nBCcMS7y8ok1YCx7yb95FTOQvdE6cijQXVkBAsAjBtqw
bfXG+hqAjLLoTjdHbG1YzB0zzvKofaeir6WlBl0O2aO04g49T+A42tqX+2eaW39L
Y7fZUS4fgGNIxXEFlECIB+P4RS7Th3vURWO4gUPTPzKIBzheNupIeV8G3Cf7JgMx
yXbxTH4gbxugiPzvjLaDoqzCgjJ1Kov3r/GJTXiiyabinjvd0UUJksVHw4lGF8ja
4Sf16JHfWSjJdx0PLLwN8MEUhiyXmwyA6ubtkOXyDKB/3v1koqd+tQmh4BBnu15F
YyAuGh6BeD+4mHRCmnMATHAdr2gd20+lmZ3bn1IwYqhEXae3qerByGnbjacTcAOQ
Frb7rmcHpzuGvLvdow5R0DwC04FFuKocdR3ECRMFtNBCRJvQcxrIm6SETkWUYXUt
O0SJEILyI+5KcNVH3188CofKvLwlAtyH1pBrhSiXfcCEGoY8axWzHC2suoxn1slz
P6/1+3mBRnl3qFxjXTBXd6vKqiftWHx9E9gS42nK7JbxR888JDNFGJ9EAY/skboZ
E016SbPFPIZOZQde6zUI2xfaC3W9Z2qaj/HEopI7ovHFtOST6Qsc7Fb+HHsgWHII
N1v/5qARmTDiOfThzzrYzRCCRopCuIaZeAxLrokznfxYk54zBHUwUXbaQbt5uMZs
R4CSOcDFXA/1nxHHdrsO0KGLD5jfY9/lkp7DcU9MgDWzLbNFbQJeoB+yToNq5DDC
o8KlS+WCfX4rTThublc0EeeKRfm56kwyiCYz0HoaLVtZZEY2N9kM8QViwQvn4O4E
v26Of5mHskCoteARVCp2ex6U8cDzQIhUptzG0rvHNreSQJ1Q/p1zVXcq8J/aWpAE
pOir9pAHWZmjnnNKmaOSywAAZytHnqMMxq8RFH1DCBV1ONZ0jLwWPOp9WQeEF99x
vQCWYL0eCKSbZKFbu8QggGPXLtRZrtxYJfXqA6wOIjJN/4Uo+X5L0alNCiBELhVj
GerLCnMcq52MH/6sM3NVeJnEbiKEqXQ+qkiptfA0TN9dP0ATYnywhe6ONOOjjNBf
pmShhL+3sGvsW+w0WG/i7kvmPeDl3sWP+2nltOTmPMpx821QXHSZVHJfheiaJihR
bwJzJ6CWoEfm3KMg2veePUHcVpNDLQFcrW15gtVv3iRGEzVOhV9yMx/N/P/8QERQ
XfGOz36N64PXJ8MLZw/ntoLEmv2lfU150ZlCE8Y4V7wkGZusQ5BpATY6GoL8Yftt
QddVL5WLx9E7Bbhr0oyCKXTvNgoQqRysidpRNtfifp6j6SNkcd8q0vlsMnFJesnG
97kIEpMVksGP4yAxYej8EOpulPtp9a0neMKw/CVWui9KJF+PXHEE6axxccc1p3iT
dxaQNgVQ6cDP1Y2B1HEKKsGlVglUj1MG5yapEuMf0qtYbcydpJNeNOJNfFurrTe0
btrrTzSGLrtN2puTosk5CiYa51GYTzotwxCVokyhigXepvtP7NrbweRrpNiSYHxY
peIk1nJaXI4x2vL9wcozmpR9t22wxovAPtqH0GnI5xB24Q2ZodFP/I73+c0npGOc
hrKwD+1xcqT4wa5yxxM88/dLIrhGrtsPF6qfUmsAylGTHlQ9B4sySO7YNXDMH9km
cA0U9ZaT7tK9TNAYlx5NQ9qQSoMpjJ1a3NHd7EkNeQxj5663900OHC+kJGab+29L
EqiHRw46aYWBbCLU/VZwm993o8W/TndWQXptvyGK06bk/ua4oZID9Cj65JMYuhfw
oJcZQsUpGRtWOFwJ2g773P1CrEcNSSqiNECPpHU4OmMhOafct4HeyjBHimeh7xYK
J14V134shsWfFbEiEll/SaEP+G88MwG7brGYuv5iDJlUFoNrEI26p1HU6i5/69zT
gUYu9oYNSPeAUueHQUD43qogq7i+139bpbLoZqPAspo9NIYK/+leBVvuBvUeSfuE
w+9WSgZDEhIBb2uMLiO7G3X4lfz/KhFp9tEwEzCtkZt61qvWA1n5x4Jy5OGkoTQf
6gPoTB48DDtkM9J3ttPmR9PBaYVjXoUK1KMe8SgBx0xur/paikz/7lhYKVT7nCQT
wWhG/CGX0bjx87MLtMcVOQ/UOl/H70xC4SKsG43nP5nk4RBS2YoPFZDHK4Tva5Z8
ym4i2OS0WG4/UFpEm/NzJDsjiuRSo7sB8SOgJwlHnSsoXIwB/0qkgDQgLUkGFosk
1rLA4VXVdSgUtfAckEaqVl5CV6F5k+c+J6X+2gptPjIhORucsg1LADvLCSi1AZTs
AVmlOZTpPcl4xUvGO2QMY0fY8UpyLEFzoZYoN/jjuWE7h6JSzudH+OboC9wxSug/
jlgfM1dKcu/PrWEk/Kyfv7+nOp6EUvgf3SIZqEPjJlVPE+1DQX0THR+BdpnIK8xe
2yvLTMmLHF5l3PNwiqfryKFP7SmxRtr4ap2U1ZeQJQ+4v95eW/jz6CQEo3ue5IsW
aItvbp9qMknSFWSvcyM3xjyAxoRWe+cJ2t0+zXf+d4Lv1pAE6b5cV3RQ11ZxBSPm
A+yP+wTDveH67BWBKxO5pRALL4gS0xpBywqLIHwV67tUdpifeUkBnrGpw+zl+2cg
Q0MJj3MnEi+CS5MvN2MHTSG2RTNS3fy5h7xEvvsslz3XNkdWZGRAQrF/Xh2A0sBQ
s6ZvQ4bq5Kf97Curdv1IypEas8FJX6yQ05X1R1FgIPVHEGC7zz4MZIsoYWDKCXO1
qAbzRjSJElLHO03rFNb03gpBwZsDOXvDiGAoMdQog1jF1jUuNRKDYmc/HioGSPOu
tgNH4y2mujG9WyzcehNQo2YsgPlNFQqXTk/K53NoM8U4XXGAl8kCggugPqvBgon1
jc0rtOSqJJ6bDGfKPc3HrfvAgfXHxjzES2c5NgXLt7VFDrfAhnp1KhA8+9xUztBq
OJvyVFEPkEtZn2ONHp4/JnzqHnKpKDL3Owsr1mpEWfe51/QLHFxdjw/U9+WsMrfD
oeKSo8sA+R7ID6JYVvCwMDsitajwiyUL9ogUT+FDFNYFV8O6u8isjTWLnV5pZzt/
4WdPmO1djoR+LU77XUrmi/J1F4mt1qLJTEIX0hMesenqClXcAL97q4ntrv1deZ6g
tVMjl1pQCJd29lFd6MhXU6b4wow0Z3LBe3JqMPN14G0I6Gn+/R9oirQA8q5DcuJm
VFJcB19eHNBnERulybun7Srs1Nf1wBCd45NNGA6ENq1AtUhK9R4FcobRhDynjbEg
sowA0+WZBRu/L6bO1nAX8HUYrPgvElgS5hLnrLMwxekWxPjC+hWp2p34yK/PUoD2
tHB5eHHqv4GkFQFr9U9Qcv0GF6HFI94WKtIg2vdmmOIURMTHpo4nyBE12FQ41keI
gxC4kiBGRA/YauVPslUL6mFVIDt4sUUwcIASgDtCEm9orSyMC26WSGRum/Vll/Tm
lvBOPbp384Ex8umirmxVfagdDo9hmgUFdyjHUr9CqNIhp7zKsHDZLlSDPlI4byk8
lHAynXW/B/JCpNw/f5kwuJFxhCbfEHIm5Dv8kEQ8MQiA+T9S24MgZIK/4VE3e+fn
NawmVCOXIZ1amnc0eKuI8UgQ8jKuFlLhlqvSK3EO/EuTIVzw6v0AVO7gq4pLc+oK
FqfhdPdI6hpSVl5nlxASufxbeVuRGG5BZuNW7AGm9WtOt4pAC8W6LqjN5kIH/agy
Urqi5t+ysItr/F2xI/7CzUEA2N/2LV3Yl842Us0RANjhEq430OI5/0EIGnlIVsbq
Y2X7CqJgpDKgpv4VARMNQS2HA3iP9U6AaXU0OyEjUepCZ2RmbVKcTOcgsIHJzAdI
FijQkPo1W8HBaYs0x9rNKftUqEEmUP638twsz8T2qmS9E4RQ6fUZecmJhGSVk1zr
/NaDyqq8b4AwidPK9eTnGjPWKUClryGNv2NSNHrTgyNFOs9Rdb6wPCqhMd3/6cum
SUwbTwMi+AYw6GrcbV5SYk98XWMZ+29v7cjFY4q+boY/OXRIyguTI+lR+9qlu5I0
D+2tb8Kf+PQnHf5wX4xe3yWbSHEQr1Ag3LY2eAtiuMekPD3Pb6cG4/mmNRwcqULP
WYEWYwc5HTjAPQH93uTlhPWK2xucZnKPdkyD/hy5YU2Nu5tPWHwUTnKvJ+bj76he
5Uj3mxTNf4yHcF/QKczfmqR/30cg3jAg3Ww8pOuI9Awy+h4NYloU0ux0LcjZSi29
sc/Yd34QWQ1FLT3EuAI6fdGUA+2VyLP+I5s17dqV49CeiJCg3LFZ1CM+6gqSIXWo
ZxVPcqxU3icGPd2jwSFTaKemDNEcTrfTb/lHhcHXnpDedgWvsW6s0ZVEooBGfWek
hebNORC2XI5cW6pHr/Ww1ULTvGanVYEnE5LVXI2A89ivA9ShDNOAFj3lGIfVrtI+
oXx7hj32SvELGsLA19LjczlM5QMZkumc8awKzea5a/VE5+DlvkgcRbXCRtdgIOcs
wZLFzUZdyxHG9dK09EWXtWpITzpushvME0HROSn+JrttBELqQyOQ6VhOxMNn7CkF
5PPnQfvh4sqIb8RaqKwXX5T80lhS2S2fEwUt6WNaR0Q40YAZ4611yN7t9NJt+nAj
fTyUEQ6w3XeZTtQO+h5Z1XGWAcJn596+jQSlFoxl30C/Yg4lLPe0zs+JsKcSbDki
SEbJWSPHB+rHLTiDJV28IwUIfd4MGAIQrCC0ufwNG7A+Led25tSwtqHHroVwoIIA
zbRSU3BPoUSdpEXrdQ2kac/byGVruWFhZ18alRZdL6KS1ZlZnDsL22Y1TKGU9B4F
0HWqLhnoPG7+FDZ4UtbLAvvB2xoCffclKJ4x5Yu0sP/OwOxcAe9gMcUwzCBCuNJf
p85SxX3NnWo4R17y3EqZuqcdMkshdY58fGwEDVoEsuCtz6VhQ8Gwz3/eiUtQpDsq
etEnJA6t0Ly+yXeltPccNt0L56MhEw+d41AwsF0MlDJMROdXikJnOPMH954E0OVQ
oVsn8vMx6SD4RUhUtmAy3TOzqurEingFo+V2QAzA4BSGCc8uKnUZDf9yvj02MvMZ
h4ygHx81dVWJ7EyMaaSyT5Wh9GetBFRE8a1+0cgwz9OoGVvvG7a6mvm8180nZjF1
gp0bXZ6wa8ce2xvXxTJvwil+ypH/cM34qsyvDAGwAk5jz8Jm+antuynG47XFE44T
3LAg2u9kVHyV5j4lOkpo9Z1DaU2qYuGXGZRf9mOPK/ml+Ho68v9FlmypVsUO53z9
If+2hXa8WLM/cp/TMRxMSgLQIiOaHHaoE81bYGqXhZPsqn6pHHzk20wfG5FlnOBh
FF0D9/FUs60qv5gXXoxcOsPd26gB2uqZcWN+O9DlNlPEZimDz5ZYQECCj0FQ7Gjk
vu7Kl196fW0hLglPJ38aeG8fW/CZx8Fzg+eDiM1Hj8IYgPsXt+xIgUKnWSFRJArv
W+l6JcPuaaoZc1yqN+6JiMsnork+ZE2dGNfN3xiQTHFNC6w8dx/5+nFqqkIyfmmR
Wb/UZnQLo0wV4vRW3ObURnmUe9mfJ2JP1EAoAvxMyOpzCxLmy4BowYsCrItv4OrI
v3xocusIJqK0KnvqyVVH0qc/tzgnFbUIC/ZdzUnCdFB2Qn5xEPBhwEoqM/IHXv7I
NcN+xGKAX30oFptsmQOKxW0F1JP8tR/OjL/dbo1ZK+oyIHrKq4Lgv/d/7uuknBS9
FK30IDw1SR2QKdWdS8VBgcQr7hWErMD0NEMi3SqiCrWG0t8ettyb+dmG8OSDbHcu
sEa8x0tkG9LVdlb2dCFYkuEol2hQPAlZTd7VsDskYpEpvqvzN1+IuhZMVEB7bhn2
uO2Vq/mai2fljlChX+EElUg9hXEbnXDgziVajoTe2mszBkjEkFgIORhvdjhXGb+H
jMPz2cPCk4uFulr/wyfn9jaVvFUMDlNzaJHhIwZPQ8Rvyf4BdxKr3cQoNEDCT4yE
6pb98BZLpt/9/VCp/50P+aiDsKsQ4qFZ79fUA3pleYYe+G8TQ3otlZ9IQI8yqhHs
Ch/OXv7Bj1TpjtnXfgHeI9k2TxJD6sFjCzPg4QiSMZQjXhJ/iIZO59O5F1RoHfIc
965YSAopgeL53XZDqMFy7wP2uk0nceKKOonkFxdsOuf825iqupfBPAI5fFtyd0BV
/TywXFLFhSD1JUqLkAz95d63r6do5vOMXknKqphni4VH0EZfiYcMFq3m3fodXV7a
oG4wrgS3kS0DVMd9BB+9ZSHd1yt2N7Hqi5QulYntmn9fbo+hyCXVkqogwKoZtgId
WD+2iMox3fSwy8G4a17ZE6QmArUlwkrE6HSzLnO2lto11ozfQbduHz7iLDrbX9uc
MeEjY/aPBtk85MCKvLjSdbioZj8BQb8JYKI+jBGdoIoJf7Mrw5PCN6ADsEXx/i1O
Kyxg7+LPGV2hF//y26ZGdi+MWfB62isSWmR8ZF7UBcUiCmzYtQradehLpIB/XGww
u+T++PHdfXjsoGRmlhHRNlKfslEpwu/mUmPjhJF6xGf89b2jLMWS+zZqd3Tid0A5
RNc5g1y6FTnwWNnM6TJp7XDm9SjQ8LMEQkbcIHJUUX17beEi7+ZR2svIBYVsdKRW
dkaTdev+Q2NGnm+clSbcyC62snuzdJjh0fFqRxxhshJWejTtQFz1cNZY2Qgw+I4C
xgdtTkkQ+2n5CjJlIYg3rks87BeeqWcnIlFjSMLoO7NsBciTXKoxxNRAcbr3xcoe
xb8/uj1D9fs5D6y1GdT145liAtpH1CKTOwQyDG/OYjPBP1ynurlC88lTLz3efO4+
9zMvmEx8MmuALBWcOByJS+OawNDof+UGdIvRYnZkhI4ID1+mMUAJBzJJ09WjTeQ1
DJ17o/2H/890AZt4tlRFNxjeB1esxG1laGZMyOGl5KjgQmHBrB/8a8RcPVY0W3SP
WiFEfHp36HhzUNp41tQZ2p2S1N9JBYQEWpwsb24ruJDNDNu95WjWlLl5/hfViUf/
tJe6+SVHT6hjLnI7fKns0H6XppYfNvjchmRQvkmZQyAxncf1DTvTK2Y++j+znBA6
Bo6ojbFwwtNto3WIqfkfVC6Yfyen65irLwoSyoAF6jGFRfaaB9a/soar+jyWKDnS
iPqo63g+k7B7dRa+uZ4OQ6lojwbXb6m4lkb+3eMS000oeQXUItYhlw/Mw0vYSl87
7Fr30LRMd8F4s8zbU9ooE1WOQ57sqQ1KSzO501O1BFTBeqw85aG8uwjm5jPd7tH0
jqm0cAINqOXwcy9oH9d4E5ZTX4Jtpa1Nl1l7v58enPquKafmANixnzKDJS42oNhV
R6Fbv4kDZ86Lw2OhZFSn0E1G5pmVna9fD7zHp/YZ6tMeYnd9xEHEl0ipFm/5c7Xu
zYlu6rGqiFU5Yd8Wku7RhDbIf3l7HZvhQnumeZWeWVfBtQVAQuQ0njN69Sf8Kl+A
AwioXm3JDlucJ/XiM+2aT5pFTVlEvkM1r8MlW8046Z1xjgwobP+p/mrGpAbl2Vua
W7VUJBy+1+cVtkoXpaCQ5rZinE+fJR58y897KkHpa9NSl0jXtWrBMDc3Y8CzcFGD
CSLI61EYiYIMqFf/G/BvOFoXZOoXBxzOiLYdZK18kRUa/Xmg7c+Ay0mKxTjKH6l6
MZZeExxQuVhgur4QEfKmRq2QM0WPlm4UMQmsKC/URuCbIRCkVi5tc1X4nynb6VZh
cE2Bj7B+9gpFFCP5kpSNdV2ZJoE8yJcnOe3BEFLlyGo7mQPcqPrZn/4ZLypr0BRg
6uKteTyhwUAskNmCT/Q+/b0MbTX5UhPg7ESndJbPe5zHC/PzE9Q6pWKxul4Gbh7K
RBMEi76eA8JZLY8xrI+i9v1Cb4bvKJRT5ZFR5Hv0KHnN4NhMl7OdubpBZhOZkaA6
t9ugxO8V5GrZytl2RCSQtmr4sSi9kghI/lnHHxaS3FD0Ty9HCxgXJh/+xeLBhv0S
BUksx2OMCEZxnkjmwC/idYSRaWQI3kAbdOfJywhtzeor/YIvUYyYBe9YL5pf6A6e
SlN94bpgOpon/waJqBVE0b/w9w9gJQwAj2zqFEDdpwXhChiA0RqpWFxPdYa9dInT
STj6q5OTTwiKBPZcp4Z59tblFN499bswoRB+I3BIIrBLowauGai8+WJHvkmJC/ie
Qu+o3+8/709Hcv+DEhdq0IpUvTrUtEEaaZhEU/O/VAQpxZoX5+yER2SzELN0vRUw
j3wYxQBhZkuJB5XnynP63P7hBmIoQzwEwVbODLG4sTDjbRHTjPGVmel7H42JwQ0S
FoQnzG41BpK/OFa37yEdputQNr4/ljYsh60nZzu0wtqekAYjY9Q4fy81Tkn2k7IA
dYXZei7EPzhhKxkhLFRWmkft+T6olpvSZXI+0/FMIzz95M+eliOZ0BiiN0jGmMfr
q46BK7SIT3U8VjpmbA9hDILcvyvXu/CoQfA8F4DJL5GrkRNVk73H3cnlGrlEoWne
AI+vR6pexBekYv0RdGe8HUQG9oTQBnzu1kvBqiSE1bqTIiqftrd7mpAJYJc0FnTb
r8bti8F3iftyoZ2b27wR/zuYbX5mvvC3UjUJ8E8bBqUY+Jn1Eb+cuJX9achrbra9
Sn/MrcNGVgPcNWeC9/BuLWpdcBSaQ7hi5WZI9q+uDZtysDLxhrUw37Wj5xhrOpH2
9/JssVcg5mkM51iS6+ZnOwcJXe/cPTjCblOQff2jVk7fui416GVv9YnnVl/BjXLo
0CBSzWse8JhROsV2baDSru6HgkSSNfZs+csxo3zNa+984QDJSERwn851kSl0bOL9
T81zirRO6mzhE6xs29RK3RCci9/y12RwsuTIsM+LrTaWaQUOHmnzh4u4Or5ksM4g
vwVf5XYhYFwoAHPVNwbTMGd9tRpwPv8SReLcCSjsmjhTvFUaa0cvjxKIoZMmFCNC
5OQvph+4BWsS29PY7vRDnca2jJ+x8SGxHH3f3ramW+rHwY5QPa2xVnAJvhwyGp0Z
8kTfb+wNYGzIxTTScBcDD7SflJkszCQie8DKFFm3IxdZTNIlzyiP9BXzg2LJkuZu
vMQGB0Ry+C49+EfmkfVLigyrTeSHW4181Bujbot4S35zhPTFNIf1qm1jLC86wuLO
qBewtKUl/kSUjmKwKn33j6e1Wbq3J9PIJL8C7MD47iAnOUc2eyRSHkIApOF0cQMo
Y37ChcWGfmEMwJbxnA06+yS18Pl0/BepZNVdUCq9sJKDEmr29JYdlRidwXc81qq4
/5IGgTenZ0KWf9JsCNGmewNXqKO+HECf+3ox8oFWfMGskm6sKASEKbj7ridQEGrs
nMqPY0VRpiBgldgD0Ob0DuHvQX6m5XJEGPnPTE/hdS8fTtJNPey8KVaQyBPOyu9B
I+v1UDQfcYf2W8H0wXvzS4b1TXc7vr4wrzxA897beeXR59MQbD4qUIHzYq8l8him
RIuGzBNUbShnGKUa+TZG/iabSZ0y4ybC9xU8rm0S3/gWfVU0ygaZEMlSBy//oWm7
UIk91XLTNIyFXLL4uDhDAbVpNo/ttSdrkRkTagFtFbq96nYkMRJXXrF2ygCInMg0
NxNPMyTZSrqOfckOAJICnpCMDaHH/NkAABX4A1wlV1KmOcAl2eK2tGE8SgOygq2v
eFwFoeDpEO2YOZWMjm/tY1UXwW0ryyB1tXsVfxcYrcoDC9sqfOug8lDAGLPiK3fL
gZh1Nr0RtLv11pGP6RRNOz5w/3+bUSf16eAHSay144uwQ8q7arYsFgb8abSaEGMX
3V0E658J/U0LE1j0nIWMEUGRM77GUqXnVYMApRuxEs2yC5cj+7kf+H1c0Pju7gYO
7Pa5PQPRQ0xIuCq5/ue6WfTBxxyjPsoWQzn3uGVukZOUppumlMGmPtYRK+es1NHk
+ihYx+YGQQ8E86GGedZB9vf9h1NP3ddJhqkLV396+v6RKv9Z6vMzx/lZusO+dc4T
CQDHGSOgLpNfT+ijjbuw9MgAPFee9e3KqTdpre3a5u5qlhuBobhM02PohPKLWhL5
wWiKV2o47q3nHzkI5hH1IbS+ZwS4sCrxFCNfoQwmiikAdRn+92ZKvzW4V3kMMMMA
RjC84dfvVkb1ya+O2lgy5N7TkNtwdx69I+oPXRvkYW3lUSZ66yRHmnb2w1z94M8z
JyFmUC+k/ON2D1vl0lEGUWx7cag4DNoc7ubpe9tys5Z81P7WjG6q+uYuf2GSN9ph
Oi3o6Cuh1c2YFpx9JG+F0y49vdQh2s9pRmpX++mDkKsX2EIpsqjLeA2FUfx/HMBq
YewFHnHbL6LCXEKL7iNTYbhBweFwtBJC2/lrGHhhuM7KmY3WMsqU9LFlYtCiG2r+
oLRg4crJWXH6Wz4nKWTT6Hpm6qYl8TYk+smWJ5rmdaeLDegHcQEAbww4wAcM5Y28
4RVTlkrt8EmIosF8RGbxA0baXMU0Zeeol2cjoUcDQd5b/DpqxO9Dq+5B11O/CoIS
qI7Phu79yX06v4H8a7MNb0h3YZ37sQgl5hLETb0oU8IcKyw5fmIWo4vAcaMCmFJj
R7eUX36VqrRPIyULUxaoQlMCc4a4nnN5lg8URFmuj9LVvIAt4M4Pc5PCvDYYXmrC
/oGkrfZ3xi38qHFGUqt25sNNluEkevzvBc1TFVu2orcuzdCNhw0Vz+xrb/2ccaLr
VVtjbOalbYS794jQDH43sdv2LWgTuXysfnYsVDu3rpi1VdHZuyZ+Jegx5sV2hNL/
GLJigws/Ypp2GMGKyJBJlxpdzqRLWIm5KfTPXsSF8GK+mA1l1VS7Jn2EbaT7E1Up
EzSFsCTFgytXzl6/Wy8JLjSsdYEFTRY0N6tBgdhNk4MMEttGufwmIpu1cYFV/DvN
+GS+wE0qrIVw4FVHAYlCQnGF991Wy52n2wI0DviqCW+sC5hfXVFO5hdoYmMkmTIk
64Fftsc3HEZU7g4aEKERhjT1sG97xAV/dsAu7VnGZ1CMVnQZOWdm3m5AVxVZsyC1
jWx4HSc3fTWUt69sFz+yQ3T71biG3lhn5yrURkaESNxfkqhNCjcL76kLHwjYe+xd
Bwc1bhxiWmfDo0W2Y4+4r0W1+hPR6TiCOOheqIClXr3mlwunyZaIfky1gQAOTabr
R4hSb2J3e57iOAPwUg4rShB8hE7sd+QBUmeUnNfmkw9bOy5dnVng4IinWgOB0XD1
qCsTQnk2vVCcoSJDldQZsTyPl/Z5vtyyy9+4i94wfBaiQtKjSMQaaz7ux+xdoq/p
K5rFu+TtI/wdePUM1upjv8abHY496mLETCMAw7y538DvZYYit+2wLXxxUq7Wl+/1
fadmbVF7upduouKlrZhKmPz4zrdsgVQd3P3zxD1FUa3OrvQZpw+1SL2PGaEWB/62
S/4jJzFoJwCaYfAIulhxCVfuN/0kahmmGEchCWJe3WCAiq3uWGXF3FSW1HL96E0k
mORrMo3TDj5E2vk4RWlgKmdp4Akq4i89iFmDl9oG0UqlBpIkeAPsq7Qe21NCg1tT
Q3WPKu/b5iiZMIQl/Kvo1i9ZY47nxFtdfyaR+oCujaAoXlKcHTo1gElXKHErq+b6
d6biKx6x6XLr7XwBMy+iVTgCmnZ16htAYZ2dRt8soDohchVw7CuXWhxZvbC+Val5
ouv+YO7wAu8gsjLCYItMBSQdexr7aYvya/7dxF65W/ztRaiHuGcl0jpQKt+CzR8o
HUB9BN+/6fydHLWDr4AvmZhwylWwhMHXNV8MFdDOc0rGprrWtZnH0Tt28xRioKfh
do4JBjvlFQH4PT+cXErEcTd+e/U2/lMrNZ9VUlUsl5AJ56OjUo4FcmxSU74dgUUH
uOy9tIC9Xb+ky1wlpvSp/iiB7eE4xlvVM1xlA0lGRb24aZCnMcHwDdTKeO31xdlc
AFh/jLMGoC6wXEIb90SFIfjS5BCqz1wtif9F9ETFV5Q98CcxP72l+Rw6m1IjkrmN
oOqkgUbx5xQW91mLULsOty0JFV5zLktOWLBNjbHguHPcZWAqQpg8HFJD0zjI+WZi
VUr1lrWddOd8G8Wqiptd+LDZYwA99XIc1/JF2v+9xISDOn2f3NdIaxXNKflVZ+Lx
paHU11laQPYgvEBHbORSM7AwzlpTELRHf3BGDIEPu+r2l4ajGDy+2QQRbci/Uvqu
ep1HVrdBgF0U9yHR20XZ6TWqn8TyfGQ1mqRmuK35a6kzzx3+n4VtXrYC3YODJ834
PGgWiYll/fK1WWEb5GMiG0qfOVm1K/9qdcVkKUjXYdq0U1SB4JyhtaEp9eUxv0T1
L6RXMcMEhXixZPBjw+hFEtW4NIM87jtn6g37auZX8SbmC8oAUyRCga4KAR59wram
YZknh/HQhlaaBQr09Wczg8/LPCnjO/pI/GK22StNCFt+s4bNjgn3CHNxBu9k+Tp7
LJzR50dr+n4RWxjNMTDHUOVvVaT8Sc+uGS0Ba/HARWbNV5R09AowZ77Pn5HKojYP
giGE34hVXRnDaeY/BK5xXGGqjoIK+T1P5hJmRvWWF9+zS+6r81KOsrxexP/U1gB+
zPo6KWIGL1FQihejGI73RrsJrriKtpKlzz/yNJ7cU8nRxnwn23EG7FLEhkB42hPj
yksRDOidgwV/BndkzLUgpER0VdrUqgnkVUdRSOALHGtGro7hqBwNmmVRzLBreVke
k3Q/vyK/0woMdjEvLL34DSoWcw176vNUcfRNV8+k58y6C+SPGM17DSD27EhxcTI5
5kfQVBG45uTnBiWmItBiWGn3+NDKrQRq5l8YoSxn+CM/vCOIsswLnVI7eATIVK4Z
RY9h2Ft3veDJSr8hu0SzBoeFL3O1BXXwRxVfnO1+aP/rC6zMG1Z5eBRZ7Bo0gC4B
0luU1MP8TSZj5wQO8EhCAo9mMYP/T4o8ODkZEIvKV7U8PLdYNp9w5v4/fBLMGnRT
GJocUKlv+Cn5GSyhm6vRvb/sVtJLY318DNaTAkW0BJwUpZUulsCyFh43fx7PmsON
0x5W22SM4MC3GY/CLCKb9Y0sx35vzFDJzSsOQgDeD26KvoUztM1zEMjWig24TlcQ
AwfrUgKevRSPK7EmWVZq2P99wWiARsQAf2sn5CcjDWZIjtHCvQiOJ+VAnnN9UrBl
yEOr5rVIYrBRVJbJP0/RoKh6abk1ZmYHouEoWPndoCXjkIlOiEE7r0ntHioEdu4I
XpBdas+afggzwwL7cU/eaZYVctc/BI99DW71gub0tNEqunBbQneg47jnvmu2DzFb
rjCEFKQzCGPqh2yoq2cpMUISbbKTPkgqk3KnA8WrGlwJOH1S6OvP0GsFlL6C/iN2
SeMlRu6+QB/CXPDMhYZ7N6v9o15ZKFHKVYbOZMYRNZ8qG7/ECbAx+HMV3qvYhffq
YI07dNH/I5nqHnek/iMbFyh7CiYBxhfkTNaPdphbWcxik0TH74l3nhEJ/13LrYLV
oDzO4x0+8xRhJhtoCSV7ISXnJhfpzoOhg61541V3MEWAmbTcLVz2w5J5lZgfcinC
sBwQ5ikKPKKxLy1jcGgCy5TuBqYv+ntzzmzuaBEJb6ph5FdCrJmN1WYZICo6KJDk
O0wza3vmsLuNwWUKKkb6lVStLzf3WS6UL8z3oxzx0SpOngZmHndBoNoDwFE5ZC6P
WP1FwOU5Upykg6c+c8v9edbRgTi1Cfs6aidk+/WebbbXWpxHRTQW7BiIglOj/bLv
jmR8KOnC0fdI3c+c7FWq+5oftFqiy40MQ+BqFjLrIcdka5EzRkWc+78HblCMnuBO
oKJemsbxGmuFhOGZmR5A5f0Hsh0TI59MJuCok+gLGQZuRYuJo1b374KBMNknswpg
o4bSK6+OD6sNMgVaElTqIFOaXS4vu0gTjmfgnzCjUFWeK+qa5I85T2HeVqBG8zY1
jO6HJ4/bMJtYoP9j5Txgz1BMcm3exzm44dqZ3yXm3OlAAG3htjZCCNNY8unQkS9S
z23xP1UfYBYFx9azMC8axm66d20wpRi+IxsgUIqqcHQaX9kZICRLpXeOcXwelalA
kKEuH7t7m50RkJ5vku8YyITpOe+34mzMy/9C1daoe/DrCiYYgrYlDZo7LBhe3GcB
lD1lG5PEJVv0XQ33nDdHSbDYg55bXvDoCt1r5qJXrzsynu6hs7OPhZ+4VfToH3fy
s0au2PJ89miMa2B/KwBj1rmUkw6nbAAZ9ZAdJp6NHh+bEUzu2PUQ/7u1bTrzO8TU
YQxy0ZusLBaGu02nTchPzhBk7HFdiTyChmGGBfThfs2p8dCuGxsrmXYOV4HoDwJQ
w7iF3pjn+vEINHlDNL2VUM8RkbqRSNOQvbo7L6hM7yi1J2p8yYj3NuUH69zMXKRw
bOKEk2HKaLaIk/dZigFWIVCBqa+TTYFdfbFG+It+0G/Q3/2j29HrHkHNI5oMH482
cXidS4/8oarJ8zfkV/SlvVgQO3rVXVzoW/jH8+OukqE9SEy6YRosTftF2uswKKUE
z62dt4xnU+N+TbZNnOGFpHriHcHEgVqGxCzlja2F9Hjo4XaVm+f2WUW0RqEgdsw5
Np2TwcNThcfRWUhUjJPbChW0aIN3B/fC7bet9jl0Y8hDNsCqLYcMQW4TITcf978l
AU0y+aDeQvwJv75Tk0jRhX915rnbr9emc5IAwjiySmTtva6JrYZvW74gPYVL57k4
zua+GQnal9jia0UchW9rtNPdsjM29Gs78VF3r+UjmheJF/QmMmiKoOODA4yG9aPq
0T0mktZHEzWOtfjSoTjBLfuSr9+0XpY/nykBFRbeBbyxsIoUxH4NdVT6xjgyjQqJ
iEArnTYOyntyzqJ1D7I56w+v//AG2tuybyPhNTVdfxeFL/xyLrco/eXgWrZYG56y
d+ooCxVejme32GKSS85IvneWmqTyKM/+sEQ3Fb0RMDXJwlMNS0u0Cb+eAeibjOzr
mhFMyyfs3eWdkB0DOblPDQi6WSZUEvgHd2EPZspSRTunbKtXE6X7GtjftIWBAoKx
urFFEJhKv7QBjwxU1h3a93KvZ+txXa2C16kbRDOcHnmBIXNo2XTL4cSpVxyOc+xi
QenchwE8782TrI8qZJK7y1Q3tJz7KCrv6+U4wW91JA/LeJDJqFtz3OV7tN+fEPUB
ieMMqjMo/FiD70NcnxlHcVukPAv+VCtBkFi1cXdf7YAarK8ugya40nKwT7I0/rbS
5jhBwucK9eKpX+LtsUTPQuK9Kx4yVf9QTGv4uCKFWV1OVmsZoVZzyemAKfGEoLGL
VmNodiPorOSWvPMuBRmm2AkOPy6JFzsPnlmTqnG39uQ3WPPQlxNvybeoZ47BRmoD
6Xih6cEVmYXusPBQiJwD+jMzOa/Hlb3beDNRtGzRgq8T50wvgOQZwIZPF0YQZ/eU
Ndz/cdURapsNypEbuvjBmZzXIgbiJtqrtWYRlB81xnKL1IWWpY9Zd7STMAhwdSEK
w4SHeyLQXykZpqHNiylUUBtOmCq5IDgJr86PJRIGCxHTSV6p7qvBOVfSD0gR6J4v
8XX+5sf5TS553ZE4bZrAn4YTz2DRsAM7+9fPm0yWUuCxl07O7pgW4ifB9/x/GxtC
nB/tzR7htNhYWJlSaHrzuUbfyHQMqFy8LR4/ik1yAaCvMJSmHy+dYe3NTiCvdcf2
p7rXP41z47+G/5iP+cMthOg0b0odpRJ2WkCDjl1H9atXEDhZvJTA08NIT0rhk+2P
WdvXV0T9uq0TtoXpvZcU9q2Savx7d2kQU/Yz1UOI5PwPJmQlKphLd52qhfMiBTxW
2NGbkgJqQYwB5gv8Ek5wV9TeKlduOJAJCdWcCiDgPuqX5fTMlSgTVZwpOSFO81wP
2O6vIhio8Jkd5glUhCJiLA4zHg3JowYmMSMfqFVDLS2oMcn3wcvsL4tvzq/wF5xi
ZGgrOLDe1QSXF6RrpNqEs2oATqQzz/wQ3qI6q+VFKIBMhUtrVLl986mEl0MvhXmo
x/vXI6AmyBt6l7qfiyFvudOkRFw5apOaE4J2g7r21Sw01QqXUcB/ejNQjsktOiXT
gKgo1FjsK7hjX6XoT1aRRhBnkJIlBQmZ3SJNxfItdfpvuQlYwVK8IJOJR1kvzf3F
CsOvrI1zWHzM4zqf3jC1eeWKDn5wL5knplZ4ysG9xSBFD/GiPgkHAsB3kkA2zLQf
owM9q9X9yZAm0HOQuN2Xfuh4V4t+wpdqN3qCVg63p+dQudl/1RYzH0s4OUFQLJIR
ThCcg4sXdeCCwtli6TgeabpcKuQ2IHyP4Rdlnb7gJ8ujlpTQljvay8Jo7ocEBSAF
kKJK8mhWAvueoxQTYeaM2uJ4KsGjg/T6s4c/681nhCju08hDQ1nIle6dhWdwjEXq
JVZo21HykKqwp6II2wEuvLW5jdDhbQXVuM+ytDtQRV++GXNPIaEpJXmu3ijZmIs1
v0Hbga9UvKuQF4a/HoGU51I4yyAVwG/WxaUVGVPv7gUFFX294hEFtov2Qw4srXnI
9T2Z1tLh9zPut2+UMCXfMXM/brbjpj7wU+aPw5uuI2tZ/igfwcojo1rxrzZ4DhvU
Q3Is/GHsBo8csxbc8YqOLHWZXkpbuvhiPURlD6tH5l+BStKzOoHQaZR7qcz6yQ0V
q4qfu1aOdCphBdfniMD0iEgZlyyy0GdKvHLxnh8Dw/KoHWJ4Ry8SIPn95XtngrmE
zRtGpHQm7ajOWE16/Awyu1xEwtNUxawnVnRA2ThA677UJ2EvV8rU/6xLrtLTtUSG
Omi4LEaVIEYgQTk2qfRmTLHuTs6RTtuH6TsYUSi9D1Yv0Z7gaIRXQxQC8NPDbC4U
N4PLiAJeT2eXh40hgZdUARfoyQ2PRhYMUkORoxxkxXoP1FvBI0SzziSTT5Xk/cBh
Q8zPPZm8zGy1R9wSzVshzqEpqpsjeanBC5ULfQznJ3oIGIpnGr4AC7icFzMiFLD7
5iPSa/rBU05oipXhJnb63PqyhjEWbBF/Yqrisx6Og7fAjQcsmynCRWHAxTlbrTZv
tSQbLX4OD+ChDEphelqy+ZNIOkJxVmiNaKx7mOLAsvZQ+sKL240UHE2YVVy/yUqw
xsnC0xNJY7VR0f1svqieVSw709Yamh0PFFWpYoNvGXBDg3I1OlDZ1s77PGZNmmfq
guRBBXGCE1YM1OnsPvkQss0GNMb6oINDCca74vAx2R42VNtFESd/oCA125CSrmR+
QYT7bE+/369UM+capnwGI7l4TA+LvM0l2pLtC9u93jhRNTnmwAnMkvzeesLv4klA
Q+O17Jts11Gw15B00LhtzwxhpsKBgONPYyFwGbZKev1gJM0ghqL6DEaAc7NX5fv7
6BbkZ6dFGqJWHj/mkdKFTI/TEigK77lRlfVJ2Es6XXevOqrHVioihP7aTqaXvLs1
zjGGYugogHwkB57DCtZLhgcBsa0WKfP860DhO6uV4R6FSJWea8CL/t4yOirKFrX8
8RVPJr3c80equ9gznhkYI3wFCi46bfBPnEhJErf0yo89W6+V8azB/YSXyWkz3UgZ
bz/JW0z1+aEatzjrH2HHDn/uZXVLfMIPgSy8Womvebjhc9PnVBYo9yIjWchivW3f
RwCM41Ykc8RdkFuegfK7eWA+1KNpqctqhFDy72+RdigfZTyHRPd0izocnB4KNsxQ
TtquD4DccYDanZdNIBkgnvN8un80iB/jVtkNKgM9oppmaghO7hhaiiNLFzRMTQ6f
Es2FHR9WnJiP/2Q4O6we+Gt4mt3eg5RgdotndcqkBhh5I+y1JHcuys/I754imuIR
Onkou/uN1lYl8QmvuWLhcG0XzAdTJpv/ojiEDgRIRfzeSS+m+Roz26/ndWzCwuST
lCJ/cY3M8HJfDR/G3shkjJeE0DJe+MkDZty50tWRmjuhxG1pJTjGKkl7laQpJf9y
hzQEQQkI/HwjPz77jvzw+nsFSS5ruNjuxgpx5fa9x/afG8I/Nmu+7RRKlIqxFmzS
ozpKxc5VyotEOHNN3DTT36F54Y3U1wEqaLU9L8O8urWCGKw9/gu5ntRNHkmeQw+7
typJDh1ArgpC3z2mev5fdbPO8x9vfYxIpOH7wdlvj6L1sOdYgGrgoW1HHPFSbgn4
KLpEONdCkxTDxjqg42lJiFj4ZUJQf/KLdhUypJzene275hhLgJepMtG98Ul2tEes
D7Hc9vv1V3okLfIqQ0kaF8m80sEnnpp7C/n1ZyUV4PgJLW/tUPiST7Mjp39Ln4dl
5MJJTBE+xebqpLVoWTbUcWDrlbBasZ0qAz6dtOkR9w2b6d4wzlsx2CWymfmyv2SD
k6ANUYGpi+kI2OkoEvsv+dIUFjSeLmIvmgvRdYRrEuexZzD1KCKnT0y8umgH8bUX
0lAvjgSYit4th9/IvwH+4kZebZZz+I/ZcoaGx15PG3wN3ekcn+NMYlf18Qt2gdYp
p1pT+HJ0ruRadfmmBa1FYENt2iFFgxlwZ8ngOoWBsF+TAupMM+MEiGeP9rOL1zhK
GTDccuZagYk3tinegQzLyqDHKWYNwnI+9z//GUQSvsuDW/45I9tLA8Q++ieqVOCP
/MCO6K0Pmr1MQTTkY04jHA+OI0tz+0IiEkaICTG/pep36bQkopNsJEZ6MfaciVjK
ZO7Yi8c45m0QQdrSacn4ny46GDRtbkTMrP74GAwK6n1NsDGbfTZzfpk4zQ5D77kI
758KCTgyvggdKxnKFFQZuHp3yp1JryXCRuwW2hZybmnUQVKTcxY49znOQl1LX/In
M0N8wEZDC6s8GHHfkU14zh6L+tum1wGSYOFNI1zTN+N0GNq2dE4i0bHb95czjio0
aT4nOgteGRJxj86nLestyqoFYuohd1QNq19eZdt0XdI85VpWkJyAW15/V7WBGrsY
GEmPxAuSu/lyw38wNnFnvc7Wg3l+oHJYAoJtNq+ehCaJshLYdeifUIlMA6uajJww
YwtvKI6leaxsiDVgGSUUdtvBzibiQz193UgBX0kjWAx4C1i2Ihx42WEYKMdZ5RfH
dCtIKo/8Ke9BC0Zl2DnQ+awApqPAuAka5z6lTt71u/AmYJOg69NEyNUT2KNZlZL9
FfNB1sPnyOZbO8maXCMm1aa5gkUllzcdaxc6Czj6QocCvH9vxA3iDvkSjKsbkiI/
1JBBVbHggFxIONHCth1t7ni9jILmEhmi5PWn23am+WXL9VDq+USEMY+b5yttTFNj
geQoqyi6KDUEWYPGhOvyqmfkyU+V6x3LB6NQ7mVHX9Jg6XhhBIX1LbLxiOZEQYVB
nqcA62+9kC/YLs8Nyx4tqRYyoRdtqGRoWlvlbpT4z6ZbPsJeSjP3ijuDD68rXxWM
WNr+1HZkQZ31Q9f53SG4ZYy3ulqjKWyiKqVb4Pb6oEJwlwlmeQY2Q1GOwXjiYCH3
wT2KX4LgFo7jD7ipIreb3OgqminEvECdSovTsOHDfWO4B/fjLc3Lishn/18x1OSW
IA71CGdLWZ9Wl4NVMDZUc+bGKLCAzuYroLOGBhDDB0DuxjWeeuC8x7BK/O/2rDAz
1oc2Pt7If8rLZM77nfrVKQjje8g68H11UxUQTWGCPztouSes0p7DfT0Scb24KEl9
/pG0p7r/9ok4F76uD28Noy3c7ydtNIIka56hx1V7/raye53OPGOvmZMalxIhrdeY
WCZ2bFBPHEa01kmEdIyR4teE2Esc5NTeVvRxAtAfOznOhe5HB4R52gZEdvSgl6wj
LVvbiGI/7jSHrPZvJuQwp9beLG31Ea+wFqa/9l6wCWpqNAjWIs83sE0IzTYLGbJo
KiDZxMnc0oc49XElHZtcPU3wgCM1jeGh0i2WqgHCZWGuURVQuGxmSttus6hizGwG
USmj2ebegzmNEt2YEPEuKw3RMP0g68T84MiB5R9u2caF0QHtzHSFhiR2/WH2n5K/
GjyrmsBjMZDL0BRrzZLctsNvsillp0p3rp8BfbOHg0io4LwNp4Kc8gafNIEZ5gbZ
waRPji2zW+mz/tXWhNe/KpnmJmZBDB8NvZzpmdfIcDFRaieRcjj34CC47TCZb0L3
OeY+vgX5ymY5HOfsw8fI1b+5ucDtI61SNPaANGpA3KNwD0ICZKd6E2hffz3UJqEz
7jEU/Y02rVYhRwIaSnSlux47/ZIuBNAu5mXqezdj3RAu9qjTp9Z1865bhL6iGVqh
XZjdZLPknLAspkIaaRxmcF4HLN6vH2SIqhXC9RTcEX5SpRMuK7AXlJqPBmDA8ukZ
t2lpIQeDtJGcBR1mldfmGyZ4cmN+JKINbRcfNDsz0bDkz5zB1LLudZ8sGMi1MC62
WpvVyJCSLW4MFnqe2BCvSB387bjCpSzx58O88zXVoT+tx0upOEdT0uLzMMMtkfB9
oZEuSa3oAgAJoxQxOInfKo7XKHswjLnxLtD2R9eRvtZxywuGofs/vTWUvl833cfd
1n30we7N6ByCZR38MT8CJMRTbsVb6eSYrPsP1eQakAOUVENS+FYzqAVYY19aNnle
VJu0KhgnZKBxdKAX+BbIEwi+QTDAqIfwD1Iw5agLTgnDWRuaibCdAS2WwHjLuDMt
+zkQTTbA5G+/JJH+XOH+17vyJ/5XeGo9dfMhZGkhPFW0NRdiIa4eZMhqpPYYNiuE
mOVumQQR1z5FivQn+K39curOt0E1u2/AqDN4DOWcXb9wThxZ1bFLOh7v17u1I6G6
uJAcfFWgo04jTWNHP/Aq+w2KxZuZ01AvAB/u/wH7RaK+NXH90X7aR5W545LGPYVJ
4rjlbDLlWga26FDm2N9K4jzcTsOW2ULDO/CoOw0g7DWDMlU6SFmBb+3m9CJrfSgE
YsCsIbm41oG0l3S2CA2p40tA8QnY4i7ZpLkIRg74TliI/aglENcsHkADRhElGUAD
oYZKi9P7XD9ZFc3DIjoyeTtklSESKVJMz2k2/tSA0EqyzbiJ9fwokZxjZdRMELko
+IzniqL8Lle2QoMEzXevxA0ne0N3dkhVhHXog630Oo47q9Aluf85+YnprXE9rMMd
Gm3FbMuReiXu/p1sIOTxFFycV5QrsN2AlRPGM4DA6wxWfl/vdsVON/4Sxof+nQeq
NcQTuQe6IaklmGNqG5ARPB0SpAl9JW6M/3X3ALwXOejBPJJoAIYRMjm9d+XECZdS
D5BHo3xTx3T4v70M2CZlo28FZps2Fd3XLNDoQUzqUeR9DHTUSONSfg+Q/ROnCaq3
70mty9b9xx0edw9WR5xpWXv3HbN7sCHZCnb85fOUNrR6oiXflK8Mv1x19IXRSZIq
DCcc+lNhp6HhjFEdTsre9NCaNY3CszxVvTnbNb0lLUHBuJEG4RhsYV26AsF4Ae/3
QMIBPWowJ6CZgtOtPcWU5mldG47OgcWUgXQk7Hxw3iGo708tT8PfvsGE8C9IIbPw
Qkxi2KYUALT5sT9A5gIi518tOMEh674y6WfMXKLOPREfBnJ4ItKVPFHC8CsBPft/
7VSgkJZIvpxzmcTluTQVwo+J65TRgJT+buF5TLu03JLluIGhf+nBR1Mo67Y7ONSj
h4l4cPvmdE25Ay+C7Y85fZ//+pvANWiM6vnhD1R4h2/eF13cyUBwZ3QoYwAq6EB1
NQtt1H5+YfB5jHvUiB5ZqyZmvXiAlCu7XWKXUUfvvuEUe7B3SFRX6zgZ1ixbNuBT
AnxRFq266pQzps3y7jn424vYRfLVH0B0P4g8PSGKSK3cSBttGTwMKpmu4pwLoVW8
7qH4PqoqPlfCa5s5BhN47TQebLlj/yAYmp33s0wxCcoVojpmfJjDwHaY4xlldqun
86GFF5c1O95SbacYygSPXhizXbo1IKHX8ADiMoPj9PrKKOrNs1HhIDx6lF1RrXj0
GBUfJr/Uql8ZmwXBB8aWoAH2bM2YP72I2d5V7QRWlfVGhattf88qSe5ty+fQRGBM
bqXMSvDvwK1TPteXaglk7rkHr6hPSCB5xiQbum0UNaCTluvUW6GDSmbgU9AcwCdf
CekOv3lvppmGF7+RgXqOmlQiC0YwtYc0EBi65tc4mw8s2AG9z2y+XGGKKmrGdw5Y
YddPk+E3LsjymO7zXQchWPZIYQ3oAx3ZZxxorNE8n4XD+8S7Py9jwVQYGxmisBWI
AlBF4F+AUg8FBih7ftWBIe3zrlJDZklVvBSe4h8s83+KWYjql1J/slutw14/Q0kF
LwU0nl+L1Te9z+qO4DUbOIC0DA7S/tZ6B3c5l7ij9Z6IQD2c71ffHDeINupz4nyY
CdhcXFayp4/NG5bTUWC0MyLx1Jo5rQaqV0jWcpECxcFCSX0uZfskzG851yFpXnPs
lR+mTZgwI3tzQmWCtqIUWcbNubu+j1zzg1FGkQAklXy0jmIXxuGi5SZTjt0UsdQe
qXtSO2gIUfUw/B+F8YOqrfURGvv4NNlLReC9aJit7emy4qiFNCxAzdBfmE6pEidg
iRuZqYtSzPh3PsKq9vFEfYYGO4zgOStxC7m2DoahZUxKc6r1ArwU1EMNz2pjW2VM
S6hR5BcMESnFK3hfQQ6ueRCwLbNuUvReQn6fBPA13O/ITUxmwQC4FK3tqt/l93lw
PRyWyZZBF9KGER8xph6CLAVTyQvdlKxGfegu3ESMOt96qPG2cBpSP2oh6lxSjIlD
Al62MiA/He603u51L3HEzdGIqQtZiYS8tNGavECQ2b44cW5RREebHFc3mUk4SPAA
Hes+bEBt99DC/0VkSQYjLo60lrEUhcwAetfUnA0Fq6G8iIrQkG0P7zYquS8P7+Ps
J8imiEHgqCmvDegThoHukhVBf1tZMenZrHI3uxKUBm3fvelPSDeQy8Ygp1P3DgB4
ejnk3wIDM0WqRY9qfDCvM4H6ExcVp9gqsDTuyt4tocdE17OLIVDzjMlhQ8wuzbUS
Ud2HWCUtrU/LE7g5ADSOmg2pXbejo54YcBjZMtWzdDoAi+deXEwAG5b3ymMNwzcw
2lFvaWfewas1JEv/Gv1KbRKynRrBDJNwWfgxEgnNSSjMZYQSfbO5AiUhIsm7gdE0
KMXux/KcnPVNdiO43uzBbHDHA/KtTngra2YB+oGAd77k1gj1FImjyLxdkXoiv8LD
6yTEtiaYbXxN2VylpogBene46jPhFqY5s5o1CsbetlT2cDNs06KX8dXOQyfJFiBY
d4lYmeF0AAH2xR73VlO5uxRdNizwk24e+qHnYsigLXMmykREtIto2lbG1fq96smY
T128EiYyABah9Czq6IrJ3N17UYjFvuMZE0KSw+lv31dN8kgR7161gqQicMug3PQh
Xfv+x3jWsXioAoOgSkXfGfHxnk2LVeMgLNRmtHgIbP1/d3c9W3x4V3cbKyXRVm3I
tup2uJVDpRuwZyDxsbChOerr5pIsgU1+wnDCyRAenWKE7/HfMWB12q8fol1DmUZd
gt0Gy6ppVyRXX32lC93SjE5p/3d1zS4VcglZhDpPJ0SNlcKK22sAWCARHkY5SeDp
f5B3/JcGFC2Fz/pnq4C3g49IwA/btcNiXprh6mJLVx7PajCVbTG1fDW4NqAlk1rX
S/wWHvv5XOny8IuhBNVnDzhbEZYu6BG11cVAJbJZvxK0BLKjynO/gU9O9NAzA0Rc
GTq+6GNNgsQVMYP44+rSMw6EK9rlkMNH2t3N9JWvH+bNuksjdqad5C6y5yLuTxax
u+SmqY0aXP40Ozbts4HyZ7O/KsbCAdfus3ze2eDEhl1PSvHtxA2VLsXCaAApbf/K
6JYrreezSQHlMNX5zVxprkFUB0K9FPCyWnPTvAjZyDMxY1xKZryomIg7spT4QvH+
ykHN5jw/sERBLCZJYbhyoLk1Rpj3eVmlrZ6mOTw9zhC3KaqpwSX7kWRy/PDhETri
1ty6aaevLFod0rVq92WQP+Vg/1VvIYYVFHx4Q9nJw1Gm8yLhCWbZFIY2vOimW1Eb
QvWL/edCbLVtn++tlHDPfAWRhMmJaxR8qM4K2yq7y060bD6y9hHsLVIyLmLTuXY8
KT8h5i2TOKDTGaMOnYiIPapNrOJsey3ZL17G23WArIDJDFqR0bwuy8u6vUEdfNyH
oHfqM70QInr4cmIkV3k666MYZ7jKazIhQzylGFuODgxIDuPWmKr8asbcXELY/VXs
ffTE/WJx2cGnHErkMTYvq2r2Cref0IgIeptEkL93uVLEtxHjJzVnVa824N61ndf5
hjxPPNC8a8UFo3juxTRMmqME3/p4x0BESOmnir0bAktZsHnCtbd3fGkOcwTSSnM+
pQpMLhz8N8mrpDiJh1VTXBvBV0I8rJdBCyfS0E9BDkwXgJM+8Pn5ttiz46YIgKRa
/cjYcOA2XpFFWZ9pwhKZ421MSDL2E9kW2GhhCDJ3Edm3jZ/Nq90ADWeJZg7tAn4D
uZrn5fquW2Tiqzjq5zxknvzWH8ELZKQd0AydSJ6/5dpMbcMoCfrV0AUiPlfSWxtN
dES/Ga/0VXulh9uWV5m9C048YWCXU/CngoMRDxzHNoDLD+qaTrnD54Z3CS8M88Su
EJaBOo/7FfPftRCDdsRt8rTQkkr9kFP8kB5+8ch5LdpQ468ZLGVPEdvKH9NI3iQZ
4hOs585GiaPAJcPVdIKzUHmit8beBMWgyTvyIdcTjhGYT2rhYhOBit0YyfqUuxkv
G3NtaSJPr+mbt4azLAR+vfffluTkoo0e2fetCncd50Mr2aD4Dcwc+oPtmyoho8kX
x8lAyDQQQ0Nvq+Gz1GAtbNW7ozknwR0xAfG5kOFtX0+ZRmDZ5rBNU8DevLpCfY9v
AOeLeNUgsUyvsEnR/pAZqPXLbVPwl/mntLbyyMEl7aTYgb9KNeBl9Q6R0xyDhd7A
Sg6HKGSs7twAd9HHC0IfYV7S8bgYCDovXmtygEZ1fuCeGUPfYVDJsLAYwAHHbTTD
ApKfpL9qY6UWikf35R7tIzAdYYnz2cs70dNnm5k2owDIoPBTIHdARItMF+wQvI88
JdeRLfh2TL7nCoyx9ssM+iik7usdkU4G5WdmvGI5k4Sc3/K/DONESSWpGIt1o/qP
GVkNJ+62YtFkSkcoY9n2SmBx4B8aHfcdXdZTJiMGdyCoLPRIkuflc8W6DJaJqTWl
01+sX5USJPnELG7l4alMsOUgqwruWDDOB1SdkgMf8rNtJ21vHQIn4VWAuz5+9aXa
yqwVDplQIsT2QPh8m49Kj2kLd7NhZhflrSaPfK4O9EYwLtMLBpbTFyue1DcKehpQ
n2q+xeDsBxsy9k+CMPUzrrGhr9AZlxH+S7VYSymoWCfiIJqORbOxFBPHPZlh4Xj9
LdPH+F5HKQ4nhsV+3hplfjHC7HUr6KJospbegzQ4FFRTc4PCxSxMVs5XSlev+pUW
OSIdnUTo6nXLDsmlQOgp4eKNancJ10PlGxqM6KgDgzHA6RlOOf1S6Ml61y5HTcHh
hV4VCtHFTP9cck/TnP5Lwl8XvZ9lVVoCHafZJt8zK3nG10J1nbBn19vCc6m+jLRr
V6uIOg1bnPpzkN/e7M/MjwOCUIyRSKqR2W1YpCvfEhPT7Ng/Uiz9mH6OKlw7cdup
rct8vjONa+aWJ8ZdkNOo62FrtlyjD2xYE3arl4wu48lxAABlnNvpK1efGEZIwoOX
4tNy9se4A4DciGrodyvxr+c6IJDkI7ROuyPtqlzbfRPVyhFGq9UGYsyHmjoMHyFS
kW1x4iKbltjsNWMzkBuDoyVnuNwwqGhYyD5QjOC93HxTj4KS+dqLEqm/Hp2uG7uZ
e61t9pHUulQF5NxkUg0bd2IBCgIBSd/yUHDNDb9zo+y+u83uPzIpqGjxClE7N1iO
pvrgmtZ2K1cocAIzHeHSNSM11yqElL3ApytvLgJdXxBkl525QMShPT1XJh7mCYEq
qbrfSxJu1wVCjGFIVzs2K1fzIuKiMax7pUAaSvBhWR4qd2H3waJBAJxzG46j3g+E
SarZJBj4QApiSz7X1ovIzjqdmuRavIErMqaLoRKoXRXjQ1VKsoYmj05tS3Lecef8
74xEa8euJncEekZtYsFWaDciFsjIytLsU1r1s4sslNPyeJ4BNNg/4NC2c3WycatO
NXx0eZVQP3Fd1Ajd02dNQq7bMDdh6v3xZe86bSSUeP6oHOQiEEX4Cx1rCA8csi6M
1Zbnvpo+9rh6jOMbObkI1KEhjIjfHGYy7+CPfIWGPJ9ZbPfsJy8qUmHKnt2YZk7/
8CPyoMZ/sAlr6FkTXYokr1BAThH4992OaR1VQnuoGLsJd8jlqi/03et6yHblk8sy
rwVZiw11DZz2yS2IuzbJTSYf1ADzxhWWFUUHGINOXE1lD2dFM/PoQVKSih8MWXxC
Adh6VIkYYsWCHZTSZ96g5+zvQ5QZEJz0e/T7O3+eeN/hJ6iAZUWcpeJehNmrUh9y
xiyayMvdE63Gx0SKQSuvU5ycenB8CP9TsdiVAPpinrjJ8XUn0zC00+LcpwcB71nr
dDgXVE2MQACvtDHKHvXJJZc+MUBCdbuyS7+XfriDjtI1LrbOO6lO2jFrrrAgtwr6
SAkZWbdLxmWdshDX6H1In5iVguqoP9hfqJXWVinl31t2InshUNdZPsQqcDPkCX3g
7ApSbF6NjXuyDpw27z3Y4sBvrI3TEOw8tSE/Xi7d7C+HrZhOnR0rGOqwjmxkdtkZ
ezE9mlzGlkaWBybrHKl8Y/m43D/IFIz3EftpG6tn5PDFyrM1nCMdA6ijZp+7BlN5
CuZCPFtozjFMwFpfLcRLVu+1BkGZvym1DB7vu/n6eQknue7gSLL6AnI9usqqOy3E
qfeu+9bBf4nwTdHgvkGKgPMYQqmR892xifO8oHGuFNAi+mETf9R4ZLXFOz7m3mkC
kUXZCfTeJUidvI8I1bzRMhvF9XhFj5Ii/YVswHgZQKOSIh22EzzZSQ7H1MEv21Jf
2OzzoWqZAN6FCGweD3UFpWJh34NieutWCkAt9i3PGvd7nVjXF90XL06ovagNCb/Y
lmV9VQx3kn4JjQ+crw777lH9N3XiQ1lsUoCjXiRHc8Kv1G1oZdcjnI6cyxh0EbPz
MHDaNusbx4kwHeuC5SnxRPh4ErcxqdQ+Zg42Ew2au0C7nsQOGt6FSjypyKYKgLIx
wvFEr3JesgIwEG53R0Ncs56BaDLsIAM6DEddje9f0FwQxJd1hO05Bu0KQ1WwWf9u
8M/2OoO/Anl1c0sBeJ3zeFQahwwpOkelaABwBGwKhknnBp9CMTbh2KkPICTVCC4h
kl1QbcHDGubcpXhG0iZpbSGyC7tCin1i40T1U27rZzliL4ofon2Y+JhQlIr+t2rX
QZiyzlNgZFIqAhsRt6pCko4BbjXi+WP8xoUK/LuncwMBamOfsIV97ap57OEhnU5P
WJlNCRSGYL/weauY4Rx+T9zMiAHB4Nbf33mCPmYU1ELojpkyVvjws/Gv2F8wlnZ3
BTsFFkbUCWq4soKwNQCSrfTyi6aOheNVPOrNujh4xi+eboYmOsWJxbZEy32zeBWm
Jh8SWYxae0EcclyYUko9KuvJTaf1jXZpZAj3pBOuhFQyv3BN/Nf7M8r8CGL4mcUy
NhEM6hHAHnSc2IbBzdE7b+9+uB/Sg5ZavbQhlpKgH1//UPOwU7OvZKmvm/lI53VY
CTVJCwW4+BkrpHN6eXK7DXkqdk7KCy9jyZXr7itgRPSL0FkFtKulggEjS8pbIyDk
wfmgkIM0DRrOxWfYbqeVRqBprLQX1n1Px/PO9eEMJd7WqNll7ndt6hevxTJaYGmN
RwM8f7LsIsgvQ7wH1fH3F5T3u1nJ8U1UoTzIsuv2f0tMjC7KdxwHEsz9byg8m4kJ
ycAIX+vwHJI3MSn8EftnFqJyhMrqKWuBbp+AKl3S80MTa7ITPkHgb7kaAX/SOo5a
RACYIDbYWcaMZ4dJlQjvT1hfWpRHRBtXIv1LG1IxUiFsJkEp9K/jVLNdWlXl4Khq
CpTXDVCaKfIt2JnSPzyobczV7TpPHtuSgFaG+t8NDOimPfJPzl//KrK0bGsiHtgA
N3INMXk03KgLPn2D1IsIR76MSzhbmXLquy38AN2Y21ZJwqiTGqjHzIR3qBMQqtBJ
ImuraAOTSeBAHa9Sm4vHY+5PKGAeAeakIw4bpBqSat/aE0W9r0dlTAHHKFns1P6Y
wspWz8xPJ96EGFDuJ6nbAuIjU8Q1GatG/6t3GfIddIdF8Mfq/Rnl+IVxUdO2chU7
DHwE4PvpRgY0m3NRou768hvoyPfvFwupj1CtxEPy4cJgUgpkY9CRbN2Gpu9lyZ2j
I0U6ameEkqCl5GWDlwhcVoVYuTWl/B4ZAlUeoDIGgaCGn9NQnR6w9uxrEW4uAfpW
jf2Nvkm4xukNIdmw2yNL5X8lw4rR2tpiX96xG6WEldQPhiK2hAQUALcmQ5d9T/my
txkMKMsVm4PPeTZRWN4U2iNKoeGTfrUqTR+89cFTldY0zGe75NbejubtCrVrxkpz
E8iOp9pSATsQuza8Ba5XrhopKjdB6yEktFhOv3uIaOuMidHURJQYZVKee4hxKcw/
1uIQhrUIoqwuwxRqqcNV5Q+aCSEBrnXtzdxTLNtWSvbuN9DPaYzNZf/838c3GiNY
Q2W3eii0ksTN67XUAfdRQnZC333W0XyWuBRyEPCfPc11GZT1blWg0kNG92jBmr6K
iIoJ/l+KSfkzJ7tVjXJsqZG1ViNfh0F6sqGkK0L2hxMjhSOEpYr8yiJIuMrYwldP
1yFEUpdQjkf432Rbd3XCwf3d3MYZKtTFuesJY0LLKy1WDzKTnTCeE9ugir1+O3Ks
+QwVmeFtkwlRqRmLlwS/RTUCJjJWPAxwrF8Bq8/SdzP0uCYRDzjTpZmg+Ono5VMr
fSfuYFcuEH+4JH9MPtFJVIEX9J5QvbVXF4noS6KIiSj65esKEIqqZZiJ6p/nmme9
yrBA7uIuV69uPcIIBY9Yv3Cyuq/lUtVPKffKAVQAPu8lbKZIzH+W5Lg4ASPyHY30
bJfgggHzLotQ40pQev+6DSi9WpFyi9BLNxqu9/O53WlfCDNqDE+fQZNNEcBdn2L4
AaAbXdxEqwrwHV60jhDgJRXxwJSQIlR/JkymXVlU0COIFQnXd6wu7lvsJvtX1ERH
CVno1mSRJXNi0BneuzdVh7yogicSZlOIEEeao8mvxQ0jcprcsjY6lNwC6vubG067
8tLvyB11MZzoDAJ3wBgFkBBhtuiK2bhJ+nn8Y7P/dICJsT8I9kq4KntSyo7SmWDI
KwjXQYspjlHVoWfimNIPvWk95dUBuL7MvVKFql+zrj5rcXwenxNF41zd7GzTHGOR
hD6/aTCcrOk4fxRuGc5CnduV0mTszF+erMO/yYcwHOQNXp0V/mLuA7NIHyf0UL/6
bn00CvguDAhP+CW6v+tPul5QXdDUEBEvlTnVcD6Ym7qO3636cjzVSLc48WoIJiSz
7eC5+GB20Yuq9HbJh5d/nc50hGAH0tGysvHYt5O4IVOzA0CxPvduG0bV4Rp+cUaJ
iML3fIxwWKYCU3wNah6LP1uafhK8rQmQ3BkQix+tG5bnj9OfQwm003ahH4yOLgi3
4E+d83niU6ANdl5mg7NvQvn3bs6P+N/dUj3xGoXmqI9pQE/8Q/J0HWhuGXnY8ook
nrkSgi4UdtUZ5sr5pbuXefhWjbtSVP1veyyhT3SRbWNxb4+NJ05gBBTU3gawir6W
OqzxQV9BsIx+Af8XnzJAZX61vp9z0zheZUg1Zi94ssJwQRq8rwkg0jLmQ3XABOoL
6CJfT2j+dXV3uzRpfoHClPo9FWktrDjSuBfW2ybIFqdyXf3pzsvNGLIeP4t9cpVN
bjfa9TGRU175y6MwI4FY2UCha2daKdbco+ZVHdw2gGLd09lzLMwthswu4eaAaSPY
DwaCbMGN3RNdzySmWThWsiQUckoKGa02HhyTA2gc9IpHTM6irNOGlPKrCwHrrA0N
tXqi+dAgRnX/bSwZzzbAJArvRQ3f1tDJY7Dqq3J/xCYUxLO9MdhjVMD/c4NaRwCy
YjmFjk1ORRukwZUprAu9L+5mzwSERwZgd0P3Gnp1RFUSlxImWZw2aIZhAowhQrsa
1TKESxyNC9S1K39mPXKxWa+zseYGIZeoKC8KABsXammTohGDZxsY6A1JIxVPE0e6
54fL90vqgNb5bwFxcDirv6eyKJauJjcOMLwGD5NjMaSuRZ4qIJtwgvB7b1nVvq5R
+OvFszfwN7hJIGUsP+23XJLA+eTp6P+n50OhZOzsHZFZpFLdbNNTT2ZRdM4wUclp
1IltMh+lQZ2He0GhqGNYLOpN4daI9U4SqtVKNvHkAStlNqp6AuZZIAfEevGrPaY8
kmX1Sp9K71LouDrTBX0xVmDpzdBT6+UpazKeVpG/qH36C8uiQLc+YdNqn4DKinSB
s6ZrevdDrksXP7lhHlIRW72s9XXVPM8by6onQ2AOM+mM9PJ3OimSfi/zGOx2mL/L
ARGdzXyd8qJ5bjr69oL5FPLFT81i09iusQLeCuHmcHDw5plIUYVcOBmNqI9RfjVJ
Ovgwrokl8Qsf27MX3f1uEUc0nT4WQQ6fnb0Df8Bsr/2YzBrJ+tFTGRWpnrbSZSS8
jIl9yTiDYl7QUrcuzOBers0o9TI5r0AoeO7vkPSRAqONEtTvev/NK6C7VneCPDxL
iqJi1mbe4Q+dSb0vnTRpRDyKljtdhYQ+VS2Q+bC5Qeu3O9Uss1ZxDyNXXL5o4Ill
C6TJP5GtkoWuTiWqGFeQHMy/Di7Hb7bHXoSiIXYOxofZu4nhqUMILVqdaefcjaYn
NrUiSlCq8U1B0CGfunkstE3sP0icy3krAC1AxxOA56mflTqfSCd2IFXA3NsKNEyK
qln9UEJ8nO7JNW/GbrC1tOSojd6csm5lUYQHeesnQrczoIP8cAv7cTcPnzDpwlwv
weRkPjP1C6wy6GGIIXnq65omief/7/U0Huv8hlYiMD0eNwNPI6UpY2oqbZD9y38J
gQU41wGlsbvWIe8iInW7/DxYpb2pQiR5kBRbWSYc2SrsDUvSPhQjBANL+nRqyuQw
m9RNLb0mlgL6AdX1lmfTH0SK7tZ2fXzvyQYsUtTBLV9o0yjsKwKJf54tV+TuTon9
xk1eSvMYn9EY11BcXnVizFYmlNnCZI6av4rqO8VpWJnL7nYHwRcUedStUJPzTIeQ
u0HJGNtoCT7DJQBKp9DtZgZpQ56/qYC/Ynp8OPrBzrnjG75JighpDAHT9IJKH97F
DtNlR6L8nJUyxeuZJpGeluePenANPJSc6E/YDs4ummxW/LgJVn30zkAr5Im0G8kN
pUOn2FF3JRHNq8simL78aH6es51iHp0OKxrXwdWOsylWcSRIm0WeCaZ60MBYSf2o
FYwaCXg6Vofu6DlEx4JVVNvOBAD4+HKTf0qMLe5WYcOvlsC1qhE+BweMKCfXBYt9
yZ+Wq0aLh+AbloO/dXYJNYnwHr6kjqxhm8ZDrg9k57sG0qz3dt8rGK4qWFUBGkx2
6VKIr9/3zecGx5yjmiva7TPhCa9Dc371iXHLcSq9O7D3dt0Ff5mhjAhaKrk+3xzC
DEKuwUJWIp++j953e3hTZqJJXEpbu9TUqltShI9rX9UApjNaRB1WjI33RLX6tbRU
kWc1PM2J/KTHq3aNGrFEodr3lmw68l+f4YE+U3OHtQDfLf20bjJScgbJ2i/kL3or
UtoANQleMHEk3H9DDvC05mpXu5JO796ixe4wNBePc8MRdutUiJv9HIhkMHh1QY8v
qPIbLV/mpVkhfdJ0ulU0Z7XOj7ru2d7YOUBhfMO6j/xJNYSP9YBy8c1ds5xgq8wl
8bali+g8nsUKoLwEd4H4zmHyaQmPDoESFDkPsP0q7LQxWmDYp9UMrsQbqMEQ4J/r
hfkVU9RUeVIXrfBBOLX25bm6DS8hJGDUTcpGkXEhZ90UWb2XlJt4syDSyIMIWhbV
IsVh5X8mAawWl+x864eEHhpm3+z3w+w3m9woXl8QW2OnR9iK1bTkUru1sdbEcsXl
S6LSNHLWvRELNebfujquvQpdtXogok4X8oy5gIYLvm4ldMcubE/Ff5ErfsNFehQT
EGW4vTOo7X30b9ctxrhw3usvMuRtDRcdJjOECmnLv7NqMKFTENvmpaCXk1y3bM/h
dKZUj/6Op5cydeU1UTO6pdDa1mWjg0oVxvgiLjxzJ0cOHT6NTZgXBlvLVjqYsZvp
j8zpp0N4SFuW7mON/4J9lP9jvVyKJ5SlTpt+JZ1JzBm6Rv4bUnkLzotFahg4B02a
ItSmEHG/xEmUJcmjPnn+t8SYU11ZSjfL9HJb4E44sHFCZ00zAS0Q8ryCmJ8fUYzG
EbQCGDP+xMFql9bUoIs8i+7sz+UcPEwJ1ODN6l9R8Kwx8v46e/RI3FIB1pq/ht6l
W3iBAAODePFp5C5cSRa+i6wiUpf7/696mOyCm2kFji5F+L0ADEEmNmvnQpN5Dnpa
oxZw6Nk4rRpqI5inuRo2ESFcFaIu2Xp98UVcTkW/oxz/T03rw50NJHdjbWCeNkXf
mGfst/2zmk3XCZakgTwfOJ+eCazPNt8dj8OcqhoYsFc7kc0tFv3+D9yvvTrpLGSP
j7J+1ToSHzo19g0dCCN/atRNZDuEwoJ9li755IWRND+Dq7GKoPsH9nyaxNZADucl
KoI6pJxuuDUlWAjUazN6s/TrnwGFHO6/ugzGcqTkOiQtmoGlIdTPJV6lDrTuVCe9
VjhOCN3oh78gBjh5CNH2w0eARqQKulLC2oYptyRrC/jMFUSKhSO67Z250jGtqkmi
iKC+0gLeliU98rwBdzS77pWH5A99LutnAQE6A+6GFw7jaTuWXNnavgIJJV3B5okX
Hs2ALgTiwJP7TWjAzXnZgdlbhBPkBVCnvr6VGH2FS5ekVPTNV2TViLkP5JP8YqRB
laPhcqs9kwT3VP2RTEoXYaTsQEU3MMFmJVycRAhEJPTK4KAf77rlRetgzb68LH/D
19Q7CAWJbcukWOe4J7KZ8zDJQVACJSJocUcobdrxDU9UGQ291HUgYTWvhZ/jFhnx
eg1JNVgp6x2VGQOPRa3+khbiH81z0XlT7t6LbpOjbdS0K0nyqG1t+i25l8DAgD/m
F+2ERSw8nN57231lVJRpRPeOLA+k+0jbtKtUCsi5mu2UAFfwOtZvTFg6+I2u1HFb
eziWt+Y/D4Z5PFFZtLvtBU6yyClt2YzfFAP0qhyOkVnrrapDKtElQzb6nEeD7l52
0HKqVZOs2gA9DAgViFyKMfyle4ly2vXN9vH47P6ndcM8pgc/A3BQfrVwlRLOBtOf
SqCTwHCmq39rNFJORKZIhOY+lpIV8pe6sT/Up2h9YUdWOPN45JR0oHdsEeNPjrVo
5l+7JSgKOuQ/iJteDztaO7/Pnik4+saF3waWTJP8j+5g7y9C5Nk5eFW1qrPpo6c7
nSYUN3x3lJEA7NFEE/fbCs5L/3QiJ8/CJteBtyHIf6C8gXaH8TZ6i660OSLQW/Ih
z158O+JXvIukSmlIZO/sir13cDtb34SZofeIpQ9jiOvXkS9KilzVwFzw+mdMTMis
RgLtXdvwQqkAfbrd2qZPTi359zOlV9eWelo9D8bRC60yWqgMlXo0gGk0sZ2+gERs
Cjpm5oIprFe4EkryDT5JaJZU7Sd6y7Wnp+imFkaPbfSpOWBPAuCNCKH6x99uKBv8
uHiFW/Vbc08BDiObLofSJF9pLMylMf/bbkmzSm3IGrMoyWf5D4RZYTxaXxKlrbrX
JMnbUwUq149j/H2T06dkTelP2cDXSZZSZpMedcO+ZsCUSHqdWTeiUOWa9N1kv+ZY
R6RCrXt4HSjcC4oNyG5YYQEfkHGM1RjpvP6umSnKkpj6mj9TqlKFT83DhrDk5gHd
FfLL2HK8JD0qeB2ut9IETjI5o3ONoijvgzXvqiKf5j+vSw2dFysKSCkHd+os1CfA
Mj7mN7LM4G6feCnYJb5GEmR3b9UdGUZlVKXNPg/041lxTXl2gO+gxMB2rMRPZom0
5P+ZWwbnNdV74CLD1LX9F1WzUglVqI1SeF0zY3pKyTn0MpkuzWp5Ywa3m5WZcHn0
o/O64LDqk2WTUYsP4uqrl9utQDkWRHFTZdleayiAOs3Gd5ci0eQe7/CNfbRuLrYa
wX4H+BYfXsQLROeiaSqKdANX5vwnZ6I7OxJoJJZSFFqmSmCmNAE6XRqNHFOGMN6K
BrX5dzo2A0+l97LqUBi/DlynqEUnIM/D67xo3/Iwu6PXD0vrkUJWMEw84s3L+S8f
QqEyqijjxemhlnXBLBjbUhVxmjgp6tqRqLmIdk8XpJ4V1opepR7A4Pa/mu5V/GVP
7U9GaY6OdzTHWYmCMVbAX7ewd5oBTAh5Zykhk0DMJlQ4iboGBBDe6S2RobOi57oL
2ejSM04LlOec76JE3r85U4d47qMD/pPD6xaudjSOliPwFvkLZFqhJKlzK0sZD7GH
fWh8UVoJeKII4NpqI/9KI4ioao9womDwwXSN8onsTx0WO+PQCpqtYG5szUSXlge9
CSOAhVtEbEldbncg4GKKbgPWi/f/hNe+PatXa+rzhZEEk9XL0PyzPkwH5nmgNTf6
D5Guu3k4z+v8w/itg1QXROcC57B/RDrKZMVqI+fIJ36xR1Smlche5yhsyA0X733d
0M27sm4FpcuxzCX/IBPjv6YW9arM+U2SZEaZXtEYc6b4V7WauSwMY+iG15ZIr1jG
8ta+BhZ0fTN30NFJnzeyaicaFi/nMNgewXHcKJBEdByLLhGeMIjxamcEV8hJCEO7
GlSw9ZW4mQm6e6lYbO91IXpudi6GSHFnXpjx0Ql/jWCBpD2om1gp/MJRQp1wK3fO
jQr8x7jywkYReAWOdoGX+QJkKs97MmTpx9axh3qLDybdTggUzm/sBFqq75Q3wGJH
V8DdCSa3uVBSfTrskPrJyHKH7Z/ZTg6jL24TFJo6oc1CpperNDNEl0hkIit6sDqo
Yq1ES7YAcdi+D9QawRSiuyknwPdatjMYnP+lJSwoUu9HCT+pxegjIj6Tt70CxKwr
LVhewQdl75KhIpabApVt9i9OjrdzjkIoS/IN024ROaiv9VdbxDUxW4/8X6w1tAUv
hnBT2KyYt4oGpOBSH6FzaODsKPs1cAJM3WVjpU+ydiz7Uno7ZUorn4nY5XB0jjuj
+lzynZ6VEQGdXOGYKLtBVss+Ya34czA9sBzcMNz7Tu9EtqkUxsK0oPxYJZVFVWMp
yH4J2b2WFS/oD1YmXSSjzkfukShah50iyQI6oNPgR2Ua9ZmyP/PovGzBHNvmuCQO
ihrQVA3iZ7SXMsC6tyg+slo/EaTvXhlNokExG8HpcsQJWvsYxHV4RhDl0gZL7/KZ
9LafHN0S/HbSR4XmF8NDP2SXCv0H+bNO1w2XusEJXS+fvUGg7dVp+M1nKbRv95PV
qMPjUyAcrOBNw5qG6jXFjzfCJrH6NEvY6sECTTDxHhwZAzGta+SBPoQ329VAJYLk
ySdUnvFD9PUj/ORzKhIBUitWT0oPMWJiSpOSODp+s4cH99TsdZ7d0I8HTXIhvFRR
uIBd/P1pfFeHYK7xWaQxU8K1/SDKQpT0IfviZ8q1wj0BqWNWizAzPxe1dSNoxFnR
VogL4KTvuX1a5tGD8QK2gZkWbXXusvOdapxd0199lwkbfE9/TwudRkXknSo4/83V
KUFuFKHFStX2uvSta1tkublfOQeniDp4RiDGogiILPHXdRrVtBg7cznTZz4KVNwa
k/Ih8FbPUXK/wnctP6L20B2BcqyVw2WqI2AresGHjSmvQse0rfLOxTWbI6SmoHr4
E6JtQC5QTkjG+/qZG+i08zcevo00JXeX3qMA/HoV8Eqp462LCdJqnEVQmWIUngIx
SY+CqoLnKiUPVLP9yr9cbIKWaunlNq736PPDftsWtTwahpwhuQRvd9k1JttHvWkW
MCMJwC6fV/0kX/1zeDd0LMQtCDz6ellXHZX1L2FYaic7pmkONJECd0uuEcoDJ6UG
vLlpuSEY5OqkFKHZknAUfCtBjFyhG+SIOydyPIJHPwPf6WTGYxfXZGEykY9Ujg2j
eFqDZb8ZWtFe6dnJLf2hU144tgq6s/mR/OzuIAJnkS4WAGbqyZUY1yi0wN5puwI7
+cyhSsJshENYpKKfLOt240yl3gjyKTmBzkaiRmD6TSjaAzJurX53wvCW+n861h0Q
hESeeWfj9raynaF3uI6031BSNtdBwbnWAK3surX+a7RMr2qkGfaHa8q13npi+Cxu
IOV0IMHY04e+/8lTUEXe7+IGaVLuAqHjF0NXuXhN53p//qd7/l22fq2s2j09EAMn
jnZM3vDTztFHRKA7/ZmxlB5gk7zNvgc3zRUoWUkLzQ7DydbFezRAeZEUP/+M5PCb
yaHesz+XTTXXxyMEGq5+/nAZM3/Job4PaHRALMaAmgv6p4PlmCKExHS5+895Iqts
OFTgjktvAbyjcnG/YvAXRm5/EjIkjsWnNRTrRyjSqNCVttTZiwRRHczCYQolS6D8
8xc+MSRgj3zWSnTzpjfq5CVpQnaPiwWoKhfNqwEaMWIQaUdEBlkVPTgRoZh0B+XY
t6BDaCErLBDd84H4tWlZanpCgj5gn79P9aO7yeCOQRb/0htxCQg+OcybgbVXdqqz
N06V2qrrZhPvYOuMmC/Di4ow9GQaeE47Jf7VdUU4q5FtbJcoa9RPgsusAIfURFEn
9U20FcZVJkOX6BG+fEyBcZAum1a/JjmjXUXvkiY+5DNDoYZabqhsvJQz4d+i0+re
23Kqh0PFTOysKmVbpwGQXCqjpdBb33Ni61lAbuWjScrR33I4Su/5dFKjY+ycmADJ
1oF8HtquGagGOa8iW5E030qiIop/rvBY04kGQob5CL0NsFkI9/zgBKLzBdx7cIGg
iqMM8z/JaaM+B8YUTDHisfEOLiA+vlxbgPAjPn9p3pyYRJ6vq9bu6EUwFBwz3zcK
49E9jvMsWUZ2BKwdcIEgxPcF8WRmiteHD8gE4adNnJ9dnDIsZkS/dtW6kFx86FgA
yrT3oPbg+y6XK/1oDfrJNS1lj/OZB85Bks7rzljhijJYaszbVUmPMpoy9dKOEG0A
AHRbA/gDobFEWRMkdNXZzBawG43zWF0aygsA3v7V9iudAD8cVnbeyfRbfzwUPT9i
EZNy162TOuTnHtLP81pDf6CaDDVeoxuGpiXuNfGZX32BwjRqlZSSEzqzOZQ2wQXJ
O6uSwGqzSjOJUVvXzSY4yXTtEJ3LsWQCYSiJ4ZtdkAIiTlxSM4I8oD1nQ/tYoUiH
PCezIxJ5t38oZpDvnFqiCSx8ALSTabuSsXiVUzB95qmOBSQeT1XHdmzupBBoaAM4
CBios/M0VFTH4TdJ43GGQDBNDOude677N5jeewhLqhJ3ewrriAQJMXQvqJK4Owzy
E1lXDm8SJxvGX9cygYOqQe37yfPvYjKyNAaWBnylTkdOYgZOicXUYBMTzHsYHWZA
rOoZBX5/z8qE/G7QIjCF+cnfTwh164CjrbcVd3/4cJ4pvozZJgDvrrQnipUuNPmP
6nfVVQ4wTGSAH7dnpnn8mihj7Dh+OchoNPLVYKw2TcPj2UPtXN/QMslUS25H9ZIR
DyyKik0uYDN4vOZwmcnlF/0CKRH8WUzrAMFl5mAScItG6DN6kCTaa/sexIpN7out
3AzKKOVuvv7T0DDYYhllzsSwxguTALRjltya0tuTDG6jtNXpb9UOS77NYeENHnqT
nxmWUT5RTMSAIh5tsyZp6ixBkINicpKlRurMQJ3IP8BnNQS422PvIciY7fRI/7Sw
J0ZfLqrfpq5D31yH9Zq9U5o6ezEnZApsc3ivnr5TimlJGz6djpx2975wquEZV+eo
yVOcjo86iBNAHQ09OOszjyIIqGd24gt02KVat+mnyKsv/T6IcTPFpecKNzQ+hbNc
M2t5Q52z4J+6YB9xJbhaDQ9MQrOxk+gC0BQ2YzGpw2BZp86/vIRXkjg5h8qRN2mb
+SqMFf8paLy0dem8R6taYY3UxuQPyF7PTiTuNIb+YaPP/4YFboAdkE4NB8CFHG+4
LaBgMaa2kiOf7AHy6IETUZ/YybSUe9mL7FyXpeofkBKYzXUOFJMt7LmUjDzjS9OJ
F8lyHlH2WqiPiOuOdz8tnbvBPCKP2BbzpKxLdqPo3cfTk27N0YyDsWznoVJA6Kjy
HVJ9oUgZXOK36AOfycT0E8yk7MXG+j0gcHyix1bLOa4mF06RZrSy9LgkShKceClm
Mblrl4Zg/9mTtQwTYWyDnV85NSvOVkkeMpeF2x9THSE0U+xfLgrPf8mtEB5E2Jy3
sxFNGD+NKBjuaDh5yMUYQCWbDlW1CIFIN2PWFIrfVRHg8dwGO3KCbtwFfwiZeNcx
eiIEnga58H1/1TbWSp6Ml63c+CXIP/aiDkD726W+U3rVrq+kCZFxroIcBOs1tOzZ
jDih2CROKYZ++65kvGk3z/eC8o+H3ZbvMYhEHXPiXm6v2xOaVCsdYAmLi9otqwcc
0gtguhO1SiVyUj9I6Cm+jGLbpBEjRZtmuOAc8YMeYBDl7hCYV2LhSN3tPpoGpUwN
+33hU+SotoNb2MJN/N/XW+L6K3Dcds2t+CdHZNf85Y1DoDwMEaTrprukQw3IOBgi
uvIlsR/jaoq+vxHM8AU0MBilq8xdUtcQGFrxpcxGH7Hbx8+/zwTCM+ehP3ygRpTk
KHY+SkPnlHtWOMxbKd5aQWGzVA1YdVoFFKMx6XTjWLL5Y6RlWx36FG7bpM0aCixL
7x9yMrUB8/TMyf2HbC4N7iSq/KFyESHoepIV+v4qg6Prp8wRbpbVdObf1apzlhoY
U5uPeN5+SHympJ/9qz7hw2Tm5xvbhxwJyXVCGIH85u4hBLcfVuXRnVKiNGw6WUgr
JEWp8kuwjKwBNwQdf165yxLBVTYPesdgRhkq6nqNwRJUmOmu0JmMxXvNAzjudkb/
0vM4Y5bZ+4IJDoj0Aa9Z9l/Q1hHRv56XOADkObat9x10h6+1uRYexbuDCO6dmlNa
SCwSKsC6DgVDzz3giMB6RebrfFp5Pq8Lneg886PIh8KXYpbw7UCU3mch94luCG5v
og0t/4XL9A2biiuwPdCA2GWy7sARvg1Fc6oM6eM4zr9oiKctx1Rq8z+wmI+o3efF
qncOIQY46+UtCd7IXr8IpcgXFyZ3unx1i7Y4iawiMWE61TBW5nMod4SYTbvPb/0B
pz69xqPpbD+i8mYILPXlssMP7a/bT6UB+Ty8RjXSrTF8Y6/Rn8kGblaBntgx0mIR
hAFm5kh47O6fTHI6mg+nZrdh99MBSK9pdyjxst0EDtQTn3GoXURGhW9gz5XHkrvY
rCs4+w+QpyU/Rg/Qr/lklDwObwLRUf5aM/mA4Xn0tDOu0hYoMiTPiN1Q9AqQRBdz
49nD0Ie7FGuq+q0cpQ0OoiOfI7JCqUZ9rHFk8ncqRjhTDF0pTZnpe14ufeQxZSq/
r3LCvAL2jOIj7swTZVK3vs1RXI5JbQTHkERkG+l6EhOX9Mo5rgztlBRK12AYtImZ
Hj7PgIaNgOGzwAqaNnHiEvoiv98JPNUUjkDDgGyxX9UIdhM31cOMeUjoaNob3sxi
yfghpZcrIHAi+YLTpkglYEKjdu0qf7Z3OuIo2fwCr7qaUNSjOkH4U+sbQpgy894M
aZxF0Vux+uaHtzd2hTLXUEjAoOJOmWB/WOB+bv7k1i8OsOJQizq/AxbDgMXMv1PU
ilj1/mP22vFanrneuSQ/KbsfgkW39I/9iIc9+t+RBwPlNUqnzrVu9jj2T+UuhiNg
Slzhjh8LF1HbzBPba21ld3EYHV0CJqavJdx1gITcUlVSnOxWJux2cqx4Ua+Z9c2F
qDn7hkcuRXU1CfsNAb/XLO2oaujdYK9mt0lcPih2J/RtFfH76FlU3kXC5Dy8SRTP
eeJJZulFExiG3uYZ2rI1ukTLJOCRrrWTVRRre9wmYJ2PEdzg8x00z77A9M+KkxzA
KAP1pO9P3SgSx802xNoyaWl/iE6b4TPMgjtrUMExY5jmdgq947NJseQzoevrJj/G
7GQfdjcuLBpvdmUUzIfkSuPpFXc6pInQ6W11rDZiQyxT6JCEyXF8csJ97dcFtEW2
hcqWvC9SKMwpLnzR9LAXt57e6ylRbnd6ENOvbaPrXCfv0Bgy2TehLJeFlwUq8WXe
0A1IEGa2W2EVFPOhKW48BMTsD/1IskXt7kIRVgrSd4eziPDNDmPBeWhE7QG2M8XR
gjuJnV7qxIPoR/VC4FdgT0E0Il2sAkfLummI4vN1dYpU+2qlRE4xrMXtAfT/aFyv
p/lxVFKZUaOdTFiDEzSrkGQXMHSj+MppvOpotYgyDtvt69lF3pjnFSAo+Uh+Omx/
yTaQMKrdL/59CfeP3RVTidW+eI8Hy3PSwR7dk9PT8YXLPJOiVaiMAepcWakwmMs8
HNSYPmw6DKeDthbcWKQs7oymjYp+KJxh3szuxHD5UPyyZJU74AfQ2UK+DzQpz/cd
4ERF8upt8Rj+LjnPCjlQGF5Ojxa2Ac9N7vEftlqf5AzvSfma+5dX2vC2vP1B4zWr
6t8cfCpbDukGSu7oOD34MhxFbpZm2x0JrKFJcNGNjLYkcY6+J0LqO6Xu+iZgyRcE
IfR7YbYn2bgtJ+dLnzzxmFBqq7BbGS7G86Hc4b2wize1cnud19PzZYGKUlYrZv0u
mK41mOMCnUb9DbOOCq93gC1D2sSEfadNg66VppXqajtcZXOFVjLAfc/qs3KISHoU
ajneVgdRIbWY2dkR9lMCGcq9Q6gQDqYJNvr4IMUUMO1w13EBQgzBBf0Pjm3m8xZu
/uQr81CuMCnbZxJ9I+gdUPAmGrqg2MrRYTy9RYFAaXuV3p8rYv390+jyU1UY4o5/
11WqdAcTYbZhYIJZyJQicEIr2Ja8oO22xQhklX5fGwJpCR+ugfPJg0TJ2lV3WGCf
dxJPjzYCiPZfSLAn2waMIjyd1rRPenBJOwdy4CvmFNj8go1XR6mGmt1665GqNLNy
aC8XzAf6kOoGqqz3IZz11tijeZOFuxNQmax+JiYVpyqyL5X5Q1brPfyF8pWlUe5b
i567N+BAZ8Ae0mfweWnH0lqR6j/gLdxdGB1SreIFjsnAcz/lrsjE/YIHpvTniu9T
H/HbuHAbKON2gA9JYSQ8zHzmkCgpTeWQN+5I1tR+jRtGqp2HmpD/tmzrljVJ2Bk0
tRZ6mOjx6XS9OfD4GaoMBUplOKrb+PKXuUUMqs8iHBspBNQNHjPF8aalydAeVF0c
nxmdMBOUNGfAOdMe6UXI/6zhuaBys02blvOVKKK3ZPPaXKC9Ye3oRT5DE1iTVYXK
dLD0d4wf8Kxy24Lj+Bm+7oVslU2jlkFnTS/SmiMz62QKnJhhUPxx5OfN9M1TpwIc
D/TZ2cyQqRtCl3Sps/h9n/h52VpAGQ8NaRk4S+drBmBsw3WiSCdE/3Fua+CCQiCP
v8XmVeUw0w21+UqQq6H+nwLX5w2Ulfl+a2dPZUepHoV4mYtIO4daaM7Sho8O2C9F
jSO/iVieC7EO04bKIrY26ZIhrM4rFWHcCcjTgR2ppuXU59aOE5L308xcixj3/XMq
Jme4b094+39Kzu2aBRONzWkFE252zCK+0wth7zZpGKzua5Crm11oVxakIMxAFYqI
/X5fhZBeXYkQumzvNKcUXhOXgpAg05M3k5KZ8SeBffwxSeAhq2ft/GcVV3d4XXYG
SSSrNsYD9/U7sE70tzl4777E+/EZKEvTc/SsLvnauLrX+oWEHqekmGU386Plz3UJ
Ejp2wyb3llxN5/JDr0FiXWRGodDk/qEJPT5SoAAJSiwA5h3AsGYHOtWGIQVh4iw6
ALewkejMql3ZfcOPThgepfr+3Zm7ugE6UAb32neDr7eiv7vXsPccghb3iCla3oKV
iubqdYT8q1uAuBDlzCFh+EnsdUk7XwNXF7zT9GqyRKs5cZxzqbAc5/3uI6mnPVY8
UcMViGFXmpxz2IzLzuz6IetSgjMuXEEhOD4C4V/+NN1ndgZqTBjbdTFv9qFIUusQ
s1LXHAnTTWhGhOtUTA+OPTlpSodlCGUaqmFhQq44QT2xNPbtypvUPLoFer8xfr2Y
8BM6QCzkx2F1QJYbcTGKRxaCiZzZ8rx2n+RJEcCdXTY8cN0Ux9nMBg2ZKz87mV/q
8WUDtI+H+2boWquLLSFJe3e3ZIO5z5KsIoS/liJetXdY3lT7ZjDeQQndmNpq1Lfe
Eq+tEUkNVWawMBvuq3gfRRL+YRUj/jmLEYd8uBdpKOM//m3ccy4f0+DWUarU8OVO
RFPrk59xGaEYktT35SLQIDRzd/4virpTFOvDQtBiXL+ht3WCUyvxgm47u4/toFkM
gYphlEjkHOpcbz/w/t9YkSw6+Rqkc2ova1dXy2YAflLmTPLePRRZ7iZUXxut6heP
j78REjx4Su6vbXmvAxToJ+dAfaXbKLHHu2rEoTRuIFozsDg/6RKJmlhwm1PRHF6u
uZ8hPxbJ4rNu0IJHNisBWLY67LvdYZ5P2cLHVEnG273dkG+JuU3/cEqMUDsTu7OE
EnLMlV/Q26uaQMCNbJq93vop8eFj6oZ2ObsZDPDeU1nyFVV36veCOLlPGLSq59JG
nsLdf3NDNvXC7ICUQdJNSfyKA71WG20j/TALmxTJ9JSDbuRcevxLGQSQa3/OQFjH
VHXx4PbjPaZYKKoNK5nN1+kdSCXivdo+L+QdLkQqDMAZNakDS7wvPqCJlGvWiuap
vJ+LdPYSC/uA5WcOZ8pJwOAYRtbB+yJCo3xR0YED5wzOnaLJDkHGlMl+Xy4gXsrv
6mfKYhfaTFDA+dWzZDlHYSYbkvk5/KIlhz+dKtNklHPB7So5LfzKdm/Bm54uF+yl
ZAvomnULsE+qo47lVuQuEvkVZLhcsb+G0EH+oSjRxgQ7y56427luADG3p/RC7jQC
Y380ZBDBm6zzo0wN31862M+2H7jGHVEOT1YbSB7n6KSmcJRLODbu1XQBmfiouxPy
y2EFM8RDDevHniZIPU7+zJSdzqZrT2mWIpzvlEWocVNyPRdMlsFKaOCKvLGEyLFb
Qkrq89yVpwMZ5oj7MEiJggHRDCiomUrES2IuCW2ks9nyXPRigeclAVyyJ59YrKV7
oykGOoNAIVMbQdpHze2j4cL5HXpmYmql976mT5U9+PIdUiP3ZT9o7Eex5s05NQ82
48/eQv1kvcoJHB81XEx8aCH2VQjfPFB6tJkqW/RMoJw5NQMEj9OXcXgSCosttMwa
9cSQioaEF0fx/B9uhJt1MAKfDaoTcazb43NmMXwi3xXokPvfAWdcDSz0B/Io9FII
LkN43iwcrllKX4HpemNk72wgR+Y82iMnKfB4gBi+EdvL69KzbLnJO8jTsl/UzPum
IyzK76IRvJ90yijgJOhZ62uP7efrTEYbMyUSnGddzFZ18IpJss+RaVuNAMkeeMhE
Dq+eNOIFIJ0HIwDzB3rCMGIz36/gaMP6tKVxdUXyZRvZZ8/jaJC6EdVhfxMvRm2j
ifz1yibWKJ6TeaeH2Y1NEOLqCigDWF/W9P4EMM3apUChpTM9d+a/royEG/1GQa3g
QKJPS0lC1zGmEpjCjV5d7W/QjlwbKTUu+Tg55MMX5xTazfM1iazXEr4yErLOB9Al
yyV1naLLF9TQiqasEnCJ1TkA7BivnU2Sg32qBZwbSYWXfRfRCV+rz6GZiruhwh7w
Qz58EXopP04xFcYzqYxUx/5mf4BLhHLUkQL6CXwTTdl9mJQVBlozM3Wq/n468hKR
TJSd09gZQnHWea7wNaps3QS5UWHtnKsPrfLOKQ+DAU9ol/2wr2yzRDDg7p1bnSTV
P8iQmC1eLhpZuTMeylpflF7jdkWUoXeSwxFJ+pwKYCOI7LYXmcL8O3sxZ2YfRuOv
VqOOLIbrzC3r7kDyJrgmAof2NcWD/MGyT9/xNWlhDTMRiJxSq6IsKRu+jRKXgP6e
R0lMmUXGWcw2v+0n25pL67lBexuSIXjdbWCLbpVenzFLmYCVLkHaWH47ZQBas9ef
DbllzzmKyGMD6MEwbZixW43NNayIhQBsrMI7O67wjY5R5WfDs+jfdVyVlFLk41US
Mmwz/LfAuj9c9GyWsdY5RnNz7eoNJYCGbH4W73Mh+jqsXTE2CjH4xh+rP3d8nS94
fUyeOs2ORolTO/KJAhpuZhbt8tSL3oA2KRlDwXFoGa1S4GB1v7+D6s3lSnNvxKGw
c8RFgnR8FCRRUTiHyNGrJOnphHYQcVAuCHpt9+xaHff3hZRjc0BOB+mhtiTebyT1
YFiLzfYhZfP/wWHRt7UqGLm3AmlM1qe1TtmiQqgCymp1Hq4/6q0jDtpeHcQbOto5
cSHtDu5KXNEDsFh9c3UMeNFRChcTnLTb7xp8ZnwHlTRmxftUvjcX2buuSNvXvI18
UBubjmNkpDN/kvsPgolOokv62cIe1foC1BtJPcPQIXkO4afMNEZr5PrmGACbsajn
n8YlgwA9wMZ5/dGlU+pxvOm5wGcgMDeSnICRZIcq+jKzn+zarOT4ODvCqJQTaKDO
lJ0oui880Z5pxxfB82s/yst5tmGFbYAAvhDOEipTXTv66zlHgmwFd648POlO5q7X
OoPSmaxU4inGZdUg2Zhmprm9b/k039Z3LrWJMnLS6a+FLs8NZ8oXS+ZZfOUCqZDP
4dlNsAb2yeDR4c51vVKVOcqeWcpZOVXuKsStn2PFjBhlgz7ZsX2qgmAqkCHzAE7k
RNJo1q3ylO0T2/ApYqQHOAq7lPar65jdwphncsxUvswf+IAT+ZqKBER9b3ucJOK/
mJq9v3urZWO5IaByfP+wVkALrbklAb6ZlGL982g99D83fsC3fC57EnNtqVeiuG3Q
8WrkY3PtIZV57s2OS5bk6NpTJ1MhWTYPOMfIKa1CLrHI41VAPb5J+BBt3vohV4+3
0TlvHc0XDL3Xw4YQBsER8sOK4Y1h3AuiHaHDByHraM8htgwVokPiz2Trd0X514vv
6dehMawKMQI/x8DLavxvcFavc5ETTWEnEpk+ZSOAlyDmZCkycaePYbn8FxerpkU9
jEMSuo79DcBTC3ePu8miLC7PdIHHPhvEbVpUi3ZDhHkA6McAJ6G5zKo+KxAIDXww
qp9kzaT0DkcG61/ke7UqO45XVnSij5B13G1ynL+dpdxqVVB15vDPCobwGzhAAXUm
+hq3ZftBq77qgxmpyUrOxx3ecoPwuE29qudn+h6+Y4Mhtt4gL3ssP1Gs/tS5acoL
5dwwxETxRSiMoNUo8lYocda+pdaE2Kxm8uOh2qElamFWpSy8jS0jv3YE9h1mMtDH
oMYYBcRUZ5DWPKuKBG7LA8h0iD+1mInrb2IOA+/rmA+iMunqnweeDNVdyHO8dnYD
4PDdbyI9u6dpdUq4b7Yzjb00ldYrSGRGHrlMv24Ni9yUPP+3Oro/EkH/sqOJdRkQ
J+vSh2BqrOxUP66mEeSkN8yQUQaKivGZQ4hNY5mCVR3CKr3sy7CMn6+EqmYCPFTu
Vnc3X2JgUC6QiP4XSROJWnRG2NFDBnAObPrHTS7YzUbxWHMQTqUCZ/+lMnSXp1v7
vW4HQX+HofdPGzehF5z4srqs3N4L5ivKEbEdPyvo4b+vMW6m75oNQnHq9e8omLHK
AWa8loWPlm3Qj5o88e3KqtsuOA1yakDnZfNB1amVz6KbC47HRvac1nP5QrpDm/5m
p+fQokNzb9uT9pD2sGFQp7v7QMFD5tgc7qaPxgfXs9TRsEfc0nSIrzziIHMF+lXL
eq2QESK7JIfa90xuO2qxWg3Vb20j99wklLZj0McTn5Z/gKc71JYLAOkfI0MUvMPP
g2O7gcOt7yv0kljrqbppWIC0LQ6HICqwE1EsMGp7fugF9Zdpj51trAVL4YheXEOj
s5ywDrGN4XkAVUwCp9gTmiIfrNXkSNQyGwr1/2XzbAfMXBKoYEIExy7a6ep+rDo9
baaTGSQInJhGz+mtnG4YGsK0BLOeWfMXagcm6JJ52oAknPk2RLXL+/TSmYaldTFl
sbxDAL2Do4hr3oc6h+wQ1Ez8x/9vL2H0mvL6GexOZ+XxrmnaUMIzLylZmOBBIEo9
ZLsRH3/ZBJcezrXyQWsnh7JwuZPRaK/H91ZaKBB5hj2/OB48sO0z6ZeDYXE7Funm
DIzaeLBZVWdluNXyOggfdte0qXkJqCL2aJNLLQuvHZnQQhlPIv/MUP/ujE+eS5sp
/cRHnNHpH3ZdCAoyyKI/vlRESOiP1cbK/tP3tbaI+rpRUeVMRPw3H7Pcr+qlg/9h
paffO75ru/rZV9ChtIXAybgafWwEKx6UKvw6IDEDDzhTmT2Jegu6374BY1PrL5OW
T8LLCgzgvaOcWj/VxBzigXjVCIsO/JiSG80HrU1PnpGL24U9OBlREUBXboQmtLeo
3hKoxYIfLr/pN6HmGbcWqO2yYJWmBiFWG2II27mZ/C62SZYTvxunXypDx1+2ycE1
incyxz5t3jGlcNtvWb2cFlWkuGHBLin17FS8ml6OjI5x4h5/KL6yzcfR4JQDdhVo
XaLMeKOUsrcNxhlAPtuLm7+QAltWIeXhJ1b0sfkXy3qz5Y3aDmeNKCCyZdpnSoaG
jtJ6clOTb0NdwK1H/4g3fV+f1COMjHxQPIMR7+dj3gaCsDn6+tvCdePmQofo6ohv
K6skO9Ek22+r660wq90JSWMk8PgOFQ6RXbfQWcD92DcxTdL92lR0UmgS1QLVt7uH
yQzUM9dW3+CcQmWijfblFJ3IznqtCQnc2loldRH5F8RGHnK7EbXTA9ZUWLZ433nG
t8/Nn75psKnGIKH3UDDB07Dj5COCAGpbkGW+bll9NhVxMfqbT6QzKGy145v3J66b
GjcscCCnTzxXHyz2Krtdl4dIOvsLil438D7MWVWb9NAFDEZc53H0uPh0g59dRgYI
CsMs1zDPBL5dGiwK0TlMkLuKcnzlFPnLoB3pNpFroEqPvsut4A4gYnbep4V3enGl
NZEFJynwP7UAvhO5IhoQNnuZxxlDMbJvE/GRnWfeK7aRPIOyhjdY0TLvw3/R6nmH
uj9uVlOTCU/9mK7s5Xie00pPHfRa3Da4r4yt9ZyaAKMwkSgWRyGBa13mph6wqz4h
HRpvqHyvqcYpla8If8VumqbkyD8Q3oVKvMhhH7mCpz/8aPrpXny2mfQDQOuJBgBY
PVMv8Ond8ez236+eFDodnFn4G0NMq5Gobqd5zJxBNyG/YMdYKTb9aviCFVvMWv/f
uVGrPAMlDrap+xvvWdedICaE+dAH5uo1yGLjy0npnrIzv9JCy8Ei8Bh8ErDSEOkl
5M/TmT3IFYxOe4+GloMQ3/q0d7rgoxCgKp4VjZ0hKCN/zZ46F4KscRpKAnB8lMdQ
Ah2EV5X1YgNC/WlQucUwV3loWDElGhUGRB5wxCBUYae7hqe/8cGOu4liHobussCk
3zUmnk020C42ygbYtJXNlSUGGCEybK3gD5S2hR2p04KohkNH/PaZTZi72bzyodmT
d/jb3qg9q4iD4E2fF0vlh1gZ7MrpzD3+pYnv8CeHc+lAjbl09OnvCEXihHxcuXV9
eiE++DtayzrPBRDu164kPgtZSGrZ6U1uwjedVanhB/f2RXC5WfbRX0lCIL5otRQh
VfvCY8PMPlSiUR/ondppt/s/AFxNjIMeLgDSZxUN3riBmZNlxPwE/lh38Bn2hwe4
QCIWnlQd6mDIV9i5nk1qYTcdrNMJgZvxxC9uu/4xU0r5LQarim8N85eSax4h81rh
pvDUKM3mWUyhkjfY4HO12eKDWVFmkI9fL2PKaR5v8MJXzmtbnhkRJx7lrKtlazX0
yCvI0QFrVO2QypwMZIYI9R/uVCq19efNCrb7+JAtWnM7gADVFgzOpKT04zWMNt9b
zhLjRsDoU+HhXFru9mufotubbtlAcVRcEkw1+IQaU5HpvDPf+hidcT2DaUJItFLC
frVGUg/SaRChgSRytvPgSvxzZ6k/fG/Pwz8OlpML/pgKllswyM4y/HXHFUXxAJtJ
T0j6ZdSPYV+3HsN3I1/gt1tsOFpNeIeQeK6I/EMlY3c+bGXl7v0YmatR+UpbM07Q
9LSYWsZ0OwIkmYTbke/fO3mLjxBieCsDNlOPuLnLuH/XQRy2ANGAFXp4tYVgqyjJ
InAV0pEklrRdSv+WEqVaMEqcQmcLuwpAX4ky2cQ94tF5sO5mytboJftqPx7rGeI8
fevrhFnVh2CDXjXMlLt+ckXllnewiMaBSuRRHstO9CDKoYdXBZ/hDMRGHUpU+pZl
3RB2CviBHV+pYzN2mRgEKTXpJS638W3Ct36+x5DXAEDDNqv7FuEEvvFhw3muIwRs
UJIvt6U1EjQu3FBs2PdDeY5u/5d+Ysj63EBzRNw0Al1HEFrFVEW7C2VH+H3dYc3/
O5TFKccYyaM+MMnkBx10d/vMELvb+2s/z1wbyhcPgCdhGPknumxyWpM/O+YF1KJ4
6zQEpQ4qo6mAQWWIz46rxDNiD1GDEf+R3aH04byKEgA5tvY/apKm2xNj0EOaAgQy
JBoARpTP1lk09P2lTwHKA+a0tK2bgL+FqxlELAHFGPbMEa7grUZ89VtN+vj5x5Cw
pUSDKKOKjrhltUzwH4mdRnzvB9VnaZ2Akp3icERlM77are/1qkt2IIuu/IPGRg24
NRx1vD7oi12/3i9JAfQAu6tvQgDFNvur+HdQNaDDyxvWOAO+AcXmHrAWPS4o1WSb
yv6C/bzMKbBo0+eUD4jNix5NcfPGmxTPs4byomDgYVPm2l90aa3OxCtwmHhIjjSq
FEa35/L4yUxJp/gG69EODAg1EQgRyJcDt5kYZsZHu9Hsb4opfmjVRLpTyJ0VFy04
MuPlOg8HChLbvXvnVkDE6g4TjQTQNeNjnPWpFJpbaYXNS+s2Q09OjtFrAJW7XiDC
MFdqqHMLLvH5e/wS32YLiokdI/Wnq6o9y42+/ozRbwAL92FWm+AQ7SzuLtS8acYC
zmufp6mBe99VwyKH5GOW+k1EFey0e4xHAzuaVXZOQezLT7451s8HatewA0MMBAhA
iSPSj1S2QUud//tPDP9Si+dFN6kpKIVEW4duiBQvFpHeFLX2AwmHKscXy0q7HROS
iGPcjxiNRRO1zjWt9bU5Z5UwrkWzZEKjTcpghXgQ/FwN51Hhz/O1DScIqjfvdvHa
7S40Rnv+COs8HVytpNH3MN7ir9y8YZAWuqwAOVMHI5Y2avDum5gh0MWet5lIALvr
X8ZFefwIcKpEBq5iwNkkO9ORULAxQPs8JE2oerSW1KM+jGPcWa+rlsjBLsoUVzRI
sG8dxSEMdhqdOwLnxBbUlvzKwP9Z+9gMFvVcrHcuL1u5/YxLbM4pkl8pBAWFfErV
6VPml+yovmDkYJxRb5/Jl6qqR0kWexWTcEvh7k5NGAw8Jt8uJiwjCb5ak1HaLpoT
QzX8NyzJU2FWPoE0b9TCaYq8fD/ZzOJ4VgG2uL++AAcS7g4rPJHjFiw9dsWhUuqj
WFaO4yrupm2FiVoWdPfF7j62Sjeu4t1wXJCc7I1OJ2dpKYqh8owiyCNhRzFYBNBa
RjMkUapAyJpWkA5wZHl4ZMIcMwidz8XeN1by7yAiMsliljCyykIDxorotkxal+wp
5o+1C9lEijSHOwZa0/Hv402Xto0TyJcrD7Q4m2Qm8ArAoEOA6vs9agEZKbi6P6cp
imoxzNx6DPCdeF8a+Bdx99FRMpCPwgxGcR3oxpm+DSFhI9SJMknoyBNkxfWSaTht
TGiyv4oMtB2VT6hn7oimdB6tmygv47/a+0SDXsvq3SDot69klrsxLFte2hwQmyWV
vXNzTeCAK499+2TnctyYJUEM7scUrVUCTeu45ViwBTkBu7KVR9Hm0uCYt4RaNS0p
Y59YumFLrltZB2RjAQB4M9taK0cyHpqylSFE5Yehpy8WxpqwsW2YKdhxAYN3KMBu
iVCRZWb/XWxhC5btk5OxM+0apcMrRtuGel9t85+XjhfFJ3snEcMQRYaR2smcpS7k
7Mt+e/XOtBd6pr7s8sRzb/md+OQtqNUsTb8is36wTWivtBJ8ErYaziQt+6bVLsH0
UNU8jzK6MEB2ubtSZfuDyROkabGzaRH2J+93ToRGieAyUhII02VkRDv3ktXI4sfA
YRYKclyHcv59RIDdOD9DpyBk85Y1mMQgsdbq2oomD/DUeLnNmUcMDLeTv+2UbbKA
1xgpdX4i5MxTuNWBeMUHUiFBKfYJvrF/xYoj2iuKz/rDATmef0AKaEWftzjvMCbA
8qaWDe6VZRCklYrAOrxYZuS5T19lnxHp1eC6f4CsyJA4ZbyXTL/3MY9WrAx2szjz
Nz/1Ic7/0yuyVLOYorlm3wPc05VF/+oJnFaBRl47vkZ/lJOCH88VXeYktqyQ4jEv
4oNwh/ZECdX4uR92j2Lx0ONy12578H5FVjqbdXZCvOGo+t+W47DK0vl4zLSKwi1X
PG/q9lWbM+MFbsgyJB4546EYw8KvZStscLwnxmDmvt0ePtwEHJvxLdPgh3dQ2pMg
Ky3bDk27oeI61dlOp8M+RS55HpJDqKfNss3IzJMD6YT27NBv387HLVI+nyT6BkvC
9lVfal8B7mIsDWbB69EFZiD1huh3Fc/GGnd4sQ272dPwaivBmQ4Gbxh95I749Qi6
zDQcyM8YF9n+TNdMeNLKBEWd5UzijQROWDIFAkzgP97aoOSQUfg/ABuNb5dVA0R4
d1q9PZLzX3eE0MZ6+nyigmzrTNIStNxlHZ8bnJIGhfBOevZI/IFbYIUDCseFoQgQ
PNEWYLyRcVUaFOgts/e/4SYP3dTZtYLvl6TL+6vLyCsbjd6B9oeB4tdJmkK7aQtV
Tl6eDLGZtStAAXdOZlASVi6vqn6YEtPvTe5wHMocH1sG5vXkzfD7n+/wvDfSz6YH
ckQBcRPWUenm9cvuvPGj21gy10psZt077dspGnX9HdZxSi2FfiXTIAgW3akD1I/V
B11PcIPYhTno4nUOmPpx4luvhUG2aM4h5TDhJi1yeORYln/vLjWS8RzzYdzEruCU
LhvohzBktBpMOLMjooCk6O/VzBj/PSor/1b+gsgNeX2mKq317QOLFbZsIgj5qUep
hwrla0hAswiIbiGk65wLPDCFd5EGzBGtQNIieABat9T331dox19pkWjHwGnLOaoz
gw7I08pYhS/QThDyxLUU1ZKgVmMC7d+qrhBSXeXNwhAT5xSO2URlzxKH3f6PicYK
92q9TOSWq+YT6x5e3g/ZuZZOCevft7oLTUrg+zshIBQPbzXru8qezglvXfacFBcA
gfLfCoJDm1v5snUV5USiXqjciB2AB3lV7yyX2uCrEFuH+4NpO+fuXN2pg3HdqDK3
BNZBUbuwP0uo6ta+wkZlSezQ4Arn3NLTRxVWFiB4RCgMtrYa9bbsdVeifclDMruC
CaLKxjvXTum0cJJPXwNHIxSRw+SdvcsaZT18zrpBU50DWVEC2SyfXCzQj/JXKPqB
GDr8EhkerAG4k8/2C2a8qjVsdPumS27pj86mWV+hqQgqeAHDDcCob0H3fNcm2XZ8
ge9GLbFG17EaSaBpF8d2csbVLXE1reFrHm+wfpJ5/6t5aBbMTbCSQyjWr2CQfQKS
t+SRsZc5vgwy7amZ5pc1NcH0XPME7LbI+FTwVQRrZ6yfjzQ6op24n/8YSjQgWIM+
sD1I/NuJ1kYqF7JBuCvgmwAG0xj0TKUFCQfww2ePl3lbQTKrhhhHPDyv5J4hcUaa
Vt69ALFc9AlHwv5oiE7CcqQfZux58AxuOSMY4fVeUA5agdCZwhV0SKGMpQ7q+HZd
s7diyCBA1Cm+M+lJy76/BmknBDbh/uDDNlRXvPWq6tHbsFH+2L9waColIKE5iGnY
15lQLxVscVlAWkcEzKeN1Qb6MdZC18fmt1ctE087lTjFSwLPDiXJoVCRvnLTgcVw
m/i7S+pTJeAGs6Dno4M09WYSzur/NgxgaFvqHwEHUOi+KIUwQnFELfyzP4wiZILF
SKzMYTNfHfQSMgXilxfHKl31j2s40cwpKU9oBOKcyCFYHuQkU0XDzbWN/xcgAgS5
x914RZ+V0Qebcoolm77U4mmKOG8nDijhuiiWYvrICBnn3a1IQzU7FfJ8+Fsii7oQ
+RYuFA4jQxzgtCekuz1Xlt4K/UiW+HU2zcLy/4tpBv6nGqIY6IQ3jIPHdpiTI2i1
6sfXCVgaIennxtZumnIzIpYEY/tckZOgsNzg+9WKy4WaRgBbhXbLO8fm6WoejWD3
95D6BSqGbwHaIzac3u6bYO0f3OqvTfyxZVGvxm2xH2GbwCg2CwpXQakI48fmlui+
fhheYo6Y7y4GkU3yoLtjX7ZBKKGP4m156lKql6BIEng3cGIUd5wtskUUaDBaBm8D
X6p1z1k0cYR16tTVebkOycDr4zpRX/my+weEr3kfFlVKwdKJ/ry6fcIegHfzShrZ
u3jU0xGlpzdG28mgnYTAyEEcDVApwOV2/yPvizfLIZez0PEDT3j5HtvzbAMD6KKR
ZoWCpZxGphOUQ171MLG9105V6f69tAYOUoABbO4eAaMQPeskTzOE9ZF3/G+bmTzG
M6OWT57kzcztnUPSKTABP8FP99bbuZfLK1AHs9EqeIHXeXMsx+PNOZPOxJZCyrvd
MpS2Hjo4tLQQiUZ2PiMy4hGGzuUym5pbPvX4QaTIUnm9pkcZMfyhrNiRquBHRNb7
nlLdgSBD1lkMRMyvLtiJ4RVDFYjIX7el9wdY+e3JTIfmUEVhZb3Unlez+kHgD36/
to2gfZBN4O3bkYXxEn99RhpGJ2uHTbr9YxWy4Y4LJ88sMcGeEtzAmQ2Cce+QfBTU
LXoGxT+7QyxYE2Q9sxGrMZaa/CVg6lbydGdO3ZpuZ0VBW8DbSQrIP2pyV42Oy8op
c3MqaYexpczWsAa70KaiP3xu0M9HAaKBYnsL+i6vzjAXgahGMN+0p8kRHo5M1gcF
niZVVqwC1vYjvSRjidKXJT7Y+882tZRYJvO3YX+JpRnpwTOyef55Lry5fZ3+cnS3
F6xEO3NGnl4rYuf8p8ebByqmXh+usaIVmvWOPlq9x1L034549LuNy8E+reps7Nsx
9D0DwN4tpnc9xZKtK2Tv0ZuDpWu2PouX1MrxRddyVrHUNNJ74Bi5kUpFTs3sE6D4
No1FGU5fJ39tJinEn/uO/bZPNvoo3PjNxdIkremq/nq+zm0nC7SXutsY3BRioPlg
c71ocuqo4hetxULPYyW12sX26xD/EUcWR97ajkn4A8+EwvuO4bfJ45TSvnxD/Ocu
vNLt1CIMXIR8gQek00P5vHt6wSPG+miRwlAtqwEpGllGcBnCC5VqoX/WSiZlwArx
dMhs6hrA19AN4Fi0PV9WI+Z/VzZezDrKjmDww9ABLm3PtsXHAZI8mG8Vt3e5ly11
WBzkD7CTsPDJiotECE83D1CvhMFrAH47OrF4fcETm173/DdqSO6scb7OZpgUxS4n
hGFeZ+sD+3BRKAtzSCf9/p+FqkpF76PWqWn0uHdojTKXNGD1wmvKyX73KD3m8oiw
e4WmXsGECybAL2wZxRLD4/cH3VHejuZtXxGB86fU9yP2IMXi5NxxHGiMeouL9mnj
wn42LXakFAfZ0aE+yXt2DU2i2YP3Doi7cKiPeMOxbGxAMbjJFkMK638qbxAk9dCs
qOnLc5crtjt7e5QcSN8yApaLli/0GQdPsPxeOFDR6wzCgeIsqUnLhaTDR6VMTq/c
8U08qmuQVZSAcAFQZZfjmDSMaY+V2iXvww8BaLo3Rs44fdjxbUZvG2ZkWDjMtVKp
cbZX+xpD/3P/BW02SWe0VwxegBf4jHoPYUGcDB8neGXSzCI669RWNP/swJ1YhlcC
sqNow5+zxVgYAWjb2sddEYI5+cIGPYb/2zpHLmD17Zso0/zMlbFVCKu5BLxO6Lb+
pqoNK/1SF5f2kpiyQXdDFkvMqr5DDhRUzOoO0iJXxg4Zm3v2QU/mAFkQnK3sjFvO
/PC9PoSO2+3TJFxf5x8Dxpe5dfOUxDVz3zHsqgheIY5kGhJfYslQTDOFeInm+XuD
nI6zZo0DS7fvi4m3TJVkLM4BMEgAVXDksYT4E0VoXKIFr83rsY7Dbpdbma2+XEj/
8a0rbAJj6a1sc4gJF049reCvYvODB5oFX0gjHJ/qxecp7H9ug1GtCTTBgl5Hfa0o
U0OH0Mi66KKT93Pa4I/RJGV8jN+ZfoJJR5njYceUrhIX0s80B6cItB2hhktvPYs4
lY+Z0QYzDDV/VnMuxL7K4TQahsAXVeeLCbwHiHwvIandUgN/JrYqa9BKAdqy2dbg
5P7zaXkx1i4J7f69QQPYFXqll95HHuZytfLn0ZtjSDFBz27AvrfyMv3kjDLJXvRr
OK48OQfKwXM55Km1/mctzVLosc13Y1iI/iWIYU1ok4oOs3nc1OLdeZVqocPhI3Aw
dQmVrkVR5hDfE2kp1G2HRb9LxeoqyNqMY89Uv+NjCJ2C4+Q6ODeSjx9Xq9EJFDjK
gwW1Hw9kGyo+jc+TrW79Ah+LMzbhJAI16XGiYQu+2xEwbYvWtXEigWtjkNrEnC8x
4smrJvM/BC41TAppg8Y+M8DLz/+evZSVHM+YmwSBWvJrxlWVoPQjVN9MsN2PeAH5
vm8H/NLjMf6lYBSkNEVwvB9exqzIcONs9KbuV4KNYW/Mgm8slj6vsqZrj8RYpTv6
X/cGQslb4E/8Yrw1jA49/QexGLk1zHyrD/Sovu2N63nQkosePJOr3btrr8BZVdlD
0KpJBpA923NOStrDDjO5Wz/Jpzxufh1pXP617kWkSMjyCNKSPsSpwODecMvStuXS
OOFRDZaiRC1nh4ikKjHADzwxU7NFe0PMhIXr9AVLae1ZJylMG0IrUPUbbSlDiQ/p
b/Qpl6M25AnGDAyz2d1Wmwt1DKq31H/LfZW9lMX9OLmhwCpV0QszXOnwarmGSIeG
c/dpp4Rdk7JhuOfhMGL2NUbQgzB2kjjAZCgjoNebJ+c7hSmhK5uxIjHK0qiTU4ze
D44eyb+1gcthyYmpbcyQNLIgi4Ho8rgIqkh1fsd1BmLrSQLTpmv0bBaPYVZ5chYn
XG/S0tPBh3A6XyWzV/1XlN/q/nOWZZYD5jMbIbbILugjHYV3max0bewnKADEgaqz
8dCF/1elXxbjPU0seVutoiSAUvMaK72NmTxENRQLqtPaLSoWPDU/Ahpwat8oanBt
OMZlTk5EiMNdrs7i1SX7Dq7OOFsxUqdxn6itQFe+owd/PamlkevEud7vkssV4WJU
RN4i/Ozs0Ihtn2O3yU5o027eE3m0KK4aVv/lBXlD/cdeWVYeglJ47b5HxsDf765d
x7OqZfl49oo0fxOu2FLfoSo/wu7peHEFuKMrLyyK5naauH2YYc1Y4NyMTXsIn6gR
v1EAGZnjq3AAohdYYTr/2FjbWIbKQit1R8JrFzEGBocEF0GuYnhiMkB/w6ATEdDv
ZClDTCvEGRCQ1YenvcLzoEOZQoFRfSSJr9yfa7nkMZI6ETaPfN0s69qLZQoRlb7y
y2RjlE1UXCGtY991zx5lhxeEQS+HtOPiQ4T17Og/hU2XB2y+7/Frpx+tdGG9BmSm
fksZv0Ck6lucT827b+zUVhOa915kciLBqUxSIq7Pxe71jIZvvZgpzLMGInycM4/a
YHjfvCRml/qyN/zU1PRY4+8pngMea4diTmJFqtqZRQ4wXZC9sMwIThfjYo8c4uoH
ffdiwMGygs8rhKP16ZUgDL0sG05fUbLRn8oPiplD68FLSXec9s7/2T06/Oc5Duxk
EncRefPFmj2X3DanDw7M7uuImSVSyuy3ju2ozjT6sGAUAJoT8fQsXZpXE0eFN1gC
Ua2N2yFfTtTyDX8Jg5zmiZ54dI9FuXAFDoGYiCb6drskXLog6+uy4Oi01N7KTz6p
/nke4MqBzeQuC9X6IenE6o20mr0bQGldHupf/U8zKHkPt+ildfH7tkJkB1XzF4eN
L2x7XhNiGfn4QpHsodgilDN7i3u7xBpJd+6CekbCjHhl54jGQ7kWCyCAHhHXboO9
wk//JmsI7/Ez4XuJ9IfZtfRrTGcWOgou/7EqJWiVC7cQtLYUcDi+TPi54mVeQSj2
l0bRRfq1aMUuXgIGjUNA7y9TJWTxryPw/SUpwcqkRz9WJE5ja8Q0/h3NIBwAHL+n
X7AJXFl7O1sCi05uTaN3uXSbnrXWoeQIK2rpRjtZFz9MmEdCib4RIYEVuZpm2a19
IuOJFA2RYGBnERWzFZv7WXzzYb94JXDtFCKGwGVUaIRp6GJGhoYME5MGkXQHF9bn
4nz3mVgbyVC84vSKt+B+d7NE+9JBlHwBMx9QB9dW5x5tY0EvMgaT1j0nc7zuuXpp
2CLsKiYfY4CJOmfqBDASMMJeW8SxeOHf1EIZtVkzLk2o80bvRuX5S6HqDMv7LUU2
KhZJfGAkQ8bvoYAsqmVI8wiHIrY1+dyxXkDhYnPbyA7m+KXTRiwFH5Ja6BWNS8/H
IIGDq0rOw18yF6RpYxgh9dbiZA7zpOz3UM2M1WyV3Id88hddpVcfoFOhUGjsYc0O
Z5emneQilmErPwqw2KODECnRGw2Hd2ygPycOmAmp3Vl6+0w+UuwF1ZrtA5Auk3Fb
lMfzZjE15CwMMnFzRNC+xiKHLak1vn4lIgjSJMyXLKsNTjdNQ/J+kB2u7VlV/MNN
SCzY9WpRN9pDcVZwdsU0g5L0RmbLMy2CqKnQi1c+taTlTsxQl4ic4g5YOU8+Z5Sm
w7O/NDSudcwJ3nmXSLI9H18nLkG1YNwlYwNA0zhEaHRceOiokaXnE+EX3nGbgUlz
3VBmmwNEhcYxrn/jW0nWzw4UpwuFPSeliuZ0gkNjO7qc14A+1Z7OSAN8vUA4eH9+
7UY/YGRgrmCIwVcKmiCoy9AHvXKgbac3DmZ8nK2Zi6S6ywyBmr5tR76YsaBjq6I9
IiF+Tmss2sofI7brO0A0c7CQWkq/fMPPL1JmkAXcDHzAjuvQA+wozuF47VlqMnRR
mAqeKPBpXAmoDQH8P+bE3QCn7dM3gMMzYH5h2FXrxC0Uz0Mlua6hLRjFUinD4v+E
IZljdn7659eUQEy0GUi2HIO51I9lTq/YR9dtkdWrHBzpYwrSc15WwYzIsjZRxZLs
SQ95s0eIFxBLqLzpeuK86+nz9k6vu4BFUsPBqARmksuzvbOppSXmahHEiC1dk2hx
p98iEiN4bfB1VI1fIV2eVNoKRHAVBFmywA8wuXAFuWDlY/iKsIKVP7wm4mKXEadB
Msp6/S5hl6TvwYm/ePmw6eLLmpHFoWpqhGISNHnz+efqMBoyyqxSJLqMspNhEcvX
Vk4+aBTCYS5zEL/MbB87xSFEGyeFTVrMv4mmV6K3onYkrL0N8fDqIGAbThdhYZ3J
1GPdENiQz7rNCrMSL8b4N9W9K63taBZ0YREvP2zVCGsbpCMQwwhJT0J4GEryIIqc
cNw/JPvhfmkfHqlGqwwifZEye7GBdbeHw/188vk6Mvh/Va+x/0F01wcPKhBKbtpZ
oNy4dP/CwyKFO7jkgCivgT+VLLRKT9uj2lEp/ZOMUa3uxFFbzSNI8w94yyP7dfuD
snc38LmVMWeKKJBh7lhATg6Mx8rGf6c+tQEGqIFASWoi1BaZeHBqUvPRDSmI4B9K
qnw8p+JYqOIr9bXdtA3hndmOtx2k8jIulV99mla1VOAxAcCtXK1JZ7CgeduaH2Vl
0/ubbMfc0pDNq1z4E0UdsVw1TifCLwSFuj2JuDuEly3x6qK0ed0By3LPk1wMqIf3
pJ6TYSoCr0IxwLA7/wLVjIgzxClyT7RgtNqE2wHayoCVJEB/DlKxTP1Nkv1GCVSH
8FMLZSoipm5LRPsi3e5ZqU0EKM6gXMDm47k59mRMAKsfxSatKpXYT9vr33GSbkUc
C5ehIIB5G7RYTQ0qO/T4S6K6uh9Wj65fdeL3YETWMuRVp0FSJAPZ/9VuGOhaPAK8
fl/pIGG/frQ1I4zlnNG9vHeUNVrVF3R1J8e/cblz4+cHfkPEHxBwhOr3ElfszTMD
1VnjHVhpGsmHGJDGCHgrSZtxe8Jnr/J2x1+is4vGX80Eh+mWfUzdQNAixGPzsyIS
jOzFKOXbZyk3dahh+Qs2glQiJ4qV8ik2UcjvTqkmT96K8OVsbRbGnCizBDkvtY4K
NjDiSXknO8xcG8a2ZVSiCVKe36kHHhqQ5QhGejBHj46Nk1Bru9D2f3wl5qED7OJ3
HEm7vo9WVABegMVzz9XlsY40SJhHoxEh6E1tg5GeAWzYvPQWjp5nU5Ux1viiVkeF
8CQNvMDeWVpKeSkk8kvTprrvizMzaAt7DA1T/dUlMulu6vRS/1VqSUjLFKgBmV2c
g0aU0Ob4zveqLASOh0LqY1kZ2/efGsQgFT9YPG2Ku0amzRrhGwF+aMsPjpEjI3UZ
dkIefkC7yK/tO1ziXi2RaraEnWX8xG8U+yPdF7bBfytxB/bbIXtzVaQv3qC2U2VZ
YqBbj6yDIXCxGvEE42ye+2JIXXK9yiPJxQjYWE8Edfj7RIgwVBjmEwBBKqwzW37K
kLp7kxo0+koAAvUUrg324RtZXFXQlpn8Hv4SJs4thFzVc7R0ktxQdXkH0A23d7Pz
kPIsOy8OLWD/q23d5b1tXw0Id65LngOhQlbOQRYuQqmayvFjewJ80pVoyC5aT/JU
ugnpDLQokD/fxYvvmwQpjE3+T5o4DVNCL1Hp5J24PqFfvtdl2j4oxtn08Ym2blvE
F3+OgX2Z4KCoIwfpyQLhxLE4rWI6EtyLLkM9p2GRjZ+Ng1b5mtuO6OlUd6y+vOIw
S2rg9X3PDPhRJIcNJlm0bpJnwtyHkzIENeHWVp6nv71Uuqv5gC9Gn6pGW8Smbo9b
7sEsaqozAHg3StmZ14w/jexYFrddoFzf8Bb2y+kvMjfx4CDfHqY6HpDAEQaI+XL3
IRTWkez+wZZsGgBlvkzaQYis6HrqZRaPyDxNIxrlqltZ299m/D2+1fqsb64gf+Ua
pGahbQai76q/owBRyoA3g4jyT1ZP2J14j4VtjJgOtusM9Z88pfDAbkoJjN6vTO/A
BVzMkGD4lECnKWF2/AzVHQIHxq/QLV9QWI2t4a6+3SAzzkw+31Rm5lxFZ6Bz8uIG
ygAa6XoI7O01Ta8fs1hBrq6kNAHzNkzrulwWf97L1beMjb8sagvw6jN1fCPhaUgt
JAY5DnMLH3eVVMyegKJQRUZCObVXdQgQayGIDjxvLYli/ZlTXO65G5ylA8pw0JW+
aI6jZUm8+WKYEo2t/L6ZINBCYFqTFaAQlJKGm4KVUgKG56n8frVuI9RiRwc3UwSY
dMdv+TWNTf7xsE7EdAwltidqc3eyOtzCYMM9gr4+0pXaYko06zDR/txgbtKvrWnb
pqokPmrxH9q+R5KWu3sQuWSk8RDeZ2Krk6/lQhp2Y2vFxi1kDC3G9b/QUbMpN95/
RCzAzgYBDNR4gjvo+GssZ9PUaVnn26LSt1be6zROpJntlikxFxDATuNfgk7wJW5n
CoIZ+lp/GjIYEABhvkT7VtTRzLLZOrOWEK5mhTsah/WBjqR2wKvq74OJLVJ8h+3O
wZd7sO2rbs53Rs1LJEphTO/oHbzYHTXhII4MwLOD/1nOrRMwZGO+xXdM/CTncBrt
rlPtKNn2DGyrPsap/JTLLF1yXrh+EcsCcOEXaPYfbIfoZ+ARxG+GwVsaAb4qQI3l
YKjZl+sdj3mLVEw5Om16Wp7colXSsXxm9256YbQ63nL5AJFaop2mM1AnLAhTZAtz
c+QXJ4WIVcv5N41enSEnIMCFWRj9asZBlsWFAwmY/Kk4wteriVuhfoGJvmh9k3bv
LwbBls53WQiD6yi/0QoY1ZkKFd1SN5qLwEkSTPfXV3tBtCIkb2Kl+EkSLgcwifO0
PuIrog9ypoIt8Mr6iIkD1pSrIees4zJwSCYDedUeBFPJjwelb3ZQAeK85Yf+DGWF
DqLu+u4JNiLPwLK9tSwPbxpSPYtaJ6k7WBXWitTGjdJsxAOSY68JA071Xmdg8I4R
cBSMxwyL4UuoVj3qtV+YXH4tPgbhWoddrJn4frSzpHlv8+cWmVku0dz7WOHsK/SR
DxWkKsBxmXTerO35TqGTRs3oO2nGYqhIzVE/ME4FQPh+5kWUp4XpnnJjCcrVldYn
b2ea6WyX+svGPdroVJztTidoNJnE/taqhT9P/VzxkCuspqHxU+BJPkeM4XS1WW+M
N+JHrSfXd7POvPecMH0JRdwI3w7CVImWMbA01JLCigS+vtI296zRHHqBukaMRPKG
v9HgQS7MC2dkaVKGifpoico7x+OTlp2vJheJnXHozmdLTn1j5Z2WEc4F08gg3DGU
r0QPKFmJbodmTH3IrUGV4vabLKUXAjfpav1wP9UQ/HQGltbT5WSRHD2g16pT/DLs
+tSW74/jV+sYQnzbTpFYHMMU379UG1twFcCV+2P7YjBeijGlTuT/JJr0Rg9tNfLS
nbjSqOxqUCmDYsr5hfzFbgm4hO05wqqOow5au4TgBBB//lPZydz5Mqy0iNqgWvVp
ENiZSZho6+nHoRnc0oditHof+znkD+0OsJiEmgpYqs4uPH/N1AVSChkCU8JzULbl
rUESuquDFbVOCnZ2do3Y9wE+CAjpt+9mqLi4ng4xvURPzLFE27+Pt7d1I2I9jR1r
1qpoYcwjzF32vmDXvcl53TTgTjnni8+1P5T6+HUhP1KDezsCgHlpwsCmayleTRZ6
H/8fqsNf7IkstNoWEray95IjI2KHw5mlXzW/zSb395o5dw2CR2GaBYEaiVNBemVS
9thxk2Nt7h2SZDjK09VidUmPTnbS7gVM8u3BhU4zGR8Ghf/vSxCgZtGIj1pyu/pO
sTmWI3Xe+f8atwyyDLzl0VID1iwq8QvGyBsa2Bbl4cUJ2Nm+AiwndQV+YCOs3D+P
0uZ6jkfB6IZ42iBIh48/3nwCRKiYHxwSMuC3uTHRNXOxzt3W+lEDkyENfV9Wq+6n
iK0cbsE/BUvCvORLFeUzQnVB1sRxct3Dv3WkiM+tBpK2aaLCMOxWKsrAjBgCsfeH
k02cIBsBt3TeF2E3aYjPzBS9GTbv6Tu0bAwV1UfwUeDZ8dtW3PJTNGzHlS7M819g
xT+DoShGNB4yc066G9e4VEBlMUO49t7xEKkzLMODEfI7Ql6B/E8AAqKCmsMVoltL
MrzGmiCZ5AfJYmiYv96yWqeuGiYzlmFXqh1k0SJ+4lXhRxzQ+so0AfcoXFEv7t9A
ZVX8rgleIFmATdvXDJCke3UQpd4Dhxkmzr4Cf7WXQ7QxAe9wo75GyRV5niXS/mAp
GjEfAAhw3sd3KK74CzMs7yF0Eb9NnEbIyym+2zcziiMZa5swpr1+vntXG49zUcz8
gc4a/as8rC4cECN8hno+B3NGbjSAEI/tCOJ4Emg+dijy8TBGmpPTA3k3oYQlIw/S
bEATOqMOkIFu+UgPjHJc5fpXTVA1C8n1I1k08raC+/cNAg7lMioamo4vVyDYRUbV
/jIu8BLCg86mkmH3tl3DKdXWhS3eqTFUfio2q8qcIyAWBcxJv3Cjx6w+IOfP53oG
yxJOeMmXeuJTWX7KIENaHVVlbwmrK5LcgNbR0vl5GKrewKuvMtAKG9It71ONtuPW
UnfuFXW2uxs+8s2az8NxhJ1mtdIT6hE1W6zo1fr9w5Fw3edzRDOzINSHNBihTFZX
TqsioLw8hiWIhsFXAyh8bsogA5r2B2iNH6zEzf6u4MsgrcVv8OL8oGG7qK+b6nM+
qJ/J9ybj9y9dd1vbS22OgkuFQD76cuGEOZPkQDWgLtNTTiY+kTkl3LhvBBbCQyS+
CGOClCZ7U5MBpsJlZzVaNvjiddDdvAYPrCDSzg+G2gsCjyl0fLR0nFF5XDe+PYAt
7+78wl6ifVsttx4tRja0+7B0PLiSRiuYn1DfKsMEv3e07Dy57xiLAN+Mm4MUQ5mL
gRpwkl+WFRxZf+HNEUvDKrxRfiAo/VG1+x6uXI6r52WgBG5kU8kqsxKtFcsH215E
LisbcG/ewoChBh8nerFSwL8XaI5PN1qFkTIflwiAkB/UZ8rPoQDcbhCpIwNX8sL7
1HcCLQlCZxiYars8pSwI4kEiDMxIpWsMVWgC0bdecq6oW/wwx5iIRZ2AN4+GNpVF
MBNchTAG/isF+HSzvEU1H5bwcpaBmdryTN73TfoCiqty6jMD5An+aq9mjqKui8Fi
xVpZd2a/h862b9ZoNXlWmWBP5G48ue8S5N4eBVHJro/8fLLRBHLNJlztryA2jnpm
uKFFiDtAWPZEZdYI3+eIONAQBIPjmDG3dKdwn7vIYZqyIKx6Jdjl3a1VIzHOvPFT
IKMqQc4v4Tp7zptHN1T/AQOAx72EgK7Bk6NnlJSccZRX7UAntkBP+F6w0BRtmmr3
tFNwUC6N3WCsHrmHmR1dnOEH3L5yQwzdUriQ08xvOvZ+/AopEF5Drl7mnUoCIHWH
MVX87ntcAd5TrWfOmFEah3t+oR8XknnI5zNS/7lVSwttNetjwORvDmKpkvh09hdP
ZfX9tY1e81HVtrbfCeIefJZ0Z6EiULg5nBNj63Jedc/LzE0dRWYq7LY50xWujEI/
qculN1Ny97M4eqrCKHOgzmfKSw+b1xrEyEmw86lTHpe0JLC9dBbLOhg39VXXkWCD
5WmGVB4mtzCNbAG60Uaba971MHO7v2oTuNjktBWBR5vUc/+6k7V2M95Lm7eXvOKF
1BUXNFnZLRWW3vn1drvIhSpGYlPmLwVBu/UozG7o74mU9r1xVew13C3XaBUQZ7sN
fW+2VM2E+XY/fn2lWh5SiRwoqFmrRhoIyHTgRVabR5qJJJUg2mJLeBHz/M/jagL7
c6lS2SsuKdtP48FfkRDWdVrNRAx+SqkIJLU9RkvcM4/VNcYGlTHTapMMotLgouKG
zJ3Pxd+LkJ+xPmPriD+5kyIFRynp6MM249x/68gaxoC3OIdqstUMGujpZZya/Mbe
usojFG2RboukmYeZKjqxdZpIB1tzWjLihqWDZMPjqiPrHBMEhTXBSn8ZbwDlNpeK
OU3BXa/4XpJypRx8ERFcTJFhKDBi3qgQjrXNfmTdzCjYCANJX9VaZrBl0vITznRT
aRPS83sNFWdMXSStx8WvsfH4va7JXe2WWjo6bdZCnnkDf41Zdk0HXKEcT8OXeEL8
vPzolehDGD0n2Jeg+6Z8Qd+4M18O4gpeONARkl0p371OHE07BjzD2Y231uG6u1FW
XIlLtEdqWHxEN/ZC4TNc+ZpmBq7cc795aL81xjJpfSD6btQWZoZfzYUiVn+hn/PE
7kMGkNKGXfGsvnbKmU89b4CGFgz05v4weDc+En/wctOo7B22/2dVtO6k3qgt/n+0
pAeGUw5FPeVo8GqwqlvH+VzIgTiPCNKavdKCRiENeaYAYz75sxvSUuQsPis82OQu
wV34FuRtFS+ehM1V5LR0m/ntY915y5o8QAVSo6RPnQRDY3itzDaEDWNMj4n6U68d
pUWllAABsN2OiCPazpJSe0QGSmF+yghjL/mJqeISnjyhE42mcpwlpBCFwJjNXuYj
ypUtHegE2cW7F9WQ82Mb4DvRDubBoBnlREuLztaLmYiLlIAKf634OdHTyA5p16Ou
qQLKNm4/O7rWM5lXhjFNLd2YKzV/aPR7Eq8HO8aQXalBQ4iBXwtofPpRenf56W3q
/NrMFAHKQQhqabyMnZUYM1NKp49YQ6bFP73g2NDBqZKKw6CqU46ZvXxV+2sBuuB/
8sLl+bn/6NSPmgEBIsYXHbuNjYASwBYIFcoe5MLbnsTEieCeY8k1J+Jq7VxQ/kYV
r90KXBD5ocJpxFVOwPaNCU8a+6lt8Ad+fwHGkb7XdCQ5d5wxPTrq6EcE5facZIJl
Ugsx9LpKBr6a1N+4/AaWyJQw+PEiMy6kE7AXh8rxHso4EnqaCEABTX0nDxf0glP0
XYtzWBk4Y3ZNrloc++QJcn73xSL/XR0Qbm0Jc9Dm2OdxL0NE4Y11EKaJ9aaYPqZT
Wx4KYIEWeOSVbECGJBRRbwLF927BeyqxsStCN3XisGxlMwBhhki3DKX5Q6944UmF
YRxyon7qyawYMceb4pX0zuqGXi/U72HxRYhXUGc2heMEoDSCzOycuT95mlWDo62T
LvHaAt9NJj3eA99uEt4TEGVemFMbl4GDXAUV6rZNNx1gNJ0BcgaMzEQlBBKSlz51
QVFSd2mJsH5xFTYyWwc9c8Ai5Nhp635CJzIocvWZeFYGDJDLAVthwwD/8mQ+niiS
6pKECn/Dzga/5IBh6Nm/xTE+LaHp+C9DSHoH4GZUlmkczKAx26SBQO8izKoy55av
PmhUxFVzM86iRKH8CMD/5II92M7T1fwKweYW9XbSqw1giA6n1JCNMQzkbvxxEIgf
u3Ko4aHlX4RGuVABBt6dH/i3VGu97cA91ZNqgsQk5v4URPl/9pVeCp6p6Zd/ImP4
JodkBYIpNe0TWUukvL3u6VYUmDa6GMl7NwyoMKo1/iq5h68N4LYA1KeZkbdum49K
1RIkza3p58AQ9Yi8zUxxY0brEJKU4fPO46POkHqNFP0g6jiUyrUd4Sp1DsIOPnqT
od86vnrJHOp020LYl58ovg1/bDx2fH37dUlKfIV1ws/E/AwfkuL0ojHu3bauX58T
fYG5oWZbwM9Z9Ky48DkSJw0uHPsrdat3kPxtIqKNEvg+/YrthbqhAis5bux91nbD
qpM39IQmGKbEnjk2NT9J4WMeGmzjNFqWpxn7/3RLTV2iPUWrvP56W2EBzuH9CLQN
ffnC95GQroONT65fWkUo6TlXHGt9paDuUo3UXc/hFmNZmilpUKKf5Hu3kGYjEUIZ
8VS4gPqpZ8z8V4oVtMAHplNR6XMFBX056UoyFPiHIYZieNBBO6zSPVodJj7Kh4Zw
TLd8EkOrzThCWzMbkJDyh9QQQ6LS/2zmY6yrg/nzqfs8+khVWNlN0HjzYtYTK6MH
PeetNefKBXoC7G5v1KHyYsbu8+2jmxTB9/E/rt6keadZBMpKT1lK4xp0GDPxVvrV
1m4JOb2NeTepzGrXizd5QLqqjBVjBrV17Z3qZECEFH1QcT5sw6PxFHR/wMHESbTh
9FDwW/13rCvYVi5K75jPt4EcFvqgFAn8Wf9gCThUT1OWXw1yXkXOzivmCHUlCiIx
/bvgWw25ch+mo8377FINvuziVT8Fik5+A+ap5+T+EN9DBBnxkJgojuUoiKBcUegR
qdPHw3TBNrripgSmJpRCtGstvgcJVlfvBiEJoEKa4n/lm3uTRmFZrd/3HUQ4w7EJ
WjdYG9gdRVrN5Icq0q/tLpfM8qyMViqog1DXaa9b89zt/fkF/Nqnbzsy7ZnV0+9Y
owPTtFJZ1/AQ248qbm3wqtYiK/NIF+62CHp9YPSkIe+ZbMmco8Gp88C9j6BkFr5R
i5maBQDa53AtYpM/J6MOUD1UL6A079H6B7+hVJrtu0X86EWqcfjaXRdAuPjyZFB0
gdQHVEWqIAE7VJ01+7gpupM0DTQXATuq3aeIuxJjsMSRmJgsiaHgxUSA/i3Y0YOI
knpx+1vyfB703+JeIdqWcLGIE7wGphYKYcATQ58afHjUz5qAkAQQAdlcaWeyN1fP
gRiOSe0QVuV0PA7+gWOtLmHdY7u5wOM6QDPWuvArhgL5GRnDE+NRvhnWpYG/mfow
BawWgboZsN85R3jAXhMXyhpMtgtqjdHkHnWtAyM0QEeACH0wIDxwaKCQHgPy6CRP
OCPyPAOrTf62J1rAThqsdrHEvFzi+iwZAE4kZGR3QB4m4EQKQw/FMcqoBE4WKIxZ
BvndHH9EoHitWgzzhlawp47chNtH3U22WCcGtz2Q7k4A0hVpolDt4inYsJw2fhNA
DqnvCtgqBSkfi6itNof2z/kVKW86Ae/seQ3BoO28wpq8oMOFzqC6yTM57528+Oen
NAl/R4Si/RaLlIFoF0lcFS1ZZ3PdbJXpVNbrTfKmAtKmA5iYZ9emypjelqTH1/3p
9bKInmIMDJaXDLWwg4oYG4yvbmbEOP5f/w4wc2bW8baOShQuymdtVNbY+MsNk8ID
w9tAeqtXWWNP1lIcVMf4goujyUfwSDjLFj3w4SvegG3589v6LcWhoEC8XTKP5re4
jHSA//HtnWB34RVr3b9SCf22UPW/yJ2DsmziOZP+SXNhepNTmbrI7m/bpUBaXm0+
Ad+QIECVoCCDp/Hbx0KMQ8SAGd2DTt34CDgu05EWauRQfH3No9dZhGWAo+1Cu7GB
17xnXoecIIBEGP50+nPhfFFG6USV94KZD1sw9TNshHLQYGmh8Neup4avmC5iqNHD
ta3cm6YzUJL+qzBOePfw/wJyTiruO1vRhsGA1Os3kSsFoh/rj2uZ21MrJEg35Fpl
WxRRRwPytbAjktYF46t2dP60cVlJ/L5A3mYc8zGe9H01+IpEcud0N7CIktliBAPC
/R8L21W89haRw73q1UkLsCSTGaH3xPTc4L/s+Gw+UONY4JJ6ikFY70G7CAJ9yTEK
8lr2ZpEru1PcQtcyipvIw8vq1dxq7welha3jCVtQGwkRyFvQAt/G6+xLaSRQ6bdJ
BW046nYy+MjgGIpbrLKN5gHkFrTblfwl5voR4biMx8Gvf/0cd7ZMmyiKkeQDHCb7
8ZpvwhMD/nTtw/WIYZ9BnAxqaESfrIblF4hOXO16PI9cyyIQdLXtoP9uZjJh0dBV
x936y5gP00HRIYySKwXB0hCGKmiCr/SjwLcX9mx4BCJvJ/g/KaCOCEMFSPKLwqd6
KB1QAwzXcKrt2pNF3dFDyHtk1THrw0Umj2VUtP4QV0RByZl0r8nnBMY3bjjMm69d
miisiFuuunfvccRX4A2YueYc79M73kpDD0LJ5GLd8MQfjHiGPtJ27uCYcnRoBPqR
1Zgsn9GrrwGJ598GenXnzV4Vz2TCAUKzWk0i737ldDaPMLavFzPsEkMV+UcrYxzb
AenZ7QYKtrhAzzWVGbuGs2q47NOQmhA00Rs9xnt3rnzK/UCsXwEAbGNAZCza462c
jICMFVdcde/IsXCvxHuvOrM8KW8xhBh0T/veEr6dtfL7ls+N5ZvjD6WFzQxsHAt/
t5T84frkhpVMvJPCRaYj5B2A3bH++1ICEKjVSf3Zlt8pebuDkWR+PN0zOQLVcAx0
54u3+BsOYfQtPBF1cBjvAEIPmwQF7eSpUqmdl1TDk1oKcSXsPnUlktegQZZyj6Fu
HRL54ddetLHN151uLrjsNHhDFUlSvrbYt9qW7NSA5I4r3VURspaQzyAxrfwRzoNz
OZteebJP82PQCiIVoPZyJrOC0MsUHnNH+WGnDnuJV45aya+gyXOjoATooTpVGWhU
/WnvlVxWnzCMqn6UOhw1VI1THAUXyFpfL+A6kDCemMwOimVgCm3p5yLv4eQKQkRB
WMa5+zC9lBFwayCG+1O6DHDGqZ/spxPuim3bJuzblI7O10G3fyK73ML017HxQzm9
gIWLlQAFJGjQs2p/OpenErMtkj1EFZk7X/vXHTnz7v8C2bH7Y+DerU0x7mQ7Y74i
dN63brNAxA10h/xc8htQqnBi/eL0P9r0L4iBTtNGE7YtQ2+BRwZKCccbA8bm+CgC
CmwXA2L1/mdXD7w7qapFMfz+WRc3/uZC2v/1EIR8uVu7wBllkCaHKVTUlhF2yKAl
yaT3b6C4V0CDjW+O+J9HEIRl9cmVCjPpPONP6Nv8DGrs5mKXeGVAX7lYECu5GnOV
1BndrjUGe6ErAGWPhY1iB3GZfwM8ydL2iv7HCX1l57KLE9OWxZPIzCdjCWsYnNCw
zbtxnnmFMYBVqjfmBzGXe0SUBdelm7r92+c9qXnPQp87kJ/FMxKrtQkS2QOQj+jJ
UQCOGKN2tn/Vsz2Erfyo/qAeRzxaGirtPmLuerKpW95qth9xH+RqmXgv6zdCaq6c
cRaoE2Ex5qEXxqcnoginsfpnLsR7Pc4mMBmLN4DeDiQEfX1BHbSooIMUVfbvYB4l
XspHBhMV3VdbLBPYJAKBOlDYM/lGMWamWlHv8Pb76jbYNw/DL4A5Ql0/Xl68L+cs
RE0y+KJu1zbP9lE/y+EIaVq504TMoi9O9i53xk7bDviVC5OOkotDQHEOzDqhsOU9
IpscQetplzPIF6tiHaLIxQ3jXTw15WwpWSV43IkeYO4ers4O7wwKvD3Sf4NfzchU
pVKS38sfufC9Ef8YTjWNqfpYn9PSU9bI/rIp74zsY7TEIzBW5plm8bo398LltY5o
cg1jy7NwfMd2M9LLWLy3JfC3BcHb0HigkirGAWct/YXCLAIMAx4SBvuuh/cOeh99
1dQGcY4id3JSw6anKLz/tGl5PCAvKp6+ptfW810Gl1lYM2HbL98PhFdDQuvmLMHv
az3V70ghJYSDQp5fZfdeVn6P6UkDUPWOa6idDnbR+bhjkCvMLN1sSbVEjMXGkReW
o3tSH1szi7iLckTB3Ki9eUdcbptwKYQFR7xH/gXOK85y+lq1YwSUMGaevdAzZ8zz
Y1Ryc3KUPhCQk16wo/6njSzpWrpXh/dW6g0DD4tesLjAQwwSMrcFXnwtoaJzzfO0
x1s4MSc3KWdSkjQ70tGXemHZRvPb9xLOHPotdMHzfwJGK+/c3onUWY4oYwienRhA
pIDEMGmyTSYsQYwnFHexFWNnPdTRyI9RhbhJGu6R+mQOKdi14aQic47MH+yiHRzy
0eO8yfzXHR6ZwehY/+cJxIsYm5qVfPJNzvlDlU+SYAIJ+j+qcV4vfCRt0/jKEzdQ
8CTGFIuOYzj46fHkIsz0wRN8x2F3BfhC7gZllg6fF2cFRBpaBHvuaG8tJC/I1ZDy
9Xxo+BBkcUzEl2YSkA3RUD6K1sbzz97TEDvfu0k7Bbs8LCvq23VklvMIRsZaYFXK
V6DtDkzvqN42M5rBPqBEg5N8tjshTWG7HFiVdR5W8KUuy5ITuKnTCsif4joNdqOo
NqYNbHuluuXbI/eS/Y1y2OT7HRzbwujn9m18k/G+3V3llnByIsM8yBMt8TJ08PHL
aNb82GmnUaXvSb+rFQ3d9yqc/LlACIPwTVWqC2M30dsWSNPZQPxzdZIatN7FVDqj
StdXvpdD/szgvVRUK7MxUOAJxJTzKrfeG2tUJzrhPpcCazKvlJk8edxhdSMpAgH3
3m+czXZ2i+IFBvMc3b9t7OASf01lpgdzvnnMP3uiVIRZkZZZWcO48Ho3zMQ8vZDi
TD2N857abvnJAzAg42qjQludoBash+WUJgk2v3bvcNURlhQ3TaF1WjarLD73kI3J
dDK6lAxZB2ZrdcTmShMUGqSVphWXlx6Xo8kkw9Naamw2Inh1Q9AQrmXeEkweTTWZ
9jyQ89d5G9ivL4/VUnFpmOJ6oay6mk1GzH3Bvr1n7yR3gHgw1SpCr+MoSKJ0Pv3h
pMWp4JslyPIuzpp7vd2RBVJNA1tEv3xVByQRsG4B2w8qZo31kOeAQnXCzNe9G1dm
UR2o6IuHe66rSPlMWxskd6Z3nvddRR61HmzQfWP0jNKRUdcz7TG3hvWASRBiwg49
U3MT3gF1PkRfTebGLn5dIIaYPZfsk57tpRgKBjz91dqIelVHmjl1oi0lp9+MWQlg
wZNPC6b1D6PiIsadc7tnBrKKBNr3TAkVq28GbajI55zE+8GjIvAJhFZHrAfGgvuv
qgS85Z/jUdGTc7dfDfIBV/vmoMPzhejbsyuEAxGzkjzqLFAnjvvE8qAu/SE2ZYsU
NhJD1D90fxr+LeZvEhJ45K7c/jZjHTe3g7Tj47K2t7B4sOWrIFPEGZ3Bva1JUv9J
LgS26enflY97cWxa+HhpmrSoSLs/9Wkb1h29jswlO90QUQp7tR8lCS6p/OvZWaox
GChXzW/Dx2dTYGrapo9NI11QKx+NmvL9SYVxeBg9v8drvvVTwN1Z4Lnvqhrt4kx0
iEH/1OTwrj+v5IipM3gMHNCpkXx7fv1DjOPrePtMnY7aD6aaOdA0hqi7DFoVi7du
yZ0rlF4FBhtKRcPT6ZCQkRiE0fpNZoH/E0gPUUorkGbxWQQgefeyjiEABxN5Jn1C
sPvCbQ/GAq1NYLSgLMMik09INzgz//R6lGZR5EJm/LfBkp1NezLnkY0xZ0EooPnp
nirdKhY3EdpBC0c37gUIsqcbsiwP7cTTUpE8V+GE43AVz9GWNdzlMFRs80R45tTi
HA4JUr3dITV56x3eEk9yLHDOd0ytr7f6U+QdDv7zbpqhg03JojFangWxOf2claft
rJ0eB034N3cM6iKfIsmKcWIku0kXbZgZo2MqLT53neo0I/6YRqcx0eLBhLYw3ll4
AF5Lt+7HQF3hsGbqmLhpL5/SLmmBwhEdZjI12cnktGJbAZyohNnqSaQtywQv1G0x
Kfzenfeg2RFwHVhSmk9aAlSdf71SbUQVIzPxhhYwwaSYMty3JmJf7qhuPMVgKA1d
vbfigROa6KtEGZMZbUxGB7QElsSyTYOUrQMeNGhBxzbsZV8iLGCiCJm7euz9bvmk
C1E+2B3iNiMBBJ9NPhbWVrvLs2jJyoEUX4HahvkneXlDiwelPRoMvHpScSVkJ60w
Ocjwf+tERdNIR/pjifLgQuWCstOJiuLG4tpcWgSDk+jq/jGAIGoopz1pcDrP1FjG
G9Qy39Tjbk/RGlUyy9ooFhtYPP7aw2GqcvQamLaxXFySLo+wExZuEU/uRZD3Pm11
gKd3XSRmw+wfP1Df4DhjAHqlB90gh/m5xS5rglopoNli8QKa2FVkAQ2rarZWlwDq
GsoDOjF4SWeyhkl8vqJyqpaDv5EyBGxIlSCJatyRts3sayqu3RSZ8LVo8m4toFJA
5KejdU+kNElnQY0IDDS2EoDUbAdLzxp8eRoIANvbqHamOeY+Afz7ewpLkvcEo95j
f5mRP1eahkKUWGge06zMJXrDGr7g/dx6W1LNM5K2++eB6MFxYtt98Sp4HoTKvH4P
i9MyLYix3gtZck7q2fxakXP/tJz9EYITIn7MTAgRMPRXZMMYzi9Wq82wZzJgjGM7
MqIbirx9iIITT5184tc7bG5x2qWeEvTyCGKe056s3iYyrqdrTlaYDoKoX0CaFspW
37kWgYRKB0MI00q0W8wlVDefCqRt//ksdETLZd2hz9hNRVLw1BFLtWyg4PQJmMS1
JLzPr9duqm1DvoHIH9C0KuyAuQFEwuh7xfYVqH0vD832EG3SYfHLhUEdERaseALy
YvNwrrqs01XuU3NtruSd2Rmd/y0zUVUezwcrjeeanE+vtICudGbpphtx3LOqHbOh
YNiTQ846svjJWQlbfTcEo3ESY3c+bgvJo83CcTMsWfaSKaK5pEwiZBWU2pYl+2gX
88YeDy4BFjETL6QaXFWaNV8BrHCTWtQlCZHN8Bki8muOR5AEp6B2GHdG9tdA3bie
qIKQGVwqB+ixnjH0KXXLt4T13PuTQkz2JTfrz5EVO78luJOuBt500savnknapqH6
q2F4LrkuzdimKWh4wIX5lrxg/O3N6xX7vc/cOF7JwnjWBSjalZTMEhpagVpym3on
RzlJ+iPa2hQAasmq13QncBnb6aO4vkpTmWJ9omSJ831NC17T3Eg5XkZEiPD2d/9o
h7r5FC/yXoolV4q7rnVfYkx5srbYeaPvOGsHmvF4I+24SLz0lpMhGREvCxS5jHOQ
jE5ra8a7NnA9fLPFKHR8GTmTPZlX7Bp7YgamU/uJPKJe0e+wPbTA7Qd+3JWzJeDF
I2V93zZI6mPfL+fVZh11PuAQKVDygjKvbaQc0HsC6yAMt8Iedgts8U9iFXLckjV9
nWitVv5uDjrO9Kv13kVGBo5Uvysb79kat0THOk+w4Dk+zYPi2DcgrOfIv1gILdQo
oUBjMYgwXfF5/c0pE75p3y2cEcyGWG2ECGRh6FGFqfOYRoiXUQWEKgPU7aJXAeMS
YLfNDH4SkYf0bhpFi2hUJHpe4a3Rm+2Td3gqzhOmlOyyPH/45b1GwratmTt4GKcZ
NnMX2ca3PErDVHt6siIBGZQKhnARhWGEIbBiCvqPDaLQLnBdk0ATN4BT4ZZXJx3c
SeYxaBgXIsJcU7kTSkLZYECofXR2h0uwdY58vUiIJYazHxm7vkkrhX3AmLoJe2eq
aX8lGc96KwTKtL1b5E6zMhIMW3v/vAgVcsXKWVqWaIRTcaCq9RObSgaug5o5oowK
dSMt6+r4mPL31HFgnRdMlkhJyiVMWC8pCLhJySpFcI0s5u/DPO1GnME2Na3LxsnA
XvYVetmiLSzMCSimf7YibpRpOHaqwLAIQNRDI7+ChdvJkpwNzDUTEWCTX+wIxKKj
z6XzuY3NBPLQm2v98wvZexK0A+7f3OnNCN7PEH5/zURpGGvdqoe+NE+QPeFUnXX1
YZtPSuWxbNc33zDi4X6z+va+BsHLQHvLK9TqTpvpFS61P5+QPha5mqhNITjfal+5
hCxLFdH66kUyUoZaKEF964NcK7LgjYVFB6MrVYL51MjBWCQc5DY1hr/TAVFe5nYw
ofcFxfXNNWu9UPovHOD2mkuu+EZ3IEflHwYoqEwtgl2u1QxUfyLz2szbcvxC17GQ
ijBMDF68nsIG3Lze+XRStwZ77+XUec0d6Ql9yaThk7v5zYwoosjvSw2ngu2bzTSj
JEu/ojif5l+hATKDXIwYW4GwjdWfEyqoJ527tHJMuUsvPRvB9mZypAvKeA/lzAN4
Wu9WZSBalmEFVrFbPJEth7SrevusMZvP4LsFDtqmagb0wCKmRsMR+4YWRQF/+unN
Rql4e4qBFhDdsoIKDuAusJQIP+L7999jYPAUd2wOxcevKg1hiGA+na/f238K6xpZ
LTHJ+TXnClAjfOI1LmrcvF4TV1Mep7wRIiORFk8oLT7ZQJdCASstf2ZxTJASBUTP
O5Pv5Ct2kKIVP3HIZX0vL8BTqLMuQEfsweJLe9UlHviIh8xWJzNlkru/gjmNHk7s
9Sf1BCX2t/e2f9FxH1l3Dq1mHTndHO7AmZfIfxBdTAgIcXi+hoSAqkFYQB0lA93x
ER3aEUk1jIr47vxcKgSwd3ZlVTLq59CYPz0pPwMxP+t5gLyy9Z7VDAZzm0BjHAme
5xwCGLGKMhnNKKEH2h5PCilBGHFjWEzcDx+2wE0bg6QBcpLecQafSdFAHg9js4qG
eeMpYEv1eUFQh/5mRZ1sOJbE/60QOCqtnPBZhGCYuYxVdxY69t8V+XVg0SRwo+2c
/HqpOfDqcMiRyWeBFqVrgcgY4OMBz3RsS9gHuLsbyZ+LEa9R19St1KGV7k7YCyIb
MSoE4FQy9DoOf3cNq41VRqvq1r6/Vc5qpbTK/llwNBIZrPMp+h83oDvEgDcwoH6f
5suqiW7cQlXWOhilmdrpsfgD8KzsYGYM5ah25GWaDEgINCXcPuPOmephKlCxijY7
AdLfdCBhPsSBZz1OLBWT993BmVf83/KAA60/Hg0ere6cj+0beMdcDna2EUbVlz+4
ro+qKsiELgJ3zeKnnYVTo8pywtyBUYejrZwXPHcCwCM2SNTkgzFY+XZovfLlW9na
haTK7GTtoCQJJlZz8A476wKnrtbHpZGmeE3Z6YMUZ9jxQdbVpYJCgVJdx+OTcp9d
6b9Q78STuLJG6A6kYxsaJjAfRz2F7jQOeSwdRmv8mYujPcOBy1igZOShHCLT/v1C
V6ifaWUKU+n/+CX3LbvOvcqmK9yM2bjwlfdNObsT9lsDwN+NSykzF43hFx1B/uF3
R93vgMH1ATYbaHEJkSZLSliN8cz9wxjVVW4fmsycAeY6ph5cnY7YpWTcopHjhynz
s1EstiVwfryrdybEp4YEhgE/K62koi70KQHxByffyBiWOeSTKtI51HYCIGtj+uFk
XDOFVRZacZdQjZ9ZrBXrd7LXBdsdN2BpNQK8dM8XACQ3hBN6SCPvpaA4Onn7PCO0
6bS3kfrpKjGjPgwxHWZqa/GANQaA/NsM0VNyGuKcqZkmE3ZrYiG9P9SPqu6oHhRa
1UuOdlMZnFKjJsYR9BrtSG1ICqErF5Mfw4xwMMBSbinxT5hrlOn8Vtq3CR6XKhrL
7r7rZzlDxMMPpG9e2ODn8rD7RghJzOF4zgKW81y9bUkUhJIzGll1VwVVeCHPjlWm
N+keco0CDaTpCiZCQlr94izpJaZUa/N5IqVOP3Dhd2TJVsO4NvqOiuVs6Bnxs3UN
XPUpnvy4xs5egoY43yVRYZI6au8go4SBr2wDaBL5EBewuIomLJab7W2Kn+manV2s
k5dQFxrChuU3yirzQQoGTiCU4u7TBUtDcumLrP5cMn3v7xJUik7IZHXcYaADuE/7
SNZLNhiMra5NZ4hoT9y0VfUS+++/Ori3876ADp2tlqzflqdV8HKwUKhC0wskYCKQ
L+10Ln/39PAW0s9p1NhdlJ6RuA1RhkSO52U27sAfE4RYTRBE8TZgUDX9q/N9hYW0
1TtQ+1BnQxGiVfCQgigqHrDVciBQwNZnF/2XUmM9Z40PiouITdqVVDQgYOodu+ts
Cw/NVLanENJddY66HYeOAkEFfqAM7kueIgzJwWMw5Sf6eifWfIclUsv5+raVgfB9
DqsPSMwJ1ocfKrP/2K3ziTP5MFGjEUDBVEqa77ImPbEoVJ3NCKrx+WXvOkApkKVp
1c6aq1XLEJ5G3TGA37kuMG16Ri2q7UbmZYp53Ffo6+xEPzyHznwG0EhOjAz/9dQo
Jt2hq/4bsRponH4PtUERjs02Vq4yyQ7gF4B/8SVWvZil3sFB8ENOgLMpwQ+B/Eee
cBfUjQttj1VE8A5soLs8R/GcTRR031/JY5ss0DnMLjhyHKuBFc7nz89I6T5Vxnhi
rskJiCdwzyOlciYoUVdJJryyjqG9urSFEzo+2blmMbdMbTY2oCRJQPLVMcQfHH0h
eoeBIPqf0/j2/QlvZlOIMYAC/0MDKJ9t7Vpdje5mZVDQd3fuVi4HcG5hZlAzzsRg
xnGWhY3m7jUnsebPYIe86P16FJsDt2oLKmqeu8uKvxysDeZyc2uAs0SAtd3KUhRW
pPQs63xPgiVDDgrNBFkJ7bJaURqWcNMTdmd+DBKLqvgdHR3DRtU1Fu/GIP0jAuA+
woF7HKWodnzSePusbvAQYBgEKUE/tCqfnT+YN6uFtml4fLoELcaJMtvTE+X68/Df
e+VQzytn2u8rto73tteAap8tU4J4GEUHQk0XgadsHeyo6v2ol2RAlrZberATGJ32
nZ9Eaoe9xCY0wSNpSgrY8RqRYFEKhnO/qUMCFQylUm1/6FEMmmNnHmcQIZzpBluk
geaaDQ8Nxq34zkDE4qs/BZMZ6YdnesDVSyFStHzxmyCDwlctz9vEwk5Ls1cyiGiZ
VfZD95rmdjpTVQ+lTS78nPgtVnvjZZFABApnaEJbJrwU7yt/jA+7rRRImqMkmG+Y
GJbapRNkBMoA5O3ah/aAmFxMtO0cmBg8OOVVtyZJdqzzyzGDtUT2TWcyIaPLEtag
w9RhBz4wS9YjFsn9x5NoUbGjK/XuhCrqBoYOsflPwg+nizHuHUD3cP2tEgnk/XcN
Juz0rF5dPumDZmzyBA6Hpiwn4c7c4WTYmOKvSTGadUFIWvNKurF1bbba4VsF+dHr
giVX/XnLsKCrkloyPnWg+QtbwjdHRehFVnG2yxSbMBK525GBiD1ct69ZQcH8bgA5
Hy1DvEOqoU12n0RRhZz093MwgkBbz1Vk549jNItRvYLJAihtr2Xk1PvnKkXal18L
4dUOxj7iIQdjWzSwW04uF7hCkeBXAefRSPid1bpp6+oZ9BMMG8oGcBSBRt3JBZSt
BiUZGQ6AE5zO6bmotx3If7gjX0fdGcjGkv1pDKdh+R9a6/wgrJzovPauj9dVluf9
PAKBZF9kfB/xxjhJaZjS8WW8LFj8lQc4GyUn0F4MjiJaTuTuMIMvzQYMNCzbwwSI
4ysOSnpXcUvwhn+PdSkPzxxpS4PZoHhDwN+A8ZWBA1y+bbRBLMUlkwv8fFDag/yN
0vBDJ4jl+ZW00xQcAnDOsISO2F+IZjNadCZEZxm6kF3MS8AYF6H/w6Fzgr6X1zPy
nC4oxrkXkML2NFEVF6bgq3tg24c8YYp9X1943sg4xhO6rmEloliWT9cmgyToZE6a
Ed0jrimKZddHZM25rK7z/IvEqIe5EIpjNsBotsHkOBeVD52dE5Op+0wVpV/E/Q/t
9NvQ31Vp5wmmfPX/c1iJswNoD31bxQOkO7AxI67wBKyyLwVM3DCeTtVUpLk8SoiU
fTgCXE34fkRKn7Gy5qJBPSwb0zf/VTojxElP4hmFRdwQar2RJZ6thH0XafJRjlTD
rFIgPGl2UjyMWYV82I6XqYwnNkmJdT0IaglQ15rUHjAJBZs5bnu7sX4ZnrNEX7GA
05M67sSKvQOKWxwHMXElYT57QsxpgwbfSamPzs3ks3Kv/M8TsNfvwvGSrl85z14A
vpScIM856QwFWWaO+6Q7jzBE1y8lGm1LoBes9yPiOgHDwq9OC6YCAeDgtx6rjq4t
C7juc38VzSwpRF5R2v1cpDvRICBxGtSEnzJTMt/+y4Ho3dt8MlVLXyd0d1n4o5mR
zEb5wOP75T0X9qG6cIIT3FPAnxjYPCTelJJWd5+wl9SKY607oacvXDQehsy2UB52
v5fioZnZrFdn8fwAxeZy3qspV0ev8IudKYRdKDF3ZYeIs0JXnjFaN86w1o89e9YV
cw8girssqZxi+6t//c0MY92rZtvzw0mIyhb+03qLP+s3dP5aISWtDnOaGRTXNMDG
Pc+OstLfxTs6uNiPxUSIH5OT/BYrfrBjTe1KLj2beWEUqsUqs4tlRPoh+2DWuk5O
65Kh5CpkMi8C6w65EHrKbk/VAB6OeSBj6zoC3qDsmFGRd1C7pM0DQ/XGXD4+vz/A
/lEx5jukqOSOTY2kPQ1n76Tr6ZcEvU12oRJoMVDitSeLQVRawiAQucideTfewMAE
TjAwETSqGD/KRnOESPo/QIWFAnF0xgSC/CCmFecjNCs55k6pUR/C9N2CVUvhKfWK
p+XclrsORwT0L9dKB+Wb+PS22AGapCBg1vYgeOgJrLw43N9eXfqhIBp/gYF4vWPt
Bc4Knbi8u5c0U0myLhioARmHKg/JfGZ9dtvhyME8YYko+Mlb0f/jiCuIu7piwqRa
P2IfPT6JJny6ldMMCeJb+jMK7m4DF6qbxAeFaI3DxFtIHn4aEZE86T7IVaB7jrTD
1ZYokaKqot8YpWdk17qryXMziZ5zsC8qjGKfaffEhhjLXviYp1s6wsIYofovSrUi
9ojF6pTm/A2pl+As9x0eZcyTvPCzUAX4WEeWxR59hqeeDS5YMAnbHoO3IQC66t00
pGbyKwnkXR1Q94qrRGOoK7fN9PTyJMN2HzBLWfAlGAdZatIftfeMN0V3tujyr69k
fm5M10YHCQMip5nPSXNi053i9yeCpydbVpqtQdqnrWhUZu3HLrce8Xvtf/85fIe+
spMipPpXYLqGUmx5kC1YAuFASnOJHV/ZuiG1ghyt4NtG4VwrbCzeNb5cj/WVrCby
ZSGJzoauSBekg0QGYpVcwB9C48NpaxG7CloHPYO8XBsM/buXz1lx6jSS/eFtSMsk
sOEvky4ozCrqviaEwRYBoDXPh46fNdEsj/c2G1NUuYuYYapsukAyjqsggMV5JtIP
7Mq/wenl0ihLOPOPWNtu+o/MKx2kOc+sOz4NgmQ2au2BYgSOBLtK+WC3toDkRH2d
rXNG04T0ygGI3dkj0U5TxCcvY7mZkIlYKjl+kQojNvNuhVhhaXOtCDRp1OvfsNyS
IbZ5eWL7u4uCEstfhzxSEZUGqs79vzIy71TGuJGMcW/7I/agTf2RNMfzoV4E44ly
YT3DtjwKxktCozhmW51UCieILBiun5ZmxtN5Gv9AetXIQ3qPsqSqHZ1OsqHMrG3n
rf03A25Gz3dM1H64volblFCReya1x33bQS5Ylf5AMemQDlizhGFNUTP/LMAIrjw8
rPJcj6BLOvfTsHsH7Pcq5mBj1r//g98Z/xx58ekn20GlIRhPcbhlE8PQ8TMUJHZC
KzVfaasz3sHhppDjI6CA8/mUtuUzqQubui1w5FrOm3upxNsTbQoCfiqDWQ4Q+T0J
6HoK3yFfp8c189Un0mPwJ1XWXoG28DOE99U69hN0giyjJeFxe+iZx4+24I0nOiq2
OhXTzatR8DUr0BGFlDDWfsdUJmIIpcKueWH13ZD+sMSbonpZFn8FiqUbSAtaoXn8
FzExVxBMEzwOQlEh2X1JtN7172ENDPg5mJzfw5yd6kNSHP7sneNTzlBztAOxHHPB
jYTaqEY81YL1ozUVN/wQFPpPHgse647UxmNAX3YNnhDM+4hJ1MwikCJPF8YRtaTE
gABxh2UOFHeZe2kSZxG8ekHAZyFi7GwiYxyTAw/R8N8TlN5F9EAgVn4MBFZ6M0YL
gFTa990P5/AbNYjvnXWSmc7EjA3klHbzy5EhViN9ct2fQh4vm4myTiglfVxQfuC3
6+372004jHfkUyWSEYHNNRw3p8cATRrnn8F55IWv+oXynndP/Htinaeblkxd++dq
FKkP0Hc82FZAl9jnLSr1sqyYCm0XVzYZIBQDEZB2dBkOWeWlr761Cm1+AkDODtZV
RbLc8pEmLCjHMPUbU+p5Af/EL4WaFpEbvxCcgyf2gaj4EUO9EmY3uD68SAdJRgl+
mMeGPR5sUrCqQ18wZjEQF15NEZFtrXTWP+aXbvgcXB00nJ30RuTiiqznMoTCGzhU
R6SnZBhpijzqIBOD0/kVcMLAzktbiwdqLfBNkDPpd7KCQPInnIdKyJNF0nl+/EMh
qfPqYLTSaRCOLhCl92PQ7Iw0M+U2oDk8GsdcYpbpWqYZZt3/gGlVhQ24Foj1BpUW
et7M5qmBgD/Xd3sf2e2V/1cRVfhJnhYU/soqETZ6sohjEV6J1X6kdI6PMnOZV9R+
TM+VoJpq7b7zbZ+rB/6YdT8ebE/6MxHTblRKl9BjM3fWorEQq+WyFuKvVP0Omo4l
FzYRq9FOqhCE5PX3x6PeYU6uUyJ/5HxF9rG5X4ggSdQgqMLk/slu0fvHWly3CB/L
/PerIB9RL3+9/sqySufre9adif5Wl3uTX///+ZIBKOecjVXYBqnor+e3sRZP3+lu
A3Y72a3XEnlsjFBwBWFjzMGVTdg6NO1l37xIGdr3B62Ur25JRi/rpvRl/zJugjL0
iLBfgngGaW4klcUEwIZVHCERelGApj/qA0gMvNF/xjvVVRA3w/0pPuMKlQi4HI0b
SmSggshB/NXoASvUbWTe4i3qU+4QH/XlkzubLYJHZI3hxBi83Z9rGicU44xFrfK/
LtWp8Ot2hRfo4GaR3gsRW13l+KmQv1dx/oMQU+8bNLZ7PHL81tL60wVarLgm5zWv
cJos+szSpBnuU8JNf+IwuA22NC1GfPJG28VydC455x+cCbSK0i7YpIA64SnHk3sk
kx+24ndxayATAvf0+tMo4dN59ECKsRDVi74MBGkZcJQ5WaQSfJVWVAASdjsl1dtz
wlW2I2mlqwzNiFLdDA4reTpssEKmPMBL8iHXUGH+hWfxGgWfXBlm71NdBQu3VuXF
XrjpXLZmXXLsYVVrzFcEsbP5Dyv3wD/m29lmyYPRo2XzFJojy80+tABCJLoq4HJF
ZmD4pDdkgI3dkPDhEYo4Y570eQG7lTWWmz6V/pDP4XLjfaHzkoF0jUVyA53xw6qk
nh/FI5nsnGzpT4PcrwCdHotgeFsCfBE8w0TWuXs6fQosb6/jMeAsmDansorvnnEw
PX+Z3fQC2+76ixOqKAX4x7d+hyB9iCewtdkKe4h/+dNdTyJ8BH1qgdCUuL1AiJ5Z
L7gzM+TeD3CAbGpMYpxC4kvkd+aDYASubK0aHWyiVCCEPWi3dmXIkTkcOfZWWnd2
+sYFSwlCMVj1Iu9fe3f/rtdYcM0rYt/elaRranXyJ814IwWalVk3kjl/VQBbjKKh
iNnQG4VGPPXEE6OJ3SV7ymcZbw/qc4oLWX2EMGHnahXngE1052D6L9Wrco8qQacc
HFQAt6ZXQ9qSE+0/zdZK9BP/uIXS4RVyY2Rt7mPvH4NYgZ9Rip7G/vTHiAxNRAJJ
rUP+ToExVDNtuxddYnqIJAgIkUlmtTBSehV2pv2pX/nZdWR8P2e2JTAgncL/Z1am
ZGmEPM2pzxXZf94J8A7K3R4bBSb4aGwu1+KGndzNunlVBjqOC7OHgm8KF6FbQkRM
GQh99ipxhmFGkdY2pI+gHu7nvQ1GXEcIhODPpvNJ5hsIFope6YH9s80QJs2xwrIJ
hD4gDQwfAV7xwTZT6pIJ60icztJDDVW1yxvouvgVg5A6oBkz2nX2x+8b40jgKn71
KUEkTt9J7MEzZl0/SGekW5xRAaW/Hxmq3ywqwj1FnQLtXnuZkSykiuAUROecsARU
XnQwRFtE8F30d4kju2nEvs8coiLDBBBIbEIfrsQgodqUNdH0CVJ1Xmc23r0nHQvg
XSv4XZrY39ZVIjlmIuy2EIzii6tw5FYDGDKnod2lEgajYSVxs6MIaJz9Be1UKM0H
fLfIEDAGPUoL9JXzh+y1b4iz5O9vHSjcS7W1a2tEwbYf/h1yb4LN9YK4jai71r83
JhpR+DlovnALHDxDQ7xvPr9PXcf3sFdWZw0Y2WUOMeLRKg5wV6pWdEZUVfDP0U00
2xJ+0covmTP42dWpV1aYbPXAgcI7W6PnaUou9vWjW+ZOyR7ARGdtevGi6w8MjP9K
205lHXZm2+oXZmX0SMwnfyp6oDOEvp6uHknTbsTTIaMN4t34CMponbClHnUetOwv
mB5b/3sh4cZEoSyhbHVFgSbMIJ2u9d/Ieq9MIDUw/3bBPwsPHkFewUP9lcMcrFR2
q4gFUAT/RD/e2USL9cpsHxmqkB0G6/IBghDEY09XtvEyBZicgP/VSVQIUSJvWuCk
lLsV8KehxWvqRWtdOCxW3rM5socNheeDXmX+UX2PFeyXdVUgEfDXJFIpQAwZEk2U
tFEH6+kgIsTfCKdOTPGT/SYpdYm860mbumA8I3gjihL1b/kEfuA8nX2HQjN9w4LR
ScjqdfNp5Q+8HbliRtgDoWbyW4gmJo7vqhtPkrIvw3ftEw1KN6FZyFaAwh3wUhnL
PrAleCi7of+YGVYjVhXisSERYlrzCsLYkMZUnfeliR9RI5WK1wsOC/4kV3Qmfbs8
yp5zAXFhr2S55rXU0tlRcIJpysxtjDufzZHVCnlggzXKV/iqq0Y9WfDnch9P4JNg
Z0zksnT37Ep1+k31Nw7EPgp8Fsh6hNc2wUy50h3zn3h1KSRZG4yzGK0UVwggbUpx
u3gIcdfReVM/a53FIGFZqX9YFfpnRoOcMGWx8YQUE3ebeC7hO1+6f528mMbMoYq7
iwaWe82zEYKOJkp8ST+NnGpXDUkyIBNW+GovBfJPg4a6C9gBuqdOpu0/tkzlKMIL
qQw1ye5+JXX9m/Az2zZ4wKoRphmxP8+owCNK02HwQJcy91l4GGgeI8d1snh5dZC4
8FjKpATT+DBvPZ8bjFBNBoK+xdkELxRuqQdPBC6ADRecKlSORCe4s5dV4FjjkRP5
DfyT6PbEZvK0nZnvfAi6xgrmp78e1MPx/dtBC3cicaks6++sIUH6LPZz3EsK6pzj
cPjpWwsIiploihIMzK4h48MCThkO6+RZPFkrP+1yufsm1Phf5c82NXBXRp0F3Pz0
/J0OgaH1HfYQ53ByeI+piW8go63FczOzwrJX6j8Je/krHpQhWHZnLvma28dEsfV8
El/TE5MerUG2ZSkOLb66Qrs0UhKsL3pjarcC5HVtk23J8E/6tmkVQHF0IDPA2/FK
9RRlPuwg2CfBKgpmVi06ipnRcBITfMvkOCGA+nmbUhxXcN6UkHC7k3HVTfmoGYzW
StLvtro/eheM1GwacVYA1n5Oo1dF48RgMfKUmjss220g71LsU7bb6YRhYxT7rPrL
/NeCAldOOuq2zIvnRB6GIXPSl1JTa5KZiavCvvyQONhm/oGxh0YyY+O3Q+mlpO6t
btcgK1CjjSqg9wuvKzunkGs166OvD5gkSQSaZQRRaENcqo9JGyaJEqx8UmcZ5EBH
iruzq56yfrTldMqoeI657iD0eKcWLVK6uLoILM+T9agzmwdV/fDW3KmCwKpusFG4
oSSDhEdU/yrBdcMigEXePoDmNQHLaqVodyEKusYO6VlqI6gDei5QrOtZm5CXs4N/
LSej5W+iU4QsFcNnR2FVLQoUSLWsIxgBlInIfGMDram7Ls1wHbP9RXKRwUGWzmk9
DsN6ygGzxHCcjB3JhcMK+RBdlxfKdmINe0M4bhtdHHaptk+p0+dc41ZhOgi4yj7X
k5V7NrBg4YFwy/jAjGjahgENesmI0Y8lO0fzt7j3Rq8VvRyd0h3xcIOgjQLvMk5i
H2rX1VYm2g7AQjwDXwam/lBu/A2P9fTIImwUdHczd81zmEuCg0ec26zq231q5knH
l78omaB/ULhLX2JLTJ4opH56Ex/KTgkveTWSuYZ2yupdlCizr/suRTj/DTdphkDY
lXeeKYCTm3FkxlPLvg2WXH6R+CaGDPozzvnph1jskHGx1m4Nn1FeA7/AQCgzLrjo
sXCnoi7hIhc1rpF9HuNrg8sY2L+g/yE1dVe3uXQOMYsYloOahJwle0wKoFOW0unS
J1p2qsSVVPza6wAklNFLfsL8cOb5NpnT6/32tL/7XoJ+TSV92/shvWE7CRpmQoZR
XAqzFtcUxQ7Ep/KJdpFzwfxk74TcrDw6p43q9bOVpjbiBk6/F8cPzxIzjeHLOJZ3
BprHbVoqZMfEMTgRfxwHapr858p4krS5SLOHwJHw11c+I0hmdNbvKTXwB+Tcivq1
TgvfM2oNZIXUcipR5dGAvcCzmAay/VYHmhCHy0NOAypqvX9kj0VqvIuFHuoTOcEp
hxk2BmJ+JCl5Tl7fwfznAdb17YuZ/X1hPldMzivnIWBeWByuYHsPhSOD22/1GRWq
ZADgTS1SKh/OHWabIGufZxebtUrm1ehikkyr10zm9TpUMoHHG+WwEwB7JTn1Xo0r
s2RDAv63gkfaLN2uuHDd7/4F5s6krNjPlhq8BsXurtNLrX82W9JBW3pnE9Jgbi9m
Nkf0253KUjptnF1Zf22JOUUoOVw00xeziarfEJnF4y7adDmqLKH8gjKbmPS2xbdT
HAASxWUoUuX6uEa+nj/thLhVWp2vUfd26I9Xvt8/hc5Ao/fKbAljL6H9PfGqqYft
+9QU07lTGzrNUJm6ds/nkqxRxgDbXxSzTqNa+elid7ss6IH2H3d6RMtFpdMZbAg2
9Bw2w5OYVwK7G/WLuJNsBoOwSjdYwhKZF7ne5iZmheIDvbd4bQSr2cscL53zjxjm
lSM3/bt1JFIkWHHd+C2H7Xiz37W9h9dOpWdK79X1rBKfBoY5t3pNXwYbG0h2OIj8
4GrW4P14UWESmGCJJ7PC05gBbuxzPlASoWWG/wanaxfAaOhd4uauyKYvqeVb2dOX
8QuhDfP24OCp64juwp+Mb/551b9oJ86S32iFrVKQu6nJCCIdv6iIqV9E2exNEql7
0iBT4n8nkgv5SbfD8b36M+DbQ92GLljkdURGXMPMBwCDHY0mvGtdAhOUwPVs5/rG
umBQD6iWj+aSOhIK575LTD3CkqrpNSUe6h/TmcmGqtCngxtIxnWdlsZ52V4IcKT0
96yh8KHUgfGRpLiOq6uxq5izoytZvAeahrnjikl7LU8EMwej+0740yvFKn6Uvnqu
gRNL31JeF0gsXyeCKIqe+yV8faUpl8H4xkyoKd2gQaSq/Y9NompIB2CrvBhf2TxM
9/eORVLAMVE8SDN3x0zNqX+JW32ZlOGHmStokfQSdXyGw2MhdZO1PR/dP4EC1R1p
lPLLXeLqG3t4Mr7tdpc9Q8F37wQcEi/5jqRYD4SbtXvrD1IJl7U9E3Xcs31X3E6b
IZURFbLL3tIxnCZeBcuLuMuiqs6qWQRsZUoVp+CklsDOfxzJf745JcUbOsI2QPPs
A1ku1LKRJTbzDgE0ZLK0pWLXC0Qb4MFxjdtPWZOiV8MylTzcvaokPEUG6MQAIHBT
F4af0ih6TWQc8oJOPD6YpzWfl0iqkebwCICNJE3WUFizcc/F1IUYzzyLldMQqV2d
NjgoZTITXlcJ0DC+knaGh0Mvkluu7aBRdUehaq6LHPds0BYu4n+7vwckenkLB5FB
281A9eqHdoTw3uxOYNZNwJ/GF+k+l7LbqNFGCD7natUZK8MpaqYTwf6U+uEWn83R
9Jg4Ma+z5PjTKSdf4sdSoUuyNraINSqZEb4lpVmubXiptMGegZroOnaO42W8m8fc
IVvpgQ1G5Zcd0FwVnwxjhMpEYifTkWh85zgKG2vfo3UXNlJAsWqJz0s4BBLJcclU
UBwzFLr5Ciy4gs0ZwsR01KZrogN+s5Pv8j3Vi1LiO09W79Qdz0PtHgGMHfSuUKWN
eTxlw0rY8aVjly3I15S28sc8gDqfd5euoyYlG26AcYKfETsHxUX0yTeQ5DLNa+j1
t0IkXaRmWR752LiZt+Gb2PUWpwQV1DHccKKKb8e6HwI=
`pragma protect end_protected
