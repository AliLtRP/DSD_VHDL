// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bXHdILr+4S6aFznZSq1xdKhWg3JTyfcBQe92oI3nPS3ntPZXZruIqWVDjVBpd9lH
UZlxV40J+sIyNp6J984jJCSQFpX2ruYiBerTMtCPQkO2WvYGG6l2o8uUEh59XLTB
W66fT8TRK6llSixFeDYVSkW1FxhamZDhpeBM+Ue6e2U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34000)
/2dPwOW7teT9RArkRX33yNZHq+x8dVRj5jmjkQkCzh3LwsfAcJRQKxj/YNIfbiMa
x8TtKvPqejcIVTdXaBFFxtApMYy/NBEHZjybfw2FMtXnwktgOkz5/C/PteH/BqF1
/bdXoF405K5tJOou2y04WsqTa3xa3OPoCt7h5U+B6WTFBLxgrh6QyxnHBBp1B/sU
sMB/PnXmoqVcjI3+8Skor/ZkEJCsg/et7LOXlhChDeYAm1yqdUh6v6OOedE9N2ko
U71a/dqkHUqcId6fJtqepWmL4O7auS7B8DZeSsnkzjbosSP509Z/NqjWzELsdVOI
02cujirRvp2s/WoNjdpS5inowa581Y9yzsC53E89CYaJRgSNLs9vPU0rQHHPMpyY
bBDd7d54Yw0tAxvqyv5wQlslHOmBlZiQBIHySAfqAVWlC4lju6eb3iPqHZvhLEUb
6KdA94ZtEFzNp6N7lprGw4BnPgWSeZ/cPqN/16IQ4L+J7CY4LuWzXvp/1H64UAmE
hYwi6Snxh3IV1F08bQiOIWOWy3+mJIRDfmlR1Z3LXUjrg+NHLuUym5RInwj8DM+/
uj+DH6dY8ZApwLUTvKy3nUw8LZqIkfg2DEIQRaRFGL4mMO3eF9ElAjA5ld5i3GCT
mAjQBhwmFZ05ncwzOS2/qLxFzQIZqQ50Q7znQUW7iTN64UvHE25z05mhLKV+E7Pk
rLKa7jyMbl6V46igQZ6oQYGaNKCXq8h/iYk849iujas3j5Msuaaiaf0WUgmBSR5E
tqnn5XCt836RiTLvr2MYL17/Zizv5j3b7w8OcLnjKUBUnoK8fsQl8PkTqTfPDMug
UXqfVRd4g6Naq2D3X1vHz3KUiOBrxSfv+aATHBDo+YYIlnoPka3QNlyT++PuNpoo
BX+r6XC9JMe9eAUgTwgplDUtiqjMtnyse+XDBL28dQelgHTDx5MxRNRguwL8fkQp
b+4XYqR44kyOuBoL0kr8VEotxfLDy/6aSJjD3M5Hc7VQRVD5gmjau9bpOQ9Kp18Z
DsPG2b4dPeRGHUdSWFxUAnrqKC7r+SMRfuT0kDWwwQlptQgEgL0BlaZHlap0pfPr
FNzApZFvshi2SnEo6ufEbRmiRA3wVTjLWcnsqwSOYoS6eszG5xI2gqoO1kp9dP+8
K28NtEepxBqCqGUnRZoAQt4AuJvIpSvq6ILbTrpKeziqhhNV6T/1E0LMWD2oVbNh
1MyKgAWuLc2yzLoV7n6czFVXm5sGUyzxYpNiOzlN6b9TYZIP15/dhVLyQ0B2vBmx
40DwC09xGDjtfNDb0pSjoZo/GwK4DXRrh9QgOY/41/X6giU5cxWW+3uUHvQxH/5Z
RXy5ugMTGn0E9Z0faaW+Hz5n+RlZozZUIkqNRr/sqr+pdpJyJ7J5xzQjneG4xDDO
dZnSIwE0HGgsZ2sWL6UMezgxI+ai9Q2my2BLBufljZWStYW7Yntaga8BOEWyxN6B
y6MbOMW8YcqqPcwC8DtfQuH+4Kk+k/WRlFZir0iM0onqWEsiPYorNYZHZMgdV3Rq
Zf7JSzWyKVKYJT7o5aTJXXzxVMzsOtkRd2RmDfz9K/HN4+5fLI7nkK5bLMZXyBin
PmVgWA33vbepBTTxpGimqdcqTBJa+enKViWMq4LrBDyyc8Jt7tax4B6oY3RSgtSH
8+0sssDXtPF+LDoAhUHmXLkRunVYZjK4h7FgnaBqMduSQ8rCmMV0ZH2kJwL7c2DJ
vNQBY6XxIq4A0Hr++dvkZGtJE+CrrGuN9mBXWImvojGu5On95+HLI998/i1qIwWW
Y5N1uo2IAAT62yUYIGblxW6VxvxbdNp1BSZs3BuCM1zPCuom1gPPBP8qXj24uMSQ
C3O6REDdLB8OpnPZ1piQ4wOSFovxdIVQ/q6lWgUg5PUre1MXXcRLEZHa4OuT31FK
tkI6H8kzZ5VRjpZduWrynYL8fPUHC4ImqB92Wkz8V/Xq0ZWSiL6t5awHKiLoKnQP
HXBw7aDWJsrQot6dUID5b8mnE9ziufeFFNX10MsMucTNAEBuUxO+bxyIYVNRoIJ6
MjCw30jDvamFH4AjvbzXTuBDtP7VonLFhrmjBXUIETsOufZxTiEnHzxsXcMJzscV
dgknnGA+4k4EXg3lEJ/EjR21ICQhDt4RiZUpE0ZHDq/d09+GnsD286ieLAashPgR
8LlH4hlgD18mFCQdngpcI074BStjmjNzJSjMvykZywdT/wjiy+sGUIC1+dMadmb7
+bQK5eV3F0O0nyQ1IdalvwwEkMecJsbtqDAiu6WsZMS7CNDH8t5Bt9IqKx9BxBxm
zb+xeHBijoGkLaKF3YfrhILrNOpVm0oecv/5ngu2UFRzRNjnEnKp85ro9r1KR7OV
iaj5fI6oF2ikJjdteBZWZ2+AifjZ/4JlEIw3FH2XYwhkafw+PDFQ/+fGSVh6+Wom
a/fY2OSynEg9bfduwO4yTIQ8n7bgMxnXEmFpjvdhTQxAInSgPDVGzCbU8lqqnqbf
+CwYlgb1tZE9HMUPb7jxgUyYRaovLq5TI88pcBkWdqHB5SzzndwMaIcms/pRics3
Kj3AGJzxrrZIpHfE68DCsjjMGXdCyMg0N0EJF1P7SP0w0KQQxZmm/18s7iF1Qzd6
STyNDvJw3Vs8GhunRT69ctF5lfLdc2yn8Iteot2fiEF8zcYvpWqU2gkGtUp/iwNL
ou+G/3WrhCi8QVllg7rYX0/9AZDjjLRWFLd1mvF1OjFrn4+8sE06BajJTGiRZR8t
l0WxYp+m4LKLngDonx/RxC/K/L31XJvqLC1LKljkKspQoGjUazK3W+1vVX3lkOPx
HmKdoXAu1nGIYMvLr8JF7SMBlDmMl91zQOJyGsXYBcWf3VDaHMIIW4zfyFt0bR4/
NGidFrqjxvn9SxpjmYlAVn6CxykrJw1DgNEe4gP2WihQElkTOVEmXhyTJROxeVEP
hibakYhK0DJA6Ko0aoLktz0tbQzvyml41WxUs5bCO5fGoMtyDbOWyngU6vuUrXGl
uSarS1yXJamSFyWrAccVwoinPWlJhXBJCoDRQRQEqT9ofVDEgCIAZ6GZVQ0XVWIY
xGJRijyeJ+t6R6FZ6CKom4nTTWF66h1dFMATz3hw0PUa4FGVWtAxMoczHVNvR5bN
E3YPwLKpVvCYu1Xcj4lm/2JdVbsLM7I0V9WBxNcTHZ6ggGpqHRzhaY3W54evpgbv
TQkmCPsxvYWj8aPS8tpeo812a3dQOM2pcwG1hrSTQfi7+EKX7xm3ax/imnrwr+ky
o3nx5kpMuTl63Wx8sT4g6jkrxtyjScdzCujEHk1S6O2/b4fdNC29jqbZW0plbMCn
DJNDgybUzWo8BLXfloXrJTloYTn2B43r+0lBWSwjoojWbQtd4QIOWrSkwo2r+Sz4
IywPsIM6i5UolwsN+IecXTZ9y4fFvLo2XMTO0kyaxDOoZM+k138JvgoeJnyJrrf6
nroSLKiaqOD8/HdzCCPjr6YI6xAyXgGHw6nhWtvtidrTokkuqDiWFTH+7RR9vrt5
hEDc9Xz546MXRXuSc4TPX6WKCZ4+ELG6Ojb3jYSC2uJiJAZNaK3EyAg4XyPY0rv9
0sSsEFyA6BmnD+CE0YAqe4UwG21vd4qfWaE7FJ8tU5/twOdx/DQLOSaHw7qq7/7a
kCaFcpk4LkeANqTFklsNbhVoVaiwYPkPs/jPHDmHq60DgTTsjQUBEe+Fq+hRIuis
T07NpqNdsbZW3pok8bpSEluF2phtYX8Ynx5mlEBnS0FenGPQ+xC58C+mF+YieYCf
mUDef8ISK0rWRaNZX/h84d/XwZYa0duC8vLlt10Oajm/ynCBYsjh+0nQhSv8YOl4
Wekn8ylN1SKVTD9wG9QDz93rIuvCVFcO7F59qsXj9T3Qndej/qkUpF0cSRRHbcnZ
Yah0MIO58CB0XC8XPqMgCA2PJEH8yJlTAi2sGfOYt6X9pF0ZzgEohj9tTGRhBbY5
Ctp0smPwFMAqa3CxyKRKYjDq2AGc0Ey+WfZ1RKGz92oZGJzSuvc6oEnkaey4JBTH
wgmT5EMaaUGWD9DCCZjxqdqEcy/bvyK7f7k6w1eAkmaZI7etXSKsEONzxUIuXTdq
xR0jFIBetpRMGeMlj6dIgqB03FfXk+eJZqyMsoneMFtZRzJU9FAmw2htMp1L6yPS
0MxlyZWivpigfvdaUhXsXeFiYCEuuWuYQDkZ9yGPArqTCUfGit86ikr7fO/E6MEB
lImgkx9XwnCOSRhucPmDPvlDx/noHDOehVwcotJdNgvVgPkSuCvKvtcP5eD+UyEI
MlHxMqQCmT+4Kp214jk1kdW3WKIEH05VCod8cVER+Ep890/3ma7YFqp55kJwJ0n+
OkB/sVRHUgJAzwAQrAJPu2tylE0bub/pMD5Y+z2xZWeLm6c1K6F7dMKG5Q6ALxzV
AS6Wd6MP+VMs6hwPbTaqOZm56NEtQO7FJNisWYUH8BV7E8J0G/GsxnmJrdcq0DhH
2AZpBEPhXGwTFQUgEPjmGrHG6OHnNhtEgKaTFR5Wf134S6Mbw3jLqsAKbMPu5OJw
c9liFSHutABcPgEKkgiqOxygkdsYkwU8YcAnut1LMVNRwAakFN2uxRGSyYi2D0df
pcbHC2jqWgvVkfqGspHR7kkXpiB883w2LlkUqQDUGWWkighoDFn1h86ZWzPxbP8t
6kp6MSxcJjcfVx/sU/tdkKXqRyLeWqk30OM8KSy9xDSHrLyTJtkc9LDvTHLSAae6
u2hmyLqi2NQkdPwn7T+BAcmJWro92s7ARz6F/KDs2FEMN7VdKdO6a5h8k+oYg/eo
aZFh+9QVYh8zmqc54xSf2DWzVU9rPfTZMcR2d7hqi3F5ITyV9511STSZDjyvLssL
zac6jXo6HfvwRGI3IJnLubBep66Xt5FFWaWsRX8SC7nFNOCDPZHGnD4jWNm4DmFW
+KDfV2qMzM3vyCzKcfrStfJMjhGIclC4Xx0m/HPigApH0kn/0vVv9c6zbJ2Vzruj
1W0ijVUXIDBYKIVusqD32b7w5MIctM0P38C3JNLNse40+PS5JRmWfL9TUVWAXGuU
WUuguFrz0n4Eay/tKw90yB4BDfrpRNbTSZgyPzQkErNKr6rnMIy0pUwxjF/Dn6is
M0vMAA9lraj/hksApe0QZ/PgAiIoE1mRRVpptMt6tbH2WOVIrwvGQxATkljSyoHx
zI40HtqAkZxi6SAkOW+neRjnxiuRrPysIFj8lqUklERLrUsZPJiABFZpGAPiFrF2
xPkeKjdYrsFtCL8h26buXEZrw6jImXkABcQnHXf4pJDIy+IW9pYu5Q8eCxyAIh0X
n+PQVa+jJzGl6fHIzNyFAZRHI7+iAQ72Zr1pvBmGUeoYgJO0P3xD8drzx6X8LPte
AYLV0CsCpn0IeKQEX74f5TkdZOSGAt4GNdmx1r64IHP6rDrikhBvz9hqZIiEwLhW
Jw6ZWZWe8WmTJkAFL0I4t4J2joWH7bkHcSn1oF2LUok4V9Y+T2zQYcBxC0gnXKvY
BQl0PuZrEzKCCUNpPVudjiJ3MQwn7LWqLS1BgfZZUn2zPCLXPFcftZXtblyulcx4
gRnmPim7K66NpIowswZQCgoSuCM6daRv5xS1N/vLGSJxy/TeAb+etOZTsh4+Jmy0
Cs/PWjkWyOoQKrlXIO59AqwtPgH84wNChFSX2s0JUMhIFg/DRLhcAoCUW/RAJJFv
qWkm9fK36ReaK+EPzVXmVmYRTjxwKlTl3QAnk6UaXOZTtRgBubareeE7f9OdzTqn
yepbWPABxHhu5wo0NZiIMt6l0j0Kke48kEU0n94zkwx8FN9PEQgEaBbc0q+J4XMh
Xe7n/fL3WQHbgzwqA1NQ7qWIe2E5+Hte7UBw1Tmn5RoEY51/g6mjxDVSWb++8G9I
k0Bb8SvL56QDe1OP3AFp/fSKyQrhrYRckhroxYpiaC7z7YTtrjzy14I1uVFL3YGf
y42yYHYET1bZMjTccFCML54tK2VXgT3ksQxJqs1tVLheW3dk0BzW0RATbASHf9aP
ymWv+M8CPcMe4xOYaxrX3Nt73Uknpsz8Hpd5I1h/nCZoe2eXxfAGFciAf3ISV4Qz
kSlz/Z8o/XD8pT66ZIJ6ZmuK4PHbl2De6hyOOhS9wWVfzHxgZ/3LKdStTKNfvXkG
idqusCoqSvAhDgvCJv+yEkuALVlx1/o/hbV7EXMRHg8QLSHzugEplzFddwS8K+Jv
BP9WfG/L2uiyvZC96IZLXn0xkTZiWBCBQyPY/60onhpDm5mY9KdL8PIvVDRktbLS
9MK/9vN1tRKKfXsHSrETWEWgf8antmeYam6CGPldvAwRQYcR5Ppo7SjouEuwS040
lBn35rhIF3gn4Zgzec34B+9PiBKfGIFKsxlWXv3pJEp+9fFVjkOqmnRtmizTOBKr
HOzFcVyOblErPDB0SQKOJhnE8wPLXS6EdkObw9mmo3QMh/7BlAyDSlWPH/ySnPfP
o/rQKv8gM060ZZ+aHHyAdM6Jb7a2MuZWwS9kSzB+0PSOirNlm0LEwMkcy6y62SDP
RV4ICgy8X8fungeZDgZY+6+wQwyGFuppV/1l0IcF7nptiG/ugAhtFsoyE95DGGsE
R59/UXb/q7lZZCK8Se+DK+v6kWPO5uCXmBRDV6m7Oanew0b7iiyiTeEfJZKLV2Z0
/J1DOmlNuaqnMGNv9OD5aWdTzWipdAIJBjWqB/Ecjm0XOgqzS2d3rHbtJUq0p0ql
7c4bCIPM2s1lShC4K8aAGcoezi0TCshJ5aVfsc9EZMhXulHfLO+KlXitJOfmgtgz
NLDGlFSTV3ptXQFqRaF0DhOQLj0A8ZBaMqFT1U+G0a7vl9pfmxl/I7gZtT8E+Zc4
Clc1qUAPuJjF0cxeyxCef3I5vEs5BHGYa4XBy5qgMzEYcHXk+NAicq53PYbnLbc2
plC79HiT/84nwn27axW8HtEuYP2RQNbtojhOKA8XcGKksW+GglBfgzMIeU3lRWgM
6TWj6zlEBMCjHhROth94QllQjiiX0kxjA+SAFwoO/598PoxKMXJ6qvyoMPyewHnc
dP7R+LUE4yg4XSHJHLie+KOOxf+K9ylW1PDPQsWCi810BulsAlFHnSTugkWwVcus
QkriheTY1iHd3k6XSGp3d4YiCV3SlQucxw6CWO4/eiTlLZAtM0PFUZUPWYW8wZqF
GpZj1CVanFIc5Vii+tlatM9MC6GkYXP/OFxR6UEU3qlxt4ruOLC/AQa6iIEjU7pB
nksugIq9XfD6SuKxxXNOcskrUfr72W+owN7LhW3X30YV4wFvzdiSe2jdlGfUwIQ6
+QO9lA1Az+J7vzOASiTwDO12bRPV0UV4yOshHZw+qOMRB6/g0+oJpGVsB9Q8+9Id
ZyBbK8BRq8vKn+n2v7gk8KvYRmu8f4fsIA4yhgd1cphxMorqNz6TmXuRHaDNmhCQ
ajNXfFHX6L85cwrAHwbiOhvIH8DAbSFqwpYlx7RJ2r3hCQSzm3KyNHYKUP/Epp/J
/6shL1CPR//6H7NC6csAikBOXgaGcMvD+Me2I77a7U+or3tVl5RU3d1Qy6HFIKuY
C2BCedELUSMm7/QQuR+lP7w0IkkKKNSbN6JffJfx1VIo/Hn8GK9Ig6NCza74bTuN
lEWcCUN+V8w8w52evJlMaofSXZLtyLAJ7D7gOiy0EPKP2Ynx9a8rWTfDORtSxlaG
HDjhDT6y9k/W5FkJBMfvZRIf41feidKVfridYrC7FAzNKSNAXzOGH5GvQIaY6UaC
SFhlRxFhXsCHKrH/fox6Q4Deq21h6VAeBz0Tt/Ib8leQWKeLkCnpiMwl4PLW1wxe
+kEY0vHnIc5OXshXJF/LOH6RIkg4PYnNfB++s2xxZXzMYYu5vorbMUk1iUTrQgTw
qHDhKShrQlRxaDwRAZPaHgzm7VwJLaBUe9B7r/EVMxhfc29tIhagaQ6IkM3Rp6aN
FWR2CV6lYMQDYOYUvtyD8sEj0k5fAUtdk2tuVnzftdCEnAHKtXT6ek9uu2BI7jJ9
yCAf0xfbP95eegiV6Pe3k17IKs/DZed31RMK/YiB1eKoJsln1vc57g7T/O+e1yLc
gZUUkV0fcBik2SbI1PKtyxEUPunwgfBpEF+KYdw2EqdYMNK0NrQ8iPkQw2hNhyx1
x+A1hQulGaWIXgAxI6hAp2WjzP71WOjpQaNIR0mVijEQWRWe53tVJs06IPXSwH2W
O8IJxs+ul2KSugHl4u4XykMAdZ05WvfRrK+g2aszYlKVVpma9FzsmklQy5Vw57qI
avwrR1TonwFjNemf2CxwAPqRVRwM1sTusgZdtcXL7d4YZwDsslRXvgS6U5jqSuA5
0QErWL3GFJHITKBKokxlXxEIlBl6RVFgishySmqFlwSQfnOHF69WoXj5W6Rb2e2q
bCglc8nc9U3lJ6FsTl3bVvkhbHh1xZIwGPTGsom0cPT4ASPBgQdIm/odcUsthBD4
gCEQA/x15XoGo28ZwOaBD+a2Rt5UO5VsPww2+Xzaag/bmr8X0L8OhSw4tkrzByEe
ZyG6Y8WU8X4GcNn4IErvqnEKTR5weevBF7mRGJW65tKxQMliW0xEdHcicxIBarfa
90e8JCrskeEkFJkhIFIj/K+pA8VDFZFX3j10WGETUg551AHX1XJXOP0lyq1LpLZf
V4TspdbxKa6V80gOll7681Lhq2XqrJeQWeqA/i+0VXt0xUCjr4cMqb9bEfm2p3C5
1Ze+IzRGDGZEenB1SJTVQRN1HsmJsy17xRP9BW0HrBQWWbjhSjAV3hMta+m2fxAI
a1pxPcNIb11HzELToEmOG4uQryKeBF82G1r02H8qVF7D1rDpx3VbyE26qLcy+b+q
8Vr3IEE0NK54E547kNBZwFmwzzdD1trbV0qsSc6E5RXCLerBKDgJWYBBKNSadG5E
PCf6SpLCP7ZMZRPZbjToH+S+kTPIWDqR9+GksC5B83nsFeadPfcohRg0OpAMpcf0
w3+czW7Or7XeQv51aVVTc+3GUQXnn49ePjmxMve5yq/jXklRz/LdVv5MrAPAY+KV
hRwk8rYHjgDFTsZSClKohTCAzAXLCOFkbdJgf0ch2qJJ9qMO4NLwyO+I4CHUi807
4D/xwNTIHgANXEsRvOK7OUhngXtVh5O0Uk6Ky9gaiV2U5j13pVVCMG3EJGg0vpD2
283weWZYDUGFIDSwStbbe8mQ3MrL8rYip7v1GdSOEkGEFIEkpyzhHOFCEYEFy3+t
OkKMOgt8KpVW+kcgZlXzYEUsZyv+2jcN6l9v5x7DVfKosjsPc4lN1IpjmOGOxXEt
tCt3kL/Whmze2daR2S+d1udGk1rj6c0i9SEUWpQFAaHeNlJWSZnpNYhFT5PnfRSX
0nHdP914X+yBf3rNRHoedK5rnW6oW44MQuTpKKv6NobeTmOuGsiu0KtI2VzaT4wl
wbM6Q8GO9BVvvXKqCygiRa9YQpiAYwE23gwtUy67lViDSHnsyu3/LnG3IQFyd3Qd
7KQtC26GhO6MutUWH9AFSS2LebGdPu1kfLmCVErPziIVZzIR1alQsRXAcO2fTtWE
WXZWBslEc5NfVtdVnRwP60FC0xHz5LlEOsdyN5Gy2fR66oSCLqXpXSwbsYF5AgaU
sYK1z6WBa7Jr9ihM49QLSi/r8GOH9gsKdwit8lNZVX1bbdGUZuZMWdVo5jAqkD76
bLap20vvsDhVKWxy8kuuyxEKRmKlEWlbjd612akvdyoPl69oaeMVux78BV8uyabW
bOwGcRW3jzkh099NLZXap5C94iuSVn4sBCd+SGn2WTO7eS9YpeLT3/uNZcOPWPso
cLMSnX/l09ShzpLEMm+nED3xwbNPjEPMZj1jFpwRornBE/LiCEGWipeq0IJIyyOZ
fLX66lnjL+UjJsjNTWlIdYlXjN7Dl2+RfNV1MVkN1jC791GlCQMCrj7QSUtkcM0c
f+FHf/R3U5qEgmkOvuPIYqhQ4pv/bqxq0zYonyqmexyvVtzATm4OXYganzncsdqt
eJAv87+ZnTe3TN32FptVCMWxCWqFRyRo4t4WSFBfFYBR5dmNSQOwtQa0SJrr/7MW
kcM2WeudOYBwmMUHWtiADfiTUWSf9IZ9hgCMCOK6tXl2i1lCfXYObLvpGjXRBscD
ghq0QXIjt/KKQsbGQdQ8DAUE85IhPOM3WteFZFM2Mlyjpz524/9E1D8iuHIeztDk
3Id82MngynjM+QMKgeH0On5KLK0VhfOBbgw1iqJp1NXGKoeecHqUrUAVAqt6ycvB
UP1owlXVD6Y/tSpA+bv7Ofdi1OQIFqLOZZAzr2Y8BTt+zPQLKc5c5w+O4iRj+rLT
jCynAw9JMumxQNB+bWsA7ADPekcgbEWBPq7yIi2POvzkHhneo5NBx0X4yoUoFrLM
sgpQpPvxUr2dqxSY4jRr/Skrd18echgXfkcME6OLTLuzy7Aq9ehkr+Bit5moxeK8
vkcxW7saBIt7sU56uFL6urIdNJrTj/VfK3PjxWZokX+I2H/a0ZQ9JvsOGMW1uYeK
VB2hreoZzlcQzgo4jJwBJeaJv0hqzJPUxbvnmV0fayHBgK/prc2KWN2kMtcp7LHH
anaXtAU9QoF2Hq6jTt5QCe7saqqnFzvZtawfiEp8EkIEHSXR4OxKNXLYsSath90S
RyL1aWR11+QwpmFYKY+x0SAD4bAikAKYVSDbOULwkQUH+Yi27eKlHEPL7ze7KAWc
G8LYBNU1HfGaOthxx5BRMOLOELLdnjP4hsctUZ+Rrx8OfRg30YHZJc2GaCEugFsR
S8oCUfjfOV4RQAZXu+1xcPVq9tx1AwlNMhD1a9Y6SgshVBZ6gIqp1RN9J4BEcPZ1
6HThx7gyGR/MYV9D5amwwBU+IK6kF52+a98hVDYlHQSATWN0OdPRpDGarjQcnLDw
T4FqtmhT60ihQiYFVpC3TEBEDkYrE/qPq7sl1DrdlA4kkUo1sCcImlR4kZdzZ4Me
sjSq6ZLN0/3R82WrOIFNtm4jYns4Jk2850h+9MeecfSGPYdrKVnnTk7qjB6gjLad
ZpbMIGiTM6IaXDaupS9M7brl9x07jhJR0rw25O0HAHO8enquU0SM1SzT1H4G6GFw
0AgFGsol00jI3ypCegVDZYI2ual7Ylkk8YyB6SIczGQoPg9riV/Im6GP12F3tBnP
qawKEV4X2otD3XEfB1WCclxDnUPdCfDZ317Pq35MCYUBt6lPw1+2QGrBHMfUz7EP
ovmxOQekqXdF9TDQ0EcQn5VXc24TOlmgUwm4pAuG7KbNasEHHkhjCR44K2vMGvZv
HFHbRCZ+jwXyrOuVMFp6UjIi2CJ120IICay8qFlle6Dwm8zfKNvRFrFDkXdR1gz9
6ZvMyHgJRv5vIa5zPRLBsQS58cLInFS5h1MsK0ouJ57f14DzMw2nJ9UToN+aITjo
AM0q6NWNirMespDLR/3eKP7RBAMyi7xp5aOsazOv4L5TfgvoYm/u9J5EIAdYB+Sc
Ew2BaA1kOYd/+z/ncLDb2EPjqtyFCCdbtQm/ZwCMTj0U+AztRJnIfd4KlXduHrUE
LkZxZKyjMyT05bRDLLqxgMcO9bnu95Yq+Vr3TpNgL1nF8s2NK1oF2+2LIiJi81bf
LRxo2vX2Y2ReOXPLdo4NJQoSvmp4prJchev+26x0IXdcjWvOZ8aN8vFmxiKVrVh0
He8197YKQm6YsoDIfcg0XY7crzvjnX8FK93qXEtC52cOb9nceWB0bnwUQvx3eJOK
alEGhrY/zhUWAyGr0JfKfxkMUMOx6vwVHU2VQ6C2zcaGRqi+IjHfk6BYgCFeU2dL
6kWukkXtHvzoTsx7/g1KnnPYAmOYx2IrNFKmeWpicEGagZ8q2kD0YvJM1k8b6C32
mAV3kVFCCEXuAGYImrUwny1nDJiIuqUrciD/k2E6bwS+vNDgK7JuZsanUzojXPs1
vzNC43y5WwM9O5w+C/Xbenjcreof2HyabVpG0xc7JlpRatoaMWDYQJ2r+4L8y+P3
B3IlmjQs6gWiWGdiVAtnaqK8C3OeGN0EzIxjAiPp326RQWv6wP9P8Tu001VmNtK4
vKqskLraQh/GqvqsuZn20D9GIvBwjYcoIUHugO2nhPNBUUZ8/aWjZB9u/taPlK65
qhY1EFtOjdZXTjzMXUOHjk7ExEQjKVugdUAJsP25ohQzOS1T962G3tCi9zcNOqO7
rqd3BW/XqaI3MRiLHrF6lxEQqSZEFCRwE6jzzp5fkF0yYK1hzWZdXpDkYAHV11zm
KMBLZPAZioSsBp6prad4PgNpUsOTpHAK+haZio03ioy6+iQYbDOMXitMmjoXWAjF
4tmAny0v65UG28SXPQ2ND4khSCjPbF5oePlAgNV9kPMA1yKQ7DvyFODU/udxjEi+
mVD7fPdz3rXB5YoGUDWV8zHFTtN6RMua2XLppycgzN0N6hYYz4R9xXsy5y8NtJad
T3H45hxwuC/v2goF7KKsffFdcYBy4TvDcwrVkGzUOuLhMqyMGlGMDvC+Uybx4x7t
/yXCwv5eUOGh2tkP/y58Fuf07C1NXuoiVHqKzCjB2nVaLF/Pp46+QJKinW1q/tOf
91p1Mam6enB6hqZcwx/fMy+5VSQv8OxPjayEjbrYLLN9gQRQ1nZzXxJd/ZSuzdo7
SENO5oe3q3lcoD64Oa/cUM4gkim3fsfn4ZWxyYLMcAAcoVebcaP2Z7qJPnhWibzN
nKb50vZeP14i6AxLBUjEOlwNAKrD+0EEfksFnRfppHsHgf4yls+FFk0SdBB9dhVt
7snr+J2ZnwG2yE4LfneAf/5JD5HHDjqiEAoFIJyg3Ap8ONVhHD9tUBuoKa3rqbXj
wzeqBvwp7x9rXzYSRu0Fh8rfZojOJbALJ0/TCsT8mUS3tXcpWTzYlYxmu/UonC9F
kOcFeACNQx+/09L62IP9TajhuBcFL8+syL9ro+CwZhhlgh7OnI/UG2upAPNZDcdV
UArTuSLWCrr2U+nQ6KP4HrRo1dacFPLKbcgF+0B+ZhJIs1QBuRzMctlUBjRZxdvZ
GM0223pTJsJKVJd8/7X9zfCMmYXwEaRtXwGcPBawjGIeHCKFOPgiYBD1BQy/vW2I
kqSw5PBhGnYYu21t3fSvN+qmUbABF5OO+iLy4WTV/NTv2bJeKlOJ6zbeaMkUoJKf
pCVIF8PXosZVPWiuFmkkOjFOVzXIFiV9WfbKiSajQhqWFNBN0s4Xta8ucYTSZ63n
FHRdXLMrNlT+TnEXlCmrgLcKG0yeCB6BM//LCYd2TvBhHeyvSS3gCuRbKJgAH8b/
2bHGObjRxbsEBFAcYBdW8X4WGyDJy3VNSQR7aWa6X73CXzIJt+s3jOTOL1nqMh2h
0GWQH2ALMNb3HPSJ8SH1pqSy2h94Ldh4J9o92cP0nuVXPdhyQ+YvOVUALGz352Hi
Gc+oz3suO3I7tYXqUi8X6oZfSZNCosnaqfq4GaAKqmSFwO5t4Q0VxMGOXUxzJRm0
1y5d1Mp6KDR03cdoKHIui/XeGq6RAOo8K8WSO1yjRru3SAupTUK8krd9gKf5bV/1
HhKahgPOpoURHvjVV5pJMaurrQewhP3A22AqI0DyuUl7sL34Y5xIjiFkOObDJDsS
UbIPhI7/lKoAix1bALzXiQB4apaNmXw4y0tfA1yyLw4Fbek3PJgMvbk2ayCLt6yC
XSVA0Wyok3hTeYL+0RmFnRP4WdBR2Y+Kdql6iP/iFRBulZzBemX9tntk5oWsxaXr
Np12g31IenCW1vYrvAQFJ2IK4C/uIh227Lbv19PaQyTzeNfmVFjiFBTXfylv7N6A
cUSLQ6LODIDA2ZIh63bO/V/Q3jzasYJ5KPo1husbHfRPgavifoV9dt50yEiryfde
rS8et4TwbpTE7mi+E5XzO74QiCrCtnW55NBv7fSr0koV0Cb+wNtMJ4QoKTvhwMeM
NL0Nm2LKMiNnP5KCDjHIiJMGAx+dNnguYqDmtxGydfKObcS7FYcqmPvZlFfbNkLy
XhLQyJfkkvMIs2isC2jcI3vajVQhFKVbr0ibYp/YukR+6MkiQ7CA8MwOE/rDghym
xerDDF7XSNGz62h3eOq14p252EryHNuqRI7ou7yc0sLA2WtAMH+m1xnYXj3lDSP1
wOUSs3X+Yd1Sru7dykXD/E0cRbjgNa6mmtN5rt204mk2KClZC9/HvTBkHUArf8JF
AnvhNiQPx8/57w+qCGOQi5qQf0Y4NpNLcilLw5s96MyJpe3E2qZih/TZekiRfpFS
+GwNtdAOnHbcWlx2T+zwhEtXAfgW/ZcW7O5xNvOUdMZjxjZynN+QUA2aNU5mtsew
yuJ/B52LkAA8Fm9AMUkTuynYBjzRTlYLa9icVWIWvyq/FF6tkzx6gm6qGLwJRweF
K0QwZwCFkIBK4aVK1rsf8d/rmI6ldv7xKjV3pfGExila3V6Xp+DbxcZvC8z8sP8u
albEvg00aeEQtZB0y67g5y7YR68njKWK/jc7K9vfJABBXWr6b+zM+SoyCVD4hDKi
k4GZ7wD5bO3nsp7eDEVAE+XsHBK8gfzmdU0/pIU2x3ZnfIvgs2+rV0hvg76hngyu
Vl2czeN/aLmdgfZo4v3oVgvHnqa8OljERlKrel90o23PscfttJK0kh9dwaqiaT8N
QOC/7zoMBlrGlO5kVaeSZRyq82lzjtlWDJp3ODo//PaIrRfGKwnLgK/vBNqnCrg7
90rJevvjb/qNdhO1NmXcEQ1uLnxftVKM+uGbvHuz9yKJ/9NJ1xpPKfoZ3VXwAQ7M
KRTvHauQYAT9EXhmcrG/W2VUJda7ZqtCRWR9iy3+aIG5iUEdwKAxG6zIejMSua9e
c5pBbVQd5uVw/g12V3yNd+5kVbwHt46X56+kvzYJQyQ1DwazAhMjodfv3UkTONZc
j3EXESiJJ0YGohVFT7smhz2zMYYIgdBVqZkjx+ri/DV4L9NyZDFPOsaLMoVbxTJf
QlDnIG393g5ZKWTp671r8z/+bfyXESqRSyzJeM/3Ym5xK76nLE0ot7C7OoVfjTIX
ihhApKNNMQIOMM/UdNWZU5C5P3bUQp/RhBBV+dzDxS0yU8LTCxI7iLhHdF8fpLhg
c6pfiwJKcdvyBNUAH9rYcWxIOwH7cI0Ote5ug2I3Vd6Kwty5PNIMHLzzvljtq4ig
3qtQKQBKYcpd+J2HzoTClwibKFJlxh0/u4Dpe94/KqwRqGGdH048YXC7wUNS6DUV
/ZGY+XvPxd//o/eD2l8LGIbu6JPofXhoAQJ7tvu+tj99D2sRyKx2h1bDphS7al2r
/7xcLMjDEqqKsKUWH/v3ocecnLtNec+Sgmsh8XQ0Vo7AAGbhbt0jGBb/et2RCDzj
O23w9srwJJ75GUzaXIqGyOM6rNS1aNaesxhlC3/V0Ta2d8x8OgwMAaYO91I6K5jq
lo+pWbeJJbNBlZGPf/MLogZjs2+UmPIU3bBelWE7WM/J3O/VgsmDhOQfaA8zPms3
+lSeBAF1Yxst/IqrdSZySh3rkm89qrOdIn6ZenTN9QC4RSNZEZnNbPSoryqpZDnx
c19tF4blDnJxgCPixoBEipHcrxHFad2oeKRxv08T0d1bUQMF0Za2cSaW3XdCbain
csUtCbcbBnU6f3H+QoUs3/9qrjFQ1WurnhltqMimmQNw34s1NksrrU5RiVwybVeQ
Yvk0dPvrGiFpCYwB5gihPHcywOvJhSgcZb/jKYJ9GE1dVxMF4ebQEr2SP5Nm8EqL
wlYyJQ8CbPx/71zfOiUajNaArKOtgAVLWblkBmxon82uiO4hAGz7JHGt0Lh71VtW
4zv8hQwMCuR5kgPZTMz/5LSl9hTt8f/6u+QQm6ufLbSgnJy/6vYgdTToXCnJIVVN
cHz5msJ+cVRiSKFy+JpbYIXi4M76BTu3la7eGsaaqrc6DVWhxptd8C94VGCEmybK
3gjwJWTkj2jKZMoM+CLV0tdWPN7/pQc4ashsNiP7booCzxpY423LmZMCIEKSijLC
27JEFbcLlzI6HLBInC1V5w1ZGjZS1bIlgLPo087MkPXDa6Opo7qIbi8fdEB1DnnV
6U0Ucwm1Z6MwVWqwO40HCFEsJjaTxVmqD/acmD2VJvDedeqjds56jcj28jVSMRXn
iuGqIDCvxcSieuQBI+gmSTNvMsSUQ22inqW5CWKGQhziUmeZWZLoWAXwMFKbSLkJ
fMToJRly6IBnUx+njBTlxAVZJUEEfKzvpAUZ8I9zaOeLMK2DKEhtf1nltauBVYmg
ZZ29j1fBK1bFrVVaIKRpEfr/oeUDfkC36bRWl81+w/h1Lp87fzOv82NSpcmiE8GC
u5v54TQ+MR0axTRjdgzmejXTVucjoyaMvdHwpGzIPNdDcwSBL1Y9P3Hv7wuWcxek
+7PFQBnIAK3DnXNzYP1v4aYSrPMELD5ezKb5rTeShJ751FduYwFG2S1NT6Ys3Emr
Ym7wXqqz+Q32FQ9ZzZOSPuEEv5+l+fumTzwKfuUC6r43LPRHTG340+MSWisJJYP/
V9KYhp6q6SS/5BVvyiOnLy2tjycdNRkSTiW+BMsGkAkahF0M6Eaic/DTw/+I1FHT
nSeQCBeUn1qcB8xbqT41qYf6g9A90l72tgRhbmAhiXrAaTxYkSHK8JquZG3+9vTb
/GDjZNYaqATxjl+WOmOSWYISu36Rxv1NjmhOflzw6TMaJp2oXu8LulmArgXVBVcf
qK5PdyJ9yl8vzoT5v/NuEOjmItLtTZ8FUAwnq9bAdjPcbhZLmUej+G874A35ciYN
dP0MTkNuxkjIhYn02pDiPA+orwch8FheJoCN9pUJVYZeIq9CwsXvWnTljmGHeIoT
0BFhvDIJAve5NS8oAus3C7RI0IgrprX/R4cqs3kJ0ujX7o1qGbEhaF9Aoq0UGGCG
Bo1o2Rf5bT6R4xeYc1MsKR34HY+2elFRFgcCV7Knx9WOqXlkza38IVv7Tkp+QWzm
ry0nakf8xOFFZzmsFZIFZGaV9U3zbc2xwpAvwLmziqbTrdyPgRa+JhfxqxTJbTF1
xMHF5UMOp0Iu1/L/Hza8WpOq7YpL3jNlCffAGMqt80bqwqd/6iY/Et06RsUgKkWe
YCg33Q1vHZgIfRwI2NeN77a1lgDloxyENA1o0lkg56Zvr3j6WTBI8XaY518ZEoXi
VKJMVgiwY0aJGLtzd/PUAluUotBkd6U8vE/F71Lb/vE2Fd8Ns5jUXcd5W/dJ/Z6L
+0V3SUcnQRV/F+hG7kdSAN6dqJKYRAwxUbfpdmIC3OfQBcPhagZYtijkoJVg2qye
G477CpBrDxSpSMwRFZqq82/lgwDDrRL6TPn/Wde/daFDEPG7lH9fuG8y292stqTT
ThZgBhJLKpSdil+R28QSEyA63/TzWv+lLTvY4iPd+aJYEUUpVL8wmxWGThPIcODH
eMH/5Vb2OBQb+yPl0t2uwJxx0KEAqF7XR4B9Sq17i3ESDXdiZGMMIndl7fVecHfa
KOyAgWOnYMLk6x8icgaQuqxyuEfh2q3U8qO3mTkz68rQdUpU8Bw8nfacCqjsXBYN
WjiCdoLpN7rE0n4/KzpUwrxTSMdoTXlG2Ha/x2O7bVXz5OJIIgTVruUqcyjEdVAy
gL9z+ZllDKrfLlsQz7GA/2Vn2s5gkc2SBrwP8kqFG12Sj3rdfoLFXj678s4bIHNU
ik4RNSu9o3cqKDmoz2dmCAUYUczLgmCX85JW8/99WuC57wb7+DAH6KrezVDQG5Av
GmWbp+vOFRwWFseBqD92TpaJ+gwlfqMgypd0y2xQTFZJlZeGebUb98IimCG94Ou3
ObkfL7quGuy1dWHNo7IODHQz0WczOp1CijpmvS9RIbAd98T3IDaot+FAYkZMv41E
+9dZoQiigETw9kIa4E/wGL+mHKwZc8dCcAJNf9pTccwMrSeArILC73Ci+rMYAGdM
0/JR1cKJQGbxyCaXvoEa0qagj8AIZfaCzq+GG/PP0hPpjHdKf0gw2IFgFEtHB9p/
QtBO39bTHE/2a1orxkqE8cgPQoNLmxE0f6EY80HaAARtJb8QUXPOjBeBogvRShVU
8dxUDg6zRLF4EPwj3/9gFUOBLB+zto+gxH9kfQTO0S5Hdti+kUe1OranHccXTJNF
teeFLrQL0yGgFzwpSbH3hW1tUDOE9yJOtDHGbr4+K0aIlqPODHg7Ts89/GFRZupw
HWgKG1F1mcfdkgTu1D/aP1/FY0oJKfPOMc7WiDH1fQqaw8nPVma3HH6D+a8O9mYG
14ZDTVUTKHkFWJ+Tf1hOTU0XUYrHe6Rr9FfwM7ZDuJFxv/BBni3gyoW1gV63fMFm
587AH0kvz1NEHFkzXlJCiE6Lm8x3rk/ZqQ80cFBSnHY5E5T08JOfY9lnAueZ26Gf
2LyMW76GLZFDkiGMR8gV8mtQ1q9bhx7CaUlx5pBL68bU/bTwMyaeeaoI1aOl4JFk
26aOVWVFpJvCXPXamaVv1uhG/klI2Bf8xWablu2RT+UCUzfMx8MgbvomIK4cTJXI
p08I8kBwjY5QPI4/aodgGFcnfjkGn3R793dZPteyTT6FseIdhUNDiNj4dGbYEbi3
iEew4ugUTe/YpSRj3V+VZh3S6FvznTV0grxZPfpHK7APZ7g+WpYsRYghDp+M9DBu
0aIJGA5JusLJUpREQcaMnIRluYFbxMjAv5WA6WFOIvpakmxMzIMJouXJ1iq8mU34
AMrnKui2Jj4RKxFiSf+0zg2/B4NAuZPZ4GgFn8DRbeARCuwwqhrQRIwQ752Ure4+
CkLyrMw2U9RHF2F+YhTfOiebFW2uS2kR12UDmlPJ1vmAqjerv1gL9TuufJZo/0LB
mJ5zJRzPMorUJzrGWDR684cVtEy7HI+exlEyG2ZceT6IXopneimpShfMaJzi9wJ7
7dv7xFruBHVow6AMyxgSmb6Gx+HhBjuKyXmsvtZXJyjpcc1EJRMqlQAMkVpnR2WI
OLhI98dHqo9D/NlnVpC+By+sIsSM9dT6tJvUcXS7embFt/Rscr6bg/UfJ1bbyTO7
RqMSv8/3QlZW0Ur1zsdNQXRgn7LLbH7QnlrmtoRPPbZMbO9jBOYa/hWGrYwaEDDn
EJorxdZdIDzPBtDotBf1AvktLVyM9pj+4PXu43cKE7hXOUi9CQXRo1slwGqVfjrc
TgBCuAkyUX6sK5My1KthE7KuS9cSPqG/65y/j+i8NaPAQ2a+JCoQvzym1Og/jVtq
PKYvGAZRdbamVCsBePg0FgRJdROs7mnCChW9XxXIV4Y31qaYubPaFrK9SYpTbbF7
rAQ/Bxei9KM66tUMvYEEZzc6XlYeQ6EA20CYab+LpWkkbsT0k2QUArHyNjswIuqx
iCgsb8RZZQvIkki5Q3aXkPQad42UNRLfiObNMjSJ/Qj7xc3WjGi55NHMqy0UGl7L
jvnPPqc18E0MSy+5JuMRnKY2rUTMDWjoRBKRKrwpwbFwMBub5oaFkfxllMeAKnFB
Bb0JjLLSgmvBvgTg+2q8EZQNPEiNxFnk+9rdKmzosIrhfCftiEzb9JenHiu+DN4m
nekXriHMNV5E5Ms6PdbQJ2V05JCBJTrXhmu2FANl/pnQUrraydhxWz/GdQJJyVvx
V5NbgipdGQWgywGWw7x5tje0Gu8H70I/SLvpQdWVFiGCmCxAYTPdBOEGJ+5605HT
Zbr3JK2AjfN5U3olK4f6v9YDG19n+vC/VxQZrAhH6dDYPfPv/YayMgEbVt0Av8ww
B52hUviQ0J/fcrrjbmboax83mDnDJhItpZzBzSthV3scJOAp0Npl0WmT/dSF2FLm
iqjKDA+ugWdg/oYvBAOKT3utTTmepkKGaW0clnn0+WNNE4oouk8/Ag6y3XddjrKk
0kZQbUZXoow1+FTMbaUABKgC4DVGoDJP1tSHGePgkjEUzCq2c8Jd1N80NEwpa/UD
Ue07Yn+UttDg5D5konq3sYKOqkoZvOGISxxU8Xrx1M7od1FPOtnBJzPBP+Rympf9
lSB8C71sv+uZEIsTkih9VXOVcytd3jNuLTtKm5pAhjcs5330pPIDEBQiH8Xk1e2S
g1g84Hzcmo8MXkZ86WGEikD4TW9LS0EeJRXtAHtcGUcchw5g2//Iy3aI5BP13aRX
NJogOaaieP+jtw9vIf44bWmbaUAAJ2+J4/YknKKrB0HQEP879SLN3rx9KUNaVV4k
AhdqDhIL0NPxXH5kpVb9ANPbgqfTWT8faVmCwOOsZ4NBBFwBFshtLPQKLhD6KeWc
zNa2B1P4S9FEDuHjOEVSxiqm4LKH8gSzwuO4Q9x1dRU5nxwOXwxonZ81l//Lo4u3
MeN9EaUHld9KEYbX5TVbqcisaPhYFAm3IQavsuhjwRhDYPI+Gjy9ofef9oM/G/bb
MrHfPeJFMjtJrp5PdqVtlHVBWRMhmpZMZb6OXA38NEg8kCEDqwnoEArRVeEtbkDb
j7309vHOtemOc1V5Gjl9hFc+ZGVzV5WC4g/mXsd4ROxLStfpMLm5y4hNOzMi+NU/
aqARm13Ll+JiJrNEN5A/auH7ofNuxy47y3v8jWlKDXd4QhGk/UgnUo+K2eNhHGpK
xRgFIfWKn8pGMbTbz/7UZ3dJP1ewUXtj4v7Pyiaqy0Rj9rpzP0U0Dw1rvaAEltbK
j6dXjjeqxIzAqveevA8QUMgtnoexFSG/PQbVDMNGS33t32Nql8XhA2Fk6gDIM99h
KzXuQQy3wgJC1DGj8h1n9NnSBgSytvn/kjmBh1aYrPJdPBxIGb9bR2RYdgmOGrKy
/dXGa7IguDmC7llWRm+Iqr13nk5qJfM2IViBPaF0e1ct5lEiB3UxoPMe6oLXptc0
1d/katxVgF9NGODo8HbpnMvfmUbXP2X6Yca67hb2nT6uxv/9FUxj97lCfcxKh8Er
uuUQB1LDl6+ET5Ea67IEJp8XK4sZ19nUZw38gTem/uKoSSRTEF/L8buJIKyOOP75
Y9ELB1/7ltzzO6dPkO6NLObQVl7OWQkos1Hl2wE9kOm2zJIDS2FLxtw82OcReR/n
N5QY7hp2N1Y60meXlqP5nNz2lYiE0Aki8XydORNTcuXBE1lc3cW8Z0zrH33NjqbT
uM7Gr5YVo78sk1SdzQ4croVAaOhT+gnQKnL/YgQNmakY2ly7rm/PMZ2vn6vwObf6
l0ErmxRTqMbwyKFxT9Fwm4mfUQL1Peg0abegpp3xtybpXShuikuHTkmeMVTOKUwI
KWvLyu4vNd6Qo+l46Vug9EhCyy7VeXzwBGswrzlTl13EcYqfw8z74Zv5EOmKMTi1
xXb4DxC6Nh3cieweurDLLRrbMY4wPfdeuM5CqXb5ulQckGs4e47gT5P+ov+tizFe
R9Hr9rcnpJ2Y1mg1t1eFJcd4xtl2GqUCIuzFYpOKwQGhKwoFdnsn2m5ruAu4HtDp
3sDh+CPV18vfoVGHdETQ4XVdaaqYWVr1LoOW8VtM8iEb7a5vP8NoJpO6BH+haiR8
HCKsipwNKXgjg6C0ipsnwgG5sCWPrNE/DZQPve1+Daw1Blj5SqQR9nbpSo7qboc8
VwQrvl5QqyIJP40P8CVZgobt9lg75CVMBP0nVKaP23JZjgkaUB8+No9QcQsKvx6n
TOsnCPphrV+4JIP0WiGWHHa81+D+Svfj96UpNCqYW1C+o4MMgAichswZuEL12368
Np+9iFwyMTWwh+Tuc8BxvrkTNIZbTR0nncdbK44rBZRgS0PKTo8ibD8pj2XT4uQW
82DZENoWleojTIICPg3aI5Dxk0KP2b9DX+pwlxnzpKFrspON9taFZgOrM1myl+hW
zc+VQj1j26HE9rErqYU8BSR9tocaFe9DzJwat6g8lheNU2uQWHnMtDsFDD7JPXSV
tMuwAKzyU3IgQqZdTEsPasre4b+pinHxapCiec/ygn0G3+/wiyUshh9b2QNB3i8r
WOg8zYYeb89JG2YzC13aW3KPTHdEYtPHlwj86Zz8Q/YVz7nqVIM6k2aevIKaOTq1
dnJZ8M2eBlnv/nL+zTxhQrIPjedUu/aJab9V4gudFL+6Q6A570kCbPNmCZ+sy3eK
Fy2ll0pH/F/VT7LtAZlCZ3rnm6Si/nWERkgo712z32nFYxmaUgOWPmxG2EK+nT5B
mQUzKKsJCn19eug/mcnsLlmuXikVbS7ZNHmVsUefNOU00GQ0FKYrhh6uHdSZeq+H
/6okNwxbZYA34qwE4Ep6K/lz8xdYjpRuEqFp7OL3Y3XPxKVDs/rqUlVVwzaBXoqL
HMWmYOQz67c+J5/oCdoE0jNlmD2zLW8Yjbc9Ch1dwAZ4ALwgVAVBvhN5S0yL9DYV
OBaz47QWvCi5eVjZzFi8VE0CzcDkk6OhZeSbVHZTFsTSn9vvh+8GyJhraWwe+HtR
FEm4YaHbz6mGxAr5OQoaW5Xd6tB0185nTCEThf9KvLX73Rlb9L7qA7bABcoHYMxg
/RGk3M7lv4PyMfokw8T6SgZ9oacrrY74dab5pj9HlYvb4B0PmpTr9DCPm8+GXjs5
LulKy9J2woBIYFomqpxJ4spb9+NOmwDCrfGQuTWtvmPCHFcg8s+twc/4OyWyOJoR
Tj67EQV3+XXfmHDQ2CVcukItelid1dtDYTClw7T/Oss1P48Z3HVBNCIIJdRojrf0
gFiNnhK1U6ZDSl8mFKw+tzn8B0kQC7fZZX/859XRA70ChmlwzVUYSj9AzaE4WFoQ
Time7EQkcFipnyXVrE/K91N6gfV2SbECFGq97fAimGFbXOkkSBm392bfwh9N/erE
R1SALdlBRjpnMMaxV9jtBrjiLUeCu/IYF81RxomubCp3Nof8xfnS732SpjdAQl87
Fcy9BTgU9v0iMCkdNE+8rKC9ApKuuTy5gdDl+60H0sQL8F70fD5g1nZIMVfb4Lq1
EGC/eHkpUbqFlIPo3SZwHhXhsqmmcd1GdkemRmosqzLWTrqi9xIvPOdlLHB6LpTx
TPED2zi9yJ4OWmV9UnPBBdfrgLeuNXf+VI2evj5jqAYluUMqUnVnL+SWKBzTGW7i
KvA+xSTVzGdZ5MH0rBdzcpkDv3TmnOc4Yj0ggkN333EF41QTfBhAZ1i6YCoPD8xV
2BPZbU2iEq2eVH8mczXS/uWdGjfrFvf+6ccQwYm63PnwV6JJP1kEU/Gh42+0BjQH
OgcOORRUU/fAo1mnOHGzmxCyaa+3YFkvY3Dj5HL/D1UzsbgMv455lpMWnTPcrNXW
hnogE0iiFTpkk5i7MRGYxB9jQc9s5ZqO+RBkeqO3SRDo6/U+1vryBYw2HoPxfZY3
rx5J57jwJOMiIJ6dgvB280xBcmKWHELXLBVKptVPURf/N2pI/DPNKhyMNjdOnwz7
BICmLwcvxfQHsi6UGu9vwAj0ppJq3+3IRkwnW1ZdO4W8FPhG+96OkfZTYJjO/x73
0ibvfnejupDN3zGK2stNHCbpjd7egDUB/vxoz/K77j4HwMCRkiKGvF9mKruG2pQb
2zebZEKPBDFjC0WaTlmGQllEq3vPlqtw7GLVoPxiWnm5DeMR0w0JpwzSgAD1wgWo
xd6Gnf2F38Hnx6cyBbU1nTqckqHw+z4ijEY52GM9mOnE6tm7aAajzHZR5HBvRX+p
hJeZZyVFIU47EgsNtI4VAIpHgnc3Q4kmLOzDHZJa5pc1hyDZV2rMz69cKo8e+tQ8
TKZrpBfWizq4F1ltYREA0NHnZRrprn5zD1/u8lC0TSyLCu3wNN65OBkXFLToF04u
AYCaaq3Kall+jUK20gOonEQmkuvRUrAqmmSK6/2Y5QoJEyzwcoIaVXWRPIw7muNY
likKT5xF0UtKcdefArjDMm8f16yIdg1HGuLj96FW8MNvaJDiCj8ZLNTx363ntrrw
sUb0iA/i9bhnwq933p8YYlcjolkcp3mJzetRF9Hw2SWufVwAabYEwcG53w+/OApp
IA6wBA2E8nS2NMHOrQaG4RG6f2YRfYXJ2f7TjoTA2JavClU/6G3IcLlya2XBQUJe
4GeNyRdpBUSv64bfqyEbdm8xbQXIXQYpTJuxKb9mlD5wpoSGidWSs4CU8qX/S14x
I+okpg3MAfyMHs21AjJ01lYDklQOcxlFE4yxHakD8eE9ikdfn8BwNP00fQiNWNxc
WfCbcCt7oVkbCGBSTScbBgtijgEvCvxY1FyWHJSq4n8YVHD3qRUkm/PObuKBf2YW
MUU0a0E7638FcAY7Ru+BgcFRoREbg31BrB+XjoBt1D9iIhkIsiOQjVFU0GtJOW0A
GWEKLuOJubh+QIN1+S5cRCVZcIZczYS0N8MPYDFUbbGoftIvbdZRiw9tYkEoAux5
LnUsBiUUCVreTEcIPFCbnyR/jtqdjhdxrlr+XPn/P6J+Z7pKTjNCXGZ+qRjHZCqr
3ZbLK4J1mf3T5JcljUWpXHA1pNZ2JocxEeZ1dTloS/hYB+NTr8MUBfYECpFwTHDJ
fUgukrSFcZmSiDqiWFtncUGGhvROqR/1Tn0f0y3MmSSZT6MO8rVy0Ssm8b+pT0Mb
5GaI+OGNw5K2Sa1c/5UQMAw0+G6rPwy2+EnaUbmHvoOy3IYSGlT+VmEeyfn8KgT2
4tqv4CPXjBQ87GqPbPoiIQf3hMWaKXTAX4WTHzdZROaumZ940dVNy8YO9GffT4Mx
a1SPvsQ8dCirxJSHcg5R11olXw0KZuQyyRyi3fqMxo4Xd6ZVajLmPfNlMhxdeeNe
r8It+OAd7fwlekOwTLhUeP7qXi3Fj+u7qOY/fqakEvZPtiC5ISCKcQTIt9fJHoYz
4oDdBVPHSRYS8r7gBZJQ/CWovbPm8yoaruJufJLVOGHbfxqIaGXZsVMkOdkzVIXy
fEZhgq4MHhVd4XD1otLjzw9HmWKc2AongesSzwgxYXK9njcG2vd1iX9wKd/Oqsco
P/0YIgZngNxO1E7tzCUIoNONuBGKLZ5wUf6Wh6sVVpGUvWvMqjUi5SfKMUpUuvkt
XToNBQ7DBe880euTpaEwIZ0ajrWp2G2trxlveOmhDMj2GJ7b7zC6wJL+SfQYfBFI
JheGczAEZHp4ZgKMKiwJZbO6FGybWCPB2T61VOJusewDqTuXK7LhD2uosFUb7NLc
iYZJywD+NllANyGPJvSMc4sxvYFPlRgCphQdF8+8OnyLL8t9yERvhW8XSGzojXnU
FtShI+q8FKbjsVc0IhOSo03GhWP92ZDTmTB1dY925ybbX86TBFb4lgphcXVDH+za
EHIUJ+xDr4+fHVEuZo4lbianOwSBTpsV/it/MLYLXDdKAGuxJAq76OCqpBwRHjea
Vc1IwY6iC+kTVN2cvepN4l+YEy1dn+D/9h1/gc52iPahpKjqt6lU3bANBCFnstXX
qliYiNbQx6kyrJyJsYMRZCCTVFQL2faScvje5dXn1n54tNIYna31csX9yKZY/Ylm
3l4T+w2KP8WXLXdVtfgLg5edZfahK2xP8dRU38KU4pQVQeO9s3T10tHqBHjMzOG3
HdVU3Z7yypBM+208dtNj6BBXW5okIwvyYb4ooV/CYWps9yQn+dXUH3dEXdiJ7rT5
3uXTg8FgviBM6/c3pdf1bi452pz3IPk8KqaCAlQPKdF/ZLuK6bkQePXMxn/RbRgG
XDiFdJRHU++VvewAKEc87Lht92jg3ki8GjTTSIN79mGWaI878g0Og3sVdM7bhR51
7r4kngViE9rQaBPt2OSqCQljAqF6l7JWqMaPKs/xE7D8S2ABeVXvGP2UTx2Iwvaq
qFbd6xxuYNkiiZu4pLpqeX5mGPYr110w/0ikh7l2FEh2x8P7JU45JlwHg/I6LB+e
Ya8BsrSfv76LAM61CG3xcmR0+xtsgyeCuqFqHbhxKvNyfGcGZRnBMPKv9BAxuvtk
EzKSOmc1cz/2zZpqFzGi+u27oP4E948NOKlx871fJDHqhTsXEB2iwfdH/QcKa6VC
vfriBOZ9AJP85RqTIM8hvldLWybpraTc9fBYYg/WrEpi2vQBDiFCVdbQrXpP4OxT
QwWOwHDQfQ6hlV3YD3mjI5k1WTSPtw0MuAl50GxM0VA4PfnYh47h7a8+f87WOCp0
zua4wu2TR1KUkjXLrZqYJckeIlCuSqgr7e8cJC+GV29WMwvBeiIcCHGX+Ges+PgU
uel8YIdrtEA7Ixk3PcBGLrl9mJ6+/dmg5/llZOVWNPvbPWWwuy/j2mTNmBYBkhU0
9pe0TyPUbzc4b0lCjc2YFZBvukSFDqLK8LnHCZrN7EKh8ucex4upzn5whJdzcveU
U34I3ib+ATeiY/p4/DDygMb5EJ36+LUvFe8uDM9JunwfVF04zTWm6aVJ+x21Nf3E
686txG9WlYSZVk2Su9AUO+htCTHgQ3IYdxiBK19sJYgicwCHIWdgp73plT8WWp9A
XVg4RBXj8cTu/rq9jbHXpBNGopgzdRB8bXOHhp1thT6UKZal5aiFB6zx+uu8F4Ny
X0ITXJ1Sp56FfWvAPcvyp6L2Ya5aRm7fH9l2rX3IlRuLgHEnJ4eJwBD+gVXTXnGf
SRzu1RWXMWGPLPLqTOaJ/I6v6nvfl/XQH/ORDoJPZ4Yxud3ps334bakm20I5kcT7
EscDdvtq2AGsqdpLjvqo06BYPXC8AShIfs++QUoTe7nrOW9DaTtZ4MKKHN/nCcyc
ZGGTgvG98LLOeRUCOIAsycaFb48N/4SijEIRzo6JaDnFBviH7MmaPyNb7r1BlIJS
R+/2YiGKUuTNx0qdFZ/jgQ/QhfLwfMRjEIa6C5Dx5mU0Rs8SWfcatk4PZ83o0hsQ
NGuZHsQ31bdzfGsIhI57nBYJrY1cw/6SIYJpRViiwWFoqFELJB0sBMSzWf7525Zo
dKGTAU/w2SFU/Ax+H1s7tmlugvs/b5g+4tp/KhH+mzNzbUMrMs4fVEOqsMUZBfA8
Sl9QK8CFZ72axueXYe4cYpfKtGzxTetjnahRzmetsQS+DBqh24nv0m3/WVySb3n+
x/lHhbdTHtvN3VjUWBK/j851pgRkSqP8cfbvI3ErtSaKT+lGjpDSLEE6GsCYd045
ts+vOyZrXWaybeh+RcTBAnPch1FAcXnpMckhMcNWjtfxkIfvMjppXynb5L5DAFlo
poSAa9JbJLoobV0Al4vXkF8EkJ3jYjIPv3kro0G27jZH3kunZbNWBDH93+Lqik4j
oYvZYRvNcm+8iQyFOcF4h/Y7b6mdAatnNjjMs4uzMcit9SL7HfUeHuBGEnJ8k3cN
64aJlPWd/4jQKNio1cfCnuRZ3tzgoxnTOFJYIFo4lPazsYrYnf6EaT2GgLYeaz0B
gyjBC6bFVtE19c3cfB8dBfukNJmrru0UftXujeODg6SgoUT62uWN2qGypGJ8MscY
LpVuJzdWQIuTramzJxlxt1tpa9RmnCJGl+ABaFsdBaYGdzQuUJg9uDOpX1zMXOtU
FlvtKXXRydGSglOVKypgFHbMlvsWAItkbTIOUkmfuirBGj28PCqhtjHs6MvvB0XG
CzE3YTjqx/M0w2HjTVr1Wtjd5MJCpvnDGoy9R19bAdWhkWz4zkxxjKFgTKc2cVNF
rRBd5YgceKZXn9oH0y47yzSfdOYdFl3WpzJ21PQhnbp0xP2DDrkZdnnuFb15vdCz
1g3QqO3v3bVAH6hmqKPivWE+ppvbKQVMPALo3G4QoWIOizhqjA35DfBgwR1E03J7
5ZEyc9hEYyp6z8WfMubUcabkBdaIUK7rbqMEYRghIIllB+JLkdUNLg0OO2p2pVhA
jvYb/XilyviwdLk+1oNDRt4F6MgKTowLcK3etNoephb+hZwBO82nmOmGHDq5ivbM
l46f/xe2YhXNJDE66xmLK0383OrEloBhyHePWc9Kg5kAWk50o4n0G/8KCUDM4Fec
u0I7gXEF6dOKlCYmO8HEkMpz589qVU+nV2RrD5CEeDMLPq3UtyJ2bwLQBHpe6fqK
wPHF1R4r4CzSLfGMQ03p+czxKBqkj05PIqgmzyuJZ2CKFHELvcdPYuTpouaQ/g16
D4z3kmDwCzvuwtndrvCPYNtsTEleMTYbUGEBjXcDImo+l9Bx6OLgwrU0xMOjrE85
wUnBnZ/Woid4Loo+HQfGdHBoZI8fMCMdBTcbAICBlpBsBlbSfKIFESKzeGMUPYub
+/Drk7Da8DE09V5bXUeIyYTCXS3ej8ldpE2XJIrnzP8VWC/wxnj+WnvhpH2x/hTf
sKN+zVDqDrg8+X6MLTrJmdVE3WH/viE8UBmX4VIyMrArVM6twajG8bPN6FTW8T4G
QSyKcorTVllS5iTytA6Wpox2wn9NOwOYL/FEMdztoWoVL4gmuAy/FMA+N4jMjRMD
fCZHMMpWbcqvhX6B5Lce/oxqatrAVdt0odcuaw2QcZRogYjVwCwtPlqfjN4NS2ty
t3W5MRTsRAkz59pfyREhB0+u7qkafwZDylO/ldd9Zi0jJlOQEDGQyDD4AQAvyECb
rgh/VumDDXupJaxWo0U6kMGv4k8gIWNJOkV1MgmYCR14jcasYX8VGPk5tiCmUiN3
+NqMPqR1YAuRgLkBjPLqSflkf0S6YC8wQ15QWPDXRcONsWXVwh7+ywTsE4760ZC5
Hl+bUSrCq6z6AKld1EFv0jQ1Km0VIRc6RKtSea4FdYurnjbm7wljNeJnUAtIgu2X
F5V2MwIdzMgh00/El68TsbwknpW2dOgusdQKr8JCUznzwHal4K5vPmcAMM5tBOWg
C3tz8nX33ML27oMAMqmus9OZt8k97iHwuNGfWON80Eh24eXK65ZqF8nUpj/iPUxQ
itLE/6tcGdTv9G6zU7V2jNZ420JNTPJ1pyRtesXZiEHJrX3wDGj5WE415p0Ctfp7
JfScq3stBcH3Cl5kQpDBYwLFKHaI7I13i0DUWXaRoPVQI4FO4FmTImfF61mrKpCe
zOWqQNLXKb9jHQadGrhVMYXCMksiXFE5XWZqTzex4oMrJd8JC3J9RhY/8n07wkXJ
bZtoyeu5IXCJ7Dw1zmRymyiyCZM0uOIOdlEA23qvF3S7+HprLahDSAoqGYlwBYxf
AG+JrRiqR2AFS9hL3T/GdrTABYmaCYvueMkPv2fHqvD9b/mt9jwY8mdb0Ivpeu0E
puHAOcFP1eQb2MbqZji9ykdF/VadYzBsnD32wEAlDXzHqmA7dufblf/nG1fLyXSF
V/MKkJzkSx2NYVnUb+vaczXskggYWkez4wyUTaM1O/Qf6FU4KXF37th1rAiX6bRY
bjgKgLyyuI+HoSGGpaepYTx8QnyMPS0uaeo/FF1av7Fh9+FL6ju5OOhpSuC7kohd
z16fKSQl0/463QW9sO24fXk2+cziCR+LLGbXlwvzpL/b1+6NNu9hsF1WsavxlAqW
3K5+H5369I9p5uq0qTAJRy5RDm52uZJSzly6GAc7lYMVh0Hmpe8O9z/UtSLgxjjg
VLurir2bFwpg7o6/Wjgjx4MyWEUyaREgNF20DzEO5C8rMDaEFyzaPdi2RVQqaIKq
MkdpFDMUDdSQ6VqjLRqLpsEX4qQEPlkX7C8iOozQum3QSdSpAX+T1mFwppQ2uUQY
U5khjgRKyH95MpOa8liYHCIwb8CU61xsL4mIG8yhp1f8hSe34BRdb+eUjFiwbppo
pRVD5lEDcmjnv+mc95R6jl1xs6YpP9dpzt3MNwQySzF+TAW8/0Gf9fR0kCI+0ydM
PNMhajhHKeqEr8HGiOj+5FBKnamy9oD7nanlBqNgfD3/nVr91qGLV75sEcQXc+G/
LI7Ul49/hQjO6UuYYEB/rZ/b9qSO6bJCUvOdRx2c0E+OR6wvxfGK5ZoOGyhXvV40
PCSzZ6bjgSg3R+/ZtpUcUq+e236VsdXkUvow6fhA9n9/oBJYfKt7pupdu6HefzFh
ebTqRBwEafmrBaUxkDsHc2nFLtqR2nRrNUnulcXvpFSVKMQ10VSwaY9WySeRvrJR
gApN5VVZwvfXytjcC7K1i6M/Ky5V8mLIIoLTkF3PWobI0D9pYIFOJiJMvwXopxWx
nx0gIR8J2l04R5xWpS1EeNufat6nFzswm/EPuVH3ZbhRcyarLopOwUX3MPcTZ/dX
sdkvMZiFeztjJqBmbQ18izyKFKvZH9kjEqkn3rp3LwJz7eAlFUxyZ5VhhGfClHwI
sw3CgO3pvznuWDkvYxKpkQZiB/fQELUrHj0e8Adp5NoQuhUnAgc7oDT5KA8XEun9
dfuyX70g6RLBNMeDYRkut7oxZ37oiSogFwYKyViQ3P3iRPfxGnl+k0mRzj4y238Q
VMrSmrNBSYh1dPSy6DjNcscbLVggPvSea8HksL3dEJMYnAs5MbIAIDIHEp3iPFZc
QZcLv0jB3o7cuGoG5AHS5tdC1/vOkWFakNDoUNZbCvW+hwqdIVA2iQdKeVtao0+c
K7Hlpcu/D0QsC77hYjRcr/LBiYZCXCu59t9+tBABm04mnZl5q0RqOxIbPNePMcAM
qTfbpTdtxdFQgsGaoGTudigUE/OfDb/uHVNcSPH7qybg4xWDgxdWInLMGT88UocT
ZQdxxqQ4PhoPA6WSHhEoZiT3dTSl5LjNtUD2yhcMVZeY5oD2+JwHk/yLXnRMn+uQ
hGS0qP9I7Cq0Am8OprZzxzCD+NM2q5dgMkENGggYLtvYMCsjFwf+Cnhvc8QWNFk8
bJxaAwhVgOTqmFbcHzNWsprJb8brfNyTv7fDgkRd9Je1hdRJuTz9YcxTs32k0hrW
MNnGsDd7RPN66mlEaAhZ+IIX2LZXsy/kwug4HOX+lJOL1wKxRLfQozDFtyUVR8dy
Fp3EeG6j3iowS3Hak/juQkGlS8WPVCAfhKvHxG5qU7a/gQ5WDSw8KJBx3BrUM2Ov
MBwQU2eeiBeLpdVOhc7L0i1WFhPu7yGcCKKtY7s1WyfioouLPKjk9+FBx8mhGZ7a
JUx67Ancb7DX4bNjtV1rsCSI4vO/anGuiqFncntkAC/oeGSe5mBWe4ok6gv/GsHb
ExKX1CcYVzE6zrK7asquahFM6rA+E6Cym0waVl1MPfhlnhQP6HY1Tl7su2XzdUdz
pgnEOdptGLzrTz64nEONi4DMw5BhPGmDi3HPVij6LYEbxb4o/aXqOJFwziS1xuuT
kTgtxbyCZp5dyBPVpNvZ1cAe54JtmYyY1V1JmI5w7AmNwxLll7M8kQ4fwYEUsRgp
q/f9NfzoPUfKbxyb+YoXx7zLnQ79QrzURWPCg2a0NZRa3jIUAiX9CJJpeJ1Zr2p2
HpvNbYM8xbEFwM85xVHyubPwLtnh6R+KePc3hWNsd/BSTNt0bT107WFNrpNV7D8O
H0wMM/eddksUrauBaTNmLfYDRCiUQnbAovcGAmoIXtq2Nz/OiFrRZHpwU2QEiM65
QQypkW6gLhIyjqhjEGRFq4KRRYC9RmMptgsvRk34DBjCiFMTZg4pYNEzO6VWMRF1
KSGHDKEHVIv9ZAnjZZqyhi3amxwflNycRx8ONVmqGXuyseMJRRa2m89Xxfeh4Vkt
zHnyH5RgOM23gbOVXqnBDJQFsTUARLa/S6FEngrG6SX5RcBRoGB76cBtxuji1Cgq
canMLColx8hUgF6Hl2XE+RcCMX4CVoeAU+AGXDwYmvzCtAHkP+az4licy+KuBxww
zq7c/RvAnm0AcD9C4B1ToAMSurBVxQfi9cg5VD/SdmkPk06UYBr7bef3R75X5ajV
w+C6xpKsR6wJkRWz31Ol/Owqr7ZM1ntDFQbmTs+sYUK2MM0gd8sx6YMdSMcRaC3C
1qP2BQJBu9NPB47tJLZ5DIvGkntmEYGvmqIA2UuegDqIXiTnYWdtypBDjclcpKE4
Iyedd8wcBLIP0rZ52qtC0mnh0MIKudwLy8gjJuTLi4xZTg7SZObzV4VuQu0SiIO4
k514EPdGrIjndGdvwVho3CI27BdSPn1GRDQbCVuQmynat5L1tPQN9zxjjIBlr+Tj
FxwxbaPn7+0cpLOcSKW19pSSPyqWxyIpy9MXhVuTI1gUShENIbp5ajg60vLnZZ8+
LtpBm3FKBDneYucVUMgmthxHOS4dsm+bNFsW0P+AbU7lZA5sfEyWHZWWvjkDzG3P
8RqvT/V16kA3id0oJopPIDQS9uxPIXIXbjfHaHqb4/qgBsuK8TH2bpxi0EmdbzwX
QQTphiJtdhUyg4+L+/GCcfjAAIWpKeOL1E9Mtbv5GvEuEiPeQJcZmPJyeBuuH41j
YnlhKVES9br/1HCbEG4WnSjF3RLqQ8QX8QFl1WB6jKnwzhoXDFrcwST+0E1ccko2
tWga/1Mz93YjkpPrm5Umg9doVd0Ztwgm3KVNx9w7bi7H5NerHpcftEWcmGRnZEPA
Ojhfzx7bC+O0SF/r0QwfeEdTVaN+SdCeJ/shUznL2y9C0cN/QMB22EO9b9ZNX6Xh
zSTIs7Ltu2bueB+aukw8Ltk546uMNwa/PbWmHEsN6JujVw6+gdl5ymavBC2wOVq7
eoGq+fn1POsAdDU8PGPr/+PbE5FRwd+vxFKiWNowmPSch36XGhAsbeOa8nOgjt/Z
7NyZgao5GhkUI8R9y7GsD7sfsbKu2TeMCY2GyFVHRm63M5Q2sgEWIizbe+poSdfe
2agQSdCHqjc/212gx2DuO9vy4lPrMl+l+D0dbYhEjS2uJHr8V7ZFx5JaRqdl+zry
NRtxdo0YA00WPos0Hbh43Tqrgj3nFzudrwDTd2zuvULOcjdGNT5p4Nv9E62sQMcZ
DElQGRgololyODa0UroLR11RdSLQirIFP+yJLcmFBKEwiT0959weMR+modmzkzu2
lq6/x+OXAuiaxeZ6AsksDx6WjX12Y6ZswSGpR6mN/dTDBbv/HMsJDhnqG8NsaSgJ
dI2DNtTCDA0Q+5+StxknMbwnS2r82dIJ+y6dUev8KQfscCdYKiH+3xhxseCooVFU
/F8Yn0ACX1CBPggOXwAM1OgIQ7UKBBh6CtDem7bjHkdheVXnbXifKMTk5WXb+OzX
pnlDm0cXJiyFMLorY1S8Gg3Un7BUUw329mDrPWOHVPhiZQzNFH6HFszdZBlowBiI
Q7ZlztztNfB29BmK20A4JwvmJPJ5XQd4InxYGeDLB+ciUvJgCbCDF0D+bRcXY+09
i/TmJOKZSBXl3nFMpbonc3ZZ865juHVa6fte61pqYW4yYMpuNiU+NwC57odoW7rZ
z4Cre2l4D/v3oz89z8i005T0xKe8o1drgEk0/YOj0VcW/Mq6wS4XU81u6X8Mzvbj
Ub4sjwcPbLQVSJTqrMsHSXrLhfDJl3xl7prEfcZTcQvUoe61w5v9ob0tA52CMd2q
tfTfI/Wi7VvGk15fpllPjvN8x9SjsvN0ZzwLjA+VNGGwd1fXpVJ/y5XyNv0fIkik
hIBviTJwRh5Bb6faPUpf60OTrq+6GQYFX9+0r3gY5vFY3TWAy6xRXPDEGWZkheKS
Qve2hWsHkVWmrkIC9i9mJoXvOPLuResrfpIl+DFMqLRF7IzA9lYPA+SCbMmqaOfb
QGbBevwM+HCnz+cMCNIV59MnLTYPaPh88V8mt7hpswGW0WatmT5QWk0uTjPZ6S6Q
j/JqSVTFSdHG/WfTJalgeni30lyOueINaVgzvqUejOilmpx/AqC7DoruOOjsIQoI
7otvWLXuWa+A8BQwk7S35NfmOafwGAZpVYv2unefS1Mdyp/7QfiZpD3+TkXpVdjJ
S97P2XIHSXOAH4AiYkIE6qxzJ+dHdQd9MKqChagQb31qHs5dNpmW+5+zIwXpJmum
dGkaJq4/WOg/bj6N13e4PrLmqV3TE41F4LnzRvGmEM4LCYJuIGMIEsxPeOyzgPzG
zYHv1WKtBQ6WuZA9kxVFu02xbuZiPwxdM1Foq6AniPMj27+pL1XvPa/sP+KN25qJ
V/QcOkn9tGD5uMSPUL+J99djXQ8v+Jn+nR4MXYjFZ0Uq3fEdCPrnkdtwkxZziS9Y
P/qz4a61OgFZd9SdneKAjBmMqYqg3ahVBBV0ZnKGW5dZLjLtO6DZmvcpD98LtZ95
9OFG6WE49FXHS/DO4pUl4g/fgILhWjBOtj7mnU3/heGdR2JsNxLTFfzXjZBm/QcF
uaGJumvzFxraQBsjOrifdu7TVW7ldsj9OE9mQgor+2OHOzgVqqsjskI2/wPjHQDE
fhAfpEGk+YPUOvstBdnIorMB72nIM3vH0A++u/N9k1ocYM0P+d19688dFmYJRi7/
2ZKvBBv0Q+qiDOScoGKayc5FAL7vhaUJVaDfuZAKof07viJ4vCMv9WbKKeIWqrUG
K+KV71HeyRs2Q3Ngw2PxQzKvWpkjyTYiKpo/x3CaqBFmVVDR2BVIVGs3aOIMNOsq
eOCsTo4HNNvFlGb6lfWCxsroyK3gTlfTQvEe/k901Q4CCI4dAOHe7syq3lv8/yYv
cd6mOmIiP1ejOHxNKhX/u9IxDTvzR3WSzrlABYfDg35IVbkvS+MtY3TS2MQYK9Cx
diNN4EssHEWzO/4KIUofGXINMLkHK6fNtfx/gFU8THSToBoCJ8TzAVzUkKlRgSFv
EMnWTaQDtTSknkRPdRwF6I8R52W6QpbmLCQ0Cgj7K/pDfkoN79IJ+KcEuAQQ8zPE
vhhJElv5gcNCatYFjs6kCU2hVrxAQgbOgZh/P5+7WTqjz3Rj5joBiT2QHeby6Gxx
rWK1XyLJedrbLZ0lUrLLDuVwqoZyz46xIuGJRKiDfekJimJPGkxqqgbgWH9Rffmi
JRK01sLVth4C81kzJokaHG51C2O5mPsiA8ihFJWh4FUgdkvrb/xYOwZRVDTJdqTh
1JgY+8hzSshz2qpTs1PJTLywt7O8qcudvsm0yeLvG+Qus/m7FWlzokcJ0vPvSyAc
7Yp0fzy2iRacTqdSHGGuoGfXMwpeNDhcU38pSjlzybJxSIR1B9GbJIFoSjsnruRT
dE1l0MXo6LHOV7pwwqx0soaTmTniF449z6l6vk+DFRaEp2WTvDYstGRf/486oTDy
uCS1x4GaSNDPayTahbEOdxq7TslR2aZgBxUUprHQLIAZdoCc/A2FQeVqRoCC2vyv
2MrlLJbMnIKrIvV88GigWKmtiqYk85/oY1nUFc+92XCjydb4pVeHSZwxDZyzP/is
zHusO3zs5ya6HGveQ0xMzjNgqQzVjWjModoBqQrF5Vd7YTlfteuPH7y6AUE7mVYA
zkK+g4/8xIEZvtImbpERvMWY/vpbUumykpzeBiffe88ZpjUyrxx+W8GGGlDe2aW+
Dw/73qO16aFyi0jRbwzDOM5P1AyAI2c+xj9nq9A+e2og7+fPQ7/fHgms68z6xEIw
Tv+mFfKL8oJlT+uc7h7AWTCbtj+UYL1VR+G3pkrfBEgq54MSyxq/oqrKj34qOtNW
SrJkASdLumSjFxbJmoGCQt5CsS+cwd2n7CkGR2LVhrMenrUCBGsZVf3UfT+1fkZh
fBV3zpJ4Xen2e6mgzjrpJ3TvYcgIQorYomUg2zIwoGrrkA63L9F3MeHwnBvU6IsP
c1LhbBpRY84y+IE/YkQoF5i/y7gpLbhMY9nyrysA6XBltjs7y7bkz3YukALpZ3LA
cyfdcvPb3H4FEtw31m6MVZnwOOH0d00dISY9LEHqVrgSX0n5tsp5nS+xcBjmIZkh
k7e58gy83k9vhbChJG7HiZ8BL779OUAV1dsZUHc6fEeYQyBzISypFsZag1TnDV9n
JVhiy4zAL7vdFeIjVCrd1RYnInPxJs/HvQ7NAs5qkjIFIkanp+jYKLmrzot1eTUa
ylx5E0yS3raA6TwfsxC4f5XVzYxuvScqCX63nyRdOBqzJh2S2LwccEVVxl1ssR8l
s7lMptxilm2cKQNhJWCr9t6HrUut3xcsR66SJ5+qjx3kV5N29xojwrPlHpCyYm/s
RCmfYK8PC6lf7kczNAOU18Dg5GVw33GOgngjw9Ifhbqwe214MQ12DsaTLBkV37hU
kt3WPEX+sE5vXp7KVZaJoqmHA57a3swaR/bJYn2C2IHgrFDe7020M/gtmUPeOCCg
dvUtidqb45s9UfjIPm5yCAHqvKXSc4OU9dUXJMDxMAckZIAeyyy/9uQmr+/97LzP
4h05l2Jkh7yiaUMV04tL4VvGZSmHJZ6FcHdcTs8Guy90JTvKTB7xedRmYP8Ddz7V
3taXNSY9OVBuwIpJPThwyb1cJeTwLGpNsLozB9AC114Sp91c9u8D+JS1KV+DL+ZT
N7/buRY53tz3pH8vGJgcqWJc0A9NnCOnHLxTyQ2LcxSHBz6uTw0O4ZYqBipYbr7b
pNo2Zsk4jNLLw65Hco/Apsx6xbzqJ4oKwFZu/B920paU0ReEKJljYK6qL8sPn9TQ
VLZi1gB79++DCxYTQOsCBR7lSaIUbQN0W7vknxWLUhs1wvHYiXBe49eASr0a9vi+
nvwvMFiWgrk5GJ398GbAJ7+yhY+KNONC/AkpXeBMd+jHqqTepdHHEFNBY0eJ1fIy
YvUHD1mbIyLAeHplMphpo7z9fTPOQWuvfJcphTgR0p2TQzr1R2/AO9tC1dKeBpWc
e0lYIi0+YnETSM4USgGM7AEEfbKHtsLeMDE8HwaA1UUQOzlYPnG1+mLP1bsRS98Z
bjKhmejM9iJBTLyYvjipV4/AUWeF72fkz0QkapSNjE28Rmlz/dbkXfcaOzVgWPq8
g8iZLKP4YJRRvjUdIKiOnCfXgTVCRK4RgE0xZ5ERLHKF/t96YXo437H5LqvL1+3c
OafBfxSQv2xM9kZHqPq7MbjHHq2x4/weOaZrbRblfuCW/zoTd/zX+aoF04se6W31
vYtutY5KA0k4thljLR/X4qoCjItZhHecMG5PXFNHSqCVyb34vwuG9N5JNNCeUCCe
0VEXYFjSHzQ6hmMzB6DVY+/D7TugwDXbT34ebIGvOpEPnu12XRNW63XjG49KnuaT
uZQYNbFJrak6uSMPRo8xzno75rUNKF8g+TcuH8WshAS3KlTn7ZZX+CQuc1aO+/WF
DfqzPqsvsG+18y7pGeEoVVg5jtDUQRTgdBRaCfQ10R7f1HnotS0tQH0SsetspoPe
mEkQePRPi+4dA/w3XNhH0mSMUKHyy8UgKfN08/Iyy4+Dr6c5DEnO00R4a4RkvzKm
SLILobvhldkn51Hcc6wp7kCDK3pAPcvKFOaTvFr6cWRD8TAYWKP502CI26yzAgT0
XEoWwk/HBKTBzEygPwIRls/s51UHpXwKnc2JV1GsX7C7794Xdw/P0kGo8YtfeBlu
Sc1+Xw2tYtvPOLfax2IDkC5ZywJsp1cIiaQ1JelYxlgHDp3Wl98yH0ZsbxRUtvBg
ik0H824YrsfOkJkoqAAQryOD9diCDIXhbEjTgq4srf7ZphG4mypsaqGrWsy1sKvJ
Y9rRs8nU8OCNk0YwqS2fIXzRUjPGCzu1jgjRu4rSuLbb83im+In1vJkzjC9DkW2s
fX3N11Vse3wwAcqdMPRSBxLd5coBDkDAvJXbgi9B3cgCqcOA1ua9d6h3gkmyh4s8
NFEnvxxmxmZVudbiWwSm0PL2j0CcoJF4yi2oIZP+VHZkYdyzBIjzgoC2qfmuZRkb
9W1YGDD94mVj2C1S4ZcxhkqtcvRM4Pngi6rMAZ1CsDf4lHGAwuo5pG6n7vYNQDSJ
OAiLuiU1R9AR2rY5TYTN++VOmy7xSgKW8G36aG2xBbHLijDZAVEj3fN0wSgdS9J9
sNxUj1TbbzrFzUB3f9bpueMhfAbsRTxfevP561KWQzPzQOqwxMkqC5CldH1aR2Iq
+66ezR9ZCd5fz9oIwrbP/dLNSHNNhE6DGkxOQYGNhA46Vmbzdj0dJoOAG9grhO+x
i1dLBe11PVhww+w6hO59HEqEfXnYbbjnoMSyiRjQhucdq58BRgZheJLZ9M7nOKGA
ySL8t46WZOESOrkMmmIdnqEzIjK9jnrUYDZXgqKq16cEyLufrXhll22sWNiAG4Z3
yH6Bo9aUhtynwKiK0mkgarsKO8ZkkV8D5zfcdH1r1KdStt6pgmhqvchK+S3wpdnv
gJCR+MCNrRPPvji8rOLcqexMLI4y7fXwPT8vS1ZU5gLxO6YR4qJq9u+alAo/79Jb
09kDWldclwUWjXTENCeU1tpDSta0Ssa+u9eyO0KkaNdB4zp2PsfOQC2gY9dTktrt
oQgC1+2Pa2O+7Ip/SwY42PMX6niexdiaLpefC+ot7X55pg1js0vtKyGDCa94ZyDQ
KrVWEc40pFkFuLinmN/0napK8MfqHISrvZ9a+iZNWmHkftiaUj4gJOVQAnDfUTjV
Z7xgWf+R37XDGe7GOKYtEtxml7zx7F3bmtO7nRDnQxH0pTrB+dWqpkJimdoNL3rT
/jHM0n6G+uY/hHOGvFAIrIqLhLhp27xNwXIv8MJdmmPjkk9RDY0857WFtJ1wlFJz
kq6mUwPIBP1YnEqYuu/S+t7AQB+r/GdBi9tEIk6DKAG3KcWU6iCdnMpc/oT8flbq
khhH5oVIZIJ+deiQDln9Mlwq5obvmyfPfCrsPGHx3DKImSBdmQmGfQ5Y9yr+kR0W
4OtC1aQlk3E0roVx4pAKJ9b52j+gcOP7EtQSjRt7JVIsjsMHXP40Ey8ojnOVPRVR
CpmV70HYbJFRPa0obQN7t1vAxE9W0FT+C7i3JZkKjWAPTrO5h1RhNTqBNtUdDrxa
c0Y7LZCAXQSLGvZUIDpUH4Kn+Sh/8TZWl9cThe6dT5yp9jHU0xuFBs1Qb7B+ZIm8
UEgPKcG/9X1Cvy3RY0YxMPbu5JxD4S7X/uUph3rOXoE9pO8AUOOM7wSry+5IBz4R
qY33ON7Wn9irJTIhWqNg6eM9XQ3gJNBqUFNVcYtR1Fb7KCyyKHCvG8mfiEK7DGjU
VoYu1o7Fh5mjiXw/L6ucwApI31mTBLlThHmBc1bswWk7Q3RGDhNewJLFFRxrJ0pK
9xEbB3Lbt35zyknWA86ZVibFhtfeTryqB/5atanClRzh+3wxVuuVCXTHvkydgGzO
YWcF9s/pEZd0JXoFnnb90XLZFbH9ETPrvz5r+IawqnnzT2K030tcnIv5qmZbVcGx
mSPahWjpQWgcHRj3/7Zq9XLAR1ART/1HvDwgpln6G18af/9Y9sWHrEz5NBLbMLCm
VB9rB1eMvP2uys+L6Sdw2izdP5HZgCuPo8CryjyaYPNHvNSQfX/qt33YTt0hdnzb
QsQMqG7mZRQflEZkXYzbA+3piIL/X5pF10ZOvbbsmTUHHg0FpjNdH1amCcAF45Pd
4T5p5R/wIFHEYcZO83nRtWHd0tgIPL4qtsyUhR0t62AEMVivRsCkf6WlO8NorroF
fBDjHqc8J1q715IlYzE9CDZvtkDqc2NiiLPPDkBgSkzGyBW4wI7TN4b3cuIkQN78
CiEMVlsACRUawgUQLgbrsN5xAoli6/mUlog4GAm2Gdi+0iWJkFZ0TPkrgM955w8Z
mkPdbk7aWODVEIUdKnKthep1gPL8RZLuKqBEkT9SL/IcRyoVgJmLTcz+royQkqus
ZXgG8uo9knrHlZSqQpzICp134HpHLRwow6fo2/H/9G518X0HjdA/0SivtOQAxC9J
aYBKh1K0/fJ2rToH6KE7T32lBASC+aw3FpeQXrqlR5oKcquKArufJwT0WDPv1Cdi
PuFUarDaxWITWdKbXZjzmCYSaGQakYtiTqYkkS2XO4RxhpxosyGxQRiFvMb6ZRUV
bUXhumGwnk+joyHp9Dx3o+W4TBYpK6HZtE1mspv501hlsQA+bZN0FfK/GrEmEJzf
xjJHBvR0hXTSaqXUmKbHCQlkGZSek5ODthxj/EWkY5g28JlMLtyJoy1cpqYic3zE
OtespO+H9vKn43v2zZl3Uz3IKKMUUW9WMtvII7dAuyZwovmbWhrFObC4DskGhaPL
fMR7baYHoz4FHy6fSAdEWKyWYpUSf69odYoMOTpCHJI9whhmwwO/LeRHQU3ux0wx
UWs2SOhKCOm07VfvpXJlC2QEl+BxF1ptt5t6bRPWIED1fE/m1U26VQ51UVSvDRRb
dSr2kLSheKSg6FLzb7shnbcANXC29x+8dF/OMszB/BY2pTx6c5OiM7qWq6XvwHNi
d43qsLN1P7inw0EHtbktc2vX9T3zP1MZ/U9IrpXTLlOp4Uc6tG6bOmW12rNqqQ0h
/leVqMigN7hPh7Zivqpc8itoNJgkCLUQqA9wu0+iKVuj7kSl+bFcFclPh95J+3yR
Sl1ssr6br45xbIjvRnU5pZfn4djrULS2RQJ4wE6aZ1+gdp2rp3LcqAgTQ7oFJfx/
OcJbKSZXQCxGwqIXRLo3n3ZqW1iqfcMUNwFxV0NAwQLfYg7GmB6nBmx5vbaAuCNZ
lwrnS/fEFJAoBkwoW3N0ua2Mv/iP2HcQYIkhQ3y+ZhxYQ6d2/uvhIF+Fg2QYSF3r
RHVhpWdtF03EYUXR1BF5vn1Jsr5O8F7Q2/BkUc7fnq2f196xGTPMRzH7LD4f+73W
jqNavPX5CxaSqF1PYAf/IXQUL7WHJjJxNFkdf8KbYfvpG0utTlaQA4Ls4C67vAnv
mYsJ7DgwbvjHthvlIudlEWuFiULD/3txgyCUzt0pPlZP9sVtoiC+mEY/RQHI11rb
PXKIKtRWoq8xCnBiz3dF413QTYIy8ay3/HR29euBgPtKxDx1DkWIoYA0vweCAFgq
b7bClcWqaT84WC8l2ahf5H/+3VVjK/UatfQEvfgehfJXSpsB5A0N+GPTBuRlh962
6A4JJhyuvjAvZuTP5ry4Am+JtgLrfD5p1/Z4Bk3tzQf7eDxxpOZ/dgYmEwRmE6pV
cbyqeoyQ5LwCCkAcwKqs8EbYiBi/N50ksQaiCbaq2Nct9pSrCckTriwzkFkIhBT2
P4iOoztW1opCpabsKTWFH8q9uugAEYNsSsz1b957zDapEIEQBplxIg5YZWOckYP2
D+xdEhg5Fwh/l3lrXbmGGLih+BcY9ay8uX+USk5gTPnRYUs4B4HcZSjCKWwGmRVn
//Z+o4YgDQs8Mee2+Z9BN9d1nHCEEIAgBBicI6gM4A1vualVhRuNl0SiKVjgnDEz
igAEqp00VLS3xTkCIwSwuTi+KezuB12Pz3hhLqCBy8Uwbcv4VXtYLQvZf7T/tdk+
5Ue4QeuGD6GekNGVAbaKjKBJ8J0ponSv8b+2eqMC2h03EL9fVXy9vxNZw7tFXykg
4bwfwrMrlcvkHMCpCjLAU5q8KimIxztDjk0OSfj8IYG96QTagZVPZSAoNyD89Q/L
oDHDxkAW022+iwRnK4GFK3ksxH3Dq45BksNSvorCdZg5LlxsDzXzqZLn+3DD5tyQ
4ejWDFCrFny5RAshF/b1FWUCEWbjRydcQxTHNkOC6x/lKCY8ca4wnBWXUfHmtcPz
6nKY0fJlC63DHCvEq4cHFis6LQzFNp6+ogB26bx9kJx9COabaUuAzwzFjFDC9vtJ
Z1mZYZ7u/Li+6GI5JTw2kpkRCvmMEfXI3yc555MYs21ck+7Nh0gcTwuizY+azfkT
R4qBl5x/J23F+qnsK+4axT+PiTssWbJg5s2NLT1MdQPWUyldtCmIufiJQIdShEKN
yV9eMOQEvigzfxb1Avc4dh18ID0LUyuV75zkZs5RSDqx2BQaXEs9QSOhfXhN9Gkb
z/2+3NZJgCrJHCo29UZlPuNI2Sg+NtQstJq7vY7jEoOHZDYzf4v2hRP6qYCF8ydu
uqvsWSXmO+ephLOsu3Bxj09jVd6Kmhg/7W2ZBdV0MwWBep8lyurKLTB3BFHDm/Eh
uyiarhFf6ckDcBWFX/ozpolZxPnDSp44PilSIRdzeARqizvJ34pTEVo8ZC4MHjr1
tBSfHH8Y2t+hw9c2/xmyE26A0k4/qEHoMU1clLiZmQukZgoIVT6DmsQC1rT1uyYG
HZQyGjxVypHe6qsCsMwpGbKX4ES8Oo6JrcLnFoGWsUvIquMKHTX6abCw0piMkmmB
fLWHNvsH8QBr4EBLtvMy7y9ttMbSjX7XHl2dmThFw7QR9xhlj9VGuJgexrSbb0oG
5xNVbsrzjkhGeg/Bbogj2TVDniFl+++qaLOkJwY52Cp8idQHauOlA7iPff7Sa8dD
+PkLQH+ON10ZSyrIxZy0I7A2XzNbsHb8BbR9bkbjoWaXF719gJ4mPxTVeVxGyog0
cuRTOfFoiHg+Cjl7WTWJm2RyIuTKiWXBXiR5DQVMt25ZU+kWhc7RtlCroKCKc9KA
Qx46KiUzSGhZZMlQCQ56WXBJR4HhxAoflnBwGl/VmTFFE6XmsxXIu3BsmKgmzWPh
0o7FPYo2xGkncl5zHeL0j7IjPp+FXPC5AnLSU0jQO7q49GDGB1OC2x0hYbHoFm6M
hUN953G6K2dl4VCJjHMCj7a3nmSEN8X2wO6lx9xF2g2W9SN8pIOMXlpASZZKGR2x
lBk43MxgVXWNNUW0MSc0tGC/4KKW+rQz+mKuqEH76jZdGJYPdS25JtkDsJJeddcO
cGc1FW2/ChwY5eXXjaiMmi39IcNvqAhgu6M6BGBSbM3W0/ao/LAFZFVib7C9A6y5
mcFrJrdqV5uam2auknZpsV+x2LybBQNhuA25j/SX2+n6z3SGlT1z1Z7ff5WmI15Y
IuhlDSWZY2z7ctJcSojpGsSG+6YDFLHl6ZTpj0EK8iQ/27umSJcErlmIykMQpGjH
vs7eC2WU1MRnYp/zYfTqaVlvDX/zzWUdAHgEYg7JpFZRCz52KUwomV7mJgA2AemP
SmugOiHqg73yRRqK+wQwnY/wyRCsFfmubqxFOukBLSPn2kEVzwjAexaV8uv9uzcg
aokHeiMr/o+vehQO2xaTKSw5UYHPb0UsWXKX04OKl/HDHGvfqfmNhROe6eUGkdH2
1S02pRPEsi+PbntqeO6hlSN1AtBfylGGjRBNtobwxOEik96qqk6mW3bbrENVVAoE
D88tTZEpoXybJyit8HcO8T4Xv0gebN9XK5aKubOrYQ1DSlvvOo60Ran1zFtrqFTm
x/WGvr0pR5drZR/YUQOLU/2/e/R6W+dkW+Nuns2RzuNXMYTfpC/dnkUbdAae4w2Z
UTq2TMMtZLm0uTvaLPo+hl59HwI/zefcStbEl5tzFARuW7W+rxBYzeXvoPi0Ppk+
eWTbU6KhMw2pf3ajaVUWLWIxsPlsyMqw+mpCC4348lEmdC0oFXmatnuKcgo+Npbl
q3OsiMl6VaztyuByH3M45+Tirz3AUVoeSkAp26alw9Y29LWiW5jwrrAdguIppNWv
NifKD2qnofLH3jJzmUW1ksr2w5PaANBPCTf786Y0MUEw42Bp3qhZC8CVbY7uBfmc
yFxVx9MirXIreZh0AjUYkab8tvRfV5iCTz9i9zaNFB8tnpPktnen34HVVp7FWmdR
e7JLvOZGRTPicYVibTfEWM2UnfcrhNpozsCGirgvg7H6Yw1QuKI1U1hcHVtIzrRj
JHzfQ9kF2yXT5CDmgJvt2H55JaxC0UmtGIs8gL5BJSxAsEq5nKjr/1Nu2JJ+Qr/r
Y0Htzb5xhEWet5IjyU8zbZhenKgM+ozaCSe/+f1v+mADniJyxfXZYDJ6aPHi5aoh
GBx0ne8iFHf2X2a6hgKsBaoxiIQrx2yw3hLZpOt+3FMBubRm7+M0Gsn7UF2faeBk
/H1iXYjWRgAIFG05rfjD+lSNbckhahd+qQrpXtVMLdWcfvnay26ZWtpNNsUwWyuz
3GYKSRvkQFdWE5S/WBSFIxOD2kmfTYTDdUGFxxQp1YiPi3GAvJ+zX+XTmAb7ibUp
l6C0Sd8U/xU4qaIppNECQDufjFT5qmdYF+ONDHttv6AxrxKZa2wD6QPbYHZhvelf
rkwBpr5q+B0+scM5kd8XnuT04d0zQl1Ynq5xId2OLC1UW51G8dXopCDZLXlRrLQJ
KaK8nzTqVmZEgOZ3j8QUOcD/TdWPPAICWvhIbQXs4524MET02RD7mDB3v3C3+KUq
09HnOvwjh+0XmzufzaXG5ZO3fe/hxa6hTpCHxFp4ROy91vhn3G4ETf9DCn6b/gdY
22zmVnYePaUG3hDjdvD9RHV0/ZQ7pe/pM9FOBY37+3YLprHSbrJQB2rmea1OLOBi
wrn2UX4FU184YNR+Vv1MVfFIBQ/zLzNJxaS5mBu587xF5gOXMgCqr7+D8/n1fboY
pZ9canlBuM4HJnSsGBbuo5LKcmVxKVlFDAijqbNaB1i7i+P64iVImqpKXCQr4IBG
uDfyVGnPh5Snc4IdlZtpRG9hsc+IxX1yygUOeeSp39EM0pJlPHqaG0rUW40O1kR8
swprSNnUDM2TLxfgBKeMg+Vz3CfyToJVNOe4nkVKnZCU+nOIubT0s6ubNBreCk6q
0Td2cDWQyJDohAEEy/2sjm3e3+6Hah5ZFqH9YMKxPBC9fPFvJsinSNz0ktdn5Vdd
sPHns8UALpoW3mITcu+VMUlKO1xeGAyRnKscvYb1gOllyhMwzZw2MD4GBqGLMCMr
Jg4hKouM6/XzH6T57lE8EKn8iH7rxpFP1YTg78crt/y4R7xu5OeyInH8+GiSip2W
6UzhLvgJZ5rzAacdoYErPpq9kR1N4M41qNMG6etmGB82k9pFuVgZMRlpZ/6E0JD9
snQ9k1vp//7cYPbJyhLBSWpKPYi286LSOb8OZq4CKyKpP4utfrJ4Y5kWt4Ze9k4H
4GM1as2WJ1cRA4VRWqbPct6ETlhSkDDRlB3Sq7Rwt/FMV6eKnzSjksKs5nVmgDWT
P1iiwkAWmsft9/tf1doblAU/7egDNX0tqDjSDNQ9u79sZDMw6eFhZS+Z3UTPXP4o
wvwWs2VKAjglPVUn611XAylo7oTekFcd4hACQxJ6239BmgNP+Z1KTMlhWOov1qJU
X/NvsONMhiOCEiT0Vb50VnLDFKHwWpwUWKEPjT+7eW9WrqqutK2IK4d/Sy+YbY0x
8lJwlOTUqCq3JW1GIgh1QFkoS1XQC2HmUiMdwjyhs2gUXv36pimKhYYHIMxnHPbd
f3Qf/GE+77SxeSJLuRTvtAimLV2v+RdaN+8cdgiAvpCKo1FaDNC1v8frIUjjFUKU
zaSYp7CHqbodewrDX4HHuUUs9dUUFC44E82+tlWIjkaNBp5fxmh64FofAIUDX4wC
NH04P7wT2CZ+teJscUkxEIrASjvsj4urhlweXGDUxeGxHRwlw/mLO5FrjrRtaIWP
h6sPBPcutvHztTY3cSIZqlA+ct2E7YsPhSo0jh+t6e8+KgnYzSeOW3JEzFDPIOS5
b99zoXQ0s4H36XSwB5JUAjIim236+6108Xoy3vu1t0r3SCbIzI21kXjlAHNJctqF
NqBroJs4nLcLuojNjKxniPHxOssey6RLe3d25qIZWi4TGfUt4VbZvrgI1YJ11SW0
sarUT3/PdEjH9nWx4cfR5ajOv5zaXn3dnz0cLbbxXA/WC5Uj+XhlgAPIaU3M35GI
0/otn2nB7swVcnddM7N3riKnkj4IQlJGD1fTB383EkSR0gjM+IUQdYvP+mXgsUmm
25WQFY3WRK5SC1HsPL62TxAIO+APtduu6kAfE21BdpJm8+AwNh8yedqqWu0auOL4
BmOKQ995DiHJQifmL7c40porv2+mq4RGAIi2uSEZ+GjIu6FGydmkh/oFu29X421N
8AVIgGSzhCEJRmxWF2bu2w==
`pragma protect end_protected
