// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tWVL6jWRb1GE/21DB1Z+jgRNpwdgE+9tfgNjNM/zaXJJGjI240goZKcQxaQabeWK
jtDi0AHbxPJ7fJr3Wk1+6KnSfd0cxwUmpjys3Ikbw9xuIiN9n4q/lYYSKjD4cJsB
iHbHXtIL0C1fBAvcsF+OhbsI3IswumnXjjVaZfxnDx4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31968)
ytS1ELpyFaWNxqF0bECetxo8aqGle4Nx/bxUmK2XYIZYJXcO5Hvc9M15K8389S7N
cBMVe4vdZWsS/XFA4wWWEdB+jKDwsaUH017tjqJtgN21le8ceyGsyal33YIeOh1p
tCxqXCahHjLl4zro9ZUKvPV12Zmfoq3aZ8p8DslQNiX0UNTqgU/sCin6U4iBqC2M
8/NYU7KHH94fYw87QgOaKDuQlTDLacjUN1cdQQPu62XnAC21l03ODqjFCBWbP2jJ
nzw4N8h6Q8PGCL9SRQD+fx/QOwHuFy1gaAkmqTcE25nO7H6b3xCjzBBX35zk+WW1
DTrKBMHaSidhZS37yWH175/rKGoyJqgcSb87lJvbV4qS2G1l6cBwkH5LmS7OXF6M
NTGAEpE1a/rSvMJGhKjrOsnz0qdn5lreBQE1MjRO01Vm5hG0YWEtMTD7aj5Z/Mxg
4b+hVFpmPNDb0eRAfJVVSWM47/TWtr3smYUYdLSn5bWhJWMgkcqoxOoZmQn4Xd/e
q+7Nae0KnUWcioE+KByuNbMzk0AQCHJq8D8XycVfMTep15Sf8K6vgiZO1TevriYb
PpP/OdcrpnuIfJUjT+z16Atphz+tIm0s4KS6N70vCBZvgi0ssf9N8I7/AfugElFr
hlQjmCE0pKMAQ1Gqky6f6Tmp1eW86Xyy5SerC+aXVTTa+HEBC7lwHXhVb9jA1i5q
JJC+rTIGXuwofzK6u9HLnqAiLi1mhuBYxE5w1xGl3nOgNktturEg/1LTX+DP99Al
GNUfq6kgbBlglv6myLtUceEpRXIXjATh9xQF8jcmb2Pe+tPefgwkRvGBzdjM6xeN
yTJy+/Cw+F2hZnpMMoejaeu8uVw84rKJKn13nsPV/R4hWfPqEe38xKfs8nDWuKHI
HmCFwff9O13lYdwEziYWBmcJkT275p0hofTnb9bL/a98gqp+oYanDitHm4OSAf7i
fEio1oDdnbvDl6SqIvreTQK3GaEBthlQc7C+wGuOIMT6i/bI3+bvfpx3LslMcaI0
y8y5u7vkvdwv33dI3sSKd2dN0n1+QpTHJiT6TXAcU+4ZnpRqKIObd2vUExpw3pOj
IM0ZEh6iN0OWQpnY5AQ+z7mx3WhiXKNuebj4tkd2MFO+LUA63YubvybNX5wvIFe4
zkW+aslAGdEagEUfUqZtNH+e/SSeNpdt+oEo+VRXfhKNdlTU+GK2njLVds0FtfdZ
EsdQMJb5VC8wRd+2AHzqrcoPqLeclZg+AKTjjoh3ZHuSW/pO63QJcAJnOOXWsJH2
ez0//zHPn1Xg/bzdiPWav0mScC725xJVOPt0uFurH2nUjrj7tF4cQtJOUNHtLM5s
qwfSYrWAbXBoFNkiQ7/jG3cXdtFt5tU0LN9e+NI5oxG96VHeFPlwppHAtBxNFfPE
AU/5weWT/IISm8k+istCwY9VzjIJxF/lNWjNTdIOiBv3Sm5MJzr9PaKOOpuQOwWd
ZDFO4GbfBLwQ8Y/zSuEKyfOpj7n1s3iOIVqKgSoDqCAljzIO1v7xF9VgO9HBpPTX
74dx3hcmRIklXmWFw+zWvOt29czkTJOJCGjK9yDX0iwVM5EZ7LUrBejRLVlfxyRN
ZkvL34p3bnjjOgC97MS9XV6HycRp+nWohEMIS28CyU0m4IFuf0B1mlHmdHs3R5lf
XdgEirGIQHtc3gGOVdKYSReNLlMRMNb2/DV9Ma/TL+5uVbfOO9uAzw71kRD4k8MK
MoQidwbhjP8bFLmu5dRDJ6hxtlYKckE22OPn9kZVrZNPr3YsbtnNhGUK/sU61v2X
aQzcrmXvSl7o9GlNKHUpG6ZmFUEd3SUt/m7/4B4V+kH7cXSzERedFmcTWxTFmaX2
2YQHOCnUCDBzHtDP405gCOW4IRCxu0GT6FtMm1H1+h3YJjC8Gb34N5bcQQD5giZd
3XjPfV7PT+zmHAWaK29XPs+NuZhv3fsgQBUOamWh7kJC/jNXod4WFF7KT5XrxNws
unihE2qUBFd1J3J6EiCJllM6qEZ2N2zAKi0nkIji6FBqkV67eK8VDsFnc+ALkGPd
3WmifqZKyrU9Sy1r9BiR6XaUjVbe4kpeAKst/NdYRDm0B+RYtN4JEkrU83u6LRKN
U3Issj8veh+naFtINdrESjlbNFxUGKMCxW12fkcYEqUZFmXAPZHTPj/ngrTVdYRd
tPhDwJr8UQX2RibzpvZuMKRBPp+AhgvL45JXfRl4yjh8pEck2fkcrxZJr4KkFqt0
CKhIPkc1ebBBhRltrsmk/MQbxOB5zzjhKDGuO8s7J9qRmsMkHkEzYGbHuBC8+O3s
4k7G1OkKZrqGDACpy9F1FqDAqxasMuRUihTwdAqRZLaBzLCPLqvn4va+iWek0iID
ap/n7/Qeqml31+SClr1B6myEzu89ifb8rnclnkQ1isGlh+PhHkgctALssLyu2J/Z
6P7TuTB55uJQL5vF1n9ewhvrpVpkw5me81p5BcrgBNuDSMPbhJ10QF6kvBucETFH
BWTAHV1rsFNtZHyhbCEobAnn/xGbPbivnztMGV0pdfg8imAXE4aEEw1FF+P+0pab
eqtPiL5/O2iRCb4TrRzDEa7VsO7thpqKxeyYpVY2aimc52dOOPWVX2df4w3g7irr
DpSvmV3TgeWjTb5Au9r1jKosZSfO6AC9QOj18oxLnN4TrwXBuYvwD6y5PcJX9XEL
q9pCdsfQgh8ySa66eszopCiIMquxsRiolGaLv+NgSBqvoOKhZzpaZ3k/pfQ49l+q
aR+MPc6mcibzQ4WDKyWNKIyYSG0mHRS7Rm5tklFlh2oJNx0r0EX3iubi0GfuSkQD
I5/dazisHkJYjIkCPraQJEqIeagXPNPALmXeR8p/WRgvExmjGHzUz3ZMCZOi7Fg7
HgezkmLLB43DtnhXJXNFLTERf1sq/dPNdY6Lxb0Z3Tn94YSPea39u9iivTkrFKBc
lv/ABDLjxl4HGkbKGBRw/WKZ2TyLAOSSoYG/Dr8rBG3qyzdduIzYoCOV8jHzodkv
85efOKCam6d/dO+8Z27+Cz+/gMlSCI+I9RuaJBPI+TgQ3fl97jIfosurwHuUG/1a
C6v7hxkcFOlun6NPTK7fkq3Y0c2X6G4mXURlhtRqivUEzSut40PkqAEmCYG5l1Vf
GWS+CnnFNhoqM+GFZcrYgKB4b1dBnMZDi2YS4nAqDy6NCOt6jUdOjRSnfh4kG2YI
bvCFTFEVRKIoZSl4uGJwuprFsuIOoNvIYgVgF23MFK7G9KZvmH6w+LWGbWzaFdiJ
kUyRsDZCTlgOxLZ3tPVXnW0Fve4dUuL8QzVtmrDGV6rCmSyJxuAf/Y/1CkJaHh47
WTlw4qn/cRMwomnNtDVpwTtW/HOOqIakowi2z3ig9Ryo3mZOl+ihT/HXbOSIeuMU
/SudHgJzyM3w+D5/K9bD8YJOODZxbKl+NOpAFy0dTGjOH6hTLG3HgNjDWQsr8GrF
SPQAlK9Oq5+Pr6ZdFeNOIYiLkWCMmtuY3v0A3UHX8ksFxptS6HPjC9O2ZY83FZAa
rlU7RTomUSg6bihRSwhSAWGE/yiiSADRSEgw82bUa0Fc2s9CkJQWYYfJ7GcdUSGA
hn+4fnwRFw3WO5/R7GBhJAo1mYcJOmIV2cXNnC/Z/0UcXRgl1hN6IwQNs6yPIkOW
bXSdQ0QiDfejptAD1uKf9VdjKO/u+VSUIw1C9hEJYpjfczCUqzMqVXIlmO8wOQbT
ioq6ytlmKDj3z2t0ZQ49i4d0If3M0tNb4hRkfsh7BcFiDmF4TLlGgzXzH/A6r7G6
ukyU9NxeB/angzJCeGB36oal5QGaorT2S9u26YdfoJ/VCcw0NOnYCfwL5bzKd0k7
3V5fISFLF8rkT0kLR+JCmKVgD0F2BufeYcJL8IaQu9uiiHbPgMUWsqSepIxHDGig
ERvFRHAdkXOUId4Mbn8w/wpzLEtTFBiyzbVlJUmjIFbxTgHdc8XFCkxIjO6Rjqrp
EVCxjm7mI7jlxYemIkMklgfYqlxgRgyGJ2nkszJsX6xkU/CWCY/YiXkJBT4RyHTd
kf2zEtCb66Kd72JIqHUPgMpMGWXN0PSWhKLEw/HWIkNtaunuj+Mh2jCpgcHmy3sb
fkCkprmoVZ6pNStVaNVKDRAqnXjrB4UKyLmuFwikXcsxscL/piGoykngSSMSO0Ev
PF1DiWmttJywqC4co5M7pZxr/YIVWElqmKqGWJT1ulzcYhN/qjXCkEeBhKV5WAjj
yCp76bOBH5SwigOauuhM0nhwe3R7/rp/OzYtobKsdjpWT02LDi/34nZ/A2d8Zuuu
SW8IO7iT9F2/bKdRqfZUWMJyRgB/nLJb7l3UfnE4MKPz8YtTmi2MAKQI3I0+NKHA
i4Z+1wSopDOR12cEToHMGva0Y77YuK5PysVPgpFjtjW2P4PuFVDPsaAFTzdyc/Y8
WIS8Jych9mgMV/bRZM8qnwBaolT0o/YLWhwHTwMj3wnHn1DxFyds7D6Zuf5JaIX+
osTBp1NxIbAHWIiyZpC8CuQ9XQFGIkGCo8SOC1a8VQ3ofnPR5PLTnlN0IipL+VGy
wGT1LhWPK2zFxWV4YKjOJnNkKNLLLQQlcfFKXFk3Ak1DPdK+y9VIfdaI/+TFUapb
Xs5mUH7p5hdLU/jmKuVDF3vLCS41t9UzBt5OcHCez+f44ZJm+bUYoscfRUUFe/ns
wQh0aYdvMUljtmbCqJD1P3ex4V7eCFV1XZlpF2SY5/evA/HXelPftNHfAbOST2lg
+XsT2IE0s7otxKMxz3kTTtRPVE7qROB6uL4w+uVm3DQJIVPpkLMly/5Ds6JrToWI
IOAsU5Zx+xAu97rNnswkzpu4vaL/tVMO6LPC0MM8E5AesEzqk5Vpriw3uDei2e2S
0psL27IL+T0lj6F2FPOG4vHst1TIGN9XWFION86PrJqopN69aqkVl/OhgtUjA48t
iaRS8vzAMEggIL04Si+28QScPzXqlWD/pl2Jm7fJel9wYyM7qBP5uxVkExNfgl2B
AQU2uLbLqMf9yFtrnHAJmvSzPA6xCCf6PMVstWR8r7luXBfb45gZqho4cU2TP3Cs
Shr/kgT1mREYFup9pJBvmRoFPHRTfub8wr3kx/FlGOlN4uJvfRIHsMSFDHppq59i
icT7gnLuhTvrqxhUhyvhfGqfr9ocGAya4lvqXOIRsiXANngCTMXB5Dp4N2SioQn2
G1qUcmODPzXWSdehOQaHU4yid1zr2dVFugwmVnKks31cMjUe2/SoBeEZbbem222A
g2JJQkDNbQFqMb3rzpHh8G1MR3MUivdc/AKdkUpo+0mWJ3XpVv5uxHaftW8zJyGZ
TUcv/giD1AmH3nLeiFPi0FfIfIiNdPWm/Rb+ybeqiOcm6ApZL+PotrXUoUH8h2PB
5IHx/2j5v61L4QcelFgd2rql1NNjKZunPYaUu1w3Nlo2ho24AdxufqkdARY14Yr5
F6GPBzCHawbhmgR7j9wRCKzctJh8VO9dGhca4tZYU4cmIjLlY4qNrpiMMbnbn+cX
k2Uoxf8m6qU/3T0nins+oh57dwp4iS4bdTNscQxIO2oHC8TBtjGhg6BWQyS7qnav
QHt7+CdcDZZ6poON7Zku3KCk8Y0wdrs227bTpvT+S+YXvh8YnGv/iuu6zXjqBMaj
+B09T/BiQgC14fAZXlr4ol3ypAjGWHceM/rSXGFBfMJ8wTYR8z153UAZ2Y88DOKQ
28IKh35JlymBOEmcMOHrz3eHEsVgG67uKzCRjL9Cy8q1Ul0pEFGJY13LXVIT6kuL
0aE5949vrpUm7fspSiTGJplX1I1gsJMWugMrdSU5Hxv/Px4aXuvzUwf871GgGKzA
9LeJT/uqru0C74guyEzIAZBiVezbGTRAiCh0E0hPDLfJgZIXmLJDfAgmNUWCDa96
8yMoPH4DWUiwWRkNVwQO6vhlZKSPPO1g8SlU3pHistFHANq65r3u3/5CQne90PCU
gKOnAIULWRqExq92e4DIf91lB/ouz9kBsInsPNTitzf/ePeHTc3EuxVYkKMzttQ8
rl1GC7dvtj9gHFC2gqFRMrrNHT4GiNp7TPNA6M8Try6YjA/YMzUwJ9pvaf/UtaxJ
ToUa1Up8wntzROZmz/iCi9v1lOsi9K8xOaPh1lKULypMEAw4alsgK8FxrYUfVH4s
YoI0SNs1Je2Jhymmb/0zdyTObpC+zPyvhjjwrQOPGP4gn2VJiFW3veF9I7trA7t9
Q/Arp0ZTUR1UhUGOekFlAISXKUIy/p4j8pQ+FMZA4ekcWYoUEoOJKPdsNxqSV719
vP2Cj99lDYdxrSKkt/oTcmGJgSlEhf/pb/D6jRKPThfTWvrQXJeP/v3i1sL279eq
IA1czx/nx2VaypzpNiOaTUtBV0ZjpMyMBlFL0iLRl/BYCbz8l5Zk1aMI9KR0rW8M
HnH1JOLp1uXKQnfPIMGpqk049JpI3slgNbVOPaekuEZDqU06trYM/k4G/Ri775ED
fhV2I+ILiwNJ1MX9+d/nYRPbKRkNYd8Z6bDR/TWE1a6ywcWfZpIcqcnxmUh6VwqQ
o26yVNi0/rPRz7IQmHoAOXUUW/8jP5Y3BlpSUfbn/dX975RlKlj9Fw1nUTvsgIqv
2MmLRxdtR8cypUzzC20fJsL4EJSMimBQO/f+Em8aloZUQ4xAtcQTtkvZGa2XTGEB
s6lL6Q2n/KfEAbEXv/pcIZnIMu6q3OPecSUMivNQq3yRqTclNQWsXH6hxMTZu54E
+0QK0RzhLUSLVXE0D3HWt+hN6u7lKzJI5ECiVDBZq2ob09Ci4j/5uh5Gm3ZMt/aR
oLFLmU9XgAVzfyK9GSfb0qURUB0XH4nYFLbL2kVnvpQY+4gixfF29ou04APWgiB3
yzjOgjfEZI88CuUIXHTFNgmcC872DW38fK3tE4XsB9SVkcyfjQcJK939AsPIAP+w
k8pIFRyxpyvS/EiLaWtbpb7SX7Z2lJUx0lIpVURD5hQngdJB61pHeluIBcnWALR3
5IlEPlSjgDH6UkaM/03IJJjOIy/zIaLmwHz6IWBdEuc4NNZr+pTm1x8dQrkB/rrv
qleKk0P/aPYKXmn+qZplKKJ40YX5UjNq4e46Uiotv6BxybD47mN4p+26TXHtFbj5
E/7tJAhgfe4YtuW/Ax737UDvfBo/xW7l+uW5MKJQNHcW2Ut1NXNtfp5RCBpFAlhz
XYsMXGtyd66XhVaKmdOIhZss5uSSxUNjQveUgUtIcypdumhvC0uoYCTHIeDejany
y2Z9cUFUhg3Y0ifrG0rXErDWmVpjb58AHC6GN3eNoxNEZhoUjtuZMJXp7KF/tTlJ
0tSzDFeZGWASc3HLrycSdmCfqQ+r1cdMNQP69QZeW8EDQ2l6P3+L5/AUAMZOcBTd
IpfyILzU/LJxZeEmo2JOpShNVEjdnsrymbZCbLXP96rJGKNacMj5AUFTmVoikm4Y
950zndUMmMITSyZMSJZtNJNsahgFDYXdB1wl0UWcKYu6dopkoaouXEoyHxc6244H
P0YLWuZwakOm3Po12S33eBQDwYtt16gFvkhxxMYc+6klnYrwKrdcYY60WS6S2CJI
WQBlZaj7iBccOkNWK0MTsBPhzaMf0C+P/XTiSMNBBhyeCpktGwM2xmxZooK8DvBX
Y4axv93pO2/Ol8AcOo7I1SWTDpBfRAsxZosxBd/p7K9d3esB6gT3zdCen9iREOoM
WsLLJAWtq8h1LRZm6ucx5MEyAS2+MHVLVwEBtLDxMKcZlOSDhia5xmxfCPeikigz
vfAddMT90t1NMjIDHhxu6i5WdMN15pSvbeW4x7AfCDzZxLiU3J1bmNnZsc9C/yb9
TUfTyjMABJQnv064IBvbVzknXjvD5qVrby9Wsriw6SQ/0F3Nb3O747IhCZAlljRo
Lua5U0FXqv3FYgn29TOE72GUIHI3QseKnSp1+totZ27Cf5wE8vp41oLPuq83XSmM
WiJQTNNx3M2ZyB3g3DFuVM3HWkfpIvK9FDC9NmQeNpJ8+isWSBOJMtDOBRv7IhPq
F2bejT77Wa8dUkh3fKlrN/hLuILLQ08SZZ5bIqxTa9zsrxhes6pLDoI4F06GOCI6
qmOyghVGSkOZ+84AwIykw/z7MRcODDi9BjDt+utKBRZRdTkML18boLxhS1UZ4g5g
XTsI2J/VC+8ekVem9FESuEGGNVmjpOtqyLK/o89uyKJ7WLf6eUnEE+Db1bNmbO8w
jkjVUmwhdFTmYJiQU2e2h3z+YNcX/02V5BzZ/QmfyVO/LwnAvwStTuugcupSCTLm
kS7gJdIddNhjXsz2DRbFhEXCsNaFsJrj+QKD9cpSSquBskF/dzXeCUEnBWf8Oypu
VWqtlt78JQBwKkQSVDHu8kWTeGNmt9mHrhJapagB0PeWhvV57LGwquJIe5sLy5ht
cav25S/izUuoOspYGNgz8O/XBkd6S++Eq8EHeE0XhJj/dhSASfRdB68bkCLZ96MN
yMf1MEAW/QpsavVLLAFa5m09DB1hr/QRq40p1PrhMoCK5RvbirHtyWqLQG7xlg4z
dzUBja0PegzAODHLKJwE8tMKVB9qJMUhSWDOvKwRG0RcFRmeY6rMAofq/X0NBGfE
yCzYvTESZjUTeno0BSRWybpAYzXlzUgxfS0S30lKtDjdscr9s26XxfVP940jvXax
+yUNfmbyJgvPEnzIisCaNu7SxQSf6ts68g3zeCZfOhaczRqRHwErnSIetYEkIQk6
SJwxR4HEG6RoFsU1yBD9h12aWabM09OCzBQzaObu6T62+Hi4QS3B9Yt95DTUsOaN
BGo3o/93gQsDYCagAuNokbB4l+5t7exHYzvAVyvsvdoROPOT9RQ3z6VyzowGaFgt
lotGBR2rI3XnnavTP0kB8ZpA8Kpb8H7whjmdPiWQZuCKZJp8RcVA5gkWxnJ1Yg7l
WsiCYBMjLPDI3Ink0h6x09jZsyxfQhpBsGE1S+Ez+3n0nTg4yczge4xyGy6cJyh3
rdCBkn8ZscYKsFA369fkssyyz1xS+r/AtDHMqxZLDU6OAl3t5yCyMQTU/jH2JeKV
PYuyyGNloiuIJ9Qz6D2so0g4dFAM0P7yVMDsI5nbPkpSkB8lFkuHeMe+BZ/4qLMq
YJTwLEVrmKaZ32rtS1SwafclyeCOOw+FH6dgge+3YPqFvi45if3ZMv5glztMjU1W
ya3Bvya9qbpLRzNd/cvHLe0fC6pC68KC1W+eG6rsWjGySRErirt7he8j+IxqVBPo
2jM0miMz6oAs2jmo2s2CuQ93pUTZJ0OITM4FUVhikbTGN/Qq0TprvhZZD84xus35
PAPt88ozjT3/7fLLEOYD8l72Am086gwVlccWnXMi4QLdxdCsTtD77jyYP232gx7i
Ob84WY12hf5hQBulnZALg1qn+TmEuxPyzTtr54egiHoWUN2nSto6Kmze3Xrnw/1Q
ok5DCPauXbrL7/KZLrlbfW/7xNPKbPvgj9pZ7dTWeM5tDQmUjRt8aXOoMbjmwqnm
JEgCCffuMyDpuJ61VPbtU52plg1do1tchVEQS/XlVYJymyWOXokoEQcKdZZnEInS
UxsH5PUi39brTqnKgIdFfpUWqDXp7nS5d5gu7Mwbwlm+JmQ5JxyKDw62zK+zym8H
NbKnQpCR+j++fg7ykbi0/orjNc7HB7V7VE1mx7KHmWez8U6EAOk+Mdvz1gznZm79
K4CPY14vrF2pqx9LJMZv5DStPCJfChlylYZCqnzVBkfo+YAi4j9aX28JQuxaSvj/
/E/QsCgzIMS40OHrWwfRRA7WeMDnxtCLZxI86KvmvLkWaVk2CIXhEtVO1r/0Im2W
LdlUgjMfDvadpY+ZwU2WOj8b6TKfJn89CQhkQXVVNhyCeKEafU24nHpB0pvlcXU3
wy+xv4lcDwuFU5kNAWC65mny02ZE0/Cqn/3GUE+ctYNaprJBfNsVgCQWcZkRjNEH
6xGU3cDdd8yfRgTtmQxQTe6O0gQ6bJL7rBvvEMK+wPNQKS+nhhj2r9skL/Qmvian
JKMtiEVnRBlliXL8AbAYkH/V882vVN3kyZ5nEYxJLkVRhA2dxGkXVSlxAj/7lBJM
pyAFqlm9mhAVdMsyWfhe5NLLjjEocQJCD+hI82ii7DsySHjpOEzspwzyUvzRdGbB
7bk/10VA9GibnUXlWFxe5itxhaHqeo3aBkGEPeyRovLth31nJEyRiD0mFCBffjx8
LsCw1clgYPWS7DqAskmM3aY6cYVZUja85zF7lmsrnSiQPODxw6dCOIyoVYuGsqWW
v6FI/UIt1kxgABzkdXZpRYhqEdZHsE+9laRYvjyJhPnqP5v5vJosHJUlvPfACzxf
nPdZCSRKn1eWBnStmyffSq+cYGmxgYXX8LHgImaZftvZih2FEypbxW1sgyBdebUi
9POqF2IQaxqHFLiHHlVUYam+t7nu03WmAKiqqjybGgslFuCLLw2cg48GFbIAripv
F+2BQbnOs5KyNnirqw42LLPOg68x/SEmEXFYD9PavaT7KnaadJcwOowA6WBpcelM
uPgwthhR+0YshEzXX0Z5sm1F328gRgapisUwzlWYqDVg36Sby0OFwp0Kk5L+BerG
wnXjxOS+kggT0Ayf2fSLYgW9G20Xd+DuADEUIz7CZHOsp1f/2VuzThQo/+iFqLJU
VhBht2igPTypNIVAOb1sTUJ5x4fTUcp26cs8X+sZkiDrYU38B8cKMtmq0/TJxMya
g88Y8zmltJHCHfgX6DEC6H+s3EOubA1ZNBayQjZep8gZGOYarBJI7tqhW4Sg5jEe
4dnYIoq4Uvtv2Ck0b9pUWIMNCnLoDkbAPTDMv2LEaT7Hz354OosPP9yy41dmwRtJ
+EDZKEXBmKNZ6tRzWfPEyF532TKYJQiMTJJ3QrS8afXfGqxN9xG8CX4KbL3xvciw
AORuTqg7ZC9rAa0n9tDazPcCCvLXe56aW3UIP+sImj40Qfkxh/1+k0KoThMGT9mH
kOWndDjTYFQNqMzRj/foCSaRXfsXnVKo0M4EY3eepqRA+UlkLxSRNAuvSj31fHPW
Oyc2kuxK2WtQ6IkeN7vWXm2eEYxsPPY0N1RueXEiKE01utWrgP8Sg1TeLdOxprrJ
Z4hHXdvKmYMf7bTRWzOCVp4BOF3a/Xm7EaOR89PfMD+IO8Kv0/R0RrKPW/zQG1yu
LajfwBQkKiAnPNbFGBYov/YxNjsazYfmBxC1axXoANwWIOTrSibyaz9EafbfvPB4
O6OYQGDwUR2XNkxUz+KfYzBHqeh0tWOwHrj1r7LXXl1NMQml4sLhRqVkWWjO4Fk0
ZvuvMVYKmbKWhPuLDFhuZs4J/EcRZyo4YtekeqQ7/TkO6dIiNozIPGkcdJPCnV3J
AbKKVkBXQaAYxiCT/ybwRupa4chARf6CjrFJvUqcLbL0vdy2HaUpf2H1gc36xMf8
yLZnUJ3NwX5yFGk7jDFY7dwIl06Y2qNki4HgQKRYfQSf9PxNlkXcAT19W1a3987/
6lf/+I7Q2tWdBhUXip8G5gYXZNC+S7NYixF91LnxmLyXck+1lEow3FPm5IFCBDco
0tzvrWbdv1b5KHLpFR4ZGY10a6P9ocCgJ/xWq4RX7/gPh9R0zKE3sXtjaNPkF/3l
pGtYeDI2gGOv1+zTKBUxgOfxAp5gVD78XRaxQWq4+XcHN01GCSJalhTLnZK7pGw9
UAQnlt43mD3anC6ika2NvhKlTC7p5Hr4Onf0vQeiujwcLUuRIYkwpT2u9wzXtkGg
pCh35/2hvWMSrwn3069oAYi35W4weqC4JSFq4eV1nxdw8zaVk8PC579u31nZ8Q93
LExNhWvvzZ6vcbQpIpc2W058O8+x+NCIPKS3xNTIgcXs0Gm3m2cAIti1lnzRuyYg
dav2L0/UjP3/88DQUwvZc+BlqaF2ixTGUO8zmeBOSf7XrFXkX1IZKHVlU+STssgY
b2ehpCebeFjWppIii9zOC1Hco6my2UwJbt74xPMXqLe/dHIXiTE6+IGyGcRNV5vv
r0ou9nneB1Wm6Muo3auxTaWcVKs0MKYwjRPF1WkM08Kgb6EleJknWTY6Y95k4F0v
nDOsjtleE6gV/PrtcMJkpTOntJyxMM6AUXbRLBfHMdOsk3Msv0furxP0J8sfAGoS
OLhFVadoB4BVDD4F5a9DSP+3KBk5BVPraLGjsW2eq7vTTNTdT/jU/LFW4xpXPiZh
GEG2D8rihpcyaUNOHeTFIgIqGYl4fJffIne7MV2sEMn0lQ0fHdj1Ywhkftffj751
guvJhMWjfWOKeGsz35VvLVMAO38jxR0JmaxFEJhXXpqIgIggV+3I5S5Yv4AIa/yb
/pPOG0ZZC6L8T9rBJj5R5hRto+mCb1evebmo2fVduyj/QDAyZ0o1stC3rUhCIknQ
O5Zjp40a4rATLaVvBhPpGDiL1goUn1Knd2Oh1JrQB1MsYa89nhB56Px6UG6KWwQc
8qnzbk07EwH2MBxkOYVlvub6aFljvBTlBPZ9p6+hK28YTz+bqmstguUQ9Qp2xStw
Bbc0bNxbkvp8YzE8BxQYWGCTvAisQ9ckC93hrzkYVzaw0f7XUQyUqgsrIa1BYscq
1X/bBaDfKwWECWs67zCT90IBQv7IbF/Kv4a4ZQDrzujEojq5499mPEl0/PmA+1xp
CnlMh8LpTbZar0FDTJ+HlRxpKs5z+iSNFEEFP7Ua0Y47sAQKuvQ9M9tvgWNbRG44
gpPcPyJutKGdpEMgTr+XPxMpwq+npffcIQle/osWFsg38RAmJZBXv7o9kKKcfjE1
0VY8jr7o1nsjUOsxwsC1XeoEaudj2cS1UgWycAGVJgvaPtwt6ap8Q5gzPND+uAcw
UCDBhId2T9j4oq7t0Nlqz0qDrg8b6eTXxkKzeSbOfNzS0ZwntmwBOF2PQ09sxS3d
RNMjBhunJ7zJKvWQcTjjngUF+wjedS2169r615Ic0GlewlTSm1A+hhUIVKBw2WUF
3ttfxpoQKbCqfELb5RhqhkpwgE6zIFNlJ175rqEm3m/vnevp8SHT8CxzkoCMQVGd
qfnX88DE0C5/jxqp6Yo0XCGqg3ppigqm5wQ1Kp7OXYmV8uXnpDoXlr748deYmDgy
LNcUsbRpX1BnK3ry+xTbM7MqfB7TzbM1V7VVmhI1x4/qU097/H41FzWFMTe2LGqX
c14Yzs8Y+SXw4z4Toal1jOEUXmYhOY0179Y9Wrfzn4LjyTgWTCDlPRjelA5Dg0/7
ZCYqKTRkA5ANKh0QsTjHN3mJb1bOQlvCVUcY6+TIlWH4GYqSr7kofXPgeyKI32jO
BeJ93OzQd4gD7eSBpJvKWWtPn4qNsRf0TW8F6ISN7c7PTAQfzVYgejEFYZFkqn0v
8yDNnqV/IrCkGOTpPIwJZWsKy3eJQkSykeOvju59qWelVUeyNVN8OPGrG115JIN7
58WtvOftlvBM5m/Ie5/NJOqMMdVX1fYWqZUPYsX5fiID6/6keYj49oQz+7pNOBBP
852nvrXcnP5uLMA6MQNHIiuPTRR9Mc87bpjDbYdxXy8WRf+IGyAZpN7eAUrc0cRi
+n/yNIHNedhsm0EuYMQF9K7hV02deUKStEEFh8VCL7LsKSv7++VlEykkTbzHW6jp
kUsPZFKVQ9aSeP5/9v9pa8UU1aiMgUVGJbpDLZCEBeFdHJxygfRGYsuHtjbBY1Z4
ZDDVYD3dEgcshutWAYNqJXqJRI4hUYqsXn+PuYBZLlIBrt8ClK68UAyJvpBVVyuN
McWK8ZUuW8p0IDFRkvltboVKUSNc/rJy+KXjiweYREzX0lnFGh+x/uI+7oTsKaes
OaSJoXa26FCs3RW3DeeuBus8X057U2yGkM+btUhJPHTnMzy8GOVKILj7kQALfD1E
2BXog9C3ePhpkMCI6ugrmlc4/SEeppLFNWd6aAAj4ZUabfyhcidLLUJFyugqJBsE
4i3PPTwN//cvtmjNEVPHTIpvDmQSoUf11DbgONMqaIDjtSQaRjVlLhc8tIjvN6Ee
X41VfuQYn+zHAftK5DVxYHnGC7cYIwoXwhIuS9nm9TxrzQ2X1WVWGDDlarK4SJZ2
t+0QoOXKw3QZ0t9GBGd7cV6wlSsjEQyUlKDQcmbBBB+dt/5Cc13RwFuAJREBX8mu
N8FHwwlMJDCcvLLAFOzdHjz7j/UnBUqDj+FShU24aXjiB3LtuHCyFCnuasf1z/V5
awrR4X0OhZtD2I+ObT9p5ECP2z+b7dy+abXqreTFF6oUpuYB0+jS4FBEptDRuYHi
eWlN4oPKg+iL2StoPpRVbdS2G/UsMuN76HXUu2IVFrPLvxhYXBv3Mi7/qfgH4e3L
ecvci4Trbi0ulbMdWnRNWSS2l4MRZCi+fu3LwIXG12TKJ073zUuzL9WVhXrj0sYE
d+FRoh3IiaTKaYe3c88+MZve1nIFP8c2eT1EbwbJ4qBZYtootYxtS95FegbjKD/a
NQvoeMD7C7VlSWmuhhcOTeY/NoYHj3zUE+9g4nsyZNXM3eU+a7h9hgYX/rPr7WD5
qlT9tRiIEiqj9m8oi0araJntr9eGizKmulTiYOenyHX935stQbbTZtWAoBF5Rqbn
wyyN0XGNEvMUgGTmIqMWwRsVXMFQjCmzoT36PWhArE73bg5FUvkxr5UWHdv8ZLX8
mT12SaSLSuBS7Px8Vlfiwdf3fW5+BBXud/wV+I+QM9U06Qn+8XCW8Lv8tXVBp1yu
sQggqCs0xVW9tcK11PI8GON4lNuA0KcIZfEOO/k2jhN6zDrUWApGq0TMu08kF+w5
dE69eMvWVcGKegw/GIrxDoqql3ta1mMgZnRnTKVjni2lAst2RXDBudVfm6eCThyd
9sz9HuA3IKaIcUziFysG5/0IJCUb+GfqrEhGi/X/dBMCHGSEAR/8B/fmhgG0ThIq
sh8nPSg0Juyaj6EUw4toO9HfxvQ+jM//SYMd+mVvL+AlD5Pyd8buIWAdQmlJykd9
akdQovAU4RcN9UarWGttyg9Ns1zA2dubC5fB8PTyhZAcxo0WYrPkeCaZpKtXoiGu
Lr1AYN24HGNY87pLPaqJqoQfmlAjqOd8RQb6XZaTxmCuwmlPCCU8OT3p8PPBziMs
HR8hNP1fIaNGWMYkqXoLsiRcUzqbMk5JVcvXoml4MeADrxx4icruESEKc0HQdAkw
vyuy47XGBrHBXp9ra/9VVDc903xpdkwmylJkukWaKO56fhDKXfLC6nSLxIUcfgPc
EsUVlMwHhGHS+vpDI7PdzjNHrU5JGgwL96m4e05UqoG10HN6AIJpeD7Jx1lVHvUN
8a299glGKgZ3tUrg8LZlcC4NR5g3iEL3iSdEFIqitvRX2B29+rqQkedWgjxFpegJ
0MAl2W5kcplvUM9OI5LflU7dZooQQyb+VH3FcgKsBIYs4n7pw9mGZTGyY7s4zb0S
KryD1NVsl+Y2FXaWZSjtID8NtqlOiMdh/+WQekLhp7cnFJNLhDWJHWdm4DpaCDRk
Xro/yYSIQeRWNeahiwbDJcLFPHF0WLE79fPAoxCkJN11ozNjgh8flGn5mYB4Mipo
XFgz5CTOQK+HdsX+3nwu8MOiJrZFs2RfL3sa5Nm6TRn5XsoD7093+7iOA+9lHOp/
HhsB3V0WhTfkGEQFWpq2yRUkGEQqXJhNvyKLMofZQ3846mzoy3KIVYvYHl29G+b7
Y1KaKx25R0nWLVkVuYv6aWir7upwVEfDbgPlKNh6ixio6kqPonX+ZHK2VKzSyIo3
U9CqGIgsuio0NGXzZ0ttLoIe/2+svN/nu8Qm8gsqv6bfosWP5Ta/oH5Ni3wZWaH3
wN1OmIcP4jz5gXrCNUxIwhfA0pHhYV2O5A1xBeYBGQrvF4gZzLrKjH8YiPNOLqPy
6NAvTmdO3TACRS6RWRuWQmxw+0ckdO6XRLquRH5DRJKKEqX57cH6PhsYt3Tbt72v
L9hObpKLTkF2tSWIQNpUufq04AwiLPlmt5onWRmktf8VlmWcNxOm0s4efAsquloY
Wf8+0x3ttqJFX558spzrIi8Zw8EZlO5m0/YXqnXnnNQGu4B5LAEX080xy43LxS8G
iVyH5s+Fq1tC1xtXx2cjdz5fD4QWfZEwkTGThjceEbGsdqWy0ERk7tTKvuSWos/8
QqVHrygv9B6dtrUGjQB5DAzANQqbt+1+gUz0DURmKWXvEENAdc4eAPclkL6tThc9
kcVWXAPv2mfNmHRc3MBcXUsAepugMGXzLn+Sv3Fag+sS0vgSmYnKNtRrEAEkMHc8
B8/7VhbmOl4lU3ALTLjAOveJQCJZEXU0+TKoRdx8HrabvVDPaaIaWZCJO0ei7kB5
n6QOqjv46j+nqK6q12dBy+Md+h/J3ooBcQ7oV+8sPkOgH5tHexxqtrjo7io8r6s9
1OScyyzMwQ7QY2ryp2RkufXNk7ufTOGGwRism5Adui85epJ0Oj4lO9mk+ynX0ogo
ZQBXIHvIsWnI7IiNc7HwR8pWRdqqexksGkc3r19eqcTTMB2E83WhTdWbYv6NICI/
mWJzAciz4S2qEHPCmeAWJfyIHaT4qBMSN6WVip03/CrUZ/z9drRsG5h3oiMaGXA9
zpPh6q7KIGbcIqQ93HZEFbI+OdYYmu9pyAxaofLm83qLolU6DhpCqPJVb61eZZsW
/HNpGvwP4IxLrVLLBoTrWNqeM6yONjFpuJZRdnj4TTGcRW4GIZPp4xb94Cc+F1ZD
QanQjkEtfDJEGud4yu2CMsOesHBMmCBCjBWW6RohOy+glJr5aJp0INH1bNO+4sbm
6GKbnVdKHfSQMVO3urvn+C/TMb8gQhxLTE00SXcUXOHaYA/srHmMZ6N4EsFmnVfo
vwGytCOj9vYm9IXU4Z28L4jQqcWAIyNDlFyKi6O0yjDUXUGVR6r9evOtsNYVd3lp
e+2C5X68Sq55v5VArcWWJjPydfl5XQjbS+HdjkVdEv+EljnfIhznffLSz+Coyt/E
p1l4ZdKCsiz+vHigfcYdwe9kubg/qyqbHuuPDcO6d5QxvF5p7lSInTdLqhFsv129
YCM4Da4q3aqXl/yilHWdD2yrTuaLKhegm6/piTs2qrQ2rMXMzk0wPcXjMhm94rVn
/lihoQ6urR9ycC3Z2kVCxs6aFgvjHwLB5NJcCjSUfNwNrXVPEhxxtw+yu85UfQ7g
4xaKLfj8pKujngrX7cYosyLgSWlUbuOj7jW2rZeenld4yWIBFwWijr23/ENzQNU4
nTb3BjDxQxIRagrBzJtGVd3Y9zP0Gyf7wiSPjS065gMpZVFnV3LQqCdfqDiONofC
CHSNWgYL226sUiBYCgU8t/9YWlqZFNzX/474hllSidS43PwGjbbsemF8IH0OS0k0
1aMP5nxSjb8YKjPaj1C7+UI22FVIgsrKV/4fbWlX3g2KmMgVRA7IitK2tyiuAxNr
V/43j51vYuFTfZ/U/FlmKo5rF0/zD0XxsHW9ML6D56JZ+1caFs73LL+NdhmhChuN
/O2JyF5xkFPAJeMK3/TjgEIH5ouj0/Xf+twzeFT9V6D51TCeIjr8VlRtHwxUTVw6
OWZtXR0LjuDutetU0JmXroiY11dCdMF7F40RjWgnSFlX92uziIJR2ELO5i64309W
RihZwee2F2qPI4MajIzTMYfOvSZUElEcI2bURNupWAsaAVskobhJAtyp1xcmzu6j
Ge16Ur9X1bLBC0NQL0johVsoUeZGlua2qMGXBwEEMzzV6vVOFlekOfgP4b4Tchbr
k6MqMtGUW+WtjVYqdTfEtscGR5xOqGuYVwn4vc2J4JqyCl5FZPir1le7UvFftOFc
rMlMaKh/z2k3+5avfbGCLQZe86J2iLPf2m5Vwjc4TRVcK5xzgsqFgYqh10QUhqD3
M6LaQQOQkVlDTxfShhdiEBiHyQ5WCdY3P0pa998Zik9WAax06RKxinbI+PGsjXqu
1QJmEIdfkksXN/rA8+ZLsJ3oRKTtyg+PIy3r5oTib2WCfFJyTtotKBAfNdXOfOqW
Xnj6oBvwsgyy66bkbxi5Bdhc3U1apdAZZeb2MvLvD2aQoL9uxqqkQCus3xVAifDf
y0gwD9OtmQ8A8YayU5F6YWIz0L9vpaSHAZnAx4cgxn4wclvgbQp84u2Y2THobP0Q
FxnnHNtRhGcl+232X+Jc7JSv7lzOW6z/SbtTFIxYCT2aPqQkQygpBSau09nKWKra
QMXgj9x438hwDeIyBIeeK9ZJ0A9IcKT31w4HSkNbO6PsWsbz8nA0F4Pc+dt+WGk4
JW3YqnPLKBofWKMcHvSFoIQsnPPI95e3HE6M8uAppza1uVVu1/4fmwhPyXPw0I/e
9A3bz3d3ypmOcmjdV+p/p2OFNNhuJ0WyP90iNEFqwBZrHnaIGHCkN2OSGPJconOP
FykBI2cVtJ2446pkOxzKR+k90XTM6L5yrmGRYoIRZ/iHG9gtAxY6yB6QncopI2BZ
g2gtcJSnIgETqwCnkrdtuz2Oe1xcCVFJHNQwXqdVDF9QDZFTM8ae3ts//kBs+3uw
JYsC2DfG7xUka6ubBMi5fqpG/NV4u7Rft17GpruhVaoT2ydp5SGdxxEFjmvSpyBL
6rYAaC3B/mIqtwX3Fjzp1P5kbUEovvbY05k5OlQBaTVLV1pxnfOLCr7eKYB7yMT8
ooXNi3VPMj2RRNi/TIpMOvJ/YozfNrbNJ6NaKyZd1fOnydeOdFi9KzQp0r2nYK/2
oxOkWDIabx2SGWjHwhtzpIq9mD7IG0zwsEqxfu24G6N+/vdNDPWoQbDcuNXW08Gy
GdVIhKz9cH2xv1sFGwfpUR+PgNygGBebD3rphuA1dZfrtQYpBs0IIHd1m8nFGKtV
nxG223/pW++mKzcb4KXB7R2FQaCmZjBa3b8pHdvDTnCr9vReQtwuKaa/uzhTKtFr
w+eV62yKZDKDkJlZhGbowQPMJ8M07ZjVY26ikQZkxCd+eiFEn2arDqLYnUQoEDhv
5DYHYMgicn9mk3tm4rw46np3jY82jxGLZIh3BM62I46+kVsr9GVtq+yChQYkBPbq
Gs/BCWmkRCPuGi8IVEiSnvW7oNRMM8NBM2GeBSyVWrWZUl75tJQ+Gxuzw33XHjNj
OkMm6RVtsvfRwGarUaaNVB9dU4mPUVdvjxbSejvaFs4e9m+wPaohuXMW4YR6DXkL
Q0/S7Rzrw4w2lhMSCJ0TuLLMSOiFmMSZe5hVgSZopISL2m4QKzFoVSw6OPhh9Vms
J424h+b2YdwnRJ+B+c/QP05eg8XEqRu9lVvdHqcJ5q2LJ3xG3zHdpZzf3eEIxWEZ
QtD1jEq5uMwE588KYD+4xmufCqz84AllZAhRbBEMkmFJHLU/FXZAGfFwRuEM/ihj
fk7SoftHpRCz4Tupq7PWqjVqxRjMHkcAJuH1KysQ+8bdfI0jvnFJdltUbccrhY9A
e9UyTvnICzphGJsb0fybkDPWv9QU9tdiNudNBiWm37ZJMXwVELgrjBT+CWNAmiSs
dlXjK0iB5uQxB340esFbgtr5NcGHcBWrODmIwqAzugKvEcv5hFcNatVQVXXQeaeg
phVgDBevs2kM5dQ2Gw9LLchKXHy6gVZHzI4xz67bocDipdlsL8PQFzkxrNSeN7/5
jDDXAYZKHqWbxO+hNJQAURSKxMDQLhN6ybquyL+brnX1pmqBcJZpzrMaXAeP8m8r
KzqqLEcQdQfjKcvyYrbTlxA6SV4HxI7eLnxaRdTbgVAQRW2rsDLjQLHKQ4ns7y2c
Tz1/8AT2h1Rgz2ex9QAEmqF3MkcpvhrqCB3WMOW3v5UmwnjL3vIzvmf1Wkk0IMtT
9F9IqeutWN/O78hB/i2hPhJElBICJo5P5QBYcRMtQdDOKgG8iRfSe8pNYQAyg1qb
jV0hBL4qtg8g1FtFKHwlYQboK5AkhibKM+zIJu1QieElfM2O/d0DcqYsSLVziGCl
eue7xeqazVwzpHDBERHA4DT2VYNjAw9SLUfnImYPbNYuJg87bEA7oeoup52RzAQt
PmKJH8pOH86B2Y9bkplMs/DBIb8uJ/mXMHi9JFQCAiB7g7YAGwS4ucaSB2q7SCYs
ZHE6zYyuz2LU7EW4LQpYoigQurV+jPGumeyA3o3xpF/GSiQhkNuiau6rM+fEnrcu
5J4HszbNQClRfqnooL1pMLVKo01Gr3sF0VScrpT8YvM+epatvLQR/9Gvp5cxERnm
EUY5KM9ZcFsyGuPzjsvot2VL4oaMu7ChURCU+464GWmaW+1FeMVKnybj47EVnu0f
tPU7rTseJTvHK7OPl3u/TFycLlX0D7mGpjqCMLbFKxmz4lAoCqnHtteHINOCnCuP
FCXl8lH6WRGXz7YCg7+bkqaz/h7WEWjOmWiit0jurigwgPLUtjxOeyaewNO7rYIN
8dhpIlY1mKphwfvPS6cYtfJMWlfELtzPqfqcS0eINLowwrd15JNlWWGAttEVN5hN
3DAaAr0nQ9FIEeI3WcgkLA8cZAjAiy0UC9X9636eNFdQlO62JGQIW51lvQp8OlOD
KfDTIU7nv8bP91JRqriUqrzxV8d67foG1JkT2Meow6KVgC+QZcLiwI9hotHmzIQx
r+WUG7chrVKTT8Mv+aR/nE7lxlqfq8a04VQN78LsNsARfhMHpS35V5YQtKu6N68Y
u5LEHsC1FrgbP1jE0LQ2uVh26X+4WcjiXTEJgAIoKrXbShWRpLDdmibCx0kusqOQ
NBm6NR95w412qrKY8yYywuS+bugJQPtbaJWKwwLWVJ4kkQlVWc8stP9qJDpZPqgi
4XOLc4je1CfDyUK0pEaxZg7/fu60KhrxYZWzeYoyQ8LF5ibODQ1IA5m5c/XJLIXx
pqgL1DPwDXwUdEW06sJkb2rb+umD3EMYF5ibjzPgL2W1fxbkIi9KM9UmywPJBnt9
L81+sKIYr/hkvhGATopueJDI4NEkt5/Do8pKfrCKa+o2bNh3T1sBCJO8ayik5CP9
EbmS4Evc7UNrlZ0xqLG61V/EusWn6MnnIF2NTExLgxlsmPMjCSCM3EpIeUhXCzgR
ZqrlxGyAG6LKWXeJVzD+iesdfB6TZwLNjLi0i41QLMSk9aaDHolt+p+AjIUXhLJC
Ivk9TGadFwIoBXTGNBqXm6aLtrpHh6Rf7rTPJLmro1owLpoeiGrHCW54jJ+xmbrn
wUmTkOamZmmuW5I8tITUdU99DkY9DLZSNr4HagSecs8eLYDxthOjL0jj33uZob23
6IIdLQsGN8XPzMj8QLS0SATMaoG0ZwuqtyCHsMNsjthGcwVcACYsTBoPjlWg1sZu
7hYP6VuD4wG2iOqvvxv2JJSWCr8XIy4XmXjPacbeW21TZfTtzj833WNhkRy5PsGv
QFh/VURQPTGd0UR9yvGJyWVYG9B7TiXCQ2YfD/vpvDwMV0XI/I6eboFTu9fZ9a5w
lNBlYdRL93u8/WmnhLjsFOVy531MrC4YEuayVeb5rSQAdSNcTsMG3DminWtzv9V7
Awr7x3ma+iP6yDbMMCZixzsdK+A1b5ZjgcQhbIYRDtrBg3Xu3xtTCgElAUyqaQN2
Q/SUGDbJDaJ1HSSu+jsVK+yGMFzgWRQIYz96uRk1DahV4R/FB1x2fgDgNVwO9hsc
elsZDFQnRxeBMWcpQ27Eoybh2cMaBWx6CpFaLCqwZaTSDMpeCmMIloPhRk0HyUqA
F9PQIVqtI4YDsXHupmzfjnUTdyILNAtIzO58/Rj20Y4dx6wJtEAOiFiP/LhoXgc2
Yer53xtB5tht7EMAtic88fxGdt9bZHFhm1vARZszdqYHRXDmn2X+oHu/ePNzgwgo
P+1FgwfUnujrS6SJQETTLaspc/otkwBqJ0qvx2nDljP/HxyUx30z4xLgGyv81bdM
PepJIU7JvoTItmM7znAwb61z3aDDpWQIIsjJrJMird763Xh4o6Ierf7ElpdwdeIx
jpiGfkI7QSyrwDeOHwefTZbPf8hhJoDs0X758+Mw5K6+wPhg1Ioy9xwFTUq3hk3i
alN10rZnYjphh2ZVLwge4SGzbD6ChKj6721XZL81Z5u/lE06eOVaDnbKD68o4XOW
4byVBGTDAQ8V4zjlOgRyEoCnWia3mnSgJ0fj7p1CjHC25ElpnwHkSU9EDKnSBf7U
X44NIT8Ajdb5lM0uJDqB5loBqYFjIvDKfjvH25Y/zoVDtkUrOXa+zBhVmDAwZoeA
yWSnf/21fHdCZVm8sFGk9f6WOEcOksiWugDrN4gEf2TSwz+Ygm3K499IAHEtWBN+
Wa0evz3MdGPtkn6stdCp7GINlwmjiYRtsqa8aLvJ3fw7ZcG1ogQ5CcqYZfzXNEvW
5Sc9xcqXolVa67yy4RSoMQgrWdtfSvsQM2Qo9STqXXZI6cTiQuoX9wCrvdJkhXR/
ynRxXb5zj00rUhFuNfyXmnUlkBqPUk9UrrZ6umgrS7LX1N6MdSCjk9wGXkr7/rD4
L2J1Qc6o7RtlDq8+/TG6O+eDNVHN30Re97SkvdX3gDHWkycHbDSiHH3yXSC8ek3o
3TlPCr0u7VJRwq2a7WG1JnL45NqdPEaaGjQpOGz03wlyoUp8CLzzFnw2HMdEgJGI
cLZVD7U+aQOImg5jWepv1xUkMjopPqL4Ep04PjARH006ITXYBZUTQsrbwAFotvqZ
K2z1GsprIh0/pnfZfwCYTqxun9DFJ7pZCFlCIuHnOWsPH9HuMV4sE7WE+yI1AHUX
qmAhg0a7LhTzNsBo7wjm0eXvFtyGyx3GqZGnT6cqMaIsHzPrDvcCP6rBoKih89xd
5reCXyHPWrKEtC65xhGO+07vpC7F/yCma79+ibtdiGjQlcYgJNaVF2YywCuVgQy8
SKCfRm1+0HbVWDkORTjH6yTlTukEhGr9iJVC/tbTsBg0/pPgEyGW0uCxjli5sqIh
IVigJ5BjfCgUjwaR1vwk47cpohAKvu4hNRYIit5L76SPtoVhZlDV8pf9CgysrpnE
emyKv/AzFLA3O33Dsm2GBRLcksTOcWNmNs/ekiQjvNez5rmY6UblSQiNcaWbsuaC
nsExJssfFfaZM7uRzz2R6BkDb/3Owu9INqZn60E/eiMgt75Fg7cWfA6P+uTm6JSF
xPDFLNpZHGyicFQlD6uRB9XqOQq9ty12u7GT4GoeTbuDt3IVSpHPzSy8+dPoemSw
HUdkGe3DhgPrWL2kZzqJLGWannhVe6CKGfN6bAry3P6O4dCHLvZqJ9kYp6+j3AsV
07WHGZilbsd9/LnM+oYU3lqtjjvudef+QDBkIPywjuCcOWww8h9B2fggUVgtCML6
N7dDTZ45DBqsCCVc9/lU1KxOsfDrY0NdluclVPJVPLHmNXAJqqDOZAece5IdVpLb
Fr4oOcR4FMgq7DMeOoOBKVrtW5tZgUF8tMTUJakE+AGTRsecnxKA0Ov8lAxyNQY6
crTfsymXe+ITowhOXw4b4964tZD+0JXSiPU54ONcMipR7pGetezI3p0z/gvvwcYu
nhVAK/A1IVEmMqr8hSNsBBt9qyFAzMUsdLuTh0VlHN85JPzz9SPjRNaTSwZqfCBe
BcMiIpCIzrWM+bt2Fn+xI7yWXiCVxsnz7FeAxa/POXjPsi1CjelWCsoLLwoUfNk7
MAK2Aj/+jCuqWb6DkK/FUTcoy+1meU0BEJYd4JUojWqu8DmT16oINGRzBCo08LxM
zj3cs5CQ4Qw6+iw/RGm8sB8UU6R5wmShgKtAMY9aTCrPF1kefSqsZrw4W+RQjbHd
gBs2fvDfcgK2ay+VPRjvL5d4pj3QbxpASRhG+EFLZ43LJ9D6xVWTA3+A9fVRt5S8
WfF9YLr6WpkO8Q853ht4bpfvk6wttqwR6qwig/zP+SC44MysBJJwCqawMabumw/e
GtiL+GtlJbAJtPA0FgkRQvZo7Z7kM6DI4v97db3A8TruIdr1hdDg1g8QIhoG7j6Q
bfKLu+EKfvYyxpfnUdABj8p5b37Y3SAigeoh4dypaNBU6TsL1BLFrpd0BsYw4rut
S8vUFhF86jncV8Gzy9AMbvqMpa04qCLAresg4lBgmC7EsdVT3OD/nGPDlaAf/PxQ
ejqWw3AtZCp5kOse9yN97tSmFRI39QfMus3Wpi4v1svLfQX2EI333gEFqBRziVxb
mttlJd/GJ5FB+/aNcTnva3FtLm2N9XUAlg8THrrAYmLXKW9UoAHJmwkTyupC4L5h
tpRiVHpa0yfrLIx+0QkM4zsFVwtS6XRtNInur93LCGZIaovHwGzYnW4DBYfaieHQ
jS+5dZhUIQicrgJqH0zJ3B9j9kVBy+a/48Psr3HUDlWIqco5H7A7hecrPmE9P7pH
6NwQXbB/18CZuXIVySAiGL+geYWbXcw9p2WdnyGdRE5blon/GyauyhkqUvwEybr8
yMTHTQpuaAd+Z9YKvWTZiegLFj92OCFBWIqf/n+mekcOI4fsMaF1TF5dS9bopEiQ
vNcNikWPRmQGAFtzzhrOzdKFC4bagwDP60ROoalje8EEjnnOrI3/1ran9eZh9JxL
tqWhPiCfJXwvqQE2wRNyRFhLZBLdDniGl9ja2hZwe7NVmKT2B2Pm28uVUde2r7LL
NnZ52lyHo4xJfu9OOsAonRJEKXHULbwCq2+sXNoHuUzDEdb7XUUWL1z5uUWRdYsg
t8fiB0NcIPxCX4gZ5bxM/T2NYQCPq3KvnXIfBvCIofqsUF8bTejDfp1Tp2CaN+jN
aJVZS84J416+KjuOFVQeWHU1d4LvgIRl6aBRKxLzrmHSJ7EyWT9N3nhmYq9NerHD
C504Tq+HygNaj78+OJWP7u+7iOm/iJXzERuVpUt4npwJPyM8QYwgN2Xix+tnq2pA
/Cl3CuA2PDcd610imyu/M9d34RmWs+QEMgGsGta7c0MXQazrtuA8FrL899mBBTzG
H11+Dx9eai48UBjNwxhBSIB8Hj7zAcEaatTZQCyZaft33tKrHAcG4okDa05Lkw4v
RdDaVbFu7k9QjyJKo8++2FDIfhzddEz+19j0zdGCMVnhk+j7j6ZLu0Adw/DgdGas
v4YRfjw6GPsQy94/dQ3wx053S5tVHD6hH8k1t8TBhMKNl6Z0QjWFJyGyD5/jMc4A
kgvEqPxgWQRTlm0o937shHY4ok9MVMSyDfabvPmKL/dUdYNMp2NZPmqnLgAmMHun
XFTZYpjvS8YkBLcCpn7FO1pGNGALLMsVXNZNkY69qOP4dnyw9VEu5hXXV1Kn4Lpw
PR7y9Icldsw9Ng35hFpT61Kzrf32bMjnm/3U4oiPZmhFmzuvQ3aLv7VpuMSj2DB7
VPAYGTUA1zr/i60tGxQ+/6S4XLJod1ZgEuqWnqpXwcgG2SqkMv0boJohv/ebWtfC
sxs8k4ibcQtjdmFLCvpUNDPwLX/QIyXBPpb+OCNT7cVh7FCOFMh5H8UIkti1JCQQ
1B1hvsmsfFi4YBUIK+gGR5LJUWohOYh7IMnPQ/N16nO486PGzfHv4X/zHObInJGY
rCq/gdVdixqMZX1nZ1TKbaTa3P5jazNS1SKRpbFSpKgCm3LkytThQjMUpTAN8qpw
a++gnWDjBxhYcm78ogaa2Hn8gZ8PiDQ7uX9kAo9drnTOGvNtLMbhiBWqNR4uUOqK
JJ3Dp9bje2p5nCKSdU47yF1Iu365K9kgz/73a6KCYUVBEgq+xgL0osJc3iOPDwTz
+Snz6+HWkrw4GZ12K6C7X329WD/6N+RL8+ZV1fjxJT8bp3kgga6eaA2TlrgXM5ZC
QlRVuWNSwuSqBpaK9ZvDwnPWIvvFExuY6Y/IwtX4vEudt33l6sK2te7ufyJjUdUP
sKdThGXs4r7zSVJXU+G15RxfpuVuSTUv2dEdmOb4BIdHljJaIjZ5L60N9I6MsA5S
UAlggnKJXMcXj00TggoAA/OPetNZywcdhIp7Tx4Cn96GtF9ELtKrDH/cj4EtOj6n
3tudpP9s1Wd7Cp4c5Qoqvd6ITjzHxqUUQ1uTHtXEJJ5NL2hUkQyxo7FZaN2RcPiy
AsJDg0BJnr+jBtY9CdbgCjyqbo2Btl4Jmk0JsBgS8oj2yk4WC2av+eYQgBlcm94P
Z2h0IohxTx5DlYSlaWNhHw3hBXMqZZYiXuH08W0Hew07MEKImHlA6bPlL/yqC2vp
RXYTlPJ7GiKprWtHTfRFLHye8pEExdCOtEVyw9pFTkyM8WZL1JhVa9wyaTX6yZQ3
1NvYjXcg+MOKBwe7Miyb7TJJxaXxvi6yn5FQkqgMWt1+QgbdCthnK3vxPjSS/vUG
X2z5y9gigTJjZLYdNN0vJI2lBLiyqckEOjJKZGm7Gme0iTzvXhGDfYARpfWOqdGW
soFDGbqg4UhhsY4jXgGGZBujY7qjPevft67nyIHs19/D9ud7XLAEUDoOgv4gKOMf
ZuvOoEdjzxrdS43ezgbCVkhhcvKmnEvG2FBLsb9FudXwiYtYOiUYb+gT1bfSpp1G
rH9hI1102ZTuXK9TEjV21wVI3pY3pcNx9RNojkrALYYeT8lucvfDey7okvR2ZMtn
f1CTN7eyurxMrVgS161NIyg1yj4BOdKeTQyitw213o/QIhYFsaurr5oX0MZ2FYkX
c9oZDdXU2Z97xOI+9oKEcxHyyJPciofvVxStXRxQEPr2xCxY7CFqkBZsfNU1Dnvy
EfMh1KYUip8zlvgv1iojE0c3O1ppSuGl1bxG/cHKbEJO4kjvjZafCWuOASjnDWX/
eEPQSMRYgzEeAe1CP6k0XL2ZGlm8Q8T8HZQBwX+O8U2PfSSTna42Cg50unywqf29
OpdO2qnNhMjyecDGJYgd/VbATwfRP+PAEZlo6p7qqSYVnzk8vARjBKEtHHkP8d7e
7kKLv5Va+AQEMUN/wy539tKyomeaIFVB5QnrZHRxx4zktyJNstPDmQwB6dbAeMsa
9PDc9fd1jlRujKJR/x+ZmmkyP/wBGSNf4jY1J4/P4Ja3tG4n16uj/3Lw8P/2R0KN
YQBIyGahOAucNS0nDTO8xhmDcEvNmHx9zv9h+XNzUIWF5JnzTD3u6AvfT+MCF4lc
CoSigCuIhGBEwS03fFYAMhnmSZ8UKWFMgdt80qFawCdP75Py/IRFKuyuRKIEmBJo
Ck0VbAqST2Fr4MoEheZFPVPTj0d3JwnvcI/3Y98ggeoR9WoS4kBtQTFTf7gBqBIG
0c5KSQihQKnueh+FhOHXZN6ca03lgVpq4ejq6dKgMOg9/1YXiVTi5F2O61yzLg11
aU/OK7e5Yli/TgprzgW77bl6p3/q1dHIMRr5QkTaFdCvc3NQidDG92GOOyfhJWZP
wi2hV31ndzzdCLtbr/0E2nwnI+wFOBvPQbl4csQihIvvee7mCZFKi0qlDGTjZbg0
yIAlfruMwAnLBwsR87AVCuW0MjyD8/6EfQ1IxC2gH6CHDwebiykVVz5fG33AHDri
UXxXCHXw/53ajm7y8CKls0hLO7vWfebD2snmYBzvWt9rW/jzZ567iPu86cvGB9ww
zEKWdwjz5EGL4kHF0Y27Aotked26l3dVUOWWKBlxvPfhWxrs9jpu9fKzijqbR0aJ
JZ1l8iC8UUqQjfFG8GJ2t+rFc9AJhAMNIg/ysUXMJRH31LRi2fw2vuttYNsNorqe
xKmRz75/oJRuvz9CxwEIO4Qkdn678kM2NrvVhdjciwiCwYO4H186YHeGNtb4uuCH
y7DrMPD+8TMY4N1X06VF+NfL1xyL+hTM8QfW3o/2f+Se8+WzRHrMqcREzm+J67Dp
/4WrY2qCJxX6/XCVgdDRgcXx2YndS4UHVoDP3L5j7+2ECaJu302NQO6OdcLgb6jk
uvwRQ3VvvBjXA49CIJ/7+/S8pCKDGYZ6qh8NydxZEV6Qr49jOFa+L2jRAmBC6kr7
e0JyQxGRReuGVRh7J2rR9nW9zj6hh5GGrb24A1v7wsENww0XAaHxZV6yg9OM914b
pV9TntgB5HEzUUwSe5GoQnrIgOiEbpkkW1U4ENQMsHL+GnqOx6ufLsujfd8NlZBX
O2Ja//1854QFkG2TISTLO2cXWpTYKdv3YHEl5NSznAf0Ov0T+LFuPk3XHCljOOJd
lvBzv6Cc/z+ZQJliWSiIL0Uu1CjsTBsfSOfswkcREwEqpu+Tmx3OuNNFYDJ6I3i8
VANf8K86Y2d8ocZM/AtQ0hpr/UZqg0GpHxJBgfm0sL0gUOOum8/5PAApDwZtVm9L
wV42AJ3HxV5dDOUVCJlmOTf0z5xzgz2DFUwiubgRXVNiEwaO9lDXedYRuPxoW65t
7jtHT96BwrRV77HJrKXC+eM0wUsCDVz0tQVgthGE/MupAK+Xv1o5k8cbUYf/ajJJ
1VXr+cuThV2sfUAI5XZweIepRSwZqAzYdrf7W0UzB6b04R/G+D+WEbAcg+zA03uk
eM4l41bzUaXaOMwokf1uQsal0wpcYHqmvPzOiOw6LeQapxwwABgaTO/g5IwZiVGY
3l/rNirKgPsRyAe3owdv1nrlY3lewq562xC5KqFpXYr84zKIXcCmJ+nn2y/def6H
gXbdJAWNudfdOmZfCrtIRsdkldeB5/JBsKq+ZwiRCcS6Yesg+dClB5MfnPEFIUfw
YYMi/ONV4J/u4+ddyBoaUv8E8blwJgH5GZmHnpQFjiazaOVcfHO01ICY+EbOpoO7
MAITkrtOaIUnf+i8xUYrYkNpgTk/2tH6nV05HnwqvY9WUQHFIZpnzFgkwWwHd0Yj
06h56T9SPV/BZZQEO7kRSqjutSIFLw6/lhX5Nu991bg768iJti3uZbdEEn5GaZLN
E0RhVUmJzUQLRgBAc2VdrGIfTBvjduRu6+EJzbpiSb7LcQOc4k4+njWQq7GQwb7d
dBQUG9sCo98v03IZAPhOMJIOeWli1QywFxBOZ5QBfQFDOi5v+E2g/RmCsQ/enh1r
De8tGWXpivHJDQX3Cj7AwSjn2HNu8nD+wTZBzv4qdLNs+L5KNbf7UjDGD9Pvu40k
JRKG8rIx6wAJt4ifuuphZiN/Sr1hy4mysxArWraXfTfACvTMNvIj/cNpOnkNY6aH
uNNtRpG8H46vzS83OTxH/rVcW0UM9Z211mIWpqztuSoFhanb8LzgcEH59bMIBz+G
C9LzTFGHCNOaaRx8WpnuZ76Mqv6aAncymAEs7MLaJIw4kupmHveDs0o87Po53f6F
soot4TqNAI2SxN/Tg/8ETVtEge5equAvGIqdpunqHAb1HosSUHLGimHOFtc3grJ+
U5gCCtqOqiqmYtMDDidiOB/sSbrkcIqmGpOTeFoLQeQNgw+T/pz/HtUM523vPXRH
AIwObNDa1iMsWTXPMBUIw4V8gGCwGXswPmIblnJmuzJYqshZgT05hGyoTdb4O0Ov
v0to5x/YgDX8QVCwmFepmJ8/PJQNEc1JKKkvYMRfr1IKosq5haRIu6PGEPy6PHAh
7iNZR65pIZAac3qj50TYfOoUUqXn35jr1PJaWWxzpuYHe3g6IY6nSDFlgtabqupg
nU+hoUNOo5AdgvoaU/kCTTWnRsLvtV4cFyb+vkfRIuIoK8gWZD5nFhqLPqsZbdp+
0Mbd9e0D+EGbc6IYhWelA/qSgDNvd1N3JWZK54cj0ZwgwTAx8QWLLKbJiwECrTsx
Ra+xztAbLolKvlsvlxfFgp+bmW5AMBbqhIjypBHm5DWlPGmITZVUN7gjWxr94GQp
h5HLVeJ+Yp3yw03e7LJrEYrkgFwQrpOb4gOXNIo56PRlY8+P1vMIy2P8TKaVwPeb
ZiiP3lMrmnWfFB6nuhmdyGSME4i7NvhM8slVBWq6f7OXmaenIssyOHIWjoiMCx/E
tXfSGveAqJDXXC2wu88JX6Hii8iHzuLbnpOkmIySRwpXeZ3b+KKm+Fp+s13jxX7i
MqQBsmOzvuco+bSajVoiwELJVMOSH4n02NfYHhF/Bb5sBW3WQYehwSrI3vSfi2SP
fPJcPbUiNYGa5BaN/C6UzDOmGyN90MGqs+d7d5qc+My8qdPG1gSba+sv/4C6IUGy
xq2Km8br1CKVvilFLZbM7xPkUe7FoWrKRF9ll9ekr2p3RBVyPMwFSEJNWxny+p42
Z8KlKNiLTMSKyMbCsJkhZUeP2eczW14vliFST+2AGAOIGwjxLNT0B7Q4yRjUguES
ym7SsZdAcnnnA1gG5fnk7vibtIPxmijBEieDWSv0T3DywitZT+KOuw4aOX3mUIsX
qkB7fdJRlE+p1UKW5+bd1il/E2ps8iNid24A1Ux+NbeWitgFvS+KI1rtI+QpdpZB
YxpJPiXw2dIqUrvGMdKYf3GRRqYq4ebhSLp/nwUmM2Hs/DAUW2EaYCITYtPihK16
mAMJ9KtU7d6574F4TeSP9Sp7glLBE+nyIF/k+lFdfzOn09rEscMivQbqBAaQ3Ymt
/BCxfujxRO/pqAcLVOsm445ATuyUVbR742IT6j/0/V337xs0mTMn/YWliIrPIgrc
UVjiZXh+T7bNVJ63MF9lzAqHPrwu9rZ9v8AglGSNPGrbhw89HDToIRHtS19alePU
O3hDhpLD2wdGZzJnwr6ZR5u1suTohYkcRkokkoI2YxlLea1cK2jWLeUxALh/+gFH
lsFusbxMwHzW7l/1OgNVIpDgaCr3PhPyK4t+tcuG2CtbTxn+DRsG4LYqSwaEICGj
4k0W0LkJVIHefBV5bxJjIeUYQBX/70cAtVQgIPq0vGsImVa/bv+ylW5oRH15ejep
pWxxSeCWuO+UdwIx60Zh8hEFTYMIj0x/xGm36Io0D65SjRMiIkOy3m8xAitiHMKY
b0eiyCoIws+bU20Adkmhy2SjCypsJq0vnSUm0pDI8pOCm1FI59Orm7eFbi+Pq6lw
oXBqmUJRMhGVoWWtRWd0jlagor92FuMO2irrJpwd6Ln6sufGTWGgUPDeFu4cD/St
KU+YyuxJNSemCDKyJ8GEmne5kwsRNcVX2amYK3P2lD7CvajxwwtlMi9+Lq4VtFWv
gePcgUAGDOaIMcS8LwwFwELqZPEjU77zh3dVhwzN/IYBT6fA9stZ9K4pKlLuFAVN
NpZzQv2gBTYtBQufvFvCjjrY71uhno5i/2HM5SVXMbxh06DQwZ4w/mDMGXW39ejF
foZ6Autfu65Hfwo2zqxNUeBrPyTsWtScbFbKXw1V7GiEx91KkiT8AuPi8h7AyUbG
ssRtkZyA2rBwss+/bDkwLpzj+wnzy1IUZ8xqPSbffwNlMtOsremDdbyK0uoIscI+
pbBd1ssM+CNl4SgyR2FEhb2ehfFPoz3l89LT02E8BsaXUC5bLY1m6qwB6DTxKJxv
ho78FuSHLYbhBv+73OxXUyRD+JB5w72ITDhtpBN7Ldb5Cu2lsIziUYsXnaySaQXP
7Hhp23S9dHa4NONyKoy/IpsjuZ0g8p0Qe6NJ0I3LFgfOFeX2NATPEqUfrhO/nwbX
dMheQNrMzQaeqDsY/Cy1VMVYycUi50a6zid5/C/7xkH/0YU1gvlAvE4r05ZJgjnK
FEHuflTsd/LAbeAUwcPuuyyPa3WbdJQZTncjKpuiqYqCaKarTctWkY1za+wpMbiH
DasbifsA4mCmiHNiezn+ccxQ79q/VG2Z55GaIBiZ72iVHKQSf868RmhhpjUyrokv
FxiebuJbj2sUXiXh7q2lxRGK8LfyKt9EUm6cQq9IQu3jSEIGfJH//+KX+6sD3QZj
XsH6gaI3aLNqFUFcwsjtXK91i7w1DJNZocbg9WNHiYzkop5KKqj/HXUVI7naJDIZ
vQNrtirgXEcP8NEajPr8pl3je81EKhjdjPvB4hdKbMrayMDu4ey8QI4rrGzKgBd3
Zp2G+q8uCZ1bmXd4d3FQOIINz2rd0rB2KaiRQVMxKYaPi4MTNQke1Rz016hKQDrv
Jd6xRX7q4ufp9/eVYI3ZlanUUEp3heqp6pOF0ON1ogQMZApEAYZ4IMExbYot326Q
xHa2WJIt4O9ueL2wj5j2k9Ve7/+xGofe0ttILBn+6FWuJ/OD9iW8gDJcOJBp949A
foac7nupjOMdtt+TDO4axeZUFn85F3wH7pbdgLqMynTWxNAeJyS95xNWt8LgVjUp
GpEJsoE8aoDgDyz9lAxmOK2W413fkECNJXtgzfESSu36vx3dXlv/sSUROJQ7xBr6
FQ8pmtWNcBPI3R36Yfj+qyunQx7uzcvol6mScd6lt0Uw+p3Cyj0Xp0T6vVn/CV5x
P1Xpt8QnP9CSBG15SZTb50G7119pQSpJ1zufpmBLEpAiRnl68vkR/D50SxgJirc8
21rhyLyi8Cnp585NHd03eapF46qM/tgFIY8mxyyH5nw3+MvlufAcjF0J6/kqRwU3
Vv0MZB6rddUUklEbtLaqBrtewNmOO68g1jFGtuFrgEWkPNOfLgQ48nVNSAfTl5rr
WfWM06PQTDN66f2IMD70/tH5Yr7IibNoZFOwBc4/aNAGqNLd7W78I0tV/AwPovlt
EZfrFqCmbdOqLjzN2Zf8+WCOvp/rlbZrUNeiEptDmqp6zR4AgqtEY32CN/yAgi+q
cBqIxdzJ2LjCoM/6u+0zcMB3Ga7KZAijfrEY3i5MYyNcgseSXTijhYtoNilX1buL
3vdcaA2rXaaJJuDywyc0Q/A4uDDxMyqG3cKuuiQIParTmSiu6orbrGYsKC0ID6lM
YWRsLOhhNdhQBAbZ0ZzId3GriQ8+C6OnVWS8gJHfdkFku6ViyvbTY35Pjo9a1Th9
EjcAtM+lFHHOcXCgBDfCmT0elmZxZSvnSTIcCU2dSbpTRU4PiD3yL3YidCpX1fnU
gQywbgue7HKyA30A/WbUgMEfNDvK7Gx374QvOR6sbz6/GE9DkGs693YSFLF53M2W
W4tLvP0GiqjFSikN+gfDA4dLTWPGi7wIAO7yV2fAHRIW8h1Xah10tOeX/akab6Xd
Zda+x2GXuAJT8By47OpWssKpPsMojGpXIR1216UVKvas5u5w3KEuSO7XfJ7qXol2
mufxB1+t/Lf4Uu6Cga6CUcM3bj6Asb0XAO5L5D461IBH2SgM+DrjBSy7gTqamthH
2FbHMgNhO7LZGj2ww1SoBI12wfRXq5wV9SF/9X1Oxi+E1sEg/U+vv5EbvB2tamXS
/k6UKiZ5T4KnjPFxqcdDrOnsWmjOWCo6OnBgcYvEItLmx4DHL9e0m9CLw58isy4W
zWv1jY+gYNhGo4CwdiIAHJL0zmeaswtnXdrcGIzeSCWqcP0Sa2yAu52Gz21GkbzT
g6ZOyFkkSMUuaMBSlIOlWQ7qStHFmO37l0UuJbmvjjK9ToM0tiNXoPjGGMUk8gsn
w0MvnxdRKAsl7fpHxSKiCJnzziMoQJk3tWz1OXlKFQR9VHNx+fmCrS0LE3ALWetn
uw6HmeolcwanbfpMAvtMEPo1C0hgy1dkMivTv7Nd3dgymg0hiwXi8WN7o/jVqRPw
Y6wq1iY57f6t4ZKmALtLnwFpV0uIGNKijOAprtwp9rAxRdiZ3v4M21mALNOPpyJO
j3Z2aBIOeobpjcUozo1DN76Sm6d8iuAgXw2FJyobYslGfVGodEVqt1oobnDB25LV
ezGewutSix5fv0dzLKbtPSBfi+d7y18XMMMDPjWJgiebxSoyXelh/QIjm95SkL00
hoEoPkQ0bPpXq+wznBrXvHM9vw9O+od4dICnPOO3AC0XWHi/EctCb8xDAyj7VBHk
kI5Pkg191uvYM4KhasW+V9JWjjzvEdbk5PfIec3w40OGUUFYAOzQ+gQ6VdfL2Hjb
kUuhJ8t3szhqp0f5nRIk9c1tpLDAoC4/hKl6lc42349hm8CyRbu1b3QD8lbEr6J2
In0Xhovs7Kp8ikCbtQ7iYCfFJykSyDbTDAgjYirWNz0obnLztv8A6Al3gwzX8kYo
3OVKn46yeeEnVrhE9v2MUPCfhjn+9dh0I9q65ABG/RU3pIIPika2SSGOKgFJLF+f
aWaUhDZsrjZd5gl//4SHMIWdknGblwz+fWQ7DL6JLMcNIzEE8yzW6IqYB8vwepWw
dpVrAAXeXljb2OgmEwDHtmu/wVGJBR7JSmo5cqC4q3OeZl6rdwVhn4BhvwNn2KIr
fuqLd/F7+cZSxD7JaWkJNP3jY13D7APezecZL3o6DTkUXdStOQjr31i+ZMIZr2Fb
HWuqxR6JzeTm7akWqGbtOo4sPfi2u3qLE4zhoQyDOn289USYGR2EnqHxgkdn8JVR
7JgjUTkwNeHgA9YccBtQPzt7cg9j1e7UJW7B88PWTX0IEuJikEcSi6DZmFB+gFSB
7COMvjUqjjpFgQii29inGr936nRc9qIAzTDcsu1WWFz3RfJlaQPCFFrUlx+Vr019
TiJuW5gRxNQwmwAYSi1A6j5fsI8JsMWwdkwTU9Y4G72MGjB5mPKfAc4b33tN3Lpq
OE9A2V5WyB+6F7UdJ/iqp6QOpeIm7qzIrclAl8c9NPptpBn/LdUcMR5GOT3KVLyV
aCT869AQ8ziSgLFSH8nR+dnQdoOEh4sJbKdzBM0YQiJma4if9M2hGLs0cCD2Mx1z
OMkSKyjXHqSkEuHxbA+8go4ckv0sQwFzZjGIIkEWP+nXX3No1L55pXJG2UvQ94Zp
FucIQutxzjytFZ/ANy9wODWJ87Lf8+zcAWgnnovJJfyAg6dZln5m7NNePLYLL1VZ
41c9jQpGX+qP8FcqqkdPvXb9VsMT/MTT2p9z1O3/6+kIZTqHfv3NoILTbZPdiz+A
9JDYJbqqxcLzyM4xyW8ZpfcHAByvL7RwgSwFKvxQ66hcjcckrBqjO/N3mnUpYYlf
/9QPeV2ArEJpcD8zozZWAKSnCVX4TYhxuNFAip3eclbtHbJrLw+H72lTQoFgcOST
SRBC9nZSynoOdB2KCiA/aRbjV/T3LIiGiXCQvPaIbT8A1j1sJpqrerrH2bV61I65
sYgYkRseQTOtTh0xD5fVXYDBYiYtfojDArSj+FH1V45fi4MrxglyG0raDb50+xHA
s9ArHI42b7Crv/Tzv3fMw2qd+3gV8w4UnGQct2nr7xZc01di19E8iAlIg5fPknDp
c7iE+GS+JhNIGm/mQozScieO0RRa2soLPtY9joJHBIWFmq2zg0/oeBTDVogq0DIR
ZFU0sAxrNSfoBnLOMwvQax+HfxEZczxfurRV/rEX94zCuzVw6O+BdtnIWoqZJL/h
UqjtLS+JncfsgAZGzilxy7c4s3GHB/HlHiEp8dBqAi5hFlOzTtM+GMY6UxRQvhN0
F08Kx31H61AnPC1s6KoSPIeSitlkId5uOY5RgcUj/HZfZ4uHj07nWt+TMimOqAiS
NZvFB3VePpDgMQVKJqken1axFy+pLYiIZLCUD69QYNe9Ta2cQooVSe5tlasyXuVW
DWrCxlGMLaczI4AWGPFkGXywMIzmFg2GE8eex2CgIbVuPBXvCvwQHi7P5/nvQ8mB
SAD7fhtyOSU31m/cDGhri5Z6xyhe6ppVjJo5cp5JQRZLo3yEMMLQvDTSB+0pycZd
IMhWbyCOMmjATj7YnJz4zxEsXJmutdakanWaJydaifon53WkFfY1FcBxxJAN6eaV
Rwcuki443j6mgYPUqO1/fcrQqslFPGLL27X3vJ51k+lsK3BKFDJF8ryvMSsRUQJc
57eLcZRAigC5z1twWiht2s2a8zODu8vtkxxOmTjGZtPQXBtWO8TiYjETRipwjWgW
tECF+BIFVxJUlOqwEq21P2LKD1Cuv80/Zf0Jo2PRvdbHeUmG08SFdgcoxgQoIUUE
4V2aWky9AUDkXgBxf6wRDPtYQURUHC8mlujoM95lCESbLq8RYGqHUtznswiOjhx5
nmOW+9IO4SUckzTarTsIm6hCXq3tCtTDDd9n9hsN3HerG00h4qXIGccJnTD1QY19
xlwACHwEpcbKACzz0bUXDGtBSGmv16wdRP5ktEImY6DKZYVDqjFdrA0cl8L14MaN
7JlLbEn94v4xSihIsioq4oh+GTvGu89qBUvxaGuea9wIqep38UoL8zlyt6r5PoWJ
ZRubcMeg7OXFaohyIBuAkuGb2+hOek0BlRHyKcE7N4umrs0sj1fAtzlqJUjofaS2
dwHaqWHaqo6hMjKGZP/DV8DF7Hmdx63eGfJqtYagdP+S/awysaVI8W6twC5F4oL0
/Ix9uHq609Zjs0HMxWIS72ysTIexQPKDuNwuMt6ah9rI/xO1pd6WibyovhH+S6LV
H0wh3bzhL9wC5/qLMSAVZBn5zW3mZVCS1N+vpNbe8uUpiUX1dxFKIrdCrfLHVH8+
hm6y1MyTAd3SG3ZFpPF3BcmCKhCv/aUP1BUuZVoAdBpeGaSv+J6xgvEbHJwLx9+9
nQdSOXsvs9yrlYxlF7HwLUm3K1OQLfx6EOBBtMtiblxl7Gs5EC8NUKvB5u52FjLn
fxSx3CVKzaaETvPWGI4sQX1XZpROV5Cp6xwkg1jjZxeljnIKAET6i7BbRs3AQ6QL
RDRRic+D2zb5jyBKT5DGfXwzlbsEsoMi3bB8xJUjdD+T/I+gHKwLx5dqJpq5aK5i
vPFCU3IOPaYx86BW6rHLQv7J9qiftEjXaAXCIYtr02iJpjzaNpGTa2Fb9NYMgRLo
rUuS2ieHruEGllZD75T1efzm89wCUvH4J2ddkWo3d2jbJMYnv0P4+A9Bww4eeRRP
JFiR7Mra2o/8phXAX9LxgDyhuyvIF7eSoNjBMrRi506OGimU2OxsgloORaQHvaWd
2U5XhrCtvZtadVZx+uAk5bNkiLmcM8RGxHH5+kdUV3RqKAIAgyzhDEZsKR3bldbu
ACciaQDKZIf9uCUBiBrFT+U3Li19OnTBQG5Ctw1U5/r2FTZOCXu8Iu0xd4UC++OK
pVrXSr08TtKkk6pfuE/Yipqsm76TZ06A0NQ4Z93CnMMcHhzpFqwrvOcF6g8cTomz
L4JV63QCHr3yhzGBVO7pMmZ+q6tYXX8P1xbWyIP5xKkLXEDRdmZC/D/YEtMYe+Xs
26JaLUEaAjoCHXCa99OB5CwwreveQxcA0cVw1flCig7JqM/7NTy/iR+nSUXx+42b
HcnjICDiJizxxvgBUcqh/BoX0L63Fc0EHgQqBdB8WuUOpl2OjNcIQ1kbMwwuAtFx
q7yh4A/OnTDII0tAhjqxsV9nOEjOyHcz/SCmmhFTmRge4WcABJKI6IhhhbHS8Ffg
zZI3Cksa+zoQhu3U2nzQzEJhBAYJYlMJ4HQjFH20VJfK7q4wblA/ZUpPmvwLIybT
jUXfQeWQEPin9Vx6jG7Ov18AQncWrPfEUR7oNjz/PuWIw2+vHBnTSlTbKCwEawKw
1/9b1f6fPosGFLoHi1Z23N0KYXdu5bAU6tAtPDv+FMibe2+M8xx+eC9ZPTPWiRwR
06k8F/ojmlCYCTT54A20zs+xBacxmwG5kTPwLMNNkSP6ZtR7Yo2qHBP+8GCpdi3I
OD8wDJb+MleDI5zWiVwRd33TO27ipdx92ghAkJsa8nZlKhTqgSCOD35HYZW3Qvd7
VR+GdGdr/bSHRCG2wMVtfsey8psGPo0GLvYR6FsLytmbWLxXpTAdkBoLEcMQ5AQY
YsQYZ7cGN9kYqp0k3pjfdYKHB8T5NRnL03fUSOxdO842p0vw/biUg0AzoBZj0NC2
bxZ1TSd+0Rhiy/ytsiDA0kFm/zWoqFhZ8V/RkDJQBhdz824VoslmE57PkHmTcFh+
ane62W0n3JdzypztEybMdWVR4tTwJUnCHiCgP0fhioFGUE7S0eX4FVsZlPXcUp9U
LzLBUNlN6pcvTphbqVfG75cSjD2Atwkgu7VKdwprlmDwAFoz0OSsTjIhrUmdoMsF
mB9guZdWT60KG0o1z8D3TskAVOCkFjImCteGXKzV0rdtXP/UOIQHUOiuQI5yoMie
ZG0U2W4lHT6SZopnK3X1uau9WReHp5TtuGM5I7nnax1vH0fYYEXxAYXJw57pr3rG
pwxzuqSK+4AIOswM1WqDnLq2D/zD4CNufq1ImLIe92VJYvny2vOQpYvbuqZF0Ubt
7d+TRejXJixHQS79WeW7I/sjloYWpb7DjVRQQprscw/RBQrlbu+5t6NRu6AO7vvz
g72iWy+OlNOpen5oqEdU5hM042/oRnSwBPYR+iFG1XK63GHCydVjRoiuSGd9RfNI
IWZJu7uGcM2le2mSCxII3POMSyVENDZDSg2RsuLsV8JAOKrw/eDJG2fkvFHWNYo6
jomoacjxOIq04bArVQW7NjWOzF8iMt6r6W8ycjBTzw02Ba2/XwGn4bKx/TxKZ5/H
KMYhtoS3UoVroEv1oHVFM1GOW4xTL9XaXLTTxScA5E9Jal4fHsAUdNXOUoyLEAIf
PGdmvEydK1GtUt7urS/1/oRW2jOfoT5F54lvE78CCvViQVyPTcW6Xrqm+7U9cnPH
5WvsuAtm/gV4jGNMxdQ9uWsX4G1IHhQq4UWux0QGxMjIkbxRezLSkKkuC+1rqQQw
Ddj5bQIPg5WyS6dA9ATdfUTPckYetOsmAUAhAOAE9zP7kxxplSlMM7Bkug/Iaeod
reglSibUvZMd7VagdJ2x27TSjoS9S9gz954vy99cwEfVxFzmqHeVuwnjo725EEQ6
8DhSATwqyJ/GLmfYm1HTvsFGAXndU7ZC+3ZRZk8Jo0Y10zhXnWP32J8AoLWdQiOv
9wQgPguEprEfYqNL9dmE7l0z/1m3VaNxJd/a6xtm21ZOHANF6NNiT61znPYVMCmd
pyKQ0tk1blc+kuc880nsOadIq5/Z3/gDZKYq2/kS7Iojn7rz9PvIRO91FLo+ekvP
k9iKInUeosWIWggRKhKSw3LD2iQKadi1sj/KYSxe4RceIBJEQYO49FRFQsNk06xC
8me40zFChStYaDCNB8qJhhHYsPZpkyrPLvBtxZds5smRfwCmnFLYAd9wVkyw23Fg
Zz1V0NN0deH+il58jE7vzp2MtrMZJdfytv5tsjl+Z0ujZFQfaYj/QFnkslfnd7sT
OLA6L7kQ1aTYbSGUuDC53iCzerJPURpQIVgqhsFlEn/JAsdURknlcgdxq+fwR3rC
tYmnqh/5eEHzpokuYXcxF838RQeZoAN44a7dxRK3JdF/ls8f6LXgFM4BXd2S99Jz
KvrF70FNLRllL7KRnZJl4BxDDLSicDHPn5tcK+1rTsUIRvPSpbEZUEoAtLp58U9z
aAzObKllZ1No33cOwR/JoD15dvYF5HFU1D+2HepVUtAZ/sV2gN2kWdeCrMVWoW/a
W0Z5J0JCTCkDRAvHML1Uk2RfLnyhkWU609rWG7i/c+D1vn86Sth8sdDDQRBKEcqh
mSpzGBcSGw9Knx43O3BCNlK53IeEjB9yUxvj9V18o4QIQlErXi+embfSqNGdhOxd
YMQfxWFg3WOb7vir37khiciLsPmSp/NJGwC1wZjPdtlOrM+D9p6ra4JjRzZTQNRs
hGddTAVVNcjsfGrKJzmyjXCzlk28WvIf7iZo1SZ50Rp4Icb6faTgH1vIhqjpgR5k
eWVNeeiJE0KV7OWNqpXVrVg2wK+gW1YtqRGg6maSX21fjs0LSeZ3ATHmwtRBYDsv
m87AqRu6kYTUWiDi5MzYICK05D9kSMMPUdjxcXWjM15nu6P4uv5fFIuXsaIXm1jD
SGOCNoizhiODoxp6Z/y0dgqFe0QGpQXabTbq2b4yvAHxHdWkMhyP8pnxGPvFske7
0R9Ti5YVok4VF7W0hVogp0tu6VgbaQLRBxemoxNWCG+NOqCZzfmhaDoYaGEmMLbN
xZ5wAbVDFukgOoZhyxiqCL2RxQwqXU2pR7iZiXuk281YPbniE/d7fom6eyuDfBTK
K0XJjd3LAzzc4/lQKdWsiMH4pvvALLfVoquNlTU78vMLgs9IfGTwghVVEmXUWbAu
MBrbT+WwiLUX/Ch1KRjAIT+/NX8mn77B5nzU0gC9Vc6M4KV6xFig91ukEoeb31Vu
cTtokg/dYgtLIYS8YZwOHuzdbZSiSteJuf/d5kHCD+t1pwtbEdTNiHXwkv04bPQi
3Tq96KrOvux1nYpZT1XE1g2YkCbRlm0Z/C3RYNXcGgnBc5ipRxS9S/VQMZrwRPhu
ygh4Xk0PofpYnE4dEwahA2FSZoS0j89kCfTtw5yFvsUF1j9SiHueNS4DGLPIAr32
QvIFr6AzP8OgL9Tvy3mA2hjDjtrpZDHKzo7A58JPI3e4SxsGu5yArWOUWM89Ok7i
bg3Pl+G0DDkDq+RQ4gvzBoeULz9APyqTqiAwLsnXDpbmaHqfiegyNLQflE3J83vr
9E2cvjN85XwaELhLMjaISeRwrQr0YwwP6dFBVjfnR1V+YhZuG/Cw3ZAG+hiH5aIJ
HuCLRkAU6yRANHdqbYsIat34k3MNsPuNrh73NtkUBs0Muz4LM9PYmbbaLMDGSM0X
Y19wWSfoZG+r4Io6KgrLAMltCVgHOmQOXFA/+cNU6Rhr4+Y2bVfd9qIh0sOy6JlX
yctPZ0LHICiX8ckHmlQfAR3Zxvi+9lgnqMd4mwNxe93kau/xGyCj9yv0MTzVZJ2N
itxPhZgrntGaicu7CQRxa4qBemcfQtCeJV2Z5Sc8KKZ3YksRFKNCEUx1INabVj7w
mE6NYHgSKYEEDXad9aqvtZAqlFgB3Pq7QeynY/afXCi0ridqsjZOj9RjJA7CRm+0
MFYC/l/MVrMQK+NLOXrvEWSi1LHvCEx9YpZY75sw4+oWsVIwP0+a3t/ZAr4CNNA+
8wgqgKuC0EpVmmCsv7PkAcV0Cu+T61NYhuUH0OaLiHgDZO4Yqh/ICtQUZZkVP155
HPStdWZ77hEGkl71aLj4gbh12TmZ+oPYw8YqUdmAjS+k/dK5gLvYLNi6JTyUooBS
FmiL6nKiCpuzxwmfr99Gd3anWJMn7XWoZnj4jtkcqa4jWii6GVyCNuqkaZEMzO6E
dQxaUVkzV1LM4E91jBYfjscKB1lAP/Hcz1wHZj1b67GpDBoplxBjPWHM9l35uMN1
LCrV0ISLNsrN30ny+9tgpMuMJ4eqJ43zgtXrNHHP/mpjJ35MbSPGYUnTe/jsWrzd
3ZJH7k0ZYIQc8GPkO2yVcdHPR3++l5BH89pPw4/pzHXcNGl1AnT6k0P3MyHi/Dp8
Jyj4DA5PeMN5jHZm1EIQBlPQHPpaiK/Gam6F27ciU/NXFdkVvqN2nKaUwjHjdrUF
qIaRxnv9ZmC+lOxqEQH+9Emm/oBOYr95y39GlPyIuykBsIMzC6mukKt+g/NrKZsC
N1TKA0JHvi8zqRJP3bm6PDdLpU5Jy1CND94/cBl4JHPLQrvu6UQVNdzTus4V+GPX
UWwEtiUlBLSypWbHnCvqVHk5J9g7O+89/JmmDUu/oB7uG5/2/O8MWvofECGyqWYO
qMJODvhnaQ0mN6ZxqXiGLEEuj4UYYn8xNaCErea4KkTrjnOogd2nImKY660eR0/f
wreuG80uMVj/3s5MnYo8RJJ2ijaC1ZU20IEj+UaLP01aRnXR0wb9dcttSGeCHjUG
WYPwC5VR5rPF7ljpzclRQ9uApDYhUcrKm7qEW2vleJfQVWCkRCWSkD/zJ6KUjkb2
1wf1PMQBmW7L0WAuenDb+8cy9rvBMaMHaDVkmNf9FGbmiW3Aj5synUWY0WERL+Ev
10cWI+tkrixEfJJ99y49PzUOGxSZYnFsNIdju4A1dMr9/mWmbU+c4zD+Xd+gumDM
mf455xK23aJYzaGaV09vg5HF7QvZrf1PVx3Wm1HnhZrK9dtMo0KROJFNOn93RFRl
/gaLGRND+mGBIt4ExzS35IhKdlE7yE3p/ib3O5kWHbV2SuwQnPdgAjVSmEWT3Usl
cT85NLaRweGwZANFtcitKRKi0d/AC+zg33EDQ+lXfVIV5908FgrdWL4YHg2My+zd
nxxxXIwS6HiL5crge6pMdp2s9N5BNtMaE2GqUjDg9Tb/iE2dIdD3NpjeZ9viWw50
c55LMJEDZoJm7XbmezpDkdrvTjPtQRBEQxP2fBXe7BB+rMmq78XWVzcCInvWPK4s
KN69iJwMftmGoHDRWchNxRkCNHGaD5v+BnEoa3KXFYYa+GfJxYxCrb5ik4Dm4nmk
qekJ8Z5Sn65vNKwiBjbm7lZOPDQ/AsUAemRJa+G2wJccT1TKdyAc570vmMnW0W8Q
EkfZuxRdp9XiZvcQqFjjZx71ZcPCjmkV5QcibgYJBDMyeT8TDDyfZCOWHoNUnzXe
aotqxPK5RfXJKJbajB3Em+/ALiDSnpRKPUaXLlIOWjCZbuso8n+HA9t1amQcPyyM
+jJjN23o4C3cdNeUTHob+QmVuNg/ymBcp6tlX7gg0Hdq9y8mzHkhlozueFmko1hQ
lgi228UdWkJUl2QmXCItRMD519L/WjREfnh+ShjeUsL5hQOYmCy4/8JhafGUrgEX
TO8coHORqNztH++ABV//9lmRFiewtSDShXPJ9oWoG/C8JrhqVLYfrrkThdT1cTMt
lB6mUbuCtT5yx59FgV7ta3dyfhNkMCgYftM77ca0IFp5C0bHwvlbJNuTZel9rGk8
ehbQeg9t6wZ/hYDamVwEQkWZERadaZDIaiTYDZ/0p7kZ7nhr/RYKgBgVYw39BQb0
zkvsgVpR8i5Iw8J1D+4xG8h5EmU4b3h+eAr1+ypEW1narnZWw13uHQlCQorpSvJg
Yw8fWkgCfca/NkHmxMa4wFqvO+1zQpIwVWy7tn1GUysDhSscavTGwcfomyjd/LzU
rn+fGSCVZKrFE54V2SYveHWa7eWDnZ78/hSgJjMEGXmNC42Qx7MrlUPtzdyhs0w5
65OCYotsZywFyraOGdJ7f0AOmzpja9En4rrtPUa/MHd7mS/8Dwr+LPP1CTmzkRvj
VbWoITXOhQWB0UuwgAG/Q2cAqv1yTRNn8sZPNBR4bXNLUpvaVJOkbNAwrAz6DHKW
`pragma protect end_protected
