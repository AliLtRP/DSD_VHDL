// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iqE5gm0AgRpIPlcgYemZugHuRS22pf4WMVU3EQfaUlmG3n9X8lfRsH5xKKBDvADC
1GbRIw+glpNex00TkTgq/TNVU2QgyjEpYdT9XO3PEjrAjqCPEV0fpaeOpxNILhVz
/xFdIQuPci0m7NsXLFvLSWtWA5gbbw/gKJh4CqvNUc4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 88992)
CxJO1KB9F1HZ1tjOBbR+MD7f0jo19u+KmMIn/1bX23x0gRur8gvVwClq6IPGhG99
GDDnIUU+KExktoAeT3dZU1jE9fLnsE60ylRU+GrqvzmARG5W/DyieAlz8yNp9MdR
GRpkxzkxSJ8eHKr4IVi/1twtEbzPp6aWjtrZJxwy/8Y+6qILF3MzXHxUyp9Ee5NU
rmWQn4GIl8QKnNG3NgUnuXp6LQXphi7v3Uav70oQJXlYMcWZiChdaUvZYTxfHmR/
MCv72kS6SG+UyYpxRYj6iNqEbnKyshIhZYXFDZmsS5virQgj6mgsGxHy7ABK+rzm
JStRw+48Zs08CkY8mh/EuBPQiMT3s59AZ+QPZKaN6SuneCxsdwPHONMjtb4tLdm6
GC7O7f1KYv6PzrABAqp7rJSxqSz/yE+mOqANQKHH1LSnqFaFM96ePI3k/vBmlQWU
VhkZZc0jGfrwdBOja7REdzuWhapcsg09AgLZgwGRd6DWOf4U+7McquifHcaX+qpk
5qPJVIfpUBKlESoXkgPxlLCKz/+LXdyRpT7mmQibJhxz2b4xzbb4+FofVg0tdk1g
Kumsm+SLlOZJJTfswYf4CLOIjjDd9HY6gNN84Wkfcpm/bADbMSGdfp+gD0GURKRq
NCzdLVbW9e7LlYQuh71Z7m7bhc6UPNstT+COsgDPiSunm+4EUEO2jXnwtCkyuzRb
5yOse1Eu0iVEI2ipxt/hlrSJIjO2e2A5QZJijfFBdM9FYv2oW/ePJ/GOtPGOvjH+
v+oXbtT/KML2lezhisydAjeJet945Lmwkfow4SivdzrvVkO6Z/7KErw6bI6JXxV5
9MwEsvTFONQL5dxcneFrY7UdtRNYQ0utZmSUuwveEoGUwhQJ8atyjo8TZxBc+cZV
vmX+7ceQgVdAojJVsnOmWot1jzgKpwxlCoK+YT9BkdfInFAjRC7T2nEjum4Lf/dm
TwEDRoP1QBbGvUVzbmA1wPQiSzWI9VuksFGTXaSQn7lAYrsaX/dphc0U0swmp+Tf
TQtc71AcA2zKhiGmBU+J+BlLjF9G5P6kAN2xKL0ECN6XEGYUlnM5dLIdslFectT4
JbboREuXlpp0pxzyGSjGFKZtTO8u74l/TuaiZE1YenkapOa1r6DtR2c3+FsnXMf3
udLj8QacXZBkIfY4PiFFFV6YPLq8r3xX2C3WQOF2u1lN0DqJHPYIFZUlqWPbhDab
ZOnZHFUw7NWeCXP1rgbBH7QeUp1BJJAZu4KrvkfWNGiTmBZuV99FVBtxIg9spfjX
lDG/BpbgXu7f71V4VqriSPTfzXRfsNyZ/zpCDn5tEMeGTprraBMWZHf1sFlt3sZU
/gLCQIMDyCw7E6MyB5/a7WXZoAWV29n+CDO48LrFiKHqCVrGb7vtf3sVdMbUwie5
YWOztlB6uwQNAlxWeEItUoIwLlrhorNKdJ9M0suOuimkPUwBACK5IGzM4demFlMk
3CZD9pGcYSN4FjmOFfuZ5btlTyTAXBkeQmZPSLUYnXLMdSvOcd6bVMERL7JvbNZ/
D1M8/IFW4VMSGdpwTrBp2RsfMlhV+sEdDFE89PWii6UXe4ChWmUWX8mhdPFTtQjq
z0vAB4KoDI7OhZwROzZ/sGYdBJYQAsV0G3qCn/FTnygmL2kZjLNBQ4oYsiX4D4wP
4sSw9vJOeCXdUv6znK+IDln23zh1dk9T2IGfYQ8FPSIiuRyGcgBSEb5aiixgRDDT
j3FoVZeMzmHV+K9yHBMP0ZpgwosGGXEu+T3shx6qZYx/o8uCRPxuXmEOkV+7Hrzh
+CAiLSx5YDAC+JE8TNVvPAn5y5ttsMJLSdZboSxdCwUhB6+qVmFri2h6w+VGAhyk
yA07QMiZNzHe4r2rijS/pjpbh/w4+THgVzXNV7/u/mLUssJE9EiuAQFf/FKaHkvl
eRg80uuczeVNMGSQIM5irSDk9SJ7hJbAMWAfFmfuPVZxUIC8cB7ZCxjSihWrAeTh
HcUPGvkaZFuCtGDyevLOm+JjB/3Z6ZMPEy/4gWh1pXKNNkNNk+qOryuS0RUECBsB
Nj8di1LAK+w1/kEC0AdLdaMr1jdmwBUBAUfBTC+HvwJjk5INV9u50oiizbr5j4+J
fg49nf7+nMfFJ6k+/4Esg5TG0v7vVNzn/3RJ2DWI5FGU7filuV8XEziCJ/g+m6SB
lIhwR5mhey7Zz5ROQPk0uH/SAXLIvVPxm+j5l5A9GQZkGSh6wZm2rrtDjZRsJj/h
Uhze+O1UEGoeshaRbKAueyWNaIk1k92eExKOfEDbMi9QlSoaOsk6Z2PvytOniMdy
/Gw8irp0eO9eg9ohVxunjZHSKLU9637CMeWEIoltiRluOZmutir8ge8ZJWXQQnh4
rYmQ1VHF/j2jBwLXfCFqIr8EWvnAEag8HpMAZgW1JgPY5eor7zz3x3aGmJADT4+p
KPIQJFXYMgUw7hM4He8ZrCEqA78DUs8Pp7co8RMhoLkH+OUrC9+IvG/r0YgJcoIJ
dKg9UA54MYve10oK5CqF7xm/jeDjJgPlkcdNuabfk74AUY6KCtbp11pkxyirQAlQ
u1uE6ICwpyLkVQYY4ZraCBXYGpX2+/DSkPVFHQoixRDSJyxrrXTMe1ispaiCOEdy
b192kvQLuDETaM6Uwlzo4ARiNuAhEvUg35a5k6UPM2IZ6/dcT4W8VQetiO+pDqhm
qQT+6etQTRPQ2ma0YmvVaFoVfplsA9cu9Of8St6roAcVTelmFlSECzjrnVxd7eob
+YW7U/4I9VyCLPcZaNN8KsFgKhDq3CagN+MuhyLAstRKUdwv9tafzJ+DoscIaDRw
rcg/QAU+1beB2snIjuCb6flm4BNTDbPhbxas7RJlP57QXGlKSWbccm75RU6GQEyk
tGcU6EIaUNiwmiDRoQivDksAGBdWZ2El3jhN6s8IPQTRh8kAeE8uHwTK/hrX+yiK
/Hm8RpPFFtJ3tb3dKF7wu5OdV5OOYQJldmWusOqUA+lZ1QOepl09IZgIS/zk9Z4j
2GEVlhBILKEZtVdvPDXMSffVMrh8Bgs5+EXumPStXd/PEc6EJa1BikiggJ8zRe3m
ZTsMWegZWjmiC850ssbHv7z7X+bYLSwtBnAf1LRHtyxcZefm6escA9qKGGXLkz1z
spLaXjFtPJNN0rifsc2pf3VZc8l8V0ciINaZhr/L7U6HdpxY2J7k80foZoBSR9Mc
WSPQHF+4Hv6ZKbXPbTbJL+dY49UO5anDAQyzNeNm9mTLPZe+B9feCW8Bxt/O2nEp
zfbaEBc35uYBl9Mh6z0wOjZEy9TDLKc5OxddeVORY77lvLdoOvzrh67ieEZ3YHh6
8wXT6fJQJcshuGMtp+84sxkDxEgYtxVMAKqRuWuhrUybQvCqxh8z/6t9K+bUQss6
NBtS73g6oV6Xna3T+PmianiDD8dFTGIfZkn/veal/ND1kU0wZiBKK2OAfaIYrS5e
NFyjdu3W6zjzkd0pbR6/DpRHIzCfGl2Xs4oTjmEfGQHPwaHE2tYu+ICVKheovdSb
tjWbBPVyR8qNN7POgitPLQFCm2RR/GOO+ym5gYrD6i7onJoUdKi8koUF1elmason
wLZb849j29xGUHbYxXP+k9wEVE0veH79D25ZSYLIQMv7NCgjl2WVvZpnu0G9nhYN
cXL8wfsuSMO6U2ziODDZzUAQOR2Ku+M3RCXejVcJBrZu/SydfPeJUx+1V3NctbjL
FLrv44HiBnpB3pyOzQ4zOLtwVy1z9vodZjU5pjHo0FIT0UgZ+xXdTqGmESpS6km8
GjguHiib4QX/u0358SYTqMRkGjwTbCCapyp93pw6BZSPMyERK+G/VM08uPGeUtVy
U9ZfroBp9X+qxCRwMSP3pC/+ziLCkBb71cfa7nXVILO5LprcwhYkeBV2Y7TXXEb1
7QThUIgH1k4HOOzu8AEJdpftZ5RycIMrGt69Z07sUkm0zwPJCFqx1spJcKdt3NnZ
nxIVBVYQzT39bhBg9DNaOo6DgTKB9NshCMV/M3XcxUCxjr70CYhJBMLc48n8mTzQ
BnPP+YJ41TnM2KGXMVIMzG9k/vM6fVWcqb5BIP7A47HQtKu4ewquc/87vRu4zMlF
ANDj/K1wN+NrNFeyp0Yw1jKIou2UCxTmbutlKhGCry9jQ3BX87/icXJSfsaoGRaP
wCvhOicwfTApnbrgmpCtPeq8x+EmJ9LaHibbywF0OQDqXiOWcuoi4FYM4V7E5klz
CJedM7aFo9AahEXJTLXu7NLrWf58oiuJoXcWINMVgAeDAjn+ckzoQ8nWy0s39Ghv
Yerr6okttIp57Hibv0aFdHnUuui05oUj7etfDbRxXe5R2SowjgFu3fsHrP2+hhfA
mo0EcKQ9M6mm+U6DcUorgIh/fr3B/G7OVy3EYz5RtMIhqeo0SfMQ1eDCN5NVaK+D
BwuwwTCAorQvPg79ItdZ04Qv12A1LdlevFvk1GLgcDlrFJ3Il22r0D21R/bEs8lr
+pr+XwHlRCqoSVDB4WeSj3wxBauk2uq+BW0d+7ViaMgUf9YFj8JatvDJ/V5mtJXh
ra03HWGE7MkJnWnSHxQCwA4x7O9ROQJqeQ76yBpp1VjZ1O4r1B/ZaG1aAUAAgv6Q
6UxfU+E3xCwKw8cxxmyUVr0t3/l32GWDgQEoVomRk8cbb00H7Pc35JzexKc9ZHIz
pYxSDvselnNrp/23UiWB5URluFulRIsCeoT8U4NMUYDn6AEOn4Tp4XsV4Vbz0IJS
YMooNSOxM8MgR12nYsmxYbi4yCsuHUWNALGx9R0MvKBpCzooXgpKN1c/ox63JfYk
o4KD4so/RBZVobvmK7N17foxeyiR+MHkOatHp/VejWPvsC2Iu+P8P+5tL8PoSEUN
3QVs4O7y/mAXfqQWdDdJRQeuGHFKMDjP5l9NCcZPijiJj1BuRk1XGA6H1Zwv1qtm
kMOU/mgr2OLCQI7MS/SdNeoSGGxPY+CUQA8N3ienyfnhXpQCdBM7+R8tkLFY++qs
vmB1r1ucfdHeHeBxK72dk/FwwU0sVFNFntVhr8/kv2bdZTdUD6ns+U5wxeIhZ4bE
jIDwHG+5Hh8vU/1TLfYEJS/JgkUYgLsBWubAftD78J7FIdqT3ZzOXlAbzhKLMLqt
6ILdbxd7WkAijeVsClZUrg3zgavbL78oetxhTMevo/bNLU2vbaiMzcFvaKW6DAbr
ePenZkTDtM8QvmxdQmoJQx9TLwDbEAbgcDkkAUTlHEoJAMq3NosepLfDRO7qfvsw
Kqsp0uW6dzYKDuXTR+mwDs8LU94E3yXsvxZC0q9Q1TAWmc75halvJ9i8Qmw424jA
7pqwzXRBb3TovokrA6yLmeeZ8FZ/9D5AXiXLIZdm3wNyffJk7n6rWrLo5g83y7Sp
NkzuKtDkkNt38kAColwALgAO8joUbcztPUDNYdaT9h0EGYa3qTwKeAWUpDJSiLUJ
GSiOuqOUD1jpNA5BYURi/gF6wmgvrB8ftuoqsPY+v3dHuIJcfAj4XWKdhvDsdEsb
sMg9hLu4KpiVHxF56EqeP+4HVSk+ZQtNJS4fBc8MGuobHZDoS8MlYO/43nx31hki
KquJ2Ti9vlAM0vUAjlc2rJOsD7CM8IGKJWszfRdujsvax8tpIhxIe6UKugNTiOri
bZl7RHKIXQ40weyZFbeb55LeJreyuHXDEIqZPyuurUOp+W7NYnaHg8+Dlb0x25sT
B7g3f0jQbsvQeEu9+xaa0a6jEcwEBWlexfxV2/JbpgvodcqGzou0bI32t3Xdq6sR
Z7myeuS9HftrmVC/n99HxAD0NYzRAv5myLec44C0YC8d4dDgKIGlWR+oJ70vwB5b
9ynvnn56sNA2YXFokRVhq8cOH4h77B1z1PscAxeJS6OVCnnvf06T8mZzXEyhPhuR
8bl4tMYTXE7r7dJMrOsIpGhKJBpiBdOrRVvSu+9L5oXatFJTMvaMjEGHN6eqnKoW
hHeSqIv2jnkpWug7aCSvOezNb5e5KYpWbbTR/O/zU9toIbBj9qy+sFk5gg2zvY8j
arZh02GQBoATg2JDqNyFEt0B9d+Z4KY1g3wle8Z+8HYUwePUh4AUui+6L8ixIq5c
HgtFX9VzWuBL5SxD9O8XlQiRLD4aExbq4t1ULCo7Y+p9blsW3JlEvq7kf4AuzkP8
RHOUB2fPSuKxD6Uwnshkg5EIAOIpfjrWfD0vXfWVVL7wmLs6FBrojGaw2S73wyQG
Skw+k5U58vn2KmhVql5hbMx+dCYmVUavy4aC6ibMSZGJWCtPoG83Zxr4iGWDXxIF
uJFRUmNeYxpzhZGRMw/Gg+CN1Qj9Vmcq5/CnCXBx+bLOjmoetRh8uKtYulF92uV/
keD2FHRIzo6pPKO0S/uHlz+VQ7cX8nAaKNFxKG9a+TtWsmYbFKAb7x0avbW5lB6M
TYBeZglPz58wKymURC0Ve8t+iESJzgf05WD65uv2BVynbcTzkE3xNhMOhTKbc0gF
NbVnjoq/P/4cq+T9/AD1IBFbNc0Ya9xOdzKqgXNiQ2DcAl6tluP+kaGuL/AimF0Q
iK5a3IavtQ3CG1O8MiDkNvvECuOogZi7ZQeeeThUN6ung1LjNcHqCXjlfj+dffyi
9BPpUgZOa4NlMkUFOomttOJh+NXBrbWe8RouRr1yiqjyetJ4H23ygkBH1CuB1u38
hm5Bvy/ceFwUIeUjmC9OyeyPneV64r79Ydx/I11bvztP1cRT0aIWiDrPGllNVN//
1mvJVj6Ij2B0AakYYwJDREGYYIdKPsQTdfeQVEYqN+bJNdMNxl1wtfn1v9368++1
6uCeg8VzsdLuU+Le9W/ZMcs2pzY1iq31BTBFZfCJ3lKPueIRUbWkujbeZBdF++pf
RrBMhEKXHXVHfiENXQFupqzDXdBdMUvxvKjm+WJ7bPD/l9doynV8KEAbYN/Sk+nF
1j0ricDSpDJDu5qLfHCw48ffa0rI5WVkCT17NSaJYEMTsded6zdM+LTES1gYhkaC
ge1M3ZVyU3e91A36gGbCc3oyySAhRA3mKJZDCFoUt1PU1hH5iuI5uM6ozvRM3rAC
BD2N9joK7O1PmdF4HnYZ5Mx7lUuwnI5n7godhMR+zAymdZ/WyTD3dPi7MHZqlwfR
0nZmyVcyAh+Di90S1yBPkp4kz+f+K/trm2seNAAnD0ZQQOXaQuGy5mPw8aCOuWl9
s0Gc61V7DZZJN0d9tSPNoVWSeSFDrXJAbFXk2NFmcJtK+pmlbYZGVVH0B+aZ/8Fl
80PVs5czC9fFTQzSX/gc2l/5GaJ1Sgn9aVdXc83UK6qIQg364oS207Qj50BPeyQg
TBKBbRuOeVd5zbdSODiePwfiArhwWOXRTFl7UMKZl6TxUf0ZuvNxsUxq32m+YAEY
uEBhA52dyQDXoLEeawZbMFIIgqGx95t/cmDlLfDClAujrVWfwM7Kq1kbG4YajRNU
XkUheBNfxStaZnqG5222jFycmaC6FO9TLmCorhCmqagRJk3iZtdX9VV5dnd4oOfr
OOWI+wBAzlbZtd1mlnon7eDrXmo+Qhhhlm5WxLJC2Z3mMYDnUkDdMbF3+C0I198A
SsiENr6NRZcTvXiMQ8Mu9IgUCQ+S8TLHiq01yhtHKVyggrYUXRL9l6AXF8c3O7wD
A5z3Ydtq0FqJye9sLGKZTIZrolmidKrLKbmiXbI7BQcio0ddhaQrgNd7IKViBcHg
1pLSGYEa6vBJZf4fRie8X3Bxk6+uHj6vFEYqrQSvPXjaEpYruFWubYpzBe11gkjX
AToa2gv+CXwK00BZ2Dul7SLZSWM/LdzTEQy6AlxqzciUzWikbnrfbMUvkEyx172p
6lMEyP+qcjPDH+RtC8367uTuFvVBHti5oVe+WCoil6211FvQArBTeR9He/LTesSC
Tff9Ns6Gsdo5sjBMIViAMatl5XeXeUYaT7mkiFSjen9jZjuf5dvOySxkC+s8AxyF
wFzsAO9r1QdGJ7gnJ+11fCocPtrU9jr8PBwIChZCVGHtt57VPA3AjPgmOeK28ppQ
U2GJ+IPuans0Cey15riLkjct7VIlJ6QwScBrMiyYiOi6Lx8KodZP3ytya1+o8tkh
A1FtVu55F6A41pLSrMdSPun0ZMvKlUaCXjxhNvIykR6sWhE4vFnJHWdCags7KYso
5N4VkdPzbRPql/P1eawkLkdgTx8mVDIV8tj21yrjLIeJMu6D1LZ6bF4pVvvpFP0x
ccJmigJe8+M13xSHsT0tSf0c8sbDACli+FxoPhg3dsB9p936/21dLvlT9Ysj+EUC
T06xpup4DVleUkCI/7+hKpRktHxJnQb4ECNKNdTQDy5639yO3+BgRxSR+nYXw+2Z
hWOMcbPVjPfkZxsYRC1HBts8/B8eZQoG48gLEi5wpM1v72L9FinEICXCK3mupnpu
9YmoMUQ9xTKOqV3vJsIp12txK8W/hpnzlNtPIxlS3+8uvgEqEWVmrHT+xcGYct33
f3INHP0ZSqjCN4U5mjdYeThR3DbDQLY/8om/RdLiBkuL+ESIcNE1gY+09VmWsMhy
lvrGQsGPN4q4JH5lwCJU0zV9yrG6CNTdsb/9DzMh+Nvwu73GnMM1krrU1Z2DAmm+
SqUW0o/ensbf5pIBiqI+z91y33TynxkI1E8DRXb+1JPxTSNaIopPEFYn1cK/+Q66
SxsgugHQb2jRTbqci+0ffSg2hJT27cAz2rQi/QbGVrAsiLWVytlKxEwr8N2lD+87
cODWqGxjvxnAUelCORNRVqy36BipOGK4bxuFM84KO2CUauMP1FHxGz051ovRCutf
v700jwe++SycmuAHN6/2GUDVxzNQ5lIcjCmS4Qg/4u0Xt7r0uxE+DNMpnsJYEzYO
M7XMtdisPXINHM5Mg9nIQMoXN+qELzdC7L6mh9W3tuvh32RypgfUYcwOuFF0SAFO
unrcYKQlAD4txlLe2E5UvkikONZE7tYT4wf/w7kxxtPRLbVxij7BAL0fIQ8aGeWl
hHp6qZ3b/ULEFLl7MfKl0gm6mwd1+eIP7hjJu/VGTfZFGqPsu+37zMS2DRRKi02X
KYtfoAcVBZ7tuGtPmp824TWIs3UDAvlH+Zln4wuCovraT9zMiCuzcO3gh72ZREIb
NoLLtgMWYuKCvJ5XGG99sdQ4KT3cQr3zkDy1iRLnprPZJpfoweU+z2PFgYBoFiik
1UiDE7F8BdPmYvsNdzywGi5yXvaRkMs5GEzd3PLcepzAeHCznP0aNOlE1dGj6Jio
U6LFnFOhIGq030W2ir+AOQ2hi+f+5/CQj9plPj7Vpi6T5aggduDM4/oIYh5PTJ4D
WE36tWjwZpKWmF425N1Id7kYN3J9vSouS0aDaqlCledvFC00bY4576jHJRW/Q52U
tsgRNOgM07j2JE4hOmL3IEq7cvtWF6ON4Lc5wkcHyrxG7c0ohNKoz+fupnKV5pA1
Rp8o4k1Kx8ER/CGaEH6dFI47DAk0qSLpCJZ6VjASBe+ragvYNYlSjxOszs6TAZDx
9nwUXG8i72loOe2Qg8Kp1oPCVgL+aSjz64+hfbdz15O/2Zctg/71uQb3jFpALBRb
mkP6UTRV0rJJSdxjSZCxBvt+3E+94HEnIDAqT43zlnk/+FrCRXZ8IQOU68r6Mip8
WCqbk45sqZWzzcSsiRiFwh3eMx+DdQ1+/z1ehGxFDdjDm+C8GgKVTWrMr1LiBTeb
j8lfYBkshCt32ElAcsLz+t8XZSVZO6N7c3rqYJD3idU1iu4Oq/Ftlue8rhJbHaPH
uJAHIWwkkIFT3k2Z9SoD4b0b6NWn1bm/GTq1GRPfWKOGrjhsymfvB6HuCBIJdYij
/dia7FTM8G78GyitT2kzfYMdzXupoL54Io2jVeNqnBn5VGrkh2gtbHv3W/LtHErV
pRyusIzSZR6dtq0uTyGJBUGPxOFR9bSrMhU+53z9vTfriaoBGkCBpnKyMuR0B/7w
G8UH94ySlQQOnl7Qe0Y92Hfzv65klWbN+o6c3QG9vxZlMT4WKDV+67PM+6GFoKIl
shocZ6Ivm6TFLJn9HV7e3wRm+LxLJfydiJV77fQqa5aB89zoIHiRstQ5JKd9O6XD
2bTC9Jpj+ZExQtbUCxzut9YzdPlQeFADsJ05UzBvmH7zLTmIjiOsZqFliy7twtQH
93xXwxexK/n2FD0bijoVDmNR/1CN5Da7jaPaHEaNubBLu8keHaRfWxu0yT2e0h0d
d4GEVS17DNzc0l/3pG7jsc1IjOLv0RX/VSLCKdzj5ta/QEu5D3mZoKJUsLgudyBy
VWb1kYR3Y9iPLg1PXYTLho9OQYTFvl2uqBRlbUOIsZo/+MQC68269FERo+Lm4yxw
Dxgl8oxnN8FDNgskg6Tjz2kBBRUhzS8KXFKd33uDwLoVvq9dwEdF2oJg8v8Mnfmw
DE4O1EHFL5gLcWmwfhdLJd7s7LWxJ1eFxqk20/0f1C434voBNeR5PQlZ5RtLe7At
zMUzWQRyIo1ZW0afogxSpRd/dxM9JGCmbLcHqxWYcJGR7GVOE6vlsaourKFj7Rb5
n55hLg4JfL3X34teilm8cZy5PEQTg+BQhdGnkCjj2wmQpz3Fye3x+DT7XDFYLLc/
rI9xFEnFVdsgVO4ykZEZb7544tRdf8+afGUaGbgLqs6kjLVT/Snvm7n5mVFX4olD
gt3OTCAujECaAkUxP7zcnX96EeVn0qT6DVPc3qUfpnaQdwPbGqSXUjNJMGnyIoGx
hUpC7/FXWSuC3V/sJ8Gdj+ls/nfd5SZO6s8M8wwNP1F7U3nH9z/ediVtJf+Y1Vmz
IzYvWS59JLcw+LSsvNdWlJD17aESDYhpNyjwnhT6+VQ71IxEqzFNwDEi9U96bPgd
TZyyl0LzLMC0npgJXeDIMdgOTIs//iSlG2vGtlc3XsIlwISs1MXjjs5MWdvfY712
HPwcn1YXaMyWOcjag6yyF9G/cM9ttG85ddjolid7eW09iiPQHITrr1Lfbctr/jb5
qM1bKoqfXC6znasmAfEC53Kzs8Xj7rkrkWIMI04W7mERvAunhenA5MaRn19JwLHu
xab/+tiEuALhYt1E0jXgbfAWxBVABiz+OQu78PZhHq64s4h6PC/aA1k1JrTu4T5e
7TNfP8FaH0D02vrj1kZm50SiTfshB0cBx7bhMFK85xAJ18nS8caEySuH9p61a+Lo
7KpUndEXwLCcfZm6ubT2brni+eSz+lESsWRbr2PMjIIgwDZuj9qLVxV97jY+HDkO
dwzWvpxdbYpYiFJgDjXCLubHsaGHHh7haLs5EBb77pa8NAFCx/tBs7TTTYQhfq1T
5MZlYbwb2n/l86GztH6CU+7b855tJRTqiC5V893HMwq7P8dfMS/NAgVzCXTk+YTT
wbgLKwEo19qZUvTdiSyn4Pb3hudkFXYtYzw5qEyIr2h6kZKGn9MvaNmov7+bydKb
O7mG3NUEjf9Bhj3cHs7Z1ZqWZfzxnOD/FSviFkorglnQzfGoj1L7RhU2r+ojQndS
2Igs8pkG6X2P2w5Q6KSFEiieIqtmRmHfaddb7w8Wl5ppKT/1B5MTUTXZkhefG2he
2tO6fvpsyVE/q2gifXgUAtc0jzA90qdKpjiOdbm8XcrQGUEG/hmYmpytwRK1Jcah
u2lxWCvVF1AeVJxmSWpdrBYoJbZSH2Ik7SXqQjNn95UFJetmyouHGuuXmRjI4WJP
3M2U2lresX8wGNIf8m/pU8XBHz64zbTsciQMFUvXjjmUN1Jor5YZ1xvy83w0DzuA
MLWybJYMk4r/2un7sdfjoM8HG7gDuM0UtPDLPyoI2US7HclggjRiZ8jkCupHOOJo
QdRMUih/piOnswcR4zM/1vyLNB0vCffCfbvcoXtU6285m5S4QgugP9yxbMuB+oGC
cqifrKxGcHg0cyftJTaD+hKOxMfFcM+H0j6OCfF7KKyo2PKEVhxOnvF30Pp4YDzT
UVcRPipNLPNAwu/Nt/b0m4wpA5Snqrkb/IRBN8g9JsZOLSM5bGttS9jvE0+UJk3v
BGW6X1iEc58UfnI5R/APYs+xyiJkgxCFUon8F11Uu0VIlwhjBHAhWVl/tffaEbMA
Fa6Y12+Q89l1nHaT7LYXvaM+LkfqjzzsFzmLjR/sfj4xH56xrOgLMdc1cwAKvz4j
yXgM9CdTo6G/4wWS4inLu8fO+snuWsjqNFpvdbbPM7AKSkrScmZFKUnlEZ+gmlj1
ev34h0YvX8uZVGw4AzSci4JRpnulE72SVMbrrmhJHqHiZxwJ2fdlD3jHJjITWnfG
+jwAe1saLUfKMxzp5/OGjE6uiA+LlFaW8PVVWOf9MVdCjWd3sVkbKdRB2qH+L0oh
xQQp6cK1tGd4vyEolPdwdnZhVsy4PCp7SmE34fj8RgZm9TT2YwyB4qfmvMuvnEja
C6pjlD6oTtn6e02seGIy+hHKNPnPgCRQDo3abSr6Ig+gYhBsQYWLUOckrF6wh4ED
kWMdvx2OURDygknXTgCjJzhNfavJ4NkoZJTpX4nJjIqQY/FmP3zcDtufBNZrIpEP
isrqyNPkDcBswqadaTOqqcjeQyYz8sXWmJrRXt1GxGej3oG56nat4PLt1E3wTZC7
UGTJ+khvlNA1quciA22djMqTEjdY8OSi5D6pWCa3mz+WNpdgGq4i/xOO7RKYcpNC
n8c5+IN3Fn//pRFXNKqFhIIUqAe1qIr8dVY/yQUWYkR6YNeY6j/d+DcTB/RCrLaE
tZgTziOcDd7MbjPuQ7I5oOvqqjAQcPVfOapkhGlaltHUpexFfpOM9IQ6Ia/TXXni
1b7GkwyzCfm3bSwoamGGjKgJUvua8+fSO3Q5t1eAVF0iXoZzz0GcchzuKd1rG2UY
jtxWL3cfP/5qTG2nlnMwyztI8FEe2QJ6fbj+eTZB+h820WuPieHvVEdrpTK5y0uW
na95JVQH9PzuYjvQOwz27QHAhicCTNXZD94+C4O3dJfEQhaSSlZ42W32kR0kY4Wl
lWUs03NBztc9IaHx6IC2ywIxjW5BLUl8TNbPZ8lBIYMCiYClMdGYjud7gU9C1bIw
rEnzOkbEoGPu/KSA+2j1Hp0hsqZLoh/9TQh6b7wMajP8UEDT+/EmpNbp0lVOqkUF
sKd6T6cd8FwhhrEmcecblL2RQJPPs69VkrJJh3xmodGG1jbQ6p/+6emBBlLeuZYI
FFQSnvdkH/g3pcmMGZjLbp7C47j+yX2Z+AvZp58vbFg4E8pXD1PBIDT8O5QFcJND
mVYWqI2o7JErFuTns9m2sOhMl9e+dr/+d9CXF335UxJVKRtl97o0PuNiywr1EKIC
xGUBPfuT9RhT8Yww1hJA8G7u4if/GKX87kd2XBfL/s18A56om+6ssvYa5Cqdq5j3
QKk5iLrUI5ahg2RzifupVjjgCUTmwjHOURf11KBlcy0e5dsOiG3XXSzBYz/4ZwBW
L3Cb9gqUvWClRNzCWCOb/v8xmcwA/0zQX8BLXQTBKoMfEvBpsXofOPocsi1QFaMX
QXQKTh3+y1DsjkSAlimOW6JmM1IcbOZEnJJ1peqL2a0NV9sWI9/NxoOJblBJxuas
zVIg0gA6x3or/umbX0oJABXDFSGU4k6tvAdqL4+7gS4iPMYMsZhX2cnPZevFgTrz
+UztFvSl14jXIPH0WdC2IoNJLHZHjJxf9+B1pBNpDeR9cfsC+ev1a4N138qN37cb
Jg/b5s82Ok3LabggNtIAQAu37hMocxycIrMnK1VcRiVudpq2Vq4p+kfZg/s7XMvf
pZUT9Z87omZQryGBxyeW0plsqmzvWNgBjtCXtKfMqJPAQEShkaFEqf09q7S7pJ3L
j1xsTmK7rLDyCEbRODtMoKoajkrGkUi6X18swlARrc9K0cSx5Q+G6d8VPpPlXFNg
g4pgsDzEFyIm+ahw34zqqx95yX55nlH3oqnzGkcyPq0xHx8GjDwT97axJwNw3RYt
Jda/3LexzBmsDn2Vr3bLDcwMGl0tyyJ64i4CaerN+BGrDidD4iK17OEVpPJ5RhyF
r9rLxmaiD92m3sJGlcDwfq7EsVl5N5sBrdgImXXxMzag6jI+VeXHaM8+/orBrMMJ
bs5yf+nnpOaHSuQAoxKaJlx93K56YDi6o00uOGdvPTLcTO0IWVh6pcfBXFu57mnD
wlhzvs05RS01E8/7+QUSP14uCjjVS64Feb/tmiDlyrwbkmT1GHHMQQV1p9l8R02y
M3VLpLQAGCxOggAEprn4UemsI0kFOK+hUOuSzvghlOJjCQaP2Ti9ZBV5STJAJ7nc
jWovuKywDslfZxKIztYcUVgywL2DixGnXJ3mCzch0+nMsRtuR0ZrDhFAQL73MmKc
Vae08UVlCuHALI/NakwgWF9yY/NwDHUmUkCZwOf8ihQnwb6x5BjnpKgo3jJl36LY
s+MKgWfR8UuPy2MEuThZxfYcahGDdQmR2mkUB9LQn0/QYHsjCZBc1B0UmCjqv7Fw
/6tbaoFlFKs7Vqha/zK2f8nETAdv7fphfzkxSt356rtLlx1v5ZntLbQVWZpW+RT1
g6LZ/1XOWAuIMJZZjF8moyXw50A7tOb7xkCyawM5dsiDC9QeiACCZH7UNM6qW5tC
wq1wVWMIvWvtTz13agnlKgo7pP/4kpk2loWC9u1ZE2da4Gu8mUT8vdEzW5u5ENeh
sNFu432N+9gOdzupmPe1R/TbnyG+3lKevkOfbWQVDMCGtIVidMNh3fj0amYw9MQW
UALHkonPAFXcPR8/TR+iqGbtQN328FGZWC+1eyUUPwqThpbHkc8NAkigXFe0xmVJ
g8AG9QSbitCKua1pmioy3iH4s3sUJuXdckFoE0K1WmE0acRajJeA145WloFFcEEr
TnH1fk3kQmv8G1RZBQeBLK+WMj+w6odY5ZjT6JYSF8P8+nPIonkGt3p0JaatRDSZ
7s12X2yHc53SFDSCdIJb+xmYxDCiwc9Hpfao3XPJ5VJ07rDofEYBX6t9E3HayerW
rhbbx4S5oB9TXiPAIqavM7zETmsNwQLD7Sg0eV2FqFY3+Z9PVmDfDtUCyPjhVqMO
rmf9e1OAs5W+Uuusc9ZlXyMSkeA1D0Epod8NUHLB9XFIuzV/nuUjJrqcuzIGBRlV
8RPLLUgIB0SdakEHTL7v5JIgEsLM70MKcOFIKjsIguWFKGWCqhsATwJo9M8D2+AN
4QA0bDNsg7wUkQdMBnhrpwCidO2Ubk8FgTkprPJl6saVR++gr7+ocvneusr6Rd6H
71PSCOHbB6BdhXm7OjoEBQPq5DeBaZVYTBcr29EeDGvJeymZPLEp45h5Igj3E6pu
2YKIHI6zs7C47bjiOgmqUpEfoZjbby7wZX77j9A2L8kUryeEonf46hvsO80sk5E8
8yVQec//ZDrw1zjcd38r3zFu/rAUzJJZYlzGZT7cxWOIkjYQQrxpZBsE6X+ylF8z
aBdXMHdEUZnLR+GTmWKwrnIT6CJB8x8IotMSI/bSyAUt89Meph3NlPH4O+vyXSFA
5nnzG8yLvZM/l86O1JXK9FKz2dl1NeVSrsLdJU2ORHhXiWIp3nMt5W3b7FTkKOb4
v/cpv2VpbxITTrAlp77UFtDD11VSrxsV5y38i9e/ndde/H0B/1wIfEaIbSPLaXy8
+1boVf4HEhmNiJTxNSYkk+uWAQTXAfuRd6Wv3J+2qFzrQe52niGs71DL/2RXOTht
Vzv2uJPZ4YQMw1mi31kE6+g1f9tUn97rJ01AMp4FB4vKSNSpbvhAYXzvVFMIqLYs
/vKW14a5HDcrq6UMomzV/h0vwTtc/nz87LiE7oH0vFCGWhizdfAmNhSPlwOVvNDl
7A99g57jakI1/aA5Ira9wd41xZseAOVm/iCu4HsNiQDUkSXafkCgMPt/3BK5FBmI
2+mE56knhVPnY3hGEiwSE1vA4j8/iz2jdBcV1yMMB8XSsFn+l6YZl7ZwEDOlM9WR
+nE/pfhGLqYdERKiaauCY7/t17HSsk9DkP3tytCdg+/7805i9P/IkdVsaD03QkMJ
8+jR4hrbvoYVzyFuvhN1llhLSw+s3Kmqy2/pLxQYJhsNTNIkqSBp/gxmVafAVa5o
G6QofeRmeRBlJ8OwWjheG3jFoprapLY6w+pfDhKYd3E6c0NVeugzPwwU+cBsbc8M
5slxoDtPyYNMbUhVbqirnVS4T255PdJZXJK85xu2zRq3pt8ToOyiLdhoWG8v5tdR
+qv85W0UHjzGiI7tFcx5pEh1iW50ae8tKt3/BYlM31Kt12xKMHtqjs0emq/t2hTq
Kb1ZilDwxAfDUd9W4LIq/T/ktwJCqEXeuHFa+ThJ1AFomMbjkhNKxNsJ1mjoaril
STwecm5AkMzN6AssNPB7gwIS0SG+trDKg7drT4rG6vbnhcZG4ZMPrVRxfJvnZooD
1ddPa6q3Q2iseE+eE5YAvk5BcO3uiWu926Dfhp8cavLnffKOBDeHzJ3QLMewuh8S
EVfccqpQ2ZWNMwP4uR3pUx37AKIjmm5lmWD9Db8hOaQQ2oqxpCPraZO9YZbaNVkH
1QvCsoZLNPrnPfZ3kHKqnXXFbpMU1521k9k0nOj6NWMaXxYsxcO7SMMTT4rUXZla
I7e4XU9Nm9eU5theIkXio+lzej/MfAsA7RCpXhkvQZH4Jp1bVZ3OuuqNA9NkVmTy
Ei+YJV+SDmS0/NIgqdmX2a+5nK58+or3/ace+wpD+brNeEX3sE1rF+dnMhMfj+HX
0dzlwUmkVmQaJSd8wRytpRK0705P5pH3lcN37jXqNw8gTJTQNFAxukAKIzEsAk2l
xzqYPTVKXgP5xnM+T47CxrZ6sJ/kz3BQVevcH5pqo25IOhe7UhnD1Kj/zIuPQNMc
O/jQBr+vvzbt2LRqL41+JkZnw5A+APEJqKzKsbq1rTUbWMYfRK4Dhit7t2SUkmMO
lcHEPy2PZMUTn1HDTy1mmgx+FIgvBTloav2Cgt6dtpbQuC6q7jZay5jGazUR4Y7s
w3IM+Ot1sIzkvkf02+uoMuwW2PZl6trVKuGyc6Gn0TXy2p1ZSq6YmQE3MniLG4GH
OBIgq2QEmXVIhcl184ZjpqQolNhfRk6mCRxUUw2oz8JiFa3rPYSYKsSKFd0kr4Sd
Kpo6D9VEU4KvvIgyG6apmwyAN8gwX17U+Cv90665tOvRBe1woQLr3ER3p2ZEelvc
djTxG52hOyUhqsH2pstfkjt827ddIKB/3vYfja0EHo1UJL7VH5ZUUdooltIVEguL
vrgXSBIJKc+P4POS1n1WFn3zDYYCJq1Ytsc7kRuWVldRhi2RS63GcnUHBL635sCd
+H6MzgEKh2t1rZnpeEcDT3khXkFUeAJp1Ykb01/d67QTheW1TIJYwwiiJmtsjy3a
gwsmv69YQgRKNHnq1yB8nOOLYKB/vlmLKIjzwW7dzeO27pP/r/ybhCYBpUaa3P1W
yM0x7kgGdvoWHXcaslE5tSQO0hCy+ENp1vasFAVfKEIDLk8raXg0PT8sZJFfDbrI
QG8vavZtVIUIfjFxGiO1Jo0ifeyQ0dbOqy4ZRq/9to+xTMBwqqNsV03zq693KWu2
wWBcDqoNlHob+D1QWx27R6Eq1S7Gtbfn+auZ4zzf2k3QKpiDB9PjVx3v6sEOTeu+
Jp/K5wRv89TU7Gq5JC8ys5Tz7e7ffsMWFYWitSHAhuNQHj16LOhyX5r4jRS7j+kq
fRUe4M7LZYxBReSiIYxK9FUXiLOY5WdCMns6LQqw6HLYBMJPf0oMNheGYrGKy4tl
NHGNisgVV9TS2gu0BCg+LAGV0WHWTRnp0uvmyJAazXPS7731Y2BvsjmnT9e0MrpW
7GYTi3jk7iQcPWAI7t7T5rt2+jM+MLvSf0nEDooKAf6+ImWHQ2IRiwymfdBkhi2r
gYHPKoxSYNDgvjMvQgKZFFXdhbVgm+1e0Srkuxvv8uM+S9re29A2EZEOIvWsCBfL
tth/mYZGTQ2+hzM8s7wkv03PgsGJRd3LcK5aDz1CWoEZprNBDcAW5A4frs+Y1kPc
ce2BrGJy4L2cYGoI2kv4DuCuKEFYqoWgX7GgzIwYAD+dDR2gw7Zhpc39ZRLUU6La
VxPe6bD5VM1MqpmFZL16QU9i+T7dzIPSYsSKYlIndVydK7hAz/G2/AwNOb9PeBvC
cKcKNsazVyLyAmQyqZ1MVf++Z2QbaYDvUrYXUu/QyHkVjSBn4KpAOznzsh+KDqN6
COtYHXvZ3UySWCDuNqBSOh8sUqcB1UP4onEx9Q8sF6RpM6Oqb6K57SBt7MUlcARG
IT27nOH5oWyC3qEYvkM6FF4D6kE/4wPK8jKjNzMpT3g0zmUl2NWygZFiInsc6Yhj
wEhWGWufQy6KnDK1kzQK4Dk8w7tQlLA5SSGcWiepsfuiLmQld4WuMx9bZ97BXodV
iB3PxYd7tqRHaP9oDms6EibEzki5p7hmtuF/4i4Q9YckHcXDMq/pYL0l8JeirWlu
/Ana/XzFziGYGDaqB1mv4avx6e/jkTONwE3F/VHYx5DcGGyAliudmn5uB5xbvqf7
ptQ1pkAysAb+GpCyuoiYCpRQYsQxEKskSQIXghRTNMPZVUVndVMPb6Vk/QKnRtYa
wewYcqDTjXc3Z9LyLXa8ZfzT5z8ShmgzB86/QdeIxA4Kn1sFHZ4tsDjTlUoYN9eE
CJU+A/PcnkWjt/EpLlrnMOQRzzZC1y0RfhzSMu5I9CcOsHLRg7kUav/E5/i7lDMv
A4tHCEwrXtFaaKQbh3r24ibNvvDfAPo8hCLim88QS4Mo5dXTjMBjoJWGpO8eMtQ9
E5eGLo5TPrqdYbVL+/FaDZVuzk+ThOj/fhTohhscwDyt+4kZjkVVHNp64MunS6yr
lW6MxA3Ft3JvYcJft6v/VytkK74Yd3tv+0ERmu1n5uvsa5NjM+DZRRj+OOtRG7ZS
3trqxgpfAu/FJvyoODUZILviH4V16IyiOdtCW9BMrYvRvJZFRUJi50Re+Mw85NZZ
zpc84u50RDzmBT4t588ddcq9DhwfYMAGaX5zepazZYikK+ZwEeEhNmkf0klCJder
OxxkAqEUqSpOk6PTNMbK+9mcPQeqk3ijwcmhNPrW7FS5Gtt55cIyKtmlJZdjkfuE
fZFojXXSzJflnkuhMoTjHAGR2GGanPIZD6q1+XMngjxiSDkjg31SqiWpI//H5+BX
5gX7K63k8QYzdQDFMnLezCAOfqdvULEAGYGN99W68aDZ4r+b2kAEc0Ls2ERQ9Gms
Oab92vXULgAe4txX3lLf523phFifnE7n7PpRYtOE9e0la/PTAMkVWjCTGpnf8cHS
6F09TKVs3dt+P54UkX5GoIYyWW8fbQgqG09mVHuAD7Akj1t6jUF6GwvRQUmwMNRG
NCsUFWqWe8B5nuNA9stHgwhhJrOqhoZKtL/rCb8549G4f7Clke2vFBMYFBBDHFUy
JFj8U+cEyR+/cSe3LTirVlM1493TSHnSrw3c41OuIboe/400FXmGuxoan8QFaxv0
z9zhLdrTQ+9YgNxgIrgx/BtdkTJHvQbMc+tZgetHBDO4A+OnsxpSooEdaWSnSJbZ
pfvPTDaM+UHASMcWwC6lBt0ZoQIix2psYDpIPRvVyFgKoxpgeL1QZaKlBfpDpJ4s
aBiqyctJ0ZMPmoogOUTDlDXd8QcnvrOsecoiJFJKUDOoDwXW7dXqW1McfmXzW1fx
7rALsTLNrAeSzBQVs1LW7Sz8D4eMUgSCVjheBL8nZsKHy9RqirwVvm72y+Ow8dGe
3LJd2QO1dPrK4njr/Cg6LUju9I6wI8xHVVgLz3q9JQIzb3f4EoEJqI5sr6hBdyrF
TAVYu+Di5qnisFKYxmYdAdn+eoV6q/v7KvzinlIs0iTk1QKTfWXSISnwu8iLpaEQ
/WZSHCY0ag99XNkxUj/I6qlBuaJmJY93CWcIrv39CbU5Udjq2gibhiYv93o9Sa00
ULS9LqQMRayCj6IwaOilrCt3z8nL7OOU0WzmqzV1OAtxztJqpwtcM7jps6TLCjg2
dnpke1ZYI+HHkxhUSvKsSK3Rt1GrQ9L9SW56QtqaOttKcDEJ1HurMx535GckjVEn
y+0Y/nZu6Zk2CvkNBCeJ+sbH8gk7xUn1WEikByEW3XTEiKDnDaY5/FqfpcrdUKLm
ShOB97+hoX2pKSiTesKmwjhiA7XZvzu2R/dEdmWtMUQvZaTd2ZbwybudLemuvdDH
9G458NgHe5dBIGYYxAXVg2TSfuywKILPsG4aqxU90nbYAEe2dTQOoMZNU3QDdxGG
v+TvVGK8CaEQr/XQ954V4QrmS90up+X+O0EinJJcecgP4p9+fWNBQGZ0x4jahImS
z2Hd2uulBa3cc18cbbhV0DySEjHMKOIY/4EPo3H8QO+fKWIngNxvKoD1zw7yB51b
cNuhvx0do65/AAkoTgIzrypmfCt/5vKqGLcKR9DNPAEaArjtBCD/bMIUwCCqYhp6
yEBld/a9E6pa6HD3vLKPvRb03NqX1yZEnjpc2w2FTnK2Vk8+Q2dU1yGDa9UX2uYl
DNZMEqK/b3sSU4R/7qbET8+UFjQpI3sU2Dopbw2bXg8tSNrhE18ig2itcliHMO8H
Y+bwyAUF6c79wz7XEhoP8AR/oDz1Vh8cEMtZnil/oqZA0ekmjygyfg/aGEQOsjU8
ZRiE3fJAbssiWLQYxwjaPxTdHH0X1P5wIAmrijVsgrRWeBzntM5fYe3d0hb6fcaK
QuiUS47swLSNa1H4C/dAJ8zgdCV4PwaaLJvK0+PVG/jAvex980La7Q7Gl3bSa8oN
WxhMCdp/mrF17Mdk85Hr8YfhiUVvOQGF5b2h4JcHLt8DA0uwc6h5MmbPYV62yfIU
hy9GxQYeXUw7WrCT0M8kXazQce1TNacIJUY9QwxgAZklV+ixz0ezk356WHf75gZ8
9dkAjKQKck/vgtcJXy85lrSfvmBoPFSF1NhIT6D3cJ7Ue3UVUP2XbvO8Ru9WGmp0
wJgRQfn/IkdHoxbti0GDO7mHWJJL7CWX+Gdo9xa/3hUljO+b2NMmY3UvkaS0rAit
TpCLacsTk58nqFX+kqgEXp8atV4U4aDQ/tRkhoseJETgCEmaQmJbTjao4dp+MIYG
7OHJk5kfrAmMysJ6AbHLsMnTMfwitVrCUC1xyLKF9gYLu6i7H4/dAcFIaGHEL3jZ
VawKLDmPhr01Gvqdafq5GKRg3MZ5zocwy6UbIW+SREpBPNWkH81zTvfN58D0epBV
j2fZwgwLO4hyYdbhp7nn0pBYe6qjquOc8pk5E431x9n7VrQ4bp2dbE+GRXZX696L
yx6EOkRDuCDUx/QQKnfqOicJk/PGixmSKqcS6EuRJSm5dru9M0ZjmQ+9k+n0oet6
Z4KykLQywg1msElV00OXgcqX+JSw9NngxGVN4Od+9+iYbWzrmd4VovdeEV3op/MU
Gei5q5Rtu+aFWKLQcFpRh+6+RF1cnH89j1zyFl2Epkpz1n8mb3MdunQ+pVBsPgkk
k2M6uUml1puFtptT/LFlxS2V1J0sML1uwqjPXEZgI4G/J7MKTEVFnM4OHmz2ncNj
4SL8x7eNu8Qqe1B7NcH7+p0g2KioQCUIh284Q9y5EY7xnV7Pffgxsyl8P5Lk4qZR
5PI52PRBElfAPZ9kPzcfWK4FK3ggB+IBw5KApUKiVS4TXBMhXg7AMW8w3kVw2JN4
XT8vpBdWesH49KRH31lNNDXeKY+LA+R2K1qoUdDHsjWl51GLUwGc+7CykTRtiwL/
D9sLWOs/nl3lTVmA+d4fhujDIch+GlTdFgRyDuitrypdAsc/KRQArQNLAzxiL2j8
lwBwtNQf7wofC9LDIP4qQvN7p2is+YtSr6XFAqLjiKc7graRqMVfArtadaRxxg98
uKTgLCNILN1Zy4wdvyPqX0A7ldQjs3bX+zrIbqPd/573bvLDBPDVRvieD9+SvS7J
DnRDQyMg2YGJUEMKCEuNgsRzDu+ZnilxGzW+pVJU/3X1opsLB2IPg3bKYREoukdv
phak00OH5S2t7etuVgBH4GMcrajpajVmhP7Rs2sov/aWd0GGcjURZbIgMr+9/tue
RLNnZEWPuuNsXpM2+VEFhXpvJm11nt94Srgm6PoasrMrE37GfbINWci02VUzehea
0+unVlRi3N6nArteQ4E2OwU99EzXEcj+/jb+biz/dP6LndsU6ugZmg3C9Qoo6BhK
D/d/AL7vT3vMMdZevhZziclMhQaP0pJvmDxrRrc23gkmgI9HsqMQfv39S+lwIX1O
r2JxbYxODngAnEYfqT8Axj9qpI2hmIdjdKLN3G+PVQEElJ/6EfM74WdKEa67F6Zd
uBaUwvAHpKJLfQpr8XpWgLacHtxijI1zT6yVGXoyKCgFRnoaXka4NVYL67C+7Afj
CAC6U6PwuFyWT+kEa4ijOq+wshvF8W6ErJvLXHiOGe2RmIgoOoobojecOdM97I04
0ILFlkdDmtZa58EFPAwBDjRNHeR1Myd8iYcosjgqQ/oENy16KcZaRsyUUBAdlv3Q
u4I65xL6Nqt2Miyn6HaYDsj9yTQsgfVdkzeE5NP7x69BMYn38R6BBL3crSP/EDsd
uPAE2160ZclPGpzkfbYek+mEUpLu1lK1JXCCxwEU+Ufgc1k+bBxpfds6L6Okf+Ok
JHvxEubduziozIpmbkwDy4oqb3zX5dPasxEGZ1DaDoEHlKFpyRff+2lkYV6nKRvQ
X62b/2y6b7Pacq4ItOeV89yC5Gjk15/zQRoJ3gg8tOSD9gGqpKvovtTi0AuMwEw3
wmt/FSzczyQGIrnJMmzwxF3XRZxspSeCZZNtWepT8O11QCfkzNIn6rSPs1uXKda0
KbZbG2ZMxvuob1bJUYh5yjrsQ65EhNdEywNm/cuza3guyoUhvbsybL6cL7KXupFB
MaFMott3F5KIVcoCI3M25uLqED/N5K4H2HVEJoLtQCNzScciJIysASaQWDrlaeWQ
F0xXw/oBWvikNYZVtcbDpg/uLhqthzAYabmra49uYxdCrNxvlGWXTg34H9xuzygL
j6Or95nUemVZV0tpQbX/idHG0b9KHXlH7gJbkhFezNYiKp3sD7WUFbElEyz7hlp8
IbKPMym9wLbCU7FORVMHwxRhzyvFe1pO5QKvrmY1am2ymoBXq4VEljqolqFsuMTc
ChV9uFRjTyf22fCvEbQt3pvZHggeXGn1s2Zc4rmahKbIScnCZudywB2YZzzfskQA
DtSyVC23aBgcZ6hDS1KBVS3EvzlqgjHvci+ThcHlVfQNlFHYyk+WEH8Hs9ZQxi/x
HSIFzlH6RHOsrKwU5tlGacwcfiFT2jSg2/QOu/F7+GwrbthYWGmYPLJJoT6rmLQY
uRBvdh8ysONsKdUoe6gN8JR5k7zsIkGIAbFKOJ2y/F6tnr8gFEGw8BoUgDKxNF2b
zsi5Ch3sqnHBy3/b48ooMrEv63k3vzwmJOcIisCfTg7oX83v4+uZyR7ANulHFCj5
CwCxidtgNVwuf4ma9DS6R3wV/DfKI8IkVVV8dugFyKRNRIwYD0thXRqudh0henrz
9xhxpFRICqMfCFYrNxXz+I3tbF56iJq/JVFZiTdEeGSYA9oCqNyYU8XJeo7iFYeV
60o/c7/wkQrSSzOuzp2wW4IAk/oatlpHzYQbwusPRHeVUmlpL9GuoiL7SKlCYf54
CDTVtKroMv0rC2yzGEZVvbHgkv+2ZFZR4Ywhrt3sotZrsB29iH2wdejnKa5+fLOp
BiAQOpx7Apax4GTH1oBD25Jkfq93iHAJRUEtoWyimB5lERip3U97d9+yvjvSbvvj
9n+I+MRehbdNRoZTURVCbWzAeMkTxjo/vC4THMUogOA/rkeCEtRNjU//oPDaKved
nxK6uD5Ff7XMgIs3+ioQ5276oeHGG1UnIrr/k6QrK71eMfpYSfQtQ2L0Suud5EF7
dkeHhXCJ4Ec2Dc3RGahVz8OzIG2/tLtbcXBWGtgQxTIMUcictbWf0mLs3BmXUCbT
IO8IBu02waT0boi5Wn4A2EdJ/zItgnfloo3lu5q8m2PLs7b2PZ8VPhYkkshLghbf
opc3K7RwmBbRNnfZlJ9GOphLWsvx9ZmZbpVjgPXmmQTC0MkZmlusNS6DLQKqkqv7
m8lLaAc5MD8BAU7TFJ84vfhv1BttEauku6HCTdOT75mHF6AljLivYTs5WxTsAJaV
Oy/d+9gdeeC1L3svAwA8oX0YXcpe7TtcVKQ4sRk8VsBaDP3fcYy3bFEYJPJDoRJg
nS1i/L0iAf19ZmlLT3RpRlv+nxqzgBz2oLVC9QP66dfP1a2MdOdmg5OkSTIF2hGU
0jV+wHkby7WVCnpXK8XClq/5Z55OnUUGE6k3wGF7nJSZC6TWFH/AWOyy2KYzpXZ7
htLMZM9rppUwKsw5XZtV3egwOU0uc2SyZJ/d7xIrxh6gmMxw5LmUv8RWhJz4n1hD
aHa3/Lf7bwV8O3Vu3oFxmA4W7ITpcqg7dbdYXPglsmaHF9SNMjZvTTyBs9PpeDYK
2wy2dS+i9Ty+d7ESR00ebXVicIJctRcuFQSBJhfkrpARjsZGUk1j0rcWZL0rkCsT
IHehinMfw9osFQImjCF1ihUmNpvsVw+w0MKYT0WfAVcwJDpnln1VIU2lmSf0lChR
kalYLjPQday50BDTp5bSJjJCdLTGKX9CuhLqTJEJi+aYCr87uim6iKfP1PQEH3W0
DxDDxn9c2S9drscjK4cXW/enKU3s1/q2xsW87Uk2BYw/Olj7mGGPqKQV8gRohzG5
EsvDyPNf3UVyXmYi5w/GQrMp2w7cSW5ZvZ/sAO+1DebJaFxhIxo+sxyD6wdrr23c
K+7Ic7Q3EmdfmIoZJRhp6cO6LcLfG4URFSkhWrU7tdaLCjQfHZLr1n9EJMbx8mQQ
SmgFtEmFEPV0NOruwdg/3YRumv4g4NqCTci8j2j8Uo17S2t/k++PNExtCRvrEBTe
UqONVCEjPcGDwF47ksf4poJ+/FPnGT/D8sQpPx2Cm6Y9UrpZ5mCpc2nZl38mHGbi
zpMouDTiDLG3Y8BWbaI+q6+6tBX17w8mBOgBEQZSYHNYeBdniQG7u2GKTQnh6ugz
XnfLrrYhZxNPgXGhgOlUMJ73zuFlmwYysh5UgYvQ9LRfyfJmCEy6FbvC3xSr0qqx
CNksKTEMie4SGNmmU9RbolBmQ+cWaEhYBwW/EZQpWCESyyVAVZm+zqLbHmYfkqQC
Iax5YYKIOmzug/rWsuCccX+Ck0d6Ev3GMBl9ATpPLpSlVpvUK/SfBf9158tuHGCL
YEKsVIbJLWcffxevLLUYaBEes/zTvqFW7PN1QZNkuEG/QVzg2Tzfnu2EFjdDamxZ
sOKJlot5yjMokWnwXRIcCUWqRiZV/YHvLnu/ohNPmr0QEqaGkC5+K4zkiWXZm+EZ
GDoKu1j3f9YeepkpCdQ4r8GK5lXEmzS+T8SafCsb6gXG7PICPNP8yiT3qjPn+1kz
v71j8lM9X0SxiKuFSLRp6aXmckkJiq1HBLNY7JUxaqDNgSNj1yIaw3IA/TI9Og1O
mY2A8/lNs9mUb3ZUuEmTUGW88/wxd+taTahqoA2rG+SynaklAZUabO81UyAdFjQj
J9CpXQIdEZty9UmMwQJu3JqE3oAbwvWLI+rx7mWToFXsCd4RoYnqrJ7FjkWs4Dhb
xCm2UnZw/2UH6YeieVW9rO99sf+cJmpYqOCR/z1cxprOdiwT+T/mQN8ahnsOqc+q
ufHYK5lEvuu0YClaaBKUST5Og26L0aaG7bQeYej8RZKDKiAP8kyJRNImq1LA/wmx
8Cdrs14cjy3LMOW5EffYLvSp046qKorWaBhqRtCtqETfa4Bdx3qvNENzHJPsBeCB
M+0PvfipnoMY7IpLK3uNillq0aS6pnVtFkn00TFErc35dwi0wJdsUu9CsaGdIr2T
LSX1hWyk8So+Beavs7tFsg6oNKHZk+dQ/0+zkJeWssDBUbSH3yFqh1HKDMmIcqJY
FIZ52Ent8jI00xUraSX0k4P5o7unufAPH11wAAg9NOR2YTer+gO+HJnMYfe5WaLJ
RkS/4jdLJJQFqysCD/kDVQ4HNN0RD7Jqk05jZDh5dg8SCJsB2K5AH462DrVa0c7N
uPcSjrNGAISSRvVdELyD3LdA2l2meqzp47/PYshoyJ8yD1zk6BR4r6btISOiSdro
0OBnnS0YhdOhY252bJcfvWQPD6uJ5Q8u44lkcp3enssbN2nx5pkzIELdjv0Q0ynS
hhYAA9rm19ErRClHdnpAPjG2UqW32Jynbvp2CUuX0p+RdZoEZVbDYSItuTqhZ2yx
DGzH/kbQBcMCGWM6a+txHKq1LkrMVc4THLbWQw+uueNVXdcbPg6Tt2d0Hlp42VBI
IABlNm50c9Xze3uiHHGbRzbJwy7heKJgJ0KIWbAQUJA+d9oE1hcU6Jyk8Fg61vC6
gbAh0S92qQPSs82GRvDVasUqZ9+5MCkpHwW0E9Nhz4GYmDq68wrGC6Y2BOizxY6E
h7cQNqiaG0LRfW+6JV1bZ6QuiG4gPfZVllq1kCWavxt64jZQ6ypme5vq92JO8Xxv
bovuTx4lJNEoJtK3HwppkI89AD0gvPTfHjYPNZ9a7irjFzZLHbqXpU+cDszb0962
wb7d1StoO8nStkHmWjRZ7NOttCZQXyck1ZqzNpIWafDcm+dOo+GobR/PD+Od6wPt
pjmcJcbRkIGaThG5YTyAwVreITdkvS3M61xD0TZni2N6yJiLFo70tyCWqtMrYLaf
KUhV5LG8LCrxQT6Rp0cijS0JdOaMg3hJyfb/ZM2SVtZMKxjyiHT3ZNrRlnGz/0Ez
waiblpO55J1KR9iZO/qdk0LTz3m7f+ech5jddO8uZ2Z8hdpJiDs5PknBRDpN7zBQ
Gcu+jPqqUkmMczMa1meTEX9//8K8GnUdlVBk64RYOUUV3dTek9U+u2jaEiy3xwKC
Xq41aT6Z/F5jJE4y7qQEvpwdI+Vpoo36WZ0m2ouB+nNjn+DDUfoIHfJ+I7oG2Lbo
kQBHQDHKKG5FpgNfry/LDhY3HRCS7ZpGumX1qItwvXJ5LQChoYQSHdwdct16UxeC
mdi1RO+jN/L8b0TD+DBdNmosPdYt50xbLqLqmG5DUhXJ6X4L7d4jbJX4kmjCvJSw
LGdg0PSfFKRQWAHyaRLE9yNJ7sHDPezHnTY8fIXSODFRZsY300GEODIkHREncyCm
zjWITvV39yR4GXnQ4De3L6nJF/EIwAzWRuUn8PEB1uuRJAQT7X+UCd4CV34CbUOH
FOGRWFGLZH5FRQ4fa+yzpDbLK7zm1PJXXNuKX+ykV7IVe8RpXTuwNVc/W+rqx9RE
2SG+nVfehlw9fyxkXohz9sEfxNVTg581ooOX1uht9+z4jQuzYs83BcgLGjw0atqn
Cekrlv+Xzydj3ZO+uKmCD7gZqVKeIw7RTWrXqvqKYY2TQeyWCeQ5O0ftuyLGa1ju
qXzKqRMt4GdDoKKpA9b8WuU7sxubLe6Os/eBMN+9vanHySnw56RY/aAslJmwAZmj
3sXoFGaStadpUWa9m6jA+Ds9xT24WHAuTZr87kSfRCMy5hG5uhU4/W2v7GXVNrtg
qJwhnQQueKGlqUz5ichnAq+BLbCGLgFZJAx8wHVAkDMdgFpR8wsCCO2UlThFGTuu
fs1G4q8RiQa+4B9KpVxu2ceBWBT00MDinKZbUoDpexzR597s5Ljw/TqX3qRBPO98
RlWwvvT7TLOeAUWbsQlgeD5KSxO5ciFkZhicn8LdurPuHsPcSzzSyyZXapizgV/Z
KEIxwFHUt3a2YU8rhAopPhSl77J7LIEVaZzuDjPEE6hnreyGHjXG0fPzTfHsAR6M
MUMRxpHl9tILucZq6XxLn/ZXwnfC11fCHI5T0rJuuwS0VmUq+qcrRfuudVuuQ5rF
NNbsMMl1Yd1EGeadwRoMjePrJYbDC+dvRDrHZZ1FZ6b3Q874eyyTRVGCmNabNrd1
Gc7d0ee+lzjwh05nyFmUQyD4hK1g7wMM6MAYuO4/YT/WqTuJP8C0zm4A+7vLMpSm
yEFejgzI/BNKthlveI3jFE2/UuQk1BklwyxczVVm/7uTUL7y0TcWS7Xr3bbrFJRT
JhJ6pfYsRzYqN/w1wOv5Z4Z+nSo5UgRIe0fqT+vilMijj65drH9TVu0XTW8vOg09
BoaCSDUo/0KKBcXkscrKLm8z50fQ40n6UbTK17ChjWo3hqkChlhB5zmIjpSETXt3
JyydR5THO9wbF9+6eIaZoIRpO3PJbvuZmZbJ6YZ97Quhwxfp48JCpXIMKJ8WAqiK
6vu9NGkYpoos1+KfDeYxf2WR+Y6b713FaT3hIhuprV9t6eL7soGrbd5nR9dC2S0x
uNMyn+wXoUvuxMl5Q9C4THZL7EZA4hmU/i1/ZkYpjk5Yj5cISXnLqCI3+rtUPzix
8ovxF8p4qrtI5yr3uvBi3JlL+3XVm0d2CnG0hqO1q9F2p6zVr1BGtl6ayGVSv2e8
HBGrnLRxKWJVvLJl/ZSmyB6XGWkXQWZPqgw6LDctwPXqEIGx0dgzdWFsCNIptFeW
stj1lbw0iFhrH5R9V1gMdKMQNLMZcqSK7p9x6J2B9BzlA0KrfsPePp00xePEZckM
66tZgDh/9gq4/mDwG7q94YA0jgYjHNhTOkjg9jyamepQ32iohHBomlxcsjcSYhrB
nH0Wz5kx/Q7K5oYJUOK7GjEDSf57LwTfZb9/EzsQFfHCOggxnZW2h7WXYxzput0n
KYRxFVbZ32petM1yNq0573g+AGjwGwM8zCEWt+pVmK3I1FOgqcWVzMh7JXKnu1Rp
qkUsv+Nt34clcDKwru/UE3jDUf9hUCru8dNxbOZWxKqbnedpLnz1jmEL2F/GKCXD
5TeZcEUruk95P96yzVbii0HbaDfV+5EvBjax83VwH/1liL8j/hUxgH1QPspM9jes
BKIotd5yO7JWWcTm+xKj3EcwWtF5e1/dr2YBf0T8gADy7hNZmYop4yl281sJAaON
4EaR0JjKH6rIpsUK5+I1jPNRebTt5y2jEYQSNEXtnbg7X4EaJpuXl8pjLMAhNKnY
otUXKp80KMYuCDb64jcOpJzKoJ6JEoXw457fHkJS8DfbuM6MpnTEPp43wz6VAi+v
heiJ+uCF4u5QXCYB2R28LsprXF6eCKd08wKbN/MN8r5LKu7etlYBoXkp8nEqXcyl
uUIP05Hqai9w+AXf4lpwEj18wIK7F0P6WHZp4o01wbvu83BwVaPoOYtPsevPpSeJ
v08B6nrpZuzk5G3xfU3oDcS29Ut8u/dMJVEXu5GcoTaiBMJ5beTzc40w+tnIw/Db
5UhopOUCfRC/dgLJQX9ko7fKKlGtA3lx3vIZMOo/cBo88Kwiy3fTCcUycreuIKWc
nLiEH8QMDKuhuHDTo/3WtgsqUvJw1KR+fH8JSVRsSE8A5M/hJZEN5LfMfgwMTmxA
Tuv/7N3K3OFMndZy45ScFGYWPs+A3If842235kJ0Pq1Jgw7NL31g098WlIsUBtGd
ALJPq+s2f9DH3s7zVkjFeH5Jxa+xTD3MXvGDdSQEvTaTRAhQAdyHiQ27IM2MZ9TR
4gIZyeOlLV/MMjcGarRoju5yhrv1Tvst2ckO0x5dPIogQyVxW9ucfwEReZZcv6nQ
d0SQ2Sv0RLHTqH4atF4MSV/dHVaqmK+rLdhAoe5ZwO+mX6atc+AjllQhr6ISPwTR
xm/RCCMG6ZoCSEzkMIjanlAub4mIOxpAOlf4H84gGO4bCxaf1JI+1JWpH8URFCDb
9okyy3M6GWaydPyG4mzMNtqOnsPH52gotMsG5/ySM8LBdYAlalMBKDBNXnlqTeds
Pw7bv4xwFSwoKAEtrvq94WFxYszyjtRZ5YQickWJbf26LG5lDyb4CWZfkJMzRdT9
EFU+YIPLbI3R08tYl7qszn/l7ggvoDC94/i2LF0CnI7NgG3eY1Pf0SKhc9XhWu0I
Hy+tzasDtEaFiWYPBSxfnLuCEIFpqd0HqnaIPiCLdtjiV4qyg02x8qDSZFRVIPQH
QCsYdZMW3Q3gD818Rxd1qLUD/s7QyoTf0hDyPrhj2UiJYbc+jaEonrAh39IEK2i4
4i6rZ6i/KOUmglcMLQXY6lmqTRUf1YRCuAAnhr2ryvt2ICxrcX8dEMk+Q5Lmn/Cu
GyOof44phe/7A++j0AccPe+fThsFlyHxxntF+iqe0zqcu3Tb+jNq7EDKQa3mtRhf
fmaVHQFgWze3dV/kQj5qf08o51p/dBiDso4SYVLZIPhQ9I+mWpdCdbGwcPqpxEmg
UMQTyznEBvUwgZxnxlMD4JE+2xMRT0RsV72GD7RIW5HwfCmz+FcKaPo4lK3UJu2d
EYTiU7Ac2grMRxrrk//eFcS+HDGwWqqG8tBFM4f86Gyo8wWnNW/6CibZpfSRLkUE
aK9eG0rHqq82YHNXtDH8/quzazobZBt6jVlhaMM5vnxNYMKi8lr5nLnsV49DxIix
PTLzHgTBCdSAq04m2iFgqj7pPUV2j6E0RQAeV9PA7HtmblVQR8FuHx+9dPKQS6KX
VP4gmsg2fWc1mJKdAM1vG4nkXrg/rS4h853bgC/IEIBmHD/AnxnJoTSABDAEHXRn
kMNbltCp7ix+QKf2wEyFSyhmEMXnz0+6DQ4mePgPuxoXKjw3xdoCOzAw8AFff8dy
QYhbKu/mP4u6dH9ydjm44ujB/0QSSYUhRZ/3tmR4BNz+HSCukXGKemrxrEWnorCo
HbbwhT24tXQ4ng3Le7AN0aq/F8MHYJDspmfnoC9rsImpJMHFbUZ0tTqwzq1qFIpp
7rcpV3hHD6B6ydpHhDb9d3do0uh2VXk6u9xzVNUD4Uq5UJhBHn4tfPXYUz+P6DQF
FdWF5FGB9Zhovc2hChJ20fvFdy4ROGTm+sJiGm/mYZxlSpO//MNfjudzuXq/YnwG
ELDFPuEK9LPr7LTHx+In/MrAD4xLrkOuTHtS5du1LlTdgm5T+USkB+GqtV52Hhsu
coYC80QILxVqIEiBJoG2qE+OLga8F+Ss8buDK5OhuBlKDhVlv5s+ynWUxO1QGgR2
zDF2gpbOGellZAiXwybdxlbAV0BeoGZ4MvfLgpICpLUgaqmLR9LOsXA4Na6uGLen
KflYILpjYBaB+uIHhLqM+QUgBnFALXsoyDb5YDu6DKFLmhHOmI1qUsHJfILqMYix
lpT9dN0NaK4fiKA1fVFDf326PumbVFUkCPhmpJtLhqGdzZ+LgbtKk+6AlbiUpius
WBnpXjot5Ydn43LC7/TnHEzRSPAZd9rJPh9V+k8wcBUrhHb91X4VLRf7O5bICWkb
oGdmL2Jy5XJmqJkrSD1f6knMFXnGj6WB1TKC9qCHZDRy69XA/Dqpy9WOM/AEcKxy
SZPees7ibs0etQ9Rt8jo6KCfVkfFEBGCLW6mzBEbqrQ7RNgNkfF7V0Ma9P0UFCul
l4fADFceq4u1zKl4VbNzZTITWx7NNSOCF7dhWdnwLdzeU9EJRCYQHa5pLmVknN0Q
Bti7nVjR8MThlT4/1so98ZCh29e65Vm5XLWCSTgVSgQAaColNlcJ25HuIestei3S
bJAZYAjtTHvaOUHoWYKMKLL/HBs3C9zNzlL/WzMU4vo7oK/5wOSQmrO30a/GQcjD
kYZR1YAiGy2Iabb2PZiok+ZAjZ8M09IG95s3wEdyto0HOj2tzSKIK9cRB3l0qZbQ
5+/Y4PFUd8393Si6VhLr6poAaxbI6KWHRTPfCq76fZsr9zT7OFLxIXL6cqJphs2q
gH+dQvC8JAGPcO1dC8NkSz2XHdZP0dodmYu5+qMURyijMEjbzLTUBw3BIlRou9Ty
9gN/XVYFT8TVfTWpRGsBF+/gJPJIV+ITgCqye25mPrF1sX654GeT4eWUu76P29vT
jUdVMJZYjaH46BfxLNGrzIalfZ7ziIX3QVV3RvLOhS3RFGqoaQWe19qOSLPhfidi
1lpH+akd/q1JmUIr3KKdunUyO/X/UMjf1D75WdzM0f565VAqNvyPmhcRSymwxao0
LEP3xjXyavBhSscMIB7wEDrWodPkaUzZjWh1jT9x0sblIlotQEVzsqN/eBGbKO22
CrmhZx4HCAdvQblkCaNObArWlvfI2SZrhzPQi4V4Zzk68Vcb3dPaukiKbdvnUmsm
hDJ2JfgMJEqUBhb+Sj6zOC0LXVaIwpn5kNr4teRzIWRJEXng1W816uVqaSsezq7T
V7/AIE2eEQnCWO4kc/eXIFmURIbJmpN2/mnxpi3iIxT0dMfIn7tZwbbvcQtjgWeH
s3lVAJ9x+qpr00ajZHs4q2ezzEHjCCOlmE03P4uKjV2nqxGjFSsUJRs8CSqK2fpi
O2B/vDwOT7GMO6IOKY3f23CiX+VBIUkOcDvRAhJvyiJLdXkL4QGW8ayVI5NdTHyP
PC4e5iUl4qNPgUPxldSHGGNaqAIH5IatqWV2fB/xrdmqgDWL+203gzOSYNHS3zdl
5lyBfhmir8iuBv7XDWvZapUzaitJWZLkJBgZZuRTFnuKU0vbCtzdu9q2Zcl05n7T
JMq3LmV2ReVrUisrJbS/fVf3iLxGxlN4gpDPg6Gyt8X8lnczQzcl3d4+cjiZJJpf
Ri7dRd05ni7RcvKBAQ50uja7naUE68E+99Qliuz0W6zH4tKHcNaas7n7C1nm/ENg
NtbQ0Ho9P1TAEceEAz4eWjyuXncrxBdb6kLLzJx1rOTJjV8OFTuuwIaPpgshqNyz
DHO/+oTqySuXw+paXC2nqZbzAP2L3EYY+kjKjvucbSdXX52DqWfgjDkHsfXdXn3q
CLiaKuM0Q4X2gvtWFoKIMJTAJ2BFcrHB1fhaDGCUSuUTzDWQjYMPRP7Ynb6RmVTA
LE+rAPRVXhYlB8kk+l7tUNm8fYR4xGXUQAX+X0xe0asNVVzg5vsOFvj/AL/0MC/G
bFClRCDh3wR6ZmAXZMEaMoQ5I3fMDC7s7qcHcb5rB/uPTtd02SL/ippI3gtHWfzd
jVQwlrWQTJTvtsvQ9Cf/20hMJKO8LHcPWpkVYyU7foM5kEkVx9atnPafU6818SDu
nzYPZLgoZTIoSlk0xDuiaMcHPS8vYFVLEz9ufdRn9+djFmaFaf1mLxxKaT93OiR9
QFgZNy/tyNP6VbkbzY7Dhz8EqZEWNDWJOJOrJU24ax5WfraVi4FSjzWs0Qa+kMcZ
7jYYAE1EkldFpoHeAiFLRhlUt5pvSCT9LXDgRiRck/4zmU5D1QeBwjvai+8GacOF
C4RRhkg3Y0ccXb437vFlVd3QIzQNbrkQFpkkXcvoqokacszmuuzEe3WbDgaL5yJP
T48HaKbjE9isupsMgS4tB5FPJ90/mKFIaJFt/AiMDHXYNAMT9WaM5xaxc7FaKz4J
gIIWFoPvFhUe30leIB8fjqry5bJJi8dLdVP07EAkcsYTzwA6exXGSY6J/hcnMIiR
ume4mLycLdIWqvA7E0/mG5RsrgpixUlt6iVUNv8L972VHqsxz4tDwA0SytKWwJO3
tjh2nVhXa+N4hCzVKSr8t7niYj5P3Zu977286DX0yOj+d1SoE0WGsygWx4kazaWs
Qawg9w9iARILZcDB7hG1x0TTKPrgbGWEZz+VOxhBF8nSBDXtrMCcDDEejBaiXXXR
NIabiR+HGVctG9uDBC+BkBqf77LP06uYUnZRL7buUVWU1/QvvNuRR6WvWGUG5vvX
LPnnczllfS8WZy4T+urTUFSPoLddjoN954AwXKHwF0uecL3Ey3PCX3q5apdNBo82
/kh5/7akHUd9ly7ql1WM/L+5ykX5GdxYALUJiY1ASe/h7VXebm7CKznKGL03b85F
kKmmfbfJIDSvF4Jb7GYEJMbqEVhSq4ubjSXEIW9ULMmkWkY0xf+I+2XD1tMatZCv
oXqo3q+nX9xT9yL56HyexCxGXqVtrLmATvOWh/I32vCOW+HT+gsf+YbkgeEhz02r
W2o0nT5cxQiZMRplXHRC50i6RtD8trIXVHuQ8OzNw7nBup/G26ZTP0QX0YO6zC3e
wbJLmLKS44W4l9zsCZlLfq2HKYSpoK6DARwxL77UMr8XDAtkWrqS8nhRJo188wHM
ek9M9AhGDtHQoKKNYeiOxCHzv8wP19v6SXPvlCTAi3RFm9PxFEGaYTzMN/5gjMp7
rWoyToV1sUpWBOlp3qXfsmPZG44qfUn2wQ6VszMMYCGLjlF3m4pE1mDlgdCzonkY
kEVb8Z75BXJj35qwObgMsi1YHwHyIUEv34gBoO+QzYDtcQI7imzUcdX/aH9GLEBE
cmyuHCq0MjjzFtqibIvd8khjSAY4QSvyvUQrytfh6i8X6DK32Xh1rto33PArMK0v
0UEubQNB8vs1e3Lw7IHscdz1lRIWlUF3PzwyBTQcNGqViaFnDxyY6CG/J5vFp8rb
8GImgzmL+gG1+A/kC+IfFT7Zf8MbrYfIYkTGN6N1pZVGfggcgqwYFbmYyQX3+L2K
i16wbKN3qHea7A9qq7XtE1K2FKMQUFjkOpDScB5+o/A2LG5vA1zcbgEqb77IB66+
2+JCUTt7GPyLYmJaarkehCmI4nXL1aDf/e4cE7wifWeWa/bSX0F0SqYS0fdgiN+n
+WCh59IaKEVhpH819suLQyJHVnneK7va/G3M+nwn2sXwGcpvQEqFulmHsWf1J3LN
miHax2XXL+UbrZLiCEYZ38roOtdSUg1jZaLMH4ZDOGXX6/cCG4NnebDElHs6tp81
GWQ+JKOeVJPY2FvFckTlijZ6sg02yObZzKyEbmDO1VXH+vbK6jMQW/Nu875kigxC
ZYeob76FMvU+reyYjmwuDqVPCzaaaLRiY5WXKGysepVTdC6nFWzaYiuCBkEuVBtJ
F3dRy4PHXEGOXZ0DXHsnzJBD053BWY7UTJtANe3TxxULMOqNjEOY2uOTsgVs/6Ss
HopMG6oD5r02WKBZ6mi22n7+FjpwLIXxPuawimrEmkAE+HolYOibUE6o9ib0mHr7
qz7J1MdO38QQf0c/2H51wXdZXWm864TnDPknqiPOMnJX2UdcDWQOCrd+0ErSAym7
DYjEYXXavC2h3SWvIfTFkiy/qpwURS7U0YArOlJnF0y0jXeFAfjFRXiQzbWYkS92
n0W9M1PdlLXm/ZfmmJYrhwYFkYSEQvCct4l3wvmaBp9/oYJFLfSe199qfdlh7l+n
idDf4lseAJabvOhcTgdmOvvt8cVZVK8ho85AmzJCpZ3cSXll7KBCwkANKfj+irpC
b2073e2nb4Nm9hXj3Z3qcfmNETtXgmMRtgwlsFgcPQS8VdycSvXbmYnsefBLjLD3
Q5P2u047cKEc0X/qf0NaeR8mzJdWgdOo/uoHXrOXzCchoHaQD1QeaySGosL/dWXM
yuc5CoggnHCNcqyN+ajUrnVLwkYpVYC7mLdKSDmV5u/tMqkyA9DH22RYGsl3OyD5
4aw0J1PSf4PFlVKam6BQbFkn2xK188QvJYSvC96wPCnojAcYTEYtm1JdMOoRfv7k
GrIruLx/KP0rHlphHwg9kVc0+vPUrAWdNbPxZIeb2YdzS99c6a/vRCpobSGqHIRa
iGI8PC79hi65WlaupN7GTDVggrvO/0PbE1nMiXh7gq3vmRij+83RfocnlBPll2tx
19IGsSaqGs+zBuNOt27OPOwu11FWEXEAXqtH6BAOYz7Ow6JSnM37zAS6Mv4VH7Ft
FZen+6mdMEmckHuf4rWuaA6YPeA0SXSl7ljy1vprBEvN9qI0RW/dPm/xYYcSP6Ju
jAvJgskHweur7w6CX9TPQiIHS9E5vJJBapj/YCvZL5KuEBX0623bZbcjKz0se03z
qBKPyTLlX/hplhGwOm9B4HCX1t4R1xLPYmTyaKAxytZwZu54B9pH7vhTT5MQ7y39
nsrirYwJx+S4tTThQM6hymCtBNiH3tqgPB53Mu0yAc1F4eJiYNHWbQlwr6CkMP99
ofPR5qqRQ5q6qo4LGPJve3gL13ugUwy8pKbrPccG5ssEwZn+ESGbdI2BOOHQYaKh
txp0Eb7flyN7/rDInGTKKDIIXqN7lsJGYGBj3ggMyYkj3IavoE6SAUzEUtcrxuoU
U4EKyRXvnYLre/rpSNZvMgtMTl2n0Sa41q4Mzu1Nw4kRjE4oc0nmtNmXLIjimghb
HA0hrrXRTz4g5EO+I06hUTxHxAUq1F146/G9qO1Ikd0rmBGrh8xoj2U0VXTgAXVr
JjncIwkY1KG1/3cFl1r3OBt9E3bJ11RexWDXiZJYU0lZ/hz3A1bFCeI2ijt9xby6
IBCbdmNnSujVOktkAT0CWYsgp+0GKWaa1SmZIrbQqg3qE2+RsP333fGnoIzUQeWN
kLQZdWLtoJVXAF8DVowCfRP/f7yq3DBb4vGjW8bhSd9MhDxshIhQIkbQ9zCcbdBY
4/p1nyywRPTfsruGVPqIz0+NCJOQ4Pg6Tza2Co2memkX8kHbG14NJ2Og+vlg5Xsq
LqYykhVkXI5k7yrvQEpTZ+Kp/cB3ZV10MiCnMqepIVYfU5zxRD5iX4u2gN3jeq2Z
47tvlzuFT9uvT9voyxGrgjZ0+4P70hJSHMGHAPN63peP/ZMp71g74w73EJ/sSUkj
xPR+ZyG3VjZxAC/7aSysxfYFO7IPzDWMCYSg7sphKI5Vu70QMQenrwjts8Bv+jEM
LnQT8tLBp76JXggj445sH/ehChYfwlMx/Ov3tXMbeKuBs/d+B/yjbPe/rf31WLwT
XhUxWiO5m9qanIzyaaVKHxdBDl+nQTv2NrNs9iGtH/6sehguZIJsg0KrUq50MlMq
QhO6RAGbfUIeNdNMNdEC4zBjsHB6QrroxDotwtfrIJiTrIVCM1JHrub+MtH85rru
Li/VtWHsFntCB5GyU/Er+hXYyg+KfG5kAlS2Ya734loZLQN16Rh7Ctex29DvBW7Q
CW7VYl2tCmZCjgqOWiP3SPrng86b6P3Gm33/D7vabnSqhor9hsn2Geg3ydusIUiI
f+M2NSEnuJ5esnNMc9nXDuAc3AUEjsvjZEN3yjEwo/T+k5bDPjp914LBdF0z3O2n
xtTIKieleQhRcI3cVCPf19/5l2zh4lqMrQE1vEMZy18uy+mCvGIrtZYmexFBJwKQ
Qhh792x9HXXpMzv9T13LiJ4HW0RcJIkEwsw2LHt8gfhXmGahseYlI1Ip7lfxTv1a
G8NRjed/Xuc33wNNW7g8OnjOndfXrgLX89PS8ibAnw38L1x/rHiC/R+qu1xmyiAo
qKz5shAw/egmJ8c0t0k5PTQRxf1NsK2rGpgS76j3vF7PWmkfpoubMw3eTzACQ/qR
+XE9unIIKQl6Tgu5IXRiRpf2uSXZfQdfMTR9zrW3huEDVis51lR9Y/e2XOun3f5c
4PIbqek2qp1DWWCeR4arkVNmInMWZphM30in5aqtLcEWBUeI3i7NAHloOgDgZPUX
3GVGjwi2xGD7a8Knp2hURTi6OPWkBeHWEhRdi/XIbKFA7K5Cgf9xmYueWj5u9lT7
3m2hCYerg4hk9qir7YxQDDt+pmLFWXL9gKArON4pvnmZxNbkdkB6H2LLXTxs47A1
7nKrN/BQR7PSmfgprZyz3CPsc0Bbj5RmsKl4DXudr/bhsKHz6zzwiJjydv88T3uB
S+3e1xCnlN0hykWvPdn80y76FL9DPYg8X7QtM3uAd0PHaNGxOCEbng0HqE1nFf5F
LrnuWhvXBoTrii9MH9i3+FUJsBNotz8TnCED5+i7vGs2zbLyuMc3auDplO2Fg4i7
Tn4rMGjqDXNUqZoCBMdGH7IatTdnEeyZuE4OQvfhIma0o7DKc/Fh8HdcOWjoyTc+
IKV3ZDos+RseeOEJSwdCreGPWsCD8rFSATrIth5p0IX6NqibkF9Z5G0UFrkGZ0y/
DudKQ/+Qh5fi6vo/qpFM1u5S6fUgQYD23njCHwuvOSUSXpiQsDkYRtTesRQyOhip
9e7Apl9VteVbh9TNTQKbXV69hhb2fhEB992/wUEmWqUlIzmYsYli53rqdEUNnB+f
oZIXQKW2lh73dagbX77NIwqgdeCEmjNFdSEw62NVxYrz74vnVM7El0JTmZ+DDisi
+GJLE8RhJIwua3gA+qwqIrW0PhZx4E2rWHD9aJwTZiMpBGPRzY9TQUp3yIinMP1k
DqlVWR52Q+MkzJ5IplTmX3/FL1P4erhGT9M7MGAgXq5ifqrTTAuHknYqMYJOt5Dc
onACXm/H8KBRZZeulAGDP+Az6XHgFBuDPtC//BvYD2BM/MiK6yYE7tKjemblKK8f
HUu7BY2I6008dZXQtFCMTdMCVTULRZ45NxUlKGncsQYHjnBMk3d64FDQQbjHPnhg
yWYqtp4OOzctt07ZOVe1SP2Pdo2kVvJSdNBL+sovimp5ej6izt/Z0828wX5Gl78z
EhuDc5HhgeNGkzbboJbNnqzkQVe3x71tn5JuoVofuYuTnwOSNlbw4J3P3zVmObtk
KCVEQ5ZC8g9lnactQivagGX7aDiJoXDRrwXQYjSmvOqBdknQY1d/vfhctwPoTg5Y
8beAO9w7vbjfIAocFCgSmHJkbHXVs2Es2Gp/65UmrOB0Ej9Uzvd+qq1nUMf0KklT
TF/UqGBBrVjE1hlyke1mprSMTTUvXp9orRehHXlZAIgyyEksapMclezfkBS76vcD
Lhh+WwGZ6P2jy9Nt1PEqkzO8eC4a4wwME9mynKYNnNZ1KPx69ulS+w0OMc4AXhuf
4Lhx5FbMNfkK3cuPd4P6KIJ7nMFyppX0SgUKubsniGV1Y4acDPxoHRoKVVwPnL/a
5cHXc+jvkbNHXYKRGPvzJe4kaM9G1YEB6cG7Id4YCuLZEqWE8FWIf72jJrr99XIe
YoZ5ioEGSrZNyOuK90BBH1mGD5rYc6XRcQi+ol1UPVYYwlpQI3x3NzRE3JGYdj3U
VoJ+gGnQw8SUsgiifI1qJUwqC5rzSNvep03H6Q/WRr+muPnRnPZag4SSrwrQJ81D
9W0AcdstOwa5WnRPIcGm+CtlDS0HqnwVA6hHHIlCeCVrAoCVw9nBxxyvxwi/xzJp
stCEmvrP8HzcMqzCRRDG4UNoot97WL7s5FiL6j+GTjcxIWnp45B6h0q3wnb8chWH
jbcsnx+RC2N8M0fdGIr4dtByAWgLrCMkjEDRNYOZqWlaJTo8c4/Sy61pk1/WI2u+
jpNDc6cXXYZh0p8lbYba1fe71jL8wn3h4HV4Zu6/Yzb3DG38AUW6jTV51WbiPuv6
IRmLsG/sgWVizp/P8z69A/4taows0dNvRYtDtI61ppfWDOIsasA4n+ehZ17oizxy
RgN7qmmSn5quDXLhQc/Aiem35TJrXmf0g2SsMm2lxMmf1Ffnjs5brRuQ4A/giItE
DTY6/dUo4HeOqgLlUw9ErdzbVmON0hYMQikEliSzsPhDhad1CqPrDQ8A8so0Jlb5
3xDCmHgquvxzQFVCmPK1nsrLMAiQaeSkTashj2Y7ByicLlp7yDcgl0isgrtJrv7V
jMeY7IVYl+fmscUy6WstDsb1oA1OFxGeLizsj8H/fCH1CY1pQgE3+QslDYCTciT4
Qh2G5Ip4zPZhF/ZBWltkXn7KbqZROrrDKRX6yNK1CjUilYaEP+mL9M5HNsjh16d5
ovCbg0RBrHUSZLxXdTcDB3cX+RKCDg4m25dQVG18QhImt7/z9rEqcYoOxM54sYxn
/R6kPJU7LUwLknqPtK4ZoVI9MU3wuNtiC0jqUkxvddHdgwf8nKnx+HYTqkisdFo+
bHatwUaTk36a0wVm7r1pme+Vbd4f5aLigk6JqmtVJpwSRagL1f7wZhHEzSOFHvCk
DApaluopeC9h82UNGUnQUnAlPDXxVEP3hdTJ1LCNKZBeGDigwB4g42jloAinYDOl
VQ2JPMGHWBFedvgrp/YBmDT0nc0iUf2jKieXQEW5u1BdXcVwu8acrLzDjZKfGQzk
dK843KhJkicVbaVAdhXZNrjuF14uyt51KPaWfEI+zSHFeYms2GPFQyKtrEWBHCEw
dqYO9aY6d8yX4wdzQHerZKyNi+z1dbrKQCL93DwkJ+3ZztBUzeRtGMwdCw7mNXPJ
60fuGtuicSN96yi5v05A5RCNx12leC7zZf+rFN8Z8U+b/T1b4PbvA4EF6WC+8uSc
6BKbQ6VNftwQEgaWHMxG9F04HTh1S1taVPG4DvlrbsucpUreZjE8f2tXoYEwHzoJ
PKMjyQN4rt9OT0pR6ONSvGqDAtLPyDfl24qnyHZY8Dr2/zxbnmcNUGnytBQNILz1
+Hfq26uCofT5Az6BgGL/+gF5zFnZZAyt0yIcfc1MyTwjXk6ImQZX+lEpcVXGe9C9
3mAmEuzxGImGxfpVPLOz+mMkIElqYg1L62E7kR6fNuAqaMNdWK8wSR6nbS6XpMBe
rYsBErYrl4BsyTi+rcLnJk2DShKoVbvf7kYvl7OdDzrU8KqW21paVnKZPNZD6dg6
Ek0I8Aet7eKPVatzdavh8wwIppXr7ufXEFbLHaOLKHA4dxkiB6/pk2i0zQunSE2g
tbMmNzm9lianVMZUj/LSH7jD32YVIm1ny5CRp2mLJ5cexc4cFiphbmm/hZ80afzc
1V5DA8KbNa0+h8YZd4MvZkSCVO41RIgCYJBv1NSHSCZTZf21aiRhOP77ddHeWhnT
/f/ylrrKu6AG8Oj4Ygfrfcxe7Up16o6cq4GhYSes/7z4C6tn67NwOtCcowlSf2kC
BDZVqW4Ii+ZJvRcOsuNdRXhqSJ6+flILKDcG16JaYG/vVUJJR8y/P+SaLH5MDsv4
ricpF4GOG38wVPmVJssPo6fecTQZwJoCdGDwiYtpT3DmVl+P+GofQHmgxJWa6HVq
9OB5WI+vtSO4vSbSDmWwpRf/WdIz0rsFoBoIYhkQthlXIMkzzZ2I66tOFWb/ZhKN
cj38UyQWUI3OehvEJqSGE6HwlKmvT9kXFDY9KvOAzJMmsZEvggTsLNFbITjzs5QA
Afa+n4V6kHfIJGLqMf5T9uYoP1FNcSaUKqISXyltrN2s/mctyh27BMieZadZgGkD
qSvnvKK2AQ3DI3GDKNxzowUMTm5S8qc0aSNjYDQxgIdZplE+QFmortuTiyi1kCaY
O3fBFAGXmePdpOYtk3y2sEreasUvdpWWT7xaZUkf/X79JErtsjVgh7dWQwbpxUNG
G0yZ9ZjACjHW5ReqpA2C0RqBKYtL0mofhUgR1J3WtA6FEH2V+GBccTTV35JoKBKV
HSlwcPrcyvQnhHc1W8Kn7G154fq9ipILKi8143iDmz5g4XSTOCgv1ko+X0DomBva
g5pwXlKGYhGvU29cAABUdl6cCJPqXOya8nvF/LIiyq4tlWfluMVlFJKR0WUs6nr6
fa6PxmiV5BMNm2uLD89HfqKx9TmS6HDEx1Cw6i5uN28GkzRjcaWjE4I3nGf0yrQE
+ttivgFP7hhFDizSKtZuPrW/lftB1y+p3BqPa+AsDmHmBSl8FgpQv3CN6xg4FMNf
AeNHceOdKlWhaUsH6Ne6R+OizVp9sKJjfNC8lNkFaOmREzXveTiq8b3LsH3wylin
EDLQDIj1+UTFdOFC7oCKmS/zdwdx5e+G/hDixRGztI4izPwIHGVqni118xleGxUW
LFEb8atZ4ygHxMD3PjCasadtZT0lGUnvzibpgEl6Wyt0rLHFbPjOTgzgbXLX0gd9
sGAtreoxn0xxMEtChZ69s5SF7K+3sOZAbRY4aWZ4hi0axbnmUoITbDPsO6RA51po
bIfx1V5Yh8vJJ0Cq7Vd1By6RQeb/0YMHdl6ENfxdInMRII7D2MWfdxmb2jttk3cf
020aktZ/LNOyiUbsa6pAMTjsVVGgM72pKIwOlACFetc0rFceUYv5+MTCb8OqSuYQ
cTJP4Ph7nbhbbKevBQSQTUj7CVqAEkT8KpR/hL3UYAZW57jaILAp3vHMW1q0jMpj
RmJF9zmIIqf/QuaNuRC8kqCXGm3oMRHqxzi/byxCEtXwLMlB6BKnvHzADGTUaJ/l
g6GIp8HzvbV8HYMhu70rPy8ULSBreR/68yNmj2U8XbkSFuxvULW0dfOuiAPSO1kO
p7QLiJfkc4VFeH1R/3y/7IvGMztSz8Q4MfhO8tfn2NmlCDomnsh06ei4niAMLEnc
YXL5Y8vHtEl3Ey9LmuZf5T3Pv+0cd86UExZSXlOTEwQjmIQPA5mW0NU8NcDoambE
HJyusmy6wTpdwS1f8PaBAg5aqCs2rAIhn6W50Y2peByzNfhvT2CPpJSToJPSva/A
qq2WXVx67XYoYydIea3Tzdd5CA+YQ2pRju/T9DrCd18VVYx60cqXLlKpVrocTMTR
Z0Rnqql/55zynW6yCpBw+OM7QVRxN4TBUPjmTldtBc1fdqNc/MCLE+4reZtD3M9Q
pWtG0Dh6MULW4XZ4FcZ3Ebx7AexT8lTLN28jcgMlZgOakChGBIemzixJXyVoXudu
+fbjeugpI4QqI4ZhxJgO16oOZUu99whXi8BVPFV6rGzvgVqrd9nNJxUweUK37oHg
ytgfXtXqJbV28AQDPbSyr0Sc3Sts+glev6KPVR2UKOFjegzaX+rhTnj2IZFbuFfZ
pijJvM/uJhB2+0mliUZop2yBWgxUke57+3hpFOY6kMTYG9oPzCU6qSt/YHDX40rf
sMLpF2wgK6RutqGuU7vRWup3m3vXVPTvGMtaPxTw5VGxiHUuNfUQdryw3y4QMZ/z
Pz1H1y9kTdroLYvFGrSgww4VJyU5Iq8IqypwPv9YgEbx+2pd6kBFe7c5ETLg1OXA
1rQKyCK168LzjhVwJZq9y5xsyKGWaUewLGMUc8PFQpeMjgBxPdIbOLTUJiNOdK+9
AJzm6Vo+TFNRVue7gajpWy0Qnu0Y1LnzWNafiTFmRjKiFa1rd64GOl+ElVXtgl9Z
crl+3swFEewefjM9sspCYWKrv2pD1KEw5XYutNb9Ily38xrtJIw/q9xW9Dv9Qw0U
9HpECO436OsTuhKr2GhwQq5YS01qWQVkW2IV5QSOSIiGj2c89ZHQANHm76c3W6gL
hVSmWxSYsk47/PUKQYay0k3MtqxVpDCQjrhR2KKQ9pkYjCyL6wlzkab20VULDXI6
umaqYutEgpKCXLEIOLDxncbdK5zyivf5/MlklZ0GnA/qxUDcnmPgv/Fzl+aq6CTE
0oHShqsc9l1rlqKdZA4BtDN6JbH+zo0NLGevEAvGahRu2APKWi8ZJk9EIgCLrMLc
YdJqk3B0VirTNCRrHwhHASDBb/ksYDnjfqITiosMzudsKn2+oowQURzbBaj0fUJ9
/ZZiq+LOhlxU9v2Ox/dVah5EfGQ6afk32EeJXJ/ZROX+6c14yGM4KiSw2v3T3Ov7
sZLal5e7GWPIliRIjZob1lH7lXlTxqsZGtEFmHj3loG43s6vWvtMw+IMVEKiJWw6
0xhtWHffNh7R/PtF4YyAWZPofIOBb1+T4X0h1hEhomGszbZAcMQQKUBvXeWhlCNz
NwMK1oMFdj7Ii31dwsLhezGbR58l4R2VU/h6xH/Brnr1bQAUJFyJKPrSI50CFFZb
LF0g6mLUWBkLJOmKblLOYctr+0VYy6aMQqc39VxqHdLcbMg0YiLfbmWa3ceRkbxW
Lbk+VWIoIcbEF9UNMhsiN15PHSjGhah248hsic1o3tMZVWEsAkPNzIJbEgcT6mT9
8rW6d7z/7No6dA7QEtCaU8/stq9jKfbsde/czLhg9YGs6cWv8MCOCguVXLbl7WXp
Bk1BIgZt7kJuHpbXMtFqGyNDlMsQUnWkBfY0mFPU3+lUpjUX3Buk5LqohjR9ekSQ
q8qPsJqvqRerIvIBctCUNkml/Ua94XhCZVGo9PznGRikfc7vG7x8RrVrxuohDfX2
baorh1n2B/2uWoww13I6dtxEcHmv5zi2GuKwlMxVnjPfAgZ8guOit3aKl8IMoFPc
t09UFxVvR7qqaqSwIGRsYKR7yfV8TG8BVMxJ42MIUjfmZ+20rKEvZeGpycE0KWE+
CQi0Ca7jPQAYazbEEYa80c9RYbbIol1aqm/iiSz093MnFxIkwlKLPhtzqbsKhCay
dpmGx+jr7EBiyKKZb/ViOkQ4/5+GOFfURxdUeCWZrxm8YiXk2aa8oXWhcx+mShtT
mys3kmnQ9lOw30MBMrZYDhSuKaKgd8snmtgWDruoFk53yBRlsc1ftYb1L218xKIJ
VeaRzGiNAmZjmxuahgJa2z6uwB1G1oU6fE5yu0bOlVR8Y4ieLpN4gHCc6LZQGKUJ
FEIog/zvDJC7qIQhcj9S8Pbs5qnghpHqxkcazZTSEoxMRS5LcEeiBdJTnjlaxEd/
AXkRHmNgAcDRi6tU7NFflMLC4uAN0GMaIsojdWgrMEW4biDdGWhAMmbderm1KNJS
9CIe1OVrjAj+4bbyIYSI2pZ0WR1t2n4HbpbUFcDINCgV/IX46Kdx+pCtNAREx3Au
DHG2O1Dwq3PKRhJACEQdhUqpvr2Io8G4ijvsCM3J87uidUrRnctlzbw7vC2Cfhmq
gv4pwfYiEGFVupGVVliyR8BJAtbbTvsl6E8PAM8OxXpsV9IVFyOqXi9YRebhKuQt
Ly/Cd1FkiAMkhYT6dxWoT6Z+tf83CWV2bD7kiA2b7sGmBzWtdnUCaMGPB0or2zat
0lzv3LzhuRSAvQI+dOJHV2Vt7Ev/Qo8sMIadOh1sdMth62a5qkFBx+zMeKKeyF5T
dDYs/s+/Kgk/nAxnZnFN5rb6ewHQ8TtwiZGmcsNjR//7iXo0aulDIhqhFEX1nWJ0
Rb/1e+HJtV0pMDk4fUot5vlQL0O1r0z0Er7KMsB2YzVEjWPiv1C3igNlqzbmQ+uw
Y8l7Jue1qhkwLxsVaoEt/E5auUMbU1hQOyt+2obiKWSf6YFEIOSd41f1DXeko6GR
KERiwvYPHxM6nkx8F73eptC0Zd9o1gI1EDMMw3MMeApWBpCLK8JjsVMdzKtNPacf
Wz7bO2vlgpQRuaV9E7I3P037YyqLwDie3GLOwlVR97UCvEBhCx7tKhq5tH8Vw5+h
Ga+G6b/0LZ4TED7grf66ztHvTQHADdKAr44tXZSI/iV76P41JLjp++skiutl8qm0
E/V0CIaDjJjurccob+nEOZw/Y6qdE09/Esqy9xE8x0vBQo6/EIyIT2KghT96SFhx
pMT1kRiT8pbR1iwZ8F/J2LNMgCcmDdlJupD4yy/DnPDC4Xv+15y0Xrx4DiE7WjcW
4u4L2qzWTCeCefDDF2rWaq3ccQ+qs8a3BuShA9mDZlbFO7E6Q1xfPMf6P/vaysOb
LgG7WhKgn3snw7b2WVmEJUPLBJnwQHDF90ir6GC6S7UGk/smCvdmGkttjSMYOqUc
AfahhJykQ4EiLJ6C+0/2fgsplhGob55El3K3djzFXIYosJrCZD3g29OLySLsDJVc
us1Qt0touwwh9+UK1ZvZi1hL4CYBc9Krx6Crya0+A9Vhu96JRbQlvSXv9F7K13aS
UgDTqgQh3xcV5Jo+nJBnVKVS3s4pTDZTe6+QErzP05KSYmbcxZs4EdlRWU76XJvU
wS2qG3vO3WfzRchvQFDFg5jkhFktBbKTJy4qxTcyMVYULraTdXir0mbAprgvoVMJ
aYjD4xuuEITEZp1hrTzQBgGto/ghFKyg3s8xGkv+0WZgGhkp+xrso6satXXvimnA
DH+JjIU2Sa9tbjgR67K6Fp96X1D+i0xYRWOHn3AKHUKFncuvJ2dfh6kS4PrJip+W
Oi0SxYVIMLhgiOJQrVY5vLOyRMO6qKvrU94nxmv2WFVIaeIiuD5GIApxZcju/XrC
BFUVtygmGBwGg7BOnkjnQ2UyejcwPV4fdW0TGUNszVaAw59xFuCC6+JWtAQycsgh
ZFBrikYfYhX2pcazOXx0jomJgzY5pTvvdtftWIQ/gUUOaO7vzw8sFSsTx0EpoQKH
7wov8T1FS0hHdYsinGdSJk72IvOwws8IE6PUEbw6li0+II203OOPyCfSGqK/VeFj
ZZ6VawKen8GpYN0qA+UA107noV9EnFyyb0DNOcLK4GBq8fqlvWzFQLi7sWZ+44PL
63sd7u3Ejl9H4dgMRjbZUZVcOnSxERb6K1/C6d2eDXJkIXW+v8qFgnHMJ2PlBEgM
62YA+5OeJKMossl9R0tjzJ404Uf+9Qnma3PDd7Lh9WgGQpSUAc0Mxo42rZ43gJiK
sK0Mqw7NsFbqSScVNznwApoB8bKryGw3PYQLQDuJwzrQxCXwnuM1UFmyyeAeRHgI
PZxlykQ3YwY08VxymMxfZxdItj6reUHE5BvFWDzag8DeuFALF0VoXw8c2d5/wsdn
UG9MLdMHOGC4xrTASdeVuhnyZtcoSq4uk6EPIPg/me2QvFxbPZBpD/cuJQBh5oXC
6uqozy58iSBPCp/ifIyd7uOHBNOKkHEPdLDQF6zHlU6fMJDRCwJakc7ApvreZ4bv
DQZcEQDeyBRlx32ap24v8zX2REZGU76HTbD1+tybpxHZXexuewSRlrRw90y4ohmM
sFuLgRFzAW3/zCUPSrqzTVcVTjl1ASLkq+TRpFtprVADwYSzYTMmY+0vkxFheY77
ntSbxLAmznxbYA/m0vh+J4juTv6+gtSr2CxXInQ3TRjmeU54lUip/kLLfPEufyqx
T/Uvh/a3or5hpJNaOVFoyEbXQhUzfWPsFDfQ1gn+4QzTMhJdrOXahqJHiTHALC0w
m7gLEQU1FNjR3F23Q7n9P/GXAEnhvIR3PzCB2lHn/niNgBsReLpNMYBaUrtiy5FE
/APBlGz6oPFx70qnJXIzLwN7zL096v1L7fb6qkFPktBjs9/nCRMuhDVpdgCOEKeE
tVmsv7QyBDkgbFR1kAjdRaK4s34st3D++d2oUA3UDBQT0bo97+Qo/CZBreEx+EWF
6zLxhPsQfjo3WII7HOBi7hpFTL3ynj2YDPTAM4275w9W6EwxU1xVWdSX5qhizqXp
qm7LLp7pRia6UCIdub8Yo0C+OSG5R6ujqtluzEaAnwCgf976r+QPF1LGS0BI6JGc
BBo4slp/v4m90oW5/Tzviup9jNU2/fdiJ0rkL6hIeSEHZkozYMZs5Sj+ONJegrOg
QP7RsT0VhIDwLha3J7VDZjuJNX/Nz/p/DIOWlqalYQQOh91+LUpZg8E2kFeVo1+6
beYqjmI+uVKr7fQvIpiEbtidZdjXBzBNfaH5VwTiQEwnFNrwJiNfqXHJYQrruZbR
rAoj53BTlLKZShej9900M9o8F/RN4H7L1Xxak27did4WmiP8ZcElMYhMSzcjcBwG
iQ9fvl5JroBWAev+d4NWQM3Ey9dqMOKwMcV4TgXN0WVBdoKuWJxVt4RSoVPq4TYA
x2v96rdThTfr+R4aVp5NeSkr6yIG3/UuCvHlfPsMp+BLlM0439xqJsyVM4CLNBFO
kazJg4eWFqh+Iuca/1r2TYvnotMQ+GODDIuDld/sZArjwitlHmvWQUXn4F4ZGXgS
zflQgDwpntBHukdRyzVQUjE5kEj+b010kSX7WS2Je56UBYJMx9/ToRFAYqpLX+eW
Ui5M39Vbp0vaEA3IfeEkAC5wRQOnXdCKJKI2lCHLZm00yp3fZIjSb6Ugisg28sX2
5BGwcndqUPCHMPYmYwlRlNGdFJYOcJOPOvgjJRvv3RdM+MsQXadFlDiqJb0eGxTj
0Bp13Kzq7MWWd5BtHbPnh8sjDJtfygzT5lX966j+Vd1cI7itkILsDA66W050Thfp
1SwUaLqbF7+bmHg8YdTYoF11yLYO9YnV2qbeEIQ2CnXSoz3qfKUSvJkctrlZs46f
Nbn3A/Ut7HCkD7CtvrYe+c8ITVMomc+uo8yIsRNatCiz4KAsngIWvGRo4/ToAfbN
do32r4lemnk59NnTjrEeA0iRsRsAhXLTrb+jQoK7Vw5KZxJwwTzVQSyIdTrZRUva
AKCRXEmwSwts7bwy7ssKv1Ju7+HmLO7wFocAmHgmWD/B4Q3Iq3bSc+lBHmoIR6yj
8siAS7BE1qxuuJ3RIvnr2slam/TrdJhqmGpWd02cxa/R/TOx8hUzmUr8mX3v45Yd
QP8TfP5ZBgMmWZqXzTddGQY4faLAdum0USagJGBgDqnTJo6fcK03rpXR0BuC4kZb
xYy5rJSxysq4RwSdRzUz4yQeZSIMdQrcxRfjIt07KU2H4sMgUhn6QcdsMb+kxM2R
ychA3Nb90wFuELlfRvP2dtiTvHJks7IEBAYaH3/0lQp/swoX5O5v+eZs22SYuA8e
4A8a4qAJFci117KsBNkI0otQZQHQDXPlr7aCGgrgnjO1iuo5hl9bbdem9aT3KFZm
WQON60o1Yp9AKYcZ2fzKPK7Rqimbv6Cm+nbJO1Kx9KaWhmfnbmC66+sAd7T4pERK
HqdQvdgWDxYYGowpOiVtmdUDvouSsiezbyHWShzOaBdNgbMSwskeiIslWkjv3JJq
HEckIR6T52JmJzQNRU3fYj+42NQi5HmpnUOWht5iDHKbnE0FzcVn0LdV1LlgsXye
hqoQJeqaYMDZ8HZWkYe0WV8X55RryujcckBEVAvNOp2IK6oBUjhuKegW8XQXJHyc
9ZAYjCfc5OeB5V7VxXXq5um6AN4fs99k6q8O1cNbB0iPqPKbxgAPjxs8Eow2DmL/
t2MIhc4hF4GH2O8DrKshwVCisXMPoykplkI2dji3RYPxPZxFWq5MgIAQCk3A2bMC
R5aXNAB1GNzOnOl+ah8D4luxz1pEGU+sOI/2nvnN3pmkAc6n4aUknmMUd7ElWXrp
5S+a8QG1ycwS2ZM/Uu0GlSfEesWpXWohw3OBXfaTA2BgMu4nbEyGU0SZg5gTYuQO
pzBEXh50UzTtSz4Z2ttt3vTka/PGGTanLpbuLseGNFNekaBsfCs97yhMw9WtnBOR
Z61CX990zLPTs2kBInJgXBOmC6joWLT96xAnBIFJLMBRnI80OEmrLexhoZQkZEk3
R4DpT1C7InKIhkvO0p+h20VjIC08RrAL+0DPY3RSfJBJSuKSHAgiN762hM/GH5bg
jO1z7mWTCR3wqNsDm1jaP29ljNfdS/r92TZROJ5cvpUZ0lOZ/0zYWrEC4nNU8v26
R8tBa+VdwePAtcKEtPkRYskIjwJfOUh6xLcA1cjrieP2kWfTH3/R0EEIE0wkpCzk
OPX10ezHNWee3+R++3OOpQoHTVixEMLDcmolDtDBerhKbYuu39cjJqxQG6+ubc8V
SJmudB/ZF5+MHk7Fa2yxQlmGHbW/OA2aoQdpe9Por4sdZorGdy+QmaeBPWs8pSSN
bA9BYZ3xUReYAVtfIz8c3oq+cCvqOpaDxpTaX2QeB3mlHQs1Bj+Vf3g+zHMgVgxK
26At3or/qkeWOvZuD5UfsMVy8ldKZ9PavHxpvvS5Ok4CpJ22CRCy/wLaeUgS7x/V
Kf4LfqooScYt37fR/+dfE0X+3syLSGUfWKQueXp8i3q1Sa3FY+vR9e6iGrhKYv12
95e92wh4558kk2Rxney73P0HMua0Z5TRHQJgGvLnxrV7Oq1ESo+xMkrGnQFxkHT+
+MTj3v6xFLJC+8kK8HsPfFIxv9rFvseemoUrnrDJ8FAkSi01NP38Pd8zGTFql6jQ
EmYeUB1AY0mCD0fCaW/QryZaTGoG5KE5nPuSGEn3jnUXbkD8+9dCIdIe0KGasMdC
S+dVco6+JDMCYOjRuT2uzNUdaZWorxukzZuETzd1kZLFTCIjvY6gZHrGBzyUuUrZ
mMljBC6k7AXxAf847fYrHUBwTwss8dB3VWW4cblw48O73NPwT6hd+HKTAlG9KSwd
mJtDiv3KITsUgVtqemELpFoyMf5mm4yeTsWjaVr6zmEHGbCtg3mLmZBDn3SFI3jJ
DO1vaF0woSumaWakbwftAKjIOI2dUSmlpTsCFt3oqVHRdRW4iAtWGH/h+OdBf3dM
POELLQ4JMvYLeMQuVQ/Y8w/O869cReRjF2wzUUMNhwcAI1nJn/aZa/sOxahH0lBr
IgFRuPmyju8bskWdlARhpR0fR2Rw3aeqDCPtixoMpiawPj4tEpWvydm9HUh4AVDG
TFABEeewo4nVgtrAlH2hcw8D6qKeAr7RccvBespxhnKppIaR5L7nBn19537u0zc5
U0fRrQ5gdMMb1KqlSZLPFMP7fzWeej/nh5sgywN3VyDPDtMmUgareXVo72q1qZoT
1bckrDL8q5skRTRNRgCiZga/rlIsgLJJdiiHTsIs28LCm8DQDa3A8dtSSZFTPE0F
12XgFnfJrPvjgw2LegEAs6ZE+y5v7zgMSTmjBY48ybNfRL2w9C0e5DSFq1Lbg1vC
BTRgBiRyjRVEenjBDBClAy9eKLmyHOpCXFLj+v5iC0xi5HZGZmGFKWlCM5Cd2SL1
L/vKbKMWMx3RZSyqNX8/7Vjk9uvd8qQaoQTvNKqBZBGArilB8KuN2kzeugDeaiKd
MkQeA71oazMT2gFExCPMytwgixDJz08hOQKoFFV/RDOYiWqct9m2fvUwKD140G+t
FgfuhqaZWvCHtxsF+Q2mBn05S4V4z+pQ8/1wWWLPmkRhQQQ6Jo92oddd0QPGAYTd
EJwLoLKKWz9K4ketLpB1qMeEBFnlZrPWAHJCbvgfW0o8ectL5JFC6rQzV8m6o0Cg
1j9Grml4L7Mrzke2mZ+woerssBBxYT86yVLN63qbOk8H2hH2sxBzpe4GQl6zytq4
BXBzdMooQUM/f5ksYp8iyDdULf3tCht/Bzyh0tfsNQF1pHFMbZnd2TM3ZJNCoC5r
XHx6tEQToJ/8AUNZPuJhA+L4s8xklV7hselDftgDosGcaSb57TJDzk1TG4LtulVi
cKTFKptBuoLry1Ri9GximUIrq30RyiNWpbiQeunLXYTigbEMoeRrgzvGR9AFBno0
Eg5yNeC+X/ZoOplwRQa8FiXha3ocQ/aRab/G495+zvxS7uN+YU8aY2MVs7smhcxO
jdWI/wofTRbK3U26wDDc3ghdkqSC3BD/6uS+u1gZzYVM3/ZeZn23D5QAv0bpRta7
aKe5crVGd3Qx207HQyYv2YAa/fMB/f/c/0/1ke30pHZ9tvJGCB1qVyuHaw0FC2MZ
WGFo6Za+zqGXH9W4rnXWnXx76Ryln2mhp7+Lt+4aKSUE3RAXD4yGj5mdJL2dszzf
W/oiI/C9uB/LLj0O2z57xrgxMHidDVT9UzN0omiyfDS4qe5wjd7mKavkjVqRB8JQ
sl5igmkle2JbnAMxohjjRmzbUOJayVfUTBfO2p6it7ra5hPYREkZQAxbR1EoKFJh
ewMAXvDXxx7wvKffQzGcwRXxev7PhzxnF71+yRTBlZcRiSr9xGq/gfcRmNNwaBIN
sk0cIWjL1zf/5c9Akpx/7Q3325Em4RrCLGwEFdoHDXWTzj7qE9dYv65FWkeMaLMQ
deTwlu5K3VMsoG/I5/02Vd3B6VaO7cPNU1qfhABtfcolSP8Pv/NopfNM6rXw5TjJ
Gdd6IsSlNOpbv4wcsxvLlmevnmZU4gEMoF0Fa4gMAetFxXu6veYuVXTCp5KHdWLT
y6Zu0wHUBKTCDWONBJpa6V46gzhjrp/fSiH2ZzURWParNVpdJJdOdZS2mfT+QTpH
sJOm7MpfZrzZGqzmnq6bFEdxihwiLXlwsDXM8uYqpBTCjxeed4nNb+b0FcVikzUj
bQNmLp9cGAwJvDaasc6wL7pQyuKwXCSio5gkLwMqce2CqtU0CZ8G1bmN6AraV6HE
X6AwSkotOXgKg1q+lVase+sozuyvjeYelQXinWgJbhuFo7Viokb+zOuJ0o4zaSpY
FrzI+0Mm/yKRumvz6e/J1hvqUbSXla3h3CwLUHosAePRaBbv9rFKJck+KvJFZfoV
Yhdt+GMDDccEYW973HrMjDDKEN8REKAxOdaAzofyx4tR3YHP6aqQ3qrsI8QabsCb
Jd1ccsLiNQL/B2Br39dCOXtPPUsBCxe7GpZmz5Ecre8/7vxxyjH0ZJGgx1Ek4Euq
Ye8dQkkI7zf6bXesN/27qNZlzELvA97LRNRJCggamnLOgMA5NsV9K4e8sTrxgeNR
8M9ThilC0+bK/XhXWYIOyBeu55VG5A+7AiF3aEt1wcw/G9vvPl3sy4ToV3hcOpwA
oeqUTbSM01X1iQyBAVbIMTQRzBUDTN3jeHbLtKPt/2nr74tehSVDSBJI/Mqps1C4
dpDtBgfmfHw90LzQnslC3s6H53pkk0P2zgONyo3DvB72WH0qZF940vO1Zmip+ESi
zCbci7qWs2ECeuxDRV3WWHwNBg6ebb5pTzLe0JSLiVWsYKTRFeqighkyh1r5OOFz
XLp3Ww9v1UQaBSriN5ymBIME9eFRLi4IEpeK9CebpfwfZRuAf6OiAKd4GxUqKwAy
GUBv62BYu7ecLUXvpGolRTXwHcucdpPNcq5ZiF8GzLvBcJ8ogMmEBZ/kJDejmfv3
chhVzqqUvzByf0JIvvxd4h9+Vb8kt5njVMMMG3sjVA7dJKdX2oZoIJHMZ1nPDM9c
0v50GhYA+1oR32ZozQvy+khsIbFZ6CSqPRKZyuUDbkspg9gDI36RZ44soWuQNnWQ
Rx0/gpGT7+pJY8S/oRD2x/HOvICVPLsLURHge73L6jgremaTkCd2uVsg8rEzFePW
MI2RVwdcJru7aKTfdsMuBHBXtatJkeTuxANjbcRKfhRQ20RhOZCudhlAvq7vA93f
FeNUZ315RcwlaWgwxMQaGIwTNY66Q5sl7agzfkl+Doww+9xfmekG0hg4CuSh7sa+
QT4lNFS25OfBL9wwD8O7AKPke5W9xEQpQ+JeJrF68hUS9p2LQgn8rCR9x/CMYJJo
3UH2OOyNpI10AdsSAisUsvURW0+JOL0cfZOqoIPF8loMVE2xq95OewOOnmJMoRu2
PpXeuWkR3Ks+oUgkv5pdfx2rhSWy8HnVWNLk/4QJHIaiBqpsLZiEzaak7Iy6AH23
WvQcowZk2crj8L7s8h1bDaly/IZQVODDFALu0OPSOMR+urS99oJriG6HKjyxS7xg
PPls0eUFkbwTrYqPrbcNYcddbPeF1qPGVA1bWOicj4yaJPnJzbMm9T5hMbIIR3gw
1Ivm4p7e9+esP2kpRNK2NiFnzhVkQ+2Zx2jPQ+Uushr6PMUUK8hWgqMSdf3fq0e7
kX7jfUqnTn7U+O9moXckcwbz4/Toq1q2Tlp1yMdh6oawbX3j+dF4voTGCNzcLmoo
1qHfttfhX7zDyg+6I7zXDUHaiMb6idYOQ3PYTY11JoiJFYR75STueaalg5EiHk0+
Z4MKpabjFpXvxC2bO+gqyE2o76/i/mwfXO8RLpoI0754wVzSOIYfray0hip5r2eM
FgmcVOcdL2prmhmv5z9BPmcpIdsfjFXnXOXuBupPS/9qUfucfhR5DU+c385LJ8wa
+l4gR+uNbUkC+rPiq7bGxyv49ne8jPqbE0O5cbXAYP1kQV1DyTB+XX+NXs3EY3EA
hot3u+XLuDTnYIln8liNnnYuItQgcU93qUox7X+dwOSoMQB9k3MKGWnD8hhwmvcw
YTqRJwaig2JiRcnV4qiWTTMqfI+Y06/Fl5iD+lNAA6OgdoOagsMXL11+t0ER/Ub6
w14kMoaH1TxamEjn/rFPwBu8jdYZXu38Jefa3DKnFNYrSzYclR06sB8QlerRTbuX
cnzDUJYy8Q2uLbkJ/83bsxkPMY0x45CW1GYF4KdonS9TLMKZlIE2aMmP3ZDncfTY
XllH9nYXfNEM0/VM/JOfzyu9PiKANb09JMT7DNQ7U8WcEqK+t2MsZvYTLTMgVtAf
IO0CsdbxScnu3U7ZGJhm45Lw3VpZFS+vBxivWim3OGXHHaOCrKEtSXdtBlu8Oa76
kNkQ3zbb3LYvbMLadbdVg3ttxxqk0zCIW1z39Cnu/Fb41lsBVAtpGbUViLyEwLLJ
O8NM4fCZafjK2u/0Yo0ERQ1T3SmLvLpztXLO2SJ1y7K7YBTl9wM/J/4y3MXoRRo4
7Mf7ySewDUD1by87aIhZP82zPX2NMW+E9Zf+wTftODDuSf1I4z0qEsc+t1Sztc8t
z/DWcajSk02V8PjNwpW5J620T16xv/r0s5QwuIYCHKqcXhJ4PBzbrbFRaRqxdlNZ
+4UIre5FfEb6PQQ6DvJ+URXH7sgUuZ4H6icmXham/QvyIJ6O1cBuAR22tW7FbmVZ
31yzXg7xLfXbpho3HH9KPuwm919M9B5tRRoF5ljeQ0UwGNZ4HHAAuHAsCIzz0b3K
YOy2qdk7Z9v/mwJfp3FY2ePtzGbhnHuY8KY7LFBk0/+nA8bTGC/9bRsS2esAvUGr
tZRBeN/8jTfEYXxMcRzQe5t4pmQ2nXcwROmsNFzJ/Z0OypfgE/vWMBRqAyTDAgA8
ZmRY7ygfoKCp5drq5D1QeseMLOknvn3MsZUubm+Ttms9y4r6RLcd/dbQHlW2a0BD
ZJtB1JuW87qUI2sMQ/kqkqQrKHrN0sZms+SW3bFMS1IQZ7GJJ6lF9yQOI9cUKZaH
YWiy/Q1w2p/3eKXYAb///xnBm0wrRmv8GHdedXAdzW1LAusNgTUZ2E9gy3IkWjcA
B87YM3rdYrWL2g4oAdWY4qYG7N8TKMvLddmHQywUPQuJMXcw4wd2FtfYifgaciBY
HLnzeBUKSc0QXJeogc6a5MiuldLUzmzh1BkY7SOubXUJt2eKf2UJuNWVuA+WMOwt
jW0fyYh/QFF8u+LAkgpL1k32bSoi95xPQUXAerLHrEzOtO+84ZrzXePbgOLXNVu5
vAbzwTcm0Z7LxVAUmKS1cMOSCpxL4ASR+5f6BGZcTdkDYf5x59EkzJsHZ6IoPDAs
vTVlwqNMyM/W05jXQ9ZFYJrumEFQL+2QACkrs35txJMiy6Muzol1r/qrnvaL02Ik
6Rzpp4voXrerg6/7GAYBk+nbDJJ5HwY0XkQTBWkh0h7w7g0mIkVeixc6qnvk5+80
V+f381JNqGz7fz6YbajnLfvkijL+M4cfo4cO+Cxu6357EskDQ0MHAF/Juzw+L1wW
tL0xIRVMF6850iHGeAXQ8BSMdq0iqT8TAzrS4EBWRtFiMhusIju8ueakHqfWuFwr
EJKSEONSB4Kc2FQ0f3DHVgx8UXj6I93JHHeRjHxT+J8L3mH3/jp9L6FXYYVcB2vm
14P92UNCA6YYBCptt4fBT/rjgiNCn7aCwsrLobymMqCzkUqoNV/4OnGr8uA72uEu
4QnrszDgBqqaFO8JEhHaRSbqId6LK+xoLjYJq7kw523a3aSU8vKNrrJDIaUADCuX
17aF5ckqiEm3EySA2Q7a3uiHQhE8Rllh27CHeu5B/T15AgBfwdo2oNVwZizA0Qfl
JEKKHn8A53xiTdwOLAa0RVuTa6wna3SXawZjAuptpYEQcnLuXMZrZ6OkvbqzstpQ
IQWnzg991aq8ZVJuI7OVVTaJ5Gz2kMMj+S7GQhn0oUc4n3NqVrj7+3IJbBabHdim
hPK7JjW06uaJ3asploN1IvErBDzhZdPmrILCsqa9Nd26PO2kK234+rygftOAJtoD
NIR4gR5VxCvImIPs6nG+JkEDi4mOcW9e4yvMCuJicrWXWl5OSP1kIincJ6SWjfOW
xPM1zyer9vp1vYj2HJd4LFZHm8AJxxUGy3VYUHejq8UtlxK6xrUQMnJleWl06Nat
WonEUDtfEzv1+yoGd7kV60I2rO+Kkz9epIA2vDPR6PR87PiRFzhu05HnbetmHtiA
mBwYVWKG7Emt9F7HqiBOGWdiy0H37VuJos8+lwuCZLgAxLCgtsh/5Z+yCiLjWN4e
o4bro2JWoVbw2dF2+XaYRXfRA83bxkKyvhU/PHR9RSU1FnZkKsDUBHQgwoz2Qplp
GhQ9U4gokh2XduA0PgKuwHN2sG/dORdXqAt0KKQtFLM4uBSrKQCXZZ6gaYeFuX8v
LagpvPEm3vfgCfnu6TX1GhtrpfP1EB2REMlFBij1EuLWgnRA1M2sQTXqu0S56ZYM
UfkH2C/A1ok9lObHI1pFu5PbI+Dpnm2s4/d7WNVNfvgS2TE4Ly7s3B+PpHmphFrA
LMXmqOYB5ZQn1cF0D43XFLoZx1Yb3Zqkv3h6o3By8mbnKmImbkQQSMpjkUzk+imw
uRlItq6UwRJ0PVYrnAtjhqd6kpSjZyVavm0SQhrU6YBQrs0Z7y+kGWFrLpjde7c8
cSOoyoiRRDkbW7Y4uAmD9uGG0urOylGlDzWryzSMY+DgIpVsL9Utgzj+mtutuarH
914xeU7bvF0hBv1zehTJ2BoRvRnj4u4Kq3Iat3mWj8qDwmOlTERyj6fZZUgrc/tT
B4SVJGZ1zGfSIuipPcCh28b2MfOuZxJUe729aW8u94NahtJyZNS/QW1BFQYfYNk7
zTgY/YEVVAtd52QBJBTwXaW7TbGjJwxHzFoFofZ/PDVktfsP/ceKdtcyekL8xoGS
PIdwcGsFH7kTQfaO9QKZfhscZUwtq9v08PtOK3+oCE8cogWsaoQ+GYcVrNowTS3n
DqWyrrR4IT5LN3xZp3eVKz2iH2Yucf50KUly65/ca285KQ8EwJfp3nAFB4U+nWmt
YCwHn+3ZA0KFfq0z6B7Nk8u06/41jFIL68gcqd0FihOkxqFhULdhHTsRl8i0qDxK
BGDdSsjQZ8X8M/6YjTGKS8a4Rp02vTXDj4GijyjyPxU6WLy5VvDbHzxeKu2Ru4Im
dH+AvyB091m728BuDAPeZsGONI0EtZuEL+e5DxOzb80rWsXEieOhRaKRyaQ4SvTy
fHkPQ4SRLwTJ3IRnSh3sg8I/gjBxetLhgEAnSPaCGoT4TtZHBVOVfuwbfOoHSpb/
bNlRvKY9ycaeK/irbBHc8r+adtfvNIzCy/CFmg+YS+iKgtINsJ4gvXhWHldWUmqj
U87jDYCzjd3vugherMjIv4JPP53PbLS/krv+0qrUvwISgRqG/iBbcXDwwl/3l8fW
ntr5OqjZCW4EpHIUyh8vB+S9UpJe5QBSegbBr7Mn6HH9AZ0Sws6HAsXpI80+g/8a
Sxcmui/L4Mkis7H7Jt+8hw/lMRcHuZcVBJPwugYICmNJSMM7984rJXkWJ2rCOj+u
3t0b7Y+uiLtS+d5UeZaqdf2CQGrNebQvIcoX3jlfTwgNPIUMPqOwAv2fLnR5ovWE
KQe4rulc640RlnxGxMM4fU3ObEKEkl0/dUZ/mkb3LhP72Ec1WPxOg2phvvZRoDjp
xwhPtdrMD6podvC90/VLj9OwXSM7dMg7fygM0u7tg3GmvvxhZtg1dh34O6fiW1mB
HXw54pfgHwAk2F6d7diWGHRJ/QsqAzhd8WHa/jYecYUO6+EKDcSAAmbiAKGQYm3Z
0SdUteiAblUPcjbdzAVOVt0hHEQpg8/7t70dm4mObFCm5XLZoXzBO1WXSj/jbvzh
cPe0vSTy4f74YHVtRTn07YSvOkHK5OmW0WnaHYvRzO6cch8uKtdFaHRpapDxDYQs
PsTIpNccRSl4W1GgnGbz3mDnzC7o9ZAr5Gm7oUDw2B5z4Xq6xBmMUciw4UmozmkS
QTsVWiv+YA3tbhiyFX2xeOfeopXf9WWO4aMk5Q4J+UGukpaSV3TJCpR3pjg27CHQ
PqAIY9efbKhN6s5zzT/TsTAMhPHElMMHTUKjvJEuVm67y3sW0BnIrbHaa0ej6M0y
h6WdfJCY3M+h92g2e0QpVVB9x2sskOBEBrP0HwqZqDcevACZow+gWxfh6Tkxn8vH
rOp2vnE4qtCDrEwXLPcjKwAARZV+nuW4QXN466p85nVexuaXEQTtzFYVHBi2I//R
cQkoqtXYYqrJZtcSlC187pHf3hAqk6iA1ogp/+hqGDOAX8hyFgId3tHdKzmtkV4q
4NM/aK+V3xNbIr2ezKC7N19S183V+Bn1j0wNwWC2GxWwYyJZG8Y3dEfSS1VfJWqv
0qE0s+L603dWL7VhTKo5ehvPcZ6Bvt9SN0idf3J9/KwJnGidIwIkBZ99Bg23Swy/
9dcj6JX7VuGlSps2dpYblvo9qNxEpCR8njZw7Ir2zvfF1GtOXEj5rSaPiFBkr4Pq
mCxyb+laSYPmqzyAdLzRmnlYXLODidwz0T/PpN+9BZnmP9X9nPgqayRFhAk+b5um
6dT1M/tAdRRKjQGUfzpQWfTAfnWD3y0UJJg9CRgu9/LsiKkrOvj+Qs0VMishGMva
Ci1/3vlIjUwAe6BsAlenzAoVJ+qCExT+RcOSxSSx1dLPhWWHUuDpWhJIgCjmgx6Z
VPD4u6qIWQPWfQfVKIvbgjIVpbpy8KjsCAuhJVcCxM3fauX7pgJyuBjEwlAd1Ey4
kCELa/8RhM+yXYbmqUkbW/1cVgyZk2L86vnfLb3jz77437K0iQzZVJK/nv7F9Pnv
7QJiOyxVt+X4MBsnCyG1KcpzULiTfH5ISgmWLR8C6cu35KHZTTYmSJz43bXRaUcJ
V+n/PD+nUrrQ6psktmpYf86B25/T12agBQEvrzZd8QRTmEfNJ48oVkKqLVmq+S+W
+F8/A1OI5d9xzLI9fAEZufeVbj6qqcmgL4ePXhW8mB7YfR1FCevLHcxnZmmLO1OG
mnlRnND7VuV5SphKosITEFvo59GjqlQ+XjQs2P1mm/P2bSxwutN5h/eBNpaRG7eQ
Y3g06k5uDfH51f1yoEvGuXwxRMbXzU5H/wBb50I31QMYIk5o+sjLFOZQUSDugSzi
qchCVFmbB3p80+V1YtOVHhzOolHtOeEkoYlGxL18e8z/DgoR4W4O6XUOMV/FiVnt
peM+7jlWMQbcGC7+1Kq5uRrFCleeMMmqAWlYA+89HTYUXizCGW6Mn6ORjynkLSbL
TT5AlRCeMA6dwv06FhaoWL1Qx6eN9b0npTra5WeZ2hhZKNjLRgJfZI2ciWHMquj7
OQGoB2KAjEzZ9pbVxWyAPYkUSusfovqK++O9faNInOxj8EN68+mNUy0CBYZeg/6d
EUwI257UKQtw/6MlJ7WK97tEULUZmL3z374MM/7EOm/bVxAQs0ZlseJIHXdBqBD6
VMW2JVK4lccO/jLnJPRvLeqp4FZiFOyplZEKJaM2UefHSbDdtDdhnX81GQr2vN4O
ScSdruhgQ+vO70CMNzwdb/kYpPKYToNADP48wiDQb+APHrG6E+jqk2eSeOTa/Syt
Nv0+z8xU0x8byUlayVC6Ezm9pxckQ6czSnPn6iCV5VFhihn6eSZLjzDgJWKdnIuS
1+1dqVmI3thA40ahFomn6lf1OVbiQEFbakLahB6ZWTTXx1BZxDuQ0cqQShLPzT0V
wvwucK5Q1adTBwVGoZiyUNghoyLR85kpG7OkDO70DyAvu4WySFi9uzqhNGMOWyGQ
HwaMD4rUrlu/Zgo98UlVh3MR9tVWSpEb1GqgPZV9GFMw4e6DjuEBnysIZWCD24jX
LkOTwjMp1X97rdRQz2asKd7DYf4d2I80L/Sk32davGwYw/UdifniCkaFL/T9IZgw
yXvbQVSjsBJ0gTatMW4hirtIAyLp5TGQ0c3iwLb5KM7B6UQG7JP7YvKHpNcAr8ch
MLO5OY3K8QvaCwIXwfXp4CD+8aiQOb2XR1x8Um5qBID77V5Kzn4c4ng21vrH6ZD1
UnJRXIGjqHoc/j1OzRNVnQVfSNY7AGYG0w6YyBeyBhsnXU7nsZ4PXs4KGISCfi+I
7+9Wd1dJ4SPeeBUPBa+UYNsVLJ9xgXhrmVcpSHR6+w9tuWR7xcBrU1fWkFw1MefA
8ln8Dwps+6tZcaGc9dUOSpL5fxFKhGoaU+fpGemYslIg5HU1uSKSj/6yHlrZyXZ+
atY9ORZrNvRTAkOVrCp7RqL5z4AX7ylzxSKU7lwRbqEZZqGji19/5Yg5mJmrKLuG
kRkv4Z934lXglbK17Fw0XYNAkUKM9t+OWc0npyll8tSSuy7fvwcV2DEJPMDW2Isl
N/VxTecAjHANeanRll0verlh2wJWiEORPru5YSLLpc/CdT80MAV5wt13j+psnSFu
fUAn+l6zp51DNgef3Pk0pbDUwhzALjWZvcoFGmCmGw8Bg2gr7fgtmxk0o97i+J4m
5U2fS9J8Q12r4w4PLdgEiazAaAT7jXAcA1U7xRSOCshxL1FvUPNn94VdaCLLLwen
5stG8SW3/xnDqurPIRPdjXGgTPmrgnptLVBcd4dLVqCNVY3nVbhpax9AultMUNj7
ujYKDkTGo3wgiYqDWAA+M3dG6UBOxIetOGi8xEGJhT1SJdqqh0oOlK4Emwb1H3nU
Du5OcMqmlP/OM9KvNv9GbGGWvaoHV6yN//d4Am565acRyxTiInRSQ9IhBtbcHQ2y
oNVB1Lo0PSM+Zoo2aI0mYMaX4LkhaVRitthVR6BztR6uZQ3UTjq4KXxDJWz25yGa
S/bU45QlvZaPPMDD3ucin8zEhipZPcvNpohfi7UKf2V8TTZIKTAMLLcxbUUbuBKG
zkW2h8Oqsk1yl+sjainjrMB6tYW5ZYPGHsmQwQ7MWRCrLyjqJfs+OY1jjjHZVrOE
+8iXB4J0+XeFuXjSV08N2DBONUj96j5cHYcOGvGlnJMaYiXbMBlAOmvLtyg72Dor
6gtiB2BIGgTShIrVddEEXcF9ZYgTqCOJk8y98kfv+yvXgTsxnbMgq/DQ89YgnB48
So41K6yTEUH4YdmSfutptuQxtpGNhOXNfQgyI7KH8JOX6z5aMjB435+5IqbBmtcv
wLmKuiYUae696A7eYgasM3QxyKI4KCryflbCwnLXT8QKi4OltKQrxK54XKNQBk2b
6PhicvS+cbHLdhyceXXknT6dzFaefOKLrCNhG3ex9qMUszmBQ+7cRJ/84qYuW6wP
rJgbnQpno5u4KZjhxOSgulEA9yVVI7SkpiIVm0/FqGHmKNQYwErOJb3KWjy1C2X4
fiGbaOxFOZx6D+tVYcDtecPBDvhnQbYIa+zzQKuVbSBxD4vh7Gwi30k11Lofqh8Y
ZFCn3k6Psz4F4y3wrfbvgTbEaZecd80+W2LIwkzyYaj7h9+Bl6m9BrHFsVUaG5di
8BgmnPdsiF7FCqeqyzmPzc1hAemWWoeKLGCZbrhtMllOMf2Y0zLzZpU+c2bBzorj
mZc/nHF5jjpMrgpJsTcLg7PB11R0/CU9QxqlI6F+/eVLk+p36mUNa99ktbT/anmf
04qkKyt2gk7LyIzRn0EgkhTtq3Ktv27X23qqX4QNJVBV+19uJXUZrx6SCd7qxb39
YZ2p3ivwRod1rNkO/7ZizENUcKpicWtgOKD9NgQNeFexaWHZ/cgcomalk0fAXt9X
Jctw/LQc7lCcdFdicImm2H1ApuN7fOU3clVLRVfiOxTPfSB6oCWVpEJJ2avIhL2n
CNgDYaZ1Z2w6/phayrceVT+/IX8uxTxULmXguwxuwKf0JjgHoeR+D9XhmmMOiSh2
G3Lz1Q3ZMRF2DtGTFiAB8hyogpFYaeWFch1h1sEYVgK3p0eMnNzXLzOHLixVUHHT
3yB+lCt5DDEJDsMp3wdaWnTADOwBtnepZsGmfdYa1vjXs7fnpSUn3eeQidr385Lg
I3dTqFhE/MfB4aNg4gXKVLS0h0Q7sCqwrxQCr+1DqsJcKOWFY8bohChqY/dF+cix
j85yfPaId3iczC9p347q4Ub6V1HrZnYnNwv1YEsLWOZlu/s3BUQX0fur3XlBNPRz
P05ZfpctLFwgV1bEuHACAqYk8XN8yb+AKpssUlhw212YgSTAl2FnFr8Us88kkB/j
As7NibjQIO/VUb/TrZEPUx118PS2SQVl2r2Mi2fSTE1+qRrTaQCX9/9uUqG2Vw+E
bcko0rLb/hLlacc1VNVuWmyewcJDWNWYBLmCJAb/D6nGybazZW8CtDikHIposqD0
QvX1cOaMfp3da9W/i0N/ZPx8DWPivx26APPWO/SLKW6hpXWGBTMGW0U0QBUHlY6o
lCDzUG9b8/cdj6q2e61M5RTfvBtaEYzxsuV5cB7CndeCBavfigW39kB/uBvQfwyM
bVBxC3OVHHn4psujSMBzsnbCs3jotQoTZKZZKyYbhnlsSfUUKbkPg7Qj8mh+f5t/
WUuja28nkig/alwViaOzMmc7E/xCkO4Oepe4BYByCxGrSHw9W6QAHLQifA/gHj0L
tpi59MPSu9ON8wESI/r38BydNrR8kI0NHgZJL6K7Yo9M1XkQasuuhvC58ZBiGVUf
E+Bqdcfs5SYnyGejMZUI0NArn3JZ5Dptvu+kEsve5LlcxxZQvq4yRJBITxSa3e6U
SM3gQwnMQa6SPgF7JsFxFmKW9eKpK4FPeCcDnYRAgPoAugAxjvJdpuFOwFrkab43
cXuilqcBmTVBiFmnGb6xoFz8nNU92OqwhUjAaJq0wI2mh1JVJXLdqiUtZrBa3dte
l4bVQ/CelbNJkPoVLOmo+LcTAsYLyhuAUI9gITzHiKdW6r/zIOzH9sjqvOk+NG4+
SED8UFHMUysd+p/rir3tfDwTtI5deYFXRoYBAJmCntPdPSFXHZH32SdC1tF3yzhU
A58FlVPVLNEyshv28bUP0bxGhVyrG9s0KYnjklJF9Q7PyMJDVJ4SFg6l7ZeJ5dT9
uNuzsZECvzz5EUJzNzURO7GcGBB5FKd+De7gLXe9ESKxZPFAJt/klVPT0W772t0H
QC7mRCIvKrs7H7wduZ693hFXQZrwNtxC26YCO9tW/Qx1a/OVtcOT4gy1pnInuMTU
qOcwvzBnZA6weUv6oezGugmE1pJjl7SGZrap3eZLjflwuOJZDPqpYndKpXFzuNtY
YkA2ZBWg97VnTaD4gNDqKYOKlWBgjxeVkvlDRYQ4egWjDHTE0sP9skAFc8CZkxHW
3jx61DT/Ven0n/DUkQCv2jTERIEmM9+pqdxg03BCnw2MKoKkTJMxUSdcyTDYdWLd
bkuM+FeAlJ+bA9O9ttcl1rO/vyj3MVof/66UsbTF21mUN97fgkO0UJHVoMBnOLod
qDhhw0eyX1tGv9lCk7EMPwsOUDRmar4us3D0XyL2Io5jRR1q1uVBZ9xCYY1+WqSb
Z3oJTKKeE6ZyVSSTxhDCLzRWo+njQ/TCWg93xpzCDK7kNZnPATbhNoPoUFw9Hgc7
3qbyZ7g3OsfoRpzaR5TDh4lJuI9Ss2a9gZNrDmJwJC4AjYpQuSpv8lAM5iayV9ft
UGWGfd5pYay6CvrbLGHNfKNGOdYojw2VRpKZZPnC0YDA72mGp9Fe5JeuopZrbdOl
ftLy2/DGL7JAvnSOrMxC3s+IOQ3e5rCC1y4J4zEk8SQs4doxHcwlUSz7v92Xkgkw
OllAw6kNZLTHGy8MVH1UnoNItR8BHci+QHkW+S+7s88G8Wcw2y3mywkDE4J7MHWp
a1VkwFLi9aMASTmmu5CQwQaCY6BD+sZsdLMHY3R2JP4qr4eJPx7GSIDErOpAEYUK
/1JCn5qDvsouDhKHaQoLXaZc4HMWwtyF5gFIR0peptPpaNB4MM4ROhLEH3lyWJ6m
NZe0QhGt9hv2J/7sWXg9UnkCfE1gmdZL2UQGhrBiQqkGWTNuMJuvMtqx1162YA8i
DWSZanliBRy64WqvNGRJW9aJbZgJ/i4jrM8fibjyNLlo0MeK6axWxeQRW9SW9s+2
3R0b6XTrLLsjZcDKgatiBNUVTxF28gxnU/mDgvf15fSxUGJUF/6OlJ9Q4g6gYsii
b2GyNqy9PTj4v/8YNFAepiS2vtdcENuZqZZBaTHVaiKZnqxUVoMt76R9qZ90QEIL
L7XsNbKrQx8aiCshigzyIt88ybD7bMXqKjHnX26LGD1IezXKXO4Kxv8YTYWYR7Y+
wmCtitUsFS0HZTYlvmIxZluC1NIyps4pPGQ21t1M3NlQTqL+gkoKzsryDM5M4G20
A3NXjW9X1opKsqfp9mt3QIXSNhudWPjtyz5kz6mq7hZUAp6pLPaK97NIdvN6afNe
ssh8ch3kSXTptzQdt/JRhqXOXcHOF+KUAjbw7wQ4NIVll72FMVCC5IHCxOoncvrc
m6CEcpp8tWTLiY6TeVdGCyWOQlYGv9UYleLiWTNjhrCxhQUhkSCnAfEt+U/toQaw
NPObWwm5VlcGcJ4eKvKFWqfahNIZBSDj3B33WNCeF+2lwpZfrjKGJFpHzZrZZGcG
r5pL6E60F+WPLPScxx937lQWtz2x61LoF+FAEIeGEcVF7qYUdML0mlpDxgQgzKE7
yMjfavxsE9W36WfhN/7LzLtMv0wzqg1qFCmWn3pCZUl9eSW7m7OZImcHCsEj7WNO
ZuySyS4P2uklqk83tOiprUmSldcy88x0DfdIZzhW/hNJFepJi4UAbm4SEcpf+5dB
qOnD/mXeuk8INF4ce295BK2Y8pCj1a4xBa9Nu+vBWG+E5l3ddWuB4MUJPnXdctxN
KoDFu+ZI/OneIsYOOyNHJlTy6Xrg8TbOP3ZVlx4DwlpMaNisH4leDWRPmoMfONFI
kOs9XCZjDM8q6EFTUKb1nPzbBdNnWJ5Q0Mhq2f6I5c0niH5KKLwqiV9oFLZ3vUz8
IvmGvjGXW7YrENdCNQ73Gdghn9nes9FfzEeGFnh08CFs+vHe5YJVPlqYkhvKgAw2
eg4TgftGdsPZ/3XIa0XH0Q/SzJagcsIYaF0Sk41x8syX4GdH05z7Efre6upQRBCp
uiTkVen5z4w+nqdEW7H681e3os5i4jPUw4jzFFdrzpfTlwhiginKwY089lFECyXa
JMmbr8EWJOQG4Zs/tTL2caJKVHZIm+Ixtis/771hxbi3PzdBjC/uBsuzBYXr3ng7
J0FfcOWjay0TaNDLcSDExHZvU3NCi6UUXcUaHbNAUnROwx7g3WcwR3UI+rh7BBqH
lUOM2Ew8cI4yyHimX6p5EWHbWHgkLJUIYDnYixI/TNqqDelEE8qNitZ0n2ECkkLr
y50kHhL0ueQctduLLn+TWw/dSrGFeP4ebxOe9fR990nwDTy1CHxCoszu8cWxIgki
6DTISDAHc89d61dQVNmchbrJ3eKvNus1zKYSg5m9gwUDCfpGyylx3WBPQxDBu60H
xhKi8QxGN1qIHZiseXKMi0zfIKTn0VEBlkzGi9TFPHD4xY4QVvN3w6bn502RByia
fw0t01KFaspNqBlIqU3h7CPbGen82D3hIi+yD18VKQtnwN515MGPXm/4fUAdWjxu
LgFv9j5VKg6h44MvTCBK0nDptyEbXEI/n/GS1BUo4ThIzDlgdJugeu6cmlIkJQXG
Yeistva8ZPmTzIyY5QJy7dCXDnuwPanOGbyQW27F+7rlA0TJkwg8YsJhHRfCz2on
fQv0sp0E2aUELqUzyQPztxekpHlXCu8HeWoaxNGKiJOHza7dxNE4eAE29736B7jQ
0eo4sYGOWkMrcqMygsqrNCEIqc2VivyGtJmmW1ptoUAuTCUPzeQ1z8KC6Mu+X3ry
2Yst/ugxDHmlzzZNe7T5f5NI3oanLDbEszEuwTPC41/h+4M0npQPeDp76oFBRPEk
vEINXUMXZADfaQDzM/XhPEmMFubZTgHysjyAYZeGwT241bVPK+ZQyMNq2S5UiOwU
+xkYjHc/FMbsWO5EYKcoTCgFkqR6z4ltL/R7q5C9CaiiCUefgkeEiwQjSErjp3y6
l3/z0olYetlrdszVWm17PaRlbUmj+ivR+fTaYRiZmUg8iT60yWmnn6MgRmPHluKU
ciNsqQD+VN5HTnrd0HwFmRx7SPUZTfuTKrkj0d2Ld9d0OchNLLbxk/yw1piqq+nl
0QOOHF/oNrpDfDB+5/1NEpYLS8Ozh6XAsZH/z5YUFaO9CaRB4TjAwuqTUy2tzi6s
dT1BG1GOzztSefjtuWpkcPNttKlo2KVTNOzOLybTNPZUm03TvvdlTF3vM7JyHWOk
piBxrwLa+Y30fAVMktrzjEAVJIMTl5Ylpx3baqXrNYhK6cDk94v8FQv3fxlPu3SV
1W4WIweOcw5pw2KZREkH6ESW0tlT2F0o7t9d6J3s5DImRDTjINhewm7RDvjAsqDR
TDvfSE4Tafr8A9qwBQFP1IAKCccVm2vFKhhWs4taFIwu91TiL9WMQ2YnwBibhuXF
jgK/dfzOSt3Al5K2s/PLri1hCC9tZFhCZNla051IO8p4uYI+AnKjasQ1NfszWOjw
4mCmMIIYgxF/0ab5vnrvTo1t6ulWwzg/UWd50ZsfX7Hn2ucAPxD5ZqTluGO+pAvo
EsuZPsG25vKNYSLto6qMgKBE2Wdi9bvSVlRDze1vWvG7hvrbQiJx+L92ojbU7QnD
yAFlgg/cDtpqdzjVy7wd8f3mX+i2SqZIo22gQRm7T2/k2JNFe+noE72U2CiLtwHl
VSRB0K/xNSDdOa+SdKSpmtOjoUFNvkm67YDzFlDSUrmofFZndvTnhsGnC8GxF370
YWBv+sfrngtvqUfk1w2zSStDNfU+EUobCSEnfmPpvvhDL/rL1XLS123l33YwpTN1
ydi52whFkfEe3LuH9rYz2M0T1xk5zOHDPvkXz7eRUOUT1zJmPkYcG0QLmEI+mYYX
NesHCNhgaTscPdfevWTmi5g4ECUzEj/5AqDF7MOloxKXXelYqLP0bd51rc+VQEVI
BtohTfLiXr4K0RhIEnt7L4wSmYIrvRq3AIGLpY7knMQd/oeaFu9FN0slakc5l3aD
49Zn6OZ0YM3u9cUidp1hvCNJZ6z1sdvCIuxuHbwVfuOOHw9jMSwBc9zJi+0YwJ3n
fpOUK5/7a631zzDvoP+F8AqBejpE32Ii2RE1ycPxD1ztysZvZYXxslaneRfNOMNl
y+gRPUjwFaTeROO2EyZTMr5w6xa/OYx9A+IcnU8oFPA099fdhyicfDntF9EHVN8a
QovkjpmqQVuYh2llOEFegHXG1DrjoxZFhEOn16E+1yJFaGD3ielH+5IcQ/8LrFbQ
4uAjeWDV8QK3p62mYgwK11i5aBvAgBSGBCTpyH0mG6VJMjnczMzhmP3upuPuyIqR
/0k3ESjveDUHkmlApZ1IEU5czVG7+vMbyKyzqC+Kayhp04p1R9sD1LYNS6YCaO1E
Ohx7OCYOp3EZD+cQaATZDqYqO+N4gXdE53fmSjjMsoimGFHSM9sUAtIhxA+3l9qq
TrFKmyrmPwUExtmXgOLEGySQCTPt8gKZlRDvJmnkZrgcAJJ/juJGrcSnTQvuiMmK
ByXxG8iI13oLtcoIMJ8WVgtjyUhK+CCyyhCzNt+5AbtN4BTFJcgOhzG1IxP/jHsN
T8l4vlRcgKVKZ2YceTCPHNO8NAnwDZXSRPX7gpyGJr2+AyC1TbApKyCsHXvcqovW
nUMhxZ6saNKteBMVCR6iX3zOwKgjNAndNsxIp/T8laFM2Haduve7zSybj2qXUiDH
nI59uF1Zj5O0ya8yNybIvBtZI6DkfoeOByuS36rN/6oRtL3ZxM7M1cZj1T40fyQl
MsQgMVzCWlpbEIa3l7HSFVQF74Wxt2Y4iw0ToJoA76vzDJstJvM16EnVDvQ7e03o
8E2Sr4fVKlE0DqeA+fu88RzvD84T9CBXIFzmqlcThG8G0DgaXVV9PauRu2S4pFT0
GWbREPaWmFrta+rl2GbtJUgrsaEzrKo8nqUAPMLTQ6puSen/T8aycyeAiWmjd5I8
mjfsPQub9ZgIxG13KAviBmj4/nBDAZ43/LQUPZC3T3uSL2in5Eleva3CNmzPc8Go
psX3BIi2TvUfBJe5j1okCxNF5dVUJYcrp1C5InaUIc5GInBrfznN5xDwgQ1KZqBt
NR8hEGzHYMCbKMCRS/WjSjLe4g8Ves1n12JTOrdUBLyvbvcf/H2Op2reMENnlHno
KUhmEqM4dcdqxHnYGBOfr9VTgz0zsSkCRcKeh4QBZpktPoGjAm29KVxihO9Gfkkc
x0zvsKIUYqURqc5mP2Dro1YpzX14UrZbHcVmD7M+ux79HB63CTfsCQHAEXJ+lar2
aWHhy5H/lxZmim5gugb+WB868aghi+FfNOv1o3i84qh+8Mp4uFyYwUMkd0o2TsiL
1VasrT7BEfW/fbEQWueDGVECeYVE+Bg8whaIsuVoH8SuZMKiyhJFRLtTEwrJgQPs
uCuDrbY4hk7u006jkRtG9zsr3Pk+mfsztdggLNOwrgbSZYde88dSEcXpXKzjBkUO
zW067CippljkxeYq16Su3moQpKgdytstdZb7yFKiabCmc5iLrp0NObN3DiE+EW59
Cx9JuqrH9hUWW4IzbTXXQ7CTxCzR97gHimzEG5Mjx9MMOEkXRUv2de1i0QkumYdN
wTb0FbLXMDBSmFSmzSTGoRztDducrGv991dkVFASPHjcMZ8Gd/WvKSe4Ja484qhI
6JOOeLTIeNTd4s4kdKGtrX1eDpBVbYCQ6fVmiAQ8cmA54zamlQoJAFx1NVSObtPR
WqOw/+iuiP2dIu16RjbS6MLCTLBeWJFsQ7Azkw/OdCJ7nL50MyI0iLcgnwEHPtK4
CPyyxekdKDgBkW22nNpeighOtwycpFuNkhnK2zJZAxJ6pykMricyUoHgVfERJqYZ
egaL6tZpSX4oFqALgEfI/XP795trtj+tGTG0qnTZX5E2QDZ5fVIJbxSwGGd5oYyC
6bAIKo0zYHi9Idce0Zxo50MUpnx48MieU5UDBp790CzzLkxqPhl3hmieQEdArpS0
qLB3qursk9hyI3JFFTZhARBiknlGrzwJ2ITIQ7P4Mj5ijhtd3Ft9osByhhm5ML/S
xqrXCRSwgWr9qj9vVIPXmVdhyJBAy50DeRs2tWTNg+i9GkM9+ZrEOGmVhA2eGKK5
uH1fCxHbDuI/6A+sT6ncl33aJ9fkzJsXJzNiO9HObm4utuTpYxcQLdObgntglL5u
iq7vQpyr2N32B/3qxQgtAi5gcixcUIcP+d5tCpKzJnKIDonGp5iViEDdS3ECRiVq
2nLgG+522cS1pL28nUDkW+YX7Fjxp/45zIzpEA6mvjHO2ufi9dH1Rm6TOTKi774n
CE4tE9SaCIPIBs0mKSoKtxfX4p77NyHJFleCtV6ZIy3M2Urq+XeXER7JADExtX4X
F5hZ6lDeayfCn0ZbyY+ZqDFIOrZmzT6eASPgo0irPs0/QmboyuuIp/5n5WBbiR/B
mhyK+YROkwF8h8TjB/JUEk9epyK9bsCjdNIIfFKdKofdSyFmA3IqBgvaKTzcloWm
QZHKSjR2QYmNrtXDtN3A9G5LKVpi+3wmh6QUlL5/5ZKek8NFQrzgT4elP/i3aSrc
Xr3U+BaSFWonIe4uHg3RljQ+9j164jXRtNaKhhlGa7UV5NMCGrmwyvSYRl4wFpK0
576H7YJnIRtCBiG78gA0NpgS1wi3i38nlcU78qZ799dYtnBmU5Qe79chHkL5J6C6
Usr6QnczNrdg3g2cjlYOQuHcg/UokvrxzYED1sZlAOZApwQ7jXQwkoP86pcW/lAI
1vKjHIkw8RtO3+O0jOCz6sfUoczTYt2pIKtcOOMsbx9BhwMU+AuW1M0RwNMd4Kzb
VD07gNVngFzhi+ETasLa3xmdTAX+0zidI6LMbpLljDWOShJv7uTTdp6H3x4rVHuz
Cc+QWBi8ClMwDZDDxFtyx0DI56IbHFr8xpzm+gtY6dzhKdGGRnxqEqP80B2ENN+g
i233HAdqN+spEAXH/k6C9iCSnU9J9+1+fveHwVB2uwg+URARji0YwiZcnor9xioS
eDxG8Sebg3oLFxqeeGu9zUejO+rRiBk79bEnMwLXjkavXsPpzLnvmrU2bzTQMK7a
eUdy4k9b3UtaHRay5DA/t7Ajt/UJkZu0LxjOIT6IllpiEHNwqkaWs2WuQTPbcJO+
geUxHkbYHNxGO2m/LnSVuhplZIDB3fbblofVN5Yl6uQAUvDtmvtAcUtw9V8NdGSJ
ueHLsavUeGC3vnY/fGIrBpDKybC14YjIuvu3y33nYANPfcBBVVJm9aG/qblBejYm
8pMEwIOb54IgNGe2X9Tpf+GMh/1E7Jz/xlxp5LhuT6zhvrlIuKvwr2qs2dR9kqfK
sXkyRqXkP9QwHNGfiEhwy+dXoeSk9/0vvAs+HwWI99dO5y3Dj/m30xbJd96bkF5t
pNMHpBP1HQmS3I5b6BHnzvcSbwA+ox1KBdLaTwe2RBQ3nn49lS1pZKk7Kbzj3lBh
f0NeXtztUZhO2cBYO5sE1JxSztRumbv+kt7J5cbMnPmmPQVeLtrgo9BA6DIXtpFy
5EVmT2CqwHB3yPNNrEY5ip2qiv6qsZa1pEUqLIMPVoOIh8WaJSIWooL1DmrKBsWq
W5Y2UJJcAHk9LAcA+jEw1uNOnhKnUKzqmxmddjiPAWqf8tSIEB+NCV6ty+dMA6bn
58zGOoQKCmCLL3QSsy7pa6Yl6HuGmrHzf2HCymdyxvaqHRXYRzbtp0TgSWcU/Zb5
JMujomfOxH8qKDWUZsGSzyjj2+BJRBIV9JrRNKoJ2ToRskM7cdLUuLqTS7azONpa
Zxcmv94TvGWw8zT5godPj2S13GRSgwAbytu4yqZRf/tZr97++iX1xtQXGfLZsBpu
iEdlR7XkkleGiK0q73sZK073gQOND5X8ks+e/LTNMFEUxS4ywByPXZCZEnrFtLYj
Vd7mOgrWoiZOT+c0YwwCh2Ukc/ByZgzDFotPnGbXLBk8R1AXcmCQYEmLzXPdj6Tv
BjoAPXMyKxHzdhS0dXkino3tYyjaWxjuO4HNZp/IUzJw1nTVdGykevf9NrDT1sZo
W+Xbx5jEtYXoQXVfqPmK/RXonwCvmeZs2+EPbTKpVLXJOf9r85dgrpWClnC9Fkqn
dgjbbzRpWBmJWWQ359zgtxlVjYGptPad1d1kUNMZBPDzJwsJJNO+iAOQeCHXDrFn
IfErl2JPPyTU5A72MM/fS+7EW4GKEJXRfXQyJtCAsEKboKozW438GOO/q+oV73z0
ssVjgdBSg30H5WWXyZUIKMzVjBlhpWhgF2FEAPnsJQfLTRsIbzfR8rhxDuhpTazs
kgiXda5jdhAGcWGbrYEvJUhl/vD55fkHKpDFSIlSCl1KHMA6KT7G4rhF1bgywWl6
b0nw/m6YzjbKsutTLKSSaMwR6WyBseIMtbvrEt/Cb6vitQ1Ky/qSqUfwdIYvaa2r
lSjvHRgQHMmhZiTakW1FG4ba28qnyEzzGd+bMj558P2Ri42Q/idp8K3vU9KHF6Kc
6P8RpEUMK6Jj3EGGX5/zLtIWTSD5jdm8vvxG5KToPan7Q/DEIAEcD4sPRTTsPCIw
y6sb/BvZgxRS5KrejbgAfXeWDvcMtu+PUqDjxnhanz7nWpm8q/+BgGlyGKikk88s
uLHgPvNessRzpOtNXjoJlkvqnG+5TlFU3rsCJo7dR30wxRxp9PBQAvWmelSDwMKD
PZbhWjXTc+gzHU1OJ1RqtvSSXYoOe+6KacbgiAt1pAL0Zv6rVmBY4++ZcKtkLfPu
6zZWEyxUQ4VcShwL3S+tL2XFoxo5dyPz1EprR8rC8yJYqXL7ck9fMHgfC3Iw3clr
GHddEpzMuHqPYW0h/0JPW6ARYFk9fGHpFBcf/vYp5wakMfNYxesR58VZ/1+gVfvC
pPqCfASxRcuaFjGQ8esJFip/M/OSiWBw+SwFvNLbPF+CkJuzQuX8C4pAWCSVHnkJ
1/PcJsW08THUgoHqkND9aq6UvV244erDu8oFwAW71qEXi7nQSLNO3mrULHh+OOWc
B2KVqvQtLvEVmBllhjuoZe3GBwmFFl6uo7zJvKxWy4BEMI04y1d5oY//zCOrswJQ
8xBP5hh8xqnPQNkDuyoc3U2d9chiv6UuPrWmmSFb/XqlCy6UUSmMhhsWFzn84Q1y
PiX3MxvaZAtzfBAUw+ytLGQTEfUejpedzzjbZvYeDdlIQD1E1/LvrGUt3dsKFvsN
k60c1wd3oj6qy4PjnaF5TbiGn/4bom030+Ekd/0F+xNyq76aPd+AXelISGmnz5Y+
tjJ+WgZx0s4xf+QNQIUb/nlwt4bA/PYc4v6JTx24kP/83+aiHaqiGCeK7X4kDog2
m1H34huT3BwrmRH0o8/KteCBj47xeT3tDnPbFDZ8A+nKrXa4QBScMXzOLcZ2i8Oy
0OccqEGX6/neJsLQ50Y+psBA6y1TKhj3oxQvGetMcEj+O2B6IrZ8KduJD2CZc0Hn
/e0Ks390l2x0HtViHZrXn0Ett2oz93/SRwvzAfp1Gvgqakb30yP+haniWdcHuYBx
g8qsr3qZK3j3+vE5fsoIeMVXRKGOrlaS9CrvJNWD5OA0DMacIMQuag0i2XmlLGwn
UvNkIctpMKt7XBnwRXrl01IyaJ1PjNVaWxbzSGWWUqqvNsvUl2CqWaNsWqp0oRSt
Il50zh49WqjYtn4KrqhYJhflXM/Nug1ZhjmMo2kk7rBbk6fvmRFTV6xYnz+SmZVd
6OZiCtrKAhVGOlL+QzwF1D9MtJKsbLARh2r2OHYPYsV4eG87hcmVKgNfER1WUjBz
5CyW1eXjhjIDh/wTaDSuoJHvZVlACjj655BU6bU9zQ39Y83/soP1w8cOeldIXIAv
woRdOY8Z3NH6fA86Y4fgzc9G532cQtGzF8ZEnJYglu72v8h54CXbEWnN7Pxcea0k
YlhI+B9BWH8OgQ9hstVbx4fVsLSOKdslYCKJ3MCsWRry7A+tl2LWgD7IPqOEK+Bz
zXaLzN6m6YP3xtWKz4u+JCmDWWAfNqCdSyAiKVr6rdBOgeXF02u6ETI1GLqkd2wq
u4I6lQCA03f437LKRhQLSL0qK6J+wjHtUlaH6/9ZsV7ffWkesb3/0fKuMpBrp8bo
jse1knyboLgHJ9oa8u7WuqTu12jbVSOo4OHhqFqtRZROsupLo82vH7wsEh2me4fV
ucYpYpF+z8udCR7RRcJ7JZak9yACAJwNfURuKL7ZJ1XyyymX18Y2aJR+H5cbv787
xn0x2kvYWWiDCSbFelBrZhFHVXc4/g0kvcsHHEszALP4VWJlQt74MJgjt6RXdKtK
WXHJtTsV3H6oP3P6ogjx2JO42CYvd09TT8DfEugc2txIBipG9dNKdjd/LQV1lRhQ
CvheiMPrs1V0muMnkHx1mzA/kbSson0Uu6My9lsoWgcho7dGGwRaJjJDfNitocaC
TILCPnQrAJoFGuN/Km2Pd6DkqZCD3itByVPU5Mf02DG8J2XfbmoMKzeq0ewD4ggN
5EMLmEQNf8EyeKY+uVNyfGiZ5oCMOgNHPVzZFsYjDwGP6Ym8gcxxqCS4bH5aFKA4
y4f1RRS0kO+g4SENTHGGYiSMEVxRQJSgvwFGsdUmf+76EDgr8jIhrWyoqWWWATKY
6KCiPyiCmwpJInr3sDSFMo4h292OdmigsM/f7S05B7LFQrgEYLRXZJ+QWM3o8dFF
IgG8YUKUkSIwFk2hE5nD5UnmrdYeNaypN6et6tjxdki75DaKXdy+6Er9z4rtDiaD
6J+q/TzLekqQ6zwmS5O01dXFhsJnNprEW+Va2S3BkY+JXkh/mhnyRyEN6tN/CNo+
GMFEmlXRkPpbIzbbj9xRLix3Qbz7ATI5oMOoS1YPEoJYR/E5eMa6TLXwxv7EK5D2
FzYXxYaaKQCaWE42HobtUky5o5387s2HPxFryFkSPeN9VHkHMSMqt24RN9r8bp9d
wniyPP3ISVrH2rEl3F9biQCI/0t+tDcWVtZ0KwE/uj7dr0Bib9xW2GTKY3rm7AKd
x72/NsgNGzF7uzjHcf6+JEbUMqkJCQft1jYAyh+CIewy7IT1wNSep5QhXoZZ/Dsc
w//xtZ58fMbqvv5PiziNxbU2Wb8j5k7qmR2N9ulQZa0HcjR3zkZPWbEWgSRO0LVg
1LnxnRaVvkYkeN2/ai5JAPc1RavkBFhx4dV912X917TYAxEOeSRgDHT2ievZt5lZ
U2rVkQCNRtsvcu1IHohGNtk+TaXGaojrXyVjN/BXk4z8RZb4kUSvI+PbboXiOh/S
vTgDdUkFh3V8Y18znts3BjdxYQMqJhTxyp2KUx2KP/ilge5x8Wx5db51yegrUti8
fv8njEcNAX3YJbkGcs6iZN89hxkSWXcG8qwA02+NcRvBr8px3Nl9w8rISRB8OUjp
q6cvaAXhFHZJw8Tho1pKBejcXP4NzZmluHHr50m0u4o+4WsSFCsI3t59dTJ4oGqH
/k6zrkRRH8C2OgLdz9iwe+8kpWILMzK5k3DJ0CeyksTgMDLEFz5jjD0yK7h+M37I
oNgunMrbZql5gIT+ZjDnkljcm+GdvubZf89HHUwR3oSduhJfp5YqOXaa7UdRlv2k
689PntAaOJTL5LhQD3xTENbiG5Kr9E9P33k+JUhDfOD7ZCLkgbBJHYIQBb6i+ysQ
OiBXAU9crVSCIhRcvDpE1cRhr3HNoGDXYZeO9nG0w+k9v8BRf6a1z54XzROdgXTC
ArdjYawspOjd42UOVSMAXxKydVYTdiD6LAnBBIq/wnGhpyK5txX25EkjvzTdrP0C
RARey5TBoukf9PkZem2w8o8sksK1dH7umZuHUdgEa1dOgZtGl8OT8aW195tFQsG+
i56NkrFDyBhHL+8iGMGbeTyqBYujzTdruD8cCSGjxQNzZlYiXhLNBQJWULwObChu
L2BHPTlylpl5ErXjkwFVxRWTXEW8A0yM1BfToKM+NTsnnLSwoZMGv0w4lm70oFk2
STtTmxl72paAnqUCHoEVzJ2XcxIt0IPXaQ7CQDbeukT4kRiZHciXJW+ujvxbzB93
kTbkD3ttabsb8ge0ZjMrX8fZvyhIkoV6o3zAif5sLJFeo+1RVa+mq2DKn0qyx2xN
GCIUhVEUVEIi7nbJp/RN9EJyGDOS5Vrs6czZ6D5tbwaJmBJUW49Mtr14w+biMHwo
TJK+G1r2874SjAf9vJnna77OPwbFLisAtuUk9MWtG0exBghnj/cg/jyzGzRzoM1a
OS6oDGOI+bMF3gL/Y2dMW0l4nQIMSjyxW2nK4fAomIhQVJd+yB/qqCCXTGWSLog1
eXfHzp0RIGI4KofBwIYUkhphHQPTr9sHP751AkexpkDd8c4ZGjDHjlBBieKmk0kE
JcLi05OBtdDKUJrqCiN1KXN5vkSULDt6hUb2cuBUrmoTKxhC7JlZLml43rSRM+9X
mT50uW3SFh3bqIJvbx++ytiSmDZ3wASFeAHJ8Y0uhWaz932RRc8kJwJMaJ1o+3SF
yMilgW3iDoaeuo5LwJjxcC3unfFQDRyUQp59rV0icY9Lz9URgKzF2sYQkhPWfvM3
oXsf0HsORRMUvFmNkHBpyz3RBQLfUyeI5FJSHm3mvlpdUMSWXIWH+PQ7Rg1l9wif
UzW8Z9bru1J/VUUC6+6ezLqQpdMKgu+6a2tKg86iBxP6MG7tSeabKHPrBHgvwmjt
NgrPxr7HL/iokUjpI/8CxTepcH1PN2SfV5Q7gHw2tU/tDA8n90pjMzV2apgiWj0d
7wnqGM616Az0Ka5YZpkzUlk+ShjrA6mBpznmqwASkPKXmpD15y3rtG7EeMZgXkEy
djGOnrAVA12Rv+7PmNnsjCFNlg3biyL3Fh/N5OtBkZRT1WFVrRBxGnNI6bJ6eMOk
aSgECP47zr2jmyaRO038ijRzoxG7TQs18TjzIGF5Gfog27z00oyZ9Vlvq820VmDW
RhGdhOPxTvRxdBtJP9SuzLLfPdSDuCvhIEH2rF9sEHyuWdy7yLf6vtYTb8jPx+BF
yQUxzHugBhU/PTIdLeMEIXfawkd7FWcA4XIz8+hfU+Y/hulx2aFfAoB6CaEZ/so5
MAIL0jectjsrEHcbCy2KLVJ65G52n80JDhptkuFfxRu5VIpPR2kjexhLrUTGECmU
cobeJ5lJ2oJKZUUh3OsyxF5e18w36/lTfYJIot3wpA2Wr96OHwC+WtYmKLKuR+Hd
TwtCwUomuEUGDxmON2bNtKhpyasMDoYOCz7WNkT5Gl2L8ejFSu68DOQKTHdgMBw1
5kfQl7Pr59A2nn/ZtRPES2oMi+CV6l3dmSeepl9DhJL3S5HaOJHv9Tubt8rPUGvG
Cy2/HWMSTvFrmyyySEjs50cd6Vtm0cBN6u7b2Lc+9KE6whdcvItFEpqiPjXFzVdM
/2JL5WRmZtMvxNq0U6GWASod5x4L8SnM77/jFIw/lv+yEZcequY77NzMnW8PTDes
GuJrBwZZ3lWfKqvxzycNdhEvsQMbg5NrzpwILu7J9YqW4rLJKjbbjN4MmBLKalDd
YA1/9SLlXfvyG55zlbDKQOn5Zejjb46AzN7mg0NGp3Gy+65TFy1VWL/C8tY5Bbn9
yWEALonhG0HVHjwh9lypWZWo3yUGIIHxatm5G9sjSu38lFM86nr2/2jo+qRz0ZUd
dRe+ex/nIatT+OFTYuIxctKWfTb4MIuLRw3LA8C1BgYjKiF+z6Z01wzTs8gL9U39
s1CgQ+OVR0WMpANCV2qKf0LuJLjiubfae3CxxWRRejLC8WpElwT0ppQKJbuQV4qM
kzQrMRyPxeTAuQ22FpjhLU1gemSePCim4YkJ0lBsajek5OsjCR4HZvu7Q3yP0FEK
V4uU9e3x7LrlOqyNOfqXVRKZ+Lwnt/j+nLpx4DHF1z9LcPFqFX2cFWX4ccRFI5ak
kcmnQaAkMtYgrmPSBOdTnXIXO8cj8mGDbJ3WB7qQ+bJ/OxigzaLIwAE+FUAOpuvb
YCvvPgDuaTPJX0tM0ToO+ZLNxrIdibdM8gLzrKL/lW/6GKA3DcD+e4uxYiWd7A8I
YLVzr1UX+JsiCVonZULf53Xj0pU5bVgbnvUK39WPtlKQthZqeM5Waprm1szqG1/4
HzRDb/RreDW8tBuW/g1Sz2TGBsC/QpS82Pkkws6OrxIfoUHbGebfCpi2ghOZv+0V
YHVFy+dXjXcOpQrW4rWWMQzr5h5eCk28mBTr2ZSKOJbpdxhcQykxsCkT4jgDqSG8
xn7rXKmXbWjh1Uwh2OBWtISrPijbVf1fITiK4wNYEx9R+bEBvsUb/BkihrpqvDtd
v6nUhXQpmh688MtsG5428lgazWb0Tp0etx5C/3qL6IYxTvqS7aTtY4HFViM9z4GH
SFyAbS5yGAHZ9R6HWqgUuO6FL9RKQ+k7csHrxre3rQ+2I+UdDggS2XGP+KoeKyFf
gi8zzXDQZzp3dzwq/OeTUE3SZ4j8Aijpf4tZt/Bb3mSDf252RBswZTVcLJbp5PWK
hFaYa4f9++AkLZqAGA2EfbEnZBHn9nSCQLuePYMkj5vsY4raz0/fnS5+YsMcOl9J
vgBbUATTzMHI9SBTow64xDrGehRiD6nOSdhUVByKksbijEL/jFvN1YPQE+JuXVpX
krqX7sqc0OmQwNkpyiJrkuPKho/p0z6deu/C+apSLdqarDBy0ILBEyK6Xc7YnWe9
iwudzHrvRMmWrvRyMqyDhfMVDYJpw+AM9G/vnng2HBdUak5faKjn1bFf3KUCiWEZ
PBWnw3RemYh1+SBs73hYG+gRWSG/K1+BOi182ZblrafqSUyguvh1jkGymahR3cQl
20afQxLsdGxGYigdoBlxDfmf7yOkLxcYkgawjEbv00c95eLi2e0Z0ekMIoAg5eRt
Qtj1PvqtwNMHhyr9yunrLC6Z1zbnX9BG5jTQn7oZUFTp4QtnfTVHusm2M8CUsg/0
CTQdQzHNF4FB1qRyt7Wv9JED6EESfu7yVdEG1paayWfcV2DEcyCZM3T00ntHUfiW
3dSTg81MkW4IynFWCNhNH1weGf5ej+AvUYDbHxnYrWAooNmDM7W1gi18+tM89kC7
SknSIYIzHa2xHTy2SA5U/e0X9rIFhs8STcUAWQOlAnd5nBAMnqYSiMV0qq654pJR
dvV1cPM4awk0MfDXoa2H8TVINMx2lTYws7mZcVsJL7cRjZDtf+o2UlErBDcxGjNT
Apj6Rg9qq4l/Ree/WcJfS3mLISiEiLdwTjgPweeZOkzkAcXCSXPaeBA8qOsZFwo4
EZTfz9R0RPMEuy5GaxfOE8hMASkxcJm3d83Zlczx0mLmg+ikaiH007RFRwoNK95j
ZwbDYQJlzQ1lx0dNoz3ZRHX1bR7LuQLdHtAMg07UpEh3AbfcTmd7gnA9bUd8ESOE
aM34yEGSIKEi2mZLSZmiyjd8A7reIPiNEGP/VQWdH+k+PfAkK6fbDJzaW7yhO8eL
cXaOksVq4vDHijZoOGq7T6VEjU7AqW3zgWOsc3XxVYhrE+VmSA2hjhw2q6l8aRw+
FP1FL80UGh1EwlGc+bHUeKyZwWA2it4zB5Ij+O/tkA0BsIWoa9fL3sS8esjevYvc
qGz/iuMLQbxCgraLk/Eg2oSJUTxqx0YFeXE9/Ku0tfydYuh/tulNJRTeJuSffr9G
kjMtxxAsif4+A0TsCgBBywYU4kNBvDHXGh5ekmpYgE1w+eNolt3mRfV+Hf+owyfH
lSXpvQGv6zapwfhWxy7HaHizOUMn1PYbXa3/yX5c2PDeLOaFa8XPHNFmKpSOmrDN
Hhesg0IRGYTuK8UHbxGS3iZQQA6Cxf9eF1hzI83zZG/wWOr3pOSnvTBzR9sdeeAw
5317RUS9/4cmrFHGvjaLF2FFh2ObaoHErdzOqkqtRNO2OiSy53WgbdxDz3BsCYQ4
5zAuhYL+zmWuf7hvFse/u/HafyRoWl3bMhC8hGr19TUM9siqkYMkRCGAxy0AndLf
4DZtM5LeUDMRIl6Hz6hOL6Q67h6TItZX5R4dxt/aUIFaYa80+j8sD3QxtyprVIV7
g+xLsi1tnGkDcrdfBXtg1wUNIJtaWA8FwwH367pBAprceprp54XshSzbNLpJL2Id
VH63k+vwBEofJakwMSQ6r2g18eWlb+l16/7GBmxwdI5POeuUr9M5ZP/1ycZUp+MN
5Yoj/9LegEmz+D/WBIpgbqj6EK2IovnCQwh111i7VJSTphCGUo8Ilb5iN2Au/Yps
FryLJlj+0SOyPfORm0lnHBAgpEzz3PqymMgOrb2B/0N1HePg3a+27j3eLUbE9p86
us6fIcCr5PoJ1rgxTzoh1pb+f3SCOUdWnRDzfGV/aRz7Fa3cy4LfMzrIvYGyrVJS
E/aYXXAfag/xmuo+Ch23pFxQjdQKs/vTb8HIN8cirYdnQXBjM4QWQA10aEl/gzjF
WFCoyXP9bdJDiJY+HgrkLXQmhQ+h8pW6Dq2SmHhTzldQ8xgxpuC8F07kJsHm3LKV
DBAbSkR6nKkwUIeMFVAuZyQGS12DVcRb1CsV/tVxBZgVCwJkfQOtjcU8yf3r8ezh
i1wdWRD0Eadn8eny18mK89V+Og0OJxfn2DNj4sYZp/laHmVM9ArKDA0rebPYV87B
ChEg1U5D9xo+h17DR/jHE2K/h3ZqZL/mxn/wqf9ewd9+PVURO5CprqAFvfE1ZReu
rXbIo59kQZOjIoD+lGTYVbq5QN4ephZj99mnRpsiXt4vwmYJxzQHjC9E2fS5g+OP
Bifhon/c5kF2KGuhy80RK7skkBt4vbNcSZIAnsu5OqD0MzfHa//HLlzfxPlG8Vnx
SKWuFDGlZ4pe9NWhdIjbjJCeNAvqII70du/g/qqziQ5uIvKOcCbl+senmRd9OMfq
tr/RaFP2D9Gs3C656hHjg0dR9PbB7sJT1Ci8B0UVr482vD1G3rDB8QnPIsUDK2DD
Eyjm51CYdZdTwb2lwmt2Hl83bjy7NmMyhOPRyE3DIQYoRZrYVBfdt8OMT/srjytc
Xim+joH9AnjaFeSXG34XQgAAZzx385pzOuGpKIOVz535E8sEHMzbk1SuDzpNDaUi
d1O+ZOIWKFN2hpXD1ykNeCKxAfxrWRpFcQyK1jH46UvakuIkfMFqvKklIfJzg9hy
Lozu5PIIiXhC5vzHKNRkFuwRakCRvYfX4y44/F+7Ic6ltDP1ap65Ps+BPC/wNbIx
wcYkYY6qZXyOQRWm81EJDf6JsM8C3ktEINskcpp53aTVlcvhr8X+32kia6QochEr
UiITEFSCUOeN/7rIetL/aECj0G3H8htJDk5/gWtLIpHKtAmHGNaExDKcU9va+4lt
L+HPhIrT4y1ttT5v3A1i0Gi1uLly1wU99Mf8kWPngFIKknV40YNRVYNwMAy8UtLR
wuTUglspHXhV0rXkgbskTRixjg5/xwpGhgWOb9XEyySz9FOUK7tnRcdocctmLL8+
FXET3vPjIp3RMCZ0T7CN4MOkYXWBToptAO+YHRXGgaMiGz3B0QdqhUCRTUrVyFZG
4lB9zeqrTNCImyVUJukg84AKJMeg2avbxKhpXRDhbvPWun0Ldo9ZTIFf3LtwA2L0
6a+Ueo8OthcqGlmAgnPHcV2UtHnm5d/fG6G/DZNeVZhX4xtpoJTR4kmjaEt7DEb/
sCHzr7wiDBUdZIp9C0Ei6+hruT3jufPUc8pLlM7DMig09PdFb1NHH2aThLYFzpFV
2pmIi6hLGN+5ieW/065l48qUOkNfJ5oZ57o69GnkYW6fzXQTL7mCJ5CJM7ljGYlT
5bLRJp5ZMpamQ339VCryCQjf68q5mjHP4D4J3Buwz/zvkdqmaY9ScBSRnNU6960d
UTnEVMcMDd4gMeFqyvcy4bMISKnW3gdNYeUa3v/KimXC9xKVtjvV6klyttDYcv37
CslhyKsfzXfR7LF+K/0y2vlokDveJnGJDXAThIhnwke9D00wsZFDXajgs6e+Nsjm
c73y8NZV5ia9E4tViiLgNs31BS6dYXEFIm7T+AC+IDgPavqjk3NIGOIDShm2gTsX
l59zEFFNWwM0i928zkP+Esare5cxrp/3Av8DIOxem1oPoABh+8O/Y7Jumiyz46hx
3HphTHz4QyT5YVW9+lFWo/tUyr++v90MSVGfsJGKywYyGq20D6KOM1QThQcV3nDr
ankDsyqYXdm23aL2yF1VgqhMR6OGIEv0PYkp1iccffX9LD6V+vrfYqZogv5FzKbL
8bDIXi1XysiS76FcSE8lOgwo8UVPH/MNQF61Tvfwo7VKvpezVqK5yFG3/XQYq7fw
yR5We11L6AdzClUKtQtf58Sfl3QOAQyE5kKJY+Q43euOyxWItt5EzyRkZbMwhW9a
ImkeNCE24OSvvcgJ9ZbSyT/l623fH+aFVaVWtW6YlxVFMfQMOxWswsn0/Yw1smEv
HytjDk+4GRPG+UCMCEVh9nx8usQtIBh6XHnDGLWuiWJuGhIegLAAhJiMsfIiAlW1
aFTTV1lny+tFwW7sbfccWTCCerPROghyomw/uXylS4STn3g++/F1aRYZIyvK62He
eOGjSONgMMhDHu4JxaWLDawfEFhAWwsvsDy/doGA3peI9EmUhEXLpOaWv2wAk1P2
PN2f8Qxg3jLkllOdk9/LZhBFVncQKcSdXTy0nxZrI1GP5XQfmW+lpfV7m6wPEaZz
nc8+aXoPiK7hxIvzwUoYLKb+VtrXUkmNIsPFE6gmDxcWk8IrDybZ/Gbvz6ky7sPR
yTQElPYSAt2olaUml2UTGzW6kezijtWiVJ7PTztTa/WIkHNOGeUtD1Z18j9hA1ox
82S+7AdQU6sghPATT0f4LmN1NjE8dM9/MfmISOms7yhkkxQ+gVIhRCIamGz3jLkb
nkrMdOJW4jN9e3CO5FY58z8ZYzAEma4WY5y8B84Pc8EpljFsaFzBz3dWT8W+It2/
mzQJdN8Edn2CzSfhY2qocvaLzhc0uGZ842c2BoeqRVQP/3A0YRhzusnG7p/Ufqny
Z/ur2gj80Up+/r8VkHijfC5BazJpcZ1BGmWgRXYhOdkj/OpUnWz43zbFktQFqBy6
8aii459OWuTCaWVtYwlUfObdQ5XmUWdReQgDghYScfs9Q1+2+r8tjpzJQc0iuas6
zNjTH+rwayzHycEA8WtU9ZHk7vQh42nUwag3njsdOc8sfPKZ4vd8vx9C6f5yiIOI
GEWg6Bxc5ScudrAD35JfqvgSziMqMpFdOnu9ctpA0hds4fbOBC0/9VscuBurjrrl
7DyW/fRODKiWHg1wvZflkaXjRht2FfJ2YbNWJb1hx0CRKHy+xzUeu7sWQwAe1wrP
WbahAYB3Y0TFUV03cfxE6gGfaNTiPNI9agFHcQj+4lUB8VavumLmXgzhsX0BMvOv
ZTkj+qEyzj/7T7rAylwTtKXS/31E/liHbC8+vhprJIEEvSquIvShEGR9dQDJTRVf
XB4vq2N0hTp3VE0S4BZaZzplrt439w/rC6EtYuFNxIuWnZNqD/BK+1HOvbbgTjz1
Y7ds4Kdcbuvppb30Uhof45x+9jDALkEMN4ayvPyAXFFnZASfXC2jwP5Fpwb4M2J1
V0HvjApOrXIkz/MZQS61UvQctaFMk82xMfr9AqQwCiq3vBv91WKAIElVYOduqkug
dof2ewCxGvWtAZ+ebH3l5Nn/dm86XeNekLdZSin3gAD97hvlG+FmFSWh9zXHxT/I
gUOvHy1sRbNAF/CRWf7RWCG9dM/jpQpdzcAVj82Qv1IEG/VE0yg3genBY/joe+Fy
qP7MK2irpUoJCpy2h8oviawqi4UWiX+o4O4kGlRd5VV5Tg31EvKtuzb8xz0UnKSy
wjA/mkPy/OGpeMSfsnlnFdpcYrUs3aJ8x1jxGOiBY2LYM0uRON4UCYeDKqcJucgT
AWR9uja7NFAPHI+EwGZhqKHmJoyeBmsVJ9cBxJMcvQtaJ2IoZ4F0mJc0r0RD792U
lW6Tb4HhE7ADH8rSQMV+gjW7f2YNEhrHrjRgQSUIpKb26DjI7YCrtA1X0Ez2Rhk7
i2m9eRYEFi+D2HuCe0+IMQIAembeZ/Fdu/r8YE98zA6II36lIW63WxTD1jb01z6h
HKZEgUO1jii++xSLCxyZDjAAjCQZoSBSlLgOqkA8F8jQfeW2TtSgRQwGHdOW+hG4
B7AYahkn40PJwBVXip/jmwPwVcSvP/Pqql36S8808ZxB9K8KIk9ktmsfIXiT0/It
bZjPmK+Kv5Q8GIg3AuW0aJlODtKQGdUhcY7vrP79s9PEGFcyCYOrM8gI31sKxqXy
f3rVylPtkOyWKr8cHQ+vyPElW7fzqRhRvqrdtNid94rUTayEnFtUSFraZRAdve8b
zWu6C6jz4ch6p6Axspt9Iepns5LSHkx7xvCXzRCr3ZUXkiL/5GGMkOJlETNa0Lls
zD/HQ4TlhsEz3RhSNV45qJGq2/RCRHBfTcP8w9yV01PR6mf+pjHD5ApwVAETQwUo
5Ax2+Bppkrj65SiQC8McBh/wrZxUYrrmX5l7fDibb+N9+IJuYGpPzr1MpFX7rDpQ
+SV3EWbRV4eaj0d46AMl002ULW4uzmgD1UIZ4ZAo+aWBu8re+kYMRfsBWbXOS6lS
B+41zWOUbjY7SUIMqemnhhta8+LJ03VLSwMrGJE2rIgC3D0Lot9p+Q5H00x3AD94
b0ZJTzR/ayUuaDOpaOmb6XD2AVM/MiQ53TCyB1uTzBW+SjIFE1FmdTm3nbN+JKXy
zUy/6pjDwbft6Rv1elpB+XpQFoPr48w1Jw8XvWZlx9CgvfsVyEK6y+SH0Juec94d
GtXv9xGLK++ylWw8mNtlTtr4qv6TVWkmdlWRzZ3FJcBFzm60iH1jEH4++qCG7rkH
2gvf4pwHgjJFzhDYwHqOqFhGe9/T88YXAeKPC3M2AtEdhm2UXysWheuM504lvobP
vMBBQL9M30GD43+S2UcHKOd9fPMzSdOXlI1d3uA5BS0EvBvgd2yjsKfc4V+w5gIb
Zp1q34VA9adAsGGxhLuNZUevaaKxzF43smpTw1SIUjap4UOrgY8KOMP9uEy63m3T
JErvQkP6kbkgV4qU9f4C/Fd8bYg+BWShzjuQ9nPakyAw7BPG7hy6jxDsqa4eX2i8
yOzCy8C+3xMeoSUF6eO8hBpJVBTaW4hkL1RdnmvKlli/jChVVjFSP1voknC2CXdh
1JieKdOngztUoDuFM6wbBNniaFFISafSyYC06LSbOJGrf4524C6m2HQQhaRqAbgE
WYcsQOvQUF1Sl5LDpnezehxagAYBnh1E4StNgSecfMxsC3p6JmJsUQOo7svsB6yi
pV3QocH5wzw+T92ggimcQo0qYH9hoJ7YWd+tos2z9SAuffnOIKmJE+BV97NLGHyQ
mS65HIQGMqAbxU+Okae2t6AkU5aYlGWqqsiYHSu/X0IfZP+TRefAhSQUtEKXTF2n
jzNCP8njVMX6meUffLD9IxdvDie7vNzt2WifHfdAr+yOTS/liuo3sX4q7gWtVFkN
iwAhW1eDyQDQPfgzmpa/4sHeZZCbHIIF0Crf7lYe1rK4Cqit8/gNMvsZXOyu72Dd
VyR9YXPT60AKYZ6YddleLDB4VcECJWNeUfQIn4uWxjZkC9KIkiLDKjaLNbOO0QMZ
NsJsvBISzd17VTC/XhFfnr4WsgfOtKkB0e/xGmvVyFcT9JWAqA9l992p2tgpZIR8
uzEmnNpJ+RdTMp6r2SlaNoIDgDKTsDhwDdzRjvwwlIbjWJuMVgEZeoxsrNBaajV1
kVZbmL64X78egX82LNbpbtsycJfzyl5x6Z3IPg1sQYbAKaBN5ZfhqGJ519f0PB4+
GEqDq7rh3doU8jvlRZNKCHAbApnHOIu2tq95/sdWvz+d3Msmpu+PLDLO41WwGixj
KJx7MHEu/jf8L1dRaKFCPvYvzrULHwMwZnvvs16Y66ZUzCscOfyW5SH81qo7CPdc
zBL5hSsm/7mpNZeJT449gFRWF9EgjAxOhJxzAXFZe6oixkS/5wVWCjmd+g3oo4E0
LwEMJBrJFCy5JlIL5sE2/i9GCiN0UVOrWbl1AR10umpiA0FhWJO43AGISCnVzb8Z
Rv6Ic7bT+tkWiR8at33IOx4XcoKmjeEx+UjzPNXwCKyqvt1f5YvfXKIjbVvqoaPm
pJbp6G1oxpw3aqGpustMeq6i4u10n4XJo4FlxVgysJtw6sWH33ELeuWv9YX05R5M
c621pLML3NwmH+bLff4B2RmtcpHKZtx4Pz/uBg49+QqoIUqa/eRSai6sbqjYRBU+
hC1Zf+Qaucz9NR8ynYJGAK7idL9pG8UbmliXDnTQVlrIio0gI84khJvaZymgf1K7
BuHQgIl7tz99gKGi0pvvgd2dP9Y5xmeGOp9U04eXBLofvK5YpL89oPwk7NsBbQ2W
wnmosGxgaL2VEqzXSyvDE0+g/D7gDxFA3gfxhLI1Upw/HKI5XBmqg6RzvIqS7k1s
fJR1DAor4fIb0NtytwuMDSymWBC+9Winfa/DzCnjrHLPr9LTKIOGkrlJcRSBWxwZ
0wmJesdRUqwOEypEIPYTl6JA2r8rG6Pd+Z5k8mSu9JRbHvDjXRrsQ9tJi+uAxNow
NORHIR2flshvzpsShW2uoB5MdQiobHJTVC8Awffi2r4wza/eo0jAJsOCwTVCzVk6
YY4CWPBO8ROIlJnVZe1wtTsU20gphnz62F5rqlfKi5gvqjMW+t1d1G3jRglaNIzV
FhJqGE4J6aU8RBXo4dA2oJdJqR67Va0yIrrW/2wz60XSIrp717JSiWTnbFbjIgXk
zpCM8dhTYnvVMpolCZ0bFFflyME5UAdkr+6u641msvZ2EllpqqEN22/fbqWzws7U
BqLWaXYXCg6OeaHb8XEJSzuY+GUHLuocj46vGqM2uXr7KixCYBc56p1IwRwCmfWq
cbu1SW9xK1FM1gMTx4nQhKRrGGgycCiWOz6Y8AMyYVMeIPIl5zp+QFDepANJvDbT
2L7RD+BQqXO3gncDTAOaJX3Fa2U53B5TvaTaedQgMElKl18QrcQuphDzNO6bW2oJ
tykWE48v8E1EsUZP+ZDbuleg820k8qw+alSe2JCo7Wb9zKjSHdiw+RrJUyDC959d
FPLB9ySArQ5YLkbkSGGE7kLDdbVwktXbCf0ggd1UIvlIBniOmELozhk3h5Jo4aBT
alSfQk/69bmpy9tfJ24cRPdLfZHHNs+751kq3/ovdkgwR96NqyHORRa4DRyZ/rpi
BQzmhmlZu4ILtnnrH3zNCvHou6Ik9HADzzM7Umj5K9OPLDHtkzTPLsN2149hhd+7
D5iha4JsrFEK+Ld1o8XxXQ6P0LT8LmKfoasF3EBRjKl63QBMiC+OqiOykNxwSbnT
RTCCA9Cn4xZu22b0+VNfFsNWyLBixswrh01TIFwbFR5tafbRd8Ea59vNWZi99aUc
bGEC1LzQcuOW05a16YsF4yrAhoYj1chvzm4ixZ8KeJ/lTQfXYzXg2AXg/CAiPlgC
97c/YK6W1/58MXbFRhNEfIqEp6Y4uIf1TmzwUp3dWFW+ntEGohXQR3peueSC8WYo
x3ZcEiVFWU1oLdli2Kyk6kWcsJgiTr5qsY9Pw4lS+g412cX484pW9sCqt0M/1X+O
HjyZensJRVIZadY/gEhh9j/OT78WwoioEmoDq5Bm/h4FScVg1u5PGvwDDQsM1t6G
620Nw3aeDF8GlR/CX/vy9ZeEoIXapdpd3bWv4TMNf9KwFBR4rR5LAF4U2cZre+bI
hvE+hIvJQYGGFk+Qo/LfM62hHIiEjGv98I4hdf+l2iZ+D6Frm8itiypNrT5v4ZP3
U1IkFW2OPliFAaMKko5JBZAlDK1T8k0dTBKAinYJSmlkvZSJrjMPwEmsIGZuZUPf
d3SKD7Uo1HawJt0ZzF8deZnH5KiDudoYbOCaSIyIPyNkUyUT5soJzEcjBnnEJijK
8wNsJTe+rBK11tla8KZqEgUGwavkD7djbWGhJyHPl4nskC+NGNFU/g+NtVqc+WhY
M5vfs5PEfIeZ+MEE6CQSSwTDhpAwWGrAEKqjEyo1+y+bfskNLvPsOu9J4kzdnkAd
sCdLQoHHUvqDt5Qzc1p5L6uYH+6M0wG7dB0zt2P2xMYghobKR7bGuPmC15ML6G6l
3/KZW5DLHNk0RDVy37m2v3k9ud8CoJVyxrUNHlASfQ0DKmW+ZdAUVUR7AB/h5Ptg
xtpnNTjDFwCxhcT32DFWfgq2MdiMz17torqhc1ccNbSd1FsHAA9AI43TK3ccNacJ
zzvVCOvAIdj5MWNdcNEwusotGN0P6ixlq7VnOjOJP1rGPSL9r+4Op+NHNH1qc2fm
Es15R0VtEnqDL/upBAZjrILknDMALHm6+TMc62BGTuwfWW+dzfspTKdvZmLmYV+a
9mZuAMpVZvTqIqm2KixAuAdIUOlQssA/k7j+C80eeKpFhYXKu2S685+REdPIIEio
vmNME7KFOoFvoseAs23nTLpcOCJVI+Pecs1hGy/b/jSSEasfxgSQURIpYhOwS1ki
J0/XzHuy5hR4V7uAwu1AtH/RukL+0rqmAOdj6PfXhbdO84FGdC/2gUnqUWWaP8/5
JVoHEX9xuADXLH0iWmAXoba/G/0ct7DQHpS4vOR0Kz7DyuDk+jmoXw3lXGfvezE3
/5fASi0qk3FEEAv2zDnSm73XOUAz0XvHJ+NtiilSdmWror8ByCahIcZgUh+pqVxK
MKJd4UjRxT7/x4bB3LIgak6oyZV4ZAeo2x/pDDccD/x4g4Hg4TxaB0uobr6X5Pc4
OECKGR9LE9eF0uUZ6YqPW0Kry7x3j85sJJvSoG7KciKkeP6lg78k1KxwBd1tp2Yl
WwEnrVIXQ8D6QaE6g+z9MLBfFZaSKC5N6xH8Wuw1qcznATXjZtxujZCypSoFI9lk
FstIfkmYGGHgf+0WAzUX4qdyjXliDSxOTNF3xx+aO89sYbvb1KOJFSSrZyqmB3fY
xDtgJ1ssuQVhZ30lqApUcDncmeUw3utx4v/F2+5IEdu0fWib7DqlXA+25bOlzxPd
gct2uz5OmIE+oOvP2TQHKSNhG6dm2KpbUF0kEI76p3gA5KxCkUSNE5Rba8GbYwKv
slU5PSE4koAnWHeDltlUlqYnWb2XztiX30cPhfrOtuqf6OIDYgeoqLjUDLEotqeV
GygCpebb/yF4UgTOIvsW0EF0b1EHDTm+C276Uft95sSyj9hlPyawd4I/hk7j8aGb
Nwo6j8puvs/oifGGp7jV02RSnjLcAO0T4GdyaFkuaiO9ZXIOakCJR3H1XPQqQ0c0
f/NzA5WzoGqbX4+T9w/KmoZqL07Sh1MgQ0XS0WbXVAaKoJIIfRJJZCSz1Ej/mI3W
yhVEKcG1umkcWvCFV003VVoRn9/aqTgJQIzwRWqx/G8U29oCI8mCfjvNMcvkxccX
K3y6mPRs8ybw0qFYVpOe7QFMkiv1FfbquezBK06S85CLrx6cqnIMzed50RsfN9Wk
JM4VMSOzDUu10dKcXq1q3hXQLzZSSNpIJruqyKIz9XvNUwbVVdJFil7NEvF3yKht
4JjM4Ku5wuVZQTqj6vF+vKHea2bqDSwx6o1Mj4Pb4ZFZTqAdzPC1TmE4XVDj6LwO
UPdA36cZcRHm5+f3OIEDza6OnIrG5qPs5zM0gZ0w+0NcguB+imacrY99AZnlWm60
wLTYHKgqSk3GubXajcLgnPmxthLTvuBgT8pm48+DWcD1sC+bY1Xp6Zj9RZRJMq3s
YJLbo3fDjGYsN86gNPr30FHWfJl0CBVEU90MUTxvLeoUhpnVkVp0Q5hEBAKn76cr
fBZSB51RdZDZBLqGZ7QAKm+gmz3xI1d9douYueU2QHKkuq+GTMcGxjOiuM1/+kJK
Kn1UOoJrjbc61KzvIN8xPPVUaKFzE1qq+N3mi7RE63QlYUNrJdkXq6DUQ8kIIR1+
iMjtS8dEVsWsg+gk1WlRPDmkQahHll8MF0IHNtiNAHifJTu9ra51WF++ZWNQ+R1M
PtRusw+Og5EFkA6a1Yn8H66ZtAsjkyszQbAK6HtKyv+Ji5XaQ2ToFIM7TuLWK//S
mtdiWVmcMHw8qJK4ftq0iP7DSwtGI1dMTmrfU8djszmdJkuMmU26/zNNshYWS2ty
JSfrUkP3O0uzzS0mKW1BSEJ3Qye/J6FYkhNZNGKbBM3yFdJ4VvyT15HrIyyNI5Z6
tAhLXj7AmxQujbIsZ6XhuNJaaM/0Cw/so1boIb3OG8CYvfYTp6c8+Xz9pxwwUMfd
AfirwBSahEdKGV5fVx9UUyLeB/FHuevAE5vi3IC3iHpQLm//wm01P8nilb7TkNoZ
k1i7mKNcI5ikdzSkyFtJlXHd1WkZh52Hz/hNgFg7cOMyiJfIGEJUTN+UaXKLiBod
cwRy5x3k5Ldftf+7GgfBXrrA98BFF/suscgEzVSWVP10HYzfez7oDUniXdcohKza
GAuYnxA7I8mcI5umGmrGsn4usTsFmDSqBJUT57c5l2dcFgYdrMk54abG479T2cgk
wJtc248YvrrYGS+6Zto3RU8JhOcTAolrdgYMCP+XzG6fnR8LvzdCrP9hKVXHb1/M
E7OARULMfaE/e5942d+kkizlsOvHTni75YuWR56ndKnbZYc9XLyViR1XLuu4WBTQ
WxAReKMNcACGAmOfVkQKBATt/NWWBgo+VG37y7zpuBfq/u9WfnZfKdeyfeEDUIA7
wlV7SCKyrSoi+l+S+JHExYNil+DTALxL/px2OFjcKHekJjm/F6LsAHy0ulL2ynxH
h4GMWQeWLC8MkPaUeD7xvN+iF2RPsizmEAuYoFcjKsC5tAwqRY8jfaTCQvz7p/3R
IycxJaH5wNhcyZilYZ/EFvtvRrnu7l7911K09vbyKUDm7anStJG+hPMd2agAnZ8b
flDYTNMQt9k/Mk7TwiXfPTj1DsAaIK31zKTczfY572prp/lw2B2MIvW0R+CmCwBJ
oTk14ABxPenCJX7KmfKMcEdkqJrwIgocmIEzIjJT7ZkSybfk1TIN3xl09fpTrDd3
9NtpdKuPSPGSf1GrbYk4ndJdbePq7TgIGRtB1EOTDXOPYV6Hru1OlZnp9O5hdnqf
UX6dNkKRcPfmTDHC3b3RAmAf63wpDAaCnYY9RbM+aK/zulaMoQsyKej8ydXwVvpX
Z+tFAYQ+UJZ6bhHpTdsnbvVgJreu2bD96tI+SKK6IxtMkFhC99NHFHdl2IGg66n6
0w+zwhFw2J7RuzEHUupPLO4fpntvVTo4u7z+NniJzbhI7sEx75yeOVwOLSUrHLWU
W5yut7gFB3+/mXv34zHnTvhObVdUZx1CKH+cCN0Z1SW/JIuenHVy+ySUoqbdl8Wy
QEicrVSOJZN/W3v1KNpC34feP0BFEXaNFWoVVx6a/2b2xDRCj1wG9F8Y5GXuvl+Z
rsmi+sLeNK9NXbYQMKneKXn9NeLDJaVZkFKsYHMYw5H2W/LO9+e0O2eDpohdo9CJ
AaKHhjEgRDYxvUHnuxBsfKjpDbrq+FJubpmJYYW2IKLSylUulwXkjAaH47pk+iQO
oPmSn8GfNvHoFN7xaCy8zA9PdhDSThsvgKj6uD0EkcIYkKFXXMhyAzB1p0WOx1Tk
y2FozW5qHu+9EplDmFaJdwyHORDtcnKaWszwh08N9looPVNL/7maUNuPGGXnlB97
UP0srnt1UITB0Z9NMKx2LlVH/dkP74jpZujaJ2duUVCGvI8feYCUTpxSAr/MMrkr
7T8v+M12jkJFhXrwHM4FtU+I0rlQYH+DnVUlvMlWFvPkBCTNc1QqK1/WI8kXGKZx
OWdvZXtnEYTvgoGi0Ba1zRuShABA+EjBCFNJeRlOWKbjj9fIpi+5SjXOZX9spvqI
sL4JFMAiwdFGBjhv+7n6RNDfm6ulCOpaaBlg5I7gG2eIEyPQB1qEuyAwubL9eY21
/MErL19MwqCUQCNjhEgeEjMBsAycPY2xDipmw+DJ6HruvViMNJlLScYDmDktNuRp
J15QnpIEm9l0dj1aEoeu6u6xw7J/gvw8U+9CfgRGR5sY4/o9iTMltT7Q4uaq3BU9
23OdJYX2P7R+1TGH+m4RjQ7BPtJyLsQnn/RmxvBvaB81W/ybQxbNUt/44Dd1bZlO
I+iOYUkP2dVNuB/9rOC8MZvjGuInKeoabAr6OzoxhToVGAItE/hdZ0zrhfHnuF/P
Ji0LaGBXQ3LHlzI9xkpOrdm5wjvB2mYAbfW6b1FJ1ysV8OCMUjJJAx4h3tscfCsu
0DI9YLTq+I6Vvrx3Xajnab7YAUJWOZ6xxMMouCSjj+KtZXmPmDAveDAsB75fglT9
i5WumKt/fActfudqoyKZjeK54RDEbroUuzl46TxKIsEzVfpSBzYz4VcNCtc3XtIg
YqvGFQnDGv/CNWCjBlCKwbVcTC6i+o5ZNis3SNiaf7UenhDwaoCdRMa7eCZ6LhYm
27BcMj24TskA/9oOmr6Hcm1UXEYhvE4/GjS4M5Jfp6k7PEzZ8ZklS8hEdpbD8XL4
L7f+U7YglRAB+xMUv+hpx/P3tRFhaC0GWHmyYjEaPrrrWGq1DQZg17on/EJpIRns
mXN+uvN0yA5WKx1vIVxWfixyo670mQLbfwpSvrwRXgmK2J3LNOr6fBBokqzrjFDP
tc5v4N6iZ3bbW6vkUnf5eppafn7Hkpz9kMAjLYdm0kEi6i0DAoSUxVO9kOsVdYmJ
MG3vyeUz2qBxCQhnRLj9q5s9b1UpTHzZkkleJaaxT2CCenssEmV8CGUMNzQvSfZ5
9YsV86KqtnG9j1dxQ3N+gKMLu+KmLQqaorqtILD3jn5A+joVoI+OpUymeMcn80wo
y27kUnuLBDmeJAQwlEshqGps8viESRVp+pZopHY81CmCMBHkP6637AZS4UFEc6ZZ
L9BwBN2V+e2ZHs6KasddVnYabiBVeau7LlHxTMLUe5kxqyQPMhxqhcOFwnicxYNh
y940jBiUxmuEdoUVtv4mrU+QGtaDsxg9aWTobR+qhUdH2qIMCX5FDKUd+QWv/qk8
H3s2tnM5pjOtBgR6WVrKNwx7FZBGMi3R1q+5I4ADL0dFGppw8XkHKPUzCxZ1C2zk
9N1HFKRXnYKZXDm/mfPFcE2ao7ZibXWl7igYGWuj2hZQRlSDmFcXI+4ejo/Nmlh1
A3H0LsO9OyRbBQHIp+jl5Gqe9L5pncgKxRUI/nbyeDqc8lasqxh4t8yFY4tjp9er
aJMc61PH+nRSksCz2QCJ6AkAbgVZGDdXD7KyFOmwdBsoxi8G+y5GE+74XjGlUtw9
9syGdWGtB56ZZRUFY5JyWHA9B3EvNqPJJgEJG3jle2DAfCTCBClawHdyp15es64P
EbgL8z0GiLh1j5eM9/+LR+VW+gc7mnBsbwGuLXVS9EZEhlTE0EhYlt6BbO5/+h2i
MbpCQL7/fR5dmAxUe/YFGARAyUJTeUf1qg5psrivL7it0wC9Qa8qTIppXGd09ozn
+uUWBzdaHfc6JLfz8HS1MeDJVIAZ7l0mQoNm52baX+x97j1EkEytU8PZegJ+C4pG
lM46HKAVJFnWSUKEV31C3HLqjp11h+WcOD70SPSny42Rq56cPQk6/O6Oj9K5zp3T
ZrIs6GLM6wS7KHLx8S+QHxYb9hyoZG/bF9FoXN/+8ndXYV7yq39QxadFnZxklYew
rCsfI6Mfd3KViEDRzBU+FJyP87CYNQhpmjQpLOY36YPU4Z8oEwhaYEXWHD31e87R
ueQOk2uYOjNHvMoKx7vUiJPOs80UpRzb1oPNwuew18qrQ2HHOCVDuFrIsaCgGKki
BIpM7eEymTEUYbkAyTecjiUW4Hn9P71+E4Uoze4tiIxEY5bfxD1Zqo+pOPZ8tHXm
s5DMQLseyJCkvZk2xTLz0oBQj3+GNxzUd0PuMc4XnzeUwREQNhnLIImpyWmm5dls
zHY6gk78KZE7m1FDXr6uvn7PBdVuHfJTeOdnByL7b/43jWeKIHARh7cmDY1ViTPt
Cc4E5bMrpOKa5RPomIYtMyw5RUnKoROZerfvgVOVvZPtJRF+JU1X1ADHxi2WynEs
jWEL8m8RH79BtQR2Kfo2FKqhRTLwSNtQ+fL9Yui8mC2uifixKDMmOY3j5X4USIpj
/q8hiNSiaY97QWvxgMtzEIDOErElNSu1ZcfqU3luucRshp7q0KvQjt31QRoXVpdg
O3M9FHxRmV4pV8nbpTuWp349Gzsz8awlvY67bNRjvv+wucXXFd/cxZdzdqu48/US
V1GWrWY3fi5GazyftVz5x5PDDH1fqMY6lRjOIqQ0gYFssn21Qe0g+LOnSOEHGhj2
V5POxAFjwUYxCPTC8WGBXDJBVImxKbThh/hAwnDvtGIjaZNIqunYQSsA3PpAHLyQ
9H8aO1tFlle1IHFaioVxVoB3zqGMPJC0iiiUR8McngGqi5BYZ/7UO9A8U9Lg/bAK
vXqjzbecHsQ3PAekWskuVLfm3tYyp9HH3z96TL+QvzdInL7JKk/YNXEhMxQK3reQ
Yg7Rw/96qLmu5meU0YbMbZhMZMYs6c41+pQEV0iBvx//tmykOn7uCbTrxnF7bmar
KV8JuQ7LHwaQzZf892KRCnqx8WyugUahyf857v1S5ecL7FWSqKmS0P/V4GmPa3EU
A3cnhlGyr4KkpaBWy2u5Z0EtX8J1VwParg7cPH9FsStN9bpNwGtFoCvR6BRVd2RA
Ko+DYk84SiFzxoQQWgScxh0cPCso3FlXL5U5F0YqCCwH+PJLeak3riSPti50WBv5
tSZWG9OyLfU/Fw1ru9x5YTHM21rvTZzqcwW99usWANIsvZj+9GUwRj6gfpyHrK9l
LjcUFyWy0hHWUC2D7yrViwTTyNGal2CJ7l6DCLOjWFxiLxRk4kzNLNnt3lBeoCmk
1oBXWeWlK93zS8UdUsW6R7jPwqiPTqyzH3j92tIRH+HlDKAJp78WqsXeJppvjRFC
hA+t3rqW1PL2AsSXDyWWpi82ldM/UGhMe95hsJcYcF6sHY1zwbgEo8kyBA6K2l4V
kQboRDK3yvqgRHDQD8DWuv1/ruvm4A1Ss36Wt7lB6ZESCFZyjvdNFgI/qpe/Rkva
SG0ElqkexQa5cgWjXMfge4M/0twUVNBAKWuZvYACfIocw2rMd34AnokHJnCcCcqQ
3c8bH0cqxm4fCI8ZLaDBoILwxsA9gysGJ1aJA5ttMbLMshj/MWc3h8nYCBQAS4e2
1ECdofZYBRBEm7cvZpaGnPdSXqbtG+2cNqSvXZ0TBG78A5LQJ9l6282zOQGXmyBt
QoiwUII6YbFHbW28fbYrrM8+IsIAtaDxhLds62g+0AswfVlDEkspOjvnVMZavYG5
/3oBFHl7/DOdjjE7AdrmORDpDCE76bwlz8Bjps0f7P4hR2PKDrW/jitKbkGP6vnp
XO/78Z+F2bAUipG9Jxpvg9HRqSEenqa7DTt6ahKoAVO0m305gAdZ1pDRy/4ddDFm
WXAXFIBuStJada79qqGIP36Inmfcfqd96Wseq7IJs/PQHgfJEZ58cmmq+2tjr/X5
C5+9/PcCGOA1wlPsO/yRnScC/msicWxGFY69lCS0A84OYZNnk5+vrsyZDZuxt/9Z
pds093esbNBrFX2f5MZ8Dli79iWDqqtVRAqKVeAI/XECpIkyKc1fh7n6DciUovcM
PyI5/5qZ9T4wOSMyG6YrbSLlPpp9cMXixeUYeXjAR+/TC3y5nraflckUumG8gM05
+uEF8BLD9vQLTBk1rfgWc5AD3SojR5GmyuVrazypNCAsWtAR7kr2O7fWwdhBVX5+
IU3w+IcEc6LO0+c8jd7BuoyqxoSnoPIrkeSv445T9wnqQIaG5jTtjjJjKsgx5qPM
HDtVVh2Y6ud7YMvIMsLZUcot4XG4Dj7REA0ZtguiquAVMtIYPAMzFXTxpBLUNczB
cGd3Ur7ymeEAsuyPIjnW2Y6fKXY7Ba7aJ4fRMA8q5p/EmvYQWEbgtRpjd+VTfppc
DvImlaByy36ySqMXX+0BWMZIDwPM8xrv2kVu6BrmtW9r2CDhrUG9eKrZTR17MeeV
oGENHLtYDAgUjz9hN+HUAauRXk1pbZ2mDC+sBqwsj8j75xNQFenr/+fM3NjOxluq
3UyG9eNfwRFFV5RYj77QvZghF7D0g9WrF+1+nwOG22EOZrOb9mFm2ta/qn1PACgQ
feCuyc/n9i4eJ3APtc5PI+Ri68EpxiZFLHqIhx1a20Xo+sZoMih+0XB0BgsQZX4d
6sg7JevtshL9vjhjhsx+i982Mrm84PSYGnL21fkYsfAObXHAYkjNRsGxOvzILAtX
6eXV3xdfTE+tVM2WfwF4G07s/EC4b4jHG2giTMFaodZo4bA6gDJ1/VLuIacVGqxs
CHH5C3ky27j3ULUQKx/+xI6FKRu0ttRb2LzHaJuUtUUbiCVzpJwr6QwnW0QOhS+7
HTNkE/5i8QLTTpMcNcDLafrGkaUAsVM1IklF1K5I/ts5g8aeffR0isa1K+HBCWyu
OXZ41H1jcgLW/9Q4/d7I0PyuE3XUNEcz/kBXX+7bx70fhOOLOMhp0oqzOd+Dn5en
ot9iugyonFZ0xHQCr2VAiV44vCNK/5VTifTBNUAopfVrA1e7+/dX5nNO+KNWqwCJ
hiXpZ9dS+tox6AsBfqHlLoCGmHyzY/IJjFyEdflDxlQB16L8PTRWHmF9NDtGkWep
ARzPUPOvrwCJxdMlvf97Hm1QjsI99qmk6oO1WmOmn4A+/+t2vtJBhpetNKg3YVAU
Ugzo0ZVBiWH0A/cxc0zeYWEbzUkLb/vHbukxd9u0piVX9+iV9Tqm3SaiiiAqUghp
ewEzY7+wf26JmLhJ9GkTAliYkVbb5RCpnv1kuvTXr6kX8BN7voTZ9Lsf3Jjm07Aj
9OXh1LJToQFNSU0fQ3MnHogAjuWqO+bjUnS18ikMVEKCFE+nXArMrjexcKfj4iK6
3VP3Jdh6u//OcwV5FXsoKg7xV5sx81iwiI7H2ofAJrV9L2QKoomNcTLk2SW8UgUL
TXQazW9l6FAA0XjNlQggCqbRv5lrXzMCFw0F6UFTQfhCK7Ll90uVVgWs6Ji9iygA
JgLBEaDPa9jYzhi8LE7rPTpY9RU56yBs6Nk6WW+a51Xi5lT6q5nzV/lXPpeUM/bc
hAvpVvN1jReV0hT4Gr8pph4w0ENhiDj/2HjeaTtVa0uh1WT5lCEEIL8273L5K9AF
8pIag9lTtTNqizXpZqNbNoeMLStOOo5AI+ebssPhPgbtQnK5wIIGtv8l/Wn4g5yj
gS7kTF7e74JP19XH+pZ4j2TWzEaRiFwzcZLTWhk/AvHBn4mVipLKkehOL4n+Ou6Z
2K70AuPv+Zy0eh9egVUYo2dnMZTv4g8FaIXtaHURmxA3jxuydKpomtXtQSx8LIfD
mm/GTMacfuoaQY0j9tDa8pEXiLm0umk+QgUnL+4++ApMm3jNLkC9Ys7JPgk5MZ1I
hTWj392dT5AiDvgrg4Q3qDKuSD2Xf8osFtMvnJMHQiesU8H4vqlClcGn5dMOxmN6
9OSgB+Upbj6VFiKr6TljwNR6M9VniUxQ2mQfxpLmUvmcUp8Hyu83djb+k2OhOT8s
4QiD73XtJOPmeKSO3J5uw8TaQQVESuZcc1UalfVzswssxoiflnJocgx58djDPBEj
YJBAEH+1KMSqHevARsBBm3aE9Wf6UqqlSxcYxx6uY3GlZsc80GcocDK7uXidvBis
C31J4Sd6RpVT+WC7SQj16dYERJH8o+EpKLpwUPR80mbB7AYK8gAKaYvrIzyMAj9x
iv34d3o8W31dY2JDpV6Dj24D5DIMlFB4/kJh+kPHJ9W+P5DHj5VHohdoNzHkAdQD
eK1nJ/551Ca5gC2h2k0LtVYNedY49CG6bZQDGbBXFyl+GYivWYjXwCmbqorVl5b/
xLCMZyt/ketfNmrTonl51oGPbbKwVM79vYwDzarYmYlaL32u6OVeOG/xQofhVnH2
epn+Ey+XY1rB8b75EKWDtgBKIzTT/AYTQVt8jppxJJcaIiZWKMueruf1SmWsFmv2
2hoiL9Ob/d1Nak68t3aZOaeMpHvoIZkGZ/3/7f9OlX4enjgRb0Fkx/ZW+naPVS4i
qU0+rukB4N9IdBPnAtDD2ZadruSZgowOnG7F7NxMWl17hr07XkLy9Mzeo3+AV0nx
mMO9ktJfjQ2UDXGvK0JriP+hwRuSzqkvyERK7UYi5BF40n6CGWRQI0XQO/KFRRvY
mpN/i0jQrHT9LwDmFwROZgzCChDoKfWB0hX/kXUmH+8Fbb1uneEWAX3RR5tRlhdh
rnAvvl7+1SgYSdrgMotNM6wuk6lu1KyVhyLlYv02kamSZcaGz90F+hJCUH0Fw1DS
WLxL3hcxs34m1HoDpf9zJl4jq8U36RvLqGYvQAoAArhTpec9+lD4r5EzpK/qer0m
IfACQ4iK7gZzRel+CUtWXqeb9kted8xTqgoahgFAz1V/Ut0uvGfTGcTHG8Kb/hKg
mbAX2j5f+HsBiqkfIR7lxtcqjnPHIVHQCJi094TlcLubSTfV9Ogdc8uJbQntUK51
LpXdXVTgj114B9lcz/8/vI50RZHbyxNJPsKD3hoPGzzZG/odu9sL4UsOMytS6wBw
UiEVK9FGS6nXdjTPIavC99VWJZQgf/F5FwOCZ72gFTOqzpXfFY1wEJiExyeIoMP2
qt6E+AgEIy8ffOrQPMaIKh4Yr0oBimmRUyFyOm+itj485obsbqM65A/U14c4hoEq
iCN3JTXhWohP1jf2Mz3FyDHWjmrZFZSziYeEsqK0SWn6svdKNhyMws0V7JpOoWNr
8HremiAlXwgzu6RX/zWV4EkKorrEQg3SjXHuayLTri8gFaPTEqjZTN7HXxYiTSu9
mwEZ0OydisC4c7uvKCcgzizBZfHvaeFmMKLo+r7M7f1QUBkToG6lChpy87rG+3Cj
TtYAye/ae+PnQlPaLA1rZSpuefA4BmgHhSqGK5C/jd7LJfvWXS/1C/CwCPZKF/qK
5J4VhTGv4DFp4yXRZQY2/3LRrWOT08DlG6LnNCtRvyZ1DyhjCX3lPYQe8ekMzS4Q
C7FOAXhivJ6QNp0HwuaaGBLYV5EkEIdBJVImdVvoYbt0d7rCH3MiPwLXVpEdK1rp
P793bVE0hVfs1reF2y5q1kv2ivL4pAs/Hl27D/bhAoywqzuKhI9tjFU0f3j7zsjT
D+1tNZbZJRyggGO3XIBe50l7uaq5rkYaGL1TCRjg/tSKIzKeugvQ4AD4w79HIMd8
UvHtt8BpPMlwch+0JGqOw0w7XWTxSVofZi7P13S6bc3+PfvW6dPR9GVpGODdagAL
llXxCQvsdOwN7sIbOi29vkzY6uTEeupniCWK2+FCDdOhH0FF9kwfvkVBLvn+sxfe
wa23ZA3NeUj09mCd2wWgolM3Lfmq77IqKOluBIACIU5Wga+Iq4XSggk1s1T4oHty
cBfXUH6VbiqFM3IpcW/lLsTsY+V5UKLPdJ8QaiQy+CsXR0rpuoPRb36fH30E5Fus
Ckigr2K2t3eATZMzo7yTX2HddSvSfffQBuoajb9LKsa0NJsCGjgQsm7F2Pk1jpa2
vd1jesGtvDep7weRJ2QpwvT7F80FqeamJ6dIW85ank1yK4Q1B+pFG1mc0YbVTgb8
PVgBEUIYVVH12qKLMtWVSEHdhyg6AGS0QqZEjv5Ui8v8BjlaydnkL5xBP8+L+qdm
RaGFuXWsnglDlQtES6Y2or+kXlk5NJMncXhsnT06uSuB5DKxGMeTBd0X2gjNfu63
MGlSOgX46zxslP/3KgV+c/yfXF0EwqejVWSRoL7B36wX8UxLMrsRnO/LhpxJydg1
UiKSfKY/d3fs5Yfilc+5hY+2TiFVK9eXc+6frknl5Z/HKocrV6fvEmzDqtlJ8Auw
Y6kt4NJY7XwDWtqaiTCKdErHvtuRpuqjh3h3t79z/H7sochZeEqSn9WbPNhkwKce
goGaBKEROud/GY3XwNuZYEoUAT5Hy8wheqnbI23DRmFfgyAghP2VlJH3HXSSiJEZ
ODq+0d6E/0609lsbvjQ1s0HqoCTW8GXG+QKwqiZy5Z7zN136v4d2BZZFMSdz9LVZ
TBihvg+d1XATNhCX2RttF6/MGT/b8VLicHKG5i9/vFxydLEfg/VtA9ImHlk01YgC
lQPKcl0Fb8TWhJ3x+k0KJsivNE/4EhGf2QvX9oYWAsvgR94aBk8sB2DqB0OV0o+q
7qxjBb7WoU943Yf4Gy1beNMAZLsbSMMxb9HOC8poO5xtoSWleuWBhaozokq6vwvq
Z5HEII+m+U+WfwY1UgT5M65HTtfWUG5p//RtuHSZEQ7rdCPJuvwGEHb9eYD+C7+7
zlpJ+H26InWeFrhv5wZSUxMiIuN5fGFq+8lWfTkfBMwMZcPFNJ9Q0mU40GfSU0bp
cj8VuDjr2urHUdtMkyB5itItYqCNQ0kEL5ghKIt+JKecugHr0f9+8yfkgltJTf+d
VDSUDsf27iIa8PaT4uSSthy/c4Xl5BgoBXt3sJTz7f0wmYyYwJwziVfZO4+hkEDp
ysqxcDcvlCqQCPBLJFYcZOBrBW8l0Rb+Ay0OVYiO3KyqONbVrfTwtRpimE3yOCy4
cA++f4+1CZu7nivPNozMFLLzo2h3+fIyD5MJDqw4kdxOT5M/UM6J+43ybCG0boWP
Tg/QJ6r4q2NuVShyx3vWhr//C0/Xs02FNXYLPYViSXiUtxriGeIJCcSb3P3iYyVg
k6+fVCaYxZh2GpC+iHzmtEM41C8dVFWtBME8W0WjCyWy0fohwSSGyoroFPkmwNr7
cJ3GonaTSKc8ciqOOBgZ5NBBRdAKAUjFLaC23bhWdr9IWIQ6P+wgjt92lD4YIV5e
7aq/3S+Lc1/VbBWsA1cHrHKav3rBp2Q7hxPM47HONQnRQCsjfVem45+qgPG3MpMQ
YDOxvFNFuM8hARGUBPVZ2hS3aCWnJQnp+ujvNmXBJJ7HMW/gIKEE6+fVrf4ype4v
6CtLREScLN9GLeHRQqlHObLlEuxexcD11vGCjsVKPqs6v41VSqEhDBxPSkfhjbn4
Yq9BCqMgUNrtrYZ0igccLYeDa/PBr/nSGF/ocSebr9S9Rku+HC9yDvKeEBcVpSmR
XD797/dlW2x0VW/Y6/j35kohn8FQszoeY2ZT3vT9J9tT5kN1lVxuLQalPKAirJ1b
bJUBMju7BH533hen3+WN6rXcU7oFE/Hj+69RsX6wXXQTFYBaxTjqWdteo4bQQWhB
Jfr5VP3A6wsP3RM/VvEr94agO/w3qV5Gg2r+rUwuFS0vHgje9LvZ7hIud2xFIpj2
kBxhTQ1BU8no49q44k0Dnj5aAa6ZS3+xvZSqvASReAEh6p7f/RMYjJKLTBbomrPU
RrhusGO4TUvv0HSJuMw5/2C29l63w9jHh4LR3acaGf0/spjkObM/EAdgsLIRk113
dwdtJ3uE46QvYv7xPGuDfM9fHwjBZZy9/8RgwQxWSq6pPB2g9x++lL3xXZXdmprN
RtdjbxZy4BZBVzAUYBCs73LNWI4QM18oZmyovCrAeXQr7H79+gK2sDc9SQF6Dknb
ErghtKHBWcrkQtqUOW5aUVFUgPrpCVpmVk1OXVqFEKrlMXpHKwr0nPoQGHfai4Bb
vY85KvTAIv54QDrBLoOIVKnF6HpelKALEu/83oEG9Y+CDvqAOwG6WduM/DHRRHM2
XRgkMOmHdZERzxMkHC8jrE7ZzMDafGYq9LOvbzvOAc0aeRa0KADRTV/76QGV2jLx
QrhxP/PveY2eRq9eT+IJ/RWfPwfXyVuSaq0LGUWf422Zvd89KO4SPaGKRHIITAyD
1thOdiRdyrHr1MgdYTIWGuV75cPuq0bQIjKhJ9wZY8XRhuH+Cvl3dwnYuTZ9xooQ
vhb2q4JZyZNRp17JmMd/VnIyahlvxZk8tdMHVlBqdVBVOV/sWBHFcMXBc20oqKIs
Dh+3tBgsrW9E3yX1grXv+MGUo/nauqyumoQC8nZpKiozmyGNi8uJP7L0kZXDCtQy
7t6wmBC+02wU0phm4HaXuFrQHJnDoIuUhLIdvjMaO9e03IPbEv2DWts6M/elpq03
bI5tLNiNeoggOFBKsngz+6FjrSxkVrfti62BB9Mf3DMhz98TusINoxwnfXmHqaZA
fM1+lk5YCIBW5R6tiR3icqkX1rKUx6XW+EKAz3QwyMz7uNIN3gPTRirVhSHmm8+X
w1rrLXfDFBp/ivyJtVp1Cp37AWgfOkoxNUoeGypvzZkorXKUAY5kT5PFQqM1k/VQ
onzr5OzFUWyrsUHKyxr17EGZDPCv8+pJoN9oaWa1wikTEZ4ic8QQg59qeGtV0Ejt
IGU6We/vJDYEzVeQGTo4NhBLEVEk5HcB3gVCfmm+3e/yeDUhhPOHOHhnCnCyv0B1
Z8FeyG0fWY/4WSaBzmkpv9zfjB9Ea6H0cOX11fXFMg6MEa+bnKdxzetmqJSMaY7w
tmcmMlJ8HgiZaZ49v+jH4qX1wmpJs4yYkOG2MLDnnkhj+bN8MF+xvZlwJQXy8TjY
8FlxPdMKapEJiaKKagOvGeF2hLwjJcTqjshWIb9GmGUHwuvKxDDRgBgRp6aGCHIf
vrgORSMJhecz0IJjQ0WM4dBAn/t9x7MpAkXRh9mLszlVk0DWKwjQ3jG7TOz1XDlh
emM2JJwnfk3317zrXTQ+prsCK1c0UecfaH2ZaGU40cScpxQQvidMjwYLFf3TUrhi
HVdOOsj0cCV5OfEzLV6EXsBzeGNuTu4z2ih38xeP76VTqpv2GrUmWlYHvy76uQzY
y8hzbY4QddHlnWNT/aYaM7NF/5ftmhbWneeT/SZ25zPVn2L6e0o4+Y7RawzIIjWi
f1UJRFWGpTIkS8HZvIvgi/e54X7PpIy2sw8L1TFcTnPNjkpTwo2VvYsHpb3MLZJC
v5q/t5ZCS+ycrbWQxAqVAZEqUPEuOWaLfcFHqvSvJ4var4jMvHe/n3pxZA0Kyh87
5qtaECCy0yQLMHLESV+nGgzbhRrVPi3EJnIxQQfJrhfi15KQPo5/2/nWEPFrNaVb
IHEVX4V5oKiq2WeTlGaODIPGaImaAuguldHVHWPfTMVbeYFEgf2fTLlOTY0x+HJB
EntMLLkfnZj7oI8pxCqcyw9yQHUVNpFF0SLNq46GoEWgekRPBGHEllS9av1ZKRzC
Y9MUM139IP1o1D4RdkBoNpERrIPJ5MNSjireGeEL1vBfQl9o2ONJLudsL2xbm31W
5GCPnNB8JavHTc9swMiWozVJlHurlP3IJ36UYgvGoV2pfkCey7WbbM2cHOw8A9lJ
Cy9kcD3riR9tLIFTZog7QdrqcRBVqpnVeIrvOLjaMZACYErUVpD2HZcM33nqgOsN
UYTgpOkKqR1GG3bZtoK43MgEJxRPmqbbjY+X878sM1Z0NGTHltpphsdvr59LuLjM
PVkKcRrcmQTT12yeXV6e5QsDQgZCF07Ed/gw0cagYWWtE+VyXCQ9lY97/fmK/Oj8
Mv2nXiUqtQh/QI1StIe1baSPhIoie4Gr7SwW7+QVcbBeovqhdFLtGRp6M++c+vd5
zX12n2DFFalk/TNfMoeCS31qUcIr6dxuzju4e9cl446WlBCW6Juqt4R8RMFc/+ua
v8KrgpqPubxImteVUc+IoiRQSSOpXUbhvROkmfgbkFOZsHyoE7tDVJbihZCmBZWc
Y9lm4U2LfrLCbSsYlQohxTq8VgCfHxyKceK7GLMVgFAQ72bOHilO8TelPig4SfYq
giKeu6Ty1RXrJsCFCe6CiQLQQYQaA+JSZ86OyyFYDb6wV66qKtyywUzZgcqMYE4f
7EI1PFiGZ9HFn3ZFpsmo91A0U2R3qYH455JjzuT7OjaaYw35BmBBmdKduopVJcXx
7CDG9IPJvzcAVP32IsM2qrhi1BccLcUE75azg82RZE3MYd7kWD0ydtXSljIyAS/R
9oBxSDGNcMDACgH84XGAjY0b3idopJA8x0vUoT0UTaLlNxCF3WydH+x46ijTFX3w
0g6ufCKpKvL7inGgyFrj4QKanqfWpIObhuR3gFHunwvuzp9l7WJKnKa2LWRsLOGL
nOZj2xxaFcSf0HWfSZ1NZM9hM39edi5F6Q5C7437mVj+3MJI+F6ApS/qGZE7CtGB
ZHvcHLVQPJsppghLW+Q0zCGqR7LSEH7scUXaoy0/prfn9BK+UxV5NsVqoyPsiMmw
GpJDUpBewj84zCtVnvn6gozNqJi2NfHgwtaCGWP6V7NHRnI9OgQkOI8CBVx8+Twj
6aHPcf+ARttkAy+Ckuvzykv6OguyVytFD4C1j5lTx/yE6qTZG/iSR3AckmmXK79S
5AKp04hJqhDYEF+oEW/988eHdL9qonF/IPhZFYYRJvGpLACH4HHucJMc8MXM5hEP
eQla4rIKGnWno+jA3LHIeJuM9gl2K/mGApM6AgXYigQ9czQpHJGkFochCqPnSLpr
Nl/kBjE5XLRwq7JDUYqDk2AhLhui/ml6cRsAQiYCXARf6//TE6tm8NYYcXsrjntd
fLqUuggn8W3hYumbxBdMN7FwfsndvgxMf6lj80opxCBLvvX6YZ/nmuvtXyrRhzr4
ken4BOH044c8taviXzuxLZ4GHmS44jj2z2O6Ca1W4WJRnyMbncMAUhsDacL6Q3/t
McbpgLDymL3goJKlzUcb2obk72Bb4VR9wiTTgPxgP+/W7siN2CUWkP0RNhwDuWBH
92gIm9AIRqg+TVMRqwT7ciRTcLA2r/KkPYQEan3od6TtjkYeSqXsq0AHk7wPwBN5
dUmRH0QTn7cl71wNu99CstHNS2p5Ibo9W1anKwW28iAQ1U1yBlvvwxIr+X4cDeL/
m9iwGgaJwItNT0UQ1LhGelaadFAso8gjF8UmrgzQMteHVxQh7BsqRzjL0OpQohd3
VOIqzC91St/r2vvIR7r3Zw17ZQxFkO7B04+PsbSe81hZBO0FyAvO2pJjSwRzfm/a
WrtIfyborTM+/BKGyxdIL5cXG83sb3JR4DzwO/VFqAoxbjiYEw8OvBaEHD8pJ8Jo
Er6R3XuWX+h7sMp6d8sQQC4QzG7iXDVZJavt6Uou+nAiNiFKcU6zTIktfsGQQqvo
iUv1thtEM3yQJtGX8YVz2B0KO4VSp6yrYw0QtJm7Ghh0Ch1vOiSBCtIhV0ImSc6L
4WBEEtd+63UbkJf4LRqE9QFjU17/9/F1DQOQjFa2dd3lwSvNpRV/t/GJnKs7K/eE
tuC7gPD+fUVXgfe3g7c2cdBKbFB6NLX+1MF47nhCmpunKfUBCUg2dxDgOBmo3gXr
2qhDb3xmD1ERqqyZxHd5Qh6lTfE9jY68a/HofLqtTh0Z3sqcJDZk1eK5spXNfx1G
LNWDpwYNO9v3nm0qduhGI4ZJl3xcTb4cCs6LbdETxkdRdV6nrbECHzK4an0qwDbz
EPljyOjABF08bdDgz47O7KHuD6tIAwQWuJh3JeX5jfUREAE0KlDrzjHDfARnPAkP
gLFJ41gkrxgBNSUQENN1oilzEoUV9fdY8reumRKwOuJIOcwGseIHBPVnARHn4pOP
raivVgIwdFwl2V28i5EcGVcBegAFB9kWtisCFdjSvjrmFc2elDubA4/D8Wgv35fy
142rbxYaRGmqKd6oQGu8I3O4FnmdmDTd3ZbtebkXTrFluj4mG5cxF94Vv0398Hbx
RUp/hsXjdU3SfNKUCk7miwMJHLZPPQGNnF5+whzE/vAVQH8fR6HG8vW3NUk+NLh/
KAFLOmiBVLSCkG1P8SIqhM6X+iz42thRO2qLgpqkYTUL9kAUV3YJCJ0II7J1lfXU
KDVP0S+6+WxrnNZLC8wpiLpjgTh+n10eSAgdDetfLzwMvIcmhO7stbUNR08rqIQR
LeDFt8XNhtil2K8YbAma4jeRhwJ8jaVrXvpO5gb8XzC/pykot81w4Vi8WjEaeow3
cPlRWibuLy1NsbKxM/D2Wti5+2Mb6g6K2/l4hdkbkrB81EGDVTLWmmKGTSfibXw/
uFX1S91/jB1jNJ/zP3qxBAIqrcL7/4ZZGCi6eMXUAIS2yQDD711+xRbtg/qYCu9o
/mQdFD9tLOqDUAZn1aerIPKJtKPBAmfADOfgJT+PbgPHapmGqRkLwAUhxhwFAeDF
DX+YbByDekUgsx/mxPsQ6j7yEwmULdRBIqZdPbi2VPwbiTZI7DqRJzxxX5s0tV11
us+4/+tf9xSufvE04FLh5KkvK0rWz+ZSp77k4k3GANxX+JxXq1kzty/PTn9iL7xu
ZF3g39ZMDUKGbfj4PuB2Ratc66+3/YT/UzKJZ5RFKmac/GotocCFQgT600VPV89C
i6EtLa2vK98vz+T8kvVkSpYEUFEdog42R5NqRVLxNrSGfQyOyz2me7Kn4+yejQvI
Et1rzo+IEwnnvPcklfeODTMFIb5O9GDUf8bKqhMa7/0hwWNziZtkmu7JdQzM6XJJ
FKJVOR+PjG87F2XNe1M8oqPu/UUBBPrqlfOAHEXEwt5mU1UZjklfjZPme50un2n0
CIf2bETOMJcZd3RdU0DMryqbAGRKJFicz0cF+DMp8fOPateTbk5zhQN00AWpWamR
TKZU7UmAbMHClv7GZIrBhxanDxZr4R4FfOQsd+5/UgU9Kb3V8HYb9T0dEaFB5RzY
L6kMdfEOnmboz6/U3rXvfppfJs5zdut7LeGjaRsVJFaKQFzPakQSLWeOpZO9KQji
TMNTpDbvrCcTfZ3NZTnYXzlv/As5Y7B2d4deDK9+hwZnYCu8lS6hHejau5DAzYUl
ku4V9xxRty2mAhxp9WKsEQCSpx3x1ITFqRoazPUx04sm1ALZbxx4e1wdU9SmklRS
2Sby1bqDZW2QBFLja2gK2NZfwIcaHtUOVQ0LlJwEYXcusq+g6VhcBF6OW4zXvu3c
2NHrknhsXezyuf2x3EaIMYmTzVrGA9ej+FV9BH9CHgLhjtdkoe4MSHKS1UiERxF8
Col+h9dm+s6BXH88S0nQ4qKh0b+GzyTcxBuw0O9IGrY91JQQ4VpdilI//KG90u4T
Bd9bXIT5BLWmrTIz6jtJID3xiIdZtr5LbBI5IYeRdRCPntrfwJob1WipzABUVz1/
EwXa6nssRXpPvIDS0p24wbEUDi1Ksfn1IbvX90Bwbg6XMN1nkI87IK/WSYdU+PrY
ENJPvcg+4NTLOHU/VEAAORhmL/OQy79YOYhJ0+dervC49A4Tk+X4Q8dpCcUZ8bqN
7vVhtleA9fIn59mn//1SxdqTTMkjeaUvrs1Io1pgVBwMlP0wWpy5f661y0Ak0aIS
/4YlC/NOoqjXKeMuxmLekvU/15vAcSfNCIF0MlBJYnG/M9oWHs0JfTPy8CcBFSyP
QfnupY9hdzA+psd0hRcavjnRbbFkfbGVKEH8okYIEfZpdwv/h94A7CHrbnVBkHeb
/NIe9AVyKnzN4/CTRFss6T3xH0TVmvPDpKM9IE9d9IlW7s8R1CVZZdFoitm1PFQ1
zEqC8GK4BX4vEYBv8Eyq7fLvvJWH+GlQULumn0751j31euJsxFXoDSyH7MkVOBgH
yP2lL1BoLxO5jDu5fQdt/OX7QvpLRqXd8IqCn/30b72gFyfgVeRyF5Ss5TuXRwf9
lPUF/SCCcMGiupcXYeZue3X5AVohHggIklmraNm1Eh9pP280qPyISjF3tvPBEB/J
d3pIlH2KJURtJnaHanOJINFn36F4/P6K04JkMHGxd/PtrenMoSI1lW5p3tshjVh8
YfVS1J1Z2fU6Z+BSMZ0p5mGEx7yQIk3A9taCHuDH6uEDRxnw8jx6kJCJboq2hoL+
ZFqfas0uyszJErFa26wlqs0rMhBOn0gdrO6tAAnbUj3Z5tRO/a6Iz1J6QHxZu4Bz
urkzUTmriMLBVKAcf6CawI32Gj64EUIBoaIGVNTamPCyirwDc3GziTv6fAqrBlhY
xsS645HOtCSpfG6EkHApLPtj3lA0r2naDPMhriIsl/c0364h/+U5YFEhBz/vfxTO
Xac3bQ3xLCzoxEOjoNxxOsVBs3nPDBRFtInZe+D9KGXdaE8ATKLEvAy195A8/WJi
MjhSNIlV3FUCy0wbp+QHC85euEkX4E5niswOFfKanC0jA3c9YCYmkDp0vGd9PfHZ
/eBlm/IR3xF/nxu33nzR7ZBrgTOQXwFVZyfAPjFgQzsWitUGULYeiigICh2tVvmH
1nKR2lHLW8tGVq9536tipaMvzRB5Q1LoU1190q0o0xT6Tr3r3fOJCxwA2kswQ/IY
kMKHw3d4DOPtS3Fhb5q3R0vpEs4YEVMRqouUfNfUO6TbgQDLqkEyZQhVqH2cH0Tu
lWA24n+zlo8NmhVcL54rZZR/3T2skPDhlkW+PZrFEtHHkVFmSxJ99cnt7kSGglE/
pZABASoMoNNWxBXGWOtJsMtu21o0v87rb3D8IuT/DUUSTzzHG3o4g9t5V1hT2t+U
Z4qW/BMRTB925oy1x8MCa1JZ98UEM9BEe02IKdR2utVsMvyiJRShBx1Xvjob4Fxt
CENbGHRc/db8UJPf8iUiQXj9KmZfPr71tXT7kjF5LauywIjK4xhmeJURVWGDNk6J
/5JGYPFwrjGiYQ1ue5MLxqgUM1/EpN8Ny9fhOkbykCe+mA46OHD78LHqgdgGXUxY
F+c3GkxRACgdIuxymtMCMa6mAvTDgPPekSJ2unIBlH8Hsz7a/ws8nKLUSb36vqVN
aELIXPQRu0J12hDn75BS+B52RyeS9VZbmvEwr6zQqWF34tbgqRD2na1060I39ruz
BWVUJEDi66FhBA0GXcTUu80VdmsB9KhjYXvEfcWbK6kkK6AMDdsXqC5FbUAihEZk
upUrtDSi272X72SL49y4gPAVSaN5VCwY+hPjO+17znUemIjUonFZ5CTEaZYyPS4m
9r7DcorqZAZppj2JnZ7azVMmvhsf7BgwuUVj+1nQJBlWH4ne/BXJv1dak+sjJLEj
ewqF0rXeEOEn0vOQmC/Kmlg//Cb8vobn5mC8F8SHmi7cErjffjKXtkC+TEM+U5n/
Ze2FTwWy+2exFxeiMGBT+6MNRFZ0XaAOBhEr6T2ag+6RjldqJVeMprlIstvtJvCJ
Cp9zzD8B4Lf6x7SFTvtChUw7KcW7yMSwyNKKM7BxKrJ0azZwKvRJTJ8f9Z3jym42
NMVpWVnND7XA8uNndk+tRYpqH1YRquLyvdo/fKhdaRRL1SD3a9se9bGtKqk4ANRz
OnxjL+C/P9WTTCLzslbUvCJmeJYOO/o6TBZXO/Wk0TShyU3mWL9QF4JgF9MyIiaX
XGO4CMzR+UNxjlNMx1gNqjgebGjoKqE7zR7ssV3zUWtIb1ynFDNu3PmiWFW+zw+s
Yz3/tKh2DIBzuhGYmSrZnDAeraicCWhjekX3MsEL/yyxgnUaxqV1BD1wpuF+xb+e
mPm05twxgwd+hCekweOZe/CJ7ZoNqJuPjUf4FYSV9c0YOgO4d0UVu0s0u+2IeeoQ
uIm/MZ+FM/ullHTo3fiogXldDcKNGOsJ2Lfwy8oi/VPKDWaWm772pixEEa0A1vf/
A6fCcXTZpf2ceoo+g/4UDfi6Xg13xPwVrzE6UGXaAmo+FLLNxkUvOUfRRIGYf+9z
IfZBdQSKrThMz06JGYKS5YCnLD1DLPFXNvzeheB8XQbZ4+r5LBAGPqmgr6nFPSQj
oVAKI0pgPTV/VE+bE8mmM3jtr9o0wYcjjCuvMXJkxVdMpncyodR1U/7kxP/3sO2y
TAnasiREnJghFXrT8Zs7LquGvT12KoxRxIjDyF1A2NKYC8IM4g5gvBOHjcrWg30S
ql3Jp14UY58ttIe0xBYfx1g8Kk8rJ72EmUXWemmtsa/tvpnkZ62JTECph3EhNX60
CbjDNpXo6y8Dg47tO75gzXRRqD9PHZ/a19Z+R9xmuTgz5ltQQiybC96IMqLVWvEz
0pWGgU76ndn05KOOuAROIYMQSn3SB2W7MAwPcb58gAyWOWtG4Ms68yBXWtuYPuI6
hCbz1AhqFXrQEQZ1n02Zp5fskR4TFJcj1PI5ZrB4Lms5GNsMuCB+QdclY9f9HK/E
Ly5IOv/KjWbwZrv7x4z/Q66n2cx7XFfnmfLS80ZNI0RPDOMv6JHpPWW8eCyEiCl0
vOUCCzP9laNBcK5TJPjwePvUrQ210yn3EUc98nLK0lUtf58+uPXqkzf+Wx6LqyC9
ggQfKqB917U0sZFYVh70GSuITvxiKZhNN9r7PFlZUQcl/kx66594fLdYVGlRJpVJ
ebF0M+Jt2jGP8W5Pf6Fd9aD7vXbREt65x9OXKzfdvKr2meMnfSp8koN2A/rECfnw
qRYtHiG62uoe5iazRAp027LGypLZD3W20BdNR3WOba0mjy9zK14nPB5BOvuijN6j
dvENpmraMsluGK/rJdNo0p6MFYM2h/rSAGAZCqshq7B6FKgleOpnK4//D6lIJI7o
uD5266XvcNDfVPDJY0AW4rAotjV0AztWUnpU2lNB/VeRkJu6tCs85JM5hwe1gkwX
PuKHG7Gd+4v6okmcm/hfYbroFpCVYBC4kGCoVv05+AyIC2/Ueh4BQc9RNYY2qcsB
rJGLcR8eGFqoH51o4XFi11z1toZ4eOYAc5CVKvGlVHWOrsR2uW/jYOw03GHkKi0W
2mJ4t7QGcoA9vIVn6ZoDWIfTYFy8UjRMouuuCAaBUnmvOc74udMvuLJ+ZFYFQK/r
NMpA/MW9oXGtS1KYLK24NAfZBp8lrExfRJMm91G1v5LmStt43yBXQB88V899Gt6V
VRvNWtsqZ5YiG+4xhhsLzi7h/gQUEbfjXIr9ThOhiBZm349UofBnRw2HQLKGpP8Z
C3A4UcoBPCS7H0n6k1J6vm2/BM00Zb5FdupceuY+4Hk+ZxaARgoqTF4blOndzYEA
wVx0eTkb74iIm+zjOru+r+xzIea9ZhMGLUoS3x1rgrvA2SVgTsavSP17l1CbT/DZ
LDKy9j/W0rcsquWVVdsIszLxMV6i4gQ5nKTXKxfH3fMRb94C0NVBSRgkT0B2S5GF
ICLygSdgg5DiJqgDAqku+Rez6KyaUfJE8I5pugfrNpv1uj7/+n1piSSQN5iV1KFG
ZafGt3vJE699emBRSXt86EY9ijLIq3qFqhW8FqdwUvndfCaYKwrGqSicHa6jQTNi
xiQ3VvAUSr0+olLuCRlzuK+JekpR7u22Rw8RvEeGVqCLutM/fK31zx0EQ0DCS0gx
PicnHT7NSouMtHbeihUL/69FeP/0JrPxAB4grGWpM04/3Q3lnib+HdRhSLBFNSvH
Ho7m4+Q2929yaq7xL66uIT9l3/Yrzaq0rUonMMrn3QVHkcGEWrB98UreImXK9Hoo
VR8Z6uEY6GX5dU5QU2b9EDYEZtfPrEmNq/Cyyzdyy2mpNZfx9M+Cl09G1R1mCNxY
IHVHBhZV12x5ZFw7mTVqLeH9ld4LbRwEh2YCRqPKqrPEqwGV64AgrHH1tU8J2nDr
mS7igCMRA2BvOipRrOu8yL/+mYRt2x0TZ+b3SWdl4gWmfDDCWFpbu/uEn1+0chZj
gj+4/Zdo7o/ATcfgTGKDtRddrEbx+VBy9kShl2zloevwt7v4nUAWk8wGgvtpV+xN
0B4JluzzCeadK00hD3YdoVHBO/RmwONA/r5Jk3h76jDl1UUN/tCjeAZrV37pCEE2
0tXka4oXZ74s9abPo/lbCushedSjGsDG5HGaEb2yxrShj0gL/oBtp3SE3NbebV7+
EAfIHd/0SYpbLwEXolVZNam73k03C+56P88W/fhGzSuGn8EK29b3HWaEgpOYVpqJ
dgbfcAKDd81yPuSk1oPPCVFd3b7XGNuN8hCfThOvv9v67D1I/Nn+RR7hIBKI2Stn
snUwtfxcrcYKQLMRmgrjaVIrGCFnOJRTXyM/f2s6mbV+ZXMEE1rQLJYTXenzrce5
jfMLcv4imKBGK3pKzJ5SX2mNY476GLNmSrgDtAVdYoUQpTcYRAC3tBLF0HL+HD4u
DeNiSrXv9B+hHD2JkTUIrsOleoqMtw04qWdHGxez/6zjVoXFX0CoBH4F1uuC3FUX
8tLItzEBdkxAjQNRyO60QtYB03GjH1G6G6pI59Wib1ADx1JCfqK8NSj1tEyIZ/FV
pFiCGjjcaCeciRflvt2lYMIoj+DcTHp+Q1wJN+k8RgY7goQ1CDSFwGkiKp07lYfu
UDMM10Q+fhNkxrHk7miEDizTTY4baCbc4vS87tr7jqmx10W1gTmD9Vc2gP2zqmUI
yPT1ZXp6/F2XExOcHLFmD7Ac5gbzE1g7aRdO+b9/vxQkIKiljWUPrPNdAME3rxqx
bTniiCdz7xS9fAeku0ofFqMcINaxu0tfCbIJObXdbH3ybrUUt0PkYVUX2Y/W/bZl
bLiMtg4qfYGa0kSyl3wKk1MipJy6JnYQNbUuRFc5yl2CdqJB1uMx2vZjWwDz6AVb
kifNDLTZZxg4LouvlrTUuLfW7CHFEWxE3AJ/xTnZQBJEv/XHoogkJ8e4HluywyMQ
nPbW8MqBy5sET20QBE8lhzHwS5hx2bjqOqJ+iYiuRejvVOtYNMKqrSexeXAk0yWk
PZaSLyDjjwYS24vOpXBrDdUoZX6X4eAd8OCm7woY2aqqwMH3nliC3fIqzs8ShDAD
yzbR/8LLts2V4XScZSj0OW2KjH3hvRd4gx9fydaaslBs26APvRXE7cgXo7dQn/zu
8+V1zqO3vkoqmivjlWWTDb4w1ivQwxqGK+lQo/ZSF5E/IOFA7t849uKVzX7UtuMm
s428OppilO5h47qK022SRRVxtKR02CR9jy1zvo85VSMYVe+C6iuXQ5bxOaLx4yGc
ydWydVGMoz1q7V/5HhuhU+im4OKlXVeX2Bm02DMjSdwv7yhUCwXzOSfCdUO+ooyO
927CUoZIjO3Gx3HHuUwhInJXSzbqF0qgaGEY1VqicG4Eo2oJmbhlw8HfbKVnkWDk
i19ae4x7cpdXSxhd600skGNSiigb7sUUL/zbTTbGhhtUDhtvEX65UWSQ0l/BwmZe
ej5GSQw1nZRdA2/jmyb3SMHUtcFh92jValiYiPhq7ZenHRWeJfnNWdybS1K0P8mT
AZhOqvpzr+rDasmJ+J4/5bpwlzaJFpvSCXWWPPyY6HmjDOMeXVGjvmWeWD217osF
YzPdmpdF/MjNlh4gaQRjvZSlc6Zzll2ADz9EeFnn6B9GP9dojIJ/kdBwuJ9c0qYB
wjDnU7QJuD94nnkjan7dwG7i6imqAptZPrvMJIDSG8dVzdhJAK+VNLZeA17UskB3
X3O60OS8/ltw0VQnbIa8bK636rbdrw1cEAZadZABJFtludiR5QjRYTsOCnMHDX0G
wnF8mLC/N/oLpUPI44lyAeVOMxIsTyqCOGy1rnWEA42F4OfN0bfPVruJoNuBV1Ld
eRgi7fuMHyuGl/NhFiLX0966XUAs+ldzITPwmtIif5bnwGN5T3OOtpMqoUr5HYeB
XSjOWPr6L8/Oz5CONdtvrh4NT0Qoh+s6Ho2rehAArOeyfZB6Eg6TijRq83efR483
JLvOATfT1oMOibLn0HG/yKGOePYsfceX3f7R0E1W75oV0n4LeQWoYuiV7Qi8WKV0
Ic5FzObKhJUCLNhyyOsK/JFXL2OSS086yboqYj5nH5zMbRvIDIdsvRVGnxLpVzJj
BQSgoQ7lnVv7hownv3apz3uW7FJXIWIYoR3C2A6a32q6nuND8Mqvnlfi5elfw5BZ
JITk7Lgc6uXz0HhobW1Onc3+6mEuOVSQNlWZRgei1YtOSBCVzOWf5WE49pT2tOqX
pnMeeCRjnm0kvPs/KPc4Q+R96FvWdnZI8XHMwSuROlfKNqbLNd62hzQgM39R8Xjz
EndZwWQwiCs3/ECs/MXGNfkvf/GcZHZIyHb2HFh1lAWefLsF9dyzdTqhbaWj8puP
pG2Ae+/rynVqiDYI8gJef67nkJN8NiKlKtz4hrg0f35rCNgc9G0swVDWlbe3HPph
01EAJiXn+opG5Cb7iQTOIZrtCkSOZG0I3SLoH0l5uYfdQ9NFEPTJJ0YPXEpmoC2L
igCjz4NU/7Xar4hZStGZdhfkOW/oRLfJGkis/5TrPmS3w2/+xGUt1pLWgUuJci17
b+cYag9o9ETTWT66j2GwE75lGO6OJN6707WI4adATSbwWrXY1MvNEmI70rzHEKvG
2cF4zmwYilDcPbhuBiY8+MqgXmpc8WMbttf2luASIOD91FTMVdGgB2UhowVQ39s6
CA5+q3WaijY3xHEmgMkviZRwie2nFU2+mHJd15Jszk6ZFV49wbR+jMSmxTgApvcX
OH0TWeWVEv6eEdXRYRdjKSYZel2iQdX/32dB4VtHABr/I7jlvbSPUsPIA2vmovjF
Sz7N2svov9w2WnzONRlG/JJFY27vMWaTPnLEhuaLkV83cFSq/4sMWyVJD3uD7Qcd
HAzpTMxg1eTjaKB/ln/Iumua8yuMaWVSo3ySjnOUySLxq4WSOgtjbMmHlIh3JOzv
wnc+y3qWcHR0hBzzHTDmaQ5y6hdyUIte7WLs+XkWJdRfMYQqAq0dpt6oV8rC23ze
oVnUZU7fg61atBbUl5WHPqA44B9akE6dPm2DmxYhrDOWJOYl5ZQk17lMuLaLvU8C
IQGDpWhYXIhanUNXW1iC/RxHuh2/7wa7JQr+wJ0ms1Bfttsi0mQb0FY12GWAbRVw
sfyGryI0+C89ABEObKBsJ6Ljs7NwRylOjggpWraZ/Ndnf1oXs9RBGe5P4MmZfbib
bfuIh6lRL5kfSBjGAMN5SyPHdzS0pw0hI7ZLT0q4be0GXuLPcW/+Whgd3/9+g06y
fqB+Z4RF3udUcY9nsGS6vWjJHh5GgSuJ3tq3N5bMiE0lHGwmP/gsv95ASFokE4KY
s45y4gf8WqQr/bIYHUtzp2Q40kNgk78CEEZpbX+uJ/mWnLu+dGYqY73weYJrrU8R
WXvuzi/dVTmGnuSzgfXMc+DoD7bHBtgWy1gV1mlvBH/Nf8GqmFoSbI1rcyN1ODQQ
PgD7gD3aGG1i0hCmp+e1YyfLv3dAtW2Odkhl9w80saTvu0kKYBLdiiDd3Mg8ugg2
BPXVA6eo8EA7JWp80Bfu9Jh85NXk5MFIdWWDMUCNMizqNDxwtJa3sjqQTmK2BLRh
l244xRv+zUXf3s+wPRVSmHLFvAM6TXatxE9zKIMymWlcdNd7yORpaxSDMR0nEI1a
6RdFNQgNosmBGjMtMAZG+xvgYU2GdQBLmbvGr9ViSiRASKJ6yuOekyaPQ6Hyuf4C
8MWSy8cYPGz9JaR7zpbMOurDYR2glk4eMtZCRGzwck57vAYkOP6W/SDon3tnYwXO
qTw4M+eToVwRLj62o+gvwxOd7oVeaalkYWLVN1cttyOkDwYCtQszQlZZ9kvrizBO
BNG+VkotNjMhbKg7Mkk63NK6fKwyPWKB21Og5ACEGGM5JxcKS27XErc4DmKEFOjI
GhdtC12R97fpVBzosplWLNpqmnPYjL5YaiaIVoZk249kAkB2H1A5Pin3Z9hkGVUS
q95LiJU+G5nKhRi93bxLE5ML13OjRBv2vjhTFOES2URXli4C8+VhX0o6HYpgfIU3
pceq36UYG3ScgRImpEe+057wemhXk4YCkT89bFkfjckf1X7uGaVLYEyuReFQDTdi
oP+Z9n0R26B//IwEgsREvpuuTiMfV9VvUUTZ9v3BZ1szNxQiAaxq7Yq99dNPDRvo
3UiOOM9Eq2DcJrOIkrAMyGwJRmpZzabDQULHAOTi/gDIza24HSZvNxZokAUN0HGE
QtzKTIGwJdBwpK6wJO1LzqWIDqQRL9RrctIXiLyTkv8Z0DNp0xRiKdder6KGuq5p
YnEBIoD9iyEJ6HJAgvCwVJpBeGZ/wQ4+nRx5nldZdSTMyBb9GJIGfRwwwoGJXYxW
ufDc3FPPTGzdKIHE8b+1W8LHBVs4ef24iHWlnMyN1aAdHcW4f7jVqLMC0v0oDn8H
rSkKtZdGIPxx18yQ1T4lufUGIJpZar6is63FnLIB67SNhv0ehNWFlX2W50YOwOPT
ZyPI+Cu9W4jMmyzIpBwP8SwFuEYaB/zNvdWLt+i43Yi4a6KQ95ydukm92zeKwI4h
Ck2LFol0nWW/VGZ6Hi6ftfHUZAnfU25JVD+lXhM3a+pp9l6uGrkfSPmYxTGKWlzt
T10OZ6y2IE2tMcpJeEOafgDhBlLoAHOAItJLH5DmHAf7G3hQKFsKJJHHPtX3nX49
XSIVKaUt/wP4rai0YL/YGfj4iRjPhgi7sKiJsEDkWdzTcS+d1p9qN+g7rCrl7RR/
kOa/sSzhSRTcDWb5kmb9YcJFzIlg1RUv0GfeSPGiKn9phV/eQeEuKhP3FrSstmdF
C8f1VhTstcZ8bNFT+fcLDYD7H31F5lROS6WCWPzNJRtvQyJREFldFjXQ+nb/blC+
X1r7Xmsq8xGBLlH7YZDupgt+t0O/qJsemKOsFKV2KJepIwqJ8mLu81km7gn9Prfl
VsUOEE9NKRxPbnDcvqwsGpHTLnB6Q9U60A8MVp7BvooS3z3YF/ubS0VT4Ht2h0Lc
C0nkpkL/2RnB6J1d+XDcJGWncxsAySpBu7S1xPty9na0y2QjmGmUXS2KISV6EHIH
0m46M2QMGkvKg9FGefXI3qkPax99geMfuTxTJ96q2yN/AOKH5mlu1jFtOyerh/Mb
9eJdmfF6ORIRzYAS0PbQ3V3NgfddXn+Z40LyRnYlTJVMh90BuQjvhusG/7q0FICH
NPz7+6yKpio5U68mtpncsP9zYkf373xFj0AB04zw8x7TLAWq12r0agJ3goc43Va5
W7SPsMHKcK9rEg5ekEat/TZysfHyNZb+xWv1h1qVirHHH9XEb9VeLWQeiRr5ut2H
z0ZCqT4UjByD7lUflMVax3gY9knX/IghSdr5sQNA8OiRAg34QhFXFXaFVdM7/tWR
WCAolkgVf+2oisglVCo3zljh3H9MWh9Hu3uyoYsGhhDqGPJCzMqax/t9D2hgbcVM
e+Fm5ek0g1AwqdOzk2+PnYqRwLaI57erCpzvunI+YmsqZQIDHWL4NWydY99Z47Qa
jwrd6T2N5YL4f3dSxYu9hks95ESHy5LjiGHYhT1a8aKjBkcD+ykmXHJD2/f659oF
rUOlBs7pIX86SYLaZbi5A9sgSv/ivazZ5u36NfJ8Uy6z5wSGRV/n6u+IN7a4fWRY
O80vIMr9wIXKs5F3HjrFs+lx57jXdxM+7g4HwzwQ7ieTXLZ0CFfBYvCtPKgYpxUS
rxvRLvM849efy6kNCTkGEkkZtWwCDV/YoXAN+9b6EB1CF5BMXSbQT09koCV6BSCn
Z/lZUqTMsDBbr7nFnX6KXcYmgincbwoq1zvulIxS2JSGtzC8N6GRN6ozM8O3ozzt
l99cQ3CqPFS37FCCItM+4PWA4Z3GSJcFKfd+UCrgOPNOUD06BkMyUJwe82DtCiLt
2NDqw9tcGXJLFkxYnow1i0HoPwshXPjND/t820qmZYaSgpzT97nLd8wyV2WaBroZ
EjJYvvM6pK3+8lA1TYqMdiRv0eInTRTIpCOGxibkJWxZmBuR40Uoc+NTXB31J+bg
BxBvAjRBwm6iIhKF3VrfeMsYKedlQTEpThQQv0YKUPEM7RUQY1XveJpn7I5Gf5xE
mFosybdNe2VnVFVU6L3ooQFYeOFXm88fSjjyfn0GbDOE+8RCuNrwEJ8iEepztfA6
k3RQUn882lV2mvs+8CWy2YSHEebfeJWTSMC9JRidwmctH4Nx9+41YfC0NQxMEpm5
3cO+qcrR4wf57CBWb63U7FxwROU7RIhxNQ9pHCVkWnG09d0v4elWeGbds5+mGodS
eCZkPQRGsGsGac9NLAPaFqiaU+D84N6/sOAh21/6SwUBgFZTe33hw0K4qpSfgZkB
3Rs1bFBAxlIuUKNtF8kJegWGOZ9murDK/KBHqV/SHtv4djA5HTm9iN5jXf8JaKB7
Pzld2fo4U9omzEBOZeJLAY7Qii3+C7rWccyuwTqVIzb97lGWHVifisObb/MQGhT9
TGg3mbTz7DpTQfeUfA55ccSDxg2MP7uJX1TH4zDwPECNLN9nb7/tWZg5uT72nGhL
I9zy3k0sfI+Nh1kgQIiPju0fr7nV6pbv+QL79uInz4BNgnhKHJujYnH3zh2PTPFI
3btdyPGKM+XloHOZEb0EFWX8da0DinVdTsQUDofTq+H53IsoUg7Sp4ZGpdWyHXpk
JdHm6e2nGbK7oHhOLmUrCVSvHSSIB86c79hT7T5qUEGZoiSbGnAX5JdTp2hH1Vwy
VVJElJyuC7YaS1MKc+iGCqq3/lHzftQgVFmwIhEkMTu8t4I3o8eZ32tM6Z7MZqij
dX4vkbKTr+ZGPWllbfbryup2xtCkWdHVEN6RyGVKIXdJFGVtqkW4Co4hEeX367iQ
aC7+qndpRegrqUYuTcPLRqop54IvrY15yt9VVktjUghMzbWCsZY3Gv+SkXMVJhgm
O6mhfKCA/cFlwnVJB6zXMQSs5RGRs26GIRwLolwWYgDPD1hAxmbH++Bd+BP/8IHi
eC37f6vfjVU+vAJPObJmUMDvP+RWy3sjiu4gtvVjazemac7NXRP3ldBxpmdPE38W
kEHh51JaM90TgoRapUsPabdP29o/M6ryrjwmjQ0bLp5mnCT5ic2w45E8cTRQcVmz
Q5efrrNPtswrMD4zjh1FIZA3WBuXu8332EVxyZ0fG2UWwvYh2o/N9+cHt+LzA1M1
JqVfIbXnsOVAHkqDXEY50QIjNq00M+LqcyipHqvvRf/Twd/PiEWYW2e993BCymDu
hAHJows7Z/3OL7tcB6a+doUQLVXTflxkQh6/tw2aeoYIL1XkL4E1hZAclkj+1FxY
t0L+cjwwihc9yGnEAxETAMC39wED365fJjTHaUGc1IgF71Pz4oCLuMjZ2lg+7GlG
UqSeDnMFk8b0XxyEJPiNLMLKZSQb5a95MSJteNvhVtYbdlXav9okJELojyU9YaBM
nrcTENR2DczXTQldfxbmBF18UTs3RRmwR3gZakrLTBE8EI7FI67k08w8u3kpJ7K6
WaVyNapzQHAHTasuLblmyHU1SMX3w7gRKXGIfIredSytujwiVQLxEscVDDzaj3bN
Kz5jzP4PubLWf2VoDnDfscnfm+losxJLRdfCc6fG9oQBjTm6LLKnm78qD1EavWAK
CAtHtWsajCTHljD94ebBAO6nEPMEOfTZA+CMTaD93bdr3vs5Nuvep5OAT/7UoQfr
E4rAd+H9cooHEyV4xKu92l9T44NC89spaP0aXiiTNiYKESMdVX1Rw5O/j8QVR4VT
0BUbq+EyxvTMeTJQ7lhi0UwFQVg1OgKrq1tbqK+XD93sFlMl9LB08BNdoMv8WGM4
QiEa6StK9AfdSk+tBF86WO84lmgxLAyPAlDWKg3ryrUBfU6QnpBrHwGKFOg1AL3G
ijrlwsM79hWVVEUD8P7lBDT2l6oMJWDlMu9j9VG1mKiGXImoaJ0eykjmOOCy7cg1
av9AMdx3Aow5DerEXFZH1lqYdcGZ69o7DNCSKPu85rFODFAWQv/jQsITxCCr9f+2
CJ4Bfz6ZrArRWa6TkNLALehUOVDfNtuQZ+zPFwcXneAYA91hq0NTJEgw6sTMAWae
yJkr1k3nErxdl00xMCU52vZHPFRe05gSh9as6GlJTYMLGkedyjG1IH8nhK++2wSd
X6DS8yfGCutt6w0gQgYkcX976yrggqHNXLmitHGfH30AZEboTkaQWaS/ddI1UCWg
FHw5YhHOuGCnmASjQfiolbe5zXxveiwZJaQ4o10XcQOxMFn7B0P0OAh5hegUwKIl
4w54O1Mx57qGgS9cYAE8KWIaiSvOxNsljComszPWR6vPGJUj/VvkoFk3Ei3Mx/nD
WE52UugEQElcvBtgiBPp2bilHgOzGzrRv8ib1uxfoRwx3ehN+4h4BxzwDzebG+xk
116V4726c//ne5pa1sWCTqSYm9Kzp86EtB/5s84TqMmjG50CTIqoX6LNur4vFfZa
jDDFZeCO1g0NfBDEOsq5WGJgnq2RFswIQeugCS5Sns+JxKxCipyFeEV2VZXf0seA
DFqrf9DvB3n+hrATKnl313iVWSGDm/lC020iwHXqqaOkZNOsVvu6pFVip8e6z35Z
QYQVtBvYyYeP6BkOKYJXVi72BTTd2+Zh/9QuZvwVrNyq2tDqLTerTxGNSz0wjhxx
SV2OChYxTSI/PPnOfWFCGPsGc2twht+G6jSmRYiUJF+NFjlYUtPpXtQeWwCNHVIG
xwJ+5FwgvnGRMCV92LpKrmaKGhyY5QVYJAPqhOAASHtNkgXfaA8tPeN3ZGC1HNTQ
NXjBCsltluhHosBofNztsPdtL92cvcgWYy/Igdz8ffIxK1ilh1U+W1m4IXp1Vjgq
RP4C3KKTNYMcWkuy1dN7J3jE0nDbm7zZUPSZj6abMEzUpIRP9yCsVn9pDtOChsho
qKZA/tpJyH1sYUmxy9enEFpyOzYdJXjlQwIqanpJ6HhEcuEGGkqRDMiSVm+ZDEat
tNJYSCJwbfrn1Nf3f1eGqvkQ0TEGY6RYhC64x5eTxvCKrK5Me5kcOdpgEfmC0+kU
OWtnWI1ojaCbZnz3PVjFaQBd0azuXHsf9WsKsV0Pn1UW0hCKgtkm+ufpyd57coXF
`pragma protect end_protected
