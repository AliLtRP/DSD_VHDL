// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Uon5KMZKlRlmvr6FTVvy+tUKz0J2FvLyplaFm7tibyCKLRAx/Dm4mZpC5B4ips17
8895ws4PJ8aKCGWBnG8SsveOPi0p/NJeEnRGemJ4Hv2p4cgo5RsNfnXLsPsnW5M+
nnUxbBiQT76imkdka9IGDSkPopV7unsFdJMpmgxZ3us=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 59472)
j6xtOQc8dZ4lJnCV4b2i/DjukYXdKC6gPyN4I9b4v9S6W+G+Bt8aJ8NzUa2d6IIY
FsWPnPzPzIweve51dvfNbbIchCFk3AUEKvB5lNFc9+Q1SUm/jhIZiAYKunDaUC6t
vRnINruL3fs9vIjU4Nr7hZsGev0XbUyvTIjsvXVolAF53JeQIKAGiSOG2SCW6K0x
l7GvsixTQ2sgX7AS+qCQqOxL6y8JsdCZbcgK1QZOx9s4C7T3Z3Vk9KSkLBDLsb/o
3TahmL0KlW4G8tIwv3QGphKubjtV1JkIh8+0CTDAPAz8uMR1xnYOsEl5HpS9neDV
R/rBPBlQpwI1lQcRqZNAExiE6pugJizYw2qvd1cKM4S1YJ7vJGaMJjtgq8GeDDzj
jlBPOXoT8FipW1iqQHxYcjYsXbwXhf4Xl/Sbk3rrKU4RiesZwkHaS4RVjJdFd8nL
0nugy5BuZgPTxsFaceVQCZNllay4p8PKnoR9ZtsWksx+YkYgcPOMN/VgfA1ZWu06
7NPa/PEQK2PIW5PT6C6RKItCm2ApyUAvlYrIxv7Tx89DeTgqTulofZbTC10q0mxv
ge5E4LTudJuqP1b1LLz07jBpojc6iHhlOiXfcJ3uw/8kb0xBfDh/cQ9yTsDi53FZ
qT6vncwLOxS7nxJ+QGNRcipFfzEu76MDFZRqvS7ca0tcWvzeM4N5sqZQQdJ0h12e
kp19o6D9/7D5lhZqTga6qPjC3D8M0g0rtiuCOK7mwaP2OHM2h2jf1WcIMmE7Q/nZ
FoHx1lbYIM9m1Bgqzme6vOXJrJjIR1pHF0DYhh/UkDoIF+S1UZb4KJ6hVeqxXYGx
Q3BFb653LfbGcN5FZOKYWFZYrZvfTWxGrXHQ/siYRmmA5+2Y3MIj58uD6NHF9Jl1
7BjLNMHJk4H5p3CdfZTVDtALV/BiVwrN6Po54FxKC0j38hxFMHlKX5Dis0Y1NrGy
ppeLusRM2zGWIoowN3Xar2WrXmX3FV7cvxZIKyBtWBkjzjMymyHssSftfRAduvR3
W/YLmUH7o+H0A5SL307/8tqYJ3q/bf3TU9ERxcG10/oiF9F9ZncbZF0zDMP3/6xu
d8eFpvomqp+4Gs5oysnN3f/hiBSeQnaDDW/Z8Lga9UhqmHlWDPdMGYXf3+DrGlEz
Bo5KDdbEVWm2HAELyXUwe48P82CW22glrii9s5+FFeh8a4MKYX059NGyBa9stg5f
b0ZAA1AnyQznYdgW6j6JsNBhnaV1wtgODCtmaCobxLh4DbpDtb2Ls0WxQC12wtYk
GEfJpPdB8SMz8Ictl+sdOUk2JsBaQKP6RFmVvHNL9mzyaTnJsHgT6vRYYoajynTB
NJaHrD/To0hVG5x1HPumbu98LWT825Qa+CRv74JfNXfiXRgR5kSy+DLPu4BwcRcI
2NTboqy8ypsdjDtMzKsrBa2YyFrArG9nvRimJRAG7EPvaM6vo4+KqXfZt/e8iy8J
3H0LZrXCQhupH5Qbv4BuXgLTDUfeO7VJj0tj7w28DIpqSbK8JjjyDoB099h3DYsB
UKsSUzhdL1L9CPlFgFCOuZbx1JUlGO87eMCyWj97yksd5butDp+SAm+kqQjuEiJm
IbEgI+f3x5HLO85SARUSN78zeANC2davdXVvABFQULgLvsrwGyh1HU/K9hT3uir/
JfaqSyKYcmjCg6VTpfzj8VTBCHoIOnN66AEmLVuaqun2Bz4/39km4Fn8c1Az/9YZ
69RkVFyPCQJJoZzKD/MTHCWSfU/6mMxE78yNOPnwgvbNAx2eNn6Pwzb0v1K/NVfB
fI4ZzAM2ZeVKJVuT/UvyhaR4ynHpRjCB2aXP10utqjdcVxbe947Zr34P4dqJz+7a
sS21uFjgU1QPstGDgvYS44Xgm0ndNAnMeXIL2FVDqvG58h6eKUvXbIn9OM1qSbEG
R4MESElXPwc7Atq1FM5BcY1ZCYTmDXJ66Z8C/MoxvVSnpuZW75Vb7h09082AAgzG
E+tnx/pAp/cdQHj7uHUWH7l7NSU0jYrW7JLt/F3yrNtsfzQ501fO8Q9gxJdT3cOS
0NThUm6ISlqiUjbcvLVddZdke3fA1yYNWJQoDW55MMVEWH7LfhGm/pxNDY/VN/iT
2qpGPZ6s+m5hEnDngUWcfMETM24nckNlhEDWbkaeuEKHu0MG97YOmST08Pjjek3L
Hl+BjFq2u+vrCw9q3K8H5mw35ZODb54t/tkWMrG7m/lrzd/RZGLAOMk9xaLEUfkV
O1fs8X6KkKdkjpAWY89QvaBxu90lxvXepiglui8RDDKMx4hrgMk/0g/41wegJ9rB
YsxWQmcLw3ut2DgDuyCWv7aPpvajyyTNmcio0/qbA0SMLo2tavuKDQlYfRt3j1HE
E8IoJr2eGuvsnhqaAQnj33YM5SYC4/ohYtyoHVN+VJ0mdhblh4h0Xxy/tj79RdaU
4WPJQXuxUBXU89OzxIqPUlge4Pu7QsTMRnpqrT4RCwLYWbr7DM6wBdE2s9NN/zWO
VBDIe1KlgzJlQaYN3gxIncvYGKQ/P4NLc26qhRIwRyWlt0grPWG55wW4z76OhFT3
+4a7YlZ/M3IV7PmRSu8yQV2zXBnY0LW2jtXYH9x5osGz2NJD6zFPUDGM5iC4C1Or
HySmAfKqa8nmm0TYuV/Pjt97sbHxm9wY7VSqgHnboSNwIRGynq8PVOjG7Au913IW
KI+dfIeaAM+EDz6MiSrTF0kgFPt74E5lcOP6hwkK4zgMvIMa9l3nwRGyAycx13xn
mc6dNEQ9Qkf/5G6inY1rIgnVZ9b2TZ+9ppIyAg7NeEDvRAn/XRWULD1oYla8fRg6
w9N+3fB2wq0JM60VhlK5/wdatcPrB9pDPx71AoTez49bDnjt7vPRqUgPll2JJfGp
jGHBP0OyVBr16jJLdMNZdFgiz5fTYgcXogpp1IYG70XobJtbB7QdzNGXNwAux1XE
VgWRykC00jxr6M4xXHT/rt9lCxf0bRRFLYbHOUlAtmKImPsgBlFGxL6+UDCyEo+a
PD8KFNJapCiPdg5Plt2hyo6AswiIDXAWC+a5ko6iTxjgCAdg6mfsSvW4VH7YTrui
OKtLXKTIM7o0tGfaRELX07I2m59MxW1/g48js+jT+wr2fC7fETLp+e2fd73d5blm
raCybv34yb7MeaDbPuK3OlFB5nh7Y+dQtievsZg5M6aJG1rl01KULn3hs6QZ1YQC
xW0dtsCn5636xrdOIdBK5SfyjHk7Cri8opPmhv3MNUaBZtdEe0SV3xZfy/FLK7Cc
B52D1F6jGEOVi4tWxi+PljPeTZJ8bIQk9WCoXSyVgydYi0jNnuavPcngsne1puZq
LJruhJnbEkqcS4St/8AnnhlJ+bkHI3cMItW3gBp6P91B5mCLQi0d/IFxeXIh6Z2c
Cyal4BQvBNFXmRGwja6Eat9B1sycQS+a/6gU1G0qkfAEr6Rab7nTgh3bIeytkhYf
Tk4feoHpgeLcPR4yHJdaYwcymqfajInZdlujAMnTVmzgEEaQ3jF7TpuTvP5DE4TU
ZwcElKXde7FXw5k1J91Km1+8wD/9/cyTbup/6bNqLsflC8rUDaFLPpEiIDqZ7UHh
jHLVURs3McUHRA0Q+FVQLJ9WbxccDc2raLtSi2Pe1dvVYJC8EsZBiTOOE7OQJ8yT
C7k3pFde7q4nSinReEIP+EPVKqgv3iQa/Nh/TGjZhFjfr8JGcgmuc0oXq1Fln5Lu
850SV25FrI0NLYg4hn0wj2rclXz8D+6VmV4ZH71Ib2fek58/6nFyj/6BoqaFJSxG
sLwVM2CQFTpQ/8PQ0FsgM4CXGR9MbhRNGrcM36YbJcTrTNTciCqx2ijgBkeLKlk/
BoqcCoUBxKROStngmwtnk2rgRit3u9SF98zVzDbfwBvxq7VjTVkM0nK92o3CBQo0
Cpz8SWcaIk+y8NTJLcs+U1HsIsqatN+iL4d+Aia7U8J9AwzGVRwLBTQF4HYcwW1y
plTQLdUBD2Z+4rjcc8ib1SzTKoeRq1DGUf1P4Wm24KjAbNrCZ4swQNefRgmdzq4I
J13zjjC6Ip5wn3yCidb0LlKKY6OPL6gin8jr95RZoKbqUdhoiA2GCWbIfMNctJbF
sWbD1koP2Ra30K9QtpvftD8/HNMGL341SjXy8qYqkB4S9Ois+RGKiWwK9ubM6w6M
Dv74fJPF2yDtyX/ZARJqMeuUbZ+mCFLyK4IhcW9PkTmS5F0ufvfPbysl/DUeNAkw
WC49ew/Qiw94c5WgqPQvSfiYj48o8o8X4ObbZxin/4NhmlEOoWVpIW5ccpfAR5h+
rdjnFv/yHHvadqFm9IWftOrmDG6Zlzja+/EU4WbxxMPVV/NtOmHTIP+QRMTyrlsS
icS09eACq89EizjY9uMbsg+iOhCNrrb/vu5+3TNlYVvco3MIp2zTEuT6HiOsRtXq
OGbYVu9KQ8kX+kxIk0/WQN6/UNuCO02TNj45bq6A9ejD70VElffyelK5HtzgPFbr
rtKu3dgIZSeOQ9teSx6dxeVxiBBXQV8Ufqtue2ZMBlO3CzB4CdyIKI8Vw3gXWOt7
zev1oMeWMXDwWWsn96fuiKFu2Tha/Gr3XwWy0+FZ8+Tp9KdCqDrpG0tqZKxLwJVG
RBxoZxNp0EszJXhiJD6xCjUIbYGDvPO3cBXIeK5xPprJKpOsbsuhV4cFsVRN8ZH6
w5BUacwthz6A8BICcvMuNlp/h6wiwBG4kol+8nIWhGjr/05wUIay0rheCbSeobrL
WpYtVOcbR45SGbIJm7HKmrVJmSLQ5IxzY+VFNxF8zsigAm69GXd/4mQizZxzEsdN
c4/lPvBiDnLzlV2ZrAG1PgVIFwN7hiXGpvFNsuolMcEbTzi7R+/WRw6+e5X9NsVO
kJSsC0DN/3TAm7wJTrmTFbdUAmbEEotwBKyQN1pchXsHEtoY/xdTKDLtMwVMZSd9
Z/P0+PUIqsKGcbHLb6enmdX5V8TzuzKXaQXU6rr/KXIzCAfJAAS0/c2yUnSOmln4
KTub+ioFvZOtdRsUg2FlqlPXbquzRwawQ5lRgTFmyLLC1aRM95A34+k20eNjC8gy
Eb7Yhs2eWs9uHbqTbhdP/XzBGdTm06lAVoZgbfZJ0jdR5PncSvAMaUaWJ71C/TXK
akRtMzlfQbF1yQXOUggjDJsoXBCHMPsWKGpTw6Pkjj5Erd+JxG+C69sShKWrRq4K
uscC4hNi4y9GrEihZj2Dm8nNCikAQGVEWjuj3NW41qHOGZKiPmatfHxzildoBlaA
+LlhxAPLibb1lzHnqriwdhKm/tHY33/fiji0Bsf4pyhZCCCJRBp0yOPZRdZ2hG1I
866wyIf6QLctN41tvYPISIFpt1w8PmD2MkWgYqBRfpY+VwHuflhhppzH6fWWCoZ0
bj3RkQlNPDfSxcCTqqo3n0ai8oDq1X9rvgYMlT9R9YiHAMhFP8yYG6KBRcWc4xPe
JAdLbe7aPyBlRDKDdA1cds6Iwr4+pSu7aohvLiX8AWvU4CNVX9pb/DksAScDpbuz
SCwzEMX01Ijn0oAGOxfX8x9tofa1xR1YJ5UyVBUytXMOVfuMbJic0SGpUNaV2lRj
0WSyCPv7l1O1A19AA3IWEOp6e4/dYNjfP3tOFBiRVJjWpICv2DJrum+NRPh0fZ9f
V91Q7E8oEgNOkAKh2MwcVnSt5rdedLc03mv3mg4X40zeieFhubd7EgEBUuJ9oZiO
Bk/IjC/D6aY3gmZrQq6DPTeAVpSGiICpHbbLovB/9sy3IrFM1Tix6flFDlyxfaMW
WovZHsQyvU1eRgAAGEQN5H/kqRuq7KFUWUxj0ShD2dh+7oWlL34K/FRliRH3jCMz
/y2RRM6SIFkk0PdTAEelAqyzSzSeDSQAouweZrs9OBTKk1wYY2VAobSKR30Zg3d0
WYAg27VAniRINGQE7RTsnCtfy62gzsFrymZ422Y3cZbd7NUKy5i2NOGIz7byA/jB
SloepQfgHg3U5onHazREJLxBnSiCKjEe+Ip7WT7+4gxUkEwVEsOaD9o1yvx4qCkt
CpeMFrG53tm4JZzp3HmyZYc+LOWSuUV3p6SZ5KPK7Olb86rERG91iwAjGmv2Zfd2
jmSfz4epCXVRcrtOnJ82BPC8LfQiA6WvDnYUYoU3EV67SelS0Mku8UrongxvhvlT
dKLaervFT0A9yKpMfSVm2XHLBxwa1cZ2ZY85vflUP8PIUoo2hDuQA6s7kngzwxGT
s10u9LIHatoXFWCmgQKqfpBTftH2K6IyGR9CK2+yyBlMSG1UbA85zhLBj1KwKElI
rNmieqg7qRIIzY19wJ7x8pMvuu39Nb9vHOb1UWtV72vbLjqGgjKcWMs0W9+zgnJM
fqSp1hevPLd7qXCbwG/cOHvNz4VuGM4m4rorz0qzc7HS+u95h9scQIG4DyHroyeL
Opk2LPsAWBXdjByaizKvFrcJXPl1509N3y4kCBVwa2fL31rKTuEabA4Q/h7Lico2
o2i7I2YqayHs7fIhcuynGF+8ZxbWLK9SY6Unn/S8EuqOmFAP2npjeEAwDMtQ4l+q
Mu4K9kRz03tyZ/utcHGmH4ZpgmsEsUDgLoW4q2JsUW94zUznf+4lLRHciPOnXMeZ
sy3bVUKwuATex+IwWK8yTkRJ567jo52ITPYIdzmF/C4rrgZTFosK2h+2O6lguacQ
uIVFjF5ZmZp3tfBGYR09u5cHYFn5Lnq6p1rytJyFWOLiWltKd495tkmZyKMUmPmr
dr0udClmrAthaLtGgsNHc+U2gCY7YO0hsMqZY7iEFu5xQuYKxBIal9VmodQvPuDN
vEau7yfSW8Uz0f6o7fpVJ/s9mAr8sDfs0U3XAygv8chGGbpBwrsxrzH/CtcfapqZ
cT6zy3ORm/b+ZM3pT+HMX1ZNq3LrJC9KckVu3Jp+tsfxD0m1fr5mXeCOb/SIPYxQ
9k5ScbgGNO15d1UJ9zrbOrVUiEbQiumc5hJNWK85ZwGOc+NMF7iVobfGfUOuQ2sI
B2wUEt7opBGYrQ5fK1PitMGY1689vbUfJmr/JXHnF8Q7dtmwRMEuOmp6daGm+Y0V
/99U6V1qw0qcpd04Ae58IIoPrkzgYHndd8MO9yx/N3d5HGZuJNW+WQuGcb2cR6xY
oNtxYoW8QWIBSzx0/jozfcs0LzhVmAHQadGDsFcxCjNQ+apTeIYUI30uYwukXZ9I
SlGH3WEZjYXvIwf1Je06xhoMLWkUUhKqHp3BccrIPwY/0PyFAvQvch1CY6lqp1Hw
CBjYXQqSFfHH1m2PJd7IlvqBBVzOhMu2TtnKRzaA5eBBWeUi3oiBELTa59v+TIJ9
qHsufHHVzJM9aR2USXnyZ/A2GjKNgVhdivXKGOKm6a9vR39bZ9i9UTiEwrxdjhjB
MVV5U9yl+PbHG4sZPxDO6FOQrvsa8Ca2+1wNikh+NH6y6H9xd0rNu/wiPEoXO5Xp
9vv0PYE8e9r6rDrf1wpPfKS2GoUGaug2UASlGt0MXG11LiG7BEq766ROJgJeVAc5
q4jskS4QyYBtnUl6UoOwolP7j4M9d3X859XKD2GDapifcEx9JZkrQeYOTLnG52Io
oCLiV+cB//+jSBtN47+uj9kcfJQ49dorC8e0tUxsuKtg55U6nfoS6YVcVbG48GKD
eVddvmCnV+hILB9M5FjJpAPMKC1BKctowW9BrCWJs6GXWwnyoxJeIU5MLRbCn0p6
rG0iNWDIYjqSult66WE8Ns4G1x1ubuF/gxIpzLi6LOQCfYquyw3yVlrymolZDd8r
C9/sO77g9Y09gf+W+Aphj/WEzKj/Bow89ghgru7znI8MAZ0qkAT3tKjUz7pGmm8g
PQVvoZaIeTxhuawOhiD7hX6pYYEnbutbCa2Y4xntTHzHm8/al4nR70AR+IThLzkZ
m3ZdROR+VB437N8BV34FLqliq2nDV2/0ACqa4mdYFx41c1XX6/1YhtzuiU48PdRL
2xBYB8kcLWyqmv20Qdd4VKf0K33goIcBx+UQEK6UEFLvvGJ3KQHj5R82bbIXsk2w
Vl7PFoEmElpsfMI2/dq5QByyTBJBTxXgWGOqKmZieQAIilqVaglrVhX6srpb0BKd
shoI0z07OFTcOJsBd+HzuNh5lTvvLM0mNIlwl3HLj6I9negqB069Wij1+XP0YVWk
DDk093F+6hOZr0etVIWLI7r1q5PF1MXc7ICKGZ+91xzJmvqv0ZwqByH4FrcMZJJN
MJC5k/4TGofivqC/AemVRevgqVEJed6Jnq9iNQ8YOxNYP0CJTq0Wl74aFA7nyXYv
Ua91EDQ1y/L4/Z31gPcNU4wUvOxx/u+zSiAe9BaFbJ/kAnUNn/BPSAl9xz1g7Yb3
pouCA7IcIwjVlnw7aRhWvkB3ynIMeZ7EZm5dEIrDux9fbe9vEfnOieSBORGrppCU
KOIZ4lpuOEL3fcdsBlRQ4ajb6isInqYjIXGRwApsp8sbSVyUnEYLDqmO271lw9KL
31JxVg6hoj/PI2AiArAwjjc5mVK5DhOTDpTplQj9kgNlKJoCBZMF66ghF63slum8
taDZWKsdtpNzbJYOv3uzMEZq6v/H2zu1+9Ytc3gg1amVJYeeEcg3LPkAgiPHnDc0
Tc84uc0OSCGdF6uq/TCsorcx0NyNkLdGJ22Vx0CmBT+eyze1MrEijsAbbdNYHQET
eaPltLXSHwZMYE4GxA5oJ8ExSo1Hndrm11HAVMRUa6ifgWyCpzlKLS+HzAui0QdR
csP5WZQ5AbmlEjmxdBLEJdx9GbC8Uvt9zjjWCkDb79rbBVughtKRnVxIjMvy6wt7
g4uRSLssgWdAjH0dCpVy2m8T+VjJlfYhR1F9iipeZ9RboTeDcTXPgzUi+rxBmg8u
vNyd/vwOpXGpXH6M04Kf3AEkSBz2xU7CK5mvyfxAHC9tXHaSM5kpWA+e6+6xPQKf
m9dcRTp06T1bEugXEcqhdj9ucH0OtNHueJW9IN6//teZDozbfhIHOtyFDJy3/SaH
2ELmwo5v8x4kKJg75fCUdHDoLpT7gL//w9C49gHeXCx8HtrnCX9z6qfQba8zBsgL
x1/KIDnG23dFHMLEKv2BbA5PfEBJHqdm+ZrNMztQvsUDs9kYb34VCdrlcroWG5YC
/FjtSEP6smOiF8rkvoiGwPOBEphYMpQAg7a1YobPdVC7FdBJIHzWnccfUk6xGfKj
tMk8DDzvjrMWpEXae88Uzr1BSr6317MT54+lM5UEJIx9VtdMW13G0Etms5TrZtrY
roeUUyn0F8i6Z+DYd7GSI9jUahTprODuNXKMKMUecyCt1o8Jcx5J2ujMOKAeQNzD
fPJekX6vIWX0E1u+ZsKVOR/cBJ34sM6gheJCUlue3UEvnl5YDg+h4m2Iz7pQzykR
zrD+hMof3DFb/51TlZYyJ4t6xfPV945XfopZkz/KfwPziILtmI7/H4U1ZgpqeuNU
v6ynfk8ylfWvZqNB7xzqOdz9/pV43Qjo+YkftMpaZDmuOTgUSwR4tKCtdwvENSuS
CZr5e6uQrn0xgjHcHsFNFy7Tu5ohTEAEpqjub3oE8oCD3Kd9EhI6TqCYNvPthJO7
ALdqvWd6vplpIL472KIYmst0NuJ2qD2GS4QxkriPQeWH75+tzT9URFTkbD7oBcbD
UC8gGTT+9RZDx/63xjXF0z6igARurpGRwC1qiQnm477NhVpAaOE6RqivbwUa5kv3
rfSm8d8d3MK3s+HMOOG2d2db9todsl4YmwR195I0A5vtsOfeAd79CKmYDvE/Umbo
ZHgUeFnRreuKZkZokNEv0ODcW4j89xXCYBN9949OdclQmsCyrjHivo/sfvBqSUWd
CUGlXIYuqH34Vg4YEKJdtC1hURjyaGyzujdhlrQR/qnEJDfDklOYKjmVXTFNuC2U
4aivm5MkU4dJUb1hM/8Vnrw/OJUp1bdD0VNI7/58FAtsnv/B/s3QmDnXr4jHyUWt
nuNxjnJYbLX/9eZtmQSeWuc26Uk9O3AztLgXXNlJ2YeSI0N9+c3mrASmCjjfWMXC
S+EODKdzIXBJLkH6iD4yXw17EJ7mCTw8F8hR0eRoNHiuiP9yhpAoymdqE4kPeTM0
liAoZdmb/LruCRcjkcjR46ZgLI1/LZ41Gt1GYiIji3iCVpCNVjnWf84SrFCKIDiV
MXmmYkfyGv/8VRN2WB5ZKUQq/eWJ4XpZPgMADEleuk+qWJf2FXkOx6BlNqJkf9UZ
W9f+FOCK6yGUhh8cJVHdGrByzUoTrNjRJei80/2sfqJNWzZ6WwfzWLPbtQP0QKDR
5ikwftKw4N8kegcHBUZvfDPAvjOa9Z5nls6A0XzrN/pxR+WpmmXcdG/9zSi6svWZ
Mk2XIURv/iPShZQUmXIoxNaDAxBxL8yQuIHqIVKT10UNn8GmsHMuRCbc5jXBzYdg
eKlfsJJ4iVosHtzXsvYa8FUp4hoVOx9eW7UebTSXj/R9aZYpV+5+9UyzhvJfJqqu
Ai4PjYCohVcvecwOAdAhOlNHtEYh+alkIcbZJu3Tk6911gikpiVrlNPIvBeJFSCO
7XQfPblVb90mwACDZ+K/FzZOsqMVMQnHdoJfT8bEJ52MYt4sG5mQiXA00Ehf/OQO
ip3yr0QZFO9P3PwcvLCY6JlwTEsoD1fVzTw2hA3IQQabVYcDGSir9l4y6bX3R21X
dPcV8qqfHnJwxHJojOjfPDu3LJweT3SuJwffYU7kEpIUlzrY9YIe/gJiELHG8WT7
GFxf27KZEu4TfeMs29G4eFmCln1oPnclsZcNflZbjp8U/3maeVsE0gGTlmE/W3Yh
7U9MMm2SSuyWWwYD9ng6BCPdrCLVSqzBzyOzzNw1T22ImOGmkJe+MglOjpgTRG0F
4zpAONCdNFNgJ8UTqgJgJqGLy3t4th2h448JV6Epy80L/UMnSxdzT1U2eAlC3xOJ
ZDlus+Im/1jOO4CQIwOzL/tLyNyy/yXjNzYGfFbiKTc+u5yKQSAgeq3AfGJC4ufc
JYQVnLvOWK/QXpszoXAf8Ez6kCdNDyRazlYAwSFdoRHGB1jSrpS/G4uAHpSS12GL
fR5GnH1Ob94Ekyem+3QP8Z2821WKwNr+Pl5+Zq/g2637M26tNUVImeGFloJjq7cQ
BQTw6NJhCeWFZy7NEljvf9AKCKK7zrVjgcHuQaGp9JwpUOl0NgKhtUtbwFX8tfdJ
JPIDiI3kJb3pGKpEIp6bQqX4zIslYuUouoZmO+2wmgTPAveaTEkKQtqY7hjpMMDM
ujsodznMoX4h3BmHnUrL73Emq7gIaD0bla98vUHgVxnjpftzaZHjcfcUSrh2nMsW
Tm25hN7EkMJ7Rp3IR/rM938tLqTfjxCwNnpKy/dEhvUknUrj+7kE9OUUXmaafDSV
DzBPMTF4GkSrBN44mV0EErblNxGJlr84Kt/AjitVbIEs2FMklStIEatS97fExJwR
eH1uR3tuBNhKsQUa758GbUX8ZTzgO2mvWu50paZdf+BEE3hlYdizEr6s9FY/dHOy
tL1BmoJyfwgwaxLzt55aML/mr0adOftDi2YX2b1Yq2qbTPqvZ6Um6AHjLy44+FDc
gXm7CBbOiBaflwAFIPSyGlabEbXdDrIFqruOFQT7f4IFmVJEBOvBg2hlu48Eb8rJ
jk1gYZ6exbo1zll44m/gIwWO+JJckz+sb0XBdUCPwUvvolwQcxQUf9mczhNgKh+g
PHI/3a/wc/Uq2VHc5nxq05qEX963pZ7Ch5Gp1c4FKhnGl4fOXgHId1Sa4BD2RHum
gufl/mtZvPbLFsi5107AtATP7tOAqZYOmquf+dlx1LjW90x+gWhXlBe2ME80XUOP
M8kIpIllQKWi2sdqVFfceb7FLCnebLxGCto7dNaRGfqLSxN0Z2zaTsH2g5uE+fTs
bKEC3/CJivK8/BaGpJZv+vH+L45y2A+uZ8NVHR63ympqrBkaWTRqBrHqSh+CV9LV
Mm3XWKWAcslqVehfLpDKekOjT9tVvYmIXWW8C6+ZqG0Ny8vEMdz5vF0tD1z2q2z1
TsRTzAdUWdTXKo595oeBhVSDNShzkNAkJYqGfBQOYsbFKxdkDiZThEJvqkOFqxM8
RM4Wmn6pk3jUhKZp9W22Zdfv/DW2ji+e0hULs1fZHVmsuBnLpHhLaZpD8Tjj7PS1
gwE5zlP3pV53B78j2WF63IQbhixC7HOU2vGDy89+V/HYebqwiOeiaGbMebRDjsxr
wS7ywMJal6K6efXWZCEPngGaLXu4ljU2DWSquWT6aTqQushj//G77umjEubC2GHh
H4EmMS/diYzMPsFNetF4FI8ClEeMX/h0gmDa29YLBgGBmvvXpuuLZ6Dl+BCs96dG
kaHSs4AXfy3CouJPNw2xYkEZJPsqxmY6NkLARxEwweb5E5veytlxeOPr9m6QGRao
4WxsK+MLm+i/1i4rhHMAA9UnxAn4X4Yp7InsrxROzoLDMk8oQPvAjgV6mmuDJD8O
4jKNmiLaOsztFVJvYWND01SDE09yx7X6G3MtckP/30GH7u2ZaQWz2QBtb76XB8kB
7/lZxSuAHI9sr/YwaLd6/Yy8AAGyrIOnOPtsXaU7amryS7p1WaDj+O0+ajUrZKgS
g0UwOVUfdmabR4CQRuLN7TWRO9HYUUTe39OBqxwkgDEpTZPROdJ0nMeAuM/zLpUp
tCIPbNa6z/Cs5iVUMnfWGOiJiiuYlqIWbwzXF3nt0Xzf1UxqcBzTUl029hktlXoq
77j29maPt61vm3wJS7S/x99dwV0ps9q9eyNXksWk3Q1sh2qCcJRLAkXGRmHrHub0
bVR+Vm8a/xqlcVrwNnRBXJ7nuKlK2VcrjNnuBAtrCG70PE9bovIYuBm07xfGWoHh
H0PLnNXwjXevtiZq1BDIiN/mXf6uWnw1p4JJW4MYmFwCE0/auBygAQhESrxTWfLW
8zlOOpSLZj1hqcUvWh6MQpMQxNax637CDeEAgzHvPk3AIuwZuh95hnbMy71nm9lX
+SCrrgquoyyhhA228y4nfMf6nclZG0cW3lLfkNQl6jbT16SrmY154rwpuPQZ4xO6
4ZfW4xfkt0ieFwCUsBxrvNGhL9yfdzKmnl9R+x6kExwMO2LQvYFGzu5QJR0X5ioI
Q5KKgFByWu7vccFtXehTsrmBWekBrW8JuvmMiEsggSLt52/oSDujjJkqNSSDkkhT
F0aR40a77f6vS59309qSgLum0xBCz8z5blfN21ICKQ5XITi2THCbUMvSWrwJWKHq
OdKld/toIaRam+/2Rr8IFGks0mTt08tCjnOBmhvqqEiZybAtxCAGmfO18aA/zn3z
igBumoRWAQ/7ih3wi+YqfcjARSzlqs6y1cqiHRujXxIrnWYZrtupWZv5Ht0hKjn4
al0tOfw43ok7jqlK8Xib/reIj2vo2Bl3ICa1WrMw7AzDrvygvYgNq5oMfDX/tm4h
OQCXn3Ktqnh9QNsSIvXcbiK/Ab7XEAL99vwXbFVTVMoTsYbuXiAP7OJQrW42HIsP
5WVxXyjW/8ljt9Y99Bep911/hwutDBmGvIszfBHUvKbEcYyPdQLsYD8efuwOgfcY
c4T7zgPv4dzJqawyfUnKUAw+O7rlEdBkzsfmsjsn1FPRXs7qloFZdSaS7FNX7d1g
ue3fMzxKGL9r1a4gqn1oJpltgCzYEnTCToB8QRh6kRSMfAsdpW94+Km1+JbGpqtq
Pr7nS/L48eZGbAbcPoJ6QYAFTstNLAaS3Ou9UYikM5xQZUyXp5qblgFm9OSVpOmQ
xv2mDDMkL8vxOI7+fOZLP8BySEsM/q57RtnEz5t7CUxDyLiFVnrs0SFoWz4Qd+XK
6MwZq+kY5aHS/H3gMlmVJVtMWAOf2ZajaeJbL9G9j8rq9A0gwczPJGBk30vCZjjt
qWK+tWDFVmPj+Fj34DD3mQq/HjwIgKno3WjmrYnVKvF5RNliz95nlPUuc7xqUSgr
T3gy8jRFi3GQtVYQT7RLgxzLfV45chzf2HQxNnkgu4XH3+ExTxjU9rTsVYZTO09R
Zwus0gVD501uPu7Wh+xicjndymcW/I3Id/ZuXDbpMb6Zlbchl6WChXBtO0qrAaF7
vTEUu3zq3mzKpmrWzh5h+x2lj++G156NB/gdDTbtAFlUk025AwgDHQ8OzQTCUc3n
uiUYlR7yCQLOA7Yu/hHH269AQacYcL0YvfR7Bwkd/v+A9EizCIk/jzE5H99eUFfg
gKhCskIMEQrsffKxq5noMgQjwTf2enPy4ZFuhIuqaLH2kuT2FuT5g+CUPypo7k/K
jHxrWLDDNV07VB1XFx15gAsw4yO+/tqe2PEiqObb59Vh6aGuci0jqQJQdrELLeyL
cu+siWSE3AZMa7hl5MocA+Z91kTfeLFuAEp6LGFX3kCSPnvk9t4osxDimapURTA9
2C9AV7dc59SqWPT/vQlW5FfZPSVmFpwNYryVTN+fcrM1SQcSgZFdA606E9S8bXdG
yS3fZJ6r40XSXyxqtRK/BNuht/Bpgdxp/A9KLVO2mXdzuGB4XmSb7B95wOm3aYJd
L1IgTCbyPRpFfuhi9evxy29kHQ4mfo3PDHFjkePyFPWopnm2viBj2qB80megRqfN
MGQl5KgB6VGh2KRUun5GsxxXUKPpvdt4NCsNrsaaJRo90+Z0kGvxVtSKlspDeBsg
INMPyvzRG4V3yRvefQciZzs0xYfZHnz1rU+AeTPhFURNyq78Z1aFmGyOipOroi/D
84xUmTaGfqba1xTwTABS9dVcve/dJqG/m/YMI6K7sB6AAsrjxsnVqQ5UgUH0Nwny
nC2tm65Br/RmFnqtOPQODKFgyvzMJH9lhQtUpS/n1pCbKX4cWPubFfvx7/4E5Ltz
mul5m0b9VJ6tm3d6O1DnAKEB0QDI4z3mvxjgQczVpRdrq+FFM98v2hu6UamHjTUT
1C4d63wdObiPPEdlNNaJFgg5L5tDf6xQdxpEmU3jot+Thw/4Be5xmXkEIgzPJoQ/
Q1guoCGUTNneUJbPJF+WqtQ/sUkFGEUN7sHb0+HEFiQksq7pzQlNvjsSAdcrB66r
SaiPU85VuSAH8cO4DW9D6h17vS8PTjufJLW1R0HqM6uWKJ+EbtOb38ZoVcr31pDm
5kQQSoGpUu86EWlLJb5pD7FXpuRfHWVEAXMemk54jibP1KfdulNwWcGW+xpB54If
gGzTTFFF6m3UgCjJDtHvlWg4LwO6TFfhxluqzIA6cBGvMPorjkpPkSL5GVTMGS2R
VDfCL/1qs5WHbrXgwJQlEvyqRZcHEZwvqPIpIEJYEjpcU323lvbBDhDcLGngTdM1
rUlRQEIGhlnLD6Z6OAh2Ym4kG7ao/1T0FMzvFcoSGK7WBY+IpnSE2HumC5ABi9Sn
rEuNU3vQhPNPyeJdtgznUfs6e5ET3DXpTWPNpKPBvTZt2HPh99tL55xD5eXCJDYg
nvQRAqirTqOzZi5OmxkWbt8wphnpc14DtxjaCxjNvo489kRgvXGbcywziK97rmlZ
sbVqMFHRsMGLh0hFaDgRm1lCAFQgJv2YIbnVhSP8+JVbR4VHEepnAlJTsdyUUhFA
uJo4bBcc3kG8+yObDoKRm7Q3JsmByA9ZTygc0DNxz59QsML6Ud7NWCsJE7+MBBpn
nLIff5WjFOY0t4rq+qE1XsiscB75YwOFrkarsp84ZYKQ3cVyI5gfUyHT0Y5ebriE
d9ofRc1BxQKy898DNNqaSoE9NuHIVf+sHn6j2zYamdpqeK2dPA3LGgXQJyfhs39V
eqM+8360V4JWZmkxejtoZj7UQSDNMSnXzgaesrwNCZqpWumpeO1j6mTbWxUuWAqt
1CAfL77Yp2gFtrJRfYzKFQEKLP59CZgynjIsf49nIYK5JyxoT8BjvsltbD/ckDSC
Wj6r93Fdiu8wZZzKwXrrtc3Eg01MBKHLoffMXhxglDzze8gBpAvfuoOvYcqZFfNZ
gLnh7zIMxX8tcvAonqfU74eh22UB39J63jrzrFh9RNQxa5mUsZNbvDlTuAN5uX2C
lmhH1//Z3QTAoazE+UdbpIXEyt9uBfCrPymRD9wAAYShSpgXiY1bfsnWeDfgSRtW
ylZJMAfUtx+Q/W44b87m0sW10A6/tQ2sp6mCMHh+h6YZVF+oVI7pNxFB1eSJoWjS
jh2boIPXqN4SQu4eUEW7qH7zKxjV7PN06uP656rx89dtnqr5JzDi2dnSln0amjfA
DoB+Sp3ROdwc0veOkPjoq29+x1KTAVIK7S4GiG2Goh9//q5WlhDhbGy8+BtU8U3j
KWW/42h6lbjcdzJu1DPJnQzSJtH2qLCPguSpKcuqRcmRlc856JrsJDoDvmqlEF/W
ehzmDwXQP+EcQwcsLFhpIK97Koh5C9P+9nqtV0UJr5trK7TwVmJ9U8fQLMeAQ3UP
RItNZg4tiSeD4Vk4FIutFQuDuSpEoPmmgl1giDI6qm5plCm1LFVwsfQRPgR4s128
RKAdrbQ6x35gnDy9j0vAmcFiKTv5wDHwvOCk0oJukleB6fuuVEFcEYlRuT3ZbBfW
CUy1IUeHGk9jGIn/4TD5MsNzVN1X7ILxenEwMQ+mqOks3BQ343prr9FE7J+4slkG
lE101/opMgE0jjiA4O9P1fvSSfvobRVaJMe0sTv0A0EuCmzwbAyLUS8qpJLfNGxi
pvP8zZMTTTwTpKcatlad+7B0vzt2HI5WaEvvY3NJ9xKwTkK+F0v5AfEL8rng0Ree
bhue6eEwcvUa9GTTrQs/7DTInCuWH3JDAL0Y5SI4rSO7xa37zczNrvVgDSoV36YJ
gMgdpULOsfzVNoqXCPNih8Kd8u6Nf4Yxj8/I/jOelZ6WA787xU+SyIYG+jsIUyol
wn7AjeG9Wan8twiAGtxF8CkX01BVxN4vw66Xv0nsigXNNCGLtCqnKDd6g4Wv07Rn
Dl7kI76K779wy6iDzngwSsDVxmaFz7eOINEtdFicVGv+WcY+GT565SItHVWlXcdv
3eOroJ8UOV5ClriJubd86g9DIx+EAROPKbZk0avd5/lc3hYsq3scW9ng3q8CzZ1V
xIY6Nz7smboap6sL5M1nJOgRZJKyxAXd2oDH3rmJrd4GGGajKmz8+QXwdgtMjQmz
jQq4i42Cfr36uuJtQe+4lHzJ0CKn/6uLXvp9LHBnkQEnInn45GzTz/9IP28nzlCL
aMIH8JqjOVdFzIY4GuCw6SotpSgC2r4Vg1oroOtYdwYcBCIsGDDqp7qy2+pVoayG
eKb5l8ny+05FK/ZSTsulRgMz+25/W1MXBvJfG7M61SGpk3fbiXd0UEP0HmH4cLMm
wpzuatkBXyJ27epMIZgkaXimbXdbEaNQ2kn1JtvrWcJbbaGBVVI9Vwbaz3XBaclu
4YEDP1TgCNe2YOBvBFUaKo1V20HCrYGISCyqw/dQUz8gQ6qoiGYvHuZbfiD9UFXz
Ge9VKRwWHDJehuEmc4uWTyXj7dt0TRU70QMEfxGzeyvQEaQgSwsN0wKhTMEmg4e2
yWMDsMqgKqKgcQ8y2gj8TsrIJTXrvX22ALWVcUG4b5jYluJCggrn7MtUOX+BSS9T
XeVoaVmZUwco+j5RWZ/tbcFiQh/5M1qv86CbRvYDz2Csx74IloPhxKMrxJPMVNSZ
1Uz8QceDjjtEZIYXxD4STAd50o9o6op+sCCyizY8sj6lr7GlCPJCO9Al9V1ZhYGU
N56yGmBISjCKd4SY5T/oeiL309DX4NunMqJeQsGIKp8fHkD+fJywO+Yxl5Ga0har
7qmWeYTXRcWDmy3Sqw7eKf80+4PkQPgBeZHT6/joCGINwMOJwQJhwGBqRF7/AYcW
MFVMY27dvdm/ub0/qNvFy+TR8EqQp6HXOT8E7DGJdbcP1MJSE+HyNBdXNot1M+qS
3rdZWDZ3qiK+jmxYl/uaCC+LMs2x6gdrNqAT5dCdleUcs45h8ewkx+a/+J1G6FRg
3fW5hbjHnSsU03aNLqtaOuhCtsRSv0CRmBSi8+RAgsQxCc6pL/JkTWvm0FIlRb3w
5M2Zezefc63xodqAGlUeGyTVpYli+y49sRGnImz9Pohe5lipm1XTLNxrXwJpP6jc
A6CQdm7nEKj/lrypM8N3k9V60GiqK81CSDcgBQKhdBOkR2jLQJCOX9ZG3jjavoFn
CvBNmb/3Tjz1gb4vul/86ugmhdxfFYAsA3pRpTnatTAIoWjtVGSkKQK4m/ebcHSb
klyl4zcZJOnaKGPs1UzrQQhAqbO9929vY61EOI/7YHSykJZxPF8xzeJ1brbZVayh
qgw/hCvW3y25bug2Y8TdC4iDdr+hPLxR/OjhTbJX3a81+8okqN7jbecd2lBVxisf
aOdMLiEGXyD067ZeDg0IFhBNAtACpuv44SMXkqOZ0YZBHMEbDIe3PKW9tcZh7eZm
XX9JTWdQxTqQDvPenZ6mlr/RAVpmx1J1E5hPC145+PItHmnh0gn+j8IYTWRhqQbu
Dg+X8H/s3seVp6xv1/dIIifC0K9Ach8W0FE2oyZQYQccfRreaeDr0jR5brz8M4FE
ncBU7WqT+jULZTg558Y8ESxiV1cuCI+d1FEUD1Q7kV8ITBYfIxGPdbS4EvF2kV8+
tN7trNkhQLQ1AUTEnMJvsD+oZH9LG7b8+aibGvrrncrLJuAoya05ypPjcWwnC/1U
RHA7T5sus4p1By/4ALUalf9cSXze+tG+pbww60CWAWItHo54lf5uIBPLFQU8SAyI
lir8/JohXmaOTzgy02Wy2th7DZ0QczllzkMiF2kud4tCE6SYxJRhX9auw0k9c3wk
tfbJSarsfMIHEc63L41iO2STA5G7jp97AiWDyYa+4OVY67jQiSEBk3/f8sJhSJTq
sR9xnmvah43L3BLop9RsSmoKXYCPFUNQYXFUHuMXbSfJ0VEZaX9HQ8QJRCZq1NHR
mVHxpMHPt+yCRqKRJj2t1t2xHzDTWPxjfQh9yHiF0ECI284sHUFZDhAp1SvYxgYb
tghPrIABvAIpJA77EP/QjXPfpVog7kWhs9Y5ApW0J+/OnbeV2Gj0fzovffd6LT6c
xM7s6zrl4kF7qWfWxm9qk6RiGIZ8T7+zTHxsr0306vvVa7yw3fwbqXDvGv/abSAi
kiB4Ipd7y2oSKnStaJiYpA982AhHljj+dTiOp4UHiaVhuhvJ7EyFuwWvlfxhNuM3
NS9xYMu7nILxeZMheg7law90OWIEedUR2SU2ir3qujZP/yG32nZWvFQE7B1mHwuW
tIKGPF2Avecje4dDXxacJm4VqTD4pe3yTNCRylDNtscnnzOLWHhTL/X6SK6X2k6k
LI938UXyCU8w6EpkipNoXjxYN4VtMzQYeeuaAllddL97NQTHc7GMdBRtVPMVteMR
6jMHMnWKnu00ZnVRV3avIMcrYNBJS2fZsFm7h6eJFYZXxFizJBnAk6dGjXvSa+gg
F8JSgmGbGdy1BfnmKE5rnnhIwcfHxD2d5T0YfMgW9SJcLO35JXKsXP5DM+cz4kfH
DXhBKn2/av77NugEIUkhneEaBM//qKrmb5dS+RbqEe2FKknqzVuM1/5JDreyQ5nc
gXzsdKKSYalfYVNu7cbJpKLAXLa++49lDd+8j9208PnUspqR1QrFjweWkkmJfpEG
KBgMe0cmQaKLw/ScuNy63Rhd+EgtZJszFakqBfuS7tddOhe+LeW1YrUhmc0eEa+j
YgVWGwx9SZQItfhMC3NwyMAK1upqUztO4H1c4lwKEvMDXSuvruJqHNnELLXFAatR
pAKjwXlCODHqLdX+Gw8pHZHyLE+dAdtK49oWTALkbfO3/aKwWTgqAdKDI8TY/pE+
YTmTHcqPkVRqvLEr1WuypHjIQW/9AFks3pcgN226wLEHKgVU4A/eOjSVLYdxZBkI
0H+BvzNuIrJ4tPr258XqbtCVZCkTZdGyIn8nFQchPZwxpIclI5AqIHSDa1C/ZuiY
5DguiuNAcC0QAXIPCLO93cn826XlfzvtjVXN4hSScuDe1Mr45L1j4HOdtaYZfJif
ZgbJBSEq39HuePzsrE8ve3BquYdwcCcaAqN3GXPdeVL+5cJZPJsKfbM/JmJQHZ2W
gdFj8Zx6UYy45OBMOtGlyi2bbaNAmDwYZkc7fGLlI/VKuTGI+ATvAVexnxq6cck1
QhNkQQhbhXJXLq2a+kbuBXMN3kGiJM3ARw6izJTmTk2jriMg+n6ByZjQF6FS7FPR
wcmKqyiOImDzj2yvT4nvoFCHlXeSyWyWgMpY7P3uAHokBWWZ6j63VRLDK31feBHH
CiqI7wNUSz4xHogAx8280QIARWt+cqrx1q4PEpXScwRNoTslPZRR4xWBYM3ZgSTq
yhS9hqcNc7u82aAgZevyNZJ55n9urR8opCpV/rT+lVDn/Of3d+vmdf+oMieVWJG5
Ff78QIexWIj2K0cnWt/SoEiUv3CIUej2F3ePIZJtZPAz9C+UwzdNRTfthLc+SAEv
ULTiwo4NGqnNBV256bVQyHt41HuA2U5xs0KZZBoLdvrhWNpLywBeXDIiv7Pw64n+
azH7T9OY/9d2CK+8z9dXPEjzS3buPd3CNP7T/3SzGssdMql74s+gzH/SjjacqdBC
5QqP0dy8WgRbPiJ39CWTiTKWaT81h5plWKUOU9iL1vzE8+KxyjrPsticwHTTsEx/
kSfUYDYljm2UEl4/Xkfzyby+veKVRkKFbiYYEmaGbG+2BrRLHW0xHyVKOGLOxX2R
ToI4DuDtN6SRpddL1Vqm0wo1a+CImNwSiK2NwsS+8d2YRckUqxYJjZCxMK8yVWye
KsXh0v5hDUwnzbVaNOOcyu/4IyfU4qF+h2z491o2l5gEfL4XsLXaUraC3NE0hBIJ
aRcaosSA7yheJDW/flciiW402hpCRnIvDB8xgEU/+UwckFD73NN1WJB38AoGE+Ev
gVsqYRcl0N+z3Do15aT3GHRSs1HDtZlYNvwBkYBLrtqRQYwDg1SZFkfFsGPK4pN8
+/0OMILi+mU7KCorHFJ4bXqd+RC06sDQsg7CgAJExjknTXBXMtnIDWPw7gTkoxCN
5PRt03TH4KQfkpLxSvYno/QlXGFd78s02ntsDkb2gfcN5zCyg6rj9/CGWFn/Jl31
dG/ZGtaZYgOM+wCRffqAgx8X7bfPu58j7btarQ6qrqOeTL51dI95g5jEDSkZkpRR
8MK1jm3v98h1njdSPNNF2FpIVLkkFIeR8dgDaAVtuku5TIrF009f86+Y0VYuuc2M
77ElWFE2wmTzSCnNJREZKwHUtL87IXX7hRlqKAT6D0PHfMGSw9NreTu3vBGj23Se
tqKFZOlo9ZkW76SLvBTGOU6cFVmqgjAiWoF0VixSDzkyU/aNTrZ60OuGRsRvcvh/
gZIbWex54TdQnLdnEmFpDTOCWVEkmRXOCZX0OFC6vS8VrN7uqvJysgIisuMKeJmE
n4S9AM9I76c243R6dKlex5US8tRBI1nrOSzJ++mazwK5TLWtmh98gCQ/NNOp3+iH
IQeTn08bDztc91LgyTLty5w8zKWDBaBO/MiFhjWwYKlW6Mt7uitrrI/5F5HG+Q5C
LsgE+iSpF9Dy2hzM5ZwKur4T/4hV4Us/9wkBfYvBpFyGVSp9ENYJ2mG7GARSu/r2
O9jdx2KPv14OoCXIw7M6/cB0h1WmNHJQltBvDsHJUOco1Lh1RXUAWGQXdpk4aJc8
ikxpOx3ibqtmb1HWbCe6sQvRO4Rbzlql/yHDXc8MdRrtbERW02FH/KpVimuRY6aY
V7wyc18LGPAcaGYt7SDZF3BNr8+nSqSzR2qM5GCjy6CJOy5Oi1TUhfvI12/iudx8
zTWSIvxZtpIxhzXvWP98FOTBSK7zC3PavekKK+bJOVKEBIrGAUYUohXjPuf4rN8X
80Wny1Lto8c343kaw2sbGco9pJ3dOv+POkhhRZeei4SmHKcfORUfM+A80aufKrHS
jYESJPOjA+SiSd3m8cfv96z07VhIb8Vz/aZG9AJSqBRkW8+z9UEB2r6pWRUcv0lV
5sJ+bOLWrFj8XBtz6XBLQytvgDXasYpgtqHSJqSmZep9SituXnX1929bmpn7sLRL
3RNEjQubphc7jWGV8sdmamRpcxqNlSygkpcZ+PASIgF7sCQKwmFWZajpALoOiu6v
v5rVgvwWzduxhmHfySpNMVudHMumbx3/pEYuPow8t2ZdO1MPOCeg9rYRX4mEUpAg
KF6mm4z3afEJplwttesj3rZYxWA1aazbgPKOG8A5A//6PaqIg7A3GAXsQkAgDIAR
d98mi1efmaxwLw/erfJ0a5hsu30nX5IRsWlf07cf0pQCX3oqEOfF2+Ln3MJYOBr+
ie9vFeih2tIPfRw0aPPihb7zThKqOvchsHfTV89jFOEttBLEZbT2/T7HpqAZQbIB
oFmougGx2tc2KdvLk8iBDgIuS1J+/RI/k1ANe1T1naBFjR04mep3quMwwP3gq7Zl
ma81LpglT3++sfmtNaV3ozbOIsysBqzWBJVgCsbcCWV/ClMqvbPCYAQFQz+w/EG1
u7B+d34+chTJShdN3WV2yv2oHISlzwyvjz9WCDhs0RwUz3j91r+fZdboe5KU+flI
ucoxXQ9ERPHSoa0gZfX4C4by568Kxb3UAdhX4bGrot5EGTzrxF50GyW/9/E7RMgQ
jPx0rYQlbZEvTt6e/AyVkKZ/iZ0enyV8l7nGO7YpCArb6FthaW9V6dJZSkGRt/jG
9DHAJPKBU0Rhk1gqhFEw/1nJK9jo5EufqS7oUoyfnzHNJpOW77iUUqN26t8x8pYj
W8sZMbxC7pAgNsliq0s3u7b+iybSvCyV3WbArZRdgtGN5yEkIzXs5mOIySyGvYih
qta86ZiaHwnpJ6CI3FMIQKmomYpvwxB1nCsS1SfCThkr7ujiU5ckuujA4gY5Z9yx
n5QtOF3mi1dq0boZVE3ghsfuLUHdxnLIQWbHkEwHhMBTgM+baLucYE9bXZcf3Xxv
VAyC8kbUZx2/AdlEok8hmK3rt3mKG5xfLV1XqVZJwyTXNggFO1/+7pTQcb67uN/I
dGWq2S9VUmuCHynsA/JJDv5Zk4KNgarWhNjR/NA4nyM7pXXos5B3qAICweaKfOHX
Caa0uu2QnEwj9dPB4irpOW6wY0zNYr+7lJfwKontXbJmCCQe+FkAxKRoAxy1+jjJ
Ha/jnLPMdZyhPuoi+5dCoYVsPIvMbkGLuFUAZar/5awBOa/0K3HxGqajNHeXZMkK
DAeA7ICAvhhmefN5NYULQIseavlre3lv3pqKxOVGfz2FcYel/NNuIG1GNR1EZLKA
4vto6lfZiebZS1ftNLpKM8BpPbxBGlVi7EOFOG3mBbBGqq9d8syVppfF5on5XYDw
tGvaNIhhTvFkiAFzd7rFJV/llk0skIogoD7VGeV7HYT8WB9b2yZKVs+OapceVocA
NlyWDfiNKw4W7LqO8YRddoskLxTimrgQpF3s/a4wolU5RsAuzjkduRfa7Mw98cv5
7YxbmjxpPo2TwHfREYquih4AqV5k5W2o+FhzOYhemq1tzDHGjokQFPxq2Dcg1WZg
DxRVNBVR2anwB4lmvmYDceRwabWWiFZLwIroqedNAYtvs+vMId7PNXKsZW1aA4wE
OTvuu67wvSHxVBi7RM8N95CfENGJbdS3dRtVxGkZIPfCb2sqzXmcQmQfuxfZfvYU
etFhtMv6O+xCClkcZgVFBjI3EMj496bW8EosQ7EWHaqRFB1hjTbk3QZMlM0xZCXK
oiucB+4WVLeLW5sy5ywNA6hMn9hCQK6geDUKyXrQVBR/gAb2pOBq7tkcdm1GrQPH
tpHRI/SX/7C135a6Xb3Gk5OTqAUpVderzppjC74d92XTIxYo2Hb6RZGURVGmcfCK
p9MYfky1zB3nR29aEYavAJuBVCgTDpvZ3Pq1aW5mKmCRQsXDHl2zq5zqfPC0qdqO
pQKUgWfm85rmyfWn9KRmrjbOy7y15DGWDt3gmHm3B/dnCT1MqXqxW075EUxqUaZ7
Lxm34HXWuMQ1forSKkQFqWH4i+G4S2tS0Iudxg0EKaZcsizI/tT0yN8l1y98UKJU
QO5bGShtf/YeJQgcnPkdrlizlEpikQGYehh0iF7U+35T0YxlyzUpEXOhBOOjpyUV
mDgHASfIgVvQIDg0U2d1lznh447beRueCDuT4O1Y7MWsToD04RvE+8k6x5bd9ZXl
sq+BRldbQ1dL/NONZelQ4PPIM6/xYvV80DNuVSt4iQEtOH165NNperoFT4cJIoMi
N63ZCY0RTiW52TfMLaat0givls1mycenpPLhB2WG4B4YOLfSc8cVWvYnKUMt3zQB
i8qE4moCoxkvm/bjyRNf5MnK3lAgC6da4EOPnCweP4rk102iqVcCwkaEYFu9LiaS
OowGwLWeew+bvtwYUAAPBMEcUzMfGyc70UtFtyL2+icivZ6vh/sOxFq0g9ChPyER
BPjVwd87ND1fO8rpcwLXb9ydd7aG0i1C7WudAhTuJ5Ohnjk1bef9h5UgPbcR7PcX
HNvwGq6+kt/5Cgqhae2VMNNi0vzz4zFSxc4d6xhSaaLYdX9OyqseDONU8kcMZqWu
w3L7OFg7zwVYhqqqWGbY8+oeVudDovvTlyOdnVn8HVIjbBWJmRXrKiQN9p2rmm2B
LnZbZ6MswkO7GlqQxK74FS6ngGYft3wO4Sc/yNVCbQLKseqx4WWAAVI64sNMMh28
kj/4zHGfO5HPChA3V8i6GkdtKr6tofAz4McAhY7Bhox37eyGEQIZNx+sBFSvOP69
pCJc/4QHNWwhIU/6F5oBOueSybMZ3v5jJeZYZafQXf3zMRW2PSuoY6u8l2Lmru9f
nxROl11IQZpMCMWESbhz1xglUzzoiqXP1qLz+Bs/8ab7ORb6jJHWh+SVcZ/LGiHn
8xpZouk733yzUFAxWUas4cNrgigmGzXTn1EecwL0gWx53P7WhFKNSwm74zUXGoWb
CfroojAmp0FX2vAr63zMm+Twcs2ldFwDU/thFeqT/salA8+stJNGnzRg0N95UsRw
07VasQp1KO5VusstvXTmRfubrep+SASioliuBvDSP2jKTFeUnIdcZujelNpfI7yI
ij22PGOx0fSbY4YThl8j7PujGt7OyErJWtO5vQb4LBOO+dKPDjiImuWNYe0AAnv4
y7tr2kREvqaI2J2zz552ObfRYFKUSN8I7qMSoe2HTthpXJI8L8pyp/dW8zcfaVft
THJZ8XivV84cY4LcVIi4h1+5i1Ui8qAa9BYjYGtFTvTx/ZPNWv9eqtxEn/8RB6i6
RuhW6bsrb/GflvZr5NhkaBgikoVpfNPHewL6P9k+pTTcSa8jqQfYkdB9UseL0HKV
gnhtU/THWPRjoV5idOplN/yAFAk0uEbM+ZOveABUJV7tUKVDdubh3bATsba3JeWX
nyYRyhmZN8+TWUBctsnO8N0aADJSShI65YDa5PNmwiR11TC520uMwlpIt7zxnmU8
FTX89jYw/AImEZyBBF5y13eZI+/Vnv4ncvDaRkZsaJK75pb+8+R1SNrr2gcpK/7d
CTaMMRYvieKlnypfMykep9Puz16qiqg+kAlojEwRcnLKEFJ/oApgyekK1aQkkAdn
id6UvHIk+nbZLvcVkOiBGbKAPxGMaTOhJHbiYUN5SfDlrdKaZGCcJ33YqUjyT4VL
L4PUe2DC51hwTxv5KVG7RghDLOvatI/2C1xh4TOqTMPzIUOTbCuEDZX1dQI2O/US
z1HbNLRUMQTsuFNGHgN3RUKkQiyBy2Gv9G2kOfcRQXK7n0thsakLEXJv661FoAEL
R1axY6oPs75/QX7nDTlUhAG03o9MEu9Eh0TgLiNHnoM6l7fKpht7EoR0F3Lwrpx7
ffU27DJk83bNx6/cw8K3UN3kYiqSfgKZHIV1zKx7dFSitYmk24ejtlwxE4nkodLL
Ol1sSPHL14ZYMrNToIbHqNGzPefOUm7kd/XhC8ntVS7DeK8H9nFgu+Gw0wIryVug
E/sKYYv0YS3KxZqVIhEfs/uJTgShIUfODydVqzVjzRE+CMelrmtJxy/09fUf1ifq
OrVnsptbIIE/iOdC/bvq8Mi6AcGztt4/G31LeV3xjM7MKQYnj38EuLQffA8NxV+L
sL/b/1aOKNuMG+zxPS2n/bycMdNY0rB23xDAMzdeWp7hYe8+JiK9nzrb4o/trzB5
Jxt/oi+29YBlsQWBcRD3AbXgFuA9i8Xf+wLGKjkxq8ZUyTWdG07zxCjI2uZ/nOG7
i69xr9JRLGR2IASUmb0YRpdp3My0yT+QNKnfFCgg0XHIHonH4gfnxZs9icBr0S58
1IuA3u8EjiQnAie2Tgh33j9DlzEwCU1rZ+JrGWeoWXbMIZFPshK/m4JjTmWGDQJR
Evhr/q0NTATGIu1G0kPg/mwQ2TtFoMdttJi9oDtMlKoZSHSDM9h+qW94SKJWxENw
g9Mxw8me/3Gf92PxJnlKaaIL/WJcAPNOJhdOloffxveydXxxz49J7hSpIimblh/+
ETvTeBm7au9jDeA/ZkbAqd46cVhkLHvGADr+s7CAP2D3C9m2jxc+mgYv93UsmMf2
3RIeixypoBkZyTXOARJzhRBafe65IIMDyJlpb1tE+2ZdUt1O8xtdNH3gvcyt2uaj
nWrvsXljuZKMMNb7nN83p7So+AteAGHgb+XyhPDkNj4hc87xEzEnFpN9Vm+Emhe+
UT9ftDfTIW8CcN6hT+IkcqSC0zpM/6mDVQZVZ9Ys07mcMm10J5NsPEd2decayKk2
C7lbPnSmbg/DR0reGeYnrMM9pch9zobWOF+yM4vcN5SY4u2UdmIfs/dbhwl0ZnsF
hDa9cyBoONydY/kpEsubUy1eloa6Nvdb9iRlaxxU8xttRaYb77d6R1CpdVEcrIZ0
6D6e+nwD1JubGb3d09Y1n/q7hFaiG9FoatRPTLbodGEf12lhPuHbuQLS6koM6gr6
3xQeqlRRF8JD/IELntNacCPtz6hMGAqNTDAbM/izFXB/EUJxrbOqqmzfvVnwNlZm
YQIAwmIYu9o39nLae6ERNZAC/v9T45UXPGMbdEq1LBNqjS4BowLt+aGYQulvRL2Y
uH63F9oVaAdI4Rp7PIqVzRVh1mLj4H9BjOP4NCgRSP27k8/Fkl/zxw/BcBeiPs9H
9pK9CxNT5gH6VYfVLktHvJym15h4ZtLRNBm8W2QfLmhtTiCAQOflNwvm6uyxAIc4
Od7ycO2+pfRacE7vf5VysIMRfi769XEm2CGp4eHxz027V0IHIwc3In6pSmNJUuY6
5tt87jAwnOolLKE45VH83Fc0zLlotozA7igpvJGkvc8de4KAmWuqBONE1Sj/5cwb
IAkmd/fQr+uOi/U2/geKJGbHsFJnIQ/1srHyYhXno1vcrfY0mQVPS5AToW6e31mp
E4SJgiuF6cTu9trxRP0u1RtQ3gzmFnntXRd1l6QiytPTTvbHc6I2AvG8uWaTmooL
yUT2wqqzrlVssWzt+VYwXhX4dfj5r12ij6uJLQu6I+DWuDsYvEUBINVBeaZC65Yl
cBxcMgAtfxOEB/oSjUmdJyH2Tzzl9oItdNzAQGm0UOAQiri3JIvWIL9CT9W/mueo
jW8XfPuuuX7NgGmz4sXkGO25hgw0RfkQrnVTHQmwjStndnoerGzcjKiikJjqj1k4
ZFqz8wAVzG+c8oSr47XxAaNElspI/IVXZAlpLmZg0XI0z+V2FhmtmtkmCRZ6C72y
gpkfxfLq4y0+/+CZz+AfUrKyc/LIgFqTHWM62V6KBPESwskar9by8d/1ObPG6Yoo
WFyCn2jf2n5ITpHQ2G9mkg5covOp7zQziWgvf/WPZLd4Vxa79mo6SobrVJ3Pyp/j
4W6TqHvyP5DRRnEbCbSgTDADCECL9rPTB5la04ckiAAuzXp7+YjO4cEfg0mzW0Ld
0kP7F7QNdCgTafFvpWTZRK8ssrOXVuLzjZt9qNvkCClBqXeARZmkLoF6AaHpX8KI
QS0DkTzaoLqlcrSEG8o1V0UH31vKSArxPbmv2kQapg3GCDn65E/ss7nlgzDQl3hB
1aJubnS8xaXNZnAN/4819NyPDATF5Q7xuhK1gEuMRAYTvG2WVCo2xxMgXumexAha
0xgu+vbyNYjTRb3CcrzZm2beLIu5DVdfUVlUClS2T0iBjilfqoTwCQ9buPD/Ri3H
lKY1cEhWyIQmEk1KNHX1lRHH+kX2feHyk6Gn+JALr7sKnG94a2ALtdwf/uS5SWE0
ehP02QY1N66Di6Wz53YNBTEPwQWLiU9tY6tAvnRNTzhYmjqPoxUrUzXQ8GXWXWPc
LAenaCKgRlP8LXdRtHzRTs5zRnfXsLcorhcsoziQkK9ay3oC6ja6F/shIQ5QxoOD
8284whyn//lurMYVuT6UDsTVqFwY49XuCKJyCpJ0Z+rtB0JQ1FxiN1Yfs6BW9e1z
gBlund3cYFLHt8SgCg2Xz9l+mzfwDJYw76snWQSGIXXEdHesfDgEWnCSBd48VT39
lrwty6oVl5jNNMHw6Q9hXTlevbZ7ajHExbp5zI2NXLw7AQV4uvmcRRYGJ4pZbyYI
PRiSNRB0fovIDdqV2UM0/gwDQWGIB6GMIWn80cP73spnCdUluPYu2TCF0UCzc4u8
pnAgIhRdmeb2JAX7VB6oHdcr4TxNQHNn7rKfX3x2TELBjT0WPArOHvJEZFNlH51F
unTDlPJo72JYPTu/4J3bR3goI5Fh9JmeIIAGWYhZa2OYC85QBAvGqyS3Tm0i9UJH
47dCcsF/JDWUnKP3iLaoFXo10AMQvlmn/rYAbNDeLe7EGoeavgURHt3Xwrywgd32
3fWzb+KYvpSSjw/s2d7qfzn5fB6E8z2AAEnrG7QyR7bW6XeH4D5c/E/YTaKvHvZU
TpzLLxGo7j4IEM4OJIs0/8elp2+f3B+FR5mUnyrum5YdvSC4bNmVwOSYtd7H6t7F
Qht8BVILLwfSKURcgxSj1xH+lQ+Avhvjnk6MyAYNda5N+2Ynoqf8t0w3KkK7pwe+
Z5YQLRGC78QYBiT8JStahY5A9x9uCg4Z7jBuu05ZJClrhCx3w6ZJIH5dM68CLSYa
RdlKtj7WxKZKEGvHiKFMnFjfdTYNWe61ceO8///Bu4P8lZy3klz2g9kBnQKUj7Rg
3s+Vk7lP4fwwPrO42veXDoAODFyxdDGq/mDwO9/huCQ4vziAiDeXOhh2YeC+0vm3
BHLuaTRZKut4412DQofSL1P+1r+a3cbMBH3TCDEQkX9lssWX20fYMaPIa335Glk9
x614QkxooqTxyvbwwbw2cSE3eBuvewCuGGlKvLY09R2dXg1Buv1nN5k6yLZ7/lRy
wXXFbQy5CGIVAZzWa7x7tyxXTn75NKdZCGIMmmwi2sWCp/1wmMy6J9klfNtWeF+0
AhnUVVpYHBK48UxceKoDQGkLmjSms1TM/cLkezbJB3UNkwLuyXGfL+AqwbT7Xg7B
x1rXKNuXUzYL/ZUfvqaCM5nemtzERhi4bGO6MfOt05Y/WJ0A7zNeEGPMkr874jJa
nG3R2h1Tnipp7XEbSIrJz+PIikezXk780EGif4qhZdqIevC3R1VtO67Iv+QX7cej
Wic3Sp0nbcB3f4Ri0GpRV0Z1oNDHxDAkdVeA2fwH9ihtBlsjsDt2H1PLZkQ9QZ3S
vXF4yEzh/xI/x8Kw/nXJ3YuiZfGtEH9bgAs5FzlViJRH/PBtYBkGKJtaf6PbBkj0
OPv1CqvvNCWar/rHNyIf44eS2Aqop2VRzmDiD6ei/CgB7+g6z7naqFdf8EfgYCUf
p8XYz1qoOw2sVOQirvmZRnThZskRp9WhCI/quEsW6JY1cPdiXt2N3RlrSsM2Z3Ck
dWSIh2pA7Rt8r61tpdqZnLXZ6Ba3qExcp33GV6Q23vYAcqU6RUw1Gzg2SuzxYyzc
QHjaEOTjk0Rg3HwmN0UQY3YlfMRw1BoGzqXn9/+mdokhWw+u4QCTwBiD9EEah0t/
UJcs1fgQ9S5nkdm7zYGDNS6KKPTO4gQ4b8n5kIgiRcjrhvVCeOWA6TM8BvOgYEm0
Uom15DdwR2hoXvdPRnSsqPct7uqq4SKqdvRGzlXn3bJ7q8th4e4ARj/xrXTVq1ts
sZo159KOnCI3Y/Y3ZZ0ToNFw+PBE6pr4yPI8nq2jyCAAl/wUhVTiLZlT1tuyoH6R
/dueJD7Fxk7wVeNuLys0lK9qGAQkMVkip4nCK9T73cdSOP3BlQVIXDlgO8SWyxz3
Kxag9XPzxUzKYzpgqBEqqq8vdmkbkusBj0ASlstpmbNgZvO69wQKywpAnQhpGiGi
sL5WJeRKOWdaBoS2tvkknP6YqOmF3JPLt21ApakwGbqZHPzdcRVeXrooU4AZwob5
kEjOJCXZvkV8OXSb89HjSmwK1yDqPaU0QjBAZj329i5CsaRmx2Zy9TGfxVLe70Xi
sESMo8V9E7PVSS9gDQXw2cKp4WQyfw7sNLthDw1BGDEUsLmqouFTGJk5LGOjToAO
/cJYzlLjJ4Zz/xjU0RxwbQBVNA2SXhNP06jBolmlgK32jOtTTA6hhCzyFweW1ixy
NS5kqqRfzrl7SfsZZuBNHsFj3nIQx6DIygCypBXWAXFoOfmJgqHmT7ns0g7ZCesK
eG3ED9R1HihnyfC0L66BKIGb1g/QZIoYyoXuAhje0PeMwhy2F0XNTPhmJBWEyNUP
cPPeE0+iarklZyYr/Hm9GUCa5IdItXMvqd4nxGYQ2rL0pF+P2arkp5KhtS2JDdsi
2eGPOSITYQKizO6lK0hCbmptKE2r6xiQTqiSF9+BaEr/BSXU0lro73GwbYeidVoZ
DeQzpl2RBkP7chciSSD31vbMft/4Lv7mBe0Y7db/kBgXSfnC90OKvx+wY26zVFfA
GRcwioqKfjWx7sdNeA3hauWdQ3Fm6we5F0uLpCONq6YOJ3ya9Lu0olUcD9dIJ0Gd
DyA9y3KRAwe7Gs8F+WlpEANu3IMd0zmz5gGH+CuSWUW0ewKDWL9s06fQd+xf7rwz
r6/NWop0/lFmFO9geyNFJfh+ssHWnZgbzLo828jg7lc8Ng7IqWa24F7S2xubgZP1
oM7JYTT3bU9hULh11/2thA/+QOBBi9LpPRwCJD5oC7184Hf16uY4R8VszsGrc4An
Fo+ZacaxBf9plPe93OiIdbeS55xqVLqPDKCwKJXjVZkjKSwO4EkDpk4Y5uQyftCB
b538lNlQm1l9LY+7BsbBbxSDD8lHJKFoHxf+v8VC5tP5zrJiO6BgSMtBuPnrNQOx
z/STHfGOxa8bCdXHKP64cy53de16izgQqcdTi/IpcR3XEEuyd0RHaZTWZsfQqL8s
fy55yhGwRb2GzfwOBftxiMHtfSwzkG9nnMxwjeqz536t30I9SbsnsyNJTyoryLE1
2hw/8ULV5l4ULBxJExrsOn5DzwwekyMLtZxSC/5LX0uRE1vkITpygGKl3liHbaHh
SUHW1o9Y61152y5yFBlaaPjUwaZOUtfD03HCcuMPxaL0m2RNhHT1XJ8Mf/SrllxT
kPDzgOOhy/iHDE5sMxQ+TC2mLI47XS9v8IzbSidYLTCpW3U2Di11oYDiPXxmd/MZ
1ys8/n/BHGmruQgJynlOf4BCvtUaqlQRC6U5jnS6bf6RfZDHk9Qjb7L7MJguaVk8
cuvrfhnyN5MS/p8zDSFMNHqb6Yc96Dsmp4EUXe0UaEQPgDoAQtKz5OJFNEp22G76
U/6v5aNN8wcg+/dsniUOZKwGMVsjOTkz64oB1YRLNuotaxct9HK6Y9VyORBaEGaI
hgtoLEBsmcdii6KklvD34WW1czRls3Ir1UCX43lQDM5kS4u0oSKC6aoBfhC65SZ5
H31oxg0xKSndJyQMF3czxtL3HgwZv+78nFUTWke1iySCH0s9BZlSqv28OO+2FBrF
kCqeSqHTXorhZ9M52xP+PGwrvCNLsitTyLf0oT49glFYYTPppJoqaQiAUThvgwmh
g45S+/XlbT5Ta5FN8OByQ8SzwC8ECrOl8ntooMNqFiEgOaqcUxPJ/8SATw/vpoOR
+qTtq+Cu4RGkoHgflOoueaEMmGFwzlUOaVjzYl08TM1S6dgIEr7TixZbCiCmP+BA
eKSb94KdBR/xPu5gPNtiV+WVRmjDiuNj9DsOle33/K72x0db+TXmtkRTXCEn80HD
SdLH/4sYtZrr5hcIINACDKMdmfKJc+lzHHI2Wq0xFP4ebBvUN7nnxKclcblPAM3J
hZkjZox4+91P8/S9NbQ7e2DwZ/1kz74AYfc43AbaG4RI4SFhVvCxRXKgeqOBeWD0
W7ewFDjJG4PxBE0JrR+We6pX75qrqhK1Vyd3/Z/qhG6qTI4R8xygYIUO5VFUIrh8
asubRsCsV/3fBjP2k30rgsHhsS0nia+vmcpdDMSQb7j2S5Apj+K7Z6I6Nfhs9AMR
FPqJZBgj3V9erkKPDsUe5kZ/7L5dsOAnbwJ5qw4lDjXGYKXl8DWQ7ztmdxBfGzyM
oTrC3gaVEX9C9ukYHGZjEAmhhQ+irudTJ0R4VIjPYoh8DbsDoouGBG5z5VFNjR41
yKc74OQNIvhRCWcp2hlyy9S6rBzHAfdfXgoyzibytLZpPxRrwD4gkiPox5sJieUc
MRjAclEKvn+4DgVtu265sMt+q4rOKq+kJOvo/1XeZZ1W0ZpMd26Vvh2UCXNZXwW5
aAMOlwC/xjAMSMyJbDChOHusUJdLIwSOkSZsLVimIpe1lV5tIcWBIWqVQ86puK7n
ONB1RTYm4/LuBKSUCdVYRVHFw3k1k4fqlJsCIOOeS556Ik40Q9qP+ZmEGSTgfGEW
CGQKaSI8ScDcTb2Z437KvVlJu8oKZJWsjwMDv6iG6jcXmcDtHGIdxHSYmqgesx8r
eXFmG5kKJF3rXnIOTNrs5DCEVCwsxPCebZUh9TSTExotw85dTd5aVAzcrNSgixBA
aS8iIwzkTCDcnSqZBRzd//PwTJTyBREFgqWUTlwMED3YhT8ZgfslxID+6OLVl4fE
SShZvG3qClT9nvbd5kECwVh/x+3RAXn73QS9/s9p7t9oQv1e/3AhaIPM8p2tbBJ7
VQ9lQOAuQnBRnFmrto+7RMDMGbv0kIa6akKeI/3Pidaz5wcq9q5v3Z6kiXJ4L52c
AC350WiGL8ubVpVTImgbdW46NpW73FRCegrbHubkG1KF6JihScXgTDql4CmtMhGT
fv6fH9q/jTJ1Spk3E/qb5rBrNOSvC+1LDuL/WffbsObTSdXYgLitdLMILkdhu0NH
LQgB+byPS9jgDtHLTx8PvjPEQyqRhTuXxtv2ZjE5pGBjBIOi1mC2q/8bOmof0LW/
3trlShUqlIFvUgpCyqt5uoBygVN0C3tXXQch8WjzyvddQtDdB/BjpXxV7c7Ruzmb
bnmO4l8Y+2X1sCaG1014J1oHywapq5noWx3Plc7N7z3goCRx9n8y4evPlLfjuwtl
54LoExK/81LEB6YCOmkJBq2/25PsOIB57B7hnkD/XwkHN7PZtcK3WBWKzBOcIf0E
wILd4dTZxYnO17lT/AXk8eEE1eCbKlBHy4vtYxNmwCXg4FqUHJR7LcbZPeQxjC1m
GIvrAObXXosbUb+SK6+rbUGWMwYjyzOd7NJWXMMo+0GVqaxC5Ax8q6DFcpHdw4KH
CGOh6Y5PyxjgMY9GFTJ4hRVWgZqVrbydR5D+7TaFvPtiX1wjbBA7ZS+p7KilaXIf
OJVMHNC4gCuWfrzsVpo9tAGA8tWh2QQVZmu3+XYLUi0zBgYMDP+6URnrehGBiCQr
dVBsv5fxikFXBAlvxyumgMagz/GnhOEY/aVGkjsoop9m0ctQHm5f/BoqF18DpiAO
AVqWT1pJfKiItP59IiyQ1BZys5ybJJNSEvNE82E34Hs8MejDJxnPCQe0u86nvSRr
CN0b5B7tBGsUOmsQDiuN4pFQyBFVurmVqQ9CjR+TewtlVMhGEEscKndNVt/yynj0
ArWlCPFFXbw+W8rfkIJXWs0Ss+LNoo83X8a2fIFjUrDG37K3gV8wY7q8s5OBFFFB
jsPXEnc8K65H6EwtUEWOa39yQSyqbobSSSpwqsMgMMjP8Y84HHBzJq7FkGOa13dV
9v8umbJQkwxovnGdotDNCB5VcWhhznh6Rf2GwetcJQIGqUpiDTDOSSS4xqOQG3bA
6Om3ZiUkG8pFEOFmR7c7KU3OqVOWuXyOerfT8gJMVa1qb+uDPb1B3KaaccvNGHq0
cjfeCrdo3y9mdp5mvjcdT6PwSKoZcHVJQqczJIPEA/xNGA32TSpY1xXIRHnL3jE5
2m9Ft0ZlBVqUyNJZRId5FnejOmrwjTuIIXXZ8fJib+yT4d9qs1tapxcYMIs5f+ot
XBOWMnJ/Gm9gW2TkPeL+vufMkJtBuy64djyqbPkK6siEbjGXEXUyNeXdiWobV6kZ
x2TTFyx1cQWcAyLZ91d3NfNKdqcQ+igMS8TndZ2uInviTpy+Fbz4KdSEJPBUOUjA
0DUDVXqf4l0lVTlL9ftWyvhQrLiztoXpBFfpcfxDL5CZrbadzmnUH7b3vcOdo7e9
tzpLuhTd1P7cFGc/5WKqg9MU0MIdm189ra/+bUVjkrE6cc8pjQqBKGdJGZfyuojy
DhOSOOGGT+N9lXVpeNR70WJkKW+YpqYd7Wgm7MWkF/pdNxZplCquwITffQRlw4ne
a0H6it0ZjowPOfklJAW55hGCBnm4yK76OKFih4MJXFSnej/K9VZ8OqPUti6iZ2fM
0IgEkdYMrVc7q+VNzpZaIZnhQ573hp9POWZHGJJ4E3RUOJvJn53BUSKqvbHu9MkS
I3UoLXelHqFIROnWilqhVxjgZfjjGIUBTWYZVYn+oAVNTmQMLCE7gfdAXQ0obJbU
zKXns0vkH2bXnzzZqlEUjuFgTFQKP0+TedIN4dSEgcnE3JYHhsXvRZ/+u1q37mKz
/kq09u7qub9G/LrP3pSYZ6YqixkHEoR4+fHRyVEj/5axpNB3XrADw72hCeyjiN8F
fz/4LBPasFab3m7MTgSvBMYKG5j1dkuYtoK8umr8ei/rpLajqlAnKEBLfJHOE+5Z
dhESywOM6xJ6+trbh7HEynHBhGmqNyBhaEpowU8PZZVOZBB7vp8YoD/AYFqCLEMG
KtOhm3O0vTvGQq2SLKnazmhlGODzIGMQz8MGgnyVbF9nrh8zqKSsLFBkK0TT6sDT
srKcYF2d7hX+TYknfpaZA8/RpfEvPAveDn/vUob678xFFvDLcbXKgATLUMHHsULt
Rq/F+az0NNTX6VfFqNp0soqeUkwVZsdiJgnJPAP67sRtZKVqugwjd0JYbQ68CZqR
US8bi8NVFblQKeS5biy2ZLnD0A4E+mCtX4T8WOZmw+K9iiJ/rnQA7BNTnQvug/1g
DLCoFQB5e4PqVQhFBVuLn5qPvMXJOb+Dt4uWFoVUuNyCQixGTEFxqILBgeoqXORh
4ff91CeLvHAKsJOrCQEtr1tb45qk1h2EyoZaC3URSQwsyC1t3qUxVm+bJ4TVNR//
TOON9Y/EvHR7XM4n4xd4UuApf6ye1e6wJyelG9L4u3w5e1Cb8776xI+AFJEBnM0n
GmCOfYY+33Jp82m9SeHwTlL+sypYnlv1TRKZCVQb+/XNxa9otkOb7/s+hYlsmxTB
BljA8b25CEINjs/2O9J6FcpLKNEFXJpxbg90eTb+xJoagcTcH9Jmx59LClA4IKmH
zNt8n25U1ImggnTSvsCQnK/MNpMdijVckTmJfqYdjXKLwoeKbM0b7hxSO51CtMJR
y/+YRLilX11DR9L8VNyqLqa9KPyb7K3+88JazZvUjXwBcml9TRZRyRKDAEZkkmvw
V2Qzs5V5Fnh/bRyPtltV+zFl7NRnlIgVbBz1Aa0NiBZUNaQ6Ba+TLJx5xe1we76Z
on/QQKQnQko3BHfrdUYLMJAXsoyRsnApmRtqmhCYH2XRccEb72/RZL7laYSMGRGp
GDKlSSZJiT8w3azqLAFts5XL7dvd8AVANLqfTiJMfMJalMA54+dzzJMrq6NJfrrd
+gw/43BquI/IlO3R+PM0sgJU9XiQ7XaZEpkZANorTAK+V95ZchBEp0m2chh1r+iF
AoR+IinKtuzHnwvLPKUPbl7mHGh81eNXXMM1T1j3s9gsAdBeFNdVjntkkya2Bseq
SnSsutR2kFtY4rNm+uzyfUjkwE4PxSW2gINPTSTHSQn9Mv0QlL7XaUIrxSPqI+eC
i699RMiSQBG23Piv2tgIz8RhdahV70eo3gaQQvc/ZHmtkYU7aiZagmOJP+btpB6r
8OhAQoDXM0AXNpZ3pxAUZpLlM9tHGhgudaBaU4IzQqzDHoTv1k1K7b20L8+QGdSB
UM3KD0W0rffTw1iQ61Xd4f59VlyOvK09gt53bmOc0rGxwOJPVvim1NjVg59+2737
Ed7tmjEH+kufo8C3VpN0iekKpL4jKgMgn4J72ix86GcNHumF9oqGNaDy+6e7IDqA
Xs2mbYWy/dob6cEJsIj2z9whP7w5v3Q0QLT4o9Kt0eIzabE3BT4LC5nqKhPUKCYz
F9lOKLwQjKuolJzY4+TbTqsVsJvHRcQlpeIaRgW0AFeMttVDlOm5uWqREG5z//jZ
21v0ovQbtafAgjWETw04XpiQHzuCEj/cx0Xat27xDRmrRnl7dc/mIQ7cYRwH/+mc
JXcr400974vq7fCSM8sSxoOPukqw/xdfPWCAfzeLqmIdUUoTVOk68hPIrSuJcbrZ
UouHHFZ8xSGBUPDNXdvdr6A7Wew2CbY8pVaQv7e+7WFMjQqzZFp9WsZhrQja42r3
QNpH+FweIUcpurughm1G1qgTGb/0Z8iORsjCXvrcj1cIaHiWLhLO4hsJMZ5/xt9a
B7Nf1JDSZAArwOOOTcvbcJuWQqNQ12gFbScmlviagrLY4/jMNPY6krXWz17zdNzR
nTf/9ujttf2qNYfeYWek8aDJq2eILmQ5H2YeKnrd/XGgrxBH6LB+/bA3Nsy7YOeC
4cQbKrkVNLwX3uXgPbZTSA+DiQP1R6+ko2pFxt5mvHKJbzRYjGgSwTlPpGcJw3S3
0IdU12JEvOUNwML92JF+1g4hU3BU1fEBEj6UZ5cNSFtneiXaYHVozaXYdPedIsY+
hrhNH8SctpjXJg/LOosFvoE7CrUPRZvA+K462fLAxPJe3/k+uOgMjNiSfLa0scnM
MNJFK7sapSr6enfyWjCUguqXMehIao1PeE7PLlcae8J6EbpsW1HljAPKkWgC9FPC
VFRwYgHvnrNm9HW+eEd0vMLxs1NdsbDxDK6dRdcNEbhnk1CoYzQjXldoFPSmJKBX
9oZUiWw3tuKwk2TfOu8/OXf+EKwjKyxn0U9HHT15QU3CcCc1tbATPXOBva69c5P7
dRBc3Wc5yS1OZJ26dLPN19oI4WO5R9ZxDhJwMhDTAiRTybtfTnslAmdvLD2CGaB7
fgOHeE7EIj99x8StwOQ3VNoXpIDfIuezG4iPurdRNnKN8v3Qjl68SQJQO3nPCe6K
bFZYzQgIhwgnYEQE2VqbDAIEe0kty3u7dO1c+JHrTU0MT7Vewei+NkwJy0/1yt8h
VFw6bODc/vaUHQqEr8nLpGQAeIYJrP1tcrTLh2RSCVBlqhS31OeoRA8NORb4Bf9P
LWSyhsSxtE6mjuxCNgDI4pKCVu0DeYTffg3y68BT13q3pZPgK3J5JwjZvO9D1zw+
JlkQNEhZp+iCBZh767xnW184jE/dvrkVyjhX9t/IXnnnCKGN//Ai1ahzpJwornLw
ew+gu++az2fOB7GeSVM5H9egmj43OhHu34/eH/iifCGMpDsvI1friHTGeF13cNUf
TtTIb+4IA8tCuIqsBLqrMciletbDEDC+zkvmw9G0x/KIObpIP84rCUmT6w3ldV14
R0UdCRJyXPqoEYp3tvUp6L0GuIVkltWi0/0yPbVGpdL6fHT/GCdrMoQscw34rGhe
6GVipR0Ym6nNgmjvnx/Mmo5LWN+7pSU5W8rMkX8lT2pmqs2IzU6s43/oIFYaAwwU
jGjkKio9Ohg4bFW5+tWUY62O5JITq5gvfKmX2hFEgu52in9EZI91yozbZqIphYk6
USC6DMNGthNyjTz1wIX/BbAQ3h5wuR+n5RSx2WIw2SPkZ3TtZePpmiIAqRaLIUUJ
r6e4dPl3Yvvs+/cm755tmC/VVHr3Q5Ig4FyBcgigkWLXef8ZT5xBU3yahVAP9LPz
ZeERyR9ucxK3MZ/TXW8NUqnwrzeYv41RXZRVK9gkQuuVRoryMX61HytSDS/CWCl0
v3KmaXawv0KL8b0nyzSY5mRCSNryAU524m1+ogKETlX7xnaZwv0pjWHtdCjQeR0o
pOC0UbrrSC9agyNNao+SLhhaxlR8reJHbX2KczkKQSEjDc3igd1HrdxObUUF0TrF
0IHneWIp+V6OoCCgoZhOJkd0898FDALUrvGsvq46PvqUUY7/Y0CzxN00jf9ciVbx
5f/6R3fwW09kMm6q2+WW38NPp9F0Skz/ygD2bnRycycvbz5qqIgcYRwux1JKdLaj
GSN+bSD3zT6jpMtXRez7X/ysp5L4YrcoiS5a1wXJjFGzaaLLdTfFvOB1HwLHRIq7
dmoJDUWni4OqIxkjT0Zm9SBuXGGNGbWlQmgb6RB6DAQvUchKqJj1icE9bWloL4I/
ilklgKCQq8WcJ/I0saBvdXqsBlnuS4MkQMe2bL4BUxftxi9DLWIF98RZ9ObCgFjb
zcW1P7zF7ZZ9DmVbWqnBg07OWe2iTMWz0qpecDO1bNQTmg6C48MwY6QyRnn/jBb9
ZA/RsbUaMwy2HRxyOW8WmbNpUFrzfcljCuByRtrNkjn3rELHEv1+dHKlz5cFj+zP
wQ49IrAyg1a9E4AjX4UKDCzsYWEM72dKiNBCv5ZCASnyN6I6/ZhdhtVTIO6JfxeH
444iZ2CNp9taVBVHe3TEdBiNlGoL25T96PzOcex98XRiJauuVT7J77FfnFzaaxNG
pm4iNbU7D3AXTyzI7jYuextTdB/z5xty3jfMNjls46hhB3ooVwONtrMNsvAJJJtG
YxXaO7eqCifuDIhn4oOhECR8tiHSvMfngLj6Q4eKuNpQRuMxLWGarfh8lev8UQcF
8Z7FFBCKxl13ZF2adnJrThbSeKrC1tHr2tGeU4STqkF+IdwGTibLAh+gReZKxE+X
HSS5SGwcmaGsgG39r2G5MDFtmCMeQV3L8W/P1ki/DMFY8RAAioABHjXTD7T/Xtdq
RQEiUuyx/O7SJS4tQ6hLdHjFoAhunFbqnkG+cySkXgGT7S69mY1BtWl5Mds6/avO
Fbq9slDWeFeKOr9EfG+sl7SH0hPMUicQ0nmj1R5wyIGW8rnOIcLj4cy7BAgt1aN/
UdtKF6KweVFauZt53lxOwRITX/qkR9pW4cpTTB9FgUJ+afjsaCHXiZ67MxJX1kvl
4i7vHt7qdnp2qCP5VrjIl+2H8BVBVsW2kOx2oL5ADTKwVB1PuS75G40xFk4OP9OE
ibL/97eNB4Kkfdw0bMVfPrBcn82oBiOTH4a31431jU4dVGBPvKGzC93YfB5VjgDx
RybeURKlIzsg2GTTA8IfLNN9uOaR7CUIAeK3JAUICcrp2ulgbo/iBg3amlN6Il8h
/+vWWA54UuAZGXmoa493cQMojbKCLC32fheBG7dNbnOFMrNaMC4DJLUtXuPprQt4
2aBt2Y9s71UxbW1RyyMhv628P/BpHL8GcfugWx9enKnmZ8SqQ9vcSfcHnK6TNqY/
WJwc0tz3DdRTvWh+16OxtsNKaF2ebB7Ou4Ecd0imGEKNe8hcxWXEz8Myz2kHy78c
ZOMkWQBO0hCtrbDZxJJ+4mZRTOuPszuLL2FB3ojgLFtg+Yoq87MbCtid+U0DxXem
AMlDF5O6d+yKVuDVQzTjiKBFQRmVFVKR+wdsQaXgGKFGC3+zMnyt1d8s1Pza3yrf
GqZEImNSpINymVzxWi1H0MbFoptItg6ONvkDLb2EIbF60eU+MNRXF90BiIoKghp4
EtEL06Ow7+1vxLFY407L5kaMSXrtgfuSyHkz7vHg8WV9UVz3NbYqNjexCPOcxOfv
2o9jzQ2WhaG9XWAVXyIueRRFxoD9EWB5P19mEIaDwScC4W20Nuanu4YmFRxUquFD
pCKuuumASthz0orihNjh+oNRIoy1uyURuEsk8PaoTN6jUFExi7XjdDQfjfTQpQrk
68j4UFlTJXOhCIY4y6lHzNz5T+Al9uMCdHGgLbvQwzAE+AC7Rw0JPxYvilmqI7Xr
J08eOhPQKZhxQkem00Oajdp/kMy+QhhHdbistMTqherPNVxceztZQ/wFboHbLfwF
q2KOBeK4Y+9Y6YyIZ/ttFy9f31xbWLBaLr9KFV844tswZ1yZDtUZzLzoYBb5wdiT
a5rvK6GXXhXZsqyLansrmhzkc0euk4w9lDGrBdkBIuRyxZB/xA+kRcA09gUlZK8o
8pp1zKQU30TlGLGH+qdf/E3ANR0MPZOUI9FCnUGwXfiDdL9yuEGYuAUBQ2Sy6r21
lQk1uVdepqkywtHS+ziNUnM4zrWT8p3zn8lbg0hY2gaGfhyumBFCgZvCXg+/pDa7
zcLIG9epeb4OQ6EYGnspyegzxCNRtajXQEMaYGUOs7KNufxY6w3WCFru6IabNSlO
1TeGIFqTiV8yh9ZjRNS5wBgEGg+EAo123h+/7dj4Z+TelnLtj1C+Td7X5uVmAfuq
NByoC7CtiQW+RmYuNHXpsnjfiEkH0XnmT9uYBQb2KPrdtlCLRuGnRQ6gFIUmy2uM
isgXiasVVgd3vYcbVf8aJeIzlbq8TCF8Mxod53MF4BRAilpwUPRoVwcfajH/aJ4o
IT0ayoB0xcV2raXxadeLSnPHiWJTRuNkYV43C479vePgckzsqrNNkjAVKmk6kZLz
HyhnqldkiGkX4xbW2PzOcvBwTBGzj93E9wByHRPyiXUgemWieDtAOyQJYcgFJZzA
hYppB0D9PP5YkNH8/slhJyMx9S0pEmQG8XdCH46XJfXWfPEZWmB0O1shc9sjKIwh
aHneH9fsV6SEn1gH368TtF8y1EDBiWjN0iaf4PO6Bj+F0VP43SuRCrd741KnAKsa
epXSAdl5MYdQcwq/Wn9P0HksOh8kpH7sftP1RasQt2BDP/5Z6iVKBPJabhFOwj3z
vLRHm/MqhViXeLDC4Omyw1cnjUApmp8Q0ppnZbuFurXab8IEHBQlNuQbnRV9r2OV
g4/MNJd6fBWlmpJJFpg2SY8oFujPHOhaNi22nKSJREROg46Sdcnw7fRGkp22ZCrp
82PIZvWja+eG/1GZGWkJNyLVDGg5hiQEa5cZko0TOPpebi0Ode+i22RTvMMsynRl
mlqwHckkeYkTCJE2FcN/kxrHovGWiNPhCtrxzbILPB6ZcBUg4D/bm+39KUb2Aql2
SQNFYbDNkJdEwAe0H2Lg7GPp/ZYfXFNPvMgwQPbeTe4cG6bRReSiDQJ+5tFJmsF+
lm4lOfkYyohOtngmFuQ/GMf2QmElQWgNnJM1Qo7UtxZeVgkdi1SvhtlhprEA+DD4
tdV2QSYimabq0ilPiFRKaHF93JqG9YeJDAUKRl6hKUmsLwRsSFrPXTN19SPAy/g1
y+zbvZDsWbySlT7tL06GyyD6lxV8lZA90v/Jwv2ryMLnkVQBBnM5huV8faGulUi6
DI/r9EvodKLKyAmhC/qXijHdiksPybfnFcZoA7pIGdvDox7ecvIXUbqy9RqWHl0P
9iKwStmYcunEN5hkXqzVt+yXrniVM7qu2M4nb/9eyjtbQ+B0y2rYY3c9vVxn0GKy
CqYLPW8K6QvnESAFPRHJfSrPRtGUo0OR5q8ecRDmbAwQRZepoEh5P+l7mAl/t0LS
g77VP7FP05+u5M5ahZlKE36XJcbhHrrxZKOpxJ2x0yR5aBFTN/khpDGtF/RnNBF1
5/GtjgNvBxGd8RNnL3/I3D2rZ85jvY06l5OX7Ol4d+yzQ1mJ02wO90XkT1RB9Vbt
9LatQhNhHbdzjsYMNhig6dQpRAVI3pRmT4W0ySuNAOsn0JwK8LDCNJRnRBVq9VV+
ZFEwmrDdIn5Wtc0OSMopgPSbc6w+TM5SMm/JUduHXFhmRexTGVtxOG+dc9pbhtL8
pRaqdI/CB5nsQzRHvWd7sAm0SORHL611Aq6iwXx4K3w4debOLVUalvIpTlA7Mwfo
u7g1J+qZot+xW8ExnKktNvucaRsJa/B+PPkF3aAJuqlzfm9/tigT//r8XyIxkJFR
fr2lfuUydDaRFDWnXPQ1V+LLOp/LUFJPGCqaXIv2Y7g9kQxYSj56QLRVSNPRFkp9
98u1l55ZnUUfYpY7vredprfiShuWm7lN50snJVtSRoCpCeO5SSqadCRIyy83fTfz
gIIh/AV9KLl3ZJWvgM+l+Meovd6nCWvgzTcG96qS/VcLaT8dO+1b+n4sRK9ht3aj
VEcO3e8WcAWVLBYHztBFtdk21IG8b65N8J4qbAp5RGqzV4fIhsjRDG52NEYLPWpO
n8cmV0yXJhPLzdOC24kwNNzTWmm7pM++wdv8Un03NvuOb+v8hvcaDkHU/Ich71yj
fBeYIpGOY0hJz3D1zRQGvXh9jbOEjpEJh6JMOFQYsPzlSI1y89L8elZWyaTt4q7A
kY2BuDA+zDGLtLiuUH3wep+Q96E0btDk2C9CGDqMiswlN9tY3mnoNbSueS5lIoxt
y+WozzG3TuOSdoeGtEwkT3cql8B3Os21WSjXl3d8INQRyNuKBvtT+30goc7w5jse
+wrpab5DGt2rYWZwF530kVbKLR5Zzy5fFx4jmiShDB5ggTgmCzCxrWc8QMdZjUWk
vHz1hTWSVFlFrwEqNCmT83z5f3/JB/EQikn/Dqs+hr+VZjHaqAWBNxML9FRw+rIl
mDR/ai334MLm8miicIQeo6bExijTufZMBgu8oOYMZ47LTMDhgdS4Gz7s1EdlHmZx
cRyiWFu6gOISOPAfGaXPh1jgRzXkYBC28qCPLWEYO1V+9YzoB4p08+qIDDMD32ag
7blEqUmB+kbX5dBTXhjFLF8Ubvx8acoKgjyX3anO9HC2NjzvwhxmrhqwzoCcNgjd
8QrzGmv7D9UB5jLQPYY0TVRl/ldeUqW7GeRgtRqTz8OejvuafJsHGM1Wxo0rLyNB
PjI4AmzQDZjtGV/S/+Cr8i7KIYmpAtQL+JljJvbnA8OV90YjOgDoblmmYgn+EEeE
p2QEzXzswZ7HgR/Bsaozm2/QpfRmUGxzPRkfcNVxthyrd7jaJHLerknGa8mQlaXW
HVf923eLAb6sW9S2yT/bm3YyCB1qiutjzde/TlNNU9/txov6eH346EFx/ZVfNNU5
G2kHn53LGJoQu0/8tQBfvVAb2hg0rMnxjasTmVQpCJ7PG/diWdPgY6o6ne6irh14
wG1ykcNkSeYIJ7+kUme69wm7Hy5stBL9V8T/TbIw+OcMbcRdYglY4BqvSdNQa1n+
DFpzx+zgymtPEcM2+MOo7wqKdE88YemvIX2xapAZfI6TcVdGG5260rW2+HqpG2eG
UBAAXufAa31tmr4D7vbu2O6tZLIh+yhHN5SKNRMr4g3WQ2TmYSfh/xCHQ8vnqUS3
pUwCFjBqO1ZHsA+RnQNDpdLDeFImlGwlb/JPcVAfbBMy1CcBIwYvpPoRjQGzCLpJ
a4SePd7o99uJ/vVD0nnYOF7x8nylIXZPE/kZwGltgPqVo/NNwfvXQBCFPqUpBJbg
YX34ZdX9QN+Iu8VjUWk5wRJqvqLcsgLxEp23xsMsY+l9uqBMaNpLSnLnfJ/JB7go
5VqI4HGwOTixmN7FM37a6uyJEtVgEk0M3yMCZ3zGR5yRNLoxK6+JCE+N6bET0zg9
BmDjOzJwh1DYZioVM+ati2rDR7jU1orvlNJp/ajr9MSQFny7O15LW7ZnadIWUFjo
Vd+DpZAGMaIMPMUkocg03B2+58T/A2uNM2gliix+bDQ3kg2UDt9bOnBEe0VgHIlV
t/n/kd83EbICxMU6cFp5Xi2lcU2z12EPTUJBehmVU72vHpx179d9eE+2bYf/EJ49
JuJQbj0HsxTHv9Nk5nPnZCZfnKZtshGMgsfxJmUOardqkJ68qBZu4FCPJ1Ou00rc
c0gNtt8CG/HVzXJC+XptiHVyNbbN3k2DPZ8ek2ixG+//okhkmhoeISlW8gkoBUFj
kDe1wrFIJiVAL5HPowkET/CTYGFeYEXQ+MMpnruOk7IbhLDxiz5KWfxooasvgakb
UmbV4hNjqMSBqoqPVboh3XAUIqgMAioVNfZNED0oAUK/yKRBDXPnqqh4xyYqq4LV
dw/yMrYiLAZYveYTzqTm+cMtli6t0h4EVgCtuUEgAGLTFtTZ/VAIh/K1RDWeAkGt
P3sTVrx/eGI5cc7Q8xm8G6YwVUWBVmsCNTusp1uHQu3JuoEmWOcwQX8ru4g/83ll
mX97gTZ+NQt3wdg7THLTs0wPk6f1BvSWTPd90A6tO6SyoTrbG5vF+jwUE0lYd9Nd
lq+mE6QF7jaGmSHUWI/oI12jkzKm5QYgzDz9MvefGePRDvZ/wnqlU1IPoKGVerze
jBW5UA1/LecT6bvH7M90l+vqUQWDDY1g1RDIRHL4Kdy6aVKM0o28ltjAqCxvwMOY
YT9kVTqoRBl+/AySkwTXXBpl/HRzhJTEpTEZiQ5S5dn09NDYb4tTGHI9q08sT8yB
HmV4f1tuTAmPgesK4ABmQIqrZQPUAVN6oP6+toXpmsxNloLYmtnf8qA/a+7t/Luk
JcvqIp/gVK435cOilT0EOMNw0CBRTmZVr3spXuYyBpzuZ2ChsqpFpjjYVZJl/B1j
wtXMyA3g1ERcehi80on/hNFIIAAhF62xYdTic+pUCUN2x6daHY6RyyECR1HSwLsL
cMAqEnR3/qAgGjkh16sa667FJPMCOxqKb+pNEDhioT63Wj/HNKrge0Hdnz+oSklM
CA7OCDtwXKS+1BWeMH19jK6TvfF4I31c5XO1koMQGGFqQQ2d1UIXrSkUNtymDuC8
Uy4klnEtFpQhTFYYc50oLRilNdVtBadkbCji8rC1LEQYdHoX+BfGx71QePmQ9Xx+
F6+JqRnTYbczihqvAa/6PtxUsAOohNCVsgJKw09pY5D8qWlkkOfMS7fRWBqB5dFS
mrpvG9N8Kw+OmiV6veg1IhWtHiBBbXpnZenjz7kvOTIWlB0tH6CgxtU9Er9RVfuV
f9N9I8qQipx+FLDS8ghMT2CH5JfCPbbYkgXyge9ZeKYkdc2MwDEHqq7Tp0qlljyg
IjtrDlno81WR2IKTIY/faI/I6SNhQVR2B/s57z+1/25O9Wyig7EjMSweIFkruMC6
i2v/huI7IiCE2U6TFV8ugcylyo64Vf1iuAkYBCmD6uZk6qHQoJRIcQ/6XGK8lgOv
gEvdF0I9ODSew4GYvXKbfqm/EbUETlUB/Au4tM7HgKoCktDLBptfoOotEsR3aVzf
grz2b4rR25SB7Pn+zSlPMIUqLsXBM52FpbgL9oJsqtFoLV+KextmKoq587MC5woA
H8VmBl8wsI7bYA5g1oXQevMPcZ5Z8lU1w2ngjfWkWIyqC6IbkvfuSvp3IHu3+F/f
lA2olsK0tDsh1dTWCUrveLiLDSx6g7V+X+c4oXQ8Y/po068ibvAD+rcNR23xyeQz
AxtAw2GLKnR8wsb31JC47Eoc4GVOymjrKi28j4TNqy0ktEM8VziYqbcxoYNAXKTg
czLUFZlTnMRVuaGRdGEdMrDRDIUrSiRQP2fpAwss5dQ2yEuXXvAIgp9ARihKFXku
PNnT2wCrs4gP0a9yEnEfk5AyiRVEq9ktMm7JaxYsXPoPKoigAwFlX8eI1MCRW66E
fMs1k6qcb3EmEMDF4ZNVgNeO1vbv/+3B+FeQGJLnoJGkxTcXmC8ATAoDHZoGY430
mSVAV4/lNvFhDK6lV2hJF2iFzmItkafQk0g8Dn8MFJzEYR9hNpDtTgdAV6Wl87Gq
elreti9UOvUX8YtjG9KNVwm70SsktDjzUFZ1SLxpNLVTTnsj/sYQpAjhS3MgH8uJ
0Pdk9FqtFlAjF3mmstlh2D8C4qGd/wq/W5XONOCjXrdJLGXHZQGzUV3y34Mbb9aA
ronkVUKTFRGbWRhbyz+S+Ajq7SdMLv10nqIvSkmI9bZTEIzuufMh1ZxN2CREytVF
mCg3MYIQ+B/tat8tVg9zOw+uU89W+7DUJnTFyFA0xatm9ykPFHqnkzmciocfjD2m
f7XQsrfbqJ4XzRchAAh3kNtMj86ybzQ0oJiMHNE3MxT92m1307L0YnLogDxVVs9K
ApK3U2QtD/xuTR373JQgeJ6IBwX32juJr+WMpLqb0mXFUtiF20gkhYqFygYKDEcw
XeWrEBL+6AQfZiKhZdUM7o1j1MTO919thFaYf8Vz3ovPOUx+naEnzbL4KcP0EJ5q
sWaAVnGWPia5tlmQW/9IZNG+00OBY66oQS2dZ78Al8iIDoQRNXXWH9UsjCJRK7Mc
lz163orwGqc7eqm9PN1Eh293u4embjpkXMSXUgfQzX2+behvx2zV30D0d/BUX1/Q
tpPSm5GDPR44o2jNu2QhJtVY6wNkVxQlFT7c9azei5QnbkOT4yOyuMkLuoMNZK0o
leSsiFPVnpgA7+PyBCPkrkEnwMKfU4FZZ25wZhMUugHw6japaHP07ESplh1D4VTc
d2ZFd7FWgvrs+EPDXzkKssdJCMdI4Z5RbZD3mpQ6+Y7FudAcFBRE3DG8NXUTn9wt
YDNAXADpxMqWXAYSPNGihUsAXRwk/3zbpjcCGZprQHryyz9HLjeYIK89k+rRaaMf
d5swG8W1VJRDr5btpl003P4s2BM52V/ShKGQ0JO0vSaBNBwLEBls7w8xPlK7ZXED
exflulWNjFZo+KhrW2iuTMhM7UqAi859rrIfZfbWR7Cu7pFh1rJrmnhRfpjrSBrJ
B24XZ9YE8RrycivFxjgVOXHUdo1nA6V/JdN1byijqNJC8UW+EtL/Q2vZdccrG2NJ
oFqsxtCRdz73yxFClmFf+VA44XnsVvkCQ9AEEix2gl4fDmOKG9n20a1kLk/d2hVQ
mFA00/L0dfFisvPghYkDElWE2Ap15SJMD+xIZiOAK6RiD9DeUqUCRMyTlcbONxCA
TEfEAt9F4KENvjgBPX+311SHjqHesGhm0bMto5oU8ZBZ7BR6pH6W8MyL7krhMSwd
fRSXlVuI0iuHQ3JoTV1PDwhEMf+LV/myHqcdDX/xEozjuKj6XkCgVsDpeHBuwQi6
5lcidsSXbap4paraZ6YdRkzdkLX5ueVoOOLHb45hJI0HVy4mjO1ZM9N1dCOxQwbB
3SjZARFwYQkDnTcQ34WsQZM8SwlvxROZr6La4BBBb1/8gtD/knr2caEzvEiUFPM6
a4nXzsmbLFrzp9VG4rSlSZwB/IXi3B4QJEZWqq/eQJEPXsC1LS9QP1Eua2gaiETZ
JpsC1dYza3+eWqnkzmXlYg9HoTqabAn/mgOa71L1E7Ew/8pmqectWjfRX70djIJl
O2KtUAxCuzPEokHNtBnGhXKetPO6Un9phCVQ78m2urISfMoFW/R8dmWDNW6Ne/td
XrlpxBj0tCJ0miO1vO+KhkzEE/Pm2gKzQMy20QOgsMA7GpIOoW6DwGqfqki4lJop
RJ+NMNIVBGnB4gMNmloFjhLbauZoBnYG1279xNuxuPGlA5Q6ih/HBV8QJ1f0Cq6v
FQuleU1aEA7GMZszdHTPrjn1Bc6rivmSwkc2+WmocY3R3TuhdpD8Z3ilU3F++Ner
fJA+vzr7XXSquCQx9dSR/YZbLKQLRJGeaEo8A1sQ3pO9ESAnkO76uLM+EjzhWQgX
bj87e2kVyLEWHU0FRm3Z4CYZDI9gryGkYMOatnBS/LZNpPfobbrU2phDxBL3KhSh
DaXS1VfQzJPa+DDu6tTdJortndwG1XdIyVT0m0n/W1HBCc6UFWrzmDfYWjz+Iqsd
WqJmI7kTPuZn2coLpdJ2Y0vBfjKBJHQLiFj8bIOSNWC49NY49HZT6/PmCXoawUGu
RTwr9AzkVpO7+7mFwQYvRMRvHvj9eYJYJpJmCabw4yEymLU5ZU37GXMd2Pz6Msr7
mdTQTUjHJMW77cDp9S45Y4OiQvNuhUDp/boiAJOvD/7iZF552z+0VvIACSpwXTs2
P9wt+nQhaoxAVDKinhimW8eLi++b9Pv7MY9Pr2kDoGSIGmUrHo976kBMgPWZQJ2B
bHLubB7H+KsNkNO50pwe/k/7d8+7nWAVwOLcOGYqJmzoQTfHXJjKgEEa099w0ByR
lO2FJ9QyRk2ATQYGirFo8suKnWo+1IjJ446Q28PZ+aA9n7pXjDgA3LvliuiKgoBc
fs1PPC3jkCzqX/O99v2Btp6yqz7X/gHz2DQucSel0t2b6zySAS5+CtIpVsr2EaP7
tTc3UBiafHGvxQ77VwKmysWqnQ0wykuHAEeIoh0I3LyrUKEi6RnSM4eCe2FJim6B
fyP/GBQmMFP45Bm/Jzm1hpz2UD19VPdg0AGPOnv3YjuKyT5Y/3zuwecim45Y/Umz
Kgk0qJgv1X2fBYx4zuB0iSanS+mV17/mCZa8R3C430V8ElihZofclYyGlbVcQJpk
FyCCCskoUqvyUkNpDcdvlB9fESv5nxZUVLJ4CIio7fXmpdixZ9tqy9s1ghMawc+n
W6z5EI8o4oISzTfLe8vaR0YSWyPLMBzaUQyyMg0M/C7X+Tiaue0IeJoj8U81cAuu
KVuU+BYqgCxO3xMwMM86+QpF4usGC+g6CvMN8Ug6b+kupr2tIVq2kE8i10uI7Bgi
djkriGSOiS74Bbj6vVi/G30f5OneFHc6XeA8KLK6hK9bABLOlovwLnZYm2jXFFOP
kI/BaLQ4+ol4AzppS3TDXHCXyFcEIuFU3mDchYmHIqe+4f+QoEyGS+KT+6YpnERg
0HbxELEM16BN/RJHXgjDLkeCDV/kDz8bFo+kJjnfF9/A3r22rJm1Bcmj+YTDRHpk
mBM/hLnxxprHzlGnySJNddjgYvu/hejBhR/gSNuJUucVdETMEmhdFrU9XAFfW5mL
trnqEfsyOeoeFLJLvy+2IXtCpuWXK24A4aDStuVTza7Vb6sf4PyuDJjofR2OrplB
QUzYuvKkteUOq563BUUXoh/2wYtoMHX+yyXr866vjFs8xi82TmwA7ekMywgZ7EVm
LZ+GHKgkCliP6CrtFXmT0eZl1rmA8KxOQgEFVO57IDuN49sMt0zZEMFxn2v5OcOf
eEuowMR5gY6/XHupde0ApertdpkgN04xYKPA46vlw8ZKbReLhsVLXdaZz7OTWer4
QeBIs84DBQG+6ZIKO5YhHmnSru2h8RVvNVZ74JN3UNZp6Bq1h7B0zKFPqlQoqywN
m5NF+3P36rhEnTciyb3pzDgOny1+tJmuBVmVNiXtoJPVs+QLG4TTKd9EgwuhOKFY
1vq22NhJHvoILDiZSmSENK3Evgf27YZIr1thiK8MdwO4K9qiOelA/4heGOWOzbIf
0M3HFfGOHPcnKHKAYCQkD0tTSDIqqvjMHZFl4ZX5jsl4GJ0Qzw4LOYfxvLkHRbq3
58ljBa05UgWIxyCovsaf4aRyaBHEvFI2wBin8xHpOd5UxBQMShMiodVAyH7SV9Ht
OOHK81n65CwVzY/k+LbTyLjfogUyGjzh2MDtUS02wAG52TYKTrIUc9GOIhQdZUIg
CW6RsVo0/VoTXxY16LWcmEDlWjSUuDCoCew0CGcsPf/22DEP6xTcWiBvjj5QDhe8
JsjZ1X/p7q0ZmAmhBrgff9prFDPM91ui9YljbKtjYuTy5E7B3ZqwItnM7w5pRD+c
KuM3H6HRDqIELlYv4peS9KYA9mhoeoLHDLgEDZQze/nYpdXj2TSM8ox9s1NEBrUs
QsuM7l1T7GYcYCFyuJgWxWah0xrLJWN/GmxXQLDw6OCMWgGQj7lIxIuNxOfY+ORH
fGpWj8FJClLZ+eHWXAruNTU/0uLnzqPXai1j/kkcAEpotmIUWeTaacyNXgMe1s5k
S9TrO74a48PAd2sHKZdkhorzMmIGIMQJT7MjFomK/MHBSOyomCuND49+OOQhVgQK
XCdIWOXzi4pnFnFVkJmssbkQ005R5oe6slyF5sJoQK8i7T3bkZSrWj1fikdLkOMS
W+M3TdkVDH8UPUNEmpZYttv0XNTCLaHnBIA0205hmJQznLBWegAdVfHoOlYmKCe3
9gGcqQkAIl/sYVwUvneZRdaD/4Bkf+TyB6fn4xq/WMKbHuXXQ5Hfjw47Kx+Vf88C
cISuOS3oQKcAPvkOqz3Zz6I8i0Gw2Jlh/YPU11LCkXjUfXU9NXsK/6A3NTzxFNFz
4H/wwYVWY0rY8Out8l5zg82vE/ZO1+2VeryLLbbJDcz1bbqMl76YcoGSLxfUZ+2B
iUpHKs3j0heHZCx0QSUnTbIhjzYyxQRmpqZtDuxUv1Q3Zt6+IMq452XXHIIlRkqW
0l+I1SxK1CbaSKHOImL6T9X9XvTBLOWUZmvrwwEr3nswAwDJiucV8lym/R6AbbvR
AQe0SelUuIXAQZLzT/1sPKXORidLTgKF3pk1Ve2FN0/YEx3jTz5aZceesf+X02xy
E+FHwPGU+YCJ086yqNefYstlC9hvsNVYNfP+hPnktriqW5J/2QHanqJbxIgIUgzp
Z3kwONegyAe7S6HLm+7bpwlxUgPcqXtQct6ZJtsfZ5xPsjbR3GoisEX+sME+XuJT
BT8Fqemg1qv1d0naLoLjp27Ka8sbNm+rGlRVr12XYze/Srtu4WNUapdDO3WEFWQl
joyyeydDzrrunTIh52sfFr83qCccwdTUc2fWj5L4Tg1DU8GaQjATS5bFDI83nsB1
9k5/kaARySM3VBayHre38Xqi8j3t+50MllDLdgvvVfilbUdH3Y0OpT23aGqXjhbb
BzSUBTo//zvpPjxclNA0j80cKKEpMALzTq0apd7QWD6FQp+Y5kqNcYlm08CS6wH+
LWSUGnHKn42knzzmuuix5boDN0PelzR/+3CSvGbUBOQQUC7+S68p+gj8TM6w56iP
TusKNE3qWc+5Sp4EpSf+AXg0DkKuSPs67tbZac+A7jv8lhGlS7WC07kzXaH1tVqX
MUAi7kNIKqpYHHKwxXwXzhg/sXPwYWVeS4mDpNTv7R2Vrd06GKqjD7smKEmkOWdo
SF0+Cx54GmLIB7So8h5+5FSKpI9vze9e3raNdkal3SvVXNQ3BthAk9h4xGqarJIh
/lGlMsauiYsVQOPaZRbWfG3kiK7x32m2FK7+1+klkwxhyYnzHOd0iNxmRkRwqiKo
HXo4VAMLKzDjka2xx9oW1t1rT6IfeuKgnZ1sDrtio0XDTpmoT/1jFOA2kCaPUK+n
50W1t4vveNfeRUbh5CnXjSBbVl2OiAlP2ZVBTFlIPXlE1wozAgUP+1ZrMB+YZpOa
6EIQE9/0HuwdP+qWuuE2JCaqrDoThyATtjexq7vT3ZkvuO7Gxk8xParA1nn9pY2G
HJwrCQzByG/BKsy5GawV7QRxCT6zBmLzWWZ8r/CuECd9NPLNh+xBB4eJRestEv1V
3GFDNhQJ3gt3mKLwf/Hr+8wt24gJX67W48BJpcslQvzOE+EhJIJUPgeGUK2Uf/k3
qOqixAytrZxDIhkdqtPxic5TgvTPGTzvhm9xYr1wQCq2yXuuWEfF29iAfRix8wD9
JPopj/OhB6aAL0KnMhOkjdmW1u5NyRfFQQwZfZ+3/5MmCJXVCeC2n5KTyHY3kyw2
8gPGfgPDCgUpiAcZxCFn984cJtwYDinZI43oooJ7+DUdstTsLEEUWbXVwkdWFCVV
F67eBKLGtPukwV/5Lf38uqo4pr20vO41otHcszUaVinKov0QeNsjah3W7NATI+/W
UvrE8o9UBkIF28v/7tWx32eO4dpHSiybgUmDUeygX2wPx5llsOAYvD4NRbmL5btv
0P+ZiYgbNuR5lOwnC4fYGb1f5ly0pPO4qe0zzeIXusIXMoxVUeVklaNJuHuJ7nz4
MoV6mia5coCUllWNW9YOvSnWPvBcn4I81fLmyIBtrI5rV157EKq/6LHMhAWUg3Ol
BUGCVSu/zDTwvtdPdNo34NJ0RfvS6DJeeZe8sw2mufyItkGo1oaKkHhwoneDgdhg
oDER/eJ79DFOoRyFruD811HffBqlC+STIIXMz3Z8jakQh8pA9CHY9vwifMo7ilDP
vYSeom3LhCZ4TMh0UTjpEqIVAuqbF1dux0D2LIOCA9lJf5r3wegeBE8ns8vOEsjG
ot/3buD3nHk40bCLqs7VK/9SEhlA12thSSNkrIcbIZb+qyN2ctxmeF9E3DOHmCa8
uL5///vdj2cnqeVHrQHR3y27y+rSNYfY4T0cZiNyqlkNf6A8kLnLs3ha6sVz6NP/
tilDLSg+yjsa9XkCJSbeNXHCsfzqeAQw2LeHsXrIEQwEVrOkPzcIOQ+8kW1BUc6n
NSUSZk5g+5VX98qa86rRXaMvww9474aoQZ2rt/wazibgv8xn/9qxZYEHfTUheosf
QBK9GnW6PjjchyJJMEDeymW5EN2AEQDygTk/ZvDe0pjNrR5uC91bZvl5UjJHWRlQ
6lP5acCxR+5CyBXlfo4VaVFj5rum7Fc1Iwt1+yvGZeEJm+ji5jrV2rxpBtA5iX3l
qbfxeU7NCWJlgNvKZ+kr4MYfLXja0VXrr0BBaK/KVKTZJRPpnMkZwOj3i98QYQrZ
beyV1auSQkU7Izr2tyBagDS/VUkfWaCmOEVKmqVKgDGM0/Ud2oUzgl2PCMVClEEu
TvVI1BwPNLF63AdgWqarTaGOnukcd7u7aL0O2M8opKSCoaqgNvuu8QNWD3Ux1/hE
ptppRHjM0zMfDd5/1A0TaJXfCym5aNECygsXZI80GAmugOwb1ZTQ1uejtF6Bu7du
x7dLF/cOoIBghtepbXaLJ7oUDhRePPZUlfItiOf68FUxzY/DXMktQDfB84WEAVRf
6PQWt1FRrCS3pHSEPVfn+enCirEYmSvPyF4MHUOqT6YL9kaG+qCohvjLLWhyCmBY
Jj1/xLfa1e8OfAzlXUFPztus8wZNZoaZQBnXrelATz+YhZ8DAkdrqfNfTYbJOs5X
YUON8hI//ueLmuQ7vQzCSTRUA+HqrCIzyvdNGP6a/3lOi49Ooh7bEWJakcoLehJF
Mf5Ys2KDX96TSusPkQCiTF21ZfCQC/gnw3cI6c1w/Ay0fM02lRuBVRsC+J39abrZ
LEHhE1LP5nBSibczVTF62OoY4JqGIVJckbKxTPw3X2ab3a11uUdedCrvnZDZ6RAt
l3r8LwRMirXMR3mKp8F9XCUzlRVYO1XaEEqHkqg/hmZghJO32QZTFli2WqK/o73Q
Dpe78P692SJY56HXdZ0ThxphW4Gs6sZi/Hz+lOUlH1qhoPRa3k9+NHwFbfj0lbLg
jSO6RLImotyCFHiFtjpS5MBU+9ImYgkfnW8zptaEftdOr7mv/lQUirGWkxk3R5RE
NcID56vWZjeeL4BOM/wZK4nIRcAMyuDwPL/9d9agQ2rVvDjVOdkc+vtYPgq60v+Q
/O9LsiekTidVkvT/so8hMxz2RgH70oMWt29ZhcD6phX6uBIpIODSErTkks/hKGgW
2SRRMbMP2ESWVzGLUbatoEGTjpf5WSAso5zv0qtQbpJKTrCVQlR7o6UXK1e5WR06
WEuJsV9VSMROTWDKvsCk6GiMUb2dbkMNqnpD4UR0Hub4Ul7cjfyFqoo3o4bO4PX3
1t64l03YrA2WpiVmKnF1XcpWsQyj+CnRG/xkxDn6l8SuahvAHfZ78R6aY+8dU147
r2/jOYINfIcgVmGBis04NKDK58RC37PWHltiT8BYZ8PVoaX3JPs0sRzL0vR3AVjw
l4uU+E60erAxjfYaUFhjgLBS8u1uHzoArA43F9NBPU6odeykIhA9dsf35qk5bSNF
wistpp+cUqvvNG7JLz1aKWyguIo+dPMOytEGAqBn0sfhcMnSm+UYpuEq9LarSyWk
ZAFwrXnQMHIruOKb6uAI8gOkWq9sosTR9gN1xBiEVLI2BmpAeeJEfO5fJDEohNpe
dQQIPrheKa7PKGOzQTuUOexSk+QDmOcuPQYZeoCy9KP3BS8yaxUMjNKBSitDGw6j
7Ug62BkfhKQrrgiq0kxeq9zH4P/svc2Sc2vx4oPHGHl8h6PCJLGAWgbQdeXxiJ4g
aVeeVwk9t0tR0DsBgEbGoJ8sEeA5VHFkof80Pa3K4zBMJ24//rdDI0mVyqWR6Mwv
azD6H4OKyfWgnME0QXsCMTagVDl5UGtuACLn9FdivBzt3d+p6XJSniZOUp/VxkE5
+fHDUjABdU6931r3VvIchwqCylVOvfrgpjZMr5YtJ3fUFH7n4vpe0Qy5QZrn0VJH
OPI6ybabUjC67oJy1DslMc+vGTyIS+t+RYsyAl401Hm0k29HJ4m1n4bypzEtbT9l
1Kn4LH5hjmvZLmvmpcmslSv2Wuf2myNFvJtpbjSLMVbtt98VNpvjEM2DlHZy6AOU
1SMpAcMCfzbxdX1Xvr0xw1fOc6uNOfY1duMlvRKkAoYVmkFm98PUHigJq/v+YZB+
TyKizqGH55WUCqnGKmbhG/B+t2IQTM0MtKA2qeikpCrTWA2y9IF2HrOlERuZkhT5
91ySWi8OBval+gvqFGcACDUzbHelUY/p+yNiflqjKYtcsodk2yp71J8pq/5mjM5V
9OPeOkxztPJwOWrjAY2lrwYYCUoVyR3wJkaJHxUHqFyhmNohh8eUmy7b490MH7+D
/tQZKrMtOh4wjLG63LnAeDkAqzc2+bSeRqxAqb4T3QbH31JN+ajKEzEKDcCptSze
6e1W7d1RVdiOqYVM8fJSoUYMMnNSmPbzmyVHpDYBCVgVH2k0sPxepntAbB/Rc44B
4ba2EPG3rAvT+U7vsLzl+MXZXtv1iMKISffbGiwk3FWeUP2gJpuTFmTzz4UILP3Z
p+BT19fLKm6vjPnpMMUpogFcenOx2ZnBw7BUBo5MGOIIr3NAIaS24RvU3vPoZpRW
u4aRIfEaZyh2zzAk4VXpk+ZXTC37moO1AAtnBnocdpoihNJmYSzRDoEP8mUMWDcH
7rPTllhTUPosfboOyNOnrWTP3xvfE0NcuV2YNY7IBCATmtMg7CbpGINJSIEggn3H
umGbhrGHhG2NIuyKo6JNYrsobqgiKfA7iPXb5nszmTBR576XqHi6hV3umcqQSZtu
sZllRpHsl5FUTBtkP27ncCAcx0SW8mUrKX6w9n59xDIE0jB6umVcUGDSQfMQ4XYM
UOAtwXongRewhb+46PIaZCFWbaXrq9kVJEjb2LMWm4qdF7Ovll2cp+nQtSZ7xL/w
FvEBeJLsHHKdhGzvIhniB8W70gxZSvH6mHP3PprsRj8/TGFLuXOtIMgl6gMnUJXD
V5uSzOsu8Q6jEJbJZhh45mPysEUYexeaH3jtNLi0GG3gh8m/JgML8n+Uo4yTKGEX
epuK8u7SIC5IBKUFgYmqD0njNkM7qW9vINpoWlmCxUxPGHv+0thXrkdw98ipqNLs
AMe3Lojg68HCiKGSdOOV162cKA3NybPZMy61tDwbqoUoICADXH+0hfAFQmwX6fNf
RYs2Lz7kSLphTUdtavY5klVXW8xg1fbBH4nNqnrkvt2xtIIBeaRbL+hbVUKpA0T4
h4kHAAVl6m1jYee3dg6L3byzn0SW0F6hXouNtvyZJ0NmZqebaSkcmzhWy1/a5jIx
Fe/xxVU8ZaESw3PG4oak5KPn5x4j2bPGkVEJO1t8ofwZ1axr/Vn/WNPMrCdajJKG
wIq55c2KHKBXNTRrHsC28VuQlbxXFsddRSisS8njWvmlFY5O+2kbduuXOY1c9ir5
wb4R7LIOa51YtKrVVzUqhjYH7H8pFLsHVuNHnSYGlLTLx2hZhzTCDPm+I4ECGSZb
bspn8oXQYeSnqKbX/MVJZa8UVFm6hdsi4QkyntiCI33XrZjS5UAfWzADxIVOg+nV
o0ORohY8tib3uO9WsaWTbHMAItRoE/jTW9Ox9v41PkWm95o5CV2p/A8WyhkxNzpV
DhpAaCmE6vYpv7mi0UTLhk8d31TL6SSewcaNgIjUgpBC8/48x7hUEI21RKDBAGuC
teerrZokejqKerzmgocQy4moY9sm3/X9ayh4CIwB8MoyjRzn9Y9l5oUaOV39CGyq
N4ZXjeW9DYIaRPbcZ5VKCvIQO/CyqP0FQA9lgl73A4BfwhUaM7C1VNbS9dTguB1p
CZpkvVuUTUiCJ0RMPbjPssnHby9wOn1fj4T8yOUyDVej7kYwu1XI0v1jt7bi8riK
Gv5+YjjHh0iwQph1JmkN/L3bovnbUqSFNYiWi6laGMCYpNC6n9SsjSVF45PGvGir
HJcBertIDxC+/6E5jKry262UbJ2ALCfX3o2RIw42wFoF71m2upnViPAGdLPT4U1/
l6L2+sQB/wWbDxzCGApaoqJsUlESpGqsvPxT6PbMuZvfZiFN394rwV0MTmEH7Qh4
8B2GSRvOpgF2abDyM20JznQEvs3OmxNZiR/0uVi8g1Wb4NdBpfVG/bzk/jolWN6Q
aittmvFj4fn4Z33WDpPKnn4fADoLVOSopXir+tKQwD8sbXUZFJwvXJmn172k0ll5
2G/Fq0ZHwZ4x+N4hS31V9g8xa7AzpkoORVQgFuDTTqMzWHEpm1GMyEylbNrWE67A
O7myzXeXFdzi1FczmbxpUZzHka749IZ5kZ4Wvi3IgFOWn6VjhpSRC26EYXwt48Os
Qm51IXFv8PuORssuqXCLzuxBq8XINtxqMyWT2FZWyGHdzwpdJPG8oWVsnXutdzng
w+PenRyy0cLB4dfZac8Hza7UqlJKaR+hH+LSTPitsIvHi8nwkINZGaMFn97wIP89
JY4pDR0qpg7bPhfayN3Ia7U7BZ2mD3LMAzPD820NB88MukegXq59fNhspK7kk57i
4xohG9Vqfz1uv3Q0PLsP/P+usO0LatczrQz3OYNbCyCN8LBvy8egsDGH9hUquE1r
0Skid+S62fVeOa/DvHBi+/+bH0s4vl48X82rHjHrbSlqAnBeesq3G3x0t8kres7H
kvvH2Va6B0vb2tp1vaUgzV2o/9OFCCtMkli6xEb4OX++jeS7TatwuZaZfS7tKmlz
mgZ+gnU3YEP3KZlobz1T6unWSRDh34+OmbrA4MDlonDBnPxQOHcKzn1jgptWJYnG
4zJhUmDFPvCz2RY4WduYHs8S6MuCKM8EYwpRAiyGW4Zn3lTF6F5QSNL7H7JgU2CJ
BJ+ZJen/rsS3tMq9vJp+5fJ9/VVFel7u0U7+zD2P+u2+j+dv97g9UFJCWbEMLu1v
tb+ykDLG/dL2+aBWADT7FQgNb+9/QNcHVlJDAMtKFOXa0ayu6IohojYMQukk2zqD
Eyhvn2ywg3nLcU0dmr4DRdgJ0SnfJvm92ilUFudokvnRGNiBBhZKm7IAXvEBQ5Ws
eiTHDuY/PceRaDvjUAZ+/Nl1wO0tI7+WSuOGKdN06c1hJopVniKGtUxwQc4vex/o
7Gj/PtP+tIRcPlYj/z4vmsO9TC6A76/NebuzF7F2yQj/jiA51r351qu5tzkzkHwC
ZTGtLPbVyBMJUdzpLJ9Mf+F6bnKFz5LV9PR6heLZ/ctz4YmDS+e4gZRL/iAaUgmh
ku196Kb2vzvyXUrv1XXrxk8h2inIvybzu+taVnGwvgw05A+nqlblq+tXsGy2YXoa
ozq5U3zZW69ZKY5urzrV/9tiZiZj8oZwzrenIlGLZ7s+4B4b/dNz4V4bwH3EggyJ
w2b/eqRvSmAeeaQbgiCIq3i+iNAaC0QxWYwq/LItIzWwWhed4YKPwO90bxMSt4Ga
8nfKYeR029uZbgHy09J61+/Juj9WIl+cmg0hnEOtpBtcJrWkADERXYLabVieDelH
epXx6qL/JaSurDQwps/3iF5LhvP9AFONcuEQgqLDFcMml2vMKxVM+5DNYrKFtoWL
g7XwI+UuimWpuRDVVGFPq2hx8Mqrb6Do++u730KOg7cmShngnvlVl9vaTfYs+hE2
EYK8lLmVC6e2/W/K2rZvkBoNCV2W8X3F6OYeF59TMCctGIsCCEdjDE3cdA3CwoP6
1I+KhLEWzGzeeqwEGGzbBW9XTglaU6iXs1CgxIXL8mNX3FzXZ8+yEl9UEeUSvLKM
ZzlDbQLWgGFe/6IsHYWCHKCOsb2ThuD8C5dkdYePIO6fq2nb4+vqNsGRWkcvt1cR
OmefF0W9XDs4yuJViF8VSidR8bzWXjAF0zwDS1h81w+Imsk69KIzgaGLCzOczJ+W
S0BjRN5Uc49/cU/4687Kd5QWEEwi9t5dtf5fbmkF93IrXMQDv4hZpYBQ0yb8XbNp
InUpSBiC6SPy6jNc/E28Xed43dt3T48tKdiTkQIi3anesTiStuiwKLrOgnmzkM63
2QnPPHVSRQxZlaYH/X6bdsbxgc6AYueicMS3JRC9iVBSRNOSWZd2rYKaa/9F22O1
ZiEbJvbqBDzSAhTcEur51vlDCf/YVxO3JFevUN2yVjuuQOtDvi09NDe5wOTv2gI3
3Eqf1kc1ufO5HQEQKivemYrmVrCUVCjNQdLJHMCHpXg4NKdqESBsf1fo+odNNA5v
/+YeDYPxjaTstDA7GrCdbYrYpUlL9fmV+ij20q/50AgvmfmYwWkRGXfMAzJpxx1t
kP/mnT1yHRDPurTUcGSGtO8HMgcHNgry0LTRmC9iQG9w4fIOxQymBeU1mO5tieOY
GuoQs2GkoKp5QQa8U0ha76ewcejPL2aVPTD9ulzPcHq47Si36avxGoUVG1WVLv0Q
nwEFyeEEH5OCN+rw37xRdrvn4wISY6UeQZxz6XkGUAUs80qQ5M4BFp1eRCXF2cOO
6ivSm7Sfa8SjVm6I6XdweWaXzsIDoCC9K/x5yJNXKX0wr2jy98/3RvOujO1U9pkf
TBuIuP3eFM0h/8RVZFdyJJORSFdyqtTyu8fC59/Q2mRzWL2/UeDf4yuD1kefWTuE
Q1lVeC74Sbz/6Sc7knZ65e3OTj1H1YEf+hwZH3+6HqAb/MOFPiam6UwAuRjkiuoT
KTezFJVbSFewlXPepJLuwMkdkCuRCiohkJynNAFLdsD6mDRcC22UvbiOC7wL18B/
KJTg8QVVXUVmD3HMMpUd+FoZfRTFJOmqEoqyyStRcn175fcJpDv453R/I72+COYE
ohEJgNnlQjiN4ANocMHeytybvBW6dowlsctIIfC/XTqMOG0uvT9x66en9eJV/vXv
rAd34A3keNjO2DmGa69IOqNkAb70D0UyTzhKw6kZkf/Z4/KjigrjAPK7wo4/PAYT
GylgBcKe95KbtBVl/8l2HVwmtX37L36GFJbpom9GMwuRqI3+hTA3QKEcpvNhfFhs
TvBdbtsvSvRFzNIokMIIQ+lBW72nA0Z7C5y+jsMb4iBXpOmeDuCzG3OXcnuu1s49
raSsVQo+qhS1ER3RcB52huMr1SQ72aU4RUWNgI0Stnv+UVMYExV980gW78+jlTaf
5R7VgRYfEDbD++xNecJE2qSXOPSj2LDdnxUCtEaqUX3zMGKcbXHw9rMRjyMNiBqf
iEEgyKSzhnRXRj6DyHXvOR0IMxz1vj7ZXcHSB4Weu7m8XQ8ssp7XNsSiHoysxaFH
tNICrgHiRXEsHQfINCv/EyktM4dvioPaybXA/hYn5IlN+OTAF0mlcE7hP+XSFKXf
ng/V5HH3fL3Hu2lBEdo2o+hQYHXzNtOCo3KX9OK1aCv7U7RVHITsk5uZWXXjEZwI
2HhSICJas1AteExM2WHY6wv8wIgX914zu+oRnYWfM5wHyPp2ZZgfSsskgmqpxvfk
ld4oZlTHGkZIG6xW2maQXGBmfQ4rhWLT7R6oJeEO2wpeoq75y3eaqzSHVqpvKGdq
wwAZ1CZGfYhe3kxg+UMo1uillM06Z6fvJTbgNjOfU4VXgwqniZsoi56n/KljIflO
dLPJgGK4gBjEU8s1M3vKbJT1Qr2mdk+MLzitb9R918TfGPpgE4pFn5+vPYpmEOTP
UZbLf0DvXFCWVS3Z7JnVHqfWVbUsp96IiSgJ9yH2ocucD7KYn69kXL6QvGZ7ziZh
LTOOW6NX8AdDeDUR3tBTbxn5+Gu68SpsHUY0Wmt4cH4pH5XVyxTuzLeo+X1JUWOE
GzPZq0hx5sriWe6B5QJKTYtO37ZkzGMZ2p2K2awZgTSMqSUVO3aNg1HHRfUs+69D
lUsTtw3AUryEW1eLKal5oAGKPdewhxL8sB4bkSQyU70S+0wf6imJXS+pO5yTcNyk
M6PZ5gCq7UOQJTqs0//6XXbYjjO2pGX85/tGENNPAeE3lC91sEFp29bmiTqn9R2G
i+cMpFPcgpNvl3FL6RACwjUQMvrv5L6hbNVO7Ff/lhXHIwZq3QjILZIcle59Dg/N
I9oYR+ouxo4u1HcgRKfiVuv4hqXwjtcvYv3BUpAWC2cbMYcMnygMv8LDXiHqz44Y
2OfIcXMM+luqYYu/exfkojTThxf6Gpn+VtH3+g46QTgywjzt+Tu5yVBxlmqiDpHW
wVRG04Pt3cqH3+LJdZIqPcq4AN86bdc9wxYHgu+tX8rqM+Twq1h6yI5cz1/yCyyN
mYpE4PPCyMUFxjU+HbyvMEph40XrB2Su9v3Xb82XVhcvT8IS8kbR3uzMHIMWDJzQ
ImEhj/5iG0IuexlBFcs/rpENPJvEG90DXYy76MUhlsJhXkz0zzpXy6QHEJUd+21b
JR8o8pFAo7N7CliH1fMgztGgup8uh6cpMWb7lRA+j6vFe5GMvvJBDn4KjcrqAbwx
89Ex+fwoOfH89s4KUxSjFbSdQX8bVmVx2Tt6vICE+a3qAYgWO4vSDjGznd3lXIdR
J+Op+Rse3tIybrWzzFV3YKw26gSFy5Yn3lfFC+KfnErdXbaZqZAyf/1NGWmftdSt
EcQ5cgm0PMYQpCLQPNPF4nDxvpH1oc7fvUoMQglBX8LU+AwJ+i+aLLbak3GB6wBO
PTJfGkOlRl4QE+6MNPvcJcH0RAYGxVqDzqL2wEz+Dr9m+kYN+8RRl13UEwEn22x3
kX31o+dwHM5z688qAbljv1FiY0AgtrwpTo+RKD85CVARV2aJ546uI+nzi+ogar4j
cDLBpot1jE/amfz36WqPkCwy9VuZf/TvELJtFzhmRrSvL0mIuw/XsKuL/7nPZHxf
hk0rASU8AdWxi1HvZsSpVVe3rzPpR/K/fcyw18bfKBaUVudEHXjuUAG63e69HmBb
K/W1/QjG48mLb8I/AUTuPaiqT6TjbOTiNghCIiMoG7DgPIzS2N5l8cdlmNjTQGFA
MwnpgeOtqDqlnCYzZXfPEQjtXx/Hzmk7Ku3xjQ0lw5wgnqMjVjdazXdgofryPUSX
A/G5Eze1d6yD36XDzdEw/7R9eAm4ZkuxsuMf7DqHveuoFlMD4jFj38mysSag97hv
hFk+0lC2rrR7PjkAfg/S3QJ/rySq5qvLWbEEDppIOZvRtZO/R+GYCqfZiUd6TUV+
J18KmyT/hhLDQDCiZqOwtlzjgoRQT1SjA4VyVBcFmmkx6GhpnMdq1W9Pka8AJaOv
ZEpJ4cDL+6Fj8hw6IQSM4gxP/mgBNc4bz4T56WHwVfnP9PeY/vtYgYInNqLauHhI
UmNT/EijOFYeP48X0/UOP5YYSPcUBNICSrxXVdZPOS4uhqvE5/PMWPyNOazFv77Z
OI29RljdeO/g4NyJx9T7XpCxc0HaoK3KMk4zQ72eaaMH6YBS8VbSmeWhkMhu1RA6
sTjdujkb6BY++h83G7HAZrrufQv7ONqD8q3S1/yIN0Eig0Hu5h/cp2haTPYZqwQz
OS3U4rNCMjvA+MzzJ+9Xu0VrG+fzhkix7BI1fEFL5NwefQbdFyViKLiyZDkT20cY
9VlMI4JJdJgvjDW+qoDt2c3fzIL+PC9NiqZWit2PawmqDPF9sqEDedrAS9cZJNqX
oEIW6kbOORVDbYIVtf7Q8gV436/7tRbFRmWBhtXpv0pP8BTjlAOtjN+JMc9IMohl
I7dgl4LqpERj6zy+8nIIshjLbArhZsFYMMex6RisGRNtpJV5FWSdM0AuKlxMwqXN
ynKoSU9fBKUBMKn7pr9L9KAfGCJX3a9mZ1Pn+NOdmeqJpOtDc+lvd8ohxItus6lD
98nwbh0ut2Zd73gaQbfpLc7XlXtRqcaZpbD5J5JqocK0kYGETKaLlbBVAojG6jee
HEPL3/3GM0UQKG2XdksUvdjzj9acIcjpLqUpRal/l6OwTF9Y1n7DYJP61y7UO6Fb
4A6FatlXvP7s1ULxZQ2J0r16MHPnJJAeDbCWJefY1yLV37luRvzwSjatmJSJN+Bj
OEUAUw2S4yuQH2OiV1YFIR0bLim2c8hdUKgYY/cAS1Z0XtQ2wkKk4WbGAnMVtf8o
THsdwmYFffNOg7sgdrcpgp43zOCNelgXYtBNZJ1fTd+p1u2e5rH0ETLz7uj7oNNH
UBNxORMAm3hO0RjLVp0dpixksEg79RAf1YR0mT94vGSuOBe+oZjs5cm+SacA62bS
XcCZE9AUKN537I9R1Hr5f9kq4iNyuFEpTKmrGBKcRAGM0IgxL8pa2VLQutuRLXle
I31VA4Wum5B4nb8OrquMtBMj9KJuUt3blsIYwzXSZaRJKzDnXRDqz/2xUsCC8tFE
aRABfaqHBbWHi79pAk2C7K7wxBl8BXVEPGwVS9bNEdhenJ/QWY5eLce95y2xoNW0
jAIIh7mRZEOw56geBCjtM/+Zymrl4r3x/Lyz6Xy8b+gGhNh/9utIljxdKcQrrF4V
mtQLjDEHoa+lJwalytwdLN2HJC5ocvVdgQEm7MMbqbnXfHw+xqVYXC3pEslop5AE
yabuUDvmV02i6tGWHRuIEpY7y+lQZFmJoNk9TUGp8TJJO0tehtfg/E9mX0QtfPra
r5bvHOqUqCle3hL5qnpEVUuolj8Hh0dQoOoYmJWpc8MbbfmpDxtpLj1K25oCoqo2
Oj8yvWFTXoMKNtD84YfQ5Kz68WvD7et7i7d59auVyvJeC8aW5NQpC5Bm05VB5qXg
5WwIzDu0mDwBnR1Cn7WwTwq4dQZpXWYBJtxCy84hB0jCQlIFuy5EfxJkE69CXaSq
BfU735ZG/AHBMHCVZo4cYlu4Pvls+taSvnKeIi+qeCvmwVQPfcLOV/PkH90dv3yi
7ooyrpBIeW8r7+DJFAS2x+M47bps+M4z2qOrZCNDMQapNvQHEyLawuYRPXLalHP5
VAnNuDZKNNilvQ1CATK2Et8AwzD4AiD8JFNSs4MJ+7s026nuRGKBKWmmJKZJebbM
bsrlhi+vmwYOi/L+uqMNV5V6yB5byfZZNVjFWNq5/JuL524p/pHCNwHwb4dzzvEK
RqH/YwZr5Z9J/qwP2WidfMMUmjMqxsTZZq07i2C7c/bM3bgkCTT36Ym3h0Kq30Qp
2pEwvsc8MG/GmrYwEGq9FeLgy81+l/iPeSiVu1LF4k99XGEWV+yDczd8NRmxAQKA
3Q+xcPin+e/dHjJSiqkSAsbnOgXPIkWnxluUw4QxYYUFxD+xw97jJFHvmZD9lT3q
RZjcSPnILF7IUUfvmd48vv6aoY+cSCE5brhn7QcNq973akLPw77FzemPOcM5o2Eg
1syyJ/oZfsxg/OLXGlOUKoxjklFiY26N5He38DzogygALCSX+rgyK4/aKUq6oAUX
K3fiRdKxkWo32i+p22EDulOUQ6GZOErEqnlGabZjxyduI1bRHQ+0gAAcnpRi4QrD
gXYRAv0aUBNYjMse8vKqjQvuq4EzhZBjM16ddRlMiO1aJLWhfV0j+PBfh2dei5gF
z1oLGdO987axY9iyeO2FJzCYJA0k6xuo3tjViMrGqZNrHRk9ZXeyNzA30+Q4MxU+
j5Yoov8mbp6JtGxFwHLB2Ap2/1VIRY8kye8FsTjeZG22/JsMfMbNXJVZjMCoGkp5
o+YSwHjz2MEdb37IBZZnTPwsOGe7E8A6Zfac6iuTu2ZSESl/Lp8bR24UUWXGyIgw
GVwwIP5DI+evBpvUgd/YKpinjdp+phreuyrP8wS6oecIdbHqnemvJRgcZ4RJqQK7
RuML7LYpsXsGSwdLfwgQAyWymJ5/Ax8Q2u89iwfXqURm69Mm+k4yJSysi67+ncQI
CKDfcDfvsphACGsDo5cVzgj+XcDTP4OCd90QmRgJEXAkICDo1n4yWzYgNmYznPza
NKvPUYElqVosM4yBTXp8yAL1gyGkyXkYNQfroH1k8ROhcJt5+osu41Rgg8PwJot/
z+qIqxEpnidsaIapYzjC7KFywlq7Tn5mGGUWG2WdhhnLp4A/Tt5sUI1tmCuxs3Gs
oV/U6wkTPe+8sf6Zzrema6fYcU2RDZFoWS765Bqzao32dY2PaJFnS6/agP+1OYuv
7pEwKZv/QANtZOAMtYHrfooBAPmFY+YcP8JJzXraW6dN9EcjdPhh0XwOdLUNbtvw
7YMQ22B59OB6Z7sGEHONU2eb62tnfz11MbyjSI+46dtFGult7XVOPRf426+g7pEk
y1FJB+w44zIFCE6IA3kiQeocaJii1TxEzDtxntAe1BZoSK5lv092Fhpn570pzr1E
ejZIy/NLi3vAFiE/Ejxx+UHEBHyXg8OMCZBPd/KiOAHuq7hOoXUBt0kw/SDknzNV
GOibUPAz1AgNw526zJFMW92nD54dItHbWkZF2hJu6a/GKdIY/B+DeYjr6sL2murI
KhT/jURLeMP0FCKgSZo5Ij8zOZfVb1HN42ciNqKa5k6CCQPT6Pxf0DHQ/MiAJ5Db
Nr9UpQooUz32IukhCS4cFTQCB51CtZuO7tvc9aKHf0zP3H92wFIGtcBzTEYWXFPt
uKK8t6o724t/AokOCB61btg8TlOasuNrEtlDqvB2mPnCBEDUA10YdGzbcMJe1tLc
l26aRxnib7W283JqKVTOqhBBvs+lGhtOisj6SziXGf9oTcGhqyQgKtZlirmfOEe/
nLc5V+235LOwg9vaLaXcWaO3Crsz/ncuUK6mrfJzJkKtxoEOTHBENjdQvDb+AkF4
caRYh4vdiBhJG2rwEHgHjampSwF2KjHTPVayVEgj0+1BJiMB0cDlfeokhJLJ7wp5
urlsHxD1l1CQ0bcyxG9gCiCkYevxONEpUJq36B5BNl8IxHZK/wm4c7MvSdBSVXrn
lLIofmmL/P7UbbOBtxW8kdmKH6jWb/jexskNeRuAqug5vPBCsLdY1ow3rgONmwmi
jEWvBaKcTwUPw4T69+ltccK1SCCnzDp8EwyIKArMKEFR1hDXKSbRlkE0wgCGMnzx
O5jD/PfGz16WcNXFm13S+epaPXAHQ446sq//seyXXZjigVEP/XDvDawr4CrwJqnj
T0Lua+VvOqbi9h5DYs4Avqkg8KJPnJCOJvo28+7pfXcmJcHZYy5p8ecN6QDjYivz
jlwHr6rJPkaDzcgvddiG2QPBdBC71jBQrDRBq/MwhLkuwo5ijGBByq7eZl3fW9j0
7rWV5qkf3a7ReLadswixZKQd5m7nBpywWPfb9sHwoHf30QNJBTa/IO9B+TU351uH
lEzRnajLsOKuEiD0SMdKc1dyTtdatSz9aAZ8H6NPu7oSIBoq/zN2y0CGCYVnd4mZ
uvpwLwcnKmkzP+3AeTHXkV40Odaeqoagh8Mwyb10aBEv+S3Q8jDmWgscM95hSElA
FkNmfb1uQVq4uLN0uUtyNs/KpWAYR98Bqv+htpWY9EctZiFKZceZqxropZ1A0/gy
aA4idM4PLRpK9GR8+KJYwTC4wBreq2gFQ/JdTGYDkn5G74hf1OIdZgFHwBN9cmzT
4lNCb5bHv7HNBbY0l+VBzO1k6WgnuxZaIcA2ik6tDWz1scQ5OE9XOXYA8+wbcfRe
/4ig5RHylLaeKVE1h4wWYxP2PVmxVTTnM1+cy4othHHg2Q1xlZzP9WyC3xD7dK2h
tCCayaueMgapFKKcmuPuBV/WqVbvBd44G6/pudCWB6dmInF/nRBO7PEEIDurH7D3
1UBqbpO7dptc0YKqlhzz4ObonPWpSX19LQAEGP3Dgq4mECHyblsVppgr8vcvYeO4
1M0KUiWUt4hLCYH2FmalpaRzvix08DquHR6eojtjc4Hx4qU60/3vQbeDUTUiZU3Z
Nuyc4krX2dI64cEQwNAA6b6zvIgnFiCoqf4t74ujKc5EeRjOzl2oTui2dRvvHyCM
K/cyu0ce9w2zSeDxnMKu0gIcbQ263CdRPhMu79qZLQ2sxX4RSs6RgZJQkZ5HrB/v
c7AhRiNs8WfLctHG5X47YcUk5alNOwnoRSilIjubPtjYvh7IlopR3QPjz+9wY8nl
nHoNN87dPb1Sr3ph5dQQfXlJsSpurcrQjP50ukJMquDDP8b4dZJ7UOPDHNRNrPA3
kA39hSIlQKucX4Aw5YJ4S8aHEvSaQzrelsHcyhsKdbbmegjq7j/rqJZAi/CWjZ8v
9NnnhSo5EAwPYnGPl0/Crl2yyzHHojSNzN+EKKSzy2gRV1HIpoYy2qPCSN0kSL9d
8tDNOjiowEkemWDglk70seSRQ5ylHdNv6zZHYaHj3sxE0jS6s9bcf3xzUaCJB2tE
Xu3z5cotnikb50wM0LEqS3UFntLw/F2m6sruejLLnLX6z3jlpOSUUUAFM8mowBbh
awb2tARF6qGgHsYkR2rxCNjNEmoGNzAHmgVQbAoetDS6aagRaABiAUTaPVlHpSpt
jzlaZcqVt6+qzLefE087+XgfVcNE6GeYwsNeFDwEyWpSHC5r+irtZTCH/FxLbGIE
QHGZeUQ7aVCaC13oo6YVF+f3t8Z3lIoLA1lDqjI66nqSz6A1MDsly6HDBQWf6nBo
9riuPGr425CPSf18iRRDsgJ3Qo2C7nCyJyUNMkqiafjHNjYpfIYTPAi9KCPWpsbQ
VnSQsYChd2gPau2qz0as0xiv2oW1U7nJZhHOWLW/O94H/R+COlpnKryDBfT5cQJu
yhkTBvsI6mbP59hHlu3BZ3vukqO0Khz2NhQousOFrLIg4xOTA33iHiys74WxPS7g
m1vB3mEvFSJAYwVk01hJ+sxpm9xfUwqR/EeWvQRrL4+wL0coEzZIsUzavAFCV8TS
0+NSZpGpEru1ztEKWx7okh6Zm/8t7jdpnpMrEI6E8BmS99oGAiCsZxcugQxfb1DQ
HqsgWCt48a+JJnDGiu5NXtYdV40OV8RzGnH0WyILKvqVqiAjemOM7qyUc8nR7pZF
qICGm7Nt50Hv+tFcx17/dYmElTxlFYRYpLHJLBQ8KfqHMPw6/NmJvK2bgVec+BEd
2doAREzTyBPOyzodA4JuP2Xm/2V1behg7/vynCRCrxla+OO4n5eoMSvLSAjMWkmG
/K2+q+ivJWRqRY54uzyq6Qx79tOQAV87dfauyNjDrF2dDWiCiIDJKi+NccMwatdT
jrgkRfAXQgpxM9qoO4SBTCMHHomSmTFhCumps+bDnHi8iDL42YDc1Q+u1L/eRZxh
ex4K8DbyEBl7ZmiuuPtgcZrTLinuX47xuIQKKxVuDDMmwSkJrDemWXFRxp/HIFZQ
hx2NFNsu2skZj7Erf3gSd5abJaPAkUOlXdvCeoNiCAC6C5xP+J3DHyDG8bzYXZp6
WruUAgKOoKtKApR8ufM6wZYDiPHSqMsJATtsFh4vjvY4iFu8ylHL1w8vHdz68G2q
Ss5iMv3aqZxxA5pamN1TVwvysqqPlKJpRLSDROZchsW2/CsbeffkBpJHyegf0yyG
ZNq+bIwGnx3+Pp2FBlnp2E8N2ewzeKC0/vwdyGekPHOn0WVFaS0yV1ww0dtD7ETz
rjtuL6naCA32lN2UHW+kXv1SUBavIiGL7htfEB+Z8otp/1jXaDebyAVyPwdW5g3u
INzTmEpmgIjrlemREGdp6BJqLN8n5dv1ls0iKduenWIhM8rNAqSfZua7VhjP/eUu
bb9bIsN4GVOMa2rJCvtIgbQEl2S2vEm2Y2hhr12tHWgPz1IGioDJ8AoglzMx3TDo
mLUudg2KLXq8C2cxO3tgB7RcrKJW5JM2kcvT7rXtEjWamox/WxCs9MvfC330MjSS
ikx9YBHxb7pwiVRN1FHluY2tjXhYywGXsKFI+botRgQ32GU47QLMFkBTMJQMKAC2
pyr4t+c38N9dfr/hDY9o2QiOz7ilrRhZ5TgreiqL6EFXmTnFB0SHmEPZ7W9zCsn0
vKNB6KYu+hRyGkOFUT78EzgKJNMxF8xGPJ7SiXIFty1aBvXtxZdGzed8/fSatJWO
rjwTG/5rS8ifzXAZ1Thx787ZGySWBnANwCsUTccyFq0GJq0oRsqHQVAVGmtmSQ2q
69nqnt65stZyhTqcn8vc5LdVNBEja5/sk4g44OzFJZvsMWYCWzWAyoi+6jRaLXhV
FbCYccnn2czaiVslkKD8kQpK+bTXdyJKkfSaYUmwf4tVDE82C7MN/n4Cs7kAK450
Z/xHxjk1YjX29DjdHlij7qG+vRaUFqUn3iDMCDwoj8DKRkLxLWxOeDaVSA85Zhpz
zjzAXWFlml9pQ7zwxSlwCsPS7UnfE2xRG/JcMNSsmrriaiqjBLtL+MGr5r8bk6IQ
g8AVLJgs+yU87mJOBx8X4o05YoA1iaF6ZeZ90TWpDug7kbTkmgVTI2Ue4n2n51l2
nRsIjM2InFJ8AS5KdXOr9o67qXhuPa1wkK+7shjLdqU/ELBOeNIwwP6jaMLgeiMG
M6+LRg87WOwhM3XFsMXv230OlkcurxWXl0/OdUef8nsLcl1KP9a7+NX1bA7xXHPv
7LUZRbGi3etUUOWRC3A+0vuZEuD82t57ZjHs9t7D/155HUTPGvFx9Yn3qIgEPk7P
PXYBg/kX7CQxiHLGy1XA1/UfvTGeGEjtdyTutQcTUeTCTCe9jdffqLO9n9jafv6J
hp8Jh4KhGbYXEuSUM5E76wXJm9/U0zOasWuduYw3B1VM0c9sUXczeNOkAd3jAV6M
iegQVd2c2WglraUPBRzt6CIK5jx02/QURtiH9AFnQtXfq9w24EBAGhx9sfu0oh5J
utM6VOsC8lnbXEcwnX5JXXhREAQKEeObRodL8uy8xoD97tpRS0s02sFVhoi7AtTv
qSn8QV+XMKcAynm7n3TTq3/pPJ1NwN+k2wsBplvwJwcx9gNLKxnPrBSdz9xW2RZB
Ta1CReKKp3s3NzdNgXm0A95oGyI01ZtKkw2v5JXjXXea8WaIu4iBiMQiYGtlMco7
RC4JY3SrvDH51+Xjexb3JzzxRBKMZtWvBbK65VLKIuqIgdRq70jUwrQwg/1dVZj/
J6NgltXMoytsQ2rrImoOsZRASp4ad65M/oK2BTkxTJ+WQVhkt8FAXcrVQj3ByW5n
rV5rEFDt6PPKHKRnfNQzvcoCVAQ0M7XJN21LdsOAzrliO89lq+3JDZWu/kMEchns
VpG03gVmcNlW2pToi4yJFBRcMtF/16WlT7swOh8S0dPWKIw6G6lXE6ok4Kr5vlE4
fuIN6rtcEibuy9oi/ZPD3bRM6dnnrZLUJAgv1uFz68ScR7Hq/IiNP+91MRjQQkKw
HZafNimoZBPBNPRvHOq4iuAD+tv+zqATBBl9ENxdqDd3csRX97HShC67W6MqjbB/
X+1SD5floSlN4KDQ+gxICuaSNkw2/QD0yLHgOzxdAGalwBSkrrcjp5cxNfV7jNv1
L77Ztwq9bbc/MyCD43a2XltHk1ykhcYMMiX3HUWsy1/bc5Y+5ZvjsrTyB0t731Wh
3BR7HwRjeGJXxedYOjnpIEIsDykKXI+VohMelBm4mGTaQH0g4/7LqHphf0kON1tY
AjN/1n4/unA12YwpXmjXwxlIPCpwolmXY/P7sRrHNC4F+GgCUKoIULx/y5p19HYx
h+YrOdeNWtsUWxKNSrM8jOjTth+wZBTqtSkQK+KtzctNn6dXBMQvSiLzTENC29p+
iXkE6qStWEbVh8nv0K3WspZpOBdQHYfkLtByx8m+M36qCjKCTyX19rbYJTDiTsVA
kEGZjpj/szEnSWKc3wCA6SAK1QBZ3ZYG+ko3GHG6wyHpex1/SufwPrtzZxZDXN39
vpexABgAPcGAUc/DSy3TGozC/yXMnFps5x7a+fd51L+PMcrL564jYI+tq3/LXFZN
+AuUbKr+1T4E/LBCchtCfQS5KQ6L4YH7XR6Pmuge7jca4MiBSJWJg9MCfjENKgOV
VOGEpoflHq9BNXZ8JJN7h1oTl6/oBKcmmQd6X5qdNJjhsB5kz5br/QehY4y4gCzE
gWf5eo6CjssUGMoi1sG3tJQAokGQPuMCAq2mIq63cJfmZbVKaVbCCBQO47X6TnvX
EqbD0glJtN4vm0lVW7B+9zwZOxlrwhzu3Dgq5+y4pstxd9KslmTq5cqxCEQK71JA
xzjEa76SLNqH+cmxadPDTgxB1yG+Tx1ju8pCWAIJkVmKTRNSSR3zWH4n9qV1oMM+
J0aMOV9qlbb3P3T9Tvycwwlu5wqK4g5R+ZsDtVKf51BEYubW5SYVF6X+EMEz2Gs8
GHc5jXkIHwCYjZh1jAbzmWnfjDSdiNipTlI9O5ElmvrxfEsvRrA9vMvDyKMONIkK
yNUuX4GScYtoQiB1Uvels0c0mdVSD6qxA9bvHNcw66YUqVDJeVJA/eGEDfr+675a
VvNTTnZjvUpOR7ZdL7pLi1T9lJbT0MsGlHua9a/CGrc8rZoc/A6K8JZpEDfasDuh
hintdXibBF9FXzWMGiicJxpv12paoxcTMzSPn9ruArga9Iy713YLOOO6i7LFcwEy
bzVWzlidgcaKXNL1qh9RYtSJY70v56vsjexjxyPWn7PNUENyt+STIBrVBHafvLja
jQ2/QULzunjhfQcQAxEq64Hj82Z4rJF75sgF+Du3/7jEsWX/sOeTBs1ucxyvOPl2
LNWwsVam7SSFMRRAT5ADjOMD/EXeYyeqnH1yTzi+I+DJ4okieHFJttHwnCQIjAaC
3b7bwPLeK44ujq8g4d9dTr5SDMX8l8MsC9iPhiNLgCIbUBl61IOd+BMqT2N/tPGa
VBK8xN1TMMQlj0cgV/Fv3kLiTFn2GouhZqN4HdNajL5KChjWhQoqaO0sDuFzfBJM
d5A+lPqJvxtv9BdPy34rA0rhMYVxEyXRbW1PPnvfTk/CsR0dPA0vtGvED6ALYl0l
eaGbbMIV5FylLNbJZzO29lmBj3IorTDQ3APFnTeQtwwnPkJTLwZr0qTLIt/TrR/C
Dmyos1k+HwvPruEjXJV0cb89UbxuVSmQSD7hkLgWWQOT9FZHcrRoIqXXRvQdBWjd
nGbFMzw0RMiGy4zQGLaK/4xH3KGe4/TClZhU0npRp/EpsD0FmOxkatzk5t0Qx6yy
rDsrjhndKe1A4jNdz49ZPZ21o2RDojKdwxruBTyRH3SnikIaYeb3LoOZ9iP2ptOb
vaDWYrm/NHJPNkc64pFGYb/RIIE31gvRALPGFD7PRQKElXMXYNsARIblGjlkT9pW
eyxb4yaHkil1ywxY3TY06AM8AG3otrtL+W5lOoSxvehzCYMCPKp/qpUcxjVKxCC+
Yg6Tej2G9xA+ngYb3O1S1KItG4KUo0trAWnjuIWOekbTWDvHnREhs6Kok4bHRcbU
HGrshxkjFldpSOM8sGQ5VwXPGFOSNvu2FrflhbA7Q2+5FwXhnUPOdPFL2+CMN0DX
EVtdGVB04WFmNk2/uucR2JIi539WmUXvJDI/ohLACTym1NZZyMfcWY0lFmVY/qAj
Rx7VmV8le7XFFP0D6Rw6YJR8gmvzynDhphzgD/Vm98ci9+ZN6ieTfwN+lVTAy317
sUVZy1ZO4EYGY0ME7B2rhkIkdWmqCsqbZSeUUTDhSR0UpSob+VaQgaPm32iFiWpW
3u3yAjVrmP3Co0iy10yKruqjAhnNzcs0rFBIigQXaAC8tDRGR40SQunGzVG8vto4
bA+/bnZT96E8gLal7lG2fFW4SCeKXOHGWPIa9+8x/82TjqeqaFh8ekoZysedNHjy
qbpO+HD7u6/dbFtrCc/rQaQBylVwL40QxAMxTgjng4JiEIRHY+D+Ej+Clygiq5Wq
QhCXaXV/mLxVcUmPLdf4W95hF6NckPnmEwWQoTRDZ5eiJ7qiFNDy3EquGIsEfLQp
DhuT177wNgGDSeVGZyZDkTobBjZlPwMJ4YJMaVj37CCms7NdZc+wMiHqW6U8WO18
vOdrud0ThCqDS50+4HkKlQSdnijmC9qJAvzFDRjPiWyVVbZsAVB7fHC9X79gnf9H
MZZCXSt3EJim0b9RQlhWOgyQA5mgUsXBmGDhJqVUQS46Xe8hkREbjJQEu4GI4I3V
ESj8YPtHIw5Z0KImXDFVZfu993vtKKkFXCiUC5e8ITVKfba2hMvXrZDQT1/IsuX+
Pn9CMiH6JadFLNBNyqatZerspyx/7RiEHJ76XONzAsHsGw99pDtgIU1h592uXF6N
seLLuiFzEkh928asnykxVtwRqeJsI7MadzZZtlExuvyTVr9sVccHf0alsm2MUMBI
YDHmO1qVoeTPmt2I942HgtL3FLIzDD+pTcSAP4F5wCnBpQDaH8ePSE0A69J3/Ehv
1WBXpZS7cave2q+MzEnO62aqHYG0NZlrOTeCb8kSdEymWWPK69Dde+mDBmGhBd8E
4E1CwYBUU2FDTJNl2BCIz9XJZezQ0s0zHJQSfYajRt0MHVGIpDqqzidprYesRQmk
dhcVrutLXXiq29kzJq+9cLVGCkb0n+MSIYSvRtwGWa87a5ZQWaqnbEFu7UWT3WS2
oge0XZMfYZQ69/F5toJ8daRPmvI5n32YO3ucHsQOaTcmM2zZEMu+S5IVo1GnF87w
by0kBHshpJtE6O5nXdH0Qjk98OLMu72/VbJ2lDh365xLWvB1LbVn3b1rAiTCrE/u
AqvVgC/EFxHlIQuX7mK7QTAaeQ/djbl7ImUi+4BFT5645sielRrawxHB85Ss/JKV
YypKt8VXTI7e92nqTrxfn+uwzFbzOoB+OgyiypyCxSke3HJA4lxdW/WHzAka4SIm
J++QFZIZ4HmbRnJoz/QIDuEoiXkXo+fgJMx3Nv7+xu+SnjytFA28Z98N9gMsahFz
W2E4hWXJKj7Pw3s85uLxiEbZEbNesUOxY1ZtfOTT/VbFwEa7xjSUpQ7HW2tMzO1P
IDG0CWUlUNnGk+xNcnMHUFjbywqjSSPDBexP9u1dRO0qubiVk1ZDlKZFD2eTOsHC
TOaLhskzoF67vKb8zRptP3XVADeEQEopjdRbN894CA56U3mT5mlrWPsc9hHnwRkC
8AqlHRHOhtvm/EuOB9iyXUcdG/aEm9VxNxM9L60U443vtFYh9tcUXG1qHgVAWIm0
uRyIud3roUzQNKBQ2fB7Aoik3YMnjW3eET8XjuX1Uk93ooVuj5QBAzYymDMxcV+h
Db0KnL3Pu3z32DWEsTWP5FnnsLrzGOBtbh1HzF6p/BZRYKBe6uOVRBnjFQrujo1H
r5Smp5t1gGPhNItAQghEaYD3PhNmTv32X5iGTQyhWgBYl6HQn3tM1QHkgTs+vd0i
SpohAyxGeEGdIwNRdFhSlVKfQ+JGvro6fEKqLkpGIAey+mJTeVqaeL7zWIH9XAaL
ZY8bp6OKpS651KRkLbxJvjxT4kcmyrRMCSB1LAkcq58okPBB3Q+lZuwRxghPhW+z
wrJxq6et2JFwjwoZBCXtmyQoLhYvHft+tdzm2PT0znBhRWjjwmoSn7x5bMgFz+lk
l7FP2hgShLV2vM/lsUHnP+Guqs0SPA0pY5x+AEKTg1Miu/01cj+Q+kT8xueuAQN/
YuI2ELgEh4Lg41sJoYQIiUw9MwIB2aHTf8X+jf7K2+c5YIw2r3osuEEvmQcXRSDB
Bdap6OPdHWWxdZxgua+pY7Hf2GmsIKp3sAprtqE7E8ih+CpizhFCA0p+gwpH4HqB
KqOcXJArIvH3HGLSupoWFiG388pgK8lcYhDjQU1jrYszGLzmnCsMvE1pBRXkGknV
v4QOmqPpHsP8YhNr83NqkSAhrKgNlvqt/OtTFyEIov4SU1gAx2oERhpfUs4uFdA4
f3SySHsxlAJO8MIlL6ESyNp1wg+vxIPPConwuhH8V7MybUHySp3ddnzYq7/j1gcP
8usHuFwW9wdhlXW7YUm9nOHoQvCrImUae6Uj7RffRxhtwu1712egnzKNwuzYG4W1
gQOUn7+7xu9G2prIMP78hqvdAMoDa7oKiZ2iqRiGLzEQ6WltN8gmOuxJqN1CLUJO
iLhxarZxB5uUgZxUw0mOaNLYNP9TQYAaO43lSA7S26cdduQfa3I9QevOzRLsSnJq
6IaYLu7hVb4kQkfxlvS0bRAz6LMCeCGnsLHDCl2UrxCtTk7oLUqWn6RUyJicUtRX
PXCinWAuKIqah14cQa6LOYPqrR8D/R/xXgbo74LpEEElqLcAc/Da1BzsbZ6ljjyu
VlZB3cENM8wNwkkfBmwXKL8jYGdsdxSUl0czGMr/gAKhB04nKzHlJZQFvsw6X9Er
NMCUzJpDO+pRx7ODev9NeWLsm7GvLSsHNlSusOcAkTYha6wWm3ySqTW8Pso6nnD+
J5psYVl720p3OYfSTeig+OAgLcp88Clk1o8aX7fpqfSR8VTCM9l0QBggS51Db7I7
Ty8ZZTQ8dg1R7E8Wk5MqXRGvE7fFUphrac9YnT8p3oiY0C1a/VrrGYXeLGbPXgxg
6wX+0x4EOBaLehpBgFdPRygmodTOFewM4C0dTq0BEnJkwtubzTr/Fy+QACEwNdrx
SCSh7WA+pBK5nWRxpAyu4cENlYDfDXEmZEX+k11llYgcuI6RB5/sw+yCEfqV7eGR
rheYH2OHkI7VyLs1wlSx970H17z4MUpJVqad53V4arFAdz9Ve+QQdvlKgdpblWyT
akjzUFB3g8Y5cL5wuIRtlRMZ2VCl4IaRO38zVIh3zD8JMOiLnv4Q/+zQv2jsoU4O
E3sFGqdfuhb2IpEfmI0PK5pa5AffFRGKVsown6B6vIoLx/ugYvH5ITImknZDrZvu
NNtTLDtMNAKinBV/lvJlkCWZYBX0f1h6U6XRROr/V+wIhAfCgkhLU61xtSmDosn/
EDdH3i6cFaJsct7DlGAjQzGsGZZ1rGegEA4KVeZMlsApZ7ctVVtmkPUgEzD9o+mf
6NH40lFEtIf2c43CbaxiGh7fFXFgYBX1yci5Ss3AKJIL5PfkrbHIJhAc28MMZTv+
zhrFf4aEeIZwNpZ/A6e/y8YD1LoZWZPd/bLylpoXRsUhpnUPq4ko7kynCeUp/xf0
1R3gc+Qaq7MSORDCjkQKeGWocaWRsMiUfiU/qy4uz3/GaosmkCMNhjxZmOsDtZOc
8CF0oaNOU2aVebdH44s9TEggPNxUuKyX5qWBbWKFFRDPyy2SAYyA9t1EteRhioEa
VrjDf/DkOxJmXWUC43+StPLLB/cR348aHdhWxe3Inq+HXbqDx9xrW9Nu5LUehg2E
3YcHoPD346Oc1ynBYgMuGzEcE4XRV4S0miB6JekQ7vm7AgGwyzwd58A3V9OUPNw8
86kRbTVTjFWaPYvqyxzhAgqCK1lnDDO8ccTCCrLqCMC0c9gyLNN9R7Rcag2BjI93
EfA7C8OyWIWdYJyaICRcf09UeiosCIjuTOvZnZi0XzB73nxUjb8fORqrnKTQKoBu
0vYTObvHpMZk8SJAYPHO6+Ee7tlbEFdkYxlin7Wq1HyWuMASkQ/g+DD+Vb7PEshY
Afb4yVqN1R0G9bUE0IWxSBf/L98Kzw82NDI+lh1do3YxmVQx4mrdkDdCkoKC2c89
SJ7H2Uek+ttTTYEW6pFiIk/atPdzsb9WZsEpDe3EiJGKDgMgjYRhTULRHPoC6xFs
NKaVy8bRfIzzU1A115mWGP+b/izQf4yK1RDT14nA5zj2UBhU9EYJJMWJVgi8i74t
JAw3oipSiQuOo1HLCutNYArVGdYFmptD3Z0NJG7lpq5RpBsnNj0yH6diCpoUVT1+
DSDuRCozjgg9znXVdYdpGOVKcRU2PbJfUAsCohUztdOQQ1I/YB/h2sA8WB7/2bLM
6bzbXjn9rF2mJilE0xvIxABFSN5b1cAhAZqt0Gn8tEMXeWKENXG2QTR2Qelil7S1
ga4uBg+lGKOfx224wWxyc+pq3WGrVKGj9byKBrFFG53l8MAJ+FqEvRs4gxWUXlOf
8Alxm3rfLyM5X/NPF76DKN9PWFziDSQY3F9QZ750wTHjiqx+1GQ/S+o5URuE74EM
5Om8NazbX7fgLfC+d9WPy8JFtDw/VXQmTYP7dGK2BZt57mUQFZgkIr69ZRHA99NJ
9MZEsK/TxLWEggTAhkUYC1cKrIqBY/uYQd6RsCku5n6ApvVrQxVUIVtyXa3BSdzo
IBoJhk8FkJNkNf3MAobfhvBfZRpcKqNxuWugtgp7AFzPUpMuEe+1l5UO0f0n7zuQ
tiznvAjbzVSoB3DMKH7R83f7CRa70yjZwMtd298AURta82zAqExZQef+V8dBfeft
6lTr2fFRACEe0FfUh2abfvXz0dikPec0yRuBpIsZykRJFFE7YkXsDCrPutYugYqH
FLPRZO96PgP9CYhG8StM4gaoj9mr1nOtbThQWfaWLEe2jmymAVbV8ZA4uxKwEbJy
N0KP/eGqDT7bwVXHrpO6dw9WJeYhUMr/JFJ1JnH+1teMBkcCyLPu8jOQYkAfga5t
LXD1Ursqwr5FADjbnmuL44R5E9estObjfGAVskDkX4fzzpb97HuUfRUTuF0EJoxq
50EynJcOS2rwu3Rr15dBF1sZyWRR6ZMJBIKHeTUK7HfZNaFRdauVmlU5zMKo7Wpf
pOhxg0wOzZNYbFaAWYyzGJ9yWb+hGKXrWCJu9tBFmGtm+4H6iS3YlJeqhqRBXSNy
Ir+Osko4/Ajhfp7EfPpHdfLFuloJtFf/cFO2/f/9o1UrtwUga2o0y0Bm5qjLv8ix
rsEhFsoXTbOFqVHjb+L1aatsQc2IpgteJ8gJX91oStjxJXUqXKAa6xRiMqoKr0Dc
x7OlculOA+4vd1dUwjNjcz/FzTTAISGsReK8WePiki8ajODZcfXLsJqD2B/a/wT2
PbUglU6aBCvqLLT/L0mzYtGnji65ahYx0XyN0OUQwDVyX9PKPExIbPXkutkD9SdE
2xOEVDnA81AFunw0gSwr3M+1Rp6cNXIShUtZ10/tlD2zvnkJwToV6fgpaxPhpPZy
lUAzToT0yHLD4QJ9dh6kUm1wQ4Pc7EB8LQeBEZyxx7AlkTbnIz7eZd6nVpKkSSEI
Ly8QduE2qW3XPHnCffmrVWJwNy8mPMHeSpgaW9PPUf7zXDnRvrCP1m0DYduURqrN
AXwdexnu+RON4UiZ+Q+5WLmXFv6yMq8cFfJxmbxlofcoDgRw3wypEuqxpXCU6yXK
BmZndOzPvY2gRH3J6CvEkjyBoxczPlFOiPRdD+WnMbNa4h8S3BdqUrINab1EClGS
875CqyPsspqc0y8JhbglsFKVWgSKhvzPiUjbSR6M+eeXFEG886t05fFINLfT1nIK
NWzGTuvsT4fuv9EsxYOQIRklZ0EtNUssWYgvh3gXDJrezZMAlNWcaczhiIEYz8ML
WMEcg8tV1i8OyJNetkdq3dMaDvv27ahx+bg4xn2N+P2xghkbO/yMgtVb5UmH2myI
kVyTSL3PbJWA2D9ZuSTG0HdBnqNsr/s7MbdFQzi87lGodi/akZB6B6o+14ns+jaW
5ossMj6yls9ROGIcEV+YR7ZPFKtg46oCNsOCNnRSq2xU327yUjFXHwdT+ppgkABM
tTw/sRwCpuAl7Ok2Xxb8U50gTRrvocnR7wVt0qpLisz09iKgynztq3zQJ+IsT4Wp
2ZOS0mxUJ8h3LNeWmhb01OCQqwVyviroX2/wZ0EbhVjkw2wFyXo7lOxC7fLWA7B5
IbeKN3iSvA/88GcrZJJQO6ygOwXBSjc05llgLYJvlWYkZ/kdlhrJBfzIKpKBbEUL
WSGC+/dodHLnJ4wfGPm3xlrfI01i3a0g9HxMGF41Q/BgS7NH144S76+ZoFYFx0ap
uhjrbC9+2LGMYCT8WeQkHZhJneEmqHuEaRxqvMRLiQLfJR0sECGBJAfhLf7v4ksV
uW90u8EnQ/YhBxkZSto3SFAO1kCyB0ZGGTiBINfczlc0QC2VDV2YQL8wTruZgC7f
nQBcD1EFdzDmj4vuGT4Nbxbe9O3S6MWVRPIpmwhUXIXKQX0FFsHQlt/wOyIWkD4m
h4+M/eKRMrSySxppma+mcBZ1/ZG10wKGk7lcg1WZkdkOg8I5tL6f0UcJbqm9ptH+
g6gRyHK4Dr6dNOo1NM+DqRyKNwZ7oy/m66pvmLCB9ZTp0Uckvj5OwxqwMx5P/OY9
c3PxfPQVhRQ/Xn+MXtfFalFcrSNnLTAG25IJgrX+OWb8c1WiaMpntuapRERX0jk9
f7XlE8IaC61ByVBuhjDIIgBYFcJYlOtXF2kJFT1M9hokv0Xhne2R/z41f7TkRnsZ
yZwsyHbBVgabVJddQlJRjnmOQF47+eSSGzR7dQIjZmfc8dB3DdRKV0EEtpSG0Dyg
t9ATzrsmhfsavuk80iPftPtHdUwZBFhCPcmk16zFX6Hc5/oK2cDrvSikZHhvbVfA
EoqrGlsZ4OKa2GgD7ifX/wa5nVpVjLyeMJmwRmqzjMdE6QIv18NV+5MisGsYnjrz
9ITG4psDnnrcVbhahGHcFOLGTloxIaTwe4VhiqHjH4tHud9tBugxd455gAAsM+aW
ELizi5VHZw6rrYMFZyzJXlcZuqKi+AYPKOw2aEcRQ8qmBo55VKn1Y9vHOKsxn+cj
7cb948IaRfVok9e17a745L7ZW/ZasrdbeK2UCbLTikenpLJ7NIkzFbAOExXb79M4
vSYX90ppVDJdghW/L22a7i5E+J9GGeue0p2TE12hjf39m7w6TrKUVZZoHbwDQzLk
iJ5ZefzIRDfvv4Pr1a6jvwRW74jIC+Hx6Y0hfhmWZr7FdwgEAXbLfgl25Z7ugUfq
tyW44K0+Cb6O3iSmD1iWJBs8bh+urJpZ626kNAM0oOFqwipLTV24TpBSbWSk1Dfn
iF9wlWwCaKzK92pFnwXsKt8R/OAhOQ3U5zG4jYbsNV8fwH6WyY8bCYU/iKcv11pD
ZXIxikykUVNxvrtJgc1lBnws11uf+f8mezpG4tfGdOU1XQJWW6zhKfvmgoIRoOGz
mgMGqmFPI7ijJTa3oA7c71lrI9XDm0KjAhqBNixL9Gzp+bFDL7YwLcC9/G/4u+3m
qOuM/5U2z79Q/AuEMc9rCveJ9YTmnfiLrUxWRpI2gODRrIJJRnlRolOFjx4ag93V
hlHLl5hVtqA8wbO9T4XeiLQ7X1wuDa2LBHm1/VZuQtlWnc+bEdl3JUEigSDsrOLa
Ez52VGk20rjb5M4psipWqoYGhx03USr5zjmJbAHhBCY86jOmq9jsjvdIZUsXu/us
FgjF/HmtRmVib49TS9Dq+cKeAu46/gypCovRVO88x3Gs9OEUvqlC25hU/Khdmofz
KCUGXx+TBjFdu90PuCHwQanUnGA2mVdG+YLrPIFB5BttdmZPwBnDvJKZ4PxKqo1y
+PNh5j/y/8eWiNUeEzihVLp2s//7XP+Sy0extK2ggkAQ3uw2qHDnOVKA6ZIvzREz
`pragma protect end_protected
