// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MDfBxmTM0FrtwAgwVgr+oCT5lvqC9cIryk9KBvRU6g8Tgwo0/6em8M5FVH2MyTUX
VPA1eV6vbuTINYDkf4ud0fB++z8/nc2fTFJbkRUVbdvv6V+vB5l+8Glyz7S3jSVB
ghzRhAXQtpZzY9nYa3PzdifrKb5mLEQ0OaE4tznFytU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3280)
c0d+hNdGizpuiFOg32Vo1wUo/oLC4c+sP0udCT3VVbw9PmF35BG9Af8JNZwht8IN
dkBsEiwmxCnX4pREaE8r08sQSAqCaOtlWKgF1psIyaUlDrAFOfVXvkyDXM2QHtaP
ncfW90tzdkwzMqVSJKrfXqoQVatcZdQ4qO3yP1V54AJEFgsXHP1YJpoEWClngn7K
USNCYaFy1IPfI3itibRr+8Q27xrG5VbJm7ARkouSEsYM8JZ9fZNKKbkxLuy9u3LT
Knem2I0eKLNcbAp2QunoW8S/DUYPhUOFLeybBJOVBz+vcjMK+vlEJMfZDkDRVsNL
daZsCKeXnNqwmOhaB6yWpqp9QSm6EEk7Qxg6hQDclYnwOuC05FJHQPSlHQEeKvHC
BbYvWzzSGj9i3CR56lfCpj97TySwFPn2xOe8AiZuHXGlorXcvjnDa5DGf+PDxSY4
C2IjINeCEhImWNpvwsf7ROCEau7o11mdNDNcXhG+wFxXwYYTZIlx5xXC2vQ4nWmF
KyXfYRC1hyrcFph8vMQsS03W+me6Jm6kgkuhDlyjIrLmwcELONDsX++b/PF11V+U
GOGRB5mCaoH/IG5i7kwTjpDmNQVTCUNG9M3zdiASUk5G+MGTcnQuPcMgCrbev1V0
oPTHQ4a7xA2q3+/5306qASkOis0E/ILLsaRs9R9buVyUbKbZR9OqWV6e1z5VA6kQ
V0n1Y9/jXFXa25NgQlAseyFnjkO7VEs2N9GVsHfGAnUyy+N3bM6WzceNmhPW24d4
D4RaInyRdMnnV3XVhBud17CPly8r+mEVExWPW86WdARu10Zl/jsR5SDzh6MZo6Vk
toDbMTmX8rHpI5GFshgtuDtJUj347Dcu0uKiUcAHflvB+Fnq7ZGgXgTL9uHYunRx
B+6sIzIkPvVvNVZT5YtkysrfXKlAffqUv6NdPEpMRuoHnXbXVfgkhqJZdNwzR+RG
Yg4R4qEhgFHWznd9xxdjGGrzR4NKmHyMDK15tGD7+e2azqFyCOOHglowh8OtvXeP
eqPLHfjneAq5cHKLrZWldchzJqujc46zxfrcIv26IxTGVw0rUR4wV7Xezh8IQMmE
pobUMF1F6JWGW/O660yssrPmoUBlNu6FJKDMTFdpmRzZIrli4pJVcUf1NPf0r3vJ
D6DnjFSXOnE90UXyQX2FslDbEvZrA3SHjyxHaYs+xHzMIGNFYomO3bfp4RwiFZrs
eHnZ8fY7iBXHmmeaRP8AGdyqjqlSvutGsrpdA2R+OAuXDYSR0Z8LquZ4x4GPRHSV
M2bzfodMh1Xpi60hWZzAYvfMZwVbL/9k9HaRYMZTbr/OJTtGpk+cdlh4I2R32s8+
ujsHZrM6aU30UjhUtC1+QQ+wUalbw3schBgoyYpcwAGAAZrqpVCGoAcGAPEkS22Q
9zg9QVLGjiidiHFmblB2I0gw8CVCEkuok/b4RqB3owv1HbSDfcOhRQyiSQ0LSv91
b78CDT0fUIXsMGwAhSMu0biBD5GAxTNcmBJLGPEBmFFllNLUcrBi9bziCi0wkFwS
I0rPkYLZKbE2HyysoZ1JvoxItAc7WD9rYcbwbQzoY7ZT1EciqA09t9w5jRLo4ksA
ZVLsBlHfUv3XIlMsti8L6Yf+wX+JVIz/QGDfPj+nes1NvjerV+fq1idV1x3H7/wo
DNQAR4ZcCJG9nuLhkZJ5qeQczkfiuGSgK2WK8boR3u65FKlG9d9PPscRPQGR/AJz
xmUhhzZ7b7iRPh2LqYpIoDLbJMUldJSlh3omnPW8CrP1LGE/IvZbDdy0ctcL639D
he6uBXw1vnbg1I6XbK3pd/2hLGXZjMJDGrvKTLDLTeD05wcl8rhBLv0CSvsWHvAe
0WvKAwNvLxLMqSpS3QsESuAegmCFlHQ2oLcO5X+tRxiAbHkNaayOLPWxK0CsZO2F
jLlZyvhIqAXOrf0JBSG5ZCPaG3iLoigv3XcEmSOYUD1wLeQBfhdg0/oN0BJwph/k
a5z1l7i/IxqRW9z/2gOojXHofk+kNdM8m3C+i3yRijSLOnB1Z2wY2Wr9FEtbsVJr
GMxfvIWDHZTxmzfkQpkdUoLBjz+LDtu+Bp1LU0+zc3WZQsW09T/2SrX3MAXzTRHD
gK2MCPK6fW95QJ4hiRz0Y7+YDbBIMrGjdSBZNGEkL3iCB3lzmAFW6EjYt53UkKhd
Tk3/Z1uN97lOs7bOiYTnyftEZmJ8QvtWs5ulWAam7JMtB6Zzgm9H3WLpXEpbEzAZ
x/9CHR1vd/bS2p63wcwMa2O4sFpQx6KkNVhCH8bwc+zZ2aseIHYGrgAPg4xBQRgd
PC40aQbG3k5vyVa44XJvKFvcaxBlL4+YFPmx1PxGnygQW7rqIMiX7vjHxQSm/KXu
IKTKdPx5O9ObH3Ogoy/sgZF60Pv5FX9lMn/RJ9Qs1cYS7L9sNGlrh4m/GpWu/x97
ahpSq8EPXcyu1rI3DRBRnPy3RL9aaX6NMTOgiz8kYU2C5UTqJ7LDmwAwXROJWaJI
9d4c5BBDKsrzI33B+cK4Ximfhgt2Cr4L+TcjAz5OO5lJh/phT/uO32iqYqL01vQH
eimFk3P318+ct4WE+OQ6WFtRAagitf7k/gbeXz6Hg6GPTsTlrQntr9UxfL1ye1kK
1DmELuEv/VO8Abk89blT6ba2y4DRw0iRAimteWpMPMfM77OyHzsv9ELGxE7w2kcW
ZGs6vhGGpn5caWAxDwpI1cbPxc6OQ2J/Rj1fHRVBp53Bkygg5zCgNPpknXK+0x6d
+oHrkxxpoGJbyi/GCnB47QFBgPa3yEAs2ToENTjLwZ2VUOCsB0Xhi5fGiCpLdpZb
QMsxtsdI7aiu0vMa636wmS4gJNlZIboqaZfDzwTjNM43J2kjUBU2spsvc8fcb9+Y
2uMNa3ZSXFfqzQNqv4N3UFII53s03Bou0DA4XKjGRtCvfZnK6QptBEXfdUOKr3uE
PoAIT3X9LFAtlaIEKWA8LTqLhLXinT+KXkQZeaZ1Bcu4RAM9/0CLOV8XeO+bWQDz
Q+QJLCoR/PQ+v3aB7UfEqW0ZmQxfjNzKHjm9Q3WRLuxU2FylPDVuJ2sCUOdQA06X
PL2MitKpZYrk6HOSgCxw4hgqUQVNjfk5rD6BnUFec0mB2mtZKzFF0bwp34wk56b0
6WlijsxCeF3zKE022vMJIQwwzghSnRqVgCcIFwvTFqvsvkENW89J1HVHkuMxMysF
UbtrPMNMz7rbgH+hujF0+BHAHSt/wK1qSOS9nkLufg0hEx4iQGM+62hYJzPCivDL
dLvSw/pws3fMKsjdA1eL+iV9wtb4o9qzic97lz3HaaA2l1k8q9y+FTRpf9fjGpcC
eJyO2M/y/QTBYjBqyWccYptm+A60XH1dcqTpri3KcBDjIADzTOMt9SQn9CkAiDYH
6DVB56fLGn8dXNiM4ogzIAp9dJ2G3j/Yf9A59oZaX2wTHcjSPLB8sIEPbXB5gPD2
Ao0RSFINR2isQwQ31e9kVoI10BhJHd1D3j0RJ3rW/OQh91Vix85XPuxyMnXYee0S
V4fIyuMnV8461uvhZvD5x/55MJ3oG9C88SgrcqCycgCsfqky8Zm5JSNJTEJWpJMV
CeNKXvTBA6N2GjnfJ6Y7+lvaYcWNMF9QiEW+oC0iLRqS2Xn0lFS2xiknznU/DKwy
GjUYFkTa0+jIp6294sp6NuXzpk6NDAPq8FKDStRJgK0zYLhIpE+ytSbmHWA0Tvyr
QMvub2sye+GsSbftvmJdO0IPGRlXOnJ/Xrs6cCeikJA+N8DSKqUhTZ7wSq7+6wM2
uInqXfjbMtTH21LnUD/YEidR+v8jkYSkuGZIeA72GWyGQsJXZpi/YWHNLQkKO4fm
k7HbYeZyCKpwwZB45srQ50Pbb4looke5bnYPxLWOjqju1jQE0tJETtwlhRUFNMcj
/dyem/r1b3GMKbxbHnq6GfCxcUV41Q8cJ0BFk5WB7vSif4c69iTrk/ffjIUhjXa6
Mu7IscOjmUlT+QJ6x4PDJUL1S8GZ0Ql2/P8TR1uiPJE9R7nCQuHJOa4nuelEbDXy
eDdes6S5U3d/TIKaPaCOB5N+R+8+S3iiH1PIsu6rrA/K6lwu8pgEZqwOztuexohW
T9gjs9BDW0L7vWx/10czcEAlAcpAMdXnsoVMnLl8fR9F0fKQiLglw1tR6MBItwg8
7kQ+6tCfdZEzr/i9VOeQzPbd/teAfWwWa4rpZke06jfh0q3u53zhVcrQdGHx6yTb
jlKh9X4WSMnmpV9e8E+eavIdERxYuvE9oeWCycbamlAW0TfITr32nTxFdoyoJRiu
ZR702oZEt7fQ6Sfa8jfdPZCuA7I0kKDpxp5YSUUKSbM4KiaazDYu8O60cMKE8uoi
aqllZGar2cg3Yadyv93K3A==
`pragma protect end_protected
