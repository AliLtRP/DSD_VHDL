// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sQsNqigXbz3G7JYiUeGtU3VC+aJHebEYBqn8Bzj3Nawc4TuqFrm80ride1APM8A9
W+3Isxg8+yQd4YPazuTlr8sOH1AZalECA/y9Vvv2YvlERk5UxrI0KHYmhrpcdxSK
QAUVRbR+uaxKb5CT395mXVKtxyviCNNFQ2+42v6xRPY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4784)
LsEuFFpcYbjxttYVRGz1h/qBEXdzG9KQgxaq6zWX2aSZXjsEvmZ0v/hhWe0yPQ32
OnkoXzMqao/BJbqBM2Mh+C16IObIKGhXWkIY0NMrt78iubm4+92LYZiv36k0VKKV
sD56ABMJz9xIVqeEF8Yc0WrQ+O4iaXHQvUFx4ylykbIoq4NDk67YgOj+vwrClDRe
K2fxFXvdpv2fot4LAn15DJOTYRET4f+Fx3UFC+PaR48ISEXJJyPjY+et3shhjh1j
RT2iQbUEi1CJQN4pR4Djz5XJCnkrUh1g8eyOIGjLinKKi/u2h5o50VxsNJxzfIP9
0+sKlgWrFd+6Qtik7BT83hJZxjRiOUD6oqauqIfoy499qQB5sJqUguaBSh2mJhZo
+Z9w+I/oL0Z4Z3iCOcH/MCQfuWgqGpU958UGvWmHT2RnW79L7gfU7oJZj5uGgee+
+mY//XZr7A2Lozp+PjRxbH7ZtBD3uZe46TUxqs4lMuB+W/QUKgK27r8QYn6aG2Vt
3vC7Lcg7ipTIEEKzxEJ563se6po6fivuZLvpIVPqHaBaXg8Y9ImuL23vwoi0a2RJ
NSgvCWlf7dftlyH2xl5+eAdB7Af2rmyu4XQevFW+DRzn0HbnUGEnhgBRHS6TH5fY
RaDnaSMvFO5VEiVj1BtT9NWGIuBQI07rRmpkqGLN6fZG1J1myJumcjRSifHDWY7D
qNf70tGrqBj6qEWmgATsYnedhLXc+o0tkBVb6G3kXg0ib5yKkvnTaRFxs68wal56
cxZOEWF+yscD28xPGDuhxpGHdgHs1Ki7sTEWY++kXg4JynYhN+awAOqSVXiEx4s2
3dv/pZX7I6dD5LLjmak0bLEeX54RaNld3B2ToaqrcjQqOjjv4X7tRm7lm79lHdJL
V61S77krwLo1nmYWE9bFNrikSWMpNsl5bWsKDEVIMlLvavSpp05iom7JUkX53F6s
k7cfgRYXpwCAbWvuKm7tIcgmGzdcH3fkmmvUobFZKQ2WvD505idqnUdrhsIzWxFY
2gfgmbxuN5RUePQzZw/mUvRBSTo98LmhkwleQgZXcDRSX9jrvwWSHpAVzcEjtCyl
6X3TwJw6hCnQz6IDGQFkqmi6MONPO+LGsy3pEqpL0XDS+I+FWKMisgrvPcC0Wq1o
JXjFElNgTLJnMhscY3WcuTra9Eq/wLZGCPMWTqVJr4fF3mtKXgOPuSWoIobccwtU
DtYZbj3cXgkh+vvfBOsaCcqb8rc5Nw/2SN4wWyg6Nw8tTZeIlHBRcfZVWHeLhZMp
bG61NnCmWmO8bivJzTJOvxMfRDhpdBDVabQBMh89DpuVW7RlVnH3cRoiPU3n2I3z
P9bPNeejXuji3eaKvj8/2jK9dmkH6NVDFcefS9YfGgFCH0CVnLHxjvTNWDGbj80v
ZtRmV1LG8QbkF/IzHsd5+9Fcg46PL/r+PYhlz3nTU/Bd9X3vFmO3Jsf8Ya4qJnfT
huW4cs/SQBN1O5+HJq8zKSGzZjePZzpMcdeAQMIQ0DZfpbqcj3tglnOCoQqZ2cM5
oJByfpDU2EuR6IEiQVHh/wNfhpjbYeM86UETw6Q0W4wgdvcKtRV3Evq+FKeFqXIx
E3aKNhFa8dL+jmFDRb6UZrf/pMW1DlSIfng9l/9jWHJbWBL/Cx3mV1ZjMWN16e+i
wnIS2123MM809vIbMAwePGeuZXle7sLtjbIFL7ssaG4w5EFSqio3/kCWV8xC6oM0
NETRdtl9smk8NYmXyPW7XS2AEVEX6BxN26l6l1GyhmpeS376t8NBOBEH5lpT6DF+
SaBuaxnhOFvGHycIESSqyCgDfOzvPtTuzZj6unlkzDoRxQGm4MS7vYkYGaxIEMc4
WOF05Wtxi83kCEqblVKTJAZK6xlTqDVq9G0FiRDSqnrQS9CKlb9BxKRa4cz6cfcW
ua9beYj+LNoOUBux2czIwIAIkPOw8c+iiSH6+3VFaW860SPlrf4LnivTBEziwnIj
8BGa8fP1NCC7TSuvQZ+Lkq0IefsoTs5noCJ/SpxuEXtM07h5HivmPs//3be69Tz9
0pJ7wn0e3UVxuYzGowIHyyofPHiHv0vrJ2E4M1YmUAckR03Xr2BTfkpbT3iBAgYL
PMdq2ivyS5nCFndk0CeB4Kpsn0d8AMrY7JT0XWaLEonmnu8Odo7PXH71HcSSItvf
sWvylMQISYyM7BSEDyWwNwklxWEpuHxk2jQjyqh/7yBTWpcvn4JHi8kY+fuaLk/U
7I5rr8WcUWGsATntCP0FCKb/zDb4Snxx6RdCQ/zg2pjjhUWZKAd5lKjRLdTXqJyK
DcoJZc5uHoG2Iw9XLqDhZhgZKZstCfEgv5LeRuC2pNCUof84HoPYDLszDXV/KhR1
gcBzasKvkE3i4a+bz/NePSAQDSViPVa0NPDg34m8sP3kcA/TrgkVx69GnFrw5dTp
BJMeMlHeKC6+29EW7oZGmL0BrNeHGlcWAlutmMQmIEDybOpw3Gz+KLgH8CU6MGQT
Umokn2BiCx7GhYN6f+yn5tZaiYv9/ALpurF9sNGli6LjKmg6kSspPUZgCV4i8TNL
G10AyMBgEuYNqxQagrxEoWqv7xbHtSCWep5BpJMnZ+3dyLryx4JDO1kuz6w62jwG
OGZ9A6Tc/UdULxNGat28yswa/lR5Lhwk5PxybyPkibIBmVDxtIWvRdabJZwGijq9
JNdBu9V9ina8d115Cg5Z456owefbPGdQNQF88xNYvmXyMhKa516+GuUyh74VyedC
Np9KLjKJy7qx58/ruggcoITq1MhsKZkfSyqwZoS/iAhYCqT7sd923YqO56O8Hwyo
ZAvadlOUql6BwoEFQEsq/00vbq5ki7GQwaesiA3efQgpvjeA73iIbmfPVbUW28rF
PkEdBNO/vxXhvcJr4YOhXeZtxrzTosMSMS5qA0uvNHs21IyqQqGMT1ztDT9azbiQ
zmoqo99GI7b6AFW9qyOKF4DF76RsGn/yYLtd5NLUXH3CyeFr4TIkwGb3opRZHmmu
fco+1vN7iBCfQO+65UwgqXh3HAI7Ei3pGIboOJKSfeFnhQbB9JG2Z/eLcn6Iw07o
o4zhM0/gaGpSGva+Wol2t5uxx0tAWJdA+SsV1jn78Ma9emrhyw2JJXP5FX+KD7bU
WzymsZEtn8Bv2cMJirFnBh5+HLohzzdWyY/RqyKRBg9zqTRVuww4GS2M0NfVwMc9
gPvEMVADx5v0gXT0s3Jr40mqybfN8LFtcBoUV/SvDeF6prJijFkswkXiqhuHYU16
LfXlXXViA0tejw9CB/s5fsnPqjvbGgw80vKhIZK1jk3j/fYEhcXrVMDh8wSRVKVx
RpiH3L7hLUgHDSku3VotrVc86Jih+eD9Hnh8Vumzt90QRlD3yL3K4s3edRzszidS
B8nd7GdyL+ZG79iGyNFqQcyyDMAuFxRGDBJvaztYuatssrV2XPBeZnUqavPtG97E
jkpKeFb4N9DCyNIa/aJkWmi1pFxjLMD1hYl36f38+5AGed+O2A6XWPuj55DsW7Af
zHChrKgxsB5LP+7G3ej06IIzdQtO8ZPp9OvwSuNExH1UjVbBa2BqzLPwpGiVz2Ul
x2SA9uZ+1YGhH4k9Tc9/gGcjzZA8toQyuSuqrxpgsnG3zbl3AlLPSEAtLJplKiTp
ZgEVQKoOxGAtaTXlpsVJqI8Xke6d5/qqvWjRX9M/iEHzn4pYOluB7UiR3ypVbvxZ
p/ePuwMsauLBECJJzmU4cLr7e2yfBH10Hhiqc3IUy8bqiepwEBymU3pp+STKEtGp
CHgsH2hxZJqqjL+MhtU9SvHc1viM6iIqXWxkRRUtG7502pEy7bu0MG3GlatcrpW7
zV5WTz0Sx0zf4DCM4KZ/puEL/RbLGn+T/ltRnvt73IYZjun7w3SxShh/wqYbM/pq
F/yhiHpMvKbqYgQFNGAab51A6HIZnpT0xq6l04YDs4JS8gSvDL3f/qpIaEfbgXRZ
gM6YQ7Cqc2V6QZFS5JkBYkDvIFuvzzG7ZImfgepbEQJa769OZ/gU9jTu4uNhumpS
8yfduhOPPBns4p/v7VJZ9Ume1H+HXvy95s7Vu5QwtlHbYyb4ti+65A2pWm1MV1Xb
13DetmLm0yUIRGFQ5DZpbrZAcF+xbOflIoeGQ24ADVjvnBLxmUMzLKzsBckIU6xn
MjA4nzQ++Y5lSID9bzieYv047SCDbiaYzKfBNiuuiHKzbOlh03QY9rsIqJUem4O/
TQUPekwk1cVjud9ZcEBCXgZWvsyJ6SLJ5O5cr2Pmf6X91pO/RDuiMBCkKb4nzDe+
yEXb7VNJo9pqXJM9ZBabKTZ8/aOnU1B5aLDQ0ZNWSYRMCkNmkOYaQUMBPlSXQ2Na
MITb+xMv2+S3TPNHmb5ayCF6WZyNq8j6rif2DBQjFqTpzZd+vO3q7d0h9bgRPpqd
93/kCIeHm9LxoO2cFamN3buw64TbNIaF3dmRC3B+7zIFUxsezQL0Tsty8xwMno61
j9Fy+tp8EPEhdc7Xh/Dk5zcaerKEg7yJqsplHDH7e+D1qRIydJk43vFoPrr2oGb3
YPGFojBAYJMxKN0+ttMnq4CRGc0S9yQP3AZ/+3aS7V9/mwWqVEwh9J6ILZ71LdQI
FgeniC5M13nO8b7zBYELpMl5bxb7oRAYvAlnNLSqBPlkWFoeXtnNr7Bkbz2dcSr5
AOiqJEcQHmbIviY5Ze+tmmzHOI7XqvFxiwkNbKKR+3RFJTn0owfvrCe1V3LA+QM9
ORJP0OVjU2n7iA90Lt35SG/EGPj+BOOFRwEGu6H1e20zmjPMpc/fxqnChrIFPVX5
P1Q1OO9OUN5m/YckFdrZzBylVS942kCXO4vbVcYO38alJKLzFX6tQgsh8PdfJBT2
LVFRpo3weM4BNWGvo9iHZhd5PGml2U0DkOBO2Lh/e2V+Y7LpbmtD0ANlyC3cE0ed
GgeCZiN0VnTmAfoXj8CZf+wPNI/MOi4hdREbdQX7yX47Ij0uIYRy/9d/Q4/SeQef
nLgSlVRNA8svmNExd76wXp9SIHT4U+ArdjjwPzwAykfOfqkCrteYkjNyqLHz0GIP
APTcPQDKMgsFkGMzyln4jq80S4G/4jpMJE6Cfu2CIx37VyS4zkQ6/SAiY8jj2P8N
e+Nx7Na1p25ihk22ChZKs7rUIBporRyomSMtAqbNz7K5Iouv03ajyfpK5+hH3RSp
5JFPSAELRvE1FOopnsZ4HPEWD4iMeZjZ3f4Dp4yGlBJQHsdm5AIAHV8BSHtrblyz
4ekQd0eluux1AxsRBaL0mc/uv+Nd1eeWEHc9/yIyn1hqmCeC9JE8wo78eEuloyuP
1wKJoFBHsUHfTIdjdzWGsgupyaWqQ4nWAWmDgTiUSBYHcU6gRnVCNCZsWK1U59ZL
lwYBJYaSRY2USvhPS92vZGyv7MB60wBBr5e8LoCm6RpIcWy/PAOFY9bB1lmMT7Vp
Xizn7ckmfqtm11FUdGleLjxK+77oeK2XYad2tjb1ZnI7PSQ9JLFtj7k4fy/+BSIq
GWwLLBCnSE+Enk2XmwNo5AnOjkgrhRtgD9gvsgXgPFP7gkidVVqPKH82qN/SV+LQ
EwbSldzG5DpV2dpjzkQuB97Dt9SyMeVYMEpxDlo7LUBJFtB6FkwzJp4/vRmXOGfh
78qjXBAj9B1VeXHfztue2A2+0w2tCNOzTHqIn4BCxDQ6vYGYgF0P1yTiQRV55tCZ
/Gdj1x0zfOkH0AGMpL2F3wGPT4DW52laV4fgkInrNmNNsBu+qgfYV/k24fy1Luvt
Sks4/9QGo4NPUjuQE9oZSCq868pJL5EerDYz+F0f3xQAVzoPEQ54yEOiXmbZv6zl
MiMXaRbMcQWySpp3KAUSwISsha0uRBTLBWPjEP9/qGfoiCqtlUpYrd1GjtpQHAto
i5dRlpFB3fe47dUnYi4i7RvlxUX7ReeL9sn6b2ebTK5btyjgfJGfkzL+GoSDWNNH
x2Cac+7RpmG1pUA3j7OSHu++M0yLVUUCE+h/yXN3NitSo89eJsnEB+w0WQrue4AM
xkj1aDfrJwxrTfv/5k5NxFKQbTM+lxlHja9XRtyzVJ++EUCcXD4pJL1FJNt3cEMs
LvCetWJuizCCPsp4xH5zXT4KwaAIKzPCxi5sHFTGnD0TkyygbyYDsV8zGTo6AtQJ
p4UEI+yBYUNnY+vt3eoEOi8nxrz0BBReZ7X6+TlHIps2J6pyy65DHOj00O9bkum/
K/Awwl0KPb1s8ui1kcftDNJfWzjBLyS9hocL/t9e2GbB3WvaJ000JWXFf9n50amB
2JQ4qzEEgZbKVXuASnBKvrqBm0BHvLrmIutGv4FSSymJUy4sXSredhPg6wZ/YPpE
K1+lm8Jd1dby+phyMMoFdwyOTwBrlsVYIkbWlAb31RI=
`pragma protect end_protected
