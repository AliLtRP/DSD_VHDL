// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:03 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gJeipWmv/KI9dpPubID6tUYsRidITAtEGnLx3umaqAIWcGFmT88CtPsYMw+jw02V
a+3Jo3GIRO36pOjjoeof5Erl3o75oPWFFV8eAx24qZSzdLknVTcsTux5xxTgi/hd
UeehxNPE5Jut3dFqPBCYJCcHcX4WH2vJQLzfTfowNF8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11488)
YEzj2wXmgHYxMmeGUFBgOBhhZan9f6rxPgW7z2sGEoGeo5vXhnOZau+8oE2WWzl9
8aPsrmXd6wFMBWo1SMaPYdO9lUm+xQQi5TnKp5m/FAvvr4KJcFfxweik5ObXW8rf
2T1OMaoXiWdliM+wvMxQ3a9w6Jy+995dQignVtqyaCQOOrX8GFcVD6rQWi0bRvAk
cvbcon1UQfpnviPcGfodTZDIsYGECsMNNwE+AL3GMYWaEW8TulHCOYY6qKijABa7
NU4ymIuna4mekjjdyuTyzJYkVM/2XRnEy/4ABMlIi/ximxW4kyImmdM8PevCFqxr
SazAOomQEVPK2nwZceegt6thCmk+bSi/WcNgdebbBT7fXkl+rQaWqdTumOlEeY7P
ZPC5YSsCWZNpRPkAN54Wu7SfJvFDXEn9YYiFd358YImc3akBWvLgtcmbPwRzxEGn
K4onCB/ifJ0LDUUVR8+2tOpr2ESyus5LJ7fz7up/+NPMhn5X/rEX7up7onb5tzv2
X9By428eurTVeH3/yND9R/d/LkhP5++YSQOZebhxZhRuG+O3PsE1GUqVRVY3o/Bf
5TFyZmKXjxlmLJEqDRXC9VqYKk9XjhlNDVVvHaGWN1t53qWvGtlxQMW8dxz9Jya+
HjKUejosb9McwPUknCQZw6j+q2HcPmhtwgMFOeaSNxD4nWy3pcRj4WyK3pDuiqb/
AiuhBTahP3dzCm7sKcLst2xyLpK0OniMDVUP5AKZGMtkmmHlbGsQLpC0yvjOZ2I3
PBrcogSEfgwltBGpU9ZhbOI9TyPZq8A2FJWwkvKzf3EHqAg7iBQSzU6bMlL8j0vV
WNLLCyhJ/VsLhH6aRIr4th1Gf8xwTOugaV4R99eDE3zJZYuTbgiKBknHQDmaRMJ4
Nugdb+8nKnj0UnhQJuC0L8wOsLE0CvDx9H7tM60n2gjUd7Cb5/cUuZLuEIn6+xFM
ItWudPTVUtHvZ6QwYI4gyr9GWFxc5GUH/0lZfRMo8ap/uQghuXr7Lc7pM9P8lXRM
NIHnv/lkuHOdGhv+g22L3oSX2UKG7kF/x68usZxc0CFU4h/xJFpFP8lt3t6EB0Ao
x2+D8vd/54oOuM0/DWME1g8iK+FJOCRg0An7uRYlkQ8z9kXNyVoIQj6ANVgsgemv
Pl27WVGa6Sc+DPunmqQ7TiKWbfTfTF9P8GZrNX6RVaTAnkL1yKLNiafwaJEdzwO4
DQG+qIR95avUYrnC47Pwl5lvHrwtJDzSHvAEJWgAW1BZMYuqIsS1y2hQcENnD0Wm
/z9FHb+kUxgJtyeIK/g9S3AzAXhwXUYbX8biQJWm3dASvx0eoQEQOHb45bHny3yY
QIdO6a/zTd14dBArPbrtjgYRqY4jGPOdBB25pbXxLf8mvMl6xdyEl8AHUUxEjPeL
aw48VlD5qri66o37S4/xrC68hFn60tNU/P4+fCR0IEd16jSColEqrx4GGjRkt19l
FV2p7zzZaCGv7HFvt1+R5ZbomCk5VfCF/UiSEOzNAvimiI2xvyoFGhkzJX5++QHb
z8CyrbuFvDzWyMxhCMxbkQFvaumkHFwOEPT58mdzeRT+usTBUuNKiSiE5xtzgX+c
IJcMtx7Us5EA1QL1cZsQw4eXSp06gRBw3ZFS06Ieb6prBnr9YHngrW/pHouPm4zX
DIMdBWNgMpwPDRKyEFst8mUX0pfeY0hGkxcwrWIf8uWSta0ggfboVwrUd3NJUzik
Dskm21cc6srheNAeHDiN3TIvTB/WVTE/C3D/8atpf30v9z8Cglt6M54WODWShd1+
PnMlcOu3nm/jJTsQOKOEk+tvEORr196t1DbsDuTC16E2hd09ToHCyTj38ZZrPgl+
WJ7frN+oASmLZQ3gvgP8iQLDmJvAf9hwMKi2pK5FnE57N/bjLno/6edfR5wnicZQ
aGxaLBsO8dAGbWLLTWAImoMA0l5QrZqBGMVuqs6uBfFsAVWo9w8QkHnUGNGjixNZ
496gDuAp36A1OrE3opgZg0YxcnngHODhEBSlNuFNSgE5tOczTiken8mtZe++R2hQ
0w1lLYEy6OYzGAPa1KWy6kXZ0Q/2ToNOQ+BK+vmWk8nMlBqis+vKKOIikpUsxkPJ
ElUPGmCMEPClVaOAX6fyvevSCflI6KuMM8oD+za+vaPl65VHqNJcaOa/pEIeZjhe
lfYLQLHL82AoZxW8t9wd8Baj/jJm9VFykzPYh+AMHHHSBH6aTN2HJBSsvHqaoGCu
im4UVjAbmw5C/05+NuTj+ux0MJxPuXhP99YOUpIROigE85bwZ9TXIePGPIx6/Yef
RlzNnRnJededG+D9LdItS5KHXl3wFY58On0CWg7/zIT6mZYa3B+xXjwqoxizkf09
hUr6uIC3oab2tNFuf0QS1ueUnBpD9CKJqqAzqSKZPDi1oVCPubQhkks+8PXKIA7H
M3VOLDtLa/YZ96Rx0zh3H5yigsGyJGXQoCywN7RTfx3Qh9z6yyI7z60qCYcQvLpO
hKd+JenFSxTyuzypBRn7ejrmuA8WQE/6je5H2UtwUZjvSw7H0tEacyB+k49JOZ/l
3NBu6SAiKtDfVAG1Fiwd6EXCEhX3D4UZi46RYSqjwnecBVf2MD4ufDJP4WwO2TnN
x0sFKbhgRW6oBHE1hlxt44s46WDAbwv22F3Vh4F0iMNitpj+NaW3Huh8dcsj606w
CpDan4jOKhj71sQn6OpL6k3OfmGIMmNB0gftKekt0V3eTv0ODDqaXv+k//isj/6X
+p/PJ4/VwiNmtDURzMJ8g2b+SxZ1a29C7QYAmQbwtWk1+MTiLwgwVNVG9JjwNs0t
Dw0L6prwyh2ucYH0BrjLN5olFvDJN7mmzlCf48+ZiHFVEmfY0fOOacXgv71NyFW4
1A9WYsfapXJ05TExKyY1HPJ0kMqdQvZ+0IyqN/6gIN2Rc0rCWqPn21X3/gpWHq1j
MY2W9s8llJHkRTAVFZpM9O57WC79OnD4j/sV9soq680WSEFqriNHd2vZmlAOifXY
/vPxjzydQUHd6kNVeTTvVgfoQ0dHYUQjhW/V4cUwOhraqLPI3hUdtUTPu189m7EX
cHMQ1FZ5XKVD3qEGJvUpD0BIJyO7iodXqfX/jRO97DU/VzPRq6A89UBlKOqtqUTG
4w0bWE0z3VqUTPByhrDq9Cs3+ervnJouTuPyzN8Sa5oyckEDk3tvINjDzHbeF/+g
DLrkShILis8MUFZzDVeaJPjSH1kyUkEv2+PefCgO9lJ4AwEhhvQ5uT6L7CkEMmcF
JL+q+T6Aw2yl1B0FrDW2/PkvXIls//CWxb9gjF/jwuabkBO3X3rMbAtU9Z9CwxBw
WNusGlLdZ9h8TRLr65Q6tFWYdASVuCgYe/QPnqtumGmDXO01s8+owRrRBFtxZh0H
+kpj/VMJDmbriHvQLYToZOTTFLzcG1iNo/SC5q43VRqwx+LZMuizbRpVA4sRn535
tE7MmFSIN9o8S6z5plDdncu+0E5wm81h1U/g6faOXqgHJvCLfebnCL/r3j4B4y+K
0fCwtryqoFNOdNORa/Ma++hRGANvPehjIO7zk/hJ/Z4olwO/C/9mxu8wPdr3Pg+W
yEFKapPuQxKjf/HuBkXF4PR9S3ViqBli8/L5KLCwWhVCOoJTH/W9ECynJrb2K46P
siskLtMMcuMLn/bGaIj7RnupO5eYKzZ1ipBD4LotvgPpEMiNZubxUakC2nYtU/cq
Wuk1q82GEA4fcy2hUgDgWH4z7gstywh54SzDjIViFim6hnLs4PjJxmlUvzqUiNu0
1d/8r7yc6GgYASuEvPKAgQ4ngCJXkTDAr7P9OTM7TM8iMR1SUJzEGFGKgYCLYiz6
gAzhSchke8NE4PcRfZa+HCMcL2jeLHAS55aLel6ZCkpAncTDWACN7p30vR6MC71c
yw0szRzzG9rdJW/yVSZdx7svhyRlWTKZo76/86JS/LPtoG2Jn6mEk75WM0C30L9e
LFzIt+M5v9ZLrbvu+e34VOGrhXezNgeEp3mkxGF0aL/7mmLmtAMItLnuxXWOllpa
KbmchZ4ccJvRmoqE9vkOjLhqzoe0AQaeFHmLIG5zIqtj/1cs86zCBA08mk9v1TX4
kK/Fl6oOdByOd5St3qTXZtumxxJ2WdyzZC9zS3L0LfXx8ie9AHlpbxCDbDpAst46
SAGcEF4mSqmaJFVb9TMKcubZeg1OHQ9z3zE9L7SDnYogs1mr9v1YXTFRyeK7T5oN
XO2+eClkpenUNX5f3QnCT4J6cNHIwfsbwgB+JusP02xSMqD7AqwYwc7gOmwe91ik
R/ohKv8hy2h04OFw25zRmn2zyLC/RU+M1BagZFdzGUlKyDseEceCUZKmfAIKkdNc
o+rw6c6prwq0R4Lmy7JL6wUjnvfqS0QP8oa7+fdoZD3A29nKZU079ER2JCmem1T1
XlxXGPQbgqXPc/HBNh6F2FZF1gkAChNWGXFPQlnOM9lJmUL02DrAOoVzCiKHEBOe
62XeBoQMcVLiYunmGhtRAERtJONfX5nK8l1/pvkCXpHVpRu6T8o/0wfi1OHVmhxp
2iv0RJq6LMYvdI2OFzTL4z6i77WGkgWitPgXYGu5M6USZzxbj9VQIqusKjG+RQ6M
hZXpWMRqMdj4AD+B7vP93nzfyLM6fPvbZ4cTHMObU1T7jH5paass4YD8vY6Jtzcr
4ed+JmvWrkzPE3Vcc4RsoXwz+KabJDZF4aiaVkrJOkAUyWgueuqIGNiVrT2CACYZ
Ezlzr3EqQ7P27x0ZJ7ff1eQc2AJ2bMWq3oNKlqjyJH1lGcKfjtNShyILylhRoXqD
3zEhq/jkCT6d6v3YmWi2zcxyAQYRn+RdhzjRlCZ7ci5nQ/LA125AZ4VBuE7Bl7NG
EszJEo5V4nwJaxWWHRWrLLYMRKlGIqkBjwLu0l1aP/oFCvnnXhNNG5x00zjwiSnF
zTQUk78jD+qxDKUWQ/5sgBLv9tjei8q0YvkyHmTHA8l22/sR/yt7yZTFnCVqASYh
eI/2H2HxuU0/H7YpnfmgwIIVf/u/WY1eEHIafpG2l79hQRM9Cqe0OK61kgfVC+b1
zF15ETXIMuy0eHqLnF8w9v6XDxTA1c/jmmzNzcVocg0Pnay/ArrGIFphdmXIB1Po
ZvI93ZCQJrtkyxGY+wOGzcDXQEGVxCx8HOssg/nSm86BJyK/BVzf9U//ZjGUL1KZ
l4PBP53Q8BrVKDwzJElKxVEXP0En675afC2QNfn8LutvoT/pjdYfra8NdNuN24oU
M6dK2P/1NbHcFy7rEL7UYxOiw3h10krs3R5SL7r/VoY0P8Q4MFGOkEZGDZ1ykYOb
5wzOooRVjEE0azY9kx8tAJjZpcCQA0/0Wx5zCCtxCU5ZrSkf9cSwzNmiPjo1P0NV
mVcIrt47VBd0IDqkglq6YwLhXc2J2dRN4NRQGGVzJdDCCgu4CW/OFK6qlIJmIcya
mvk6gyJkgR3G6UBaiUi3mfweeKZ+Xd5KsP3gn3QAg4IqSNYnU/LTrEbLXIrbEMrk
2c48tXwVGNbb9FwY22eHtNYhwIi2eTQB4A1jLv/ltEr3OCI+mOwU/TmcPQqXwhKG
YQhzA+2m7k4qEVq4kxoH2yfrjlho4ULI9HPM/c9IeUyXdiMoaEnx92x8v5RGNdYp
w+OQrCpuMDDDb79wSg26JVd3z5jCuD/66d+LyzQq9bEdBoxns/pEFwZ3r7773dXK
JWe8bkqbGN2Z2IVLcXgDFviAZB6ESd7EGQCUhmIsYpEoLePsxLgXjaH16DuT7TfG
rXPAPSuGANnWgozq/lwKoz1qMBiJsZOcBkB3NXM1QPInCfcRGlw4Dos7ACkHLk1M
1YIDVTeB8LfDlxaZRPjhCF+0JMtIlLMXlATLRG7TZ0BlHvv8lZeXc/BS+Asu7XhZ
sfKBkartGKvObbFt+jr46jIMfpAiGRBdiib6mQcTZnQQrXd1weSiY65kR2ULjYlb
U7/2zqYRJ+qGRaZrBMCfohFq5VrcLikPlaAiKnodVfAclB/DhrHq4I0jlpMioYUT
FvlsStbwJWU3+Aq2BvSGZjEfDeXW0j1+7be6846mnm1uXI6Ho9UjUbHPJcDsCugh
vUvMGBK8mAYKQVH7mQKdAOx7D8b2luMUBoeWz/N9ReN4N/gyhAgpuKYymuwSU/zC
/3tD5gMmFJkJDiua+VPwrddBnWgsSzgx+g/dgce87sdy3iXOCt7NtAYt1Je/yd1R
+ObokHvGWI9yqxrCbX3RM2V0PPpZtewC3QZA+2mzf+Wt5BW+OqnECmW3j2kuaRAh
fh7mACBR47ha46fKkve6QRqZ0a14ruj7comh7i4FnTQ0kSAlsqUPjnDz2719k7JS
oYnPTfda/jTG3VT5HqZXAVhKTI8BikIYuzRow/io+6j3wH+jYuK7HQeAB7r5pwoz
nncct2rO43YY5PQAUYkgOuG5lmDzrgaF8ocivR2lKsyGo/02Nj4YfUZGoYJmtukE
KAFlmVueMTupiXnRZD3mK1hQeSVm0JTY4bw6Foe0oR8po3+lwprQKrdMZQ7yC28h
9W/nbRQRK1jRc2H9jHFx6GAAGiqmkZ4AXVyJ3muze0O8wiceoFS7E02hNcZ9k+Qv
VvDNiDkXfM+bId7vlJEZwXAbFl1dkLFd2X7Yv+NCubcxrgOQ/RJ8uRcn2iAoB1Xi
Xr2yicu5A4LoKT1PPLXNmQpHFzkE+GEilHRtXuLYqUueZy3JnU4SMW0k1pEcBoIF
KAFjds4Ov1zfULp/sLIGeL3/e9LTQ/IHKkwwQed78JQ2wYIXwvIDboFueQugBWnm
obF6/SpoCDNkR1o+4eWOmRXwOV3BnIlhwtd/kKFW6IvHisSS2nzX8uygRJl9UyQ3
TZobKyOrfOqKUwsQknHrsNakZXna+2+f/5rnqEwC19tGPr4d8lSg+baSSDoN+fVW
JQ4SuI195hizwHw73DlKWlWI8vlv0Kf43IueUxD7Y0FViS11Cn6uLIGICjYznhPK
T2axYVaVmWJJztsTxinYu6HVHLvsfBXKoNMRRRq294GHmVE+976EDc64+J8nPa0g
igyEzGMsZmgCRqooi3L4xiApEE1iVyOZfGXXsicOQX7UuCLOpYEzwpcGRDxZ4V42
ag7lY19kLaFXz9yU6yX9WbtTIdUErVLZkQgvEpAJvQWpa8VMchSBY4abMMvr4n3d
QgyxQChjKfnT/Ok3DsuUjbijz+h+CpkXxx0M/dvUm/x593lNqfSCNfqELyBIVWiG
+RKRaEDbCAN6+9QZczSNLtphr1z4E11OTGDLM8GsDpk5HY3hS8Vny/SXxfduXR48
kxPf01nv+ztVNCA9K8GdEVlUjhU0bkOfCld2fO8BsNI2sALdANYQa/0mwqRRj7jP
ErWlMj9K8ggAR+heSKX0j8GhEEAZJ/iB0aoX73FC5rN9umoG82OawyuGEYDtERRh
az3bxYPDW9yQ7fraV4LwtvsJ2LPBkWN6r0VXTj/0aMy/i699ZDgXQErLP7+klRHl
WCNMILI3gopAyTjtZlmVR/do28zALCIaNDWmzPUU9hBAmY8SLstocIyC6BGdVvDO
epXfx/IBU8MbSBrB5E1MTBXCHNKPciX2FbC7IVcTspB88NLrRdlVoKGevPwavUu4
oFvGA/3oTP+iaWBA5gF0krAUGDjvKyE1z5ybk05U0bzxGCF4uABBOxaDs3csNSDD
HrVuUeBdW7Ttpk+b+YLJmecUu7nUjaXeceO79MT63VvzSwimia1HlIHu+256K7I9
gUm8IsC9UPcoZ/sS449HXIl1/RL4N49kf6mWFwsiFRgLcxaYOi+ksdGITY42ds/X
1W0/Bg/UVE78FZnohAQt873No7Sesx17tpcfnTMx65bexkqyU2Zeqk+pYv5S+xkN
Konknn3YcVb5eipQ+La1hqq64W/8fI9BHS5eEr3Wq7USBg5/8tV6skuPCAtaXG9M
EI/lCBUUmu+vpeifkjRJ690z5NCIqD7PymKfS1t1T/5YkEc/RvAS/6k0xdmvOk1r
Y24CvxDN70yTBAnQ9aG4Oc/Vlj8m/py4upvXzKfJ1KhKj6yVaV5Ffmdqau2nyJhR
TAHagaZTHQ+S282la27Uxz/lwZeu3y7GeEy9Z+zXBGBv36RMkoT1jn/vVUTaFWOS
0BWL6lWDx5h7KpGU3J6rqenYwE3Xp/O4XoYuAB08NVT73WhCtBZwH1RYvb/NTMvt
WJBwaX1ZPNHWyY5EH3KfiUKGYUhFkPqcbeNGAGwT3Uxw8RHIlv1cZ1UmzwLy5bUE
DIiRX4RJV3hHfIaO712h9lgQcnZcmbrLFTWtUEhz3oCCmHLhblqV+vLRtjuFfXFi
fYIzTAmwpS4wIRtNWQoLJku3W1+bonDXcsVgrcSlpwLOC0q4teBQ5h8FEO39fc53
kslNA/ww4c6lAg7QTn9Kw/k6iN5+1wRdkG1V4e6oUu/ckDcgUHCW8LrOiNOx8wpC
3z1BAYJZroCCQIw7Lnr2BGueNkmdH3XPGcWjDE8AcXdR733m1Id7O1FBkm73E7c6
5I/vE+j62y1BLw6J8ZC43gEys3v5cGPtNxtMHsMrQuCiqsUtsCRZQ33kV10SUgwt
4xZJJFAXznCoXHTV7LQHtaryxfjqaJEZgsFlAc7uFcUWMwrd4QHY/aBKurkgmirp
8MhUYlPengnWqrAPPO/4bZcXBV1PhyD2PXLB4RYwRdFGc35m5pskcgbxXgAqa8na
VHlMlXlOl8UVNfzRSEPo+ARC3Ui66pTWofe5AyV1aQPGjIzAYrP7z3J6rJlOaY4u
sJJXqrfYK9heAZIK2TTy277drQw++7UWuGp6Y79e3eNzxAsEM3vd33IlR53rqDAD
F1VrlVl+LmuyYlsWrd3TrX9yqQ97cH8Efsz9Gg2O/oAclpF+O543JXGwfxwTOG1t
aBTfHePc78r8un6OnAZ04UwjDX6DpLorgcDFgmF7+1+OdxoPc4cZYaDVbBpKVXO1
XbLQ6pvY+ghShH//NJiN0adxNoI1BCuE4u9ry5Io7tQHM7iKSi/NcOdJaCNDRCt3
VVGDDSfRmSqsF5iLK/EaNy5ywsGWcGF5m5C5GYt9Vzhh9iF4kBEXu+gKuObDFSHo
vq+COhz2Wdvnl3OYUbXMi/PaaihKW4h4u76P8xO8lRv7m1fbQh+Qb5/bYui15fle
n5X7NTz5a8R4tJU/+lNVECI5Qv34WWLh+F/kuONxrvLRFo7OLrr7lySPA+UuShtj
DI0aFVMmIzXoA9D4pj5/b4c7DCC0lbnH0rRnFL3g1m/PbCVORtzSbr/Y3IK8jH/b
as2/NLyTnQphJOgVTBQAQVkcl5c7LVU2QV+SZxTrMUpbyvJArkFkmzKIswpjBkdV
o1XkxAm8RcqMJ6tqyomv0MbE2TKVDTTsqYk2v0N0KA/nm5CKDnO1Tl9agVltoFBg
Q3PnqhsP+CEw9Y3hwXbf/EynjMd6I7BQ3huE/BjyQARvxEfX/dnptRVmZq6dQFFz
nws1ulkqQnGiwSdzIRA2Vq7LDNaDvkn6Ugprbt/xByX9XZ1HJ6ekuHY9z12vrRk7
3Aikfkkrvv8GuhZ7TdewL90Tw19EW9cpKti2Hdx2wMed7V0IXyr2s0yVAwKL6mnq
MM7IK1asE3LbScPSDRUxWdKTrbYFf7Q+bEDy9Rkf/QqTgI4KJeI2znLu7Sjbn+vC
8H2CV3MYXBsqBKuy5h6VOS9MvRFAdarY2mWDz9pA69bF6vmMOoUczsML1AURTmo1
ZsgiPi7Zae1KEjTWU+LcjyV8om4DW7R56oNz8iS3/pMFKx6tkBSxzyEMTby/eYNV
tgbyy28n8XReYVfE8MQmrxZcyQO+DB8Mzhd987FS7dD1ny0z+3MJGYUPNHIJcEEI
UDnbRiHa7HPtdd0+hEPp73hztWtCVKTVjVDbJ0Wr82zbCSheXvfbm/lNtMVM0+TA
QrANrvVFOivagGwPAIhuMALUy9luWMOAJvvZPfmmDKK087dZ57HaZcQ4fMTYd8fF
iRTj0ytbv/zfel5THvB+Mt4pjAu4ert93zjrJObaS6f6JRFpX4XbfUnXwTy2LF7s
+SNNaaAmB8yU1bba/K3pisecDnbgo4Y2nPrfaV0TLenVXge5h+VHVBijT+MIsoLj
mXfA1UseNue5RUA5jqR1ZgGHzsMMfGzZCrdF/tXrE7y1+NwEAx+DFQIofHGmT6I5
92vgeaO4pq9pRxRGE9LgyS63yn51vMQH39HivESpu5vozswDZtrMDpSiG3HrnayB
dH6jQ4+lCiWAuAc7gpSn1cJFzfndBd8mQHnqT3MoDuuIfEtVggIoktpKIu1/bqoe
LOGKglTb4k9pE8E95oTpxFSteH3KEOH3PW9MOVLg1JRUE98tE935qs1ZkVkAochg
fx31/HRif8yd8849eJVQrzSFtU+KF5wUheni5oUGzSnlyAGNd263yrP0v1VMwFJY
RNElO4XpoitKDdbTnU0ToeYcDYxN55elXG0IiuFQeQ9lOYfciVQrkObAw59d/dGy
3USysYlcxPYqKaavRw90INwHvj6OIm/PGwuRxptf5pTpeMLzGccYUSEOjHQpkD9E
iCfCF3ZrIl55vTEFECwJvIFETGcGglccnycm4DfDQIU4a/U9LmagNdSqWfjZGtPG
sxWyLIpkRC5X/9g7kGz7LIXuUAZ1JeOYTUfhETlsICoToDsvg5Rg6dY3DP6IwBxx
C8tIuDPIVj0k/PYh86ly8JQckWqJhyToj6VumHWfQEv2uMEwZmdlhCrdzArv9PDa
USH/iRLGipkhsCblXeW8ZVahoEJt0a9WAIyMRnfe2e01fxsXRn5fBkO/CGyE3wPY
zlb6Xusu8OaRBOdgm6BM4qOL94Sb2cmOay1J0IgBGxhGH1oCAEkL+nnFMw4TPMUs
GatlE3iDb0HY4NlSh1SjwfCo7MPvSulVOVTZyL8MFnEuDww5RE0nQN8zE0NS6dBi
81gp79g6VIm8cZZwsF+KUKgOmKr3/WfjuuSoDIC8cHG1q4cHuglTS9K3cOOA9Gwl
NYoX967TUIHBr5b66vObmo2M6+dtZ4BEeFfUlAU6JuwLOI34WcUscuQPLbxQc2R/
bpkZQnFgB8FO0kD07ZUcg5YBunNvNP/g4bnza+3Dts84mdxpBmZD2BLVN9EaC+Qd
kxMed4+lCuQf0WQ9SSmwGnGaWLYd+sh4xGNl4g8kVvEcT96OZjOT+Mmnp0SR+fg4
tEwPxuo1xcUeZm3SfpMmYCCo97uPG7gnjk/8nESJQR/Atg6QaN0fGWvDOi9LCN6d
IoPMpW+r0fQPPnr2o6IwQjiP+m13FA0+nAjvoue5NFMnYcjccD9sVX+lqT5+Uiui
DAz0BOAZRVLzqkdpEBJi7yOQFNqXhfr6Cui/zYjGxRSJ3HMmDrZchV6bs4lCGmme
KI8epB0utfwDO1h/XlSuGk1XaWTcFxBt+5lzLblZALRjhgYHiAwCnebBFVxcphWE
QANrBMdKdEQZdUpXQ6+cIyvLDFiQ2NiUDvFjKmeaam76iQ2AVdlcfl13KN79h155
gdVERu+HQFgH+QKFI8Ut68BGfqr9mWcgqirjifBgZlYtYiz1SLO66tsNZPpPtdh2
pHdYhWPYwdOPX+5N3osP0gACePon/HsQDk98WBELq84K6y4pHJbUCMKXjIn8/AmH
NiId066XijgtJwIFvXFiq6gfnk6jat6W1oOgWpVgNlg8powsMQK3/9RmC/uEOjHp
fLU52keHgN5Z4Iq2GzRkFJZuLPISj3DxUPFMKCg0z5XKV6LTzL7Yd1x97gAa8WvU
zeJ1Spn+P7cXv0H3VARtK0Lj8FiEbNk0rA8SKR0gqiWHdFBPIkdoc5WG/e377k9S
fSlVBv/S/muWRagx7IPYW2WnzhVNx8PBc5swRslRcpsQTox//vAzzISko+ISdymo
ff53sCW0NZWX056i+/N62zk44+KgByJG+UxKq+N3TWsR9K0WSuspaPOemV0uo1jx
OhkX+NxjyjWsCQ7NmjFPFIQMoTy0FGzmVokNl491Rxfkk4mioiz/skavXog6/7DA
GT0GZkopwz4saAvilAtr3w7JTo6CBbLb/Opm5ssft/EguOA0ZJRuULCNkhFy0fKE
NTwAd2Pn+NokllKZTmNtjEublbMKUTGOn/LB2k1NjOVcaySmzwbWal13JJ9yMboq
F5YZWTuN2UrPYb80jskNbKW/tWK6lLTr3FDCZQ3c0cTp2317+7DxGjRjGF7DiOYA
BfQFGeTiu/uh8YwwA+ZS5tkK9v4pgt6gs5OSoL2eDNs6QohwFpTKhKNrJEeyWGdK
XNhtTXdcsVTc4VCIuF2KJsj+5MIfwYozfSxuF3h+MXqWQsGN9bxbBR4rmMBK5g1B
lsXvqzos6SC7GWZMefOPFDO5vQQ5WP/MMzvjQW3yTSWe1/QVYqDW5AIwZtX/USyj
SrfV0xLqKDmYqioYSNl4gj6dL40TYckrKH08J1iTct8KR1RWu2Czbyt1TuDuqPmg
kxdpseBTYzNz0qUaRXYPDVApV94fISXNZWYrg+L4FUQGau7tqA1gnPyYezTjX8QO
NZMeyYJmbJL7TUhXzKzCmsj0iZLh/nRDhxQ2z78AvosbC0lV91G2NFAoN7rEA+KX
LrzS3fPwq/GCPDQG+l1im659w14HDAyNvg9pEA7gujWyqQpy52Xzzh6RbGHObSQs
sB0q5z9ZFOxO8F/ww/eQ4OVUGah4d07YBRmmVT4zVQ0ovcDG9YfcAX9e21+7SOQQ
4uKIZ7IUvxoZt2Q5F4EDw9l5IEusOvXlWqJLXiPYXMjiO0p/AXgKbhFW5nuWXwlX
zz+DUs4LQZffXYfZwuHZcDCPsVTub+VePSp/Z5OlA9z8DSghTGgHk143RqsORpdg
I3kJ8ISNJ/YlBWtRjNa6VX8aGbeyhYPjwMG2CK0j/HepLas+K7MD7jEZBnIZr+ag
weNXO8tRgTFW8VyKZurbqSh5CTz/10xJzY4GX1wKIT3IFSPnMZ7PFDHUttsJ1HXf
5+k26Glvd1TEVVNGO7NzfXB9mWTjcqtE7Y3VFlrMlhGnSCDxqwkzKVu1SdzSuADf
MbC94HOtjeGRtfI6PtRKD4cBwrlzcZHX/oulnCm2fWlpm583BNNFdW0DDS5zxQqc
NY/hl0H4fwTQNWlXiLLI55xyY6Ufk584ZxalePbzQLU5FHH40PkHoLoTV77Hbz3Y
dlKXOxtKqhsqT8WNVOw5s8tA7SqkoAdfCn9CN9FkzWgwJN4lvTlHvqCa9L/pGAku
AVa7qFt3N0H6qcriviCY3sG9xsfE1D/3EbUPTrufv2RykS/70EztTXgcld8xApNq
70PTtGtaCF3e1BQU37CSrcQi5R/8nPtsAzlFxmX6QFL6DIVV9yLyKAvzu7A250ss
XsoOL/F4rwRbZFRfi4Y9bI3WOsmnrkpWlGPc12EH12OYAcCus/zOgoGDz+vS8Ofi
6eZMJ6s/yXGLtQ/dofBBt+BeqlYgyce0Fsaa8AocGs2gQ2ueoE0KX+emJL3a0Mb6
3nw3dot605XpA3AkbxiTSfDiFV4+LVB2WdsFa8xKO34p7/jAStQHReb7F9PAVUQ9
pyy37/ToLHlalqRj0vR4GGS/ubBng2p5b2oKdScQSv0PmT1rR8IV4+wQnNRY7+G+
vQeoEoG5U7UK8m/VUlmQX6X+C+eRIpbWlHJf8safIQyzLv+xlGb2vFIpFgm4faBt
ZE44YU0Ugz588ZjC1IIkJJRdLIPdthXNDpRU08XuD4Lrow8weHi+yeGmbWtrP02l
51ifJ9YgUc6uX24Suci9oRdxKW2vqQgrlrY75VkoAX7rpS/c+anK/d4ZYhx4BpJW
qmUNmap2mecpD6zAcHYNuLxyZJr1k5fYrW5BpsdHedEPqQ+gYUyFG5DZhceDRF3k
hfOxNL4h0G1A8Gp47k17ht8WcbsI/cgpzXveAfKA/NQa1TOILJkZnO07DpsurV1t
SJdJeqQJmdA8w25pAxfafzp5d6AIriigbp+tYHt+jraUy10Tviuptd4V2nFuH0HZ
KEMbGX5HqNHrjiIxR1jOB/13ffdBb8FlrODuIHYN+QJ4tzG6l9s7lJI4VjU1kMLC
BcgNT/Ozxe/kTPrQ3DYGaSPWwLimVFJsdiZnFjbu4FEtRcnaKb3VVniJjIwQHYyo
u0ZMY0FmFlfh3LtpjgmXcaXwEJZZSiOP/8MnbS6DuzUu/VJL0GG/sl4G+xnlf0XK
oUmsM6OGfSMsliYm6lQNSaHbAb4SQrLWtHlNio60vpPhHPK5mQ8xYID29zrvzAPh
zPwyjFJVagMV9T1Pxv+tUZCzSY3B2Vylcxgwa2SOITaBQeYlbB8OQrkr7G4Ljw17
0QJbvCpWT7qa6ieKyiDG+2wUidpIn+FZEmaEkGH47gthwNCSHd04RCbfjXYjuIlO
M9OoECF3mMOsYnwj8gaxdYp2XnmUIYZlcOxeaHfwudixph9RiNjAEzwD9Wm4gDpz
ArofTjBEsD4Mzxk7t4tZmqPTpxLJTdYQEppJ9/gMz4jgOikHYXNj9z7h5QYeCZOY
NVLy8VZ6Ec+hxaQKZlbsSqhF9bwaKj5851rncaDtG2JZGCxngpKO/pXr0zvxb3pQ
hoOT82IkilbHGnm7xN/n4AtjL9vKJgWXgPNgXLm52kMQo47qFaJwPVFiplekwuOR
RMMx3hU09ZyU0tOBfFpDzatFenLEZnmxLItBP1a5tx2hi1887DhqD1KTibOUtYMX
OLZjWNHeZIjGCkgIq/0jeVPiE7qwYwhZQS2Q4+/carQf2XVyXqIgl77tyQ6OJ/wY
p4ueY/xU7eJ2EdIMtPy6cAg4bptDvhjLStyIYslLNwel+betqmU7Xybfgh7Jt1eN
1CcdKCoC42Eiiitda8HgYm+kZi/LV/XHe1EhgDKCDNC5kXuRFzg6gICjfhA2lVc5
zLCwi7mPM7D6pX4UGGdya3s7Xw7y/w8in3bMjF/4SAxrFwY1ZXN48jl8cb0PYH32
Egdyd6rSDkLsxothssx171OExzOHebjb5IE0arSHac8dkILZIdF8EyKRZjuF7em/
eWNGN+GGQRJ+9SFjd2fZDeXPFhi0cW9HbRG/9MaJqBQSopvstneh1x55ahJAc44s
+39WPnEDZ5gMrqbHA728RZk044NQxJefiHW/8Ki8VNyljTOjMVA+1nwW8oj4T9qN
6tZSGGb40cLAOtvo7qZsP7sZCDtCBMISsF9MdJ7WtlilCcXqcM8PUIJPvZzi2l4O
/TBzQR3CEy4zKvjXyMmc6NRvMwkfdhuyBrs3kKJ8zcDQD9OsVoM89ywtQEhj5HWV
b98rjYp7rJF7D0nTA7VE2Q==
`pragma protect end_protected
