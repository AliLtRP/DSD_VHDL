// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:13 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hRSJYEMpm/HOUBJNHKdsI+VD4FmfXQqt9ScMq88wU8o7z7oEjw1r8bjrtkhvL/0V
PmkmYBGh1rE0dZqr9ErgOr38ZtupGfnaq8okiCHg65ZPEGTeF9pY4DHF4Nxaqxnf
motp3w8P87oauUFggH511qBddqYAZekUtYY3hwvhJRk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13648)
ZoB17HsAKCy+ZSH9O7BvB5/ZmUKnCAcigi1atPO7hHIyVq3qqjFJEhFH13+WNNJd
m/TV8/8rhSmqASxxzGubAoIuadFEXzGLN9gYggWicqhkgaJdhTQAeb31THl2Lg5j
c25sUVO7845rKNGrOUOC/+lbo1yWWr+Bg4r2bWy16n1NKHErrUP2wvWtissenObz
bUHvMtqqg/I/VJaozII2FGUBSaSLMFv2q2ZqtrqPdv7Csg/+exVnr2UVAFAatMT5
+GWHXcXwJD0NHvzjVvKdDPVAjn6QZF/J23AcpwLKdYT8J5jwjMObc+ZgjeMQKzFl
8XetjjyPz6+8dTKYzoN6TBnfMm+b1HHfdhC/qqzIV11pwqaU5iMENVVKx05MTxT9
HUoriso77cp9eb6SYPlnvDsoEpw2Y3mc9vylzTsMzM0l+4tPqajN28oMP279nktn
RAfMlgZEoObSHoaziYjZ5djfx1ymtPrJGiTj2CjuDReAksEx+BZNeSxtLQTjYqt2
+hfAXdeg8lwVbttFy07o1//OFUT31IL2TfoKBkjQUYmO8ajIDYDmF3BV8zLev3a5
34I+FKThOS2jY5UUR4go3+Opfxkatk8WhF22JC+uxW2MyHqTq9npuXJ1m1KzmUP9
KrBc3Mm+odNm/yelxphKGficZvLRzbO9GwXDVFkHv/I/XKD2tJQaMMfKEYB75EW2
dTZai4E76T5u9fU3l3wrvEmB1EyXMisAY6qQ6Sa+xEMNUWF3X1smDVZd0sMlzjLh
OaeQrqUPPyi7tV76hzmY3KEMllsgilw/kiXnYVVgd60pyZpC51nUaGa32nYUxgxH
tVQT7XZCpb/lnKPmoh0jON4lkOKXmMsegwM77GBmQCj8kkB06/7/HHKzwtCRhmJb
4wUaliMUtFzZBXbywvZnxEkl0A212W7N5DkkkjOEtMy41nH7j9Uz3Zup2xpTdpRw
DkAiT8mQ/ZT4ciJnosLMAtI0MtI9ql4OUOlNDoYGTr7hUXD20t6zFhr2FHr3V7Dq
qFkV5jjvyou6no36TXTDJ/WqlgctDYNTOVNQpLpPWCY0lso6eiR+c/JCU/FbuWd+
O4tZ/CbvtvS1ECe4vkoU7Pp72YaCihP53mYPq5eeF1OHdxNo3uKyLEPV0Cv4Hz+C
mVopnIed4ughqRj/76z+6nSyYqBJTE13lqzDTCk/0CkLZArEm3bDejJcH+9kII09
1Z2wU3qjn29VNVIs9KwdnCqxLdq5GMbX3HWXyndegV2mzjhJ0B6NF20AjN8gIEoJ
YIopjtg0oN60cP6505fCOe9S1FePV/s/B027UTzkUQitR2TNNcJsoQbBkcnShQ3p
tdCLG0OvczTk5BDL/UwM7hk80veKZ0av5dd+WmJ9oQVVEV+QpkuI1/KmazegWVBS
/pZT73fm2LO4p8sRJckikO2NYF/ybyfMhTSQqeGnDRa+YW728+wqA+602+GoRw57
SdFiHiwIdGV2aMIpXYN0S5aN0DnoMwiNpadw8VzzZlYEv0WmVZKleDf+BfUvA+RZ
IyqdOdOODtXeA0hGdjDm3EYbiJgdIotAah8N+DkBS90NWaajaxLdzcxbE8AQgrmy
9GJDPXgknbk3Sb/D5/qtBSDfvt9aBKA1618X93op5j8wp0a433BqWDVdVZGAibOK
K4+ntWMtPDBJL4Y5KZBn9AMDi75hvKhiVmYH6GmUkWk9hA2udwQZUDaozCdRNN5k
M7CQLrLr2V+sY8srEk/bo30mzMVk0dfSZYTGDXljTLbKV7rJUO38Kzpc8CIzaOF1
ASetjN/cuv92GmlRAdIjtfbHhbMmTLyCrtYJUwJ5GSaJqRh3ygm0RWj1zmGRa7Rk
zzKh9u3yeqm/tAQv7MxR4tN+eTIyiLDinkxwFv1JADKYnir7jq0/1jIz/n0mkJoc
F+M6PCT4cGxBXVyd/JrUX3ssi0PONPUSA5kemqPtE5V411m0O2DFo/70sm6sWv7+
P/3FTLOInVGcEeItiBE4Luyh1NHnsnHO5PD+jrVpPWZX4XFRM5dp1lJmLDsgtdH0
eFAifLLDdDxmnzY4dMByXxJVtO2FxNQN3y1T1SZAQQ6oCxh73sz6P/RndBujkejX
oL48dLQtMC13PNk5rG9b1+K6J253DFIk4HxfH5Swz20qT/zsaOOuIcl5PC/1HfxH
rlJiaPAKSYq1qLDVqYNVhZCWm+Hi6hs/TMtnMIwa0YDK2xamvJ+xuFF+dJi+6bWs
tH4OxpuY2IsCtOa7re+Em7iHP9eInXuEqm+H4QQW4030x2yH8dsLHm0wFYrrozoh
v+g2im6nfwcj8dGOcXV3apo+U+Qu05r0qcabhUeLWHnTqJRGGRW6ce20Rb8UkE94
A+1MoSOYDfM+ZsCxrbv272JlhUheKltK92ZSIqqzQOWHEcwnuywwLU3cWLjeSWPe
ikuJF6M5MI3vEdJfoihlVYIPTMIyoU+Q1jxvV92A6FuYOCRHC39Vk9ATqdtxUBxo
JUABhywH5qIZ/tyhWqFQZ7TpMTT4B6kGI6zYRTUoJHXOr0w12e7LWBiUdd5DxjIJ
LWYrRMvmJqdshJixeLPJ23ouxCMJX8bbp4N1RfsxLy/ia+62c9/sq/7IQ1TIX7+d
KeIu0nHyxOd0AUQ3mQtkETowxzXwOCqWNbPqJKZufJ2Qe91nKiWhh/QK/5ZT7Dt8
4n9gQCi2iasQZ+f7nG71QXXzy+tExptYIAAk6ljDlVd5OZYhkt9odz1WsfVJ8fHu
vSeGBcxz1bBC2d++VBEfJ6pZLUgw3LBUQ8idAwt15F3m3RyaVwmCht683KQ1wTKQ
KYyohA1ymTjzoVuCtHTB+2dWXBbVrpC9V5fAFg/pHpbLUFQqyaN2FUOKKBey8BmX
bR31t2wV8hNjHFAw5dXO8NdQh8Nfnij/fvPC+CZgnFYhprG2wi/nyJdPG99ZWqbD
j55X+Hn7aZR5aexmicTf/fIEmfyczo+KDsO5+e4RfCXNcxKHTCE86CT1AAJGMvNx
1l4NuyGTDwPTL9f+gDmmla4NZmyqZOr4LpS7jy6IQw77CBjKdu6u4RU/X4sWl6zD
Bx6vqbUByYLTVn2sQqEXXKJzCc5c850sVvt97Vd2YsiRRqhnpnIFGkFWGllXsXKi
bnmYsXFTRc8P/RYFZhkD9PGS+etdNz+28YrUx4FwKipLBNW8T0PvhK3LaGfyM1zs
VSmEto6o83/GD4hsnSKR+tMf8cHcimg7bJQ9gsgs/aVdYL9pCz8DoILxqDssWx1Q
SycyRHOb4f5gqPRZsI00EtmyWopQazB0kjm6Mrnu1VoJZXHVrVrPR3HSFCpGA3gE
3fyNValbdaspWq2cDxb9368ViC6RBCRAXcGJa0YJhvbIUkyUda2TWD35Z+d9FQvN
Btg61MOfNsJvKQ2nLcWkTdiaiD3GdRcpkNpylowP92f/9UeJppWqS7MialZACApg
0dEwlWyyqYIv1zAeMHwRrdVtCi849rrk6eDgh3Rab2P+0bZyEhAI9I9RLiF2VCoR
etzXvhb55ZIlsTunf9EHCdItmj+Stx8Io8f/FzfA3G/R/mrN3E8yg/tbyqLiD411
hAwzcSKg6wpo6RO+vWwQnCQDp+CmklqOP6HJ2NiejS2T4gZJOzLAChzTkoemTjdW
V2wKt5irEbqpq1I9+ppJ/V1gW/9Wrv8l+HPPDcJ9EMF1ekinJKJVyeFfZk0S0jFL
vLjbcjetOM19kT/bkuGgUjiwh4cnYXiFXkTNL4yWT7ojWW0hWEuC2C9b1JA+XxKE
6EDZW/TquWmdlxEbOj3UE2Mtl+uKPZLZuDFwjTxIeuC/COmhlX1hktN7NrfeDAqr
UyEGi4nE3frnZndRXtwmzy9n3oYDwIijUwoQXQhf8qZ8XfLzRqTkHMHiOs2uPW7L
ThJl9FB7V2LPGK1IVhFbGcvuMIObChQPXCIMwxX0yZPrGiOW332zxdIWc356tqjX
LZmyB7YlJU9qeecT55xPgY+iCpWJgedbrNedWWSBfwm5OYvt6V4DXSNVIvuQj5PB
k1lK9Qt11q/xbUfoOxK4THgxvKMUWyrZe67nfgLEIBO8x7aO1XWEkOOYzLZr0V+2
2CX2tGuvkROup2PDZaD8vWk7hGhHdpFwxAr+HJe9oFb/iehoeRUmT0o5gZDzv06j
eEDbfKqtmRfqMHbDFFeRucyvfks2Mjs0SybcKPMwmF0/c7+HF+j4u1q6MSzHMr/5
l6f51lx0IEjpTYd2Y9HNvqxdQwikSwe4t/59pN6156sfQygjJdLAaSFe4FJgnQO1
FKaHflD2Ba+AFs7TTDkANtOsEDTeKRGX85xK8zsY1dldmAKg4c136Aqxod00cx5U
amrFZXYbUMPuUVqAbvzURB+AjOf0ZIqQRXqoK9je3qQrpL/jXX3YNCkG1sDtDMI6
X8kLmm73NbxW2rRzoRD1Fv8TmSyWbi2gwa2RsQu4XMPejzX+uzXcmhv1V3Bvw4+D
V8K8+dliWb2iIRAhbgmTMDigvTrhiZ6OCZD0K9AhVMbIqZBTSen2d+R+it2TMaDM
S1EXZzSQdl4ztDwL+6k2IXiAnsdb4YfA/uJReGIBim8rBBjEiqzVmb7K/Opy0O8p
v700/VLrJfmrMIG/q01M6z17YkjGzHM3lper1R2yFO7abATWFYqS4MQDSQXVfJB2
xtZtTlz5CgLTE6+TF84FElJHnIq+LE3yUiMp0Wv9n0rBHgUF1i3hf7PCnv9OiM6W
6WmmcOuiDxW1CIEWwuc/uEKQx8EspQX1B+XVry1KHW9PBS4dAKTqDcn+QWjiFJr8
dJStCioOOPTkIi09nrfZKyzCxQBDBYYnHuWwdf0cMVBLClkxOlgwANQcRQFn1uXm
SLv4AmyIEbaYcge6dhe4T94LysS55OgeXYURG2voubPu4daZizNesv7YiNKYEsLt
MV+9BsgFbI+YHTe3zR4RZzoVaB0eHgrvS3M9KEzd9uQPhiqbVmBECI1yhOjeorNf
VvfiFqvIUtsGBTqqjyW07CNKSgepxR4DYnBAzkBKZYGqnIQqELcIeu3CI7VImESQ
lRmhegn4PCyOouOjKUong/p0mxg6NcKzu7awv1w4enXgjc0Ot6g0IyDoY51WvjT+
5bGrZTIW9IfkzN8xFOobf/rZfoNheg+4y9lyls5sEQp6rbnSF93KIZzv2s/Z7o0h
Ubr24524wa5j+83LJ8EGv29MQnzbkYE/ON6HTbrjl1YrFl1gqqzY5262BiWIAJwR
6eq/laU+nD4Mx5jCNGvPYzPSjK4DQTeWUsEa/vmebnuBUEaHFPpyvgTLal09gnGc
vkb6+hLTFyJLeuYXTr7sh5/9BpKUwAmH76ygPE/I24kT82G3J8GiOXDbthIn4ory
PJzkTn350De9NdcIVHBRPDw7HCuLPifAGKrswFrWsC65LbvAbdOoZTLZBCsVQUCj
crIzYAsJ/NddIbnqNJBwgmLb9UOE5m6d7WS7NnA4N/aZUa+0H5dNzsKeprzFzDW6
1BmRHc1nKoOd/1gBnyTgy/xMeUlZLV+UEMQcNVLel7nj7HntC3lPuOo+KbfmbKsd
PUuFDu6PvfaPzSB28tghd9L9KEMXZFNF0jm8bu+1NLY3Bj8n9g4V6lp739m6c+Xc
70Lgc+M1mivMjZRn0Kamsgd56OJ62sn0oLemgDfQCl5U1PoyNQqdVMpQG4xVFnMd
H13atRR6f3fETaOIlmzPHo0cNJyafAnugzIX9eOJCjbp7HYIrx1XVkLUHAf/ZXRh
thjUD2j1mDmg8lF685No14QWnDAKlz+sqBVLzU0qObTy4xjAVmPNVRXr5ugFSViw
Qc+bNI1R2FjZ+xD+j4FLWc4QxAh2Z7NAMLtITUpeL7b6RrQUZbQbMI9YEHu632Ny
77r2w3zksbimagIP90fyQboRIWxxysAExSRjYHdOJcCbKadXtbDQqmvT4hhTQz3m
j3fcxi+tpgXrNvEWAEEA3kML5lvjhWu38/BgQoEEwvFMdM+Gt5cPXc/m6UdD05mY
BF2amm6enBqHaXBAHOkvDykIkkcHUawkMRNh02pMseerkf1WsVoCA3EIYh79F+lj
POXxWmAPw0b2ESdgRBLHE1cAM6ENNBL5TNBT0th40kpke9bLRt/XzqPLtbPEYRO7
WdNbfX6Dl0qLdMJt3b556WcLl5tN+FiCokR1QQ3q/tt78kYlaU772037at541oAb
bUvz6kn+Mip00AOEzHhNkLTucGecvRNFVxpszOKBcn3KpVhf0287srlyFEUNJOgC
PBKhygeMoAx1BTQLa1m5MyfruRf5BhSJIEaGM5vLdDLXcaghy+1rXa6lYtgNQl7k
Cfp5V5ZWkny/1rM4ePbzEcXq3zQvAdhqe8t8wIwEKOzf2FmPwrB/m9mADFS5dG1U
QGFx3Wmkc66F7hBbb3aFbkvP+CLJN/7ZYgglSFfjjHrFC9TuyfbBxrXD7+2JaF6u
M0MOKOn3IZsyniyZRICTwkepMKruiGFtzRd1bfC+YguiBxuJI/BH9HuLjUIXsfxo
n4uO7b3f0+3bQZo77jUzFeTSHmi4Op/JL8pmqCRkaBUMxZby792fqkFBveZhzlPJ
+soJ50f0WWyiMx6XZRQuVfO5+4wtRVTWqfG6ehCGV2+jGDSy4gpsOSDp1+jlDMS0
q+Cp8sNMAPZ9ndvxBdAyckfP2p2Xn8NEc7FK1+xWOpCH6xV6dbaEcrQFC1BKkePK
xI9p+g/1Hbj4ByJLYoYsL8kvykJt9JMbug5aDd21eGKEFb2qe+zk3ekclzg4N/8S
/OZEA8PLFwJzwEIKsgdyHqwHd3pbiC4OG6AuRcGXZn7k88OMx2jcbIYfBMolcCUn
X7gxwFY1ivvRL6qmh7nLQ6PptpfBvogeCq3HpdnBWkLWZguGze3C+JHzNCLOIJhE
IubE130uCbVVr/b4hdz1iXdNkM6XQQf11Lar+y/YGY7qslOtf5pf+twvGqrMsYMe
u+yb3hsydDLV3+SMGj1Spch+XZ9E+O5cfIQulEJKsen1qIeKUIrZ99MNrAXl/022
4q1lo3XjzvRTnuxw1QnYxk2OapD8b97cUIFmGnzk5KfvlmmoM6SCwjqqMfBBxvce
lqkTdPn1PO8mU3hif4Nws3GF4R8tRGd1x033DMJrQgM8piu049tIYMSAbSjbAKUn
x3e4wXD8nUOrvGCacuGYOipKH9vV/Z5n32AoL+oTLkA6Irynp/sb020djsg5iUcs
BGq0kT5zGU3JF5FlZ/MDNcaRNrBCuBCsmYflHAZYa9q1gUrDb0Pz4OdCQt1/VTcu
vQG+0z6nn4opTvct17K/a6/vY3e6xnTTgutkX/UVbmlQCRnVbGO0ELOxW3mSUFek
zV7Hh3klKi3gf/E3HsNrv2DHyhRXn/Q6kMhPQsvCaCJqJTXNenwjFJ/tGLSYbsbb
tEPkWsD9lSXNa0iFUSx8RykBwhlxRK2Msy2yx6NsqW5dY/LpWg3ANBcp1kOMHPEv
7xwa44inf+ZxBGuBMGw+qB91WbWQquox8Opp2lytgebeq+oqhEEn4bKflpIf+mBL
q/0vnVGYvPHmul3yx7gO1ZHjV4oqnNTKD+6ii0/bEFVkyqG4+Zm309YqNfL1R0U0
FNUmhnXbmzF/6XB583v/mEFQ+nLGl8C7M5FMlsJiK9lApK2ECg2QlazT1dHsc6mz
nLltDjeOZWwTw0A1V/6UchFU8yHmEzBkEGVY0lLoNCdxbCWttjIzd+1sv56wQxsb
XJ86UAI0lJNfAViBj7avrlh4hZN6wIllclUuKWBn6wArftj/1caaied1V4up4l3D
qswibJyt+M/7e66sZ/HzstnYh21e3C63AJhYUxIJEF1ZerZYkSMeTTU78TTxbI5b
/USENSzTyZUxvJ9r4luNQfjXeJga0wbnoQS/WuQM4idjxPP9aco30LzoCs3ps290
quSFbddJ/RJIC1E5/bpGWfQgWLan2Tnoap/5OI7mWQidttuFLLuXMwOBLzwNVgEo
Oi4xBOONGKB8ISzyCiHXaGMRC0GeaBKp5zHcO6IgXdk3EmBCge9tX/aiQ8A4GU4d
Ib1aHN61alUMXl0Hem/dL/OROKGmuY0lyBmAAPk4o9XfQLq229Xe5uZVDRnSs/m1
8ZVkaDjtFR4vEjv1GbU462naDMdt6dNP9F3UMHUBiQaysRE42YlZAirZePtDQ8zZ
n4Dy3qFNkL8mFMizQZ3SYk1TTNDbzw/S3z7d20ls8I+3PWkLwRv4W5DSgxuenylZ
hx7icOOoUUBaGJjmyIPeLp15nVlaFIJyKr/RfFhDPUKeFtdyCuCEr/mUyLKyhzyT
AKDq55TLfQxJzWfdaFUlfiF5aMpb1aXWtlwPTmeY7nBLOi4bqjpz8rjfjNAzJCPW
1bx5RQkn9y3GypbtSgpCakxmktX3GpaTjNhuH/QF1UnMnKbwtMy1nyJQOUgV15oK
fP4CtTiLdkkj+X3aXnoixpGJOWCsG5iwpNy54/8ou8X3zhkUz0oKVBh/L/xO27bn
+P+lm3jC7nV7Wr2K4LWiMnOrqebhy2amUpB0f7WxgGXO7h+d21sBTbrLFjOZ7Ltw
8roc0ps17p4Gu3jzym0vUaepezRg7bt4CfaEJ6Hsh/bPjXBm4l3pG5y/0P7Xqb2l
KnHHy1J4DMZExONEvxYP84hCqm5qCug1Zp1XC6Dgyrq0Z41mt2++8PrTY44xnDBU
Gg1fzHJwlHt/D3+VetnoEqY2ZuFkD60dErdIoxmLvzq8zs9sH0bjvKoZdQE0GJ4S
ah0hyHbuRqPc0yoaIufjxbhrimSP3etg+e0vWpbvXH50QAxy66vJIojqBq7QeI66
yqkQp48VCL5FZ71clcz+9qEQHTN0rzf9kHy+AG8JClHsPlnYcLA5CVuVO3T5ynGr
hK4TPYFx+rEj54mf4jrcZsfjn+XoBpW/F0u74aGdzY5slZLAKt7F9Hk3Q9qjo+z4
KOaaIzzIhPKvgE1pieWClvI5xAG9ov2k8NBKbM1oRdjlYPt6YLoFvCySA31KCwc4
nxbIdDdRREAFldoWQ2nFPYWXRSy8Bx5tYDbFzqq4ClCHR7ACV1cz8SVBYVaExi58
PoRxv0I1xb2zD6dTa+7Fy5kgHSwTQUe2JiWG6tf2cGbPlfNHZ7bDwT75+ggT/H1Y
zG7wfjcEQs1ey0XRt45g57lbsqKBXQ3RckLzeyvKkRW2YXJwlllIDEz/WeLV1UZD
9SdZvBFNXUxzMA/yVQ1s92OZ3JFX+mLekCJyhhErQpHgDonupBiQTlVzs9bl+hAk
MdpPECQAEZrUMTQi6V5pdzEiXDOKRUOfwVazTNXe1gk/G2Ls/1LTfwY56rEgllys
RvYGxrXykT/kmZ0ItS7rx88Q7gIVhqas+joV7GPpWcYqQN/psOCVUPhGtaSnwoQJ
gDozDdpHAIVBX8rkRn2Pzo5/FR4WyBYgW/JsiHEYsbtX6MtJQudFTRkyLV05smiJ
qE+GqhCcQM4RFwpaWdWF5lduP97xeM3N7FJHjjA36NmMcXYwLWkoA/XUm7Kc0B3Y
YBncrSx/4RLz4ToOmS12bYY5HY6as72WEWMWJtUoa4tRzfzoytbavw+XksXLS9IA
0/9ou9pkJFOAQWJ6vk+qkU2zsSXLgv5zlXSIcX6QkoGdhSBb7u3L7r8tqiEpnKq0
holtURCQdbT42F9lwrkNI0P3lgjU793FuFI2kgrmF8fzfeBYd9gycTtHh1moBwYu
hp7ugl8qhC0YwjTKcxpSK9GkAVyFPgnoxVfsM1l6eppnDjJ6lDvE4BpSNzRXZxQM
YjLGbBE+dWyE7FrvxIx2LuWvBk8NSTBI1Y3SKU0TKYiL6fWPOWv/+vHAP6QslE8r
O35RGHw9pQu47k3mHafRh/WF2L3lA5riV7QGTAh8up9LCqNJSK/1t6USWFzaoonN
ANvdViWrGt0KxX1bPFkO/RYofTHx0p0Qf44E/UAa7KXos3gv4JAUAlosuX3g36N8
2s8J4OgCwoXLV7dhiUvAnQf5l4ezoRZBZWcxK1jPIpCxUJPEPDHsUtn9dEKOShdW
orLVAJQQ/TWHU4+HRWju27r/3YRYUGq/skozYnBd9Y4ImstelztVmy9cR3j8gycM
vDVP3Rtqy+4NitaF1Oyj+rjibjD0CGeG8g9/zpFW851WVbxV83aB52O2oHLMD+ZQ
BjxV6ejolNzLDh/GEpo13zEpeTHVs0sD+IsQfR/PRVRPUskGWQNNg3fmDvgoDI6E
EB/Xl8HumjFfbHnztglMcWn21jvuJDLyeW0hzRhmC4CR81xQvXkCIv8sWHsJETvs
qgHgu5LCfXU1GpSqPHYmmfRIUCzeTNZksPBYk64dED4szhgM69W5bF+LFjp0oo5n
S8+kUEpSmrncNCoKspAYrimLk2wnfdqsGBiW2A4HTp682bBD1ULxZfN7b7pH0oaH
RFwR6FZOJT3c9H5hKyHT9OCrlr5KL3feRbqQZONwx7Q/GMpbPRaxsLCGSY+onC2Z
wM+qXNwmne6b1vuWYFX/RSXt9CZFD41cv/dugJJCSfatTboo4Ek6nwqjuBdpp6xi
pyRNDeTcBnMxJn9/+bzWD96E4FshM5m6NMxLCBKvVdOAoOeLJMOqdsNwqBPUp35Y
+HFBYN3+ReU160GbRKTcAgTVBydfy7Gn+1qgwvMg76DqgrzsBGTQf64AG0LHn3KD
y9qlDh8BoYrQ8WkCCgNnHM4BW/N9tqIAXsX7LE1qpZj7fMIvQiND0SmPe9yry3tD
FC0+raEVIbZZ+shUbVG3Ae/Bq+qH4JCXvOe0XP+UM0RyuOPbFuGNRXUiGvJPl+in
O8r6+l2Dl247vhMjwu38zLQ0KpZ2kTApCQ7B00SFmeE5bm6GPoThVxkYcAlqecRW
y44zDqVa/7yk2ptnVyKhHhKEE21qKRkjY6VuQzgkPAa14QaSozawgnN34oEbgfLO
9re+PqxlldBdvOdOOo01DvEL23jsd9LuBxGalK5jbYEhDapDA7LsiRBjDaRTWAJJ
7j9bbcUqU+B2pIlS+2Hwc6euwJWliIpX7Ncge0fTEH+F76nq2HjMMG9ll6rwB+jb
BltgAhlEW0gXXMy8v7Ls2e7KbyzQhk5+vTdPW4AkijcONcEI79GNuzK87JkJIrfx
kYS1RXSCtsz7O/tYI0y6p8NE8g4Rj3hwJ+yAw8T1gVqRizFyunqQ2zlcVSzW/baW
Xap71lgfhCOOmogz+YcZuA0kL235viZkcXHCjiT51NQ2zsGUZEyhpoc0b5PGCjLw
beC7QBZkuHpwCJkBAYGqMfmJIkzY7qYN2SAt+PPTSU5PG6f+yFaC4+ZmUDXhMvxe
AnL/1Qs4qAJEGxfc3TuivWRhdZ0AtkZcl655Bc6ABj8c/9MKd6UIOazlKW43FqWg
L5/qgEFnJ16BtRJfHsmvqIuOyNQ5clZVlU0FnLRWRDBl/nGZQVTolHb6ftkE7x4j
m7KabgjRqGmbFMPxTLSwumWBR4eXm3/cjU/ZTz5cYK69Z3tMtWa/02hA52UOaKdI
SHStoqONtmTWdRvS/kKnuukLSQkScOO1EzcLFYB/3dyA9Z1G08Vo5RiOPLcRcx59
ou3A6Xh8oujs1K+YY6fXF7PZoQvBY/a9MSuQ7ZE1rzDu1I/PgWOvwRdiqHBTipEP
aVDDP4QzfLCfdWRiOhcaCvl0WzhVtuUAiFP5xngmRzZEir7XCno5m6MHndafGbtH
Mjw43/oz/7l6b3q/dTfjtkzj/xP9YdvCOJND+fPF1VLBfJehSF4pPEFm/0TNnnZC
JWj0dlu94rM+A8p1KAe+Bbufdczp6hmN2c/fetv73krTwe8vb7TDe8gRZbHwMx+p
o9GB28mtvGq46gOBIYfakcF7HRmdMn9YtI45GZpB2OAUzSYcimjOmXdX5CRD/SSO
VtNBWPpmGbTHDWWKslRbR2yIpMexAQG0M1JfqR7oFtHPL5EGlt0v0rlurW06IPkL
vuZrjtsnZ7VeFHBAw8YcMGzmor9NZJp1Io0+1CjwjKn41/8vnbMNCfIM3KjbtvA7
V7pdFmSdrMzJX6st/nGYJFVoG7uU5YNnU9GIMNLdNk4H3WtBN8HdGTrF9FEGNxIq
EeiTybK/CJL5aHKPOLUmFmNQn7ddmbY4Pv/xM3Fzz2uyi2p1+jfpu7NBWFjd3YR0
frowhHujV8BucAufbZaX06yqaarZHCrT12o4LsM3Qhoez3AaxJoxjy/F1eHTGw8k
TZfv8c82xhk/BMA+fogy9WXLRIB0+FdSVlvVQUgKsyXmqomLbvCHeNV18PoKMrFe
JcwqyuqNyY/g714MuYjTGsXvu4Kcs7bYAUnrtGnDlS+qrIak1G0Fsb/Ju2Jc1Y9b
dTm72m2BJNknBYMJ1YJtoBBcS5p0MhDtvdK/ht8D7UeSf2BiLeFwPVttgc25QOLo
SOakNk0nByieWi/i5S7y+PWNOOKH5ShBTeN6typPtBhoFnESK1oGLYoiRVnwNu76
HRuaGbzRguGT7FlczkAwXd9xnbqzWpq6U8nHoBAekdlT2j5+/e8w3NtU19yxRtgc
koWbcdhTGRgpiixRgUXguRMhusBkfOK4rKC33L+cOz9IpdwaQTGisSylMyfxwCcC
U9xO64XzDO7UUChluK4/p+QoG4Ilr8T1IrQSu4FpUR7dxKVYgQHdVKUaJb1PLI27
wgiLbz/WcHFWVEgIcxDP0kVisJlow+rTtDhrnZU9oT1mCvYl9w3ZLT+KIU2+K73g
0zzFXXiqNbqaEwkE4LfxeypLs03RoZc41V5b+INVwqgsAt458jH5VsZ1qhQukERA
A48jwfqtuitMJIbr4QnnCmYiliTH9hG3rsUIbX1hLb8QX9fWrCwBF4p/Nhj4HrrO
PdPDWp41zYADw9afWtdyRIuIF+kb7YGZ9MKNxkpWwxfZi8ttzvSmlntDdSjeqP6k
rMNrSxEFqT/Z3IZHX447/T+HnPsGTrJmkvH2dicHo2fPh6Q3CuFx32cua2dWzgQU
lcH8h44ZdeOHJkdjImEYMSynY1zg3NPex+fXMg+1WrS9gvcC07ifjjtDdS07uLyK
drwynJ3Ths8iatHDJzoqeZEvNXR2eJrUANUtGycwbXBFdQcAb0Wg2JiqRvefIzSo
sNTvrovoH7Dx7+TRVuMiSeIz6RSau1jDSdqMH3qjycSwaEsHcY1GJdEza5phE1CQ
rUdMQtO87SpWEUljWPmlLlydYxhq7C2Mye0WReEXLeTUs+Ld78YOUVcFs3NzNM/a
iS5iF/VyaaL94IAVXkGAyovzJP7MQOHSiIKhST2l4ekb1yeAVSHA9npiM+iffR0L
uUdeRGEeNQAdz5UzWl6vDoFHWd2FQ3fe2BSa++vMuVl3IDiqObQZhr1k3+LXEcOs
C8f2TsVtICCcsTuWqd3rd/irclGh3zyD2hN008UAFuuFgo9l3T0/j2a8+xk2FO9e
qeOQZ4V/lTLNg9deEoQGCCaECc1k06nHMENET33X90iiz7zG1Kae8UPoKfArb1Re
Cm6FJvinwZ4q4ezDPTsO8UDWsJj92c+ktNle93+0ZChbUXSSqNaKptzs3Du/wEIJ
QedskrkfhpXK85Wf3ZA+s1WcL1hq1VHsK9YpNB6kWICvvSa0rhcGBemCG0LRoCpU
GwBny1OeXnQMMjTlrkzoaTo0J0lLBc+aiDXraWGxqWAbApsIUmFrX3g3Wqek1EjF
GQyixGr8De3T/0oR8DD6p33L059A40Hw8FK23aEP3Fsx6GNLn1wgkjR1fMV6Q3KU
URqqW760g0pqcinuTcM1+CbASRW7scPmZO37cdYRaGe+qo3JXMxfNNOsHUE6QZwz
xgrTO7JO3xUvzA48gmlW/tsBBtcMEy8fg6SAVMwCSTNTPFJ+OVDWDp44TGyh3VZH
MP75tN+jguPhGNsclPJ9zv9otKwUhUa3de5u80+dF6VkRJ0YqqEzIv9ZoSlQQn22
WEYlQ2pRfHL8jNYzMbjP4paVtPrPXfTB4SjP1tMfhWo2eBtiOq7uvqVxWGXFOozo
yESXCbymaIX0UotU2lQFmGp0wkbiiDPxGTyxMQs9KCQgaose48LVs+bJ2tj3M6Ux
0bULsQD4BplVTzruZIBp9wdQUpLXU5u62bLP0sNIpv22fL4CZAh4P5D0Se2dFf4u
U2muPQGgyGjZRevRZZZJta1+AAADxwa37HKKCzFKkaIdPqMPrdOaCc8COiYIXm3N
09ipoZGZC9rv6l37buzVgXJYkCcaMbNMz4nFmG1GloDnpuTH6pzTtw09wF7ubSEX
XRyoxS/4zRTPHLy4OrXoSpVKUePXP+XrDGpDD2DdYALplmhn/+4km+XbPAGTbdW6
AlMtVMPi+trGv/bCSCaPFTdX2hBlc7AheE0jHueioMtnytTss6OfVwPv3Zrh/Hbu
r09gKTgP3y0Buf7WL0TIdPVZko2NmknKBHUglmVQ8hW7C56u3umtflEqrzF8mLRw
OBBVbuL+l/cRmwAG8gAGQslL/2kck3rwFAyWUnKosrK0Kk9CWOPCzFjt/6YQ5vxj
nwjouWmOCalgGIxV4w4OhYgrtmNPglEgSExL+vVlB2lIUVA7m2Mo14O9OL4nO0i4
JYoxLo9lTe3Gh3p7MdDOyWTE1IsJORYxSkc0IHYRM1cYypRx0HxVZe8Z/esC0buR
IIF+/p1D4wsmRWlEvPJPTKv0RORjuAjwCtmdBLOdBpxfO3IdFmC5zocaU4LZOp15
bFuX3z/aDwiv29HoYsxN61DoQd2JIBitUu/CSlVrL49ZAG+NMv6+6PD7s3KQz72F
pgY29AKNgISQRoe2x8b+UpkVr0fJp9SLMY+KnufJjrKiVhZkD0/t8umKPdw9BNwO
NkObEfRDkTlbmdcjGyzrYIVlJzTBWNqyCDQ2p9LBlJHdd22Utag6b/FAun5YAS6n
CSZLPEOcv/cIkUIWZkliWuQlOgnYU1YkvhS4HT6HdGaEw0Y9f3eYnH9Jt+GBkNA/
HFg4ocLYRwtJVwHqt+J/+OdS0G2aPnuJsqNXmgJKHzE+sAva4Gomqr2flV5eZUh5
7ydRCvhTkwcGsfCVgvhZ85Rg8IJwRieZ1Yh2jxb6dChY9WKI813wjVvgmHakM07o
eiyKSrQbcQkShft38jzl/lvzoQRcs3AQfFPNfd4zfvL5YYDAi0S1T3xTyLR9a+mj
YYbXw2j7jD15627ENFM8oPGGUxcwph+XCnWJYpYE/Q19nDSyDEOiBS682b35K2Cw
Ewqo/tBPrcEYIF7nvQIg9kPRSLaYcwDwToMZaNswvpsl7/mHJQkEYMK2MVUVGvLj
qdGjXr2w7RSrFiUjD7+ROm6+kdqltPQzWGRsU1PlyL0UMym8Isg1hDbwsPWu4iHY
gtwf0LSt7b3314ol8+RsmSMI9lr9Y9GiPnMU+i9YuGhhZp2kiyivsmqeUb754s5O
a5bkK2uEMPOsY+ByI/e313EVGZkoBn8M7WGeIxljX+B1w1ekss7CQhiGQzW1yThS
zOAD5gH7xzRC7jIDvbsAPnBskB0Kye0uvcemdxQaztHGHQ6X9S/WUBFYMM8RvlLT
Py+bnWRIAcxYXUUDI56UMzS19UrRuQfSXWN2DtWL5j16Zdi0PKhuP9oEX/qucf+7
UoqvtD8T6pYORzuMPGYPeJjRkf4/gchMFI4SdguXSY3kFyLqD+p4ty7CTQa/WVbj
XtysjAYFxBpMgQFKo4jV2+Sp1gT6h8FwzW4e/YzMMeYKDN9ULO5COuozk2ABJmba
TASyla77YtE94spEiizF5qVBwDsSsQ0YVnaDeoQVCikYmuMjSkF1ujYHAh8zMOWZ
Y0BT5usQfvkwNxKtBUL+bYXj08tVjuAGV0MhYo3l4/2lH4Y3N/Y+DUf5ZfG4FCuF
/LjqvSOiO3OcwPNbJ6aa6QOBCn4rVqJlbGFUwxGQN/Hf9IunnmqYYaKP0a8iKDDx
4Y/cD3JMIy+Cv6rS2//4Vzf3EbaQfFb0pKnXc66gMeeoiRibjQX+Z/kyXagd3rO4
2Hti8bMa4AGIMZpaHI3VQ/YLdoo96uoHjccJJpUDA9FoC0mjyVswqPU0mf+me8G+
ZtGsFcz0n1I6i/kBPS23R/VRPjWD4LeZTIa4sj5AkXiqmaXLbPkPA1TdjobbNGFb
SIDidpkap7kwcxOlkYG+hLxhggZ/97hiP56CK7a9eKSNQicoT7+MdJK9b1586JCT
5SOkLsu7v7pyCpAXSwELREmMdgrmDdfaI/sLf+OKNAG8cmg7MM9tmGdsYHpbTh43
vr8p2DkIhzbZXddDzaE27+cTAFgup3i/HOni2bCXR/SvsWxLuBqAglyA7ZYx/V2S
Xw7lNlYm5ndx+9Xdt9dXKYNLNhQsDB45NMDJz8mj2drshgWMlUORlge046BL2XCB
dR9o/jk4SuyvaVjqd0ITovNCDbnKG6ndJL1P+91aOtAe7dyT+jfu8SpfRdf0LRic
/Xa3jv+ROU+acGsHDieBL/7y/eD1dyPjYoV7imyS8U4UHsZOG5MVgcN1U5Ry7J48
MZ8hWvhu0tzGZYHvGsVsbNKOnMR0yLDHVFz7Ux8Q7jBef/7+oDA2jM/h4D0Amnbm
SY6bsSS3jKkqBC6GDuUz4FS159YBYgBVNzQiBR3BgHnJ/+42+KTiOdIZm4tr6t+F
bKmKQNbDIHGCPqzIi1mqki/E5rB1RWV+veowFvZRoDwefxeEVHnJfVSNii8rFKkM
IpulMe9ObDgrUpIGAV4KKBGZo0TzVpaMCR5pwiT8aAGMBXF78RktCjEL246n9uhb
S62qyB/hilgSiOJM1ahy7b89r4nADZ8Iy2QMQuzV5tXotk0H/R8ENLzt/jIwPG4h
h8Xd+aZmM9dris90Lw+Ymvdk64YX/R/qGcQ+EAhsj4ealvDOCVNGjGMdkuhU9Gc4
0Jry6iyX16isKWWGcq/ieScNnYcX29DZXxY7z2K+jmM3owIGeRtR2QVaUiZS3iue
IFfCa+uJFwADQtHKOyGZvhRWRBWqddtXYsThBCZFqcFv5THiETXnlfAuR0UeeYGx
ABwnf6HgXdYBFFOC7cmxgP/pRM3yEcOG9zmuwtPCFeQ1pJqZUBuAAf4L4mrZQIQy
LDTNEyqdiXnY2aWhXw6BJLIhBo4jnVccpZCX62suade7Ds43o2XTcCv2wsClePQo
PL4XF2yrOltZGcoo97ZuvcATj6moPyYAHR1BNM4bJ+sfEiX7/4jDCxOHZT8r+wrw
bDjQ25mIB8i/l6FcR4k9fG2uwsE3jTOq970EOR2ZCl3BySd3YjaBrhUzWvxgAdo6
iif67Uh8WHu8kI69T3OlyIWlrerwEM3I6B4TawRqeZwgE1hROVvnE8QrtovFH4HQ
SuyKiwD8c31q5Wy8tmmHJnQVo4nyyV9v2WplBkvwpxwmEBMYLgZTDmT0G/oiDTMP
5WyHnWJKIhUdIFlDurYpUc1p7FudZK7pRoNaRxs6XdTOdeH6sy7+LsSOmGXz+LKF
0IFQuX15ZMROfn7CuQNYv3CEYhESJ4U0mewrLN4fKnL5yOCoooaRbIYZEEscyLN1
pP46+nHFECBGWeAoZ82Rynhddfc9iZj6mv+eb7SMqQaAnpGY+DQH7tvy4q0Wud/q
K3Vs1YojPMk3GEcfZp8/tZCijO8XQdBcmDVUuiGM2zPqm1lqnbm1bbP6PSfAm+ZE
Mo1j3Pkx7B1VZvmeVXJcyLe+tlpqTKJGtBXDHFIRIuSDRtFlPNMW7C12QsQTB9gn
y595+nXtTzYS/qsJzT7lHP3BS3dx5dZ2W3dCBsRWFlqR56pCiJBVm0NtSaf8AfiJ
gYIHmFtuAGRimA7Pqw1E0/jdHP/3s1GSRWtqOJx+EHexqy6Jnoq8/psNOIvM9Isa
6jIc2Z/HxRcjAN8hfIqCQZpkhzoPEXVGTrPp3+qyBxdwenHzt7hdwt0Zu4HFYQDo
3853ua2Gar+6m5Gr7MC91VJaBqktjlp5v32hGDIsk83c638swBu+bY3cmX2y0mO2
Z727HlEGggwRybfUggZSwyQNMvC9KCSiPqHrJ19bRYXSFctMPHcB+5pvwBj/lGhB
BO4Wt6L1ZfXjhG7cfdpAMF4NXNQL6LdNXFUFBEFwqMtN+iBhzbAct0MScVDPHALI
GZy0ZYsQ16bdrq6BXJscFlE0WHaKTZ87fBm7V28FjbCd9iGWxV/mAaUcK/J8zN53
hFLoemX7OWhNDbU5/e2a3w==
`pragma protect end_protected
