// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:25 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Yooia6ED/bTasIn79Eab716y/nQ8oMYlTuG4BK36H6fcHoy/V++uprSuOraCLUAx
t1GZ7OZHT3S3B2ixvFlDgMeHrfP/pUr7gzQKmZwGOc6kMtYmrGWsBuXUZ/j+6+OJ
9V4PY+b6or2Jqfjy4lBAAP83EOq++hzGyz0C856J8uk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8864)
LcFyoaQrpmEoMz3/FZzbgAjOISO4PoVIjjsvo8d469OTRTyO/NNXEwH0f6qawYKb
puigK1JORPbxF4kmJsRpYeYUUYxtsuZP5vLIFl/S6wHW1atceTSDueLF7Jnm5yCZ
LJYf3Eyo/5Xpmag5HZ/85TythKmY+omGy/rfw8lysLXW3RRNV2l6CaFAk4+GMJXP
wml9WLcXQ0SlR/sO1cV2annUiEJ0LO7SWdjPvpXVNcico7GlAUrMAkm4gyk2XPSH
rX//XYgfOrD9G9qOOzQ3J7SWbLD4JLQllbHZNZic05IWo+w98sBFtCdM10AY52t8
uXjhYrFV+2CBZNCcgGEOTqf2M5ic/8wA/14V7wqnHGJLrcfNrcGoLLM0cpKdKlBj
xdSxsNzqmMDyltO5jChtzcAyXb49EwD9uVPom0Y6Kaxq9SNoCMgzw8eZVt4uu13G
yj+SiCztVcEJV3O4KjIj0cjiaErmy1k61PrVrF8Ps/fyPhMnFfavWTw+VK73fkWL
pnCxc3IEoVRlJs8Ml0VytrdlhK+9jYVI9F0nQ0pcpxxeyZJLvJBUqMz4ErjHQF8+
szCtJNv8wz+jBnwuNbOaSg7aIgxePbX9mWCk+UiZg4aROsd6B8milfaiRuesRBrL
Q8zBvAG5fkE4gAYXLUcFghFWJhPW0EEhZig52lWqYd0WF20jBgovnoKFIBXWpgSX
KD+fBDs/plDo6MmndGBQZDxzYYWJxNnyHR1DVl54wA2U1WbDjlGWb/YkLGkCIQzU
hCSnoqOfJ7SeWtlX+eRSddcZ+GGzCEZTbWS59jQ1IItKhIs1XCG3NXLjQp/F8p5X
2wmPH6NVAtMZqqYKD0Ez0Xg/eAG8/u5dGQkPg3WGq3VFmbbxRrx5Sk9CoBwJsAx1
OGXuNo+5AE1Z2ogF+ET6Jmb/dZN4NbeGpkugsyYw1UYiHtW6qKR81fGB5DzR5h9N
BeCPwEEsUZiqzPNVdlFSvPe2xeYGJi3P5sS28SCThX8A8SBgtGQrR8hjAjcbkYlu
frjAdsli+AxvJuK3+3smNrVIQzSDe5TJst/mbrQpAdS7zcj4J6wkPYGQrQNctkSo
ZE6EwX8+kc0v7Kz7hwWu3jPWwkLa54nktt5Ehq0szDws/Ia0RR2WJRSDEstvj6QH
w+RtURQdjWbXmmHc9dXzI7Ijjwb9xXTazFgpL//Z//lcoE0BZ/uhfH/wuWAwdRrX
EwrUl8tzuWUPMd7to5avny3yRTdNBb8DdbBc9JPyl1IJSKIV9qa+WZVXjZheni1v
ESfVaO2iMuGpkyRPG4QMbECFrLH9dvKg/I0QEINODeRgq72OE3UFeCsBKIgEgn2W
CGeyes7i6aIRkuCZdchpyoS5QjXxfiJEBcuVmydLQt2iQcgHEidpO1PM8U3gQ6gz
WjZhWLBjlnkII0fCy2upUBF7Aw3dsXCPN6FVXqwnN9TiJB+6I+z0ah/XvQmjA98B
S4eh4ASE1ckzMA1ep6J+Wrt2oB+bvSdfpGFHnIheyJkaGBvIME9rtUJ9TJ8+bCMd
DNNCDyTUkohwTGQT4U5qkvk0sk33xU7cQlhQfZL3D+y3Ad36VaitbRHBaUOEGJMj
PPKnoahP2QpVJHS+pHEhxCeFqPV3n/czv2jAq9Rj20DRB+C4u2hlFL0a5RJhzyDp
+dYh1ou724KVbBVZrW7JcB7puYjp0SE4Vnro1qoJPDRUa5Dm+fAnY8DEPQBWL8vf
OR1qcK6DB1yBFBf48sBq5OHASwop20hcWA0PLDCTB38F9ECCIJh1NnalQlolH3li
jspP9J3S8pGoO6WdxDN0fzm3X+OIYCnV9Hi8TvZHse/PclHJLarDG9vrlRLGJSw4
3u3ZR+lThOWI0qc8GiUVWhwhqyuQglCqnGfasVf3w5XieN2LSu+cs3YHQN4rCgS9
Q4aO+MX1RHXpcynb9j6HIJUBB6htd2ZoYMd9CNS30o01owtXzw7TDAsFIcoMxGYY
duZn468HfD5vnOjTzJKklu7U5Rxa8WwberaW9uNl2jDcri+1QCyKv9VB+PO27eAb
/NDZB1cL4VdTWooCIPzaoXiEiP/54W6W4vAjKFull+brv8E4HF7lfwmNidmEiinF
ZOECBEcLIUHPGfMeanbDPtcja6TDtE3nyQLCHgipKpCclGaKem08zGzfRMH75qQv
LWKWM16vK699if7h5+GaSYGU9VVdx0rGNiqrE3nWKCDVb7mtTSioekgbCsZjgXBA
jqtJZFvRk0kApTd2rvHG4fNUUM6vNgGOLTyQEKlZI2dhKoOyiWHHtmXMg/45iMVB
vasi5kAzKtoKPn44irEJc7PlBr/bb4knoUcY1Vk+MYC7KiarTRST+s1D62+ZLvvZ
VmxCqdW58KjpugeaEVLxNETus/sTUGiEjeH8IdUIbQe1nCDhOn7PHreK/H7eSCIl
Mk19ol4dyAJ/FloE9UpnEFq3alFFjPGADHmMquxsxqZGbeXONZ/RWTa6+rtQHGhv
Ub/Do/FWI9R9ecdG4uEnO0CbMdIroaIZgtzzdcrHiErombeifw7nRNazWPgKalMv
aykS0P86HiGM2bPnrW0lBHUIejUNVNsgsfkKqaeZ/+PsjkytB10v2VI2lg/wdtq7
7LmhMnu46L+hVPb5eh0Y46pkHxnkjY/8K+bwu3vAoVbKJ4xmdDaQvlUEjXY/1SJo
4vDgv7vMIdSnky5tmK+6heYJ1a8W6V2xX9/duJmz+pMgu6JaUAw10wYhANhcVkJe
NXH8b1nbE0VC/qVyCjm0DxewAhEkFpT3jkl6r5wtI5sRU+fi6k0VdMMn2sIBFHE4
CEkcDBoN1JBFHpgN097o0pvLO4AO4wYLyt0sYXgPCapN+fUm7svgGalfoepIpaK1
BXJUm+rIXt7fr9zzOX2ZY+nO6uNgiRfwW6vleKLTziLw/6NqskORFT2g/rFmcTzu
022Eq097Sj8qx/XUIvvVqPxxIK+9v48wJBG17Nti0vmc20T3LUMJ5HecB0sLJaxN
mgsU4Np8ogPqGulwmFuKTXTkgzT3URwjSVBRdkt/YvHuscc64xr2VKZE0x02rgN4
PRxxHFccZfe/UcWrgHEFLS0H7kcaYJyGOYDT2rFxveat3vxVBo0oBh2VIW8GgQ93
dzRSBmUHE2l89r2HGF3zJr3Fes7f99wr5nC6DMG38yHaxP4Jm7bmtmYx8E1TKr4p
YDtply3U2elpBjqVAUlnR38gVk8SNR7Vj+RGpMDm3EeTNk3C20Sdxz+cAlsbxs8C
8VC0CYBROMmwBcAV9bmAet8wvoltxvaDgu3Cnvhxw38iL8aj/Fyd2aVLQRUjDsYj
jkLi/r3HSeilcYoLaEu3Si51WVDLyDw8PHrGdIn0EtVOQs1F7imMarJ/bmDbbF6d
SHEZ+ibhsKsiu53fU3C4ymycQegvgRECfTpPYX65F1FR+ZPzGghNB1eD3OvUFqXz
+WNU65tPKGhlgWArR6yfA728Wvzj96+qoJYavceOButd0LarUDfNZGIr6G7pMAFV
wGDD2KeD2/eakS7u0EKaF9Clx/WY8a25LFR/ewn7YWc3FJJ9l4K6Mv+Q7zxQDF1K
YIf4Sfs1DBYidZcTjpJTLhJ7HRB0QcvW60HKazr+rkijfCSAdVcGWTSRJRPtgVny
tQ36+BSuDhmXxMAN2qVmfdDTSQEH9XEZsGLEJW0qjY6DIAQScSpGKKmHSQcu9F7I
3uHSN0MiZaeQ+FKKItmtFVuNrkb7DCIX0D5b75d+ZyxiWu/P1HLFbZWaSI4LVp1U
CxePXAf0t6zHK49+PJKdSd5GvHBBbV27WFzQyjzGuf9BewVvGlfq+OrSHce575ev
4IRxUkWdOQeHlfc4jW8uPPDGBeP90JK8ebtdakTaUZ6O0TDauHYa+JigdMKnLXQp
3//EURHm4+GqomD1qEKgJMyWKb0vQQ/qK3GKU317Fj8MnlpmI9SUUlsv6JteikDq
UYIUUZ3EsBi+gOSmTAN3LDW/6pKvPks8IY6qMMaWIAeWAFDB09//l34caHuf7Dyx
HwgnsVRIdpr1Xq7CmilQKdnFt3nLLPW6P1AETMRbR7m6rpI83qn/KdGkBjpflx4k
depdMbNYH7CewvGQl76MWuQIEJo93bzPqW8XEVfHd1Bpgg8Tg+UxCpvKdblltBLA
CFwtIxv5N0eYKjjzxPHDvwvIDeNtytBdva7A5zoFrQHSWLWdoSFoNQvaw701b21s
g+1MSuAeFYSEdk9s/kIet2g2JAtuwwURb4PV5G6wST3HXxMos9tlnCTGxE1AdiaI
DWfWyuLEM2djCqJIH3cAp/jDTLJbcvaetgynDM8YesP4I8m9l2YNM1fl6nP0XqmW
H93h8iSB7xQpY8SuCCaKvAWznrrhjigYwomP1R800A26kmr/8CwHnEX7I4tUp3nq
vG+Vz6TcQvCSLDdC49Mp13C0ftsFQxeHXZbkO/0bddyvZaESqFNt6C61BS+eJ27T
tH6mXsUL5k3F8jUqn2s5NbjzI9dlBhpGfXJSUj7E4PraYhWXY8Z2uIsuV44MdT6k
/u9gonmUNg9+IEk0+9edszdb1ZFKgus6XjScSXVe83TdQ8Yd7uU49P4PO3dzO2E5
Nbjt+sKaoTWK5z2cT0kNnp6TKjDFx246Qkmx3Q+HNOngxfr9gbDJsvuMGaKMfMCW
otJ1TRV7+GknHgR1QUrGmuUYzHgRZ7C1qyuMqpKT5/qv/gbI86UT85x95ATerNNg
KarFV27Ajj0EkeRYQ16BeaTXx3/a+vlgtb3eX5XmkPiK72eCzHsD/xji/vQNl7zj
iGKBLNNHy3HbvnUNCyvGb4YnIwzMRbZSosve8uh5/iByJ923eKB6J2PaeTwuZx0V
djENXTM4BrKCMwzWe7XoLoQqPW5IykKx9kNnT8URAGPFYBwsG379cMjryLRUHwmi
woh0ZE18EVVzFW0qFPE/eBGISxJNxJuhvt2xxf3/mPEZWpGLzIjVEX8eG0Nq4UeO
FwMXBy+7bx0Zfjky5jbR/XrHumTwHML4Ebb5AzUIauYPeHZFEQRFXbA/hzGAx+fy
iAMnouRMwhE7N36vzlJsumZLUOP7lcJcuFKqjSFZg6QN7NctWaqSK6ywnvtirm3s
b52wZl3mVJqJGKirAQmKxkYQHdGZ04aRwlDsHGFbhF1TQvXKOhTKFkBNtcY6uSuJ
3Pp7ibrxg4/0P47c8QM/AtrM9XW09t2pfg2OgriMoCGLblwlEDe9+izFXd9x8mDn
9GJQRCMaxNA4Zbn5i5XdhNaiA8a4nppKA4y0v97tAT15wRqpVx3obuEwSoiHQlqi
gOPMUiJ4jQ4NB/eLuYb5oP/A2nwdIC+jfHFFMz9JOWMj9/19fmy3E/KGJtOvP3gw
bAgP/2pra2+1CIpnrL+QNTyDgJPB6o2xhOagXP4BLTJQx5Kdmgsh4x/HPIXwIBcH
TaPbWWoJP6rHBw8CkrYW4RBYEqAt9XbQ2hwUGV7LQq6BqceLJFjWLzrWHX2ZLFQd
DnymtL3eFo2VGUHj/ktc0Q6+zLqwl7mUu03zm+m2yW7f4E29bm2Wrm3+QTndSX9r
ORZHy/ULKAL07b6HuJ6TgEVIi4s7DrgxkmRS5EoLps3dL+0h5bbJsvTVNk7u5Gvi
CJpc1p2UjCFu3rxxj2n85/3jrahS5TpaiRSKc05iKxyF4cPILqJxldlYJigSoTXY
cQHjpC6dMx+/5xWQ3N66iSyTsTUHGHuXErb1JsXtstzSUH6ySsFMFj+DacZczk+a
kKT9LF7RJVQtc+5L0vHtNyIncPfkcMNlzMvL1j82GBgNo3YZTA19uM3Ho3QgJiOT
jaSYzJM5T4BztSyHKexsmfqTcUHEI8P5e3CA6Z0Tm2e/yNrcpqwx5DEyDJAW7rI+
46eg7LlIH1peJHU/GQ1gPkqTvBVaYkYAv+/zXqsqfQOWSijAKKS9GQ1i0wCX7h1H
pWZaSTdLZcxPXMajPf5SyTJ0fjnVfBJrDJaZM4AJgoZDaLbim7mEB5Z/J+dzGZgj
IEjg2xexIQ9xPs+f5YlGxxeBmivZySoGdEj8Wp2YBPx5GnZh3IHynGgbBzwJnwrF
1SooHWF2h6pofZCMPLr7b2bvfT7dypHdu/GaLcd51zAddhquwFjtYUYMIGtG/cCh
62RU11QA9LKAxRt4O0jOrBFUHhcBg0z7Ds+TUJ38pnYxzBRPu/QEFUpccs475jJp
VjasTZZJI0dtcffTge7ef/uX9dNAOWcM92EPoy6Y9mlr1Q1kNsz/tW2pFtHv99Fd
uBBNCrF3i6qwj3Q3c3nmNwpDkTqXAqaQ19ivwnuyMF/qytzG7Evd1ivkmoi3I/wh
+FosqbPyGnxILfVUCUtOfyp2rKFr9icPKAu4hTdni0o8dGDbs6z1eToaJYhwj115
3sBZksIW56a+AloFLM9LFQVoQ6EUREY/EVg/7iVi5S3OUImDTcaGvCWdShnb7Cij
I1FEQDrx6pXoCC0du8wHLzOLkiV/XSeCLUgECOpr1vSNaUvdTIPzcPoPgsKZXzZ+
QtrQW7bh+Ita9PhfCoSgX+LbjPKEaXPd2366XMPCj3JZODIeDMV2FPrXofVanSgA
t/Eat4i36VNqWb0cf/avru8JnHcu0Cw5CjA34DK8K/La0I8uchdHhsmYQAhrET6R
QAS4jJ1Fc7wvkxdUQ1ZQsPsoisotPIobd7h3ws5pyWbi2fRRGS2aGMV5bL1mNZXj
puA/wlf4326ebjw6FqzRNk5x6fun+e+frG56adxXd6B3W2xrk6m5BY459M1Owmik
PDEqS+Jh2wAzQDENnxu4ePaLLw4WobVl7ZzFGXii0QaV5cxWyR5DFogSBzdKGoTZ
dLALMM1v5AtT0G9L4k+DpZFpuKoV/bUh0BFV/N+2yTdi+/ar9T5ZAJxOuNehWaSc
Y8dhCKKrz+pH/n0oqS7gkJ1xkT4dqH1g133Am6xsprfVh82NPcyeJFNT82gO+7KC
Uqlt84CMD4Hg4ISGW+6Ne23EFHLfyACeSaIjuk8lvjqTS7n72uklmMhyFi+AFBA8
Nuq1/rAOb3kCkev2BtHxqZr8MtIckKGUIaC47txcQTXjhk7Dfx37p7cIsICHCAu3
PE4E/h5Aj5hNpGxlcrGfcIQMchpVng33Mr/ydTcaTQMgNU5xYwga8hiSQT/5/fq7
wHLUXHeFw2KzPckj5GbFz33G3lZcOARs7JYYPCPApP4F8a7OwlGF3yfzjgc8sBwq
HElusVVweG/TC+4SViKUfloJ6/5DqQhFNClFmBHfOg8Tmsuc+tFQ8+/rvG82rNgX
WFnxHspaINZ1UlBFQfabVqtJENO7jw1cj2DcPobDY+UzaDoIpnugZbw0eq1+p2jg
zmL0Wq8TD4Do8at/5TZb9wkQc9QqwY3ljK6ReHJMZbD65yjFQ/i//ncULSuFE7jW
4e7fBCoTBrMxVkJW/RAvE1EnSJ4z4IMEC9Ks8IV7IBfMzPV+OS0s697VmyYh3880
QF+UMwn/UOi0saXb0foI5H1ukVj+WWiF+qGXzCwfqHZ0INOBRUofMbwWQ8PuTKaS
POJWjylwf0M1sYrSmsB+HXBujxubXt12v2E1YNbd4H9PIpVQJDzbJBb1XJ/zimQ4
0KrS949SIk5RuXcP/jhJbNcUQSsrGdrFE4ZFQhE5hdCsS26jXAH64ZfoxDqCBA9b
8W/C3kW7sRJcpfMxi6S0Wdc0GimwP1+ndRsD0SZcoKPNCnmhqfuJiqsAdSIMPQdA
6/iHmkHU0QmJf2FEuXoSfLNHwMgvldYkcx18lR82VbfWzpdFjvVt7oWSYe2d0mF2
PvUq+4/aYaULiJLIniy6PPPzq+Ro90nVIAEjSk5zBLAaahsI3u1n9p2cUyrZx0Bn
AarwdpJegKzYlbjF/0eCuQU3P9xR2a/aHfgYlukaJJRuiVvtQiseaFAxHwHJ/l+2
v/uHNZ6crGQ3JxjryVuJNZAvc+1cyxABuDmvcbhWbfpgLR+prIv69HI2MYM1TVjA
NUeSoFOMeuPL5xSLBwjXKXgOzURu5JKeuv6lMuGjXPoM/cM3cgqnBiT8KwYYQupf
mk90ywroaw6TPCPBSfPDdtp21VkJ2k6BU6fjZjzlc0VqIK/FCn+MTEN/vecHf/mk
zjVlC17c6xH/4oB1YqrAlZuA+iODRqHojDSxrv7XxDJ9hOpDDvkDhhIjVxgEHKsm
D+haymZuMPnjOhR1Id2y+ZzfTITj1tOqnWzHeykjIdVLbYl7i5WboQ45Xk6mgQ7x
KPbpNvsKxkBMVvms2rXESZPFLsRdacwfg8EMG4m1HrFi8zS9R6z4Vg59yl5WjFqZ
cGimBIFJo1OFsH52fCJHFSrYhIgL/T0OY3Upm1t1Ayuzuq4bxQXhJt9uLMkfmftC
ChdzKuPovkXw8AMube/mdakv/HhpZlqgNaMAIH7oSPKCoF5QIY6+qnr3Ja3SgZIg
RwJ0a/D9mCM93PH+V8h/hg2iE/XU/3TSeKMPfFeBMXqg+oKeEcZYX4rkERd4kEZH
0f+4emsIEzZRDAHowqDrOLrSlfKd/Ex27nJmwV50Qe+Uda741wrW5yvPQm1Gyje/
IdU8pjprmbSqwYuzd0fazFWVLg0BxNEblpi24oVuzydsVjTA+JV8GLja2M+nwMyq
7af5BmdxdptMCT7wr4bftVYMNRym/5JG368K39waLj5FgDpS7qFd+BezsWoY3jrh
pUd06fLTI11RVT2xB+psogx7Kvw+o4riK/LLiUWp7wZ2WgXV0PEV+RouizVORLZ4
P1JvnidmEg4c3o2cRhu6qMI+E0BryMYAOLOgBhpSsHorFbT1IcZ0bV/cdbqQXPRW
cxaod5OmUCZvDR7WKVbqMp7g1XbUGqesw+b16LmrHkq+gTSiw+gTN7W5Ff4lpLfB
uSQj/3w+CGFsetSn1xgOdpJxk4lp2qpsKOfem7CpApwXFAQ8SDVyQZEoEOOdiDj3
gsw6B4T9uDcKqDXrX+9YJ/y0sRamBxzbPRF0PFwjYTOZrDIKBOZA7anqWuR5flUl
jLooSokoUiGYKTOj1MNfj3ZZnMFUk51B3EkAO8m9XQM63G/9BgsZ8op1etiEfpx8
KUKkmxzHcyM8+yUVbpPoVPIxrtWpY4rduhQFf4ZhO1PKR7peHga+rIq3/a7SLJrr
x7H9svyKbVsTZaqxq2IBhUFIHRicV2JbWQX9lsBO0qvsDQFp8KxH844ozfZ42V1E
D18bjznv+q3YGIALCtkxken1FYUTXRquEbrxihij7ergCVFvCa7A9iEYWXiNdw57
HY/D7TX3AFawLDLifsvdhSoEA4p8CjaS0Etr3Oow9aml2wvGye28KltKcfz7Or4n
WlvGpeRpa1XXX7pjZQorc7flDxJKO4qNVYT9NlJp8rif1m0CzTUX4hLaosaK3ket
eyfNssrd1PtYY4Oj6eQ8rzepWuf9hNLB//e+02aclGaHnFBNjxuunj6ThJvy61ka
ZEaF1uCifp/rHTz7Sawpk/gxf7MyVMZVeAWCEJUwYYP+3DI1iWhBBEb39ZDOuvGY
HafRLBB2Hc57ASEP9JskwvkddL1evHD6nIAuvU4CGg54s7PcmXjrmX7K5j+1jbc6
aTM054D9+r8cC3Thr8jCTXa1/xSqshmV6LTSXA6qUf+8UG7gwLAPy2K/BVyU668R
KjhIQWZO/SuWfqYlUOXDITiz89FyvjFxb5H0CNyJubmBXti0kkHezggHbScdYBEy
yC/IytYTs/9vj7eQ926l7ByFUT/Qs20pEzw6vw1gxTo2K02m6Ev3+SJ8+KczpI5W
E7+APjxAP6ConJaCdP7MNyQs7/AgdwHso/n9HV7Nl5QGr1bcMLgF38a/GI9hqJRg
Lo9zp9O4RzBmV1B3s/wwTImpYwfLPVzxmxpYYMt13qY7VlP7VufqIYh/UY/zcRmZ
LYDeTeELIBC+cvGN7x/N8DngTDqV0rOIBQBXk17vPDyC8/GY+fWEGbymKeQEGdlU
nqgzWpag8s0ItLs1VK8InLXG9AccKVDHgxVUkqZeqZxgR4dCWWXbAn4ZWL/Pyw6l
wjnnuT5vW9u8Ne2dFxI4Z84q/kt1CVU8AXAE59fb1KtgzWDsY+QFdV8Lbdr4BICt
GfaTAKeeKXlX87qWuZvkg8Cf2xgbloCaKEL2SGiL480586lXEmiFXIWsKS0l6uaS
St3GtlgPd2r+QS3krnnMgzDudRh3u+c/+F25x2atgvLEGcCfKYsDU65EzZLieO1U
HanZk0JNH6S9XEqdOx4eWtxInHGjjJ3XtEim2dGXLz18BAVAy553HUPf2j4g2z7m
0vCN0gzZjLEeMg8erjsQ7GqQApeFfBNNpJMWNJEKyaCKIdzUDzf7n33Sv/gif8XU
U5oRKnnJ10mRJ49yPQJbzkqZOgDd07m5OnRiCC+RrGzHLQgbfIU9vJb7qeJG+JDM
wG+nApGKkSLuvy9O6qHy8l4uTSD1tea+w2/clF5A8C81TUBxpbIvMQ9vDe2GZD3i
otmSmJQswEdQlE4gJpPTI+Rq4chBxCzLO6GFFD3uPT4CHMX9cUA2q00n1SIwoLCq
Q4aQoT2fwBawQZHX36I6juZOWIUC+xQDPc805MH0NijT01Mh4UUqfBTlFgAJga3a
3g6Ze9mbYHRHt+21vkv0ZVpbrbJ+l3T+FCx4JfnQg5TINEJkusMDwEhVYRIbxWYC
zg/tBJ6SDXxryJGRExMUALmadrOqZCK7voQcU/3kPyzZ3G7eFnrZiQ2iZXdQwCeG
sW3vc5Kq27r+Tt42QlrX/PyTnzGl5i/yM6LRNnrITEace9KfZ/tdUUMTtiwLmuBd
qzcWBsAnwRWa4e1C79BlIOa/C5B9H5j54ZTELJtcKvw/4vkpUYOxiyltJ7CWneW2
NQ2Nxnu0VvFRC/Q4K/P5ZDFl+JIIrpk7ZXD5Cks29Xol8orkPM3wHXoQqy/ML/VK
5c7s6YTcB0jB3DlsoCtxEfWmgbF+K5i0YUEgoFeidS0IX1WmqZ9b3/TpjCufoTSi
Y45kH7YvDmioDa1g3C3sgvcfIR31/HLRvBIs2VT1oXG1S87BhoAjNGZuTdcuqJ2e
N+DL6+4MFACLqZ8/xjS6JXfIfv8DRiB21QC+0WgBr7Q7vTX7mrOx7sKWWtA2hrN7
GdyUM800BKDmYrVGa5KqA2RJc1LqF7EUVMHbJujEBlrn93rRVsL6BHyNybDzsc2f
UfvxA0LVAHt0QrF5Z+TmwQX9cB6VKbH4SOdsDcn4Zq/SzcBreWMpnnwEv4M0Cnal
uHqr0bQQMut30wszOuQA0mAWxuLq5ez6EnNpHyMvxwG84Nc/FHRUGtpB2k5gJnZ3
yuWcN59EwMZ+BgLgHTXo4PEjQFWRjbT89trNYAFGdsFGUIhZncUHMTC3V4fJ/5uO
OPA20DrWOnL8V1EezmU3rKwT8ibkwfanRsbZekgKGqSKEVvwe9S0QT0yDB9qBpPX
/+z+BLpxMKbkZkvwVH4beeZ4FOmvgGYyOrOZM3DqinqiqO5n0EN4OX9nGE84InOq
Karq0khCEZI31X2eovTuKDhvbH1D1yKZETYPLb3EywozTfO5znDJzCD+I17iVg2V
oWrYQkPXssUDk6VjVEOy/8YQX3k/dhzDMvJxcy8L4BL3Scncm48+cRuAZB8pm/CG
VAewidulZ5HLdGwkMxMKX5C3Fb9NnuqnwwHmkhG4TRXaSL7qqphWOHWIY4brx63Y
HvQ4HNQhmsbWIwIeiixws2LXmlNxzKILW1Lc015E+kQGE0piT8F+W+m8FGFGCTrY
CGHIQeJktogu+BJedC7Az6ywagkVv+tWGLdv5Hpssnk=
`pragma protect end_protected
