// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:55 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sNw6zNzZkf82CxMvTsf/KAHyWaSIbnxYFPnydKfmUkUtcS1gLG4MyKOTwDA+L0lK
oJmwzSVnsUhHMqW7UBWJWy64qS5H9dVpm0NMl/isRoULPr+3YxC7JsK2jWS58Qzh
AzDN8aRl3ctXar2a7J77EouMU2vL8EfPiUtfLzX7/Z0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17296)
TIuIBErzFISHKz9QQigqcKElKVR48sGHb+R6Qckhdgb4+8wjwzg0nAJTLHTjjTzG
iRrfW/LovZ2HWXpperVvFm+hb4t7Q4mFBxxcu7++MGdciB4wDQczGeCfa3n/Q5OJ
UFi3WRVu/sDkNFvlYtAPhsys/A9MNmfIMDtDTJGl0kuPz2XslpJUqC6WmcfuJa99
eDBIcpzRfvFS3WfZXFpOGjQrS4HY66U09+MpW/24ynj3D8W20YR5Eq9kBdiVoMEq
8zIeRwdThJ7fMBQDnZfzv3BhK4T7JNR08CMKNuvik3vJ6m9IRrbYtDY/OzN07Snn
m1mOaG+m3Sw8M1C9Bot/VxYLT4GtZDmTH9fW50Jn6mgyUjHPJasWtToXfSkZmTbM
asABhB4VYSigugWwzaQf/lQxFpIAmhRneClIq0soz7sqSzRgOr6irY8sasJIrI2Z
i8xYQr1gjfZafzmvFoT2GSVpt5OcmvyalqWMNkzEoDGKcb+6OAVpo0YMm5nEeOLi
J9eafkTxt6yNfN2vcyPW1jn52yBZh5WUr70qawqJeAoYCDXnldyw3fWa0CZYKtHH
Ck5xLWJyy43d9TJkyjVj4a074K1ZJbs9d3vZafkXPJOPFK9cqhIf/KaR+NQXilme
jfarMw9dCaBIZgfcA1fRDmZ5Dh31pW+l8HRcxAyQonH9EOeiomX6+yvtO5rHEMl3
L0YR8cMYKZpib6DOpbZfwn3Q5Pslh58werx1N/fm5Hb826s3r43pXhsd/eHY+4+1
2x0SQkfsA0CzP3Lbjmu0F7PuljnFB4PCfcyaaKFZV19Kl+LHykwF/mA1591FdHMO
dp15Io1LxnkdVN86x2ondv8UUQX+LM4Il76w2FE0TFhOjuNbERQTofdYlygC/EQ9
+Fsc3fv21PXPjG2JHfeeQPIxeEsQIIk0zGHU+4QY8b657erZBSyqsSK8IMJjYlMT
vdUQq9Fjb/4RuqSy31wf2RrcD/2MJhUFBhEqp26IjW/uCoXIGANNqNgr5V4VVCU6
x4idbkMsLY6mT226cenlHJMG1FT7QTNI7LiORzP8kHhuRJlUWvYnKHFKOygKjGmC
d0Ck2blShIHEP2iAy/YBob89M+drlMVNRkTim805bL8ZEQsS12uVrrwJnx2JrVXq
hnAKs2ee5o1rahND+mZbFNRqWqHVm33fJJhsojRK80bmoCgaj23FMZGLhA/Vpb1z
z1OAJSHqjeky8MWYCawmedyj2AnC8ic2PKwyeDuJlgOpwf+3gMtVH0+1Y/pEGJ6p
NjQrDFQHzQ2UgxBBs+r8ollOHEY9319InDn5uMy4uDBOieqOjQK/O3QjDOwaOAnD
GVzP2T3ZAH6F9jLBV/Ub3ok9gSEX8UHEw1NMg/hZ6GjmUOdL3g5UJUxW+TahdoFm
MPP0cyqWSA+Rjrkequg6+EH2ttTPZl4P06OTSTCWm05VFxvdvpOG0/wqpNqMNC0Q
NP1p+xP+qxx6Ows1cf/gRbwWXgAfh/kcDQgJxIDo3Uu8HN6gVL3lTAZsBYeSIg0g
aQg4yylFnU8ynVYoDs750/W1AaJB9i1soLKPIXzxKt94z39bTz8UwO93X0NeIn/P
EXqq3yvdaonK8/juCaETBd7jPXGEglHLCz/iP8ujOhCcWSQkuH3DF798jsYc7xFz
Z3YgJQE12aaaA+RWkBFYGl7WSa/njTobT7ntpiYOcwntJwd+MU6QHUAv8Rb5I4vx
9MWMzsCglLhkvN1SR3I8qWs6BrSlJeKyZKi1f4IUG25ZlC6FkDpPmbbCnpxYn3yF
et3bswX+N04iprhockAZvRqx05kvJTM4xFrdK9apxGIYb38M8e2ohL2LbaEuGoK0
3rjDL13Zy1Gln0YMSXd1abuIflpOecsQw+K/JnyJNzIb4GTMHcpxsHUPiBZKuata
K9540dfdK8zpkuPTX1x0uHWaf9AaN4EG9BBy7oqQ1vol+vUH3YzXeFJU0OKn7VHf
6mPo9USPFYf2E1u67TvLMDORLx/5D+BubERKBOlqmgiPiUd5o08Jgdv68qBZPDFz
wB0/Cq7U3ZXL8buyF0w5HRnd3LnSFtG/InyWmoJDGlaXxECrlF4hYtEe2Yv2qn3a
rHszmx5T8oFzDmvg+Nujh5+2L2gQq0q1FA1kz23UfGmdWN/JJaSglGT7Br/j2rO6
fVqmzruHgut+lLQyqO4phxciBxrSkTw+YrTc049omTfUW2RRw4l7U6pPBRe+gBJc
KjgvWwcfB8oOrc5DVopCI6IoY3l1OU8zomAV2hpUN3vzDCLTRj32k0SNiHU1kSvt
nKGB6kG6mQqRHI1ysfMzfVCSYXf98TTHOXEbNiaKOHujBZc9tCI1oAHYd59hv3lu
kU9c8USz/GI/lAAtYhhoXLkYUSz8marEDmm3lmnfipxqYIUQwYt/ziKWvtUkifkr
T3en0baSDTHgu35D1ataSHrnVjHFTNJEFvN+UnOo5VRReXDa1/rDORwMHYrHQu/4
rvYt1EySS2cWDF5J53k8nthPoM0kTUCqiIcHorKTfnm/J+fib0gZdxupljPDwxxZ
t0x5bexctskCXIAu7PfWHrQWlyjKOBtr537j7laGkCYYYawnXDVfg7vaUG/5KmWp
Let40rzTKpQDHkYtxnz+rUqU5e1zrWhHuIylXZ5dU3Yq1w2JwHUh0+cJDezs0Mgh
Ymjpbiwtpv+8lJsUGVayxEs6BVjPYRVSNowBOzxpV+l3Gisu/souxqnpMqGH9tq/
zocmw/2C/E61b0r/Tbo7wQJGOIYEIZIb34/UJAu0rr6gBsAMvOZhOtIrSs2Ok/vw
Vb9epPdOsxx7zdnPy8lUA6oiDDJMg6280JHqbr1lsaz+uQjoMV4py87HkZGc+I0l
jBdxzXru5+Jzwiq/Pf1gpWKPYYhqzJCHuVHq071br1gDRcBAQ6y6JqaQZ9EDfnpA
Br2psigR8RtdhXaYHJy9wxpKfjfXkLovVr48dfryv6/YfWqjhl0AS1TvXz4C2BHf
ClmLsVLWfT3oimJKcoLx0CtIg+h42rv2sTdgcmr5qyYNnOzOH6m2T4p56AZEUP9Y
hU+CSVyaiQzT3ttLMh2wP11w628FHeiMkCrZx8HEQkzh1tSiFAtsYGrrXnb0aB1p
veuFE9eyF3QIxuUCevi5+iwB8fBNmoMPgIUyL8bxu5ecBK8dS84xRGXhGnCCmLL8
Waa6IXJVUhWClAvPJMbHSItnDnBxQXrBEPBWLg9FPalHu5IloLmX8+ujiA0kKPMV
QUYBlZVUjK7DgrWXZ0Izc0GFOrAvLuCeBqOrXXI3tvZzxkjq6wBrVrWxM04eIVFW
JWtWVqrHGTY8/nnliTiFl7AUzkdxFvYjwEmYpVdja/PFwsB/GxCSQVqj5KHog1RN
mF4yAYtjMN3kiDFs32z2YyUxbgy5IcBPH/DzF/eIWUaPVLIazP7EYC7mhpxNjNwL
dyDnRZUNSkD3ZToNUJ8S6JpmzpaI1ZBhqGhcErSnDLz2uzBHZ6KZx6XwWQsLY8pN
ZEeTXO3Ns/HrcBdpPHYrliMU+x2wjOfIwnmCRymn9bxmdKTbeC24kz6x83IxpowS
hv5YngTqk1m7d3MEziPC2gmFBGCV5ADLndsehaKtzKnLf9oC5ILdovoiRmD1hOw4
RnY0CXY4QQ3yMQ1FiKNqJBE1YTtffM6Y8EVgvwRTrzmqIJbDY52WMJ59jnyooCi7
kRXiayuldruZjahig6RdOl5QPBz1HxDCMvBJB9j3IY74JIwUJnRoPFCjCQLVBnuU
gy62TpkVflhswxU96vtxvouGO76FA3qiCq2zdoggeSBdY411yMWa3VKVN78FYesK
AuZC0kkKlKj/AMVvAZXRESzr/VCAAiabMp+PYuHEh+TiqMhG6JxeFVRNjts9ZZuW
8vWtpi+DgcpTrugUqcsNC/UJaogdIvIBtg5Kq/kpclLZ+SptjQMdvHqMZbLzTysD
JrCMaUwo9P8sc90Ddj7hrRFPezQbTrOccEdr9LdIARVTumpYlvgRUKsLtqbdAs60
lI1tcN0Oux5K7zZRvUYzK3RTkpBUIjI7OcYDj7HpwqGazZuswkodEgC71+//5Jl3
zJqtvqSB1yvkfF+gpTt3a8nOueBE/SMjhJu3wA1aLO8QsplFULH2cLA5cVx2H5sw
pU50pibw0gUxC6vqA8upoF5ncHSoCD3Pou3cxwWZQevXmBU7fY9Fr4jCQQb9cVWS
sYz/b1wHqBnWjpLWZIpkW615z5JEu/8pU6ASh7JdWJev7RAMQDKMndbJg/YJqjBz
dqNv4gAOLan59RWrXbZXaGOA9ZEt1cfX7H8h1mz+oPf9jClePD5nRzSBZRbs5Pyw
fM0bSSNxRP9ySnB+Xvyd29ZQmS7C7h4g7uOQD3pDYDnWY9AvYBpOOJJWu+CkRgEF
/s3vAA4R7fVPZoIJSujWAqfBaUbacDgyvXEE9rL0TViw5FbBJPIJFVucC6hhF1cX
YDVFxi0q9bJs6a9YuPpguYTnrp4+m++yzN0SWEi0M6Is4gP2vocVotuvWktiIhLx
9ZtmCh/D25TpJNo28O/GirZ39GfDVh3lnK/ogS04U0Gvfv3MAmdbNAgLUu3fGmIH
n5bD+9meRXbgkhUTiRMx8f0AclH+hdo/FFnkuDN3aHVTXTpoRQaglPtWX1YE0zL+
fBQYabPXYrT+bSwlL28oI20t8m+jWuOnqzixMFi6SfStDMEinMSynNLlr2FbNAfl
ZaNUKH+2R3m3rI5l14bHmSkULfSr+T/viX8+2TdNtdoXv+vh3KchptVB38j6OQVr
hJtqZPPCsP89BzdrjGbSyvJ/wM7ZZsF/3iWGxwuQHUzqUdrJDbI504GvYxeQsY3+
yLtkPpASdzp9XFTBSK+tpGegorTbjgcxlQEbrWYRACwqd8nxIBuQsd6LX7JNitoZ
Mo1tyVHOILyW05OrboYxAr1gnUL/6Wra2mjoUVL9PkFGx8dHvSQj4sbOf0p/JDXZ
63Arkp9cZxnJp9HbOGPgtGu43ArFOnKSakzFlj6mw+Gy1HOWh3dWlqoIM9EHGdog
JgxLUDnSPkux0TuSkbdVXo3cgggmonKPc6nGbzF4MN7kt+UAyQiQ0Jcbr1kmFe2X
O3ZSzWQL7o8nxl4YCn1qn8TOmSlhjuzFuRF2G9MjQrZ+2ilGSCjs55bhOq3qAESD
66qxm+GRlQFjmrjUhMo/YbD0JiQOJMMtzxG/ID0F5zGtOuVeQGJl3vlc2jkyOTHc
FLrVUS5eVMVHeVjNpQ5Q8fOsfY+EZJci3g69+V2ZIez5F7aEr7CSBjjaZY7jeoIQ
xlvvrLLWe3qlRGTKn5m+3muiEymoAVwDajYfIPykE7+jLYEEsFPylzW6QZEzEsWE
PUXhsChGkZlpe/DdpCmb9W92+zR4ltNU7FqbQM3yeCLpduhR48cRmPfzhQEhpt2u
i+x6EydhOYlCQAq/KhqZKUrJeqRrHubFFlkIamygoZcHgIHdebgwR6iQt9FUFJjI
7MHNzPkrqHAnLnISK8N+CGQIKA2M8D0y4ywr0mlS+ucrgxR5IL5Fuu03xWFgEtpe
G76oTp1pK+o1Yr2R5zFsYs6bt/kx/aeWk7pFZFj5DaYChzRRpaaEMSJ33ke8qS8r
o/4TFnS5bh9c7F1SBB91BhwUuK3m+0/LarB1g7LF9nP7jbFuHutAvRpAz3za9eF+
Ktcak0SQTidhC94e7qLko8GYl89quX9DebVqY1UsBRdqbv8ZEq554+ifje+khw8A
lRUAqonU/amnXbqJ9oAC6q/bpv0z6ZsauL4E8hVO66fMGdr1bouWXE5KOkEvtHgT
s/IsjSiJ0kOxNP0bPDLP2a9iLUeJtSyJWF1uu7BOTwe9LbVW7I+LL31fByArzYMk
d6dz2VywCphpESGh6UQdRyqFcfsvUlD2p1nCNvGXhKUWvJAn3pxkGmVHQ1yFCwDS
wpmj6+SRhAtF6a8zFctvU8w4KR2H5RL18rPeQgEdkyacxxeaEKTLnN6nbf7VW8/d
pyNNgKAkrCGCvOeAYp3gPFYM0qqE4ngwJvxmdMCyleuJMeWErVfb/OoByP+YNm/T
1iNJaVW07GpBtsShQkQikgmUVQ0xuuAO93wOIMao00fer96DmJkt2xTcnb6swF9Z
/w871Ridzy714ZzcFw5MEav4Bod4kY47TmHXMrKkZU4EAWVskH4PbQjW9hOitRGo
h41XmGqzysHg84V7JPs78givjC3+eZZusLgJ0PutcceUwpzZYM8tQNOPctdoy2YE
symij/yNllaDk2JvMCQQT6+dsZ0rAh47LC4uKJB/EKpQT1ID+c4out2RUrRdDZIQ
BcT1b2/xqd8f54Qh/lgtngYghvwQvhnWcXx3LAPiBo+X8mxcIxQwuZ7CYQ6Y89kx
vBJDLlt8/QqdS/2CzU4DLTewtTxk70qJ+uQNhXiLgBtf+oHT0xEo+jINdsfPe7o4
HbXAOpXMnLTYJL/PP2JaXiPur2ZrG8+nthTMwqj/reW7VTnOUaREy05LjiStlZft
p44VqasHVPmRpXJDOKQbnmZgkNcE3XMZ5D5I8J7JGi2rgTCNDybCwdcGnXuqYE01
uh6LSVOGVLswtivb35EUUOgsC8IMKFyB0hKn23XRcoeraQFqbhvJA3PbKlpND3ou
KPSJYGADp24TubHDIbNYtMgTrf7qfYLMZ/8RZPbcyzqN3x0U2lnQfIE3F/ntmI91
qxeOKP6ebPTu5aqyO8SzL9pW2aVGJI/+e7DYtCjqFMuFueI62G0FbbwVUe+OfY2r
WRHTlIjnNhA2FWArE/k0d09RxQgyFYeJXYtjUXCibxxYm3orsICrUh4yk1PG5LSt
ppbbd1NoGqmKkxVbobRRHW9KiKfh5D9mQla0E8SZMWUx7UKXpQNq753lk8jwWmT2
ZFaBnp8l2fguAguVvkkSaP6lLa6ij5LQbVJbozOrUSw1Yony90CuqcoIGNpcP/pt
HAmnH0eY11KfkZcLUMG4J+bKS4OUI5x0nvogSx9lXbAfIUPSneFW+xpShIZ98K55
1X4Zl2vGmbLIBl8wH66V5NnH/DQqktj99SI6q9h0FPBh4QFWxw3nimHPpOJACL5d
Y/v8RlDlbquu5dIu9oESxBcqeHz3mnuOIqY3DZv9AksaCrKUI/y7Xi3fKNdw9BMA
7emPMB+dXYsE9dodEHThwaiPoHYsq+6/S5T/igaB/UNjy77sz1mPMVeU58dumeAy
Z3njELpL+LM2aIXiK3LDjOcwZ6jc5bT0K0V3eAfOvCKm7O2gbvx8WrT1SGH6+p1M
+0QAaNOY3hSD2VhKCCyDysbk+jbT1mkoVXmElgzmUwrdRL6DbSkTtUmFAa6Cpp1T
J/7t3CwuIJ1U8nSPKpLfsuOyIjNm1pL5mFH2Fit4dI5F6A0IdXLZF/FnbTrcFMEC
OiWq+SORDMmOi5InDvhqRGLBD2RqAWzJTAG6m+so39WpHL3RkFOcRVseccF/3Ymb
GSjrueHKbdbwag3hbL8Xmq/dpWjAPAjgPKgWGaLRDgWRLXYiWkckv/0wM9EDLTD6
GGbauylHxobkklrJgjypu8d1iSf545DldC8/VsetZVm1z0zFWMsp212VYi8yj0DI
SqXUdpLknLTlWsPM5zwk95uvEW071tFDYcVEZ4wdMoPc4pNo1QuYC01YdtDOt8OA
rip6H+dpb9OTtcm2GPIxk82NktLWFqtTql2QckWBIGAnoHDl5jBMsi+L+IrolhGE
0FWi7GxDMf3O/kYO9nbCX6XupEbDJip7jGiG61jWKfAMJAxeqwltosQunDNlAjGh
pNh7HJYDq5Syu0Vj/3n1pmk2myc4qFPILaW0LtTMmf86rDuXfL7kA7nBTpzm/4iz
WPowauvI+1ft95W+/KIZ49v+qJpNCcj29VeHtvjDY1OjPvCqd6efHePRO5egihzQ
tq7IvBmNsLVyEAWQ09mzgcza5t3zYfvm/29AWpzd6+DfuDHBXe720HkxZteNjJJv
pRqUNIO2C635mOUFgzLqbYKMqIdColD7hTkEH6MicIxmNjk1PxGf0KWa6a6dgNqs
9o/jFMxKZ+6pZPJ1cnxwB3UhXKOhG0G3R1k4adC8RFEqhoKCSC86j7+AEih8MS8S
czqEmjox/7X7SqYWMJHx3nngr03ukMxpmSBFdarDvck45eBO7o3dR/EVoQqYP41A
MOvNI60whaDiI/H3lbq0DOr4l+IX9QDAhdAitM4xLGFC1oQGf24zs5lcyGu/308a
VK/m86uRUOnQN+yozP917BF+3fLGJTcP7nXyTp/shqkYKrBeFCn1ukhKAcKAbv+E
XDAZ4CF+b7xCnEcgWp/DD2HEjz4EbBdQ9V9yNCv+DFwiI22sjOkFhKTq+W6gWQH0
gSKv8LARP4XUzsdl2ggkFmEKTIaTOctNHyBjIfSEi+DRPrM5/IucHbTlNUHunSJ3
qzjC0dNpgYcji5DHq3BHKKQqDNAqSDnQWtpimXQVhnc0bmbLhe5hniRSYIzYdM1i
o+6wLgKIR9RB+i5RsHXP/wxaIb/DFSfy1gXC+x7XuELjUp5RXBf6yiijNLucnYWp
n0M+WP1hNDq8mpHgM1xRw1cvwOSBb72CGjHIpFwlnvAyMB8a+NXvGhcMuWOUgB0c
i5qDBFhJc5om/wTy9c4ab+3bC+hYB96TvDG1ufQrxDoedytHpwzb9gHBdaG66Iy/
py6NoIDyhlMsBoypaDjMFREmiweUwMUbkJ8hROjYMGCDskym9I2xnxfOq0WLzb3q
+uESycNHWInsvOPDQy4GdO5A7H/8OEmXH9vKyOfwz1VqLe22vcCVGBMaB3ef8KJE
6Kp0AFMX+UWzyaZ92jI3IfZKoOheJmgDRY9hGy+8ySb4YNxDPAHbvh/Is887mdoy
1Xv5TO+onVC903/o7aPGOIrPgXrJ6wTgAmnkDkGjUpc8FXcQCdQSOJHtT4VLOLko
IdnHNhzxJq0BiD+/munrU6N9ZPtDns5gLTnNIOO1QtB/4xPsPsobV/iamYxzy3aK
+a4ufrf8SYSAVgyCR1ch6NOVA6WcB4SN0ARSEWxAlJSjnpPxEwNMBXGvcR/kWa6f
qLB8e7F2h2BLBy6+EV7N0z5fd2ttQwXGTjcBIJr4rBIspP4oaMCkiA8/pM3PUfYK
HVV5mDTb22D/ckJUO4Du2kXkexdbed4IVuyUtS0dsrc3CN+j0ZbvW0ktW81oyBfj
m1a0xt6cf9DsB5hXrarWaAPVUb0ojVNRRVTCHKpWbEj8E58evITmxZEP5gB7Wyuz
W/gly3cxPc/vZTzeIlGNXfTPEzwnozA16ZpRVBftnAMGyiUtGih+4lMC+9Kg2e9E
ZcTBgnHc0FdvSiggmx6CQLktJEc0GjXzHRuHWIa7b96dlBcBY2ynzHFG6GJiz7Fb
/CXiBRQIaePGgSaV86tt5QpdF3HKbIxoEwhywNzrKnoalrvRFJUpBx9jUd5RsqOC
vTWfwvwulcxskXjF006vhINq5TABzxAX+ZDIp1mHGz7qG7TX914sNWL9r9pUEel0
7LiXRWkMLLkL60Um2bOPH5KvO61zpVonn6nnXYIXRLtUS4kXaY0N1wgXbDdxAXr+
z8Jp0xsRGkYf5rETrHfpK0ZvxnTGXOide7iWiUsed4ju45i8EuQmaTl6Wz4Ii38n
iepT/6P8Lf6NAc++1x9twTMAY7lDMU3SO3W/pSt1COtnRvWumtwYajXziml6rBnx
o+Xd3Hvtk8r03is3rU0EO26Irvs+d/fqoQnvzIoRdn2L4R+yQz9bP3N4kCjRNOlx
VQ2ycDlrPsgNSdgC870aGSUO7Afhlk7vWrmW1hQhK5jW7s8t/SZJWbaH/pqIM4dr
DNRBxXXPwBui5fvt2Q082nvpc7Fk3Fi9/e3MzIyuk9VrsY3j+tiJFT/EQMtQhkmI
DaOI9sDi6yUIe/DTs0wc9XfkSpb0AH9SxPLDe3cTkkFKA+LTSBASehDDFuf/cOX2
/aF0TwD9nFlgeLhtPQOZ1/WIwhFdhkLakVpzUw45zCmv/KqC9x5cclCNWXd6Zeue
FZHQEVILmsB3uqVUVR9Et94oic8QXPvslZLMLsop2vofyHuJq35tmbitb2u5anAL
Yz0HV/j6iWf6JjSnhK9RKbZT5nXo0uKXdvIGKVvpTEA2WKEkTxX0vNnOuUImoIL9
ElRe53J/76fMF/P2zT5NQwKdMKU1ifqGEAZtBODib5aNzjCocOeMy4oiIOM1RjYU
ZtHvqWayLu1GWihTv6COvLvd2UJLOdYTSG8aTje7vK6elPWt4vUuh+102gmhTd8A
QczKxh5izZdyt55DKG2zJRx8gTth3FjvZcz4bFWzOWZVcjyoOHerALOfgnAEYKVA
qreJsA3MAZnk+h5hYrLLf/UKuuS8J7PVmLlA7y4TwMa/7CGsdwF/upNzuiy4RCTz
/o+dsjEfsAKzL6EeArEOSiL3tzNN7Nz85GNXoOnwhVCN/huSP3yhs+io5lDRHX+E
aPTtYaKzCdNAwA3PvvdEARe7FQUNimz2OW7rVMh6yfbGEukPUT0QcmNj7b16U73m
C2o6yKedAUi8FWlwJ2xtoDuXA0UC2tmY8uUh5rDebunM5KzCcz9Gwmk2hXrdBMfw
leTj4QMmR0K3o8ULbz/C9fL63dUQmNsn5BgVU2haZF09warsI1DDBvFWGGMZ0/J6
fnRmuatBMg/uR9ma39JqN5ZDAawvMbFs7SitdSeIXDTZlVqDsiJez30fsXWU+a2w
a7ohchvcoULuzrTHw8X/beE63DwkIht4DadqTeOumfjcWgC+3m0ohto3sjhM9TLJ
wTw9+9DCUQXNFq9KAfFZ+v4nNwNb6Xyq8c/xxhXsMHP0NwOhnenZhTzkc8dIIdOe
rwEDFhcOQ39LnUjR3krflhX7ehWldq9AdrA7RWN0la917GcxvU1z8rNkikQ/VXRa
g22zyoA8ekQas1yFqOBF6uWoBsB8WMyaHeLKhFZkR9Sb4DHFjq9bd7cqgca7D8Pe
k2xoCJcoUM30UBkubNFS82eRPRoQkXs7K8Oe5GjQm8KcuYF4yW4gekGqBGPWdiej
vsD0Y2DdMrBGq7G/XrxW3zBzxAMbZhgAwMd0bzWu8/w9EhffEK4/IzCnvC18Nt6e
tZ4h9aTdU09RZC7sup3T2ZjNqQ949DyIhovkqKXAGUI2qFnUppoOGYklNf3SLAte
NrTODz2qEO7wX6oCW/EK0Xaqc38GFjwU9/EZh8oqoRhtSrI+aEsoAFgr8Vj5idDf
9bHFIVuh8C7sw7a1fc+lPsdRYDBOE4hArGDKr/p2c1wvfgIXhdLRk3hBl6m8uuNC
Iu9U2dlf8QimmclwS/YQjy8+erdwyq4KAcpDz+kS8bCOHfpD9KNuwZt913Hbjtq1
YgOQN3QjeX5v17aj3f/vxsRgN2/G7lXng0gOa3SUjCIAW2rkiR91Ep050DdJBqKX
y8CxDgxfo8BF53djGgVLoyy/QLt/70PNejQ1PjW0zmFkE+OiFLx8RWUBlnFgifKq
r6EnVbvvRu5OfiZ/If5V4JJHuWk/kx2SGWPa94abR+K9NMkZ+rCDF9NcfkJbVxDn
cs7lhYlG4D9QVoqyglW/3lZeflXhmgC+NhxHvUEg16ZQTqIWb602lqnORj+CRmei
dn/oa4msdQHUBrMVdUHQjoMaurGZYhCgFKpWaVd2q3cePDowxZ32DGNDJ9Y1Zr6m
/ATIkWIDZviEZ7h/LCqdRbtVOwgg0bb1MVfFIzWsp7cFXWsRFlyaGveL/uc77U26
UeTtSANedcQ8CatH4Lm3GNCbXVdHxrrpGytUovYVyr6wauK2IhBY8S5e3naNGchW
72JpqAOJWJ4hHED74HA6Qt8JI4cPhTWQOgCrvsJvrBAlhUFZjKSmzYpd3ynjcydI
Y8C7hOPXyLAwniIW9x1ItqK2HUW3sIXkUeVWrkF6PSDiPSQt0ucI7tfi0dHvcDBV
UqHKO8wpJqwQU3N9TBFO6CY1B4h6NbxqbiEyZUeQUMQi2/O/ME7DwvGfxJFstc1p
UAUkX/mGxjCd8H4XM9cTjBwJMOeBXcX1VKbPvt1x9Uoj4D+zEiPRGWGzfgZGypRE
67/UnFHyr7Z5L4gTXCjJSULnulTOxY4FTt4x5fxoTWh/Ycv2dE1YFWA7HfoIec1a
vq2T8G+7fVI/AijtfuSGgtan/cX962+I81Jxz7SnE4ct/OhEqMLLfL9zdjHXMetz
JIAJvmrSglEqfc7a0YkuA774uZ6pHxWnCW28dcyk0j4kLnvmo5QEmYm1eN8qy9M2
Bx8cj5lYwSsHXYM62qOJ2PsuWG8FdVSFsWIbGnGKNLvZo8WbkmZxhFyqj+/zsLOp
dSM1Wpxy5y9xFJjxyilUKkCshrsa/AWeDJsd6gBTRMghgEZc8TI5DsmAmOXkgrtj
UGxuVQdW/ZOsYtbEZ0puk/zVxtRErISn/L6++xLnzYfFBor7zo8G+G1m7emefC21
ewHcECurvS6zToytitSebfEpSpsFQ50X4HGZRjJjozcYVTUCGYH9ZI1B0BQz1Q2O
F07hyWSfgcsh1Hm9hEupub/yQArCo1IC5gGdakQuUSjVTlin031dO1tIs9DrJnFe
o2ZXtRqQXk4c+uGKlZtOFU1lO20J349fWswB1LtoYyzA7n5m3SCFiG4Kpn/8anN8
YUBjqek8584Yz4bm8z+GiixExc6mtuszNlbJdtCy1LMIZYC4j4wq7X+u/TEn3oAS
l7CMehnTV6+sVnyDcpdOgjpIL35pi5ayNZ90vCavRjnjdycemwEbA90vmgJ0l9Er
nSmdYVT/quezmHMqk1k/NXPCCiXgSjNmwFx05K/HVck/DQ2P4EdRw8Ke5aJD3hRO
pLJZGe3z2cDkJbfFn2zIOYGD0V/nq9NcfJNPsqNzsuy6EiuiaMEYYjHBdOO18kgb
sOrJw6JRDxoyGCeWXDWjduedeSICQosYOkUfVUqFMa1OMyMljmg9cEFb2gcoHoui
zMBa/CL+d4lZ58NuWqP/LpckF1H2sq/wRlg2AnpM9SPK9pncDGxtlKenThH2x77O
IeLs0X+J6EVJNlNus4Hds61PAoKwK3WQUEaDoXXJnH7Eox8hVBqJ6gKYyxcW4is3
0WODKAfUOGSE5RQiaDsgCo6IDlgh5vYtnc3LONpy6qkHLLFoAoaam3x6Mrm7HOh8
KIKnQ3lY01tWG8qekeGU92gj/8nY6Zo6tciOUbQOcP+L/zJI9hh0/V+NZjCKPJ59
2dvpOURtPtsRf4Gx0gR404ynOxfXACNlVQZWbAoboHgDPWYCTQb0LD0inok92WmF
Qm2NV856sgFgjM2c+qlz7VxH2H5gJaIBxjyZNPE3xjtGCHayyCeWV7RUV3+jJHah
3gNEQoshhzC/NF76Sa3cSmnvMBB3OWyjGtUUXdMrPgH/2xlWquo8BMOvW67dQc77
iPK0rDi+H6w/5sVVO9aCtWUq14biO8HZEvlAGtvBQB7cfhPTzOXXHru6HWY3vXtG
67nFCEFgThdLCTA8TgeYwPdpBt9ThD8MdSWm5L8tI8em6vMELka3FmUe24VnDlAG
/D7y//y945qL8pjlERZqpFG17yeaoGqu5jrd3NFZMR5MTVsI2L5vna+IDuZGVUQi
2Bftw55DiFewImdq72P9lmVhTV0bcoATVpoIuwzi0l7ca3TgPVpXtwsW/JSA6gs0
MWsJ9bO2pIdtmpZ4n77rsPfw8raaJ/z473xq+61HmRSrGCAzb1wrQOPmAkLgfD75
K5N7+GUYqq2r53MUF0+8M8qzK09Yhzt4GuJhXR0iAe6SexFc8ephee5s0ClY7MvR
1qjMYWFynrTY4NhsHHjbDKaqpaRlZYtuz9DR1PYMOnnxYcMjLmT7Wm4HonxYeXgn
nF8f6QQmm2l/AnI1Ll1uYuPT4igto8xMWSvDI9PPp0ztOgijXPr/X9fdG4LNMEeV
o5pcDPOxrBndBlHXVlBI/In8srSSIyHx9SsyJ5UpR+BTcU0YyINm+vOa+ORlXoH6
8lwjxCQXkAds3UanftYFnKn+HdvLdMeMMC4F0YSgFjMWDfwGToi4XezysVg49QDQ
+4r7XLy4vOVcm0yxtYvm9VZWySV9lbB8tmy8o5yvJ2OXrV8mGvzWmDJxmEhKVgRZ
nbRgcdZ+4ou3Efw2xEh3HGG5zzZTuoaXrggqZoY1B+j5H2OvjZlMCuEhUXQUxfZr
tCmhTUXkM3U+LjvJB4oZVRufGIW0F+3WH5hnDna8SmAO1gvZTQoZ/egpKmje3Rxx
5jX2w7EwU5Gjk/I0/SYWD5DRJBi9IX1IqdTR4caiQY4fYLhXABhHiXuZKwvexsYI
bhQHG0+UgC83rX8xLN7oXcWPaiPMJB3pgLCDSyZeajZSJiR9QSuoRupv3IeVzbWL
ptH/3fvdIIGDMIZSkdIdoXXGZoRMAEzKJ6/ZpROgJ5CDXBINYPbW0AXOFuDHWSxr
N4UpjaZNNd5BvHY7Gq6jBfjOME+st/LezQ3ZhxjXEv30+rBeWS//k+6jbV6/kDeP
sJHxUX6w0j5SPmLoTCpY5PElhBauX1Gn4c3z0Xbx64lU8GtanJsIMXG0InXl+w3t
6PBJvhh6dh3P/RjGbHD8th/On0hTyT6xj/uesvy0+2vyUQsWgONklrN0+eAkW/5W
fNVRGKzrs0zzf+9aVbALPK9+epLRdaJz+/tyKnYct4tj9fqygynH40xNazpunKQT
OGawt8Qr6udhDg+UvHxxQ9dn+hX/epK2ywlDL0DQCLwYiHU0SE+TwuIUW7haN9LD
lg1V/ODc9mJC6HhzsrtAZszRZ3CndPKl75tZiK6RGmYiJnF2NpWFMi+vkMCCAq+F
V91uYnjfls2DE2CznR2X/VAkv70DQmvxo2PIIPv+BybHD0Sitvud3OEk8OEqXQEp
ElBslZLiK9Mm6u5IRU6GkeBbu/f1MpbPZ+H4cdFaXniPSQMgVgbVD5Mk8xUg0NsO
WCSn4P0CPv1L7zcEejmbQGiZNseEfP/5jyOEnUo4Tsr5j3LqX0CiBOjyM2CB38Dy
QDQUKovAa1zWJiXPAx66IHwtC3wN4ekUc9iBCLjD6aK8ibgun5TnN0st0i2++Wz+
+qw528kW0virlmBYqylmmH8VGEBH2np0+8CqxKrsciqPXbJLlUHIvWLP7jSktNY1
ir3Nf3tSfZDDl4PN69Latwvavg6sEO7kho6dnUv4MZmRoTrMe5uKulCFOmxeUinC
wmLVmdFAkSDl/TkS8NslB6PdfpW0ZKNFI0tMrDS5dQLaJjhfBMIDJipoxCS2hxzw
zI9giEtLrRZ8y0ZOcwIGMiR/XpbQikFkpY8yOkO3HLSX1tR6b6bO7CFRA8EbVMTb
HUGg3WFl5+7MS4kMDOFeXsEFyk4i7LGPPwebLR4F+XAiB/FoCHtsd50HXzm8WXc+
HNSToPAlQeni5/Ex4xX56puRwO7Jf2w+abe/QTsTb85jKKxO22YsyXoZQ9crwXtz
p1a42+EJAc66v9G/xLzLNMxaFS7gxM5/O4X/W5wFBADjp9QinbkRrEZ1NXbFbu+6
7vs1WigCtEeLdvWG/QaKYc4n1qQnqGJzSo++sb4C3/9a3kZFpZTt9DBCT8/3HksQ
9nZ8V+gJeZDZ/DGCMvx0MjFkTGfzu5Z+p7argF0V0SmFYa0RktA7zx49dIXQt+3U
xgMvYK4Rx6uAeLAZCWyO1TT9mDYhrSPQ4GIizePUUhngtmjNHXDsXUGhOoYonV86
3NUPArTFlFVujLM2OZ8ikpgPxNrJoXHWyRN8mUQzx1qhlCQcEBBAHZo2WH8qxnWJ
+dLt3zosrz/faJw8AjrMQdvJfAKJkaPvENSMR+i7NOBhLZfNk/tVUYx8b09A/TTB
+Px1KGHmdYUarptyqXW2dWgbUhKXq2pdwb6udZSahpIwOXrQOzFGaIkt4/zZiAbb
tbJI5KegH3OSHfGEj5a6zS84QDZ0wIklH7QC0ub81+dS3BFW8DZOaLzBsrHPFqtx
7zrkaXczh0Q3j4l9Y/EeZfnYmS+9tlWRtJLbvRqtJz4dYi+QiABbSCYAmmJlgPp2
21mkGojbGIhL6FSiNOV2JeMDmepQcCOCMh85U1nGGHKQDPTGDtrdnlEfYmEGUDnW
9CymCTSpK5wB+uq/YKe11rZasyhvDr38FMhk+L9hx5sCOPQ+BuBcj/4rYYb0NMj6
asXY+ZCCn7NboFKIceFa9+CPRL0hoR5oOgieG6lCy+AM7Cd7SfuG/s9WjlU/Dq/V
76gucbIGO+imdVdSQstPdQwozf7xn2Nnqi6PJrxxbVMAhBlngLjtTcY4A7sAQ6sv
NiN7tk8BfN4anejvvb/q6nc6ug1oBSQHjkrWyzk12VD/5O8SBsBFjmRr2izp7+LP
XyQ1xIPxoaED2Hj3M2Foa/O1IlUknXC0oEbTX90FHdtismzJ8JDdXW5RGFDh5U3K
/g31bxjgivxelFXzj8IadGv+/op3zOAWllqCxjXRbCHR14CYhb6xSTwg5a+qCQCp
vcOOdZgpqidB1FBVeDaUIk/T1cwfRCeOK7Ii+85pQgcZ/Kjly0QDku+t7b3yNz3P
WiwxYqA2t41/2ckGIC0oKAoWMHK6bZPoRf5rMmv1KjMnO6YQUT7iDVkpPc4OU0Ls
7r5C2WBM3FB7WAudqLS1Jpl7BCOhuCE0CAV1VOTfIr5YfTTQ9EhF87aZfEq7C33a
20U/wzzP0NLah1+Dlm6CoO37JfctE8AEGjlb1+yrtByJq5sKim8LbkIOc6YHf6P3
nUeR1OmKxOdKhB2fRQwV4esT9FpKDi+FrRJRRqoEugrf0NffNTA+YD5HBbP7FORE
MjolXpECC1iPVQEegOW5ZAgKnBlJ7UxAhZhIj9QV4WJON+XRhsv5VlUirucvHyoG
lskS3d5vek0hOLuo78bABp6IaX3S6iM6jrA9Q6h5pSGfdcnX8ljdiS5d2psRMwsf
+5txcmjQ1C1dZGYaMa8D45jIFSa6qmenWg7a46FesF+zuZVlW26DhODmfuEgrAW4
y1+nnBoujyB5Hhzqi4LgqMF0THflcUI0aJeWeEX4A/mm77cTM9zrhNmf1yvHjtYK
dfwNoMV6ern3msVyYwp0nPg9b4THlKo5fBROy+X0XhTu0s7lWRjNK6D74n7Ho9gj
lK7vFbmBPI6RtT4r62wRsfiPRukQW9y5WRlvi83YNha+vAb3UVzm9prmQslwZ3gm
B0NgS9aFbHiYPLYtP18YAyKyB6XPXIEj1NQzpl1VjSOpaeQecFec6fnVt0COVC1S
AF9+RqSWU/qXok37TJCVbrhMigkm8IsGyxEM/YXvcdk4M1zjaixSqSxlW96Km+jl
mLH4tFvbq2bYYHx2TAJr0XHma9gu219MdVNq1OMkv8bHJxxjrPEXpEBR4RQB7XZW
zzMCiHeN0X851RlF2EUM3HK2lMpLdUwmY8OnNhi0zKBP7D/DZKlG8Xo1G9fvI7dg
74Ihx1acy8xCgLpn4LYQaQ6HBT1IzK01Cwz9urp0tdp9LQL+nWLZghKElUAwEb3k
CHlxfakghDqT874RDV6+VDhrbfsUCt/fm/iLVJw8iQlqL8fzVb7x9/BcabftgRUy
7T0wcKpN5Pnln9nf88I057dRhHd0oadqwrvE3AfdUMynedmu4oyGhusuDwmEfkMC
RT0umQh12Ls+L3GUZ+vB3irS6a107H1O+LMVWTNJE4vPb09kGDF3v7OWlJ6Tdjl+
oLqTSMq8wqXC7pAhhjlsfjm9M1/XcL6JlpKSvNTpWlYbiPXKtaxXpnwot1+GpI6O
ueXkIKOGYL4smIb0NfH6LxXyFjnCY8FFcB9cXKRj67h9fxhKBXOBgmh3EbllUdhz
uf8FdCwCYSvIp/GxAJ4+WUrPgO5rrcsFgMmfy0RvcHRQ5twu4TjIbEaJmGyTYHJy
uNM4roUE8fdSqWJpJU2rC22PZKZtcv7VZy6VI0QxgYi21kg8mUTTRitUSUOTaWi9
5Q4rkKtsSIGpKdg+tjhu2pWMDb3UdxfOHdWcVWuX4Q2RhAzW7c4FPpfJEnx4KUsx
6MmkqT5pYmv5EyD1Qsr/wbsxnBazZxqfhGnmBIv8ftTJsLB8R1eFWk2GgfCg0gAO
4nKlBCWKPFZ9IDg23VNHS7WOLwLwMzraVf/nWNWBXQx2qBEYFvYjiPRJv230Shi1
Oqgb0bxQQ6cBkM71UII5UaOHrRIwx7jhBiJJ3sfYLKX0C+8qWR4aADk6fBQ/BGU3
noaQ1ILVTTX6CAmdL1Esn+znxj9po8+rWy/M4o+jIlAlQ/BmUyWEam4AYAyze9MS
nc/E/tpWk9BZoHIazNLL3SCp5T3x+8u2UuzmOAt4da5bKfufKIUox7JHUI98cDlL
t/8mMbVHBm2B6AivjK3nWGOphjBrTNegFDNZSedh/UabHESdXOrRQesYnH81KHuN
9FMV9M2hEC+UdJBtCfyadKP6Nj6ixLu4m8oHIOCzzEmJB0S4fs9SiamHP17Ow8wr
oYD5Sx/glJuDobYXSAflBvQvtWRof1BdbdCg9+HXQHcCpFmxXiGudpITrH0Eq9+J
uTljoMALrt5Fjfe6HbBX9lBKemhJz2qKtsm/SrHskT9dImIgJjU0UQDZ/N4Q0W9s
a+0UAyRKcOM/MQB5v2j1BF3kxyOnuRzBwjk60io5nTPLPlE/xpQ6JxPuH9RIga8+
CqsmOppsjKNVPEVJgd4grgkljgFw3nN2+PIPz9GkBrljsk3sdliP9sr2tNER0/2E
hgg6jknYhsGo9bC+dPNwbmklbIFKEeFd+jIC+zlXnmHvzH6Df4XYK9DZloF5GamF
SYKjdJEkvfnaTeE66I9jSR69dPsKnjDwByX7ZcbNAPfoHm96n0qAGyS2nJu6xsf5
cuMxslR72UOakcvmZ93MrZXTlIX/I1IwgIEk7/LESWe0MZxAUGHAnhqAtXmpXwU8
DFYa2GZ/TN4DYQeeNYUfww9SkNWd7aQkJo5IpUfSdpH9rZukugnXsmOyBGVqxe16
A8640n1tijHMIEwAFn56xrM+5v8Vlk/namuw0vNJugl5MccbqgIpyJ24sIlLHHb/
QAJBALDle5gLeDlFKNk5bUur+kul3LeFYWJmhpp8bxskcYXFHmtEoTfm79XrDqJo
Je+YWPeyYmLXi9ZBn/JVzO6ujI25Adt6NrhpF1PeWhsB0afmLYupxWDJaEdr7mqa
O/sS1U5DjkuHotJ1QootoSqoO5sU4WTlZRUXNmKyM+OUknwE7xveMsHHh1RrdxWH
Z8E2+22zQe3k7BvcicDMfnit2p0C38Mn8du/dK1hT/alDzzJFBMtwFLfIOC5U6Mh
K+oKMekPRce0A07XsNx/dgHGYR9yxt17irYnSWSGlXs0wCeeV4EHYKE5nQ73+6Sl
58XQGVG7WgSoYF6iOBG/O9CoTU+hGznfjKHfT0p3CUTQ4J84xHDfFS2QfduyqL/8
RIr3SMY83BRLYSwhc7CNV6DynF+ZWmXtfI4shRrh795vF/dkzEupVmD4iuwK8QIO
wIu8J3y+cyv4V/RHKQCNP5OfjkdHishaPmQeaPE3DWi16bbTumqvjq/iI4Ev31oG
hu02jtS7Pm8JMCLav0zFOCxVBIziAijEMu2cJ4CI/48cZbZTemPXwcwvpFTAmYkB
dsUvS++6UNTHrK81p55DIvAqW/YtyrWoawAWhZaGnRXFztE8XhJZj7UHzR+YpKAj
x0bJe+5wagF0wCHNFmCgV0w5cGXJe37xdX29Qprpg7y7D9qCH3ExO5q6hTeOL7am
TqlthCNtjAwSqZKeE3Z96xXbmhaplUW8G7c8VsSNBr6TOcYIAAWv9z6Kgv+zX9TM
6T6Rcd4ahTzTDb+NSyvK1DVDBrxQ6brqtFeuYYEMe2nTeiOB9RqpkaqDUY9F3Ij0
7CJziVT2RXUNfqe2NMoALMUukrZsKcpoQdoR+u1UG0Ixy6b1b5chX/6Sx2Q9RGRe
4loNyetsfKafdDZMrEvRcZ+tu4lmX8z2HIP04zaPv2AR13jgryfsGRtEmk8zZ2U5
8uzEVepq96WJTi6+GzDCA33TAStCYQ32eEdpA9Ifb2YE172SnTjGex8RcpBcEjva
pLOqYmuzNemsN7hYY+YIjCc+YGJB2YM05eUPpGOPiyqkmAhyY0xpTROL8JwpILBM
1xGfSVnGlDrAAkPNhQny/U2pRFQcJzz59WLkWvbd1nIKZjsNPnLvozXFc9JtMhIk
D0rCaHIhgphl4jE+icfVT0mXjpAibf43PqsHzoIQXYLFzIpTXkZGguIDtbt7a7Dj
kG8ma/uCmZyz7fTgk9Ptg6u0uVAeHxkeM8TjgwwhmXVbg66U9WD6yFAknWWwssUu
4uATWOxwmLstOZk/zbM12QRjIwVsoU8m9KLc7sCvbJcKwpsQY3FoXTUjof7/IUz9
3AhqyvPk1lHXS4SyCVYmnT4LUNd4XAKTvo/+NxlFOAT4pwII7k70Ib2o7UUFwWSK
bhhoX9nPO7XVeCUpL02vacx6BztVuIDBGoB9Uar1GLBeYCvx3gq4QrFFCjl99sa5
RnOnVZ4Oeo8w41XQ2zj+aPgTrel9zNQv2ts7ApFg8hDBSzoTx40SUOFKq/JU+k8U
1QdKIiJnH/kXhRczUlIBCtfk7P2Gnq6ITWCAF5lwEoFG4V38d5FVTYeOVMjAHhze
Fw9WKjW7YI9TPv9LhsiiiRaens5hP4Mi31zAfX4VcIFzbO+uKFJrinKlsiFxI6yV
GivhjAeyZI9QA/zZjyM1v2hQL4vdrJUhYTpvs2WCkJCwflUuMaJbWOE+e6SITqz8
WOqTRCuGyjTsURPT9gL0GkrtVvkYY44vL8WCFv6xKv3fv01ZOr29obbSqha4IpDq
DmyWkqUB6mcKsWM/AQotCJTuza1+C7ND97945Oqsrq8JonvWpI8ydP0B8L9F+Thf
GF367YTC+T6NZobGqX+8nMJAg42oqFC414EutSIscLn/e3IyOlqK8jetKjWFxI4R
+w3WPGE75dN5Bl/3B35totNOrOgNWT2+Hpqdn4mTtbA44efGTN1W3KB53fRG+SPV
dwTxQ7h+kOH+q9LAUp3c3CiR98f6v93i8HyUO6HfNXW81P8bk+aGxBKt4LUsKyH0
D2867n23kFYjXx/HRGYglr5g1t5BsQ9csJ8CwhbVZAwGKLGl1F2KMj80S53dCMUH
k+3BdktHyYijwt6W6krVeS6MxrlKkvO6DJXE7RQEdlENLgYLDF759ErgtBCmUQQR
xyxNMw1wFiFAGm9k9vPpPvBXElp0wQzKQbbpnvAvnKgjSwKfBQBGk39HY5O7qaC8
AHP1eHfhlr4dbGEHhkCTZ6g/ZUBwDL7LZgELJp2uirfC66wGXJP/kcgG/JUEcrQ3
e9CkMz7NcIwrYyu/mQjiNzXCrluXpcd3kvHudRKWc/HdHzFKabraAQfs6iZ2LnUV
AZcXvIp2i0o+BkL4WSrcgITukrdUpdgwchS3ULNN9tWJvVFYgG31Y1IIuKUjvsMz
giB98iTQZPU4oRXITSufHQj0Pvhx6VyfcgEwSJGsD/iJ9ZM3ZOHiUb8QRVcALrsA
HjFMhMMV+HCohFoAyJEFLnbUO33mFibkTs4yRJxLtpLtlSPB7nKNRrDhBXgM74pm
LNFqxg9VCx5yd0WnWNdA6Aoi261R7fimUL1C8UvIhGyzezsA9kDoCdxAH29Qna3h
BWlgHF5yGcTsm2fuOLCbtvT6YH480x5Z8r5Nx4LmUZ42kWkrCOaUAw1c3QMNJUIv
qvNLXSBz/qVPDvu8hGeZKCnuLnKPeyxnR7jSWubFGlJ7Rhk5kC2IBMYHmpo0wW2P
Oybg//TTAf5xRqpdOi++WEOHZhkcsNselw7vwilZYCQlibjkinau3O/vDuCFVeHW
EsfYYD2M0KOrqjvm34+zo3ilSipM+ESr6l/v67jrecQovzru51A/2vEKdMtRU6+T
TgUgqVCntrQhKwuVvsk/b+m8PCKNy/6ss64vlBSpG0wZjqPAnHtFyeOfSJu3led2
O8CaLYCaVaEI7kO4A2ZrIY2jXOg5o8RdHrV1Mx1lxosPAI4B5tgUww6PMkZe0uev
NQYAs2B1Qqwj5M0iaPrT6Kk/DV6BcVde7TwS16wtvClo17HUBLUezvdINPiNizq7
hjcQYdZVKbJK7QUdPZQ7DhOISF3BWsUK1sn3PuDbQS3nuhdolER4sCracih6RXOj
V6LBRpDqv1VhkLVWNbZ0IcQFaExCYJc7xK53H57ZlHBRogTgNCi6/6RhduRxsS1T
KOn9+V9Afi6RTqqomC5W9iUVud2/SSqG5Jwy7WTG1Q8yhwtkDxpnAyoUr6sZ49vE
6Ng6QhwZVxEgclTiyb1UvIt+8BLi9rPOngDikxXDBrN5C3hUh727qyzDv8Z+N7S6
D+iUR/rx3H5Ianxn7o7jmxYWMypABUU2mgfyZ50MWCa+PgoTS9SUgzojwOiEYKt4
e/AIgClYxg/BOL9p1BJz3J/wWsghZZDeo02FInjygwTM2OOqGLitimECdpZb6Ji0
BiScCXEIGECIsHI2Z8b08M1kqEqMNTaMggFDZCRS53bU9cO3R6nWHRCJK9UrUai8
8GnM+cE1PIMlfJCugDFl+JehMbGgX8W9mQUWZndQsxxDyOXn4Q9YZ8Jmx9945ccG
RUbliwfVQhcFpoQNfu9C7PFmU0MNZlmS7IfiVLH+NBWoqL8t0PamfoQ5rAXMNkj1
HTzQf6+xSl62rHlE0wklISeluERhcQW0QWi1Nm6Lczlozm9meWKe4jZ3ygselES/
VlyCce1I5SjN77efC5oTGsM/LV0BykBA6EX9FPJrOMRPliQ4nFMv8HchKFyh2uZQ
CbEuUcOwR+f3RWA/0VsRd/28+s2xxNOVFU8yn+OerROryZkUNvvhLonDSibdYaeQ
wJ1BEBB5J9ZjLGR5InQNIIbPwF58VgCq6CA/us6Rc7bdU+TjZSPXScOlYGH+t1as
upibj/RefWsYZArFq/DwcUrLe3h0YXvbNeiteLgfpMj+B8PnomdJei2j9HdkG78H
b1V5YewvddYdzib9vR7kNA==
`pragma protect end_protected
