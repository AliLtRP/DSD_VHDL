// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
CR63QRG4+pMbiU2u0pgd0eWz2YOubxDDbVOceBckONtz3X1hkYDp8U9jEeAHlxtc0dWJcUvhODkk
mUhXCe6Hxkq2OA1AdG52gdBDYO47pMPPueZjtfPZstfjeBh4fO4EgmV+KxrD7ictwFPB3MaXs3zl
qGTD1euyoMMI9dt8ddfLihB6OEhvjRtJc3+OPkyKSu0OQsgLRIiAb1A8mWHlubzmjoIYtDeZ3DXT
RW+2e2mnhY8s37X7iAjrZYv6GlfFXbAaNtAqPHy0PsEgKHL8bBeArXsm5lkvmD9RNZrbL1TVPcHe
rvb6Lf99Ak9KTLUtWSA50GzneNwoGMA4WBPXeg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
WmBWjw1vtkqxikCJbwsnrhGNIw4Xudfddb6qxjWG5uDBA8fWWMK2ZKdbKjWTHyqxC1RW52pWRrsw
4utJOykOtirFpWZNbx+a4oI/QIttlSa2M7q2sTUM4a7ZhMYQaXG3gOA7vVZliYcmlfv/seuNrZBH
H9XzmUdm5qaYZAWq1YPE1mo6p329xrCc+/XwRxJAXN5YuqOmkbD9wQGqNmh3ZiYR40jzj6cK8fqa
OM2BHWYxrL6LkCUD7N5zdc4v3lJvxBvl77/ItACAEc+a3uw21xcOy+9kuYB8feKhdpbgiWKC95Xq
I+DYaql9acC12XraSqnpeqaw8dN+0ueSSeiC0qWfx43dRgD+AZ3ILSzRLXTOoOC7w0QH0XA9aB9+
OUB5Qo/iLpSL0hCLPDYos96D7VvHmikixPqtfnEX9Q95mF67Oil986+M3S+cJKChBfI8QutnN2yx
W7ALxytmtmwqIP1eYDQL9PwJgwjUE6JvcdiBmucQ29GhZtBj1i9VJQpZEhdT+u5wJZ7dYMCVYLa8
CeKBVutC1hqmR9razkBSz1ywjgFSu8m6YOz3KBOSLSvEgPPcXVr2uHpxO6L5iHS8IV9gexBscnxw
iPP96sSFDABgB2i3IG5LjMICyQW+5gtz8XU3Gt45//h/lmMQ3514o46flLutVVNzUkrVBf1ChX4Q
a1I3l5wOOMD6ooaJNB39caQ6p6GJxWgfeOuPVxLOXCL+FJzpApzRLrr2N0T94lYXR3T5yeUqUd0b
XLu28fPC24cx35bAOjTujmjQ/Nf9JW62RNVtIAIiM7K9Y/BYgLGIEiUEzAfPo+KIEiF1s0f2O8My
SHtB11BNpkLf/5dK1SyWbVB1peSa4FHaq1gMnqxzKLnsdu2oYatXvA942ubDIH3jj8b3DJi309MA
eRV9DMfcieubauh85Tmldg2huBrmP4gHU37whphlmGvW6QKU6zD9dfpd/pTkbIFT9MmuYD1MRgTU
LSp4HCmh6FvfxqE7ffgJcdfL+3+vo5YueDaPkGvJBzLa3hIn0iTjdZwaZ5Y2ckpL42E2rnCR00qk
xHFvpvWR0PiZ5AUws6SmBC/RZpNPdiY8/tkBJhp+0pHzi9eHv8mkBw/1UzP0ylZ853xH8Zh5fI/B
ov4uQsIzJ0vIyKCZr6fpwdtOfNvYYlBYO/A54Nndn3ZjjU9AKW5Rfqv6wdKSmhDIk/wZv8yj0pj7
aiSR83BMDH51/OvUWz5+9jEm3ZpJ8w2k6tumBl6XEf0xy2lnkg7Rb6jNrT0Ei3EiPcW1tSCcd1tI
/MQEKl0dI6x/7fUupfmu5mvLaDAk7zHlbedT5b+bIZk+aDvYGefGXd/er42mH7uvysAyvfJ/gMre
v43P/Mwd1NqAXDW3IK9ZV8aolJDdKjZj+nkbIBvodJlMXL7aSm2Mt8KBxNObWXiKks3bgeFTl78i
T77vuMr8Fzo9tpzpae0sJI3wtiNSCmRsJexLT+lybWAKSiqP1XTJNRaQoyEV0qG0cJUnJn2V4JhQ
RlyXLQlAO5SjEktqW4cpeCyqyW+1uDM/2uFFuXgIanqUdNAN6apkv6XO1qbTZ6+Bj/hEPtxVkk29
RHSKFWylzMmhw5G1Xl6zzbPhBle5+fUUn8CO/PDzbxQtA4Hm3JrOVZjKM2WyVYD86MbR5r0+e4F2
Mrt0fqtuNi40FyQDqukYR2d4KArbBk/u1BeGdmNCQoixDiPe2CxoeUUH8Ks00CSQ/OevcDelzF1P
xlYt0/83we7GSUS+5wT6DqGKNWNBVYK5VXNtnmwvy6B6eKyEvbMzwWEArRX5huSkfGuR5a5vWzV3
CQAJjZ71H7GY+0B3eGaNVNUWofn51rl9ZvFOlTzsVmTWxWAQMWa0BOXssgXhwO6eIrgrQ5DsUZc2
U3Bde2yxxGYrcsFdCtFcj4nDUAiytmnJK+ZGzE3+CxcBJl1+xiDimqRnNxXj1Flyf3sr/t/9WSpy
XOU1HYuFADQMkx+dsI+ZFzxjfDwIYCxyIPqr91H3Ry/yqPKibn09whX0JB0+JvrcCm6PfSwC2BqX
uLGBB2cBa5mi/eyf26ye1SlJ38Eh7v4CDgzUsZszUhOPkJcZ/tI15MGl/5T+/VMe+bnwALNeL8Cf
64AZ/I4v/sGq6qS3iaT/t/6rPXlhUlsCTETbQiz1uBU38wNdVFJeIqOpFTFqx/rgfYekMFXwGPpq
ryl+vrktZGBsVqSQZNl99nnJ9MNM0pD46oMuUOfsGvrBxR+HiK39bLmMSeeK+uOEme3h4rSReSUh
dUPMNIAcU+7HkmQOrw8PRVsEQdWbPkCfCECTFB1m9T9YDxtLVlIMsONwD9oSZTOyCXRWsu9KCFYY
mtxtysdiAjna6aeI/DGPd1eRqVwMCO2FJIwYFvlovMNs8drHBhbLCTarzd9v9/AxxrGOmsC89QFA
qQ/+D2uf6UFgAwsTz7zYR/7YmDUQsQntiGVSoMohNgYMOl4DKEcU8PZFsBVPoPaT0iVPAOh70PGC
YYVCiEjo9pAegqSMYXSUU/yK9jb34abpqPM3GqVgCEEO3hVKZRtAMl39c4FHPOt5VHyPxmaQvKpG
l9GBiwiDl4E2ZEOOx1EnAIplCSGSzBJ8c5Xv85nSHJ0CbpGCgOQvNur+iZU1VIT7VfFihVxwJCeQ
QhhVbqYZy+ysqa5F8FiffTHqhGU/kohtq3q8CpazVt+0x+IPn0u55xJOtxnCdgdIqn0EjXlIDsZK
lyewV8JGA2R7y7JGG7DkqA07KKJrxFP6ZdjyG4W0DMCfFCd3Bm/E80AUOH3efjjPQguGIHPnGy3K
Wx7E1v4mcxjiTDDnwMjcfjzi3Bq/5acWDAseR1j2WrhVFRcMnVpdXoJ4lUgkvobarfZlumyb8cA7
BmAU+O2M+UGVALPxDAktNNOgt4MC4TD6fdL5V9eeRg81qwci6vWdXKHBBInXEYbyRexfqFczKZEC
4TnfTsA8LwsSEdwvkaL1kEpvt+H/hZMeOW8+RcV8u1eJEqZE6K2ISoLmpX10pweDbQ+7CloY+IYj
sitRdD5hV7moH9YU9EqxpJShdRsoz9GNf03KH8mXSHwGN2csZVKvSvQZnq5/Wilo5xZojCd6ZxA4
A+rQ8PKwAZdGTrdT9JqbE03hHXEBWIRkmWjkHr+wP/Gb01zmVjDBu+2Z4jhYvmdHz6sXOHjq1mbl
mOyxDk5L+Ca6kttyAuKHAdjqKmTPxH++2/E56vb90F1cHwJxkqjRtJV+CTIbQxBz1z70MIw/XhS9
+DVtFVAW3PSz1HzMTuogzBr6Tt0N8Chr4fjiz2p5S35zsRHjPXpuKCN88+aMNdgRQvDRI3x07uNt
ABV/T35keNc9wYeqMd8HvT06hAhiLo4YkggLoputF0RniIzyN0TUskR33Jpb1vvqujgy5pYfsGGq
88ZWH2c8s7ssXjFb9rZCs1dYhZUgUMnTW7vD0skhH6ybRlxgulb99zyby00taXXgswzf+p4IaXL0
UQprXjDeXaXMqRDKCZhVXbNcWHdr+XPZfh/gQr14EPryFyZOUfHOZbMbtJK2HtdfxE1Y0dUj2yfg
t4s0lT/cRw/QR5KjSVxuWR0IWHV68WvEo1LRAZqc+I4W7Qz0GVLaU8IseD0h8LTCHNnztVyVH1oc
nmHcXU+M0N5uas0hc9louASm7ICBujE9Mo331aBwk1JRCMdhvP08KMVH0r9ebaeBIGjARbe2YIcB
pfqb0Vk3Swvq/3yaCGkB4fpZuBtOspnYrR9ZYp1gyoKpMUG1/KOb8K3H147cTtBOT/GMgfk4n+9o
q05XkIaBkVq+f2sQZosHQIoRu76DeWrb9UyfN+YF2j9p9AoURpf4ivinhtG1TlxFnXSw+UBVQtdO
xUrwqYPEfT7r70bARCY3vY4StltyjCYhd/9+msUnY12WZpPFiBGvtLcdUsfAAnADxExx3Dryss3V
shkoyKXIQ3uaagraRVXu09C0S51J79fSvY5VwW/6W2MFjMXrE4QD9YL2dFo5BbCYcXbXtoZj2HNG
ax6myPKQ+fb2duTxJIcDhJxAuA0iy5JpqBgiP9Ili0NmFyyBk4ME7/7o5r8o44Pd7OadsfpVGJWC
nsCOdGwktU9XtgCMupAuY8zwGYFDUdrife9UhRNGh6SRt/guHKxC0R/lWKD/SxBf04TqI7CZ7UNo
25w2Vgq1bR+AGA6T+rD1Ghtv9bvzi7YlrTv+WybOb8ggHW+H5FLygJM0b0sb6BTxlkIszL4nq7wS
pBgisacsqkpStbxVbZDXSRG9PFe8xvo03nzoZFjLuT6ZBB4sCG4waG4vb/rDuTvh8D73pKcK1fSC
SvSN1IXXWLyY4nd8CG47W6QkN7FqMfuaT/HU8r7AAGDS6GiRlfKZXUzarc8CyKh69J9oTxeQ/9YU
RGDBYg2vVYQ8KUIU826Tw5t0gdYe+j2WvYRT5AeFwwZp29VVZqhrOzttiiS480w5TD+Z8P2pM/2g
MGzg0e1kDUC9WY8ZbsgyZPniJ9TiE8CGRXkTzlZJt9OEKHBHzqIvEOHiohJvZcgp9ruIySIrS+Q/
m0sDza5JjaHY+OgjeyvhnYK5BZO322FodS9J2g+cGRoGNihfJ+NxjNPtJQKG3p+30nikzr38R4N9
tJI7Qcohh9Npc/0hF+d9O5WSwZFHiIHr0qfAm3A0VoZtArvAqimqCGKerkkuiHSV+PCfWEwOgTIn
8CQe4PYjHcfngniWirUKpTZ5SuZYtRV7d2EWUS1SdJeh46A5hWp7KNBQsgkaGLgUZTRBlP+lOyww
+ercgj44f38vFBd7U6j1l1UtCDEB0y3towE5U35uMd9EgwsYiSwHFWbVu8PhwUgpUAkZOcuoxGJL
De1ickQDVD5N4Ab4z1rmMJj1FXtAgzxAjlePSDYweSgIOaRoN19G87+3JrUk6uNyoY8l9Fs5ztlq
MUNT0Xn5ONMTzDrgFGXJxxpUwOguLoxshDwtvTv3xC+Q0fO+5AMPoJK6iwavTSB/uhGx+6FW19mP
EtMdl53kymeIr/HSfsKLDZ01imMpTPz95GF/qbD5AjnjXeh0DCTHNndWJ8LSKk7ZRDYW4TwB0g+U
fXL99ImS6lrzyl/0f/RUlM3UoJQq+ksB6DtixUaXHdOLE3VqvbQOnMVpqOYXxygo4bAUgwNY3Oxg
MfofO5qCYwq18pfzolWFSkA66z2UBTZMKlEo/eR3qrqfyEqdq5YWQzvqnhdDrt4y9OjXqmk4K0vU
h5vfCP/iutfdWnEEJvmnB1w6VOL1mKQ+TFy+8rM+RmQ180Jtf7ZyN3yeBMXFfifgJ3dskkDBqVQX
PS/FW+BR8LRqnJjK59jV2YWdXtPi/EXNnGNELgqZXN79qNx6iupezHbjBXjXTuc8Wj54mW2STXiY
bZZjEyJgmEFfe5qiIegIww74kNenvzNd+fUfEI4GOLn1P+e+blBhMXgnw/kx/9CBO996GLQVIlfm
Q21egJul8PDQHkS7RjVazjkLrc7T2Dn0OOoiYc0AKItxHROknlgg674rtYvaaT09yPgjfjWkMtXw
N8Z3J8U6inN6DBqaMRfEzQsJwJssfXG54e73fBOTD0F2Q+tsmyMZ/WV3Nt+5ZpQK2XcIXj+D/eFJ
bhKB1KXnXMUWaUd+AZcQyuY9Rp2zGqvv1Yqjh38eBG36+No317v/E4MYDOyg2frm66+BXx7/Oo2l
JyP1f2clp73CxfI6DNx3ABn7XmWrsYnAU9M9MIuIUB0MXxrnRq0f+rSHTa0s80bLlHqryATx4E9j
D7acpx4xX0ELOqATnKoN8yUgQVBPpaHRL4SUReaoZhhNNi3CR/EXQwXwFAEdhTKlnv4qCv75KqxV
R+bSEKDOmkuk1hXRJ7Bux7Ja+ougHSlG1XHHwP89hXoV0PtjbSjTByuk/WHSqKq1u8D2+aSDc4f3
k2yeTzZaHZBiLnTcwW/dtJQI3QlEfKIrdRZ9DTG1WeptnJ+CVeglHQwYWLI9nMTCqUwldzm27psJ
h9Qze/NSuDu0UwH+XIiWRgL9lb68lqKZ2VAemoiCFvmJ2TQSF8isctTEXSHnto52SJjVm00Qln1/
dRoxfff6dtl84vxLnMCVCIh9Poseqbw6k6ybgMiNkTXbkeQIlzmtdTuLvEXnzIs4JUmDXN3Eq6JH
SeqP57YmmFMZKxnoC3jMJ3ILHY9vmybcdd0FC9m1GIDfME77GLE52bfOrHtdPMP5sjXG4UqmfW6d
HEctWgRqAPvsLkRzLygAiyVJNCDYcb7jvi1XgLb24x8zAEo1QBjJ/b+MZJhv11Ck64WwKxNnEXis
TMjk9D7PQ30accZlI2X85cfVg2IFwNn7f88VOu6f+MJIqQ5Zaq8V0dTS7xyh6d2LJkmrYVTCXVUG
+pcmX0e0GakJ0q0CjubDjpEjmzBKkwSqR+iitJDYSVcs6aGrYsbwbbZuhIist4pTRMWf9hDXb3Hh
7cZwMYZKdF2qRCs7G615UzBwWPjJfmlkTqzsg30iEgzLdDIrviXZAh56tCVPvO+wApqdGwWgutul
XorWc/FLZLYZoL+333fC+WwIkn5+YrH+V8iXt3TqFckcTbngfkHBOlDYZ7Okqna7HrhtA+hnQij9
EPXGntdgIf/jsGRPkqZhbx5y4/K4bIB/rB22NoD+Ahp1Y4CIo7DC5S687nutLSAs7E0ZkA7IoBiV
4OZtmtJzxLpDPDE2+1o5MkDzknM0CTiSLuwTHgr9F+Z+sVucLeILyU3/zESSXNEz8IIaahglhb9A
Kz69EllctKLXUa8Hs80fEsH3PQ7lmJNY81f/9XAdqo3D4Q7y7xSX8BBGOnwsGQzXgEOMoZiDL1pw
CU2KN2LCToY3LbKYyqSUUW//jjjZGyWvC4la6tmEd7nxJxeX+hngrGGKATxxono7Mk+2M8TpKnpk
UsTgDi60aqw/V/w+0oXwkytBxXAaJsmM/GotedzZK8VjRHVV6vMK2D6adeVaKEyxuY6ay8/VW88e
P3YAsXZrajjgo9Pq6PY8zYkCRbiw7UEaG4DWByEj4B7Gc3uHwPHE0KXDNRya8t5HIOUU0tKi1co/
TAV19NX5OZjuMHD1D96yHL4PKO+g2PG3w8lxSa+PJgPu1JCNVthiJZCyAVKFPOxtzyfL3E/gwHv7
yEqUys9jf4+xb6rdCiOpSbl8YKX+JYKyyHU2AO4sWykMejnhcmZMuXtNwJP0frFxwE3FlfAwI7Cg
PE/U5jJleVIkoPEEYAqaj9PfRj71OmKfoWsXIMPRoTosZp2tq+r97zyy7/FfH6zljNAlzF72vL6E
WExrX/ttOs6+4vT9p7oR5C50tP5JHs0qtYSIQd8wH/FptGNR74VFTAQzHkj7eyRhlhMuFtayZhl/
enamCXsadEjdxo6oQjrrvDSxX0mWx0D4RdMWoKNrVXvd0pgi7UzddHUrV9+2eIQKL+amCTp5Wbxi
jwXiX3WgChfx82ZZknXXUPua8R3E25/RekqwxFMf+J7cb/+ZLApUlH6zasKYbbB3w9apWtekSomk
NyUjSt+YRfhuJAJefbldCFnUVRHUR0+546cGcF8+DT4JcAXs9JEhqY6BjQznDjDGELt8IR7TiriY
+bVvFeMstQuHEn9b+Erb9PM36ikaPpSj2yrRTsIjJUVkFv7nqIUtrnAgZmwh0N5+puplYEaMHqNz
EQk1ArG+xlcwbUWQnInwJmYaM6eRkIdrijERbQTga5G2scW6f7C3xbJDI8u5IqF2QJsVV9F0rf7Q
ZHtxjFQE56iiKnI1j3vGzI4X9l6EDFPIiEUOvWbDWM23zRuUK8Y0P63in3oIWMkaqDI/zMBNBkCi
WM16FOzS6sEmeBH6l0E0QysJkp5pm7TZZWaICXNcLy8hf+axaQoGEGcwKIrHAN/k1kDToVIMeb+0
xXDXQS0ybZ/Oln0ukKDVp2An6Josayw21RYTyT6F2vYzd8vlZW3Ja8uQ81/2OLN+2vv+JiJFE+y3
XkCy94YybEwRWrAXfx6/1gZp0Zc8ubzwGjGSG3SXxjNdSN6lgz5ulnZINN3bRCOp3mZ2Xwa61xvV
XZV76sxLhVyMP3Sh+LblDUPkjp4oNMZCx7hqUPUqvwkRc8qf/Fcx+Pyod5rSW75OePX9ynVTHCeq
ZJTa7htN3ZyeloeyY9HIpktW1eASlHHElY/PJNjc3qyee/Pm40Qm2WCcqdk5ybzuKCvGWpaMi+7L
Yq3wVKKTAl75IF7rzZOTXaJvXrDpdD7nTi5GeJlLNZ9v675XCTKpberha7L0YPGleal/goCdC57D
ZUofF0imM+Ddaq2U5sro6mrcqTPmlHrA/8dahtGLU/qwl6+Yrj6yYhioI5CtboQqezaz/mzRrnZ1
9um7SrlPxdXHFu8oqluAl+tX0SmGI1kUjSzJOsl+GpxxBCmJMb37LSoTGvOBrGJloD3aouH1hoKs
ZKbrV3jjuYtre7Wey9yqf7/tGVWfgEVj62Q8cMUBxxmhaQf4fY6+bbt8oYIJYQi142mzr6hOIHZC
9SC3yJfJuTboO4p7aYfhgeOaPfACMubU+oRmyo2LQ4MZpPui47z33PuPX6nQcgiJHCBKB5AzVMkI
ruyi3PlDoTSkLZoRsUJjmHXvy6A2yMihQAP70A6g61OM5gUUZvBTWSrPSu7Q5LwXhf/NWbw3cXPz
WTobCbPAW+2o9GDLunkrNnEZKhiaKUG96CC/bOOZhwq3BvrXSKu/VWxg8pCmNHQTiF6CHgPqXW04
ptTDMM/QD2zHahCs5oV0+hzDJzdVK2lI6PnPdqwYaSgTa8kUEf6g4KNM4MgIExeOtT5Sjhx/IB4R
cFInbVIcgOGAAbhoPAfapZXjx5DQGkETW8L5g3ZiDuGKHmEOufhxmCYHqix60uGm4dlLrNN6mLjT
ZKI7FOeBG6pQLG1Q80uLioVQxYgPz3YALt2+LbyQbERFA6IkDJcxzIDCLrQj25vaXX/7IWHH3TiP
x6OLZ3GNGPKT/8qJLY6HZxalZGtWZgWauAcgydImuzVpUbkrpAZrYwExx1630l9lTlT5PXhE+gS0
fLQW991rOm53UqPqGpaeD0AILoR5+90cjTDmdlwgru90UmPCp3+jvr6RJ3x0KCCGIUqSfLS0nWDU
zT2LSNyzZFqv74lUQVl2zFL6pOUMSNIMZLmp1kXGibWypq4+qi4TRD14OFG6ZYYYxnAJT1bRNUVP
9zKulXPDg+d7lHvYpryMIg57Dx5IEEmIhiFDUDDZ8ZPBDpnDocSQIDB7ZFjK9YNv8Qt7gfVkJB36
24u8n+TMzeHSR1ZlMtxW19B+2Poe/Oo+dpJBGCz+DO/QQQPN3g5tH6UMPSnafBIiYlCV9L0oLky6
49ess04FvB/2aCihyOlSCnaIz5heIl3g2Ksji5h6g+2pzv27G7KSnB7pRz2kKd/IVjQRe2uq6lXD
7gs+1mTGlv3oDB68Mx3Ym8iYLwhphk/Qu4mf7fh5U/53/Ch4BHvJ9sMiHF/7iTgeG2yi2cqj+LUz
opFWWlYXIpG/8tgbwgBeCHA+e46cUWE3AZb0HaxlDBTJ7Vk/fYdoBCirTFKB3sz9q/y0Nkw1+klY
nqBbfpRxOYSkJrvB/oHBxD3+cDoX688uaCY75XmDSLHa536xmyzvyj5JyJ8nEu/yQHHYNbV56Jx8
FBLGAfUJPQD6c04WfrfGBdRLy/2epPJR/p56WksbXA1aN45+KgT9pY44ymZC7eRifmcPX+e9P+5a
fRuQqWQ5oi3SmCR9J/Phanlb6yGpw2oiK2efTHA+eTlTLpRilK1Rm+k8zoACEukNSE52kS9XYPh0
lZh0vnbyra9qCQ29kmQk/k1av8Oaq5wG0N8ZGgKQvWReTWYt6I40EytrdrnssZebt5579i+WnBc0
916j50tS67hJS2pq0fODKQf62xdq2gPKyMNDslPH6LtqsFbGG2JRw2+RoF8Zu8oT8no+p9iotqx3
IQ8374HwKfEvNxuej2xmgaWiylkFpJ2X3ZdrntxaMJUQndSlYEZq+5/1oHxmS1fF8qsZTdYTOkRh
6ALawBw87O0oBAaQe/8NXDspVGSoEnN72LTRSoSM/H1sFROmerliF6TYP/Nu2bFEKkGf3iLY+0yA
N6+dOHwZxDWgns4HMKpq8yRQrfyU13czshAFeXPUz4vuFX9ERozCk+FQh9af5Wbhy08atRMuA1vD
EQQuzHPMRGpQaItgiUFTrfXK04uEHMbFDvlLEQSsWCxDXN303U9zjR1jyABXmNWWqac4Ry9twSbh
qPWMM5VqO8q1LqgH4HUQnJMusSdShjkrZayKgDNXGDVDIHDSUcZ4wq241yRQcnZiqzbnPXJcVrec
1eSCX5HTnMIcNwhe52MHtP8mYhs1T1IY9S5aRQrRNQ6IPRdjMjE1jhlHzY8UwYXzbT3rpBodgETb
oHoifjtlQoI3rokkOgf6jfwQHG89PCBSyB2ib7t8mxxXEzjiFKLAw9yS89KloKU/b9cTObhGVzIf
Q9PLUe5p+fFsjEdkQZmrFMtcDL4fokdJKDsSUlNzZ+E35EQNA5D1bF7aoeP95tArd1swUji5Wm4l
o/2O5MDZWWJMURA7N+cfNGNgPMmVBGkC2vC2RBmG8I2rxvnfAZFr6p5xphSFOLEegXHDfpBCkEXe
Wro1K0RwO08Uq3HVq6KX4UGOBGTR+r0uCkFmaFs0rXmX3J/KqL+MX5EbnG0dkwZADPF9CDFRoFep
Op88Ivxeho5rnKxVepY2CtVx88AdCgENSIaAQppFp5DjVsONjtywfbowuNVkM1KKYCmX6OG6yVHv
oFlwSrhtFhIj6RlqzoXPb5SSugsUvS8sa1y8Hkox+mi2d3pHFjXPslVCzGHYic8Cu6J09K/1v6W7
JmDA/uIOLmTq/e6Fg9v6gNxsYH4UKAbk0tgiNvRngyCA12enzl1hcr2rVWN35bkbY88bbD4xiBT9
hTPm9ATF6HB7eFKGqxhiQZatSfKQQTyAG+w0Oj3Wxrq+KPFe3QtFACSBfZ7jrfdv3ZGJ2r/bX/Dj
muhC40x2fqI2nfNWfbEHLGW4FGceSANCzWt3D0k5YWsfStb/TVC3mcE2v/n4iqQz0GYmmI/CsTwL
ZKIoCeafpMqDfCRLxUnoemm02JAwHmTUdKM1qmOrjTRWkA/TwAtyBMM1cZpoHg08HCok/LC10WGb
PMjqCMEz7acRfEUFjv7MzxS0dH2spbXLYHSbh0UOEXaCnF47W1gi/mbUFTdWoTSSWRU2pjCl4BjO
Hl81dOpZGPXKOTJ3VH6gr2MGxzCsQPjKOVOojzzTaPrC3PVmbU6L8z1WOCarLJnVX0nulGFDVEPh
iG+/wFmDM5BHLtRzFVcqdI/c+lN6An3H8qWc7REgfn3cODaehavfleN80CSOP+CHfk47i5pT3jrn
mDTAx8vx1mObYHk3dD35KgtjTJ+LTF/EudKFKFmbKpVOleTwo9MZawHzNSV2TjT7uIMaJU16fXML
Rb372Khgh9SvJwd0mmIVJSsuhN8XQO9V4h+/6ZUu5dTkMFdefBTIH+qHPZisDtMxZSYCgR9OBZ1u
9ne+KWeROwv0nhV/nql244SpKv6n7ELU6T/8sOQmnEXrh/oWnuaDW1vq7FHclSlLnmF8e9WqPbAM
6z29x8b5CAe+ecN054HRQMgF6OwFchqMO7H3epOAxL22jY9lim04DlOUDZO7u2Gj5zjln5kBt1zZ
UnVcqu6rfs8Gh+hcnlVuGkx7AiRnwI17VoP6eBZiZfWIEUTgoeJSGyUBs3QB7ZHfu7DqwxCS0QBh
A6efwUudEicdskvmGCJNwYpf9PMwBbksm2Q4ix13SDHWSnJG7S6v9hHQoewkhDZRGyNgABL7XQha
IRxQncywvngglTZl6n/YYN3ggit+MjAi3qUDo4HFZm1BVVNAtZH0MMYSPeVAl/oqdKTjWe04eo7y
JM8Jk1qCpi8bGONNrtcb2HvjhKjeys5hqrJrR+B5F9u76ah/iA2RTRp+WmqHI85XXtb+lrlX5gXa
O12KhKIwncfXEM72PpiUGzkP+seeIZvst+CNYSrEMEENT9wnr/sGISBol0qVaeJyW0aQqQtb1iGv
8N65X7pzNP85qoZVP2QkuWTuCQHKbpCLm1cfmCYJ86aDclVc50IBDkBcl5fisRwQhgAbLUw5O5Tw
/KeOA7rLvvIWwZpP0M2eUsSXIH55lhEAiJjxJ2tktMKk2q/JI29Feqv+ZGweDa9hydUnCTk7bKXn
g8/hUP6c9oO03ThW4ZkMU8HzGfCfQhSvp2EZNEmSogy6GrzGY5SQt0N2zZ+LSp0frtXwvj5svwKz
NiQ+RKICZ1aUnSDhXGiCVWpSFIpe5FMc8jt0KG9Uo3cq8mMHpDV7fej9cKz/iVwAvqIcCkOPaFXs
RVdEcz/gmeAIazvW1ATPHlIDF88NY0O/ZIrSaBl97NR+QoiCl/bLempopvO73tXUjys7M76VNAZu
WyDnyqW7A8wwgE7sRvDRkcHienLXroJdx/hmkADtY4ge2mPyCyWsTCQaYsOHEtfxY0pl/mpVPl8q
qolWgEDmjg/SR0C6uJ8+1/QZRxwyvAwXH6iZQtsz+VLKD8ct3pRqEuzK7s7fMKj1NIfl4xlA50MX
rNMPnN3w5g20Hjg+GN+jNWJdiLVeJAQDQmPdgRsPjSqB+REnaG06Cmk1OspRwbS5GRh8Bp3jMv6/
vrjmRCR7XFetPETzud5ue5+rpnTjdy+dijFUQ17g9QMn6To2sURUZBHf5PMQvZ6al1YXd4RwAjY5
vv4Hj+j/MJkf9wZJy8Rpihw39MS7Nr5V4AouE1Zg+c74hJHwdsbrSIxWfu7L7Xjzt+TxM+UrB5XP
9wRxwQONVsjm0G5z7DyIKp5cikxYjgzxIDkCm8rGpfubYgPMJD7ZvLoBAOnCMt7MepGPuHV7XmfO
fGmbWREfJzgFsoo8nESdYSC/kCMIs1eyFD58itD1t27P+jvEYRqn3VD0RjCbSo78qkWA5mHM8WjB
mgoKQLH/jVQmrQaQNuMrcFyHLUzXz2SlQ0MqIl0c9eUMjjr5+rd7aOsdKXWidOpnkjz1fJcDrN0y
lXbubASVgm3kmA6Xyhh7GSwumhw1hvHEgu459WL0ydxPS5MGy0juKtE65wvkUD1yEEuZyiC0Fqok
FNEjEtZ/atLK6zNq+1UwS16T26FNcHwUzzK/bIcAhuGyPKDiYPCc0DB9iog1qISItBCrKhCrVOAn
TuCUb0vRz8MvyPxx1GllP6p5nkwMer++FGwcu9AJKT93kuoD5LbFhSuIIoqNkHYrU2eeuzu4fQnr
PuJquMksoGaoGrZ9FZUIAN5N9VFGrTWHoedvI5wzSZdegmCdakfvWX/Aw2uVrQBql3DzhmQBl2tj
6leQnP01u1NGFRkvwPhyWOTRTxR+omZUC/b980Kia2rNYla2d3/7B+opvD91o2raA9FUWXPrMrr+
cv2P8udRF4kED3eeBboKhdZsLujhnfy2RZuX8bRDjcz+jMtqyD9QIITGWz0fx2dYUvXv58s5vH2q
PugeH4sHE539faWBjaAf0sep2CKZrEIAlpFD8685/VFFkigQC0nkijXnwue5W+7QWFXRAKrezaGp
3S1k8UlW82ihvbbb3oM2YuAO4tTeLoFM8LWbzk3hx2CAi34Elp+DcYy0mbbxxo171rDvrYfqYjYh
6HWPtJRlZGGbvMDtD/+xhCGaxAwnGBCj+xaxruw8jCWRxuNisL98S+96cAyfgw5OiAYKGZHVzwyD
K5gnty8pPSOta9I0Tv/B7eZVzI1Ocv5jDwjsF4227JXYo7Td7YhKmeSSJZJBALWPzNgDlaBB7/Xq
bRCRLBdFOBIltJ2qnktUyQ9sBGO35WkPwD5ZgtzB/5KIZvhIZfmFutwgt5xN8H/tB0lhwBEdde1N
ozfMKp883Z+gAtRd8HWVWpgQcci8h524MM4wQ12Sn99kXPIBWt/fg8lSMytYFC/T59Kf7ZZ0swga
kHwpKfr3FiCkNJg2ixbH2unn2cJkpzGbbI9SwrwZlgY5p0UrIIOfRe0tHBxtYG+OshTM76Xf5YGk
jYXhox4Xt22crNYH3aNeczNzmAEmvvNfLB0foLdubRXLkkoYnpUTgg65v2fyhRhDOdzApOr01QCX
ymm3Qgp9KwLI/HzMzsmzw1HgpzRchBFcxcmPCamUi2f5mupl8ubMk6AOxhVg5FM1AEV2i7KPf5T2
3CdEYarJbo+jFqPyLVurCtWEJVOg9nkdA0R6HBLwHzNDS/BWbEmG5EwZ44V28z+aoibxe/FVWU8U
Ec8G+N/QLBZsyIZFMJlLG6Q6BUpzr95gERhAAirutZEKt9lnDCAYcHJPNwcEe2QtDJfolPSF+iFw
7cz9ZjPyC0U9rRf0G+Y53KkvxP7hWOh0wEmhYXBF9wbzGmHcXO91MW9PH5cJ2OeU46fEvQhUUx+j
tzMCPXomExjhjV7wJOuFAZIFCKtQdwkBBEgM77exJD0UGbNZ/ziJWEgqv+CeKomfDIeXEhcfBoRm
bufkz1KnQfJAWVy4jYFmR8Zc0xYqdZb4QyL16ZeLZLTtT/iq89dpYuvi+Csh4ZecmjIJKAitNeTj
f3Dyqc3LWrGpWh1S8kgjbZXih6IutN2DLlK0ygWduqJ1lvV3JnXwottDBnziK9c8x1/LTxM3HlSy
o3BLkhkFi+0HWZ9f0oT+sIVDWoWN1xt5eD9zoCaMIn+j4EtJKQP6CmfWXr5VAr2hy2NuEcFXJ8El
vmSQ0tzwiNSIqfN/9GdctYA1xnDHNRQ2d2y5zfEyBC7Tim+6wHraBQCnyNHDN/XG8+8Oh5BD0Zrg
Du872gLwUrC0Qm6B48aO2/asyMD7tebmd8JhO7hvbaV7zkpXBavsE0hnBqvdhWaRv4QizLjipUv1
SYIK43bjxjCWzC0VfTuEfz8iZAJbqPUwD0pg48jnrNvfkFLAPKgV6Z7pTgfFpZbIbHxPNQLprrw+
3iC9EK04Je/u0pn32bU/CLMi+q5bJx1eLhbgeVZB0JCqoi/XZQ17NVVmPlGjOirCh3JiPlbQNQrc
1KpSj6a93AP9XPs1D3WE2gMX9kvEEn5ZV5krWXmBRDYxgHLj2+WOD/RasGfwJ4Gm+gZZKZIY1/OJ
QhHGtFpf1+g0NylMGOqWk40RvbmzjkxvFZ4QDfUh5mKLNZuwELGJSWjzY6ixteyx+MvnqgoDrPT8
UNYuu8vOk3CJJ2jNZE7Ihy+WV3CsZCVoM0FZrCl3SIWf/6800Gxbp3RMVIpdt+tgHUNqVKXukde0
LNm36x4J/jSfe3TpF7P0KCVHj/66P24up9FKJE40o3I8rQMTSPnuthIg3gCRLv+jYmwKjDtKCEnz
waJTUtC/NjGzr8VNZHBAloA4M2WvtD390Cp1M+I7WvYM5VqzYouH22mtNaoO47dS8o6PpMBP+u9X
+xzGImShC+Zz5ZHkFwN5oQUkcjA9IenoVXvDY44vmik0h/qZplBr6xvuHAJq1n8hRi3ifyEBYhY3
y+tRyUf3HNEMWXp6RXRStlDdq3sigwzxJ+hbCy+kT44eU3JK9J87rfLjFE6aclDIJCyyH4CaV3jt
wO/HaoyV0YF6eed89Cp1fP0/F4yF1ZFwm4xSiTG/jPa6Wb34LHSQOrfvZH3uXLQfpG88P6Zh37wM
4Q3pEmlQLsXgIzz2g7rLZXKpNWC2fXOmN2m5nXfqYsf7C12BQrpVCeO4ihU8QszCsUHAlxFicZtJ
6u2ECc27uuEqMGZ2TQZpD5PjBPMZTyNJeonRTevOfh5e7C88ThEV4Fpb9GRyyQ0E7hTuNY53qnVg
I8Qhyij5VtJoivpt6KHB5X3lluKRsMv58etLGFQGrOn4gZwoXTx5PTpWdka9YrNFFTvnWOBxT0m2
lmzLlwlxl7yYffnTkprfyiWKeEpyXSyTG47b+DEZWpUc9AvfIepE8fQY4pZ+Xcad0MGLiDC+UbAG
AVVn7QKSbq7OYOzNl1lhGojOWzBCVd4tN6xzB++y//z5cYpHaNFtL4uaxOpooRSxgDi0A4Y/mGDU
Wmf+lq+aisPUo6OXDCMAVr9hdjnWShNGLMa9tQ7zHGJX74xCI8RplfAhHTiyt/vW7ipffPQFX2fJ
FeY+0YPhbkJgx+HvcfCtqIwsFRRylq6Hx9oDyUmFf9q7xPgGWfMZAZd29qR5VzynpuENWOg5rIBY
1FPJxodBMBAdUzXcGiwDQRLAoMR/xaJaOEuPHZvmY4o4DDYLv6a/VC2OzlEh7eRR2tyZZaxs5VMd
gnqsKrCOFDvqCvg+zufRmr9Yno3CEpwspbWFvAj1JcWd2qsfhqyoFVxYmAkuKkvgIvUFIgT0WY3U
+9xckfB5V3rlWTivWDSX+qw7S3P16zKjPQ0QQEioNKW6ysqJvY3+DKH/3ye7unEchfAd5U09ooOG
miLUz0USA+Ax7gPiCNhhqrW5J0BNZvJ0W2xSxvOjlzf2+LVb/o+cyv9w+7baGTTQi2cZrN9i77gG
gIN7hKnwNxu4XdAYxHBZTrWDHXmo8Jy+h8jSBIGp6kVv/H5SmyaWwPqEK9gI/BbU8dBq4of0PEWZ
8pc2HmrMgrZsAHpQ1v0a98WBBDl9UWWer9mM7ZOCjMnSoYrHZPkUCofzL1FDd+DojtvW0VEiGMYr
FTz+2MDK7o9ybbVbgC/Caws2Vnmm238MnDLyCNbyy73kfjTLEb2sbAxP9DGA6gHCTUvMi3HQ36Sl
Y5l4hgFOx+LNiY/r9fY4JHfPpbLbFCaDdoaoWAloBs6aHPyzhPVonsJL+MQIc1JovVfCr+KPyvgk
6oKZN4RJWCAlSEjiwsx14ZGk9Mu60T+U5I8lewvwmXpoNg7hCuzIV0oHnDeDl7shbG1JXs3ZIY+8
sdfmd+ooKdQmPQnUuiFtgHlVEBBFiK/WNiA9J0YZpiLYpt4V40fgi9JsjC/6GamioziswT7VToCa
4ABZ6u2t3z5P/hgLpiSoXtUTNC/q2/m/AyOoPFqoiQLq2goJl9oyX/pULosPNK1/GCE+tqBMNgVW
xowy6kUl9AeAtcdW2n46c5QBC3MJfwDHHpo9H0P2eZqQmtNMxmZVvhEK2J3Bvf9irkvlPDn2xvLa
0nDagoqqE9NxoNJC1WFBneiH/keZDyIAkK30/DkM3SMg/RD01HlJVUW4Hk7VTQomdF7D4zwnMOA1
cvOEJ28BEv08iiMEs26WBNuHTpxNlh1wEXfXJ3XRbVadzcQtX4gmARZoDp2tI5oVhIMDO9zm+C35
kH495EFhpRfui/pMx6AJRGsZ341nyzbCZXP/eghvYYjyz4LClraDoSx3o4YtYNasD7geVJIWbqp6
3wOp4acucL+az0MrIa9p+krrnVxN00YIXhMzlW9eiE9flF8UTJNdMKGOBuE/vTxvuChoX3GPK03Q
xcuY2NzDu7Z5prlOOJcFWb1xa8mnxQHQ+gAhO90523OB8f2dlDsgU9auydPdVzscwdGXgHEo5MgM
yr5wJzMY4qw+XyM6KilPlix6oCgsPSm1eLbrNsV2oGjxGQzN1AFZcl1ygbU4jrz3CHGtiYn1SBVj
ZWIkQikdNRIFjALYId2I6wEqFSlz2ryRLfZIIGXFOWsDq/FKABNpd1nt0Cff+wfX7+80mFqtlYEX
u981hoqyM7Sz86P+wLFfuj4UMyiS+tPZTuHwnka6HhaJVkMUWUOdZ62w+PraItMhbq+LLEIMtGQ+
slmFAEM8SX2OPeTYb0MXGBFyCfEmCTTsy5ccZp+fRQhFMxVIWiDLmI/4LCm1uvkvRMx3oPTfj8ed
XHuS/ruFDuBr6st4RKYsdTTkYT2q/4zT+OYQEk4LiCNM37Mjhlweo/RFrz7Em0FNdQOlrvehUNuu
otfL7syQy0S1UXb7b31CqfRl4VM/Y+20far/prRNsE+Khw0f1TRRFpf6erEnVddi5ahzY2sSwvIK
GhVWRZcGkfhKD27Gqq+zyTQGmeAFyLQhLNa/HNf4EkQgpZbaCSh1jdJcNCRjgi11SpChvTglUSAt
Ud4yGf8mJEdamlokku2Zcona216mTNTjCZ5f1HSAAZCaVMw7B6H6IVejlqhKAVlVDvLjeQQegfXq
CqnHTAF3Xi+B9U7MxaUlNsCPnFHNKqiR+qD9YcdHt6DjULXW5HjaUyySgPe3LrbnHWgX67kyTlW7
1BJTPRWdaqQqvBf7ULZHVenZfI5jznrEYHO2stDqcg7EctVJHQbDG1YSb52tr4Zu96zawKXeQGbM
umjeX8KjxB1/6R5NIDQ54lLc4T2uDBikYza/aheWo74Hj7ltoQ96sXxzRJl/g5ipZF/wJJ3GZr7y
mGwANZmbf9goMAD4+VizqS3Ix1jH0AJt/pyP/4IEW2zVMdJEKun4ta8BzeYDTL8P9aqu6rcOpp/u
Jt2PZjBYJ0s7hUYFGlWhRZ7HYmd1112TNcmJzNv9yibAdny58ZT+vW/lW2Re0GnShnb/igSQsR7y
XKHbR+nJKwxED/cyYPem4YfTWZiDeSoaUSShfjAV+nIVliiKNKN4DJdJGODxlylfrkH64OTOAlSs
zXRxBzjrQTacz6JRceOGzyitLJ8ylzGU1kHUMQvWS5zKbq2k6FBZ12h3W2gQeHeNeWnfoyTtH9L9
d3qCgGMnON5zBBGO2dylCrV7TfKa0Bu4IJcI3pwWmFDLBcahaSql38G2qk4l1YMqXXoYCxz1jluR
zEVDD3kOu4QGjxA4E0xK8jI1AcwCaSeBDgj8q+exOykVtL8kVYFFCdSPEg/YDahlpUytRBC8LxUy
8h9FNEWiY5Xe6Vi2a50As10NvNKysbtPmJF2naOm/rnNZ2AnpnFOqS8CSfANIZT/Lv1eO7elajpb
9ztyUAsW5HGUWSc+Hw7EGOwuGgoaPppINc2KWz7ZhFbLchwV76KyavRqgIhFB1kUQfyN78fUf8p4
yZn7LeORJRkUHCJUb/P4S4o/CpIcq3aT/kqGscPWr8tMFdUGp2caQ+c6bF/rPcZXE06U8xuhFZxq
D2c7Uzz4UcK3TR0GeSFaSLAxQOp7np7+bPgLMg+Okq9btIVasSh7Ggeco9TXpafGjDl+fNXTAFDr
blCEOEioFbvhFqn+JfhJlzOXybwiqlP31KHN+qwCKDDh/rtCTUSt9erYdidqNkW066S1839X+1lw
Y0+umO8ikYzP6KO43YF+yE8gfoBFlyooTidynUt7WA0HfNlFALyr2NTo2ATMUNpDbjEsHekgRrom
wTfsGFZBgG+IvL3uingvWA3TsS8f8Fqps4C0/nWi18tMxj3yTDTpBROFlrgGgLr03J8wQResULSt
zkxke2zO9Gp3pZ3dpxOVuR+EfsP3v0LKWbXk2MpbWfg/fZQHVfrh2ka3u23F7qhLsDAeMiBZGk15
Bp2ML2qZ5UuPw5oimSd9l5JVktJmsifFLSJiwnpDTnwt/uIdVjT50r5rzJZPWHh4Pe7GWcXywwCK
9eO5tzTuM+dz3P6cT12BiL9yV6ARm0AB8XPHdsCNSbOxie1yq4yl9yOVnXb/UNBIu3dztn5AjExw
VlgFUGgftAWGr8yx6KAqemKB8Ela6xl1D9YNyevIRrP0pLtKJDx1pzsYtzNY0wsuadBQ0h5W37nP
ATOwhotzuh76qyAeldTnEAvWQCUUXxxjMLJPpgGxyvpA/BfD/WGaX3fsg428/jvUGR4B9sCvOF+t
oVcNjAPi6F2YCH6pR/ov6hesWfsYvyNLRShkQpsFpydHuEgV5uXmuF3jsIWMPQm1GZrNysRf9YRM
PvmoyJKlw8HFshzOTqpxPeNUybOWV1rN08QuDUEtoi9Z/KwWlXn195jKKtAwk4jJfFayAp+rxNqu
gDN152J3ZLG1Wnva+co2Zv+Ho6ngSngyATTq95mZKqc1ofMg5SaNO0o33knA4x4fdD2uM4P55fV4
jQ2byHgR4fmMwlDIHqfVffWjshWqdIYXGm9V5y2G7Sa8NQNHrj4zIeQP3u5eldThUKBlpzi3UsXM
i/B4XIBTQdBzCUNfABOCFvBw51/8JuiFvJvAUrgC2Qdnhw1IyY2fZUuTCocVeo1I7zymzEu8rH3Q
dZM5ubU2Bzz7q5z/0iFRuICwUd3YHroHeV7mW4jaY7Xuq08OsAa37e/uHlXoP5QXnqF2+m/DBGo3
Qmd1o0bFUGNX4vSc3dV2z9dkdV0esUWhsoOMm/B4ESdMM8hxxt08qjxXwJb9DSX1KHfOWKK0aies
2fQAQjA2N1ORFjAUYMKymsDdTi8bHNu3v6pEHqZA0USpAfXVewv8U2CVtOZ93cm6hFyOwxRohvKL
kAf1/ttn9i9/jQhud0YXlupfildPsW1AKYAvQvmA4RxeJWtASPpx2eHF706cp+LuE+p+bGD/YuHa
IavpNBJeVcBWcz93BqS0cF5j4/KtBe5NkSQB12WY3uanhzUZ8XoQuZaxuGV+W/Arpd+AVg5T/013
fjFiZ6mChmOQUxQt87sbTlBu815H4qNoaPKphD/TEXZrZwSETKk9CQy1Brz90uqw4CIk1qMyumuh
BsLjvEafnJJhdLcY7Wb8pj3WUEkwdAambnFp1hehBsw9pAhKjbE43x1xPFUldsG5xPtVi2VWMe62
lvGGmuxi09DFHPy5LRdyGdBRWBaQol/lmjUoLHJqhWWAMbOVf7dFQ4TlkfZeMUV7WBbMNTJjefbK
agx2GRg+kP5Ad9ooRDGuOCGRpQVHJAg80GtpAZKqxHhmRAqLiCGo0D5tG89K+XUOVaXPMCyFzms0
AAbYAkcSJDqLnXPsZMm/K3o7SEAapnuOS9OiolmbC2KbDxS/FLIjzaIO3KIlDwYT+FZTkRvaGgDA
HlCMy7+Vs4+rYpSumgtHkoEtQUvekiqFZxvSV/kC/jmMFRh+QvnzvOwLgPYLbXubJ5IaJZVA4W66
HMbRc71psQtUhtCQ0VkUNumt/tigJi69hz3dVY4S3pdQbTHiocUUOtHtDvas5DyloaA4VqdvXZKb
BgRW4Ldtudglp8gI3wbL8SqNOR8/4dMQKdgMvwmg87YPKPb/ea2GfqDdWJWLZGoOGOc4FPBQnnVU
MspZw4g02e1jZiddfJr8hGOGFEGo+fV78eRcgd4onPnLX7iewPDQmDYw4T33CnuhoScxNq4YsQcV
nZxuq6A6ICuYC7vRZNwBv9Gk9+qbqIAiWvsV0nWo4lNsN4pjpbtkv0D+ovKv5LQA7btYSmw/BtJ5
JvdFOmd1n6wjoXBrQLpve5W2qa4ZGdMmFAI8JeBepuvShow8AyE9OBhpYX8HIe1cnA6BsPNiAHNw
Dl7TC0Uvicwb/6yFFVtqU1m31R8dqbedbD73F7t1pOEiOaUqbo1/7Es/oeBYorlVWaDhH6xgGav+
WDRucBRe7ywGQ9TmMlgzQVlfZclTsiqYgBM1PJ8zLqdE2DgA6CfPzqVbQEGl1LpUrDOn7uIO+GjK
n3gjxKZhGAjTlnFl/T++0ayG+hooprFCZYuR5uep1aYuui94GOmNwLuyhOEOKelp2FqTtg27X/bF
6GhlNzRWn/5Chck1I7g7WcrRkTchtpwyNqn7Pf/L9MBUJ4KDGgM0QwYfUeZS09WRlKbY9KPD618i
zoE7hLjTdgNdOiX8KCbRrakceYdNWJtgepCd0XaaKVmJGEdpYP0Hvp6yz2vmWb/CikTsT/ugyksP
5dnXnkZoFFDXU2YhR2QnwWWlkFEc8LnrXXHLcc1JesBZzji/lgm7OnXm4pINYfq/ZLBDK1Fb1lEj
ZqMWHUOk/xAQc0OEeHtbyrXt9VI2n4DI4MPXMtQN9etNVJ5GLxpzUORHDl6npHxRzt+e5jDLJif6
hFsoFgOYNtQdV0HALVOkPbQSFxmpUd6Ufo1NrMbkIbFpZ+k9ssoDf/iBmjHsfmIhB4AiQu+Pvedf
2StSiELDju3pmap2iY5v0lKlH8QLlNock9RTcM0xnYHKDXgKiFcz7oxzHUOLu1Jx/9+eL1SLNued
4F3LYbaxDNJ1onRVCI8Ht/HsR2K9xxK0O0UODxKIe5BWX3qeecPlOCE1BLgBClAhH3RYOqLNs3mu
+q+3Dp+azgprr3hHDY5KNTXrCAjXRvyzcIk00cw4L4nMAlisfFNMzH7eJz12gx7+PFv/rbROpQzz
6cd4wrelJLQSMWQ81bXZm0rERfTSsUrtD9IAxjAa0dgUONRItbQNg99otwNEK4Cp+t6pokPKrZzu
SvsjdKp0XZtrSwLYymj4VzUvG2IXBzGWZ5DvnjaRPEk7vG+fdy0ORZGchjKLNYNxlA9f+l3rs/kH
B2pjXv5VaO2j70bn5y0uExtsKRLL3NoutXH6ZCc0e/yCaujx/hXwT5tAvCQyRARZHp+GZ2e9ojFK
ruenDk42PBkCXEzVHlVfPy2XpYq8vpByT/h/LmyQUyzjsrADeDtAN06SyfXPwKn+OmZRw48K1slW
vGJAwCqa+WgCTCwn4fjlPOfQl3sjIBJ86Rl+RCJHD6y3IjtZ7CRPR6sqqz2sJvmY7qsLpoIGmWla
1wmx6FO/mODHV944/jhBi8acVH+EUYxbEqtlGrOeWILwrBLGWNERUmok/i5KBensN3L0c1BTbrQc
IxXpGP8eoURKjTZWWzrRs5gPAoj/RPOptzwn4V1u7xYnmPYMDjqu5/BPVHjjfh0NVkzAPbnWqNQU
x334QRizm+cBjwQrMtn3xKu4HKIrxLVRIbmRAnRGGN75wL4USwp688dKP3J2RgwxJ4NQ6n9BhdBt
b3+JLsCuulsx7My6mpHSBDCNdE1dyZwyhi11Yv34u2s58fNUfCDRnXq1jikJTSDjRb5tTNbgeW7A
Xe4XUFhGPvCXQvpFhyYVCzi9OpOB9Qde7iY/VnFvW0It+z7HICQhd+0/Y1wYKgQYaTL1LiiqYVux
UYejM2fz+BXWrgWdOVtiGPz5GvKshmhgiqqyv7YDPEjvHZjl7CYxOr+vmbbdMo2u77Ko/VX8znwo
A6Zi6mQYT/siQP40Orf4SX+pGvw2jhVALescPMSwhwFAuizrZ6vulcc0+Y8bbgqPCSFO1PbFbB8Z
a55yFFVmuKICfOFySrq03AwWyzz1A10hKvA7WW6Y6TshRlEOFPHwa7lBXRq6mBQBZicylXiBsfiN
YMQvfM+JlZ5xVRxZV0XtattpqvJU64xp5+iRz8YfgwuT3hnfE3Z7bZH0gmg+p0gciH7mQAzRytfc
9QOgrMDBvpV4qmDQeqLsGblLi+vRoGLJO1Q5b5i19KH4fEv4lubTCSgBv6rBMRvlyUDmvw3UPGKp
rFijH43EFg8RH/PlbfYUeWnX+uLSBgLBcTecyo2sJw3obOlsxsCSLdFyPTUGUOSqrM3qF/eI00RI
u6vhtvoxYZzVSqv+gvB+C/By8RRnmjbnreCbbWrte/8R2bBayp4YsPAJpoVbLWU4CX5L7yrGkCly
THtmdRmkjE2mzOiCaH8GIeYL8ahOBctM5CKoU1SlkWXMQm0Hzl6Kif5KG0Sy2WGMFSaB0TF1ht0k
E9z+K5LM6yrCE+dgCeOlyfZamy5KOA4Mi+eBORVNO+9cQAIgAqhQGgYb35CpXJh4sSPm8dNKF0+T
OyO5RGFqEfO1kVl7yLHYGcF3sYkEqarDVivK864cZomu7WWTCcfY1b9c42+HSQ02yZA1MC6/93xu
GC8Ed+IzkcnAdRg5UDLzbzIGV70a8rII7p0bwHxBH1femncixztaAAtNSkBCQltxF+eDNxUR0I8G
+6UccNZyKwxcV42S2CDt2vKYA+wNxA3wxWvwxGrKOTkTpfZWs2HP91k1hBe77uKBAGEatIdWPDNY
Uh2VeukuSdXOJim49ZU1o9v8PJWqsMOpru1viBUBkSbUX4y+3acjNT8A8/sqCZvMqUHCGWi6Ucdj
VwqKpMplUVNV5tvvwM9j8tQizyrYeePnGFt7k83++/Maf/yx3Jgb7hLr7mu08gJe3MZHRg1HwX9Z
BZuA5w6O+uYWY/6OdPiKSg6T5HFrjn5hTnTHm0jnuSZ1Jd79ck4driKBwN/M7OslBVgDfKy1aSfh
3vCacP7hsjRqqXa1K3zOFmkt9kQAB28yYNDc4v/deK2rCLx0Bm69bw5Ran+C1129rimRhM99Q0nP
AuI16nCMT+BWzrEMDn4ldJUghBL0RIK4w/IN5Aad/C0I9hboPC5o7JmY53gpST0U5T9dBrEJ4WaA
Ie2tapbLb3bTWlYQ//23J1hvjfmk2JKIt2A0Oqbl1TnRKyfLLtaba8heKcKjBbJPM1xW4s62dq9B
xXNqywFwA7SVFyHap+YkjEJygsr4mYr5oRYdXiW8cQcXKYjZU/Lsy2737sO2lzJtXvpJaD0Dlun7
rwnirGXlqedyr87jkt0pHzkwxaQ9UmoL1P9vCDNU6no=
`pragma protect end_protected
