// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Mun45o0hHcfPACz0zJNXKcXOCzX0YwX2z/JqeWYOSBCM1gDSt8tSQzKZYTWHZ+ZX
VNdxRk5moT/VYqLgngC1QRW6sDdijDRZktuo0TpZ7S/AMz3H0xILmVd2GTYe6zaA
mTFp3XN5KHSVl/e2THp3GL0mcSQrzBSMUY4NwCsBV1Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20544)
l31lclMShvS0H8GIPp/6slEhpB85i5veCzPOaIAgLFEwkfueof0y+7zaCxG5j0H5
v3KcdjBDNe/g82fKI1cLMqFWTmxzWSncdS3K5AmLFjHChd1U6TuNbqAcTk0gUprX
QGFOwFGdy4nDiOZ72nxW8ESePrqt415Uhms7llm9ClZgXbPA6gXmhHbArW3UMO7X
z/673uQXndsFLiS2/3xZyMXMcMkcuuIVAmea+Af9pCzB3zsy10WvdGPqgvGdWQIr
XBROZcqouYRDCT7IrxXpScnoVyJUG/b7ivso6Iih7xgodge7tkRZLSkJWUmomwTu
WGDaVw93qiZs5VvA/58rBEc5CeSEZpJnOGiE3Cz7/iL26LqJ8u6SxmL/Wsm51wVp
Hzz3A8MVHVG7VShUGaXvBo6wV0aF0xiK22VrWMpmzeIJK9Je5VFm+hxM9ohvMaar
CMFn+gCyOHsvchPd1ExguFUbvvugbOtx1D/7LJMlxgKpC6pyUHy+m1AbXe2Ny9P1
9AF2T/+RVl8Nd8apRMyF5MvJ0Geh6Wc2UWmiFVYPHyALE+hH26/1g5q5p/CB6pIr
CbObusHIwh6aPNejXpvJs4C/VFoeZZwSYDFxOTD0vhS6PU5pkwgJlbgGO/pYfsQM
RzqtPGVokTBAyKOxMSkXHASmPHy5pyVkaOfmZ9ZqxCgLMhGg618WjXLLXu0Rp56N
M8dKH2q3yLdbzajwzUOXZYalh8VTtyo7GEFoDUrMDCpaPZOzFdZcHQg4xq+XCh9s
e0rEfg/ARS5Y9Z4fuLKzLyrRPndk6S1xLd5blLimzqtRdb/cdGGC2AvyyRkgFtCi
zDHJjtyJQqSIGcUimhHSCi5Iz8/Sql8uwTELUU3S8pXVKLIjtNSvJP8CtFhj6HMY
TtHd8MEoM+dsboXHriBqO3msi6kaUJB41oAROw9UADq9rYzZxMXa5754wDOgOleU
RwYaj46fF1wkMPURpKKNjf6njnIxN5+6xfze+Ep8WWqS0n8OpGKp/paK5RK/wnm5
brK6cm2MATGNvsNryBSNNTPY/pEOXLzyG3MATz3mvuptg1i8qdWLXBG2YWmypU1P
vqhvhOrWwFMzl39jb0KGspV/B5nHBJRtU4KhC1AemFlPcolq5L+TPhtk3K6dwz9n
z2iJ2wKD9YJslJyQHN40qvtKSoyI/qPyaKLrREZcob+aGOvKypwzLSHm3MWuvMeu
TrX13BkKuUL/tCAy73/d4vzGsGVX/yNW8+PCu6tSpA9oWZn31QDqj5ZUbnumgyx/
NVAByFP4hUqVSoUjklZ6Xq8E6GQeFGtP66yRmkNvSseUkk8ryW61Hj+tbZgEaTlS
wKAKYAeyusgHAXl+fMzhmLqI7p/IPffukJDPt4nZQ3Og8e7bFrCVYYRHrZv0wIRW
1ENJ21sz070E27vvdz/UEqWhu3vIDr5MUQkwA71XFTsLuG2+YgRHO5qJxNv5v5Pc
a57KX5faLk3Tg0fAkUnM7W1TM5y8ljS3tdD4rxlCLqXQyMmEIAEDpivjuDkL/zuR
lqmvNPqj/vg5go7JcU9xk9bKRleI4YAUmKpNwHyLJ9dQP54bk69yDuuYTWHrB48U
mUmlQ0LyG5T5GgirTbzqGfsN9JMEUigLCuIoV5BCBhhxh15cnwR91Y3NGgBHj0fZ
D1XIWR9/tVEiRGDteiNmSixQsCwBoPcs1CUMPqUMpAsH8CrNPaZwHX1hYwdK6Ci1
43LxhMArnk99iXqM0i41Up0IWatH2Tglzh4XNgWpKC3plBlJ8184yCu/UTFrLOLg
0CcbjMknEfH1hMyEzTo8ockOFfUhFzYiW8CJ86gVWy2wkhNiQPzSFzJJr2ISxNeG
23L4JKrOjJuJN2MVY4D6s8fFB8ukuTB4DyYm2zHZpPB6wYOoldRbG19QXGNyCJze
7RXLr9E9FjZq5YzNV0wgoG/4Pbk1Y2mZHXfFpx4tsPhsZ8IILHJs6ZQn4fzVmSpM
HRXsU5ybIpExuRrDh+qTIGEaHQ4lZIEFPrQLnwW5S0UMLZ9JNlKGnfdwSVhKqtky
bX5mOUcu44mgxIItD7/grr/QTRsWaMmyVzzFmwMBJI68CO4oVwBTnizfFiAVDroC
daVdKgbqO7SEQmpaW1Hr9gbSu4sIbgR35sxSFXPUGE1eTfCA9q6/E6gqwbXkd9c1
jYi+VJsKS8RufRU1tD9bHevvV7aS1jUi84NYdUOoiHPOZ7RuDRO5tj8tm5puuxIF
yuCpbjHut256zAhXvvQ2Zk5MZbSlpdGRdGp5tH4ad0u0h3n7IINdz6BowITQSOGf
0iCbePq60bqSg22szVzz2UckFIuEBoPUP6DF8ylw13OSqWLfdB10Jctdi7hagSVh
I9hMLkB7i76Y8esU1d+C+3MIXJ4SL4gRtehm8TpL4husNb12WNqeiYVNmJITHhsd
LrkgyUOlDdb0GkaiOuzoW9RvnahxX49qemwKVVYN8RyOMvneNToldeASvmNZyPqE
6bTdy8dadgro3UP4yQAcujJOLwzkdC475aH9eZivqsCrrMe7DDYIJ7aI8lZ/fd6Z
lSLND77r1Vb3Qs0jwXPQtTPxCycU5h5TYa8u0S+QlUFX+mrs1Ypyaxel4qhaOnPB
Y+fo5j45i1cadeJNbNtdArLMYt5K+r3AqXzbmjGvbM939tkluV17AkThnCiDGQoZ
gk6yImt8VHAgVW21Wer279pE4IbO1Ori0QXo6SGdv1u2rvlYxcbgiLBTpZlva9jt
7CF70Q0+ifd8UQnBeFUUbWANw34jBcqNn2SRTDLwtZMeF/3LfDXFJMlMOXANQwAP
TbTlwARxnqcDbZO/z6j6dlfPQUWhf1L8CgD/S0573rYsY6+Ys9Lho4gkYejEjFeW
R6vusfAUUfw3U7xYncX7dF8Rzw+nsqNwFvcQCT4DcBbmjvh+pb3/12dAwSY5mXS/
c0qPu06VQn+TiygZFVwd1fqBuYeUM2kpe8XWfMTJbGP+zwryUszWizdx2q5jqQo4
ubE8upazvDNFnIXEk8FLackfGN0IABSzx4p+G538NOdGfsdpDVckZwZHPK/BjTid
wsn5egDuPi3XRa+G0lr4OxHBeFoPTfGK0UQH/mvAQamztSDXPAzrvWM7FGkFv+WR
EMbMtNDCR/AfkCRQBT4DzDwCaKWd60VoE4u5/9qTMjXzHlaWP/n8w2dBRraBJixl
foefVf4BoPf+zVfZA1IPXDOAtYl9b/ZP6KWbvpKjL0ktnpqYs2LwqpozhltVMqkl
wRFqxU4VAhDiS1UtjJB2OZbPleu2xmGl3+lZdqzN3toeDEmVlF1yTCLZh921qc0X
49cbZUT5uAK9hix/q7mvsKKaCz1ovA9fPPz9EJYBnvp9MLOqKR8J2QEF5/Tn6jCX
V5GWti8jWHtUMNvKuFVPbMLTtV3BHWdw2SQG8pVJeyNnQezqeHLO1/rMdfiUWQD1
WGv7ZsvOAJEcv6I4fopyfMveA6+B0pByovWkBvjV369aNQaqV1D2UrAsjfISy3/D
ez8yt5INj2/OH1Wg1Y98lUF0HkbSDa1XTUw6zIzfKkWVSbmpqEuNAC1hwDHkJyJc
vx4nnhQzGWOjRKDbmAhbKRwfGerJdZeX5IOIunKPc+GF6LABTxD6y2QPs1ELRO80
0ooGE3o+NMkxSADvyGlGddKSgQoH75Z0lQNlYrPFgo/PC+TCeGuOYy4HA8Ph9hlu
9T3TXlV/Ql0dv55XaJ+dURJKupV47DcFtrXUc3fytFHVJhwn8Wef7RlP7ucxRD/q
4E/l3DqeV9RQcFqcBXzSIEFigajISrV2vpqAWAaF0/wdy98HIq+kfiXpmxV+nmfn
Hsxg2KUeD/V5rpnr7pW3aHLli+cygm+7XSfq3zh9FipsPb99tl05eiEW3MlqcRlt
qUxxkPnRJe3+z5xGb1fYqp8RTHxSv1XgVnUVusw0zolofsRouSMXYV0G0ukSl33q
jS0CRJzEo44fg+JyplGezF5Pu0+kBlHcqf188fAz+9uwQmLa5/Nrp8OicLge1ZHi
ml+vl03CgZxhJfUCjPKSCip9owjwto6FS12CaD+NPNAgA7vD/d58W60SxsFHGnkG
7aXkDfagdfeYf6mnOKBfJvuy65NMlqd05HLLhfoC4+dmBJc+Ljt+95hDIcvCGQLq
bxK912TAz/zWycfUqK+8ON+8Ci+6Z83drCflkHeYjLa/FCGgEAMSt+/we8f8MlFj
YLbK1cssFT+iHt4LGqQ14+/Vok4VoV/wfMXIEiP1cya54/0zHZjj5vImUwWQxa26
sHGyB4l5LB6P9by7rtxrWgVTqSk5ruJ/cpwiiyKReEWOowXbu9dh28f1KF8sNWSn
I68y1yrC6C17Rs+Ygqb/zbIKETR0L5Z5qgmlEn4qp1tULfd3WRZGn/idaLWEjj8x
uDQ7Bcehe0tHZciI1Be7QdsSh8NbD8pH1zVVztlv7TbObeKQJUyH9gXKIYhBGTo9
18ujHVESqFVA/snWt+UEiXZN6gl3IslDjxzmehmuu75JXrvGbdS/7Na3uSaTkeKe
S3aNdsDfUQHzww+RLY+bO57v26n4QidxA1fIHnbmmqaPlsAYtmtsa09G6e1S/RoV
3fkeBbb6u4eTSOaH2XQ8HiYtpIQ14E3CpzuvlU5bfRbn5zobLLDAL34BuF8uAbeq
13FZH73XkiAfzSTvvQmoTXIDk58mDSDlLoOfsSttwFjXeibSZNKl02x3OFZaI+pQ
FijZmbFDnOjBa9CVe8cbT+vEBP8DLta90x62KaWcezZOGICSF40QvNm37v8+3oJR
1cK2kTaa7EY/Kx4/FycBBPpx6ia1JgSsRkjR4IoEljBvNwOk9I8XisWsPLv/BriL
jcB+65q1+Ke4XVCb6EowRJSpov2jT2xI15pHMtuFr9zu5Qu4QFwFvfQASRF/NFbo
qICgG8GbGPVHcojGoQQIgxHhKkSyiW8PZkoIQGEXPCHseTPfvuiXK/+YUPzaw5yE
NJoQtK8v/0IbbgH6TvmLmNM5qX4Sr4nN86ngoEfNRGc0tDjcxYjRjemcX8OBMLFf
54rGJmmEz7OszpoU4/w9KJNhGt74U8DUt7wffnMvRyzRbUga2/nHedxPvNwbQt0a
DDyfHVzdL5wk5ycZonxNIoy3TanngDTozMafMbGS4IFekK4U5RvDKB2tnPNzQ6tK
n/Xfg2VEnvoAnoAtd1HeIY32Bmj3Rx0Tn3S/CmW1OdyTGI8ZkOL4klvRV05Dmo40
8BuKbkxllDE/cPlGJamscKwXSo6fSlv1+QpwzsOB3cncnLta/uPtERCGlIE84ahY
YK4bbyB2mS0/IKoPFSbveGAOywoiogRSBRXITxCCPseN7Va3XKIUxaAjeb1H1Rum
FSUc8EBqesPtay9TSeep2erYGJJsFAr8PicZqDABLzSnv+Yx2b809tRaRiuJLNZP
qW+QAVSRlQsDqLl7zBTfT75W4tFPwMm0QUZ3Jw4KxJQNQrubFumymbXHlR2K7m82
Pg+4vP7GN6W9f/jxIZo/YeG/ByYylEFSjbfquVkLEp0+UBTxMxi3gyrL4sIxmsrA
CAAIytNznl54woB0AWolT6GPVZ+YtoTi30qMyQuH6xJGaTHm56wNg4cQuKygTizJ
4xczYarNYqp3QaHL6SwxbXKQ0qjobs0wjPoiN2vSwLRuZh95Nw3CjheNPuBnTri5
Y33hHh0LwTjub+LBvJG7T7jUzhryaFpiqdRS4wQ6VU/AWkcdFTQovdjHurcd1xfl
1+CwXVVZxC3/JnHPTm2UTAMNXkL3epGG/u5XQnSi0a+nxfHjkSJyf2zpcCAAfLm+
pxk8YjXMFONV6Ql4kdegxEPaMzKlxoWYuZPYR4Iq1lKYLbZLDtMCW8DoUj1DsNL3
sh0rH4QRLV25OXokq227+ouLA6O4z/PkY9Yk1gGW/s99844tstu90E4zBzTZ3q7r
GjixTylMTpZeMwYoxT4aIGRAx2AWnJfl6zgTtG5F5XgPrhgs9Oy2toypPLB39TSX
5KoqFO6XcssUz2RgXMpKYMQO+PlKg9yoV6LAZ2veMK7Tl4JYNEXfD7B88nvxPuPO
lwMoTwOUU4DGZjDgH/zEfAsrY0ILvXZ7o8MrmNYPLVHNTknzK0holsLU/0Xh5dDP
fDs34z0yRKDKlVGinBQ5jJUfu/0TUmTS5t8/ksgjaEsVkJzFowvR4gaLyHzaibKY
Q9OVbXm1mln3bcwvFbWAV3efsbXEeANk0dE0yH4vCgvwhOc38PbZslpKMRypwy3b
LtHzCztXlrMdGjahjXW4ardaxx7Kuij64EPyPcBCqm4QByZIrplt4vIMebFgI0nK
7D+YiEaGdG1PhlLvDJMfsiyw0Z3czGe4Adj97QXCSYPZUSAHg1P17ZalnGb4PDFp
p3X4Yy5NqqYOvHRkMCWPLvpqLFRBThl0yXshIoXhQrvekrfVcMSALLaAMvEpGOP2
4qo3CZILaL//XoN59dP8GnD8hN3NBKTGuS4WUuRc16z1bLpHMkJFXd0Di4AJFFj+
Ujb+upu5gZg4vhBDgE9nxHc6eaCwuIATEcqmla+CrCwXSuCXgX49PsN7pL2p3+Sd
n0ImwaPkAQvEYaTIJqCWZJucT0BZ9oVGfmLv4jtiRjZtM61cE9CWahfWgEpKkvIh
PcN16uo6zcZzogLwFJKglIFa56q2LinBBiFjdQ+YpncdWOV+Waazfs8C2oUggJiI
7WB+bTeiPcxRNipNi4xVGgmrswdwzK5LFuga6P2awdfylvcnkchA0NiPoQ42fRF3
I8CkKFQH8mylgmZQeNnsTFMNMDnBZiPQs69yOensoHCVBx1wtaxRx7frnOe2zPAj
k1I0YY3/AusZvQ9uGk9QVj/DjseEVRCPyIjAmRwRR6jG7LW8fLFdUOJykb2GJOjO
62+qq0aJaHP15Za2jZGhNyoQOi0090/gVKY1jI7hjDsS9E+m6Nflaxa9IklWOS9H
cpNjYcHHZCp0rB+/r76byee8aKNNZx/jKnAMgTxCyiZ5o87oLRllrJ3V7ddAlvac
KMFob4nVhDPr7mF53QKHhI08edmVovE7sVO6W4KHsvrKW4cQsckOTQCX47Ft72/m
EToFIjLGB+ATQamndT5IBTmY4Il8S5GNKoFE1EnYAMZs8Azas0YqD53YdaJxEUb9
D6fmEav+c1ryA3T1n8AdZcHOeiLVruIesTwqsqpYUnQ5ATSGvavlC3Y9wgTi/khB
TmfNlWxS7MPzqqVYYdrKbeAGvj86yafYC3sKZQNpaFl0vqsQMFYzGs9ywa8JxCnC
yDlgqTh10FjHFHUW5+dcpNQIwWIt8ZHfTX2Uinqld2IP6SDDmZNAHaKAI6s2hZ58
1z5JEWF9EjoXmmjo7tT49MC2motgu8sam7UhgCmxHkmhZnKvkKVeRahHwAtmwm4+
O0wIt0DWowHxnu/AQEy7h2SXpnT+qRAp1uBBwGrM+sp+WLWH9psOubV3J786VSF1
mHo6yiGCCkgqpAiJ99G/MrL9O1OKPHjxapJwa0UzH+BpSC0w3QaxTu5MDzpBaUz9
1dt+/24cHA9lS3LoyPUWDuVcZ7PF/kVOHrsCuJVX9+DZoWynZ9WcC26CKuan9vUF
I41Vt9DU6yFaJ5R2CiqU1mbwWg6eo0bSfHQ7cprBoiSr3dsRertJhchlD8QxyBIa
6wBQLJu0tnmhsxk/8uaN8MCWjtNm9q9ygRy2YhyoCnwy/7KncLWJ97QexAjQlMA7
lIjAk8og7+Y9Ipoh3VePT/seEfUGtpk9VjPLOO2TVvlZUAdv4vMdikrbph9St7HM
laNWd4E/J+FhChX3xOt6+6FCAleWiNyBhQCZBeac4DxGxTSMYxjeIAJFf4qN/fp/
ZAB/Hf+ZXVojmYTlxI36rY73zp2MVIP3J2OJrvbt3N8QrVxpP2rbAwAlSvzD9YbT
xQjFG/8u02rop716pVstq9aOWIgXYm17cQXZDiPbuowjcTXVDD+ORExkozWI10Am
fC+M6WU8EJ4MdxNbfCsCtT9C8rrzQFewTtrlyppUWqriB3H2/gHIVEwbSzShqQIs
cRwzxRqIN3aqUBCHQM5NQqV+39PsiLLaozHOLaBHxgnHk+oaCMRx2EZtlMvBrh8q
Gz70HWotcqoxdnW5XuhLt6scQyqIZV6QePmoeh5Qz1YM+1NW4wdeRvJ2SsH9kNT+
NVPFhz+w1uZO139/VJWCDJhI64dL8mrAxwDB5zB/inaAlACdgUjDZYENJBFYt/y4
VR2nNJWUP9ioyyF4ve0bSAfTi7n1jWN8ylP+0WwQzgj9NShI4HlUfA0QMzec+MtY
yipWTenubyhXF6D4q6Ug5oxYWcutYMwWX95WwgEGaPopTZXEgAhGgD4ct6e726lN
iNNQYDYweYVhI2eCNE7/GF7lGAX/a416yicyo11ctg3V0fUSLCzkfZ19yLwTS6WX
++ZgmXIrxg0bCIl8nlR40AB8fhCASjP0PoZW6DXgUYNsFV8TkG3/iZIDJoAUF3zk
r7gFIL2nlicLZaCRu2yecatics06ZdxMfT3wM5q+lXjWQqCgn5cFWd7/lZDmztJF
LB9L58nXavXp4yh/mGxtxAvoqh5jTg3dBh9O7gPUidyE32vLHluMWCEXOCPAw4iN
cNK8RyRe7jcymtV49eaK6ENnrPKeLXcbS4FTxNdtufqwlV4/juFeL349KJYPL8I8
1rIJKf8GTF+2YyI0ql2TUtuV0C0TAoflZgz8M7+20Kizm0emvM4m5n4WfZRSiBp4
85Fqt7MjKs9KDH2DFkDuxYK5Ra6aMgwNH7HPO9GJpnuVG4FimgJNEaINfLb8LHdZ
fJtp7qi10TWnhe+5JsoRyTipK0VztKcbTSZNUzxv+LA1YaqI/qd+nsIK6yEblaO+
7mrMssI1W48UyP2nhB0dkMKrpykKLIz5QZXNoUNG0Sc9LLpUbVgw/lqB7yawplOw
fxpcuQaSQr7y/n1lvE+mwAd2XoiBFORKmw6DzeaFAIT9+vk6hHQubzugRnVZp7cH
Mhhl9IN2gwKAB9O7AxeB3Y0Z9g5JItm99NGxRHLjcN2iq42fraVkdiUThYn9s+HE
7l63QoahErkOPsPh+cgwTyBnX21RT7QKXshwTqpEBlNhsh95WLGJuCN2p5AWja79
aRfOWeGdA6VaovQE2BV7q1vAaXgVvQsRoaOtb7/G0opw7RgV6BY8XTA1N1IyEcyj
mElvSS580hy7DeW2EY5ku+kzp8k0OkmZR+P17jK5b6H6iOrCibKj8nFfPb1tkcoA
PiH/2a2twS9e4JbvjCY5Ean53/E4bUa7bxJw2/FSPOY0wRK44hIbTQK9W0RRKWeH
MbajIwuDZ4Pxd4Dl2usr+pukxFFSJ8g8NKIRUTqQfxrIDjRkt9ZOz+3Xyieu9x1/
GDzInKAni+rRthoyouqjvLXMLRc1iQN36OQG8ocYOu1suHA3tOPgjjdzA2HIF+wC
OqUjx9CvRfCo5Ty+UCvTa3bOSWlPlfOiVJDnNk70naGTGwyXIEQH/NhAyaMeqgz3
E6nbgZoKEolt7USjhSttA29M9mHBqpa76pI0RX/+k0daZkMXccXx6QLWPH7mUC67
Yu95o9jxe+bwBs8wZ/90Rr3U47n/apfsG0b2J1/Sn8Q3UXpBubv4MCx9vqwOqnHk
rmUlHM5+1o0ZoNqOS+xw3aPs+OuUdpJjT/FmcgMohfCI1f3zL19hY9SgPO1Hrkcc
V5xcsgSfyVWXwXDfPO1GencFuJl0Zq1v6pbUV889ZQztz2c9mBrT6Ub7qlnOKIZt
3qs0zWWGEgv+zFTSZs5VWfxPf527wCGo8NY16XpttlzhJD5jHWV/QsaaL5G8jd6F
X2QFc+bGmN73+93uW6gX4YvkYpV1ulhe3820UOF0wCP0SVD+MDQuhdH7ETjLvfEj
KihAh8+1v4zS6KvF0PdpVmnDTOMz6T3jkDr0sCBfLpvZCJ0mAmaqSogvxWQ2UfP2
LXsadKiPkt03z/5fsNLarDxRjhvJKxiro2BS8fc+IM2lUQeZRjalo4jdri18L2G3
WYYAaxJSZOMNcQPihKIITnXmXWxFaDhbWx2sblgDnvijpxXUuTpvruL8WmNScA1v
wEJno5N54wRpLGOzZzbTkn/pnM5yj17x68C3trWkQkP51xCLOQY2pra1b4Vjyd6F
KwyRfKqTIBkDuejOIgjna8uAReckDTqzBTaqh+erQrWJiaM9yuBhDUdDlOSynuCG
MOlH4uH+1hyTaWAKgv1k4wzwrOUceMOD+f7+iMOmFQX9xlFDvLnLPj2Qn2ogkymW
jOvl27GbApmPfEZxwAlFOEeTZT29a3rFox7bTYghtkfg9lErZ152M4AkE2Qqqajo
IG2j0MCJobWk0lD5Ht8X4I7i+KVDe+wPBY1V9cYsqMANrfoeVa2vJzm0thJ1G6nY
wWZ7cjoEMlU09iJmDDWnhDQjj6NxstW1yK3ObmoFugmFhCD0OAjBC2d6wBGGqsQN
sWbgaHeIe9XoRw3X9sezqNwCnHE9vadlHvrXGDoC+IcY302ZY6GusQiAqjt0lZ4l
fF63sFPxIop4cmpph86FP1H5tawzn+0FcqFm55zbxqxIgqjztRVr8HHLosp9BV+X
LuQdkMXfSHEq4SXT3z3tYbYk1Jl/sBbz663qE0dAN34/UTQCBVOH1Te2Iv/L25du
q1diyalpEplbqYt/3F+UINuS6XaIKX19afcmwC10GE+feSlgWOODT7E7Tbn7w+3T
yz6X4ilxx+kCI/cj3D/3I1/6RvkAG0EN3vMHoUfXGwurRwqFlWe7DCfjfxFyILJx
Up1Rfyd+XUoBb8ZgY5yq/PuDzOYvBkKgwM/F88SXgNxhWLGMs1YFgL5S2e7hy/gN
E5Sic3LC8F/q03qUglUNb5ev3VMOY9pAFQRtqjTSolhsYJjzbjH3ZAPS5jDVjMgY
FvZHJM/e2Y07+kM98pf3SA4cQWbVlPW3p+Y0fXnk3X/L50YvfgazdYXYw0piBdPo
jyp725ZKIH8lO9du250b9LnEeIUt07U8hQs48MDWyEgup6avKXUDWuEDq+MMtvHu
BEpjrjZ9SHN9wx3ygTzPdDTNOcKzswrwL4ZisV6l8XT7fFpac3/ycbBQImz8Ts3A
gLzZSv0fT7t1VIokt8VwTH83zyMTlXCjZrxicXxDTBpLuZywdrv7nLtuOXjd5Lq8
QJSsWEjDPHEhL6310ljVscJzfAIt3DxgkmsYZM7utLXjk4W0ZzT+WLfADRdhpcY2
RWr7SWizL+sq5lMcBkn5QTAdD6OqW+5EB6l5AjGPsAib3/iadjh3S8EJZROdpTMA
tVNx00MywZsxUdCegamI9vddd/GxLRmx2NQ5l6N4xagOfss0zGmdMYbu/QyIft4A
r6nQwiPUuxzRfRAsXe/m/1NC47DBpxhIixSRgWlRdHdTEV92cSnCGj/uV0bML7zJ
H74XBjwbbHl5pCttH8x7m1XrSqRtxOAwKhiebWzCzP9nJ4wvq9RdoenoeRbuzBLq
/IoM768RJ03Rg4gdF//8sW8tRO78J28T4DoupqQMOCuV6IEABY3DcJuQ3aSTvtXk
wRkdsv84+MpPDIzwXU+6QBx+7Iqydmu4QdbRLz4ueL/RI6z/lrMILVsCNELeiYPY
R0nfv0wgUzXfxXV6mvtocaExnilcYBzxGyvnkfwhjmLsDbhQ1AU51qFaKhSdTjUz
CzTes6ntmlkSPCn0Y9Wu89ZKVbuogYggOJdkUiTvi+SlV3ePWmHRuDEA6/gahcY6
3Gsun+iPFC0bdzNImtvga/MUSQ+sOlT/UNplAN+kxW2tKpam6nZMXWA9ZIMVFYjS
tKwQ/ia8l0i8VIrIz9QQcqP595Dfvjnp7vmHhM1ofTONn7SDtmVbpeyoJ9d++5Mn
nciO2Cx6PKdO4U1iZrJ9HbPoJK+tqSBci0pby2Ur56r0yvTDzvc8/6ycCpnkDlY8
k6+rvoBa02bYwwHMZrETldrVbCcnAvT9opa1hZkJfCkyvL60FziTDMeODhlC7dK6
tW7MNa50u5PDtPqmHx7UgvlhTMbJtz1rZgO4znj1q5vGXqZt6hRi9JoQWe88todp
Yagoaex83a/QGTY5s+xCMNvygYz00x3+0YoY2SuJJIIaV58SwuXubfzBu7ZzWBeC
B9Afuv8UydYRqVw7IlOFZw3gXmpKaTYt2FHz3AtVVK7N0bPxHcHW0OHS2sz1tqTV
zXdjkQZTKapodoXZUL/gIQskkzwsQ6/9R/p60I+HhRjvdzkwWgfmfg6a3jX53zUo
FruM95brA0E5jQItDrbpwMIgwwdAHIrKPcv5P/IDWKf6kacpLOym+qF76k1i7KOm
duF7Hpj7X2gPV98lk2wlb1MPOCBsZqXWixxgz7pqCv9E+4uDkCsyr5HkAfx7L7wk
VOJGCGxZBD2cpFxl2XV6zVqyVdgVsJDAQelq+YSUiQqwzQ1fGiJU8FDtveJI2O9W
Q0KqAzZ7mbGsficOhfOiLff25PmwEpGqFFrxuKkheC1tXtws7fDI88W0es7o46AY
vKgwqUguVuGxecGINFGgSzGQ+4zE6hDBQTNdCYRvLTLgty6OkLJPo8pz9Ee4UfvY
NpqxcPRix7Eyyay5QwQBKJ+yJV6X8pFFW5deAxHlCZ2FD+ml5IPnn+yJVgm137vt
4zQHiTBnMKMq5WM2vcErXZ3jvRZkEZFjL3EfyilO+Tp0GozCUrf4ffQuDMKEFdwk
8LvZjW50rl+x6L7P4M6D5kAQXphBJV/7ONvWEuwkWvX4kT7aZmnNnQATC9JS9NrN
rKFhGfmOjfBBJInVaxNNp15iEnlxNvyTGInFPe7tiEdkK96whXK2Mk3Kp2PtepwZ
l4KEQQmeICrJ4k4lnUHCR/94CYKSbiT4VLrXZRAMIJwcolq/LIDkvM+inSmBG/Su
6wqUqyM5U2pi1oTqP2BbkUin13bGJxrAorsa6tsinolCd+EOyEi2SEo+JUGKEfJY
eIz1t8dbEzJcre+6MhxLueVbVpNpzYp/UXwsF1QGSR8NClzgETdj7fM40MMzc4N7
o0R20MygGHe+aHiqJ6l7G2BhBbVBkCz+WuWEBUFW6eRc0PllIx0X8obM/N/GVvIl
ayTWFyPbVe3/kO6ExwxhFqxwlR2lUJBiWO6Cv/fHXPLypqo5g9nhQhUrF2nVh90T
62pWBj1WnXuFMvCWxbuH+ff2LBA3Nx7IoAT9HzHvN8tMeSxbLL+1LP7ZtggpGqH4
+eVXsWWwO1BnMjN/3BTwr39NDCNjKIRP+B7gyBBG3kcPb0SreaBCab8GNowl/fp8
dG0381NkNcKL+fhy1+5bnY/neChV91VVD/kGUuxzo+xcXcNpzE4+EuOrYPnmp6lf
eA3VK503nTvWFxmo9Tl+wKBecrCeUPWwI+zfrGHCpJkdznpUxV504VLlccbmMqAi
mSShOrt5oaqM4x+f4LOVoKUKrDbR035Tpho8xfPTJU8LxTCWcDLsUvbMHs8GtTxI
iJ/1A4EvYKCeHh2Na0R3Ioy5KOn3g2xvBp/3fgIajf6Ztfh0Fm/IEDw9T8nIRFtV
UFbPFGahYuALz05O7woWlNxYHIOroyKDFBz5cNGqL9Z64Q9Xpe2usLT7Bm2jHfX6
I2Tmx3Rj6ESgqhKkXdoFIrBLQ7uS6UenCIbD1YwVarNQqgCycBYQD0leBk3lZups
83YIDDNdkT7JHaQTw7FMXIA9wPbFNMLVowmBUIMtN6LC/jmjqr5bexOkqaC27CO4
jIpSAcsAduNx9IjkAHOAPpdyFzyfwzGtcxf1lXSaCZ0UvO9wqpMZb0JsVSTojXEt
yYTSBEoeSgYWRoj2nQfAeanCeUCsUY4Hj6PqhfaZ7ABADCwQVwobRzAiAOW2SDUf
gW4tbp5CEUBy3mdRUtB/USsoZrvDemZdeEwM6Rp/4u1unmzYfL5yEN2HUT/AtoMj
wEvRvYTIHRIv12b2T2F3pvDMRNHRJ/LGJilenRlkRTa2WHwIz1G96iY55WyqEyNK
XPRoAHqLO3/RnJR3SkqpR2neRhoOg1X8IqiIMYHo6YNYrq4Its8vj/CVV1Zah3IZ
/1LSyYPdQnyruOTbWt+ktovEfcy3E2RdxDtA2oj1qKyXSCYIQNPa2hEt3MiPpD4z
lgr4Zhl7FKAvcpBZatOrnak/sgsPU+jJrM99RQ1aaF4BuiK9fVA2liu16/h8YRrI
fHC38ItbsanBZe8gbyrUXlPM+sgOGj7JhyCb2K9UoDYHMgpo4fVfGaBrgZI0EaLe
Zsuvom3ylONz3ce6nmEfkmf44dJh0tPGfEUvifZ3x6CxsSX1Amc4DscKLS9d+yKK
Fiz0OZXOvRWvZnHyyplpNKRT/c/iiTy915IpXC9bVrOVII7Qn9uuoFQVpbp9qfZs
GhLnrVp5czzEjNRIQIgxVsip5iV+pZQ0mdZN7/SBoikTiJcjYkpVSr4RY6o2yEXP
dQqF6837HxxiC1/0e3h5EvbrB+0zLUiU5dUfqJn9DE7gXKJTbA31QCclZA+1Fqyt
V00D3As89ABhFMqbI+xJJOd0a39uq/TjyUlssh5Sa/lN5joVP+j87xBYEAQZdeJW
sPw8L+H62BbhHUQi3tlT86veilzP8MbMhH8KP5Qab81IZTa52BRoMto0sMsoo5wW
a6hICvF4bfkFXVz2d4w15ZXbLsKxIN/R4qnu+VW0nBmUVHU8ag8EZbf+508y5up7
PjSAvWeTfO/808wFLchsD3t7GVEB0fH3lDb1G1ydlb1d6JC4Sr+Wqk0WZsOYo7Mj
kld+Cugj2SRrOU7qYbn4PTUpd8syoL8kRnPgW2zS2koFs56Rvr6xfv7X8TS1l5IV
ftKmB+2qVwXNGidDZQCGeDO9QjNqRVjdRYZhRjgdGtXs3nXMYJm/nwo6dJAOWl96
eRckr4zDZZctBcc5808/GuH2ZAzNXF/JLFjGM5sjTL1xq8RFtYMqN9QJ2D6bKL8k
fnz77Kfc6HCc5DyonH9yj380B/c68mrD0x/jn+AAiduq9t+z/hmLiYbCwADelyge
U+mVVfpHMlaJxHpSlhkGMVowyABHrl8xvLENvJ9gMpXR+qPsVvyl18n/zPcadcOh
c0FvWJw8dEn+n4PWoybw8KFOPMuRb+Wn83FjD16t6CGi/ko3Od+uoSSNj0vS7PnH
6E7FL/YD0gN3f8uD5/lsyCyZCd81pVzr0lC0TfJ/ugbP0eMtETg8PWCqTvbxEUgD
V8cWlNpSgJuKfXcOeRwR1NuWTEUUwHEaSTK3rQNb/UNrBahjI4FheICyMSi+5OPX
2LilAZ3D3E+o1DtB0DnZaTSr5+MhSbU+0KQD6vJA+lJ5PQ3sQLB6ETzHieCil73M
rHIyfmtb/p0da1TvDimDg5qr55psfmQcpQirt95Vn+QXNfivQaNaLxCOiPFElOmF
DIquOEeKfskeHopnxDm2vH3oErUd5biIZM4KAAIGNyOtRlv7Mgl4Bkz2fE4kTJz6
7tj2JzKM3RazkR1iD+YvXM8jxxL+g8oiac2DbWm8y4pizfWhxST+kxs8RrEGCMGK
3IDTWe6lBSsnwNQqNNHSNB7t1V2ffEr/g3qUMD4pVeCPD0/Q+8aZvM8iLZ99olhj
zBlsfcpVfU/29b/iwIqpzKDoBSDCPmiOJHk0nQjEPwbqe+0+/1vo6GaQInCxiTQs
jKydxa2m917n/LY6y0M92ZdzQPLpRdc8diKP5CYymD4DnwNkcJy7MEOZHfUdyaEz
VNOxXjTD4lXz8VJv6rNTjNTKvXSt4Rxnm3+IVKmpCWo+ZauN2F9x/TS1F7AzqkcQ
jHZAsdAjunywNa4y2ZgLq3MUj8Xja0lihk6ZHyWmwbhggFSRyMSef62yuEAB7Qkd
XsUBNd+pYRtV+Gl1N6PHOY126HX+Vn+fFSlDZvJbhsnvq4A2/3RKNZS/JIRRbJs7
dmAxLq/ncl89iNCGLSMObKyYrNNKRp79u62VX6PrUmEXCjY+QDNOR0UfFNNqtc/z
ke2w3WtH3MYelolkR45VJ7eWLmoubKqIemUAPYdh17ZRTujaFm0xJ4eJ1jinpZ8x
gKI1cs/EgNbWdXD6ISxlLa6Cv1acg324uFDx/YCSiwfvVMvFhDUjzI7vr1k4J4Ll
quG6bs5ySaM22YtUIsar1dXcxFQsmBnXPPT4LRGq/2P4iSGNworl+/skS9PHVp/r
nUPr374PhoGogECJsMBKLpRpFC/Bry9cpPKFzxfsF62sLa4BELUB+4RzGigSn21+
FjhkPLX/bzP99NPf5pUYZhf0KgZGeww76dV/FqbmHAeg2VJLpO9DwNXpzRAXTc31
YtdyE9Vy1+tvENVbQ+sEdEVFMwpuOGfVCVth1lGTDLv1gcUZeALxoKkRwNML3dZO
Srx4UjpbUlUrgveCYyg85Dphy35aoLZQKJRWiMg33VLQOvLweKKb+TNVmYjpSg6V
k86J2fdI6xb9wZ/CJbFMfZnY8vfPeKrAxqTetITA4sAUdO+ZCQyh5FwIz113tV9Q
q50AcX1UukmZHsz7jdhdK28bYVOHvQpHfAbdOhsMKSFPbfUZv1H4tOVlSp1N33fO
a7jlw6fNLy3y8nmJW+btVDBBKmsEZmAcOvb/kRKjVUzfxXE5RQsoZOsfYuMqz1Uk
mEeqiqThJxBuQiVex6VyoRTksvoViCOpeduJRYD0ncX5WmnrWdoNUwlvTmX3Z9QH
lkayUQ328MrUkU6qGAkFDogXHKVprdUqA2QOaHTON34DhfM4UdQChdbXEpgpIvhU
vEUH3cRyx+UrnEF5DBpzTuk8dJyWXYclACNAJ/+rUtv2vf0lYQd0roYDcJtCSQPt
4jBAPlS/p5A8Fxp02iKhKiPmLQNLlTHxgLHWx1Kq/JZ88k4eMax5zJfIL1gviHMx
666nzb1VjXXCul9BFa66OmDng/wnyAiU9jFFqlct5YOxQ/2lT3nNazfmEvSZsvTV
gDH29EK6uk4EQX4+vB2mM+1fO+rfBcCklA2oYcDZrBc0WOauE0ZFp+Ow9PT6R20A
ihaugC/nj1iXuIeV8cD0QWlnRvOd9vQ0Gp6res2lA2hgg/FuWy94DPapM6JNpLAH
2G8ofJu/eZCunrsBYFmFgZ1I4xK3fe/70OFdIXs+FR/3IVpxWsaRM3Voq4dNhUqU
yFTW+v77HiEqlk7jGXD4e1gYn10Xipqpcdf+eZKRgNmzGaoNO5JT/PgznXl5lF0j
smDZsGYoenaglRbE4TKkWCQxfVF7rH2NbB/LMh/H0vJgqRI0ymiX7RJ5jteXA/i9
NixErQSnCCw3BDpB6BGujaBgRXMdz3JkAn890yYa9CJT79Y4FsL6mC9agzV9fo/M
y46zaw2FqQPmHWyqrusM3vU4jTAZwn1QuqwQuL2HNCzviSKguUU97XwfQg+0hB0i
qhbuw6qBckgIsHUEYnbwp64W0Sc24aE2SI28DLNehhRcrlXhvOv3o0O+awoHyEUR
Eeg+T2RVXhaC92qMjJL7BlnfCP4Jt70VW4gA+Pv8NpmA40BuvrWgjkRgFzMIOmMI
AslKAIWF9zYX2/KJtbcYt1w71GB4Z9E2F6mOnyCyuDo7OqgYLtmPO3W60ZZ91VlE
npk1DJCtBjIJrZf2I/o1BbGbPUr8O5WmlFn8G4zfkOaXjmuKqLmKcvOWE4jqg2oN
o2o1Wuze80ONpAYv+tAaUEvIl6BgaRLVTjAb7CDNvD7jtxWro+wY0KbtNsUXf/HI
lcUBYETIiouO/Lw6j8xES7oHD/JfP/FWQaQkA8WALS9KzDTnEuydE28nT6ZmytR5
/xgKqYI1YBdQN9nK8kk4BsBllmegoj3hoRLEtYxfFX4csufiedKzHqTASAuGSP7u
3Kwz0/E+iWGmpXXqUHYZ75ZZURoS/GnmsUvYRp3QTsoCX4pUOWgtVZr/pwaX4Zl6
xycr69mGWEtKcz0HKSxZkag8pgRmS87af4LuVtoGo1lqFpCF0ScH8y3+4L36cwoA
MHlOeHdvOm/29WmyN/ThFunYI6wbvWx+pvWdMdQkiQvl8JFko5gTa0oTiO2UaHhf
geDWqlmyueEsguT8yZfFYG6jCSNFbCSHTMCHxyOq7jDZ9ZUIznxrz41Cw7jjwQRl
Z4gU96IHBZoWC97pp7OR3P18oQApyBh0mAta0GpnhlXlvrg4/2JL/X6v2w+vCRr7
oC1pE1eHIATz+J9Oa9L4DXiLWa8iTtMva3LoE/aOSnWJxK/l4CZL87aU6Z02bbXu
JheF8rOZqhtrtNwFQ7VzmNRh+U9iP9gyoMY6ZWlZs+rYSdEjSY2HIz2TMapiGF2d
2TEKGLKHyEuZ1KIOuUCr0TqfGpLLqJYHCgXTd1dWWHyiB/dOAo6UpfQoiVjIbydG
G3w34n+2W6YJttbtc/J/TeAq7OKvJGSCETUe2JgRkqABlO58DVLQLYAfBek+BMUd
Z3H1RVAlSIDDN5UtY4VW+VzuV0HFa5T9EdJCRQOh1Auk0FmBCSVZV06kUiP92GBE
zqrVsLztO5vDIeBXqZnsHBdKI83Ae9dgaxVxE7Ybj4eBMsjEOHiuyoIicpmxl0Tc
Q1HkDxOuEg0NpMwcKQDkPMxF/KCuAwskmBZ6eAEfXjbjZSLoqxA3waWU0TSLZRrE
Y+HNgs8gPbSr8F+19acqHusdPsg++pVrl56NJjKFUal7KRzf1bFN92sPAMlnHqS2
Cz0V/7x2zeyh9eKd6DPwfC6XyB/6r2cnvknB0QcnC0MBLeRF2oA45NGeb/TxDBf9
g+A9xckOUIWqy+rjYjKzsroNszO+2NwC9xRHk09B0mSKcuMIt6qtJJfDWXFIgtfD
nNuqFvo+KJLL6qi0dusOVKbuHs9Xe7L0hVlGi+vOGAsA+G5UbbPt/vkOew+f5btR
2uu3JlE3zVveWxgJvHjJvlh8L8om4aHt+D5KsZ23dxQM/ikywyimKKigFo9h9Dgh
fURrlXTCKnEKVQ8PaWY2vtoBHZXc0q5YGrj3eZHVABdL0iiLlkmK5+Um9R4lRo0m
iMIa8sQ540u9fmqqHc++FWzsy9f7H46Xoxp3WB+xb1JLjnNK5dbPnkBUqDcrxdm5
F3L8L9/2tQIiP7b5g+NJMIBpQY4Po3Cxvzm1dSxM/Gi/dHD/fIEVXqG0zpD3vHfP
Qhmqj8P90797SEPrXalQSkVn+Mpa6nTC71jmNbofkPd5q3FjiKJcmz9pC8P2KJGQ
pk5uErNvQ7VupL54pU6cSHA7qypExNmdcsbaXy3GpbG2qhQgc2iwHmgAFRqLv6Kr
snvvACffNAt5wyJvmvMmyv+t2QAnEFM1LXQv1/onodD55J64/oqHCZFevik2e689
7/9FVF5mcx/1uwgL7cvYdof8rq+mLkb8XDeKus//KCnGPUGJ/yetaZltsEi7HuKc
kEDPWeJqVBAM32t0/3jV/3uTfZNBS62fVGt5S8xOelstAy25ZbJjXPmfN2Byb6ro
gQjB7dC5y5budp50Qeg7uN4m2LAcsXR/dNLfusyWlO8rPVBNgk7RXd+LGOncMlEc
IngUFcHOO/Bp+OliN9wozZxTuWDURSXKpnvaIIeY2ZIw7nxQz3ewvV+B/9qCO5DF
ZcXefIJ37snCQCwbaMQfj8xfuazrTLexRX9y+d9jXalewvPRxL/l9OzjArgW4Jyj
Bpx+o3Ev9DHB1q3NS2Nhj6Ar5S6f4Ik+vO5DV2VoQSID681lYmv6F96aB0+eXEJK
d7rQZRB5HQD9Oc9aSfT27ge2ULSFWqI/kr5FwkNpw6iiI0zLrsVqao9rgfp2DP6P
hFp/ctpqpuNXTF46AJ29cNpVBtFJYnXg0juGjuRxog8ji+l7tHZdn6hKHzR32AFV
g13ikZ7e6WlXkRnIdqzwjXDP3GJ6idvrTaGtY90owgv/PFtYePJFlBTJydeowAJw
bwpphjISB8Fs011xdLAjZgdhaYT6d7oDwiVjpoY5n4dpE3db0hgcs8hEn7syvcSB
oooj6SDOK5B1IfoskE6RNNzyDClitqMeu3J/70lCnW6QDmfAX+sAyEKG1opx0QJZ
+oic7E06XhAjLtz2GCQnsPft7PXMxFwABQXy+OkDEjAPoLDHcvM0M9i3scOd9n/h
1tmPiIJ3Zp8cPw8R1GorJ7mWc4G//LVU+8/YA7M5orUxUYMR7b+tHOHxqWNMa/RY
HjA/rX/olEOD6EmRq/U78am2x23gzLkFhrKkk9jY35gdyplGnqxvWEVVHCvvh5NR
MSDyEpemrKsR0Q5TvMLCqMt+b0rRD1+fKPtm8aNSbPzKRFkB9tNlnENSye/Gv2ex
w8ymw8xrzO+kcXTzhXAn3iHziPkHCb9ODHJ9Hkmio8Nv3odrIecPjmmiwTEk8un0
pFNA5PjG+oqkfZwr8k1XmtavDwtQ0J8sGAr+fwzAnpXvKOKsk5ydmI36tW4iK2IK
38W3HLsUXlYjVooLXn6RqAyGZUBuTBu537B1ERzWvHBQU9/+sASZAzow8T+IPmSS
8e9c13AJqpf8MdCN3xenkDdMVnpIF7R9uo3fIZpNuK0Ik8n0I/cXsC3L3Xl2mdFS
7APjsPxAKCYIAMS8NAFDssfUj1NDGTez2pbuiceeedpk1WjdC8fo1wCyBzs8Epmh
LCwZcSpGI10uaKUWlpHCEPpaJ803hzKG3VzZLMXeexGJW+VtOw6lw2ktUE+QxtMn
WCtmkx63YXcS8s4liqOTb9z1sR4uFxx14vmc58UNbzg/R02GzYbiShStwg8OuAGq
8odadXPRbvPQFeeiEIOQJ+YK6DZUgDYC4R4kjlctehYhzkLDiRFf/ZKdEQDw1yv0
npYecAfeN/yNPpA0121hQYx6pDfNe3NRT7IzI82OXPQ8VBPs2BYR6rR33rvyODyh
reXEcqPZLGhQ8c5OiaMlLV0KBUQDd862O9ad4FtqkQeumfVfCMfhjGvq2qcDnyIC
pcSZKUzxBpyLemcKvb7BHlEG5oANVo7LZywtN8gx4EeTuIujxWbiVpVoXrV8Kf17
zobbdCBKBdSKVMjoVkt+WRdHoYmyFz4Edf3RtXX/lq6H8JBVXAtXkRtHIvEGJh6h
r2MPSWTq6J5ugMAYIVrnQELQEYyhKhKywNl6MpBgfjc80DMZrN/hfvWO21AmvlbZ
LAgF4iqyKbGzqH6qbn+nTdkFr7cNi6D4ESKORtuqDAJveWF3YTsRfRVONBlyjuaf
FvIzyXSx6+AAuAMINRzmkxqfoMhsYIdUNLNy5H4KMeWFjMqTR3OKMd7XKdulhggv
pwzcR1febYMaaBvKo2DDZ9QQXFii1icVQGkykrPCHYAvTDur6wgkMMGHOu27m+Wy
VlpHva7NcJAMwPvXwR8DmKvDj/2BuZQWG5XWqo7KDgz9sJYyrB3RLSUrvmnccjUH
YSfzh5XgHxCJglMEuIi2GEOtdvinsIgVbrRYQhdZCD8G5+wATYZoD+8R9VojVQ+v
PTPJ+TMFVHkxJZ2oSr221KOJ9lxZ4SLAGQhWR5gPj+PrUGoNyoi6v9samBLvBsee
STZISIB76svHWaBEl1dSfRX0yyac9y0rw4XKT71wje/rbtmsm/X/O4/F3zd29/6C
uGA6ouWEqqZ7JwRITSg58VRZI28FRA6yx0sqDu3C29RPqkQkUkcx7b2TIp1Be/1Q
yP3ITMgYeZw+iiiEWGFvglVzIeF0ZHPPmBpb9J69diWWpQ1WASHueqqDAAXjpKEd
6bPz5UX0vqqQqnQJfrQAlSTEbb0g+dEVqSe21+IBw0f8t6lEB4kC2iBRTGWsxCkw
DSyaDuND6nC/9QhPyzAPnGgmdew6heT8Fbp3oV++7QWZTf3w4lp4fOXnt8ZzEbbD
rO9GgnQUshFj+AQrO8VJUtOQ2bjCkdw/VnVitomdhb95JjXnaZU9KSVDT5Oijdkr
UyMovTmtzDG5N6PpGfm9AX/kGz3ni5dYFS5qIya/oS/kmGbXTfS7YULPFrktjEHh
3Gw0vRiN4rMYRPSGgG7QfG4g0nsEtsLxFKaaxtq7qaoLH67W8TyRbVbY9YqD/yYy
a5J9xuDLC60rXH7Ea/9p82HDnMgb7/D1el9cZ81tLNM3ZxgokwDG6L8K/F7C8uSd
EN5d/4SQ+KsnHmf4OvAN/GZt0AKF+ZahEhOGQjB4z/6plcRD4Zas03L4ryVRBjuX
al1L577BJQ0RsX9+vpCjrUtu+l70FXkkpNBjsd9wsnJP3a/acrRL6w77f5ca3GsL
r9g9vVtmMPgvelhMyD1goKUAIgzqPAtQPSJsav1guyioGvkP0AsOdOivJ5VcIPUa
mo6FwNdMDSuxoY8ihV6BkIKd2H9g5UOBgXgl/lJyOe8zBhJxM9acgDOe0XmNYvbJ
dIOd7ODOEYNomxXsSJ2Tp+s9U7jRpS95IBLg/E79/DwtXVxPQp23DvQvTymzN4pT
bijQS+sEz1Ah6JfzZg7GFMw3e6bGTJPJ7QwWiOwXxu0JXdwIoNum7JYbOSMKsWYz
SAkw5MfvVWHjDs0BgUbtkNjNSZ3d9j7JogM57WG3YrS8k3kJAyiuulIBblO/KeBu
rNqkXfQM4TzKktSsTrYzlJ8TtrYof9aD5Fs1LB5GwfOATKAJzsCKNsjTXVyQ09wR
rIsJXSAWkPs829r2L8LVeebpOFpIntgBWznTcnX5fOVwpcEjRGUTNnSQn1JBFHGu
itjeOmZCoX9wQ3qYHuKyRUq2LzWHy/2usuSBLyeb3DfCaqOrVBJDL0Cwmy+aTBLH
FeGoajsa0i0JILjgRgkVALCRrwMyReAHC0dusKPmPZGGjG+Xim8tdLiQIvUKizAZ
SlBu2GJEHeXcJjqcy7ueRvVq5Xh5RD/zKBqsg6h0ABMlbRWFM/0A8HmnmKfmkIWO
YEPoKdew5JUUKLYwiqcq5Yv9sz9ztzHCFV6P9CngihT2OUCPzg9ZmnrjNQ++0Ihr
0nMV2mGtW8Le1ShsCCQcqycEVocdEkPDnIBMyxxTh/10ExV/V2qvTAjB0CmbCY4A
j2h1HVYjfXJ2qJk8YuoJIcpgtRevgYxz/ZNdh8ii+T+m8CUyYA9D04zZFDhcorPC
Gn6sfv+HvuAbPIOINuJ4Vb1AI/hXzb87v5eoU0THLPpzziLWJaOmNCR2l7Cqsr8A
ynqz76BvhGgXO9OmWdOXWKYESyRNoYlL041L31sxMij+nKNhEPBqmeJOUgF3Nd0l
P2A3Oc0EdGFnJQJkHyqnYVAB3DDXnsZgwJafy8IQnC7O/mJh00FKc0zyIyjCqjsv
B3Q/4mLcDRH8f13ttCL0OuEOLGxFbB7MaZsZ1cIY07JmAgHxnFFUtl3QVhGDySCr
sCJPxcTiNXK4t0HqWN6Q/ZwqbYEoXyvKKbbcsdvbdx1V/K3z8zpyVwb+YO8D8g2X
nXH4uYBy+nLF6L1PamO58F6dtoVVwBlou8YC2+L9/PfJ10GV2Hyz3rBYxV5/dk+F
hneNzu6CUURuZ/1M7lDOYdPqV0gm5vOkARDli6WaAE/HUvoOEMX0EbE8CoaoChql
zqe5MdEy1SDFOFf5KfUGYvzRAatxY74zNwFfJvi7e/eUNTuHvuaE1VsdMcbD2HEm
Ssgo8qqexEW938LAJVyuAwt2c+TFn27ovx5Fh25lfghADBJBKBgziQsL7V2wdqq2
wOGpJdoUYhXsMFyxFeeox12WRhlwpTjduYdGI88i46HieHgW4cGymKX2OLKRpN8u
WGynFAG/YW9fiic/G6pVE9zS1LTSnTpYtTOLGjWdehw3ToOOHKfgmw0MZthZeIm2
/L1h85oVdmfOi+VrlNc7RJVLet2sjaBRo565Z/VwUlzwVHs22QTz1qYilWAR4ymM
iPjJmHEnwI19gG7ohrND1wMliFaihNPT/V2uoYw1If7CyjJJEW6nU9F3+qP1OGeh
d8PMzw1fNGPgXR5CpGAhETmZUGvRlmMPgZhX4gtpWS2Ynxg/E3nqGUH9y77glTBu
+jq3mwHf4OVQpgiiwsvAuCvvPUE1MXu9AoQQCDo9fbAA9k7fLutmaozUnsr2I19b
3Ux7as0uysy1eZqXIR8HBCs4aBkv2nT7GbMxWTe5ASlty3xPOLCt2ED5XtlWv+Ix
mLRJxwRnPJ8azGiF/sZOfQ9qNVMjneVxFqhXaWnyFycmwKs6Y0E5Zqr/G71+ofnR
JQDYf4yMY9pfF8odatCYFSMmyPBhIxwRcfI33+0mIPS9Ct3V/DJbTkY8xfSqskf/
q1SVBIPd1Mu4poyvVTn7fpEm3BO26M8PWDr+4qfbd3qQMaPVuZ0ymDWaJCt19TVe
x5k8CpLFpaZzQBzgahkkBtxHvnZqdNtrpMSX5Ab77kjQqMtuDmSwujrDFVVCjsvw
QHJwBreMfsGai0ywW7P9hvjP4XaBGTOiAi8aUy6AIehWXKYK+5xKMnTD6IvMuuHq
3p+2gJfKDgEvz3hIgxkv3mL2lv7YXRaTkcp8P400R292wa6BSslLkwGWuNa7AEkx
CAsiEaU4l1QGPEndBiy4qaPmGQiBDLNzM8knDNEndJlSnnfelho6odk6lJ1boWAs
QmmjO9L1cIevx21yPdUdoaTk3Hr+Jzx3WGS2yW85fD9y1U59xgnrSoeNiASMMA9V
skEC0zteHfLjytljLv2aGKd57cQTbkLKNHLvFaiG1fy65MThkS7CFCTcYouaqL2y
4g3O79ujItCUCRf5Qm2ay6AYQHEEeOk40odyK5vkBXhw+FslD5770J9Bq30Q5ZuH
jYj/cU+eTAmhODexXMua2J7Yw1kk6DBkEwgFqgUJmrTyEVj9XhW9w9wUEQey5je9
os6GkIgEY9ZTI6K8GP9twFQvWKYt2Qq6VRjydRCwjf8+W4xSRVOQBbuCiYqCylUw
3gy8fMFy2Ahh15a7JCSeGsJsTnj1ut+VetCsKfTLm9ziQ8o3ikTwtPJtacR3JKaW
yNmnZkNHJ+w22CtXD1iG0vyqTIzyz9wZjbKm6j3jxNvLFtnqVQMXlVHgZewAFj/T
8uLGcro9V5E477qA2KYFrPQ97sbGWR4ioPJRdXSazIm9Usu9ypAOcMo+ntjGx9he
Q2xqB3KpU3clFXJS0Ec4e5TZDOPI2hG5B+nQQeBPniR7juoFapGb7/Vb5jx9Ozci
7SyEjAOU/Fwp/OTx48uhUFCZ16FC5RROozwoW6efQQa83Go5TLzNQne6+pwsFbQ3
XSM+EPuVCgNxwP630bweDIpTWJ4Sf9Jiwm76c9wErezoi37zT51um9CsDqjqxP5f
hlgixBL0dCzRsHzxizFzXMcyLhdgOxVvXqyApARlI/wB9niCYb7SJimXKHN1/JU6
z35hxsodtyDQ+2J/rX8f0bYUwOeneM/UYtlNOXg2IKpc/277VmrtqovxPeUw1PS0
9yxP8gxoscLFJxCYzjcrc8IscGTTXI10pn5yAKIxjWkQrCUpnxVSz04NjUUSUmR6
sqFCAoHs1KfTK/eRMFJesTtYa0aWjj9Vda8nid1Ya2FluExHn/76Ds+2OkjJnQJi
MyAJVo8phM+wY1eIzfFIoMvDvvZbyjVzZYoKHC2TCosOiZzUk/KENy9EA4QLA/OG
VHCH0G4Vp0cCf4xm8LQ+cvHpCPgZuE9xfFV+mzbLhogwn8v4hyuk6m8AgNW8zCis
C9GPBO20crqcjbtXUp+o9wLy3+2Rf/1zOHZQtCv2ECS32kKhon6OtYG5MEk7h73G
KnVXiL7KEQOXnn4R+ehKP9q5vazFRdU/XA7+yFq4b14jJl4dyOV84WFk1sAO/4qp
pP1fDc6JwnK1jxTxfgB2vj4HJFpZE4h8jLhCEJPaT1cNSf6QB2PCxvQs5rRjvHSO
M/vlRlb0Aj2cCmP6w9YPUyBPKQUmhF2TTM0aj2sy+aKzSrD6czECBbz4//ZnWXax
vWJ7FAImsB9QP6ZyYZZCJcxMo96kmp4nD0sHPMri8KB7lnqf2xWR/nE1L+iqOnzF
nbRKcDmJvt7obHs4qDNS/E/xSBOKC+WAdkU6zRsRV/t1dv7+vgRKD3liazRvJ3sZ
ppHPyyg5na+o7EuqypfNV63G+5LCeJUDiJ/aM+hY04euAp2p9AMQHHfIxPqTN7Sk
baRnGMksathhRSIMX9gYc63euFE7A245rtN9WAMZ2IPAVCbY5VMph98fhwxQ4Hn4
eowDwju7dzsJtxEE8GByblhXVSrYmgvSTTBTXc/vYn+CbBBCmlGSEg+GtyXDQbYu
N/JWW/8+3Sm+PD5Y8slIL4iAqnXl8oNcATTZ8iJPHshXb/hVpYbIXitziXCWXr1s
UzvuS+1Ksr80wfdqBhEkd62Fni3KUNF1QpXXVd7v3eGIkeLszvxRga03X8oMWd4i
/zRT9t1G7itiOHsKioyvHNmpQ6K7U7HvO4P7lTKDCpMnWYvwbVecT2XeCS/58zD9
VG2qoXYQWTGTy1GF6TXM8nEMlX1MSX2vOpMtXJlT761Zi+B16FD6DGracw6TJdzq
dEHupIz9zFo1P0GiRynz56AOMZFTjq2LLhpIhm2OKzNjVO7oAw0uo6BiAXiMFDHu
4DD4x7y/a7T6BOTHY8Q0ZZqQnUUtsVX1UDfGmdOfJrMw2Z9Ql1toHG5c6oqz2ciD
kB+KKm7rCM5U1jcbj9BoTbicCc5LHAewQYsdBFG1UwF3lBnXVfF/aJvTujKSHwcE
JvarkLXLSikMt3V7QWjrGqyqtsRBKlgFu1d6x7F8A9JvxIqwnxLaZdq1ZNNDQAps
6C2irPj8pXEoZ8AO2VcPmfatFqlwNSQPE0oLqouMOJiqE3GpT0AYylWs9EMeadRs
A8t20/5aivDt/4/YHouVenhlEecJNYav566PGs9A63j6bxjpXM1fD3VSb33Cyimm
bZu8JeM2h83t+XnH0bv13DKm3W/Yw7O0RG2eLriLFmvzNmV+83teDdRQbt9M5p2J
gQGsPx6Wg68Nph98kK1kKbop5SfGCZUlpMXazXr+bsn2mYEEXrZa0huHsJY7FVDS
7wVXtVUwAre1OrVPDKeFA3OgwHUxwgNUhWRuSLLU8MnL8h047QZhdL0Z6C0/wFKT
Zhi1rEU/AOCtjpzG/ynzyAuxKIMmhKUlmN4FVFuYGgevLNhZ6/AfpQmg1wZ4zhY8
AQp2V6lVspFxWlsBTuHyLSOtu3nsCNhciMROZxDVtIZOD/7Qx4fV9Ys8VnYGfCFd
MP4orajBADSfRy3xMKikGfE+yeoO9f9pWcGw7SySuzfBgWsrH+vWVZi1bnMsZdmn
qAxBfyIjZdYfYfOi1HTVN/uYgBPwrkRF1xA8LVlpC4yPEvoKlpnhvpm8wn0VZkAg
t5r8bCPMHghYJfsYiDjTrIdLYM4zoOxTG4eML5rAUUerW1/T1Bf88pfP7gKp50Up
Ed5JJ00gkcOeljmgnA8pk+Avr0rPdl5/+RP8RP8y+ljxQBQgDnY0b5tYmIeZPUcF
`pragma protect end_protected
