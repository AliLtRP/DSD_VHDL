// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
EKfGQJV/zhbeVTee5eUivpVXSHm3xJiEfbriJ8HF5Oj1nyj00XCAN+7xx5uTHkBqrb7tjRyJh1sR
CcFRiScUpfES+jtNARYoirX1r++03e03WyQMgIXKZhPcXOmkWLhu8nKjsLCGySJzIxYXwYNFZIs4
kU3gGNY19saSHyxw/YF/eOKZ3+VLmgYiuVrMPgcRe/RnXIwB2bQry74isjdsw6YOxkNtKwjGuTQU
/57jbp1Ms2pabtJNqEUZnGswNwkysV2aUqxLftKsiH0uhFRgnTPuQ4foDFzMYTP7FT+LUtx3qs7R
5jBLx+3oaiTVtkDAwnwEQnJqhnzWj65eX8oc5A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
XeLNOa2qjz0ny3yDMcHs4PzBBcMosCluCqwU0ZCRctKaGL7ZPa9zC2lPg86pgxPt3Z2S3q52XjQe
nyxCQV7qrG6Wa5/N7b2P749+akjya2fs+OonpmjHqMZZng1ODf1jUktdeLyc4mxDCaSrs7kaB0Yh
0WDryVeT9lvCGH+zS4UghAs0l2wnlACwwPjU9A9tdY8VLBOIP72sQZqb52zKjEthFtA04taz7oPs
ThgFNahSCafucfV/L4BP/9ks9/+eaDHr82ZY+B+Agx7h6zcNy6GoSAIO1loA6/6YMLBouVntit5C
E4CRgs5LxR142MRCxV0FBcD5pi8rfXsOrpRYSZg0HGKBYT0EuJZfhM8r2bKD3+py6tOUV/PfAZCO
hmFeg3RQTgtVg6rEhmTK7NLizLebG5YMsuxuWZBowsfqIQww9SaVaS57Rdueii4DXhh4Qe5TRcB8
B/uJa4VpcOHYmxk5pgTfhFrcqWMv7NLsNdYkXWSEBOPmyMHMhZFUYv4RAekH2iXfKbksfjkSf3k7
G/l1EwM2uoQzz7JfnF3yBQJasqf0hVCI1eGhHAJ+RlHB4aZr1wINVSTB6fLShp6oKxsRKVJe/KXo
pSz4TqfvJNbWUvjhQEAmXNEIFOlS9hF4YDLKSubv2WHbY+bu88KWpmq/zZfm2P4H9Z7s5Bz8+wBl
L5i1jgOmizS2D1/QQbpN8H4Mn6sTOUpZNU9/u8SeTDV1hJeROnR2evfOSkXK2uitYI4/BBfIFd+Y
ncOdpFUcaV/Ebs3b2D3ZFum8FvZTRxGUEHauFzAvZJDC4exSNIpXHFyb990vCMlqY5oTVfiGHUjw
3e8BIkvpqftXBPChysSYl37BdA9zM9hJB19k9V/n7h7SrLNeEvFuhY9/wEc0AitaT2S2uWFZxsgn
UAqmZ+Wy/zeXeShCZKTfxp4Gh7VbkhC+5/+BsmewgIVJUhhBaUOnGEo146mH8z7qQO1WxIS9exj0
QCKZu6V8BwAmD0zTUhMZ4KykgRMqwssYoteZrZwitgx6OGRIjyXDpnuj4JdMDupNCjzWbiz7kcWk
5i9p42Fx6Iz69Xr2GZCMc2yrgWdgc99XRs7d45FP4IhPrcSFfOGvadd2R2Nhki5x3dKZZ+OnF/DQ
vXmrNSkHQNKqIYAN7ijm93FtQtn1bMjtybwJIYn9NgzTiKOmfghxskKKCnrelu8MzEEYAKGyaffX
mt+FsBAh5ZxwTs/bFjsTGqjogXTMlYVRvGxe/HDWENmOsQdau1aaoqhjC+JRn1NSI+vc1vb+6LIT
ZWUDT8dIfb34Vsejro7N/JhJkvhkJE8gdDcH5c8wDJnW1qYrSJIWp940Kybjdjd8hO/1Bclmp8No
+9ZS9EOYzKkizuM8VnMUzU8mK97Wi0XUkjedxum+pimmlQTGw+R0x+tr920TPoNIcuMhDFkXsK0O
9axsJLsAO60s4PFFXGxeFVbAE9RHsmu78SqtQ84fGFO/R9l7RkWSM4uhl+z5kuMSvgBBDMQx3PP4
c4ww0rjOgscBIo0w5FwaePeEOY62sChujandCdEzuESgAG1JUA0z38sknbELF/cAul/jBu8Uq/cC
8kUte/fihiBru7y/9Mbcn0+9Q7kInXTNVSFlBw9UqiqQbpVDyM7FwxZRO3YwkDteBG74sfdP1x86
WJzLq0yAMuqNz+FDV52+SISl9mU5bM+TwQNsFt8RdO7G0AjsvDfZxJXNGfwLajx/26uxESYXbgA4
HvaKFMjMSpFM2KdpLvUXRLx2i55LL4aSnQChs77O1GK/oul8cHpulIF/pkmCi3W3fRXTrYiNMvqI
QaYuBlHxRlX2B4ca5Xp/6zz5gFT2V019+bawmCoFXB05qVkTJ/cFAo89+KM/V04qAKz0Pu4aWDqJ
tr5XWwlH3rRlgI5hhioMUhNS1Dt1Oc9pzFDSjok0JhtTU2d6Ymvq+nOXAUiOF1bELfDVojoNPLSG
JefSMqzdlG8scLouplvzMLWVp0LRys1c38AJgO77vCBm1KC1sVY2Ja8m4rGPC7mCtuepDS425qNL
uypLdOlrVU5uV2WoVJZA7mgW3HEnGMc+/ZtvPxkWR8VfoiZzWNY7Yzw2yJSyDQqCHRAuZeiJjGPM
rxQc/mojsudVY2Pp12vaGLATrMwFBnmc/IhBIR3fLuDsnbW1pJUNoFab9ge1Xh5wKLyhSdYDOofd
LHqBo3Dn/a3HtSMMnB6qhVHf0mRp1ocOsIJiHO7ZwxA9hQgActyPXMHjMl+k7Sk9Ct0/kioezbMY
R6HniCOQKELLkUROO5VhKwwlSIuGGqj+7EkEwrXn2GZoOiWZTvdd/IFQgrpczEyH3lIVBugftZnz
3Tdhxk9QqNg1OV/Ho353aXZcQ+DJnXEjFYmhUBbPP0suqC0sjZ1fb+qoPybEzaITmJPAlLc1nWdf
ctoCdhwP0Wttu3Pj5ADBgr5zgjyZ0EwXbuwhcgUytx4CLrsCqp36HzfvGO2gQTy33i3eB13WPxKq
n1+iCI/c32OkE7H8BXKbvvVSCOdU/3C2J9KHkCNl2YqhyBcMtNcZKaff2AmLIcTxZfcD3MzBaM1E
I4/Mp0h1Xdm4yFwvui43KT56ZmALgSSNstenqcwpw/7uI93zw9XKUfykIzdbCXoCmBUFiORHBFKt
r+3XD2WBkj1OtIIpfJnjfSQmjzS+YHOcSTsLgtEl+1BPgYaFj6zDIu5tvOO1n+T7KyVzrTzpzKkv
+wyDjp711N7VXFz3znRDdJR8uoR47/wASwYm0DJ4xwzSVuBurAZYpKDu+wQsrl2atdcqfE/leZIx
m3DlKajDWxc/k1ZxkKlKSxIhFirqV0hFTNwI0nWjmFfcJBUY6v8Q/Hi4EJrM3uXrQCwNPFRjuZhS
eHnjY8k98gW+OR7RNzuCuu0kmaZffM0aAcV2C0oLdQUZJETiHNvm7PJgYc//FP/CNjiQ60U/lRdg
gE2QC7MVQpPobxB76BA0a08TAjeuXnJl0/ltuKHHZ5M/EZEnP0vwwe3L1NyYWRi0LsCmHgeis3R/
woPMcwjaf9gUp7brVYfdzjotdODLfDoelwQmab9U0Wn0igjwX8zvtx67XqgBk23Cc9YHebLqTQE4
H6OKEsfGtHKToseLkJ6r4FXXlCBNaKvGCzmlL6IR73zjf7hbTQbmcpN4XD1VbGsK9U0DF1fS+pC6
t4qxF6FEo7xu3OxxnlSxjL+th6uAxf5/6LNvLjxEXKoe8vpJh2FH2oxPdEL3jH5FHzqCHctuvHXK
5X8jJJ1DdhWJMj6rtkr+1Gc+LItLIhjAfE+bNzVlr4cDTZVdsMtaAkVAhZg6yqqzL4ef8aTDQ5ek
n9phWlFuVhGadJwPp+Y+s7sZ2+Mx7WoxBvAlg3uaVfsUYtos0+QhhTDcU52YGgZ5i0l1dNaHO/Pv
fVOYa2y9JIUEifqcaHE3q4rhE4erY+5mi2N5y9h5gup6OTazq10hAAeNY/ivtswZMQRRQUFchcgF
rXSci5wQDeO3CJLV4W3UWiyTgeLAQb7Btxvt5w7TJh0PJn7geh5UiaJwOTcl4jrFoTQAE5MtBERK
cdZ+qzKg/3xGlYE6S2U+wQtHsHnpg5OlPXL+lZ8KvthoUyd0RH77fv0LkxeENYP/VDOeaFLTUtsh
7TVD7IyeavFbe+yixlz1sp65iW+b0DylkiKOYZIbwRygAuLg7WF/bsst1pIh50joOBodZfXtjjgk
dGYtsAxoM6bUjnPxqbCm6sf/jF/WZO2WhKV6495jci2GFyk2v+S+GNqaTi8KgZryxNKvdUisMed5
ZPAmrhXxJBWB4Ks3kxOiWrAGIrh1grjn/UBX8fEsx4Vd5+t4D660cPNZZmYtZuZpG8fjnEFS16Rr
+rJqV9vqPGM7+Q14CY28fa2maPdmkYmVf20E9pIYbo9OnxqNWM/r5O9eotkDfe6iZIDK/7/utOl3
NatHApeUlEewZNFsHEv1cl0jsp26bWLbxFkH1sobs09zF1mTe6YCw2Sv5YCIDNx95WzCce5fiCBk
B7WKdrnGbWP79evBWelhpd1OS5yYu3ogetFHuO4kFLRj9WC7MpHAfUCClUg7qhIwr/JpAO/3KOvQ
/C8OmDLbQ2uXnG0o8XmdvgpC9W6qZU/KpFOXyDWUkJirY2kUFiYIqdAIpocKs5FsN4am9o3BjPbV
aFnd6aGuV3EgXRpE+MTXB6FujKZUfz9b53ECwO9jfEKtZHDBB/QTFWjpXz/FEIaVYIXoAdE0L4Ys
ewzt8a6aBGk0mLk06JbQ/at6hgs+e6ptyA2RkzwpDPM0iA4musSGu1JO09rn/ekmP6d2u/1zEVZq
18vVP3V9/eSWEMLMGzQtxP/yAGhD9L6wHnP3fZTeAcSY8Gire3puSZzgf+Z4GKsorkqKGqjLnTpw
UGgwurxWtPDeJtloIYG5GWFtPHQ6RhAI755vkEqearHuPY03MYq/MGr4E9XamqVHWGxgsb2+kBGS
isrFYzVH3yzSqZ4WMv/hLESXHeLiF8FDXlFCUn+Y7JI5Z6P0Qygk1yYiO8zdwZCGKCCqT/zsKmJt
jamjSwSSUyogZTPWEgBHxGpf0AEZhLbmrspmaOcXjZdgzO8GJCpIpSzHnyBAOwttGyTpLYvMr6ta
GcLUZP+tQNx33I88Ufi5EK65eVAz+es29miXXvwb6jau1MZxt0sua6FmUuOuK7nacVgvUNWEI3SU
NhiKHTEcLuf2yW/Tht0p9FY+unPt4rW02fic35hvEHLeWms/LXTd8L/37UzQbtzRdhaL+fcuM4A8
VG05YGSeHvopH7f9TXvKLokwAtPa4vGxSwa3VW/rUg1MBbCRKqD1orz3N8g3UywTHjKeZI4YMIoQ
AGb/ZMMbMAl5ZgP874qyt5U/gkBuNHiVYq1d2xoFK3CbqhCHek90YQ5we6oiN8IRpaeV1d1DxpMW
MTxveO3T5F+rbblZ0chSNWV6L4cJuy9lYSB+q0YS9elIj0we0tT9LJt9zXZQNm886i86xzbvMSn4
nUK39AlHUdhvJEerCtz8bp8eOaZsT4Wx4jxZMf1HcCYGSVBU+Vc9pyczxWCUcxZ1febNnueabL6n
pjw1MzYn2hXL+dcVXTXcNGBaZIoIbJ2q2nnq8gzSJlD8+shp8Re7oNoidtk3UF5eos8nV7/clre2
I2+y7TqjQd0Dm7U2/QoLk3NmpqwqdlsUmBXJC5MYQB8NrN3d8JOqWG5dLk5NVloP6US4FydWy878
jg0E9FWg1iDRXOo3BQcbEehZLorBHGN1n90sIg1Dz2RAi07XNCXVaeCuMdMjSIVbxMhUobgYqc5m
NrtY+gsyTgL89C7y6IPnGm7Z7oU107lgB8Gv5gkurK2zLUWaEHE+Y5PVps1gAVEVXC1iYVsPpRuI
ZMgt/QAwCnQqR98NBD6c3L5TtaiGJ3S88XUZLexXfWO5fZysTPoG8INcJoOVvcOMqqmhzDRfpCc8
fPN2gpcgG9bPA4xQgVI9clm3gKllY+CBvCpaKMD4hR3OV7ZbgvQo76L6wRjyyqwhpNxSn0smLmr+
cCOOBMnksYxenC06nOclOwjeDiED3RBctgntspaj5DhC4XwIbl5b4g7aQ2P3u17PSy0mnM5FcvOj
isR4/5mESm9iuvcevz7dIOU3QSMI1S/c8qMf4pVvPkn8kGf96wo/aKf0F33O8nKhkJsn8r+IQz2B
qQT38BvM9oQx0wxuHKmOLouL9FxeL3aoqDSXY3ZrJVmQNFb6td15M0cwCzK798PyjsSSo00VuvxY
UFYePA7skJT+PR2j/+k/AXPnQ0gL2StAXHOTwJX/nNySvFKxT/zmY46tYK+APqnhZWecReF7pUvB
KqmAMOVQeC32zQmF24eaolpn/eLZFuKe2xCYciXfEuRC6GJMfZIj0n+T0a4RsHpAaBjkHdCucEAo
Ke6IC5oXWwgC0k68V6+bDZrIW9gkgmHeidOXj96V5Z8YNIetKRsbtvFNYNoOlbZ9fkD7yFXp/ws3
CEnsrHZ9cE0uKZxfnkTDAhSu15AiORYsO2rFM+CzMB9rfNESdjlERFAoesZ5MMhmdM/QhAOxFvyH
fBOarzqVRU+2noUobwORHrMuPNnMDZDV1l08sd05DFFzJ/dfZlSac/NOdNkyO/pBykADsOx+Ohph
xqhchJhFN/ovDhNRglK5UfuaeAf/WlHpDS4QRYPNvrv2xcCCfAbcSOVD/VBxj+dlbIzMACNvyLQz
NRKPmX6C7z7QemsMN+OgzKWWjhpUSc1ZD464AOtc4Yb4Trmv8Ekv4rcwgnH9+7u76p8heo+Bt8xH
wD1mOSitvNQ8DUWtskFRhN6GWC+xkqEPGSLLLUeTbseRI9qeogBrWI3lxR0varvDDGZWH3xpMTyR
MERWF0ELxdclqLh2W8qUzy8vGSfap0spM7PILf1hw4EEWyQ/AFHJWa/jkHtkosHK8GbgPBI0E5NA
C9ibc2a8BWatxNyzoP8GDziP39koYkbjDW6dATabCDNIi333CSF+0AcuxlRzvkanNGBw63VdwS89
pgqFZhgsfsRCFjhi1KS9En44QbX/RMcHehVGXdyxSyhFufe0SrdNi7wB/54mJjPledNIYEXEOJ8w
PUL2EmTDNStRqbbFZa/sxYvEoSdIwv6c0GsLUqAuAS2q+yd4xwdZCGITWURoPM5jDAHV6kVyWkfJ
hrkLb2oC6kd4K4Hjv2mn9wsDQUGEeOEUIaccOASUD5PR+RXuwMs6T77GuGMHx1N71wudNo/CaLXM
NVgjq4m8NlZPGfYr2LBVCObfa0rnMVZ4J5Q/+rzWPW8Sxl3SsxAr+nNpInGyDbN72nLBfvQnxj+X
Lb6FZ2u9Y9UimbIrqfpmHFdxSaXp/AEbd1pQqayuyCCokXKLFXln8UEKxJjg/6E5DLlmbXrLEfBn
KHJLefMssVnqyRg71NHQiukTv6oMHG06fKb5fw6VHCa+zFfKNviJ9sU1gofoFhDvpcHUqdk5oDdx
PG1CtqljhtBvSN2l8tgGxXDnk3JGiVL/yYobGaCRC5IlFZ34+Pgy8Xg+CqGgO9YKYE+M8IqRJlhN
3Ct+XwSXlua73IiA1ORjGYwWrHfJB9KAfxa/aDhP3bnGXUXqgHGgczeYUtBMAUNpkRThWfy5GGKW
WDd7TDy021UZmM0jbiLbKXrfewUPT6brhaPwDgx8gb4VcRDrLpWeDL7y5uHWyEw3xTcAj0TMOveg
8WPIDpaDYVby2HP25kPLQkeKDEMwZ62/dQFhUNxGYserHwus+n7Qbu3eEJ3vLc+Ek30qYDU034YY
eJ22YJ2glyUpsNTF68JhOd/yKLESrdCp3TJnN+mtfczMw2gBR6DdeukWk49E+caVmcwyKrs/uigK
if7Fd3pB3HyQBlkDNqurwPKfFxqQeynvOZ6j2Jwjos5m5e6yidxyT4G7My9fzwW6/2rcK8xSLBQj
ItNUJuiYQxQXuwOWh5+eWWCEP5FrQEkzOK7mMUdva8J+LsZ4VD3MbwP/AQOAmUeX80f5ANyQIJqB
qm53qOfMD6guXF5uQYXk+el+xvPnmn8BzbBglrVPpNxOWgMdrOCzmwSDu8RQBQjKj7Co8O9iRXBx
ta997a+bctCtYzHwR1oAtdjXSbg3hJ/xVkXXhbB2hlkpcJUvCb5u6JOhQwFtvhMSv8dfGL4CODPk
T4XHq823CGQT8XQ62B/uOAenORFC0kEku4QFEi4s4b+vIF9Yrni3Lee1Q8VuUHcfIhMbypu2xV/E
o/Po8Yg5UdEik/jfg5zh+7dvGSMzCDxYtqIAARImdH+t6iahg2LhaLMNud/fag+ed9Rwa9iP18cK
DANm8q93sHPtNfVT4ufyTWZdVjDI75x5wtVBJHjTGli3/l6UAiyVJRkFpvYOB6rIVkTq450owwOp
VrJm2gZhn4HKprX9gPXws9NXtJ9H+hS+kTb/x3G87XyOLoyN3XeV4swet8DVaf+A+6zts5t/oxmY
jQbp8QQhs7M9yS6gvTNy+QPbtebr+lByBsWEgiX9eEOFyUP5zlMklm8iICAXPtkhN/SrgDoQVJog
d/+Yh4mQWGwLfTzKIk4UKyFvRfpKNT1Vbuis0PXNfd0tBnBkeZGN+gMyo7cf7qL8LRaV2ok3UV0W
6BW3R53FrmBf8VqDKqFqW7EKdHZll9C6A/1SbWcBF+syn90OiGVapfOUNoMspxQSJvTRUQGNCxWT
wEYE5vmDC/Uq0DJYQ/zvRijZfq/3B6WrAfCkXxr8R6ZLmNOwK8A2NtFkG9343IUMXYGzwkLWe9yt
BhLGnT9USnbq06RGCF3Rq2MDWKq/bkrN6I3NzM/HTQm7W6hr78lFBNplC3B9engDewvoGUSXftyS
llAJaibrVuWq1quBZFFPkiHo4aM5U5c5YcwPC+Ddk6ZnQ7/hpTY/8HJSNz5R7aGHO89yOt42krTi
zCur0KSD8Jxs/NplIIgQOxfr1Kzyv7JZ3WW7XdI1M5ZYDxxqkt3y/kT2+x0tQLGEzbi7FhgMgXpx
WtAbplchqkN4Ct7924buVzaHK8Qs2i1ME072zyZtaITPI/2gfE7FYPqJlaubr9ibyV9phZwTn9PF
Ax1xMMIg8Vj5A2qb4YcFvuQgGtRa2ikNRJlyaj0Uk8VdB8ywbDGn/iW8ik1h4Gr0WV6kQkmG5oZm
oJ8ITbtMvYjX8s2jX04nfB5fAVjFrZY3oa+SaAdbBD73aoJ1y1IoOsC9I4zSlK2BEGIrvv6MHAfc
fI8+TqvD0sPOfK6QicjXSmY82KUqjIvVGRyEEqwTCWGLzMBMfcN/QExZ15o+6v6uOh5Udq/AmDLO
aOX7mVOVUBkk+Tl2doK5GoaupKQmX0akNATw7VpESq/t6Ba3WOrUNshBhMLYrJwplj5+oyYX9j9W
A5rnDfOXJriOz9fbsD8jRBcgnHxSJl9KcOj1IJQ/dGAYB80D733fTR1cSJxbBlOZGbuh6D52u9tG
CSdo1N2fLKNWmxmvdAqJKzXWl7H1s3eMvHuucdxZur+BqlujM+2iIqCFOKbr67XnrktPEYzS7H38
sjnNEE7orvU4ntMK+Hb4AKkpkvXGymZMZIaW5S/Wg/F/pybPUUX7MxXC5lO58dOtyruKXDQer2vb
FVasowtlLzhbRPC14I+/t9bFd3+H348tHn6GZ6YcZziP7JY0W2HKeieCmGfxpNgsvaUcFrSdUD9n
A8YXE/u9bz6vxxlP0PO5aHByCLWSQRGqaCZRZ/UeZ/j830akmhhaGmET2gIq75/Z/WuPQ2vZPu4B
dFxOzC+TSWZhMhOHwQrmIxLTIkmrZ5dJSUrD8mlSZ/eV/j/YMa1vId2yqwnHyASJspSUBjM4GUT2
glCW7dInENZQv9Fawa5NFWI9p5ZeBhnYIySHjJJmHycoJrketCDPkKvld+ihdXN95f1hz7rhsmhY
hYWEgcXepvbx8fWBv6LDKpOqloeuRDtT1MmtdiLBGvD1+Ms+51ewKO7nSoFpPGqIKhVDI/mRrcBW
LkZQtvC8ePF9hhiJn3rSqjimEQZ6WHcn61bjM5UqGHViW/la7ceI50ENuoAO6z0lkBAn8XE0XI/p
qolfpD1Q7u0BF7Sq3hsvSQHyQwP9eJGbNnXqyI6vkqtaV7t23Je0met8iM5z3XTR70BUoVDV2h9v
p8IlfnnIPtPihvfBJScu89QGom9u2WOK8tZgC3peIoa0QbKeRKiMph+PrGEJUPVxsNVmHCZw2WhK
axPkO8wj85nSztminBKv3iUiicjJwy2nheVfgq02hTiI7X+15zMf4LN+SmGEFtAUfzdwxP6vP1xK
vtWHHfjvuJprtR2o4U4pZCch4Lkfdb3yDaYAb0nOA7wGKvEuxuIgQZ8xSzrJ6IrsiMdvH7y3o8aD
0ZpsrzPXov4/Etu6cJ5eHU5lTbKjva0y0g0J0vUWNAOI/QJcxlcyOmx1+5JKUMZSDyHPNV8oxmti
er3z7Jl3ZW2jemNneGh6BzY7/A056SAsY0W/mTkOqirnfcsz9zE4v1TCEczU0DmcXnEbgj4SWtUg
W9nem+41QKBCEQpRm9CIiMy/6kj1KFvUKuwG9uOkjmAERVm8x1Wr2kgVXbCa05UCu9P83rp8o9Ef
VpajcHajBs5o8ysK22TtsN60yMmZpE3py//fOhbiJ1VNfiP33ssHSDjZTGQ6Qa0/EmnRS8x07HOb
1rffheQwJ57Wn7M6Fi+oaK9iTVCddGojyrD/7dVZ536Ivw0MAt1fOfkeslNJx6orqS7XoTGfmwUD
3dsHYedi52MPOUwtt2BBignsSXgJF+JOn8FacDoQ8VudoG9uW1F5IzqI5h4/mr018qJcnOiXaAlw
5KKhcEoYypKjZcm2lSRYCE/JRcYU5MC/A4bdlr9yeiLvv31o650Ut6QCvPUQRgMPQVvP9HsZlFwS
gnIZIAnzKlbUncmt3HGFmdskcULtNhR0+wHJ87K3R4SQ834CqdfZnQuJQ+3wFvxy9FDqK1divLX5
cxYKvyy+TGCn4KA2WTS99INty7GvAAF9vLj/9xGwUzOAS/369/SwG2cVermasEVnb0RCi4nLgtvb
Do7JnqGdpFMsTZUo9rfjJwEkfcapbdzlgRyQQZs9xcNEq+zZUBeBRRTKBZ18V1flzx9KYvxr+kZg
2kpu7rCyApOFWhWdeG9tHY5Va4ESnPzMmAPWWcWi6Ssc+pHzXJILQlGj0lmbzmpfGlUrREg0rtbg
O82RH8mfx8Lb2M7fgRQ1X0sPBGkzdqyJP2oqcFFJ4Qvuicp2sUHE8rVK06quyhwFYxyXTFA88I+2
v2tnn33xAXrqF4ZkV2zdiyofBfZ314i/4iiFiEcnbSttlN0qdpaDEEKZMJqzCjGyqfuHu5AHgCf0
b5fvOgqWIglda1b1Tyug0VhaecQeEEANsjjn9Cf+2MkpTsTq4G+7nfLb4g6toAswixhlH1YSljdn
qPo29DuN5AEmRcslWhRp7U0TXpMNrVd7ZKNe1NQRYLML7/4zxy3hnI7lQAr0wwwupf0D9xjbKT3x
ntadmiMRvoXmUmfvm4nBUHhawPavZWazIeBt4JiWT5YaBC2GEo3b07DA7Kwg5PPGVdQbFO+4dP8h
4EUKkmrRfq7OGoahjT1LAM57AJp7P0b3qCahHNovIgKMTDhP8iJvrdM8mTBxm44na+H32ssYaUw2
IXazgTKpUkZEy7qRbrNAKZMPCqgnFfsNJvcMH0o+Y1fI/P701X1xFckBNLafAq4MchgZtbeiJnop
b441wmGqcipLHetmIR8Cc16lhT2Rl8yRXbbOI1usybOBOD+HGCuNvlyd2A61vleRPIPKjZbt5WkC
fywOvMpagJ5eb4+yUH5dPVnbbb9UZDKlM/Ltkgm68V8GPRr0wr9wR3H4b1AV6/iivb19WmFZCbIk
hQQcpTa6VhVwjDEB1sIOtRcAR8M+eGctHGYvUnmawi4BhhTBFgGTvCYBOodywXJjB0U97ECld/z/
t8lr0uZ7q3tj6ryywZdXUPR0zbuDwIpmryseetN3nPyRcYF3XuscsWiOCRzzcBaMx66S7DsVaX79
SjjJyxesQeWcfFidtjjTrJPUrcSiwXthm/wfu7CMHFqdAKyEloCq3E+kKZESQ4uGePszVtZoENFk
PGYtgBr+VQjp8lzAoRNKmcxIXrVKnR5jMqCDSuvPC4rOzRDBlJFJwcTwa8LZA636g02mvqcavlCF
QHRL1do+7E0XZo6K9S+vHuiuT2iMNWwnsXFRbvshJgJa4bTarLRO4a2h7/GEa3s6xvOVzDBhM8EZ
h6zX711jB7qLTcTqLpb+Tt/N9qQ0G3PFYmI69JwKUo+rBncRLh420oJwlvpCoN/tTXDazQky1hhF
kJb8ddOuaeM/iq3415rS2dvrHJkgUDpAZ4IpuDxaBN4C1EyQnv25GxUwb+dcVq9mcSDWxOKRkt15
YfdoCgWe+3jF4Qb1dkJIG680FtwJ4yPJg+InmWy87X+G+9dYn26XqQKhyHRNq+oMmuE/tZSii6iO
FCbsHUyVWMmkl+1N2kXkU76lC4FhP72Rwr4o6R6TPs4FTBxQlyYSTt8RoVOWZoQ6G6+RX/g3pmUu
GGnBO4jz+sdMLy6z74QDB2XIB0neqP5sKPbb3y3mfRuLBs7T5+40oaE68TfxgTfGFoYczOM3wKIw
rRGdNM9eRWeNixSzj+6aLxOHbFukMHwqKoFBBoDchgFBF/x8gquZhiAM3rcE9aqWBR3dH2iHT0x/
j0/TYe/ik53fd/Eqwh+7/SfWkdvSxjSwX7qfznQ2FboZWVD7VWAuk8ccl4IpbMODWbmUJTLN/6V7
jqRERoFb6QXnIhvh8pyCCAjpQfFW6YOL3Sj+3snbTi+zp9WC2Erl6dYY9ELKKmKpQkaiT22y+ri7
FQMlWxH5AadH3M7lbNDgvsmgsKM1cwcePXuTZeg8sQ8EJPl9aUqyAlbdy4YEBI4FJw4zfZraaJ8H
NvOrionGWfOf6D+fvNmR3/uZ6ykNTsyhWE8rDesw0k3XnF/vjYQaNE5pdWoozU6hiLstQoWLlA9V
xcJLj/gTLV997BPBloBwT15iT28k3LWjmUwH/xbq7i4ZsgLhYeM5gUlOF+TR7CKdlTTAXSgk+aG4
lQ/uAFaYFLdLS1W9eTMBy+GFTjEEu8u/FrUxgodUFbZJb9l+tP6qpz44NFVrB9duRw6Z4+hjbC+4
sr/Hem66JnIMxGjlgAauQKzuZb+Eixt4WzQffZwiZyG+RY2exOWcu3RJX9574S2hPeTBrfZeTw//
akUb/f10o+k=
`pragma protect end_protected
