// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
A0mW9Liou8swJvQyLWIIKRNGoDsdbZ0giOaUlpuzvM5DAtdzayoC1c9JfXTkg4j8FuvtjKgapKJi
qL3OwWgmChtweFJ2eTpQL0YtLj0i2+C2J3rNXUyvM2bw8UojyrZLMsJaZZGSTQSyy2zgGXMbebl1
Ht+1opCFlFKIAp9VpjcwXAzzZdO3y2PFocbaIF2uJG8/IlhVdPDIoiLw56DcLE41GswFiodefQqY
+op4+H4PyEfP9QEtl8bdK3XM5jcIDAaE7XH/wrbV4jPA8W2JCFKaXoxzly2XQ0NrlI/2Ch2C5ofd
s7vM/CRYRJKzobGBvxN6rS5/JhH0llpk9Ebmlg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
hZlxrhxiknaj1eP0LHPQRchcVHEGPP2G23FjC2x51LBOAKqiZ2ZVtScSmPU69WCdak2fdISX8Y8p
pll1+h0MiE1Zn3WyjZ5SMeBytWyYJGaImnv/n31aD0bxNBctNTSqVs40/O2iYeLMlibedQqLFzkp
51F0ICF4GruqaVr6WiffISHwvhk1t70t0K2433nQqtOeVw+QSuqjSp9FFFCNkD1Jexk6GeknMA8j
4fCNwmXgXTr6oWLOWTz3LU7WiJlsz36Ps9O/eAIakIyA175j2bGrn1u1U5mbqQ+HvIstbBDYS9dH
FSW3XVzMvKSqpavnZG9FY4QhBsug1NJ10DW4/x94F+BTblBefBiZeexlX7Bxf/yQYhMSwy5i/+aZ
w0Lkcjz6cFLoZVMprcVedle1ZHJK1PoFARX7e7wmSZR2141X6ga0NtD/8Rstb5ZCGG47utO+rBRL
IGT03+r2VbaD4L2tJguJeeH4BRbE1WUM/YtoOk2YaLMPX/J5z3TlIUsgiArpg44hIFx/V2SJTI8U
GVytpG3zCvjdFvKQKWiqAXiDkxD+Ho9n0saKgoDfQ/ub6KIcwqQvnMpOI87ncE+3THp2c6oprA/r
LH6yVbD9vc5x/JpyqAj2+IUZd07exxcoJGVKTHExhovSC0Fxjjt4I0IT005c/uUSwGYgc/RufkRK
yNnrP1uJfCr0RSIAhL8JWAKN8sAt3H9sWAX1IKYvRxlZECXgaaoCQfZ+7IWrBNXZ/Le75umjd0D1
NfABWqNbjuY9Cd+HqMonK5XUU5jTaSgG1eG8yw3xLcIHBbp7zEShZiJ048ijhjavJR/NGVwQFytr
LZTUx6M3R52tZbVCENAcHLPMKxUsfg/Rl6oMguOyZ8PMok0TPzsr0I2H7tz93lBnxmbttw33cKg/
1SAZ6kFZRNSa7Nz97jhWezl1MbEKC58/QzturDEEc2CEzDqk3+S6ZS8MiMox66l9qoQ8ZwtAZ+t7
XbS4k546s5Q4FNkgV4xsa0UxhZU7BJD2gkk4j/L32U3eLMbPvH635JNHlqXp69M6Pen3kFvJLmOD
IokB3sO07GfRrB9/BYAWWjAC+ZHEW++kNoKGO3UOVCFb92DVvZlU5PZb2rooGc4zsp1digpuWXuK
3U1zRyj28kYph5SKpJfbsw4GAhsNTY3FbcVztJzAn5Dt5JHNccWkaoPCYd1aAOJNSHhXiytJNfsD
D+S9oHEmSex+rpHUcPwgNuoHgrQnjSWR3m/5TVIe/kcZVoylVz4w5OhLoFz71UImkO9/bZMIGhQx
oG+qULIBsEaQL0zRyZfyiINTCZFPmx34TslqDDxfYBifIEI7Kse2c7zEfBrfyV8m7+EgQ/PK5WQB
0mqsvFX9uJKJpZ68lfvhJDDWT5N2QGVBUZK8gjiek0r/OFlU6+Grayc3Z2rW0NvP9lWRdBTc0ZOP
DfrwGF989TBlgUqBWmef242ej+lQCPgB0gn1S7+vXxGv5InNXTjQJWVTsGR8cfHBKzDpQ8averZ/
qIVmwBMYqziHWZgvv26xY0llPIp4E+Pm436BXhH/w9qQyRqaZqWVu01UiyYzYOVHMLT0kdfweFeC
/A90Xj2qEXywQNdK2VY3QPBH6LSPCyuxUPJa+3QZX2NRaFSv7/bxEA1yLrIw+SWHWPSEfXxZzDaE
tMbje5pKNqt2lAVMkJTojmjux1jcbTUX2bVpPOyoB8cGcSPMukzPnGUtniH1/Bm/BlTYtYxFxGhC
SsD2ZLQZH5AOJjXCr8NSL04XUDzeTSEFpAo9KEusRwjeurLav9T7o1kdrNkgmVkhWvI1XJmodpNC
6xpQeROG4ue+ZJFpYDhBHv1/THD6c60by8jjyPMa0k4LDY5f6ncEv62qKnwkTq/cdJVdV3KhsJHA
2kZYyvHkXrh5YSB/R6G/9wzY1v+ufi16j59dlEuo2wszJVTe+3TmTnJXMpK/d9X/q+F9c4vyKHtb
RzKQ0fvD5JAozabxZUGtF0xrtEjlWs0TETsGEZYxnKcGHEt8XFK+IscUfSBt/Rt+LetW5OCq39u+
K3JMumMzlDovi0B1dhu/rekwM418UwDBa0eJ9ji9Dj5/cuoaWvQHh+iWntTfcjRDDaG+iKMQVd7w
R8C8sm54sALk6b1lFZ06If5ZKi06Zetdtayhwb43S8kfq1MwV2LbY2CpbEHBJAdDNGoTzq5s1SKr
kA+9m1pP0JHMAU8SdEfTWXYDoyCkKzZUMxwrl7qiyrZLuKnV88pfZjV2cgoFKWRybwYw2G+3gwrK
Nu0W8ff+QVtJA9tgalfcZDkjp1NpDiQlW8heLLM8y2Jf32tACgJRcbxdB6ieS4JkWVYpuhc+wu2y
7U0kVYHzcaRxGvySYKAuJhe3VboZDC+WAuEcS5WbVlplWyMsOXm8Z5qsbLlF1/e3e+TSgfvIGdzf
IRFoLCYKGK3gNKeC2XXMZMqxz510BEeoE9wqETddP+B16EoUhKYkrfqije7C+c3GOpnlfSAyM5JE
XcZ4n6PEFgcu3O9O3vGd+COYWoHDIKtlj3p3VGEjipnKC0rkhpvk+xO2vrDz3HwrR0QEjx5HpDLt
7uLtNwy839yewrA4RF2w1RMQsEPAkGJnMWaB3ycpe2aZLmItiLuS5kYTA7jFwar0DMxiLXf0i51F
UpS3IP3zsWVdTPw6/VbEyuIH6warSngGbx9ir0YfdlZU3ljNQnD3jOSLUAmbeK26dj2VaOZ3cDuG
DN+DnuHU66zZUaF6XMmW4EUNNpe9hN3pA4ARUZNnhLrAO3P+JTOENf6LaXkEWf0hNpvzh+KMtcNg
HHevxP//YBd66eh+st65KpHcxoPmJjxoxXFyib/1n214SVCg38btsV7WtSr2tKo7ZFWu3qFr66aC
G4Jsm2zWhwDBcrrUTEroQz4Npe0JH/Ke09BvY/uzmKP3EhUuYKWWrdcJbYCDtFhN1rLkTUrB0tGN
8mz8WE0T7b6oT2tNWn54VJ9t176aMX7icJEsTxOcTyomOwSg3b+FaDxC6aqmw2uGCW79uZbro2rQ
+Ug1wua1MVt9Kss75LD8Pln8TL/9SIrHBwkXVhTycoym4GZ/y5bymmg1HIUKnYVi6lLeGwgt6cF4
XXo1yTq1pXGwl4AAnxBmdKrISqIs0Ak6BbQrGVixGqHaDWlazpbp0D2zqqoAtBAd129hV5Pm7rJ2
QO5PGNJCY1pqFvxDwNUo9HEwQtNT8peNzsoMTFzYMpJ+6bQBABEAx225411bFkg8TEbrthAK1/M+
Z+NGw0OiXyHe5m3f5Kk2ZrfsDS6eXgSUJl2PET3qpAphchF2pC74JYHzTg/O5KH88SBu6IyuEV5C
ND/BtKl/yCheY1xdcVFq8XKi3h+GSjVnem/RtsxMEIrNqIcVcd0kjau+RUjdMZxIJ6Qn9dfFLjAt
aSEMeXUBYCzCmVr5RapcrfpQDvA9ucUL5UDkBTeeU1rPQloHPhDNpwFhUWWBDm60qIZr/evTew0M
pQhwzGQT60lLCC1FsubjnMq44CaNuEtdMP2PhjWmzr8L9pSCAj8vUrybNXjJ1RcRJxnov+ESMvcD
wjJVXxiQcvAGUAVkJ6lDX8bL1vpKGg9kFirtQclOZcdWJ2mmNdPUvU6uAx92JQcP4AhdWFJAxxnU
ZvrKgfRMKqcTL/MRthPegLAGlbJaqbCMaBIEB8MaMdhoByEiFewYJE8Hm2LZsd7qeeMhGMSSBVNq
PHXHYEvZ1GweAhs3riR6s8qHpvXYPauXeuH3FRdH/wkB2Ojw8p3Cg7wQ17Nn19h1pWMqEtVhkaQ5
KKH+fSl2VMhaindy0Zk/ahZ03nhJlhg7fqnhegegOUB4a1A4dQsKrZGWHnUH+GgJvwEQOLeS1f08
Fl0mtgALeEg9N/ryVuUp3At8pSoGermOw8fQLYPzXE7M2KUmxnvqebamjvblWt6KMcFKi82jOzVX
TSOiE1BhPRqMyx5oQlOEo+scvE1TDIDeBVjUvAFvvzV89r8g6OEnfkf6s18wzECbQTkQ8HfTMEJY
mbf6OyzKy6Ea2KP4rATE5GapiT667/HGUxcQG1RCKiP1ZRZiQ+wiCLSggXkMfsgpG7AEr19G+fko
gNrM9roROOzfNdyfVfhZngTl6KOwb1ro5jBnkZFfuVJUo5JLGs6QO0na0HynwxD6T4zeCUwGXJ5l
ct1BFesRgXnRDHaWTlc7nM7PPToixclhEMZl+KElSBJzMc/V7DgmOIdu/IHo3YLKGR1aHKrJN8i3
XeftYwLYH7yATdtO5TioojmaHNYV0pHMSf3LxfhcxDh46QQpx1SmiRB0iimU32QwBm/dLHxStF5t
WRJDoomLwwQ7ei5++VofBPwq45FP44XI7+lh8zMkAVUqsANk1Q+WoZLFD2I/PKIQWzSaR9QiChgn
hFyHH8qjnhDIBUDFAj0yIbk6cGaFE7bDM4YHd3xpbxaUFhdZB+VZBEu0mesD8/C1rIs0pgR6w5ye
H5x6MlRF4sM9lCIEPOVgIBVdRtbpco1O13FozutqmfnKritRUXv2+GJnJs/Xr6ypsX3lSAmj6CeC
HPyWYm2arf3fOKSVNP20m1MjudcC0Q3nCgOPhVNeSB57fVE+U51KxJsnRLghwVnvwgz/Z5130CTf
K7aYmYCYNxZSanhNirbuzvidMUvrCVjBMotYFYRHsnNdFyxZm7tGz3mqfVY6AEmoR9M4nCveDk6R
u85HWXCBhfHIsHmaNttKdufC87ybZ83GCMPOdSuFh1ky1DtKnPPs+B1DIaVc9BrkWSflGk5qK6dr
9lORbz2pPDNY7JSkIk1szH6bllwb2Fdv6MJJIC6LdtPDw70b7u+BH6EJ7l+Z3/XR1pnok9z1gPEK
WCwEquT3/EzkPEIQOBsLR2fmH7JJ2hfsjzhWsgoEG3D0Koo/leBReshksOLyf9ZuNQOZo/vnk/wA
Wq1BfgNdDvE0MgsMbnl+uXDERI0uggVlTbLteFqcnVtjId5p0maTx2w06hojZlQNsohkiFnvh1+Q
hGe+jUatKl9J0qINrsh6tSNAV3ysjx+sUT3YWunzUj8VuKL9him7mXHPaYmBt32J3Git1uMP4Aah
MpsfOIO313JxcNClXpmc104w7g9qenWeivKIA6y4FMI8zhjidVwYWmx4/bqXE3BZ6b1PP0PCzZF+
N5CwFPlwAquzMOKvuEjHyfrWjnVkPKd3J7W3kzYRkLwq9Acodb1VpImUXAQtYYCqQqg1wXZiEwx9
XxupS4qz16rq/fluL1OsUpx8tgpkmS4LsYreiNMIDXaFgXCzn29HVz7sJJbIG1fcIaf4vXkmdThX
lsD/U0MR0U9o5tNFIbiSqmgRYU7UJgcseNl1CbnFZvc9kW16+Bz7AzNlZ4tCS3IzgORbrXd1jzB+
3LesiXhm99WGELrsjheFo2j2imJIyMjffNpXuzzbUWavNEDJbn+1w/HCQLxM9nHeYi7uA48NkMAU
SmX1NgRoEpozG6amxrJ2QvsjZzXgrbAobvxHVzmLpxvL6dMJ7M75+SPrXQuK77W6OJV5p7rP9YOl
Xp6ZwfRf2+Jsb2bdCXvlGvEAIYk3d5vNkz2PcvSt+TTxWSYL5lQq1LfN24g5UtYcly5/yTN43bBp
8LA+ltdp0cC2ZLfBmAg3x1EmDD+YaZhPDqTCQBdi2rLvWt81RnSCiMCzJhLwM2Dt1Q/bmYW2BlsF
CppvTQR5im3JkFmUdkc1vUvcXZHQ2I0KFSFpHI61n1ckX9cjO64nrxSgXgbZvRIOVhn/7iTPNf9N
8gkCAIHdv8F1c0HIaLKH0A2KEz0y6Kq0xFbJFHZ2mWpfRkCxDcip7CZJlxJXOzfp9UMb6HzRsWWK
d+3GbG/qrla69zQm/WAxrskaopkP1IZD9wmhWNlojh1DdMfkR40U8mtwye9i3S2lz0DrWi8sKpxr
nDMECbi0Ou84nyPIXRtKzoMNatAE+EcCLX/FwQWDviC7z78Hzr4tk0f1yI6NLulNCHqEzELQanlj
iPls99eRUN3rkSiy6ABGCm9+fnTz7Dw34gDVsXL14nuZsPRoytPLZ03ybr5r/1LQ+6JJ05GbcQ/O
npWAajb1Y8r440GvjZBtRP2d9Nlr2yzC2bgq2WgYK9IRhgmAtDLaob8psf+s9sZcGYhR70CldMlG
L3K0IfNJMZ1gvExMVyT695DzHo40zCT8WcCiNdalb5Dl0lXuZLbu0N3hD6pSD2fVWBn07cgpW6Z6
2OltGIVKFnVk9Rm1QfIUS8svRSVPEX5MrQ70SzpuTVBZptVYz0faS8eRM4Fdo3jWYD4b3ip2hto6
Caxi0YegmAy+g0LSIxTdfDx7kxqDb43XEhGMqyvfB9ui8EPJJf2rowNXFAkQ3X+4lvR4/pUQOsBM
W1/ONpPPjPKijJNIwD3D6il61A9CigLg8LfIw0PjHiBhm0VKABjBbEapabiKQ/9bJUUdRjFIMwR0
QnV+5W07LMGA5w54jXjLLqJq/IiUycXc+UUEqrRYohN+xPGkvUEaNt0EChk6bF++aNfImDhGfhFd
Kz0+oEmozXCcmgVP22kCTGpXQo1007iK+HgY9sxgUYzihlpgLqvgJZf7aiBRn+L/VuUwr9RZavMl
5tYoBDGYm2AO5ALVmddQ+5tCf+I9k3bpUOvB4lMq0DejQu7104jQo5tedOIuNyiemkg2zcsaiNlm
nwKt9UNUPgpTOqgvKiSecKjmmrIRfiTNi+YDPAThZTZPV6UBkrmSfiLe/TpEkBrCmCCQ0Re3vVHC
uaQOyzXEwtlm0381aj6nLccsVALCWKgLkNPRwkLzecuxyX8FNFWI+qVa5aaywxsI1hEouvbI3//F
EkabTz5qZZeO07wK/e0mnvnwtD6OJpDFUEWGoWu/2TkjQPJnm/F99hM34gJq6nZTIiIxmrV1ke0e
vDv/f0CRm5jPS1RWorn24Ix3DL8fyuAScO2PDPzQ6S5l+aeU+C+ZSXk67bW1uKTYqLxzzeJJNCjH
hwhVsjxFUwvASUq6oTlP17dgaLZqhCnAIbhDlXms95p3a0vJrY3LeHI8S5IxYe8mgQrcGOHw5fUl
9FT0QFb6vwue/Qt3g/XIPZbhnsP+5NBUXPiYD0lGCHWom5Y5QFcYzmWsFMh6r7b0q21PulvBVGo6
48lHpA4CKztW0cRcPmk4ZwYpAzSFEWx/sSwnRmAApe2JV3TfvV1kwHvRj+VFvOwB3DF18IxwfG5b
GLRPdRzFnKoKRzSS05EeKMKebr+5w0U3raMvgjs5zVobkUowyqnzmKui7VMMBzFg4YsjMNfU31Fd
t/ui7PI3PXgIDZc9vDVy2z/CY1B94ZC4Kg1Sd6JB1Uc4c73Bxssl9RP46wRHLg82+5SVqn8I4fE+
lfdpbvN6qoodyHX5DUBvYuS0EJkwFb0dM6fQYqhUrM5ED9kyJYScxpcbTddM7t3Ikg2wuCvHiwKf
VMOmHMZ7YU9UlsqdWgaXcNPghYvfrcMWSImrL7Z+mmsl7t2fb0NYHWbDPuRCRMxfrpkq/B8UTrGK
cE8pVtJ2puCHHOQQzB/vRIT5oift0cfz8FlW2ssO65kdpUNs2OCqkVyeHihk19ybkN1ioe6NQTDH
/oEuE4BwKOadIlSwCQju2CKtC1aW9DYwJ1HzPAYsZzsS8qR8fDpcLLuo2lgBMwm3XBKD9JSdp5d3
Qub8E5XG5lO8Xk//j6gaabXWf/xYv+cq33GlrConJHcJZ9UmDhD+fUHLLu/xojyAjEHr7Du+NIoV
xKHWRqj4jKAS40eLctrGz+RP9y3+cPF0kgXZhSlb8nTw6YFKP9YaUTrvjaC5yBtnR2iZw2keO2B8
kwWv7GeOeT849Y9L5cT4hFLpe0WfGMKebKzpiHJ1v12EdoU+2LJTcV7XZ/fq5f/yRP04OJOs2wcI
JUu9Cc2VQiwPR18tBx1sQo/hMWXBDF2FegczSvpgQ7mUBDO4Q4XkoxF031DF5SjrZ9Xo06RxK4hN
kYJP7wVSn47CIPk5EEavXbQGnDn3gY3GY8LiMl13F3o+pDkVy+oB0wmGjxky6Olppyj0imAS35+X
UhI3dscS7QggOkvd2L5qgBRZeuyEdPbNUg2eK5kPVkMupbd7Fl9MYhHOyfSIih1QSgGCUAxFK8aj
DSNenyRPptUZm2o9BdIw6R4/9Kni3FMBr/HJFEG8plN6JtpmcKUHYOHnXiEqgCmIKkw1qjgebe2S
zRfTublgHXFr9GZOZIyHEHZhRUyQtGqbBwWCcmFFLxWlnvBaxf+m/sqAdjXIj2eWG73ANkge8I8F
dnmhLWPiB6Jo1uP1fiUXNenlYaMM/tUxohGXi3WTft269zRFSmcnknc4BWk4q6PTel4RXwhBYf6T
hamLPZnVJLbKOM4IK7hLyR6Qbrf76SZXJ11lmHMSlw5ctSlNTBbdPYPHbikEboMwI9NNh7RXuKTS
v1q1UsaApM+fCUWxbnQMpeOo/QWvM3cNmvWqIPl8B66qW7aWdDgFM4D+kfTu9RwxSm7crlMjuT4/
nTsy/mbVQ4jeMyLfHYH3ifC/0LIuMw5gRXxHN34iyRbVRKEMouzoZprW9xnemcC+WIgJXxdpTZEO
mBN+mW5m5h8MVYBHU/drbXvy/7a0nJ1YTccU2CbQxGa/aq2nSigQunSO5PZgeKGe2xDN4EHXcIz/
upfKkyJ9Dsc4WvI6KJ7lSy+9EVofLseA+3VlKRDbf9s+LgLRe91d9+KGyb5zrXCTfoBXYJ4A5GhS
MHYfL8YSClOrobzYQAm1CWwwkIkK+L+55hFRksEltZobOL7UBK51kYbN7ibTqi+vsmv6CM9stze+
8sYR4wsmYtCqoaEIFrIeIOIsWH9Miu9OmTIEDYS6KWYxuqZG4bb3iUE9+uw20+c+TAEju8x3FU8O
gbZgA7+3WkiyKN517LbThEraJnmmXBxQv3edIVYd6ktRNjo/f/XrZ6IheWIZgmg71VLgsOlrzSq0
5Q/CIIJOPpPe7dX6XOEOM6VcGGN5iLlk27pHhCzT+xhu9QEAB7tgJutXELHQMYNs1WFoJ9zWZ/nD
2DRQdZhwC0/SAIZwRBQld3T6Ac/Q217rVOHfTyQ7WakccTYPsL2rul1jH/cPfxrGD4fw2d4d1xt0
M/Gf1iPTAJtKTT5/ZtDx2WhiqBW4WGGNuEO3VVR7jTgmySiPzOiFK4/tSJ7AzvVQc8JY4zzG2NRr
U3v0X7udSw0Mv54k4zW/CrJhNL7E+McSf+WlpqotAkiMZ0zzsGakwfQmT1nj+3DapIP44ZPQnIuF
a7ha4oSHYwvPNArZuWEnu8WwykEWNqs9flgnbtVgy2gSUjcVDiva0Xmo6lIDdMwmVtGwK9B22KNf
NLhsY9TG/2ZZzkA1YXryT1Q2HZo2qODFi2sHZSaKmoea8UVw8l4Hvx5mGFDRUdB3C8B5SrmUCRxw
rpX2mRbnwfR5MVlweQh9VzL9TqP7zkNEyrgLUNJeQZ0jy5HHZKOKGX42j7KRpcdxyeuP4utxBSvw
i1cpPpfQgTxQ240hj8RuKtj52sThC2fXOfJKA1CbboGE8qZHYedORI+vvxblWtFMc5DcK6HgD7gw
tkCEQjCTiYqZqkOwCnJ34vGXkanDEgOyyPqsLPhx07tdYz9b3g7XnWUn3v6oegdGpQkyoBL3R8JG
aVadv6mpNnqirUOE8Fh1H0vTTLJzbeRgUi6mFTCHuaMCmyTeETHB4t38T8CW+l6uxAkwbdQiA6qZ
nQRJe+NgVYuOTTX4fqdlBNDgZ30sTkVbOI9JdTqMY7KdN0+jOO/NKcgeZoOoGCfv
`pragma protect end_protected
