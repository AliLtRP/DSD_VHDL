// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:01 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
e9oQdJiyqGvntBxI/dO3df0ftrSsuhE7oJ1xas7QfEvYlOEao3IETeejuY1d3uSO
mZTgUas32/AlIKI1fHBLaegP7hQ1iqiDW7Q4YEFb5Gd8jI5W2RT+35O+4OSX7cvH
eY+89g389gQvpTYfMJcQT/Q4JdJT6exTB6QmL+9Qv/8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57984)
oeBvR7fAkN9dmvpFaQJG7s6TcTA+5uopx1xvi6L6RSQ6voz87sFyPab1+9v1rIQ5
y9xBBEB76b7BYZYSmADF7PaQkBFEeylroqZAj28oXLaROX861DVybdY728qCNg8D
afp+MHBRi3gN5z1QYhc9YUXL8pX8YyndKvH2aMIyxSULXUAcUevjZfnfKeD8qNm5
rTs0Zy3WF5rGQdHjurdGgE+aBJIyLiG6jV77OR+EmzlDxOsckZWRUzZ61IH/zdJA
UXt1bDlYOUD989fQgsE9ZS8gvhaz/sdnoqIMCL3Kwd61+iwhLoN9Vk7xl38I1YBf
q1JjICwDdqT238zRdgbjo8gmb+SG7IeFe0hvAPX6Qd/Ju7pJWBwzjFWTmtiWerNK
B07L6BJJBHbMFf9BwDAVLsMvR6pH0zgEpaB2fXtutLC0PNCqsCUjJaZmhtUCTkNh
/wJvULqF9CYPPlP6HrEWjs83mQYvhMz4Awdu/wYeBaoYY+gZHWk9DmyHl3y/PRzS
3Hp85o29/mynulG7lG3T30O0T0MiR4KF8ojdyUbjYFExadYv4w7nR5qIoRVffXum
We/hUoGT+rRjv6zi7iFjSrL33HpBxlz0aVmgdF2ixoiF+wJGzROHcsVhfOezmF5c
wgqwl+eeFdI1Oal+B7644MGQlkRGMJvkpwNIpHVNFwyRzn2tEBYWduUN7pDUAp5X
H2VMKQAS0fNkCvmjLAFq2+y95uAWqGruNIDpqR8HnLiqDgsPCQIJZD9S045fAnYq
xIa6Eb0aUKiXRVZ+h9iFglwE6aqbXmW6XIo0dtPtnSCHRwe1hn506MxQkGiaSFk/
mf2d9pH0wKtIVH16jnkLh/nC7/C9hY7VkD8tS0WAC1bW0f1MMnlD0XU574ksLRlx
b55EPj5l2EFK6sI0kxaorCyQKlrpOEYa4gWeft727iU06qq6WvLZP23OhMOgKWQm
77uJjaPO4DocCP7UL6i5ySRKBUkH482eCRP5W6XaUFEvsy7tpfd//4ThSJ9KVLTB
s/LcDiabfR4RbxVoGwiZ7sgDwQIgeiQtHPPRIK1rjIlHqAF1JD331R1+dGA07QQn
dua/xauJhrDQaOUE9yc8LPJJDTdnn1sd772KXbTfMHP2zkVIAy3uEmLgUb6ay6cM
MZRPw9dQx7u/RYRKywqzycW+th+aZ/PvtkbCoCsoUUGk60HiFiZJR1UKZ+qP/B5B
L30oE0HA/Z6U4IKq5P0jI7Ed4WbOjUNra9fYbmYXly+b8/XBWOLOtkTpTyC+R40V
0my32jQ5DSvAwSMAxV+3ntQsoPNiTEQHc7svVEDrcCPR+BelWFci3Ppg+X4Rzt77
mBnGNM8ln+m/vRu7N08UGHXg6snlJ/VMx2dmYYNbku3hCnibAuHv9sBiRc/qz3hj
QrNO//HRKk5pJ0MQpdW5LeFu6eVcWZyOfd72Z/nLutStf/1m9qee4XPn4u1ka8aj
Ky+y4vOvtMYv9PgHwJxHzh2YHW5LPdEo0kdBmx8VTBVbDe4NolVpeO8urzzjrx1c
r7NIiVkYfy70UIXOx2iy45PZ15jGT0s7pRYXSJW4WUFUFx3cXMRdwfwYQ5iKsQ6X
wB1arsQQNCC213oSjNc4j1qiQ63EzuOnxOUWkgNi+UfB83jiQFi4difBMGh3WcXH
V/dCI3EtQBSI5OYv3y2Efn8ac4wghLjtCZPXkfsbQ9WIPy2+aDDmMZ2jRfXZVfr4
BYghcEX4i9Oq7Qnq3i9irgcUS7lXK7Fn5cV9oTNmeRpnfWci+IcvDvMQr88HrGWY
r6od3CCrQZmTwttRsXhRn/ATPBL32+0mytcOpwScORPbQ2o25Zj1b5AyLe8YdWCd
mgrLst9hBEwACkjQSsus+bj/RIbI6uc/brHELzUDUn2uO77G+Z0s1hkLhX6LOsqc
fEBFFhRgydNEFX6ola8rM60H+X89HayYKZkbol8WV8enBQBo9P+Z19Fn/zo9wfjz
xdlyti0seH65BQtdeIjfaJmMXhjLeaizzw4zNy9XGCGemzYm9taOWw2BoywUwFi3
/TknmAEp9TDaVJHsBUxwtgv/1V0rmF//36i5MsdHAHL3AbaRmndDQ9jWy+Kl8k/i
uPw/dRvysnnbCg9d5O7kdqbyHlf8IatcPVCThplM47ypBHzRsCqcEODUsBgl9syj
giZTpFpjgBB/vI9MlK3BpGWqf3oGJVHIBZoHZ9LSDG6RNbU9AYBP177M2z068qAb
WLh4BQEjAGo43BF3G7JnBc5lvdg5bbXp04SDRaPVecnxL/w+toMBgr1rm8JL7enk
zamyxc1DtTgeGqAOZqnxXtzR3WGdSEhwUM3Fa9DN3WBXhV4U8P9Qja68NnrjM09o
lK8bKvEKXtbKofupMsyjrxQQqlyLAiffz7d+1yqGINIRP5xDBSF2hVzrrYGrx4u7
SdgZLGfaoLvFtULOrZ8E4Pjqq0rFcSNeqOb85P/oZ7Bt1WxEfGg5jnn2mncg3J4a
DDdZqpqfES7aOB4UJ7a3kVg2MmzaDKKBgTDCa9+iHrF9Mj25zSQWWYLftBQtj1b6
kFIhihB/Sby82p+qKjQrxbGHsarAN0kJfgdUAzqRerWjX2sKhcpVzyhIy9koWpsj
TDNeZGUcLEUHtXZErnsVVLmHKRFMt/n4XLYqhFwksOjsfQF9pFoydTxvr+7PAivI
vM16ATtSyKx2E4UEECmIk95A0j68gWBfuW5vsuiXfPNC36VZXTDV+zot9+SH4s/O
/O6l6uBXuGLFhL2o9kIPckDZCtCJOSkEgjJI9BRuFwFHJH5+Y0jZ+LTt3+cpMCTi
gsMma4/SRd4kAAcGCXdUQSHydLqzcQ4lfOthH1Od7FXKk1Q1iG0CB4HMqhovTRFF
mz56K/D+IxV7VWQF4NRO+XUuMdfDLYEDKcNjx6fuMFxkCGaWPhIxwC12YUQH8yS4
Nj1eiZ/hitb1tVpUMZo9I9I6n2yohbMXV8vKDmsjISTFOS1CcSqNY9I5hnwGbOxM
rpSgWLLYI+szMyZs8YlHbk2QC96LMVEF6W5XvnGnE3CJNCbRrNktLJZExHngAIPV
Y7jbZeYlVg2Bk3weMgLiSuO2ZGlzOGsYK1zMWdOT5AWzr9x3sgFQVOtRg9S6SslV
iZFx/cSqWmU4ukjbm7gg65NTAHz5iURxawqxgzezLrvVKByOvEGzl15wed6wiZXQ
VClBfcXGQuA66JZ6K7w+ruvm+Ok4LVamq45m/YKUjPp8u0/yX5RSxXnxG5s21/pE
DsNCTwdX30InLTqC0xWaXqORyAnln2W1VnI9kyMuUc8H9HYVMtxoYUkrY/aMvb7i
lMyJKnjqjrQ9ZpjBRvOu4WjuFGJoA753tCTx7yWn8CTxaNoPZ4Wov2Ja4uv3g8eD
SlzzCEIaxIZr1R+d9jNWm8C+dYfT6OFxfQVLfgpxrSPSvcFx0RGuVPdhxyImhb+I
bEpaJKuLRDjBzlyA3Ajxm38eEL/LPqe9/wqTMuM3NRRSESw2qPe6bMkO64L4NtC4
aXScCxnhVXztrcV3hW8p5EJ1CYcIutM+wzjtRewVn/fHG5BoL/9lxIBfslNqP2UV
ugJ9/UB+12m0mgVhnO6MTG/JdQMpdWcdswUZ1DJ6kqHTw98VYZJJycplbJa9iz14
hcM/HJbXZXitDW2XpRX9NRv5uf9nlE58MGm08KB5Ur42YP0O4CK9eyDG28gT3qko
eQwu/AT10AcAliYZs4H+QU2mar1l1IOO8TV4ig4GoCAb3GpinEoaX4y3qzsEQmxw
h/SiBFX70JCfrMeO25IlRITF7AE1hK90iCsppdRqVGdNol1Ul4BsyssKIVka96B+
MPVQJAJYc2NjDi5/my/xljY+7ibCEgHIdV8gJbnHtRwcthWgZwLspAPmZX23uRK4
9WLe/jtjuVDG7e8GFAqeUnY/z8onfVPgXSsNvT1ZRyNugwSV+0gyM2DsFM3MCUiS
/bZFOlFahdVbp1iJTxmTSYd7Bq4cEMWKzkm/hMTGciAZo7P/x4CzorDDXLvMI2uu
M1xcR/d4jnXWO79vangHqpz+vGZ+zY+heGUT4SIFQ04wFmk9IseZ3x4DQW3BCMoQ
/yts6QzM7bmYgFdQh0Ru/qFCkngFsko0RXmUDlRkQ/MORmu+CaXjB7EnbCGwMJtT
8iRIan71gojcAtgZz67ZRYmrTXcaMKQVQVhbF+v3OfMmlXl1YYUakIUfs5czWM4a
SM8XEv3/xhokO9qX4ZPm8SbOES/myEws9Vi6UBkTTbT5RxreBX8gTw4KM5NlXWW/
p7tGLTnHlqCWpFVqDEYgKIjpvcaU5WrVFs6xoskIJOJCStpsSIhzMexKMGikLmLW
rV55Ed0gv2xzG+OlJD9w/+o+Po1o0/d7B5Ln/nO8ouWtXvaI/NPH/kdyNjJktaVi
C4G3/AMyG0InG4do9725cDNUnUCAx67tpG/70+zcGZ0QUcjzTT77cpeWQEuEmAZZ
UByZk5mlaUCKilP31yWIiNuSygpv+doB0FY9MXKHsDAbBJ9+oxVOtH6thsDtVSFM
v7VaNaekcuKHost/JS8W+gPrWomkstIOjP/tW8Jk/7tCYqK4G9ytcAk8odqR43ss
l5jFq6VSXNvJWZ84pumnUOagl2zSjOxU1moI3/5WlewIdk8OnqEf0fAxCzzNkKD1
0HMr9LJFZ9w1BjUEPZzdT41/JmCgJYv5JFyI++jwzWLnce17NNL7/ks32Zx3hoU0
ZJEcoQyVaHGNJlpmVQCF33BJZQvvr830yvhQFiswRRPPLA4+L0QX+mv/OZJDC3k1
gRQL+aHC8z075LgAHgAnyT9DB+2/TgeMJ2MkQXWmOpyx1+B2wbhvKJVb1CW/a5sG
kENbj2BCdO1jEi2bKSsnz59hhnW0aLPntjqIAuzZ5tdQvZr621h8p2VnZPxPm7Lj
BIJKBkFAVuYUromDHrm4nti1M1wQzCrNfXZeQVfwPZWM/oBkroUUwoU0hqNHs1B/
PbAQSQb5oJBeTF/5iklwPiE0Gl2KSYRfU6LoIBn3LyxWwXmYyB9yYMylFaMH2ZQl
wIF8WywjfYq4i9TCLEFOl9jVFW+MV6ThlS9qR8SgI4DYUvhwv875exKNLbQGDmoH
c3bLQeIoyOQpfpf4YS+kUrk2kBgFBl5xHJv0/C4/sp0m61PUQ2q5Yi8iqCOt+W+D
fSMzYgdFuXBcniiObkUuGGNk1RsgeB5UljBorQI5v7X9cMDWWJ7jQnS10ZM0/djp
Vl1w58svYbBwmwmgOTo/FWgblSs4shbReBB8qRt1Y++qa6QijwWx6Z1CRA3yZ+zZ
SJP6WJPEkt48ZGoEMxzjEgi8fqPIvUCs2pk9sjZ8gx25l/e13HuSXVpXj6ic645a
JdMHxR+IWSC+er0awA90UPZHpUCiFoFqYYcidPYZ9eOFFB54e4sUEcO2TqnVZim0
tgMxetjvCPskIMOhd707Tv2hZ93SYbz0zVkEyQexpAxIqwCoBpgrWaeeo+aRfHRV
OUNmjuq8jqhEZgdHEJgtBEsGvOBp4dZfiTBNmCZ6gC+J9ZWByIxsjmxmTAutmckz
hT6PdZ2WhgV+QZVZ7XlPfyBYPkygGvZBe8Rj1ubZiCIjFZNUS3Jwnz50lX/+uzy4
pERV671u9p4G8IEpR89G3o3A9O+3tb7170oZoTWrW/cbMx1gVoSQRDaD8ijrUMvO
RpySPHk9ueTUAsnHSg7JS52RmazVnROLXqjO+Hx1cNIFl+G7qpGiL0KeATjPh7+T
lv4hvSdXSBNGs26DcXOhHPO52wgyojVpE7v+RmD4lVd72mm3+8I8Met0aOUln5MV
4n4jUjmyeLkl3WGS+GNeTwdXm1aXCrH5RQl85+w7K9ktIcIjCNPFWL/+4+3Ne0gF
nvPWs0nkXw3bovRbLBz1nPCD7Atvftm7k+Kfe2uby5v1dw0pZsQt/6JniZWI71Qb
GXjQ0ywlOpLideRq/HkRIURVFaDqVQVulJq2Z19eZ+s4u7x78HVDLUDmznh7zf1z
WFGuCWnvgqylSJYUFnahb4YMyacLSiLEFeyvps02jhbI2vBQX9ObdwaGnQu9ffNq
gmO6kqV8ltUjcob7c33D4MsJpiJcHT8ua3H7wjJFuK80TT1M6SeUsD0utykn4n0a
39WQ7pG8Tkoqzz3pAaXn2D3Nclm1N7Cl699vBrtNFmPQRiLKrW+iF4TFPPdZ86Sx
IHz3lBJNMswGxeNgd5iugDZ9qdjHTccEDKWaaVnZVKjdpPS3a110oPW3ef6vRt+8
FcB6JfR96VbMEyfksKZflNW23GPXX5FKTdwC9J3hX8t+//45KSCS2Y4/PlghPKE3
GoDlOSq4dLS7bZAc/dTHNwURwzZUepBTzajfxYfOBnmZNv4HeHhHeFuonJ57LSnH
OJKYNjUwgM9dMgfBwTDPVncvfxeQEZUsvyXoq6uz7YY3zVWgLy5KWFgAgaANkRbc
xJz6iSLgHQjAg7aYpta57I0c5hvQCVJ3dUI1JL3d+H5TGKiD7+h8sd2uny+/QSzk
XPk26bWRH5nCeXajgcVKLEXNo1meqWvFR3tM3SsNS5UCnBWNm6ZaSkv+vZLEH4TW
HvpYh2fo8LT/c7C4yVffAU9NNilnG8A97vYCvp7ifz6cHpKkKZDum+u0IwMGmqah
q+ULJhE1RZA6O9BJurE3u2YyQk1jMVn8fCAeXzOn6NyAS+fWyMc8jhbiixY7vLR7
+xJDncX2HWbEScWUarXKILhV6sl81jXP1XsYz4f7gSgoQBpPid2gdfs088iRTzmc
mo9lmT9t0PhY64HiMKitcWgRFaIxDAH0ew+fboO4uc8NA3o9DhYQp9dgywUnq6/K
1o1oqxgx9lwU9Nc5i243yJwlFBbYhJpELy9rFbfQgsPbAevK5Y2nMDlf4L6rdOdY
Y1PjNyRZM2X0rB8JBJVOegeqOi5Sj/yVmw+KuI9lIBoLol+E/BNzMXhGYtPpQxZC
X5A8ehtSENLlNfNQF0v7dC2p7aDXTm0jEWNv8nrnsWFGj2dGMoSjB3og3OuguxOm
C8/hilD5rTL5uIc2pp4lg7kSkeKIHpvgm/dkDh3p/pe7U2eGEAj7unTLUmv3V6P7
dzydEXmAT1rA3FE77QJwU1yVqHyg5zpUjOv3N7FoBGJqj9PD8FJl8OmMxGhWLW7E
N4yfUwS0fG0HpwzZTv5boxohyJpOf9Y2LJ2xHuyKmKCLO0QkT9eXhG69UTAaEtvt
GzL55MPk7EZg93ooKGtariM7XgjKa5DmOS99dLx8AWVahS16Q3wcSRoR2hvej1+K
iGvpVGXKjGp5i3QZE39zD3nkjy7qp8RvHQoo/pdGErqNWRaZ4oTHn/j9UF2zEHzY
LdYeQDvYdRzFT3gyHEDtwUMzWe4iKe+JOigsZUo5/GCH5N/HiIHuCGSX4OwKXrPh
8eWECh75nsxqsshMXVgpes1JMOioQvJUVFDQ82iaRIl59zkhBvHm4qyztV6J+B0P
6dfeEnW7Do91FFrr/0sHTUNrZE2IwUDXrzoECYyZyB3SsL8v7iEuNfH9iA+xfyVp
ZvBtWapOru/YSzOJZk6aO1g/PV2iZ3o7s40A+DDbuZjiBw2J9TFqh25JIEQLhHqV
+9mShzsaxOWO9dd1f/+UFEF2fjoyb/5yij/gCezwy5A3zN95HvZjXuIrSBvoDMZt
YpkcvveE9ONTNHJ4Rbx8efBIfH6BzoUkXq5wBB6SqkyiUkYfWBs8raFz0Y57K7fa
7rEZn8EjmgYLD/wMgBPR1QcPt65b6lxu05v5R7KwOX3PfB+1fcrFMQFPTLBt3k6/
nPgGhNcQ6VOAvq1F93M5xf1X2RpDyMD70BMlpsNdGk0pyej9VGr3o7orND7g0sKB
pLTGZ+f5p0wG1O0Z5TgK45TMg+g15fOBkuDkHmO9QO9B+SB274U/Begk01ulHCte
D7GZL5P5NIHQdFLS7rL7FwhZ8yVb8SCvOErs1TJDdoToAPwPtpiGipc3L4xiHP/5
My241UWm9/W4wAnWZnP2KGamm3EbfkmdY4v1jeZHknnmzqcDChzhCpm++GvQ+BJ1
tQSvDwrHl5AJP3f1XgFtXoOxg5xYGKepyo57QltB4/ukq94xjvEsUUVkIg5pY8qI
eq8965vLBoU5LbUE1O/wtKtetiwjPHzydqdOjAEmZXeUNIftvglMMC7DZQcNHWbu
RntOEXY1EycTOcDuzFtbwWwvJslU1rkIJdZk4XQT+jqikRbjetganmuIyUKKMbb8
9x7ULNR+5RUQrwEUUam/9yA0YOIztwYoc9bAKHI/N09clVQoqhjYdMse/YdLBjjr
HSvWHvnisY4kXR1a0jq9cJ8Ta51pNZjBwsKKaMTsyNSvYYqKLHMQ/Hp9Zby7M3ui
aAcIiDjqmt1ukz12bOIHij0OnWVMO/+mDqHDEMou0Mxran7xSmU2zLhmWZoTuD+A
G53IxqWQkPrq+jSPqT/knlj9o8FNPp/Dpg5DIvMOquCLhb/61If+bDGHNDLXe5+c
JMcgj/Sh7TqoLau2zxlMKH3BOg7bUXYHzkgy07QzEjhymDNwEesBwTpZgPIY8L/W
NdBqABh3ls1gn+cFsW53Wgib7XjmDChq6o6DQx2iJdDsO30ydZW9jOhwKc2YK0zx
rsrwZE68I55wgkWJsKo2PtkB6ErPhTFxtM+tEHlOtvNg1PV0r2F0/cUt2wiBUCPq
Eulc/dFiVLVyZHb57jXzL+Wjjg++4Cd4a0W9rxDmGvvueOf+yOGoat2QL5a2pxBS
We1TkKjr3n9EuE7QcjiAj8oFDJpOEAzTHZZrdoUs+uOmccsrBsnHTl27uGbM2CUE
MOd4Txg0UBN3u19jJumibLvyI3oXCEWe/Yd1oVBPdDl4VNVW/ku67q6v2d3+dmSs
C15RNjtNq1hFH1/mi64nfR+5kSvZd1/bgagG58AOT1wKaS9hMjYzngmK2GaAy8Qj
8vur9tXI+8mI1N0RUldxxgNmNx11qgsh9ck3m7eValFqi/nY9//JFJoOfzon74FR
8+i80l7fVOYfX1TXPJXZ1P+6Cnptk2rRS2SrzUuQ0F2cxUgjZJ/fe17GPziNmABM
yun9EP61M8hyHYFdrVJ148Kp3D00oFa+oADYRR9PnQpP0Ivu400L57DQXe63vDO1
7a3Z9wyAM5orGa2OZiGmHJGxnc7976rTob7FAU2Jzg5Yc+8ycm8iDn8nI0uOaPXf
sSOtcf8/mgYh8d+JzclRi+bpioigE/Ze+GfGQAM5uiVFUQhRVLW6FHD/ptUhCZOh
21gP7PFpbHkYkpTBGDNWUxDhuS/NbTRvkWRT+7TAyxCFooXam3rAAJm1OTGO4Fk+
agR+WpTHxfd4iCTpnYckFk1CJ4D4jYqQp3Ux7RfiNd2KdPQOtPilrEFDpsBOkHjh
iCsF1DDpSckD/8xk45m9ND5X1MouzHL60rYFmA3AStp1Zr8SRvzO97IHvci58ZQg
2Hcaly0qMDuPVpxL12U2TsvdQ/B83N3Y5RNtJXyzciSE/U2UhYAGkQAJXhKI5mJe
zu8N4uckqryRGOoT/cuwbcX5N6Ywsuu5iBDL6I+ThN4oY3KW5JuP6tH5HOcZLLm8
UL47p+YfSEXoGVHM3gxj2/J3bjWX75PUQRAdWnw2l04c0Tc9GFJM+bPydIXTzkRw
w5al6v8hKFO1ggkxqGRHyDeVQtAMV2jI7VrBfEeMDTDb8ETj8aDIqltb2UVrKZgX
wXLRhnQAZaeC5IlAkqj5q5OspmVtBMmp6iUQB6SWw9e3btbwOs2UleoaRwIpQ3LM
RPerZvcHobSWnNutROZwQ2oj/Fadlx8e2qAUggSv2FuYGshjeVJfLdkUkyqrEsGB
khtDQgEQw4tE3Hhh/DKooRgrsb8BwPtmEVD7i2tFA1gKIFITm3mfXtSYsdC2otxR
7EXvWvToh5P8s8y+JxQ9pD3DxHPl5BxdQcPrSpvredzzQNb7xr4xtkx6pJ9ZThdq
NDQdEInrBNZAviGeAtjH7jBUc4BM5GXwma4UhJarLLx7tSY4Qf4iEVauWZXOJG5m
xTE61t70x1+HY6URRay5sCbRBelGd/wsdf9LgiaTzD4d1fHcUask1ZbQoJw/vVUi
UiFVQ8zFK5Pxjv7KkiIOqhaRVG5LLjzP5xVuHhAJB94hS14jRWeGtRkf7I6PTyJX
1cAtGSzTRGUAsOO9U7cXR9q6DRx2tQJ05czOU9ZadMyY9ImHg9MsOcYhelfDr1H2
yjLI5wDRkmUvlFPRRL8qMmVZwHx9P//GGTfPOCNdsYE7hHo3nr87DP1AsGsmFxL2
ixBIHgJqAp2JyN5GFWewIhZLI4FhdPg5Gxcd6aLiRXiOacxBNctr0+6t3WoR6WpB
34GlODPSdoJTLeCV/+GKpdoDdPfsWrLvNfKsmms+6ZwZbVz/6MSPsq9NOAIurjGo
VloIDGri1HKVIRYKP00D3zjU3/rnhcAR4x0CFRcporUOZNKONUz5P57QlO7latau
EMFJNvKoVHyu/QpGq+/5ppHYJyCAqIheHBuqkySmFXQHomhKlPu77LSa3D7qpYRP
bkVZkBkYTm3nZTn1xvp713O12mfExDHsgSFk+QjQrBvCdhpJe5deiOiQKQug0xPC
mBOcBfyBCdGVgvPRWDHVA238sDuR/g7Hy0A6R4rdisEpE1Hnxq4/G4CSxfOi09xH
rC3xXBEeX9Xx4Xw7RTeT5gehyVwKUV7woZXZLeccVM3pmAsKxniNSDtuOh/fQTLa
m6YNtRVI7mViaoMUjYB6JMJXVYD9OslA7KYKjH3Sp3texsC+u6hU3gLMgVaMU0W1
TS0Q2zChqCRW9ylCM6adxHPde7xpeFdy2fsH3WiSRvtHark+YNIz21rMYS+Aab4N
obC2QZAJemjf53cI3IXzb4ixVPVaclqs04IKNUEDUcQXJaa37Arr6HGGO2tvYTPy
649Emhu2GdjH4OmImL+Q7amAHwwwKgfpafw34UBAF2WX5eMmTYWK/ytkAhEAOnV2
V4gGOedQKV+CZqWrE0YeoV29N3H2VwKhYJMfRTdRwMyhxcnY0o/Hie0w3BI7dlJU
PXtzHhg1bFa5B785rdcufWVXcjPMa3Vi7S1VvWIqMZclkOIEYbIJ4t2SdIEcsZ3D
8dcY66UNSFp2INJCkIPMLVai36zjgMNxnkHcs4YYaYUSkTKRRM2w8vQixzEriaMZ
7qzLkA5hy/jaHN0hd9n5iGcDmpG1mvL8kszGODM7rkejfupgUKLm9jn3fcmEiAcx
WhIQ8QsPiN/e09b1hdOoTAZuQ4PjUVT88OJ0ybQJoUT5uIGZr07FBT1WsXFDCZZT
hNjW+BGK8v+ZO1J7DIVrwyNHExT8UaeCPeAAChkXyxD6hgRkuXC7lY98LgTMSDvC
5KGcWG3cUNATvzW8/uBA0qixvcQ1485zWQneGmSn0QuophJObUArfA3bjsneb824
hqWVBH9bK9jMh+qmPpNThaNLW3QuMiREM5xfvYNbItrOeahP1vEbrO+OrYhhCsVg
lF4cou4sSi+w3b9QrFi7H1g9xMJRTep9urRic+E1hx9RqWlEiT/tGO/BfVpGqO1i
u8O65yOs72j1ZuhKv9xYhUjlViIit4pEWs99bBcpdeTEeXsX6Ctot7Y/l7DFMKuy
Bi6hEQ82EAc3mNw6M3ID7H1sV2XmWoKLKLdOc19sPmBp2e4k5bh5BE/1lXw85YxC
G2FF6V549kmcyTgbPlfei/rYmW5qcQWisK8P63DB5GNBmGTEQiDPT+Gyy0bvCiNy
7FAlWs+9uCXnlze5pb+uw4B5OwI2sXv84jLHZuvFyu8FIr+L3jxeqrdIoi0YQ5kR
PCkRHoVr+95Uicwm4JNJamjHoXjWqDUVe/+nUXMHXtDBntqfLI9+i64Dsrtluzsp
vRPDgsJ8eDy5SJCMdM/yYutoR7FX4uL5Zk7KgR2TNeciKZYvIG3GxNMDtl2HE56N
sfK4D1f2bqHGOQeQHwOm7HDzwXkXzNPfkcfJu05cOqyno+Bm9drfbx6Ejr4VN3uk
X+btvM/Wh2cbYLr0ZvWSg5pJmlDQicoYOdmovzR2H7KoR7Td+FXPHVVPjt7zIrLx
ekvBTaQL4Ty++Rv2GP5lCD2bcLcG33J6HuPf2+2pmyU3BuPvNfpzTHA2aHtLt7v2
Ya+QMxHFkVNjP6mS0DDOTx5U0WIRWYkqToDcWFgIJUKR/dhwE0IJVw8+Kqai/2eP
1ZJDPgFqpu+Ag/rTI+k7Fljz8m0jwM4en9iIhQV8d34TD52/Dy99QQdguMmShV4S
pO2EF8GecSSCMGXJJMTjxfCmfZEYuNBFrmNvXptBpUcKeREuqwUSeuXc6KQNunm7
1fgAsZFU75QL2fglDGyOemvPFQWVif5l2RHlFykmsV4q5aVaaYxeo/eiUh/QCL73
ToRhkZ0KXvKnXCSeHsC8gMNWVuQczz33ygzlL3kKpEdYiQ6UVWfEqUHowS/ffY26
gSP/anDyf15W1pnGrHg7awRKtFvrBXg+pDKVwgWo6DIio7uHYy3fYXZz8YqqBnNE
XaS0+MWsUkaPLyhV4K/jFpeJ87BzVzlzpiEoPUXlZ/WY8iqy90nD+Ul2KGaWALl6
3OjYhFZ3M7PQxUC9Xs/MuZMA75t9fSN2cfJJnSMy9Pd+MY8hWj5E8jDnhx1JEYvk
rYChTF1blHRSBZQwxzHjHquTNh/xRiH/0FV+M4aP9u5W2xhyoG9897ni4J/Uts0A
yazXJwIQFqdTdKlM5trErNSjRQR6ty3N57HUHRNBmMZIUmHeDcx0bNAxADOjsss2
snuj1wHp0tfaSn9MdXbLOHnFdu7273u200EfZNSST+S8MbbvN+k7vQ2JvdfxSCnE
u+nMmCCHgDyKVohXB8gKue1XZbzw1v73JFzBH3JFTDo98HfTvJXfU2/kFtMmdrkD
kkMi2ehQpnwz+WqJAfJOBIGyQ8gcRX2iC2Z91eKWX3F70oDgVS3VSB3hWIKnfGvY
DqLdlDR1Y4iRGtsq8w74EeokmCtJtNqkKr5mvPaZCTtIGqe0xuFivVGcgcHkSEhu
lKhmkjD9OXFL62cJvbiDMrmaTkRO3dY7tCwUFnnU93BdQ9yt+/HqsdU5TAbia62Y
A3RdjZw30SzKblktiuloH2VEdkuxNJH+AxSZK+L6UI39EVB5QlSxWUGNpuX2N81E
7RF9XL25eHUeqZG+PHLJw9QSTBFGqp4teh4mWyRCMcmg9GYsOcSjnutVc65Rcomx
z5aXRo/zAkYh7joVx15MHy4hfnRKfJht9Cty6Uj8ChNrXS1jpAGxblB6KoXeZSL3
MGmymfHhZXmPBglGEF6bvnDOcY/E3zM5wg/wRa9TfwcpcWee4e1cPDWHPMthuB9S
TyCKosyH5t9JRT2iShLBzvW84f6bi5jEBcvAR5ugHgIMLqlyMQ3sNCTP0mwaCeU3
FJ2Rh/IjQ5G3HaLYgfkBRSDO/QkRnoGDC28WOA3ZIf/JCoUbNRP4uSknMWsT1Zfd
NdnLyNxvbCE3L0ScF8Rkq/LT1L+46jEPehuj00ceKyJfaTfwUkeOeFVmQdrRN67D
BT4k4KpRsgWewjEXxHvJJrG6wqS1ijpDn2FkBIqCA1KGvEdo6zbIR8Zgc5vTRhFf
8mflTfmoJ3O9LEMsULgHLV+BUoCILCuXsx9qsQLgDskN/5GD2VQUNzIvGrIA1f+b
KlWIUHc5CUsRANBRA7wvTf6E/2UoxoLUuiC2z5+by4v6hC9/9+5zLCqOueD0Ee7Y
0a4G228Pe19c9rbroppfjPeBfG6gETJ/qjRzHh5kRYOyaRd9QVmkk+Zq+zg9kuNi
p/r4c5sU3eob1yP9C20SUR1hohDrFQr4F+aj445hvT/UjykPLNFGzAwFqEN8uhpn
G78lh6gIWG/VSKKfiuAJvzWr0hp+wJttynwH9Bx/O3KqqtMfgk1nMkj6rjJAuBl2
0ewvXDGr6VbTruG5hysx4AQ3eEYEIPDhPfkAuC+b4LO9d/trHfNiBVXzSL+JDcUV
B0wlIcgSB4XhVQuptxaTLE2k0MO1mWvlEGhj/E/HdLVZJZm+2gCD4df1ObFhuuCT
ZqfPbZWC4MYSEp/lPRSm50wp66HhdTWHGfcMgkAHNBcVdMlyDq3gEpWqXYn/VkUn
GsL0PFGJopGGicp4rw8l87jVJn9ARe5QVAPFI6fGB7p+TLciJUPM2uh7hUKiCD7s
edXSCkH4hDjZQeMu78tBmnc9K33x+fDI923oEjqGDhOwIexpMpW0AIbc5MoZbPdT
/Q+wPS61uvqw+0jnMqrdc/wk1TGza0q6NdfIPbjhCqmIGUxlxaNoYHfmbEvj7Yqi
CZJjqAdDAj7GeLzbHIYQd9pRwU98Esl2fgq5TWOuhlR+ORCWLVKPnQKPcoDb6XZN
XherTwJeSchj8kAG2hFIudPxPc0PxXZYvkU6zXFmgSaC/nIsnShUgm7Rg5aGqSup
+z3UNcvXfEM2XV0EmM/CI+o9+qutT3ETuSN7gIEQLL5aPdzY586JkGaJqO/2/uqm
KFIyWl1vyWRm8LENqVfzv622JWEP1z/R8n2wsKLwDVQE+Dvtsds9KE9KbYgxOyOe
w2mzEK65KDS1daWzHcK37Zmq6OzGUlePYD0BGdB/RF9f5U33P/6lVit8NZkMLEDk
WntNVK3rE6Rc+oFd0TqZjmMx6Y86o4ba0Q9lO0XdVajt2JMTX4/+VkDULDINbuX9
iE0aw1k0tDikQ620aubYiiBI8h9sjAqeyXzkOAtUtn6FsbNyjI5cCMO/Fyvg61Pq
W3gjMcrz667oXG+4F57b/3CbZ4YA5X5GRdnnufARtJFiw3/C3chcFSCngDkWoano
NssHkiBhjyKN69P7rgvh6QEVRQ3LGpqLmJ0bzcmPmE1jk353CiwE2zE2t0tZMyKn
OI882V7c8KWNxiyrRybMzYBXWR0EtgMCDzSnEooaRwM6vxsvf+UXzEWrzB3/sEGh
CeTljD4CbcBxGBd6q+1yHFCM6vhfVCIjA90mfkhPYtZ2cE/YaFIJ+iQJ6uBxJBg1
jJuQvcqiJHmWDwK93jDbq3i8AXcDt5w3LkRfuUR5j/c94VM2SXcUchl8aDpL062f
1f1aTJWVHkDP+ZL/e8xZ/WiASBCqxW+BC28UIsL08o8PdC1jJvGJjzVPuDuZm9+/
Vd1CAYztMUdXlMzAc/9Kg1lFzyjBRj/hgYGIg2jRWPbjbKgniqHRub3iiA4ON07w
TKgtH30b9IwmBf1qrg3dMG1d6O/DKi7+zYUfoEidJrBP5kIqOymAH5aBOK4+QT84
PE/vix3iNw3O0zsNNoPQ3Ylvig/OMlPd7KtgcUHuzJz1013DErlNHjTKGo0sSLdT
eXI/oJOrmjjcc5D2bxVv9C8T3js3CI0SyAjoJZnuQPUz0KtSSCpXt3t279f0Ejyb
DJUv5q8fCKrRVCMH9vYS9nv0M5ZL03MNSBursOzU1W60mCNSgInM4kwA1p7l8LzK
zIz4IBrqjY3bQC1awSPhfriiNfqeTEjV0OFyarJrsWvjyn+SjK86BjTTu8D/etdw
CmbDu5QyKnqe1SZZwAVDHaNa8/B+SdOBCrIGsLqcSE9+8jHTW4MNNQ5KuC/Q0p3A
HgtS5hQ5D2zaFRd6W9c8bJSED79HIUAFfPo0HifFiHflu+jiPPO+YOEHZZ+zMJ6w
4Nl/BApBMpDj335E80i2BEXTwjdGnh5FIX+GfuYMA1RzIB8GLkWxxaMrjkMa6Hlb
4U583w+Bx9dQ87hPqLtXF678H0PayvilifLV/woIM1gWnmUE4AV/T3KgC3G72gTm
ID6CeX0xQdNKIJGFEquGFOEscOwW5rieCySDmCIwY49vRp8DrqVI2fDDfop8b5T2
jMSzvS2ZUjqADFqOZVUG/YJ3R6Cf5g0TFVVx+oZY+aMpfZL5RMFiFVX+Xngfaa7Q
qVZgDRBh0nyCytIXJnhNgo9tIlNPPK0IUx2cYyHRiC9jcPsk76alGCHSWWH9xcEr
nrRIks5bSSaxaRZkHVhLWk6WR+GaC2dguzQOR8ZAMc2ZGwKtd7/aDHZvDvue9mdo
vaE5I/ROR79i5WJbJ+pPYcMcBZQX4WwfX7AZ2LBH5tbHedTlCa656UO/f4o0GSRO
EDLZsL83Dq2SlxnPBVr1gTiYQdJYYZiV8ffRo1XhilgrSlUABBNvvHk0pQ0tL2rg
6OLh8QrLZkT3GbTAGKuxeVnW93INS6b/i2d3L8LctzADDZGwyZWiZ1Mc62HkndH9
Yhk8PY+RQrMo1bYRZzNYVIB/D8uxWUFpTXS3gkApAtza/BbTva78BywrnlPCoXBE
cak/PvARxQ1xEGXyAx7mIVYOfG1F+uIGpB506A+0311XjbHnqVthX6qc+w7jYKlu
9WMce2ngd0H+A4e+W+kbacGGmxGLUzuYQAWYt8kTgtL4iHfhWp/S0raRDAlF3AsQ
C4n1aCYm76tqQ4VY9Ltp7q6rPzq0h9JxdhukUbhtiAFLv9DWN63RAKqsoKFONDP7
4IZIPFmtFJb3SPIzou8ixRt4rDCwBIidlSUzjwEad+MYY8+ySjvXkMHLlzrS/1RX
unhQ2hnjq3EQXHHXCIH+OR8oJhJPjBnV8Ky9MKaNbVK3FHBLpfcTmLb8wZujnIC2
/egCFYIRC4Np+fv8zRP6OmRrPVIAlqZ9PjIRtYWmT6IQ6nZmIbVCiwbHcVcyVUdh
Dp3HrsYhfOGLTyKM5sux144hFj+St57Ph1FaB+45soFNB86/72SFla/kzJfBdBVF
KLxklA5dLq3j2zkVUBERXhBwkejYgKRkd53uqaypSfFKBi81bzHLY1BidBP9pHkH
PggEOSKjydSIFbuLoIyTdixNA6AdnoxFCr7MIAdNM+6tgUdv6u5KcsRK+aVyTwBO
4qAn3GzDpnuugRizdnXbgubw8+lFvaDsdtNclhA+pm+l8nyM397JVz+MjneYqd9P
Oj+JHUcHQQca+SupYiPsu8AHGnYjIcnRAX2Lw/PlvO9qguA+lztZoRIRthAi5FEm
8RMVWcR7GXfoqpFXtCC3Nt6How0Es0PTexGxBlBY3ntXt+Wh0HxHpdE2F7QO91MI
GKLAKo5P4UvfXxhSsWx+ZcCB3zk2libXp8+f9OKaiXxnjUoxIunb/jgksD//fUC0
XfdqypAf79Gmzm6il9PSh1D3Qtn+V3EeuycN1whjF9UiHI/OiPoV/CW5wdXNWy+Y
gepISnqylIXnYUgRNuDizQpGXOh0zM3DPRDbYw+o2P0vIKw2e0zykaTjvkUIJ+B2
6zAgGZWdftTn7ime5q9540+KfmxWAXOnNb3+6F6yN1dE2Zf0KOpBo7/MWK77IXT3
JBwF3mhcVnBdhQZKKLtkxmTbK9xnBSxAPAgyhYnAqmNNK8fvoF54MaBg7A7oXF6U
+LZxBCeShWALx0j2YGiqYpwDbjI9ZkJG6rZ3OC4GbKuoTsa7aQdf8AhPI+AxnnK1
FYz5FbE3ywX2BkyI2BZd5t76YIwd5X1bQTRo9grRWdgqF/nyHOQzof4zm4D5ladq
sm9SKSMHUficpBWpUFVTwTEwtxf7j3xE3WcWLlH+XBeDkeYfuLJDCPZ4TbMW36K1
Gxtx1B4cO2QK0iXAHMN2WZq07+ZpVzE8JSgSyyQ5N/Q0XaqdNt8JDy8v9MFTsenQ
ujEFLZBDBFgkIk57otFSJH5Bk2QVYIgpDKfepXbFM7sLpyE6wLjOndgsYo66IDmg
QI8e7zxO0dEk509jBuj8zr0XzTKatpzqeRNAYYebrouGhUJ7iptLHpZFZ6WshZ7h
eBP99+IxRu/MQV2Fbn49I/ItXs8yxMWtGTa9aSWkUIt0hztnlVdQl6rot8g2++Lo
7WysbVE0YjSebWkHGbe/lFUlTmhbrhztsonyLZpqoSGiRzTmyAuBiGkUssum31dx
aTKhXtX4E+o2oHALYUEpeVaKhW/cAVcvdg9Y9duXFPvGlEZBE7lHW7xFgOaw1eK+
QA6bU42sZePQXLsybuuopPBLWbPp6WG6HtT/3B7XzWakOrdsD+yZkF5s8vvFg20g
Iz17EAXHhi2X9sRlIbMnVFwHEbpYaP7Iex4fd13OrP5vRb+Nb3v0kSH74msIS39I
S1MQP8RDZH6G6dN3lROf8TG1JaMMmf4MLZV21kTT1PeIpfGOLrp5Zjhy1Q6qTOiR
5+BsHBn5OmzDsGYw9GFMy0SHWYPjFexYGoC90PjG6VVWDgDiV2zF4UH5W5BjbP5e
0SbWT+2W6Fxrhprv2hslpi0/N263d7d5tn55UQnAwfk2QlH1RnGWeK5gdtjVNMA6
GJaKkv6qUCzuUyJzQYsvVSM0h+5B9vAk9jyl8PUVvA+1AIwx+5V/kI6WJXN6Pdtn
+22rRzULdOYOXU5V1EGKSYyovrdEiU1CaGqDbQJkeTTS4LCs6dZtMzFiECukLXdL
dPOYv5JmwFY2NELTfwWVXWKp4gx69kJTTbQRQNLdjrrUbeFAXgtJT0/LLUjA2b7w
bvYrGZ7Iz5aSTr+6LfwdfEgj2cc9MBy8digN8bnC5Ge2Cmr+/30fEgicqGtOkXNa
xhpyP5iue9J+CGQ/BOJbXs1XQ2h9yIUEmKkYUWdf/IyKSpq1CknulhzhtactFLWe
jQsVNMcu+kp8OOIIiS9EN5MksYzGyaZ/DP1vCwOLMEFAhrlwDJ7aIFo1e2JKGv52
JtxmHDi/SIyuHI5U/CMFaK+ormdvqWrQJU4Jcu6VncDjxHNkwZ+RX7VlBPXM/P2m
xwAE8KKj3zv6YELXnrSQa/IfH1EhtP+AvHR0DtslQep53WEo9P0z0rWBJ59OrwUi
Isd/GNER1/CQ8FfHzOgA6hpZT9tNfGLALPP8BlxOZjPUbFz/bPAz6bPXT+YFTNtS
hJ0doaLAhDo5DUuwV+5xCUbENyxfRGHNHWdFkxSC/au0H4WthPuEv0Tmw5wF5X4P
Xrwg6M90pKIIi6VRfzHp/iLcBmGfNVZ2+zHhUYgy2JBszxUwQCoG3bEL638GnkRu
zNwS2o5t0HgCxHP+STXIJ0Zgw6Fa6jDFOVcLBclPjCL6aYa32ND/6hIBEcy94vkU
Mgo4XnIwoVHwSUUDg2i/6eH6CQ984iofOP0ffB+WdGHkBaSMRE3prFM6Z8Txd6l1
IkLmE2zos7hC11v0az6bISxdw0dNaeZHVORkry8zMvEKcfhTTYr2m95MhoIfE5KJ
SyEGyJuTRzNdSpzyk4i5OzOEyMK7OFsP8Hd4qsDBbt/+BmEziA2vPc+1ovmve5c2
a2q4b/IfXLn/cIx9/Yb7ZaEkR3x+OoEMuA6elgxkFAYozk2dxCL1K6reGQiqCjdU
N3aD2QYoKDDiZrG2bL1XvDwThyiUc0hztPCk1sKUy/RbayldH+IIECklIIp9qZe7
WQbCVDIfjMFFSKyg7OxWl2Gq8gXoFAo6uzS9GHlzRLrVkw0k/c6GaufJe3xrVK3Y
6yWup+ZYt1BvWajIKiMQqileG2XhfnGq53HBLbrZkfBgZWUwxs5SbfTMd9tZgo+E
6pKdwU/8vue82taMQ/LsWRaz0t+BqTvWENHjgkKdKV/gxwyXXxRFMiU8EKw0Q+xp
UPwn9zYL1ffn+kwfEVEU142T8ROxfO8sRMaUbo2iXGWlrTTFLIsvpH+OVfEgL4/R
za3J0OYCmA4YKcBahVknfpHdw5ydXhd9CkmJrbOnrQNTzvWWNLkC6z9vWwrpkpka
fSlm7tnl7Yj/SVVw93h/qwKiy9E22uAmNfiEm8JsxGM4lF4uLFQXzdX60qG+7K4/
VAofRmoYDoTzxHSnReKS8AQkC4/cVqwdqnNUOkbuSP9cjqTIFtKBNgphI1V6tb9X
1wNhRaSlh/QvuKp8vbimey84apDOa67JPnW3Ddou5DqWk9qYoTr8WTpLwiayUn+k
ab0IwjQnwnvmRIsYhcQ0Qv/rJhAezQ4/sWgIVhMGu4OA0aYcsW/1EM4ZUtyPLgFp
Z6FHmw5P8hsl6Bxq6jcajLmsA3nJ/lBJKpl65pJCzjF7xgwVnw4OqEEtCJcz3d6K
AD9f8KhE3Di6Axgew2JvJWkKUc3NFt2DsCzPbFSrlRBEGZgNzY32o9BY8xXtcMDy
zVS8Cl6le9ZzGUCAX7ahn1SoyYC5WomnyEmx2JN2ENlbTNLLruDl0mlu4S+eWLuP
dfHVWdHzjY6QFBaE6A352Gtfq4mKzq5Qn+Yz0o57Eg9oHSDY6FHmttKYSZg12mQW
TFyxKdrHQKM26lG7G8JqCcXfiGwjhfXIaQTjloEshvE/2+MBnu2tBnwamHYsjfRa
fdMjvWuZCy/vItM+iBI275vwL3m2wCP9CwxvYdeoP5OPG0+djhTAiKu6c6dUHUW2
eZ7LCnH7sS4caDDzUA5vXK5KoBzqTNDn0JGjJQ2Nl44WKid83e/Pzo7QlrPS/npp
rAux8IkEsb0/LbRFXTrW7o5y/++8F9w0knC43tw72DbV29k1uIPZaGMde/WrXvPQ
nFjaF1Aqc8dHWw7+sbRzMz5saGbjQ9BnshDu8pXTyIQ6KRuhkWm0/kUq/RTmivFN
Z9qx6ZSAg0xzxXPIqUz12dw6Sz0LjoSbHvgDpgU+zGa1khNQpUcNYCI2ZJzZthQ2
0+HXRaNNDUGsj8D7YoLZKzRQBZWQTMdBc7J0abi/iwVuP7m8pgsHHVjdJ/hVhakv
woTImUiZ5dwEa3frI+RtlN8e5ZrNewWTF+x7QqrKPCPDvMYIiHOY4o9srZkpZKEb
IPaBrX2MCfY0rnvg6w1cyVVQFv9FnWQ8Nwd5UUpVdOQyAwVwt/74no1uBB0qKpGV
1ezNmdn4qFxnWVeQdFxms59r2wYHiBEKv2m3Db/mGKmXoe4NKz4eTd1nPF5/KDeC
hZsqP4roOZPvk9Kfcloj7KIP5Cn6IovRHyT6NKIyjK1rz4LDgxmaYOKVmOrbxNfE
Tf2jPBsBzMkxYs30d9rpQ6hddKmrDwuA0FIpsJsLUVCFw0KdCJh1v8IIkjtUP8il
cpk+rGvjHD9oRwcWP2lMkypAV0yfX53mQq3KvPDPIOGTvTALGDNnptq8z04RaoGc
Yx71lD3sZvGD/VIQ3UGWB6rTRcloQT1uMVaLtiMeaADVhgNfz9gbQBpwUe3Nfyc1
xI33wRc7FckMJgU6KlM1lPXy5+EI7FqE0Er2ItLO/zpB0eaR4CufnDKAs2JIv7Vu
gl42aO3xMnbH7bbDu8nlABjJWrpnfGadCRVZaAVCwdtCEzRy7g5eVDr+YJiS0mo7
ApcmyXHz8LSFOdQ5yWWQhaOyL2SNS/90G97xkSshtoWOWLXTTF1m4P9eVbx5wKfg
VZ/xgmxmtGTFDY4QneKqB5QmE9QBoLMJjvepAe5mHbNQo05a11geq5rJwfetLOt4
tujLWH4+QOVySXJEN2wBNV7jjWcdxuoZuwkFfAU02K5czGEaNz89XL7SDrmtSBIw
OUgSlMM4kMXnyAagjCCv84KEBftpKkx5uSGMqwzPy7+hmafxEB3+8GOTWde+OI9T
I8G0TB879Cmie55II6h3WzHy4iHb611jpvrl+3SxCrzqVhXYz6mddIxn3emCfBWi
A7uYK47jqn4DZOnIXGmueboTzK7meBq8ZClCz1zbjlsidwoDsG537Sr2qfLmFtJP
e1bcoSFpOLGV5mwJTHamb/abAgwY1WVtx4YSpFo52t+6DgaF7/7aLVcxD02r0RUn
5P9i3ylmmlWu0pcNwv9yZAor49bmnIW5tpEZxqbU98qaZ58vQ0Ggq8Jugl0B+YfY
/bSYe0syqGk7UZc5fpOpSzZXhQL4QcgffcZablZ5gNa8JO0LiSbCEW6PVcrG5Lsj
rb9odbU65IzPj5eH+5uOozcUhJPLKQbksADCiVATz7yPy9cNxVctEUNlLwWaP8c5
/q79uMzOCAKYLz36XduxGX+zZr4QOdWFHyOz79ueJ6IRQkYgGd/2+JB2quezOMQV
7fv339BgiajTBdYXxKpL/YYyJUI6FscmzYt5RNwuNu5PEyNOGM682GOrtpX5iWrg
7crTK1mbTUQM292wLIppUB6iMJgI8qYbmqagR+HH9TFCFv1x/aDigeYqHc7tgdhy
bRTuhk1/frFwuIMKhUNR2vDBj0dAvxd/49MrUmADBhHGwJMOG+b9H2eNmWivEthW
tqtWfMAP0CYJWOMUs7s3fpzBJOYz1a3mDDxv2I8vzvD022J6gxqwoyqejy8ZjCFy
ran51gvUH3pgpFM9OktJvRLZ3GwITEj7DR/XasH3LylcChKrN7Q/A99kjlNYfKDG
KiaIn1c2FNFbty9T1kPaMEEZq2LRj76T2j1cHs9UDFnwxUZLS/mlv8KuASH4VgHe
oP7bL/43u6jCQYJr5rXF9oZ/bxgJO9ob3px9ypveUINj6MQqHszDI0peLzuh8WI/
5UhvjSoN7jSGcGiIIiO3cc8Sop6njwaRoYi2ym4P4dt2XM7rqzC+SPMAM3EIVdYo
N49zXy/NWVlwwrbHz07LlEdD6Ty5blWLyizKVSpvm/k08sFWpSc1Fx92yAAhW46Q
eQsRo/4hNjmLTeVKQoKXZDir2SAOPc5J68qANFhSAFZMvcR130iiuGpzdfW/tgsB
2gJ3lGHxqKwivojo4ozIkzPrf9zpwoLIZpjhWln8hFehJjjtugS1fmUsPkAChWOs
7pyBgAVeNk2EnX2olwH1raOg0So8uTXiNTqM4dVabYoMi7uQoHRtTXoCOYapQs/Z
bH1c2cI5WooEOEHZ11YMo4wmKO9tzd9Yuwk/8sR6H8wqh0arQPM6RSnYZZZgT7G/
3DWgqv0+/lzBqJ6+OhvSOsm46kijRd7VM0T//XLO9kFtNE3ZFH1GGIwerWX/NP+v
MUbsjesToj8dq0E0AY6yjaZX70C/T+lPk0Vk6Sn03sl0C857sxTQwybV92pyw76N
DyUxiXppMU5RN5ecAXaaxtLufTxVYUz3f7ye7RfsOFArE6gQO5V9GEvr4quDW/Q6
A9c9rJWGzRAjdzVrNpbmsOLx7iwLmoyCSiNYrakoVWxv/BbboVNweIg3sLCujzrJ
+tIAkL6V9RCtMfLa+azwetAXduf92dK/JyBkyesS1ccsLQIQ3ntRQli2j9RU1I6B
FNqY1v2JTUbzno5PRSxMxxe2skl+bXChdWEp+kNJH5mMHuL4hZDz49KG36biayO+
JPdeQAtZc+YYLj8Jc71KEeSRKCTpZC6NRIc+VrvF/iQeOfAX7DZhXouJvfaaSLN7
AkSuop42jfI8w4gMxNRztffbQMb+vzZg8yhD1CGt3JGXenALb+SjN26mh5nQAO9i
pT4yf9jReG9jb7qp28JsmyyNgMXo1fivNO+aZehPgyvId9yZCz3AgaYC9jw/fl8d
WoVTgtZe939vAUlQE4hrN6jLq/R19AkkD54V5PI/5v929xR7kLa6HVVwPB3oBG6p
1zmIfLIVyXulwF49OfEL/eEq9UPgCbkzkJUerxWT4hI/ZlCQ74lNgx6R6ULgC3+z
e+cuuUzMgFOA1RlVkacCCYykEMqsLG6lyyFL1U+spqsW6IBthCpdJUpETfiyc+6n
Iyd661uxpEDbXv+TSmGhpSVKgGI6TblDwboatbO9dMmdjs5yuDsO8F0P84RqonzZ
bSFrlzr0tdL0/xLsIUF6vWebyCgHSF1H1YokBffY8kVZGdHSxZjE8ZVtOyWncaTr
uO6y/r4xXXOYNDPKi5x/bPUjvxiZzsi5AEJfIRZLnI8JN/exWLT3JOP6jpnW+hOk
J6sT605Ll7RawiAoA1B+LvYoMHN2Ejs3Bl/IL9UIgv5PdhX4UchmSVy2kJLRArJZ
cVgmppxg8LWmGKXV/rBjEsBmZmfMa65jzoPtatY2ZAsSt2Ji0wr5jkhD/3Wj1RFv
5CUIXSt+z4glQAujnNAmXgkhd5KmgX/ZOrmPW0npJhgUQqCUsPVP9jf5vnAyRegu
n9cS3sFSf5LC2Z8G2isT1mroXnyK0+uHZS+Zr9FMnLAnIgS7B/ohJ/F+Um10cGQ6
sHPIpDgrMdfFCzMbfV1O/yYXKI8e8habFOwIv+0bM3z0k3jTYEMxEuIKBuGgrMEk
j6eheVveOZJFw4Qz2XFbzvAyUtyVqmkf8a6RrdeiIkfV/VTOcqZA6PBUopfHHTzT
0ToOxCv5l7o8aCAU+ye1F3Q0ETcIU5VI2KA2lJccsTZIUVcxod+EITobtuoW7Vtn
7Ba6n5DjQwSi/PGt/iIb+0/tMW61TzB++fKFGNeN5Z9m3oHqDcJsaWUIqePQfWPQ
3B8/oyXFP3eP0OflDxqsNZraxgDwIk8zQMKQyqD+/ks19K+yP28vp2hUFMB3zKiK
kVA8TDt5EVw2jej9XrHzFgeE669HUnl8mJFDoDRSFpBistbPyhhCrDnanW5ueN+H
z8nCVLotuXKCFms5zpEoKZRhrwcjNvN2RSPmdBMj4jf43+XaQWwQ+6lhc66NzhUH
bZjzxiugPDnVE3/cJBZa4fFjWYlkws6ODPLWbR9r871+We/6rUu6vrTVBL6E0ce7
2u+9D4xBvcGtNYKlVUS2wJSQN48bBz5dBNhDdc5mgyeGGJpTDFnDDEaPbi7yBKfd
mTK4QyjJyn3FyRdOsWvbvjA3hmLTqWgNLKfqbtmLJjm0WuefLT6GBVa62YXbFOYO
pL+jPcWnKadnE4EVihWp71TT/Ub59ATHlxVmSBbGQrkYxnQhQmU9gGrYel1UScDO
0b2hxmhA8PGMFJGAVMuoIKlDTvkzi6xb9AiIsFGZ8WJsHxpR6COrt6n1BKXvqa/b
n4KTfcYutVQo5RqtbuLnaEhzRx0EgK07Pzbi1f+krH3vBge9tuRqeTsboRQMwftR
BUTedPylnwPL2ZizMyxpQO1ZQknXJxXnlEhM3r6K0d6txSk9mbazfpM/3k1B1Lay
E38kq/pJpBHLt/QerrS0SxHoLqw3RDKFDiTOfwGad1Ac1JZ+v2YNaFi/gHbhTZpI
FuU3P/OyM4kptb6z3DfVXl8M+HGSb2fU4ULztJgSOgn2UQlEaaPu83vLWR7MCf6c
iDLsfjNfpeQpXGlnwuPgAhUx0+ROdmfongR4FbjS9xFfW8W8hx5tfKHCvx+dPOOq
1yef7/MRSp8E5zTAGDvos5ZCYc+lURK3fEpWFYN/yi7sGjfnLqiAeKvu2hUfTIuu
6YQw8UTL5f0pPFEqmaHB/QscK/oX0WQAVirR9lyWHtaAs7kZba0lricQSx51PR6X
QI50EziLw4sQCek6Saw39A/xu9+ZDQIlKqY8wqXpS7UkFalvEGZmHN58bv5Xla0a
lP+26wfYIVrP6A7JHqKlY9QxM7uVBz4CWwS5ayyuoSNLwgnolkiMsgapJdnbHD5P
DeDyapv1nwbV4l033cJBj3HdNW6DAhdf3kEJCp3oHbdhxFEImAhGsC0Eym1Kbg1I
X4dCtbaWqsYAcFLnLIxlUhyZdSDqJwRVnBAvROnWe1gAOnANhuqNr3VjKdguFgHh
jR0yME+VCtSoyiNpMBCbQ6zrBUnYFRv9QQjJFmZ+7hYK+pFUpxbZRdTqo6Ce+SQp
jehowHGVmijV44RuyjyZm/CmIfdnADcG9PokBdGg0Xin+69fZHIvB0j3/GXbnUPY
cnQTc9IXPpXmicnz9ycquJZRWGRhWWeK15C8taFa+zs7V+cFxADQcfIRa+2s+ycQ
E+of0cU2zDYaWVI/hmPGPY9U+vzW3334+MpOwhMCSu7/tUZNQGd6vnzZHbdlXo2A
o8tCh+BFC8Fr755i+9Xwh7ZU34DmZb+eWSiC9j6ogr01z1JnEc6YQf+557zwbPok
R8/n3d8OX2krebIHHTCBxFpBJzwopfCpl2GVfkUfPPSyahWAnz1Qbta9Yba5K8qT
2lPsk9FnuaXSyX3V3PcYh2I8TXkvEBAnoKs7mK1RFEs5UVUeDb/NW/OzuZ4aGUqw
CZ8wMr8l3PRpK7Goe7OWiswaEZ7o7Pnm6mJLSG8ydyQ/GKX5mxpl9OSOUcP+H7cP
Mq1QKhEZLGS/wU/Ipny7jxU9PduKe5890QjYL5Q1r2qI37qB38gy8jLHBYmpO0Cq
XUwaiYa9uLiEFVq4SOTaUrx9jwcoQw5AhtsdS9byyV1Xlj6IUSs+bzdlDNywN7LS
DGnJrFnnJVFIMex/Ic9Ako2w4Gc2RPezAMMjXATzIMCMLDwNIrhTpGEw7goYN6Jz
yybe4/wXONn8rf7JTy8p3lYOCF9vBMEFEQIq3xLCAx8p3ZjEOonrlRM8CYujKOwx
doeQEUuLGXK5gOUZ8xl+IhvkNStk6Vg/RUjh42zymn1Pv0pfkOM62v9HbuwQ0sCC
/FhqhD1ZGxss7qjhiNdbXczLYQby1zBt9pXn2qs4ALxhOk3IH09cRq+WEoy2E38t
WneAyomX+oq9cdsstJ2Z/TUoCmnjw1gLiWZLU8h1OvOtH8Mpj1KLYIyW9WoOOuiR
AkfGwUc4y3fmz3dOTGxcwCZ+AUXDsvFwylKGCxdCuOIRp++MhygxWNZp6PCsz/sx
/m9ycqkUEwgawIjBGUkF07eX9DTcSP3+ItQRxI0zTm0i1Px6zN4znRSD+V4lPwEH
cFxrd+SoreQo34HxuoIv8tQNQqmNgbD7MDRngcFXrZjuN/9OH1i5mi6O4QwEINgM
VsNrYDWlhJT7iGDTlvluptq6wVBySy+6FVYu+VfsxK0RCOd3DGkUi7U3OVeDPwS8
O5OWKTbCgd5yADR1uOqj9ri9LmSMwTjhifIrAzmTM4Hb00i0BwH/sUtVhvfpuRZv
h/aeAkC5UXKCBih6x0FbSo1u5u+cM+50dcCpXpwom030SXshyuIIUIvVAv0mpX+5
H7IH3tT523uXbEmej1rjsLy57H9cC7L6jEAigyeRjeSwlUUbxmsm09swnoxyzAE6
sBLdslUtDiRomUQOxLB6EGP8AG3WjSshsPuGlzRHb9dG4tcmwzbqvqnb2jiq45Va
Awg2q8gXxbqt4NOI7sFwbboN98tcqxhyeEdEohc/nbTk33W2XCUfO5NPIoWnBM0M
DjwuRYZn8XvjDXikKqHX9Ff9qmKRNI16lXj4Jt3EwUhLnRWDV6xREGjLJCS1U0ya
ia0d9EBu8eV8xFT9Kg60YRF5YsGsJ9+iU7ewr5ERTDfYfx+LEADkS+d5ZXbMEyIL
EOHZcgKBUhlBiGfpVwBotiGbKZ0pbn0F0AxxI5S9PLhsJXJ4i3WXZaBsoVICB/+6
HPm3a84hQYyC4D/HxxNy7MwYlf+awr9kbmIJD/SWdg5EmXesIqZhoeO80AEIarfP
H94unF0TyUZ8QsvZ8igD2jbaDrIrt8DFrvjuzhfU4shfk9Ww5Id2gKzQAdJS1172
zII09e8GkIUqIdr4k2dxesjbZ4qmt00t4tqoHQDt3vqseUsknOhY9q5nOgbWCqYu
r4g+aFrRM92fbS5G9lKiTvNfn1CsOrxq6TioajQJ7rT0op3b/cDpp9IaOoGoEfy9
EqWvAYaFK7/ACPGE5d2nrCCf5j+ABcTbKbbUiESyNIOxP7Zzu2YNOQrmAb3jbAKP
VGGIN7fJ9GVli4xkLZM8OGHYl7VkHxW96bEOrADgQ9rxA+Cgqt/MrtywSU3a59dr
mth9ptjjcxZV+cET7liiCedrWvtr1XLw9xSzr5vuRe3YcluOSWXZxUnCH3DrOcf3
hosfVxzwS7Hvt8rsGnqJoAxwulBTmErQYaVPAFhhYl7X5fCTmguEX+HxUNsePjT4
wukLZ1xELrLCkox5redMp/SzKh38MJ0N+yE7KY73dT4+tDlhBt7I8whbCVuReyuW
q+/UM7QVy1c2o70cyoMhCssMuzCSgO1zVttYMzX2ic0U9sgQ1trFlWsQKdDgUeut
9PhqFoChYAfKRmJDFIdC+vPQwBg/0HgSjRf7psOTphuGqUAESBmNZNqvJG0Mw/9I
vij82K3q8uruRJC3Q1xR/vzRmMBZkVfzD3RFq5sQ0qwQBZ1GR2kgV+oeKw9iMfqH
8heGgW8yGkvn7fTMaArWcQl9SE21d0LvKpMiWCpH7chuEkto1QEBcJhfPmnTaIDk
F952VkAmntcDcI2lSwdrQ7YBhiMuXeRTs/3niqKW7J3nPvIhaJ6BdZSih5xHGgsn
NRfi4Lkg6BG9gIqKNUEylgXL0qjDe5kq3Lq8PEZetRbitz1CKCztLQoWDt8bL2Xo
3cBseY2RUHFiWdg0SQjACJ3C6kx+qO8gL6Yxreh/yQ0VohU4xxoQw+fZt13mCjCZ
EpKoQvAdxPHUJ0fy1GRskIK8h6d/+tu5vFvJK6Ik1mgF6AmwPXAWPN5WwhmUm1Rs
30ORtae1PQ4GyFKVta3o95ZbpodyJB21shRhstLaCj2HNhdE825+gm2qVG9VmUw4
BT6sYOvpT5q5KjnYqQ/AKsK/zrPZHotGvXeNkptPOlBWQpE9U9Ofki7Ly9/BlOqR
9HJXPzapNTHWweJvrRlqQeSEk3lFajQNxcZ+tFW8g1vv9Ka9ortx4duFk0NVkLKT
DYVHkfZ8yF7RnA9mBzbyT2u9eysXQaoyQPM9b6xGsHi0J+sNtt5FpmYaLw6Tsf7W
y7CVr3MpP4T/NCGztIYvUsb5pPiJdRFZPwx0BXEAy/XHhUcM+ckV5VAR/sOAFJUP
wcTTp7Y+zZx4lGMx151dyXK5l9ynvSrARjE+qoEwlk4uKN00Od+5I9Eyt9jR1GTf
7HC15Qo+8SDxLtHjVnbCcsXRl5WgQQUY3NsvkKgo5O7Fs0dSmy7Vary7MdinaAXP
qH4KiLS/YKm7CyajGAxak3cIS0pY6+Q3UrzNh0RPTuBulzlxZ5NhSo8wrlMdWsOs
RJdE9aZp70AwLLBzTDE+jv19scDW0Kr8mESQiVCGCRUilez41PBtqOfFcBg7jgnk
nS6s5mszN1M6XCCJRUkkdUXwI8jiXmF1uCNTRgWercvRsu28pt++pufuWQHp9lAq
fM7sJTgc706CUKZ0hiMZamJW00ORYXyhUCBGwe+0dud5+tJYoSN1g15IGXYbmCFk
1zOKZ/2rOGpmQYlxtsbupbLrNSdfpTFsG/eUwW9MdLZrLNOj/sbeVceLdmrHnvri
utihT2o5pXWrYyfLL7dYDXu6R4i777TtdcDDECD40EHlKeT6+OHJze159Z39XuMM
NiWKAYHggRZJWhbxvUm9dk7aTYQaMkRzMj8FMpKsTZVBNz//sVZ5pO96BYlezmbl
BA0PDP1j28jxugs7QJ1W9xHg+RkuQc6v7mWX0CSDJw61uDSNgP2T7jLcmV22Zp5p
yL8FbJLGSt2T2LXA3+tuxBCGECZ1suApHTCsR28w+aYz89Qv5kCqlzc66HsBuKZE
CXW9AGFsb+b7rDj25DaC72yooPx0cYiyTRyuJGoX21q+/xX1+RtWXJ5tfLP/V6P1
04OQd0IIuI3OWpL5oFZiaJPZ4xDwVl88OJdlHCTfBfCelF3IgV80VqLpRZ0PVDqm
0SlYe1YL6+5qbIv8F85vdZ3A+qLUNYUcg8HnjAtKC/86oFseoeuvWFGdwR19pTCg
EHHAS4KC/Wv0Y0myS67aJSsvQhCeb9rwwqpWSHaT5LhdYfFMZiD1bK4DnB0nv/PU
pElCAeXKve85GD2BvHaosTFoa/PKGpBMt3/LunO8NNro6n5VnfxskPKsT4ztd4TU
fkUU4TaRCIA4Vu0l40IQ0lwZ7idoh2jj/0dy9r02GKIX2VBLk6aXLRu+z7LhU9DQ
5A3oNKLX1owB7Lh0qxc0/L0hb3hkb2KLp7INw+qDkR4bNha6yIuh+TdpYddRuemS
IxaSxp5aj4/nAJp/mW9/FuM8yNJFGFyETDV+12bpvwvIS5nWysDfyuaiILgpJvo6
rsgG+bxtNitS4aDjYsByLREUCjTixXlqR69U/bkI9CqCL+0r7yBXliyiSWjPj646
LVTHyWlaOl102GX1JSFG+DAI6dmuHJL7LcuvganZXWiwWBkGfbCItM5oEVwAQn7D
9P7ehRBM4TZ2Lo4Jo9Ke8q1c8l7px84TEx+ThrfV0mJ4D6qTodyntYv30B6mz4lu
RycOppTSPmha/+rLEtnVt69J4wCjgjDOrHX6VQg0Y4uq20P37ThCmh5/UVKkpZTN
baDA6ZsV55XJUpIHki8XQYYAKPPjc1CqIOKuINBIPcFCT4IvMhQjBaaoOTac+9Fy
oKwQQICfUG3tyITIdoBQrZYfUCO0SVx+LiZIfPUZeanftn36w1z4T2FJXDlkIgRp
3QnlwKb66goAuDyealZqZYuuRtqRK4UmAiMInihkWWEEKuadI63VkXaAD5fxbzFy
RseeGi8sZ/QZn55e/J/gmhvNVRdbZqi4piaMgD9iyM/+ns8J2gUYuX69vQinTNcF
9hQew8TC7fvjprzSnO3DrnXsflSYUbyIuXefhqlHArYdTRxuyqdtJT4wqxy806Et
gz2B0Zvosmi/zYSziUu7y1r8B7p/ea8M8tKLWMIOvAYnuO7vArOEF6zfwvySrlNS
j2SFmBd3PYZ8rkeICGf70yv/p3UCYkNBfBbU9yaIRkkQfWV9hoBQxKC71Si2ghWR
sba6QlS7+ouc8fnPbdp0Cx3ulF2zwb0pQ8Xa5YmTBhrSjFw3qYQi2sSH86QfMThE
VeXGT5UN7bsoX4F/f5+/NXR1OibCVrFyxCsADSFL4ZeLVG8BHxQjLWvXiIFyaqFm
ZKmYJaJd13BgShKXwdFKcHJR/dWiPv0BlkZD/SLQCmhZNEqXvlMpQHMauUDQOL8g
275TYrVqSDGsJ63wlWHCqvPqJ5KtziTutWFQzs/nUH/yERdPwXACOKYmkozpV3oi
3X9dKWPXHGmwK5U1urZS0DiIzX5DUkTYtr4Z/KiFZJPEutNZA4iJC5DIoCCoK4zO
9bWa6glekN05RduqqaZ3hriUNF/EnCf4iE92Sjhe+T5KtS6ZHShoh0CmlaZcaENw
D9chd+qGPOxY+xoqEq2G1XW963MyMJGU2t4fk3yjqAFLWfOY+EqCwJjzKxmweVEF
P6xDWnZbLekFnp7uD6EQDZoHREpAss8b3Yva0Qp6/L3L4Ce5o5XBlWqo3yL3pqOQ
2+x0BtoZkbg2w2goIFtzCwXNrJAmBxBskN5EM72XXqtuVLIc2Fmylnv08UU0MYib
RgBJ/llE6dZWGXqSk0jc96+eOVwAHtAlcwN0vHVdNDBq+VMBYRGMPpSsYix2NCEL
lkaH4vT3is+PHD/ckM2fzr60qcNNaoaUhz/RfXUhzcB1dz9lAKa8x/S/NbvXtCQn
T8Mioc9NIj6WVC1FC+WcrT05IBXW5Ahq7w0WMwM1OrXQ/5g8qpYu0qES50a/PVpv
Nr9C3TtyBy4RXHreQSuCbQXuAlwiofJA5g2HEWh5IGWSSbjCGwMPwVCn09c+h10/
btS9oFa/VecM4KJADbsAdK8OhGefdiYYO/24fLUH2UC+0mspk1v7CnE/s2nUM1JD
IbUzYkgZYf2+EzX+Z5k07FaVGEyehEPncVeyx419ZP4+h/9HlgoQYKuPUZPFMdW4
E9O9dfvHs01sBkJY2FJKAMB+YefkC/Mrzl/vFFDQQfF1Kk3QBpTLMVGy/hys8MY+
phBp6ZLm3emmXCBPqaer7Ig8CXO9l1D44166W/F2Y1xa6Je1vlGXGsTHKXq5P3mq
R0xupri05N2KhyUhpcCTF0voROd1LKh+GLGiSv9qW2Z8q6YUlmbRrOv68XGz01rp
P92avcbg26/uc4vpXdJPkzQ17LJcy1oH86t67kwXtJR7tURO8I6W2dk+EA2ZlxQv
la52TFMCcaWwre/IFCXCHidNVWefFL3hWyXzSrnDu+k/H9Ehh+IyPAdWJIhjWLN0
qLTzVDMq3nzfMYEFX1dvN95yjGiJ5qI0zdE+v5JVCRMtzIV/MCMbBKlZ8LwmvU4M
P69BZKEF711U/tPkg/3EmD1vV12j6qpCfwTvcVfAoWSvVS13uCSQF+2z+ewKky1b
yYakPN4wq1F7tzCV1XslFrRUGwEXG1MADKU2xBi/JTmIs00w4Cf3XyGrZzPfooWd
4DEd9iKqaNME6S7AV2Zi9xbMPcI+bg69ITog0O+jOKWR50WABDxJbi4oba73N6KU
O1lEXxgWT6ApY79QKu8kVShUVtL6pXkgrLCRMJtoetk/e5CjcuVBltJ2aOonLEIc
+zdPHVMLor5bjuMiy4T7NK0lgJDeva7QKzIUa2EZcydHEH8HCF0z/bDndnsD1nrK
iH3BNZVukWSkx5BqbmU88IB6Kpg04YN4TjWORldT8eu5JauJDbve76WPmkc5bRe9
4sPuxTKQfAzpJrgjplSO5i98b3QN77poY/uoSTc/UmCiSTzaOrGWro6Sd5MA5Ep6
1dNJL0rF669LG9ghCS7MgQRdzk+zO7lZnKcjpc1oNNvsI2mTpzvw25qZRCmADN4K
GnzpAzpFHxMMHNqQSQRwM8uUuzHbyXNwsQq1jCEYbjcwgWJu5GGNI+ZT18HS04xt
WIR9zEjnEKyeQzyOF4ht4zGptXRC6z//tFX4IpRUaiFA8ohsjfRcTx0EpRK5kFzh
qctmYxynPq6ityjJYqEMRbpQKg6Sn/g0VbGpSIONDobM6pAcoIjZ3OXonPqqrPJ2
stgyf2e8k8NqHI9qFldAw/3MVwfXLeVVVx61PkEZnhAsQJWxb68KCHtidZ47oTsy
1YuPZBBFUD6hSbZ0ypxG+rq68tALuZyRHzzW0HMxSabvMLpphuakBuzMRggLEMTM
v8V99qqqxBU4TymZ2WJRE52bkl06xvRganCB4PzGcjXZpvYzolxk8ZCn4jW4BPE7
T/yGRrISI3n/o1NfLRAe1K/a9Ha1hAIiyVc9pfcQavT1pb9YJh5SvabBBRnUKQoN
RJC41+xxKhNAX5vegp+az3/NGK08IqLd/XDnUsXtIZDMsN0YPHtIgH5F2/GjnpoE
laA2D2/+x2BukWKIG/xI/s6of/C0W6B9nskgGMs5AUWm28mNaI/ueXYHU31aUAQd
3nWQWkwFQHZABXsiWWfKIphsYDK2dQUXd+duBgvcRNu+nCSPajqZ1NVX+NX2rALo
Ccxh+Yez0Eohi4mXkF7LMrFxcQ+M2PR8IOMb42Ndrgqiwt7l55NH8D9aeh69SdZt
riRA1LY97aQe8qvW5ZWHq5bmbJbU/WbfuGAU4pRPGMIJ7RqwonsddcWC9ywyOP0d
aApAMCtu6sQ6/XHx154I3707NQv7YOpdRZmb0tUpwzr1JCPN1QHU2U+oQwd78g0R
wwh/daVg6MeoQ9bd6CLpglXtLJbxyEQ4CPeUlOjCOCLvNRVKaz0Rd6IgLYX8VRoE
XcAjgNvXZePdZsYM6xW+uBCKeDm6PGhHjHqwd/tw3mP4Ktc7DstU9dOkijFCOYbF
K3ZZajyY1rlTRJsYeU6jQc4aagwnu5G5h+g8ztRqqbKyX3w6rOp5oiUq5WgXNwWi
dK7frh/RqFg0fiKq8z+IUeQHJosUI1jXp8dYE7bgauhVkiKosT//fY5coJrwGDd4
4T8yhhBq2LbLnrlOnFQJC5NNTYNKpLlysnVfjGLWNyKd7zs0BIbIVFm4vZp0qGtW
Zx+ZrazqBT58BujCLHD5Xq3Sp8R14vL19oPqiDVN/570Q4WmZyTI4ZG+YBSPeIXv
FxxnqVoK2BtLBveHUu+kQ+yYe8LKW6Ol8gMqnP/1XSR9/2nzKcNZNiWZQ+dThHoY
NPaTbc+NB1KS4cVzXAJ8SiBPav2doHpWxB1w+mWdJ4IXY2r0wU8xO+MjO9BpcA3a
H+T+mUqiWznzJOCE2S01kHAyZqyI02HU6ICuJxoC4pzIeCuElQG0aLmhbO8HF8Dn
QCqDeRcuQusmStTPGdPmPsR54zblh+sT8Ucr/56UAtmFRnyzZe3+yT71ELax939Y
vnkfj1RlStCjVsthotxOzR5au40KlWbDSifzqDAO+hw0UZVcjKHoBzlwIFXberRP
Dhkb/I6fYnW7c6yjraNneR4aF9nCgK9a3owOPjvxDfmOtHAAnUdg2ZT1cJ/nyN0U
QeRR/GI1wj5H1VpWb6LOLd/NlHFr7c5Xro7I/6L/CQQOrkyS07zfKs1lqxxxFA08
4f/weIXdNqAzOPDLKvjSHBgOF3IDyuKUvONljLJH4SJG50cp65EHmKhWKhNsAijK
SZRHkP6Z8FXPyW69OyoFskfhAJVPLsWAlOgzi519AVRvVfSTA4c4FHPBNtCpOELq
dHRGqhnLYHVWDgMzNnBC/bfxafgFA+2tOgEJTYRHAj1QblXK5QXPq5QmwOf9KR4S
b7V4JTnM+Ql2d8bJdukcdgCxHB0FP3hFZEa2FRYlzDgYOrybrDcvfcCYMEnWH8ek
Or4z3+cSTEYHMUxH8fNWosOv7VrIUsFJ/W+z0XTzXICUuEEo+K/dE6vbXJ4hVLyp
YaZMLIvZiobCrZ3BdRQsycul/hT4WKqfPFVJ+Z6q6b/rhOg7oTdtEqANcz4+9iAQ
RQu2si0l5HNbYVujQqUdqwkQWv4SSmTKFqhme7l0+pH/tlo0WVu9viicUxyPhSJ3
vLEEDYDdxB/QZvlh95J9gDfjkQpAZOm3iCjss2Q9r4XYJh13ERny0/TE6cMRmFrz
hhe/q/bfR70DfSShs0AHquneHIMdR0Fmn6elZ061ypLhQtncb5FQ0CkbOaZWlMbt
nBbSzUtmpTwzB1suViYQxvZ4i5d168sCuk5rSQ5mK8DnijHb3ZJiMC/LVoOUJJZb
FYpm3cEDwo12rZfC09p735H8oxjZMMWxyABzogBzLGTGimLNfWxwUHUpMVbNmcMJ
xuZ20Ose//u6kRMW1DaI0BNjozqyQzfuwhUGLZxd8jmnvJLQYLDhq8/IBF9bJd5r
UQMdJ9R2sOFPoc1w2FMSE76anjJc/WdzJFpSKTI5Obs6oej2bxlx5IfMIFpHSEKa
vGnKDLsHs1SI62zBl8su66XqXATkqsOLvtvMBGk0Px3vOQQrINmy8jPE2tzwdRdB
w8SBT4iT8wcb74LFxkaem8hPuvW3QnbvGlsjUutcRF7pZbowgt4NvyeQmlLClL5G
D50MtqIzVy6+aq0psMBtEBEfi8LgUIHYDpwWbkfOYzR9FSv87CAlNn6u547o8VIA
ofZg6dcGvJ2UcjECo3uHqpBJkBgJIZr2+xzwHaOQO3/iRSNJxBYErWebkbRXdv6x
xh5AkrkrjAEYYseL14bZ7MSi2zj68lM+yFFlndnAxD4C7b++o6ZPZpUF4VllM+xH
oMECsDrkUDIfUpt/G5oaqizsSW5Af9egVUIxztExaEogPHx/7EHH/n4Iji/rpHIM
TZJV9WLzCJsraOETre21iKyRiVAh4b7vcUWaCQNUfgRBeQ0nVS6TDPTQoT2Ro/Pp
vInj1LmvBeIm8Q/1QV5rrc2+6ATVrvs1fKS0FZHzx1g27H3SX83Gsl6CaNagvNQb
nDRwoD6Nil3SiLxWCeeemIDZMirIajngTl0ayhlOlPAD5NcqgvTtDdF0CgfJQ+r3
an5ugFFqIWgGrHduTy1U505wVMWqdwlvf3SZW34TGb28I36/iB8iWXj41hlvHzuq
sRVZE/6Dxc2Qekp2FHX6w5fqVRWbOhkoJ/a6CCNDlZcbaE5ecnCSeZh3u25gaOqx
8fmElvpQx3qiNMvu2uap0ft494NGROKb8Q3Fq8AbUhWzpO/qYk0hmxs1cjCqBZmk
eChcso74M841r1qrXBO4QHD5ymjifahEXjqD30asANDdUHtJgJcqjD1FUdeyssYM
Dm2/xOvJMt2P/j9hJ1lIwdXEp/Ck3wh/po+DXWHXraIgMqUUGFKHqub1LQjUFX+U
tZnuCdKIlx0SBsCKZRZDy/QG3h95txwSHE+jOZ5QorA1piy4VlTlocta8a4i8/7n
THPXs2MDSh3kAUC1V5kcZTwlX5LxpFFnieN41oLqhmHhvAFt9DyHyiDUOCh1klSc
tZ+UjLHUG+nDhTBwLiT7zLt6ADvMg0z3L8ej6qBFeXcLuhlngoZd/oAqD08Dkma8
kKOb2kR9eS9Lp69XMuJUL1ogUp2bvlykmjZtFTqHP+hZIrK4P8vLVErxfcZlmY74
tluOv4hy1QpymAsnO2gFlhm/g847XC4URkdxlsgBQhLfMKZlWm0awDlr8khspijj
ofN04vdGsvU47RisUjAjNL/+ykcx9D3VO1X6cMQrEDAnHzbj5mdXl/ky5vGwc0de
bB/vyNpeLZsR0sa2e03kjwurR7zIfBIkAFudNWvBWgt2dKUhHNuQ5hIVCpMGMn69
CcZ3FlJKYTxJpLGE+oDuTfuECXxbZ5GFaIWrxFzVINQm0fVOh9P1uKArOHZjAAbm
nylpJ+PPDxYKMSBw9eArEgWRj8x8g/Cn/6OEnPT+H8C0dBMCqofPm5dx9svDWBG6
5wqb3bVYCKAbTVJdJ6+1QO9LiO53+WZQLRUiOqh8Sp0t0euEH5F3KcgfIuQ27Hbl
9XYcIKF+hnEVH2u4eLaPCChRSxt/XXqgVsTgN8NrQR8idhPcbqHUu07Ld9DqVYQ3
hI03WxuW/88b77eRjVRBnp+BB0GbdimTxOz/xnGqNN7ADirTIyZfl7GZ/zG2XaDU
WdaRb9wVyURACNrC73/GjoJ8jOiaMt39513SgqsbfPjoPZMkbk0L+SsqVLjt6gxh
KHkrzQUJoSNnvqdLP03VI4Rw1LV8E4U5OYnQR4G4N9N/HY5KrNs48IMivBnumwtV
wNMaGLQwPSTjrixzkIijuUOEcdnPqqp5iVK6HPmSmyz3w9l3wbzBO4klzVY2DHlm
dz9ms9wpXaFYt/z+JtGUXs3bLauz6sAulDNmpcRh6X37UJ9y1vLihYAfi12lNMQW
NR1n8Ziorn92fSDcWIIcUoyNTNoHnd1vqAaQ+rscyi7jqlh5Ph9vR8yCspYuh52V
XiuUoYnpkgXsUkPzWicy1LgFOuseU1xuWwG/gTgS8x5x43sNL4B+IreRDWoNRJGM
rFYG2h5i1KutFKP2G325T68meiPYXvyLm6HV82q7T+04N8I/5e5TyLpzK4CeqsgF
ZJh5jZGJcxals4GSOzzleGfKPgliZKBUDSSXEPNkg7pZzFNPcmkrpyKuaiqKITbX
dTbGWdw1tWsgXSjo0+pxRQg2cJ0PMjgen1p1Md1S3EUzTUwWoL3riqmU9ugPt/sh
mVrjPTPUsPGgWuT+7eMIKtec19X+hJcL17rrlnm5CY8fCrOMeS0X4O1zX6ChUo5m
7GlIvwAhCcgHJpntQU6BKZZ3y5PBPHuZD+eOvuzKBaAHbZUzl9JDzbbzMU+pMCCo
P3hfdLTEny4IWh9er3LCrv+t5hyhX4FSyZQXZcvitxMmf4UU+RCiAyVbVSvW70gl
eH926mvfCH4l+NsqJpetoIbXHvtSOxqFEwEf5C2pSWVWLoWLEHdjZS8q/SvnRo4b
c2S37o4Xg9h76zyXgI7qIEwQ9LvHQGOy/mtUnSeM4XEIDxNSu6/KOZeAbKAR34fQ
IVbMWXBr+CNRsYCeip+tlcJ/py40XH6FUwSsZSz/j77vtTLZq1DmX39WVWJt9iLS
8MrEs+hr38qeoGTSZL3iTiJjk6z6+YyQf2ZbMEpOZRrcYF9Wt+CqDqekMoTy7dXg
wNNKiNnvvdN2F1PMN8C4jSo+j9ct9IFMij4fGd0uAbFT33jO1z3b2x7Bmxp5Lut/
+bDr342xFgad8AT26BHVrU9cgbqzWjtQwvzVWYngS2AwgakvWp1tFyJG6p/4LWfK
5glNM7ewoNi8WO+1ybDXlvtEGz0MyWgx5zRUHkGUAoipep+SQUK/9vlVtceoDfj7
Jmbdub8ODGi47H3AD85yVbuOOOk8mjQjFJhQK0otwdN17sOt76KeEtjn6PhoH/fB
frpI0BqAOG6M2zFUMhLbNx9MGbahg17zNQyQkFNtbDX4A6C1Wbj2XQ/s0KZDcsB9
y8+dqpLxNMXC1LA8mXmTDTY2FmMJ/KAbdpPxM2zZuCNQM62hQnbtto8fm5u4BvjV
EhCtqs8UXidNlIomOph9vAkNGiMWMLwTWJjQNhWBdL7+K1iY3FOnfJDB9hpT4Hat
2Ie4V+ZlWfXpO2Wni9fx7zpmIzv+YTPDo7ZmMB5zFvdARIf0P6rqg98uVoAMta4n
Vufd1EpOIClLT3vfxh4J9mjt3z1D5LfbL6/927rsxEyMy0HTAb17ZV9PgzfUDjWH
akDjPBZdxkulUNvojdyq2ekmc9Jp69OBLu8fVJ51H72a/DuYO/SxqKsfeh2RoKpp
JX9M0q0bqrcqom22B7xpA95OiwG2g3zgChTM2RJhrqNJqsleLzjLsBsVysu7AUkx
X0Q6W609fGZKjwxadTciZ2jVABsxdwdudX7L2Bqqgc1NvdgWwaivFpCtjo9w1q8a
k4nmdA96fuFCdY4Zq1pH1noxR8fwTAwuXGFuQfIZRtp0Bb8OuYmIYUFWm6vQV4yP
Sxjs/bh7dm/tFbI569w6NjBTv1rplR4fmNHaBZoLIbzZcZfJLJdqTPaJl6SifjgK
XxGsaIar63QC9GszczcjdfnJ6VndA4ZPW1zSbfqYBhnopd4iDnb90yBoTunqGWoS
Pj/+urMnlbvYnjo/mvitajX4O2CugFgmuNToEhoXTVC8eSPLPKVqEUje4J2ci0hw
x9+DHTF5pCoI1S2SyxIL2uvh/aji+kig1TYPk0xUf0lRr38VFJ0WmfHRRyozcT0D
/JM+ecGiIkHRaRJaZkTFH5VuVo6vsgVrebv0r845ZN3LnYgASV/m7jpqULw6wA8j
Gp5s9+1dSnHcrNyJfvkiywo28Di53Hug9qapM0txDLjerPIKKsADCEOvcFgdqois
9cDL6Q4/NvX7R5Pe9kf8ug7vfOffEXIH/7BINcsF0QKXzZs6FNyEqxlqqX31Vt2P
npcDiMrJJ1Yhcc1X04Fd1ZapEkbuMxA6zZjgJg6yZK4nD6mbWajwcKGOnxu9K1Kb
8DPS+XEMRo7+pz6aFKZsjYvMEapmS78INKlzjXd6LgOjbJVfczPPl97qQ8JwhkBX
v+RYXk+SjEF3Oz1utuGJTUPbH7AMp02LCwzDIGh1rGkO7WuBBwCdYEaWCYZ0EQEK
80vgTD0cd/aEghYZIVz95z+LYmjMtiOKrIY9VjwtbnHYXd2exjE2y3AN/h1H/VnX
rXDq9+E0mrmC67sZJqXZBHrOEkTlAS+S/38OxS9k43ihN/1kb9bohyRYrQGRI0go
3QpcTPBLlqZuuT3BlorypF9f5tn3HcQTd5f73KTYk1BUStSKnuWp8hrqOuVwIdK7
1S1amCUuX33IZm9d2rWjNFL3XOM3/I8McwgS8R+AreU0karIChfDY6mRUJjWrymT
fqzAtFCzOpBNXbHtd/NUrnGhnEgAOQwexEP2P4/Or0Ys37lkMZLLltXTlSqE9mUS
LRgSoWhg4kdcqmWx2kAUNNxUfNjJv+l/GqGUkpBTs5xVeGqO7FiYB41/bG2m3jhg
W7Hv0ewFX7zAq/56BQ4p1OWitcy3AvJipxIiMA0Lex6X4+FeCE9y7DUmpsHtsshr
VGtm7RADmYpOoiRBdNHOJ/UZzuRa6DT4LpzCdKWTU9YLFlXVoCWkkbwZz5OureVv
lUXEZtkEsDoWM7khF569wmH9aFd5wW+NSva9OfSwRS/uLAFUpFCTlFR4R/qI+Aap
6cl7+eaanznH92hn2lKhaRq5zNm79FOxRPBtfRc5gzV9JYdgmbT9TJyvSJMXC21R
LvK+j6NLZspdISOKSQDhOmJzGzUHp+k1L8YRQYchP6fnXg3BqAeYEKmWIbbVoZmF
Aj9raJYLjiAGXhDMrFRfjz38oCU8vG/f3N0vu6C/xpqOmNC8ibUH1S+mKJ4Q3scR
MjKafchQixd1D4D4FnXW3qIz9id0y1+UICIZftYkqg87b4wPTxeaKab5rCxvxd3d
WE+MbigQ5an9Xh3lcWFWxKCd7TtQPohHGKDDCw2GFwIZ5dxBz0VVTf+O6R5fBlPv
mBLHX5Xpsquq9LeFyPIjMYB9YJJ0sY3/ftWAZLZVr5wL1x50rfdZJf4WFe5v/xNB
zgatPy3xuzjP8nyQYuJLMk8Ab71b3Zb+CT0MYaqkrBpohwVV6u7PIT30lHr07Enx
yv3IX5euRgISlDYfpgh3c8xQmHDXDTcpK+VELMnLdsLsVi9ZJWQ9mmt7CtJZBzpm
dn3v1Dlu2dNY6cibivUgubQEPjZOCqf/ibKeQtr3ZhdTjwNI6KDC4r/OLJgbLr9f
E1M5Yh1sGcHG3u6txNjnsMceI220BWIQVj4Cc2ZajPv5iAby1YDTwnZ/P59b/c7m
EwAo6nrLZSdmkjT86Kr+OD3PZn0JpRN907bciCTfUPqjxpyFIC8jImmfj1Mt8Vv3
Sy9BkNW/X3DIG4XJI0n3Up9L1UdEwKjYaRgEui6Q6CMTe39PpwpRoYmg2PyxrL+/
QdrH7XEGooSk3er7FOu587YPjgtNZGmSzZ5qC11DOR2PqKl/wn5gDeRqIc7h6D7N
vUfvNLRYRaopQ3e15A2kOAqt0Uypr8AOHTDg6w1ZKe1pf9a1Z/eOizF/dq0d8uft
g+ncl3F0TiA4nWfTRcC7qc9Gt2lPxSBxIyVVKFvDD5CwihargfCQkRwzYOXbSdfS
dABSnTiPO+e1/L31a3feNZNyqIUFLycJcbDHA5ZHWsc1WFZLYSW9zJklNb9AIqcb
dXq93UediZkpngbgeZPkrlsvAGYzAH4sgmsGMzI2rNTJrNsv1Hh/sB5D9qQlmyit
pLFdGXsHa7Unc0eAgUXsmnnQGSOMSXWq7PhZXNggUTLefLs2UgODgYcMEiCc1YvU
ZR1/f7g18+CnSd404mREc8r2AMJ463YV065pd1eo+T3w68vp94dzN0E3434lsgeA
VcbaioypgPsYtMG+J3WJzc2mUEg0nRji2ua2S6emJaPMF7gd0x8ChLQA/3biRSbz
VfdjA9RPZ/ES9Cl/gxaxvHx9HGBSqDe96h4GJW60P9vqUSoPuTpsl1EONErhzrFG
PK8pYeqmfauYhrv+vlCgXv120PcGkFRfj+jA98Zz0e+hrscZTybscXkX/zsl0aXx
Oz8Iu/wu8MkR4UYQcQ50c7k6z/9GNtHI26DLJuJpCypGS2kwRSIXY96TJuKaFGdV
xeFq9XIugR/wdZi6bYwq5DjVOJaANBBID6hpx7FlAHXPdVQvEZ7CQkD9AmQCoDk+
CUNfWZy1Uwiq/OMCzyXR91nsz4n2m491zORXGOUE94ZaQ/Ha/DarXVstE0nIN1UT
Mjn8jN8+1u5t1cXc9n36I78uO8M36F2xtQId47ovCOF4gPbSYODchSS6I2PykaVv
UvlDnsQs9/FcOax/yiWu2ssP3X+qEDu9DDdM4zBPmmvIQd2mlS56cmYOlX/+D/85
g6jepO6ScCdqz9szSqQ31V/mKAkwp30LG8WJteIQO9pnwpN8OqQtnFpk0z/RnWxv
v20il/LkSpW8j9bqKPk+uJHCbTPy70KH5FJ7bOzqqre8xFjYiF9mCnQOyE1Q/JQr
XPfGnYpOWYC+PNNUsIfCk7gVaquYOYcQryyQ/y9KM+5iYgNl4u7qx322TF7WP3xY
VrvtCVyceAnTJvsnNyUdm6F5Syby4WWHCgHMIXnK4wvYQ0MbEHRdZwC4BzDSR7G9
NN3/jVBv6XOxXf9sbGIRAAQZ2x2IXcGjp+sqCvShOovVeaAUtmLTtudaf29Eh+3B
GwoGuL0qvUctCQFXjzONOrAtILpJiQ+1VAIDTxH/yGn2uDRSZ1kZzMLoKN5HSD7z
AooAcPjaEZ6eZG3OtLKevfdTfUJkFEfisAOJfhqxK28ihjfvFLKHMQR2W4ETOlpK
EKWZ/+w9dg36MO0AUPD9UvMCzobwzZWks/CbKWmeEDoycyrlulDJN6OU94LPza8r
mDzyigYxkqXR3i3yDDxfyVmDOPv41yhfhWvQs23O/GkexvvPzAvTsxAkrSUWQHNv
S+ah9qwMyk1DP5xXIh8eakA16lt810xB2crVjGLoN+YUWHFFFrDJmJJkbBSxN6RH
5+pURwHv6nF3SimEg8Dm9UGqsPB7SBIg3FeS4yhYa/OrHs6Wap3QZByco6S22FRf
+Km9PyAL+98z00MITnNN+QKmS3x74K3iEy6su/1Mu2IsfXvIDMuS4QSsm/3lOmYP
o0Bzd0CLlz/b9EvU9tT7S3QW3d23xT7GBkkGcEd5h1bfu0NhxoB2czEeNjqpkUL0
YFYqUCeWn/T7itzL7ZW/I/1ViFvVyDZ7oGJnu6EGWxE8dKRZFy9kJnnDajX6mmIz
bmnFhk/ZW4t/1fkSjcuZhqKRbSFM479i6U2SD9ZE2l3Owj1gjWjty3UsyaNL4HBJ
PvvLLIPKE6Lan1l5TwwcuknsKgAl/Q+JgXkQuu0I4rP1h6+3P7mPCigQllol+iGe
95y9dx43ETyGjMX9mycpSN9aLnZSvuvaR+GM9FkTBC6ywm5hXtpQy64fqiagqTW9
MEXc/kjPcuwxVN5swEroyJYZH87Pa43XC30OZaLVuiLUGeNKWaUiDkIelEEQbaxG
ychRLYAs/ScfVdC75zEEP9eMU7NQVlhi0yfduThelp00j1qq9utzzUV7baXl2DBx
a/PG9nTrVPu/6sgFoMaIN46tUmw9qo/ZeMeCD58mgj9AJrMYh8oB8uWma3tPVO4A
MMVx5gK8Rhcek8NJSXSzFkFL+hJZl1dEHsjqn7PZh7AP7wQjiO8NtipG3RjSSXAC
hUjO4hwEtmtrIYl3ER2nGV9xD+/JDwyQ+/Eoi3TNeckTj8GnuC+ADjAlOLUKCz9X
QiTmWawh2L2fk7AWU8KS3m/kCItTiB5x/U7EMV1/LrEU9lNFGpDlp5crGuR0bng5
E9Pj42CjFPwtN8VRg7vb2uyJ6F+ZKjxMD52owNFKK0Xz+c4OTB2HIu/bQzZKlQZh
eLnwcDm9gDfMTXF73Jzi9BQhv2EZPVWrUDBQtZTUyG9YXbULAKiBdlWYxY6zZIfu
6nhFxoG0eWwGic2LbaZKEnxMVwCKd4PIUwaT0N088WZza0M6VBlApXNSMqRMHRAu
hrRhe71ujFd5hCUez7bb6OA51KEs93xvOf8fvY5sgg5V1mxtqJKjkH03yJVQa2/U
t2MM8Df/S27lGpdUmUFSqiEGDBKdSrSWPLrWn9uOqQ5Dcwz7Z+fImStA1lvY0MRi
oK2WBEwPI/EcBT4NqPoy7B7iG5bXCme73Ds43zYYfmXIUOiG+cKKtvq3kyOsEsU3
8k2h8ewicxQpD3HHhhJVazgEzGCmiGKwnHHvvihZSDE3N/9wPqdVimLrQUhn2KgJ
J5cIbcWXR+U+fK8i4zr6qfwFKhSDtIHntfNsmgBa3p8gHZfKuNPg9qNUafnv/iqZ
KIqZz9QgQ/VYo/BmGzXGvSStY+BvHDuQgqQIqQ7zX0NZAGwHqB6NIKfoQgCOwHXk
bM+5a6/uAaMna/ZVrqURHXDI5Bm9sbMEsW+SGVlHulbOz+1HZL430I8nXQ2f0HyV
j1Hxl+Jh0nsiKHYRq8QuI8zAAbHuCzE0mlVvrluDRMfMRPNaAbSzm75rbKuUAoyV
QUuDODfADaT2NDqknasTGeQEkl3boYvHlKUePLnlsi56Aw750VH+ArGv/MBfmMAG
wtPab7UxT5bnj8Qgxue3+7W3K5HFhkYyZLGwEK3R6vKodCCvTvqBtXTu3iVsVxB+
YhIuI89Guzv1PL0CQ1cGqm0sBwoO+gACWYJLOonHnTnoon2ogccJiosEDLLXJbXI
YehFA7hOUQZUhyIVYFKzrPitceAC2vYmEHJtWsjWAIOUL1R2EwBIPIscph4dg+xR
YH3m8WJYTci2ZV61zY/Vjc/akd09NynsTELZ8v5FId+FpqlGAER+UN7X4gSXB+N6
k5tmZfqXdQrZ+6XH5xTT8MG0lTaELUhPz7upQW+NQshwldpbXe6cBgwPGKkNz8da
ggE6mcDS98fNUKmFAhaUQUgJFXyGPkYV2z2OWAYJAmQF+YNG8PUTM2GCh7dHjByc
v3uo5+khqCPhHgtn76ndo2K4fP2sWsq6SMyu1cwhiICHIobo9SHM05ymbugdz2Zc
PKv4K5xi3lklb9qHJE7O1JKsVVAVebe2hKMWD8DwiVYH4oTqGtlWK9DzRQkbA2/m
Muyvttqxe0UJ/oagF756F/jBLeK6wkajsJi38l6q0vqlrA2DU/UkP11SPKOXcSEt
hYRKSDaI4IBOwitt6Ii+C3ABWH2mNppR0hQ+/rziBFjgV9ah43atIdEJ+W4No44v
Tp7Tp7iG7VgrgAVsRO9DsHmc9id+6635q6fkZkhOWwrorVMJz3MsXDDZ9VaWmWdI
+t7g+2kDnJNvrrUEx2k/5oYfO0JNfpfsVGm+tAiHqz3Z6IWGzeIO7Lgbjpa1BO5a
58gZw3foCl0Hp9GP33okyi9hCXjfXuQcoLSicPr+6nJW6svabyULD5y/e0i8UFqp
VSswUsHvboPCQvEYY5VuIKeUXnOcyVEhS3N6d8U9buObnP8izSmV42Y6ANyORync
yH8mJ//NR9if8EZ9oQnGwR8dxwLhxw4WeD/Kbb6KWHoq19/tVgqKt101eM7V+GhE
gjRgdTNqgYCVFkYpeoipnTBTnv4r48Lz8iGBvZAs84GAv3LnxNGRrEgjlQaSMf2D
jaEVIC5ddiEpGVn/RXxm14tzeL/Q0RkVFz2qDJtFKI9h9wCPU/MQwGgrQ6FpFRz0
0bASrwSiP6WDGYVmS1VlH2ZUOzXCgb75hJKQEqV4ejbu6+1mfzigRAUc83ArCwC3
GWBeNoaMXkRXJDjTVsvHG2r/8uE+lVYbB0N3Jy8QTu9nVbJ1n1k4H0pM4/+Eemsa
Kvs4VSRFCJlKVz0453e38EmtxUr9ANJrpdeZ5Mg3JS/YhAnrcOeNDxCCSRYqFuKT
Bdahkg0t5RLGP3r5JFKhY9UJKq/Q9NmTrF2+cICMANSWrkJ9ayB23b64Rcz8O2sh
YQP6wXTtRvqnTgBLjftSPZMK1FyU4j7iTwdoX+OlqdlpzXgwb9MwUVj3v/cm27iY
DDvF3UiKXOs0TqS78TqXXjZZyurtixScWSZGHy6TcGpaICD5biByLOO270IwfSP7
FIoHhB+5TGTg1DpCx9xIhXirT3KPm0U8ZDuSqZjCfsT+2VmrJdSt0BVrGziF+y9S
BdhfDXgXdWp5nFf23rrA8fBJ8lBF5F1G0PmOtE5C4L4YiJoPKtf6fTRO0f3ZxcSN
6fOSBU0OMSpllEzGd4321qsXYpGdIiVo2EOs/9RcqbW22byT8TjoLanBoGSZzQav
7k7hLXNF1eYw4rrNcVc2EIUWl4owTceKs020Oq30fnvS//JYX+5rxT6IibtPrPm6
XLwwGwbTDzQo/Zi2QfAbXd9EdDJkUYG1RNH9TWFVde2o8QvOB2joWRAixsEsRuu0
wmQMoY/KcfC+fLkVya0/iL8rhGI8Ka1JnmTWsKqjKQA1F5jUBeTWGEpSBLKclQkX
qhY2TKaGTtxnOeU5hof0Tys9wvt/H/M69v5WhJ43AS4JKcF+DteSzKERvGWR/uo5
JtzeQHa5ch5Rm5IaBEy0SbgDBf12naSiQjAiZ1/B7JQ8K105IblVE11o1kwh8Qxv
d1xAtTPBNzmWfWzi0rqUXYXmnrVprvqe0Lez+f30LC9WJG7GLjbVMHAU+PsVUiAb
taD1mcx//BPbzrsUbAkqFzxAht8/YVAg9EoskrbXO8TzpeBfXUCgiOIPnipfLdEj
TGDYaLTRG/XEvCZNbcmKu3IvtUJLa+FEc94yj9R+OWtK36sVg/Jiybpist2lyZny
sViFYkxaEuCyJPYd5fjGSYQA/pLyl6qws00Qbk9vaospU1aUg0fW6iNQ1QiRuFcb
lJp+t5vng13jJdp84IoWPO+OYvRmCnmFjUANy69JZqNA9btgojfJnmuESG4foRVM
9WI6Lqlc1mvO7cAn9PZKOrK/Ma/PBjTa668OWkLEYA70qPi8lqp0knv54XqwN8BG
1QyaulU+ntU7sOxR+G+8PzT3dj2Fn/oMJW0zZicILKd5U+4TYfkUBv19/eC9Dh4E
eCUoIz1jmBQBfrOM1SfAQAG31ee+vZ/WtJs4FXTuTfGpjlQ2Dq5fD9yexeQS63Yd
s4QR2/o+R0Ky5CkqFd39jKXFRsx24MNa3MIK3uLbdvyEhyUa1KQydmEH3rX3A3Sq
gjr8HcV6qioH8WxWQsRXh2Ofdw+xY7ZG0rapeufhzEB69On0KP3DLcpNviRZ7MIz
2cRerDIZgBvHrIva8pobDUTKsxME5t/8oKOwd4MtR6ASDicqWEQ+vHrMKG4tMZcR
0bi9p4Sn+PByLOynXDc2/u+8dG7p5bsJifZWhMFFpsajkVgkB9LG4SfAdQz6vuxT
45s+HkCz/hTF6cdNejwgbMc6wL7UvZBINlpsju7uLlRdOtU5sTRbSOZjgtIojkTK
KIiL/Ypoj89kdhgKk+PO4AsolvsUMdfiRb/MDvZFa+3/nCwhGNZPQY2dhTh22cly
n9PuWGNkPoB8OrLze8KMrXsRl59z11Yr3frnUx01sZHsSs7yLBLrzDDYBteYHmOw
hDx9X+olxgyEI2QZAPT5rC4BuTkNjV8xW/t62PsGIj+X2hjmJ9pBkQbPTWTPhQhn
JotV1RrEwyFtSDiQbFjrAebYL5tIf2Zp3XCBNlM0kLYCtUUwzbax/SHIGxwBz7Vj
iHRUvA9QfsB37dUDmKp6sOOZNUpna7CKwtIIJkxRyQN9qeA2Awvz0dBEDP7iAxLR
k4uCEdtJvN+JfiRhn8JxWG+3dvwrcPb61LithQvwgLTVFsOg660E+7c5FVrCe7mW
WGFcIPml56fc+qJC36kP7sxpUNDoP+Hj27xcJ5g8dkcr20jTYVf14PHYWPaUbWxq
iI7sbjJlEa/nWI+jzhrCtUpF6nL6iphlmcgvQ+LmqvpcF4feL58eUo8JfbJAYVDi
/sgvC6sH7tJmMUXg7Y+5EA4cXuEwf/TDC1uy5VMbxHDP4Tr2/XZDQFf6AF/RQpga
KN6MoG5CoICBRYf2rXmsWXWWujH6bpzXNO/HSYLckCQuTSaAgVfI/rTVdBXRnah3
egp59nR1aSbaseobpTyFhReakCGa4TFIj4iboGZY3EYrv0h97zUFX17pbQKFv+61
67nEHWnUfFMCnu06FxPKMeCLDSoU0zSuidwIlnp/LI57dSODfavKJLmLg+PyIp5m
Mawhgx/rgTjV2Q7Hhnh78+ttw5js79uj+7YGpSP07mr6+znqYC+lCfoo7PShdEP+
tRO2RaFncOKGglYkr2DiXaMf2akGBLGS4kOTBGYbaiimOzyTelNmTfo+b+74soXh
mAZIm27rwbxyyrO6n5lMeCdJdugL/lXHX58zphIhXOk9WaC4qdT/3CmSMh3u2IoH
n5UIqi6JldyIThcVYH8BH2I95KwafEgt7lZoM2Trj5puwY38Xs2cktYsdqOqCL1a
fMtNSQBukNgEmn1164KCASW2dgfPaGqqNMQ3ONbwNObS5fTvd2muWmb8hqiPOVHL
v02m94VZlBMBmLXvseWtju9iDYjCn0+iTskHMo1cy0Mn3JBIGSIhbFLa4zgdRzzx
NbkcSLWNEABmcgwZYG1yf3YttVWKhOng0Oby1xKMzAWu2GMIvMS/+ffq3Bpyt2R6
AdOkTw+gyGxf/ojynIm0L03wBUWfuhFoQq6oDKDf53FagkCumSxUctcekKoFz8W2
3JBy7tpE1v0cDcWQZfB7MiM7V+4G5bejySanqXobSGyTvDljAJLihVRgP3zzBY2d
VJkxGK1q8fylX05NDZR1xuMltFMWdrVFaWY+ZHJFnqraL4srZc6FgeLBZTkfYMB+
439Ggz9qCIQj6SV8gJZVc8UPJ6JBudSsUhjrP7ISbCljypQ2aDUQb3sr26mXqe8P
eJIGb7sKA1wNNsR5nGXGrDbNpRf8WZ68AT0R2eEj+NqVyMCLad40SNN+JHAiROkY
bYANIdd2FTXaV6UFrmtP0SGDTC0WJNyiyGFICG/MRciiB80CS6Dic9t1gBM06aYN
cTYt/U2M6Gp9NN9gxAt2ygK/JQn/9TUSuo6YmfdGtWCrfX/MC2hM/IJoM4p1yxuF
8meOvu1xItA4RoFiVnV79cW1thxM8zvAS7I6+feIR9f4lL8MLsESypJK2v2vN/Du
iWcaCz8XX0G7SR+aiP8GOdOmGTp2FATvukR/EK4QNy/i22V8OCAh7ZwghCw1xunr
wC8oivW4QEUCikWxlbYhq57BIRjbkKyJkGV/7jP6DemMxiaBzXUnbxMun8DB2KBs
QmdVthMfjy+cmCd2b6lAipxZTfj8UXb+g+wE3vYfuEya8sK4bj2MeZU5E9s/oxWh
lhhX0sBVKgQ/z4T4JIyHnSEVtF6Slfuxn56zl13zXD0GKCBIUmprCGQrmqbQ4mzi
st9JX9rGHwszGk+a4G5+oskk8khqd7rogw9YcAloEcH0ZY9J3fYf2EdfdLDM8W7t
6vmyefwZleocgprw7V9dMiNrraR07axFbnwdhVEUeg9eYbcCFSGKGlZs+1UZtMHV
BTS1ts3iz1fnT03qdB9TllsyuWjHtbfMu69TNesWuSJZ823I9zMN5gxFK2xmTykh
1IydaG2t0gGJbzPeiIXWfL91JpowP5fG/TVnBireKIoNsLpaGyb+DbyNcs+HrC3V
tC5akpQQJNk32xQQgsAo8ng/lCFZ/7w8d70ptAug1ASOMWsUSzxADDo6qFtVMhjd
yb7Aix2MylyaSFBDA3V2INMgDPCJNP4N3eMKr1d4rzF/5B8HDy/N0pHSYB3arGBX
RIO3WGS12oB1voG+En/o89LfIZ1+WLFO3Q4ENiOxMf45uHeWHAgRKxhDEO93mwhP
GUuEDBUUKYsub7UPUQKthgBNkc996UYjbXYUMlxLpKYUMFhqBBy6lojc5lhrUQBd
RtjiYV6CcXyXha51SDnEpVzqNKfrcVVViM/75e1iYg1ygkcUuZoAFcSWlIOiletX
LxOie7C3zqMMPzWskYBUbua5Gp3FHUrLzoS02z2BD0weRrEziDNJhes3aidHjZpW
Suzx7EWtlhGlYiZJvHHODJFYSvELfcTBeScTsmjVuloQ5KAKDsmhfsjqTIH8KGTe
kYCqkpXo9MLbrTw9h4ccSgchv5Sigo2UbEGeGe9HAUw3KZCNp2kI/c922CcBf9RY
22b3Q53e+SbcXCmITOZfp5H+MIaXXTnHDWvoSFvUWXVWzV34UalUlr667JyFaRve
rz5PJaO948KyI1AuChUjFslN/HlQnf+cpot8471ISFQKJG7/k1T8ikN+vTC+5FjF
cfcz6BcugNe/szJ1ZXU0YkYW+iHxZRHI0uKvM4qjpmsCn8rgeBylvHB+gxN8+IN9
zXYPvzl2B1V02+Q4EaZz2x9ML1+hf4ZGow3+iz8mw90aw6qlYIMunK+Jf6+5dfqy
OXhZNmbWIJsC362dslwWI5W6O5k4d2P2FKUQxJTrYMbsBP/tu/gArESPbiZ72Z2T
gFKgoBzgfZ80pJxAdtAGuH5ePHWrGWNuL/vpS+c+oTjyM4i2pGQqZUlVgsDlsyrt
ygN3jLA6/wpC1BGGl0p7OP9Zu4IZCy1W3LHtO/Q+Mo+c0WoB7oq0hcty6mjSizF8
TiKRpptxhLVf/XWdaiirz+tL9+j0y+KJR8EC0TtfM7TdsqiWPwkoSpYJMvjNTtUI
nhDTP+3sWmXikaFd9/i2TWtnV751Ekr2CY7yUDtRTN8TP7+AzJRHCmWTZlh70Ikl
EFP/7JCDkWEkWGNK8Uuhh2vkefJLw7RudIBGxOobKq8+6vVYlG9Yrpeq/b+EMBRq
0vhwjvfrccXnGQbCeNWTEIoMkZAYsXWJ2MN1CQixS4q+jy4/EUE3ghLl3Rc0zFzQ
DoySoXm3gloTss93E7sw3oNf7rNLf+yaqQYPh4VBObazhzNpQVLohI2RwRLGVRUR
TnhDw56bWZmqT21ROXQH/xT5tE242XE2mwOnE2/l8UWEBNL58OWIUWKvtJDrolhu
A9t1ceQU6u+jjKLA5zRuEqIkqXPGA9ou1ebxAn/D4e/QrkFChCaklhssML3K1thJ
cRMjZQLBDQzMvYMg38igKeB8U/yYW2jEThfYlO+pGQQ7ehI2CbyNEsMy6xGyXdzg
9t7v8YUSzESb5UlFROxu0nIOC6zdFkWBhT871Q+VhVKE2R4vpOMrWFCZPKGkEfbO
FumRg6JS76Rfl8Kt3RzNZwkg5bpsHgSpjoLKBY4U6pAtGfgxjxJG3hYpFDWpTFK6
6UIJKXG99fbBq7R9GSEnPzu3NLwMyvj+mO+B06O6dLNKhuRtu5VfF/E2WuDT15M5
ncJpW6xC7uSZp/FPCyV3LwD0xNbDgnq5JuL6Qd+YR3NQV2RzJEQApKdk+nLr++nR
0K9PyrIBGyvyamOnrlBid0GhyjMLHzDcygzkIw0uwjKh9o02CJJ5vdgJCCLgU3Nc
+Tpjy1KQ66w03U1qgczPQsxmdKNShSEdOaJTqw6ImDeMbXfy0/rJZty97TztuLeh
XCYg0zvcEvFpMCpKkPQLpSJjwcAhRqwpzd8TVe8/YiQo8ISqwfn6DxuQM+QYvsBr
gsC3ipfpsgHstCMpzzH3m7B4smV0Ziz8NV/WoU8GCIgEJnwfPIrYY8gfWWQDU+D+
bWHeZIOqmMuVCBmbloTqG+rEycxrktUU6PPewJyBqUoesEbvi+wDsCCo+EIWEaS+
Pu8vC7CDrvun/YsTxULQQwnyoAvJiuuzXDl4PNu9xBUIH91MgzJDbwH1mlaPfYUf
BZdZPppx6L+St+zh9g04yFfu8yWUtbPEJbFCWDAKrZbP/lRGFGtGzpUisvR7UN9R
wu1Nju2hezZl7EkpJel3267rAP0Li704XpC++QjAZ71xGNJlE8VR6bVYz+QdZW/y
MUP8/udgtizY1TabAgE93MMw6SeH0xZMmNmHHG4BWeEnGdl6AgpS+uo9CQ02HqK3
/A4bwBRSQmaOsjsTsFKEfKs9xhIJz+cJC3dn8xdf/AVUKEfFmaijXZldmzo3HCj7
+b7pjsvHLqzAE+gcA+kOw3nbgQnazEQz1j5l8QjA4tFB5xBI/G67T15X4VA99GEn
prNrMQJNJMMDQm7YrzlJ3QP94LcdzoEZNJD3VbfbhRZZ6rF8ZHDVILE4ACNNgYUo
kchfIPk2m0UNJwRTJ2LKWMdoQMzvuMNqyk5FdrUKNmTHke0IVqk+JqDvMDHk0QxW
KbGhZfaGHB1RzlisDP0RzLf0DRb960/3eCxsmRHUa1VuMF7oY9B9F44VEaH50Of3
+ePWksj3AL0l6Oy/MbjIw/k6KOABAX6CwSSRl6p+Ii5aDhzIIaylBGX1pk6r+pNU
JyuaUVUWD6DC+T3BFD7ckL35A9Jv9LxQaiZgrD2Cd8SgT7Y4KmbMDx8HWhcAMupA
NuG+5TpFI4Uil503cTLWQmqHsptEJKe6ATfR4pVbLjeO6Un1wzebYXfkvOVEkUNl
nxTzxiVWPPk+jSrY/s/JtlMZ8zwzu96Oe4aUOFAtQmzZvN/OM7TqNTsB+65Fxk7Q
ZVgcA4aRS6gpkCC0uXQIKMgzMcnef8ZHV6MNrlieFVwIE1FELK39ifKc8Q6c3eC7
OAcvjlYtzscEiLqgdCxzWCFgC8clOww83TLAdND88Q3WzKLx0/7VDuCg4EHPR6k/
snmdpZg9gEc62LWt39bal+0XCsCivdCcIzaCNHRuhOcBnLHgOUkM2szuLZPH/xfz
ThBVltWtKwJxQ3ZT5XrH8a39PXVZfDz0yA5mMzZW+cfkAQd99p7ZlvdSe8naJVVd
J8m296Ylt6JK75UxBl6UBgQ02+eJJIPEmUbE1r9wLhRy1EUVqi7n2tSdOs5MSMsf
F5Ae9GSpFzuSi30yt3wWCXktGhS5aw/MHBeddjhsHSTxrEgtIHbmxary8vNyq33v
7X0KG3+EdfL5Sv1qUkXhIQ8QoOigioQd72FDMiRuolq1mMMaQ2uSqzI3Ieu9WeQ8
+REt07cZZZDg93q8YW1N7olH7eQKpM3jdZcCoEVnyktBgXVZIe2IPJWCkaIWf882
dQJ9KYiUC+GBt1xrEBojPX2sBgG6dRgBAP646dbDG5OSNYdL/269IIwbRgcUuqQ1
y3ZJXiBvD8pO44YVWaRpFkESCNr9caMww2CNOpDbOZpL0T57fPsyDie04YDOB5sh
1hj5zSz8ny783YqqoJN4D7bcrTs4wE5GeYzEBzUu0gVEkRIV1YkRBJ2WD+o4nk6p
zMEjlhaPp5W7rRQSsAAjw4Z0xjzFLE/Iue9m85SE8uCHbIpqc5nN5F75ww6lQeg+
A3dKp6l6JrxQeCNe2/9ubbpMT55cfIgfAo/fWy71l9wyLJNFSjUYjbPn2vVJfKhm
UoQQY9bZFpTFY0xCsgfcfenAzk/YWEjHWTrC6XojDNlFkYjrmXEEtfwmvtutdm6G
5m1RPJ4wbOBoRbR9YLLxVfMnHz190T4H047kMAQ3CcQFMPBue/DSRNkr6K4V09uq
R5tY1d9MnzzFG1eD8Q940TiwPuftu/zaSwbD3lnFD/UzNLGEnNNbzY0y8erK4L17
aFPvepABWaKygitQrG4iQ8NkK7wyCAyAdxbSjAmF4bgNxa1yc88JuL+VKLZDgHQr
XvVDfS8WgH5M8UFvYEc0DnqfyEyAZl4u72PBN6mmbAONn7E/NDfL1Mg/PD39Vg7d
kv0E7jJquBOXICXcNK9TU/g66TcVnzRmHodm70tNAuMjNBExjXeIaZC0h8KCyas6
hRE59MMQp9PRmy9qBhT7jZC8FNLZ3HQNmH3RNcjigtteyh6ognpewIc9cVST+k3b
jgmw7PYiQ6XeN3wdejnLeshpEQ6BDeuNG5VlwuPltpQVOZWngWIannIyS62pJD/9
IIcFZsDaSMdB9FcpUZYc9T1lcqvZKNuzlAepV/EIRKI/Mgn4Kr+C2e/JwZEQVJeH
85On8EtwOclFzN141zRtNExzhJDoFbBhMMehfeIe1kvUoZKY2NK9/EWw/DRdCHsN
vUiG5fm3PVVgRCoJxhcbzusxhcaDuIikUUGeix7mIvgvfPLsYSA7NtJcEh7HtCSX
2sStVrC8NjPPIx+YisQjzMFF0nKn4ERtGxyZ3sU8RuI6CMnqj5Kok2yRaBGc2dWa
0jRkFPK5H0xukaRepU/UiwJPw9eYDL9chmxW/KEBU/Gc1DP89ZXoDHyq60I8ByVJ
Ml9GQD7grNN9VnVoQxgQGbI3Lv/95WqdTwNcRnMTLft9ZgHFzBuwocHEZi4j1xvP
+34geP5F+KwBiNlZ9nBVdK4z+Uw+blryrNqyOUb4qUjNAapCeJujpe1EtwJGikJ6
16vdymOcvxjI3BEWI4RWf6zPH0DwMaeFiZ/eyjeFPUB2BgolrOAFFFFbfQW3dsED
2LTc5g+CW5/p/raMrsezLPFq6hvmt2bz4kq9DgwnRHnCUc0EIi00RmngnsZcIL4X
KnTeT4AS7VG4v/PoOZHMIVzfWnfNZqJU1KBo1yhGwC4+ttrPdVUB3XBonGJX7aaZ
8DN+klG9XI8XrILzBuw9r6Rj1S4mE4+uOVGTQpWXIJd7C9eNqEefo8oikeJSQJhH
yB5Ui6iFn1TGNrMymnttpuoZMjdu6eXQPKWHyzprCJI1h5NenqSWXOuaZ5YpzCmA
eYU550gYFFgXC9NkBs5ry43m1WS9g2vhUZhIsPNQL+iwhw35aZblxvNLzqwrD87q
jmIqAC7gB0XmuDNnU6ceVytqyyXzrZ8ejvBLWcjXRlXySpKXFxKqDVCa/7JyoqYl
jPHx8G1b/67vl4Q/If7S5j2WBw3OY7nmNysu0NCbbgcmtpnhK5SgA5andpM8CHJG
Ac8kMPsBCjW5GfAp3cZktnS6KXJcnTW4nNiGZogPRZVEnkolmb62wyr79uk2D/tN
vw0X/mXLFE4GCOSAQ9y64T7GjVbumPPdoHHatfRIyzoD3ks4XvncZTAVWfVj6QfX
x/5E7dolg7hN2gb31zkbb6XoJIdXjBKJnPU2HdXzHlrKgS239mW703zKSFAm3rWg
jfPkJBQvVSG3FUMMWFQyGRG3z2Q11GPgh93/Y68f+c+Vgf10EzD3KisxuzZpOwAR
joHOgSSrP6MYABm3b0n/4B252ldknmrybK914hRsbrAuMnLRNXOD9yiYj1ZY3DMk
fpwxT9KT0qbg7dSnk0Z9RhE7bq16wlRn5YKyhAVYtDvVGMgZm7VJjdSSGgV1Ox5k
BIfbUvGB/Mk6VoQ7mkXzfsxz9I3KHUWlVskyOhnlruQIxEnSEvzPBSxSDsBf7+di
KAWFA+A6+AwMdBwi/SMeSQI76DBAStUWvLxYCTFdJuGZtV0sUxx7ay9zxdn8a6Eb
qHPl3G3ksYXABQgCqfOkPPlamMQnYY/BMBWdqRbFWeA5dF8l8zunXrnOC+tSVCjc
Lv0rlnA44Qay6yQMOPCYHbjca1hM+hWINfv0Jss2ZLaqk1Q60gRZhqbTP+yUoOR1
5/KScW4auvFkqY3/0vhN/hYHd09gWY750fYSQ0pKqS0Jli9yqIWTeqDhNDDVepkd
aVvmfg/llfS6vW1Hj71RjL/2qYVs/Yd9kJjopc49uET2et/xKYKMNrbXIx6Ge4WQ
YBwvFi7r3Tg03kLM6wXAFjg0x5jk/EP8GI9DBm8mO33dG5LjzPNFh9R5k2QeYFXJ
S6U0KZaK8K5Tl3YGCA5tQAAXiqortuVOoX92VzQAhSXrjNBSbTdgN8jxUkAAsT7k
G2zFPvDuhpaThjM3SxYxD0MVlDiWZVsoQa4RD5mhbbgKyKxcrcmuU18ZPORjdzVy
irEVUoTFznUn04wYLibxM6+7wHWPLUGYzbH/7kjlSAiS+yp97BGHjUHf5kXHSeAZ
ACK/Ar9NA+Is6QmuK6KE/ZywzenMspts9nADVggUpgTrfqyZBy3LfSW4zTt+IWyp
rKhOkQEK+wUdyGXdJXokrLQxdKEu9heWQ8sUBnhNxO64YBjAU5AS1c7rsKPXsHjT
kmGE7qeEyuiFLwPNz/7py+ww0FWBWZSnGrkQPBLUeG2PCtf+LwqaEcEQp+jOqlhI
1Z6bfWadKWtJH7uzNYUWCXvIUrBg9IBFBmGKtpFQ+fkKM2ox00I6TC/hqqvxuA+S
G7OkpNOyvXfuyrr5fAAInRGtD4riIdoLDUNhuBEobV3LO9IwEtSSngiVopWb+vqr
FzMkx3dG8Z3cqst+/vfcx+vo7vdz37w+/idta2LfIXU+j5zigx1oVkrVnLYhZ4Ph
RvVcKu1e24QuUkHAxVEH0B7ijzYrWW++8iMlR0l5hj84pwozlgjUa5Em442DVFxR
XmPQDaED3tgt3RiZmanNuul1/U1igSg3zQpc4R4PDxMzicTdjoW0kH+r4CHdDdJc
mmzX+7rK1mpNWZbZNwmMW9NGLgU1ntXspPV8yAYwVl7K7xYLdNe49gqpoWTEszy7
P9cep1uEf8DEDQZ1O8VRswCiCYKqRb8uikfUQH8W4S3PbWEbTN63focr5wOrOjTm
a+MxrD0aU6MXDNh6v3V6zYXili/QaDebcyT7xfwpFOZB5ymVs9C4hMkm+RuIf2FT
buLZvF54ryGanr42IGljuMaushH6oIUYIifc0lvLbDjzNfTHBsVkCydPKoaW+vUz
p9/2p0Gw7cm1MEyOZpHfgxxYbx3Z+U0bCiCrVKtozTL18m/OAWKx/A6mT3epUROQ
rVoXvPUUf9S+GVLffHTY9tE9dDI7rnHi8Q3z2sxLNzDWlNNtc1xLKnDnXKLHoY/D
n4B/S2d4G4hAudG+cBjmxa2xzHkfWJzMVOrE7a9g3vgYX48BzVTuE51uHUFKQZhi
3s3/MNWKWmlHg+3ufw6kdzkZfjAKbfigMoveKRfa1pLuexu3IlD7JaQvaPN/gi/g
r3cfIXwpDCRZ6XOwwqy3Rh4uJaWPdj5QcQlhcnmZJWududZZ56EewSoJDlkFPtzC
cm2g5zeGLewExN/c8kLNsZTd2/CEp6z0AK+fSboX3MW5nKYwx5p4hjwlZ4CZ1A7k
xvtImCHY0YTDRsRNK54DjCLcisMejdDhUO4Hn0x6+DPGoKfIP7MMVLUkZVLcrYKO
AzNZJ1UHQJAjHfcHFKrqnxIL/yoAUaA/3SfUsQKz/u1sZqpLS81WQsA7eV1T1HLT
FUFZ9vDz0rmYJhlrM+fMKY4DDzVeTeCWnc+YURS4tckZDxjlEG0scgkv1+3nag8y
JIKaAIUkw5QWunJrZBUQVBPSzAa/ODwbt06uXPEWMelm5wps7w2JYSZyRqKwiN2S
3JuYcFeKVAGz/WWJT5Erf+hTWmKX4i/E02WfX/rCNusAbZOE6fd5aDdSkueFlpGM
0onmGjLzOPx/xH7ESa2ZOFBGKoICxq5T7AJsC8bkYRkb+ELDSNr4E8IvS3Kf5Spg
5b+HrItS/s1w6ucpuuGNM2i7tbaqrZBrsivCQ4DHl8XLxI0rg6wG7+fzXgfWzT6J
tci/dR5WtNI7wOhkZOM/CP7B2JeOF0K5v4akVf+ibqsCKTYTmTh99O0dqdwDeP6d
L+Tkl7lKqBC2yNN4fKw25NFA8ekOi19xq21to0DGgPZs4M/+vj/SgEpel04KsrVe
TM5qo9cyryfKjpup6HpnRrNmgzxGqmUIyp/tUWDs0gwV9OZN0r68RmyQl1Tu2f6t
rlxr4dE7iXK1zS+Cx0iUbVTCpX45DySFLNUKs8fjGvnvqbiQ3fIGF5pQ2H79M31x
2zeQkgSxnykdk82BhTGGDg0+TrX82gM+g+VicVBrio5Mmiwpf0VReZK3bLiz0BRB
iHGdSBSQRCyDyqVwyTVRCKDrzhIGG4+itSTz02Ihrh+i5p8zKmkbhHtVuaBaTccs
D7jVLYm96YiBL5ITeXny5WeCoZ7UaaH+RHAOCUNqt9KHUayW3ais+tZ+QDEbYyq3
2ljVYvwAmy14HG8mF7puflbwzK4sTqRaWlZG8HX8h+5L2LbA20rAsCXoj5oEgP6U
ode3HIXAK8ifrt+bF/ay0JW2vLg2FA7kEiFwCrJORz7jYc5q+Gbk6QW0ZBJlRZRq
GpsaioxCQ4LrXXSN/pyRi5JBMQCXaVm1tDkHxryhPTHL7IdeXthO5Mz73uvqZJbr
lVaNnqFnooZCBQ5ueS3mMVkHJNMG4CFqLLvxIrt8lsJyTNTs/RANUA/0oHoBXEVY
ltyBwslkE29wZl9vGD3E55NNz4TXlrTvNwyNIKO3iD/wjbUmyHuLcU8JaN6TVGPP
OjKEDTF1eWpEFmnWu9fGhkdlviU/a9XhVrInB9C9rRKgQMmsLLRsMMAYDpAi9hrL
LzzeX9s/AQBdexA3NLLRvvJp6R3wAzbXEn4p9PbQQjiTFhkmkwoi+9TohgfLAm4G
6a9+Z3pskg9B57VCdBkH8jQ4JKDWkwPNcKyYRFeIrAwX9zrfvA8VeZoUOigyF+nF
/AKhhJKHmq8tBtGfJYgG/xhxWmQuKwIbiGGJATe1UngHruHjPydx0TsdvpgFI0V+
/rIv9eHGk5NYwDen2eXhGkkNN4Jpsw23Z/dRIaXY/RXu4WhAuhCj6oG4I30+bjPK
66vedONkRzlCOEm8hbxYgnOhGxZ7B7gq2CD4E2Donclq92fUXJjsjjFNfgXhVoR8
BId6Y7MFgdjgzHfPsoVeZuVYFiKITyf3Lu8kw0nJR0BhyYVbHcTvHmyRjok/4kDm
BuNnj+NqbK3iJVw7q/DbF9K+dglXNY0vbfvi7NF02KPlSMR+QkvnwEVGblzUEssG
NhxDN2WfQ3sXpS/Un6Gqc9ISh+E/b3UibT+H6OnXiq9p1IQqsXTO/FLjEIo0Vhk3
XKx4RST5MmCEkWxbyXJxG3dTZjXPxlbs+gZX19dtHUTGmbjTTiu8kXSGzGvvBHJd
WIY1VstFH6tFCz0ZE6yINW0ncPseAnAfovXheUb+iAJ4dhLVWAbDxz7dthtjjDT+
Xpyi/HSVs4VnIx4bz3f3XSi6IUSPp2yr+SAM7yX03C+DHFEtCTsIpqOFxlWwhZq2
0/fgvMkY3aAToZX8UEdxbYJfYmrKQRhT8GyXx6B0s3uHiuGfuN0d4OWUrC6hRJjz
xjjvza8BFH180XMHyga98a3Ry/KOWLuDMS9FAFwo/kUEiAOpW/pTMSbE8B6K1vjm
XLwL2+isw9WkbxiLCY+mubtMn8YHulKDYYO1F+ZEHFrkD5akgQT0uA5lQpGqkLTo
JC14coyr1BYQqSGeeQ3rMQR2QDzlyRn9l7Ooe9keMt8GU4goE3G2LwwLkNIzOlNE
0bhuKdelTO9wmfrKXguLXsAQsT1K616GP1j8FHu3G3jddR3/DC+hP6ex1EO47yXu
WrGMZJqvfvl4HHwVkkbOcQY6DHknFZElsbvsT9DnrZxNOQeGpVmLCdQoFE5oWf7X
Ng3/WC/4FiQxUJt9Z/fNKQ3qU2JFZXzvYiKMjNBB2xwMj7Hj33vEso6NYAiGvG7z
FH8i07kERwGkSwGMowfsw4ngQIV1DNEW5ZFbC6EUYtCrvYA3dHaup2yamcTKWdxx
RdplqLasGmfcRBSuriNETXXpUUWcXhFH5alKhM7ckDzoupc5Ngepugn0ZupF0pqK
qvN8FS4naZ2rLt7r0zyDOSE5/Wkx4XHUhqrb1bXMdsASzxIWcf3p+sM9uRFTHUUb
2X2KsFKQ+AH6pxR8Bb3NBa4015ontuN+0/2/77amkeEUEV/VeWWZnbI6yHhokDjP
7XSfZmQChAgw9JMewnAxYTRapILfSIS53Bpdz6Td76Na5kMZ4cYBy6TqJ+zo7aFY
L3vf1JT02VQ2sF/j3UVUV5FMkozxdhDBT9vOErrLY9qcl9m+XVf5baRE5alVw5GT
rUTsMCGdecxDgyPVY0a/sgq1f7TXkOS884bRrv/CJki/kYdzGL1qUYAbtRBDZ99x
jtQcIWnhbUyqFr+ZSJtZLFGGuFs4B9JjgsMRMZbvapxcV6603/OixhvzH/un3JUu
Ad/YCRgmkeX6uUrCgAP2tR0tq3UM1VX8LooSclX4000Skt/Ah1J875qsmghP1bLT
6Ykn0we2skjzW0aoqK+tDGxqGlPSYBVWZh6X6xFmbJIr/erknkGrOE57rN4YQdE2
OPudzzPLgxQDc/I/eR12/R8qPNZ/BeXU+EorxGX5mzDekuKTdn6k1g+/UuFX+o1q
CksZSFNnV+DjtB94QTaq8WmtRBjvVdV14AxEL2EgWLGxL5T6qRt+sMuILWhQzGFa
ntbsuDo9jddWeGoK8kVUsIVvxshN94CLAtn+GugIYL3CtDXLNWa5MfMeEV0HM9mi
HsObEHTp/3PaaSgk1GQoCNzw994A+emQlvpfLz7KjVi58KoLv3mECHXi4d3AHCnM
t2/XDkJtFwanLWFw0BQ8DVFewQ1lwnR6wnOHXsUkA2PZxu4I8rO2SaF++AFK7Z1D
lQ9ibPMt4isVxDEyZf5dtx3tVnY4wZ5cDFMGgRnTA+Duut3VtcE9Bh6uAlA76BlA
GzAfJkXdPjZCScl74IVeXFBUI16eqOikYkTNl5h6ovo891Yawn58GMNXm5/WKcA8
VJlGXrMfSaX4CXHrlN/c6c8QnR4o3THDaqWqgp4ZrDN0hT3zQmdWqzcsQSWLYk1j
8cB8zw+5LMcpYIpG4sL/tKxdDo2VxVnAW1QGwWUK7+ItOAXAIEy1vLjsEgWwu7Wk
pwQDllhD1WulEzZGEztPZkmrLQXE2Lq/OUpkqB3rv6V8xc3G/bz40aYlDB+jfyGc
9c/oE4UeXj3uf3LMbnKJdNxtgCiK2G0v0yDpUIL/yNBuLtsZQ4ZxLN707E/8Uhs+
iQGpdOyxwALlCf8cB+MlBOrXxxYT0JdEE0XtJ3scm/ySQ9VBGnWO/oUeyc19i92h
QuriySgR5yZpB0EbVr+w3ZOE60wwCpln+gx/NqIwilnO7m78Lxhk4c4rHUoi/XlU
MLy/w7KQNQVVRQqqOokPDtrBP1945ZHKE1JrFBNIyIP8MbQb54OCJzvWIIaHtilk
yoVGVGCiredIwYE00cMozpe7RhnneT0ejjKWDuieOY/5yq79gm5Y1yoLkXYGDv1U
au7r9zm3L7DqLTO9XhFIGYKm0bWzkRod4BWc5LLlTpx1s/OfCCfaM4mqXa+9G+7y
5IITzOVTVpXy/N+y0xWvi2/rGGJ/wosB4PkxVQn86H9DmMs24zBAi434TpiGabOR
W6XWzPaZXu8WgBIgUvg/1NHfA8MBzBWdEenhU0WGE+sRCv5cmk79L/qpPNRBXwk6
Fc6x1b/ElCH4in86tKYbKLe4qgd6szolvhCaQEnN9++d3p4B6ib1A5NIbyIPtAYe
nk0EjShpUmTWjZH1y9FaRPqIzaBqOLe5YETsp51+OZ2C2yZgZRJzQgQb7m3onkGn
PidgYneWjnlQWan9n6DixtktDK0/ZK7Qeax32ZCO9A/mGbn5KtjQBe4lMrKTym5G
PptTrF6lulrK5AwBTpvbrsWSrUnVekPAuRgxvJa+fzzlKMkb1JrUafCk69UN9zJi
jYTwY1OD1fQ7JhJeFTRJHNDiKI78Od3qDTg4kz5lp0zUqb7uHwqrTYBfiefBHHwW
sQ1NiOcvVreyRyIBr5ydZVxqJ/koABXNn2kY4AwxeMpp0ZgYqMdn8K+svXDzb35N
hfJbCQXDq2djx+50vt7GuWyGeqSvRxPSd/jTexJSnPkBDqMcl4qP8dfsz1ZRfWq0
cJnEkXI1IclGuHOd+rJEQYPI+0oLtAxRLuB4/Xka/dVCo3UM7E/ZUnICiQhvGFiW
GKfj/VSRdSYO6xEg6QiY2bi3xNmogOiSYoNEiHFiGrceOwPA1mKW6OvSIVSkUynL
heG0eBvEAj+J1pJlLCt1cVR6l0YLfb3dCSowmmBbNri6qmk+/p40d7Wt2ts+HM/Y
e4hPCOAkqfvTFdEFRwgsoJ5OEPPXwUmB6YuCY5DOrDmH2lzcjCNtQfiPJD4ReUcD
5vZ80h78GNg66Nq9NEp0n8vMIp7R0cFFqhLT4FM9EL7K3kvQCL0caeHr4S2Aml0x
pmlSSb4gLzO6clnKJyfEJk+JUUcSQ1ncLXtZ24Bv3ejBNYn9U3UEYa8QmffsBa4t
A1tS6SWmKVCb9qctToAHwLi0EZqhKM+wo2qxAMlY2Hfz4uoaUXdJqyLxMnuHrlWW
H56fGpj/4wpmD/mAEi7y3RuvqfMzGjQWVywx0zwUbnLwW5wZ2Mos0wnwMx8KEeL2
fg1ySjLvLzLtubCA2aa+3GC17fQk/So7/nIUNHVBy8QPVkQE4JXEPnUQi8RRu6bc
A7a7qpjFql9X1B80pVXTbVrCyfOyCYx/UcB82cijbcNkQ2odawAR5GOIy4/HDJdk
ilK0km68csCCV++h+br7exhzqsZAeb4jptNUDdjNX76qAdoW5/AcmN21MvJbsHby
CqcsYaubsHIHkaBDxJsg99P5ihH3b58yj24uyiXkw8p91BEBXd2nAULfvkf6Bx/3
F5CfqUqnyrFFxehaRPn7k6/MnVL90U9ri2XA2bNw/doGE14SFZZz8HRZ4+QtESBk
AeRK9Y2QzQjBuPsZlmuGnaE2VaBnjS2GP9orP+7SHvoAOeVGbTMQQC6Q4CTs/tWN
kZtAbcQfoRK+zDqvJFyDXsM0TRZ8R61OiZNzrzuDpgQE81Cd+ETbaER0tb4CnbbX
JH5ZNAsQXkiW5YrFIUfLDkIR6S9iDKZhJ5740XT4U0z68kP7E5uoUnvG1dqO28Ay
6JHxeLEfgiQ9ZckDCBebFA6zPrNoXyCGXl7zbxIurVk769e+bXKATi4dndbSv4Rd
XafHH+xuKrDIyBwUetHDGmFj748iPYLAhvNwMFz8t8gZ22iZwPz5Ajq6aRU+6+jY
Dqp4ooD76+cvnUYkyumpM6+nWgnYKbTiQaDcxE3DukyEcr3rXl9adHvidUna30/2
ft462PLZ6eFhWnbhsa0bVsrVpbV7o3akOGML63vlNwYkI/ONmoEMFz4eNAkihFCV
yjxARUULtBAO5q4qbEW1Z8JMfzMOBttQNduPTxH1kq9/zZm6nMwQfs23z8MB2LKv
2JUU1XcueXqtCaS8wow1QoK3B64lAr60fPqA5crZKiqjCUdFsXCt5rAV6rlE2cCY
yJ+4vrauTnf2ec0hQNpIZgsqBN9nIfp3NR3Xc10Ky8Fqtl3rDQqNOntm/YuXXNqs
yqUkUTgflwjaOS0Bhp8XgZYlceEbWiPbx60CasfN6g7He1Y6tG4pE55tXWl/a3kB
VKlY4Y/t9KG3+BAg/pP8TRNftTpDWBBGJlvJo8A+Iz3JVb6UtaZbgsLxnd6/VcrL
bpqECPlud6YP8DzP0lgoaX1A6Lk0rOTP/JmSlp7F9zfizNHVR191HZNzfSWf/Fue
NlwqiV8sLCodYHt/YKrzqipH7wZ9WbJCDjLodnETJPE8/hHmFvd1+qXVvNn2d2OQ
EQmXU2TMpmalM63dNSrI3dVdfNZZIo/UCycbS4sDTZuRVKccDR+r9l/xV9cE4PDU
OzntzTWpMWDrISUs1vl9Z0GCz+T76Xnqfyevug2LTJaB4f8ExrC1oAmv+B3rwrvM
NumFFIJRP28yOy47EM5FCWIqB0SCI1cOQYcPQq8bxNu5moaYOsLZD4l7AE3R/q5y
RlTLDeofPx2Z0tJoG++gNKmNRqpduDo39rda/OHRD532vHfPoiVoIdn9TkETc0Wx
CMjiSGDIhG+u3apTpfuoHFwF9bckrJYw9JFdOMVcXN77EbsXKYV5LLfxWgP6GiwN
4bhuxCKnuPHAX2aCWxgWt6vM9upb31ryurBhKgKq4KmMgo6fkILhEA0H1oJxvNkD
DOsHf8c8HByf5hrHxYPJGSXN0pmfwAoCkanrOcodjh80iWDBYIgzPCg+clf6wCou
lB9tkr7uIle9xob1zsdwJ7x7Fjk3pzjCExuZ7W5KL3Xnrd6wj0R5FJ8C2BWWQMdP
2GHaocyPqT6M81OO52O149yC3YaDn7DwHX4lPO3Ip4pozXcCfCaadoBjp0CGg4vd
WZMIwnK5tNJqRyqYeqdR27hAlin5ux7ZFBOwKhvIvtbMMEauscjm9qmjvo0/Gwf3
4zqQ0zf62YxNka3H1lbJ5nFd0RjFvi0XV1meQ1p7f8wrfpg1RTJsl3zGO15NRIN6
aES6/yTSSQj9K+Wk0xbopAlOTAIrenHlUSQfj4fKGeUOneKqUzWM0Ze/c4TWORSr
a2WI0M8iFXoOTujRkp8d71xy6P5fnQPrPOWpwMm/lsjV++5lmMp7F60bHRJBrRTA
rEzej06gPZZ87iJ55DVc/Gk+CYT/M3K1ksppnlS1bsBw1iRpNId893QHNBTI94a+
u/747ZqYrIM/Kk4urngyGGwzjWU2Df0rXTTR1iMwtZ5G5mrhK0rqhZyIOeXgsL7N
cV5YMf/F7q1sWKEurrhg9zq6K288Shq3oL5urSYoyfHFyEW+VuR8ENxYsTMGLYiI
nDcLsI+nRRYB6EdUvINqAgt6d/fkBSQH9uXxPTTVXqP6+trwGYIBQ3btA67bEReR
WlImx/qjIt6M6TIPTkcu4/M1aQc3Td5dHKh6FiM+Nc5OmpY28N3t67Kb6zZ5+DpD
2cVgmHQv/zW8RW0WSDwgk5UJhI/X/hjZBsuRxM9ivgmTdBj6EBE/MjyS+TAKs/p2
8yk11CGldwemjy+EeffSylk930BUGwoxuf9Z58DKdTyc2U5JAsVme9q+xgAdmuy4
EtNrfmNWMYWeY+h8Q44NVGoCqInsULt7YnBPd1OQuYztXS4tsVAfIBhvFSe7TB6p
rz78C8Y6d2ITJJqmipvfe1ogV0qlJdjGMcAX2iYbcfY3cPFxhYscKD0gZQlb/Qbd
Z+K9EKPaTacRIuS33xUnhd6UI4UFi3fQfmq8jB5KVDwU5xGNjeinPro3xvchl9yP
JdKolTVv+0UbKssFNACOyXs9H4b2bdCrNnvqXTBA7LCBwyHMrQ/1a2rONNEdXezY
s9MzcZHktk4JeBD71Kc63hC1b3SZXTiqAaLcEwC9VVoYSRhaegj3Qvpe2GRBOgy8
CfEGBhfltr+oeeNPmPO711ipsTGWfowXpM69QiwO0LXAx5kysAZzpkqyFaF378gI
bkIZ8K1RbOjxtkyFdEwFfhM8WxRPlmUC/F6Qrg6l5lNo6LaXETwtZnFkUdJ5ytG+
yqAu+ta1rr98NTcnkKS8Xiy3DYXhwx7GX3gOT64ugvrgMJubcVjvDeDB46qHx/Uv
LgeKikYdWcu/HuM8kr11t+J7iwI9zidI+QSG3CfJLviwc9ERxYQ+3r1KUe/qxAgt
y2yLqfIX9veOjwTp2HczBI1DsDZ3XavmGmCXbjUCbgmHMgwo8/eGgUcxeEFNH5vk
Dse5oToWmPnzvChuZAxI6S8Z6GLiO9ihpMQP2vgHCt5XMRD1ek+o1zW4WW8aJ6m0
LatlqAvgklfQj+LlJBPpbYxvDpRh+MA1c9PxCvOPP1cZ8UgKHYr+I+lqJvZA+h2i
QR3ma5hyEAGhwnCfBjxczDypFoFPn3R7er47QqkwkQ9xzO3H7CfKgTJYBpN2p7EI
ABkFd1NK5WXDDix2SnFzbDLETY7jyXQrv40c2kfwSYKmGd4j7v1RKS/KleyW/OuF
kG8hTbn4G5BzQ7uSoPL5w2+ErUf9Z3SRFT5izgou/eT1eY6KJlTywKy9Ci8ACL9L
2y/oAdReAkL9aHq87THDRIsDW3MRnGWknewiWnOzATHYBLB90jlPpoZNSfRtQN54
hRO4Mmi0Duqeq4j9x9p9iQ+d8a4cpjm7YD5L7j6h20BXRYPYaGkXkBtxlRBK80+6
f67ED85RZpIZoneZtFQ2+bWR2lk4Agl0BItHFsp1N4DX0gcwUBqyqGcZ4EoJRxqL
3okIodDic4i8ZWiYeyoELEXgr1T0kjlReY2+6rDBt+qhmnsR4rdksDSou5kWyFdB
pn7pbKsqzbjxRB9fA1RNB2s0nWyQgNKsPZAY7XUOvD58s9FaAqoIFofiEMkZVHp4
dBNsw7bN34wPqD4OnBucVqt4HFrEi9SzBPhzyrSVg2k6uGlr1JpCRuT4ogzCB3Pb
k/h8HAFfZDS1dNuMCYJRJO5JPaeUuObIdIg1YTVOogPliM9/i7vC3al0mI/q4k0N
M4/5q6R69pVzkE+dBrWNiPpofy84uIe4U+DIg25UTrVEG8O4ggM7S6mps5W9is9L
iESm+K6G509altLwJJAImsy3Q99cjkipxs6j16uvafBOgwZHSaqCC2soiFkKk7nU
b/G+tBaT1ENjxkJXmSaLjgtvP7S3Yk25waFSx5L5IcsrJLf+0PjnSHf6SxORVcz2
DKodH/ptBx5zlkY0ZN+gJzp9zK+yY297C8eljH3Scqdz5t5GEHNQDR7/6KnJCzVw
eJlKMkLMD3tEcyzrJCe5Dh3OG8f8UQ0xUIu1TIy+JtT9rnwi7e5rxBCQHRLiptk6
jPB9YIrXRNMlmEnZ1ks4iDaSd3eDONoFVuhHvs0d9Gt5E2+o88y4y9swzZeZRilS
G3A6EW8m4IhPWTxsh3PHwqRE5jzzHVD5G9OSHpMcGxof0hRBQNqBx6j5sEp+NpQg
WdRZTBQ/neTPjMOA3vgbS9malV4JgXgIFC734/2o3834tDfMEqSpw684NNBRUy7K
DuDqmRC65LwFBUffVBX6v9ibEeZEpX//+LDm9KSTQlzxZulLoL211K9ZT5mN6GWY
40p2Sv2r9Kb/CrsbTEJYFncZaN9xXPTfEpmWge8E0SfqYZbhzw0JwUYaz5RpCQb/
0qc53fRY4sgZbTVhiniXuv0PMfgyWcAGUt/GQMObNRHTHi3Pf6yewuMiNXJq+zso
agtV1v5IFtXjyWMOxkWUFnc1aBo7yhe2CSo5edZ+dD/8Wj+WLfT3Tk4e3SvVEatb
zQcMZBo3rmAn+ACW3yoag+Kx0qGS+2/xFGGBMbnkeEJQTQ/vDj8hW3RkTt+ZoAg8
ZADZokp1y0ERASGKMN281fbmdsw/6tShjyl5SC68pcPyd/VyJK+itUDWuFdQkoSU
yWRFxUWaZQfTOC4j5xZBaDJ0ma0zQKNa+utdOH/kTfQfQUR05her8CPOFeYzIzta
jgAdNOkZb+aU+s2NjpOkCqxvaeIxuxFNwqvfW94acKbPRzo2jX6LhsnYtONCAG8L
PRpB1BMBcy69DpEIa/ZsPxK/cfM5+LxJggh1WdGzP4HkMOv3uB/zt9Ou8YqKteQy
LlT6WW6hZdYfHmCHhwifMb1e1FDER3VYpUoEODX8wneRwxl40G06XexfsKUAwc7Z
/3tj+IG4ekY3XEn/YbOD9nDJXi8e6RMTG0qTbl1SClUXzYtRyQsXQ9rI5R3sna30
pbK2oYInx+FUZnxFYFNHZ/92y9vlV97RBsDieawGRZNkdu1wVmw32sYj7o098aE2
4F8BoemLAXgEQZd5PEyV2Lva5MReeNoTWTziywLQvu2cp0LvK0POe98NhY+YZdM7
g/SsKKBA6Q1eBNVSJ/PjQ3HqEZp0ZtvsrIGkvQKCUYlMmZ24+7krrrXSVYX2mHdL
XtfnWz5viJDlY1AtNc3LRFKmMfgr97qzkUUpAC7GRf0GmsfQ8DPSB+Aogen1nHBT
JzjBHzKZ6LzSY8765IG1CfnOC0Y7x+pj8JKkro/EbcjiobvTvMVM2HfSZ1Qb58TQ
D8VMcTd1nm2PEuBGPeroxRWbGpsRFSu4E9kxeW4sQk62xWEklf0ViQjZFQbwHUsi
o5aOedFQU/J3iqFbscbjEo/OKnWmi/Jp2k+Zn1KkDE5medy+FxK4wGnyVCRFVKnu
ce4jkagTkXgRcHOf2TZLITnpCl3jwQo31Jt4XOn0pG6o0hBFkC5j0z+qmqYqqaxB
cYEC0U6uFqUafA34p+jJwfwYMKVsPGDC5xpEKdFyWNYbVqAEKAmteFKfE6NAVwuX
3m4BMxsusS/xoTHfIBDbkDtMUdpdArH9/pXWwIRGvlSaS5R1hFX6+R+LlU2/Oxe7
g1tAYJhqGb21bBwFvMgLF8a3LgeA6MRDWoqiC3p4IUbCxyMiczFUsPxJbCe/oA9P
tI9pNzB9UwXptMUE8/nmrKVV6vg1AochA5hs5zfXGzJs+u5meT/Ho3XM/iJ4Rrmh
fGLJD+Ofn0RF7kSZ9CPtr/ClvlVvwZNg2u6Nshq2N/Zj2zT8nGBGs0ILoGR7tJoR
G+P3F0BQdhhlQuRDvYJ9A4iEk3VHEqwKVNh7qKLWOF+bOQGbYP1DVuH1YIoxmY54
Vv+3GYBDExu0Gh7BtpSbhkmuXbPleMMeFJ4oaAT0rZgTikz3/s0/5ScrmxjIFMAq
K6CMHth5mignhfk5KRqGqNIQPA6yqSOkFnNv+6yOs9/YUNqs1OoRq+ehAQVgy2Iq
VCutj5o0kU/pbJKklpS007VdGhv/7jyvKaNGfhc8TKC0sFdU6oo2V52ZJL8Vk6Op
IN+hcoFP9J7EMS0ES9Zlhv1QU0lv+3KJBf1ux/lhKg+xJA/PC8p2W16KrfYH3v7t
xiE1aos7fWtemANAozn+e4iiF25IRXigRPSxjRCDCmkwHMuQ+04hTH7Os2RufKCI
hdsVsZIaIcDGUKVMTp2JTNFaz0hdV30bc6v4l6R8JyNSmK8qM3j9w6QWhOn3btBO
+ricO2ihadg2zsBgmaIGs0/kQFq2mZ5lFiBtD8gbjx1HjTGr5oVwbX2k5JuBo3/Y
sIlQ0TagMoTZ6ha5fzkry0W14TgwYa/4PWQujG74tYyI7UZ2OV+xaI54Ez1vSh1W
dtADVZDkXFBOUTxhPvRnAHJpgy8buN+WSjide7bRunN9jXnmQPOQ9XhwdFji9fBR
6XcT3e8pihJ0ax/cKvGyFxB4+NOvJCuQKjodlNy1deRPhMnl4wsdyPuegLqsHYoT
Xp/WHz7CgyTqB1ovkKkeEd9Bdfg6KUV6f+s8BUETE2oKx/xVWlIkUHPcRWom1V5Y
XXEMRzA87s+bKas3b9orPZfLuW0KA/lQGsQWmj8eGoNJ/1yaGeL+6v0yfXwRf5Wp
AVCCRPHa2nTBd0Uyp1sdl3Hz6GZ1oNG+tEaB1nYjNy4mlIEY6J57FL5fVh+ExQtx
wOliZrOFe0otPPwN+G/zrgDCF8BqFWiqNalaWHRli0rxStelwEO8EF24hfTebw8+
y2kcTDC4bwAHt7dfleqaBWAtm61VkxaWfDmZ1hD4/HX+gn5RZFiRb0uoPv8TXufc
TthRj2S0CYpLBNwCn46Ue32KsdFh5Vf64JgNnWrJbPCX/vu7oYLzTZb1mjlqHefb
oZbHpc/dZtYf3kVQMDri1rZi1uC2WSoWRrhg0ZZKqIazz6zU3FUOtDP89ndUZona
Eh0K4Qct70G0vJWRQuqqCCNz/7pS3a4Y5U5CcATKNEnEokKIga85C5Kb4CFr9FhO
U5fPAjZMhQ3WFZQOLPXNtUxMq38kEWhQ6/JfVUQdZ7O18G6LPbooQ8LhPGQBsOaO
k/DhsjwPr7SvEON+6AMULjvnOYvtVYH6tkIJjC5Cckg5Guvye4tcvdLpBllii/Ta
e24XckaS9j1zawt2f27TzNF0ABWpwNWFDAyGlrAhAd7AzzF+SrGv/JPWzBNzCm5Z
k1JgMOS+dE+xXn4eSt/CzFsSlf4Za4EL9wfk073dkASrl1UsYlO57hfhk4G1B0nu
WuChpQaYg6jfErOn/XW/9y0rOFOypg7kotk9MYZaJVMcM0835EyRGTU+LLJOn1CL
zROUiUOWpFkYRbsoCpMu7JAcUUCbB/mbwwZ4rMBf7WhGOoy9IJZDXMnTKX/a2DiL
8sl24l+HZcJ2qK1BoMugfoGSJuEq3WM65ewHAXi4ENM/+lCTH+VTrsXFSAcqzedK
ohgwexxmQHProlYSXki7hNlwCkUm9AgRYQU6FDgGQV1hQ2vF8dg1vHZMye5n5MlF
WGoTKKMzT187QKVFe0rwqOOwuMjm40UgbC0x66Ucli/glrYtccKWQQ4KUOtrmufo
skibaooSsd2XF+Sfo0ukTeXQXs4GoTyHjsM2cp84Akjo53jJGo+G8TzV292uWyAG
Mlqmmc4dvwLxku6uQ4m9VjYl0T2dT8Egx6l+GJztPRo/xJNcmGWUxWOHSYhBMAfO
B9jMvtHTitS0HpxoPW6Z5I/UgiQkS9WczK2tXKynGvJWXdE6fFWVKmWwwY8GCdgU
ujrNoOwZg9gH/HQtR2hhU+yyWdCucFqm+TpRIeUwxxHGzk/XrOHKNMx5mQ9B3cY3
ubc0zLQLYtTzQKR6Ju8oa3GaaLGcOrZRNHN/0hJYWplcVPylaml35YacZz2OubRA
7F1T39gFHa18PqYe2zRjNPE2Offux2h7m6LekdSgfNFTft6iHMTK/I074/4wRmzK
wx3VbO1nDWSasTeYz0x6AP8CnGDPJV3FhXybjBfskE6JE8riSkagd6XZCW4oxSPf
Km5lYSYAZ3giRhe/6oEUzrN9Dmgok+t63Jg/73Td19N5HjQGPvi/lWzngShfrEn9
Sqw/Nux9/8sf6uy8PESA8WlQSqhqCr991lt5hsMMCJWYP2nRNucL4NJtIAsknpya
ox3wB/T04DBqAAubn3rmQliUrBS6kOh7RCyXQPJpToEK7yEHXRAvSUJChpg1dYlb
swfTkeWm1wlAIx2ws08SXsDpwHUWCjKJ6NKPeo7u8UVVLof4OugAJZznCKXoUDCH
u3C37lXIjoBclxRtNkOV8qrLn4bMK9scowoVbe/A8tHbamfnGlLpJUn/3Z55EeZ1
zaX4X5HE5/RzH8Ilj/3Z4CAJ0L2wBgz9HhXKoGZi7Vs8BWSfNyK9Rw+1pUGDVvxC
2Ek4XE5wijg/V9erWVaQZ8UEz7WDhWgUKdPSgaG1jcpc569H4wdPauCOa82KnhIY
jGR2aG1SnpxOee31jZUK8ji5BbaIU82f3QnFiu0fK8tIzw3vg1CtClYgXJDJrKvB
FxRaNGOPFVEIc/oIsu7N15JcoDLkSGmFWjz3esDnHd2X1V6bl6p9lBdoxwG/mXnt
q/jx30qyoRTCpF3PS5/57HQmSClv3514BCL5ONRLbrygHRvKTXRKL8BUm+yJigLc
KPPRESse67/dfCfitoGA8WHgaCWEyv/Fb/74z0J+UGI22/LBtHA1odcRMjVsiOJf
NrnQJzS26VEQ2tFBz6kK6gAZeti69J8UpIKIDB7egViKP0Y7e0fPl9bMJ25H/FAm
b0XtLia2zDdQjfRor0yFl6kqf7uoyVYliRWi5kjN0LcX7SicfRLpMwRzWn1N+ZsF
4clqmqXo1pr42dZzxHOelnscFrXhml8sWd8QUtncUxqLqaTv8NFACGbvBtRmMwvh
ypWKggQ/i0EWZflyw5w310F2crHjHvpAGniBb7pcWAljFQnjCj6nnSwm6oXmGKmh
tMvoMvs2Ji6GR+32tgrsg+TyF5k52+tvCNmookgP5L8WchRalib/vqf1IX71pnQU
eQgC7JiHXFSd0Jiablhbxc3IcjQa3hcQ/Nk4NcLBM0wJhS+nr3kdcJduQQ3wlEGQ
ngsmWfr1beQWyytW9PLyVN17bq3vIkTsk0fgXrqv2ihPoH+f5UyQp4gZaSe0fcwx
rBVXQBJK4S6nI1ge+Pwe/oq2ZxYxKWtS9EifZpTKIvpN8BLaloNGPL/g3Uj6LSgq
2o3c/j/UHz11252e9gUUFf5DLRPA3DawtD+6ndFNduY7Uin8cixbZp7wrGwQE4vO
hz+7gq6k3RP9COdjjAh4Rhqj8lNS3fy10mjFGd1wzFQratGFF4LmqoyiCy0cxrDg
xfHvns8TTt+Oa6JFYeJHDJEC7MzL7rlC18vyE8mMbpWeatNX9Kc3irzbMl5IT2o3
8hiRVMQjmkAUZLOfNp6BMKtie+wtA+3PtsGy4RDFttb0VkT+AISUVgIcCDII8EGz
GUbhFxfV2EqpT2qIYlmff+Bw8ydRJ6S24Tik0b2BC/XUk8ObCREeaU7+3ox/4PpW
Ne50jEly83iezd47XGxs4Dq7ByM1u3nQ+lBjDiyFvPRBXJ4zauLQi7B8HMZcnGAJ
n4TnzJTDNsvdXb48G0ZMuAHedbZ5v+LJIFysQQM/y3sk1x2GHJmNimsGObfMAgPz
wnHFaOXkDwn6Jz9TIfUrAWwLeozsLBGhcR/sP/BQYrLgdERFF0QlnzEku8lpbORF
KAgMEkD0mwLPsbui3Bf+MUYWCA6R7nv6bdC+GsZgfovzvXgD4AtsGHxITf1sJMEF
/cNPWYAH0HzaDEqstVSPTfMZp5woIYsTRVcrnYrSfkupkiY3wq/nrHZboViSkF2l
xtxpUtRVteHu3rZaeV8Vc9BwVkX5+JU53erKL9JFRBioqUJPk6MI8JMMXljv0bm5
10h+/3vf7nZH87Pp5Z60CarDKTcLD51ipIH5TXHDUAOZ10gdE7RSu0IeCJojjrAl
0v6RaspUe+Gbpk3L8JmNjdXZnusApB8odBc9Q1Yv3FgWKX4FVX+r9W9J3VEFDJnk
iUwKGZHm1y8tdxMK9G13JSULYUb83kO5ZnV2c2JY1iyNuEmPre05J9d0BdptW/Y4
vJZS6r7aJr/QbxWON9xiKrgGpQZCATbr0SfOt+H9kdtc7u1s2FKLRUIxPxANFqGT
FPoGWT+tdr1iehnF38jajZpZolsqDwXtFdZjyjL6nWxPCMrs8B63rceNwrsEQ3Gg
Vfnapq+cfgf5j8VqsLanHIcxSgvJD+4zM5urYnxGAg73zpnCIOdOXUI4Ef5gi961
UWfzstQN69JA7GtmsBYiR6F2tF4zG/kj6nuvQFSJ9lVsrGiuFcL2O70mUAnjw2gv
br1aaXNdNA2umIpv3LThSrDdsHWDVFql2VGKYR7Q7GBDKqL1Nea99Ey+CiSvVoIV
idEhA00ujnXUyRRQfWz4zesZ0PeX2ibq2auMtos20HQL1Af4cLLUIBuVirWAbGw4
nVtqfTn07u3kxsP2RUwIuMcp5dRWP/wuOS+LKh/sPHZEyoCxDOTWZ8IeZYBCR79C
aYZSx5nwMEo9/hKg4qmWUB8HpAMZvbGFIFFyOCnbFV4i14cJzDyjqfugTm4PVVbD
2Ie+XF2qVIAbBfepKb7Ggf/p9nVhAK0rS3NTtfD+UEhmJHUmhFS64cuxRAfaeBNg
fM53ANFuhUwliyK4qMwPopJdCbRf4n7ajxXzCwhmTiPH9k/GMju522kq16MHF8yj
2Ds7nrg+Z0MbS7wele+/kCdvV3gGHhL9F2kNDs09SSqI4IJtY1FSIVGBVn7LQ9WZ
53aYz8jLXSi8IjQc2of4qNDK4XRjNDPUm375Fiy9W0m58WfExThDJGYNdZjM6Vhd
ffFY9vYCLPzZAAJyBecvmQlMMz8ZhLDdIfnk0nThF2Md3cIJWvcRac/75BO5aFhU
8eaytOPleI3AkmWYxySFtIeaN74mUveANxgColj8wSsVkmK1bsg1D5fcDJSwrM8y
XtkyFkZ01NvzT81qDfbdkryp/ndBzmkVl5uqahOmZMXpUf/xvXcS/7EifcPC5Lzn
jdEfw3Nsni/QR+QLz4BNe47wnzCubSV+IeSRPPBcHCWn63sHpR51XvDmw8mVWtVw
3/iQImIjQsRLU3eZRhsCyP7mskL+nfts5BsVAZzejTZ8WnJfq+0J55CmCdSCWQs7
T0LMP8JFx5cWypZDeU4hXu8hCODgunMu5eTNTdR0Ij1tXedfwaGDCxYEqEFEZXl1
OpI2nmTwW0JEAKLPnIAA2R8/aApqHfBGbU65k8a2sYQzJPQoDk3c/09/P4UYoxo5
FCrDCVzjRCWb2aavKTUnpKoBKl+o1uJmlO8w/FlN1PhjjUrKL8621/kIZVXDXu06
UVje8I/c1x2DvKtJkRFBdCKfZ8mShVVXJjKUCyrsVod0sJJAr/S6tnQOdVlN1KIi
wg75/jGGGnWMBGCMRQuAElqmSSfKm8bgvOXoKMyndgMlwS33DtHnnycy7h6bl9hc
yjv1wNVA2UGWmtQvjYrT+vT4TmCxLvvl7tfUGDFbOjLYD3c5KvXJenkcKOwfJFNB
Uahq4bSPYyabtRAaLDFRfMN0dEdNku39noSKqhB0aNQIgLDnNQjA/1Gbryhnmfpt
773fYBzIc8hDylNHsFv6uzGTzt2EyLBvIolBBiyalPa/KGHumgUGj1R7MTz2zYeH
IHs4RjBuWQebJwsXYFpYysePG+JfPRmRiruo1DTP9vXXLwGv2tyIFbEQtXiv6uDf
akYy3gf2xoAQcAqx6sC9dqt6I96bSEJSa2qCR39rA6Kg7SKTom7KVoOHhvTQjDGB
RCn9K0Ari8fRCc0lFKJ5gbMgZsdmR8VxDz49AXkOqWc1W+fSrz08DxsfRCULEUoK
TrwOTLVVtSJAtd1u1/9KksVoiOSwe1VzGprnM35t4Fo4PseQod8dTvDAlwu915Pd
Xt5Yk1CEjHW0jgLktuYxnrOAkdQG8DBQMTV1yKOZlxH1/tkB4RYX/GhGN6A7qjYk
g/4lPiSHT1/VDxPKGyAzSObRGGToGK6zHFJm4TMGCeFy8N5oy5nJ/D0VJPeyGpyS
K93k7rMA9ECRw4ulCPLmFRIoFYpLeJxjGXoe3W+GyE3JGw/1+ygRgmM7YynadR4P
jeUw3FgajbwXt4NLPFU5cmBeW0rUMph+EZKsDAkbYsMh02bEf326yzLderxTOr4h
KDq6F+nM30kU0VrUVPXHJzFzHZtqCXSpPXJmY60OC1E3ZDPNmb92zZpgICMioQAr
3g4MuiKIVODKlzRC7q6VCGhhqffNaZ3YG3HYRlkfmAb0WdX4fyIZdfvJaYLN/MFT
z5XVraPOMBVVHxDgmkKCY39ZGcuSA8ZbADj0q+ItCOSwYQDfXFS3JpWVLzbos5Y9
eaz6aAAP7JbcrLBDPuL0j9v43HdBSo1vIUsc17BGZMzkw1y79g6ZTJUBAlW04WGM
wRFvviMLo2fOsMkvhIMP3kycuT1dmAk77CbZOm2ZyXbudqo+M9GKsIOnt26UQu5h
NdpbToQM72iGSAjHaIL9WHMs7SGcWXIgfAp5hXyMPo8TqTtKFzWbeeAcJdxc0sTA
dFuIs5vWqgkDZMBjx9UUnO+btv7OOpfDnQaR/BGnd7MEbXAHsf5SpjzQen8p59xg
EPRKUhLAGj05QS62BspMfElVBkjY9y/F5uyDJI5syS8ltfJ0hxJC4WM13Vvv6ge1
0LH7hQLH14B8sRnA7rHScnvngK0gar77VsV4yDuC/fUW3dzjkF0fz7DPQ2t5CJWa
QtUhyljYAVqCxAVPnVl5TQxy8La5rpZHnOnEXFghWC2VFtNpQZjYWKJA6E72T6IB
vSZPAMOuTzDUr2yRGO6vd5XfurNxpiOuOVd9rDb/vC6h7/gBdK66HUfg9J6Yvlya
X2j03FpQ266jjHiJ+GytN4lspsbh5GHWGy78it454uvwCieh6MDgh6UaOIjTjnFG
rnet/VLvrr/goQKb2497FNaImmeF6byk0aiXf8FUEOnQjejH/fIHg30lYlex4DgC
F54qiP2h/kDdlQKLTq/+i3cJV3Pwm9yOwhGmcs29+oelrcz2EB0lWDJiyXNflWci
S+y8C5pwHamXiuDMlWVRHl2BAfuICcyyyXS45CXfqVAH5mc7CfblpF+DqPLIT3CM
GxC1PKSJNtnRRIuuRcWoaPtOff3D797ATWIM+rn0cIPw0BB6B0kJmrTn79NVjjX+
Tk3eNPDMmX0uRE1W9wGNbWdrB9csv5PXyxhkbuBhi/liCMaCxfK7WRX93/WGauG3
i17F5YEKGuKoOmJBh1gE3Zntd8IZuyCCjgmh7pEGp0nSVeRrC/ngIRyVheYcmTN3
lo+8bWF6rzIVXkGVB/IhcvxU3q6X2kMAKSGXzaWCuwStjeANoTATKL0qbBBto2qy
xOwfsSutjDmHfZJyOh6uxugt2sq+T7F/MKe6yfbpFC42ZpSK8HfkIsazgaVmShSG
cMZn9OjV8Sz7UOxgMyM5YoX+EW8b7oZcWOwnf0g94x9KxHI+wF7n9gCYTBkniWwk
b+Puj7hR5S4df4EJFu2p5TLnTAgrAnJjE8EfXcrunrxww0COqi0kcFMPY15nsTC1
RDzjJ5tJ96KJ5xybDov8vcDfSMK6dJRAzO5oDVgtMCFW1wjisSQUs20nj6lst+Ye
15X34Aau3qZc6xUZ49dog5SrDA88dYr/gRCJP0RKst7346hmHkSApmc/PyA8Y7bs
1PRY3ZrjM/OpNzR8lbMJrq/IFxQ8NIZk+1sw13tcLC8gDX26gL7xpf9Yj+Fo/30t
Pe4CpawDTG8hMLALH1/xb+05vOhociKYWKZqBfXScoqWhhvKy2gN68srol0ydfag
ScLPvpN1U2iSlDQr1Xx7xSsyFXOrcwHgl3LwTTM7WkCAJbDeCCp0x1BC1WUnxW1u
/eG3koA0HVmucCd6UoW+wiunN2s+xaxZ7DUJJFQ+VWIycNtThiJyGs7/6f7d75jh
jby3gpAKezHRJZ77WSU1Q3X5rMrLS6f2Gf6/XvCrcSmlctdLIdc8U+vPXQkAiLB6
5CXtQPQF21m/iFULAiwa4lCKdyF1OK1PGXm58AmwwA1Gfl1lEbkKgo3kmJA8G9UH
BQ8j0EDh0JgRxDr+OoKg6yIDt7b5/gyufmA5njtn8GjJ8oHZtbm36pqj1/qqlrEt
XY9tWzHzhzcAA8uw2HWI+lEUIYBbyz+G0DqN0hjdkfCUBjL6uO6wq3NVGIiFJCvv
O+7JvypSJNhrKedVW/1rAEtZ/GIh+8OOhQZTbKx3hB7+lOsVUyaTc4YSAwKe593S
AEuNKc5a0UhMPsvi+Swkv6Lckb0oKOCX5oojopXozD4B0EgrbckKuDCMQKVP+fR4
EMxnUZpCbPFCQpfIp94OGhhUq4ysamV6FcvunLJ713qAlEZIGukUhqPNtOILbEeU
O7nwOiyFjepz4iccBh6bUAAO2/dR9Xzu2woNPhgCT1X0CB8gLf31f8GgfOThr8KV
e6Qmivz42h2jLwyeb0lgjSLx7EvHyt0l+nasHPQWTmxdsPt0Agneyhveva/wuYGb
6/BaclreWBgVMMOm5QnGDdw9GiLtjvANy428M8DRnK5LyP6STj/Vn0rh/2oQ4x0Z
dXlPVQAViBraWCrAb6zl3TtPCVWtwSno1gx3JvttN7K5jMan/V7OcqjqUZ/wC9Mb
H48nOL+nkxGIEJigiAejTaDzrJkxuwS8i+25aZHe37zQD66nxkL5j1xqit6HLnB/
ZtiljfLllY3kU48GMzpWtBKmX8vcAGq+lhogpVAjgDam+izCV55AEABj8NpFJLE2
1Pi2Dp9jub+Hm+atJ3R04Upf6c4+/iKkVnt4UcVlujWbxld9sZXiHK/EXhyNMZUY
Vb6BCwJPbYH1KI2DdY1RtfRw+FZf/UIPjiIDqpL9vSveyJfaa0pbKjnpJFuI/Qun
Wlivykc4wUJf/ezYeUwfSHf/I4IzWJ3D3xMW+xoL41BwSrnXNofHjpqDLW9dIjbj
zDz3BSvmfrPRyIN613/L5tGH/Mk0odgsCPJ2RMmdjvn1al06zb6Xz9k3bBfMmTbY
l17X3iSv6/Ely8+TeLLqqRTNNo6/prE+E/xsClnhpiAhAsaqrK7eYyAnNR5WeAO/
ZFvAEu+A7RvHRHnbxQss6vDfFIs/B6RM69iv7z5VfvEvKUuxvFp+W1TdLs2MAoVk
Aqj8UmwIiB3wP0ilXxugvYBcu06aibysGr0reskdCndpdFQTS07ohq5jcE67WdTh
StHP1yb9J2hYzRZ/LHuQJKdDAQkbWfRed+6sGiX5SlIvENmzCz/V8sGpWr1tlfhF
jgrwpy/1rj6i3hILQIIX7ht8/5+kpHRP24hl7sqX0d71EClPejxYf1kS53x1CCyd
nilntjZhrJY7YIgXBXEArNybxbKoWggseZUP71xDjxpg6R0k84+AMPpnh24Bksn+
6SiH96O1LXu12k2sPFqqOOwcpilSoliLd2C2W2YnQmeG6Fqr7O1Y1DWXE+fSG3Vp
gw8Tijokm6wmeYU213GwaLkAsDDu4M85nGZOz1aDLqXpJzVyAlT1oeHTnOtE8Hcs
e/dM5xjdw4Cz7LDsnCWm3DOgc9WU0miolTNKzNNCcxmCgvJxQ1rVzYpheVJOsFkx
tIW8madU4fmCD7gEPzKnDAny8UfIUAxX3+b8LRxGJIYg5aG8rlDOdsdfPxcp97Ib
YHxSZcSfc9InR9p7IYm87/rD5/xRkti5zalqv+ZSgb9J8ct32IzYbqZSxT1VQEZn
S4FUV5zfOF+i7kqaGkA+bKpvujSgQ7tnhLjsPr5xc7TZ5wIZAzmsGS3+K0G4nwzB
7YDULEa1C4V1xMjmTQHS1FfoGDE1PnTQnzm14unu6TCte68k8ZyYP1VQi3NgD6bz
`pragma protect end_protected
