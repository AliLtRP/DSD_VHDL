// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:41 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cYDxfLhXvznWoLBZgzEcnmuUUcp2P4gruD51P8wWUJpwlas20M7gTo2NEHOul776
36YIvgvP4XjOt7mOBgx2u8gHinpZUxAkVdntvbkL1ZqYGFxvWshfrp7/XFw1OVaX
/zzYbSOUgHhyaQmEof+7SYW45XKqNye+wOBjRJUKXHE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18576)
AlwvxuVhSaDs1HChhdxiOnp4yaabjd6TF02Ox/Xu+NnIhdGmE9OL3alHOEEe/x57
vFM7QE0xmsJdoimnS/yQqirUAbt0paTkfFf/pxAs8zW0WgZ/TphFXIZPgF2NLbrl
nDVULnvneUYFPTMe2QLpeZSmw7gs0B9voB3voLNXs0+GTuOc7UEqCqDgy7CocdTU
s/ja4DCZQGUlrvjdoX/VtJxTbK3QfKPz14TsZgQsIzcA1Fz5VZd3Oqjzi1+ER1Q/
li9YcS4ulxStqJm36DrGHGl65e7fQdht912yvIb7Z2Q7Ys4gZf4m8FVrOyHXK71E
nq8nWd5gn+mPXCSj3CWq1KsxglqLqnHrPkINv1lKP9vX+O6ntku/jO/4p/IeQaYJ
twr8IwcKg086EAUJij7/aXySdNlS619FKcW/G9C24ZvZlgXL68Xl5i2Z22Os6/gm
TjphDLEyBfsDrZoe1sC1p1fCC9Xmyz9m38nbaeHe8cYslmE3svFoL8Nu0ywi7yQK
sxnuwAoGb8iUG2WmH+nBeg3vjm6AzeQvJ4PqmjxaB39VYFeh4ixudd9fQ8ZcFrZ+
gcj0VKkg0vGekFK305oIS63iZ9+ygYMD8OpsGk8xAMfKDIYTJpIJ+gUYPYVW0FkL
hftV1DV8QRa9PM6GYXQHmftTj8ceAF2P7CJokY60WOsZL6YXYc5k75T1jsc8iL7d
8G11evBj97gADv1gcCE+IZMOk2JPgVepHZTev7vhwcU/en5t9xsSKMShGm1bHSbj
NUp2vEzmeHN0Ps1Eo495LHZ5RdGvmJ5FcnFtXn1x0iNhrhIDau/EghRbBkb32n5s
xWjvSg8XdWVenBZWZzBdAqFFxW3mNCrST4Cq/eX7bm9P9jIyNb+ylAEjmeueb1Le
+A81KJ/evVvvlI9QpZRvLonoPeQhDe7TymGaNSULwpJfkntDghbh39yoFmHy75YM
zoTJDYKW4jzXRDicUkfc517No9APD4bee3QwItsT+uDWsf88zX3qiBUQO8eYzZcb
cClidEscRDMERRMm8/LuCTrK2+HxyCYT01urlEn3Q9Jigqua0NfaXN2dv5JJYklz
cGAXxI9cOZ7Bq11+IdPofKOKyjGBoric6w+0bvNXAZNWERS5Umqaw3A0MP4WetFB
gF2cn3mv9ytHEeUz+KfTQlxGW/2+6iF+rDMApKAKPuDWryFHaP1eg+9Ds+QMHS8a
Nnvz8gQfAZdeLwMPbDLkJXHZ8VkoOYtWXmLaP1U3Un7uCqlK1be2G0pdotxSHQF1
BlfU/3i/YGkt2vM/8fsWXcmyjpWlscBM25pRFifJeoCQ2E5t65srv1CWiY/eXJxS
/xbOl3R6iyzDvxyl4uEcUaxpFaqlRLIbCXd4xJFOI8c86dawR5CO6r7tFCbE4wLE
tUWp0FCSHX5MjBph5qUfOAgYnQp6F7Ww7hje0OC8LaydRKy36kT3b5H21woHFNr+
Uw7QFbipiQCuYLSTiIoa1Ay3z0eUm5yTDAvagLD+qtqfe9RFZdG2DNyGKWEVwLyJ
ACyqfkFx18hNyzc3r+B2sx1oE0AgkHCDlENollC+2XmajXEeWz/lJ8kNhjsIjKle
10jkP216PMYEKX7lJ9JpP9aEfAy5VSQdgNncXN+m7OSzNOS+5AAZEqhwsEky/mmZ
uxx3q5+cJ06mLkwF9YuTxpWqfYKNRMajXT2l1vNNoRixV93ky+m8ecD4acpHVxa9
PlyIg0k7Hj+49gFXXZsOp2TyJ1ssFqiA1EVYiurjF/Ox8xNmrmG+9w3YkE+lIxrY
a0xe5b6UZXUapF1k+bgPJ08saGPtubuFgAdyDorLIkDQgnAJOCHa6aAbf/NvPLcC
k6rZ5wOPE8OUcdfYPBAOp1usBjoQZ2Gkq4CXvfwWg8yV9Ig+gjjTcCplkCf/8Qlz
OjSeMm1G2fKY/VvtdFFyhh+DE1qYHlCr5iBbyEt/Q7B+PeN+DA/V6W6lLL6NR9vh
7hKGTzNoJYlVkIcwe4Cu1wSKYvBJUDaimBpD9uXJxOU9X8TioRHNYt8zhseQjAJ4
alVEvsRGkHUL0Pd5iJZRAbKRjuArRfiu4In53VrqGOM2Yfcko7NfrILa4QITrQri
nLCnZPb/ECd01PqWvLQ5BkfyWU1cE9n7HmUyCMGLv48+DH4uBwINmi0WMrMnbPCI
8k5tFnwllw5HN9+NSpmJBG4tpulNo4u6ACgSYO5LSFLiOVO8c/DvJk/nIxmX/meP
p6o/qQwpYvqCur5OiRydqBzOV6VIfmIETSBTaK6R9Bj/cwfUUvpARzLCZBdVwh4o
GArrsOXpOn+IeDpydC8gSdc7Kx2EwIeilVAcyKEPUHkP7OKgssaFsWt+FPj/hpMG
0w8KHvY2KhEfq/7tP88tOsOUHHHzLe9qkokiasbhhaBagunr+HXubFQowpxGLv+a
LLLLitUJIVYLi0g2mN2ma65Tzr/Nop14J3/v+xx5jrpOYhBFtsjymMXMuBjxElGI
yP3c5jWm6PamME1EcgyiUmw6RvVMgqEeLAhBmuuMOsFBiPDGk3xN6aVWC42rgdEf
9VbqtEhkE/3zycUAYsZ7eJT2OszDZvkOfuI6Yi8w3rBeh9czj2PRwyqT8iTMJx2+
HIjy7AXWg16peSrN2CqW4fehWKxCXFOITSU0GBfwiBgP472y1WGaPY/j/kcUcVCa
e3CzjpHLoWtEoNFuCkiHYG7RxD+RltcAt6HcC6eY3fdYBvippBZro+JK4RWw4m8w
1tWKw+75+wFQRC0EzEop2+M64fEYMwTBRQ+v+DpA1HEDbCiC6fRJvppOPYP6pPcM
zhcuQPvSWF7Ka6+lT9LwuBK0RkxpZ++D/aXAJxNv6jRakU8DJR8pYkxyqL4MR8Z4
o5e5VqyPAixvvr0Y/YeyA4Br64CM2OWi6fJvp2UiYPyr5E1h8V7XB/6S6bWfcnkf
el5LyVnhgbu7TB6q+rBrVaAfNIC/O/3+LbgS56WROfqZshYj/H6Y0sb7ZUTXoGy3
3rJmK5U+8hZkO7Lmuie642a65eToWn65kGTRT3ljfvJJfaURQAOa0NSBQEcfhEvG
9VqW4jQwfGdhw9ourlszQUCV1SFXNC1TQxIKShe0ayE95LD5EslJa4RRMWrMpwmp
65rdPrXM2ZQUoKZ/fJgq7zLbtnHgq8t2ud6ABfD6iPAVbcSvs/QpG2LNfryOhbUA
SZ2mkUa+MjbKA9G7GDn4k/tWkbe+zTnun5cz4HCs9DmfqObvpJdVBZDCDLgDHOFr
Zat0L2Mmtyf0BEo4e+sfH6c4WPkrDBWEKdqPwmI2HgsXq7m4B+CD22GZZ+Z69BEJ
Ck+N5M6t6T8MEW7C34hgw2QdfRrUfb8AEax6kAohTvGm+lv9UuMAV9AeVwbed5R2
sG8OaIZ3k/0ffGWhgwFt3Nx6qak3dqbbCvTJwe6E+b2xcUWmVtzGLd2NignkwwjX
uBaXUyJqGdrql+20gMkdkUhhfP5/4tWww9o8jGkvOB1dJaa5jOgD/88vwNW3aTeO
jdN/8EzVLLFnYQ/7ayeEkInIthtW//Dx0eL2Ylef47m2SayZcVVvFUBfzOxm0B+i
EfWnpEQOVB036In6H21ng3VWXNvntZWN+YIDDmJ5b2y+TeQ45WWT2jna1xvh9SOi
5sUsTGNkCkFnd5xT9JjU6iDKyHO+2rTvFYb5LM6Acp4v/npBwFe6Gjlr77vaerIR
jCm9Zxlfqdn1c2gzxm4G8zyzKPAYWBHoYmRi061IRYpDXjfTjwnTfAjtc9ozSyiH
Lotyoutjlg4odu2pTEGPgFT4+8zLY3geW57VrdwmMkwEpwe9Q88f8jJppFqUlxP0
KKtdetEUpZxz/4PMzf2YKIqw+Ox5G8Hjl+DFjhD0G8JEdr4jUD0TmGNHmUye8OXR
ZQyl8c29D/PWPijn7WrDFT1ALvZRGlUIA/SjiI4GnIBwqW2FMPe5A8Zx5J93j2BI
FnajnG6TBiFcCs2YX4KBWCpd3z+fCweeALxy3G4pvbqU3nGi5BVyc4Z2p+648fLL
T89+uHuouP5uPTaUQidtXWm6ppZguvoFJLSLKSWk54T38DCebSfZMKCDreFEwEwf
fzSXyN+4N5o1JtAVp2H8FgL9dEn825JbYuix2vEdYDJDZn3+8OUvymNlGo8rXFzv
J5hWq5lIIbspglNcegzKDN7fbb4eMwACgaZ8kipW99viL+B07I2ltPOEetR79bzu
xKlcfTZrOGF3gE0AFrlqXnn868k08A0jTn0lBJxQLv4L+6X6/MD1pDsCRlXLRb72
uXa1BNHcCyoLIfN73hDJo7GtzBWU1I8lHRJiVOYMA/kWL/GCTVwrqSmJhGdNugJO
CUhK0BQh4klBBEnEWrHsttNvzyEHdBVPzAxmrNlte1O5V4HQcMgayAOGmUy4ZNRh
NJZEkDmgcldTbJzTwYo8SnCKZX3hUboeUWTi+OncE47zbG6oEYhz4HfiP2ojjhnL
y/anScFj9DcFjeX69aq6+WLj4/DVYH8tA35IyKEbb0DkBTv/gJ/ZE5erXpGpHlQR
vlTHhB1TpgJ0dvczDON9bL1SOgIZYxGXl7UERHwnS4R6kNcVbjg9xnKsdsA2NSVZ
4VlrNqHrWD4RnqdQ3wVJyusVfkWjWBD/mAnweK0mjehso1R0fKrauTMXqdCq8SqH
qDRKOcf5NE80VrPXCnCIA2RaxTNZ7yyi4x7jhekB8AdhbFcyAMYlxA0TKU3jEyfL
DjpMIN+hAVDViMTt9RoNA3ImSq5JCVa+bmfoohrqFlFS4Aoq2BjmFncKYOnVUeiG
xA2hIQkmzWybunYv5MvqzUssB/momkyHtAUMWrg9K0jRENAqJU3ipUehiAGHLd4k
v3S7yaWXyKYFW17NpIjLc9aJanQkX8fOHemKK17BBWRHSZEGy/uBPJX2wx6Yhrn7
WQ5ZXxSPCIGGWmZCKTMkc+YAcpCSItQODQ+tlMzaQTEYLmWMO6mnCOurdkkTkWAX
Co5wxcupzFZtgzrXtlRJ4lDKaCgQxBwYflrCRMvYYghiu9TGmBfgTUfDosrYit+E
0uBFA+amewNNlpeQ5nrnprqVmNP96JShNup8GWc7PjJQqL4gwr8UVhlSt/dkSenH
y8ZnzPmWd/xdT6wpoX+iiYrK6NHdudLc++PuuvnRxpnpRkUE/OMBVqaVM3cYcbv7
W8VvAaCdXqmCZgQfnnGaQJ1zhV3jxdH9k36OryWSrPFsK0a3g8ou2IxOwgzr/yFW
Kft4dcEC87fzimG31eMy2vOR5/H4CKY8fMWjfjsTsOa1uSfFngf2M7eVhmPRL1h6
Wc/fNldNIAKy2QF2KSU7ohvmc0BlSMPtRI2jGrBC2TNYWrYPx4l8uSvyHwD5MVJd
q5S1BQ5IHfR5V+qE5qHLSbHEHA1nnxH7dXAq31uZ7jsij6R/bUcjYywvZXoyRNR8
TbEXovwScNAdaor2Kj4DOzVQ8w09XTJUHfy2xNPWTWhFslkNmOUQZQ8QaF917HG7
1IczJYdLLQUnLCq/s+2YksE+/wTxzm5O+sJKYskbj6MhPH3xMxrYxWXFgNzB9Gs3
JVIB1qAPzDMFcnsuJEHr087G3CLCP5J9T0Xc9qu6GG6aoORN/sK3E88AT0ps8N+w
REPYXjDju1sFIPzjC6/U87VIOPGAb6VBvZH8+1kK9Df3fvgRWlEVogrLH/kDflJK
ru0KbJhceIdKO9xy29KNGmTQH+rSwvFZT53jLCcZGu+lX2jY+b5iomPy05UQNDim
/glZEVzZDUPHPJz4l4jxDRFQdVbhciUghVEojAJLTVI0gBGUxL/7CX1LIDiuNDbr
0SDMtdWRb7PyM5nahoKusAwIt+P7fp6jHXS7pxVxyI8tRVgIFxps/NrQ9Rkwgfst
O/n6vrhLO7yuVBx1weZqYRAkavnmRajObnoNBNon8MecV9E6TbHEewXGQzhOOIbH
3JcUMKND1uZjFjokv9xfNpvmo+0bNznnnBbOGgzbGSSrPNqUhjMWAJFdO9tGf6re
At2Sa1eP0P0VNHkTHy+tc/sMbPhCYiVPxEI38F27bDEjEBuP+Tuj9sZutQJ7a8MM
49YgC44mKScx40RyKgJ+/PoM/1svvb+VxNI3XhOiRJf77wAYWmppQg/qvKuQThip
Aih2Be+L9A8u09JCbNNPP7soqKsinNLdktuxUn2bkuO0izMW3/HwftrlJZnHI26v
E8HgadnlWEPbDCtIm6oXqmeIDx60NcWoKO1gd8ryQSc25nTSdhKGufm2HAKBemCE
NSZp/KnN9tpqngHoxbFXfekpUXrO3rA3lkoMA485PmUJ9Hc6+XYA72/V7XQfTpDw
GYwbEFzZaZMYN/vZOjkN56YYDA/ibzLnA5Nk9+BmG7cts2dFletqBAEiHEcrepbl
TMKEYmM8VRirmDV7zotH2sdlmNNprPXnPHwEmRZLix0GX6lfgT1HuuCa8lbAExdK
3EVaSMuizw8YjMkWeeOi1kolXkoo5Q84Gl9JEQ+MImm1mMu2PTWb68boh5KI9Hpp
PHio/mjwHUvAf+ydxkSL8vLH3Euo46np8AFu8z8O+JRxnWP2wUGK9hsqX6G5zrCU
tVf7VZ3Eabv8z1GLw69U/SaCEwULmBNnRjMX80yS4VwWNDHQGXCUumPxEKffpYfG
quf2v7GGX6A1AaKnVvc8SyJdX4qnqKD7FpxJYSyitXwuGaNeYPd61DAtb4ae9FTX
fcX4+P09SCgkPFwUriQZ/X2fgNosJhm+S1+Z5rnN38RM2N8H+ieeLR94buCH0Xpb
AW78cJZsWXm7Mq9JBQvPjKm588NeFdVoQxKVmGsgbVRbpsbqowWFatdkg+DhDhdH
tJZ5kmzPzZ1vbxGL2vkGFOZYQY0wVJ9nd9GJRg6RdxQe68BA8yI6WkKDa8NowbdB
CbS3m36kutKQfgtZUaUCD9FTQP3grgZ0Rz78zU3IIYKt1UrPE+0M0bnsVIikqHga
6CJU5/U2aJKQO3Bm7lQsuiI7gUOF1t+Q5mk1d0tTKKmNEtyRkiFFqpVRfwYZEvtN
uetkOvXraFJ4JDVkEKMJag9Sm5w04DyFK0nXvPuCOV5AL2AMNDvXVAYb3Pg1f7j/
mgBt9FtHMCkySa10JDwvE6MfO4V5Z9QxVlaUpOvLwjjJOK4NAx3h73MfmMmdu2bq
M6IhTgVKd33GHzILsHPnToDHs4yYin0CvT4fnTjhNnTIU6zjFiBJB293pkhGLZtC
dMycQI5xZoTMleTVSonSbz8oQJ7US/zSx6QjeT4dee95nswCR6dpGEeOEE1+BBmJ
EtYeru+Us2OlqSyg6p3zNrC/W9py11t7e70q9XSYVPYnW8Xyy31Vgf1XeDj1S3eC
Nte93QUis/u5BPx1b6P7J0NgOmNqcGH76kWOFJxdjd9lIEkFyFUi5bzYXpZrXoDH
10pypXlg9rHZC6uaPtK65rn1fZE5vbNpYG3b6yKgBMQRq9VjNPkqRjObEuJZlVX2
r34wvUv59ireX1NrOEcajM2SLvE2hnFXAioHY8/BIzdIUNLFMnQwQDBtoVjjOTQT
Yo3eqBX0S11Rp5TRSxPbn16AsIiI0WCdprKDU4HK58gM3hbD79BZmUKhegUVbBxv
GCBFNb/9f/Aut6G3683CdzgqHEPGR5YR8BQ9SCyoroimlabFj6UGMEOdBv16WOXk
cmu8C8rzNaoa3FOBMotmYz9UKez8+7N7pevu3EXE5uZqWP5X9T32dPOv+3EMIyr0
Gm5JBLN6oCcmpgp3FEe05uAITTPsdUboeR72sa64cqYRb0oNWcWT0iwwtIqcnRPy
jMWLV424en3lebMDf0L5FREyxEIG2WwjZBakY2fe3rPzRyjrop5K2vUpNz7pf4W2
H80cOPxyuj85KbaUIf5o7YOnbzCjyY7HctyLani3y5Mtkbr2jwbkHlt7ijY7WcV9
4kWSyDGpzixX//Fe8Ud5O2VdTtAIIIYLkUoKmPZOybVADQn+N8g4W0vh2ax3mxwC
MR08i/UKiROAbJVnyAVrmD+PAFT2I6Mz6/lQto0XqSQxMJE43bNM9vdkX9Qv50Qi
QWQdG/V8fydmB0qbLWkFmvkQj2x7zrGmQ3WCNOryRQGYtAb3L+4GCwZhpf0Fa2sg
/3Fv0dZJV/N2/xEwtxuDw02m7RgUxNYHzT5sMysPOlXcQpQ9Ow2GGMyRkPN9GKDO
XIOjsVk9Cz3hu6/nMPzItd7IWi3S3nRpxk/aFfcXKtraLiEbcJi471LD1tSuXAwn
RzgRaRbshzK6atNStPkJo3/wDsfAO9n+Q++eH24O99qYna3YCuNhWD8TJode61PQ
ZhIq/uM3QzcoJLhQWsZtk7c+VP9TENP1whnnVCu8x0STa3dECM1H7GyvjxbBckdt
A0P8ovx1HWOo3xp/S2oT9uk+juXuo6laMXXhRbSy41Z8Js/dprjlA/1PKf1M4a5+
rFlL6IPXLP/hBD5gEuFivI0pJWL1npRxm4z+CVMtADKtxWdjKkYmo0LZSKsUkWd4
zFjioJ/nW7F+dhzOXGAFWpXvFZ5ji/R6lo1MxMuj13Pl1ql/7x/QuHeTIIcKAoK8
fUv62r/NQFmxipKyLN8GmM0VncN48le5aiNQ+4TIclN/uJ54BfGQuGOCN0GMu9op
OXpYEYE5T3EZI3bgu5YHljhe4KqmyV4uSmtFYwqgANMVxiIoFlE77nIJFrPPM1iY
ncLBvX9nlRjhRjwSDI0XoIovFvdYoJJ7DjZuoEcZ81DbLGyQ1hJwmByLPP1I3863
XDjkeMa16h3zjWoACWwM1J1Ki5x1MWfa0uCQOnimpAM6mE1yKg3TAS8dmEE7dmVm
3MXht/FhOkfkXqrqo8ggWd8+MzM7dVpiL3GpnroobeV0cKji5X+Qdw6xtUnhNPFG
DeCl/TZ3vCs7QfHaPryo8Kwi8Wb/fdQGbxaYI5I8iYMipSqCtTHqklFujP0xQ3jp
Xm5hY4DWwgvKzer5KqRnCaSpITHZ7T6JcSKcRiu1N+/dMeeyxKEGDOvg8Vn5CS2d
pqocMGtg1w+JuZuH89AY2wtmX44qmQP/zkyOrKjl+afBvi6b8p6fDWAf8WZzKjps
8i0cO9Zonw0oVzV9ntSZF7VraJGvoWMEGh21HQz+yNNyFc7yKbl8+wOvIsSUnFcD
iqiQF6qSgjRptrJHwGbeWw4XudQTb6JLuCSreYsLGahXbn6gMQJvFhIvrHP1FYrE
UcOcFZWiAlx1TtbhSKqkvtvosVN1I94qb28pLF602ExKQuHOBDkATy3IQfz2piy2
p6M1kOm7n2dZdKknZrPMAW3QOOodRpSU9SXTYaFUZ6t0OCZeEOX7fNJ7txegsFTN
QO3z2WVF8sVWIlMNepP87H0hI6zhFS5CRyP5J09r9NkXt22E/hmBCZtaZTjbD+MX
MOKtvckshqtiylKyuO9UZkkQRKiHluCIIWhOWh4NV+Vr31iotouVyGLQPTMQrLnK
N8S6RPHwUQW1vI5KTSxQKFNgYd5ZR9Uw7LXyXcsSIoO73HcKztZfqCgWz7cW/a5f
7FllZ8oHB0oSxHlLjv7P999kSvy/khefFtSzAjdQn5i9bXrWKlSTAtfz8Y18SH5Z
TV3y0Fsg7huV/fgX/Jf5wb5swOpht+5k6MSmTkFJbRs94T9d3dSHuBdl1kXiZanw
Lr55uOniMzdiz+D2lElAd88xGntcAI2kDRR0c91yUzua7CozTf8EFyzH6LhvPZuz
gjQA6rWNu3D3NWmGsYae6dlbbqpwIJk/JhIGxuiLEtsEpJ7pZ5ly134kmvDYhgGg
hm90jfFN/ky4rqyt79ddKsk/QWq9cJMB5cXOyuKU4+0+GLVVEzzTfkvpvULSZ4GA
9hCH+IXFQ56mWdhs55HyWmXpnSQ9sOoVB20UXTgjTrEZZyDaVnTsA9wyKy/b/pK+
iPFWWArP2HekhkJAr3YPtO5fRmsFD9TmACJxJoj2m5Lu5CAn1GRssNhVvlABmm2y
GZDqUcqp2YfBSg5QU63CCQzcNLEiGmnNItzwWeI+Ef2w5qJO4wd8Qdj0+r5p3alu
IcYPeFROCNkIqMMvHOPVczYXxVlbszJc+gI+pJ7Q/ITb8Ctmv0GlN64sgl5Gv2Th
lpFmPl9/YxF/IuZEOqdg/QyreTxT64LjpPbapy3brFaVqk93PsAL3M8HNRNG+1k1
Rr73sDziNGlqCL8WGFrhmBFiU+ZFm/AnhRyGAG/DiWtu1AsB5FxyAmLYBkfSLnch
gYWJHcprvGz6UUHlWTJ1P7p5ZYZ+vTLzToFgyAgJgibUBuOLd4Dm/e/C6xoNMHQb
RDtcVx1JXX/HLV1jUVazy1E0XSNWTL1L3q2x/X3qW5VxMDAILTPrezOi1L4LVybk
AqbL+HCgbCkFtK6BSaNSV8u9mx0iPBLEjg+Wn6yGMqFJyhN0zojGPtzKFYrcvsXO
VTbHhaby3Byfo1xu0rcxxTwUwO+Z+8tLDuXhjUV0UaRPHDXnpb7RvpAH+Y/iwzji
FppTycNhjmYLRaVYODP2ZnSBpTir40LidZY/PYoX8G4oqWSJ1nNDd5ixrVeW+ut5
JFCOydAi9/oY0S+JoeusDI2vmEtZ3Im6LOEPGDzZQHJW6RhtOKolBbnnFkpUsG9F
Yg7diiuf7/qdPhTfSwoWaEBqJUkUy2wejepzK9LEbenhBWXPUjYfCZJKyWQ/uMh9
xIy0PX6aawEY6om0BGTICS+uOVvX2ttDpQppl16ofKmkDMYxRwsXDfPkTALXBzZl
mJWrCIeYpqbwvkyWkn2S7APqIgk4DISwkuELO7YS4q1e0dGVuRNubsPCGDrRzsG1
gkGGj9EjURwoioyKAEPWMmliTX0Shi3PoxYDQ02/+Uoka+R/BfDhCxVXE1S6kS6q
iIJC9aLGPYj8HtTRLqLndbYmy18mar4+JdOtBLQcbj6P625GQ1TdagBqPCPxL3tY
WupRZJiMMmHjFVcGXy/n9SFlAi2J+ZsiskcrDrIcp6R7jErT7wVFLKeBBu202mGL
b/rGNXK+PM5A1kcqcVmq5BtT4fv+eWB/WpeuxxXC/WkSGNK4wibJBpjuTwJWMdwf
6WKPj2rQah87cwF0oAehF+Oft1fDxeYe0tkJw8MAzJemwRAO4DS/ajaqiw7g+bfJ
RI892DF4VcpBACrd5Saj6PQN7pHJfz36ZViaKaZRpomuhPZhRkiOtzyMsqGnEhio
+dLmEtVA4Htkd99bOWdZWnDoo1ZfZD4YMYQlpwt1Yu/AZdvmW+g1quH/SnxQHbED
rQhUL0WGfgBOWbfmIADeIU4nkvEzR6OM8vptMb30710jwZsEZ46QSCfLAEuMY6RK
b+6lYd+6beBpSr9pamDo0h4YvQ7TJ+V+Rcdh7jeaSsZ4oS5Q6z3tPqEkOWZaxdS/
CUwUIqT7UK8SIEE13ZO55bPshYZFUxD+owbuKv//1Z3p85w+ivMSmsHNagA8ezrf
5kl9jVMCViTq6Vohig9RIvNN/j/NVseNbEhf/YqsEbvR3dFQqkTbbdUQzNIAjzZS
yqJ5okWnec4uyucx/ibMS7pMnh4+L62Yva4NOgq0a114UWjpqTXbwkQdSU+GFQHu
I4lnT8aNHdvGZ4Wz27bangEj2QLX02RZobSMuPjbrp9op5SdLTJVxu/o3TOPBQiy
xvbyREdEsVhD1Ust0aI+XXLkvmEz7lUfDATPrCIltYUYUzgZGvzzYhMELfyE3z3r
YydhnzJ0m/ZJZQ75gy4i8GkVZR86BEDqy4UWnaXOC/RdTIJfR2fT/dRzvCLjyx1c
TQmMT7DJdsK+YTOPnb3vOm23M1MX0Fb/zLnzd1OZOiJZnteCXJMNXVNz7qE5EdIj
uSlSElz+3wkUi7CQ38eVuInGtcoWNIEpfdiD6CAS4i2PE438+7U5/s+cXGeLoX1i
kxDvkpOVYuilS5/WGifJn9R0oliSoH6vYH+hIbf+zvccfMUYs914JOsvQVfQ+yo8
QSuQ+c27T2qzzE2fNZ2Qh8cPrp+0uucUl9NAyzwhGx6nZfYcGvoSLwfPNBXAM99d
ZLwrwM3N0gkZr59kgTu4x+p7zqG35KpWxlCC6PNwVzu9ER3+9cZyzh5CblZ9AY07
aClENe4WfQ3EUxRTYhP06Qow93Pf9zIYo7A6hkUthfrp3cuCwYZ+2j8cI1MKpZ4H
Sgs753TQtbCQO3i1hBzaK4H6K/5/VP3f144z4ro1HTkjZydVmpe9BFx81rql7J1Z
VzkpggEIg9bUJxk8RLEYMt4wtI5KOESowybWR4ox2nOtqPNVuONsnjq6SxbhE+S7
naFBqfnaCTAzc3Ns4fXOZywvkdm9XxUTI2ZcbI1WLrb9g1WRu8ksblKO6ZbOp9/p
Ix1RQIY/zLP2zJ3udVPCJ5jRr63JpaKz4M7Ko1r4hmb9yzlf62V+RmoLr2Zfh0wj
dgy6xxPcv+UffTwtQc5TNo+XutTu2Tl7xH0XeSjVosV9O73jPsCRL3BPDXlDGivA
FGz3wFyUf5uMV9VeAlBQH+/NHfHO07KxCGojgKsO3JebSezwxRc0BFTeFXU4yy/s
5EOn1HldwMNL5Ujvu5onEno1lecz985NKjD9xu069FJOm/xo4CTN+c9qHeYaeIIQ
TjCiHoQLGeIA2o4zyQaiNEzljdEyWyumpbFK3a45xF9IzD7bcUPOsXLY9XyLdsnw
OfuZzTAXniTmBRaopPVUKb/rRSseLB17ZnqsrvJ4L+HPojebT4fB23Dul1L3vWDG
SfI+hjKExT+MKzWPkxHONOm5a6JJQGgjL9+xeGfaDgeiTOu4c1xFGUMk9ZURZsK2
ZJrL6dnxqopKOns8jsCjzLHn2fQcQbJ+NhUeIEfOY0sMLwVWqpiJEEqzXkh3gqxc
hZXZry9G9ywyt8TJ58wpXT6KTYzsQ3WEY491y5aCwDbEs//ZyPwokfqdVwvxBYRs
vnMPzwToWnVf3IV23+UYLGQjNQGgwvlCWI/a31ZD+gLB6/IEUSuRzGI6ZkYdcTuz
AHFnjRVFm2GkuvqjtozxF8Eoh0kUPbcESHg5pH/WDv03epx13AmyfKM/VfRo4Ed9
AeigAEw0/rLSSKCsONgmgzr+fYSNJOp4ufr9XvA2v2Dgcjldr0v2Uwo6WaUaVJqb
qXip1pzD0NO70ybUcoEDyzGTsc1zAudS7rj+J6er4ajRvsAXZfIoXGyDQOPrCHAs
qUzAiKKhclhgzi5MEdrIipvcqxYep0fcuJXXpB9DVWSbqm3U2OQOHAH0xqGBnwEq
2XCac7xNLlq61DxCJtwxQUbnAqn2KwoNjsHvWmH3mEwXhLwIY/A1QqqQhspVHfan
160QFBJcVpslc7ThJQf9Ut5IOVpQXr4IS0yToyrNZHQ329O2QM+CN0vlhHQkO5ye
+lXLVr8zDzcK21lIFGMqwBFG+ASwvz6BhUxMcN2Ki2scgIZ1UH0Wg8CP7T7r8j+G
fLvhYgcbhR3giMU7Mt6I0kH8ppylVIzpFOASB8wtEACa1p3sS9iS01dCKf94NPIq
AFhWJsScQq6eJq2rg6uDvuluHqIFFj51oHsRqA5juhG+6lz9BjrDWzjStyrczFUk
NEg0kCv3QFE2uZVjBE3JPc+NRPIza8oTc/fVOAPG7Pgo31iGv7yAgCmxIOFMRCF5
d5WkvDNAzXij25XuZGCv0rTepcJ+CugYv282XKbvKVQP+t7YwCalyeu7uvEiEUJJ
V/usLdUHzroD4KLvd9zZUAk56M57zy51KkGGtuQyWeqy3kVMFclx0deOX1DJf1yn
amrVnXJr3rjiZEjl4N8WUbveCg8zdXFTC9iI9r+bVGPoCuENIctIJM5zticz+JCD
MdRPj2KLW2ScndasB4AcHjod0uhfUB5o1AvKoxssx0+aiSH7WwdyolwazB+NDoBt
GQHxJK5URROuz9MWwYCsfetaFYCFUzxvG+6ndvqLZdqSzdVSXjexclYQ0ELyl+Fh
zkT81tvB4uLrUdkRqK+JizA3S1xwlExoxVjj0JBiuWWLlV26lD219keDtqe5WkAk
3JWOdKsL2gFag6pbNR3IFmYNl6qioVvk8Ts6jVJMvInwu/nrJwUzNhncripeDAeX
DTqnrkTxBsAEYv/lAUW/bd6q3LyR1nRqmAAs1gZfVdx/NAXOXFIbrck52hmTYs0r
yaqWhHleS9GlGGb9nSa6E5bod7fpY8LMTJWajnclDpfjRGn/vIfgXlqMhxUKnyO1
2GbdlM0hkusfzSrzI8ayak1Niv9TgHaVzEsmpYegJ+SvPuJscESSzPwzuwWmcaQz
1e2l3+EPLhQZlRxwTWYDX6ICQRoDX/k6xGSmGx5Jhk3NPbCWkI7mXljkJ69+2h9A
jCVGknkn99ZJ5fkMtv4aFthR2jMTG6oulM2DRir+sN3v/lKnuax3U+ztZ+N3l5EZ
ClSPbDe5k3b8JAaWdgdRGkE5ybU45A9rv9bbgsZh3fjnD91KmatknA1hIX4x5U7C
18CKjPyMxWlOCabyWv5mIINWnKcZ9ktFw11YVRSe+2snbl1vpqWgn0sHLq33xgjQ
TnGvdB5GmdMty+u/Q/DNxWrh9yQrv2ivXXotYY00XdTa63pCg1u5xmWHGCkUOks8
to/hYdH1LTSaOJ9eL4rBYYgDr2YsZBTyqTbKYDv4M874XGRVaw1RpwXAtCBBWBYv
eA8JHX8FEwtoY/RkQNATQPn1aoGRjLwWXJd3/DniBN7oa8r2rRNM4a2TPj/734tF
INZLvME93iIlpyI8Ucc1ORYhBWRnQCCoQ/9VC7fGXJ7hScKy9shWDBsWxYydzSOv
nfOJwUQDDaiS4R5/5KMTaGTR130ctfRa23GqO4JfhTF0M+ogZ8qnGBj+CELma2xB
Lwtk29F0ImuL+XaNp3ZCZuKCyMrVcyI/i7dQo9+/g371iY76X3pt/bktkVreoCEp
DH+Rq+g7INleo8ZpT5L5hifkpw7h0H3WhXmQ4/xxao4QV9dnwcfV5fy33JfHusne
O0Tv8Z+36eelAq4qEHj7s2WVm9ME2k1109Oow54lt/+QTC/U3FNxOfTx5d0hL7vw
J4cauBpIZeoHdkdrip/bhqlCj/gSrhi6/b/wbLaAP4lfWX+3wZCKIw+UZg4Sf6UM
ZkJ2hwE33JDPP5tMekA2jUXIZ6pjDKlpyb7XbaO+HzvjgBsyX/dpHBr9ONCwcEYo
TjBeFdDI9dBgnM2CFMHafNy2cZvNGtG4rFOdd1C0JbNd2aj1+iwtEa3vH3ewAniq
7ah1ZPI9qLgC9RJxsWAnHgzJlLBKotqMhyazzULLdEgzv/zHkw/xHf3+qsjauOxw
zEyFg2+aixyZOdXlrcVOMlusLyrqS7i3+FmwrEm2sCNC69M4xg7oc9obWEcYUxje
wMkyKH7J8FxhuQ8YmPGHkzKzNAvNy1r3e2N9pC3ESGG7xt4eyFRFRy/KuVkEZb4L
VRwMtBzzWD04ttkdgJfzb9lALHx64guINn0YxJUDGxGb3AExI4tvkcL//skPscG4
ZuAvZCoXb+zMAHT5z4+tmQ67w26FbqSfc8tkjm6rXE0YRFfTAlyvLWq5gvzU966L
lSWdsnNPwMTQvnBNyJyUGv2OZCyrnYT7S/0/lHJ8flTDoK70u3Iy6qpzT08e9hkn
p8DSdkEeVgBAQzkHhUpB1HVnZDIrsTY9zN2UKpmIfu9rhHjNfh7xi3YRfAiUixws
3Qw02D4mmHpWIohZLztUtZT7tQqH46x+E+XCvS9n+bDU8K9KljIqKC+agng0Nrq3
2xQgddEqJi4GRQLqDABqTGF1QIesKBrI17UCsqhHuwL4FciGE0F92jcHHISc9WdY
2CPgH48UMWhrVtjPv279g1K1T8o+fRvVSh6BcgatsgkU4CE57IvYvW1FmykN33XE
fKntFRag+o9oFo4p7Ur9Z2NrY5J9my8tv1PbjR6GVmrD6baIdG++NcEYM6yMzrqf
XHfUzxC+DXBb1H5ZcZ0JyV5N1PGuFBR8nRNe4/ryMkDdRMrjNzZteOTLA8XOfwjI
xeDkSdOVtikl4RoNcTKx3UxrbzxBJsJdT8YY+xMBXNQvUmY235Xx0F6esw0KF/oX
jKJaoLav0Y/qy1ILduD0+63cW6ie/5opEhP7mUjrilYSzIFdpVdKZeISaFUxoldh
1mASzcYWcbOCHOiV7VmuUUsmyzpCjFGfopgaLNBNGPcmAdsb7xgW1sooTvaEmWHc
VvDAAGnDtX3DAN5WdvhgQwWrmPioHhN6+oL1LFOKgqAbcXjb4NZLQM+s07wddSeP
OXihg0CB543MkbfIM0CQ3IeVp90T1tnZJ4kURbLl1ZXcPdSIZqvwAG51v0l6dq9l
o3JpBWWlZneIJ6Rxeh2G4KpDR+y8NYH7W7CMwmQaNnDk6ArQGAfAGsfjPL9PJky+
vSBT8cgeK+iPU52R18mI8Mr+lKS73T4fUXzy9vNHRsA4+thM13CP4WbUWo+74lLe
lXMZDinD391oFcdZ8mW9stDB/E7Mb2ru+Y/YxTJxolSBUmJZDk1HdtWhG3c7F51r
L/5bHWSj/nzOQAahF51bU6QQhH+6iUOHHV47eK7M5w/P8lgzoBP64flEqvoyNm1h
bE7zQ/TyKfQ68iBvusu0HG++5USA7e9803ywC99EjRzX4hxrC4BOPvV1w8c2ViOh
oYQCxhdewG0i8Ro10aO2ZBQiCv/w7ldaoH4IGGcCWOYoXrJqn79B7BB6WBjsD3Bj
Lc9f6VJ38hmTph8IKJKE+d1si1E/KdJCKU6776Su1Bz0AA5uLsf/5agcAxoMkytb
/Z4U7e2v2OD+fO+cxh7wzZJ4cn4e7pdQCZXjG9P5BzJg99ZUJGg7Mdh3ABLSHnK0
Xc8+iGqVFZzh3Dqco8a9Yaura6ZXSJ4/u+BB6FA3WfoqvWUeyp3qkZYJAKO6kvyd
r8G85UzxZ+ziIPAaQf8MOo9evhq69WyClszU8ykhr9xj7cU4kPKa+VmPnYt7PkQf
3t89d6eounVoPc1ZADxUm/mYOSHn7tv7gnsd30SSWCmTw98EGTnk3TdXcEqmkf7D
uEqW1zvxvgBcBlCsjwIg5GJadBh3lgqXTHno+YdqJ5+CP01f/KPRwhnI+A3cB+EW
aad2YJDjsha6J0mSwg9kpoB0BkyCAPHWRu0v20+IwO0tu+z9a/MK1WQnx3iB1iJH
CzxrGSR+R+FhTy84JSZ8lzIF45E6AQF62NyTvfAsEMsoEIYCyfmZz7ptv5wszDmz
0e0Yi7x9Gf7nBYPxUbPs/XSRx4cJkc0tRi0Mr02iiaG04d9W+nLaGrT6rGuLy6YS
tBump4xxcPeXkBSHkoDSVas1eEpEqGPdzL9qo/BC75BZ2AxFw/QhGkn4gAMuU7cf
MI/aR6kNRZDQYYZiDnen44dvyQ4iHiN6jChf7MXUmyzTvA3dCl3YZVXq/a6RsvM2
3QdUPYDwW0rBzgU3FfSYNzM7pRWwG9KxHc3lLiUy/ObKMkArWiHvkv8ujKO8Zs0+
TWRB4s3fkyYXU/Cb23L6hk5p1U3tvt5XfHLNQMhcCBnn6vxEuXEe8ybTr/io3t21
mV8M7Iaw+PXgY8ZPLh7Cb4p/K+T95brMyOnxfGJXPzugyVr1TdnWr8M49jtb9wbR
UBNe4gVtDHr7aiUe8VspxibOWG8bZ5NKekcowsjBTJnAwPOzDsbpfEceLI3nliV4
OlQ53u63fb5c9aOzXkoTkw5Jjzbv1gBtoiFDSXCKxYrwjEewO9fZndXa5ZKQ8JSg
prnh6Rqmq7rQEKKWDl/1ZGMg0wJQMoutKxh9ESZy5HN6Lnm8cMaK6CJi2aQg9VgK
FIYqN4aDhNmsEguO+Kh45kjrizX1hHVzQ1NsLuVRqM3yBziCOy84F6Mulg0tEJYC
rJaZBehAEZxy5qGVfaONUEN8LxI3l6RLVmwUIYaOolNN4GW6d3o73I5ez9iYwOq/
QZgxVoaFLLYlpP75+vKdXhNfu1XCgaO7Cz6ny+Dt57UD7DkQjv/BBn3p6/uD3Yok
Y2BSdE9fDVhxphiw1/TvuVsUNYpqGPhpUoOhcu+HOHQ0jST1lISp9lirLrRFN3KF
y8T6GtgKMu4suMGnT+L736g/7bVR0fFRuNQxStUR1d7u6cL+rhk8Fk82VwqVJ4A+
5Iw2+O+/KfOPzMWr83p+1yKV/cMO1Nxa/ntUsS35Mv8GKnvauuGA3/ugsiiddhG3
+o96uYpqacdkBIaRvl0EBCZ+MfY83Fd6pBswi90ntH5iKkWog7zrh3AAhmO2IAho
MV+tcuIW10Y71WtHTUNuSVGcbWzsbXVwiwGIlBycPpcHK0/FalJ5vicC+J27EO+6
QaUOJ/MDmAJTDo+mJwj54wlHRMHJOUmOfkhOEwz3TNBlP8/5qpliTmk91+yHjfic
TpNGlQbM151LIT0doiICnOwaePc/SMkvXXrshk1phRRuMetEoLzIY7AIf12gSrTS
8EW3IKM7AQDab8va68YNL377iLUmpMuN5OISo48Hedjdv5HVzs+4Vs7LpvEKVlTv
LArdOSgwXmkWWvI5cTYWYw6AwLCwhmbRCz80SnGchDfVqH7cFuDucTJmuM4iowwy
mqgRMKiSIRNJiwapeU8gV3nB3WsLdDTTWUJsxFo9YcVD4m/hUP+0ojOOW2jYO/Ug
MQTsWxesxz4O8PP3NBEGAEN5IGti1nE7TUHMF2wNB6aI5Tct3nMMnMKQaxyUb+b9
De0Rihcgj3wNBY6ipOSVkhCwQqtadP7tr9ze+UbcW3bcVhynJBMa3YlYLrnXEjXM
/9ojrZXkR3mVRJpasdovzzCOXo/7P9gK40ZAHF5ECwdZP2+P9eWRoM4xt0Rx6+HA
4VUc7jVfzLJeB/8TromANMw8VfCyWNsIJ/ysKkOrpouO50DcZi2wx17GEfBlnmWB
AMLshqZgC4yXSF0K3KQpL+f7Q1CAeUqxqT0qKI8NhpHyEbKr/fd58QFqme8aG3sr
TZ0h7y0s7Kb61ykiHxTxTZD1uaHSK4KvZ00UbAEJB9x+MHSCbtSil0M8+B0dMgos
16plP8hU0Occ+cVMdUR70+qMXFzPjcQGqulVJXr4JIsJyEONAGSxeYxwLyu37U3I
WQ2v2t7M9fiXTnRwdvSFZz/duj/JKIErQlym3Jj6Pd227Acjpc2rfIrYUL5kZaNd
GdRWONa43UdSXiu2ky6vc6zdXgrAtxSFCl7jb3Jz2QBEAEh5YROAS89NgBucVnM/
c4q986m35OTe1q2J+AQp96BOeDStmpmojx6huRjxxcvIZKvmeSk3jaDwIn73i5gL
mbkOqjGxG/49JiPge090QPXjqPCgrOapdBgalOUJhDOy80+yLN+u4OqboRoK41ax
yLEBZxhJAPLKRb8ZDFpk5yrvvAIh7fFp5YNc0hBXMpWEb5ddNoSBwYq0stE0fneJ
NnwGX9EsNsGWBo6Je2UWZ4d4LRgkcnxdu7srCyhjd7lJflXSuVWW1CevAplTlQ/y
smkVg1bGWXXYmni3Xbh3V24IBFHjcWwFGr7bOIQ5cF7HDhlxzWtzQ6TkvfUDqVMb
4SWAtXr7mip8Z+N1gg9tikc9MxWX8xC8SBNoRyvs1QPFfrBs9JLP/N9LmkM1NsY4
yhA8saicwwBl83tl/yInFUaUTB++NCvxIgxV/ZP8w8iZV8gm2FX8k5IgsCLzWJwg
cbukUXr1eJB1+3gW4NifO4P93xiGtJrBX/qkJEsh2EUBFpUYl/icsUZ4uwQ8LR3C
SnJODShExYfvj2P7+2EtHAMst9XHLqwn7iikKE1UsqOr9VGGTKp6/EQToMuln9xM
Ze9GeLCvrc9EvwZQBq7TxgopTlatrikLMcByXiVw3OCrUk/mi4tO9qzrK/H9YzW4
l3nFqL/I6FrzOhJHkdRazbDPWE2Z9sD2u3bWPAYRj0kMJ6u1eqC8iMUzDUm0OU2E
nOXqhPbMhtXkIqjh6IS1UeJ95dli2jBjgPyfmS73B5VBKXwkDFZgaRuV625R3asQ
xTPchjDspwbreV17CvdMfRDtnCJn83CpfMndrusMYb3n3v4369yoYttyO9PuDazf
5MPCH/vT75CI4LPGX9cKKjxur4sesJoTxdj6mUxuNrcvn6+KVdV7v9mU0wl4TCx3
0pPBDSiMjezBAFMw4vsSd7AqHONmUApngDggXkqGoC2+oYbUOUpqOznxE7tWTZ//
LNOen6zaXqGVBdBRhCE0IaHkzruLHhRuD5mDZbKVAHCCCJyBTXJNPRI/uB5dyNu7
3u5S/yHasxuIxUQXs1clJ2gAlJ4v77WOsrfKL+AsWlKXT/1lmhPAWXRDW/yt7Lnl
jXbtNBTfWRnQT0AFtNBs0q4cPKe3JLRrcdXkvPoVVCqMPenWVMrSbrDelXU63Al7
t3he026LWHRJPmJYySeP1/3zxvGiLfXVCMOYRPzk+gH5qUGuL56mnh/ai0dXyusO
87LGAaz5Ru5tgZdtUZj9vGwbgJmAbrOSLJr4FRMbYiwZv0xjfGWT55imghJXNtXj
chAdxKjGZ8NoLjIE8XDDGljWoEQp+nM4RyJd60LAfDyGUPrj4xzGN38/fZsDTx2O
5fvldaAl6gpmIx8qsWCqJqsj32YogPfaMD26+XzxRfhMx2o3pQ9otWc3Y2L2meIl
CkFsQK03mXMestgd46IvMTEeqIz9Rrf6u/jz7O0KFju3eFo8jWyW8S0nX+rd2KSR
jGEVNd6vw7jWiKjJGhd6eiGIDH84A+D1yIbJwf6ZO/i06T6hpQEA3eSMOPml3gH8
l5pubSpp4x976ewTPR3225fkNivwQJgFhKZPLxDQSxw76EHLF7W63lO1ZjJX+pjZ
Dh96HdjgoYta5bLQ8N711KMitkNU360hPPVf90L0a3jXXJDL2Utb7xfpyA7BXWHw
MAXD5tFC57n6dSrLfbMLwnn2WzO7U9vVbhnUGVwwBUCIKhB3gSM+ohi1ZCSRsOQ0
mMSvWZAe562Gqo7fBD9BHZM0AD0MKtPrlIL6yJhlevMG0/yuRG5lATVi80Ghhpw+
YxQQHTsj24C2+1nFCSxGdf+lXN36aAjHY3M8tcyspJv+0KfJOqD0aLU84UfNjaA7
p7VtiTGP7Qg341jowRBT19cSPvbibngbCl1kZZbmem8Jh0hdntQpCGEOhmKH0cd8
dH1gcIic5lB0SXqoQhPOkRom5IvtKfPlZ6fvsREx8/PnGIzoyz/JSWmHgI4PdoKK
UQ3OUyq4Ol+3C4zKlvOpZzpjTgd3quvpOQCLYi3J1xtdrsMObf8E12e41E/fGSTm
TCb2CRvoMDlJTa/iSjzDlq4spk/5VKUU4aPzmt3cl0gzCWDwC+HsI401xYgsYz7B
dH7TbuET9rZDvl5+TSgC9icxfltkU/VIWcjKb6lHvEfQ22gWciAILRcrkylbQz8A
ZFIol707xNKz2orcg+SZpF/wIYQTjEXTwIVb4p9/90miRx6E0wkXAJePCNxCnu8d
duSJ56+6MfLpFEHMGkME7hjjx8cpNk0CF01hOnczV7kGzxjWZ0D03R6kFGAlU3vb
CytjIpdmSPlcVUJTAlaLOTjB44AK9a/OUREe/A8XdFW2gK/h8ORjHdse0gHTf268
Jv59V3Vaxnti5n3U9Fv5b76XfQMwUSnTC72qvWDy6ahmU+RS4Vbw0pZglDgv9TWD
Ochy3VqweJpOP6KQQxdFvIT7gngW/k7buMxqU/1LtKQDyB2fUay4YgwHrsTvTymI
aoXFmKnI9+5zZaC51WoUgJWybij1xS4WC9FfDfS9YXKKaAi7GJrR83OqHIweYHDo
GLzgCYg0qgRnQiqOEcQmt5rne9cAkcJBgOK0oDJRoc+PGXiFYjnzg20SdGOLh6f8
BT/zIlndkOIE6u6YShx8cLWZzqGBxCj225t1LUQ85DQZawSRl7TOffC2mJyF3Tay
bNNOhiHJfE2YV/iOe3kLJbce+LSs+hg/FOD3Z22EBEhJoBo9gEtiqzVVvDmPFZs1
rvxuJTs2KiuOOBCvQKo00yc0Jy7qibr1T7lqaNQL3H4tDGNOCpX47GGcgilUNyE3
C6RmzsAC36WVBWK16vbz/9nbG3lSudALkC7Bj5f4NG8qaE1/zmYo3d62/tACnm5m
Ck2ZLlRH30j4ag8eVjzF67581YpIGA67Q2he39AjDITcEApNkdDe2bOPgcMmQAt2
W5e9F31rG4nk6zUFZAnGZOnpwbL5skCpWBDMgCCskM+Ka2qyJ2lq9e2oWHcl1ltS
H0Aa5qCMPg6Il5gCq6LWEbtwMXe3YHGA4eFOLOf2ugrOVIXSbEmSKnjhuOZMpF6V
6++9EUkfQxlOdz4rd9mfVx63Y84Q8NXxGE89cgp/s3aeTqdmbcbQDruJRlMpaFhR
ipf9KxoKY5HNQlI7wJjWEouVxmlRqfekfwBqddDolX8hZJK3VtEwb9QJ1X4pi4Sk
I8D+mGwZbC6+t3+WVSQA+7u0wHQCshblCbVsFS0mJquBXT2ev07nZzcgl3qhm/jb
VnErKJ2vUoqK1K8GwmUEHRYzRSjNtC6j/stfQLSkuM4EdvrUMn0U8kSJ6sCUUcEd
HgilDmKE4tr/+hWc6vxhzY7g9PLDubxC+yHl1lBTY6u/vU4h8DZKVbk1Q/vjiAEU
3JbcN7sVtby7JJeTj+aWzPVNdqjIVhfXTrEUFwxFll8AdLFriRwMrf44GTy3Jja6
rgnCSJbv/3ocV9W1469+kIADVTtLiqvBKtjbnFFE4ZR4S6Uj7pP5TWA1nF50etiK
v5HY0sR2RocI20MvdXAaO5I9sLFaSDTHFDo4DbGDanaH1de4NCzWy4WOE4YOZ3p6
buB2nofzLbON7zz8M13levNJ80WVi9nPOf1CohH/B18p8Yw14fV2EclKNlVV1o1P
g5o0T7v9OEBGXIe9mEJPjc3ZF01sr/LarHNKS1Jo21zlKbrfyKQ7nNVw3tvrIlQW
yLnKNftwcOT0M7HO/oDJnHyMAZDdtD13QCAG1SVgOV9ZoFaPAs99BzJ45ErLvZPC
FN/JZr9LvtV2/z+aNiJobkwmgTyI8dDBVMhDu0In5kJ7OmmG4Z8GHLfN9lcM7aoE
KEk36OjZidGjKYvuYD+/J9KX54Aohh7H8O1L+fTMD2YlhTO8mnDyadNXuZM/lKU1
9keHSIq/3gr7UwpYzzo/TSO20mAnOfyePLCEHaSETwGLn/LNnq7A0DHvY6DFjsLT
/VUkgqaHKzY9vUszp2LWy21j14FAfBAKPVJnSfEE8LdJKLazwaWjJdWCErLh9wCN
K85vwa9kD4psalI8GERme3wM27ISs6GU1m7HMLr1vsnLyyrwVRLr7JeraKFG2udf
IMBO4AD+SmYrBAYe70pOjm3DMqPITO87z24qq17rAWBBwdANQkw+lo4fycRkEmT+
N2NP+2RESUVc0/G4JrxufcIVGelC77C4eCK2tQ55oM0WYQYeP7a4QBlwnS639CMx
SeWzlzpgXxjAz74KmDnDBTI+k1tR1nLfkkFE5AbyeLXcTFb5PNQh4Y2PhEy1JyT1
KbubPZL2p8QftifS3nD/laPfpFbelK9LiN/t1a8WE9N2rrfeJ+aIDhNxtKkJMvwr
5fZWBCxePqwje/TjDVpdJMvByVlTsvU0cLGGfxiuZvS+fmdPS+OztYqn9l9D3u/N
shSCdvvCCuqyzsAHWEwj8aKZujGPbmi22NAweMoPncCk764xhrMSn7ZGeOs9ViQx
t/L+FUWmPg+oEe4Km5XSJCHq2BKB269ULh4+fP5FSiRhSbLNj7pGqjVQcYcDzzpI
G7qc5HVnwsrfpdkys+jbr+0hjAnRBtvzpHRk2K/XVK3M6iAkDA2mM2fXvGSokBGT
6MW5uEMBtswkF4eXbvd66Pm8uooKZ6gC56BH7AnB+hX1LCgEKaG3+c5S/HdnP5a4
dEOOEbGBPhOio4M45XcNtxJuIHqg53ttT5Z5dxMltXswv3RD/eITadiE6q1MPAI8
W006kEUuE/Y7/2FkPVgBu7Fvvleqvpq53g59EzSI7GtvcxCvOviQig7KP0ngzFGS
Wk7iT5mXljSEHsVa8JysrJ+BuC3eEqeuZJIGnnG6sKmSP9D68msZu1koP7skVntO
d+yQ3lCHCB5tnsa15ONALwfa+jo2djwC1eTSKFQ5e9nWTfupdUgKbFT48l2V9/u2
UV466PGtoYNtDAf+Xx9yPGDPq1zQ3Zk6IImvJDIEXakI/KUdBD+ulHGGHnT6/sOj
9TU5sb3zRJH0lF2FAnxRz139dhTVNBe/cZ+ZkcpFzaZ3fCaeFF4P7ChwG4I6ZJvR
ZAnKRSweZM40U1g1DPWumjriz9rUDbxYrjS9KAtyz260K1aTeGX+bMqmaeFqke4H
Q3HJN/PqBtTwqXv6UwCSmyVL5vemMcClS4OcP33vkQejDCZMioshrJBEPlOzL4vA
Oga0wR1bfY3V0q58zQU5Eyw4seQbjQHOcOoYWs0gE3yuWJ7DSk3f1d4DCkMpFp8c
YKtco9olDgH6P9My5VbZ1fwS9cS9BL3dEMLQcQlVklizsVpQJJJwCJs74FV2IRQS
Jc8tUpyleXHxsKaHqS0iDO8vaCPuso2WQwCBrrKC2VGUDE+XTX2hVz6TyDoC1D32
UbXMDHifAmSIxLypEllXqEcsBqgUqZHH9ZCjc+lavO5KMSmUJVK9fTt61CcH57DD
Hw7d1wZxJnZiO0Jrka52t6V8l1LZS1igpSgoJqGT45XI3l6KPw0TlMPAxN8JE4XQ
ccoIDDVUXNLac8J2yKI1wlTTTiZcCzKalndYutmj9l1V3oxY5+GZOb2fQXpsqnBz
`pragma protect end_protected
