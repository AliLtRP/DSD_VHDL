// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
fbNf26dUR/hFd4wW+uY8VMCeLg+cCt/0S4m++U2uUWf6NhSoOzIl7aSUzWxiHM9QHQxQRtczfdKT
itxpauyUR0zVGQFs2c56gJ+kWRQkD17PbYmhRj6BAnp8/tCwb+c/JSV+KXu14gTGYrmIafMZ3puY
NgTBdWgbkc5oB5NsmqioyQf5/W+elUr+Ig+CAua+aQgYpn0UW/JBaNSfblLLo6YNJovW8ESCe2nY
415krErLSjmSHlfuUEocpqj+xHJqG35VgIJQWB+vXFySX44ZwXlY+L00JGE0tRSDcnI26QL8+bNx
k+ocbG+JJE50O6jMLU+iFayAFvPuU0WVlaRGqQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
y+8M1BV4HKK2J1X7B0uqodm2liPIpbcwfFqWh/omxs5rPBwNsC8d7q//BeirYnfUzVfF29YMyRkM
FDhsMlvpX/qSsvtSNy8Aab5/3uK6tsBJef4aUr3tAfsKVbj4ntreBHzabY1DZHDOaEvLZLc1p+JC
FK21tWMs0gi2f1fUT/S1D7BXXLS/MVBgEwtm987TtetDVN5VEmw5VxTUwSH9gCkIasEo8mdaLqjN
cDGzJgRbnMqdMXNh3G2S8bw1/VslUDaXqRf+kSn54DkMqSHPueh285yAmxyVsYfKHCIck6p5xKhE
eCAptBTNkfcbayzUeOvaLfG7EE1v6KMTT6GPJZ5DN9uRsnpdXBS8W1v4/E6XzjLfbWZI3/1511vE
/nlV8gb9/dJiuJAHx5+MRzaf65nEuqqWfWY2CQfGEdVldUf9FO2z2DmpZr6651UTV5ziJ6++zQRd
QO8vIYm0FB+m4NPmECuo09aiZHpAjIJD+dMnt3Uf2f7/ltRSZvmky9a3nj6TVTX64agmyZGgEF47
Z0/xIAoGyGDrh1FwdNyRoMe6xa9KmO1AMt6RYzVqWrWh2CxPSNKbZKQOb1veLC65ejQ9hCa1/Ujc
W1pawqZySPZmGGxpER/fxNBpbKHq9rB2mwRLKlFLw/yMSbhE7PpK12km1oVxQWiOLeKxehe8dRJg
vZD5vSaoDgSMihqROBUDyBq3zjLsfjza57OSXySEjkrAHLu3+9tg/G5/GNEsKoPEJKSZHFfYzlKP
CB3gum2x9oYyFCXz2fb+1QV9b0PrBgsxKwSsC+EjFgkuKFp4TbY3eXJTlwd/fgRaWmX3JxXXqfQu
NrXNnz0SSVIA3+pSN+3nCHhExIP+vqdWzO6IEDzYkQMR20zG13DAtP4bjlJ73/my3WVE877PHHaR
lEGDSIs7PV7mPQMnt55ibIP7epbWsPTwIBchrUyb5pJbGCapS0BOc/BklOHgOv1evfqUy7oOeu3Y
EI7FcDWX0jGNJ/AO95b0Alm/Ra6o8vKZTNKbIDh1JvFYFG53ufIq6anKfwiBtlNGbmlbaVcozr7r
o68qxub0SpS23a/gGQe8L5SQ5GD61GTjUUwUdfCBtqyqhsmUXuKhF6Lgh68P44reAIQXdbJ6C0kG
51bPN/qb2Upd2/s0d90ngr4m2Vx18Nn23Mzrd6tpB7+mD3craLsmCWsS+wC2J4gdpd+DOJByzRQB
jCYoFsu7hhYA9hZrwHz0fk4val2XeZBy1t6RMHaNdRpJ7cZO5oGyo1QI8UAEPlDgf0xQlWb+SHhw
ILFK4+e7T/0Xf6z7BwTTOI3M22cdRM8Y8M/vxH6DHNvzo3Lo9NBz4jgAZWbauo1v1Brvuyg2RW8H
BiVn3WPmU2DNYrmq8kd34O7AP6g2MdPC15iZsLXnGOfyILM2mIBDoK6lN7bBMJFV7Gd53Z4YEEP/
ffK4oLzo92sMCeiSyYEeX2cXTNo7Mh/xwfTXYXcqFOlIU9lsCRji8SMHieVY8DDVaKE23zOfcC50
01GJUiond73y0A3ikb271iBPc/nNlv/RsYOvFFNKhsfKJVPCxUyM6llupikBZlX2vGPe0fAlGk9T
4KoZKI/qlq4woP/Ob4B7iEtn3tsvCgXoQ1TFW5bGgBlE8DVaObYbIMMhsM1sXcjc6evsjJjBLTIt
HdyJJAlrHK6O1IIwKqPqpQp4CelRX9dZQNoPPC81SzF1BxOnC5QnB/+HJa1jeRq9d9lvZyW2s8TM
+HWsb7N2MV8VJiiy+/uevJJyis5ilItP63zBTgUg6pKAZ9WBZJlnlkKDMHdnjXuVxuG3zGYuRw3W
kLbpgrZzSsVwZBenbzlq3ifuzYmFgNM6iudkHQXgSftoHCN0lqNMi+Zxns9H1XYolbMSavEn8kTz
N0/UcS/Hlf438LabGO8zxDd6TWNDA2d+3tzfi1yWwACV/dNCWEe2tr2CORrGco+n3otqwcxuGT8g
un9S1RK22vsKMqlFFV4Dp3kAAuWBqGSwp53AY+7klBBsXMOe/Rjaidu3F21L4Iwk/WOSzK5dOpuA
o2Zh5cGchp2Pb2uPVYOJcfLfWw91oWzh+dayLnVZaZ+lSWU25PeUFvoxQzdQAxt7UMiM45v+/2SZ
+NmoUY5nUiKcsw3h0z9MB8ACT1uDfDmC3q17l4gEhLQUCrdwhBka4cxPBGx42BhytxkahOyyFe7g
w9tnCf70aV8tACJxa17dauyoNGWlg3N/XP3SmNO9sEsyfpfazyH1oY4ob/j9kV3M7OAnbScfaPjI
i9Oe3nxSFAse1KsieUS1QTXRPgDLLlX0LkJM1UEe8xWuyW1fRdbPQD8PgabwbHUgONENJITdonHW
kOF3GrohjIznwpZd6cNJEdsxQiyGGx9HuFOxxMCVjpX3ZdpH12oN8Q6F5r1hm98s4EYUukS+xmpi
0igN61OC4AZ85JT6VflYC6mvtWbP1220OHtxBSW8AXeLUUaSxGZ04vDrfSsKs6G+GCGZKLQQV+tk
+RBvvpWWM+yzbA2GJJClqeCcQN7FVJkerKz7/izbVaICxHkuDf8BQUgBKlWKQ1sF1688j/4K32Ut
t1FnkXQ3nooob+/h5ZOM7StOdGP2YQG6mfa4ZDMwIA/CL/kB99f8aROyo05A1/Wk9g8kb+mTI95E
Ia3U8pl5TPYR7kUgDjpcPlhnLXHrySpUA8y+h8SEy4ZV+qNgcGW6D30FiqTiUAKpUhCp1l0xjXW2
tkCJsNsG1i/RwXjqtCw6NwcJbHqaibVqzX1FF/B8SVpFtYiGhE5wL3gLJa+MtK0x8F2EWUhrS9t4
AX3wgJAXMpN3thYHZrJj3xx5EaB2KnvbmVS2KDar85cicVpaoJU7cu/BAK70TS8+eL/4QhaNG7wa
OlQNPhsV6oW/v9HZYPyTUTrRtZnY6j5s+1tcobvC9qcNvvmZpxpSxQPoAh/iZudkw8Y+LPAf+/4c
3/lM6zdad+1vKTHnPGhYIHHd0UQ8oM6pouZZHD1Puz3kdhIuIQ6Row7hEbFgTNaBEma8yD6IDvdM
dmi/yoMspdWKr0R5N8IQ9LocAf80SEi42EUQ97LUU5FqiPueQr6ctuCe6KZMJgs5wsrlPTNbN8l5
WZvSo2Q7PXwyzC5TivV+0NimBhtMOmt9h175xIB4VOP9q1lx3Pei7BE467TxV+9SsMaDrQlPkcch
CGn4YCHtFXgHA90IifPhs7vmtLeHjYdQ4+q36we2AwQq3B0fUXbr2LNilB/ED7iurkk9I3oJmI8a
0dH8WM9mWUM3GtaTd6eB2Nn53VxuiB95FldzuZmV/gqlzOqHcA9er9ijNQCumGTGZmFSSU3BKN6l
nF/LoVx2lmgJpOQ2JIl3oUIYU36kn4YJK0R9PMnFydcuZqZntkD532gQkMetAe3MOPIA/eeGxdz+
0FyJFoflCDR8Jm12APBZpT+S9qeQkBPSvWSJc9sOSOMM3sk+OF8AHJzF5dUAR0uyrJYJ3WLeh+rn
uWzbTMyp2aDZptZdsg5FmIlI2TAQAxptuPNiFUBT/HA2Zlr3nlkyHUeLpL2f8CnNZax3BwN/JBd0
uE3lb99S6K1Oo7l0RJt6a88tKYu7ZVDLel3CSaSfuNUCC+qySipQQqXInRau8E6/h9kVxyc7Y6hv
tyPDJGyLxZhixs+j5HCqK5bTTJCZ1q1rXUg+3Gtd473I4ZnoWgh8Mg9h+B5+/nJM2/sdsQV19z1/
KnuPgguo+lQu5Lzl/lT7/2XQrYlqNnbEfgxkAdKuOoC1MbdQMW5rrnmjDXTZjGBeoMd4FBjq5fhp
OIlZvK33qyS4B54PT+EmdbhuyOk/YodP2/2otiXOmw1vBpFwHfv8b81UPLPPRYAn3jcOXZF70kdB
4WZzyV17oBKaqGweFDyuKfW1WaM3TV2dGGQKXGr4hp/wJTvGoLNf8/Ts1WFXWMSVEW29EDHWdyMB
IUwWWvsbFJB1YrF6aOYznOZPgrBtb5Ej8iPsfsSFH4nQJ3j0tKl296/NQFl/ctVGa1slidoa9ayy
qDhKn1Eg5g4vGwGv64lIhzZbVgAPk5BEkdNdSf54AktCK5DsrxkEnWazOAiDEbzh2CIq9GJR+/fT
3FKeoY0MNu8hY9ZMDP+DEt7qQu8elm43JHJgoJSSx69EgheQvWyE1WODQ7EYQ1Xuytfl5ieucCtz
FusSQDFEYxrgdNLJMKD5X5ulzaVWlC3Ajo/7Dp8zAmjr+uvQAHMGRB72TeS7xLAPo9RJ6+b2OgCB
3W8cVoSL3HutQwvgGYdDWzLqDx2rgVFhtuP6flIVtKwfNIRka0OUIGEHhV8HM/g042Lhf4pzXRt4
6j4yaMPqtA3cAa9BSDd1UY4s2x9yErz3tE4VV22kSKwFC4wIIN2EbKe8bhzRUdXkZCIHmx6s+Ryu
vDLS6098Q+BlIzL+/37juVcZWBWWYpy9EXg4lD0q4KWLBtQYQY2Ul0vV7hZpMz5eWO+jktefjL0x
luS/SNYiwfrbwRu+QJbJDqTyfzYnKAePfEsGvIbdGPnSaGx6zI+RJRINy5HlN0kzTLcSq02FQoMZ
ot3uK1qfKX69WLIXDnYqlYJWJhHRYRtMH0p+9uJWjchmqSS6EkBXmpsXu747tRTSoR1wA0qgPWOP
g4xzTPJRld/E6FKeMveB/KYhTasIqLzgkOOgA8Dv2ZjMYVXzwVGdvhNSo6bZWHVevu6dg79Sz/6M
3VvAvQP9s+uqkdf5JVYGv5LZFdNPjcRWOffi0jYiA/zuoJYwi4+Xk6XP9natxFFIfPgFhNMJrie7
M9uaQ6HXFFKpHkL6gIvSqW4YVRsMispVEnDODwJ7deCd1be+9+OvZg11V9dlzkKlBhmWlYvLcrOi
pQ4u0D7w3D2FSnlLvBjcGmVWMBvEF2pvIugUsrejy/eI4KoISvgh1dGGKQLtJ5GxWqCH4Tk4YMXI
Ofz/wcIVbFsNmilNVuIRQu8zcgIVt+1vxdbxMiMnCoKIJcgEUOLW5KGhQYtaTuGC/Ffzae6vY8mn
W1tEv0aMZ8nt/oVRUNHFnunbfa+7XDw+J+tF/g+CiShLvseEHyg5s0cgp8SAqLM3Sfb6SV4VR8eU
Kp21FZcqvGJvF+WjHxLJaN5K6XkIdL2CIFOfzurX06FBIYjGiBH5EUapIO4CL1Qa9XizkEBt/k4g
qh78gmdKSbwkUrQJpNCpAWj+l7uzMbwMeCDmsbOgrQIN6x2l6Z0RE0iPPhPHEM0/LCMsySQQ8ttz
5Psi2JW8UlFgdkCapx7yNQ4Ql2l5P0kXPYw4WNvs2z2DK+ddbe40ou7PqzAyuOyrD3wovEQrkl+X
HXjj2DSXfRBb4ikeavS3ymlp/q6k0WKDJ2/VKkyqo/HpwmBNsOEee4vceAGE+Rf4IdykuSOPrtbp
bspv1t6nihHaVegx4pYuYlZ0ZbLlx47th6+FfXbrYyLQj3gzyAFRc/O7zj5RERvbdeFJNIMoDc/J
4hD0ntGLWJJ+TOjT1QrOJGMUayuwg5+qwhMkJQdwAzBIoOrpLOboZ/muPUwTocpN2Bt2fQKqknyh
7i/ITtsZkbiTffbqYZhpaORq9Bk0v+L8Zw7funQjqlaxYxdUz5X7cMcmrW05eCie1j0YU2aze8kE
8VarkDdRNZyocnQ5u5nSUi8z0Tc9xYw8K/63FELnQCxJ5LmgIuhqTQwFsx7Lzyh/XrIExSwjrk96
Q1eqsQxUBxJ4xZIGOCWjQ9VwpalbLd4vv/IYxHtz8dOFP1MxAkuiAhMHZRWWxUqxdSIF0Js2m4z4
LBP5xTvGxbM95fJWute95iXHFkUyBwpshtx0Dm5rb3hpz7fabBiZ8md9xLXreDupmBrYVFjFF6Zg
uO0w3u2NiU8YOnrSq7OTz5Z+pv+3Wwdvm46Qp93QasjnEBJ5txcJBp5TdYZeFyKuaM/WsJdbb6l5
gJWcNoDjS4jK5AhFnK64b+zGI9JqSbz8rdr1dAt3wYxG+x8pVg6DgwRKuofT08ytooagGByPGdG2
DIuvcaCmJxA8wVfW+O6/nv3+5GUO/8a6EcawYzSkmvHs2HVKq31Kgc5fokRKx61yy6YoSipxVVK7
oyg9Qmboveed5xelovZop1trpzNvwpM85EcKshCy7u+1AHdk3V8CCMTjof+YFr1rDEvo4QZvcSqk
84/i4frummvjK/n2LRefJ2gE8zap9pmUun8tPMc7WdQnIZpBWE7/G/4DRtR0iJa067pSVJy1bYxP
cR9TCIdiitjfLI5mub2BFbrXIt3y4FAdg8zI/WHehQPfgrFQOJGTZdMThjo1DonAXw5n2K2yAFmr
J0zmokBFLSHdncKrPzL8bULT9Nx6/kTGY/qc6SfTUIrq2DbzV3jKYyHsQpzkavTRBzpWBVLWb7Tb
MSWWgh7ckMs7ieYiKGHXBv7nsrqvmMcsfYWsEt1yK/8foKCGU85hlllU3n+0bWB/bu5pxRUtrYmX
YI88Ctwi9WLLlXMM3n+Cdce9Ih8c414HQvwTifAXXqvaea9QJl+oWZ+vpI9OUqmoUie3IzNbc6GU
Y52pJkLEJOaYCHikOCzLtrtB4Crq30FC/0djXA+8AmoYxEFI6egz3JvA6SYIufhq60a9Es2yuQrj
wXc436dHd5fWw+1OiZ6KX2m2ZpfmM95HzwpiQTiVHi8HBfJeAMFNjrmznFen4JO6h03dbkvROG5x
nBedmUPE4T/kAnynBBFs2VrOJ6dk9AZI+BIR3iv1RRXQ1Pou/C/hE4IpvhnHZIZ27rAwI1BDnE5l
Hj7qpzW5nTiuIUlGfu9KTDmgjXnsBJvRVSBYwlgrbNBEWXX/ZmwOQW3tr6RplvC+Omi7i+A377sd
zs+ygnDIxdGW5hqo0vrcpAGEPvhRrJ3eccYeM5u0ZciBMN3SNJGwHa7k1S7hSqpWfJsJ/UhS9THP
5fRcEmPW49DaNwCz50qCzd8nSoBSL25JNBo+kvEHetPmBP9qPMRHyijkA4wwhOGvE6GscCijNmuJ
iGaR6y0ieKZ0nNdOkmBlZwPirmQf+t3LZWUpcqw/1xOflsq2kbRjUSHPl3/SDYq0hXmK3Aezmo7H
QkAj8z9AcgDPql9uC1NpU2MAVKIt5iqPEKNW3xrdtw5wkOCNBGKhF+LRju1Swji66XsL2btEcXeu
nQ7T0Ib7cjzcfhSyOVNoUJiKKp+/YnBOtRrYG5c1XjwN+adWpjvPmhJW2MNJ+4J5ZucpXSq72u4a
jmx27pcHio+yyscz+hJp7JKOsMLjkJJfmchbYnbKFO+SSTdCTZqZWyt65HMwZ9NYJlXzyJY3m5ch
mMj2775g2byEtiNqcmnHcA5Red1T7NmvGPeJ37pU2hjdPPyQA4BbbD3ZGtiBT43quwgKT8VQ2G1m
8ouxleeub9K6mv+vDjsW7se/nZCn/4B0su7TH1Dc60UK12jbGA+dvIwHG19VSJA0V00WpB3wqrSG
Em6PR6sm8VBM40MB4iA8a13PQcRPPH2Lc796utuBS1thS1FqzAodcZ2n2WKI66Zt6e01NfLsDeJu
iNpUOQRNGykCMX5lwW5+SvN51ulWKCj/Uth65lQG19QSwS+VcFE3CuJXLOclamBdgVOIYnEudEyv
NJZn3QRqbZkSidUMI6eJoNpW4VJC+bs0zCutjfddwIoQByI6S77Buv1slSA3jC85L6HczZ1NSv2k
9tdU7bGWMJzgAY4xygQqIK/4AH2g2BMx+jpD53OQtzmkl6Kvx2EeW16BhUP4gYVnR1AbAdOl2tXr
EC/3XR+7mXD6U7alYnzBWZbMzc1aNP1ItIw0IOtFpdsJJeLnXS4E5VHA3+31eiMgkMmmIbPOKSzn
ECdAB0AWOLEU0AXsVCKkYWBJGlNpmUADMAO6K3zsfNM/m9i1tm1/pJJK/iTYU+1t+N6JFY4OfCci
uTRY6T1VCXu/Oaqx6rwgrYjrzgrlOletox83ARRCnGj2dixdPV9fAVL+pM1+rOGJOCiX2qUek71E
4tjWa/BkeBwa5g6PMWCWbL3WVtS361s0iFdyDTIfLbNaAZlE2mVdPArBH2gCToUXCtd+cinHT8wB
JLtjJXCFSQ5y6vRv+B6rB2Ek9vlPdXRRANwWVwoOXK0JbxZIoCD9Ma37JZkUiG20LeJIlk1Tu/lU
kcf3Q9vpvISWX4jciXAmTbze15yxg3AN7aSvQLG+g1AzCeujS3t95hX1937mNHJz8USAkvBLB7yb
eTIpIn++oC8Aa0Dfym/oAHxq1bHIgCXnG+vNkSLyybKTWiVKjAZsQ3xc5i4QfSmwjQUrNjv1pVsA
JwURIa3lZNDxo5/X8YZ9TStWfNdbUOW1Mdcs8qJuYvdQ7pBEOuGz8MIp6JO87+18ui5QMgF5dh12
iZufn41aEoBQ45lCFU4zunsaf7aRrTTmhTSBaLwIaAUrmFitkvS0Ug7BtsgdeEAYKzuVR2UqPtq0
FsQ1KDr4Gu/STbmpOIRafCPX/beuvDHGzkq/yflbitOO5/kX4GUbpiVKkd9eG4KGrtaSqae1lXNR
X8dZyof32mvv1OiKuAQpHXw+4PEX1VaITK9MAHhRtHQzOPra7NrZFsFqIvLBO61pDiaEC54gT3zX
ETmdkBSpP2PsnuTPhqWnA0onFa03Ax68TM3vuVYvwAKtb0tbb6czjUXd7PLx2r1e1MHpYOXIbnfk
09kQ/qqFaPMN7evG9wzg9KxTeadUbE8mjBs3kOQXrlivzWpN0RmRmBXlTdHuHI+mhswFglmHnwgw
rCdQz1BqlzBETFh8+1fLz1Oo7HHIyt7cm27DOTSdEj7gp9I61Da44P4kexp12gXa+iuddhyaCpNO
mTXJdlXDzcuTIsbx0mQXjBpGqhpRvrUuRqEDizOqnpCM6p84M5btxD7fHh5KOpZgLev7QEPww9Bz
ulFc1lXQqkFXP2UHJB3er/RHgNAHfTimXPYglxbBjqTBYe34voU8qUa1xFMQ9YrOEkpYgA2CxT45
WnUX0bOs0brjxhc0pDwYqavTuXeGPYXj0w+wxBZeMNaDxWdmnU1N6rs3M2lsFAjHDglYNrSYKJLh
7duEsEFTh4JDOtLS8+0H1//2vAoIflItDMkff6b6u2aAKbKiZ4L3ret+uw/lvQ5EnGGlTBT11z9t
ucj7sOpVBH32WtcFIyWUHVTEchsMmXXYTsha1xcAM2bjSxQ7ATz5LxoWR9Hin8kzeZwsOsc1ROFk
dlJ8mCuIqzYLydIzpvl1NY9CFSbeDTBbubZkZOq2zlIvnNav4HRvtn2jwtvNsOZfiwRwpAy9KOja
mfulAAndoiGA9nkgNpN054Hmrl0SvT2mXKvY2apRaXStx2k6TCRkM2b+z/8lxbc1MQ9V7/5m3ccY
xBIjCVQlIjT52im0TYubvRNAgjy/5QVcCx06+1PDCFeOyQn8lwIWi4S95EbVX+JwSLlL/4LQDOQo
pbb9naHG4t13nZtXgaJvgxbbvxe/fhUthTpUU22Rf8eJ5P5AHcF5AJLo0OMs1EWx7wfxC7emzdHR
D9ryIS13kZ/w40MMJk4s+mEHl8KKnaQz8nMIJYMqPj6HpiAFY2BMesO13CV5Gar0q+z59zZi2BdS
Wr2c7kVIuMEvc3FXzT1cvdlcQBwEvfG0MvmDQ+frFkohFD3CbvGkTY492ZzQktymu8ntj3NPGNX8
/cmSJNVZ9/gYbA5vsCYwpHJvqeuvhCe9+/RVYuji6slsL/XVXeQrCCJK/vr09A7vBZRdVRwcsBEh
PGenWmYKmbVemvHgbX7xA4a1fhsZG3kQ+7TSRyc7T/Mrg6aIw9nUQ2nEixcqAMytnomfGzvsrsYe
7j4ZaUO3VnuoXeWrQ5M8fGU/wjXLnNfbxX4BJthdvHmKeCI17osuaTdp4XV/7DTEmWA56gr/+ogs
H7YECQs2J9aFOegQSbgoZIXjr7822lI8HFhrkGYnrU7TE/wZydJIYtpo3l3sQhN1cEOffqeqXeo1
vIC3U/CbF3SPoF1B4YsR8CJJvlqwvUBbNP9yDoXJVGhsneJbmuycPL+lnEFnOnpMrEv961ccRZOg
3ON1LaONG91oO2tLXth7fWHhi9Ofb/xe++1uAMH+gkKVE/2gzOzBEE6RCaefkYSixwsvIQrwYVvC
M38+qNkxDpz+f9WxznlMVAkSPQBYR7YUqmx7sQ83e2VN6ClcUmf73XSa7nXjb2glCMUucTLYYRxX
TheJrZ9px6xhVE/45vDUbzbXq5cvlRuh0lOoLtbWXdSS7uXaS9BPsfatWul3kjco4rbXw6LVDxyV
xaXbcMJKNJ7B/BLkyAqQMzxbCi1SLOkFA17sYM+gwIn5hgFrcJV7Bp7ANL/a8jjLnSUQePKFd3q1
gf7J388Lg/5RrwtwXvRzAY1p3RTI4E0+tF0ByOg/d/NfubnVlzMcU6P0335jmcPInpg9FjxtUdJU
ULL/uEUq/9nXMZdor8tTjo0kUZAac3rdySGTlI+Y/TiKReivzGGkAMJvRQx4Ja6+CTLht205mObm
ghDIhwOPD6NhEUEFBAE5TMEYRtC97cADD/RphvO4jl5s6NWAqq1Cunyh/Hvgdptn8v/whxKZtLtz
g8UB/f6F+zVy92eGp4C19WoLcj425LUCgkXKwJBtDcwbAUA07OfJFlT7pcyHUryuGgQBeFR3/8P5
HLohjxaeKBXOXM8uAGIT84IPs7qz6Yuzju5p6VRRPzKaALeGAIT/bG5YgvaTwdPWHPbNcQzraUrp
kxfaJH9DDrPfPwAYfLOabdYEz35k5paynl0tE2ENl5lYCiJlLXQiwKS8Ew8A/1U7NyChk8P3oVKv
Y8uGrVlhKfLCWMNXic53yb+GGuxL2IU3JDQnWOcTjCzQb6b+jJXyosbhjGE1/QV7bNYit7997ihJ
gtpN4PETBblRRNKr+m4xH0DRjtMRVSev/rL6vuLYwbtgfSX5GoleGi/Ve/PvTE7HsVwGLRsGOyKZ
qk5kRjIsJfDj+2U/VE3uZ7/ip+N5i/TS0SMr2WsJKy51BYWYKcz0fhId6aVst3k/qkU/4o4oUcNH
GHC41tgqw4PYhjhNgr7ppI6EX0HGim/Umz6vxHK2YeXuDj3hCGTrAhPd5TYliV8Nz2BRGY34hg08
W2LcqQKIsVOEyF67/Toh1SJiWSZiuVYJwExdxc5koSzTzSKJP+FOrLXDVo5/A7+3MrS8V1cig4do
CC/smlNEs5dulgWpUrWcVMuwJOzlIhUiCWP1q7GN1v9bYIjhK/JD24HHZHFrptkbZ2TgnkJNen4y
hyhsCwehhDMw3TwCVOQiiVA7OtCCy/rezExTud5dGsvslyyednZSOcxTNGtN2v2pW8SovcuIuoRW
zy/MUVBkUjVRCT4bQ3bv3TseRBjm0pDstWPfBplM+kpNf7HveBRItiwpUeqb4qlldapMRzO4gHcw
dFSFDBhhy9ZPVLOJ+/QlqkwET9ZSvhvidKY52uwft3r468LHeFQi42NM7Pv/T0p3CVcY/mMM4imS
gkCGkflKYse+6rI5rT17bJqIJdtanDc0p+3wGJsSja0Gy1dEOi0/AXT/JWCvBvG108vw2/29LYyf
OFap6Ic7wfIq0NaU7MQSNWmaZkeAw7Y2zBmp4aPn9deO4xO1gld2P+ukvR1nEWQlV4M5D70km8Po
1A5fADBPQjkmK8717iX4tsUrheghswPzEdQn3Z7jZGcarfi7i4d2w+FHYREGZWz+AtHXPitHuWM6
qaPN65TkcUTPulhWx2vTvuRJf8RIHMKSP4e8voSYIX/GRtJXj/9d4eCQu1s0e6X/ul6JTo4WyjUT
OqVBDZ/b5wODp8JdMFsDfUCDqSJ9Mfe/pV9SOuy+8SEnOPAejQTuIbloJ9drUixcYuVbHCymmBeq
Sq27AYY9vGoPtuAh05pfkluOcN3k9sh1IM2fCvfVj0CT+5Cmh4s11FQtePKJBZpcArdOD9Z0p2fq
vFEhITtY0uIB8x0t2Z3dCiHR+4TNACskIDKcDan6kJAxsSnbUKytNnIYd63aQxCVH9k2KF/3EtpN
ZgFz3kkdwBKPZLzfKZmW/dxmIzEyZcHLgsbbDu0xvi5447NRdYR6rAllmJU1j5lTFJXjyhrHD63z
F9dfMZjn4SwrSrLhibgK4JvcyQ+MZf+41yfGqju5MfiPOUYkumbOYygQBIkwxtJdp2rieov9GohM
KwXEklY8+LadfFCrB0V6scV0TQTo5IN2IACxnGKwPvySP/3msjFyVmoqp5awGprVPeoW0zTcf5tA
2erFbGGJ05s0qqAXmZBQlLE2EE6unJUkRqlePuB5P0iDoSO+SGX2FTt0/wXnQZwaLtdkpDsMrJD8
pPTELTG1J06F/V6kkw2i1wWipdz06/rYdO8IhcDGXygBlmqPYQHE8Iigygk+DFRDmZ3NVO6eMMhS
dr1PgW9txobDAjUqnHlNQUVdJJkmhn38davVz/v66KymsG44mI9fVtH3xhy5ssc1apyI+t39Jm8Y
4cnWlVXi36sj2WPahU/FinymkJHpF3EF/Wr/qHpyllNAx7gt4h0lJf3dg7+iWbjC4Tx7Umc1mWva
xogA8YHE33ZUx2Y0XQb1sl9/bNcIOhB7T5MIBV2RYhztndkmDQef0KR2NAzyXUReORc+2/Z0WP83
VUelfSviDFQ2Unsafsda0zO6OfyvedyQ/si0u/qu4NWZJncC0qvbj1X1h/NEMmf/pNgqgrYHJsrB
QB4g+T9Z8yY6ygYWs6gnGrFg1OjqnQbDdNGLID5ageCej029mnOebZmgvheZgVjAnuk/hQdgTGvQ
COFE3ceiLLsXw+WZtxbycRdnZmg8cyT/8NO5PzJ3lCWBcVonJvPpIwiBph0TUh+x3T4epn0P1eBZ
5NRD5rCktdv30757zLaOhW38GB72naf4d6qmYCtzDklZ1i1Hcen3zQ0Tfycuy9J3B4XJ+yEyn2ms
Fs6e7uNTNV1yGJmrxg6xZyjICbVs5VSKwlWoHnIPKdQQFo6TyQIOf1pFm6d+zb/Rxg201L8LxvGi
Tkk4i2f5mnn8n0B2kQZrHEGGVhbS692ULU0GNkoL2S7BLVN2UbmGyXHxpllzIdVKYwhNi9LK7Y4k
qttljl2iLMXTUM1Mp4AD8yAFsvxKJ0+OONwZrG65kVYk6lhfVhx8PeaMSWsImJosmYx0drO4Hoeh
BrJTxCsBcBUj65RdoRLXoxyH4qaiyNOjbQNtkh0Raw6KPpZd0tXzf5eMWwaRrpCJVDA7cUKoGjl8
uiRL/LXlzFENWat6y+bm0EGuZHUvHGqW+vRdsBqtub4RTuHm0zewE4YXZTljxcjlv5WB+g6fIXEW
lR6Er3Tci3Mj0M5HcbxovNghpHsUeAnjjsFtKU2tu0O9+C1L7joBDm2T4Svqoc93AqKbL1EvJxfz
f/vLazHBUG9cL7RsYuZRR1uKykJNtOIbaFKPefToLcv6dpkvYll63mMTfiwrqOM71HvUevQyY6ux
REKjNXdPQnJreWak9JvVoo7Y21kMhB7/oKrzrVzLVO6yRYJP9B0loI5AFrs6vBwy4+opnRXgVn3y
6936QIcu9+6CWFogGC58G4pM4B+GPUZrwg9LIuFtogvrZncKeLwYIfSYQ+VnIgDvj20STIbNtQbP
Vt4b/B08MUvIo875lCUdwUplzSWIbZ8JQ32g8BnAOdHsjZP3Fb7X5XNpjK9/fOlnnCPrv+dpIIDk
Hr/ByNXWcD36S8kqpLp5DS8TJl8mx9vowF95pYBKEV3rEkiluAsh5bQnRQi3t5xlffo9oT02zh8s
zLke7YyvHh9h+kL1DanrvTydAOlnfu5Rbc2Nri1Lx10GTrEYc0+f6uHVK7KNnedLk2C6JNlleAZy
mhCCUK4+UOGuXxVUV21h9baV6QZXFSLUDzFdh53rpTRw1u8BZQdaOolMKTYLmg+Kje01b5WhchsR
sbrdU1RZ+lDJGZhVlyMs8vFAshQoCgcJSABk2YJfGBywtbwXiHPjyc6A6syTN9yshU0yhnxRXeVl
Y8/b0yVDzDWkrB994HtxLZ2B/PgG41UG4AEaLGCsA+tgrvvpY+Y+oAHApbZNovzmpdgQncjVAndV
IdJPF2jEWDcPtQGLPewpw7v+wIdREt37KKnJPKXg5NXOFU/8i8rHkBuImSMFesD5Rm6ihlr2tsy9
HtwCScEqyQ+vegSu1qTig2zrRIY6Yh29LJJWWZYRZzW/4OXJFaXrOCdAoRuef0WEhmZJo/3BIwuF
dSquvZqkiz13hOTC/xkmrGj0xljfNAZt0uUVREplOogEiQ0zzK17MPcAKLPsn0Dkzeia99BQcXfo
YdMM3SuEU5Eer1srzVDZYuccKezq3mtyC4kptotkNA2rN46StWx/8VQ5I+dgo8GzvqZvKEbaWMJl
Oeu50iOku32Z7PMikLWvWf2SJX02XkDT+56+6mbzI0V8Ay5KHX0gthJXNZj6WhX8R9JvvW3CZvKt
7x/SVkjvZQqLujcsAsIQuEgEC08mV2pMTifRYIalwuFtJOLhsw5LfwHJt+uHRu23I5GtRmxFus7B
hFvbcWV6CM+3iv2w9cb+uw1bKT6PdaNj+5JYMmO8UzJFa/+neYzCyUrz0veJ2cBON7HDzZx8DiJG
I2eb1wtpmTSSuXeHzr82WIr5GtXuX4P8IoIOqMYTjprQDwpd0JddmhyhO1OKwOXT8CBAVBqnhtRg
B0BJR+K8UDrwyF5NsExQhtNyCf1FJi1Q/VAZYidYboScQpAMPG16vekTPOO9i1SmDeo5K5O4jPtQ
fWzEjR+mP4KaD5Q+b7nTiEDStDkMYapgY3CcuN8LDuvUd+u48HyEd01noMtDq+qtuJFRXLlTSF0e
vtBhwL9+v54ij+sRtyH1XrUAZm4GA8fqrUVTHulTYawzh+eOtpABzdlbnCi15111WdFled3knhzw
GfVAICOmLgBY5BTMs0pNaN7HbVuJGp1bEfB91q74UY6PGSUcU92KUBYNQOXRXifJfP1WrKjUVVtb
dlHxnxZ7A7Wt4VhvsOjbBkKSGK7ETXbyOgfnok4ABn4879myhVzKTfl+UlJdMqk0wjpEuMCVHzkc
jkAUJME1vp81vdmysNpH+osKE8Nd1Ji4S2nXTtkCuJCuUyzruXQ7G+gTSosKfGTRgdOdBhz6JYNi
1PdU1U1haTx0BmpBHIuuW7JZC/edfv/uXfPdxF8BoJgwjjEpNaw/+2tDnhgDhfMoR0Mu9s0pAqQP
Fynhny5cKaSXGbCWEC9AsMsT82Wu+NHgrDlS2zc+xexO/CMGl81yASXxXOEDPB31OT6466Z8tbWI
6FocY6uk6LXYju0D0nRx6/CHqQvc4nFFhPjDb311DVv284Smc1cK7mqF68+BYTckHmtQZ+NtktGB
weSEWUIvEPyxPc+Po8EErjJgp8GA1I+kuA0Lb6rDyjgSODGBbFLoYrdDYjv6AntPA5U9XI2OkMDm
hU6uZachALP9Q/m9wcinYSHs5Ku9ZBAJJS9xBEHTU8/3CCYZM2u9agr6wWHcJUHQ70/3IAcJFh+N
jJ7gjOCxdijV/vQf6AcrnOBo/ZexbkpIuI2CnsKaAojFf+cmYCdoNzfmPZUELdwCFFSAMRXFmHKy
cg9fvVr830fApgIJFcgEWaFBug+Anw/4UcahbwZFOuvJ2apjw9hHaNqndFKQVdu7uLJnOE1J7FZM
xHkC/jd5JdIOz/HYFR8Z55Y0Pj2Q5bW/+DVHunlVJ/6uxaWvSD6NmfeqiNx4wzMBjKm2umIhubbV
lNH5lT2WetL4Pa07jzOgVT7DJfmqM2FWnY8jOnnbdHDK00NUGq0GaECGbYym490Doxm1zJLDAor7
D4e+UwFrNBbCh9Sjmc2JcJoYxiWbLZu5Pmt4zd4JPMo7cy2xf4sOMAFj8Z1YzrEuwM00iP4onkE0
NUr4uWsLv0w9rFOgdG2en4PLVam/fdEVDZ5kFsKRUoVKayfIFQoWpt4xxjF5YvJ7XrYro9WKxZui
Lc+0lvtFqK039FQgIViDM3FX5EpevW8QHdZoghOsiMULH18LA4SInApVd9UMnd617BkgZ/zcRGel
Sk44Iny/7OauE+FdsqqOuwq4lbuOVVLopxEDHsQOQ7I7cowrOJBWpGIP2Pafy8rXs80zunjtdq2b
ouVd0fQS9IHsXO8UZ5S80V7f5cpb2mErvllUk9Kc1C4KYuvU7cEUpzLuLu4ucfjEFUYQYgGv3tYj
gANTdbRdAhacc+sSajms+jtwam6vKP7iGI6+uQHwFiCucUFgkKwFTDmK9kUfeo5DU0BmOtMaOEjH
vTG2btPKxVAWdl5GGXJM1u9Af8YVXU1jiq2qQC30WNakx2JKHNxjKpy0p5KpTUAunKQO4bfKrZKD
XDIyGATSFuYk1QYBseZIUA33I9pk+oRZOEgunSAayCPqApRidFkHMSSt5Dkk0yhzrgZXm/JZM/0H
CtqVSk+hqSZZmqcwsO9icTBCPmMYsXnj8w4poGjvmbYV4l/mtmZ23kf1QplORhrmqalkollYam98
k8jGhGjN9y74AC9IG9qIreGnoZAM/owHTvMjyfaVIxcaaBWqcT16frBvkYBB5ZAvBdGpswITBTg2
svh5O+1C+1aBdx920r9roPgJ1zK5gbJmcO1Jp9jkzB2drXtLAuTGnLWiZXkYT0u2EY5V4pXPjGrr
4eVVpKC7JvaGGQv50IJcwkW43h02E7Y1P5PiRpUf5E4zqQ0mTaKNDuogHi4dX0YKAjagkqISThOH
hjXOjs2g2oGEy8V7ws+zm68+Hec=
`pragma protect end_protected
