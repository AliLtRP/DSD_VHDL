// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:29 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
j/km0IPx205MDaTbCHrChTYOdE7DiqkFFKPsAhFkKwmLVpBBAB4Fu7yj86Xd/3xu
6EwZMB1O6U6i8zQFCDWeDqfA3ZkyPJr1XpPQRXWCY1CGff+mqr0k8K0/Ch/3g10Q
7l2iF/z6p1slKUi7zri80WWlOISsthtxTwFU+2/10vM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10288)
0h2ZWlbVU9bP5D9Cf8/nVGq4PBuWz4VMxlwCCHMGCCvltrkL9Np6E2RGFT/x1fsx
DhDRH42BkqQSPdF/WILdi21Ebr6uNeN8QUTNc8A1lsoYRUV1Vi4C9plPXWEk42OS
Uua0AqIlBq478Bgdtyt9MDAyDfdLnoBL307b+luo9I8IvBiFtUx1akeYes2XNtw8
6FqIDPaDUNURzhBT+9vmQKawQLVtYsbFddstyTmbKArBw6giaNhRfK4lnBZHIVfT
c3loDwRI+/MNrIp7EvtgyUy+8JXlO2jHM0QqVOBsyQLYDI+oZhKnAYZQVzHNVpra
5mKenAkdVKhOoogO+3XmNJERq7Bx3HI2v/I0/5r0WQSNEKAaQonfZroaf7GAeCja
ozM6+ESTxUP67NzSPgM4gmTl7lMTf4RgxodytILcvgWSKyGpTia6ZQcY1tcp3xXp
95M47nwKq3Hg8M206KT9dkNJMMsj+VmqvBHf8T8fTJSZq5yyKMM+FJRGfrgFgMfI
qtZ/WQ9B7qiTrhEHAs/h9lLIWInTpjWqlas+6FfEgETo66aqk/7rK0pyruSLarUD
S3WexGXw9COe867Lm33fulJJarwWczYBJRdHDUnpnhc0b2wcBSsKVCMZc90Y/t6x
qkMDBvkiXR+AtdMSRXGDqc9tZMVx9D6mmxUmmv/kEAFrLmFaSvbMruD6gakuHnUd
udGM6FsU6qqqKv+dgJCcUVts8oFvnBkx8iVbdZ4LpEYWcMQZT/Y/xb/snw1hP8Yk
AN5zOjBr1rmzqcoKqq+dwC6ve0fQxXaMZSWKcq18MMZSFl4SCMRxkacV+Jr4R11X
EfkYdKXpN9wC8y6PjFSuGO97fnq2G9yZevDgRdGIhFM8smUkmOatxRN574A1SW6B
rAyWlASeHIaYOmP7yjKmMN0MjzQX7wXdMzXMDW4NzhwmFc+C63z5f5UMJ2SbThoy
Rk4ckMqG9gS7PDTdcTMGSPFjiuq1qULiw7T+VV9AjJ5/8Ga14OFRzsKUtNrCF5yh
cuJkborwxwaSqjqe2Bb+VpOemuCWXuMj+L52fR8+TXkDQtkvNTX705/4tKKe3+OF
8fZ2kKWNdgg+4PAxPNaCdUQlHaLdRSnOG5/oYMeFkO/X9F/5H7PwxG1MaTIF1UyM
JCTY788e0NcckL8ZwIR/QICa3qYF26ughHhbtu49HxviGjurUIXy3EQXiJdV4ngU
+ukdzg8KhAxhVre79JdfOVaqjY1cdW3CQ7oOkDhWXxIqjxlzjhF1i1jztLecSUKS
UjGBBi+rEBymVzdlNSHWU0WbXYV6XzDuE+T3Yxh1jYlBZhTHX15CLb0W52tb/xZ+
OW9htfzQ2w+eWaxCrJ2t6Q4k72+6qnpM1aMMpZ/w2JLadsUJMVt44LqhSQCBeCQT
pBBuykCREt2eUeKaEASyAgxQBrHNI2Fn0Z2cBToP3R4NmC8wlTn95o0OVzjjo/s+
fAUZjyjKOg81xDYolpSttbACZcZ9K2SgdC+o9iLKX7vaVYTmTKzQ1d26eLb5CmCp
/3E3VTk80Fx09+6GqxbSvCaYH66qDqVMldujqbuhFOA1MX/bxOd+LFBcvBeLWaB6
MEPjHGs4TKwlXH5u643XLxIgnxf9VFTxYWChHqQxRmUAkO1ZD75WvD9oHFzN+qvn
z0KmBxBOkoQI9wXck6tcxN4gguFy3GrCVAf7FkC+6nQFw5zc27ymgeYX8PbYlLet
kVGcBelGfDbGuPQ9WdJq6C9sTQxIDZSusP8zBEmiTjDgEfva/9XrYc64EPSEfLER
0RT071nmKzgAVNA8LpXdVbpZ49O5IAvxXULJHGviWGh3GUp2ATQXdUIefhRt67Db
uuTGCPlXiefW6nvuzmBZ4JAuPo5uNu6OsIbMwAd5FTkwvlL5f+dl36HLZ3jNVIvF
hJ0iCzbEnvKyVawsvIiJOPQl84Yu/PLqztf+sjY3FX9NoIUooAsq9iOFY5SrETdU
OfiJ+c/cBTBPAYGklSSKGGSbrXU46hYOdUJTuBrNFWnlnZ0mJYtoCBF2KSG4Yq4F
CUPOQDN+dmHEjfJcVFIWIp31Tm6A/tZvxQSitGRT++mPCXRxOOwehVWSWZFXDl6R
FDGXghT5b5j8kmJtOn3RUe6pydTuSbuOENdSDSAfMNbAiFsDqVYaH7bdeAjlTAN5
uHm0kF3ctP0pFYo/7KAfZwW/Y82fHVuFMLg85KgDaC/nzTBjtNxU9MHIzkkJDMes
u194pyq802YNbx1U4OWSEyD0vNfUTMlZYEl5jOEeGGNQWydxly2z5ZggJj6R19yw
xpO5zJZhRW2f0K2ieSxz5ZuQrqorYrPdJwpVGLX+HsJ6f6IrhFgx/JCXq24yPzLU
Ga/TqeCASkBaOaJ5ARBdPHAWVsw8wn8ARQgrEC/bdaEtuOPIJVL1/tYZT3sEtphX
TwaMPy8In0IUQAoGHI1eGzi2SwkPcvDDdigJCNvurM4KajQF49/RN6Jbcixcx6tu
/npy8UZa59D2wUEs0+jmQneV7e9UNBLDCH23aFRVJk+xBhyLiMKYBvDvkAHY/Z4M
yue1hUGf7AuxAJ7A6RE+bTnKoqGYp8LsIPmVQ4rZWwz3orcvqohS9MY0U++PNFpL
n9x7R+T0s351AOngW0pOUGP/UL8LM3QyiTDAg2OEv5YfKBJ0jJ7hlpZGVRAQKCMj
SbHuJe5gO2gjT0tP3f+Zj5tW3PkvX4pzCvUGD7du7lIYQGWpr7xGpxfhUshbliQr
9+2XfPDzUk/Hzq61kzNfWjVSMIhDkPbDgAUl4qoDJu+moZWZI5FQIS5FgPLYu5ca
kiOFAr0ke9vz9jfDPHQXwOOX7Dd279fxIbvEq58dlCJZmlQlPQliP5Dnv4bhOlfS
eHs5J9seNi0x3Vou4LHwRtoRoBqOez+9ECUtostwfuxfl2GzJYbyU8eQ4gClZSIO
VqoP6K0hQ/hh4ag5mY36mX/eYHR86U6KXgvYInyWxsAA84tWJJjOeq9UWq12K3G5
obU2GMD8fcZrsz2lAHee1Ws7lVm/6nyRKACsoNk3vgqh6m2+5B80LSEQUScaNC4n
0MuXmDi/Z5etdNY8+t0LUty+vSY1bl2oKlyE6fg4VNdHT1uUEIqxubxlYgPSX2gP
AYid9LLtV1uLs010C7/w2OtOiE//lHrGiOpXjrWpJa6f5REkuQlQXOyq09jWJKqK
0fRftAVlYFmipxRQ5aUkhknvcAMOGpc+5jN5R08A7WeyzOk+S758zr9c/4rCZLse
BZG+VsW+2VeNRbEJ1xTBLioW0/ISwrOYicCLsRdCJPBQTTyVJVpvjgpJxxucEBaH
t9w3Dp7BUjZUBcCN5i4pq2wmC9/s3khcroYQ92nEE7GUtm/sr1mEZenfbKkO7BEO
2sQjYYzHQZLAprwHuQHHwu7IsOptgei5GEiJvSq4Iya8sMYMfEbrafyjFWjFAFsu
csNa+MDZbHmIHMVV1m/MVCX9CkeZSx9aAa5fAuZiOeoLoxwnO0vfQEisy40U4jAI
4RLIS5LKx/Rw8fEAibjUqp/ciwUtTdeVE0RgtovaryyiGraZ4UEkqYplsCIkwF4v
6VUBLm/CDeqB1kSQfNKh22SLkpGO2qftTAKmEMg4J4XtrDP92c91n1Vo71BrCjhT
nrwhZkWP62q1BKAUIvDBqc6iRaaIbs8xbO12onlOT4M1FYHUfF37TQgCcsQWfUED
XLNNXIsQovPl5Ddqkjz+/hk3n2BgLT2jj1LR8vKSJIj8E/ogrsuYwF1kdG+jdyMK
0lptncbYd1XpU4i8liyyU4bqZdF3AoCc98XQiXQ1OLm1G2rouVdnQoMOmmdlkn9g
eYZuJQusMugBHpJAg+tYmi/zeoftqY/NdQEt8p1f49gK+9k772p9ZzTiI3UwG5HY
PiGDBnPPw97OH32NBNGWTlUPBKh9/Y05a+0d/b6AmXura4shEHjRAGkaxaoDiRiY
azlmHHaIiKC5REVFYJYElLYTHmf8E8ZJFMbJBGoIJzUbd8XMm0rQs5el4h7RVzks
f9iBAWOQ4D4VuJ+pUbmHj/6r0Q2QOVpwZCEtIHSoozCTs1axo5ozTrQ0xcCU38BH
rtAO/ciKFK1bBwpezW9zUA5nnOxoz4e9H681CHevGnoQQhmIKrGxghpzASYGp4SD
6JI19DwSlQ7HIlXM+UbIGW2bOq/UpVkRztpSjhzKJbtoj3EJ/anTsBhTHLlHsoBA
S6/O1/IaqJH6P7euOYc4Fwop7tivo31bg2XiWF80qfU+N1fet00NE09zYHI0pAGo
etcXnCgwduRprqa36ReghB1lZNEZq0Hrns8IIu1ex23p7pBwq/VRHv4JDnGTXA6T
QvjZNwLI0yYFYBFVyGvnkxT1bbu7whNjGdWjtN6kid2uUqYxo1N0Cy27OSBfpj/3
VNnnaH2TnuUc2Fh43wWRgzC8S214HkzpJUiDUdyq/TC98vjVUT3kR6PsBFXrGLpc
vbFwSSg7CA91Rw3AwQK/NEMSmKqD/NwotjwwBGDFTUuIqQK2iqgPGZ9vFypGjJZ6
atKn33HUeRVMXx6z/WZzSAM63A1KRmPnrzvv9gisLcK4BnZR4v96Uxz2+/F7eUL3
7GaC32AsrjmdxeSShDeZSjNqQ4nYBNVFokg68eTT1yTmjVcxxSZa4TUY1k5yyWmn
OWFvmsSURl4M+dWPKPJ/wcWbbaU9L7mAlGpe0qQ8hgj9FMtL8tvI/Ga1/9ukwMsa
hScqPszK46hL5vGYNHsWZHE2g0bR6RGE/lARfPWUd4eEczyks/TCbwSIraDvL8tj
/CGBHXOETV4cbXvfuDFkyZ2WpeG4be2IqqMk8+bjjQ3EzYVA3JMdSg8UmjvxGqjG
UCw84+NTRxuR53iesfYh+3pxAC6ZaCJEHH8o+yHu+Y3ktZX4fbGOsaUS+Q2f1PKr
6+4iMYR9RhBFRiqZU800siGsUV5vYs56jEdYp1NAWOD3q+/gxRyiMpYdMg9M/HyM
gjxh+TA0ig/pNVWFIRxdA7Anifc1kVzlraLjoJIYEVR0o1Jvl0SNoG8jzZO8FYJy
9QgfjvZIpXZTn15oUK2+GJz/iPrUljteH8r0S0HxBrUw4Gr+5p0RfjLCSG2pgMTi
gF5mG5Zdzm5/NWLDNCVCv9ejbmNQpIOnHhQdwc2Gv3Pj1RZYTAOFhmNML2IxpK1q
Rsfd41cLZMXWKmRTjrwA3fPUWIhCDO4qqBz+DSha7uqqKE00E/XfAKNzYpynMY2z
1RXvCAalTWnab1o7Txv/V/HiaPvYjCXAsIJ0hmHPWwh++uWaLDFUtedTcEKCK9X2
oFyEJlhAk2OPbAs6J3SX+RdjbO1H1DkFMf7/781xnEQ6G8Fjs+E6K99A/OEhlAjt
R3Mo1nzc6CnVXX2v7U9C3ZWwbKqjO/20UdMJZhcbOtpmaeKhlh5YgJK7+27VfMkz
pYU8TBt3pDuoaNOdFwPqMuT9FHqzO4jM3QSuqXOCt3UuDV28sI8uqNp1FU96qlNp
lozhy+zrhlRGvTlhJuOkcoo+liWssGlTrygFkfAI8IxysK90caxrbqTZ6L8vJ5+k
pLpX8vfeXOpbfcGGNOBBax7CdMbXfm0g1uHjcYSRLEFAsvVzp5Q8bdjmrm5JevAr
EQTHuOOKNo6YPsFAfuphEQK0bGkzdC/jUe8Qo0SPAhADkGbpgtPL1RuZjizqbp6c
V2z8Lz8sh9HSk33EG/iTqhAaqygMUS3GRMd0LjJ1zCATfMjnIRxyBTUXj/w8Mnw0
JCWbHMzs3GQ0MzUkTuwnlGZWJWeWTIbx3ZpFzPQbKbSeXJQgdvCRgudfjVuQEUNN
93mR8Sk9XedYYA0nROdqqKL/Wf1o2UMvQpG+2Mcm7NuuMDb6i49L8uXuyeFKZ9CF
Itu6SK6sHkoh7E4eJEEYk5+SuynmmWVF7HAAzPPyHgqDTkNd3ViXFiZXtOSBRObY
Z94FlZk5E2OdsGNcKuq9bwcwDNKq5W8NYBzuVtwYV8vYVAN62k6/0vw2UKQhxI+D
EzLZTMM0g5GJqTAqV/T/KPKvnYqOjkBnpk4XHRoN8q3DDy4ItlaYdnUDItIERLqd
KVhydYWKBiUBmHIYbJwVM81Oz6smPNz4ojZK4Pi9B0+ovRlIW8aeKJGan5BJpex6
OujTbAvTOnE0KkGXDgtnSkRX5EoKIkY2c67AO7oNGdjzpbI+/cpXjvZBDFyDv/36
aF9fakdhPKCKG36Y4uNmQp3KuCNLU0WcIMUewvkCM62Fp0x4Msssei8NG+cM7hZG
Jgw3AoW919/Bc7bNnDD64Ci+CqVIjiYUoYRrxmX5vbzSpP61uhZDGiPUaSRS3OTN
Y5ga1sG4xoJbvcWXatfFX5w+oESKuRS+cL9rTIzQGbjifa6Zz6+WOrT1wssEHCqr
LNXil4AaU+bVOWPuVo/J868DDuRDQLkKblmAV+I0D+OWs7lSKBhEBRlmo/HQTgSB
t7WBgkVdJQ6HQSG8OmaPyq/OIfLFMM12l6mgH6NB70wxO1JYlAqumvPvgN7rvqZl
rnHxcIonrgD9MYVzFG0H112yAnLBl4cR70isr4lrrj6tU9s8edUAxm9cgFfuj7ZH
9Yyg8+fytj/ElbV2Xcxf+Hjx4HXKEb9jBaUL+vNJn80+xAy7bwMWy6PTsa2MgLsu
436LPDcnLrcnXk62hS+AswWHTuh8finTZl7vgTULdOizJz803Aptia3jTQJg7YzD
PcfPG+U4vz66Z+pg4dvqXwLgouY4U5QphgMdOFVi2zSqM9b6MOW60feNiELONyRW
SqFiann9ykYawCXUB9XYwyI3Hodw4tc7wGTmGdowsLq6AmqYtKG2nkzqrMtLeJyC
V1D29eIFiMAFFagTq3SLkoYJ0TqoyvVxgnB6e0t81h8U+Yy8vosfDWmet+/dgNRG
lV6gL2uWJw2rQWexKcOV19UTCUFV1lZTdZWzdJJp13fWBpfX4SxMmGNOt2smumOM
H/LDf3ZhbHgyc+s3lMrAgLFNFx78XZUELu6Ex+GDACQ3DtO7rATGCq3PMMupYMth
tSfytpj6r4SZiq8A3qXA4D4aXkAfjcz7jO1xDZdVeLcpaeIGP/eUxHaSTGm798Vc
haRZS1uyPkSrY35p2wBJAWHfnACVcF9s1PzZLMto3Iu5eXt2C/52UZ8o5MFut7N8
sdcCj7mGOPQj1I4KQ9zMyBtqTA2azQjCYxlY2CpZ/iSI9cJvSAqgE5lHGwX5EtS4
HYY2SoVumWU/q8mdK3zk7YNr62NzpqcakUZGB5FYieG9QuaIrqfVG5CkouhREyYn
csiGwwtBCWxSzL7+bo1vwA3JMQ0zvUaMa140Pi8b26bMJWhxlP0oidjnhyM6Wf8a
Awe46blFOchYoo39guAWgKjufXIyEkJro0W4FN72yy8uJKlwof/dRcAXfkBJJ5TZ
fFlCKjFPatOq9hws5DiFQaVBMTQ0eLDIzxXsvfmLufL+3gwrw6XjK8eqfZv9AWa/
GXACtXUxvpSLMHn2foLW8m/lo5ecQvxNO3WQkfP6eaGqScd4B4KelEZSC1le//T/
b04ibIkJPswyETIZqBAuvUUXSmPY0nR2zotSjZ3Z9wORZNT/Ce4n8NjocKQy8ILd
R4WtOBkys1ZR35NJ9z7xi7NxFLDFHMG0QVYZlEroxKQ8fvCqRfeCVUaJJ/hMgJHW
9DMYi0WRLk5FjYqs2rno30T+YB2SxFdRd+vIeuKkKk/B/Cj83NydtNejlsDCBRmr
1OxNfoekp/gdg42bP/xhS96YEqCiB1iUCADAYOfTtLkYMoq5rYgaETZazCodg9R+
JsMtQWQ/B5y7P2YGBeRQvaVhVIeZVSrhcOuSm0smHzr6FKf1OlgxoJi9fMpoQIJM
TxvdvwmCE6gbCQqXwTf7oO9FjRKjF1BwKV7hmCM8+0W90SHd2vjnHXkl5u84vuWi
TjERltkqqIBhB+PdxbHOeo1Xhy/16/pZ+mtH9Rog/bt7Rgirb5pIu96VdhL8wUbt
/AZczjhsKVG6qLmv+z8v6vjyJIscZ9NSbIwUkh/gZt81KV83vCCcZKFspvg3vQV5
lwChKxiI6Ci/hzsPrW2Alx6xuAmaXRSELJJtmQ06ezxituzijTLwjC+EFhaPArp9
ix4BOWzv+sIuULbiscEoTfuID7oz/40CJZ4dDNnseG1jkitwqAJ5fn1Y1xI509no
5q0/KK0uRZfucHziOkqwXyANDi+P2GV1DNP5/aUS4YB6ikohiDB1DPX/JhCJtGjU
lP5CxokcorOL25+2ppHaDPzwoa6Gh6ofpxVy79bO6Fb07mevKO+p9Q704Ynsv9pe
5Gs2AF82fv5ud8PTwc3ohqjI3yWMVl0jwRwEKi29nQGUbYctFA7IEjo0wHuMx1p5
/HVi+KD9sGsMwGcUsFA1qheKJsHffbsAhIuREm+FxJam0N3QH5BOvyPxEq91r9bj
o0tdILyK+fCNtSKKnCI416d2tm16FA5SDAp+/DvJATRl3ffV4gBoiAKUZsUnmAxf
eGF3jcj7WkBtCUX8/LeYQ2rI7NjzqL4d/Mz0JbatK9f4kk1dzR6x9jci9xaszMlH
SV3GtrIvk6FHZ4/aDsmKPZT+XZ1/qB4JJ2OlMx/J8cm8E1t73bRFzhr8y42izIL4
82BXe16RDe5f0KxL+zuPGOiMQ0a4g7/etWz05cUAOXxt0dZJCGTx6XzEADIjICDu
GwUJDnRIHDic3pa03lF3dtMWfVDnH1kaDKoYGnDagS6KmX1yb9pJTjBwf+RB9XxJ
wEmn4bn/Kq+UqF4UFYoFcdnDzUaxo2FqDD/qurVC6rlMQ5zP+r/DNJ+RURsMvqyy
1gN+O4/qObdOm3lVO0Y/qa5FfKD3BMzWXY45pqAsQVs3guk7WWRqCN2vwVFgmvwH
BVPhUJEwVqz6sXXvheKg+fLJk9lHhPD0OcVbcYI8VoDVR9mmx9R8KTQ3foaHjHd+
4Khwj7VvRpZrnhTglNqE4Xu+9sD/dPeVaDa4wQIkjDumuGAMgqqUnCoUf/lxg3U6
CxvXYedGsc8VxRtg5B6ByVc+P6vpYkZ4yOiACXKonT/Abwjbzdr+pS5qlNLzRPet
CmWHNmkmVVMEm+ke4E/bCagx+1AVP73w1jqpuSAOnlocvRQ1+JdjGI2JWdlS3b9V
sZVVojaMPUjC4IJjIZ8ZbX8Km9piChvc/lUpoQkC0UXFtmd9ZnebUhY1Yz7uKpLR
5967F38wFSB10hMSMjTUuQ51Np7c+ntR68Sr6B2jrd0IBxPgY0IpTfYNcGGcTF6d
86nZkZTT2HOFpKMoeKUGaVP1wGXLQSni+9FpBfFjbuNcbrmHBPtiSv2y+avGxxQe
QXg5WKg0jifjD5gqGmDAWuPWs+x9EhCnMdkgYDXHTNYKBdqf9/3j1pBH7/3HTT9e
60eAphptQdUB3ATviT7eIOYl/XQ+qSthYN/BQ8zaIXG+CRBlwx9TNz6e7ptDPYQw
zsE+PDVkqypIVH6/ifdjswTS1OMWvGNPGMEWoX5F53SdOvuICoERrljr0MIVb4EV
Hi/TLPhavCCHaaOULI3kbTvT9HhLmCLCimIFBbrhNfX/NPZpRZ3/hgSQC78pdxgH
H1lVxT84E/GwMbbBh/V43BQty1gpcAlPN5wQPZ08QuFxgDI9Wp/qtm4B5W8JVCQo
Rzbv+pKvA4eF1mozboKwh8k6s3RYSnWb+M9yNXiCjPHAzzPgtueg8p8WRJRt6ytl
VN0o13MOi9aCwMOhj3bD2BlQqo6LhGQ9malqCyOezzh5qzWStQJZwml8i7jQA6L6
wk1rW9Xs2/oVZUDGEpUZLr8knUY8+VRBldsQagaBKrWaGpbZBhaoeY1dsGzTHGWh
dq1PaDDobeJxLcPuwmwr7jYRsAVm6oqXeCDyAK6iX5+1pShS5K6atbXgzaeW0UT2
J5i6jeoAlrgFpAgV7zCEDaFYJTZyurv6oowriIGON7ynAPH2bCr7yEmMrqzlY5pt
hT2AYXEPvotfbFS3kD+WaSU1muvuceo156+OqO39O1zByLx3TCYwdMHAnrVHgtHc
sMeM2NGD2Ix+40CTvow8/2r0QaBmiOjwnLQUrM9wzDETkotbB4yIm5b9YALe0gX4
UCq0b7tkuovl5+sfXut0/9xfFwewoUInxu7tADGxLPGYFyhOr/sxPlJ1FLfWhzVt
pNZVVKBp3UGsnhIwRKIL2AV5Mn9z5jqzCQms6eF3fXxVJHIryRr+8ZE9UvBo20T1
vkmbHSvinHSchpa60V3yt6KcXt3WjqQNs54VZf/HIAU+wiOHHfHRnaU4x60NNJkM
7dr5K9AObHxwvoE7ume/K5OngKuo7DsR4xxl27vmiTquqNpQ8/ubLKivh7aw3wQu
1Slmlj5wDn0QwmMGey+HfciF5fy9Lsz/di5oLfdJ0Pm7cldgO7amQJo4JTKPZv8t
6B0m2nJvwBD4lKn0XL40lE2/fL7L3V9BAkQUJ+tV7NPHpCPdKg4rD6Kic0RZakH0
2qlyI+Jj9QFcrqlBmmYo/izGCO2R4eSdQpoAGAMzbLpeh2c+5TkVZuw7n3I4f3Fu
FKljgFqre/HsSoHfKdcA1Thd0zEjZTfwnMxykxqTKk/yuHDDDZqsykiaihc6xHaA
710+uSDAgPx0UnWbHBASNx6P6D+4kpkXv9WpTkMn3QCZ2dn7RSK0vdIfcHZgeHIz
mVTaUNE0S5N1THm67tPm3RgRS7aIjU6r0aYy8A43J790ikHIljSLAoY0KLdX3MY4
dPzxK9yY1gU0wKuwD8jAfK8n9j4NJuw4FOYVGnnWSuJytskrjvkZ+/WrO/F9GGRt
pXUDm7lv1l1oAJmBUwtbGZmXvJoffdcSLzPihjN0fZ9wc75IaAJfbJAmaPiRt3P+
twHkYa4wdNDDhgw/YjVXn8gVdDBaPuTwc8FJ74DeemwXOxiGhKLE1zWJNjhoJOZk
oYAk1Gf7sSgPtOuBW+wt6g4NxzprxTydqlJ5irxPTz6PuPgDcOzprHHhMYW/aPq0
j0VqZCME/1agI9L9ru/7ns9hZdVi4IrzbNlYJvd8HOo5Q+EePJ92uENQNTKThekp
NfirZgxUzLnusnXDwx6h+LZRXnUx2PAhiY6JJjCMYX+pGKrNh7n5hRneHDe4b7aP
A0GFbIdyqzXWoTWL1l+ogzaAFHC3u6qfMdhMHhe3+aLkqgQE97Yv74D7St4HEeGt
/fKBAZz3w/lFPicirkrTBCWe+xM4A8j4ocjWckpO4RWRLXQdxyGl7PEu1d7v2XX6
9DCJaZGX+PcUgyzen7E82bnRRwK7dSiEWZ3Y8wu2issLFbmPL8BlJyiAU2q/lJ5R
keCd5ksni5g05W9QDtrWWPZq3+spUfp8Fovp3XhdyQi1DJRYDRdynPfB3EWnvBRX
MZLR3VVR5FM6SHAvwGNZhOcNhR+YsbmKlSX9QELsMrr/AyCMOFYOlzq2h9hcv+X7
VvK7I+JbODAh0ZQ/DqJkHwJ/hX/VJZCRIEvFvb/HpYus6JjNFyHXIOCL9G3GzQNn
ZavNF3zh/NDL2dB8IKxnqfP6SLa5IIOQtO/LeG/mhgJo4lnAbqXihsXRz08me6AQ
zHhYXU3HClEwRGJVP8UjXYLBHWc8hVkjOO6lfs5X3SspEvIIaRwXY36oMLOtED9o
14ONsG/mMH8344fwgPYeAxvUllr9AY7DifdlpUqNCj64ONQaTCnzELmsaQBS224+
ty1mFf7sEPzsixF0CkeZglKCWmaykxdmAAk5WXCFtW4X1UUDV8VxIaCwv9yE5ZC8
uNiBoQP58KxSybVUQtMgjZIQnRIkILRZLoDyo7YpGb1W5byMo9DnLW8+SEdDnWrn
kJjW+rK6noSYdrBp488yS0IxzdYUoY6H0FnmpWhZtNx7RHVn862D9N2d4EuQ77En
jyqrq1rG8xxXtwyLRIRKN9+O9pRFNRRw2dTm34UUz1YERUwvAZ7M3Qdl1w+eqGtY
O7BMKdacWsyLWwI33RiZS6nOVVX4Rkt4P/0LZ0ILXG5ZQM03aRreS/FOxHadUwfC
K2+hEAR+xlw+BTY5tTf+CCJ2DLbisLkANBp6s7JzwdzbUZFa6dIixHCIMKroUO8U
oRz0vy/hTstlqy/dvdhma31dKw/n0psfvIVtAzTk5oAJfj4t+bspFXd3jnEzYEhw
sgHV4tCyixiH9rJdUvMes91eyL4OCznpnBB+NUgQizlSEFw8P/2pjE1wHUqHM+HJ
wOQ09FHHjdkMqM7GTNFXPgZ25GKANuiDzWFWTwmLo18kojI9sHFXXkhzQEyz4WBY
rGjY6LwGOsCJvIqygov0xUiO43hXJDJdNNH6cyGsS4PcD84uK2PG+IHPiXEWsMjY
Plt/JnWNtqlLNCe9mtmGCT80S6QQqY/kSPbjgDL0suBsY/9wUmkHYGs5cKR3i5CH
zBpki+uanWyFBZmtVT4JwdNwrBkG2DGBWR33y12M3MXImhJ2D0QoRT/yqHAf7aCr
ddpajpTKbuOucKTkUKidd/4Yvrlr/sRnFUfzUaMc0Ai4cd+RvJAI1YYoZyCtYjz+
eTlDRMBexdqjOcfxtH9h1+2qzds+f36N48zqXZ98oJVEKr1hAF3OmMl7UNoGFPCA
ToLGQJgX7E3EdEhvdh5l9N84rM23rP/tfpPjmtxTk1TGJX3qFu1XrC/VG+Fd4jwj
xdSbgXEo1vqkOzPY2SSHH/LFCcSKMoSAkqV4ICqrMCqITo5d87rPCIpU2IbL0Dro
GuypDdDMwK4IEW3WVzFplB987Go1bWAJzRkgBrmF394SZ+3Nc4XxHcDHNSJjr97W
v2TQF9YuIOfAUQDIXP1fFUw10OXULqPTfg0j2+qykvM6okfBoVXIUIOS7kipLX2S
BFEsZ1Cj48KuMgdW/yiGHWXr06W1kWQ/ibW5voycYiqvC1bzv+tkf7Ych5b/0Pc7
h1Taa0B5F7TrjK9ZozgveW/lTKJvFWtj24MZ3SoFSiSV0cuvXW2GPjnNj688V/sH
OgED+oWiB/9+4igmP2jKxOn4ZFry/+YqAq3qYmSrn9qSfxH7ByVd4+CHRMzid2KG
coUssKsMcnMjM+s+a+kalJwslgT4TWNlNYs1mcIoU25yw1h7lLy6eOwAD2uzBF9p
RnF/2lYsj5cbUY5FZO828NcwSI127n+UzgRGIYdgkUr7HhwC9g2aEMreAS9IJNL1
leP5sJfm77PNZXC5EPmO5xWIUviK0Mdly2MeXQ4YCK3o2szEx4N8yecYI6Ck9SLU
8ZM8wYHdIHYNoWU1uWt/htZWgdcEIpIn5itxtK66Wa8In9PAeY4RRTwJ7GtkThSX
3LQjvKwTSuKScn1xlDvdHnmBG2ijsiOQGYJ7uCqhqoz8Ea0ChCGx5KTX44uUqS+H
fsnYI6nL4AIrjZ/mjit529ekvHAYBV//SYQTOEmd1Oj1qw1bgY3wl+R9H+m2NiLN
EHbiYTA/qicfzLTYIDTVeZQ68rwpTs4LvNL03qkAK2MsHasBRmuRHvWpRT86wGxL
LJnmYdJvbDunTGTqsZJ8d6ZVAgWfTNnb8RdCnCaYBKy/i7SwZIV8GrY17Zza8b9v
zxToBTZ9nDZJ9nn88hmJML9lKZ+899WjuJkgSvpQ8KI2w044GtUDP2AWwZ5Zi7Pf
qwBf5c43Tw0IXXcbF5b61eczERNU1f8bOSht2AHNBSig9pIiM7Uxzj2d4gGj8prj
MOrj+2VyX6KwOmDa/92Fxw==
`pragma protect end_protected
