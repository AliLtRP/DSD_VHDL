// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Ivm7DV3vqKcnGHWKqKS+h12ukr6WsypuvLqWN87acljJaVyynEqTjFruFE/f5adtYol+DMzbL2sy
4lR2iVPLAUgfPL6s3ndWmn9AGizyI8SSYatMRFGF2I6u8PM7EbKAiHIadMNv4vlkLPjg8K8dGmGg
pv+8HCC+LD7212HgYbNcIsggwtMu1wpE5nd0lqGDHyEKwZUozhNzVSYpwij7eDv2czRTuwz5e8zo
3Q1S25ZDcZ4bM2o0H/7Qd4bTfQVIuoYliCvflnBFLsaFQFwqPxhO3or7QySvWZAZbeTM7KGaiQm3
kFR7r209tbVEzMWXjUV2TFqt1yvrgB7+0zFYOg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
zKvC/0brNgYOyLkPzMUAnbwdqY02DBNcdc1uneUZMxDHstpU0sBgAElkirG94yizTM3BVp28hAFF
ISG9JZYqqdqAiJkiJetZX+SgyRq1EQVG547bVlgh1i2JivwB0oIAWJnrgMrvxkIYbUO350fNKY6q
KP9FPQppvvMuz5xixTmew60WG0Bf0S5eI74kTpSwLkM/8IXo1L+yHdz7Qt8vMekvUTCklwjyMvFs
HQw9HU32A0g6co7uG0zNO5ND8tBX1heVDL11lqiW5VWTSEKFEmKIS9GMHi5eUKpkEeR1CKvTxYvF
uHntupK/yZl+KFDtlta6HeRWwotLHczxx3f+wkj7HpBs50/EecM7bJwZ6KGVW2JJoUA86tQ8croE
51L4U6rEpP6w62xH/+q0c2w0IGsdWWc84GbRe4qbDqYubE/mW3CfQORCGEQvyrzz+ZVZrJxRlE8E
g2wnfSsyLsFO8yOArceunP4+YSpQBiTyrGBnxhExpSDBA1U5BzAZHMwp0gqdsgYPVWlqG1GVvs4T
kWjky0LGzT/uY7GyWW8PURshjEh1VI9XfZfz3AtfbAg0k/Ho67AsEnKkUiF8vkfuB3liTZ1Tm/IU
PZj/nm/adkiKBEGAtTryMjQjJ4P8rJfrGs9LVxYvSR5FMZPobL4n7lguaq7luYmr0TuYFfz+g0UN
ZG86ZGGv4ekyPyNCucRAoB+kD/DAV2i40EyF8YURsz69wGcee48gK753tCMm5Gti5HZzAP7qJxrS
QdfcDBww0O+mFS2pjUiQ7Gb1osFd5n/3owR40KohVPwaavRaJrkzWvqn2OzwlfbS6sL1TCl/HInh
ikjIqAXRhZcO5opRE0h3ZVH/jss81OcWbWmQ7leueVCCTQ7iMEzAhwLA0Y3UlZCiyVjHkUMlN99s
41PayVMw2nmCBH3q6d3UdDO2QfQ13DHJGNG+pSwYkzWafDCiiLXYO4dlejPAlsQ7tJG/rqECEC8P
7rVNMKpCKa2/Sfy4ua1R68MCm0Xt7IZa8mM2pXoX+/QA/Z+y8FOw8j+oQ5RgJifVutIRcUpJIv2Y
IDb6PIxpcMbV3aKW2iYTuYqV88sUKOxl13gXGnFPD8WvwPbYdjowFFMUTkb+2DKrEMmnNxq14aU1
/xezSu6NwyjzXJcKzfINho0yA5/yVqYmY35ieUEYJq4z1pkLlloweVfI6UivHlVNbU7Td3Cu5gxF
XvhiF6rSXplK0Di1RmV6r2QTjeltbLqgSuJkWzNIfdKruPjQSey7kDzSYTjx2I4LbzbQdDmRuX7B
KqMkzSTBOkjBN4i1kU5PTEft7rK3svh4jV86IIhtvI12GWIiBmzG5NUMwkBAxazOSAd4ei/8xacH
wgP5sDNU1bbLq12Uoth+BP1PkUsKujOS5ShA94NxzynSqR2znxne9zed7z7DXk1NgjYFCL12CdrB
oo1blPsPlJt8oqMSJ82mQoLoLYcpDXvNwEDBzCJnUgQYh0n+Ga9aE7BdQez9F8pj7X31+FUHIGv5
UdM5HMZ++L5y5N2EQa/fpo4AJZCrRhOhnCL+gg4w85iB7YiFbEszT6sSCZYT+4kK/aL/3iHw2G4p
X18k+XS9JUsr1dTDw5t3vedOhveHixohgnOXYqs5TL6difB9xrmSy82R01vOKFJCwahKNRp19y4L
PiKnXmwKx6JUu1QjR14NVaa+JbYNI4AePxHuPfnZsXvkQ33LJ+y02i92SErqSpyPQvZdq8lLi7L6
9NN5A2gQa5kRd0IoUylOElFzdS6WpeDJQbAdyKAgcmdY98Rl1rICUSyzZZHrvJyeLsXMa8rNMTLJ
RyRMHW1v2ealZU/R+D/ZETyoC0PxNAuvvz3Ma00XRMpjSscK47UMV1jUuJB9zSPKxRvapc/b4iR5
KT0004UTwGZeqe7vI/4sK7cQMU2+uv7/lSfYNgYp2eibWPtq/3sO0KoD00MEDrgTNSST0GnMxAuM
c8b5pTO3bzEAKWUWiJhhdMXi/MvnbOHjsyvkhP40bQdOf9bkiXwTnMz3QbF16BHRg1K7lwjoLZrf
0bf57VqFxvlM9W9ePzwHwcxA0x6pf64Ruou9X9g4Scnj36yXZkTB2KMhlAWOv/m9LhTp7pC2BKzc
Eyj4IUkqfw1VQ4tSU2CrPHKkDVbTZASNGvJrdKU2xNr61x5EqQqdHH5odxt7UNSQ3kDPDAdtYFvG
oP8zKFI6CvXji+y19m7pTCqC6A1JcUL+28r/Y6GIszI5Zk20xqS+09WbiVsJKfhykaJHihraq4BM
UDAXPkZO4AHv77+kvEt3FRuHbjrAkcMSKg3vRevnR2PU5x/kfi2f7J+bKHzVLJZx+FkFxXtDkz5z
YtVw/IAyfd9jJH3lP3xF7e7pwMQHOo9efwOMEzADn9tUS208ZYMqaJyNDZORuNYOp1vYIW5aIZTs
Pg0lLzLpvhnJVm9Hm2byrMzXs5l9PvFmrmZYg3gAPnlWZoZKFESAe4DbnfUQAsAG0IikYIy9PXPh
md6pbMzELgHYvmgMp5QEZ/5Te8rl9J2Fg0BUT6FuO849smd5C+DFdjnq0lutyY8cH08CeU9mA1ln
qqpNHAcNx1hvr8NENlcfBymKxHGBqbUlUFL31D/gf63ulcOIEJc8SiXaUlSgEXY4+qEZlC2sNTg8
5QB90R7eVUtU0naLhW7V9AlQDF8TXywrxY+NPZb2SBcBQ4U+/P6fVFUFKeLM/cunWpL66S0FHyFt
LimHn6dEAeO+mNu83Y2JPcIvpwsuDFI0i60Q6cM8xb0wn8PxOzGh0lB6VXcP6LRBvi0jM2uad3Yu
vxdqgY9JWbv14OKoztwJ9kGZWVqosOI2udaxECgSjyfNYjhWRGWFSvQSqAhc00Gq7B4qNXLOnCjV
zLLx5tgTiyCg+hg29Xabfh/4a2STJnola82B9CxqcOJyxwKgXCvPslgmYugaXQqvAe81N7UrjG+F
6WJCUGfLmmHDDjVYFgy1pPu/xdtxReh9/Qm0b62Ugw0v/oHOsaFHzzx5cSxq1gpgdg2e877PylbT
aFrmbPlXpi8qYEvOS812gTHSKLRx1SIWSmPHlcPtI6PvXPc+QGnS9LNNSq5sqDmyQrzOZnABM81N
QVCY3zfQE5SVKvMCVo6zcu2dsdD1cygODhGUaZNjZphUfr3FU8bMdtGweM094EG/4wxxPOAm8GyJ
UcWkacqK5o7KoqwWAiLQtoNtTSF3Ofne7FGQ4kwcZPTwx2Yo4XvFWJ0CGnWfFa64pkaFy+0pSQgP
JwQDJ3hmBSJErt69dY3/1CM3HfaZzbMhMQrtkAUaEOIkXJTMddD9cibRQ35GPqJsVPHGGwAHp2W1
RHh2kv+Rh8xnqayAyRKEwWoDzeCC/gbai5teijf5+t/etqLgGsYv7VRLFNQhHo+wUgOzuEXL1LLA
NKZsSQtqlEcxSqEf4fGxxs4SGPlgwWmbSyn1z9CiX0k0woDdx3gyQOvW7R2orZeG3P3yB7dJZa3H
9DliWL+nAg/0v2JNSpq1te+8l3RnbWw16FybtDt7bx4C2xDe4qXuuodFecsxG7VdhdiU2hEzdBsC
xLw90T6oX2HwvMhlfr77W8Vq/ZGC9D8Cvtt7jmZYzdnssOB7M5Bcm7KBWwUvJa676nJovOgFYqWN
49BU4YsiUn5nXuG4PeW/OMihFeshpZAFE/FvZD6wMY3inbBbc3RN7PXDIyWpQZAQ8yzN8arzrs0j
hK4Wt0zYz8+Dzy7C2XZ+ZaQPqwEPRZEqH8uvrP7Ian4Ds6E26/38Id2H8WfBSBcY4MD3vG4drFc2
xV9cvdJavfjJT+kiQ0M3pzUSllQq0jjcOXNBNgGH33u4yxFoJdMgzisl1uj8jydYOviy2nBzCldo
SLf3HTtbWrREr53zkWmMF0yDqugCaVUIkoBVg4KFzenstYBxC580liQ66IABYX8oaeeOGG9wNlWE
+ogsfr1nCm01CX0m+yO6jKXCD6x3ILDxClZQhbhtoEk6NhqdMoYCZiSTC4CC+h9s7oZIGyCnLh+5
ywODkXb7ou9nnrsRc4Zx5qiVVUjTOwnOdkGdfushzhTZP+t/WOVbl1mgKjf+SOaQxtGgBOcQ9y7I
4j00bJ1nX5YgYF9wz0b84HpbHEQibRnOkdb7cgt1HAQZkdgaj7s+nGs29aZBefOml3xAFV+w4igZ
rrghX4a7G9MUXIdH1I4MbgXAa9LIytk2d5D1c/zjoLuEO5ZYsVl1zR1oghZmWS97ToRwSN9tGiTm
Q87Fa5mxHUu5xOTrhtjYtPVtVy89rfBnSEHlSnqWilY7u+dqTdXvna0gKmiW0wBDnc76v1Q8vI/6
0xQdugwCWVW8GRQwLo+85sW2Dj+yv9MTck1ZuyPpI88mu3cHTcFiOJRWxzAHy+mmsNgJE8luSxbA
eqGeCkEJq56rK+VO7ne1zck3/FbniXKgaDbCSnKyloRXHeWSA6Rw6ZUfkpDgBAtfYjc67uVCdIvS
urzX7G4TWDu5zNg7aIgl2hzgK/PrrLoGN4SklKOyB+ZaZQH8g1xh3zq600id606KlChvaxNp6g7D
oGQAo5KnBYNJYZ28/7LJQ/MjEYFxXGZHnQSf/9Ews+VzFtrq/9ytD0KuwXt8AxyNhFNf37gm6LwZ
OxvWw0knupCexH9E1n1ANbs3RsBYVIGIelmjtUAL3bakvZPO5RA1X5nEC+/QVb/2aI3cVvUhudAc
VMUORpgvhw8x6XXZTJRF3fMHWe55ELNGo20sikCUO1viZgBb+20qMO7CAkWeGUG6aZyEUFLM0lpp
TQ4oHKV/tu41Ad8nkIJB4mp8If0l9D4ZxRo7PDNdmOJaCBbHgtVDdq6WfObqVN8Z9rg+3+F9Hkyh
qrk+um+s3G9d4xwAzyZbbUxu/yqmLCWKmWLaOlgnvYwf7WNziyjoDx9aLlM17zEJ4RyRZO1ynKCV
Gxrqdszum+xu7f1A9hfPIcYX9P52QDK5AWjKzjl4utEYmdd5yrmzy3iIzjxOZhbIp+bfhxkSTcC9
AaSDB69m+4Twd1ELCVA+RBCuvD4u/P1/GmFcMe2rfyaxCXCbwqwCTFkM+UbA1GSEEujBlug9Ad3U
05Pz3Xs3VTq7Xz/OxV4sK8Z6ZCEOuZWKKU+F8O6quEPRiB6Ttn6YAuYKjwh4rWrq6UIXkaM66/xW
nBdOyAEe+qZCLPgYmCfHu+wWuHamIyIHwSCbHnBnMt9Ygx+PPoxyy+MdTXrAdlxY5gWmyiA2ZrXv
Iu0GLtqw4HPtbTEXiWDY5rspekVrR0ZqTTOb4cyC5E0WEHOITSTGPCtW4FxwZA8xDEHpn7icXwVQ
tP6cMIbj7IdV2L3DRds1fd41RUgjFYiUc+7kcr+IaTlqK0F+dZgmF593XIV1UPFr+gF7R/g5PatU
o/0rYkvIX3M49btAEKcLRrjouHA5lSClRsrkiUA4Lfx22apbonsiFP7xb0b2u+FP34rZAi42zXzF
6+HLHsR3CwbFtRpi3FhQM8fvxZR39hh4s9/XgFTUa3mqMUOP0AW5HJ1Ur7N2obHvGC3aADkrYZNL
A5gCAw7oeMekN0HQX0tyQ7mr2rY10Nlug8RcZECuoEYZaPCCcYRXADsC7+NQE7oqU6Lbdz5y8Bpy
X6vCt40SKMeZmYJgP1hT/PsShpOVs6gyYMiZpTJR1ruysVraVgfwFsMQEQF4g58xc6vlcCapaMLt
tzII9gPCt9q7yBTuLjvRZ5fk19/IjEgq8mBonk5Z7fFQNCJ3WW3I9CUQJCx4NULKTNykfeoyLUHg
PFoWDuGcSMrE1uncV0bhoMQvEEDxxSU+oivAMD0rLwkmYw6KZHAiC5pz9EDfetOTwsUS9MCwy77U
x3WSRQ1KCntXWPgcD3gRpDfPiB/boZ1f7d5BX+jLFpcwdsKt6eI7vZofPCBVVX09mSkKHNCweIOq
YBMRXaXg/AqGGnjtsZsMX3G53rk8i+1h1lXyDGj7Aw+/eAcNsfoWaC0nKeuVZFUCFTqW+lxhmTSb
aZRsG9iZ1sW3Ld6Bre7lm85tNQJPcDU8zAk+O/FxzvCvzvuZcPkmdy7uwH0FloYcZPyvvi5+Q49U
oGpzu2lsuReJFsTSn/AAUkmXZGjmBtMabC1rKNRo+3eOB4Lnaahhtk/OaDRGD/nBBdbYT+lYxOJs
7NO7JcD2JXY3XR2Fv1GuBEBUYkwjL9/q/7I794JAPahKm4dTV8DwSoRVHXmrggbLuAUkXRHy82Nu
iaLd+JuE4HxRkEMqxA/PG9uIfViJW6amPms6uXeUUBXosf1L+l7Q9SQMk7zQdFiq+R1ujYl8TokC
qhURk/xCC6hc04Hd+WeMrLLPwRrxvzOvGLJndYv4+yE6uW4xPRohF3w9M4uwv4arCstG3MgABTIC
YKuGx5fptLROi5vyTnCNsQ68VbebGZ6gtjfj/xlHDZAiir+Uba8k32MWjRepPykS2n4syIki9h6O
6MQbxiE1YwoRtjc0H95WH+KRNuQpE3r5+B9Af5AdD3EP5YFzrSg7KdD/JX4GqsGLntgqeZ9x9DGm
y7HErOSAhSmfqsucYDD3XXVGoLtsgQAh7ipJNkd7DAQ2NISlHaOzX7+qbzZQhJFhx2vx7DtacbHk
FzpVDbbO7boPQNxlC7k3cVXoBdLjiGCqTHWm1cmJfKgycA5LS47l0SfVOSWDD7iveM8IwdA04kkp
CUsF1Fw1D0QraKGqcav4EHkodGBfv19rCDgIfVHdPRkASVJQCb9TQKMVtx1Q2AyfOOWNTdApbz87
QeBdnUl6LF1vYdYysTd3FpObyL8PIy0zayBxLPZXo0m7RpX6oVhEuqWUMKJeNYRK1UaQEB6aySp/
KSXd46e++ZVU751jKPwkgSdZkG8pxQ+c6ZPNLNxUz3YvPylXYzqSv3v24kHMMYy6Cyk3b6W4mlD1
elpDpPVnvxQMW++F3k7ZuEJ8g/905VKgAuFzUqXQzArv3FC+cC6Qv4rlQL3KFIchRTszOyUSCwRm
T2nxIVphjn6vZVVd40epribezNMd7ICykgCI5UNm7qTgQHJ42Qhkn6tHVATf2TVnYfOx4too1GqE
RQQySCvdVJl93FhwmzSE3j4GHvHKGiKT6tnbPGYglMFY3+KfXlmp7D6V3Js6f5BdGtH6C+WMvCIy
wj7DsRG3iN8Lx/augkhX7nNoZpTq8g7Mhnoy9IOrSYpUPSxN9we+Cw2dn8srUOQjcGwChZRbN0He
0LbsNPO3WyXVU8dWsN80qY1Vk+zI0H8TyhmO+RXlEVONgEjwOmiAoz5o2jZooY2UHStBs6Groy0U
tZwX0JWbvQ1NbX5dtDFF6T0/7SW1LEyBLkVtNG1zweYyYO7/t+Q8K+hV0BOK8y3pwjF9Dom5HOcE
hI0Kq89ZbZHIVWOEDauEgFRu51U6yByCkwLetmXnTzjbRwXa38OszfiVU68A3eCZKdbL828nHZWg
GNYURF1lmiOQvPTdJ1XzC+hTIEe7s8+uTJrn678vaZCxlcC+LhfAVCcNvuQSIvK8Q8YmX3fN4MOR
97qkcKKFlKrMQhmZfSz1WL+n4roH2VF/jewasXSxLOM2+H3MIqbzQ+56FU+ZcsUjtOGMRSjR2VmD
Y+Dv9vW7zxDPRGg6KpTGFrkOQFjiuHsG49hgn5YF9TmGpYaCjDkutAoh3YIG7Rm0ETAYIJWtW99Q
RyyE7Cd+tWM3qUNMvNIW3jXmhsDftI4+ozgsbds51nbnSg1DbshKAXuCV3ecyEJycalWhVxCpV6Z
RJd5uGeIbZoSyuWZi4m5TknYwz0Lwk2rbiTCTfAyBTTefV5P+2myzq1vqpcOqD+OIIc+uIaA3r5J
VJCw8XltyYPJHxZSyLsqIR+drt6OEcRlqwFtJBtsIq/X40dRs6gmOShSAnUaFlErd2bNUdAzz3zt
NZ5v1ZotNDCGJAofvGFzLiOTrgR3fCdFnOeB6cwDov2IWP9GuVfw8e2PogXggOtHHSAUJP5u47Pw
JuNe+4l75ttRw0Y9kpxNxpYm5jsIf58BJl8gDy650Qy6IB9n2AO0C1iMZ630HIcXKShVIkePis4I
sVBdee+oyea2iYU6v4rzGZGFIa/y+scv/EdQ1dXJc6T+vWCvKMXs0zR8e/TWylw163FbMf8bX4lm
4YN5YUugCaygnp3b0f2mihWi9donzqa5hYgDiW3qwm6r2pRrDHEWVTk+sFRpQFxVWHRShOr/zako
jPoBUuNmFX3h13bzS/a33lnzc0xQCtnB9iyFoLly5fpXMmIE7lo7v4gc9i7DDqngWpNMAIKGoLfE
5Uvo7/bXKs0yrESnDyW764T9ERxoM9m7CtAqMs8JdnlXQ/xHnXemgSBscpkKYbYNE8/CbqTM854m
6eLNxrHVt2lX+H7pKPGGUSF57Q73qzWKEAyazkOBerE7zvfTHhiX/o+vQiWRA3+CinDpcbgt4LlO
q8CzwqbtetZCBfGBZJSTPCmz1akaYWyPVll1uxDhhWsbYEmstzptzU0xaZczD99agVmzTr1LFY8q
wpIyZj+DU7D/j8IHGkScy0lBFNOWRLjbdEX+bEmw37QJraY7GwCRLfWBA5vX0km8/tio9+W4sGEk
wdIMDmQtcW5KcCnlGoZuabdIKZCar1z1dff1BtOOMWNrPbu5VBU1EoiuA/bCnTNU9dC+rJPPl4Fr
P5QmjqwEYtyGoKCWGelYf29X6XoQxmkDrkeGyyUlZ71F+SQQnDNPdy3ekB2bpAvL8nsR7ThCOdha
XH41T1sXOTDgrUV0kBzogk3ZogewdH/Vlgp5+FK/EwaklJTP7WhT4gD5K3z+MZKsskPn/mt1yaaB
YqAwWr5Abfk011quK4+cK2x7eERNRMOVmqGhV+WosMkHhqHkCFrZWfIynZka+SAO1b3cpnF5wqGw
Ec2RIJSlN0Gd2M3mG4jDPjD2NJn3oB08m2AkKZZ6qbor6SyTo5O1zcJRIncfcI67lF2Cv+6NHbkL
mYsG0yepKyByB6sTIv2C6qzs7/79Kr5Egl3zrSpFVpzkFXnKN7lO0mUr7IuHiNhsf6k4fIjmDOAo
fgAqy3XeRIAzW4bANhIRG2C+EczZ+RV9/bo+l4UbbBDVsYVRTGDSvds4S4cu1+wleelDeTt0Bo1f
0SpnS2jyAD73nI6sHrDJ6/OqeX0msh1gJYnlxshZx1qvsVh6RsqTm+9YXfylnxTDTaM2vr4Mubkl
pSlB6FD8fy7kns5tPUrT5dj0SNStGHuQGAPZN5YgBy6f/G2bRbYMPwYdaMRWGOLdNaCb5obWRbpz
BbePThxL/j7kyC64hUhvics3B1wftVUnZMniod+eMnW+JuQ6po8GWJI+UZmS7tfYYhZfQCtAZ1C3
/G2GdWmmwBdJPFQjJrp+VSwfOzH12iPjSAQS8F5sULpuq4qFzfKPLITJjJV4sKciANBT6A0dWBPH
dMwz8m05rvR7aISsK2HcP/OxfWrj0LBSsaEekfOCDwLfeoOJtUobdQPGWp0QRKfhw8ZmRoE0oa4U
20w+NEyCOTU2Yd2+HdPekl5nDKwthCOSWjWQAZHikJ0O93AlUxQ48oh0x4cUMCDe1imalCpk0IbN
jZOUt/C+4GrhOpdQIGCQMR3gy+8nHHkrOisd/vaGYMNZ1yRNkKWsHkUNf5K5M0/Ts9Br/hogFXwn
oemYe9YgAT0Nb0tesDRUG+8L52QFpgCzqRKk7VeO5DzAsDuwoK4s2jpxvShh0D9TEer4qIvxLWtU
AHFvF8C+YRBIByYtEGz0NB7nTGryfQyQ3hlTLfAoESOWnX0R7f1W6sca3ZsTcvYcyLPOgL2ivcLy
p0cv6QzC+gvLM0Lc4vVXUqh0R/l+sDoHvN9hzzkrU8d/ZGXvGwuF2hN6/lfEaVvgX8KB9+qSH+Lr
ezFoErJ2cz70pBs46NqL9QZslBGxzGofntJSiDOjlrQ5R/cOBwFeBtX/C5yM6KWMplBYQEO/2NtM
A/7uegrHe+8WC9dgHY6kmB+1ATNnPeRFuBeb2suKrRhcM3/Y7+ZAyR+r8oIsXnsBDZSyWaJeC+qt
unCdE8pVO2gZRee+HQ48vJdaHlkL7DuNdWHESwL1brVU/QX+/7CVEE02tJQSoAUVqiy4xDL63eCl
OkYrMAouh8v5QK6TxjzOWmmXbnIBteLUq0eXPG5VKr+kfkkCtayJYSkVrdtBqSU97eOHw6v8agBr
Y8OKH+RG+bJoVUcLT3YimkID5o3VfUzkcUahzKc7Lq2KkFdyPD4HlCtKrgEE1tU8JN4SLhtRqD/m
59/TbaXr44W/qc0UT0FjECMQReWH1PNvacb+BAktz4YE+SavstEe9XLh24/T0mDLaajedbJvuGVO
MgvK+VBzmlQ2xuy2y6vhaQCfLCXIgdpEWgq5G9QyNTL57+X3KkCJ+aPJ4aMDgswZeDt8zBDmCaM3
l6m6vAXBD79Mj/hVPEMIy/pT0t+87Q8MTLl321ph0MeYe0X9m7rfce+5izBHfzO6K7wKd3wHTjdE
4gDNCYcNU3i+WcDAvQ0p2wjxKXyzdH4pSTs2570YAVrVDBjkXz7L/hdokhpyWCC2qd3WuVKHs2jK
/lZk3s42/OBtYYa0rZe8x9xnS7PZYIsfSZJkabojYYY+VgUb+j12wE/TYfuM825OOpclL14Or7V0
SNs39/orLf95F1cQ6htySQO4L+pqUfRlYzzvPekjHyoFm+owZp7saKJms1aIjENuLOokHffFOcp/
TNkUu/aCK5ivrqFySyFGidHMZaBB5NKi6qP/dxwMz8Xtjasf3TYQ+VVaSynR7prQd6gmmEZxIS1U
+1ZgrmM56ysCfsttxMMaBfjfCYS2sVBc4fFHUPtHSr2YIlMydz2rmkp7QezoQqHSbaOGj72Ga1pT
cJ0+dstLFXbI6ze8w9y2KFIGNIDlSqpZm9mjJVbMVqfP7jdZiNVKxkC+yNAQZEVWhqrlHDVGdA49
wXMiyJm4rQjeWK2uQuNXJSmOupR6jHMNNf5hNs+OsmIRXDPRci6SA5BbevHc+uRTt5AEefQWIVv9
qoo34GGNUl5IKaesxuU8S0no5xarw9j+6f32oKUynOre1puviY5qhu2//YP26Jl/dKgABaaj7K/H
LZTmqOB61SLX8sx1y0NaoBKZxA6SeMSfr/o4b0NY2cCPzJlhzne7hGkp+0Brh4BlZQJW8Ep3Zz91
etXoX1rOXKUPHJNAAy68bMhCxa7zW4Yyu2Bb/AsHyly4EIOPPIfrmrz0//6UxzpBMQipYKWNqNQD
4B75My8ffQNTXc/5AX25UPInSQm1TZDRlgxTQcH1LA3/7+z5Gi50TGd9BMsbFa7SLeVHtPogxSth
ve9bv+f/hX5vvVF5Y1MZs5OIfKesS7CVKtKVsNZqV4NzA7jx1usNFpz8p1P/tBJcytsmht1VFgd2
Q3GD5Z13R3qYgLxpP0ZwoaTkA2G1knMOMA2jp9zDsdOvWhs8m1qGa+oE+2jKaNhqpPbXC2J9N7Hb
rROEfWvnOWuvD6RC+OJoUP3Rl9iDyhAhBvl8Wwn8/wv7gEG0wx7/OR6REK80LtFYGdteixnwGWri
JywOMMHcw4sjX0cEkL44PXpd6swEBmfDfgxtBNGH7uY0Od2F1J72SBTJDW4E9PDCpvhhNakBhlt/
J+J2Bq8dELhVW3w+ohEKV0/rYNJWhUgL4VSSXS+O+DRHOr8IrZGQkVqyYMGW/Ig2eU9INy3lIhcL
lfr8as9fKj8y29wJ5UgR/orXmN+9eOCxilQhUS0NvVEfqVetXJkQigBYG0jqL8aZRU2qnXicsMlO
9SPzBI8nsHXO16cyzR1M+W1LxZujGqcRUdMkNzJ8oz2UnrkL58jLzDqaAxg3
`pragma protect end_protected
