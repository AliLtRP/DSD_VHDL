// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:20 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oT2HYF3tx7969uBCjJ9WE5YgNWrPsJkgrvR/g1auG9rmPbdADy2GhFgjcik5iLOS
fwAB9u4xmg4DirIJynm5QN0gXwa3CPs/xcbDmva46b88GI1McsYdXvVCZp/KBe7O
AZE9SMvsniRWmdya9eSWk1P1e/qsn1PvBcHUuXrPCKg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 71568)
rX2xxy/4b9i7D8in69KpIh/VHmAfy9UgKHl1QjDzcV1XMYJ1tgDPGz7QhrYIZO3R
3qNNTN7aJqRGiOY0itUmlIR1qauludoGMqF9H5nfS1c4TflHjGVvkDEqIDqbKtA4
0scAEhlqAYvOiw7RNkIiYN6eLwyqSTUdv9RlK2mU27hvwNsIkpwTRdkZ2QPmc0ds
769pLebgyCY5Culd7BactjsiugsOevI9tJPgccvlXFTzfE/4Av0mWHOS75kPur6e
kwreWLenJ1AFtE9xK8RMSpiRWCReICeq+cP6mb+UD1v5Yg0qqCni0htQDaoViMbk
jDoVNJ6WaeYhklS8w5N2mrYOV2cw8u/9HLGo0MD/A8zH5v8IxxqyNsqN0L0fnwEk
W7uoXS9fulX5GBxnXteedhnLEURJLXw12v1UIOcAQOoPrVTIGXivjtPhvMg0Cou8
YeLpHaslgBbLZS+6NdtFvA+WCTWreTwUJjnAykPcpiCCBNJBuxKkVbGpuVMaz+ll
Xp6v6uO8404oVPfUytQMtS+V6lk5CgzW3sncH/Kc/d/WcVoXXban3UDXvXkNPO2/
Z9x+Kzhc+/JHTlgGnK3r4XxDKbv4UgdB3DGmmBh4ZMSwldtfvE9qPR4d6Kn32CHE
kI9kwQTS45olssv6pXrZ3Z9nY1pt9+t3dTvQV2wVrWXqjCxly78GysTwFAmrsfjY
0u9WSwySgg6XZDlb4gDOVs1LWYyC3SsY7Llo3fA4iGAUzXz7/M+8cPJqGahsVY5H
U2SdUhDE78NG71qz79ZeMq+sJ9RRxJ3X+7ESE/PKED3j5MxRZtXtbCPwtbCacxy6
nrT4MoFCiPantv1fi5mV8UDEeR5xfa432nFUJj1PuPeBcJ4+EbsmCNXzD6KL+w5/
7G2u8wXFACnsa4EXH/hihsvvXEzEnrtyJ7+V6PJRQ+MDltTTO3IXvmGOjF4AE6RS
ZEwD0dja2UBeUvZOFiubZJbAIkn84dY0ZqasSbJ5JBEhcdeotn+h5dP6iathZ2LI
FO0Yuq5a78HCvhcCpgBh7rWyE2fZdNBn+N1EqsWqn5uAClCTPMHUwT8iYeTPTdJG
PgX5QZekV5sPp0iLkqugkiMi5KP9ZZurQaMNzbApDMBJ1gTJS2s/Bdytj2U7WKQ2
cJFHEMYMBzvK0wmAkhTvtsBKVeIpGhaqSNR8jvXjFgU0RcD1WmVnItyoKJLpRRBO
hjCaofJOasoBIIto2PLC7mUcSocUgN8maiLX+IMn8ZqR9XxltaLRdo8bM8iVXE2k
cBUPhy2oOK9JW6HliKulIm8ujywziEvhcCb0wzD/HOMXMmlfyXooPZznSiDDbE4X
G2MXkouXnIw8vDC7EYc8kR76W4BoWyzWnlKZGkWEIh9ztXkuEr68/yznHeSV/glW
LB5wIdv2b+dIu4unhgh4ryzEr9SgPO5jXd79suB/uyVxl1y8jGUOs9TKWlxoH6rG
lLUY0s8VjXKlksRBoYab1brqKBWOhBJA+zXoC0xR1hejVXXnL3j1GkpeccHTEZMU
iLN0y/do9YJoi1v+ACbaH82p/hwhEpfSKcq+uf34n18Pd7UYKevs/zwXrW1wbvOK
LjMphM6oFvUUjQlAHFpt0x+eiAbIklptl7qqtxu1RK38laMyNOnan0LSBsrMNKtj
CpbOzutpU50XQltNP+uVXFoEW68+tu7QAbjE6gryP9/YD7TFyFXp++8pmVh8vKRM
XqIkP+LyIyMekQHA6wqdav2UKVTn5/wWOPNRy9EWFTaPgkJx+zu65BWSrlMg1YPE
UkVzpbi7nxq5tt7CLenY9uSsG1pCY47UkHz8T5V6mLhIszsFAmNZNpQ7FhQK22F+
Ef47Hfxw0mYhMKFkDS8W9PXPe6dVpHwh68chGkeEWEOOZhBSU2fy7k/mQMtTyIU+
Wui2JmzdvMgFPWjWa5qms4/14qGKyZI2NoPtcGr7c8fvM+ae6FgWUIkRoMceNf7d
SnQ2bNLCFUhGw0wFaFk4fBkOz09cwtMZmoSCOQVSGXoaC2gCyk7tXKjfI0n0/DkA
mFxptAtcbOJfqjXdtBEA/o3CRr1Z3jSWv5SRdVmz+ybrMnVQKliaQc3CzALYrFAb
+0ZP49znk5i0nIJZ/DlBioTTNL6HHDWjkK5stsNUCobd3HjxPIE+93UcqCIEChMG
lzE8H+fcQwAOi+Q1571Hz65eZFO4847jvY57L8K4IGBnzzqHP7X3uW8HV12c6PHn
ME5WglSuI4qAm/70kFGJ67gM8TjbPa7j5JkYdz2uGskeQpXj34bU2FXhpPkdDtIy
fgj8YjB4UuPxRIQj8I+OGmdPd4qLhioGrrUMRrZwb0PvFGdr0jNnhtTpY37xlKz2
p2WyYrV6iSqHuXyS/q/Ne9VRudkRjV9jw7tHu4GDKVmOXLnX2aFQQW+ELB1l+LDa
vpL0pOJopI6NxHiZ1Cv+dy1avIZjGs3KEm4tzZgFtmK5sp6nsI8IlkGu5G3kmKZ6
RQoooaOzRYirfdi8ueC8oxlXIlPxzyfDLiPLh4Kn+XM9NI591EnIn2pdgqSKRPky
qLhdv8t9IWn5iu/QqszQGujBNdBsMH5MugYKrLBV0X6suGpFkIPUiJkQdQMB4i0J
mit5dK99onI03unyy12tTgO0asmcmjLIJGP3cbJMDdqqBelFsMiCRGmxknHn/q9Y
bjZCdpPXXVvYJL0szVaF/7a2G+rVk8CilEO5kxUTRtLdr4dAlF/oOVBE99fBh4LG
yXQxfv2Yc/4il5TVtNVBbUgMnzgjOat+3FecboxxoreseUeZD5P/S7J3kT2rj8nF
UTSdRAwoABClVBhITtRlGBWIQuuZ0R1XqUJFSyD+qJQpgrxdW/y/aTBXQgFTrUR/
R+krx+2f1yBQkTxGwUkg0xAIF8WqpvQPycwEh+hDO7bmB7YLDnN9aOq+bVxUs0bN
Zb1WBF7UFYQ9G5IbFbgcLEpPVRp2fGFL6ROcG2qsaLf8oYJPGybbp/dvBoz+DJAa
tN9cZOOF5s3afYjNr/1YGe5uv9EUWLQC9ElAkiAVAKj4sFj2xKQhBn4GeX0aS0di
fFMwj7Jue46h6v5S6queUz/6/QrsthmnmbaduNN068cDAzflEOiEcm6W1bVgaE1t
iEAxduFP2eQseCMDkOPXC2thoQkA3D0RvwcfJdTqWm2U9d5N1sacLwZnQPVeDIPm
wwZFTPGaQY3PmPd5ZXwZkp6l5q3cMwZpae5Tk5gwpXasWzZITRIExDfOlvFdUZUd
QzY4lgDuWgb7gqsDk4BUfVEeVz9VISeQGFcntJYO7ZkQyUaCt3ds9OcGLr1nsTB2
rfIV12wthqy9ecDLPoOtzI+uyHc1VofeEHSOlN4kwxYRlb/cZWY3FXenOyVxuP5z
LSUlfvik6pJSRQQUrTDTg3/rnALqyCr8utxGpeD6CYp32ZiDSRceFPxn26dgmZDc
l3ON0v5jWMQEMaSFtsCHj0xRNp3n8FdoPWyOBIq/24SvL1QVtgFrZfefqcQe08d0
yQ4ZVDjWJ1SqAZIDb0qCxyHlgDE+2FBy10QILcGNrmbjQM4wx9JpvnQf0uji/fUy
h/Ir/v9TU3kRtZNAOzdz8+IwNtFmnTe9FKuKDm3+O1augUedtiUDsgwTGoo8PpES
mqbtgnieQJWG6r10n2k2dHfxPYV/O55xPQHl4u8Sh0mAXVu4FUmPqAQlGsBh4WMY
2zxaPRS2NcljLRqsZBL6aIkzrlZJ2dh37QZa2HUIGiKc7loZgxe2FqeGphfHYwuv
hDVcMJ+PBsfqbjDAEb8no2rPtAv0BWeblDAMArl1K1VScIfceEyPKPpFPUzhYjfF
xrScrboP3UYqC1jPn39NbSzwzioTrQpKPuUBvQ8/ioD8GhMtlyPaRsO3vQBDTglQ
vJ6Lj3rJYDh98+d1EwUhbDaKIi8Ex5vfFPExV3WWvKTboOvCx6yQjSaGxH4FSpg6
kWmSQ9h8NXn1u3CsqxYou0Oy0j6uNEKoFf4r+DgaFDUXw2OH8wvqm26+6v1CnZOE
IXhAwHL29iotZ+YUTjq2TQ3EFL+T8r46TWgOdI4LkwzA9QGXKbEmPQOSUuAqdmMc
XfwPRb1Ovr3aOwU6pKv1UJg5omi45KQqBkSEGyCsEgX1te9872F+4NYILzP77h5g
LED5Z+yLx0vPOHepBOngPTOnAMrXhSfChqg06chyR0MBe7vktO4IK+Qxmu4i7Ecg
qOdfy5FfuqFwjBrQGA9IYFTuLz3U+uKDwqsEbZeQdZOuoBZZOegO+f8axjXHYfk/
+/f/S55HDAjsF7GjHktCAT3+eeUfmiNLliG7pgMJmwX2ylDXOTT+TIgRzvBIywOl
oRfzAH7no7JQP5DFtuTw/5EQ7C0tKRu8xWC7TZ1u672jPfaUsT6oHoQtdzbvoUQT
EacXg9Y74G5YR4bz5x1ROWwa17nDcQxy3MRhdmQLlUr4d4yit3kRcagkmNnEV1ai
1blyBA0WtK3a+vQX/dZGYqM6l9JGNqQKY1He13hydRofrEDhBdHUxtcVjnJkTaE5
8oEMMgTTo2ywOrbdFx4D17vTg6nhgBp8PmVYL3eoeDOPaUDH1HGxL7iVbCW08g4R
czcLErXFwjTaEAtG2zGW/iu9nXwQFUsApOHPmn1Nj5V8ZLr7Nf0XMi8yiBYcrYoT
/TdqcRleVKeqOGqxoA/CTuCUr8vqJ+oebKZ1DZJpXWdQbrCUtK636l0NUaRHq9+6
WPFTTQL+T/SgAc40/eJ7aW+NB+L8+hknZEAx65G7rC/nbSPAad7JLWhcH1mlMtTP
A0iIhqOqoAFnQterC38MF+/f5aSuDS4SbouiVZiTOIVrmwLmXDnm/9HZP4jjtDXV
QaBesK/AjlmlqnrbBgXEqOHLIGYB/nYWFUbPp3u7teUl7ez4ZThgYKVJ9XSQqQ2q
1244tJkG3JX3gn80GlFSRYB61LrIZmKAE4o1uB7AGJ3OX3lp+2QoKXv0ZYDInwn7
vSgjtK43jKPmHt3286kzabgDOIqsrS1u5SnfezSXEenB+lUlBypCYpxhhSZ1sEjE
oKNRnDjfwkIZrY0hNvjKf9hkt/wYVdGuT4gNpBM9nCD4bJ1xrZdCIItg5BbUinHN
tO9eWq6nqdeg5h1nG5ioBdH7idpJ6VfgWNqLVvdd/Ttk4MkUdXNc35rio2PGcbaZ
ouQXcOKtFR0Jol0mdlyRxEmcWet9Dg94ru9iM1pCq9t2YvhWawkb1GpDW1HsoiAi
pj0H9o3pK1K5SCmkPrs9DgxecsqQmhOFTnBewnUdOkeTtQd6Mqpe9eA9alADcMLw
wK8VYA4+UFDrD93rnF4EkDY1+X9bW9QhG79J0jlWkLgkaruM3FoI+KyLoMdFUfXV
405Y83+MuJbeoDly4pw9DBhSiVCtNKSgqWTwQyjxOFREFVU+AUPjkZWvLq/eIDTl
1C1wqMj//o93fV689o8pUcGeXEGPtcJ4283+gKvpvArTwW4QEHyfX2QVxABkb7by
RLMyXLWpI4BnzbneqnGxC68C1Xpcbc9NpVaJwwMP29X5IBTE5+dajhT8Pz6wk9vQ
zURfjweMuBR05DYSGGdoNv0DM+0pb81zUqVFoZxLtyqcpOrHGVwTu8aZiw2ri8Je
pypmajbAnjhqAX+W/yRiPsPHjQGjxqPdoTZU50pqoaMkpRJb4BrRCZqjSUrYsXeL
AB46qFnXh+Ee5MowhqO/jXYQuNOl7KOiPc9PFBJzsWRuIvP+/Tl4J9Gk/eX4WCEi
cX9C736AbTLUwmQGhWex60LssqpoOCuXBtL3N3XVXoukVNqBauUZkGSezal934wj
sPHc4wuP+jCAPgCv0rIH7x/NIoyTQ8JjQopMawkKFFRuMfT929RXocOxb4EuGp4c
X1qWbtuOUo6ebb67ZC6gT2ROjXyrONcPiHD1VAR/FZespn2Uqb4s8sd37fCCnC0h
VfmmUugVAW12kiOwjC9JD4apfWeUYXa2s6KLZgQyyKN7zLUF7owTDMd1E/8LRdZ0
edIF7FVeA2bkdKwd7am8Ayv3QfPxQ5F+/my4q6ogCY5gYmYyNwfVp5O6Iq30FJLs
oiJ3W8ju+mQ9tS/14Lpc3C8z7GGmQEgWwM4rwEI1nIfuBX3aiuEwq/WtqbLRmjm4
C1wpQ3UNDP/hnyFs/wTSpdsji7NZIIwY6V/Ul1uN787/8VJxb+jiqUki9pntkodg
dfxKyBXry8jZ1ef8uIosGg/sw9FFVh+Ig72oGGBe9QWLWU6IDn4q9mps+Wf9n4uL
gEDschvecznHJMbMx6SN/vM3i98+X8gKodwVwny+wNKU7/DPRiMggmv8OTKyU8u6
TT+q7UBKufVIB8nC0xm2gyR5duKt71c9KQBPNn9GP26PDlviB7vm62WHTWTZQApR
o0mrY8Mp4FuC9r/4ZuQ6hDCz+4egHLxoXhTzyzLMkyuVZV3UARsuNyZbVco9E3Fy
c+X6Pgd4u3RG3e/3LZY5nQ3HUOc45k6kyBUSHYttlk/lj5G5hDet+7umJhyHtmbU
uy23tWK4nYOMxlBr4XR696pKdcj4sCMS97uUHlCEOZp5o/39TrIkB4NW9XPVoO49
LX9aNWkpS5LH5JSQYIZTZTcYn/HSVAJuqQ4NkZRjErlwGCqA1KfWDFNTPMiRfAxD
NFaYOZuMWfOt9lwvwhbDEzBPi55Geg4IN6H6h7ajRI+PFXV/7HUu2sEa0u36zo1M
U3e6aidOb/CryXK+/Oz0DcTYOr+DWd5IL3GcyK2l9wAnlyt3+/yyhTGzVCi2J/b6
G+vaSvWgVXPIU7NA8bk40CHq5V57SeaXVZnBuBKK2twShYZNDgpTzNJZ8wFLRNo9
76me7ZApOF3ZBYpcVP+dcbPxNhJzCx2VnftlI4SISB2uInLNbhE7tj0G7364cZcn
m1oNI7p+/P2MMbMzaZUb/50/0EHxVYCchAOjQLdI1jqIxJVzKkzJAKLZtX4phkYG
8QaVlXVvXOMNrim8mK/cY9VGNDThmCJwbRf6A/l4AuOT4cGRQNAdQaVqMfAP3I+/
t7hsXruolThpQ+W2hi2sISOTT0Rwqbo2IXGZsKzvLYWYuVom/D9DzfYajo05nbnm
pGGo5IKh1g1yUcsLjZRo0AYfzBebdFpnTUpfX3n8FdIBZ4Simma7dg7KacvkCI8e
T/7AFmgb6p06O7c1PFrhQYpBERRe1QMRkoIlR9J8/OTKs8nwRSdJ3JJmYdT/dIqI
4yBbsJmMyyO40RN36sMlln+dpAhxrkRDjcXqfdrIe4v4IQdXClsvQQW/ezXgpTUy
TUgpDzgqsU9a9ge90a1OCNTinRd9Ut/ZiylpiihyLQoxWjPyDB7JQ4VyZxaG4/6g
29A0RTfIxAzb4KjNRvx/0Q9cV1+mwF1ZhGpUN+7Sw1UAVQvMrl1LGz68UJkePO8z
Ixe4y3l8H4y5/qFvNdcfnjO94U2xMFh4cyYpJWoBHTuO5Y37L4/0dWF8Htkz3OwZ
S6FAa21/6RHcistl9ZR7oIzHCiWUw2TBAIogyEXw9Qu8IYPsmagi3gF1nKIhhDTP
M/K/ydiV1YseKYc744zDrvTNZLsa8Fka4vijhaZf/paUOK/N77djA2zNmamcxPdr
M576SIfd+snFsYo0BXD656ZHBURu1ni7lVM/2WIM9aIYUR9fiK7bM+WkVAZ8FB0U
UG22Z4df3HNC9c0rd1YGKhp2FQpoR/hNhFU5aXIoVvoJfm5ga7aH/unhzD6k9oKL
0WH4prbfM1TV5TwUm4/HOVzLHKJpnm+nHo+R0eLHHYfNWMlUJz7kRkaG+8GmXzdb
VJ5zq8Wfw6ec3/if1vT7OTWTnnksmj6KaRQh5wl1OlQ50CpjntVLyiDvFcOMnx4u
S6yYbKKuMIpXbII5wZIOibnSJ8LspcIY7zph7dis4SbTvuiycqZkE1jOb/IjjtuY
7vCZWIxXvTKMgoZniX52kv/XScQxzwK4Qs1lugulI1d9nuDhzrHP2/s56IeoRQJI
tMGa1egwQu0h99d6anvlFWdz9O2Ahyn7Dx1S+wnH+KBuOvQuiYCO7n+VPZx/ks6c
K5h0XLd8Ev05umENTXy3QgNjgKkIHxOVXaz8nG9XFHlkleP4cXSMh85yc0fDFaEE
hTnLwgZH5JpNa8cxuYEYSoJyvr8XBHIgb8Qbk0TmJYJC5QdxJQbqiGsEpeVD7pV4
/Evb8apWP/sNq/v2ZKK2pnFgcDmpi6HCxh00WjidJ8tVR+RsfOkB5CAg+TM9T2oZ
k/feWD6u0LLoU4XWtnehfNoBNCPBlEncyEY4uOcvEnWuDkWUio7lPlmwFAetX2aI
UWMnYnhVUtayf852f5P5QG7x0FpkNtHNWuNDbdBYwtbk481yjpvIIQgbwyIgtRiq
Tcw1hmswcwqgM5Kmeu4+80x0DHJDVMEqVj57CKxkzSzTlfYJ/BaIOqn/k8QJHDPw
O+3Di2U4sCI34L3pEbqXjCNpfOwRlTO1nneOENZlaQtiR7rMlHzWKyZjJTqOCsvS
fG0QtUCGCyXH4ELwJeSoHzGQM4P9DZ+6RjQA6djy+hiZcWrpDTAPB07RnZ4JucQ1
OR4C5mwo76Zs3DpmZWr6dWiPA3ELhROB8fIh1CKhe4b6wIgojXmEpmc5hJix2bN/
V89PcDazTOzs7iJK2RZ9xedg68Gc0FjLOxK5S1YXkWpzK58VmDH7f+5V0RUG1mGc
RfTnO3ozw+DeS2dH2s+kYy4nltXsj4QeF9dnjwiacjQi6xW23Y7x4cU9tWxM31OU
BpsX04ash2z8kfL1TngO5cWXDzF4gXxFFtMkpbaa8CjPUFqR6vcR8qHmxDSkJssS
IDb8GOIthGjIgvnEXPl3wCz3ZiOwva5gywMmwu2o2phichBqmjocD/K27QoX+CUO
fKNz4jb/JmQPrhg4ClHyVwu5hhukhJfOh7/UmB05MkN15iNGfXWdNrTSiGrSSRo3
zFBlEXIm/PnwyT5Mr1A0rH6hwQwAN3xacI1jinEZf02y+Ah4POL8Z4OWeWvcv58b
TfBXnP7Fa/lHNveikUzAEmDA9gs8SQ5FKEtW9e2RbwIxfgQvoEI5KjQNz04NFXqR
9acNayxPiueSn9aEOVyujRLafnV3+Ret+UoQsZu+Qrx0PpSWCr+BAkyC9WcZ4XDT
UnunQlf0wl1ZOOeZtaMbnEIzMYK7QEzPF9q8h+8cnre+u116zV3UOQMQO0uODPkn
bBnRxrHB/wTgO12cFHM4ASBH4UpqoVP4LvezoFHDIJ9p7/76IidZgkAgVGia7e6g
7QxWXOE+hPZRo/WTSybMOPBCrb+8tSgtSus7wLJVb8H84WZsXvRYeeTRYgTzFQkH
f+cqNcQYNCzzy6DXovZgc8ie0HF2DlCxt6d7duEiC0RBxDiex+notEo2GpK+5Lvm
UpLjeH+9VKtWb8AQuC50ODOE3AaS12bgoz5tpL3Got1IKVOcZ/i/723S10PsUdxz
RJeObFFqglQLuSEoUG1L3E6r5ppUZ0RXOrzhcfo1QtLLXViVArQ6iwezWxaWAWSa
MldW6fULpfozxMwvEmft0RjpiRsE0H/UnkFdSWGCjY29RoWqmTA7Uww8y0Ki3MwP
n9yZ+TFlpxw/K4uVX9wV0JRgxCrotG0TCa9uJi2ybN/fjmOHFPpmPzR9IDUgpGlF
oMJ6/DfkVsrIDgERgix7xpqpiXmhRMQtZBhZLKsor9Fy0GYBqSvkxLEb0ek7BfwO
nFGjL9k6iNM8VS92Gjvh/ZBY/Hv/gktNNpMV1dbXe3Rm1bnxnmsXIOZNdN+mSpmy
GcNiPq92sSqckJVCfVesCrIcMNAXKl8vq9B3XJxjN3tETKCC0n/V231XDbnWnqm8
1Ree847NwZkgFlxYBTHFtl1tbBI7C2h7PTl6HrUs41QMZJAtionm1E4bMt6boSEl
mSN6LhzI+ObzY2gkDRovmQ9gCcfzXnWllaVOwP2biBOAzTcguDFnrI8dKoG6LtUG
Y6U3mCZxxRXxG2d9nv0F+8auKpg1089SIvKMEbuhq48p5SlFa/eKXsrU4/BTw0OF
rbkrz0EotloIHzNF8OaxYwKfSAjsiqEttPZSdZ8sg97c4GoxbvKMNcUfE+4ghKK7
jkb6Ne4XM/dv7idk/NEu+0ZLuVcg/+us4FhGwshDz8h1Fbys785hLle6nn4Zpudb
KzOlmgCaT+V2W/suBkJ1ce17nKlvKncts16rUjtB/uHM2q9gJE737AiekXWcdMhc
RlSGfCdHjFHh+gP2GL03R7zaesa62UeroaGXCrXi1IMpcqbmwvs9XzcOOAc47VEf
hsuZs4gKBjm91amwWtKKg++IA+Wyyp8gsYmrkR/3pFIXz9f5CK5v9K7QH89zK0Or
iEua/tqS8Hsn/rgvYRXHYUuVFz4Zbsho8VU+44AUn7iSXepGeDZG73eBhZOn8xb6
suj8GkX4nOZU851fXI7yhmb6ypXQGz6ICckhWpLh5NzjPquwA9YppvHp2rsg1TpX
Avqvn28LI8gfIiUyS7evxRuTeuPIHV+YlRmCpgcy0zEj//z0Yws/J0Fv3nJ0gg0h
KHaVAISehVEfKMEBIz1/oS8/E/l1Bi2FSXWXBOUZXzOVfEmDuESynymbH5A5S5JF
0/c7GiMdZgGQPOx6TAwbTplgt38Aj1aqOjwaB9ng7Uy4eh2dvErTxpTJxSAlrU8e
1F8GiU9LpPDcvABOojhGttZKiqDwyS2agFJxIrzZEJHNrTpa2HgHnjvQLY129Tpr
sYvnA8cNS/+y5N+NU1UT/CcCFtEann1S/76zZlJtlKa9RVgBIlU9TmCaF/LffYjp
lVzaTQfAmiMjjMZrmDRvzrIgJ8GgxyqEvtLpux23FEm/lDrJGNRzXoHXCKpPrPU6
m/lLjjz+IylTHwkyBZU3cE6QgYkllwJFEKLTM1FXs5csvypNZ9ETedcGsuMXU+D1
e0QRcgwvsKURPSH0IRvOViCPtTD/tefEb0nyuG7GQh4OWbidVZCmxwUbPWPautXz
BPnuwkoGEHLGymnN2koKWBN+XnitCwIC3zFAtuQARJbsRdaKY93MN66touTn33UK
sPK1TF+8ROtWx8c9rLMzrJghgoWWxZ+fjoPHVqs+4Sv7szTSBdykVpch+TfC+cPT
XEU+HEfuy3kQ8LVfSOI4CKg/TEqJ7IeNea+HY1COV9vgC3fAeNKFRxvaSUJ3kv2z
tYC0ssl9e3xGCFXEKFSRvIYvST/r5uAOlaZMShoeRcDuFYbhr1pEQ2ypinoHi/pk
+j8WkmqRE0tzPlwYS8jGZskxT1LVXxHPaLQl7F5z/B8MdiqGa5fz5na/OxzvTcpq
8BXn9R1SY0d2YdKiHbxphoceIGWiiTHMCo0GEnFmpsh4XbiStmXKfL/1sN8fCYkq
CzvkKE80uRc2CDhil32KcPWD3SVSzrDroTr3bTdWN8OipwYitAObmJOvHxkmLFQS
cYSW1wCHEPVN1YPnUC2M/yyau7vs4djaeGIamlCooQIm26J6fp9nl2mp3WuBZb3r
8FGQs1H5vGDsl7ThAaRMM1slCckgJcbSsFNNiWLdlmRWixzFERd9b8y0fGw8QWxV
rLkC/j/HWKs81hcT+eb19HZupbfdywfwt0QrWQdIA9tuDLSdlpnkJx3lTavAT4VN
WeQU9WBkXIDITJOWbmSZhmw99kQ4gHXCRtpxLUhuTWUXpKJqQk6DW5/3/1jXSeH1
mDmzFj1IfRvAszsyoA4didKjlKqtl0uuMdvF9h5IXr6tc5SFwkNEnmDd/jLmBtYt
jyxNG39w7nP5CBo82bel+p7X1giFHUnCBt3awcYZI+Ulb32ijMbXUTVqrRj+sxmJ
pv2/bWaq1FmLs9rFguarMRvga9UVIjXPl3GqKVEFLDcoH/qsPpINUOsNoy5TYjcO
wmzUXdYZnbxmP0Q9oYcj9Z/i7cBHKiTalryg+tqR7ur3fPaNNnksDRNTuc9bJVzB
DqQaSdNcw9mhz/gHa2Ittk+kUt53BmO1JuGPVXR5feI5VjooJ5SACL6lpvBlahvc
ItuCup9h97LTWdrCmPSkjsrarLis7e70BYmp7cq8hlImIlU+E68Mczj+hF91ndRt
2OsFph0Ld/oQ1qCk26CLKKMHl1iFgrlO3irLQGUOy55x6TzKuuPn4HFAAD7vd23z
kO0lPKeotlU3YChSswgqShr+OS07UptBOYbTe3tjngFdX9yPV0m6EoFB5CqcdwoP
pNy2YVVcWPRlOue+WGPOi+kI2rokPJtOv6V0WkYrfdURFGucIj/CTPH7YHBykhK0
ZAGc1GR1NzXApYB4gM7nr06ee+zArTSofmUs92zWKHj5vSyBwBBzMEmJTRBUzrii
ws7GwjcpW6JcP9yNoxYB7Qvv22EDay7FPQ1YcwT2FPAtxGlMFVeQicbrZ+U0JjMh
BPDSZ+nn3SprEx8uIgq8eexk1pf0RDoeSNJG7/pEvth4T8oF0F2dEoC8CveBOds7
YEijTk0fyEkJLWhjhCVwo6KWMJ56VgQs9aY2upaFzN/pbIT2VCyaA+uT/Cb4twxt
kTPzF546d71MFS10iYi675ZF9iB5JmIHkkR23Wa6sbWjdXzXxPL8zQqs6nXxxys2
5dSFXnmXX8duI5uJGAKtV/Qzu4J+zkdrMp5qhie2V4ZQC7rlARRmWSmVQRzJvH6N
7eIQLWqRA1v3uPnM9VguPR6trtqlJvx/i/TTnmG4SG9tkvPmBFUepubuqNAhHjNL
btTMXSzARtC+aeI9wvrL5mNcwLP2Ar0D3xooimluRm9h9YnO2u4p3gJ/0icpproI
7XlRo03FrWk81YNMeclqopy/Wai/m5R35/sP0+foXgSg6anqTJSn5Ic4F/lYbU3T
qcyfh2w3muihc8Gobbsrtdutzz4JuxdlLWCcyLMUT47vI38NcU6GOtFyiy/Dz0HV
dqqfsmwee7697oDLyK4xNnk+DX+45UCG47SeVtCY2z6ySMlmnA2a4xnfoWYyDMTB
wtN/kA7J5zJPteIUXcTodbCmFiwsK2rstmusUdYjJrxip6pevUKZ6jLqoqHRM/+l
6XPXL9Yi1cL0T8N6qZbyHmlDJ44KlFWXQxvIhYK34kIZIPpROLcwQwl/Cvq/qAQZ
fhBeKB05jt+EDqH0q24JDd0uK/oYYKj0pS02OSsB6+3+O0OmaJl+Z/TjA3fuWYxh
w0QChIE5rfjBP+lpIv53amY9St2nj22aWhSNLe3QdMbvy0p1qd3LL7/feij30NUQ
OBIRBzKbi2+m3HbZH+wHPx5W5iADK/ArlVT9AW9X/49u9jLVPwvOvXPkxehADvLu
ZXZs6BspM0D3KpwkIH9g4jZCRKYtbC1tkBaK8sJglwELPEtHdqwS1M2C9ikEGfVM
zTGH8JzKq31nHqoyFk97Ux1bIRvSpqQFwSPiEwoE51D2vCfHf/ZlVfLDJrLuMZ0n
+uIbdX+H5lY5ruRxNxja7n3+VWB94F4vHhPX+LOZQWrJneX1ZtfTWBkvKsL5GBO6
+rw6GytHuCdKbwHIELH/TgPQQJ1qSJEgJSBE3vlpJx8ZQ8r7Kp4wrWMMH8FN2ahi
2joloK28/wcS8b6qhZWoaPwBFrPracnoLmEY6Uf2XlFSDEXAywdx/Iux2ate7hXw
qzR7G3XfBFdO8GbDWJwOEcv5Z0WOr15snomt/Jc4ctQvAL2q3Fl9FUjP2pzPWQxZ
VGvKLC0XXYSzOFFvQ21ssOpiv1/jieXQHRRDkLv8cx9ixVBW5dIfj1OvFrHDvyjG
3IyfNMmDfnktHtAC81ttDsuVQ9rAUUViNOpc7WPVOpnMQoGnTft7MKQ9QUCmM8tA
mlhtxiFCs2i+rYoNMEpM3kUWDN61EU3C3zxVceDFczIqbjQ0JDMYziDPOs6R3sbm
jiZfgR8nZp4yD2KhXAGvereLIoYoV4nTWBA9gMpX0v2PNrz6/qQWc5jK8VSA2lhr
smBguPtKq/QMvpgzFpio/smftzL3WVHZK4vywXFBZfLFBz8+1+gbjdod4sWGTbCt
ET1TzRhYy8U6ZWkFnHFMy1hPx48HRR6OmdOWbBExQ4JgfxHgFc6se3u5SyDNjfF6
sM8InP1kLya4bBNav54+Oe2qOERawRi3lvv+JvvshfNT5EC0VY48vWV0Xh4ZJ0WO
9/KuRTHW5n2xAGNvF1TlhS2yN+IZhP+qgAtiqxhStlrVnxbFQn7O6T/NLo8tZntq
WIXVliuSsYrbgrlIs5Tc7IVm0oRn8G28HGkKK4RJYffPTh4M5Uawy+IT0lSISavR
0C4H7sQO6ylDwSHQ5dSmOOymtBO9ml9IAIYu3n6dZ0bElHAJK4p3wSZf7i1PtONI
VvtzCApI/BoKxypz/yZUoLBwJvoXfn2cGkHzj61hoSgOX7af9bUKGBJ7IUJRzieo
LZA39ieItOmca8DXE16Kt6URl0ozeRzVsBE5Yn9sPrRrPuK7oSfFgNQVChdJsmZt
yCzlXvcKtq8osqmgLWbhRdpwv5ehwfoaIyDwXT19k3L91/KPVaqwkPmG9U6ZdnWp
0HB8/FwTmwvMuaL0dqvHV46NGFdxuydbzYfYHuXKInO1a+3A/2kjdZDT1Q4zIHB2
KbfxGflJu7jcBrCpG/dfHDuUzY+7UXR4P76x/yL4JYURpz9aQtypt0aIs/bNz573
V84kgfku8eUwVJQ5rycu882SYWYM7Hnj4nOr5XXpZhXet4A3PKe46gLu448JQXW2
5E1swZpUoadCi+8J0NWx9blbNRxNLuYTVGVVLNImRp5pJIpWqSgbzczUMlaD54HN
iujMTAFJCDg0fzddNxDUL/Ncgj+o+wK/wr3RnKO8f2Xn42EHOc25RI7sjzsSwgoV
ZZy2Kl6qp2vVzlE8RPyaoLae5G2PqrnTWqmQKCVJy7C4015e3iW0wkDcijpwJiVt
DTKCGdzTFMw5UsknVmDthKzfQPjEMrDn1hneCehflrxTc1nBItKnouBaGFTBF3Ox
lcJP0VjiAKSHAJBjAUzAMy+HE9cdjB8BTw/T31wyyqLliZaS1q1uBBIL0koyC8mD
3v5CCkyz5tiFHHvZMFgAYcx0qxXFy1fLas9CZFKdA5tLzTvS3kO4chldGPJxAVMx
x7k6tmIqLZrRcIJ4PzAOIBvG8+sFVpckphHetF74vcvq3dfJQCihX1vQmpCfEnUv
deJJNNwnH+SRadh+mJbZWPSib9TfWKaMhqq5XUUR6xQVDfCcnvANPvOaiBFUqnfk
sO2L1Ti1jdXhuMyg6yzNU6plu0QSvUzOpuRHSNh2Yfk7H0OLuKWbskvIVr7Xf8e8
PvBgtcwNNyKETJ2sLH4ktpFT2Q5G1hurNaiN1gBu0yu4+uxa2csqgyDNs2op64aA
9xuKJGr9YnirtubMH8MdFFyhCkLXonD9aCw2nzKZBJF27SCk1jQGnfXDFnCx6f9f
jgevRBhXi8nSSpaHtTx530lcFALBuS/6rfHL0S7GfleFeD8aD5D18pCEfcEYGB1a
RszS7VPWcHc5X7D64zRr5WcD5nm4U++uxRcHsfbSROlUCDwpAWdsudc0J9d2Vynt
7XhBNw2N6jNd8q/OBEedNEp4k/6s8YjOIZK3ykPv6YLtnd2yA7U8B53zv/QiIDcq
hTO4mOCpfqYilPdWDxfMpQeR8qfDOMtklpjAdg23lJRJTf6EOe4DUP8ujxOPolHF
0iLasrYR8mlVr4P2nhw4KqZujVh9eSduh2cd3qaaHAgiMhXNz4+sdkr7Bxmjkg77
9XVOp3mhfBGXAe4GHMOYyJtXiS98yu1GD65oO29eSrPGUF70AXEKHiteg6Y4r1e5
rFzpaOcRw9KLXxcKNewmX9UOBiSQ3tgHmdpNMMFYiFAvttSWKlZK661BAbgb220H
+6mg2q/SYcG6guGkhTzvTY3WjhfdwaLuW81ytPzCw9YLeAvAgBeYKPC9CUvYay37
A0FcV/iZVjTb0+kAC9UXOg4FR/7nu/oJopJL7Oaepl6qhJ5JVeu8xXjVgYCuiojw
R48q1NU1dXTktlZkjgSye24cwme+xf5BEsKmk6iCkXh0G0eSw0hdDxu5DfNrxLgP
HaaQTxo2ohcsk0b9YPspaEHw8HD3n5BuXxYEy7IsaXSMeF3Qfcb40f2ARv51TPeO
G39OieqhGqfjyoye8IJNtB/Gf2BoF7GwbJXqob6r++JECvOXWyBQPienITnyIaPK
6/mXlbwKL+RSnIxKhsFDUDQWl3tF9k/zvaEJpRQL284MGKxmE0Dch5e/Oh2xQIKO
Q+DoutJT6n4aCG+FioF75Xl9dfLG2waVSoapEIHo4x7xy8nwb8+rDmWKuHRQDrV/
gs0Ubt+3Qx5NDzydn4Vf7/kBJ1KF/6H0zX9XyGO6xAPAu3yAoiE7Xqb0lLuJ4WAS
N6YSn74JS/giK4+ZwAxHwnoESQNT7WvTr7FLaSCrEb6BHLLU9Dlek+4ybOX6IL+Q
yeQ89KVQx66OiB1x5m8Ks/UwzITtH9Cm8sIRNtQp7MudhNbVr2Azf2xIxZyD3CcB
miY2xyS3nz/u9lzJBcMFderGzBjJMjrteIBN97oC9ehNTCc8mMAkc4+c9UFA7amG
SjDWu8Qr6RqCfPNlCpGgNgl4mhshO+X9p7V9yw5IghaVzfv7/NTmLRTtUrkZeVGb
0AB0kfRPSmheAFvTk3zsk0HqEgZQPSfdqh9DpSFv/zym2/yJT4rcxHtGUK8s2uyP
IwIVqBxEJtutsMuEi2AEi6SpiFM4H82YnNf4artza+QiDm44+hQoSWvstKwfOF3/
YaBejJbnaD4Fw8DLpcQzk0EfCY4PEeFGEE1QKjY9Rn86R1BrGiRUFy66Ju7di4XH
ZhvU9v4jMeXCCXnr1immSUo+odkF+0lIa8GvBAK5E0rMyfPhn1D/QHRxaDdsYjue
oegAKwHd+QvqC0BB+CV7/vHfKYyn4Q543Tk3C4VHp6ViGkOA7Dt14uGTvPNxTycx
yS/ahSN97c/S7YNaJfEB4dpPp84+sYojI60LOqzhI0lwQtrAElruwyjxH2S5pJOC
pnIILvx2tD0s4eUcFdpohza/2PsCoakIgFKJRO8rqiNOA/nVGrlk4nWzt5GZFtQ0
QI1dihkDya8nP0kcaS3zBbWnjBuymG+7ekcVD+mOSRbRmH2BAkZszykLzvU6nKt5
9pC2C7tHNfVU0aAqkyxLsvq8llPCvDZ9iw6V9koUFzcZ36G188jgfPimjgtZYtCr
NFtAzHlG9ZoMGE07GyhgJD4+StcFfSw37RhunAmfR3f9dofpuTjbSSoqZqWpYIJI
68+Of91AsdZnStIhdzLmtckPrXzilkUAXpaxjeRZvImyb+CUHZpbNVZHhATC3N68
ZwTeLApYpyYE3Qz6+idZENw29vbeAB8QpNyTj/Rqm2GTq8KsazdNkekWLsTkKKU7
zwzrbd9uqcBCr4Hc2eZyWW8j0/yJ5jfSZV/NJdSUHPTnYARThZaUuCgx4I+PtaDw
ETLlXh8LblwPJd9ditf5Vmes/31MRZVQAA7vzaaxME28UaC+Uq35AByCxq4ZEiBj
cE8LNLf1BAOi8UikC/lg/Hqxztw5wgBhkm5j8x49bP6An0qg8AnyK3n/BOnko4lt
ti0QBtrjMmxNxE6MpBNFUh0cck7HmrQszIYeDnuVC3X1vQZ23THjp9vMn7sHqJTD
9Npa+76SBx/+5bJwO0R6n4xJvcTNqrtIcLNI5LxFWDjU4BDN+q7LE+ewS3Xq/QgU
ppy4kmuFNZJ/fcTvUyKEzAZRuCEQrHqzFkf8/dK+LSmk3Zvc+qulq4ECs3CTjBrH
e3Kru1dHohIKtfw4Z/PqYoT3X9kRvd7dMU8UMEJRu8PUvzP3U+c4L/ICBNnsdyKz
zpXxMD4CTrbOdCiEd5xiMpj8ueUiniHbmFlyaqtfdTxUyxKSUjpFn0cPBIf44Y9H
0dJgS6BgvmbzQn2X7DrlHl6TR06vjwazDU+SzlkCu8ZHMo2SUWoBpxiAbsJx6Cpo
HB9snlhQ11APPFwOIoRUNkoanAV4DmlqFT2u1hsgQxHMOA+Vkvsm8UqbrBOdBrE7
hEecA8TI/niIbrH4t/OzZ1lJVmxwMwZbuLS7o3DLDqYuQ/t8ySUN7DoZdy+ING4Y
E6IxP3x54JQOwrq63Y9QT1OX3gsGTM7QnNILsC7BUA4Cnq47skuHm4Y+3MI7qq+3
9T6Lzv1AuYnA0Kr0b+jQIdECDuevyGWKyYr7q1C/NDlQv1LdIxWufHQ1/2UyrFtY
JhL6QnHCnVZUk4lHByHPII9aizpVPXEm3oXhdjVRzfaWKRjnrbCT89m1VlGGf7SS
mXbufSyCr21kJPsCuaAa3WwNjoMbLu+rMYtXC+EqefGH8WrRGE1ZVUmfqxlM0moR
Vr7eOypqIrplxW8IDF+2bJuaOFiyGLPo+tsE5xgMbybGsrHKn1j8vgqMai33dhic
5foFXI8zHvzqFY8RxH4dvOaPkCZbRqvuJOwmKVTpw6fZJOyqJ92KShaWcOwxpxqb
v/VjO0sPKUk4X86jBdty9VEkwDfcgYGfSJV3Ia6DcBAsq1FzOCbY7QpyTCy17SsX
BhvYU0QKEenFh3lEDtLSx7rykMmHIepc+tA64njIis6P6oovYYjoKHs+mfqXNf1u
9r/hxWoSJM4x8NvWkZOHkwo6lZLZfgW3MDeuMHOPfGoinPTM3AWmBr+/AjSISCDu
9IqVPM/hR7bSX1Wx9D1WHOH6yPj5eYHH/+muOmQgW46aXivFa7exQVzWA4BtuxQh
Y+B45ZZZKvfa5XtEwA9eFcbRa1B39gKKf/ZeoGmZO2DF7j4hOdFEyifVy7sHL3A6
aOHQmet4AlXbSaLUj2LBX5pRn5DsFyEDRPM1ydbfJ++N+vBd7XEJlZRe6DUoduMb
NcDa58pCZkISnvM3oh3V1Q//Eatts54Qsmgst4RlTG7N8uUCk9QoEE+MvGwJFsT3
loOMspMfXkLmSWhTWLzSe2y2ciPr2KE4xiFcg97RL5QkHO+P/s9tyYMX+yoRTDk+
wmSn8wIFeKoKEACCWFRN+u80PX2rNmyEqVfifFbeCdEfD+oS0lgbRfaU5kAHt9DD
PcTH1T+/rDub7B4KqMlaBYjbCvrO/sgrwQAYNEsNvNyUnMgCb5On0gvmqZrxz0YF
l0NEnpjT3PZuBwc5cWAHw+Gzpyt972ou5/jY6fydDCckjU6dr3SjzEDOapwswR3L
zzhDoXiTZAelMhMh+ZNldsdBCwkZhrrYsGllzJk2B9aOih1qXe2bwwg9nNuT0xTl
i/Gw77VrdRWXGNzjGXK6yF98vUThpKBj0X3lK/5kiwL0PhWS4xZT/J+KHRvXprJ8
M6sf40RCRKiWLqdCVRfcFmMaSdfri105EAos07NlnVWGaQqTi3HHylzGYy0VX+uW
qNwTUxroyykot1mt/aaAnSiop+WhCSUI25OJT5v+BpTbhd72WzNLiAslDUW41851
50w6HBDW34v98WFbi/En5dWam8NKgzpYK1imbRCleCpAy4CPPM1sr1mdVjHpe7j6
N0niLxOCuXMPgIUR95QPherF00yhLDUpLRK1s3oV3Xc9B7TEuAurs/vHanCcNlyK
GlIh0t3AdPE+fzGcfnrVgwrP09UuGq5n6SxaIZrjIEf1uCMBlQGhkN8x9gBcHQ/k
+5xkeo2y0s9VItGOvbam7fzsWuhP4SFS91Q0ZeVkmHlCOdgcySBlFGlsvNpFlKJo
9UUOp6e+SdtOJ5E/sfSfsVk5uY/+vk+mLbWD16srYphdeksbxZ4E7r0JaQ9BgL1R
OD8TYz0ChtUz9iLjxuyP1hBwdBtlgH8r+muWKeB/pAhTpGDToBIZZwSdRVESxD6A
e0n6XNN68FEh8jZFKTESP6RwGT6JqpIC9rm4d4wwWN4e2EYxZN1YDXW+99WhKSBa
8KoW+/5CNEFQrOHoUo8Foo3M4SklZZOrg4xH/RemMrZGtkA1gi9/xS0/OtA0CXVV
fbzGUTHkaYHvpJXFTclaPwPr2CQxrq/WKMqcfPvmrweGCPq+hSV9nTL58KkxlKS7
j4IVQcLoOK7BluK6rvfnRhoCsKAXG964FI3f+w821h4nhyoFkNdldoCddZRGtWvl
aa4J0cZCtL0i5G0x6sYFTBR7YdN8AxSvb5Mfu+9/vHK4n7ZEw4AzYeUZKx080lkd
dfxj+dW1KDsKHoQw+PrCF7DkxwYLUt01aPJS5umBmtnnT+2wb5MXgfGC4Scj4KZ6
hSyBJeZfsquKSgiOG+3yDigtvjV2I3gxHSk4ULkA/FNvgi7rcqAczr4UNgsr4t6E
2KNVpJ30/cWQqJWj7Xi+CVhW66wdQ+rd/pUwiuW1WKt8ID2qihxU/NXbPOrygMLf
y8VL2c1KhwXohbMT046+4Azl1N9pmOQF42EulotYOguynqA3e6SB2GvvAqMX9I92
edZudORZu/OD9KrybUoNaQzIyK74yGXArIeCEa4/NBaCoupuOfkYTYoE7IDP+geK
47sYahC5LtLEponK1b/haShPgj+yg6RXbwG8vvGd4IJbaBZPcKHlJUD655K78WUm
1F62BHRGC/KLPROcB327/sRblzWc2OgWngckIse5WkeBt92pUBqnd7w+yxZP1eRt
3iLypZMRcL2E/e28xD6LgMo9bClUIZe8aZFqcanhVYaIr34e1avRVvCvdle679/g
UJmx5S8a4NwaxLBQPuOfdHwrqFiROwdrl45Pqg6L6MwSufbYFixjo8nx/ax/3ZTP
rxzAb5VMPGXTEOjvfAqq6rsbTsWA1mI9nyAB83bS1f85qOwjY6Ak0508Wz+1/vzy
5nyA6I5hdg/dxmV7yzkoP/jqfps/+Bv+uq77tXoZtSXPoar3eo4jSOI9ityEbsgW
b/ONTIKMUkh0t0o904QXZGD3aMbnoaHZDZETTvgZCd1Fjf4dz9po5fGbjIDnPUNP
kec+jCThEZVTAA43JP/c4waSqvivjAYRkJm5NLjUv1gwQCFZ8jJDoMPY6SJ9tnQ+
fbllU2gDkE3NPlfaKNH1+nhr30EPAFyiHR1rzZGEEIK4WtanMICH9HGs3E3pZNPq
ZzHAFDaYQCiRTqu3Y6pcCk3L34d6fYM3I+aV7HlWh7De7wrS2bi1brnHVf7Y7PGE
rsAjrSu7DAUewHlBmdZZ6rMtZZdVHRkAONFrMcxh+OehH7GkeRJQC90KsHnybuyZ
USUFGEA1ltdqJJmZNrXu67FDmx6bkwqRoZIn0I09wKOgwDbYZRlplO3YkBcebHOo
fwslBmkpID5tH2o4IVzTQ7iWOCLYiKUTfE8nw6KKS/goAJSMtkv29eWm6hJGuS5T
QKiL2UtK53RiHSbniwgIlKk8isl8wn41v8jzzltd5yKhGkStE7MOkIqJY04LmLNs
H05++pRICZYTMKjqEa73vG90Y+hmVomsEVnRVVv4QZSQAuR3YRA8SbOP/sNpOmfh
sFoBnxrYPNTa/67z/bkNtk85/WLeTAwy9OmNkLFWpvrxWt8Bvmt7cCybz19DFoiI
AHTkiwMsgOwlSGCPEIBmSAB9oT/YBF8K2v3wvZC1SGLPPdOXKuB7C8a54JH0gtbb
kt1k+yBqWeDR91hMlNSc+CTkqNP8dkwD6NKxpJB9Rx2589kVgtTQDyGOuAaX+dbF
zVe8430qRo6lDyyiDLjr+cWmgYrb+tb+hwXMIuNgJvrcdBnFKc97XifGG48ODvdA
+tjKbcJ5Y/fOmSpQPEtuP4PDzQ7/E1r8quaRW5Ro6X8xa89OUpPko7x0WhK9PQMt
K2QWz3uNYUTAyq2/iEc+DHvIYTJHwnyBZgdEKZYUSqmlCIICcP+EHKMkNG+9qiup
7VHLiDlXK/eoy/2wp29zQV62CLXgQQLV5A92Jtiiw5xPNf47a653TcewOsm5wnsK
AgLhhzkhvMSWVPIqycXWIm82QGixjLmy1TZdcAES4mB+VLu7jK1RtKVpttVi7nfB
Ukr8Z5QNiuYbaQDhVKAEzj0cKsrU8qOWtuAZesmvTxUHJZ/i9DqCRir1KhOR2B0s
RAQxy6A/k/umqnSeiBIIN6MfE0jFnvDlNhjPVToV67USgdxSCuFQ9kZGabI8OnuW
LwSpbnNn9TTXAH0fcp825ln78MBIjktsSFCzGRv1QvF/Rdd17Pk/iSNoOS29mPiy
WidA12WskoppCWqecIvIfzEqPQ6h2Zd2s+dDd08U/fwQptFhnivOSpHv7ipnmS0B
hGZKiSMs4QawIZAIGJzRj/cQAzbAgvw6QlnIeog2ucTrNSZnmaf68GGw4QDygrxz
tM6tcNSV3cpeHgHEs/C0WB2RFUevJhCedyDrFJqOh+z8FkmQtok6bJxpp/i6giqy
nkcroBwVTparUkRJb4asFBJPaqz2uXRzA3Nwd0yQlrpqjlVzL+FvR4UEtZSWTFGD
I1XHBgsEQFe+/J+6UDLHToEChba/Fx2KmbqYs7hJFdbfhIycCeGwWhBTTYpuT4CC
YOY+B7GgFeFoujCsO1gEjuS4l7kNtRxdSTXnvPWfBLGpeYT4kiaJXjA02xR1n8L5
z5avCSyKnFATYrkxxUF5m7v7VZE0ghfQCBo5/W/Je4rFKtCoka9L3d8Q7yj0kE8N
oGx7Rnh2fhThWupvPXEKcvuBgTC5L9UG0+9uZtl760erFtj7PrXDCuALZt7EDRfG
Zmu3X2CHs8stZPFIjTDNI3otsON7SsNAGPUzwhlYXMGYDLMbtW+lYoxDm6BNRI56
vH2DhqE06rHtFOB54FLrqCcFaZCCMjLgYrHuq2xXX5UFYevhxmQtmHwXCIPZTYBb
rFgS1o/+iqchMSG+0olN7Q0KscEsZk2qe/bEa72D2NuhKp9onZ5+MsV8Eoux1aiu
015jxiLKen/8lPMQWf4tsu/8jOgol2AqO+nw5OcH9ee5CLZEJkCfBHN/in6zGpjR
1KgvfD88p+3rV+goCDTiquqzUsEumxKU4Bt63qzIzWWnmMsVIQC3b5jWtWg51kLS
cZi4Cn2YJIxog4CrDVGmyU+2OCyXthR67pOmAdFSgYMFDUnIbaX5gNdXZsbTmUgq
CS9uzFX++ngbMedk/UCbfXRY/TTJ4/r/gNaVZQMpLA0g4zVIlsRE88dZ3iXWtDZ1
Tg7FkRafsg7RrFyrJ0I8LB5RjY3YUu9IgYXjOMQeU5cL2VIdAJvxHgXEW6A9wxpq
HOurOiR41pRD1L3MdDr6ClxmsBdV3ZHrxgxctdWsIjm7j8S7clKVsPBaNLz+PK+O
273Oamkc2W3jCgo2XcK/NuFqTJgcIvfqgE541kLMCQTYabW1NNp5mgpAhv3Im4lM
yQ0N1lBWeIpPNNyfVtZPUgLFspJGN9nvPZDfdLh9bZXasAUxlxF71tme51r4sr5c
hVik5f+WYqOTZgGcl+jEoDjAJEK07p5sDJaPB5EbmiudykIUhc6U3nucfhoEHiP1
p9PNCCqRNwZ5Jmc4ua2Xd37ul72x9xXGdSEhS36GS7yqihl9tGPIRBOpxjVcElGj
TgIhFZ3px6wAtKL9MXL9dBmUKDyYwV+Ua7C4uFBwmIEK3CdAhdVMJYAy8lo11TC4
TZuDza/QXkWzwQW1O+UZemPxML2dyyHwB+2BGNZOCw8J/x+Vf86bZuSTEtvZrgqs
eteUvj7H37Ck6lGffZvUuodijQkclbfqACeI+CpNW05+7Mac3W5aOpEnXbJV4cOl
r5wmMhrQeRfwPQqIWjyC/YJowHLoWOy70wZaqSrOkwkQIvbaS8SJLNQqsfrULL5s
IcK7Ygnm0GqNDcEaN4S47fZ/RtutYqT19eIMxh4toOzNCDxRJYuQxHjsbgAZW7O+
WVik2ntLQ7R2eD5BIRyCzc6b4MoK3nciuQocxeiMkCb1f3OWhCp1PtujkyeiH3M4
nMlsOK2z6EJMIdrDToCnbKiTaf/Sd2ZC4YZx0KwYp2Xgs63J9ZFb+s2q2tRTxSjG
QwHJ0gBAaCYTzmjMUCi1+d4bAtQR6tmjdDKZi+cwRsYCbjuyvTyvJnJyonedKi2L
82wO3Y0XDJR6KhGzMZ4wp5FLF1To7hkttN5ZcH9dvM6dkbgenDPUcJSpyW90S7An
hk3T4X3052XuT4PokIxxatMhK8S6PeFCXVTmQl8xTFBqsKtRl6gzYI5HUvuJOqB9
0er9VAwxNY59FpSS6YNrGoSENM5PSLbdye+QvsRpCWYGz5BhV2Vro+IHsgU2b8dH
D3/ANLvpLPFtJpaZVO0sW/imkV/QzrJsYnCKR8ToJNk2HsA1n6IafRt0v3/Rapyh
asQY4N5YGoeTfM1OrHYOccSQdxr2K05XViHG8AfHBQnyxhNarMy9Jg5rXSlS1QY+
HrsUig4ZrVFdD6Z3Lf5crXVGK5V7xMlaFOfAHqykL7/myXFVyvAWqo0SdxrzUVLd
UNr4FpmMyZXr+fQA74ansLKpEBLLaKK68TlY93hmb8SQU21ZlIFnL4tolBV79HS/
ZuGdrzfp4pPm3zqUT+iFQFau5MUgDpv8++Kz6epviKEV9jY7c/YGX2rKBAlR6lBG
YKV0ptmJweoNDwRei4LidzUTf0YmsR42Yhj/izx9P20ITQZniHIaMkSc+EGxSf6i
5Ie+7oMFQYaIxVhD+wp0hSJ7gEsnK16Lz0xiyUGKfDn+rdtB/m/Ak5jyNjrT0hNw
itUjJSB0/VSxpLWzxykxcyqDtbPJMercWIQfcpnm/p9DjM2EgHTl+nbeenHhAmTG
nmz7U1tOkyP9OTFh5R/UtiEuiK4+bQApddyh4ZnBzCZacIUnsznhPBmzc/tTteGK
nUgtpao7IyWt0hwSvMaWvidmu8V7LHIEODwpQvM1IUpr3/OJSmiLMLhzEZO0Py2Q
ml2F9HtbqdyWzMQg402YQPSQzRl8X5yQNvwiJcmHrM7bBDuKLlC6pfWrHFET+2sz
FFKtfAqU6GgS2BjYQpz7IHV+BDSK48hHWXBUbJjGbYm2+zIInvaRnfX9ZoAc4/d/
nqsLiMiAyz9QPpGKcTTQKDH8Yv24u5oe91vH+Qy+YSojp2qy24Pga1RbgVlsl41x
34xkwHBqWcGmNas09w4A/sP7zR9UAe3sDFcpQdndTYxiYkMp6cROI0/FivV6QS+X
M/uwRW+d2x3qqce3IbxbE2j1jKVMPcy0jz19K+kd0sWyCAdDHHUm3tdqaHLkAnSy
9HQeOjkMobDL7n6nMI07mn+ogxMRBM/T+EzwauD9nVAdm4ljeQnzdWIU/A8F+bUc
YUBJAh786txWozt9RwJp9bruPhhuuuSP2hoCgYWkpeCQtb3Vx60tmxAxEfCMcZwo
i3TyHjqbp3DpXM5hIYwnJxChAorKCADtoe0NpvdbfmpwEr8zXh2yQf2sz+LtP7xA
g2c5+4SddocbDWfLBpc7phyoGOwjpVUbfAqE248r1nf4+r1a8utMkVMb1Ary6TNU
7I6PeZj7DgCUxcAzOnXPvF1+mTnTeBa//xwlSvCtI9H5o5t5kHhUWoSvAlikMuD5
nJ1E0NIqr6sdVbZV1aThrWZ5sLxWf6MuaCX4ZKGFPOuOO489lr2zCVO/BpUfpHz1
ca7vpWvxQa9iWFJzYb5xUgOwB35HZtGnSvig++L4HlZDPlzaGh1yOSfCck+T5OTp
nidhAsgWVkANnOTR7Dgfei6ROsIfXE2gnyeLTpst5CiLGdLrH3tmh+tvAQjYN0TU
RXfsywVnfQlrIZhf+ycprsaWVErXEgCYbCdA5E60bWBD1hwEg4XiJhlIBhEB1tpu
wVcdxVTXGK3d0f3RHLOE3LGYu98hWCbfZPR5ON30uJ1GjpO8vPgxi5YNJle6rToa
hjV3JdTlZxf+t+q5KfkGmT8p1hYP4Fu/tAOAv907zEFKtfn2HOmt2fAFTpWt/z5v
yh679zVbhU62wTNAX3RtKFrJoqXXIx9zKQIFN7n+W7I+MbBn/bm2nA/bRcce+nqU
cTBtrYCxKSLRT1BwCQc7d9btL+yM0K3Y9kK8SyEwNRnOM9ZE8iMiMDp7JV2lCx4v
LNNoyliifbrbN9ichW1lrkKDMz3cwaq/X2eiulRcjE0ucOT7nRELsm9xrb21ELS8
dx4+CeeyPLAeeVSokl0yZKFESYGi8drzO1n+bCvn2koB6KBqB7w2p/ag2xC01cLD
gZzTZr0t15ZtmVAagbrmrPKRRQEBv31LLvvlPiRrl/gJFcPt5Fk6ys4r2X7L2oCr
ieKf3GprMZ9vHB58eZpsIwdtRITnxwRGT5GFgcZkeGzeEUR4CtcR92BDCuMf/Fwk
F9D+saIojRo7VZJSHInmIBKU7zieEJo1HHFHYrwwUyUJ3DyIi5tvKHXa5S9VtAJO
ponGQbi8jRmvgcUEhSSckqZMvLcIQYyaclBAIzNNq5P/sjwe5mqlPMQ2GEzpVACe
wYCqe8vK32q/rjgsbN7Ld2n8zndRUatKYih663WA44L0ujYJjUZ+lR0spDOE82BM
Csq15X9FveQXmy9EXZNs0HBQrq7grvCFODL/KGOjLiF3mdayE5qPiIPFx+GjulYn
n1B/AKUj7iK0or9nyjKUnf2ReWLf/aO4M8qSF1Cbu5a4aRlw7hHfCsAtH9LZzwzg
CFKUBkXllQ7Yt4meDVtxu2TOFrT/RuMHPdThVno9ik3LcPLtaBHb8nN/dU9YAEg1
S0w5NizaBI0f6M5gFQHym6Q9qT1NVwTnwshT+YfdlMzLpfdh4OZAp5UpDLXE9ewG
AtpZyezr7aaIA+rAzXDDV911XfVRM5fuDWdCewwAaD12gttT2npY8IM8NRKnxE2n
7iTbaL0hbogzm88GPsQT4io10XlzsObygUwLY7vbI5S7AyVGuJBZP9ZqmAQ7R+Lz
YFbn691WT9RmxSsFKQq40qKiddatJKplrQMc2sxuM9553Je6BWGRNAljT1wLoDry
7R7oRj1gka1BXZljOZLrye1WOcch5z5pFj4UsIMTv+grBvaEiHKEr5naRvisgR44
avWeIqSWag7TK2G3MWEpYMYyn1Pspl4Qjnd80VrvRd/dw9DlmeaQcOMBFw0jCQIs
OSiGlN0fsojQQRQwn8qMxw50SZw34a1dAPHGpWYjZ0vn5f6WpfvvD3lYWRTfDg+9
AR1KmqLFFBhmR9P/Vq2UUcmxYiQSDvAXmiKBuEeCVLIu7UlG1sv+Avt/ZhQw21l6
CU5KnO3cxKvKzzXetoKpdDnePVdrQdUiY4uC9zHiogC2In8BJjzYoRludU3sLHnH
w4D97YE2jkHKwqdxHPplZiNGD/bn+rx+sAAlGp7N40pW1yDkfPnTy6uNolkZhjJ8
ei/GQ6nyeogopNDf883tNZakNAEz2n7ERwkC88GGQAGghuDMMbr0zQU7mcs42qrw
DvxmVlrXm7cuxDjjISOqOE7tJn1EbVBpGwGBXo4OYs/zbTF5AaZceyzaEpXB4JcS
YmOQeR0giJhBgXNqdkkgAX2ZDDKLugOk+/Ok4QQxLAuJy5NNz6Am4iR64Y95tbvB
SzquJqf69oO4efobJjoCGFmsgFdCSJjtgQHEe7RWdWl7D6S1UVV1qaeqQ/lOIB6I
IxYftDDZx9hMpVYJJmc1w3ed0A0ZZ0tkJa8rCGhquDuIb1OGoowY5I6DToaqD3yB
dwmyeIyk5z8ACkECzzxkQMOt4/sYh1fQ2yFrfxMaq16cY9ieRKEO7I1cGKpOz94u
UOKuRYJQRVOsroJR7tMt2bnCchSeG4oYqTwUT1s5+LUf2BY7iLIGUmN7W1ex6mQF
5hFF4U5vn30iFf+Z0PngQFTH5gUptc2bo9riHOe+iB8GzivFZelT39P8ADJbENXU
m69Sr4fBF4EUDRgZZMnMuvacaqzM1Dg9VUQJ7zWRSnjMW6EJXYsfo+ttJijub3Ni
Hlbw0cKTaovsHCZj1p+GjZk5NN/e7l3PTO5r1wY3cIMf/grx7tOR1i+WezwtS94K
cKcXP4OGUW1kAau7TsTcK8ttIQ/DLp3sfTQysjyybuiI3qNSFxJdC3jJRZrcoL9j
AO7OcH186smeY3bWez8wJt0EYryUE0t8MWGEpbExMKls7a5vnwUXCvjC6gIdvgSY
xemGEnwHEpDJN585D49JLgtlOjbnOPfAHIIprgErM0mZpy9VodxqeZK47JAdycoG
pzZhyn5l9NKgkMdm5rXfaSXrYSr0JQFTV3NR11KA3swP0NuBZVTtqzMKIq+AX3lv
VnYWvcF1BusC5J8nqgGYQP+9ASIUWAdRaeaId92vGSLl6ZGMdq2qUKgSRVL4hqhq
PMj2cdmJApujNqc1K/M9/YucZVQBa60Msko1S1OroVmrSQRtCeMY3uksaeZ6AHPn
1H/n1QjiqWGmiZD2fBA3wD3cgvN61hUaZ3iZ3uyU8qHREXL/9jtO9dV+3Jz4DTni
2oixuqJg5zAO35RYKAga1p9QbH+OwkZOmcdGFJbjMIhPI4ETIdgDUU88HjfZm673
z9VhQXJIkxlwK8GE+p7nuKHCSYg3xzwD0amgRnqAEBztcOtZ+z7D8GKJZvdzJHOl
4e+uZwIGmijCXNkZ5c/PKXha68Gu5XLaVUVoz7yktGiagm+BPp1bvG66Alg4zQ9I
FmWDCw0vEONe9pJgLHNbXY8dqaSlVAgrgZFupIzhEfeA+jJCkYA1KeYrEayy2Ix4
HWNs918DByLBOOd17JkdZkdLIIlCdz6JusQw5YSpAxIOss2zbNKWrbaGPwSCgfGs
MswmAEIhxgdS38j/XOJXU8wZAJBDBJ1TtadZBiu9Ac1XhCOhw2Prqpbl7XqkvjJL
8ADPjbQdkFFip8Gnv2m/BDfWtn5lFAajHqvWFTitesVkf3G9lBrrIQEz6qLjKeQC
YZ0CTtTGQQ2Lw17Wlmcck4fCpP2cdU/VciAo1uAMV3zVDXCxEkJuemwYAWJU6Y2m
WP2PVQshXCpfKRgHbujzLQ042p9ZOhEi+jwe6NEi884ld6bBDsgjIi3jhrMZs4JA
T50Rm/7jPxLhOBAHllX7drfo8xXOcErd5ew2bW2DEefpUDdIdhcz7e6dEiOSTQSi
2caAPA2wTX8V1zIk0ds7VR2Rty4gy3+YNqWGm6hgZ4kgTaaIu+jDi8tfQxPjVTg8
63Bw1/bNoOuteQYe071Ew2fbN/3L/nLmXw2/B+v8jxqvVPb9xPWOl/ApRIDrfryG
KPm+GxgIKIpLV/MCbSNAzMJBazGWyKVjvvjqAis7AWygPW0jNX6aaZqMCXxVIC0r
szD8qLgLmw9YHQt2JCCOwS8UyIVZx0COdkqxRxH7TSlkNSlPuIyyitC/wNsNw88j
pDaYQZ8i7AO2wQQgRYjPtVdSQ/Z7MySHktgbQO2gvLwI2HxvOasvsl4jjVSFBojY
k2sGVNi21FehnI/xDSKVTQjembCb6v6qE+c48DmzWUrm+ufDLY7OzRyl/fQPQ/vT
4LTQ4WW3EUYM98o3+kbsonEEB5f9JM9DcEgm5aERoG3XUE8b2NgqKOp4k36Mtjzh
5h6PI5fyAL7W/jhuJPyPQWXoj861JZYCIFpfw4k2WEtF+c5tZKMbbHJeT6+dbwpu
6GPRlJES7IaDGCvF8Cjuuq79iULT28xdRxjd0ngAvWjZA23KbIk7ckstSmk5wbb4
8QTJgj6XAk8Vzf0BaJKo4jy4sGn4HaAN9ai4k0Nu3LJUcVNXz5vEtH4qrpOrjz5y
Mx5Lzx/eWCwZTsQ1Q8vbJhu3fDtj81G1FDa//ZpA3O+1peBzBzDn5NZLEjaMuVHp
e3OYZc9k8HLKk+N1Q/8oltdYZdj6VoGLWuNlj2r2ISI9UhtCTgfbDoF8avHzXfI7
ZnB8LhiEiJI7s9itpqbjtSA1toMI8KUM2MnpWj1X5HNg6OHzaWbU6medtAzn2XDW
3/uW3ZxnZezpWw8sMUlKEwhHOl0+GzY+Rny3jFdjRqaG693Ap/XWMBiLnt7Ll1C6
6Ip00QPSIIN+CVd0ENgBfzUa89e1shkLiLyjv7QhrmWjL003EFctO2n2aNDDKAjM
L6qpLIR67qhlUeqYoqpXtCWX/Qh20iAqzJyYGc1ri3OEct9JreVmh8QxUdmT7wxF
oBoJX/sDNUO3wYGSPc/y9X9lKfihsf4RVkro3b/hKhfq2WbrCgpSjaoT/zVui+zj
/sYbOH9dLPgefSBjHL6g4T+rtNPkjsBILz5fM7qXtBVbpqDae/z8o4S0n9GCq9JT
VvLEEwJddm4QHFjkKPgiLNxoJf9DWraEsvBjNdlmSzZYQotGAIgeh5OaWeXIk+Hw
M5mt5EEjlRpIer41PrhWMjAXiQB8WCi11yG2TgTaIQpcuIbxr4oBNn2yNFo6zDSp
jR4gv7mUcTeZ+er0TTYWUxgFlEr8EooXo2h2f4wGbzQ6JYRvbspwPjmVkZe45qck
BwoVwpxQ9vnVEQMpf17uEDv/0GMZnzVQ1CSCj0gkVVf3BD/wXVjrj4LVx5Imaj5a
fIIpwBCFBYRH2bU626a8CxsqTbpcGudBhFfOzjVrGIQdPGkH3eedxYIL1quWe3Gq
pPViq0Rx2B3VQ+qdw05BlDjv0s99nM73mjbli0zCFgYmOCW901A51UbsZvMSCYNt
iqXZmYLeYBCVYdPpliYdxbQtQj3rpEgh/kkDi4xTbsGj4blPjsojFkSi1jTf/Qnw
XbvR1SCiBIjWtNb67MYfWpdpKfuCoeN7CfYoWI3USt1dmGkL666TjStP3e9OmNDt
ayCx9+wN5hmaduUqduWpQeiIYIxlwJFfLQ5lRj4pRV3x8WLKcS+MN/hW5agjj7/J
HHePN68YXPX+vdlrRVq1uPmGZp8oZMEwEuO4Q7dv0mPvrBnSKYaxotl6ThtQwTI8
ThuFdF9idSWXg8WUpOOnIXAAjgesN2Jax8BrJjENmZk+JwtgEiDzdbycAp8I/GpD
rgtpjor0ypD7P9BBBamjlrkHdvU9pwDy9FQo1XWKQaWs9MCQFgaebUsJnLtvVzXg
4vEiqNRNo7iq3cwijGe13RStkluvwanP6iyVXev/JX7F1W17taR4yNwIX7QNlEh0
MofCwlPwsj7SuPZ5ZJfJI5kj2UTcXpJ1pdxeqVgBj5HDihuw+zb+XAhZsZs4O5GN
hfy73kvM8h722vyKvrZCyyDRk4GHC1WP4vE5nVz72zm2UBG6+2aeZfBtN4H9UDbF
j2ZjL98O2zzfNSSJqjCI8jQG4vzkzTsaEfmvbIIX0oiJvpzFlQWf8rHTwUYr1FJN
ANYXTB497SoozQldIvKvv5Je43o02xW4hwo/Ykypv9RITd4H8bQ3CjKp/JD+HynW
Xey5G4nLCvWv9UiAu3q/ZFmgzlPqdvhtFJUT2534mdUkCSGyzxWd63/J6pApPvA+
l3Di1RHCqIgXSjz31OIYwUvI0JI1AAieybC1p2N2l5BXIFcjZPm/j1u0GE2lkbEE
UAlU661Gdc15RELuAkJAHenOgK1fgxuVQZB8xZwoGWw6IJF25fWVQqa89QN85kYt
l4qPefLCZXHN1GF8LOve9Ca9Odvl8mthkpiw3afC2feZK1jguC0WvBpxgm3Rmzjy
Nb7pEvoRUP3qoID/TxcColGe9QSsGEl3ItxfiSoYe6/RHeFWt/zBXKn9tGIj/rG8
fAd0ie18fIMAtNJdFzCbccDco5tFgi/L8La1fSkmkfSUNk66spt6KmnETKX96Bry
r0N8SNPRud7XPVvK+yxAG7P0A+5WZFK/k1chI3H/B5Uj/gNT+O7fLbftt0xtM8ao
esfwdMplD1ZqTYdstIF7sLkawlxxc5Qh3oreoq5lvbkfofsGl/K+saWygtHrD0K4
mQlOCgPJXFLYb6y0Sf0tkbcwQUwP2QUUzJSwGhZhBLeU+5qvUmymgaMfKryVZJ2h
CQOTylskIqfcu+1vBf4zgDunVsCry0WIL5iZVICNv0tacE6ypRTeYs9bhvZe4zyn
l55zWZVK4r7/+8XGBi6uiatWznAyPbx+BXrmwiKoogSmCZZOQTqmsSHoYkxaIQlA
mbe1A7onSd0TABi3BeZl6qRGPer4Pibdo+qnoEMMyPpA3dtcEnaxZMHKMAoXHjSd
2pKHNCwvKb9LzODnGqMq19fmuwAdIt7PQ47THkDFFGzhmnFKmcQOdthTrb9RvIJi
5Jd47yIx5IOpawC85mDA1yATug2DPrmZLouQOTGhyGtd50Lnwmk+zFePj2LX8urh
0TnGiJkYHpWNeGNSB3AuCmXbQDhmjlgBqqJzbC+rcG+x5/7JmnaGd4WXwqDUxCQ4
cbG2TG8ZjDjZerOGRsV0EuWT7TT4qbbPp5sf6aH8DxW0he+Ua8D0z6KceEeAc0yB
pg5s63IpW2eaOAf95GP+nhLHNLGz4j5nhZvDTIFwJK1Bzdw7bOfPe+mjfP5hl7Eu
VpvxU7R1sFP9lYLJVZAKDNuHVRgCox6O882D/o3DYhtNOVN+szaZQj8KRPZBwcjO
yvYscnxMjKYAEFIpA/bsSbs6fOuA31eOgOk52pFE0cQArurrHSVl0WS8DP0ZL3NS
JwNyTpA8jmi+xn4VCZXcRN75AOmXwZ114AARSed524n9Tt8aJrf7zPcvEz4SIERW
94d0aNOkhVTZwMvlz9+lzjE/zBsweQMhYa1gfYrB71nvXZtASf+2cwR1ByCTBINI
XrK9z+Q0Kf5yukRzfKhA8BR1EgUlNjt5Kk8N7nNgCqv740M2NRBr2ZHPD/rEa5fR
/iASgaWcrGl3Fef2lPmlQUf0l5cALkMNg2dokbuyeuIDmW32hMiyKScNWtOB5Huj
GUDKVaN9B/ETZLXv0dzdvW8T4lgnIvrkbe1uNxROrPDHRA5Re7pDW7Ev49rHJ2SK
KZjY6Rv0swoC8OCYCc9DJk4AViW2VipcIMtLnC7xM9XQ+f8J23TP2SkNkemjvrnu
GjPXr4NTPbE1hB3vkhW5M328Ia0Rf17HiIxlKCCKPVAhls0HsTBWcrbWJ4w++lch
rV7e93l+VroZjBUnWdiVrsFOPQaYjQ2ivWChZ2SFCFCQCXAnuywnHnOMBNW569n6
WHU6JQtIWCPTzSaTqG0I7EVQktCLXpynjZOHePAH7h+WsVdmXZCbxLCvx5VOgdgF
aoBHNfQRYbYyEqU/U4Y1zj55p6LA/SnaJkRdcalE4JhLn+c5+bYhETcCiwAzEzpr
U3MaoxpsgSZd7/WIb23zmW48jNVe+zM5OtFjBZEHflfSpwH6zXPaMjxqAAvHPRsY
b6twdk/0kdEs6IsPM1bv6BKlgfcH8PEbsBggMzV3Zq3OAr4HQT5sP3Ya2CTeo/Kq
SzCW1y2WY6hnZePp0YTqKFvkvwf06iziM9sQUcWscHC4zjo8G++UMur779LAWfOE
3ds08r+cgd69ONCOVLOPh8uRTpYKJg/vh5d8x+r7v+/OGT8U4UQjQEwKE8QJ3hIB
LdsA7O7jmMs2OI/+TQLd+RkobGUZdAaVyqc54CJb3JJV/OqR5LdYIT6L5dnQQUmP
dQnAxFjngEYfSoukDM1Qn0KLmQo/5Q7BKDpaZaIZr7hGI22Q63t71r11v6s6fvPH
YwNFdeV7xTpX8wI+bqmLhJvf6mYYxQeDerAaEGPI7kOduCFnL0Qw3O2ZCaKIKI/Y
p4mlaaq5WM350k+eDlPriStJrOhz8pH9YHPhoisJ6O1QLC8ZlrvcMFtK4PjzgNjw
kOo2MX7W4OtUPhS2kwi+pkcy/LERI6oW9EB0Ib0r08+eeXEb98ZJbcun9plgH8G1
Ick0apJ+o11M1gSB9b/XHTcS9vJzcaQzgq9CIsgM+y7nMk50ExeeA66rX82kKvUB
hJ4ElFwbRElqSBcgG0TK+plHuc/lRtTcBdGHaX4P6iDivFCsfn6+yLrYcDc/JxZX
z8iOXGtV3G5CHrlKTiBafJh3ovt/+18QflOM7eirB4IpufITPscKvGEi4vU4q776
13sMikSbFjtuFiP3Esz0vG5yC7hxpx1R9CwdjVHHzpkh27+SEAXMq3qHsuuV11wE
IhLe6tm3A8SY9Q6zXFAcVqzkXGEZ8bJiz2WB55cTt/Ht57fBf7FN2pyxyrxqz3Yr
x/nXQBsN0p4hC+ZzoLfqTg5iOKZsVEnamw70+VizAAV3QEOUmPhJK3zfvNp37/kS
p8847QDe23DVq932giQ+8ryN4XpF7x1rtaMoj4wvUByATeBQuuLCm11blB9YSr0P
P2bY87FJmXi7RuqWOIHBfvVPMA0mshl+dmn3F3Am0bfpsdSh8CCI3iOtLkAFVwCg
D1UMx9i6XvssnrFBpCj0LuiO0hqRUV6HjqHhgm8MKP518Fc8W/pz1WSD1mRZJOZe
VA3+xRqILYBkczDo2QsV1hrkOfwJ6kFBHtPvxoXztclePF5GijwOfaCcDAVOVpYW
2vF57FlAs0odkaf4hgw0E6WhtvvXuu40Zwv4voYLrg88hrxByy7eJ7QpTrGxuYVY
pJiofuqV8c0YJUW21IKPX0XT/fyl5sqb/do2JM2Ap+FPGUvgI25EgaelublNXuRp
Y69wUpLKP32ceZOa7Crc8HBYQVzL63/Rc4jqtB0lZ6iU1Oyeo4hmKREZu0jYsc8f
7wbZmiiBFehHCGglJ3pZ98NJF2ZdpH2Gw+MSnGRjx+T3QyckhRJOwTqOO6tuIh1i
C8XqZwbAzAReB9fahKQjY1QGECMzWg1iALp3hx95nF3ucLhXWvNv8YHg0ZCH2ewn
ziB5y9MtRGFoZDuAiMZs75ATBk/c8H7rMq3anTVFvpjGN/C1ZgdUN7aJ/ipI4h+M
ILM/Z2kpxglUgT12/CCvlXUWq0Cc7X2Xpb+mZxR8cECr5r2nlJx0SdBADx2o5Fat
/0lio86ZFadwpcw3cEcP7iDD7Fd1euYbGhBNlslq5mH6KXQp+6VIC9muzC2qM9eA
2brBhCmQrFWM/BXXf2ZBb8omQnLi6kPf1cXfhJKdksgVnYqMfgyLOPeVkJIl4wiu
IyTCOhqao3dC+5TEJgXcbPeJ/+8VzvB5obEbu+kNbINmSBnLvre9iMFTm84mxNEN
s2iYXI7byWvg6goC4qGjhAmQhuI4YDGL1yPy6pkns4FNfsSFz6VFlYQnPHHr4Bs3
fixvoHK2onOIF6SHN/UcYes1jm7gDv7KDriUQJgVaptAOZv3UTzdOuYRsswepMIe
mU2nKU5qIUNRIOZgeCkqGRzNyAW/QrdE4T9r2Qh2CkiTxuo0hryqMkuRYHbY2Ctp
JxBS5PEXLfhLMaPMJLFviU6IbwMQ8pWVNMRby4nALs8z5hvyfDt/3iJKEn6dfhyZ
48/Gle+NPWerCIquwWQc2dd88cP0OnlzUPormZ5mJw5G4R6lRCg9XxZqmpnF1Tm/
7xDZVHvptYTL4qsc98QrLw+e/DkMeFKpbthBU7BV1Qv8ozq96zQYyw5xyYfxVQ21
J/imfaSVbdUaGJ3WVR9+58s6BGLS00bkJqLkfySlaYH7u0Ye8AGGME7BJxd7DKh8
swXGEp585B+enZxhZTxroYZkDLSHeUUAmuqHoukQcMAaTpLy09nUaWEXsaNbZV3n
gBJlfyM5VsD0rKy3XxUJOuf25zUGGLqhcl79AiBkeKXoctEKWhR420Yf0wkFT1b8
lXt5p6Wbtude4bKqy0FUt1zmDAuNpkYiK1SPLOyk1gpA4Im5ji/iP0Fi9zNMU9Fq
9su7zdQAWUa9Yzqu62FnzuM27EfuM4j3vOgihLiWyB6ImnquQ2eWlcXc8Hd2T1zW
fzkyMxxp7g73IblYQIQ5mpOtATXzo7APcsxM5Mcf1+7hOu5EDg1avgeWVoIe+OVT
qmjU0WB3PPKit5V9ruDWUAXYzWWS20OuNnnha6ADPeUmMHkkscDN4KdzK4SFPDyU
FIwsasYUvi50PhkIs1E5SBJbhyNwUbeZrDeJiX6SH5BVHjBm12ZDMhOE1wxoJXSy
vOIxbnSiNdHmcpn4yRCCjW2/nL01G80s9oALvdBwoIs7iup64hxkGU9QRmTig1xE
WVttjHpkKq1wMaAFtH2YAhctHgMau3T0v1qlF6TRM/hSy9d4dxcPa34yqFSEN0nL
XvwQ919Lwtanvpmsj/WCF6WTIHviWV7F5IHlbuFYkuG5ZW53evUY+lHiFOFpKYpd
pha+2ik6VRpMW6Id4feVHFpJPipIdNu3ArXjnEgHrJCq8/j22LT8rJAF3NPIwtcH
16alngevxS2nGxllfeg+gcdgt+MsW0sps9usoFI6FZkTNoJc9sm3Z3neQUpMKc31
lObD5mnHXif7rf82wEAetmH8n5nAbZpvC5YiXVdN2rGikW687HGvZDyvbh6TT3KB
2mbv3LIAuv7flQ1rFpcrpWW+OfevWSgCXGRQVm5VjdXhu4sIlnOLGNNsRW9OQlm+
81t93Y1NbpP/P3AhsDACFQMonVsnPConfvUbeTt6mizHQzMSqfazuZeGOXEQOjOK
epVcmhzrAyod6oER0Bd5HRBXvfNtnDxQopTUPs/XTVmpV1GvWIy2Mw3Q8HaKKt2p
ClKnDrlz5MeoIs10VqweJ7w8BXIPVz34JZ++Dql06LnSvVIcBh8a7/cwVF9VuO6x
Tn7Uj7RblTEu2kDfPfdFXSwgcZXkEhkKdx7KJFr6Jqn1GW4ZTA1P/ObP4erXfwGi
jd8APLO/ya4vd3+xj0FzKUNE0cgODrpz1vx8Q3JICVBgOrfFTJUkVGHVbDXkGIz5
CvhChwtrYNpx1nCVKRnfiVG11x9lTZunpny2xxBkhoJwFhzpY48RglNWq6F2LLlG
ajyD8Vx2BOF3XQEn7G1FGvn+O0a9rz3f4Fr6p1vwSKblVe5hSk+oPcxiFUDxfABT
sEazV21talcjYP2MgLT/E0/r7g6EHcW4s1dKTdLoSmDVb0U1W7mVB5DhzRpfoSt3
QooHbiCLlpzeCdXSN68GdZjsXwwztTeRMmhuwlaG3ZDdF6QKXgj/Jkb5M0KQU9On
RYGQGJgDBag9TVkPEdaHh0rOJspjImtcGFo4WjIC9MNKRC7UD1hhUoXJ/hJJy9hW
J+BHXPAV44vqWVznJT1g751i+/KJ73wuvZPvDMfDQ3cPM8m1AFLWMzPHHz5yxRc4
qei2JIx+1zZPyXFs/l+kO8OyygZAOpIWmtzIc4QZo8wM0pWtRpcwnfBGeJaMd+2k
HcyNgfUnFUk+3WzOnOuDDDP1Gx66zLaqav2u3gE2wen2ZE/HXmQDmw/V6dwz6Bpq
xoA9rdxnnacebhO1BONr6PTuOSktDc3njRupgNQQgHW2vt/jQOubnG5NRgCWq0p1
zOYT+L2HYKhYLfhFqTaVHIOgtMOHxe/Hj1pg0++z4foU0NHfwQ6Vz9WAsi9AaVFK
q+Z61jtodsFb8VqnKrC5Wk3vyLC6+81FvhpWsAOa+qdsstG6+/SofeRHRhzUZ2gv
u+pA/owuACLnoSMgknumV9jpkIdIh5CqKbsxjm+/Wf0PKr6etepYS/zoCmIPmIV8
IzL/c3SlfHTQta0wFmY+Mg1YTAHWuOh1eTiTOvIKa8PykzQKeE9cPjZh4WgYjidC
6GB0hd1k8FLxkmv9AP/PGFODYhR/GH/7PTk5HfsbeCeQfhp4K08bTzuVx5xJqRA0
9JyostQEWBAHAnOcfnmCP9qolDfru/DPPzt8ultyePQKn65zPlH2auLdx03fOPvj
4YBEjNDEAO+NPjgj/wV/dTHkqTTUXDXIywKromTYSno7svcac1pGgaHmQfl+YErb
KOsrJKgrHBy6ThCsSPPy9cINv6PHfrnxLaxQ8hTSrzOmN48RaSsOCX0cysSpTVdf
jXB0Wv3EIbOM2c88o/ORrVasSxjKjdplN09quB8hw8hKQdJuYmYk00TE7zGxFLbT
0vZTSXDL4zJemUGKBwHyKmvMNm44WUd44AZNbgtC1GCTaW06u7bKusAu0hX1PtJA
FmJaa1+DAn3OFaNzKLdFjsJ8iPLr+WerCuiOAPeSuYU2hiHgkK5VFtcLPwtgi/GQ
3+D6xYPBaV2GH7wL+2c2d+EBTKYMfWjVIcrKQI95jIPiVC1HfhnTdOONLVuj+5JW
f5REVd5Fb9uqfp+tCM92l9mNlgP83pv7Waa8yvzus5AbThS3ExSv33T0QetRWAwa
TOytWJc6rz5hFGdDQwTm1j9JZ0HrcvbyRBE3Qjm/at8YqsV9eD52lh+LuZNgaA6z
F0BnjilsH1ndfr/DhZuOwXznwYeQrVWSPBjRVx3g+lvdqVUFXhT98LRkMgXQf4VS
Pwg+S0n1FpPZpvy5l6YJOLn6rb7rj7dxtvC9GjDYB4QjNSWFXXmKT5E+3iW//PFg
c0zN956MFqlDJsI5+7RS/4dN1Aw4Shd18ytZlYys1N3okTMHq5avpHYukM64Pa3Q
vtv/EqeiDfnxeWORIAeRqXvb+oKqs0xkgBt/+iOaFkbcDFj6dnGbQhcYGUWe2EWZ
JZ3jLBXufW5P7IpD1p8umlWueU8+V4gYx2t986/NDHOIOtgliE5MNNUs9t3/Q34N
SPiLXS1t9m7UKelXObt2E2c2xREqjDKKVp8LjWzdV0cATnfIumJw9HDSub/CTNi7
4Qtuv2+zYzSMdqBRPcTIAKOjjRNKFySQRXLRbnGulN/WgPXoc2OSBFUKBYK7ROHN
d8EqIF/fhKA+M6qEOUdeXJJUXF2OmwM/DIdUg1BubVZUkyPlRn8X7m8mppbG8z2+
V68GeQebGluVV0lBVznJ/l2ml+CrxZkV4TWM1RhYdsZAhUUa8Z+HSkfXhR4zYbZk
dF5RbT30PNEMIVaYrb+FTAbqOLORkFJDdO+/dUHEE2pe9dpteFO/FMiqHAZsYb0f
zbuXFUps5wbKv04Wwy6uGc7gF5n7V0PBHhHnPVSKXHqQ86CcZaYNTtF3oOdisnCF
WhrkgxlaBQadZh7oza5jBhdzubHtUayG82kIUe5zbMEmP7y4Z/B094aY9tp995Zi
+nA4BJERCk2qhoeLfZZflwZBD4Xw5mpOJPIe5pxbRK8tlBdhOz9KXWbtv9Ck0BWa
xM+8Mx0VY2ZETSjXPho3DfYY+64u1tYHcBAQrVU42onw/gZaemd7AGc38xs7lhVe
eeXBZXYlzTAZ4VZcf1bqukbRyiVrvfUwB2gUUjbzDXfr1MMzqCggvKj8FYYZG2DE
iaRiANPTwlTYG2UvTrVkVNQETm6FlwxADxrafm9WeqUOQCUE0HBt0sXZpWf/sTQa
hneSz+PXMq/OuJlBp277EulOWtZafh1WTs/PCqGc+R5sYz8hFPbV3AJIXIChwTWF
aHEcmezQ4s/9gj0Ujic4orOYZ/avYLZPiuqeHFw/+LXssk2avrcdauacM3dsYNPL
985S5RDB0cG4iSdacVyJRH+4vCWSMCAMu/szi/XuEdlS4x5NhY4KsNuLzey9YosJ
HlxKF3rg1IU48d8mOHh17tqsmwBEkYTPuvzr7ZNyo6pjyIotp1Px7ANhdg9ViTvy
AwD1x2BgIYm/qiOhfc4xV7WM1ddK96GnJEas8g485WYFupoKLNVw95InjRqCIKEI
DdrioseBGUo71lW2eu7HtM01DQXDzAUWgNs+ChU3kL7aI6/vTCSiQWyDmFUyuSeT
0eabo+Ki7QauEXDgFHsPkdDnJlL/KuAfZzQgnhXYgphpdaIgflJiUPaMd3nwmQ1C
/islSqcph+T1lhy2K9iTOAxRcU5fdK6RcEvteW/Yf4qZsE2nBNUQjsEAuAgMLBjL
EcwUcCrnDu6lIFfe4HF8dGCnH9M/oCuObVHcdNqgtHQ/cvzzQEc3D9vnVmGsVuUD
mbFehuOHG6wKgImQizUrn8a7x8rvq70pQCcwgBrlL/YYHy4TdcL4amI4a6gh3x0x
3lXvbJPxlyW7QdyZpX4ej0gTJcUIqCnQBHaJcpJ4R/Oj+rJqZC59vHcUAU2eJkqP
mTzjs/yBkBV+U2kNCDFqsEQNBZ07kvdbURwGRQnhWubV+YF6sOWvcifWOWOXZQVA
FG3VQg5NCpPN9RzVz3rSVMt/NM+p6rfLoCOseE/pXSWnzwb8Fu6nVP2cNuZuymsh
Leiagfp0BXnJrLUhxILznNZidY8iA2n8fQl9bQSdc+syRKMNZfUIP7Sf/oPdMIWE
maVzCPdRoBgL+fFGzf3UTYyb273Pr8vgyiRikNL4pFK+nEICJBnACNq3lxR/JYVy
0KsUByUpfm7fZmvJCQn/EdmpQzctsSKRwsw8d+sXGPU34v9n4S4Kp+cnWmVCuHGe
aVHvcJHU6Zpn/jqtbZgGFWDJZhGaQNXePeliZelB/4koCyIQgkwTv79iJjjVB/63
xzmIKAUMGe6WDXawU6O/ARMnkm9flT1yke27Dzdms/ianABV5bBoYSZ4FkuoWQQD
KMO1SbDtx0AE9tlMsglYYs/mfjj/zuEkso9pWRZIST3oLxaMB2jHWvbWFLDLCNe6
DN8yr10BPx7mOyryBPxU+9Yy7NIGiUznSg3agfdtjW84RpdNiGiW3tl+y9V1skXh
4dhAObFwSRK6PtQltqiOp8qRZLyqSiWj+GwYqZrARFTPteOplKzF0iqoIb+1Z0uQ
PjGuLFwojdAQDFW2keRfe0Wz8Ahg/y4GVejeWfylu6hO/6QZbQrGNhOK4/0OZnfz
c1PxiAJKT4SMtSKMwS8Z+FaEYQ/Y8V5wOXbw5L5EO6g2HeoTlwmfgWaY8amRItUn
lJFFOXDWy6lB2TR5pGsyc8PTVNj6/+mTgB3YbB7UkIdpXfI1oWGdcRPyWs6zsAS2
ai9fDcOdZDCuxuOeYZrQscnVPxpHc5hOmM2ix16vNQ+vF2kiQpaYEZMwlFlpKBsY
akxwXBjRatqVbg7z7mUIs+bAum0fZX7kkq1KzVOgsIcTSU53+/wS2obJmjz+B7ds
cyvowv3prqI8/Wj+YA1TXV5FkMihG8pA1KAi+cI40vYTp48qyPrApF0G9PalCWQX
JAGrH8DtAPSUB8PlDqe4qZ9sTq5zkbQ9BLjqxSZbDUTROwNZ5Cz1UOiCAswq5IhU
v6mP8tdM/3Vt3Z2P3nkmMbk5SloKDSwgDedWVb5xILy3yK3oQB7kPOi531m5udg8
gii91dbM0nJQ9477JT5dnY/R0YLTTaxS7w1CjTNk8koM0oGZvwA8zJFzYeBdXbWT
5WQNktbKfc9mAZ8IBG5QLWNU8DfUMkTPmZrYQwyC+1ejmb3Z6iwaMN6LTSU0c9Ap
w3WzrZeiWnzE9SlAIk+G/qxclCrPvJbQRa1gtiaBg7Ek+VAL7tc53NJnWCfDE7Uk
scyq+enEMPRojCmeX8aC2iQTkO8RQBTqUENpl0WdY71ckozwX3a+uazJJZbRi0d8
Rw6TiUAnwK6ZU4o/zrRO/YPVRoWJLvBpKwXTMG/vSCpdfi69cOsME9nTpOU70Ad/
1JwO52W/HNYOaGOqM4wvsxEkcUqPkxIY88Xs1gRuls/nsGV9K+5DFsoLgLODcsH7
NL8vU8EA8t3LXeK8y7/2q9d22qXqQ7t/8uzYYQPQ2a+hQbvYhd78HgEnRCP3tapU
d42ePhq2Ph64suCcYwvRbzeWdOmU4CkzAtansLz7SM7jOI968ag+DPd4QGHdKFp4
ol4B9wNOiVPWeHS+B0q9g58nadIs/dwNglX/eDdKRnYAbdpq0RBSYLTEcoB4YvFd
TacFW1Lp0wSBLBpL8dGn1KjXPlo2NUq0tVvF+Vauj1A0toSrjrwg3xXKvqXN6qLZ
dqIBR4EqDgWRojSSV/yOxmwdTqyUhqCe9Ij8EljUZecHTzOkQLXY+Anwk1S6Guni
NE9rlSjjNDChRyStI2HJz6OSGnlZ4w1L2O/lPGA0YvdnEMLBTrhYLXVlOC6raGWN
/rJL80+75gnhnisgUDJHzLSNbquXD9jQgzCrC0NKGu+tPt/qebnbCawi1Bsz4E3E
JUmp0j+daltGluenVYUznEINkEDz8PVGW1isTdxSzZFrqCDehbwOiGThsOzYu2Re
SzzpdsAE7lbRH3FlN1IROzBFeEgYsgmpkg8qycc7UuwBj9FAulV+QiroSb3/vbg5
JM7UONd5Iy/nPl+2U7oUD0+HmLtwcngpaFj772BEZDiGSt98BiLyRC0fhBki43fN
qPGo97RzwuPPj3ZnnP+Q8N30M9n6MTQhylP+1QqQggMPRQmYjtZiObo593E3XPlt
KmJ/U8hJFUcPPz4DHhkVx7ZW3UAJAwUmOBTB71q5rotXcmVAxJQ5fhlOuQGsZe8i
2Sv4OTpdRHkIo4WenUj7ru02Hg5cHHo8b4ec4/GfrIN1I51Ao6o0G4pkqQpkGOKT
+VhLXumyXGU7/krckrwgUkJvp9cIkH0N95IHdjUZsEiOVUFXXlZ2GfdrvRnSv1P+
QlXyAhuH5EHxWJgMOrSYZWSOYMJqKOiYONq1F+702hl4NjCP9c3nMTtvY8rBuOWI
OWiQGBkw5SuS5R3UwLpEdPN8ufT1VxV5pRITQX29nvBGpuWiRffDTQ+ZEemAYB+1
42mU4BFjQlm9bFH2mnbvfgLCK4w5ysKaXOPf4peICqFBTbA+Mxi4tXI4Vaekepjp
mWtL655Pki+Cmz13+Uktz5yxirFXylNeN2v+pM6gu0qkLIOkdhmLYNj6NGcSpQJs
aM/Kh4oEdyIudjLsKgpWy4VXcEq2PK/KfNoYKtY8MQVEI/XAbq9vqEBsBWtUFDvO
Rr7LobjzqOCkQoo5LfMhfGT89bertuy5ppxx4cGGbsfecGiDrFhLdYbZX28JekJp
ErHmYUoOubAnDgUNZdbly1Og8ZG5mLj3E+NCxHWFZDXO5bCEBuBUi4H+F7GQz8EU
2oL84aTX1KjWfg9imuiLIGo4viy69javI57dyNwDsuBO1IVcwObiXGy7G3DMcngq
pz3nHhCSgCXWG8Y+lBCwTDtlJDb7Vg46ydcF6Bu1oyhSt3l1zCQc4yMOnyPJ5yjU
dekXcN2V1pIL83rsQQh7GD941Hm79yQb1lssyaYCYqWvqVTbKy0nUPu8IcEKxg2z
a0uhKgwURH/VQr56pqmC8SWt1vEHHZCUp2nzYXSW4XrFf4LetX+c6zv9b5VMgX9Y
S5ue+box0zn6hUQZk+Sd31mqqvGvFo4Tw05V5AwUi4nNhbr9NsSoFdtzVwCq9Lof
nnqXOz2lf54VNyXyBOS7H9YQLZRvNi4Zhwew/2TgCy0cccwbp/3E4QooYB41B2r5
SSzKqfRo+f3CnA8U2Un3s+lI6C0g4hDytXsGHqqvVgBUmEoqlYt9PCNBYc+0l493
s7tmgNdk42gM/QCO2ANWmzj8pWzvzQPA4NKjRnhAdPZkDtdwUlZAaNg5d8dl3TYZ
T1+SBAJ4lEww6i7tIOMUQyn1nnPf3eO4ijrpmXttj53FWmQ2jhrn06+bDVgEKJEG
/A9aScKJbq/QojAjUjK5K8+oPZpOP0P08j7aFCLwRutGNKT1GFKzBbHuwWVRIYpC
2ZS3AnHy+/QVhZwYhMakKBqwV03Po+Q8V3ELzyp4to8hd8sGMMkIMZRHWJW/l3cH
psZ4A/InSmzxcPCQ/Wv5IsYY3dWBR9GUOTfQiPqVFRBSAUn20sxfGOGgkgRYP00+
uaPcD99eXsaxbRh3/ocJSC4eSu/xCLZJgjhveuFf1dxWJLHtBYdbr54OsIpK7sKV
1RhyA5WZPMdCWiPkCtzmdtfl37a3QTJCXiOLqZuypeUukqInTpOjL6lPemveqOcB
Gi75KjlwY2+2ONVZbDHdmurcVBN7AbBwuZ9BGPHslW7TYvcqpHkYVUEuwxchm4KO
/fRP6knFz24zsmgtKX+qcTlykbWMcuSggSOmDxVMaVqd5eQJpLC9mYwuoW96YVpZ
pydHiDKM2TFbuAYOgmuEY3GRBVS9lP3757UEZoTzce/Skc+zNm8rP96WWEpd/xyF
kXhe333BXU1lc7ZbIbMFBn7wfKmIbwL+OpsqgLNSFgSvKksaNR98kZW43G2Rl5pA
o6wTlZKiQLV6WVMvGDKqIZJB75h11Gx8bREMfEUGnqH0xgfaJ1q22hAL++T3ZBaf
lQSc6kb15ltTzqYWbkHdQ3ah0jeRSljSyvgzt4uSKTGRxCECjwb5zQOERxdBa+WN
XaOM/+y3vYF1Rf5KjGO1zzq2XZI3g2gdY3cXdpw2oxqz7mc+1hJCR3jjBvCvQp1z
tuifaZ47ny8qmv2OGa75TgiIcdX5Bhz4t0FppWfQR4NTDA3QW3SZLvb0Fz/kl659
3J2bFnmZSHW71AIskAEP48/sTnb9FZKx0rLgKNRAuSwzL6v2Tn2Sc6si6NTAP2Zz
wXPFDC+TQnQlPaxF9IcH3HM4HjtVRaifOLToU4xMQWSJ7f9SzyOtPGQxaIzw2v0d
pEpX+IdrBKTwMAEr/JJoiiATGyYnbmg+o/pk4ZMoj5RD0rJ2/26nbSUyDMLY26Kw
PlhC8U7fLJeVI3Dw2Xd9sclT+7DRpfw02BgRywG31LtwJr+NehiJ36jWXMQJ6emo
H/XFghuV3UWiGxkf+GebDhyhI3fWMEai2oz01WMrMiA6rN9396e/ZWC7XxA8QhW3
qfEaHgDLVliZrZ7jh5VjWMNp6mIuWDOpr3hXIUP8S0O0FJBr9QZWmm1zxQkotSNN
y0SbpC+gl6qEcqNp6oq4a37zQjEuYEqXLBZceHgiWxLkmhdKZAPQuCOGJTIoSyuQ
N24A2VpwJrQH1GEox7/IlvM5ehfAkRYNMGWJb2oYX8bsOMDo6s6x/+yg4lEkgwDd
ABv/v0czUucdsYnp9Nzk35tWAQ+uO44VeRtm8Qn5Iy0zbx5+ILbU+xpQPPP+ib6s
9yo5Y0c3xXYRQivaVmm9bVSYtg+pOs1hu8EtjaeLFx8qyBIL7Hf9tzxxeScPzISA
c9e0vxAAA7Nwx4gEmF6EWywYeGtrvD3Kr0L3y5HfvNGnRfkyDcusIWj5aoevCn0t
jwGYpOA2uCbVtoVC0zhUoweyFmTN/qJYrhnt87IRa2SEhG4VCVFMq2KJuvL3DJDJ
MM0XiYgsALF8RQxP5MVP0qIGFpOL6hwRPrD6ghXwGcHoUBDu8tiND7VOcLXEUecC
85+6sRVVqbUQI/et929BnYQjj73IaHaA1PWX0leO+i2sJCAr5Ksfrf6QJj49ldzx
dkWQofGK31oLZM64IPcka/OynmRPfp45YBQEXAOxS4qMn44TxEpeDtSLZB5g0ihm
zXz0WEagR8YosEIcBUPKzV9wX2q3k+gpPCnIIrpUUo5jPNr+4cjqe8yXOCpiW20z
B4q+D/xfkC2Hv2CpFhiIg+ZsvM5btUbpI31WwO1N5SejThMNszaOM5BJS+svZvDC
dtc0lNTNtaVSEmb0flFoDi59Go2nMk+OPxgV44cKOKUi98/DPYFLO7pRDoyscnM7
f7WAHl5zZT4NRakowZHNy3dKdboz3kP50TqoTr9jXFzjv3RRGnlkvyRIvL9oNOYq
2/623acEPR+p65e+VtMFjzKszajQRwQn07hdwMYpKOf6jWSrkVH5/7eHF/JnZTeZ
OGuOuEXrRiJ/o28hrh319iI1yqhs+sFMAWNe0D6gEBtLc0e6q0IPVqGFVYS6FyCu
Wq9YaljsW2SvB4SXRyno5O9/zjh3EDUaLk0HVCjfFFopyrQ/WEHJtCI4BzpACW4p
q0UPDV+2bi0JggFvjSTA0t2TlE5ZEx+r4Nbp4WUEZhdC1UGNM6HJflsQOWg0uEpw
j4GGA9232Zq5seuc2HmptMaCwdoMARJzkSvIc8cOh5Mr9ZiI2XqS7zs6rlsWtsfF
rR9rXK0uNXqn1piJ5g8vKmPEwDjV58i14SJ7Lu32lWg+bLoncE04t2jRs7SEdHVI
j2NrqimYvF7BzYsyNB3m70Jhj5sgj/PHyzN8yAfn8t50jE+lZEsKjoZyL+8v/o1i
wFAVr93K8lAsjtMA4hbnI+2l7fqLV9dMGAlH1FJ/ulf/pMl2vUvZdPgGDE7fq6Uu
XyQRse2VVjUWwnbJ4TCkm7j+zI87mEPpY4Intq8Jjs+0AYoaLQD6D4TxWXfd7NZa
yPaT+a/mC5hJ01zJkZ7auj/q2LiOOgU+W4uBrHxx9r3QLpe0S/O9PFtuSzP6MR5H
V/5JTClLq4GcYdRe1p2Fs3PQKWrzqio5eTm9Ydrne8tKAgwYovkNIPNFTlnQpnWO
iDjUlxGYPQRXgVi1ZqVeVo32HwD2w/Ysj7h436WZF7/cDNvILxSijW1rvp7bEmpT
wr7ekbXetWBBuTX9nSAnMa2W1UCNsvv75UjCoQqlU+MVhyoQRHhTzU8NsuV9LQ1Y
n7WKn7s1sHR2WdF2IVgzitCVYHUm8WVy7zP/INzzHImw+TzZc2aAhoyWWDxMetwI
uUB7yO94FyWF0xyn9jhNFgwETodmHGs5DVh2ToJeB9BfT4DJa4wGZ5HyfzURSBwL
QWb+ZHf3G+NX7J5UxcXDqZlP9DgJ6FaLcEnoX8I2hGzy95LgxVOw2qzcE/vYMiWT
XmTgD0fDOTspX5LBCsGwl+qohwAfvkRzKIa/C18NB645yDsccfxPRXSqJQlvjx5P
FR+Qi7BKDRIjVeQ92Gp2SgJ77dSNeEBo5Mh/Vmu+5BOq4srsMAtLk4cWyL2XYFxy
5PvFX38QO9ot8qTk/QHIdjr4SHD+OEJAfq1i5irW45QnO8dqfbO1kLHVfIp63Z47
Sr67tdChKPtX7XYIhsubYFcK9A+GFbd4poEl5dFyUwSwf0OALFHy4BkPQoM3r6ou
kRWvwS0uBzQfW9CHFWdOhaE5INjFrECOQgA7Tt0tDQb6vLpW+OTSkBGwaoaJlseu
/g/a7T9xlGzh0MI4dAvNjc3RDN3seljq0bjpCXMv5dINkZtaEVqL1Fb0qT+IUYIS
F09YMrVU79JrZXQw2aVFPG3EbnmN/2prWDySkcJM5Z1EKL2c1ZxKyKx30mq/+7X0
IjOzmiZ5JN9bwxCPWuIPx6XWsPGc+JBM0GzmDEMwUBcC1QmUUhAm6Yz6K9CYsXvv
5AbDBlH/A1Dkrt4wTJEb2g22uk9aLohWF7P5cxjzQHgNFGakd+XuaxL+KlBPvMz5
4KT0zmdTpt5dOS1aEjqdboNV9XdUVGLgYoTRgfRuQjqOXWVs6NiZYYLaPAXv+c9y
y+urBfyt3lEzJyT/OyqwEqHQ62d/54bfKyx2ZmiCZ/HlYw2uxhsCezu3r4KLimOI
KFb4TyHbmolg/Yj87XlFbZMvzYr+ZU3hQfvpX4MJ7ULa8MWDVUwRxQGD8jgBp5Sy
Q9nHtgDLU9e20tj+NcrdYlhEqREnfCYwpPAwXe+/e8BVmFfcMoBK2ENnVRjaXAES
0GkCtuhvFHeFMSs56+inRbYN36roIPMSO2BbFz7/dklL8YJz+RCXmBaVY3GiU9Mn
WggzATX1fi8wxxmEK3WAvsSHQ7euT/gjm8yB5XIdPZYaUeWPtPX72tGJZPTKaPwr
dQM4fjaGRjStq12OHoE5mQ0j/8Al3u0I9hZqzUYos/GUrAN2din1Wh5Lszm26/z0
WfGJiTuSSr/YUlSflWpd4lm9hCkGnW3N6gtmfdnl/jqZQJVJHNeYA0e3/LwUGEjN
SGGnBJg7cEHiswFBHumaQtQ0vV3ORasiZIpF0/cLnNvor7fCZfessOeNR/Sht8E8
s+ZhzH13iS5ZPaKplstAv1cMUw2Rtm/QNt55hsqD1ORRQFIO5s2/QvfbjbNxN/Ic
k5NxnJvUdOFDjwAvS/JxR1CyVZhwHV7paXuedzOh2sSolzzUtRrG2biAQXWLoj5h
xVOCQrCxLBRIc708VkouclEgXvgjqfNpnna96fuHGhp1ymb6wLViGqtI8W/UGtBZ
31EBKpECYMePxGujBhHSfM6CD/9eDaV32nxLstT5d/+goyivkkBwrIX1+SghHoHR
A/e2kms1nEbObE5bhrjy/JvTcsvqLlGaAe201Q1rnoVXSsr7GTlPOVkuqAVvcS9x
4b0JApCo5XJHUe3ZayE33Uo1BkaS7Ytbj3Dj06b0qxb3MQn98X3EfkKnopsvMvBJ
RiiSDE40411/NvCA0JQCsgK0cglXzGgVDPlHvXNpXzJ3XqpyfQjQfXANiZQJYnqw
4qw5oHcWCWHVOajcrybybwr3B7vFwbHOKR4V4p96gzJ3clvdgjw4FvjTGiMb5jm9
JdEmc7CulxQuViV1UgvFv9H+1MP8QOxnrYiJQJ2L3KPxcvKlaKqYu6KV78ByRMms
DY/HwxXl6rmPhFXH2IWO+CibzNfvOqz9WQV9DbCNkZgNae9kXfbLv3Hn8NG9g4Lz
PjE8KtV5IV/Mi2Q7PR/wINprGOFwjVdQSPhKxf1w45uUoLyo4YuNZnlYLlR8uuI+
t/WmPaBln8x1ZLP3dcgIrUKUULDU3y+2vuZw1xgBTU2GAReK+KU0vtWBFtKm5aJM
UeXr8YUC+SkfuRPy7XxpKmtKVP/PlWkSLBcWpfArrcepI2cppo/rGp6VYDGzp/uq
UghDpIlL18u+0ie0BLXzkNM+0ZXsfXg9O2oye0ZDG/C/RM3uaoCFinxN7/GEf9mT
PidTm4/bgwtTdfEPvlIoy9cCc4khenq4kkVkkFGiu/u2Duk09ohWSPwjAzKvNqv6
ktCeEv6qHhhBk0mwOAhBU5lSjdkkP6mG54tOEFGCnG8q/ErtrhqFHL3uFP9W49mY
61lfq968oKmvXkSwkmME3W3bOIgd3hllWyrz6YDj3GaO9H62rbAD/gXxTUlazSVb
JxRAH5URO9PtWRKysiAI4yF+9iq/lXyJ/vhH7VFs959OiKwWW1bFIyipBoo2zOuM
inOwJpKCqdl7uRQoHv6N/iaCh4rmurZNcyLfY7GHrchKIFS5hCNmLvL2l7E2Ev6d
Kt/L6E7bmQJMSGF48iSg2FsnuxcTHdZ/uwAGHia8h0nzHSIC0aPyJUOLUUv3YQjD
niJcLenknizOFxwGZbBWC3yEmjkgG6XoPsKjvwtcZiRi0gBxkFEH7hzRlaMmNQ6T
OthwU0vUlFEvIVs6uKReQZhvVjyv/5ilFFV4niL6MxRJIw7U3r0CXHAu1AqPhU+F
z0P+5FhCZKt+HQYZOcKuPauArXfna1e5rTMRH6lv3UQm36p/NZ2etvNPyHEabaRH
4FdrZuwYSS9bEl5jKDwdY97sH+u3CQx0oFrcIWHa5LGQQ4/jSgpP+jafChAEkhH/
aqjiVQp/cUBNVerSGA6r69kh/ntTLuKVgLT0xTcpoyVFizHc+0h3pc+8Ob4t2jxx
SvQi8nsDddD8lvwQdbCsUYiv8S41RNySf1QuWoLCgSdYFoP3iEKfjo2cMuW57iZr
kHFS1PVKHZuzAC4FRzQ1/9fRzUigY48bhrVBEJsId2N5T3akZsm0GQMghXioaJRd
dzxSfUmv1dGbRJazgj2kX7Hjay6oJk6A/3DDSpXD12gbnjR/cqC/y5EMgRbXrLhM
GsxQ7tyz3/VHd5IUluGNBK8RoYJLMNdg6QoliL7kbINRasfxGc1jFzpyCYSrU3K9
n1pKvdM89+qsD4nEz6GhF9P2F4l1OxEvnABQytE4gYr1UKXiQIjUKSLj4zjV3i8D
Xqo5K/3glJe6JQ3iEsfJjrE502Js8gfxItvoB5J4NewtwzhWjrpj4BimKolC1Bo8
krBLroUG0HtF+p4SpnH+r7QJxMNWAd7fxIMGgD858yq8jfCtmX67xvkhr4ynn19a
fXuLCneX43f7ecmCtaoQTzbr5cxaVgqXxIC9vZ2iC3AedZjptsjf5yT4cflAZEb7
fbOtOjH2dG4u5JjKUdCtqgul6tP7UOJE49NI1AynR+iKPZU4BqGJPSL+RLgD+227
BNYa/S9dKdvYvzQ/eHX4RtepbdswN28AvjeAHQqUxc83cuIh/Z5lyLUquHP8wbXI
Z0u9KxI7VnA4W2JFrOO2fr9wXOULGa8sltcenOG1EOIo5xALNZp84BpKf+el0N8K
EmrURXW7E/0sRfsK+Yilex2Ac8khp2RQAiN5c1WWop98o7J16mCl4K+6ilb1Kwvh
PLWW0YQs9vRtol71sQAGfLIM/eXj4NsgTcSsPCBUKO8lcsrXfR/RyJMxftetVE/g
qGet8i+ZJwyRJO0+NU3JEs3SpXooNGFk6DH4uFVTvPwJrUoUX/oBbp3hGxypT8sn
7IWo66U80QtONTlr7+1EMtG4XgyYwAHJ5WP4evgGeAJIQgRzCmnsOmwSdnH9yVOu
Zh/9eIfezxC5ZqJ/tXWmeaXVcpAriN33B/L9ppPOqUbJb/63L14UhSm0DuiLUECB
L9NHJdC0KLyvGmIn5IckfvDSACCE8F3YNzukbL3v8m1eJd0an9NvKKmFsdqwvan+
odkK+WrjgIIe/qiB3ZPZrF7Yei0HbXF552n0Cj8HzAJ86Gm0jisjCivL/WoNyWEn
LirsG0AmKP9lBpDW7vIWVomdM2UbGGWOcRtLDvoIIYmqebmOPgSdQ+EQp++QA54/
MX19PgEDbD4Jo6h4YyoUUkj2iWqWuzhGZMsGHUcUzLj9oe7xzmNCvx7fTYagn8Oi
3AU9eaQJBLP2VDoIb2wAYjk/PRPqciVcN4rgi73WgsV+gBSlTZ3RLUT0fkD9WNV5
+1Iae/VhbjjoOksnF5QwvDD0pOD5kHV+43F2d/JU6qxLW4R6KfoRfbhTv1Nr+wA/
bjukgFd98LUNyJmfxJWz0oWyK90xTMyoX/yoOXWG5i0AymUqBWYeiWpRoQwZlIPj
Wwos7WF9zeXpB47Ivm5AiG9L5uj11Vj2Q8+yLkFQhJfDxTGWz2pRJ2y/oSQ3ganD
MPcPVQnWEuRhs21mzGL6FYZqIN5tw8JI3fHNlWRTIBiosRVucnV+/Z6s75RZDVKt
45gKngUm5zsjJQWgD7pAWbP+e+Bc7VviGUpO0JcdSAU6PhTw1Mth9GQswlYIgHa7
wpqhrF1yLrf4GLJldhODXuZ+FQh3S5CrwdkONeQGdviwZOTeJTSmEXePu/stuRPi
MG1lSSxdYThzvHRTy1f/deSHnk21jfRuGoa2c9ivlokRYQj/HW3bE9vNX6KsV1RQ
+rlm21lx1jgOR3qVCUhlLzbgBlj+v3cSKG9WbaRlq29Vj0S1L0oLjgjS1RyWKFs5
HoaGSwSTJfSF/RzY/+lN0X3kp1dProTek2znEC0rfaVPIswUVu/CdqbNwp+BXpbA
PxFwsdfMnWaSwFC4qJchbOqP0LXlQWXIm06S+C/dkmHRowyinzz1L/RaUPmh2U28
gkp7HE0Za3NO6dyebb2U7XYPZqJLMjKs9f4bhqJRikuHYNFBYlSYl+PCJZ+qU2WS
aQCj7jm94pmc1CFQszLZUHC2GIHE3t9h0aUw3WfDgMslrqmYOcso6Ucl9y6Hpyv/
ZdGXc9rmCvSgN8HgBHrOcD2EtHVInNo4coT64s3j1tL+uNiep24KAlU5oZ00v85Z
Yo0Ky+ZpE99zs7xHGdXSPUb8PSAvWOeeniaGN+asqV3YyT70pzlpD9Beg+QTnlRp
3eOgm2znWaunReEkHsV0SmsEFPOBFV6elscpsXgkr3mogvKvoqY4yYgbblmoz0ms
cZbqVvWSDXERac6xAJfSMsURKnOc3uiR5rMfe1Cz7zbs8VkAfxVpfrsJZQhGmKA4
xl3jaeGhhqq2PtImA/UGE7hSVX61LIMyKySw69RqepNfMvTo/nJpZGjUwcmkzE2S
KktMRX5um+BV4p9O1QdQLUB9iieaid4iVDWVl3ueEyrJiPDySGcYRmyqodW3Yo/U
FsMa7vvYq3pxupbvnunrhlMJ93XPZV9snsNwScsqNzFMVfXv3ax8RYmOFanrhhP9
6xMPMWM0RLeTcNSZDj4FJXVq57VF7ygWFeV2YrJQgMcauwIDMW5fQgO3VcqJJUxJ
N9rnc7pCzZIcEiUoSUpHKXgAOd//XL6gMNX2j08o/Vi1tPD7uHoDhYja5jk9med8
lO7sOHGms/KdTp9gH2/1aEiM2v26yJ0R/EACOhw/zDQHwQT3MOOdo9tjGGIQ8a0x
eqSyVALhM4J+KwqVI/NCKIhFCruJyCNmwQlqAXr9kJuDoSm2J2iZgZ9Xxw+yg+I/
gmSW39ArKunohwRiRcr7pdJsMUsqA96MDMXz8PIz7J3JoazY117jfvdqG3TpdM9i
dz9TCtxu6pgZnICPKixj7Og8/9+Qla7bxQ66RBEFd6gJF8zgWXgUQUz6DJ8HQr8j
p52Szw8TDe+mC2DTCG07ek1v8f9trXGw+jK20guXz1XlMjxjO2hrtsEouZI0XokT
/4J53tJfVuSYNIc0XTKO5+jBy84uwUehP9tfREEvp//0y4Ex/V2pb1PygJ+vRTVt
ah7IeyydGhvVIfY6iWpUbjW4imoRwSE75+2m4UUwJLWTC+37yvCKqSNKdevV6cDH
OeAAD18i8jbVlin+3jE8te9nGpTV9NVSJN2PARdAi0TUKFdSg7AZGzLLDkhxrfp/
/8y9ihZ27B9YSn1fF7RpR0yo0ZVTdYsQBtccx52c2Qk+fr/UaClqGvtXQAcWW6by
GiyVLNpxewTnBbab0R+77BuItplaqGqHgLtEOsOQeltSvdFY2umMa67yKM171I0z
/qigUh+sjampE/jGHZyIpYuvVxezmVOlHD65rrI/8kGRJeX509Lv6Opm28fxJsPl
eZ7XNmyecFdM/UMK+Yo4cMMbX7QLyYeJXosOv9gvynaabkP2ckRMK35OwpbsFwFm
xurg9BvuS5uDTlAi1D2LAhIBIpIYzXH0GTAocMl9oj9FeyRLyy630qp/6gIt8vst
A+Mw4MK/+jg96IhYlr1wVH4PnJEqxw+Lyfm9zUS4h9+AXKoDwuc25D33gpWMsfik
KsR4G1s9KyhTeXUEf93bGujZyHpEuaZh5MWYPaYMbz+dbg2lOSu+GWt8J7s//+/f
2GRWIJmVH0y+UaIjNTg/rjHEhcRTBj5oafiu26Lx7EuP1yJlvadc2WK5jCmFR+Yj
vVWScFSguiRi6iQ2cMtJofBShOU4ymnS0eSJ8WfcbfL7HFVSu8rLmJwGxo+4lV/2
Ps8K/FHtlsYNwrH+IXXV6AIHJMYZIPDNcF+YRSMJr45ABkZyzehzGJQ7oyLjKZDX
BLkRnzQD9vj4R84ZO1kg7AfGPAqb6JXqxzQ4HHIOy04Iccc8E67Bf1dvLo/sUjws
qImpmofnT/f4teE64NRc75u+QXiDS5ll1nbRr/9oa/Av/v80ueD9DsXiJFSKWGYW
rNxBJwYD3bO1G0VWRNXZkcy0A0M7Is8BMJQMzEz4Noypbf51IWKS8E7X879iysPn
ypdz9iXEiAROgOPLfIC0X0x7xXMGPlyJyZirjkP06iw+2l7jJPTuHK391hxdBTIp
NoI90KhCO153g+vwDJIE5HoSGi7rLvYHZ5zeI7lF3B+rjj/eVxFm3Wi8KheOkqhB
ivZpr0CyOgB0HXXLPTP2GO1FMMSIwx0owHt6mhCcFu1vLYCV+pb1252mDoOWHNdN
JAqivAY8Svl5iKsIV0nf7TGxxkwX+WkPU4y9LndaX/Xhe+Us4tUtQPh7+CES6ZQB
bSvjP09kRmo5ddmoz+JUlcr9zRN8iEd5FdXvoVfj+Q7ccDNriBJgfxKzwiUeRNGt
BCNNSQP3iaH9yU29JKnD1Hss+zuhltXMBvQ89nPfBBIbpZlaLToVm4xJDKsq6+5h
UW3RtUN2h10ZSWl7O+k2dv83h3kYfpjXR65BKGBzylxiRXaQKL/WiD8qCIONNNmy
SQrcvzy3pJLCGyk/Vtl+85BvzrFnr7wh6Wk8IM/GT+dOPLibF5kJPI1bQDU94VdV
0CT21U57MmVKLSyLc+Htjepa2XgQ0hg/qdKFzEqbgmu4UfFCDctuOYFhF2XiUVR5
UxQgnTiP790Horae8Lqdd9ipUm+n+n02u8C8wXYT55wFeSzQBswIpnUUv0N/Dsg1
Dl1ltOwz9UNgl0WOdNOOtGr09sx5NL2sCJTFJP4YnGzDWeKgKHl3LMaFpDaGiA35
HHVwGFILZbgj0NaTB3vz9dsXWoSJqULJqzLNWcjADl96kq17UcoZnfQbXlyhKxfn
a+Odl18arxh2knsr0DksYAqKqZzIQSSe+0QoLl/nhXmN6paEfdR1zgZCdmBJ+1X/
VxPrlqHH8Fkx+o1auWUjnXMrY3C8Am/9wXgTQsuuWIRBYq6ASe20C+9lJy1KkLu5
56TQA0yfFYJU1Z7FF1TRxQX+zTvQO7b8ZAgdhyUTmxpFTKcqpJGIl7OXgSNeTifN
UjgjXE0F+19jHjVJe4tLJO2yq7KXxVZNZ5xtKO2Z+/nDqDT3eyV7PCO0iWlUx8Fk
qAGvnvb4a59ZlowPWDr/ULozhXq2mjR+luKJRD37ijYCMkLjpuW4Kb9aI6irPKda
7vjRpsQyYxsXJMu6xXGaqSyX5OOhc7snFeH8iXp81j1mBGpWnuCmnJ8NiW9QN13d
EIkgHcWTc1jKJsNBpWex8ZdjSz1UGt9iqOkdued0vEWsiCfZgpMn/kJ0tfxcpQX/
eQVan2Kb2nWLeEM+78NSXHLwFFFgrXx1bJSGHFbCRt/dOxRErub8KMdQotK0C5zc
Ht50n4N+wvshcGmPf0/d2xjJm6qSVWDLPtPILxngSEvg5j3RQebxvWx2AjcLqJaa
QSz8AZ/e3I4l24qtBvLMaQGloAlVc47dkPa2IBNFRCY4leZNUiO/6l72BHlSJLwf
C0Q4UMZ8otKGfnmBkTYp+jO5bwLncfYxeDMwtWTBFURLhLsGdlFilenaKyMo65Tj
JX9E3kf8+hhRCqQCQutNuJ6u/xsrBmJwTuHqjcXo/a50MFDO3ZBBwSUVXEtvm/d+
y9rI493bjan57mP6HwwTR/OSeUg/kDkWZcczDmeXgHvuLzpvRBOx/dftKXbT/d4B
YXS43WRYmMENIZZd+oRiNFx0N0QIB4TOU5+qrZXzqz5LE5RwpNgOeWU1fYs3tDAL
eJezubGL/qplGAVraRbmvj0uZCrYKlrHzs/RSrHOzBVTINpqJIwQnUcapH5duNeO
KquEN0unwFLqEzP1A3ROM5D4aGeRswygCIXekg5h7jZUs32kU4HFGIgE0bzCMLel
5bOkmr9/Bv7tZTQjdSaUn5Phr75UkeXxbyjFtcvGXCDn+GezzaIN/koyrTQeT5lY
re6ZmdsdAcOF4sRjWgBV744365nSdt9C1n9FRbr1cDjaLehi3IBcjIGU/CGq48Vp
7r9sfzb/b6frjStZJuCf6hfCbA+udMLj7AqyhRtfHmyV7OOi8PN24LNCD3ddthBS
aUpAJL0ckL4uVPX2zIIvK0ZSFG8kf4ILOa2daYEhQ7GMCm+uz+S7irsdpkFBXuKB
7rQlwee4k65R7GFmN5jZ7PQDoARt92D84BZNB96WsHupo7o8CB/XChYzvYN8DWWK
i4FxPYXHM4cHpfSZrNbFtA9wrXEDj13lWZLWDI05CTksI+nIHkMwrIRQwxphv35a
LOLlf6qavw4eo1kixK5Gt0XESXP1XX0ggcKrIJsW4sCm1uXnL3+QKyfUGq9W/3Zp
pEtvlS99aNKV3o2S4Lh7WwR03F8kX+HupsYkIhir7AnflJTOeGp3R5HLK2512Stc
MqmeyjNzKNmYD7sttiTQXb+VnGJ92BayzUJzY2z511NTS4duMwbAdXbKT7VRmUdY
qsGJL5Fdxq4Rr6xptGxHmjAenWAn6YIjZrS7SvAgUADr7Hbl23KxgzgngzvedBZe
spJlUGMhmLIzp3WaWadLjSdqW/vidNeNcD/+5bOaRRQPwGxbeooZNvrk7ojZ9UGU
g6ZQyO4hPNIBsKcbNH4gEwTRyXDX12wDvtgAwzHvPF5YUDGAKWllZLTNcvK40pIu
snXjsTSVec94/EJ5ugKqIzrKDdglUgwudu7Eu8vhujyPNZ+0VnSigwKQ75SRCBNm
NDr14cSYTrSl1pS3nzn4ncmYDBT/DRGegtbs4z+x5hOyqwq/PF3MNeX1MCrx1MTg
8Txz10k/xccQeeExWrF2cDNV3GPWL6CjSMhocDEDkqGwKtDo+GhPME7M+9YjFlzN
+yJEA//Chn6R3SKS4cXXTQHk0xnF79nZ+JklGW0+A0FfSTRP7u1cNvppl8xRK9/O
SmGduI11RaUXn8lubSUY8OjRz2g4Z2uvj/EOjY/njS1+I41mLWKp4e0QewoGSGYv
qGonGyh0tZE9fiY6SxzkoNa2ikDKZG8srRoKP/rrkgDkgXSw79uBMdM+fjUuKB0r
xZqkISHPeO6bEbfUGPFW/eINBP1vaOkmhbF+PUXGuMJxV4lyGUe/ec9H+yBOmn52
NVp6ZpqKc2uW0Yrnhg6DGQ0d6YBOmwD0q3S/mW1iBAfaDPOYCqL3dsYjnFrYX1+V
cM+Ekr909+oKDFqTRPAS9UWEf9aLeMhO7AbavUrmlYJrKH4Og3nSAxcMeuH5wEpx
7/3F4xhin0wBiQAv9qxPwGEbm+jsM3DUhiCEdiw91i4Y7+7DYyqf3r7PCokYygp3
AzPnA6d66KrUu8u+JiM1QfSKhpAXqPWad14qHk8dZGbfi9e4TH0JciXl682ML4/I
/PHO9lnQzQsSGrGZcpcJhIIToIbspuWUzwWGc7XtP1c9QbvOCijoWB0jlwCLHrH7
B2POyCW4Y/aAICcx3gQzenRGDbSMfKT8ijgQtpKyyEw6GLhqN3YWoL9OfBFR5E1Q
/jO9Ie+9p4vNYy8hLFf6yAUhjAhsCvEU+jSnlD/Rw7UzNZJlz4Lvn/z9nsgYkPmx
rQmsauClVY+9Lqj3WkDzbjoR2rnBPimrbOrJeWOoWZBWECqyOYPvlOyhXd0e/CDe
FdOQXVQoN4e35EpdizMlM+LcOf+VKtZGleNBQUXusklvFegY6UiV0dAxWoEl7wBd
sJCBL026I1OxLZkfwuluVUDoWsQVerNGfyya8IhCmI9BIc4g1YPdidBcEWIKThDI
ehqRbaqBz+/cHzIJ+ZnEZe/BXDdaPl8zIjj1B5lxT79MSnvtEQN3vKePtIpsFnVF
kifapYKmAMCl6yiN35XFVD8/NKta6POmXp5hXIsVNT/XyGRkdsXuiNwhujoc/+Nx
dT3Wk/wVBeLOixayzDbSSWJXAxXAY7p5ABDw+UM5aB+v1YnB4KdFD9QckjnphNwF
76Jtqf161OQLrV4ozhQqD/OOWTnXpvFl+n2fBI62xGXZ2b8WSxb0BN22deK4eg0v
KA2QkhIzIS164Taj/rfakJ2VSnxznHPxLE0FCeYghiphN87vbuSdKkjDgj4PmIg3
BX+RDfL/6vAMiI8X6Q5JgZLVmT2B8ruBm+rBR5Vs9dl6rr5rtShVFWVr0YSatYLG
lBgaViWKNpk5LIJDC/9oVMG7vKHuq++4vswO/5LdizVMxG/R9ul7LV0OLmFpUl8d
JLXPzYso1jJ4KICPQgstinJ2pZj+jWMAMhrDXcZ987G6XghgaCTzUt+NrI2bkqsm
2f+BaC1MvzTC8Zig6gWIaG6OaUeIm2VJYZsr2JrPO301RmUdp+1R+yZvxgnC5TSR
F5mpV5c7te6kfbDnEI/bfz9URWv/ra6Cdqbo5YnJa/aqEq7fyMuO5NuFvVUkxlbO
Nqu0ML/DcxVf9ydX+DdnEsvFuvoGYK0VcWVVRTviIqVErSlrdsRijtsWKOXAz2h5
ZwCaLvo+Xh6Pq5ZbMYaozkYQtMeyx6Db47GKyP5xYrRY5JEYn/OYnbtXj3jKLVFv
cp13b3ylv2g3kgbzwEr+Sn7vZpr1aqbl7K+S5mkKioBzIT4gAYDcPfGMV2UPnZo7
MeZ2l8eue6oTbb41hJNdcGWXbluDOtwlwH5n6DvD2RUmlwP4dSZNtmABD1bjlDBc
AiphaS+ypUPcJiEonmMl4VkyliU+bGFRJLRYpSvLMffZBgO/vY5/7E5vVDrm/fgN
M9EJcBJnwDytrhQ/hD+gMDlBgdL/aiGy6Esq5rlfEgUlmqrhf2ORrD65SdVoniN+
FKXHtsUGsTTMjgPCppNtROFutBIXO2YJoTnGD9Jwki8dvX+modCVTKXbZwm/1oFI
sKhlGcTd633tiwsAr+wLzQhK4POpy7IyvmjEUaQhFdUTMn20STiV8e28b0QR4FiE
Ik0u1X9ZOQ4ELgMtkFaI1byQN5fdFTWufiSllR0Pw2UrzPv5ClPbspKiOZ/uPyP0
FUMtPEn/WERgptUvPohp2nRulEvEgYpzNO89AeYns/TAa8RZIiNKjvCkrWX5ymby
N5owFjrd0gBdhaCzZ6pko1faeywEMgSA59Gn/hfX6ZRxcdnwva+nPLzqMyvCyh8n
1O2SlFzSREliY55b29ZqGkHVeid7kSC8iWi8A/BuoPV2eRtvrz+PdzPO7N937u0n
kZpFWLYiJDMCeCCgqidpdGagsFFUfke2i54PSCdz7RkFEpbqV5RpYqHCQ22ggHbb
p4H97AmNz9deoMng9u97aSvJTnNkkt7k/qmmvGXqWOv1KiW9G5zLhnsOf0hX4pvt
YV8INcy9krAICO6hi9AeMFLLltuFD/uA97iUNcuGGugINJudA8vNHJc04wL7/zF6
xl05CQByJxifJ2cJzkdhLGbEhPyiVcdOGMxeU5u9whUUCbkfayVA+xyhClG23nya
hLlJ3UiFvQ/Z16feoOELv82V2Jg++ZQ51j4HDrW4hnFF8BA65N9sfSLBBQjL0Tmw
UkRHW29jlWbBswqgFPhf5J3ctieEGnb12MKsRwkzr2v/F0cXTLKp4ZGzwCOmYrgf
FuK/Xjc1/CLOvn0duE6lz+ytrKmMEALs4UFf2l0M07x8TSCEWCxKba0EE2103VoD
57Hgj/Dc75P2DzGyGEHNF3Dq+efd2deqTlvFtsNbp3P5xWduyf9OZb/qt0oa+PTV
VLTS4iYuV8VY5GUe4sNI55O04DGjdVyj7PiSvo1yCkYzZAgakr8vyCJWq9SLQC7j
j64QXXk+0RVjSdnj4eeTP4oY3rwU9SXVCvUlYEE/2haWoC1lT3Bht1R1uMSwhdII
z/Q3B40IOXGYoqRgnbtImzmSpCKwDSaVfSQ2JgHC2tHcbxaFY2iQ0wFz4sDkLVNL
gzb6nCcb/rcge2UKiFXdpXN/Y+fzWpK6gYptRopZZKSqRNJj43NGW/IgxvQORqa8
8SOA1QM3/fJ9qoT8Yv5uPmSD0hgAV/LgykK+21p64RGqAhh9vcbBzcG08j9gFy5u
rQWkbEgj/GC+MaMal5zoFZTZkb1mBs4BlgIRDSmOuvaH4JfE4sPC3ZT/x/R/Gov0
/1drzoB7DeT9JsCaL7LYuLxHePlivZ8Ew4T+eLY7VSvWsHmMc22xB6i7pD7udaO/
9VGYAlKXz001LhZxuXFXd25IoiU6jfHKGY726+Q7JnBp9r9cz4YRJ9snVlB1tAwc
a0mS10Lu+F8eSG3utvC666MW+THQ1j9VmsvSMXXWTf/ZPelkj/4VvNeJXhgz49QL
IvaETQBdnr+qTFDd0ls69uGyL2DrHbx4tn9dzvD6twWN///AJajxb3y2r97RlONW
O8dX0bDL5elfACNppIRKWtnM7WQhsBhznmSE43cjp4H5EcADMw8k2tV8fkDLtHVo
9rnk8ILl3Ah3Z39o7GwNcxEAjTBVgfCXKxMahk0AN2c7qP3VPrxMoV5/xlMPrm4p
QNpg9yuaEVZzd0NVavUiHVQsFVeXjHs8DLjjVMRbHrGHJduRQCE3edPSeXH4+8re
w85hxlhq7SA3wppMAktQXFhe8tLgNKD1FdWbICQrSYHauyPPSvSRp2pS8q0SGxZ2
pm6OT6wIbtHfwWLAyCKoGls1xH4MqLO98Ac/XITriPGNGIkzLLYUoNkWy0fbep47
buGdYESlcuLCg5HbtKSUzfvkoNWF9ZcKqqD64KgAvnWgr+05pBqsGOG3cotKofdN
EihzB5Qk0c1h5Fx2D3sBE0lHjGGS/54GSjRvX2Wj/kwxcigD5AuGDUexDPIOOHlq
fxwkPCs8OR0HAbpESV8hxiP1X68+wUfbSp1MAUF5FI0LWYi1WF8M/zqfmEBteztd
VeMl9p4WH6DtDM/menjmoraswcs/rcOIlvP/jUQKdYQOK97fjSAtTpHrCJd9yrdh
iRE5YFVZ4nhJ5QPhDDXWC7N1EYERmcoHaEO5xgMCy/SDXCv2uzADaoZt5oEIHbco
ODOL6KOIwC69IZ7S9UNtoxGlcAWjkjmnK1WGk9nWsHyG2gvjSHmYT2wnUrjk+g8j
270dUdto/c+SmLG8Axfg5teOIyf95KknL0vsoMBe5MKQJCpd3W2PQAcCJWUTBQIl
81AWbNLdmeLus1VdWdATZa/AQTuJyP0IYIjgeHvwmF255dgNqXZ2N+ZN9+3d2HId
WPRfpqb70sGk98JMTndPZebzHBie1zDlW2ZvasdpT5gPuqjLwRvaP44l6VX+E23B
FWASqDBEPOCLQJu+Y7s8HbvHkKxjqvTN74hbVptCFCMPeBFSz7v62rgEfFwHYbdT
G0rVr8AZAuGI6cEK5U/2eiWneHnwoMiH/9n3BcKid8F0wrOWLrarGRh7n+ZWTuKx
l/jB4gTowFRHwyZBpynffG8dP34Xq+GRVuD+x4OcQayfQCI3n9R6Jn/QPK+18X97
jRVWrijD41HDKfV71+sIJTRXzKk7uAzysvaV0jEDtxK+kNVwLQiKJ5wpySCcx18u
1Qt51WRmdn+tweMXuEDXuU91KdallrWYvF7Mf2FIhYVf9lEGSvqz7wWEwax8W1W2
WnRvx1/QhYmUtVqR5fc2qVQ4COQLv3AmNZyghbxhHz06zsrLDfTc7/7FsoIOExMr
5lYu9u8YVHCto/kvBoVuhkP6v5QWY531JcCZe1zfXFZLG6wnt3tRVz/GVUZzdglj
Do44bTmuU/go7/HZo2zdAXan8cNLxLy9p/geJKb3k/ibfd0bzmFTMp7eT7sVrx2P
yQxcMiNq/fbPpZYb0UOQAJZj3I+w/Xx1UXjwu14MGVo/haDSnGqjwLMV0T3xDVED
8chco0Vn9pUbyMlQOXBwVjzeS1vXvMKDkM2O6rGpMrTWt6HQcGb+1Gwq2OVAotk6
O8XPQSgtTAUxcJVHPiEU5o1MfwsjkAMh5m0YT/ASzW4bhnSBKF6F4uDV+gjvFafT
Hxv21+Yl4PCSbMV00Qj3QiKI7fX4HvQU/IEhVdWQ7+1mFIXQo0ol3XcCTgUkKh8S
En+Kj6dEB7lDq1L+Whwt33TAp14qmWab/7lPb0fvIZKFkvKR9b61fFbD3axPakGd
BSxBH18wjhL4xofUC2HtrV0EvtpvwUGzhXMDpwK13RMU1TUBXksNy/LqzCgUb+vG
A5j8F1003+mrmtHyyl27epfVsG2VX1yz+6sJo3Po+c9z2vghXqg1okB3eJiTtsJ+
kU+1Hl0B1tqEh1xMnhITEDjWWe3RJHxTVUiayTTbh3IAnRCJknbQMdxUiVYDTV7G
poSXJdIe6hSzgEoNTJ6i93SE5AAhJtJILRwm4y7BU+zrC+1nA2coXaho5yqgwUBt
BZiIKOwFsyuVoQDkaUwMFbQLwsDUaJEBiH9Burt999wO4HGhAWltrZFb7IkNy/Ad
a9uToesEulLCLmfjEbaHeljsR6oYp19mTJlGyDYC9xKBffSbcLfGAAcQlmGi+krd
kUmxMPfDv/EF+JzuIcBGsEcIM2OAhCfXOQZAl6pZdysQCo1sR8C0l2p3APkllrQL
lOwZIXFxPBszQpmfU8r+PLjP03BqqCFLajvqIxcrC1sr+i+F7BKL7rNjIdMWbGY+
AQGEBCQd9iIO7DITtOoJ+nKRAaOwDhvxHr7XVzoQ0yVax4lm5d2JuvSF2CaoXp/X
xzSR3XDfM0IiY1jK3pwx+c9WQ1gaTdkRojpT4ON0v/lId7Rd0F0uWJGheP/vTCjQ
pUxTGx8cMh8LwbHK8VYfcUE3Gjja477vfNQrAEDNCsg/R55Epl7g2rEhpuxznwtc
yhZOuZrA4Iwu4j4hoxNHBesH1UvaMEu8OU0/gMIkaTn4z+/1RhFIdJ8PDsweg+MR
HAzmnn04Qqoq3lpsRPz+DpG1yx/dnjvAB75lVHiR7q0wFFyeHT+mPOA+yYHUVqDN
sCeEkhlN5SwC6H/uOdVG5olmn0LoL6YigjF0E/6VFj9wYyLlPXgeX+9zzYZ5/da+
xrXcXe3zxir2cvY5PYpFngXW0Yo9jc2NpyN/Hs8H6aacFBDyE1PgT6aLNLf4tkWB
YCaPIZwyHlKLxVkq3hbGn/KuKYm8Ln32rpEh6YIEbqCadnlQp0ELU8XQ3IXWCvRH
4Q4RzNdCfZrSXg7OjsO6hP7ib77sX1Em7XY9QH4X8hZAGBa7F6aDyZHcdMeH7PJ/
xlJuIf+Lw3dPQfjA86LtLPRjmqKGbg6LgHhhyH+CcqOLu5lXuYtwWZJZOJyiE3hr
0claJV0ML1Y0bK9MvF2WLHOxTSS5d8vQZB/LVlluLJ4+wpvd1S8nktWSXP0FQEJP
k+VwDG0mJBSMJlUS7L+AZFjHy2hlFcYOFsnbhku1FA6anWg7/P207zch6xGWBkMj
okobz+5tXhPeY2bGR7eZPEiCXb+0nDPvry6EFaLXyn/XJbF9RVLvt3r88lpV6slB
XRl4RPPCi8zcFUHPRAegiU3F+S/UJfx56b77GHl6q0nZtLHcRi0fOC5LujQpJ0Z5
uMMr1jaRaGrrSGA+3ZQA7tv7ePNnO7hcYy/cXAZvw102MrhXvMr74OMdv9N8QALH
Gb7h6fAsSgl3Tpitofs5drPz00c8Vcp5Cjv5Pe2Mc3KGYVh2Yhssbfg1HTjTMSWy
x7j+VcEJyVP5D2dLPJQFdhDHD6y416BYckIfnIIV6GmDnkPyUOs+NS9KQ1GSNnM8
8hhJf1XDzh/j5VtgehkeOeWYNxt5aKT02hCNdf92yt/0z8Yuspdu9JgqEUcH0nLA
kFHl3+9YNPtQw3M1QbtbFTbgWvsJ2ONUUM8YfCk3rANyocbitq/QV8E4BtpHzWdb
0tNSXLep8RSLp4retpNeWUOabu6vi4sj2Njo6wW+hVgeGMEbK/ZqBx4Y1iIliYgH
wvNU4bE/30zQmxJ+cBk5wdc+KqXxYE+W4PBpmSutzd2aj5UHxkUdvceriPtB8pAP
ee3+W1qkWOfnxNE0xhyfGkRP/4ObaYPnOksTGR9rMJ+8QhBs8i7KexD1FHvfFmge
x79rrQw+Izwy6VFx91kAPCvRoYQ37z6h/AVTfHaU+rIekyAAsdRpQL1EQrQLKo+4
2T2CpbUM/0BAVoRkZa4ZBHJXr3D6j71ux7J1X/bDZoetIS5F8BsVimHcBoMSR9Z+
9YACpB8unP0hmhb8sL9ys4kIl+NJeRkYXY+bLMw4f/ian/XqkvNv+MrkGoxKYE88
NSPaDvjzOFU3IDoIMlih9Op/RnXfL/wcreyoAGnFq7BeQggamUyskhnP1WU7sF6L
HdcKfRwhHwcCHF1iXKFOejnhjOshvsh4nqLSiFU5G6/7AYzaLZWirlrHkX1TGhz+
iFriG5fJ8S9MK3N6ulvA7KV2CiOm3931G3RfkXsCg2cvFkx2A7OO5qkOC4naJV4l
7kFC1apbtlnqol4KVr2PgYYVV+uprfj8Sr1exmOj1Muaryc6+X7if2DJ9D+gQrTv
V7cNAJa6j5S/TtBlW+x9tu62eaNFOemcHPIXQe3pljK4WaK0ipW4AgP9gi3jFkEN
KV2H5CdV1RV1JNYCQRBNZANvUpevSxOcaonwI7P+QNARCR9trvgoZHN8dyNvLGaF
li0JGhurg0IgOSRUcQKQ1aTEZGOi5DLGnz1yH4IZI92DtDWVlXuV9PQRmiDbHHi3
AIcad2ijrW5Hs8QkK3nt/f9w0ngE1ziQoqQY+jKtIhkzxtJxwyXImp6U5sc88cve
Tg6rG7j6GfiXjgqJX+6r8tcNAcWa+lGLky61YnrSYGBIooYkGakqTo9ZmzmKWgKi
Gzt4xzYeJRUsePJHVqvWNUkfwHs945q3t6HINRVr1tPOlm/LMAeK585fohWWeL4R
w98G9m4UxxqtcwS6M3B9yOwP+4drQrxsQbdU0jaIQM5s3iaIVMiP4nTgP+q7fLLK
deXXRFhizAj6yQNnH4AVrNdTNap8alOwBi/yB+iTKUWM5KADymupZtoQc78YO9lt
EYtTMsyWfejZF1H5gYxywjIp0WRHk65Kp0zqOD3a04PPanDGlMdz28vUnRYoxgNP
GvTf5jZeGlXlhm/UdNkRgxVZ0gHHEa9gfZhlV9kPa3pwSA50NLLxJY2tJJBkd9rF
69kwnq6zkhLaxtNdPKQPhdVfybFEAwPYt12PzeizH3eRA3/epiFT+r8F2qn1I9Yj
J0jNeVg3C1UOmffbtrNci5MCLdcf6mfnT6WpkNkqLbEudrY60PiLJE40BofU9vud
VS2XGU9Yn5VgcTq/VClSb+B6AI8Ha33Ri3kzCaDufJ99e2rAyyGA5cU9YqnX8JpZ
E5iBmw3V6GdWnyl4SH+gA2dD08GcGnr4Kksqef43ABgE9peZXwci8+4/j6wjKBFZ
vb969vLP/BvmF0V30t54dzbBfiRs93ExHkO9ZMohkNPnrjyCnb+jkaL0GOkEu+Fb
QX6Z7+ZmXV5LULF6Xk8EsNX+tpN4nXWYN28KRRnUzJM1ALusOmGuvIohHTG4Q3Gi
lOgaxsbONIYar++6xnwQR3Tmby+dd1OQ/KzZXae30wnGQyhszAjKwmhn013p1nGa
iXgZzlRuzoCJX5fciNkzjNKPasrM3GiiUUSGEIKgdOiVR3cD1orzSmvR4aBCqapu
DD2o0mPRZTj+58hv/MWA44q5ODIBO/4wI75yGylTQIq4vrX4kQH5gU32vH7eKDHP
w5UcTonXrwfc6wVRBO81L+kIdKP2TgcTS9Xu4FHXA+FiJY/IcQlcIMSPmjDKqYL2
0DlE4VC6ZqnnseY7g+HV+PxFkTdNdDKmLut3yANN5EWzsRKJ9MDye7dy9nIBSjOP
rHF88/cN5ypZW7nZoXlV9MwQyJrzlstUAsJJPuCZ1hxlvhe+wX7LoQ1j85dVGoLJ
Pm+JOYarHf2k6HUCsfOY2SMxZ48AmtA6JI3Lo5Ezwqlx9elYe1lMMbHsGYtQ79W/
5YjulipDiWYziJ4TE0X30alpZlaW2qgXDFI2Swm6+BMgHxAvhQfhDugM2+enomXq
tSQV9nfLQkvdaJ0xXR4ZEQdEbMr9tSfBkNqK4rZLPjlDQra61ZSgTE/OVFDUdSmi
qf04kB05txhFsPWBWdmbY6UQ4QTouTrSrO+nPQ5sczxTAjdJ8FoMnvDY40c6TrwC
SL/FSsxYg7MI3jYtlBCaXWsc7/fm65V51JyW6guGK5kElbXGTT7IPtTjqO2pC7/A
LlFzY2G2KOK1vTfgoRc3dZGLtlJpJL0q9OIXD86qA4nP6iZl99mkp5n8jofYF5ZN
01RbE4KhlUutEJ/9YmmUScn7DKNfOlHWd6uUqOqnkNUXeTfRij8rDpR7648WY6cQ
+MBKZtumqAky2wdW1V0D4/THWEZmhmG+sbZncDaHv49gbW6nmTVDwwhErHH5QLfp
/YVF0Ci0fMhT2XFAldSA82VVfx7GiS6tBYtY1YyQ9p+dzmM0FXUlv46FU6QGzkOK
9g2ZaoXIuI0tzHKg1yGpZoz6MUBECsPziOMsk7b62ZJFS7z2SxyPdUIZD1V8NogB
ijLyrrsHDS3xnJo4lEtkNjl2jGH5lE3AA4M/ujf87woI2OZYxYT2gkO7p3RyVseH
R2iG9/yKxfoB9TU/6z4zg/etWBZ1Qs1KQoy8T3OAst0HcmV5stWuPRrrE8TligBw
btZsUt4oWB+tQbTNcSF2RkOLe7WQw9wVynKEsY9LP9tOdztcvf85OhamyWw/A2uE
uypLTvm6vV8u53cN1beScbgmEN73oRotii+sU8Rrp5QR4FeijZmvM46XnASR39sC
VsqfYkAYnQ4dsU5rI1oQPlZ1jyxoS76zvenkUxV6YFFbAmD8WLeQf7qGKEoJGkbV
qo4mNQkLJUU71vBciH8p8kYBuKDhCIA9Yruf7Ci3gRFJmzSgQGIgVZF2Sq03zQB+
6vzNNYAFqbgpkjs/7ZFdXWfXHZ/GHro1Mk/Xe8urpJ4MGUciyDcEixr7kxbLd8sT
FxFaN54K9QFifAYxg8FccZJNgFIoXSkMyiVn7gNizy0HVT2hGYTFNF1XNUZQIv4R
ycfaGhWvJgTu2IsRigZNKyVeNIjYuwhix7giRNwLmK7H+vwxyYbFlFlg95yfi/is
MyEl9d1pB+augzT2LhA4gdKTX1p4IQ4VDwF2tK0Ck782RDLwjs6REt615ywWH0Hz
PnTHiOCiSoWcZBSwGW0e1K7+Pg7RwkOii9TtS9p6aFsy/JSrBfyHGrgpjCOSw4dV
SG0TM5YKNrWfpS/VlNcBlJkpzRr6ERu3AClrM5g5YvAzsoQ12q0dJjVKoUlTJSq1
yq0UXMbQIOvGlDOIeqxLV/yCa3AV/2k82tXQYeSSjJsOL5S/erYWmGG0tK2m6EuZ
dVoeaTzPFf4e4SXkw9/BTLbxEMXYu3lUr3Z0eQfxy+S74FIEGj3kmSE95qWXvI+8
BkLOEGIiiosGRJbQA6ZgZXyo2sRa3UV03SOhdWialfPVQCeJll8QYDUflkOitxrX
iKUFnt/UpLsCXqkuLPgk0szRPvfpalmLhKioxJasEEsgHShuYFTC+WkMqwtlwH3K
0c6w7lJeHfY1Txa76n5tg6Y7l87EO/WmOqj9RLFtbVkFi9lmccoeMNMVqbBMbVWP
kvrusIsrFT3F6LNnVXWw9SaSpdHFPpP3YihhtO2d6z3vhUq5APFDwml1Q4epSx1c
sgtqUzNJOTigjVxOtfuODp331PTCcWoxXfxhHIOIZY0WPhOCPl6/1BtYLQbO+8Ul
hKgqPvnGkZosiC9hP6hpj9XqQExEVIur4lRifsXnBLFTkwHo3rine0PFavE1gthO
+kbdwFA2Ns6j4mAHQyZSErMjl5Xz96JvpZoxGxtdj5eV9riQ0Mt1ajI+fbDhgCCV
L4K1PdYVokgvI+T1i5rTF6F4zGky0zq/SB1pT2jEpXCuZuJBYXwlcE6gFe5h3hf1
aI5GgXIHbJ6S4OfX2YVUQOja0JpvBKivNWOzEaifp8C+PdP0OP1mSJDrPa2K0bxm
gAEX6I3Uf6/+65R/hiSMoJXT6wliwYKk8zakVQsKOAYHSpGaHdlc4OFHqtHojTtI
fFx8rvSZ4wMZcZJUlSUWdRSR/ViLnbdb4LA4WGILk0o1Gw4iOleYaGoOxDvEDynZ
9FIcQ8qzqBaVXFyaG696l9oxXd2WAhpLEUqUt/nYQhMrht+oloU2vi+j3iM1LRRh
OOJEEZxVyJxT0wnhtE4R5eMX/v0PZEx9dM9ew2JWmFFdv1YdYMA+OuRMfxwEfYZL
kc2ZpD0WC4MglBdHr2vTuL9bymDs1V76I/QzV7hisW3hvvLoyw18+8ZP8Jcks8fL
VwSBtgfMx2ae0ALa+l6GsR8/rYD2J0suP3p0SwqzfVPush0I07TB+/TUJAo6Ix9G
6rc3RiDqMhY8sMTXFAuJwxBwlr2zjtrQ5cSk7Dw8KCHnbPlPFhQlCNp45KtXhvbm
Bxvifc1t+Gn9+JC/yLbix7b9qpEq9DWRmAoUC6gmZIGQMlKDLeGmL6MbrsiScP/n
QIfLjMTxlL4Aar5hbV8XAeauVJydkXqajAgwE4ceqs6VlIZYEHco+tOe78nFpTl+
i4q3VZjTybY74ZGtT4XAKDZmDm9iACpxPoEbRjV0HC7F7CcynzP7b4G1XKUfNL3X
d5nZ/gO1GMImNagDRJ2Sm8+ppVHzIPhJQ7DJ2drgyCDe/b1sqtvKX+WfGCOCELze
gQj86TT/uY7NbR2X3dISjwpuvFsrQNr/E/Ip7N5N86mZR4XOfmtf7obe2wIXepcd
x6AYArbkIGkZnqUwK7ANr0qFyxxuoVOf+zNz9ijI3PcUCfEc9cBTw4teWg+UNd3r
D2VbePaWOzZN0hTuifln58405ZEgVcom0aiRRgyXBey2PMX9mdQKodVlcfjoXMEV
xWYw9F+QYFsW1KLIoA4mknN89xAgPXSS6WcKiy9mK/fGrfPc2agJ8WaTJO1P9+g3
Xw+JWGBhptFscU7UIEwzMZoylUtq4L+vIKQn8xPN6eBULTm5j91AlL+eGzEWuqUf
0laYFBmd0nO2S5PHIqDmwZTqdGbAHzYthiZKdRSaJr0Sw2t7yOj5Z6GcShEmVTtU
CZcitqOLtLxh2oPgg/0uE9zZNxRpKwD6ICKA08Fz/k4j4BhRQTHxEeywuVqv5ocK
gmNZkSuJs0f+mbWx3y0ks/OV6RHpwcuywMVyJCKHruPTkvWsYLTkgJXlTI3KScyb
+5Y0hCqQy+6cV4r0dhFftyMX96dAgVGcg7QVQ38yZHvy5Bzesx3bIgpfl1rYcIqf
iQSYCCoReQj5duRskaudjYeW7pVTWRNyK5C9U9m0wm5nhI1z4fkmASw0tuTZYlh5
zZrbLHJ21veD4Xc3jHcPUwvzrm/UP40e34fq460hCZVEe91Q3TlKou7OHwmYAX5v
Sdhm22mQeXuUaO1VwZPsg4lS1gUbWyrOUAhhotWkyodMEsgXWojz0Wa7AB/03X9P
Sw7GiokHoCVTf+SeDDLlOmxm0gw/qzZveQJRcZjvQVxlXFyVU+RuP/U25qRXfonJ
+nRpwTTcA/NYmN9Qs38HyVgP6Dq2uAgGliS0dOFk09Pv7yXaQC/CRaO6nRukAsi2
AK27akEecdOl65yoLXY6kFUCjuAqegwljbdoiaOEIb/1F3oArTp/4QgMv2F9i7tk
LLpV4p/sbjXBMKhQEsrRIQddtGI0BkudeF/KrUxAiRVv78xISpV1P9W66x0+xMZD
4IWj19b1gNJ4Hrur2s+Hj8lEmzBqginQlGd8lAT1GjW5LmsPXwiIXRZK8ajFd6ci
XhKKYVIEupLQfVXMZFOFtpuG21OalObtJScFgCX/scjtD5/DOeGdDzbuX2Obe7VM
wvF3Csk4TmMMh333/0GDNqaKV4CEZ7bR4yCzhxtl830ldOp8v9rZui1i2p/TVdj4
8M/sFvpBnzeRpABbJTPHDzvFuOaaJcx3rbFaR0cVpE2KoE/GYN49GktBqtJwTAH5
+4ODf5tui6OknjNyK0Ua76S/+YjVsONB6tM2Ka159IdIg+C3Upx+cZ3mnbB/SV1u
QR6mPfAPn2EqHuV7F3hGp31rJd2QJq/ooiG6utgvEN6TXh66Q6mMoULh87MhQymi
eNsKEq8mCFwKEMvunBvK+dq++lCane/amJo9T0wz9a9+rfv8QCko+ZYYBynETlwC
7K7QSQKJNFFWl49YchnvzvwHy+NpVQxI2Jiz9ySeLzUJgKdhQrm+lb2ZaDmhYJ/Y
y8aJugDmdPPAAMuwQLOzbH4YAm0aPuOIsa6hJI518jbapmuli1s7ShAYj1VOY/Wi
1nYk+T1NE5NX/IrJaQM/M2SvmD7lTz7d8dvhOrKuqwhOLPykUvgA8MviwiZu2rnD
aIwmOilYMJq+mEzYfuXWCA38h7E9eJipA3gtSXvaxXuV6+f6mtTZkxJwFB9TF7G5
PR1r/0vYv1YBREwbH0Qcqzw2FY20bmezkgCnHAuAjpIyKEkzHh+h+1XKAFkjbygj
Qkc9awaU/uu7Y2g6G/6f/4DxK8kBkakvGTONZPp+nSLEirS8/ayYfgexi+DZg9pQ
8GvgMcwdgyA/Zn9DKaV/t//0oGR5aSfn3lIFw3b3hmDHbcX0kbakjyhCcVfGle5R
HpedV1vUrBjWHCvGdSn90G8GJK/Ny/ZK4iWFRuHB9h5N84GJ6PiIj6zvqNBWJYg0
sOKl931+WdIbkNZ3dToIy4PT4agXzlzomx6qlDDR29hdp9AH0k47UXH69UMGwRm0
S70Dj9gbChojq/yeuaYi6v1BCT9sO2P7Mq3mHDnd4Wy5jELex93b4POCH0zi31c0
G57Ftwk4hnJla71G50dtmjD5ipBHwt15yhASpCEBh1t0BJJL4o56EQ6Wc3ktmR0M
JRuHEfowO9oHUBjewX5Fu8gjHcFki84NX9jGxZIxyudQnB/0wqTzGRdHCjnGf482
VUJUMH4JYJMOhg4TdfpVECajonOWOQbo/CtxTSnFOLMlo596CiI+n7C7X0Dny5YN
Sl7l4EOPWmJK3EAQTeBMdhV8jnnAM2ziHKpC/Pomlv3L0Pz03bT2paIZQ8N7GSIp
nUlz7A5rYqaRmx13boxv9rPxJ3EnMWSaxETqrHcBT7m6ykJs7N2fOEvtg67SLC6G
jtAuQdsd0Ek0kSlnmIHmfZIk8Fcoko8DnHu6nk07vEodhp0fBYyLPIPekKDU6rD3
W1QbP82i6GFxgCS3LRWvgzI47rEXxoAxX/kVfNist/c2ZAStLmRYcfYVPQmsE2OU
dogcA0z66xaAkLaRG7wW3olOk+C/xUXxetEwVWFBVzenwJ4IJr4JdzuuV6Cr6LWl
6YivaXIPdfFiVHBA5egoowX1QoQfOpLgAzP9p8gTc5mlLBZD6sBR1xztyVfFkCaW
hZrpMTMMm5Ny0vmV37D5SKUdc+KKBwW7BUY2R0IgZWBvmzu7ednPTi9iAxe3KNaW
sVfGWE9aEiYclYBAlCTv5AVmrYs0Dib9pCfCkJ5oSl5TkXx3+rwaMGDmskasA0eQ
mdtoEIRL6vpevTcUYuDTgu8GPpRZHH9bi6OpaK7/oYDbY/otjshXSTNRJKk3KxFi
MgQxc3LCHidu7ace2m0S9Z24FZLKozRWDIhjH/U2fWqrGCgy3tqocd/cgYg251hI
3xvGcA/pJSfdcvLWrY4tasKwjmdd3L08hjNyCOiOo8XeRmHDOYEwF+58uUNkFACv
Ui+g/8wafCf0EZth/sHGuQ2wSdNXWB8yY9DiqoeC4mScqL0+n/8m8JD1qDPwXctt
tqaEbylVfb7FKh9dV9KfGoHWD+7eJ1LfjruBFCP8MTnwbSa1kS22OEnKSu3Mfazb
PPs2GnVBEauNqnDt4M4e13S261pDU2t6uSTOilXpQEvOuDAQpAqwqxeom1lcV3Ce
sl9qLSKgE38UyaVAMTC5HkPJxJO4lQq+d7CdQu6dLaMX1PCFFMneFGGoMTdeoxVi
L+j3hcZIXZG01tUS35U5Noh5tl9S+HEsMmmkl4Z3IH61ikhr68Ag5xMGuOmKTJ53
+cf2C+wIh76tj+eDsvvV8RxtifQSEB0q4FPIx2wr0URgOgBD02rQURd8H5wuK/O1
QgMsgbrtc/+J73RuzDPLb9St0XtR2Ttsxi4umEnWRnYr0rGsol7A19mCxQ0ZqvRS
TuCs94lezRvoIliv8xKgVebNJx/yrkEQ4y8E8AWAcBE1oDt+K9uUDw9IPV2cHH+9
duub0kNwgwY3nH61smhea/Eafb6Csq5g0FC7i0uw+Cbz74rVC95GQtNhAnTZJ5Lw
F5n14n4/PctCcDgnphaY5Y6s14tsBNOFguEfhvmUaRBzZ4JpyvYj7p8b2/TM8SFG
yMgs2/drBDBAPpJcXuOu+bHOK1AYaYe0FANPcdt0u0xGnbXkrJisET5BANye+/wj
pGWmtHkdHLUsnA8NYScqUoivifi+aBMc+xWF4hQqHFiX93GCx2j61lxZxC/kFYOy
jPcdLfB2pPFZR1bDxVYm9wQaepDWsVEcXHoMuQfgCJrdwQ/O5/VuYuKrVDCuRYm4
AkVDByiG2cwhVns4bCp1EnTlW8jBhDX6bAMljz91v4s7bWV2fZWUBviZ0HgT8QxM
FPfoBpie6aBjVpj3dsg0FAu1HYvaQrzkqMRmWJ/EE9c6AlxN4I2DFXHXkCy5qQ3p
5RdEn91CJfnFRTNOtnZx3VabqGU81Sxb0/YA8DomnsL9kMcwjpy5LBr/3csNTJS0
dmfEJdhuBw6rYiN01X+sLh6V01/Of6ZQPONrTHJKVHzQUm3UGfzbqoI5pWfEHNXG
yhFjnplQLnwBxlNv2Z/JnpgA77GNkWnHpWpkGVKVaTTxk7BUXT97hl0VkDf9n+fu
vtJVK+9prvNsFW/pYM6iaplIB6t5hK2hV2Dn9nO3swzJFHGrBOuLew4uUkTRlXXk
WzS9tfJV/wy6mgpAz9vh9mM4N3ScBHbNkj8r20Ap1/Vx19qRa9St0Ug2+4p8b68Y
SjjxTxm8PY0EApu0K4BhCBtPKO522ft7tlh17TpqESRIJ4gebgIp/T6TLLBXDXBo
f45WOxV5yN49Nqo9SkglmgrqRNtUeTjQxAXN9t+BhiGVzagUElfw4Skg/ZGfLXqM
Bj9iDpOCH/Q0ggvmnCBzpsA6i8Q1kcjKfqCmvUnwT1J234jpbDFalMHFbBKhn0Jx
JuOodARbAx1ncMpLXz7XwJCPxv6k+6VYSmB1LD8hwFDZlH06b/+EgY88+5+8pL09
m5QJr4vi9Fq3hseamfOTF45CoIgyUWtS9HEoPxpzzNIac7CYEWGmSbfNZ0dJ2MoU
8rnLxgFzbX8vjI3g2GqIJzl+VZ+hViJO57Xgh/hHPDQvtTxxUlMMZX1eJ1M2mJVI
Bygs0cSnt6V+PCdin2YLi6XEUqyyEF4oMrGdKzj7qC/Y2L1wBAnAHOlPtVx6tIsI
1INEw1MkZwb0BnmgFwc22n6WvkzKaF1jKfDuQdhfp9PTKtbT3IixJaWc0G5UhTd1
Fd5b0fXXMU6TmAc4WCV8dnlhTFQpQu0uMNBZL77G5782LdFg3fV0IPe3Dsfd8j7I
GbwWjWRL6AMmHLBCZQmc2+xA/Fc4RDm3FXshqRGUnp//91ShEokuxjo7Fd3ibWAB
f5WUxZU7xj20deQuXf85Y/AB1AK8bXd7tgT/nTS6JIa7d3sS7vSggzd8pdG5yCkd
lfUJc0vE9m0YE6+BjxB1TR3y1eN9Qf4zIHNEQlCI3Nu6V4MUtdliVR2NDvHqd6k2
htS7udUBGxy/+OjVraZIbNbPwFbUqE89+GqYD0VlJBtZzxIrxdcE1+o4l1xhefU7
5J4iTK9xdYW9ZsOs1Vv6MLTD813cSBRs83lFoC3957NKl5C0S7Be0Zt9zt6IflE4
2cHRpChKa/8pElXdDfkDBz1MnI++Pd1MAr/z74XD8cr1Xo8jMNofk7oKb8J/pLzu
8wUTid8DmSVejwH1bxa4wV29VhwbZBf0gGswYCQHQ80TZ2EYXh9dHszEdnEG7DGo
KK8OlYZISA8ZFBJ/nSbZm94k9PjiybWmjNnjV+01X1tKvhJahcRCiC8A2JJ/9ZM/
Apu1B9VVZGYdFeYMyZhy0I+IA+RSIz07RdXz6L4bzggk5fty9FN+iONpWJiOqbAG
Y0MEJcpJSykVz0SustGsYO7Ag0Rxwmgz4VmPAnBDLMDz+ta0giISGt6kl753AkHI
AwqaUdXF108QYmQvrHIkWg2z/M33zn6rYBu6xL51YvkwvigtgS6kHO/B4qJ/pYFP
lTOeMgcStJ6t1P5uEcnp9dwYJFyfzdXSj8F8rVayZ3iZppXiRPEbjarDVPNS9G2W
DsqgADVvo+fuMt0iWtmPuqtMu4KfywOi5aVZDKKIsWeUd1oG3z5p9flsvulOEkmn
hUM+lqwUZGBC9zLBGgCA9ym+eRbolpQdgajGMPZGFdWUNK6j2UJg8IQkrm0j/Oth
wrRivxunCTjPllQPFhU0qLoNClsfMGOzXP+zZoEBp7Cu4SFG4Jycir3O8xJWqVWI
BG+EhBKkGIAWGfIgVyGl6BU8Cz1lP1pPijRTzPPYeQHltjheg+H0UrwE+wg8hqGx
pqQ/wzd5DEOElwcz0msSiLtLb6Rxzp/U7kNzXyTX3tbPRKhwk7cPZXgi3FSkYgo8
hoUXZJt5336uVQisCzgWCOMkAUBOFaH9IgpkKQS2zJh6dOy2OvmmVDVvgiN5aFI3
n2DNIXVKesw9JT7zKyks3kaQS1x1sIQhYw3JwXrwzlYCTWJLr0lgvu2MaQpzxEJu
Ok6UlHUhLj5JnbUHOX7CHBaBBIp/GrXYw11FDmpI/tBCIa7UOEZl31+eR9weZIS6
3gNkQfUJ4lhKT9wxwIVMUuDLo+n3u6dsMBbV7jJTR6RIPYnzqG49sH/aIzefo/HQ
BNsy55vI4VW7m+3YRAHry4+XUm+f2KPKYyc9EUFtNJgKmMv4iUJurjz4wvuLqY1M
mAzWZIQzPXmU0VSIFcKXjRmGk+3lzRl5nzc6DBX3F51Zk6vvP4gflmS51lD3yR2L
5srg5KbRuqMO7Mnze5F20BikKRBdhITeKY1ncsnPFiTj9P5KjPK8z1+FD1BKPV0H
374AlgMKZr2E9Nl71e86xml7s8Txf/9BFydamvLjOYgZ1qiPVVqcUOpwK1fOiixH
Nvklwx08FUsFGU3ei21PXg1bh9kZyaogO/LXhS4R3b/NgrpB5LZFeXaMM3qf+gor
FY3x0qSsLiAP6bfzxLJVYk2qba8VhDfLRHGf4NPPz0xTtFJDTJKQSUxa/44k+epK
SHxfN6h0zpNpN3g6HUyM2RdsOfGoj71C1tk+66v1siuKKF6F6y+iMcURsFimYOcR
QGb23DeC4XQwTwVDeiv9TZ52yiN3VrFDg+ZQiRjsA0wcCdM3MCP7MqPJ45XYBpKj
NdBb0r/CrMsbC6rXawth4lxbPReTsOYzDftO9S9/T+OEFz2MYCYaDpuGbSjq2A3X
j1KTWireEd2Qf2cs/G6EUCkR2znC9SWlJu+7bjH0KTJzz7wZlWAH9y7czOsutKwN
OFSvhhKudp9nTarXE4zCsgsi2R12rXuY8Yg5Lw7zaEbwpwKSv7nAXc0Ql7ipPsGt
evAcShbFRcjLOKGwvj/YiBALskEHJGMCpSGrqBAJQX90MkPCAOA7FS7rt8wPgXlf
rUi8h+wjkMCt9oI/PkWkuIETg9CWQcSoVZE5AyY1jHaj03QmC33fzM4mpWfloAs5
hWVZelU16NUGyuHbz85L4Mq8NqLfSlCXF+DDlcTNHozdWzU1yrr9356Xo/x26A0V
ShyNXOBoxrOpaP1IKQQoiDRjYaGu+Bd7EymjgJgVmpfCQ9dBSFHRf2UMU0bUEkpf
4999U+zmvJkX4RM/e7OT+NpA81bia9P84aRWyRHz/Wgkc1ehOKzjHQx+OXHKyMya
G578aQWeo4ZaMmBOj7aVeKeSz9EjiPkBIzkgiwTyYbgfIdwfyf2iHmfzbFvmMppj
JwLT2v1o4cnj3MG7f5pVib0OFYenxs367UiMb6MoccRs2PtrU+GW9Gx0wQ9sIEln
4O487CsTUuZmq2zV+OL7oZEQq7GvoUNMFaQ/MNHTpH5W3HZBqH5X0j1jAWK/9pwu
EvlULUc2aeUgS5bdoyRUrlRkqZyFpWe9vLOi+xmL4dlpK8U8BrStVHFzhywyKeHt
uVMfTnBmQfYWDY3V5gilfBgShgcvEm+Z71t7MnTzYx4afrRO1tqMVjUGA3KdXXZU
cCoGVLtPsAmAIRbFU9EsU+zQBZ9PpM+scybxWVfM9RuXTt3CgLpkkon4m6Jt6VMn
JRh28vACbEBZCuk+I2yeHyBH8fMVbQE6C/l+gta7fQ7tFZbPg2+hGCMe8jXn3v/6
cRMd5WbViJZ3+Kx/YDe8OSlX6QKOphD6iu9uW9EZ2gPM2s/cXQcMTH6037+kYlOW
UFW0Kh0ACDPDX9EpyqM8GjDaHBVe8JOmejiytHbW/U4JtmbNJ5xWriDlIoXaG/7R
k4a8iojY9cxKpniFPXQdU0Ob7ZeqoYg70MfTktgZq2vBm72vKsRor605wOn+6W90
cqQkbZcaovRYLi5QCFrNvH0B3Ywk+lVIJKw9hoIBxlnKgUAltqxMjhyaex05eP9J
qB1+iLUfe4ZCrHi2be69bjd6THDOBYrO56gcBEY/uVXVLfcUUjFqe3e+L5toTypj
QlrhxxWdbNsGV35WEdPC48UFLv4hwlpZDgTlJg8u2AZLqUhZK2+yowNYw7MrdLpe
6AdUV09wXu1FgZ95BKMFAheVFonNvO2lLcTaT9svBrXgIfuu924GUbiRB9bymQ9w
pdfKINTjB2TOstEkaxxKHwgwT/be86d/4D48TaFggQYF/g+a6GjPOwKTFISWI1VZ
36ha3gwSp9xNo4/IG8G7Lm+6qRI7+tvie8qSCp9hT660FOAmNlzKF7GACiZSgHxi
LdqFmV9Iedp+YwzPK12PbS26CBy1kjpoxaEunYXfcyN2KPCsSX+VNLl4wrDvnBac
irnZnVQ5kHM2S5pa5/SbCZRnm5iSBH/3J6RduYOD/dE78BElmnmJx7Ka3+ErKYiw
9g27UgDP+FjSyCxsnXS/uPwXvJSWgnhhn/+FZ/zyFojuYD/kW/tk+goxYtPKFQlP
tlW3oLBzeacmBMl8F5abRC52rWvXA74pBwYXKtoyPFp49LtiDTJlzNXeG6YBHm/M
K5xOw8eM5JwomPGwgsWpglgXeXdyHycm3zJg6ywj22Djrk1oBVj2Mjxhh10T7+0b
4VylWO8vYsYR5RcyGmprOpgbgsi3uGSn75Res/5xIKCPfZWO6cPKRCHjUKSCtzaV
w8FCUc+C19NMjgXLymlsWw2dZWH4OoEzDNZqtX9khdS3yP8u4p77AF7WMe5LzyDx
+MoaQfAQvdxxZ4CG9Fpc4dvNmR5jg1b7HZ+d3TIlmHtoFWZpjxK40z/vtIEfvn5z
yViXySwaifR43+DWqmLEFxNny2L9lrpAmO5vJvWNApV83msgN1Y5gYZHJ2+IxrOO
j3G7VPIKjZv3Irgmn0N9D3y7C1eKeKvCVkbcI0fqSbO+R332krJS5Gfhv4u/S9lm
dTV7/fw4ImScn6C/xqtTO1ARbqrpQQWfxyHTFfh6jV09YfUxzyV5BV3WfeBwQISu
49ia3ujowKR/gEFjwFcpD1CMAi8OZwsMxVOu6zbt1lXft1RNAGK+b21gUZWjt+uR
GqO7zxWXrGfCamggd/fp/6fkk6Pv5fsGtYRfpNHJl5YVLLRmyPlcEuqT/krYgRxG
ltv3AOKH72BOhKje0aM3iWDvCGSlxS3JVu8jrB0Yl7cBalOAdtXujiuvn9RGke0o
SFjchnERAwxssmnC0GXWXFICkZMB70YZPwVtzKN77gNnPpixL+1AtIK2XIbzdM32
5XzGW/3sgrrECW561v0Qbgv9J0gy+OHdWx0F060gL70/LmxH9umiRB016K9FpM3D
yKrlzzx0WR0PpyclF50lIlizCibdCB3W6RoQ6W9VCrucPzoNKtnBz+T2L+QCsTfJ
9fstTP3qDZkWMK8Cu3pgm41P5Y9V7dpLGvGK3VgMgb3NH7noMyiXc4l3wSC38sDA
E+zUCtXPd3pteCj1uCanvSOUJ8fCVkoFMTpS/u/5l2RjCIDoY2A2bCJK9ATfOesp
6bB36T3QQWFTIAZX/FeNvTQOIDyWaiW+HzevN7kG97cJ+2qY/jhR+a3ek4LN3az5
YQKifeSz6gRTC1edD7IicNZqh/wMeCrtqj2OAiYx+1ek7xjDONVwk6CCG2LsJfCe
gVg3vbl1hiSGPFnQTEsZaEQsi4zUBoUfe22xMRoFsXycZswvOs6z4RdN1z4Mk9z+
xdjKax+lsr4z8wuSu4TKwnF3bajwKTr9LXC4VY+taAYr1w03keVzBtOnQveW3KlZ
IFS1yNag8A55f1kKedYj1mGkp30SBefkg0D2Ug2B21WalHpsTaqkX0fF283JN+8H
SoZB78daD5Otst6R3STJUjkcfJ177qBu1EaKcZhDMJfO60Db1yH30PtFNyLIB6Jk
2jn9LS+3eb/xcLzjTKtFbY8Ndx7h8nsyx8QtotG48YDrX1/tiyqOhiuT4ncGDexj
JgmmV1Uzakb5dhMznD0QDTbj16v+an7Nbx833q9Elg0P5NhXFW67TTXm7aFdnrwF
YeFAmguUlk4c3oUZXgiuj0iM7hRaBl5JZnHvnK63Q9whp4iE3h2B+LFien6e8Ptf
jFgxIZkMZ3+G+CLS/gVu4q6X0Eb1ACkHIEVDBuLBE+KWdFGwk0EJX8o7RRF4wvRf
GzRpyUlNOCi9mqJKn2V5RmuFbtS5f5UvqZGBKpHjbb46Flc0Gpts/VccAUfgl1GA
usL2WdxspzXtY2hoJHaYlZf+DmLyq849qIE0I+3BZ1t6npM7i2wJ6TTmZHOJv1gG
97QPDQAfVgT0U8RPqxqOglHqKoDH8OKdfxbn9nsKOkByLYKDYTRDGM1VMWaXwH2k
QnwDOPE4xpGnyE+O2yb9nD9ztI6fJhri8M8BpzzuWrfqarJPY5NeApGXuKJTquFy
l7vjy19IqEH3rI9lLUFr7sJB1D9i3g9qtbbiKDtb85yW+ZmAA3KvjGBxKTAWEPHu
IIFXDEBwBdtSc/Yo2V840UPgl5enbshwzgBueuf4c5PbUoLrv58bP9xCCzjx7YCm
OH0HTKazrknhbWOOQfYVgw2kP+7cIClVDGzLpnOgY1yuXeCKu7O8QQWO8dMQQHG/
ko59FwrhQjpXGO8Xd0HcdkrX8vfGgwhXpYNZb0pOEbg+99c8bSBuxr11KXxMXSwE
QCdBgaT4wrdK5U5IGYpBYau1N1GI8ZIloXZ0SmSsqdmGt5XCu9MjCuATSBqTzg5B
C+IxZNuEF1qkZrkXrBaaqNA0scjNKitDpGduC/D1EyutE3btpeXg4uX4GxWxFPB2
+xc16fdLZNlMqequN5X/ABjT1ifVU7ek5dYPjKctPYmfDlB4zJUeSmePOx0jOjZt
vh8RziWGco1JPimWEYyFdvaEqqJ2CAcVm/yOu0oxOhmAWwYAem9UfgZVQbdqN83D
QRQT6ysEHOT9HwT+bE77VkB9cNS/HVwPkZtdu7+VAP9Ku4YPkwpLrr/8jeOzu//z
m9639WvmiXjTXsckw+q/hk5d2svpNhIp7TzXC9DvbcnoSw8kEqAfV9Uq6WHP+uNd
Ctlbar0b5o+yueX6LlVScz4yZchFB7dqG+eoVUKW/NnYgNW5nEwhJ2qK4tDAPDAf
iNiibVVIxGiXRUuOncD1r5/di5QeMlCQtEt5JPuE86bil6oq2MtiebivLY+Xw04B
D9xPvlTz9quAYi8Ihqur14jdIz47OCFaClBbnegEGXOgBkWE4NRF4qD2bYz2n8j8
k0LUT7w9gpJb9jQzOPCzKZusi9O3QDhYaR+r7Y3A/AqPqY2b7n7PpFCEX1sdfa1o
1TioKb19wzGasqoYbqrBqpJDTDYA08nYVbX3/gkF+XBIyzou8D4iEUJ4cRj49m+v
KK1d/Zw07RayXE5W+vhbTWYUZA8HuTP/R3N5dl4522pSaUE+JWGjlskNOuqRtSCy
qkgkQv0p1Nkkrsev6kcVRhNdTK8qyYcsMSKc0W/rQMd126xE290qdxM0DnyT1ade
e8XrqEhmVfrOgDsJePHJE//rkTKcaf+kGpkBLnYWUfX8fX+ln+4YwO5dN3X+E4u7
xr65apfoHwWJBK+WBqORDGEKz43U367deZmr7SJ+jOTZ8eGYDe2beqn9YWTOEIlP
slGkps48zn2unpTBdh3v0SQzrxUJ8Sb99HdWmY8fokt7WygX1FlcuML2mACzIfyr
a1yYny2uobCNK2r0EExCrDMX3cfD8tvctWcKSTPc/pVZ7mw0Im548KdGeUMzDq75
3LL37IRJx/aJS0WuK5Qpq5vc1MRzwt2qCk5hjEHPluFv3QhARhybkQakHFbkSqNA
jx1yLg+OG7frttmKoUmjD36517zC3rIwu1ZD7Ny/AHM2HWzOAAVyqRAofGlBWJlx
9O7RdtG4rgOyoc6K5hNiOBDPchxhSY+cK815xVjmhNmi58yGSm7P0kHvtjdEKOXj
ekeBzarEwbkcCFjM3h2tRMIAlsuu4xiDRzmvwxCLnllTBK+exQA+/m6Ym+mclrrd
EqDcaInKnAeCiDzL3xyvxmPO1hyUu9TKolrFp/r1F38esMdzeqMVzG0ZyM6FWpBE
CQSo1niKJVt72WD4a/QGAde2tyII14d8k2Bp/B7vN1QNSjNdtJR6N/6Z5Cu9MIV1
VAQL+J3BXrut0h9X2tsHx2EJpZrS7O7enbz46cpMLlX/hw5LrB3S0aDacy2mL+4F
viW6Z8flT52a2i+8GxjGmHzfhGorg02VFJGuCxHWdLS8Gi3VvrKjpbHl2FwdeHl2
pZvwWHpqGviM21+G4GgbVrAFToc/37SWfeslbwqKPg4ixtrHCr+Eg9uiaNflik/9
ud3qZhcWXuDKH/WSTjsnjgS69T5Gnra/k3KfB17jdJRx8caUeBFbkR+IObdfyqKI
ZaiJIU4+IuccKLTAJzXYrnbFwXqDFkRNnWYrMFioZwS7colUOjXHqve1PFEOQ3L3
9PDHZhQ4DU7CcXnEICTwNpMfRe42xqzEk6UKal9vtcFa+1umyqhCdeYWSlG4b1X+
yA63ozSNu3bl2StYOMmvVUUgpcAszIIK6fMMe/7txET6TdEyL6fL/xZsQk2rz1/+
yOKDcyGzm9YQntD8QbbvWXd5O0Ac5pjgbG+8FMagMse0Vsa1Bv0O8Tjm/BjeJgtj
XMjgXVyTXzCSKZ6oIhem79Ayaf5feGrVdDNMTHi9ZG4K98NsDrQuyMsRbWImdL6G
luu+4kTErF4fNsR7zusOmRNHXcouxIxc1Rb2VForGwvblbhcMkWImfjtTb8gCaj5
1UV65G6TQi14CjW7wil3bJJNhQwWzvgZI4SsGuP235xI2U6jY3nmZTfcuXItwi+y
bSpypY0+cTiBDpGC1KNYPHKE4AZzutMpmZpHiTeIvZ+hr/zXCLPTuXd/U8xaNh4P
NQhF3GG72xvRD6OimAw6NxnGEMi37N7MnS3Davy60leUdzo7DgQrQLqBklYf6Rcn
+m215nGyiBKN/L4glMYlq2N2jTx2xp0H2DUXk5SKxxLkoBlDpfFenpDFND/Rksqi
vTPpE19jI0CONJkNer1oiLRamQWi0jA5qbd/SqFnokeOaMPps12ligpRLZQ5bNhR
aSChLVA01qZ6qcVRFrWLwH8+yR2QMNSBtCLAtFyV3ZA6ZFm49q4c0ug+5vxavq4u
xZdINN2ErPygS11qtUMD2C8Sr9rZtBwVTLLDrKWPmtxYeqNhVE3v9vT3AndOUhFH
Isn3putFP+XZ9q/+/s2jLIHHNbH02Rq+8W6yO0Rlwcj9sMP0aQjLgsXEFrGmABPp
BvK86yM9/tdwuDSDPH7KaAAblDetHBeNYF1jDixOf/o+6nfK3lx8Z1S2SmXN4wNL
ujce9XPj2OA9/DwtkpNaX8dA1gDMLhyR4ViL9ZrE1v8j0nSFJffxsErL0FDwsFVs
P8zEyJ4IH/2VpX126O1IZliYsLhmYZKrNTq8vT3ry5vS71qQ0IzQu0p6t5p3EKl+
n4zK2wSfKlOpzfUVvNx/JPUsVznfgXsSiScuL/cOc+xnXl3ADTVjleCx3mEir1bp
vgMiGkXLK+sJ2tYp/zzVkvDCCjfbxOqjXEASggoI355M8Le8/HrtDg11gu6f/rRG
ivEp+y9ybp4iI3iRAg19pmqtVKe8Ybv8nMXPOFeGX6ovvG6/YicXcO8q1j+ZvVNJ
e0df+ohpFp+tqtkaUCZMM43WZCFB7uI2yMnGOGBU0YDl4c43IgypCA1DRj0R0bQ5
DuhnXupImUSMCcsQ+sxmOCHa4xP+2uXvzqo0ju2bFEja5AId+wiwsSddsxPDePqs
Q47D4siTjr6zSrbCkl2eGlY+kmDDUmmk/pFzX7yWHXWkhbXQECRByfGRawJTEjnl
0XVe/Aps3HnjgqS6F9TpFzsV/MDXbLuKUiDDIcQu0qnt0CsqKUAQk9P7Ff6VTYMH
ZKZ8IubxtsrbDm0BxxuKnZK/V50jzbMcRoQPDH/BusZj4lU1uRNznh/+pWxuGCRl
lPxD37iN6yFdmRS5+l/v6hUncxLakxA7o8s8gXPo4pRbULdoAvTZsYv53cQFBnMA
JvFYMvWzzAwhHnrnEIInUn6sqGr2SwY1OqKym0nYZKK7hlb1GU1uc73Lx9WbEjBT
wjKzfgOKsMCWX3LXYymVvtsZ0HIp0FOqEXBEfhsjvh8EJ7T7vErq/ykzFmiKzPaa
SJIntIBhJswrbFDjkowaO1UgnCXVzpmSsIEw81LpVLKWmeXVI6HPb97VsdkeiL+K
ayL5FMZYU5hi38TZTf8Pc4OKXVzLxkIFrMIYQyLhi9+CWN/LX+u7EkfSSmgraats
hjwSCjd29Z4kwe317sZPJJqHDuBuzQ5tsLFlmQgKJs+o6uBemEf4q51eIDiUCCqO
g65+V/sYHBGdo+EXZ11DLrj1LEX/ITm+vlLi4MZKTnxXfSJSXlk5ditaJHpS1ahn
mWLf2f6BuePnao0JchB7KfIHy/VjN75i2eeDOGz0avLwhQqnJqywEq/3ELuJpE0X
XPKdeoJap8rURaiZqUfvjBiVJ21y+vUsBcn6BxjNItzy54oaeagF2ISmls3uMX5U
XRKmmBy2nDjdaQu74xVmFPSizX08goDjZhTbJUR6GxCPGvbbXG19elfTqd8cFI5Y
+hh7KSTr7h9djxdF9dAKVl9iNIEUM7zJoK21xgMHunfHKA8GhiNVC/+vsRo6wpzB
Tz9nNIvZCrrT2vVlb1keal1THKk+uQWYaqVAtHVCl0GzAgWzivkWSo+LDZKha8Ds
4lfSnaV1LGStDEvHvXgYEgboRF+/Uu5TvY4/0JalYlzGacIE4GUvHy/wfr3g87XG
ctv0blNg905ClpwYbCRRxf+Z9wOKagjSz3kl3tVzH7DRKYm0YlK0JYcLlAQdGRM7
42/z+MEXPXikUU9uwT5yM54EYPEd+Fg100rNSZaTl1xdIcUhr4QAgfImpRH9HNgY
6GDBBXy7mgL2BJJFXAs41aOJ8mWk86o+mBRHM2BPxJ6twqBqen3DrozTZtFAVEt+
ztkbe41VtKtW8akZgQ05elD20feCyuZNbJlLTm2k1YRWxxssS+XvmzdQeNBEtdo6
ZEg0Rv2M0ez9a2ou/+gtWyZZ/o51H/xzFwIi++v0P9lmEEQbl09pGO8o2yayVQOd
u13JZFBcVZfpLi9uHocL96i47iKz9H9He7AFjWytIk3+/B+jZVMMRGyxcQhzHPmT
rl75rvemmWrALhVO3L7SW5vFLQxAPg+fqJSXWspP/yQiQPhPSHzp9FngsOe5djje
8fS8dWPA+HOQ5Vik6VxOyoMyKUVv3XrT1B1trz0LXkaHQAa584O4DjakD1SxcKRk
zpSytcYv/WnPfPXtsP7u4b9YW3L3EQ0+PiHGuDjhvo8iiKMHcK49PjMrS2Cqdj/X
WYLyEL9QjSylajoQOneBW4nUt+A/AFoGKlPWsn+95XW+W78SPFUrjMbGgTV+KtLF
opqeEpuRL24yht1vjh7jAz7wluhoXHCkMLq3qgledA4sRc0cEekT6vEIGLhr/JxL
k3Hz4Kn05EBEk0w/GJoHhMlvOzBnGH3wUNr7ExZuv2NgrlTvqCEo7b9P9OGJjPu7
LyPcdsjFye2CVxWfm80xef6i2taorQqcbTsbwr6SG2ePf4P4eJzSoF3U/Wb80hOs
dQPDmr0KHQBeH1K4rpKWVHjqnWWZdIg+e9XJ1svl29eJi1pP3dBo99LglN9H1l1g
8wAF8kvndRhszBT+BwoVEDTGP0wtOvDHt09lvlsd1T5v47wuaRiXP2Gp3AaBMjml
qBKl6/FOIZPmrmEFPo8iAts+/axCVk85MShUxP7rBwiA8/ALTzlJWAKUYMu9DoPW
tQE0Dzie9EdujrUddNiPKsCoq7wqo9J8Gctc2Ou2VI07NWD2VLohJnlFVKO3RsBk
cZE93FeV2/+Ysxkk1YyYRQm2evlAi/3SwwQhIyXydOuOe5n9GlUhy4F8r7n+MIlA
P6qf59bKR+1eHe14DkoODe5W+X1DeYm5MT6Pnbvl59hlJXEONZsndF6V5mN/Wk/c
FyhOkKx7PuldMt6WpjcvNN6JWc6C0c3BF2E3pRz1K/Hm3nlI1iunLamcEfFW5O6b
rS45ZXj7OJIsMcu4npayt//s22l+JUSAQ/Eq9gylWVqZ2ORT7ruSgkzN4RPczVwe
L7IkgRDqTL5sIulaWit6JOlKIwTaxZqZEdbbrsC+HggaXcu3R59Bwv7g4sAto/2U
j7WJDeGumouZhufP3s7rIsF9vKJ5ndH+IgPq6FiVXpKLmGaly5qwtWZVkf8JQdF9
iBsC7j5xTWyrelq8ap13962mKb4e3GDSBsnEDQwr1VQ7V4WIQpDgcQIIycEeIte9
LLNhEH4KvEJRx9qx0EiW+6nmfPp39jGUSzlvjBWxwSsSGEPDuXFHOkgr7RIwW/lu
6UTHBaRGwf+cIuyhr364ZLTy5HlItAadRxZ6TqiB2g435pEuHY6zJsS5fiPlfb4C
wtAYVzEOJ1+T4V9wTnPkRsKJeQeU6bNDpGnG8CrbcDR/T5o3S6ykKgXKubEI6aYP
wQLXYPlu5CeGbdyLPFN8xonfvujEM0TKohES7bNotCOUWKtV+G1gjYS86z0HXdY0
f0OPmIAwxgPc8XcQuB69X+gyE+s5tGv3fY/B16uaQW7FfjrOHzozeXoKjUdeHnSN
eAZ7D03hrIPk9D7f4BGxTIi5FrgwnzJlOKzp2KBnYXWd8maGipndb+6L4uj/UAW6
2PmOMqidnMeavNPX5JjD5A12Mu/nxC8WPe1eoj+nIw8PT/TL68AXgco5MreBgb7R
4nz+29EDP2ku4uigGRr1AN7Ot+0hq2COBe1b+Vxpp947N20/w22bP/9uKNAu0FeZ
9M7FR+48uGG/HeonGdVYV6nnlWyVbEUQPQborf6l7KUkVqvns1jKM3gnqyMz1hSQ
rZWQgXUun/HvebTtaT6MmzYbdzksGvJcRXnm4Ez61KegfB2xLJ2jLY7VQVTecbb5
OzoKtdNnCwahqjac6TTQvShpE2uLNcWxeqiF/xsvHMTHUuaA8RWava042yzzk0nB
d1IAUyvekm93sfGehocllz9RHvfj6j93X7S9zi0XoLsquywCcO++HA/4/sPIXv4p
jYQcV9zYR96sAPYqX679Nzce5Up7EieyAqgcfRWTSR+kaOUSsgvrwQlszJpgzhMf
5oCmpzgdscCPTfTExIJHWPBpEZzSntTzRvyAsQv5xw9idF+giDTVbrFWH1u9ZqNH
xamfPNF5FbMCztsaaJ63CWXir5UFJb5LvirBoeIPoMGLsBEWmCqBxbBqxczpaxYM
c6R99/ZBnPAOFh5fUJzPzlLVt8xR1/wR3FFPmmojmuNgVHajCNDrZJRPxSp0vlG5
PBq5ECtclBpIKfKHAEB5gtN9KGvFcoJe7iQikww2MnDTisVu5W0jgBKoCYLRmN+s
OESaIZ3EPzSx5BY63q7SRJJsHt1iaG2h0fFvRwWSpdvAiaISPr3WzyD1bf+3Li2O
DNmp3z7dR2ypF0g6Mxa7woeo/8UglocNx8Sm4TAyJ29ajZN3b9zaESR12i3/6+qW
agR+nMb+/C9tfYEoBdzDBGoJHJ7Ii4Fo0doqOVMNmMVprOsdu9hCGiI8coRB+8hj
wkGhjj3xvNut7wFX6W8Gb4wHE5Mlxh0zQpt07Ll2F9o3e7iXnNVrbInPLPw4gT7R
3B+Pzj7s5PJhYDmIsLG6Zqf2Pv7m/oUAEzMwaMe7jFYnb4xY3JxrtKUfF02bc0bF
gEzWxrvgksq43vKOACZBHI+Vs5jBfL4UW2mvsK/WSSZfKcjDr1cN9nbMOcZ7U9f6
VH0eZVG+56jYuMsSZz4nbLHNdW27YfwNBKxHz2ED12DZmpG/Xxjer0jdjdbIVw13
KEJ9VcsBVrl8m0JOYoPar6VuJc9Fn+W35K3yGy1Re4LSmSBXSl5/XONTE6nPyEX5
5+y3ySYGP6NHCHcKu1JvDJ/dBMCW8Zkg3P9hsWp0PpQtO3VVkjsE+h8imceovq4I
HeSnt5xdC5XlN4FJO1vaUF3xThv7uNpMENiXkDd+i44qPAuDIqtLzipo1BG72vq/
TXSJAIgMhPuh+nP+5bobNuwDitXgznKhqS2C+w15mwGKxvxvcTSQ5Myym3H/Eg4f
U9IaUkED6cWWMz297oRi7hwluIp/hkA3TWSkdxuDV79J+eGazs6F+kWtxDmjtW9d
ZH5tCetMtfNmdE0n7Au2/BLOalvlf4w4BI1JWYL0qBpUBpx32uwp7h5py2FGsp7j
G79RFH1p1GmRrCSeQd/SuYBqb23tfTxOhTn6ftvuf76cU3ONWp9ui25vIKPMv0rC
gpxFKGcw9YEmwoEea7k4C9XddLastwaFb874aIJ2ZK3fU5l6GFSmBsZQIW5MJN5A
MXorMIRZv7J7jxUj+ujAuUqKA4qpxgbG7dupIT70G8l1nhYbxIae4fVYf/uO0ZTq
z5RIqXUPqHB4KMITzqbrJd44V3x9VMNUEbMKGiiiYl6JkmUZ0v94oedDPDbRDou9
T9F64vBgyNLk+8fcaMWHCQN0T2CWJ+gU+EqJER1x4NWso67q+2qgBpWuIsKzvd+C
GuoWu1kqNf4OBU06QrHQ3OaQJUWrTuTpGQki1STWy7k/V6WjkY+mIm1bIfdHyaRu
t943+Y0urJN1/wIr/cVSDmhtE7N2/7fS7e6puH7u/eBU00F8CX8Q6s6Fs4F3H2rV
5SzlBlfFv5iDhtoAk3C2INe2BJ9707+NS78Fbhm1rR3q0PkZZC9/LdB6ysGjFY73
N3nCbD1dCCT91LUlt9oLIMAevDVadN6Xx7FG26WCmFQO4XIXLALgMHoTvOnOiVxF
DBl7Yb7/gOYY2HDrAA0bBrIo6SAwNw3q5PKxYDq5b1TqOb5PDHUf7foeK2DraTRu
MaJOf9xMAGbH/wK8TvHxrn+lcpb6FPHc2kJQe5Bv6Jp1UKu5kHOgmKeFpg+fKUrH
UJs36jRQMhOnxWD24gqDT78psSSogXRhnukSSSCWKeIExUqJZN5SsU1yNFojPHbo
b0ieDWnNPYvZJeVENEdePCmmkqMrdSC0kg25is8o1OA2M109lDaAcA/5W3JjE/Fr
Dd9YtVRrUnr8qzOvLu4fUJ06cr2A2f+dGoMfMEoaBD/e4TRVdHa5jjnC8jsUtBOS
KQIOy32JzLlalzaeRFjIx3T8lBLhIlo4nUDRAEiRSuD78Vi4cP6WT0TL+fZqsabo
ZtfVGpgZEjcZbvP5tC7+3NFw5aWzjO7j5YYijSGWApO6p/7rVr7jGyzQjuxCaql/
Qv+WtLqTP1foynkN9+QaSTQEv9+3UHVmBmnW9iO7lOw67KS9mreHjUBBl6B+TssM
Bu5tUrMACR9hWHBwlKmImYUSHLhf6TQmlcCWjKXEisZADvpbvKUVQzodzq+LR1lc
B6eLOIIIIzFb3d/UmM3mfPr8ILKzUC8vmp3jqto0NgH26F5lfMbKlodsIzjvYjAW
9KubvulkhW7qt8AW1ylM7DiDT5m6WRopoWbrgDH+u0++8RisounV8hilwHnb9BPQ
kS/4ByN6UYLni6N2hvHjGY3ojxgRDj+8L5bRgtEfGsXVC5pcvc6w+B5DK81in8a8
M4BBpx+6UEMR41xHqyqqkBLTbqfhqPwD6/PjIEULzBGkW7hbKDnHNyp8Dwjrgn1V
zewcNYza01lm/gF2td+8EnplDT/IF64DMk4yCz5gFPCTx80pj9ZKWLAE1Yt50vBQ
xhzI1NQIdhUfMFvgYQJgnpvEHd52AC/fM562F8lsaJwHuIPduV9SB3FPtb56hxw4
28nHVwYgEZbLa7le12bJoN3qaoyNZ2k3HoUZ4pYehUAWVB7IS6AwUZM63tgtTJVo
G6XcQD9gRGJsfxFhRiTIX8VZyRY11ea3kgvhMr0/IREXrhjvTWUUExuyDNP41wuD
H0pJfmaN4hZKyu0md8Fxqv/87gd6HowkEhTi/ut1AajByuRiNwGMy+KvWmxV5tzf
L14sgOQ/5ExPypYj4ZcptxAnxkmmCGEJBoXGxMucQjBkubQBzDkXntop9obT8ooq
H9fqcJXscCzaRdnASdH8XDwjItDUzxzYGPCdTFREeBbj1hPVwC/oOZRjBckkOMQQ
MiY9p/skY/jBrLkSOGspMTGJsnhYfYaEMgIo4a9bRqLit8WG6tLr54Fy5eWyrStC
cjvNJJNldCOxPyN/D/hob5XBnCh7llE+rrWl+FayYhd772yVvRqDldYj2iSVdjpT
pmFlCa0mhkxj3nDW9iG/9W+Ffs+JygnU9x7Dpwxos+h9qTBA4TC354JGe3P/hjoK
DxUPs+8wIR1JRlUI3YTE2ABRK680TKcxVCne7vToLTpEqhK0TMYcdQgSRkQ6i8O8
+Gh5Q4cuI6bA1yNnkW4Wfy2VlsmW2u01c5c8YdR7oMethKm5So+Yqjkpb+mRj0lm
zsoklpVzpzw29hAtYk2YWHCXxJaH+b/xnujCCFr4/VkJzlu5BO82CKdCbqOlyoCK
LxWCNoVGE4TfHXugYdXA/4JyFmis/dJ/RxeZwvs1S8LoAeF5XUlirDkImgpzmd7h
hIN1XaxFL4P7nZOrFHsM2XXrIsoH31esQc/eP17TwCIbZKR1n+KbRCEK86Yeo3AO
lmjCLdEq5iiTRO2sqg57S8mv0CN85KsiLm3Ja3E4YQk/MoPEDEpqMwX0zdhGcgfQ
xorAAgu9bcNXmHnpQnwlLHa3F75DAQfBrdTUrn97Mt6OffN3bFExiihewlhVxfX0
21o5Zgblhhax7XM8hdi2z3ogtCCoe2SN5yaJJcVmDIcNCmy8GksZSDCOVgIE1XEt
tJGnYAhTcF82Z/S3P/z5KdVROEdTxhVsenlDz3b7OJBj77W3k7hnPtVyRnloCWqt
yt4pfVj0ouJeIBURsmCL5mxQghG7y9tL5O4ta4KyHJ15SY3l1CHouxS8SuLkw1t6
hI+4pgpnBFE86Sqz1rgXgnshYnT5FGOsKk437ID0HYqihd9+sSdXVwJS5D/gyfDd
3CSd5nIGWmGawMcGLWxy5ePcMqtKxlqY874Nlso1UkQEDIwhXl/q0lLGH3rg5LVZ
Gk8KyK/Kii38zjJGlB/N+/KYqfaf522gyQd7Z0Qqj7H5ZPyIcr/UpyjYak5T+Ymm
UZhGiuIqOT65n5F4Xnyaxbe9fDW8nyif9Ricn2zjWeuES51UDMZNts3mCcBgajrg
x/UNi8aLGXkFl3n7ONsTJQdVOH36iWFMXRHYPVe5uObuqfI5BvnYYg0WilqKSgzS
BW9AFpWDr1Ufs662XG1cC2UB/g4uVmd9q+e5+fGR67UP0oPnHhUl3XGpml+rJu9X
vQ9H8ycLqyIGQXVoJz1ARGi3aLJE5Wut4zFYN1XipQn6QMb+aHKiMEYgYD3gbdS/
QI9d4pvJ+FJG/e2kNFBGq/RwY22y8IdnBSAWYxW48+qNFoW/ccqIoMDKTIBFY0N7
DKlR1uIWR0fYg71DvJ98CpIMU45Jz5fc/MsPqeh4HDTylwSSy9u7FsShqi2H5K6h
q+K8aNJsxHWQLjgNF9hM/DN/iV1cHJnxMyp9IRjLGMPUIuQb6cKieMP8+wtSNxia
H0QWQBtevef09T5eVrcvV7SdBo0kasF/qHYAVfrCcdbeJeBYkyjBwWT4KoFh9H9y
L6hA/WWLNUThshI5QDj4yc+nfJ5bKn9cj8E+RU6G3jvLhz+kbookMyyDT0RkDYiH
fCa4w/jNJqNnD37SZ3RWXw504lOjDVEBbGnRnt8Q+cXspOBzIx2c5PVOOx85rsR1
uxDLFp4nMZDrTxmRN7zx6iiaAZxNrD1xMbuSWTQPbMsvCsNKXwclkTV3Bg21tbwI
fpuQeU1IFDM/tu95fb05I14SFwHDJOHQ6Voa724xIzlz+YQKtsMDhTPei/4SpK4l
kL+7AnOzFRJrOOHkjCPzdp2Iq9WsUdmn736Lj2+5VapRiKnGcAhj7pQjUW/T6dpx
aOh+0+LvP6O6BXDPz4S7eXBXLFuFmkodedZLlDopwB87qWCu/07pSc4YFoi4yhZH
BUfPc67uQriXQ2WagDxW0nPVuyceW228mdXmxDJWwhLpZWG9JSeZ4p1MVVbmGhQs
kqlRIphkt6AHWrPe0iL7JR7NvrVfgS1Wxn4aJmUTVYmnwybIA7booXfgO2m0Oov/
F5sFuwyyLa13zKeydIzKvqnznr2WazZPAaG4chw3rtZAwbsgtKDtApbCFxuMtRtz
HHXeY10KZUaKL+pLVyDrPE7HXYDm7Cw03+F0bz0/rgKqm2BnNEsGvqTEChuApB6w
QIpSubXacpDe0OaqQod1tLiM9U+KHnJdFETwNlDk5oeu8U3TGpoJshvfEQHCKu0N
5mvS22UuMKVDRTkbWtte/GpGVis3GBWv/bsDt52o/IQbleJAcAw7cVHQLEw0ciLN
i6+WRuK6jGmQAKGK7DXAhbiDySZZpkB5Eq+ZmHeNutiGM7vufXs9rk7VYeoT0LLJ
PttHEpTxhx2FgquqWOD9ZY/aDrtsrSK7pVLZs7QBmCqg1H6/99khIJVqAUJtk98q
GDtLQxCTjYUigfVyKvSL+kCVkDoclueZ2IY2BsnmQ5DqNjOuxiVBEQsbc7CC88wk
K/WT6dt7+TNMufpPY+FZlayCeeSdrXxqMr8PszhfFKq52o8l4TatSN8iuoVHeSaC
u/iDQtdXk8SHby7ScSSSmXn+8DZoObC2F9jE4C3vTv5w3l1MRZgcyviJwHqUg+f7
JyBLTYfCmrTf89Dc/phV4vFuHjOdLdluTvH1RnGJgSHEcK8HMo8SpzUkjUQFYFMT
vur3QXc8a8HZznjuqQzk170/BcXK/aJDt9wJCOMSJ5vuuTiN7T6KphUPZ6SGhVe+
njKJdoy99OThkmH2gmG9i+LXDfvXm2TqDL0O05mwIluLDa8PNJ0EcDRdhpGfr+cu
cv6A6WlfUmlM8tQPhBJyDITsGZX0wNUdh1IzpBj3r4Rw8X3eVflnLOXmtSvjZ3OB
RwaHxRQKIvFnmsQDbuOA5ZmZw0Mbju8+G+BRKLw5xVj9/kxRivm3tqCTYY8czw2H
ZioMmrr8qTBhHq4V/eW71FA+pWGxfnQSgl7Z5KGKq9x8uYEkhqBZzQiswVIyEvyb
+TztHpWC2ek/WYWMuwg64gPFuW/irYlRRyOJyZGNeOs1cvJ+lCC7wAS/RYECuq5r
vM1mZpVYVbu4qHku7JCprizrV2EHS4gnAmTGOKgjcLP83RbNRk5cjBJA1NWqOWz5
Lpi1RDlUVQFD0Pk2mOJLhuaIs6iEmtiwbc6PO7e6IUy+ai/Lk9NbahpBth7IZTGw
J4u8GGdJ8WMjDTzkJq2G8xv8GhY+xdvr4SIaLk/dcpJnAcSz4W5cP/yto/Md+0Mp
Q1yni85mR8bkOpfoDiy+uFU2+8RDkyZczA2Opv4XJnXSDFjs6sqduk80C+VpMLRT
6sgJDto7pVi64CnV5GqV85JzoqS7d7SODJcZnw6d//gbQNh0bAd+WhSXX+Z0gxNb
zZ3Zti4wAcR46TPOtVjZphSgFJ81b/KcQ18n7pXqlzKjUweL9HD0JH1IdA2meBRb
GEpZt5kQ2+9pXh2gUN1ZihEb6v/Uw+dZsU4eTKZXY2fVAootIOYj/GK61qySStBX
qyEcNN/FyFwhK2qpdsOJqZX3pZe/2wJo+fvrHLRK00mH1hWLoFNQ1cuC8zUdYQmB
IsBQRoP7d32NsZ70ZIh3aabXKRtC0t8Nk7lRlBAKRJLvdmKFRKidLcb6dvpTiTJP
NKvb69gVqibS9A1IcQp6RJwVWOkLBsVwD0cV5HZT00hq5DBvtn/IuEl88QGQBdpx
J+omawrg8gMDu2f9GRuNWXQpDRPmB6vU7fa+O0dHQs8vVqQB5vMXgCb5jzEe+Opf
M8u3ajRulZ2XjSmj9SPf9EdkQxm67/WHHm3brgFmrMQ+Ddq2bg5FNOkK4hVn4Tl3
ygzSZSBvVBAIPGffKcwm5ciIKlm2J4LzYKRFhtCIjlCOc+BjiqXc43W+/1niL19+
tgU8SA0SpNrr5XA0nq5p8wS1OpOwN3xx/y5jBVJCpuHM9fhMYbfcS2pVrGTefb0L
nStZUpCgPmRadsdFfCUZfu/ZsJXoqHrD28JrXpzhufBn0VG5ScD1X7GQHjcnt+NO
ER7d2QMo/qKLAdLQ8ids/WJxxCFLjPIYkbvkVjNnAFJJD5L7aOq6aHIu82EZcj0H
nbgoDm/R/BVQbfLYtN7iOlTH0AkuLzhPwArp0H1CUvt3eyI2J4gfl91GK5nyLJov
k5VExmJS88xvr5KSh3gCzcaaq68GQisU7RI69DmZ+bnsG6P/KKbkkteY39r2VUtf
sfoOckMJKunSfZ11x6sQCseaB/FUAWFERN9Oy0Vgnh4g/OZN0dSlHYd5ZHK/UgTl
IDeI4+1rb3avzScPdXgOiE+hviYZn+SFpyXBl2ezFnvxx57z90vu4hmN6fXY4cls
5rSJ8kikVmSlgr8VW7Ue5jYEx6DkZ5WAdYLVNrlcy71oI+BPzaIABZdsjOC2KYo0
PJTmaVG6iSbmZHTTP5D27j0dvA1tgJ45i95Tjsj/UtapqYYYag+2y0JO6935Sa8F
TgPLa6tnOrqgkqh3GaAIZBemjDYeu9Q0w2fT1nhsWGZ+mVMiuMZi2Ax0O61ZrPfX
amGlAFTT/wVyvBiMP3cdV3rf0Eevv3PSCb4jDTZfAho8WQtAsoI0DkXsCfaQeTNj
LO4PkYvNFlefHCYQxH7hubwvmrGW1ZKkxvWnNUOx/dK8ant5ubL40CqefQa8upH2
JU41fATihQBaJbBzsPpmEjyVllrBDMzC3/eUkolcyPDzV9W4Lu8VBzty0sD9sXYQ
TcNPkyM6Pi/UfYAqcA+GJAFxhY1MPCRf0Pk6WBqnf6bu6TIxAx/QjgAWTmQae2yp
bVkAd7akPPeeAF+Sk1r+iLqxWvWdYwZPiXdB9mObe+wBP/3TJezD1l/i6c1r8JXO
YyvmEJcvrLQMfJnIAkgqxiDJMQGC3IaxUN53rz24Mwcl6tiEfXmPysze4jS45hNx
cAzB5pcQOsPEtuYz4O1tLHvG15EC7lnfAc2OrGkTY4/dwTVQ87Gru33qSAr2kEdu
QztLD24by7G3tmm/N5iykU4a2kjbRWqsNJZTUdV3N7iPTyT1V17APVl3mEmsZmSZ
8YwIdeaX4CcrJCGDZdVeQrkmoV2HoXG3FjEYykCOutjLYlM90BoVJl6/mxDw/QTJ
WajkRTfcGm9egHY7Fm5qibzkvaBz+YjePwiL0REEeI1DOIsfpMJ4QkG7LK0kQ63F
RzYOd8gSDNbkTXdkGVAzZ0TL3YlobjaKQ3Wkhrah6AihbctntK+NeMQAmMV5YZbd
I44tdy9+Et6JFFH+4eKZraMLOwfFkNMMr5SNML4mRBMAkLK3uoqX0LXSigBtgh/8
MOy4+9Cb8z0pRAEfh/Eqzi+8y5yX4THMTU+rt9Be+EIRWuedOE8V/vvrYmWHjUaF
LAliTtfuywkZw02UcgzI8/2fwIq+WmWQ+Vj9IFYid6mi0EhbMbP9ULRHi1ye9eIt
TtpmxXnk0hCwFLHbTW+M5unuenPjV0C1Crj12uaf1THQeXprDpi4peXJ44X9+Ifz
8MuKLDsJMyJ+QzEctU0TMWACyeCu8egaKE2+6wuyNlM7SLMMDylwUvrleHNFIXcR
j7uVZzTvdLxdY0nyS+LN3jbw1NYBMhyAeFsLRHD5g/diDZsTp8o9HAu/Lq+DYm5Y
f9UaiSAwuSNw7sVBa1ABfv1oWsodjaaCl73bl3I3bbwG8SSIKPMj73WzPyQ4+If0
OAJWo2vz4m20a0GFy+7HEPxlS/PF5aR5a9E4s1kqOdsdXWcsjOQKdKLRAT3ikuPl
kytclGNT97oqw6GGXAaVGQ8djDxWJKqWvaUp9da8WRkSZVATrktGAhjUKxtiioJf
ZxKrzaQAyozoWIhgwSfvAfjRm5I12mVRge8wRG1IUDLaOI87nIPScWXekG8ypAgg
x1YsR/+uBuGn9ct+xP7tjllfcZtLZ6tyZx2oW5RnbtKBZy592KkeuMDtiPV6imqg
6dbrdMwvtu+Wtj08HaBX6rf0JVeohCWxZJ2W8IGHHmKYUY+pFSFilqKQv8PM1gxw
QUaCXlZG3nHYn+ilwpJEMTL2aEfCzMMAtfAb29nhErerOqcLFOuF8eplCjo+pd03
jfiS4ROhjM8C5edBJpTMkVvIZCRSjMagmUQy4RBv5olbquN8tPqjqFsogkzRBPdI
jUP3NZSuh17LLpseulTMw6zUD9TRZDTg+PQUxwiL2E+SVGmGhmbN8KN+hlGKDmfx
UpjIQcE/9wlr5MinJcmnPuD7SF2BI+13z7i25SH+dxMcV/0dIKTtVz49ebsEdo/5
ec5sScrI3IGcYY4mmtoADR2K7M5jSYFSPHwVnXtl2cnJ9hsVBKZ7/+jd/LfC5Jui
e5jcon6bZBHZEdCRdkcz+RIZfkpCbXW/LYSCV8TfaNjwXaSSX2xKPMpG7y9BxUrS
rLA0OHPSwIcjQiIBGu6BFJPub/1aCTOUpa/nE2uAJ1kuJIpSlTGPqoWZAPK/D348
XKMFt5wIJRG8BQn/j9OF/M9gv3oCXRbyKag00vrrVaZEJj1ItCA9Dz3X4lE/rTFn
43G7mY39kw/xeNm1M5lN6e1wCgglnybBCqyzGq5fC5hJjlJLntLzmVWVrccbtLSL
kvOg5T+keRDMWQwaK3vJd0EJXrDr8cHG/E6CbryzK4sRydaG/LetEbeFlpf8AXJ/
NR/PoyyXF3qi3c0zEWfzNneEzelFMaGA6lfJf4GX0CNa1UI6oqCixrWj+t8+XTXI
/FVVa8kTKVyiQaklmik/y0f/b7V540Iry2z1kKspBYUDQbBiPQfghYOdtgD0COEy
T/kwixOhWHkv0eK0yHVgcquuiVBq7nnPbdX7GeIS3R3p2y8A490MDsAHo59HnF6j
T7S0Dndv9OUB4Xujhe++nmXHd1BDpXy+HmmZNPB3T3zLmAXZhJWJEYHJ+e3aeVXm
OoKdH/9/6EXdMqouhHe4NIgxKXGI6xj9bz/o+fIiJLvQ6ORqyWh96678xTfk3IZI
fkgRnOeUvJVjW4yja3WouZIA+YwMUX+tYfdt5IAz2GgvWZcJ1qgnoJB6QUXYBFeU
B4cMdQBU9/eXeBBJSl0AcT+SV2LDUiF5QpgBT2OhqYH32UL7FMjqMfFGV6hwlBpm
ZJMYhNUwVAM4o+X4i68I/91nXy3cajgyBC4Hxm540c5q0xgDFKUvV4RnQxGyOqnm
wGRJ52fFBCHDLfpRKIE/SwlA9gfeNyeGAh4GrOoFR//D8IJ7pwH+Y6FDWirlkR5k
4HMEkNhq4GB5jL0XXrA4dCkYk+7XKH020NYAAQbf0IbOQJD4QNyUdGItPIVwFPAX
L8JCbAi3B2kY17gC+XPeUe+kJZGBDjmlfC5ZUvcyH9Y+1qnO4eUSuOh2464qWT22
D28KpGcOjRgaI33/L3HFP5xF3aK6Reu6T8WGRc80TABHj+7hUJzH2G8ZIQPrJpGg
lzQ5gVdeF3xHUEQNyuty5DbWk4aGn0JrgSmmqvzHCoMY6x9IDI0UNKjVupaxMs6r
/iZlVNY+Rtkq68L6grB9C4gJgb9zyKNMkqXXxkDXikj+2Pq11YFCN6MinuyzSfp5
w8EoHJ9z2Z02PCWR/CLf6XvlIafR/JKa6N6Db5ualujHTuTAOEImLcWM3mOLyyD0
l+0OXkNXDL3ByKa1Ozx291d1lcvYjaNJt+VLtFH1EliQfLm9qFDPltHRy1R6HJQS
`pragma protect end_protected
