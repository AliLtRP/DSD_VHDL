// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:29 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KPDokxdjQtDedk7dG0sap19+hRc6/xgGtiwxl+FDnmA/kTX97ztD+wYDlxgtoD/z
hbnCUdie5vBv/C2byFeYPy/1rM1ntI4LrwL/21t/8LPc9czcIm+Uol0n5OzjtJ9K
/63PnLTdpNKcnakNqjMkHD93EqV/rIn+gHXgTgBBGz8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 63216)
w6lGLleTUhbu0hmHuVgTyOsPbJODa7/+VXDnMCfOIvSsaokINIIDGhAnAiHO6op9
IhK5RybuE58V8m9Y0qVF3VJDWDxHdHLDKnSSYcGUpn1l74mpiVBxVn+EFDey0FCK
8+bwMLFmwN2i/QySZ9teAqh5lv3kErRrJZteJIukZoyXfqfVYTw3qIrAi4vAn59f
AMKZEyWhIc1FhIINPbVbkfa1oqcB6K0N4GjPjky3i3rp0B/2TSMhm3BNKBtH4IHO
oYPrveM9HRub04xcUzjP25zc3o/31lSj9OWgeiakFuQEEwCnwt8YbCAypOpmkj0Y
L3hIe4fJZ5Q5/cJ5pqGtfwhE9hlemzFADc/ZPCya9hfi6gitENyL9WMXVdvL+Voh
e9hcl8olSWkumoIgHYXL7FTNtzzdiPadx3Q9GBG5QyPAkt7IKz5xuSBWReHbC2iK
1Sh9zEUjO0iIMf6S8lFpIGXkGW2LCX+qgueIYaBQLwWTP3caGpgcd0+++3SN5obC
Qq/Xx6xiLux/ARmbh1+OsapFxsl393p9C3mZTgBsI+XDEwJeXJqnu7+JKscgcQp9
mqCRY9DIF7f31ipc23AF8Nmyq8SihngqUSum80xRSyEGV5hRau1AHNE9+zAQ1pam
6GD5ncZZkItsyomMZypHmE9U8NAmMJIgAqqkdDxqiOfLdF3fZwCn0EU+0v8lYwbM
6jP8izKhJ1oqJpWEYyDok4Wq3meDwtutU9VoGlri3uB1ETRwafbPH2lrylcayQ+B
+eUa1SKcOAhckcyFsFjy2qIWsY3aXGq9okMYYMW8GOW4JUIbbsBWCNuuMlY6FKWr
aLoWrXkwqMBLtk5LEiE6AuwcgguvWZpszMPrMApKA6Bjfh64Bav93RSq6XiYseVo
afzXCK6WaMjVgEsgHtMTCwl1p4+yZ2jPBQnhPpRx2zox+YUlXW2P+Ty/FqOK5wwL
Slm4T+MafUj58FYcUe7+ze141Fn9y40iyaK8ViLTk15dyT2uEyppSUY1oPOrhshf
BHfAXp37yXJXBQRgsOIQ+mMZW0nq56bFuVeFYQ9nV2yyTA3qXhigOP3EiNancQAt
x+mn+KphYwYa/FsqiUGqrB8IjOx09k7sOnj6JBdxZtBQB5aECResh/R59bWSSmek
RKNvkHDQ4+zPxS8sNnpGcAAuel4QH2Uiv6VkzPMDxalitV9aG88IiNcztoRonV85
G66cbQgrC3CKIZhm5Yh/or0u79aLrZVNYQB2j56dKtvZXVEL3UFW2U/yYGT7v3PP
n9CcYJXDxSjPxMUdH+M1Gc9P+ORvNQ2+vk0zgXjrb69mGQE7I6WUlmbnzix9dEbG
Wm6/PDLLfpUuRr1iks7AkeMp/NCmZiY02pHZCg+Q6RpOz9mwp0+RIpNNXfyGRpRU
8bIwMOmZPz2wRY9Fi0xIXYs3+P1IXX6uinBBn8u5L5rmCIvao0wNdV9vnT8XcSza
emrEgLhZCYODNDlIxOy29gfwRT+sxvUvu7DQ/qmdRSOKRZrM82alJH8X1YlQlKuL
9ibiXYlC/kKB+JorhBAFAZLHbsGpVVeUonSlB7e/mIS++pCm01oJ3Ajgpryyvbdi
T/YXh9ORdw/5Ro2TG4ldWNog5+Megpjti/yCEh1MmTXBwDeM/oXhJAFHXeXJh0+f
Z0UQjggqHte1m/Y+yhYZY9SC8U41qLELYj1UNbJLHG9EMxKOa2WyKnHN5m3SZqRo
1ZDTbANuStjYkWq/zOhty4y6hJjj5xSD4zOG7+Gf80/iQH1iI9tqsdTRMA+SLzmv
47QItrSssKbRWcKgKaUB1kq6/tYgCKl3jq4+xZP4YZrXOOFNkZ8brvL+kUZm1dS0
L3VjshdEXpHELNfJ33Og7CZWRWpdxJJJn+UusSb1UguVuseAD7WT6/ezCsFxhUJw
z0zqi01KrYKS/gqSyOCWNP/ZdgF6kF9vB9Ocw7ElzMjWqfDffePtGhAR0GzcNUVn
4bZ6XD3VnX/6SkqRaGVg2q3EAMTFh6N+WM/RlXySFRJYVn91lwrInn4LJWygNOGO
ijZ0TJBEa9C/YymRfYO68OMOQONZegdyJj731At8b9P6w/v53PyX69JZkQaTqpg6
/RXbvZdPe+3EVsCB9nVwDzzWk36Kt8KnbTz35wl2yudp+ds85pcDdmmVjoCnG5bf
t2G1wH9S7v6HaHja8nN8vovckJGuqEu0wjz58fbtyBgYomjGVJbiNlIKoZWUlk4P
S/hofaj+BhtJCGPQALaKWxu2aKKv9yqztfATy/Jj3LRx0Rdu4u9pWoY9IxTjpbgT
wfD7c0rfIdaInlhETgxK5c+tk8nNTfAflwLqst4rWk+u9Yh63tBoHljQY39U/QPB
/fuunCCy18GV738H6aMYRj7U0SjN2LYFyVbcJc786XwCyUG0CJesi8wjHkcdTflr
jwdQn8w6XPNPrNLoMKSJtBZAlOJeT/f2MVeQlWrixU00/Utg6DPWy7YkNRWVSCf2
eI2gCTwB2c10FChSSnYAfoM/nCwpapcb5RrjcbierH5n6Wp8Zaq1n+8UEcLmolZj
LpTO43opb1WA1wnkH0ocuIXIki2ifFVHThX40rIuRaz5YhEUT6nG93Kx4RvOhXFu
LSd8eZ1V5ib9sUr6z4ScPbOd3FYd7IVCHXTKMmx5ZcX7AZPjg3VGjVGOYYwXHcty
rAdOm5dFnvuts5JOtRjr29eOWA0Gb4xYTb7YoTGOTeNH029hTPQ+wRa9irUPFClD
PEPo/DhSWe7VjvHUFlA1q37rtZqcfAsPgSYvg3HXNkxp5yvzSqz045PczyBHt/Tk
NX19PUmRl+ghUvjh1yvKMg8/COZaRnbRYUsjIUcaUXIBYEZvOZcgK0bqWKHu0X9Z
Ka15otth0toZwdIaLSW5MxwQxjz/x4duum0s6mid+cfeHQx4WE1+bDoJxGLBnIyK
YyMJrflpb10qw5/Sw89vxvylQU1MvjBRwwz2Z29TevA8j0KgMq7KohmszTvxIxSq
ma98CylivtgRltHHTsniizsiFZT2RsqBRa7Yr6AEX3C5u9d6GP2AcUAX2S1RuMiv
4hzNpL8EnGz71g8cxwGKalludUOtkutUIaEEpb1DaWM+2htFa1RkvsRuMgbDP1ed
A1CAqAmsXDQQqgPuZhF5Vf4qxViiCBol8RxJdCjvF7J+yyxr8J/tNe5gOMqWkZwU
I/PJWTNpiJ4xegV8MYFJ5MDoBN02nu8bIy6utbTA8jOJD7QflTNuu7b5pO0cFs1l
weiQAW7ADbpAemVkEVF7iWeYPZO0yQ1eO56pVn7PGf4sUuMFwAWDqUc2ys14usAP
dKkcaGaYNhAk28gaHIICU2vhCQdxfivQ3g0La2W3Plx1w3wY6J2k/iNmcwMmR0cG
IVNZuIAhNdjhqiw+UVq0pmpN8x0UkA7a0I7E/Lp/DVTJ9ug80BjaqN58vy8+CPAh
dF6/sFQ/BQCk1p3qJegOYgAf/+8VdP1ZK/4VgG+KFOL6CThs8reZEpmFqWeuLOHw
dY/73R/bq3SqfUY7Np69vbsgx++kcJein3jkQZvvyYjHlV0wLUmwJ1u3Lj+p3yJO
/3HcdwSAs+frXbIaUSp6XI7FQdW2wliJsqFTVnTGqtZeYBOLMX05C1qiol//IbH9
IakBreptMk9XQX1C6Ts7LT4M4n42ZkLQs4RlkskCstP9CIJ0N3ERJGNnVoVxo5Ab
7NVe+3isUd7ae6iLOw7+N0hnQ8NFQ6iRzozw829+EJIU8AGIOMEyJ2FSfutbp1an
RnWrMyQiSaEGUcAlBUTX/3v782vVP+Dfg6JV0WGyNa7+C74FOuSjoqywfOPceu/5
ZUO3jtHmpJrXHEau6HGKK7xvMAOxucoE2e/gXrSz6HLYa1A0g+R0I21n/ttnMtx4
DcadVyCBnkzYO4D6sRpU1Vd/ip0qvQ5xUWTMcd0QjYIX37bVZcJW8ffp4y0Z2cHQ
l+TpB63mXBpwkCNbmX02zSMy5WvEZ0qcbe3qPeOp5bPJ5dnHPj5HsFY1DSYLmjnT
lAfrHHjXVPAoDJtHPOkHQf47jTZ3B5JQaynuYcyszOePiW/ksVDiRXfwcYZJl4Cf
5Q8hug5K6vmUBx37tDua+xtfzPY2aPMuTsWwq+tpxXpALDME0FPL2obIYAyLJnq2
C0BS2lsZFvkst6x82ELP3CCayU8tUh6cirsjHxk2glJX7Ie2ULrPDKMlw+FT7ajK
SS1EghgrJl8+hZOxSie/HZOfW0PzIDiAgKJ+8a1X1sbXvU2owm8srEWsTcT5ndyl
QCP/l79fgkt9jzxL3GwuNfKEgr7W7CGguSHFgl8q0uOg3zcaWPAJF67r6Ojlh8aa
+VFPu3/dTUeM5Xq3w+y97qbl6ClMpOm8cdJcAHSTUwwcI3OgA4UZetwzmmAI81mc
nGficYJjvrei+FGdyXp8VWsmcyeZ9Z5Io7f2UTNosyGNDecVz0WbiUFbzNZCZLx0
TnYAXWM27JCmat4C89Pv7v5DIAShM79VAoWxDRLaDDCEJtm1P7nVmty4quWbXSee
y5tW14TRyijKrZ4raKfup0u/yVaPolUJBBSr5ZN+YVHpigJhAhWUCCaoPdO22lQ6
cY2BK+bT4lJaQLI0p7rQmxJsjxAM4ZCZuXMfe5NEc8LM9cb6H/YPgpuZgPZs382r
K3SBdNJCUMESqe3rXacIY8hG0SFO16yT1wXbyJ7BKLweOnmbs8KIapKsCX/Yutq3
mQg9FLZxYT8iZrIr7u3UFpsGdZxm05WoOYTkbS1/jKpeJ8e2do7q0bqHR3fzgHq3
Z6UKeLV93RUiSeS8jZmwboqkSphad5xcJazmRIJoq5C7cCGh7YAAUx7SETzJyojj
jKRsV5K4Vl8u1HMIFfkZu1jM2jJgz6ohi1o3/ee80NybJch080nksXPtGQMRhOPy
+nzKZVlDChlJovTqMq2bVE6uGi+Hbdd8G8P+fQztGM2KwTRs4vahuvPsRoDHwgL+
7gge+BIj7uNCL/yBi+OcGkwhJjeq0CCEz3H4ANM7lfoKPUQilwGUiV/2OCPp7nzu
zuhqU010ItlybwAo4n9paz9Y3UuyIQP8aCjnyrMi5ZHw0/pmSzxX+7h52CebdcAV
/J3PzSDE4lzKWuIH2Wjv1sv4FIGNKIZ+MuZTxyzRT+/cT+eVwDJwzKEFzgIJ53XG
+i97uQtPCnHpru8I07pnKvZnauB5qN0J9WzTyTj3qbuLbiys/nm7J1rMAcHFunNT
jI/JrJ2dTqaMhmwLhRo9ZiZtPJetS44LFRH5dmanhtWg56f5dfAnIXYq9WN+u0/2
KXO/ZiI61QxWA0uXEwsUlVW6jZIqkWoa+n4ALDS/zMSk1yYsgajROh6tGDOVt21s
6hnIGGfQttTuoP0J306fVrTcoTP6QmG7q6ZRnPllQGzo3g9RJFf982Sa0NXZu+HV
QEklVYB3AuyI1xZ7kyVyrXPHjFe4rX2rxbMzlmO6qEJ+4eEfo+a9G8xArFBaK9Zk
Ses7J/O32x1VdUcyA+ZtgD4mUI8XdKJs93z04eB9WoiF8cX4m7lK4pjgLD0P8diy
FE+8l6nEiLnVK5oseisAm+d5xVzYg324p3Oa6buReSCEe4UG0HGcoOO4JTF1iuqI
9RrJbHk7Dw19FfubDyS/wcYuxmNEVw1lH0wZZkFZpkz28Wgw571jAJFrOunXVxK/
zf7V1mmRnTzQs24zTTJvIz+PFeD0j1xrMPkB4K7OIQsGSlE1jzAnjKjGq6Z2inbE
2gWA8TqYIBzrqbqz/wWPBrzrK7u5HVf3w+/Abh14V4VHzzXiRVOkr/J3BveoE55j
kEI9bfWmzHpSAa9f38Cqo3OzcGwDhdkJZ3AYrJcYMYAFFwZAjyggwcqGOdUPVVaF
c8GuBglhY11Gduo/+ff9lpzHmYfYuOlQvHwF3g2iYt9Pj7XnYNtfLtwCaxWMdjT3
B5aB87fAl5j7ya5vg9aqB/Ztet/KLBo9KKTYBnMs+WjDJoUjkajdoC/+AOekfbbw
OM295d90VTvi+Bq1kMfd1GOmCfn6VEGLKPbxAJ0Ao9RpmA/FSIE03LJLaY05zDVj
Yj2i2vcRMaG5iFCAnh+GxVvQoC1WCMyndz7ZtX+QFePms3aTIkSWIDp5It7/CYnp
yYkr9qrYlxe9DZjKHp/fCEL6SWERdNZRyUPYhAG/o4ztCH2v1TCkaD1Aaa4fBUQD
uyrI15ycTGE0eTxTIWCSGSB+0hpUDiOiQlMymPPsyoKuZtgqv8G4Ijwigq5q6j3m
hMxnxs+RD515vTJo5g8wNy9KcqjhbVvjiYqpwwF7axnIYK6ddQuM/x1dqURGas7S
k8S/i3wcDVubfEXoCDkge5tFgwyL6hRfLDqxBP/sUngNC6yV7ymErPzx/tTnGRB4
Pw2b2a12L2OtSD56v+rZyTIk/+ZCEBJyYlXYzs7q2ovw5R1Df14youhQKjSOuCVh
4pO6irlwSiZqc0LVMuxepXq4MuFJV4CwqsNq+s1zamJhjjasZX3Y+QcCzN9KQrRA
emawUbGUmN3OYC07Wt0BKtVESbndQSKS+PX5E71NnPG9kGqWb9Z6Fal4XrpzLzjM
xLNVl7I84B6mF62kOcoxPIadrJ6On5+1qflIhjxUNEj9IGo4FGH9t1o6hPo3r6R/
Zjm4OPoHAF3aQKAZYqnoqlFw/w0WjsVCeohZqKiRNylrNx9xjJA3pt45GXhqK1w3
ft3vJkA0x95WW6ZjCf1x1yp185+tBe6YIReTJI3dqpwbI+xWh1aRX0IP+Ys+ay/2
lWPdEWTfJK4I/TH0wTSFp3BeJEpSkjS7Kt9VBPfrPJcl7hr3G3OtMKP5wsnI41Fv
v/odLO35LOlIHXbBEec+s/iTS1idKNnE6mFNIUQufkhqaZYgKYGFzqtNusBh7mU5
RT59sjY9TSyQBxehdhZRgo5NAVTHwagC7l1F7oDmhO/9v+CYr24AB9xfW3x3S6Ph
/TQgrRbIu9I0icjGgj3rJWtsy1mvf8tN+k6AiT+LrUM86ZBN8b9niDARNk60pvuF
rRnPGm7e0W1QGDSszL6PzT4CgeVEITew0nnzL1V0pzD2zMouGHiVIUZoflFPoO1L
92v4RovvZ1167pUO+Eu+rCKQLxq0rw98cebP/YLQYeE4bkdIF1F2NFzacnZtQrp5
iKr3d/EtH3I0/7PfTwSqO34OJgJXcQsn/KOr55IOoJUnd1Ca9QD1xN2ucftIl+YA
1Xyz2zmGJGdXC1BgBEmveHEr+oJlVbf8hmtdm+Sd+69xIIMaGpsFehiYy9XQAiqP
jvUsU73tVKP8gVuh9kq5BMBh+erGa82LzbEFEhaW1uoIkivS9MBFgYXK7ikcodLI
WKN+TwQnj1kxSyHeFVyn0GMfdSmTHO9vBgZEuXeVNxp6l1jXL/LmejQPLlYgjtoW
zTAVLmiBE6MxaNz/XKkcz6uCktzqXG4AY4Vbmz7a/yB7K3AV6Sgxoyjuoo2XYlPg
TJTHzu0bcEp4RmjXBtMzRiq93mcYAJ129ovOGkxvzD6h71vclMP5XYFMhRVYysK9
sgDie4Tlmq4PxIOYcPclDQFFJiaj7t2lkOi4fMQTBO7a+0Xog9BrcfEy7r+zZHZD
EegvHSqQyumaQPFq0P8cXFFF/zbK2ICcsJej8L3Y9zJctit9vMhzOfl3IY4nyZ5f
i2bcnPTfYAVYY/BWanioSbQ0ktNV/RPGcREGDCN5sDJWxggKOuUQsgq0mxCCMRnU
SclGyvgI8iE3e4e9PSbcORMSgClX2W0DNUXyufaJWZ8mA0Y+6lgM4l+OmNKA2T8T
Qbade8iIe+rEvVlDUpIRJXJTGUzkZN9bvUE4HpkkiOOoMgmqFRurs8WK8JZVmcXL
ecpz6ZpBGk/8zwufKbnmvn0ZLlFHcLcIzdZDpbn74LpIhbiEX8hNp02mULjah0GO
HKGvxsiJl6BsJ+NT8o5XKVx1qM3DXTkbGEoMM0VxoGKfnJoOaImD5M5MZxDRPGno
xFMSyIUG+HIb6jRIw7ow8j4jjlZTS45NEH7LSnCpwoEv+0RXUMMUP/neCcGsbmSH
kGM8tSXXJ09NNQDu+tt4j0WIZQ/Z3SxIYOnWiPidUEAETfwyXxotc6I5Ibnzj2y9
J2K2pde33RX8LZGFFVgD94aZ+EU4dIn09ckmjlj6tAUl64nS3ilWUx7x9ZeUZPig
qsG8TrzNhU6nTjhshqy9bvX/+BfRROAVhsnygGTj3sKPsQpG17DghxINwwY0TyPD
IXV7Ib5JHeOCrlJLmHWHTCI27Op5unuKdIzpdlqe51IaQz/X/27mdRg9D627jt/L
ecXtECnpzxycBPEphaC9Dy+xmBxB4FuQ2klLfiHzNq+iBFitbnkeY6D+wFPjuR42
dpX9Dj51gASiqDUvgSYIcKnT+sj52HWbtBUTORC1/PnGn1mw0jhfUy2xj6jrxTz9
tMzKo96VGrP4AU0B/W436nQ5lZdhXGVLFd/W8RF5guDjGRxVzA+an6vvPqZcJHnM
+PkOxA7rKsfvlaq6oDFJBMj/aMsLfvttMtQkrTQxw8O80sfVS0F6mG31ooEsyfYA
Ly+PCf7sE09QClmMHCyJzvKmbVJxyWfJtjGliumWM7l7/HjQe4n33EbWYIr7X1p5
NqsYu5Pq35Qh7rtcJ32dcnv3GIHQ5CcjZqN4l6E/xNJdQ867JEkVwIHepSQMOVZR
b+Qctou3kUX1TNLIfIJKbfpfEYYWye50zXYNyf3UiMtcDjV2xL5DnsRNPl4Uq8ZM
I0qHBWXZ63kWPApB81eaYTkz5/fUpaPHTKvR1F6mbmMiYwo62BZSYS93drXpKt6z
KdYwloYp2G9yog8DyCq/foVWrmeZgdzQJrzcxMMxRr3xiPf0IAqRBqlwfT2l5nbf
zmGSFKS6yhHQJURIAVejBp9I6GPEEv2igHqx3TfpJMcUbSF46wjLziHENzVrNdUX
+UIVCDBe3wtkEpYMZ2+24+So3LbRzNlbrjBFSMpLuO7j586M9ybQ6UiKj14q3JFb
2PPq6nfNi1DQKvPMuKpBTYgpOi/urivz8976MzXk9WnVZN42mGwQceJ2FjtZMB7m
8ndRWDBTg+jAnEqEqpSnguGCNiSg9FKuod+zlfjyaCz08EJzT+SN7llViOZhFakj
AhsOMzInZ96ignrJbY6W4tgQL1GNj09YGrzPIsC2fhy+1HoEQ1+LFdb7O96pb4pk
q+cF6H4gsU2DW6wm3GJgFiUVawDbAqdoJKmKxp8OBua6GblKTILf/SLdE4UwdBQp
+D/dS6nQdt0YF3oxo3nCyyXvvpj2N77nzQ3ZicRy6Lqd2AEguRATDTqltLaxklzt
evMT364boCs76wUEl6AY5ErHriInMXp3mhdId2bqReR1o4TCvHPOBzAdj6BppCWz
jh9X0rqXczeQ0Hwxq6QUh7NSfgXrBTXoi8uDLtnz39YCRlI49wRC02yPY8osskii
GFpcaO8yMgos7Blm90JszwLopEJHo4N8FXG1gV82bdvEW5TosD1Iy3OS3iP5DI07
qJBxaIA6FRcDSM5bbX6vqkMBWMeBImJpFXL4eypOOhRVm8rHvrCPbWcPGR7enySR
rMUcSQrd/AKqNS7S+PcEBgil40bFM9/GsMdL6LNBts3mgjOZb6/my+kvRu58QESE
BY67bthVNzfv1QclhDpKHwxR/jRI4q/yuml5wqPN3MuayIusw3hrx7nsrVmIcPwf
uoBpLbBchk4/jdwqQasdlHem5yW+ox60DUvuAQjIcKF995eqoNm7mo/GWjVTMxx0
zWGrvn9/6vD1kYMC9kjKwj9nMyqE+w7eVKhbq4iX9Ed960UBjBSTqlW9l4JS/dx2
YxHZtPJEb3JN7xyUq3C0OQ4CWxyYXeMpm4dSGWta1Lf8Nu/YOHSDzIASQ496VpeE
J/zWlm4WuYXvQJHQ9ek/FA0Pfnhu9zbwPkXpPNSHgV9T6vKFHC2ZfJF1Opgz0Bpt
Wlh8WjXJsk1prELjMt41+4ei2fht/3BpP62YLnm5SYUAZhAvW8LMmIoxwjz0/Jot
4KIdckJRlJXK8fEIdmc3fMzWsIbiojowbmhSaGfGB9NjQkLc8YASScu6uuTUIR97
oqQT+JnLDjcrqo8tq3p1ipfhTUHsnWjUCRRnVS7coam+CAFdMRgDk8P0IVTvA/iG
nROzyVb3KWOQXZIuZw0wxkX3ya5xkpgIDK4obHlJPO/whEsILSjl9E3VTVo4UdOw
iJ07813VfvHai0CGYAM8dx8WmCGiiTdx5ZTHjc6409edgHp9d3Wzu08Eq7CmmPOx
F+JShlA1RczW/Mz6lwbTdrvFAAbyXL8N1Fat+62N5NWCLx6d2mwN7WZUI1xtNizv
DKskGgnMQD+VFLTdEi76jTy+hj8z4ld2i4sGT4R0ws5baNTNVWu99jIL5qv/bA9O
r9n4HNMQCMtmJjxfb4RYFxODSweEzktA7A0xkuAA+AM4XrAwmrRBjGsZ5AnJP6Yv
/PyPpUaWIWmc+BuucD9LVtjVlYKu8ys1LaomxTNWhPQc4U+azRwyiulgXZsktDj3
HGJatSkxXAJrWONvb7IXD3KjSmDyxL+DkNyB2C/Zzs5WVKLUg6T4CQxlNYACvVrx
RGGiSp7t5a37sR5m0VQE/PbP9v2UWrINnkvoXrBVFdVJQonyX7VK3K/GzwTCWSAE
5PJHNb6XX1bbcoU6cy47+sKoqXVgC5SRVSWKlE4R1NtmketzZPeHZRG1vEKEt3fT
c1DOH4jgC5wMquFYkcK6GF+J1+rcAvlsfrhTNTu8lkWiWg6Wy1edxl9cL8qIF9IX
J2efsytz3Af91l00Ryje/fLtJPcXP/UgbmSYTCX/IGfu03ed3P35/eh7GfRxJF99
ltwjb1sq6W8A8hUg7ZaUpnKvC8/LUAQZJcLrjvOrdKxP8b7j082qLXpYN46M1V9P
Jjk/RU6sQ8E0PylCwUqW0uO8s4kvyZaGbPS4z4+o7G9EwDXQF/yf7CCJSPsvKQDD
xwBFVg3r7FnNy3Bu+L//wlte0TlI26aMHaptl1wOzYaAdbQ19g37/ne3ModoV1UJ
z61ROOePIrQ+N5yxIJVk1g7HeP1zC+BGPedo1A7FYOXTZKOAZqIxI+gyDblVmx3L
INw5TqBs6PW5qkw4lCYQ1CmM44z8BW8EzX+uwVkJr8H0YZ+8v2ljWE/ERh2mjJc4
dWx+XFIGNPMrppcsLi30hZ/oBZo/Cwr55F8nuKNZvuJvY5gmifBwOa/eBVL4yh/0
9xdYG35DWyzLc6zmxacOcqGJJmJaKigRin57oWZT2I//7O3I6l0X+Ob5ogYXBEpY
s2BC1fKRPkrqlWk1ndcKS6sMSTdF2SWS1UYlx+xQKnhpKxXUsCsgeoMw5qu57pXI
i0wdblFr+kXFKXEe7zr747nScTVK+1WYZ/S03raS7Ti6x8gD9U0VIekK75B0kS7m
Glbd2RH2DbwyLRgXXKmK5KT+HRYEqhIwnLy7DsDOTUsaiwwpyQpW5HMchJoiAsD3
JJ8nKOyjETo2zMvJrz8iEHH9worTgoykDfyqgX1/TasHtZ9BHInNNirtLGwl6FJj
b/F/ne1R2ODz1gSo4BZuO+ZztYhmdugXEWfHbnGMT43py6L2wZZazGPzIgdbHo7I
mtt7SkjdFoJ7ND+pr7+Hr8hHr16Td5BAhDeDfui0DI5rkRjxtJuzaumRyaGGFcMm
kVYXx+eQJrt6HKGgpRMw8n3w5w0atBhkx7o+Ht3ktB2lE+x8SdSh9JoLv7ilouEf
pH1tJR8HI5QoNQlaUbRKgpFRKh7mtHRvE97wgDUYXZZwFSem6QfFxstx+c7vCJl5
Gz+P6FxNJ46Z25+LUzFMIsuJ+EN0Ts/30QDZjdHbwm/a59CosoUwyrXuLknse9oc
VqJTXWfwv4v+7yWhmMQI1QIhuEoVCUpPxjrWA0YjOKuUPZK80s8w2WT9BxIPJfFt
YwA5u91SEU7YyH64olW3JNziQXT8ekjVKBMXjhassPCc4F2ANlqyyp8NlYNpTY3Y
g96DfcyFPu8rJAgbelFt68igSQebZmMpxAP4L4x/9ldCPppchAejTLofCKnUhAuH
0ZmY58oDKSlRSro2RegmdgrlWobwJ8ueSNTZBhXIdQUuVI/Ckvgkj5SU2MXGNfFP
W51EobNe4sh4HF1U2FNyU2bQd4wb0NJodH+4KXk8wmhuH/xubJiJP8LR9pKuK4Lc
xHFX+ajUXlhCkCR130HLDRk5UwKJQ3getI7bRkULxer9Pl2I9Y6DaJEX8dMh+EW+
qRUvlyEBJMMjFLWq0ntVPoZPN0+ssr2s8BrS5AP18NzTUZU+cEtCm4lL8zBR1SAu
VNGhw0AmhpFo4UcHLLC25bDtsBiEsUUoTUr7cR8Hsg+3XSTLCLolH4pC/4Sf0vyK
zlotVoZZmrEE+VbGzax8pgxG/X4bBh+2xIkI+j6uC1Kdavr+BiXfq6bntBBPfnDO
8AL3krlWEZIDr25M/SO81vJ7365ujEWUkebrDUacV1F4W2cTuhosGJE2/GLAGKax
0rbC7bS2bjzjr8Uk1z7E30PDSBT2g3c4v7LEn+3Vr0dcYxaOxq4//UmkH5dXiw+U
Q0PFy7qNH8cGOXZPD435lSu84M4gTh6RNlMpeNHdWV/XHf8io3RcKLKaj6OHe+Pk
5oBYqKtHwQoNgg83gFPDSIpfSa6MTsNkqpA4vKFi9X9i0Htqde54oqOhTvY9SExQ
vARMx9gmvSYWm5pGpGxxOcT0KpKv65yB7Li3x2/dCnOzNcn+MBLw/sNA5IuYuFF2
bmJxsQYj4Z5aosLsh+4864G5E0IUJUIXvXw7Y9o4Y4FEAFodCXzMtV4+WmkHBG11
KHtatr+SeiIXTOuKLmUjUGMJIkUkoeE/xZFx4hI0p71b5WBWIOc9oSbZgWiGh10B
jm/cVLtXg8ngEowd5oy0QuIAA8rNcvlLBSKjZYCyCtx+LGTYqG4DlWcnPoR8g04n
YszCmi7MT+L5rHyzcZvOzLaVytbjejj1K1v3iWYCTkAgu09oj0IMWtbw92Qx2NUL
/ynQsh3Vq5adhIZkJQzyjXMPVt70N8a38Yltg1RGAw/GTmlqwMQZ8xEvrh9/tdBV
/HvFnULBzDEY4NSWQMvf3HbZO5I1AYT4qmI1OSL2LVH3kGlB1bXEdKevFBT/4yd2
Iu6RbR9dWsKLOl9+PFM/LW/5/lRLbK39FrAHx0fFb4RWvP3nXSBHJ+EwbUaJWzaD
9Vr/QpD0I+AYaudxxR1Fsl0FBqXIHhFzwsgyzEPZgzED/7mNCXYFCX8HUnyVyftE
WvyyciRdeReiKXRaBla4LJ0BI6VdQsu9JrxCXMKpOnx+OYcS8lJDt8+Cce7vW5lC
oPGqhSE3HQAyEzV5MebUTZr1c27aSu7fMmZFBkYnLyeRBYnsS/kGTnVcASOE6lqy
LBfc4wj7+N+QJGhBuj5dSjhiuoZaTPdkz5FxioYPRkR6ru19uTVnae9lelfb2XBo
CZGDuIckutF+09awjx1kymSGxHKfWSdIhoOsKojB9YiDUd4xqSYAnU4bQu4dAUpQ
wf8hj5IbNqM76rrpkgu0ssxs2H4RqT5bE7EqcPbpAP7NCC65XphPoH+s17KbkW99
+WsSbx8cFl874cX/HYqJJ8BDrE6P9ba7wKL1ossut4fH6IG11K2pZanQTm5+ua/Z
O9wtf5+9YtHVup4A1pFDK9AT4Z70Zm6cq9bqVsHZ1/tUZT4bTwBNjySj46lJoyGk
4vlMIZxN/PUxvylFgyx4tG2WK/xxszgUVVGBJHy1EHvW7OtAQ6xlrHELXZdVRT2/
zU3DJKFIkWuRfEKgp7/6FxhcCp45anIduQRyHpL2u37ci/q0NRq3tsj+2cQ9Mpms
hHSDaFc5YxvPYeLfNK8htKjZzPc/XABo9XO8f9HB4kjR8JXMPkxN9sWXJowoEYwr
2lFkIxpXH2Jb1DwwBZ+VvjTahM2nlUKHSPk6VbXkyX0dyeg94H0C55IwCVF7/e1Z
hR9JX+R2SXrJ3MPyS5Po8Xzv0B+e1/IW2hUrSot/kEuBy0f/gog2v99MWt4+ZtS4
F6dKtNuBO6ZPIpIc0RP1nBVEeeLxhzRme1r4OdqW5Si4OcD0fTXAzxhJiyFAaSf3
narDKo7VjUcvFAi8auEQC/N6sfgZgsvKj/ZG5F4po6Naj1IXjCUm0CdJe9Yl4sLd
N3l2QYcdZ19NwpSqwas1G/wkpIQ2ynctgs2RekKFmk86xCjvHVPdy80LJbtSiuC9
TsZq2UOdVE9P4p7qvt8p/NBDfUjPkHiDzkuDieDsOoHymezVnVzarpMwOia6fYlv
JZt9ZhUJpPylEgslq94oRkI4PQodvYy1H/Cz0NYbM8SWskE+HV6cN7vx6E0t2ZlS
rKdx3gs5VKezL5KB/177j4VfsqLM67xK2P8asKkH+9RLWE3jYn76/fi6LjuotMG7
rcICP6TvvXOsD6ZHn76TCB+700Aq2yJXNo4p9EcOjzIDgz0gSsitHdS3GJInT9YL
cJMdMQ/vmDirSBahIW/1r3TFd0Uehs8YLI2a8RTaTxvsw77Ejne9JKInyYfT7G+u
n4nX3xC7cTwsW3fX/gocmAIrBord7gPdpZX5G36fJ60c8GdbbYD/GkyTKNttFBbm
dnS0Eiw6B7t37pCGTDF7VrVLNsg0xXh/CDu1txQkkbWZsCnuKeNYZZleyrL3lYvB
pfgrXxoh7LlaPpWIc78t5qYxUVAJApBHuFsJcVWCTE27d38SyivmuHJ3XZUXMR6I
87LUa2LWnsdMLKsWnptneb1o9OIAa0wZbvSz4S+b2KdsJlQK0e52fVlBddfNKYyr
SWyUtMuxsRjEfe1g/en5MR0lwVBR7VtjC3FdhzkD0Tm8HYIYxFwl2348Q4ZZJIr8
BqAbZkiFevz6dofmgrx5W2YJIwEi6xQCy8jBdLOJ/dLHTnuwuHedegGQaBVYDQTc
b315np+rmXhHMJbVmSj5IPxYIvML/bpqTHmgEpqxo7nmejTBRHaaHiD4+pjR5k97
2G63HmSesfI3zkfZGEggBFL0cnUwaurOqzHC8OTqpQByDcEL2Aje6z5zfM9XUdC1
SmeO6FU8+uDVxIJhrnuD7i62WOpDH+nbZFmdTBF6sTD/pwyKgGapV4AWFbwnBQXY
YRuu+jc08sf+6V4aNk+YeUKvZQ1599yoB1G0EmlVJbrjodLSWYF1H0ZPvn8Nx+JG
DLNOHrez+O8B6dUf0wx6IS9wamMvXBbI0UMyLHIYOl3sZTYoTJu+WKDIlqGIBVEA
xri+6PaC6uLn7utwP/TfgN7OB/LXUe5e06v4hKCbbVnXjzpQa86WAsYb0/t4BWE5
MCvkZa1wgy289Yv9UUYEpy0oLFfn+SZ6gY6zk+YOa6nnXtUtrtcxcT7rcAu9boQA
9Wq43oRlQ+Se/Px21WyALFSHgO5q3tb6ZUdGLBLzYMBCAg28DXCfScJuDwt3BkNo
8kZbZEHvZWBWzP+uZaVIRGpO+kmYJxCDn9VHrelsXYs8GhDdaHb85zBnvyw6WSI6
dR647xhsOwfzLpcVL8d2Fn+SKIReQSGb+5lAoR2rpU+c/K3TLKGWUxbb7SOflqIx
zTEXWbfEh3WjVm+lIVoCiR0QQVwsUx8g2ohBkoMtbecfHI5is021X4jvMYF/n5J2
0qS3gHO6A+TYFw+uf0g3sBGtnTHFyZ/BxmEknSFxW9GCtgl7DkPpX8mDJKVOOh9m
5SoWxcMoiaxWpzPJnrmlDWniFj4CQLko1NaSh7TbFueKzfvTJWckeYmjKLuyS4Yl
84tdq8uaNbEeNXyMklScj0KmUqEoWsRP0+7CsOnngyR4AVOGgKVwMr2FkAm0OL+u
unO/HoKEWBMWMDGI+VTTb7Sj755YGnNHve7Z+EyLgddMbYoocb7AWQIrZy9CebVZ
Saof6JvHxwzsx8iAyCT9Q0zus8JTDvXmoeHnSjuqTwNYqT2XLjPPkxTRiRBDjYMe
y0VFt4h3KVsSqxPH2kSF+XIGj8DZg1TMEWBAVBcIPGyJ78y9twzsnEv2OJEsPY4W
v3/A2IMFLH01LnhYCPGt2Wx33MBGMfZ2fNZhU3oIC2n6a98F6mQfvSVoF7/ayU9c
YdOD7PDIk9no77URKPh3FOy0P1D5sccQ1wrz2FF3OLIg9qJ7uVOe7bdgPHs2+wZX
UT2Zf1XOtKsFjs8iAaoNw/0QFj9UuvrnX1L6PmEJHk+7YGIAJJOYkwAo0+W+AzMN
GJ7TXy7yr7hknpdH8dynAxJWNRwvMliXkhbSClUFbLkrTdAbPNRoX7sfPPu5Ovfb
BWbudpqRqMl9KxZv+IEMnhYzKj+zouVK04jJe3CEhPf5f10A/wQBgl5Nkzeqdpx9
4cg8Dnb7oEzWi3/dsV5Uz1qQMepg/7WjuyZ82PMUz2Vkb9L5P5G8gRZqZcQE0KDe
eFOciUrh6rgDvva5aagVEKbyg5sKWBtAKYGwy9btFnNkeRtXZCtcgSa6bUfAj4WZ
n5WWLQ2C2AYZUsrqg0pKPbTxUsZE00EVfJYEu45NgJ/s6gm5bUHJyFl/6yxm0vVl
/QvAKqqCU8WCpebq7tkErhSHI15ZkKt6LZ+Bwo5w++vlRIJoE0c6mVoibvEi0S7X
5PC+nRjMIHGyM55E1ODTjLl+5SMsWxbieyRW4jFx8P8xU4/jOwo+xTA2picojgO3
V0cjg+t12qWFPo3/JsP4EAnMPv8gbfcOlRu7TnpPbC+VkDMeBlmP4cauTkYqkhMk
Q26VBtzXYD5FbVa27gXwtRoIDwYhUd9G3wnwaiD4King9vX9A4mkKKa8ab3masny
vGctf8MmSzW9SN4Dcq6+ZbUPsfP0Yy8OYwFhbxUQtomwHkVMxZmtOaCUf5lcxWmL
AKwG/YUhb43FhTgkjBKgvJfOnIbmuxaMaFFLOM3jmCTZkjsLIN1Pn4xF5a3wboEr
LE98EalWrrzUfEY7tkZSID9wnEXI5Xgo9lNQG9Bz1LIhew/CmT+TYCX0HdwFKdiF
umHDDi8rU3PRHif5Wxxdq9CcKslycKSHyyuoqHcZdb2F2kGrXXBoewTlRv3rAc9o
e5aTv3klax8VTn1WX9DaSDxX7AqS4J4Y0hQJKA2Be1jU/SUmNpZpB1hBcl7Ztfa+
jP9apMNnlEFAUjJ9M8WlgXVq2LxLl4s3nDKPWaWXc3rTkCTyvQA13rIalL4qRuNY
ySyr85OKVBWqb0iIAy8jELxJZMuB1bfI/KLGwx383x4W2eBp507lc0JW2FIKc4tp
u8+uhtKDZDEWuXKaF5I8WDHELrJpwSLK///3KipxRn3uKSegXtOEZXMv4EAeH4Le
B6sujV5LLB7BrCkw+DTk4xX+T8sFgcTD/pI8LlbLVSvujnAO7YMbke2mJMGe+wFE
uXzQFK19fpUinShRDtU4yDMnyul2fNk6BVOLeIFmqTG+9SRDIG0Ao7H4HL7gRBq1
9lu+Iw4KV73xqY68lpbMTae8F2Zy1lqvzTYEk2ewkHfgZr+BkvWW2TL8/Ofp9MEd
782Kv1xXsEW3SiNswsISjHsH7958JiWA2t8XeSetqLCQAz0P8v6afMKquAwTRNBT
iwFqitpkdiFigcdJnqiV5VHFBrZXVx2xxUYUYWOLg5uASIqIjcnaYKcLsi8YOEF6
tslcH1yjiEJ/lRjKElyHJfUHvEPygyMZWQULlkk3etgfLid75c4XRa0u5dSTiV90
6XuolgjLLUsr1hGcdWxnSpwaXZuzgiun5LoxnGv8WE+7ifpo9L3QBHta18IsnWOh
JV3SFEGD8RjLrxtfeLx085O/jSXdVlbD6Wr/3N1B/Zl1INAAbfyfM9BXJRff+3L2
QGpXWPD1hwiALYBmDyEnr9bgZHQh/09Ze6xch0dLqqGc4V5EJQHS1qlamK6utt8z
r54egwIaL8TZ2Y5E7piYOctciqj9voUsN810WZaFpBLjNtxzFKVXCFk3OwD9HNIB
FhP8bpS5Nd0IWTI9n6jX7e77NRu+u1ceIz4FQzQr1Yzc9jA/QRy7yn6aCAGy13mf
jW4mMG/aO0sa+oQdAOMtLCfsASy13u3OKw2Y9Ct2RVUD1WMhMhgF+UHOyfiW87IQ
UG+7iwYsIVbJkQhdbLwhNWN7WWSE6zxHtKLlKCx+TD6lKwLJOl3lwS+m7+UYbD0w
aTBZBBwvPhZr7wlZv1jil7GhVYk28eEx9LTyBEDyU5JJZ6fSAUc49XTkPmeMqTP0
d7FORRKS9sFovoDBtOWNTU2bIMvTTmoG90MKCYRZGF3z7l3FghA+9/cs/+hFh31t
DP02HBzlZbVw3M/8FMNVLq1bXPiKFczOTjY+aeRGKkPGIvGu8uMTCEoXEn8nY0x5
78dxcXGQRbj9HXkbr+I11jrd+Dy/HMqJn2+l8T9ZdP2RTZskybui746bnrqdwcx8
4fodTPTBLKYkmKiGNzLrVcnbfyzARya/ImUcRadY3auoujBUNa3/SOa6T449qgmW
owavpphEYMr1Zn7ve88hsmSD2m0iLAoN96dKSWfzYlQemvkkdRNV1OgQvd/rVhna
10UZvHWsTF2up01vsS7K0tPQdtWd89/zAvBrJ1iIgz4tMRik+0Q/8GdNh+tuq1bL
EduidY3uaegEX6n1zqGuHHJSXRCmRE8PnkiIUwmXg0hsyCNUXLEDH1rT2Cw8jGo9
dI+nFW4NZAMdyUJsxxz9mnV8sWuLygBAq9F6wVQryqy420ArTd3TWIl740thEm6J
i/Nhhk9d1JyscdG8OzSLa5WmYFk8vkqlA9QA59O+WvyGEuOSRd5+K0L63MiKUQdg
ZCd0yiu2bYHW06+B4DlPoSy76e2HpIJD4yFg2JWdsbNodxWTBdcvPrYLHQ7PG/YL
gv6aYzPmZzOZlM+71IDJgqgsvjNlq+b/h3wITGUcRaUFcx9OzL12Rngf7KWSuQnq
eQMNSOQzIZ/JL8pTbtQgzDi3S6ZIKSuTfwmJJ0iCYp6KnoU6uZGiw8/gjc91e1bs
1X9LfJzR9T/6aFzpQz8z6jFScbeWnqMq7qZ7zRTfz4qOQhaHdwwgGNy4bEydoPa2
WcZsAGJ83/BE8IJ/xGYclm4PjRuCJvYjcLL2+NcFJCWUfvSmM3iUZ1jSQ45CAy8k
Ibwfm9EPX8ePH4EQPKDT6UAzoC2gcHAr9cBNZMLjL13ElHvZSbDKX0BtbEFAZi4D
MH7Oa4BGmJZe5NCA2DuGs+XdDwdI3rF15ZVDrzuUTCsWOfAlsXXOP2qJqoDPML1o
hPRJ/+nPk8y1L/M5y8KbrcdEaohKYZZxlxmYd/VnX7bXqfpSAZ69VtobI96yvcOE
nNUN1RMjgT+3jGa6+GwvQyilwc8aR8un7PAM0DQ648agCj1rCM8/bg5zpU0L8v1z
8sYUIY25bjGoodXToHMTm585D//Qu3s5PxCZCQ+VzVFNWvsJJa/OLzOurPAavRjU
lUk/h165b+yV7YymllzsLAUXbZdu8RMzA5iw9zXsp26i+i/uN/gQMxu0MjXisJF8
JpuOaj6urPujWmTbQjFzXfXhy4UKL8c7qXhF93g0OKO2a1Cwk1VQwKzmX60nq5Jf
5VO5TklPzNNkhXRGiQlMaLieVdyDRNsCGh9edIoSUvxuPDthI49N+SlF+cdwJ0Ax
FagXlNAJeLnwMkFOipmDt92EoymFMgYz+AeGDWMjEWHnEiLJfJsLXl9QNqo8ymSl
jxcC4/uEGV8ITQ2X8VFiRmaSUXvfjHQRZlaa64MgY1sTdswR1U4WcSEzBig/hN/o
u73J3YHcdd/fGPGTAb+/t7mxkuwGa6/qDJMHo7e70iXIaPs0fFGYay6/uIv9bRhQ
0V9JDyWJfgWo4c9G0ymD1LkjgR16wHbXPqPfzoSlR5RXnyqfHdZha5xUw/3gZzhT
6wYYikQPE52NaEf5gBE+L2E9iHktvDwrYyA948sUQM9fmgplz1ZgfAmYPtJESFe7
s9SvWRq5hwjw7Taz/jHjIB+hy0/WTl8oanbtTUXbHS2pub+tcF+n9wILEuxopihO
w1W8cKJ35bGc7PhDyfnzULDqiT0g7B3uadltAKpmLUMYeLABJ8fKn+fVf0I9W76j
YTc9RdS47fCPIHiOvq3u7eJlavAQVak/P8BvTHneSMBM8dPfwRnU1RLCgpyN0QfK
JmQ9Vxde5SdfZ+cDbPQ69tIRw4sLnvv2vUK7fqXOa3GCMgikoruu505DE214wT24
GrFcnl0MVe6uqywKHWa7Z4XKxBtQNEOfHdYnJd0oYibNphHDCKIFOwfYiQx38J+8
w+UzxAOTL4UhA6nJxtmITptA422TwZa54MYWrTS6a5VjIbgL8JphuXllQB35FwAz
LPo+I2FtTOs5WaPsglbMKa5TUeDjNp66mJIWg88t9dlNgo0bQSbyeYZuPxIgndcZ
4UO4o9AiWihrCWQJru2P96t1EDZ5O8VvtFcmG6hHEA0NjGPTWf0KnrYIlKqnRZyV
hxlEm/YYd7Imk8ItpgDCjuKviUtIOJVkhSgNkwOyPkHXhBx+SiY99TIipipJxjEB
4Kw+WEumKZePlRwvlc7c0FRtPV9Jt9pMxNuJ6lPqOZEPCPVmByOdyV/vNbpGeblj
EBxRaPkfqaxiEbhQz5BjsMnfxIxqpWUXiCazhcw0PPH3F0JAi1YFiDHHW9R/qIze
ta+koXjrqYSb4MhjsMYSTTNcpUohuKbkA2b57nkM5+CR786HCdsJb0u09JwBClUB
OExoIir8ICf6pHKdn/nGu2z87T+QGpc0WCb0vz+b4j1k56iN+JxoHxWF2T0VF0UO
vc5OrWSRPSOZ3HYypspXK0bWMy3UiwY0iCv+841cdZ3m+QC3HKEfWRmLptfD4lBM
2acVQuxtVYlOtJDmDFFAaeC1+xQ32IVVNxmi6UD+CyQ8qZ0L/Cv5YocG9svNan9f
vWgL8+7VA+3Id1pSNoWDeRfeUvGXFSd6Ast+o5RqOLQiC5Em3EjHD7LbQEVswKCT
M0+DQ7EflHV1S7PtlHrWQjIAiKTrTUqAZOg9mhx3Gk1q2BqzsS16n3L9jBKHRCUy
kZL1QF6rBMflZra8UQv1mICp0ldyLWmpNPuJyXqSMHgPR0ZKs5nragi0UP/POsW+
zZd7WoQD9epzbGbPDupiLdMJgPQnm0iTgE7kndfeC1iEB/aA/EU6trohBEsRw3Qn
RwmMxGpna/D+MRuw9r0YUbH2nbpWp3lFTYcgCtuNWltly77LXdeni7hIS8bEfDhm
Gk3h4tTTCnIxNTF9XuW4xaZW7uoS/C2WocBv9Fxi/uPG/fNu901/nplZDO5mKMHL
yRAoFOpKliN13VLtH9asp/l5kjzBS7kmzfjL/G+OVlQ4Ab42I5/J+O/O+GwFbzhT
4Pw8tGvbFaIlctI9BPWB0gAohrqn2/wfcxZ3lcHkREeFDR/kF2I1slexGKceH7H/
W+v90o2Lr7+KJBqpzdL92WqS2wBpcQf6sa98hVzUkkibYnZ85oF5s720wo0DX+JY
wVImTGMtxybUN60hon2y6pWsyt6jVC82MSrUnMBCKT/hSgDO87obWaVY/sdGHM5d
L/0QqId/WHwztBR98mKrBExvZWUwQ04FIxTWHdjeI7FGMR2ngD4cH12+iSWrjtmN
K4DFxz2lzGNYQby+S/UYyoHr4CGpgRntGCFCOmqUZIiZItRNJrHJOO6TATyGcbMo
bqA7IEi35GXO6EIiI+yC18IgX7RCwvMUHr7DaU68PQ75KpyP0kxKFtOk2DztdJkg
sn/VEEl+41bpUPStc5NOFbDTmUoYwWEBdsf32oseTR7uMA2CIa0ncRxyO99Vl5RA
nXA7HLrgMowPSQWN8eGn90toQOqQ9zs7DiTaAT7Q/gTfgxbSJtY4sb2A7zRcCv1R
Yuku2B1Vi3wlab5SfuKc01Du/llspMT0Qq7kzYspg9u35VNlISltAS4y8UcH2DTk
amf/c4GcxXstT1khqCgLnpVpIN326uUNog3y/Wpg7L9Uwe9FlSXRF4emOJ+ZMhkf
aHxYtFWmNxHqTYRE8mbUBSkuAAG5c7j/g6Ouioq3CeyfN/LgL5e1sWuFDJhXrn+E
sSWvCBzPhjVai5VLFFGBZDECeDS1YAjlqFeD1ob94LOfRTzCHa1t4bAp0caD3Plk
UGBA+y7kdnVAJ1c9F+dtDHO1hkqr3iJaOdzb2GgIjW0Mkn8qGpVmZz+voq+zYqRO
SbokSOCRmOKqaSUhAs5BR4KyxQmDmQWBTNt5YtcBKH6ztyvbugOLZfYratX4oGa6
NJaZAUa4m9t/lILcUnYcRlqMQsQrFPTo0aT+6hCY86yeia54jlBHHtMfw05hGpz0
fvpVQRfqUBRnwOyt73kwKEtif1drrPNM7Qg4Gndj+J8TU0XsVvKpK9VsP0kENoDn
iqOgMiz25q832XWUwemXrrRukEd8r6TWKQ4hVuzkin2isNi26SIMLzB9Lz6G9E+r
Ufue/BNn5epFJrG/AtYrVGg6izfiZJg/xdrMdzHIvyACqJwMOJDgFgrenLmHA5pH
YS5RPV1EpfLVx0c2oVIdIrMIdAax/dHyktIwo0gO7pCr8L8wHY5imf5/gU8qjaI5
JW9Gh9KDFCtvR0uhDrHF/2zizBHGKy3oToG4Exl5a7hnc2OCIEGEMDhgVZGSWsgS
zaTsD5zKxNHBBQogbiy3ZExboa4AzXh0qoTPoRPpppwEAwdyJGFd6hFi7emeW9Zx
0W7HffmNu2hzGrv73OszFWNDCZvAxpd4t+2MJr+1Z744FDXht2vzv8VVEdMj6u4k
ZND9TwGD5NcyRIWjDyjXyR3cesow2lEUxRdme70mECE0bBY3Q3nEt5XlP6unVxoy
ZI02g5obkVO+UToowHXnLk5CLnDF/rXXdZ4Oze9E2steBFFWEtkpC6DVhIah3pQR
lyyLi7LjHOwicu25jX2ZpSPb2v8bIepWWyPGLB8AcNTMq8qsA+4aF0Tt45coEGRA
xRh2JWOJBRQaDaaJmyTkVw41E5XthOQGuAaoVcWmo/dCTY9u192z+Gn+IRwNiyqH
40R3tczqBBMfRQG1E8SyggnZCiUznK6gC7fx/iahQiljS02MKTUnd2fdtEQS7tTr
qHV5I7lHSiml8imuWfcqwrB/9z2lLcbm94qXwgT2WRwbHgczVCnoM/UNcv38VyWt
9GD5m3RlX+irLoLIhu7Ac1ENkW6wmE90c2UaE3fxdqhJ17GUoJYRq3B0uBYc6bhQ
1hKqkglxushWjocv/mZFgKMolAczYR8bp7AAI3mZ1Lax8rA8yL7N7LgRtiq32YA+
ph4p0Ap9fVV8GDEgE3z3I8ZLe71eT/4bgYD13PRspyZcH1t6OtLyaAN1cBhmywLv
ySBSXj6oLVceb8v0Xq6WgFkbSPv3CxkD08CCke15V4amuGgThqdKOKsRhWJLfZrH
hzuo4z+IYgr5RP99Yb9PsyoSQPz18ya3NVpV9idhZNBxiIpnOiDLvCyDglTCc6Ao
9rzIPb8ewrxc9Uyh0i3lTUE07jOx89YVaBvHsmvDYBSZpMi4XVKiVVJHKsEpn52C
Iw4PxuuxUCMrL0H8QzbT8J2pDEEgMHNRKpY2jReldir07+u5Nw/KVzWcT3ZGRytP
4AabsSiPWrYR37tnYegzSvp5ZOyRVtxToIfGQbDruzQKkqzoIkfeyp1GwkiHQvoz
Xpgok+QWMYyUz9SRdcG5p6HfgR60Iew1ZU/C5EDAkGIzu0aPsVhN6sbEOu17LiwI
ArW82h6KEG51lCji9WBK37SF5GdDtUAABsCFAttKRFcbOqA6PL6Il06ZaspDyXYD
ixcjpFLl/Tm05kBoVdDnpyZCagz7qNgE7ZqXKj2XOU5E6m3SbE7SLLB4W9WpFnwG
tNs584lBdQJXTOYpxVooCU2zhGivcWw1n/5haiNfFlf4ZGt0e2W8CiEJOo7ffXLJ
www7RErVtDyy78O+jdFIvn2NSDsYh9dG8VdoNvXSg/2I7PTff4f6oCsgbdrmx7Dp
TiNF0Qdz9lSyjuZtRsPCPd5vt1EAYkP9Akvrd80/M9OUhPkqOYGlIZg+gaiFZV0h
uPzNUrgEVha6toNYv9kP5AV+UDcWdyvz9dFXqkdvKqZnTqUSJEPtglt2yekLD0IU
WeRf15NV/GZJ3GAz4TIzH5REJ1xEMJsDuJGoGaRyYnXFdkljIofZzE+rj5cSURRU
5mBYQ24RCBcfF8cWYvE4eqFPc9yPSMDWUGoxIePXrdTICic2F+ukQFAlaieymOUM
nxg7ws58pSJDQzn+LyVyuOWdOwNhkaoDnoEsMn+kCf2HHCBHhYkSes9HfYdFNrzh
Zm9ciym3/gHq570UGrIjo+/vOwEIITKSeSM2Za/9IAedXgXgXqk41IqyFvTuxw7q
/5C4Plb3YaUXIaeaIICm7tgBWShovQR4Cbr5xfNxgClhSk2q0ls8keRkrlohYzao
eQWsCYCBMaNixkFnp1J5zxuDxj2E4ZAdvY20tOpftGgJJ8IYsroZ4kZIOHxw71Fm
UEaEmMb/14hob9HowLg/T3uUkiNF1FJQX3nLmyufH8e3hdicn1H3kyE47U6rMszo
KxgoukqxJg60Uy/Sj/spQNqEK7qt+WsjNHziVxmdN65GFwm/UfmZojhIiAkQWWkt
JfAzG2nf/ahe076CD1nzoKyoRQoklb631sKMegnfC7Uae7nd1KWLe75tHHp8MCtY
ZnScO153B5FtY5aCe3cwPvfNHVGH8kL0LLNnqbSqVGFm1jRs8lMRy7QhluchHCoE
nZYlYlOlcZui6eYIxEoXNzxQ1g14bvsc/I38D49/9FT571Hf11onILPr9uCX0wcQ
tCp1fJhhOUEBm3kdVwK13Gs45uznDJp9Ddo4sxSEwDH0fb7M/C/jQ32+msZYT5C3
5i2ipqq+XFoVPtiUKcHtR8ViBSeiRfk1ijesSLfAQPNkYM7fEVNuEXxI8+JPv19v
MUNRoggXNxfY4q9K6dX5aK+jpcFqrMKasv1531HBjbIssJioQiD6I3gbDIrEFZKE
/2+zPJB+l0Imb9o+IDjZCCzSNVlnaM9ue8LvNRTze9XqWKovHpXVPZr9qWoNQw1U
eV7tlV8E9CV2XYYveOvBpAGHqDwngzXgimLwZZ9FaEaILkIqB4wEX6Sfa17qibTh
NQf8U6wvUOSrKtvWE2VGYxufU+8V840gsH+vuF5TJdVDjlGizIW11FHC00bts04k
ezOCmaDtthvwdOeRJq4E1e8a5nQmPDGcaI7TRVJg5iX4ce1n5zrk8c8AiGnsVaYh
dKLz5xOV3N1gP20yjjqk666aL6yrBZP+COceV08d9aLd68gvxzJBsbds3NMwqafi
HhMNmn+dl+waBVTBokPNtnVW/wfVJ6Uhb9I6R+4sYGZRaNZh/SDbSLwtgs+yrflD
tmAJ5WDLB6Cpqb09UH01TSaVVv57sV5sMQE6EZB78TDvz3Y9soqtTQTx5OXOMi2D
QqGTNO4MZTKXsz42eT7XZkMZh9E21pq7i5VKhuDxTmK3aeGmD3+HTFav/DxJznGx
ciWIcaCP0LunI7dxlBEgOCOHx1keZ4fik/mD17HHPeqGr/eKKnzZYB02RIOzTxys
5oOgPAkt5bZ3I65+X7zkRETq5TNHfD4g7DYnb/ih+x76cwj++7nmGf7q1bJWAWgu
x2G3lCin3yc05hHLtt0VhLyvUZnfVIVg8LJNIrJb0DW4c31GtsL1nNXV8YD+U/IY
h8TszZlb43rv+yUvtwNmLrfIV6andnOo3b3Pctj0JidWjegv8j3gf6u+qK44oJYN
0gmUp9126aaR2utR4cBxNa0XA8T3KCz922N3QxKesbPlGZ0R5mGBsOLtnb8ojK3w
pzIyE2sywxi9TDfT5tuHX6uJV7FUWbtxIWv+7OQzISY6uwnBXuSJpljmhfhw+qZ9
R4bIB9LgyzY4O/1bMsThNGLYbqqHvZI496Plll0syn6+yHaI41psRemJFisI3lUH
rQVKgdzhfpEMaCYK0bCIJbwFXneZ6KJkTazvLQIiVXQtM9awrVTxHqowQh0K9cJs
lh2Yda2nyPXGlkP25Cv1cVS+kAhhAxAL5QGlmtW8FsfHYNeEJo2b5rziD5vqR5K3
SX3BFv4BNOKRIgHNv7tkoRm8807Bh70KN24pbt46zVgqU6vESxv9NvVwU2KwaEzO
e7ceEb3MD/hlK9wPr+ngJ8zqJ67kSAPDxRO9ZPieIZ9TNhfoblOnv7ytt5VWnrf0
vtcXFdw/yTX9APehGsfxvoTmXAUpkhgpM4w6pLyLLoeXyX6SFBK+d2ddLsOSxqVO
vIHjJHNrMvJR3U1HCCI6sqFFXgMZOFBKm8DXs+gvyQRMrXYXpeiJs+L6lhlULga2
VPCjKbfJSGBkDoM78uKujKv970oCN6BvpbSMIoCwhNjFDAkee7pQR1lkCmm/rmHC
Wsuth0WjebZVCVK1juOe9sVcRR9lX9hkhxZDmDAFAbbdGy+I5q7DvuTITw6xr+Vu
DbW2atpItQLtmPXUrNKi+ZXCc5huO2eUnbc4ymN1vFFj1pgi6B1X8t9cUb+voE1+
cwCb21irz8AAJD/01YJtMcm0UyVHOblAWYBMXTqGHjuQsI11ZkgHWistkKRPH1ea
Zv4/GIpoDSFKMFzpyRIjsAQDJFWBh0fTN6Sk84bGUDn5PLW/OB2sImWyzjtfM89u
eISU1H876S+McxXBbK+tKPJkBXLbDC20VFilhLURWSn18yh6nyKuk8oGkK2qxalt
pVQQlvEI3OhlExO9BGoBnwiBOvLP7kUm2KW8ImtdbmSwAKL6kpKRqGfyF07fnTfG
+NcNmm8D3f/DRD9VBWRV1SCgSKe6krkv/s5BrGClME2H7fiVmmHKVB573pHQgWHt
Kx+1QXH/oZZjIrXkqzNQZgkamAHKFLN089Y2zOs7brelohwX0+1LtRyRKOJ8VltD
aOHEhd3zioTtyXNElfpdd008zmCX4MqmF/Y2csErNAMyIzdSSl8q069erbghYFGC
YLVGW+Oaz1dXOgtG/I6qa3fJB1HPxW3cBQVVwIxaOlWIKozfKmEAEg13ID7md84o
G4hggdFnmQgh0M2RCHsp3HqhfsEkh+AC+Y1yiR/Z9JSZ/6ccmUBfzPGhABQhx/vv
uZB0iLzaydSejCGV0HFulEBRbqP+ApUq2x8jeUW5xcw9Lu6FZa2N/ipKW/6PFdUX
RQLpt8TFPsmMTwgT9tDQCCp5JjeBbMCiSi1shuV+RzzUS6YEewjMCZ+RgxyC81rh
vFP2qIkpb7Zf2YhMEDn5+TtFnee4OGGzbNxy97PArWBW/TOPDtamnmo2GY5w9AcG
SrOqLdEUj9a1Rxx7dVMepfPm5DETIC+HCRfCQu/gazyuG9YAPaNbt/2WB/ZRDkmZ
uRG864O0dNOB547f3mmgFf+5fXLQJnVdehIyBuszZ3REAJAo4d25xm3BaoaDOV1m
bKYjvPCJ7YxHMAruej+jXzgQVRGc8r/nuQ7SC9YAEk8pxIu3gt+8niFO/3DThhbo
5A+j7f+hLZnYDSYNgHdj5lFfvOX3O73JmflZf5A2++2ji5jrj6qp5lMqUyWD7WXx
9rlSFojtCAMaC4vIzKlXoR8aW6xkGgg8+0mXM1wKPJaCw7vHO7Wk7jqe9vmZCqHe
xDSlUUXNzJrGFXmUA63dX78yjoUl2+9W0hwLiZavdfHwTOG2E/3h2/RNFGDnJXXr
IBnRjaSXo9BhcWUpAL5bNTLRFzHjyuAW4/YgOrmMlrCoS/uzq0NBkKZ88hnkbh7D
cxi3fuqGNtR/k/6UClGOgjCfBdZZPD9RgUOF5wnof9Eu0FFD5osy84N3LT6q4Gpe
98wX9z06bswLcQErjLU1mOa0qAwa8rn83Hq8sOtGnrfswSmXMHPu2pRK4B7Tolkk
4hncObqXWRHqZasEBq1pZBaqqMTMl0CbJf+Y/7p8JcR3ZNsttt9L+Jt2xQlF/HWx
JoJNb8/zPjPkJgV74wMo5hL7G1U1ePoiSjJhfT2YL1U3q4YkX7ZY5fTewarBZArJ
4tDZp/X5VI4hyGxBSN/26cVukgGXWjSooRynByWFHjL0pSjqi8fWSc1R4KGz2rQj
T0cwvU8OJQtFwudEuOM5wMoTJOKXzvVvOpyXm5C2jQnUm84uLAgmQiTuRlLP3fBy
mG7Uz+BIHax1+JHCZnokKZVgQBwyo0C7+noCyclqwNUci6Wzm9xP/keTXSvkPbur
peVyMo1i8MkmR39Oo1THIo8HkJA/21s+GWhUw/vLikHGifi2mq3xPCXC6ZEfpkw2
qH5mPKDq3tp7TKssYfHf7/a2cbKFkImVylJvb7UrAKQ2nOobepMT0Gtrqi96Q7mF
AyD7MYeQ59KDctKLtDhGkVZQdI5k8lm3qVHJ2211qRxHybp6uySB/eCqhRhCfyTl
acr/80NaM9ijsgWv04AzAJaR0HRMYcCau/7gxLsoPVlJ1THE2NL4+gImgpOc1vAG
LW/LpOVsv2edAeHaHLqcFjA7uJ1fyTvpksLiH4D7Uj80ft3PhhCG+UkG5gdUW6T+
Uva5hry8/oIJfGrZRC4d4C7zoLq2XXLXhV72F1ZYls8MpURH9gufPcKXzVGv/+k6
EW/yBYjd08pnfy/Y5EeL4HxsfCP9Qryq0NNu1WMZKzllALNUvBXQH3uTjrXOzXD+
PUpDaoC7EzGm+Ysg9ph0TVHhcO8wDLC2fmzMwj/CeGzAIWJeBptBnJCB9xAapw6+
m5ijKMo7P3dqcfEy1V3sWRsQmK35+RPvGnGHc2Snec2qDWapbj7HD8u+dtBCF9/5
+J/yONLkPUUBGyW15d52TtYo50CzMeW6EKgPkGTbasYpODPuvkgf2JFbyedSnG+z
A5/i8lh4CDFj9ZltRFdWD3zz7imqDIJXEKW7z+ZLlsQ65HVe4hYoXsso/3YNryDv
vhLewmZjsxGBopZmI+6S3eH7ytc9Aqm6A/HMjsLQzSv0CXtb1cqMW+Gbu0UGiZyd
HtZ7SQ8NVHi4Mtkc3hU+ri8yniki1Xn/nzSuagmSNkBQO4BhG3lr5qoEj6I0z2la
PY6SKIwfwNr1mJ0H7T/xqpMKSg0Aeu0MD9pNMjRYuITPeNNtlm4CXx1CPLrr+PRM
KRAKQMzKT1BgJvreOHWNY9aZ9GY0yjhjJDMjAofvq9xp8lHRg3mYfH0unr59wrnc
LOtftsPHFaRKIH1A4X6zi0c2GNQrPReXQFzTLDGQlNlh52mdlTVoDc0l7Se6o/Bw
P/9VjnCm0J+MeIBshsAh9IcRMPjOyWbkOkVFUVc3+tiRA99y/JZ4jA3Uy5fu2IAy
EE/XeSCoCM4dZeQwLndJ2YtA+M6JGLZsKWuZZQR46EjuQgNou5PgAuOxZa96Outo
citeKWDDywCx9vHi3vSr7yx7HNGh680aM1KicsanZ0UmfuWEIvyAT3yNSb+kipPP
BbTeiJ5K2mD9q7iuyjCKdktFD2T1YiP3w7G5JSMzJpx5zARMlWChsuXLS0fVhHOr
eR3Yoa9Hid6ji1Z1JD3zz7rEiwtAYyYz+O27L/kQeh/YEwNOKXXRZYFWjxzteKmF
xA/qp6OJ/4YEtnT6+cVD8R5e24rbOXZXtfF03hgX9u5J7JsswVRrDFt2YYnAznfK
JATFrVS/XgjTQ905OPSCpgEsJqVT+Y5lgMJoXLOzRO1aOKpQw3f4if6ZhqAvtQam
0RkfTh7BDot07gXOkWTxDySXk/y2eg8v/5YBtvhm8nAuZVdbyt/4k5+Cb1yVs3E/
w5fjOrYACU8HS/79VNenZFwYj3WH4c2lws3ViEkKgoGnP3Xi9tZZyjMdbn0RBXZI
Lj4ppc5prTTCDH9SIyNqmtBmk/ORDov/2CwCi7hGtE/lTkgKqHQUqp2yuVB5u+Zj
mDf1IKc2F1jBGoefJpH4WUEjoWkfKgLZcqST1nAENXjx9DVp1e2nNZMzE9cNsoQ0
25S13O5xP0kITosv5mVw2bO/dbRhlHwwKA9/eNa4v0nnygirVl5d2+366CwGdQpT
WY+V3Z28ZjjV/Pjn2JogOz39Y1B/O4OhK2q8bgceyLfBPitbVGtZ2RLNroCEWmXc
baRKtrcYaBhn1kNPy2dzCdS7a8Z0FB+MKhoGEiXKsbRWnYyG+D7AucSawHO+AHt3
Nqo+0liMWKUubXv+ZRI3yjsAgQpIgFSV1kLrtxtn7LqemOp0reQtKRuFibTInT4K
/EyxXh3VE+xFu7HiCrlfz2ZZba71PsMzYQsYSWuDIqkzTH1YzzXwW0iFOHFoiL84
Rb5ow5eD/Swq6ru8V34rVbYpt5oUHBVORRUXvYF7ph/Oe1T6TlA1H+11rmxC20IZ
exdAyGJkAhz+d/dJMXXV8ejuIs5R5AmisvImmPgLkuirMSkOG1z2f5YcPyLYuL2I
k8CTM+kQDoMNatgocbLnN9C2p54hwBgw6rpEuWam4IzeT9yw3NNE/dGG0H/QmuKI
btNPPCWdD5BMRx57JKfPhP83rkQWo1dUiq+OKeXl8a+TVmtIte4y0+m/D8spI8QF
WyunQjwVbg5k7yD0wiUXubhZspaEgczqxdk+DvizRQ79Gfgfvt8crOhTKxH2dFxK
4ipF8DaVaf/FXNnPf9n3SCCxBfdOPmXMFr/FUOVOwGGbbdykpdaaHw7CFNNHkeu8
T6vAS5sRnwOiZhuFQ/0mwAmmVKA9EJPrE8KiWIx5NCn/Ol4FDQ7/lg29WugGfQrg
bqZWsr68sPy1Z2CxUFhKAh4zlXsrMu4O1VRU3rFrJk6e6xCYkcfORq734geK4zXF
KbZQnO1Jgd4nUD8sliNleq0aL/zBk1N7Td1V5XLvx7Qo9x+0xxyuTA02yEmH2/wD
u5m5v5rLHoYWH3/ZSG9YgFlXlERve1Gu3ICmdad0s327LWAYNhjgy9ypYP6K9wbL
kA4YVBrXvnHQRCHIOjd0RCwtBF++lnj4ZCtw5FVciTibnVzP41j9lH6Gg4Ult9ju
f9E/A24SCEn+8SUU9KKQPCdXjWTwyUYVQFAuXToSqk4i7kYiVpe/LUB64iRWgZj7
Vzhjp+lSTDxp/VVWSjFs3m95/DnJjsRmQNXmcbWm+MDgwOzRouZAq4FpCT4iPMvs
NyQZm3fLNCbIm5kZYsxdJRkdFsTuwEWx96VsiSbFJk/mTf7P7qterNTRyzbJLPl9
fOGRvZ3UtjUekPE6sBC//EBXTVI0z9EY42myMi7tcGHL4aDhWhWMU1dyUBzQCWC0
u2bRMBLsLC0RGikMq3HJnPB9baJqemhstEHYgT77uH9fQc3+OJW8frCq2qXYIwlt
MfRz//ggXgfwkiLowCddAHHtU6KdKH9JjESomTkHuaEmDajLx9t/ajL0LBL28FRa
20Z4CVzpq3JCEgS1fIyd7jErKHbdT6sjdd1EE+XjSuRQtzirpi6Iue6qrdkJk/Qi
l9BauVY+sWGnGHXJI1ahlN7nJVDZ0K7v2u5SqamN7BicXpYt5f26a/r49B17DA27
V4W0uQgDyP1ZY1GGbnIe0GhBh2Xus6q8SeTQ4I82RYL6ItySYS/b9LK4KrZj8zq1
AKctNTs/28535RRdRR9dntQDfRuvuxjgOJfjI/vUwhwfoukMlcgjCZegZBqpy28p
TPiiA6wI1EeCOJ/14vLImUtZ8URTD6A8Ry9W7tsGlyIBREutSP56s5KrSbJMuCKN
Db/DfhvUj5NLvnle/C0IdbVQ7qcp66IpQw5oH+ED6qSz/Bswqb4zPgUPTjdDi8EY
Zh/ggK867AdGqLfeiBaPRX7PNuyQU1mGdlEL+8mQGveykMRI+qQLtK/rjbBOOSeJ
FibXxI9zrjRWqnR5youKJVyRAjx5i5rqN52UsV3fpxpCt3gdsnPQgYGxfwQoxg5v
zKCfXPj+T7ehhb+PDj0ttBUjIon5ay50gPMj6yEwpTVbBstxFGZ1A5Bgy1xowTLs
pr52jk6ti+RqieTC8D+yDMjPKTqKfj/VYddNKMP9iVX4vy3LIwqZboqhbWoaIRQ/
F2PMNARy89HjZjylQ4l3z6MeOzsFLdBPK8kFxMYnzGjyFRwtuUYIGmppotV3/nE6
jDnDZEbBGmFwqEPefUtjVc2SsfsSXhD8L0Bo8oh6Cu/JH04eFgyJ2O6V5sfJgWvj
WF8SOMDUA2En+SQNnAcg86r8b+YOIf5a+3Q4nb207+iwqGdANH43g9M3zHj9YLe5
7E9O/LOijE9uPEoB+H2jVMkyHJhjmObfGm0byKM7vgKwZzSYRd++fugfjTmcS3n8
7TZUWZ5XOB/Z3pTqzrdJ3F6fXf+KQY0HhLDip1ngc/QBspmqjETGoVa9ysOa5oft
55WqWkWfCuofZp0k4SOsNTKfpWmjY5pTuzH7FA7AwdI1V/amcgHu/1BjH/ZE/bjD
aoI5194YiYezthgDkrUG9aSsy3M0R0+rxgUNFzthOd7EoVf/rWqp/uKhEIXcAQb8
o+DWUaXBCDRKblaX0RZJIyFXwzhZmqmNHRfTMW88tlVYcBW6cfp8cWPqZEwKFLVt
oESNxpXMtELWAtJQZBXLY93wFa04kGrdCJM2ZwIdQIxhveMaXmcUzM+tvcUIH5FN
sp4nPpGS3qHnHPXOjLoJssJ/JVDkLPSf1Ph3tLpS++exKbsRNeafZnbKWVfsIM6O
wUffxrmyrpTQqn8LAy2GbLdjvQbvU10/RnRYASQNv690YNXTPKPj7QQtxu8bU67a
DY9/vI/dhighEKIQ6E+gekRF1To3gjXFJddpAdgvgv/AtKrcXR+ZIWlKRrQ0Sbyf
7x6MXcq4+DDTXX+Che/ip3d950qND+ZxfEIeuCrcYVHxn9XHPA3eljUWp1W/zYeb
XIvTwftESPXGN/A2FrQLfnpDXCloRSD8XPUJUHcY457fBTbUbS9wafvNpHV8cXPm
bCRRx3i5115jLFxdYG6JeFizydqUb4PgSuf0tQYRleXmzM38tBRagB+ljCYtcSp0
oxktH225zZ3XI1EeL/3LGKkPdOOzizx/HTMTMXuY+CKBSCjVwtrfOyDp0S8F9AvS
7RxE2tPvlDSZqVlWbQPOmutlMmfBnE4zuSnDOB+R/Qtz1dDQySeVGJos0tRNnkxq
6mr9nXWsMmHchDw6dczJrrF7msL6A9MfTGWFv7iR1KrPjP73pzHv6qBK2b20WP89
WgvDUnrZd1sorP6pn8NTqzz16+ja3Qk5IWlbcHr5AqWrUfaTyu0BrpZBYSYp+22c
rJnmXOtg2iPlkiVVUByHLBt2nhNIVpUR/SFJ5q8lN5WictwHj+Y04U+cxgO6Ldfc
oIkCelY+Mt4ExggN1Cw0xHOgVmdBnKNJ/Hv9PBO+S4BVsQIvRsrLUdpb9cnecUQN
rtqFxqDwWxq06i7L+LxEdx4dwQlg7JpQpr+9XcS18ZlVHIr+VVYqawTML7I0PJS/
NXQYCYeicACL1yaA7yAayJIktf4O3y02DIUgAkeBrJ+4GY5zbIC0jrnYIDZxZCmj
vjKztCo+mZyv1HhfoOiy6pgOkMLntSQj4h3EDa2ZdGm5muySHKUR9jhqQ+kRAZoh
YdUqb4TIUFF4aOpHRrDcN62deyOkU4WktZkjbNZUmL0P//KJWZ2MK0V4EZJp7j9U
G+zAb1r+VsAYpr2UzCLuD0JuL5YCideJPYBjdp3CNbXdDN+CHsn7QAk+ffUIz3wk
hBzX9jeN5bz+BtM7pQUBmqQ8xL+vbTDGsnNuXtIobdJWCFTInkmynLMSq9XenhyZ
6BW7DqG+86+MNgBOfqS/Z14kGZ4i9Wnh8cBbXxePdzEMTRvV+Y/yQixINvSJOvvp
XovSxQHNLN+YXQBihrVRFGN5ZIMaSt6SOyEnwz4Bi2OtIFzUElBN6bPWEMXXsfFd
1tUww0uIIsnaYYObgU4s7EQqiDKxU4BL6wP/9HVD4rKcgybDIS8mJglgBYXkahRQ
M/ngQ4mAxqxqPS0RT7J1vt+cvgEXlbCezyVcN+GJqdVGlTWBAkhiX41XoyfbwqMp
s1N6Dy+Qxt9TZqWf++oPpT3JQZqRdp4tjHBeXD08UgCwi8GmdZ+1if2wNaOSP3CU
976ZOUv3zJiV9XsVuFLStZlnygpI3mPhrY+DA75yLJm6Z7u0lbhzhcTeneKCV/da
bgauc72W/o29gzvqFauiH0Z0uhNWCRaTmrkCZkJIu3yaHHyAwXDUVdbEiYDu0ADn
tmBaSAeevIEQ0/0NWju8EGowePyFkyDOGWbxRJdq2decUeKqJ6S5uPqx6YTgA7FH
0G4glxnHDxyHGl4pUMCVBfS0DuRfD85DwVdvmLOYeDLk11YybZwwxZcohS+56Xer
AE/VknRgEtG+Sh7MtJv/POsNt602fVXt9pe3ewSVRxOO/WajzJB+taISCFBW9e8X
Z0CsHLCfzthai+vY6uEiNGGggYhSd3rxFWczBq+jbSU6lRBjnUBt0mP36/I0UkDQ
OFR007406NaM3XyvAT/KOzRbVO0jwlkZw2UuEb6+bhQVAOGkkb0Sw9iXLIukI7q0
9iUXOdOg/tEMBOh2CLYCaXEJ8aEloIJZeng2GeEah3NXduRET7T1IUI0444OJm3X
+6yeS3MgxCYRMGi5RzoKCnFc62ek7/HlWevrjDqPM2FNpOj9wQszd0OEsq3wNvd5
y3+gMvqrITT5avnaPzzDPfk8JTwnxr6IIFh/UVUVfd9S95Ee+35yyYHR5w0w2Ibj
r8F9ov8S4LEarnj9ceu0jXJHfJszqjwzYnAIm9OhQJiYcNYTZ+2HmiAI/oIyS1xG
RfjHYIujKYDQVycYSB1ov1RIPrzUTxs99QVvw/02IW4+/UNR/CjbLK48SPrCTzXD
JbbwCOh1AJeG99de+/n0w1D1RIDS4N+0vyptbNdDz3ScsoE/GLPaoz2KKm8fTbim
OFjRFb+7U4ziG+y8o+ID6tKQdJQTbb6gsZEzmiYesdY4NZ49NR/bc2h9iQMjYtFs
4g0TnvVc7Yy0RHlhDWbRY43cxBDh5hEejQTAHm1axFxabT4tnMfgUAl78zZJk7PQ
AobaGpv53uwnPKyy2b0veAU1GnMvZ9yS63+KhKC+iaAOu1PcVLRJaoNUMUPUbhgf
lRUVuI5gNtSrGJV7S5GVLcDkRGrBKj/3mKgNs/fQuGDP1EFy7d0So25uzsxKm0EU
ZlOexX9NmlbWvmengyY+qdBzjSdsqcqjcrLJmwBO8BdqRZl23SBHNrInTv12Mdab
Bi74kDpm8hIm1UooVlW5B8l0KiW6zleCwpvoAmRiHs1z3cGukXQCKHjj+08TSlul
2e5vrOf5fWGc0t3Kq7nEvhdUOFXmM5JnrGArZTyzEtxkzn9mdHH3vXQk2IpB9MKF
LYWx4NbiQsU4Ctlq0FvVZLP19M8rzgd0rTTJu3a9ffUXnv5C/qTT1LTM2AXWZuDE
VQw5Kf9ghroZMOJgahA0NmJzRoJRb0dOP1xhCSYozTEigosu9g8ZLZluyIOnoWh8
EMd88G+1HXfSbH4vzvENOxPPxqMcB+hW4okwlPE1lGVhRFqdaRNY8D9iUaGl2tjQ
5jgBfYLyjoEf5qKvmqza4RW0qJo6Q9Dkkg5ga3ErGJ0x+T8N6PEXr9CoHCV70nzh
ub1ddUOnoxPt/3bRBmel/0CitzPdBzBerKctKm78w131wtRAppqHJsF/2a8tJxR3
9GkjCT+Oaje47fbwDY8PRGViDBV4dcnEfIl6Rx+dY5+jvKku8FOsS/mzS58FbFbW
xIJOynRXhM/dmUOnCI2PCXszWuBsDgg75Ud8i2KvaB4ngfsEnteAS0L6VtSHLv1A
Ni1UN2Q2pYIDaSAqhTqVfwNDlYHxM/ksqCMVUnd6MEWM9zAqtbTLjgpFANIJYZSD
aueG6C3pc4SDn8ZOYwbee+1xiOKMwbiImQRxk9J9MJCtorCisE6KBV9RF/cWzafq
Z/dp2mQsxWfSswZJX5SONaABbmp1OeHmC8Odoh4cQwVWHknyX1RReA5v9oPNWJVX
uiTCRiAexj39+zBCo/eGS1uXvlgZPh+2Ba1+LkskkogG/jU0QoSZ9p2/zWCagc2a
pqzVtCDmpKL/hnNZWnojuYJRrL/D2K7W9KpsLITDGxZnzeU2ezgvn93uVK7K6mMg
ozkgQfQHUQP+wUh764Dtz3MMZhU8Gnknk8Ldj65STwBlJiBxF8JxIoizqFm4LXnz
w2q+lI9EqMkczsKS1+MtUBzH2/RWt6vfcSZJcGWDMyNmXCmzM0V3wk1TXNhqxAR0
JnKx2xJ7+fUpxtENETYopijQtd8ULLyl3nE76fYCVmBfTROp9QHJUxCxeIL58G9K
Nss6s+pu/qjvz7v42HZkKCIPLup+P6nG0vLRo+OySOjI7AzJNGedXxRfzsTGUrq6
cvDcqZmITensz020ON05UjL0cXbSNLmwaEuN5zq8K5e08N3BwDakze4Rt5thkkBc
0C/ZHVGOTUR/JgqiGAyPg73E8yA8BK9OzAMUabtzINVtg8MvPYf+x4qt+is9DUn5
NpLVC/941Z5CfwstZV/Nv7fcluJ9NT+lmbmMIcBa71ct5IFKHjNDFjBjAQVEhN3W
5ZCLpIzrz4eHHwco5kuq606b5R8b0AkS3Qs2TE9Xf/W5cjH6PukKquTkvqVu4Y6J
4vflHO32JkICpAl8VorW8YBWgLz2n8l51pABr84xeUDrrEM/UgBh2AP5U0GP9HGN
SrVuHz2o77HqKbso0GZqQtIM0uWXeMra0F8+hdVVcI1FuZgpyHxKcHRonM76n2u+
2ORcT2BhPoljFCO+esmCGViWK4HVvUM9qnN1QdhGwxVOAqpdtKVtqfyc1vxjJ82m
MHzGT+9+BvFpb3FjaCWZLwQikid8ValG1/ew8+sQiGdxij9eS8ckSQrHSN947VPC
AqDBc2y+gCP+HoVT0Tmb0y4f62KKt0A+h/wiFmJ7cD8OnRnNNn7ayFJc9NK6g/Mm
BIQix0odmB+7Lc6b9nfkN2HMwGzSS9AkZCRTyRkG+CGz3FfRA0r9AirnzCnKfyZ4
qn2Z2zH9bx0bsogNkggwc/aKhFZIHeWgxRSEHK0//NmuQEpvwr8he4sfmKnJM6Mg
1tQ2tQKGFIGla3qfOKbZ50hgFLxupWQGOBd+viL+3kl2GOaR52BwaAFpA31MaKTw
npbeAZXHZtVdlkvF7xTpFKI4h2uhU5g450/9rEDDvAVaDu/oK6VNtvppI3556C82
bBXmDwEVGlwqtJkHHDM0PXvC08k7XsFo1oaQxg8WKDdKnTTg7dBkygqhNIXnfaEw
YlM6BKgCG7BkAnZtp1+VL3HPwzeCzCwWgO0CtN9eZwhI7maF0CeULufw3HUHQMJk
bcPgiYgXMpvZMIRAs4E/EDf5OI3Ytc0ZxhpWwTheaVNG7RLA0HSfllf4yK4nCbrj
FMIqtiygnnV9+xGEUr4SYNNNamTkUNZTLqbH4a2BI7PnuTofzG5yLslfmLG/xgSj
dhl4lNsBCeNibBb+u4pXB17HRjefUO6ch+bp8Qm2KqYY79jhmDGetGKbhO2DE/O5
c7sP9KYFE0HKWzFVgxItGyrhTWJUkqej6A3WN++m3SzmZJjPYc66Zi/f0Xwy4bJ8
K5DiIsmq4yFIqU/AUXFlWEi+IQzA7PfacZ79yo7P/sO/QQRDlwanY32jTOyFot/L
yuSTxVxrToFqR4sZBa4VC6vzFvh0NTACG6RYmi0Pi4bpwpkNOe4zS6M7Rfk+QiTv
OHDFGlJHjR4G1vT7r5xXKU24NzhM3y7lUSNNqNHtPMDrx/npN1APanfZsrOHyk6O
FArKtVrU9l+DXMULt6bH/uXKOJijQPsHwpz+YU661EilmGayfAVfa745o5ju3IJ7
3C8vdn/gj3Euf/oUie5cdkoLZxFbIfVgBdLHKblCDU2elozJ5Lr9/cpENkpLwuxe
UTUKRWo2qiZ/qvIjyH5mc0rhLx/jOGbF5FddkbKsQfEeT+9O51pTcioeKqtO6zCd
0kfg5zUG6j1qtjPnX8XbIWZUzSP2NHnMSCQYC/7o5xrdGbKY7zTweh9dkt27kHos
s6bYLVTIVz7zkn8xAG37r5vkICQrsqrun31li8sg/9///MWZW+SSwe9neRft9hOc
BUWu2yHdHJ2qPHqvzP6lAx0lEZVRl85DXJ49e8YK8x4iIOWt1znVq/KboQYVo0sC
s4EXxB/jqJ9CBfDVVA/V935yF49pn73TFMBjYh4BkcVdQZpdnAfD6yuz0KpO7ro1
SeuC+0anFpPbUnbHImcNtfM1npWmJAEWn2zB7IQG1Sx6GX/CqXnMpdm5eg8u0pjb
o3Rh5I864Z8qK5t32VLXsafmz64jjeZhp4zTT/8QXlzbYk1CW7bSFFxEVPuYJbHg
0aKHlXgRBYc+WfWdu5g6tOnOyNGSCjqpcwHpUGfP1XHX30h1JF0UCPCHmqRiSc4e
73EO8KBeB6SWeAWTKkX61DMa4QVwqIBZKCapGzzlVL+WvlTJC8j2iMntQb0YwKEv
KAD/WSWs8XdXYP4/QS+zoj5Tlqn/RPiZwsAz0fi8c5YBCStpgFiSm/dPpDxYx+dG
UQTjJEvXMaQlJFKMtkj8neZaHIjMCeL/vDIxp57cTj4+AzWvIBGrWwerMKzjspRm
NZQiC8Hk+cRiqj3VnK1PjyWIhDkGMW2wVW52PIdLq1Jjkgh5GSdoJvW/y87yAli3
ejPfoLIfIm7A1+CdzHxpM0zpH0GVRhoiZh9w6pnxMLa7X1wqE7QuhKrHNXpjAzNb
oMLQU3gGpuDXvy9lqkj0ak9lsLHtDUI0SuBIIJpru74zxiksuJazJRa0o15S2Ib7
lI1IE+FUBdbPmz9eTPoE2rCUVlBo8W5zxN8Js59XDqf1j9HO8sT3eCDDSWVm9wEE
BII6n5ZBAKsz709AqYUUydFKSiry5LsH82qqigq8ItaeDgCk3pF0uicAZgcIUh88
prqkvG0r8cJVpIoPSgtwkXvQpS+VNXTUaIvMns65KQbNXWNCiuABkb1hO3yryZpa
UNjEg5jAjoEy0Wmf17AD5KTv9BTfhqcUKxRMsGOOl1Enoo4cLkwztJBmHlCWIM8G
H6+3azG5AdXtI18vAsj47N9o3IL3prqruMWRPuUFS626vPO/I4pLWp76yjLEnwZk
ns/hDUoTMYwGLec5R1fPW4m2pMOax8tQbXZ96MW/G7CGxNnAx7wdVzaSlNo8tqMj
yGV8uSVLUASbyTfQw8y0CAu5XrsStWEZDJEwGNMiSl6FCvfa2UUJINp8+dJlTAl5
dVbrUkH0Cf4ZcJc8vIflrjx9Q73buYhx57y5v8qqHSDWOIp4Na+Ta2awdU6HuffO
Ti3WqmF1ktv0qtvB4jlRZ808E3mN9BRb7U3KAWeCkcywHJyOUsGQWmgKiDN6QuGV
3GsoaWKEtobNzFlcMjfvW8KXh1iW8+mJwBpLXM0mZwaas8qo38O4VGFACI0uUcXo
77/yMsASwVK90FIkM66fpw99EmWhszDBxPxeO4bhHyDsregtDjOhI9rSaHzve7Sq
hf4D18sk4j9cqJLHiIxJ/ta340H3sgumJboqf8Rqq0n0tS3iFwzqU04z4vQ3HU/u
rdqrTMucqs4H23hV7dPyg4jxolJu5B4utHGi03hxzzfM5yVqzEghLwLwKc63eRBa
5n36DftKFcvh6uen0oR/Tl8Qm/IRLLnE7SBT8hthbrdlV1ahCY8AoLx00kYS/M5W
Zth+4g7FeK9c3CwmPkJzkOtOGWH+EYrkGv70cMy4jQqtA7wqsxrl1uoeIepX0xXH
mqn4ZK+N/fsc/Sfx00tFhErgbZi4VUUe3SOUfRQeCrECVgSOof0gcBxgaZ/dL3+9
qpFCWzEVLQ+26KuueBfrUFQfaKNkM7PolY82N5GlRvoyo0K5EY7l6nXNmyY9qQtF
QMPWvZFGIBxZc84tMl+kki2cbYzvtWqtc2V0ZFGx82igs87Lp6cHlFyEUFQSgcQP
nXRnOuI3UkD0xOaBuEILfNIpHuEmRwZMztw3awlhw5k68ESUFJSF1fyTO83jDy1u
XtwKalE6e02+669+L1qCafbvImmw3h5oxbGNOOkOSe61csSCMtxpgAxsGxC6V1t3
VmqSJWc1wboT2wgqkaxUH8PP6/yE02V3AMcLXH4m1wxyn5e0SE1e5ccNARhzfdAG
5et+OHdrdB6Au3MqsaCQnBAV1r0UIHS4IGKAobI6UsQxoyqU34p7DEcfw4hSucp6
1/f64nB+sAS+U5f8pnFq5TlYPDqboPF7jyjA6T/V20iGws+dXYXK0/DovTeXd83h
cFDDjMhTXZR0L11Non6JNwnKpq7pGbTLPHJryuynHscz4x5E59/weW5UB/xKWFaB
pasTUSB29pOkO2NWN9P7mVktj9dr2RMdKxbXkfCgq/gGx9aVGfBgP3LWcgr5477u
YL5ce0aUCmiDi3LomkKuDSn7TIzP31B8FxB/U9kBZ86vs7hYvTfk/jnZbDmT8KFL
3pn7DuqKoVnOck4Wj3dLVFROKip6ytkKPfXKL8v6YyHX8+l5nx/cf/TiAjlPIodg
b1xK+2fVYZbVkr3OQSpyHzMPQi4Gc1wjnsWp/k1IG0bcdtAmENZBjm49m/udXaOO
Yt/n1Npc+8J/EUj/LxRTGY3TyLeKLT1LY6GQ4X1oSK1kfWnzYpdWk5XEVw/olxUs
VB9JARHWlDSrpxj4C1R/hxXDgJ6mhbwv2E4ew92QHQwwOakH8lpBMk0gashRc74s
tyw0froVxM6Zfe4C736ckiipdO29+fSYqG9i/Rq1VMfL/Xv0rorMRsQeH2icZn4F
DBjggi0trBUdVsi62eAbnlbd9rt4tgS6x2HOx+uAlTLAT/3sfjSiEV1eZkAlykln
AWVDOBuZ1NXnx9Ja36nVvaSsMroX9pTkHriphMI6QRAVwM8zFwBb7b2/gqFMh9dW
GImWpmZcm4c0vHlNI5beeI4rF4eEYN5dfqTku05UoCnxgf6bK9SZKPSbdZfFzWhy
LQDqWwwsWi08zWhYzePwMkR6VtNByu4fmyTXLnWR6rRe2b77UwyC55ubWbMHlLF8
9AlHMin5S5DfaNdallRc2u9GZo3n+0yPuI0KC5fIyahR+DKZkQF0Pjj7+64H3+c1
p5o8q5URRWvK1vMWO9ZuQdC0eFYKEGrXLXGiCJ/YD+UqQISbQi0efiszjYJTKW3i
SPp4+eFyaHFQQbeYctzI0i/RpGJEdFt2uuYEVwkJvu4VWe0ED1BImZZNuSNdQipD
bxv9M1ijMJua3MOuvWAVghUpi5ScB/TRduhiAnKN39lwwyXu5ve6vGMDLVZTjaNc
EhvT9W+TJyVuPNAIow/vz2Xu+Juf1uYDhWMiVHTl/xBKl56Zk7yTth4/P4iERuKI
c1EXk7A5QRXchM4rPVcP6xHO8umCsklmxYU9wFEIAO7ZeP/uAR8phvIsTU1TTtLT
U3CO0ZVWtHE8lyBA08qTQwpyGVgh1VTxCCtplWZVe4BYGS9HNnN4J3dxX8VG2Wzm
CYa7Tv80R6gExllMxW4CeLeQWX9hn2TXWT62hIc5RlSdPlH70k6WHP/e5vIKbjKU
+ePOVJA26+ajfvtnYSj1XDV0lEVgXNYOwYFBTsw1tZyB2kmlTILmWkh8IOyqelu7
R+PkKmHCSsy4fMexjpMEhgeLP55c2ZX2n2ATmh5vNii3GoJp8hgstYhExRav5ex8
wJMctUpy39nezGgtX3E0sLVm2GWLH+DTYQ/fedievsusAbWBaagRohRV6pDu8G0i
TzhnzCbiGi2Ncu2ifCRZXZsz7teS/hVoUFEW/rsm4BzCgRu3xcr1lzNWWeRfuCbQ
u1pBIgb3GVPQFpKjAebC2M82KzE+IgUjdkJbrBfvr6KRcUvGNfdbETe5ePIic4go
ucN3ZHKTh/5vO1eVuzEwVLucz66SksaC+oON6QTTMvXv3+WLrzjIXgmnmZ4vyHEN
3d2sczOltxuvXAzLm0sFIlY4cL57F20g9gIlExDI1qIoEbh6eMRcU48dSRDoRRnl
exwsFAwvRNSPSDngs6VEAxt2+Oe0MkIUYsXfgEotag2hhZvx5MEncV08JWoc6N2v
OLxNJSlBc0Y9Y100SL7MkDYbIkZ0DZ/42wqwUVZL2l4LK663/4YGBdlOKTrrTrrk
v9E+C29kil8y+9gfl3PO4ZJ0vaaHpgj2pRshitBcwlj+pDcqsQnQfTAXV1a8pWFh
uzwKq9jV0Wfpp9mefqXnnSarBM4tmQHOIeWGqSlh1TOft1kkngoXpjjZdRewYK3w
J2nTj22iLp6xln3FoTpJ95fJV/I53wY2lUSiz5CIyZPmO+0zNX3ri3QMCyWqaOHT
W8X2v2nj5NyD/8gbXbhupnYfKho0Nz5TePDqIGdA2RtBVNaqgRB2g0fMXr7RC+c1
yxlTpwy1jDiBRocKNb2BVPBLgGr2QGSBCF9CKGMiTN4GGbQx16cjEenlDM2+u3p1
BIl5s+ILnKnFoggapoWVYFIOliP325LXOsA+zKrqUNccCmTXXCRU97wF04Hs+uFB
/f8FimMWy6G3TmhnN1jb9WN5Vw95Xqs+d03BVyLi/0tiPrQ486v28bK+QWlMyrQE
rfm1aXLLPZv1G+3O7nEq12lsKb3XS4wglm/5OujkU5TldRtT9JGdGyj9Qr8WjxDR
B0odVGx9iY0KK8BhLtcrYeYFmjSR/YXhg7KDLvyvT749f1ph7LiYO4blKpymlXQa
snG0NOl8Qimrc58tGagkTcHOlHEFjUK+CZF320mIx7JL6L+KPP4pg1mVTOYHzD5N
P6H/mVg+BeTe6fHNTAndF+dajCDcPhOpeyktdvpccPj7vfzz0Did9VjK6N4DnKpV
SivLyovXA7jsmSmqFAEr4amlh11YUxXO6HPNQOfFEE9ADGjYoXtFJibt0lGeTt0d
UGDAmRYBF3/Q6HRj7g0JNf26Gy0al9hcShBOssno1yRhTK9UTtc0i2LmhljBRBSp
4DX26Ma8S4Dwi4AM6cGVKzjef6lDRLEZp4Z6KWqN0xar7vpgJxqmTBxPj4raUQWQ
n3xPmmKllM93ArUzf9yKft0LVbhO4qHsP2J96otLXriBOmE3S2Hww2W8cA3C6qjs
RNAmjaDXtbR54lnlfPdu6JYn+gL24tO+uDGpELP9e2nd0VQ6Df7dE1yYnDreSwtZ
lWPS5wXdcmCRv8KqIn/VXZd/2fq1qKKNucH9yXtkkocBewkgsrIWwjcGzeNVoQ3k
w9I44qMDtqPddE3Ccj47TPfCoIpe1HHSMnUJtH/z8s6rFKMRJkpVXWrUq4eOL/PM
7cfol27uUE5Flhs8PY29yt9pDXQgqB31dG7zRHuiXbmYQ7KMlshccCZWsvhi/zd0
obF7b2xKMkUVMxWDmvryvjob4gSzfyRH8fCv8TLdbaqOIGomjDkJ61YAGp/gOd+k
/3jGgq6le7Amr1JvRXBLN8+v92T6PWmWYNiqbsPhBDOsnT6ypUaEDe8n22UyDHJ+
RQ4BVBzq824h5IEq48TqGxgu3xYE9lbIrXTZ/qYxAiYXWa6hnJfCDesrm+AwacmW
TMMG1Gn9vlcPs+Q0bKrpP1wwq6IWPDn9k+Jodg9F8dtBRwJSgwezTVIpE0jmNwNe
EiT7BZGYDt+IrL4alPNraI6kv3WDNXeybvx2H8aUoVwF/ZjCBoNNvdXzNWfPlyMI
oJHV+E9KGPCFETW7TX4mK9cOiGhKYOUUYJJzljjZmbRUn1nL8F6FHSqRQ5oQqml2
esxRK53X9R9zIb8blero0pvgU4j8tpt8Hu1Wk3Ibt348hsuc8isr/kqxhp9Z3Tar
RLfpDfg3FjXQpyxFPNVCrF9HYUO35US+Ar7Q6R3gpMKR9LPFdV45HJYtRIbm2Fem
PfjXO1M8CKro3SqxXK+QnPG1M6z5bpeX8U1a8iiuUpPEEt7L72aZs1IDv718Hztt
xYYf96qiwxgQ6MS/nrVGG2mYzCyUvQ1ksxR5rcCB8uzzS4hOVZ+rEo/tmqhadpFA
fAQ0ehvFWcoLQplTpyr/EIhv0ccNVJvT48UxVgsnuR+vtZh+V6U3jlwoq1wnV7T3
wmy1jEE2CS5c/oTeYcKrPe0xXNsKbFDEj/sTzBq9VNp/be1fmJCmPbVbUlvh5jLH
E+UG8He0/OHBoEm0KtuJNjmpD/0gM88chWUB0qtwq2uBrz+usrKI0GVhnHznYh31
hjizpnEZ8Hdjo235wRJss3kJNQqf06yrfluuy0GJjtKBfDV7X85QubnJk/DwPnWP
XILkXKaOWFQpBsXbc6QsUEWZ3LGyi+TJ6j633lyd7lTBOAXd+vvGJX9e4XUUwqNb
zzzik7jj062ENjL2LYLIJaWDNJ5MoAE6DUP0342Ao4kdPoVVk823shqQthU6E9yx
C9GOWKxfnLx595ZJXRGiG17wWkWyl+OczhenOyiGZM6GWgshRtkaxo7aZ06LpM6Q
abg8T1AUoFRWd57TScQJ4ZG8Yxu2Pc0mlWb0IYMYJg8ENqJ926aZjZin310Ib/Cg
3EddWYCLdQSMhOM2+Wn86ChmayrrhgJz/z5cJ4w+wdQfUvR8jM33ORijbNbPAoDh
1b5AS96VvXLEl13BNjIgKJgxRl+a6JNnvvVquIN2TC3CRrbMQdTrj6cqH4Hz1Uw0
MA0OXnvNSV85StttEQN216iV+lMDDhyUt30CK38uOHb7cgVA9GU3W2HGLEuPqTy5
VwS6u24R6HGkxA/qk2fsqVIu4J3i99NfZLC254lNqaaeAJRNs7FestoMkdGgol2K
J+woVo6X2ElZosvwAwMzhPeBEYV5F8sUxohUG0xppAY4shq1m4zqa+AV4jWU+YHP
wr1VnQrFgbF3zwx8OQ4z/ATBPUIk4VT2HrfkAKn5Yr1+nuyB3rshiFD9uohy8Fqp
pGlFC8QK0aahBRuqbHbB6XoNN9x58mF62XZunyWrri2n5UcoHaiLKnzqwPlCPHBc
KTiWtz02aWxeIB+ZmhrHVPnt5F3+1qMuxfuhXHxuDb7cDgCdGqm4Mx5F/QeMQiI+
MU4oObqonMmLI1tXdYQagzOXxowfZOfmSCR2+rgHUJhcc+Dd4k/4MsXoLnVee6sO
0glyHwaIWHN39smm11LZzTS8e9l0Rtxh1nm8gOBZN5kcLsW8uIVlEbH9jKVx5nEI
Gcz/OR1v+iwVCGr/I+J4onFjpOZjvkdU1ljwnF8QwB+XmMaZ+aXX3GvkwbQvpld9
gJ3F8lZYeiwgUaODfTyo6o4GHzPiSrK7VBeBl+h0p143QF6Utrr7VB6RnDeBYxn5
AOeDf/fd+Kdwup6WbQlAzgB2NzcYF5DFp4U4r0IqJgtSx+tmXpt4ZLEUmcK9KVyx
wNAk95ulYBQv78k6FFhWZJrRbiSjl8b1G9OcFFBUy9x/W0Smg17yY2yoZFgXI0jD
XOm6BIVE11o4tZWaYBPA1q8+oeLmp7RwgiPU4GTX8CPtsMqlXByUl2opNHGqeHEn
d26ig/pKA0guWw0m2+nNqs36i2QiWIrjYneoHsxR9Z2vVUO2G4cQObkSi/2qNNz1
kfceF5rY6vDhhQeCj28D/hKCD/GX3IclySId3eN3LqiUbuBeE4fR2ecvqTP8CggD
mO2ly4PO1GSLtRDAMWjsXAmSrhqjIJiKPlwdiNZUlYpQCqba+Dqn10ZjGJtX/cUB
HjtjptGTTUjepr98WTq9veL2WcWVgoKf52tcoyIO9jv5BMAkmDcugXLQSisyjPsg
DwqVMowY5BDidXV2y98GOIJuyvWzWYUiDywQNgVba1rmSgUZ3oXj0gzOgYcQlrVp
3MXZztcUIdwkQYNGFRcrxyOKGZ0un5bHsZestFSYhMpjGlP8IgoTTP6VeUix8gtZ
Hnv+5od87zKzdZIjiRl6SuiLHgb8L+6RxEnVvrlIoChgtitFgSNEF3mLmRr7M0Bs
5FTNdbZ1ZAxTy6JyFXgsJ5PT8gJ4XKlKs6VW0XZGj5446iea89x191F6BvBj66kA
jS/BAu+v/KKH8scb4Bu2PMy5zKyvOCQZ95b2IuVPHq2oIpjJJMFfNzT/s/Imb2gD
OdHe029juAXDcYW/225QBv9QKyeFj+GaLyxtRAPQncjm+ZxgFbjHMI7hG3uAq3HZ
Je8BGvhrHAIaHCrwXiPAZq3t+WFuand5ozZP4RJxg79CE+0DUOR2JdjoifZIhpNS
15hKSrTOAQdF9r5qFLy4ai0nN8RmQL4/aOdlFcpChB8VSoUvIzyphY/14uhEWGso
6rCL3yFFNmd6FyiS+BL8h8ifZlSHYlL6Ua955AGnqeMGowXlLp+aFrsdM2pY38Av
GKmNMhtDmQrxDeYSl7gC/U6rO7ewhVJhGTIAudby6XRdZQqMpUwh/mSeHvn/OcB2
8NWnM0h9keC1czigCS0sfZwhguNuTouUDMFfSQgJXUjh1owymbELRaJ2cCQtggpu
6eYHWc9FAonwiGioap4y32Fp5QXqpS3swiCIGkAVUo33YI1Ex6B3X9DIz8IyEcoH
awukK3Lv51WfWcKeWkpgrOwGpXmaICYOnvhOmW6NI6PAL3bsxaXXp9BGgTdvTV8q
cK6Oa9B8DMxWRZcTcO5RKNj/wzFpkq93C9NiESEHM2o1lgzgmdpuQtiHTd9Jp4NA
KQsOtkWbnYd8AQXlSdZqWHRAP408J2jIahsIk+PjLL0+78R9AAh5N/hUGL58mbrc
7NmAWtBY0nmlri99DLw4jTouoLTpQOMK3y62p+pTeawpMDkFBrZk8jpnNCP6cnIC
e5QbZev+P9smACYibnI2JCKw/GAPxG0bkCS47lC3MGRWr/KjUH0djur+OSmguzrJ
/UbQNFVfPSDoPB85uV+RvObhQwaOQCkzf2t3Rg/zGZVx6bZoSC7MQdYlCw4YDqEU
LSW1K4x7YktMdkVZcWrFEJ+ecvSl4mLs3p8vqFEubETPZ8Nu594k+nn+vbWRkP6F
KeHXNRkaWhtK+twOA8IcxVkRdtUG3oYWXwtluyOrhmEBu//dOp1Dp3GIJ6Lcqf8t
lmcDZwGa3LV+A9ZI8WRx7Zi+ru7g1WaoxxLtIbtzLHJ4Dl6UELyyctPPzxQNjA3z
wiBuLn35PvWewHE1N7swc+i0V+Me/+6ZbL9g69Vt/2KLYormmJk9PRndPiE8kUei
bFE+PvxDl5oyso8FcyjEmGNIkbDAXTmba9oPx0qKwcfqmmKX/LLk2etJZC6g38Fl
eoPdH0+P3d+ci+14R77w7HOgN7J7kimYvzAmLshGZ8BRAnieMdX1yk2u6WtEF1DA
2FuWe6xz7/gdbIZFh91dDz7BLgDX+mD1nrvaDncW8NGjHtJkxw8CDmCMmn7OUga0
v7A8A9JVAk2D+xdoxG8Q1KEYU4La0bo63hwlCJnHmyQpJqgIN0gNvYM58XsoBay/
dat/ksZedR+CBLCMUWcdQlg2FMwVKuWdmqLF/7OxvHQ/VGuD6huCew9Eke283mVw
WShkSwPGQYd+6TpxdA8Up6Y6uzEs8ep3gYEQHyXkDZs1WHRb9eAhndjFtvmrk83S
zPyv9QvHhgYe4MQ2h+el3UccCnjd5Oye8P3Up6WiJ9A9Y6mG1e/6ZibMAdVmz5IP
ueDnil9hE9sfBLSWYxFzkimklQpMaUtE2wend1k+XLCbX99pp3IE95y8+OYIdZT/
/B0bJfZq5EZuAe8kiqNfvXQof2j8Jkez03fEn4dQR4vRRphTfphjseuiwCrak2cE
ycdPOqzpgIFAzbrT+Dc+oi5O6bBoWEv4gBbBa439t1eG3FWxEJhtK942Fnspl+re
Pz8EpOXC0HWWdgMvTygor4FBKMFsaufc3ocdNQCYwZr69PE3XiXgY7W6x2C6IZvk
7bkK2ILDZ1wF9K3Jdx8ozknTGWp0d2iVrt4/GvwdIs8sx7JwawSiReZskdIXlpmK
3+cyUTFHtxKAQonJxpLuOO1/ca3drECvk+FteLFpXT7SyMad7BVbmT6ZDdlI8HAd
KMF9VgiLXwTsGF6sGAJhvznWeEHrtu6pWIWmvOiB5eflw4Gz39/FYxv+u4dEgTer
fnG226XNAZZHaj9B9VbcfPjd4vV2g2nHgfkoGUS43rqyU6bFouaNECoy4lK24aqo
dG2gzjxRsfRbuXP0GnVY+wXIZk7MEEBW0F+0TdX0976WKdngYlBkatS3X2eBlqxu
shLHZVqrU9kpSv8hZd3Qbxgl03trXMmqeiSQsDw9ltZfbp1sJ4v3RCFDStAbO6XK
f1CQd2A/00akZubbvzPGxW4j1ocr5Rt8P+fi3pInkvkIb9h8kLHZk6aX3p7R4Wok
RbQODySfHR0Nyx07Fm5u08n9Q1D6o6Jm1/OPl2a2B/p7wGA+yJIGsSK1z+ZWNUlA
9BjLwIpJtagfLVlSFy6+PZ7fVv8mpBE5z+hWSpulaL+fuNdNZcn6hJiOdzqFM0yi
ZdE07CIkxI3EYTOFp962CFfhBD2j3J6z7FPqO8TqGBMk8H/dXPUfP3Fjb11med9K
KVeIw9FdTqvFjrcfaSNckMWSLH8XXSbdJ1BAERBHGqcsAi9giaP60RfvbuOeA1wJ
nGkRp9ow54ltbTSUG6w2WhvsCRttZrQHXdE5xqnmaL81dTlJ50+kp4azP9bfdts7
yFCq2Eh5gAd5TenfQoJmFhFeAftxWzpoBn63U0p8gDVJdnX/rMs5ALGHMd21gfh6
P4SIhtWqYXYLoW9Omy1QM8M5Q2utE2Cp6vcrsxVD06dzX5hwqu//cJr87l0ZPZzX
kBgzmQdL970Hqhz7WxDv2clt+rJiMTOIYofr6aR8aQ1oDzzvr93OA8v+lokoF8UP
5g6QwpYCs4WiaCaxdcgIdCTOcpCz6dpiz2TPVsYpYXkKhhgCH6Dd4qoUAWJN3LGy
/mj/vMHryYJPjzPXpH2uAV45ZRWKPr9X3mjcjOs+Br2diprfZmT3h195HdGhO5lz
Xyg3Pd9MEz9itogI0nhbraDcUoSqdvGHEjEL8SqcaNDJzEU+js3PMyL6i/hWPv8f
pxDjequw7IcMonvE+FgcuB4nm5VeB5dlocD8/Z1t+eqQvkLPNO0I4YHVx5LmyWzf
wCAJnRmcxj6ZY++Tdk5KfqKE7Gx6mk/C+pZ+89scbF6iO6EZeYdh2tgsDpGuKJ3z
cf0+J01Dh9MgepDyZHJdPbQ98lkDMbxXA/G66XrxhPsxANIO2+t5VvEucYXNZecX
bVtXjE+SFJIWRg/xFEq1O5uf+Zq60HCqP8UsuzMO59pcBgMIybNvJ6+Ag9lEhSEn
B2SVNwKkr3Es8G27jp2G7/8588Nilmg3kxJlteeO9hVTS/Gv/wI69H8ofNpXHmEy
Jk90kPCQZvF/Fjqlk2FM8mFEQo9aNssS/TBvRFgxDG6PKd0yKKReUVtthhWSxQVG
r3Jrb4f+5r5er4KgFn9n+tMPlaLCkwtR1I51y8EJ4aYJzXbu8/4NWVGL7Y4HQYw0
y31k22bXC6bYdaLp6IFT5A45UjxdvBQ2nKHLKIHwoBNP8POQqK+Qj56/t0qwv2Gm
dreF6G7KBTnUCOS+MsdyhLiMyPzRgfzxf67//SazH/ZEWPBfE/21dEDuTZdPIwI6
hjKJTQ9A6EX3r9b4y2ggxPLx1j8gEGw+Sngv9m8wscsaD0VvZznKFofY9VwJu5CR
chjpKNhwn7G9+lPwTtn/JeYzjDUqRCjOhd/QIen3DLtLssGqtIrcMdJofU2Om89o
j94j64XmAZLKpifAxmV+M163w8MyXEi/am8ENAioSA2d/3ZlzC8GgcDbneDdB6rA
dt9JEp0V15xzzwbYLQcw2qu6LvOtTxMn+nde/cXwjZKltps+JwRsXREjCVwSCmbj
49W0iwG90SgFwS74lTJ4tSUihwdu8g4L0LfhtuLCQcQn23/Rd0Z9NZvfyOjbp7VA
57+8jSmfoMIrAx+q2Mien7Qy/gj1sepb6UkbAcE6LahwfJHjpPLaVAAYccx6H1gb
Ahop8eoqOuwHzabsQjVKJ2w5s3oqCsPSpEmFV6YP7K/+mT/+RU+IL9LBP7w3nILO
cBFNA9a4bq0E8OB+vRte6DqyaMG/C5kHYaI9DK7bWsETK6SaXYMZRE9upS70ql1q
vlelNiPVUThDtxeVZ/2qCYsM3MinvgfY9CUFFrPLhZQC/Y9xgixAwxcgWUE8pGWV
Wce12yLzj0FVuX0ikPz6XWkduueMa4526NyB1fxEkLktoTTg/GMJHxY/qtPxWZ8Z
/cGaLuhWzocB40HXB26A8KiXv0bTHvAdYd8WnDBTHSyQjXiNYHPbSwDwlG41u+L4
zCcj+39la5HknKvIxg3wyZdU6wRyVrvim/qpRqlxCKcuiMp3AG+JitpGH4d/O11W
T+Pg5tH26jrJZ8TMtsBEWUAakpOkVlIKn1Kgpjv3MisxjL+xqcYYhBHmKnJDGSSf
5ZWDyfrQVGhISfeGvaYUGkWTpmkA9aDD/jv0W9oiSSk5B+FEgyHayZPiK+HkOAst
l9r4tMopgYo4zkC5AHL5B0gSLUNrOOBQdTpWDj6BoQsad2qANtcUSxcLGGm2FrNK
zKr/Gd/wB4MOZFh4zFzph2xSi8kEooP122tykPbfJBIvT1GCAEJtjadqc/eboe6i
TEvOzdOad+7sRJpCb4/rxwdoORTJ9W4yDqCNMU4ymSsFotks4oKo0kP1nEyF+tBp
8n9qlzinP069PwsJK/LiU4yHtA7sNftZLS7aPQUVj2VYK5+ZqHyTszX5GLLrHZb6
on6F+ADTjA1b/j6n9DS0M5z/IO/RyGpdKBClGGa7P9Z87D3OrkTcr8wIZ02qazJF
qIY89shGL9jewmjmyoLUm652fl+YPaRvHdkH6J2UHmj+64+tRfYRh624A55xLfsy
UI9TRjC4GvJ9nPiYGymRwHQUgxnDDo69us4STEyRD8M0gruIJ/2CGa9POBx78lUU
9/liKF1WEnqq958afZNqQ/LJcFYlX+2UtyPezwriS8qF96Nt06Kq8gI97xXNpv/a
R0O1wejxBpt05VKGapUn6Z+qEzFbQLbAriqMCooMHYiTUo7h4Iyld2lzjsXlTsGW
wrVvDzZMLuDdHaA2EUcfaMqu6DGymeBfU7bYws9ciWX/FRQFS+otCZMcJcuW2LqP
eKqT7volWKv6BgyN4pKnHhscB1TrdsynqelXgDF4ZAqA07a4YU+3J0yF0XFZm7Bv
hrNpNsPGKTuLImJRQWHBgo6vXRaeNOyfe7Fh2x7swGRwGbwwQHr533xMgCA+MM5h
yDP1/YhqHndNRW6JL3VtMeaVWVgHu8WTz7iWya4V3eum7481qO400PygQn102Ks4
ogrIyrg6aSEIE/pQeNdx1Z49QwCLRVnkXFnZLfACRChEiFTD55yUAfPL6okr7xI6
Z71t2GKwWcKgVhC4CZsCHKfsY2e3kqgt6onKuj7RIudTe2KBrwJ7GBGpWYZGeZEU
zAAgKHijQiqkYq02HqoBtNXgRSmgxAjc8Bz/0Hwcrcm8M3FKc520vpA3OoX1fWMp
/aG2zKxpLmEsVzCMsO8iATunKEZl3r95DLVh0tQ3JQ3PoQzdXeADwK5gYG5/+tAH
AbLO0fFx+vqJCNlrDGhYUnumcdiFK6Mbq0hrM8MUdZrm8P1XSwwjwtULm9ZpjMBd
2NHWDdr6q5FUy4mnYNj7yk7PrL5lUVJKCnjz3q0oal1oC9ai6mbywN0nIi0UCZ6h
MS2f2JhuRqVnr7qRlGWkolXiQAPFvxE/4Sg49DH6aaaJI6EUCC9XFCYrQEs/VMrX
QVQRK8+GBjiWm65ITZGqcQNssm2bWSswDeXx+r6qDbMUigpIUl5Cm7sMjNvXHdKv
8ZhnxEyxSw0HZKgnggbo5nnYI1Fr1xnjOd3BV2bnPudzc4uV/RmEFq0jApgByMSF
Z25WlFrLCpPDKDvd7ZS4Ok8zvJOGGmJvmx1qloaPH1tGWveHRfUJ4C/25BUWHWZq
NkFJ8vgRwSgNoVizTbJz4iNFODXctnyVEmSF8y5hVpqNMx1ZDzBY1Hgd/y9dhY4B
6nQzEv4ONfMthCizCO+eG07khC+z4A035oUc5cXV/8BEK+TDGeNjavqjh4a379lb
g7FkgmWFAi2GJAFtdqDU58+Fd/x4dR0aNhmo2po3H87JRdiTHA1l/gd9MXl/lW43
UXhkf9nG0+XtYg7hCbn8ktxRDq79hxbfQ1mGn0U3cQdT49t4NslJoKbdgUUIBH8U
06lwkkpI0IT9kpn4JCjNQmCFLYqOr0HzMBOcYi0j7UnDofqv09nY3gx6PFrMA3Fn
okSxQcRKdk5eBmG0dN2ZkiXz2f6gFvIutzys72LnFrtTeVXvVM/jcq0SWoF1A474
zX6PG17zdQ4b/e6gFtLuwvIz0vPLPdJr03eSFHUSca+8hrVy/rmgRcbra0WUhdU6
sSC3IvIPybnePFttDkWWXQeh+kTwT+uKKJrP6m2JN7mB7l5yu/c3VxGgRozLpYou
WCOtZlP9A/wVpNnXwKGRtcwf9TPCS3ysrKRrtI9qXQraYPw4bJ5HGmwWakjZ4BDV
UHGYMHmCEsZ6q7FSlE7LAtlJmrfJjItFgwigy9pMGeirk3huQV3QXmeoYoWQ4SJ2
s3GOy+U/kI7FbrsxTX3UaEcXouzr/cwyYfaJ+xpBkJyM9WiXGr/wHZbJzlo37G+5
88WfBmi0cXiatHQCnQuUCdAdKkU1Qy2tUY6aVtXdK3+XGxuYZq2Cri7Njv7jfc+8
i9MBTfikISYp8UXC3ywOKLOvvARoLtCRPynqbpcFypU3/OGeMYW9w/YBLQhpIxvN
/RbNk8xBAev4NOlxR0B2K739q6DdeleRcXHtugbT7pQ/wM6HvxUWfns0SVcDfkee
6lEvSCefCgAOdzIHEO57TnG27KDCxnH1wkzqYATTD0a6Tk53Ua4QJhlKvnO5IonD
UX9F3c67IWJfqTC1KXiwdgXFXkO51CPo8GuQM5jzH9Hf1kdvhM/4beBhZQNNiIOs
uOhR/wq9NKbMRsk18ZD9rbmgQCQpEkfwrAS8G4CstknqxtWdoHXtCkBmU7g5bGCi
p9cbiKqHD2ilhTQFO0z7OLG2paxJpp22uXCBCDfTycBUXERbhHR/kz4pRaUcXxxE
7OoEXJqWWgyRHV8AJJQcnm2faCFrT80S8BKtmWk12o19dObU6dJU9WxdSpbjRjjf
D5YXFcbGOL8hNytLjPYX8NL2Lpw+nRiQrklLnNODtgvYJTRBni8QjF0MhGWO1kIm
DdsAn4jNYWORgA+LlSgIaScG6kOzqbAP/2fr0xO+QPbeESYY9JOKT1cKrKxpPakL
9YXEky2dqELXli6iAvS5Mpn5YDSbjWijJGr6NxokhiGjuceRmWQ5Srnq+Un+6bbl
vClztp6yClT2sNCDNAqtwIg53Irwd9hCAea3t0SnsDPnJ6+JMMQNX9tM9auWnSTW
SUejwq1Zb5ZTUyDhm3BqMvkrYb+80fpjUgkO/jDTmpputflK44KzH+Jhg5GqEF/S
DUfwxTYJO6XOtKk5t5ZQBvwWwWiKi4UfnK9p4N6jnrfkAmbx3pbuXwjOTLKC+vjO
d0nMectEwRSVjVsSOv9s0cl8JCR26j090+hoCTVQsrhZSsZ9tXKsS1BVOtMOhnC6
j6tKdcelTKCg1ABs6P3pR7yNfpkMh83Ga/tmZIOXREysKDN1q6IvRAQNZQ+PAwb0
bzVHB5jr7Ktkfm4EWz9Bry+fs12eVTXAqykWhpJeLQoOa1WUGoV+ADjgyOeOLxcr
/pMZxYhHn9m1Oc7E9wdnIOEHYAahkwHQB4k6XrLQDXoQe3dga+ozH7QoXfOHUqMD
U3PsMgTby+c1asgpXz854sBB4Ce7MOWt6QP4kmqfhscxnkCB4loHuNl1XXnrFS+M
UKAfp3XzymliUjMkQJoiawJHTeIIubFt8colOvT+2NlnTSE/X2yDDulESsfbabs/
bw5KKXHr1pqb+jKEPdIJvS8B5DBQu0I+O0mnPhXkRHFZJycuDypKJUlM4KOFO0UV
TajtdOJmrmLW4YH+lAzROthabvXUnJb16uNCqgvfDofSeMCKwaYiLPs3sYHMA56b
Jm64pYrj5Ue1fhU27iSaDN49CNhi8ilnLiwF/riwwDYfFfuFmRm+w/KTW5aJkIPv
m/8bn0EiV4v4u0jjD1+IhPtiAjfvqZKx1LWW3Qlbrmz7P3i8SLj+jeHyzIuK0Sp8
hWye/o9gjVQ74zKgNNjQABo0s6ZnR66LPq/ITsDSGyZvva8eu0z0SGqzzeejs8Gz
L9H87WvQQhFL4hWyzixTa6mESBNXBNwzSrJvXAFpbfrjQt8KINCTNekPHTBBlPnT
RqLvyOEJITQfkh8mo+8JV81MR68TrPFUCdgDXTq6M5Z8PC5+fWkhW2mUsFk6IGyY
m9D2UuFsA3cscrZTe7F2l0qMnrlpMVQI9xi8kHmmkMKRVaxCo/2GSsOOYpyg/yfg
t7iLjhJGinrZq5y+HJCDcuvf0X4H7eLdkPWu06URXQYeQdZQiBw5vltYkCfPHh12
Pej67lPWQ1VotIVhq7pp6euPt5A1qb6kWooQLrMWM0wcaI8EcVWHx9yqeZn4BjCV
cVgOwbzjqyq2fLAjgrDXkvnSySWW4jNBo+uBanqaKAQpUKNzI7Zr3am9VjXWA63C
jX3Dq0XuoKaFxBnZ1N7/8TefG9795C0iTbZfVosDc56t3+3GDKRscZJiARBiXkiQ
2Hh0N/kELyCa9f7l7qYXK8hLU3pCU6aI44wTSMgxMIdJSZdCxVSHyFxmseeAzKpZ
zNxOS91Pu6AhbPyiBB1bLOo62OGXLtPB+yfYZPe1WyzGbkDZqegPbCSzvvSnZ+ZW
Qh4vzBjfvlyAQK3KAKxTN04rZ2N4oYlDJUTLIUtKBkkWVKjtUwEgi61xCT9iQ3Hl
6xg+z9yGmOWKFc6kamyICDqqZo2T4TnCeUr9LzwgN4BnYjrtCCWfiKjjV2uCUvnK
RPd+azzdgvcq4nW3cz67KN40syCO0rIkncpb1TOSXjdClNBqGj2AOh+9FiRkJK7x
56CBm7wFTVgIZ25fbuaCFIQ5phLIgRepKJ441fW/0vFm70qDQwNJl9TANZIHb7Ze
xNnrtkiY189RjcULIGPwMU9qQ6BqPIHXFbRonPvK8X+Hs7KuNE4x2x3pn3vI44Wl
kLUyUeAD8bZi5lXXpowv5xY4S1N8Pv5XtYvqTAXmAC7FI+ZLqo6OIB8xqDwEFVS9
wn6zv1jjbBu1q+gfvFqJH6WnwbrIML8Vl1BjN5SBLlllRt+10dNDnZC/x85rx9PV
/mWyDmn8B3ZxwKUr/Q5pVbmWfTre4sV/4Td43vYILti4oCXpfrj1tYyW7MATuFn8
eVANFeiwWLlP+jCh64shIWUzAlichBTei5NywfypjMxYBggov+rVOxtmUD3frbU7
GqA3SI5UbrAiaDBTReGuOvAQtX0Oyg43rWadxcve8P+ihS2KH4nNisqLyqXMPUcz
isxG9ZqKeD0UWku4fxBvPYA5uDBlDzy9lrqBEI2tvGFN+CIPO7e0fas4OzyC1/ux
oo7WOuKPJVl5FeytG4ffDPjpJtNCnztf/cCQwiF05pa0cYQ3vZ8uqL/Bn+8dyVIj
0PIvUnOlYBvH349KDSN4vLvd0F325GNnlVzjfCGeqPbUDGOE4HxdlhSDNFq5PFFk
donDbPqS8K+jGBrKgWDOoIPuwQcQyFPuJSQxIW9Y6EWzwLf+HICSm/RwSyZ36Kdz
h5YHtgsGSnsxzoCLdpLh2y6x97NlbJJdxCMsVD9oeuFvPtn/9uH6ZrPSWTCp3Iw7
0Iego0bh4ntazUw1Y376ocEZNd71EaYUIZgQnj3iUJegAvDeRRe+eJ68cSsOVfGF
jVqvjQoIZ3iQsZn9Ch8YdB5FJs0fk+cSchPxnr6+0xms8CQv8KNmhGjJhOzB/KBM
baA0RZYFjmZBlxCOiffl34tNswwR+QOXjxULnQ2764UR5kt6b3eJrJ48nVCscLUD
Sd2SNRLZr/y+/2z3SDX7GlVKWlF7TDgaQQFWWlaVj6P/+k97ifqsmVG0Bmlg4J6f
NuJ0uC4qmIW3DNG2NI/fkdwNzhtxUZ/YZDnwDWwCeIc74VnjqWCiTnOtjd/HlDSm
wor/2f8obFgDcxZC7PYMhHfHmBPCv3dCzgbxQMmAacxKZvzqj4pc4WfT5IwrSTAY
6P7Cti3zLwQzJ8lCZ+HkxsW5xPglHoXoHS12UWb1sorFQdCMqR3dYtgcNG7J3QFg
LPQK6XZ8H+UH0fFNN07vdu/BWTjqTRCZK2wi19ldXHEMb3pX+wl5cG7h4NUdDq57
2DfxxCBzTANwTTJVmnX/MXzdRIsljtNtpX/xVcxVhBB62djUcyoMU67zDhpi938Q
cRCHc1PCbnXO/+zYfx0nBUPPCOZvr1zm7W6gswJ6sejHRW4KMJTFljqPXf1gVdCP
I8gInpb0eZ/CIciCNnevh+bZzLUTPJgnNcgEJut7bJDxTjmitfXhNT11HF7hOwsS
JPZOELDPZSAaJbo1aIbaPjhGKiClMxvAa4e/i5hPx3+boCUST444raY37m0oRSoS
kKOVX6PrTsdcz+r3hnWinPnAMGch8e+/gRA7UHkDrQRQTzVS/+wweoslETd8vkJ6
9ftiRtZvAlPwXMiqaplzNHMMpblXM/yHCvJZ802gJm9RXEoSrFoAm97dAAzemBLm
SJq113CQ0v3kP1UXb5FCCpd2KO4QR2R2emDJZHVlBVBLRuNeQJcF67Zn3+DmAdkc
+IEzbK2yXCufLz8ex0EtGdzAOorIXTlD3qYFqflTB2iqBN95Md1KihJXe2wSPmQw
/6pIzPXz4Rz/0SP7MgHM1JqJjqhnDKOb42hdjO4BN+VUiBZiTeYP+VHrBkoMfBQ3
3YGcNUfbnxPlboKXx5yIIMq3m7vxZbsu0AK02DfGVAo+mxyh9rX71gWYKZ6Ns5mG
usn1xlQ3QI2+3OAP+NK2nSDzjUCNt3/VGAGUsqhjFK29vW38oGMbM77m7OpVuSkm
iiFTVTqnHMRbItvem2+l3ftxkYK6aNYIFqKd3cmfT8CqKdoe007u8KGUr2uKPbgJ
+YlEiIS/a/l2Zhzo4VRNTbuHlzDJIufLQ9bIFB9XFhNYouQj/fdRH/Pq5QztRXCT
Q8T/GETbGEhmCPvjP+Xv15Q6ICbIdwWc8zInr21yi0KCKPQ1eyZ/pt9J9sO+1O0X
bpJdZ4NZ2sn9hgeMKIREhdL8CjtknJjDV50I1NmadnsuNQmZqZ8BJ5Yyzc4FrA+D
dOZIB9Bt8GFc2t1Sy4w6SLjCbmhgRNaMsxDfy40WgO3ZiVFwA1pUFLsEWQbC0jLd
JniD0OhSpFfJxnnLOJP48yDJzbkpQ1vW5t7iSdSNFaoFAg5lffYszBBuNcZAIs8f
z4NV/y3nmTwcs4ZUNF8N+syJkE1WF/n0l/pzciQHXp2VRBCRT8QDV4Jos/Bw081Z
YzSs4voWOQOhw/rmldn+tSfXVB8iq2ajEXXFX3esUHijyBUOFZeGoj32bVZfjue/
7GI8HxB/uUIr2YYPIEiNwHdgSaapMhzJnuULVvjCdXUfta9D22Rt8O1+T1Kqo5r+
X51IoOfx1X0P01loIn3LQUNH8KVctam0jq0tZH7EqavI492sZNIn+8aK2jNlTepB
H/KaVXNWiC16IRrH4iMgV6f9yIslmTHDaYs30dnblt1r/8CDrJ5uqacGlvALAHr+
tdiJyGIAPhpHMFeBwnDn1oD6KJCNW2OwY1bilaNj2plOlErn7myfup3jjTlASR7u
VttOuFExiA3/7Z9eeh+aj0b72FoYjN1Zg/g1U+wG4LxswWa7hay7fKf7hdx5IGfQ
mCMQ9Evq315lz8FE64IV5/yvr9UFXFOhodskMsE7y1vx7WS0X6Pc8tfYs1G5SDOu
4PLDDYfg68dUsd7kczZj+PQy5XdQKkZZKG9AkTdUkz9OPT9OBbmGh9qEVMmFyWvr
0Y/13nowlyoXtch8EevDDy9DGVbm8Qt5WT+dAsWsGT/KH5RAskqmQK+iUgM0xtGm
ceCLjBzYjk98XpAJPfaNSg08MrIfWTJtYbOlPJILDH3hL23CJDouCnTa9k3LN+8A
VVis5AS0jUvLY3oFRPaQZ9RbyrIDHbJD5YwTLpzzKkAxj52GSn0iEMIO9c9oXS4d
38fgAtzd6iGA6+3htbhAjBWnvt6ZA4TBBajQaFgwuJFOF2NLXNAPFz7u3J4+kC1Z
Pv3R4JHHAocZMwgJtVkkkREFTlq91hvK36Us2M3F/7ElWuaqfMLEjv1H7DXc81J7
2YdlXFvfZmqHXGw+xSqOYZyIxebIQDtIEMKy9/Lgq6QdiCsb97Kblxn4lEnO09qz
r7mv7x+DRfQDnLSD6+aM67qQF5kcjDlPdkwLya7806dx7dsd2hDWiIhptV8KuvUt
6YMWRZdyyWTGI2eD0wq8akYdTSFtW+g8zDmAD+WCPQxw6PxA7unT4haSm2c7tKXc
65CDluTScW39mooi+QP/yHF94o2gO5XoUUWzdMgahR+NxOOWjOrDLk8YHU/10qRO
ffswifn/BfpPOUhkuzy7+bwozb7kFTrbcd02OdmKM2sO4jAgB8sP6LWX3si0HqE+
PHKVHBN+KL/5mcZuWMSdGqJyQ38eIviwAQC7lADlDvw7Oqi0ziw6LEqZaZcjZc7k
vVR/PIlIZEpeA7NhmjOZEYtmz6GHZfDNAsZ+yPIZR5o+S9Tu35GWniKnbn2apTUQ
ZZkqhAXZEtf1ePhc4FYjtCuBhbmD2f17wXeaTAX+SJmScISLyp6W9g+X/Ath4yVw
8pv2u/Ta9BIO0EKDFzhWrUifpKhm8F17ig2tNy5wIQyL2vqoMiUFk+CW+eSF9rzt
RJLfq+oWxblrQOA7FEMa8SjqxjXDjl1vQvYXiRmFrHzqIG9cg/dLfJI2YtBPPGFJ
N5pQz/NFD+j4S35BRFAJrRxQL7lDffBwVIaUzI+4YN+VOEa0YnzPkOuk4ozv6bX6
stjhw1DuDNrsV3HuZalWOPx8kOVTplkwIZ9AJ3BnDa26Xpy/Gj+9V2PNL+/Tj0x1
wBOiNJ8JtaTXQRfPbfIgsE8q88cEF5T9uVG5vyec3C3WhYSuJuXJjJTHJZD7qFg8
u8tD1mQ0zqCeux48IXg3TTawdxzWg9U2glr8lSBtLVk/yH0y1hB+N35DGER5iUK/
4l7C+BCjwavOflvcbYeLUb9MwG0az0fInOIJWrv5Ug+Xg0Iqfr9AyrH/5/pMdRbP
Wvln7WHLeoDGvdDziMggnB4Ccp/xzzoJNOPN2E6l/HGuq2Hs6ypk45R2vV4bRRn2
HnhcGoy7h4LU8BaD0a4a2gKq6xfV3/dksLuEUUIJ5q8Q/jMnvx3dMcyEY7L9xOne
8CWMx9bw61zO1A6eKRGhn4I8F5TMpvLtvqMTUHCr2q2uVrbhLC8GOA69l4qCB21v
70hK4+wvsYWmLPpdrxtNUp924xx0B6D1ZV/AhIZ9l+Ie6Vt9VvwlWmK4tcYZ+KYV
WX+/x8/gP28p1h3WdXQ+ibP7mR0HohUnyaVty0Q3gCwunasdqdOPr+x6AaKqL9cz
8yI3U12vmzwfekl4nrJ/sd47sHNIEKDfrRChV143QysjK34I08HduQfRTmBZFHED
gwFmvdYMDD5RHcLTa+GEdQihJZgHhR3VBBQdHCRbJUBUuXhhn6PYN9CV+S6xS2C5
/unT3AnBtcLrKwYoSgpWtp60Pe7eL/xSrLbpVTQyL4/9s7zL8aezKAslluXRGObw
LODB0lKjelwLEImUjHaYerLV1uwP0LXFv8PwP61BvBN9De7GOigS0ALMy/eRDwHa
L41BFP/hPHTVzKP3YBafxwOsv2Vy/EyW2Ce3BK2CwyRFg4Ro/5NdgCzasUZz+Msp
H/Lxg61AQCq0N6lFQFNYybh6rlDwNvkyJM67Loo6V4557NuxGiyw3uQP0sphaUib
FRkeqGVBVB2IfRlBz9yV7ts7rxscLlPXY0LQrPPRbw4/LCulsEVL4pF5agCQU5wq
zRLW+osPcoNhcyhHeu7BOynAFtsVaFfBoC78hrZK+tNdcGTLlLjpeh5ogemx4ZpQ
HVcSDsA58Q+XGVLTE0JCR11J2GM4QKp3v8qKzIRvyoJy439p1MpODabUnuO3p/b8
XFOjckzO5G6c0iZjvC3QyjN0F+IkywE61mvlXYcghNhX/EFeCbDmmUJXEzhcbd3m
U7uugLCxlfxm4q4AAqUQRXqS0awPcIbwuEG/Lw15RSmtBm/yvlPKJW3dd/aaaBP6
6M+/or38trAKRXE7VAsmeWHXEn8jnuqWD2E+hxgloMkNFv/nOIPdTFKf1Yld9YdL
c76Gr8Y3veLTckV0VVt3pMHup8p1cU+pEEi8kNtlz6jH3J9qfWZMrp069ct9ZDbH
YgZmlspyeG6w9SKWqle8kAeViEK42FYkyygxxUxvpLFnFe5lqfHRekDsLcaWoHd5
5q/qYUXWIcSFmq5GaQ7GjEJpQeM3oxYalc/bQD+BbviH58oLPxbQ+czXDuw6Njdq
N9/86qBuS2OFuRsC3n/u4aAldfsSeoMzkfxsF0aIF1K3+6cxnAJkz/2OpJ5kWWVz
ayvwaOez+JTgrDZ7RntSAaKGNQNWC484kDclLS5CFqFHruMPgIPMKzRwgbsq/CgI
3RHs8a+Xx6c/l1WuGtZuK9bV29t3dRv/03BBa9l+jH3OzOz44CcnExXZ9sC8IWU9
qRqxJBqoX1pw7XSGmi439YejJ8Dtvcej8FM3mM20vdaJCY2N+lVVcl1+fH0BCyTW
Gzzvl7Cpk7ghm9OH18O42PWYneeYDyoW+G1QRzasj1Tti8JZM0Cp/tg/n6O/p4MS
azFeKR7sszsMxtQqCc1W70IzgTGvCrGZbocG7wGiRnFMT7SNnCTwOBEN5THkX8br
ffZEowgQ4hdoqxXJUrlK8eNSYaRefBBMR4qfKNB/osQM7yfxjxhsm1Sy8UFBFffQ
dUnczqd4Ql/Un3Tvvxl4u2cHgriwYJaIk6qBV4o6X06YcFcjrJoKcGPVko8nvHwR
gUNYvorMcfndxokezF3/5b8tQnpepN53u6AJwWUb7m93joAvLw2khGy9vASN8wuh
YzsOd1+4XDPXIH7VBjGui8IB+kj65TOvJS4zlj+Ww/3EwrQ2sDoEUXBZ8tYg3Bmv
8fjblJPqa003vpe/7RHz82wW8VqOLIz/UfvYCPBK4Nau7+us3rDJimjNMmKZBjZg
UngOCys2oqYXzadAEQsfxabwgsUoSN+SvQ+RK5YSkt0gYgGy4utI0PORXymOwC+k
9soDWE2EbPD+G4BYM5z7NKU77ATpwICcv5d0aYots4GM3iNSU9OaLY7zXCcVM6I6
fM0lnIIQTGoVA1LU6JIno2ndp1856KbJULZpAG7Dap3dVYo7csrjhUpGTbwCF+U/
9kXtb3+ZiFCLCn6l/3GsS/YMm9DNaJLx29R+YUETA3QtlcVW30xqPjwRxBeFIJLl
vK1rMfWj3PsrCgqZ9089EPZyNlMP65EwOVXQKc/VP5ZX30oZjdwerJztjVLDiLef
neZHnQXXoSSmXz0QozMumF34cF7QdUfN32oO1Vylc8soFxJ1BCBJ0CDoSmUqPSSc
HhTief+SmMTGnoWHWriPzXzOHpdXYadlxd8DkDE8kU96WoCHD6CVDwMOAlXEw2+G
FhaVpWcb9itVguK4zQqaAb1BUDe7iJc6uz18Kep6GLjKi3lRyQgNBmqiKDGRtRml
pJ1yQ6EQpVuqIIp+V9la58rpoImcQMFNMoBzYswV+QoRCmKAi8aWrFHSbfVgN6O8
X7oWBcEhzvW81D9qUhPXbpHS6QYEC6z1lUBWdEfZKn2G917lgGW0znfVl9Pcroai
YVmnM+Kl5qKoFm/yGJoWzTaEvGOO86BjLABuZHlWmYw7bBwxsCyFhOiHRAIswIGs
pX28bpPl2+C4WoVxNENjXFJF+QXLA7Vr4oq1xxWGQThbZ9YNRW9rEGBYs5jzx20k
y+DarvAGww/iu8GXG4mY24Kllp/VHnAy5WgF+9Q56UTxSpltJ+6K/o2M8IaQJ14I
AikUZaBIYosduOCj+O/8Y7IWJMd2p9jwN+3IKOV2bUNH4B5hOdbliKRSsz4dcsfL
6MGLtJi87p66la9fBbIXbBIyJ//RSe1/QRCt3+wKgaIOxpnZZ9Gf9VMUb5Y+HG90
at5XEXfPe/ZyFcm39NPNDSuxmxn1Au0qbkGhI3CBy3EgGjRpzgjdZ6sOEribs9CS
QdOhILVL4hJHqxsIqRd7AlObyzAQ+AXXuY+2X2EQ69uKmrnkR8DC7hfv9lb2i+Hb
ePFzTfMcrUTGpjFCsielZk6gbaqIoRvClemhw7DHFepeMR8cRqMLOl+pPw8ia+Y6
NWZtQFovBi05lfLeM1Y8/AF4zrKMClajPCL5B3V1fFQLJXkcR0dh3h+9QgEJNu1u
qEXypgzOz+hw9Hu8/kdTUfW8DLsNyISXmAtNMJqEwu9ayXbPi2U4Vfh0iaVxqDb5
hQeMAdrde7nVuo8hJF0sIkJiuXz1B1a7nsWF0WvNzbL3kUspQxLVVJIsHVVYgkxn
jsuT0yTJiIEnaCtOP15iYY81sfawvcC776wgt1FF3PRzVjh0iwg6uiT5fJEXT2cB
mGs6R9Wszo7O+mMcZ9sisVfd2ljSYBVYZ1PVSV2GL8KgNPaJrWDW1VCcxKbwEvXu
eKqigaUc8c0YjbfvEDCLW3tbLs64j8aLgWQE4a7kkQbKtO4GQt6W1Nk46pLmW4uQ
Z6Vj2BJXyZmFGpjso0drfij7QT3zbdXZ6F0dtGttP3nbYa95wrRc3/6C5b07p2Vx
nix79jSBskVg6cuBZSzIRZZ/jhWADXXGKGDXkvfJcd83L5Na1ynwGjLoTO3S5WUH
fma2om/58jq7gJWkRLfRwKue4qr6kO66UPDrJpAtbvGMtzSnxpGNhFWJ66ZUJtPx
1wv/EPp9daX8J+sA5G94faocWCWkIHdZoLoC9iGJiBjIga7BLgEiEWdekrpon6de
S22UtuSSB3jmGp+srPow56vYcUng2hagOoJWvI1aXAFlHgRCq49B7n976as6zGdl
0vyi8byTFPdMzLyAD5/Ld1OAkNlH8+ZcUo15y9dvHEGfjXPB6fw8qUAT/LHEpmwZ
buygM6Y9mrBCFdVKRBLQlMaEScqKJoaHISb8uZS5Vswcr9iMWyJhgR8yHlgVKUz6
xVpftIiA/XIXSu/AvCai511kuSFiZcI3TllV9lKMh+sqCR3t5vpzD+0sJeDnBdUt
fidxNnBbRc0hX1FRZqxwXDa7qubjtPGCi4Y8aCeBaOKLqxO8dk2qhZcMaenI85Ze
GUbBnoowcx5FS6vbEDsLdtIXfIE510FAozd93WxcMzkAVI54v2dqC8VRTSpA5Nel
EvjYN2QLe9uJd/j9RB14NYYND3YdIOg97CCRTdUvynunrQS708U51FDyfZ7VCKKL
YWR2eRflhYFF/bm7aJnUok7Jr1xlyWkcFVUSD4PG0EAX1ntA15A1MssPxHXr6Ae8
Tc83q+ScGCQfSrVeBqeGX0XVgrN8EITZpB2YpU5nPdfpqShwJFhokNqo7JOo223O
enVol3ayV1vY75+eOzNOyjQBvSj1uqsoQjpCx1HxHDfA4zqF+96f7PXl+8w2IjwF
uZoDO2RGWlN2ujwYfdZN+lT0W49n6pF4vZV7b+zglg94NoaqtZx+1UZF38FT9wha
IaypQFLqVlspY1O6BH10kBbnnexDGBwXPi5+Wa0DBf8OYXVU+P8x3K23RpFxvoUc
iFtgDosCPa+wDkadsqAMkFxQKLZvKje51pYr/oa4niDOYcx4pmj8uoM8+3V7JRK7
xP+gdgoOKZuQKJ5lfkps0jibrnr1tKi8M5wpxNqcHSNEssf6qwMKmTOMDt6w+gSG
EvHydURPsmzYoRpliOTiAvmaGMfOMaFLF7bL4l0EZawdi90eXQqKK/4K20diZkSR
3yEjAvqHIIVFwm6k7J9NmgnQKswTrpRt6VOYCm+ur5gH88vI6rzAjEz0tZ15eNo8
sKOyDFwoEjYlEoarICFehrqx7tNWqu+zs64sdPw85WW6uwX6BJsXByMY0+j5Qdc/
nmAkMxw5ybSXSXNdRDOHu05U8OJbystDlH3f/mkhnKtrwemWsTRPB9gDrsp5KXCm
16MQWjNaZlVVKks/f6MPu25QCAtDGwYpj/4lMXtFVKYn9OIzV3O3KzfOanNUw4QP
OWcBhCtdQDUvwG5ydpHrsNrZNuaa8YNZQ9cSdOeq4EwRYiNNRY8B9Npt9YR0EWjj
zrwd6g6J7JI//K9Br/puqZajMrjT6pLnHXT641RUUUvLfvgYoh3m0YfY28sGJotq
ONrfGHl6LI5z9wHtY1dU0CQyxfgSGhvrKVH6xc2Ju5kvODBExpy/Rdxh11HtkCBt
8i9nCSjv43I+x0vkZ4TchRNb12FEnmFHCNu0oL0kxFz4OPAQlXy7jJNgxcvw4Cd7
SV4Ju1ND23mS3/L2Qcn3cLY4df58hTVs9g/7laQLyT3X400DITiDNEpCq5a4j8gJ
ny88wKhDDvb3x9Eqbz9wyFDqrGRgg+V07sEcJObLKC4u6f7NzKnJODR88yOi6VDM
TwrmBSpuqNWlMsoADNboRGk5kPDDP9x5D6mr69olzCRY6lhdxEnS9IGUbwMtkdv6
CBwndCNNvnCqb94t2QPBD2udj4bSibKVnAVB3/EutL2jI8mj/BqPWCA3McahY414
XetmZxNFTLM/WDa53Lffa5/iB+KRk23INZIy99FLfmNHPylqivEgKmsM6J22ThKY
ymZoQFwbnhSxLGyC5RqTlCYUvzv3q6pxyWnnxM+fVX2LFKmv9lYoHvjpOOLFGIzC
cXQs8/CazcsPXum6sr90oMunHrtyrxlD4RLOfJnkJXGP2HzX/kJ/vDx/tX2VEhwJ
RA0ir0dzbp6Qg6nzTVY8zMmrLaG0kJbk3sqKF7tuxufU5sxe8k3hHKrEUocrMIER
pOoAMczOoAe6GUYfMv4XADIC4LkbsqIXrPagbFiJGTBHKFJw84JvprQUv7fr2hzl
Oo0bTBeXLZ2wCUIz+jOVwSxSq2dv9ErLW3wolG+e1iEQN0F/VTaOe4ZsbpwpnN7V
pBPkvZCoMldeSlKJBuTt/KDgEKvphb0XiTR7ATvYEk56G5B6C5uKwhI87j3Rwgzg
+6e79+OS1QNWLrYYJn2gKF3m1yD62F/VhT0mc9fj91ObbSxCf/hIUtO0z2H5+qHh
bsLFAXNDqkz4MkethCu6hCEQJE8cIxFuCmhQGXHEvsXJvtQTRmKo31+bsz4ejtKw
r4AnntD+THQkZUeS8uM2scERYj+iB/8X7v/kIlYpYYsfBO6S++EExkkiJgDRofSG
vhyah4SF3xCB+JWNtPWvtzEDLRup9Fjx8cpL7jhbmpxIrYkoAbnlFNuwWzKtyBFG
ngpBaNQzDjBnKiEpuv59CW554DQd2kGQbOilgV+4Ni7UxhGuB1sv1mgEfOQxErvp
YzagfA1DuNm86Ngp96yKArJmprJ22LmQrDb82rWGsCcsQRZLp7WjTll9dF2eZlXF
k1mRoFaHT7v4uaZxhY1G5fXG+aRmjyZhhLsSvfhoqdQ1eRGPA7JzI8/erY5bP08g
AnugBYMcIorM5deelYD1o6Y36PcyKnPn4ftaduvVq/h9ngvmvBZvkN3/nx085CBv
1n42w1yf86RP3AjM4TYkUQJ065akHULGfJGyCTYjm9uSjHweyFmfpGaSLXXnJapk
0sHp5rIU0k8fpbHXoMyHCRwEaO6w2qAyD60bL3pVz/m20ip/qzYFc1aRfuCmv71P
0IPppHUYokYP3AFqSfmQ8t9OXvFR0zvpyaPD2CW//gzDxYxuYz2Y6a/iOsYF35p8
CEJXTFqSRxz4ptzLK3UVVEMr/8kS/rwTW31ZoFr9cj+BAvx+4ub9emFizhcxyPcQ
Exl0S/z5JVWJyrGzbGASb7NdcQS2sV2KAplnEvOJZoQEebKfZpJZPLdy3LQzaCp8
c4K3BzooN0g9Nn9O28bqTGziELduoFd/vrUl8m9JqSn6FVfih+CCiqaW23sG9Hgo
uhUPLgvZgPIIZ3UfpvKy+elA/lH4QDupMDAjLyc2pblm90WkVvY6Uq4tq1uxtf0d
O0gMvBMQbi62mIxT3K5/GnIcGFjcDGJ4itBoMvEbPPHOJBucI6SkpmZ7NvanqhAR
qG4evve+KM1kYg4TYE+sFChqdLDHL1sUwIViuDHeNb5WSQrUnm5qN+Q5+YU7BONu
GNE3nV+8hjW2WJfNEJ0n3oTODC0E8sm9M4wBUFHrkIN0c5diFsP8ofHNU7VSmMqZ
PLAAZX+hwVK8BHxo1UzvY27sdKvepfFVKMW/zRoyyDM/9bKw4hUMGCB+lBw7bUZe
s+WS2434WAuabOooAAv97r7yOOdmtwMW6R+Bng6fReH78JKlAy9t49UCn1KWrjzq
vICJEB1bO57furkfnarMnqhtITZsPcivzfRyurQb5RB1oH5NgBu2LDMM9oLC/a4f
scKaDynYYcllxRvOL4eRMIPf6I6gBO0PxIrgvrT+ULYfpnXkBFwYFw7qmreyYdrO
xo6nv/vr1sMdrEhZndt8lnF3hPi1bSq5Nfz7+P940Kctw5ycMYkyfeZyogSJci3j
7Q/3ho1Ms512elJ2ssjK5L65R7VB+Vs48kiSUHikw2Ce+5j9n/u1PK4hdzMI6Zf8
j5Z1vMtnj/2THpzIhqv/fqm1DAGEPdqLKUb67H18Cm9qV+be6VEoIMixRIrOn9SN
6bgPzsvr4ftGd8nmVdDhYjm/oR6XrWv3XB5L8z2lwWDdjTSu/z380FY8j9AnBqoz
7/THz7kBRl0b2dq/tYU7aiBp4wiiimR5+5+one1/glFH0UEZModk55DdjMKC1/RE
n9zVTuiQlSH2sSpk9Ue9Ts2A2/TEjtnYJDedmebrZlvgBnGlTL88tWnoHskdTBrf
JtfT4uD0YGUF2vIg2o6EIEeBdHOkI5FtVMHedhBBe+YOdajVfSKvaz1xoLLaR919
inHL4IoqOZfwdCS5BQHYcEJfXn6hmhsr3TLaa0WyylTtcv8AulmJmfZ7L6XctQJy
IFplhDGyVgzONACbPOE+hOfJ805DUxltBmkC9Qn5FYF+4AzoHOxERgS0BikSB2+b
bSQfKHBerhrE38eofJpH2kxaLSSgykfYNRVaqPOtURN8M5N5XmiXXq57pfdVMO+F
+ohO9dyM5/gURB1rb1yyjtiKXMq6JMeOxr/sHdDKmgayRx6ROYqBjUIt9wlH5gjs
0FsmgwaEpt4lNY9Zc70Be+OtFzqg/8N64ZwT3VL2ZljmeaHQnmFDEokb+N7JZYBI
8sPWJj28Qpo4E2WKe6Pvp30MdtXt0Oq7NWK1ZJI3Zr9J+wKXcSRwLLIpOI0/SiYz
qZ5k41gZtacQPR5Biof3FHQxqnsIIm5JUJW+s3BOdGlHICAxUce9d19Oyy2lYH/Q
uvkiWOYIUojGYrsIhZjFBqwcNYfqps9B5U8OB4dawkU2SoYJjty1gV2FMXdrNLvY
zJuPcMVdM5XP0r9k82/J7yxHNetCGRP+lfEEnF8iU71k8qQ2vEPqdiul142TtMvw
NgXPtHgQzV53n3vg0fU4rYiZUFSCP2myJNuE9PV/S6BHUqGKtQMYjTMtrY68NVJy
DMPo3WPiAFPYPTwp0PjUmhFX2FmCdMouAmc9k3yaapjPwHJtG4fBfad4lSJ9H3Ay
/EjdEdDj9qcNZqkQGoQzrGwMyEnXF6zCeM6ilJCWzNcS8Qx/MwumCkP/GPf6y9wj
gUlVgoXNoQkMnemqo1i/+h0R+KhkNqh7JFCHlVw7HpmYXwC3DYj+E9Jn7HfGC7ps
MKxkXLGmpa8fno5nxt2wc6w8cok9xOE5Ex5dlIx3WPoJBED5K8cfi9kXTR2uh49T
K8OyHEcnAQuWtkvE6BPdqoWIwn2ADhc940B5JglMxz6q2U9vELk/zxcJq537TzfL
Rue95iYMmdEeKoMyMVNz3R/tSnf27uaEfgkTKduZBs3DkN/BAKbMYWHFQg5JWAq0
6kwqULVfraXKUSm4YycokK5VhByTdv8clQ5QXV1rMhFsZK5USBnd2h3QZxHqYo6h
u3bwToSjWYnT7VuFiQcRI1+RJbispnU2ZHG2FsFt5TIOD5qTzQN5Tiy7t8Oal0NW
5A4HRVlrszuajXmBO9fVXj1ywi6MOls1mMGbXPTHU9X0+24oB/cAphfb9BBCKa7q
jbFbfhenIU9dfe5QfmZ5qFYCxyFrobnNdEBFGhe3tnypqwmrTbTTDlt4+fIH3pTL
IxAlbN6rezhxX2GoxjxatSESpjOoWEGOmrz12sL/zXm2WX1DX7Faivo/TuGzNKTt
5jnirNZcOiy3spzwuvxEuqsw5/0LYS3aPVVMm0QKhYjZWOoPYsCIwYlqsqbWx8rE
VB2Ls5FKJipTVzZp4CYvFh519VqvJV5Gy1Yk9XS4PvXcIQ6QAz9o9eYOck3Pmjv2
wSy0r7/QyEi98at+HxqCIccp6FxL+DK5qR74dtRvt1p9DqneOfrdAfU71xL4roGA
5ic3anvr7cyErqCdhD6YvnS5TekD+7s6vQavh8Ygph6DdCASlt3v2twsW1mk3fPk
08EuiXfdJ5heZbFqvXQqyzDV7ArxReKaLJHko31+io3cYcQzmikRjvg8mW1q6Bhg
nH61oDx1ubBPm6aWwoMatmZDQIOqKo5K/hCgNZ4Vhu7jOLOzHqJkSXVMTS0pQwNG
yjMOCxsYqsibZRJEz1UCIAhc0JAfBHqqsPEIAke7aD4U7r6U4pFA5IorxKxcRK3s
SIALEmEaj7rXDFVSKINJDIzPTVwW5jg+81fXNMTFw6R1Dul5r7ncqxbwB2jy+7/4
lhefnnhble+Sap/SfnDiqrR+fdluDlaxf0IAXF4SkK1dFzoRnSBmZ+X+2LzsJFIb
ybyH59U1xUjDrayQPjRGVEgEEnvP6/MXYLjyLpzt7hJ7xY4otNqPyzO/tiDS6acj
KVf5i2szRVLRfgzBSClq1ZWbsKuxKAC2wr0Mez/mOWc3o1rJ1+EwiDi0T1I0xpum
4884JD9soG1JC6WyzmLkRfDtIkYmVvHDVK+rWc6rRZXUUxhmRTMT6ePINN+KFKid
RH5z7HpIIRMbQb2a1xgvKW2Tnmc+LqseEgqJQGcMfuwky3BLlcqskPj+HWK08a+m
gU6Yp5aNinE0wqF+2KZBXOT4Zduek7Ek4iQbSfQPWjmjez4PrUIJpEyOgYlDnt0W
6kGLPes9oX6A40XTKKyAZgd7WYr9SV46Qa0G+fvPELKtMdd0ElRmR+pj0pNmujeM
1ZvkXmmtHpvBTETvBBUc653OQrRx6WOeEEmJIm7FiD7Hei4sCHqwm7EkBN0aDH9V
RF61HLbdtOT5SxVKBhPdabF6UT6SWvlVbcYyuUtO4woF2AQ2rnxSFo5/cCpU5UTW
R+R17rPhm6kINBVva5vegWf0uYs/j3eH0Zx3HbzX+fTU3LeNUq6I9n7x9cqY02tX
foFt3BAl+bLkhoqsuJ3KI/Oqip21xnl/fY37kfP7lbMT0JhaOGUEBnJXhQsYselj
KTbO1zZsYw3HOej9Vbe4Pabx6jPUcULehyptV9Ge7/ahv/6COog8NHU4455bBAvY
pUQrSJr5KblfItXb8FppFHP3kOcsh5D2B99WItm17NNxj62XC4wlDK10X0qnyaKo
tBxjwdOREXFVO5L7DU31ZD6ACTk6X1RPJIb1XNqOLh4Gomtip9bnVFDwSSnkZMAZ
W2xOq99ulPlaR2v3sIawIhCaUcGxm8n167/OsPROHAgyWlVV4+IQRm0fH+S1lUoa
ZcskP8SUgvaE1hMeswYVNhwe0G4ePg02DtVCGqXKIZcPWMNGgDR5gPxof5fW7xY2
A4xGavSRgaT9gZ58QorDQSQ7L2GGZem7mPpkI5vwduV9bi6FtEcKusf42ComjiZL
Rj5EOJrkkQiaJ5uM699VAGrzaoWmK3WCiUJezH+OLcUaPIjHFHmn4lFlDz4yq+nf
GAeb+9OqZlU5Wn4YkzihqwwB9Qgeppv+ROrJE0MWha2yV2tOg7cR4OJ++aoVGQNx
bWVTnvLEwcGE1zhdYk49c5O7fohgGFc6BgwbAiyyA2zttXJ3i73oQnU/CrCZNJ/2
E7G9hS7P4WckcvLAyf1/Mzgn7a311vRNHVnQVJBr8nqHNGUlcSwxfV+9c0aQhitD
nvO7ckgi46vJEj2VfuoSJbELnc+ybE/U0vFw3dZXrrgCfFL9gN83+uuI0pVAUPVd
iWfWN0QH3UKVCG7aWBCxvwXXiWtD0Y9HOKJtClVNv3w/UJT701zboHIG/g6YifGy
L2lQ3sfY0zIxywppLDDCppDO/M8BwAFE1ZWknpkFO+mysJqXx5k2ETI0vtPo7vdz
9yUuWuriPOHs05WBDHdar0CHfJgGuqMJVeIgs9rs5WldYhBGCJiLyS0wWHwBKZ4f
dPr0YIgBgwSDje5AMTJTwH2OLGoLicJ+p7w+/ywj4klOauS1MFo6qFcBbL/GICw4
HDo19/qY9GcUCOCabd56/091MiChgG8RUsfUk4eTzi+4RvJ1yF20GxbEp/ni7o2A
WgX/yDCErN8rXevgAYZ/hVvL2P6C9C6+CP5qp/Augiq/6yqAzQJM8kbX5c/qr2OC
NpTlfByrOC3GmaLGezJhIwWDK+wWjXuurlD3mCj6sW37DF8s/uYaw6zzwZ0PTmFy
pVkMa7/zzgzgGXJu1nA0UEBMgkqW6LqIZFl1xj2+F4BMQmZmNz7zYLp+sNzRVWkS
SYmCt3wxoQP11sWmf/ns1j8W5JFuxThoImHcd7WMEP1Mul+06eBsZUOxblnCnWhc
Y/UA62ZBrgpn+qgARS4kik0ot83aBIP0wYknhQ+QrUGf3bflkcZ4Qxv6ifk6Y3IV
atIOCwE9QJeJrDgnDhscoc6BYeIpmUBWBIhtL2z1Jf2YRn+VvtgOQV22VkxsoOw9
s+bS7GWlNR7L8CO2u7VjjXXnzbTe6Irlwp/tQ0R/zEGGAaY4Y3CgYPM00HfMlopE
H1bSGwdmV5A55RKvkAto5C/BrE/PDI7iIpiSIJiavfXzUcrbTi0UzjigdZfypV8A
Oj+Cr/6Wzsz6iJbHEXkUZZpCtVfb5tMMRwofwtL1fjUdWHGLLmICKvd5CdMBRsqQ
WX+EyBh0BUE8GNqpKKri7LM588N1eZsmmhBfcmiEFW6DpuNwrD15beftomuAcoRO
GJ4PSN+hRzP0bw+a7KVVsU+MeITJgNDz1y5TSHeGGhr2bMjqDvSe7jIIQp57N2B6
2YPHMLYik4jsLWXIQE13b0xDgee9Bzh6epRtoIsBLEX/RXTfwfNdqozHt5xOAawp
QyEo5zRZs+2XuIXXptrL2GijkTdEiJReaMeq6ugiCmrZlCPbdyYBIO0eRlC/EwVQ
sBj5ztNYoGlOy9hKvtpnT2kSV6VnagIfOZhbifOONfDPpZCvYwZub6tX39NL8G1U
l8m8N7dNVJi6hajIM7xqNLRKV6oaC8/3tvCfR2WrgZyBw/HpGu0OZZpJxWaIDdKT
qTt9/7Ran2LCJQnO9lunOPAhzeOMc5rGJZAxrKLUi25Q1HntxyiCodw7ZHoqeLky
Ddujdg6IcxvCeynaomI9GJ3iaMrFqSgy55OcFBEuNYJGdUN+MwMDBS6gj9RiYlfL
mmGxzCQe5657FG1b7Cm/oY2jvUqah7LoX0dQ6qKvZkPxHd9rjGvJgIxxuTV2jhMG
E3n5l933q0wtuebb7b/rSAlyooJEAPd+Z8LzsWUW2m/mfaURdt1kYpZ3brTYGX2f
bQx9yv14bhhrNLGklt5RPfChLaKhZZhZqh8VuMkWjJPKDk3NkxbZ/H8U9RTF6LMQ
8UX16yazFmAFwbE9GUryYXz0/YvTwckAg3yDoi+S52iAV+sFF5rK8pNPInQBeo6o
8Bh4OPiC3mYemvSMaMUwAJRpWOzRm2P5OQqEOCxkrESRiDvX2IRx1WbT76T5V1jH
QE6X9sil1djU9LxC5mwhm6/RHyK8KxFP0DX0f0VRgaWUk0mH2AHGV6L4vhrTKhqM
Ctnem8bJhYjdAirscOKTFsbNBwIbYcibgtuNGC8JZydujg+S7/WZ2fl6yJdrEnFt
owz+fyNyUEqKGQGrttzZxD4lWEDMo5NOkHRIYYK9BgiCqNj7NcQBenlpuyPpKUlW
5aKYdJVw0JfBd7rhRiBXlZoXGKRIJMHwGZxSv9K7gnv5QndB4dk5l3BiJfBuLa1p
85kYY2bY6TZJwG5xlUuxT7aXbNWtpASPE+3fmTfN9wua4ZHx82A326MONyfECSpG
g2cVd+tj5/LY2kSeEpavEtp4oBXZ36IcObxKe+7iSxQ+4sDrjM2thGJKPSdsriRZ
8/EKssNhEsoiB4sh3K7Uu0HLU7F61ucDuOeC/5EUsGJpjXODMF51VpWZTd8tM1Sk
MWemhP+fuTaXwVp3BU7URho5JxxjRDqjHYEFGuGO2u8hab7zXpEiXTvArOP9aPNa
Om0a47d6bEK6+tTSyPpebyKwETk9eGx6OJfnIqcFY+Z+Fs0S4VS9N9mfCfncJOQ+
p0mP/8NbqtR+Bp44lozJiXSePsuqh5GrA3AtR87tGYzGmMVQ3GsksBIRmu9Z1fTf
1v9D17h82JqCgsQOgub8YnWrx3vKrZ70ODchmKnrr64s8p4H5uVviHrSgtAFcrq9
modtDBOjAWHyUBsmX3wk2V9FgOvo2idlz5Ra2HQ9GDOBTmGJowDWUO55C3y6N8tB
/Iwmn4kLrURSCWKKsVf9zyjbILhQNsvV8HQcX/835XYHdAso9auWcuATGBXyfdkD
ga4EPsdueXtGjZ81vlAb5BaFHoBv9HGphgNYaZ/wZcjrIROVWEYFg1yp7KeXHXuL
DtibzORiM+NvxER/NK8IJLOD3hLWeAhUvexbw97apsFOsS/rcKgtZbPUFix3EY4V
AsDi2l3PySpBYsq/vpnzZxHN/CybpmkboWU4kVYlQ4URbvobjgTWcAfQ7oWaFf2r
63J/QK8ef7sYE1lTQGHBsJ2h5vV7ipO9iUXB9PePjT8L5K98eJQUFkkV2RR9ouxP
8qCJUXyFn9h3zOC70m3EL1mO8phNBZQEWHuK+BmgUgeHOuWneQy2b/SSWB+xsyFq
TM+9E/PDY635PndwmxHiFL2xoI1PG2GOfqzXly04Szmma1zJ5CFaXTgOMdPHwQIh
i+tpJh7P4WCIdyfqHdlKZfIid0gU5nGNUN+7LLuuLTOllNTPqsx7rJ7ByEqVNpY7
Bb8PdN5ia3uJulGdazJYnvFRS006SwJeDhK9CIqrifO97UT/rAS1jBssovk+1XVW
N99/UZvTCxYoNOmb3DRoYkVDG6jpnVj4s9tVhaE/xxZjBryPsE1rdTF93yIQH82v
tGRwSIG/pe7b+fncUAd8x3H6rG1QeBl9ohEsynBYuEjLQWy7XWoXULBN/+dm/+Fx
gN9JfHGpIVnZscDdRAU4RtLG2R0yx/DLmnk1XV/KVHuvAl3rkOP2zrFJtJxIISY/
sZ1aMohr1Dczb81Yir+5n+am3Gvg1Yp6vcbAhsImrwpiuNJw4TD0U1tAs5ZTekJa
bjXx6+72EcVt17z+qQEzHIRWdP/nqzLQzIGcwdmwe+MIfybG69BNOy8QbiyLAI5f
q7Cbkdb89S6lySKNDluH0lUq68WI3QvgmIBW0dzmVAQhK2xs0xVnE96RSQ2ygfcp
SxxMiTr91G633GHnyslUktUb5I5YANWOcY3TjFuliFIlosJhXP168Z+1MjNt3TI3
ZayczLpJl8iTIgh2kC0O27tdY/AZnOKsMyS4xYC3XfNuilnTpYu5arytxG7+FWqQ
RLwR9/bkwLOW0/O3eFrT+i6sXWznTUxRRgi4zvd225NW2it+l98o8HFwIyH4aJQN
yOsm6SRLvBY4o2DuGuaQI1NmEjKsvBbFgl3YHuE4XpwkaI3YpMT0L0oiSb14ijmR
97/A01ahvUDBL9mOVyvf08MNRHo7s8vG8Pws0QLNgCfV79+aB0f4D6obPi47HLaH
OH5rzR/h82+9J9R4nxSb0N3s5qzRkST+ix8/LzHQBvuQhAQyeteBOpbdQv6DByWj
H6akhNu9P0I0a6+8upOvjw2xem4mRDCTm1yB/ZbEUgHmxpOYPxMY6YKY1a/7eFpl
MuVagVWpc6WSNZi9tEuJFqh82aJbQHOn4L5dbQmqot0jiuEYuDltBBnFKIYeiTxz
kD0baFvnxd+TyhUSobP2DYenu5jbiBLiW0ioPoRMiwtsWJRaF46oS40/jeIXiS/l
U9vzc3ptleWgJVoZXeGtWJ6ASX5V41d11yQdLPy0DGt5NRU/gb2SBHVr9m9q3RqY
soPUSM/TLV220fj77n0k7s3Fix4cq+eq8UH5/H6jP2y5pGje0ubHh4b6O+R2UUc9
N3rHKsTF4iSLJ8cugApBRSc/F4LN7z9E0tbzK8qK0Llfae8+DQXvubgZXfCk6+Il
Hgqvvx/MU9oIJghYJspkHb+DgcYQEGrMZKox5BXrKowJEI0gSJlu6ljYMeQ5Grjz
AyMSTJ4TpsuehRhZCXUb/zRqocZrxkMkptB2Q0jF1uNXtzir4ZIyx7rF/e3zb5F3
MsiNL0um3cVvi14O+HhTYWAVG+qzfvkwa6czr+jGXnx54fvQlNrSTUMVZznhvlju
rsuPN4HsMU8CU341+m8uywFcEsYNKQh51Wv8r7Gg7SYOD3L6uiLd4FTAxmCMGo3m
IErBiAAHoffhoAtqRk2f8LY1fPRB7hB6FXIpSfi6v73ex+NZPfXo63WlGj3iXnVt
TAN+rmZqDjJDwXWFoSjx9lmKCJAS1H71uAAX+UTQFynXtW+VKvk3HSDaBjUg/tS9
lXCjRBhtcvzQI1IRJMvWYNFr7m8xo2sSYSP4oI7d6J1TzeDvtwKGdMto7T5hku9G
j8keO8gIByvK30HcMo3aiU8spVyiqpS5JvNnuq/xK9SaupW0yKQLflZ8Bjg6qeEn
bGLkghnfIFtjswRkNLfmCFcl6Rkf5/ccVcU9EpgwbRqZq7svMOi3AowVb+WA7G/O
xmlkSUL1/UHv7tVowNJesyoEJnC7xZ6lqxQqxjjNqDinTRWFVB07/C9QO4oPqsKX
57nZ3htQfXQrBAn1mmNS8hfvLWAMslaCRf92EhOHlnp9usrVvQ9wWm71uXyppVQA
O8AB4VG8omtdp53JRQ9M/6ztZrSqmZyH/n4u2FKA0iAEneZXDXIL1RPXPPrm3Obu
qmvYZEXBpzHwH5+z5tMd8ZX0sIuCzhNc+v5zPmX0myU9KV8B0nOvxZvoFFXqmQuw
4/AyXTpVkd6xi58uRxwOLQzvmA/G7S+azamifp4j9HL9IuZQBpF87ZF0xuOqspwp
5jyTrOjw5nkqmGosefAGGNfrRAPf5dXI33dWmYO6aF7z0AYSUw11t1iB6avfmD/Z
W5xAUGhXg96GkmtcNn1g7bqBQYDpLQgulmjmkya9Jm+RlONIzU98zH0Gm+bTsLPR
hkdEgDLxAGuVroG1S/0IKMmvT0ZVoPhUaE3nG+TDRRwGdIHT4448AztAdims9nOh
pt1OsIeezU8dkAl2qqF/4YLAMwM69g/ewPfO5MeUNw66Uvsz/2dbw2HsykE39NF9
vpg6CsjIsJ/xYpG7BSGR/gjbdxFMWAEFwLua11xVgQ5V3Y53raU/DzILFeGqJZ2a
8+dC+pCM+1AgC8SH3K2Qhy7pTlfiZO5c+o9bho3zyDHaL41CBGxe/bVYj/tnDH7+
sYB34SqWQFSmX5pFtU3kDv7LctMEF1IcY4olLsg0kUPGp8WNjq+e3OFWhYTvbu/9
EARqs2343gZqfi0OMcmFnJkRXnVrEAAbzy+FiMDBAMr3nYOggVlWz6keZzJl7Fuw
EfmU5r25V9BmG2Y06px3G4W3FtVbYj/WG4QAcpiK+N/kTtJZaPDvWJMMY/xfCgQK
Vs5b9wXoiksfCFwQwzEfe8YD64ZxIac0PqC6WvKrdWyHGgbI1cqXOxA0lhbXEjp0
UzQevdTyasY1P3FGncDcGGvjQ8Htw87t7n3ZPvv1fBhhLK0X6Fohaa1zghu11x6z
hBBmKjhy6+NTAZ1JHtr2D63athaFt/By6EfSgTVYfglZ88pV8Z5qpQKgdz5d76yi
5ZNtADT9KqwNjf+KoVK4s8FQAVIPV4yaCdQUtQoTi+b9zCseo7EL3RA4Rf3Msizd
cBCH3fFB1dwdoUkTNLxNFQqArHQkutARobGlp3zevcg5WNi0Vp0vPsG+HawjMKsy
r3BrGLCr6nwD2NB6PYQhMK0MyRiKeCTezW6fY4Y9ReTKzBbT7Tn843ddHnM7FYYA
k2BJz85aM4Ql8bWRpb7LBIaxgl5rV26B/1EQL+zal1BASr760Z7KsEIuw1zEzKHV
ZrwKA3ojAGy4kcaII1+wQzhIWs64LTddscne9INTdLYG6ug90zMompRlIB6jydnd
pnf4gtdYhPnD4v4FMvZUDskblDnYDZeO0oHr3N1FKrDJFV4mSyo4wfGzhzJ3f10H
IKKhYkA7rQqMqhOER8M/ReoznrZijzp3b1vT7m2+poXDkS0Y12JyDQt/dhMH3Ttj
DxGRq8i1NAxhWJZtnt3V2N3Fd4medfoSGZHpJHkgwG/iHgQaYdj6qiDQ4w7eQqF4
FE3p5Tzt1BMCgF0yyFDpMQ1ZD7Z22TOfmD1l8OBX8eP8PsTjzCDHcseUBn12Uzc7
xdouyn7crMmBy9cGke+9J2pxGVY5nx0+LQ2NbQpRfXKKZDPOFbKxKb/EwnMzNox0
qcbhCi8eRwybDCrcqYjw2YQCAIE1m7r4CDQYKj28O+xfKjTZ12vpjD0PVRXkfg9s
o4kWorOx5i/JlW+123x0T+FJSuufsK5oFVypZgJWOC1IcqEf6WbvbKm93wbcg+bm
F5AgsVsAee0jmKq1Y49KW0N7rLLK+YCuNXEOiPOIBsQrcRn+vhElWOqpeJgFAt29
ovlHXyu290lplEt384oBOeppH5g7R2oPgovO2CN35A+Ew2f1lAb+Hoj9Yx2pAc9y
7BrR9l4QiXec3EBPvsQmj1O3s/9bCcYHEmNB8a6tlUjZUtlcYsfO/BnYKSEXOmGJ
P3zd7NFIomgLb9JAQTMlm9OKwJA4oN6UyI2ki2OHG1JlApD1PBcjkw6nd/i86nu9
pzQAsmWgXHG2uitVSq+u+wTrBisAO/c2u3tx/6kmb7UGFC1RI1Phvm///ZPTmZ1O
FNc1ArmNcxf92mXVyGJU5qqjTagrEbuE2Wm4hKrmMKD2udFxEYS1t0K5FfmCdWty
JjkWegL1ASaTAOOzsTkiyf6opcsv3hl9Peu6pc/u/zHlQabn+7Mln2s7W1Jiqi2P
6TblZX8ng8UhcTQYhMiIaTO1/oNPftxo7OkNka/UNmrd4N823XIaVCPjdQlbtaRr
JAW/Wm4Kec7VgntQF5l8ycoOjo6ud21BpW12fDjzwOdsnXBMTiPWkYiwH7V3vpDs
iH87undXG8sTezz8mqkd9K41c3XH7XJXBj/8wgT/uG7CEM5r5iuj02u0DnH0KEeb
/IeCBqm6/x2kylHnzus4nOmv9u5cs+chDr+fw4eVDy5zGJ+cwweHYmnR40eedjoq
E9oILAZ5kgkcsztaTj9OhZXJ5BGpWdRubQqAneDb+lqlJxTxYQI0ZMlrgZi7Fc3Z
EnctcAK6s4gvvTQiu0ttFr2t6msMETWJz0MRQiYBeoqLpE3t1D0GVzkx3GUgHegF
13ADvsM1mu5bTfeYOtkhiYW1Tc3IAIRcTm3AOAfDeVwf9q1tJEUIvpkeiaJ+ud0t
y4XYFetJQwNnT72s2yJos49mz+upgCsIV1OtAS0Cbdhx0f+EfFkWXgnKiQm+4JJ5
QqmN4aqYTJKpXZafDOPc94kgaaGSiuW3HqS9W7XS0Qm9oChRuT0AioOz1edujBsO
TPoVombECdUQw/fJy2Jlx86iSayY2mnQ6ax/mxd0+cug1XrMIibpM5HTME/nHnnt
KRpnxASJcygJNUzmH+GdQjJfCcPWNpMgYgWHlak1NFMApYVG3SdEZTGZB2FW4BoD
JONyVHOhXYtvi+8TjhSqBw76m7Hqr9AVdtTgcvckDtw4MaCAmvHOFlFFI4QK2I9P
5wGNc83lXnpu38VA6TdJ/s9WcBxorWxNd5fG1jY+YjkSdk7EftbP8qfQ83orWpPs
EH8kYzg2OGa+rxs047XNhUhDT3e0m93mkPf20laCrDt2JbO550EaelEcOVu+EN8P
Bci2ck8HxkEU1xvOdJUmDoYbzNb5j6w4GekGakz8hVhfy0DdVYsq1PqjSOGe7mmj
bRtP1yHd7Ko79TDuZ1LV4uAMauRFZU7TsAM1yzAU7t3Ps0xBPJh6bzqNkr4x/X70
Q0odjSkF9JKxqYfAlkSDgmXV7AueOiVpAu1FZEK5kzigGh2RA0ZHeuiLRVvbHnXS
4RENKnD60PMgG+XGTkR85P5hU1pGijnq7RHRWpkeLmoEuu26sDh0CJtg5S++nlnw
Llpu0tksGxwioaibp3U/8VFrkyuL+kQfuWV5GMw8pQt4FlnEht9Lo3JdWeFMj4A3
Yz0nZqS/FXdPEZo4jhsJdbfdCWWM3L6US23CKZpwvR5/KMayg+V2ompJO0X7Hd1x
gGej1yx+rTfJycFjZONqQsr1c/2+MEPnGJsvivk5bIoSqwnlgOQeDnaGitibTbI5
3u3+TWC7Nus90hdpmoz6fckpGA/pjEY928xilmyVStgqSblqQg5ZPt0XmfwqdNiO
PuhKonaooe8KcyKAUZHJXPYoTUL28+eKVGzqXqEhJ7w7EVOtY6AS5csSPqxVGSpq
H8wsnvcYGmCYKHs+u2A/qVXC6BtbzRk6+h5FdarwgJQl0iRdVJ020wRW4xSVki4o
rzXb5Ka5t12Ksb4aiZhaK+pXZ0K+F+NhZ8dE/KCbEn1ECnbyJcGYSuS0myLILlbZ
dzXF7LK2IHXv31YIsRZfWFzLnvMvOG56V6b/nftDlwX6izMPkevy6w89gWF8T+sW
ZMrNVie49SL5UZK4J1QgkIAeYpUCV0uViZv5rpVKaHjukug/Tg3JM2CJekbUxo6k
iUvVaXXpDLWldkNOcH3S6AK83Lim6uTn7xRGDvWHGyjAuPA7mhwxwYwXu8VWHsNX
LYTNes+hGi4z1G/0rDG0hDxYjJavrQcH136jc1IjBfK0DYg3QK+vVdo/V78wl0op
9OdCuWMyubQ0VrPTaeWwPsQhaU1NuByoD2IOsmBKD2HqRO6C7zQ5dIcCPmzQDDI0
bzOwk9ecgizHe9ZAsP5c4gdLb+EingYv0MxOWKUFRrZ4yFq+4qb0JepBG2hF4gag
zqajcqzvH/JBchoJiX+QLpz7xe3tSWsW+Z0GsMWNw1xS9TyDRe0wxfjyIuroeLp3
a3K23wImtZv7h2nCLWF7hNMQ7hQwONfXmQ+fGH+KVZ0AxyH01Z55ug4zxxiWVlpk
gg6sqfRHTbw977tnJ3l0AWWVUmjhuDqZ6Y1Mx546HyUeg51iMgu34zF4lRyKZnQp
HCe/I0txElbiKBnplCHsvW0ZeqjJwqbfpf9ekKek+/FTV8ohG/LeTUQuU1PRHy3X
ZfKhq2yTA8drQvezLAw0SaU1I+CO6+FWcX1nVAqkRNG0ciHuvrcmlozsQA4705hy
PYE+0jmSF304WLrlxzYI4kpvICujeHSKGHC5nWzq9LVQwbzSwCF0bLyquIA4SsoI
8OSXjJIqfW9Jt+yI7x1/+qfjhU7fr83ClTiAE17PadOno1OxDzhYiSjb7URUS1fS
ZcJqFH7Nh6/Nf2xsqIxKUCkF5dlFdy0kHrgndI9WSfcf+f/OMrTPY0W8ewsneH9O
HsqK0ztXHNAoaOrBBVbFHKqT9cCF7bR6vVJ0dm5eYjrF0H/c0xoHH1x7UlimUFV3
v2W1J96EHPNRun/ke3/gM/EEAk/pau88HGJoM2gXOehhCp2rWmRz2vMo1ngo8box
fl27hApV2rRYn6ld0/L/t1H+5mbOxwjegL1HKovBnBqi/2wbvkhzN6qiv7u7NkKz
+Kf20sD9ILH/omJcdxmJZGo6FrCPyC4Mfz/zvJ6uL0Muki8RlfEPnAkAa/F1gXYT
nHiB+IcGy8LlWB9o4GzFajM6xYkhIQ2uqBJ/bMYo/L1KWsGkhnYZjLD92QQwU03U
UXhclEu2k+VIIgCqYNaDh5YlHkl1hA0Z117MicgTUsBIykvekTH9DiSzl3eiHq00
1krz70mspPogDX8bwCHLDT9XIIsRLB7n90AtQC539R/AUECgLjfygd1yCN6/HjBk
jOAMhaE3QJWXrUMv9CR5V+SNbVP/0t2tKPyxDAzn6EYRMTsHEsXwMhV/auKW70Uw
ZdW9iinYRl/UVSqUB6U645BPcVtHX1rPnQia9Fz1F+lyKna+ydZzlWsClxgU4GFp
FZjTb7zNOHQlvsNp6kl7YTL92yNOTcR+wiOiW3Yt32riJi39C9vBg/oSwLsdAfgA
GhSFaTHD4LeuEchbJY0kmNMlFJbSC6D3vbOSMsbva2FxbGEUrKlbJZ/S6yY+5Kvd
tUonw4e+y2YJKR7IRvPlLmlyiiPs3vjPqd2IE+QqCt7YU0lwzU0TBt0LwT4pyaoh
Qdy0rdCVKmiGLrkqRGf8dObQ2BsRoc4ydJSmhReGvpF0cTj+RG0fl+9rxUkOv5SU
4RYwn1geG+hC+oSb5amrkO9zK97DmN8t5s5FLltqiMxeyUor5TNOLMDI8SYGKoQJ
aOhzAAgA7nRPx0HDT7nQZrpvQAFOZFGOnAcjm5JyNBjgJcgL8tiW1wkI4IhyGTyf
ohUt1JFt0SRahUHSuLWxweFZEsPN/wM+ZLL9XWPHMomPQQTPl8YlbH+qgWl5rnqJ
z2HQ4Gqrj3M9HKnj3EZG7qxKII/PlsT91EPfcnATws+AvVY516HcdDBOeKb4lW1M
hu6oB5G2ZoV9n83SL/jFDC+T7KQEvr6KagkvlOfFpqBkh3GuFsVWZysXGoYVydFu
2oOrGu3N+8XQBxuk4/CaTh4rpOp1PHuyqn4t53qyrwy/I6dOHauqKhjR8lDZqT6J
JUzAgTbql7tnVAUwJXN83g+tWfa+Gib6kvD9j75/1bVa/h4qbVZk7pa5pNDlACce
Np3TFbn1q3oDsSx6WzplWNr8DMooU2FNmTQZnNMewayEY3ND85uMXZsxcT2RI0zX
VcZLLTW5mTX1/PxmxESBr6ISOpw7AVe12iRNEtAAc2u89uUTJ/IVv04gDjTIyN3g
d/B9y1KpRctPuG+xNFpAfF5VdZuMCQw/6ug3S3H8dhUBLyQyAyEpD6HxSmE/DOeo
vqyyx5DrNChbkBB7fgX2bwihVgU/+KAK2ul1Qv55oviR3AHct6VSgunh0WlxMN7I
dI4QbT81ok1gDAxZjELpLEt1V3ttnqiL+DoG5W6rMtxYXlrZkOpaRiF/9/3u4zQL
WhfXzBhaPYqWEs9RceG2s6WFHMWqrj9px+nkXXwGIrsvZZBm3kpnSj+a+GJFXZPA
AoFAN+wg3BUylbwRw8ChZEYDstw3j6oQBpC8h1Efl6D223mapsWwPA2JJlyANS/K
0CVjZqXgUZ8BBra/YNR6tqsuiHjaaamXfOEKd8PimFA9RQBceLU9CVO2Kz3QF/14
Gz5f9tJPtMGX19ClUccFOzVzqxQJgi7CK5PL15XIiB7+JQys3HJGy78eaL+Plptn
g/R3jDr69fznHcPTj+jjrhHvDMuu9ZzhqbFVmAhpcEy/Ldzj6tgqoOzwqZL7oIqO
hKlk3yRTj/pAZIPYs4aztpNIu2jV2qMeSJgyEi9HK/cu5tCULO7nyHF5ESxOHLey
WBMm4YIXNSLaOs4OJsRO3ogsdBswRLUlT7Msga1JHJWX+s+48d8pEZUSd3J9A0ws
ijMledv3wc8ddFPs8cDK/juTQc2T6EVOTkYM9M4EM7/q+7Do7cxQBcIl1WXu5wnO
yXG47GEkH6wYTifJv48Ww7evZLnD03TnkZsHuZAl7aIFbDXkwHI6ppFk3RmCmpSJ
R0J3xI+z0BYg7jqsZl7BV0+Jk9BaAVz/GqQ4nJd+Y3TJBCFZFNO1HqHSs75XG2Dk
P6jl1iHBkp8jP65OD62PThmBNb9G8IFImGFhlJHDNKscy7CBpnit0+Ie010eKCJs
+VOzMXV7TaTlgt54TdCiHeJ9RCV1YZNkMoWHI6SKVZtneq4+s8DB5uoJOardUoO/
G2UpWBPJ6d1VI070hZaw/kgZBtwUPmy9RSuiyGYKUT98HMm15EzsDSOYYNxRML1w
9731O+rc7Gx97haAtDA0spwQ1MCW1Mir8INTsZd1S/lIyyJS9f+yK3G20A9D4k4q
R39v4O4TfxeVD6i8TkWftQFkWBTyWU+LNRn2ck/fu4h2TP5JAP23OmEBMac+f0g2
n4byyUXq1cKkqNBe/7YXe2QTp9pNVWeRYCuuKX20KdJMTVB5/KPw6e/pIEuzaiVN
efe3eKA8aQrSgDyOGDlmcHCZB8v1P03BPwP60fCXgznuoU6uJu7ZNpykBCRoekja
4m3nclH8PNo1p0EDpDXCOHchrzT3louQPBGVv1+iXKd6bV+S/5SuceWbW7jWhvbV
2on2jg/GPiAVW+3WCP+v/KlSDMGnNXNXzq06zKwl1T5g207IS+3PTk9qdGUJD1iP
KQcDgvBWJKWoeIyKyq7F9luEL96lLzEd/qJZDLckX/cWkb1O75pridLCctL6bwXc
gkisVtgNkoWapeiYgfGg3rH0jQ/PCOoLNNP7CE1j4Hr2aQBrb5Hz8/J6AUJQqWOZ
RhPwQ+jMoE1NHfv7Co1aHKc+6bVIYeknOvdCBDwIBPFjY9hBEYjb6g7fXA78J5VE
s4eXYBDKqSM1hnJR9iJ1lVRNmBDr/4myopuZisJ1BfGkw46MmZyOEhWVLqA75aml
KvSWGwyjbcO8iHUbD2pH2hAdfLQuQF4MWhllssr+GAfCD7/2YMFOuuxRXFZ6hNmI
4VVH40v4SpgYkZOlZx7tKpfKW4AqI2jkW0vQMv07f17ZV2Yj3bGanVDyhzukrsyJ
BoHIkQl6uNp6bNkajj2BHkyJ0J2V/2RLR+oT/x3tCeJ+SmUCfjTGCCRM54I22UOh
hzQ351h8J3MBIJ5GtmGYtKHCQPzJjsKp301wgkcRrTq4fhleBMzr2z9q+dLFxqS8
YmKXWZkGX5jS+4hcKiWDxl5L9h1xzynXejCmArmBvylolSpI815Jm9XmFuTnNAgR
B6lttG0eyQm1B9lv5fK2h7AjUcFgSf1CDCkVKYOlV5SLNZcn/u7DSK/2h0r6dB36
tV2L01mGk7SSD8FXFcfc0mf1DiaATb0qlPKBeBjzFoFmFVFBF5xOhhcA9axkwICM
l+NuEfloehAd9rZRtqS+9x8OQvxMUHDlVaFCrln+C1BuT6d2p/7cHtBwfrIPAgc0
HWBU592qKZdv0FRIkUECJKPaXvncIEr0XmZ0HBlciJuU+tIKye8NzeKmFyVj1k64
Fz4/HhJJARXmnckRxjLYq79gZpjtM5aUSP/3fkY6qzYWa6JEE3ookQkT+rXdGQ/N
Qc4hlrBMS40vUvUX0B5iY5Bbt9N0l9J0zNPVers2VxTsCllNIMc4A9hu6OFtKrLr
ASotH2/GnbDH0pFlBk5PZ6ngOkVq3X6z8E6DG5kS/P7wS7EUef7/uEOTPCQH8vQT
Z+8wARHyFeT89gfV+4imlqsn1i5Ji7fldNFb0CahMICNBDj6lO9Hzb7+RWLZ4Yk7
Ma+pn6+/B4rWJUngQj7IxN//i/u1HCXfVGNlC6+UK2qNQ4m2rjOmzd+JOGHsLhDM
OAkIxefeTHhTAEpGzMEHaVedjAagb9LPn8C/E9iKFUxOzU8EYJMA2IUT6bD6uzND
VkRk874IqibxW7xEZaVSwo6toGIcDsiCJ7zG/bAZwdRL897POxpvZk7ggeh421cy
DHGB7IRwZbkRjmtoSwhaOkAQdY7oMioYEIBy4m3oAspttC6m692jqUYQgGsO6Ekw
10VxYt7qCL8MpnkYZGPsKGdL8KzZXTsVwudnJzJyjVwjVolfzW9sSiYOfQC/KDcB
8oV2O2ZYsJX6OWvQybtQkZGNuraDKZvgyrPoPWRb9RsjsQC3JhR6ZFPdJhSfGjt9
tlJUcxVTrnKOPpZRuP5+sxPzQP1EkOYBUETmuB2qQY6ldX9eZP7bpYFGYNX6G5KP
Nm41pW1Q6BsYhEqk1nrtU7NC97dfxjcF0sfOjamkCUnZty3JEl8q2Cp76Fc/bSLe
`pragma protect end_protected
