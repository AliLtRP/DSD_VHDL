// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Syj8vyrD44QzcylTmhMoOP5cNPK6YHAWGNVBXK9NNc/FxoNRpLYG2HLiliscX1bY
y9CXb7qt77JkovnzddRU943AmX8kH1+kACo50QPgQH18HyOAJDVOudqtVtZrCh7t
lvP28jFUEbjvYX4rP3XsLsXbL3eCNnGwz3JW9a7Tcxo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7648)
f+xdSfqzZOAY2X3lXAw38d49QG+gRr/5qrlUfRL7PeB1FCKCa9+McOG3Zzl2q72P
4AoNnbgQb/YLb5UCf5K6BlkdfJsEdVkWHSSycDT09J51Sb6gJmLcARiPjfI1kiLv
YCkULK+/vqobMmWGnA85T6QDemyuVei7l1p+QxWvk1xWGopMcJT2+uKRYK+FGHJ9
aa60H76tGqUsX1ytHWGFYl1z4bGjZN8ZC4HdgILpXkvuUkvKoVIxG22N/yNvBemW
E8OPmCK9Rq/FpfjZ/jpggqQ1mvznK9Dj0lWmrrjM2zAvQT19vpvxYjs6UvzA4lar
GPMBA2tP0He5c9Hbz/RM7FgwADw/upoEBXeEXNMGPV9qnkG1fX3PSVJDuFiia4N/
WMeogcBQ5fG/BqixC/4sgiume10k0ldV8wMeMH7ydFBFo8iXUgPtgxyIgZrbP/Sp
u17lEg+L5yDtd/yEfffsfFePVxIgBz1SwhuWo2eb/+jfy3gP1CPEnMInAqfs7oZd
V+eTl7vC/ZPy75XR58UriY8Y0RNANj7booeiEnWH1dKJzkqOZ6oP1mk7eGwEAdEk
FdA6WqTx6JKjNwmzIvHeWXdBgqnRxOoG/toISDxXbBeMsBMSHTaNMSxZ6jvabsEW
ZI6MGvnQffo1dZGEdEjqezGnz2psnVt1U2Tvfh5b6Kt3MsZZO9KmVmLCWKlyvf98
o8mb7PTYT9lEErif7TMRiD2sXiMHzGrQGY6zyjo8Xidr7NpM9vvCu47Kk9ccSnGG
bYOQlE85Yvf6sd78PzCMMa00moFzI9pIma1ZeTUDUndDTMmMg2gVyMrNkavMNVXD
ejphpUumpm88HafdDRrw+nA3l1a6Euh5uUgunUjQrEmzz2heK+CJl90jpnNhwldg
JYPM8iuyewXKMThSOeMdNY7zXwh2WXK3GuTD1dLDUZ17/zE92LKKzd7m8xnApsXk
3zdG+XjYsI53CBlNr86pN3Hmc7wET87Zdx6G7jYHpqlFXLbA6MCkLzlWHTHtkamy
ofMx9teGAX7Fn+yvkYS/Mbgtks6HGAPzTTHkiP//S/OQhPa23eOpzEe74ujiAp4Y
hopw9n0d1isMwkd1X0wgGF9iPK0Ae76E7o0MobUrMc2hXKQxCBuO1D22XBounPIc
VUP7F/ApkmeH56LFKnWt5a5lSbrrkf2hWciismxW6gObjjoWUCHxkBTSTIsI+1w3
1zfcwT8hniiCIx5M2ZyCpBMzevawILWhFAy/ZltKel/rz/NF5X5ce/zn6gNP4euf
Y1yRj20JMj9HANz+mR16kDiaObYK8dCAT+7ek+Kuilmkh8QBfUT5ZuHZb4Q7ozMo
y8ezhcV/S7iR9l/5MLmZ20cYkW3P5t9l9Q5xnRvDwz+xjgTJ6FD2kfKK7BA5D/cr
O6NNhhEJg6MFaPaF9rymWGyvMQSyNvS+kliptHS06UP2AD9ahxtkz6h4YEyg1r6s
bsXkrEI57H9vfXZ4+MVTgZFSN27unRvMj7Xvvb2cv4GVmQLT/4DoFYVYAYULyoMi
UB01t30WIIl3ak0HEAS9Zud/5OzCY8iWjlf3qCUNKlKKyfs8jBcARau901QWPlUp
WiEufPBJZ/faDCKTd3iUwLz8k1Zl4elkcn6JHZ/d481JwWC4d2j2SyUIq/TIRKiN
efCbuqelC1BXnQy8O7ss9BkGryiUrhBqvRnFir8+VNydzJ1ZsFBH1sq3CCbo8a0i
nZ6cDJUT4javYhcVFc2FBwmRA0aGqT2PjL9B702224wt8NNGvgdCU/r0t4bz6cXU
qldkbwmgw6rWUgJco7N5SA7dlp5Yn9R9JaLFJGkG/QkAimeMnDNTooXSM0yvri9m
CIWdDBhYB2Mmbfkzu3bY0mJc4Z1eakL5yUZLwWraCLDXuRr93w+I0VM8PqoOOAO4
0xjMPAkl2c3/oFVHj6iwkJCuQu++i8ki9MX3KbuzxF9Q1apVmnCuH81amGInFs8N
TbHByiDqJydBMcALL9mRMetvOI7c+KVx1cfOoASKx1hoOuXnAxZP47Qta6jQDBhg
UxeY7eydfd8OqNnypCjpFpCGqE6ZXKeN0KLLkHcm4lRLi17IxgxGJ0zBRtHR4j0G
kst3onxQ1RdgI+yMlMRfXWVZPe/vSUc3fkCTpF0CuZtn62Jtx2IesHFkJMPTGaYG
nyt6Y8C/ENk1Zv1jyYWYwDug1YnYJ4NzluV9oswx9qejVGyQwGPKM9XabAtoixfn
wkRu+QVk45LuqscS9thYC9DfwRxNyxAM6N9yle+nIMU8xI7BUgXGCsyDk5qebDr9
VhZvp9IrKsYlt1xqT+2WwckzjOxRh9BHn6BFsXYe8WUFYRZxIMpSIkVNXEPcxRnc
j0Nxle7H3ZCAxNW8D6TsoBkouQSvHOp7w6BR95yRcWqGbe++RV2MQ7hSre/OKsrQ
9P7QqEoLXG4GpEegN4DGeaDNQ1qK+6dv4h0EjmqP1XKXOxt0FM/Ns7I++ZNSlphH
/unlOGDseDKd4AQeICarV4Af0Kz0GUrJpnoGmMNRaLaCRz8akjAksJJEsD1mc7FE
ADkhbwUtNYE7ENluBd9/CeGgQOmLbETRt5CHfojLatt1L/jymhGTm8zGbVuKvRyv
rtWqXhDITuYKvM2EhwyR5bsEiJiG1Z78/Yl7k5gmndH5QHLFeMIJENESZ9bEfYp1
O3xsJYbe8zWnlHxupR8kYz0W1l7h0Z/632nev0VKL+3TFymDfn71W/AN9dDdmHJB
Igoq9qv2x7rHznMi8BJlMxQRloeEfOdHKG0zBXMwzqQOBhCfKZVfboGSD9B+X5Ya
zm1zWOpUMDR0LgQTTO93mqDbEXrgfVdlRbhHEmM5uH3ddzF5KjHaE9iZco+jlIcE
J3thUyquw/ebSTcSTe6Bh3jBqoq9Q418uyRkLQFa/5wlXBKqTY0zSxpJ7RdXwlDb
w4z2SqhUXZGCqfjbD2zpkDjUC9v8pK753VMiIpf378KN3D7EssMcoUzBMpYz0hIU
PAX5sq+x2iuiyuCbfxQOoUT225Xpr0iNmU6q3WLRhODcKCMe+GIXFisIQTyTg49d
AfS0YhIx7bsehEn87ZFq8/LOVXyT8XbMCJ2qZ8BiI4Y7CauMBPpQrUAqpTRMArP8
s9vGraKWs1fiZRgS/o6coX3PFpcb5QOwhi24ALf23tH0pk3eeOCoUpErasJodOoY
L4UQw++8meQh74DFIwZxUPDnTKXnMBsAETxXCEkVBqfF1jgUAoSuIAG+uK9TA2jO
Bs6ugWr36buhyQK7g25OzBjVas7IbyhSgPqzTPm5HnoQ/tEAW4S+ww45KX+U8/kA
NUCShsCs4wm+EdCkfia/RYfEEaBhk8Sv/jgwODR8YNDnh4v671KWmsq4rJgq5Hnk
k/eLh3AJBJpqEC1pYXVoTSl5La+nDl8eWsie0b3rN94RIftvd335fpzjTMHAaDMG
GTVewzJiVmrzmcTHUrVZmjCUMjy4q1yTbAeIhrITn0oxpIpfdb9MNigvuVpbd9gP
tAK5ZZuWW6015HPwEt01neD1VgFtD0b8njl0Iy7HbNZ3NuhinExLBWfs1TTgkyuR
UUtZr+FZ2KyrUn8TgdrS955Qqan7OdUfkUqLUtV9QiKCnG+SUrVg30ifuFeY3/ct
rx5ywS5SEgMI+V/1Vu656Opy956rQuV65gWUakd6kBGA1FoQPcgwZ2U8X1QUteQy
o02QiOdHkiCnYN0QUQJd2kEKygiwZ6uoqoRInkOYqwOBY6nDR7HYLma1BhWk+7Ba
AQ9oilCgKOAw/adDSwqel2Wm7oHvhoWzxctcykBHemvNJ4zKZFWEC89w3C9HyK2p
suxGhhwc2FGMMpd47slnyA8tsdR0hAgdSu6wV/jj88gud+ThjTA7avZBRbFDneYK
LHhmEK8/Im49jnABAK7d3DpmZahIJmUA1dHD+8TEZJrQ6HQm9CWfhGkIwZZZroVt
JkRsYjNvjesUpzTyj0FYIvslZ+kNvGDqxuqcReBuRmhbkgAfxf8y/YK/ZZpfG7Vo
dcuX6lmNl5IFVddgw2hjN32iCUk2wtNaspvBS/gf03Iu+M7kbYRWhv5YozOZskgz
P4t9tIxNN/dl46RKPmKIEZaBdG0Vv3XSabvZm+XPxwk/I1XffYVZo+GxPF0TgOEX
SxQOCvUhVRIu0J6xfjkYLpMIdjp9vDWt8KCVbXvRU68U3WP93nzAwPTDb3IJ5sYf
GwRRJwapOwHIcUqvfuIe6BMpoxG+2Di5gj+3+nXuahtby06sZKRf1LvcQn5nvCbc
PD7KYPUiq7HUUj9Fz7kuFUQbVOqgCQW9PUMiON/chM9zWgxUdNk5Rhuk382+M5PA
GX1C5y8sL6+oNyCpP815sCIFPNGTGUIBZquPuC0jM91uQErStl2L3auDqkyFT9aj
t+ByJphMQ/eBDO3KCXKcfcLzzXQl/pIReHztgkRBpGur5GsowLfmAVB8danV1Jw8
MBsV5a214VGQ1OO8FsrSIGG9hZcv+zsUT0DAy9bu5wYodU4CXRnl3CnAhbC99qqN
rG2ZToB0VC/0TVJP1mOGTaJ3C7AOFfLkBlMw7vzo4KObHxJbg+PWQjFcrhAEIG8r
ejluclGaBvhkSAauA5ejGS5hq7ymrplPw4u2gtkYmHJ5uP2Pw2obunLZj8xXjNFm
YI8QchcyoAyCU4KC+AOo+Zi/J6vUjSiF1ph78SauUKRJvt3yP2rY+WlUyfrrNTbP
UxkR3Mtw+AN8Gcf3nY70ycjYCecVH7hGlHOgqCh9B2xpk18F80HGWRYQ+FnMGQfo
4906akj2NijRlWPrHahJJnnywJEumgERMsHRkoOGw0sHMzG4DddUFY1CxKV9/ozd
3JgXxhMdtv0ux6LOq1NBsoZSzwsMADTOUTseXaPA73AS8qKG3cZg/7WXV288Ljng
t+t74LEhdEaSMSSCSZInlIhXHOLc1Pl4uMsvXPXA4MPvtgCBLffSxFKwXdh9wRVC
DfDNMfikfIilBA9670umdv+RYJat1gwNCpVt1ehC1UbuAClAQibDNkIBQ/edSE/M
99+TmyKUv8aJti6COjNHxRKoiwlyTGg/YrP6qFFs+WbbruEoHGyzviGNQ8y6RHmv
6Q+wuhjLZGkadRBf3HTE18FXzLfElTtTnksh/reRfgO/W1f3i/iYzbydvPp9EvHV
uJidoqxkrxyj7grsFcXaCRqCWqYhGCGF7BMQFDoDvV5KizcLE0CXTKLSLpNp/BVp
6oWdY2cnaWBHrbelaiUy8vYFUKetY1kvuDgx8fVYxpaN2k+40N+ntZC1J479bY9s
2pmp7EFxWGvdRM8XssgEAbRLBGFlm1JuuXUndJD0+1ZUBAPoFBDcYZ4/FkcPUDGJ
lfZig4iK9shH9/Nvx2R0a9Q/gkm1q/vxvKzXI/XRTuiq24+psH3DOEgjESBTEtQm
vQk6kiFVeCnhJgh0DQARS50DhSLgqRsg/+koyF/H3tnkTUhwMZonlu5NpBT7GqJ0
Z8G0YkhFuN+DRvxSKXuUU1H7Ch1EJxYz5vZqIio5lZUnM0UPbHibSL484vZrcTnw
cN8T/gx7Jr9dtYZUSq3pzaulUHIbVOeCHTax/22iX/5hJtFYa6ut5RHC17kN9104
y9GLPCl0sH+lRnHzyH0sbBrujzUncCWX8VDjU0gy/o3b1aAV0USBYoUBW/QZUBl6
ZuMNuQOAELUN41E1Ywvk+fOCJu1m8LkEh70ML33NLHeMJnSrqILy0tTqDSKMamsg
QF6lxzue23WgaGYTkOcspjQA15WQxrNH6IWj3n6X26FXrMGe3/LC1SomOHUclRr5
he8CqY45/lZCg2jXPUWTjMwUjmEmFlt4mVIGDcyD3p/IO/K5qlKysvwzLTV7Es/v
2ZHoxA0w321z6Xm+07jn12UQfBhJSsvAD/yVJ2o5BO5gP99Eh2whORK7hFomjPh1
Tuihq4HY46CsmpNIr9vfZ1JGMCo3Iu+hJxi5aFmo7Rku3BehKHcJ6XigewoPw5AS
9ObinNgKQlJNjhqkkMwMSTp9BAOclpmFpxMjUExUjcIye07bmmVJ5B8Qhsc5HzN9
ipSrcaBvh5VAVz2cFP7Zv5fHamk34O+5HS75nyevJ3fwMqcqLdKBsVeRtgy2rFDD
J9cUDESKauejDCpiXQR+8gGUqQmiCGzcjhTyS1Soz8CK4qJii3qSeNcv1deItimX
hnG+lZ6mMfZFjYY+1fg49iKVVoON7dkGLBaOdrj4Aighx0YNVydr2tZ8AThzmjm3
n38VpiFRkYP5uoq5Oi8aZAwZOkvk8Cda3J4k58qBeUd4eHcCmXhUB6xz4mYnSa+g
H3dnJEIt5ZWwf9NKJWc5qm4HPO8B5TLLjgBeCjxAnvghqTZobSSh43JleXtC16ZG
5NQOrvPpa2e7oUDWNzbpXwGQLDm2LZau/9hxIX9QOcHDJC5F0E3MnhGf69idkEYE
D6Awg+PDQvVmNCJAZKcMZBtu+nGMjWUBiTfj4+syvvn0J56qywVSdZ93lPPIWWfr
t6RE3EfTbj6FkM7IRph7C9YDKd9HpxcvTgLcLpOZ+5VdbWhh3xvhbpiyJ9i8/sZg
utJO9si4uiLB77TMorY4LvfEs6TpAh9vA975oSrNZdgJCJxkyXpJRYAiTEm1ENeL
8tDIChQc/H7NgrbdebrtOUHVAyJql9BjLiNNOwhpNZrQfOVxYSnY/laq4fUQMwbV
sUvmDMvjzzzaEJjvsphCij4DjGkRVyCHMMeZ4hwvGuNHpRivdlNsFabPuXd8zbNV
DcrqQveqaR70MxoRFhZHEqeemyCVM+CLdAWL5FAWkzzFyPrZwpFUbfcLA7GI/ShK
xx1o/ZsKdJGz9Po3uhh28NX02gJcsM4xLByCLM4sqCEpuzLqNJ7b74kEIQMPari2
MY42bnxdmdBJs5XrKtLOP9s85CWzEQ8n7GNGPS5F0JK4FGChIVAAyietVQMHHC16
M5bCI96bxoRsNL74R8f8n0BY9RZINjgsub7W9qOGe9wsON60HrLlBKIgYnMsJ2y+
x2TJ6DPeIx6zfIPLKObrPxK9gkfgdj5ra63kB7qzCn2KsXZapJTaOHXNoYRDggTc
r8mRyXLuzbp7qbgAVQ1n5U6Kx98WaJ1bsblGK/9M2g4Sq7bg+ta5zj87W3+w8n/X
t8Z5690uhsWd3jlVlY1GNPTcbFRyxJeCX2w4r2nIJnpvhahzC8D/Nko+9f8M89Jd
nXWUrhyEpxhrBNvqgNzlmuBUTp0InUqLrhXnGjzZxjBq9sIMiGT8KSHhswYqt1dC
584nCGUWp2Rbb8EvhyIP5Pxr9WNm5kQKIUmNjQB5k2skDBYetpgXk4gn7HYWFq7I
SnmcrVMp7gzzt0WeLodQ0GyHY2D+b+OiKa+G6MkZQDOHWFH6lewvHo0MZKB9wGQY
8FbV+3sauCULTWPG9K+rFzG5APAchW2ueTJFi/Luq3JBVYB8Oz/M8B5/TxUPZ+Kl
VWASeqmywPLmv+BQw82NzUrefmaRSGxceblFckHdnBPvmSfi2e9dY4GCG/wnJsWp
OH+6yfhzAQxrfzG7G3Li/HU3l/RIyt+Qy1a4i5Be2sqIaBCtltt1c/iCE7eNb26h
pRbsXlb9zC7CcRj2S7C4qKiuQCpU7uwKbse2c0vpIMMBO00XFXdTWeuAIc9CTRvX
Qk6l7OQUnT6p7APxOL0UqD1tlRdftEL6+tfyAFIKxVHvAGCBW5ro6wtZ4wCeziDN
G7vSg0DPG1kCHqs1C2pRERvsVS+HwXW7XzdhuHbDmzPAJs895D74z8oL/EkmQvlz
TE3eLcSr3ihSo01x4yn4gXxZ0RYi9lo/YvJNjDT2awH75Vux/+wkzKTnyM8HzhrB
OCDTX2gjbRous7Sxu4elh/xFmOxMJXd9gAVlD8FZgsN+e4Qnolw6rLg4upUu+c4q
T2YavJBjKOtA3UWG7j1Q+qd6OdKXNiVN5BhCn2JSG/JSIUVkearQitF6yJEDIMTU
1pYnBmIdeqKljT8V9J5o6jVxnNV7V0McoGSO2kcuKMTVJ65MYf+J/cgapBPlqnbV
6ozeoCsukJpewhAWc/ul47jF5ARXgHVaxK3m+3Ltm5mopCC5z2TjynA0UawjWOb/
bpTSpfljo21c2Nit/By4nVM/hC+DGf8G029rxLZnlDh2ZiKfENBBjtPH9OjrN1xc
ZdOzI0q+1ki6Dv4KXnws0JPo0W9FlCcq6Lc0agYZeoDGg9zZ+8zEvdi0bJt4pQ65
ASNDO4MnnKRl5+OHiTct6ici1N1P8qPd5m3S1ddCEiMEgRqI3jToHTpinbknKF8e
LybZKPNJUPdb/mz6baVOaK4trtmL456IA8Xm0fpseT9v2vZJgoATSN/6iMzDPf9v
7lZFV/uZJMQYarqlok9DLWliuZeu/Rrz9t/TayWkMTXRy92etX2LflgWByilbPQo
nsaqvWTe8S5lM3SQXkWQPiBuc3Xgcu5AuU1YG/6Ql8lt6H3saQCm4PApbvwnTsP5
sMms+mm32DcJXZjn/7Svk6Qu3+MA5quGr/fMN7CeYKOyaSrvA9/uszXPiPPEoI7B
O0tPjO9arHrDFDnNMxIbCDSWe0Z31zFXBuGGc0lMLGL9C+uT6tQNckwPwRCdz+LV
eGutDLDpeRfY/vKolopPsTWQSiClEpUFXYPpEp9HC+tiJrIxk/IXEUqSx7yKLMAJ
zogWN/VTWnUpseap66dLk5byZ6JWXHT2+9QGeo0pW8guOCoDwNrpJDu4yaewy/eF
v213WHXtHCykkfyOZ1i8vHqID0wn7MUZ/vUi3Z6s4sn3zaYz8Zh2LMS8qx5SGzAB
g9A1gmEFeDu4ai/x6djkRn+Lzpp4Bs0Be4XsH/P1CBovQeotQMOGA8nYXYOlXNdH
utu5xvZfvfWxwPX9hkAn+j3hM+lQ6PEtZ/Hih/lUiymzlahBK/3kZJ+XEGefolz5
YRVL+KpbeaI9mB13Km/I97Pw+Brvz11KcPuH1uuIfOA3Y/5r8MwIWzpwl3ifVhLA
ikYCYO3dbPYBM5fa6YO45kBRpBGizTQ4/J0S1BQ+U7F1XIC20Rn4Tdz8IbilvnM6
RSuxW2ItfZbt6cthZyZF+V2RjDWkDAzth6lpRjQCTUXCyf9toTAdICdu4/HWsP3m
3uzb+KerGxRQbQ9ZYDrvqEj9RkWTPVID5WAEA9XgejQcCXu45hR9vhZqTBOqlDZi
Oy4clRm+2C3K1DBoO0o7460JnYTnKFyGYjnLkJ9i5A6oOAziX4Xne/aLsm04rkFp
FSxX5kRM4QP6bH78y2IagvFW887l8geXSAM/tKaAi1jgwrZA2Mm2x577noCoLTlY
ql1dM64Qm9w06baQ+wYO6GML/lxubcr2ctz3kgS8db495LWWVD7Jqg54gwP3ArU2
38LuxJuolSHpqmLSTgoCbD9++pKaxbpnd1hdectmmzGliXmrKZzNEUwxh6jkMISC
K9KIDT7asHJSTQfNPcW5+iXMBdqCu/mSc+s0+SEiyZE06qbx5zDOxNr811MtUzpZ
F5xuN1k9FaMqLze2OyMZ9TUycvzt9y+PvwJH5XFbQ1kkF2NvxcdG0nH0nZHMynOV
KfaKlDzaB4FtCDT4AXbfnVNB8v3Tx0XMk/D72mMEroj/W79OP8fqLEAI+UxkhizC
cxSy18FAT42FVRBMBxhJitJXSF5Gi6D865Ge9qav7e7eejk5LzfI4mPo+UpGV3wG
Re8/diSZ9FOSv9tIWowYSks5W7jFM7K9hHCUzuqnheYx/P6nZ/OMztQGrXJxt/AH
6dsIsZuza2tMmQ2oq48eHwOiiN9O7ACK7LjdHMVGEJPqcJ0iT9sgXgVKy9S0t7by
Y/dWD2T4VcZyoBPuDoqzik9cIaRNllTuJvdnrmuK+wJ8fmUlKQbDcWaHkETltRzC
6gxLCkjhTPr126Bj/2R/P88wUU88uxZ++aEdrxonBwYc8xkq0DhpvtZ9CAtx8K4g
Z49A08qUPCMpVcdrCkk5wTESI2z9x/5o1u6QD7KKpw939QB0FUFDotlqmwzRacnW
diLg/o4Its3GDJZVffeCNnQ0cVzdRhmJj013+7OAG0uI8cT1QOG+Nbhm1o9lp5wT
56p8puYrOKcuwb1lwwvSqvrE+CCV22nE3ZMxMR5ECUiVrah5ZrZ0oOysXsjCx0F1
5MEQ1uiu5I5CZEoMbXaTlA==
`pragma protect end_protected
