// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:31 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BRYzoiLCDtsogtOopPmlsNXWNS/+GzUU0Xk9C4/mKrmkfM8Y4H4/oE3DUa1u38Vi
mmAkh0A/TIys8X27nrpOHIagdYo1/xYhbWPAZWAJSkD4yseG2wN2gouClzVKxDeh
w93lq3l9ABGcDBPy2USeOXExUQYp+IkZQOEkuVrBSBQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19376)
hPg78N+CFLiF+JltEul6SH5gLsdKnMrMC02P+SzoOsHAMaRSK9EA8G4sfhR2qUlj
koq4ogMJhW1mU87C1GM9NBLP4HQEVmORxz1O9blHEah6mC9zNkjgQ7TDKJvVG28Y
da3w1eEBkXQ6AeS+suO9rWkszJD8uKMq2EmMCtxPtfQbo/qUciSS6iz+sKMyzUxu
Lexd3zQ7py24d1+DGIdFVtVuHJhHdYbdsn1hClKsMmpD/Ks7yQFjiuexeIzDbA2b
2gGfqoVsoDGpmcWRQcMPxavmFHc+3pSa2FCsvCg85IaEAJ4oyz0VntsAXfRT1Uj3
mwgFcLpH7ib9uPfPPvTqTHwV/BlvMJJmMzoiquC5xmFvUqWSmv3O16GCcmGfZ0cv
lI3ZtZzin86x/dECnQNeusfpIvpDKbOhnZNG03OIfEfQwCkOkqBGW55Px0i3ywqq
SBlz2kzIpdmjyqVLGOuNHuXHBPX9knQeJxXtnPY2pcpoglEmNL2/UC6xS6SEy7j4
WZDBpBaHxSLZbYajD5B3QIXdJLRsAzh0ctsEqPe2f1FpzDK3SeaPPh+Iw7j3wEww
9CxD22ThY+q/s7a6hrk0ZNNvvtrJXQlDz3vzOooH2qjPOnj2Zfx18zONEIM62EKO
Zgjjw+qU5tAPF8/r3+GTMhc7HH7JMs3XVKK+cADj6INfmqKLVjwZxaWYHCpYrDT2
haR/GTLvI6ML/fiUUllciejE69vpKef7sO6OcmpDH5CEr85pgK+8WmvjaXpuGshP
q0D/7dj6od2ArOC+0h6EuRIeNtOoFi58gs3qJEJQlrbQ+OEhdsfC34fwDMyiEaJ4
XwtvZWK54COe/snKoYwqBgmiCH2ZBJN38v1haZmEUJTjnD9g8ZOJ48q4sld9UkrU
jCU5Os9ZQY70K6yPLcP+qdIxbQCq9GpIKilGhA91YBdtJQdwewLZYIOApHCKavph
MzFxtDAQIsq/jB8Rn1Sw6Cjg+cAklnqYM3/Te1xs3DNBJQ0m4ZLXmqduySp33AM2
GxxFpJFyMxkbBrVFPT7yX8B24U5Wegk4TRJU6dSD9mGlage09FSWo00PkfTcVY3q
sTM5MjR7cxm+CtqSezrA9jR8qC8CigSMzMMZFavXcvDsJItEkULXvWi6X9KX1o19
2J4C+Ok4OfyqJny3Y4AUScLFYFcFKDeGAsV0CTUgq8TQWgfGZvO7X0BdFa3qI9gJ
AHijXBwH60hXjOGmGLLawXaE6kQ0s84lqX+fvXph/ADxPkMb59LELIc0YRMgywmZ
I4H2O+Vm+grJ8kO1C0izVYBptoR/sT8vbPtyvhHlnEdKsJ2uHMiCrz3O+h/Y71Vo
yK20po+7IWAMpudc0TudF71rF5titOXRlzjOvxObY/8FNrZgfdYWku84CVtAXnZ7
+ue2Nu6e/4aMiQigdB6rlecX7vVU7aYwmpBkeGAHVjNktxYA8QV2GNK4/1O2qln3
VDvST01mHPiTJ44UU1+aTYLylr1/Cd8l1K05EzS0NC/1JzAjWGOqrTWx/amG+DWE
Q9wlXyNsAbwrkfW2wDuE71mOrym7v6e1aWsdCpIaSz78Gk4cM3aGBSERNGUlHY1Y
c+22Hsej5LeEd8cLqGWiJzmXuFFeAE3OEiEcl029Gee4aWqOmCAikjont+4Tt8tJ
Gr4OS/HrSuuDsWVGf3dBqUVoGH7OZegrr3vOcu61Etigx3AyRnEOguQxA+po0eTx
diiro6TwR+QqEI9lS701lBe30iDETbdJepmo/04nE6uNExWinv7SK29T1s5xv1lY
gM/eJmJMg9MbOYTkmIFvf29w8rTUMhRiT7LQRvPUYfMyqSIkJVzir0wFSfFRlBMX
7XC6qYPGZhXf1yYik2g5tNGKrbWmjRvCkJ/GiLBD5eQZ8rxxmXhhrmyKzXje5Eyq
J/Gl1P/b9M2M700wEIoTw5A9RQa5t2+UzTYtgZxNgFhpCXBm7F4HyJe1ZRWaxfxa
1CBWoAB/Sab6t55bIIGekfp4499CkU7kx/gNPwFvuI7eedv5i9pXt0CsvACTmsaQ
+zM31m8DZSNNHjbP/+4lPSZE+e+/003jqDRWm/73bGXZ8Uu8cKxgViDgvh8c8Pz6
1rdRUwIfgtijz6yoO2WouJfeIxE+ViWXEkAe4AJRK9kwQcBsyE1JXurKyf0m6T5/
m4VueZ5lOrv6CQDsQPEfgF6t40+R43ztSS62S0VKwHmJX22X+/39NHTr5LdDfVEn
bEip6RM/vXth4w6oRg3vgSEw2PYI1wnqzWUqQ88DQjQuOGkZG8jwKBxmqab7jw9L
9vT3po4FHHtyuebGtdoCg8VPPThv7mGqVdp2risn9ajKnarVzHIaWYn+dH/nk8Au
0MUKNLuKz0hF42ZFTMHCMXqhT8Bmjll7QPR8mvLsrH6ZqBqtIDZtuRsrP/ZACRIS
o2efsPtViBvPtksNtwmKr7BYIVL+MVfE1L3Z4hnoFUFs68ng4+IJIvs7WcUmNqIj
3upv9RWdmJ5d5iWXznoJyvV3Ds7vGVUl/JITnr+1pkcGjp5YLiGEYgKPwQMM6m0g
vMQY5wAsCDllriWnT1eancMAuj592tdo0qdIgqO/ipWWRWKt4WjJ0pYfrCih+H9f
TvcNdPF/xVIvdfGrl8a+TzRu7eridsgHi/vpWgVehmaTsdb20XAq5DqjZio2QPB5
dZ/HzexhZyjjp5/aarEmcvaI56Z0x7qeYi6v2hOl9AQ9RhlrHbSRVxsyNXph9U/6
h55dDxvpd5IcI2UIvPvweEMo/Ryjo5IdStda0m9bVhfCF2as6kue4E+/d1qn8PFl
619QKjm8T21h5rliLuJ4vVCQWeokGnjkpR83MPykt/ryNuU9xG8bETYWslb4Vb7G
WKXiRFDtzGC9W0cn5aQQmZXtYQDlHpRBco3q+uA952qOSGcusS34WAI8j8gO1N+M
F/WLkG2Psz0qpAmGL4njVTdmraBOuHfVS7jIX6Zx/hVqorlmX0PWAxuBeKjVHtPK
t+f+gPr/xD8sKibz5XG4e+v8IBgT4mICv1BDavqi8JWTtOUPQgxQ7QLGCnxZho3q
WOmJFbBP6ZSyVnUpQxVXF05asd6UEIk8+nOD06PqptULRx9VgWhRNRn22f6uD7aA
p+61Sl259+GFISaSvtVnfEhe0V2WGSapzTV88pvrkmtzMz85wvEZtU3uGCJa0Joo
LxVVU79QpH0o/lOmHXalN2WMcl47FP7fhBa9UzskWyMHY93HGfCiz8XaHueHxwQf
Y1VHL0EMeS13ui0tM+pp6UGuBlAAwT/ZLhjWbnCDMFN72/RSYRfsdAc/NpEQkcYR
uFXm7sJbcIPrICwlXr3EGfQLVmvZ2R6axKn3Qaq1JPcAOC5aBc1or1EjNgEpda+1
tCBUVZhRQEChEpok2vkLfidOa9iLCaUyYRFrBjJodOMqPB0KOE6ScbPVGiPqkQNs
JUkvF5jWhLkgbsdpdKmc7qVujAXoDsE9m3ajtlfq/chYMnDPRdlxr5cUROqxViuB
willaXa0SPu3W9M94I5E0UoFNDO73B7vpHalvjFynVw40U9W4xHMiW8bQIGSe8Er
BMm9PR2U0Zptm0MPKv4DDX354b8vQIiO01n/loK1sjcwlpG9b6EOweYgTS8MCzqY
feNqP39Pzt7s9DVAhpnkbnWpzzR2ExFqTPhvGFmxby4OFWqVsMk12fj+ayJwStGh
siyLz11Az2zBMFNSb1PRgwSlV4vDGRdEcLhRcv2Pak3l6Vnt9LcVELXzFqzg3prK
dovJK6zhbW5kkzQqtURM6Q/w4S6VbCeG1XPQC5KNWKJXjnlJYRsPruC05AqIb9fD
WDzgisIV43xTS8hNEuhuw3VDv10MaO9jLhSLhDV8rrTzXigjYkMuFTeI8oLuvtkb
H6Koie02F9xeWSMQTfdd67q1o/6+cJs8aqiELzeU5F/Vmzswvfv7N+t895GhlmEh
ra6eMJctHV06dR6V/04SK0ECEa5hKNnRlEJ9Y9IqqJEMR9x8DsvJ6hRXZ5cY0JSZ
TkJ3vOaZcs1Y3v3DwdYp2m7WnzDjxVOR3aYYIsq6g10j2d4pRaeQ/GQy1laiGbxh
3YWufv4unDGaJs0aQnyMd6KQ22o68XDCp7huu4zcn5n5dMA+U5ZPdPG58UNIOcjB
ad2xUyQvxMyCowpyThZuebzQqHXu4TPue9lltc9G4SONkHDZ1eVooDKHCC/II1Sc
UDzmwyAEqVgdBUdZLD0B6NCj1Q6hS+KjfH1Fgmaje/hwvL290lT8mksxQaZivq/w
eWCNZ9nwZsvDx+7eiXEoBAR9bnYsHOKnn6S5fyDgqiQfcxTk3UJmpHuOZA7bOLjZ
0dY6nm7FOefZZ4tCKYVi/bspOkL764LfgNzW779PBzWqVN4IcPepRO7Xth4F0a5O
vTtOMoPU4n1kzfxSzAIb+x8f5xqS4HHucCBkEsDwR5HAkDyXPKlTdJVOmPAp92cA
VX0Lb5JTUk8yx2xdscveYmc3tGdDOyaTwoDyHn14ZA4FDAHeAp80PmzEnsmoDmK2
ItYIwEaokUUYr8alKABhfQORZMVIezhoDcADQecSKz/Kb8jb9CD+C5z4HTsBaJMl
BxgvVH+u6dQtodDGvdj+9sMFhCsOy3bGLwFOOWsUB/w14A11B5J+jon+0fs6UNdI
kp5D1T0R5sjPAIvLnNGRMATmSF8jJ0ekev36mlHZVJkU44Z8QvAQj0ITJslTppLa
aTn7li027w4TxFRHMCe0W4Rri4Ahyx5VhWLRh5wTZo82Av6q2VDT1G8R9cxKPsq3
KjPGoX5Q5On8sn/ur05i4rmhDT29N6pHNSFSJ+Oa7bpYNbJrEtDYjMTA44szgh/z
70QVK4bRsOGDVTJHbrXl0dAvcvpVA0Nq+LMjt9pmQrxb+TsibjZ52jE8fbfGn2cr
xLv+8tUmWcZIjmXnXiJPIzM7bHxSB4mBUp0uQEejyIP5Uqjymypy+LY2mBOSmy08
SngMl4pMlyinH1rVDnmS0jdVSDVM0XaI+Xmur3/qii7r8EzWaA9IWVStkUpFCEWr
DfJoMwXS/MXZDQj4vtfUlMMxwE75HcSCjz01oxtehOV9DHYwBRB2tiKdcSBnR6yG
2RHFnEgGxaPDuDclNm7Hj/nT5YLSngXfyOS199hemil3qVuoohXDIQnJI/zILmxF
xlmbdhVsCCwxEaXvEtx2Qoz+uvqE2aMW7OWVmEnRKBkZRckPE2PX1uEXqPNX5myQ
OrqPv37U7iTTgIUI9sZWy6AbEvDQE34a36DsOyJo9kXOUpW2Al8mDBiD/8LBdLye
FEoYW+VBc/DO4a2rcmM20kCunnLUqqBoVir4Uv7lrEqBV3UwTSBGJidJJZodS5Zu
YH9MI1QUUJo3/l3PRh8d9j9D4SBng7eue+MVQzaEahIrw9ThloCgEME1HdLGb5RK
UOBHdo29JII6ia0IMDZ5Wv8dYSAhHa8FHxmmiJ22Nkr9Rq7R28mfrSilVv6UEFhM
0Tr5toCy6RoIccqfFTyL7X5kUp7NwREIAP3f1m9lCXQTEZjL/gn+m0YVOd6ozQJO
P54qsoGyNLLPY4J+t7OfMgTLj48vUj2RqpXu4p+xh0hqkhJTM3VHrX4dk0cMPeJk
g9PYXha5XoWxST2RY8ptpPtvqe55+8agMnq7xh2Jrlf8s58lZJ80PEHfOeKyYEOs
5RZhY9MFcSosbcQASVPQLHCz++dMejurClEfDp9NKxAzD6EDYXLHN23uRtMVQMPO
8siv4tzEoGfGIUmXKSoxJ7AuHgQaCeGG9hmoKoMavc096tDgee050RVB9yCVmpVp
zZE0xH5eNaqY5TLrkYgaah5XquGREEu2TVYSgIgF/DmeOpWdSOJi/hXqzVGqmSmh
FVp9Xvd4t8HfmHWnWyUByQcfrJfi2sRVA27HHLPMQUdDeXncXSAaycZFUONaxu/V
BEfyGw4flDEp3LdXTlgroWpZNskHBBckUtiTimA8XzsHG871n5YE5uC2pQgpxSUI
wT8l7en+CChHD0tcc33oy+Wef5t5qfWVSdAbyM9EZ41ByQbBtDhUZuAOk8kBBhK/
lJB6MHtGupIOCDZ1UiGzpEq49P3oZ9bRUu4P7czDafmogaNmsZLj9DYZ9d57wHmE
FiqFXd4xadM/K6lH8mT3uqx/Pi+YQTw43Gr36cypC+X3mWHZWmHxoIcjVfH2+0gB
E2Udzze3Hm+YdNgs5TM8gb+6jMX1gvybIcIY0h6Arrr7NMLiSoxlBXHQ+a2J2Tyk
0s3VuKprcibOxPMWAqrvJGQ0bZLharg+NBZa/gDgwUqHF2mJ19m+XatVjbdu7RRU
n9Y8ASkdf6Yge4tEC5WeEK+czLfBUYuLid60YApVAdp6/qBwkP//cj6XqziP9fWb
5IdUxsCBJ48nPzUz50SgzM3FNfsIVjwdyL+HgXv61y5ZI4iWDU22Nrw8N11C+H1k
ZOoJ8WQeia1rLot/Y1qIvexQY5Klc9V0apNFBlC5NDe33O8zlCiW8TiBKaNtqsDB
6IzrpFUIs0Wr3xHIBS7XDnXcXDmi6CN3ZcXK0gOYdNgJ3eECD28Uy1jCnx+xEWdh
kyJpqbU/UFbmMQ7BJyPYuwEZMsxEsqVOVkWQEjEKvVztzdtLTqprTtJmbHcWM7T9
kEo29WU+cQKlvFq1RTijANa2VkwSlDEQcYROqg7m3JYmM6UU5l+DyNgRQvouYUBt
qEQS0jagWGMoHVXvZOBnorgikTjPsa28AuAtrhY2gZnVYtTNXsQdzCS4QNb7SBFd
tPcsKvR+S+n/pUQYbmcpaPXbCAJNwkOjr3eNpW11KF/dWsq1v0AJ4OCa1zM1yZPQ
2QecNX8Ja3iOvDAtWJ76GaUM6CXtFBoVlMWyZW6VaEY802urgs+cZ825Boxq6zwW
41WFocXe+nLcMjzEx0mY1aOofcUPhChsU/x6CCNoGgMxAbFdPYzETNWtnWBLAQUu
ky9SAYEK/pjduORXujNBspBHQBA8NNJQW2CGVWe0f+aq+4t44+UXvnEWLgZwWjNc
XZpvhzwdZRxJp1WwIWyGyzRFHVdo7RQsPHmYg63XSM426F0KbZEHY00m73sryGc4
TLlSsjDyhbiKsPaODn5jkiI7WMXVWL57x9rShS7R/CCUmzxIubgb+qpFeMt2Mv7R
5h0nKrYssng32pffSgCl8m8rZ04sR7GDvJrgspIzjTa/uwYshJAxEBrfUf0y4MW8
T/m0GlRwSifwOQNKm77WPfGHHkjPmMdkeONdzqKxcdx05iWuKnodNLf7A0GZi9NM
10ps1qyl0NpEAphkWEIEzjIhXKJBj60FSBNYpvjcuiBNa1qngFDcrBrYzOByhx1Y
/Er6nPp6o07CanDlNygwhxuJQdNZE3EzK4fsQn/XEoEDYyQulOiIlutIG6dNvlZh
ydwVDWDplnQw5xBpCBKkeFaftksgHtzQ/6W+P3AgBPun2acjN4HyrKOUChw2imq4
dzOJ1elblseMCSiy+KyNEhdDym5AT/QkCQofHZ9xmmNKQoUncewUtXXNITCyuTKR
gwtw/P9yLc0H6DlHg+p2q6QhSH2kdpkfNKBOuiLHeMdk53pVpNq3jKsjW26oTQ7D
aPX0IOTo/1jpIs+fY2AnOhKDttS6cv9NFUVlLDKlq/3UpPRPLc4+8dTjbtgv3vLl
ap+gsDJcfnzVAlALmV4h4fYwzPQRbirkR+QoXk0CVq6WTug2Rr/RUIUxOFqwlc2i
wtohwBMj6VURNF+DHZ6Z1Ntmri2baCuYj33MZ9D2p/+E4YI0hL04aPBui4UOMFj9
+37Uroxyxyw4OvfQEDNVvlVRggoXtCwlwn+Q3X6hK135S+ZWXVHn7CPZiY+YGQtB
g8RZjQ/Wo/xYChconC6MNm8hwU96/aodGStdHdoY7VIkVbnpxng6TrcwYsAZmjkl
h7ZhmdC7EgpQD1aD/BpJoW3A3LLPZIUlWfnNrJQ5P07nFVSel1lQwdCx42CSSnh1
7uuuy6CRWMOm6s7uJveI8cMDK7tw9kEbymhWdCgsuEEiGTyAfXIrMB+rGicXfAoB
w4p9i+ub0e2RaLytUKmlWvPZvqLqUtOxk53O/9Q+dv2/md/BWMAtyTGO1zmnUH1R
EJtVqOL6SRzkh6JwYwX06M94+jJO/MElQZD35scUIrwYcBcpCXcwDQB55HCxMj2L
9dug4p4apuXkfbvl9iSg67wEDn8JnPbYO2gqZMMb1ThY9kFurg1dU7owtcMZza7/
Ahl2GeMUlLaQ2WQ1bT2yQMF+06Oodkk5y+WqCYk7LgrIcZV5F6QTJTM1wwfixGBI
ymjoCJTmKK4L2iOTaEfkfMp0zbNUQU6kyrVdIeKWEi2gnBQvhfvtKqme+Ol8IYT5
8wLjlidNWjaJLgPggzW0vS+lRoIsKfQYVuBGqYPC4OZAtMays0p+bzuulvhSzTMy
ASOWC3j+jwpOLg0Mi2I+PtBFrIB0UJ9IvMqW4CMLegjl8aw5jdZvcOkIktv6tCji
klIUXZ4FJ3wfFyWV5m3jafH93fUcYdKdE+z3ZSHMo/yeW1wyQvAFX2DOu2HtoZca
/KW2kO9X0Lb9F6Hvsmyrmy2BNHZx9Onl+CvL83NCiyTiuAp+9zeoVKRZ8R7M4uxV
VvU/X0m8i7FYzFep33Dl5vwiL/VkS+O772szTaG8OqQaYsFvydkaPmASvgODr6P7
VdjV0zshQhxoI59Q8A8rSdukaOwOEwIBM83fAcwe+BSHwJvbcLqeAOeVlGvznz8V
uU01msSi0MZYAfaN2jih+7je9b60TlR6CAkJk5/VtKjAm7iPCIxTL/TB8+zgPfUY
zU57QgmdlNr9t5299ijLc5IAEBZJobqH/+A39RbPOJnwkJMmrf25Jt0TaDRydJ3q
7SSgMIx7RDuzaxiSy1Etn8o5gd92/semzww18L4HtHG4AyGRx01/s9Ohl00HiGkF
P+ZqmrN9cCRpc5yb4kHrkrJvOgZPOgx27navfUAvDibUet7AgiI0zAlin5n5liRP
ziPK7m6gHbih7gt77BZU2EAJGBZFPChtrNJs11u6JieWDJaltrPH2kHXtC3/hHPt
5IM9/sNKTxgGFqeyHgozzctNgcYEkl8FDMRwEC03kjJ7PQ+Anl4yeAR+Tf4QNGYd
bGBPdKJPEyxO/Xx8gThhbG0l+vfz9Bmbmq46DP2K7WuXVWLmJW2kQ2ruk2W9UISn
tSfILVIVaxypoxZUWI1BBf8EDQEfkFvkBwOXuFRfwJ1u80QBPrdnJGCHv4geaFqm
kXvgSWgaLk/OOlzba174y5bdrAKm4PLRY8GmvuUcuu/0YSkRDRBbThK2y3qGlWEv
YxOAegVqu/Yyg++JH4vJhbYhzUfhCNA/ynIzHDF76U0jrm9xM0C9BmCSn0H4kVV+
wOkoBXg6vou8b9o+E5ud2EuZneVF1oqENBBUFdfYz3HpZe1QaesxUQ9C+LDVwI6h
kmJWKSgDC6LlG499LyDLNphudSxhHeTAtioXgjJssySj958smL+b7sbpEgRSuDyK
e+VCVRuicwKHoT47Znvaf7k8PV0Ol4QGW+ZUm1cZE/7axVueZtTXyqlk4qQdDnXS
IHmm57fQ1P1GoN3o0Od3+ORrGQlgK3Q4pjYuh+Pr7QaQ+AUDyhj6xpRxXroImzoQ
gVcxnsDxm48DwQ4frO3ArAqWUh/7y+6ZKsg5MBNJQKKhFWdDjXdZrDNEEEWgQjkf
XB3gQbvxbiYYfZNpkjYVmS8sy3tFpUXsE2phVYwQ89VMkuhA6TpIif3KiL6OJ+cm
YmeJCe3tgBhg/7VEOz3qXvfgNs1c142zmstR2ARXaN2YxxKk9Js0f6AlgEhqSrNC
MTo4QwckId7Jo9s0zyFPsiOugpNN43gi2UkYcAv10GNX+XInZsaE7iTO7dGo3tH4
AKNb9QrjC/Min3nqcjS+JnGQwl2mG/uHzY82L2w1U9PPzxJviSWMhilMVfBTsDv/
Rxbq+TosG1rkNPahxXwDpHTIMRg7nRw8s2hsiDV6VfhLI8lQ3olxzzCJLinivEQX
0v7VZBpfnWUETMjWPd8UXJkI9r2uOpCk0U0r4xGPipnJGLKde3zDRRy4Z9g/fm+X
xkNHewHrnjFxPQohfpI1Fc73OXb5y7vySPZrla1LHtnCetvPEyo1lAw3vlDNbAkQ
iazmW3ZOsGaFpOFD7nmFgrXvGJW/ywKorFMk+jJINE+pgh3rfwYjTRURjcJsKR3T
p2uaBHJrqWAbJmc7dxL95eRdKaEndv1rsD7aEhC6e7tjoUo0uwuEMyvM92sIpsxa
JuyVA1+bdndhLTI3zxyHU+4o233a34qhWwUIn1wY68sp956QHIHjkib3hyx1cAk8
7BXr/yCUc7gE9CVfeEidTDcCUQP3ev2oTnLXdzkRCkw/jridR+zio/aSuulx6aQy
M3l99y6Q5ynTPZzbjLS1mOw9iTzIuN3b8kM60/LJoy8XfzTprivTaSxqUXDsMXDu
TapNVEG+WVbAyjonWoneuLKcwP4t4VxBvWfrkH2YtnMJD6qg7X0a+5JCXs5BeOwh
hpXXjEBndx+xooKQuQl1p0lrv+XtIzyDZHhLdAAlddncldB9hJRC+eZEr2DRH5ko
SucRfxgsqW7VEY0D+cPHp28G5Y6DEq+V3S2oOd2D5CXjtqPz/8ExjjSXz7oXIV47
gLJB93P/thONBAILBumw/PWTe3umEYW3OPLI9QQQBPjcCD+KH/dcW/MXyLv2Uw+k
RF/blwoMEjn1Mt249QUPhb9/Dw0B3I+OaqvlXkOhQgM9QK7JTnZZUuL4A7hLs/Fe
E3J35fbVY3ejYYdqFEo3g3FL3w0NUWGAXs3S7KKTO3lubub0kskVPiuV/28QJrrY
29mb3CoNrGpw94csUzYDkOcRHOUYF37B0BKBcocWwiv3fSgvHdYmfeWv6u6ZKgNS
ODRt1u8ZedJxDQQPXy6xBePKelkEuu+QyZgGAcgk5vJ/+E1TJVruHdovJ8vBNOI6
bSbKJ5g1Ym6ifvxmWOPQXKs3dveZ7vRVZmFdGwjQvE2Q0FpCEyv8wEjenqOc7TzV
m6un/26XgWm796dGXzVUufaIx+35OGPqtM94TF5VraTqpZEMLCfuY0zjHDieEqY+
plFd2CWfcYArFecR2Vc5/Faz30bKfGKR5X7RytkDgMVfXyi5cZF+21xhDf9RVevX
ejcMyqYZcdn45cKTVz84Z8h5sxIKP1v/MkPStstb+MmB3roo+ARE4vVFSfKC4HIZ
YLVlpe8V2JAtRVQtFsRre0wG5ptx50f1GcZ/uBYYc34TDvR/5pryhOBPGdvqkbbE
CI4VQeip+NFOXhoGUIB6hx+7zeK/JIGjwIXy1MZFqvHJbi4JXlucLj3h8cBMAsXg
MKjuRO/LABAFM/2YwcnA09An2FPx+SJeIm6fHXRcfp1Pus9OpcfUKOAUTVTApPmu
lW63sb9r8Qe3ZvcHM6GavtDquOr2tA8C5uL/8hFkTyhSwPlTDCrMTOZDsuunmPM2
7fJ6+rTgphBNbJ7YRVrODHYpZnAtw92O/coEssx3aQvRfnc/L6nJ3714PoAJKrd0
Wpbzv53g91uVXA9OATfHwO0riZrtjt3WFOHEQ7w5PXFjL2Yi2Y3LZzdljWylOQlZ
++ECtY2o4UMDMC1GesM3fVU4rtMTBdC/TSHPcJDLT7CrmyrgKKM9cJKGox4Rb0+z
6nfzCu5PLLR5AdlwuxWizYElyiB9na816MpTlCE9Gr5xZfi06xsAGsHEiF3AyjWi
mtlGIbTG6ZjPpAXxOQKP8dfYsjVFUlt0EVyo10B4SssrsW893t5JeBoVI0vJDP9J
LFQ2bwVUNdV3sv51jTxLFRDJns6TlMPN+UiEdof7SvQ5mzGZBuhD5FM5mc/s3Rjd
mtheI7EYO3+FhD/8sMoaEeoYZgGmmiyWJIg9U0IjnltPmgJgQmxQuXN5XrrPLExh
E2sIOq/yWxml3ViyJrmhLLJL9PvD+uusxioZ2VmQ8Ljsyx17pjL9BwD5zjDMUT3o
IWCAsx+pMpH905i5i/X/NH6mZjY14/gfmuE/VLQuG8c2RlFRv3XHEablK70AqH3n
cWbzdbgTzUx3oaLBaoGfF2Zl0hRNUM8tHYyK3Yd8YNl7e5FvheJ5V1lmoteTmU2R
blTRW7jt6l9n/dECD0Y7QCvcEQYAOqaY8kdcz9HjTgUGY7e0j8yCA6AKq4D5Ec8V
M72f7b8Non753iYXR4dfVFAMIwMrnQVVizDIR6n4EuJKw/VmM/X8Dejt5dTxhU9R
iNNKLMK5/IIVQnvKOKemxNcZuob8+6i+OBIit9V8knq/jYKXPh0vgzIWz5kYange
ldKuXSM+L5xkb8sv3dYWvxDvatyFD1iXg9MD0986H+KGeQRhk++2L6d+fs+KCjbn
t5CUdt2n08g46G34MnYe9ShGEVvCTYaHUXPSG4Ma8iT7wqh0d8/mZ4WJmOhTabTp
aA4DcqvRl7ANA4/OoDrbgPbqhqdo5K5L/xlPJMiVzvjbFBIPA+4WzxQIxehwfY0V
LDSbCA4mW5bOL5IFdlPBQsdgIxn39wAa70ndgHVIJgGfposQKk3FQIifBqrvn6ha
si2Moquo3DKSW0WQB8TNdkILPIMWdvcQ2G97S0dGq+2hoL4hW1bmq92FjpXOpBEt
ErTltwwupwQgJYuj/Gg/nTsspe1CAoDaJUuKsSXv8Cm1/5mZgXNovfucnNB1UzUt
9iNAoP2gozTQTdXvZexf3rp4/RwxcSsCf0lLotrL1B0ki9JtOhn08Bvmo2WTSGCD
GPeiS9Rc3DLJz9zLlQUY1N4574qqSiKqGswDQv6h8cb8QeYdKIXWRLzQkGykz+tq
yZxKPmIESbITxWaymKsembno4aRaWaRvIrmqVxdMO7Ha98pfQiDD/Up3uvg/VJ8w
sNJpFIPyS2PQFDsZofEEBfwPcC1wPMhehQg8S7g6BFhtfkQ5AndChhL/b/3agLYS
u3W5sDMGZ4GQvHkoil9zie2//8n5jlYTsWjq8xqSjM570/xkTPGqSBoRN632/DRl
5rEvt78EjveTMssiAMnUeeeQdGToRKHBAiNRa2y9uRKXXm7aMNs39FTkYyJjUrOG
80r8nK9dzAtpNlg/qjBfIHPvOI0rbYAFCG98UiJIjRhxGWTXIcVd7QE1hCkpmDnM
EWHGtZf1xX6cEqs5DwsTSQteOLcCpLwK9Aajvh8KB9Wi0Nilcp1XpLion2DPCDyL
nR3BlBAahpk5rRxtNQbzrvD+KHwzHywS7mOqlisfcSHA5iAEeo+TCipn9R5YIc2Y
y8YlLiGMmCpIA3Zct2ZumUG1U1S4MwG//aLEPgTIkcego/Dl2STnOt+iIian91m1
jCGVW9u3GKaIYqaTTnuM7taokUJj3P6hgYA0NCivtF5LHyriPSQmJ3n7LoF917+8
38i5zIczlnfnCwP6WtbNPdmsuwyOgBedJtQR3iz15aAAgtk/FMBaal6qlqyxS/7e
oY48Rk1+rMyPCwHfnbWVVjq6COFqRSK/RsH5bI2pdmgnEqn7xwgUMwjrlayEpQzf
7EXXp0E0RbjdJzIw8Xr+MmKeSZdmu1gHhVj8dZKsiNwPMzSF2o2rGGEu0yUlCA9a
Bw8Rzebx74Cr2WexhQKy8tobFe5d4hCBiH7PY9vJe2zLTBONdeE9N+wdB954qzXj
osDpwFJgNciLmpxK9mk3/JcD2BVbInO6FgWL1+xlLwTsf9mU3pp1auScoq++COMe
qYv2GOgTS9hd+ZAntT92TH83d7Yb6isNMIiBYTvdcl+55Lz6lsjtYIf/qZmYjY6o
UP3niaVtAeEnJHjn7julUZEo8asiollfKQBmf/EMly0it466dIwgFu+mOeI5QUOq
NNTMcUiZDIZBvT3fIy9cCHZ4lDNd25OsRAzCAPgXG1KPQ32XeXHS8bQr9mZivEht
7rI7T7qp3OlQWJ8CPpaPEWCHOyflBEoPj6dRV8bOhNPKMiQs0pW+vJI1QWhVZK2X
0FMe5p0EENVIlhAAQsTdtb8LxjOaRtwQWPKXPfufqp682YAkvVA4y9B/4ZJXA6ZO
whbWfJjYWdNv/HNvWBRhPRN+/8WC+/9LgyJTxSFc6B+mvbWEdh3sUf2OXuaaod0M
+KjgMAnrXAE4uiD59Qt7gyAWEHe4vtjMJrWyoLrE5j2+j5bKSlB14fJgz+7lYfC7
PHm1WHlRexRkC6Ch++OOWInO2pfyI6xy9WRYUNZWrJF7CrJm+tX5Rg1UT5LYyMcz
51JphPHX3jyTbb5M/HMnMc4BNkpMBoW2bdcYnQMbxqrinsA0dcjd/RZE6zbFt6hg
W0nuqkQKFqxTbW0L9jAcva2N+mvG++oYJCEQzTIaTE8wbU68uSpTxveIabrxRjC0
5NcfcYph959yWWP+MLikZx0n5ku034v3HEgw6ZuS+gK4mKfXmvRO9wwztZCSmYzL
zLBErcnGa6AK8dQ88Bg99SeCP+6AZ4OlhTEJ4Vqfw50KdYcGgzRROQ3KS7LJ2An1
zaZzGPVDORhmzgn4ljt4IUHCSN5ESzLmuqZ8UElLa7jLWmvP4MQTWXQW32lBXvxX
ZlSqoBZT5rVX1duSjH+sLyQr+vLPQ9OWP6k8YUVCfBnDcGS6C+psY3nhpAazSUDU
oxe4OYHQOQSRNOeaiDPG5vFkynf3IS+BJ+ul2dv3T0HPjznKfEyIBSZo8C0j0gEv
L+qIjyl9cX7Ch1zE9D6KaXYdOKrkseXnHKrzKcdmTtU1jn9+0LF50Z+ySiegVA4Q
dMvctElNyomKssGU+AFZ3T6cZnUgzRHu4K/4OIhWCdOMNRLkB4Bob5C7+3axMrhj
hg3A3EX2p122iIFFqa3p8n0UwR+9VLKYyj4EHya/ymA4i6BgyAB3bWYBq5keyO/t
ilfHLz44ZKM+WqENtNQ5LrXaa+bID2mtyTXmE7F3anekOWZtK4jLmPc8f97FTTvR
PreqOHgDU8zopHr998v2ZvhO0C9/zt+fgO9itO1IogidDtilamhgBKYoPeexh1Vk
0HpygW08dxLsKsV/T/l6s7qosLdhKIBjuuzJPMdEE5gV0dapEo2hKXwY7NOgiVJi
QXHQm/j4kB2Oe/vf5N+mEIWbQmC1FBOvP006EnA3/vlGgJzt0B7Qp0vmbMOGA0p+
SCJfauA2olvic8rQ56PUs9t4FxYrWXB1CkUR3biqAWHAHXrU50R88rtdnSrTO/ne
k+z3BjOeKk+WM68Pnzgsx2BJ01klo29kZahwe2W2mZ9ZIWaXw5nzvkHQxJHimi6e
wt9ZO7I9Ga9aB+AFk7T90XwF2auCXLg2rz/X2JYNX713sfJCxRDiRqIvPlva/hpT
sxxbF7YdCtRzbi4fFdgLpzuEkNuR5VNN+nWXYymB/YxiS+HmMAXkMHUvSxIy1jz3
AgYlMyICnLU1cxO+hEx8fH5lCADoZkVQspMlJpVTDfaIuDbhdjl3rkNYj4g/lcje
oVfIqirEZSrJMTMj4vIdiLsz5f91qyflfvkvAVjg5UwwvUmkHfE52Gd8/V7c9I5U
694lKK/7sPA/s2pe+TJqfb5VwoaZwtkW31jzf4O3JwNgyOZOyjpJv+7MSgb6B62S
C+CxGRB5lknJ+e15npx8v5lQlAPzPweDYywnqxK5Z28yRPy5BkYoSLsHJbBZ3TPL
Uo7ioDLXQoFeWY43+hwrDWVNR7jr8UHDpyFTM7hLIhwpQ+4O7TQwOPwbqTmCG8xv
5dy9ACcgLKqDbbmwgmGJgzujrj9/dbSEd2xsKhP85G808LxysGTaZCbxViGqYtFN
gAsXpntQI5G/IpYhue82CkN+kVcEq8PwfSOuufaC5PK1IdeAXWTOI5UChBe+sfHW
wD0flg2ibTYLg73fAER97Re1EwJY8iM28q4uh2nFykIsbMMa7CAJZqHk8gsDrTVs
NdAVJPsFGYE7kIOnCkI4H2N8oPw7ftOvu+5TQEDfG2tt3N6aCGN9kxuUMfwYcR8Z
zzX+OzxQ8hp06Kq6h21R25nnMu/T4Egf+X5x71vLQGrGcKy5JQ8cA4GaPDvJto3P
1UhY1rkhzAukWHL0S949/PQ7VqAB+ZJ68bwhEBo02GdOnGKT6di55KRt+sc05PGr
KIz7gQ1hhyhcB3KkAGTdCmDhyhELS1/+6u3gjtc1Uwd6/iT6AMPUXkvMxCqiY+Qm
D7Sg5VR0CeVVXRCfpFkegXLeyaoVAAJXgKYM5xuasSHWm77E45t82dQbRsbFA6tI
aTVK9S+GKnisvxT+JA1PIDZ8Iq1qurcb5gt9eFS+QjbUL5UkuIDJw9udvMAcbyzK
myjgiXqLPMf+P+P46ii+rAUzLs5wtdqzFzFVGFbiDtwxXTlrlMc5TnuEHsINqd36
vZMsHk2C52RyNHvvzrfRnJdywJ19aP0Ay2J7r+V55iJn0kbIwFMgF2ahUlZzGKqZ
klaz7ImN+T+2KByehi8ANKFiX0FD/k1q2dcDZVe6/szDhPaIEekGwnplmO3hjHyN
ld8z+BHfw9F8VwytqkYixYaRsBhhmFvRQEpG7NHlUsHnSDdeXu7p7ScZACLWo5vo
LTko1OKnPUNP9u41oSO1QvX67j6ddnH3XX+MdrF54VPIPB7WF3J/ykDEbnak7oyM
dqhx+IIyeDDKeY4/q8X2YTaSimfoCLrymDSEk4yJMuOQ6N65EvgyrgdJCb6asoDh
113yezu2K7z4xGRSNud5smt8VYr2TaNNeCO4lmaBv8pW4+MeJ64D/l4nBfxeVkbT
gV+J9LzxH22oguwptoEX+errmGNKPxTCYpciQ7zVGgkR80y6fPgemE8BF8yJz4C1
09PVrTFoI/iSb53yGm+URdHCXOV+K9yQ7TvfTbY6p5kDiEd0hZv6FTN86liRh57T
KHy1rgHKP2xNT0U5CVxpWy3d3pIF6rmm0tsRQh6sWoRJU6LoCBFM7UVwzeNeps3W
/pb+BBTqq3vgLM5ahziKp8gCcoqEWD/TyUAS5e9/HQtarlCPGGuDNpxYCowItOj+
MD8Ehk20YDpPj/kubfrTjirRTXpOBkh4vHlGzQPC3gVC1Ugz9JjXVl0HJ5u3mMr0
zpVoCbhSY+gW2WHMjKu/kBVBW/Qk6hc7D4fa589ClW4+/W78SpUkaSo1cfawf9yf
WHl037y0wYFubGaO+Uh66NUJN2W3KFaDJRRu/5XFIkUHF21jNOOM8U0fB8DFukqQ
N5fcPTX1PETnVim7M0LRIgcXZBnF8eYxIzU2YRO4onCHSF7L9ygQByMZSPw5aSaI
W912Ta9eg2DJS7yMDXlY75G/mLpV0OwzUu5Jd41LEMZROQD/rPNliysHq/mf5aMC
Zf5wsp8UJMQWJTfTYs/8m1XOnkQ8hTjZtZz5a7g5pABv7YidOy1/0lgTPWoKrXUA
+Fl/yZKpVyQ7tFUd3DLnDui8VjEP8H4VRVEYS/3a3O4D4q+MDs+0nBPgqQkjTxRd
va7CULZfhdGbEVt0QE1HUUEGCO8WRRXcZbmAg4hjwpEcFTuRdbC4Sy5aG9lmo4qg
/uYszrSZeydLL0KAfJgoT4rHV9Qsc8PHn3kSRLWC3cx6aRQaXTvO6FbKplDJf00x
OxCdjPDjN2ZCmgkqXOsWiyFN0JWB6URQO/GMsW8XiAFnllo5fMp0iUTfesAc0/1g
0vjBXFj7CFuTo9Xde7wSZkrWvdiJWvyDFRilMuKvl0loc8vMvcOYi+H62TbCpdNn
mBps88hvQQdbFw6KfJiVZu3DQC30kfFUYfI8diDFZRfMuB3mQd7+jkgUd9SFmg/w
K129yUUCi3Tzxer3Tq7WV34+sBoxdOswtnU+zaf/BjaebeJhVr79Vu5LfNWd8HyA
OaVQVHiJ3IUMDiANV4UaiXExUfsUuXLxRgJnf/DMxj7JQSaXFPhItmyfokJZBZzZ
WURWCpFKalFnfJCddcaIkjFoQvremOoY7YA90DD2audQ2cEPEVe4ZINaygnYDeFh
sc+dFXaPf2qALLUQvFIgWWIC7wzplsT1sz+8E9dudgVXbJltI3LPz9THFPTeOQkv
G6dyZYGShgmHvsoc5qIdH178CwUX61IhaOiWLcxY2CumONE8tfWyZ+uK0w2HhEpT
cMzX6eG37sRm/STg4vfo7CHbhH4ADwkLwWamYbEP9suQKbdOkuhXIewqLHz8DnXl
EDcQXhVjFkDqGkWlcf3ZSXEfRUuRmjlrjhZrEG/1UKPdhE1OFLzK2jivpAobnipO
i5dGtNgTSy2nEGB/8rqeaU4KuL7WKQ8XBiz8C04B5+ZMv09f5mb37aNF6U1bFFRJ
m41O9h+AiDGOpmItf0FmOVMQknKlXnPmZ5k3Pxfg5OAa4J/9WrQUKNRdTzLwU6l3
1wbvgH0QyQ4kmZyqfQ/Oi6iZlSXE6JmgwM0YhVqcD1cTYzQDpI2+vpWGHRlDCioP
taGb7CRCxIQxENpWQ6uiTIq9YDeExHhXEfj5WmidHLOrLzqs0Eoemhs/OMxwWImX
Mii5Qt9RKL0keAkph7r33N3EU+1BURh0Fz5suJlKeBwV/6Lf6Ox53ReB1icQICOk
iOWWY5pboIcZonrqAc4kd5Jo61HY6QHM7GEB+mBFHP1MXYknW+sEpY8XqIDEr44M
D2m6BhaHjQpvVeErVc19fMnhXSuNgJuowQmFpRAp95NZGNa7JNojf+BCgodwjFi/
Gb8oUYL9mvKycy0U6GPm080f2rf0NFLy01h58/7lqaxrN/LAzFjhbTuVUjQogLlQ
Twdm94oCHx6kLh2awLpcvUgRbdBfBGJjwZtJware/L92bTzdNWo506gJUwf+6Kws
XSq4kOn8y6KcG0DvTyJGoIi/GSZFyprOemknzHZFiZA5MAIYRUdyu6L3iL8BCqpj
vHkKWj4uuAYjbCWbca5QBNNotEEaMo/ASbTigB5fkCG7lPQMYOAn9Hv+38Zvva6G
qJVoh4pAcah5Elq0iDz6yGhnPJf3nz3jJ8YVfuUdJ7hccUv7cbWLqV9JCZgJW12X
VTzl6nOJM7awQQl8E0CKuY+QrnkwVOTx+5c2/nKASSMBVIAh8f4SOpkCogbAvqu4
tWufNSSXlpO6WK9Fx27/8oLoP0BufQ7KqtfptfBme2flDDsffzNlETQ1b98DNrzS
+TEy9VJ0NBa5fNIsajt5zaeY2vsv2DA9KUGGiAnTxaORwzhWBwjDFnPq7vEhj60V
dHImYhpXmWVET2nvB4Fe64ez483oradawDFFPAFxneYlxOXPrsCDeTuVPFf6dceZ
Ok53fBcpP3Ao7MglfDHoTHTmS5TejBeYHEz14Xb8RXLOKFteJNFsGG/s8AljeD+O
UluLVgO+8NkofUspIkpGjdbwS7y7juy6L0ZFed7b40ibG6k7qTzL/Yb+DXTgYQRL
BsOQTfwHnpC2MvSuhcJEVecOnEBqgOxyfX/1AK5imQrihEJmoOeSTkq2CQyari6S
ZKpHug2jTcSFZYubYSumaQCQ2js8Q1aFb7SnhAV9e3iKjxdSO+hCh4SwCnreTr0v
jymCSWZnQIDCCuusbw+2q+Rd40nmpVhmkbF1RKpsqC54GwZFMZKNVp/C18ffdf0P
dNRt9GwVlnaNFJW0fkDkP27uegiy5Kdz9HpHWoUyxCILdEnP2Zi49L21AXl8SatO
ZortdD9vtYpGnNqN85UNNuUlfP6tTOZnbgn1Er4w1lOR3+BmlN+O7aZvDAvT2MSy
2fOCMhAd04PM5NYPSk0BmUmUd/dinU6gccC95lcIlhC9bICRCce1bVOnkiT6YXox
0rpha+sj7PfmsLd7tPt4sMABO+e2zBxrgNr7RcHZBymzlo/4TQCrLc4uMIcYuJY0
YtRldOVUAkkGjHOt2kMD+WQXX4Q3uMLheDFKKsSBvJxXB94TtWuvhuHXq8ISHt4C
a5er6IpeLpOWO3VS31pL1PVSUco+W9kWc3Y0IV9lPjIXrMJIm9y3EMNJyQiTtucA
Odp8B9TJ5y1uu2d5AL1EurWmO5u1TYgdcUFCeoacg6inOHq3QWybznRfewXDoWm1
dUaMj9SEtatC4b4hTd9Whbhpt4+wBBPGq7kCMainP1d5zVgVmtmIIyUegyThsrfJ
dlBoPBQglQrp8+JCOJRg/tDIYTgoTek0GHPuIt3r5kVPMfWa0SztjJ1Y2EuAtoay
mpO9T1wLxUfKa8UVHQ7PhvlrQ8mQbJj8sOW3DxXHQcNedxGFbc28xhiPf7+wcthl
+9qHBGe9jBwj26lBWUD1DgHU3FB8KuBF13p+h4P7Qdk6UUlgW6ap6d6jUzDRFAL5
9Ve5JcFqhkpNl3aWIYDTMtg2aYGjTfsVHpXIzcFCuwGL5gQ+scXehIHsDm50hCty
t6aeZLxqwmuNP70F6d7KkXMFr/4SAqxqJkjQtACDvaK9gCFbhf7CA02M9RKpXlwd
K+dajTlxzrjancMhHIu3OrFQPEzh7ky6x3f8XpVGKpt8mm3b6neUrbcXuusBWjKA
Eccva8pEW8KGvYMf1q7VKDx45iiVM8L+OiZtVdWwSG2OCadUIIo9tyNS5uir4Mu0
7Ty3j6HpB1JEtQN+rUeO1AjRBBLpRQqm2dLCIUXm4hjvmE/JJlW13etqBKMfdq7r
Za4P6EeLY6GB9WztwEaAoGtuTyb14mdS/c3nvb4Npo/Z3mbAgO2SkiiSuIdne57V
OQ1eV6R77+UMSQGK0GQQsm3n9YCbGaPnm2BYAoE1+WiTY8eSHLehHnDa51jvq9Te
Nt/b+10OSZg3tlBdOJ6oKmadUi3WcBgaPhHWvKa4kyVfGVXc2sILKud9kmE5xRYE
vuFjN7tm+bkHi9fjuES/8CPXprtPDcGcqe+wF7CyQVhrzOfFA8YFMfBIZepk5LJb
tOVL2QDSaCEA+oRUXF9iSU/GtUI5EKujqpHuyAzN9ItBEfV2uladf2hxOMDAxiU/
3gU+Gq1FiQ/4PKCmtyJZQuO5UCxkIaVoTZ5kvhfoXbfrFOR2fFjL0QuEzfzVMRbI
syStbHFn8iicCcAR6QyEVKe6ukkheG9vo4AK9yvx71DfxHdx9xWfwMoATQrGgFGY
bqSI89d7MdjyYGnirxkj20raqJD4QuCQsMFR0gvsza1DwylbBIHbE/JIMrzxNV4b
+adXLrXCUX1/21G6/pDqP8CivlYyIPqRI2txXMmpqoG6uRPHpOjr2g6UXsbChBAy
pVutMxKp5uH5X1E9714E3UmuAmBOpg6plQeXRc5rfDokwL9CCriGIceFMq6LyeB4
jGZgbeG3SofWCpsN+xV0PpRdGBiQBVfNxkVlSUFUtS17U8AhhX+wUQjnjNFbbSO0
xGVitaZ9uNXmPkj7QGRh94GNcj3rUEq3rkPBsfgW24RsbEFUl0fcUoiPrcxK5K7o
GwIej4ejb9DkhNjC8j2pdnP5DV4S7d1fHtaHpQy/CLLQWsdCG9CHkcwDxfx4o+UV
yUNKQ49fA1l5cYaavwAgN+UN1zsBftTAWIEnHcjB7hJm4hMW/yzs0222eAZegaDX
D3E2Psfcy/Iaq0xMCzfRTgOu6GMlG2wIvcX75sNNNl/YTt3/kU8vA602JqJwTynM
7fVd9DptzTVWTLBH2oV3txW8yM4Em5vM6MtQM+6v8ErJXgC/+SuyL+rvHb/W568v
vso6w1dQk7/JrVtTYQ8POUPzpXbIUs2TwXPYEZ6pOfeQ2B03yML27ctQoTTtGL4P
tTutdES7Ol5wIqlIYZ/wp29Y+QDQnRLC5+ulLltaz3ZiRVTwlrC4aAfFcBUzVEOH
a1R3/xKDZamqelSU4JaOQYd+As+mgNgYOAoZHdQHeNZHkjl4DcZomKn/lT15NsMM
r7aB+1KOEi3q1nwonoU788+6wrpvZ/ttUeh6ZJNfQsl5PjyTIH2zj4058YXZyn30
fmM9o6cbAgdqWCTsDESRX/AStb8xy3wp64xk5CyVRpymq3I0M0mRrTr+QJx+FXUy
U34Oxh96mVdy+YoBANtdft4n/k+flHIaGKH3OGSdWKzAWxKzqy3oE3mmmndV+MJo
Wbib00pDfk+Y/P1jZb2BRoTCLdsGhiYDOaSMTG24wNrl+KTrwvY2XvwWJju1Ri2P
erV1wlkNonAuvzXFzWMGUCNX6v/SAdaj5DCG3JoaoAUuRTwLvGRQkLQbu+uNf5Cm
9VvQSUck5zze1rzhvYJ3aZgDB/RMoPTnl1JpXzSVoUXXVSYokSF0gXpjreyB1oTl
556bnM3kbINERA01xWedibAk0/SdCmDy1Rknl9Rv4f3z7mV0tX9/1lCf6dh1w64d
NN1EJaGT3mj3/aqvCcJvq/etslCYT6pufQeiB0wisicts5Ruub7pUse51jNgk+3z
f0BOP1q2LOzKuiDrD3/uJlHTgDwcnvtFaGM+8/0i+Cx8/OUZAe2pZzDu9S0wLPEs
GXKgGaX4KfNuu20eemDJGyLnh1SA3uEy7eOznHQN+ilpOucLUU2vqOwkFMu/LCtz
ibqhHWOVtDqmKF3Teqv76PwX4/dcpLMiMEyocl5fYRWzAL0lJ38mCDDNsrfJle8M
1u5kWJAW6I0WRclg1vjlI7sNbj2JTW50pstDXR7N2TNFf2/MWHAf2xflpprN8P1J
6C07DXmGFchXsBavBfIgV+BgWGjnBGU6tx9kDlPIGgIApIiwunS0EZC82QHNmvmw
BLgxye6qYle2arrPfebJg1/4eo3WubllMhRRukz1j7EQUXcqsyCXKz4YCX2pQR4h
dcNR1zv8/K4f2BZd2v3E4DKkmIEqd5x9/Vpr15dn9EJfUWVyE4rBxwPq99xadrs+
Acdn2MCmipFo3wUzU/DxTNpo5C3HwsEDaqCfkRXro07NquHoUlJYmOPKEHy32EuJ
IP5qjdR+gQVfkbJvAwj98EElkKDbaCcIW8CJfoz1ts9G/omdqYFlAb98AFfsADG1
ZdmwQijkCA7lJqgROx3Y00f2Rf3A6gpg2SXsq6CTtbSiPHQ/iuohxERUuqU4VY29
8eLxSebJXVPAH5wTP+hPohPNHIc25RYcEiFdUPDt5J0GFDoEClmH+4l2yE8qmJE0
SwXlI85H2N7WfEojzMT5vWNWkfzJQ5pPgO6/vIoeZh9RkBplSVdk/mpSlmftMGbu
0wS/8Ls7lNPmZNMSzXBy2IZzYoDBcv5NYBUXFnEbOR0O0p61qGLQE/bvHURE/THB
5KIsGBA9gNH9htcn7d8ETp0Ffui3dXmBK87dDijqzeDxJzcIk8gpB/kcF5Suq3m1
kmx3FwL7Z+fImxXohnWWDforJMyUhX8cm81NrOkb3AbimpsKRH8btsE4xsQqX7Op
LZB7XwGgQmAIc0xru7bk3IhIHmM1vVuG64rJ6ujBR5mpNXcZ5s5d1hkQkR2feWae
MwSfbcavlihQSn4CQKfZxqxueQyN/JayrL3AOSN5FcIH72jMrSVKJWwZODmL7hLW
o8yNbr5/sO2OgzB/ItooRhh+LIUOdlQWz7ovwRX927endGAoSC2Isfh/8IhLQOI3
evHwaqCiFq3qGB1F+0EQ8SS+QysIrDry9zB/199igGy2Y+AVtGqNySxZKbs9hwtT
urZFadRqBv1Wz8dDzLPjGdhKWypXjisUrrcNYgXSRAMAJq+w+DR40Sm4gDRg+3Du
i9gn/+5minVbtOK/qAIY6PDNPn63OIIdZq7LYEMQQQ9OjwfQoUr/8lb1XwfeQLTF
mbdmQbrZD/izS2dALp0mqbF66KprdQ0zq5f62nZqzMkEQyKg0of2QxEG7YFfPYHY
JF2EcWRIUfhAFJjgxOrsZNmbCY3rX+j6NFet0e52jDQYdyi3SH5MA4RkJHiaJWcV
nv+Us2HCNWFi80owuxo4TEOsuUL4SN6pNlxQPo9RYrLuPX2zlkWcqpAsfTtfcOJN
/z0HY4CvPYJD/YOStE8oMXz84mxYn1M5RvVMRZ0YVc5h3T58p1q8u1s+4BUM+I0T
YyvPOdc0gQebZZTykWRHhsAtmFc+hXdNxa5kBgyn9r6zCC9+7WC+AhKjKNipS44s
WkoI9IYbUbNNC/+bCve0TBvC19OoC3C1OjWeJMqkmgJ5BqELJXwWrB+OlxyWobB9
cFFGeoT5/eborHEGTNB2l+r4kQcgOgBxwBOt1WzW8hTrpgxTWM9pvzf+C1xJq6HC
LYlixJmiNpxt+u4Mm3RrPcerTUL8mPJxCvJErRqK21GRY5WFhFjNuaXIR8J11rDU
CcKQbfKdHxl1nWBFBX4VpPiVYQwd7bmuegObHLaHgfhS1tX5wYdGE8kQivn/cwqo
hn6Vrw0yCVYgrxogC7CY/Cs3DUOzJ23yxvm6CnPQ1PMlrDMNX8yWuMEEBp+0RZIn
tFOHoOFqkNZM+Q+E5HMaHUq0ybhTSMP3B2NLMgLOyvwMSIjhZOKtaO/b3r/N/j1K
04ojuuWc6cRFVzBmx3nt5bTVCTW23XfdsozIAL4X8aiMXiOBh1XzprZrBKg/tkkR
m+3ev6it992KUeROrmYn0thp7EYJjtwQJ//8/1zpuWurPU3KnfIxbLSKlzeTmROx
xAXfUP3xR5p6BvUN2+5S1eDnfuoo6kNzTLj3lsUXfDYnHRhVp5xZMXzdT8lIqVyw
vU9kU44elpPP6fyCpDP5yeYrLFc2zKb/+xbic44HxCtJEFcTaOSalfyurFwJjzaS
X7trOmKPpT44aYcq/ox0um0ZD3Jkhd4oeokR/xnKfY0ZqJwB2v4UiEeBhznVTWK3
/s81LLxxlUj90P9zWPlAgC0E/9pXLkwfJw/nILi7gR6zO/jiRA0hBNzdVdL/48Wg
KZZkaW/T/wBtCf4epsTS561jdfmep42qGj132+qwTtRAalc4F/j8VuDHQqpGi6oh
pOjJTTCn9lzsgj8ZWFCumM4uvP6p2LJvvLvow3M9/Q68tAOLWtBtBCmZtrSn1pih
a7nzluwGP7ttmPQ4GMRH4UUQg9zO9b2egq4EpUFh2huf5AfZoq2CUMLL1O86qdLN
dUZz1ckl0S5KgPBwGNc1hxxWF8ygMPhKUyse4W9crDwMhrUc8Y57uMRzlRqfpoaw
ynAYtzHzoSA3MJZ/wmt/Z1Q1EUkB90JGKPyNi9qcuMjUk7vlI8JnaXVrOCFFJVF1
IsffTNFyYoKuxYv1tBt31fmh7RrdeaUxt8RzX6q5uRhOLFSNOV6iFXRBxygqhq6A
IR68hRhXtkCRCWnwsmYkhVzXeWQBW3aEElyOva5dy+7RujAQe/fyG4+xxJrzZ2bC
H1AbwCiyB9kAKu/fUr0WUeq7R2Bahe+vL8zwqQrM7PARpgWSGrNVC+O0+edLL0g5
myK0vPw6KhSP03jOPgqbBMfCP5LSnPoEc6LjTEApD6GY7mcnmZI8qRZDMlpSSBjY
D6iTssucEVNScmhxb1+RCSu624S05fzpJlyMAFwmtZ2+aJgJhm8VfccAZiLkn5IP
QR7wlie2yo+PWR2JWyG3TbgWJ+pFAFdRoR9FuTOJf+uHNaRcjCpSRNzDqVdcn/Hn
HLZD+yf8YCIx309wRJWD/CqFOligZvAKeXNGArt6clnlB+etvo+lHIp4W7qdiNUe
NirGha3oZdfcfCeuesxDxRGpqEijGJeWViGx68ivANzlDkVv+gLqHX3qZTclM88k
8mhHqeIH88JPBy2ru5gYLrhjHcfiYKiYOdfCPlXMW08dLQDvlCBvutFgyRoz7Z/C
OTmr504sM3BBE8DPZwY1v6T1d/1YjlXuMDMzeTkHCz/cdQFJkx8vXkq7s2QRbKkH
MJgBsymIexa59yPSRGeZAIROfmFnhKfZbeODoAARQhH9D+bXdUzspZJG829uUBq7
FnJcL3Qgp2BxBCQgyRe9mac9VTCri5uuQHLFWDhtGkY=
`pragma protect end_protected
