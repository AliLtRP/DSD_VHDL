// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:21 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OmGs5WiihOEIoXu6U5q/2btLZp4QJDZ9iULugfHzdgAF+7VLZsK/vPjgPDBbd1Tf
KdK92xf2dn9HW5wEhXGzcxvQZhlVwLqDZdsGZBiYWWx7It6+W9UHttCWLoOt0qct
1KPSc8T5R/YqGZf6vk4FBgO+UZlZSCOmNDdlRuUKNPE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26384)
m3X5l+5o8Rue8PF+UMaPlppWchWL6b3us0NZV5G1gNeZKEvG+X6x3AomLTLieeE3
ff5WLZeAV0xoRuJtp4B8jjeZ4hj4eRbYRQt9QmRI0li/04NTp6eDFuw+/NAm3ckV
nolHbUOOQ1q2riVGCLevzrv9XF49xrcBeY6hL9NyR6gPtDJKVAsuUj6itXzMVInk
Hw4UWXDJcLbmJ0YKdW8WTgXYc2lwz2YWzSywA+i9eNmpy25/xRia3xrFdPYSVMNM
jUJrY2CSLUpjUHx1d/tS8+svWFvn2yBaO3+vxokTlljV3sZTmFnoxncRhNFUvjLW
EkimB0LiI4AmuWwCshoPwUgtMFOSm4vgxDmR24oJRgra5V3GwQb3dR5JGsfwOOeP
DKw88rv/AmQUWqIhT4SfPJlFdB0oZzkzuurfd2BvsWgQRhX9c8x4Dn/0LdNFW7LE
PWwnZcyHRToxQkYMTW8XpGcHk0WwX2IpEFMtXTgI/GriQ9+EO+82lWTTZ110sVYs
xfOqZxNpbYwh2PivE5uROmoVlUHBOkI2BOFWbsHooppmHAnIxmE/TBIM9RQg1avu
PdbOPf8IXmRUtr2G1CjfsCBVe5ocdJ4C0Wi29fi4m2j8x76zN3V9/zFGxXanizu5
S24Mp9i7NtK9RYUmIYJJRizG1B5gxFde1lIUHxRUxXb99ZiKc0ouVvLdHIDp8U5G
nPjfQR7aQs1yo+O6POCf2aEy4mA134SiNDCU8fRJ/feywstmvidzoRIAKvsW1wth
5aerI3stpoPAMn12aGptCriW7Xba/Pv6ugxjAwrDFJuqsmvvEaZ+pq2JpdX83KfN
+vMPJlUwIINqw9I9eDr/Mdc20MH3f0zoDEeie/3sSWfkpW+iIs7yxlanKktwemJq
xdMZHLycJ1jQPeJVsqetpF/IGeJ3IyNNo0TOdXDT4O5/8iC9uZJORt4qafq2ZwGa
uWLHFuEKJQzUPOS3hs8o+jqPmP0qaTJ1A93TE+ADIX/aK24vhpfjAJzFKrZEZ0B0
GeqRc3QLow2m6SVawbItBDFkrGLdFqbRZwLBZkgDxWtfx4km1WwMpMY+pWr35WlF
j19yYuRPzUr9w1Ede4vsKxuyhM5MWWqQJHMIuxJSBED1YRanRUwHa8iXZbvtTldQ
GA4PcnqLRq9MYqmzxcm1KPP81WOvZuQc6cZODaXHujLBTMb7Z2cQtAMVU7Hdn9rT
VYt0v30/8+d/SMsi32XEdUkplyPtHNd1JbXGYmFXl2hFmhGM6cIaOoUKE1ACI/hO
l9S9fVfuW8XiU2rxyteZ5a2XsZ8jN4bU7CQudY6JfxrPAXqINAJNMc8ws9nNrQ7x
GDu+2P638kAYJNq6jOD6E4z4OLRuEKdVi881dj8ubBH59CKSEsuyW+KPg3Eb8aWv
1tIW8zwx2nB+aLSI4r42e2hINOMgX3TWOxj6LyVBEikhcFX7UHWwa5ha9ETbx4FS
P5Qhaq3E6Hdyh1yCHGuqePxlT9dVmFzHKRb1QY1rEkqhAbcBAAH1pwpB3ZMA3Qhh
NhNXK7oDnYQh2XT7J50YNJEDozF1LCpnZ16YVjQHEZxB5A8lu+NqFFHodwd8YIMj
QnSZfet0hXc1vW/xbynAepyk/gzfXp0Ja+Fg4FFj6X060/MX/qr4FSzBx/iVZoU9
HXqrlIzYDOp8lv33vMthlSeLcm/tzw65em+ZloujvWH+pnMb0X54XHpZE0rQ7r/o
+NJsK00BKKuenPctXymAxh1J2Ar+nbyA/HMwSRX638B3ro4t1Lxx/9Oi4A2d12sP
ZQx4le4RWhHawRBXVsD389NAm1PC6heKT5xfkbsZq/g0UDpma9M+K5MZgs9aGcLQ
AMKCdUmYrzc1kGEBseMeb67zgHtPHTr+8Qew1TJT0W3Hxh5FdJO6Z4Lcz61fHROb
+Ea1iHzn3Y/5kjsc7mTbsOnXqh0QIXmbucdCGDEoX5wgYn4ah1QVlrFW4SIdgLId
htjaWjVKX+s2qEHzhF488Nrm9cxVyQanZxUPyOxRnErlsEQIFzc5qrp+nMyfbdPD
kb8AjXcGIuhuJ9tSL58OGUOeVHV5vV3CoADacK/Qf2d1EVm9luAAjSoYfSaHd1NU
FNvEJMaayqW2DL1ccpzfKcK9zRYQI80VKDVMV6Jn0xXUT1wCY5Gd9dC2TazSVFUt
Uv+CzOXNagG0YSk6mGAoKpHkwTJOC5alWloI/RiEjTeiEA9D0s9cch15unx+Y78a
TALO8UvPPAUMfcFdRNVqRqoiE0gftyJiMs+rWFacDCUJLNdFwC1CxbpTRY4aMixK
6XgtkzFnZi2UxTjrQW/tFQ7iBVOBM/UvP+zv4o5mE3kXUhaGpmWIXnB+/UTEIYy/
nfUb9zRc4tDxvP+ZyNSZiXO0L3xNtTeQlEfLQz9xTLYxNzspCsXw+ry8B8vRv91R
DRKff9TdHhJUZwLUIdqTMVORyF9/5SpJnQR++8FF0Dr84s4R2p9inL8sV8gqS8xd
3vywt6WNvjACBB1vP5CD+ENIhS1m81HXDyAVplVgM+X5cD7AadDIMj0nz680dPGt
mTHgIqtqJns7imzySRJYB5iM4OwxkpV2KU0VyNrL4tPXPP/Jz/t+VkVeke5wybbI
W6FeWoS/axbhdUiK0uO2pHz7fVPVRCBj4n6PIi3zlIFPXraIolRFnGLmO80lyu6N
Y9xHqLAX0v4zbhszFRudtF0dmhElflwxr2lSoPTHriwcI3ygr9XcnD6Q8riIO/Qq
GYXAQiggBjUyQTBgWA4mXUioHc7yrkbNAUhypz6tvExWLycFeAsSqVUVwHhJonJ3
ZjBh8bdk0UuhBhenkEs+9GOmagb5zr6EpKJPlaodvEQdM8x3q74oVzHCibrrCon4
A3X5Txotq+E8IV049Nk5JxoJpN0k9yUq1FSBTyJ59pICpireodmbQhqzkFeS7wNR
heQhHYPjn/CnGNjSrBOIX7e0UOh79TDkrwxk+XOqu9t2g0F8ZlfoU6GvTRJHvW0m
5Vd8qqffeJVe0PuYemmXJTKJgZtxSRhFpjDFX/fg6LS32ZLuOgZz277QhibJQArg
re9JAYMBzRFzAunGDOk5DIf0JhZWXebviiWbXCB2x4V3vlqAgR/gRvyOG5HMJcdh
8M1Ndi/FtxveNf6ehhG3UPh2lETikumF7DOwxKOv6T9+4SrgvZfAlnA/CbL6OrEU
tL0doA0Bgw7PjRzwsOhk5lknXMGMzpl0hgvaEI7ydIoyWVwUzUh66chOdCzrDHq3
0jfScVMekHEZ8e2u+zLBRXOkJfUOTjvLutuA6j7KwbERwd4O4baRgW0/93UqKVry
JDLbNN7EePH8jmk2dlcD04aFiH4mFcIKrjAiwBWCWjQRCfX5+RfrRdJNOgqLVHew
2Ep/zANqCZinfMJ2qINqyWaUhTP1hGjns4sJGmT+SBU784TQsoW6zVdrHHW/HnZN
ZqzA/r65zZ4+8zpJffLQuP8c+p/2ubkpMzabqSkR0Exwu4w0f4d8eWT4NY+RBEb/
KR++5qj4IfqF8/zPzTUqO9YQHGDAokGPUwBMyYCfQ+yN/EfJlz722fB7LTZHe7/5
dJH0ORwZX1W1nSLc5T0GmHn6UfmTDrhsutEwUj4tDGDBfqzlGGtA9xqMQBY/QLRL
7k+sDGYhDioOpW2OOsPmA8zuA0bqLk9kpSnxmiH5mg6kKD/n/Zk560ZsWJLIlPUM
MCrItHE0d/iA6snj4RLOiODGmZYCZgHtTSh4WrL2vA8PWYTtPdgjzTbC1ssGNrW4
v03VS0LXqUzn3RPsAfOcIXf71E2sAONp2DKij2Z0HDJKsQv6U/gun96uQ95+Xoat
i9n/U/BWCHt6A5g1ReH7duP4opQHa11jNI2PH47jq16j3bzdWPcaqwter6Ni7zeF
KsMJSOTAPA1kWJZD9ozJfZyZgZBt7eg9Mne0iGGTLmT9KS3Jd1f58thaB8Hne9cp
xH/TWDcWC++/UsLnyRXZJqobmJEl2SaDhqEpxSO1dTDRTwdMopBxWm8VXxCvm/4G
3lKwPjiivrnL6d8iDQx6T7uYIP5Sa315oqLqPbYLZO/yGD5Zee+Dgjx5gGqhZ24k
b5j7f2Ew0tQKTgQ83kvsXaKd3mLp0ziXJoa+6FYp6pHdnTaF2Q5PylBmvudW21T+
b9Rbm/NndZKRjpkcXLQr7ZE0UVyAIDP8UFPLnTkxeMJPqaUDeLrcGibkBRM8+TbD
apFolrh47eSe91n4vlBOvxxFcwQVMQjlu7ZDKa+Eff8hZo95cU430SBe+BnJnrNS
6hPF97nux5KKMGVyJa3l4CDTx7XcVD3uzuww8jeazi5aQ/sYHP+d9TKP5Tb/W0WM
l9nRmHAJwvZ7iXi4lo61jKaqn1sVIEBaleHXi6TVGID491Uj+ehobxu5f6lqmcIi
YTY7buxi+CX1dXLXqY29zM6dFYi3lDk51MvWQ4K2a3snJN1xwbHNYd2Hd+Cziz+0
L7Pu84rS9zmNnQsLioJrL/Hr9YyPtC9jCqSaiiMCpEyeTXcCE7mGKD6vRoIv+uCR
2Gy/0X0DMFGrOFwen0fOsaiBmjUMr4opVpJxjePD6EuIuDiEBCm6pmw4d418MAJ6
dM9rMRtXBkeIwSbIdk9yR2iVuO+pS4tliHQFJAdtKXXQ6D2V9SbZICdo6IhUAHsI
6t1zN5axUWyEDFVpk/KkEdIB5/ZyH5S06k+ruRC9rHxHCYK58kvs9pKFiRRyAE8P
pqgt2XGaWWcz+i1qQLpHPba0hJ/ErJk2orJsct/72l5oKkobG7HgCtax7inS4Qia
K7S7cq6C1b4qPyp3iSSJuvnS+dW/Qe7jjdNV8M5xIeBrZldiMqIfomDYYTBuE6i+
pRwdD14Age8SbK3H/jJQ7eYooGeaIAjO4op1iPZkySKIMbFFXfxSxQkSM05nsuhh
C1sCwviuhs1yDkYFURhfgyhJoWV/NVV//HzVNtLwPUhZNOnrBaw3aLawOqvRaC/O
qJYQlD/NQ1OYyYSYm8HjJx0TvPZBSJ2QJA/oFGGJQ0mT1pNeI2sOESjVIm7gs5qx
yV7OSXYF7Doc8Th1S4UBwmeFfjSYKT+6C2d77d3Nz2+OeB+Mb5x4R4ZxdNWYOemQ
2OiipuSMI+EZtJJjPHyMGxIumK5WjvKhjt8pPcKOgrfXjAypfwigUwK2i7+5kCCc
HDUVr/ktR/yB96pGkEY2BW+tesdqjRdhuSZOrQLwzWarsDpNrGhIqev65d6fcMzl
8R0nsb+SAGlKUIpCcQFYGRcvVNlt7v0o8m7NgmG3Gmln7T0IA+rGUTuRXNJEbKcg
6FsWl7pDjwKMN0XJ2qh0CEOyT883mVe/IUfHS5nW6QrgFMwIu/f6cNUre6sGXLCS
vgUZutA2CndXoFVeJrEwzjFc/5dS/UsSyh27O/ohpuQ0CMd8hnSYY0G3z9NAyZPs
YlRRYehX0c9aZukvqrkfo+tWy0E+Uts7urEKixyrA5x/QIL/h9kbZDLF3c1TGBO9
F2pDtpYy3kqI9zPsY0jl8MXyUPbr55HV5LEvV2G6Ox4HdiDheEUx8PmVGVIQBN12
/6v7/a0j9OMFl7kKffiXl6kSvNG3d9u1CxIwB+RF0HxoRT95NX1H6M+fBRF9i2/K
kvbZQRqHLr5Jhdz1h/aLEG3m7CJDGJMiuyLFVrl24CTRYeKntGpMLcjTk4ZrB89C
eebSqxtlp8c0HM7U/KTo/ymg/4TpRQ4gDWN4cwmbyVF8+VpcRJOLqVq5FY2cHKE/
BZ27AuJatxBkMeWdGaMk0Bs+uL3TyKJMR47m+HKFgnmGTy/wv1YO2w89ZHmJzUSs
3MdI4QK2N5uc2OowjHiyht3asisX+NnxZ27EOh0R2CkRAhyQh3II1BEPYRSW9zGD
cTZpOQEaQyn/rlZLIGAb27Y/MVr15ypdLrfKDdVFzLNXxMVRBN0mztrZ6KoO8C6t
pV98p05TdyrBz+ft5811MPYCIoUj/5pBpk4NKtaCPj9D0DAPGTeeMCokSUlgpIC7
/PobO4OAkSPmsRi5EFPP9lGJKB2ly67rpCL85nKtxjHfwTvJ/0YFX/YK2SOIOYO1
Vs3yXjwebBYbGIeEuaUqSo4bU9AUqXk34FA6TPED4Qn22y3mQCu24i9LNbFQEtXH
xWJ4kRqe0MqsQOFwqezlvEFVWzejexTukreakB17twxH25llNM2u8ykgV0ZWPAue
cROiSZViLaxyqExwk9Mx4LkCh8UFwlGg85qHtlVSDB58yKRE+1sRX7zxjy3kauxJ
Z7g/P/5BSeXh1HLXSWfaj1zM9z707cS5zY48sm0P+LpGpPiMY/3sQ0hnW47CpWkF
7elEHASFT0NThnIrVMwshGhDqpBKBB/oggbSm80bL0BOYy4fteUmz7f06pZZjANx
w0r+0YN2ETQ///InCUfX94L7DlPnZ6Nxcyhe37KHPhtMtdgpphAGSpNoNE2HTAu9
VI8AqRumADePDqUdZ+zSXokgQGpoDPLirbjNj8gdkK64eZs03V2luzQq3XmuEfBF
JgNULOYkThUSmgtvRp+RzPxeoqnVl1RSqIYdH9DAgoMGfu9qMpMxpykwHCzIbK/O
FN1A2JWME7pGm5qELR+oonaEWwgdNzQk6PcPj4DclU86hgIp8whfMNk+tszsp2ui
Tfo4HxWMJrQrbKdhZjErQFCBm/Wbst7l1lxiw3BCvcOKf0buYomRF1O8qmRlUbK9
VxUk8m5HEKq1tshrgqZTc7Lps6qCkV2YjhFUIkB1ZQNOAw02w/uYSXWn4V33xmC+
dxWBKpWd88/x4UTOHZizj8+1bNYcLW7hdads87jstNuvL6ZSJaImmgScd5XwM27B
dvuNeBcCUqlCwkuxh1vC1cjbyVI8YNJAMr43dgiMUn0xVJdiu82moGPT2CWT1bwY
tOhHE7wym1YDP1agFnVt+vGb3WTlKjW5IATR4S6LVieYqryY2mCRrjsgIbjfOK8m
ezS7Ef6mgRnXrNGJHIsL5ZiDGCjKpiFYQpipi6EuAQbcgpj4lkBIGz2qNEZ/cSZM
NhEdzExifCKg8eCxdotz8GiyrHrb/CnzshBEIXCENONnLLQpt95jL7k5fo0N7ShK
7RmxAKOyXL0pZbTsR18fn+4ork6zjv89kvHgs+cnppwJAzSAdXHQzEFYRLv7Y90H
CbjEK4OAoglGQHud2GqP1/6rPyVNcmQIwQVRk9EsPkqUIBuoTGU4Aj2C1rJCel7c
uqYS8etodZF/J0WJKqC8xFn01fTdMXTFvUkcejw2hBF6zHDU6TaYAiie5tEsf8+l
IzTks34EbaGX8pZdwBT6gkofk+/+kAKrIu4Bux/6J9M17A8mfPZvDCiJTrjZEBWm
Wrwe7amHOjV+Qq6N4eRfTAIPM628mtoVEJoslbCUzipT89Ecap43Zn04kRQWHUbi
3i39t9hNkIOooKkuLL2w+ZYClelQYzkXnxJA1qsazgTVNN2R0TIzXwhkM4EXNYs1
Oq9RcyaXcevKhkUQ/N+Z3lb5DCc+Fl/if9KdJFHcj9md1QND64ASQ73UTYmq+Edt
G6sHYkYhoVY9hs5Pxb5ExzWM0cNZds7qwMZCstQiwWqFvae4fFXP0XfQ/aKQZN2M
GD0GKdMeSHTxVfVsE9xnk1eTTTJ0y2HbHk8Tao4OnC/QSJUJBDd1Tz9oudh7DW4z
ybo+dkfRgfErNqKwPDNJuwP3F0bTbYU9Mtt+RkSmgEQgaU2WZoboP7gqC9PPt8yw
1uc+pkahVCB6Y0ANiUgV3Nk3MrPfbXNDmTCVIA/1salN3FUuujf9QjFR7zyG3k4j
1XvBrdy+HlkV6fZ7xqrE8jtNPrXUPYNGb2XSYE9IfyOsE/EhlO6oPcnSM37P7IVg
e8f04OGIz16Fwr7i6wOtP/pbOO5iqSC2L64/t4XBMEPCX1eJQ38R0yfID4P2Wvln
HZYVINis5ZS/hAWkMeUkIhoHRVK+Yu2ifSegpsxmuYMjQqc6Zj9TFyhstQJ85fJA
Ln8SatzFbx+hP0Yh0IFYEKudRzG5OxbiLOva3c6Yex7cba+TFg1fdkLaPFUglwi2
VR6GmDJOGyMEoRzhC6zjKhFh7Rda3byiGWaWUFvFxbAKvhk9DDRk2cTkwms3HoNK
T8M2da7k2LZsBa/cqE/zFAgkgdu0BF5xiqidlS8q2aMM62yZg2ECKOM1GtiVqJP0
kX8Ss13MyOM5F77xHz5bs+c8GDy1Sg174fR+WshQrGjN82RAtt4B/eSrHyTcHaHd
rQYVuIiN06gY9MnxAXjwnc+jbUyl5tWBF6slUkycySLxYrr9YjfL5YKetSn6mDrB
cDyJloY+jzl/nQwbV+7DTaK9ZOpHTpqmXVw5oAIrwLMAI6rLeYxH1N+K/mJwYCMx
29zW69/zMBpsdq0VC1NHn9tHZ4aFaaghGhDiXt6LyJ6EZUiugz7DZgCuTI1EKXBg
lTBrrfW9O7VFSKueJBH9o7xaPe19hntRuPzurOldSqgn9QztZjE+Ju8SJJoo/u/G
NaGgPkaYEmo9h5dfWyMYN+YkfoTXJdwLNMWQRgZNtH05dn1T0DYwVImdP7A3ZSbe
f1Vo/zNPFLIO+KDzTfk2xf27zw7vx5WDRMiwNXOPwOy3/5PylDaEMXrlt7isUwsc
6HepwqhrdbVO+ztpIzQ3sJDnws5ruP41spxTrrijF2Hyrz4OUstIQ1mE44ZDfsAH
MxXaPpaJgtrAnX1CN2MYI41kS1uZWp1FAwCeYDKOyEql6VbQS0laBiuK7WVN5lAW
ml6lzoi4BDHO+3Syw/obEI4ba6DrB+4NxFbgBV8ibyWjAy4ahfy7xs6+0Doj99UH
7eT4B/uw6nscx4sEm5QsEHggQ6C7l3fxu6HBcpzdv9iVWgyG3iAnySp1hQusRBXM
Tmgf1XOM5ud1yFFzwrm+JIrmsPQhaWPFdObQrWz4nSSIfHOXlvkvexCQ5meMUH4K
F6MeylPzNpyPPGgKzWGaRQAsLCE0d58fD8iapFrOG/UBwrfslo9bB0aFqJtbS54D
zxPVYDCtLPksqL62fKSSi6cdiGdHOBrTR8m+CE8JK1+f/1xSP5dfYpECjwHVoR0E
3mRv40tFmB/9F6tvMSYJAhUYcB4QUY29Bmp+mEvJf3xCYTEhxUikPVfFO/Pg2YXC
PnaLA4rcKdbAGyszf7mmmjWn/rAe2MQZ4oK+gH+y7DjnvkC6ib8W5TydCwQaCoPL
Sm9LGt2bpr/nzyli9pzBanvwDFBjEXLHnrDQGz9VVA0WU3wbK7i3+VNPttnECydl
MS6H+Q4kN3UDiMWbIe/WBdKKMUjCr8Wfxd+z1bjyXBP0KvFc+fGIM2/qQzdQSBmR
zdFxcKegNdkplEwT03ICwoyecoh91tzzDfhbROpBib+v+32Cf+OUdzT90+wij04d
VUorCk9F+lAC1xPP/+e3CPYICJddcpizCVB9UkfzcrBOkpw/pDdLOXYPOoWzTL44
mv2QAbf2lGlQpWKbDbga1Osr5q6JzI4Rq4FisHS3lR7MXbaIggVqBh0qmrWfguHS
W4ktXATtJLgkTSZpFMelmAhrPYUXDUlIYj3C9660UGk+91wdjA9Ze8Bu5viDlz9i
1wMNnsqljUgNIneqlmMyoCFgSuX14BrdKD/fNbxRxRUsXXqdPma+29LdADt4cxyp
sBl9kA3zXaaEqzFJgA7BzZp0iH0s/Nz38K+Qn4kMEhUunnOwj7oR6UdPThQrL+wY
ibXz/ay2GQv1l/YDY0b7XhpvDC0zjSik0jm5S4HYhM/6ZwycKut/YYmP+EO8xY49
1GkMLLtQCe2mid7ZRzmxNkBfTFvqgTN63KNUbOCwYY7mWvZ3TTEFhBVfPfEsjhhR
9z0XUmAbGZDt2KrZhR7u+os4FgYeni3JnxoyPbKUCD4db8GXzqm8H6uAnqE+uhc1
91QEvA55gdwm6YUsLFR6cTsPC616xiISy9uheuYYb6DPVOJH4322LcYEgjlfd29S
obL5jBcVALCmyn/XkxJoJ7Dn5nhrVvbP1tEhbQ/kP7gXcEYC5NSJkbDv6dGVXZeZ
5rIqFOrTDilt2MJvKkdPVps6GCwKfa4t2S2PDQjrdr0wz6CCC5WYMrdOoe1mwYzm
p89mlt1KDy6fZsxVLJbaH10HkApHIew0+n2JlC3cLEZ8QDd+ETQ6zl+mkEDGxEmX
lNtfj+jMtEvPd/L0S0CMnjnLaahUTz6K/UwzFWF88UAgDXJwBCk4mjnKEM0/nJ8D
IYYWZdcQOqYvkS/kNaek7hXJvCGbkqn1DgHBmcJwzBPSAZqzxWfemXGC5/1PLYJG
cb4cZKa57HhaTJUD55PdHeXDEN1brlNbr8I398g2MD8reCiMexOCLAW8kS7yVh6r
Z8ayFdS0hfby+ZKZ6z8KQQ5PCg9RzIHvPmobMWQVEnAg0/hYW7uK86KYzP/SZq5W
V07qnXN8+dSUrIdsSJGif/hku1cCN0zTS4roqyAPmxHFe/kfwKquZpdBW5ZVrrtK
j58oQX5fE2mexOaU+XN4mUdUyXWKgQfaUjNtnx6Sj3ODw5ufZI0h2i2ADAY6nBMI
kPG5eaXmoDhFInjaXITCRPa2sibwVV8vR09noJvXKtoQ8kv/Oym1bBkCkwqcmjcq
6pIUqBeYG1zOvpeWJfKS1danu3L6pU27Hbd8ghPBAOnUoIiHw13KjAhOc59zzNDg
t5z7zMs4j3TwGTUVUL2U8JOUNMgxte3LQg/cZRMcm10LUOxfbHv+va3/yiWCM1OU
Yupd61UL1XMM5SoRXp0PEctMYtncXNM/v/hOVfGG1Fdq/7QBeCKrl5/yZcvOdenU
TXDAhmobTcevOanarCvnQtF/88hesUAATRaCZwkJjxWK8SRe4r3leg0ZOdvsBw6L
4MdqhGNAfbYVGj4EFg/WJHalQdSED+qnF6rCsJqlmhY44K4sN+lsPUINtI6eksxh
OEFoUlePjwvtqWpO7IXlFWflkV9sqoqc08q80c4OZBxh2VgkyOeryT7GpRgK0M7i
MsgAMK+SUTUw289DJ8VdUkML63JbbGOw2pjvM60qWzO5Wc/R9OpSKn0kilQLRs5s
D0IErTzV42JPdO7W/Dw/5ZTZtcxFbvv19pBohgr5MMzmMHGffr2FqlYbaG3/IGQM
G6av+D70CaZqXQ0sbz1ngNUfqI5Uzkjre7Y63fIZdmA5L6QHEXlZ5fCpuNS9/QgB
ua6/IYZcCAD2SrR/nP9vvqc/LIqUj1Nx3dMNNNntFVjE6sC8FuxARqqpYy8I5CLU
vFlqD3CuqcqNiNFbhZCWv4SG2cor+Q6LAfS7EK4XfAqHRzbi7PVy39/RzJ8zxjqW
r+9uweg1nRLcOTCINm8Hlr+3VO6g9V9ZP5HrNbN4k4MeXHLAqUGdBxcCivuWZvMO
PURq+kw5UO0GCOFX/roCar5p7GX3Ra1kiE9HPyFXHHmJBf+h4H7qaqpnL39oKWC3
YUdd6CCDIMj/783gOGL/lRpa/s2EvMV6QHQy/IulJfsMOuX1yeSFDT49qRu8OPo+
8RwwW6Whf5OPSeuFCSsrzoBdDZk67MHvl1zT47SrgG3/xkJOpNAfnKJixb0cmRzX
JMdGvtTFZDVYqTNhUTsc3asm74Xv/RmrLcSrt6uypLfOnewx9G2pLwSHbKF+0Iux
Q4H2Lj7GbK3qW45eP4/pY5J7tEyjzy0UNZC44JTzZzRbWddQz0Er256kt8t5I3D3
iuOTItAxzKeH9r2xtrLcvqESyGu13p5vOyhL0Fe5QW6O/iM/O4CuH8Mt+xlOL3aU
mHqsXc90Z1A4mrQJ5j5hNwBAiLtD/vDmP8NtNOceMY3jA1och0E9/fh4oZuV0tvY
4iJthGdfRptN9B/yvqeAbKFXKyp8MhZ5YtkIQipgLjdvTOsaTGFjfGmvvvv2l/TL
s5oax8xc4lnKru0lB9XF4Z+rzY2p2b0hZ0N6gRD+K4RqAuuJmJXAKvhsk4a7b8OD
JkT+jC7+tie978sztNCuy+chN0r/zMAK73h6WrOZRYXcbf2cyKcIGGFYUtFImmTQ
6yBuHNMMYXiBGCoSp322XD+tSHUSBhK4pZMOOXfRXTKPAYTW0AQAuL69QnZLJ9QX
/7XMbh8uvaybcmbaxFlSnrApcuiGO+iG+KEIlnR0NfYN6C2LxB/fYj4k+JfBFpSU
1jfqNydsXWT0CjToG8UntxqFt4zZvwzl1MIoVOwqjddgf/uumfjUWmeo6IHXolmh
FmbvzqX2miXyZHUUymZHSRO8w64+vWU+HSsKQgmiy2Dt4rk0ph8WMbe6PKSAU2QC
8CoMF9oR+JCR0qR0nUe03eX0qtK+ulc+HmHNSdTLEfG5GLtxE30rtYPHUSVSd14C
BxSVui1ewodmp8OSEcrh2tDWEmeN4yKEFIynt/MRPo55XiEB5jYNXsN7ZpXNxsgB
pSzX4KIogt8pWCBr75/+OwPQMaljTN7j8jStzvRcY9ytf/qxo6cbcd2fFRmkwLrz
P1I+kpodqXXpTiBVJrwz2WDLEjtswQALPfatUzHBQpjt8rpbk1/UCcW2icio08Gx
ilGKZVhz6AU3E1Q1lvP0g9mNoAws/SNX+AwDx12Hep5lctUHm9DarfBoMH4+a70G
HoNrNWwKMB6lvjeChz819y5vs7bh7UizD8QbCz13D2vdOLushmyPSPunRlqLE5hV
1O3tb0ToUOkQxldG3WZi3rteQVqkE2WLIi13T5hicudtxJ+x6Vlv1RZip9qOsCDa
awIYRB0cqpCalt27Rlwp+l+IlMEwU6TE08VmOYUYhv7m0WlOgCaqNwQyi5Db63OG
NK0gLxzZQolnjYxo0DycvoUN7iGElcfrWEH+inO/748cr4nLlImfLR5YhNZXu12+
eKjxRqjeOUxCfM561XOIMCQvM3yqKXluln43rTeh3X/9a1NrHrx4DbmoV3m8tZIW
NlOAjAQersrb4WJ3Wy6qXSAOUHewF3iiUvq6GBLegDTp9j2vcgW6Bo7VEfBseora
ola/yCMHxyK2Xg3xCVb0bs8eYXM+N9xKcKO8+JK+PqQuvQgqG1PT3xjb/a6RpeGo
7EDVRxVSR3RbUQe6Qo4VbfQatDhuwL0Oe7u11HJpogjpBgTQ5Nvjo2o3RqP/Hnea
Jk1avsN/c8JuIexUZWETpGh1kz4HYGvea6NFCsONlpi2jKH5taYqokOlydl48te2
ji/djkqH9IL6r70HeWH8YQTXD+Ex5eL3k036+Pe5YDyMqr00ZyNycN4SUIY0Kkhf
jO+TXKW1BA8plLp2DC6LUNVfspnnhpWICGKPP5OAcFpcEYITHkV/vvxMgsRTmm1o
cCXTY7Zn7k6qr8pkRQe1V0U/JQVylkjr/nuxR1dkX1PtamsGYB2c7G1rhy2Fd/H9
sMbCIz93GJsfZLdAgVYsVVIf/XqUyZ8dcR2UxQEsh5xFr0GQkCiMux8kHWzoLT/g
0Spmjysx3sMpNE/vW0TW1RKlRG4j2iRF5WjfH8gXXznTOikxqiu0unHFePTRUAOL
qvhQE+SLJa39tGNTXa6I/JTopCXuTGFsSNO3ROJIRYTp+Scq1lwoeE6/vwXGHsRf
T6So3sYRG86ucvYyESl6+AXeBsKr5KmON2DR3jdbDUYFo3yt3JqRo9tCnYIXe0lB
Eq7h96x7nBAqotvKx1rnyEKcZ2osMrlg10bR3MvEzEjzpchxWP99Pcs2I7sYzl1Z
SLDBTg3f4qizVZXll1pAK7xHLMcYpjpn1SCLrOmWmnm0MEXmeVaLVTTXjgcMuaaF
o9sGSjY8G6xW1pDP6suru94GG75daG1M9qeSCUDFjH1CQ9kgXISseE4JELDlzVkL
9bLnHKKN9cghS6piQaHW0YL3GG8TjxpYn7XwQRpocNlE53ueArGqTL9Yze8tNFKF
Gb0SlhVXMiqFXTIdXWUl+0LSh55TCIzTv7ZFdZGgX9drbSZnRMYyvw8mI3YP9PsY
sfK5gV4GtgIknLcRB5aEBP5VScVLSIMfloMFbeywF7W0qwgS9Td+RtBOicdVQPbn
SMRdM3ozoQJrSuzPqC6w06h/Lb2NOOGnuhM0Em4dhQeWpF1a/RCg7yyBe0wOrRAv
+x3FjCcuUXTIFsdSZj896cPNfoGE0NJfHqI3m3KvmJ8Fwi5gQKfmAowxzWQIgsqz
FrbnreLCqpRqhmO0yz0VKirAvmyRYx+B+98E2nJIpduWYUFu9WszxkFiL89ZyXqK
0FAXPhZgX180fcWXRSFO+CmwxhEgLrlS876MVdxeQjSyZgeP8d8qa4I+KaStNuBi
zrd1ShhmFAULUrxOZhCJuqnZ9hWkyOFCyLw7ufDKiiySfrMMsi4jwkqfE3IXC6Da
tMdEZ5c7XKUiX7K5ZJlQfKpKSrZrJQYwLNra7fR4m0DU7ulGHAoJ3Du86Zzwtpqh
q7OcZrF3MFhHDSo3UT2TKdk8zKPis5/zcQXtOCJxPhNrSTHdkiqCoUsjXECICwXL
I7PKrVfGXKKeuc+tfAh6/azieQ3VCQXuokM3XA4G0tW2XiX6wiZ+HXk8kj6AyzTT
aUFoTCmJjOv1w8KqlZM5vady4i0abmQgp9yQ1JTwnrRE7HPyrmQg+s1dpKeeqerg
Xxh2K8MZtfTZWmvgTBj8P0Q3HY8hOouqrcej11VhSQ/k/HB8omnjKWwqqgoLfjBo
mKWN/6rP7QM/w4GFNRuC9BVD5G0iPnYrwu5JMWYHQvzHruvGLhqWSH1rTbcZo3VM
b7ku7EV3nrFgyvM3fPSqVUFtlbsCFXXcjdxUukiVq2FN0A07a2dZDIw/vTH6jX63
WqzO2jgwzDfg74JGhL67L+onc338km8fAyAl9cqmYG0+3PItEWIvDgO8RlW2gAG6
0CrJCKqOn2JVVkeYDaMvkzTykXG01tZAXzelRTX6HIDjS+Qq5p8WKJ79RtOjfZM0
ATGJZ6n6gaJhhSKRDC5tb5OlLFYLFRQLtjwjNFa5/Szpfyha6yG5tcZQEHdUcw5j
3vWwyablaz1hMTd+Bo3W0zZrvdo7+ZB2wSSd4O7XnYZHGVGxlGknmesJir9FOAOm
L1BCyqcc+s+9rJe+gvJuwpjyu2tyDHejNw3D1JGEQWTTPH4+DrG/BpW2OVJhqGJt
XVpLPmmyyIsgdx/12D8CMNYKaCaEvidWIktvUZCbSqIH52c7HEGtLWilVeJo5odq
596FR4U/uKzbLdlrLwBe3044exhbeD/rvNuetdiQ4ZZliHSmvu1G+/XhUTThax2V
l1lk3OZMKqzElVg/ekcCNNpjhXsJ+uLWrHFlko53AIJZc/6ynvHThbA9cNEGBg9J
P1/8oOLzRy+EFcBIf82X95faSejY1BeDJCPrAtTo+/PU8xE4/VxuPdU7X7eY9scM
0rGEhZYlSSQN6qP5Ax0TbgN0M9ehcoYO19GkBmy8LjUWvsJQvkvrDqGfZsv29rx9
li7mLcUAcqcy5XCCYYlHGdvYSYGc/06qN/MjA5NwV/hP02Zg26dOCrfctfAYG63s
8F8GeKHzPyWq1ucLTaf7v2Xa1FyIdjmiviKR36ETsQ2cpdgbpCAYk+2FWo5ReSRh
xTkQtiSB3BT/lz/JkJK7pv8ydfn8/eFGkbR/3yDs2sMK2YGhbyU7hRiOe5aYcWdG
gJI507eHpTPVyc0IOdCj/G+63RAVancvYPKOWWfgvJPNfl35W6ocN98XAuMEKJUC
dRWPnerKzshQgGBiWnBxUS9p8H3FJ4vS72G/nBafe8TsPloqIvDnzqVJUnKWZBnH
GJT0hgEQF3bFEltRg4DQm9Ql58iNo6aH6McjX1Z5Qvem8Txf3a+MsCXFr27FlDsI
0MXmdARzIq5ir+VUt871CV1yE7zTAMWzQxxh+dL2q7cyIzuPIvJ+OAVGj6j0RjQS
ned25GpcUO8gN+M0t3OdWs9Hy3LRmZq3QrGUx5JU03uj+lgrJihMtmgNy9oF2Bi0
TZWV68jwtd6pcUwvDwmEMXq0DJ+U5d1Zf4SrRCr3UVEa42CA9as7Un6/07p//XCm
Jh/+YX7LdUN1xkuQuwiBZumMent2z6Jv2Ro6N045zWCcW72Kml6jI7T8R+DkVgEl
PHnRYqEJ/g/8as45O0Wy/0Wkg9C+8XZk2K3ErsVKvdGWtn00rANSH2RYR6rCNw64
CaU/nSgyB49otWgYA8KC89bYGteffheCvpLgkpO2VbZmN+lJDinJ0LL6Z5zsskBC
vNXe8b2PdrvOJxlpNkRRlP2cnKtb/l2NeENvOKEwVpe3axU4ZuVij+m4FBS3kTJl
zvhACRNrSV11/nGgyNtk8eU7Gfnk5MmCQhBYCTfM0vTAdgT+tSd4Qi+f7S2SSPf3
bA4I96K9FMpyU6FF0IOqqUwfWBlAFQdYt14u3j2fmvrmFOx+ZVb4Kck6bo1CnRKm
m3OjpYQQkdasc8dUyGWUvrDV7JzjuxGSfBPr+XIlz6JpSeCsLMQ7E1ngdwwa0XUx
WOHFTVUMFJRuT7FSOLlYBPjTUT6EIEiT8c5XGjdPfQMnldCOxGofic2NJtzf75/v
xi3Mz2Ewdz63juerigJ4A7kb/SbevIs3sQLQf1hShncRZuGFraA6o9JQcE1kp9xs
SXZwY6pEnhnFW/54UVm9HzBuikmLD65RCRmiHystzqrYaHbF+MslFKvJFKyjq16e
uBFXY7zW+/rmohWR+lcjkfMzZ/PEOdfBYshD9QoxfoC6xS/ynV8FRRTRLA5xdxOC
gcl6GybmWfNzWMz1BKH1XjnErTX6C9+ehhSLtBuVLtwZTpffeiFYfxydA01VhvMK
MaM2iNsLUEO9u4FdB4MzDm5zr9dyv4G6YQ1uOmi+rg07Yo5/oTyhk/7OAIc/pQYJ
No48IgkUy2XZU0iqikUPlZXEI7xVYOxqK5ftGqbC67Xe1pGzldJw+/vuGLcxp41v
4nuGQRxjcrD7/4sCyiQ2VbKAqy6PAFXwNOJPGgqSNOxz9sYaHKzVH0ibrH4T092W
9BQubUqU/Qz88sgLf0N5N4frD8V/blA4/FFQgPn/Pu5m9i/qB4BmbdoEZgYf0SRX
E1lL5UW/UL1JAWPwPPanYDtBUE7VYQvJdDnTh06ANEyjzKvz4Q64MiDsFsrEEJa9
fK8hDar1gOgNNL+E4xEMg5dKZ4UtDZ5Z2S0vn0/IzK1L5xvntRgbXuFDUjcKHocY
9nYqwUncMqWGt3uwEWZMELkSImBR2VGi6NOlMbOhFOphJtDuLz39+si2ypvjFdTj
fc3FaWtx8gEhANbSGQig4gE73uxPZPRd6RHIDeUHT/xXQ4NBE9fDFDnXlArQ4eX5
NTBPe7qNoEtH21B5L82ETrX3prMcXhaXpwMlNUVzJmtaJlFt/StOwRjNGtbPZOYu
MBtM39gKTteYCxffvLo08LPeOX+1WLm8AZLDZk5v179YQlpESclrfCiRBAzSbCYT
tbJO40vjkZKKyEXIiRaBdmpwYVJs5BQm5GYBfPtBxS+FDU0p5mgz4lsmcJ+9vH1k
Fx0dcAkTjrXOgDxWrPh58mfzvFa+SAQs0qtt2owypEamRw3YGKHT5VFPjHBkZIVu
mF6WMJUnbLSrpNB9WGe15TtvnbkaMKSzS1XXxW/K2P027Tj+GzO3Ugt8uNbrzLV9
Mx2mM00zsJpxgKnR27Dxgi7oC5Ketm6X6Fv4rYQchcIv8wRtSU8VjiDqwf/TbUuX
uFBQ52JcRJ+1tL3MmVuwU9CNM2MZH8EwTLSFb83HjF8ZnCO9rnmY7rVzRZr7PMav
EkZfZjoAhdIo1E5Aqer4zbtoiFQRUsxtV+Vq7jMm9F6S+k2SqRW2MLA5d1iWVRGy
il3usFnwBq3P4N+Rd5HdRTryNbWBmKpHjMmwgkDZivc/PbijlwbClxWXwQED59Ut
rexo6cid/YLEL26qhgdsQ3rN39vtJlYxr980caGQjNHa0yhnk1qMkjICqRfhXrRT
ZFbZ+SidTzrnka2b2Hgy4rbip9Nhit3zaQuVizHjoTi5jFO5KwSEQWH1R74WqCZA
dlWPElsY9XrZ+tDEsZ70WwtGWdhKcEsXlNBiLAwvp7dblhj3free3pv4tqy40SlY
bt440/bbSN+lIUsvWII47vgWIxIjj+F02/yUC0Y21m4xEiJvzWoyzH8d9M6mPjFN
iUx0ehqhQUjPaqBvO5s2tqaW7IwTIkbXbwaED9RcQO3/C+IjwVu4mcbyaGL1hb8d
6ueesXsJMX236VvZUNWHKNTp4Ik/vOZSI3cipOPd1yNib6yneCnk/Q//Ao4oWmS3
/YYk5AwXeAfv+Xa+jawKyUv5sdgLuuCgE0UMBoqZRlZkhfk6wSsyAmjFO9Q1HkY/
jw/jhRV/HLr8LL4APwxn2wZOacjOOZHzwTq/dlzvmCD+A/Qj2YIZru5FQKJEmW+U
JHiab0stX6ih1mtxuZ4y9vT193tcPzI1FnNCFFV5QCnh2pfbCWgS8J3E6oo7FQqL
pmsJF6V6seYlDAY4JxpmmTy9y/TG8vK9VREIW9s7wlWZH82ZE+ljRH5bYyi209jQ
UE955JvBv9nDiP5CuV3O3JQUkkGdaWUCCrQcHDEHEiQBGzjhidEIqMYLhnP54Hj1
/NysVbnEglVmfTd4xm46jQU15+nELM3oSVeDj2Z3Yg9ERhzambOd/xmEW1+GmrLW
kFDYdoHOBER5tFaY27wd8hLuHqog+x02/oxZv/h+s1/vEE1d64m/TkmzX890kmZ+
dsAz0WNQF4HshzG+hfKNWglGw3yvWyi6IFXcSR+TxIFs/PjpxYUqukJiws8n/yaU
VMgMlihlV5pplOa7AM/nRgZVdBWEKGmoUoAt5cL/mJDc0Q7CwuX724IwbYDynhAT
Fz11FDKMeHbK9WOlHVsmic3qcgvFvq5yTcc7+lII0yluDspHMmYf2f6rC1hEEQiV
YkWaMv01+LmxmYtjPb8DgeM2vO9Zrg+pia076tc1Y67cfxmztzqGM7ADlC+Wyz4k
r8R9IewFgs+/IWukK3VN3B07fxjYALymXi4yjKO61tKSjbXFvsWwIrzLjQnz5kJw
cmKEpNZx/6ZDf5sQX2T+ddciw5DCO2JaiErk7ajjrhZeNxHG3oTUkAZg7zUUFEwC
Ni2ij8+CPehgYwEGTjfwx/CMRO/0jFZML+U4tNrS/iMRPF7DGhCBFKeHeHkDISAi
A9UoAm3DqgwMKFrmeu4XlMZxZInA5vvaEbtPfwZ9jgYGIwchzyDa/UXOut/s7MhH
m8oq+46BH7pZTs0WhOUJ73456lPCeXCdxPl2ipq820+d2NP5jlDGrGsqA54zZ5yd
Yhd+g7vFo3QvuYQX+i26DHsS/ANxia2QY1vorpDr70mCkzTw+oxdbOR0aWr0wwCg
EQt5yKnDRKDq0qOjccKKw4XWf2o34urJUAuJ3T7bKEXGSG2yWSJCPkSXimxaRm5j
W1XrU5OiPnouUpZK1eD0Ptmv1IPl32fh16A5vmq4kIZ6S3YS2IhZMWxNggaJYILC
Ol4R2bYNI9FtaA5+G7rql4atIJBZZvkALedX/4kTXIpAaifnaoMeSc+q5X/rj+Z8
skHieBo2kLPZSasrQPidXbT8Foo+3tNW+/IsP4FtSQNZDIhcI8sFylGa2YKEMx2H
qRy8UBIeZCPOPdAt5OqxRV8dv9C0eBMdopF1xQ+qqhQO+HyyL+ZsIIWFw00jtXVP
9ejolDaLGavbgvW1o3++pCWXTMVn0mM3LDfyCUvNUi/A9liypOxZIjAW1wO9brjk
/7w6vS7Zv/fm9aZJimMyEuMXXd3xU2vrIXJ1ZOC0+OeX5yh7FwDIpDHV4H6SwpgH
kjtTmVYnsfyR3IAJT11q8hZ1Ty9HnvSBaBJuFeedaZo0RoyVugoLuK56eZ5AgELt
vcBaRSRiL5/7XUPDP5J6i5GaAO7JLN4UmA6dlZLuCsSuu56RMj0crJvnMrBPwga/
zBhNDrMtvqOYcmj4ugpSWfd+nxWuYGxyHbWNs258xDaGHsuFnLDKLXymrk2znU9e
dCJWLUbBLC9ld0KCWwxoZq2fbXbLdctTbn2RqMoBcLjDNPvh2IoNfNcABeYfOqmJ
CHSxO/yPTVTLs67SgfhcvO9A2S6w7M+ikTzKLX/tm57+1JlG+JpgfMJbzmmiQsUW
xcY4CZUbhNlfXrWWHXG2LqRiwlwy7rtgjJhr4EhPKLU/RxF57vV5hj+qhaXPLNRO
Y8e6T7D4wznk+QosjwWVWHvgytuct84jO0w7fgdWCPocfUXpyJlVwvZ/R5RFbxBq
O3AP0wab6a223F+pWcvu001JqyHIeR3p0+HxYRtG2CIILKImfcjXq6nbdCdlizw3
HD5qbrrfjCmQHl6IK3KqPmW+8aq33FlLQeuYdcynn71VduvuvNXU1h7oslkxT6l3
IkZpmy34DtSYA1gFOF0r4XKz3mCpfmaxvrN8xyASr5v7p6ybP6Lm0wfqvXPIHexL
jGdhuT9GQVSkvJu5ymlt4MOAzEg2qdHLtC2PajdZlNDvZEQZk8IxPUzqOj6lIIq7
W5ATq9ILr+PVRRvsQCI1KJuYSKir85TcLxuO/fUVJdlpxFZ1xK9EdcrUWR8UpY1o
J27QoeTsPpEwvcxxfi0lTf8+kZNhE9otgZdHxfoLSPDAoTZY9OacUXkOw2huFue4
3UhUynHhopsNtFWweWcKnI4IZa+aEztSlNSDTnHvj71/Tf7LOEi8d8ugsGzs9O1U
RIgS9dAYrZNLhaioBy/DM1aTzZtIm9mkQ7FqMrlr5Ayns75vW0YG4TUwVi/axcEk
Jqslq1GWGwYsHcVRjMafbz1IIvMVdE9bilYm4X3wvvhYDjM9FKIfVUnQcWW9N5GK
2hJgffYZ8ORP1Mu8CMfjFtJgAZ+tBoEzU9JC6IfTSc9541XJGrvAcu8rWrfUnc8g
/9MDftH7h4fCjsINBdQ5133++FJ3HIgyj8eMNKtWqBehpsSDX5SHe4OLZHV6uqi2
b4rhrD0QA5hqoRnL7CwYxJT/G+gEy/KvqTxCvG7neRLszrTjNWWJe0wuC2AAzMgU
qCXkRcE/zpd0CStSmTMokof/HpDkqd9YozFLOt6Kz5XbU8cuW8znjSzpcTpWfBRW
u7riCt/KmpJbF1J0S8xCNwlggIb4lvTo8V2I1epHxX4mfNGUcinBOLoFlA9OwpWw
UeD/w3aHPgIUjCG9zpDdQ9Z7bM+TdocOXyyw3PzDyvGXfPme1KcU/jyYNMXEW2W/
uuGtSFdXY+dD69Sesh0BLjb3+6nfMjQa+cvbKJiUIxRX15IIQ/s6uXsp5bXOUh9R
gttU8kpX1M7oC5AA8+qUZvUTZn7yMyYv7f2V4tVERF/h4/5j/AARljUnNyZQeFnx
D445voTJQSWwrKr0lyT1Yx11v6picN+I67LuI8Br4SiLfyznkgWF+plw8q3d9QUD
zAs+Mo6eIgRZ6BgdOADubqzJhB4Q0K6MIAIRmfKSy7DGZvgGeRc2lRDOuB5RM7zY
oV/j4FOHzqHERq0KWOHcBkTvtlWvhb9wLKTt9WErz31kmz7FCq/HqEixOHiXmW2c
ttRVdeQ4diHy/IdMGpyqaIsdfffIpb9rvRnuhJOs831h3K7zDAdiVgLf1y12mWEF
cOxHyAnFAODiyPYEfL+m3om1qXdOYTFPx/gfUR/F0fGvT1d/rPLC5sz/vYrH85c8
t4uhju4QdkHPb/h7gys6gUw1NUO+9WUNITzn0Ue2QIwCQOl7xxdXhoWYKRst+aQ4
oS7qUVrOzxkJsd/3dJyKfvUvj41xHMAE4+6qh9VzPYAC2AHejVSfg8Nl/VKHVkXu
tiV9MR2dUZvcKqaQnraiBeIM+C/rR7dMmh2iVbNA12p49ua0Yx2Otry8ABNmau7A
xUgDVQT+4ky3YA15Z9cjlrQbkEafGtB/WfQ6w0EkhDfgtiA4P5rosyQRt5pwRzZP
JUcpgqEvAkuUFsQQUyLIB1pWisIuYfDPi91kIUrvGsnX3II/k5wvqVukbirJ78O8
3zaifsMPuVEM+oXfDfVGKB+73xDm3kOwT50Y5QRY4HE0PEpOpxxDHecMD2FWmkUp
E9l9/NpxQ5CZlYV46tZPgaJwYtdJ/8GatOrbyuyzrWpspk5vwEWrW32YBXCSvxjc
Id1Hi5T4AOUkvgCd6ZQmhl1C1XEnUwtPsv+JN9t0a9pTuoZW7XGvSj8qtv957M26
n0dmjPwuKQtgfRgJB5tzrAk/hJXhwKdKOEymlahC7ne0yKa95gSuFK6RZYcVKUac
eB9oqOrO+TrenXaVIt7Kv+Tj19Ef19I/KbJHDvxIf/rNX2IxXIU9UYLc2XI9Z4v5
152kLe676VnuqpxghidpfRCGtgXq7jGefde3QocuzM6XR6UQqFpdGBlVj3igDbar
QokCdDhZkoCZ+VqUICdD4nn3eOaoP8waBGasX888VnsLjtrFxC8CDXiT2jGkTBa6
GVccLMEdMfjIaTSGDFtcE0o+mAgiNxkyldcc0YyBzeJ3AtEBFmSaugzfRbZjlYBq
OOd9xeRUUvg2NySfQU/kah1R5vVerCBq8gp/jzwRdghaw7MS/P+ylHIcyDLZQuqM
QAdCQKC0m0T7nfbOg+D6ql6FwQV0Tsly2RcQQf6l79U+2hihmo90yVB4w19V1Ge8
31DHNjFlGhbD+vHGDZvhRUUaPrEK7cbfzRRHbpEK7RaCaqbhoMclY1CPr/LApWx/
2SLWczLht39rlEAbYVUoJp16ZIEeX+ousXKJOIQPb+PJ+TQdTA83nz9xUTTKgN4r
NiW/WA5VIdvIxe9dueRSGfDcgFWcWVQTxI5PnF22DpTlq6IxWkVuroMB2npkZYuT
dpO8dkdrCAIoXwcDFeUl5z1s5StklqyumXRsmLHQNhH5DL0OH3ModfvZsLKxLQiI
Vih69Bkc8qUcRxi9GobfzsSUnHbDdcs94XeBzLNghdg0SJ5of240WpgW3YfElRbd
yenZhVeyMLaMkuF46Y25WN7PKQ4vYsGyguYawWz3qfNNXd5doyXE/CDBZt6ACnPG
KOYo111ZZkYHSVIgr8Zk4gXOvi57FTYCWgD23pFzExBGb+rEh9PYp18TWD//QEU4
Nfu0X2h0zRSz3gNb/4vpDLxQc05Xb7VQoq18Ug6/H04Q7m6e+5wz+mxauGC2U0oI
ZyMMIZtQ0eZpMgFBrDSAEJlX+ti+XpuNqzCLSCoLvt+alVVnVaOTFq3ivfVA8+YH
6vVadeL32pFlfOo78imrUM6jrGEyDSk7S5xapfel5t9HmAk3YBJgNmMC8l7H2Z9J
lLbX+1wxTBcWgtX11GRebeqfMcP39EtDeBlK0BQdHW57NbiavobBs5qMs860ezxt
lpRzPl+RfJ9ePUx3WlDCFQ5F4HtCcVKea7s2fik8NnT41oAeFo3rKMKwhIcpSFo7
jqD0/WuqZDfBUF1I4mz721d+Nxnyw0yIJaDawkfdmRyfth4e2wqvnghkxMGOvi+N
Xls6O4Fpi9d+JcGvXBqdfuhZ4AVeGKzXOSmY3Xx7E9LE5B/fta6W3eiov1PQ66qr
KDNnB632U0xLFFXt2P5PX3yk8fj+zm3w+mSG5drp26T7SOaRO+6MlgK28NhIrvKD
Cye2A2oAMos0D758MMeucj2+VrYdebC7vh8Q8+5Yk6sBTCKLF83MabS5U12QjwRF
8cTjcSTn0GbRsPEnrq/eTpatiGbli8h2i2xamJkfYmCoYGR2QcmK0SEnDJUBJvnx
/s0++RAckIQHibvOQxWj4JKqV6SOzKvxoeAzHU+CKlRocthu3Tx8bps72Pxr2aJp
wItcFf8RpJO8svNTXegLQ9944MbDiIdoHNHLg6IHu/jXS1gizU8vkuvzEKJ1ditd
pRaTHasBCOOZe4wPWL3qTQjagL0XQreWSaaI/hcK3BTixDpjvbS531jYhv70PPLC
DAPHqNeLjmKtArF9IveK6AaJ8YMETD8kdGG02EwXK0wamh1nTRB2Jd0LFGXxOaOO
9K3S5GLwM8zYWR7jpEXCn9hbKuKJR8lfoOCVS62NJmgGqBO2NC6IeTAbf0i9qo3u
vrJnUlrFNU+U8xF2kj7gITNpYBkSlqPMOn66orZXNLHlDVOfvHwFnKOfUj1GZLLP
IVCq0lTWMtkiBwikjhm+6qvxOcfZVvGIya3fs6Xlea+EmxESXfjtU7MCQ/EtFsBk
uHiGxLkjMudOFBGc7+Y+wBIIl1dOG9d5VkDJ3+QIQOKqcwP1MU1EoIIMPm44kl/X
BZ8pVygCnR03p8UDgfNn4Em32UzPaRhPeRkTowjc8HfwCCi1i+7LeX6mEXq2kX5r
t0qSLaSsGeC8P0Z77wL/dLHaobT+DAVQpfo9YTDPkx1kM3aK5XrgrkEe7WYYb6+7
ez3vWSP/FyZAhIK1joiLOsE//v8BW1k1n5A5WjxMRaoJulwfWx3MG47GGgHXRyLy
HQuGv+KRlv9EygB+Vzrbfc/hRHQO9LINHKXoW8n/+qD6wyxvVzq9PrKVHU/pR30G
gZGfhJYCTj0XDqL+HhdxSku3G8Z55RAHhfW8sjJpPSeo3H5R2al/6D+sAxKxRL4y
MW/XR0cHyOmJ1lGhcZS0UUDz/3lEwvnmnAcQoegb/rtVqgWDlFuvaXAWAV4WxAwQ
AJmvmr5xXPVnVs9sbr3totfjf7j2Yp1aEQLMqRY6Zae3fYmye9Z4GMTJPHb913xJ
bjHytAHvO9VQ6ZaWBqZS4+4txzC/QWbms4k6qixFyR7PJQv0/gkxzLmBs1QdAtRK
7Q+eOHLxaCTcBuKtOtw7rud8W25FTEtKD71qh9qJrF8boCRzfZHjG3RVtI4XqwZJ
K/7qwrydvHS6ITH+K5WNH+LBEVeGgUfF4SLPUcWcQw5NPArumo7M6+BAp4pvcysD
uJf4Ny6BtsFGb2jcsGPR+cAt5+n14necxZPxadMZEF2sSXUNoV0jRt53G1bh2GFT
IU/A3aTTBmnxAuGtimbc5GurlaCod1jv41oJWvPNKaFaZWi28koJ4BXSTYpozQMp
ogHGQ82E7xbuupQAX+tRU41tnjaYY4Yhg2maO/w3YtHdatyYu9lsxmQeIeNCPa3N
spwm0rSzeu21S/fyi7VsniIwXJdhzPg335Dko48qXEwy0645DcjrnuoYFxNngVbg
rT0A0maq0bWVY0rwkvKInL9IHKVAZTdoF3HisnSaT6yAxz4G0CN9b2VF/V/Pvtts
VBbtS+7o7vUky848AJKjA4UqK+hktEDN4W9iJQuPkWSls9H9A87CmbABPaU+zlpt
9zQbCYjglChCjNfroT6FeTDl09wMDMalog1fAq2+D0dTvBE0exEQoyYjJ7mf7q2q
4PB3B/XTY59xMXjrycD3ZxfiuOFBRJ+gRdvpboJqybxx+8nvJLlxR9waEV/ww/Nq
2EKkPxKcWZxBtGrQdKFgPkOoSjZJr6ji99lWA0J3Svm7Dwl7RkajBi+jbHKE6N0P
jkDV9cLh6rDoAKNxztbcpbsgbO4p3GfU+2Z3WY03w//5y6cQR/GvtilsenfQmwQ7
/T5QV9Gt9NxLQcURq5x+WlB++MKVKbb5eVxLDZ+/1SQRtJsEqqIMvZ8a8JLY+pPi
AAh+YH/V9nCXBwImXcmpcKOOV2T4oB3KAODjUdjjGkOVzCRkNGDqRevvHAaH4Tbo
gjIUg6/AcO23S9Jrg9ZKNhAAaaL2fvnf0dcME5BqdUv90s8x/NUTVvYP7KYhzIF1
JIc6/aXDzyUIZX77hqNJ07d2o4EcCgDBmobKwIBAWtiI1RRxQAkZSbjTO4zwHwEo
ZG2YqJbpzpDi6Y+OVTx6HjiCsFc37VPVvvRrtYEXbSRUeYfYK87apFCn/W282DHr
j/5P9Q+F+BLeALofFjF2Cqfm3w0ycm9Zy+oWdCc1HJOw+85TaiviWTweJHRXR9Z7
sVy6kYaqAtVVErGav9RQCxnvHI7223YrDyPm9KYkazYEUQI9x3IkiTPDbdd0jpmW
2Yp41dl2p1Sw7owpM+/S1jGTdAkPlt0FiJqgu1NioLmYdQgLPvu8nMgm6ETCcj+/
S7494HJM9YSlh8x3h/Mukwv/nRJoqm9Sc/JDG5eG4elLFnYx6Dwvw3GcCbiiX2PU
fDkat3hbYMiz5w6K5wqdH1lA8+nacpTfg58FNdabABwQKhWb7ja3mpuJlNKQvjmf
OruB4eCn+QrYVJcr7TTz9jmvfswI9BC0jeil/48vEENAaY653zXMWxGZ8k9WNSTt
BYUd/dQbTi9ZVNgNPUwUoEkMbW8Vr6NgUfcJDgVQwXJcPJtsnPduh+RtkIPipHl9
5PJhyOxdw6BjRsr13K+3uJ9S6K63SnBzKOqAKjarekqYI4HoArp3OWbT2RDW88u5
Ly1932TULD+Q38FqTUhKYR9zHgnYRmQ1k3DNVFfVAAcsrDBJzzln9PkUJbEVhPeD
icE+QVS5W6g4dm2a76WiAFKS103dIK/acGyzYKkywUk97fdHDEh15F5qbuY940s5
d771rywPHwKYTKMICE5VPzumOM8F+7HK0u2zCgT2AKxsJokNY2QXsGaG+GOp7v3D
ZWCLCJHWAkXu5XKcDeC6EuqHFoHfryKWlaAUvy6TenREtqQfzqsoxLw864y6ezzt
ARUVXHIa8EZbZu38VznbYzghgdJDsy2tZGB4wD1TfaynYslTEj+WRRRkyF/57jS/
uGdeJ5TzwMmLV0aJb5Vv0UgrszdmSSXECDL8vnE+SAeIb1mLoYiqWZWkZzT9jUf1
TDxikV4fey66pqXqWqogYQEr0E73iMJFREuoX1wtsMwPy7nGLBcHj1oFKiVrby9M
JYf2uA9Aq2acHscrAi3cnECOD0FgnhUxfLUlJRjuRAAPpyV2+zHAbUt2j6QETzbT
C07t1kQCCHA58v1odmTlwt74KMk3suqqOckwPRncGEwfBWWHRWQLz2cL9c30YMVa
C0XT8p3za70Df0nGTMxvL8Kpq84hWBCc9bfb9q/hurMlqL/ei0uswqSXKgISkmDP
tbttYA44FyM66HqTKy9KbknNrY5CJDhohXz3bqvq2m8R/5/KmIBR8U5p3OLQkQaa
E6rys4VDUakrPbo/nQ28jdX0HNHarHAI2fcPamftbbVerD6E2D+Z2TLfJ4J2i4f+
c+jy3qHm9VPQSA6DM7Y+s07o+TrRv7wBaLNpjMMLfXJAmM0hVifhY2hPZebgOYbI
evQUZXmfl6lGCUpewh4GArTrkAgwjE8y+DbekV4rRKyKrHrwyybg+dQaa4Rd47K1
r72JyYdgOVHCW34tzUIbqtGizayUhTgzibTwXA7Utrh7jCBG2xtVoPea168FWIo4
vrlToOifecautu+WZMT4vPeMWmrboz1kvAWqQzQXd/Zhw+l8bbd0k9wq9LGhQ+Jb
0GeziyFULd1vya6JHcIssnE+m8O/L3QF/lJz2y15MbSGtDzwWGas8x6BLtXaEi8A
sujyFhavuyY6fqo31g5fpFSWUH3NzMOn+kannKkFB+U4PdWRpfUVd4txafL7NBfB
lgFYrfO5Yq1j8L70W0FrYXnlHniNzuk4uBxQ+QbUVlf6NehJoYVQHSKmoieR6rNc
cE2M2tOwn6WILsbfQAeA40VWE9gyeRRTuNkWgsfkqUoDM5KxioUGDKyjwnwyKinT
4zeKUEe0g7Lq3TdbR3w9Vz6d4KwSOq+7mFf3xWPaou4JwvWF6J/aODuNCDTPEAHw
ZGqZszxtDGwlFxc2rjR6+OUlZ/4msPQ5GCXtQoxYe8QWZRWM+GYmUBV2P6xXdTUO
mon30f013vPrSlQgOHaV4Hhix5ZOby7sV4wOCwDBosrkeciEpMyKhAu8oaUWzyUZ
RfRhIzVnTrZzMSw6K2I1QhAHhJPvIS15zUt90ME98VF+hHLvLmbUsiG2zkjSi/fs
JwqzTsVbp6Q7SPygjwVRNPeBGJF3gRci2HT02pLSZRl9Ox4sbd6eme+gmvzs51GI
7T3KrNgD8NN6f/6JeVSi/L6gYby8b5117Ze+RMFF/hR/Ir8He1g5bmasdELTG83K
1DlpHFV6yDy3a1Xe9rgS6etQBSNaI37AkBcZh3UjJ01wD7im4G8xKFSokwUpTwJv
f4k+kTZTATqVWjJsiK5a7WN8lBXuTSuIQW3ajtmHTu8e7SDbu6pr0Ueh8nFoEZ6k
5rj7rYMM2c3CFmuqThKTPXHv16uvb/gd1Zqnvc9O+GrYRLaDn716x0YAe7s5wU8L
BzsuVIO5svOVNA2T4V3+TOu3R/aFijI6sAKMzb9wOQQRkbUlnUgf5Bc2ahlIm//+
8yhsIAwoCj3mIfVWg+OQ/yc7BOEaQCZR85kaPnoAgoNXEBhe9ETUXQodlmtKl1nD
/I2h80d9mz+6S1icSb1ckxBP5vpecKqEvlnjLhrpd3SbJs+uqfNs1i5LTwltMgJj
bl6tfbBBYWnlosoKWDsUjv/UqreXqB6/57yyOciwglHaeUh6E5gz4d42S2Orj+AV
HRsJrtamI0Te/Offm6xe0r5X9f+dYb+K5ete3M06DGxC+OzRpUXga5bvwSHA7466
S9IdUZ9V47j7+9AGAy82N8HL2oVQde7LDLWmgkYLWpILswp4bAXWHsIXhNONHqOP
w5l4ssQ+Z5xUWDDzv5+U0uL6jVgkHIQWCQwnS+ih3s0Pk7PuP+kkCyQVnwlhd3II
LCHLtw/GwoMSZvot7jnNhhitomldM6b6HWZAKI4i7qBn8j4tvfCG7mA/0uBAbXDU
hwi/hWiV2bqzOeExS1NHlKBfDONwHexakfVgG/HLCTGFdv0hFqQWdHwsLjsiJ5aj
K3YxKfU2pcIazury7THuv02L3rfg70R+zuXa4FVYG9YHDA/kA+4ov1ASm9kXX7wB
WCm0SPpisoLuB96pGFke0HFqJG48M/OgUeX7qhjZ97O6/LiUlm+h6N4vfeY7Swj+
CuIYlMGPmZvBTFHRFT9ha0/UPQqazr2aXoX5ouHmBHPEcg+rUhC8pw3PxlKIy2jk
GaakH6ll9VscvhZk4MPQlZ/3ifw6Y7q26ccUv4K65bnVGiYIZt3AfKsji2dacajk
GMwxHBCgceDkQDzzqgtl8AZBxiQEeuWeZfyUhBt4yA2xexfx3dB+dXWZZV7p8TIM
c+gZVyV0YWzsulo7Iy9AytgJxXqKbasmWS+0nzdPIhrP1y8uZRZHnEt5JmAOt+4I
KNZYm8Bl4Y16P8fi3aKN/bwZEGVEXU9Jar3EU25P4o3A4Pcqu9GdUtEzVpWa/9RJ
GvIiXPkKTq39liAdEkMfF6uu33+2YCy/Y73c5WD0xOXtu1GCoj0s9z+tsp6kG/7n
g0vrNngS0cGKoDOGOqEUzW3ciRzHgZMz6tH10tmRJQsZihz6XZgpbVkwmRbBS672
fVQAu/x6yhJi+HtaTLWZ3L/1prVB9ndVKogSii7qQhXXc4tOXbxIEgn3xhwAvTbN
UN0jzcA3d9xJoUe6XFEjtVtIJsAR9ncDlsAgrMPYURBuw9GOm3qYK7RKm7nwmAz3
j5KLh8oW2g5VgAcCprHbY917u6epY2IT5ymr383363UsWbrb5MtBLZ0ue5vcEuIG
5gpG40KO5CfyiXlu5JrX+yVswt3ELJUgOPR3l4s5xDLbM6HM5TyHdL8yOihTmI7G
FynEksNlHcvPYQkhYFd/K7L75xhTYsZ7phx2qYCcl1wTiJA6EAsRNQ3JpnMRM92c
YbzG8To3R977886ETpyOVdL1tXC23htww/pd7CBJNTtTg6OIw8DbYLDOx01G85FT
fyYrfkn7UM2/HEZa6Q0aRCYlYCS2j4BRYgzfH0BOWN1UtogDUwfLpTfhDpfk7s6N
cwD6k7mzLgwt3iPf/bA3OpwyDFmU3ovyH9xCzV0JTTfxNP+6M3r/83aYzq3LtAKw
fgKusybdyeS1YFB5LZkgjZzM9oCzUT7uuCxdQzzJ3WQhIXV+SXbhYFssWiYPxvaL
SiNzWtOkJFdogZ14HVZyH6ui/Id760Dyu/2lrZ8CsaLg1Yd17cUPJVRJd17iiRcB
gVJPB8sRnwLoL4q4jueJGOUimyCAHWU+PGusKxVhizvwDKJx86P03E8Yd8fXe1Qa
2azExxflw5Fkkvv0JFrMMwk2BpqXuGmKXwXmfn5KvBnfcF4Rn9vva4h8rYXnf7rE
nmTu6TTd6cll0uZExEn9WpnxL8bQf/Bk5BNW+bNVGrZrYSZReNiKeN4DCP6xY9lP
98QkfmjgkO/gYZfLH67IXQRT0EJH8XS/LBDQ4UJo2/ywQZofZzC7U49HGwY4LVba
dXmv2pvZLM1Us6bwU24mcswdFPyVS6OAGxr0KjqDVzlnbgdBBW3r8k5FGahtWzAi
Ts5IYsyzSUgxJENjBXwi4+B+I3N6qgdgaG6OFuOinCfRXywh4cJNfSBAPaU/u1i9
urOvaWahTNQqjuWFDC1NRBFtKD4/ZCh/ciasMKTh6fqJxce5Nfj5xePbyRMj5lYP
ekxGxJMRtsSa8Vv4Gi9l1xwJlmDmXFbm990d3hTrreagR5sMlx6JD6A7S8deKVQp
Kmm3NDkN08ubo2lHIoYsLdsotnZhdtM4im2853rsstaxSc6CpNT2NtF8dnx/U0Dz
cV/UJMFW0FvNuYbOy5Sj6gt4tY+Noc0n/n9AJlE57xm1dRzCUh1MsOCaaAWHhy5W
9jV5wE6S4FiRUEfIiAmerlbzTboTBn5rllD/bcz0j6GhNzcAxRDGq/QSpFQC/O+H
D10uABbD1pWg8oo4HeM/xCRKQfO9YNzKvcLRiyQ236b3b9Ngeko+/zes6T6YutEc
PIj0ClsFD5DOVpEuMC0nkZ4hmxZVKRv0dwfEGBGj8ry183X95TzBpPfnv7hbHjGF
vJMW6ofONXntGPz/RaONiCj8dPka43hy5sZs0jGbUm4N8Lc8m+9eCvnN7z87aPQa
4ThX+iAMzgg8VsS9MF2TchckOBvVntFhfyblebMc2rPyUtHe8ZDxqBXsIXQgl7d6
3ByMhLygfBDEqYd7EVFh0rR351YCA3MFdTtSDXfR0OoDvjgnF4GIiEYq6YQs/04G
Hs4cN8g+UGQRxiEse+zjfdHgBDHkM3hpi2DyR0p2jNfATzuyQMvqrfOPOust89+R
JN/qdbsM04lec142UhgicdC12Z+8Y6Vz9r57iGllWdmqFoUP33mIniEj4ZcO3OTR
unbOUR9lrCHW3gfa/BbhSYrMr1mEhJQp2QlUVrqSmpzMH1wg5EzwEz0kQRrsGJYS
IWzdf3Lku4U6suncySA48NGpYAL0jpJb/J+7QcoBMl8w0JtRtWxmUrX24FtnRx4d
+FKayw/XO+SSKNYJk3HHjAdsjrfdtdTIh+IBswsUGa878Phg/vCy3SPO/iijr3/q
RuHTdxFsUcT9xf2snnS1dBZbBslDiQeJ2M1XcYgK546WqHUkO0EPRgr8K3mf7IsC
teuM51O9Y15eesY2QdZkJgkuJU9I50cfDeYGf6Z1KHIRxQmEwHEf+ZAFVw3PzLqG
xKVn2j8h4IagLXb/A+cn9r/QBlbksZC4wnwjGkzaJgov4LxyHZzNY8TKobc2IzS0
tV3yYjXxPuebrG5qSrMp5AT7Lh0r2oN7x7FbeQyJbs8x7Fzg6gYr20aumLWM6i+J
swkvMvu/rNpAPSCFQfzRZC2/VaYgXg1hykH96/AHT/K1Eh1nAgW2jj6BeYxXnuZk
J2v1ezIvEZl8mKQMO/MWCvQEBxXFigy1k/qzKGyFGWylpo0OEtlTm0yNy9EyJHRK
YeRYuKM7e+nEu9fJPDujvvZ3OU8xJ0a7QQpyUoNXGLkQ5m7o+BRZLbF3UE0hPSAF
J6cRQJR2Db0LXaCzUwJzCfgjOh7LGjMqc7e34wHGgamXLQeIRr4BWzxn/C7VlJe+
j/nQQl28n4CeR+zq4m49HQ8QR7LBRwVFBeOvayFBQfflpj4W7MlOKR+JnyqTTypp
Y8lEPKHF4tgJIqRl5CQBIKJ0FGBCRp0kEghJK3HQ8NRhJVpspypTlqzROcp4CLav
rDMyFCLZBeCx9ETPNC1IcoAD16DcblrqXKoZX5SdJVwJSu2GgzfwmCT06achelZw
FOb15bYe1CcnqIYnlSiH9Ua42FROxS9QLwmUF6HuqP/g7xyoPFjrrOpDrbe7oLLM
AJhX0croOZe6fb+SWGINQslbFvhe1z4zeuKf2SrjJhiUhlSZZjOUZdJv63xuVTy+
zEoQ4AN1p9kNWA6E2qFvi3of9QyzNboibJYvJl250XdPlbui0Pk2w2JFfjXTjKAm
ZH/JiF7mVKMNkSbdNPoyW7SvcsW2Oa8TV5kczJHC8v8k98IBmAg+adjHShGWDqZ1
0D/T8DPl2pYVRN+No4bOwDS5IpNI82gsptW5mr/GGE2Md7wKQXnwTSwvKLR5/k9W
TlKP4ibS9yJHE545mLoOUZ1Hpm9+pY48xe0441JSCx2qhBqjqwXPK8dMgoE3tuMn
nht3UglNaa6ESc+w/jCaHn9w1DOq4jCesg3qF5uFqdHd4opfT17xZJed6iSsIZeb
UoQXam5YhcLp2OumQ/nqGP6ZzpHlfipLTmWLRNco694iiko48sHgQquQxWEDqIgi
428e3gKtbSqmBBp1HQL1B0bOQIGTjvnHG2oFW8Lk+Y4MshfZczk+fdg9M/ZWGvw2
XGJU6GXITrfQvRMkh5zaVjLZbggNY55gdFW4vBVNapzc44LzQuQ6QACvSoLUfaY9
4IsD79FoEKXQFdCwTTSiAxs4dC14Rm2BrJNVLjxDyvvlxWfi1x5GeDsYZa4rBjRy
xx8RtAmmwSixaYs0jHXKVr0XaKi2+LkCK8yntmfQsD/zMz7jaEOY0FrTlBNFAPQL
pLYmA8N1/sH2PJRS4Jfj0L67cBnxI7/cBezDx2pS3D/lfO/mYPCm/B0Pr8kU2qKp
J9zFhAjRri/ceq3INh150XfMzSryKl4BkIyFHmIGzUwnA8mdNb41S/OtR5w+0ZB/
Z4WO1z6/jRYhS/KiHzcqBo5x8aIGlI1qj6XDJADoqgGVBEgu7p7pCQaCoN9dtG34
pYuW0LKIgpL5ANA4ongCEt+YtHZfWXgFeOia/KkCA+dhXfpAJrRllx5TaO+HOX4u
Kuzai5vkXVAx0OnbqP5jhEyUfmRGwXuk36kIL62lYyMzq3/QfRMkXosITyoym8Yb
Qx/1GOHTiPZwILT2bHpiLWFTCDJ9aGszha6J7gY+jb22F0mCooJk1yBZceQ/4d/a
38HA7u++rvW2rJbGJdaELlF3t2R7rv5pxIGqA4Qsn+U3RFoN/9oFU+zmlC1zAI1+
HpXYuFMgItqKfb4eJmvD/mRFnypadhCPTJ5kiZ1bDnKMLqJCxCiGwAMNEKNKtlK7
3Vm7tDchG7lo9xJn3VsQx3YpyWs5nSPBdSc8VsPvPFVHcpKUxuCmbVzUt+9Qe56D
FNglCRT0mHzPbJeiJGhkYDW5goEqb7pt5rIgTAu0kboQV5OHoC4U+yFjcC9hd8JX
iwju93TLabTvKT4hrblnaqa4+R1wBEOnPlG8uP5gOG5ZVkIdK9TCjbOPgsVoHVLS
WkjHXfmJeIa1SXGLCI37+jvnsL6MJSQb4QZKPoKrspbvP9GXzaeR8ngPOBrijMfD
3LJpWj2ok0BRARxIG0IBaOGs3cWYg7Sa9X9u/psazzurAik1bRutlzDeL1h8src3
pDqqk/JmZui9rR9GCN5mRs/M/EMvjPGR86Bx7lkr0p6BIZ8aEP5A28gLJ10jEC7z
g2IHM1T9zu8f7gs0GBiuxIaY3XgIKZq6Rk52HYiktIjooS0LbaJ3rDblBUTtPQxn
eIzFNpdCVLOdtcM1ir1opJG1AD2y8KUMRYkftmgEaWxyJppoRPWA7K2wx8KTRbdu
xECCPon8dMMjacnvQVrGYi8Oqlq8WoeX2n9fKG9b++bJwJsd1Gcd9R0gLuNIc72j
IeePyIrEFqWXaQxKdGcz9MBbZuSu1LweNaAIi8O3YIvVc8WCOgaRHVFeYUiiXmei
vDZDpPjHRpxthPstb4M84hpcYXsFy4XH5spxcNCFXutOirUCKi1Z2aPYN1yPbvS5
AtDD0s6d1oIn/Qa8PkUuOECXE8KYcpvS/Fdo/1V38nq/jwpQ8ChQWswxJFZ0QyRs
wrSDYnfXlrnjctha0NBbdLrB2TXxnb8jzCMSKXaHE28iBz3gXnjqIJnTGotCoTSa
7foK2YguwZwcLPeDwiDnhBf/soOd1aIlHQ5mw0lzoTwt6E5O2dzfEnPLztgUNlUm
+UNoGImiBe/WgZrhDuVJ7bu/z40dexuYkwBRjTGgRWkf78OZqh+XGqco9YQTSxIr
Y/7J+GbPiOHHHI4Wbo2IAKNfTG4Koaa3Cfgn55AkiobQXGhyLffHYhPmmh6hI7aw
S+SNdhQe5lGtPikpXdv/NQ6yXAjRMQ4qpBZc+kPHL+0bqlU9Qpm0WJ3G3tUPJG/s
EP7owUllH+DzBJf/t2fH5fbOuuZ6Sg1T0ygwLZbPUvzjxly1kHR/XUtkUJz0gij1
u9LilPoxpBYrB+OyMuOde4zVVxl4Zk477aOsxF3JO7FSgVzjgC9N318c9NiaIg/N
zAUAGvzbBMvxrOpDOhITM03Ok/WWy86ElRZzjYEipY1KXxNTRMENsnFVFLcX9QYN
ZXqvJG/xLoikavG/ZQPgYdLYeYkKBxHxcDTX6P5j6/01Vav7ESkFghzhWBbM3uTc
OpuNe7yoV3/sAIt4difR9sO9qoNdn8uWX25+vRxmBQDcpQQ6Qzal+FjV7Js9SMIh
IZWOqFOReKeASzpwidRCD+3/+WEZIrdrRhkhTAWXwSYU+ogLffnLGvDLe2yLsdZt
uxJc80sW9Ui3Noq9jezIlUpJiu1NcTZPURmNUUM3PhLH4DH5sHVu4YXjcPBBQK+t
bg6b++hr83+THZ7FGgJ3tgfZPrmXjpzfn8kdUG4iX5jkcx2Qdafih1t1VBIwqQcp
Mn/2qD8MFURcIMDPgcNY4WNjRFR/teutOTDwm4AN7YgKEOkUQMn4Ai78vxIuhHma
X+pPZ+OheDLABorMWxXPyNz9QS/lNzs1hofVvgdfJZrWF02x3Mx0qHHlL9zTXzFX
akOwCndsyjNCk1B1fC/fvw16UvsVC6f/B4KPjeJFNlYVThk+0DWinEMvloJmEjVw
BKP8DRlyoKRVg8J9P1vmJBCI1EI29Qpns+QG9LgBgL/KjGau3+bgROXvL5RFB+EV
Z8SCTDT/K45kuL61JC42UN+2QxBMABFuH/vcLjAGs2E=
`pragma protect end_protected
