// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PaBFK64q1p0VMs+5F4HdFwNv4+DfPjfeWpB/GauCAq5QoiByH/qkdf4g4UGwEVUW
PN48cP/eV8mn2UbW2rCbxqKoGus1uI8YBlaEyzbW9r7vNY1Y55s1+6sx8vzKVTBi
8wEjSawzavB8+mANWIFaYA71qa9srhwuXkKKifLes5o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26400)
kGTdJZpFSpm/RN8+aSZ6XJ09SKvVf9cE7+sowUN0jFJ9zSSjUlL11yL9DneTRDq8
GF51MP8TF75CnKEkugHTepTuqw0S3RxpJgb3YW+w7hMbc+czjVioCo1Odq0D3Lcz
wno/2/kaoV0d3O4Pu0g4OGNja5oKdGwwiTtp8e2W1/++fC3aq11XkclBdQD5l7Kv
UnXsWimVDt8TYzWN+zq37JGe9L1OenKx0XaeDOiAFUs1+3gwZK16YJs0zN9XzVy2
lGzVGrmZaFIe7vWS36zKYG2p+D5D5Lh+2UQIHEpXTgRvB2XxbVE26pwuzJFGL6hY
ihiJzcOg3FVS1I1Hlx6yTJ+CAMHtpnM4fbxQgGzibWC+dwbGvbT7vgmDV7VQK0To
zVpgU9yKYscVDO0WVD7pw2Q4evvHGkf7iQqVhmMTzaZrfqPSbXXNApgFRIG9yFlt
P/mHXQtcsCbayLZNQaZyjBoIjeIZuGkTyMC6VphB0CxAJymQ8dBR4TSalIUBDmX9
TiK4lup4CDMWxh9KdbhAbozB90IwOB8FxQTLDnfHcJSP0/XueM+MTi3GFxNqHc7/
WZ5xagrlh3VqAco8ElBpSf4b2VeYTBhvjnHg8pYwxL3ty5A4eDeUhocv47p3xbzs
hrfZEtqNGBhmPZxdLqZth2OH1EJfdjFVe4hFSkAowXTlJia3H+BKDyeVioF+ajcv
a3onvj9tzyndZBVkSIsIiQynQFM4wBOLvIjMOoRFpL5q9yXPXN7kRzNQZzNOTeir
DIx1ZYBDpsKEdHrrtqTQCGUl1OYhdnlt5p9hhNpylc1ntDwS4hqbiNPUpVVPF790
C4+46E8EJk/G3m1X/qWLdk109l4OE9xt00VjlLJX3guL+Ks1A6ytFZkAubXkSbvR
TMqQeu0u6tU5ydw1ozgmSA7wfbItzOfMgvtN6vGREX0Sbtg7E584Ot19zhlFsT+u
E/DYmFd7n7v0k47N5B9LhSqsxMSRGgo4n4WDeGtTWWZZNJVVscDF+CSc/wHIwTFw
6VijH/ud1BhW/0Vyfy8N72//LKvMggoLWM68RMebXNn8cQCKYLxYrC6Lr0yEq9H9
lVfREwqlIHLz9E3vRyQQrO+ZhhLWnkW3m0DOKxmjbf+iDoWF7IKtyCBu+Gjn5/61
Ymq4p4fzhE80LK3oEfMLiuptoRhGn1EB9aJ37jJkCOsu30UFxaDRxFt8NKWqrIo/
s6dANeDNK54eDpPe1ZHHmp5n7CjvfnrTr01S/0nolQ175qR++g+NkVgnlbaqX1lp
qm/nvPosR2akwXDlmyRl0JfY7HtdHAsG2GrQnrGQ8DUQoPHkMQiRnMRVobCRN6DR
vSFcTSo5wID6/FT00OChBGSDGOoCi0dqsx0rVAolJ8VRvK8jIuu5lk0UoYD1k0Cw
Bw6zU0OPF6mCdMXDNlw5s0l4IYcAeDTjdVRraRjRDmjPe3Ct2L5rd0PIVrmAzVde
N4jrcDWTdQpaYMl+ov3c0dvZmHh0pCwxzlkrA03NJtjpGLE3SYw/7XMy2aGirBOh
yn5QCNYitjUXjQjJjiXEfnumCBWxfz3lAN48w+AIoZVAS6ZfEF+fTbbTeXQe0jKb
pnDBRiCoippGRIK8LoHfZhI/GTRHoZu8hTAqvxFyh3cFrtm7WWT/I4gVYdNjzzv3
M0h1HMnh/kEMffdpvc/JFa8frXMzUiOpCP+NQNxMot7EVXTQk3VKOdCvMVbKnOld
1rGxECP/Ixp8RC/kM/CzcrmUerod8O0pliR08m6+HLP/VcllQTpLQt7XhDjtwu+5
b28VJ0qw9F2wpEckglt94WL1RFWJONfrI6KZnDgmbwn8VHewkKpcVCWr9h7oFRyv
g4lIUM89F2cyU88HBiRWJXdiiYkW/MA8H6X/EZWSaJridPxe+nNr3nRswWDE6bF0
iZzMDthmCdeHU+wMWwKjT6KpPmDIdnfMoh1yZIXhNfKoSONqoApMLw3ED0uyMZiv
Tb/gfQztHQkAwI/qLMkIRCxSry/uvyLXjtEKD684gTg3Z02ZTAIRsGpwzEZIgYa2
XzA2Gz0eMyqh+VPWUGjaPRN4CbHlxfGKyRzQRINvGVOGasADnWyHMUkzfC+YtIq1
Meio2EE3AZl/DqCPA8WeqYkZDcLcjGE1R3ylqTDlrtG5Tq9HCLel3P9vfhZvzox/
tAYY2cv5j8PbssY8D8For1Ma7xV177auDtL/C3EbXDNFBngjZEPkUmnz5UHzYl+t
aes4gZG1KWVtvgG/s2AVqqbIWQ+YMVWKKidrPjBD4OxvSvkjBaxME29ZJ51zyeCQ
LXlYJS1yRVSnbExV3FkDCDmmJQ1fkPlKvpqTb8wzGIK+Qn1JaMpfG21NM2joS3tF
LnRN0LCxSMN/mp97XulHwOCVnQEmKX55kRidhNr9zBXUfRpyLGUgeLLQIRro/5GO
VSUzt4ujs54wW8uua2BvUWx9rXJWKRgnVZuedWeybkuMHeWExD623sLbAXeKOmwz
egI0y77YGZj+VuDJThQSqqLq5TKVnvo9Jul+ft+qGrOxEyN8nkYPKMbhRqYdlyzO
YCr0jBaIWISPoOTHBW5W6R/yDtlZh6ldnB6Z+r6uF9sRL+/QhvoD964R+nAdGaMF
38ccmCg1dUFy6Pr2b0sFyJBmSgDCf9zrayqXLEVt1dPeuQoJ5y2JgD0cAmAk76WM
A5gzd6TL88FlaQ3OI2wwfSieOO2xbhfLQL4Lg9lPspAsPjaD1fY8pR+6ZHsspjgA
U6BGV/5f4d4JnvHjJUvtmJdP3Z2SER3C4gT8YbNO549gaBGjyesl5l96ZJoUuNeY
aVY3OPAgTC7NI0nNCEd6Ib11bN0y5SnFwQWd7wC8MKoOcCFaGx19+D8lKfbLcbJE
zF5fq8KIX7XglDfQcyQYoh25zrTTblBjZxNLDkVAUmOFb0E830wKH996Sr5YJSHC
kNixYuFs2lBIH+BtpAvPSUfVioM2PYA9sAvAZtZsWdaCtRLV4XSAwKKqo/7QzSXT
ehmJKzr6vOSa1xu5QPnOIR61/ba3dCiRoLSZXIIHhkXXsR6KrirG39J55F16xeNU
UK0Gvs+BfdTXILlaMH0TtCEIh/l4OiIkgGm0DOCuqfz8fBusmGn0AuquFg4XAp4O
hZcboeqRYIsDne6PkhuSUSXRxlf3m2FvuoTA/+M9znV8orphwlkkonop75xtHtPb
f8POQNjgB9XbWwxch3Hk5yWIFtqZuEK0IvpU9IW24A99hxF5yX6nYXxMMGgC/sEN
qL2lxhAHqhlPctNAIHcdf2+X6X1GHOURqlJdSkrRqxbEif9e/b0xbU0AESG5TLlu
+nwIaLPQhatRPCOFWZeo0RwYBJdvWBolwSIXjIxvyqGXBIOCdW36Mf3ptLWFOLLf
5Ko9jnhrSlpzxVqvdbf4nKM+g21/m/+6xbiu3MIhzZWjh5W/8CyBr/3MUW/JC2Ad
RlgNSjLHAHmbN9g6mRv0aiCHTQFZemY1fLSzjT5GKHh/w0jwwIqTIJwphnciCdA3
2S+/b6waTpeDuHz0X8G7vlLE9CONhQi4t57IEXfXx4EbphWSLXmwYh8pL9KDaqcw
30sbP/uiZdHP3vVY9SIWi2JcboXzt6Ks+rubisM2qE3c+x+w/Yhv+d0vap3lsrXm
EUtZ+XKEYsvCQo7mApARsChNnobK/Y+2oNi9F5uM1zKgQFAn1EPG51rVmloIceFb
RP3YLkDHVQaJd+S3yNj/h2vgmH/9qHYI2QAeWgImW1iOzcWfodn3QfMWpuwFuCo1
pjOYckylnx1hObnfqjq6pi9ZhSc6DKBDDOh5E7bSwdH1oqkf16HRXdhTrtzSSYEX
a3hidkVtC7VHTUYnIaCYmnHNzCl84w92Bl3RQRJBV7CdmGPUjwkMvFEwGUUp4Of8
WlU1/im4n94du6UDJOEyns26ulqhl+QGEaNvXFUBvZPHcumj4t0jzkUHocAQLrn6
Cby5d0S+JT/pCBMRE4S/GhuNSrEFmUGJL1al6hLySfEtPBQZudpagiUN6PrT6K71
2oGhsCf4nJrShnMe3XVJQR289DVBFoxLYUb26OoX6a3KsziFVt2Xg8V6+kBM+Ljx
CqfBsGVm1CCJoWvHgomrZLZIRW9QIil3hhInTDh7zc/uUa1v20eZIYcSqllPc2+S
GK9uH5kUtOEJTNiNrLt0/yZXxh462du+Qt4vG0OgYZT03PfORqrNW2E4wUDTl4Vq
Ma/fBjACfnAwdI0WiBrPyHqPZ6Jdj6KVuPAjDM0pzfhNrknCv0bv45TcftiynHl4
gxbU6rZ+AgUVO8fBWloPgQDw40dbhjLRL/YZG8at3v9ulEZkg/Zz9YL8pDnBMLKY
ZalJQl1PrPNVHSu4RjkK/o5CfLULqBCVpmAiC+rq4HIpMOoq3rALLTHXgLYTS6Q0
sjzEg9gF7N230gJ+1voEcYbZXCIzeWFF1DVIFxQwSxc+S9f4xpc7ZuCCoR2Ig5xo
E1dv8j5PPEKhhGtNco96A8ANOEPR6/pyu9HO2yLUEc8Cyg4clxmL8Ta7xU+RKT5t
5xpREhS5KJ/9Dwdt97LhRUUfkOoaoZK0e4uOFyhmL0OdSnW9n9tqJZ6wf2l1CFL5
v4aM003JK03l0CaTHvwkoIIvKflV2c/HzErd6SxXfHwo+52CoKdVrX/haGELo9kN
2THF4iyjW61+bytul1bjP9BHPSTpkSFaUAxzuBNtUGlaXs2KyuTzuq+SMbAxfeTV
RynsVGLc8oEXC593HVTmM7HsFITArUQ/Z6FxPDzp8Wn1keF5FJJexljHQF3egGrr
xw2Nc7kqjdwIKzFAtCgfbukY1ISZQPNnsEUpf9QDI8S+Y3hKj8KQ/PQ48lHUs79Z
qNCh9qVDLI3/fSxjfjdP2Prib9gAIAN4cNiDxBeodMi13QG5MYDKfP9fBxTmcupc
k31PW7YBwwet4CipFgy4fVCK6Czs1LdjXwL3enAvteKVEmU9TLA0rOsjUznehLgB
eyZHK1RZKAkWhdcnPDMJeH9myDhieVpiRrfJotgoTKTAZQVPuFAUJXTz/1vReYGO
wSRMDRrjC1pN00UgKpBjzG/+rwsgbXMZdaOI4kR3wW4BI3lZkDQ0ran07GGNkVFL
mFAH0uAScIBsnZKTrduNRJTADP3DkjOKakXmcJ7h+UZPJDgYQKUu0erd78i0aaaC
BSdl6lARVgJpoLxK54XzN1zD3Rio1ZYMtDG5Gk+iMBCv0EYVxk7I4/CyC35zyA5y
F85Z36ydr0p6JaBnZ/t7pQMw92796VTxl9GMMT4Cc1m7xHFvksSaAw8McHNDPEUe
1wuTD+HSxWH4K/OW1HcgkF0jIOYpXY7nyL+bmAReG//CVCHWz2fz5HsMlFzRXmo/
Wy8DF4vbxDQotLJ58IW2M+TPtCeis2ipkw1YNtbsSqqkvtyA+Nf4/tJ0/3kkloGG
XUhNh1RIv6TqA+g/g9nYItJ3Oux/anpURUxO0rCoq3AMN5mEtxeDSz/hKQAWtOzd
q5UKQoHbQ7+iA02dM/YGmXBTIs/wO06GQBGDvoI87PuRhdhWlWTINddsy+Z8Ik51
OBbAaGJp6j4ZqbtmHSnDnF6MC8/n9NyNz/s8SWwmyQx3w6Qk9xKqlFTTlkzwJ58j
DMQFbfolmR+lXC2q4VpWbx3a6TxV90stTLMhYkZMjqN1q245Rgaic8fgbJLDeAj9
/vEy4Z0YpwnZQrGPrGzd+X5IMxA7SadGT2+rODQ3zt8L9mxF5RHNOLlACefRhGee
TCeekZgz/YsJCLVp1XMQel3kp9wdpnIs76639xArXNyXZiWVwBKRQGAF4x+6w9kV
c1DETYxV9R5RIalQlkyYchxTKFLnFByL58awG7G55b0LZ0wLNb/t9TL6Ti0w7O99
iwZpfmE2vwWD2hwa+EegphAZsY6JS15GAAfl3pC7m8K93kAuiDgmOOGV20Vti/7s
k0BJY2DdGAZovh7Hl+1WGO975/3x7fM8E8QxzaRyeCVqiBIEdHG/YMNNQa/FzYit
yx1x5cn02fND8GLP1ga79IJb7fCx5oBSe8rCyNrHYSi0HXISPJbFTz5VFkjoh6Zd
+8AeeD/bq31U5rrDVA+qf4n7YmnoEMWT6uDY5dvYQllNsiV+aPTgIApkY4N0p6o7
xGIaKjD+88TEUTWlDZQUjgDGgyIw0N2ZaZ2hrorHAb6O+C0gEXeGoftaGijhVgQl
XhCbiisoECPHcNzIwaHgN7bQ+050M1OkR/5t2juw/p3BEcQhWBA1DPzzO3lh02Ze
7NbjIOJyGIRM3Mpy1xhwbT1IYHx5swHdL9S7WOD9tog96Ri6dXgG+9cVAbuAT/+g
06n9AreWMi7nv7hwBTIeGP2gxHnpYis2MHypft+NqSOlGL1q3EyqQrWYLFn9dMxe
VSPKlK3kW2VsWyM2aag9yAf0fkF9b7jFxff97PrVwXqH/Fl7548z/XtmXtATbJuT
MDYx5w+H7CjJudz9iv6z8kFS9kbG5q+ut3IQz2KsyhJ4y8vXSIbqn5LrqiwRT+46
+94eL1TjkJtlViyvXJbJhy2oyuJ3ocdb9R7ynnfzhzxGEE8Gz4LscgxRisOSeoiW
1HwY8YkDwULLWxiyRkP5CCr6VIoliR0Nxl+jDv7fgA3KkLx296qbw3quvw60t2is
iH/tR3N8fj5tuRvSK5QYU+uyLmcl82lMK9ez+cVOPqT2kvx9XzscvOD8gqcs7ktW
LT1ySFN5J6nXyPwZ4MbfGD/WPsHIcDZUoGdTRyd3WarvzT0RyroJO8wuKjgD63Ev
U6afOT0r4lmZrMj+zzcMx6noPbwklEKDa1NcWz44VmYjBpVBA7UM/axtsW17yCYa
GX2wMH0oT5M+6Ha0ncfYSrxOgp56NuZH8hsr3xuB5JVsF4tEvEzzyYn3TKRo+KjJ
BK+mCHKnmT2K2GobDrib3jzKpS9xlZttwbGQqh8p7goAvZLdYG7cAoA4dzS9yqMH
NGu24vmyMrasQ4b9Snpiz4ZvD4xlrwv5NvOSMuqKp9INZ3LPwLghQkmEcC9nl5xF
eh/jmJ8FRt0CxBtwI9Yu8CCNaFpzCC7vNjuyIpPM/mNI3WF+MnLE/0G5saNjadTX
biXi7pc033S/TJtO2WxfhcsjbddXh9b9/gh/qurxT7aV0yTN8izRV2BGlWNqQFBO
O0orfBNrAliHQfzTcjr7K/wckrZgWoVdrCidfK9XF+FW+QOWrYmoSGxc3AoNfril
Biukfm98XB+ZgD8T4VCDJIrap0xlbpwQKvUv+pMhoxckOXbLmXu1RiwFC/ra8s6C
UuA232InDboaFdi2xDsQrEH9kY70VX6pteRbQC50EjmZzofoTCBOnUk1CREM3w3I
P0aGWsusxiHe95tF2UEQM2DwZkKt8GUp+UERw5UUOQPFsoMANyexJKGFmobRBC/e
xkcEr6GNdmdOvGYT79g64STrCJCcdCENufddGja8SGRF+j37fHwfsIvwQ3zAB5WF
90V4/jvQoUAuj7PmpsqBQarRunpH6NwEX+YHlS3mRoXlKx825GZFSfZQ3Dpzbcca
TnW1ciFRrW0FbbR5ZbEyQoULixNal4KN1VbAacLDCVqJFbfKQfJKqIWmrvsvcDLh
gmnBfHD4KhuSRn4+vV8ePt6qDmOcN6RFMBcKiiiPCZlfASjPYz2s7GMrWXawUicA
oF82CT+ySNd823MMnEqlfq6Feiem6lw1uU54EED1+7PQdWDrfeBQ+7HnJAPtQ7t/
f4RLy2ryAONTHFJ4Qf2ZsbCS3RJMpsoqQ+dC0EFUZGfW9gOuULtZaZJz7OJnC01d
9ksXaPlqCzEWu3CR9YUhL3VBNmgIkcNSxZheqdKO23gns+269aLaiHRHQNm/zk3P
dp87WE7JfmmnQGBuR3ljpU+BAXS40xfc91ILO73baLuSBUii6BbhyERTnpz0r2G5
zRv0rYqSerUeVb00W/MqB/QM2lfEi009U4jnk+cFV+Qqo6toq+4QKOzi422mByCn
kKwEM/6f0kr/HgJdiZa0aYbyjXg8NVdBLKeURbO4Lz4mcv/pHJzgixHq8mbSHtaK
KTDza4BJ3tvsjGhBGxzCfULZkPKDUVLZCTSfBZKaKJ/55jNfnJbhHgdR2ZCpvV5S
R9zaZ52MCbrBZ9bFunWNNRFsVwrADjoeS/I3fMFJadezrKSJFI2xoS/ZaajZKv4t
g2NjYCbNQtgicnFVcbGGaBHFrBuHhvpUcD6gOieSH2hg5YOfQQ9H4Z6NfCQt2Aox
dG5d06SURzd5urCq/gjAKO7CwAUOhumHOZcoXS24/nzmoX6UDmBn02tSj53HgDn9
YkbaQxxLxDKDmCYwPERdbdMWaNXPiXvYvQoe/NoJzt6Z0Bry2o8Sn+7Ia7nTasyv
ofxhI3/+Ba6GIXO5gnLutGJ5kvnw0AWUWr2025Zp7YHRfa8FTQW1KzRav0sGxMQv
M+SD2SBhqKO4ESXuFONQcPNI7b6iHPkX0dF+sMxv+0BHto9yzcuSrHDQUlRg3ngv
YuKPI8m9gc/J4qJXv5yu+QSxe4M4YSYYqcsG0tnKMc/xJ/HTovWUaw1OZoeQ9Z9i
k+7MqCpefUXKIipUMjeSiY99v1pLM3FjEm2kutorvdMvVP2AKEMjN3w2Jn/qYqPt
kG4VBE7foeidzUgoLsCekW3UIl/kuxywgkSLhKLDfiEFGX0edO45+6njps0sU6s3
4fuy+yQ0TSJ4gckFMgEoLWERurI0NlpqP8OS97mYrlATkcf0QZiawuY52wVRPOaI
iYi9WV9q7aMqa0ma7tcpHBEXVQEfmLYIB2svKKGwDZaytwdlLEY24RkzMpGw8ky5
cjxW7jKxf5o5I0CYAul7j4JwFCiTHHjvDIMefRO/oahP8AjIpT5Lkz65WGdkQ6jS
BrQ6eTujUc8hnmPxdpcf3OQwYBfjH+hRbmusnbXvQUA+Ly54tKfs/t6bXjUdZFdI
L4Wqq8IDqItZxn42RQbF15NFQRyg1LOH9L96mO7E9sFgCncvKq2F3bbH22gsRlNN
sK+BsN+Cyuyy4dbn0RynP/tOk4Pk5b669UgVgO42K4CIgRDl7Km/FByQkRXSVytg
LM1VtQUFncDnSaLPms24hQsxrqjle3+r5J/oa24bsyEyv+jiKtVa0aZrg6Mvro3G
ezYB/V89ThzoGtEPdp6Kb4KoQa1tpQTZe7DXsu7uLr3Ghf3EGX0U8MbcmTDOnhqv
QBzq6mQrQmlnsIjEE4Ae3BBMULXo0+CLimGUAGOzZ3MnkdvfFKDBB/+LrsBel8bP
0+8+CHoZhA/zfskjquKvOXO6F9BFjmVmTtP7593kJ3tiTPQ8fWOn6HZqOiaicVlQ
9nd+RTLRtnXr10lJBZRSBZRBNqg3Z6mJzqD0vvCTfx2tmSdMeDz3/nGpjOn7jORq
u4EXzs/3AyPaT0YN1Lc/QncZA1JxjyFuX5rrn7lflKQc3KTD4VnwTgTq8ZVb5lnB
VFIAqtlIiIFFbr7pAmreN1nylXDOTFL8mpD5Rg5Rj9kpQsl/rN4vWOe+Tahkel6P
B7aepIYRBhTJ8ZkXdMR5QrP8fYGGay8P5B5W6BrVOm0KLmPorFt5u6e5hdwU/pD2
WHL/6hrniFFWG2/3yBnG7ASbX5q0iUF1UAcpBj+R911EDYxW9ZTC94c8LIJZdeGM
HlCglr+fQdIyTBoTyr+le5+dEsNHUfrCbUVvK1U4ctQGkgoYo4eTYxw5JUtPLPIo
N9GxPGGTXhDdpWuOcMrppQPZwGcTzn7xYkpBh6grf+MLbingz3nGlrUZcgKwZb5+
q/Oz/NvpdhX+bPtmz6H8hCsDSS7bVD/FYcmzl+OMa5g0P+O5hwoApAhTe5NXoPdd
o9nNKeeQp3Yq85AtGsP8sGUMN6jSSYJawUHpnyA23xMI2TncUzftVpECwIhCo+oe
KDJybIk1LUDvFEd0jHr7GsCM9/KOMkwLZmLHZNpNGrHPaxtQ5LNJ/fZkFldsOFzC
iiuzRsKeinTNZpGYxfhSoAyt++7ggj1qUKXJnxkHrXUsiLloZOLIo3ti4gVfKqqB
AFkXHxNdJ/oIK0b+LExzWlva2An/FyUtWF04lOBGEh68rvaLlKgcaMESN0Ya1SzR
tAUIt82ZrOf1GZY3QYJTQ1v3RHoUOJhlfBg9UbsTlsIDFoH+4bx9J9XBQQd+v2SL
XHWeb2QnvsVkxV0EtYipi6KNKwpGWE9c9LJv+dV+1OXzEqFL5+wTbWgRLoziPSxe
R9+wixJw8mamaLXJHysDlDP7xxPoVOrG6JmGNBVixJp9pLcOiiEnVF5y/xDcm0qQ
aT8YVxrCmqQ7tLj8QVioP3rdVnBH+TFGfWV9NPlJq0f3zeWUShKHNgwsU/BlYxjp
Qj8Xdk9T3e49A3yWiGc2BT3jH9xPJwFDAN4ZyOf26kJzl6cd8Xhf2IkgA2XOMZw7
1x79BXIRuugKuwikWGkAYU4+ru4npH8DGiSCfREtb6n7aZH/v1/bwKGhUnWouLzG
EiKf83yg1FTTeW2MvnXmkd3AODw1BL50ULxQOvY+W6Mr33IOKZCYQdh1OYF/nQgX
ncRKyath9Hl95+JjeOlkgHY+lCnJnJQbTsk849uo0AbPeWIBhbkG+cl6V3Rk0bXy
oJ+ApxdCsbIEBmSxmHTP6Pgc15ZgNS24a6zn5+rK3B7vwIkgPvgTcluZpsu9qzdp
C+4vD3Yo43MN4BUG+Sy5i7Z6tQIB11t5twOH+AoULebXcVbLCzhrQQ4bu4BxsxGW
I38Msi2VWPFka+C/T96NUrIXfcllxU4lQTArgDkJ7iG43rRX7UmKKiTnBsqQreSC
y/s0AI931Au9xTaffk/h73F0PtsKUNaGIq+sB/W8Ve9KNIBX1wG9TxvH9uypVFMD
xqaTaExMOybO6/sohkXl2fiV4I1n1eW2MSV0+y6ZjRjI3CeJiBc8NIwth0m6u1Oy
N1XStGRc/zQ6052mC3/TjWN0aM/aEkHSWtH3zrKsBFs/CJ9iser9tXQ9x1eKblcQ
lXA3owEmQGHGmL98hwFpfVUQzPgQZMt4EWWxsnhcgEcYkz16bumH/HskhTXONvL3
jUJWHwJRNEvzwfDodEIUjYgc314lfB6sNbn+lC8uozwprZotcUYM5aCBQJL/ytHN
vPxdijxlDkUgLboPOIHOU2oM0RMmHO1e6JpPdgdJB7iCiM39SjnaIsBqjreL8dfO
D4jsZsUDh6SNCshpgJp7uJWkH6pKY4XD+sGBokQSex5nS8qMvu80LCTX0WRiisC9
kECADudTqosVt27Ubka6ak2F2eKBSDB1smRzZG6hiEVBt49nHsT49X17nL7Hs/3G
BQ/9JvKXex6OK2mAe6xN4pX0lKxYJ/1qhdhXgxPeB6aHcQpL4RYEA3GKOgCFG7nK
vTnMF/InzgPlMmnW/GjA04yJsCWxK1AcAviXIOUVnYCU/GL8LyyrbidxXw3+pBQ5
qU8uMQTcu8Kkxgqjorg8KEjDVZtU9qJZLIbfJB91teOgZumRuvqlva2Pdzm1xDCn
GZ25wGyePeL+UhmBck3Xp7QCHwU+nD+c3BR04wuGa8N9sev+nxa0VfUkVFGGgomR
ORyc9FNO6QR+IAx1TbaV6kpI+mMDzylv7uS7cW18xGrv86dIfKQGqcOUvDmvLj+G
PGy7BkQpdkXIV2YXupi9UgyAXseZ1wirYp550d8VO6149ccKdtG227j16uO2yp/J
7xqQmecMny/XbcXiCG0Ff9BqZ4scJMYA0HGU/TFsBZcFq8VnGy/xq+xqgruy1HW7
gavftm/Sd3aVnLO1iZCmk05y4lAvMt9loG8j1Nxglv83bZSvKaSI1TcHof7QcJHT
vCADT7ga0Ur18yVXG3pzkTGzEX+BRdwqCGfIzApTC6Grp4/hBqGE0jplabO/5pIt
2Ni8nytmfWRZ3cOV+54kX3Y83cDLbBb1+2XR33OlFdzUbniJLJCU1/yMUoEGlMEV
6Ez0est9nbIs9iygAjRbLFrxJ85JaAPHea1MYtfj4dnrZqGo245Acn4se1nhU8eP
ZBxczbjcAxEgJJCS9pLcqacQdZ8NPtnRMU8252ytO5vqs9M4GX3aNhMSi1bijoBm
4yuKZKROzBALNxYnHM2mDcGRB1VSOQdH+L7R/R4k8BlbX9N/ETIb4bWmoGhEL9UL
g/ulXv8v643zBXFTOmX1ZrhPfz601DXMw4UiYQ8jVkQzy6cDdYphd4JhCHczybA2
3HRHA8wbGTjz3JKkagOQGO93DC2HtHiBy3+PYHGnIrsp7wtlOshj88aGmD0WuD3H
WR7pluW6UkohpbvUArjxHQBypHGCisherYnHb/m4AnHTBoy4XqR4RLjoollKneqP
vbEyMI+yScNOToCMR5A4iIiSCE64cEQAECMTjsUXqyDLjc8zUGWP+EYXbr6cfJiZ
BJcpJ9d8jtLMnP4zPycVxYcl9ZF9/jXeegGvHsLhvL5P43hY4c4JjE1xmeemyaO7
gByzCQCfN0L2oldXMhzVqUE+/wgdv36foJtySSGXuUFKZ3QCHtdqgAPiC5YdQkD1
UMl6pD9XKfAqlEFWy+1pxLfPDQCpVThp+qsfL2dGx+E25xdUxPUKP1B17kluHKx2
jbyilHQlSqI5aDYxOkMst7LJ6fjDI6uOn2Qfsqw2k8YPNNFB77WEIi+DeMvZU+jx
yMR+Dqs09ogNFV3L3PlCQmeqNz8slbkyzi5yjOZe/mskNcCXxiqgRiUKJS3QXb55
RXhPL4kjSZ95B4AOAVl3orNEQIpNo0VbECaMxqXYqx/gWv39IkMAJfp9ThGuUjiQ
y2XPtgcxOjYRhl+veZe2doyZZfnZNZqm6bZzsQ6UFR1BtxigyBgx405I8cecnNZL
QWPijpXQ6HZZW4AtNYM7amd+rN+25+wohCpqOHaP+3wq9v/Jdnm0UFGXTvKnE+cw
LJCRBmydo05R5FHyudo61SnEfTObXnzoWHkdxBUkvEn+1ZQgrUjJH9WRgMDw+aHA
RbXE5OICdRY2qkkyTalMqhHVOxpadf5X7ioxIOMxlFaaMJMndVWYMbDGAU1Cnctt
Sb9u2yM4CgJCbVCfZZkh7b9L/kBiVmj1BKFSq5m8QUB+iNXBSCeRPiBT5BO8O2BO
ku3RrgVO26WTRL+kiBaYGmKClO6dmUE44HrgFew79HaeY5gyPBAhMeS+LnfWKX0l
Rhhhir6Lk7ajHWnBgPo7JgNMaYn/nMxD4oKwBzoPBshcfUY48qEskzJ0mwr643/3
6iwE1lA+70ExLDDmkjTTJCi4wDw1Ydwx71yti/LwZWM2HSuNbg1X/ewf6464NhvD
vKYBxgYmQJ4CqZLC6u/c621e5VXqaIoswd1wu6+xP9CHsDDpTSQWlXhg+lvYQN7q
R2gla5pu8qiRi3ShNJikGhyebgXiR/WkFbh7T10szMAw46HUjACQ0R1x5rkKnZho
4MqreuweTwkAPwX8FBPJxkfyFC6paQ4D+lMOzxZhYp9GeE/SjKmD7ib3/HkCt/qE
DygN5VMsAMV/GrPpuOuvaOsH4NCVFYReRRoXheCV/Cud3V3ojg2+oiCig1SilEcR
hYa79rQku2HMZ/q4nn2HZJZnQ7/92tAZiyYnbVz8LINc4GXHW49ifj5O29tTT1SU
7cmXzJGQVGTNskqwi9i7yXqHoOtxLoTmFUqSHIonenHltr2yMTnDa1qDT1RQeoBC
KCRLvpFxI7YzlzZ9ghb45/Vf/cvo+ncNfOUKGq0jiXSQfkQ7qd1d5KCnk7tCKpuE
BlFH6K1/16mhxv85LJgaEsdA9MdQds4QMC/yWQNfI1AtXBDm2kGurYndn6o042Im
vwe1RCd7bNZA/HbMiO38ZYbfPr/R+iyuRk0N2rqo40fw8SzN7pXlw5kHoSMBtS20
2zp1Y4wezsdp1hlLiJ316A9RFeOZtbyISxAoby0A1ACPVMDrKsLl7VRj+JnMwB+S
Al1sfhveKC3YgLoViLguumVnpSJu2m2ukB3iH7tuebq8wfip2kd/F4itoLOKk2Xp
yR/Cfgr2DYDm39yZ9iH2hc9/SkptxoilYs7EKps3qywOyKgAqzcAhsO0RptbVRnB
csDnHUS3ZLBOP4c+BqlX63kritTSjB54XEqu5tJGO8aXf4qW3B9jLMXgAvKgXb9U
KQ5wiF/jo10KHSiFKFm0D8BQ+dQwU8S2gjgj5UGxMzDJFz+7/Qh+Z5/g/hNRMtOb
ewGrx25jFVdUGIcP+MlCxOcEMb8XnbUB0RxpVFzkW80THV4B1R60iNQWWnZ+nRSb
qkP69RmUK1i7jdSPI9QXQXrK+dWflcZ3vffBm0ktJnH1JA6y8XVOVIfLtW+Q+9Fb
TTCqxetT9e5aVFUarvUztNrgGm8EY0twibYyzdxrN4M2YuwgDfUvLewLw6tF+m/f
lVgpKXE8xuT3IqGWnZpNewAU1qZnsuKlsrUCyEnZoCGe56uRRZwPQ5d1qkDUWcQG
ZpHClVQYh2hXU5nXCMXrEXR/Gxt989g096DiQ3kn5mbkh+LWWe/vBrmKx6QYZNk8
ShSEIuRnzSWLarvk4z/LoDZBpGSB+fpTLSAklwEOlvb4GooQITmlgH7pRe4Ey42f
kBl2rSCNGkBd7Hp8E7LHj5sxczQe2pTX9TyeAPm+e6BukOrF3/NKhyatxL3LuBK4
r7wk5yYwyt7Tyd6mWrS7cuTc9h9Rg8/clis0FUQ8hHAHa+7s10V/vpyldfLpl13/
ECo545U6ZaRdiPcxZ49Rke86pf+Cubw9hzCZ8Rm5zJSEDmquEyN0R7MQTKSwKatY
i/YbEsaMqj1Com6eOv7faapFOXmAmshubj9nFsrjWjVU1v7tjA4UsOm94zwt4Sg3
2nmG5XLlw/TXF60D+H05Ac0H8jY2OQW6OyLjGNCTXsKKN9QstlV6awCjwoflvjEt
nVQ9cvfaMzqJQ6VkHUf/Jbc0ILphIA+Chq/RQ7shL3B1aBqOeB3gHWp8yDXYi9qE
8SMmJboyMyne6VZXVxEC5Vuvq/r+F6IkWkzwJdzP5848S28TDtipeVaH55JAxbzH
4KHv4PHhVCXLb4hoB6yxEBoRxtEOFPB193pjNTVBlL+ih9H0AC/lj06DULrYuWrJ
VlmmE8BHUI0viffG+tLqbq92oRI2eH9Xb1RPx3R2M0V54+WzTPb/e+GLVnUtLA61
G3BpM40IvrfQgKrwDPacMb/gYQIjM3BiEKkuQQsOnilSYEE0DLJlP6Kv2YIPrnM/
P99s1ZDoA9bwu65yubxPJg3EdiktZoYCDpnp+d/3RTH7yOXeBjqSn1DEVV86D15W
P6LnY5UqQi5UOrDAVFNFLMTh0+T75gyEIZ8t4QPrm6UGOhuHHpocUjE6nmb0bpgI
cwgkXmDnLIdzSi8WElF9kAOZ6BfOuYzL1tmf3EPFzyuf+Kr4DQuU79TDSv7NQRio
+YnBU7474TK472ZhdwrL91zcED15MmW/iSRP+za+nK0Qp2cUDZ/JufQ2kEQd+Lv4
/9AOzwwyzDOqFxtyjRJRyodkPsyohC50WPYwzo5vwCFZ4hiPWYLimtgliKldT36O
dBojdcSlnLr1txm1JasijgAWJRG5ZNtvwcss5XwQz4dOXdpOgUi/BcNv/M8IBxu0
F7hDEnbJ1mGpctfBUJaTwSSbA4eC1AxasG8WzI+uscqnelqVA+QitZ1cm79hcfd1
XPcFTyiYDS67xxRPX+arMDZ08UauzaVCYMB0ExNaR6PFdMb9HfmYZ+C+U0cVYwMt
vE6PR5rWvWfHtjAvO0ug6JFRmkAQxSXspPXrUw7q0iq+AumGkPEHQM22UOj6ZuJk
N7TPCMw8yosvMlSmHPAAnoP8VDzPPIib/dC2F+8qrP6PsPiI8DvX8ZFEe/WiChPv
roRzf5QXuQnqDFA9QyJfhQ2SRM+zqT+unfkKzn/njFvtvWJGRbOByGw30YBKIerq
COS+SL7UEco9mOl0rOEuWMa6pu0+u2t/A4+erVE+2pxCZrGDHUW1xZ2werMnd+6s
7HP3JdIlGdqm9KNyExabO8AmJo98CDOSDbNPKZA/A3rRQKPRV/XONCgSvtOgvAOT
gjpTFzbmYyGGCe4pvT0N01qeNqbo369GJbbVWExUrD6sn0fAObdtQyVglNONUGLu
6cyt2YizqCLJw5Yg2zuVpKIWBwEJYLuBBaHkHwdoPvQvdKBmtF4MUBHGcFnnBsW8
pmY2IT/ydfwgcnVVz4m/ZHcDxVKPiJVCrqytVSsoSeO5nVHhwq60SUK/452UrZLG
dUGHFDWFXz23cOM822/H4pazGL9CEjm5jG3uyYWYIAz1OwIzg2LAd+h35H06D6rc
4UltHWpKw0hTL25jjGC0vM68gg6G1AjWvw0FMD9wBwd1PC/s1kraA0+hfHKXJXNa
/FpCpBQ2Hs/lo4f3GVG4Fm8OOwOfp7jLrUyU5PTHTBR58I5IOGIA9ssQZbRyNHav
MHHYlkUkXurW8zt/sLBY2i6bBgNgKehMOCmYpHIjiHW50Ll8xezymQMSvWNjyc2O
DjX9ozE2Dt1/JFryCT1Kp5yq6CrSj90igluWjRLGHRG7brFN8Z0w0tFdj6HVRitI
kAfAwJdo4SjCdit31FKoSfX3uBL6iap4oxXF8bPP3NPSvGHT/+S3iySPYRqmBJyV
/xlMgnIFEwrdwQQXy77g249iAwHaCL6jn4rk6/WZe+23i2V5mpqyM173lroh9+5X
wEOd2HXFDZK+49oZOWpHrPEqskMQr4vFIq07AvZ785DxPDAw+WgYuHK3dB59QEB0
nOROvWowm5js6DUsv10kUGCwBxhcC+krQ2XT07z0iB+fWn8rPlESjgU7sY+WB7OZ
EB0PSVxC2WQ9RnkqKed1C7zhLMIhPcmkqGeFoayWEzgQS8HPI8EqmQP1Imn+aV0s
Q+IaWEACetBFG/ozNnK40mM+Cy0HAyU1YYx0YR+De9CLYKvU4g605jh6nDUtoypM
cL/aDzK1Ic8RGAYMKC2cPGA94hMiaC2HItTzL8fXSSLmO3AI20UYkLNwq0CpK4GS
gwfHqtMxT1+ZyH0usbla1ltCYvKC1hNFvLL3gCjWaI7tOJIm7wNOpN9rppVrrH/o
1Pu1mpLuB+OD51NIfslgozczosCZwxnIcjmoQpZ/h7+0y3Bszqon7kY0IZd4kMVM
dMfsDr7EyLTOlyDc9eZdwxg6SNQdG8MRxbwDyQ3cY6XtrzTDOQ8oAtmqwQTNna8N
vhYcyHXzskxlJclrXDxcXgYbOh7YB5BuYMWayuZmdTDgC+to+EntDOXxUc7eJhhz
TFvH9wpymGsODoOleBrix4TWpaKnPqPRCroRZMEbSMAKR9Lk/hrMRMi9LJPR3OtW
MWZ4xkYQrlkuqOP6vsYcavkoUPP5ptx7UT5JZ0/JMxbgMTtsQLwI861uoOA/dDk5
8wREN6mSuVbnr2mLJuDbpacL3rpDgjCIQvz9pKEqLY/7qzlur+Ic9kIt13mU9v63
PNrhO64MGST7EvkOvq481JSFrO/yMY7uK+uWJGD5FMzjS0vkCz0HZ0kigugOnT0a
ztqa2/A5CeeTzzMJ2B/KzTB2t3l/6eIhHLmGMZsccVkwenZqGDsmjNT1jBHEa8pi
xlZK8kkLHEkgmY2bJdMECqWgRtfvSTr95zkMOOsNuH0oV9VxdHkSBwd200t0Alh8
1Xi5PRa2FsYIT9yWR4y2jKB/Na5LWZ6czFomu81tcpwDNsWi1xpDMBrJiJl+mehi
ctZAPgVk26jT9c/ea6dBv0n8qVyhAY6uKUhdoAipL/LgMyNHucnkCj0gNuzgRE8c
NKNxgTC6q9y7vyCOtiQJPvm8xRbFmb3KKoZrPY8aPT46ME8Ia1yqT9qQ3gf4Su7z
/q7GNYXZ/Zt9S50WaoKnZBsGX9apoicyWjn/RfwcfbG9JZ9rnPhxYP4It+Eutl8u
YLHRoqfkWpfX4jJYQDVetl5BxmjLdN0LXWKyujCZaLJhR2X6QPmQSYCgyBPjqED8
sU81sQDroiL2yQMDt3aCS0cAixKPKTOuA97QuRMa9OA9VCSzmVusnAkcOBcV5+AQ
PzAW4f1gL9oYqW67mSlg/kCfjgL79kh+ZwPQsYf7nmWfDhQazKpblGjYW438/AX6
H+wvj2a0+Gu6KatkLlawQ9xUweGZrbxnb31tBh8SZwlyTDWoaYMbDwksQnbC1ptM
ziBbypO2gMLNuhwTym8mODuXonGM1gV6D+iLrmpHPM7JBdEtmsa3VFbRALleC0/U
qPfLpQJaaIeWyGn9ym/i0cn0E9OZkKoOp2XlntXzlzf+hCP4c80b1Q1zNb40emo9
RWFuCsMwDQN9DPGszpsqENlpmjEL5ukDg9528LA2/e2KgrS2waC7/4FEIBej6xkW
n1qi9NfloNbPGsEpBNZk0V+ZxtxnBMQFkcJDBJxlNNhVHXdNthPvFwx/3RY4r7Rt
wOaGzh+1VWNsDbMoUPLFVIw2EQgk/33G4tC4DZXA2kafy0DmzW+LhoQYIvyf/Saz
t1+rFkToONAOOynHmm+NHj62b71LL4Pv7BPiIqHORNyBgcEVkA72D+1FYTg+OY6N
4AJM4ttF4C2d81Rvu4q1gcwigp1ta3ruSAhkCvCGW9fuI6e28smQIbRJY+5r0XjI
jjp/XO4vTDz3rE3KFgidaVD2YiUywow4oRpNi+FVqQvXiZN5NjrGrtTa/KE2YM0T
pRXl/UomYcIezIR8OUpLM8lz+oz8+Djz0yqf2TmnMRvmeaLmBQhcIyasgp2JuIwN
8o/KjGgaFl/xMZ/k7xPT3NOGF/ZYNogSzvfvrTdtc9Csga/Huyuw6KpzyQHP7saF
4z4fjlOkrYxJ9O+Q4QhL+IaYZXm/eoEhAf8BflVfbE581PZE9D2zIrXQ14z7CiAG
WHmylszBCVagY2VHO5M0OSosnyNDp4UzZEoK1zquXl6cCF4PW06trgATSY/u/Kks
mQZzvqxDsyxGowCzsXr0n3FMfC5jb6Sug6/tmk9eL8uKzmpbHrGb7F2UIWdS+whH
YU5TjkGsVjCQSbAHmm13zFw9wQX7I7Jb+R5UiTkNXVc/k6H++c97U+C/0tFoz+UF
RPWBvucwHemwYMIEN8cOhWMHnuS1H6zECwQhKKuxouooLMG1p7lU4BjlY8lUR+Xv
qOKFc6Cl1iWSia/dS+yjVY6pqjMjO9KsaEZxik1gO/UEikzYvRHrlQx4LVKRdHCI
Wb7dwp2aVKvg1ZeUDyIZBHRaV7n20BY3zVwrmW+5CIwlC6VaT9ZBYIbo6qmZssME
c5t//7RPg/wsEsaBIHHOxhoSw+taZ4TqWfG1/Mr0MepdJrjQHpqmho65hQ8JIqOJ
r30oAU6ejOChxlR/E30I0gMzN9wT/a1fHeufHXWxnR93Ek4a8KBvnY/ePxaaLWjw
hyraWPxeHa9qF1s3Op0FmOQyPvWgO1lCDW/Hr/yyalK8exeubYtpw6LxCTJiJIPh
ZfplD96s8wnSSwyA2vyCms+IGQPBOmmPwEnZnKfOOsSsc6HwF9jHWb+YtIUYE+oW
QElBRO2NguGYPjvH0O57aihsn+6HKxcWodO9X/LRlSkLGwIaZU02m3IANNDJIOw+
+MevgH+f09R8oSF2USqEsO9RgcwTZ5Lr88rTziLDLhU5lb80wyIo0mE1lCwRGgXN
zI29xaSaRGQgWexC/QnGQJqW6VWR6X+1su71Ofo+esYOza7OzCaxwiUexn6lX5Lg
BXebAhJcJUkuaXQaMfoaWdq6eLbC5QI0GTaciZEycnpB2A+VDIXdyVbByda+K1RX
k5iqFVfI5EKHWXKrdqU+uk3SlMli1Lyo7njd6eHWWUUDTzhyOk9KnXuYGOZ6DjRC
0CzZsGIa1adNnNTyWO8w+B9FjdeCpTQb99wpxdLMZuOZPObkIn4JouvMQCoSy/lB
F8J1oQPYNGE/Ni/I3DP9jdsUO08Yo2YTrAx9FUApzhXfRyCN0UDD7AFeNvHkuPiV
EIt9Q7bmfeNs1J+pxRKHs29AU+bydKshHQcTSeAXiwq7CRq8gCABjrGnKE8y68y6
cNpYgWpzqROIH0GNGW4FDIhVp44UWlhpjbFsI09L1QIY4L5BGEinNMaNJfYaxAGH
cJH0/5+QKuvxb0yJarh5yzJpLr/Nxchs6MAS7m3npTjjFRc5PlOT1h7uRx0hpcrM
Vecafvhv2726yd4VBVpEEL5G7LkvQHQ051gjYRLKJeQguQDlau1CLirn4pne0HQV
UZXGNFT0MIceprc8lcnKCt3jiLRfuyYWheAJ8878fXiq8oTUO3BxjvWIblAhkfak
oJGiWmISuUu919sncuQbtGj3adPnynkYzrc+UPmbHo41d++nJmHezlXGfUy5FJlC
aV2Yn/0ipQ3MSrthiwRoPrPcPjDToUEwfPd3w8Cl5jpWTN8Qglcc7AseJu9mKO1E
kEmy+nHRxhOpVmY2OQs1/Kea49+JGV/TSXws2raCzvUJt7zcRVm59/2WboKoDiqm
CshHf6A9Mnyz3GzZ/0hZbfRdT4LL9FDMTjMX/1KyJa0vIw9mi0MQhFCNjfIcScYO
iGmlUdN2Z77pJxPZezkjBq8+HGsURq3zdbVlH3PTKuV0HQmMU44A+i3CaOBVTfk+
lYLHd4rz8F5YxFENsR5sZysZrxjLMj1EnxtW1NeePDYUXBsBY9QcgDPqNRdNAcsn
Su1a92zpr2AtFKbiouczkO4Sb0T7futA+gwDKM5i1lXJFaK8wxWbCytehxwCvnUU
X2ColcbubjdYTRL+a108hs05h3SQHVKcemyI/eaKHxpmN7sSRYYA8bjv89vPT1lX
LxH4ev4jDq4cAMNOJzgU2pYs1NrxqYaBRPFl0EVTXBuC2S8xVHWAIE/IV99JCx8N
qBTKSvkIgzrFH5nndNRQYJECp+aLuwjldmTfRCgcSjPh8qMd2SNlPJy3HA96UF3U
hVtNccRFVDUvlpg4xhzDy8IK1VDC+RFG5oDDVJbCsn0A9FDlHsS7m2kkO6CLAKum
wy0aKZHLCO91Z1UGfCqOwfyRROxLz0yPebex6DgUh/+6T50hqDLJJbO8dhWGuDw4
4nOZVvATl8JqtXY5LnL01y4Wos6Z651AkGOX39FG/N2ZQwzbPqkUjFUnEq6ZxxSX
AaZdCm6GIjgh//prCA96ePIlj7quIvHNGOevFMDHx/xPYFuoMQFJHFOH9pfQjAdz
zN3za5PQ/l3K7FgTtlJQvVfOy6V5i/1C8E1w4bAzc/vUYazcjerdPTS5zXHTHGKK
jGWZCJqFLBagRQP+XZLByretV0KDVFz8h8SZlUJbGhgnCc9AiB6YEScLhffUSnV+
5gwDe4MnUvRQdN8dJ1kC97HJ16oyaolMDRq6wA32C3BDrSDJtAg/qbtyv6J2ZjCi
6owkYYGrWoeKggmvC7pa498tlUl5jjzcHK7Ey1gR9r2AoSrojoZH4nSEtBQhYAtM
3du7EnROkeZq+6ogqQK+F/hdNX/Kl1Xj68fiWcSvzBelKLoNsChDtV5Wh1d6lgxE
mRrMelFi6uX/HTr2zGwodwIlvFd3TORtqGopvEkoLg68dOI2OSAcXueTlA7/HJ+K
c1D8UcZ2JjBPDh+cPNNVk4p5gyeiIQ3AOREzwh9MXwt7dO+awXgYffI9UF2h4acz
XuSlIl9SCa2frupI8O6diiNVCku8Z3UebbyEp6k7YMpOF9sD5EGc0POTxBJA4EUu
EyIEdjcXjn45c5VyMROjn+W7ou8588rTzOCF/JtyI4n+XyvTTW0sv5wJrIa83Y6u
q9ONQn30KxikJM0shDXxmSZiatUY/FGA6Mam2lD6G+vD/i0sm/pRvFumIhtbFO+S
/VMVe9kfv38+0cgiyff3rs5RMSJVy6iB6KIXKHpg8Ia+2vAjqGS55V0EGe1rplPR
xoKGW4pldeg7/t281FjrE5tJ80l0IaMPIbuGrJBXGtIFxLEdjn4ZiM+SSOLLSJka
tM+6lHvwL7snva57lDs+aBS6daPlySGRBV40OTNzJPYsBEy0SsLZFVrZ4e75THeh
V47DvU3nIeUm8DtPkzXGfKEzQ2Z56QaF3J9SDfvRlBcw5FTkAnVjvgpwuljN7dHr
di/crEKlPH8/QYTWZbr8+Ev6CpF7F3nDy6/QgtU5BJzn/CiPTomOGJFcXMrFrk2S
9axWCs4mNuERGcLUa6I/4QWRvsp3V1vZvaTtf0VqarQoJYiJCJ1mUkCYkv1OfQDx
Ic4c+HKRYDt6d1QTPo6bIObTSo9LQNPDvJX6wT9vwPQUJ2pOk9baHZiXwk2Bjein
EcPyuKrvWp3S0XdyndhkGttvDgxLfhQgeMBrI0NbnsiCW17tufgnxp6tmUvpMcQx
27X+kOEGELbEZjdLGATBjH/XMqGwChubdJqyocPF/vckyLHxGdIyGDqEUZGv/sss
lClreOmzlsM/Vhdrf6o2M/D/JhgNoc1CNwvMMVvh5SYxgj1fATeR+xjSgwLpYPCR
olUjOTDdhvlXdT0t+J9jtN2ozhc1IFaPndnjA8R2L2sPy7SPDp8c44C/rjrZz3Sq
RTIyjVqscp8oCNIKtvi9By8nUTdP79sULJW4dOLbxSyFO5QcbMvr+U07lw22bYCd
CJq4zHfeEUCe2G0pGFR/vlDyEGWGGAQFBg97085vO+8qUDJ3tIkI9LRgdmrfbyDe
VT0nnJxuDiAmCx4+OkNUhDMByhaa/sUpz3vjzcdMIgSHw0Ci6esbM9uk0kySMCjX
5pjvMG6AOAgKjkz49OLZ/L+64pjVEmQYa8ik3eJn3Hfuz0rcFfDWpPvs+lDivNbc
7LMRcXZjY+2zQAJEzeOqaaqUXO9ibKsaA3XrTFqRVScqaRTICUmaFp4TWHkvaQnf
6VYc9v/FxA4EPgC8EaHFfQNwlB/rk4v+hKuuhSaSDXY1r5QumvMmg8O3qL/b8oPR
tVmo9/QaoT0URc8tgY3hL1/bjTIdlHCow9ac0n+AvaXeE8xjj/LNYX5PDDY/TXk8
cktBgeS69lphY9rQZOQL/qq0z+pmwui2K1pJNhe40u0XO2pcKuVbQUCvOYVuzu5q
0ochb8aezhuTnYGkUAzWfEkGTjBeK88WrJ2mejbwl3eBYw1eqzoBHs+Eo+p09cdC
hHR9aWcOPzw8fKWE5iNpePZOczErW85RPJ8Jq7PpuiLi3JamSOsynZ3jtPCeungJ
FxyegWbWMQYRdLQCFjTx67dIOO2Kt5KTRJ1PlTEx9JX/ylawK4NCsLGPPEETQKrc
NgeYJF6a7s2hzYG2BA2UD40LlcX2rCPyGTRdwSnSIuxNnpINTGByln+UxCeE8TNq
P5575b3ZSvjKakwmCw4raQz6U+SGJmF7KSgmoxPNgb52EF+mKq8HCdDvYAY2mwVX
QJBSpISk8JxpA6pxIj3JWpi24eKY18uJ7b24POZr+DNLXlSznGerN/asuZzM74ZI
LOexGhQT38016EyutQs6yPSJuetar0VTfmY0MHYd6hkfAfhncCj9ghtoyFViKYB0
eLnrt8+++fs+mA2Lfl2kF3mT8xYRhIJefuLftt+LfeTAx4sGnVRRySltahBbquh+
ehdqOnWRWBr1z/7oyTOkpYzkQWwiUT/eG8fcKm/HKUMCX8p83aF/vSt6fEM39oXV
3vbjbeyRSEWibsagAbzZ5fWyHDeenwbTL1UdjNMVRhSSR8eMbp3OPltlL8iK3I8E
1aFyaDmxOOZ0O99c7PrJBdEUL2pUBoU4X4IgLAMUojTBUvgGXJq7Bh8Bl6UDTVmO
v65WX0hRbJ4l2hwOGT/Bw15VgoG9W4pI67y3Dj+ONJhBm6HwJ20YZDCU8t3E97e8
SRsENnA+Xl50CObC+gz5O/fP2G7N1ByXXIVjIdpBtGGoknQ3NJxJxxad3oERzf+r
Vkl/X67Wq1prXiG9IB2ZVoaLEzfj4dTbNfVm+s7HFpecsFT8e5fflU3CAJewBV71
dn1trru+KX/KIQofI3Sx8Ue9wGvC4hfRcIvWM3s6m6vHR0pBOvq12wt8G8kjTkwi
dusAAXf4i6ESb3hlBYpZ25EI8iQDLVcbBP0ihre5s7R8REUpsAKbLfbP73enIDB1
HIriq8Qnx+sbkwoCw1863xgVc0q6XH03Un9wZ2R9RHJqIaJR21N/sgxjmj32H4/u
uWRlAPrdZ1n/U4uAXVWNF/VP0ICQhAOGVZF+Qzvy82Oq7k/xQeBAvBp3HsKLsC+Y
JbEIrQhED/Cbfgik/KUMH3IUj8T2Ej6uLyTF/Jq4UEp+R8E3UJdjmOJnMTHzsRgI
J27YZRbsXO3l9B0r69MYduRyRQlalGaBQjIEf/3VP59yNXFn8CMdsx3NrPlqZyO3
enC0MMkq/k/pbGKHHcId+pge3mSXo9KivT8Z6gqWm8pMeSg7gZfLwhZ78hdvvUR8
JAm2wKG0h1Yn87mySw/Cd2EDYTyigw/3RET03bF6iLB56jGRYb/LE5oYWmdppFRU
a8lFunts9Fpfgmliv8utPRROPz4JJBC1Xsmg+a+kBjlPEMEx0mXGvfDyHE4wFjq8
2tzMsltpdhd0Kxm9zg0Msiju5ZNGHs7hbZsoQ593Y4/a19Nfb9pGS8i2fV5K3+QW
Yj37O5G9xzVGKOTfAUobZCHGVtxxC+mVkheRQ7Z97iYkNf2+zwNIZTawER9tNwaU
I6qJR5YBLzGF2wIpa2yJywXrPB0G3qjFjAlGwGHqmXtZhqUnf/x3kabWJF7uUT1/
7cN3/B+M4NIvnVpzrwHtBzplcZcZDt7G0lq4912unY0LLgxUVk6LcE1J7v1g3+e5
nGstx90xm36VHd2EL5aNiL3Wqmx9PtnCsQUfBQ/8NK4IGlqfN4Oe6SG6KPUZVpW1
dL/7mzaIiAzeHYMliFUB8qE9XAKG1zV+kmipLV4skysEyN1wL9eoioDAxGr1xN2k
rzXiB7aN2e4JZWC67NIFbSd0dEBvowGZaj9MYX1oqcZLvZ9yBiK/pFdVvymvtAgS
cXTt46gypX5T0AgbEKwNQL1LqoZpuZ3/+8lECEnXSH5mRPA4SuNjGRCR3ptzxgFb
O30Huo5Zhlr3GR8XsNcCTFHkAuHBVM9YwFY/Balgh0gesenL11kJWCTQbVR+hMqT
HUgjNVPgumYgY3Y48Ojt+fI2H7LDYrVhkq8DveIz/l/2En3kyEyIWdSAcGEs8e21
jpI6KTmMuKgfCUcUWPYELOWRcDYs9ddE+V8VeYdMv8ny+f3n0MkqsdNydXsbR33I
W+Hx5E69somZoxBMyqlIvzg0L4983F4sBPGk5+DDqMyBMpZfEbGzQjsIE6Q3IhEm
Pk8Km466ZG5xP4PbcxLeMe7TLoo95DoSjjA2YNoq5MVDhbgUo0VVfkWi3bMez5rT
C3qdsySy/5T+tDgi+yWOZSqOHMLmKfOF9oEl9XmMFi48f7aoS+gBdzjBUUF6NEKR
9QXoYhds0LqnBuNDpFWU9zUWIE+RZFJibuJEyillw5c0d4TnR0Cf9aD9npv/9rZF
ZEEwO95t1GN/M38OSk6EQ/R32kEU4x/Pi2o43skvK6ZCPp8zhGY+F6aQ7juFOXuD
w5Cv35l6TXxOmDp1fcQzviyyYdXkJiNObwx0Vqh3V9FaHyFedup88ZZZCyXUK4Qj
KwvSaESmLuXlXxQb1YZDSymYhkXu/rVdJgGaea/ZMnS5yGtp0B9TLGuy4j1rIxx4
brw842FgTC/ChXFcp+oiIs8tc+cFsVN1L9zhGYrb2yRzBYTWDi22XNUqKrCc5VjM
NNwcHqdFIsVkPrEMRNFSIvCThhNv/io6ET8/4Q8LxCUvyiRyzbP9106+eg7jXRrS
WlRDRwN+zt22pHbsmy7Dgjsnu++OomyLzte5W/P+wqICyRheTBQLOZ8BfeTyvAsa
OTRKaCt4JHqWjv+7MwNjAWRhaiy8tQSI2c8XHJHOCm9AjyEuCzr14C0OUJIgZNXA
G58O0DREXiAqN908AYFM/mnimm2XLp9vfKNyGCR89umvgw2NVjAa7A5QKHeqV2UW
ADMrjQlnm7QMOCdHCKzsuhm+z6JWugTo8VsmoPwqCjvEhPzisGiSoP0TYsl7/Fo+
6SDyqWq23hQg/ziw4K4Ix6744YwyD8EpOzbMms/m8UdNcAVd0wRHkRyc3fl+NegE
PDYN6fpRzP9ZaKHwahfiB86p3KeyaKl+nE95AWQZfGh+zTf7pjwJd0nxb9MD7Ch/
h59AE6BmHT8nzqjBws7ABHZPr1V6SrhRpNZm7TPdbqFG3XqDs4YNLAnmMZp+cJ4C
NMM2F8yQr/0Zepx4Xmy03Q1FIswaTjJiQBhQHDI/ZxSfXewOPx4uYwDVUcR9Z5x0
c8U2Ru9iwRpl+nfIHl2WSZMqM2bPtujK+YVnqhy0OYu8yrDRxKNqi5K0aqpLs3a0
itbLoU9wt2gDvb1fCMTHc9hoIUd5CfLy4shqzmDQesl+pgHz6KosLsgmcrBUeHvK
efnswojbSuAw4kRiGcDq8CsUkk5/NUmqqmRB35+UjMwETS0ulabvlK/akBtKoSXJ
LU/eOjvHDmocAkQ4AinTKOtMiubd4S3lmng4itPGKxoDxZU71jlx5B0c7oPuuu/r
B8KSFtorkTEKMO4KLLKsWTdTI3a9WBRp4ntHPAr2NS31d4CfvogFAIrz2s1K+O+e
fUWhzFYqh0GmNVyOyW0qEShguZMeDsqhoc9xcwzurS0Sch8yLQNEBg0nG2Sz/ThX
dNd3k9wfiUo2jUxBg9IZbFwviN9pzljYQ3BH0/zwvtu3JhFeficqc16WF9w009Iv
gLpead4Jp+MMwYwtqrIWMgqiaQtXjLkg0MzXs+Vp9IiZ1fGzDlriY6uAD50IM6ak
jnSKZK1W3qwPlavSd6FKuHps7gsDD6a0sPcX/5ry7yjkJhj9gQECzeCXwG4wuCaR
ew6bdAFOa0bX+igf0+gvt6VCyk5dZrISGBokQAqtNBBiPwTNYiezcufhMAJIklYB
3to+FfL2DoQNv9GALZwNP3EBk0PrHSDyMjWufEE/Mok1uvQnDvj7AiWv1R/XIRSA
RgDafgiwfPo/tq+G/XSkyfXPZLWbIOeL/HeZPwx5aS5RAtTNqWBGS8lRczvVWXG+
dTjlv75c22kXWNpq+7Nbou+oFfdvVhvsj4r0lSP66mk2da2tOVCHi2sndFQeCrZL
rNFL9vw5YQf7qGwL0UhNWXtuXOFOojZ6sF7OTDcblaZFgb6lIx6D+2vF5YFkHU6l
05f+DcYHgTFEFiLmmom0rg1SC+7QSP7slohXRC7tcgUfi/6JPKP0dw5z35w8cOC1
4OrVKatPyfwiYJj+oJ/8JbEb98Z1jbWB9U9kZ1mRhCYln0zJFsCK4XuNwM5RErMi
jz6K86Ge/ZLPwIzE5bnWGq0aaWhRLAiYhB0JNZ5OGSCgVGeRFjZtbSwOATElnoik
Ac1zrNkNCW1PY2Qar2tzeWaQq1H7wdGzbQzjjBSHqOQ324RJ0/hz4XN23i6k224d
fJT/3wOs3TBOVE0Jk+jfTDsbstJKB2Nn7uYf2x1Bib2AJ9FjCXzKRAuI863gV+G8
Hm9Ek3t1sZJ1tg4wQ3oTasWPLxi/eT7CCYn4mV8D1Pc+3bc9JSjNxfIJ7O7ElVu8
dp4M2n1P62ckvTPnlwxU5dNiwZxCPwYZdvsAlHPy7Uqhzc13qgtk8K2NmHOCjgtm
ouM4Ydgyb28FE/739ezJetvhyr4DBCxjnRE+D1B3TOFnjG5OuG+J06BQP0eF2P/p
XYDf6OocX9cumyQtLMuS4aRUIHmkYnyyJhaMYA7oPyZObGezh+F+YQRSC3sSrPpS
HzLWZCzugsjNC1i+CWLkLhB/uXg5G43kn9aVOSSSR9LxRLnxHIumHbnZh+clgGBv
L3i2nQpUA46350oqDN1n7kFnmQJ0MRX6TRgzRzWXgAjOWkssyhCNH9uCSFTF70el
1Ai8wIRUcslimuSyMYk7fbFwpCtPfCW9ZaSsqN5AOIKaHncPkX3raL1YzSYKoQyW
J6OkFpalrdaICnhszTZ5HMQAWLrgpvvZOFyLtirO4vJPlUhqUZVAdzLt4ZSNNlQr
t6ay+Xt6Mk5guKjT5l/EwIhSB4GQg7d7e0dt+c0tyGqP4I6WoWfQC0GOK0ky0ytZ
aUAmfpsFbPYHiXr2zLr4wRF1iv9U626prz8BAgTIsSFMoqra7wP0jucojyYWfdbT
Jji+p7Kugx9uL/r8SbvZpfkdA/oTabvj1Gd/At+a9LVMatShRMTx5INI6SJVXj4E
cDqa7YBDbCyzLn0vCJp3yv32RFKA1+PKeCedOhCahhL5aj2uUxYLB9aSAXylmV1P
xVfHCFflNBCoBg+bn5BXf3zrKrLEIIpjv6C4f/lFZS3oOGkfKBEVDnKUB80XrLl4
W4RJy5y5QQW3135yNA4H9awkhnKWO+9he9W4fpwqLPQe6trBXpcgJXsLVckYYmcu
gdlXExat5crwYnXcOoNdE6na4HoYS/XQd44Gvekw2cFVutoUOt6cUUMBXinjwq3G
fK9bC3beG6Zd/6HKAElQZI03v5TMzopxV4MpH3l0yo1czsHMkSGXbaPG5HbTeWNO
BGR401yny+G3cmLop0g9oQxDLVfzuzLud07S808N/Ek2g35eURVGzash7TWaBOaT
alMgXBSMHy1m1AQtJIilnyiMhUxjju3BsDMRrRyDd0FP44PZ1cvngUWbddw/MmwO
b40DvcBAQfw4Z8tshTLZE9vP/28K8jTEAMnLknSGrfGHlSj0hFa3QsSX35X9hbUk
gyPa1Ynzc44x4o1LRKlpf2I1CgpGKg4Mv8yaJOxofJJvP3ewFkxxE4iKddSAxG3s
jksju2gqdp/MzLpR2M9D7K3XnhMa3C5Mqv8H+oEBx9senigF32/tF4vPc1ntxENJ
ULcqyR35Ynwj54RZcOa0dhA3NPfp3172FQLzj5glbIE5o5oIj62DY3VVAOApym0g
5vs90GtvPhkh+nz0Q+H81xrnhhPr2i9Z27Mr/MH50ZMH2B52dHJayCl3ge1o8eQ4
koOzwMdbEoM5IdVrzZetD5RSZiYw0mhn9HmY/bCP6nDEo03Er5TgYhS9jIwu+bXV
7hoBYKmSUJSWJBRKkHQB6PlSKzGGqCpBlMymk8KjxCG4XPD2BktVberWt86Oz9NQ
K9QudIV3jRfA2X3isqhEVz1b+nks0EFSnsKsezFp7B3ybbcMSlEaAYLvuVz2l8xi
HRYhGmoplifqa2DLf+pwXtuwl6ZTWw5sI4xDidMZBNlaxOAUtX8NUGwBVfjPfy2o
DQMy7DelVHJsVq22dxRMV+nT9J2KVtFMRw+GI16y/c0uXjmGGwRKiu8OkZZTWCk9
NfywYIAYbVbrEcCvtNkQ0BBvkMzxQRynCPo55Hwf9vQX8U2RjZNMzj35Ae0iRn5/
WIFPAwzeH8sxFXE6cwkUYBvCOE5IVMsIIAm5uIefkYBWxKO26ZPANhfbIy64M9QL
fKz+Tedoa/Z+NaeHpN6vriuVnuiBIdVuE1k4G3Y70CO7cNJbfZjHNOcFATtJCqum
dOkwHlWjmL2sxQ4z6IpTzzPhKGgaPjsmso1IOL0sF4KdA64rRpxqstDT4OCxsbRt
DA1NKa0+wQvSP8ZE6NHuNRXQ6jeRsVLOdcTYB+EF4FoHSwkbkoR0+nE2e1m+046f
UePHn2aqE6fcolKf90ELRvOOJJe+jbkfjb7jRJxhobUlN+A8ADLwdMz0aw6EynRO
W+qxZkrF/hGLpmGtYljeebU7BHcBlDrIDGzqhkOgQExrMpNjPrwKMSBKgh04zAlC
GDTuCJhaCzKvjhTJ+tgdt0oF6Xo6xfughWSppEiP9E4Sb4cRihwsbA6gHqzQRPQZ
CfGVGA2HxT97eLfhcdww/fBhxZO/iZkc43AAclliAjOFkWckeUAFWZ2pwNSIeb9e
0DM7pbXS0lSqTQ7DVgrZIQQMw1h/E3us4xESo99PVFnCfM1gSXCdGHA5//BMOgFp
iL6gufecWMwWYqMLUmPHYhyzFP7I+C+6KmqTQv6EoocTwjzQhNDAdYrPkSkjsDjp
/IJBaVn5uWAi7p+tgEYS+SlTa8HkW11mq/3zrhQBBrHbKjCfcloLW7L08EvTN0Mh
3ozElJc9RS5NMTWv8noeHDTvY3+xsjHv1ts4KSBqJmBA93tnk+iWZShdyncdTu86
jJ/J7HeNQXhVWBhhdsCmgxqQUN0LvkPL69kZGFB1UqC144A8QED9uNP549BUQusI
y8Aa0iy0wJwqttzJHNWXEAgG4dX6i+vF8KrhohX0rI/br/berF8E8YbiOpH9UIsH
EIHluI2NW379AutW6Bc3glTbZCq81GtOCLFVZTUQ2EzaB7/IOeA4G1uMVWV0WIET
oPJDrqU22ML100075afVTuny/u5/6r+L97aLgTFDIdGPUg+RWKbpFtP4tSipuPf3
q67ReamgENNOnQvjw85XPEEKlX2JaSL052F2/77JjCcDHWpKuAP3cimWQLMq6o2s
1JD/1o/mydLLlt8BC4GhRx1CZ470t16Vjl6crcBshJPriShuwdsOSCoMsn9T76SO
yPqq5YXG4SP4O67AupFEWyhu+bOvTXLupMDw4iUXd7JihVyC7XfE9X7ZtBJPmSix
I3fkBWdC1VfjkINvWaakzB4J3kl0UFEW5MTxBflwfl+kH4w5osJ9nKCWiS6+Ph1h
objMbVd3y4AbF9IK/s/QTkAEL9LHgKw0OJKTVeK2ZHiX8CFrlojkplCoAlmkHuIF
z7gDTUXGjZCpBTDzoWrS5es73N4TVywCIc1M1yTWN9ZplKESkkGCqntTkmJlC/GG
Rpwn2sFfHbv7v7o3lgm796cO1woWQbm1KkpxsUcCuiHQLDtFE7nfPYMkz7wEvOOE
FjMuxP+0rxHLn/7a8DIS5OHD5xvL3EUElgNw4DrKrigVWt/3zmpKWbGGkvbf2uGg
WiOCSrOoSWF72NeQ4Re8FQESf3k3iSO0UZaSHwsyme71DwJZRjKDtheVRvNGcUO8
TnmK65bDwUqSQKSyhFJrU4ZXs2ea2xliVl9MSnswKPjEJrTbDYpnZhu5GSsbUoqX
R9zW8XICVuT3TChIh7Jg5EYHAe4ax3GQH2XabcwpWCdI2ISHvXy8bc90LA9DhCHp
0iS3jBMCZDnNEpGuGn6As0DzObs9z6JRtP3h2WtGglnnr8RsopF8IEKXU/l1KoeC
BX/sCS4eh5UWvlXsqmh8l+osY47iS35d1gsrPWnB86Efj6PBWefT5NWCyE84W8fj
5zcRxP1fH0uED7xm1WLC0jMY5QZZ59Q54uevGCCgMLB2jiz8w79IbGh5Tml4IGgr
A/y3IKeVamjOu7OL48ABKR5gxi+LMv/1IYgOmPY5MSjIRi+vbLNHWaZWMD1zuL8n
GAYEpPRyYqJ8QpyAgz36PS4uWYOEmAYIfwIeuEHH4YXx5mMVZVTLsDWq1X0mYOF6
gkfBP/npYMAMjHlSujQ2U257DjxveTBUdM0/iwEMDFUWDn64WFezVIVNVdXd/b9F
cC7p2YdyH33C2wAVpRksjCZ1Axlq51EU9bZqkNpP6VZwflG0mQmDLzrWigYw8K/6
ZV1fmg4Xm6TFxkqOkWeDCy8xTnF3s3ycOJc2odckAH4DfUHK71ntuMIEw0GOvkHY
tpzVhZf3BxZD9bFSnj/DLEEGPpdye7R3pn8LIC6HCGAfhpscwfANuEdIPymy2xcy
2SPxCr92yz6J6Wle28AEc9PSBQABan4RsZfIpSjj17Vyr30YWtZoa/TIJwOY1S/n
oL5EP//jpRfmUqvOMWfyZWfS77Px1Ty++wzeDfNVRca1ypPrPsb5EsM6rhpvhpfP
V0IYTTS1P9cWQ2c//rtc2144CMHzb9AfdYt+SKbyfC41o9GnwfHL+GyCiJ0w8rYk
zRJt2GxR+HsecqpKCWfqx56ngYI7CMzgkXYkE3PCk3ofIKle1n+I/so+/VRHEqa1
eQznBLi9Lxe97GP5RBke21UixPyl5Hl4WxnsSHzuSSfgoFE/RCsE6ccIVYYZGoUL
/tqPI1a+Tuw7APJMtJ3DB5+q5O4n6RoIBW8ZeCZQ8EcqU7cWLeTH475Lvk5DKukA
54SJxoHladVYV+sRHx4wjTGqgbqAqxpSBL0VjEgKLRhWQYBiF28usFn+t5i1UdxL
whwOeC5y1cNmnyKJvYTMwggHJ3ePsW7jVfl4TYsedk08v/QvWWEMx50bSoo6CYIQ
A0KVAuVOiIMyFehW1egb+UePu3TgfIeAdlp3KYKkuFM97jbKom0Sm/fosQqHA/Ig
YSj9Selnx7xTAHfjqVegx+sg11cMV7fKUvAGo2hYv814EGdP9OnigO3xW+oe0D9Q
oNQV8HjXuaFVVWYt6qVeRbdDXEsBvCjF/36IO2glEATJYkyXxMrIG2v+veqGZA31
Lw+H9sQ2wA9v66YnLjesHdzxh0kzat/ZCxOJQ8gWKlZPngb/kMNGcxInyLACC7Wk
q6e6Bm9W2/k+G8y8Ow6jawIZHBrbwCB+iEeBeRVVO9qJ3SQisav5w4nJPAqiT3CI
0XO4hJqdRCcQFH5Xje3G4rZ8CjFb9TsOk8cRX40Uz1OnQo7h2arPy0ib65w6xqPa
NUHz37KZl9E6dy4kMF4PpwO89hfG3aYJmNZI4g0PPBhe8u5UjMGJlUf4Kn2jh2fK
3DChdkOHD2G5DD/yk0aJXqrH4g6ZF8lPHE7Wu62PD3QIYX8CRhEGoTT//VIOE/dy
HzlOfG1C61NbM3yytVHXUYcR6AhJqr12gIWTQKxppWYVP+s+5Otdd59jwAGWs9MN
MvwlDTAJw7ytpSC7QFOx00xIeUxDbximFn2foS/dB6LZWVUN3pm6scfz1lIkZyBb
Q93wq0lGO+GhKsnP1Gg+UNvbDLz9tueMv25ESaQoU/Z1VlsMJaiD2qrdMWJRzToB
UxlOOHf2ajFtRDeyWD/x7RK1lrKCUhHj6SgISI/zIqhdmye2z2kQFci/aWY5g3YM
9SNttK3d2Or0e2eJKT8JcgOFDHLrq9vaTeHQrPisnY3rEWpFxNV/phjyfsi0pCpk
c6SdMVifRUGtTXrkYsAQr1tkK8MdKNkh1KV7vcMlE2QQHOrJwa39m39jUA6ZFy//
FvsN0fsIyC14gIl9jB4Z2CWlilx64bLuRj1gL7mI10xC8Pfc/x+ZvCba+wCpNB0p
4sg0XSfJgvAprQbHKOeZFu9iOqT2OGURkwN99f47Md7tNb7IQReH57In/HKfF86P
Ix1Bmz5R0RtdRmBsMgSI4aumEgX6X+uGePAVwXRvXlWmVBkREHhqu3a1Q1+lyqd3
jvCgPhzTg95yFhhGiccVEmxTHwyQPQYDPfPOaQd8PTcM6B1+9S4Fb4INZyow2zR9
XA9SsmPsuxky5bOB/BmqmqRgriMNPB8XDp9hYwxkrFs0UqDl2wIXTBp3lhxGBcM/
f05nVsWZeUwiIkav1OFfH8RdZc7DTPOg+c9lMUilVGC2Rog1Bv7cwodw+byfwvpq
tMg3cGoI0/Ad79nGhbONmg5igU+BOC4LHG8KPpdNryZ34b4GGGcHlayzPTumY86b
u835qMoDPuo1qx8Eqw0We579UuzvswUl/+R4wQ0S/dXVfoneViNdcSurQdHEYcQ9
xOJT/fZVodvyBqHDxSnSntGgxbrIuollEoTV0tjk38NLSHkzeJOvviAidgv5iXHE
PYAKQZwZYbXSBaKGHbuAZGWIFte7Zn4MuTFPDV2uIDWCb6zogP1JQZOrrjpfE43C
jmLP6hfaIVgNNj5H/MUGY0LzLpYlUZX8m4WqXsQSm3P4kxr7/lI56rk3Uu6t5n9X
u5vov37sU/3GXs/psXpKBjYK8TJRX0YFXZw9MPe+RPgjtfI423JcbiVB/esLveTl
/um+fCa1zY5OuNGvjBl65n99ZOQOVmO0wAte93n7j7ivm88eguuDtSPGKOuxmAh1
OI85+iUb4W22OuI7Kl87DCvmdLo38eRas1s9qiFl7yxG4xr8FO70CX7nOf/0cux8
h3g1InYaU4Jc6l3GnPy0/Yce3mnNe9E1f5+QV/WFRNANnk3GUCOPAyh/E3ImgUln
YAA9J0IiOwjTOlIuzmR6oySxqlsfsA8AkRj85XA1xR/pR2AuDKEcr9eOOwrMX8Zf
MLFCo99GWjQ8Ftsuusmb5diSAEo8ESBQf3pBz0B+XezB/6J0gX/rPNDDFQTJhkG6
CSVKoFA7HfzGTskD4pTEaF+n6Eq0G4oS87Q5OXHl15Fbg8vbVjlEZLyUYXO7eZ/8
RHmR5MPG5EST4eGgpyyoKb4DJxI+41mlSkrgvXQDMHlBbd79N/eOvPSO1atD4vUq
Re3EvBMCEDIaIVuXwsuq2fCh8xyWrE/MVfGqjPkUOWsnQpAvOuHHxARg3QpArQ9q
mGDFPLYjMO72Rqd55qSZqQ0CsFx1qL84glAlCgyAVO/a3WA450R1oqR1MTnJxwug
SuUAo+kAXa8oUC0E3WfzePmjfW6WQOMVGjroKLt6OIAh4tLtbZE15K3Ktk3aVmiv
amcstEW1UvN250659nU8h13HP/f3TcWAQsOHcGhswEhLvJnkK09dAtppk6n2qpmJ
BrqxwaNGEvND6GBdJkC6ghlTNAihpl3lhpgGltLVyv4hL64NOJTCJdqfW/4lE4nJ
BxNiP2/2qzwm9kGlFFU3beCDlubP80O3qf2ROMndbfPM1soF06Zy/MIJSIigEZ4a
6aGcl9R6KdDgiYjjki1UUmNjh4Dz4LEqED0c0g+2ZdjSmeurHggUvPZ7dNAUIXk1
K4me+/gj4EzdO/KrgREwRkczjdf4GOZPZJeEDV/KPK22F4UfvKfZdGA7Xhjtezs1
SFPKsPXxLpzuENg5Ue7D1CKI+S0ZxbgvvqeHMiL+1lWi6atPbW2IN+38NjUxJqtw
2y70wYH0UgllDoij47aUAHj4Yh5QtQl9J5Sd5+BKFdwNBR0HrC4hmU6Qi0/RKcm7
LYbOt4Nq/kpBQKFMGqPWRf/XEnBoVHtoLj2g24sSTzLidNHwpooJfgdY2E+1pySc
bniQGAWzHt8lxNXT42n6F9+glo7JGLgLuy7ov8MTFmwWzwRJCYS9wvhUQT7y6iES
mpwG00T5eF4211m9yTpRVg62G1RDUhSzIfHvcQOKkeepJR6pZfUt8r6JC3kIxybs
jwtPMr+TvGWwCLQgHXEbX45A/d2skiTJsAe2iCTmuE0h5gd1HsUEERcrSg4SSSdc
`pragma protect end_protected
