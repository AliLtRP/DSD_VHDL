// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GQeegqwedv3PxrowaacNn/ijK/1WqTU7m/vzEjYDasQ/jXMQCqlIFiCWHpKTsM42
e/qkWT1hWggEycK91Kr8anpIrcjzbyyEay7ugnog4zGXCkLi3TrEzwMvTgyBPWOm
FXZAiMRLz6exAZ7jrsyxbsE0tXvV+nfTtSecFSe2794=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19888)
yaMbqaJOU80Y2BAh8qod75/JoH5LEAKSsFfTpVrTTGVIJH2SCWMymPsuL4ATB8uB
+9NcD/GFstpsbitZIwQRuepEdx/R7bhB1lX0WnQNGl1wCnvjecCaSWt4C+omWVaK
Km4FvJJmP+E6Ic3IvdEFXKbCDufolFjh1/Huh/5G5ErENdQqjVlFBlPcmab/Y0aj
/Jhpy1/hJ8FRk+0BJFW3HJn3rLqy/I0rn6TNu9l38zbBidZ6MXuWLniiDRFOgt6i
7el6BPHh+SGaham+ddyH4xCr0XW6qLuYs8H4RnMdWj9LWcJla4ixeMUUE+2PntV6
mXWqZrGmchPBJK8LZRcAwNlI3W/XOf0K/6KHI9DFWh6FvMyG96c+j/RuvaULcBdW
Y02lChA6yDOr9lX0485WagfoQFk+4IVXblP8kfRpswltdMfgea15x2AzvT3PEQdJ
iLkAHGOpJ1SAdBTWDGzAUK7qhp+gYBXRTNs0pDRmnNdpVyH4VYX3PxkigPtB7KIo
xbx8WZshaqf92lAVn3iyCiOfXNDbSLYs3GUYHQWiF1LGRVtCrAK6eEYaOPAL42WM
VepM14mV4TYrVWYQ7FIEA6WPRyjGJDLkwsz1SQK8Toowuf7DD0SZlbELEyIeO42C
jWz5/4qC16kDM51Nin1f4vGrwCSDfbM8Y907hpcXjmxuuGBopzKJMQPSA9a9HUEq
n7fn5XEsqN/vNXCYpJ4uo8zP9+0U4xRTTQxdpIAazlzVaNNzxdp0wLJW9rTbuydI
09LWHkSKDq7smOtxPiJ4x3KfkbOicbzEMqRD/jGX4qzJGYxwfsDVD5p0S/xKtxZU
E4gyA3QJgvEyWmpd/Aw0Mm3pTJxPBdPkCZe1NVdDGq3fmsqOp1mTN6bSXp8Skf9+
Ndd0sXk3gm7YVwbO5RPpnvVY+mn67AkzRi2dWMfqHQoyY/EcICgeASSkQBTIHTb+
HcHG8VH5Y/s5IisLGZjqhPBCxaUtDTuNKzB2BUrJLw35g3uU33STsFbx3FipPaY7
Qey+Fp+npgJyXCEilWUlg9253vVZiXnM6WrKgAQVWmZRCWUehoumWWFx9bzdh2dj
rxwdF2zaO9AHLiJ6xczKOCKeONKpjhgvDnjVD6iDKKGgADGfMEgqg6IGNviRakvW
YA2VeuM6KBEN9H4Ap2fzsu0DZnluPDPeBDxuZwBUfxJIpLUkPyoQy+05YOjLoNOQ
goobjACGqwT5oE9MPspXYGCk6lPORG0G1nSeE6syI4OFvCMLsMwsF/6YylADEbva
cSqHE4zkUWgiEFOaOG0+z5RrW4niwlFgz7zIUnNKkjK0bPQWHDhBhrlq3f0oFqcU
dJ5CmmqufiLEUW5L5t2kHr9CEDMSWmNUgAVxOSeQlVagPu2ofVvM0gMYBgNHFEal
p5ew2zRehFsKun5mc4I02BeBEanz+3u48SvUgVyx/L3nAv6/h0gVaxV4VTUa+sbn
Z44aoRz48W278QFiz34jtFpu4LJrnp+Im21me4XBVQMKG1q+SXZSfTW+n3n5HZaP
RiC/0NY/XBO/D4xWDjV4fjl/G9i/iC917Hziyor1Fk5cXq02PM1aWDLGocuOwayL
59xWQYrv/Sf8TGoQbRjdLeJmHzhNKrZTw4zgvVp8qyvdkmBUDow8VSeqjVAUVBic
kohvXxCgY7lXVjunLgY0N/x/IJbQaeq3ZEPzq6hD95GETBYPtS/d2WvtN00FtE1D
KxeSnhBMmT77Vv/2qdegsztt/6bPAnsy+71b3bj0i+HsrMUnYzf5QebWXLyLA/M/
zOz+hDTo2y3FCc/mjKX3BI0ymfYFthZbeV1iz/c9xqvKMMu9TN6BfaXFEbCB6fPh
8mGSQNXCNLKUAe7+ygnQXEfbpL464i7fM0dbmXss/ml1XNj1FM90VuuWFVIoYWKI
dFqfodlc7q3y4HX/4Nz5A2DADz8iFp3L/8qK/VRuuJvLdD8KClDjIcdtHbvgkN8D
e0AaCzvvvaULb/axgCZgrYvbfRm6DTvkaCPxKYzBVL8k1KulGRPuJjAKF84tN/Bf
aGTxD8y6b+/weAiagW3pe7x+S6MjYn8S5ZXDeqjMMH+KQzuwrmi7IxhVRIeNF7Ql
ZqRMtSGRkO3DNGiSBdYlmgfE/9CsC5dw4jQdL8rXPhMaha+yRHREdKCJwhyJuloF
y/1vXyY1ZDoD7VGSX2zxnauZoUaxdy8oKnYCchJDV2sbroUNYyBB7+ViERjbrxmp
Hht2EweqEgLKmTUqmKdZ/Ua6SnTmj1Hbkd55SCg26Ln+k72V4hpGLA0uv9mNgF6J
F45ySwxPR37qMYNqGYSJ6HfRdQfbfC311OvEKFs5xT+nHOZbFqcL9VLUa24cCzrb
XQBMZDVFDVL+UClvN6Q6YRkt7EKpWtzeMeZYqLubMjUULTfEXDuXFiaEAlRCKh+t
LdJc79nuCgJvoOFh8VKc8ZvsfwEZIHZ+sp3gcLHQYGlE5Fv0yI+hbJzqnZqhvIFm
jpYDw05p8vRa4aqct4nhdN2V5SObWfjprpGQTEpdEDflfyFzI6V1adlNLBGKB+/2
AdwRMJnQWyrYAb5gOkNIZ1YFj2dPziS2SbiWv8T4ljPIW8xz3J8QbUSJho5Pdya1
bJb5UCd4Ia2+Bm1tNNjX+DgXHAsmAPOobYJeZyxvXnS8cpdPklZhEOE7S0YIvpO6
G8DwKpOUfOWBR1ehsnkDH0+05wG3ARq5rGzWiulclg5xdUugoMMR5U8QOg4GRelT
lEOgpeb/cgfS1GXEa0Y6E8vzCJhmRKE8Bw/vetjPl8FIx8Tq1x4m+jUZ+AbVvTyz
YqylgFYBgYm3ktvBBYx8NmbV5531JkrpwV0okBU8cVdaX0RJSeNvyk5DyLhAa6KZ
qbz4dHC0WEpzW6UHqOIwXQZu+4R6yzyW4ag6naU9EawD39bLjESO9KAGg0mTm/rS
9RtZi8tCtDfjM7Cf7pw5UKGoglXqV5S661VBi1vIhl4AHMvrKx9S/BkkmorND086
gdy4kVs62P4Fi8mbkMBNLusV8F4iBkU17uGfD6lcXnIZqpjER+XLPd/Oed8iM1Is
PBT86ozcYVWxFaODvp+2kKE6TMfYrRaE/gK1j5fcvROKz9MB+v/yLM7vOHrXriQJ
O+GJNzFyKiMHHUC3dIrKL5gcxBL14cnRc3djEgI5xtc+JODzdlAl2ovRB6DSa2Vg
R/F2TVvgILP69EW+soJdm8emOJSY6BXzsNIqbjj9iYsJK0Nt9rjhiuIM5A25UmFA
dedx6RQ70nuw/dra4qsSJOisFMLOMTvnCaD0MewgegbhVhglVUyuyQN85F6iGtae
AXyv74BP2rsAQmM5DDIz+S5CkeSrhdrZrb7VwfNDbH/Nu1b0V9WrWtsehnCMrT3C
vYZrfSGew8npCk9VRejjt3Un3L2MALwBE6oZWRx5a/vdkmFJit/W+Tf0s5LMu4yj
aRfv5sCtLpi92cRLdHKYYZGCWDgUSZpU3hYrKoQRpt3B9IezUZu0OKCUApgHl8cW
lKypUU9nbMj/MMIRJ/MOee62/jUpA4g68nD+m5p61j+qg0cJ4O1PG3WcZZFa98Du
M+hOkVDoo066cWj8tv/A0DEqrsvNX9qG8q/TT/Ent3DYRvgsmseKF1nr/rGubq26
6QtUjlv6VK9/g5s2KKVZojWBYWOjjMgFpbP40jhSD475ckm8mcyGuZBizLA096D8
0h5Vbw7btEesAeIncvwEbIZSg2KNA6tksjkwnbfbNRt33PQxd7FiW85y0lqN+JtV
122sjFZDmoG4ZS0LWyE59u2ljo3drPRjo4jcwlxxZgob2RRVuVDmKVY4xh7pZkq/
nRqpdVT+eqOPaupM1e+wHkG5Hob+ZqUznDBTrtQDHI8MyhmVc6qkVaga/akgqwHR
18/f4iAfHvMrkS96hXCN2bcXKB9NfEVa+/UpbVFWwu9pwfKt6k+wKKUi52gI3B6+
yiVdDfBEHSHXyv6YZgkwqEnq9feuqFMlzFd7E+YW6gIS8Q55NJtUBxavy9EyOUdg
87FY7f/lK86IsghnuK2rUo8nvSHpFGrCXVrJXh6zdqIq4QKjrrB3aWO5OhjnkGou
tAskViPluBj4AInKeWIOV0ni8uSJSvh/GSIgOUQ9KyQJvLwZfC7kusYC0/GYmRU6
Nm9f2MNNZiZJTTRTlQeTB8V8dd7WGY8Oh9tt1/r43ll5HDKyAMYw6Y72204zWd0L
wA/UKJbaDEE4pD5ZS1ONgHVl7T/lUJEB+kG7VDOy4nn8ZWRIr3i2dEXyBvqEn4Q1
EeseOF/ggZuFvxNJF4S0Zu7c9NeRRBJhXgiv5J6jNqffugil9t8gh2r7dUY0mZW6
gDSgIhPtC1clo5rpWK7/OIPW3OjSQ1VDjsVT7ujfKIrbKvMDQZHUVUQyLPzrVvcm
oWPQ46VHsddWHtCb9wpBbx0cVHQrrqTXjkvLrDVrf3j0b5MDqguSH0A26XXp2Ivl
xpMx39wwN8jF8+B9EuqLMLnhdT9ILCGcvTqTffgpIy6xKJvpuYTwn49rFbyyBH61
3Imnz1LcvPZ9UmXvEA1qoiatu8dNBaBJJdKtiLYxwOnRcx6yDWy6Iaa50zWoHPE0
L2JZm/Bg8owiKk2EGi01dug7YiiivZDdtaZ4Z/Kj6kqEYpfd02Z1CgOmFYJSzW4X
k5tq2mfGleWu/e1vjHejmawrZ98sC+jnA86Zjj+MN4PymHGteOMEg2J6gLBL+bAU
wNb9nZlkKYikrMC/a6dobG6WKBZZ4gGgo8smedhhK+BOyLUWiMUyyCfVkgQgPniH
tNjE5O3L4oKJ4VNoTGJXNZYaSAVm12lCjzSUt/FPUP5TXDtzgiZHB4wB6/BFg3Pd
T87+w0c4BzWLoFunLWi/3/KMp00czVwq6VlkskR6Me4hejUFOo27wlm6BlzTjXFv
7thMeHA1thOBWONFhAAVnJsCXoH3KSzg/MIEabmjdRnj/Ecz/t5CoB1SlrIUhBOG
Gd/ptRC9jNpxQPOu/n3XZwBeeRFO5hgjnuvMfkSe2g0bN12hfgomdkTuWE660bNw
04T4iI5Jk1tWa1vt7mggyEFcqj52llGjgM+fzN+VZ/7vkZrOKlrCQGsxKgR2DOoZ
fekXwgQICkexpCYtdTCpE1D/+4MACysKWvxkNj0jMFY3zKpEq3B/F7qdCIPTLGId
IoC0QxwBbwbhznfolSNpdk0+Rea6/KFS7ASsez3lYXq3ap66dz0DpyPFNnwuotaJ
EewoNvSQbtvu8LidQ4oy2VrIu5l/+B5dI2qBv97vK7y8YuyIQnE9RdAN9/fRCbFv
7MDtaIycWnR4e69HH4x7hgan9xcHeTWb1l65RvkjP3up6dZc7w7/pORc3isMPsAA
i4g/xHGfkUSRHOaSdoGeb1XjRSUjt36BjoKy70f1dvt2ecxkCrBgI099bKPqZotF
uuH73X1J7Wt6XC1C0CbBKQ6PdgeM7Ft+p8P3aV8FaziPRsLD0Tx4+IN0dOXQoAwZ
+BlJvOV1yHOVEDfxtbKFHDXdfelW1WhcnrTfK3Fnwo3imGVMoMrcOvZisQ6Nz5Zy
jqcd9aT3saSfFuWTEeejMMHAXyOVV57LGwZb/DApsbO6K2ENzWF/NF50mT2Gqr3b
/53ERwxDkuUNyxz21MV/xtkx+clhu8GhEbFsYW4aviwhcpsfDhNF5M6knpQ8/vB1
AVxI+MVQc/CJUYfWFU1inziEdk1Wc8jLirT0+TKyqPPbJZe53cXZqib9rvEiqOrR
y8uozNXuskHmjwEHtwfuO8GzTT9veNUni5skrgZW01CCx1jfMingTolTHfSg9FCG
YJA+WZuq3mug4fDM+49wSzE+nsIJMpClmSzX5CdabOsOM4xbepWuDoAwGqYm1CdH
GAPThrB/X8G8u2xLLqMpDX6LUQHFhQ/+APEapw4cCjf8tj0FhjHspG0Uj/JV7gCv
yCgkBNvKZDZHDWsJPN3KICSKEtTYyxvnTqGysqJ8t+ujsDBn8bPZrRUayNDNwHN3
dbOxP8cAoyyxACnBRl5Uf/GTV1pFIXOyouQ+HZBV+nFhta8XfL9CY5pVJNrt3fM6
E1Rjmk6vEHmk7H56hnWx5gAA7HybRVPzQl2DAigtw8X4QdHkgQWrGNCpdl+3pNXd
nhoGptUYT1ZYb3sSA8jLx9VSSvcdrN4B+RbTw0qGobOrZXl1a1MYpPa9aRrEljqi
/tFHljhXkL8LqF14H5hUpQc/XdWWKYtrbxy1CtXTDpU3YBjnoJ0ZIjXFNObQQq+1
DiEm705DZYDdBhxmw0JjHf/k0fGPX59y2HQcX+7M1C0Sbdpotsn6rIZL8YrOnZtP
tXfUtpPhnDqPUscKLsEj5ARIz6wOagYSXlCUrykP4mDTpb+n/MCipkU8E5U7G4Hy
mCqhdmtcEDOMT4t4noEMymcfOohJ3teCxd/0gUXpMyoNjegID/JXGYwQLX0Cnhg+
bsPOnsJT0Vna+H9iqCfwvCyuv26dqaFzupSEOGHSlUD6+DW7wPuIHq9cROUNjdcE
8EoVTa5X/WUD6Cv1UJAg9NRBN5ZkXtGw7h1gcGxaVX+ZABvbignSyt5ixy7DE+Cm
mobcMJc3E7wGSTbj23cDN2+WalXkClR4Js4CZ3d+BVpdu262386oFt51RjpvurYT
tt7T4HhzeYmO6DBi4gsRX1JG25yL1cukX11qj2D5HwTxNQ4NnfOSMR2p6kooW3Ju
gj/noo8vuCOHEw+a+ulkfQa8Q5rsBVkxj9ta6RQR3y65ueMIv5h/+v6xQf60ASjV
XK7YZeonFTk5y+i2GFygH6CyX1TcXWJydFuwqgu4zcNXTYlrSDX/l5W0nlt47pWi
aRS2Nppe8e3s9ZPY/SRQGsQOXR2FT1BXVVoP/ST0X6wSRV1QI7MAC9dy8I2K4OpX
xPfyvJKGk5tEQWXvcfMm5fpwxxGRCcJSYS/QEKX9Oz4DdN+s1xBB5YCFmsKggA30
y3aFjaPIPYmGXPJDaYugnujQWZRsM5l4ypuU1guClc9r6NCZHwWnhKcirWPZseKv
UpyDEVgqkgIs9iLMnqN9T88a6z5VkWEkNQ9WQxLUzcTvQIibLcixMAbuWzVV8XE6
vnSZJ5e9jIedkQQszo5tsFiOahYQ9VwVFfTm8HWZXk5uU7GDikKlpFX6IpifKpDA
Jd3VI8bpUex1YpjkKWT+ASpzWF9ubLHE6mJlwlAIKyoDJfhDJBiWoea/u4wXrgsP
u7FAINqb7e9fwHLc3lI68nk4KQOWcmb1D/Bm4NyHE695kKnMsxIoO7q5zVPwsrAV
qIOWZ9vmPYe6iIQz6o761ZxoiRJ7XP3pBK9ZAEzpvXxTLNF7JnkIFcr/J+92MlpZ
paYsj7myloA7mJ0Lx3sJESCXsyLrTazxDGGWmHtAP3fZ/9TH+wh7LjrF60NdHQZf
j7hYHsgVRFbJ4QQ2jmNTFqY5iYgyCQS97iLHaKtrlZYtEu6cy3BUYYXCyHbvTQ4I
wPy692zPAoHmv/v02wkf8Tiqfh1UZhJON+JEUim+8sjU/JpPcc2HVZaqzoSL+S87
7SkBa00zgFq5aQzQ7NVs9aC6wKBDZQHFKQL66h+iEiBxG8jDOJ9rS3ZxJ/JGfOr2
nlUZ7F2kEicNttUL45jPkcyv0VsMA39sirs2CZBGJMunWgE68KvOqzv2TLTIEAWz
DSmJFUXaMkQzRnZ/MV2btwAQtVL+VJumrGwV+e4dDLfYZeuFX0QibNKRl/4Hed/2
j4RwLm9btFerPCRc6d7dWJlTDKGDFvAAPO0fatR84X9g98Dize/9L572pU4oajDj
qxXAOvP+xKyQd0qGtT39KJ6niBNBjayHUvYXHBSPqu4RxugCHYo0YUe0f8PNngdt
O7G0B9rGHDEgh+aPa80TComMpcNhKQXKz2ReBisAglv7YSN52kcd6Fyp1DwQQBvX
T37XS4ZBfRuwihnA/foCWIVLdpitiJiOeuiCNjaDDyGkkRlK5kRnMfPoFRkPhpDe
VzreP62gPq9Wn/b9Lx8cSwDHeyvgVbwX6rRpQlNwxPP+O69zWhNf8GkYd9iTdK1W
VgonaapJ1+7X+pnwQwnsNe9wYtjf88pEdwioKorL28pdEMmKD5DzR16/H8OtO9M/
riajxxgyVm9wJwJz9hHZx4RTEYzH/CroZgKfn7t+z92Da+2zNk+1R1b2qMRRBIO2
sgJIN4Bw2CA0g+6Kb4bXXBP+3HzyGkHwa8x2yh5iuTmgu0AgUKIIOcrHEC4izwWm
OAM77G+xgyRVDw0i2qtr3mfnXB686tClZM5wouMArzfNXOZojdicou1yc53cfRaS
SF1rohEx6Z6aVKkpDsZzg5tTZGQ9UlELwxk9tqza92PS4H+qH81KV+hOF4dHeyGZ
QnZ/2zgSF3wftvLt5ID3apqPapER+YZG7A1Blf3Y7Vrh6D/QcWFGtEBbDO6hixYy
mkHYrg2Uedgk0vb+d51S/mr4eiqegUm9wOUo8k94CFH5bV9GgPQozOGwURjhZ+lU
K5h7UcNZQmFKxEujaDhbW2lmXg0fSzfKJlVE8JV4lh0Z40FwQrgUvwr+wynUfGFx
Ua3yPSvbyaRJG4+sk+vti+gipc3EVADI3u7LEHSNBTua1rWYmqxQc59GbutfbzXb
VAvLFBtZxvLeUJsW28UVneqwXG0Eg8FlkW9qI7kzc4cXkyqYoPtLbNrVoCDPuEah
mJWtZo6DQggpEtB6gE6M3Ipv+n0CMgkpQRYh4qWQJZvOq3WK5wXOR7W8mDkfsUO2
dl1ie0gIZ5or7z8mVrSx6oO0cBS3h0+GS4dQjDVUXKs3WxPMRvGBDxe3DiUTdDo4
f7Hh3qelTFmZC2vBa6D59gcZ2+TmuTiChHAtfmemoZNTn+93390ajjNarWHYfhdE
KWGkQXYWm8mSgzBn5RccBm6XqQiZPNl+bCmC+jwPiPL1nPsTe6tv3O+guN6wRx4j
XmX+qaS27Jp5UurO/MB2rTXPirF/0Z4AlnTT7o/Me1++iOh0t0KyRL4qSWJQN04f
JVNg4IqaOtj+WjCPMb3MtvKXClxHDxEuFl8Hrt6BuOzHanIVSVkP9h8ZZUPc/oNY
0hwJpFrfDBAevoVwTkFDhJ5GUwghsoHsWoI+qZjw4sBalSdkrK5V6jWJ7EHixXV8
uXaBfQWyEd2abP9GLlVP+px7JC7w3yJqnzRZbKZdhyKWK8/XX6MH/IsLPtdRmwsg
6KNwphF394w4ObuTa+wwGZ9K2G555zB5nZ40PoVnWrFW0nzRciP9ykqR5V7dqTgf
uTefZyBcn/rdfRxEpc6R19PYpNPTV68NudxgA+ukaUSBP7TcAAhmDl5h+UYhKtyl
ZRLNVvpYY/WkWX4JCYa2QYuRhRmAZMMRfB7i2V1eg37hNrxmX5zhAUF8CIzCZsUz
IxQtqVBychm50zM+8v89AT6kWV0xXgSxAUM1YRUfFR4/rzTmOR9seEfJmt1SnVT2
IpsfKSLwAxkqd7lKqfdWUC5AA06XfU6oKqDCTRlngCHU15wJgvb1AG+QvdQYAA5k
Ri5YAoPvO386fBtvNqA1Eeg8Zpn8TbI6D5Qdp1SU2x/EM3XmiawVR+jKd1UQVA9L
yc0smC0B5I/H/jbe5JrbFPXkvTJFIO3zlr/hl22dkPbDo/fFNAlJHCNPviBm0WrA
ndyQw1iWDopD0HRZuYF1ybAAYlBYtk1FJS2rv/Ek1DJRV3IDp3BppOicYS+JrxWB
4bFmEtHI9DMh+LshXEGDaHoqKQgz5qjAi8VXWwALlyswyDwdLS2ffuK+zGOMCXvA
P+Xg4PMJTLfIiQUgDj4Epbu6VUe3e+02RF1FYiCYnDR2ptpv+5efRoqC3q8PDe3Z
edbHnK4cMlgWSs3ugQ9x5Bsi+N6wIHFOh7Qvhw9NuHoPONXu8n4u6tVgNvxqO0MO
MaMeXsgvjRJWzXFkZuwGHAU83JXU07ecB3NK60jZLgTzfUDWjEbHMcuz7uqgKyuu
66BKJtr7GyxmV6yc/1DgQbrJeNmjxCCKHgfLzFp+q+azXBJtzNIo5YegZCjMeMMi
66HlpZ1MgZuNVVeFBcS3YfFZ71FSdzCFsz/A/Tu2twNi0NwqZC4ZLeUED9WJhWy3
Q5P9C5X2ZjPTgUQjGgm7uk6/jCiA4AgP8+QZRgOguOYfoGG9sauI8wSS5qUohYZ8
dI24NpoTcLwcVEjfdlSMQITohQg278r2mbMdbgWU9krYapnYyyvJKUWPJAH4XnS/
bJjkvBm4+SS5G70LqaZ7dGv9mltTqtOH+JeC3nIcTxdIEh421uAVQ31umqX7KOwE
srJnqHY6ozvQIw/AIUfxxnb1zffMUs23aZ5DeN+QXbVCORauoujPTtm3U41X26n7
Kis7baZBgDuy3pXt+mltlSI+2cWeyk21nTjql/2ZyT2SPBopf2h+yVmGTYEzBM5i
qFeekzcbaaK2BeCZewuNPDFfHsyg2xLBC9HbUBp1+OXVprVnCwK9gvtP81FUX4Ed
PXWsue1NmeErmThkHnjKImHH6ojcfTOHAbMroHzyGooOlFIXBqSGGFXHJGYvjkmB
rKQkmGqeKUhvKBClVQr9EkQdKmoWd9mf1a+e6zgEyF0Ml+Dp8VPy8NRfyLqMqjM/
GUspArmu7AbMw5N9JAdCjGumVCVwfMhqpQkrQ1UiMyWXXyaDs1rCDAFAN4OpSEt6
aPECc7UshcdzTNfykrko54xlrl0H+Hh3+kqOKjn3EwpVJnuDmaYLl9tvtGH9aUV2
OLPy8Jz6S6lPZQYGpN+YYsPxz8RkiSyBQNI0EBE+8scvEyYwHWCw6p/FnIXaw1m2
LXIksWw9SnlPTSvAzoMfjVgYEX/bXLPWMalixtRcguHtIIafkJiyc8eA/Kq2R14b
fqqlwUQN+ei/kqLwnGBxt2m5Xun+9cccmEIjtvSnLcxhVnUpxmN5FMdRtuKLLGXJ
psNaq2oigdUwbW8hz4B+S0PkXp5Ug2r7AT9W9eJf7VNXBsOIjaSD/qp5Uba8mL4S
VXIxQnmsOliD0aO0XrNzWXXv2tjGc49BhT4oUv/ba2179hpoif1roQ0Y9JSbh+BH
PLBXK6uenkk8gryJv5MoX/NkvNv+8xddC7kjTExKJ36qOcro8X/kZp1KnCGVrHia
YIKKbC/ukEsPbDD8UpXS+m8hhbgkOmZKc2rrMjYo/2Ag7jwAUg1F8XmKQltRVs8U
kdvph0jOHfN/cOVhIeFievaVu3FwkISICM54kpqtC4ofsmpMX77qGpgu/MCRj4cs
cUcXJ4ElZ0LK9wHjpyUjbcedloDfxf4+a1z/y0aN9wsn5nHA5yEOnIoNlwcLZwEH
Ww2/+jbX1kB5mMBZayoVYjiewyeJicnY/hgQM3nwFXwIwu91D0DQOCBe2ZWtv/YO
jScXzz7aRxA7wLYC8xyuZd+VMyBed2wlXpPZuemEQwgwf2pm+oaRDy8xzdCC481Y
8wp/sNSJXwEfxBPIg2eRF2fSYzgBYJLDHMtsYcVzPLu42DoPqW50NmO5kjDlQSRa
jncXyrpjTsPnC309pJMp3wDW2csNokNr+9F4QwMNlfJdRuYk37gXpxHCVoF5ying
s8V/aT/UqvNHa1ojmqZCHJP3bwbsMxAU6gylGWteDnbEbediSduGJtSJmhGOTQAb
wwAvpdMBvYTuOJqUSrDOZwU+e0/2zagJwVeN9owXQw+CKKuV/6OOpA2yd0X/LGz1
hHaXdOKliPJy8rW5ZfLA4a3wXeqtuc3IxW+2yTUkDKWvb29ImHL9BrFkizBqktK/
Y5OvSIrPc04BEKT59hwGzF9eECs2B3IPA3XSiL5q92U0Tc8esrxsy3Jw0W6uI0VG
xhssdERUmqeiOJeEmd1lyBPQ1f+OlB/xQsVYdfVOAtzNKlwNAga16xHbe1DPq0oq
sSjeKh2aDEVbswbycSRTCazW+ELxHYbImQeSEQmz2gRtC3tY079b+8qva9ncd+38
kV1rHPlryV1IDTDFZQcL/kzz6OUf479cBW9EfK3Q1JO4ZkV0SgfVI5cZPMJN9BFQ
7UdeYs3RPkagjDq4yDt5SGM8Y4oCalHURsU2AI/7Dnsps7UYZurVc+xNabfuEJZ1
S0Z32nRdDnjQrTjxN+iviS6VVxaQgtOc40lvDzIYxcRoqQa1xQ6FP9BggUo3MkyC
LIvFK2JCCxFp4ZCjv+c05ADYzrg6aMfDJeW/Cz46LXyWBQeLfKQA9mAGh+r15TvJ
vEC6vijXfuHAE+zr92aOht520/GLCGE4aOjWB45sk5yFFfsEsv4pQTks30KNngUa
nTmGmbeCHL019bCM9plNwvyudEQp9C9sknDDZITU60H6uOFToPEqmh3lOjhi8Iv8
6jq5CQTq+VjRF9dC1MjfJDeR1n8SP1SuyEw720CK9yeyxWRflbOZMF5p0ooCuySU
CjVWYS3yx/lMCjfdhbaYPeF1Wku76F+JpZfyWafJM9bBbAzotePJakWtmR1Vytxt
bN/VWgO8xQf6DW46mS8zBN7WMEzOsriB81xwqBanSkS2A83koUXh1YyIs4W3i1jY
BkFmFfZGTTlNWD160r1/Gb0aa1FMzXssbKsctQqapqMjwg3POuOz8AzRI4Ww0fV9
kwXwVnHI7MmHc7b8wjtIORDnc7T08s4gcAk1qVSjihEmBK9si4akgD9ALQDnEZZ4
e/ECpX7HtMF+CgdY1X/R4h5kIK5rqbL9Mb1dYmp0BNaHNfa4hgz+z3aaA8Xygemz
T1Cnb6krXNvpCGstO4xHKS8dSO8a28Cx1YqdNCE9B7jFG3EwvzgdqAlhDvhQxKm4
GkWe4MTuBB+8a8K09CZuCFQ0OR/ZK9L5JiHTak5pp00wVgxJGFK6/94U191YFjg2
EujqOC4Y4qurryDHQcFlbIy60NtvHd0/O/atyfWlRAbZDWGdunE/x4AaTNmxXBkT
cdB8oYQPEhfIYpLBYwv49YVjt/JwAQkqpD7exWxQyTV2P13vT6ApA/sW8Fb7IUXn
ZQsMrSLF1+XYh0w06j4YRAJrqxHQDprxkTgyzaXoKzCo8RYh+OLUXs8lVZBVkIRw
wdpgCAfzYy5Jjw0k3GVHcOEjfx5KualRQttK6WYzwF45+iS8JbAN2Lsxv96awf32
iiwW6jFuOHhZLRamNR89fdvWt7CfpkZROwuspjONDoGku7kf4JwHiroo+LkUGOIr
971zlG2muwNTOBa44w8nefIJ+1kxXctFrb5nXbDqAJ9MgJDGYUdZC7PDO/5NZIMN
R8cpxftmeBgbnI3TFd7PO0Rx8Mzj2uEsjyWtdNXmdcXUKuNvnTD9H0JcO7BYKksp
sijGbv2Q+jTMfkLJwTy0nRCQxuYPfsIKB/1qxtVaNdHH3D8y596QXNbfktE6Ai7G
8l9eB5U9a0CGrC6KwNHvPy1YjCHs8e2+mvsXhH1hT1XhUwydMwR+OIAt43bvyaoF
YdscF9KPCjNF9qgjIrqKa1yPVAKAcV3NO+WHd7zF9zGu4eSFhzxL/D5a+7/lgtKc
TDt0iefWCW3UqcZR0viLzPjczCdDrdyRF7vKVFvAyqCJ9Ioej7l4JNQMBCmS2L6p
FHus55zw4ncXP3AXz/GjSRPS/8gbdbW0R0tpdMBuwS7EoQN3wSVh8qwrDna2fmN6
+Oipe/8Z0l0OT2xYLcN1FKkcvulYIbvwV1jIl+vgJHbmCuc9pKIj7jCBKioEylWA
r3np9aDxUXiSVIPMoQbakpAQ+QL/p2qg1dBQU32BN4OhoQgJOr/v7oPO/UCM6L05
iWDKAZhd72dmFV7aks4egYAJIbz89huIP2rKO51l5y+MJvB+Rd5ywnhQRvtd+le1
/xK51F9XN29wzVZ3lQR6h1oFLYSsIbkvBFDZsWrehRbCIymVuP3EC2ZV3eTI4i/c
GSR9B3kjmfQEcvS9KdgwvwlJAlPYACwpPxMWXGE/fTchhD7ZSf/DGQAsgf68cKKZ
2eUohkwgjwAPi/CZc+kXc0V5P1jfXnuS7km3DHFYJL/nYn3Gm0iMC0v7zLAyV0Bd
tcCG8J1LgFFud7TV5lF++41X1ms3EWovcIpevu3XdODqngzcOa5zD+cRYYv4sbFW
GnoTVIzd7djcru2G54m37d9sDlkjmLwb5tmfh+NL7RDb6pMk86VjX/IrTSv8n6Fn
H4NC21F3l+HH9H82zwdovRJfNEzsOg/gy7IotehDNX3Yregliye9y0LtxrCSD7cr
ODz+nWT1z8MghxdSAa1yfkQqaUgeLFFYCPAohY1fczeiURWLyB7mFuzO+3bHowk1
DmcoR6VM4BoQNHKSDTsUs6xHGNvxV2UBYoBZ1lgcBQ6qaam1YqZ7r3R1HctppOH4
3hTdr5P/LpO4cL7Qejx5nCOZoLr12q0QIfXJG/Ym5yoLNDHF9kaG8nMEUOIzlbu/
DhnKo+GsNkXe5b7K32zaES4X5yj2lmondMnqb/w5TL6fLENGtUiHPJ7U/v0dx2Oe
PXDPpU98GBXZCyBXp04GtNINbsupaGMYD80NKTkFv/uubmnJY3h7+r6bKbD+vvZD
q9L927eod2w9O1d1g5DWdPcpMikKjNwBPiWfq0uRhqEFyxwZrxF8IZQeufALgFUk
rAf/8BMCO00SR0SjuxPQtimrbZZg4Nz+/ewBHDIPgUP9ma7ZfI/sy0QxSLtT8pjU
JTXr5lLYQ6DmqPXtjzji3K3UJsbBitbUoYat3yLKw+oLLQNuse1O+TPf2VvbEFjn
mb4WZ94fJsRB4tZPA7YgPNcsNGHHdH+OKFRQ0qXBn17Byx5BCkYuiEOWMhPWv3mx
5PWDLoz2+na1wqav9zmTHxg2kNDTouLsUtxtKRsdZRDWM6h3wGk49FAmxr634B50
nw+jygZTELwToaEVzUTt/IckZa3RTEQeaO7yCdiBtcXdRaO8tdMxvNXD5zKi0zed
utrSZJ3BkJZ4C1aaW7X/JT3Wm229b2I9tkCgCjkGN0JG6xb7XCdVW3G91054nrDd
/6ZXX5wfRlvBMShtHhL74bREDBYA0Q9b4oiMFRUgccFtvUamHYci3tnus2CruKJt
2qQUtLMlkgRLBvpIpv6F3weq3LNgNK76O2M3Kq3w370FhRXRdZn4dX28WXhB64Ce
N7n6jaYjshl1iqjbdk6LGP0otDXwB0sSAkS1g0PJ1I8HcLPsdExD5KaerR5hSAFe
mxOfTy4apdB+g49IUciGBl4Ajla10hsfSHpvzQ76lqQtri4hWPBjQ8qONaZeHrcC
sjBjmxWhQwq+uxs3zy1/nisEbnU8yzjzbMAFiaRb0+T4jIP4bGiRt+f3SeQrcr8M
bNqb4lQel/O01ACZbJbBrDJkVhTnDL5sJqQQkvXUCsHYZgqncSByUviPzYkDY4NQ
OOE6Lu+O2pKh+GiW/uaI4rDE3e7Ds4m/l31qtcM86bHSimJiWplXyh5XNjNme6B3
RRM8x9LuWJ07mOEJSXnVYPAE0znHVjonPXBiDLkCQR0IPruQTwgCp3YIorU2cuUO
sGL8B38nMjprH24nOc0Mh64RcVykNv06hV1qnM+jhjmfGjiJ/FC495vz/2lON83g
KHTcD3mCoc7BV+SLyndm4CwmbW7gx9+R2C6UR9JuIYmnS0dxFeXWNEcdyeDYjkyL
7zAzvGLNrLJ1AluXWjNprMmbUTF0W91u7lce9nNRgDRCq0l58Fj9cF3gV0ArVH+M
fv4kRcXzI3RkBLj4w+rb/HnyxYCOxaSdeu/BBzgT3z6olRWma9kD4Jr6N2TktlPB
YxUOtRNbwntqnBIXAc4goG1a93FIUwWE4an0idHXaJjSACbE+bFvCtSSLtDJZZwi
xETsRihEVvhGpjCdikkbyX9q/1046HJqf5GR1Jj5A2FRff6YYbTcGbiLjBEaO9St
R8RVdWuJaM42hxcDExR13osPc0nzP2Svn7rR5mEPDdsLiagIaE50orDTmYMEKMeO
8wcu6mQHYuNfEmP48DVRxls303WirbsaPJ7npQ20KugXQ7ZQS+jGGTg06Wb/Px54
uu2eiQGMnvbufXEd0B087/dvtmw5QyhVpgomZL9ZdMA9mGs+S0OPTPslM9pwRgkA
L30D5lYbLg5EBcj7GBhg/bmsj4RsZN56IJjLTg0z4YitepO5bvBA5CGNhV5nfNrn
kykgX/9As7O4TG0fJHMOpWQ+Ti7lPvqE4JViWn1jAya2nVT46X6tPgDYka4/osAO
a9mutYkv7QQn6ZfyX/4U/d+8miS+a7t15WmzzBiR0XUJMccSRtD8p9qy4YJrrdjA
IRss+LmndE8R4yXdBC8VKIMYfeI2LOCpge+j4f/AKcgWkd6NOFsRM9TPYv+YkVJU
qtn7xUElNLKYxTmAaRA5tu1vy8COJ4DMnCJEMshSPbAtF5twCiDfHJ2nW4YYKQAn
+9P2CYljLgND4bHItG6QL1s5onhcVTBMTU/6IHzem5Mz59mWl1HtgKwBbKpViFJh
xL6uFBE9D14ig3Q4UDcKHLl46fPN9UUaeNn4Xo8TfwaMcjAjFGWVo3jRj8LAVAWo
8BSPQ0nuBnojAjJ7qpBEgfjLtzvRCqfus9pyIwZR5MDxMCBq1giNN3PvzwO62b3J
iMNw6z2/civqmguAZukvG7rtz/Y8TCKc9jp3d6NoDDGg+GrkGjNEOlzTPNl0+ClK
TjRqOugQmEhIe261lp3R4Og7ZBFhCX083sCfz1OJKOt2kCM3+r7h6CwMDP6tMFmc
wfvHcKY4YKh7vff2muK6shDyJQ9j6QNQZCeKjJBtU1Ag29wTafj3SibF/jhIl+hd
Rzir2a/nsGxPX1n2K9NGUqiJ/1bjbFI5CEPYdZwRDvYUN28UqmsI0QgcPJPwLnio
9LBhQpLD479AaYR15fUHrSPP1ojUO9zitkzBdvAlD8BMxRSntdQhyBeOKpb/wPrt
FSHyS7D315xnqY5eA5UD//ezKJjRKR0e1mprIdfsCYQ7gLbjNMtYDQ94g9UbfmMt
NYklxN82uzwdWiEqIjMj2PIPXCvIl01ygQanzF32C8mGCAiHS1R6VcP7mNNmQ4te
+TLFvDrXXmInVMTiwqM+ZNRRQUkggJDngOVc9XvZYJWZufDHhccxOX0xEaY4YqZx
WV7DY9LO7tB9KH+7mIPGFPNBZusyFazauqflgTDvlrY0W1qzQYEy9jd5ddnH4rem
uDX7VcrEmni6QAqe2o+Z4HazUF/RdEOo8oT3TM+7WDjM4oYxsG35LsPlr+w8X6t1
hJ5KKgEhFjlU29H8m0I90HhUFE19bxtYSwgUKZhzpDuRmeTafiKbFbr07nW84JBD
rvg5XWE2K3D5iWuTNXlQ5gHrSJho/i3Uf00Qi/d0sEXI2k4/3u3vlTbGsB2KS+2R
2dNacMI53d7qvOUvBh9FGRZmyS9ckh/zpzCR90tz+wcZcFiqa9hxzpZh9NIziTdF
CYwMwP7Z1MrsxUxrqSYIG9lHFmaaQCwU8GEvQyAxFPL/9g7NBRx+KMMMM/oyR5Dt
tMa0g5De3NCLCJ9xay3kmarP6Y9OAL3vhvr/GavIkItibm20dNi/DrUv4tm0gnhY
v5GY96BwnO7uAj06F2H00rdVJ5Q2r/s0acPD1C8JBZ+l/nGiSBQ2RNBaswGHEnus
eX4lubcTxjMJwLxUlvtW8TL9doEPA+zNuBQpz6hnr7LGjEG7yTf/OFwKNAIhN23i
duoI3wtnOdYA1J71Ca91GDjhffY9JHb13j6DNI2kNbc75lH21p/ft7A42WtvUJL/
05gTocx9gvvjbYlG47BfDrtKxFO+2/w+v8IIufd5ER3fORa3VJpTMw6DMRulbd5h
SjiXQ1AP1mN/ZF++32JJEhwMwTuaZbqONy+RbLKzXe+zmns0T4/jMCLYLGt3pQIY
K4DH41GKBYZyrsXOo4DKwPTuzNth0Qbmk7U8LDjcltBsE9EuMjXiqJT3nDRqNhrE
5zYi1bW7/KDEoZsS+ispxAid8oRvESpfXZXW+PFsl1JPD7W8PQN89Pi6Q8xsSNw+
Q4SRV3j/uzW4JavsoeDhJ1ni+KVdJFA4G/KEaCjynXzmPTTal4e/bYcsSjjB7ojg
4bXvo8c4Zb+HXG7uDgZK4XefFAda04XXFKsN67XUP9tYYNKzWEptv2o7QF5/oXS/
eBgw7I+PZyefoYDYISQIHw1Etgf9RuRNy3E1EwUQqDB+UOruVhGpzXIzV9xWOhn9
sKdYuFrR0N0XlgHcgDA//u1mfmw9nxqfg+woiFpofwd0XLU+VntPK2I+kDAU0ytP
QEiKPbLe0V2AE0x9h28sVSGEkALN4mn4drPyf7dJvele+6OWGr6Hll8AuLzCSCLQ
BJEQeOpKBye7ySgIcwBN65uL3Xcrj2LO3Lrc4Bh+QswZHm2K6C+3pHr/v50DQWSu
xd9pW5qlUWoLliz1gK8NOcxRT3/9rS+Ic870geTX0Zu+/72rLhZ+ruedrW1BjBT7
N1a7X826RTBHKbU0ZkYsb29Dej8Qx0QA0Xwk/rhCgIMOVnws4bLR7RXLUgJi+XI4
UVTEJj4VojqUP1GpyLdLT6buTvnVD9bMM/56k79CMXRaAY0XrPV/aC3nr/H/Eya6
e8Z9IKF3NkeMTLnkUtKxLOEkGYvODYbTtJUH39mMNGnpmsuWbR9vbBWTGoy8VpE3
VPFm46watq1FLlPQeFaMht6MgqgZwePBTrZ6ANisMtxcmUfN9Kn29o/PRcSQr5id
R+YPZa7R0CtvuVkKE6anCL+dPIHFM3tH4r4hmtEngdtKdl7XXfK5vem8M/MTwLC8
LZ3uL+SXEPkv2ak4Zoeuro2A7b+BmWC4sf+vGCxKIakuKWI/OFmqR5D4auEaLM79
ZRn8+XO5SjXwGwtId4YzEd+RIfsS2NOL2i8f6/0Fs+pyA9zRDMIg+IcribbSYem3
J4xaH0ktfZHuXtIrc61fB6D6mjgTd6LXDmWz9DZsj3XD4SSiqTDBlLpJwda9xd9W
xMh+x/NPvIBKUEJBgpA2elWf6r+WqceYE8Oq7DxCtB0+KnQ21A1suniML7eYDvax
5K7EmH/wJ1TZ/nZnZIKi6x1iLC3KHtI4IlX0WhVAygjCik6g6G+Cw8zGFRSBdfxA
HOn8meOEDVzyhOk8zSkx+Ipil00vlgKxQt3lBQmnSZmL+x+9nF9wg0+lA5cOx8dV
7YB/hBeSMOR+PPMlRurNvnCQmWv2sB2bXMV9mhmFmRqZgs2mzXzYVDLl/1DOJnKw
4duE6CDE33L2hrMY4LS4Ps+SHxHQhyhOQQUF1KwZiVNAHdjSck25m1BdUx10Kuak
+808y1KUYEiNIh77GrYZiH6URdaBljGRbGfPO+hPdEjs+c81mwBZ7RqNXCX23eZM
JJ8PX/I42qcrHotFTlsDTnaomqwBKq0lMONGQYeEInBA9XelkXFqwhgobNufd61e
/b/xqGdTOLgy/CqbrGKuHEHWTUaOjCPiAGBNqzYBgw08WeQJyDZ2ilYBfnorN/rG
QEASb7RbcebAk1+moPvuUfVIxgLSTbKIBJRtUnsc5xFKjpDz49PLSYzCe93VoXN8
sdgUOjPDkSYyyZEOCc/juk5IMyCx4D5IREfE38uk0+Mm2cz/wkIPN5qcts3FMpWg
pUrxipqJngE5ElAB9k6S7yGVWTBY17NlhbZ0zS3qU+5SkJlSqalFnx6zvqX3cThk
6jg1vTyFwHxF3bKf8yeqFs7lgJ/EHOPUq716flj0fMEBR5yWq/vY7aVxDBQMa1d+
4TZrYjNWjJJgs22o8eW6CfPZ3keTxLl9i5D3FcLkqvbct0tLssKrja0cRQqmFa7B
hrgjS+rf2pj7gQkbkEFZa5GYt9pUJ3H467zH3d5Ran78QrHH3KXrHBZs46QnvZhY
88ltQBfb1apa+D3FiAYJt98m3OJUZG25Cleu2uSNGCUIEn3k5PVY5di6bx4OEiZZ
9eCY/UinobRaa6Lkh9n5yxdVm4TD+Ng8QVBkvyGFqZn3RuqjDn3fS3MgnTEu7FnN
iacEybmFBn48sDXePVHQJHDFvyzpRCKXCD/0DkdkObZg043llTjKMKVBajwxw1Ja
eiRK3wn5NAymBeWZQf199HyHVx0SYsy57IUgIRe/qrAlJzGZuDJujzIAb8DcmI2g
r9oq2Iu0VM30en2ttvkxvcosndYsuet/DGvFiGnX5GKnLT2yR07TRxQcw30Whd2i
fe8otdQYP14j+zq7chWdR1taA8uFkZh1oWSeAXiYFZBXEqPYKcudTLDsbMRESzxL
FK8hewq4r1db+aW6R+Sh7JMpOGBu2qd4MY8A/kN8poTgqpg+bVBBBdRUx974XeVW
s6Ax2KUhBTMkklR4bUL4NmVb5sv8gCuC8/X3cCElaMJNJeFcY4gl580qcxLtbDTp
srRrZWv2T96y05N+Ms9nx7Op3d3FUUSKpUuWXz+ks9sa66D15tKRr9fEnFwdurN2
ddcHvY6In19iYooRsLW/LNZzyMcjiSCzLbda2zBI4UEDQlPVTQAemotLcakGzDZk
uzeIy4BKKJKqSVpiRYm6p8Cs/7AuQKxxmhefXhOD7yf3HzoicDogIFLHeCc1iPQ7
LAXLNXbeo7COUPszGR6z+avuABZy1QhyWSF0i76TaU5UHdwsMEh8Us10nZGWa11g
kEE3JrgDGiXz8g7jTsuGY7mLWkFdg1KKI40w/sV36BNrPCrBH4YkEEO6LFk+/YDR
Hw7rRvUpe4lwAli6rAUhcP1T6hobLNFnbI99wmTBGHtVQ3E/X5wfgMRhX6BXv8ya
Q0nRlH5IpXrl5ZjyKGCSk94Msf4stKvxjLc/gH5DltwCoCTNTtdfGgSoTYyeqpC3
fKxKiTVUAibh1hk2Li7shg1pcF/FS7Q2msK44jg9cMF+F4kHDgyjwpXKpghaYgvb
0sniq2/rE/jAIuNZj2X6C70XZdk4QFv8cenKItU8aXg8TahKe2IsC681ZmJmiUz2
L7Bzt5A23FKdKVC/ZZc9MYgEEEH/HN0wZ6PTMemghhQFRNH679EghrOKqBwcoW15
WE80FD566/3+O/SFlire8lXFCcNQwnw7IHJRYLmHwbZr+bwr5Wo7LW7Umyq2eeYE
u5V1ujftsWpFc5zPEDq65t8jTplC4OK2CuhUt8a0dQRJFUQxQNU6b/pwuAF0s7Ze
26kKkPY12hiOYIHEy0Ti4tHLH+SfwS7zKyASvhF5WHYUxrjycCRcUuCUX9M95OCh
YqvGJNfaQU088i6RkNosO8gkMi06CoQhI1Pd7B/7xDbcdqXmnOXFGziF3bCniExO
bg5Mf/RVp6TeYu6J55UHKh9TK9Ag1NPa7O7zfZAWt3tWkDT20WBtMRMdv2qY4ROL
uKQ8Kiqb8Ap1be1xN7C6wOrKeyuaDnmwygHw4XqDfSmpaLMnylsacnfYAYxo4nrj
jzxpz5fATL7gH7F+iEeSZO7G2lzcaE28S9EIqUleoUaRqHCJKAMjbIZ0OLdx6O6Q
Ejjy+B/lAzNutP7XoI71i4TepA4mE3LyWLCPE6rXMJKz/dUd81c8X/XjEKX3Lgn1
9ootFianVMJXH/irwkAJxGMxIBzmU2Zq9aYVTjdGstMqYw9xaNO2PDX/qjqcPHse
OFiUo2vxKPjWoVDz08TAn3kKksxSx5hbcoRjS32qJQhWC/4xotekF1e6ORgipSLk
7qbC7X7o86b3K6Zi+B994f9Y2VfdMlYGv79L7R48bCJLvFG9jepQvxdTDJsF0cJz
TujzOMF7DdCIJ/EO2u39YYl0ZAxevITI9ah9Txx9oO6Tnlipt0trsiUUAcagWkeR
Dq1GVjQWugX3Nwivw6nR61p63LXT+WalUlfX6bR7nF/MYcHn3OO4vGaFcCDhKiTd
1tp/dFKiO06L13BW9nRgpz4N8y0tfCqDzbUlmHa3vZX6SaMpaTXlCdbE+V3h+mpa
kjP+DPfLDIih6MGpSRecAcgNGAE/jZ4f92r7NR/21+uofcrkFuF6a6sdTMPwIaXD
msNtvwyG5udAJOcx8Kipp3ZTRUxyGJa8r5tdtvvogWm41IDckRijVEmc45vqNo50
0eQxAzXeJxytbUkTRPE76WKxkEuPd0KhrNzFOztBgZ2y56ITmlZ0b74OPkXbtRxz
Skj0Szi39vycNJTLhIM+MtGl6V/XK1564pXEkzAhA5aFxL12sna7T5nEiZPgNSCv
UjmvtRaCvScQ+EcBVoaoYnoiHMrUgR/FynO2nMeg4RUoF2lrF3eEGVUp2zMITvfE
uBC4G2QSJxKh5z7pmZ3A3ml2t6TrbvVmvh4l1jL4HuMDHzRdx/YS3V2HH100pnMr
x4AT8BG7g5Wr1R0kg2wigDCxw8vhKfbcYgz67sVaasFBLnBSPcVoIoyoBssvI2/Y
8+SmcIYhHT9551dxE8Gw8g4fm/hEJpFcGvy0N7ad/D3qw6Rr3WjbQixfVCZ1Jac+
Sb/OqRxEh1PaxYl4CTKV+1CaPRFFTsfC8XLsLsfhM8AmhrIr3npyEK31AERSWsWu
x/Vi5udCIAP8dwRVHOUA1tzq3CUdacKqL7SWbn9al+aoNX30BnndExEAEJBczopZ
uCW81AmaG5semZcIDe+oe8fHI+2k8PevwQd0N45o8tP/Gb1NVeOaiuXQxv8Z8gmo
ZSSV3dtZVSseUXHCpRfjZ2xhV8j8FqBFDwOnG+sRsox5csDz6KNCA30iT9Yj9Kg/
4vny+I2leuosk6pDnv2teXFgq6sSb8id7hHnYbbVA8I4/gWvQ9lDDX7A1bhv998u
o46zUzyMV0zRa/Y72ML9JT0J5cE4jXNCzE6y0ioQYV9u3myaEy6eWORuccuE7iD+
gURnxzsnTt8+Spn3VNBQqJYOctkwg2BHYJvOQTlaz/Tb3VAuJDQOejRnLrozv/S1
0InXMWvn/6Xe40PFT8dH5UcZyQcMGTDm35SZBHnbx2e7nWmGUEOsk7HDJew87ZkL
MydgFcQoLB94m9mJiZF88mkrxMM/FZeehgmeBa+rPcNRYQ/PAC1pWRamRzk21/ci
IL9aYpRM5IJF0OBJVhBdX55EW4vDf0j0RcLtiMBsIgF97msw9xWhkjBxPLYJF8VA
oNrF5/lDSaIBn/KL3QIN41i9UzdgrQRs4nRNql9HgTKVlB76409SQ+9/+49cP4JH
OP9QZqvdVhFTyhKg1VRiSq+zkgvg4nmrvk44vkNrQeuTsUbkKjGvQDMnabASji0X
AcH0mCqxX71Sxuu9bGxbNuhoZMlrZvbGnI/D2vmrI7wJDc43hIoW8MKakWwQhRM3
hfavsH3vQ9y2nomb6Li29GZycl3CMPr/QZia7twhzI9RVoHoh6Uiem58vjBv/rY5
Ay4S5IW4V4mvjfJoLIDcFESGYPtQ3ZhG86YjEEXRYBbKSwxc+tZj+pYyc1yakIp9
qB+lhraa+1+2OP8EpXVNIJIJljZ8t+SsM5ff8fn7I4y50G3KhMtplBXZqfs2uW33
5RbVUVDkO3ObY8yu1HuOzYXES8i7wLxefaEXeKSUi7Ad0FdQlnZ69YWMmhYfhapp
Oqa2eP6SI7rz+602dHVnyCUeFMGXFlN/5yOVGs4OFZLqDQGwfsKBK452vvcEhy1p
Dz1XRjqnr30tIecob3W3i/z714Vg33YfmZtfEb279SSxkUDpvEkek29NVifnNwiO
sVvOBVJxnBkAzGV5e6AyRelJkITKWQ4SIuEah6TS9ujU9uMTBNy3rH9EkkHRfU+o
fO7uDjmZrAUumi1G0XOWpHwsHOzWJN8YzGNSO9rrclDT0W2fmcrHFcHkZdCathGk
cn3z8LEL5QNim9mvT3WWpRVyZTk9zkZbGtoQaES3oFSJD77RZne9c4+1CBOhzuM1
4N/5ho/Ir10u7wVtbrvUgh1MD/U+6de5GXB+N5CqX8DqWrzMwzypSAoEUInOsyon
urqZBGBoFEMgyt5j1mdYrE//gg/xZ7jB9FmZhrKxAro339aImyYO25eoN3ob5Jwv
p9m3kGPjHEytZWoV5r8sKh3KbNYhlKohb1DEK2kHTXJSuUS1+sbSHMEcIOAW4g7Y
3i89lzVV6xvZRc7TvSsOsl9zGcnUFlBKc9zyYzS31XMeMzN3mzdZ59Z7/ZIBumSa
NwoljM9Syckz9/8rTiEVwGZZa7+0be9PdhRuB/eNPJOtSCCk12rvbBtPPcCTr6xK
kW04ma0zmMaMPPdaRrmwKstNoBeqHmxscECYWZu9nMM/jQcu+tbg9LcRyR+6JAOX
UKjGcE1cusB4DlMOjZWRKFdiDXsunUb2Zm7hHQcDXfs7ZlAqJUuAlhaGSLkpH/P2
6k7X4pqDZwaIrxumY+9QQwRIGMmRK29SBVqOaICU7EcNpOmxcmczEkSa87ssbS1E
TtjHCPLtymmKsfoegtty/4yx5xq1Q7ndm172B3+x1aWgYtiYyN4k3vHQApS1OJNp
GtULPv4F/fVW2rrRctt9uznNeIGP/hvTC5Ochfus9+boklJNRSHbh67iPPb4opu1
AT7vxSswJmxwekYelQqN6dkOepKyOdUzzUyKAXh8Bh8O2YwBxamoeQd50I0z38Oz
Gd5ENzl0N3aIzJCZsxyEn6l0w2SvxrTxbQ5NsIYxBleremeFFWiMP4qSMq4IJwAB
7yn/qSCxU+MWDgm2R7F1NH/qyuNXjG1CtnJpTltZx6ZY9OWPko+k+MnJLhKv2ufI
a5q0IWuxs/4lef8mE1CP10T2BdKsuAwdjgBDKeO6jB0+ATgJPRb8gq1YoBYjc8/H
3Sp+fHzohxJv2rlA48Dk/eeF5cwmfQYQ7TMIC/zZViePEV6mqeniJC+f8At7stVY
EA48h7CKi9I8ebGKobJUhYYVi/xBNj47HSvEZPsnzPSTtHXIaOEuU8HXBlKDXc7T
E7sSRl2TVveODyXNRD8n5Qg53O7pwno+FiMyaW4qVTGY/W8wUEqZlfTqVOFRkq+x
LhsqKY+Sd0HhTQyW8RVXFiZEsbPRLIjUAU7oNC+xhWx+H3WOST2xv9OgrR4okvtT
9BhLMpWrpuBQ/wtj4P+4Os88nRoLXRXtQey0zB9qni0OgBYfD81JSKeE7OFCxT6O
HtMnmb7rrvi3YXO6BlGxSCq4RsXPHfv7+AMiR54roqJXyexifbZ3RVDWi0YEb06E
FxYoYqmX3PR3v4dBMNPTqjk8Ey7QxIIsCji14ZJImQts2pFGHCspbzXhFeTpzYLb
8CzaEGmxMfTG8MDnof1Jf+cmO7FP3RNt1Wz0p+W3WEXLF38eN8VV0sw/TwW/3bXX
Ln2keH04qLEgRIGwQm7e3U4XgJ4iNbYnuwnG6b3xj/X2l+Hte54OBmgdZZIVqXfa
O3pEQIh25tGont1zPncCf2EsPcVNQ2xNGsYGYpOh5TGAJkJ0f4E/6t2X5nvnH5qB
WEbstK7kmUKmT7qIZNLdKBvF5PIUpWPQB0WBhGDGU7w/Vx3wzTeb9Wd7YraBIGFT
cbyUeHmn5IkiHFplgm5VPbPPmAf8ajUvJVUljXeUcY9cN4M3c9O6NRy2zEDhJe1e
QEHBTkeHTwqerQXo8RPtpOcAVDesIQDLglssmAY7n43pkPHcVa9iTE7iEIxbWPj3
P9VSduQNUqcOxqkEwImTeOHjkXl+Qo5FN0nMAA3haEpn5RhBg0t73IWqa4bSvCPX
2IoBUSVFb/1Snr6+8boz3xxnFNAnj/3qtYh+FZrDtqsoBhnhvncUN7zq8QCiVK5y
JOHIR63HOv0i2CrNaQMGkatJGIrZDJ/qU+7u8TmzYA01AMBPn6fLVjH6NiHDSFFb
9eC/KreqHijUpshJPiQX0RbJHO5RMR8oDE+dJ7KlrT+nrVsSSIjxs8Q7WS9BcpZx
zLcuYAUkEo6+YZNrnQC7P8bX3jz10GvRyw20ciXFjmDGatKxY1HppHhAr29R13Fa
PBEAmfwrEMuKHcJh81d6oR0VvsMNUG3/X/KURVQOujqEyEgGzQiXa7laS4aI274f
oI1fF95iEQFAmZ1Alh4rCMb9T8OF2IJ9AVBU6W++iLt0NBTCAcXWeuebyXn2XT0U
Ewk1yMo0oJlaHRn+Bku0F92/WyyUuSztk2dtteR42cfzQOthfzAxDz849F4qsA0O
/VRcFYSSqG91sXJVE1StrF9IECDKDYHrXx0QE3QKn7yEfV2ml+eImMz6wDvPUrBs
D+zqNjxeWs5mVtfhhZ/KSMJpSilB/ed9CMgvPwo3//Km2DSfZRxZ3NCXiiFwmN48
3OL0g7O+IT87aVms6jYPQ7SQIVgVEY3++RbA0CAFwnJF+C7TfSjow5r8Xn5cVBRW
Xjxnmunmvr4k+2KXKxbrPI64nO07blSfRO3FDQi0aqHwnGsAv8r1bpl/nChtCXyI
ZagXAcnI5oC5/gnkSRf4f0kdu30mKTwJeCpLAcPNZ2a0fzJ3P+FTpTE3/yJJIbTL
f5Emrv4UaZG+K4WzkAypq3aVrItl2HZrVVFPoWohFB2C49D7G883OjWeFDO4Z40R
gOOrAo/B2HSmzAo+C9F1+sgzEzXNUsDYA/VTip9L3jdP3zKp3b7r7WSiMuXt6ces
k0CUjONd8e5h/NloNdxhrw==
`pragma protect end_protected
