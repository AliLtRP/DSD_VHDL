// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
U1XmZwjuv1SUjNFY7b0RY63aBhNL/lyrPBEVzqvnodf9lTgOWmlQnc40NiH+zaId6g05uKltwmFX
KtYRHZeOD2JzhvzdJRYzib77CzFn3bSU/7zWOm3kAdnlpUrG3I5Do1lTCsSOeoOrm1jEWoYe9FP9
+7oE+uodi36z+JjCUnoq8Feh/kWBFKdvC8OjFXDlOvkOBF57UbDqNQlRoWoqyr++aBPrNmJ4isoQ
QneeHfK1g6VFh5XpDCcM2zHvz4FrAh5nhC8Jpt7b6BfLJVAzo03YBuuxjRLsoklu3buzND6WNHpF
jaodqILpWpPgoHjb+JR2+zVkTIZW/Gwuy78TVQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
+eDyOGM6z1cWgOJ1OXkqnWTf5cza8Ax4Tdu6BmS4YlNRx64fwAqxszb6XRzO3mqY5p8kjhZMzTaB
JiFVmyknJLH6XT42LK/SYiYIrbJKeNw9hCUH9NpYbNjews2qdGIRk2zGelMogy83CEOvS6+IefiK
LLfkhfO2baHgXi9Lcx5cOamxXdUUkXL3VK8lYWvlL4mP5vV5iLgTAY77WfwFEIqw0FXiGZsFneAl
gDtPlDdf4+dRIYUpkWFc43Slrr3VRq/rifC1sUk3076h2QOEeETqYTQQYHk5diiYVQ49EHZ4jgNC
sTZjTfZOCPS3oWqWyVu/AANv7jv8B6XjM7nMl33QB21dc1frMMI2TpQOlpCVT2FMpuvhCFPBIZCZ
nJ5Gi3bRUVlgB7EYwi3XpHWFJWU/g0BoAMXSOnj6tFKT0Fxpp8pTUKTyW8GsMAnaKuJEkLGBObuR
DUbkF5RqAJtqyK8oqmCjbyie8ORXhTPHmeksllgFmLo2YJWGvA7+XscVyt3EeeqF7Z5gSGuz2x4q
gFGl+gSPGFhbu6gz9TZ/zoILBNa2RMmA8yc5YPYb6T2EgsLRNItmSBgeuba66wyzTANTkvAqc6ti
wKCl3MBZj5f7WyeXSmQj2YMAVHrEpqA6YjvKQu6zHyOstjKGbOj9XC5I4P64ti0C5ABm8XtQZjOT
asCxK4tzk8vYyQHwW/m9SwTKVgOTnWw6B4uJkfPwk6XEbV+jWgz9Bu/nVCY9hs32O5uAddatknHE
ZY7/P5q1fFfq200ykRbSXUdvnGfiKRgQ7QzG9VjR0JEwkZgqnWBAgpn0/PNWYHxec6VBjqDQkY0s
Eghu54OqpDvvVGGLQgKCvJsrUO6e3S70yuEtiz5XviwXz6OHI+1gNsZ6JnSJmMDks/73m6fILKWa
XtuIv92rrridZWSS9oCuu5/mzH6UBIGau1QR1caTpjTFJRfMI/6iPyCfB/Xk8CLukbkmW6lzvaey
8nQwNfRJ0ZZNdJbKvXa26GypT8eT0tzgbUbjDP79H6YzWJmcZWdWedXhjwvb9/vq1r0rsGiWMYZT
0Q8s/9fguI0s36MOjxchIbf2+P/LP54vRQe7nUhx6BJ7lGa7hxW6X+UQ4kEroTujej6Fvu0E1LvZ
npLGZxSLzQYL/8o3wID8n9c3Q33jYcDxztF9mWVeUq855yCDdQ+H095VwwOPS3CiwESl3O2Bo8u8
fa9F6AqqR5Q+yMUa1+mlpC513bH8Qef74vH35IzB1W0PttXK5QK/4PooLoC7lhaMgKF7Z6BFRore
/6aWNEJPgzm6ZdhViUPITa1VJrnEsRFP+JGXqOKgroxlNFNAzd/Kpbc1VMnTTmme6rVlNzyo1Wbs
fkEG9vxd0x3zXEVwIrIYlNzIk2YpVz7x9HXWfC8OzkOCXkhmv1uHAuVc5OiKJ/hqdJg/3nTZV+bV
/rkbo8B9wZ73t0c+zXMC3fQlIjNTsNaRu6TYPQWrsemW5QQRBkkFDne8UB8WeSiOe3QtFeEznAYn
YfGy6L6yeqsNq10Mp0AfzwCDpMDAQK5iXN4rMGYttIWctYulJ0ZPu3NilT70QBfXOsXL/7nHdBWV
fpenXazNhkqotd/rG/B5S0zvXPw/8UqjvMdn+Su1t5+QzCPiBLILrTrJTkwXwZEFcOQyxyfmXi00
/MAWVjKQ57uBGFLBNW5pw7kQjj4SR2/eoIZUUjxUlu9gUf/UpEY6jWbYsdID+ZZPhx0WchyJdS1v
uAphH6iGHUQheU4+fXKR6upNUUiPgo/cTtWL+3eMZtk2PdF+UGDviSgq3h3CXFW64lt6s4KYtyf2
eUVnBWY5KiGBJAnUPhY32iipIQ0EuSegAUkibcff1lT/l4LW+PN0Xm1BoGjFVMo7hEuMiqd4AzZH
r9bqNfX4zaTIpiOjMyzd5jFvWDSmQB2y7F4zaZq1mUUvhAlxoJ3iQZNZQly8fU0OamZT0k8VYJxB
3G77N3L+xFfzjfwxQ6VJ5txcOSnkvUFWfBRnOlEo7VvYIkx6IbQv9mRxo6TXGBwUZDIU+/LN2fMF
8sW95IoaHDmR6qOBvWARtv0eJViPAeFTl/oMK9vA9j0O+hGnRbwa5BAh8MWOIcIc4GSsYd5NqBN5
AB5clXVaa/pQqTFwq4iMkHGIQkBLHHb/JlXgRhi8k/N9l7vMuo0NLblFd8SqxiidfAsu09RoVo4Z
1UfjBzmwniKzDj72c9+PE9C3zzg3gfiLvpi2shqsU2EP3P7R/q5PgE6Z/U5nwy0P8EHZJFeSM1sH
X+tutMpwXjFh1IWoRuv6V9/31UDV5lhV0JCC7W+TX20JlNWQMsm0qd7eaGlqWfuMpk6T9MIHTGte
qCAmRBv1vLLcbdUfCqlL+Yl3oYgwRef8JfPRuqHNNdezIonEqv9x6i/75inbBytLkpe5xClWeJ+G
shiA0a2Kbp9ZfPQebrO9vcAs64ycB6Vhutal6vH2CQuf8PcRsck6w7YgLGs4IDG7Qy4/w6WNUN1P
7tUq/KVER5XCsqR/Y9wqgI2NYdnjGZEVRcGFdbIrhOmsAGdaAlRM6TXhlG0mt3Mt3a7QOhS8QqAO
xHW/bDoQuXTJKtUTTxhrvuFBB6nBKPn+rCKaDFscIV1jmlKy8I2BYEfLQhXL/X42g1egyjTSYizm
7Ax/6iuftl4YnsaabAXzwQhaJ84PDx8JuWpNujz5FwGoTnT1tgB41S4av/NhPdKs4CnPyuquvexR
hMXfC365+6r7s1oAW2zg1w+dSlG15CCVatMImNZzeS5WgJRFvRw3HR5xYJdqNHx1tt9ssk8eNafE
VOro2Yn6kM++qA+WmDysb9g168THl4TkqqvRCSHyxXhgGVs2bB02jSNInTevaNCIZqdtnk46/egT
eDcDi/49MhVpRc4kfRROSzrdylRNSI/EZ4Qi1Basr0IuCrPWlTDniiBZungsE/esiFU+nGaEcuqT
uNZZivyQWKBtdD5eGi8Imu5NxUtu6RTt2/S/32DtSta4Gzo5Qs6Eje0cobk/Qvby5DvRAUl7azP2
6ttTQft+rWjFwrD8M4UIJNZSsmDGpUIcBuhJa4NonuKw50HNvdpmvnPWix17YvjSe9+C7nyzD9Az
pslll1nOHkjrD+6pBzGHocK+yCB2lQmeOc8fUZlPsoxq4HJ6Q8Sh7BovRhFR11zflxGzzXSN8NzT
hPF2FivvDjc2zKHIUpme9bCzco63nL1ao+QTvedBrtp53BqcT9rfLiruUwQvX8EWLQ0xDlkBmPrb
15CjX07p6RtaJdo2quji4AABPUtqQ8Q5uxwvha6h4fRrQ4f6b85oRkOZtNj7AsTHFZ6oUZ5/iGpy
51fPKCzMIaz0FYLZugG7jhWktJHZHA4klD1Wuozifhes1Sqag+x4I5IDG9VsjD+Ny+nGzZdsreBM
4nhql2t0UycJcGz6Besom8hnSdbsdB5dkV5zIiW8R+AVoDkFfhAGGj/xMILrvnS5p2TqCARAPwtA
5paQIFl4L1d1bplN4sexOSrBPK0ctGn4hNlAvb6gnwjsNH43T8HMOYSDBzji6QKQgMFW1lJtKMuq
RUev9KWHr8ZI3Ck1BiK58hk0lrf5+3w6ZBFYIKVUe5RviJBPmfEI/tRty83K8sA+GNMulDMRqd8m
Jd1ycUUD2GWtCdVHb0k+ewKnAifySRhSaQFcxl/krBAcANHj2/Ty9mI3rCEAStx6aiW++aOzg65s
jqHzwSftBTWADMB1Oj/WAz8Q9TlqwIY8D5NEbs9/p3tE5jdQTbd3nnB6abSb7GN9vNXJu7Vou43Q
4X3GIY10mcKbDkJ5vESIgFMGyEMchYRripDpotrrjunimJc6X/hRsnOryi8EXFBDdGSHx3Aft50v
rxQ9NkgPTWCJtbr4VV+GUPdFc2k9pYYwgjyWxj0y9wIutdHyOaXOo4jTGiKcMoMp9bZ0FUPGeQ4u
XD6X1Ekyn9bLYr0USlhx37tCuNF0VZ7bHnjlIGBF3eB8legYyYKWJX9nF5HhWDr8twp36r1ciN+V
In7s4WBiHp9AdYAcxxA84RY9TXiwV2IMgMONP5eqWyp0LwZvbXTjuqpkry3IO5PnQH2A6Kw0JVu8
24L5IC4qsEhpz4bL0v0h9+S3TXBos1ZV9v1DzWLrQLvqQzKZfRp3AcbfMCytloFk4HDcnpLj3LQH
KaW1wWmtzSeIpBk+PafyLEibeOK9eAbhlIiCHaYVHzCj39HtRPz/UhFMUPsRJzLNsD6pt4VTWwqX
pXQsC2Q4efkBHosrpCuXb84BOFhyEiSjg+irdlM4pAEfEVVJOk/ylhDDyuBd8itC0/D/0Y299uvU
XoLxoVdev44lwu74W9nJQukBDSWN23I9B4WzjXOmUmP+SK313wuRsYJaoVEXdyp/4cCM4UCWdCoA
RQO8NJEO2CVJ5sNk0PqJFhdIW9crGLSCN7zGoIRzPHmVgd08H79LyHAgo2jhn33mNvtiKGl9NgTd
SQsJBXJYdrsQH0Kdv9SgiIuZ7hBfMoP2eXVI6qemRBSffN1e5UPqSUpL50EAcBvVOpu3V1nuEWe1
51GR4rNV3tZI4pgZMD0YgtXz1VfCbAt5NXdL+N80sPqWi3h2BQYu+vjrgXUYFRMGGhKdcT34wayH
rv8V3AfhmlfoWRbePBHpDPgXR8X+I7BExLnuWG6Q4x+MfKEDJ/rA8T2vrOYYcowGz9NB+mvlhu2A
NX7r3TEe7I8tCfgooMKCsD1zjYL9YRoz7jdHFYmf0XWWJPoP3hLVfNYArEASoYk7D8VTRafksQwt
Pe0SeICwkCQgp4+wySW4bVuqiuCcp38/Wi0qpU5nk81eun5jMVrfdLuAn4nRmErPeMJ4XN3/oVTx
uBVmwvEDPb+CbhMyFLueaNXS+YQp0YOQeNWUbAEAtVy9hS6KjFgdciixakLHlDrY6au0LPMiGgWX
itaxYz9ERrJlqFddDBLT9JckTbLTNbrqv/34dYnj5EMzB/Uf7cRWCFTOscbiZ67sG2pZY05ES/D6
/3KqPlfyuoDeuiwnubV2K6jDaSSfkSKDXIljorbp9ctcqsOm2aDwUGSpDtUj9cKCEwXquNu78y0o
/+rTxGgS6VT2WQDAKHOJ+63b3zLTYdjJGUhcpytTO1R695I/ZZPYtxoZyhHQC2M5DNfpX9RMv6Hj
qiHG+xPJX6OrdGuHi1GMTMlzMkHegDwbTElUZOjczi6Fqp0F1rPtLDAd9NGfP7sE32mo0mPINN3k
IJQHmOMYR5YHwPWOGJ9wBHwpgeKHHSSyv9wCGnTt8clax9+DEXrdv//P5Dm5tT+zooqC1WrdBo0F
7xl6OBMl28WT4ateq9IT9BQnNYQviNVnwXrHtMoes0B8aIUtQDdgWCbHMBlCdXT5/FXhgYAM/1qF
TLbjKx8mkK/Uogy/WU9SLoNIibpZdj9FPb1lfEfpHbr/Zh9UgRH/JaK3ia6sVpG7busK9mOBwaJW
UpGlNAVekJ+gbdnnQx1MIo8Zfqa6lJ4O4BmoMb7lS3BQGi+NjjMnlV26vlGQefuDsaoLZib/BwWX
MjP79tTUF2qTVQMrQTHoCceanSvwDKT0jLQ0iPMm3/Dw9xNTHOQPh6EBTLvBbMslvL2rafS859+u
gqX1Z3ZMd8GE3Hdzgw3LwTZ+/TnFHiQQrNCugm3lg8YYVVM3eVm8KqigKAxfNWOgqEYuYhZD7lhW
FXsahnorX1p0JZGQSeHiVL1VIsX1b++xIhKtHwWY6zUhSIbYYnGnTei2lbYR5/oG0RGAj29WuuUs
gPwjnHq9RKojS7HuzAEqnZrXDZQla1D8+ThOZYBRaEeGX3jOdiZHIANjTSqtxb1+LkizD11cYBI0
C+xH1ye1wbKFLrRleUX6pON2k4wdYsvTxI5wso6Mks95Fono9QfbdoBQrnM7QDGL2eImj/PZsFcx
qFOJCItQEkc9DPIGFRfTvVo6qIZG1T//skhelsq80kRNLzTosXh/s3CLEpjFxUzT29Km72B3P8Hl
shaKSqvZRxgA1KF5hqlJIlRXXgra0uFMtkTHws0E4BOdbcHv//hNp7wD/ywiIWoi2NWf8uF+4i0Q
bId21ZyhgbWwvmRxmjmt8IwFod7mYxrnuqGgDwBw980Vm31wKyKtIvm+8tcAvE41nm3Op5+Av1Pj
DN6tV3k9U3ro+7mqSvXn6ozpbj64X5lnWQ9kaOBAKU6sdiVGr+tKyASAdnde2cZWfqmF3pYz/l3g
Y30xOfsWCH0SRP49ykHIrbeG4fdASbHD/RbyKhsR1XAZhpiWSrGAvsEsr7yhNKfWXoar2traT8Br
O7GMIUm0gvNVBAdQzrgl2RE5PZg6U7B7kwn0JTqEkZlxvGdUjsP4r6+DrfzFMCELLn4doSC5/MvU
TGm6izr3GklHObYSte27/PMs7qkRSD4KsWKHyPFv/duVvGc07/KUirviR63pmgtEiGkVx1DVEIj/
9bINMDaRMfsHJumRf/3+nufKSevIK65lGanRpXyarkFz3CnYVSPqxnDAI7E4egnLWPEOSpCD1oXc
5Q5taGiUy3l4vhqI+LE8qq5Zr+SPpAndVmGtK2bKm3sdU4aKUiF0AttCqh2EZIL9VSN44ssccSa/
c3194TggCfIr3BCeNQI/gJJDNQrXXPndZJnhttKsGRs/++2ezvshD0Fu1d70DWacgF9N8baiywzY
u/j3WI2CkrgenSxFN5rWlqeu753sOgd4R4yJZ+ATrkCSckVSMXw6FE1+PQGTb1vv0J5s3226hiGj
tNFIEXLyxR9B6L2HoqP6S1QGHkkQqD/xgHVGawyoR0vjEz6mCh3Z6EGSr7LaGeAqeb0cZn42NK2J
5WnguD+qvET+/Y+1s2ige0HoUExrBdkEFx7S36fVLG/boRuxOATC2kHBr9SkzC090vdEzZIUA5K6
rSWYQa4LdR/FqAJXPb1AW4YYxekLx46au3sh/gTKnhnvh7SbgQZ8lD/Y0xEbsBYPytvuOGosFi0c
w5Nx1L0iDeYJlaAgtU932EaROT+fEBxssY/hKnXR4W6mAqh/Yg9yu2UBmyCGT+ATr2KcW8dizrKI
y/DsJzCTsSjGoshMA53TurUFsb28BYfnGCgmSPkCrJPHrrhEkPplljXDyvJzZgwdwIFGdEVyWHQX
I1XuDwyfAL1Eo2pH00Uj2e+iMNFdTRVsydPyqCMo3EAOYv6hCY6NNISRdMhwIHjM24NNohb1+E5r
Fs8phKUJtG1oRQkqzuDn+hn77o05GGen01SuzyK94Y1/jSoaCmW9XCzoMfoPQbqtii4Lq+FtT+s2
0uwZEYSQgLFOlhLFi19QpmfCG4tJZaO9qUeZSWdn+Tj3lr9aEEqD3VdPhpjpeSenbwxzCU/RttrI
wllMJAv75LTCw6RbD9gX9xyx/7A/nvUrJLMESdY22WA3Eomj28LnKJGw+mcDf0qLIxwPXeGdmUqj
+RYd2H5dm/0hQAWBjALrpuYHU08e80cacoVOapTeBimt1EbQ54oiEYKBzxLUQ3ilBgbRkk7LEbpg
EAD9YTvFEzOtTrzUvgPp9azp/VV6b4WaMGtJEBlRh3k7gs4RVT7GLuEeH/rbb/g+hEEes3Qwdcjl
eeKrBaeDWoEXfe7Sz5SP4f/2L1dIwGcHB/F5QZyTk4dI0iJBoqy1nTzWh9G4nz8P0TA7Ia0HFY95
EvT5zomLexdWBs4vzqCPYiclxHbJSoMPrdvXKGibfO4Lv6Ub2PYyLpjkjG6w3DpeoHibIMIWM0Ta
ULrtKbAFjh97qEPHHwRgEns5m0B4wbLWUz0r/EcTkkvVd2BauZLfMmuzBzbaR/OtdeMp2ki0OEAQ
f7wOjWcM7OH9rY1MSyg34Rvh/7kPqdCla0vM5b0Y7/P6vB3KCz9m7l/SZdmzP+adYMrTTE0il4TG
ElXhFKt8tHr7qy5cUrgRolSVjPSAJBXsOrbkR3/iZTZcNY5ABFFQkFKTz+mSos1/cYpeZolofZig
eq3bgtCdx7IPHfbt54vseNCh6J6UFBAEvhGEuPwbJCbWVYCfyROrmBxJv9uV3TA6Ur8Bo6BUCyFp
QUJYcghIhMNXgecIMhwlHqfMkVAtC79xg+QUSquraaE6ij5TObEhEfW2D43bQI0/BIfAHH61XdxE
/pFeg+v+ghf0SqldzgPGykckRWxbP5b4AtFXpBNrODow9ND7D4LrIyYPqVz2Pv8fOwW5HQWY4yrG
zPum7vyMrmQ0JnTrE1FfEnhWAsNPYNn39NHfbdvxNIpslqLpW/N9sdc7ZeFvAztUtlossH6KWlZn
PBtmYXiqHiBWQv+L07xA/AGQ+uqDkFw7+FpQXz6W4MwNkru5CNPsifrw3piBy8ys6llFLwq7zPnC
Gxt9mz3abGG5UT7ZHyT4L7ei5S0sYsGVRTc+g6AHBAuggvWZz9SsBxPGKM41NDJa02POnmk/pp5X
w2o96CUNnUws1evV8fMA6W6mR+xPuTMM+IEFuw7FVPw46I/PWvv/F7o9cKJQQjcMVRw+oruSDY9R
TEn+mA6YSQqx7Jfxc8RBiPNs/cexQO1dWS7oFKh9QrMUotTr0V7hBVQV+lbqyZBz7+JoBGXG81vx
YOdCDK6FzuSVfCxymJ8Qx5UMuU9tVs3240RCh8xD1vpvvwiKpfUnFIGP/wAaO7meR20hsjcTHPk+
ibWEbdX+RIdlHN+RGt288AaDvIb4hzPpsCWRxRvJtrRUEYY5Zbzwb2g8VZPbQ+4tiisJJnj0GzQp
ROW8yTOpKQtGIwWy2IWtKbu6j8JUYSDB9WafVAI3k8XBUsLOX94OwS9HprLGo9TzMUrMIboiKR5i
MN0wM6wYPUrpia/eRO7ToydtO2HwjEVbSQbp5qocPJy9QttOI2A60mTEgJJ9xmoyFOcR3/BSoWB/
Ov2uPe+5VvZR+F0fUZh2cDj68qbTIKYkM3uO5212jP+NhYXWR6yV71m9cQ1wRhqICzu9PO2fn0Tp
1PoBbsvSg9Y7/yghRevqrWqRZbmNyZOy9CmCf6AD8elKS4QndetV4GwZRy7zuVzw+xmYLqrGVMh1
h/I89PXa2YofrXsGWfpbrUf6JtDFVyEtrc75EGj08NThEQxInuiDNtibTwLUrReuSSXqYcV5gYWh
4ifOGX5S4stHZNsZOUHb3C9VlFq03Mge+wzqA0V/jcqpwcFPjeNPlW6dm5v8tSvGyryMyLgf6MEc
7pUA8Usmi7uxunfrArXMgl3xkNHVplOs3j45Dus+QeTWEh9IudeOvI46/ndTvIhoW+0nrMB5YhNb
V8n9mVwRx9R3dbngimkQq//GHjLPPCWCLnKqhKubq+uUhHO/zgH+z6q3+qxzwVR7UjnDJB0ub1Fa
Tn/IH4vsmMwIo8YCiBY14lxXVUjLXeCl8+4KMScWZWdCIjRvE5ikkMXw20Ocqoj6eMTgmN8BvZo3
qc+VPpHgoga1hbwjrGomne2GAfZkUMrDly3UIekLv/Vf5z+i+zbf6HPDxH/jpH5jH+xxedIquHZN
B6pfAbpmRltmevVgkDIchhZEZ3JkhKOKwuHqUEaisekJC82ytjhN/iVnh0hpFJ00kn5iqNDaJxYU
zqk/jZEJwPj0Yq0gLhpRN8nAxNsKKhB6SDyBRf3b93gHF0dXTxemEW8K3brXW0F+ZDzWl1Xn7e3N
ZGLIMCCBcNZn9iFVNGaYG+3u95NN+d2ZWD2U0Jxr8vS7nhPT6l99jaLW+hobbTuOLXC0zpol4FKn
jgALWAeptq/UYr6g4BedY3JW1jB1EMNHv0mZf01Do3tW4I9eoII/4LpOsEmomwxRFmNwzUxxWRKr
bZ8XrEL34HEKxyc2bm32rxx9UaH/RniAybETtBGzOdiEJz3+jHT1mhTcqNp9hYsJ6GSs8xpv0iiK
uopKYQ+iJphRZ5rhbmrEaIj2uRnR1SmNCQDdvaQgtopVVJ66UVxVKtN/Mjw0Pdq6JlEqXnlSW80N
SRsJmlBZgknMfUMabyGuPmg/a/k41O9bBf+Tzzmi5DWMNJhaTKQdlf0DSM7z31XeP3S93RC1XOVg
ufTDOi5gYTZcCx7CPsyKMvUVfbqAKjv1DuT9lft+ZXQrSTWxaUN2t6EsYA9txtjq+cbaSr8Hmhgb
sGYk6PMOsazO84eFenOngtr56TZfR7tXsdnobjcEZt96k9HlFCpDui5N73aiXuS9s/GboSA6qmBz
kD1zh/rmbaHKWqPH0C/yKfCAIRTbRLCsbN86OTaDQkBhwdbKQtEbit0a
`pragma protect end_protected
