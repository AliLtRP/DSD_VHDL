// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
b9NedOngg9xBc6T/+DoyabN52bj8gqc3oXaCHyAjclR3szz1zGtSj8X6go/LHVWr8ppWdv2eKQW/
ZIyDr05dArnOxF4G7pKLhb+ZlfunL0m9if3fBX6wP0p3OFyFTC2Wn/+4xDgXMdJCEAN8U5z5BnJt
AfGiQtafDuOeC3hUPTxpjf7zyENGaJYF24AI+Qlv9q1eZdeNNc9UhRoXcbEy7WgnJjbgtXSPwxXh
Ef5wYdKRPfJITACogkZNFArfkxgrDRznHuVo1/s4vAJFhaQtmM/8D5y8DrEktmhgIqQ73Aqix4by
LFR371EZ08pEs4WHJsMiKVW7/d5Op6KCX3VK1w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
7PZRFdiUNFtx0u7K7cmw1Y3MzgifRokQ4/zYeX9bTPp0MjKMyeYo9UPMxeXFJ/tlLX5dqV7ODaIs
sd+HZ4zcmFqG2ErEmvqzspu6yAIw4bfOjnHZf7sUw5LcahSEkYyhUZ2svYNR8n6V+6464D4TSier
mrC+ESpQp1rCSFpeEh1lSKKC445TQE5TWswhP/g7df9e2sur36oecMAa3+6za5uuvA5wikJIp6yM
i84vZtbX+0AETMK7D7IqLSP+i6+mEqZ/h7rmHjBK8TlW1jn2l51KRCPhN3m41rjPlyNBUXvzoKge
sLPCeNSTHAzOL6Wu7tBnRkHeJFALULtcFV0CMFDVt13xBLsunvrJf5T/jXGXDcQ2LsauwCsgE/xO
gP2jygS34j2yzkZ8WtcC/fdzrAPMWDV+b11m1A+DPsUakCsyzl3FXQAlIBx1gavrmQf1E+dHom0w
U928SmounnEIr8oyEiLrSh1xUgNZRRFLLdvybSIBfDco9kPllEIw0+mzxjTYiiLPeUlP/Gl5ylgw
cu/O/X2Txm8uG+LJJ6OivRz6egff/fZEgHezHaMEyfzOddAMzU96wQH/TqOjLOa+uCuIyQ1hBZ/d
7+P9WWiFqtmJlV1PYecVKaTm+wcp/gfZXG/dM3PZBirLCCXqB+JCq7saiDYjJeEB7USiwjgZEn39
N4J7JHKWs/EATcojME49XHDeKBMaDkbqVr00pESnK1pN5+sWMVQENH6KmiJzOIwLsXnb3tIrgj1L
6e/IGNvKQBv2a/l5scR4/mR33JzBTjRX5/UvylVp1x01b9aiLZVXglk7mEp7FlNwzK1CyX/zII+A
b4mJxhCKWr7ABgLtFFvgBeg/1b4LIR4laFq5ZOVE3VBfqTwL1vP3KAD/PaJ8YAd/K8fFAPK21vCG
95sUG9Iqo1O9yEi5KUtObvWOucKPthgvDbyTBspT9HziV8qpQkgujkbr/WozR1OPPOoMVUEbfjRf
co2mLz9CbEW1oM9ut6razI8MzxlZ/EA+xIE0DVIIqhQxX7xFCcQCXNDhHGKUcrPxyuaZpvaSOJU4
Cy0WlGxoj5G13II6n9LOLB7VO0sYs3vr7XIf/MpZZ485ORDj8XxqpUIE0rRwLhy2+hewvUwqFz9F
XeKPJzwCJNyrGcTelLPTwGunc5SecGoX0QYoiu8pEXjzoAkCGPMdArxUvKwtPtCc9prwHQKCqZts
XInzduYr9RUB8w6X8Lo+PVBZA0J9AEI5Z9dE0yTU3G/mkHlSGT1kBRKHxp9ArSF6XjFARd28usuU
IeBsYTG3vG7huHeMCQWEukTuPQdQi5xWheXlucwBBNsl89OkCBbumqk96ED1VqZtjjRxmmyzlFhk
sLDqdjEFN+iYbv95LxlpbWOEsTH7/Of8lVj4ZTHDiMYO8J7fbi5bleHC/jrHQYBqDPfL9fpuZSh/
B5yqVzbnpE7s9TSuqY0e5+d4M3XwhGQFyocImEnnqDIsGvWl9WviJ+Li0cQYhXBjIoQiUbkad/cX
J4i7bAJo0aLzmNU/pxzJrkyGhKf+ThRK7IDldLTGfXueaAnOzkrRXPxYnktzxsDoaprBROlb6Q+Y
2IdNE62OALNTNFJfAJXtkMVkNHEO1hiY+axnvxO5DDQwm+SH0YMtFyiJsye/pHwTS0IXqkvA76yY
U4Fzpa4RSGJuW3QY8Z99C0r6W0oYiXZe2JYBQ9cFGTsrf8E7wZqYjXWl7bAIvzcBxivqlPdmXX8F
22PVv2ga1QYkKwgICfm5ygzrCtVyvW2wA8xPgB0BvRAY/IBpJYCaXsYz0pg3byRjNNypInftESmG
dusOF2Qs0sjinzQySEZZt0Hy/EPm9FfJzPvv3O+1VH6X+8V4GGDAId8ahdeRM0kHZ71z/LTpoBO/
UcThLiu46TctRrUITJmV4ynQy+by0A6tTV7bm2HL4aucm+ud8N3OpJJ7jlbgIRF781DWXq9W2R32
Q7ZV5sGAF0j/qIyUYqBVkMz9rdEIpL48d204xw3DiYQ9xtDIpoPORNHjzv7ryGybtHQNjmFFc36/
34GoLAQLA9EkwkWcu6KSZONmLmuORIOZRxsIQ48Oe+v1AQ+K6GsvS+ZKricfKx1h6HVxotM1qINx
ZgaWfvahWp4jCSZ/L8WtKAOM7pIAldAxu6+V9RavSofshG2ZMknaIvCYSkrofdSA4S3dmEku88Ba
S2/SWwqv3C/Do2xIK7qxGo6hdVavzZZBVwwTmCBzx3iTToW2k+lIsOHj7gK5ettp+fHWPwi79AF7
8CTrUBqfWUAe9B6jgArYHoz1i0h/d86Pf90LxjZCfRTDO0PDT/niJjHcAEbMaTyRH1da3smd06FX
sRPGuT9d/btdEn5wwK+yWTpf7Z9XPLMIA2xsjHnEcBf2LQkRvYfq54EYKqCs/P44i2AaLc5Wvt4s
kCpZlmNAiFV1Ps1GQK4tROziPuynN50fYk2NcUXUpv383usIAzgQuetIQFdRHjdzlGIs2bcD/JN1
yJTPphB2IkiQ8yYomuQTQr88Noq4LnmJmZY29IytoNU3j8StpENH9AlW9EHaQeVHOI9VjC+giv44
g0lq1YARbN02tm573RZfIumDy02C/FMZV6tQf3YMAMDnXdDFypYBH92H6sBIhwDovZdVL64aDsNA
Qe5PRaLOke0OIjcSDufjzmq+pFnFOKpC+LXXK7SJSIHB0QOqju1yGR7kMZoYxc89I8Hs9VAvGsbr
FIWBMFhHLIcXaT8TGjpVo9eeIwEljUNk42DHbBZcvycKdebChxTGgddqoHp3HTnbZ70DITrrD0Dy
W+ouE/G4KAv6F7NeqiEWobpeTiKTGYgp+AAtHc7DsZb6sbrfXvvOYB6t3vdGd+LfKaNQEA9Wc1pF
7F2zdrx3YxPoTVxg/gzzhJ9nquEHl1pLE8yXovSK5Kz+P82EfTNivUQCCzQSQs175XUfklvqsqhQ
KUsh72C6HFqloMPy92Vd7YSQNqwKn9jt68aLULbtCbyYG3BitAnhqrAE+N/8oMyNjf6SPMsOb+8i
aPnIzJq3/ZQzS9bme0AwHkzo1X4OFwoXt+RjLWaLY0EKYq/POVFsmUn/i5UU3jWmSUbEfT0SGcSL
PY1Brn6bam/6zeb6p1oBW7y19DVf5qg3Cpx7n4Xsw+j8kzT9ci6m5Gi4HrUOrdN+Xl+IqC37nI6f
ZTZ4fAE5WivWp8DoxRGANSZdrl4k8AGHismcdQtmbS8EgPE2fNbWI1vn2coOn1mk6cbB9d3vVTms
Z/1arW12NksQVxgmcCjdpblAo1GmFkKTLifBYCI4Cniw49q5fbJMceyn3PfJXAGR1GkhBzrekPzL
Z46sKE6sCjar1YDMD3b6bX3hkL1P7pEmDtm/Ttek78nWEkbQaoWGZOueAMCIovbHjC3sTRdSfIUs
ZG6mH2uMR/WihNCFBtx6mugcgw7ahZkSgUGNhlrZeD0K+hmxCGBMRIgpu2cS9kfkJ2rMk9VnyXXf
sSVTiUYdwwHevcZ/zEtDAPPsJaOA+3dcR6r2SiX2wA1JN0KBNuqOcnPMd8ZIW1Kv5ditzJDl3Ot7
MfK6jwNZSsBKPXJ2g5xNvK/9EjKy8w0q0jD+r2EvQws/GoPBrV8ctyJjkpT0A59SEAikIeZEQu6E
W5yHl+s3X8ea4f4zpqzP7DST4I8Mg5F8/nuDvgyNJuhk7rrrFlIKrLde5J5YZQhuN0nHH11GeIWS
pZ8ljs3gqGfWVPKt7hHtQI/QOnRIDRTg/G5yFqVVcEC0TWb5eIwScgtytW7kfRmUjCtRNaF7ufY2
cvibxTX4ssH9pwXKeds2GZuTpVSLXwzhHhTz3Ogx3VLMm7x+i3ZYfjWfgZWMIMxN4Vp2tPYkbN1q
mHZlY1rw8UXIX9aEQpyk2kb9JBboN8MoWrU6P2T6WXhE3bKkcGz9KyWbN0VywuzZiUBqIKTH3som
YyaHsucMtvnQVuqAg8nhojbio/24/GQsc+Gyh8A8f+z9AYDT7faY9ncY2CGmhFomBN1QHtSQFpIa
75hj+aHThRUqaIK6YZvp3a/37q6dKe2XkyqqHvXIvDFUhZSf1iMdXlSumrq7CRoCQyL7xGgPWord
8JlWULjYCfMsAHUspasJb4X/1hU81jxA1LH3xUoH+/tsfergcHoox7RhEwT0MKUC8nPdQgAzTplE
L9BtfBroQ+mowQy7ECiUSgeFhXUllFrYxkEgODLgO1bg2JOqDnxb6uI9cdvm6u9SZwpK04V6V1Ra
zLmauQ+O02x4qYP/dlxeS5y0HxcSgyI6tZI7ABiQjH8mjqrRFNrah8ay49mLp2UXVDUCb7btD0Ln
xSUPO6OztKdeLfRmtBvF5XHttYnzFSFv8rYazsAW4Q0MdwCjYnML/cKcf0zFiFTVJQLyKXa4QQIa
5/DdEI5YxUd72zBsN90pgCsAr/OXq2TjBYqnXWkPhQRsWPRevoNVZUXyEi9/eHaE0iYI7G6/2i0F
/39M/Pba4z7r2C22oKoZr4f5qHaU+c5Dc3XX/9NrwTSaFbC5X9L47uWunGOT4ak4EnkEPfshYvU/
EjCoRkqoorRyi9cClQUuc+9ae4QjOSnSiJTWGGIOcL8p7aQLFDI0kE3TFjjWd/OmX33elUKRoQ2p
PvXHua55lpgsscWAFLw1tHrKtsM1lE+foDXw3hvsxRDC8H/HPIGcHsaNTxBXE+YHqup3JICFEBMK
W6UmbrmKVv8tHlZWhPG+BKNet3xhI2EP2pdRlcFMr6xKzhOH3XG2MFNMhphpczx8JCv3rbAPX6y0
WebVD6kzYGrz2NFeYV9/2Mvv7O1VhGH/u3fUtDFyDBFLk3PAZHMyMfoMz7KVTO1pyhjRiB4N4UUs
Duan0EuQP8j2C4dtWYZWX69VZy4zzuDO/SvxIwYn6qIsYXr8EMaDhywFx+NWWOlChHaWEmCKcwr8
fsRTwyC+Zb/hmLjfRqdsVskkUBp/y3KlT3sTR8Ad/8XfdGP/jGQ6z7iCdWfsVrmyAtKBao45Q5il
KZL1c3TyuVxlAZuFs6+a9DcT+lcEdU0BtjOQbc/cfSrM7L+CT6FKNpwKXJ0bkbPhGpwD44gs1lx0
LnkqCnpZjVgphvg6g3/ndxiU8XMxUN7Cs21B9ElvjQZGIxYRuDrWbYV9qlhDsQiiSSHXhDXeimgU
pK5MVPmJA9yhfh2FX816cCU2QuZh52o0sKokwIsX8RLbC6/jIanHWeDe+cpxN79FhCmjfTE7xG5F
TpUM5ZZNqI5u2PMCO+BJ0CSiUoM2i8rFEU58HkOmjcXOF7uBx+q9hE05Cb6rsl3dM/KgVmCVQdFL
B7gHNGlTlFczCZyGOLeCmdR3qTV+HXVpjzPdH+2NzNn6XZg5KrybgdsyulBnm/WIDuGohEYOhpBB
P5do5gmTUHUXL4H1+kETXL3n4ryeM+zbKRZ/j5StegUFzVf10AMLQBgGh0MYAugWX1G/T+l1I7WR
AGl7tF9bXsJ3CP+7x+xNEWDy41fHguZdwUYm4OMKsKuvuwFL5Ld2zUnCH4S4MIXuddSL/pbW1ImW
+Y1fom4N2wwTLwlEI2gj+IJB2pB3y7TEJGRyU1RcyHLrFVu2ZkrgqfNDAIy+3I3SVEp6ywky8mkK
Y0/MeAFncm5WBOAslyRyoG+cicF9+FZfRUTV9hx1lfaX3evbosAMUV+a3Dro6lREx8kI+O0TvR3F
/kQSe/3eH0NvA5Ye66RRYi18HWLFwzphdRJUrwuvLAz/hA4ODo3jCqW7hxG9WCafHDs90efbRqkF
bRKm6G2d+hZNvKzrJsYXQXf5JyU8UTGpBJ0IwNoDbT7nEzJnLzFMSSPa27NGc0lp5jQdoKbTnud5
Kri3Rk6GxLCgEZNhumipRhotxeDA3FWbNg7ERX6YWGHvsJY9W/8TQjhYc3pQvZak1ggPID6q2DgS
Xzg5jJ9rVHz7UT0K7eLeKHZWhpAsPgAFmx+hNaorK/ugQS2eCQKr/uais1aOwATqCfseJo30S/aO
f0X/dfeGQPhSsq9yDU4f8eA/1h6xBvJh8geEOXOIL+ULvl88oPoQzEyb/d/YiZ75akAb50QV7e5t
3kPvcE4XMgLwrt/FYnK2iUYXcIQRuR7KG4gef9pUscfxQS9WWFvFPyqBx6ytbx2R2+JHggnsZaXZ
ruKUKWigcTeYYF7jfgaewu3+yfu+253Z/ycYXQVriKFc2fX2T5cXoaAOOlotmNrpSPBO5QL5iYO/
PdlG7mRBkGPfsYsWCVKiJnTjRlLEnhfGX9lMvkFRTfjwrAyBTovY5PMY63E3BB+UG/iYYwhUBXuj
9naUp8JRvoShamq8vobaA0FhjjuKMrEzG/lgq4k8isNnykAAgvUmJM64+A+lGNflofFxJAIfqZzF
FQkUozpxxS6VNZ1nq55xEcp2fC305GwfK/jzm2hAB9ziSUWxqvBit3eGMz+gNWzjYapohcPfMSFe
sBs/kpC38fUyNaNCgD6PKQPA8oooQE+nZX5k9NH10gqIfB7Kttz0YTPIuERSnGzfMAEcTqIynjPH
Wglb3FIqpa2NnjEfDg+l2kMzfALhW8OuteHHnwpAMn+bH3TrPyyQ9gr3FGAerEeIhMaYgJVaGmRM
zX7f2ZR6yuNKLUWHmEEznfm782FCUC9k9bgkrjhLTWJ0h6GiHMOdXMSavlEI7eGYD9VtBJKzsmbJ
zRIQF8eJh5lUNer1StA5yWPwNFRestdzTLDaQXc5kgUBc5h3JOHFoPfGyde1AwCgMOT55Dy1vaQF
/Kbe96eK16bhXDpVmaKPGw17QLqAE+NTKgpDJrUtK/Z3InzBr6kBSuQuAZIupM8UfM/+OQweqjOu
2I2PAJJefBLz5wcvfnlCt7GryB4ivrnwNfMFqaqONQcor38NZeO3y4gnWcgsQaiYcU16DDA/I/5x
8oiabaAC1bSgRIzPm6fw97Xov0u1Kh24Efm2x/DOMoEQwgpBGnxKfthY7fqyD1N24/zNAzbVO3YQ
J/O1xIKqv+AyFywW58CZbLHcx9fd+ytRhING9klA50MQ9kKulaePMY49UunWZzkQ47PdjAPCn05n
cHSH8/3O5D55+SzWCR/oNQ7EDqC8JKSe9Nu8TzIdyt3jT/Ke/SHPUlh+bjd5rFg8Gm9jO2OLWhF0
xucAnM1liZyTaXAgmFs/ZX6akaoMyN50qshjFuMMfrZJtdkmDYvc5mucFBDINYBXwqxwX2vvbJxL
F42mnIfNFnSwz/0+PC+YYkubc7NyukZhMtY71DZ4rFQZqYLlI/1Hm/tUH4PxdPNkNLVbYS3iygEj
SJMMLW0qx/HB7wHCIAfzt4xRxjrRNhyDlwP0WEBA+K+pIIdfRSJrbeoB4ykM9aC7PNXXZoOfs8Nk
HU+lBqef8b8stJ9jTGhejdjDysvJX/OWY35LMAqOrapB0Sxa+DA1vCb+CL1X3mHeNeY9eg3PT8s6
62cQqtSeqWY0a6EdmF0226xPM0oGmovRS25dvZcX2GtymGcO4B41Gk9qnzIml7EnuPNpNPeqp+W4
hgQba2g+/VFxl1JchCuC6dyRshRDqz8zXvTLUsrEhrNo9JqOLrChrs5uwqCKcnhR1/6657mnU8Sf
hax4UWBvsnYU2pauTASWqliUwntPTJgkXPMyvcpQc6pQS7qfnmZrafnHQMckynzxlYZu0G8HyE8q
B79wUhRdZr984rN/wYvSd4HajA==
`pragma protect end_protected
