// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:03 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sqiZ2FKBHsGiT1UCmlOkP5s4+5xn6IH4bD7XA+76j9BUctyDjCO7xP8fSAl1OwiO
m1A/qtukvX/mmZx+/CNFcSo6pzBGALs1Le5VioUWWXLhNnJPNk46r4dM43GbiirD
6ougDf3ppOgWWG1S7qCdccT2hP8C5SfnAh7omQ7OogI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16960)
bSfm6vEehAv0tdk4hUOLTYALwX8DbwGKsTNNMD0B1wsbUEh7XjBWZO2Qe5uWvkp6
6LZtg8+LtYoewfpSGOeb+vdur3TMpA5StPu7aJYQKVmT6xZeAsl67b2u5fdloMjW
5e4NKw/B4kSw25NDOkv18kUsAJN8kwFw/HbBXlUGqDOCE9ZONszIQ9rm79O2alRs
bL6626NhrVKw0+fBcdXra5q839Oozp9zFz5zIFhV+wqiYF9MS0efQBJbuUjUU7oy
SGOHrtC6r4gz/izBDbcI/GaLzIf0DsaLB+x486aN5vJT8dGYsX3hbKZjeQqmNoJ1
QCYLFKndAtMJ6EL+I8qyft6gcrSoMhf+lrSOWYmhEUNXmPaySwJV1Gk0KVHjJas4
r6CarKoaBpOrYOs9Yfm7+fOTWhtTOenibXut0Zd01qI818AbNd+sdNtpbtqjz7ca
UEfTS08dow7GVy31y3Og/mkhbWamKZQ694l/2OHjCm92dG177a9o1358QZpcVU7h
/hfBZKkDlSb3hnGM2WuzGSS7afeTh4A1qxvbZlCVahQ8yLjty83G/d3EGt6w5Cz7
qceYqDbMpQR6jTAeCs+P9UQ2Vp6ugR/NoMQqewHuFKAxDSnFMl3Eo1sUPN1bMeP4
8Y6aQLNzdwwyRfwLXXFVcfClOdkrpCJ/cpILFf3SXuparJE3AGtwepde+pM6vd1m
LPE2P6jniJU/0iKaYEV62dt6mmIzVy9H5d2GJ5gRmd8u0+jmzf0AoR++iwKeAMFd
uCqp8eNKsbVJCHVCJH/zua+smrVTPlZI7I9Frt4xiqohf4BcD/yXr3lOANhC4yry
i4E3XhPDrH5nQBpA3rBA4hTw4oIAqTi8VJFqROloQfVQraUXUCK0jMPdGtCDeBch
8etw3gN7sG5f6ZknbTmm3s/IlBxtb10XSTS47vkWNkn+FKtwIA9ppn8YKOYHjL07
+9tb/H1VWnnbsYcYdkqMQcCMKYARK/AVJKMkqUm32PLpr2gax6naN532y1V/erze
ouxlxiR7cZyCNjSSBU/niV8c6YsyhJuLfUbA9N2e4NPhAggVIc/towK6XYHgImr0
4lzziGpdX4zflfNWAgkm0DYAmSkDflQXP3m24hLevlzT84pKxrekmrjL2xdyzuOi
9X7oZmDcflvMgSSSUGbXA/FlCG0Vx33gVbkAuVaDr89SOdJcfNYJ7/JqdZhfHDHg
IHwt6E4vOq17er2Rb3joPuzagck7Fi3M9YBoI1M4P2UK0vCHHw9S9qiD5kIfx/gh
8XMrAns4mffcggLwDwtkBdd/rd6c6Bv7XoNXzOlc5vyM6v7Buyi+53y73vRDBn4Z
v0/TClUlDQg7gEghvFmo+G7tlCTLFvpprWfkGqHnFi88FgkrkFfRhY0GFXcuKUJQ
CjASr1+GkUCJZ/Ig9zi4Z6lOmtchCbC4f0SOjuA9bJw20ILdpbJByE/hZ7UtqCzI
/wpO9Ky+wSLjCcmuZECtUWxCTw2UvNCS5AFpdwY8fM0TqAjKh88iu8obIbUBVFVz
efXUXiZRgIupZTlled88HxGPTQCQ5oA3E/P9m7zyH6y/aYm7eYOhrEXElTd0OFSL
W1uWTAen6lsK3H2SRzNEfuBHpAvfR7SryPts56/0hXTmqQmRJopMsbcucdt3Meoy
CC4SI9Kj7l4iGL6Pu30zabN3KUESlUyvqXqk3akSX0vFbaK/HOB3SfSuWj3aDgtz
O/1/tI01JmCCyxt0wJWo4XJkP2I7fkR7hgN/SQJnwNP+hxTeusFoWD5TTjvm2JRb
sSATatIijburxrqtnEHlbbWXbZ+HBHpGxq+zaAkLM9138UhLovXkQjIQ2foENKge
re2sHAkQaDcy50tWP/ohPCblyuqgRVzPMAS0WfTjFFh7AEPIUDR7uPO+hcx3gK1+
lwgoH+0HhPuSQx/pbHl+qxbbDaHJyDICriXt6ELLjAJyrpp2eFnEM7a8xwZRsVVq
EOfXZAvoijn3wu/Dth3N8mrtcHNHWvTNeN0GWD2s8Bc7cwqE1oq+5+mXGgcrYr9g
drE6UGKeZgpU5d8i8GcUPmevpq6lkRORzwRoaf8MY0FTnuhR6AE3XnCsd6yWDXwW
O7cTC83EupiMQJbNf7maoEriVmf1dK937wJwwdpNQwgfSTsHqmGYCkMxDRgrXNir
2BmJHHLHZ7UMl6lL+KbRK2nxp78QBs41xKw8SV74mfbpVS3pGuwKXoHMrJHgiuCZ
Nm+3DUKCyV2+U6INzDxn2v0TyZFcxQd0CwF/JdLNVXyhxyYwSkDYL72kZCdrwxPl
JNLBhVe0H74y1WnYx62hRGsmJpWH3DsSELSxXcaCdowWtuTQKlyv/9a27fT1Hf0Y
zEmnww5wCuSN/ITP5VBAAlWEl/MFm4WusIZOWJqmgFlY7JugTMY4ZzB0YxKf93rT
sAd3wRr98n8fxPG6RxvlBmtMTyagyF+UngZ/MZXrIQLa9SOmchACp7d4rAGR0iZh
DUqp1NcSUZnnBSWRnA2ZjbDrrG1vbwbQJqUiVCsPZ5U7wauAeaVnKtZHGBGCE5Ds
sRpd5jTiuc13qD+cv0Blm771ubu8JzX4D1YqaDZNFOgVTvB0/1kjOXKt7z2mIlFy
l236K5Pr9N1dfAWgYFIr2Lt53CqJStITculLcKxvIlYbXd8M4YfhqE8JAoiqoh5I
45hs7Rp7jvSPAdnFX4Hz1GHSfeKFXPAxV3A9cxl3LMOQii6xIVRFvawEVLf8QWJH
8YXrofDyrqOglr4he1YJdA3oGspUnwWcJgXxK7jATVFf/we8HD1pWFRkYM+z8yhX
lsmp2qeAoF7rpYXqLhuPrfCLM3SNVFuFiWK5RCU37mbcYhevrff9CGd/1xSPqSvH
YOvkrB47Kdybu+AFE8m493phjq2tVAOpH/SVwYqBZpcCHZyysQJQdyPpDDU42Z6l
OE05A+0pmHrwnYLsc6KR2D/FaJ5gRYUUdiUh3zIOWmhjZzNt7fJOdlLKsL/EqLhM
2GuM6HeQQcWoUjYEqt3rqcOJPlDkecgIGoiG3QD5Lh0fhoVvH3XSNEcFUz0NpZfV
L2VATFycXzmajyHUafA0o6ZCHF2fa37QR/x6Hy9vT6pc0y+iVzDHuCk4qBkcvYEa
A4PLF1H9gZ4EvrH3yknLqhFd7MxDWGbeJC2y98C2Hk2mqmw+qUFVXrexdcvDpu8i
WqHMId8cV8MJG5d5VjRpSXjdbaqA8vNp5ZM+cw3jYfdb00RKvpN+liF6wzVUCUe9
kjq10+RJew6f5MNFWwgmLgBST68tf2+20QHBe7jdNPcu1DMX3oSor/Wagea0mS1c
XG/I3f+2bui/gSKZWW172oaPlc7U9gSnWHFbHp28lV6VXXnkaiSW6Db/KpbQ8FKC
zo1Zx7WFKdyskclm128CjwkPgzNfyDb0E9Nirc/Rys4upsSZtinFEomAo9Bs4ql8
0uA9Gy5pWuJRlkg7nbUgLGuy5Hh94Jnu24CvGtdIXp7DmEsoEanq93N1YYuh0bUX
jKNk2GaOZtaaXezCLuLMFsPVM/F+9Ac1WUL1wcrhUKM+okJwkbLp/K1T7QFK57zL
FiTiXxiGlTbFtIVr9JpCdvGHnk2dOHgt27r7DVe8yxmkmHY/dKrtc/CukwLa/FOz
g5F9huG+jx3HFfIAc2VbHVrGzOCjyR3dxa4PqlO5E1NhRE38qkQGqS5hs1gHNlPx
ttgN6oxb7UctYMCPsYEbSKKdG8J1eUQb06s9i81QqHncxIK7rj0T5pYnZNzNRuTc
rA4WnAeAb6y8F37WiUID+KDOANe5cjk3REpO3aakOjp5ToersKgbeky+Aq7TXy1J
+IBMuu1XsnPuftia79rn3zE2jlsJjH8uBsJLYRdqLXkPSTfWjmaQtaZzwbf1+4zw
kaFhXofAYxpNFTF4HMN2pUa9HdFG10Str3EFFBBmsCdaE6iVfaU2dS428yHAvCO1
0/lzcz2ucKg46LwdURdF9eN6EO9URYl34Gbykd8MTOOjW6P45Xd5SMGIMdaZ1luj
MPCQ5PiG8BoPO7SeYlfmbMGbo8184JMvkBigJ7bLNaohvU72BQWuaa48GE0DvDi4
w+Adpubx1fMtjuGzFDmrP/emQsIDi/fSccNYu652FyuHQ0OyPc2NTT2SrDTDtixQ
jd19NviQvLJMcySo5zDCVZ3R3vbGnUtZt3ATtHR7zHo6tfW/V3ybLHUyAy35HfcT
SeBI996REIEkckGhYthDVpsod12/R5AoWfS4IgEiRISK5/nl5BlDRhH/4BcOtB43
TlRH2FX0Vj15XQpAMYkBjcMkXUzI0zAirunmbQeVv5NSkZjBDkfsFQNkcps8EesN
geV52W4JGBOSP6XYX2L7wYvbtJN4pPm9lGP70enEahhSrmsQdfKO3wLUCoVWKHYq
vsj7K2/c7gez+q2iMLxJLlBCJdPMVps5IZUonrQBuF8R+W2MfjCGHrtkL9VsBUgm
EIkyvEaLRsD+BP42ekjoiohxR5QmWk899cLReXzZWcWehkFqyhfm7JMlBJzbRsSc
CUFS5RCJDRNOKnNAre+fn8IwnUlHbuy1fmG0JGYiogPnztphpwWSgha82dv2h5jd
i2/FC/q4+zrOiCYHTO8m6GOrftZyjDuNjRyB6pSh5r8SAbdUVk+rYgNfnpqZrlry
LUyKAc/bzDdNl3G6hzm07aMrI/M/wA7DmuGB1RRcD2Wxrsg2tfQSWmxfLlsS5a0R
sabuP7VodTQecHJRBUpjppZXFV+MnZMIEqjiPHyE3leJctBRhX+nloenNxjA13+H
aXFTxFiZAiAfglq6fAKr9heWGSuF3UsupruJjvwGJZU3kUV6ZEWz2x7F0jQDXHsI
CjNENWdKPFCSM8wDLE62AbbQPYTh27f7IVDjMVtd67aNWXD7e9oXrDjbYm2mXzFN
4UHUHzqPCHCiwoIGjZddoyXPXEgX8x+yIIJpwkyRrmyYgrHCkZn7H4EelRANf9qw
HSAUI2lxvHXuPKpJhx1i+JUAyZIMmmLy0s2pZE1UwL0rfP0LwBVUm6BYgLreiZxC
RlV0g7Zv+omSxFm8ExrTyI/hii1XjMUb8gBzGH+rAvv4Gu3B/U52HLWOo9feTJT9
fJlM4Aukdk7dbdQt4wO0Is5WAap86Ac2epgdMls5GLkBu5TYMC7jLF2sfxOmJe72
WP4MUQ0LP8BHEj/9Tyrve0REgdmCOQJ6VXBLi39Clh3lUzTKOgclAQgEqON1ElHD
4EEkvxplQX5Tzgo2K/kvqiTRYgByGT1Zna4Z2gnE67fygzRRFTpYDSfaLRrVCVI4
lEkbqHf7cAA44PTD8Ktn+bMe+NbSr8DcX1FdClokRYNR+ay9aeqARl8v9JJ8q0Ql
bw7DCfpv7XczXjIpaOCvIsQZU5cgoNIzqhfv7ta2U+FG/0T7x/SmSgf/iv1jU2x7
dZhrSlXN3NrJWXL4ZDVq01w62ws6arI7nigKESKEVxHOh135HdeiEhWvJeM5KQXf
856ma/H3JGDRIbj5zHB/Uxw5SE51vVpCJL9zMg/DSiSEdO4moDZm2nis3pPcyf7W
D2wPLuGddcl6W7y9gHi7rrnd+0DCwHbW3d9OPTNJrOykRA3um7jmePN/UmF8u9fV
j/1ro3ZVPjp77BZ1+f0+zPT5npP84x21Bsz1/laeHHKUYQV23FHpN8moeUwPC+hK
Rv1JQLVzb877x9khirqvnqSHV1i7g4aH2VyVek4uJhh7TfQ1NyuiXkqMH80dLRJ+
xPuOGnf0th5vCtBPxIocP8SKVE05VBDZZLrZi1FwS3ddhF/TSM6wvFvtufhyoLVv
KAwXBwozuwQ4QGSFBwYApWFVLEBEx/D8+05AxDzPSas0wV6pX7PoYLCCiT7BiXuC
KElxSK2iJWYHJjLswuw4DprXA8WMNtar6MElC4DYPZtWpC0qg2I8nP8Jdh8clPyD
v6C9uJwJ1/0VSFbznwxcY6I96BNafFQrbrHZhXPTX9iZ5JbfHfVg0Z6QUbhOa20S
b461DNM9SLj1OWoxDpc8xrmPpN0d4P0wrO4PZcKBtZe3NorrgWquX+9QPFVdVFVz
tIlNwoTqrRStAvQomJFDIwsz6FIlcfb+8XJkZQtEjMBftdaTKqpP0jdsOdxbD7xY
CeUDf+dNhTrGzQWSad7lu/ADo38EK9GP+f+VUFJ429NspatqX6sl6ipPU0aE6olm
vJWFSMuk9X/sXAqwuDQzBFRJ3lwg7qEvcRM5EqRtFevrlGeX38KSyoXUgTLoBzU+
XBL98igPM2pE46QTBDY/VHT2ldiGn05akDn7Z5s8J1x0V1JrYA0NvnogmFURJAa+
OdLrstfYVLc5Vxv4XLSXW4+fEkRQn8NfT5U3gd6Gu2ubzjcT6ioK+zthMvsbE92w
rjuabFEK4g5x+GFJ8GEVCZltt+6f1zxzedDN1bW6opM6gpJyj8emV1zdJoClNv4x
QAspJIf0O1mRoYr0Rj9kAk66bqCw/GgiRGepo+MXgF5GN67+QK6QnP2iEMYlz9B7
H6/g4SQcN4k1iq60rsIUsJRGt3mBM/+Iu6UJw5pMJ3Q3Hl+uGDDjBnbqFs7zangd
f3mmrBx8uKylNju5aq2yTrl/Ypg+8a4TVuRvDhhdJLjVB4Win3Zb+Dkxr5wmn9x2
3iBSgN9NcYDJVSkORARqyd8WWibeZrXxNcElTUHa1WQOkFcSxhgw3cifDUk+jRCu
ULWTza7O5LM1IZNs4irgffBE8E+EXjccD/8YRWYCNigitgYLA7+bFkaQ2DiufqtB
nV9hWnLIT8TL1jIG3UsSUY9z4KZ4F87AnhjAn7xqeVIUf/SwjQBKYA2BU3oQmN/p
Llsve0ZPs/G9c7hRztob8HevnmrzMIOhPyLFjmzzytmcbmrlvS6Mo0qqe2u2fe7q
sYWD95ofahvyc1YgLkRU/vAgurYLR8ZEy48y7+IXMkYekMiEOIPg/JgkvvX5BcTI
GnXJ+Ainnu87DvZy/wEDvSMYzTXYnhP5JjvPf+AsoOOrIlKC+fBuaPmmXQmlLmrU
Ew+/xD7dsbV+I42q7TPTaH/hwG+5jeuaMrENg5WB3DQ/QmK0Larp3dBvl+wZT7D3
fRZmSmuCRiIu+8kQKUkkoDXy3SGSPx1NDMOV8KQ03ZphOx9akzFaqqoKzsgaLHfu
nfxzesw7C1fHnn7FPkeEpeg2w92Wn21rIohlhTTF+QOC2HuPuTMPAy9Ujy4Oe+y5
zQT7V6oM6dq43XZSaRFqlPgNIhEfHdpL/Fo5GosgBMZIApq+mAfm+SXboNU/01Bv
+iAJF+goD1CTKzawQS/tN1Ugdbm4NEsPJN2fBcsrFHMEx0W96GAVQmPl7OFpUCyk
5v8DfdyjD6QcbLPLhijB5GUD9qAzt2AFUla+WLGULp/4KpaicMjj01HC9oZWpYJJ
+kbrIiAdyh2qO+KO+UKoNHcf5hMle8bVgZAIu83GUM/Gac5qTYYuDKVVjM2hg/ec
QXPJ2NI46/2h72gkBlUZDoKGuuk5huoUsSFpIF5mmG2dxNRYGn1lF2BKRqHYZE1g
bK2xJFu0sfac6v/DLomHAuiJjE8om08fsvSbT6rCq/UiIfY3SIRFJAGQ6cCt7Io+
yqroDDdY1UMsPegqfFkNuV2gueVX34ZuscduKRzcCDggODC19pdgiGuORiQwpQe7
EBXxzZZNIG+DZnOgjT8Sf36xdfxO5+OEPEbeiRWoQbXmULNsBvAODQTHalYqShVn
x0d/uAx+dlOwBnJsOIh+8fdGchpPZjzUHzPM1fe3W8VtqeXASL2dfw206TZOX5Xw
HZwU2VLN02RNZ8AuZl2j+mPwmMx6Ff6kAOqbN/iFxfrNpC77uwGZMTCZwKEuqTMK
OnCuNAsvtS2bCRw3NEULsyHwcFnqBPqH/xS/2QG7OJfK7K2FLuo29Or4qPJwwFm0
plRNw4OrQCaETEX6RLMWIoVQ5cdr9TnTTaXXU/mwDt9klEaiBly0+cM95naDnCqo
kjt38sBLI8MCIZ2DrE4bPoQg+c0PRiUhXwwkFLZqs8EpPy6k3rejxKBTEDfuNCiH
baSYsfXwFIYNZTn+j1PGFZjv0IwMbCRyYM1BayEGk8BRfUe2XpsIbjuO8CaIh4Bf
2HBO1m28Csz9YE3c+RqHypAo/+7CzSwc2Mw3HyyKmLN2YTvV70JjZu2zHUkYlhmg
Zwv6YHj8Bkk8ca/cV52owlYsjsIp3Tx7yTWqukFis3LGTrGlqy3xVMhyXcZvVwWs
0z+tnpfpI70CKtOpAyIa3tbVaYYMH79SoRbx+IETZqINwE+MsHH0buGunjpY64uT
qDmBUfaVcrW0n+LGekhgG+hVZ+n3OZq0oXwvFbZ55QaC5QrGofZBR+GyCJPw1UFH
xK46fVn6B3qody3IYRZFUHR4hyEMNnM4xxaIig4D5/cgj41hYxDwSuvf+DhDddf5
QmJj2cpGNRxVqzHwU07EyOKJbqWEHGbviFu2mZvw3ZNaYLLkC+5SbAXjuzTUcEWt
onhGZz0S1iMILPWO7q6hoQ33gbIMpGvySlOepMF6fOiDUWYLi0CFqhMwFYnlurZp
3SoWnlJmlnUs9hXXq00uT/ri6JxQORRqSNEA8cMvVsWQgIVkQ4ueclTpAFhPrgEI
N5Wg1ssaX7rM36WwszGLRGi8D0jnjWRanZK/DcmUNXtC9EB1ZiC+W4Z9DqUUJqvy
XpKqo2xQ6+xyzQpw8Wrn9ArLaM/A1+TA+bUnnwSoMmU5pbrlQV0UBT7EC2ij06DE
qwxyuZEOBVJ/gfwJ7cyyQ+M99wj1VNf7ahbTNRFoj0EatJmxY+uBunRQI9YidV2W
UbPLvDtnpMRQzIXB/K7VVWsyNd+uYpsZ1nHkXoHLLVGgmTPyqiHBBGPblkQkKAx4
CvSSoriBbH73jjFYRnjaMA0IHuDScztxJEAs83b0cY48RekvdQSm7WTqek25QAgJ
L8A1tXMAz/XuwvCF5H092T4X2w6XfFSKv0dQpMOOHvkIOPtvcMt4nZ5Ov5FAu96L
QLAZ+rllGEM61LblIJ0GzMH1pwKzdOG5T90HcsP8seydbCIdkjNWuh9OuGn8RULl
4yRFkhOVNKJt2UTeGf6ySsJz8KA7Uwb2BNqu72bdm7qTlTqYaZ2ceLd+ElQz9Vqm
BWkC1f4WPTFwdQw2zkQLfGeTtMfH5vcy0skbPBZq0V21iKJFnJL8ej8ms+oTi+B+
lIVo+uQjgvt05aS2CDO7jQrHZq5zy5sC6M9raCxUmJrm65zbaz94zHj/sQI1vlGa
b6HOhwxrIvbUqD9xwas/WXAkgt9rM1H72Qr9h41LqWx5TZJNmD+TnVQHfuCeJoU/
qHMMFilQ4srb1l6Cnp5tXNPJf9uniK3SzGuiqKJY9yeNQCAGTO7IUQzl/Ep0lk98
eELIHkG4X+iL31z7IDeucBMj6jNdx1qeGNQ6hKdotcdadmux9kE3OmLtpSwmHLmR
0kSagFNgOSrIN+zCV2sIJt/20DoWlzEQMif4wWszpJekPfgUyIvRHb6IKVrOAfHm
JUUoWCxN3iy0U1KaJMZT0mSiU0/CuNjckX2rGT9KYLOC8Vl1HtLyeMAPXv0L4j0O
5FDmkzFo61tP3bi+3cNaS+5eZ+wdLXh8wuMMQu0a9Itxg79BGFQIeDYWZJz0oAYm
sqhndQLkleNjSMF9t+gumMTcP9e76HOk3gtARTFBVyR8Y5nxTWqj7jMRDTmv4hWQ
sFJCoc9tUVWWKyrmYeuG/gcAyzhctIIh9Jmi4mGXvMtJTXmb8Cz9cIDaGfhBh1g6
Qo18qVKqocnLM3kfgM3z8D2syaRJBaBzeXXZQqCnHqxh933HWyInHhIVUUrW4r9D
h6YcT9XpmZiiRkY8eGl/h2zRvJpN3FZUATEjS1En3MFDgqzgkuHJhzYjZBsD79yw
wgl4VheeQtzvwFmHwvo5qRL3oPIE745MvaH6JJYfFSmlZYcC4XVV315FfALh5uUG
avoBSzJt41KXmlhnu2KJ7acxn93s2Js0LKer5j9JdS4dRyXaUwVTDwZqGlEbVGTJ
PfKNVLdJj2iIEupDwVk+Gf02lByWnjxlTsRZczBdgQiOxwzxUuA/neT+VBswrA/g
JN+4A7vnBLAWWGHx3PKbB3dSE+JTdl83p/QJtXkQEkik/D5BNdL+viysZklGr7Dc
RWra9uR55Awe/pyMMBxAI4tg3iFu69O2WiTqYfAP4izn29nhDsWZ0zBBe8fJp0+A
CGUY7aP7ODdHpoF6PRQyn2SY1bqwciGKY75Cl0uatlovfdp/PA9pOwfEV3tjDz4y
iFogQskwo9fGRWOZsg6mCroYSJodWxuTm12V3EvAEHmu1lZ/+7D7+im7jdej8Rur
fZF4+bz5jJA2cuo7L3KnT2JX4u3511ZkbjipKUAm1kHmE05qySJMKTbt9mJxqUwo
nnzMU/xLy46pTijjcmfnLNAXnDeoCpiSKgHaxmhxIS+Cu6do44aREQPIOKvMSfB5
DKy5DmhriUji/5tQM31im7lGJ3rxlgsErtrjvDs4h0+YiqHPk48aateBxE+VsgoW
U31Vg60AWMkRWwh5rWRV7mh5bCXXGE4z0d7IJazgQiEpJ0HnF7bYXGIxQKATaPtA
HLu+K3cc/vab87XFipR/ZYsaqhCB53/tDSHJ4TZI6Ba2QE+vU0b1XDisIIvn7PgW
06RdIaRQ2nFE8hXQAONhnwYfC6bH//vzmWd35ErDioAzCtzO6AFHuGgt6nx6yewt
ERscsqSiqEca1wGuNl2U9tqXK26mPHrz8cJNePuJyGB3mXTUJH5gkaL9LhOMy422
21Iz90wppY0hfNgfGlvXRLbsbiat8+UZn5kjX4QQYScEzcrw0HPZVD8F4MZXiQu1
ItwiNOv0IDLZuHclwPwgydEUgrRlQMICVq7s+JQ6BelGU2XRk8S7DiG/CwC8pPYJ
C9EH8dGkBMWb8Ou+ZwMCOF7oPf9l/exjXYJgQ5X06OK0QE+4a5Gno1gZWk1LVmFh
IGCK5C8KKdLg4WLzyG6WD9Liib8tqQi75+47zBbCGyoOvHexmGjfTfYXu7sF3e81
HCt71Y0vgTcKJWpN6EVx7cKF93YP2BGeLsh9sLELE2KYv3fbP0Ibrw7IHqEkB+4y
Q4m6ae9IoTUV29y1MS4Y9Nl6ceUFS8+rBsh0cgeGAT7yjcL98VNA/H5x8Ql59wdi
Bb7DHCyQWmIgQFv/6LMIkOZ+bRdZw4nN2zzNbVjZMdzTjoRLSHpRiyC4c3T3Zo3I
pmsrx1qYihM198XgtZzL2hg5vw79BmNTOuw/OSavNaIZ+GkjMVC5Div9no31cfkB
ZRF4+mQwf+K8O5kWjS8Jz1KxiKw3WIW6TPDXSzx3PJxRMaMPOQCD0+c+DaM1fFJI
5JRvnqN7YgYDfLlwclzw8jW1wmVouTZ2URmIbwxKrwua4lY5zrFI5SOIFVbSCxmt
VYvAUTUzHmO5ccPHmWNZYv4c+Ygs81511gUYTHCqnC+2FAjqij8djGN1mUsZLHk/
CNKQV6ONEqitIax8hsH3lid7nq4AkXNgWvNB38nSIu561mrbUwuOh91BD6sH19AY
5NO8JjKctjMr8tmakUsgVyPrKFHiHtHvd5slTr9AHTSEnqhXhTbvF6GF0gDWmNMV
lQFTAFiKyM/F/tMql2kJVMabdihR1kcMpyngv8KYMnkRHLVH3PAq1ccfwhfNoI3y
yC7QQe4k5ulXxupZ4cCjxKomhQ27AEjW2cD4Vt/ocDr8YNfvhXveDGdgeycnnwcd
z9FipSCPqzPQ/FH/8WsHJpe7Rjwk64+mEgAUwkQ8Cj3LD5/rjxeCGWZfrJOZYYc8
a510+1MiqWU3c9nCmkWZnEvoh1S7soP+rRt1591+DK+VNqv9YhPiLhlQgurkkA8e
p1RgMJHZm9/5+oJVhf50GpoDeat87cvW90PUvdfHxhKuE83Ny4CGL8vIRr+9Bbpm
8rAqmbIu5C9/+AGmYu5xfO4XDZV+2mrZI8c0XoZqhbqlTPMcxPJUyv53d/foAjGi
5W8oBOuFB5uB/R63b7IGe+neManc/MDDinCt9vGXjm+PW8QQu+E8Wb1HzHTlAbm8
joe+f8LEmrLnuM3B0c7hyOVRyEEkEoylYZQfgnJQmZT8uGhQezc0mVTXTcHZ3i9+
Kkke3caTo4zfU0SoWqw+fFcqHlpvelowmoKC8Ui8itMyGHDteEPq6vduLzmozdpj
iYxItqzqkNUmOVLqzs/r+Gd+GiUHMzSyXbUmvkTd0Iu4Af+zwN7JjqYhYV8O3KHD
5cj+Mwx0WfZ7YNZ4AYjyDIHUIF7gsvNmO3ANoSlUCsyBWLKnN51RFHDoh+5CiOqI
In75lpE54276ecDcw+AOykOzWdYtMOEjwK+Efr/D9vDYYIfY716fa41mUPq2KRaP
yuNNtOxSYImUdqTO4KQPQ7u+o6Pt97QYxvMEtl3IY7eSnY+94AP069b3HtkW3xe1
BEiNmbV6geyg3VJTet4BB2oXfDtNx+EitrZDNO36nMjntuhiRvBj1CTCbznjMJlm
p7FSooMWiF81/b2p1yixestkVodbqsftF3FE5o0N0335lLkN67XKqs4aEY+xYEj0
Mz4eK90P2y5cRWDPepqEhqU5s/uU2EowfJJ4tQtlhYDvghNVCfZfgXtLBs/H2gjx
KVEeXom+LfYJKHN8jMYyrwKl1EuWS5wzY9QtYrGtN58WaDMCCzyE86SuUOqjw4zV
PL7oL/UyMVyJrdpt6sJAVZdNHSb0+GxtVkaREY7ixF9cCXgGxcGhoqD/lUDVd/wz
p1f3sqxwb6BzKLur46TVaBz8lyRXI/7rErlxz6O1sG1zQdpsj1DOaAITTcqOcSDW
xwq0toHvz0LtFHR1vTJMesSBktkPfh4JB8Ixa0fpJhIEASVbioJlqw8r2gpKgCHE
QgxI+XMDLvPQw/XZuqpHyi4j/8zsAafZCjcnASXHaf1OCZi7LPnNq9ApEJl+ND/L
9MY+cGXgvi7fJnw8x7utpRHVo4hWjnEDmW96W8Bj0fH0IICrAbqP//wrrTG25YNh
w0Vya1muWM9wyDq80nOfLl+//9I6Nbk43XVHx1c2cxhuCB0mlWnbBgJ6UkRM2Uhg
xSW55rUuGbDbHDn3jrEtK5Zgf0ncE6b07xZ492ZZAHiWRiEkz/37XFpp8Sn4e4XW
EdAYbvI291uhePT/rrdqj1Z9BqakYda4QUoUSUWZt3U/q/ughlFUkZJwqFg3imLR
ArpBliMkQZfwqZ3uLaSMYqZi54Qfz+2T3JdIe3IrQPDlPjN90i/oMFE8aWmCgwdp
VGZ0jDUD6pNbeOraJ1+CkXB5EfbenuKRfvc4pS+lCGHSK0GcftWzrTuhyhpWFWbu
WujCiWfVwCX9rrLBeZM8gjyCic/aHHVAx/bm2obssFM4KGx18iSIJucdzwtgIWXC
hMghUfPiuiVXAa3UjVNsQqrp4igBvTwv+hiNAFxgohfSdl7KR8H8jlBquVnLIHzG
P6cr0k7z63xeN5W62a9LcZTecSKXbdBb2VJoXV7/gBafIUEzHALJkqb509XnQ/QF
tTxVyoDwQ2rTKkJ7jMk/sMIJbiF49YFcgttNqn/4VI2SLY9qfNUdRs/wlN2FauEp
Y/2YRgoCe0XNT+VAlLkeeDV8LL4IcO4RINQy3RH8hUTiwqEIpQmbZPhLjfE8AMPe
PBSrCjNwVNiojwaqF4L4hhMmEgheF2kpqzhul897/UniZn5jFDfYcCPeMNW7aFAh
llj3MV12iXP9bTT1QmokLXDWKoJlmDAxZplZwdoARx/5/txnY5OcY2Iuz8580dDJ
drI6253JIrdA/xz/bloUVk9k5xTcVC9m6ooCkFiuBJMWzMe2eg6MP3n9ExrlivbN
UDOOUpbpgaey6x85EbZ/NGhe5eLsHHw91FOYazuynIiVQR79eAs5MVbT8yFPEuhc
oSr2kNdkILlRJZlNHLmPRHTB9VfewpVsIM46Skppy73IDw2VF7peFlf9IRpsF5S0
Kdw48PYcU/hNfwR27vyzwnrAIiObxjFfEuict0MVNrqhGyneDDHZEz2JA+5ajDdq
Tu2mtNHh0GQaqZWvnbX0isa+r5Y4a8v3lnuIvMwqYy4HfuJquTxdACjR5ehquRmI
WFz2U5NUeJSeIQZrjaXRty/7dRksw2R/KIIn2PjSRtLaH6lZ643Zkee4c8gYvXWg
51Gp9LNH//q8wb6+HJC1zUR7q9DdLjxmyf6/G0y6uboP/ybJCG5rwVcNf8INm+Ci
4iGbkEiCoEQnz4MUvPikPN+gzV1Be6wipoaMqiIU0ICQDN/ANlrG9y2yJUP7QnDi
vEx6dcGFpoi4VEE+DdcUhUxcM+jYloDHNs+yjtxuLaRBZyFcHtUhRZ/ceK3KnXMK
EfCcOtjmRNL1ivOQDO5jJ7u0qqBcWPmCGtiaP1rrMOz3k1OBfUt0CZd2Z6DmFW5s
aLSwotR4h63F/fGClZjUR8UqdItVYiGpINM9STWIB2axuJ52Xj18TLC7GbXowC9A
BW+hK19f7XJ2mwSOAhHUlUiKa1fQektxEOb8W53jaXpUTYBs46hYIke0aDNvlr55
sD7X/dCLyicXQqu96JpL5a5hD8HF6jOSVXU8Art5IUJdP14I7mC6wy5MEu91g+Pv
FirrcbC9Kd3AvbeKx71yl1dfS7xeC/kvl6iZp+ZBZRcRT06MEbeBv0IbxBV1I7o8
YW0W5YHOVqwYXaxDuPcIaaWkzCLz7FVoS8HKUo2kbR2U0fDkNROHy3SXvHLhrrZw
UeDwuBd0PMlKSfD9yOMLKYm2FJDdD3Ec+c7FXqilZqWGxP1D3U4W88A2pbjMeGCe
UT+yByAsyq9SEAC6uMQxdyCqM4JBihkTzFTm363+g3QxWDapPdfEvsT/emguxjma
uTP3CbnESMshf1U9MvorX7KUrNDd2r24LlgqtWbkF9hOeNOfxJFg6SyyfsnXAlC3
MkVPf8x4XVwg9cESJDKC++Sm1MX5z5NkO62vmFVpb2Qic1yOH/HA5yYkgR7bdWIz
XmLlAZvRoWd4o6r+wYw6EOrLYMP4HoWtRUcu28PPG6KPF+Uc2JcyYO60kNoMpbzn
cs86bVyQssK25/g3Itw0LbEsOVg/SH/cb2be5/mQaPQtMt7CavQu6FfkBS6ghKzE
qCH3YYM5+E7mU98k4eGGCcBy27slA+H/DwCuTJKz6vvnT0y38WoQ+n3AzGQ7yIkt
5vqdvQOFu8P52B/By1Xo/HZJqd0l8PDDKcYmXIiNlr0yiN36mJrUv0+puiqL10Mz
kubaxaTEEZlxqtLOJ8Mz0CT+q6CgKN4KC8KGb2lLMsY4iNn4bZemEeujnHZksmhG
Q1Pz5oxByN2tSmFUb0cZb8mNQwDerlwmJwE4dN1h1qzm2oPBqV/F45FPfer5jswM
0WMcgDzxvhMTUpSQz7N4GIDXTAqvQD0jI1XUrBYN5ebpT0qPqMYT0FgjyoQhKCX4
QxDVpUYMGdqvCxy1nUU0jHSpGo6RfPNPs4YaTm/0TWNDiLCEGF8CHCPFlOY8SBHP
qxldWtt21wXslPULUCtfu/a7bWHoHxXDU8mj35cgnO/1Yxz+qh8p8GfedLwzjv+3
t9asqN6S0Wwbs0JroyRZdRlGWB1wjnt1h3pjFXiE5lst8UxsnBb7VBylIa8S/Off
6bFKH/hxomNG5xMW9FDNepqchHJ0sPe8QkV6kSUp6ZfonDiudhg7YHFwQFGZTMQx
fJ+i9wpbO02yQvBzKE9z2gWgQ//av1obq7cFl1Ffq9Hml0tZ5NlEaMpY8s/S/IMm
C8UnwTERpDKcj200tavChEMGR6otU/nDeeWiM7/AO074HEv3dY3jA1kNkuty6mIo
Axj3eulE+8pg3zZsb6ejSTxVlk0rWKrID0VwxUURXj8Cwgxr+6Ffe++MlCbezUvh
0URijZw9Twq9IaemQs8nVnSPtuEuY9FfT8NicBB1RdbsM7Ir6ea5Qk5yfmmgYoss
FSJWeZ8e04tf1O4q+cHYnEE1hL2UviC32/gxFKaOW1FRyCEESVvEgkdshZ5Ycgqc
A108lS26OZcn1xJxqjHHVPLK2Zd1ENyVQOIueqXMyiDVM78QQk0f+JiBGGtsPQWG
zYMZ4LM3D4TN6XuKn8Fx1TMeV+FNoqUByOw+YdpzH/Wy0QNvIanFkSIUg4WdyCR0
LFgk3JH70aCAF254ru06k3Cd/Ax2NouEFJuydNITa6ZZX1PSlB+vJl+e/hpX47MG
BdN5vqBfot+22Qxtfsl21xqKPv3weKKShn3w6bdtbgokKKS6lSlgnKzy3/atCfLM
WjwfozyfE9DUup+vaLNc5VkdbJVGes7Vrf88FJ/rrkRzFO2powo3ZBROzgpIDx4p
WW+QQeK5Iqsh9xK2cU5KXF99+NZ3LViVx4b/Nio/AGx71PDE5IYkFh7Rja+AM7Oy
GHk+L6zQ3KSSyLNOiEMOf7qycPgSIOdazFgC5ZmnTRb4tkBBnkTOijnG6V7zyy9V
i/mDVBBk4NmPGIWOWxQnNp5m9xT5fUyzmtQPuOVHD4D7Zf9ZTwe8iAh3IQllW5UB
mi/5WwMyL7Hv2qCQaKQ1e3o4AwN8DrA2by4JIBpI5qI7jLurFgeR2iPoFYyJM0ze
cMJzerZpZi+Y3gGsDmMznUwWubne5C6tu6awg8AwbJEQayCouoMWfNcfuVenMoTE
fkrmNbQNpGztT6V4vN7rRZr+Ed8CTEo0sxXanC2PCmngibZ9lInORDtrOnRX0tRr
3S8rdFfG6dQbc5Mp85U1K2Vg5PnBAiQHELqZ3Pw6wNmdgWvQkP4JhfVqodcx3WBe
ah+4Dnuw36UnTKA128G6+118QrzFzl7uTBqx6xJfCSjz0J64jXHzUfQ/s0pXf0Gj
S/QDu72LPgjvGd8Fbj6MadNA+WIvawG6jHCtHarLi27oyb9K0rb8TRU4wDDAdSrp
ioBrDttF8e1gG78AYljM1fHEd7JnzM2JbjPRcZf+Gv5DOhvH2w1XOkug2fnMtKbf
CRU8QXnS58LfGEIdHGheqYpI5U1NOnEF7AAbOdeVDNDw0YvI8oWFyeLo895DNTN4
Nq2jRRaDMyWgdcUglR363WzsUoiK35CrXxrvB1OXrF+RAtmxHfbS1KiX7dz0TWjt
j16kDpna6as6oTCUaBSgPTYNYw5sGBH6JFsI/2A+ik6AhM96IJTFdS4D1YLLQphh
SI6GYB1blRrFYAMU9XUjo4Q7yGL+Dopq5oykKe1F8panIpIFRF4cMLf5CTgiL08h
LFW4CeqiMcG0l6w1uRLteg13KVqLp0flumOBVuRRLsZ3JYtdFlp6INIfdLQg9sA0
KGXEdJoyHC0WRQi15/0TT/VZZGo35h2Ltmn8eARMFolT0JnIlhPA7Ux3pJawykP4
pEzG3VZ47X95YFlZ5YUwQKjjWqJQnbLQ2NlmYTaMEqcEukHtRYY8y66IlPM5+F9k
1RCyHWykqS0gFXkg9hpzdrP/t9Lj+sQXp4ZiwRzwtZcsrtkFC8tGDA+0cIvVENfk
HTvWonGvmtmaETVTEzWsGXP6UFCf3Y7WBeZc41VNPISprP5yGOn+tuzFB7JDmy19
nCDkSmqj97qgtLCSShsd3VXqcMmD1/yRi4nC1wa42ZNcyvHTx5TZzZhVmkFAGAe2
alj5ZGa+IeorfnsCDFnapvLpL4KK9yuUyfklU8GXPGy/phvlYn43MlAWByzULIwN
6pIN2dx7eBNrQum4AP9NQYhAqPpjvLy9Mz8gE0CIdYUs5xU48oU3jvFbE92h7kct
TNOAhvpcmKuOAa3SQlMQGG9yxEuxGxBGbW9T4kSHV1ve7RyOux+OUUXec8ajFdhK
T3mArfgA6yeSa5JXVwzjzbJtnEKDxbxs6YVa85/4VyCIBQOFg8nMR9V6HRvrRtup
dWDpnGYY1KBP5xEcWhCXR5sYM5zJjvdmlrwB1ruPQGCW9HnAYiaXxioT3EUJypXV
Ve5XnRlKY3C/yT9l8jItGgIuj8qnWTNCo8e9PqOmDBbga/MT1rycOnN54rYVL2K5
mzzXpIXYlOMRVC5ZchViqFJjnmo1Wb3dIz56+/LQz+IjGLeIWOHwaJUViFBP5amp
R9rcAq+fjfW5b6KmCkmPUz7Pj7u5pAYt6u540wu5rdMW6HLhAs3N2oAduJ6FS0kI
xHPg6tcjgIsPsvY6zaN9gIWREcihl/5uUGHdkvYRO4vEEObl8UtEDjiZ7oYeR8I3
/v1O87WWMCHPuK8TBultoDXEfECim3lGIP1uXFOBQa9fJG6Achd1kvKXouXpVghU
tx8LjyPGJWVV+awGX6qqRXnE6ab9hEFakY/NJO4o2yHCREPGR2LHSECwDOR5n8ka
nNrrqQK2foNi5dVUJ7pJ2dMMJn1xRXdLZmRI2d6tjnFUekhauOuhqSk07QZlCAUi
jAYhXl7a5yOFYooSZsR3FL+QU7c2SzDOGCu9k5YfXf76gj17UzRf5bqZCS1G1L9l
C4mASwS0T8ctdbT17DVHwU9K2O0WIeRJQoH79prgRtHS1N41ZwhW1swn8bWxqdrz
uukKsRAsxmd1QINKiovUEZw6SseMRs6m2tNAtrOMLDL3SjMZjRx0jfA/92P8Y0A+
UoiTNKbr7cjT4P/daWrwqD5NRRj267r+JkXjp8M984xNEKez6vhMBhJY/i/gnbbH
nlJRT/jEaPLoA2lzCQgdJQWrWcE6TfqXVd86q6i+aij70CqTUHMj69zpocKULZsO
83NFsCn5/jn25bxC8HeotTQJbJCX0rswSqt8nfKo88upB1QcjnLskwwiuBjuXt4p
2c4zc12GML6edcZ/dGU0IKMI0hoBGs+wzVm1Z+SAOSFaqIRTdINBgsoGxnyQV99I
9Z2VLXcF+HCIMQNNpIpHCGRVE8urcfJljz99+fe3p8gXDvIRugweCAJGkR6cunSw
MtO+YUDBicj/msdcN1KHm9TKjwUeJC6IgysxoFdEUSnE8VPR7G0mU9t6gv1A0+mj
VeTDkOQ0NKhSGw8rPAcFKXEGbgQnQe4oKQca8hcHlsZCdBLqckdMadQlgErU9/Ms
NBBWi1lpFg+eqDj/SxoChhgdCWgdrASvixvMBCqoqCR42bO5rzLLUNp9EtQyJCH4
fcq1iRRX42PDKPbquGTkBJb/FT5kF//SrCBxPWIi+v83xgoaK0SY6BOd2yHzeSrR
7I/YPKxkmO6J9Sfgb17/eOHNpMEj0Y5abz+77m1Gk2kmDIRwhLc/XMslSYdb6kJa
zPivQpQwD8HYUwaovcjQ1v7LpNktWLOzCt0zWeQaPrTMmxZU+SeLug88YYtraI8R
bBNOl50sipoTBHU/h6/EXW7elQVfpoQ3LadKXVg+/cHYNnxzDCrPwTJq+6cKsKSK
bdEMe6Hb1vj/lqTJOwEnHGoPpIY3RZ6HTJaCZPlZk1nq2jOa8Fvi9BprYtZgqFBm
2Nicq819fi7KOZT6oA1OehLidS4GgfMGE5/Oph+x1LSROEM8Auu4PikbfaWxyZG7
ySemO6OoYWRwXI4JmnH0sh3yxujH0MmbNrL9se7pqOBSVrCwQZASPbzr0tgVlZB9
9hfPbLE5AdxYBatVVnyQursXMHfS3M6hD3ts9jLLGbARqiaQz4dLvnvhjMsLLZJp
L3XaBrdZHvwNpGBSJ3Ct1tVeAbN3e+9pwLDQOGEZeZCdbywyUKHIDwHZPMh1gCLM
MlKYlPsYJTrDDNDozpBEg/BsUObDETc7kvmw2C+WIyr0LtP7dz5zYv0b7waYEwzq
I1zJ23i2nS25kl8x0C/gWQDoKh9AR5k4VaggdXx8CeO9dZ/oeonWuWEbsw9/Iur3
QAFhyXRYg9W6lOrZxhN+BBvjQxe0TrJv9VQyDXERBtOblozEpH5+E9+aQXVkxhXT
BHCSqnE092mTL5Y6AbbgPCGTCDkMkbQ16vj10dq8jKbuZn+7JNqem845IDtUGM+k
WzzXAJQZP3kNK87qnQn2NigE/qrG/MT9b6XOeCT/b3HAfu/lgLITU7xXiBPPfT8/
XQ2bKlSGRviki9rXxVnnBzmrDuT+ULiuH3LRoEBgTQhs58nzfUWyXixjnwhsH3vd
yufZZYsPfmYeOZA0sHp996Ry7Q2YWlI1Ik7yhRvx6EWuaIDV+ZXoCdoxT70M/NL5
bGvbqN8/UIqvUd5jy3F5xRvH86fK8iy6JZ9oN21QfxvLxC0wz5+jIZASYMRziMl2
PWCTLvWfxBXD79xIKFWfQCGdOrQTn/OzLB4KqBcQlgoGRaDGeoFc7YQDH3sdfQKz
AFoDSaZEKZ+TndGqMA7ryWfYqtpetIIUKM87bwMMV0k7m0pF+tRGgsiPzDuox8yI
QGEwa2WVx1/p9OONvOtjkn5ojWBdM/Tdx6B7aMVgy1JTZ2siE+1HocsRsCxVUslm
0XgtNgJAzU1cnM4jwFsLGa45EHtEqypFTtebqUwM6ilD29o3zM6HSTGPE1kR88cc
GU98feK5PqS4T8iHPr/Ndf3h9ThGC4tP0HkqQ1sNNbpe6KV09SHEQYWSQsW3Wv6H
Lp8GwHeO4x5TqMma2+tCOS2z/xmhTYuFCxab9URsUMZD4BQb5SCTZ3qSYzf3lF7u
1nvpa1QUZvjZp0IfvW5H7yhdwDOc+loiRb/cmwRgOGhUEekPmzhHcLzJtrKkOp0n
gBGSKU80hbSUyvHBCHIrIFOjPRE0ZhyTTQLgCKlAQ+5K9KDcy8U9Y1TyZw231ctY
w0A/0m92s8a04NNcKtBG7uBqyqE8C4PKpoKhG0tslfN/0hATan5DcVDacsbzu/g9
x5Hz9oaVf3PsOzjIuwOU7efe01idLDylk6jpKoSlTyXgzMiqyrkpuoMhs0W9lH69
IQBRzI1rJufPe8Pc1vCkCMLZFRChwXdsFIhZulB6hQnG+2bA14+h7PMAPGAOok0b
cMVf4SFi8v3OKU9BkZz0vXJ0JdyyeT210XNf8KIk+cN7nw9j8pfiqU8PCs3zCXX1
AgqUv3hzKeN7hlkFae/xJ6NC9iyKNUxunJLDwFV1rlaHpMKnFYbe/FjwHlvSK0A6
v/TecSYNSmSrf4LGVu0UwNt2UYjITZsLEUrMfWNbk/qOE/rNZHORimCcgSM+vU/d
2ZEF0pZuqc4P84gxFaCTV2uwYuF1fAMgf3Swurh4gRZQ9J4FoTWxgM81498WyxLS
Syj3hYg4CfTjWfos4FveryzxIBiWsTqZRRFmz0yQtGyuhFn2oEBfwAsy7Rde7s8M
c4CEaJ6wSjrxyhqUEH0wy2Ws+1yxS1j1QUbo6Z4Ne8GxrrQo3v1LxNY30OMezOtY
s0cRAJewIJuD9hEFCUmnarU5xcMdNRKZ2TJYQFUg8vCGQAHv6EscAo7I+hKTTy6C
fEG62P9Tq7khg+38S1+K97gPJx1cUa7mAyzGsbH3LgZMdLYVMskDpGAXM/whxvnx
8uwgrTIu07fE4/6ly3FYY8iwomwhIEbfw+1RmxFELsQGjtZD+D4kDpOkxoVG+1OC
V/ugyjQ/O7BTXGV6mExw+kc38vUWAmvUsSgd1ZXYFuu3iyV1rTSxDuWunVwUNNew
S6FuJ5O9yft0xmO9hZIWuQRijHAGiSKbsszPg75nXlV1a94ChBx5I1fr9XB+k1Mh
bo4Fbg1xA0wt5z+C3Qp5WjLgq3fh76NbyEfHSduk155FzkqZxvwaBFjd9gkF8yS/
TW6dIj6fAxIo/FDFfIT5zqTnvwp6B3KnA0WxeytvuHbPJ0MlnOMV6oqT5zivH+9l
V/pxmWH2/Zs3YSZa7xZgZ3hV/W/PTm4bcaJpGi+s+D1d4XVeDi/TbHsQGALg6XP8
YlT0KEf2iyxQT9/bFKHnaLOGQzhZ9fRMGF7F+t+wwLdj6u7YBxVQTkw/C/r04cwC
k49exFlBAHi059glZyA4upupC5mPXFo5/CXjMwp4jo58RbMhcl2+6LxqmjJx188n
tZSykzlHCNNpCdYDT2zrxolUEgCNqlYBNJzL90Ka18ihao8jnw9pEzmcwxrIZhlx
En47rU94y338M7ORxKrBRzNt9J4+ZEokD420lu7dBDtqoCaSQVCGptEk+FF2j75Z
ycRQkpw03sYN6MYJYhyT71cXmy4ML1AVb+8UKLn1sEzANvX56cSmgLde4tkvnE1z
pwGcxkKsw5P0jsSrIJIxbh50XFbOkZChq/6lSK5Uii3HmxvPgjiVEtloVRCtY9sB
h1dc/b6U0cVmt0C4fjE7YM1t1qQ8gXPd4sOC21+YXN0dA1bORNmBR4wXDTvapPCC
2eWrR80+Eso74TB1fZmu/4iwV/Q7GaI2/pWe3pJ09+OyqYeUUD4j0TT0iFdHOlKV
vz/Cc+EE1/keHhuHwRL5G+f57ejAhPzhJDJe5/XxiIAda68ADpFLC56ixAl1WwMj
UCiO+5l4tVWmoa90WlLy6XWMP3dRiX17s0ymTysl8j7A6bsuspraf8Gyl5IQ7FJo
23ePxh1IcdGYlFvu5BrZ9z8g6i0qEotul/+TwU3H7wnYK/CYwP17ke+LPef2KwYX
cs9YjYdxL8ti4oj9rUnAYUPFzLNnRRTKJXFDkGAUfsFdw+WBGll+QBby3awYZqPR
UeZ3NRVGrqLZV9IeSaNY0g==
`pragma protect end_protected
