// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Sv1TSAVf7nqNukRZYdX8iV0RgWhqf1KYSPn1pMzdgxRKk1ZjAY3cR7jJzMQeng2x
Gq2t0CMMyDN8ZOLMIrHUvICdgdMTgEHBjPWBJL1kDNr11OyaSJQhVsWC7SUXWFqh
EoF1RXkcun4BbzeP0qSRj4mHXrIBKT3PJklvpjZv11A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16560)
oXiCfeVlZNNgSwhqvcTDvCZNe7ga9hXCcaKnbGA0Iz5D0snDw40aRPmiDlqBynSl
GLXU6DkjR4cPypprc8lslRkZy7o5jF6qDJTXptDWX+9Tn07HbjuMem2iBx/GkCCZ
8HHyV6NoSd4HQB6808acCkYZR+oaciQTCHj6QztNa9fbRct6Pzjj8lAnxiXsgWNz
ePaQuCWg4wPw0/COk5r6kipQJPj/swokl3dTsMgrz/BiNNo5Ocump1LuhWLClT6o
dD5u0/jlCw16B9zhM74zKElj6WF9GdthoQUW2uHHSFPZWhZAajiLaQxce5S9qsyq
mb4QQHsnBIJMGTqmvfFY1zTT3GgAmRVPIrvyU1Oewphyel0+xqFU8o+VmqX40vzc
K6YayZn/86BxfrIFdsUS3I0P1R5mLKV6XDvorVjo97DQna6e6VRe1SH5lT0TCDfb
q2jLiISzYVXi3W79SBS0otFKxIRdLaLMkzcdqZil0VTJ0177YE5PGikVtOTfZTuq
KM74jO09Kxh2EG619PZzPh3LMFZ94PK6ENw4RJiPVyNAtATfoiqunwDE78AhzvCL
qvE3UNY7CBYNfKvG4e67vFmN9P6xFU0DJSslvr8tFoNWaCBrHJG3wTfZZsY6XfYL
r8+p3J/PRm8P872vUyQZbKeLwlrYFiVyTiC8GRg1dW8oGGi7/c+Mg/rRBmCnz8fr
LuB/Z/yoCSlHJ6G1mWIPtzl1OmRXwhBsrEi9XRnu4J4D7ssfUtl5ZAF7h0B0ufrz
DZh9Pc1Xhun8Dm6NWZmFuvdWYBWngGtRg1dx1l25HY0zQkL9T0/nI0lq7nKsrjs8
SnpurtHCA2TqbFl2GFrhvIdB6IXcEM+I3+tnBN+7gNbCf0JRJ6QVFKknxyXGR/C9
P1BppZGfIfv1CO5cTIMPgrwy/YpGHMi1Pa/jP99zLcSeFeBriIp/ZsIhYHrjF+Xn
GqNXkX2i3U4Bw/4GgbLWkGh34Z+9AAXtkdQPlX9WmyDY7dL1vuqOzcQiZRt2Kocb
o8LX+K+3y3TFVBPTYaxdOQTiOoYArV2LQQgzY4L97pCmskmkfqcJiQLURnamiO76
M5pojLwHa6tP9f8/Gb0QRtxXRhvxhV2JkGj/8xMIrSj+wfakk7J5qZjNNh+EbZhq
d1XoQL5WVBi4ocRjBbcvRX3CA+W9rL7e8JfLV1LL1wg1BWgC1T3AHEL/JB+gtloQ
1MhMek7DXMLAcbB9pQNicBKTwQkSyF8VE9YsqmbcRO3gv6o2/wMKs/sIj47aUCCj
ZSrFeOkKcvF6SfXBnu8J9eUTY87/rbUalIfU6UG3OKL9zOaE4GklYpnq6zlTzL24
PyB1GuiECCZ2Z5bcuhHtY26D/7//YrxJ23p68d+nFyU+7Znisnnj2QHs5iAPGccY
TzjNDNx0o7cLINo7DqUHskRTNHlMFtkqrKgzCX3zi8cJLH4IRINBDDywrdkmEo5b
l/LKm0bWP8JvA6EHWUb2y8D7AoAve+zaKVVzABkVTzF3qpbK2WqTWtzMmZRgVThD
ADBcJ3ffP+3h7BjMVZQUajvPWwnQShX89EMfJ4uQkmi0VWRTjtwD24DUd6gZv7KZ
lhwGPEAnLggZyJ39b0vz18/rfZoV5Yc6OeAqD8yWRHv8CVF2VW1UWAQIK4NpXW1u
RkyO2Kh2AmIDxf1UbHVMXlFwH3Tb6U857/7r/IlIJAHtgBoTo8cjFDelrhRoj53i
2RJriidZ3ZIPWVPKSnxu04WrQmLiXe1foCwGDjGg9DgQ+PZm4WZwtbP9CSipeOal
f7WZ7lqjoMRBtE+KVYiWWoR4xLmFHsm9C0C8pQnSM/nGGSAJMcSSisBM8SumO4zz
MwhqUyDlxuo7RmegxirpJoPAaf32/BNiLgXQWrSUI1/I26VGSSRSzgWITxdKBxs7
cltjRn5z4P28osVlXM4g3G6s0gN1haxafPUas0kF7019YG3w4PEAqn8bnYCsyXYV
pW7jq0I+hTv39s45wz95a2o7Fr/ogBc3EbiY4KhVyksd9u6zmC6ZU+7GV0Lmi1kc
iOP8eRIMM2BXkJWzjL3RVuEHkvS1h5WYVSw8NM8gctnPBvM6t7aWjhz4uVWph8xS
DhmyxJZKuzX/Ge9/gvO2dGpECYS8kkAdfmvmzl8HbfDUnwxpS0UxbpxjgmcZfyx2
FMKJHFz9m24JNVk9Vs7S6BruEz7XQz2U8An7/8BJxtAbtgL2hnXcPh0gbtznkz+B
67c1h8WZPoX/LJGtI4zHaFFi3OGSEt4EccIKaH7Gr448lxEeOPphNv0YfCP/hRnI
XOSmhDwMkgoOt6ezVhGGwCg+36rA5TulAulh7BpqIse6u8OQCHzTvbouHD0ptOBr
lVLTBHpDcnrkdU3nPSlcq4LttDcYdmGbgGB3QkjeEjsYvfhX+/U5P9sSFd5joeHd
UY3mpJ8YCjJL1n9FNoiByDWPtavoEjYjToMmPfDlOCWfsEOWBk9p8AXXldpxTacI
RZn+PZi9/4+Z6vh69797tutlbBfomUOnFnFObq8sIRLybbp5r5FhuZ7xM73lxjzt
p/iExTjShFVVRNbj9hLRLlgmnZISukqAaI/H7nf1iGKIMcjCt3Un/eUg+3w29RxA
tW6bcai8l1vwCtYuf4NpkdEhbuM5SvQjUK7y/2wZnB4n+EOTgrXjd36+xSyLY3gw
UXAKfvDPomyxGaT7QHi2DNkCSuOLG4heP6kyBg0rjymKULgM5P8G2xR0xmXMvk44
LcJhOXxqA4gXU6w1ViKZr4WwV7ImB9LI/8RgHvEonUATOPz9L0G+yQS71cDFW/DD
HU00zg/QlA2LcyMBUqDPI7X7oNWQdMR+P359VFEK2XzgFUd2fSbN9bqYfjMzyLHH
B1zNRnVQBnU3D6I6mrGnsfcUEMHKQQByWoqQgX4cxG/jltHA9NutKQjyyXn+roXB
6rTTYgkdx10f6BVC5J59J7dv+PEP9go79+S/X42SJQOhnkD6wz82V19cAQFqn3RG
749RWFGYKN4JIR6xHSznpsP2hdVkSPVB07zUvqV5mCp5EwpSsUz8iIM0tPGEU84J
kZ/rSMqPjrE6TTz+c7HXwIy6ddtz7TOuZiP5dojIyH+pfbE07WA2E5nXOCanOT+Q
czbze3pivP3nwU0GxXkivCCD90tualid5gyYBHFOlgvlU4PmDgfTh3wbJVr1U82C
C3f1rhibbCAVhH2CgQA0jKPzZAjLp4MmoA7i46UI0ptWNLz5w1ywUOTAn37hRHuL
FH6bAgMTzNs6EUQLMlOtRvkRGR5NkF/soy3zCo8Psh4U8MWncOZ1UNmF5DdHYbAo
7nHrW41/51gcCxsoMY6OAcL/KeMlBopiz2ypWbs5IQNjioS/XJyt+PURqcKNN+cd
+WAeosilcH98EVr/oxk8DJlfkAdtwYRJjDOxKym6dG/vFXy1Ca+3V8YlZiE/y7BM
DjddZBysIDCkHgRm+CgDqys+L651Xmy/KMpCi0Pf0+pdYiR/i37Yvyw+Cr3bDqdC
lJJ6FIAn6eQUTmdKgpRNeKZWBoe61yEBWxALlX42fADxaB0U7RuQfN0am01xjgLQ
9JUOacvuSndjKlaXy9dV0/aD2JsxqQQKsgxC9AWhCYsj2nspVcSlXuqQinI3Wx/p
v7b29BWAhpiVUjrI71Chbio/SB1kbhP/Dv9oKw6Un4myTfk2rVf3VZjcBPbXANBj
oPLFVz+ayBSzXMVcKirGJ3M4QMM27ECT9QfTLRm5W6MsxRTCcpIhvNqOE81cv4SY
F2PkjuIizu+uvUZmjFTvlxQa9g+0AQUFsoNJlmIv35ZFm1//IuYLE+e9SgFKAGCt
rx7hn7IOtt17c7u4aMggx6DRB+k2o35eKGiZ5Qnl4SobTaI2knaSirM3I8/m7bA1
a0OXAHneADyRWusXUXPeSCgwKolD1ASjYqWDt/+FcYIzGRcTAxg6TtYg3O1BAg1c
FK7grNR1YzRt9TgUGV3nQfkr4LeBIMlqOmXRBwrJQWlLMjgAQJ/zHgjzVkniSEER
HslPSA+/e6P96CjnVDRE28PGNapmfjUTnsFPDvub2TpNd+zI+rCRtSaEF/sPaN0U
NIVnMUuuGIED3NB0v79InaS5HCc5z85lWCcNv29WsW3q+QxUIBSPsrPeNiEJlH3m
HdUQluZU6KdLdX3mCbYfdMnYc49n0eAMZa087ucme3tBFv24GkW5/n0XhvZiwqsc
wHlWk+GZSRXjgGjGo9hcb9dmB/OMj/MtWhahJrH+accRvr3KgO7rAddAmJUdeUUf
KQkViHOsZ1Syz49BnuM6uvb1FmCQq2BPhVvAXiyToKqhdIfB8B40ETT8WMs4WPHC
yt5gMqNuf1uUjHggjHwiGXeaY4gpuPtiHkMdba6WbYk85j9VQv/yP5xUfEjSyaVm
Xgvoglb41KC24m3BNm676YtD8VC6Gkbc/Ew9Ym1h6q3swbLibggYNEsgPVEPa7uR
xrrpTmq4Ap3eRxUGKkIF0qjB8/VOPATtrgW6GWNUVgAazCW//Mfn6cFIZTxy5CQN
PJ/bUu7cGAfykkAnzYI1s89yU6Lo+5jjaj36AvK12H5nLLTJCixQqGJSt8UfQu1I
lf/mGx0PPSB01vIQMCGPuodib7H1QtbtvY0f2zJseKE1lTrMdtTdIUZNtwrPS8qp
3sf4hsHA+4tVG8Xa2Y0my3Mc8VHGRwyYFgua2HiUwrg2h4iujvQYk3AkuSp4Ppix
NxbYhfnkz+DqiwzSh5Tk49VD5DxpTLwfrUeXg9HYT6pvx7SW6U1ObbodzS3dqUd+
IzPLKxJgElflJrjfeIFg3C5gAZh/Xi+yXMt4vkWp/wUmS/AfXqJb/crwkfQ4u02n
GS0Lcdnh38bhgIpUEhFnpwj6DQeOnNJbb5FyA/6rm+38N6ZLmOyXLTi1GgzoefH2
E9qe2caZsO1UGjVw+gAssa7cvgyuXSX+qWWziAXbNizNkqJluSVnqZyfG+G7BYRZ
2lERdCoOIzOfEEhZ/UftZ0+hSU77i4DhlYXcg/REpm5k/BSZnpCbr5nFFOaACzdq
4pwwmHRk1T2D3ByuwrLxEWqyyB0WiotRyhaUFdxhSZBEkmr1nVI0ZPEWggzKJbMv
sfYuFn/Fct2SZIDQFHGPTNDVFZWaIWBDH5jiqnAiSDoiOlQfdHP+Wud85bBsOvfo
Hn3EjZ+i4MwiVPV+XSIZDd3zqagTD6hX1yN9HdnzD8xdykQvReHkP126oz0dbvVj
ZwtTew9glM5YVWQpmJJvKWW3ZPThMVBL0edO1pUWFGrDxjWHVim72e57ay/TjELY
FBlU1hFWkbg2KAISH8HtHwHKDSLQ1ShceYsmTb7Crw3U39+N5BtZ+6yjZiIH2huL
TtA4FpB5e0Sx23LGqFqQmRWYRRfgF3uOJ2340R7ZNzxbtqwJWLlAYEDuMzZ0Y4k7
TWCE9biPzB0D8Qs1dH3uUv9oPFjM0bXa9Af7yUYYH1sryTPRzWhErG1IX7yOaRH9
Ca5B+rxpwoRA9c3EogRRNOu/0RGnz+4xfbwvCnIinOZNVm6K2X8B894XwzX4IxjW
zHRx53Y16Gdn4T9XpPC+dJyV3s5jI4VGic/LVv4UqDn/qE/GeNKKZff+htI4mVk1
POBBKuqERp5nQ8PhqNT2wpfFPTTHvvcIMkveuK+3pTgLnX0Ce8w7kE4bTilSJaAF
xc3svydVtenfD27p25DmrnmySB4o5x1TaNhbLMEo5YqtvMJ8J3JjyWsKN9MHw4LW
2W0EdgNcrI7NuUwK1Zm04ZMipanFAoAQBn+vN6Br0neb8diDAJgI179/XB8qH3gu
kBF27o7WNH3yW0gUSzTtIqq5ZlMpj/NMQlcxt93vb/XvmTnjDGmRZT73A6WPfmn/
7RJvtocbvgTqQIheqSF1NJAvrD9VLOfihCNJIpb2eelLt3BhggTUOoVrAx95EfCE
BCPKSmrPBIvHywOd98w6bjBVrFaL6cnGsoQJZDCZjixzEJPbRinJMXBfhTQCKPjz
ZMRZISef5vJ0HWVBTfu/X6BO4zGe+8FBWNfEa6hkE2IEAmWoGQOW5cow8R6/LY7t
fvwdQDzJeu+DwKbiVjdHzz/0/21u9GCM7WIyv6snviCeZOd69xgdyvozdCEA+huy
+KDkVuCbPZq+MrIFjgOiOLsPVh/OJL5kZeN8+g1s3eA6854zPGmfYGZt+I15d2zL
zotGEDcjl3qUe4Oks2r0s+bdIabL7M2cnlrI+VYboC7eMPbhCd4hRlFLqU9GGpmU
OVvXdgfvU2KzOpLQIEq2rqmyD/7qAIirXJB8VprgLZq2hGXjoVft6XNptv8cbkKx
AnfM6AxsaEIpB0FmaxHesja4KCuFQwmyNkomEtodInauNDiIRpgAmeAGN75NFjhx
hswwcKn5abzoAgXf6RnYFWk8eiOXxk/PEpDfFRQacx/u8PjSEou3u6DbJX/wXkPa
PwZmNmJ4fdw4TaXtWM5S5GDUV9oH65b1EqbOqnKXXweSjpPmPYjtRjRVFBOynEpf
OyJPyaX5XLW5yMg3tcHg6wMRbnxqRbmmZ0pSgCSijqLnMos47ybM4SwkrBDVYDoX
L1l2+zVejaEN106JvF5ihpr29eFcurC4FwChfzyDB1/ZlXOT22dnrnrbS2amzX7i
RfqbmRZN8UrRqh17sbOsHf9xC/zBEvUzPsSaF8/sFoFD/1ag5+o5rEGDnHCFIdA4
zkjIw93ufjiJdQq4rs3mQSTnXR84dGzmt3Rrl9Fa5T9xi8bgCEmKX8BMqRJ4hojQ
x1M+2jjpSom5YDT7u1fNgQpGvtFT94kuJHfQfDRiyDP/9ePRRkzDpmo7qFQTmBFi
YUXgnht+hBZR73kVLRnT0tHtoUhs2birL4M6cED6txX4LJ7Se9UH5830USAMFn8s
/fkrb1YyxXOti4ymQ5DowTSzZheKnPRekm8Ru3J/Mb0Znz75y/34SSSc6oa0qasm
xmZLDcmeubdN/SODTqI5n85b44SymPj1aCXkqk9Lu3SOuQfkYxoWt6N5gHiJEglO
rV4b6zzPUoURQ1JL3HCa/bXTvXCL2msTznHD7edkygIwu0tzjMWAOj1inNU+KqnM
hyNe0l30ec3M0eR3WMwYqa2Bj39cG0xq18fZN13Nl+bG5DLAn462e0tGMwlC0/es
D4751Uo+Cd9zz+qj/Y0XkWHwhoujWE1RCPSfozrDY9q2Ud/bm/xxsHheMbP6EBe/
HhP1Qg24z+xxz537uqNcvHDG8Bf0HuBalpEU+gnztWCGgEOhUAnLSWz143HcNyjf
a4WRrf77rZwcPleEGeOQ/uL/A4A9kMcy0HThBMHjaQzWoAmEQBaPm9aUZDNljq+y
rpGXfeJEL0870PxQHmYypEFj3J3XCu2Tlw/olkFJ/6ItmOqpmr+SJrFqre2QDKut
OsEH7qqcpuTM3s6UsP/gD5CjZHN4Ev67qlupu3dJ2w1ByQLGutQh1Rxt5EX819XC
lKxYwDIFhDlyLsUtrxE4ABkHeUAl12co9xFXc/wcHn1LOtQGot6QS5tHOhdE03qb
Ka4fv8JfArHReUwH8CvyV6xHVjDttgBGsUT8/Sg0SBtSkdzjTWGl2cT4Frcs+O2L
Qo2fZFwGpnJ6NK7Z0w8WY1vWiE0cr8JR9N/YqIQ+kLOvjTrXDGyoCLjvWSvBHDDd
9eH+NHRlI9ciiP80ejGh3XDXC9MGcgynaKAzyz3gFupfzLbrsmxd/+uZtzCweS/g
cA57dS1c/yZqXv1Tgtq5EcpqQR2ddnPWgvOSprsrdXTa3mS/WsxtcUDasynzLtqx
zxfBI1ydK6SBsy31c1kADsHGxPc2M9wxu71kbo96b4fIYZgjbw21teNurb94CgrG
egXLXVaRkyB31LLSMyRNme8Q5rpyL7l7qXYHprtciU7NztUrBkxX2evJDsKEnMcz
BXvdqcH+9ZbcGvHe4oCR3YswnuAZzma8VHiq7HFOoGhQXoBEd1JsWZvBPNi48dmi
K0Ddye9ya3ZwC0eIQw75F0jXJ+tAWbQsWf9b/6xDUoUXvr5cHeQ//5tzeeuXTTuc
2igK7TgimEa9MKHUsETqAoLt/myi4IwIQ9jwk+4SHhLdbKiFGhpJ07CAtK0dRMlK
Epr1eoz6gkzVkt7pC2OB8Bd69OY79XxiX2JNRrZImiFzzTWPH4esjc8KFsNbtVoL
0RgP2WZTviYvcMvce8J2uX4Pud5rE/8TUeQQw+hiBXXdFGR1wgPJw+yIHwTBjrJo
mIB7/DcoeSWGV6NKv5CauSi7JBTZeq5B3ZsW04nmlY04sOtYt9d+w8RKdXTOg/V+
Vjd8mIXKjdrl+SC5iv3ip4e2v1A12ixQ9U3tEhI9wWYu5PPkOoz4cd2trhtu1ELJ
VXD8xJ5NpMW9Abf/mekyuiypPSil8dRVHv8jnhqRbkH+p9El0shUofGzQncADadN
THyXL6x6i2QXPBvA6+0BVMZuoROpkjzUz6HBYGbwmBXwy9Vich+su3OZdit2LuFo
KI02+RESChGN+zRHMPmnI6ZbLOxbiwpQ5NTEZgQfyVtJAUppwuUy5LInLUmUq6Mc
dkWaqzTneMVWgiOPA6UPPthFzPEL4YMo+RLkpvYVvTMSSyr+alHa2nnw2hv6Ix1E
XAr3KFGJUNx/ZSFZaMqILNvJs9f8jiC5DRthN0yxp4RN4jqemugpO2ZJwukZxCrw
rJAaI9KxIoDflGv1jrY+vJ3LZX92D/29JTlk3BGDC2C2hnapwhePTPvcVmShpVzX
x442E2sI2/Rmzzzc4L2i85kuOE9LymOWimKAeOxyZ0sGKe0cl/xdu4QtkP5ieZO6
/qS7jMfdCUIr1ofmt4vIFaHYxU/Gc2ACFOvAdwiHJ3fqpwbVltqIrFgvAeEUHDeX
lo8bhGPdX6tuFOcxUhCIdB9ILm2rcGYunCOlrIrtsOnpmupTD17aFt4/zApt2Wwt
IXABmAKUguZEFWaGkS5owVGicLakqLTh8TvTbAY42bfQ/5+xuBHSzuGiFqrZ8XjJ
r8M6iBFVQioYeDD/BMyt4wOYBDNrhnY9CTpULBnzQggktH7cIgikGt0nNZp2KBLO
A9yXoRsUnbfsYgNYS5iTckUYmH1YIloi7PUUgJvhKlMW02ZZpCWVda1JnMI75Nwf
a5r/pWulJMtikNlUPh7jtQ6nmy8Y0HzPwDjMCYTuUyBpm0br1HFfhdmk4tyBKuy2
REneeM+WKSBrjX/KBZ1P0yQVsy8I/B5EdXGgGgb5U+J0TbzT6WvT7aQnHhy6j4Ua
yOastPz7yrAZEA1oiyHRjQCjQtTTCi8EUU6rpEOUkzSVqaTbLHmWZWKluvmF5gmr
55SSfBw5NOIYkJxwBdyGWt7JxhIIbqUoKgLigxQpg2/GwmTbnW4npOCXSxAjXZEJ
ViTk7apQB4MyXTq9orUsDZLuBJH7OlHCfnKjIaGpCO2zTjIDvkCFVOIFFoXp+X57
WPg39CmKkj5F3Ah16E+B1EumWo8/OscKmFVLYI7DU+I9e5Xq81mHvHIrb8eroB1u
jVbM544CH4hJvfRUnRN+9YaNKGlSbuyeOLtrEktf+64Fqz+rvmZSesX7xfvH8mka
02XMflYsJKZ7VD9rVwPo1wZR/VhkSAf9CL6ZCuVMWy21Y/2VqGmZ91iX6UzneMrt
w1nmxtpsm6Uah9Bi4vY3B0PEl2R6FeR+FvWSKcXvE0SFZL6LoLihx4/rveRZGjjp
l7vzyYEoAnJDsPtDsdhiAH4Z6XngpOKA8lslSNboIOBxJtVo18GiS8hNzC3GCxVB
lu7OHX6Qcj6yBLw+nHBJ2vziSEohp7aWZNvqpNsURw/Owe1xTTWiC/1uxuNLnuUQ
26bB4LD+PDMR5MZdT2H/uWZ2HsbTqOYQ8KWop3IdUu2/In3F9YhCRKsgEgWPR6Rh
0TSANDSWCE9pWzTg8s2sb0C1bFb6DnQSb3KGi3qz9W4+l0LsdfrqPVdZpTSlqroc
rtcI/Wtznb3kU+BIei93gq+lWgjUh+kIhd1C2mUJDLs07dIbfig/flGYbcpkO/2i
0Fb1oO7YI6AwPRJAU3A1gDjDQ/yqidk0xzc7HI0T2dvR+fe/A3XvEac//tiDUcms
Mi1pW3Gv8tRsO6jE06DESdecELGjDlPhPWOfOsTw+PF0e2LB31qChUkvDbjRoVYq
4IeUkGI0H9/dG7y1NWm/o2plJfU9665JyH6JkxeZb7qb6OrFk8tD/HqSo1HbkxZd
ohtM0vutV5Z4wi1UJPdgPFNANMgs8v2U52ePVqO+1tVhJ1NaIC0JGrU90Oxl6KET
AwaVBdw59Ex/e/k94dhSS8HL26rIguLduekPEsrxjBFAB/RATNeCvHHAQnLYgQuz
wRncL0ZhF9UgUYtdXCkosYeUKbp7gcqWSWVa+5OICTu6G45O0BFEJqYn2KIBG8/t
GMCYtlDfxayfypiDv+JsF8gbja7AZmo6OclQ/Y6gFRYWnk3+mHti+kqFxpeqc2sG
2xJMBGrACXzQ2ZbysHjSll2NcRMAQtyLhsOTht1YDiqcr8QzF2cX/NmqpPEuAt7t
DXkFFwe2d1AeTU+zlT3EC6vPLnxEy4KCokzpA5jSB7ssIXgjzbKB2cT0SznxJGt2
lLv0lSe8izkmvi9FuXX9D0EjcjLRr7/ZRAtubvnULkZP1Oi0wzt+BsYpqIp4kOjF
vq268r3iRHa6+cIco6cbpBjELJVZQiR/szbqTMkLEU6B8l6PS33SoFB/EAI/vqRQ
BXk/V3dlADIUCAcIKKVMQ4kG2Y2dsfs6DOl6piYPAnYRzZi0QtlFshofNVPdXxM+
IyvmAczGTwxnejNr5KphNdLPJEDl61AsAPz+0v9BQODLaozHqDsiUnSlBU6qkpEL
PGRhFaG7XFUwgCPU/E6Ss16g8nqQ61fSXvpTizUa/x0FHE1Xwaqclb3CKLgklr6h
XPS8PzDhtLi6emTuD4vJLuhojUaFF4gX/G536DfS0TBISeYFhHaO9s6Xh3F2K+hu
pXuyuZtl1HPhcO39Mq0tkoq12hmPJ76YUR4v3nr3xQENhhvoWYBB1dfeXSs3gjr4
nTCLf5tunq34Vv36sca/qmHpxlFX1a8IMHmiaeoDYHCpOr2/lIJWiRRBEviJ3b1d
r4+R8k6lf+DXrLu0J/N84Z4PCvNmrHsV8eaTRpT5tJF8Q6j8kof4yPzm2t3ky5fY
ZUmSC2sxjtFS84rxFifPnYgmZeufNyE98LXE1aWcj8SehUT3ZQ9R6dN2WGTrQdy8
T0B0ic5AeSGr9tro/H4RHBDeO9jo9VVrv6uzq8V+4cNUo9bWLRlx47g4We51cc6T
aEQnbiQ5xZLJInou/bNMtZLWV3IBjyflZoFUMnHLXj8P/pAWkIOkLE00FZTEkrkf
goFiiPd/TVmy+tDDvLlf4QEPHYHiID5+ltOPE1n+rkfFcNwxOfTpYgw7RTlCrEb3
39l60dJBGOSQ60/aPk3Rv7jc5vuoeidJgjtW/SHpeLky/X7C0Y1j3Yjjy5EpPqy4
N+ZD2IUgeeEf3vWsAjaue/CYtfLWr8nDr6xIPLw9aGWSlL5muRzCQpgrkbx4+FZ0
bkElyQvafVSvsAMxEyU3JU4KphfImmyP/fZgmwUxRpKUG3yYnx+csjBo6LLyPdpp
zYBp+ZUdAvJgBcaQXybZzm6mE+2ZnJMKRlNKzhagJIufSzdFgYVRhvTC9BQr/zpb
GIzp9VCcGjdgTueX2apIWFpjrJzcqVV8CXO8qSctOmPazTXl6Ja5DfY7QEy0tzsl
RRUz+b0hf1sexjA7oLLv7Wh2OWUhst5CwJpy99QJ4P8cw6nu/z916Y3kpGlRVlU2
yYCz9HnhpFHNT9Aw3jJ/L8K/xBWAjmmp2bNwSr9XHswwtwlA2bAdOWb248peUUeF
/QQ0CBoRU2C46asRhx1S3JJaGa6GfS6xD8twnOhu6FXSAxO/O54L+2x8pVyb7lza
viKlxmOd8/sq4U0Nh3MkFoOsEJG6+84uGS7rW+qd71WuthL0xG0YigtDWfxcwmDZ
hx33a1dmE/JgdQjdgwhcSwTivqrVWDvSzWb140EE0YUGr+TQ6JbrSZ+vc5jeb4m1
sTW9KlGx7jKb7mTQxvxge4cNI3lO7aSY4WzwXdhfnhDaSQJDxcPsEEXQtqmDR78p
sG35NA84ZkG7kyQUInH7zQNl2YZNDXRni8EshxVaJU7ULXsVF5X73iVwF7h3VDQd
ZsZMfCxcbuqirxOYE4RxActl+TPGKCu4EC3l7LMSE0GKcFKVrfQOg1SoNowZTTKB
qKWMeDLBeOm5mAbRrQK6XtHiUkpDDSpS5dtUFKmsuH1gOWZvjr1wbkb5AkrAiQif
/q1jn2IQCtKKyU1ffPw6bJNzqMhzqHl1Oj4Sbwh6m2GumGrU5ShwSB/cAdnq8GBQ
2445OJbXjQ2TKqB0aoAEF9fiWLYCuxqJ2I/wmumoSqZO9v/BRyimjkKpM3YYWV8m
KJEImkmyrKcrOGvfaGC/BPgculRj47g/nXzP8KUioeNlT7ZzwQdGafdfiUn2VM1f
18jZBhwW9oaW1e92xy40EOwlI2sUKHNi4vDygQ3yPQQFx1pb62AvF84RG5f8z+a2
DbO4QTJSaHTbiGjvfgEGZGOI/tejTi9zc+KDmIeGTMWi+vy50uz3PIfwg6BoulzA
LBYWHyaD4CiBORfETi7shreJkErDws8tR9iaxMgHPrdG4kT2FixCon/4UHdDIO3m
Pw25ApKsJaZ1ydgZ/UZrP2lVsfM1bqWE490iFpVflMd2w49AnPV9sl9Q9OWB/Ypw
rsuQtX2UO5sjdIw1ykPI3Iq23eYgg6zFnKWuj6pcgLHjtAUH8LwgcnrFVog+CMLj
A8Y4xVZ/+bRycFg2D3FNpPTXeDC2ofBKr2bryz4yjyaDb16VyWr+X6jU0ULc6bA+
jmTmza7PuXOGyQxQgifAlzT9V5rux8klX3wPi9LKkf6xRx6iSKb6T21Ui553LLJW
KhkEBJ7sxlGV1Aqxd0m4cNYJgHgdwE9vWJNOSIAMCZT3SK1BIwMye0/3uFMqL2vj
fmEPCoXk7Jn7Z6LKy6SKQvOqwECg2NmqSyv8W53YJBNjlp2oWPuhpHaGz8VYfp2G
XwrnuimWNYflrPCwiJnZBUo3IurlLXmhJ4zhWh5/14fhSfVCnUMNBVAYYnSFr4z9
R5jXUkLTkUx9pZEZIQVdvHTm3IJ92Fy1+b/hEdg8WYQhneXEn7KuE/EVeXDd36bT
6aXNIOJ6g3T0egg6WDwiPSJLZb80BC85CuIQQ/mtICEtst+lOkeMBS9uYtdiOHN5
BKoMcXcKVHvghHvbI7inHsd5nxPB+0QojqKQHceAICy/K+Vb0+d5OONtIqTZKD3u
sH0mZq6OhICoj/WG7s9h6ufCXSOfaGt1eTbNOeEevXtrUw5wzDOsS5/5h4folDG8
gpLHJ6dAfXdvxptc+zU4FkkB+zdOQAURZiUIfcBVuMpxPqQi0KT2H7PCOVPJq90a
kUE0UO4yq09n23BeZDERKyH+ayX2+vO8Py/4ig7W1KJ9ni4yvm4Y4P2Nby1pQk2k
AxuVsPIpXV5Qf8MNRlRyCb5zyVjFDQAFG3T/ejYFLpWv1FD8DuWBx7HjWo9NZSfg
kpUTe2Zev3sb9Vu/mXYJfaifvLnP6CPVvt+sDhfeZcKjfRkeggpdnMyD64yyT/yU
+O8++W1H71GYT2Ix1zUC0no13AsTnQbfjjMEhw2LxgiIEBQPxApy1HYpdTl+C5q1
mtOZswWGkMDwBRvyW6rHPO9JdlCf/smlxOjVSJC3hX8KEtuAxjhBZxQlLu9i4WeP
TZ+vWyKwM5uT+vhe3GhNK9+mxfozNAebV3wOkxXuBt9kBkqe3D8NHZcTWhKUGhh4
zzd+29Xu28B0cpa3ZVBEGmy19rA6FQia/fOIK9MxVB/aKyQoPJaj64uNdOk4PCwq
npjIdKVPTXS+gvFUXc91YYO/ztVsy+DcIjoKBS8Fc7cyD9Ok9/ZiRVajih+Lp27n
T0gOCrCxbDRIKSLLiCU8Hwi+YIZNEfdwH3Ed+PRwRPMFCm3nZkltf7mOoZGTjxyp
V6myu7bUGtPlM48/CwBQeEf+jp/SNJ+JtXwUCLej3Z14d9WvvlSncZdjBxzvOiPe
bI6GIy7Vxx309V1FOZHhY/Udw71yzjRTRlCZgI+ut2x+wCi/EvSTJ2NkZ+5Vwhbn
ycCRt1/IYKifCr1HXAuUzIm3nJxNclAwzSmYWmAkzdxQ933WiRfbHsmXuHE1VhqC
ptm1ZXEUUe+5+8+8PCjxylq9jw6oenCd+99xNYYv4G7zCPBC8y3l7q8em/SX6mhh
6UoHa2Af24SgAXlXP7LEpZedNwehazgWT2SPbBIIoEpCbC03YNoiDNuwwXYehoMP
gYUuFZJmxPGg5j+2sOILLFZoQO0JxHwJbThvlJEG5SNE12ods4m62/+S7yqqLrqY
/9o5a5JwafmeMueIVINdVOya02ezJo4RSHizOvrxon0m5yh5P/xGtsW2XPspXbpG
p1RcWZUr/xB09/8r+BoxXH3UT4CjQlE0o6lCAD18QjEpIRgXF61O1ihwX/VK3Ugh
NqmL4Uu5TdCMGAYdO/koNzktE+K2Jxwiup2LIR5WbIZaEVpHC5OJR1UMtOYRgkLH
WMIoa4FrdN6afuf5gKT17lCHe12gKFYot5zesMhyTBpkn8tfChO8g9kSvNT71IsF
GO0odcemY2t2x1Infaz8T3duAI2D4gF8n8sJZZdA/4F1NbOV8XYOiIBjvZGlhBh2
zrBq7Tad7iXn11hJNN2xrLYsaSDB+Q6h+5FUXq1XtUkfimz1HyjmYBk1IrFsqUH1
jqYJsDo0FxBJ9XhvRfi2kHAaf+PGzZPxgHpUheri2x4C9xbJi1VWgzJmN3To+6gu
WwElzZf7VhXAigteLbCfD/0bCFA5vlqWM9LfFonlfLPSHWX3nCdsBPts83BX5uIB
802gD+1b9Zhp35Tj1ePSZoGvk5ObrT8eB+juQgP0aVYgMKqhVqx4lyNZJ206t/Ol
rE/h/rerNkNEBix/WvzpgH4e+mit5zRZWXnvewdfUsE5NqDkL7qVeK7QrkhSD6gy
2KSM2iWmPP+dabOhkrLnB8oNH/r519XSpvOSp8iUmlkU5WDXTyUFjNnNAXrwcTff
u7LBacZwRRiaDdxgqlndM+t1Ftlhirv6oO7WgVks8oJTswQ5GAHoeLsluPjC9OIZ
B254sN9vihiqcbIca6GhacfZgwaMMPSPzcyPeSVcsNa2GkPrg9iCuVX8P3aWvMWj
MyQTXqtDAYsvmMDAGf0LinQ9AUuQ4ZPCbzuYbVT+g6jqKDIi7MGYDL51M/TLellv
rR6WJaXH1PKR90C1XIvZPNuG9PJclHqmpE6lICk+kvXvw8sOd8GABUb6WHszGy7J
K1D1EdiyniqEtkFDlJzSI0Zg8M1ZYZnJ8UoOZqM7Jk/oliuh0UivEhqmmFg+8akc
n8XXCX6xmO4Dhne0RnD/kRlbyKvFLZWF6gs6GBaCCbpNWO2YJxpMkMP1IJ3xo+iw
DC7gOQPN4pIKJoqfK14/WkS9FQfVh8TzSIkkC1USCPHqv99pWRAjUpvnSw1H1u5l
jXKhM6YCNek8NocCdsD27M/ickG9P+nV4BpDbZjBRyBmjFb+yNvaeLBLsRVMVvEY
Y4sUkUbK5DexSAmWua0vchoo4aODLdo05AzOzUsrVfOAj183kpo8ji4s4BVAIfhK
PntTJuR//Et6xG1kWdkesamcKvdkoHswB1IwaXVBoBATtq4BgaRuLvgcWxFp8FDo
3uud3yrrihVzbEdt+/h/nkkzuSbzK1S5JKmjxFb9O04vh9d3rOX8tGaOI4t54/V7
KtuNv8TMJjcd60lu6n9uk7O/JqXcRtXUOedh9VwO+FXeUTd1Ba4AQkHe0GS30fKr
0yLv58+oeweIadCiHAH9PAMgKlqYt9P7Gm/Ah7ybe/HYG6VyZCRuw+I//ZRhYL0O
+cy+ajLm3t1+ASmWNMpU27EyxN3b1HOMgAVGqYFWzhymCfw9M19DAA3ZDtep2Rak
9zck9NcfqAGWOaXWKdAtMC7IHH2sDRRIkaqlddsIESUbwCDrhS8XlV0o98tfvWFH
BqqwcVOmC0/6MPiRkwgITMW4P1Ro3eI9/lFTEotAFkeKMK71W5TObeo8HBVTZoqY
MqN90KwVaglZ6xzBtRBCa/8bA+QwknRgujgJcWE1syBcY8pZo73MZfaFEBSAqy/6
PhkuZHq7tATv/5CFTNxUdq8AniiweE7PwdiOsxCZWFmrvEGxENP5TDAOjQ+spKUd
eisvzxkIatkCmqwAQON3oa/UEPW2z0T41LUekAsKyerDRAXEpX3hYFV87KaGpvl4
7iQ+c/AO2/Y5BQBmQPAaGImbNHJefZ6cu2eGleR/rNYFxSrkPPMSHcpv4RjzixNy
s5BRjcD7y/LmeJdjJ638s3AZBrwdO0NC92cz5BBGOY3SHsyMfXjzRvCEKZCt+gc/
oK+xN7DJSyzat8kJrQZGm5U3i6E0PJLqjiETSRS3HLIhkcX1nn6ZA9Ct9cEqCK2x
P7rYgI/XkNjcEwfUpByOZ98brbOlGqeYb1oxAat5S+0hEC+gbl+XFONFdu2Q3w+4
VLTiDMaBPypUHU2f4oK15sr8YmwL/guCljoOohN+NFm8qsZPNFEtmefx1IE1ZkoO
Z9qeCCL7h+0LtebSZz5hIF6bDdFsqgFiXabptpmy/OMW9qUdBtYOOqJW0dpLDJk+
4PpE7eyz8+0Hcj3sl2Ksu+S6omQoez8TVlG+qeucLCiVQenDyMiKESq1X8MK2Khs
b0VoC/sAN+3rmVDcSZ5JWmH2dlc0A4PaelzbjLmxCguwUEOqOVtZlkfB9KGSVw8Z
wVJtWp3bu5NBsZgamZHMv1/iyNMu8kt98dbpMzpgeH8B8zmbUCNZRrvNA3Top12C
pUClKiQILRMUq/helpqArM5mr+prKVLa0QYCOOlftWk066zN8bmPiEVw9Zn/hUVf
+esxpcT3YpVsQTyHzq1MRH/L8B/ncJMd9FS+au6bguadnvtuGdpVCGmd7c0jETI1
6MGE9axlpx9ZWSUfYfZYnHBKadbCZAwNIh8zkgHawVUiIem/hO1zlkRIb+hJMrBn
EEOE1btrVObgHkUddopNy3/s776O+BaSI1DKrb9HQgsjxP7KxNVmvhPnmhtOfwR5
zHXxPwPb0XQW4PfG2TJbhubRgOvdAxIIyIwy83NddKM2zkIdofs4wXfJlCI73rnb
SgG7VWBgsHVWAFa78MATpTV/QuPiwtcvXIec9vTz60rA6ku//Oy5kFW7Rln2zL87
UehuN+vUNuYPJhGQB6G8pcTAQukmhf8fPvjjE8QmrMUuPhQxWfhwBxI2MnqO48MO
Suoxwm0PydAMs3Xl8xC2C3fzo+bjUp7EyQgzkAtY9JHP4u9TOcAMaYvr8p7CI0pk
Cr4TzcTurkzQ6C2w0oEaIM2ZnnC4nl/lA0ic91Op/o9j/PLyn+X0RN5BZleYCEo3
W6a0LoGxIh3V/agDgkxZHk8c52+PgYw/iSP3Ygw9zkAHTdSGauoHBXny4PYbJIGg
jjy6WUS5h95fA7tng5R/sdxI4dkk1F8DcWSsVCiSUVWqOVTdYVkpN3bB36AaafDx
9+7u3f9na0EE1v8CghOyJeWBDlXEPcqWsmospmxkDD6orL6Y4X28ivRKR7urtLwR
oImKZMKIZFHCfzgjs8kdgTq/+TEwJyjij1iMJGvz9eZZq24a856IHwRiSCLY5FO3
ouXXcxgbO5569+FZC/FBThdqNLhJGSgc4jE8qgPsbgQpWHAxYLlgCYYPVnOoWlRb
PHtVTUzeOAZdhDoFPxrJmyIKZUk59F+us4Mqz/qYalpmeFpvgyzs68D7NMs0O44F
Oyr4xIrSs3/ZXXIfGs3OiB72Ojis6qVIbcj+RwnUDaqeWwtpjfBjLkabNHRvubCV
5oDqtKk0z0IPWdZ39NaURwusOaVU6IkX50veI63CYVqIRTFcBXaw+lxvZlVFn8cH
K0G7oO5s6ZoResyOFqjanTcZVzhxlOateBXmobQL66tWKelaLsvMskc3iWQsXlPN
pN1Tie0of+kETsyqJFFFtPOE49cAR09YmXVHduemWsP8Tl8BP3BerjsmnON62HBu
W5hQPOS+rJMcz3dGqZZut8D3cZ40JRnBiXgfZwHFrYF2VqtVeLv5xCel8TjSIS++
iJjx+ygCFe5+VksAy4k9b3M6llI0sgK8nrJkmin7jNJmUR8aMM9u930vCCoggdMA
mxpOtyKTknp4kyVveJ1iqrj8jwGN+wB/SbesMoJkY1EO41HivorPd7XDtASpCZwU
USs5uWh5RR1xN+JDOZXx+MR1L3YYQrJgc+aWGOCRAvfhyCt2Ng3mn7Ie2Nt3PstL
TpPQMVUn7igQaqeH4akRz9W958oBUx6HLH5jGHT7qn7PiLPBmcgUJMNoL7Cl1plp
70RDCWDyS3WTklX3ZGZOdSFNPWLY9z4lsP3OpfiMayV0Q2+t8TGgaYsdK9NZe/6R
tabhGKOFeKO8Al3GFyKJEy79zmTcA4nVT7IheEbjldiuWsYQc9BR7oRmseurf4SA
ZC0+qSo7xOci8bPN1ymg5tjSoh574r6DqctIs55pHrYNUsLAM3Z0QDl/PH3iA6as
F9yqctuEWDV9D9R/mHla0ReemQjkBJXfKByUgB1ShGK04rl6+Ovx2scqVHGOFctj
vJ6est/6d6oAicy+GFONLBJWEQaPQnTttdA300p9zEuy+yN4XgMXcFAnBI10doKV
FGdXrdgXKn1YejggC5I1f904nWwyLOok5SEdN00xdEbCcl8WqRi0KSTMoGEuutR3
BHvxdK8donfZ4S872Iw2zLwn4lWMPjM0+0O6a1q98phLMZ8flOqAdNZgyaJ5KsAn
+3+vpu5RO24v25kJJ9eVZluPmQicg4yq+pbvGpuMZhLlWiR6QfPfCRDlVEYm6ha7
b6aKCQnzHDWQefGFJIycaCnRgEb86maDAAqQJDIjfJ2qjyobpvCPHJBduV/HOvSe
7YDd/12tVhpjVAY8VQPJL6R7GMVE0Z/TKnq8hTATbA6CuiNx35clc3BG/f2hZEVU
iCXclZ0kMVLlvu4Nh3Dq8ilGTBsi17SlnGKVuZByKk09gFo4hnJlfl48ud+vm19j
3KgwqYobf2dRwoikkW0ustIkSIU8G/NAxEzm0MLcF9/iLydd3oIXc/lDjwh80KDF
Jy1Toh4dbWs3P2aSvet4I8CHvYX3d6rWpeza5P1YQ5Ua416nVcILpgKSr3EV3y0W
rTs1jj/KR86R15tg5e1SnHWZFgV23Lj6vF5MD9BM9j5WGTZBhuYIemeO7n/51eBg
+gCPfQzy+6CCDmZ5Ql0n0Npv8WXCkLvYBvyTQViqvY3LZzrC+SpfIE58CzhuytPI
b/bKQo05S010AliLY4bNQNUG0jr6jNKJys1Qk3GfHAxwsAl11Fs2pjQU8ZBaLyKc
jKSfK9dV3OGkTJ5Fwxim0b4DfmGomqQxol27FIew9rBe+ArpPXm9N5HjI+nFrMX/
JTdRf+ws3XSMYB9wbHSvxHPAHteBFAdgmBTYew/HPCBrA2xbA47QnetRE7rUhw8H
LZiB94w+siIyaORBdqD9xam/VrnOL+4Unh/L5i0uqUECAcgHql/a+g7iESwlxDKz
Q7BHdxWwKqhP6GkgWQQVZCACExu6tZH/VWbhU/BUKesOwf2/XxazYrBWLA4Fewym
QB7k55W9oAirN0LSni9FKVV3iTpwPe4/Vho5ODqklRyaLd+PsVEa23FbgmsFJmWs
0Xwi+ypFX49uzevKQI9P+MSQ1yWrBXK6kug2vVo3DYkeYaULAXPbO9hS1D6UKqx6
ZCB2Ixlam3yURSUHCpqj+c6lZ4AEeqtYJjgWBBiU8kfmKyqTI+K+ecgJqyOh0oLW
v9CNKhFwMyZ0JVXpQqACD8V7qFIy0UBro4AI01RZAtblW29cdleoTpObajgYDyCN
mVguamLa8w8uKB9UtrgViNhva/tOiJCPrSQUZ2E3fYditYc4t7B9WTfST60lFSMd
fPoZSarSKGSffg46/uCJxzABQ/OoXKYVwQOgeZ8p9X6mGLuHSGtaLKSrEjMfvcs3
huYcuSrEkZeXVt47rrX82prKzXq5rPkJrfM3c3j1sMxooCUv7fOGM/UAOSHMY0oX
vfF6sHlKwWzgFMkm7rUONa4A6kGcpVIWzu39odj164Shj6bzlPfLD3Bk9v6bSK5t
T6bfC1N1B4oIY2nx50qbc5GEWdzK95m9GpTETHaZfUT9RC9HS3SeNQH/peki/Zla
IdKAJcfrE+LoXpGaC30/GDy/2b1EHzR4nspYQ+zTKtc6bn5gKzZaitccz0PrQP8j
p0OQrDldJD999JLZns48Qsak+FWDO3Mvqy20OOXE7BAzWDpiyupNjTFpS7WUDXsH
/26niHFg6v0rQTlG/oB0pyrj04+Hgz6XtY//eCwXVu7In/ppTEXa0DD7iK7V3/F/
m8o8K5PMO9BXSg98UL8fjVAxUmEKwwE7ngqviZNmxDIRY9o5pfTk3dBe9yTCrhzr
o/MQETInJG7q30lqh8NTzh+GNe4TPP2tXtZwPtyq/xjVn0bmUctp9sr8iDtNyA+p
Khq+aDN37yZjvxjQAc67H1WbZ7sKU7sG6GtVuS83x+2/NMbEpzdau5SXV2P7LfJQ
FQwdNHhECGkn1oHR+zP0An3VDwTB9L+qtsX11gCJSfTlq1XNN0DZGcIY0rn39Be/
uVnaAGUOyrJ+xz0PCssRcLMRX9juranh6qnrqFslcAw2KmDyTEXwP91By+lRlFFF
qcfXVt1urT0+poriS55hNC1t/2BkPdHWRs/pzUVu967iY9uvfMKSdaRkMsTiHKIH
VKNTtSIcsKZbYLWosGHPLLUaF3uuyxb/tBxVAzAOLHy7iBcKO0sOn9+1DNzMYFSR
0Yr1wOqjRNYTYcKopykfrtxqMkqesZceg/4nPeykdGPlzui0h9fOeZWdXHjOAKf3
QlbOvJS3QfITRnq/CNTPwD/t0ir920j/ix7gTnhOnh4jn9wAMDSMIXlLBgyZtWaW
jggfQbmCvtBzyzx1/BDdgD5wW9YOsK71+/uX4gs7UE4qN4R95u0v6GMBDCm+JB+6
vAkf3rTpBpMb4xfShZATsuTio/gUdu4eDXGtRxuLzcaywBj5zMRNw6uo6WwSRmRE
aDLSA1OCRdW9P1U+9AcvwkZLMqXF/kMUIQhnflIpuHyB7LofDFnb1w1N1w1xxMdY
nrHC1lPhJeM7LjQ/3lXDRk/a5SGPhVQ5QMwHp/Q+M+DAYMPY7GD89fLy54kPB4IV
hyyFID4XWILeJSoZQsu4s8Um3xW9di0SzYkObg0QJG8KA/f+OU2kv7lYQ0JTVInx
ZGvxOdCj0GIebAcQ+6Ph6hrXoJlMF/nUeIDCZ1ELaEb/mKOke2knsmS0qHIjvoMM
iYUpLr2iiqIewGY/xaMs5Klf/NzNg8wMXYgSk/bGYPbLC4vjlKH8cHodSuvF0I2a
3GzDy0QzlhbEp84K34BziWLzf5KeF1j/7R1Sys7YuWpWzO7uBg5qPOG6O1loC9IM
hoWYyUNj+MHY54rHBuFECEfEmkkE46kKTV265gWI2wPsJgIBibWzvokza2lT7xUN
4+TeDsNqXZuuPEWhnAiLv0LYsVcxRkzizusuylW/be04p6MnPvnyTYGOKosiA6pt
p7pd3rcCWtBQMobLB5hraO9I/IP14/WXS9NV9BbY/xYVl0vh3K16Nmlksg7k2jmn
IRAB1qQ2f/7gLF/b1uSw1QRyYdOgfevl7SwxSQUaaX2ufR31JoXZVsq9yFGTDXAq
ea19I1QO0ZeB6DCBOsEfqfKZaZOzU3VuWk3qIVPr7R53hUJFie+G6K4u8ZzRXjl7
JCNaPfJSV+tksJiQX8UOuN6drUYJBQxIjPBNnAQEoFY/ZHhda89zGu42uUuujv1f
g+An9ERZ7apznm9zS/oA778/sFUn5Mw/r3xU+cRd4iFXa8EbXSkvYNIBJ4+QZ1Nh
`pragma protect end_protected
