// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
bGdqeFNdIOsrMkl+pVoKnr0MMGCzwVgz0Nttiqs+NGL/lhvnxonDg9txmczwju2Vu1sWaUqBkovl
T6vZf30M+O5eggsP17KwsQPhmUzRMh9uaFZ1rusJzlMuas9GeFPMZaIEAHj29CWpUhMovxYjgdR1
NRIHNL0t2z9eNnbbEbkZSxjsYjoAper72UoqXzq1vpCvl08eYQHIESC/RNCkt1q/bCbWVwnw0530
lGhummwH18qd0WWV83oGHPFJ34HtcvmujEdJYxYMXVPk83Nxc5kaWr93rF6UohIxY8GqHvDJiYRD
vVQWLdm4L+4bf1W6ZeufRwetIV+2iy1DEA+ukg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
VSTGdIw3uQ5zhune1AJOlHxV4ugJhcSPYzwNlrKKPYjWTP4qlG+5UhSyzz+mYPzZiDCSEgrp9QFO
xbZPY9kjsc0fZFuaKTvxiwkbF44T2SJBDg/ktPEpKcfsZ9DPL6iZF8+8JA43go1+jks5DSLFHxCd
gUC2sytYSHOy4AHUQlPAftXJPjdmv0vsz0WI3Win0aaNBG+nrzCEWvTSvP8MNnhVi0FK6Mohno+O
H8EuSiBKpJTCsz/vc1vUbkPcys8V5+7kH9jBf/sOyRx2w/UOVGTQT2t4R0rYmZnSUCH+e2ZBb2Gd
mpBwazPojADdT2JhavBdlBzBJUoim8hTXEwls5oEGl6LlIzZLb7D+NWUHOeOIaeP8heBaOwWLpdS
ywldyj3nzx8pF9W6v366nCxmWT2rL5Oqzew+kImaZbmvlS1WAgm0Rfs5n4DySD32Lt1Mr/GxdQzm
Kx7aHQ8fszikL7ztH/xhLHT8B0YK5QTIvCLW/I1df8MG2xrhvLyL8vc9ukrlt2pqh6WWjeTFVd8u
T9zOTnXdiWb/MPioqyJ4ojVHnK8ImyhUv+iwQWjuN7Xqn4Ft0fKE5fAFCvja1S/rB4wVwv/Oax6y
EF9UWI39rKwSNnTyURKQV9p/5fjS4I63XRv9hxRw0CuCqZmxvESCXQHHLSW0bRsMj/1TKlBJIBj2
wG2+36ceA2f760Zim9S6es/7BpW7n/92ww4HUzIuSFLia0L555bsqKwon0HJ/OSR2DyNETA7YzJj
X3AyApupmYDHnpF6aHDWSvtWsuXzXqZXHWnGwBfdKcCqvGQQySBLHDCuqGPLTg4xFFlJjfkW1qMh
cAiaBoPfGJ53Sgdc2LER2vkABQvojkelCieA84pvu13d8Rg9qT1OqaK0P40hE+UZ/Tihs6/gPgoT
SlhRRIJzRqQHyXFKKTrTz7+ZQjxk8Y6FurtQCQD616VPQrWhCtMZi+yxqv+MEj/OxRgP0QDhrXM3
dO35r41D2pMvBM3qQWw21AuhcOWdToyxFwoRvwCJ9zsLHDc+SdLxnjqvRhiUbIFsEVV8+eRRWmQb
TikKcpCDHfGRYA9LCUSy66wnRm6De1cjFBKiWtK3O9r698iuYdtmE0XUhAgv2yJHKJeHvmv0kRwq
r4vp/WjTmd2V1bpZgyfj/4z8eC772J09iqzaC1kqD6PwQP3+SdxzwB56CFwUQVYQwy0chIzHPkLx
7LC64ITbzEfmEelfqreqxkzCFICZSY47aEFDd3Ug88lnrGO776/KZb762xlhgAvacVZ5QoM1cGTQ
IGwX5xrK5Mw8spEpSmmUwmAE1aCoMOmc00UxcDHRNjx+5MMlckn94sa4R7UlX7VrNWKan45SOSOv
55xtEGkxcflc/Bglu8Nd0aPqsNGADPg3SiJDJAJLp/PH+/RrV9IMSFkoaNQ7/TtxSEKQvxK9Ur5Y
0vpKtsJh+8JZ6o8lxQ4WyZMvtfATsfJ2QVcOPdO/xcRkxXDNAye6qT0HrMZw+zlS4VCUcEEZ12Tz
0PoErfFW1edVzhmNvz370Z+CheRHU5POPcr+/6QIttxZgRIf0gD1iJydbL+uOnbuvYAGQX7NbdRb
W5ilU8MuACQNyN0egzbBuuZaSRwc3pT81WgvAHzmUhWdnybFxmnb9Dtl3I/Ua4pkIThQCM0YQqga
L7SPM9BUVo5TkBI3MMldCP16NcDlAzbEIPiryhaHvp7pEmoI2DJub4iIDmDypHQquhbDkz03hiNP
MZMXzYYOMtJZAv/Gjls8OiGu3/pnVVlj2aTrOAOeqVvNDpSnG9cNbL087aVC/xK8InHyJGUZKRP9
cjax8BbytBuNFnbpmz1jaLiJFy9DmrGzW56eUJGi0pr8pr+fIVXumbcTD8NHA1hqh4BHgQVwCfvM
HsbvB0nmir7zJmI60VXexAFdnQFKPSVOUSKP0aRaTd1O4ZVnsk11mX1EyFrsBZ4Is0mz+P0zKsFL
aTELdxvzPMDw0HQdSnWyKP9i7nu4BlJPlemWvUblimx6APbUO22/OMjQ4KBwkpyps5wxOo9YwKEd
nl3L3wQijPUIcURpXWCrwB+he1KyPnDN9eGI1/6RPTu/o+kFAxGG3+QNyC7w5ZlsuuJgYlnH9ROD
Hto96CjhG33dAQ23a0wiWysGYmQ7uhjUhSO2KAQ971b4VTW6GMVbnrPZ1jCwQY3lJpPn8Rxj5fY5
ul7pgeqnkP5QFyRVL6Q07Pr7K8AyYHLXN19dKksV3ep6x8KIcDhQDPXHUxf/yTVM8bMnrJ8nrnK7
Nf/ba7Kyc3B69E/xyNiJwBHlnvXPG41ZzTWBOfWDtxpz7vEgLX2sL7iEFhc3sH832EDSCGsV1JP2
1xeVOmDLS57UQQqNvZOi82u7AiLIBw6kXdIdIbjG2vBDjvzyUpahfShOAYuVcGl71TJQx6ehHVWo
LfgrwxT8g1TwHKP1sYn9mlRYErqwYvmzYnPpDzzrVQqug4hl0BywCqHvlA5Bu1Gy6e0joJDvTu6X
X78V+JNdBXS96U6eiJaukeidcLpzJnfpEOzBVUFDcqGp1S3os4rL3ecSsJKe25yHvsj46QJQgeuc
ADiHf3HDZxbv8/n1aQaaS9dX199tmO98dZIOv0ll7zdykvk77IHgEawa3NZIPc6CwMjf498aHEHb
tACxuXa2oMUb76WlLHt6qFhNSZuWOA/C13EDy1GIOQ3kHLFVBNvyvWbZ0t7XWGu9NR8R0W03+5Rb
mLd4KyPgQrYoSruCtV4cPlMxMEWRKDegQ5H1AcpaF9E3n7tbjqyXvl11/17vGVY4Wz+GfQ5KE/+k
+6wHBR2Ut+dxGfyTbUGhz95pO+J4MnUbWAr4KS41dwYPljd15VWIl3dpBxXJaOzIV3Hx7BJ09Ffh
puJ6vzHepZc1yMBpRyah3el2crQd0sm7Ijh3Ptex2tZj1sMZnCJh66lIgHUzljN9WCIlczDYZr+Q
NN1LiMNAGbrJv4BMNoFNgUnkML5Zt7sRoGkzYknQFRZho+GUnsFWwEtsYmUrV0BTnXXibTqXVSfs
TcP57H9IRSUdGfXsvk1szcRyQekJ0LHuwNLgnTr+Knr53/Fvf4sRk5yHK00VwosFPXuadmzYaZ/V
wJGfIBhjmpQE0W/zYSNkXpPsL6sdyAChGwCrEsDFI7Twq/vq2ngem+e3ErB7uffOssYlljroCLdW
OuK2zME8hKkfGxMxy15/ZJsEPloyApJ+U4rQpTStE75KF5mnTbZHNq2jDcIw5gEviTngY6lfDY5b
DFFOf/jCn+OVe4DxajAjN5IJqeyEl/l3V40HMFBkORiaIRl6aIwqDfGQ/pUw68C0ev2HJtoGoIMJ
cyEEPY29PpjhynG/J+yMk5BbnjnsgDxB4J97O32Sbq0Danu4TBvYkwpGjSM0j7bFCsx/iGur5rHr
6ediJ4sBzrIfso3ObtVFE3BFS83jB84mlJc4WO9tpR6SgpHpPRq/TfySK0OGMRjJPDFbcVL+8/68
474YwwOhTTpyhdFUyoqqtFOy6ZgWEyfR/8T1ur3eWPFaR+yjdw9G6QIGszYneeVI0u9POXbVmE50
rRox0J2IjnQf0IxmlmesXBJfvOHueMBhhGmIngfmN0yn/3WZTNQv82HX9XJ0VceDmJ78lcPNfEYK
/Q9aYPCvm8UwEn1e5UmifbsKRQ98gF9Vvq3U4tw+hHv9Dkv4uTAosEYDHW60fy4+TGZTTK1DyqFK
EJRTiX3vCjiDBGUx1vLneZBKRxTKkt967As3DrnKzrQ+OdTmI1WaABaYu6Tv90o0z/lY25peSUKJ
hib33icVBwkRjbMiWx0m+TmUmaRG9f/A+/XzU6BFwjUpXg3LjrluNKjeHWnijDqCo5HjcVn4DXaJ
A+0dz5KKgzNS2zT5Jf/a6EzVZwcTVqHx6NeCiVa8jBqxop5oOEkKctgBddZaDuc/LN0V6tABiPbW
1zrgPLPFj/5UtQUqcmcG8H79alUaMgRD55hNk5k3H9xxXnswTAE/HGT9dW9YqGKYSb+GgmTcf//n
RKy0102JswT/5kGIjFDftYjOYvCnWpgjHrPN6YvJaqH9gU0wb1k5st1nbucg4WvbG9p7mSB5oMxs
PtWKjBPNn3r9h6uMbl9IRoDGpBg+yHRX510LwCfbA0eWcCPGzDiH2Rbo1lpYboxm5LV7CIsM9bp6
1H4jEKqeuthotJVaxvTUoHATJn5H91sHdl5mDW7tAvKKvTWTehwIW0misIT9mC5/aV0MG1KvPM4+
+Rniw9AomkESxZzHTVRR/LNO6O7JY2yongeS60s1DLgQqT2jMYd9e0MFgBv6MyO55sAZlXX9tajn
VAxFKGQXsJsj4jj+fQwfoM0mZt9HkZMj0DcnWwVWO1v5B9K21dOB43/pOKZSIKOAYZXgVa6pUw1S
DU7rMFTnagFSMpgav7JLDHnbmtBKlRAAZ2zZwra+EtoGWX6XbuGJEbSXtz1mg9/kaY3yD4wl5QEd
QSVD3HknZ8DaJpmzOsxM6r7kga1rw/t1cPaty8bI80+NjjebJ+GQjBCU+/WPEpDuOXHlcYLY4hHo
WAKak0qhSkBWR69aUNC/7EVYvB1aOMZeMTq7zks09AQA8oKp9S7oaF0Tln+jakXwTRE6poU60F7r
BfzYz8dg5Nu+gnKqFLJ34qZd97mrkeDaWZMQb27ejMmQA1HMYgyQGfD70vQzVw3Uy6UFzrVZHUks
uFT1J8D5BYz/0+qMof99zasM43f3QwHa/GNftqLsk+Owy3RMyiNcGVUZ6dHuQ9xcgV1+rISm/NFx
/Ed6KYomLje0vN4FNdYU9ZA7UPpZoX+GiJnhg5swyCj5YkMn1KSiNMr10k14BNjm7/FFXjcP3JuR
sCa056RVkkrJHdy4Nyu8NReRwuZDnayvFZ8zFQKEbUtly+PUZDgYHI7cPglDtUNGp/wHyiX9dQ1l
3D4DpoFHe5SOVt9j5BNuC917gzs/6oXZow30EoorOQg5cvktYVydIM/Jf4MdXbnpXnV8zywzPZdb
gFQbDtyqCH5QPBMTwkXMxjorTN4Wf2cnfGeZg4iodAVvqQ6NJb+vRIjqUixo8mPrqkrmpIVyDpL1
aSwunc1wOCOu+21SpFPqpBC4rC0SmO/+vJ/XPTz/+WmATD0umH+MbsTCSCoRSdMGHM+S15TDKRNf
Rbha3d0dVoMRy24MeOGi0mA1tXoJXTqtPM7hquECEyQi7grkxEbHAso4s/+tDLji4NMMEJlOYyst
o7nOuB0CopRsOQpDlZLEe7zEQT8ErTmA4KjDvi6POtj4AaHCTT7ZhtmYZ5wZP1nJx5rr8KWF8n8R
tTukiEFtVrX5aUGnf36zWzrFoO+sNrUlYb+tLa4AHOU6262el9vY3fctNAzdq7Tr9iecVNECuzA5
z7p5ScF46wwiTwJoYPFWdF7Xse2VYVSAh0Y5VqhPwkoFtAGu8bJC62vT1csprCgE0urz+A4cc+Pn
Qwh2LkMcecP/EA63rK1jhAsn0migotCFoDLoAn/56RP4xC1lTo8LFUvoMoRS2EQ9/niGVsT+Pda4
r0vbkPMiMmF+Xk0xU8LjQ/tF6Rr+lWIH23OSOqXKgTb7EyOPbeI/bRvN2qJJ5//7vtxK5qoxAS+M
H6ilU8Kae+TUUVZELT9PVw5zgQoPJKDi/sWNo6EON9a+6KHD5WQAgnnJc7ySuosQm5YUVTJiS1mp
yLgz/aTuygBw+alQB9480FWvhaoo/roL6FPxqA6lxOD7zVDsgcp2jcjskB1iEwtjk5pvMtc0fOWp
LFmVsLLvVEZaKngS/xsRxQX68Hcu+lC0nZ1nVs6BEphICpVSd/cp2DxpT4qPZ5UwRddu5LeCyqQt
MPI1c9czBlCK0EGESAB7teqYYC/rrkX0/bZiUdjdiZP5lwSCs/2yYSme19AGHNcgpzuSA2qndTOB
4gUewEKAWM0yPTu6L28ik4B/b1Hoj2AaYqVty+4mM63SNngQQFKEEAmy3EIj3SZrONxXBBVWIQSt
j/gIkkJaFS+vv4DeP0DpJT66N5uv+OqIkGeR/gmnbnCz1m0/aff8arG8kZQIGJXbwlgaWMUUMghu
SEWjvbSrHHNbYKD1Tkog/eoOqrEG70XTH0Np1CO0PuZyvxZhIuCdF4Gnk7WshAls7DaaQj7sZUbC
aPY8I0f+uAD0bRs2OOQHrTHsvWdJDrkB2vqGcFFiii9QwXCn2BrUpyIT9zizMu5nxO2aRKR5emFe
iJLOOB8ozxdVfh2gdn0BhJYdg5IrxgoDFGeX83m7ASD4f4MZgzD/tHKrLd3Es44BKMKxpHyLHGuC
lM7hTiO8oDIkgIY37eKKdmjAcMTN9kVgvc1MpzHASFsbPe3OsvUMyWY/jCG2sZ4ooaNPxAplZMVu
oy0eOMi+Ntr77oXKlgSeg3XA2v1uKinhMMYBML8/cz2TF/IIZ372PrKiKkNbmoWNh0vcy1d7ozXh
xsWXz/Oa6mOIy3RGK/6VTbWtq+h1Fl1zrtD63pM8h/raITxdJ4WVrrPusBUnhqZHIAHvUa9nKUiE
eYwwA4a3QOgiUm+V/joK/ghs1GNiHU6Ubqxhr1ReNaqwPvl8229iVkuxgjn28z/vb6HqU2qUtCHI
jPPKNTaCHFRo1FzW1yo0MnDa94lx2PhpGoDKDeOxk5zLqCJpwoQLVBHCIQKj3T8aDksdrtRdD+0/
dD9vY0mj3bo5LAYRHqC7Gee5YycjD8AFg00X6ZRqegAZLjAn2NyOMhtU9xeprigVWf6Hro3M1srJ
a0hdEs4VeVuGPV7rIWGrkvIGc7i2rwOfeSm+7V/G7SBowdPrLArd9/WLkKfENleaqPNJmneaMNMe
/XUEf8Ld/JwBoIyPLL840YA1pfKt3ypbwq4SIJUPSFAi/Hmox3KXVxGETtQSzoCFvMYVxIzZXQiW
eHMjM9N4AR8+9J7SRjB+acECPfMy+QVIAMPuwCdW+ofpC2JbyDwGUkkIPf06FJCit8Hxz2HUf/qf
FVek5pOD/tEAHaorkzTHTXgVL4EXHdwGcgAxDvzhEaSHxrdFVIfB3R2elXfL4aaVUHzeBTLIZjTq
Tr3g6XcQWdujnm8X+yYZFGaY53kEw6+KKdqQWeFuMjdwcjXPtLcQmL0ueT030iGlNJf218hKdIPn
ZazIDh2fAaO8Gmt9TGC/9OlxQ8fQD3duTh7FnAEEXcLhJW+OPMKY3jvF34Ie1Vmr6VGO4zvD2Rga
MVgBfebGORzTmU7jKEWA+CZ/BuWDNPlj6NcBHlo3NsR3/xupm+trgStKv/UTfh5I/FFkrPnrjaTS
aSZfg/kQedeqGVDKPjbUQpV37hAQ48ZQL9E1MqIZBVisvTQzeCxqPG+xZXRbwmqsrbPIB3WaU8+j
QJppF3/uEY3oOV8cUHh7DjlmCSak4RaggX5xKZE+lb4tD3X/o1pFDHNt6skeUssOZ1ru2kzcSRS8
SnOmG6vk8+OwmqKOkW/W24AwEnP+CKyvdS3JU6byTt40cDTQ5IRSZvkHeutJ2jSnqXm+GXZLEUlj
elGgGa48g+EMDyQCpVC4RLpN+18ccDdCMLhbT4NBJPPagG3o9Ze/iwvdQDJXoUriwCJCBK56FXyE
4KW5IfOfyJ/1dSusiiaOWdrNzddi+PbC0/lZYgbuzbCkdDSbgu5pPSlu4TMOda+fKgc339Sw6Uk+
lyEez8p+PcoLBy039zw6VoNo9a3JTEgtieIJwwyly3a4shgBW7bnNGeehlYVwCtR/rjwfzDrkqB+
YjKyw9IyaZC1/wkuIHN9GjvpFPQljr5Twm8EGv1Uxfhp6jN9Sbu0ZCLS/hJFJHsVJHop/7APS//w
4pVxP6yjf9HugHTvzM7XzqDk9LFMTJiUBaEvz6JkZnpv8fMstG2jDWz7elHqijffW+C4bu/wE8cR
t/RbpOoas6A/1EGgdqMyr/OfoLcU0QicmnF5UJbbSMvgMrkgQhab1CkHbpjhsvNGFWLYDm7KU3uB
B6PI/Zfs2hRtFNECD5JThEbYxMpZ7kcroow32kDKl8gdoT1D+OyWbBRzBZDRMoFrJvweQk65ft2U
75IppyIMsYpQ0GaiJcf1DGVnGPTNu4RXzNb3vtzmszheq9pz9vMvlcxBGd7zzxdj1d/sC7yKIZee
CLZGSnkre5W0ikNAWUgdoVOfnnFANDFXJlsgfAIvNu7A987n4vgaSPWQqnCiTkGpJGPBcqZeesRf
MRTGzuBr5Jlc4Zxk/c8zgGkTz4dJry6mA93U8DnocQrs5KM5gjMKXTdGjHerZAKvGsHMHQlyqFTS
NNRbW8/JuVM47Dcu5jxYaid0WT0vgYOih/H0xKNKNUln7qig+KSItRRGrOVsVLQHDOEZ7P1VnLrg
jCSPycceBXfSCbUkdTxY0bTfV88yn7+SkObNFSWTS55V7zfGwW7SUi5kWRUR8dBIzxshfE49Oe3w
JADet8XhJchpURfLB/nXYq73d/A7sSw5nmkwQt3w/v+vn6//qT3YPwoBQxbf/y0bZ2ABxYzzj6cI
LuC7Ee3sCIRLqzW7ikzr2DPoSYvCQnoPAC0t6i4u4XblQqlOqinqaOPfFsju8Nub30Qa0oGTkaIS
tC1JIctO7G9bs04EF4XN7gq2MtTZMW7CWMZ/3XiKCdTVqtjkx3/91ouP2g2VNtijJh0sTeipoxk1
5R7CyoDebC8oqRlEMPxbvJru4VHpcSUqwz4eHOmSKM6qtIANSIyyF6gXtb2OShIccUQynSHFF5DS
weuLfrb1ldpVL3n7gDHG1M1sX2XshN8tgf9p50v4oKqIDsO5rXtEWCxxEcHwI8Op/qhBb4MRRx/R
I+qCqjgGeSZfJlvUQLBn0SCfjQ26X5k7/o8+K3zURYwA+RHE9XFLIhGOgMsXeK6tFdoJw5FvJKCe
VP9RX3BR4/cEIjc5mpoLbvJgGKEgqSqPEO9+3/UJ1FmHL9dhgxXprHyuh2IRqGo/163HQH2TapHr
OtyE78baaMql11iVp0nNhx1ASHMCwVuuM908mFcB1GJG1IlrI5OXmyubMjPun+VL8QKbW/HhxIXl
P+hgeajkdYZ9hdFq2MvWpFFEbb859/f2RQqSI7+3BLryzUvKD4Jtecmr4xVUmQuLaF+ld1twuehZ
ySi2NFqSq05ZGA6XGCWhi/KmF6GxNnFDgJKFvPwMlOrIorRnKGz8ffyoFzgyjD0BMzn3Ihz0t8cN
9vTPN8nvI52g1XLr5KZetZ4UmHnakfaKiOZH8gtJJc6fDldJ95CKlYFXePJ8MBXMURxFSWTFf1lH
8UrV6LNCuj8vdrZjcMLolkWsorzoBKwk8vBt841SmNbkijnbb+OG86WJfZjmC4KDRve+4KPRyBUO
WnlhRz+HxHhYVsxdkNx2zM1DypL3AsBa/4xFfHw4lFZcN4xSbIAGxsGATNvmf7eYAFI7H68jFVLA
C3/NSyiWZgWpFKoz05SrY9aXDt8b0UCGOSIOu/3/EPQb7qWywxQYW7Yd5dcg8mKCfynj2rF0l1MQ
sXcNFE80lmJV+nXysCL92ke9zAAAzBwpBYFIJbVM/e0gne2ziOpsq54wn0+G6bi2RgzybgAL0ix2
gXlrowgqwhzmYksDJfXWSrJcxFiKiPaIpH41chdtMJ+6KexS9B/TJ1iNQ9NJAqYuhPuIo6hdTC4P
05roBZD1spNevaboOJ4JDdvQVVCTEs5wmCludUe9clGlyjVUyAkyWzLxgY9ZuJcfwQASlziBUon5
G9DWcqV+n+F18vlg7a34irNcNk7MeKzZ1pVpJ+yfQSUH1KeJrybDw1Mv6UEgqPNNbyMDHYUtCq30
+ERkPgAdyTeu/CrYoQQaNg3edwS6p/bbHXtfaqmCLt+ysHPxHqgWrvd1rOFaXMPXtiJqXdrtCrAX
sYkhyU/v1tUsEaem7bhfbxHbfiMTaiWPTNnZelwjwhy+arelILHZZRB6gEfzpytlt+kWSvJIiLl9
pj+fqbMQXo69D1bkneB114QoXWquVXOGG14NtdrdjMFqiEsPzp9k+xGOn23uYw4+8vfN2OqtbF7Q
2X5PkbRRO+naOQyM/KOM84/AbnwVcYgeIZOvngfj372TEtIR678Wos1pQs/qYAVT8x+x/g3WM9H6
K64m8KweUFywfmR35l50kSvU8wp99NR3gmqJVUuVp0IG5dlR4pQdmxxxOK89NaomXxkxv79HOfmP
hya22jAAwmWJBZePOZg9pfJGMV/N1xQZMbMALaIYazr6KLnjkg9CMKJvvicVUclAwSMBPIJ6ylLi
Vcr74o6X1ZZDZYnm+2JjWOoUN4ur0aNgBU+/hKIq6ADy+FhW7PMSFEo8QLKfm4XGChBzPVwLCULE
ErI6d4zRQtftBqpW37LCdRCafOMG63lD8Umv/bfEnEUMMWgiR2wufViW7meCdr37UA8rQcgiK8y9
fiDoCA1UIC/PfxB6dF0wOY6hCko05x5CH65e6L26VqO6OqBHrwobqNPApA+KVrGBhdBPHadAA/JK
8mALhlCWyBRzj4fK/hm04BIKc/T2wzbogZmS9uUxtLQtuow5LtnuZMhRJdNBt7gTEmTfd8xNfA/T
clOmquFhoCfAGGNMo8rZNeiK748s6UQ61Ogb3UgT2sIdUqZrklX+oHlNxqFut2knpbTZaMOuPGu4
uJgWRSM/QobOqkbtw5pb5tAyq1GTtbnE3lXky3YsbQYOg03j5iIVF0/OrWkXJwHI4Gokq8+y02z5
mwe3xKzo6X7xP9RAyG+nZvJvqrQpT2mJhk9LMtHJLavi58HlMuYWFYQdJEwCFTikQT+/1E4rPXaN
zOD4HrMVy3kTRQ2XUaPxRzxgLtlhlQk+YvhX1gJ+FIBKzV8PyOQMx4IuoKWc6J08Y27VrPDpz/y1
BkUzPf0FwEohOCdA3StgeOTPqqogj5WxA6xuO1VitUsCvARRVlbrc2+zpbsD8wjUz7UIFLufkxT+
WxlZnUnh7YwyhC+ryxEg5kPCezHD8ly9ZKKAKyn2om45j6flanFNHsJaKlb9boqAI3hdVNQUeLpo
vugfdVHRM5h8Umr8Mzz6ebvBPcBhkGcvejpc48xjllfzJqI3jcC5X7jJYbH/pqDuO074sBrzAJnx
h6c4L6VGZe1SeASU7F12fJWi3NU4u+1/ntuI4L8hMbR7q3hxiazPTK0wJ+7nSAJ9qMaVlVApfV3L
+F9KKwVEz9GcAMGoU3Rdb2FUXvzQJ9YAtuOA1MFQTfxC8u0wEQLFoHmhET528hR104VnLUcgQx+F
PT132oaLIYCBGgX6OM4LN8V5RBQzdQIhOkqWnMCMyUvvJf3ZVJ9b8cusyHnsHYDgjXBVjBG2BqFQ
k140TDW8ZsWitV++HNOiwAD2I/sYBJ+XS2cnUS2oOw998E7UNy3bFyV4HwWtVY3krndKsEgb3Ytd
7TUOwPq2j32bNo4VwIAaMQ/IIJSasRHdhAs03+ufbilXhSfrDAh/MI0OTu5qVGba5X9evgj6ubKL
yBcj9S+ZZe0BWnPlXIoNZXUAlR1+ZtUr3iSM09K33Pzbr5sntU1O6gyE8+GI1lmxrqTm5w+AyuXZ
3slRXJSj3qT/yo/lvMskg0LPFxFpH2jQmePRsVQDrAuAxXt4F/Hhy0UurrhQlklVn5j7+VfUxmx2
6YSLkjOSq8gyP2o3jRRtyQiKpm4cV8JQp6ucjVhgngYyWFOvzMrQQa77APONKEYuGG6l4jm2Ki4w
P7VzXTQ+HKl/eIpraVTEw92tCwpVib/6naKr6XNuzbsZGP/orzZwsUQOrYHePBAQ5kmUUDBDFDUD
DHK7iaJHC0Vo+BctB/aR/+TEMjt5DepqEqOR0M64a5s+0Slaflc1ir8SgvFFlNNEWcyBYPp6/SQx
R7cU4VQpDWouh7L7rZ3Ly4je3BZYuyfACnIJG9KIqL3jyj/1bIeZHG+Ssm27JeR8j/mIlnMCheYI
nUDWhIeZdcvkHd7NnbMvAT1flGNUTJbAfnKCAoLJ5SZt+KLSeYRFKMa1W3Ll0UjEnl7INH8FJ/Dm
0WEM3YmnG1OI+qf+PKa/GTyvN1FSQ0cTo0Z2oqQ7qRjDWKvUAaF6VdtY1BJY7ElFMmUCtL4mMlpa
/5Gh4iXN7GBve3bBZIaM0qxh3n/i4abl7W6MBbwf5SF3cctfn7PKyzGna2jTBEPkTddeqdIFoUje
9cOEL84bFxxkusBAjFmi/x3s6xitpFoCUyE5okiFwY++QdprSCHwQW5Demi6efUZrTV+8KZSCC29
fBLRh6THgPNpTKzx6yOkw0NV9/fPnt8eW3BHotRq410BN0K5LN2m+lsyoAQ1Nlg33Or4MLljKlBI
g4RwEGNLrimxSm51HP/BfKZTN4TXclKOWZB6fwnHDvpElG+BKRgKypAOKT68getFamFUNnGFWNW8
/f1bsq4r64ZXNjFN7Xfb18SS47QHYHyD8gxNMHVpi1ZBVwKwmT8q6I9W0kt1pPkeeEVXyUar/JJw
dZbSI53alAZmJ4HNyEWEX+SketP3FFaOXR3Ly8fmyL2CDy5yoKzYbzc04FD9JXJyZFMszP+7cruo
HkPEmdrLHrYwdMGjFUr9EVGGtovZXzayt1TIyuexqcogAO6l1Fh+K8Z1nL66LTvF18WM9hSJyrGl
/+4wNyEFnZI8R8sp7WN6X5VMe5jAaOZqNtNcrw6xpdRgYZhxjFdVdId9f4WbJQOV7A191S+yCnKQ
D2ygCL1eb1ui7LqFRDmqUdx3aeKIu/jPy/qgoCi8ici/YKHRksmdItCRftD1AlLL7D8wFiPHLXqN
hzIUVvqGozbXh8fjkRcZbAzczMEfidDdRsEoEX0Tj7+XxQWIGpRTaZD/wWWgTITt2I1IU/ho2TKp
Mk6cxryAeOBNKpAYXJC0gk5BBTHfXvCveMVN5vkXFNzWhPdhCAlbTVKNqFHHMe51XjCKhz7lT248
uuNxpcpbqzPvnTGV0uME4MN67R6jpMl39I5kFa9Sn5GXRRKPR2FmHrdqijy0jL+FA37/Gupj9V/q
2II4JJvNzKr0fSTadHmIam0y1FXEqaIm78eM2v0/BbBoiVbimBW0EH9cs7ejzHg443a95yVp11i4
0520AegDw4PjwNlwXHmoEzjEuRjLxxperEoXwum0+UtI2owYiZooHyWxbmrmZQSwHBbSbRq1QjPh
SwG+837nqJ8cQZw5W9qVpm2IAJFJ3teuwcodzXXE1UIlfU8mNhUf1uiYnpLOwVFRGLZQ4T0hfmM8
kISTjJtpyVY3Mp8UtNsg1w+HFkEdMmrn4C0ioFWMj4zdt2H7Z3FkIpOUjhjadLg0UgUFCyLEdey/
uAIaAPs79FQzUoU8nV1H8skAHIIQr5/DE7NrGRByaEcGMDTmRQqK9uEf8+TublkleJvSDVJmhYHA
OKCp6iMBUdzfb1Q3ZjGWKDIpNppV0h2dmoCNWsRk1dkVhWJK+2ZSBcIsxH+Bi1nMHiqlMyMCuL0z
p3E+ykgmPBT7PM+IYVRYJQycXAmdcytaaMahfeayKnR6V/rfw+jIVdcl7bmypkrAE2tU9OD9uEZp
xC6D/G3n1RxidDA8HcaHUpyo/Lxck6fl4oZGx0tMFU5vxD31duF+Zniof4bWikJlYiioszWU+CFT
X85OGkHsYzNlg1//9xdlwzlpsN1WOadK2EZs0c1vH+Fz3RiNV93biCW/TSoQYa/6fZc5yXxUEIiR
TOBw+tgxlkgTThX/nXHMiA69LhXEEGVOmRPeBYNR/A/ap6Vf4wirfPFSUm0G2ZDrCsN8wPURm9/m
W2xlBag4R/59m1drjmQ/TARyS5b6SmrOh9AQRcOpQW6gWmHWCFQuskZYjdDtCRT1FTDm7WjTPGrB
kB6Z4YTDQrTsD7u2X9+7/MUcFjHPSfl0EIirOVX4nO7DOdB6gpIA7rCqVaodxQgEA7QeXurYaAlc
g7/ShPrO9JcH+2ehYj8aMSMCPSY9LAzqgnP0T2TTm/ZgrBgisoKOoQRdK+mUI7HH+hQTRd8olgnN
+mO0fJCks/bWR4zc6VTmYeOIth0LbwV8BYPCTHpF1oTcr+6TD5kJOjmTTHu1Y5w+trihJIUYJ9jT
o6gHFdGRKr75hx1hsht1rGvI71awb0U8aiRABPvRttxreUJZ4D4jPZkGD+IGI4SC+I+eQUPTNaaa
W3p7OhiTJ6XDqoJxgWzcAP+Q+JvxrWvMQxS4TPADc3+8zyWAbqzDrfhhwhklIhy/geHL380wodhm
L+pGjo3wXFwhT/3KaM+b1jP9qYiZgqK9sksxHzbXLIigzMUWYGfmdH8j7NX0H3xDVXg89ZBOhWdk
IPmV1OLgRL5oErkCl5ShkqwCMY5GamQ/LO0Tee3vKtjh7fqjGL12Uz/Y9+mrCLiQ69jzlcXI2waH
b99BEXMk2yaErh0LIMq9soCm/RAVVumtCTuGw6dVBsPOuYVCoZ8CGeyYYlMONoJwOXtXPhTqbqbP
RE1r+AuYLsB0KUXIsx7cC4C6pdX8iXHBXsFlXD84NfF29pJhD76u7C5D3DS/cC7TgdeJl+THRIox
DuEQfBYSzcONZcGuzHySkhdDMBXm27qtqH7juligkPRIw2PpNMOLLfCWiJZCwH7DT8qV7O8AxSlF
4uOZCQ7ATKBkE4rr1GlsllK7pTcN2S0Dh8hODn3dA2mowMsyysm0LjQ9/gFMAVZ6brGIjki2ycSN
XV7uNoak35NyExafnMcNkxWWzlSZ9N1B2AhW8IBkGZhlALjiFEmM1vb5GXX7bH54BcfcxzzDD073
hOzfPM6TJaOaUc7/ALNVjPZmBeUqK2F9JtaCaARTlk4tG2sTkrIqTiqBvsjaP0YghGNKbfG75E+U
nHL+g5FRMvWwqldhGdMA5GOmH1TKYW7mdNbG2OdN1A1WZweHT+WZID9YFCdson01TR2rz6nef4jX
8cowOXSgXsh5+EgxBOofLBCwtECeeBg4qJVIhQFJEYrUTw6ZWbMyHX2zGHOvk+gJYTRBz6cu3NlA
sVa7A+3s9DbTWlPY03jG9GtEF+ETFJ/gEpceupWyucb8mClC61O1YYY83T1pqunupFOePuGr3wou
CSFu+mlaYrvJkAe/txPvwTmhQTlC4Ju0ZQ3xnmNCWFC6u4a556IcczsBwb7MD4KMvk9ijRhgkxzb
ErrDvppia8betx/gJKw30qWSx5l0+I7x/LgY3RFf0fD+wJCAp0NFeFOXJ+99IkeWDkz3d0Is0JxU
FIcpB0LuBnaACOq2YtiGCmyvC5i//9bC29ZqcNx2IwUruHgv1PzeyHH8nbfyubXmNrrS7+vbKs8v
NtHykCSgAPfjPTZ7sBs5J1EUQRSZh0xcsbqyqxtVDjuZE0+gb0Ye2xgPrYjP/9h9HWVDvGLzp+5w
jTWQcyfWpGhqG9bjf5qAgttr7U9PJ68opdNPrAw5SPObt3joKW3WGFGRQWwp7dZ+8DgjLTg7FzZb
wMZfFK+xi+pUAgRkcgZXUovGjfxn+gr9tuU6C+PlwXAOBF9tejksrxn2qr+dBe+0BzFlqI5eaAeQ
v/S/NspFjGTgs05O6NMmH/kulH2PNpqk8E+H1WBEo6pGbe2C8+N87ZsGT3LgH5mhDRaIYe0YblSY
Vd9di5m7ES2u6ykIu/C4G20vGzvEYVzkwJ4qCh3TEfwaMMosVFLIqrRDY7ZWRMtjxGYnfvyLgyGH
8QrG9efWoq4BzwZUWiXKyMts13ButNFm+JkAUGPzNSV31hweuNK1mXPVEj18h5AdL4SERdQKzFRL
fFF2lx0pIrRTTzsi+8zVGbBHmBSOA4BZ8PEX/NSg5wG74/IPbc4l9/obMcuyYxdOijX5zFX9TNA2
fNJBVu8fxnnlEfavc8ufp0EsUwmyFnJyQtdzDjzOmnyqcaPkWKf3s1DIE0qjryL7NJcnHRN/F7cA
2GsW7IhuEhj83wqWicUwCsiK9D8mu05x7zuetBe5SA4y4OFeWRmJNeioFIeau866j+2ZuYZBA7kV
WFuyd4AcPYygr2U6kB6KnJ8tFGUCFlPArhGjFQH7PrUCkvlAzm9o6cgwblDaGdG+im5xtwuzdl1B
xFkspGYQUdKxHEFWFEjOlTEt4b02W4ARfjPOYtcU57Rm6CZAJoSForM1UyM/qrlP5E+GRXqvXj8U
pWihnu1wUaLa7BERy6GtQj57ORGzYNjXTvlmD1c0Z2I99oHnhg1qbTYm9rQNFRAjy9lM1y/uDDSY
MJghkzXEFCRHN1y8mFxLppvsGP82Wp6uJvsn0DkUiIrQFmVgU3azPc83Qw6pnMGru8Xh4Po+J48L
Os6thzJczDZRxP83oWjS5G0IoO+Ln4XuDqSocGvpldXteAgZ/nXtOp9wSPXTo8vNMwfDyEnJ+Hb7
r4dZP/95KsihLFHWid+8GN9aD3PZiaWRN0DIbXNW1+0CXJIaqJ5cNNxPTL26B2kmfEml50NmBVxa
Bju64wYaE4OucYJGP1UCxpZ3Bb/rEg7meCnufUyknlv7llcjNUvAfgmU9NBsLOypf6ixTUwxjvuU
gbRxgbU1OLcLKgwxSNeg249nwUIybC+8WOjpA64Hpfi6g9Fl3PwWOdEsnGgc2wf0bHIEBBYMjP1z
hiYGeM6qz8h1Yd/0bv+UPwCARx2UyDxPYL//Hu98vWprx2NeWSwgfT6dOgBnSBcSt/o8oONYfVki
V+bxoHIePC1AjJyj9fgFl0sHaD5YURQwAnys74qJh18uP88icntLoJ8hd91oAmPTTen1Op5S7Pka
OZS3uGv8+7sZ9oHsk2hFNJLkEFmyt+YtTjKFv95YgHlurpmR5AUaTTf+Z64ngeC0kuQTYlKRAV08
XzzTOq+qij5kv4OYzLh4lPpISsJE3gKFDjuOmr0BQwZbzQHFe+TyBhvtuDI74TQJVcGPEqphGmpy
oVEcxQXeeDtc0CxP7qMxR9cPJaWf/xxpNUDCi+TptcAnOXNYubv7hvwd5xTZ1hlXivHPknvmIiCp
bn1gqotkfod6ge3Q0ApceUShhv0CXCtgk+LlfZjDq+eFeu6Wm3IxsxA0W/QKwGzx1b7O+1bSmxt1
TvE1CaTxL2epL+PoEIq6E4ewN8mS88v+psdlHTP8CAqMHHcl5o5+muxAxtGiBeWrgwFh0jMiRQ9f
0hVkqtX/GtqadvNrsIQr+/YyJv5TI4XmhqlxVPt996D3Gwycond6K6IExDjfqlwG94DakhrRN0K7
pvkxM9fsUXLuAOeejkjvxAr7bO0cLxZbY3yVkBqKC7CjeqAZ+LRS4lvF/7vphjN+8tDDmx6tNFxE
kAECMfdqckifPjb9bsJrFagfn5gaxYtxdhpU3fiVdJ8oAbRixxHgLrOGy8TlkEHDDcTTeZPjZ7Ni
mtk7fXoEEFUxYOIm5n+YVoGo0ZCExyQ6G4GYm3jR5J4ekURgh3zb0dbOYDEz2cxx0QmEbK8Fs+gP
6Z3C0JeAeurvxgs6N3FYuFBQXPwXfvTXG/ouB80rGKzzxcg7W5QohMsDO3cYtPecltrbBNA8UyQU
zsjacj08on1Ls9GZ1L9g1aT7XOwb2KkwDOosdMk30j9VtfFevciXkOfF4MzRGkcEtDo/xetJqrdC
s7x9OO2V/ht3ogWtWrZYiMVZFaQHUmQfIwOi3ytFICOABQPISOVctkg8ZNoN8twsvhyDA2XumVj4
+iBXxIpaUF4OMW23fin0woeC6J5DLhPbpXVuF6bwgubgPD7fVTP1IaRSKIe/0CoPsLatVRe0y4KI
PxTmKDxo/ZfGMa9U+rnmA7axqd2Luf6SZSfoNcZl1dpkZPxAl+gfvl7PIR5MOEHr+CTClug9ml7E
YtkysfuMOy+fnJ9lXfzNRGBkHY23xw7iFDoONZ5HMhs+JvfYuLdOiQw4PTLjD7wD8b94zK2EmXO8
8UX7cBZwo2KyO6UOl6VPkCAenm5G2kMwGZJphasu/u6MYMcLrz8xDbwNw0UAEcs58oq/gYuwOzYx
CciZ6pcuYJ/3g6mstsRqrc3+XLKJCYYwusqZn0ZTrqoQjB3zniYsfeSuVctRNOffzhynMCouDGIV
3TbjPTQ2faecjGPLYxGtKo0I/KgfguCfkr6w15QD9+67GFO3fHHA5RjUKARF510kUkRz8A9CKQHF
02KY4MV3S1Pc/OvB28Lf87Q7I4bYU7YVTKEABqCTiDtCkQV8hxJxbIvg3Etl4E1Qa23mnurbY3C5
S25bhQ+ICLYK2sxaCS9RGTunrookwgCFyATnyxGebRjGgMFsQu4xh5k5+yiu5ix8F2jGUx3348vR
BoyQ47aazXlNcoplEK4IoyMvvyBoAoGNv7Tz4RcQ4gfqdtsWg7lyPsyH78uM4D81jvJX+JmmGb3n
mNHVk9QzTjtk9/2eRKrlx8kQFYNXtnjEjDR0lk9JjvL1kuk7KGRY2eP5dZPH8sTP7QiPAv58dlCk
86fCFbD3ukyB1zhgLbnFSidfH/C7571qIRihuWuNmHjjPPvMP+fa78E2hjLjllpTroU9L9wXQR80
CeVMg8BbHE38V8MuxkdaPKkl5FZ8n+VMVtEUkJx7wtR+IqaPHMZwARvGk9C4Y3wRyv/BsKOH4KIF
qEHCh8j3uKQwOVZgDFS0+jog9m5ONacaNG9F0UcLGojL2h5kQ6+qaqakdyOqo/QSlIm56FX2Fy1i
eIfB+4k8rwk4HDM78JSOYw2Uhskcj4oz/Uxu1+PugjYslj18QVAlEIIGq6E2OLGcQipBK08gRG1r
M1fs9omqPrKipQqN0XRHg9Wlw2+NUCl3HF51iBhZ8OerxJyfP93oRU0ewurFy3q5h/3ULb7yHjbp
A1MgYobUqXtThQdcmilHZD7lUQNwqe1O2j+6vqoU8qdUkB6rja9cIveebIYsch+WHVxiG+0FojYX
X/fW6eeZJE24btFDeFtn/8VgGnz8iuNW6Jx6mr5nlD5QIPo552wkYY/wn+a2Z2i2f/xHE9UVYirB
lMVKcWBT1tMCnXqbSnxQK69U+rNhH6tPE8EKtKfTeGeIOZE59BV2yaz60zdZCJxEFBsZlx9s6Vug
9o3OT89U2/COzbklGNOSXi4U4mbGvTUZe5ZoR1dE7uBV6l94DikRhhLQ/FGsHETiC3vdrCLTSedT
XtIub0YXj2CTrhdQ8DxK4V0wa0t0O2hBGTeDvsKBoo2l0zKTfplZn3FtwcHJNblopxrQjVJvzITo
QurqZEY+4tCXhD2p0qFl7oEeKjIqPkLXKW7c3W6TOHtTQRYMxRvA3A2AD9XOVXvQ7JNNVyND5spe
+svO5/ptGnFW25ORZex4DZTT+qdiW+hkiUZnn6keQh5yRZKztTxL/2UMD5GhcDFCLb1VZ5iH7FqR
UpQHHn0kxrr0p1a1qN3T4c7qFT1MBYoAZHjkfkYzTOiWCNxdVXck1N0J3Pm4vY7MlJjf3JP4vJsy
z7OZDH6A+z7mge9WKrSTNLy3DXbiDG6RDg7NchB8tAM++/PJopj3GHqZ0MMUX+INboc4/xTzy9yT
BjpNNussehnJWASZ/F3ebhnEDBnDQ/uuJELLKuaxmaFDtnf+1oKaObnTiOvsWwCyxywn0bgIIe9w
PKgGn7O+NNZYFyAZpxGeDZocCYJ88D4j2n+pe787YjPez/JkQHCEbvDJ4+KtBvlpGIpbaBPfJCfa
FOEwI2t7Y9LslZPLiPUA0NmZKSSsGk86IzFFAI5tP2xiTcLs9B6H4NeJkQk1JMFFeVBfvAGG01+9
Jj2FV8QdpVPPfCNaVzMg5ZKA+E7hvl9BknTAX0+WRcxuI9kp3p/0jPFbqzfRAlguYAUpzoMppgxi
8ooeeKkW/jzdcVUu7LFjM/sZem3yNYk2xJZ2OfCIwEQooOva5P4Vs1UJV2gRmrZhbvfgvWzEFG3U
n19fQemD/R3VcWFkS30De3ur1Zu0miy9dFEOxnULzfn2DZTcU8IK4VNUFDWxzr3XCBj6646lxOVD
oca91SGLFafYJV92270YRn3Pl1+xaw9STQ/6q6/vPdOvUifRTROTfURQDxnvQF3m6orkN+Fsc3kM
53EPVwVWa7ImJL0RSL0g7TUSUk2693Jkg7RW1h4COtROW3Ue9Q7XERqmDFFX2RunE4Tob9TP8tXh
lCu8+D6ZpTqmuhf3z6nFLQcyRmmP5JHh+00p3O9W9L8ZcFp+Zd4Ku6G3usvswH+ZPQzSNDZ6Mynq
+67COYimt/kn8YbPuAF0Yc9c+BKWroQtXTvhO0t0Z4plZMqMuoKPmOw+orw0x3Vu25wYqRE0k+uw
KHN0cjm+u6av9LwDpBOFj2JpNAtVqkbAmTRF/TE+RE8zDnagYY5wmHaNC3FQ/ggKyScsNaYekFCJ
JdUQ31JOHfOg5HFqLoU84dU1RD+EK1fNgTH5tFJ9RWiDHiaZhqC2dOwGCJU0M/IVc0FRdvEbPqYf
4yJKqqnKcprUmk9AF0Xv/Ln/5te6iXgvWXklvLATgSDT2PiJ9FnhNwHwVRYbv1V5wLDVQkcCE82y
+vV7HQXmh/fcIIh6R1jlahCpxfCczjX2OPCjSLbBBpfpgKJwUp/WiytMvHKCsBi3umej0c2bm5Pt
tyGSKJbVayB10LkI+LwLCW7ZzLaSL3uBTxyDyO9HD+QyPeHhpUUD3LtinZVllDKAImFyCPCUQ0+9
IQwYDpU+gl5CW4GFWmOa3qZ+4CubrzTxIkOErzh3n7Qy9SU4NTRaHwLXp1xOSlLaAESx4c8dmweQ
iwmEsE5LpWIvUY94+Vl6m7q/XoquEInG+3R4T/xEOoNAktHCEViVzEYSoB+PSK9KFLZN3ARPoQDA
3hibVHp4SzW8Du+g9X3O/ESEAvxWaQ8nz3zKqFHeq4DdfPA1RamEEu2NhHy/AaffZz/9t00sozjk
+K8byf6FcBzAfJdk4F/+LX2JQ3xYN9WOx8+GR6yDYnly4VElD3f9ptZWIOzcySYB3dOeURhGA6YA
252wULobXqQX+Khbw861/Sns/f739/FUUyChrvlWaaNPSIMpvsWr00VUOTWtz43MgJ80RFqKuvhu
an8/5tKwEyNMCUSvP/2LyjOMN/36BIBatUAQDMi58/8WvzxhtW9QInbRCNZ4ZslcUILuNOMG28/Y
YN4N/x9Zx9eA7yfvmqVqGhqTSXdBqBmdvbccQlMqXuMniBcEu/mZFvYPh07ujMUzO3SQDx6fgE8D
M7CGD8izbS44DotHbAlhVSbScXZtoUXazpgwxV+GEXVsfAN5ba2QL8tadmE5xCqHTb6/XteOIkcs
7uElk85ZXwibQWFlQBzPC7agh7CuNSTO+YlgGfMqOa6P/lOZx/6UBNKq10OjJN4hTw9wmglshXez
l4nZvxo69MD1FN6g+m51TjhjJVuNFF6VmB+e1n4jR6/J+wtvXOr66PQSozTmIRszdAcEMawe41qj
zHHjFdF6bte4yiSxbgQbMGP3yo8sF7506VrH2fC1eZtEu6/TsSVanlEXFvDgwpqeSIGWIUPJsDiT
qaj4gzAzMRFCBEFR5lljOAIkj1dXNh2+NaXZgZyM1wTVcn6xg04XHtDyERAWtx+2SKl1ootv9f9i
pVpecOGjGKzr5XqMV4/0pdsGhKQh9/fk30brAzvn5ByYwZviMxvrnv5jUCR56xRDS5HF5/9Tj8g7
0nWe8Rafo4nLQWI7I829DYPJ5SXo/O8sCWM//KAsf6ihVS2XIrTps9rv8ZwJNrlcfzx+x4KBdoeO
1wBB2rkSdwPa+rFRw4VeFxTaAJrXXjmxefP9O78vubYRYSZiIqsFTXkirl0jWhP5gge59X2tv9Eb
2jdR0rxOOFOI1NEWT1y6KM83MgoYfnUjMvzQGO+ZJZquOC9BObt64XaDr7iMndmIl10pPZeu99it
RIkB/mnMIlEV8jr31l2TrwYxp/J4CKKnWL+bjH0FsinWQC2NzvzMw3CZLdVBO5YDlzezdhEb6PcL
6AjclcTsTV5MCTd4YQ6qn8nhSsH0uRmiX1+F51I1G/lqj9ZA3ID26oigWlNUkvbcWBwm0dfk/ha4
rKl2YHYBB/AZGgZwrgwNGDurgH3AP31YModKP1r3YH965q/jqQsHg4PM51GXzqKCO4DL/GHfSuN9
6cPCkFNaYsGMzRhMrQ/a9Co0e6+VJrdb39+hgMrTk+fMr1rkvtd16M3lZy78GtnfVWZWCAJxEupq
SqridqEJhCm3BlbPixPLgwdJe2ltghSV4iVAF6vu6I7CMX1qksTSCBIo1WpbzbZKiwV+tlyJQXz+
fnVzEt7rtPLLn6bAhJXSwGnm1NPRtew5XKdCkjtGrbpHlBNOOX1erBxrNTVdJG9DV3wKj1B84wzR
d2kuefd1Xovt2pvG+AmMUsaTEBTFqmswPbFBOpjOLSK0pS9xofia/RvGU7MMhFGLKBiuEJil2TWH
QtyG2CClH1bOuKgFwQHrgtOQvn77206gVu+bsjtKsnWAeAYfY3D4gDkpmyW0KuWZwchvTFwkon/K
Frk1z49J7E2OJNr8TX9zloeyuRM4JUE/ySVPmwY2PQ63fatgu+aaAs6uTv3eYcce2byVunFjM9jA
eMD+ck65P4Z11HOLIlX0uHvr1OUowJIkbD2bfwg5Y700fiopej1S8RBpGaEnrjOj6Iao5PpppjJb
nQB4TXElORRaoAgKFC7xfl+HNtqj7N1tUAOYbqnUW7f4EcktK5yG27hKiQH3ujh0GbDSwt7zy/R/
Djz1BTJwYGckBtG9NT9pP4PBydm79od/8z+sZ6rbUYHW0C+wSA5qOy8qDGnlXOdaPN7A84lMbf/4
7c8S44zgppMQUZQqWJDMlAkpf6ZGFqPyfryC/lQk2k9FELnCTxwqO+/cXtw+1iqNhj+jsPY+PSsq
KIcvv97R9cWgeMy8gTdsTSeDhqUGsWHlfz83P17gXKCNdZraRaIPCvs706joiqT+udq9Gm59devr
tcNSXg4iLsI5Q3SDPe0rkYtKol6Cgob17iwcGFv/luNnrOcCTqg/DsbA27teuZld3HjCPKd1Rm6l
+ETOg78gIBXVaQ1O6tIumyLl5tP/XTnmCLdAkrNnpIUAdu2MSbPb4F6ME1YzmZye+XFfEvqV/f8h
LJCorY03BNvftwqwXVJS6MicToyrOIUcIorDHvoohI4dgYIQJHepX+lOqK75+2ECQTDWduEkDman
tMDGMWuyJDsdU0p9edcRhBijkXtdF3GPoCajebWH66pE6O/XTdH9PxOJVHipw7RK4aqI0qVDSbEk
UP6e7fdkUYj7q685VgUpV0fsMQkSjCkqcTBZ3d6Y9MF2cN2XlfH8uPBtzkmu/RpebEyyhmJkhPWB
2JmYYTue4DznpHuX5qkN1d94CgAiW4bsIA0tq9g8+j9j5KzApU/1OhLpj9rCCT3QWhB7ej19X//F
9igqYL6JuSSVCkEMacHdGDkBv6T6btB3OQr2Z+SaxSEhrFkYFu0Z622zQFvERehT9SyLOYlOswZ0
/JwAqggx8IQ1NS2koO1MU7e/AYr0FaWRDri2pCj3Od4Ju3Ys09/8rbfMFcJRlu/DeodEMazM+Xue
NR+Bf/jyL/VkhSp0PX9Y0FQm0IOmIq3xpSuJQAc4EiOxVMHlHLOUlInDiHhWUqMlroNxcqCS/K92
yHXRxUoRwoylXlfo0EMQFntdUtPWaW/cCFknqDydGNjOYBVOUCDn9SnClzEuD3ZxSsb138++6kkg
90AHm5zop7hPnf77WlR0G03YtlKh7QFT6qGyzPpipO2aUB8fRljxT89+7ziKq756KvulWpajIET2
xXU/WxLakeoknDds0X86AL+9VggTTfTFhTWg5PYoLsBoFsW43HNTBnzLAKOPTYqOT8DfjItZr7Hs
JASCpC+ugcHbhbQJEU1btubyrm81tBVEfA4wF3NV1oCK+TgtPxSdQzQbj0lGkRvRPapRhRcS3FHp
R2CCT9CM89kEdXgV452X1rFl2ZTb0udLb4DrzV8yxESLJQPjf9aj7BWqYL8i34n49H263H7tjt+8
t+yCZnrRFKP7Hx5t1+Mq2tpFFiV30x1mDIBJGPX4m++8ZtRJjtZc51XsBVfd56e4qnLL+t/zVgMi
oqo2WPk+GqnnyufKGUmMU/8mLLdrm8tPyP8zm+Xi647kWXqrRutkdYCqLczNJMfm7MiCisJWx7Vz
sSUj9wJujyvYTPQEcY9xN4/zCNDK+h1tjzDzJDATcbreOh99wZc+0u8dvWmXKahB4rnXlcTfC/Ji
WrB3aNbW1CtPNW8BmRU1trB1W8N12saVQ5C9JkCDyZO1RFrZoxdlX4iSUp9X4CpbHSFaRX8NWAcp
i5yF2K9buMGbzfigC8jtRjGliQ1ZE862ZrBUphWMXxdf4GWdOob85uDb+yZB0hfR5pRElkh8HDMT
L7rxZ1d5FMLUlBh6Xs1B/oG1TgVJYzLN4ZjpdqNjYfGwJqihrqVpXAxrcbUS43P8Nf0byEt9Ctfr
huoyfwlChQMSQaF+S7gR7Oego3RAzeDvgSd6fdDDYWqs9zILz8h40gUqt7HAwCAMcmPItLUx7rlI
bDTfWvMCUCPQbfnB+cWqrniRYjEdUHNPBBDs3uvUZrSNPtomdPLCxZhVKlW+8UFfOeLHKMR+w91a
ZYexY1wDqhrt+CacQJYhIZc297hXPafXso5+QDk6CRAnc+XyJTteUjo0Q4vW4lMF2Bvq+Ae/r5gz
Y1DprsPcqiGu/rKe34CHT5RERoRYke4k/MQ87C+JeQYOM4D0oI8fFHJFU+c/LUIx7m0E/CQMrWpQ
IsSAyt1JuG2f+wciYoOlK0JPNZ7Qwk9gHE3Sv6xhGTQi1kRJuLCYZiijaaUXaMSiXem93hzcjZMe
hJa3uH6xgl3A1VSOwbwXeGsIrsHHEszXnHHFPpiGeUfUQd/05SVqa9UcLrsqh1csj3/LiltmeI8C
QkL4oFISsqBRd8so/CocQnz0TemjbSTgX+aR1RlbhUelvMnpmOmf9R6fkDS8r42iYz/ysIKFAB/3
3CiYoV8O0YO7YnqR2Ovx48TtiSEraI1wMeJ+fLpDlsHC3+NWjfjeoqLsb1kzzcFf6CIVf77+M1FM
dHIgDLsEOv9kviVbZFMwspGdr+kj8DpVcuNmSRngSvPmm5Gg64M4x72A7nWlHK1qGiI/Hvd7kslX
QHq2J7j10zRZrpv/E+n87NF9z08VN6UlpEx2Ofp4R1GN9Bwa61txoVYridk2G/oZpDfEIuO7j6q4
H8Ydz+mv6tbvpDO0zyDFWOmeu/H1shU27vo+odbqxUUYisWj2PcmiFujq9l+FUks6v4tlI+M5sSr
g9e/CtuZoztaHf6AJ2j1beLMMtwdDPdAf2IDcAqrFvG9mSHwdmcOob5T7WBDSbD0dryipqOxk/ci
UzrRpAFQ11nQ7mDeI0VB+lwImu/dFgBfjSMVkJ1NFC1ZGAP6wgQDPdlkI9hwm4PNKSd0JRa3z514
vhWvbecTyf4sW0zYsgRFqMvq2oZDkhFsf4Q9kWCri8AZXKgO8URKQgjxpsqIl0/aRO7bkjCR7P2P
a756gz+pysAv65LRSxSbfL/MjmxHCKbNhIrDYUS3iAu1zm3w8DdpHpuEPgt9S9loe5SynvnV69cG
+LJ7p0IYzt8994rX+ODD2jVis9SdiA6CjLv+Gm0xJfuEJ414K33F+/ZG3fdw7/bdcvCLz35HEDlL
WFcbe9wvlLVNSEZ33dK63VkWXB6VxI0X0Fx20pEShsCWmLHdmuOf1qDuoNesuWZIQdBEoc7cWcAC
zYqC5hSgRnOA0FNSdXfY69qTYdAXrUJSmI/pbo9Hsdv1Xv/e2v9bu0Tof260eGhm+dYFCxPmrHil
Ps03hBPXnsEst638pzINV4bdBKesJNpx2j0OIBSByGg1UKELKMUCgmcUcKS5gfNvfIEnxGulV++M
wXBTKS6EZl8Z8jlxyAB8jEJN94MaP8MOta7YRf5eC0ZSTxJCm66gFOu3p89DDMCxQM7mGsplapSK
rwA1/PO31Yxe2hnfokcwA0t81LC1S5GynjgdUrddSS6JvBJ4TKqVh8PRLsEjaieUP7pylCLbOMNB
TmobSKdJyKDgUh+C0tv4P2i/uoLuEiAKUmhsnoMMKdKO5UzI3Cd6pcFlSA0iUzwbc5aSJINKRa8V
4e+JWy0vK4wR4fAJqZYr6nntOBLQquKiH2qVgRqFUdzXVfrSBq5t5Jo6rM6oxcsyHItcvypTg35L
aoIaOrW7IFnAKVQR55uBVQkpNIwpXKZqIqCACOxK6UfkUleTBywk6Pk2UMk52OJkS8jwIA1t+0as
tFE6IOTwlxH15RZn1gdxllKJMyetwK+tWXI5sWe4B4VspDXN7KtIRGjlaJsw1FsElru2A9LiP0AC
5k5HnSVBbBVe6Lz8njwkYsoJRFJMCmTlBwYcQ5K8CcAj89v+IJ1fsfmCY3EvbLy4oFIGlCAqvuV3
SXJ7MfMIEqp7OgbmQQiGaPqr4s9OVXli9EkdqnHq3XXZcb8JYXKVcE1f9RdPc8GqNof45vaymE9Y
lv+fZq84LjnEnrOh9Y106P5kFqyAwLCktltzWTjAwUgyfpa0uL8T+kDih9vCjRFg5ZVr4iREXpXl
ygen8ae/oeFmB7jjVxSaVi6AAsGeJKETYb/R+HSEJ40xgikxoE3mdqH6IbiCjIjy8Tmr2Px4mw4C
Pflx3tbe5COz6KyItUbgxQJHe6AM6QNa1xI4yPUeQrba3FsddhZr4q99UqAffGv5GkDY/bv5WrZQ
VwZBRCZCELw0slAEzw0q5AD1noTK+4xwuDaDRrpYiwW25KW8+q7cl/dsXvOLZSell7v7KiOqE449
pOzkicLKoNVUjvd9vDGA7Yn+p8Xkn9xAwJXsoqILLqpZCvCp8NeI9AFZ+UUcts3q/f/ECBzGhFj3
L6/bHCJTto4JIOcnBAGmmJRup8KNBzyWNPpLQD8WEWGcwWh/FkU16FQPJ8rr7l30X3P1/7tSc9Ks
K6Z1O2Uh3EqXuBES2IKWXOYHW2RNqfCet6JG48kZB+czBIkWiN87RbqaUWs9rF8FDZeX0per5x0f
p/j3u+qc9+u8NRgC2H6LwmkhSMlTuGdRCaBO4Z/YpRI/kKTJ8xTjcpXrzCOhf9FFztBggD0mIGZR
NBYBWS6iPiUJ/2ZokJIRnnO6s7AY7oLz8OaotD5NjpAgV2+ZIh2F3pdDH3I0d8d7XRUvc2a5ROo9
YKUD50Nhkei2Wp/i1f4j59CEfN7VsfvU/nidj8NlqXHu2afj7Nm2G2P62bBbXvl9g6IzsVBtlf/E
JRoS82t6Elh9tmJdUPPfoCoSrGWOGBWcUEOjEEft51swD5OttWKAkSgtcjL6qmc/9TVfZxrbHk5C
AVQOaEha8FvgbPt4D7h0prew7KYUnCe873eS52xQxJdsjbmzX/AO9cte3vsqlbUUeNSqLSAui2Bq
qfH3O0prtmhF3jSw4oQv+ccFRXCvDxQI2zS68g5HU11XVzHGCJsPVv4Fdjo0+a/NZQxPBQf/jwdw
azWnFMeeVO1NBATyYPfOOIna6pDUWUMqXPBEuKiB7sqDxH1oCWIFOzaCrgSvzHJVzqxL1cWszxiK
lySkLI/V0lcKp7FnYgAH7KmM4apIQV2+nw6a6HOXmxJDW+ZvnTWMLwMPPHQYGVXuIURD96w94E6A
QSY/Cnsk2eSWTzH2CZNLN5GY329ik90nsY7/cRBqzUKac5/DH9Fj/jHYqDQUClk0Oq8BWoh8V8Bb
3nRD43KVUIMz/NsDl3s2etgkyY9Y/rl4wCid7tMD0uuydTn5i3MrSkHdm/avcLJ7srU1mAxfv9fN
JLchyak0b+lxxwPfJOZk9KJVT7cUWD6c6SjXjodsrQMPi17S4aLWuF5bphQlujywe1cFjIxjJ6fA
ThdlRa8Ahp+ymVjxJfQeP5sPCU3sK/fD/5GO87AB8GcQMt8Qfd4s5bQV0skAlboB6GbQC26/2ike
2oP1S6viFChNCkY1Zg19J8FKnCZJeXcrNN/TVLMfheJ9wiXd2OSXlvhod4pFCFc56BsykEEO6EwA
qR7YwdLXE93ag8sbeRkmv8jHGnHfsvUxD+zCBcU6Jnkyb1LJ16TfnK/18/JziaJiVl8QYfDTJC4M
N1dUdQahPFf47BjtaRmw8EjxUDLsSYMLucL23dLZODNqjbVv1WtTQOBFSlgm54csN4lXEAz/MCHQ
0p/5hV6fAAs716JqpOv5NIPIKztfUkc0yXaAyBODo2aBxCg4GUK7JdMhYSwM3rd4nqtfLZyG1dwz
TPO/DVzJEmz2vH4tqIPrZbNGoZBIk7ARUIEIZB9EN+GeDriyAbznUrAsutTXUdRtHPXeIW7jABrC
soWGYz991gh3uPjhF4bdpDAt7mqKEFqOl+RNxD98wlbGUaKUleK6W8rf4+Sny01Zc66XEa62HoHQ
xxIxFWiABTnBSJmk7REhgkbdbVnpm0DXtb+a3FxFgc8uZmFSf0HhYfLbCGfWg/JpPCSjMFH+sBVu
bJz7dma0ao27odoqjAgIDz4taFndZiGnQSr8r4ewY7MVeEu0JKj8dsWi7kX5eqg9uZkXA5Ut+3oE
oYFMtrAxOxHb2YMfkfO/kWO0mEUJPp0bDYu4jrde4B9PhgcanEi+ESSkVFgZiT9iQm2hHve9tRXI
bgwJug8tnK3nDI7Hy0KO/kE5yh6KCqhKC73Cqaeq5gZCO4RuCYrTMNmfZdYsBltG2nFu99SH65Zo
meN+4pA8jc8W6VZiXIU/zm10lNDB+MXcSQbOopEq6Lw87DvBPsLw61h21MOToJQfNzjsXiX3XWUJ
WdSzdBgEj0P+S33DIOBWtivs/xkVMmyaWHfrzqm9mlU1LuIHWhOujzdclraMy3WM1zuJ9vwHm8LV
5egBSkTHiRHin9T4ODdzZXbnnCaiwZjYI6lJ5PxhK1pZr18YAQcRcVDRYJvm+srKfZ8CdvVmpH/B
RpJJBTJE2/Lpuzlepm+8bTfhJXfjXNCO5AxSdirMidaGRyjP1ATpWtDRa3EKffkkyDyELEzwlkbi
asvFLYbvERjuQBouRvFyvqN+VLI8YFBSxkgXxtQTaia+tsm/vyRm+NezPWx8WfSjzTE/C5zCXqPp
VCe0P2ST3iIMM83V/K/axOe8LIsNxlhcB2V1hkWOtLN4K0sDFPiibzHI/RYanszoOkinjd30v0dZ
wJ9Lzc6NK9doxsA5Fh0xy9umfJ4pMKclbDmyEwz++WkDL00o5GVXm55mV7BFZi4Rni3HoSWkte7I
L6ge24tsTm7X7RRkuGws42HX4hf4sy2xwxQWv3XMat9crOmPp5bu0tMn6q2rY6D9+Hg49wUOfaYf
q21OvOtgeLLhpPcpE8FZ+6gWrBFDlITIaiSIJO1Ju2sq0ij8FfKMeZell0MAOFIXJHmOCJAHlS8e
O1UxZLR2Qq/GZjgaum7RcsHGSVHbJ9VS9JKXrR1pi7gsQt8/LMW4qWdsU9TlY08z5lLNl0uAfIz8
SFT90ohUu8/WrNG011hO/mF8mG0eCxPR3r7mideOGqVcBBGTmOkY2CbDt4jg06IT3GMLmuWCE7nJ
ykT3ONBV0b3BqeWAQN6NBoUrJ6T5mNrXLC1hzDX7PGrJun7dpm+NlS6ejFBn+ypPph964gXbHfN3
aV8R2UAFK9uziViaElvXxGSKGm1smT6P4uqt3w74rx71Vnc+d58s7V8vEs6JrY4dZyN3ovNlz6w7
rW852t/8sQmE5T3gdz0ozdfoFVfFX10C4JDOSr8iAFhapHtRxicf8ADYZiXYi55X0qrcTt8Lgjql
RaJ1cQce04THfL5LycV8rMTKnQfU10xfWqlUNlux2NsxB8oyy8kachGaTxI99p/jS8UX5cmrCbAP
T801mlfpIjF44owvi83VnX2YAyrBIh/g2cVtM8Nmh2LRrBLblQsxDJyEIP1D4LMSRsjrc9Ush+tK
B40TRh0r1Wdhap1c3UMLnzn1WZ5V5+LZXUAiqx4LQXem+hCcEdF6BoCXirDyEZdoHrgbhCXQrL45
chshvrKfNGEUwgAkjC45ncLtC/2k1kJrBx0DEreB7uLu6y1j/4mqlzkg+A2LH14YwR2MTyo/eIJ8
umpNGhnnabbbcFM+JmlA7FFrdswU4/97tPlxtDNzSaWIZjlmZBS9faGnbsG1tzeXjpZaYYQsNAxQ
Iw3C32c3oo94Ki18zrZ7G+xs9AHziz+XQokJUvHgpucfcC566MaYSLneRVCraQymGeRe7Q97lZt6
W38mZt0uHkaX9eQ1AsQo/pyFYHoiRqmnxHghVjrKismvRPTnBy6kZGogGT1ZxBjq+XHFsGw8tM83
3TaLgXP9KnIZoqaw6rTAgmgcMiGntYAT5cjUmZDbWBxPf3y1or4AkRRm0vx1nZiyqM0+JDL/kbWM
h3xDZByTAkrZg0W7RI+RYpVbC/F1AInekpmB9ry7ArjDCDwKnT83sbfOiih6B1QksewBzkCVW25A
wx27v1HCXXNE7N0iT6J7wWdXSYPgEWVACSqpJh//ciSDdk44+yhFWvPU81yhn02Ky1G6uMbRAJXX
SeO42kOWLTTY4e3ivqEH29Lbtin6ttu4OdjMPkua6H4fNYWHXhhVB/7MKzghc8kejJdOE7zJ1PRZ
nAnquzHnv7hHcd6SjwUoOvZPoATNOnGNx8fYgjYvwpPAxQj2NIr3HQHVwFNZN4Sx8dd+5hYRtp5x
rUOGIW4B3J1FtO9RTTRBViV4XL96CVhQeYrBc1UbE+HwFZwLgmqIvzeF4MWkuEU4K3qYdU7OzT3x
6A3oE2nm18priK0fX+AAo7pRwq208JacPZErdfYkOdrS8El0I6sKg8M6N4kZdxtSWtbHWaB60aVo
uC5cDiLVnfJOgZwVtkdcYetBkl6gIk/t8F61KCpidbcFJhv9aIU7lR/rzvMlz3vPJKbLHPFrR5aq
8IohyzRSJ9wisCy5zZEudZhyKzokECw2IhZDllxWEZLvrhZpFkRRVyYhVPUeCHPFX23ytG4S+FpG
/UQOpp0ZuZbtj5vjB6o02XdtdOzrm/xJikSkJ/4xPwNiwgJW7w2H6aNPnh8pLw7APnT/4BeBck3T
XCLAy3YAqjJaaA1+QjN9En4AUBO2/pIaNmQPoJMldJFOCVyy3nWSlu/+MSb7p7PzyMRtTsCOJ2fd
EeW2lZi2KLzKivTl+n7+2cwg77bvFKOWupxouvvHgZgIFCCMDLCsbZV26PZBWLXpEMxITrAYSky+
P4bsSntIfF7c/eikOVDNe8l3NTJ21COqgzX5MPJF4vsNKg739B2g1cr4w0s8Q2/BdV/T4wSMsTOo
hHpHbQ66W1SzDcCY2aQKKa6/Y5/e/B6e3G2pfPYLnXOJBaICmrLLZjOVSSFktzXEO3dhdzrQ+t7W
CRoTYHA8koTXqc9gpMiQMoHRdMJ1MQVdxAikOXIuBdwphOoM+4qWwxND4llxPbBtOJm4chprNa9B
ByljvlSBIv3QLyj9TttaG6rpLGwduJa1tFo8t0nzZGTJWHxJhToDgrT38qVJql59ZOAYnyQ4NV5H
k79tfGEBxH6piJLeYUNbICw7rSQK2qBOF+hGl/OUqh0FHcxpYFKN/GXIHPzGcrFyWqD38jHbgWPy
fQe0MhlExQdLHWEPTwo2S1R4JtxJ1abjVy3EfpHlx+o/hENtRVVhlXFQaiIAfxWNPcZomOBTsMF3
UYZnsrnANTP0xy8uh86AEVJo/mtEX38+eAIwd+zGRpeYrGW0fBNePVc6lnKwICOfaUH1iee7r6M8
8OP2kABYQBkCUFwl147IrWdQcjPSxF4M0s9MLrCohMqWyE5uAF+Uz0mZZQsQdasRBw5PmKIlnano
TLfJ/ukpL9AgV5vaEp1YofisnPiVWiN5kKF6S1OT1RRGjgcLq1rTqhIU3QdJzh63Pt4IU6Un+Ox+
wfl8DBG8zaJdB5wokAeQQs+72N3Q7hZRMr276lyZsJQADbcbAHPBI7XaemaybjwjH2GL64X9BERO
CWLh0KM6EyTGAbDZJWWdBO7RZVS1WSkRG1bUj977ESh2bgmBUMFiSjg1MQ+eGCH3//G+w6p13uZY
vrVZlSXslORLsLShV6v0oThFsLDUBPUEVJBFC1kr0Zv4z89qE9ott+F8pQVvxwrg2uSbuV3DwZxV
HTjvZntNfQAz/EYnj9OsvTK4QDze1dpqTKR8DgLOubg9XjB0RiauHktPgMZRp+n0mLawJ0KLQuLU
U7RsO0aG8riwTc3QCGXqfqr/b8w9ffYJAvJOHCTd6XO4LuwNHmbXaPyjAfbTNvshSDu9amuwGxHQ
Txd4zgqeXjuEuq3fEf2BPXYo81Hh+EA2NRuQaZfRd2a5T5DpqfkV4IknbuxxG+in76QM93hKpK9+
Veq7bnpKPwVAHOqalafDxMHTHr9dXQNo/MVu9XgQSihvscvawdXwiQDvGJOMU0H6GhpGIy/qq2+b
6nHGb8idX9aq9FOlypANDPMdB/OqTndDxIKaPy1kLrJkQiprzPx/DMzkEP9z6kBwY+tzTiikfatj
iuQvWuNh6m77rg6cUCLN7xTOUf8cf/Aho6bGQWj2epx/k6U2DWfeiOqT9Elc+sUQhzEBnnOLz966
sYyqtYAtMSmMNoQcFZXAS9AZiIV4Q82zHMnH+eMXmQ0xxv3dpZ+fPRi1r2aB85Js0rbBKNkkSHTM
YEQkE44SuOc4tzQ6T5XxF9nUStrO6YnhuwOuFnOejT78yZ8HJ07oQqcPkZ/S/XUzCSwPBf5D3lKZ
J5fDpKK/SoGinphSgCHF/qNwedbyRbh1Px9UlBTTZZt26VuO5IyrXE8wUFZHl+a9O5BlnpuBguVG
tGZGBaWcn1X9YBDnLqhTJPemjrrlv8QvQlHBI5eeQXZ5xaYgbe/+zzO8cJkb10GiW/Zn9+56YIDs
M18ShWNk1OMbAxu/geXbi8/Vv8fcf6/cJ+JNvfr9UsB/GiiJnqynpwvUxGLlia7xgULWFF9nRd6y
Ftp4ayyM06e5Jmef/2gs9pYcdMbgd8XLEGcuvqTj1K3xFpC66qsIoMBrD6OKdDux5TnDVUPtLkzc
LIQySFtdlqBrELMo3eyEDjI9+8/TxFJWUqq3kxL5BXH+XJ+BmoBmbPdbKxjeNOld7K4HINKrG2XB
Z3vDwuDlTTQYAxnQ3Rrclph+LHCGrolne0DW1/seFN67L2qXxiE24uJ4L0fRQgsKXhTW8gIvczzK
yIOWd82CBHbzGG8+iE6xBuc/XOEzk/kpnf5+/6qcjLFNgRcbxgxw3EPT42evjplGzYjc5CBO5DsY
OxOTtj1LP51bNuPnNZkvoMwIcyLCHpwMlG5g0/VPYN3lahC0nPn+cd32eHaoz0IQ/0x4cS8YeiMP
PEyppXOYoL8QxjTykBoW4+RgCqwe/s8BdfCuKj5/obsDitdDo5/5mbyowf36ziZGtohtDjrdU3T2
q4ovmbazMo2+cgnEMW5G/HtktOkkFnly3bqRVt3z1bvcX/4MdlKLtiDi0gx1G/4fEts3tC/VmNt+
HdLzWebvaj7qcJoAzbrUY2QQCVJbeF5CT6kmjMROPmRG+5FWAC7uVwaNPTEvQIu1ZCZ5kkHdyAI/
96sWXQOIlNG9c6ENNmyYDMgX3LQljGMD6qMd3qBsclVrQ4RbsInwNKbwWli325Gru34w31ko2Bpn
vvnkj8+uNCz5xK9VU9e3hoF3e7pa++xo3vnTN4URuBm2vpa+ukA89W7zdphswDPkB3CUPZfbLPM+
XKgShUKGqeBKA2xFMMxsrpRPPX7Lbud8GpeDbnvK15D3u3u1OIIol4/Yg3CkE9QBtIxHTyUbg8c+
WsKk4aeqPS8RYly46IyaSAGum7UJ09WYhDwcvBnFDUB3JQHUBGGG5y0Tgd97hSTwflKKpVkWg9In
5IyFJ48fGyD1jfjvwRdpzuUEnaB8zmsSuEorYsfsj+HL78dph5DXUBzcRz2UE4AEcj07sR8n2u/Z
Gpb9xlJffDAvfp0uW555X0uTusV3LboqjsmeSRslaVFw2P/lDevuP+g6LcR/88bPI4yQQMjAospK
VLzJIQmRMi1ij1bxwXLRIuWmHArauke7CQUbqZv92cb8zQkGuHw9WOMPOfyky7cMsAMFV4odqWfC
k19MEVpYV1V34FpW0xmORN9/mtGo974BMRDH+JCbAyNaMAEIcd1ZZqQLCKONcpPO6LxNUYvHqlQj
uAXh8Xuww8eGr0otUluY4YYfLHzBcCrWQWfSNg4IWsDmt9L4Pc+yELfoMnEg6XA5tt79yDz+VIO6
MrJHEsgFGvnoTuVquJtRvP/Wg4ubMIrk6IxSk2I0XA8Whf8x55p0QbPVODxbEOyOTyR14JV2SZ/X
qgufmYBKiJD0T62Cx8rUrPTaVAr36gj8Xexrlqk2aoPSMxyxkK8kBqBr5XCeDpdTxDiNKhMmw9kE
vkqldBqFp1V0SYwJJ/0pyzzMLNX4m6UTC8VWNOIcSVpvi2xcPXiB3WcMKnEr6KgDxhhbwx8uHac4
l+16qT8jVq1HDwH5eJc/rz8CKmjqf74RU5oExruzr3m/9NUIz6COqQVMeObGG36b4jx6OKsQBPby
7mCZsoGZMniyA2ZssvcDLOVDAz5f4S29cP8zt+Ef+YmdBcqlAI3sczURCspx0vpZlCbdZMeMa//x
HkKlEk+PXFIanJgtLTLZj7K+dM9rpkRzd2rF3eg31SeUnUmYA4kFVRW1rsEFdjgby+L2ihKfkm8R
Z/0OPMhI/+Y6zj54hhc8RTM4uZBCaBj+4aM0rDx/bGGnMTN+AiJcOQlLi2WFBrmdU8+E+z/ErgjK
FWVMksbVVfT4tT2sT99vb1WaohMZpoJJ0gCLEnL9AQa9li62D0OkW2E8F1Br7HUNFagyCpXT1KM4
cd0/N6HPFedmbhpADiUAEXp2+GroQhsmskV402BaFOzjIX61xaW9zs6d0BHdPYBbf0symkx1ndox
W6iyRuwULmlfrOMKuLZm4ibm+f7fJQNbi83g8+PZi8zk9kKZvRfuC5x/zJeykK6/utDnjjauENMH
TYFgc1oxCt1awhnZHxyG4OoRextsVKaxAZvdse4+zQ2bZ4+MreRcE4l+B0d8HVbFgUcmfx4VNoev
Fa2pDLUgIrvlbkILXKHvXic11zXiFPPvEO/dl0cJIcn9PNAgPyk8S4u/qYnxP/8nd1XG9n0RD0DV
y4IDuVEURt/lKff7iWmx6ITNyoyMUzT518UThEg0umHiN9du0V0SOVFJHnShDja+Cc1BCq4R8tqy
aIGth9391kdWs8TiO0EJvS2BpxfPYnrTTFmlkgvocbqG/9NomqC7g4O84EF1JdPP22KKx2OJ+27r
XGWMzpcKfGUCbW1DVmIIzOrdMEcku8e5vMsqPvHWF33hNjpCAI4CmxMy1XX5f5vZqxvAhrRKZfOU
H5zqZZmKrN5po07Djc3KEXUR4OcdaRRnClCPNk3jwhE1IA72dm66L91X911Hapm+d1Dk+xK65qqb
qquoPhHkO3QsYQega8NQmDMbD+F895DNZR/pVfoH1nNz+DMrr03uvwC/l3afiTgW1TLfKdoDH2rZ
vOCJTpXQVbAvCLZGzqnO+fcEF2TViSTZhJHykAu/JjiXSv3H39QiWlI+0WvsXZNPgb/39ueJDma6
cTLC03LqQvBFkTwgogpcCY/MJ4D/mLvYihswM8SnJJVioonPc2YzVxxlJ4w9NGMURvu6fPyXIUoK
HkYVDT5BZKlV598oZVOBfsbWVY6iAUCOrzxtp9HzVQ9RhBC67fJ9thix0hdUcBfHQotKtN/gIRiQ
2EMyAqh2rKaJOod+0rhS7Fc1pOWkHz8MszQiIPSiKZDHIPvFQynkiWENPztfJNUvzDcoXtnYuSKs
4gG5xWuLU3XnARyEKJzDSHpXnQ3CEB9U9fl6sVJhikzO9tXdTQurU4Xd0wbkzrgsTaVLNTrdUIOz
2os3yzcUn+AoDeSaTuFvuKROMqrQ3R/IjvHWiuQLAI2sxVghOzXkF+oYC6/Lw0qEc+4HDjLFfN9j
NX/DaEO2NXXQXSMGdPm4xWy5QMFavZQ/BE9CD05Hc3gDk9Z12ZQSJZoiWJ74u/b1b7QHYZsiCYTS
0B7l8kcIaigYEGYpAR33x3rYfg0MbgTUQRwCcuF4XDtpa96w7IA/M6Y2lwZJDCf/j/DZR04wJWUH
VAfInxGzGq4vJaoODgWsvLzLlK/0EMMcT1mqTAXYmfcm3KolKGkaijsgJqfRF2zMY4BlyFMagz8E
/CpWYFG3CosL4Yvpr7YuQ6UvZ1ah39p6g86bE0cSJ1peEHG1sckCgy0WC86wLXgCWGlqjRR1GnxI
pEOg3c97V7uGr7o4sTqDBZVJgf3DUB5DRFuUamIbMa1suEPbtNY2+83i3cLZOAwhJZMam/ien0Td
ZAsI+d29o0cKOUDIBnezRkapG/vfRf7zXSp3sVdRBxSBx7jjGunNP9TkEqixe0phhuP22+AdJiXy
rY1Y2sWOM1FQKF2lmXO3s7qBi+FKoyn8kjfpdBQvlCaSrsoEuNNZ+3NSDO2ySe9bVsxInXFgUWcF
2hx4nZFzk8lx+YfLczsXkRvjDiTSd9mnUoLU+gH8oeULOnBDMD8fls52vnIcHlSvhPKiMrgjpm4x
MH2Sj7OgUTfwcBL5Fnny3C4OoTywj6BSr2oBLHCcBk3PMkDd81D5L7xyOlQyEejd+Y9vpI141EZw
nGRvhuvDGNZIwcbow2n9gpfVFnyZqOgHWblYBAyE1Kt7mUqp0U+yFa1zOgJtAdYmDOa0Y94Oa1IX
tEOFY/yWYZ0b3L8441fsjB27cFGljD8WDNogAZJ8GKLUg4DwyTwj6zB6Pc7e4Y7C3XxXg/GfphPv
2ndg+qv8S6b168hw+oLAFMRTcBSbK+Jza0GafwmAQzs5lJLuTK64mgqqyxbANNEn1Xoz2qknHQn3
lmfv5ghzHcOSfU0KYjNIaX+x7TvnreLrVkDBByRdObY8Cx4oZW2Yq2QLvcFKOzu/v1T9XnhnSOyO
fQ+Fmz7G26T5w4PXWto/QxY98MjZjAPcwEH5UEOP5Rib10xdMIf2Xc34s+07nKgekHB2k/R8BL3G
vkh0qhwMynWnqsmReQIehOgA1cKi/esvd3RI5cqIGyi8d1r3yRtLxkzq83zY4PssqrLBwyAEBzHG
+fmQPkn4LPvfReHDTIiT+US68MXp0wIBTRxUWbSTY7TsgjFIswgCKkSwHA/BYHqJV6tYYka8nFw8
d55JloBw1LNfYeoVZn1qQojji0qqgpiGTNiOY/IdPoN/s01M7PnGjTuSdiOQ2XEEcX/7aR6X56NC
8XkNXDn37bewp0p9uzNtKlzodspXbZXLDfvnTApIUEsfxcLW6kBS9NtHSTmiC8w0Qh884qlr2HRW
YhfDkwTOWfjZRo4WsG8S7AtoIJmmofyVR8NukDEV1vChYLDnw3Zk0saQ9AwaZlLAcpGOLPeOYC++
umGK6zbAnyl9s5zdzXEM5+9e22oa297kFTh6YmevrEjB7MHq42yJPxsgdIO/VxkDZ4jxUqZlcWzC
t2RCtwZF21oS7rwkkZxjP/NXVd2WQLRXsqzHWzqGlRW1cgKMhDAF88gysKAk3f5sl6byDZ3UC4Sf
M4b3+b0n8plmadngSwvXkFWJgGVCEfF8RhdL1GvMBeUpcEO/0kmUaltkHT2RzaOBUOCeu34a+I11
nxSq+ePCq1vprnYJcB7DmEf4WVKk1ebh8tcT+S/aOD6xdPilJMMq8PXuYP4jTqjVfyQN4Nei6rpC
RWE7yBhPSwL0r+MQyDJvwLtze99acg8mOMlM/aig7uDxtiroKyaeCDK/NEx1T4t1e+Ror28GY4x6
os/sVJY8QYsKn/t+3fJUMeZjUu96OU1rxS1gbMFyQU3rJ116vJGM2dO3PD98pJIrZmWNW5M8xwJD
MjMPE0E58DLgTD3DTTtXmTryF205nW0OkWYQIGOysNcStsdHl4GWVD+90jgMszyx/Anj0k9oGMNv
TyuuBiGkb58gTuij0nbPSM04kbL05n14P+TfZWxJ00BHb85GGO1iEoPFeQxYyRbq1nNVtCf7o7VY
IY48x3uIKF63+Ah3dX3+NL0LOFDCVdRYDku5jJT7fhQuQAw37PG7KeH8I9QQ1h2KXAxVceJyp0Ag
ljTuavU1Dk5Yp3NJvDK/Q4zuDKNAlLTCOWepnllFHFVgLVBfQJZnpL5M6oex8t6ZttORNYYr8Php
lLf0c3EUV+FAKlyQsnOpWaozMuTU+UUyB7N59ZiiV8l+zKvAS8zo8sdrVdJfx4dzxWxbgyhLXMGj
g+x1wbACzpw9y4HeaTDOPbZ4F8qvGpOiD+RBKobSLZrvlY/hfJnE/zPjCGsdQOcsqqMoTL75n/7N
ESy3I9qm6NfD2/z9qloD87vgpeT5AebTVROAyXO0Z8PVPMjCKqxdSo8cwVODrH71ZO87BpcwGEH3
gVBxVVIoxjubnIOV1e8I75OW94XY5MRF/rRTlzylIRpuit31pCgCmKPUSdXzdLfx4A9LRGD5Wsfk
4jMWANFprSQvfAsCh5y4RWB34h+pKHSxhgiRmBSXaBLlcSiLZbZMLGdDJlhM6HrfhoALmqccKKOK
uIv3yxYYQ5gj9YrmdSoxkKRNxWoUmwhy8Y6lO2L34qhECIkoI4tvA9utJZMukEaMY4UDyVN7LO2S
V+xH6pFAVDUcjrfpy2oaaNRdXZHZxEHtebOAWEzcHAtMBddRigh7RqgTzHrNGxidTDwPj/Ch4neL
NUG3J75DB54Ylijz8nEZbLnL/tquF12hooasLIigGGP9W/vaAfRsmeusnhpwtmULKNwzDibfk7Bz
97f9LNvE4V74iI62k5QBeF/7GFpdXxGsXtMWXy1Vndf8OS/wJjoX9Op4XqjKPWR9xBF7F1PCgLkR
KF+MYO3Pu1l4AcrYaxoTugKHyQt3t3AQbN2tqyMhSMttPuaWsedttD+BwPgU6fpOx+Vp/SF5u9zm
mQhySoJCT6sF3KrWaFWyJrS6o1OtLvqbvRrs6f6cU/Wcjl8fREhhUxWxbM9EqqSeqUQ5q2hj/Yc9
byrfhMe2qusyXD4T3S1ZgS3awCTrUgvgR2b86sWlfF39fHGM0ARiN8Swung7wgN3Pb4LaeEBvcYg
KAuYvx5Ef3mfMouxK2uY7l9gpSqnOXajsgeozfRO30oWocdCI6P/AXtvNOifspALAAv+fKFaYWyT
Xpfos/ogc/m6XSR/1jWLyNnmd5K5lE4mrLQhwRuQs6ASzmNzbw4caE/DxAZ6XnNDtjxaKNe8PVUf
erV3HA4FFew5n9uSma8G0nQUawbKDmbUvRoCoXrl/66t3wv7iDHzfJKseLczvWMUlbco3H3mQfKB
pK/J7S+Hxj6pCnpYxa+aeKJPZMGFNeRBCImG0Hcip7aUvIUBZpf+CyLOgyzaZuoVvP3iCRFY7RdD
srJ+RksxNDuSQUm2M/csSinM3fSncX7uRCrlVWIDRvtv0S8Rz4iuk6cYhmSdK0UjyxO8jgvW9Ss9
1ZOvqOTg8mJN06nIq/kMqjWU1NP13VAvW8TShruRg45B7MSbL8nBiITAmu1s/vh6fIQsHZzlzmsJ
u0c0mzBKyHnYV8HQDmVY342FLFFinPbImkxYoG+pcs11msnLoKERWd2rG73vn7mJXLbCHWfV5fuZ
R5o0w9Hs7PXB19Xx1Ge7L4fSOei5bbK3UjBhbHn4MzNfLa+spvM7tgJ97YU1axkIkSyGplgrmnA3
Q0Bo0sYTSfBWcpRQO8A4Kol7+FcDlQTwk4nFapZ+PuFFz8ECJg7fYVvBPoPcb7Vvvdolm0JYT4Q8
Y3JN3oCIp9e1XgfhW4Gshv9byRBwoO1jxeHIPWFjqlodzRRYRapyEBBiB+YdZzo6WCawmA9a8p2x
nt2zIabJuk03QwAgi88XodGJ++hcSf3MhwlfZdhfF9XF5fzteBk1BmopHbTOIsp8j94e2+a/Lxno
nnRbsEXtRwpwbMgAIfL8GJB1Bh6xqwXdN8PkmYQUR8lyrpHe9dMlop1Pb3NsBDl5vS1Z6xwSfNjg
YWszZkue/ACMfnUYKrClzaThnW6LSY8jReRQ1zJAVFDq4hmMnI7aTBZXEEinH5w/2R4JEbw1ftlg
iLzCBBMAhJJtfrnglTpnmU0GD80+oJWsoxnVX43MACzeWDLoMX748obh0cci8Da1nd+B8kWBhorN
FMSOjII6YJZuibq78W2PyKgd4BL/+GoRhee1gdY0LUc9JCFYll38ftcxDKUfrbu3vjJRD2Ed0hXl
koM9PgDEfSqE8g61U8b9ITCTm6XGe5Uc8xRYGaUHhJwZAM2EG4xdjeodX/ghB5c7bJ0efBBqhDRW
o66t1LwCFLD7awvhnG6HePUY1UJO07XjKhQN7K4m24p+ZLH+a4HYwHPGfgafFxFgE2vLkYhSeRgE
Rb0FZc9FQvYSEELsD0RX5wnnusSdD0pyKfDpXZMbv5Kg9HPfLkfSatdtN0hFqRA0UJKEKVv56GT9
kWPskyXnNIfjE1W8/ChC9htswk2Lb/BMEWODDIrsBrlmFV6QHn6/NtDBQ1LawRBT0r6QwMoHb6t9
+v+bgP8bmx37XH59Sg8Qv+LLOx5lhSVsu1/ygx1C8b7hhun89rASPaKhfLLMOLC+UlJon2Dk4Sr0
FA7EgMme6cxX6XrXXHnHHrSz1TuAUMmBf9cwJMPU517CA4brbXEkTmUjReHVD3yXS4IwNu3vo4d0
yABepori/dLXsIS6i5mY2sXcAfiapw3gZTh5qIe7qJok3C9Fr9oybSKaDzB9SDhMYTUaphlvCOTt
038AMsv0aYzV/azpXEuNyObO4t/SQ3M+oQZsW//+aS4+/+20GQNAvrMEz2kMayVWOkkSj+A/Mj+b
3qUvSBR2fWPDkFlVRMia53T0c0aOVYmsjUQu0YJ4Lm74lk2Iefk+iFURKJpDQ8Dkx2O+hUe9CuNP
+B2t28OtBI2dFHc81rdvOqChJUZirWJSwOzxSgXzGW3yf3p9QJ/liMK61uVFUHkgyUhKDTVL0tIZ
JfRlHH2PdljIkfjbEmFkZbfPLaLG8PlqWg8ieAueAZ7Y+pZ/WgMT6jtrw7Tdasfg5fRle9bMKhat
9vNEsKO84R0RoifjUG2v25XibX94jj0UlfYNyII3swjytN4QShSD32mpp8UU8oGJBV1I6/guntfJ
xkDcp023IR62nPio1cjrkBXPLg6Dyjh/2Q66l4cNFsnx4B/CLmDFBwWDdt7ihKdc5gYPViKo/6aj
FISd0MnrMbIVKx8RBsP94CBqtfqDafDh+JC5LBgbOb3yUX8F6rLACvsqc3Hf/Ucy+LMrhlkWylHi
5Dtu4T99tdj3wAt0wIihCOEe3s7ECqDJ5i/WTu1K4cae0W2xSyxAbTv5kI+idtBw4tYdDLrVytq3
9HHYFH+NTizCjhPfNUb2yPQ6L54ADhvOUGSJLeGplwcAcLXydhtMPqR4PQfZYnk4oW7lvyNU0ush
hb9GCSO3r9kNNZALfnqhuQ3HSYBzHAixDk/9YxKAjjGxGf/Bpg/z9d6wcTECtHkyJGHJox0zrHnP
Uf3pk6IHTpyOXVrmvAkRj+SMBNuLAq8Z5MNEAXJkfPitIs5aQRCG5iA/bzfMxDPDlrJnVrn6Hct1
BHJ6q5ykXKDkfat5KVeuDJNrvAs4Mcy4AN4hJ7OyHNXTlJHkQ+nNQwBVt9ZyLOvAKPLlQAodbjvt
x1g1xOyklPyLv5gNMd58xZ5sVLN5isqDjFwlUGEV1h8BXpcfaMcaix0s3q3/nFW7OILv/UARs1RN
PITJv9sEF+YwbG198wNyJbXmIZ9FUamR537x/TeJvnH7rUS0oVlcB431ZeUhx1gLnM+7/BlBR9JJ
jM8NErIisnqmJbyWYcEMDw0lZx6BLIKPVlrst0ajFOpAt/NeHrk+VUupVxmXDD4Vo/kOi1Ui64Gj
7UnNcDRNExoHf+T1VY0gY9aIPa/AmslKPSWQEkGqz7G91YwX5PhwJcacU3nvaFnWpvld6tKDyE+v
YVIiFIiqxZsD4kW1if9b8eoklK1ucK9aij5NHx4j/W2oZXjETAdJht3LhLQnFNJ6//lt3sS6HxhT
qp4eyxkP+EslRAdIsLi7R9tOBuI1BoS3ZmPNXXL/mUpJFMT73aL3Wu2uNAKWoOsmB8ezHPoUDwH4
mT72NIurq/4zEjBgkcWNPqw5/7SFM/lBYTr9A8uxv6nC0TX2rMjwbxRgWYZ1w4OmvUgoFvujMDQX
/YpDSAd3veAWLN0SnXuAJnY290u+gYvfoOmfSEhaUmW4aKzy6s8befT+z4DToeumoQiI8ePvHNXl
ds3Ccwx65ngzLnb0QQZ4jloSa8NWORW0yGA1Cwbhh145c/DO+8pH6S2q/8KA545SiPUGYUpP3E/j
Xb0pALIPFURoRO9snHIrrf7SwxbdouHrbY1DNB1p2od53bFcXe5UCuEEymCuX+OD930Q6QYSlGwE
L3Hq+ZaVw5QPdTTuGv7T32WOEHNwD4DJkrPFZy/pLneCmAb651a0XzTBnPUefRn+7BsR2tJLiEwU
nh6m2fhIzeEJNrptxeVuWdn2ofTeCXv+EmPzS4h7XkgbsGysKO6MCJQHPCPFMvCGddvGTH1fahU2
8NwcBJ2d+dDn0HazBE85VGtGk2aLnIyOX4/ZSBb9xTTgK9azjcbIIUYmHPgqwQUP7aOiVUFbS8AM
aUg/NGEtvgBHdRMnpZfJTSrN0sOBHARm6pY9ZSuje0qTEBMJpWd65/jsW7jLBahlUd62HTSaShYX
FgRML9oCRPUjBYNNVOcb/1k+izGsr3cm6WRk9jWLMcz/iWaAqQ95nw1Ps14Ve2Ge1p3aGFHbRFc0
0ihoN+ub6i5I+5VqsWlPi8OdmJtmcICqaF+gmL8D2ALES/BFD7rH85b3wcSBglbPhIwICxlf5zdE
AXo9NxnPUxRPnvScdAYNHQ4XXB56kDOEh0KdAsW+HfchVq+/Q+2o4MgV7g59wsNdrjSK2ux9s7ya
7DEO5hJAOqQESgkhgbFE17jkCTAFMEpX5mGkdPmskL3Nb6aibPqnhlH0FNw34vOiiQ4DlFdBYY+O
F6J7fPEc5CW8vu2L49qTVm/d6w9TeylRPwk6Y0x2Zf0eLnQ6KlIUme/eJVp+WXnOblPXjecbLLBL
RJ7N+Frwwh5jdwgojRc9UueOhRamjXCh2wIiiTOFahyvOmXeTO55mV7COFpmXFa2xv1q8i3AaCTJ
tk+uaF5GUiE2gggaAHTSpzRMJvc1U5D3lJx3zMTRzg3sXcGUaVTI5PUMw1VfF6NbAx/CLTGMW9f5
reSaHuPfLc41W0tFub6bKWdxetF0RPKf5RLme9d0t6QmUmPOVxY6nk/jgs2yrFTxZi3XglPM/XPw
ONYHvqA63KLpvklBxHDvQGqPRQgC69lBHTTw2wgJOErjAV8mNIHk1oCRPnhcs4CS1BeNJ7CSnUQr
Y1+q/aWypoaPHcPp+VjplW0wEYiF+F1ERLde9GZdi39OusWKaiK9wf0cce0wupLkRViqUJFlCNca
D3xB3Qc5Flg8of6OhDgk4KpUoWtmjgN78oqU38kbKkeW0r9G5gV+J8l9ypy7USPZn7GySJI/in3G
JSe6HVK6KwZZMQJ1X21/dlYrN6QJb2zwPQamaSBRswEG2rqKLwvB4N7x2ALJJQmJO2BObQHemBQU
c0++Mp8lLSnGFRpd+f+XU9ZelRFBlqvbfRqvXLNFu8J/liZ5rQ5tto3vCkhgD3JH36c8F0I4BPYK
92w+jtXBLLa8tD6SZ/4rEBveWRv8MqVt4U0YIsB1ICWLIuT/SK4uyrDICUEq5qzkniNNSFJamY9n
yKMWpYpiV/cp2QOyj+SkMTsTZ4PfjXQqP2ddNygIl8/pEpn/VPnlynYCBCDEOlxv7TwOWUL8ySfA
L2FL0SGGlLxf+APR6698XynjPvMbONYxk+y3AvBYfxyg/7rflDSjacVZmw3YoPkUoLVPGJJMaARj
ZDEPCxJhmrYHVmTqc1H+GXoZAEuf5ZI2/M/EiE/DcCewSw2k7LvS+YZQyzwUV3KnaqOrzgVq78LA
+0nNzO0ch+Hok4S34cfQf8G9z9S3TTb9Fp7l85EouHgWN6ZNok1Uu/9EMoTSmYNoc+9r0qxNWYZI
MerJp5i+/gFWJr4Ng0WfnUJW3GNmkvGIquB7xS6JZYcbUbvYecib6Tz8HgAPa4/YzLTRNSG2tFR2
Au80TedMc+NWTQ+cRiManm3z+YvJ6ykcGUqNpj6vzrhGbY9uo3V+zK0ljL6vItdVBWyhmrGKi5H4
PzctkCMv3doi/cn6Ff2x6pP9kw4CxUyIQFdprVeo58v7xnhyAjKICT5aabAB+ki8w5Wtavzer1Rt
CnVh5Ni036qFbN+q+fyPjPa4cX/HjcSDq9F+DGmht4BCaP+hPdT89PAMjodIHR0NJSWi0vitOayE
eoOhUNTJ1dKsofXAlgR4A10WXd9axebqhg1QGVPxSR4ZiI0D+W/AAuG24nNVsJNe/Jfz0dIIbiL9
VgXxHSRZk5nMthy0OYMme0D5i0Yu7ew/V2Fvuq/RaQtvC3w6qbEj0jz/IoE9mfIHakPOrrsFvSSq
YmlctRQGSSV80swu8fZ/uoKBhnBNrMAWU3gCEuLJBsYIlKnDbDK7zhOpVYUf3SPRf9EGUKkslpMU
DQT4oDQUFy+rvfIENxbsFfbmsVp40BQEVMXvPaMNRizUCBfbYEkdr9W8RO8KzFrsNQuzi0RhwuDa
D6EoO5pDZ8sbMZImJSt+oeSl9ijHvEeP37rXHZgH1GhB9MxyrJHagTHn7F0UoCpiyvWgeGUDxx51
A2FcgrLrXCei0JFzQEpuOjMllIBxEDacTkLdICbe+MJ4xU2+C027LxCoDbj605EsV7NCI3GC16fZ
56zlO9fseOMYWHu15bfu70FkZmYC7UyF5jhC/kQlK4QSPSbjzzvDDh0T4ws/QBpC+vSdQgEpIUVl
Pa8+uK+EFWDnfzKtO+L17a2rugCOyaozHutj0/oM3b3ZmZt1ikpGHraJ+F6r9WQI1Iah608+jmvh
CQHEXXNvnxUmi36WkbaCo4vZeYdjMRFFuful0Wsqb3YNvcLrMpan7vcVsTjCBwqmCyHTnKqVCkXK
3vJV4OZsgoj51nuHidXyPynodYj/8UVqUr4WXeEghu5Sp+nOXjHQG3KYSmuMuNIw7S8Jwz1BjPF4
nN4nn/032LoL2yRCwYNKjDXbPVwUJW0KQ5h9KtSH73FJpCkoxsHuHFD3zkPq/m5ahL8MDStYJAg4
ZUbKPEx6lNun8QmiYzUZc3y1FwvdVcM2MNLtr5DM7aABWwpTtU3fSJBUuy4OhJqOq60M539GwNYS
sK8p8vr8WrfLNLO/gErzaVi1fOv3/TdkEjZOyKSpjEtw6bUsL0d/mBOxeatKw5kp7fpAmVG4Pq+C
OsyD6pQbFdyAUf98/csa54dv7jn6/EwRXkkmz6YzuE7FdI4B2f3rzT5rWywlactEomkCYO1pFJaG
JEn8DYmIQsPuDwJ1Z8hSkIKjD2xoRe73S/QzQ4/7Fo0I/c/DRn563qipgF4XgXsVXviVONga+NQh
yOHV4sMo0Hx/8JlClMiFkOsyKhhzSdXuvr/yKN6ChqCD2jQncRM9FfuzyW6W9QfOsFsYxw120q4r
rwxNv62IZskZkweJsVGI09OEkYa6AqWmudLUYz+Irm3wv1RY9VYqRqk9GOpW3qs/+05SpPque6ah
LLrZ0hdlmJ0OwnCSJViv2CEDWkMvMweLbEOpWEIEn6RaCunwc7lKA2Q6jhif9AvlCmp3xIiRfNLL
ZOep5m1UhfF32i77SaDwNCXgpEMSW4CGw/eVqtQWh792iyVNXr4EqQshrkBipKj8SzQRy03yhWvG
e96y/vxw0t/WdW6nj+fAAlxvtnbpvQtoRjmcQbMOhg9Wd0lXo6hPvXRPT+WSr7AoiceJFevs8gFa
OdXSaGPA9o3bHbG0SkpJka4K1nwx2EvEJ4YNSnilEE7WWxhrzb4GILUgmv8+YWhuhm1c6FLkr3ax
vca5ni2Uo478pI/XV8ohfQMbwqKnjWcLUfR7tpdFCeAAE1qxIW7yYfhjMmNZlNMWaNDJOhRG9pWm
z0fCrnXQltsfvzRy+GrwyO+GTUXlz6ZfAGLHCyD+OCjcTH0Tm6lm2RL6LyZlhsTUxX3FIaPWX01a
PCC2EptL4DBOYvP5vFi28dNWmx7OuMs16xFMwi/DlozXKnY5Rjloo3UjNJ0MOMirJpH/FGVo/lEx
2g1VOcx2kaftpse0xlJGhVZouj4HIuW09CG+u0YTT6qcLUSc0LQDuiQTHmAJYtSqFM106vSiffvY
rI0ixU7uQkqcD9wFZLPRmNj/++rP42iBxSoYXyXjZX5Khq+zqK/6fvd+kaw4jBHxX2OLLriLhOSk
OSSs8Wq7lMPohjzcbvkJIu9mojRuZ+mRKwZdZLdLOGJktduT96vmHz6KA5eN2DHnJ4BOAmcZ66tL
pQCn1lI/c+6NqpZD2BS2oAlF0sfrqRHC3O8aiieTp0yV2uL5kf2bV33K6l2MoQ7F8IHLu3cKX4OP
MtA1kWdOuA8wM10J7Q+BsmkPto+PPYztXkYwmlhiMOnXx88s/MYH7gaeolT7e96JlpS8xXs7bSvn
8CiUJorcD/LDKqLEGIDNzrr1RsXmuxzagfp2AI+nlGkZGHfvOkcgjUphFx67eqMtM7DyvR4l0/wP
hNa5RZsZZswG1W8XoFYROsCgF3mV+QxrPyfrbO4ziEs68c8W3cZrdqq8JrJmac5pMkmAy90vRFC8
QFfG6VytpCWv0DOUferlSENxz92ZmprsSqmKtPPlg6uLyXVFZZdP8a4rYcAV8kTeou9TpG2gY6Fg
aNPa0cjiTJ/Ion2cyJ/BJYNXVb24sozfWsg9nN/olMRDHJabdD0ZCz+CUpojIJmjqO/EUDkG8dhH
bi6Hpfl4pXtcULwNAq1U3wjEbn+HXDmo1D8eytY4BPn/5Z8rGUarWgR5ORdTwS8VsgcxrxIhbZGS
5yYV74Qn8tu0xseOPxz7jdbT0su9AJ/l3oQDPh7dgrHOVlTctJQ7iYm3VML7Y1UHpdSlY0gpSq2h
iYpeVqy7CisFzwv9HcRIu0uLSLfUeLkLHRCoCKR+nwLgxLWr7mpYoDrnep0gsRotneH+Qvb1i9u3
RjLRGkuEGhtxkYtXGQUzsiNYi8ebVvX5QybqibuS83IIfaeHEkeCBz7aUNUcEQBSMsQToKSDVQ4D
x7DZJvVefvieK1XZVn00nxe0dG6MbofW3csg3Ov9uy4X9o5ghuw+8AHAj4DuPwCFuOJHHalm471o
rRwbkd9OsJAdq165VW17fNJN0VMkeBdrSQjXH7SabUCE8JF3Um3gFClJ/Nco0LlCo1RvzojHf4zA
ZaJmIxAwh3lKbd0/JwiEA3YJEO2Gk/jDl8g/HTOvNn1Wsgm2Q+8qeKIpNwKFFg2LOjKhyf/77Xsn
GERBARkWUYRhHGLMZhBAVugiJSeCTrrxW/kZ+WE8IBNTo5evyKIbPncFJqjVmN+bdIZXMRrrsgjv
EN5n471CS/vsqaUZCNMlVz0ROwQb+XPRhfb9zYHmHnvXzv77jcdb+SalLGtaKNap+ap+MoVQ5Ch7
YQmyiljebsObyd148muvufPI4QlgxskW02GBbDTThdoN9DroDIdGbZZ42dJCtpWawqD0h2QBdlba
V1y2E4SILVuVXn7W0B1F14FoGYrJA0KY+9RmFzPPejoYC4rIZdYKQjv8usyX7eXpPGfL5iPMUwPV
cSkQqigFWI9QseZppU6nPYqTL1cTc+Y3qqBvd0b1eghIPBbkOYaLJh00vwiuZimPVaImtRQbHtkD
PwAhjClg4RTWVoQEpcWK4oLGm0QtGFZzGuuFfsH1ScIPq6+S2P7aPr/96F/y37g7BpIbOAbJwzwi
nb4r6TrV+NPe93+VE/dUSzZtTHtg1fSthBRU4djiXJmdhFJsNvRoL5aRs12iwyhjLqFzGImCphqb
eWS3SAmlsIU+cz3rdMXyw2AnYeD5zf5bCgx3Zbkh8hDH+1s1XqeWnXNStOc9+j3ISwBecAdcHjbV
//Vmf4sYordJbKwlBql2FrziOmK8gUgGC72qS/3jsJldVH68sFubvH+lA6fHZussjA4sEaFxdyf7
mmgC8eLfb+KFrBRyo5j1qsXYINlH/V0acVDZ3+GpsLrYO6bt0qLrFKPR1y/AfC7zV4e6aLhyItDp
37ghyaF1g+kyRmk84w3npM9e1QGLI2G3Uvi2WEp5skhSzavD69Tf0NaZjY554oUlFqmbSizv8/vp
eQRoz4cy4xc+MlD5Y5c0/x1AdXAY7O+C1xkTAiDhbF0FCiQeUOqJ9f5MRUN32H1CDVH1thbNFKlp
J0Iz0LaiiP0Jz6GO1S7//99VrK+zjmGmGxgzKRMH2JZ8zUZNPav61HubhBmb5QHzdelAH4WLrk+v
EsTbNFDjHuDyc4fXOWEJxPbygUIzAhsQdwQkBeCI/9qIubrqVRVUfZu8O6d8cDOHuK6bPw+4O6la
L6kPCa7/bMffBz1A/yBynt3gJYQZCZktyS59shvnsu2Jbl5h3A3tDzxEZ6cyNCTZfsUaAhVfwR+E
A1yygMeCD4WANpDhiJG59LlSM2svRcI5O4vaT6VmuTRc4jEHwFcmHjUgyrLiUJMTYGaeGHBO8dJb
kVc0EY34fEEoNQ5rTMnmkfc9PXZMaFfAFXyHloQRMBSXYF0T+JZzSi1JjHCb2YcIPQ7zXqf/iPWj
5z8V5nhNnXAYwoN/F3Z83P47CEsaYP4hh69FMQLzIi0ofjAXr69vAivdY2md4BqE/3oeLlpGQoF5
qUKnu7IK9gp9dXPvDPXQIba0mlzdHGYd+ZypM7K1mJ+6OA9daVtU4rJbi/LvOFCx223M41xtvxPy
gnbhZCjE4x5IvKHscisMbXAWdR3BdJP9d/QfNoNdCgaRyMMWjFGy0GGIIMbIGN4Qz8cBWpvjm55r
pBcMO4g2mIJI/DbWHj5f/43bGfEbvXNidwdgNZ/asBLmhCe4c/4/y8XlQlgq9sR5lzbrl0UmnijA
tBYxo5JWalLLOroZZN/BF9Iw9/ixFpb1rGdj9vxWWoG0th3xBQ4dHGSUpBbqRUaW/E3C+YsPCyAL
jbE8XTjnkRte1GruMvtCwqbISZuxh+P5Mpfe3LcxYvE7LHxBGkhVIrN44+9rPyYE1g5OpW4EDO/h
tEqeucVMrOGEnRFIocoS1M0vZSGK5aoFpCgYRRcJgoh8UNa0ZdIv3iYf/zy0AU2ak1/xZPpOogOu
h5i04k/NsklFjVlWDbW+W70ijdDF02/PFzXsuBKSpSzZdISN3yDEgLEOjV6VmE/GzT07GHF2HAp+
wXMf2PEVvcu5mSKvPVeYrbBuMaabHyvmHFk0yQMUcLdd0mGmLA9HAXq4zZlEinEkWeKdElSJMJon
9eRuqxQ19L3IzKoRF0/9Yn979Vfl6gUBJ1E8OukfHTu4LQSFle/sczTYXSNk11IUMLvXkvWebHzg
mUjPATCrVH/SDq8h+DkgegiXrZo0Fu99Q535Fad0YF/+c1qdqMgZRorJvun0cWDwkZdJtyRGWgwo
vIHdnXgY6ajwwm2f4FuDvmJ0NtpWr4wWcIU6HhXoP2x6sGLzHkbS7eA7z0Ng33hdwITq3NCB9e7I
9ZduiREaSEuVbIrXXvdw0/OvrfQ/rWw8vMEwSNLhY/Ib1SiVSUW+NQ8rVCE5kGwz5Q+6+KMH944N
8TsmetNlVu18s/on7bWf8m29btqibIH6Ix3Kitf2qaCfFcf5AGqnvVtkMb5z2zPbsu8U7mEdJAj0
zdFWUGRAZ4ZOErbtfzpVF3ui5/iMv6Ujds1kAV3v/sPBbXh+ByBDIuocxQCK0PKNvCkRoVSSsSsK
vQZEYUpq62LqfCBNO/rVEenA+hgg5k7YGWW7fLQU+OQF6HhDxXSs5PmSlidePNUVreY8fJOvCWf5
g469D5ZOZyqq9bMV11v607CUuCFNhPUfO29V2d9DP9w58TtmBayuLAL54kVW574o8GjT2k+Iu1pO
dSvgt1Y6Wk70X+0pX4Mlwe6kjNm6ZuwsoeW8AizfRIYM5sElfnD4Fb3L8CK1n6aMyTyxSubhyKzo
3O772hkiZF6QwjgMIaz0o4O0JYYQsrCvUUjQhKcDlCfKwyisxGPw8+nZsNxT5u6ACcnjDYF7tYnO
TVwX2Vu4ljdbkP1PNtLxcgnUjfc9yORf0fao9lbtt1MO11kg+bsd6lQ/6CVASUkBc+uwNh8+H05o
eLMBolvDuwTB2uewXQbPw0vYfCWf8TlGPf5k3sX4+uKFM9wTTPsC4ZZ8KvOn8ak+hstgNOhVQr3x
Wh5XTMdSKWoRjfNxORvs5NC46mlsvINJbBe2k2zLbM8RAnuurKrY+FAf7NVQhJSLL2PyIDk/Jvpj
vFFOJrOB09cLJAhbBhv2KdaqrAJ09vGVTp3WJays2/A2eEyWtQz7bSZm1zOQH7ZeaqTx/ZbSXpOo
HrDxVQMdczdwk991vYMhe6vXJnqn2oeZfrZzjAk505McrVD7eoHtW07W2wIRc3XGEqDZjWDGVpXe
ARFgJqqGUG1pBAQ1Pmy7JMF42iQz1wqlLi/+bKInj0U932v65ywtuQfSUf4KmK0Ngi/U3SBhhdJo
1dOphJb9vjmqz/7m12Lsk48REvLBZHV/MzPlpDLs9GNVcSdTxjzh2OsA1w4QW+OTmKV69jNAZWD+
gVgyGnFQPODlXIhBFDHE70Yaa9znu8Y+rUZ8UOaG1YtoERKRITJlIs1HzAIyjpoeWZa1T3m15To7
K3psCAcTCFfqFjdC32AEEsIMHid8QNchvj+Qww8V26a+gug2Tj/Pv3qOWkrESeqtcqaOKH2XMksY
QSWo06HCUeDP7TElAdb1WIoqygBc8PP2A+lopiZrh2IpVO8FsXgAqvhJiSNlYs3GeuSVQ25vgXe6
mmXVlAxb5S2rfm2vLYZMuUT7DrjdkOUX6fytznEYCLXVzNz23gP8tdhAhJYpWKUJRtCPZbJoLPDs
/L7NzGwynI2Jm41+aw/+RmNgL36pBBVa4IzuUQk22nDIVJfGUV4oKg/eaEuYB4l7kLHBg5WC314Z
s84tyuf27ONoPVpm5mK/Kunxsq2LkSLMegOKAMckVVvmsjo5NehgjK+4ofbXspl8dQnrUe4VRCrA
0T1X6dVR4YBijEbSDv9nkcXz7d6wmB8B2dix+louBv99MtUQwcc0D6QBLBBET37RhQPgxnSeM0qN
GBfZJGUakBggMGe+WrXrMdJAKo+/XRrvTCZPqGrlYDTmodKPZQSj+Qh7ebaZHqArU3BXiPSFS22v
9HpOfIcy4djbyCR2ecyfZIwdFF3k4XLLbhCnMF94iZYflgVJdnZ3Bl+2DebFLTKnSa8bZzS7/TL1
BzYFmkphvX8ReazOHOkU0g5NB9mNxMP0zAWp2CtGIm04HY39WfeUUkn7U2VDFb8da9RNKnDA7gKz
eYH/G5PSL64It1inw7b8X9FLeMvm2BgTSZJjYE31Q5kEtmcSpAfWIE04KCiVcezI0hJhDjquivh2
1K1/XccRPtAFd41Qnz1UZFv2Zcra+izijGrWAYmhn0089J3XOhQxpLM1F6uUpToCfWlo3K2asL/z
X9A0q1tlGitVIV6p9Ms/nIjQNsU/snFcc7k6mOeFA8CiRYa9b9PjrAxgMXVDasjOn/dpdcK61b7+
B6kTqxOX1wxBgmCZBH+Xr0s3gmPCKAj6XrhMprv0qQftLR4RKhmC/pP5p8M4ZzdP/InmGchGzhCs
2dRakVL4yCb8AGHHf52jPxi8CY3f0OCAtHFMzK7jOft/zf5wQuBPKxpQODo+sljAXiCFs32DHT7f
GChVd3uZsf5YSC5ZQG+KHL1DXvXsdJdiu0pI32l5BG6HwCTPhT+wOPIi3EgJ6d7masyc7YNDjt51
2mdPEt1tUt5rNcCFLh7A+GKARo/9if4urLGFEd7jQK8zVXvZhjoHHWI88I/00AJF/TRd0u4EwrDy
3aaHJE2luqvPExWkvLjNk3o8OiAL8X8SHVxWbls9796PQKLZXtX7buvA4fPu4HmupASEokPCIGjz
D/2KzJY1n7R22idRxk7sn7nfQtU84Qgz/DMuM0ZxFABVihjpzgl1zxWP16bKEmgQTIdydptpZ5RU
3BQoi6toEq5hVc3434dJfaqcl9t1wWLC48A+YcehhHsJe6aynWCRLll97tAWBjMbj9xqBkfN+Bzd
Iyy8xqJePpJ7AstxheOlb+l3ff62dYv6fJBJ4KofAAhpL3/pPKoSlYIK+2oXKSSzJfYT2UscbZdJ
S+zBt/np0Ojcdvkcp1CQ0XHA5/kgkVLy65p0JwbvGDzW7XpS8H+SXNaVldkal5vk0rG/ObCWfoNs
wxy6in6zGIAGqS7onVeyHO9/+49UwVIe4A25ldVEwa0VczxnUpK8JLtDlPmdYPXlozKssyPjGz3q
lgaW+qIQdYdxU6/0NXhpiOaJztZMnld/DTx+Wq12lFOpp2uAQqKiQtiME1vYKpY0fbow8jUlVDVc
F8tp9lwe6ENm69MtSizWZaMxuUo9PeNKkc0JETMIymDqSzGM1JzFJh6cU8xrZGOyITbtGlNmfoa1
8/uxqdqhN86+8bMNU9sgdE67V9aarzDTubpPHhQSPju3rlhS8wWqkTsCIObRP1X/4t/MWF/hc3Ev
EuOv/7ajLvy2vN3GMiHlRFyYJk6hxxRLNA2gn2qZL+9FoYsbxXwcRzMCjl5qA2vjHaT/NMpNnaVS
NZRUZ/TSUjZRXkBXbWwm1tiZK3mcEi+KE2zG6coUlyYQF3HpiDZRZ6TcIk7GTdIxmjrXPWioKej7
78QbQLVE5NnldMn2OmXU4b7oilr11RvR5HpuE8ezQ6g9xQF+w4N7razN4V16UVuoh+3h3In1LMrE
iTyD2QoxQTINRpZrgeyvPUM122Hf9QJm7HvQOfB/3u8DmadgfqDLkWkDFKhUvdwTJAwlDQKNmyCp
HwdoPKb/Sv7yqH69AV4AyW1Ocl8luhPBvJqEFu1QhvDyZ04NiZiPJ31xKDgRYGeft+0JgWI4+gDv
E83QweC/IF06gd8uowvk032GMRC6xhkw/Nu6uJaoIMZH7KD4F8nPpvKctSMUmDbMGfM29hVhKXcX
w71CYdoafLy0IH7xZwQR6M+YVMG4oL6PE8qExS/7kSGk6QsWcnvUKWlD53g55JP5m8WtrGdgOVkY
w9PtGqG2y6kgdaGKk3MPwXoNKwE6EbKm0Hmh6+WiKjZMogEPp0hFIMXoK/4eO9PulrbqwJb1Xe4T
vhIkgcYAKmPiUKjk3WduD4q9mfdveXmWHWgNppwo4O0qFRDhq0vGXUdBPnJLeS0ni6AOLm74Gjb0
otxnJPmTDMYCugx+dnN4DcBOjSQefSTZdJ7vxzHo1+5PTE9Jo0lhFl5gLeJYJltA1DFugkSw+PXP
0WF02utsktIYMsspiF19BRmpJlfbFVc7HJlQqY+rqXRGw/U1jRctCSG5n3NmZTLHxOWWqYGa9wC6
UJ9MWbT13m91D4r4T+Nxh4RnX6BqLzusOQRybJoem4uZUd9uCqMgEplS9KJ9N9KasGPE5rWlKU3T
ENJWrHq/LqEmTSBA8Kkr1Ubtlfv5MjQjTGfcqGX9R1v/1ZF57UKC9YZZXeNOQmStHaRXfB6VsAZX
RTLVOZRqug6rGFBm9mNI3d7W+g5J5CMpi/z2DWQpaNzTP+SPQpuewVqX4RiM47Udke0U7fG5PHCI
y5DdLgj84cfWMRMRgN+Rp8anOcHtFNvT3Q4cZN383K3hytZU8kYiIMHVTsSdQi7c4D0IxG7Lz91a
5JhXj2cPPFMboQs2s+0vyWCM7h3DIEoTwOIeCh5Uq45/HkdefC7FbPXisKLFquRrF9rBpEONSayR
bD6Jw7u2UBxkF+T1+jZOof4SJ8gaZ5yEjOI3WAl1NiFofPdtIqYl0BGxzZPbFyskJDlnRDWgR4UE
dmEhdlKUVE7RvzxE8B2BrjzSoFZD7+aEpZu8my2rIRE0MTsZqdBU7wKiejPRQB/7ZMDz9V9OzXeD
DqmzJd9dtuU6KdjiTzcBM4hNSamnVBVT9taRD6XbUno2+5T6WPEykCUZ+XjzJU3oM/er76eaGw+t
NhZan7y1/GF4pUhgwAbIndaFPoUPgtQAXR2yAtDJsJHp0z9RDI4bEs+qZzbN/wZHNxx7Ry+ihJSt
Gito//FJioS+DnQurEGnf3Yvlxlu0bGUZ7xBa3sILcSsSxN541vbLAc++RAFfCJhltjomMp7Og4K
zwDkrwmbr9uhBO7zUPciXJa9FGse6T+xoofz9onMwcnEBvrKAsJT17cnYsT4SnR/LVckAOL+xPfN
O0vb4igV3CQtO/sbVTeWEwWDM5PCcCllmT92PcdnqIqyHtDG7HfZmxmxYW6uh7jK+5GmLL+cCEa7
11Iw5H+R6x4ukCYWmmU6rrpcjYvsSxbEQWtApN/tSlhdEvW1Sn+XhSmFa3tMco1kSMpTWRFbViGZ
wQiwjVeTiivXOQjSJsLknw6WpDyGFHluOc6ol2LmeSxruJBqFA2Hs3k6otYKahDQgaC2WYuAsCRh
i2J7OjSlsm9o9xAjB2rdOglHwjFQw0rncBschdCwXpa7Wgo6cncuRPP/CW6D/iHP6/7BSYo8BMMW
UEvmli2eDxHSTgdKAVH0dbMg9STIbvGci13JdSCIMnXVCJAb+Vbxap6/8+FTYHLcf1bXsuElGNJO
lFikSVmuE25ur4qYFbaN88VKx2q8uO3GE1K78xFYhsWOPN7qyirq47IpBpvFRmDaAHxN0+ZDsqtA
mAarhYujGILq/Lw9Y5wqwBhzGPA7JbGlC2M14Oruj1LyQzeLjJXsyuSPIJPAQb9JmMTbkO7xga8E
oAEMtBGT4aav0x+jLQlKShMWbMH9e8i5c4AFH8AO3eY5ZEZHO7tun4iGh0Lo5ZwIhd8ZJO05KeL8
cc3QikON/gf84Cqqik6jDle7Jf4SrB6EHsja80KmOTDVNZrw6Jircy7wCoJX0YOOc8UofVkYX+eF
J8thqVewgJtYy9/qZhF07RJ06D5m+OO7kuNkzYm2fMeRou3hfKcxZSVMdhf3pVHghwp5JTyU18J+
8GnlQ2K8ptV1vI/rHszEsxE2Max59sqTE8WcdPaY7JcoA3GzunxlrZlW1QcE6MEGSNUz8e9NyL5D
bI8FqN60uW9F51GNKU9nCt83Ggy+DnOb06WnbSCJ6+UicvYWbDbXjrFy6b9sTgMlvgMBYYM6T8C6
2bcmR9G9NmYLOzhCGXyXo7aqaMUgIsvxONScqkerqkaTx7AqLEFfx6Ug/CHvHQCMQEFI/ErxIOB4
YsB+W+k/hZan0hV1pig6avd/Za3en9TPOWppvu2eqqMopeD/TwO/LvZfT+EsQjMHNP/XYFb/x3yl
qPnbEfwFdhF/qwiN4lrssIxLBc4dojORtrG0KtoXhN+fa48sJZ1id0mWnvahTOrxFmbpYAoq6nV2
l6DpQ2cNEhVV6IokC+6BC3+lEUheDxOasOrNPA/01BeNVXTAqyleBgf0RVMK1hGe+6a2JqylEyPS
ql/eGbjDvJ7iW4D+Ic5wqThrRZsAWEldvmAwNNjGlR6Bf8y1iMrs+KaOe0nmyobyt0MPDMVtO9sQ
/DHeOVgyJEuWfga+Vt6s/kH5lTOSADHm5laMfzpnvvYEgGib8GJw8BIYNoTlp5VUJIAw9kST2nzr
VU8M3MDL7FOy7tVJX7yB4i8XppjelTuXlZe2yDk2vbPdcdD7XPtuEdmvrPG56amZJZgINOLaxOq7
5+B7Np+ZSUSQC/ddEyEM2kDrEGscR5hgfOrhdnd13V30JTvvzn5wmJLVErJAqM11pwavrOx69+dc
eG9tMu8KU1EWm1zZVeikFrxICUP1t85LFBbkY9JoBajDSQNoHU+DzCZvPAwQ2ZAe+/SmbUqTXzXD
OGDQNmk8E79ntDzW9BrXGGn7/h3DES+vWqFLCQqaUu2GtkHPojgcSgqSwxs79q1uX9Us2n0psIQM
OPfh5KSj4SWXuafLFqAuNPUzIyukfPtKhPrtRRqswkuq4eI8O2trZlwOWpCk3MfwkIe/88NKvoIL
be/KQbSBB2h6vENZRt1DTag7azD/h+FsQmQMBAzrrGuCrEMgFfP2Mfqqk6ew/Q2baBlD2dTJQr34
MEs/JbJQdecz+7BkEAyWyNRsKChgTZYOTTfZ9JAgAznne935pXRBLkaKiRsPH0eekOMQVX0Bb9Fv
L836nHM/vF6n1v9UBKUSGDW693VXGCfL2fOf0F1X58IQsqhADp53aIckWj+auNh0dpMwYoBgkUD3
azlnL7SgmLNj+QBsYGpwAABDyDz7Bq5dGO7XuFJRum0686sNbymu7a5/CizZ1Ui9dHQpvjFt2tPI
zUxC+EYcMfS2SppUse79REOJ/j/mspMZw8btaBcEi3IhfKLXXMbdor+pa4a8ElLkL+x7FLfZSSRv
zCvUI/yJeMXZaSfGeODY/WReU5hR1IK97MUzOAJrcYNkmfjaf+SL3Ml2hwqAZTz5oSXKYDzbimZw
joy913zuVJ6GTzl/pDSnI/jWl7++BEhbykJ965UcUWzJuE6s+OqN2PmAM6uhCtvVMXkIfBfFU0+t
NLFBT4tUlnGsdKCXu3g4v2uI40FLKZBb95r1q8CkHWZPSmSxEEk4qie8WWO8PipYrlGm3182HCjU
Vt/OanV3UcgObBLpVFYtzZ5e1hqNNJIgTam5lrQVmoxnttUepkEN/X1l9aC2xshZ/l3VrSwFJj7F
A2xlYPGENHcGpLduwSWUszkY2hORG2lKoplA6klBUqCSU97OPTBQKS80L8kk2Wo9L72HC5Flx2w8
q8NnTOrBqkLAzl/PIqtdiR5L+HAu4kiuh0TmEb8FUbLNTlMPA6pLefDI0Fg6xPoj/rklV0octOFo
Cy9mmyDw5rLbmryonjhJXa/v3v645PJp9OHsB+dsW4wh1CkX4dmSa8a6fUl8imsQ4tvBJi6RFxwl
zIUW/1FgEAZ+l3aaWEd7b7xEbhNzWV3YN41RJT7sd6oSHg64L9qfcunIDrDv/h+XgI6IzJHWI9em
qfaQMXYduOu6yE4PMB9+j02aYKrWjX3DrCBPFFh8+lwCE2SWpi8TQMihd7uEz0SeokiM/ByDLJ0T
QxZetnUDSUav+KtEm50joj0lwgjtkioLb92C79FRKg6Ha1s6a/hcRH+41GIlr636YLQiogiYcTci
kgvnPHvBZjvQg1UYQxeWH6+aG1h7mzKVIBqPUPbCCoP530jGuGeXqwu0x2uBdRpwsZ9XYN8crPq4
PMCu7qo1+2a1Na7pegvXjYcpKCRAwIPWWO1CPpuj5xs+wRTR6pG7KNsF0YBKLCfNuq8EAijXnjXS
yLyeWshdlFFEKooy2D6InWY3C9FAEv43kjr+2J7F3R0kPFfGx+iXFnoVrBU7GvIKQ+jd4WVaLo3W
6A3x9FOKjRtSUxFP78PaJq2B47+Muw6L13Mnv9XkL3SQlboYmxF3TWZBZhTYG8tx0ntVLCkFZImi
e7HuiZb5C8PIIn8v6dRx/4uKnGhFbwLjYsZp5Qe7ld9uwPx2NIft+KKh8oCLR98a6nmbHouDkO8W
RcTQ02ENp+fXCVI6y4yApqMTn1oDvFyWQxtSx5BFC811t4aa1g7sVBibNFx4kl6eyeBo+IoV8J0A
AVqBdRri+rWTjN5cJ49U/sfKssZqC10Lm95Gh3XrwZcQGZqHJ/FpzlwXHf0yokeA49zbDcbCSYaK
/481xEUeOQSgsJHKL9b0Hbp0KxuIcPS1Up/N3Wsoy6SNcl0zK4Gubb/exGr5W++dupiYdX1jgxbR
mIniqz4qeegj32T0lx4ESHBOGpdQP56VGuKaMY8KiCgj3i5CupQoZP2omXi1h+oF4v+EzxLGshcH
Qn5lrrbPMEH6IEJ9pfuD3gmHuRrMWO5Zv9wFvI/Tw2T8bMn+hYm76uY7hxq0T0fPHNMrk2+jszDC
klotHPMXmRfX3DfZQJnfZCII45qcy0M5LvUu9aHmJoQ5gEt2gLtd3odeZLib2szKCoxC1is1FQMC
w3dPkVftwvr3kPWE4TmuB2p6aru3GP8gL/C4xSX2iATbDiiyBDkFh9demwbRwjmM4wUP4gmLN9mq
cEYVBwxMbK20o4maCNubPeADkA+290guMlbFMgspvP7nkOKwy70Lgbi2DrmY4rl/BWPvFCAql7y/
xUuKskc22XSlDed8f9yAe7L6SeoPiLDPT1+20DP3ufUi0tDK3Y7penSlR8RtTSo0Yvg0gM3w4pc5
qSF53I11uZ9RfZFkyTNqLhApyr0/eUKHuGRhU69wz4xBJ1QlmhelokLbtJsmpipVGWIdmbpTkG9c
B6R9t2TPH+tOSnNPaG9vM1Qq71Tbv8ZVVyZO79p+ZigOD+YBFg3gXsJGe4nPuIGOt9MvnJ10+iEM
xxhL5ueRVyh0KxblS79j966X2qPhLfvVLTOgL3upEOcrdDiRoyRQWGeRaEFuL0lxIYIrT/8/wsin
r2GabaBXtCKtbUt2tQZ5BVsMgUb+V14Bi8Nnn5RjgYWJDh2k+mzA1q1JpTf5UHaOapxuxbc7YoY2
FJeDITt/fs8f+EGLqI+gQcwNpseHjxyHzyLpq8JdV/wG0OV3noORjBrPQlHFIVsUB96XLeB5TXjO
xPtxgDul51CoXmEV9DcgellN2YuRrBpI1JhtFx75bEI18LnBWAMhRn4KYZkHQ1dfbHjO+HjSkkEV
lh8DwBs5YP7LpRjeht5k/inLLj+DPrlBdvouXzuTZgW1JRbnHC2xbm8hm+6Ks71m53HsUMxb9lZ4
9LrE0U9xTb9F1CEwO9a7DC5yqVF8cfYaQVLL2/UfiiNyeA1WeIv2vncPHbky6l59j5RizJleGgSm
pygo2NQ2i5T4kWHYlzywds1HQXE1oxnXCCsf24IJ5NdbuQdl8PQp5q38FHjmHQ6P8Y6ci4bhCfGy
jRr0pqDH4x2AFJ70hSvi/SvTknDwvOtRy8HNl5osRwbpPQvcjWzOAKZzAwhtCUwDskl7QSua3NuX
OLr3SMfbb7UPBmzzl52N3Y7QtzpU4BCufoxnP72kfOs2XMYDqQ3uvoleOCNwodcJmjemGeHwjLX7
5hc/bBIPXmAOsNOy7cVnYi0BlkKMkXyMSYYBGc31mI6Go7KeE7tpyhuxgFAR5YnptqObcXbNhMMx
FHJz+lRhFjLKWByYYT1kE6qRS+cu9b1T+7K9x/wA9DxektNLA7a//f3728juiDz/bH9EU7X7fmxc
5ygpGmgQtPPk1Htek8PFUR0OU0tHLdRCEqmik2YA0xQ+0uyJNo5oCpMceB0JwHlrK3xTyJVWZAwr
d4HTJVKMHMGNO790UFfoSUKvRqafZVf3ou5+YOARWvnSaV52U3CcEjgc9s0y7LTdKL6u7ZWzpC2I
lP+Id9XWEtV4XzEv05u+etZeyQLfOR2UoVl0OE/u7Ic8GlflFjj1WJnEW/X7PUFuWiEnSlAlF704
vUrmhZWXJosY7Bfss5nfDd/vRP20Ji7OGcHtD8wbvyopNmCw60MSrOq46D+zj2zL1iPl7BdboluJ
bqsIWMcs3B42HBcXJ9FclO/PfObWReNJ0Iu+Jdfbm3OISQ1QBQKpNoEJ+3CCFzhd9dk+c+lNSrSp
Yr2PGvk/UJ0HI24SOB6eVtNTTu4lyB0j1HKYBcpu3pfisZRU+kS9ecJI7la1hk31zGEF2QUntrO7
6wOn9toaI9CQFFPLyz380LQTqfGnRb8xobF0wNvvg+eO1Xp+K+kvohIZnI/xS/wfIKEHqVHEhZdG
5gQm0toU6iKNlxJcsDIEPpT9l84fFZSRIwZLnOoOT5jfOQEXPOVUWA+rD5MQ1uG9VWnVOY0HqBZL
J5BP/cPFl2XvhabAzvKOPahN8uca8gZB72/q7g31Izz572SRW5XeyQ4IM0aFkRrh0pCF1U50i702
UXHcb6O+kByHXXlv7dmnV0wvWnxTpFPUVBpDSllETQxzncPaH1cVc8y0dHU90nLsw+f1PyOGPKZ6
8M9bnmsJlIRm04RuxmIc22wqAdr+etRg0VM+nIeMGjbcavDQs6m/RxFTrJi+68/lbV0lTSP/2TOi
Q4DP9A867+Z5b3evJpxKQrEBa7k83rNPZvCypW0YbFK/2jqWnNMOImGHW4J8Z65PF1hMPZdVa29Z
LNZ8O/NKbJTBNE8WLnW6YB4yNuuckJywbSkKl7B2n572/F0zzKx0jdMpJX3cTtaDGrew3THMtsTQ
S5YlgDw4YXZn/PqBcE1TKty8ZoNpk2t2+iS3zeipDiYPeAEo5HFWmb0L2tHYK26TLiSCBaTluy3C
HHNRZCMkdqzTvWnjBvpisMl58UxLsBfBdhZWPzia9VmjkkhbztFCDMYeMbiAeBuWXjF86GQZmhNa
Esk5CwyFgJ+RL6kV8ASkp/Dfnl9FwV5CqJr0gV3X9/ym4PY8TxHSfuR048e5qD9xNPMc9gwEferY
iAkTEcPBoTvSal5JKz2yXaJnfOg8nxpf4IWjDFnqbtruS/7Lfn0QKbOoZw4hBJEJoNdiQFom/9xe
/mZe0DLq2slF9bsET6WiYuN568J1GgcRN/mDci2r/jQ4kO1DMpZEVAWnuuwZiUqyclsxpwnbDEMO
0EJxgwrrB0VtDITH+pXt61wKs6rz52jnWIutLWuIdCMj51RtRBYw8Qqc/Wry8LD2vZIH8yz7Qpoc
sMFpQTkWxkqL03e+CNJZ8Q8yKUuC0+3osswv03h/skLM8JQX9GNlQZZNT4arsBCCuXaGcuiI8RpR
mtQWqC1nZVn02UbzCxcgVeL48edpOLWsYjJBEBL4pCxDIMR30FTuX1fTJwBa1LgaJpN4R3xx/Qmp
maQN5CBXILXpB/WLfFSvxkA3QIVUqrhBZ8e9rtEmN+8tm8zXEitlQRjDvsajQAz1ZfTwhB9mVlPK
VtkFqgZc9UI/u+oAbtKkssS1KUudoLIs1sfLHb2VACaNug5UduEs7Y5X2ANL3gmL3LkIXOeg82i6
uGeCGwSMzMYfELg4zuarpTxPAa6/vAnY2xD4FiqvdZm/nG6p6awqEgYnJfYpviaOjfEcM7y1A4me
R2Uccot65Ij5ivCuVT7P6b66P5QmanBNhJz/lIlB+hHAoGlUmyMdzluYsl5OUAWwofT64CdeqSWH
0KzOEdY39HbeJxyxkTi/jjBkrwGHIOMi6mlfwBPM0icOVhP9XmHxlMdZ3VzASi5PdXWedcJyIJpY
JWsLLzDnAGC3Q7RR32bcHHqMUK3DNt38Lm4xEmkWCUCP8qOeJXZYpPogGM6rE1vB+19ROzy6t1wa
ExbK1gKi8p2i7OgD32x6GHtz75Ba77Fnh3zX66KoxJlToYlrdXBGS/rGh4BXMdWIl7haYj9bvg6G
fvIneAhFzwjRXgH25OCJMuN6Jkz7mbe964triIPHHACkKh8mMl4ozoQlnuSeccvpz+8O8pN0zHxb
U67VJaDMA+VV0YHl7b0zaAjgSsQ+9XTQvfjh+VaXrGHxAuUD2rDBh618kmHlyuiKcuRSM5l1njd+
dfcNVFWR/sTPkObSyNBsco3zHIHSI2G3Rww9gTLBTOwtmLbnfJCBoDxvfl6O0Uq9xOogG1Aw2Z9v
HnArsyG7rZo6mbJ3CCdYVbL2fXsIihPHzF62q90Fgsuw1EQrGhWoM2x9qngK71ya0I1rhDgUyyYw
r6rwoC+UxWNGqhLbIGY6O0jMUqtaVVYAi52TskZg1NQKcz/523+GDh1gS+blW0mSMd3S12lk56LJ
906iJmTG3BRUHz6UAaZnS6YYBEvnCb3+ZG4SU9VngrhNDKBLoju0OnpGR+kVu3lh/bJ1CK3W6D+E
Wd7Iv7CRio1vvW7SvAyHCTrtNFY+eTfI2PB6Ra56j7X9yMhxIZD0U9agQkSZ0inON6a4xe8ghDRy
1MoJws1HJ/dKWbKdifSP6cRq0TvC9Jvu1lTGKVCEeAvUUsFvZR1w+GaltAImtyiUQ7l9FX12Nirt
e7AhwadFxXnO2MxXxdHOsKScGbjtDUG0vIz9PYf5aXN0m68ABmmjuxA5Y9iwfuB6b3TuHGX8Z2wz
7dbcbdoTtiHySSaspiLwedympUPZK5MdvR5O/k9pI1o8yXnpeXoUhc0/2QpKns2sf8ewMqQ84mqt
62GExZuCibUCXhmef4GHsW8vO/5u96+3asvHUBLhr1+N09EJ86wEkieT36YeF2dzOtcVeCImR4sm
I1XLr6q83E22YWTinqYQqV8G0fJU1Xj46xCtbfNXOdNyCg4hTalxngaXhuKoYUx6BMU/RgEqE5O8
OmJf0fvXE2YmiIlmcekeZK1c0ttrFwaldEJ/lcBzkHhvZBzgy80oB5ALsB8hv3a9klDv4HoqRUUy
ZC/20udSvyDpPQ+FrvZGk68rrhAgLlVPyq/108s8QpobupDMSneUPMX9bd/cTIDI2g9ii30xM43T
efcGenNAL5veyaYewdM1IKbT+Wv1V7vkvVKVaOIptx2n8Ri5MhKK7ddzFftwHwA/YSvlwA/xBrO4
mtHqLoh21SlV1ME61wtkeDhEO4OExgqTHbYkqXOtcjkpM3C9jzG4YaYKW0az0ywRAJbQ+nXtag6B
8Jl4EBxfpvxfMI/4d4Zd/GHdW+69PP/hDwTpiWUGL2i0/t/5Kl0SfODZQIwLwn2jIH725R5lKSYD
ysgU2jKdrfhC7uDAPuxQG+GAVc/TNpC+JQRXsxRYrJ+QzWwr9dwx5qHNKgbyxj40jH0ZXZEtzL5r
4C27d1UkCEUv68DcWMEmvvC0ke3gYkGKi0MHZDVmX9m9pdoQko2+TCjlycNqlNrKw85tbAbRZXRx
WXKs4y/DsHRtvZYFg5ZP3qN7tB7vtcwdke2TIdyW96rEn28S3j/lrjEb3Smr3jrJKzwJ2IoT23cV
HGuIaYHTIFoxZKAOUGnkbkMnzz4X0nXQFzes1zzb1QZnsUO31d9aI143AuY7YEHwx+zjxnprsEAz
LhFgFnZHPiUlUJ9w74fMdVwBlUbX56WieZT8yTwvrg90GgN4ZmcYxsgbz3KAHcLmRWdbBzfbnA8N
5iLbGNTLy3l5IQI6W8oqe2a+P6MO+Zg6ta8shxY0GndpN/d4v15K324gG50TD+QVMCRuquDaucP9
c9fZJ4BMF6HlsNHQ1pJZ+mi6SxRAc0a88RV1fuRUMi0gxXNGEXHXOQNFvbgzLgEsGp2YiTeO5Fuk
NYLFtK/m+GkE8Vq7VFXKyYT/2VwLdD34aIag0QBApuNRWLH0ZMJZHUD57kmwUvwJTQgp+4AfNGQA
br9PDLavQwwm/dEYYfQ+I0BA6CMqerOsT/VlGlAXCpFOac37f+cT2QheS4YKF/T9Av5U0FkWYYlf
8qEhNE92eqF2FufwG8igoa8XcVtStGdyBcHUBTpHbIZUZmnMV2YLKc0mkIMIPtWsWgelK1o1VvTT
snM7nGCNRwj5xDREe2J2V8qvqGXTZ0hXL4N+BqKawPxVWS9tsNE45FoDGIXSKu6hdRkD9o++I6cG
10us1RnGFFrzy0ChDtC7wDIdH4McWX7hxHIPFBSS6ifs/G+YQdp9I7K9JUj7YsLz+7uJbN/FO+S6
tHx8Rfi+PpZEraYF7F5OyIy6YO9qG3Y21945gw/w2KMZlJDlIcXLQojwt1NtUll/IwjuGu7XpdvA
tH7ymE/ok9lzhgl9ezDxBwqbhGqcm+MZ4puxqcAXQ0FsmfYZLDaPqESjy7IbqTFJJDgoizJtBcMv
BzZyscB0Y37n8gXsboZV2OdWOqJKR5g0bD4A+1Exs7m0Blqpo2EIoeZo9WcGqFnGbizRd1Dp92sC
zaRA97WiGU1viUPUZ5UiVG7slpxm/GYvN5pw1APcCaLjQbeAoX7+ZLwNp7Xn/hprgkKeY7gvQIY5
xTo9wPa03jmcPhxJEpiM/1phUPz2t9500DQaT+b8U3lG04RKfMsSwBGEuBuHAQ7p1fiKwAZepl6d
QBlGLYnnOkmunvvIk/yYl8cuF3EmrxXaG52JN+gzJ08xCWOJpENi62JskEHq7OLm+HywAIuL//B3
Wt+eSFAM/5uDU0Ux16utWZv8Z7PHFxXn2wo6tvCzEp2+xg/S3BbvBUfepfpWrK9QcXBs5uIAxRan
vppPpYw4i0HJ5d8CAfW13LbuXHtDNsfnodPmM9Hql5kPypxkVTr8erlGxc1Xoea6EztqZWVYBbBi
WGKL+2BKVEG+CvneHRJQvUwd/iyXOLK9V/8aAW/d3JdR/RKcwD3EzfY+28i5A1ZOhtf75iNY6hOP
Uhm2FAUl6hxr6y5MmDArnTGSnW4A0aCuA80Z8hl8P2A9u9Vs3y5U+7O+rlrCTtusla1Mv3TnzfQU
YvsC1UKB6NVnuMhPBBqnnShzSWqec3Pvl1KnMzT5Fbdy4gapuno0z3ysk+aSGtbwIHFx2OO7Fw7Q
2R3RczEP0tA4SPLCj0kAS58gcKVAeyXa6mqTZWHGMj/saVYkRngfX4rGhkKGZEcX/vgKkJu42p/N
olWyj/q9AOdE7xUwh4H/+FD4Zy3fx2yAlo1EeG1fGUxbYamhA2KQ2Nr4m2WP9XItQT9U0c/DRJcm
BfWahkuRAtsWkPbkbiit9tLSNcObHFpSo10XgCPUiAp2wWnlWZAR7KqY36ludlvWCbarsTSdKuSk
Pq27nRUAih8bi83QK35Vfdc4bsw69tGhtTFOH+UE8mo+JmR4eCBjWXnzU9vnCGeqDFGhHPekMY1F
B7LF9cVGdwLBFNyjAE8GWr7zNxZ/gwHB8E5A1OubnvvqgvVjQzcREUo7t2qq0W2u54/X/mz95SWi
zNNJ6zcschq4LOHE+iHPEO0LvLKlKQY5TqBEOHUM5c6IIJnJhpD5h2him2ky3J+t7ieKeOjA/JEP
MZWgI6G1wDjDuHNujelk/7kxJsCapRne9gg47w+7IqNN3BLC5C7EzQ2FUKQwcGtwTYaENIW2HS+T
ERvsWi7FUL9jmxiPLC77NwBNEz6Ga6FWkWrWCPloLCdWMSYu1HMMglXKTIp2uvIttlJ1Ce0yJNJ9
gDacdHteE0fxOyolJK5J34T6WHVhgHsYyoUUIBS13rRYVOoriS2vyuqpHFFh7wIXatk3O4+OTuzr
G4tuwOs8zRp0yf4Lt8oNlwxBmO8hodvdhixZmV0Xf/govKpyRXU3qx/tkBot4Qgl8eibjuABGikq
uUgwUSaLSC8NUcnxcRUQ3eROUHUy95yuBvOEy36q6Xsyzbes131uyNl3ViPfIec0C9x5BmSFCaNE
Ff0VH0nW0cernI2XHAmObqQsvhs+n5K8bTfNA78vRs9XDrDtBz/1694wuMGzZlmj2jEJ2ni4q1EH
fZIRQcBsQnKnFTGWJ0nHWs8e3wCuJWoF6f72Ry1HKpsc7oXUqkCQZGjL3r3+4XGfC+FC5gvSri01
4L2uSB2Mi764Ep+QJAfBN4LQmEz8bWOVDfF7A1rzqDcUzvW6KWxUNj/NNiOXKFimP5uSBro8YoeO
GQkwHYugsC6JRQkgn3BYh43314aQvRmXgmtkR0VQLcvhmv6ArLvUvMf/p3N6t8W/9QXmG9TbIP9X
G8Xxg2Ksh+L2HFcu5TITmcMHjuW3D+OCuh2ost31QXK5dEQ0NbF8clACljfzHFJues6D4bJ+rSaJ
8cY+Z8L+2oT3QSH3HdPg42AeIneR0xl0gpK2oDklB2mw5kLFfC0pQdjQjFZ79YJDfs7k0iVZhmKW
jc3+4ETtCMYXKUwfjvJmVmDGuYRrc2vDxIIhlk/IJW2LkhGZg5HI6RWcHO5/6anbctr6QdMNDI0F
I7hdh2YbfXzGJY08XYMOZicJdnVH9F/EBM2rikGEowzRsra0axMTs7nDA0AUfvmfrY6cFaQFh2PN
qE/EtfpyCAT5Jw/ZmvWxN4xa1WRAuQgNB6cO7OFnqShDKkuVOFZek/4dmO1IC34PT5CaWk0DIoye
3vLStvVj1pEkT/ZU2gffVccLldOGakQ/XIDqXkLsLS4BotQ2eNHI/9HuyTO93eYWalWQQ3a9+im/
YyvI4NwdzeS2McvJ4bdThlQx8ldmi8pgBHlJKaAQHXww/ElvbntWI6mpAtTvaObY/IP9f4eGOOMY
sPFM9Lr0D2/yXE3/QPgP/cfVY8+q02BudCFsLxxxAcaKyET+Dy7JhQvY11w27rfobe+zVF0Q379d
icysJvvmL7kvGtkmybHOGevSTnfze4s+8Pomyk2WebF9WbjVmnISae9UvMdKjefK2Is5PEwNL/1d
/Y6coJg4GGpS5rdzClZH4PQ5gvHvxqJQDsysb1yeyU4/H1gpUsnbyHun9NU9KfLr7/laCSAEu+Ax
nekTrA15PMnLJ2ucPJUbpsnaIkTxnjJTmtGZlx8hlx50IWXBl5CQ0+kyeCj4t7xlpiNvaftXtDCf
7iTqhJwGniFyEppxbDmOR8O/7pz3ZKXK4NCbgma3hH6OaIECs8ejkpfmk2ndLpeuIj3WqVFjZVY/
RY3jnI3uqqS0O1neYHuQcj3PGLZV2KpZvjRouuivVNOprxu42vVsKDZi53HJrXNIon5JjqIf8C94
zaqKqtc8A+yI5RvaufScj3VnYF5Y5NMjRJGBr49IO5F9KpV817RUOG0myXWDh/BrCNT4jxXE4Gno
IhwAvzQXSmdyIMGsIkTLaLTO7bwU1RVTlTd7Riv59hG1X0IP09S8FOD1PKyWmRgWC22DdhulXE9P
fkq2rycchtM+hSmEzsXqjX7jDRB3JEOzx/naSydunvRfsETN5YQBcQzJ1wLn+5v39pOXWCceQWdq
yWt40uVxzcg6pdeXs2AP+l97w353HR/HamTzE5v8enc9kVMoLiCtvXiqky04yPFSD0wf5J0ChwH8
rJ5IhJlqrKf8eXlEoKJS1iKR4QUNWTg5/YT+EGjc3AvQ79D2Nx6Nfqjf+O57LDSS81cxVTuNXdPF
EwAa4vGS5SwP6Yeea7sUeRzWymNE4Z1R6Pm1u21JyxyvJ5OUbwsHTGvlG+q946pnYC7eBFqQRLCI
ZSzc4ErjaR9EfoPUiSUigf64ZSNOotowX+va0teLBVOS0bTnQeowhmhgwm4luRfciI31807yw+MP
GhpHfnLhU6Ri/iWBoThAeQfF3J1aOfEt3NbLyprsmL3KCYQlLQUZf50gIlewggaZF+Vvlh8nZwXA
gaUQN+yks4nzSqIdc8GNIm4cnJjofKWBMrkcs880YPgMYzwpj2b/gWdx0SnqATTEwhtRT2r1Qq7v
AUFEs1X/vELkyILCwWbxw4I9IYMiVTaq4qeQJY3YTIHQTZtfPdtSY+YJ6Y1sU7+YrgJnupaItYo+
GEdCOYZWfzDZFM040Herr2GNK0/CJmRHrxKkbtz4FdhSVosQOJttFMttfWf3yijDc7lZ6dxcXhDm
YByv6Hnqg9s8cJg0nbH266ArzUh+ifJo6jDYDIRWOkJZ23vBpXX98hCvEaFY4tJpGgnIpjXSkYG+
L3XxPO8T9YCdLo+AfJJpSbMLJPhiEeVE4zxwwEOCGL0D961Lu52CbFyTTpD+NFM3U2tf259vPDyy
vvlOaeJOj+vfaObaetrpCNmCAaweeEmdsfni2dT+HEP0tyCdqVWn9F9lsw9yDaVj15vTWemUrVr8
QtBdoe6ImjQS3u5wSQ6dB6BA/lhTsxXVm6XCxOACACHfAHfi+3c42GJPaWMQ58PtOJ3xMdF4tagP
buqlcvNg/LIyrULYxwj1zabiRtTT2vtgq97dLROKmzObvLEZLoKaZcU9nZU/j+7yuAMwj6jBdECE
yinsXwCq0UdokwAYHIy8Xj2+Wza1O/J4ex8SZVW21zC2wkGgRVwav/88PIXw+Vq8OoI3KWIl2PaX
Cv7/3FNVWzM+BJ6pyYsqLTvBC7FN8CUpW/B9uaJVKDKTCBjBijatJH33yy0lIcwIPTWlfN7gq+eO
XbSWyQdyL+f0XHucXaNINR9vneTt8IF8pQEBeBKzOuDK+FxD+YaTtXI5tA6csqAeuYJrcVA59CYO
lr9Aih1W+6ZXApD9OCP+UD/1qdhDdx3HdGhMYLuu6rC3t0SOAaZs3d88X+oZtIfvOx2RvvvAomis
UtgjaLC1TMDxONYLZOKNTPP2LUhhORXb1lNgaRiZ9Nct/Nerb/Pjcj62TCES5yiN96TJQ3sa0x9/
VF0ja9zhZSQf0yoiq0yPNYfquKP6MHEJUmo/4xxZMwTa1C19gmTzhp0MYrG5YlJmwiXlGyVMEuja
Qv1xRHllNyWCw2EaY4jWv7P1bzFmelbm9U1eFoNlkGgBRIvXBnFHWw5z1U2q8wdq56tf60JlC6PJ
sLkFwscKl0HyuNchRu6/c5Rn5/ePVEg/dmwg+hjGPYhlBf9nK6nuq6UglEAVG1EbAmo68UzdMqLN
0pWSszZ+ZtigYmQFqoM3Wr/R36Bxp42MnGng8jZ5H4Njr4QpIE7idiKG1TZyE8F7qJL+WRiDe9sC
dGeGZvwq35JTz+sFjgcDZ+XaWKyo5kXlqTUDF+2p60MkDPUqfY8xiiaBO7bc+bD4Bjl9AK06wRgK
ja+k9R9gaFMXLdKYBY+sP8jbTz5RTeraqI9lpVJZnTHq0LI3K65502B/u+9h6++7ub45I9Jq8ID2
qQh0JysBpCnb3E4HVGz9wps2CeCH/qpyXiT9WyRky8SKI8vV58O0pzyRl4x2bPs7pUOJFk5XbADX
GBGmeMLbJrGq4gcsAZwpfJpG7PdEaw5rtz8L5+x54Q7xwIyVuLpH5s8rCAMFY44qGfIJ4T4MysTX
AI8zq06Lg9/rZrxXJW0EcEt+PMwNa0rt2aA2WSjkA/yfqkWzjB3H+/9MXEF2/FnSJLLWC0dL7hnq
LfavaGcImpihAsWE9ElgtudW92MbK0OYjmC6usIvV8wkKpnFi95VDkI025wHYN/thffBXp8buj52
/Tq9+DRH7r7iHtaHbVMaen2kmSpu+hBvHdahdBoS5PlP7t+qBjd6iL4gNiOI1W0CFJOG2MG48SA1
WfV40/46NTQC97ga9hPSmqOsOO0KEBZ3KbYkX8rMY3chrG1u2lKspb0iMQNCjgdp+o9xYZlue6Wg
lMgumop4cQxY3xTnEDynoI9yllEI78DoI1JoF6UVAEbJeUl22Xb+rpkc7RiIUdqIJuIxsZkqcH/x
40KB6hSNIgZAyijMjUKMdb1w/vNURMGO0eSmB1NaGKuWqBE5PmYKNk1W5RFhfOuI7lYtPLu924vD
A3YA4QPKisUsLTRvf3HQBr+TlGVDZvKCc5fReMeaCMWgrfDNynBJjwRKax3rZRUq3tGNP1PT6lNG
4VfuRj8Pc3mEbvgN5HJAF4TisRcMJAlNaLuUb01Oyh+2vR5CPTebbj54cSjYMda33m9mYxMToZYQ
MJH9omfNYuw5YiUL/HNfaVnm0j3ZfaC9z07tEJMwVWws3sJIKgjHBjpTJUJzq0hsMC1vBT5Hjrc5
EylD9x+ONvZPeVgislwd5A23kqwdbWrMo16gKlj9dwp3kXfhpcNLV1GRMmBpmlqX7m43wABd7pj/
EtfonfsPQBs2z9QVMQL1DsYvuR3geR/tWxeVxEPfugEbWfarKiu7WgCEFfxB5nx3LbKXyFg9uVm8
tSGJWEnlvy+AJkFsAGhEPST2K7Fdg42doqckvZHS7A9JyHMIX2lIn0TJqQwMHBjGI47StoE0zT6B
n1lpIZToV9KWdzS0S36TadNj7EbMfVbRFl9T2a4vWWDd5uQazq3fNidcVGKhOiGcm5EZnBf21y/i
XTDAz9J8aodXpioPTZ7/wswb37+s0E3f46zhBgdSZPagJmFnCnE3Rm3bq3INaHja8ObHI/QokYj/
MGJ/m4sNhezotpEOXH1lwY760OHdEzeKCmxbfxRgxDU3Bho5/Vo1r2ffR1kLYEOKV7KqaO3/Sh6i
25AkFjR51vCaSxPExyP+dHJ+PKyt3SeezsMs9jTC5DLPCS8tepY8y3h093NSMPhjWJzh0UP61bho
6rzuGbtBqPa8aZhqmoJAYq9ApYV2v+EKAkMUqAqUtp22wlPKLnbByg/PxHLEVuvFIHk9L83D7HKD
MbW4dsQ1nNyZwMRLdOJJ7BC3B/BS2gWsKiCseZ7edHw5KfoRyuCObVlgdxrhL4DE3Kl9XmkZ0TXG
9T3UOgYVH0fpm9nn9NPpvj/FrJcYVlOMPIuumOCeRpsNFJ8zdvfJ+x9ZQaPtzuRRFMSxhS8OLiet
Q9uib8JUhbkEYD6QndV5bu7aGtggKI3DPeGX1I1Rkix81TzZW5CjtsNmjpWm1NKk9aOoyD3iqexN
XuzFAV6+q/ztvzhVbloJzaOKz+woVWAbXzFnB8p9yCrLtr/FkZpHEI8B9Cs9G/SMEx7fSRdIhMwl
O1Aicv2TqlwkilltkasgZnb+0U4h+dkrfYdIyNYNsS9I9mwgSj+7l5kZTXGyhiR4iW6kkFSvomWt
1BJApLj13kVDQo8jtUzioO4k5NsiRC9bwOrfdZY07vX73n9ZtOC8t6JLisRUeTgiKLSPgOQ3NG3F
iU9bHSFZq5WZP0Wk9UJLT9aKuksLT6ZV+bh+up5K3GLdhVKj36jtQoxwwtxucbgpY5p58xgH3iid
hlFuivqkInFiU9DdRd0ID9EWBr18KFz37MAOO3dzwkAHkf8YqBffSFkdEVgJPH5DbOCfyyqJVJwq
jG1zPv2HZx0oDS/wU8qP6QawKRX16feHGYMxHGDFvqC4fArjDjClfpRL37sO3oHYxkF7CnoLh0Gg
nVg+2b86Qfj8ugvJQdIMdedNnunJhPRFm72v9CbQPlF24idwTkHjk49ioaKBIlcHELaDqP3kWJ3w
SGNUPRdj9VsDM5l3SP2jxQCXVPHpSmSdVwjb7/yWBivlXGAmqi9XCoS+cxdIvLEN/QiiWbgXIc2z
aHO6Dki96aRSS1KBKdFQcTWGVZ2r4NY3KFkzeshYdJbJ1/6KT7QOvyam/BTmVn3w1wyqKEWyFWr+
a37h+4ti0/Qupd82a5lOIWSW0Qd6A+nFUG9nR7k/vdh4f/me7CckPb3f+hpSC97pNcU63Ae9bwns
z8cMjvqmhW9MvYwQ47h/tQj1gUri7CpR7h3HFaAMVPzizlXdUdfaImhqlQSiLvnkrWZVyNc++VaZ
7e22ilW0eeNcdNZEP91wte3YgHM11rRi7sApmMf+bDcH0qhx4qzEKmAhG/9QfrM3d4iZt01UP+vw
dXnrSJq/G8UY7U+OJOwWdeol4sgngoHIkv7qZRgQpvUeRS+0YCB04DFDPmf9Rbp4KPtM1Q24mzQd
aoVWmX4UXRLMr/u6O/focyax0RDAqG1HbFrMzvhgSaku+c4ze1fCLOGyu31D2Z/Cm+LcktukWrAn
sd/npk6e6xcVKdSxdeYB5FkJcCzzzzSGXFLX5srgnyb9Y1ZVV+xvtp4WH+xIP6EMswxoSoiSkRsN
/Cw42n47eO3CJUx5Ak6EyeadZmdqHKMSsALB8c2yAbvdLEa4gWuxU/QDgzkL49xIPk4YN4bWeW8b
Ditp5yTBLIrJ2sUll0im2grNZgF/vHX5kKV7k6vA5mMHFP2aU/Mge5lBZ7rEm20wN1tkhS4cM+sP
XyWhnNsVSpmx4di1ha9NLteJZjHaxTsxlFUQynUOjSzJLHRxYeOs+N293pwYXGFo44PtsIQ+n7ru
IQ8qGta7SM+8zbEYoaOROaot2MlBMvo/Me/+quFakN3inK0OP30TgYPOFmurK/h9f8YyKEv5lIFq
FPAsbflmEwWvvavSfgm1OM/DdEhlBZ8L63pMA0h5a+NZSgzd2osAo8b5McdFnV8LKl2Y/vIN0A2w
l6/r1lJsZsTDYwCvmEgDF7l5qY1tI8oSL2WV8eerMWWsD34RVZ0gVxcOv04VtfDGk74VEddkOolT
P0zvX1QfdbgtrmKKnL2yf3FOyiBayqk/8MFawFHQXrTE+It49K81C1aBgAKFuOXqnh8awmyqzeFr
gVw+rlPokcpL/Ns9uQSxd5iQozSirDTozHA8Cz6fVh8wwvuU2JgwI1PeNNvae9SOYZd8QnAq9TW+
Zg0YMH9oVcQKtuvQM3Rg1K6+M4BFB4zeQsiuBtuL5IZNQUTjxRAxByEYFHr1/yTLXmJ7EKGVov3I
hC/du+7FLreymkGVbS6fnP7iRHWoQCsA6NfqaK0C1fKFj4RnDicUoxAnzL1TCuLjA1VMFnJU5Mz/
F66MyX/GUUmxCAT1lGw1tgz1eCvLkRcDo9yR69sHZ8Zxn/1U6G3smRRCt4ZvmBqAe0IW9twiSMNw
Ko1V6J1rlrnIJAhxhM8jGYuHMX47h9omKJupqebGT05Dt4lvfK7ECEBz1cRuAYiciJKsBgyZ6a+K
xZIfO2PbMq/O1EsWbBk+H64bPK3s12JCuhpYdaUF47C74xUoI8YzfYCP460PluVVPBppBlrRnT6h
LyxCYr0pkPziCV1nwyyyGqviD9rXpyujGR5Y/Ga14TaC0LYXfzrEf3uJdPBm3zlNXBSDF5JWAxuT
Ggr6BKbCysG3eGP8ZQ58pF3QCbffqO5crYKKWELqlG3k7fHGPuzhps6Z7SngV0Vm70oWxjvxEmX6
M+K/V6PrhsbdIwQkk5Vbj3Se5VuJPsRbruacpTaKozxIw+KtQf+h45qb20ArvTbAcxfMsm9mqOub
z510L15PJ+VWkGMnvcDd+mfHoxGuBW7SaHvvLJ91j7JepL8dyKV/70QVU6u8JqcZm7gIjtZBEKuE
iwfGu7vxlRmekRn6X7Zq5W1YclYF6dBtZDThITfnnOdSLjcdIsguMcTLinXYso1YbRgiXMO/mT+A
FchGbTKd0EDdZVoC3Qsg1E2gRCBt0oyGpUVZAPEVSTN9T/1EEsjKAya6HUL/ZicioVrOyQt0xHfi
F62/JiNbZ2JEKtM72LVfvL0M4+6HQUcb5d2dAZDojpxP4dtMwlfPjKVT9cpxynVE31YCSGOmR94L
oHKEJVV3EGYpPlSczili4sz+x65/A3t94CDahr0ti2v+hd0jttop4pcdZrr39nQAtg/tjJbm8/no
QfKgznXIsNXvsrPxtkL6Lc3BjpJYC87z5VhPbPmOF+TfdQdb583UO0i8a4O+oQkz3zCAhvafYsOI
i/K6rzhk+ln+HfrJ5gMcHraqf1GNQwKpSdqBK/3WlsovqFd1wOozWbxyLft4W7xWSwSxQJwlSonI
6r9grUOUCqdXFDrs7FAAxj9xPR+QaXHxP5bAUYs0m0r8H6Ao77V9WwXdp/xH9L4nW8QrJiQ5HrV7
SrVvRw+DzplZMeTvaEU0nFT+sh9mquje3Mi8z56WQxWtApYQl/IdOJ31PmuxDgAJKB+hso5vjgWn
nPMpl8sZgEsamqSmpBXPSPJUlfU+hgxFebIzgNid0PTOtDJ8dO5xTTHxS2ldGWhs7L48aF/2b/gE
iXuoTTB0dJnUPsYh4BhfCuTIzI9aMe1agYKi3ALYohWsfiuMFAOX5TmVF0CSmeqDJaBBjXuLDV7V
uS+IBOZPHxG8aPBxHo67rnrSN1KO4QRge0aynmyXSTr2Ea1Kqnwjz9tG0QaPyoUJ7kI0YrDctapD
XKLioo0J5eh48ylhPwJw43XnzMv18Nyisv2Fi/APOC32x1vQd0O4UJqzzob3fnATd36DiMvRBNdR
bC5j42ABvrcVHHX7Dec24nAdbyyGf1/qmjtH4rT70ndk4156M7OPWsSO6h7cYhfNsDtQDTNRvnmo
n2CrJwuAL97lmnvqxmRYWGCSFqRBgGqLp7KowNxAOUf5A8XFia4AvSGalHAvoWo61hukys4PAXIP
bfVmkroQOBekkHAYKIeWeZIUvjvOTKclAC//x38PnnsqUm7x6XJ3ivg7tqrfcdQikTCGE22+f/Ti
M9r5kooHUU0+MMj19ESXwQulSUR3XVBtbkhpoPy65Mg+tOnIzvgYXse7d3cQNrT4fOpNBL7vYqDf
Pjr1cgwk8GGnAvIE9EGoJpuhWG7+rNuLLG3cMIx+7t8Ty0N86QLgIlv5Wa5Xpej1R8tQTtU9ldkB
lwN9RRRKMVNVvZ+yr5hfHL/21gYkPuFe9Mmn4s33OxXZTVxk7QEjZufNJ7w64YmuXc5P72D3mqJJ
yUSO1Cwg6GFuuH2Ia7ZB9i+cOb6YB2f+UY4qG56WXVOvxDmp/pnLvYjXqS3NAVeFOg3NNit0nR68
FwOFnDTbU33gTCdTG+8N2Lq5CHGMJ1gOdu+OdICOEfnoWi/MzcSdyQqGzGZlN9YooWf2wuLv4RcZ
jcBzE7Pmu5FVdTNBLqqD9J2uiL84Juhvi1NXG7RSjXXgTjNCRgx+dk9Wb+m54GnCQzPI7EWtToPA
RoOGdL0bwF602+/it8P4pLsay9uV6wSwNElYyfrasMuZDS+rtG8IAJA6wJ7kfsdwwIs0mnikHpAA
eXyM0JPCHeCZEgVenykuLSGOk2hgE+ew56i5CByWa/C2HzRpxg6HBFQADuQ/IgD/T74IzdWcToKY
RWuDDrlpzPJ9MLt+HowWD49+jCa0ycj9KoqS4+Mnk1ZlgOwGOWLLc97VUJuczdb6wwzH3H3UfmVa
6+zTZwPY+sj9BCYtuRRl7FDOK+W/y8Ovkfrb+/uyGgTITICRX6EBn4JYLT4n5oTlGLdaUjQxKAdz
/jYf9M5QTbKSmPC5iOj4s1QBqVTRbnBQAVwdccRPVUya+wALyRcBC6BaDDybrP5X1Z4iStrdLXZ/
/uaB7B5TYjHWHHzLtqDs95IOInd0Hu8UBf7WuFklI+c2CwGZnOPjvO8hHiqq3ETmPeiC74WBsrCQ
qkuvBPHa8LnDSZo1pvw6XqeyHrCYLk6BUri1SfEibjMZjsM+dgyIazleTG0SxxtV8N/9igR6dNeU
IubmSYOCGQpIT/+JapctReuZHlgzKvQJgqrQ0zpcLDQUu5FcXOPb33iweD2JBdH/b/JFf4ZDPCeP
mapHNS06FXYuwvCC/gl3WhCTXJGpTeEr6fvod6+z+50EaSIP90DKy78MaXr0y2qFewEQXW+C1db2
VieIusVDbEIQmnYKaKepuezyxfMjzVCGBNgiuMzd0X3duR5CuCGmjWmbpJZjhIRrq4ZAJ+76FzGD
/1NqbnO+OymAFShjV7Vfv00AGhxCZU49bN3v1N8cP/cVCrBoAB55dzfnJnDgMnJShYY3gDWbZzre
dHKgGToOODxtkN8U4AtFIwkvaCcEzfuOZATjkx9qUeoIl52XWF3vbxK50oU8xwEbWX1ViW2yoxqf
oi89oUFnhvBcoyMK/Sl73X0JQ3w5wlRj28nZQ/ZVZLk5IIloSQlxZ6xCNUvTdvGXNierPvNJgLaj
q22deEHzUmk9U9NX/1uDsCU9DLVVoBCIWRMHjlQSkgffqR5Q6lngD0Jt3RBC8zmdDS40swz69y6O
9JuYVEkKPR2mCG1ORuE6Ag1lGHG16tGs6aC91EUT20VOOK9jVCYY4WUDqyJCI9y9oLibvaDq/fEX
llY6RnAP4ocfoK6lGX7AnWvclLEfrLjUIa3jiNZG2MdR/e8eKo3nIm53Svd0X6EhRFAbOkyi7YWG
IX6z9WYvM8k2riw/i1F8UrnZMW4qTMpkeeTEqpeKG/OWQWFDOUgBJKYr8AMt5HgNKIagaNT3nvjC
yfY/A+EsLk6DqFcl9uKrXn3rPGSDz5JtQ4B2jcgFGld4SyOONx0jkthnvPkNoWgq2nlcZdEakahM
Ewg0yXd5PpfOQGomKV61KfMzB34/jlVrobVi8+O5FZn4uxic++3Rm7zG0IdGX4/S9DhyDyg0jwLJ
K/LAWebtRVJBWb6m1Tt1Gh6lSnCiyRHXPBl+SoecyCUD8gKBKZD1TGTEjNFt9ftjeFjLo5l3bY6y
B5V7XA71fJahHJrKZRqsXUUh7OZRTFeM7RDYh4l3QzF8aIj+U76GaSRoPVk4Y3WKZmK/nMD4RWuL
lfNqkuPQnruR6P2vT08P+XDeFiPb5nOUR0YseF++FaHnBVqC9+5oS9gex9x5rdqlkf3vmUTauuY7
M9soeHCZHQt6eQvzKI/lNm/7PS92K18AK8Cl4SWkUynuO2O3iOhjOccpODhPmPxBbmVMhavua1YN
PSHs1J6rVnDa287ZXWIybEDXH1KlcCceQJx0FhLgLh9k90SA/0jYJXFh+5weTwGXbaDct/khZqNT
AWJ794mEQ9+UwZSzkqCLFtGn32kRSpYu3eMHrk6PCb5UGjGtLXVC0i8MABKYMi0jjy5Z+LQC/Ao0
0/vcfVmAQABl9aoqMLPpNJscYXSdoyCw/I/dWz39l2f63Qi85MWioO8HPBBVNQXek299DmAfoQXY
OWcZYZNaTNk2neTg3l8elSPjEp+Q/GHEZOjPZrt6JVOtUhOEr4KxwXYMy0EwoVyhayd3GO60p+xK
nTt0kOWLgo5EzXttOaH3NTE6YpsHujvImaRlQErFUfUBQKit+b74EFUoqfL7bslNOdcu4FAlS7Wi
hKnX52e/CWtwFuIQweJ7w4PbEK+E6gnUCs8m3FCmZ5bWZloBCtU52c20N1XI6l6+PVY+Ul7ANweo
HXNuDQZofTZ5jreryTFgMD9bdyx8Z7YowUFbNcXZc4tVveXZGRivUBlBXVy6eT96dGiu+h2O8gWY
wzsVYwVtt7BcWNsi2VKiS9FFbBEWikdP4/TozIp32XTfZ4rlmTF8FCvr+t1iCJU7PerlohcombWK
L5/h1sNL5zoh5g6lq0e3twEsAXu2mqEzAIuu9Xvt40QdOdWkg8/pFBZ/byQ3nV9BsgivMyu4DtUz
UG4NnWzGqTUfKaRUcC7ExbNDXLhx00DKRCjnextElzKS+mNUjl90TPQqIVe6v6XMO/eqFQ6j1xcA
hT/oL6hlmglSyVlpU2r+A6DBeoKVhSKKKxUMvHofGv1hfHeozdlbP0YrvRq/QZ3BI8G/Kgj4MMlh
otdWQTrwU/HV+B3lOOAZouH4AnrsLgCC/YzvPReQW2qrsoIzazKBHfNLuJqIIWMHi7fBRrCCLTpx
SxA2gTcApKWe8wZR9OMDcoeU0vsKAAy0k9IXyLQax3qBGlUP78lZJaad6cMn/6u92v16Ei/fa01N
HYZpYYH7XdsCq69YCT+1VAlTxHvb9JdN3DIp5tUFS2dWfCBhpgJV1Y3GIu1OaPlcj3wl88x13e2I
nVsnL0B0cjpRuJcMc+9MLbojV0RbKA3ujmUmDvrFfiO5OTdgmeX4yX1T9ZdjP5ypexvBXxRe1Gui
3RN39Z1Zi9/+E1lm5G5fGbQA/dmvHp0KSnONv/Hqt5DSc4WqMmFSfIur87u7USUuNZ9CzR4TFL10
Nng2I8qWoc7qAe4su7b3fvYdRP+MI6oZZTwuJ1KTG/4INXFSLG4l4Nm42pq7wx3cryiohSaoL8cq
UY1qzeQn7S5vzUGK7TM2ZAEwtfrQUU2VS9ld0kHwKXJ/txGP1sKo+Ba3PF8zPuN+CkHWN/O+vvAH
ODgD80FaqKcDDRKQ94R5jq/cRMWFuXqQqAzUCVvISJ2hXGFTgRUlYiYrkKZ8JSBlOgPcHFq2/JFi
ybQtgv0irtMb5w6992Qe5nKFnieVedabtOSLEYeDFqIodm84+U7tpxHAsQDqi1W6MkD6UVniAZ2e
I/hyNHVbnl62KvZwJF8FE32PxBkWVVd8r+oWI3AvNZwsO7MZ3l3VgUwVfZhXKm7h1M5JvTz/l0iT
uHfb00Ksp+XUQuuxhqQj7tzP7GPI3GpF2nuQnAAYJItoTAGEbZTtUocOcYnra9h9qNZZea0rIoCO
3fP0tWaxRO2MZx+OJ8TDM2inC9X1pfbZqgx1BBE225SWdO4uZESrfTnW+gY/b1iF0G496hrpTHLc
2B+A832XLwc28jNYCZqAoE+v0zAFaP6LUUm0Cahf9xDARviPE37ShtoYLQGdRgOT1yAcISIx5em9
gO1udPShXyGAdSjSL1BFVmr7ozrBRWnfJij5+mnN3mu2d4HHfx9kyRaDJcoav0URcHT+cZeRDjAM
9IG1quwNIL1cyFtE31mmOQJGIX3XZuAdu6czyWP9g/QHx0BZpLcQVOaku1xRRUhuzs7HevXJuuJX
NbYZFoBUweL8WlCXFxzvNd23sLB/mOm1QT4SvaaAcOuHo26MB+TX8RlJLKSnEztbnUa0pSicscMi
rSzKzUZkO2BnZiR55mCrNIerOcNY/i+5/Shh7Cr20u1FPLcVDqNroxHHv/KZxUdmB6LwBH/FfTnl
0cMfOAfylHkoOFOJlaFHSWBRR7lsNnFPRbDkJJPD6P4OCvEJge+fXG7vIzMiqeWirfv+YwskAraf
syQ7iblc8vysq98wkBpVSBg4Xj+Qoh/LzM7NwM4CSTKNfBlCkoWx7YvZXf5nlsdfCIa5IDjIiEDl
Iz7Vo45kJ3UwSfx0D1RnDMp/QH8t1I5XpMGSajVxXak+UcrP9OHUxka9V531TZgw5qcJO3m2ncH+
/BBI7YN58q3oe/ar6M21bCKYBOJHZBY2CkRPFw5iGd+8MjY3GRbd4YvDFdCzR/w/Vxs4U7uXXfAc
yL078A8zkAufP/qR9Y7zuo39TiYIFw+8elyYFC9pqGOdvyuiDOV4Jz7OW7JPuvGPYsk+iYmesrjR
h9NQjVRp3LHKNerhEYlX9WoSE9/dXrP5CNLyBIscNozPZ1YYflw=
`pragma protect end_protected
