// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
r7luE3jgLgy/rLhChxw0xcGREIqsb6uS5Jj4z22zBRqPl3e3aUSCZ27SDfV6PD57wNnxM7iBRBfW
6RnMiXzr7XVJSqo2RwcfX4vk95SM19QkjwtrV1m4pq84MdhXGCO5R3SnbgekeeOiOBfNGiiF7vXA
Tit98Kfax2RO1ISC372yUJ1ulk9uzrX0ic6m/wH3YQfe5c9YgEX4pQEOGPp6qWvEG0L8JngRsD5P
07z29td8wz4AYCdmaFrfOZd9KO8s89UvMKbMdawIzHZGsjbHrliBOrdi9pY1KRLHxBmrHHrI8//d
8SPDNft2IJGVI+AXnTYvw+wBiMGvA7tw1+3I6g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
Sc+bbcoO/RqSTOAPEJ/UEhwUBF10I/ZpIxxYvrchHsU7iXsCWacfcLGD8TmDGgojSYpSuGpPNuqZ
kYkd1Os3P2UmuntB6n8mocip6XITBztV0xx2hl8rcoeiYSCdBkvkoqdcUFP7Tj7KT6ZcPWlRzaeO
wzhCpw7UPioZ3Ctm1WY0JSipCUVuoUGda501gWWX81N1ShiKEg1ytWfP3ooMPz0Ql3bKw8GuNoSZ
SlpONOBk9dEPjKJPxP2b1KioysJwBdUnMH1BIzUUN7uqw4OgY9SwOs0cl8FJyVhzcXTWEWlx5fmd
0S5cVkYRNNi81rIDqYrnDjq99qQ7tgyhACZMcTVvx+iAFETqRaZb82AoSNRvzsupgRbdggqzeeC7
uvo3+jbuBTunNGFzWGvQAil4oSnXaVgtAWCCkZQVP6iptnJHmm0oT/46S7iYRZjLp3amdrwd36qv
y2rhJlvhL/URiNK1WJPm2/DTZDtqVqMHdX4CAAGysZSGBmz9hf6iG8/bW4wgHzKgwTqBzJsrcf2Q
eKLXXmaoGvQeMu3DCvj3D+aXzZ+Lizs9CqupL3WpVWikRsdKaLUf7z7yg5yPkHhPJD603csFiwHF
HYvafjbz2GmwP39p+u3M4FQ7W6yQSHnWgUJ/GPVAs40yLZXioBbbs7iJcIO2otphOUGV7Kxj7N9l
cNFFimFb0M6FRG42wXzlXxGbRoWmcYmegdf0a1ab45u/yo3KF5zyjpE0CGysh8jvybf4lnIHHq+x
Qy7/Ei2eHFb36wBJYJpe8Jh4bhCrja9ue4W3G2Ybh4P2hE8EbmyiaOKKHcSg2BWuLUHnQcv0BHKu
sntPiMyhLdYDWj/oymK4UVrveFrQuhZvVU5u/TA34yu0hKhlUoD71NrCMv1GdBUafA0BqWBUEpx6
LQSbOhuvsfSnB3rhWDaYSGMJo3ZY8AWrjU0Z9dpt0a0K6/V61zVQy3227Z44b0vfQJYxsd0dpNy9
aRGqCawKmfRztOoe8iSimBOjijO9M11DvbvWq/vnoOUCmiuugfaqqaIckkdMoS725hhElBvH6Y3N
1Fjs7dL1auJDTZjnYbDrYA08sYTBO4heDEgBgshTysNIB+eQApcrcwo2KLJ7n8X/rg/DyzpE59L9
UbeEnlsAsAKm1Os2SX6otm834pkV9rvQNkOSddTowi6NmQ8dcDKiyG14iaz+4Leg5KUGuNZc++mQ
0Cf06Rvyak6fmz+uoq8udfT6yO2nZ6WJM9QbayYPzbeDEW9aEXBs0Sw5wthGpWMqg8Zije0cGJDq
faBu9mB09C/0PZPjgkHBvcT4Y87+RgSRJ6XMC+xd/h1CrEWpufTJmeDctUImcASDbNyTe//rehg3
b6ZU4ez9rVtPCpbTLy+z0wJWT03sCGIlYAh0G32Wx7aAsytadUWQs6/9v/6dpo5fI/FAvf+k7Th9
5qLFP9PIpkHaSQhZHLzqaRJZsBviNAwZD2gl5EvoF8Dt66XTDrtRXQK7kmyoUPlMqCIiuJH3aokG
7mMWGTJey1kRl7kYUPYivXrYO4HDwpQy/s7JxebxWp3btWF/Mlzuyt/xJCfmIKvDhLNWodpbPoK/
JK3ohdqtolQJ7nV1KMgM3gQ2LWkpFxNhB94y97YmA7oVkP08q1jEtuMEafDbVYwg5Xbmf4TOcCCD
0UvjgoeQ+Q0qJ4F0KeP3KOtjCtivIhXSxwmXNyBrVhIxmgOCQxTRXx0zLNDGVl/f05Wdt/s+BnT4
tVdWRZC0CjuYJgXQHPj6JX2R7/YRFNu0BB78Ii7pMlFs1EMLt568EO5wboQdWexa5IPnP5UdKBT/
1HhkVaqt6GDlxjofkflgyveDWWye3Uij1e5aPet2kc+0iUTBCXEQDcnfcmAfa9wUVsyHKKtCysU0
oesLqQQDRGVyeANWpVa+WKi8Ucb+fO8jYpH+allSgQQxT8c2QUWbi2Q69ieK/HZKXyhWOWPzvkAS
hhbGspwfoVel2dWzFWch4S6ugOjAd8877Ssq0yWx4ZNqOo+QoybXxUw1ykvZ8lkU8Xt1QSmX3teR
Aw5o19Y6yWwCeRl3HBwStVr41eIMhFIkjvI2Q2TakcFEcPKPgp0XVeCs9b5v/zkUo+OpWm+i3ayf
aPSSqixlE0gG0jmQE/hmuKLEc8hb7h6z0CGgz2rFjRCUZn4XCNZWb9U7dM8T0Rng87+qxYEEBI/0
pLz/Zri70mMLlmUrtIZs/zS7/WV20TIb6EneIkEXuO+QHa4thKABiuI3awxLPCLCIFoylvqWbje8
Mrq5rBKVt0gj4fFhiln8l0Y2mJAzdHpaOMKhhZ8/anTTIfZa/t3pRY6lZbkfQLFf3O7M1a2rsbsi
mSZoUT82r2T3dpei5/bs7hSk0jMr9i56RBXVA2nf2kqyh1gdLGwPxwO4zbm/uSHhZ1dpUx1w1rtn
ugrGk1Bcr0lkhUBN2oi04rZiZQ70RJy9tLhsZhjRB+YyCb98IlEcrBi5P8Fv2v9+NhHnuOIa9Q75
Jd9IG9oqVVY3ALUYsWIqWbh8jOI/bk+YsQ+wFyv4LZ5JD3gOAZdRS1gfn8VEwk6OEomCNf45SHHW
YK8kYPzToR3zmYGDeQ4Hr09mVEL/n5nabFZ9LuhAdD+/1D0kQKSeau/sNQd1Ojyui+39xgyQXc6G
lTGbxxKvNnzDh8SJ3l+f8Bf9lsIYAtScWIJeDeOR3axu3z2J4tz4XGETUXwD/80ORXDhMYPYHqJE
bcBBW068MkEJDsXR0jlfG5cINxxxHxiamRtWPm29+DqS0aNpoRBrCNV2evF5kqSTtL6OInVPtTM7
7PgoIGvPP49ggTP8aG1pflNRSllQJh5EcIcwHhy8vX+khGJDw+hqOGsfBexKTSq3Aq0hcKIOsXFP
eKHCNIjYHp+aOrRPEyrmAWKb0axTERRl8lxoi/Ogqg9EtqM/ba9ZfkavmkTNr+kfCujw/NL4Baln
6h6PBeILqOijPpkXN0W4uXu4i4XSSwKC485nexm4TpZh1fCt40ORpPMoiaZ7YilqG7klXr1ILAb/
T2QFRfsgT344FLQ6C0aEJ4hCntS5C426jrSKLw1VRA/GPDRVbCGiy0ev3lL8RNdjB3I+FnyQ4+g/
IYXSC6J+4NLlaz54WCDueNoqdXKdnuTJRVqzMgaWZnmUGs7zklee59IhRlkMggZgCgSR7OhybO8Y
sX63bKpARLdIN4clQezBL4D4pY5ofXbYI/uiuumxCzXbZkOnD14ZvTdFPY3PNn/UzYICl6D3SVar
cov/z16Q7gwJtczYSpgAcllgg8u+HTZYhB/AUmTOHdn8NorKtjXYD2iWsq6Rzo6iXIpGCVC9izG5
p8rIZyTZA1s9alVVVA3sIknE2BTs8Pf8+qT1BB2HreXHLpOPY9EJrHTAouPvlMCGSq19wxlD+aUB
QS1dl2xSXUhy169lnrqGLyjmVoYKrWIwBkIgaatkQwYOgZXwTUJJOnyXqYPpkPEBhbhByP3zy80l
VH/5hU+3MCRud4gKKwdAc/CGWA+9oDCNMVXZm/rt98jdQcGyTNBty4RGRfXlTa5PEGjXrEu3lJci
OsWV+IRJHwl9vC6xhs9ggTUCzWxjqa9Sl2SKQoktDw5GbDPLbLACwd4pFQa/6+bupNGqN/u6u+ZW
srS+mHhb9PNdKKbRGdVSq0m0Gbxy0ibtsSwTnUZmn6Ikb1LhimFnEL5QCEtoaMIQP5gmX6ypJx+U
hmKIWgzAnCiGOX/XUjQIDcg5nu0GY7Tf9bmVywycaBZVUVXYnSc31imby0y28caD7/pbPWfOob5r
Gkj9qxwHQQKE8fOYuIJmwfziz+iaOh/uDEAnayUzEGi9Hks5ig7lCUZ9nEn7em66JBkVULkbVZdZ
46Ny+teYQX7hAEzxEV4sM+1ECh6ORKLXvFu3CBf17pscjp3ykO5Achzdi6q1sBD27p9Hc8x96vIb
pthX6lEcw0rczAXGJ/En7meR3Qcv5caN+dmUPGMKYkw5c39qG2AM9lhaRduJjBLj+hI+Y+mLIHWK
3mOF5zyW9YWF1HWFwODa5gEzKHvoe4IaBjg9kADYmTorXKjZRZlNfd9KIN/Of9V1rP5Ktps9ODIk
IErHT3hM/jHL+BJZ1qCrtvM0bf4KNmOhLBCbNUZaaSRTfyWYnZYKLQJOEyzENBV024MWaKuG+oVg
DNrW1LDf2/F863zC9mQvBTTiZPxErlcLH/GRWmBjX/p1v9bSzwUrgOltQE+sIy4Fk1fDXx38rOqF
DwdlQNhEMg0sXCh7wC6oBg/ywVCqx5vnRuHiws+aggxCOvS5R3/CmiC2Tont+OW1CNfO3k2M4GZr
M3gjdDnOAvjt8gweMSr9PxiVbmWBgG36hRZgo9VE/vsLaQ+RXUMwpXC/71auLmncjFInzMYCKW7L
6RbB9XPBEJZdmNn0ICuryp1Nen5v/jsV/ax1AXjHpZ/bpQ9alnQ3tk/8uEci8X+siUGye2/zXhYS
2a4936PY8jR2AXt08AgTcTEPsDtUCW3Bms2Yc0s2NsSuWRR25mRcdwDzOk04Sco3Pb6eI8MhoBmD
gxxXIku9GlGd56RggrOG527TjRPdtvFsoggHHotHASCJfSVBb2uwEBacWzFb37IAzm5C4Vea3qWv
EePLvtMyiL0wcthJq8KN7I4/nnBCWhNvf7r7G8Al+wtOyICIMiua1UIGaRkgQEp8KUg3LTQT/hyF
FYvFHHGNyjOMElTgVhbWuvqPLHu7vOLRZDZgdr2qAVTIzoJ7sQqt1qfN+7Q5xc60P9NGmJYEbA2z
Jl0z9rrgHmuuzwmERwNdD/Y/gNfXh0K35H4w5ZCyzthqL1bGBLV8iCJWrhNw2KmpwBUFLP3yP/cC
OC1pXmdVzblH2Hcm0r5V+gkCUR8z6H9rOQoNJ2M2TBuuK4dluBij/WceA2cpfJFu25flWNRjw0Tl
vGEMvelPEUTJqoeh5u8TGvgvb+5cNttdRvK6dFH/JfSKR7/ZpzNf9luMFvPAqg5GqsddWLpkBDHb
qso1IKrCnFRtTRDThBTk/EcM1bfB7JQQeFnsVv2sk+J4QWeNAimymlPOfn9op0SpyuxJuLVmUdew
if2mLoVoplC9iQ4S15UDhoMXTON42goZqnzGYSRYe5qghZ8AJdn47srxVZ/3t1bS3wzBUurw7rsh
PvxOl/IwBmbJJI6dxAyCR2Q6jmCmWdMophuDJYtjQBTYs3XUMzPce6X2Ioa4yEAwyBhPA6y1qjmo
WMiwyEk54G12Rnc9ZYLWbvC15WhfWcJx5/DBUHwJpBPXQLChKeltIAk4ir7oSpcF/2mF8vuVuYzO
FSeI0bkGE8dbLjM7vQLrvJthu+uE7afHxfYyvp7fsd5B+O4d47fRGrpyF/ayPqfbg4ADxkvGilrx
SBZm8lXIAsHXpNz2khtb/HmWqlCddvQCU/RaoXFCLJFik+Ei7DhmzU7Ib1WFXjVIYiEXPdLuaHlO
xAPpJ6JlUJ3U4tn7BU9vGzdiNrwh4a7/dwseabM1EihQtjRTuwY+kbqdtL3Qj8N77KnEBAdisyEv
MHxXcsn3ouCumMfa1IiTzh9c6x7+Jc03/fSUUEzUT6ydEO0SH4crMF2FPw6wivvxZU6nxk9/QMvo
odvH8XntqqyBD/91riFtk+SCWigQ/o8uuGRyaS6EFZcb5MoaHsUCaInn1PPWielp2QwQ01j30L22
vmJciitffuqG5JqxLZn9v3rcd031C1cmbECS6WgyieDshaE/ZOtYQSfr+gK+wN8qkihIfmAKB0la
alfaIzaZirDiIuKBDIZaeKED4x/+cz1Bw/ECMZMUIDWazQxK+eUKiVNl+dTOFEVdUlxS6gDyVm80
liRdYG/uoD06NYuemch4gVTrxXWYJxTYIoxxW/JwECxZbTUGV+NYmdAQL3LPKqoGVMNkOv+KI7aI
OZX5apG4NfS4ulaxtnRNmoMRt3vas9rafUe/djW0lFyRl3b4iANHG+tr01IeBS2gHJa5kHNcMgSb
NkCu4GO2d3vhZquEkl25cW0ITL5J9HUNw0+LpA3v4wXTe77axf6mLWAJYZNz0vMMhrfnmffSNsxV
QVE7T/0kqa9t4R0ytwb7PE4aoH18xRPILncR1M5VyiCSuTVONxFoTC+Uis6oTFKtv/ipddLp9q4U
dJxjo1rgHlba3iZwH20tAdMvO+TVtHEUTNL3DdOnxQhlVsluP7/W810A8s2wXGbZbnIPKKeKhXHW
znUs9tUm0jUe/c8MdvWsnuSmVsyHy9hFCCXmIHBRs6LSUnsnX/ZFzAThzB+TpmPF40ON3jC/wi22
b4JeKofd7CFcAta0Jg2WWHH0nI9l71kSSRyUBT3kyPmnirOlCzocSNRiCFu1ZNIjwoVoqujSUD8G
tpaaVvdD3B9nxXHmSfN8jhadnWc3FbK1J39Z+1oPEMpEiBZj6y2DS+Rbym9JnXgJd9HNr79hWG8T
LmIhdsFJgSDic4GYdqmPUMrd7SClccD2Wj1ZDRhRg4+4CPy4BzN/7uCtY3gDgVIZjbNPE21nZFdR
l59fnUR3yNBwqPsui5a1mH7sHW+sfQzxSJaA6fnWilciAz7s1ZGzKrCvR//VZxxi2KxU8Mb7Y7JA
EtJ1W/OlW6y90K6IeJoqHZBPNzQduFRjarAI3tkQdFHWM+wmpiPQo/NbehtopjM2zUd6jvZhLziO
L10aIltS9fVF8ATdn7Yeac/UFt4iZdNm8jtB0qX1/Kfc4U1prII5Oz4EG6cQO3g9vK5+amOG0KYm
3birMKzWFav3laWng6pKHX+nwvlCKtxtD+yi/++LBJoDsy7zVrg7yX4Tmch/MgEzFiqmqkzLTIfd
BGCX6zs10kFfBaT1ORCH6Hil6WdAKmUMt+Cg8nh0vmCW4HbiOFLdRb6WTQgR3hYVc0vYnE+98/aO
ulxwo4T+MvypZUs/AvGIIuoa171Wn1Mj9QFe30XRL6axi/P1CR9pxip3xK8f57jZO4N3eiDolLis
NvG/wL3e6m51Av4xewa0zkj3Lg/vBwYH9YZxJUgmZj+NKjTuSHyggn1/NhtXxR8N6tj44ZMvKqHB
xZxrJ5NgzbuccM65POcu6oiGd+ccOD6kubGUl5Q2W8StsfgrPtJu4KyPuVEYF2WRgH+DpOIQPj2c
Xdwp2G/OJ8FTgj7wZ1Q6dOt8HiE/9VSoDKyKpQKu1uwL9G98WcEzH9HeG887vLjonuYQVkrx6vYs
YRC6gX9FnSESOEKJF+5psPPcR0ir0tvkF3kMfOYi68aJAFuAokkbA4UJEac0Rdx9kbnCLG8CyYkR
WpamozuFw6SFb9U/kToHfw==
`pragma protect end_protected
