// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:29 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hnkwOZ7gZQ8AuP8Z0l4+FG5DVDy0qR0Z+ZbEFpJbnrxMaHZ/5jDj2hFc5u2U1mbG
SIF/bxHWdwOK1x4mvHCSkY2Q1a11g0el8Z3ecmN+h5fXc9BBAMAQLbFjehb7vTNX
pepF8o9FH0+JKi8v2R1/uosrTsJA3EOX1C3fJhfPYR8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10304)
+lqUVPDmutGBvrQUA/SvEssTH9t/KSSYMzfcSsAQzGvV8aL2pnra3k2I0IEkf0ps
Y+j+yo/iN8A3n+Y1rJof5hHd3bzIXgYwPMFK9DPl/oh78oXuj0tU+FnhBbya1T9s
d6ODBAjxdQe5mCVNk1x7zuu1vQ4EVfGtmR6rv5kQY08UwbIeP+Z9ZBqHStI3S8Y/
YkjswXSD7KdLzwqfdRwMGB/BNrcrpY1RSv5bLRIJd565TwybbJPYYiV0dI2yR+Y4
rrEO6VrE9Q8ryzOfwsYJ7u9VfmEAUS39MvLR9jRXD1pGn2SwKjqVphZ/Y55612Ue
IHFu2FklzoOCshHWcQIPtvCoxh86pIwabJ9TRHw/vetYEDySqy5yhhNGQ8PtUE2r
NZGLJ/2K2gRDxFOKUPqX8tGJLK3IPadwgOo8vr4+Uv0l4qul2bPveIQqR9QF9f1A
HffiZ5X1WA35D6UCLmtq5zF62VxBicd2kkh45eAX3HDhY9dmlO/n4MFaYeC54xN4
0JoSNDeqgZ+9jl3Jw8l5173ODUh2+wWJqCBGHdQQmoVKdIKGU4flT9ByxjqiDgqF
e67JTd+JL0JOL8e4HxtqFZZItqEJ+bNFxJi6PsCPhvH5Ze3aBbmit/1gSXaJhmZw
V/lENzDXBYuMNl8ERG8JrmFxpHpgXQ26j0brluu3G+dKo7ZA5Hyx0fJ94AeucyOS
e+2+BOtZDn2wKBSxpxWXJEplHM5oXVSZZ6FwawPD16dNzUHeZWYjxkzIICuH1apl
t45rwoQrNLHBagZHr0DN5E4woeqtA3dw4J1aTCV4o8ZezjvTg+m9nbly8sPai21i
l5jDbbFguGGLJyKhuCqN9zBYehrW4DNEoyixle3sgm0Fo+uqTI3NCUD/dOskb2qK
lwmTy2e+hXYuqOz3vrYKUTogzMbb3yUyi28NTJoSqk/m+l5wfxNy4FAk4o6em+2C
MsMUY1iCh1NzSf1iiuYpF9NXixW/SJHQPkncG7w6k5SJKleuTNBWB58WrljoLeOR
U5owiXybBI9XxWERmWMVMPAUpgTWtuCl+gfE05YHW5RZJq6hEmrFsiUXN8Qwn1Cp
JD99tuw04eyuWMBpMrYijb7OitKfEP0P3iUfik388dsKiHw1000+p9kKHh7O3Nkv
nYJiOXl4U5M5jcvr0gty53yl8NDx6FZ/JzTEZ8Sk8WAiyvIK//0RqVz0ho75vOaK
hvlsutu0Czc55BYO8GPaS259CqN8tPdNQK78NfkfIlgAWtuyNyn6e5E2ZugrZ5SK
VNIh+PpchrGVEXHVO2HcMtKJb40orLfc+Uh4XEbDYG626XAGXOGEo1VSOmGU4Nnd
DPukycdZHXNZIBCjFry5d3sznxDaukj7hOdYly2ZkC44TQRinds0Vp3k/vtOaKi3
c4ci1nLy4Kxkr+j0MsNnbGJazkGnUXPWrcJQQOZ3oq3lXZGb/xPJ6SuibnPwhAFF
N6YHpr+uLCrJghzyKyxknRtcKa1esxLh8ckMpm7ymyhJQ0XSBxHG8C5LCghKOcSk
/ppX/H7riIBP2nhCJsGVdQL3wmvDdfUY6r9Sz4kzE3B72vU2/Q/IyUKUbWn3Xquk
/2rs1zdcU726xUJbQhmUXazKZyx2zbUa5SrtdF2MiVZYwZNzS9m8FTsIudWGse7C
y2rz+nq0wevpXGQMoz3td0pRrpy99OIrridMRVoxbxb6+7zRChXbs88EmEJKq5P5
nsW5c773btKA3c7tDMhDz0/NvDwLOOlyBhZLMpLF3zmwNdBBcfoxt6zcKO8lThmf
HUgFbixqs21EfDJInfHvii93X8FChu5DjJTjzlRglLa07O9joCLzvIBqCfdAqPBI
7Z2qvKAV0RvVIgNHpplI2tCWWzTGTZpTbqO0wd4f+9LGX7pE0KsgzY2xzemvlrYb
p9/t7sG1ZCsQyZug1U+X2yzVEsfiJh9ZypS5NMZu1fYXDgn94bMhfWnFTBprxW/e
OprrsRdjs8nh3dYFuN/scE/DHZ8eQr9oZQiWV+IWJwWdZxZ2B2AH+3kZX81iuAGi
DYvvzBB6wz5lYymBRNgxzv1BjTHTAxogXa3HSz2i9DxPdZXMPySs3e98r00vZryO
aakJY7DK4uygAnBpnm58qE/KgZqlIRrCbJ3YVjyyA4gQ3IFyknelyleZwcIgswMk
dCnlSkWvf5tze5wzXzLoJs+v4wkCZ2fnM30YoNs1/g1jREZNGZku9zY4FeEwAQIV
m9z/DNUBTJHqCy2bLYa+QfCwGISdcK5A4XdjjP0E2AQALAfiI5pcPd8J1mqCgzG5
CN7v50jv4FBrCDV6cI0424b0ydQ79I8LKQBBOmWjrboCDs/gwYkkv+Fl5lxiqDLn
J+BDPKpwMweSKq7BG8CImGnx0lVB6p0DUWrvewYP4ptRk20aiiQy+bajgmRrUG4o
2ehmgxeQYBi456o/rF0QxWZNSBx9Jz8iU3fZOFy9OrutC+XK4NaDhoJcxTCgPuv9
ZPbmPY9Nm7KyjT0uGuzHvKjQAHtwrqU5Q6Aq1rhtHX1pV5pclEE8ZbTm2ol62Nuq
UCLCOiG9e8N52TfiwdfI8bNdf9MXwPqOZtczgGTZwq/p3ILF6tF6OOBGXCcmFBpc
A9QJKsF4OaV51WQTkbfpI75BTf6J6jT64pOGTMUaevsv8D7oxKKW0aA4Yd4dX0kV
lsuq5CURJIHiaOMSgF5ZxDw44U2904pq6zM48muVoLIU4Zx69HtukNanvus70fih
D++Fqk5WunUn0PrNypy+2fWHA5SzeBjH2kl4i70HT2cMybVjtLgjRwk595HlP9dQ
C6lB4I0PtgY7DzHVd+BzrC7ZcI8pJNddkGUUqzKLxVM7U53boyjxMUfzqnB0Lkqn
5CIptZK+mwB2/S5gi3Xx2ahFEeWd0Vo2IJaXfVyDSGYHla+v45kpcUkl/3EBjTfN
gDnHWvFJgrGl7T9poxBTxfCm/PNjIx5aqy8vOfY750cPYG7A0ikAu/4Z/KubjKuS
UYQ/yeWsuBbDB4Q3jARreUI1605EvivznFJZJes6/cYjqdZUe9bqNUgeCAoVQPZ7
uV0+sRIZgiqeA1DsvZacBu2SpWwFzubOH+VcB/zLdnmfCBSrk1szBIu/kJ6G4aiM
d7FGMZsFuT7hpvyK9mAGumcXuCp840tb/8kAS9914smF7/XmTpkIS9R3A/xrCuQh
0y/YLAds5Egme+djD416Hba2Rj9rQnn1AaCYml5+PTL9Xx1zMUZusmX+AKuc1SzK
PHfosLU9S7oqQJZ4E/EWp/v77Evxd0NEUdM7Iy+4Vwdohi7MegTSmoOhd4T4X/Tw
uofrSW7i6bBz1mJ56XttGm+K+7huJ9v/p6Q04OUA279xbhRabDwJsLwauMLPHWLf
CXtg17uOxuCKB50a21o4CC4iHIv0VW9qwBSMO50FiTgwPYqbUkknmK5WQ2vjBzoB
p3AuSGYe+yC3EnI7gK/tfs2N0q50ibtRt/7VDk3mKIrbZKcVBJxcNVIdXtS0S48o
/SzjEK81P7Q+g0nf+k5XXBVjDXOruQ6PhpUXEUSd+iVbqwLOe55npgtDTFTeUmyM
Pp4QFqBjADHJnjqlsJn6I4zUS4wFXtrSgN+Qfea1TgGS2qwP+kStr3uLTVXW4i2L
OcrPcXon2IOu4p2ysOxgsrKG4LTZjDwDD/y2Mqp6Q6Xbxz7O5qC4+Bz9tgmKZ0u3
BEr1Kf47YMWZ6tid4oJg0vdvXVAEtuWIG/STDm02MPIy/Ny1EuX5PzacMB7p6TMh
ydj5JGWnmYcFu7z9pMsrtEHLUXt/5XYnVn4/EtBsUfHiL7UtLfIRV6aoe3IgUE0l
K/IBu7hudsKiNSKIHF1UfcT5O0fp2Uab854yl7l+l3vJ+jrs+UjIQrHclgDeGyq8
IHfMIUEKLr8irGHFeX7kq8m+x5EJdFJ5Aif0bSVp3K624L4siqIs/RzwOv1tHDet
i4EM779Yrnt3zFqn8tFQRgyNfKmhmGWpgnlWWMtNfAvN9odS23WYeLj9MX5Efh8S
t08+IDE6QhgOUTSa3RJ+pQLlr7n6U9Pm4eFqah5p5eOmJVu+NgJBYIjIw1ErpR6Q
Nc4DTAzfxEwOb15g66gjeASRP5hiKuyyrHog3RQpKCDd6xmelghteYsZ1fpZ4gos
XH8xO6E09cQk8NPTvUOzff4NQDVzBXdUYxomyEXxXD9xCyC4ARjyWS6eB/W8RBAY
bszVMyEvKhy4lmbUctXBgBJMnbUkg0SMp4XXWGf9fm5IyWl4GqBa4HcfmXknwJ4d
1/y77nLnjLtkYYJ/1ggydkYZbO8uKRLaHWKoWF4fQmcjB54DHcIOL17ZIJgOaNqo
26wvF023u83iVqXxb/1hWwpEXkosDoCF5MolTeHFvdSghzKRi/SQX76xk50y/JIt
hBkwD0NDoYku4l/2xbzqPASNBORXtKmgqe3dPh0JXG4KWVUhDfArn8HJSfXit9Ls
8sbiSCYABTwvtp71mNXplAvJMnXRiI73kn0FtR7uCMaH4iMFufOR/NfBzebBvYFt
ZTVD+PdxzGuMsVVpL1ggYOmNJcApaUK88fn0bVcGhSAIh4vmV6050Z+ediV2DMQ7
YHoDHtphcFnBaFIJViH5E6f0VMANmL90Wmrh3Pa8tqq7H9Qg4SGztVbE6tSLGn/L
JrswUSeh6Fpe3UZpEjq9KrJwHS2FQilhCYYTWiYKgZRYUJGhzkMwQhVAypCn5xFv
WTDiz91nLO40p8y387q1Vr/ZRRee/hIAdYLFn2wv+JzMBFao7nSzm959e0NZiAho
n1nXegP1I212NpkeN4vuCR9fdFt1PQhAe9WjcyTsKTuKu4yg+TWvTy43prWxzIKt
6J7IbZSkVWrLWzpfQCkLP2CqJZhRHHeeILcFbc9AgMsfD9D/CF9JaxszH5NA59nj
CF9zX4CXK6ZBQvXcsXnzShjiRkpGpIYJ1cOPrgu2MTbIQs2wuIzzgyfnh6cwbaUs
ouz/Lr5NxykgJ+tPd9Ra5RUz3mi6R/J4GFaxyxB73G61bEWHFNlCHWXg69QB3ws3
St5ulxqWKGmjb4/QpWgjBtTYIrg23b2EXVRt4VRKSthBusoqYwfjsfpyg1W2MTwR
XL8fEPtBGZP2mXR8jjFqWB/yiD08surE45Y2mOonQzeAxtNTaNOJV1yuu53R1akP
1QDXF8q2PX6U8W1B3z95uL8D5isfkPuVCZ2yiF0Rbqa0l9rpvrK+mA5yULU9cxdx
bNpEM7yZvO0FFgEl7yWCkHxZ4ueenZHxI8NhRv3RmW88uyFdCClHvvZxQ+IKoDus
Afi6iqiVxMcUK4YKr5uES0PbhfgVjoQk6wRWNgFvx3YSsy0pe1ZdEaDEju3CDgMg
ce3AyefYoh+jY/x8t16/n9QLlzB+Vvg17fidiCddh0Bhq4SJR0cfFnDv7uKELDe2
8dCeaF4TlQDVEjOlNCP8cgiYH9CZ3AGpDNvni96VxyP7Ton0J6kw8W1dNiRwYSsB
lTYutiyQRcYhwrjgfBhFs0GjYNWRCzV2b4MV5euEBm/VrbBJwPapRiDvQxUAwrAJ
16aqWjC0ZDmvle7BQqPTbwi6E8Y6hi0UaZTuArVGv/NS9pGA330QxiaFsvQUgOdD
3MHqxu63rkrXleAQxPCpEhJtrL6bzl+rsdUVTuN7q8s4y6WtbsIPjodDgxC/4b4e
OoK4uaGg5hLdJ4TkaBTOhplj4hKRmponX+jJbxLouLnwzOGAhZnbrM0fLoJNhkKh
spqMAON0gzz7b2W9v3uQ2FxnI2/tNZY3UBMS3QsVcwJeWvIBR8/bknMXDnX5G/15
aZkcHiCzf2o4v9ph4/VOVYNwKDtl4Fxa85Anr9f70oEYZ0z4ADfzCsLPXH2JD26U
ZF7n1EJmH/hwow3ODEENm+Gk+t//ME7em3Tm0ALoz/DM66H/GQPh61Qs6K2Kd/aY
STu9T+XUSBRLAKnkQHETsx58ZVAFb/56tj1TOlUexA3nQk+gYpfvWt15I32Hi6u1
+v+C3GiuvUb3H6lTRUtE92oe7dWDWJjpo6fKtOEtO0kLM1El5TRpHj1xZurJbs4s
1jrev74dHgARhQs4ZzMoO3C/Tw2y/mQB93/D+xetWRD2ltObFR18yKUSOSXTNwCb
QFraOXVKrF6pb7Mqh/8XK7i+S+IJM3b/yMPgUsFsHIDvjHUH5NTyl85Ndo8dbgbl
QmGk9UhjccbdbgpdmepDA8IbzQZfyPHRLNwZIWnxQOBt1ayIUPh3vdhclmhzyelK
ABC43Lr6Mex9R8Uoy9LpsdPVhphdmxdV+WT3gZ/Tojr/8ClZFPxMz3mV0KhOz7UF
rkfUv6ElhQh1U2hNjO1oPeQ03+fnHMT25m+ZcOTf72yt2Flk6Sqc/xOZ0i6eb4Dd
GITa2KpIK8CfxjK7mSryxB4auwviieua+Z4c67Wrp6yAkyO4gwKFIk5ypXEE+MKl
BiAA4OoWU/qpZVyMIcllQqC2QeZcz/4gVLO1USveJ8MFsyk4eT1iK1Vr7pJaFtZB
JqRgAfnYXKMDI3nHcGeXj9Ax2RQPVm7Iq3wWt+Ill5QOa8dapLsqFKwXs0LrvuY9
DGMTAIAZJnlaWBz6n3O2lD3LPHqCD1VLCGFrJ/Yb9Uaf9805qycR3FmD9SvtQYwT
Xe1xusZHhQl1W4q5+z5kCr4fJPkb2VJ0OPZVGApFRa8U6wdGcSKWGotI/ZMZyH2k
kehsaH2Sve/tz5dckmsW2ooW2vgGMighT3IPUjqlofVRtVC570HTmxg34GaZQcbX
fLyiSh9QWVEQ4IpzsG2ku18OrhPiWYYnQxPqeFpBSbySKtzQVpvxCAMx11SwI3Nh
rlLkOyR12Qy2h55B9OnP5NvKfkySRdEKTL2h4PLMzMo0vV4Ni0bCf069PlEwIM87
fWJKznbg8qAH6Uhb7DvXf4CvfLQXInPfSxHfmcqFK3D0SQWIqNYZLauoHbRYyLPi
0HpgikhIbEL1UvdmC43f2lCC4IMITx24pLrEKRIWzr2uJOdkR5cYRk6U+LUjH+9Y
AVCVgVh+TjstoV6d5x9ePZX/fkURSixHV9IsK5wYW0iv5Kc1i8VCAuq+3vlwkh+i
7yUCAghLCln/sHe6th4KTNfz5aw73FIz4LU0d8AUHqkUcvpWaJ4FjG81rn8DJbxH
hGERhC/x+dDr/7rfJa7sX/tIYCC41kG5fVOMDviXFCjyAjmXxhstXqwmsfsA8vzl
2QH/LOmM5p3nOr49GyoF46NcA4gxdZ/bZGt6kskI/H+AomGxVAL3Cr2db3CiUDBe
XpneUSRDnMdB4ATrElr9w0/uAIogrGWZC1pV1BaQTrbSvEhW6gNUET6G/n9V8dGR
P2XxbImFbd6eF4ln68LLXUAloTy9FUv78Dx7MKKCV4mVcpGkAwrjzLGqspYE0rbO
I0reQEdNVp/v4om8W/vo+EVvAHM/ZmQKCZScg6O7hLdonF/OeZCusfqweinAeAcR
+EvWLI1H/kOR3GPG34RSNx/6cUkaBWBca+9Y0Rzm5cC+JF6kL93NcA7iaJMVO64j
advmVKHIgc12UezchMaruOHQvAzZGu/y4+FyzLaICC4/g40wKjgukNSATCn573rH
yyn35pKrCGSiZ1CMMN47hxopXNXcHffljYHfFHCZK3NOSyvbFSTyFISWUbmUM4I7
IQ4i78Jmbmey851qqvzJvhB7/nbZhEjtdjvCqj4Io2uTMQCX0/7OLFlzpOka8/mt
ZWQnp6KljY3jbse3YmfhbIEGKRLvR74EAwtJK0Sb/d7QFxny4AUYrty2x3GB+pyO
obZojk5IFkXbAL+8JxLDmOYsiU9X3trITrYhMwsNJS3gozjtcmVXO1aWltlcZOEh
1lqA5h/r2XAsZl1dZmVvacIu6WXLravJ5EBsXY6vZfQwPYXQ8OYxSEfTuDetpAo7
ziZusIXFSxG9krU/N4KImtJCoePtz2Vt7w372wyzsKfi42gJ+V/yDSPi2GIw4ohy
zSYl4khc2s0MsbIv9dwKGviLZPKRsQUPsrIS8RMZTaTFYPYPCXOC89/XxKNfEhA0
AZiteHXiSr3cRyGBP0KiCh0GWSiDaCttwub+UdJNzOPHltYQ/S/kmnRQwxVYKz0g
Sbr/P1Yr/Eaupu5sAf6fj8I1bpuDN/mS4DLu/5CEOn7EPeFN+ikM4tU+wL3yRW6g
pMwtDP75sDjhQWmCGxBy8QVb/AuBIvoWmpTId30syV64p1IAgzYoYbAnIvMcrlLG
xqstMMOeOoyYFpLH5C5rbK/4GUwMph9rhG8vKytyvHpO1WaKBVC7DP8BzgikxGoM
xsW4lWlyOIsxruqhclW/sc/c0HWk6T2smqdVU4L1I9C6cipCJKlqLBe1nshI4dtS
i/2K3+3Ojy4q0btDi1EWDsRm2C4Q0bFpp8Zs5eJRAECrelJPxY22no1Z6dESghLm
mGsoa3BZo4gIHi3PlmQ4DtHXjYwzmfILbWpb76OZ2RIu6qZ4bnekYlDoQvCPgO6H
3CRiqFb79JV+JpSrEbKZEDr6vqXYyAWFPquja8mIe/zkFBq2O5jzNSfbmMIshZgr
Ra6eKXFpos9Adnvq8UBttaE1iBbTre98r/+9lT+xETMeYe/LUJ7ri+MJO10wqBQZ
Cj2cSAoQW10mrJAdCLWi30hBr/QYYBeERf+mEMM5Hi5y27AhF/Ap5Ecn1+9IOZhc
0ZPEktsN1lr01B7jRVPU+hi56hOQMY4Kzv/6rDo7k+FwGUFtUvkXgLLKw2pPdCui
b5bwbJYgPtRJGUEAbNvZW66nOguEFzXQp6zcGRjiOyWqVRn2o3M1XXICZ9SbIFEo
5vXEhYsq+fOC+mhZUwC+AQVNxqoVcrXxfQdVvIDTgSI+W6kBN8cf4xuwhluI292t
mXGTQ4FczDvbFyKNsnTTXQhCeqQxSzEqHgNwbyz/m+HEAj7F8abY2OCnGgZokH/s
9HUe1vZ7zvS+11OZ0q3MM78kcG4jv/EvwswMh49ptkNx2lY4VUDiKsIRQ3n9F8Hw
Lc3H+2KltyyX+sncqpZDw+trJ8zcoFkssB1oDaVY0rxaKCv2fVU84sJNv/6afXW5
UBroGOPH8sMtvcCoWYHrPgoQ0PFLzejtvOHvZ14VDz+2KVafznEPl5AlOL64Tj85
OThwHeEoMr/MdqUPP+5ZzMRe3LfMWZNBnhZzxkhVdjEnGjJ9l6vXaodpY+F7zLC+
bRM0W4VppnL073nTnKd+f+ChsdKwG6FW1lkYb8MeAC2U2PeSpqXdPtR+Z301e7Rv
Qm7G9/W3qWFUrPYCUguwyh0oaoVtRG65OrMcIvHa3dD04y5ISuOL9pKIkkuNl+hm
taBfuRIXSw4fALFgl8Ee/9qvcloVFsQyUl6+IZFR1BDh7hR37IGp2qwvn6aU5YOp
E+1da4IDWYbETQ7u+mQnlLxT3FpcYEuA7QZ8mXFbOy2fpwJsdqBdJkVXdoFo26XV
3rhAqqFzrr23PesJy/cyxAvdplf/w2cCXjEMv4WiYhM7XNxIRj6X1oxVqKqg7JiU
T61vm5EPE6FwLdw2c/YuQhI26RL7E3OpS6gP5aoAtl5lkAQodvR9ReZOPtTegfi/
2pp46OeKRKiYJO7W/TUHnj1goR0q1tJHuAsXrWTSWAIY+VBMsknoeLdN00I9NRQU
YaD8G5ptZ1rweNXuB4M9zm760JwzFrURMC23fWiFdD+9zB05DtcHJO+/pGwLHyZd
pO2+brJIDvFN/jvqLLgdPvxCkszu6wc+p0NZXPjjrI3WomBAIpxUVCK1iXydIGjl
0z3oIBwvMjvuMtq8nUoaIN/fis31XeGR3SONUi/CkbAPN5CbGEV/eReuGJ8lDCYH
hfzAuxqyrMpXYXl4J29RUBHBXXwrOY0JcTeoHkQR1deRKjEc83c51U1LXOL9pQyl
HuawqVEHM1b5CHku55uBP4dqXI4H0WkDScifXjrFKrRHAWXdN5kr6daLbCk//AnR
UNsNnpfZH5XBC2yZ9pit/TDNWSEfvgoWh3T404y32dvy47gsOExG8UpUn5FBPxre
9Z0aYkHA5jARzmqqZc3lYJ8hDA+kpvQd47x4p02k69WrlZhIqqyu/9eqD4fE8Qxx
0oj635QQMi5A6HuDM0SswwNU2acJ74d2wXyJlAqajsJ56dh3ea9lPx7rMhSYn10y
ff+jSbnCWpQIi9QwPA3GqeJfpSH5xUIzJcPbCaS5xkY+ZsVS1oDor5+ljCA8JS40
R8aqH8PkkVlAeUCFZTxjjgfyetcANS03T6x4hyrVXcRDEVBTPerWvplD+T7iq4Iw
lDQa346seEwpbotHFKO7genCOTs3/PqrIyk+WrE44artffha26zNn6YT2NWUqyiq
2tl52rLWfbszhlrasgL84DOzCBwwDFrrd7Hp2q4unnGsRrh23keyr2kiMlzAmj7f
fjxWTsaM/d2fRQkGH1SrimrHGzmdq2rP4duNiB35T4IEhAyqfxDMcyCkV05naWpK
XhPvkb88yEaHYqZXoqVue3eoPVWZqygdYEEM5bMekd87F1aUQimxw1Yunk2fu0Rn
8oJC1mkPrGlUa/M/KiJLq3AmPKJAWk7peU1+m+p3nDO3Nze6mRZSWrmgXA9fOGoA
MFEJpw+vmTSgG6ZcGsoXe9UFoC6eBiEDKZoQoVFfOFXRYydPikK/1OwWaxOxadCs
Ygb76uvusQZIh48TRERG4Lh6dS18odFo+NJSkprFz19YFgqWDy/mG1+s8LWRVhCL
ru7bB229vgZMqDqTooROMg9UqeHnVdJleBCEC3lNpe5HWj5NXrCHiwSKV91+6/oK
VSNtPF5eUdufIAW+1av1eh0baIAZaoIx5EWG/fWB6o6H5OTrlcto25zjKUT05Lgz
4f3ve4ci8hkttLiQTg44Mwz0aBBYJBrm5EcAzz1y1AanfHtCyJOT3+EyoQEe7pXR
LdML5rB9F3LOcy0rAYFLy3fsp3j0ynQSm+2+X4rmUnJNXNgRpvysL5LfUc00IShx
TD3xXCxfB50s7JOTXFlSf/zXiGVh4073eswNUsaYxtKA0MR/2Elfw9lk+kEH5Q7O
Ya6GzG9TqFR+UXJufvEKntFurPU6Sbhmp1K9pOeLvSgoCbiibegXU9mwshz2VaBr
bLLGX7IvgtefaU72ExYfnunB5cubv88cVo3i5yvJeIMwctaQiQmlR11fMiSJosG5
7mscM5hxB+dTNQBc08/OXVJ2Vhp0p2+Kj/YtCwa9UvXUDGduGOM47/sC/PBUqXwO
Ubhn87ubgbYPub7Tqprx3Y2OTKzvn4xbDnH2YMeYAs7Apz5okrPajc5jaJ0VTGrS
mq+pbC7APRb3sHJmwV1mzSTplEpIG7L21+eB8eBFqf3+HOOcwiPhFJyth5lKOc4F
ItnemOlhvn8HOzLfoHSDDZzoV9joZPapPd2mL/XZMkLeCx6mPJ1LQw4WWnNxoWdG
vx+b6hB9D7dvmVZoOgXlLhJlym1jL+AlbK2qXFYf2t/bna/COrAQGCOSAkY9yRxk
pLI/24vbUYYrVy9U3jMWrlBDNMqz2SOySNc4e8ng7V2qMExElbmpL7/O2/dzUwR7
R33YHb43orkDmKwjWBkjqy0MUhwQD2J2n8/3sMTMkuG5vsW5OLwHulp39/BVjSOF
G2KetZObDwtH9aVr1pgm7su4oIyIU4Jd8UFsL1rIhO938ryaH0HthIkZCflYtO47
57nshdlESbG8wSEtn6Og1xMiumHXLHTm+T08g/VccI2qrf7FiVMf3U4nFyodZlWC
G6PPYBfpjHYB6wktlO5EwccJ6oeB2wBbxOxKTm2ajNfPnQXp9N57ZQV8AL7rXJlO
6hliBmWnUDD65UgnbogLB9fuqbVzcKHuSUgW1/SEjkrbFSPLk+ZXMsvna1KrF3CE
bILOBAqodrcapDGzfkVMPXcTEAwojFxaGAe0O8TscwDRM6XA9VvvOvn77IbffkrN
D3aEZEptva1TqbOaaP5MCBknLjTaxV4NJ4rZWCDFeJzgm/AI6lAoyuZIufkpaJdb
2so9XdxcrBtzQZmYpr6jps1H4tV/tx/LaWP01UjfIMJnCmU3QxRzFjdLyCuv56qP
4XjgKT8JycWf8d4QJaeByDTHHaBMmqHpD2HLH5ce4p3oS5FPbwnQoCvP28sH9LPL
z8mNeASWw/x/bmsYSVJlEJCoQfYYj7A8Vcgj7LYAmNTSgMldru19nNnUzov5DDFa
Kf3BpQu9G6RuD200cOaw9iC/mILjfGEmGcaQ+gjUJkrsmESYxbPe93FOkYU5ITW2
o+jYyafBYYuFRR7XIg+9TeVJMaUcBlJXwhGnlQckGig4J9Xjf6yZHj5V9LHxthpj
sOnnkYNQyG1yO9+fupcqu1ap0IBkhUX5SkyrYzTD9rIuIrBAA7uRycmhFnPqTZm9
N96R0FXiQME3xfHgHa93OYouVZ05xsaOYLPfNjOMeb9mNJ1Ds6E2VmIRUi5p8MU8
R2OYu/HHGU49/eZAaZn+N1Knd1L7aTMXBd+8toCES8LMIOP1NJbvP5llzeVPLQZN
0CscS4brano4C4d61Tl3vQBe67+QIBYlyiKtez/nKDTfePQiWA4bWy71DR2t+P1V
p7G8NQ9q+CRJxm/f+HyF+00EwXklfpvfdDXpT5d89sruD+wiUf3Aht0/oc02Dsqu
H9Fe/5SNI+9zhv9Eh/BtBkzl+fZnqAkhk2eWOHaqSGvPGzUqt/7CLNsBsvNvqCHH
p6yh9bHI91g4/KmaEb8yrJ8fXlXUtP4xICJTLAgpPEifXI7a3ELTNQj/Jd5Vzabe
P3IsTynMYHu9zHtjZnEGKR6ySWfnPqr5IZxwn2TzpL1HEBCSkb7mY/KwihJqVjoe
+qF/R03EyrCAQFiRTOsIBWMHwU6PjldIA9nLmz1wDxK6UUo1F0GZaM1ein9RmfRq
W4TD/q+++4Tyn7maU9c+GDTcGsInVmJnmbNZQx/iDxg6avPG2WFd8aeQgKidDAh4
acu19L0fvqBhXTeSaparvLe2kn6uGIYBxXH+X3aP8XEjidGXXDJDno66NKdIeDiY
UcwI+keYLoHNfpbckil8PpuwSAHegreniV89qEp6z9XtlpFYuQCrplJONGuo0azA
5GKW3ZI6BqJwBpVGevRCxV7RN3yedOWj2H9xIDgY37/0+sH/al0TU4A9v+IYpIEX
AGoG020t/rqxuCWFy9BLVpSd9ofOlvFxWIoaTnbJw2HoH6YaxzPNOcHMnlfOh25T
EJzRcZXJkXz3n8OLmNHs4PaDKM9+krDpXrZNmXfklFvOuUVRuayauUT0CpbwznQe
VOAYYcQriHyLI7i3BYrQRmcGKsULvav5dk04I4BhTcWuqtqyTDKiwFSkdBj2dfrr
bdci5PKcVDQntHPNsssrO10BA/i4PoA+rI1q3k8Gq1g6gtLt/+cIUzBJWvuc0rkH
a6pvf334ekIX0GIaEqZZRNCT2QQwIt7o9U1Ku5TR3rpFUeNtzvNoGzsAvIA1AKLu
hJ4pEU1Ft3Ts305DCCuBc5Cg1bebOY3kF3KFpCfvIfS/9VnWAGKLyz0vxU2or/Lz
F+jZ5Le1sQyEvo1MWoHrVzScQJANINb8UfThBqwNJfOi63mU3yRJZeOxmVzIkzKd
9thABlr2O8tGcEdd4s3Aii2dS2NSofZBIyIWyj79VCZIBuu7SLqdD+l4kyeU7Khe
7r9cFVnn4k5+dIEAWu+cowMpgIHIV+RKBRZqDIYGuyA=
`pragma protect end_protected
