// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:14 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PubN/eXUXWufpzBOOIG3EzCaoYoxK80qw9mSIHivG9FhPq/l7j+I2fJsKWinqkWQ
s4oVcUcgW3eJCN0sHUIXSP1ohbAH1Y9SXw3lT9vSegJeNYy3CNbmuO7XiPsgC0NQ
2irl/a35ZtqdkEHFYJjHQTX1cgroyKaRs2v497MVfJo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11728)
QisPgascAO6tJQCf4XkvCSUMoEvuCKSN9uVYEdl7mwSwVGwLH2JkfxPES8f/5RN8
mnOOAPgsSwVlc/KchUEs5PVhh/yNALzDMZH0ChhNuSBQNzGCYgr8Nxs+XN4tsn2p
X139yg7fB6n2gjNRbNx/Sva62WJaVhjAzZu/E+ZJ/1nDMv475I2ecgaaZFPPmlhv
p+TwEbGgcuE/ySQ84yn5buL5hNkOz3C3nHVrFWRfEB0j94BKzPaXekgb1yT4613A
uifwfFdj9nG10K7p83GfyyTbRnuD0rcvReykZxAxhfMqvd8uWnRwZEurrbbBcx/V
4g1LT2+HG1GKihk7PyssWgFtGhY/mZ/dq58aoU3DX9kyuq827imo7cqqDkSkJSGj
vv8pRt/b7D+Z2veIo6OzTK0rzN3YbDyVqzh9ZSKXpiS1WzVFeKufXZYk8kTtO+Qk
sNHvTeN/W6RnjvKaXSNVGxX2QKHm1dmivBPUrROxQl4zI4YTAm49G8kOi9iE8Ifc
sU4iD3LZNvUoMkL9trVaM5C4LGjr2KlpRFAQCRs1k9OgLB4tPRoQSjLJHkOtSCPO
LUrqNfYL8vL+wl+4mEzRClTPqbM9wzAcKGgWlkswHpYGtA8gcnEc0x+uaPVOPU1f
pmdWj/CBRCqbtW96G/aUfonXs/hQ5ra7HXJIF6Z6ijJ4I9q+2BYwP4ZUnGajiIVe
Gt1j7BX8AbZgQdQxuR2SwfFyETGja5/qMipnY+DzT5/9RwqYF/1zaaHrmQo3ALCR
0/xBUEUlF6nU8fuiXocSRtqhZSy6AU35BaaVSC0cdmzRaYK9v/bDDJeDP+w/rZ48
P5Oil3CrOEWrcyM5xmFQxoGKZikUy2kV/0ekvo9BZTcTR+6on82xF7Bg155c+5Jm
qKCgs+gJJn111hb68ANyM4tme71VSHHdo+KS4ly+KhQgozZtjRQAicgm2u1Tk0+K
b2qn13VZzwvoI+ET1o61UtCrQvS0aiyW7nOS63HtV0Rvv+NI6yI/nqbcKHYxCNkZ
fW7P2zjmD13c2Wk9qBgLZ2RG0l4XJHXEJM22qxM18A30Pv5tyZ3pvg3OM4gulWas
gsqUXAgnSmX2b39XGMXjNZElT6bWlD/3YDnXHf3cCX2NIEqg9w+N9x7BoeoW/WGp
XCuq1B7AB0voPZhU0IdJ04m/RmAt5lC/O0HGU07DzYTtqIYbBXKeKcM2iGBYQ7jo
g9FEoirrRxT2prTbdPp6PBvGKlNGQ+5cPPSV00HowbDaD5yohI2ggW9mrVCqmQtL
SqoO981p/8DQSK+BcRFMbpEGMaxvvT2pwAqXYO93wHmLkpg0rX12w9siWAK4pC2z
yRA/7ZpRUIIABc5Y2rJO1syxoeuTUk7mIBVYq9R2Uib3AWEkyhLbE1JkH8ao/l6N
1Wm13fYMtV5DpwyDL9PbHUdTbGq3xogxXAZUXOR1mfWHHKqATnHUpGx2SxY3/clA
aH3+muRKpzm4zu7vkYT8w9EmQ3zu5HRFTeXd1cAUuqwUguXp6/11RsDDgXLWyS8v
wKcyonzDdCCZwiDbnJb7+9ybSNb3hvklNm3By/7CuRkaeKDxxocWUVndhu5jDAYI
ASJ/6MtPbuy9y4B5aS51Y33bbGfd681YFpmHIfIdWW0F3kZsPBEna3hF71zhi3ol
VH/RLC/Uhd6G980Pi/DsflgeUlFBcKXq8bdm4DZDG5Raw2uY/DoRcrUrwu6jiQOo
cnZ7yNv2HHkN8OBSWYh9W5PFjX9VCpweqsCmSxfZrdvVXVWT7g4H9xKkeR4ZqJIS
UyuSj9MTGrIDalaG0mjIvEx4Jy5H/BvmRKp9PHJ2ZAgalO1cV7GKDIhnAEr3u3ME
GeQjJX+/c/bc5t7nn6WzPVQ8v3LNpSZMsMRHOuHgSCWOeY8Fmj6hO7sMy7G87p3s
L9hAc33voP4cJp/YcMb0Z6k0943qCkdme8ZJaQ7usAL3DwijZqLnDaZg/39HjjR6
cD1sww19iMYLd7Bu9Z2Y/slZYhy6XnFWna/XysXpiy27jebx8pe+VR3ydarav5WW
T8CyBAIIrdmbpl3gvx2ZUmfd0ADSJqJTuKfaLmTCP1aEFJFKSp1uoytsazqli+0x
STMNWLKzqOgIyYmMCo9t3KJrD9kM8Xw3LufON6gYfWGvMEksY/03WdgBGiaVHjJU
hZmZSL4kcTBXU1cm3v2P95yNm+bPcIn2FEgoVijah8rDq9c3SK9Rz/zvKY4kE6b1
qdYi8g132GJok8b8mO9/PuiKAq0zOU1yzOWUuzuh5ZBM3QkHnYT5MGYY+H9oOR2X
hrw/YKRs0kfaMgNQFrkbR3TwfoSMwr8u8Lq0ERgngtMDr10czYBDsaM1363pvEn4
yfi92MD2JtIuyoFfIQMCTnKfVEAPPXEVGRK9XTNIKe+jPu/5eNfhqipgFDCaK9gL
n9hmnezjbT7k7fsAuMJAsBrLAwUqpBARTWj9QGqMaCSFSgmlhKguKtah88cyj0f4
+CVljFhjWpH6ZV9CKQOaQm16ebpa83w4AjYPI4Mas4bg/TX80h3JMxNHllhuAtZy
WGOtzx5MZg6LuMLlMKv446D4yj5RBeKQ272wR6QxDFZvuFgKx4tQRAikLTZ0p7bd
dZP36sCU5Q4R+f/Srr2sjunC80Y28/sI3slVEAgHvHdLmM4dG2ZcRfnyE+E6X7xM
vqVncnFKKYs3voYPXN/qsKKnxluyFoIRTBl8h7wEAyEO8gFomqrdnzYy6pVjBrW3
4zzGrDkbMNV3cRBxQoC26uY2kD9CJF7arB+dY0EnsXTotsLRKiffuARF27HAxa7N
mnkc2Z+BdAb2U/xA17xudfYHNBW/Q30geykCG8dcFYaO6sXVRGcJPtsv3BMm1EOw
QXAD5wLjS/zxm4ZZShJ5LdU0DSChVpbTGZl+dsSP14B7RF/wK7S6GwGk0eoeUF2A
8OFtmZEQpb+/bCD+hra6MJXTMnve8qBUeKpclPpPrzn8jk+uIHsPyTDHhWPqZ757
/KNrGDubFgaS8jSRvdciF45eZQjH6Y31WAWpIyu3VdTSLN4zisC1h0kIhap6wqA2
eEqUoCSiCxSzRTtr9fVtHme76Mi5oSI9jY2QLwuFPpHhjRKoooqAUDYRcxBzcr9m
i5IKBoC1JSL3pfhgTMpZHLser81FV4UyIPpW6ZNWgpTk+/ZHeVlo3glqbu2VJsPw
lO/GpaU1HJ4K9bgjaXmnOZEN1JGfVrgO8oVxZVrEN8f4r51C6O/fBhWmr7mXstM0
EitFxNU2ap+v5fnGz1mdSy2e0u7VIAZ6N2l9wS47HvFuqyTDS0P67h4ZfC5FYh4T
SkcNSw6GjIw57ZyG2J6T6juiscT1Kl4P34DG1hD1N4gicYAGZmY61K2zfOV3uDao
hpVVk0KY8M5l1PqRk0XCYs9UKsL8F1LT5SyCJi12lC2DHm0+WGIGRzMrJhsCdVji
0nKfogqZoPuYi9nakV1hFBImmNUDHTyrnfsKI147u0j7wQA02pSFggsCgQbmcBAF
iRgGEd5MEroKFP66CSUS4+PxGqZMsFKgudWulH5obS7TJHE3MvxxLIabuk+0s+12
6cH5d9F5qDaGG5ohMgnCrxbPAnBI0Mo+jGb8X1izJAavSAs1HniMb+Ow8pbev1MP
AdIuoEAoWYjk6hB9mZ26fuZHYVTuhSvd1vOaV3kUA6SYhlV5heTBhHI/yfotTuke
z/jPx8/RkYtov6i7zXVOnp53H/c70NCC6YN+GZbOzdD4NFpFVoADwdKpMNvjslSs
Ha7+dHtxoErRwBFfndo1ZHdtUDRSMLplcQ+tv34kAWjxrSyVekvnwrk9LwmK9XCn
CCaIFsyfZlO4RFsXQLZX+V5k26xt8mfRXtydOPNYl7AhzNh+Ot5z5F9YXp79+7ug
RgU7l3xW5nwPQ7sJryGVN2KDyxDBBcB95wvv2kKUNc0+WOLaGDM5HRqidVQlbqNu
t38tY7HnYFUDjEWXVMZeyQJXXU+65P7MF3cnIjq+8UkD7OwaSh+c7nRFdb89PkD+
AwepOFyJb/LqOL+fwXTRb7JrmAl2PqpJXaTF3jTXwTgzISYrsjXHppC9gDZICOIP
MyD8L8CQLoCnWpvhZC2scObTR/GpWAYoZW+ZR3evWBVI8RAl1U+Ab+6/VEy5DIP7
NZYO1aNXF4QqEkc6bIvfTqDeJLP/QFtcZ+Az8T6QCJue+JApCqgogTm3Hl3M41hD
GRWKt6QK8CJ9wsCXZcgKWNpJ5X+LOhJZtRJPdjdJktZM5cUB1L0640F+eyyEQn5F
WvASuCLqmifo6Q+6sMBjss7J3qC6o7DGVGHFysLKWiSeY8gYnnau6oIJdqRehcH2
154+YeiJ03ACChbGWAHWuFsFwHqlDztV9dFUyOnGzx3G9WMS90xSwhXhquR8WzQS
ZEVQuOLwIk62+KgQrMGDQ6bgn8PBmyQkN2gpc3GNtpnAKbDH0HHD4D2yQbacn22m
382hy5gx7uEEZv7IjjqZGylEnp6bi8MgGj983WbiVmZOawkLTXuHyM95udOXf0Zo
C8l4H4zagzqlUjU8goyv08tcKCoAN5eRu1MQ5z1J1al14fPjV/1m1/lffgal0N+J
tqyhZlK2zj7nbYlwpUy4+zzip133A4KMafo/jAwc8p1CNWEXjoQkc9PHmYmfW8oq
Io+175OchJ3rkncg4ROMt+hZa7yB+ou1g68+gc3DWdfU8u61Da8Mt9OVDLljgo8o
4trACXf7teiuqM6opg1YeiYD99lNC2WcCobK0rYRJPZfrZ2FoSLU0ZQXs8H1oHif
/KXTYqEcVi+YHTmaKsYuJ/wiATyLmSM7mkrWETlVzn0PsCcm2ZYhX2aM/y4bIgzE
Ccg8pS+czZrrgVuxLAUug3uhvT5rggbMCRIZNpxcqt1OGfia6Wj/KInlam146mXa
xJ5Ua76dLgaf2oAbSVhpx+3IXpabl7MqJaG6cP2R0pSRAKabIKzAMtO+B0ZCDTiu
OLaQF51ACbFmH4l6DgTlpwt0urO3ofW6pnQCWWMZ3S7pyAFfUxnftXbwvrhfXDLz
plFy1DnYDI5wureUgYHY/3Xd3/JKmCN9aAEjrIXNPShrBdmUTM9tSwy1jEPO5eb/
E+RQYOA4hUclhdB/ifbwReFNoJkGYQ1OmKnvI9rYrnRc0nFOhPJymsB1rq/tAaEg
pOqIfpNE/60s7TZurRBExIyqPEgQklpvNZ7BSe9+rzVQh4wc7HxtStXzT/Y5wO97
dk7HyjE/4mC2Rh/tNH4q0a76hLqs953YjiEOZkXbXdFsqOZ6dBShbVEaCcusMjrq
NHwQfgmvGIfLxHrauYzfPjpddIrYerqsiYnvtT4RV6Mv3I0o8MUF9mk9P/k05Uez
7kjOqtGyForD7CjWfrq4nr5pgoSCjsEIiLcYxmuORMSyv8JjQbxuXwjwXL4TRE2N
aZ+gL5A6bnQFEgYEmWht8sVobb8fSPHD0A/Z52f+c9inJIFucj9+RRAGxorcnKAe
qnOW2pMt+acfh0UGq3aPudakjYAMfdufFLcObnkHVhEFz1Ag76k1vUR43nRSqb13
lAujfntJj9yI4Nvv8y0a1eZd5AugWxfnvfgaY/172cBMvLgAH7K7h5mZgAR3sohs
DGXIMrwqDH+vp0rKVxHt99aGn48Obfa+yAS0UpdcPwO/+WebOsLuJa15bZMrohsj
jY638bQbU42cYX+x8r8zLUQtOPJESlqFXkmj4dA6DgphN5xylG0We5cSm6mK0oEp
7c1FGLuj34gfUXEsGvrvU6T18cGHiK5slM7Bko6O52edGEezDgmBWtaa3dlZshy/
R5BF74VBLCK4x1gekj+iW53YcpuFPUfEMNVTULhdOcqVegvuPh2J/9gBCT7J2V9L
G0R+X9opUbjdabb0irCBiZ7pqnJPF2VGOY/WXhUnh9l/CZ1XYHPHJhsZl0EPYtEv
hmiqbNmdhOuuj/4fowcfcwbZBctqgNREtBXTnVy5EytOS+ohPBtRyMfZhB8g05Hh
9DPk8Ftuhy3AdVdbienHqrsOGNCrodmXJWAFld5EtEGruw3E/Uddlk00iVmj1tZM
WLLtPK9GucXthKThXx0Llr2zANdcmEp4zgYWI4YO/kgQ1Z558lAhaSjFGgWOPWAx
7KmAlusapLW65HOl+kVTwPfvbzDym9xWbVHFByCrh2/3iXhv3MXPnjXsrFQFEM0b
K1v5/2OGUqZ2DW7r7JO7MXyKCEF0n7ERs0olEHnUia++aUkW49jkqYZw7apXgCWI
LCFs4KX/3NynGDyIX2N5CPmXeeZ/p5aP/LBqx5bYHmzwbmzjJDg/4M7llexV462H
d2g5q0+vm+xP2Ff9lqbCDkbRDXgPEJQ1bRwS0qHfAXm86eh5vC4FMe5arYOIMIc+
ihiaJv2Emeg/6uVRsrnLn2uJQsZmubJYFKjIpP3UjxCthPx8ij1YWG1jPKJmXxjY
ba0Ye4aagdJ+M081ZbYxR1f34rl7Tg3aXtoUScjtNIky9k5Bk/p877SdTmJ3cUWS
Ngr6x6OdsZioKO4fORA/sxcxLAFjDS0w0IMlFOqHXOpfgsxFgTtTBV+78oxmV8Hv
ZsIit/OzOpsl5/iHoiEXerCvrZ3A+USmwrzt0xK2kA5nqfQCw0uVBUtiTLff5klh
7v0hqdJX+0TiDgEMVGJVB1FUTctNvF9xmN+T7D1RO9NzO5+cr3SxmgqeYiktsNec
Ly4st1dDz5oAKPW2ZUfjxCm0K/pKGzaUqNTyeBucpnhLuXnvEFZ0OF+fUKQG1OoV
CAUovYKlRbTcfT6mTyJylD+W+MVKMbXtXh5drGZ4QIoeve8Exowjr5dSf0ABc8GC
/qkAJkdCh73rlfq+3dh0TBnCw7NgG2hARu1hTjBjM8Gj7zgnCvy+qfOOgNCR/SdH
qy4nAcMuF3dq8stg0Omb0riXJDcxe98xCZ6Wthw6ZtCnpNtyOFshIsdXkn5HJxZ9
1RQvhIrjrknypGj9tTra6phSOe4lLne/AGOEkP3/6j52niCSra+mZLo/5/Z/0fpy
T99qwrEq83y/ZJfOkQmJjfBxRTP1Eed+i7yP0bD7gWkwePbi6Qq8fRgBQehxDsy8
UHGcsK1NvbJ8ahhkdtsv4YjulqbsTf3sVjrtk/4dPdNZ27Ih6F51gS35g26VjGMq
cftDDQ06/NOb6opvkMGoBoReLzlVtQ3hh1ZMu68m/21gSDNufsFWIhAFzCFi3v6K
80O4fdkzRUz9Fy5JIWpEh6BBJ8yXlqArS/5I2iiB0NsSIhOUHr2K6ihhNcYbpR61
QAtq7L8/DT7MA+S9ukvDaKoUTDs3EWRUHkOITNAO9HJRCzR9S2r9qe7MR9fgkMpo
b6i3N0l9oTf605xIy+a6vxZAS2CDN25J/imAah/ijsxpVcbWt+cNktZxmcyvEllK
E7Rn2nsX+Epjcdhh7sfczCUwDMVHIpt2HKO7BxtMVTgEz3Hyr6L5+oSkHb2x/rKV
3WVUmmg7mleuLpnu8Y6oZyeq1Ewf70zJo/t6yVqTZvN3vDA4cia9t/r0br+b/oT8
E3LvCqMvq/83UpOIsJnuMfg+rlZQzt0TY0LS1deX50iIZCnZ3F4a0naGDD6af6Qv
aW2IGJFfYj3XJjqfz/r5ETrVlT/SygVCsCMu8hChxyd7rLFz9V5bf5px5QSf4+vj
Zr23f8U0Qrbb3Cw04m742XGgLo4UaRcxIK1OerI9r/uUwDIR3Nk9CUgs7bChzOhE
CtMrKVJ9JhfiR5r6fd2dTagvnFfTxMI7h2kjsbCDbUE66VsWY4S5V2eziFm0136y
qWerMmhb4YJ2lnjnmC2n3okJkw+aXehnW3n0cVjmNdSFpH+pOOdc4ETMd6g5JbnB
jQZMoAX/xyqhMN8REyeHk95Hjlbw5Nil7LqwaZT2IT+9w2Mf4Wt1xVd1+uIl7TqK
3FjjU7fi8FUTRMITY2he7B7dM3rmGXm9kPlDlUVbLt8uAjK5Pajv/BM+ejoA52g3
CUzujc4iZNRrHrgd8F2Mullb6+X1xDirHbBdq3W15uG8bqndpZYcr7ouAroTbprz
GoG+6orxV5iYLxp4Yv6nadO2USH+EUYA7xfAnjj/2txdlBupjIIs6tBbs+y8mN7d
zdy6Vn1Pn2UKQ1AusGIZif+xKHwuo7WKQeLDh1do82SgmPz5wB/msDghHqkdTjOM
GAUEPoXEe6e0Zv3sttO/7FQEO0Hb99NTIJsBqwKQzRJ9ktZzDbTW11cOpPxwK4Hn
sLWDedFA0f0n+Zgq0PHi5tll8gyzEMa1F94DsPTG6bqt85p5LPUEfA8XlJZFvyVO
NMbZuaiFRWiTAvrIgbTg+OWy29/ps4YVLkISkrPHTRN0OlFG4bKJOgkI1GSRss4r
KgYY/ilpkUX9Pr4z7Flz67fJ0YRztZntMlflI48KCkDkQIdg9Rs2dhUook74O6tB
1YNtvugvbyR/W8v5uy78VFXHz+2z7Qv/AhKJu9zjpZ24XpvzSlFwb4WAZ+YxgFSr
RIujr1Fp3zt/ElLks1ZtyEtQBZTlQeW9Qm9ROLuk+3kvqWbMq/Nktm/MFy8C4bPl
M67hJ3aFJmfHtUKUNbRpliEsdgnoCEm7ugp/TfxIm/Aom98hTgZGIEBbX0w+WCqW
2EFBXHhcyKMuSeIZaXky0mJQOAqhs9xlklLX3Z3LFLniYBBT/YfdjvChddJ21jVC
V0dDzaXNvV4dS/6853RuP3pGzV+/y4MR4qkQQXj8AadK97fzquSVK5MX2qyi5eHl
CE4vUyD4YzjXP4eAFK5X+sISX3GCPiJCL+bLIwLYL2kVIawykwImrnHcPrOLv29B
3ItVhdw3GgO4qpngbbVSTWHtPMxrGJlXhgUci4Bq0Fh62/fb1FdK6/7mv97+Llv/
2zsxlLH2OTPeF1Upjt7Z87/yRXZBNgmRDoR5IEPrpb6ZN3AYgOOsGfMOqnudL9o2
lJyTIEiHQ5iImrYz6ZycAqSWY1QQPzLeTCIjllTSV0HX5Ho1KsHplAyIXc+jCENz
aG9esHiOKLTqHygB+4IpyZEq1FhBjcNPmXC1kX8N6hSHKp1chbI6fAY3ub+gLb+/
dGYcujYdRATHHsmtCUb9JQFFMpP7SBkK5X7NPA26QPcURwRPknL2wFaox72vAHzs
OYS+QAk//rpTiIcMKRTubSQvAAxSFiJRFv9vxiujFNc0R+UauXkZAgyyDQzbWoXj
RiLH2wr0jBjdLKDDH93Q1TWTerurdIzqCIXifekDM5DtX1UJ4cjW0W8ybXgTw0EC
9JrfEaBchTHu4RlSXh93/erwlauUjapHZJIkPPWI2E8GeH+og3rT8MrrbjC6JTlI
Ylmor/0hEO9a3i3VsTmwc9WdR2lCt9gbSFjUNO45o3mxjEZOHWCu8daUWLiT4Yh6
KCl6QHCp60rjiN5/Q50QB2iVJ0ZcieaUs4pJ5V5x0l+/pW7yQQpWrAhAurtB31Uu
5+qgRje+PAxFh9dyWo5tgHW0vZMB0116udQTyw1zt8gTwQycRDC/PVMXXONg9I1z
4HJSRmTlyU3vWNFZape/V2YoVNPgBNOobjzXkMFRjDY3U1G0JZXJUN4PCz9oXCc/
LZc/DDrTtmj9cpd+ff4mz2sN2ujXEuA7cKrdkEp81KgFLec+bodWsPK9+jwzvzek
PiZiUWFyA6qUjylWgTc/LbdBgnL2uQMzTLxTn4OaLsPRLDAu/Y8B+2ySwwoDgC9F
LzGyyVOgT08eY+c9Z8IwrpsdVH2ygMQ4PC3jmFVdiAioAn1rTOxKCKKTFnvPzSpI
6Yr0GTBHSHspbdrjEj5j6+BxE5t2uyTtCMY8GQzO6q1ibE8mmd4dpxhO8uo4j5aN
GTdVPPCBHpbarIfTCxcmlPUth0SMzMVi9n+COPxVPa+ZGAkRAKuMeN0Fsf/ewU8Y
TtVNF3yqRqJb3SVxYfaFgASaQ7qxVrXYr2zD9Ez2Rg53Xk/kYr/i+pax/i20eQNq
5Ldg9UTE1Sx5NCgb80ThDoFIgRzYQCu9oWSjcs9v2wAg5DF1y/9nC539VACzZOB6
yITG+p+mk/4NoUpBD/ALJhg8MU2H3iP1GcgSxGSw6Z/zKUNYRQcy0zD4A5MDNBBM
BekoMb32ncQqcYKxFqv2eDqm8qOiUxMaXUccFXei1xftrQsyi+QbrUHWoyP3MDD4
UVf71AsRTdAOXYHZJT+5KYm2jd2zp3XT1nqRoQH7tdZMQdH9FW0rSQwxCCgMx/U+
ZGOFI1r0IudUiCGFLKJIcX+4029YbBsiIuTDh9ehNHzkSkDnojzaix+a1Dhlkw+x
RBJ065a4LtC2OsMnlul8DfDaYcbM5XkiN/wfRYLtQJJRyrzNbrSFHdd6Jfwh2mgW
Ffyzt/JNw+1ERZFnPEifDypnoiaIkxVtoVcl3rWafQdQ9qeKyL2mwHpgu0GgrZU+
dpW+gyzt4IPbsH/JwDfPz0WSjihY3d5CcoYVlH1aCKM3634vWA5SLxiJ/Cr587mb
vZvXTBmtUde7ugZ/a6FHwG1cv2vCmsPP0aqhUHpvJPggbvLa3NtkqumrED+xe7Cx
7EoBZbxY29i1DQyxM2obAVswP/JLK+/q+eG7WMtV+cG8OE2sO/Ui4PV06DEp0cur
Elwdk+VOtzIxfNXRahcCuhi5LuznFoK2CR70AA2WLk80vR8MiJy5TMB9ni2aetEX
g7/b8RCXygAt0mQm+vA87v1HqSiIXENMkNec+AWh4zB1evRE0hzcXEoyeGWfQ76U
bY340vBlUsXKwaN+6zcwqQGZ/0AX4Zts0AGXi1YxxTttc89/TV886e3MoSVUjYQD
TE58XFVRDfrPh9ZeqcWBxdttaHtS661hqLfGP1HPxoKTS2Lb2r/SSGsAX2YUBoow
8cD4rgC6Qd2bgGU/UF8fl4G9FZIzl1yZGm6p556bmjy+IeHQymAw2lp2/AFd21pS
fISaiR/rhgZwzIwc6qd5vWuqIP5H3UgHbn7BW3n+He+exW4N/IwP8EvfVElBMS9N
4EJlvCBLR9D+9kT+QDfwnVpc1kdXRe2qkOpgZU5o/ZByeHbLuU0VS+02/aoIzaXS
UkUZILv/AEuchpe8030v7fX9e7R7JSUbg/nmlKU11EMkm5T5wYi5nlTFFM8AaabU
lM2KrzKs/bG1ywxNcsg8RvEEDIKUYtxoxakMSDXBAbvx21MPJPR94rtNx/eRjcc0
Y5IaVKTEISjLr2JnuVbOL5VIPYxIjo8sPBdP5ykBwUyK3YQewILGTcaMl4Ewwe9O
wtqDVSyj/73P9oCQW/OBgSYKFbBMpBNTP9CQ56cQ3+sWcfEnvotuPLQR6kubB57a
C+alfSVs2Yodcqr8wonalXzmJbRcUt1XxnUStqOXLIC2qJZjlOhdRUZRlGQyllW/
aX3R3m+2QMUsDGU0ERx/VfM3+QmltECPAGIeHnSMGK9NZEfyvNqU/e5mJTbhooXI
nth6K+ivyr6906Q5FMcaHKF6qjovlnwgC7POdbL8wplf9kwyC7xS7QFFYhuXWjYG
4UZ6vxC7QA0cjJOFuo1TIcuCdYBYcSXG9uVVDxajWmgZxeNEYfvVpfv0pUbQRY8l
DvTo3qrxcA802jOGz8ltwFJngwFfWoSyM6GWI+8dR5aOFCNvlmpS2o9FMFejj/sw
4DB4zlztDDY4drvx55P1QtdzPTYeb3yKQ6qvHVQg/muRr6AHwo9y4+eze/xDDWjN
/FeDv+gyqWvItRJS8Xoe+ECO+vP8OtLONG8Mer6RGN7rYO/uaT5h271/2UTgriix
5cG70RoOd40/cmgKe1WLVqUPNeRljPCuBeRwJYSh5tw9AjkRdsXe4EwK8U118fdA
MjJEjPzmSHwALQU3wBfqlZlr6ag4w5XfDhz4dpOhIwEld9TUW28SSDykQBOqGVR2
44U8xJcrfs7wO9LE1+d3zdnTzUL78Ic0Y18AtD/Yd+nTKKiFQM8YtcdH0w8n1uXV
zY3v4DfS1BPsT/9o1IDaL5Drt3XGqWnAFvD0apEFTZBWOFvsijvQtCMPjTramAyJ
Chdu7YireaDG5pPg96+o4M6fM4Ms25E3FdTH57ViJdYllA2J81lgm1spkuTfTIK2
IV5JVVtFWtW2Cjjbqjrs12isrNsrj2nJwFMsaFmWuKu34x4zT1X6atI0rBzG7F4m
2fmXNOrO+75WevI3/YATL6VItwCXiCNk3zccZLlqGnc7EtEYGXDLIjS+r41RuvIX
7JmIKgXUohFP6Mz+bM8PayPKkJEOBjgXiFyJ12FHKxcFMzKncqFR9IgUqvvdvipa
IlKjmDfKhYrBOK8DFD/DUJnxZzIqTip5C5TmO8OAve1d8Coef4maxsgH7iZOBsuO
s0seky8BC8YRGqcrlzxh2BoqMsSXws01eD29l2wbmhRX6HHpDsmdekweJXGM/snd
Jp7TMJwa+90nDbfrkZa/ncPpDXYasbXBgdqHMSw9U/11asypVpWdgZQBgq3NOZVF
Pi+CLxMi4xW9hinVKvEv2LXmYsCZd0ozLCRRKpE/TeVR0JmpKUc1DLtb6WAkrdkm
dDx7hp1OunzxtnXT59POz257W2o0Trzy1l82OIHnxV01UtoY5gqOR+zrZrRA/kd2
O6IEN1D4ifo+OgIlo/2HHoeHELCWvcZj2xbP+9+9oLzrNmDeDxikR1y+yqx9V1K+
F0ksQGYmdtzUdclPudqnUP31Ga/Vlk41aAGJZ9pjp2jDy010JB/h61ZXAF7JPJKH
jesRkbVvXybm0N2bCS4OTnA/NR5TUeMy/4do787qa4al9SmVn/dapZcqjH61R9go
I4s3RHQ8aek8bgpqL6IoERx/Rr3AUxpZbdx43uciIakXjUZHEBnHSCQ7GYllNvZ8
rCHBDI+hqRZAIz8wXVEtDgO9L94uCv/euPG5Do72NCUkAlxsOL7Mb+yHsb6HfyGl
SUMSWV1kae1aq5+KJQ6oxBnQQhHIyXjIgAD0CycBIKmJkwaiVkyQztSdRBotO4Ha
98ug0oXe7MG8THtlyzQ/y4pXs/dECfQxuUT9EN8onWtsZS6C3qC5odFQSzfP6Bb+
YFGZAcomjNvgFW8Mf8d8AUKwVIX5N8NhYQ8hxGXiqKcSSmNKefsIF8RnnF22HHRo
Trayy4BVl8PVfhhcSx0esoxQ88IUGFc3Nj2UgaKNYeMSdET3MqOZFcHeySFNZ5Ry
pHg2O0HM71QrlhoR3C3xtXAuw94sn+H1U09yZBLjlVGw1s3RNWKV08xXb6XroJnH
O+X4TcXaQSqsxunVArEI+qlFM7HtPSyGwpNqL/yDCy40+yX1lxDKiqgKHpxx6f5t
iWM5eWYYQm2vfgxgqpyctVhPpd6nOg9KL84uAmfzsjjNTqkXeBdFXHmzHqNDo1En
ocTw0F7xrAMK505RuBvLev4lAUeditAXbZrG3aVIXOvjSOm1+eLt3wryYub9SqjO
axQ6/R9ANU2xPyK88obRd/GZBj4G2Azh15QiOqFCil15ahfkhMC0/sbg0Vrme0LB
jIV3/bKAdsjcrnPHzO5EoBmajVfJBSN8tAvHLDpyb08TJeaYFxxD00fKwu6+xKeb
7n5iAYwENrcbxczyaK3JoNhbxAw3BNIy57UZyi3MMR/cIhQSlledeQsh/Gq61Tf8
5flIMZLCykIg50S6lPQ3uuenbi/HOqVFTmwlAb+0GS72hKYXKa4Yvxp1Q8JXPdQh
4trPcnCvVAsDlFkmQCsvKBKXFnl47wSJ836yzKDmvU6JpYagmlEiHsa7G+3ZxofZ
0EwpBn2xepzjV90yuYqPPWG3JRXHqOtJrwZMxLfB3FPDUceGZzqcIvo2CJ37NQrQ
INGBmynfcM0XmHApFR1rZBf/TD6l1WT1Wl5yDJZYDETvfGXP14Z5JzOFzVapnwId
SMecfJPyZ6zkgWdQQEZVscZWLTHmUu8Hrgh4IGTSqHP4fX/OvybZfyZzfFZpsvZQ
jmRQq49qBpq+WTC33dtScOdBQLFWkamkvj4YnT6Qgw7KqaD2r5mu3yYh61JdGZYL
ij4kke0V1NAAMK/3ES45FLa1uvHWAUhMze+tJgIm7GGzqisSvAqt/qz6xzC/qXY/
2CHVIzf1cWi5GeOm6ZNpe2ho7YQberKkav6wYDFyM/PACPopl7HSRMuk7X45xZte
aSwVJWOEvyg5eS4gx5Tm0Kt6sHJzLtb5/OAspwKbg1O2vLitRSnamz+N/+QDTTx2
E6fy+lh+ENxQU/P7g/6Ec+Ww+esiQAvWL8pQmbZl+s2dUP3p8FSiOarPPClUTYDP
/p3aKKQ45KzphRwXxiqFDFG/3/CreKlgMNjd0J4XZDJy/znbpvOJTtBFMbYyjGcg
P3E2i9P4YLtto9cifsrROIfMCIBIm6npU+r7iQUcrG/mQ4MaYD0ZQOzeQQet+q0Q
7kgHKMlznQgW8pTOGI91g8EfXwWMz3RXnsipY28gi5EuHyMApxhgdc4al/p6HvNV
te1O6w/CgQEAehFsKWVI/nzhdqJVvEw9DmfTOfWRO1BK0DwRpSiQhvKwfQLMPxZd
QjWSvraLjWD+NUxk5HqgsZfUyr5Wg1cyN5tumkvZPlQtkdXMSpBhxi4Sy9qKQHm+
Gw0kcsPI49OU7NtS698nweTll85/mEeI+5AYWV+uCIH/GOu2cV6ScaQki9Y+uv5K
OZMAvwx/8Lrp0qwi92Pi/mgQlXxwBVVr54j2w+/bHfeQhNhf9obE9YAffQ0ESguU
gVsHCeY0rp8/rK2fwhpbDbXOvcBdzrJfmdm10i92BCptTsjTYrUibUjIW+aLEpk3
DXYy1S1iBBSHijBr/L2VjU4r8b/O1ZiXY9yKAxRWrfqKmU7ndw5LWoFqxV/FkasL
lvvTOjes+KjZJ3r6RJ335DyjzlOcACIz4Tlq/axJYl1ms08UHxRNKtTRNTIANRnA
dyC2YpU9OoKU3sdcJUKdCWRvirbgmw4hN8W35lIWwK4Qj2hRcTsiSF1lRxKkWbek
E0upCkd5XHgKn8ZgI50JpyZZMNmfZSDfKyWruSRSktbcXVnQadMj6kL8UI1PEOEQ
womSF4gLf427/jHqoFpBZQXTXFxbUfTChjXufA+iZXT46mYk1WIVGyBE+IpkbhpG
u84dKd8ueWiCclKHxkm5wwmcJ1dMNvsq7tCPrlsa+ea6pRjMvzWgTIDVO2VdluGv
aEy9XQlrBBUP07pKB29Kn/cn4BXJHMU20KHX0RsGihAwLI0ZTRfXM6dAI8rmS1Li
ZEqKaSFerJmRTYTQzu1mT8VMosxTZ3I24hgfDewcMz8wwHEgTbFxV9iWpJjsLvUB
rY3UzRmZuMWYUhBgCm/TcJ1FN/bkKVBp9GRrA4RqI8qqvfYCbDZpWGOoIIeR0NPw
LPZWAxfgTClw++expCcu4pD1v246LEvCoiCpSjcSw643yT0LQ7p8Lt9axNivCVmF
BfAsGL2/q1qyNz8cP71MZdd9TKwWH8S5XNOgvLWCqokdfyQZj2oZIvr5SljFhs40
aMSdN6q8eYt83qHHRdN0qFGq9YbKUcEsGngGVAcu8EAFRD7CEKDhXIDEgtUr67dO
K6spPfvNN+r4A2Nl6YwlBSUNtMU9Bwnjy5HQ8IGWg+d6eQrcV/Ql8G8ZVYkUEVFz
7R2DWj3DMucKyP4pXcU7mw==
`pragma protect end_protected
