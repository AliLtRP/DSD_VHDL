// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:52 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
j+2PEq+fAO5s1+l/U5L/m/wTz9xsLnUBq1Y5y5doP3DfEBMlwSUjH8ula7WDJDVX
idFiA4X26YjrNpfIKUoK/8Sz29t804SoeMUJerb9vBWWRat3CD/AoBUSwsA1oWxM
VD92q5f6SBN4+JOyPqJAeuIwnrKxxk5WKrUHCY7oJ6s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4464)
AxD6JEW3z0GE4906hk80YlJnJZn43gpQybgphIGnNA8+3UTlTszWuREB4HZZklgn
rTSqT75duX/XqwMT4t3uB5nPUHxOhLYDSW+7MpufrjjRDGk594w+SYkNaV7umjLr
qaZnw6qvW6PO5HoMk5YP3ERzyyyYwgBS65VIMGeCQ8FYMiCPdv7RKTM6Q9XosZNM
I7NgEjIkqHt+/gHWvkRa5LmGMjbHokIXySRunEBABNbXLQCQQxt+2/IoD3+EfrUz
UtckmX5m8nZh1n6NEH55ie3EPM64ddFmUoY7DPGNAgjyp4H49xuY6G1L99lkx0iw
8+5pUlPQ/Bm0zy7bFrvjRGohG+YuPvcQ8yTkcBZqSbxQgzP48IS2rUfAaqbNWaQ0
MDy40ZymQeNkwxLE6TKn8bQRrfnGYLCQVNAhwWqSkQ2AbW3QJ+BFqbMusrg+X/ni
LtYkIgX7FXaq1FsAF8NssRsmQlO+9o+oRJzWqNdj7Du3CNba0H7Wxe10vlxbH1Bs
wdUExrpi+yHGzduNZo6bcV5AH9Rb9P0J0edd3yIxs/PRIT0i40b+eGUiZtAA7jTV
SMVSC9+jh/mU2UNZmrKaxB/VILD9yckJ2/sOuD1CNdV/VrTESeYLQ4kTW8O0PQd9
eQORxVMVNwv7vsOa4QlWQ4D+ymGH3REM+jq7cO4JFnAEonnDnbMWTbMMLOJLgQ3n
3pdq1juYA6fRX3HA+oZcW+FCpBhS8RPJxLp1ltu/0b1xrbfOFVPSXfuvfqeX5JFS
+gh27szYE5zau/OygSwzkzoBeUq5Z1tLagFo+E9SWqmkAiKXKBMwVF5Z5cdx40kl
HRc5GwgXjwgIQJlbHZEDcSsj59DSqxAWjUydn9Yc5cyEpClxolqGo0XlAWeF4oK9
6tR4U6PjeQJvKMoo6xeL9tyCV35zpdUuOaeAhZ7vKxfKsm/+VqoYO2UIQ+1c++FS
96dTKulEG4XNWB8B4Bgc0gKjr8QqSXhFReNNGRAc4RAlBbs7Sdwm472uDemev1C+
ENokU04t79PmOfPdxY1xo0JK28mzAzjiJiZ3pwQsVLiX+ZPqasrf/MtRfUi+2lbi
UPN3Nes3W0IH0N+V40FDdbv87h+xYpXYFoXIucDEo9USSYOh3NwcmFgScCVqAS4L
GoDPmHsnmnAnzc+jma+hvLyH2dYR1oZYqpibi2/4oIPtxNSKtuybpj28XF9/XzF0
8FHi9PpMIHWsx19bZf2YAVMl779jF6SiLTtaIjDZznWWw+uIyLmohE/AxxR8rPzt
DwCe/CTwO8b+Tv5koA8JnicOuEmJ0QE3ZZ//3dZVFm8vwgFgmkga3WOmfEHNIlBS
rivlOb+9/ydkW8qyXJ3y3aIyDhakMt/W2NWxBhcOuBBF+im+fAFEuauB9xWoq/RA
xXLYrnO8Q6gIetCzmOqJKr1ZswRJXMxYPe7P6uNQ2qXPsoXA+mANYUzbW9VbYPvv
5f8asI5lZ9mVU10yUDAQGxspKasRfwJJrR6SLS30I7/o7mi+xexaPsm5iJgua3WC
Jzi4QqqLX1zPo15XwP8QlB41zCosF2wIkNM3ZHpBzPITC3uDtkrLh3d+aUgrX/oo
t0B1j6SZnj9D1+2UmJOzF+GldXH3m0C80FEn4wItaiyplADrKUEmlZdBSdQpeFT8
i57pZ1yLqIHzE4k39LYtmxmIh4ogqZLeGOS4zWJvBDPnR80ekq9Kn+B7F+obSmfS
dDzRHUKiTsTgabKwoHbX/1VX/oDd3ErDIUYajZ1vEgy4mfFxXS6YBM1o95gCALLj
lzaVjT9Ts/NUkOav+D08ToebudEhdQ4/TLULpfnIu0j5QyWOFxo6p09qB1aqlL9m
fDuvS4jEaKzKxejTjw9yXg/sA1VMZMOcfkUD9Jm3SibQN9OMV8C8FmQJQ8nrPyLF
XXBp2bz4SB1PMi765COCgeHEjbDmCzQ3rDOP3CaKziG+J7lxFI5n3QKJ98NwBlWx
ym+/TTrV1dtJuRSc8XYMHwv7COsPhJfyXpVbGmQCeE7IIZx0bF+LAKHg50obXeuo
n9BUiIrWpyZGi9jKZjUgDlnFxKgF1WcuBT5obaqhpW52rH/pHgjBfZkk26t7TB1a
4pLEPrSJFpzcqVEM2kRLgkfMhhAobL5SSfqNRJH4lKzpAnWVmjOGTipJ3ExWJnIi
zlosR6YLn5Hu7xSWc3vi++IeqVfKdy3Bxvg8LWZ/AjHRZA7m74kYGherdlchgpxg
x3joENeH60Qua1c4XTKpgoAtjgltnm+p0/7uyMyRXbUFMKyerUgWD6nMMJnJph/t
lrkoG6pGTW5b8qry699W3VuodeL2pyS9Cqwgy0VxH+9WBPMr4ka1loxdnjmvfKjB
7gscNXD1cnoN80VtRAIntWiRXuf7YznaIOtgEnV6KM8fxFcDkr2pgQTHzaCDwoW7
kFFDxSO/ZfERvApISJiyRbJC4VP2MHsRarK+pHE8xsBegX0KznTfBmf5vP/mzggr
hyuuCPCFZsb4x+0wTxpsskVpLlR1H3qetJMkAajCbIXhHudc0Znf62TKCDU3yjn5
vGmUJLojU7zx5gdMJDxt+eSpXUhA/jxsB2ZGnIBEk7eBLauWCEAwDjufhT3S14Y0
CaL5xiAeXeYgdTYYI0ai4YGQIqh022Hi8F1mDv+hWUJBbvZby/shZH2W4kXRI1PG
dv7h0j3Ld84g62eMvHxIZyizyC9RIi3DWDTCM+6Q4CxZ9gnEoA30BmHhdPgVDI1/
+kqHdW+M/AxU5IHk7dPINA6cng2cOnUIbuJMucUCayMRY/KXXdS4opus0Hy6Zu1N
9nrqLU3yJeR1qklg+yQqdRR2kyfEm3jZmUEzCuGaYjsVIX5z26g3BLlnLHF19UZd
8HcC3dBguiXfYWZM9DcFbjotHnQBr49Bx1Id9I31pYbNWMtAtuIyYz/s8zlCLgJO
pNnMSwB2UX/dOcg8Dld8nRa/uEYYhMwPBR5QrJbIzU7u9NOWS2PiBYWhKMEDFcIF
XzNLNDRBxlSJKgnXGAJ02sGDT3fzx0RozcSyuTMfp9m9l5vJQX9aJhpssR/L6+NT
koPjZxgyeSTM8thd6oa9h6cSFWw1sHe1MONTc9ttH1NM3+/9kDAzJgFzNAkfWQ8m
zLRb9QXuYB7mdRbvm+H1fjzV10MAZp5V0NKIZVDp1+DcqAvB/bVcRFWkZGBYTAGo
usWbN+2dx6j8LKEWkBLpbKTA8BYXqwO63zsDluNwgY4wKqmPWDEbao9yZd/zge80
QfKH3hx/nmU+4KMyDPiTeUydD2X4y931H5D99+YmgYdGEXwD8iCUBeHoGdC+KNTR
UgkdMKUZcwC4yyPkNPZTpQnvgzAeBSsvIBj0VARDkjCsrVELDtgpE4rr4BYomsLu
JPwZgGTXWr981HSofWtbijl1Z4C9kXTrrPg5SEJKGlufT+eaAYeA6sm3DaNdekyq
e+uxws9mNTY6KgBEX+EdJV9GN8rphs0+QeIIJvmpZoTO8lfqd3tQlGwbo+XYuHMu
8gTJmWqUz4EvBuVqC+UTAcKxSENRmzH4VzwyvDrMWcVHokxcXEadqQyc6Wtwlho6
sXkZsOMg7QZ1rxN3Xi3io2ZCFRppbLzcK36n3EwHdjON1ili88+vTBBfmUyV5Pt9
/d37Wi4nsqeYsjjQgP+Pra0nkxutY7xxLgGsWsrDZN+IevZRYiFcleXGX6vLSUJ1
R1Zp/Okz4OrdbwQ7b4ZPA3ZHGH+nHAZuQOtM/5UB4Srx4Wr8KczJ5n37WdYHrU0J
bBIf/NVgNO48fivAXWq4lDo8czmGGbyixuVeZ/jhUXcxDwSG6An/fC0Blo4vxf47
ssmhOD717gFjhV0xeeiRVVoI6IFJ3Ldu6GUaqcSCGW8Kf3u1t1t9ESJpbNaIQ/cQ
hcidhY6aUPyDYfpqU/NJKi2aRmmKYlSamBZyodoItpBkypK7M1/FhoogVkZ+FzR1
Nsky/808VLeKwlf/3y3xNcHconkw0TKUggqnAfgYW3V2oH9cCnE4Jx3PDMvfO9kA
qjhrPnQl2EeapxICDuM0R0t+StbDYUFeCp0NowFE2099G9SUq0kAfLnXyYp+8aXv
2Rv6jYSURmlIyjn55CqqQwfgB1rKp0IvOU8lH2uOCpO9mZHFFh+jfqTd5jnk72Ci
YRiV+8F8Am3JjYuwqr+JbyhN92cM4Dr7jPeoGvgRKOE8EYtdA/PC4fe4q8OAc4GM
hkFJKBZCttO/hPJr9mZ5QdZQTOKgx2vxva0Mm/gpcOZbZ3d5LAITeskQ5zgxDu2k
9BZZpd5FJXHpVa4oOiHPOY7F3tSokJxIwkHwsGt40dTAUIsZwWr9vUyZfHjaAx21
PgVlmU0opmqXay03bJzhYjp3sERIgRAoJUcMXyZ+6dTuz1jgp0UeBIeO9SNDxQ08
SyuBjy1aAdLulk0R7GE3W1FGkMXeLycPT8v5mgEdre50TuitQitB64G2z/Nw0a06
1nViFwI+v81OWIK6xh6K2AHcns00Tx83XBoug4zsbrJwgQhC4/O0vE1+ERr2f4Qk
oJ59KJRi83OmP8bRtZdBy+4tH7wX0Y6JQVuKa9Kykh76nDaiYQgNZcdy6f5dvlB0
U6mRHoM1kmY8fVqwdFyQS31tE77qwgFmYWsIjdk7TCdb8JSzXkK+zIriqsrwJfZn
8rxIV21SW43z/95viAqJ9y2oU+8iuvWNzn2Rex/ohSQUVlElOg1W8d941Ry8LAJ7
+GBpr46x/gn8ntturftkdaccLWX2/ClAX+JqYCihOt2PSim37P9m7FAKCp/kIxDY
pkOiULbxip8Qp2FCmiKFwMaSdGsZqf8gygzwgWJtA0O+xjWKGgZzAxyB00kIosxl
FoOXB7pMCcUecL/wOMF2JRO/kbwvH/Owab9+EaJVtNx+lfYlifP0OiLpip6Vw6uV
xmtxUfdQTptOapT0BwREvOI0DhVLfWOc5fo49eDBhtl0aVhSw1e5+XxW6bbKtEaL
wUqw8xmN4XQR2slgtrHlI06bzlBBisuLtJ4Ve1Ix/1TB26+gIXOhZ9PRfoQueEVD
98eb2cjRxX8JTaYVkOeI7okQaed2InK48TOIh8FxQeiFe42oVFR3OVKmSQyK9vd9
ignaKYgABd44+g09COb0AHovFeeUGaYUhLWuWUrDt0Qh4+PHptMm769+/ivuh5kq
L3gKOFCW7Ym1qHKWabb1U2PFRq8LBpGGxJ9jJkwqPNQk0MIyKQ/CATRcZxsCkdXi
hZb+mvMEHktYTFHxMPt7dHCJohYOhwtJ2OB0QBal34beJLk85cpePlly/AoETUas
Zk0gKB1r6Az9XGJcCbA7eFrtRBJlnMrjWrMSbh4dAvspbcjBiaxP9nZNPpiDqpUU
CBHpomsVN5/oM7bTSC46GVddWqX+TtROr05/PKbyOwQk5GSRSUDs/DVQ2vhW16S8
CKxaNudbsVjAuk+tlTsZu+giMQq+sro1aUPoVdMEDZ4v+E8cC8XuHu6byXrTJmwJ
3FielonwpWNffyJH69e+CXss8UjF7+NeqGlhje8dagP9/duwohzJ+Y55s7vkC960
3YLOt7vtwTdA0P9ImEownmJuyYa4V3x73Ry4cgnw38xPS2Caz+AJHhHPgXVitm1a
M8LOBEM8hnygGCLWlEJA75PTvvSJxtWmgjGYe6N08pacyUFO44oLSVoNZanLolQr
VqqiYwt0IZOWIp/5TVDA77JM813H3JOCeAezeey+6wVgKvPfcQvdo9Hu947W7Z4r
uC05LdilqF0R9zHvFn6emqN5z0h4531k17U2M59ZGp38moTQafjuw4NCBrf5gYSD
ax1Kqt3pmpNePFS+cQ9mLDQWuMqzWhuUFanm+8QRGJZG9yhrimqUdag7HS9DiHRh
tk3IO+jHyhLJOf1WvoPqgYlB7ro7AkS66dBwMlXmRVV0P5MP/6TSdBqnkOtrbSd3
`pragma protect end_protected
