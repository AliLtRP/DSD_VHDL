// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
GE8fC18qRBGwPdjFT3sv7OCo5fD/jztPB5wUd34a0K4G0wjQzm0Jq3NH6SgEeEmVBOHmyDxpxm9B
8sWZjWQ0ibfFhzF6Cykq1x+ISBFkKb+zo0liA+meaw+vd/wSWhhiNujScN4WKXN9jcI76IzE/cjc
o0AZNEeIpheEx7bVz6q8VsSPeyEuFM8o/LbBkpWmfU/fB/PUpwQ1T8VNtMNsGOfJkpQrooQ/QHYB
jLRxRHv31dwaCoFuy70mkPjgROTuEwl03mU/69dLYt0AVruQWMhNIkn8EdmQF59kQ6qITHq/ROea
UxEUZb3oOUT1XcCYqD13M3DF4X4bre8/I9LQww==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
Z2LZFBa2KKbrcpZ9/Cw90WbKrAviXQumyq5n753gi2lBGm63l39TJ0UrfUfFM2MQMTqnmjR2DUKP
s6LY4xAMXRuT9Yn4vD9wxY9YS6ZVV4myhlSdGoFuLeQ4uJFpEGk2TlASCiY1f5uASCAfFOT2B7pu
C/RpNFxYs/I55+lF3WqjmtmQqq3woC30reoN5H0TPPR+K8tdIawYG9vX/ppgUWkWso6v5p6FJrxn
axHRoXY+bmQdE6Rlmrj4NLbXnLmhkaG1q+4keKi9CzKwYC+6PRvG/o8QACEdybSi7EJ3x0bgQwT4
7oQSE/cCS+1DZBuECwxoz1jUfQSM/yr3+vLJSVaRobGODkorvFHoaUsT+nIPPr8cypPH08aSHIUy
JIMn9yz95FLdPxmJjZ1i+93Pi4gffdKOV6kbgdf0VyRipD4OIJ3t6qNzMgslX+SXfV7HqP6uvGGi
CQIJhrPodG63tWhGjiSYq56C3QREj13alQJrtUI5q12cgZBcLURGJBY3l2n7Gbq1jhi5Wi1UyhA8
pShQbwbP0TI4g1OyPg2rRsjZEYh3W6CDYOynMYV8fyx69V0/VOMU1tB3leaG5tjJ056GSSZv1sKE
6gr7iEBL5diLwkpD6AYIAf58zs5g/CtxUUB0i1RFQSM5kXH7KSN7U7FxxhOcZQBIh/vH1SoMz1NT
8LKfgxQSE0D5j+5qNjrvMQtHBzStA1q7d8mwG7IoFUvl+OvQOQwUxQEpT1J8LqPyrd92aiz5RR3x
7In1VWRgzQJRjBoOX+Zphjkh+Pp+Ds5v3ISYUUQxI+wAHDH8cOr5QviLFSvSCIpccM5NrlXAredI
CWLWHR4FIOkEvng1HOmAFGkXmxXjaQeF5xbHlLQChIHNhcuXTCzi4RozRXR4f3DpF6OLRkqPH1Mv
NOYkBWxO58ZHlf2kQaPc/l/YsRWkpoBOiArCi/hm45QA3YJPfq1KZ+06YoX8Ouj/bH4gZFlFiLJN
O/kEMxxP+5v7Zg7JBOQTR4Q3fP2/j2LVwmT2IXUYAKHhDJjsMY3uOJYR/26lolaeSZWnHO4xnneX
i3B6tCXVncq3fmtVgscYm1P3Zh+RrleTlA1xPi5k/P9E3QZoM0ZthA4fWdtebQRbwJi1wR3Ss2Uw
+3jZYCPrrMLIkp66oiWgzEMK93cMZS0KZtzWCWaP1xcf3Dn4DiCdEgpjYNlfpjWBYDzlRixZDOTe
2H2IfIuCbnQoFXPrJVNj4tDx7ARYYBbF5m+cdCInXhgkCNQe6hNbpZremLj3f8PIaoro5bsr35YI
TO6v+gRUtDEVxXC0xwJ32KxRZ4P9DFyYtt1LfQNeG8a0NoGZV+CD/9QrOd/B09iW8URa/WrE5yuD
B6WPsJuFSJ6kfNTYfiEDbLZtWEQNodnGqWFFaQVsFEejGIe6793EeZPUgsNFxZJUVOwxTYOTKKEN
WLrHV90/ysCyWbK4c2uZDYh06GBaGlKfYOAGZrKzYdM7LpwwqVVP5PKvGDokAU9nitAReTpWZHBQ
E9EeGF2R1YLDe6t9BQ8C30L8uTS6PTNGk9hXgSyPLYC0gIq5O7ob31CLwbyP1OrEBC8o67Ypo5Rf
7BqxTcHJN3hS/VXvPTWEbQYAwyRpFuBsbLMFLSuji0SBx88ai1zOcYBWvjnmsK/oTbkInJqzvTEy
lXZ0s8AzafOuJ9+jqL3xGWELyQimQd91eNU7FUdjDOJ15TUMWQCL8Q/Po+06uIUl5KSm80zEKnzh
Ntbn6pjsfU6xm/p8faUVfQ0KBLQZZ1XeyZlvxD9h209eB6l0pzLdLcBcRDQgGTas3BYOBNAQ2bmp
akWfkJHji1tg4l1H0TYfgT+Q5PQ2j8ARyRLl0BzVLoIaOR/YmVcN5Z7oL7bbtj5jLYJWqknSN6pp
4YyspiSH8hw1WqWS/hCe6WRfd+oq1KAkk1McgHlEDRP1j8jZEJcVVie2Mef961qURNqkhvyLf2pX
xmsY6tWgxYpQtq7ImCsP2iDWP5kxRs0UTuTYK4l8h+/chWD4N/wkF5jdHABvho0oTDJF2kc7Bwh6
4vbMsXQajhGKWTInhe+B9qshW3sdh3/iYhNTuCHxYw2EubPsQgwtpwXYnRkaWZ5IZI0/yERt1DZe
Tkc+GF0UnpeBsIqAdvE+4tM23d1GXo6QaYlO4spqBet6m1AE37c+9clhqJE95gbqKCu6CBUNQa8s
4KQQiSc8VPJF0MmEE5gblMOMA5mat5P+j2c1RtKmiC5q2MGaWEIcZxnEh/QnK6v559dsBZ2FSiqt
m5x54I7kplY4f0gzrFk2IwjpE3L5nhVN8kkdQUe1VvEU3G7iExta/+dO8mj5S8PRF1r9whh+To80
b/AECfhmsOZqNBGkvanNBAozwSFgZURc/Fxs6SWVS191NicRArdFiIaJr+BbGiNFfQoaoApRPH09
pEMcfIYSfpQdVTIK4cXXIih6MMhUFhvibUNQDvU3wIYGxz8MutiiZMIH9iTlA4pCBcjUkhDSOPCV
vBSPlvHASHsKAZ1R+uq6752b2r0afa1nGuhvMHfs6hm/2I2kTIq91aetQrZp0kGKW0QP8/zhQsXz
AYLYMSvYvZX9aWOepKhwWuAI9UlfU/WVrlU0JvXBUHgcU5wutxMExUNA6UXKB7+CE7YV/i1tuy0O
X1E0CDPp/Qxx0aO/jJ+WK1fciiwN9ispEn3+qkV8L9hChleH09XAtpkFMmcU64jKO2+oOxyot9TS
mEJq22twuEMIW0zh4/6DnCREHYZdC7e7BH5a/avPPgXKaChl4v1f3wmoWC6rdK66DP6glxCRBET5
dEZZQab3GJTld5qv/mky2CqUjC5A5o4u7ytmj9IwJQRKNAkOxYBEdPa95KA6TIpGOkq9tUVdXmET
hvppzxmjeF24Rcbb/g272XipnR3XpbtfBj+o48kq/9W7EWKdLo/s9Yu6TNBLWw3Kikvi2qg/Z/vA
u2U59OPX3TtB5tCsBEVpXc5V0M15xo441mKfZcgYNtbHDD2up0WOu0Yt4Y1ZFYkdkjbpGTbmbf7n
+DsY5TkxejMettKftNRVipaWwboRtAWiiCdNEFMOXkFDyBUjP/rHlizRu4/POgZ1yBhvUAocS4IP
3GEhll5+BbfJqa5fdXw7AYXQsu6t5e1l3IIol61y6loBrc3X+LPMQfccUe26ueyTpwOHKM+5be2/
afEMRIAU3mJG0d3+B7lFwiNIkKKiucK9d6oOUBnVUY+jtWGNb3vCjVicM0fzaw4N26A3QAFJfWWQ
sHh1pxza2RXW1VUPVgyCrGfpZ6KMOljP0k7qLWE5xrRZa460cYWSXlOSJwiHIYV/NAcCkiXMyEDX
83krR8P6yl2+HJizaYZIorpJ2W+gmMrzoyt7FnAH1m7s0vYjO6dIyJY9Ij6UrpP0kAGFprzE63IK
+QpvMLMhn5OwAMBlwcqlIU+H0OP40/sBlyM/EHluL1rImZ1eIy/6iQ1A6LAy1QKwC2O4n9fEyWeM
270xJPz95naY2jockkUw0u9w+0nuj4KkV0FErvBUd4EXYV8wqjNkfDs9Z852rm/T5t4kcfMJy7fe
+brzbw6iq61W0DBNOb6vo9M2iBj9uFqYnHKwb5a66DKLoPyZZck0c2mGXUNjgROVcswKja/mq9ZI
2V8KtFBElS0YE1AseCGlugbdKoqDR2ehEW37BZwU55coB0iWMrnxztaPfAxxAE1AJeGI+66RiZE+
42KYPTyMIEaTjg+gHE/cRGZi4VkQumaK61IGROicoqwqdr0igzcQ9AhJJ+jkId8NLVN2X7LzWSRK
KYnX8qhtX4MOZwq5QHmetIBQTAcLMimAe8ithXTYWIMxFalBSWc5yXZVY5+44SL3o+soumpQXrdA
1fnip+AsfKt6FmwvLg1N0z5vrvLOxRT0olgE3lAh5M8PimijOTXdB685rSJfik2xRfmyfC+GlzS9
LRlEnvHDd1qRGse8qAN3VF+22TJ+lbv93HkW4VwYUXfNcZfOVQDn1UmNsjhz4EDfqvviqfjsejBW
HH3YQ+KSEL0gV7gFidxxaAf6hRywAVkpKOyWhUCs7LO537HHueXNZzFEBylJzTBJOAxgtf+xIqAv
XxD2nFFczsO53SzSMPln0IzkIrHBUPgCnJwiGChKllpNwfXOfxvE7ov6G5l4kbhztEhWQj3I4m/D
zWjH+ZC7ITsEeWi/Ne+Z7cIVmb/iK4xlklNBvFz7ob2AoK3IEc32i1YO8gt3s/AKjW0oFZaCTWlY
pJhKhvyhI5hKNCa3w9iTa+A7t/OHoGwTZp/+GoN4EZ102s9hc7crUqe916p2I7sZn0TrSNnyAR12
FUdkXG3qkUnIw2nvvqUN5EQBLOyCs96NAfGANPVMqzqK+V2/IJ7ugB8Yz6GsSHN3blPK46NezPgm
KRfQO2rhxyQhg+uqsv88bJfkok7lXcA0E/ftDUHFTpR+mJCJyU1of+9ck8igNiV+/CHodWVZtpRW
CSZWqlqNa6BC9DJJlcR8nxc95x8WMCWUPqO/gmqR8norg6War+oB4iCXgBLF4EqT0BhKng32pEhY
B6Iyk1+wA2/fmxM8WyXtNNgzlIKkjh6IsBkL+uKqAXGRvpFE3RcFpk3zqQK35YL5kK+8FJ8q75LF
kvtZ+sNMqOErtLzpCGy6ltdh3pqm5G+KEbaiEvvQerxJt6VWXMSUuKIE1narsZ1N9/LXqBb8Vsh2
VxlQkdOdebIylqKSIu8zbIfi+vD0sIcFNTVIZ7FZSP1jgh96Aq7phywrWot4v41yF7J/V6bVE/PO
svdn43IA4RJmokry3heyQlHqR7wmd2ey0ort0PabMvCzTdIWVe3AqIYKz0BivXx4DSQWcjUo0lw0
g9T3TChiwFz5Y0CsaBpgqFHy72cNvn6CTLCDTEhtvb3nfHikofqSKeBS5DAsv2pGNjkrGiWMUmeu
UhKz3nlOJdZW+gwUR/GADpoXhcWkmOaMenkhEhGEb1ZS4ILTdL0InW50qxfVJ8/FFoNCID6KkRW9
pTekahoO8epBUy8PW5wWP70DzAer91LffzbZ8AQgQRz5AqXXCcL/2RkekiW6uEqaTvTtooZcp52v
ZYvydNlWGvMNSnRpTAEpSxHDgHJe/MWleqOsv0u8B/207ZG5VEohrROv0HSfeEfrVL0EkPG1f0ek
UfrktyxWqHUEsda68TihOYjq/aVrPFhOPgKVXAt7b6BQ5xzhqgpC31PRhfnOfWX4nt/zk/zKkAZ+
5/N7S5a35sppiKYijhgiS+foeNUOSvgWTTfpzvBvNOO85fORC7T2otmK5+52tcaQlquTguROAW2T
bYTDS20sNTg2Mmc+xeOS117yf5tWpBvzbwi0M48f3v96nGoql6x+U1NVTc4Vz660aIIY79bafx6T
FXK88zscbWq2DYcqpyfAQAS2CkB6nd0k/1fCnvI52MUmJauU9TWJMM0Gl7Mr9imzcdgPjwR/swi8
JFkriiunMNlKQeQS0d7YDcQasw5Rorytv1DJ2uFn0e1pjxmM1YTT7FBJd3yuIhxaKVeUgqKhaoxY
8LXLF0rV3AfCckT9AsWx/6e5qVFdwURe8UOSLL1LTIPgoZuBLWYl8fjciASNszvFsKUZ3Sytg1a4
Qs94nDxQOSSQ9JtNqi1/vOb52mnuin/QGe6Zs+TVFRJ78+OaSMnu0qvitL2AZoThvwogHuqhaH76
GFuGO7I4yaimITe2t3KaXor24XRWo4L+K8bBy2VkOCdmqND1Ckwibg3eNUzK/C5t60wRLT33W1ac
26imfIpWTzi+Ep4+vrLakaUMBPzf2Twx/QPy74E7c8SLgeyykdqzCTwtnyenDQ3up7jgJFM5edbS
IElKFu46h4CKhBsdIId+sKUF0UUeRo/Mr6HRiVBwqoFFZ8qyA8IoDbY43mW89fMWPCLPTWl5fB4Y
+r0IQI7ZG970CiQR/r2JTnQipBhdWSuqgkBxSynhtXoQooFgTUGk/fiimoEPRSodqIfGmfQJT+lo
gyyfahbltnybO8RT9gt5k/R05iK0FJV9B9LHwUmUYrea9sgJDFZokbGnOi4wiB8KrQ/+2ydrJX2S
piiCuDbm8682lmoi7HTpm7ddohzehwish6bswDVhAauWR39rL3lZ2QZtzDFIS9j9spvMRpE+wzgZ
DUWBNYS0kqWcfjqgPzcMhEqkapRAyhFm5cn7eM6KeRndxCZ+knSeSG8fv4DLQR9YBnYlRf9jLtpl
KlgHwduov3oG47tA2Kfk9BaMkD6IOOKedvNIigZoZTmANJe1FlQtE1NSKfkRF7P5ADuE4LbM2vjv
grhIVdRpaqIAKLL7lNwglS+f34UakHOh23JgDoYhuZCZ8O3j9GgvaNtds5X1l5DJWsjK3HzNJ/rp
bNAo/8feHvEZyhF8pi+ruKcXUhsTLM1iqKekhIvP8y5UWvLyvkw5m1bFLGHO5ZEG/Wc9tfgwIIc8
NUKj5LRk/U+lHbZ/XfOPqfC4SCZ9Liq4vegvqdW6htQRZa+fWEUjIlnEgvYJ+tTb3+5dDocqE2xq
COWX3AnNvHWbFCNxvRmF1pVR0q9ndGIQ2oYtzzvWOdy0ZItxx3PKVUBksILjB4dGYKsuajXWf5e8
oFm1W8VEmNKLzM4WL8iNza93pSHQTfgM5r6U1QVyhK0E15Xyvaosrgy88U16oxZCbjFFx4gmBRil
yv9SCZiTgzBYZNhDU9gXY5QsTQeINww+MqFFW8pWym50X9fwb87SfZdf2efswZaHloyIy+wW+sTP
YdWiVNa5sduVevHBECPKDqQXQiHs8ZTOnOK4MVPg81UEoxPDvBE5HfNto+VmQmhRyaGe4NebKeAE
BBSijnCdT5e29O+ThyW50d10s7Vk1f89xoaeu3IAz2Xwnc1KIqLTDxD4GUFQ/8dUMriVv02lCvVS
Lhdunso+6CNTOM8XYT0wQZr8E3VY2ZslN5AL5WP0FdPblrGaUivIHr+X145QNNzvJHPS+KC2lZuy
+/jlAnY1N5Y+VdUFeqys/uvLiH+vm7eug9BoN61/K8BPIUXK5Oa/HeXt8xZiRBSKQiW+1+0PAz1h
CDXPQc4XaZHU/SVNXtpsd1nrbgbHTyOyStUxionz19GlucJcAhJse6BOO7IrRFpf4sS5wit1ADIZ
cJMdwNGLvOUctDA4jYQ4gq4bkqrN8VHvggJBjze29bHFImLT1cJDro6ZwxAHud4z7mIwDBxMqd6T
97wpQSWuQVK08J74G2ss4zZXtVPN+REFuJEdVD9wkEapDegt5eNYI+/7C5fc4o48tFOXyaWOUUGE
ZFmeHT1+ifXbKc3XSUC1PIeAUnJ1GDPblfi7Tr81wVXGEKZ5LCkfn+839Sbt3lR/UakE/u1MOoYh
fraTp74bkXI4IIPKOUc2fFbl06s4GwGT2wKXVeo74dIi4637EbSWuL7G2QB0RVJWRT+BjYQbpOCJ
ZQqotilA8QanekaVT0Ju+O6cK/6ClqrPHsWerjcjTvZTWsnQYivpwOEhF/XGSPR5lToFcIlAn+nZ
mYEJFbMRlRGMmeUmYNtxDELqgwr4NY6NhzmUZllaiPh3XQYysx1nmjTzUMAPrpg8Rj9pDvrmE/xm
p3O+2Fu3qmwAoFJW97Qqp89/bwMMQHmHU3FqMrmozEBzbOTrBJoCHWUe5C7+DmXbGky93nAI5TFg
ncnQ4RapDFAqd0fv6p6rsm+sltGPs3EW2tTaqrYcLB6BJUVmWVxkdyNhjeZQNqJb3kGHv71bxB9H
FY/wtdygujMFuV91X++0hlLrYmMz7iG+65srWrU0VCZ/fF1ZLyYLTlGDaiiEHO9mbpfuNh7xf3En
at0/Ut2SK3rfSWB/DDsQolPLQaOtkqwZt8nntXrMdr7fEK0PxNpRpSkWtZJNrWAMXLPJUHYU5z3M
fBpGRtGWB/Vmdbs1AJZiSetLFsywNYMnDLn2Nqjx8NgvojD0jvSkMOM/9nuXc2oL3ZqQcOrdZ+Fh
/vGezf/NBPUmMzUJLkRKJOTJzadSFi8OzXM4LGk998IawnjWeN7CB6oVHLbOKgAWmVGHQ2GZtanC
8qnzPvz6HD5Gsb04G31iYPkL4OMgKXslrkFlwYkMYLpAw8mA5VaqjTHadbDYBJ+Uf/p8gYzbIos1
z+YZ48piWNAOgNLVpGvlFx0/8kGZHyp6DvQk3tZI6ezWI3yX1cj1rjpScz2RyvvjD7PhBNkaScmm
bRiWYnNtEjhk4NSjqR8xG9iQjxHTRqgncDB4IQEmHyF+T1kjrFh2rCnnqkt4AmOK3kLfd2DDL+sj
hT26oAD74lVdySv3FKv3k83wY7YU+EM3SB/7HCoqAgBBH04UVuPwjA/g31QK87lffhmzWHy21rmB
4qFZWbustyzbIDbyUoOOyeUELgfbl4H/UOSNOX6L7HpG/2fgfTTA8mJVrvzqpH+x3VBhYJ6EEqxD
IAz+zhEDYaT8LD7lCmVYRngyLmIthtkO6QPIq+Rri7tU1r6h1i8gyLAevDcp9/FL+Uw57BDpnYBt
jGqU3IYfM98aFMEpbO/ezfQ9N10vs/TGAQEXCdgRBl67nc7htxIni9KvRhFfLuAqJSA4B7odq35b
c5LiTWqaqwaaNhC+WeuFviQK7sv02xBy36nAcJHwAsbLoE2CcOTp+PO9/qW4DYvIZNrXA/97/+JW
z9dwdDBrYp7dX8JjTziT5ZNM4BTUK9/Hgi75hNavhFyNuyURqPxRbUVxf2eUWE2Ueujhon6Fsv7m
BuZ3avHEnpY7f1PceRa6HWs2j6rBN3vBdAEqOP2GLGQoIxWhV5u6xfGO5rzAXERpwq8T0pb6kLVd
Qe/V2A8ezKUwaBrMxNS4fVcBwaGjvEE6kMsfE64JgRjkILYK+Tkfm5Qb+VZHZrbSzx/VcEICbV/B
N5bWBz+QgR9Pn3Hzqu9TYXGxbInOJIqB+vVYmqCK1HtMMgWtK9Ip0XeLmllZ1oFwFwjdLhfJ1Lc5
4DHO5QspjJN+m9PagIp+nG0izgBZ8IaG2SpNN6P/cLV3+G29185FL0xWYL2ozZPZ+DL3sBAezgah
VxqpjyjVRmkOe/QZlJwTTc1VHwtFqSerMfL7hVgIDuFo5+2Dtn3+tUkTYT11B+CkH/ZfBERAh9d8
wKVPFnozuFPEqeLqnkIbOzgd6uo0X5+hGJCdxLr+VrmI9zvFfq7ZI9AdX3+gtipTB6PXQJpLr3ae
irsxaBCtxN3etP/81fLyvdbpmr8Q+mifsecXC5zInhZuu9DoM1tIki0DjpN/m3oR78M9hsk89QwQ
k9PSb3jv4BdufPbu9VzvhmJiFaD2YH+BAoQJfS4cD9lmFcuVDXPQ7+qPO6mSJvN5AzL3TxMzL5rQ
V9HsiXE+TUjvIIoLX3hVq3vrhh+PymgUeb9xu1gCabXojr3OFMRL8ua4umF1IRahDs62KwrZvg0X
PWUaWlrqOgqUOpVTgXbPNUjGF2d6/s05fQy8NvQ3o+Yqzu6Co2TyFgvmvvA3FxM5D/ANUGUAc8kK
9Y2i2hDZhiI6JH+abQWGIqS/LBVBxSlvJbf/+7/Jj8kZVrd7xMYUTxgVKlfa9rc/t1Qxcsat2fTZ
+K4ZYw+w6U3ALIdhoOHCsmk89Fr/IW62pabWngYgcj8vlq+FZZ1hr4x9BFUjFze6hciHemekAFcG
RLrFjSyrzaMFmCeSTFIx2wmQwD1jEuXxSdrXu3Lg8itqme9n09ILfWegKbGZo9C/HLqCamHTjWyz
K05pwu3cO0uWZG4sWQMmNYBvNJM4FfrHULz+8G9T212xJ4383rN/bqZZiEbZCR/DSHy9dnSy9Wlr
xdnyUYLkh2ul9PAw0fmqbA0KAoVEx2kvpMepKB1plzl9E1tTtaA6c3el5FgLNRWSAg+jSpmuDQD+
U9SxFnmkGwepEvyJJRLGehqA3SWMwdKsEFbRWIVVRYN+hRdySE77hMJrzAOq+kFr7cWkjRH0jpWZ
PS+RtNaCE9id5bgY6JS3AMHDo73xfmedo/qI+TCcxAwLH9S7pEn9PjR22oevQSJ6xh0rqZKrqVAi
i3F4DW8yoYD7XYywW5kpkLoaeqjRXlgqwgbTCeSaIHSOiyZ/kLXi/+6kS+lVrIOhlg/ESygBLPfJ
8GoltAvfiEAJMNmiKl03SAbkWi9ZJ6hvokihGYU+a5BizwGWZ1uoGGM7bG/1QHc27ioWEqxaFPDP
xSX68ZwcfpKaBspttE5uSYnUh1skKWp97qnGdU43Iqt67PihcbQTpOZ23MUN01ExwqeivoDW0+JN
lDUMvKrjeJPopOEdetSA48/SBq2EtHKCWVbtqTDUTEuN/Tc8/pcvawdGTQrreNZw8e2hOcmTYtqw
Lu5aReGbYXnajkOVZLqupuxBHmemxspAsfFDPfd54IlN3IK/Ooi8qTMRpa1K9s9+4iGd3r2Rh82o
vtxw6Qv0RmhiPwJ2O7e9P3PA7YToCjWikElqzVtLPJ0VvTGneT5WosqmndaS3oaGZWSU1sjACwWL
E1vriHaEKzLxF1OTLe+uDJatDAoFUwxinFjgqRMoDFePbs3sl3Uri78PBL92SF8a4qKuIF820TpO
Mkc29jpsf4+6YQl98J7K8EQgsOTdlGy261/OEBiNzaHlJmy4NLC3O7n0NGFzMZCHJB2KRDNBnCWG
S3IYJ5+QSwFz+gPedV5Gh3/+4RKJWfBOcUL+ApsDHJGuU9XXPAbm1NDdEElXp3/JxBr6N5/z27jM
rcQizspl80zc3UTi1HgwOTysfr9COjLtUcQaGET1Cf51WgfQ+/xHnL60FvG55WxgEvN7eZ1+2i6/
L0XravU6oK/hkc6gWi/StS45MGIXI5g/lozBxECcPIoDLXJKmlm2BIAfhVYl+wuQo7Jr/DyIcZDM
bKkxE3wKTbrMKKi84mJI3SgHINAmEu7SYUQjsgq2KsTrLY69PHhrMFJf0+GX+fxnIxis/bKkc6Z+
ZxjIamYLRS8Pu9oK1IJm1NyN4kZZ2GxMyfBnfNksTAIMQ4ClONToANP3PQMzQkmp2V1adHgeHNnp
D6SKRBhv1YotnYePeTto4EZoxou4xz3SbpyconOwTZ0xN6bLrgV3r72dTYZlDo77/ZM9GCx+KUr5
DRI34b64VkeNyNBjznj5N0KLuLHFz3FMOCjD15n7hOaN2Fjj8wwZtmJuNFLNaT/Zlbu0iMr7SNmb
kJ6gZbb2dtOp8uNOWs4MAQEqyRXAHQJJW9Cf0XExwG83qNa1QZhnpTfS8wyWwnb2c7ZJJ8eYwcPP
7SiZ8wYLhv4wA3EwAZ1VIWYvNxxgxvgQ2j4fRij5DAK4ck7Wtmqq19rQdtldH8NVUUoVIQX/bBh+
MD8Bz02mEGsT+SPNn2R7QkXUj/b8JfWZLKYp44U82S9vvIJtScqVq5eRyePgdi4UdONbeIr1Po8/
QuRqnRfGp33ehvV8aAO+UeIoYEC6bZphxVRSyu+3GgK6K1XouODL+/oGo021KwGqs0nfabVmrWEj
nF4pAxb8v8qGJQxuiBhiNxHhZn0GQJxjtxy/x94VXCdYVj6XJ5zheSP+DSATy5Yan+5IQIBlyH5X
cP31rgdzYO7WoEQPmEUvzSNUyrZ8Sz69n4HNtJZ1IuvQPREYFcRXIWCCQ3frN/pNUk3J5imro7xc
IqJDr9WyegNR3aCmeIJprMIfgQnzUd4d9VemyCI1xlReX4cCuOsbLcDlx8XoE67ka3BvdgvmNqRk
h75N4tsp/Zdl3qCjeTChDWMnY1iarn9QcCnlvImRkupcbLBeHRiuFsZF6gfp/yO/G0AxTWBfo3ni
U+PDh/jVr6dHwneRrJuJZ60780NZ5RH0WE1XvOdeuSbNYomFCfeEACwn8k+6t00oajjBsSqPUTv+
rQ71SeUkwWHJmMPDS17+jlF2/GY9raqBzY4gmc0b7ekk/joJmQDeTqZjIXkp9guCwhD4SjYrgUNk
srb1ElORCc/0izK7syyoY9XI+8ZEtEWxcv82aDG8wPROmgfP/pYlrJw854GTdPI/pqJwQ38Lycgw
FlthV5AqhtkszTfJ8wc2Cj26WIVeJo3GC+VSpbvkBrltZC3d4FfP8iF00zdFJAyFQ4SRZnrU3pKE
JuKudMZgJz3dw4IBL1kICRIYSSdGQH5SrmzULGxfEPID8T/6SOAkVmFIdsHTQ+FvWfISofN9Uko+
oMLgZTUOPXDPB66AfG3xKdC3YLgKR/qUobmT1WXRWo3UMQVuQYJshsYXIyAGm5UucmQOyJ1O7M3j
EZcwmwnLKlJCe6hVe2AAPfWZnF5H759CNGEVV6LPsjQGK74+s+DTyY4BkSwkLV1/5PKzQQPI75JQ
dNdtjVXS3DXQ0fsaZEI046z787eTaaznhVKUXZirPowxu8o5dj4uodpksm+AKxth6hQtefJSSjV3
4Sg8nakhjkg+79rSLFumcd1BoQeUrm4zOajZUEFrgeWWkV5BJRUpuJVC2YBsEE5vWh2OC1caBW4X
FyzA86FSkvS8NLDte5S0UiXeA96K0tdW4eosPLmL8wpTu7lREC9XEJ1Qc1HdPsC291giUXkLHmJt
JtDMneTB9Xkz1uTnyT0OZahXmtsGk8/6VN8Avk55XbzG7VVAwlhGVMuGmDwllqBcBxOpW1+Ob7iY
aGGT1wX4R2Bl78qRzjorbLnLKq3kI3+iAuTiollkU7GS63vEU7vz6behXs0hSA5sTk+fsqnql/Q/
yvFzW48s2eVq9CJJQLLgz5OYpL+NDoJl/DNTr+GJEnd1QDI1LrQase7nFkg6DZEBGwF/KIoCfNqf
7W469lwW8CbpkOjkFe7bjHBrO46oRBjOJiaGvG/ELYV05ZszS+M5/1R4/CKy9pQnQtYDMNikK5uL
w/6L241sTRqnETzbh5t2GUdkO1iECAYdBmIUcIm28j3FEe/7dkGvjc7F987txVYvDWg0zyt8yRDh
nJpZSklG/uiiV1gnvHfRrxUNgdNlJaUhsUiz5I86XYeizOBoG+zSBm3t0pbU71wlBf3aN26bC5EF
1UYNr2Iz8gid1Z+u9erteYh9qV3//tqwgKm6zfgQW0kOO4gQP1xMmdLZBZgzyVmFoAxcfraFg7kt
CBkO4CohweEkth+prlGuOaR4H+B+VhgEZSZJVweJXII8kwaNAvORFWImfNEhfK2Ymey+TLw2iKpm
7OOf7anlcpQdaXV5YIlqJSoMm1aUw384eyiRekKNu//wuK1MlvBmXviUiADpgoPyMTy2H08XzFpt
CyJblipthIQyNm0VeNbrRkQSWiIMB1dEkOcXA4Soha9GGtGxL+hZ9eEbfWZ2mWNy5rBjYndpImxI
HPdMdpnXdUk32tzRYIouZgfy+6KbkvgK/cFYVs2ykTIZf3He+a99gJyUeaRRRvVJ9ySdNvYEEttd
WKACjEU856Q7vBxWabjs76Hit72eIHSDMUFzGFCCR7IFcjWg2QNH4C7jLfA2dtgOIcrIsFKwpVtl
MPkTOhTGXVGohwPO4nf/0il6DVElmkyoW5nS+DEQBYhgpI170dCNszJJ/FqyiHsp2Nu1cvt2E83y
bfLNhcz6wytIS3Ga20i0WC2F74MvIO2DdLUM8p/Czn2t6veykZhTdApun8EklU6JxFTOi8ss+imb
kELof5XprRYMca/0RFI502CaN1VqNAnmWzXN8qUja0jERQSvJ+Zm0sXXtUrcc0pd+MKQDlr1YzEK
Xx7yY+ywAqMURDLrSiSur5m01nhBKCbMxluW/0rI7/WcWJDnNaovm//R0HjSKPXH0q6hln044Has
dTDAsZDn6tstc8R2A80ERp1oz2v0x2zErwvO0y4v8VQQO4EtV+scSAv9RvOvtcYTlCriaGcgJWPx
ZfTp7MIwPw6xD6ZW23DRrLsXttsY84AexCxJ5clNdmZB21aN6K8oOprWvropZGeMuujPohEkuF5R
UuWxs/TO9wyJT197eu21ofdRWtRJMU5mmwFDCXr4rnzCgWAbQSniMokGsgzsAoyEqZnWYp+ZLniN
74Dr7WXM5tzKgwUA9tiGD4u91QImtCenYgiqjgsR8bA2kDiUgAzDXRhDn6R+CO95W8FAaLGJQ/PY
iljDvh/CFu6jlpNNQJbfpxeY+SEzwptKBGGuLJNXzkQbUBLcPsQQhVHRfNX4kDLdagj/+0aUP152
h40UXYlY3QXMGaFmJ/BIo1fDO+oCCowpkk9D39Y1iHVIoGBlIn5mmBuf2lkgd2dc5H1kMW8Nt4+g
Ir11eIMBvb9Ik/S+cvpwCTHQ4PjbM+Tb+aqP9Nu+453UE+7yC7ffve+7tW0spGcHFdt/vJD9DzP/
ndyOHU2dYzWYufCc254Obm2H0XxaBGnK0bi54UPDovRq5RS2PaIXKz8tKrfDdmjV4sc4jYbHH7pT
nOcB+WUUuy9EDVIW6x0piXMboQRXn06LXpQ4DD0XxUxZbpBIT0r3g5AsRjj8c//bvz+E4jnrXCLb
1/ezfVEHS/P3cFOOYOPqJBEACmm/3PvKPC0U1xOdBLy5fcCENee8CSTrbP+LdspH99+XdRBovFQO
eEGudFprgq27OjFohIKlVIFT2fdt5bAo9iCT+HA0gJmVHIIoq7Yt752B7Mf5aAcrHiKuIUQrNlxD
yzFs0nciP3yKucRxECyN2ajECbzpUXwtMiYe56UUhFfQMzDwwHTz2lX9bAu4htQK1cq/ljpupkzE
8KtXxv5LuQUnqoY91+MNhFZLBGPm7on5hoyO/OwZxmAiLU/R40tfKUEmS+3WVv4dk2zDIqRqxBjE
ZPEmjP5XIUDFcjIzvNOjWZlHfYziqME5etDkpE/0BLujAo2MdGshozMWdzdG0+3Xj6R/4JPTN+8y
KUCWvP0bkdKIb52etm0AhXz+Lnq6/D4/Lc/3XX1agRVtyLAySeY7MPtGSYG57Ep77ALILdkBtC0G
p2XqoiAoeU0nY3JhtQPqcHRiZgjiMoOFnyOPf9dpSwEm+DVWEonxZx0JfBhD/UAaW87Y6s6tp9tn
8sPBwkHCVEE1mCwWCnB7veKqlTU3BkNwPamlQXoLa0zpCnpbe2s1Lxutra44oz9TweZWt+VkFApN
YPdE+ijNFc6WChJf6tvMmQWNfv/gqx+MI0ZVHYCw3ztErZ1bHhd0bjxLcXCPxzT8YICeg23Fx2ig
PrQOHnJp58IQXenkeDFrsD+vSIl8HBfHZlDV8d09jX0+i290bSWM2tOrmcPT0v2RuAJGuFagj5jd
B8jhiQ63E1019eu7Q3FXvrUyUw6cbPdNtkUaMXB6tXMc4A2B+RWfT/tG2Y6+MdvX3Yz/c5E0D7SP
tONF9Gu9qd0XjPwRJ6IdNZ4B92nrRxdnRVlyBhOJaSeWbdNN9KiS0FYwit5E+Xen2CMm+ook4IM8
YZuKf6HXVcttVDMMLvKnUMOyCk3qg4C2MVAQrevqs5wgjkEGxfAqqktgUi35PolyPppoGptKv32Z
kfaKVXRKIvzTscX7sULAfT1E6A+RTxj135tTXPRmM2RZPbIBfkHY9NM7EfapTHyArIq5DdNNF29E
1/ptBi1NFSpw6aCuEr/JkKP5hV2yzp9CPfdNL5jH6V+XxK93S0Pi8C9eUQPuuF2QjkAW6l0HOh0a
6Sfkvy1TLXaYzg0MzaXJ92BouQuUn5W1H3rpkgciP16no9kuU4q4+n3K23wggDKERyeRttX7SBop
dnZlPIkvnkZN1Ygf4u6WCGMmn4pdhgP2QEyeNCXDj1lHWjP87KNjSIsheHEtixZgramGM36u/hL+
Js18m012kmseUkk9gWPvYN1kufaVbGgUqDe4pPF7GAkrN3gykPh366WglUrlSQh8goJzh+qXQw7D
BJsI71bBGayvhM41mO+ORfAl6v6NSskkiDfU2R7OticRuRRUxDB2aixxw+gjMrw5l2HEiRrDhrO9
sr6Ru0MsXSaoixHgFY0WDqy9VSA5olCDLYWbYArHZhe1v6nTBylUZZyKMnmUnBgj1c0pdDszWTiG
W2Ah5sYphEXZWe9V4nW8oN/qKwx4qCnG6qG4jpSVEq/PKI2m6rigjLkxjR0VfjBPtmiLA+DTWPZ+
bH839xqvdQI6ohelpWDimkNrdwnKCqzm8tIirTLKirrUOdqaonb+F+5QgUS88fJVEzf2vvU2PUvR
iHKLe7tHIzP0IQUq7ZpZmRX7/YVTS2MpcslDyXmxdu9Bje4C4hWZmdhy9Ajw12v7FSdkyl9V59YI
Gh+gew0Z56WvJvLXSCo4k/lkBzKeEL/Z/aAPof8gXyeENN+M3pA7Q3kJ+jJuN1Ci1HKOYaPFexcs
2hVYTf42S/dCVz3MESP7EWq2PZ/KOwb57jJpabaAie7JGD7HFW+tsQJD/156g6MHlzt2cZA4eF/2
DgDumkwfsziCl7TrmgCSwC2Fdr2QHtbgiwkLtm40uV2cRvMwYR9/zuDISAD/nMPf5V8Toy36U5Up
RfPvwJX65hyxz0UYBHLYy7oNbMm6Tnvcc2z5+IbkqJ3XlP8Vy4ZBQgGyKyENoQAa3eu4yPEBEPou
dv2yTAtY5OUCDP5WeWohXspoa9XBgaIFeDA/OJ7AAc1whRYqlo+PhsV+79UdVbq9HYMQGIKP4WNj
BQWzb8bfHcuVfxSeEJKG0UNv/Iv6g6qtp0b3memzL7Y0vFXKDzfwAsYsuRLfl7piFFosgQuU6IJG
rgK+FpISC/f2Q2EyVq076ouGUpxGOalNNMTwhI8YnhujFjDoBNfl3wtJcGBaBG8GQnczrVH7Nsr5
PcdZ7K6SEFnwdMF9BBkBQ3+TupqzTKfTkOZePn0kSwymEeNSuBIjPXSeeCStCjtxXBSbu+sR3CeI
2m7Nah5NX9NVK1jaH/WTEQ+apPfmXQZiOfPGfsggo1+eHp/I4Li0poxCb6IvNsHnYr7UI6IWH7gi
k/mHCjYDPIJdjiJ1m4c3Eje9V/C1t8tUN8IyI3b/bixJmhMI3emsH8LbTGb515x0lNZg5Hj+9o7O
x9trV9gXLulJZ6+GuZihJKOfWTRus2sMSwWndgvzwwT9iRiSXuHFzO26Z30p/PNWHbMgnH+dihpn
ohBGgrc+NEIkmMWESQ2hm7ySlY3AKzIaoB5kI5AFsZgcQIP0j3oRc0tjVUzSrEw6lipCOpJ26gn2
WVithGMLESaRt46euCdb8DT8OVJNPoY8R03j6GBr2i7X0RXs3aDdCtrBzUyjhz6OK3VtjYNFsIHc
+YI1vxzXq2p2IEGb+crwL5wgjneee9+gOt1W1HSM3x1ZlnqFt55HlVVEkW7Hnf6G/6SlIrUyy4tP
zsZHESPdxzeMXLGsDAE75BhIc/9uM6f/Zv0A6WefePPCfMkSPBA3xpPHHFwoVtMjMWAqyxBFNOgT
NKHopyMoomrwYxvJWmwrAB3PiRz6Q8tDrTTLhp6csHqG7D4KODrJxS/IKdwj5ZOCv0w41MbJmOcm
eig6nOrgJx7KQ4Pz6XQVp+haFlP4B6lFHBUd18F9I/pDP6kPLp61Sb6rWWr02BCtoAFahX9zuQAT
ZZeKhtcGVz3018N9/a3jcJecncr1KxnTCBSlshY07lCJgzqfa5HCxCzWqha7ZjE2cCVJDv8OdrxW
PchSoUjmU4waKibxrUEfBQXow3QCkhpvvOyPPOqG+fP9AkLZgGwghzL0tPCaJPiC+icfk57Npbpm
qkQUNUAgOWpjsXNeQaAo09mGimklCwuhILTkzwoOuQrQfeJVj110z7o4Y3t89Vfh3zzSYSxyM/k6
cAUx1qeRrbF/ofaZUADUZESg9amVhxTrJRil9YMSE1tur8F03jbffFujJHbY48jTcXXetlFbEdMJ
fQEhXyhJ6BEdSmBOxocnJAet/VDBeoIApV+T0Dez6an/biQjp1wk/1EwSQ2RLWnjOkT8g/cCjpNN
Y/HZTWuZXlU7fexzt266vvN/0vYwfI4FINoxUXToJBayY+eSnJlTM2CzpNbbEzsYcP+eRsicwndZ
0u0mp5fgETUgRfpLP8Ved8Lk1V5CxYczoYzrVtptpGw9TIfYj+XbKG7lK98qdeJirizW3vrfCKC4
WOSMp1tgbNu+MO/npzHAKf+eK2P9TNzaqkXV1f3dqAS41PG6z0FJ+dVfQCXAKWI3gh99/sk/OPgl
6+AjiPD8pNcbCjJU6XF9KJUlHFYb32LBpfizLds9mTIZvRnEXLJdGYxz/LnSIn0salItHGuRyNwW
xvNWS1uM1CEoIqYWTcxyGnjCIM0sbI8MgodpVXKMJpDmAbuK6kxa7CLWk6Kw89bOO4yd75JfUKVg
Lmas0FBgCnq2MO7gWS6QqOoofhabClQyQDf5wy5APqmXxWuYLzbucKxSdGqZjIJmkjCt7lij5Y/C
X+7GueKIdXCJLTd7tSYnjJ2VWZCwUSaQvr73lIhtH8EQ0XkFUFm5hHdFDrFElGbqiGBam+SOTV69
4Htkl/HHlyKQ9yXKzrwOhuLsKSF8g7UWDZzJIpAJQZ8bLRjezoBxKK+FVmqigCt4yM8qsEbOqOnX
Fvgc7METN03IUA/l4mLclm58lg7RZHd4llt2xG9iYMkkSdbF3BhyMx3xrDCDwqXfwEoRSrXXO2KJ
sznhy+qW6ENmZO4CfE4Dfqkih1Hala+TeZM3nW/9I586MvkQ1tn5RM8Eji5ppqyvceInrdr6zsAT
ITW+6ZuZyipmjmlPzdbxOAJU+i1ITbfvizbNlK+kOdf3+OUIJ/RIUUzTJSvubrTxuPwglosu1iuU
NdxWxG8Zs/3sBSzvrOqvk6wOChZ7DGG4PVQ8M/TwvYqveeVIqjDAzML8asE8Q481R/9Ah/cDByc+
gDe23jW1l8oB/Tsnd6VS5ftUoU+rI+YHS0Uv4FSIGUrwopGqXOpv6Iqle2DlzkX/yAKIgOZ1nsh7
Sagp37EfteyFm6LoO4+EA+y63LKOli9EWauYkEfy069ZaRomLQRFwCQheJCA96c6i6SJPVnCfZnN
VgwXbi0mtUUFXp2P01LhAhW56pKm3AJ95KgSw//LYTSt/W6mr9Fh0SG5MR08HEYkDzIYboad74rv
n8FfwQrNaOZrfsZGKuXlHEbKrgpb0wbnbmynCa6lhJCODMqFMGnlMUW3uA3ItZfymFwy+F4YEfHD
KniHY7ypSNr0IbFK/00GYL8VVAcPzxZr3IIDBW3mIsIbMKxXp4yQyRYsG7AJmdyvqnSbzPJYcktk
n+YuLHC6/tOx1O2HSlAYaXtamH6mNxtY/uO4fAwwyf6/f7kIib2uhcViVyVqEUiihrXaey9orWgf
xVryoFOY2XsPHKHBbZzUr41apYA56AZMXQtDouk08V0NM/mvHIUN9wmBYAfbLX8ltLrk33bS6MIM
t4iPnDYgCVu9800G9Qx92eqiNT4VCwaVHbcTHdyn0gAnTcHK2lCTHcpZPwWs1xzEhuMpPBbq5eYv
uXR0zFK56dRWAfjMQ1+S+L9Ow9GsFNyhUsTkc1Q8lN2p4tlPjhTaI8vUg9adb8oItlYs3jDsHKCk
8yWeaKhvnBz1njcygO7CR4SLJtWC8q+765glqGBKd04m2csFRtuDDKXEZxp1xhyhkXXt9Q1z9lV+
DFW2UVDOc5Vk6ldECETtqL5yyJxSUCtLYqvbUE+B3DhRt6LVC7vHTYNTkuLwCx5yYjVeuhFN2UH3
zWcmLs0er54V7Yk8Biqf4JodQPsxRZyFOVNAYaIr8QFQ4n0wrtXW0/4dJpIX9OqlKNtaaqm1ZHZs
lwa1bh46/dibx8Q/W2RQrAmCCD6fl5APs38XeODE6NeiGwk0fUM1x6UAJi0kh94QbNwANIWAMT+n
V8aMOzsySl/WKLUPge5r8l+KDpgPGhL7+OkT8Y7yEl0ccD2/L5ogytRsESgI6vEeIZRY3ZMVEiMg
t6e3SlCbewNccssWHWmwUjWzc8l4IqdxTqmfvJLElOnIr4MValp7Ebf6W0dhxjW4goN1PpAi89Cp
6s/yMVzVrApgq0D0ulL1UBxXVZ+BNTGW4TW42ZwMbgbagtphTks+PsjhdgRvJGdMMdXhnWnhFeVL
b0MhL8y4PFmy04uxDwoN8DJ9ha0h5IWNOWjavB4mBRBGbE+o0SYRgJl5MqHEMIKsCx7cIjMJUZJY
EuUpXcFLP05aSOMZBsv3Mc/ITuOQwQPJv7WgYVSGBWBvX9+/3T1/eznJTbBW3Ro6If47kaHGIafi
rvpFKdJSqOeKytppGXqUCE3OohIYs1gVI5J3yT+EU0m49LB44+HpmK2iMGuz+9+KzaK23iw07wfl
hRH1UGRUUr0vWK1nkWyvJIavWScvlEjWFLGE5pc3kCJJMIaHwPrmGX/YyncbPQH48w2Xtvt0IYgB
1AS5Ji2SWhBJ5PciJKvpoqLNP4gsjZHWE4QMrAE1X9Wxnmg1W2K4SBekg4FVvhpm8f5ar0ydYSNJ
ExHF/C5KHzoG7xtlbJs1Y6dwnsoZ91ho9IVVOwmwNoyi7YBtSDXT+X6q7yA6j7+BtaOnHn2zgrNw
rRvVhWvBn1jQG62F8hMsdnXQg4ckG07i0aX0ze/5EeDj+xJgu4Kf4USJBn1ic1K+ZL80p+Dl6egy
7pqIlK3xOzHaP0EZeef1B2Z2Gy4hJM7+ejbL9/XQBypQCMWW1HL+hGkdaWc767a45FxaUS7RIgi6
+3yFNU91KsNonL3t2uvmsJnLYI37doAvRBj1CVXhieYezWAoPDEDpotIUULNPnOZKBr+2exIPd+p
Wv8HA8KeaBpP2bu2wX/5EXhuhLW4STBOwlpTkG6t03QHgCAdLAKCTctcSrWKLoZvG7RNTklvEAPl
XYMNTR4ZVx7f6oDgsQ6Npu+lh8uYb10dvZd6krJpI4nB3rFfnljfxmM6KT49Qaofq32K5GoR09/u
ayMQ1uhS/vWJG/j4qeo+vAzrtSC51YnuC/wY8PoSC92MtIql2AK3i5jt9j4y7gRJf34Foq7fUDoU
yuy3x9zsEi1g3au3x/y6Ed/BPlfTz8uLNVUMZSf/I1nbsTJUjZdUx7ZqPqCOat/kq8H9Wq6AB/0w
PpxjQM/rFCv5Yt6aIUT43naREMfzgCu0SgmNtdRfcx+Rwip+YhmK76JA29P1nj02xlUtTUJPIRBA
JkQn8oTgvV0enp5GNRhU6Wdi4Lnx0uLTeciMH3EqOsUkYm9I+5B94Af6arwRcSJfrEc+QgbBX6qm
UFsJ3Upo6Ncc4Coy8/k+eV/OnJgAyefe8aN5ByDoagX0BqmNtwu/fVIDUTNqEUF6O2BSA4UA8nVF
31IbjDoF8b63UQO756wjBFRb/56832P4iu2aWrxGddTUM+B9qPvzT1mwZiHwl2LlK85C7ti6dw7f
eYFHpotr/3YdAdPD60bGzMfHHAzq4arVGl4nW4fS+0OONwfQS2Xrou+4DtTPFJZmrB/Z26OIhkHn
VSueThGyVgryCV4YRIo87yaLTqKcReMaAmo9IK3kzaeUOPi88rKEdtRCrc42eKIw/m5Io4XwsYE/
GdogaMc4Hm6+swksscbqDcozV8uuaYYXuHQH+8yZXnRXY6WWpRQ=
`pragma protect end_protected
