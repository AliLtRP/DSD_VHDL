// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
W2WfZtgWAcFsoe9+d2foA0t/XHUH/m5G4m/9jkV3CoG0IM9/pb+UymOYTCZfHVv8
/4NDSnOuPQw2gIigB6JRKKEnb6eQx97nI7tpQ2mSPi5qME7+LgRLtwz7a5J23DNj
tJ0iGzTAIZU5AVkic8y3KwnRYGubYepEZe0TFXJmbJg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1920)
kIT4FEKtdSX9J7Lw2Krqbk7zBf32hNdx+LE8alY7GnU0H8GuGUm8Qg+3AEwH5Gjf
IBhMFuhu75npHz1tRFyXVYi4takjBhp8ar4QE0eMJ/slCuzoov6b76m9zzPprIf5
lhkqg86+kz9u3DOB2EPMuhs8VVHTeGpgQlnGsYbsPihIs5oNViTqPwp4dL4MMFjq
KZgWIYS8nzPiO1lTw0Zw3JmLYk139SCH6ELgfyv5brZuxQxeS/WV4F2nXj2OugBR
soyUIhIx6iCwh6o5gIkiWXnk9IGM/aLLDhiq9YSSTVUsT8zHKeVwefARJBVqgBVF
JfKNGAravymITOxX/nT365yDphZggB6whumEt5Od9mewJcyF5anhc0EDVJw7nqPj
qRh2lbzAgEKYgdRucYgVcnYRqCRAxPOBWH7rJNNHnT5oLz3zWI0BNXIAZRBRjmfx
+szZMhgGuq8jUCIOpJ7Dm4oKqHC8R2cX4PAdTM967P/+hEGmsTKRjiEfYkiCoign
yNhsxRil+i0N8wHMfdPtf6xG5L3pesmnJ6mzm/gfb4X0WBEAUz5KkP6WLGK+eHka
I4i96R0goC+EL1tZVEMfOPgDpSRdWPAyVJeM/10pJRZ0j5sAnQVfntByOW3pCPwC
HOXkjq3WBYevA3iqjT3W458m/Kf+H2ZxM36KoEFwNQS0k9TGnDAC2OirgJfuhSIz
542wC1pcsv/Jlk0EvXeZRvNoQefZu1psry5TYkEc7v73fgNMxLYRc51G8e5NLgoR
iR1cpiEavl5ggk4T/927+cWdhP2MfPjhMgw3wumrDXKaeUjx9rvcKgeYhlT0LE+R
ofjJLDpR+jbj5QDMoK1O03xy6nA09cJ64EFfAvfFf39zr9gzRCR0bYCCGlDRyOPR
rqb+ne1LLLJZLx929y4yt5yxCsm7edRF2JdEP3caRTb8OwO3TlLMAauPdSSu3IEv
nssRbHcf3JDosrMsCFj8OATgpRmO47rRQKNJx1So+vDIWvu050JRIAZ555lv5c/k
1AXyjWjuknXfy4KlGbX3Ob4NiA2raVBwVFBJzcCTZbqdO2pHWaFqtc/E9D7L4WVl
0X95NBxXHKIgR15csCvYdbVtJn7nwa1+1NhCxry7vvniJ2QYcioIL54v5zo8KshA
O1/XsKJeV4TXLGyStZGslslX+e7AawgmCZn3RWooBVm32rsB7z9s5c6aZg7ADb9A
5MqnxjbmgQNPJpLprYB1ws9fHsmWVjna3UjmaW3su3STAsue1fzZpLzwMcIBjaa0
8XJecFXJg9rhTDYTz8vTN938JXY1zo/84CqvfW4IHKpC/BJZxR7pvLUsxX5ajT+r
hjHV+On3myRbLg7CkVY+GFKDHQ5VETwf+lMz7f+SHxIbrtv4GVmIe0ZUL85pCqBP
t9/9kL/R3MvfEjSMhz2JYlufiweReJ3hcEwF2RvkBvU8hl2KUNPjAZpJ0bm+SrOY
0w3ciVNgSg4ulBsK4jw2JPw4Y2yGoOzWBLEtoudhulOUh+nDNTomsBEvQaNpF7Dg
G5L/6uH6azjlOHwzvKGvzVGzBIwMf4/QQBZuTnDdFkB/cjd6VBuPOD4hsxxjKdBt
4pwwfpDyqnkPipFV0917lOP5UfFMruDfh2FlWzQVboF9LKaHw2xLZxcmOUf69l05
Qn2+iJ8I7zBiB9jr8iEieKlkgZVT845aEe8daj1IWUV1mQBjdo4mKgxyWINncHqL
lhGPfDixB8TIpoEWQPI2+NWpgTTHylRnH2A43tq4P6BagWovSlgJY6wNhHso5CNc
aiGFc6BX5smvdcpTR3v6rbd8IQh0U9EGdH7DPIFl5yARrYFOZi0WUczTVvMm8SOk
eTQev4kkeSlVvUe59xOt3DBrSm61HbgcZfXhc6x0cW1NuTpluOQPZhPs77Cxh1L9
nsVnJFnSQAZOC0hZt3DXitpwYZg4OFbrdDZf54on0FT87AjnPF8CLDU/FLTbmApc
ZGwho6Y/9f4ApWJHuikWUivJnnOzwXbStjtt+vHVu12Svrea0kzcpuwqTGHdPgCb
QYO+Bnpi/rdKHVqI9Mf5vBV4+kMcc27MRrft7D6xx+ajULm+UPjJh7J3CKwgX4gC
zjndS6qz1eXmqz1bIeYp097QpmROdcnj+BXzuNlscPMNvEeRYTRi7Thc1GsQo+fN
jslWTRNV1BBjGZS1PR05+p+NMgAoqNqnApVQKRcFv/1UZ7zQEH1fAFzyf0oNJuVd
xx82w+g1barA958+3+B4PHOaAg6ttkQDdy+w8CE+e5e8pAFb5P0Q0p8rGxljMAf6
zSeeWkD4kdhVmhbVXmNIb237cP5IZ00NBX7oHiQZwvoEY6MzyKIKPUoNncF65R7U
Fuj0ru+miZ0xFUvZkpiRvOQstNq/3tJ7fLKxbxNCgoKsBH90kS6oZs2QXAsE+26A
HpCzK73GWjFJv0RMbZZl9RMdAYGJwad5AD2/asYNN+xcW+Sovb9dc5wLcoPUdHXT
Pysewi3tAJru4BLv1AhayNLBFUdK8tuKVHMsyoQAt4iQBqlwAtK5+IVsOvg8lPkY
`pragma protect end_protected
