// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:44 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VJF3FZ35AyQwiGsggM7pghYvJhJBJ/VVbU+4JZ05msQUiIh04ht/LlMtTCdqKzCQ
S+UPf6Fct4arVY7+BD3JcJSlBs40A192OrZeDYgtqisisy0nCSB3MEhvivz5T0Q9
TXD+iPN/5muoUzHrWiXOASbh6PhvlAPksUmAg898o2Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17328)
IshbMcZB+DPUDjP0y3W25YESmds3eHOIyUp/rmRd+vjUsxPDaiR8qWK+MT3DAPcj
DOfP2DwKASdZNpKamYyzbXgGZm2u/f+QCfPIg3kFPNAZgbYJ59Ep3luZp/08M5/J
/zEQr38DGESaUbZgcop3xMtgPkvN/hpe4S8d5spFZ2VV3SeDSC/xHgTGt9xKj1CN
IHdlRIEc5UkyNQRR4f7li+1u3c0VGwjSlfPVfT1JAWYp3R7LD7ly/wcCa3u5C0L+
4WzoUY1jtaMnaGKb0gGAGJ4ZvnimJItvb9X/eba+hfifzCwXUDfTt9xaYcrEkFWh
U2GQkIdIub2ijg+gNd5iHePGpEYolFaRXnelbRcek5Q+skb1GMK/8p89JOe5LFfS
dQbiYsXvHj7Bl9lp3lf8bm7h+lIRwVZCCgVH+YV0RcpIVkj8DGZyPNumspa2HbNU
vSZ9gFLTFAxoDrXWZPO7Quaey7A0uYqNv/MlNQPCBOKNu3FFhNkTFmqW/r2r8+Ub
Qe9+puqg5xfNz83Qn6+kCXdBRLJjTO0YfZNFW2RmXBTxNTGd+Ox8R/+m7h2HSzGA
fK5TyrJRxPXH4OaFRc3wvbfLIa9/eXaLT+KSYtgfK/yh8kotjBmIRuRE131VX8fr
qjyxcBEi4xWiRTEUznzj1sznzjDPWT6IbGV0XKTo8Yx+6Wfvl5JMaitIB9JIrgq8
TrBRNuSEPZr4aQYKczqqpiFf0jMxfT0GxEpzLM+aZkApgj9MUKwYui+w02OwQ6jc
uS+zWSXGnd5H5f38WEmyTgoFfUK/XrsSJBfDhMm5wJPoyFWjJj+sYvcDjHKSYreI
yNJ5IkWoXiYpnu/2V/n+C7kBzaI7iDT+bfutIuKliS6efjY8haDJ2diKgU5jcd+h
2/e9a6QojtdgaD59vkxyom7jkAlq+ITFd4KFvl+GY5mnJRe8S4cm6QLJUZFQ3AeW
tCdLiiv1Xzxi4ruveWCKwnRncBdt8xJmm/qVJ5SSi7KTFPsyP5aPRscrTxQ/0PMR
0Nok+AehRopqCLZfle1Ynw2oPiMsov2HpztXGEOu+Ar2zkIhAq9exJ+1xJqn2Yd2
zXLWdc4oYO/gCYsYWi88mK3TJGCXFcvMGHBENPAyAEclXqYMBeMZnhSyRHNKsFxh
F5n8ob4T0XDrp/rlGznE8ip5zJ+ciX2u4QyHNtWJQX4reQFIlYa8Bnm/1f0hr9fH
h0So5Vfn36fOn4XCRTwlrdBygUHcrHiUPToUkUs8TPy6tW7CwZvTRRh8mUwCEgie
M9Jy7Dd+0ctOV92rlTSdqKVtimcJz5vRxe/BEL9IqRgpaKWhB7WDchMnzRaoqX1U
EKYnfDqpqmbUzRU4nf91i/cihNz8GHKDzCNCIt0Ud4duRe7XYhJvrIeRc6rzqOai
BA71Qm5ByjJ64mYiIxC9DiyiilpmyDv7gTcQeUcJt8YLO2jQ1Cngcw642PNV4njk
+XKmxI1Mq9kDO3EiHtqK0Qi39SrwhdN3QyMuNlnLZBE7vzkzJv3SIySWNXzIU7cD
gE2xGF7TIUoGfky5cb5A9jciqP1QqO/YKLNRKKSfLba+fKBhfD3vGV2NcBOk09ns
QWUHzP+qge8XLzmNYs+GTf+bXAY4QEJlray6haCGHnJgDIifWyFaDceX5L2K/VoM
RaFmo1pxzYGNbB2OCzfP0W6lbcIzlr7wsP/HMA7W9qG4kFzI4JJt5kRYZDiNzRny
be9ZPKwsZ3pEPnnpFTtiuXFM5UXLxgx2qOJmYQdYVuztjYj6Jyvv1UYmPxaqkqTb
ogIv57bakiV/U8Tzd6Nie9oZClcf4zUacwzLEk1H/Mc1a/WLZeVAPhcYIrN7WOpn
l6fJTpUgGDs7nRgls9pIREBUiYjXaQffdAT+SN/I/YvLT841Tlj8bSYRjbQzt5YS
mTejHzMl9JclFN2jS/+NVi3C4g+h7Q9lqA2l4wIsVV/JF6q0mfcx21oGoSkLLG5T
8lvS2sJKzwc9Si7+8Sd0d6ryv7Q2u1baURpbG2GJ+g57qOfnBviysqD2kDbzZ3an
gc3fBV1jEYLNx0z/Oo0Tg0T2Dd41s2ewF0cCRDrJDZX+XUbHOXYY3reV+zDKUi8r
B66NGe1H3QIkvMNvzZqBq3W4ZFcfh2OIsbi+0Pfz8OGHC80pOZ3a+Yj5gaoizpVo
dKuaKo+rXZ9DZV1h3m2pyDVspDX5xapno1PKdAUl2G+qiPwS/QzVyjgChhaeIevg
DqI3mdV1SUuu/OXLq7XG0Ch5CLBSVBwGuN1CZGVXxub2USZmNAR/mcFU14iD7i7W
Gsx3rjvt4fJUA4clDTq3UD3lzH+veqX3O8z0tvZUm74gmnDm/D6GJ9Oc40+ml8AP
gGksbBU3rV540T4BKyLaQhIZdMKe4aIt3G7BFvCV2izXkbs8+eq9JQLW3R/thexO
T2GyivVR8tSW6PF512E2jw/TZBIgpEItBToucsiy7fBOJcF1t596XS1D5DXbqFAk
uU/rtwz8lGwtJwK8469DAERfy+umfOhJJ54WZYPwqrFo84dzcD0Y26d7wyho8qP2
9WrY6WH0fYjqWw4juPpXfHbVPzmVuBF6yNRUmY2bW2AkM2HSEKjvnDfhMfV/dfJg
y7p39oepubZuE2vs/Bs7jchaiLllEZZmTUk1WryNY9dTi7FsjQSkAkoIx/9tw+IY
RW/SKRZkNhbrtbtm14IZYwUfc6anvbAc7Nz77yWAlPHhtdqv5rliLNygMOgaHTQz
xdljmmxo2N6+/QkP9ByiSNk1WymUdZQplc46v1gQmIk3yZhYB5M52jWZru+6RtJa
0nEZxFbwU/n6oJJ5MWrCWWyRsnbykt3RZFeatIykbFH6Yb1brXS49JbW+5+GCOog
cSafXGD0ugnTN6IYpUsaFVWVKh42s7cGBZR6W1YSTkaV6fLLEQ3LlVYj53FXUIY5
RSTAlLmTgPO8xTsBSpE6BY+pjgs4c8fl/UkLBsAhGJ69fyEyjZb/HPWOxIo7Y2Sv
et8KGmsknJ0nCR6m0g0n110c45NUwNcq0cIyj4d3pQatg8mk6kTuFWdzmyntcGRh
VguRV++tGFEZ+VhJaVbL1SaSNnklNW2sEjv/RTEwqJrNWQTlCJCz1OY5mcwMHbDa
o5x0F2qlOi9Nlkb2WIGPv0QizHUz00ZPHVm24GnRinxWBX51k/xuf8m46IlEYiIK
2bDe8Xr8zbIWQAyBlS9cqNKoRMFlYsThyFlm0Gt9R2AxMB2If/6XAcbH0DIt1cZO
XL/GZuqNIdXaY0z97yLLxUDBFUAibQRonuM3h33haXJsR6KzEQR/lPgMhSIFigfM
snpLRJDYq3x8mxMAHW/fCg0lsjYUcfqIN6F6Pglixvjw3CBQ/+cw10keLqigzXif
nGoMr5v1Hq++91XFKZny8Bpiw5qD3mVLi8NwABJAOu3C6Wrbg6CrJv5OYKVFq8os
jephZBTD6y4sT1KfUbslBLp800z6mKokyLYDd2SUrQXW0GdtmzZZ+AlJlaUZat7i
pd4hqi46mf0ZiKJEbRGbRgbEwrgzJn5fKAYRfOAS+XaKt7lESnzOJh0MA4wxmwD2
3afkCWYIeXpBApNjaUqABZVnmpNSIQiYBXr6+yRiSulqbg8bPrPA6JESPzoLtAsc
TrouTKA3FQTBAhFjUNHM0kmCFfr+5QJUVJHVDP0/KQvUVxJM0uGRCiZmL7Ft1qQu
J2AkKTenm2QVu3v7ooZtD7O8Xmhgp70Kvc/h2nFHmsd4Ql3zZYPGuA+Da86aGOjj
VVohZXUrBYPgJDZvnIFJSPI9+H0gmU12Ih+l8t+QZIqUU/XXmLNToZfQO6Vwn9B2
pBANVxqgB6X10UDC5W88R0ij0jhWUzHD1K1FMvCjRixvTGwcuoLTp7G8FRerx0La
NBleGMKIZOxZxSWz0e3nZTACm/q3tpTzmZ66WbdaIg1niYnK+NthD65k9DKLS8D5
bPPt7bKyc2CHFIB3eJ17b90ao096L7wXJgZ1E0x65bVQTADdXzGfhrXrJGJEz5vk
7/gbVwao1xV8r68LJgZEyIq6lVI5rndHdyLrXAMSmjOFaFdmtd6um5m2U101e8e8
0ZOfaULIrryLWFq+hTXnlqIc2h3UjpqsxZqfCwypFaE+YXdgfvlL8KfbiLWFvIud
e66wkLAlvFhH3oq9FyEScc5V83ss2kSlfgJBDv3XAD/q1lqxZL0dvpQHrpBnuyf2
Ai4T4spAMSXtdyppkwg7esVTEAbaf0skgVdCdEEX7aEVZy2lzBO3GQuogCSA93rs
4foiNFINWG07WLyaj3/WwRUOpqSJjuAbYfogfz7MffvkVdvTJoiQ71mFNS2Qw0cV
Ch+xpucbagjwaN9z7bY025bEpLGRq8xOEUUl1ESc3EijVaIu+D5Q6UGS602E/gju
JubGUX6574D4J4GS5hBzbgAsvwY7T0SBiZfXrJ69vwOwGsR8ZOtPTmFqlGblRddT
XHITt+SAUSiJGpgxVW5L7GN9YMxe2ep587r5c/A5Lf7S6+88sv4Nevg7j0Qf740p
eQ4jsGuHx1rMPm/MVfPXNpFpxhUNmYvD4L32stOXthrdxVjPygjHQM8kFSTI12IG
5cgktyK88+xSNuoJ8XF/yqfYo23UwrBZfP9MMxlUFw0N9AV+pp5KG+t+9fQsv87+
XPYmdW/ZO6cVNGqMEKTVKsb9YzpG01vjExDniGxAusJqjSzSGFkc8rXS+hGkbqVy
6BrK6apG31srz5Iqktxwic6zitq7M5OgXqtwEXmR2ydZjK/ySmxh9VShgUyrVzqP
HImH8/0q7E80WF0ZtZN+dalL/Mzw32G9mOgNtkO3Jg4sy48re7TkIYqENwntsoEL
bCIopkrllVLOwiaVLWRH0rbFvdKiXa+HeBvlKpM7EBlXZdnvw12psFnl0MVhbLWQ
5GaP+Yhkz9OFVXHloW2/fAgUlMrJXPy1tx/rW/3jAWYnUXbUuiE4stO3himbiCtx
JrRjGHdPE6XlPFZ9JfYMyu/S9vWgSS5E52y5tcGwcAXnhVfw6ueyCc+cvM2lyksq
cGTCuHFJILcAQNxSX7hmHeT39LDbPy3WfgPqrIJT1mqNnmWKGZx0pc9/cZcMqVd3
vObOfnCEl5T2Poq2oiYn/CdVdNn3Jbj8ju0gQlV6jUDzFpH93q2jSoMkEYQmv7H2
8OJ5a9kskaZBcj0axu7v38ZeMbzKZ+0LQyab+ryPT6NjpAzorKTN6Um+MVMcKYgb
SLQNiIa6bxhjy1QK4E7b/N31VdUmT4UAoo+Cus962s0Q69pzP4pNLNQQ2T7ftqJV
1w0ldwgThgtsHf47tZbLIj76EZcXTvDfGrE76sLUebwMZFEj+LuoLgkAR+xtw3a4
sVqVxoeDl0MuNOmfnMA/+q0R12+HP4GDTH5Wm7Oi0TgS02jurctKpa941rNITd+U
5vZvfeJVQbKMb0bybADLh9mtZZwyrnhztTW/BHJK9r7JhYLzcM53nZCKcc+wIn1z
dkVWUqNGci6jMWcp86ecPv8B3ocjsajCSconcgujd0AufZVHj55LUZJ/yOhN2Ivk
LlXSEB+euJcwv8zUq8ehNmUdU63mPcjUtNmUdywT/qeQU0JoKoVCyxESZSwVI1N8
bwAyln2oJUcs1D6z/uxKiNyYHtVkAEO9PoPbuNrJUW+1OVUcR5q8CRku4LOTdyS2
J4294Z8nc49bCxFfMNdS0Mev1/7dVhNwN9/6xWTJwEk/AVrx6EKCpF0rTuMOO7zp
GWV1IeVRb49O/oU+KtxfsJRQ5CQW7l+OcdcQb0kfcTkVdymayb5lal3nLxFb35Xj
JnW29T8ILff4uadpWs0/So0kK6NCZ7nceUwY15g9u7eCxOfCCvI4hYZ8PwFDw/MO
0a1ShRuNfCPR0gqBY6T5f7BXtfDVVfMqgvadJ5UGsX9EokiZPvGQREASFwmqemJf
gtMdElXW/wc22zsLZfYV1vt4D5i0ifXYUYo1BSR/AUrHtoVqKUELqthyVy9U22GE
rDlDTiiaiOtR4XyGZM14pOlCim9FJb01QpwVInAXDFKzsVZy7Q7ba4E9HNWCHXTH
Tr3VfzovajBi6/m13lRZuMSwZkRSIuf86BBQyAkhUTDPc8KBgQdXoX3vMJkTZoLS
t4vfsqnBAU7Z8/7gfE+XkmjwFr07nM1hPiBq3mFQp10+Ct86QEQGXnp+jFoYyGRz
rBJjKfygC8Yod162iZLY4FXHx2WtBDdsJa57W2ivAVDiPUT86S7qG/pH7q/2SS3m
X/xcvmvxoO7AKtWAAIkaxRypw/rzHYftqbyQAPqyt2fPWDzyKj+Nlgh4PcVTUSC/
t6KgnDeMFgkap8ATJSxLMhP5KoYjTh7v2JKmWSy+YTbS4bNO9ZZyOPw43lhQmdGQ
jyU8SPbMs7KOZIiNQu5uRJy3ccgGqgQaXTXU1lnMcHyA+1pbnm/yzwfPMiIcBoE2
/dLdkU2lJkbI3kPICDJgGkHFBGTdX9QEkV/zBcTEXwjEp+7VL4I4MDwmdyenp1Es
jD7aQrsdvPptsqarvIhii82IvtBC3KBiTVMBnYp5ZL489h4bliese86gh1PwAEoT
CTGTPV22fyhuAcomFi1L8VNM5iQyCZVAWiboaV2xIpf1H8GnbcJDSIeOAgetDYar
HeqIg+0zGEd7VDbOf/52bRETkdqtz8/X12uXrxxzJCeamlycej72lPyWB4rsRfWr
+F71SwH+zDyKaDNtIrVluhxK8SIW+JCgAk7GnbK6Hemswk40Q0FaUvV0Xyakqi9F
HDUjG8gUTIeIRf/jkZfLuMfrWz8QJDmc0PT9q8qOJR5DjBohQ3iiYB8elM+U65jB
wg57mKLidBdWKVkRRphopSsxDO6IahUkx7RYuPHHyeW+FgKGAuwCHy1zUTAjy8DR
Cqk1/RpPUrLgbEBnNtlelCFmbUR/vJ5NODK5QgZ48JETCoWPQ6G4CUxvr9oMKP/Z
FqHW60BUza+IVAm5hd6HtVZHTaHrpKYdce7D4M6niGwq0nJJfRy7fxzDDR/HtqfR
pgyYUOhEeQ/twa7QsxR7H2SoggTkq76fyhgDI5GgPCqiTed/A/lNmhXvCJCy1HTr
dk/p82msckgQ/o+0O+rZHOkFujcxXY5R7yngCqvrvqdKzM17FTr+4AjFcMgghZt1
NfirmEl/lOcvZkpD6ZqMIqoaSzfDxMDUY7/bs7yhFWMqpRgpoSjHdyLPtnvTKLkK
OlKaeT44gUb92dRFQ9V0kUaDuDTqh9wZHDkmryr4kuheeWHBWO6Nw7e2LBcFEgqF
F9JeKxP+52dSwW78AzKYnxC7UkSWVNcfelxqX+HYKQ9dLqCruWpBIq8k+hk/qudV
EdO1WKeQiCbupLwqaPwBiM0cVmF9bw/P6WHToCzi4QQ6KjWkzdEg52RTi8VIm8kY
GGXGyQoDeJZeWxFRKziy0XvwKPUOmVsCkUdvdqzxcOqMbzZZVKMBIEAiAkc2VQo8
F8cmfziAiymT+C5bkIoiVI4ckpPUJxe+he2Y1fox3jjicUaNEvR5p39vmEcwouX5
EgetLPhtKxuVyZB7rLQf4GIBuFu0cn39iMIhAiUQv+ekaJJdSmvaan9ODhW3IXTK
GxvoJ5y/x2sJTwfMvSUdUIgrJRFTSWD0y6QugIrWT2NFqUwbPjAuB78/Rp7IAuab
G5cCZaehXEzVxa4LoN67vaRLG9UPXXQ7bGIMM9PAaQjjEexHoIz0Y0cg1MjTXcrm
SvS9HjkKGNOqYJtI2Oz+fGhQTTiyx2EAJ04gMfIVPwTsxMFyiEWeZ2o0pJ8dxu6k
LJOkcV5ecpvvUozLaUmIXPsZ/A6vI+d+e50nRIHVZEkgdN1c7DcCRQI96eaXBWMJ
R4VLuF0CGJEfbf1wZStBiD+cPuCpk0lA2qGmRj0iB4PdndAaf2diVLro4DRMOgZS
0YBugmnaM02mrkLLcFv2Y4VOqvf5ZwdBUc6gRS0bXD8VAxgHTjF7RcPek+no9Gi/
Ylz+44QY31SoNxt42xcB3/KYa/+jboWN3X0YTwqw5vGvclr0Tn94/DYcQk2aYF99
biPKbYZnR4lNzSflORCmpv1F1TL0F0qYWRT99s3HmHo/2x82B0JdgYFa1fc1ISvW
SofYU0o0oqMF+BOMS6I3AMnVasUOl0ISaomrd/nE5LpdQ5a9bD5yrRfKEaZrF6U7
0+FREo++BWbkrb70BeBq6QyZdYgeep8yzGUPbDiXeXtCdAKMK1MKXurk+dOOozRG
6B6vO1YKQEsL2gzyGYpYJy1sOhinpCQJC8fJl7MKOSvdaM12ujA8g7K/qfQjoW9o
4xuUH6qQZn/URtKTg+bbrvZsi4pEjpLf2U5zsmCzFP3OFFHNFTFb1kbkwexXL9TQ
m6VLvTrGKHVbx+mfhIjkVfa9BxCkc+7/JkpcnHDNjXuTnvVoEgTAijy5zEPRRJNv
4eU8JZLTK37FF86QfGcQn6o441k0+vJxnENaUknvWfcQo4zLMpZUjGvS5hXIIFcW
KnpXvao2qovXfTj1UWAwADoCp63ZLDZnnaryYvicUBU19H788/eUd/rDeO06keqp
CUGksztIYlzjuaNjf8DxlDMccQoPOoRpDUsFDMoRgXs/5ERJ2n4sF+ZL5kY+Eust
K44qbrXMiIC+gx5xCXqOpxKFaE0wf6dsACRrYxPKxiKgCncdKNa16i/HxF0tPmvU
Yfw6pTMljlCd60fqPwb5gMaxvd6SjqTt/ULBuWI8+ldCcp/8S4p/Mf0QPtdn+Swz
YVZKxiwpILETUToE91wHAteJWxFYy/fWtvzYQ+9F7MHnz9QLf36ATMWmjlbf9HDa
8/rS1N6Kpgu1jSTjzrFjNYpY+W8R1nxdoMVxxrXiIMyQo4lnYNocNS+2HF2AW1yZ
8yHoKQdxiojeEvg2Z6sqiF1Gb0eHqF1epGXubQLAVGtEJjkLzcJi3j8YftW6Rv+P
oyjLuhSPSYfa/9+ij9RAdZpgr08uWvcDakBcRg6YQy+bXFKlX98MZsYFAm3G4zvZ
h72uBN1ThmWiJ2dw7N06Nai0KF6oRfdGG7Paev6I9P9SdmIQCzP//jm5jbjX2gzA
OOsvLQ1rEygRdQJ86TwsSuhuB/wcXZ0XRuEptPGmFk73vEoP7i76rED590LrOKnK
47AZxtRC+CB7xdQhMr+LyK4cDMeaLB9dktpjS9gaA+SVhEd2zml6z3J1TQVBnPj/
bGH9cgZkEpisfluTsPF8xQmJP+uPG2muBnV2CqE3KgETTTF+5SK26YKth3z11jlp
FCoDHu3flxKUGTtKp2q+Zxa4h366oUpI4zjZEVJEzwnZ6aH11BvbArVv7eBt5vlG
3ApftneGjSHXTx8Urxp5xOUV0h4WcqtldCHO3cG66cbJp4Ezw0QwZXNlKeUj7Hcp
7doSdSKImx43Qd4lxA3y3oMd+DiRBW0JF6GSIgU4mEWRJIZldj/TC2kELU3yJviN
hgBrQD+yGb1Zyyv0i1258lwWegHoHfyR3m1sRVW64DiOAL/DVbx2IWV/zwo2Gq9X
qoAI9e8vvCsS7jPdVD66aLjxRDtjXCzbfSZf2/VMPPoGzSZnboiAsrFSJNMXk0T6
OX9m5nQPBvBctyAM2Wgaaon9uUObjFdGerRnMAUV9QsvIL0pto6vY5+MAE7KIkFw
tRADzjDX5fbMWZVwu7rT2TuMu5V6s6yUSdiJX7s5kfTB9dX1vht84a7AiN26MMy/
C9YTPGfzk0l1NVO2ZL0h3TUSo38JsxCI931j4dwh7a7JL3Z32eGeAOA+GCrcbEhA
6S6pJhSACAyE6KmmkST9MeOKQ7rHzN38dkjy4iEL3QjM4Tog6XXT6KAIYpSOcGN7
nsP8taQe0yBq8Lv0RfDV5sfVs0XsLF6NXe/CEQM5Dc9PBbgpVRn/bn2ungW5vXHJ
OogaPHpLaR481P2ifgmrb5MUR/EucyU5IQ1eV12kEDUGiJ6CA5xmN13Fn7tqiU2L
2yOxHXEQZWD1UZXyyz3HJ7yY0RGBF5I7S5Kr+fXCpdz8YI/I4lMTUKafZl8+ntxY
LqNGIf2eCFWMki4TB1aW+92J5vg8cWZW1W18xTYPkAf9NIcz8a5RL1tOKlVB9rct
IDkJ7ycGQXeRxFpZEh01VqfLKDn6IoWox9KPomEbyUiWA+hKdwW9PtfjS2d1apal
8vfcdHMntpOoOhi3dpaL2/QhAMEAfOc4ohy530Y0i8bUyKlZGW0MKT7qPf5nVDTR
oAaihyskJo5xA+3akS1NAKyRQSnHgTYu4suv0OBSF0zqtzT7SJ3oNoE2gGZckVRy
yrhyD4erPQmcKA6zJmpUTZP2QJUWa3BZ+B7Z5NuT2SKwfcjeVWVLIixRRnOb3aWf
pcEWwh4esZTFhw18XOS5GK58+h4BIgKUKnYu7Kh9Len19QT/m4y1V3qCvBEawhqm
i+GRV4tFB+e3FcnLCqg5PYSDIw+PjtvBatyvV0Z8Rvhp/gUUFChBmvlHjQm2qcu6
GhGxOaX+353RNLsy8rshg5WpeX1sBFWrSErHzwKs9BTvHJwESk22ZrkW4Qxe8u5b
N3aBlbMn5dFjDL2jtkw6KUrIU1JeOvenmkAM9xfGQYrzuqYM8gu2lRvHb49utwv5
ci1vL4qTRDNtJvPgZ1ld1THyh2rmpAA35Do2YDNaQIpjb1dRK+BbJcuVFLmZ1Ly4
1eyELim5KIwyZgNHN/Hmy90mDPtM8JV91u+tFaaBjquIW5aqxH4K64D7Ctq8mOT3
AEBQX7Dsw8wH3XKNXzFQQZf5mPPe7eU2ewPRar2VA/jsPRA5iAKrMexpIuSOQzIT
QUz+rEfJcfTpBI0nOS8o5uKVSKaJbH0oBkaMqodBiFRF2EaRtYRkVOz31kg7DmQk
JJcC2bjudnJWF2hRJSHfthnrUQlDI9+1UcO+CunW6U9DHPCxRIu+JjZHSceY46+f
DrQc0Lhx82W3nzyklHaOSnXL7JAr0xoQAbXZHLkT+Mzf+iczlbHnw8KSVmLp1fz5
7P32gJPxGqsbAtjAL9K3GMDveEOuagHDhjlnc9XkL2vmTT4/NxsZpDk9/F3kk0Ns
+6WVzj28vC7Pt0jaYSF0ZJBHsVnu0ZIkFOyVxCRwsEXka+1YKWARxhcdWLgNHXv4
7xzDm6KJbIUSHnA+dV7pZaIU31ha1lJB+oezfioUeWYdHyX4UpF6r1YzlQ9mRjw5
YpFoufbSl2DqrQltvwwQt/E0Kz7/D/XK5OD/mY+lLaYvfHdiYbRGk5FiF1Y/x2uq
yAKltPgoyAOA/t7I8MC7QjyGVVZQ2xSLUvpf1qoEK+srLhFu6lbsXtKl6NE52Sks
fMNfCgLo/woik0fGwfVzmpNF7vC2D4MPVkAiIaQ8C70NbHh9fUx2eqoS8SOJ8S6A
lcyKXqNuJvhelq7y5gKFfVSuzg1LY9pD5DD9GWu2tt+t+9puDxXWr/j5zzVcL1LH
5P5wk9QuqDN+nN2bLQlUZqDvuEidM/B61QLti+Jacyzw24KRMmXjivSKjWL7Sa5D
8JKS/g0v7Vpccqe5/LQxzinJT5KRJn3/wnpGehDOGySYz4yPXY5eMdf+XvozUmvr
ztXZum+QoHrav47Kv2gioZNN/L+bN/JVB08Ctx+4LufYKpx2137g/0W2hDPN0R+v
L+0B/Vcl3OIFDTuaDEZuaDh9hwChBBVmbORRBHsqP02GlGtAJvfdzCN2J44fcuFe
qEa8khtUUUF91iCTuMxKn75CX25htCJhckqsfj8he/wcQ5AKPapYCCHRXcwCMQAA
WS21BKvTtR1M/zseuZ/ngjwbk4Q4D+K6118cUHMvPTYdAXQdwVjfxUqj+G9L4a0w
fGTcqGtmfgAF97EP9/uDnUIG3yKrWC4AIoupBHEI4k6/IIQas91G2gTfu1Ml+kkW
h145vb+Um6FWxoSyopvPCCfoDLD21jGY2CqBvGw3QyluIHsTa7h+CLzv6XfnF9Es
nsWZZQ16ypytKqqstMkaT2FnwwpgGsAx+1jfM2PahKRRIgxIJLdgLFz6Kiw1t4TI
DamrNgXmeOq9hiXCBts2H7yhnjey4N68rDAIrRyM2fOZlp0Ub1JacG3RV6ZAm66q
Bms84GTsG7BwDpgq8tn9coBhVkBmAPCkSPdY9kcJq8c68Rx1J71B9OZKveKeaSzs
L5fOH7z5gyj40YXqkzL6TRaTBYi58e/LksUJS7CufH6It15Mwq8peag/Rurv2e8U
95IAUfhueAqCW/cOAdeUUmsZSlldpjRNTqSlPGiGZ/4xunm7C+uw7idfYqo7oGgw
LpJ9OlWTGbKVP4kJRSRNCE+9FYpiw9tC3WSSNBS0mZn7A4+1DGgdQXuUxAlVDaTo
5DQ/vnwrwHFSYc50NBE4sl1Wz6BlfWUEDrenp8NBe7cVT1spjnsSw2U50fkWgfh7
AaAD9ZxE9KaNnBZjh8Nw0LlQTs7d8vT0ryuhti1zpCj1Ylfda9eqGZtaYKYH6kST
56D1yMLkE/3mTKFImBqWNggbsztMThStM/bFSlWKz6Poe0PIRgnavajcIlJfcsxe
vtqqLZP1OaDjlXlWd1dEOo2kU6Wp2llRJPONAVAGq1bdqH+RLoAmZJOBOwrT0Jg2
T9ElWS3MMOTI4a0EK7ilPQhBGyvgZWJXgfoGRnYYa1nTqHbgt2X3CXZSEFPgF5Kx
95h5TvMdN+2Zk141qmS3fskIh/HD9TIN8j/iuYyPev0sg/+onJIjdPl5GTZGrd+z
RkPHcdOO3c5eI/HR2empfDXuCHCAGCVyGG3woRRx8phwjT9xN+ejNqF9XgjvHYHA
a5uAMCgGyf7A+6WQiaxvO3qXHl0jRHCnxonK81m+cYyE/AMd6w/phLWHtoyRlmzm
Zb/3oMuBdcpOAOcNI38oY8W9s+FFltqNb/lImp4LL9ASIyMNp87JuFm/Uz3h1M/S
hBLpaBV2tBsRinLsuMGN4QZdPFhAlzmSt1Up7hEvu6n5f1TPTqKC7yJxp4JnPdlF
zjLQ6sgUWA2d8PFnIIWo0qZ7IM5IHu+u4zl5aQUPeO0CUZ/M5196VJ6h8V+O0C1K
ZKY0BzGyUTMLlBlL+a8BYkVxooVEWtVFgMfHjrDPvPA9azqU1JlbolI8PlEdYWQ+
kIszkos0bqQwDLzY6GQmb2yWCh1xG92DAjFVkeGfDobv/KH+ifuLlaD2rtwdE2B7
bASFeok3TVctJ1GpaQjPM3T91kFIq1QSPsxyhOM67xJKcs4nfpyHi1NaLmwfIVPc
ArKaN9vi6mG8wOWMLZRHyVStqnHQrubOjSCGbQ+afDmqm6P+CQk8N18Appy1EZuF
q7eeusujNG2zA75kXO6wCFMSvtckDa1I26JcpmwblDYFW4k6X4CSmzNjwCgwwRCg
Aes7s9BrlplzoouWLpo4oqRIQ3A9aW908ZT2CfrDzGX7QeZ0j8D4qOII7PKPGqi7
vEvul6GMsP/0my8cTPLss+NDY8jChtUJhaq0T/U55LZvZ1QdhEujg1HQs1LghTeN
Zk5GVFClT29fubBbcRcD8enz35VuldrQSe8Dd0orOqUyNILc8bnCC04W9pB1aplN
Ct/ArdQfS0uwp3z30hRgOvNUpIspzqfHITaSSeKiQG0z0d5b23cpK+gldk4g6IT5
tE0BlHmIrnmhcI8GzNkcH8bwrxQJSaCCAg4nOjeyEPNNUapVqprMyqfzlsvjm+6h
KpO5/j5bZwZU7+nF65CzkiHxSgVcWaL7gOXMFLxObZv6CH/azSKVqy/FcD5xDvYk
95RdF/BH8Quqw8NgDmAts5ikv1f3HrtjdHBGqvX5hLAZTs9ufB72+tlsIIhU02n8
5Jj8xyGWp4e9OreyAzS0khM9tYdbvs9xwFQJpHZWWyLwtLJzCp2lv74fZi3qyywb
KCqyTTkZ7+gLu3BVJ7qUVxfhHAHrCMMuQdXrhvqq9kRw31By9VeEfrwB1XWS4WLG
NMkk07sWiRKaOn4d/AaZa5GcoDSAzNrdP5VWlrnug+UnXakU2RLfsUQAfvV+3RWN
r7N5q+2Zb5sewx33PnZzymw1dq80RTI+UH4IIDCNiEK1pK0VotMqLeQh0o2yySil
eMXwI1zUD0CZsMSmXa2tDaEal8DCYH1XL9DJP5otFezKPeG4PLJphg80voS04CqN
tDU8EDmR7GbVMEygXsd4FeRoiAe07FEUlXHTYTk9sYk/ZUWLnvaLLlslZn5Tj1Tz
z7+WXPEnqr7WtFFISeHJZ4BBFN2PGyy8VFCDdXP+DD7Q1HsQTZSZJ+lxNdXMzT/m
QZLjiWqjcnDG9uRFb0D98HxXyEp4n4m6VoB4fsThtRImskN6Z0GSTCf5/BKBipk8
o9ZopgwAzDgHX5JmtYo0Z5Gi8L3W7k4dHeHbY3e+vCEkJj/MjtJA9G2zbWSsZ7fN
+kfe5NxJ4cxVETP+4gP+gDgsuInj0QAGfJBdo7+FQJckxQlmZ+26E3EBV7MZyOvw
lAbTTabqzn9ivO4mXm+s9/ZIZ3bTIXakEBGZbeXUiJWmZirth+sO1I75RzJUEeUH
F2Zmw9g1BfHDJxDJDj0uEB/g+S2/JSfDaQVSV9sh70WRwqiQOs88Ganh5i433s6S
fkkPaXqq9wmNX7jEujGJOxHU900VWEPVTM1s3mf8XEFpZhjGq+DLEnO5A3BuSy6i
iO2ZQgj0H3oq3H7aKNkCipj9RaLvPUY8VE5pDqKLr3zIgRhk5+FJs7vDZ1IYbkNs
ukYCcSZgc4Kal60eE9VbRQlg9wr1EoNvDGYMk2BkCiXWPKl4oNCIFlU0fjlWgvhj
mq/W1ZIhYNQ3gS+A6k5ncGt8Clz1U4qzlcCOCkc27LvaddRlGqvV3IcaNVG+F4uY
rSgFv3TecaAzENkHg1dp1VQKNxso1V2/t44gm2czsV7Qz7tJTLElc//ScklVIPUh
CXZYgq1+V5FoCglnZKDCztEhECYeHqfeUp5d55/45nT42T2kQbvw2Vho92Qg4tUK
XoP3ypNC53O+hIkiOAgfn7Gnq/Ej8zDWZpSQYAPpcubvQ/+4kEIpDcH4r0AFToDb
k18BVNsb4VLvEKKGYYA0rf0WpOxSFznPwhDD8NCS0wmCEgwLqX89+uLUmrz6kB57
Vfthlr7fplzg/ll5NY6shlo5HK3TWXdcDMa8qwa6RntknszSk4r4WreY945+Pvoc
qoJP9BhTRfQZpi2jbTG6SFpuTcltEJ5QNWSnYnyW3vcLYkn5P9HQRK2jPeQL2feX
mJfBFLA7aLfjRehfQtUmn/hWEtILf0lQSRiUq0okt5CywDtNoC4ZV3TVZwjaLJb8
urWZwMtwqweCmJLO/PdluGvUZy6NBR9p5BnL5BJ9Nyg/wY0YllMO6KdHcv8hGwBX
LqSxiZGmDZlFj8jW1Ppg2gpylFWAyLPTxy0eFZNAO5BiKUdmQKyZu6NrLycrbxSW
7d++fBk5yiR5ojKhWHLvvwYHyztJfNvbfxcbU1zxim1QRPkOPVTrA4QfxX1Sfyag
iZKnG0u7dt4bD/x9EkPnRiNGZvF+DZhdspxSqsQ6xtN0IKQa1ChxuM4khgxajW24
YM4ECdjyVjVlMvO9PPZ9KRqwxKVpjk1lfGTQ0HMgmIfWaYvZtebuXSS5/iRNMFtm
WN/GrdYM4XJVyZyZR8g7B/pFWoxC72z0w01BEl/V+FnmP4m9WtfvwJNr2bQEYJvs
iOZUa1GVDGxfg+PR4ymnWS7bITJpi9HJPi2pxDEHyvkn1CRH3EyZduzM3HhC+5aX
6Uehl96lSna0+aNqHFXIv8vvKIkUanz7PaAvtGW7SKIac/wVjQTsJmptpS3h57E+
cNHspZRlVx715w7fL0Mu09KkL2DmACoFwOKFDwedc92EsphkDtrDk+QnRJm/lRaR
acLkhlWBYrDk4xJ32uPIDdcxtVxpGlubUda0RYY1h6HhOHKxnnWsV8AksB8tSlyu
mPwm82G8g44jdTZOxmULSy16GQG7c3X2MHRwceUoKkRd8WIYJHsL73MzPySyo6Fj
iGzKsdVDmvcBN/JiBOm6pOLKUzLmUtDDzuhsWGL0CQTxqevGpKNO3hE4vZH5UTx8
wilrx1dimu/ScjrmVj5BP7wT485X+VF1AMuZqKRbDtzzhzXlBAHQ9snY0kQGJChd
WFPFdfOEAPf4a3S93mPlCd39rv3iBY8+Dwfme34kbz2NrGZtoVgHVJzLGQ+85vrS
2ruYHyGgpf3cRcNP/XRY49yaHJZfofdo8Q+7WL5VWC8YCN2FcyPkdbRhPYiHpBLk
ZpJzpYOwJv2hY8zyOsXPPbdnUiiGXOjzqucC6Qk0cNsx2Pm+w5RD4GAXl0bUXfi4
3vcI1jNBp7kLYEOcyqFGOivGGlzf8i6KYO9NyYw+UQjv3PZUIzAAAhBwx+acH4oP
2hV6F8hUbKqS3SRnu0kxaf8ceCkn0M4qlJOMPxmLvMSa/nkfplYL17spmqhZw6fA
0c4ElemEmpdQ0Ena/LNKgYTWh/3YTfSCivgY/52N3mHTsmWXGt2Sja9aMpqYilkG
OIv4WOPhdPUu/WEz2UZdORzjOfazXqTG1GlFYF83W0mVOoAP4PZRVz1tOVlFrjlV
1QP4m6tKNQ4QB9qtBfo9lDEGsbWKyYFPV4KtYBSZIoSAyqhCPhW8kHCneeVsCupO
4Q/bqZmzC9rXnrZac9hi4wRvJmv8QAIz/Vs3l2yYiT5tHNBqFe6pb6X39/Nhn7Xk
JMHoV2EmEoqCZHL53ti2W8pM6Sp/pj5N8B/DkpgDViLRVH/R+yMb8CIE/NZrl5oO
adNCmW9xamJVnZi79dbLaCdfUQbJ0aNLKJ7d54Bj1E/l97u0iq2mqAZABFUzFv+3
Vxmyv1ohEyvJ31h/Y4rOVv+XR6qM3+raHgH+z9L39aYmfKhI52Ult57pq7etSe5k
Azu3lmGvPaPq6ar/VfG7e81ihKtNIEzIYWDl7qxLkwjuvvl+46yd+XHaXyFHrmXA
o1Mwwpao986O5sqsVYPo0UL18LIJOoUFosdYSumuG8Df0zWfwdoY8IvQUUI8iSxc
nFcUroh3J7MHwMZUySI26HZc4x1hZabO80RG1rN3t/M6P9ka0Jxy9J4YXyTYrFFA
XRQAqtmM49WgyLpznriDeMpo6pOgTwGaBZwoQEi1Q4v27PHkT/LoyiIvs+2UXLyq
oBoBVk65bwKs/8fs78w2JagOhbVgG4Qe88RGLk+HkAcc3YmnRzS5DqmA4sHldpEz
rDYi0/ZbxBI1BfVoOdK4SWnB7J1tL5stvrI23JDZwvM5NY7URJz/yDvTD8UhAssr
5NS4W/psqizfcaeaoU/JI+/wwnSSNUCQ6BnePVxkbDrDvM0hWd12/0eJurcugAF4
O/6YgIJpA81Z/NAepQY3iVO7xlyfnmSiSOEynVh0O0v6747eyaRsFxFlMeXN0XcX
t1GCQvRqEkcXEUB6ZbFVtVauFaXrXZwbjA+ND961hO1iglgDnZbdtnqySXWU4k5f
Anj9FIAwqubtzXIQOoSP3/w43IImXrinwNwOMLElNAMG4uHIUcnRWBTMwVuvi+GA
vPuO5VONEOVhzxZlNJ5HYL3cpNys/KLc57k+qIlAiMLwVxD3Kv0SJng13yhnQGr5
uTN9zBYfWKKpr5XDSjb+GStKz/yZNDyuCzMTWSIHR8o82UbzYMBl7ET9VBVMABQb
iHTBrZL3N6eb5S2qyt0Nvf9wsAFu0wm3wMEkmId081zxHIrJMMRn43BPDmY29DoZ
4TkiaxMpcsqm90E1N50hfStjry7cJ7aOrnqATldOUh5uYWdTnRLfsUMkNEfpt9PA
eIJJNnXv2HGgD08W223sLbTYF4bA2npUEUqTB7RHBO0Dm2PQAFSyNB+2aK4cB2O/
NpsYX/Hbdrqg87NCDfuNsFFmsce74HBgjbRd4AVZqIiMTA7MFdSnwM/ct2dpPAWG
td8uANISqzaB1ItDZpIVW/0PC9Bx7wXZ2Zkw3QZvEkt8BDYr6Rq9kqQHeInOJk1/
QknmmcM6exSsnIWmMfQ991z/CMGhQM846fFrMJBGMAeMYvOdKvxBpPVj/j41DQHh
8qvcytjVr9t6KMdwV/Kp2z0gquv3ZPB8bgY47J5v3r/1XJIfu0A7eTfTaY00jMrU
GxRInDgzgxgxbc9jdlOb4qKCdQ9hnqpXeHdm/gRAs3xPbnPnQ/dvG2US0/d7ybLw
/VsxZ9hvwN3i/szLPAeDvRFFhVLV5DKzJ+0e77lnG6bEyRsqBbfSnznZxNW8wZoB
bOUd00Yrme7YbxF9Le+gzBZKgCgB6oYLBS5q0Vo12e6vXVDt93rGtnz5C4l85J4d
SGf1yr4LFbgVLLElX64snSHB4BTHBqnrUdWkVV2fEh5y3GefRtHgcFMNBZr111+K
Cz0NCip2VF08leUvF0wSIwIexPcuj4n+LfRyeKQekXot041K/8R1o5ed5fEyckV+
t5seu1kCEhHogW4vo2j529P7CLvQbPBoPfxjUx7iddZYuNkikCVad7hfMvchHz9l
f88aJLcr9CitlOifZJvoOxd8LiZc0l2o0qxunxA5r9jQduMFBVKzpw3eUN2bVqQ1
hCXFZzHCOry14qPrikmqzqCGpVMNIwlA/H2m2JmieEtD+uPkx9aOcTeqQIJJSqWc
MEw7ZjBhC7KHf63ehmTYYkzJdjRftvdN8RQFpaqoJIhQ4BBm8aDC+R0mcUOctlmB
uLB0AAtWlX8glHu6Q1E8xE0GIDe2nNyYZXGKJmohHC86kvV5qVqKUtwU0LpO7c4C
dhYNVHvjCu6kdw5xJTiqRYa9AWmtFtnYk/tqW6hICCtCftNcqQCpmAJJROchUump
AyyDRLu4Jite0bs8M1iG9dzp43ZD1CF9183KTrcpnPgrVL5oF2vtG5jmWJmXZW7n
mKovHrgrxyefJIPJehdkkUpIMvZXFHXy8WlNITzYhz/PKKjaLkfwxPkJ2jyNLgIm
DC2T8Ir6txeqH3KTQYT1C/HwrPt1sHRhXFVp8wSFTjkNrSAkkPaSYqNkPuAjeF/+
04FuwmT+W4wBRG+rdUXvlmKIGRSeLuJef37cnRXyBcIQDhophwwFUAZiPWIpTz2K
tiA8UhXlsrRTkyI8s9hBpacU6ojXhGSNlNRe+X7sTIX2oWCMgoGfVyCh/YIQQ0W+
j0pc/k5zIywg/7/VTs18G7XqMPuEunOwbx9wiAhvDe1K8OJrI8JvAidLIvSvUHtU
w9549kEgB4LfV2Q5SfMMmLFoBo2QfM2RKSZQfeq+rIXyG3uxvRkNvjdWyAHhE1kT
MdxhQI2v/BzWPln/8MYvN9SEP3F6ETHMFHYApAELzQ+i76ZnELjyTcS1KmIpspq3
6bbrhzoz0qmAGAfjfu4KYA23agit5Gr0h37+psPeFUlYhrtiSfODWmO/d4vN68+H
22PjpFKr9MUwwUk0CdKRtvDdr7FNZ4kajz55AK90S4q3t3vo6xg73lsLlcMGoweT
9fiYkVGCk65Fgh6ICrugoob8n3/CVjYecWCPb3Q/xzjMeLFolxpMSe8EKhSzWwxA
VZ9SeplmOpeAER3t8lneltWZaV9TAVeXLKflv7pTZakRx/LrC4M8WWMgCMZnckBa
ECO4k3eRF4Q4YRU1XGtwQvQp2+LEJEcnANBODm4doXAWQ9p20CYaTTaYjEzrlRgV
5TyGqkzcYzFsA0/vv6O4W5OABo3fMTw5lnSBDBaFzBdX8voVha8oN468wcin7gFa
GLT5geT6guf0tALAb4tOHkxWsgv6uB9LO4kRKwWrdUrO3spYL1RRQAMiLIznd/xe
lpNC9xvEmMfy/VsPShvAU/C7sJqeVyrFQgZKVdYwcrzM1APLf98F6aLeLEGwdD7X
lLnCpbV0+E5pjnPX7JrRJNrltpnWjotGnt/BSSvcJmZMkLY1nNBJgTV0MxR/o0T6
XLdsijrX8aguqVZe9OLB5K2Kl8AytwWAkFTL277EZyc7sWIWEizKCqcjeiZwW0F4
jXvV8eo/MR+Ji7QkVE98109sCcPFVYKqrx6Awts1g6wX8qxv54IoFfHw1tZmMM20
H+3xYU6dgb21Y+3l/fSscz8B8yE2WD1/zxwIIZNXhPHs1DjB7gp8J5GUEj6vrmkj
5E/yVBADV6MKQiNL8HjkUtrfJelzRpyBj3FBrg9petcRAZyzUrrf5o0/N85IjCwZ
HQrAA7O8Ksvo0PNRjFV+dpHVVslkGqjp2IrLagyFpBY5Po5EpdWuYew4g+BkKHi3
ceObVuQ6u647M+ck4vW08uRzzd6YnDSClf3QSg4bZ1vWU1a7Lb0UjGgbWcX4j/Hd
oVWe43AZDDUgvgGGfhNJSOyIAeK2XN6dA54PQQEmYuZ3b2HLAE6QM0f7ij/swMD8
Po0kHtt504D4H39RKJDthN3Ttf0kkURqpM/us6FLwrtd5BloofMcGoVjfeDBfIVI
PsMDqI9gJCY0bP0diWcSiKBUIeL6Nrwqx0PncqdqFurbh2Eqt/jerX+piEJzgED8
k7CskbjKHxOG9IyK2y7LHRdu+XTiWHJZZQMyC1t7bWedxfVUgga4M3qyydZLPqca
uJFgQLGrxH0P7e1QcAAPodhF+GbCoIdE4f19IH2v77Uwob4qaqsbR7taz3ysDaan
fEfwXrqdikfFyk3oPFA/aDV9wS5CkdpiaSjBnOPImKub6KT4SZLXpudlr2JQbmwV
JeId/kHJW8mELqzl5xGlyHDL3MLfwmhrOx5LZ8by3o9MBxQfI6erybT/9s/VjKey
cwFuxTkmT7jHO5xzSPo6xY0NvCAkcjWyqDvGMl2J+lgX0viUWEEM0biEu5WGWc1m
IWWH3iir68GONpKt6mzH0Z/tBO+9+hk1mYGw11mM3GjBKflE2d9G1hhws11HgLcI
aHNs7AGDLjKMGpqb8/VcVsd34eOC1uLSdeoDiVenBgP9zm4hSmAbtFmUtfqVFpRj
Q8eyeTZHutIbxHRM/rF6K5hzEiaYdn95CyGNgn8zPfaDAsib3vImsiSnyo4BWXSl
RrxVVfeDRlglolISpEtPJ8E1EkbZ6m8gaR1zeF6ArmC8Za5VOHV6+hFaD18gbH/8
TkRgKrDNDB7eIbct9D/oCJeNFBGLRchXQiSubzbWcOMbCG2k8UpTXYkNCHEL2+gJ
85ju9/ETZ9GG9uuuXh0V2AfbcbJOTcYH7F1ZwRQUMa04L3kshnKTjy2zIpj1n3Q0
vpXDhoh81CsJ2Id2MmTs/lSeJ7+zsayldRFvRimWuug105/U3r65AjeDDi/PXn8Z
f45DLeaIS5CT6HZtw2yBL0hP2fdfrPZZJacpcpwV8QXiG1e3Aas3/k55wO4QphxR
1R6iubeuY+buUEqRnkOXWjV4TzWxq/fqRB7w4iqcNCMAD99S57TrA6hMoko7UaQj
xPArBMVwQw7/zB3hGfCa6P3bKIOrmCjnS+eruFcICQDwe55ftBn6bsVanlT0xe1B
VP8rYGQ3w9cD1G4mODdYtGVXYi7Rbih9hiGHDCq+kaxRtWTSgxw3XyUJzUPhi+IA
HSB9aQZqDqHEpbdTvbsyp+c0zVnpAR5UYXE3zXHL+bsd7o7gu4BxSTtQYsI4L4Sn
lSvwSnhPjeERex9kiDu3pesaa2vHloDBjJozUSw93tIh80X7ki2E4GaoP/Ajlbn5
X62FkdXG2bPOVcMvCdse3zD4hbTz3cia7TbOCjYEqMpyrxd9hhOxyCQ1Hbze6Gzz
l3wD/CGTRxOgKR/TjlCbT6dKCmQ7/zJZyrMFtZN62MQaSfrc7FQ+XjSliO5GaUHV
CZfEL6o5dD6ku5MT9GrdKXiHRb65iPn/Zu1AUGguqAPET0bQJEj4kfTCwWdBhDPJ
teXHXKEmCybehmcvr+6ITUlghjZIlOjS9b0BliA2o1CJ1f/dkxjmE9TxY2u4tLHy
lPy4ze+1ckLG5AgtOtglb6PMic7Tq/4Y/JPIVl5+EXRb2pw28XXx2Ies88SuH0qU
PuSGvtQpzceKuwRMDzvTaUwqJ55yfVNA6wDNRvj5S2FYs4IpGsDCmW32LZxCWVyR
3rW2WFkEZQUg/s3+aKmGS6o+PPSXy4AGHYrqWstp4tknXzMBC0cFBTJ/pXQ4TmCG
e20cEIsvIiVoDJXQXVLe8bmNkUp2gzoxpz3ydkDGN/LMrFmM28WERfInI4d8vWL+
htwytwZAcwQ6mp7tukVHYbyg6ZeOlUZ/rzeXa93mcTU/mufonWJ1GtrNavQAIKtc
aFGnvECyKCyVMmhcsuCO9knCB//g4bgDyssM0ZvCuFqUYul/fFTq/pPTl2jtkfvu
bBd7jdWAgWSbRdMBUVnkpQAIRvK956L/kzwsDbAYCuMrVbZadBoK/sHiedhDLfCs
f3w+rNJKgvso/dtRosP1DRllXvTg6uJ5VOoko7nnCJV0QWaxVugywtbq1nUyPh4+
ikB5JCFfT/q/L02xLMLtsVT2z0Zm/NK8wMIApL7N2RkfmBP9c0DMpwE9zFbRazcD
wZhEd0LnkvNT44nHkuV6/TBwGvzGuH94tIpmtB0tTg5aDonm3OhpZ+Ng6sc5RM45
hYafqmp/Vp7F1UWyEbCbnKmnxYuluPwFvdlA9c3eMuOFsQkKDua0xuEESZ7vU+/m
01L6GX7Engy3QW+qssRyqsda+saejKPoamaffRtBLGIFoxFw2EVe32EsnQuMoq3J
mXJKE7975HNAILw5kjtoc09znzzohFafI0fOJBgdGngV219uPaAKM8UOEQE7/T/N
9HoKb+GeqR6wJwmOUnUamfg43WzGdDm3wCTwgkS9qAj1pwNgZxjwhTktcIjybYP3
CB3v7lEawivjwxI1Dvb3Ym6zEwoUsgVrk8nDjgISqZCJhkdu4djZfUO48VP8EC42
C1/MuH0sQOComH86TsCx+5IBQd3erBwXt/admZYUQHUC8ZnZxSn9a5lD9ZgCRGuM
+mQ6+2NXnoQhj5iu9n2aVIFsEUWLK7EMq+v7XEd3kjRbYhU1aJnlTNa4Z62XQW7G
RYRbAcUM9EV3YsUt12HsT2zJ+BR1OOgnyKMi9GxJILGSTW8HewhfagvhfDRtHUx+
qYd0rzqGDXrcY+1P/L6IIX5wOIiXsEKJkmOoIFSJ3kaf1WQh0K1gq1T5uq5z0dHC
`pragma protect end_protected
