// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ady6/PwcXuDzMYpZpF07Odl9VkC8s+IZ4fi3HO4kvA7jYTi6mamLLgR0uFu1XLG/
ZnXSb5yRiX5gH1O7Mj7t547mt1jqKUwqerxsabMtLq3otwzXOBuVY8BtcN5ZdUQf
bML6Y9NNlI0WTe+rgblqxGLv4TeHgtDE8PQ6yYG3wWs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10208)
AH/kD2/EYXbnzjKhirypnJcG/iRXX7wkPTXrrQK8CymrueJRYFQrXkpjsIJkCb1+
L5kEwMFNpV7HqAsu2Bxh+DGmjBwGVBX6fAs1YMMWz6CfT5F06K7u9uqs2+5y1xif
lkZ8e1wMwLthItlyVZQjIdk7f/jRk7cRdxFaJPXBDK6FsvRTMj6d6Zq7GIPp8mDM
PTjHdajVzy8POXZJrg8u2mNsJ4YzF2kgsbwIBbWCqDtLZLp4Y3ygebEaSBRThoFb
mLcbezMuiGECX2GAHg/w05AxMaWAcIHZyvHiDG3vjvEftgaZCOZ/fX7E893zx6mE
alxaNiy9RHQfQ4YJNLD8CBPpGLoZ8kWBC6+KSD7AFiOXWT1gVQd5flKLn2dKHNUN
orG/Np6S4KVnQJcH5t+1WvAKRX8YZsN6q0YUkbxZnSzEqsigRkakh1kgh9EOiEIt
iVGY5F9WFfRyDK8jL53YWLKA5zfTxnX+Wu5TPyCTMunHTzKh97vnqph+OrEv0XgD
h+xR5xHvklMlkjNDw3VrvKUSsxDS9DSpiTA7fbTyQktlPTNw7hzy7Kg6KiuOZKXx
Pibolo2iykwpquA57UbD+oIx7Cv0mxQ8d2CK+EG6rSS20rx6TkugA7ZXZvV0NNqf
Drjk9zlPXk5tBB0oEInbs0iYAcIyaSpltZocUWFRb4C/r/y9dKGn49kTVLkJ/XvL
wJUaqhOLbWzjuhnnppkTMAWevLSluvpXry0eVQo2ZLfec4lpCn7qId3rB7dRCXfr
WsbKZoT7TdtHpWzPCbL9ZikXMOeBaZw5yNB5EREOWDPs6wLJniTj7+bmIU51UXZJ
pdJYDJUZ/blWXp8zAUb4QBGnGkIziQwaL8aCeUvfLCLObJioedMoCJLFMX42hx20
HZBR3TCQEGX0ltGKZZlhEtkOfQZuLA1u6rHx/maS+PPBbte3clYwQYruBRBD1J22
G0naPg6LN5irtHf1HqrNVl9FcjnK4zwiAggRD+YYXWf4YQRHEjmWuCZLDoqRdadJ
JyUd35X0TFAMB2kdmW1DBgUksG+2aYXkeC/zP+fj6850EX2sETbe73/IbRn2MXKA
gbV7Qk06mhs26Yia2Iho9M3nqfx7iHODez3KfHV/uGJy4OEPo3h5kPcpV/ALyzz9
9RVQTKMeCw+U9u1inlGKKGr6Qdr5QNKB7DzeZFPQmdi+wycIqMk3XefL64Di5qMA
N2aFqBlm30xJfsILOd/GYE8z9dSRkqp+7B/G31afezylv6Qc8PsIpawV5AyC06nj
MBT6cblut7tKO1gnD96L1m+Z4XGmqMekrtXKRsggNDqDzMM3ft3+ABjnqQSMdUvz
cBgkHNQ+zbKy3rkA2micdVhNA0830tZy0pH8SzcXnfi3kKSQWU1L3t/3iI0qeWme
pS3qDanNsCyLQa/aJaslQ95OnvqvyKflQPVF4of2mTtVunyHuBrB4YVsaaXi4Be/
uT/BbxfU74P/lMNzLI0MXUpWF7EqHFoyuir+afVy7bs/dI9z1TW+k+4M8ZyG4/Mg
eMaocn2tc9yueIGgvDKMNhMWUHL3x8K3RVfrTkx3mOa4CY3ljZmdXRjtMBCXYtD4
t63IHJGhjKeBJ/cXzzVI4sLnKpm2KxUvlgj+l2uB0Y95+C9aHEL1ZgWuu7VOvkkd
zpkWAr+X5pd00J8XSWvyb+f5DD0SFhWwtadRDYiP+mlbkNGxZPM4VpsrtdT4Muy0
gBJ/MwHG/lHRlpJFR4e1Y4s+e+CNN2XQmqH7YwpCf19og/+y6IQqoenasaGKFiw2
YCS+3NcQAkz0tAgSMhVGVaERaBX7zIbTOhRZ1I9MvlIYgmH+l7+cKTyvH1iRbsEE
N8ol+LQilx/ruZhDY0tNXGUyGUmldMFxyjYJ+uB3QYBrIVkMWzVGxvg+bdXVKRnN
OOp75ifQyvTF6iD/Fy4ujw18iaqy4fhwlwx2jGMJDguZ3VkvlLinFTIpCS697ftf
yplWg5xNPs6UZATTH81tXEAyIA8Mi2HguC6Lm1HSAlvUygPwpvKmm7442ZH0le3t
TqFEuoN5UvbPaZQI7ZLkCV1O/LsZjTNRxuaJYUKU4p8REJIV6K1GmGSURs3UmPkM
VY129rYle4XXUWYx+2xj+XWbuE4+AVWRaVlEC2G5MjfP0ktK9hVyVUIH0PRKM3jP
B9cLPeSQKXoBpK7Da8i6U/pmk+5SYAOvVuslvHjMwtc5KW6ubnR1l0r1XsttqInN
NjvfVwtGGN/hhe54VcHVoxwZFRmbsr0nqMY20n1OxlToIsDmzWBdaVTHQin6symX
REpyfhIGeqLWBnSpHVfDlZcOXE3FWE90MOfyL1ZIP+FsUMncFkT7JOzaqlPyjAki
W1L0ykoTYP3ZXV5VFGfPmnkncauS5r7Brj8U+RVbb4++gOUwZvYA2dvpDtc3EruO
M+npIp3Ai7BOE+2WM190rhfUBiF8gGbCEg5ReBhaCcxaDO1NZ2+JS8iaBVbTtM5v
kECUy5VDaVOSzPhyhXubb/OtnBmpZSEF9MBmnFlJWtjjyGQPjgBhYoxvcHKlHNLd
RbXCaCd/BFB2EDqfkB1JBnzNe8LdowrplDtbPMo4X1B+6bab8xO4X52GAI8ym+K8
Q8i3zBigeihPA09F8tCQ0iptt555qRzu8chlac0z6101QWyAwEETr9J8tizc354s
IOrsXMSLMyIgcBqcuAhhgxiDZwJP0ETlTgUgdCq/+ohNdjPJyIeBSJ9cfylG5gL6
oqGMNRVrM0hS0VQeoDY9yM1SZYR03Y7sqcH9uZb9gn6K31bpR/zaRGV9lJLuyzHM
6n6aWE4n3eLSQHUqbFgS9noyY6nRNCdrQ5I+8dBzt7P/yQfpEyUD857+IEv6PML8
0mGifMamjoH2BnGje76KYkaz5CxXoz8kqyli8OSO6gBrvTKZVG5RfBb1gjxlD8xZ
JxHcO1iBj6VQ89I/523e39DMIUBF6ICzmpj8eTZMnWO+7THH+8BfDpoMmOXCdRXg
yUhKLY2cRnnUp2nYYEGvtrhv1Ek62tYYjq1CHXdSA+WoO9HMHFCGWHqQ7ZlEhBFm
eVeRZJxK9/ZHQEEqvKDDApAEEK4FLBWtQG8XtyG2E7Avf9cwS3VsfXIwH85/rmw4
5jAtoR09JXsoev5YJNlC3OoESCNz/NoUz3PCu7Uj/atGss1Z8kBmcMXOhjc0eIiu
T09fVO78j8HCNNz8Fct08/e+L1wB5D7zL/33bl1fm2Xff+R0VccqqCJMRCiN3WFQ
Epx2fCKFyjJbVGqSENrkKIdOyB18s+4WahlHAVffgLMkod9PFUYaS5hsjpzgHkYd
yFaTJo3V5r94A8hF3+lEeHNdGxwubZEia9TuqxyjlZzFXDWc8ALEgr6xPDquPVm5
UqEthFOPFj4fiKj3VryhK/a2f6bzep3fvsONSPVGwHEExtWEM4kHyVE4jWEzxk5v
UtGBNaPGQ4KQ108ieZ6ixXIt1hpCYjx0wdD0/dnpeZy4g2wPgBKisxYNZUkLvpd/
zTwfk23sXgz6nUvS772sj4R4NUBxV5G2gnpwme1JGaVxs/BRfCus4QJieu5cyYvu
Z/4gs65HR9gJw0yhF2cfbFAv1wppGZ9qiO+z4FZkVfmSbCDc33axrXQXeQs7h+gT
X7lXQuV9oUm2xx1rRICjw22xihn8EwcHtys/BByICvycx6+tLeuq8mcIgb0fx5RC
WCPBKcbD+JL/TrfJTxzzqU/zK3WTJR3R4fqDQm8uDkfAXbaanYyZQSP72OlEqHWJ
xtBjxv5DEnj/i36eoI6r+KDE3actp7GclK+NH62EM9r1OJrDk/q7Jr9tLYcJugNs
G1DHguVO4eecbTGZk58QmTNX69FPvre3uO3xlvY6bQMnLHw6TVBryMmmW6SAsxsr
DWwU65G/IPji6wagReaduNH9VQIurLLpuLuHnhTGWBFjRNNk5PLr9iew329Y7Ib6
se7Q6siHDwlM9eMOT4dRwPUJwUeoRM6aHidvuMNQFbwxMNtVm1Tva107AA3nh0kw
r5/huTmBNkKNPi8eoXBz/vNk1KVUg6UjJdgfCz8FkGi0znUqaRZQEBZXusr2HRr8
9eTzXfHY9G7OPqHDhNEZ34HmQy24EpYbBjrIF/RiZrsYEQIkS4eOHwYYg0OF/0g6
JpUVmDdbI4hCxWxjFBP0RPV/CJoM0wJE4996LkDZIIxNrIQVCyAihWpAjWOY0kAf
CbeSQGjQeQEx6Cpx1+XCViIoSDnw7ds7URM9IblSKS7qW10/bA5PjXD0Ygbudq/9
gP09ATKR+MSwLLSG0ouKu+KKoocji/oi7GfMv7VtQ0p9PJY9nKWl5QX9dbqURh3N
wowjKjlk/vYjjjvuZ4xItL9vMmCH+FobU9fiyWbqHxE96EdJMa2PCHZSbQqmUkLP
TaU2T37XrF0Lg4EiWC6YZRnyJZTzA8K5k6L1djsGCFJwuUyF3FCPeQB0u8Sx5GBE
sTyHMAZxZLE4VqSdqe797PxgqTM7/kGsSIMYR90xjHzxrAzTbcPy6Q+vrVVKf3P4
wLs2fIyyU4GniMwFN6IgmCWafniIuvmyA0Ia9NnSndUm21CcBsAblzsy0SH15mXP
UMkZofE1Hd2me+jhl3iODsDKT9iA3MaQ0ziO1t3+Ula7W8SLjJ24JHCvZFdBy7Ok
VRGrQqJJJ9MRmV3EmT+rMypHjlXcFbJuFS4CbujaMNGIEXwjenrc3IlXQYVplRvh
kSxNjFNESpbV09X52p5FwaTQMpuiRlhncfHsPlm1XovaamImWOwVnjfG9U1R804u
/jb6pu2fBbhLmlTxIrvEbl1xHlLUIYKaGNGa4iHwWK/nQTirHQ2vF46mhXtNwcwR
pFor5Wr9Qyu5OumZw+7NEs6jALSgnVrXo1dp1e+IT2lKIan74BvNduYcumHWVX1G
WDfQx5S8bymbOH1SraF46D3/H5mv42CIORvC/WoYOc6FFs3NdsdcmuVIrPxjwx2B
TDUDX4Xu5iK2iNlN8B6z00qMqXG95fc7HTQmpyqgbNG11QfHIp6NA4+N0uTLoh1E
RBM+DuWVpiMF4CeauRajtO7uEN2aKQueQtIme7ULmElUUl2uYlaB/3ih3w7scDWF
rutlTE6BdSd2V7BShro+yyw50rf0mHT25SkQzJFNuEp1ygO3ffoStNNStGObGjxb
3novH8Laqa/jBhk18syZPxF5FebP1XlN4VB9zByWaJUqt1OQz24oxsv4W9FJUAdD
Ft+5v7sha9s5z3/R+JDNo9TssB3PU+l+wA6OmEIkdzsMqnfCkhPm7/wkrE5NOhDb
YbDgySom9CB95ena3rFKEgtE6dxbZ3NJp38+WaEwQD0aPtQrQtHPbw1+JPFtYyFN
bDza1Zcqy3s22Z6zghbq5UKf/+EhtRknpcA/CtUlWQlR+aYala0zM2cZXFH6anZC
FgnTuJUWQ+XO0pAJO5YPUJT2/RgLJtNa1NyoMBB0V0I9LMUBarOj+CRI7uXLaGzN
D8PxQ0qqWkDxwl6OqjcJclj/gpfglZf2bxlYrnwPiPruvZzyxKo9JIWqkBn/1TvX
Sk08BnwCtZCunWXV9Bn1Kb8AuKBZlE3BuYLuDubGf5aSRQV/nyWJz6+chWvezEDC
gQfxbz0towayi8h4OARnxAjomgN9Y28lobTS2V+fQW2PjHdPR/P5KP7uERQBU8cN
2I8OVBDHG7eTwx/SM3rZD9Pqfi0dyHW1bbXFB0d57pwC0IZpQa3bTnS7iH35bVpl
unvTLesIgO7MUfEZeDFc8IF4rGMweL1yVYu6XnqrBynmrkaazw+4B/XkFepcgxVE
TtNhXGMcgPLtfnchABikAU1CXQpHEg2ZRa62uOg8UIZDRUV2fKrYBX6ijRrJcaaH
VseFcjZc5Zuce8IDsK1awPiwoDelJ/EdKxqVW+a9V7cDBcKL7qZD+0NanWMHcWV4
USWil0+6X19kwHbzW3k2xEl7cF7oKxKN8xb3WjxTv9Ba3piPevXNWvesCkKzmCcB
rW1UxHGPOiitkDyg3d8RbHa9S58L4qUI6Cuc5lw3A/JAmSdT41oM2MYs3bFPU8in
Po1UB3WNeffd6hgGCeGmPaUWZXw9JPAvXNfqKli6Mf6WfNgotGpqjZC6bgRgRl0+
zQXJlJZ/Qjmj8fFSa37hPFKtAUvQUFstoRZmrMr8EwwmwJMcwki3Do+6Et9YsgrV
MbFtcknXpmDyMV91Thjcl36HlW47sXphbFPI5LGnXiJCaYoByKJUzVo2B7ALPagh
l4WyxPyhX7OVBgOJoP5pW40tV+/hqzrfZ3jdGBBtUZsLKw9Y3rkrmCqB7/8VGv8M
sAmZzOOCkLtGU0xSnnEc4FNXyTRd3w2KTuXjgy0UCpXI5jX5yH0tyMpY5/9Wo+8v
HwbJlP+kwXJhnBKOx36PF6+xodeejPtHTWmdK7xapyx792IY6trpUJ+JySCy16K6
+Y9VT+EDkE00nddcgxH56y72W2L3EysWTD+LG50sVaV9/uyZQYGQd3C6ODb9/oEc
dWyzClAhsf99wIWNtgP7GF8ELVKwgI5br0gj4LIxoKKqaTbSQ3DbZppmBKGLsWZb
p9a8OpdellOnlyNmi9M4uTeLnO+GZZbj9Sbkd0VPcCASq3c7v7puU6dWQ69Py7AP
KYiPXPpIk/MoPDCOrJpfXYfE7pOwgB3syrCotzagvMZWLpogjKkePvPzjNFcG0K6
thMSbaqVNYjnxXTyJAWj2Mw+ox3yDuw4pZAGPhjRGmoajr9IhwdW9n+dCmFoLRjX
eJUolDL+kDIAsUIZVHp60mzzB5Te+on/CDakjMw2JAwL3S7Up8utckeXgejyrIKw
1cJvdQHub/w3ZhWeYzGY76lu4wU1FGBwbPdOrzrd7a6UuFvRkonikRUeIII30gQr
jt37taRpRRCOTJDOt//RB9BvaoWZn1lLVrjVcHgdLHwq4djbPPW9xGL7ZH3dver+
BT4Qu3HC8tCwsPhOythpd4eD+Eim4Ped1jgsm4t6Dbc/K6AgjLoG6QBqfOJGGvdI
8ZBGcBl7Lqflr9dgITN+6rmLjKNrw16D/lKz/bscksg3l91RH4dxNsNBegOEvt8g
vmcNr6lZ/9QHOwr4YpMmXRLAlJVkLhCMF0oJfdVK845iZiqYC77Ik1GklEPSUSVh
QsERq5YBoCxO7rrhn6QmtJgG3W9bOxbwzDOzWVnptIZMlqawvkj/vvfm9GMj94HV
7Yy0c7+X7MO1vymqDN9PzHoCTPcKN6nRoMc0OSe0KLimPzc6zVVx/4qjDEbSRaIN
l0zTgxj4VdWwg+9uLjPql8+fQK00qj5149Vx2uL5DtJfFwm0O6ZEs9oYCfGi6Cjv
cSx8kK2v3IzVlvPLzWm2ySOQtlDIpV4bXmNkhpsoqfjMbOvGfxQ8vIDkmJd/FK/+
/ehVKF1wXvjH2Ue9Ngc86QAjC+LXqV50b0RuikYU/ax6gqKWhuIuNnGoSslfD1R9
DdFsfH58KTP2KdEgonvpcHFKr0uJOIi5ww9cwzrvKcF57R+yFSASSb31MWNOI+O1
gS9xeU+bHcDZSq/wJAejNWKoFBXndmDUOmVhl05PvVjSgg8liOxZzkvtxLlDhTPI
plKTPlAcL7i2xEvwwVcYK5ac5f7CxnPQK7g8avstZ1/vOCk5+W/TzmSgVoFZjt+Y
MvBhBDdOk0PkQUsaUB6AMauE01zxsyfDEijP10ALXlxROafbbcnfkCtHORFI4xod
z8rJGNwyxbzT4Rb/aoLi/es4chbyZ0WdTrj0m8twSCa6ytfwGqjBUxFFy/61cQnI
MJyIH33vGpCmFBixMaFdqe4a1pKJACGaJgL9LZ8GAPdztzI+74cwHvglPXxRjvow
C2BA8bo8xVzsZqFV9fOSxiyn8zrKXFswqm6isBvjn1pcgOygdslNEl2mnp5huj2L
h6Zq5LmKoqR8j5yJsqGrKc/IKKDmMO+bkKNjhdSil3oKkobknQLfsrZGM1ebNpkg
e0EGJ1o1lsCyxK4/69Q3FQCZqc9G0aqMa6aK0FDoNO5bTqF+O2uSVvuyAzy9rfl/
8jicCg7YVmYDotCz7MaAnTkSXT3KKr8gjb8ZbFYw/fJbRxFRJkyZ8ZM7bo7yGHEX
3zapuDxQdAvNFGbJ/rjGbuzruKo9FZJcwye/VtDH62be310FmMkVtaMR27VcNDDM
FWgiLyzcTc7iOaBW7ORJt4F+1oK4uygg+cjcIwQWEfcnUR4n/6qx7CUeh+0z1Jnt
9zxiCcbeu74dvu1rV55cEJzukXLprJtjj+nq5PIW1gLUKODu8e+CKW2IZSjENbx/
+yNdRz1GlAEsJz5punQy/kpx2ABDNU9Ty2ybN0hWicHDcyUc7/7Ej+1NABYGkUGW
VrW8CQOP7gKxt+4hTOJlfUWW5nPnMlAttblPaccyejznqGxupPd1Dyeb//1MY6bm
56atY2OvFketZN5ZFfUAkX15KW/1OPodwP1fmUL5y+pmH8oBek4+cKT+JASPmDa6
Ox5xJIyayJ1hEfWj9pxjZuamRAy2ovBsu85geQUWRT85d5rmNDO4kvnRamBIHXnO
1Tn0C++MNfF2CPepOeWwyMpkhWCW0UNvZmSpflSlTXCATRxibOBVc8OUOBTeJ+Mp
kzdD9ngrObaTlLuw0a3xv7B20c7ZDjnkvayuT+H0IJ7S6JfmlTxsji8Rf9Zmrv8d
8xayxQYn7alOawAc5P9jVyAxJElbZ5EHDZy1EMnoV4mW1IBS9ha4mL+YSzbqjaaF
sel6El7/PvX4Dx7pT9dh/5SlYmOOgjuCfrd1rxUQZe/O0fgtNQ4rGHFTBz/OLO6A
pNoQf0LtrhwK4QX4IWFWEkLZHsJ3Cdz62843NjETVjpKxH1vpb2Zb1qAeYHmgJ/V
uOI332GKm0Lwn6ZZJ2hztFxhmV9oFMS0oVxQCDNsEo6uRsph1lLsOCv4wdbB7X/e
RSmtiugIZNqm+pydaf8tZ49FaA+7ehLXAq+eNSWOAY036Yp05GwjgnuAB9ZVCbuC
ZpsSzWoeNPtCI+GlZz290tm1ShK3Q0yT6ZO6AE6PLwZAokhlscYW6VTUHwvgAjyZ
5FNnKdoaxihg9B6DAQM9dKn9EZjgSZ9sTaBp0z2hpOFdtTPK7TyKHL3U1JvUTgVr
gKaGqtyBaj/v9Es0R4J2zaRlwDRsSwL3HbsuhfYV6eO9wfKXtwCq8Ehzu1WGM4WD
8C2x+huxTSp+TOifyrmYPeLGLSR7iRyu9+CYzbpM4DBcK97xvyXaj4urkjPBltNz
gaXsLV2myT/cQvJgdXOsfMYbGMZQcc13l9V9bCaEWkrdSqc0NYlMF3T3QgoxpsXy
r8AZx6YeIlm6cXcOqSxzR1Dk6LFBDRkuy5KBQR1UY6eIP9BcKMplQOlXcgwoaOz3
dXyYBgVvl4H8kLrw6y5MwMK5jZv/F7rOeLQbi+dNGxmp2x+vbvEpjkqqsyrjmQFp
3+CptRpB9Kp7ws/6YQVXkGW3rVVBY4WqGoAlu/YJk4VGjfXuTWlrj1DL8i0JEbNB
TOSeTKwhhyid9DU4fi7yRmO8t9D+SCEBIskrSfys7al5+Gt7e1/Cy38/l38XeNsN
Q7ru4gwKIlyAqk1wRJzVamNwHI9yVhc/ouw679I5TAVh+jxLlJ/2UZLygXw8OisH
sFKL/mao1LgDBMiZajt8tJBpLFgAM1OuKMr9bjLIUONwJeuhAfoK096lj2b03I6R
ElXa3O12fj5FGfDkv1H/D6+Kanr/HTaVVa9BkHFPh0xDeWN4sErFFLsX3Hgv/FR9
tcjT7FklAgQGudG2mfMB//U4RDIQBpoHlVn0Z5e5GbwsxMHCwsDjfL7tNkQTNKwy
EeRt207eMlaZf9uqt4mmKZxwMNqq1UYxYndDEd9P+b2TvMbJFoFlMi6jRLAJSb2g
mXIvfTN61fb3lH0MowT+1tfNjSYvoUoeg0tpUCvoB8gBZ6w1dmbO1MZkbtz/Kuao
2Jr6B1kHXaNh0C7hS7EyFcuS9Z1W39p6SqtGbj5cxSMGhp4vc5zMoDF4KoNEYdFu
W7aCPVCOQbBHrv6SwtuvZozVXoDqR/H69mVYkz6mYixlKyziqD+An75FPJ/02oMf
XSNSie4hGVAklLQadVVlTb4sVKCGiEBqtBgA62hX7N3562OXJtbOQJun9TL7Y+qz
y4aDWN0gnKbpIl/UJd1Ecg3We5vNk/qvQcCKsSh2VUvOfEPacU2bolJu7AU88f29
el4KWLHJ6gIQwkVzQxyDLdhffosVEKAgnrMYyXqmj49mG/xw/AG32scroBOIGNUN
/sl+8KnYFajMzd8pzztNPvL/HCVB1R3jh70vf7G8G16/zHhRLPcvcul3ajqAplf0
fqIZb3ubVVvqq1lQVTiIYtQUkRSyhEWx/iQ28UEI/gHxeMH6rFFFzrXe4O6xG/8a
CoJFx1c+I0EH0Zty1WQjXTXjZrQ6mtxDMCNcI3Hge0EjKdieZ8ejVEpOOl9qE3oU
tXVikSP5mJC4cwHi2NWN0CrOnS8DvTlwYuP+M76ybulwPoyMiHSaWDB+oOmco4Fm
KqtgROQRVMCuStFv9mGFp2NZx4oJqDrOWU3Sp21Cv7izhIxG6Cvn4dm7kmxq+ZZ7
j/hBJuVXPyz2RMoNoHlmOB5/9ARytAOEkn8dghuZ8HzWyQJUV5zf9saxy8TsYcRL
+GuDPWIIeZLP35yq3O/adf+/7OW9b1NjAD0X+kOAEXbwW8GtjixYBP4YJUe/0aNl
rQa8I/6K+dPyYyZJQmkZnMRqilzNKMbrkQATw/h9MrepdsCZmv9E8J7PyN7Ekb1F
AnpMnF1SO6wTIVaCEvXwrdJQVRKjcOO4leP5jNU9Alpy3KIaR4Iz2w/I7wo+U1Ga
sfjPf+HvCi2zvuJSwNjTQqtf6pMnsX0WjbWkS/DISbdZ+W5EllRebxtE3KHZTTTZ
X+Ewayi0dEimaM1310/PfyDmbgiGD7diB7qSeZGfZFfV7USiQA2R4Sk3zW0ujTyI
a+jDVPi+ohACfNqdI5m94cDc9uZAno8jEbE36t/XP7Tj5SSODO/bkssdyLBgOYcC
mIKSGm6OoJSZTyhlw0FEq6bPIk1bn6zF1Gh7CDdtgjN2/F2f0mdmdsVncdb93P+e
708Yaj5EFqOcIPmeMJR2d6t/luNr4afk7DWBIlCm0LpQbSxqgQlYzsmzbiVhRJ2r
pILy9fV6ltFKC54+Chb2TMe/5S2YgNh7rXOtpJS/sino4EaeTSbNWMADaYXpFZBV
5VdDeKWI0dbviFedsv1lRNR76KjE9DowTk+hJayHkIdan+Zt2FTyDrvRGcJNn1pu
bRTPgbpllNbN10Cn7yjtVpPKxff8xcLb/jPXZXnSKZ5sny9YehS/t7GDEoZ41iZD
LGEvQtWvJFSbQtHsmegAT5P9hyN2G1qut0AoPwu2J9ZbKSkR7q3E694N27f2lN/k
55ZR5mMd9tCATtTZTvNLom/HyAHRAx7cBrz+JYF2GVXQFDs7cnTDXMKGEEMRZvQu
gS86f/+9zZn1KvkOPZxVmUtosc4rjgI8LTC3Yiig8PrCvlx76oQ3mgLvVlVVbsF+
jGq6bQMZf/0NPG/odUVndIB2RaOG/MT7UxzfZDG2avXHM0CcV/tAcyRQBpP6Yg7a
OEfcmKuk5v7xu1463e/mrwb+yXUaIci8c7ZXDrpXPCE27l67PTzNyv0EMxl+25PW
eu7AxZkOVvoZSNxyrsfsLBIc9XW29zuo9F2urCQLnnqI5RROfqQm8Ar+qd3pf719
P7h9Y2ahlksQYdcQiZe0358AVk92dZ2dHkGfIDU1Aw8k7hFC89DUjIYmNM24Yod1
QHmVL6I8U+Mu80N2LR6yceGpCLE/K5DesEncgAoMvDMqvlTgNgGI65ACNUWGMPzs
qRHug9tazWg/McA+TwM0jJrxgVRHTVLm+89wuk1rA8Ft+yJ2VvzA4nW7F/sNPBfp
1gIpWOtcEUVCEL7MFQESj/DaDullL00xyN3d2Ix/A71/A2K/FmF636xxqhwaZgZU
TIV/iNaa7HOe0LnolYBBbAbOXvTwFMNks0/5DxGMKxbw+wDuLBmCET6OuU/ilnvA
TBasjzNnXOWqwsG3CnHu6sSqgIPf6xwgWbhPngNFgPyD2wpxmWiIK4gS7ekm228B
vccLPkVdTqHxlklC+qvMBB7QDrs3xLMOGbt/zjhCszDO7G7dr6ZHGv9jR7LGGYoy
uc/K+DJFagbtFvy/7LRpktzw/LetJgZetOyz1lvs/82hWUToKi4r0GJ0roYXVz2y
YwW1Ax4LRprOoXY57vvawuE0ftAF7tpFDYV7QLToRsGb0zyFAUGTA6If3Y9umTo3
OX4vMGdadOAjtlYtYoqAfdatkJXqEWZRToi1W/3JiVgH7+5NglRFGrh704ilPCAL
FOxPdurP5OX5GV5OAoVjNMM9K7yX/JdsMTZdMJJngepzbaBt4Ci/8zrzk2lIEyth
VV4TOOM385KjuUclL0zRbcxKgrb5bDs2c5DuYBTnNhCjcbqtpGZqadE+9WNDR7Kd
F+z7rop9PrzTBMtzRVt85HuKeMqmHjBqmWzn1tl4e8LDrewNQGkBRSViBf2aoKrM
eQUo4qpkf/4KeniSCx1rWv0UUi5umCYWxcCpxY67cJnhnRDWhcQrWEm+WdWKfHHE
94xZB8w0NJUwVSkJrpG4LGSKGzX3qQhatV7xwJmpKfdU6D5phvIG+qFSEqkWqxLJ
OMARgahllFS4IQfmkArTwg4HmAZ5iWtvUKISPCaeuFHQdqdGH161gi65uhAZhZyV
cZdoh6tPBVhmbIhhf+odTUViJ90+gLHsQjWH+HP0ltnHioLQG3nPekbtAw6O4OwO
RY8rfiuI963AYcIwYh5o/ye44JJGB9rXUHqtV7OFyIRyuB7RPaKSGU+yjK/v20tl
Pwh8RPXKzE3n9JJal2PhmCrN7XcWcTGHaOdK6ogLaW4aOt2PG6CWxx9KdE0VzexW
yCpQrmCpAD1g1FTOS4cLr4bnOgkWNWcmi/z1jHYYyIkOe9s982JBIRN1cBH4qxmj
yaeSY+leakqycqzJtBlEeh4gYnpq52sGr46VTcZQNPzVUH7CABMzG4ApBmEpY5vs
YCJ6LSnk7fdvpD219KqtAV7O/BT6CFx2N3kvRP0zaW7pmjCQ9zXV/MmPgwXM2RED
X0kCwgZWSQw5JlJcp7qRE87hm/TdjLUiYZM+3URtFbiR2hXF40SgodK80SfLWuPZ
Gh0MCEJga6xCP+7i/PdbUKFRozswrrmm92xBFs2ndpqU2cN1u3uSOfInLqVRYRA3
RblR94ja4zYYrCfoZwst31rmZjhemCuGeSSMnritoIwgOXyr0mERJ6qFSP15S8sy
TdLvZfJjqLSVcQKlT39XXjuSz4Zu72KIqqUOlet5byD11AOhsBaBuaKxhzefK/EN
iBD711KK8rb1ICDQ0cEJHimPppPBRXNkY8oIzcQ7JRqdpCXanyXZt3cmQBtCcVMA
gKXM5k7xj1q49I6FscEfz/lu2h7lhysH6a7sitcZ3rsOeSpbWZ8K1TaaUk0vWzZ7
REnLxnYK5WGuIvmBkOSd35kIxzKuISpxz2C35kRKG88=
`pragma protect end_protected
