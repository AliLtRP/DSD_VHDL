// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NwYMhnW0LHItiM3jkoXPpZrNXGe8qmSBelcQTC2RNWfjTBHlV6BpDysFZZOVObCL
Y+eO7+o/nF/drMntY/qwnbgzIaxQK98cRq6rlYnM34ddgDqc4M0mGjNL8Bvnp6AS
GnMDTLgmr8ybkXhCiA0BWU6LFVnbvF55iJLycJESdRc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8336)
/Ixfl5Jcwrgp8b8A1+CZC3MQx/N0VVqp3oCoT3JfRPdXyLUaOPpWqmx8h6hf7qf9
jRGM57T5E3ZvwPhitkX2aDzS9478h8wdU7iedcNBicSRl5gYF/FtiTr3gzTCtYYT
VtCmSJGSDvrH3Y1T51GS1caigqMwnWW9bLai9fk2jYmpv3wGgMu53V++QCJnDFkF
b96Hv7sJ/MoDktSn9AvZZtQ+EU+jMz8DW1b1ImFr1Q2RF8KyxfOTmhj7phawbWm4
57zbETXTOC4UAb4W+5E09OHL5b90DHJkhiJHmqnIlD92v7LlUaVvVo9hLivH/ljY
RQmGxe8/baeoxcQqMNYHWGwdYLiNPbhwAWjHDqpAECJzAELe18rUeY6yn1HqQWqD
/+k8eX4Up5FcThyxvT7UjSJ8UGdmDFbCgarvC9Wo4WUt07G2EgZLMAhTHNq35YjC
cyZ9zvAODu7MPHG8bM4bFTN6/KMJ0Hx40k5Aji87Kdk+Onf/Pxm3uJ2MxXWzJmBg
RTFUSIdq1zzDaVTfKqOIA9ikjoqjG7qfDcYLBm0YISNtZIiYA2hNpEgsr5fFai0h
9LJldQ7QUP5JtBB5BjuNj/kLyd9979tBtMp050TvB0JoTF9pa3LADT9WoP02imVO
ttaRGIuSmhKY62zQLiY2Tk7UiUT7rCISal0TAlPjJLlCABq5jCbdoHlg3qZnQW9E
B7FNRUb7oEXo8QOa2pl4jAKHJfdRl2buVcMtDHZH0+xqPJ36J3gAR/BAm4XIJDFy
m34ViDkNyCrYdf1qciJpeQevtkn+0NuLL0/KNj9bnzNlqA6OirtMXyBM3lI4xYWJ
qzyshBoA13w8KsiSo/SwVMiHf1U05YqWNvRoo061s22mzsloawTAtcMaO2fEcmJl
kmkz1BUKqr2nAbBhTI8rAiy3cZrv5YpPW1koy85suFm38eAnWCjDWgRwBS2o/bno
G10L4V13dGjHKdwUx82nOo9xrALkUtVNtDxxi2oB2l8ZuLMfHet1tqYBSyuOUr/y
GWpOhTtWbGGwqYahqnQQi4A5paP2hwH6y9HbXNhCLq6k+AbtMRfydPYTWpLSStFF
E8SlUORLVHn0C39DJvEKK2rLI4qiyg+3yDxvvRpprewkWTiuSC5wWE0vjDQFBpqV
eOYv1bEt8x21QwuXaN+PqSLVCx19ahK/dRHtp8DVr2OERoiajWbtXWlBKDByopmz
8nt+PJyMfN9k3utIdtGz3M2tL2EDtf+DzTehhjS8j/OtAv+6OQUaDWXte+yOMDxN
dJ4u5c5j9Z9dKQPULYZxtyYn1/RgSPcSQPvyIkQnThsBXhVRVbi2aG/ZhWzpyXy4
xuFiVTBLgdBrFSlWBgMxdpl2D4I5VzNOUZxe7rfsF30Rg03j/TUCTRYdkLJHx4kh
vk6IwT2/mhrZm2isjKb2E4+PCs5/NfeQkV2ORuC/UFWNw9Ip9K3M5PCnOS5Sf6mV
Q91YzG2VGmhsIzJKyrZTvSv++8cTI5YTu9JELDCoX0NBJzvyhaK1P9QmMfWUPRLs
IOw0bKo2NU+nymLsETxbAuCZ1QKwh+6Zd7PIu/bI2kUBr19sSmUt43sfdqcNahfu
xxNzEWLndQKQ8WmzWv11ZJnMMp/r53ST3qTrFOA1CgGPxKNvJlTZCxJV75kfsYa7
RTe5REFWNQgZ43fjwmbnzqef0LQ+/qvRG5XXOG5ySbSHfxd6TXoGNwDhq4HMwtEc
In8aI2vGa1Ak89qwDCnbpZadezG6UV8kyURXAwR2Hf6MJAuDZSefW0lJX+R4sAkg
pYJED7DSJ+zrueLZe8ZpjKYsnNY5zmwmPoyeG3RPOA82aEtooq9ijK61B45nPKMC
23x7eglHA6a9hTvPyvScy1+WY0xC73l4yyG+fC3q97J+i/kBq0Vqb53scsJW8utl
bL/LcpTJlOR9f5EGaEt4Z9aHKNNYBvEtuSZjNdmafKnFFY4ULhXfBmO/IYQ16iKm
FoBOkZhKrEiYp4iiaAN8HlK2CFZIiYEgIPwFFF4otoRxuoR7n7aK4eOr6iTCCRWc
Y5wsDUboin9bvVeQLyPat05ZqsPctB8D7h9I/qAz0jGuLEOrjOkviKLs5WgK8HE7
lW1clFWg6J5e0RR2kbBTEuxiPsSeahCEdqYDPG6AG4Xpd6+W8VOaaaBSQSQ60Ol5
HVz3/x33lQ/Ox7XOBaTAZrw9LRo/cjOjbLAAqKBkd7hl9LIri+NvQiO8aLQQiKtT
MuKERym2hJHvkvpn7y6vRUfaJz0t9j3wyn3FIG65A62Fww6gQExJ7Kuhhqw+lunP
8GIMyCNiOsULBEcJrDU6mK772MaUi0IpImAUAsd/Avrg8ejE4nNTCkpYp8cTafXk
673kaSwgbn2hHK0KlMUTsFLQSIEgCcHLEMPVGJaXfDlBs9P+eMiAM/e9rmoC6f5d
ss8F8ylGuoShi7NdM9IASppSW5FOiYDAOLYhdynZCLm4yVW4UKF1StAwgwVLgPLP
2JkIB6BBg6+MWu72z0u4/KY8A0H3SxA6ci6pOgLa6XGVdfr3YeraK25/b30lNzls
9NQbq48G3atLkvAQjRJl71O/L68a8FvPKz3xfhzc3Hm5D2PS1zn7v/nUYvS7+olf
calKVFzAQyZd1fwjmqCghtVWeHvvHwVmu9uxS/LhqzogUExXTe/xFQm4yl4K6n2U
IsjNwD/zIPxOeQwb7D3eJi76mxGcdoVohvapaUifB+GE/T9iI4c/R5iE4K+bTGrU
uMXrOZY7ghsObF4f2H3wJjUw9mmCj0OzpOvmwqhI8uVKIxXYZAXRVmq2YV+I4sb+
zWPRVhKfoquQStrhHWhiWN+mLPfbB6A6fNMj+7ZWJStx47LOjB5qJQ9l1bFWdbi6
PQLF8UtLAgeL/xtVUgSko5+Y0v0sDkWB0Xmjn4/51BYJRgaVr4J2KhBKpa4MveXP
PCEo88cmaEQ72YZz0amyAvVK8L5bMhOIHUgTlkeEO7peGXX91HT4uRaCQ6W5jhiz
8zaiB7b++9pDxaCxRee65Yw93dnVK6iy+vcxHnsaRJXdFmxUkvGe4woFzm7S3B38
odj9IywgfuyfkjNG3FCnquKY+JP02LY+KH/LJy2bzC6AsMpz4hVmEN5Hckcwg5HG
ruFewQDDPa8wB3ez7hx+x5Q5RniT1iEwMDV509jVUrZm/q4KFsED0kVWTKwpNif3
ymdDjJFjOIbeAmCh0iJl1SFK3zo5XyZJh6I1/lzi+nuPNZjjyMZrDQ8oOEYOsTv4
mBl/j8CRWkYHnEUBQjMKzpjsnCt/hKOJf/WNYzLDslHOM8TPut4bBFysBq50z3yy
mRVYCc5rBtkn5XD+MZxK/fHIW7/BubGWMH+Y6Kf1gYmZtFLGSrDiM9EYBSn8kYnV
zRIIeF7iaZys832HaY17BybSVyWo0rs3oTeGoGqxUbzK67G2aBNpvfTu2t5YgtvK
MmLYo7EXjtpkhOIvFPNoJbg+YoWmEM2K0Ypy4mEyNlHZUD7A18PX8xJ3zbbp4NX0
EGWN/OuUCiGnwg/Fu3W+mNzojHFu51iO8phwXBG4HbLcb9zgtXzUVOvb6qQ3jFgy
Rfyst083oBDepVqrS88RjIRZUsRuwYpzxPHefAJGduqhGEHWIq41e2Cz2JtWHLik
AFjSLyKIt3VZQxRGqH2N67AeOpSefCU3SjrGi4Ub9TsLfp5z2CvhPAee7cCgzwmY
u3TSQ6AoPAcf5BOx5qNcv15n7MclVl9B4ZrzDrCsfs5ix7RvzOY57MYEdQUu+Pq1
kDv/ThbANO2FDDKhu+RE+SCyJfNdZyl0cRmYB18icxdXCLeiWiWk+BdkmPUmAtn5
e///9ZLzqDdtqCGqcsF6D0rr+Z52rOkopJjLxDO0BhVC1DUt3HunwXwqDr6Y7pDL
Lrw7oofu2WctpOnUJGbkvZFGlRGBH1sO+9uPphwOGzdQzwCYOlC7aXC++pzPjDH7
S/L+Buq+zzC5TKxbkxZ9KcMCg+fZDPPe00FOUQeKC6559Sj9Aj12IpASRqupA24v
zEkk9LXiqc15QBYdF8Ly/mjdDNQCj3qRQ3iThT/ndjSDOCqCJHhS6MS7LoOG5UqQ
FIGXLbCH2eY47FZjS6FF8BnrVD2zWDKHAwqboHfXEgfsst40fdXaq+L51ENgMM7Z
pquGnhUoYFZl5vk3CFnWbNov1Uo4hwf/at29hZWV6IByQNhmDA6UZ2NWG7pUfhdf
2W/ZXSgXJCk9j4XxH3yIMdN3nLBsELTESIr03QvDdqMK+Xn78vsajcJU83Zv9AiS
jer5NfVOa8zXo9txo16/VQJQlSmijz+1UgeA6q/ULjnLuPXlHe0dPb4CNPcQvTGQ
INe11Wyhny4f4eA3ArN8zeMfvxLIPGVCgDc2zte83BVRuVgmnG+JKu+AtY7j+dCU
91K07FwqjsVKJcmd0T5uak8ZEAtmFb4ccfVQ/cArsrfwHhb+IXNY1/OjqrpOt7zk
5PC8N7YKyCA/jgBKE8UuGltqCPwNSQ3s8whb/DbXISUknwy4EgaPCNpIEIMqmVju
d+Ybkszep+t33ZQhxjESI20wjzz4ftWaCpy4GV+m6Tvwk5XJKGJ5XD7QMKfMwOzR
NjMCHkFiIkeVR31pbmPJLoZMhuuR/o3YRpEnfIp1eytcIz0Y7IvZ5zQOkm7k37o+
vT/kFk6otKhZCUQ4tbLvONIl7HAtyof8yKwHI1kLRXoirxRw+CZ58Oyvi7Fdk34Z
uj+fiaVqwmJu3nem3rt6j/u3keN+NVMBJTuL44+NnbbSp0H6u6ZA/PGKim60VN2f
RSnW3eC1X01PjRo6dDPo9xXV6cMVb3kmPrzlckV39rsIOUWw9fg3iJ1Tffq6EKms
Ht9bzWqwkCkJc6X8MWYTzy/WE7rp7uYKfoLuAFQ5h72cO9V4bIgIMkVp+DDo+ZQI
crooRz+CIWX4Vm3OOJKzIioHEBCWpyWAadhWGR6CQKHCdl1A1Z6QIix750hSopKJ
HwreDbrdBriniyXb2l1WxiiTVPQfQdKFS1NBsTHxsz2w1CshiTNJJf5qFauvxeK3
7vOvEd9iM9fLgaIxJ0bSuBJIIhj6s6jgDXXCCIYRsoI5XiFqR/aQmbPWo6MIJvyL
FFTcq9yqGj85avFTrBCFTtopdAvE7OP3dENWZbpilizYbA9MSyALp/oX/m0RdECd
ftHyqNZnV43QluiiG2/iPaqF0TzLvhZVN5Sn/+FOsxmJlV3it21X8eNjsNt8Q7eZ
UVNw8z2u0nqNBSSat7vZ5V1Kg2WceYhcj8ZCMUNi9f0gKG5ZVfqEHYucmwlkpfjC
nJY36hPcUYXBEa0aBBeqx9xodABqCACP1qEiZqc1OaSLRDfYO6FJikdkhLXTUbD/
Xu4qQc4woLymspjbXXXlmHFSn4vTMd7LB2kf+D3LJuuaj7Hbw4/YqDT6AgzwxhJS
oWlWPPasy2+scOwyoMWbFCjLUrNnDvN53aiyDJYt2UoNZhaWc6dm4m0aIwX93Lj3
/6M8Ocpb9tRM5MXYFJB6KStINz8F58yxep81miGFkAGv8kS6FiGKif+hLPpN0Ia2
CecAHXodsa0Cqth4b1QHZMUbHD//NJVJpDpTjzv/4fxSmf5LIXx11TK43lmlW5NC
ePtj63neIXx2+RPZIQzsldYDHBsC/YZj3wcjZvsZCBwDT5s0oa4kUSsqqQMfC8MF
NMDLWzigyPIrlekO/+FUkme+AtrYLLH9I622T3LNPEPLipIW0Dxx1OegoaF81PLj
hMNcMzxbKLZrViIO1cpYA44EkZJU7rcjPNVRsNMGace3iySXsJkFlgQ0EIpw8ZCT
f6EFRFxqXJZUjGDFfbT0KMD6AzhuYr7SDvrB34wLOHPHXPOFlfJSeHb4olSYIoGU
+9MKpeD4xwDm/cg8km6abLPQgv5g58MlBrrJ3TryZwIx2O+sTmRD6LVVRKPWlR7I
EeyeXEB6S0X4Kk8YNlEuyfyoY9sfIpGkXsc42ouSjoJMl9aZWbGjJmLNoU5QIAdP
KfrLA6ZvODFy3OqLcp6kXHEorbXKEF6xMG9/44faOI4KS/cRZ8zS5wLXgmH5W3tP
/v2qJoPCKXY1AetYYrj7Bg/ww+rh5voTy2zA8bW+drvJTmoNAfnq7SYfYowu0/vI
YDnz15ZBMPBymAmJ6etq+dIHd7NDpgZ6lVEnWlExjTXLedHoNT0erZgSdkbkBxnH
EXCXFHSGTCP67d+jujsbRkuse05Ky6SWd2HY7i54yChCjNbG4t+IPEboRYpoYwkH
dWxhzqzgTEyVzMCcv23yVXYi2cKJJz7hcz32O5fPYWu1RJihiodl4NVEn0Ew22ci
TVYT75jTnmZoUsBemkZ879QVDAWC5AcUc5jSy3Z+9J12RfVKqa3RqP5FxQzqD48I
h3SQzlcStFm94IEz496hyudfqJ+/3H8S3U7RA7YFpWN1Iw95eb0CskDHNb34D/lE
KAS0X3MVz5Gs725BwFR0CZH9uGkQIA36I4vn3BEchhLKOQk1j8/5jRj59NOPvwSs
Mz4I+BoDteMtEoL5bNRpAJVhzZJJrqYhNip/Dld0pukl9tZerF72jRn8KlzCABOF
/Gr9eVscaF+cX56gJhqCjsa69v7R13AIZbs0A1u87AwcmbE2OtgFmU7TAegpkrKh
SlaxKWsns6IPNxsfIPFjexT4apJSnjn3Rypn8PBc6cANyVU8IOtWt2FXpNq1TDJP
ojTwftrsvnIE1gdiu4BCl3Q9N99Rcc5WKwhFyoxjy5Ja8SUDpFa54S91rCd0IAMz
RQtmUQPYzRKHbgZ2WjJWDl1qk/kRW03ZL5kqbyOJY++F+lRFWgfXzQpIWxU7Kdur
TZI6Sy7cwwCVOjEEKPMERY+7lO5QWAI0Di07kRPUCmip72liaVkeaBYzOCccmdpa
UfcR2DE7NzV7hIfJkZ05XQrQ8V5CiDOG1DG6zCcO6ml5QlB54y2dFx096Jb2nJ/y
hHtvop+fAfSeo3HN62YOzxSHixntxv0Qlt5O9l4gqXsVwFr+M9zOtcPNZYUIMaKB
YT59QSxdSf3bKUKJ8O47m5qKrUDII1MaWf/TcX/hVJ4ksU8ZUDiNJjOq07J08Lsx
CfKc2nnMAkjHVU0MVF7bW5w2nzYx9Ws1Lt2jIL3v2496EEHtpPPMbPQVnrgOuUF0
vCLl6mrpeAwDlRl/lm6yv0NRVv44luhJknM0CRXlVvay4N4bIdOGAGrRDv7fcRQa
keGYyFCOk/5BkRfbNvJPfd8to1kyjUOlx31izWXxPbhctX0x7MDV5/c6MXujNfV1
L0BZBhNwHMM14yaUj8sUcl6Hbyr5/lZNjG9TXfCgXxHejdvRL3B5IGXT80AXXnky
u4CehgVBewZc/tRH3WYzcmD/8tuM0uylownwQL4klfL1kEVuR3s4Lr5NmETj43u4
bkyniI24asFZF+ehKW0BURb7HQGuTsNF7h2HwnSn9h3MpuJwi5U1ydOH4Io8AWYo
SUC6oXzXMwMP2cobg+5UH3OQs40UKoOpX0dSSxePRABnUuvu7ezStYhoCSGhuxUf
551fzhKHf6UPrYX6+34kg3++oYi+eElw4eX+ZzhpVPlJDEVwg2XN2ifyHDaMfFIY
y288IYE5ifhr7XejZPi3QoUj3L/qpZHtOpl8lhKsJ95QOKxfq4MNqpJA0N1MkGvt
OP2i/+dzs2pa46dF3Bkb9YkYSBIe4WpOcAihPbomSphToTfzHBKFUuKDc+V/E3bJ
i+z2v2GSVyDgJ/1dcE2QEaYw6Zzk29gdSEeAqeigJ04h1O6w7nqLHRVTQZBr5bkx
fR+QFhTNPZafSGbbSvQ9DcN137nE9FCftbIBrrIHenz5YJ1kMk4uXuxUN7UueoJp
0XFiw4tfiag02TKOOh7CAI/J2VetYIlq4GD+DVZ2tWRuUw3B2xacBWhyK7Ukvzdb
E/0bQAeTF7WzMpExPUpSu1YlZtoDO+87cjZPAQ6Y40csBT0IqAbKpde6zqkdGtme
35pUjeiM24pFOgg0mAy6uBeIzPFPbLyJ0/fL1SG9ynzOmELfVznqFeoYGYcqQDt4
7kl8wUzbWc89MiJ9CAjv3zQXaoxxIkRId56PvZEjGQ93R1N1pKATjwqJDgGXF/Rf
o5EGo05z7qzs1aVRnwYW6JZUGXzmND8bjh9YVkMiyG/S3HQ25G7MJ4friReLsFc1
5N+DMMPq/xCndLWkKqgh0yoMBWBIyYbDQ4hEP5V+9NTpt+mPgxeeTSxt63aG9BH0
kpi0Ozqk39o6oNOhbGqvVx9AzcI23CaABpna4ptrXLkVMV3ZJDrS6DIHTqNV7vL/
fQ3SGc20q6EsEN/ZcAuT6u8Phd+Cac6TiG/5FaG8pmRaHPf1+vvpVyjOWIFx1whp
Gg64ekF1Vg7Wuk8c5mkz4rWSfcJFSLv82I6yYFriILIJu8xIsQqzPjWRyoKCfxDe
MKXXnylkah1EBj7zsNDrYF9FJkDuDMrWDr4jMaI8zjiCRVYIsTt5LFHK+aB5i73c
+fW8OH7vIJcN4AomlbvwELnV4iyjlZKqVlaLP0qE2szhZG/dn1hhwspmbo9H1dpl
xbdSvl+AtzHjTjcMePQBTFU96V9dYziCtW53pkvRDeQgltP0KiDRH4G2sWlABMVr
ltEkySiAKM+zLWkS5jgJuJJZNO6biFP0tyYxkKoiEUbF/WLwNpe0bp6YF62Lxyve
bgWA0tc20QRNV95D/HlJsqRUiAyCCs473zhOI//lSfaUKHRBLVr2bNV2iLPQMLvN
QkHx0ZUR390TMuFXUpXWLhNMA0iG0Nv49Pa9ueVqNtmUpuTxYRafFPmhdeJoR0Z7
xGi9oI/xOpCCqJJrjR3GPlj9QUCovy8HJwhLkU4n08w8PxmgrC929cbvMpuLOcdv
Napo/8Hs1q5asIm9UL+HCH3zuIveAAUMjT8jhTCB7gC69sP0J6bzlfNdUp3PSmWV
u5BWBBpo4x+ymtYCIca05wm7iy7dCqkM+2Yw3ouPErMBlvIkVJLIHDjsV9Bybj0L
bFRy6gE44vFzk5OW00vnfpmGnNP6RsYSZMXmhT1ItkNcWrCCMP2c3wWIvcmNKpU2
Wo6CJXGhQlFSV4lAwYg69XQSLoIGn3UhEdhkObv6e/RHAOIUmjPKdGbPXDUpjnTd
XU8DAc/LUyPYxCD5pCjJMipERCRLYxvuNmVHjXmdrCKeFRu73hoRtUtCvOo9LGJW
ui66tt7RqmAPr+e+v9eWUy7jjj9A9RORldrlC8R6fc38leDntAtmoyCNn3Rlc1nj
Q8+4s68SvgDKGf3mihXmsND70cfMl3zy//+7ZFQo4WUY/sBo5MHLfX5Xsr/rCrRw
jJXK62/L9PLGZiCt5jEyNmMwqKuXnU2Z7hBqIu4aGLTEUvBRKkA/IMndcLDb1uiy
RjQTUx8DIr2XtyDxeMksiBvAAyHQQ0imKtHL29bBRRKIlRNAwe3JPy9HkNblT8c7
0fGiBrcoKs+dmNTOSkdeEdrdskGdpMKwvFK8qObG2flbOy4zZGHWLNMaBdLwILk8
hD0P5EDQ8ddM/i4pKZLnek/iAxVd5pzFvpJsqCbtpSuv4tUZfsp7AFpVwcnsz1w0
jfQy8gZ/AjzHL2o1WBC7F7RO94wU9UfQDB3X0XgyGBfsMJLplxJ1VCPeWL3inU6K
56CG4LT8NaGLFdxl5gozC5Q/uQsDbk3cvpiPQuO2SO0iplk2hCDwn2g0s4Mg6bwq
tr0ssRqpYRd5A4YD4l/rm+udR/otNP7kCmS9anjsFtX/z7d9IT4PFYkeCL9Iel86
ncVa4egZAFFzH9oMZtznXumcChEBBM1Akbl0uXEGh8kZ2Ak+kRL2gu+Ly9YaU/8g
KFEaESxiExdfX3sXA8zUmooXvnvTTPvS1w/YpP6cwPz+nCHWR2e/02GFs7LktavQ
bdm/BVe7qDTM/QTYFQrSGaHMDpX27kavh+HowE3Cg2/9po9VdlnNLqWhcmjFE6lc
ihx71/OD1juJeXHh1mZRvpKBOyZ582pSgtyjKoqKXNbJaekGTeKX2UqsLwFo2oYo
koCj/yej1BfP8ERSHZlPegcbECjhR7bRrJYzyKbS2PLOgtGBzUVBU23qlHK2vU6n
vLxuXU2ABm7dy0sbYqYv8yB3PCSAr56E1sUCkC/F1A5oEtHchCnBfDwrG+9NcEk0
lkLTJ/B0j1XGrnKM7tr5nNWECNezoPuC/qHAQQW7aOmf/7BysphBi8x8EbzL6cRc
IAR/VarUwtSR2neB42XiqRGLmC0yxt/MPNw5+7xOeNOw78h446E2/0Rjlv6Yr+cE
68NZlyvnR6nwn4d65KulEpS6AV8YT7mWjry+dEyq703rM3RCfB+Q/jtOzNtlzBBj
fDqn897oeuQGILNYQJN5wGAzbfgfXnY9bbvGfW2QZacTPc9uer2mZ60zVdLoEBf9
abLYUua/W3N24w5tGNblzAT3Y7xObJu05Itb1cuWZwWbLrWoBjxW4AofIQS+sUaW
ClNpxTrwx4ongAd6kygF/olGsePR7d2OngZk1FOHIZqWpoBQQI1ydCO45t/VQ0R+
4kqcA9e2ftN5zyLBqb5rGKSfRWU4ABWbqUMCXRwjaWFXVGZaSVjec2efdtxXYNYB
wM6QrCRZsMe1z0vQqCD5I/k2+A0k3kFv9miMmuoHenCrBsoea5S11OMel+mtZs9W
2VHmrWZYsO3E/be0stJjRUwphmxibecRYSCtU7kJ97TS3gbZuSLsdWLYcOj4txA0
pHiV+1kZgQctT6z98yBOWLzZ3V5+QRUTc1Wl3RBHazdRGId5Whw/u7YbPKQ/4UnY
V2Wcdnav6oz89Wbmz9TDVasTWihnedkwh49kFHyYexPB1rVPi43LWKqmnf5cjR94
jjj4+jGtgkdarK9NJfzfmN9jO/8q9ZdDjfMLir9dnSCHbdSrp3doxkanZKZIcdRJ
8gT27y1dtWi4dFF3ugNLwgGTH5gHkh7Jh4K0bJ568P8hq6v23mWO+2Wu0r4+m45v
gbxA+WatM82DPhnBI6Dn3vDpB9PJpHEWj79j7+Zx1BLJiveSbViHdW+Ei6AsSn0M
zcXnwChxRSvn/u3rSmNsYbZmNpF7foyK/SlpDT9RPPI=
`pragma protect end_protected
