// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
E3HZigjPK/UD3kAo1Zf+Ly72/k6H9YIJeMGGclttWjuUMzZDHpsBS7/0byNVY+9r
WmtbypciJA10VAm7xFh06YpvW8WbNIfwa0Fs7KC5pgvL113Ly49wbLkrSgVj4B8u
nAOu5s1OA3epDr/Bgc6SWP6anvcYcOQ2OjSNEDkF/UM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4816)
fvvdLxfRm0TClDBo9y6gs2Uc/qznuh+EvEK4K0DtUeFadZK2yLebpKR8bdnnBsSu
M8s9xOB7youQ469ZqOAIeEm9HUsOi7mlr2YeYNK40NneqUElpjdoBmI80FxWA2Kk
HRgDSOklHM1sseblSgr6i3Al8FZrEgaTagbpZ0PAWczRDfvGOMzzMuNi108Pv8qt
EKCSeQZ7jg/SVOP9qtupMKZjHCYZXgGa8lg92tblxjAsQLoIXQLIoCHPzI6qRtyv
af8q3JDacVsUNfHvQoiyr9UNJLnh0CFmKgQIxQXkK79EUavOmjs4OA2hCwXhUfAt
Z8IwohmXtJTUZsJTRhtZXpaJTVfBWD5Y5aBCI6qXcUu8kwLwukpwVWGeg+1Rqd97
RDWS9wN6Fj/A0OvgtZsQvMiSIw/SU376NZCEpBF2rBfF/bIKHVaTsRj859CHxi4u
2r0BMIKR7sJmKnq872x9OrR+Uf7oP4Wl/5uhBaV3zC5XnbLerCxrCLgho2C2WaHG
S5ua1X7Sctr+zCl2rBE+DD9Fbbamwt6k24ITmTGjLDfqKL3yzjnwvHobTGRKwKQy
6608pE3cw1M1QrhurbZ1Jfm/vsYVV7mkBkhaUm3xAal6aAcXe0AthcrwyofMdwn7
HlkxzSPjlZeC356LeDDNvDd2SY+3h9JADAmhrxMkYXqwphhINOMgs2+E6o3M/eF4
C6JfdHHw3ZXIRyC2enndg51XRUEVYTGGTgAKMQxMIjjpPjbAliNZONcGMWbEPC+w
z9fa4ZqLrK+8mMvaRj2PAB4G2FdI74HUJjOif3lq2sTxy5zI+zIdsiy8TrZyE+XA
/krd1py+5tTRLriahLqBmaS+3Ksxy9ddRzqfd9sHHfbC4XgqeBvI37u5EDCjIm1e
A5VxGA6yjYhSCK85b9wiBmGU0wOamGAhsXA0Wp4IqZTztFy4JYqRHqvI+FdcHRVb
3hF5PjgFDnIg1wqhlj2laX/zwTzuCffDYjgo4itY0MP+tx+DYwE74u/xr5lho6ow
DDxS9TDyUoZYZIVs7SclZ+cPN10SIjZKZzT37jJfrkMJSp0xoerTh+h6v4nyZkt4
7PG7LA3ry77wTwx+o706hRZo7DXCNP74i7mUJIdHxBn44bhPd0dHX04XE9r5Ph5b
GTMltMDNF1+J0vv51Dm3d68L+NBijLmPVlwdBlCN1U3ppFA63ZuRF1aovPXSBUnt
TOr9Fz5DS8RWbY2WU4wezIgl8V0WVFXn9XXeHNzB47rbS0Jl4vR3jRPhV1/sJoNQ
CR5Zxr6G7aSZGdFl/O6ci2Drc5fhwhUD/UM32aO2gWF0gs8Vec6H5bzk3tvDthCL
GcN7vuljXv6cge0z2I6/Bv6UmShvuEWKyjEEBKWRvakhJiEhEjvFb4ngkK4oPEcw
17xTEl6yPVRsW9hvowTpSpV40M0dPLPEvW4QeuPpVwX1XlsJyYCXDdXNxyDyl+IZ
D8E+sDYGlQqmEUUHjceLKaBCcbv3qiy4Gdqlx3Vx8bmjcx/l5YlqW6sXQr7mKoc3
ZOOQDPc5nwG86s5wVnyMtvS/rFwsZXPVzm9DbVEHEiZtr9lqgbpKP5F89CinUebs
QFUBSECwqABw+B4cCqBlFoQh9fDjo0hY9XzU3irpTWwezlVQV6tPQ34YjuYlibOu
cjlkZTZElpYgO/8gY7j0U3q8V5KEGJPXn1x8AMkhSkk2QYJwzGNiARD9cnLpGkYm
/vPPVOVw8fhPopt3BfWLBqo/IhKDd45hGTdz3CEhLNNrKmdgY9hAfbNG3rb6QJcO
RrKySYvqZgw8F38/nY2jL4vsaWIu69UU8iIXipTdXq9SsYOR6Y8xcj+edQIWv8Mt
FrGUAXZcUrCBWzpH35xrhwfhWg52Hq698IkOJYdkarGcUu9+vjiYBDOzAp4UA9qu
LX0Y7FhDLM5gWLI5fpeDAjHivTgfZFsTAoWZUezmnPu0ee+Ax2tzypCgqmgU0iqI
/zSyPifV9Pgldvd6we6D21INlxIaydsZUbb5cPXVSvYNv6uQX/zEWGdTSedoBUYr
u/h4q4FkCEmXoVzrIPmbimZVBzZSP9EYpAywUvA0LYMJ6cfEsj7HoKaVzOt8tuFj
C5X3rWnxQuaM9VDOegpZFsYUYjmaO7j02F9R+ODbWO9XdcOmbnw8TxUaNQ8ygJhN
T292l5+i/kbmz4Xu0KR1DHPqIAsDr2S17O+tX00maR7Q1f79GxO1eStJ2tPsimiS
94o8r/lr/H2UVjM3XRnsQK3k7bhfK0C6smGb6kHUDldUBVupE3t5eLlvSfEvHwMG
bga3qywEJMTiiRiVKMjA+1LIG61zLfabWIewG5msH6vBWDi9bce0+r8poMag5L6V
OQaItWpy0gBeqMVTfPdw483Z1QxJg71iHtQT0E0lvLIrKUsHSLW5dVikJOcL2wPg
AYjz2DBZ4MKNs/DJymmOiDuk2OgCvZRmxtVoxgEZqo+8wUDYC0yZxBB8RuoafGb8
uRwLyPmdEO/w218IfF6iV/z6ic8Vh3RNkA+pspLQuIao0sVuND1sOU1eeZFOG/9D
2gmfC/zS9WSO03pD8MaM9Si/O90L05U2rjmbhxXMHRXa4FI+hT+tanrfnC4bhBMV
S5N/Y1knVa7XfBONNYawt5zTorYhdH4XaHeH8I6jOQZ60jG3bd7ykpHsa1gaDBgD
XpnlhLA4yy4WXGQs74uHUjdq6dgAMWzByXx0nAtkrY3xEuJzU5jkg2PZQkWwOvmN
oTIjYZfxH6Uq2Zua1yeI5/A7LUukn4ZsQhBWIUODkIAvvqRtu0uyW+LDMO14lgi7
jPMJ0cJjrCFTNqmmQp+JGo3jytp5B06LGdyX6ZsIva3u9+VgWf+HNkXs3cjKtUB2
9kLCEav6uC3b6A4xmPaWc4H/S0kzwQlMyIvC8VYV/uUKrpugW4oAVk+XY4+OgB6C
2EZ9qguBvoDry7FcFRmZQHCbMupyF6mRgi9qt+PxEyHb9OqOJdYOfz5Cru9EAI6T
jE3KyaY875g6WUFGyaNIHVqxCg/l9LzjH6hspXZHW1lpCNjHvv4Uk0rtjDJcyFVA
FcF6VyfcSVbDZ2yMQgTPEWUlp8v1oQxb5fwNvV2j6zxBczPceOADddTYCxJfEvmC
f5O+U2RAO99RYyb/J23J4rHN1rALeJReZ4n6YM8Jfc3rH31c+5cSg0lyrwBHOgmJ
X8GbJ0iZEFwMt6ts3RGEXHd0NCwQXkop4tPyfjG+Y6HXh8/SXeR72mL2NOyuef3u
MzgNx0ptoGR+f4ySjV0pz8zo355dJ/RfPct4OTZeB8qpAzdyGFZNYWNFUP5OVJ4h
nw1nT7ecmaJIQ+HEOFab+9MfUPxo62fAOfU4jLuAxAdokuWkng1snB03YACTRKgz
nZ1HCvkomQDXUlw0m64HL1eJOtwJChp7ovfc4/OXCVwXzIE20/gnZxeAiex15UXA
aT5sG4jW3wfQT9Qwje/8m43GB0mO9wF9gs/BthRIc66G1kVB+J8kDKyjzhLxCM9c
a86a9ZuDxXTz69RdmWVTPSZSZuMkwzxuLlv/2LWjj2fXT+9OOsNB/lp6p4sAhS+7
6GAEh45GTUhiSHh8jAdOdwiUGjzhDRMFi2WUmN7yVXmQot1ZIwvBHE8KNCijlZnz
9G7c6g6kp65L3cF4LyphA6VUk4hRItCeudVbB5aP1+GXDa3xMvHfvQhsDza8Q+hS
R0C9oK7iqWw2ObhfwhxfluDiXF/1ceFXoICyfxc0CdOzcQ7XkIMp+dh1goeU0qkV
vUMV2lMACnC7+a4TcyDuvLakhiiMWk2f/nxRE+63yOVbPRHkTrr3gLSQlLDnAmqW
UUXd+4LVumntRDSIq6nPfvxJ5yDqQzLNCURCUtU9jnNdImU19CQuHJ9Z6Rs4rff6
WUNkSqehN3c83JBwQQJ+/JF1LDdevjFIE6hcAxe20R61KR0WN+wZu2+mDXhRJJzE
ZiezHJjs8R9U1cmtoknErEBA6UxNDmsApzW2FXJ2BEAjVAIkKV+7GAZbWbnpnvCg
6JeiphzOtPFRbuEMCwExsu597mN96gJP0Lp/gcFEO4jx3mCDeBr9+u822mdVqdyH
iT5MxParBb4GXNYoKuOcquwqpc/x2UudwL/Uw0hD0E4jqV1MCpTa55mmOYLVeZcN
M1HgsZzb+63oNwG5IP37VI9o9Hpm9ZI7hrbYRsdTdubpFSlM1VPx/rxca44GLpFG
FICpuUgZC8uxvv2Njx4hS2D0g1qnfcOnWt9hKh1fk3qHG6CTG3009SnYjgUzDNWH
OX3nQxJ72IAx8SfdNsehrbtdy5F2I4Cuc3yGaw0yMSv1u7w8GJn2Z4U7yQMzIldt
ytsx56ZV6g6dAYpuXtvlIng4epjTxieLNwf8UGGDL1Rt80QpqxRtCLfS4Xdj0eVE
HK3QLvQgQoRfZRWl40F7xxnYykKl75yRHA7yawaLYbQUeNUOoYMca0ZWqhbMFJCq
pg70orl1vo9UEtaiyAt1UNYuJTlWPcqDXQTMCwKrJz0s6lQHii46a+9GhsQN5r1n
ESibiUUqI1m3wN5lH2b+F+51mVFbKpErLcxRjOO3WDGPjwxuC5wdLOil8tCTlIjZ
ZcwcJ3i/GNRj8xzpM9SrYaZJzXkcnKbb1p7G0UITrQyFp2uKB7Sp0ts2fH9kj7LJ
peqmH7ejCE+VT8L8OSm95CL/I3qdzrSrcU0U6aoxRiZtmjKvvMFFvot8gEmChj/F
F8PiEYajJAdd0vK5RFOKoyh9bAEAe4KdsCu55mMzOxtairjkKqD7ijuqlOtgDOqO
Q/yEMv70lnHftqflmq34hEqtnEmDsK9FMCYfv4Z3gHrYQE4nLo3ZhnhQdN2Ycr/w
RUrT61XoQNRqOIJ4hvchBtv4Lk0KwRw9Fpoq+Xk9iYzfvu56SDLOo2WMxJJ+41pV
iH0HC3HENQHYyVLGJgwcwbxdYc3KFC9+Bd0O/dlJPs5dtzZlHIMB+Jfgc58y4KE1
9jZ8TTomWEKKcgdz+l77TRocRJmtCJvbRZ9slfmJ3+es1R0SBfbyIlQUOXI4ERjo
r7GVmRRzClR5fDxoZrmkt6rE1eHUOVIDjaY5io7HKvEnWyxyM+unUUGqYuOUJMpB
/jzpdjxicvNtxh6SKUmHuIGYBZUHt1Qo95hdS5TJLa4YjxrIsgKg38sJMQ+TP/ad
8Qzrnf1PvwM1eTXCWYYLucZBC1XE/sH0JxdqLyj1AzPcXo0EiB6CIaV8fVrR9WRQ
hrPWy7JeSsLQTOCkTC+CufHfIT4nstyprBnrxBi/SkFxZJ4ObCdb50ptGqDeubBE
v5m3ANDpDi1rjW7XgbtMxzMtz/8OV/4adC4y/4cOvFGLPBGOZ3YvaX+M+uGNrljA
ukTCbJMUUUqNwT5nQjVIrfuhYt2IOt0FjIEYOXZFeVtjG9xHI7f1k5Yc28Mpja4u
psyMkQvK+dhisHMMfaliXkQonimXujc7nLP8t1vaqalu7etgORXOhm/+lysElAYe
wizRQ0GLc0CevzaSg74VIX9n77bQDrR0b10qmVvwbZaqOgEo7RvenDncYwzOOe0h
8pzAG5iIxhPr+fQi+8ZK+0ksIyWsrpZGr+BwimEZiPPcdqF0SWtiCCshsDjPPnpl
NNpSEjEHjc+VWL9luHRUq2NlV7u+MsFHOx3wfevylkVwQ5tVELve956IHNwcqPoW
8lKokHeKXhqIsDKOzOt0+xBZqxUZFXjf3G147ESnifUfd46EbUqpsWKh2/bieJ+v
B2P0aK7xjvuVuPv1iiJFqwmKxwoJMJVUntfH+MQenHQlEkS3E8JxeOClkXfYWTKh
fNuN9MZ48ljYxfIHdmc71A3TRx1VV/RC2DXDT5RqKXyYpUL6qdozvIWNfVUxE3oQ
94odNhzLHfXjJjG/j/Evd6NovGzETTtREeiHlajiw0eEcP9GnP88iOfUAV6TR74z
af/gw7NsxqD3BNpNxh8do0CYIPT1bbDic1TF9bdqgMPEbUOj7esG+35hldYetHez
IBzfg+0BVsspHbX/Q318BwpthRmW0T3HLmQwjug0nysK3YNA1/USqCHwC45zLCxB
QvxKo4STnFSkltzcIC+zWeREnemUVrhmVnZxpbB+wNhKtDWeMEYdUHkhySMJO3Be
a56j2qF3/dDdrn/6opLTUs3WJNVN6sMW3uCKPHbkXYH41IHHGC4eOjTWwk6rUrgZ
iWJRT0wxanf60EM4k7mfVNJqT9F39XP/Q+BWr8duKHzKkXnLnp7kZ3qUeKLDrtXB
vz4OZsPtlSD4gySVoX4edFKlSxJYSvQO6SbAB0oJ25p0n9Dn3kqMvIr3dPpScKt+
RoKbRntD4IBRYSnkWXk+y2ohMzFJDGUTHYV1Ne2pXwrn3f55gPPoSm751wSSeLwt
/YCSzCFy1tgB/OWuCPSbyA==
`pragma protect end_protected
