// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:24 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ga2LKuSYoLpinbONvt/meUOZxWYMtpv4HNx/v1T7SYZBZgw6tpB/zLshqnSku6Ig
TsvaGviTvevvKNrRLpCLl5hSmItf10tKX+6IoIta60G14cwPnSUnHI7o7braJ8y7
18OzCS4ON1Fr1dMzbqwgpgZntwbxbp3qJx2GsXAppls=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 114512)
5n235reW92TiSK6oiNqaU1H907reaTeoDtouLMkJiY1O9Zkl6XyNdnq2whHXn3J6
i+KV+S6LqYi4tdnp49IieOoUOuyJVbnqAXUEA88ZCzRWZiAtN3Iq4Ka0cEQKokzk
Ysjat+L7eduNybC0NNwCXHZk4p4A8ec4D0VuYZ63iYJWr3SfxfGVAkH9Cjn719AW
kM2QIOdeIexmeAd2VRr9FyIzucKvKUGHEvQ1i6gEKRXFeRXOlJU+8m+OX3Bvmjai
I9UvC4YUIdX+EW4UkWc0nJLbvqR33ZCRpvZ7IbGj5aFxEXo2/MZ7bG8K6IKNSFx4
QnU5llnAzFtj8QqIGfAOUoJA4i5Tvw9KTldnkbif/fK1D+/DFB6rT6LtpbRjZIuG
8MqN1rLD6xWQ+tBa6bVenVI5xdVpqrFlP6SSzqKTqL8V+7F1o36GWZPO6DaZhrB9
TOacLh1uOjbdBsFbecMVKVuqZ5XYJsdDqjrVnR8HcrQuuvNZwObxub58IteH/gFW
LSQIBBIHrNVFYDF4oclPvhUhNViI77dNn2aUDbUvv2FVuqq01fJ2JP/NjR6+ubx5
J+zUYqBao6XOwMhn436D004k+VQljjVmsDW2Jm7F9mOlYunggmme74qF9ytPJ40I
ErYmChAusMRLiFZrY/3KbwpDlVlLIBtO0B5Nlww4dnw/xUyn5T9BPt8IwNKkkQaO
PZGJk8IdAy7X3DXN+4+8g/OTgrpoHsFNn2ZWbbCLc+YSjht9zThm//ZqWOAGSRrr
vV8kg+kNfvqJhOG3sWFyhPWey3/avZth6mZdEEAdN1dqxsewxgI3DeNQgWZGSbPd
sMDfHBJfCmM//lgZIDoiHBjNVCdGp+b+ys/3LfF/n+MvuitzeoFgaS6uSA6IxYdZ
CwoW8JQ1lnlrhCdfWSYhFFw07sHR64iubQWKz7j5wyUdkQ6G5Ahahf+svBG2iHuq
wlnD7YxjZNCBQrTDCx2rCOekbgJcFUVsasb24i0gwjgO6p/ZvKvvM1qxsBl4/HWM
OjaWLOHEeGpH+jyLewzaPbK6d1Uihk6Dg2hlUP0KrtmtkhThWehizEAbcrfWGWRu
J2bIWAIEFGq3sp72IlXuToNywHE+PGz7hOUaYomi5RFbWKQ1bUoG+xpzpyfiplas
NoLrSg4L7cBDkfMY8gxQ9ttrEB7aRlENIcIxG7YxQxCmWgFZx5ntDIuAUZP7E83Z
34DHcYAHLmlHYskElx6K7hDhgCRlMiP69zOGr6kG6ih9c9uIptgIMEQ9m2hj96ZL
DBEJXvNgxdZdEygso3DjvhKnX2Qx66UGbsnyyhudqVW4ygmdW82q5YNCrIzqIULu
hDegWxBBjyBNvg8vqd/Sh/MQwSECzE1Ydb8WljEaligEYHPFkUc7u/q44SSMOsvj
UdV7CeawtaIiO/72t/1aumAtQMHXS7JoXcRTgUVtoPdoex6sKhoMAd1lARrzV4QJ
PunppHxmjkRYGW00ha2bx93U4zSc0j62OEVxSxXoTI6tD0NTbgkSWxuK+XYfS8vs
MprEHlvN1uaXisH0nM4ld8AOtU4y/HRZO+yUb7raZgIg4gQn0ZO5gMcvgpXhNLtT
jTB/LJrs11EhQaWe9O5DZb2G9+iwQz0l0f8/cs/5Fm18YbGy9REtYoD5VxTNuMHS
46bVCaIS4eIbfAjc9WCrmQU1FQPxnROxnfMtcyc8nO9l3qrc22kT/KnifMq1n6Cm
bqYvg/pRfOZaUiZeoClaV6UCorQgGEftZCxN+PGWSogzYxLCKGnqDVk6DJZZKoza
VeLkgU+jsHElLsXsROan7nUImSwOmidKa1d47qkbAdgdPMHj0m8BYXa13l5VQzIX
o+g65f8W8CihWiIaRk2Xlo0JaTRyGfjbNqg+4G5xHPTLLY5U7GhuhFTpr1u52fgU
zABO7oeLKMexVN5HSI3lwfeNs+gmd08B/gXm1I/rVSkOwtUSthXCHQQePZ38trOL
ZaSEp4JD/kjPI26TS55/u7fe3nvxtVgUattv/Qyx6TvRVXMkghkrWChC+o0uiHiI
lEyExyPkINyER3jvuJ5KsoSk+b0rIKwWeqEwRGNdUebOB/4jTJvmgFID/X6HeXgK
zjvRJ+iwr5pUiL3LTKoQaoxGE0+XhBkVE6ExncDSPp4pGrwEMaiYESORbhZoBt0v
blRyuM8mCv65vjfnpwrGIzFoWv2+2fSrYsaTXtu7vlYm0Nu8sub2aJmMUi2llChQ
sJYYuSvOwErZAxWDquoL/0f5/KcRmv30B2dXnNS8QpkAtSC1Q516Ilk+4nJnAysR
mee3Tou/H8P98aVcURanwG3Q+oNvCvh0R1Px4VrnqFIn6ov9DFChQAzms3NOaViv
tVE82GWOvUFIu2n3gxQV9OCOosAkYlCEXLT7wWrnMtC47enbFT+ufUx6nNC+LGLQ
c+U3T2zLC/8ZwyJemEeGGa6DYcxtWEMGKyHG9dtokD7nDC46EWYWuUnbhoUBLMq8
QWmeoUkiKa6JG5LLogxuvW9B/dZB8ha0W6zIeIZvTaL9I1dbPKc7qBc0Wr8hwWvs
5Ia8iFIZEBbVcFYMzjNagK/LInoVwuwd30aB6QJs86rvSqikt+SwtZ00C3VdVfb9
Y5KCfYv+XXFGAhofE/N6J4S5QEcsKiwc82lsx98RTyO20DEQmCP/iw3CuYa+YM70
bK5QJsmBfRsvTL5YsS0HqU+W0Bhi4MgnyH8/Nlf1wTCzTzj2XfKI9rI12UBJ+2k+
7z4HSMt9S4mIQfksA7L8Ystc5HpREcGGwN1MUCLr8wKAEs48Y5Wx4V+Bn9uSYKxv
Vmt8ns+L9GsTyfMr2DIayT/kZwGJASiNdDd/a2NSaQA54X6n3Dg/d4rGcxFT8jr8
kVAb+ZtnTjUgeg6Z+gHA92n0xOE4tRSC8WmnYXitvTVLmwYUdnosrWUkgTeDvfXI
67l3ZXTGH3yfqnwmwUjCqyCDz5wH+BEElImviDEEbQGTZgWyQHeUO2HLRnlnoqzC
UznqputEiPVvWm4+OZhezFOWlEj7bC2Eym2ItTeiyEKVOLaqzBCi1cB9+rxlTl7H
YWdueHdxjHuVEurvkyuWaqtB44C4RZNcPAZvi3bG2RU54Zbv7mUencNTNYgiRB/y
f29KOb627iX9xq2iyII/PmFIVtp5052tLjTAkZNEv7plQ8k6YdUhJtEOwCIZwXBj
Pnb4yYyUCjsFXdsEHyvqCWoAk9BlCRJaNYFu/82B9h1CXTibWJoPilSOpFBbuJWN
jDkWUDJToc5TfTc23IjYc8IkfsDMGQQ7EoNGW16/CARM/U/Ajb/CsPoubjhRhR6l
LnkV19f4/1TIvXDc7OGWk+avTb4OBTe1RvUoLTiyVmkPQ4l19bQa1uvOFaNLBoNg
/x+Y9Y0aB8mRgaFEloM3bsCb0zislUyJcffoNLct8LWX4kWKsboHNy43hlkuhY5U
lNCeeBomzqNPlcLF9bgBIfcg8Y5B/xjpWOKUyw4HL4rZFt+cD3TD5loMDweHbeEr
W/7A+Xs/p03aMBOukfnPJVwdnPt8OmQw49TLk/JDN7fu+3LoEIM8NPkV8Ld+gEfv
gIiOj4PPDNqfJv1NbhFpRnobIWMEerxW14NHRPPySIMmttUuf+7q00IyufN9GLNI
JLid5mN0g/2apA3PzVMMPGjTMlTCJmZhsvC+zEciWS28w+0WuEBrWQLjRNwPqGaX
nOACBuJkObyfCSzUO3mp1th2Qch3HBCBuugw8yfSaXkyVgZ3OeJHASorW2hz2Fps
lcDcODdXOxuKWooclsGTmMDn7JE57Megqm86cyviBcucF7M08Gmo+Q4Lg+kW1gV2
JflgtjL1qVqLxYIty+IiOuJ992spQ4GIkLlf8jnCOQbJJVdWdvJo2UUWCw3GLmf0
uIqNgqI1ansV4nGNIVUWrUy04oYWSmdN82S4tWWPJxdE6YfswfMcR5Bf/jrgkwhb
GL6DksMRCtTibkgP83sHcB3tzJXWIAiw5Ac9IVKuw7rsIl/s6Jp2s5Wvv19ypfE6
yj4IsL4z0x6SPd01IC3di14I1MW1Lr6zfe2K4EJwH0cuhGQuRqiRsSoQb/H9qStN
Uoj530TUNuR0KJpw76QZu1A52zcr17slxlMa5uBt7//eXVMOoxWeW4gQwP62PdNy
tlxRHdNz+tbfQEZq42s3voCKIItUXBPZklCB/XOjutMYKJGZt9BwZ418WITTwR0b
L37WRq71LaI7mgE9Hz6x+JfSnKW8Ok0lwdbrF9e8yNRBcFU6ys1DaBxn3cV8+Ekq
JkHFQssJf0pnADS7Fqw8fEpVnAypcs5RkohwxLkwuDKMtQkTX2DIvJx0P1t6WmJP
0vwwAdlMaFp/TVcrJU86m+Cb9pfmHk7kkw5ZWXHNd/TTuU7gXgSf5w0CrMC68uQE
1mu5K3Y7TsMKIYLNGXvPYCwm4eS6Md0c++5pXfBKytztk4ZqPcVQyh0ln1+EqWYQ
LbVEOiOvB6M8Cz3MK2I/zMY7KPv9gj4xk9jNELO504G2TKrAKsQm90bL9LHKio6S
4ld5urEB2vAAwduuVeDBkh7Bz2gk8VdM9vV2IRfqPKjkP6FsG9LzuwH21KlGSJfx
azuaFaCiSrddXf44bW0uWu4vZ/tPV0FLiTt+Zjh7QmYGFg2QLQYO6Hbk2Z9CqyGl
6MIXepG7bCtUYL5z7t+9x66tnkLuyK/9GIcBU39JboOQpClwAm1nRB4xFo8xTEQj
5stkK6l/gAF9tQsELbUKlkNnSQhj2XIRaCpmnnuhrPaCQlgC56PWz70H+2aGUpt6
j/ubyi+lkOJZ08pYunyk8ORm6e8Yh5WidcNEf/X6OeB/TJQNJ3jPnPFT++WyeseP
VemEfPStdnM1ww3iBZTl4uptlCOWJcySBSWKL97NIF6+Ec95bXUaBLCBI4qEc3gK
HHtCvN+XtdOaZZy+UP8r8CQAouYOBGJK7xGwYgjkylSmcu2ItNEjCtWpXqMyk9o5
+XNixbb5nLQKFQ+EYOUwSEp+wBTAbqYMYd1E48n5Eg64z3XooeMy8Cowvt4OWrHX
0bnb21tFgOKKFIva7RVkkcuH68u8HBBKv3jK4WnNSxGIXk3RYyo6n0BXVoqszteJ
ZcLp56ReJazvKD6enbanBiG4Kl39u6qFBLHlkB+Tb4jd7XR/LxDuvV04cd12nuwe
jPzXzcdjBjYYYobuo2VF+XWpy1G9DrhmzQ7HTCjVxa8pJyXyhe4jDCs0mwbX1Ayi
NVoM2l9s5r90MJabCQJ/R2g2GCMiaX5nKE4UIr0Ekc2yVLTlnOxPQ9eaIx3DgDyb
gJzQgiU8BF6PGdCwA32dAxZQfji1NkCmSjYOUbajAhe8G6vI3gKj6nZtObz4xNBt
mALyQ7u3mphxl36RPrxzLFe4p0nXuGuhkx8hXBBksyOU3mxxMXlPapu4sIG+b6Tr
7NM1Ub8M3ehhAeNNunF439D3F7/ew1N6fAguHee5jSUOihGkFmpdU438FOSzgKcq
K6/a0mdBbufQQoBbb0DJdaks0PI1kxM7vldlecH94MGNb0YbqGJ9snK/b/SNHBzp
QODqwQw8nUhxZ64mk3gM3g5k09WOblRPc0m2BJ8vGB12ahbgsXlx9qoQLnJNXT0Z
MdxkljsA9Ib5G7mDwrmNvklCKwBJluER0OmCUUiLXRMEpWuprcQTi+ki1sHm7MXj
0gPue04KdD5c+Yblhka08dQeKLAnoryOM4Wzejw10d3doi+nmAmPwBnMLeVxCELV
a4hIk9+c6Tpx0MqCLIjkrZ6lMohVPh4Ds59EDaAEwAOfPoVvS+vYEMDxzzpXZRDH
tK+mGc5Opflp4vfgruulaEXdk2Hv/iAvBPtg/FbDra7rvPiLRcvO6btRHQ7+x/hT
fERxWnRjMC8OYcAFn+ac/jvQthICUBnSYb7ZGamMYf/YesEBpWOWMMtlPlOK+3ea
PPgK8mdnYIuHsyX5l3XDMYUNG2qwxZlblpQUl/jScxsj+G7fml/xu7J4y6iepqxu
eeUfsbA0qshNhELqjGVvIjasWYaPL4cmUTUt9J4W9W1tlmaOGMWNGWlq+s+CAurh
JbmjHCjsYv1sl/vNh+Zk7UhQLE+ffyugm1Uh9uBd2zaH+fRuI+qkYwD1fwKs9uXs
tYenAQ1hu7QpL9cuPhUibACem8jEtMEhCgO07HENYvbWflZE/fDt34eVOlNIN66B
pQTA5n2nIWj/sJjbreMNSKPfPN9s8Q3q4znzhp+R276ZVY9mQPDYgBBvVqjCEI6D
mXuz+MDLas3tka5AF9aU5USO6ZyGWBgC2wnp09wlMGfp62a6/KcwYy4dMaf4klXh
JdtdHT66HlM5udsPOqnFO44rZuUpzg2L2hAJpS46sxwaiTRydd3INp0Jig+xB3J2
KQdccNcl/Ab5svRlcDDcVJaoZetOkq6OPgPl2W0nE1NKodYxfUBsQnY9uEJvOwBJ
cQmYtzUA+SOlQj616O6O96dObln+3bVYB3YHwMtH/LTJhCgKcZr/uHcuO0bj4n//
NYoZ5z6SrdyoeHVBUgDdG03AV7ffMfV+XvcWw8xItwY4PXGRMjeCCFtunYCea7kv
K6wSxA3kqSQyfDPCTSLFQu5GVypjksIQJvPjJO/9JKUZND5oMAlz3hN7VfLr3GS+
AqA0GUX6k0wPD6y/uH8oNEfJoGwKN2WYG1RpFI/2hubeycY2jjXcvhSIUfrZqX1S
muzEisErfAOTzGKAov6Ph1TRkDTUL/KNKAn5qCZNdUEGQtV9wvJrdIXdrgUNFLJt
+cmR/YYLFMYq7Oz5ANOkzKswVIKsNZvr/vyUrmEokGLCfvEY8J9GTktng1t6yRAf
36Ibnon3TMXpbdU7RHoaz5T5bfHYbRR2g8EMDWUk4TBw3ATr+xJLCzwGesaoIgPb
CveziVPVgXRJqxjX77JbDv8D4MxfqW9L3hR02wOvZiPnGWswjDZuVQEdOqS0ukbZ
qYT2UA8rcATZ83Yfv5R1L5HudCfGrZB6De+voC7b/Z3q5pFnZfBlmqg6shIAx4c/
g8O5WacgLiuVRzU0I4fg24YuJh+guiHzkrxLFxmVITaZX9QMhe/ePguB3TwiY+wm
EJ70TLTGeyzAd/ijdFICDWZ++Ohi6fcRXscNPfXrjTWiAIp5Rddb0HXAFFX5FsKh
uOsa13m3PVSwOrz388DpvVw8sB7wqkIOKHdX05kTk/RiNUXyOu7DvIA9Nq3S0b9E
Ncbp/mywhMjbknucVm/iwlgO9o61FomoiqyQfzmagzguTaAekKdHkZr/8XEBqCto
1wklxyqxSkf2i15DBISpXXb8Z1bErZ5bA28j/LRYfrapOk7pYtj6wETVfyxtw3IE
0NDMicGzKw3BsBkCYPMOZlGOXEzIdH3Uav1cFdro6W/kGjcymFYL7Y5LdfBkvnGc
6qyNl74z4SQ59L7H2OrWFgMrFtCRKlcfGGqARwbq95qASpzJAX1EGrdYAxiV07dp
6pCq4EZr64sYKxghuEZ6fK9HcMwE/K0ZPZMHU+Ip1LbTDjM4GU6KJ/uEVuy8h+GU
/MoqTkXjucsGMFkdsz+N8wclnLNZp3DyFagZjWh/8D/EF+5sR1kdCMvguOmQQChc
8RwsZ+vlFeeEbeH+N8SMWWGBcEjgtpOaiYfLDPXPduaq6SiNtyDcGAAxTTh+625p
B+PsZX+p76ERkQ4Ye+H3h15qEbqyDaeObdJRO4JinY4lsX8gwlxCB+tkS/xY5FBQ
/HNCDIcA1EsjsyqB4mJ2Ej5Jmi1jWRLyhHH4ctD3+2w3a57lqFzvQQouRtDe1ScR
klGh23VDrWD5zcsjRzJq34WjR/Q/6ueKbgMwsgk8IItVojRfT5qRa8z9/rw12XDZ
jygbcE7uxKASh+UBkKADr8hbFUm3NS2+TU1znQBlfCbV9G1t1JkH2obDVC6F1HbZ
xa1qJzM2xtCN5Fod2zLdJHcQDlhVnSICwV4DLPKcuHU9ZHDG9+av/FqBcmXDzh7G
LetNO81SPHnaG43YMTM51FmvEHNeXt4O3wgq3smO8kHX9912Pn+qBmRh/3RyUT8x
XrdBd7vYDcb4j4JDEfBSuwN8OvMQMWPO0FGisiWoaIGacVU3TSv0k3YgGNV3x9wL
AKF0FVvYQ4rFHkVU2+0Kl7H7WDZg7JAEG6UhHJT7gMM3d1f05OVyyYAaqCTzuUJn
o2VQueGAUsaOaLE6QWq0FFtESdZYpkYJ1sAFAqV4LUMi8UfG0fLUb8FI4DgeQfPU
JmKBqz2B1p1irf66wpfCYSO8ZlBzNn9Q5azPbEaCPYMDYu04C0D0HIxQYAFBWqQi
Ce4YYUKPD436Fqe2OlbrHGCU8jk7k1mxF2PTkDSpV8XKT0j6v5iZEdsO4OL5mc/W
kUEhBpNq1wY6nRyhX8EiClbkGdl+jWzD44S6TjaWDOUjjn9A/bPSe8pUESX6w+s9
xeau9g9o4b8kNq59voUJOPmwVntJ/7qnIUAixx7TjRaWJ3R9TFWnzB6K8ojUBlwg
T3WElm5WLyuXNRc656BLrMeCfDlGe9Auc+2acnZAni7Y8kKweItzgQxf/DoqrJIp
iRytARUhzCZlplSdReeckS7uVFEcRqz2fXg1eXIZK/BBj38Zw5QFtiAT2/z7tlk9
+7YewLRqSj/mdQDQ134AWINNKeqvqOYL1AT5HF377/Gi/8oHEFhCYOCHogBKY8eF
0bPj3ekW7m3vdmuU8RfP9mE5Tkz+CoQELIY6egsgSZsbXDuqcYcZ7fFfCXxeGL1G
YjLimMajBkMRb83IgZxL+ghjZoclCIHT/3nEH5rbT8ZunlNqaLhdq3vOidqDPiw/
Y8dNy9Qmgkj33l0Fi/FSawRAHmMw+T8Yxnv6PQZKQOXkoA+jTdXX08e2nnky4yN9
urgxM2P0zMtKnAT19WsCCPROQK1zFTBnzQo3hPxCdTxwS1Q0mYOgs+x6gIG1CDlv
0vNpbparqya4Y/BwuL9aeZ9r+bE+L4EButi+SrfR7St9TTunYX20qksjFJTF84Mk
EI75olBN042zMaOFXN0sLMjdxG3gtJGHBN7Ktwt9lFJ+jBBUQfEo2oP4/+o3f5GS
oe7okrWLplDXTwrWElPnyUzV7tc/H1cWVh3SwTYJUL2XI7eQmDeBXtQ2MVJX+4wT
fUOuivGO/UPrklGQrE+LfHZfptdcsPMa1U7M95UFltR7RHZve8RI+GKonHMzq1Ja
r+PC2E0+wviQnJo8FBV01tTgrG1irmASe0V1zxKezwMa6FQNEXOpKoysFRbY//gP
99L/vihdh6XBxqtqy3RG6PMozbChAcj5D3+SG+z/AVngFDGLn2hIHXFGCDddSLKO
i1ZYBJqVmLGmthAIhjqOrPouV1iXN0n7a8V3l6zaxoox55QdRuQzF2jSRkzRjQT8
wlMNbebqFuCnpmeOthkA/vgbbq8fZAlorDtEbMHfD5dBQ47Pi2ei6TuwyHY7bHSY
IUWjRgXI1iyCstOWLJBWUN67GR4CtBpkEEYoTMunTbjLt4YvG+kEyg77ek0YUE8W
FgV5R4nYdFGmYvlYauAg4T4pf+Jv8P5/+ucxE3lXrlJ+JRm4WbKDrJYG3k0Buh8o
Z0cEc+O45ynggMwq+Fca7rlr/Dyv3oug2ryUYxUCwc3zSplpudTIqIdInzEeFrYB
HHkPIEVbAQB/+PNDgGgNR1/Dl+T5H18yBM5botnBz2gZWdH8YOTHPprXf4p3lVb3
mmB7hSQeLJnWwHlGbSJlB1IRXxeSxU1K0/qlGMgOn/LfWKMHetNBqScfzNJdRG/Q
kFpZyD20/26oC0AXL3u2ydgwK31Q45bze71FlvoNSS/IFOBmBPsSUiKjzaKfajuM
6AhJQcXYCLYeB3VGRXSQT3D1AKe1G2Utbhr840QKu/qY0sz4P/NjEiOqLPpOZya7
Qu/QdHvF73opTlDfO43l7lTvskxJf2t9M4hC2E/VazD+My0DQJy+iHgzIRIN4BDP
UN7Cj3oM4CKuz3lr2NVmokI/Z/wzOJgsrqOVDRU5vxTCqE4M+VLIQTA3ZGi7nsMH
cPhKW/Oyy4D+TW/MVnrfS7QFVma50bU+a1w+HPJ2NQdICxKHtc+jjYs/CQYRAW2X
dNBQx1okF/f4gTt8xEv6KAe7yggLQqDZuMYEUdgI/9l4YdE4r4KmFspPlHNzpT4o
D6ay5Ux7ll8ELuxhFVhV05Cqgf1AyJRARKkcpgC3G9dJ8bd/V6NupbcM9+Iug4cw
gGvvdbuSxaCs1gEQrgxdgBJV0T+IFWKpX5JJeRB3Ko0Mxqq+RSumbNSjR4mpmo3k
HA1GfRVdZlRXTsGcvhLMqThzNypkmR1G/LZd+cklIwIxkkG86XOZN0GPHifjFHfR
JJHeeg3wBWTL6jB22uAnUIkW3KcHavxv0ZhluopnfE31lkjodblcGUL/EtLsidk/
70pAhAXK6n2ghRnS5NuPFmyMy7Krw+idGUheLoU+LluJacUKceg+uK9d3KXNjo/c
qOyTWZcMCWdv9NS/us4jv4C7GRqTMm0JR7gLzSDUHowDm3hrEQNuOxmZPjCMN0ac
Ko5P7y9m3m+hfD43AFguvMArUZoeIygi9IPO231THc2NecG4iCXO1Er1yRs9cOHQ
UTfKs1mYG2lIhiNsYQozOsjrjLsgN7gQTCLCC5xNpuAtj000kaY+PJvrB7wjxHes
yHNYrea9oyl+D44yCiIM8hDsBvZfF8yQTzfpYzfDrWp5gPYgslNwrfS7DGTNe13K
MA+GjR2uCkHg2jsIEIxZ23AeaUQRG37+6qHl8i6EBtrw0AxVtob6hIhlYjDYUgpU
xve4PynDu6aEaAIYZrWRmMBLZoBKm4SYCDyBOlcZ1sH++1ou7QZ2iTO1v1/MSsF6
mrmOEplD13wK5PZrQAv9FA7QwJ9adYmx1mZKANB3ID3K2ejU+qfufBFIAhZ5pDQf
WB1ptaYRLCiJngTtcOZQV9biUKujUBWv1Hp//ziI+9ONvWsfAbMLwfn4vq/mz5uz
JnA6/qwdHnQArEouiNz6WWU5ETxIeG4vgCLzGsu/QNWSqsaVnhM1VvfpPyzssGUh
1hdE6Wxu+plzk/FVOe1z6M91YYK2scRH0+4dCz8jN6Xkpt3jL3ztOT5cLFXZ0Sel
deTZzGbUfae8HZ5DqyJFwwl3seYatvUbrwKUlRNp3vpFHpvWcOLa30/CZXZ2fWMH
YQWjG9iVijYhWeaZkudZnvD40ta0MmNFAc2YJc4OeEpCW7ell6enLXIMjxQRpTo9
99heeNtBEx6Yp2MFT4l0StaZr/bGeWdvMohAaYgaocnLdOmib6dtcp3C6aEqepcw
Y0qCRhsBmAsnfpqRN9RJALIvJ/mUxO0zpwy54rMQ0gqKOd5mb23aA0dNFK1Q/Nyr
wAQ6tEe2l4rbXAleCDZl2mEgKb8gtnSNKIHVXVbqL1/qWIdZZOjphmtt1uR50F8n
hq5kYTvfnS5IurSIzs7eQ9MXnV+6EB2XJmpxeK6kjVoP9lzt0mAMiIJIzo1ECZG5
+Vw/IS6eNtiDlRh6NBuALHoZZc4ceSKSHYaiL2vTbkT88sjLXjcCSYkTJgJG2XPp
4EqThpphpLd/hJr8ocRYuCx2FoZot1FUOn1VxPA2rq2QdjV1DakdOmaImp/upHik
A4rWWcs7VgxTCIU8jiHp6XkY27i1waOtM6RuyNlwRLPuXTHYnOs8qAUvbB8zgXSz
OyLPYCzDZJy6cduFZmOP5I7d+QjRgyyZBxyM3avuJLQ4wgpeCUaoo1ZV9P/R2vyX
1sc5LoN9MWG59YlTA/xJq8+oVEeRk372R92FzY1X22tAxgo47HBwd5pYXxQZGsgQ
Ge7fodQ8Qc4lUK/XzXJc/obr/6nu8Czfjg+N0ly/9yg/b6MO5Yojng6vaWHdb4+O
2MxuOyT1rgd2Buo+CuZ72gD/87pXD27ynYe7RUcLtI9yeuHfYKPCmkF3mhHjXpXS
Ewtja9WfYb3UiisZvkLw4pr606h7FcZTH/acMdVijhv3ev7hl0FuPtsQGhicLPpA
6zlLdCdQtUHEqBDPqc9KgnLxDhQdEUbzUcXRnL5NaABeUPQAau0lZYNE0LClRwuc
hMDWbWlrPxorh2kX08TvKENRY0qRrZoWokHXdpYDgoiQybv9qRGKlPvmYPW6YmV7
jx6fvuCxH8kENf3hTVW8K40RRPgpeDI6rxbexTH4WyfY7I2LmWDkZXw1tbl/2b6h
iOX8m9dPnf9zSndobVRM4jrZcgowgRAEkn3zdwn4HFMG/rGwW3yOocKm3/tF6jnM
CXiw3OAQ/w9Q3BPaYfwWxZrXnQZf7r7Yz2A5AM7xESK19pijTgNkN8env8iozptf
93KXLmfS9mlEbMefCAo1TIcEdMxuf8aD0voyaGRAxPfKWkMJYGMu65WNPWoiE981
GXV4T2/ui/o/Phh2MAKdkGPvLDMnc3qCWquaIzQ7x4lqDXagcKvxaN/CIr1Ar81B
xGYbSFWh360AZNDTjB3RUFIhLG7TUYbM1vxtbqSN/hC44y+6HVGrPKgaao9xZ5Oh
jjIkSv3JTXMVd9FxpYFBBdUOXTIUpL+y9n12k/EMfN6mYRyicWw73/giaNet//ez
8lDSa6WGqah4/vTvj2sbEohfWenKbxSTlXbiMJJ8NyKWiYud6QwI0VCFu0QXWzfl
Rms0XdS/ndrS7dy6xwiVbrPi+ATI4liOy6YOOTZEPPJK8r4rzwMXtpYtnW3T/LMY
JLwkeXTCE0xRLZgtNB8xDUdbCiHndV73/aQAc61y9cbgTSfIQG9XeO22A43VzV8n
Jnf0QV/OfITkSz+t13EpgnZVKSmYzx0ioMzGW1djyeAuto3/kogkP14Kk4AZwPva
ZS/yTL2T4o8LLtPcaWWs29xdQTNvkIwyM53fWkM2Mdt/LL5/RdoMj+kU60ztFg7b
rLFbZW9AytS1n+1oO6kqP1gvxzYoRG6BqUp+MCT4hyvxgcb3or2z+Z7YYzBCY6sh
yT3otxqD2l/qYl/i6GlilCA9FqeoAM7bnRLeHvhdp1xWIIU4A1pVpECYgbMMozld
8gSEkMKXN7pVC2yQfw6Cu46kqeI9wYB5dw8dlI2l9kDUJM4WjwiXrBhqVZmSkLpZ
IAjMFvuYs0gg2jdARkFMEpUHn9SlRAD/EIO3cSUru+e/P0oWFx3MBhpk0KzozZ81
vK1SbW81tcFjp69FsyAia4WuaSHwRAojN7gvfUl4LAICeziiDwnPIavTFtK4TEQu
t/xiv4lyOqfvUJ3DIMMVZQAOmVpCOFlS2D4zbW9hzNYsg5drbhFFBUo7qMryDTj2
aRSURfO7l6xsl9V6ZBwQ7phpyEiKTIQ0oEs+rKzSkzgl4+MnnauKQu7eyewM+mZe
nauuzDNFAeOurMEQvySz0ylUm/HtAter8HRzCSjc8CN0E8uUSLFo8meH0cMaRi4D
sVX2IjVePaGtKODrvQIOZ0dgv4ZiNC5p9c5Wi6r+3Vj7UlzmeerHTkOMRb/YyJRr
nvNO7VeADAWCbseSt+Tpnluj8Fg17ZpWs4dDEfxDFYQANko4K7LciCdezD47qY79
a4eOh3/iLNA9D6U1wAn7Rf75D5yG0NmiqvT6xAvMgLRMgmDKDC0x9sjcWKucGjtW
z0OSEa201hz9Oq4tNXeUGMUrwK+jOgOIDLVn6/pkG52JN+HByJTCZCGFRKR5yDM0
tdc6lQsO/ifhTRCHw3eqcDF3bkUv+qHI3rEydLcwOLCvTKzs7ZJWVDNqw/PBrDHl
g2W2XafcFvNsPKOD4pkue96swEEh/OYHhGqWsuVpt/imElY/CRl0Uot6Htww7QXr
i2RfTmNkuDIRY6ODSV9DxJ5NVA2kboWesddreukA/g6MI1/GBoGoomhgt6hapRAr
V5HMtHGZuSm37BfOwuwLd8yS2jFMG/MxR1aqQutpMuNo1Qdz1Lx6DQWG5kZcERnW
fdV9Xm146pb6VI1Puc1RABliYo9PAqgmw2xWB+WMJEXvTdF396kaVTHIxaVcmbvk
IEFZDPV2kBHHhvIB6cmJmDnEd+bqtH8cxV7Ud4ZkoqNEMKo2j2ir76Lz/RHMQsB1
8ZEJXUo5qr4lW7005oi1sSKKAY9M1GiLP3u37ENb9wP/e8FvNx3hsCs32DCiu/Z/
cHezFrhYTx5fAXynmhPA5UKWvIVp/uXBgU80Im3jM7tp2wOkquF3rn5gN01uF8MH
7GpvpmVtYe19kB0LQN/1WtVUGn8ENpCXGLVwOXMy4IdO/+hv4+eEI8EqRM44YPZU
7zB4rxgwQA8lSeZJqaLUUUYCKX1G/RDDHJJK6eIyWHdG3GRQsspe/QSLj7oGHwY5
Q+0vRcraixBBdZnTELVujn1zvlWRqm9PTr8FbFwwPDldnVwb7GV+M6Tw1SbQxRWG
n7y2h/bgzkzu/al2Q8UECZHBlyfpOJqFVl0DyGZdWMpQRP6N9u/IzErl8FENPTs/
UZy32okQlkHal9MRpNl44dB3QK3bCosjpPSjvdMotguzS06ENp68AMbigOi2E3pg
fYXDiYuLt4DRFDkrtlwdx76aHpjyKAKYtTrbfRocGeEHbfvKlxa2eQtu5muRStzG
EYobcW0txf8vRUleN9JlLE69Sb3OzN7MBsyFqXjWwACMbkEzxV3kcnbtm7+wPzaR
GDdtz+rxtpwuXBXa/6zuPCmJTHfaLKQCq3lLmCrl0i5fr9J0w5R8EtDCUSY4gnm9
tA19hotFmaeKsPE2HRpoRdlomBK72eRGHCMbN3mX5eSqBybueIAahGuz+SWhy6gt
2jYP1vZDH5qOAFEQAJYS7jmN1L2nyYnN93wsDsissW383IQ5YMCiBfX8Y3m9HNsz
xvFCNLAgUtfg89au9T9Thsc08WWtD/F8Lb7ULp9zPgBH/GeWbERcYA0zHYxERJUU
p3X6qMbgFtky7uJg3t1kcJMBAAGUo8/gz7QC4uhucCrXQ9Qt03fV4WHqne7eBDyw
bvkplhFOsP1nQUs04Y39vsOazt7hmuNRGvv9aG/cZVL+u0ZvaH1znqlxzNqWwE9N
oRM+8iFXrffZaceuCLI34W7Ier/Bpd+SrF1d8srh+18ydCHhs7XZfsdms7cNK8vI
U9UbdEDCE29ClE0Z2iFTEqrCqhCTpNUVWwTQxcsYHQB0A0kXXTuEX1nqNlxJXDKK
It6GW+dmnZM88DIvCk5J1arpSo+2cqF8MiNJCrHR71CMMc14FcT4Wi1JdUB5VRoN
eOYc9s2DlzmrFPSVb/ugNNrjlRR3ZaGwED4ya15fRL1wCECly+SBe3dYwCNqEf8D
wOmg0zidpEnNfhcNJ+rMHvFOOADqdy9ng1NrQXHwdA/goBvYQufx8UdU+BcgY8Gl
9edHlWAFn59lCy/HZVR5MM6f9nCzhK9ggqWKjbfQt3rv+43vrQzXZT0KyNyPqZzY
2mUAqypLJCo2k6TXatfrGTy6fE7e3CDvU5s1/oVG8IH9AfXAi5OZvSNPyi07v8kk
iJqbnQGPx6/EVOSgfQICbPaxIf8L01FQZGTGoIQiv9LLRmOl+CC7/Mi19eDFOlqW
MYazbxZdgoYUJs8wTAVw5gtFoTf4R6qdhpzgsjb7+5EJDaH0iTkzh76namN33uN/
geyq0+KVhskQ54mwXUHSXnNOq4yc+IwXE+s9R2NXr16NvGl0U4BWoGsJ5SG57PKe
h5CFz4AVqWsKMAiQyW4fuiL8iFu/rGc0wnoZvmIEsxARV2oksgkJkF5eeSk5MARI
QwxzrACLDhB/6xMOTrFdw6u/C4kklATGezaz6Xo4HXvMVQNR99YJ30DzWq6v2CXm
fSRkQeUmfeBowdksY1UCG7HK3sChyEASGrqzMT17/LSrmqxu3k6RNBVCvxr65/mN
wY9KQ/9tGISPeJx7NknIFCBT2uuxBKzaRRcvymVdR9qKLVjJdIxtCDzTTwWsNxr+
D4qcSnBfstWxpNbugkAu6w1x2c+okwTVSjuSoUrKbxjKqUPBYo3tfmYY7b9f2Bh0
Xaq1MVue7oZGfRntxlr2zGlzo0Cl6CXPKwbm55uKtLOjZW0OxcIx4B3xH98e8B7q
whuSOrmyRafv0DgaEYohlFhAaRDtZViScjRt255W+wJ6X/FTczUK35jjoJz9xuOP
5KgRXs55NA9Eh5jIb1Av6eDmi70AJjQmpICNK8OU7WINY5RZXetZw7mOE/KzaVA/
9bEt5hVn5yNFDP7+fsy03tUaRlnCZbEUTN7nErYFrLUuuvGHEylvKLAy77EUCV/y
tqKFs3LAPotZwfWC38d6QzrvZLVuwhyFNVNz0+5+mPjMPjnjOPjJUqkywRTiiI6/
Qa4Epmmgq8F0zFMIQbvHK7okx5Sn143TS3mGHr4NJLRXr3c/Un+jH/Me2HKXPvE+
29HTD4aIEc8KDVLspHPWlzQze2JlmISuB0C1BNtTeOBrEePZm4uexTEeMkXNJ7/g
mQM12amqkusCKptH2A8bI76qs3l4cEmL4WXP7cs1X53+JGe4SX8SANIC4jMD0Xx4
uGqgBXutiU1YDaG+fcOUaZwcAjUpD1K+FWLG/q6JsO+tW3QxqBsCmtyrnNx/ZafK
UxJOBv/oEZ7WZeKpS7aJK3une0+uEjvhGDD26/p6rHwuBQOA8JAyqvuKYsa+Wx8k
1Zu08oyT3xI+oBjvlVpQ/injYG9vzuPv1aDzELd12Csd35utV93He2mvpRrRZgp/
B5CBrdPlRThzQ3RM4Qr8tnvtWBZaELKiwlTqK2YXURUMYtHFmw5cnpL5+rtFJ+0r
0sglDqCGf3Z/uUNGFFzGblcr+YI8GvXfxi998YQCtIxsCG2yPBu/kukZGEQMQS9d
h23chcuWQ1NNKMFkYDpavaaXVwC9dHOsbMYMS+NKmQdZk/ktyJiirtPrHZiZT/Hq
ZUTCaolgt5H97akcsL093R/LaQ3xsd2rACWpYbgAQPoHkfzeItxJU87Vr+3E1QmU
HT4GWCqqAXfxKZqs6xpSZ+5MVAkPaj07Y31YTzm2XLgIA5XvkIOAXH2ZC82LxXPL
UQD8v7IT5t8s+UK5WiJoOCzL7nmAniOLMJ0j40CIu6K+TbItFziz7ewN5vu4FZnz
/9tV8YIIDYuKvGuUceHIbUOwSM5EwSEA6J8tBjlW/vkEjaXBr/JzmW3ysoFwPxnr
j4pQZaR80qCZvGLlguZCCGbVWg8CGBuDN4E5nFSsAgD6bns+tP7Z1JSy/JO2hgiZ
dkOJfA6Ov+60BD8LERb11YG1kFcXm7vEOZZc8QtW9DW/G4qj8vRSlsHkd6eIvAbt
ZdAld8CvL4cIqluejEE7UF0molVliikk1sz+jOMpSzMm4LAHOAGlAnh22g1LsYvW
fgoBSi0A+ARvJLdQPcfSRZDfqTg0H3Wt1y5SsCKwmBiiH4uOtd3jSrfJNtDPz1n3
pQUWoH4a4N+jzSE97jqpikU4j8Exo4Q0ZxDMr1l/oXP73picfcpGGCOJuLv1S0ip
nTws+eC7x7T2x+OTGUZdQn1x1KBMhxrfCINgNRWHvJkUjuocMTyQeIEWX2Nlf/0a
c5e1EQG+qLzaJUinlH+QmFbjEgNymzKE1ltWCJLgQbMgUfs7NSCJZJEYFlFn3JVk
C3wMLiHR3ZoeCUWuuqnefhmbIUgcNIGCTm8xAH7UwZmP20d9vX0OPz73YZGVOwl/
vXC7gwQLcMOwH9WwJwz5TZTOUGCk9CkvuqWQA7EHmthMInkHoQKDGJWOf1QlnY0D
unr4zSiTN7pR9WV2W6kntfAZ/E/kk333vmvbdwXIBgKA1YsuR1bFgmKZJuS7kJp/
pjp4hYW2yz7F4YxXPxHiH2G+MEgDREye6Z0mEvRHrB6247iVRxTZasJAHhvHFlDK
LjtEdzjXLgLgJlF/7bV8wStnZQxDD9+nlH3p5oxn1QmO4qaNbpdv8LCAI5OSRwPV
obcWZ/TbevfuVImmppd3I6ThzJOBFgFETbeFipOgtpmO+XchVCG4+MqiRPf5zpXI
8QFGxRbRSgXDytG+D8O3iuuYlTRMZ4wZEcTHKYoT1MEK8COQSiXGvkiTDhlcMjj+
WLcBv35FNvXhbkwJp3Bq6t3JHoVdquKn3bcXuNid41lHY9kbcSjjqZhXD3KiYVWV
u14RbD7Kngp+XbnV9Vhwou+AJmVtr5FKPI/YLBXhOoV1xNVCs3azXyNNgmn1eKCc
YfDPQTXdDLBODeX38cbMaFADCIiDeosSjUbNP0NBHLnYEFjdtZGSbEux7m9boXm2
vGFsJ2ohpcEQeduEjJWH96MBDJPOB6Bw2OlgpTebExaa+4CxJkw10kpYVM4HhR1w
8G5uU0ygLjzAmO+gXhnDzhIE8Us5mdMXbR6gA0KN+Y96w8vg1ZhPKEO6k/23QI6F
CkKL3HUuwnAhuH86QxJrYydqh062RCkE3QdHosVn2FrPAe90qL/Fwb3xWf3VfuPU
URoXlSWxQUzVWaBsVpqFxPU1a+3kCbz40Hb0HsLPM9J7aY75+CcCEsn98eoqWK44
BWvPKptABPDnUbMuS75ijh7qt1SzzjzEoYm3F2eYooeOb2Jf0yuWhhedgFoB27U2
zEiwlC1/xKZbmV7UGucINnWlHGdQTMlXcoWUfclDW4hVMwrRRNrlHoQaqzRmMe/y
L3UcYF7coKg/5aFcGEVAZ/9zZjyO/FCnZOfN2HY4jZbWhRG3b0Lrub9/DXI9BbSp
7qEJ0s+Ox/uWnNQCq/DU64jaa+qeQDzmE0j7qOsKJZvJ8YJOWs4P7vJ5LbOW+OUi
oESqSc5vz23CdgAZCaAp5WwHnE2BGtIV9iFXZpBndZyNpTdHTFest8FjTRE0WG2w
C7VwXFmkg5sbV1hWHhWu2mh8y0CuGGk0WMUM9uFa+w5HRpDQ6B8vYUB7HIBs3RFU
Kcdg5dgg+VyFsUXkggX3TBG5GucQgVoNEk+TMnTf5QUGFo01p3ZSb8dvw0cJMNKS
IJAB7ER32EM5zh7c+x5QPDyr8+IkXDySxmgKDYLatZGnYjjwb8lcRE4Qj/nvLR8h
/sT9vUvSNtLrrGj0T/Vb7a+unmXEl0MiVZ0kSGXgVZ3OfJqUlnLHihfJkaCW46T1
UesyXjA1FxnPyccGOULcBD1kmulf5KmZd7QagckPwiEX6aeXGOX5ntr6ozNFslcp
QiYkSJd0rr9O5KWxO28O8l6pe6x/pIqDA7rWlnB46ilIqmwDjMKt2cVYZsiNkWmg
F40N0Becn/HewLttt1yTjPzRDgxUEE0ZGo5opsAEyLmBmAv0Zoq5cTGIa17mn5CR
YBqBksAgTB50cxTdoeBm5hyQ/fB2cXr9FPNEPSAYUBo/aNtrkRvhGhDuQmIh4vQ4
dgm72bbaRZmiP/mbciXzyOpDH6iZWmii4srylP5u9EI91x1mjM8oIuSxaAxEaQoT
RXXTen7tElHcSLT1BqUBTWVBlKiAQaSwkMC660X34bYdgdGHE5u4lySWb/Q2Uw0S
AlDmJH7sd7Qrb5MmOSsAVi/QugyDu7sUJ1RosQOxZzh3IG8DKTci2+pPV9ZA/3eb
Wb1Xv/gFF96im08w6NitZDsnm7flfhSeXmvQ7sKxD05mmnAeIbbT4z4ftFu8zskr
96XGW7bOgY2yJoVEKd9TBQRPiqrjtRQ6m0B+KX6DtFKbRwRsBv0rrvL3kJNc7tlB
AhTiXAIyf6fzwOoW29NoNSFC5maQ+1HLH76Yx8J4MWorSAVzvMla9DXsxpbwr/VE
Gtts8DLEU/DPv6r14/18OIMeJftpB16xjhEZLIu2pDjPsuwAJ9ka6Ky1yuVLqsg1
SNQZPQg/QFk2b9xkN1xyooF8bRhJ3zDx14rin8NxMHDOalBFdHiYla02METOMANC
Wt6hhH0GY0exb86ODtvUHFGAscW52LVgfT07uc5tdm1Fg3dIG9cns96Mh2RbyJCZ
l3G5c0Bis1cTzPTGaKCPdLNAEqP3ESbRBJx79sWhpfI0Ql8Ec65Y2zZq7lb5tCIR
Evs2k5G3g/8pZTkGSgmSt0dNTx0XvM/hbfZ3HygoNmg8xC/DtfqPdwfy+oI6Bm0s
elnOoSYtK9oqic9v6yMmYEY3y2NSN4rHabPOcTVLLatC1yPk6j4u2JtqIu/Qh4jk
d4v6hz9wGd2kvIV3wtmja5QpQlfddZ9Zt+YvFXWakisU9nkZUA43eD+IVc/M1XXk
FLO4ftNb087jSB78l2eYkFPQl8IcRX4Lp5Cck5CA22x9VConqn301TnIXrRJn8FR
86BNrVgKSM7SQcUymTafDg52IVGJ+0W6OeyabNnc4+UBw9ZlJIXPZIklHT2CH7gQ
xMQz6IJkVTnIvZt8a8L8FaM/uQy2gEZRDNql8yOiEclyGQY4mnmHDgyS+EWElaSU
pLaI8crMnC70K2sl8EWDiPAT8/W8tk7nhr3SZs4k3T3LiNxAoPCa5u0r1NJvD8Vd
2AkkwSGc46knLYTrRNCFSdhaNtDG/L+FRAZHRC6I24lQvBZV+kiB00kXYdGh9NzT
Ijvh2VftbPlz2ZCUfYMcTnY/TJpDtmOXt/LYWFhAbzswMYpBZ5ZT+axpxXPF73Gy
8UNbAgbkIUP5yR152Dh4muMnbHCGet3Il9D6iEArjFWXJXdwBZb0XQdJ1KFl1ZkM
rfSKg0BxMahRfm6kkV2dLGYWPRG9wrgt+SGO6XqJCAY/h95ZpJh0m5PB17N0T0c7
+z1agOA9o1q8+YXyK48h7Ds0xoWgLnE39f1v17q4wUtBEYk7WVKOHKuqmnHI29oj
7m4yymGNCb16zU2ICUJWLjqr8HPOYTz8y9qFpvYO9PR4LGMkNm1HVZbfLhxTvthE
w4dBgbQKcc3HfR2T4aCiXkWdgv3BuTnzf8qPatx3sLWnQfnkLwn1wV2CR7I8HZos
nsYQZPwO6CXFRo/wqZyOe9TzopGoz1kZPI9gwAI++IHkDBzSDHGwJJIQ1bDPiK0O
Zyrr/L72Zy58V6j1w0gHnoBsOYilqqQaRdGrnZMMikXBylFbzSJ/DYnJ18Um2GeU
1JxPGqLqd/yVEvjqYYzGxeDGYi3SgUtfBXE+xnXf0n1LPExHkWGQR1ToU6TxOlG0
ciPSCqPAZyTxjxmsk/V7D2EN7eK1S24Ca0lA0v/NxDgFiUko3fMXEXzm/Tr59WTa
eiibwOi93/kPQUy73itfO8mH57NRJHLRsSUT1oeFyJUYgTgshsPxFL/CKuQnrg9q
iV2rDESR4wv2Jrw94hZbkgOkOyIj8K+e3CWAn9dD/T4Cj4Te+ayg7T0lnUYRgLQZ
PjOKwQXoctDsx+Hxq753GRQ9GGEiZmaufQzEXQ1U9kHRv+oxspk988OJ/Gh8mg3b
Un65I5T4o0cP+Oc8E00El9Jn4HDveY4+ndioMQNQ0c+VbCAG6LkVdu3XtBHDIDAW
QRiHtUAdFP9TtdRI3+E2wHfFpiLyH0Brc9aXlRv9Ng5gY/lAJE9iEZUdDLL5PF+l
9R8JFBqSbrn/5DoJlgUfPzE7KOTD/QACAHBpNWmfC6v8yWNFW/RFpcWJOBaLehja
1HZvpr7Ki1kqbaM8PzU8Setzcm5nh+bGh1Tt81ZQRS57dxYzQdvDusnMcp/V3yGq
ojbmEazjvApT8IgL8GsXxjckzm6uTp7uMfXsFbxu4eHm8GMGY1CAeZ6bqUsFIhdF
XEmn1uC/8XR/iMN8u3mmSb5UB74kWD4Hm9rm1PJU4M70zABaSEgv1gu7KF3SKs5G
pvDlXilrYlXGbmH6ECttpDIV/5tt/tL/QpwF6JdC3tO0idjKxSg2zYBvIB3rgqLy
HT61zvpwnEAwLIJHOpEp4dGBma8G81vNrtfkwTzdD/a0PSlrMFg/0ZHVXOiUgIid
1NA7Mgz1UWZwQdsfzUO7YUgCwTnBg2UBgqEjXXLX0GP7ju2/9mnnZ5lcAfV1cqPT
RPJunxcgui1CNJVuNQ5Yj4XxuAb7UzUxpU5pWBbarQuDyFBQoo3rAoUVKOfLwafY
sQz/cASgZ3SSrDAlyucPpZgGCLHuevmjKRTWgBhOSbQlCZ87AH9ZrskpDch7XI+2
g4gjIYX7KrQGqQhwixH6piWeJUA2OB4C1t69bc30D/PM0l5mAj9giEF+CFvVaIuo
XUReNrn96iMswZV9p5JEJdzzY+RdaKvQSgKh5oEl1v4oA9cJPLquhhnm5zxNgejZ
t53d0lma3GQiceG6KoAq0Yd6ni9wxGtxNFg6v6COopFJKELofmii+EW1uITvUwpT
awiDk8dZ/T1RwQ2WOQP5CZzBlQQOSdSaBKoS+VpD5BV7WUQ5bR/SpEdXqAq5WlSw
VMTkEfpnUw0QpVPmRb2NApStMnUyEr4Pv45GwrqWMlqF6KWT8+d5GwDIn70/ii30
749cBnNbvzAhiQM0GbxSQ0p+ShmQQoEGOytcuhQqDMJ/shRDSPNsRU+IvN4L9ql2
Fytv5IQjfhl/QXA4re/QfWTWjZMWxZOoK5O7cCREk2hxlAXAfDWINIbZ8IakPOmG
StMREq0ug98VoS18oBxe5uq1o4QQexaOxG2pFEC3nmcJ5AL8hbdFQ8SM6K9k0gW2
EYKyxgV0dfQNaH1K4o818O24d3Nm9MJddh+5fBwwqTLmdm9KouoP9PD9pUZcs1IH
FCybireK/03HckXWDJUVN6gD7O8Z1ua/B7A1b+iSYvdfhQu9UW9DSNtjnUUhvNCq
zumALSUEIP4ON8wXHnouuKfFrGI17F5UYntcz+xJON642ZQj29+IMcSCHvJGKk9A
MGKPwFi79zViXuvQUti9W0Ig157yTk+SgcFVk1k7weh/fnfOfQUFuvpncWK//Odd
wevbOjvxNlFXb7N4KbYc0YWxcthpfB34sYmhQH5EU5UVcH3GrKRXvJm6CwEczZAN
sTJlvv9fxUqdX+c5HWcsL1d06CZ7iAfdZSkY3G91rVbTx2HENMMbyVkw5Cbi0zD/
me7RcRyxAcT7HnDlqUofQysZs4uy2IxljYPk7Q82PFAl1b9vs6EHKgZkFHTmx2xn
6rynQUPUpE+sTH6RXQla6KTeqM5Guq1dTP0gzSZuA43XKwYSwKjNlkjjdRxZBEeT
G6SGEfHNAeHhdZyKXb9NseuUh09ilRaibWwpIx6kUwO/BlXmvdj582XaPl6xfASF
+0JlffPGSsyI4BdwAFB6ysDFXqdUtVNiEdPyBZAVb3nYm7ZheSJwrKDXjlVD4/Yi
i4XqMBJ2hx7U77PCNnEI+emdR6PqD8Mpj1h6MsvLJJc7/F4SknLcLg3Zpf1WoO/T
fmjBMhcMiDFauXOJBY3rSiGzQoWJ630/w8kzdryW2B/6gSTh3DBmzC1o/0KSu0vM
DAWmVgKZfVWOORNWvO0/bOYba76kj5Qw2pI4iqOnY/SJUjmdLFWma4upzvpOCxtL
FfZQOnl4ncZhIwZw7FXpf31GQoibD0gYTI3w2/BGTQLLmw84xFn8Whtnv6CND6EA
x4lI270z2GMCSAzgYPINMnysbM6CWyLFZUNTLb98lTRb5j0kMxfr4Y0Vbj91VUMM
gDPWs9DZJYn/RrkkDmjr/VGWYNJJM3Nk8hNtlfkMYs8ssfqS1aMiNQUnl7VL0uRK
ROyQUrpUCAHVilZsfg1MpyVANKmQrGeywmeokO0dicHXXplC7E8YClzZQEbycdbH
buaDH8xd0rfFKUIabNvo/5FT3qk7xJVpFHN74yVSAdz5x7rFS7G1bBXkVbUpIFEV
QWUkFfds9sob2KYzeoHAJR5v047UsNBPb0X7Gejlw2Dq/S62wYzLyWymfhOHofN8
Z8SF/f71+5bpG1JYrWk/IkSlJveup2OTDj4tEboDhCBnjx3vWLb0SHyTAJo4bjul
HLC1XNxU8l8KbTYs8vMXOOYFcVCvrnkkAAPHf2ffUub4yatrST0deaYg0eBTMyee
kCY6UUQu4r00v8R4EK1cqfiIsd3Qi7sRzh0j+Ky3OtWBJYnaaQyKX7U+9dtcjYfi
hV9TVl08o5GbQzpAIcxthqHx3ovnsmQ5+MWujDg5J/rYODu5m5VYa2BS4aU2McAm
ob86glNO0gzoq4tOpC/fpLD3knXaxKVBxdMMXe3CYrpk9NihIIfQ+ULjvhvMj8I5
lgLxmis/JqisUz8eD5B2vQ2l9daDjKpWo8sVBseK1jteBOqi2/TV4Cl2n3BeSE8i
a60TMZLdvFyiIdgM9ypor4JRctmuUWBIRA+TC+EjiiedMn7ZgjELoZsiqYOHbdi3
j+Cs2acFOkEd2DzUjKwnTL1jywb1DRHRZacCBjHDwkYVUAoPmOy1tEzGrPGJwkMu
OLsUHFdd/6Hgy5XHyV80q0ZczwhptNAyfKhlLezpGd2O8MPzq0MLl1rmoYLCYoFI
B+hmpVBsI0NcRzI0KQzwgfAN8ht0qoeZ5QkxaE9VQKjeatT5csCJk6P3j9FIj17o
MBniTFAoHrRmBuDxkhvbGaIGifl5L3pxhtG52iIlUmBkJLRm7hQV8Hq119rNLMaj
N3nYhjuin6vedhuFcHX9dKqZ6+7lNGqgX6j7BEUOzYML5qz2+P9HzxGJ3UllgzR2
xqKDkju1SdJ6vzg085hvVJdmh3FhpO6oz5T1aTK8j8mt9pzXMsmieM+pS8BOa0c+
FC6PJAobu5PEaB6eQLKYTJAUaEDqeZLwtrtWobURkiIwwBY8vyP14X8oCNjwVxpS
wOA4wXjCVGYDt088VOBTKk2VSNEqHKNpj2GiPf9RG9jbblLVJVTzRWfvUeb9IQli
K0bgcexux4RR/D8LqcmSK54qOH4/hfNxWuIQvgNinHXQrQYm0//+DI6nzpVifERO
/t5nYTzL8JCCsNbI2lGG6Z62Zs2sRGu1JLh+JwW9Lu72o3BQFuayNc66+T4fU+jE
2757fYqOJGzZeaf3+M7M8pAZCJy5KzkKkA3Zso1fEqFot0g4iEjcCbDtvZzR8Q9F
aTcB3yQYpYGDZrJqu+LjlDq63w4bSOt3IwE8zkfqvkEz0Bgk74u0EGhBxog78vUL
51pLKAmFzrafbmuw7OkMDl68n1eV1n38rQMFXSfC6IhgKuOCy1bmqZVIW8P5z0/7
YrgJ0wXjNGbiEkXJ5dMJ7qvoVBCUFJfwF8D4iu/4H5/4zQE5RZ2Bst+7WybqsrAv
Um/DvPVr2WY8flpGK+tPhGAEQdcXiQYUSXO/DzoPx9dKDbYSPfJPPImjoixnHqqs
g7K5y/MgbP2Nw00/pcQaQ1Un/ranuy58j/aAsd0oj8LfFA8+GchYGzei2Gqrqq68
N5TKfBdcy9dpaqsmegsdLOxm2RfgiOL8xngZFbVDgoYxeLMbWq9WgQu9V4Mw4kyp
iDEubvoDWxwalqs45CS5dZHseFrvTJijpprPeUif+Z/pIB5FkLis3GzneGJUodZ2
HhPNPmbC9uoYMYnV0wF+LtJw3p2EnGYL8zfmsf0cv4EMb4xjUDYtUo0okGPT4NKv
JCnsqXrAbHxS2Wo/LvozDNlHqJxVaifbqt3h40xDrNLDTPHzSrmscYEfyEu4FL7N
WeQ/0B5X6AW+HcQrzJNBpj76q+zqoOTxWJZha6kXPjxERVkBtnfxzKJCd4zhbqI+
FciYJMp7lfARWTfYWqyWxgk77q8T7bUAG4ojR0WrdJPT3cD6N6I2O9dkzcxjGCMw
c9DCVKm+UfMi9jqS0Ax6yM/fEmWt7KuT0KgG9SLjAXB0lAmUeoMXD8BdFbjCv+xR
o3MYKRXvys9gkvSQaTCBk4tVnWgnCqi+OIfy9QkmCuEiX5+v0vGbukM7lQ6Kv5mH
T7z+cSsDwvRDp2dNiz9sSf+PRrsjbGIwFNERbV5xiWPrp5mMpOCDepAGjH4abkuZ
9c/I6i0kbW1spGsohoWtAt42PtonnN69mRV96bmSUWDb49UpNxZ6H0gjI7Rl5A76
PDJnho5j0JYzvXMaxuKyGTgAh5pEXLsDiWy2+vqoSyjXPS1/PKD0YP2Gb3CpCp6J
vZVHScGCAeWGCQexixAKhZ7hIawxWitEQ+RltVji1KVR83sr7ufvjbNx9rYeBobo
KyuWps7emXABjCw+0BKsU7tPSvjDJHFY7p+BuQ0/a4/f2OTRqRZp+KPlemlJzk+6
ECupQeqf8AaBUr2p0rQEmNlgYJE5E51pG/mniUZGtR2PczcJ46ibZgXJB6Htii1Z
wE5hYmYsuT6OGbQQGLLH1xWwVq+gFqTFR8/52zXjSrvGLV/5GNzInfI7it505wGa
hcsvlcsK16W/0ARJnNEFsDvazqdoRef+l/sAwtcHCtLOqXQuPOGzqdQ7HKjsd7Qk
fzPO0S19xbw0MNMOMT4iyb/UWoAyftVsjiT3rphyZ11+gXsz4T4A7qURi0HJyrWg
K7E2T8KUsN55Xswb7kcPCf7un2QUqvcZgCmfOobVVsbMrC034eZdC/+RV2vBX8Qv
wyWzxsN1ooFiSK7AIAIb4Mflb1E12Ora0cNNi1oosUdb8Gf5ipeJZLN2DLyN2awe
HRv/LvFW6cwoJxJkYKKFNHAmnf8qC78xIeFyN1D8ER9lvxC3yLFOs3AbWmO1rCT1
0+yaEvy372ND07H63ZdbFdFtf1e1xaDPD6Sy/2UjKuymwlJ4xeNWAdxd1w11yoyO
HCxPq2oYAxiKDCGX4mAJPKerd/gRn/rjN7stJ6fSBeIuESHmS3lxKFribpHtFC5W
Z5Ha0ILMjE++q4E7M8adShLjURlr0qi1Bspf33RziFOq6vlTEISsNFgbsm8+tSj5
dBUaAwC7+SgifgTMqMiV0wSRiGHny0LbWQiW3nJUz8x7eigT0FrSBq+yLuIj9AwG
s6ijaDj3a+uj0bc8n9yE3OJaPK8LVOngwWerfP1RXcpx3ewNGX5pEWn3/jPjGkig
UOa6w7tOeOdRT3aTjnecizVc2LqbOCV/5wInvOdKws2jvZ7U45FOiuEwHoVBhZAA
AHoeBqIXQB/Ml02JfIWUdeU8UUx7X4loRIYV0kx97kAdJw3IQPR7fVZNmrILLkss
NW8d/ZiWLyidN0Q/luTjhkaff+HoQQbDu/a/DPC+DhjfBZM9zJ5Sm/1vkAy8ciEE
VOS64J5SvNfvdOLjwtauYpetXLmR+3H1IT05B7aS1K7yoykgVgwa7A8JzZcyqbri
ejdtQLxtX3TvAaVe6u1EVkq6CbANPg90dCDHvbDDm64Bu77ST+ny7elaen0amvn9
Z202yyh/yw7Rwdz82Rg/uY7MrC5GxPuffaW7gLHdD9fMKlTKtWw0WPubicuNVdIT
yvn/iczuvg2cjAlZZ3ZnltC98F5AGqiyJMqFBP+75wnWEM/68ZeA1yW81zwe3z/2
Hvi1FVBgTuEIMIN9M48721aWW09SWwFGybDolH7k41EkS/6m97sM2Wn7BNmG1/h8
trRSRZdJYq3jsvCdHY9ZZS+U4RM/7GCkbz/NWtgaQ6xxccGljqBuyrr0Max5YmN6
7Q8mngXCS8tcy3TgaOamLStJk2P3wcni10DWnRKQdBocq52MkzbNxvFxEeWZHA3S
iztGQ80r/koAoZz99B+D6q+mihuXLHoXiwYOwye6Zn6P6l6FbMjBgj0VlDKmVsJf
IeQbuR+T1WwP/nqtzzlqRf8lbBgfkcglfl5tnN10w3PK6lQDhiD+Rj28aKbfvDJT
bdPfPwst5zKiZ6y3fc5PgmBpEZdQAsgdPXj1eVhsr/Cy3pQtiiJCXyCVPvF7DAQh
O+ivoT9uMWI4livutNO10XxvyamCL9fv+YMcZLJS9iLB4wWLsnVN+/tE4mRZ+xmf
zy+XpK3jdWs8okMy+boSEUJ2BGVSTxJPyzHRrqBRdL+o5EbW8d7jkSxDDyisOXj/
INq4M1XwzE0m5QlF8nTyDY69QqR9tg2SawxLyDYeyyWmboJnqj+4y5R3S9h4G31l
hJA07sCtkQnsqtmRrHoBB70/9AjwlLKT9XbPWUt4EI3OmAA5ZD+9Lag3Cll1JC+E
dMjLLfsYeqihZzQI2AvnmURcwEIxazp+ZvA4PRWqaIu+nm8WxY5/wPJIlMM2+oAj
iNlNfKxge7gfBr4ui/58qo/ULovdW3MD1IExERjJ9hb9nwH/bLdRPbUlIxETxfrD
R0uM1O76rDYRlJUpDzf4V5J0p+3fibg6QItHyhFNQ+qsbfpyI7z1EqT5s5B2w906
jKzxHjLenAuGxRbBnS3pdo1IAxl5f22C6gJ5VP4m/pRzNWaY3FHSeI5AhnUcnGWg
CHTBQJOmqBckAUYVTNh1ybLhE173WEhH2ggI7TYeaBQ8I3CWcaklecKX3otIhhYe
t/FfTllRYgT4GbwKNlr+y//0gOuagFe+N0Pt7LP+zuCWUu/Tj4Se3+GtZscMpcLU
3n2BP6wb0Os+yh60+MY19dOrUls4AyeOreDyynX3wTC4zf/AYe1oGzxEPf/7DN+5
+0hjrQABrvj/t7ViiSb9ZGiNdKU4vcdfpPbaTB7zjEorsRv7W9mfyPEbp1rxYrzG
OLxgR/oze1pe8/MAO+X10yXC+fDrl7nwldoA4VJTk3WEpvd65OZ+GoNKZOZ03ZWx
Tu7x73/6OShPFEVo4Kz0Cs5IESfoza/Hl5DQnDG6tU0/IQPvqmS5FKM1qPUzg6l5
0Zra+NEiuOkfh9mM4C3Zsl0r6/SyDEA9pSy5acj9czMSjDHvu5v0spAHx+rw8D67
3LirL1qsEgXyQSFOMC3bRvaKYeAwwKJDB5bagKjL0VT1kzg71oCUsTjVzhEaM9af
3mI+QqzxVWwczrge9gEnva89S9S3rDwHttZ0gZE7mNqJRZQXnI0pXa4Rziq3Z4pF
ObKSAadZVsnhU98NsevKmMXdWI9K+9aM0VJ7T42MfYh29bxFb037iGt8dsL3wEBh
JX6XXL1FcxrEsQ/uR3CZ+Zdbkdb6VsINcj8/m2KrphKLlaQTldlWk2YLkfcTwTGu
NXkBpUX6uDYzHjTOkF9rrERZzGIDww37KeEtSvhTV4mqpO7+KrRFHpjULpZmnAu4
Gb+ziu3IYmgp/U7so+oiLejquWudCWEivCWJQUlQYzR4oIKc+nOgp3NDIYn3k2nS
RiOkTxEmWFK87sxqngeaKDxZ214Man17kqiolA06GRJHqlzcQFrPuwCh5/yBdGL4
L/lEv54wW1cK7D8iJgqDXoL2xTctMTj1E7VaoQLxruNtjdbxPtHPSsOswHL5s9ce
YeQrzsB2F8uRdY6yPSpD2dFFk62jTD2cqcxkOGI750ssWwdzN5rlYiZ2YcEcViY8
ECrUE9QgLcOmWESUckN52ozBXLLCJm0oTcLXbrMuVyywlbDFflVdWiwQcqKu3Z5d
MLL4Cpk5IfO/LaBI4Odg/4YU0SHqj0r3jHfVgeL6gF3VoJxanfBbg/ivHs8Lukai
UixEv58M1Rl1cKVVBiy6v7yCwxiZtiIlC3cwUJLxlMsWADXQUqnXSiPj0+Z3QjWZ
wWlzTUjMQuZcxGusE3OJ5Pt0/Qzpkp5GKfZv3QwzB6PDzFWZckI214Y7gJ+VuvTW
AYbqaWXinyCWz2ARokrC7oLlwS3qJz+x1f7OEGBjCkG/SvhTpRvNzdDXL5JqP1B7
vDZYTXcfTN2SDTymgH9S+QAJB1MJMKkMgZWZ5C299B4UcEPyjUI/GL5lbQJl/+bd
vNgdwWSGyqSg/ljpkPfaVdksjf5XHVDKUD+c3YQwcKOQZkZhdl23HOSkAOQkxVIC
MmO0IgyHxu/qkbp2ZfBL9ZDMx8tW/Yi6Fg2ZbYfdT+gITBTZXCjSZjKnYTN8IGlR
+mHkLx6uSbqRwWPkpahaobqiY3+G0oL6ljBzsvuGh7/Gil9Nchd/NY/VYR6o9a5u
ocZiU7JLulU+G24i+jxqlRvcBm9mIXtfPsM1BL0O6QZXL2QEzJ5fUBM9iV/eLX92
mn4daVbHknb8bGwkCWn1Ps4j9yakN5LTEYQPSMIzLBhkcanlKCT+/YMnn7TKLR7s
CT8PIxxfRneBMKvyI7HDsi7EcxvhR2efy32ojxZJ+qDFlYZeHiCRqrdc2UZRuv9Q
aDgNDuZ8G9QLvLZIuMdMeJz/jo97zdvuXf+S2JU1Xe9wqUimmq0ByP+1OsgAGJta
nM0gbuy3nx2zxzaYygOM4qROuZZOAlYQzeSba3echv+zzNktEt2zuNbC4uadzGHi
k/+q3GJk4ZHhsH2gSLfD1pK3Det0HI1g9mOgRACHUKC8CVJ0d81/UrGWP/BVyIkB
RLTS/ltLJQpQkXugaa+uLvJ7byVTrvbUMJ6n1PjJXye8fFZzRaku0TkQXMFKSMp9
oDE0pF36tyY/Qx+WWvy7rAEOfLlLt4i+1njWKbRkKxYyDZZ0j3ZjHbj5C2ejNg2N
Sh2cAbXFQwduRJF5XxJjMex4kegEwHD/mK+JM3YRjkatdagdQdAMlSFMhmBVnNfJ
5ebOa80bq1SZGlbHBDhCg1cKgr5HBR0VqK5lCmToD/mYN41yFeGrzOLd0N/lnw1f
s4opJGC5cTEO+NyfbU1eG4obbjKqlJY++KqKyC5+UQ1WrvDQpNzK8FqGn+9MyOLb
PbAfdh9XloWRUmBx4XeD0vnBizfVVIgWdeJJMfV3BBqjqWVT/yDVEFWtgL6Wnn9I
xcdEKnmjaFbHvu7zRYv2vPZTzJKLks+KiTJlTVMHEpCJ46f6zZ5Sm+oCBDaSPDMq
wEBYInAZe4leNJZVpAXHlt5/UJ0UrKXp7I1vLON6T4/JJYU3aH+E2II/TDcvrW2H
clbkyoQERRdEB3x6b/R0InCDPZqtERrr+I3GesZWJEsY4hZinCYmgWXDX4oTPCD7
WeCMCgptPrRSOpnRbNYULrnfFKSk3rPCNTQQctz5rwK9a+BB+WE9/JQYyB8VVcAF
iFm30yEn572SkjDuVyHe4LHDnuxuciqZvDCj8KMKPNTcdol6JjQYQrUAX8dLJ8Uh
K8iBCF7cCREie5KrHsFNT3IAMjgBH8CVjW+ftZMwlii2fnJP9G0osdqj21G2Mt53
PbegHHJynHOIz4hPuuEN7k1uA4GE25/3KeWHiXBTFiS7pzxCvK9PyV0u227Wz8y6
83tJoNeJkcXkI7jXAFNRJ8//3uy2EoIFl13dZUD3DJ8ktk3ynOxY79FHlH8GpOEP
gqQA4bp9kQR+H58cMJBPChJMAcVRqD91WBOdARvWlhQZH9ROgP7+uHV10ZwBNgP1
xLAKz5X08Ke0cmnujrJcOqfO3r8PCjoxvUdzmAUnnPU46XgCgYqY3uH1rS9VEDOx
TXqrBpM7fDWXqfnyw/KvfHXrAiw8c1knRA1NW5qgGtxQwGoy+c5ew6YZhfExYqq0
u8EuG/oSTszVniypOMxiqAjGnI/DzJJzCpoRhduGlGytHl4SNnbIIlGrvpU76b0s
FTE8orwiawTUVM/CpI8lwKTBazBfcm8vLuKOTP5LFvNtensleP3gnTiY1+p2o3kJ
ccE8jI+6WYtwQOMm20GT/1ggAuYOyEdCzPiapJZ3ONYykM2C6lddh0YOn7BXYlkR
/8JOL84JbVJAlmEhHTyE1YDnKmxq+Tn4OcKu1GeM3Cyj1mMf9z7JzHs3l1sGMa6u
+hOzAQeVg0Ryf6+YIVUtFmtnDB+nyU9yUciGoD/moJf66PJwLaLer3s2/2bRRoLH
3IDYgIen5V7mTX1KOhhXB2ph+2TZnINWe54gEZC6t6+vlgJnxYFc3bd7uTiyVRry
fsezBC+fZ+/9iLtYreDle8SfqcXwTZWzSjlyw+x5FafwIo13Ip4X/wz65WXEwHM9
aB0xBu8cO8vUP1r7HQxQ7SAvbX0BSLVBQmdNuuxHISKvIMesBd+pytfF6WqiE1HJ
bzG/fjB2Eu12PkPWFrIBRSUjl5RPc8GTipTR6HDQzcVa7Fx7hoR2rdnQeqgaUIRx
KCKe3igNvjAYkruj4+6e6+RwhIf+H9XN9Hm4wlPC183ExCjbRE2ScblQ0nK6k0eN
ZIcL4cjo/2WwlG8E7riNJMK75Z+IgTUiorM8DeMRTRVRsO0Wre97pVLI3L+Z1EZW
G1poea3x5s1m3yi65AXGKT4SLdU2mF4/qc6djqeC5jfkB/As6TKO9Tv1vaVpR9L7
4KSgZlD1Hp42Nya3gFjioWMp+/i2ki+UbQP5uyQOLyPAh3uCJr24BCMbvuXNUDuc
dSlRS1L0XM7bVnMMgmEx7z6g7KW4LXjH0Jb/jdvgl/2UGwUZhmhXGJH3dxcpNekP
DSx8Oxrq641+LiV/VLlyDeJ/l0SI18oIz9Hml2mRfsSUyzwzAlgn/QonfPxiVBud
V5TayttlSjb5NkFJKY34TWGYfJkH1C7Vo04fZIKodJ73V/7la0dNfopehZgMh51w
dfLy+ipRPKYQGpkffkIpJEHI93JMepOEHsPAQ/y1J2LZ0mOKgavkI9xpN/HCkWK7
Zm9OqWcpUUA1RkaohFboRjfCuDGphClpgJ5Iosamt2kGmnWmnXAzoHc1q8S54Ar0
Jf8rDZz/JHFWg/AKzkUYMQxyqZqvi0IL+JVc9p+Y8B72LZLcolucnzD+oTVXWtQZ
AFxpWqjvqz9cLvc4ygA8HhNjrTxKAMSwtESlQKtfjj5HIdOwBQUBu8CcVRAsXeRI
3NO3A9wThchdqISjkhrMXzQzYha9QT+JfxOmCtD1v2nNJqUfvnVENZZ6ZbmriwkX
1kz9OjPwwXDcIZ3pCtUsMQY64M/y19Xkn/CqripNgXi3HsaCbdRw9GYC2vU4pe5H
MO4hvbU72clF9ObHOV57N5QM70YHHgXTjThQmkjf1vXL/lTsB1OSMvse5t2V0UM4
/Yjg2gb93X55lCQG/ak4spoG4NoHuNpfdUU1T/FtvGx6pG7uFSFNOhewRABswtBS
mDy77DzGgYbCLZWsGTZLnSFt70K1p9VeXfajS0VpTGZQaj4BhRCl4L4IvuvjVbyU
ww7zfVkw5WjMU9I8d1WwrRtyuMZWDGVWORsarL4cZNSIhaL+D1dC0zFSPwCD4k0g
vQK0w2zTayh0tkDVBvg4MG5CDIYyfDUqT01EtakNhSawvoW1xQCGNhEIbQmYqZG/
NhAPlTkrvlrdI9IwFwqQ5mNLt+eLtLFbHD5U/tfuujmFj2fCccRFUYU8ecrPxFmK
MS9qO32iMpvr8OZqxPWCUMzU78PIfIGggSMxT53dClP8sZNx3DgBOieW1PTUybsp
KNqyR8Vrrqt/xHlHXhlm1WDX/5ew6Z56h1kBMu7seZNY2S2AvFffRYRAdxJThE0i
3yYRitLivATt1b7X842w0nlmelKUFcIrGLhVhSR74J23oojx84Ij2d5HjUQ6xrL5
GMwCMrMoayzh8Hw/qkeitNPXf5rZKU+IZhB1us08mLKnRaPshiVoP6Lbv6adVkSH
wQYLajmh9JI8uvgPRWhsdnGA/xMkf3PnV6jxvvdkXsdxLlRrOBZyDm0f2v7aPfjm
DE6mgL+ItPvGh7fk14z9IyuVSnoh2lA+XCiQ06jKcC7i4w8hWqmSoKKx+5Jg4zRx
CPZ5NskEPe1XAVDtuA6691wZz0wo5OobLVP6mNd3lVj7VbL73h9owKdkUAmasd6N
yLI57UeuJQNKeEOtOIe3MyUidqLBP8SVxtGMnKLTul0p2KKUKHpzLcN7VXaFGWAh
d1pZAXByEfPiL080wDOnModpj+o2Rf4fGp9RpQTVn9SsF6cPq3/wEjqQn1mAA06v
Md19jfFauxpVvk37M8AA5Lane3d/Qcs1cwHR15luD9qa0SxtgNgP7+YPw7CoR6uE
aUQbjtSaeW4vm/vY1qBxHRB2U9EwNIxLbUAyPhUHBQoNjBR7xMHPW4HGdbL691YC
bNd9dUGnmKLoHV4HR3nODzauIVHMlSAaJWb3sJDorKUwNVsVSN6qfMJ7pk6sbQ+Y
VSCPNr+a+GL2L3JBp2wW4K/Ll1nQ/evupyYiU4WhZX/nA6cmHYUzTdGk0eMXJkWt
8W5pI1O0NHkyEZoX60o+QxdhP2QXKFwu/lSupGTmZ0ZTXLJs7hwuFPO2a7ujS8wO
tzq2Za6ZDprxnwQc4Y16FsdTIwD1j6UACyCx9EqWoEN2XzsUm41OqxxaawhGne88
EY3VdTpOeO1CqtVicxdOl45ywMko+AqbX6NL9Pp1F5Gl61mAfYL7xcWpGIrzUklH
aMFHKShobm14A9JKkEoFw7KonYgw8DSUMgRUxi2iLO7MbcpBUcov0oBVG2gZsBSG
bTnDGlkaLTwFHKIZK9BEtAT2/D0TIv+qtR/55n3NWthyAfuYjQE0r0rd3gG04+3f
FInvJA9UTywaNWTAqnu0/NAKJnndUoNfAHgmpYkN8FNd8xjbi9Teu4suWPtCrI0w
Uv2kKuEBYpuZWO0A3/lAebVh9d7hGKZDlGbu6s+4J9voyaHRR37Wg9VSdT6+XMog
m14Xu7K7YIUQ3PV7IHLad28VCZpje6xvyQWEPcRQfWn3pOIn+4vd960tEJD+VgzH
utfIzRN0CpGMWRmE7dFquSy2z0yhMZRymJQeU16ami42hwqbm4sXru58gJ/LeByf
Fp095msHsqa95+V3a0Kq1JH/9lbb5mtHoQcikfv0oUCwXgSeroSk+8CfqcgKvqxE
z+6negt2f+AOuoxfbOXILfdh6DcwwDz+t4CfO0EmJrDQ0vWUSt3koFjrZJiivW5L
F3iz/MbFqFX/wrucQnRAFmsaIK44UEodDjNnNtldJJgmqFxHWjhNBBZ3QEwBpGr4
2FTTkP8vK8J4F5HagWSoOUcxDpukOIl8/8lYtchOWEWzk3uZRena4Mgx8InIrfAx
Dudl+8YrraqCu5u5sH8kREoFYof9apy5AoDnqSOtoDrhL6dyAC7xchPpyVHFd4ge
7uwMzsb42XlhRijpalZ9ubGgE5cgGoEjPpf2iMC83c4YxdUt3+LFAdIg7/7+vj+X
CKHp3628nVU0e+fNqB4IltHZ0n3JOry+MUKE2/uGxdXlltvvv6z8IK8jTEpxzibQ
NGAvD7NnqHgPcQPb8k7WM48F+XjzwVENGIFhmLwTSeOwcIjiVwpnwMvn9HiRECEt
+3QXMLdQ7TVFOHoU+ZmD9n1N9eMjYx5rMBb6QkijorTp9uSQjXP5clfRa6wy6VL5
qTgGTbF/wj+JfVpLQzD4hFmqdwY23IVFPcaxvahCTZo1roaOhPz16HTQFGt7F1tz
OTzQJIzmxFJzFdgNWekkuyR0ZCmOFAlXHTBwd6kJ8Ky3Cr4fw6DcTpmxuzxneZbT
fggyx/0tongngnaO7rjuInzMxpCtXP1fuW2cveIyuOvKyO9+2jPzLHRrI50m5tpf
6elbVK10+B1V5faoRytNNpnacp31yL38LSUdugNzRurTTzLSYRIB70/MInmfB5Db
/DxJQ4MyucpmI6qQzkS9xSzLfXdAHAlCtXjmyIuZLg19ICwiLAkBIkU4XJMPSz1b
TZfT34PslkTzat9ZhdfKp7qCVmYMUUfQEzzdoxg3KvEZg6X0fT49rOQAWpL6sNVY
QiPymCFWHAFAn0EhNyCyZxtIEc4SVn35mvHtpY4KMtfMOhnCQUh7DpCd6dhLiA08
sjCQcDzTq/xhpmE63q1hvLrqMqtD0ZIjeI9492W2x43zFS3OyAWwhVxZE3iqh02M
Q4u0nee0JDjtwmQ9v04lqPN6OzCn7tVkqICMarGOYnGgHiWUhTC1oG7lUZlibsFv
n+6Iiv66q4TDCOKIPiY+v2WTGA6b9vNshd1Izq2WFDWqrBtgI8gp3GOo36DzILja
oiIkX0kr63+3Admk0D1qayGoU8xx1tU1t4pev8LkMYEuE7szKHWPkKFxFx8j5H0n
lNj2kh5NSfxn6fWuvW6EWRoHw/8TaYtqZmLqP13UiraOEEXuf3S+sV1RbUxmm0Z6
jwefIJjNc6Nnebfmq+wYXU1FWzY/6MsMbaoq/bJRkzqHR71Y7RJ9Y/EGbMQ2ObXt
whVYNWaet/peubXw6RF85aCcML/waaHNeN6lF4m4Tm/ntgSaASGcwYgEPxrLOuWF
irbIWBfaM5IuhPFrA2oDKangMOD9YpFO93v9gctkn6euNGpTQZIW5F7/u+vP2596
6kKJC5yl6qCaAemQRq9TKMGeYXgRkTYAE1Xu0Fce3QX/zOZ/xypBZE4KeCsIBw0V
glM52kccnk9a6ZjYoZMHAu5/rnPIPMhdoSqHT0k8NVzZpDWtp/Fp6bc6cmSPaR8g
6+SjUpfE+W+B5kStZlfvc5Ub1IXNgkt1gFoOF5Hh92/GVY0l+9Mv2D2zh6C0OZWb
dkazcutO/xpNQbH3wc6zt5/EfVcWNNZZeqa/HaRF3QbOtIW7GtVIuVRpqjxL/WLM
O3VHXuGTTP6UiQ7I+rYBKpvmtjeOy0VlICIoEtYlu9mJAGzcMNBDiyUsec5cFZsG
fPVvmFvSd86vyvLKad6U27whMujFGgx/9NnyEfUNYBwDHLkwJKsQ+HuQG+tzMc/j
INpLM8a2pC82/iMBwmlNz+junQvBVx7QMcRxhx5vjZg7+3fCHBqxOsdVHa2wjQyo
qFs9IXlNTn8/8FKU1Wgx8mAa5c7n+LoxP3ilAcX699LFUT34NQlgab5Eask67ni2
DLWzKoMcbpZWqUaVAD71VxAEMORB9bwl/M0dtzwhi/bKv8n9dpA576NLSDu7BUzw
Vb/KTz0CAut4rbp7wUDdYPH7CJ1soj+0e/XbKNPKy5C8PMc1QFWAVyvDFd4fKYdr
oosJ4C7aAR0gIIFtF8b/Enm0dzoILwNPQwEY+J9Xnkb3lDGv8Ja4igzqHGhazXVT
jW4Trt5kyKZUXUcPVIf7EEdXMoXxVJcv3OlZjTfnxo77w6Zsf+kRRH2DojK/cK1a
/p9+smvNAO8jVqtR4485ocYwjDNCEDCaYzeebbYdXSra+okTjFVIrjLSO84NWcTH
nkRcSqwzUte7+9Z6NOXEm6LqYaoZPxCzT2qNkP9pwv8Mk991vhVNBv+zzsqh+7Lp
zxkhF02r/WwggNRIyppUbM0A1AW7Rbu2x1+Q9BeKTN1C4jshDieaqbmRoNKkIUx9
qxqtjzNFgYTuRf/nMk8JKXOLKM6MrBFQDxY1wMl974ukmjtKOtiT5cPJCHVWWO6Q
744QJhvlshkZ9ECgjIdulZoR8bGBcKokk4tVCpmI93Hr72LPfQAEHIplhkokM18v
BCHk5bSDix4rBLiRPu8dJ53chAhwk7v5wsgkDcD29Zy70wNL2mbXXm7RMR6EQcgN
gVaRNsahmgCbYv6IekZxHkUz7/xbfKetsKbPs9uYypoCSXi1mYZbi866myf4M0TO
+WEsH0A2rSb5dTVnJchzLe4tUGuxRCOqjpizLMDE/rF7aeEIqYy0raUJgK90i1bH
UbmnbL2aXwAk9hWLxWSkUYVFneAG4jNtuk16MGxtw3BYOoAGd3CDTWBR/FcLKcDT
JULJCeDR1l7P/TiZcplrufcaCZcrSA0TltqV4umi80Z/diRkyzbTWrhcnXXUAhki
eIXW+6pbaerg1xWtlr4Gb8b8CrtDRiiYB0YC6v8VMLsrJmMpobid+jvGCV85KDfz
NVPF5np/dyRc+1V3y13vBYbRc3ALzDM/tNxZVW1J7OXK1LDFycig4DoEdty/c9f7
YiMSk81VAz+vg+VnU4ftGCeLV3TKnLB9S+WeqFbbx6e7/g+NLb5kB2uM2P7Q0yD8
BgNFrGEVQlmmBQ7LFnn6iiVkgA5mPgIQ/hEIcoxhAFRl21CzTQHSpc5lOergWkUg
yRvqKbrFrkNe68T0HPLszTjS5M5oZrlGaoOVnKV0bxBiu5HNCoT37i9O036DSGce
5SGfdswdJWeTtuQng3AT1nmkoqeEdxd0V69CE6S/Pj4zHcfo8I/NorGL//vof7Hl
DnWQuLWvQ+o4ewIWeKUeS1I+LGfQNGJrMc5ibZYe9Sy8vCQDv3SiKyM9rsVxodZ5
/hvJbQ4ZFdb1OHlAvE3p2m/18jvB6JijQbKR3qDbY6YO2KgWm29t/5YniavCI/RS
TL38HrvrhYJVPn0+VmElWp0Tuou1gFcqHElV48a16Fo8i5xe9RZ7BHwq5SpPLehD
vrk710uKlu6SO9wsSoDB95u5ID215te38UoEfMzZxoV8S1K/L0goqM42gL8ywou4
pgjX7UcFLadm1o9jERCIDdBO83s/PckRoCD2YVkR6L7a8/T42BQctWAsqM/Sb14/
im0dm0uOiTFwYeXXy7e7Q6z8a+rbOAuRTfu3FBj0JdyRXgbcTwKX5nlXASkaFqST
gBMK+lnUAja2qzuKFpKpW9E+X2I+9FdYZFTEhM02ekJiFHezVrmUxW2bidMIso5F
UCxPfvVd7pQKFiqBm0AoBYLux3dDl0/CDP5w4H7t9MVELdPE17Bm638dYVQyqVgr
aAU3h/0h6kzdvJk5B46Cchct5JydyUoYA8d31bt4rJEuEVUt5Al5F4g96Pohex/K
z87+sHru14iVhxcdkgN2gzsAFHEBD8rIZJykVec9i9y/25T26vadK4WF/AhRjZY9
HxVUPhFJe+cV1IGWJ3nxmFkdcxbH/CQC1gVaHM6eSuRXmV/QlrcKLv2+SRR/1OcP
a3f8MnGQlUceZ9MllEa41kGHeb8PhsawIzgz9ELfLWdtYWfFxMDlpNOiiZsEQCG2
QBb9zkOmzEVF8g2XvIDmkI2KZX1Tg76+BqYR3QvcEiZnsX87trX9jl05zN2LWlNJ
H3Ob505k/owkuT0X3T3qz7WpkivGhdYJNNRoiT8FF2+ier2Kf6iHGn2R0+jJVlKl
PkQX8lCkCAK2TnNHyPGXOStdCEvb7QvEULCEvJMTNKmy0b6r+/Yx/ECBUYR7EVKW
7KFk/wWBRQa7qyb78mi2gydONrMB/7t40veNR+w8VUeshj+FzgJAxgAwqiD3qjlG
sshxCyFpej3CdKMip08Bz9caCoox8yRgT5JXCWsOq8KJldncIA+gQbMGG11mTos/
GN2Iak/3dq8dc1ZJP3oO+1lJpMNSIf+4WkIGI0ITh9cjfsaBtWvd+aft563eYPb7
B+hkezSHTKPb3BLEnvpM4c6veUnPK3HhmGS/F/KIYPgnwOZpLgBytPjYubo0PEFq
vsZIxYh6CDCSCKUBQhvNU+Zl2r2mY790nO4NGV5vceFQOZhXNLQKrQxR8wmaIRaQ
/ow6Yf+DnYyG87bIv9vE5YrI8Do36XiZ8WVTT3u++bHhcEuGfYJY8SST8nbjnOsX
FMZIQYo6Uav5ts3SQnYU1RdINASF76EWwfvoefKBWvuZcZN4OcMl6P4CEPJNFuHR
Otze0A4pWbvS3p0sBIH8AgWgo8l9UOzkhH7OeadfbdpZr2HtLNJyjVYmxatPI+ey
BfeZ7V+Hci3+Drahk3LzcHRjdoShcA+2WJygbwd8FvX1Pg9QNqh+VUhS+eexfCCI
ibtJHLeZbHdHwmtusQEWlGw8e2p/BCybMmBSz303KBZYgFR6e4Yhx8UCVXKcuMd0
bkUqhQXquv585WXImdSiS57shtV/YAy8jAfW9devgNYU1S3Inh+36t13mxfe71Zk
U/7tyOhYef3vm6OOeOMCjy7NYFMmAisgZRgB1eyTzgkZ9OH6io6h6sXtUJXTuW/9
gq6QOSCYbT4aHst46sPNuUYtDbQ35cvBFT3Ib8CHmacy649I0isH5tBtJqdieOWg
u4hqfabQ+nQYm85iH3EsWz9MA4/WR/WY6CKyq3BF/4oeGN3zTRtGxoe/AIUocIAh
xLo0gDKywiHy/f28dhqYcLrDuyHJ9Z4chlB8jfrJ0hdF2V+gF4hDGznXk82QFWz5
4wgydJYTtM4f4eB24augo9AJHucEGN3fVFP81iHOay056mS9gnp8qtTtpCGFVwd9
GoN3e3efjWnJIXT/IYnAxhfsOxF4N6t7j7aZj/8FtTs7IJ5Gap8qne63I8Zy4XXp
NaUxnuHaNTGc7+J0mat3eOKDpgv2ipVnwo0Sgj/M0sAIDg+Pwbs/ijdqVoZl2Uqf
aKo/nk3b43PzmJnzYXQGgjrB7X5z8bFhRC9zu8Or/H/Gtvp0v5/f/n+p+KFQJ6Ef
BvQ+kuUugOhIlRHLkjErcpOmTs84KZ4K5D0mtTkYMERkF39Q0khM2cd4tkwMe3Bp
0mfwzJ9PUqOerHUV/ejBjY/vfB409+JGXdtoYSHb+wFFSsEDzOAJ12lzahzjzThd
IDMpAso1PIG7gE8ccf9VkPX9ucOYd7ZAo4b+6YPzhVHId9J247GEspQM9vs3AFNV
JdOYzqrzYD5H51uWwa3veD1via08vpQQOA/IxGe1bX3gJapTVY/5IPEMecSRSmKP
6EmVDwfBOWVEUon9w5HnAcGQOcuj/1D1+fnlYyo/pDeoGnKvkyp4aGPeLklcmYsD
uB8ssj1eIWItk2Allc/7+9k7iqoVw8R0Hnr93I4rBolUO7tlqAFgBQjx/TIbjYAH
xWRZWDWk1kk+Xzjj7SeWfSe0ZC0RPpGRpqxj1Zi9dZgTXuHXTKVnfvO9O5JhC1H5
KIEVFFBpd5PXfwXhiAaxuBhnGCCC8t/SvMpc36dkjPhlkv5yWEyzRRxwNWM+QoXr
T9ovYIWSlqETYRoqhsB1nHK/3jfDqJoe3DR7qy60712CDmJY1YkPzowa5tYDPNz6
xxeovxPnm1g69QxbtLjBGIcTPU9iCiH+zvdK7ZAy3TXjluyPvB0LsQbF1pSCktlE
TxgboB6pX/XcmINj/dYlHOgSl6N56cjZns/ufY4Yg8x1wN7T3k7gt/CWPGjbbTrq
/zEftZOyRVBXSmcY2F/AOJtgDIsrniabePpGgw7nIIN3M4ZO+Zzj4/IecIhSGBTX
Jb2Lcyd01RBHow16BBvBeta/SHJ4N264qlGfgqHIbjC5+3xkD4DLiMyvneFbRYAU
4KQK7bCxYmVLTFGwSX90Uu/a9Io9hllbRn4S6oHwO9kStDx9E48ZLC5MhFVSoBGL
QB6iYUixjCuGvMSuU5/VBDE9rhXhLPKuksHnWoXZZy/y7u/GbT7lzuq3C3gCyu98
opSngP+AB8/U+LTIMzk/SOZXh1CRhjgskQaUL8jF9iWFZ9nf0yfKGs2Eway8bi96
dzpwABvZfKgypsttt7gM+gYGDGkJMnq4bGhwx1pyZ3aywBIdoKU7s4I4HITyPmNx
Mt/bhX8fx5NuEWHDTl4J5rIW/TsNlwS1Jw/P3YinFg6mEJa2HCKQ2AGN80p62bF3
Eh7XO+II1rvhN8LWbGFISMgPI3XDqHSBfPZa+xyPR8H6tIFxpbdlDYUIkUKz/upU
UPppy0kplzwDhqDFEKpEKps8FUaCcwNy++aQEZsXU36QHSMeks3q19FNo0iJS+j/
gZHdL5wcVf3Hmog3Z0Q1+EWHWWYPG/FLps6x12qpiLAM/63M2QqTb752VAmyl0Fk
/r50NDH79JeR3Zvq235hjdkigH1E+FWTKFWFUGkF41CA1GAMByPp4Fl/UfLUApvU
m9CqnPYn2FMBU9GozlQ33jJ8/hqaKC5PtZmS1YCA1UfFM7ZDjLI3g0OC0VsEw/g9
KZLm89MgBF/zTRR74JluDjeifhi6sbHus25XqMD3DZm6bQTIG3fDT0MxvNFWVPPE
mRFreIDxlxDKnbPWiFhOhx87rMc+2D9XXV+et8Jg+4p3h19VdPV05SM9wjwn/hN3
o8RztDQZe9vkZU9VdEza5/alkaMReOj+BA6VQJkcAArOqkQKQU7Whl8lbWegk6DP
Rnfnt2KTJhj/MZZdd5OTuSP6ooq+JWk3Ho33p37RtfR4LBhBTWNxkkl2FrviwltW
E0fc4fL0hG1sbFMhQMKIbHWIIuqBplAu+GzFcFuYgYCqLbmPLn2TajepxQpeNjBX
MReJ/jj/6X4BOfk/wWjieOck88sOvml4GVLiQCjWR/bAf04CLrwNtCAId5MCUDBJ
FVTg43Jg2IW8/nPjXyGqx8jRA9++fNmd/bwU7ugxlfJwQA7GfOOK4RGmW3Ga1iyh
DYMPoa51huJ0CqoHvKWOK9eMwgykvikpFNfV6oZBLJuMiKlVrejBZyQjhmRiy27b
nUCtMVajlCxrhqsGgslSuO/coDl1gwQfLOyr/pBhOIOCylBZQ4d7B23NkNdyEaFp
bBT0hrXewP+7gubfwOPwBotXb+cWjWD92d9hSzxt+HNI0pDN97/CyNydaJ/Q1rfe
OQKpySGXIuA8gkblKLnT3GqZmi/dj+1MTfB/ei/vf3/aIEJxr+imSAk793xiDMNc
UW/kb2K/Ulvbp0WNwlqLyZDU5FB9jaZSw9b/oxdNVq0mgq2ZsQ0WdiVIb03xzorg
v8k001ga15HesHMuXk4uc+rO94jatmOvfzX8bI+PDtJUNJmQ6Zw/7WelEIhA6KoS
LVGw2BDywMMuHs+Qy+VhyRuNupAqwFfCmrHXdQcW+RaiK+5aGdkbP9CNM+AfQAon
nUd5dPFEAXO1Z6/9GKb/uQG9rMtutt8+bqQMwp9C1c/vrizZrAzbOARMFBWHMLBJ
DJldde8dlzHU/2erW+uftg+n8KCj/8kujetIko+Mifrbzv4+HH1Bdmixa0zoNo0B
9Ohri1BNpy2RD0ivQuZ9QvhKxYnYbyXdMQVDEGZ9CM5PJ7TVXWq8xg+1tW97fKK9
uIYVWTH+RS+uJmEx5b2PY0C8uVdRSSIKzfn2U9oI6HmtOKAvlC8ah27AKnC+ZzzL
9MaioHNi4K7CVpqF4y4mbCA0lGM/5wnhu/RsdbY0U5FTAuomZp9JF0FQ32Tr3RLZ
wGhJ5qQRbCO8/L3OoLqH4eF1sR2LkuAkfwM3shrm/ThuDMMu7Fdrtf0OKcyT27IW
DapObua+gbCQsyiUIoMWc9mRwgXuJaPRxylqR3mJFl8WUVz66v/iw+vlj95ZX2cU
DWQGGFn2E/JG88KHANoTV8UH4r7kkkQsbv317jMPtjl5WpksNTYxfeTSkBg/7zZp
M6LahUQ8gtSffSnm9ZDHWI3IfqzWYgnxEMlwkGxCGwZIO50KySrI0g2lfRcU4Z01
KnrsOlbzEi7PEwxa6qjN6RpX5ZZ9z6EKH9L8B9Hcu6/n23PhzIvFWRiAk1TprWtk
dWW0JzhhkD0atHZwvjkHAzKIPyp9DOJd6yUr5ViWDXYomAztCRXWrDMrUp+1LcqE
NfrR6rBCkbvwtqNIY4aRfqG7Hy4pJ7EJVWkGh9EIVH5vV6BFmv4xvZno2eXsVOgZ
wjSxqeUi2XpCEnbyLT928uqM25ETMLefnBqzHnlwPrCShqtO4uT3zpiaThG8sP5H
pfWsfq3ZvfgnJHms5Bx3XRrMGoFHmxFLNf5wxOiSF+rEDdYiuf4E6ETvmRahbpS3
VzKii0iFRp4SDqWHffBqiH2szJ1AhO6icvf4Z1hJtBsX6jXwDCUwBTgMbTRe2KBJ
Xa051O7nPZJuqBCLEYE3ok2FUjDdGjy+OLWR3GN49yxbnLQ1+DEK4EkQQIsGZXsX
esgVT4Oygz3vAZ0McPWHYWBfG9Xls9ZmCzGpQAkSpmNGltbl3JCT4REGwVDDsdAm
P10MtxabDrXcVQlBEVrAj4r3ZErxnd3L0MAPfTNf0xwYLh0ZZV15u1GlOjcirwqC
/isA7aYLAVGMQIyAezFQqEsA/yU0HnYKLefLm0NOD50KKwwo/jeyVCcEM8qLz4lY
dxFTYuvFgfk8at3fw4OBpic947iSo4w1MbZJDYcPXc3xNDoQTtkrU85p1Lr98REP
/aWLpxtf2FG9kmlDGZB4jeECepkeFfuKf7eI2NVlEIuCPka8FhfSsxv/syrOPpFY
6aKiIxMK/LZyrZe55j8KXDBjbliP405ls7dGqZXpTzBPM4vR9GWRPV4AiJiZL0Tg
pRd5ZNk9AqEtNJcWuV8wLAAP0cR59cQPgb5fEPF2d1pfLOim9Wm/Fi+Wai/UaHkf
O+2GVcXmveaFDM5vKOExU3vD1sT+gGh330nGvpRCrDaHCVrn/hwokrtp7+A4VNl0
oZMBCw4/yHMmrHwu7Zr3Hod45tlI4gNXFtw/DxEmev/94+PBcT/EgfgE0qAJf36l
yjzBsUhq4FfsHZXNkjEUgwkPV7Vfb/TuwWOcq8lCocoQSDSb1YdPhvLEYwQ5OrNO
ubt7jV6fEr7cHwrBwl/LbsiuQ5zsY80DwuNRsPj3D2BJgMrPVrx+0jEYpCdiEl33
RgI3QwNkTH01vyzP2C6/K25IlTbYV5digT7QxZqssIsHqHH6E1GqsKs18iY2/mcs
0FlBFq6tkNWxNCJzwGTWvY3zqKTHbqTZY0k3XUFlvCRPQw8zxpBJkS/vLs0pL7Zb
c3lJl+Kw+zCgAKxnh4AJCbjJzJxyyQfS0t8olGjKLtHELNWeqd74QjuhT3iJYtzO
PsLCxYEyVpeRlCBbgziaICXM1Cb8aIeagAxixZ6KqyDgpR7tsjYmrgzzaFdesgGJ
g9Rgv1oHyRos4/VjbnBIYSHGRO/+pYGszcAd85K2Ap0EsGhi/1B7p0xwIZJIMb7C
VUmPM8GRtxarcgTRWsIIP9cGLbszzPYe1gSvTelYuPJC2wVw3kVZfmYsXl6my38X
KaECqyEvrqZbtszMTjSn4eg1dy51d8V7ecqKyouFEFtzvSaePvb4aVaDkoJ9YiAQ
ZCHGBCZS7dXdH3fe60XarQzBZkTg6DH6m4GFjUXKG7RJSvCiswybj5Fb1AB3IMbx
2k4G3dOpbLi39zEBtOky/sXdfspxpIxQyW3bDqTGcsIcjKY67kHO9pIKu3DM1VaP
prpQ2g6woXIt6ku//fQ/jv/eeyLiIT4C9/LnpHTgPjmu3nW8ycwzURjCiglPVyvt
FYfP9fGBeQGUHvMIX7atdaNlj7uFwp18yvLyGpGAc0S+rtDYxLCxaamPTfWfnDWR
P/ewVhrdoySYMkeoo4nJsnUJKSwlUhzf1wJ9DSRK8HwL7BmaeOiAM5HLJ+M28ZVh
18CZMMNi/U2bXk4SH8yyxSyb4oglIUF00yPXwh2KE7V2Ko5JENd+L0CcOCZe7smC
xPU+MJScQN+IPKRubE5CUO9Ycq1QQWhBty6ou7qTaE1oZONkS2n/GN1T2bUsKFaR
Byr/ODD7P0D8NBwmjNVhssfxXa7/QuMdSYkOBwNwfty/zrKSQADKRiTzTjAMwzzo
P/934zm4e6SfyxaaRCgx0+AnFa50xiEKWwsfBR608BVerJ9mgThqoL8wC7sg3bn0
iBV5u+CoM9g7U9sVm2PhZKP0deRmPjxlEfth7LzBOIHHd2igcOxuD666ZugzmtGv
RHy0evc/v6Waec+4y4mgfHDwXt1yaJ8x6S+YpDoCsTLnl0HcNHAPts27kjzCekYB
BHM0aZLD4U8E+cjD5dBbjFPtia14flsn5aFSN7BvDHXGPFPM4vjceT/BCM+pCZM8
TcAqKjKNulDQdJk302TlKp9rlT4xUTda+WWRHE9LT8T+VoAy4YmI5BLorBn+GlLT
4RrXWxlVeuFTzBWj5cUyw5gOSNwAHFZJNK2bvAQH52ReRNLXsSzYC4sS0kumDfX0
iEo1pJtSKeNIIGOvUHVmc4ud/I/sa1c2lQ2KB0yPZ9AKGP/ByC1o5Ix/YMJoXmnG
N/g4vDxSIrZGo2SQE50bp+WxK4IuHLbkPry6O55aXNW1uX93ml8hQd3HVQ/UtC7+
fEbejOeF2wBaivZ00KSRUd0q683+2tKq8hztdmTNEcacUxp2+vgEpWnoov2ocZ3R
t7ddkMivOYnMnqxFu7VG9i258WOoJ+rfL6EM/9oycmHNZkgGwLwXiRA0sRcRnueD
DNOUpfYhh26rbwHh1cuzBeJV2dUadH0oVVz//cTEsQ82igYKYhdhzZwNz90NdxJB
ywoouowhuKH/70/VVx4flMiVaYi5p4NjHUyD3vU0Ex6Pgv+yVOCQ0pOFl6dImfdy
+Ia/pjTPpBB7OlN44t8bYtovFVdCzMrbCxyg45nqjHfHTIvx0lW4U7H5TVzy62zm
JfQUzAXZIULQp7GC4mrY7KwfketCSnPVidlEilfaAWZUbvqriUv3YKwm2jDlxPXm
QUFr0dq+fYrrVOW4JeYUjKrCpNGPhqcBRnx0k99va7vbLDjmdeWuQYq03bDK0nxj
+nqeYlPT4I9nZ7vtcVb1e5RDeVWQA746nB95W5lf6JMS2tpsnXCcurSnncPDE500
vlaBVjgyZR0o+eNG5V3JiAmafr1kjI5s/1f0jDAomkuyB2J3zY/ExGOiUIarmUTW
DU6dz471DWHA66mIbj4pAGtMtfh54L0zalhBfiQNHRbJpDjio2e2+BPWPEr5c3Ow
EATYI90EpHiL0opTu+NaEMvghFrRVp3EhAJlN/vlWyTEXzzYA26U8qNmRnuGp6ir
+IyXlROadGsHXNoBTKFTwhMt550esbz/vr1RU0KEhqiHPhTbl6wwC0VSE9JSuXEW
PWm9oYeCrAXATfX6zlOpq+klIHiOamlp/ZZNM8a4v8ZF02/B38Q5lH3mh+rAbPk/
QeNWN+ZsrPmC3yyvwGRkogLLqidqdsNvZe9RxrpvXP/a+ITWapysjd/bvhGaTPAM
dXOaxA1i1b6b9kTK0pzFyk3t7fYL6CgbSZzu9fMtgF4V0YMR3rIePgl/cPFFA4D6
zmE7mS2RDB4OaTp9oItXQKuCBNG3nG2/h6Rt2tukPFZthfqdUEAL3EVcpfKbFlN2
Ufs+crToubh8HvUT9QFJIq6xnwe3Nq+XSxMjlVaUa4r87iQ+XD/mVGu46p6JIA99
r/6BgB3Z7jtEjHoKbA6OL4S0keW0cGRJNH6LLIsMgiKhxVoXZrvP4HQb3CCkBbBw
rylo7blc5HI4NCFnfTm4fCVod+5VkbxykJJ7uj0X7Rc7gLoUBCW7cqhEGZIadBjt
PCKi5thHpUTF+l8tb8pgMsE6sKW1JLgRkd/b2mYLzpmXvumKzPG+6OPWDIL+XiW9
3Ca9fvsVYoIFTCUCOaqPM9dpAWkCdBugcb6A+lCOySQa0BUGfLinmdpr2YZ+E6QB
CJ1YTtJ/iSiuL/ON4Jj8PCp7oAE1pNni9VSawX7Wm1mPfoCYLh0t65IaMPHqxIW1
ZibaQOHN2522YF1HiJxk8QPoY4MXLO/HARLeUk/WQ0Fvq1W2JuoZi91+nN5sSQF+
QWQTRrIIQREo88zU8X2VCiATnyRvNae/o+j9Hf+SinU4dfC5qhq0Hai6A+UpyZH1
zteHoY0GlQ6rJlztQ5hiKGkF5qRcE4Oe9IHiFm6notvB57Ue0WJnSxg6+crsZl/L
vTAssvsLKOD1a1ZnIslnbZTSZFE3q2ylxuMHJy77lhbiP2pMCk3ht0pha5WKMBVP
h4xQvkdx5c4fcL2jVWlz321udotgJu2XINR4AOznLBVyqC9TRA7GaygPJf94IqGR
oebDWYsJqOBVxC9ObFq7H5JP6tyneiAyr98DESMmWMXxbSHMMVY7IdymC3qXUcki
EvPnZRzNX+j3BwWS4dfUXZxMSqz6OVu5QDQLomkq12sMO5ftBLS+FdbOEg/I5uB0
ZXhrCGk7wy/xD204kFgo9bphWpDdkFZSM4k9Xr94WyufpcLadvepRAKQIwJsMqZ2
Oc5HBz7G+YG0/sXqdGttTT9uiGoVYYFu6lAozErjwQksPzqmzYQ8P/wuntEEasiB
Svh1uCozXoS2ec9dItZNg9wUPOWvhouRsHmsHxpM9HT3NCnrocq1YRRz1qWco4BF
U8FZST97hL2CuJdHPFRQSaltMMXTFB9gBLAN6Yth26d0sPkMcGuV0E+3B0Xy7FjM
5yhv7Iddg+LzEWRxbx+bwMi7CTjpK1yv8DtETr5ZzisnjXWXOcNyUO6Vd+7v80qO
0W3zriblAX4UYv6T9XFGU6rMNjlM4rfVbAQMnvYG03SeWaDjch4ePHPDOGy/w5vo
HFaar6/RY4bEIHFcbbjhVeZH/uJDK8GQIyacDyEawo1ls0lF7GGMF9V381otimVq
aSLEODRpWckZoMqcRnocOKSoqxcbhcC8ZoR4Umh31YjzAk6G08kFDEwxme8q5vka
eV3Tl6QSRF7SCrVvTnIgH3n+FEivCBkoX2sshqGkve28oGHBq3KEuQ3a3aFlPkcW
kSwdW1TPrxd19tSy30qz3IKoCeJ5w1jhwrEHHjatMAdwKE3YSYQ3Lrx32fvrSVaY
jJc/petZBPgz5KTsitEd+ta/Ha3RNs1BkT1Esl82s2QlRhkZC6FwwWs8gjLWQWOX
WsGybz/XkvgjcUGbqnXSfcWfktLYn+M4IQTqIy0NY0LXmTWQ2VOex8d6qy1XWpQt
K1ObfAJDOBdF3XBqYkZr5dx5G6gZE6qa437XPkAe1KCXpRUUtWqcxn/4mr4Ej0lx
QpgZjAp/j/56kzgLUPAh5JLhsbYoooFfI94p82w+DeS22PzcEBMjiRc5ei4CmnSA
DVne7asZZ+885isPQcAw5CYTnYKwuy1p5CJLMEuhTRXxjx929VLDpZOzy5p8KpN9
9j5eaeHw5I54f9zuby4ckasmGBoL47kueS0YhiHg1pTfk6uatasBb7XBDdBgG+7l
KBDoygrbLXttek4hoEWiqP/FSoJ0JkH+huAkClWh2nTOiivYUrKPa44gDscu8KkA
L4XXrZrV0JtWhyCDxAqlaAyec+V/3/mypRLFy7bOru++EOhX1TtOoRXtptNdBonL
3XBDW01/dSItyKGUyCLnRRdVweC+48rwm+kuXzu64ggyauVq6t1N8VWuO7tgiRhe
saRMYjZhSIHBChfPdiLCko3xR+edL5hu3IvboSvTwDmpBQHRZKLvMpgTSfUt0q48
LIR/p8SD4gIs1D1ga61HpxYsivshSnG9DfbONL95qZXqLY3Gm19q1tsBKLy+3Bq2
HoqRRG0VKEk8ysVYoG628JKZvXGA8Vl+LHttOzmOVYJLX9OAUcQcYChUfAdawlnT
12Aq1FH4NRnPAYk3NmCoWRXiU27L+rXUK8hcUQLh2TFgpgN0zCMcaLJwAHV8tkZ3
ZMAfnzqvJcOcLSGCFSX4hzJXC4vxMceJOzC9+6S9jBgTCYMa7fbrH/r0UijRYdPm
8gDS5Rb+jmcV1K4Xnb5khwF9xyPp4FrRT1T0t/92rYQgE5t1S5HMTdb5umdInMrI
h3aHNhEitm27+pPABxHYJqEKmBGThNFEsFBDddnrx58I4IEVyaVGyFZn9jtZRt+e
M5rLIxpd/a7ZHLJoMPqEikJ+YCdx5M8izyKdDyiAS0A2doY4ZPdBEI8Kr2WCck6y
Z8UXv3RacAVkxvLb0hg9nR+nL9rl+fdUNy770zFJUw8BxsE5n+85jhHwJSuOpCfd
qcw3EpsxKED2w/5zvv8IQs3VA3ZksS9S5VPULqbE/VfWZcUBvQKKzsM4RV4XFovM
EqFUYBQsIHLg7iA1sRt1mkgzfmG8DOExWSxyYeBrqjfWZCvOrPGekC/5C7SSHYKq
znJQGfeRpOE75h4MXXapJEUvtUqoL/tDPgOwImrPdfj0GbNLzLPVmp3RkAtYcy5J
+rHXA4UUiX5gTqIffP58BP4gZKA5W3gLR+o/QhSscBEMLWm9pbKb8bGUFERdX1B7
ddrWVSFZ8hKTB9lj8Np1LIfT7NGKY3j+GwSORlkyrQitnQgS2Yp2IGaXrhBEFP6u
pZOXVDiZvq8bZWa17qdWNoOO81B2p2cHyCXxHPAd9w6ZmYHlPoBzEwWdTCVNKX0f
8ZX9CklzaRZT+xbCVElBoa+8xfFA/P3dRLCtewDt/uOQkyHKGxlp4O4WOgOu8xoo
edEj0f65vSIpQBP1Yo53CbLeKl96hP6RC+cX2GJQ4ieY7m+7MmwT1z1S0je1Yb8A
JqcacKwH6G7bMFs0Rkg6RljrKvJWf51PborYK3mmJNmTzMc5SlDaSWbwziE0aytx
aLoT2B9PFpbQ5B4l/+JPS5kS63cFlCIEkFsM6nUF0YRW6Yna/9lNZvM+5M45lT+p
8Mng5kT021acGQ8IZK2pL87V5NIWSYsbtpOtGu5TQ9J8g/7wx868aGpM06nD9wxN
o6JgyHtf5S9tBnoupciZco0TpprmxIV7bYu29StQ54CMku7NTG4SN7dY9NkKaL0I
Cn0K+UL+9iYfrgzmdfyq3ubW22tQkwVKEEPcbHzRYx3r+kQ0IgnIgW0NBpBalpgM
+d1L4m8FOrO4wvXC6rbQLcBv85U81JJNUnBb1EGklwZA0Y0DoHvT0Q/McUPgljov
rjx/as6Qv1ip7z2BRn8OaXhQcjMaFmdmyK/RPLPJlSKpLxeOW5GJBwidi+rRWHx8
9RxPB7SD8Z7ma0xIkjO4CKt2cuT2vkF4PBzqTJvLbJlBNrwQrenm0ZSCBjp1hZi9
jbBmrBqGzwKB1tHLUX+RtJWvvszk6vhxC8qPUU/SKQeh6zGcqFHQNWhuO9ze3+G9
0LDLC863DWIM8RClRkv9eCcBbA8CbAioG7hmD7gzFYZ+/XFE7r0hzu6QCS7Lhv81
OEICQfGqaWtKzwnx3d4SFAy/3re2yP96DxdUw0wVx5uDJjraEzvMkO4YwvkqiQfT
as024AKEh3BPQlHab3JAt5CMiYuyJSsDi2qvasQ9ocx0o6RNBVdFtQmmZZtamCOM
Ux9xU3S4I10meH9xDaAs6irwmvCFR8vRN4fxd+9GQVrtFfgJr6UEqBkm7/LKJ/0o
knMUELUMPq86sIXKNpnN/d+OEQFVesteSIYgRsuwJKFE/OEZ2yHiO7avP8gv0WKX
BIwhWgSisEtCH356fp7hw0EnAUQWanjRkdMXW7zrSUxWdY8Or8fFpQWgHHGBiJ2t
Ht0zaUxJS9ErBSDCGAb6CqeZ8RSjJx5hf3kNMMYK1nokS69fQLT5sZIPnSRxC75a
C2dMne5zv6UkiwfO+ujfgAtzM/o/ULG5M+B1x/pL4DjkORvdZZEzWZGKOZZekyoF
xHnsPxvQ/R8i5GuUM1J3S6mCthu6gnafoQKNySfFZ9PQTKYlOlZy1oS934s1xP3M
6p8g+FzGXDl4qCX4InlUZDirt5fpj6NIPHM1soAqFg5voghHEe0Hsihoi+S8QbrM
79XlGWHKRCS/8P5NOdmhHwaBBeeRyirTSOTY6JjvdcFSzz7hfa70Zsi07b94sDZC
eHZveLKX7Lu9UvzjuEdvr34JUWdfWoQQukVwlGb/FddziCr2tU9eH6Zcv2pgJTQ/
pE8vuHlJiflEadSjhbluInizEMxgtFlWDua31FoCvdA33bpjfFWMMza4xtvOXvL7
fqgQDnIRco93uu544uUT2XZu0wkxFq4GOs4YHvic8VCDy+2vGxVOcGnCOmzjlFW6
tzF40/ldw1k/T26oyWIBgOUz2e+lPsfBEazq2B7vG6uwl58w7FwJpC1Stnq09s3G
udAsFQDkl7thjHUQxUWBd4WxaENNK5AvCKCzDnMb8FQmxqBs6LT9iLQE1Xc8L1na
/kk/fUkBA4yiHLGDCHkjv+3NaCzktlo5LFlOkdq//4Mhs66zQWvnbv484J8E0MJC
vn3t9Uy9rTMD82iGvjIce5kLoNIVBooK2Kw4w+DNtqi2RXsR3gtENIx6oC76jRN3
CzTjNC9ZpJuNiLaI/wFlZHQ9jsRRHtG1pnnn2bTeh2Bhak8azmnFMWTlw5R3BtMi
wnVYy0V29WFg5dKOgg0V3fuRjeYwVr3KDx2mOpY7yrj6xo54v69nZia6JXhqgoSl
drCe0SvDCcxLIGmIIyILStKnvJYa7kt0NGyOOcRJN5flU82Jobc8AEuFnldZWMEx
T9gE9oze3fZSHjmKSBUteJC9X1nN7v0no5KLoa1r+/WhStCWbMzLFb5T8NbBsL51
kCzF3cOMM4W1qNqrf1X/rkRjy97pCcVKsibf/72T3L4Kt7BRQM0TBFbeBNIaFMMP
xwiopmTj+wImQ4LwX52+5uYkSdJTxYB6cnqpMZ1idDBxxc3I1kXfcunvBsZs2PaX
os9D0vkEnvgr2jr2rEhUmRgWCR0Puvr7xm7nJOCUWAwtD8QAsa+TOnzCPmUnDEH/
VNu8Ngv9+nOUiWgspKNnYrSGC6Y3hLceSrcy0WFzQRcBkkc5/8pVa7B+dnayi63G
QIrO7/XPoJnx954TIBvvaWZ0vWPLGQ0rqUgQyNiGwMs2srHGMcrPY9FKuUC6ccVo
CLrwG2zV3IzQN7dvTXbSSk2MTVf/4b8Tgyzlsx4yCL584k2UEpFjzNOb+l2paLDn
PXzhZCEgvP8MRDykL+WnqyUJNg03RkLXa+1F4b1QM1lnsFAojgpph1bPkx/pDes2
R7d/QC1xjQQJ7C/QDO1EMi2Qde+kjiMy6IoJ3YTU7x6gGRB96QeVxwEqP0d0tGoP
b5TDQHkPnui9grvs+Hrsm7XGeaRpPz6V/Xvcvj44L7yaihumAkssCgVT65pPDk+X
lHzPS0KKEc9HrTZtx7oMdEQVqlJ0u9isOt/S2FFuhFM4A+kjW/X4PS+dc18RWNNa
5qS8MCq8nDo0Nz/kMze7oi++xuUAWKetgvUDgrv8oz5JYD0hEaAJGL7m919fqIkS
CNMktGJ2HilI+6gQaDj28DgAO+AcLmTL+AQOsnGXTeIRApm3/Jadnzf9izjg5F+d
T6c1Bu6IqVqxEaHyfunFQRz0y+LtYSTvIi2y4+UNybHOiThzQLRyGF20CThVd55i
KU2qsjFSM/v2edOKzYhOWuCFoBr+MOv7UAjgAl3PFW2uxBUtWs7YZZZbwD8zL+Jq
NDYAaM6J39wowvF7huLq6mUGRe/PYCobCA+k+IGf+VOmINl5fbLuyjB7uxR2nSaC
+Qe0/pzkmTHHwJyMrwHobfs+eKbFQJupRoh8ETlwso/hrYiNaU9iYdbm05OYVFKc
aIzWA+eEdhiVzrKU7CDXt/I2uQCbYGqS2M6Oa83Hb6YHpydwCHulivPDluFEz2M/
srYB9pwMulccpSdeoDxJmRe+CFGt8kY617JeU038Da8+gKDM8pX5AsVpmyi1HbNj
HobicZYGvGkwWZ6Ap1lSP4zYXo/gsK4XvqCWssbKx+a3nNtFY3MV7qU32pHvyV6f
rv98vfhI6K20704/Y7vhOd8ne8qeiOyAfln8hAJXdWLk0s6wp0xefF8VMnC+xkTZ
bXkKvoHVDZYoUuCXi/A2QXbs8MAVzVQGYBaFz/f0Jb2gs6U/p0/5c6f/xv1UK44w
sEwWG66cpnCS18UQBVyPdy4tvyK9YVq34sYReOAy5bjZdXLEc8W5jxyH/093rQYc
PfdDJOdfxd4FHgITNBTX4/Uj3k+F8PnwrG3vys8JLZGFyF6KgL51G19mqSmd1ZVu
4MqH4Ck6nKnx1G8Yk1LoHPQF+9lpW/p2dOS+qLsy/EjwUClNF3tn0JN0CnNIFeQm
yKMEF35k+ZWf8pACm7sl6vi7mKDjNEo21boT/1qn+wgDNKzfEAW6NV1TCXTMzR3x
ot6lgseirR4ut+crXPmLMkpXsgBVMDOmRDTImH6SpJLZ2uX89roRsy5+EEp/5PwF
UTkCcoy8S1ECx5rdI7Tdrt3IjZBVi5r/QHbGjNj23V0AaVavKgsMW6tObvUgVsK4
VgM3U8F4w5fCzEqjOW1Vz8AEFlsmQgteg0unJWcva+CpjQdlZgvObzYxX3HsSvbI
rm1RqtmptJpdDwh76pnjLBeo7eZPfIaDu1Wz51/NsCz+HUAbndPv2D4WdiAWmTqr
t4C+YXnBKG9iryLXWgGb9UNjylR38cODmvI2A75zgePpGMF5rR4piLriJXFr4+pM
7aKdkFJtbxiyEg2HGqlSmLV7hGaPvA5IrFqPUjdz39hB1Tx2Td9PY09kDOkCAq83
cuMcz4snq1m5zSgt8W3fNa8ukRlzQnUsNiGbjTTzmvI0JRKgpzatOPdzgnjPjcUB
/t+oc1Gq2R1/yUVGe4AaRInflIkoSeOj4DPfdSsaR3lBjidvLnAw9ZYodhq9mnzE
F0oIWrXppDTFVvlMs9jMFckgUe0O6IOBHOve3YIHCgklLh79PSo4CjWl8bQWKdgn
ikiHN8x3WeaMA1g8fe4eqmvEiUXlRrJpheI1sVD5tLQeCIKvkYZd96aAGiuqC++w
kj5uZHeU9zH9t3HIjsWU63WelYv0rXdZv54llC+Q16ZwE7gDGqFpEp4qAxdAID8j
oilZljKmtlvUaFLcoyJvw7ir8mMz5wrcIqlzSGGegIUt3ngjJqKhlHBJVLp9yA2z
gi43VYkEa5z7YH606Mz7Mtr8geLJGnfDodJ4H7BEsKFv0kefZiO9lWCPlutzSBSa
Qw6P80LQqrX+f2227/2ACOGIoyPj+Cj3lgbLAF/oaRchQARakJNziZ0P7M7YE9Ei
I9z48JNnOdK4XGcpqUgN8c2fhPdCB4L6jCCqCT4I6LNSRS/AggUEWArETLgPELev
ASlTuC2fgVLFPGvId364RiynjJazfS1ALG0RqHDNrx+xOu/ET3mMJAzOB/5LYLsC
IoinAEA0enAOTEia+060/3aTd07mO4eUr+3VYQI0lnvziICzcpagI5+lJ/1EJOmH
IOyi5YsNdUE6dKPpwfTCUvVYMOg9/uQxW5slGpmsiiNPKg2BL2kxEanlaV2rc/qN
ZJ3+NXewOQXOsZVi/KjndsC4F0xFCelDt7Zxzg1NAtOlGNOjvBpxz1n/GW4ohRbe
8xsdat44yXF6zAQQH7ucOO5sL5p+kB2VZjcxqgZAa30IGdmfF5DhryMqDuEj9ckL
MqJFv6rVDt/CDQqftQ6C6N9OMkiJV8/qPVa8xEOYgn8Fm3QIO4T4XlQ1Cm9vPo/a
oEOLTgzbIQcjfA7ZFJfjNGotf1irAw6Qw9uNErC36ItePVxQmDx/l18L5dISjC1R
rYcPSo7OpI57iuMr8u4lJuTam31tRZdOztoFTZ5zkvFd9TdhPWoWwis4qWDfbqYK
/ZGqmbcJHrya7YQYJdjCpmAUsJnz6qIvUxw/MQjXkhRGtvhD9SCvCZwUeG/Sti+T
mURHS2eE6ULB1dBKuhkzSvVUuuSrYMhh0aN+t2MorVZ9ykmJxp6QQlCD02iWvK2r
EAh8HL7yAL6qWCEuZYFaeqmFg6OxS05N+6yzAGwB2VHWgp+jbsBPp9Z3k8qfAuzr
dVJQhpGTxGQ8TvBEDLh6q565+FjNxmAGfhFEr8MiEwkzEIyOAwCHO0axlKhawqov
jV8kiZKQIDj6hZruTnI7lOGJsmPDD1G5E6Zj7infHFToy4ceZQzm40a+GH3VP9cv
x1TCP67GDWG1p0wvFGAQL15toi4B9GIIhMATwHv3CQ0a0DM4H78tXZKjelPwu9Wa
xNBMhb3yZSX/kTaxK9Nw4e11oJ177SpnF7weTlb1pIM7JmR/fFBinFopuCuzH/JP
OhdgiNLu1zLHdZeMKYRiADWyto8QVxCuDbUS74mvyH95O8WvvcbD1nOFnkCyvBSR
lfvhkrX4udT862SWb8uZsqJ/GB9PvBAXVxAHe+aQpbgu7Amvuu3j7EckDJsnJwOl
8JGg7Q2EYOK8M3Uk2WNhvzMXL6sVZcnbrZ+JZdZ8T9UDlk8DSYVmNgg8nHlXuaAb
1VcSZuk1Zk/OMjeVmuKMbkf+rcrO6baTxEfMlmjgrEUjERr0t+Wa/jnpzWN9OX1n
PUrYQNenBl6rxL1rWwPkjpPqZOULfshppvPO3+dikc9HQOftZN8WEH09O7rJFzZd
NLn5Mzcx041z5UUz79ss/rCT4uPi5BZyRs9m3q9vx6M+M8k+PYsQ8lr5d4FH7/Ic
e3+4ybKtx61cGAFd7BX3BtbJHL2M6jhHk5g+PNKJ0VnXLOy+ePJ5jm9p4mtdXNf3
yOs+zJEAFQ8UEjQbK3eRybERNLATp2MLNOiet0UaWB87FPkVZHPnWZt1ZgbenIev
XsMtzvS+IZv3gzD9hylVq68avuhVbEcZuaCwnFpihhPHpB4ZtN5KZ57oTrfEeAqg
n+LtjX9bYp2UJ5Hhpxx7BRdD5ZOXN0AU8iglmy3/0NJLSLIf4iixsz9izBT9LCHW
Ic/AP1lQeQzNvEfXuOzwBJMkrRPe9i0eWvkBbQUBNJ5vFKWPGh/PT8iOJVcbw+ec
B/FFJ7fYBYPEZvP96g8ncqTQhHyM9EojU7TI1hZI22uf8W7kzu4kW6EXM2Si618P
bGJTj+XWy95CLJXVBTmP4Ix3Zpc4/4U/2ZilNu0fhwK90NsH6tCCWX5dEMyBu6AV
edobczXoXdFOQEf/DXc5Jm1Kyx0cS63BLNJPP9TVj3DUwy/vpNiG1R08E/mSUvP0
7OJ9HAT9mVGgidiFAem6yikr3ciRWpfyq4BWZsH9cD6uNHRWohv8QxT36+DPAC3Z
1xZm2piS/dztpCBIWrhSlGnuDpPkws/sF/XvC6O/S9C+MD7qEhQX1ANmeJT+Ryvz
oIC+JH5FyScd3hpVummnPZtq3iol7BlP0tMBiMPuAG7n2GP/ZvuBzXzwZkP+494Y
AYWr60LGNeB3HL8MSUnIXNm7g5TxNzA/oqeXTmx6Ob6QLNgUyIAz2N2Z9D2ecR0X
1b8TF/R5dm8nwFBkS6bA3PpSDp1/+0TTc5xufskp0cAxcEEnzdv3MJSHIc/DfkVy
bo5tm9UfApG9mzCRLILjigjINjdQ+1GhQkX3ozJUrr9pji6sMO1wh+yUmd+nb/Hf
WJs5K0MJst3d48fXq3aRhNMUvj7AKpjcBvBisjnizpE5w0LSLTzGm6bp/U6RRJqW
wLy4xbh+Py0m//3jsa+Ynp9RWtN14GbpxX30Hofy8HpuI45oces+DC6IvX86wFLG
i+5jAt4Q+yflGT6GPqcS47QHyhEV6EeeFZe7NMZiKLw28oIX9/+fcXp4Qi4s0vYz
vIQIIswFUlVvjJasvJx9/if4EDPRqRBjdsjPwm0RkKlsH8lodxJNRrwr+6/SzIp2
C/mRK3x8JDpKxmtwcsb9fMCgZNCeHmoxBwmv8BlHIF9UJ0OSnSnR5pYm0YepKm+F
HJ/4lrae6EuCgC3rmACOUnIxAVQNE/Xo6HDMEV8Httd7QjJdh1B9uiCwx1n/Hyk4
jxwxOhbyNZn3Nr/qH+YFXYcUNU/RpN5mWrlPNoTA2ETwVrHwjqGTYmUDuO9s21Du
uhMaahJTOE7hvvMDfKHTIj9ccfkxBjyzsMdyCRZM+CaV80X1lSeu9c1HWwdoTkCu
mrVt6fcg912TwA6kaXsLQJqLnC8wCzWbZEbyuqZsGQqtVpGqeYxuPqRp1b7hRp7l
rLfwwi8JzNmtVpbSaoef4NXXNHW9h5Y0bhQGzXbN2Oa0o5fgnm2/XKCGVfd5klIJ
xnp8rt08LCs6RGHFSe4wjj8rBthz0DEKBHeA93yk5+XCFlt6dkktitsaU4O6AxXo
d3HQ0e/63KJAkWm5rYv3y4IhwAbWLlIb9EaOseFttQnrvHPOaoEj2yEqVe+gpSev
S/oG07KrQK+dP+4ofKIVrogI6cFCc/7fZKCUxQNjnVZDDQcfSx4/5NjIk4c6KVk1
GyrC6olp1ABpPca0Xbe5BYv4SJZi3ykND9f1YE9XfUwQj6lyLl3sDeRbJx0Ww1Po
+4GFO50Vg0Xhz6DgI+1XWV5UAjsf2AoTGyWfqJET0TmuGhrKKQlkRu12Qml7yNau
W+JSF9JBnkkVprNq/UjbiQ5gh5amcefXJ2Qe1kKtM1SSIlJ4cc2+QfPcyNGyZFLU
RTjGj/c7dKr/ndlam93z/K4CB4Zbf7COn8ug4+iNp6o5/udSCpDwbHRH4jXMtmWH
a03fDA0Kjq/b/3+EjWgZqxHp9bBT9eRFXrDXQu0d1EFP7Z7ve2dyu5eeGOZiPtD6
4CGrevS8UYaQ2uMDIB3QzMklvyFQUDT1V9Jlw5c5GrVO2q6hmnW97hLrMxvbmzU2
t1LeL6DLoEslzh4hexmNCbcr1iXWp+8wPehdcB2ZtAdCHU/Hjq0NCBvUebGkqBb5
Rzn7vbSJkBV/zA8MyrM2LttVy7mU3h8u6HlyUP9Sk9cQQPAMKoMUrrmQRqyPyWq7
poPuEfBLFZ5MnE8yc6x6RqnJ3xtCdFKivq2KLs0E3ev4TEU2qaN4NgS4jE1GEViP
2ju7kkGaPysJNQAZLy5JRlGriaLvWciD6mtsCXmJ5QUU3awbUbs3w7KCJ1y7l5Zt
6BM0t/P1FOwbLc6j0CkQN3pl5g0TA3axDoyM3b/2CmMk2QO4hGV9LtWGuBJFm5mF
XpkQGqzkJ6crO1+ji5tpBYAGLtTdIkMdCyv+PCBTh8klDUbqI5GXjDt4bNK1ajT1
le2Ikwf5PP5eoLYyjaRrAAIYPdM5CzjoS1xqZ7D49u3rf3o+etYCEPiaQfPD7wqs
rmtyn7JUU/wTJu3K6GTpLQWfg8tf1OA16DXxQ74zE9PxYapaarUTaRDZVLpETbet
+Y2zy6zt2zXPvjIzYWsmvSVgo4ae+rRXM9N5ym42XlCciISPn9dsqgUx6Nwoc9xK
SjQqSJv4KKdepd2d5n5tKjFNy/+GIIKnSY/F6+RTYS4Pxh1wBnPglygHraK7nZ0T
MwiYVI2Tf+OyZ/WYeDNqYMllt5FN8sOa/JFcpGSSr/zkDqkvYlzVgRTlY/9C6huW
x4MFW0wQ/Dig8Js1PgxdPNJ2SVNlxa6tadPBF14TATBcNPXODeFA+nnTijTZh86G
Am5eN9+Eg3+OCdaSK7z4ABWHeNSEIvmhRYoW1J5lsvhu4Sf7j5nWAxvbjOXLQxnm
e2joZ6zrdZk8lgLIbT8OMlh2azVUHupBB0gySJNHyHRkNJA5Fwe5jTEusr2VZsME
FqrNCbXA7Nw/w7j7WFFIVQFaxNZDkbF0Xv+Fs0a8rAoosnBTXQyzHakVYDcmSQCD
IQpfEcBtMPagbl8IdIiEzTNxOvoHcWx6U6jaPOWXa+w5Ns1wJysHPw6Dp2i9Wr+I
ixISFD52Q/TvalnVOy+lwdjkG7eQuaxYhRbSMzEXxy/qN1Y79OYr9tOs5ixsfGL/
DcKceM9nj0YeFEwVPfFRNpxK49t6JKLF6+VcacBzf7llirDyXtDml2kIqMMwouFl
vWPhteQN6FvlhaXa82MXlS6+NV66BLSOU4bYkkP/B2ldR4F52RCbbZCUlEnNiwsl
6HmYMh3C0rwZnR0VcrTZaxTSx+rSIAdYso66IJRFyPu766Toqs8BlJQudWeszGxq
Ncskdf0EFabFtNT4DGn8SrR8uBWHRKF93jXjZG5iy+Inyx5Eqz17TtXCMimLh2je
wbCl1b365KBrBz0cty/2jBXEE59aq7qZ2h5My3EQtrcaNDVQAmsn7E3eDifiGb02
pJQxQj4nFoP5kkB8DuGpLhME75nPiVzcMvo7+eB8ITgXFDHNOMOlN9NkdoHnW1Zi
cKOp2TCdkjWKyuPVvesq4OrtW6TQ7M7gRazSIloW0KbqNTY6jOR7RKD97Pgi8yUL
oOKElzUse52q+vXzqyFTrGb/N3ZvggFMTOPVja6PrdurDPo13QO5js/vOhZ4nMHm
dFsXxAvW/qT4a4//kDUG98QTSs4wAkqd/J4KVCuiCXrORRNpTlhvHAUoTEkuqfKS
csniPsw5E0vZULxubM36DLcR7TZ2SLvUFYIznM+u2GDDJEOesbqHTsGoepGTL8I9
QykVoEUpeXETapJ3lzr8/nBLhhse6XRjBMJlPIUE/g33YivC4Bd7k/noBbKNXbua
OCP7sslF4BTW56HOkRFWG0mbO4An1PLOi4Ur2yQfERVxBfk/Pfpa2kBJaO8yx9an
XzY5MkcLLCR549+2ba+Q8BHVSf84iUQmywlqrPEfUN7UbUyzGqbzBm4/FTA68r7F
sQrDRae/GkE8TH2/NOpsIjotU7LJ+ADOBuaIR8fbMJQhMP6zZ1R3z7vosBJtX+fK
ybwAk3VDtpqvCBmb/za8Y7BH5+vlu5tjdB9sNBy2QRz3HzF6eaqLaVqM9T8AirgL
9umgr7/OA0iI+4cdyC8sSyJsRj2keQJegBcov5pZPF66VYJIUcc1c6oYDQpTND0u
n9R68Qt8FzxVG+iJ2eYMp/3rX/ypvuR/01XXAHFdY7uWnn3jJuYBerjiOF8cL9kk
LAG9hA7iy2n9Fx8QKDg1uwbH2Ux/1BxEBsjgcPJe3oSJ+X6KacS5OOUM4+IhzUSb
tjiHwqlL9CyEMOTIAnUzXOoKwh9CWy9ugS+3Mz62w4LPMYOPj9T4n7jIkyyXAFJY
J35K5Tu6OSDy4Ctxg4e7WpASL/YM9Io9S3Qzf5uI2bnRxID/+fPuNTrl9SuFaTQx
bP7yht2FQ1gsUAtAA7z+YKguFT8J0KgzwtBYFiphXp7qvUYr1QuYs7lhgn5pA5AO
EBW0lkmHbChDYNqs/uh6lvlw+yyrkw0QAklCxfW/ww040Ju7oRbIfNZHXFt1T4ru
TLC60TmK9x4YKlTWI3IzSt9jPJwXKnTB5koDrR2edbiMeMem4UMexMDMBJfCPQBp
Xce28emOGUMkR3M5GGxhhzmpc5Z8fOKPQ+kJwpjK4KgCRHGSHraLebexr64zhZAK
l/TgyQUgal+zhuchYPCJB/SzN8qTRtErhy78Ad6kYLw2Qvl5hEGAeGMD94D496/s
MVldWC6pQKuBOsjzc8kIEEBB6nRb+gX/XWSHApGSToLTzaJLp+UlEI40xWRYA6iP
of4cqrwrUdAeL8QaUUCGHcQuL8zoz6yhiIDrdL+HzLO+7FuHNYc310JcyCnDZD0C
abs8ZvmumSKolJx/yipa7s06Q4m3sb9a882MJ7N/xzIgpsUEArZOoLsoeN21Xz4X
NeE8NwijapFgGbrBiCXUifuWbz91U62inCxlLGCSwBNiVX3k0ykaKBJhhovTqLeU
S22TLRz4JaLAWXlkvWIFGxwG/RDSLG6x4xtlP+uLvt17q/lxLQSMqZTaw0UD9K/Y
g8ITy2LPolVbLBNvYCYCImkZOgBgXaGmVvAn5yD2byHtc1Sx1Y2BQSnfYa7gpuKn
VvtqeF5QF32M3rl4hXBXWI0cGVYlp9bdwlfyltjnFAP6eOsDnHVdFI7vLaCFBJQK
dpOMnTZEH91HUPhI+yMpR6eK6GBPpFHEyQDwEnoTp2Cmq16/5M3k+bcLXogJBEOQ
9kr1r0+5PKr0+W6wzS5OqgVP6Xj2TZdSk3XgFdXcxF1nuFILncs8/+DWNjszE2NI
2WJd41UUV+J2qEKjhHWPcjqiJ1QAppUpb9MfWIZmSlxWJrMhBpBoyrzVUumfK+6U
KOouMV29xUGCD721zGC0JipFvO/+sok5Mlgef58c0vvZbWOXm7Pdo/nFBFVcAlvC
YcNULNhxYrw6OSxN59wK/TgVZwj7ZrOOosxreBdzsGvGaNHlHByIjJK3jyfqgLrz
9BAtvGOPtbnQmHwL8IoFqo4h3YjtpMsEaeUQ1xwKjD28wueCStdNnHT4d6O770of
5JZFeSTdHQLT4zV/uLBoUvD2JlM9X2Phv6DJnQa878cl6iNBAi0tt1JImC+kum/L
kg8MHnCbha1Ziva1+MYWgZ37RVkjHJmVnHk8o2QaEnMYAZKrUUqH4U1OrrQ9BNxh
jAI7jU7wc50ofNMMT0R+wgjJEpWn7a/BCpZZ1OGlfi7Il0Y70LzvC4peNGCGGsoM
TWFx2lNvbtSjeYxa9rQHNcgGcKiqB6HdSmp7MK+muumo9Ht/rh4vZgVbF5MjAFxA
BTCG/mX3fqp/S4ES7E9WP9m2aYvCmFNYTpqvOyS9thKpDsYEUwTGob20X16mrtAE
5TdtzVCLeZW+xbPLP1DR1XGfIuA1ElYKkZIDtyzaC0OnGks5WWefR9c7rHVHlGbI
3IL+IDOikIzBctubl+6ZTDgt093HfUz8bKU4Ff9ZZdsLb7TYS+TwS3SP8RaPSQ98
1VwQcLXMvyRw4ZVfGIXi3g1wntCFB6s2ISSF26b+neaMSkTQEW7/LPzF8ycZVXFe
Bdgii2jNNfjURZcR3Q7m5uZh6YWB0rE444aPvvFxbha70sEPxy6/HCFGzl5pFreD
4gsn4+maBZAVaTAL1b1aRh+McXUcKz2fh8ZIOzaHGTS14ao4VO1Drrxu46PdydGB
JGLpElzi5oPOtbsc/wtvwlRkPTOZuB5CgMlXTv3UiC04T+IDXRyAM2zKpoSrHQ1W
h4EGwmhdVoq/HSIScNWoNhCPHpYlD71ewzQzb3xVpLW82TJvGl2EpyQQ/FR7sXWj
2yJ3m8qRx7YOlrv2ihnWh+RKRjp0mlxy6UPocwbyk+V3EngHrdAcZAPiZ1heZ9DB
fOkEwjdYP89jL/NKRLJRweJ45HBwk7vJs1ROOUDIg473/xAgD/IzF4r32JOJZGMb
p28oPt+YXL2fVazGDySpxLRjWx3h+UhjdNm2qahCXKl2K+NrbDjZN6vI3AEZ6kFx
Ma/n4Z9hgO9obSxFHSKmHdYxT6V3PAaFeNeDn7PDSUBTrPkY65v0Pa6BXQmbMBve
Y6mhnPwlOI+nFzZ/g6bseg3wF/Dgsy9vegSyRXTKb+VxOXKGYLyDZUvRW+bdEeNl
0/9VWSVFwS8yRfOQ2RujfmP62Q0+jccfeKtdyCoeP8D4p3fqHSUvD9FiFY3h2CkI
s0gOyESPzLT4NXE+5vvKs3GuzmVzOWiZjAamYBEb+dhQvsgo8IA9BF6eXJAwydEf
7kWnXwlDdpJhw4eE2+frYBpo4KfacCjwe2ieEykIoHaDpAtdi1D32+fljhsE7ZSs
oJvxdwrv47PPYw1fPrNAfrZXTbslt2zk8FH/qTYgqiqzzsAWpLlMp225JGJDO1gX
8EkENHNp+uUtvUVSu2Ci19Nk3FjntxF7ciHwfPAOV1WtMD0IaVC8sg3qnJZKQ10o
xzsnieloDq/DaB4UhEqaE22en5UMzvsHXmh+JHwzN6hCHyt1gjUQFbHETUxjYyxC
K3eFz/hjhZD87G54/ewqSx4dZF7bRVN523ma2+yrPBjRjNwxSe3DeuRft4VjeFtQ
GAElCS7j/uDslnP0juCvJC8rANnecrT3SGuZO0WQm59NjiOCXWqnZzSKu14dBSyl
vlY1E+wzDFbNiquGt6gfaWl+/yXzx+pY5E/ssjfSqp5GAalnby2beGAJYQ5XhCBg
0hB9SekiFIfbGHDrLvarEJAKceufE2E4IYFXL98usPWjLghu3E1BKNfys9EmmRrg
Ywss87vq7K74vcAo7WV+7HPI+RZIAhUTG9vumTmcGKrEDEhLReDvF0tNDs89uk6M
YiQ8DJm3uAsqqRdtkQ/Tb+E0I1ELKfFol70IXZAewVh9QM2HbnUVC1upbcMQHx4f
+biM9c/mddHJHzMw5zk+YDxEi5y4qOLsPbprBBLuXNr/5VqexMX1ynNUBjYMZ0er
gd7bTW6Da+kK33+IeC5UajpMNcMgKfET37Q7MhBOhQygGICpvB8ysKRbD+wqN6t4
zaontKJTnBnAfgUZiLczrdUdvZKvRbnvh67bfdCBaAeBhyjKCL2Rm80XbeeWEseO
nFSYYwSIs4rJUtCGGYu+VhyLJU/u4ZjGtDIFaFjYefnwE59g7tggELAYCiqnjKzM
bPwmsKsom8JtgS81uxvgPgw/6YsAaaoZ6Y5F102DI6zEGRsM5KNAfAfd4wEcFtRm
RYJa72vpzdI5UGpjM8Wl/6wkCqtDcrKTbm2hVl+qknJnNvb/ktx5l2/jBIbLCxSs
R3rLrDtdeEbsDn8hqtivMh35RhR1kWjQmDwE+6R0fJEnm8cNK3FkVTDndwcwlTjl
UdP/Mkg3TtWZx7riCX7zr1aIj8Ghhnjx7WZlYObYHG+wvh9v8Y+v79NSgJfnB6v5
sJt2YAiO7a7/KzO142bKU1XTRNV+TMxa6e5r46hpuQL/DEYUeIJU0MUCfi/rkWq6
Jirk4x/GpTWg6i2qOsAv1HxE+XqFPCOnXhTD01lJ1tqgXzRUiw95Y+dnGDblwxNB
fk4Mm8QUCR9WgJKuDZdejsUtuQuKcoYzae+oAYdwWlU5lXjN7sxSC0cxCAQQ3TxY
sMDGtRV54kpxIOigIAAz8sncFDOSPyBgQEgnAHO+iEm3r0J0KWlLFw/AfxwEvXrM
LI7mCbLUIXqkG3jcaw3wRQNLNJR8l/sXuRbpmT33W0BufrH5vEQ6Da+yjwa02uTQ
pKr9yOxehv6jEpJnZZY6JLcCC/hVp9rvFfP6kd4RZjxeMyBvVx1R6Snj/kMqA3Df
esuJirQWa9+sE03IGyNCt4+QmzpiIzXfig5gLUL+07AKbIzs1uqppwCM45z/jLel
jCF0lfv/IEO9CeKcdHzERVKv5hyffKs2eRb+Kp8fVrmXTb5y2NGr0AdHS4cJRsM0
xNF4a2vnrVH1+AWRYq4yKe75ZrUKk5Mtxff6hrmy7/96ITALEAyZD4mKoeXQ2vTP
IhxrkexAXyquTb/bU/99Nmqu8vHzxBMI+tnsQMlYqDEKERB886GyOqwswRbBSX+E
S6Mrh3h4AfnO3uq776G1XJ1ncw6oscscnT3pbYNKzcP65Wow61nPJakjZqhWnObR
4jreOpjGkA5/vmhcgiZXNT4KbisgNAIixr4+IFEu8Nz3f7m5tVgK37eFusxWbkd2
v3UxHkWD8qf8T9UzG/F9n9HQIWIc367zbmmo6dJylqKSIoHOK28jTx2lXIUUOpqD
q8NM5Tgyco4r4PJ0IXOwKH2esCDY4+jY6tsOx7/ruVn76CTT+9mKkEGK/HfWlRG7
el9C1L/jJi7homxZ9fBZVrbXnPfpXnatr0ReP0rGs9LRcLvDHqJjHJQoH5ayjxzY
Kgg9vNhggND91oSg5h51ZrYW3PXjd8ekVuEblVao7s0pnGjy+GKTNfky8DZKGn1o
5Owq0O4RPRPpq/EfU2ixdR5wMVMknctdfRnnNHI/YYW5qxqwTMqKfYWUWcsLZmTF
b/4JRQjdfnN3F44ZK6KEya42ioW8+y3qgvxM8cvXGcDA25EPhBIIC5zsVxBVGPJB
Do0lT553oJA8rW7ukbAjjDLTI3bpVLiNji9Cvst/ma6yL/Ydfqp+BjQViKwJLFl0
Y6kmXezXyLn+2b/IRm71naFPNHbaNStXjk7RJPJoGMSzkzhDPbk2nLoii0ZMih7Q
kzEeSMpAIGLqhkV2CNGGWkBMCf1LMq9bQ1hHBkrHYUaZ8+LltbBsaslprZcdABDE
GR4RCvzmn/jpf4i/GpMKJ4xv/5qIdno8r2pk1HbRMjELAfcMewcYlQXrx/X9MibL
DkicI/h2PD+Z+mfzXT/+c387kPzgSCEJmoiI1mZCVdpjfBMoPEQcv31UuQtls9T2
X5jVyHvSNDb+1pOMGSv+o7nAEpfaSWFm+XgfgEoyS3EtlPQ7ZPxwoWbEqkDH2TVD
C0XOQVvLRc+8qtHMyTX5yiquXQP/jAiXojbAs+qQP0zHf9WGFN+UsUOH2ouXwtOJ
AIeA4rgbMZDIe5rrr+/4ep+6ehXAFG1Kl8WP2EUdjsLKMZXLhEkXXfpbrPc6QALy
jiPhT8mptABHvXIpDKD1ryVpQSug9Qw4gwNsgVY6EGh1pZnKTIadAyblnqwMTsYk
K78Nl4zF37wQ8eI/DiXSlCT4FjnXbWPz6Ktlm3SoDwtI58L8KufpXpInku/49AJE
lZmwmwr6aZCNGBMVcNyOvLJ1hvUc3dva5Zh6h0Wd0yDZxkjBnmi+UHR1S8hsBnfR
A8V682QX3UVFRGIp0mcoBN0hd43pu6yiIrX80H8ARUsVLiH8X/yd7Eaj9nsEtEWx
5Mh3WZEi8vB2BPYxh7Eg5UETjodcGL6dycqEmTZrGaWTJQTmn0baaxf4cuXu8q0x
fSB5FUukmve8Fxbp/DyIheth0OVsZ4mCtf0psE2qYvw4z+nOu5q4Jpkqj/6WI+3B
ninbhyUFn4iy9K1/5zp+qgciDOABrsx8j7Jsk7gWHv9hqJLefF0atzNpeCF6yMKn
oE24s5fSPoLbjh/AH4Bxk/DU4mcgFIVrM2xzKfbxZ9dC0oX1mZjSyA9omtKBmQ1z
xGKoIRMuPTapSMDJlciDbS1ICOUyh/zXxKS6RqtuyulKYl+Ziy55AEGCG4/TxMQx
lJFK6VzpUCRii0CZROCprI6QbG0TWtNZyeNB3tlvHRs7jWZ5NL7dDZKiavY9YGyM
zvimkuUR3zQ/d9ihJeEupVlx9RcZDmON4ReOUDacrHk2bskDDb1A921+L2VjL2Z4
M049cq40Ijhv0CQaQ9sVvnkyhtMyhKmnlMp881QpASNtgArJkmvl73tIG8AVIr6B
d9MT7v/jG4jsNZMTxP7yU0B+YUkM1t7BHM4thRMlXFTWsAW4jVhwJF5dlLAYWUJI
ASmRDUfyYuIvxNYSSVgyaUhlgHOjmcs2CiSIwIMUiOUmDgccffeQhdGORK5eSYm+
KHMs3jJmy19gF5rZXABDsvYGrfHjP08TKApkzo3miwUnwIO6TbOBA/nREGKbrNxr
/S5Tln7gBDsc8rE2joqyX2kJoyjizMBH+/q3VZ0oLhBUpXkrEf0GuhG3y0ySWd5a
OAZy4DTxlGH8sttI1qxiy2XzAVXwx/BiTBu3ZMOWhC0N2+/mxez6Af1eeUmikH/7
vLiVZhzonhRoY8+t+vPQUH87nx70rq9/jHtia67uMscBxiHpifT6jx7aO2S661lK
dDAyrVGxOUW3w5fJq0bZVqU38HPlkGxvbpj2sNxM+ksdIC4ATvi4dQSBWlWsIH3y
RoDjkoeOu0szoGXWYAuQir/leExuyTa9umF+LMAPQSRd62d0M0z6sKCJNpx21wma
YPbb2riW0wqWI5qYr7NlQhWPpUjM5GuDsMre7+3xcRzB+cndai2iW/IMWn29t/Bk
V9bJp0zl6b0sf04ZkPIv6jmvNg14/IyP1r5dUt9ACBmka67aUiUQUydKChUmGHsU
Ti0Yl5oo06MFdmwJosD6rzATxc3+xJhQ8xB3KOukDKvnhmroPu3NLS2H/n/pAiEM
Vh5Bs6mhh0rn1ojvPUprDkCx2IQ/C7G9j3Jc54b7TGppfJtPKUDGyZ0i8pfDaDMK
H71U/zvCQDSBbjBO29MNPgcwDmHyvLFNwXnira2xPZrcAq1eWgqkYz88s7AqI5AO
hX/ij4/sXq0yKZ6ugZ6szGYWF/ZF0UOtzcJO6teVMZHX07XmLEsn19cpDWrPtSvD
ImXFIOJO7ziI1N6aGyVWXwuXfZUMU8ypMGqHXZbOGhaxDHB+eswU1XtY5Vb9W5sW
xUeyaVvz07gutC49psKk9kuGCHA/H1qaRIkM2Pnv8/AIYfjOajWQxv/EQNw4DcTC
ovrhl54/Mlb4n8CnGKbPFaiU0+AwUE61e87Fs20BJXsSV0y6eb3vz0Fd4S1y968s
0TtGA2drjzIadmdai/yJPJpbLbPub4R8wzOTTR+LX1kvrr8IOxR9twA/G0hM0SyE
7L3Z+/o/3nHur+btcPFASnyQ9o/LgnNtHZ9NzHq41kky6pnygerVAC0bymD4Wksu
O5oD5moqW73pd8yL9EEOEydryv89Gp2Wn1SicFnWGII3PSZtGLj95iZwJ7lmNzoT
qU+VZRTcjvScaL6P+FlOc/FkOHeN94yrDY0zBk88d+cgBFBPJDFYMBMunxSFocR7
R4M0aQ6WYDd/ViW4C6Lu/HKTgzXs65B3CWlHd00OfuZ8y5LlNMhU+7xHYfOIApXb
Yq68TzgLLQ/39xTr+rCcszPjrIU+rPbjEOFrXW0AUd8dXGJm8mfjePuYJIz71cc7
2xPKpC1eeprsqFVsV48/ffyCIerNNinAcHlolIVjUaErMRKlPAi4VhU91FLB8iFC
shDyOpak5+pvHtDlRgtWLe979dHjN9PP/hnkX9Yjhx043DEN19rEZMj/awrQF9bn
S4lPidkFeGzNJZufhXHX1C3e3+46MHhn/3HtcMcRvyFQrTMlhIVnSvTy6IV3iFMC
KuXZVmUS4XRNzd7IxLkWtZENiDXLQD/oEQ1RO/65E9LxFC+zZ8PbTZdT20pPitq4
X/Iogz2jP1JDGnOz/ohjJ0tXTuhPEVj4x5VQvJ+R+0gDfs5K9KqfY2hQckR5nIG2
eDPh9FLWPaawErR+1FeezSIFrV9tJ4ZkMjOvtyzniWJfc5BpwOpKoXGy3BVhEn+9
k2qlKH9nisNOLI+2Xqp7mW9wTMxDJEoJyAgqSGwLcskr1Y5DnBa+WknOmvmHAzk5
Ht/8ELc/m8tDgjX3eGmBDybTtjI0FkfNV5N9FmT40Bk0eDKYyPg27ZDl68YmECp+
UoK0TbOK8ZLt9tYMUMRnwrZfww9Gye+f9KfBvlwhciaH0W0/u1D0zCM0FxuWDXNQ
KUWY1rgDziaiEtSmiOUSjnZEprhFmBCBd8mNt+N5LbnvNn4aKZKTghX9vEERf+Oa
2mudJl+IekUY+vTpthFGqUfImy6XmtHTXEBfMY7n2Wi0h2jBP22/Oar5y6qEVtBo
oGNr+eH2tGWhbKkNYzsmAeRjLVko5hNGNy17oj055ykVhEiBBOIGXyZT+oGMGwKy
lT/trSR8/ZbKw6g9A3gaJZBqb6AGNpEQTSVFfS4aRP7Ut6ENvCYxb/OuBxxB9n8v
ggSneiRUt9d7vxl2T/+4ZQJ5YJBNkOYZVTXBFnYtwiSutyyHm2awMhptPRIH0R9j
Y6tDmwXx0nk0yS08ii/3fpyVVCZmnx/+SAg9T3aWV4t5c2/Es6pTkhQXRssULMhL
rNjEGEdk5PJBceuLF3CYzYJa4JwGNlkzwAbYlzzsGzvCtUD8skbb9KkERDos4tgp
aQHgPG5Q8Z8SV9k6AItkGro1LtV7M0Ey7Fg1f7GBRPqnn6FLAbvNquJDNh0A69hQ
Hptng449FosqRncYOamC3dQwWo1tvANqwWIsDsx/anag5jN3O4xtp7+XcCwXIeyy
5ht3Wobe/X54XqHWk048QFElNvRAhtECJX6vxBS4fdECjeie0Hf+f+23IIfsso15
dhQTnPsaSIOEAop8kTaWb6YMNuzgTgf7TOLCkpSHs47Eqd4K2JlC2l3L/OmThtMM
lNNl2aeD644puvcCt8Ow/qkk/dZUioeJ0NU+HN+p5bD1Bde6yqdsa4gRol6bf/28
dT53pKsOjrhy7Ar9ldmJRV7MDYnK7DG0XsRFeMcLM+Iy+GQRxF0Tok3bWCAnsj91
+Vft7qp3WHuFXjhWvo/8d2gXxRKR5YkBum2uTelNqaZBZM75nq3LVKU27u6rUdCw
lYpgdDtguNpenW2N8G+KnxooxBxakq6I4gJ7FY1CWumhNKITNb8PaRFpzOrDqFF3
nVyLDhXnvLCdtkj6MXuH6N15zYQe4L7UnX3xYtsoqbWMrf9z1+LevZt7NgK7SftF
iOvx8GtWUUigbo7ImxgzuZtSE/6oB/hOsze8BH9DLWXt33ZQg+kn7F2oNEEZisX/
QWhIsdoFbBEQ8eP4tmc+Y0nHZBe085w3N6h+B7I8P8dsWBJIEsomY0NhZb6c0HvG
teBokChxNTlgXJ3jje/+H6SFunW82KnaHvVoL300BA2VMt3l5q/3HFq1ap0+a9Q2
XXyDaYfqGPXuIQRT6d2hXzEGDF8DAZx0RIogUQgWz87LN17zIx/PWoi2szsUGL6n
IYAm+Cbx/L3ADM5efefVetj3X5tKdUdNbdphtv0YN2AvJH/71OBCeKdbngNOxgy1
ZOmB/ieZv7UA5F4eCTgf8dOHLs/EBkDKftD8SiLyb+GLGkBIr7gvp7kZ4m2AOjoi
Yg7AjSBlBEwyj8R7SD2RW88ezpow/Su0kOO/v11bceHZ1skzLbl/urZz2lR2Yixg
p+5OkOS/1ng9vbryQqR7Cy6qTVG25Qzv8Z+ZmRlCwrYk3zYkxCN5nfAnS5ayAal6
GiaWF+ERUfs7leDAB20STt/3RdFdDjzwBvizEF/GtL/DIQCnhCvRzQ3LOUF/lHDO
6883EM7wZ7HrlunOFwzm9StlJ2mSif9s0/+F3DZXqHbBTO6wzgCMr2wADZKP337F
pjNYZYyrD4HbaoG1JJeu/6zgleCq7w7KCSrGkMmVz/0UJiiK3dfqdAH8rD/9YRrm
OLdgbgdktmhAftd7d1K8s8WdX1gkyYDBI53AX6or9SYxV2NEm72WYtCGOxnxjsDC
b9fzVH21UmkKfKL6RG3N2C71gMVUp1w8/eDjfa3W649h/utdmcg60gvXCT/7ghlv
xLbqTzPxG23x1dUgjYQcv63Z7AvG/ccRIPS4P4YQqV/eE1H9zO5pgUkk17eLLUAn
5o1sc6uXBBJijwx9JpO9AsLAsxrHH+CgRVjKCu8+Z40Qu+G4puX4ld3Z/kXxSXEf
7vs8hHUbFEl/DyJyY5tU6aYBQz+W5N//1rcBNJRzRkwTlXve1k4VC8Q5lsExXsVw
3y00ENFGmHvLdzbtYDJbNvNlloygG2XrhEFbpbMiHgm4vK2Vepgh4BURgLdUetYu
E56+KZx94opOmzkpMDOogu+oUtqRccCH49lo8wItL8R4ySId3OZ1wvfQl0NSr2rg
UOLRgIjJc2OYQJOIeCv8GQWUfTZhy/+Hzw54mgpKchkRDgSCBec7BJvt78FbfToh
a1VUH+u9E/u/s9JFg0KTThqbXrOQjiUxJ+K7U0MB3eycNCPNRFRyAO5dK6QnAzpW
PkoH+yGKjbx411DT5tEaYTYy22MoMRDxtB47SHHp/4oU0X1rfLkipaQp8NaRxbzU
uKUlkn7GLw1X/25J2sPp9wB7td2ULstttBKb33iiSgfVYcaJbyEU3bpzTbhE404T
lWU0GSNSIZN6cTGGhS9Yr/K/5Jt6D2HR0U8fHtyGUY7OxF8XWiDdFk1+RR/IXR9S
mUT2sekbPv9OjeXnaQPBP4K4/oQrATEzTXLDZo28pqbqSCbBaAtUx88uqxXepTx7
Dq0W1rlRduV1zRgALjvOevvqZwe00Ht9BFTh1OICQLhvaLZ90BC1WmSwGa7uF2pv
+esJuMzTJyQQI1yhooIDehd6bP2CruXMAQ5sGct9DWr8BuEV3Ucf6Ks97bITjrpd
rpQYJZs7NQZNvcIP69nILnFAjHmHy4ALlZXugbbu9/Gmb5E5xSrKY6Yd1eoCg+4T
cUoMgwYK2x+wakmG90hxa/vxLUqMl+X96bfUo5bLGVboz8umwq6xRg2Myw96JZfC
IeHI7Zh/eqYarnI0MSAqYVQMg4Jl/7g+Y4NKqf9k8/cCFYmN2xyQbwjTPg0N8dLS
nA9VT2Y3A9CvP7Sz39ALghSlKvc5WL0l0wGDJt8T2VVrJXA9dc1PZfjLEjlPfv80
AppHfD288zFBBO6MOlDYt4oPcQtKiwsm7wjRDoh3fIG7ZQNO7SX1/Y8v8pPDugbn
+/af6pelqROQ/NOkcS34yyFtQJ9NYz/HxNGX2gMzbylNl0WZ2DfHgs3AODVKx04y
RPOpnXoki0FP1izq7JxzohZ2IDW8DQmTFyCFIoCixPcITnWl3KTgRTLmH08QJ8cE
cpSAfWYC0lEWb6jwH3kD7U0IBDGybaTkSIpm2rQwCmhrREHRstWdocRPX5cCq7Fc
is0gGY5eGEAuHygJjAWCKPgWFVVgiw05uBf38aLLfHui5o4AUGJRVWCk1qprerKp
f/2YmUkrProbGNj6t9fo5UJRy53URRsYjOxCepX9Of1icqD6mL3X9TfMp7/VTFEH
IoEsfoarHjgAbCoFkB6qGil+A2oz9CJDS+PrL40HQxYYMgSqfgpOBOYS+X4NvZeS
In0LyVyhjAc1pPHiYswEPMsaUnpiVJ4MebOBXFYHF/U143qy+4GeZkxqyND0de2H
UaPsnq04YNh0cT9vksORYeTfaYkT3STQ6N5zGwDzSAOAOwV6rakPsbSu1mXguCe4
/tjOOVwMC8Yf7szk3V6soccHVcZauYpKJ7Sfrz5vmDzgDRrRKdOddM6TSjDXP0c2
0zddh2+FHcqnuA+Jb1osc7w2K/xzmkkrgyda3kSxHpmj+AHkfTxE31jcTSPzMlhq
7oBNIxg/Fj/dvs3D1ZBonbBFWIJFjFhqw6xFWm8t7OQt6Dp0Eg+03oi0xSBAC2g9
QrgY7oMAGwlcasTNGFgK6LH5uZQoqP27Zl31jO//0+ID0SCDNe9pQdsr6hNCN/Fx
0V2p5bafDen7EJOgsk5LGUb76AZ9sJh/uSgzo3Xl9pAtmucnWEZTjEni1X02i0iX
7Q2UWs1Mfwvr8ZTSGx+uKwmyZTig1fkWAKO4W740kvHs34NOaAZJNEKkuuJWT7aO
kKp2u0XELyvQ7uzUSX5KIFXvbzq/1D7ieXIrRjcC5ypvMu/Kqa9XYNv5i8daR40j
ZXHKqotn48Sas/R5pjHf3JsXK5/tmlVxbC7zKZLL4iYU26HoO8FdjZYvb/dbC5F+
IsSO1bIRqfFI3bkZg7M5PCPOhP8WbYUwHfKFGHQT+vT1rZRV18+ebkFbx+/vv3aA
xjSscuFhcv8XCn9fP5xOFz0huVa7+YL2n3LVMF5Llb4shsfkR7E5YxgCtLCmeNJ1
q1XQHIuIGwf6kpDJi2Ds02+yZthAhDZ77O92miYUAYRzJ0anH2xKvSNz0NFtUah4
uLjrhZ2RqjJ9OY8hj1ujLJBOpCloOu2Yjx4v7rhRxXjvjg5QUVJNCSzMToI7vQy9
qhoWhXI7IyLBYOfSaZKG5xzZmEUGYmGBJkfUMf+Lz0woQIpBdUnC7YGvhzCaAT5R
0lr6PHItZDbIi3cQoe03U2ITulB3lKTkDUQp0XMpJ+/PUK1Nxkyixw8wKYtW6TTV
138/SLZ5EXa+oWIIXrhI6sp/QlS1W1HQ7QiUUkpYlTUH8Y/+F5LSSKJgeeld17ED
xcsDTBAD9LLklDGC0dFBWTTig2wbIWN6PbCgshjdtebHvp2K9jvTvVuCVM1mGkPr
4pwZUlUL1IYhWqyLpHd+fMuANc8lNG3tR1uQjh+5iCj55KqTCERnFbYaM1ksx9u7
DFtmZ4oPKrzKdw0nJbrcn6u13Ahbz/Iw0qNjbyuY6JNyLITE9vPOXPDro2t8aa5w
s23x40ajvVRsHx2D5kNq1rgBZzN6c4VWiYqqyQyS9F317ZE7w5M6l/r5SwumiXV4
36+puw/9WGjypoNorlmArQTKFdp9kjD39w8MQDsd1jxoUm7lPGujEamcOWr4+RpY
U/FYKG5qAhd9ULy2Tx9+YXo/MpiRgDhEk73y1UFQtDj8GKMDlKUBESMy3dfyJ/wj
HG35uVlKCzkND9QEMYLl8/WaMZkXdpKgDJCnG1v1clRJ2M9FZPhbgsVU1E80ZW9O
4f5CDdLLTON9KJXdH/JVSufBAfc9GiVYa3IgKXXrNsS440ABLwlLOd3rXxx6kWzY
supGbaI4Qt+IpPIfEMW6btGEqnOk90CJcffysMMJo3vHgzHXZ71h9Zz0AJVpZmLh
5mBkpcqso1iHnUVYYC/UmIik/zeobTktnO8qYGMTzrU5qCOvJ+26ryRadAUJ09sP
QMT+8HQBO0JW3tNEMhSuN/tOYjDHX7/tLIgF7U7vE7BpW9c+k6OLix2r4B6Zr0nE
fD0yvrZqjmcziQo+eLOsOloKz5Qyz81CjppIeBVJQF/I/z+y0+9Vn5ssdJBTA5P1
BR15dVKWJddZQYLdQ5Lv8fG7uJDMlE1l3o8nCYNF+t7Wfw6z6pOWbCbyosQsuv0c
dmvo7Z0cJGxitgqWIyKLP0qKkKfVkLfzZpee+JoMZeIcWjDhkR07MFGmvWGxbrpS
zQHBdarSFLJ2nE59Fzk7kEqMCyV2UXCiN6pcDuHF+WFS+n3cIjwkr5lIR6aMj9d7
2RywLBxdoBYQknuA7Gke9HYr6tEqslRb0bvZgM4nbNG7kAHOHGdSYXRhGYiXDsly
HvCKY+f6ci7L5i2aBe42Uqol+keb3wxKUwnPr/xiAXOYG3I/LOeGPNduNjZe2321
VN3XQFNYAmBU7FfL+q9GnHTeg/m7ikuIREu6+Ky5vjvMlH86EgHExIIP3teY23fh
DmJDwTCnjThRHtfqb0p/LDcTP0d6r5qu4Emus3kDMqH+vSI9Th18B7U6swwQNshH
zkf+V2SxYvCrgUDEmpikjBtjkE/NtrJMC9XtYtXyooj5f0wyw61GtUGdxwPqUsgZ
bowbp1qB7TtSBygMy1PvzZfCROp93guGYLMo5D+t7Dme+KPOB+XFHtQSp7RvUxEv
5P59XCKwEw7r/KHaTcLmP+nfGwu8CKnNyNeubph2nhgvd1wupIuCFJje8Mgatqbc
rxj0dJVy/O5SEE3NBZRH+bXffYdDPz8q/El1EoH8/WkYYR0xC+Pzh8pEWGnmvRt/
YkeoR++R/f9FlbzP7E810J1yL3KsfLkzuicXgCQv6LRkVDCnWC7y90Dv0dajZEKB
FdnG/GwF0JanCoUNYpWnvf44Eh8OtH2pQCuh9IceRPwY/kJj15ejapL4vRQnX+Xo
Eo5Qg+c8Cpxzw5vbGk+1hBH0YTiu/MqJa3A4Hood8VQ3+0c6uDJD2G7wSbTBooq8
RanD4tyjJOlt5yzAJA36kx21lvZaSO91eUumtRABWutAGioPZJ9i+ggONRcpX8ci
QWtxDQEzXMT1xmfFsKbjMNSItU0YwbHr02XN9zewNXpwOd2slzSoI2Fco9vlFx1v
HrpsZc9X2xzRZiNodnw6bckrKDMqPqadMGh2d0U7jmvTQlPL45QYdj/Y5/bkeTG8
s/ibFENT5JURzXtK+Yb8FhgvEdQVPLjfnTc8/rG3pofs+rzj4/HKV1DlUf4ms8rX
7Tk8ejtjMNviEGziv3POXASlfsuLu1/KTTyuVBFmRZT6s2Qa1mA/wvDiQ1qwLmQU
ZGCW4TFitstbxhtRBnwwdHU9frU+O6SiIq1SL5AaixzOdHECSd+Olp5GGfjGp1gB
wVkw7C8dISKFya/XlLaWz0EW9VBb96FnXM70NNkYsYWvunmdqoMxUvK2/jpfAGw5
DgLgV6SlSYiqSgXYVB2XD/IN1cOcsaQDN/LG0+6BG3U6MnNdL77zPB/c7Viy8TAT
XCrcKYBNNOkMY+lDoUKNMHbS3/VcsHTM30TMYPszXWnR2ZJAI8csdHnTfrD7AT4r
8ADh4bfFoQTKosav6I/DqJXGsebUQ105RY+jMeGwQ8z1e9zsVoP9B3dmkEwbdOpg
S3J1Y4x5hSzrKOVl5wdbui4I3FEsXgJXPdUWNuQvBn55fnnL+v2W8vb8CjdIErRh
MniTyi2pkQMtl/VK5weZsOwu71/qGhFGsv/Hv5+tgqkIqeGgXdDtHiQk+rZQ2uQu
h5KfABbP2Qkr2Cx6rNfRSbBVAcUtNKNzrHhc3BM3vClSUTx/xUNo5UEaD3ACDRrc
bOyWYx/l4XE/GM1x53x4g1sDBETmCU2HbrowmLSAovoFTlBMCXGkY1Kh17asC1cg
iWED1zIKYMXNiOWmp5CxxuzAZuVG21jUgdGa70wwlgBwKTXyYiLXaZMd5hWTwyGb
8IONWZNJvgOx6iNr4zAAc7zgLXBVBKS6fvRdOkMFEYk+nNrlZ+z0kTBstW+qGJuL
lOtl/Gth7PWtBzZsLB93Eb03bZmRFJ6+k+VQZjC1fOWRvcNfnZNMkYWgQrHzocvA
nSN1bOm0XzV5jOrCPEtjo4aAroEwMpxmskbMfD7xQLlCpkkN0ZNO+0kvJxP2bw+f
RCla9eDEf3w7hRKvmNvVObOq3Xn+H6bBzEslIQiikI57I4hMe5jnfGYzKabIqWDS
FTQ5i9NILQ/a4/sgVb/4oqp7p20acefoXGzHi3Bory8JWjibWGtHvZd8ZVPi+ZPp
1WQqUcj+dBlk/QqBtDpCWnl8DDwC6fNH0Or9j2ZTqpBrGLHjPWQXa8PH9Xuzf0im
hcHFBT0h69gZdFGcOmVk4Jf7zoacsLHL4ewewyK31amFVnesmJJPxXw3MJL9DBmk
9w6FroQHmUL68Gpevu4ysn9YbD9reuln+dXX/IDx2Iv5fyYkFBnauG2JSgwj9tDG
FqEa6CDUlsGOKq9vtjBFetPuV2ecII1H4RakcsQlyt+Ta6rdpX/mgGWpJtQGB6jl
s5aDHGESXWp42zkvfMn2xjMMhHLNmPItTQ8NGidjrSjGaDgwJ3QIoG1zTMzmZO0L
sjpXvjVCA0BFox6iyYKLpWnuiQDviALkLxcvgenYkHfJ9nLncAQF1ejZj3/8qvjh
WerQWMJWbesV+OQ2SPjNJRomdbnJKUBW5mFut6gHvbIg5dFKiCHLQpS0YaK9jbp8
Q+KB+YacobncQ7R+JSOlCr+Q23ZkzC9e+82nxByuC8SCRCwtU/P7uHQlRgAtMlMl
oOX5L+8rWsX4qhBHrmbnohGLCWDPX6t754PeqJhwzYXwnfMC+Vhym9T+cl7HUOLo
nvn41iw6B62CBTCk1oNxj2D7h4/tHVoYijMsN1ObtlRXoVUGvKXC+x5RKf67qvK+
AqtKwEvtPS6d3Zr+nQ0Ch0vIPfiCW5aY0ii/z9rDliYKY3YUCJ+XeFMCGAYnT0wz
lEsZHA4QEE6DJ+ggQJCVnz7bnYei6t5G0FKi8++vGRipK/EACDSERYI4XBFcx9Y7
aKex7RAFVfZJdisVscTJhrwnNOKfU9NTFLSo+WasUTQ0fyk4JtMf1OFW9TfJGsj+
dKChoO1RMvqqW69G94Mk2NGC3FLCJYD/xMQAQJ7x4MxaWKcjPEYTJixUdCM1fMA4
LBEvNrwXJlm2m66EJbB7omPq0UdRSkPZbMkm3Nv5TKhTIRFDTBd7KYlOjLjqxDTd
ixCJMkH+tguJRsn788t5vVfnAhc6SWZsnAIbA6T4dAptgaz5LzvKxjXx72kxYPSf
yAPHVuFDbeLYdLtCSjjPNUQAF9UO0NyVEpooVZ9i9AtRCTm9UNhYl/0jhsd+nlWu
CYbVw2ly3JNUcQ35hJEl+QXTMOfRTwrIgU6G/wStDeHD/PV1ATgvYdmHqv9JZ/YS
oKNbrHNGQbaMBQGtYkqEpYRUfhpJ7h5izBZz3KxQgK7Ht/HRYP+dOj1rqPA2bBdL
Zabbg0cj9UetMa7tq1EDQoiEsVzbumZZY9k4Ln0DKdP733WTDVrPrff1xS4sNRIe
hw1xEVOvVPjYtNJqvv9b+qQYNgIJHp4kh6kjVcM4Tt8AnUy8rnoGMoNc/gef316m
UEDUVq1Iv49g2BA6byDTLvaVHfcirduKrA0unKMlbclnnt1u1zhKs5AsqjR/vxCK
gD5/7ZUeybd0FVmYJvWxTlAFScohe5UhEnj015Zl2niL6Is7VFup/1jrBP7x+Faf
BV+ofK9wvIVxA0ygSyZE3UrNjYRpEb15Jeux8Mt1CPchrR/ZO1KGZEqxeq8GUo1P
Hd0eHTSwSMOM20Wbi2PLkoaeoy10ZH1LGuiZ0S4ELdwWcUg7015tjex331CuiPYw
AVi+/7AWxHudt1OjFzo07jeQPUn/boi5L33vQrtHvYRRP9ShOFsBNUtU0Iju/h1y
P7moFTnO14j72YIyYCvqGEruztmd2ykZy3ktOaHoOOstKauMBmuKoGRlkCEBEmJZ
P24lA3CIsG5sYPIjTV5zQpRJ37b1PKgtYE10NWk/cDJ00Ibur7wYT3PYjVf2ne12
qmwWAFObpxLXwWKKZfAoEXWhpAoVyA2Gq67Igss9tKfJ7+RvDU35LuAQ8UufvPeV
99n3gCBRa+VOhVWCf7GMKB2MZKDtTSgVkibBwcPPqV+GnjOWiCr4g8LOiWs4yyLB
I/ZkvYpU5iubjLF7gzNEjtJ6U1a5hitcxAS6IJ96shvUy41h4avkQyS5DqKdel+1
JFReaG2WvGzng9UAy5Pu6svYRwwo4SZABeeVT1qxIkORRAi5wo3T1thn1DT9ctlT
V7kEZSOrFiJ+Z9HgBb4aXKnkL7jGmwhA9xIB8LonB9oQcC0gJjsoILHqqshl7V0j
6d4Kfvjl0vsohyCySWf0PJXeyJiMSxAN6xOnLCBVoKrx0Qz72xxHIr9M6RxbFoMW
huPrZncoi8BMCtqBREzFRc0DhplknSUmaU6DlI87Eob8KTKWysr354K2Tn3UgO3r
YoSF+BJLRjXeLb/+cogWBsngEcfUxgg3XICnWwOZ7MBIPbs/fcrUywf4rgqsQjE8
beSdcDTwQvDf1q7ZH8ZnrF+9kOVxLJ08tJTyabw8xntFS1dMyk5Xb9pmYxVUyDwz
xaFSkeyIyie3b1fEYbAuDGBVpM4nssxxFMtgM1fn1han7/CVn/zRQCmAQEK31lVx
EIr3WOPPGJ8AmPuXEHlnVzh2/WCchjL1zc75A3F9MSb0pMZ8JYa2W4VLYupEDbuY
nlQWnDD3zNckdcrHo2Rqu+7IFKPrqYcOIfJSJzITpD4J5TJoIduE6FPxfmqLoH66
KQHiaAK4ak2UfN9FK1DJ2tCjx9Z+YFiWpkpjpUU0W2LDsBru50+1hr/MGWBJVk7+
NjEx//ftYpcC8Qjvyig3QQNTZ5fZbGWCbTDJuV0q9AHnFpsDitp+0AWn+U/S08m4
ZFQiMZwX+0rg4DPY6RW70LZX4V42VekLE/De90NDIQ+SpRXJVrSzFMZQGPRg5rV0
kUOkeNNQkgLwUOL758FSr8qu9x/LLriTQo/CC8MhObAImyGHVSmvn6b45CNl3N2W
rVJYrWsKkwG85DaShofSykWQLIOSKyXYKwiXK+DQZR+6O2p2uGCwbzGuhv2ATy0d
W1jXustd7YYz1DcObjnVHmUzZRvv7RJHK2dOP1e2aD7zvvlKG/z2HQ/Xjy+zyecI
NNoErqzfDfeMkmnnbIe46nMceRJVNDaEPI2qceXVJABwZIiEL3yATC2t/CX4N+pq
Q3209iBkQCQVQwQhRuGTn7zcjVl+L8cKjo6617Gv5RSB9CL/ccPJE+bGW3ajy/V3
c7Pkz7CQEM7TWvhPrwFp8IZJJ4Ls8/kk5bd2DHoPJD/a2WIMea5co1nklgFDLCmF
INOjBEDcgBj2vxLYV8qvmI1KlaRPIPaFyVWOKhaVV/TnUhiFSB0y3QUCnwuWeX9s
RvnZPRL+DCdaVM+q8xJEyy+jiqGYmM3TDRAUAfBne/tOQOSLyU4jUda3w0SqBaTV
mGosj0i57PVdmlxRw4b0quon77VmElFlWdktnwI4PJtMIKVWMa8QreLo9W8dpIxZ
2gcVnwNtq2bHmnQ6HeyfhZtsL6OhEFU/A63q3l4/5aIy+8vx1rLZ4WMHgAuBxjv/
i5IddV8C9cc5XcQvoV6+y4Fx2sswJoIWFTHmoVbh/ChTyteP56HTc46hiAWA2X+N
8m04vRHgXHzD3GmYLr05g9z2Hop+Axr5hYtlqsR/8rAUqE3QtxsVmogpaVG7j3YK
TE+o8wmZQEubjbuse4lbjQXJRNnopXMLPeoGClJzUBwJlezqSviwl+KlqwJtLsgW
4xkCVVLPVsvPlMsLvEiNrhFZPMjouGrYIm8kzMIaULVQ3kSVmXFPUedXManlSsi+
OvglAF9woeZqAFBpN052jbJL1Dki+Ueh8YF9LFM56l1kKadADzmyMlnFArfcss8M
eJRFmk6vw02VrBWx0YHJ4bpCztHb0JERQ34PVUVwkw9F2VF7P5Ho2miraCtaYQmc
MKoy0GIEPtxhoNBxbHrLRvqBxYER0dazdRytT0iND9JSfa0eX7OFE+vk9s6I5U+I
3aOw9uCRt2xfdZWHgLIE8heCpIWWN2uIV/qRmMpY9COGhVSV+a+gCmtAhfLQZvvG
KMoV+t4slyp3xziRt8NYyrriFz+CpIdAH3GPXrRg3LbQScNVnVOgeK5MGNo0Aj2B
1Nxr400X/JExQ/6vaLbV9Y0NDEq9/k7hgqAO3df86NplhqKKvZV6FVNW/vuD6wz/
R/PMykHeJZYTfap21sLKMOrcUxwgjVo3kD8XIf3E/C/lcaAKYe4yk57BjnChvekz
WeQy/Y4wk5FBjSI51tPnQ8bCh4U9GkQSH77A/5QXF+Y4Z6VCPyvSPJdDZ6OTChSB
iW1sYkolco5z+fq9AGgwLFo9SHq2oc+0M7bMJjYICNH24g8OTVlpuDfaaTPEz4Lf
1K3ESZtgDbb74kt6fwyjW1Oy6OxpOHGyo8s+J14gCl+40LF9JDOj/jl1junnRaw1
FVpFAdZbYVf90fXaRvUk5agh+vyaq53Xe4oGAxlMed8pzkBXbG3zivk8cB9PaJnU
stRevlKzGPy3NC9C1an2ejPosu1S9BgWKP72AEjhs4ih4er9zsD1K2TguG5KoA9n
0H2hYF1mutZOCLhZ2Zw/l8gRhrr+c9VJwCLzxh3jcw9DzsWBtp/nKKPZlIYwsSiv
GQRa7+cZmLjrsPZpC5+5xpNwoEbbNMM7qPTAUXeQvS9+zYvxQngvsVccgD1ZgQ3w
vXE8nQY6aR5fry7gQcFkO/sm+tO0+L+eg2kMnG+KSzdjSyb4ESTaVuewm3spbvr+
m7c6YX9A5VVOWE2G+XGsV1QM2S/f+pwESbCCIwi8OLesUH6czFCOm0f1EFxBxuaf
yd323hevY/nnB8m4MHPaBuZtRKdlNb7Q7wp/PAEAcZgpwHrQJ9JeaQGOqdL3oDJA
eH6QCqrIVqWTtP+Mh4ZDM1OBWIr2vhDT+mmoGjo/dUt1DvhxxU6YKCGCZNJS/CVz
vg7cOViHT34XYRk1bNzb1NpvhSzJFNllMMusHe5a6DQsLYoLU8IAufifgOckjsy8
1uPWUBR9WE2iV32zuMduvX2lV3FWWzY+7BxUPcxnJ9wE/VwBgJKZGEJouI0H5uiY
hL2BcZT01h/V2YPcVxixMesL8iVLhitlJyjjdyQLLpJw+sQ56YRKTHRwmLtElUP9
ws6YJp8n5B6nefbWmQSOFyOoAGmmugUgH+D5QWJ62vRGbkbNnVoAeYcxQ47k0v+Z
nZqXn1jcuvqCOEp3CSm26b08R61sNVwlMZarvPAy6pwWNE5B9Bamp5n/VZRfTJij
6fHWwrSKvN0dxGmuXUw8TwjiDN6m4PIi48IBDiwsQeyf1imPjTiAlUrg0pTElC1n
maUic6iQh3/ecmlxXGbDxTNlTwitcO/Ho2O62rVV6CYMjDuV7tIPQ607mcFoYZa5
rfvmxvjLHNdVrl4Jsn0iUgZWWKsduZLoZc5f8oVaJ+08y8mVy6o1orEEeUoiQjE0
OG3g12m75hR7UpAmCT8jjrCrUxbgSJle4ivHoixSU98VYjCcwv00Bn2Un1ikqlW6
2CeTuZzG8AoIB5/vRvz3WsMkfSHCOx1F5IrjSyzYNt7RVQjKlMBVbLvyXROjfn1Q
1sScKrB20UrfUiMMBbu5i+oJC0cnGWmFNXNWYxPGT6N03nvuUHBrhtlX8dHRUxFw
TFSLKR8UUEdxDeHsldrzP+p/6JzNnYmXNxxShX5qtcQdvVTxXtJAnW5Tx6Bby01M
yV2S64FNjeNrcBDSz7ysWw84HDmSk7mJi4aXv7W5rws5+htgVoDRyQoaR1q2KbmB
JShwRdIZd6davzzV4d8wMxcTCWqqCJlw2WS5eRseEjhvy2giXIo7Uu+hEq4yG9FB
gtv2TmfvcJgzEPJyY6gHUBNmLPgdngAD+ZLNRErTYO1iycQP13erd5laXh2CsocG
1WGzq8f9KsRBAmlr8cKZBQaGVE0AT5KO4+JJRA8F0VX7Os9usJ+TcFR9j+rneMjW
73YFntGqyUI2JNqY5d8MGcflcULBRVV4eeuL3PJNhpyrcgeD4GqFd7pb9uEmVCvu
R1hgwOyWNAcdDhbA+ENYFF9scYHGJhDy+RHA4jtXGgEdCwIU9zQu0vTjTT7IbmCW
LW+SO4Q+0vwrGxw0nkAo9hQlxIlmAYCAKtekPkVa/xf4SU+9SkoMnWi8tl+zzD8+
KghNrODkbJ//T1LWBTAJIbnnBewa9NXdTUv3jjNL8yS/WF2xhXnOWCDAGOLdh6bu
ufZb0qd1hRluqocmNUGU+TfEnW47gUulSU0cdMy1UmXAgUel9G8rjFUxFEF5utNJ
O1OuyHwfwN+FYeAeuTpYsgrJdbTx0HudSh+bCn0UKD7GIo6dTNcJpDq3x3pZMxcI
kd6JMXdpJ3Z32UyuTPIEUorSAfmEfmg5H1w/YFta1pbD2patYIn+el46+JeBbAOB
o+VH+CwUcAOktlUP1XPQJ2e3ov9liNOijcGgpf68pnhiHesqKT6QOj9r0Z3LV/fL
rd5KprNVA168ihbdRTqgGapFkWpIIAd70c7mdjTN6kJ61fsiZx9ArxYvRGadWPLk
5ZKYcWgP7NngJRpwqaHEnkEawF9CSOc1K/5vdcVJQfDICife5fTpYmiBMDe+6nds
iJhnk8YSKsNT8Avf21b9UZ6BJQRZDXdbx44Ix2jPCUVv+EvZ60NPs42JEUZNRDC/
IRD4LUagYnyAoU8b6TL7KqU7FKB87CiUP/P1TqC6QRtvJcNUVuoBRKBQDZhviQqc
dCNicUn9xcWURAkzANB8PDgyVCJcqVZUkQCnsK1D35C9CNSDl7juKq+tcqO+IIM3
DUquSlsRXx6lQ9X06N9CVYMyGMthAYo+31uSZFF4nKEkdww6+mNcIA1/GornrFUQ
xeUd/7ap5gi1qrp0eolYTUKVmmXnEbtSSjqW+I3KYu+A5xt9uCsH64Ai8DrYjqeA
WGSwsISVYCQ7L7Y3fjymeRCgR/xKiJM/UBXO+lI5yLluZH1T8Urz6mwSvYSkO3zR
opUHkINTUZ1OLrn7S7qa+EHynj7svbOWNaohQxXQS/cDZLnMuZx3rIc916DdZlWR
rSqSe9wKELyUd00Wq70iwBm4202os9v55NhuNFJsFOK+tylZOvcaPYfWU+imf8wy
NErcw92HAhiybgaHiYv4qJHEvPTd8v7cad/CEDYC75irdnYxtWaQgIZ6in6o83q5
Y8o1U+N5i3EXBQsMEiJ+H7Y/kEkTT1yiSrZIGg4/tsynrz23xyzfk4trp5Gjk50E
iivi1w83tPeW88fDIKEb1BXWGgTaIZ6523fIhfqg5GkCcNY6pPymFOqfPeEBLo8m
/jIccnRDrTa9TxoTky23WJC926ErSGrmlHO+jgXB28L5w1nXHX9XohJyHdSTa0+i
EUr6u+66lvaRyYZZshOQ2MGMfXs2Ysbz/7uIb/yFKKo8qsMWK0Akl5CKwJVbxGip
/zoBpHu2WYbFb6squyrcXXgxne3KFQ7MaySVHFeshVe/jAM/GuT63Sfu7rRFObHa
o3TKZpMOMRLeMSGVfve8fLCb4vk+cW3D3uVcxbIKV5DG3yrc/4rxbTkoyiU5VH6o
0NEOcTYFbFo/WEvJHKoBP5ST97nyj1nzU/vNl73U2omTqQntK1+7sUk/OSIKDgxL
DvjXKgiMHbAWv0W8VTU01ypGQGcTfiPRrApV69QQGrTdtEJmsYd/0LgqmFhtpqSE
vsWbAi/JUH9+Y/YCufbDPFixU/FFo4v6JdsvH6+L+UqSKCvigeI2GWx7pCAmApst
rCQCwcrf2/AqzQIXV14NjTo5luB2iT/fOTa9+3scNu15zjev6UJlX607cU6LBA1h
O+sUUAN5Yr8FRVndi2v9kv2VptewJuL0A3CC3PziD9I89HxNdinjdLvKrRmU0D55
TRcUrPqlVWTxkhZzS1LO7abgBB70bnIsS956JblGoNgR8DPtSEddCgklZUG0D00d
OFXJjQsItzQ7u3pKAM2eNxIvu8rV5GeuWTRtahbampoR92zZglwOvVBgRjZqnmDz
kgeVxS6aCQp1gVs+vBG2TZbT1eShQKiajBiJ0Y1jfVeE/mbl+n8oC4Z8lkZkvBPT
Pxdqb4lg+sZ7xtC3LqgunTa4WLn/vjo9X7aPqtMl4HCEhVvqaqD+fOpRVEpX1VzK
grppRZsfBrfcTghJG05YertMmw7qOgyfrwuMevWDyXSe4z4SgcQf+ZrzUCtIOdOZ
prZ73SrjIcHjbA8nK+xfLhJ5a5/7Dhp2hCeoVwMvMVz3uY2v5EBsIF+cxQnu2YD+
9OC0sT4aYHPPKhfgsPACjIakOcQ7InzE4woePTdLHZ9mg0fJqLPxmEGS6Bhi+6rj
sq5Ni4/cQ9XdTCID/fFzrbvHdeRGgCz9fmlBn4h6qFK3uKjRq18s45VMxTX8Tgw4
/QGgG8WxAuBWtj0exVR0FFdqWwYilaQ2EmR4wkVnukxDqpF5zAo30/NxAi7SQOzK
IcOmz/MiL7jb7WROlwa93s1bjuXbRO/iASkHFrjDuZR4TSjay8u5JIs/uAU68A38
gSrnO9UiY1IKCH19B7lkptGL25MlhOCF5Xip75VILcDOVo3a73CUnCEGPhN0CBMp
O0Jmu3/B+3ftNS8zFx72Dfu2tZJKhnX4b59VSk7WxhIUwyXWZgIBYy81RTg3Qr6m
Em71GrS+gQC8JhZj2YvjIy0spL/KaK7dwXCoPmDbGur51N+YfTETTF5+mg7Iznq0
yR+vLBYk5wmlMOe4nI/ZY63uwWGCyt6BZftCoifMsjKRvXbrz5DwfaMIjHGt69rD
/1F2XAnjbhhAjujVbUV02guF20xjKfpmVF4Wpo5CebxjNOREiIEqoSOgTAkAk1zs
q/7eLjks8FnDSrc64Ovs1kOUITvY12UIL9Vh/J3AHjXXWMaddDlit4pAvFFgO/6n
aqxda0WCfgkF9PYGvlM8Vj1hN/OIfzMIHSLMwY5AGciRwr74VyOj1KJkVURzWB9S
ucDY+iijNHV2wqQm+m4hhVAjp5ARZ0pjp49I7I+KNP2EczmmY3k7GQQcc6VadfDi
1yx65fjBNGb8je/Vpq7dVOxkvTfpPcdYMeFopW0WVSP9yNaO5GRJOUbs28ZS5TgQ
Lkn+XzGAq/GYn1iK1mwtUypDfZ1H9QhiaKXW4XnWc/sGXNRsWbv10bXuXHP74uBK
Cg7Qq2lX/o9Bv3Am34BwocByDRLvaC8iAFLVIAR6zp973qKMxRUHi6C84dXAOeRX
7LYSwO5sC2tSgsBA1/Z1JXPji+lhxz+7crcqgNJ3cEiy/1XvvUgTOrYl9657z1j3
7qrbHKsArVsqwvCRKtOb6zpznXVOoz31h0/iQCAm56l7j+DcQOCCcF+fZW0sm/VU
6IRGOykwWQd77JMgcOo7o75+0u64bcqZD0X4YnchqB6XIcb67uJgHn/0gYDCAoD1
KmIkyi2tH39GTDhSFKYL1UICA6biNfQU5ao0COLdOeCMBg2jMLZY6ynxM9nHIPTM
52fmm7qD+Swn9mGgfRfJG4XARYOzPIku9aZvKm5D0j6vDkM5lM4HK/GfDI0cBv13
YqgK7UG53RvU/xRuRBtIcZUVhl+GRomNBs1BZVKQ7uiJduU8YAbiXXNA1N3t9YR1
O+GxebzQZ5qp6nc6mdxSM1a3BLlR8O7gacMTYuJU9qJTQ2KISBDcgCGRsXusSJXV
OyD6mDt5p2MtPaQkpdkULANy0w8ZwNkvq+sabarmk/zCo0i7whi13t9oi78uDkAY
lu+FgXKG/8FOIOKT1lEwLHpZtL3xbs5ULb1P1R2fwU9X3mUQHMAXXVKCyJSMTjln
RuUnhs47QnhWaPdgguAzngUzr77D6TBoR9GlwU0NIXyHGpjh533obduNvrnLglhc
wi2jo5QQ/VuhDC/JjvUfVTbso9IZ9K5Vtwz1bb2sBnZekIj8YTYokQ7biWApBwr6
pD6K/js3Qx2gfKfiUZEY065xDU6x9blgIF/aRtcYRfkmmQkrYDO8Syv4IZitP2gX
IeYQWFZFeWrXjs8+95ZsWhPiLohcnLyVGH02Z6D0YCBRfITsfv5Z2k6QzHWeUTkU
1cc43QeFLHX/9zvXICgKrICXqmvEFPndB22agVpbgeyExs2U3XSZHBqWabfN3z0n
2easNT8Q3XkTeFNwqS95NvxZzMuUdn1axHJFyH5B1ToBtgcBoEvsuzTjOxAwFeUR
Nk20oHycRxRhOoj6qXEV+vGoKEpakDyXFgpBP9UvOMszLGiXRVVn1GwvyxBmftwh
h8+Kb5LevslZU1hICyY4eGRI+QXXlz8/Oxn7Ep8Xtjeqf2a371pV8tBGhSqwO/v+
Li89RghjOdPP7g4jmOlkH3gUnl7XuINGJ22H5n1KCpwaxWac7wxQCljZsm+C9GxX
L2s2wu+AA4KpDTGp5immPet4T7YhjXfNqByrbE9Q0tyVL4DhJXojinuqG3VgBvXm
9je7AnsHmSo5saCVrSy2Pm4KZxUp6jGI/TOh6CWn+KGVwVy+Wwyc6K8fuB7+NEzp
/F64oakMlPnwOUF8YLFUF+7dOqkQRav8wJlambsH+arq2Kn4EALK/jCBixqmmumd
sUxMERzZEr0mak0Q1t0rMMWdGGwLIS2rsjV3P3hFEhElvwo4UGM5P3VNKO/ZWXPd
+FFpOKVIDQCSiHEzYUKbBmHC7pixZlqWhla+nT5TsGn8khN8bD4itr4thAd9CbU4
pMrR9m/KGPgJ034x2TCWWqw/61mm3LLLRYJL6+ND5jQ8BvFJxeR6pPJc03QmJp1p
s6b0wfexPoz7vp8/FJ/lHLq7S/hed1+6UPR/fmjuviGxAmckoJuoCv0bFxBym71N
+bHMbd2prAT4qgzTnpHrjRRwsxbPAJdZ9Ez6oPoGhwEbQ+HZ0yT319EjIlHGO4y6
iFjceMGYUpFKPbMKXJ1NfEy1VuZ4NYcN76GPSMM1kbcFkjt/WlImwjJoBe3eURB5
vnrv48Gc17H67Y5AMcWEIfOwiwU04zP9WennjWvfc1oEhncO6R55gfVJIhAClG9S
IaGu0jCJtgiMVO9/OGxQ5NjdxD/kTNoFlD4s4oaJpsqw8HbaHJzHrLDQ7b0qQC1u
fkiop/oCZcS8OfZe63n5L8OIG+Yg1Svxh0WIyh36utaLyCzckoTm7kSu8mkxYbRp
qp5jcuRILW8kRRmry/AquiPD1dKakm0fO8qzefJjzc+Sm+jZqsngvXcmEYzzSugP
5NgHkZCFReNLegpZ2tYFJnUwSicXZ/9DMzfdUsIJ69xlK9xW7blijd75SuOIA8ff
Qtpc43FiWXzSpOwYnFdxXzbg5DAcfSJ260ZV6M/Iia4zMFSoxFwyYomlzeYWIifO
JwVU5loKF3cFU+iSvGsFDGIVZhokrOYymrgX/iJKz/gmESBdtrdpiqR7pqSAMHNF
dZN3X8/pvsuut7R7o/JzpCi3SWyD+qZW21j5EZUIqrRhxV+IfnDmCFeC7v1fxoAl
fFAgl1+p54bpFlX0Zs083gKS3ZAk/ymkinIEdSNpvZH/XyCYIKtKEWJ0ECHoS4tK
m/mzg2HhZVMoH/rLDOP/mf1gGui+5zDlTIvtxeVXA3awNuxdd46hqUcP14ugCTFh
4daoKG/DLdfHiFm/kxpJD43xVkdo9Ixl3ewUsqV4zXx9HF97Zj7zDn9NWFYZ4QVr
N3qrkYDUfk8FioEsuaVHn+Iea2N9Nhxl09qlP10B00mP603ZJpHLKtkQmGIYVwcy
aOLha1Izukp1w/6yS7tGD52+r3/as3jOGcHVKVcOpCMFCF1BCF8CAQjl+TGAcHhk
Xp19t/BQPa73n/mMp/9bkuXpAIHBVoH2hM9w3ZpwFPc4QftgzIGTZ9UaUbQwI8ih
7wX7VX9c80P1ckp1osWBuJVMvtEX5KAwqzFEH6lt8mJNulx734yTVwCvyeouBfHf
YBCkwy+VI4WtwORJDd7G//dOvrW5Q/lK0PHUUcJf5wxAMqMtksmDo9YfZiUCI/Y1
RKim8Z7Ex+0z50zwPcPk/1g6tgAqS3loKkNrhjFelhvs2A0mxsaCkZKBMIXIDhq3
N6fJjZmogh414Ne+gpX/ZIwPg3yYzE4YnOVFNgIZP+bP9TujXqvpcfwDUOEsTqc5
8yysmKA5+supDEHpOOVbg1k0X/rOeHNtz1+85uFF7dA7PXg4+kXtQiqCCOtCR/Tg
MS0jIx29hANa+ezQ5KP+P50d7wl53fyLA078OdWnb9HFECsg9r0NQspcKoqZ1zAR
VX85kuReCjPvC8lDiH8gevoZJNaKDZQRVHu6jOIFerCLVd49APdS3DRMucKpcw4r
c2YFtNMv4+WALFKXiYyzw68glxI2w+Lpx3faf0r3WzSp9RaPK3IPmMbhElvKBN8M
cdbHLVDPQJ7L3rHeujnylRJxTCP4wctoVIq/y8EoPMJ8YIM2XTtRDoMjrGAqp4LP
qxuoGzpF+eMu+nly0XS4K6LF2H0wUtAlvLg+aF7GNZE04NjoQgOCWSZTq+Js0dbf
Ofeunb1Xpi8slot+d+WKjxQlCOOI9fAV0Xabgw0zccTettmDRC5fIfV+qvluggc/
u0WlfkQIrcYVSOwyhIIJcvjS61XfSpThoNvg8NQYTday9b5pj45+s1OGnXF3flBn
TwXz0h7iBq6jBz8gf5i+grjR/WEyH2dDQaBxdfKh2qYI7WYL3AZ31lRqZ5aglX91
envP2T6W16Aj7rCHVsUn/6qgJVA7hpTWb2847Fwat6RwB3UYaovZy9jrA0TM9haf
BO5J+oRV6FKW2BtIFglxcEjGX/3E2LkJujHLcdKqhQwPyYOBsFOnnW+fNPtyHOZV
/y6lUFaG25+ypez1FLtvNjrqVAtFD+45cGp7aOUpdBt5TwO083gXCjnBgmpwVTIy
giVlSdKxt05xT9efZp5fUbaFElWfaW6gXQFUePOHY3m6l5tTbySUIDbBp4i1pVsa
8g4pWdwac4am3Ezwu8WaGq6JAsyvcqio1g4nnIxFuNa3no7P2O+5BRW8f/F01nRl
wW2GbJOrobwXtlBomNuiIGWfdUfX80HIJdKmhKvrVii8alCLmXOVETl5m1PRtojm
as08/bspZadtw83QB/J1LkPGNNj/PJMZ8MiMj7xNHM08fxtiKQiXFs5cG8YGwGqJ
lm4DVMjZ1xJ9cnCBssErvbEdG2AIodStFCCEhxWHyVV33i64n6J7rtaNXq+tODNO
4t8RqOQV4NKj2w+nktTtaYuFCYiIkdyOYQJxg4gBbzYfX0ikstTe3YyAF1BFzO1M
oZouZC5qxBNsZyJSpbymCX/Bw9kP7TmSZx4Fd//j1b9OT9WzYD40aMRZg5BmUkFy
DFHJVD/XI0SRmJ3DAoiIC/zFjTUqG8FX5MIvJWs0vo60QlH9C5WQ8b514DyEF/lm
DFmL3Z8+dlt/VmgF3ILMroNBX9JQUxir//wd0mGbbqcNKW0CBNpa5bTWUj97hasK
T3HzS0gZKdZY8kybsaMRp7He8bOcpBwj+e+gRmZJqh5sp4oJ7Z6Yn3mPbumn9P+R
qnU3DTmPzv0UUNZhtcWy+7gfwmBenCGeDIDggkZ8I94idphN8ybD74Nl5Nup9Uaw
7CP08PypmwgpZNHqJCoZC16QJErJcalrFMq88/gK7iwtmjs4+HQjSagIf8lpZxTO
X8EufDPTxjfYOFhAstCo/0BBCBcKRKEGAkpaha4XF3QAJ/1kstKu3o/KhtQBzykq
4hwEhEO4YK0BYPI/7zdcEGpJD8m28gdWm12unNfBY7fCGdhHPuq9IDHKSp14U/jC
EhD90A9TOBsVxR7EJKNwDgKQCmR3BYQEQgCzSuSb31nIWQXZbnI/b00HyyQwv19I
nULcoWfSSzw7HsWI5X/trSH/zXp3QyQKiMooSsX0sRvP/6navO+qmCPRttFhEhig
Gn4K6wP8u4LBYVX16vlDdbJuf9JbNoBGeayFdIgTV+ara4s51sedSwNARAZEw7vb
nO6OPP0D9B0VGDQTc/OMVuQiSy7sHhwub5ejYNo9WC9A2t9rQVNkUsHDCpwE78vL
mHKbhzHw1RsEH/S1nfqmovy41kWy+1wIZpXAmkX2C8VNQ7WEi/kcH/5uYVH4IfLW
ruVzhPIvRQ8nvUOHWqA8YxBzy7R2fFLxIPhsnFGhxOoYzUJPuEx10mxLAldTmxYq
YLJFyTVV0HXuDEWKOSyaSGGGvmsx0k7sOkupRmBUVlQmGvPNfBH01LjGH/JT+Yhq
kNvryQzNG8r6KOGVC2RMfUEHfwsxazIDhpWIHMorHd4Os2EKuR704g0NAFY/32Nj
eI0UR0o/b3UGwR7TSXwYgvd26F+sTQVGD81CQXxnf/uWPieO0AsFA/XJYv385cu5
T7VIszow2IYBhCvCbT3Sul40+jgc0ZA4GRpdeBoHn/O9jyE9+9JSMzcqc2dBQFDC
ZYXf4G5UA/1mRkeKb22ycI0nv0h/q/Qrj5OYKgYkVe/r5EpvuyjwrP3pGB/f6bii
uKjxKdOMT79HbaW1/OQeTkxEiN9pa18E9Z6+xC5mNVKhXiwqsyBjjgWI0QfR8fZ6
mJEL5Hip5DqApF9qRzedBEc5q92ZfcF2w0JJ3xf0FKjQZD+vZYxL5ZPuvXud97QL
9xDxGtmQO+BXCakLmJe1u4sk93bCa2tV5oe1/83inNiRrQIqZlMw4G2e41LfWu1q
Xik79hoI6maVEvnTmdU+DHgn03c/kDn49FvwIQaBS/F6csrTYwetQYu24oaMvk89
FfUUBr2Pq6jDtAasWaX+5jS1UkSm9WNv1ZkSFZz5y80pmxpmRWHoVplLuHAbgfI7
zevmJq6h8DEIUQVVK6FD/KhKWmQOMiYGJAy+Xt5128p9/6pG+QnDnHvYD3FoaHkS
e1J0yfazlnd1TZYUdWbZ61sfOuC5L6GMurWVitUNYgnroLvlTj8djHHcsLN7RN62
Bv9uFcc4xTKjg3ksX8JesUr+Jlz95ye1zQAyKdq2sV1l7T5e88oyiCpNth1qnaxj
jOxa0VcxA37FnKpYLuBzc7/0VSVZufDPPzJ2ORNfQBAZlDzWGEpPIrtNvwEKIct+
TruE5Xt/+DsK+RogUXQ2Y41DlFWZiOHECw2tQqCZag9kXuibOOUZYXfYENV7oW9C
VZkK+H0shJ2z9Yi2QF3cthA31XgAz1ydspAOlL8Kpz8uIKf5dqqiFUAV1wCK9qr2
hQjnEdKlLUgxRF+uaOkc7zmahIF9ed6yJnHE6wxMHaV0cmL49wL4qbgfQ9C1y8Ir
zcMyX34P1xRSLvkdintpkMVPib/SmmqFOVR+pV4N85EgcyD+qz2G1kBBc/GAcIH3
9K3vyv6Q2bHY8trqsDxLM1oPTM6SlrXNj7SDvSMrkJQkhl+foXibKQuJ151XZjK9
1g0QU7lxKkyRmQe3mwDeEVI3yAGIH5GjWB6cSWSTeiEae1y4iyOEhGqbVF4ir9SD
71p5/pdb3Hd4x0RRj3KE7VHgPjfp1VnLKFDEI1LCZGRTbagCi+kZGE1CC3Od2LJg
QKxbyJN2Y5tlhPuH9gGOvLir2ojWmE3UO9o5A42LXK3Dd8DLD7j5MeWFbDdTJuEZ
TE7kaMOf9HdiV8caLN904adBOHugcL8lEOPxxa+M2Rz3pY/EtiTUEn8eaY8y7BEf
65pe7fJYUghxRvmfGXS8+boN0x1P7DSbctIJyIetTfB/SWGW8qs5S2pZ4AVjMGvm
eoXQf+nKzUNZAjWr4ZX6lMw5i4kdUCbNZZSMh8sFrjV/eL2CVklnz69uX2mwedoY
mbL28xsdeNPUIjpfrv+RLfdroL6UOUTeWbl5XWWJZGaMD6Vz+5kvu0FQu8obIq3o
vcP1BPk1Ee0YckIzfVW4lb72Bfh7mGwQoReiGKL2/CW1ggvMuA5xi7vYGI/gc4zr
0HFHE34KOUxNAsq9p07X9E1t1oFI+cTmt9U3uY3d+YIycRKA81rWl0hDl5JAOBZl
vxWnLVVkv3K5gbQ2qUIBMbC8COcUptRKUzbBhoI1W3ZeQ89AyTYjg/IebydayhgE
TTtljxQcuNpFgrFuJoGE7ZhPqj/kT8fmu/vNG9v5UwBQ+2NaAtMzf9Ug653Rpft6
o6jHDI8xPVC9GEt2o2F5F05IRS4pQNm7mg6mvg5Qn0JCN2V07SScuSbek4t6GhnO
K449SzNMwGYulZVlP+/vJ1Qnzt6jXTRL/ZT56j7VsnuecTVxRkJtPalRje/70nth
qFoKAbBr5QQO9YXDTZvbL91ei/ffBlNtpwMyyeSECAUT6j6LISB2qlSXpc8uoTGG
lI8TVgGx76zW9LTNi/CkSbnOqBNWjMl/GvViqO5tMdE8leUeFqG0wESA9m9/dLEv
Tqb95JBrWvCO0DNWToImU8CERC40Y+ROiGiBXj3yQDm6xYGCVmA04w5vpUAJUw4E
uMsY7BXgBFNuTkUw992mWeXyfCrxUJCh8SIBEvIsmtplo6UsbDn5eHzpPmwbzUkF
u4Er4WkjvW4DN/vXugnLT+zWug8srPWlMB9gdY63vfDOnbNRhRgCQ8gVi83Gu4kS
n+skx6KHsV8pJsH/hkIOEUlOZuizKbGKb95oY5IiajQow+CIojg5hKSGCbok+Bc6
ns0Lz0ayo6VfKQm7QbSzhD9Mo4gERGrofx1vKY+OdbRmux+xVU/i+K/5Nop/O1BJ
QeTOpLd/0MKf9CKNY9B3/zvqsBk/6d3kkgrRmfGJI1saybxDqlvc6ui4EEegLWRx
ueINYqBdZQIGr0qEtHIVGl9GXKO/69FFrBMoj9NJrNEOLXBtPaI6EGjL3mDD59i+
doJle/FkEwO3DxAH6yBA6SHxdpzEySeNQl8Pc/2moNvPGJEhcXDzERQMDAk8hrEv
HUfd/yfHcXjpE3jdL5g1tCfoBd0I5zvyM8Z/cTKKRSXH3bqeSA7nJLzMgqNRoC+A
R6pyZwa478v9lgoiLompX5obILSI+ajkuGOdqT+u+y6Yp5dydZykE8J+qG6/HoEO
JliqSdlmG6aqBC08FleFyOlsi8alSsump6rGIlzLp67MSrFK9plswaQTVSJa8Sae
Mj3YjeNaRRmEWC1R+7GRPBTtX3WvRCVbzwTlF0mVDvRWqJ51th+FFNecEm5CwVVj
BglBSOq10v6FFNhe08oltVF1DXMdL+xcXEUsUDI8IgdHn6d7qgozuMyxkFIkv5cU
MUQqP4IeulXUT8yuNgCgc8Kss0klHTFSO13f10S3+R+HDEiKLPG2QmCiB3HRjHWK
TfrtT6kSgF6ZXAeHpbKPWngD3asRoT5D+x4YOY9M8tQzNet127ItUjcv9SROEDtq
l8bhwXudlCjh/pisfgZtWdjBKVKezMTYHlEGUehUNRzT/qBgcwgGNpvPV4q+zDoW
JLyuJCOOAJwkWdIIWHlwfL7dWzzmUGx4yBIR1A03XkPdRqWk470vdJJbe7aK4ZC1
L/w3zFXE2QDmVktb6i2taZBLhuVHjS3thARGgTGzFoF8iBabmvvbOMimc2q8IEsF
ONrQEIDVQkx/qxmjYNMrZXD8nJ2TfC4ORPZ4CwrqlAUIOHYhiuqNalY0SyUpTI7p
cCVrOsK55vJ2ZsP55OoRaatVbdh0peyIlro+nHqhfsat6YkjGkLemYLxtVTUw8Fk
qAGkW2ovt6+9glOqF4S4sKPyptSzHLvIJMqC0/MHW9sjkqcgduTWCD1AsoVuSv9X
KMnqbd30uycjhtxyCOR+eMiZhB2iSSbqDJXdmvZZRefcjZhDbC2ichlPhJGukYOJ
iL61fpCl7E91f7416knWEkmgOr2kx23qmyRCdD7uWQ8H9sPklRLfMIJUNYIveIOe
ollbQB0UwpzDbcHKaXtRP2y4KBhdKW8XQHLgrX3SZ0z9OIXL3QEsJxohzO5l+nd1
yhfY4RTIQrsF0nAWVT2sx9s9MHA03h860TlxjZmmdXDIVHNAb14HcPRjWJbmuxPu
gpyM4Yx0j/UuLExCqowNBPaSdttZDaxHebM4MRvC2Er9TSFaMBLUBJI6Opv9RsOJ
L75rJCq/uOWFmkLaDIw4NE8NuvKMi9iGOt+lnw6BzZqRoCUdh1TU+zbWRuo/xVvP
yPG7NddOx4jeux/IUrH0l+EYeBQsM5qVXznc+mhfupMO3rO7rHNqX+j/epBBC3BR
RHWrJAFAifBNjBzXTIRe08yaWuWcGYvgIto1/cm8D2OPQ2QMxZdqcvIHh+1KjVjF
t5KlV8oDAqcm9sYlRKA2rAokYiRYtrINY2Dl1fbQseAuyjDyIrFH3nzAu6o+dnSG
VTkrS9Jsz621Fw2lyhtFQmVQqYpSuaiLeJrjFztEC8DwfCJkQApttSIZVXQqGal1
R2RN6pIAfmzjBoMCJhVcoH4QrA1+/OqUklo6eGJV8/zSPdn4z/TbfvTfuWYheqZ+
3SsWiBODFaqxyxuWj53xTjOm70a/KW0Zvx5agMpBiG2vhZCAa8MQdaT40oy74kcP
2qUokYJYwrtQHn12OPbJjtuThdVhkHOl0EleXQGI0GE8+efrbIZ4+dPEsf6S5GvQ
IJilqp0M2lPekUXRrkTJIqcCxFlk4e3YYIk3X3M9cqkWYqyd1RzGBv70CdIMRlj/
nf3v3l63yZaXgwM21QVSLDzuK5wcRyZCUMu7crQm11zoEE4jrlUo2bnFMq090JgS
tffPO5KYYsfJdo36aENBt2aZ0eZaKrfogC9e6536NV4tl/1qmL5i07JDToWsYoQ0
Kk070CjXtnTiGCmyLBsXzvUfOU71RD6lG0bsYddiKUYfRDuliZl9dZA1niEloJWy
pS3c22LphwlmKd3CMXpw09JV+wnL99oTjlILEciUK1rFwp+KpMGidAtaxfZMOBc/
S+pCm7MUISVXdOP4B86fRhMik3M79InyKsRYeYSujyRHbZPojz1q3HxFRMB2KA3V
MgnA0R3b2DvGe4R+qYFvVnrvE2CzcCTTwaavNvH9jFBSMdwTf4K1X8ZWKg7oLRYp
JjCr/S4OrvRg8dXi9hJjtKZYqZ+RN7GZSNrzX0PuJXoBcD5wayARNFFdhHwoC0Kh
HvlFkugSZx4Uz86ygYjHqNaydptfiYnb3uma6G7wS+AZjNs4U7xSGr2oKguOQUE0
3TXItkECKHvJ9HWDmi5v8P9sdcJl6+ThQ1nXWB+rhJMJ9efBPF/rYrf3b5Kdai8F
28r6B8fAH4eREWu6ydRC5KbCBqYZwQFTyHlmsO6vOM1IIYFlhUdAG/3MYzTdeaoK
rH34rLw7HRCuH/YJP/IrIZHEVV+MJHLykelZ0vDKIV+h98pIYwpOOGbUm0YekVYI
8B26W7jEC/Y8FH6ol8f+oJJUb7ZW3OC4a1UGiPF8xAZ2yf9Tir7YrfgUlTXuYcAH
ZZlUrNdKccCT0aSdQLDnnogNEddoRrq2VLGeDO3Oik10bhcS1lrmOKntBHTIR3qO
W163lbr5cL0QY835DV8Z0G5W5UROkvIq4suhFOYPsu9hTXvYEgOkh9yd+p+j5vnQ
q3yjrwyg/ONmavxXeTN7V4amQIe91oLYiXo8em/s4GNgvmtTtKcFdU/P5SJcF4hC
YUdvECSef0QDUUPAMZKqzcxeaib22coYBwDTC0eAKz2NPteQpoKu/bMz/WYqkXqm
3X2gQSlQzBDWnYYm5gVoH7x7meyyp+wrXMWWYXhfFbxOrS4CgVKt1RaoYSSNSI13
v0ABmiuIUaGfhafht60GPRLPtfdFyEXFtckCCXJ3P90tcBARtHpfvIbQ0yFNCCyu
xZy4cYc/tWgMgS/CXOctWhbsGA2+MBwHqbFibOYu7k6v3RS6juujJhSJ9MGuEKTt
FLamLDZ5Ixtn27bOXLpm8VcDj8Ll+7Yza3eGyeec9hZVO0cGfh1a2v2adg7CTLHy
WawfkgJikXULAIJ1pKXjGpv4sysOKruCDj7QyIoCEqAxnNN03wNom9lak90mA54Q
WoZ0ojeh4GZHHJ/O6aFLVCIUQC5r44LamgxRDcNQQnZw/UjCbPD9rgyTd3s04f88
RyiwcBbp6DpXI76guVU2qCFTYCWXs7vi3Tr1NxG9i7cLTSS+FkVuj6RC5QQwZMqK
rRirlhWZyykhaDnpkeALtbAoQGAlPXpEHUqBjMmpXtwPl28+1eS2jBW107CeAojt
3XSacjloOsP5SVqGr8Ut+mxihW+FbOGaRd1ZY+kbDcRmS/zEkeTlon9LoMW0irfP
AXa61MPy9QzHuMAYHRTkI5/xbqtJ0NK31R1402gwk4RiTcQu5AZNFIGrn0CWu7+n
aL46UjA0BNgg8DLv2b1lUTWgYe2fw17bo8qjtjyVB7F7iwB5hwrmWOxlh+gD1aW2
FujBPPunXuxc3nRgIqQGfA5lVtrtQlBNUL3Iii7HCEYn7/V8yiDANm7krRvpdJvR
2tyeq58WMzO6oTkBslCuaD8c7ZTw0pOI2KQWkxA0hf7v9B7gz3I0VqKotTJUv8tY
fMl9+vQLTc4kp7yJ0MdE24MBSzcSFoVxS9LFVMp8Q7epnKmeQt0zURLYPtCcC4va
nMmeozs8TZO51MQdv2DPcjmAvoD05Ch0QZlhwGsf1gxsoSOTIRHoN+HHqonLZvrg
yq2bEQSLdYybh3tGF3dlcneWvrcQUgEQ31ofzboskBj2HQYRLEBEF5Yv35RNYob3
KVVPNWw791WLL1Qg/AfjUIGXqBFYKGLICzglZF0zX/A0InIgHNSUb92xJoZT9CZ3
w2PcEOtUYQ27DMvCnj7sCflZNBm8QER90xlGN4RHNYJf1d0iaf+cplWIEos6mbEL
Q5Glwukse/Xxfg3Ve30CoGrRgb9aNb5ygGWxX1It1jo1qnPNX451xF2vCzfiEuv9
eXR13MC/6+jIFis4tL+fcc5ncHAAssirJMTfhJUf2XEQcstiZD037bZhhBnjidm2
GGQFGz2GmhNxv/XQST0R5e7tWbwxGbiWbWhJLsThvee4wx00upRusX3wGngjHe2x
jP++QqR4vH+b9LjR3x/6FQcoh0VJX9CP5LlP5fzz3/U1bPp2qCM1ixMBEQMoYWcP
8SPj5qDD16i8NuAMjEcqW8vK08MRsOdeOlMUiz5xsqDR05wmK9c2i931f3JWrBij
LNb3GzrnrG0a3pGXBoGXK1jesKq8akJsA9swX/8RF2FU4wwfGT+Ci/Gl4iBLz9Ez
sEgrvct9N1JbXu3Z0K2Rq6tIoHIVs2vDzZ2KgRRuTGBkm2BIkO/akmmKpicegDPG
Yzr0tA1Ux/waKmQpIbDSI2XEuaX/f3DAenQCr8ncFQ4iRP8OAnYnIBVq62hOYNGe
IufbUj3hmS0sR26QglFNQROjNoI6czNNp1awLvLUVZ8BjRrkn586kmzv9LTlts1Z
4OuLiUIdCtwL16BFHUIGFBQ1WqxtrdWieGnNmsdQBQ21FtsCFVHO69WLOtsBq6Mh
1iPKKlcVQZc6n5+mTXWNQ5whNK+/KzPC+CgpPw/iHuPd1zHrrzQ0BkC87Qnd4rcE
7zMkoRdRVk0lCAiSIX3NJhAIEKuJhqEvpgmOXZhMiIkjo2x1WP8dvKtnMY8POVbU
RjIkTSsyJUV2Uaizp79sjZiu2W/w0zafr0Kyf4VwJiY4RZUBqgAD+PIaUkODtLhf
d31nJCoNlgqkqeRKZz5qxVFmFHKO2LXAy61dWn/9y8yDHJElmAf4pJzLk1vX7ZOA
NbUfXM9czFCF91mjqWp9kea4c8bkvYHKutu3JMPktmVX6RrZ5/ACjKzxoVrk4W3N
79BCRsP8tr9QeWMjmuvom8ZU6veunMpsCQZIxL/MIM8BZxdXXo8WnaI4S3Yb89kV
KrU0IchA5cBgeLz7TVO1aGY72JzQrqTqRu4ycgPTTSz1y4sg82yo8SregZDp2z5t
TOzOs2URsog5WIqnrVSpv/svc/8tGQu8H4u3pzjFbdPRuCh5nO/h4cIaIQZBSBPC
/cuL61idUA9xHUTugS5XJGCYEqNNT7mHWcNK3q/5bq+oYEBa2ohcarUyGINK4fUK
W1RK5ba0LwhIPCo77v4YqLKOB4Uvdkfm4VTXOE3OJA3LfEBKf59Y+Ot/GEAdIuM7
+JtzyAMfxVHdlhv30BWFKdDeMacDcKTQrFbMXApxhopwHHJnWJsIoAmzbvBFmWAA
8d+ul93sM8KOlrERNANmUH5FWudtFGp5D4nNdBnglZ54EME119SXK/b3E3taaWLy
yMpREgZ+PEOTTrHwy1V2AJbn48ePywmcxaPlHFkCcKGrSPNfisFklaYNjiJU5MJL
nmaw56H3JEmjJRk+0eDSMSvFptmIXSnzxA415X/YIi7vDXk4ZWbhjcz16cMS+QyP
pTrHIEUSkv0jwsaEYpyLGyZWROOnsVeRlQ4E2ceeH1SMZp1dA2tJXKqUHBYnAyjJ
c0xHXsPDvJ51RKnvNlmq735S1nB5eHi02OcEabMpAtD8+vadBviUIcaIzLZdf4RY
xTnNEPYgpR45BopX6tct+rr4TYAuQb4qNsKIuDamg6+prcCJ9OJ/yOXZ8i4A1OL2
6UI3ogeOdlMKu1XfannPfflwMwbd27LsqI4qz2cP1/smbu8Qwsr27Smyrojctgw9
weJogIC1D6EvXp+H0U0TuRuEJ7Es7XlkmDliD0lHhQ7uz5Y5hRwsLlfGi3193DcX
sUF3FUCmIdS85Tf3nK/txgRPvMB+iBQSZJJ7R7OY6LX1wqE8UGr7eB5kheU18HZ4
3QZVVM80zp3QmUPpb4IqxuR/cXJgbRb65FiEBCnLbEWGncWOxyuRmB+QbihdYCqJ
UOSHDuIhNFQpZh/XsS7IhwtyzxBRSyZmKrYM9UFP/hkIyPEyPUGKA0p9A0+Na7xY
4aQ+9vlTex/ZvVSx2Ynrblu2YPRR/9kNAajMjE9SvZsFCRPJqgnLFpFgJ0sB8lo7
V2SLI6eaBFhNe2VauecthNz38J1Fo2xMqBX0GM6uxQwaFYkC+k3C+QUYYGBIMl65
O+BsKXbH7PDL5QM8y7tiATuo3X8wLvBu2dsM3PPKQBwqmDvwqiGSH3ZUiMkHOl1x
ykJprbWpe/Vg06oHL3FxUOtCyqqNs37hgBGByeo1T+Inv/S0qfHLY0EQHAQoTNVx
PsaEj8ud3huqOflOhzOqwjO7nh3w/N1m37hb3Sgg3hqdhZmr+zTad1kQT5yIuZZC
k0dejhzdck43M2Bf5WiJUngLixmm7JHiELL/xggdkJL12UMUt7bLpCy7rZ76TlIM
wpuzebceTuqSWqkYCkUd73c5aNw0hcD7fS2Uf0a1nttL2RRSlqxvm9WAvKtp9d6M
HMG//J7/aoy5EeItg0BnuQFkKwSbT9OQnrDfH0nVY4Fa8ZqXew5iGtuBeZTskrf3
PuzfgSB+Dz1Sw2NnUxx2h98mliKrrHdyezEg4jFkG0Q5gemrF1qcBZPpnyAt14bh
rq8Rdmis4dKkgJjw9oTTDDMoFShX5p6DAOy0XFjl6fHPWJM8mfA3ns3BJzTLgses
YRz9aTl7XmBhg9x4//nH/1LUJUDmYRRSYVzhNOB2Hxd0Q7XErSIyor8AQP0Ubtfg
m15lj4+wWiQmooAVmQF50KcLxisuM3HTVwO6AScDlb28JcwKVG4zSwwQ2Pa6RLJn
EhGBlEC5YpneAfogeSlAOJRqeDMELVlyOLodxWo4ArtHM0wPkaZdDkKd8v5ZIgff
h43qn/HfeGEHLukdcpGOXdHGFAaI3S7LazQLsvIiBzLyPNqKLgRIP18A4yxYPvFx
itUAlQA/8e+AYFY2QsRARGsIOnX9xDw+jRQbFDsthJnoLeiwUfhcqh+byyMq+nec
C197pjRKFn1yKDNrhfIiRHWV7ScjEfRhPKb/OwCprJlCw1Xu3WZiagtm6C7ttEiJ
aoSiFhWKByszP9anESu4RdUUfreVLTbAALf2h1qIg8Wv/MipwSXDizmqQX36olyM
TBskgI/7AsUXvGINiCRJN+4nCrat6Fzugh+n1EQWHj3W28EQnS2TmMKo8RPg/3+v
M+luKMjGj1gXQ+rwrEsu3mnoFYnfWgu0nEiNsv+/YRVGbl1OnambN2EO8c+ocADl
Qehl1gybFxV9PlJnXyz9X6xV5Bb+7gjjL/hmYZAoyWOScPvAMafJakSFkRDyItsQ
Zy5gKFoQdd0YQsKX3GTyJWW4VJRXTnlMrgDcTa6PV/J0WW65zBbThmMsp4pKbkFE
XP2lmOrD7ALn6cdQjcyAKTiAyv8HagRPTf4WXn4A5Ws8DCsSSWhY9Hn2xVDAoxwF
z1LEAnzhF3H4Npt/mCKWvGbMhZtU44vwNdq66btE7uy4cwqHDgqnbPzluuf7pvpj
xmlJaQauiXFZllTl1aZ4YmLnU2blV33mmFTlPND+Y9vQDV82Xt1rdKNj8am0725u
V/CI2F3CgQ4SmdPr56qH87PNHSRo10XT0FT/LwfFGtoKRmmwlCk5AUCIgU4JqCH8
aSAEp/v8Xb0cnfKrbryLZrJqWKadyMT+2ShvpNvs4T9n4ozNm0n+2LVOsNR36yU5
DMWjbiLY714c913RO0RfzXEfLr1quMoigzrFoSZgBSHYfF4l0sc5lNk4diMoWeg3
hqTL3Lay6GJk1J3npyajjw2NayK787+9trIsacx6XBHDy1eI+6Zxx9aVl6+fcdcD
DrVuJDb8sCIdKX5Tu4KhlR8TggB0qIYM0TqLjwYldSlzFWwpddzfMzxd0BSkdb1/
A4X42HXwBc4QB2Li6EyjYNy6TvU9fz6nlD956b6Xp+7OvbjOVg2lSEEQ9VfQv8wY
Z33x/TteeGTP79tabFy7nKiIFDb5p/j2FG7PeK9z9t4xUbCxsryO0SbllsAzFSpo
GH5JEXkS0t6eNaTrJXTgldT4D5z1ZyGM57MwqowYqTTktyeju9TAlPcEyfxtg5xq
Wvma0Ks11PzyS6vNjfO56dtnQYKpl1mpgBxMN2ovIsk+E03Ok6J1ojHD8K2p7oQU
1WjbLVoGXO4zkT6np1tS+LNIBJOf3FYiviA2+KsGtVeCBFtMtv7JI5dBNX/rK9+P
JcyvELcKKZzy6/qr1LGuRJE8AwcfgAJP2HshaBXVMXN/fFjONJ4MZgdSCgrR84Ks
zlXLSrwFmN4LhvFrR5VaV/Z/Jhj8fir6KAeEQBOZLnI8wce3dRmJ5fe1ppx5wxXZ
wOZsF14IvWP3DeX+52q/9nKVH+IQzhjAvLvKEjyaP/mNlh2O5CkszGiRfIYeugWb
I20CdQXTZCRl58MPz8941MycJJUw8pwUtwnayrintOXFECsRbN3rdnvxCUiN0D/O
uadyOTOVvZSPTEfsshr4i/+48xKNCJ8/cHlNpvWzuVHdqjkhLHdF8fM9fmKTb/zJ
j0LSVi+yWPLctdMT7GuopLyKzGfrgQyRrys+k4PMAPHJGnTSaarWk8W/UA/mdsil
ho5rYtXEIDiceJN+6TR62XtrmbUdC0bIpt/1ILrjGstWB/jBFl8LBKeODjBS0lh7
PAyMWb0nbchjRea0BJepZAn8VrrOu8pCpdb5X6/awcLH07M3Di594LkwBDMtlx9A
K8vhdufofOFuxRvpfuhYOVwhMeE7h5PuHoFEmeJjzRGpAGMkqIMdDDumq8Ur/+Wo
X/dri475Rp5tlW2+fIvfVzHxuatnRavHOzUXFy769gD5QLebj09wcQGPly3HMFcP
jJT74QTw8A5EP3Akrq/X0X/srLVQZ16MwG2V4O+mv7C17T8Tn5ecFANhlsJrt7vK
HXFU89qH5m2rY3rhINOpl6hq95epigCj2wd8PmYCtpAGxR0znNwk1fjDTqqAYwAR
HC0c9vzeIqP0UeWdwVxvhUo0UqXIThkEMFtDZtanbvDl233ENwmWTKNM1IGCPWo9
2/tsgcqGQfc9mMQvasXN1ZoAv4cF3L2WZNfRr3l9WShBVhkaWpCTxBiw4quNMq0K
ICbGuAMCufLcYzY/FAvSSODHmlVyWreBL2HHz6uUdn6/f+NEMhin0ypSa2AAEm8V
NovDRwn0TMGjgeYBnTjFP7mZ6saE9RHB8+6QTW/CfsgFeIRLoyqmZoR7U8y+mLjg
DP89I9BvZ4v4y4nktRanF2uKme/fGdvRf+Hs4gN6EsGnEcU/Yf1/oVE2omCBLVrz
BSSXhHot6v3KCZKW8itR0dscyvVKjHFBQORE+DKFdYYzawLFwXKYt5ssEqDL8eSV
VC0YbSzW85a4fXRQbbYD8lfAngj0Hbf5N2KPHGhY6dIoC+7DloSR7luXCJLePSH8
w06wRoz6Iw1MJXnWnU4MnRUlnkPGJIvagYwOQQYlJVsU1MR2IHfndQCU8nnAd1/n
zYmIbZVEOZ4hPSfZbkVmH3pSKo1D8/2u3Q7dIMLbFh6z4sGripKERTSarP9PFEdp
F80FOLfm/IG/m7tcmhGZLyFvqpp/Obfp5Sd8SvOdBDMPwKuz2DAInOmipDZ59L4v
5ahRK4TeOO/m+vOdxTeQBla3I12lu7+b41zV36t5/A9WIhzcRmMqClP103Zs5D5o
MLSNc+bMzxayFn8zBgf2Kzv/Df7b6gmIo+5k9Pva8w1HFmwzVE78b5GrPKd4Z1HU
Qqc+u+RSQ3wx6MaSxf17/HAV/XyoNdAFm2Vw7DbRkBRexafe5tKXOAjyxcrOR0hg
BnDw7jTUBBtj1pNHxkvqK8RTKRNfKNH656lRuMLQzgLhUoE34fBsakPznTVVf5tD
9h2v9yRnAtNUDkTsDS1HNt/oJDnGHRL0RyjZZ57vsaOmv0vYjcYdYhCLBvguNPhs
b9Mi/bj3iDrxNp8iLYw9skbi5uKvbQdZrrhctmz71s2WoVkgqLCZ5xUnPwBSGuNS
ibLM7quwFgc1FvnfNaYzWvKdhpvfBZI0oyLb4NahBBOtFHOov06fu2XHbdJ3P8I1
HlQJhpnNumU9kM/9y3COEeDXFt9boCLxlXSFvbcFnhnVzDxHbaQk6bxdpZ/9RLsn
7HiZQBHftsN25GwLxAwMPZKmCGXkZhkEJNPOeT2ONq79Mvh3ExeZm+AVpoQFZw/R
D+41UEzsFN2hlKDEcmWwAx+YQ5Vm7QRg0tEXOGEm27IniMhtPuZdUqj3V7cE3fL5
gMv4H4dDuS//0E2FsUu8B2Ldmox/pXm//NgvqGlH4BtdzxEg8tauiOUPZpaIOBEL
LBWNKdWFEHqL3HR2UYEArxhOSiFxfjGwRuzs8WI9arbaw4NMufNRV6TmAk5IrJRt
xRj/Y1YN/NwqUIJhmYj3ebhqBjj+JRbn8bHXlRrVI/vlj1BpS/1qEK5GDLcefkws
K92MFSeP+1LsY846OvuKW0CYEVJ9BmAiGPxEwhcATH0EuCHXGjfZNIoknZ0AwSrT
kdZiNI57NUCcdah6xQGE6ohLIuq3fJn82LabwyFOnFDy63IoiaRkL0p0Kdprol1q
OmS2BjusrNke3JVcpkHN67xUsIAY+mtS8xz10oyNAKyeXsB5OX+CzQPXlV0LjVZN
8Ojx06upCAMgCG56yEYOAvmyZ0isJrXY9tJXszZ8wsXZE3C3t8Adh4l2DM6mDPzT
Kfek6BiL3yAQH9YpLkXAXrTYGwWSYY9IF2j65+5/uHLH0gcjK1g9J/gLUT5SvycW
mAjnyU9sn9t/kZoRxzcQms8YMEdDSpIbZ3rpJnll6w0FECMC/FF9okOHrUEDgpIL
c8E6ETOHn6j3PDDV/ZCUl/wHGhdBglR0Iqcf0NlqZUkdX8nFfGyC+WJgO7/GJZSR
SN+sr7WruBHzaYoiKQz+Df0Y3aFYKK26iZcUve8XvpmdmarJmNc5Lrezoq8oKiT/
Zx13g1o8bTMoX8RUTDkzU/un+e2atSUAGIQxI+rfQzuPltJxeUVSoNWpu0/jcHQQ
Y76iZCGTdK4s5Qbl/72qHaDMALPUaWy6qMb7lMKRdicTW0dURc93HAmaq1hxFFdK
fyuDj5Ezkl63dNglegZET9ml6e5yHjrKBLahbWAzbhke8+IXcx2TtDFhxWkV69cn
uhbDYklfW9eQsjzDVhkjh7VazN2jjVYXIBiwpqs+DillH3xpjgFqQN/4bpBhkg7n
L2t1gZgHVK4gkNonzZBmMKSHyWaSMu82gPKAyLZIwuCUQiuxosmC46tuCFxp0raC
z99eG9kuX3679mMPxHii0eSMv3SLiS0EyAdqbocHzwIo4/1dnSTOB+uHM/5Yjogv
xU9FuK8QL9BbDAVphfShoZGjaJ+DmCRepjDfEEV1Zf6YT6zKdl8d9ud8urjTuD3D
HlTVLyLsvqBjR2IurJp5rLNf4XStfurFbUGiJbXU1y9up08NlDdzF2ZYYpg+AYMq
xW++y8pg3FVm3zQsF7OBFe2+AsI49K/lRYqDWXkwocbe+DNACdZ8xSst9xbLaEVc
c2A1euszrqpQ4jMKA4C376ytI0DP4n3JAMw89jjYmniulo/yjwvtks/ZvyK8VNQM
1Y/MnnWWxTlF3a3Am1gKphjAmstYAEJzHSGD/0T37iAPMi/YQUF9VjZ8WgROCJO8
PNQlXsL50crB6QYPFU0Cn1SnpdYPLgR50Wv2L2zPSoO7xAHE07BES49ZmgL/tno1
nhxLKE1+rWqsIEs0GTVY+XrU/rlbLsNf/xwbpQXaGaD9kiWpSDYmZfhmB528QM7a
scI+poo6v/Odzxm/eKmEUffdDaO/h/mtF/PoLS2pnjUP3akWTEHEqUDz4tjZ/aRs
7mAeU5L0Nf6Zle7qVtDiJZPgKNO6/rb6oOIuE7V/XsltfFpyNess+EeywKA7xuWi
9ukm9AQ+K4ALbx4An4cBHoyjBVhgPIYGe4QIIoLEOshhp/s7DWWybFoLp7reC6Oi
LONI041yo4nbDMyxtvy1hYanRH13teDYiOF4yivM0UCfKkY1/1XbxuaZ+K8X1Drw
lQsl7bmqf/NQfYS2wHdo2Vqi+In00L6can+p1qkKxg6zOgzcjyZv5tg6iXtmAbKA
kUVOloc/lNjx5jQV0TwVv8c0WyJktjd1AZNkA/QkDgWQPw7XLR7xh2etGDhChTmZ
1KQoohbZotONeoXtOXKx2mUnwcbiHjjqII1A5OIWzJD9zjOFpDEAoyAhUFYUBT/G
VzmoKH66WILbUrDt01JJnBAfVRnXDBedTo4EAMzwAOIZCRD31IUHE1T9GM1He9JR
Nft1/lsrwNJNsudhRDjYDyQBbGsIf3C0NpvIrEifiI5b3rxKUZDdWqvPeZU9f5pf
cy9/Jh707lcEfhCi6JvQefv1tb2b0RBLWDsRPgU7BiccACgQuVQo0BgRbYLSdllZ
VMHl2yIREsVkLZ5OoptP80lqgcE3s2GeTvt1AM2wk3D0Mjc8N74N9ch3ByaEJjr2
6A6odwf0rXFBk232eKoMeFcW7B9DclwnLnQ2Nz7EoDuaoio30a1XP+salZy0BUcr
oHsDGzhwhZTUBKgILv0r6CVqCFMjW4O4mM5RFX7oBjaOuiXvycvb1WOqGARncThe
O2Bb3RErnXw52I12IVEUjob/l4aUopmhMDMGFZaXiRN/jYEe8mK63Y/jxMEnmJXR
dZGyLHhU1ASiOP0+8mGXxnh7rY5K4qaMxzAfSPmFFevQPUX4JIcfz9D2vZOeg1RQ
Awu9hzbRcEY52911Ye5asRdIWZPxKK1Bc5MdW+v69Fd2PwZfR4wmHwqhfne1STwK
Nqq2LGfHlZ+Tm+LA8NJnl21ma+w2ir12lG+UHYBZd3b7i9cOh7JLJe4aLL7c93Bo
AyHtM8a8POiJ+Arq+9d4waou+RKeexaip20Vt1EWjH4qkKInaKmPcM5+SS/DBhgd
alCOLJ7LYRpMOgIs7gxm9CC7zrLJ6ZgVfkqGgxg1uxKjwP4w92IwvmJfmCoEMlkZ
kc3EiVnV3bOwPUuVtd3rnqVyhi9HTk5fK3Rr4Ae2a9AuNn/V6mETc3n8rg+/2Bbz
ymBB1eWob7Q9x0goANSbpwmc5BBXX8onYvBOMYGUFalEmByssa2mEiEuCkBjZO63
1W85NEHG+Bm5Pj679r85PmVPzRw9s2isKvbcnymBe3gcQOLeVseny76YBOJh2wFs
Dgvm8oykoq3zLJ7xH8u7nUlz0lJqHgneV7KGOVqllqV71ntXKKfh0Mj8ptW/PK7j
jc7IGwZRSwJsbgmeJOpKpRqkeeeH6tSj9H6APlE3LhIyH3+66RAp6HJxli8VnJGp
w1P7U+aBBb0ZEmdGRXzJgTXACpLbT+x9SBmSRbYP/Othdvc/SAwGm58GW0yn2mi7
fkZrGmsEJAXpdMti0aCZlqcEi78aVWI4iMnrjXQVhU81FxJdaZfUakyMkxtOoysk
A04iiwyJJoOVrz8ZRdRKaEvp3wvqj6Iu2xFMRhFYP6q4U6WC/8y/5XV4DyiwTzwM
SgcGMmhNFI/T/q3pKWm1Ofl4iiKcy7W+LXL08cDezw2PUWaYfAM+lIJRd2vIxC0S
dL3iqpV/P20Fw/G+0fYlh8ipGqzln7h2uCDz/cY0K/CgDINT4pyI4O2YAdHIf2ec
hPHjadw18ZYQKtSZ+fHQYC3fbukflwazWgTWohqAd2gZNFVDtEBNnT89I45LAnHv
jJE3z3HNhCK5RNsCLFQ4KOuP8yFUJPlhAR+WxO7TuVi/b/bIjOBkGXZs39hxrww6
/W2KOSSbDj9eB7eI35KnoqXeuuf1quSgQdKfnTo7cIVLgP5x9r3RVU/TO8jY8Tmi
BwG3XwgVvFAqr7ssfZFRxKo+31p+16TFvB1lwsYr6iWNj+CZ0DmkHOzpY4WwxO19
+/ZLlbInFMiY66b2upZ21cKvup0uZto+kPu3cNy/MAoPUDzBqOhJybFA2xVtz1jm
I0NGm5joDLLctRzYPUX2fEcBr3m0zeHef55hIhoyf9I+9MoezYUHoSCs189q7b1z
xtKtNkJ47MpyK6GOutOTTadBR3Sn0aQ6MpnBpUEQelgog+qVFRs4b6muhTlHeZhb
IC7A1z5ohSXeo4aS4P8diDlh/nggoH9gfn+5Fya3a3nD55DSUJUXxa7PCucZiw2T
u44aEXy0ep6zOYr6Or0DFa3oe/Y4k3UogwaupEuFKVLkONPYQ1xcJoko47KF10H4
dkpUob0wuiHluxY+f4wOSosZDOjRpj5bvhxGad891Bk5UMDR4vmr8b124+Kr28O4
J1hOopgOMfdLWv2o/37eP+tOpcucEo0fX/3mqu85NKTgueX1FLtlOLKUqjg9K5v7
oIU9m1iHpFzURc/YMfBg+wHWCcQgh6unnu9fVBvV+bnd+s+0PMRJKJpsrde6JJdm
1a+wKugsQFpe2gb/vYHUpYcH2n0ya+Mo9IQJY1bQukSOjzS48cvU9deqpaxL+ot/
h7cQZxFuXoqgDLGsRxJDjTSOvT+S/xFnAM2L9w6wYSyWHHj5z0CRTA2XtHX9MHSj
+/+1aaPrg6Tw5GexO6D1fIY8efMC7/kijjTvsAJj93Ms2jwqek4R1Z8LRHC5EDgQ
4iXqKepNQ/CueHQc7bxXd871deZVdWKaABq0MvJFtoOluJqma9BknC+LQAKz9Xu+
SpprBbBMPj+xzDZdCaHP9+Dcjm/71DC7kXl9FbvlXhALcNfVKxnMK7b2ks7FlG6k
rvDnGl2iGAZaAxSqp90OwtAiY8MeN91TRCcdUbX/Qqdtgyb5VjAL+QycF5+VZFif
PIidQgEA/hTHBLSujmzo4CDpdRoMUuYg74/U5cISIy8n9pEyU/l5NgXCYHHj4Z2r
66lxBhxwrSw1ETOFKMlCYeE8m3HzAVP3Fixj2Gd61yIBUED9NontepU+AO8GdoqF
+jVMaIB4x8XEdJCCr2NkTMg1+QrZEDgZ+lLHf1rXnrBvKQPOzxxrKjLGSknX0ViU
qgzeLkD6blPaI3U8MwK8NP+HDwTwUPwuQFxFYW+tF7JpZh2ub8j51nMpYiTNyjAs
2shrtyyT20VQa7bVa9t5enHwMtoKrkJy/xd/sTtc3dGKMvnI3VbXv45kPiPjVR9V
RM2WQxzUWmWhFu7xDj4+2oBbtqYETOkT+PsT01eXrR/wXzgtl2hn8yacPEMEv3GI
5I1RgDAh43Xb8NFs1y8FqmJoMOXok0AJpbwin0+5oCNCaO4ml462OAIB+oS/20si
4L6KEpMoFHu2Zz0Fz/TH6UAL7PCeOWVXFOFLtrU/51tmHPMVLN50w+9Ov2Zfun/h
mqrRrEp3ZnL25SVkVkAWBs+vJPAPbMO5Sukq5Vj5Ya43bltg7/rH7cLYbdoHS3Vz
NaFLORtEpJYgbnNKsgquLaxgRru1P4BcJMWn0DVQDSvngJxE8SSJXG+dPY9K+7E+
dwDrExpLnw8o4J3QwMHevot7iUxEF11anYEnQAbifa2QxOQ0KPM0DSURIRTLuPQ9
2dIrSiDyrWFbBYClj/FX4NxDn3M8rJBlKV6HP90Q/hKovpJ78JePIs34zHTHjtqm
p0EACig5YshsLPwc1roa1TPvrpwXXP8GkahUdNSGsDS4jQb3gluDM21ng4vV5FWi
qKf4i9Y0O0xqqYPhL2+k7LX/KRSfVfLWat8ztz8RUODedjJvNOHf9yUiRuQ2HCGx
2ZS/erDNqZIokO++AXoQmg0pPNqian8YWuDyUQgRzYL5/rf762C1AUNHzpi+XaeN
lbcTiNgt4Qf1M6afb9LSO3K+/xa4GqxXrq2WGZLaPZsm4zW5B6E5230cMhQTb3qJ
HU43LBmsIBy9doQBu4wv2ZV+jNBoplm13Iw5Or8uxZKDLqVGthbJXDIWnH0Ijtdf
ZU6vkSHcsLCoibJdpYV8m5HUorLjnJihUrmzShAtGZhaJUjFDWM3SAryJ6w8Kq9F
r28Ndr5msHQ9BBEAIBleTjE3Hrh7d98HzBl+kK7YoafdvjkQUkeA9kqdOor2PnDK
EJnX4pX7YeghSQNTrxqH9BbEnRyvrkb5EA0l1cHrmNkTGgBfoRLhY3nERf5rXLAg
jPDbFqFEkOXI4m3TGGcOjpETAl9bHVcfTp47Fj8F68OeJ402Vh4zqY9v9hq6qgbt
wY7wCc/RNsVMBjLMSjwN/L3HMfJFuDARVefDinMK0G7VVd1fd447NoHTZ7X+OKoy
t3pYz44vIME4Cal+mJABlXKRLDsyXgCEqahq1emz36Wfk8qIiUPly7ulzvxPwgTh
R2BOmklH+a0TaEzG4IneiJpIZ5pIv8KAfyTnWuDoWMW9fFRr+wMMq4Gr7HfY05k1
hY6ypP5dRLrmrLe/09B9/8GDppyENJ5E6HiTy4H0Vfhop0xgW9wZtwrrTTROLkSt
w12wLWlTB3tnTF1DI1zA/xvM6q3cHiI67oxYXQHFJ/0SKcHH7tenumyJJxLAHeR1
1rlhNngelrxPHWfFvC184xBsWXBLAAYfga8puPsjGHWLWliBIQFsEVpAxPf4vQiI
DJ5VKHIKAhv2HKaupW1qcpbhcaW1jDKFqkMOCy2tpaNvk30WIu7E2XKOWcz4gW+g
UV0EMZTCdtRkIweVN/FBg8i5JcZwIY1CytRBbD39N8vVDgdkZ9V2rcxxRJSxlSLe
32b0DQzRzAGLFF1zBZH3bnVqqIS08ueqALBZdOP85TygtExnXr+963ageSxmKsjp
ITkTb8QCTzCSXXcz01zWwxY79qU7RphU4diutrtIk9pRF6vW0J1Njsl8EBXD5unz
maKsTCp6H8tL/RisgFPyKEhZMSjngQsFKTh/Cll1wA10jlNly/d/ABIli9uu1Ey2
94w4t2uyhXLWiOFxKrXfCJvP0LS9j7BeEVLMz66iW7jauMltcnIq2A+0aIBRBFu0
LmAbLrcy5KznIlsjyih43/PpGf01X0cDXiuk0XLdkuEZW6XyjJHUNv7My6GiV8UC
8R4Url4pcJ7SO8RhVd4ObnReuZeakKUyPg/SEh4//sE38rpdH/AxWXkR8FtZNpg2
hMU5x8exOdbZ5g2qpduIoPR53JM+DN9M7s4os22jczaBE9PIvlGt0XawqpF41HgG
8eDR7vo3akMkdIjkcw/bPvFuUif89Yot6UnsGhj54PisdoqJ3UzeD7EzOI/hshAD
y3IJeyB5LEc9frWCpvPQxDLD7AwErDslS88vma9xTytfIjeBrs5bem12MOOy8YAN
e+O9aw1QFcgA02KklELoRQXE0/yTqUPNXqZcFbDLWUihKXYAcaNrLdxKkxYPzpCr
iBDCZ9w8pY5PFmJZeNVDOZi1XQqW/Ly0QMXoUvH4+XTBwzw8h17gJ4ATULkmRwVR
Pedmebw4eDzo3HA+IC5wcoUONTBE9G2OwIk7E631GBaSJ8ot2QbQPb3/GauJVqng
qcGaiIRJLqUIj3kIzcH8UiPruEfI7cjhoFIoaT7QWRPgCMRMRqwJAswMWb02Rs/7
3J851AH9p+HJgZjgFOJjKNawMQQ5oyc9zWT1lssPjhm5LhuM2WGCm+bFUhm0SvEg
Db/5A+dVRlnLFFC5QqqxCDT3Dn5p5Vjd5ysEczmCRlfIaEnXZI6xzMQSUikpgLRP
v7Db4RQCygs9qRQqWpzm9yP8VpOpaKyl+6IBdm3Dq7TUVJwMSBEpLkcRJirHl6LG
AJxj/fPChKnfId495bL5BPLlj8Xpy9q08zuQKaWzB5lQzrmtr/WMHLaTNx+WjBD5
aNoOHV0PImR9MvEwFf5FUw5ruxh19swgXZycIQ+YScCa/71r+8SHWTio4K6NrLY4
N3tkaPy3npXm3VOneRIyKfSdfHgNuYEOwA0//it3WrDh2b93vCUHp+QyWzOiW+MA
ufUZh7LYC/1lgBILuF0Rq1xpbbidm4ZXTwxRSqEGViRLdwtGt8u7i52xMq6FKzZL
ssvDn95PQbl64e8QY+awquHw9U2C3RYgGQPbsmDI/9rm3otWfudxovcDsGVVNqVT
4C/IGTSEiqrOnJvnOdOBef6ndhGGho4u87Ns8ivnYL5Z2hOTh+RwAiAJrvNTsxgx
lL9PgTmJogMjpoKgpBXk9vtpL3ucbm0xGkMkMGN+x9vZzXHk/bTH3pQLBVqqzh8R
IS4MDenS8YLfGg8ram9fpuFDsk4iKdpMsrtAqKYGgleC/7W/QsnKVsMRR0QL5FPn
bZ/mhDZ069UniVud7z9pvmeipYwQBUJ4wtCiog4RnKPMq20yqFVKRv/ZVVmwFr1w
bk1YWelK4qyrBSX52MqqT7JaThDc5M2OC89ZM1DpgDWeaSHm3t6OgGLeiRPr2PI0
Spat23Mc3absZl07odkyJTQ1K8hmgfiB2dazANJYTAcbpw9/+rzYY6xhTRMYTPyx
X+pLZYfUhJxr3TyHzQfVhkCenBJQUphOEmZPCapdZZc+O/ymFMa+Mk8l4bjs4qn8
eNal8JSduF1xwoj9MfPENN3WCfUpyWWJUMR85iSx4ms5d2qjwVxKGDgbbQdbZO+K
1eax8I5y9i5IC/bqlS6q3ty6mgaI1vRn3fpgBdydSREQvYiT6hzPraQq6G8wRv3Q
m3ICIprO8jdMAJSCazhDutuxqmh1A7U0VtsgR468x7npb6WAC41KaxSH6WG/SOvl
RwSTGAEZsmkXbKZMhZ0TV6g7OgHJy78qz7QffI9knjpBHj7bURr7+bLlxKDCf2Er
XItH2cBsErHTyRwGOZUGXXwHQ4hTJ4OcBLw0ipibRReRPiEQ8VOsLvDvMWqe188o
VYDUc/8Hdedu+2kw1tscfTTBkpTco6sY3ZuEoblF7qa2CC1Qo9aOu8j4s6dw0any
MIpyHibYuiyLoFPEyeGnyjd9Hs1YBR9dksYsfEoKO13gy37b3jicwFMH8Tr6WvrB
2vaHTWyujptoEUQ6jkrX87Fn/DFKTh+V7x4T8dy9SJP5K+NMTbbpp+lJg5za4548
WTTYYsV+rWEJPHfIjMdaaGc0JB0lFfzWMO65xPRBAYZRKk3FQJSqTYpBU0IsEBJX
BbXaF4m9+EcIyXlS7xougyrGz65WkIkpoYSB2nh7LsEDoHBa/2f8L+7bfSUue+5M
Qlx7ly+H4CZRzGSpHTzfR5IXWpaqDcZ4VD63yR0dyb39fnz8j4s4gVr1otVdvhKL
TgCXWUXDYL1+ZGpyexLEO2/TOTk7H/eXMaidW1hzxJw+umZ7yqt5m8p/j3YOS0Ma
6BKtcmZ2HOQnPaZAerxtSGErmr0IT63DoKTXnq+a9E4g1Dvs8eMYPkWv0lKbiQmE
7xqPVSnrF0vwxGqVCGKC/NhAMzQj9IFFe+ThiFl+VR3AQKrcSNhD0/c27FcpXjXa
yTqY1LqGoFQrKf7Jya+wVPY5QlMdvP3QSDjFJtZ4I+yyOszkdCd0A9l/Vih7lxwz
UKmMjkRuk6XCbf15HxPIpUSMhWmcRJn+3I04Bqw4dtBM/x8BkzCprEc5sNuCQBtQ
fdxyFFRKJ5yuigb9snns+sDPOOd/EsMcOUJi+aPlFwR7Br3Bp3cCyLUA98ijWZeo
WtpHJ8xXQkesY+qfkq0l3nIABpmjDb9NuhMBbLmtGPV1VEGjJ3z83T8fOzfV3Coy
RDCvHvKgHs0lBYnVcy3Ru/L/0FGYqR0nfq1WCKbHIOVjfqj8AC/CiVl7OSos6jBw
bkQVEFxhcgycDBTmrb/Pm5BEMpxVMYbPa+mqyYL3/3MxXEzp+D5TgwKaQfMc72eY
rB6wFk/eLRa3JKntU9tIpF3a2IbvkSKWaHbEIa11Iy8xjYHsxFo+7xzfU4JV6EAy
EYWljhYODlpplX9oDzlqeWyT0T502AUYPx10fWNChOu578/Ks3y6JOJ2Bz0ib8JI
mEBtUIF+uv6ZLUSA87pLMIbw9KujjmaAPQtZMfwOLSueyz0pz3sutuFmSeeHbZQz
Dh31K0LgnHFx+zpXcRUWSjJ8lcANVGrZlq/qs+dYqOGr3c2BZqhhW5Gj6C2N6cIL
x6CsnTcf7bUUDrs+dP6pTa6f/SET9u1llkojuzL13wpwuhsCHkMvzLqAu3X94tm7
M/TJ0q1XhCCJO5HY6Xy2PtPENq5XgCJTOHkBqYagFpp1x30zkxVoFc37BwMRGniR
0LbNDpcEyjbecRmlWDnM9gg4NoPyopnFUkZpePyl/NLc/QL1XfQ0tVq8og1XjQ2/
zxvMNgCOIHNQqXJqHtkXq917F6mWQdqDdQPPozyguecVJ0xfpbI2acBlShIJaa8L
zLKqVTSQX9XC5cmbLXP6v0gtSzYWhGKlFoN+ZgCoEqt8E3ldzacj/itVQzMnFvIj
br3aqkZyzsN1d4TqEENAxP91Kr/zjlEKl6RtWcwFMByozjauH4VfcF88gT1KG89M
dIyrZivyZrvIOAQtIfissFoifjST39WP1m6DFSlNpSb1Ww+LJGpcHo6rTtLk8h+H
yUFo3fo4lIKJuFY0jK4iMXzHrEu/7jGJDIzxqQZYqXnaarEvcnWxXERIK8eTbujo
iPWKTjiLS2TT4O11kUoePc69vF17HjNsfbYkzlDenhwtWlPgLyqZVO3bvCBGxH4b
ROGa9TpdxuVJHLvlH2g7WHqZxmj954lojKFzlk58njyzOYb7BEvJxv0qE1fCIaIM
w5XvAu6BpLsUsGBsz1/LrexHqGbtGJ8PcJa0+qRSKA6Da+8M1gvVyaxMZQy8lNof
Zcodf6XwnyZ5IpsM6wTclZViUehcmPyzGJjVHMA26H4tvH2A8MFZvRlIhLEvS+ij
w7DHw/f1uIrLX1gp2gvNMZpt2GN52kF7zw9Fq4MHw1RO17gmsTWBK8w9I5elThnh
Ss0vUmzsXqk/qFC3BrteOMZofPjbbhiKi76kA6kqIVk1CLH0tFEphygSM/jCfRf7
WoptNoTBfP5ccL6s/v2pYTlaxgOW3pCXhwwOaNwTHhz8OxXIdqSjPjwwxn+mvtPn
hPoIvCh/aKJ4AUqZpumeNOcfHzzS9w38ekciAOHQHMSBc06e3j+S2jQIo4SsG8SD
GFgQkv/kCNDpUq2SMg1j8lhFB05wWzP3oOhGFnUwjBFjg7N17pVInCdSTququ8t1
YL6s4fd/s+sVZM19pjdE4EFcexni4swF6FNfZowiRmeu8MW10coGHrfICZJUo6Pz
DQ1SunqwdL6EtKRQvv52bqQHH4LQVctN0UuwaNTObw3wK4YWI13dFE5LTkW95yyo
6ySFNcmH8XVpB/v+4KCmPRgb+McqcsY/M3ZpY4P6fy41AibQUDqgCzpBVkJL/lH5
BAgQ48YUGGNbfZt5mo5Bep+qHgBYxpxF42oF8wFhDMUMsTcKHIz6JO4EexsUVNwl
7F6DD/qS4cJ6x4K1ued4bqkNhaUdDz8kuF2njACVfu9ytnu4QzTt8BVA7DKwfgKd
5fsjVmsJdehx9UYHkQYp75b7X4LfhCQJFagylufkIL9kR9etLntu39YCI42juknv
b6NEfRwcYirMUPnPxy0dUaSje5sQLt9kMs396dDpZRxx0QaBlwGllJZ8a1HMavfI
oeoh3OOQcoe05oNeEK6XK2N3UBEdZdnuzGQ0wyGw79MFcpG69bNAiXZXXQSLPDfA
MhN6KsLyVgeHmEWGQw3w+0r3uzMwrnhyBfF5/1qlrHS8JV7Ph0KXgN9YEH+L/Jem
AeI/crQY+jnK7wUCz+BiZ2X7ZSBGkKBOEkW3IpOGodGF+/z8Qj9q36Sr6NFZrGcy
kpt5nPdBCDfU/OvQQESR8yI5ca9ws0OsfMKKEF7sjr5nEk+wzej3P2UzQKiZBAui
iZEWumHNrr8dpXBXAV02HruJ35t0ps85dOYz1MRTquVPZFrrtu44OH1Dn4NY839a
RFvELnS4s/X3I2qrifv3gjQgA7H2FTgxvneRoRzpyhcjJxIirARH/00R/3idr4aP
j+A1qulBxHSkLNZ8KH+vFKaCbMUEX4wZoX+b8n4N1LZ58ytgZAxrSpplAi5esudi
RCiH5bxJmWF/ool5fakds8WicGNaHDF08sjtA0wE6LIAoTWoUT0rwMjNpeG6SqCf
sCkFQtrzgMN5LPLheMrI84rMLeh4s6sKyaMsirfO/1bv1sr4F55ezgy6aSP7QT9C
UcY1rZWV3pYIdlYYSjSqieonJOv891cMN0uNG/+IKGnhkEdY3LZ1TxcpfYrwVP+4
bvMsTIdaZKQJ8jNqo73swGlgpgQBhEfWSPeY8KkjSqP2W6QEj0NrgmafN2v9eyBQ
reC7cAB4gWsxF11TIxvrSObigw5UFUf9LrNhW6r7rtNE3ayXlxj1bMREk5MQ0Io2
5IF69Uh+1HwfPQ6HIJeh0+kAOFKhAw0thaaPVocn6Cw8xU4Z0i79rLccmGh3lBqN
nCeMU/9Iq3Y5PpMtSWOWMdEIKoXiOZrLo1PdiKcoQ+KKr1xg5gQ8Jrt3Vc85f0Ns
A+L9qAeZySp1ZSranj27aVdbj+QzoFKQj2hQfCNIMKnUUp+QvxnQnnX4ky62EFAc
LNnJHRcXPCqUcNG3lt2tFYquqKWTHPKA17Hga0Y0ft7cT64sMWoeDhGeyIYJatQA
uUiXcQJzVdXPGVRkmMRHIXlItSg4Kdfuq5HXtLgGdyPqC6rFFR/8u9okgodvHHz0
jL5thJIAsSugQREYgypOi0O5saHJq5zE3Q5dkd+q0lwvffr9BXy1xwmIVlQflT+u
SYrH6Mj0fbi9oAjC7BDcg7yd00eqm54ReweoN1T0urOqpEVv2hqc7K9MK69yXYE4
XlE1z2cTnej7Jva4dhY00Ag/a4+KHTfG7atmhT/Lmdk79+/oVBUmMBuLeojqsz9b
nfiwdDgBoFHhriWptW0Xs+pwUWC4BtwAojBY0eMqym0Rc3Q/EZAAilqTuDww/ppJ
f5nOaoVAQfe/qqEKBrVFRuyCSbIugqraC6Odr3U7Y9WqrCMyqbX/TfeBJ33pDEYH
QaAZID9y74ebiWEjZl6zVbjUAx3nyaHfMIJ/pbgdiSp7gdvqI1CcXUKqTBFMv2DG
raOlBlfW/JuKCT2BXTJs8znEMxtA2NaoI5nelAvA1p3YrFtv/kZeX//OEFtLdRyg
6dtz6DtOgmqlR3dloNf0BlghpbB0F5YFnEzL6Js2BXN4LF6fDdsF3+0TleHnG1yt
yOIw+yYSGvHNbnLbTUV64NjGDA5AudgHWgBvUivoDUDsp8BG7bXiNgGGzNQYCAJ1
Ja71FswYzv9u1Wbk6OtT4AFIhYSiqiRZqFrtld9skNdxlE7XHWUXvYAIZ1xM/4vB
eJSqMkqbEQzJMnn1VKM9Rmzt6NpoI/RpAcp5RIAcAwkTT6PNPHKiU9IjuRHACknN
e1mJFeP07sIOvc2KNO5VxmdpadTI4cOkxxM/55UGlH6XBfXA0Kbf1GC+J48F7Rbk
sGt42UMWS45ZgFGPJ9KWwvNOtEIIVaBJd+drCGSpDfs2JMEJ0P87NpNzUN+Dhqd9
+ApBUuMRk4tNQy5YA6VYxxUGSn7Sh63T9M0xN6SExPxq3UtOTPoRs3ffZNDwAIXH
ACYT6uCYG92aVdvbSGw4DVVdv15HNbDICLNo3AQOlG56kMl297ijXQC+TAl2ZHIh
mAAh8mLq16GLkcZh241wFYIeB4jRwAavcFVN8CoCaDWo+a5PXvgh9JftAzRHL/MB
YMCEAugMOwPOYTv8o9R9onWnt3+YHRjoXFmYLGiTMkUkKhz42ADwSjlCq4KOzgbl
7CCtK+CWW1BZr5Ik4lF72zRat/kFy3naVYpbxcrNI5Me2u47XW8FyxKHRIr2qhd4
zkV1vA6mWqbrhbgH0+HcH5UGDn31jgG0DuIiWs7qFQ2tvcb5M6IaQKF5EKjxxKDz
cBPi0BxjOvgvDkeIMLUugZbxvWqs/slWfbkH5e68Ys86C/AJNLFVKMWhfRRmphpx
VF3C9HaPp3s0I9mZbSs8fqTmkvmdAQBKP3uKPYrRduHvUOjCSIFpRmZi2A6jvH4G
TK07lPf8OLWQVDlVowGMaIW7Ud7xxYABeRqHvTf9VrmzOdoMwg0Z9AM+ZMisPSZI
RZmcQaJukAvi2nUpguFwVjGvg3d/ZUCnULWye4jRcVLdYPPTPrNYYERLNtwa3CpO
cz3l66zeZ3R6jVvdlIbasajhLcVUMjH7VR6QVAnMsG78lXaoyUKxNHsI+4rDyfkd
MUYIBEF73zpH+QsUBAveTjH5t6YyDVQld3iQkS8L31OyImFar20d5bJaIXg4q8lA
z/tddhjd52I6pZ4ZApr+mP6pgSSXFF5TrrdGXTA7VrwuFiY29pRRWN78ggnU9KLZ
XHP8ctCA11MXr73y4IAmVcJpY9kEKqMEZqAXLJ08Ds52HNnQ/s9WTeveY5lC5DLn
lQ2EwYUiaWUStUx5o5ezhtuWCDR0ccD3VvCagE9jo+1D1DOxHgOKEvDwqXkTGJ0M
dxD6xSaFwOSSgaohooRiAwNYqhrtGAQwRNSevvhBHitRd/DoS+rW9khDEGD0SHJ2
s1L/m23Ghtaf9u5UAl+RJo7zxbRHnn0BEQGmpwNUR/AySnKN9QTL3TFzu1eay8Rq
FMYvHxy8v3PatT7bxb7QZkvC1GLyr8VI7J8BaOl32EXhHiX0/saKtLFu+/5NAACy
rsrMZmFuJrY0UJPaZSV5Bt9VzCYw+Fkag1YErscl+6acyE4EmYn5pHQNQ5c1Nmgh
WMQJTD3/wm2WN6wvLY8lj82HKKGaPPo+pTG5nnH3D5ezTF/96/Bq9pLjOeqQiNUG
iuANtegv8p8IuJRfukpgHZnLmUTq9GD9BnOsACnotcVdPTbdR2C5URwJFygzyLTI
EK+X86ssBbbHde1IwFzosA29aEeQyD5zo8rWxkdApB+bfuDuZ/uqh644MqZRsUHz
eANm0gUbR80r9k/gni5rQhxu9rNw9e08hMR5EgjwOTEbPNIFXV5y9pVvZDVI4f37
iBSaM9PsqFHaE9fUS9ncHYixDeGpSJATG6xIondrCn7dNyA0C0FxXyUwCum+QhKy
iFpd0R/MNXbDkU1mFomYgKsvPGB71GnMrqn6JG+xYhUgrMYB0UvfoN4IX78Yso9A
RMUvxAGCKbCi20oVK2uvAMES7imPn29dFossTFkM5C+NXON5wFSiKrsJEp2xQgn+
Q1ZIENDldb15+ZXRpqOQ+N/xI7O0DBlhQKIKiWS2/5Wzh3Vr3PdVt/k2eFQxtOt1
ikKfaiBpxh6t6QpLHjTWJxsTAX/fafvwwjeMd2CekWd9yVCwLE/GUm4gTLqTS3to
A8qA8mp41p2blq3s63pXJcY7SzOviNawGt5SOTOgV7P7nn0leJXB/C5pvI+Op9i4
/XSIkr9lToM2LZUZivtPmUtWwX1XJhCMSDJFLebqQb0n1rMblRlpJ/eds2AfMIJi
Wn6chIGjT7iID/895msHADVVYymaRN/fVuIiU9Wa6zSqH0Ywk0cpHhgUfPjL+i5p
BraccnaUKEixt1bRUyKSc3T1VNi+aZpJ61J6XHCcLsHGnUYJdjQX2WvaR7wZNVz7
j+fbFd6ERszQ5oR/23VNGn27SJHS6ZBcS7mEXUyj80mrNb6DYgN7Lzx///9NOHOB
bJroEJJfPUGx611RoAZ3rWXqVHM0+/PyrOW0Ka4qYfhU0xwJnwHx8vOxqkMN5lOd
fPOPImiSr9h8MZ067c1XyymCp7iEFexnJqYLknAt++pDq2xQqyDqHMFUi1ZFPXu+
r6PwgiiO7fSChS3uTg1PmcI4Tcq4wnc8+j1WqTW/dFgrMIfeA5ih/OdFi5KFSRSx
TN7IFMcYgDPdpC69Nf9fQr5UUlsyr/+SxpZxjKwNwbkLaEQRvByxkF5OtVGoAGAR
vhj776QPF8C1tuRn+cmERldILA4fr+5eE5pQn9FKsMGgKy7zwGilkjLme/MSTdov
8oPkwP1V2TZrB4Idte8Fh3qnHPM662eYNYSXi8fDOoo7OmUnq21Sch7H8jeHaSKm
nPr/UyGg3RPiZjO5sYdTU1donhymAqfXnoaZ1fskdq2hm1WP+DAnT1IFc0VPR3gT
aUb1mCmJ+UDKyRorSwBdbXNwzbqR2drA/+/qLMUzeOtCelbRc5hj7NE8F1m7JMw2
opFNDCHkqcxn+gk+32kTHUTxXJRsU9AJtH/NZXWVvSL07ZlJMxQo/N60OeE3z8hB
bfz5wIDmTYdxFeEF/Ue4v/ySowEIDOM7ClH5y0C73Dw22//2YPhS/jlTY/THSrDS
if6WLRfsLeq882ufQFk2EuCS0aAeT8MkIV/ZsOMBtMleVvvElKYXUx1kdOaCgi6d
DsFN7w1fcTLCT+F4SOpF5f8WRNJaAheUcA+vHB/M1d1aNq3De0TSM6194poVZeW1
bj6dk9BaSGxtt9XDS5XbZufqWUvVCzVwf/K8c0w/5dcmp1FhLxC1xoWhKIxtwCWb
rNq6vZCuEOJIevE7YPOXY+mHaHUhSuLq0W9CTLlRtf0dkGETqRwHCJRgdYm8UJYb
foPOOxx3KOMDPu99AUui+OZOp5ZLaW6fMBaJpQ6lT0F8d604uz3l5zRToLEq7Dlr
ap1MbnZlZk5ZfTxcPupbPehg18K99BP0GuRzxmQ54tSZVBBK2bRGUdDbupWjouf5
USdPP8FuLnKCFc94AZ5j+ivHyr5/eBlbS+InCzooDWN4M22WYfVv1jkZcERiRgsV
9ThMF/sa5Iwy4SVFKj+j0zVsDu7j5f2tCkuvC6psyhZw9a/QrB6J1bMSdWsPZC4j
WjwLbhf5KmHNS6LFyQo4huJPwOoU9HBFTlGB3mc2fi5Su2GEx+D+EcX/6c5x8jtK
y+XoNq40eMX4AoUcq2+wMucaM19esRAAI8S08IGNZsm1e7LMoyoA3YnT5NPFbbsw
fcquSkN/tZyfiHYsgI1j/BE+y/QiHnXQNZrMXW5nIomF955nvRxgH6gDtV7I8ukc
ZmfgiMMkgF9BNM09UcZv1B37EXvB8KZ+FZmkDjmu3SX57tvzfn9/0PayLgXuE1sL
ipSigxvic7/aPZf4uo/TtyOHr5E56FZc0OYyLKVDOag9I/8X59H8sHQqw4wek4qc
l3N2xhrRioCUqJgFnO54cwxHUFtwXz+rX6HaWZA5r3Nx2uRkLqQdu8vdO02q3bTQ
E+8bAVPzZ7tVNsLhjLxsfnHGPa3INleqNUC0zDAxxhJzyRa6S5ih9ajpRZMgW91y
d3002OitOB+lJRqJY3z+i6UBcIE8VcZS9Vk9ipmwyFREaGdrY3cMUyStV/iGwy6+
9Kz+FlFA/E6UcKT/pYLqorbgk30LUmUcbkwk2bmnMhGZSTNGpz7IggrjQeumOT8N
9aW90sLtIJEQPif6ajPXpht7pmrSEsSpA0In5+MCfa+SQn+1SXmAvWae4qfmx/KA
qaKj2vQIJXMJrCk9knJxx3ubHaOh9PCrgjgm+3ydCqP86paX7ST0uomnPvTDbfCv
N7reiaMNCkGYU8jR2OeUU9UADWAQRhJc8Om/hnI0RUkQGO2FcCYosvg1Z/g0NvAR
Sd9cO1MY2SYKVOW00ICtn75wITxb6JeFyPzt43NXBAQ7NB0RnN9axkIUHEwUb6Iz
MQrgRfjQu+uLSpS2silxU71UoVes4RQ6e/9/y54CSF1nC9y3sUdAKh1XTV5cq+bP
TiqOG5Jn3nAXZ65RLJRr9j+HzTQoShGnTFRDRv9xHKKwRtIXMVKdLOl+uGclmQZG
ESVkcLuO+E95bOgOZa3kiulgwqjGJtFDsyBrMKwH3+cDmjMNr8tarldezmyPbh8X
jdJtvauC/i3Waz4B9eA/N4gY0omsIGcQdI9RCN4V4H9/yL7AtmjS0PSc1wHEMLK4
oWnGtFFNc1Sva/ye1Uxlz9QSzIhC0wCzyOAgkW69q6iQxuMzeBPo5nZTHnNIcF+e
UG7Rch+hugHPX7CF8n+rt7/SYy7UmXJdY7WEycXFaHBWhhCqv9wsecPb+MMnolq5
tUalecnWvCLv4J+U1Ga85nP5MiawIIyzyJFwoCVuNAaq51ZDIoG75m6UWTlWSLLC
cJQDjJNdw6T+URH3FRMGHuAMvdKqehJyldDTqoQhta6pRgEXqHnwIQpwKCGdTRDC
kTl8Vzj4o+Magvmco7eUfZp2lDA6lSqBLS8UjaM6FhO+++dmOQtSOqQyrh0xGaB6
Ta9dtvPVqVXSobA26x+Apr5gdvCNnwhxyO8MScsKw5u1T11KeSVToKJ53olTy6LF
I0wkAyInf5DEOVVgH04v/E4kprOXML3RleVk1oYJIpr00AFCAO2tkCbsjPmOB6Mc
OCZxQDnxpInp0QQ1F9OEshFV3UcrBFvBkLrBD86jE4I+O5RWdBCzWMp3WZr37tRJ
dTdMm8rqb46M+lbl9Zoe8hMUkW1zQB5Lssn4dui8BzXw83g7spIIQFtSRY7bE7Je
TLcvJIvQmFmxLIPzgLdkoA9uExqhUgKbhhZxb+3s546+xETZYAFcsHJsDdrpONGl
fslPvhErovfXJLgiHhqdQGZ1Zbs5YSYKr5q6/SfukGXx1wU/GdA1kN2INqmYi1YU
FuMXwU2CycfYi6DyZa/LGKEBvwjuXDT7JJ+8/VR/bAOMYAKXL+bb2f/90W3CQLW7
/Tpq7UORPgT9fl3CX0GySZc8ZHp/N4csedscI+DjsauSiS4tp8h4PF2DMnCNNnY/
b4oxIU87FRcglWpG3xWydMKodktoWT5+RA7N7xvkY8USyFF15zTdm5Tf6B1l7INB
cIgawYM5aYzR4NFi+2NzQvG8e7X1zBwXRRP8MC5Wt81cIbH5BjnH9P8hCj8RdAfn
qlDMeHOn6KO5WSvcVchpO7FE3gFcE9goCpmCe/LBjxeOOiyEOCYR9wv8OvtMX1u0
vMcO04z+9BOt3hNiAfF2T+FqActw8xk7GBL0C6EoQkYopz7w+5x9i+Ifw/FGFIHf
BblbieA5qaJ0hMJjPoTPTZGDOVW2CJ6VX3URvDrtLqzMBUdjxWlc7Wa4Ug77Fmlq
g2xRU8xg1CXqLzEwCmIjlmmYeZykqGMmFi6UAYi+rzl+aeZe0xICfmir37G9v9is
RRY4n9EhmiQENmmSz918BgQaHeTmqtsxNYkhpyn74fCkbAQZjLO5wE09DfTbs8Y9
AkzfauiFlqhbqbPrd8t5u5SzXnvictH5P+vAokU1oz5fQ7Lgt5yGOaQdPAjg7bLA
cWBgUUNJhx26WhtOc0NwqrXEcUiRJji3HgDWdHU72wcXAJmmVfdn5lu27dk28yE8
TTyLeTYAtvi183PCSXJtt1poXSu5jhYyGH/TDV+IFResVp0UXeJZCyNL57jYLYOU
bhANqZRAUlx3A1g1VUB8lfRpBPbjz9RruYdvCfukpgTdtFx6NoIwFj6JbMprAGWd
ljUJtYmn4c+Sw+aC4w24SWzkTFhrF9nz5JqgVeCykUds383IzbXdW5jmUY4EWZF3
QJrbrtr8aVMLXuN1/LPd1CadZE60WEYZCJsaXUI8swabh+sJfo6Hd6VtX2gDT4Ts
kFrY73ZOvo1jsjKBaN0ZP+W+BD+0pPP21l/EJRYXgpFnWDOhjoD7PNxfSjYZVWqT
hxzuXOpiO3F7gZ67OApyImuIt/eIz6cjclGMAfsfZ/QGZkKfao9Kd5N5kgQN4QXz
6AH14hcvu4SbyokpWs4sgxveb7cnCjfY9njlv/Dis2rzMhoYCIxC77ctpFC6XZhF
flZ28jHyEoRKhSvNgsAqP0qe95MlhkrdlCqarAZ8QTPtGXX1MKKq6lnvbdQufJM+
kIqRfi7TyawF8JXrFQoBelAEYHJN4zXrH4ZlA1xT3KF13olJGIsuiB7w1M0WhvnZ
iKMdNRFIQYUHHSLpteOYWC7WYiO2cDBKU34W3vnxVc11u+VEJr3nbYGaVD1ROLjt
ggIJCLuLqwjiZVNbZG47btzmyErr1J7GBwnQVJuJFZuPVB72ftzhIbe4ltTSnJSZ
ZfBlGG9MNriuSM0S6Q90+lDHOMQL/ZpJYeIrIASdFoBnPx9hwhcQ0rASzS/2Cb7s
QizvWdL2WZtrusAXv8qsmFrRBuCON9wNP4QIbuX98ZQQO6Q9t2TVqG6p195geCrv
ad7g+8XhxdGfx+m2pVQgmD2oQd8BsT+LE3Sef0tnMyDgHJg7L2rw4kXYpwYbUHg/
Omd9kmytf9BO25rFsgk/T6itqjxphZr5EHyzH/fF1nW7B9s+XYXIL+zI0aAktIcX
IGLl5/6qhihB+yqg/smmMaDjG77RHFiQPU2rU/Q3Y2lKya/oD1AIFHvcTQyyEb3C
SqLILtpJQlvhZBhHmKZfBtfkd4lkShK6BiGBqurUCtWxvWAPSWKvdPVAMU1yhxlF
xWgUDNd2CjhHgdKz3WB9MRskNq0sIqYnxwGnfShhKv2krVTn9bpk6lzzuDaOeEnA
HNtFY9Y3ppFwxERFEV/fbKP3E4Q71/8Vc0MtgdKHsVUokOuEV4DFVeDfPazuYG+M
MiuZTRUouQUc4gkuZgex/SXWdImooUb/ltl+Bm+IjE/p/gah6BMwP75kSKYRc1ba
LQuKuArMyBeaJjNzRSIMKf0ZGbqnDKw5f04hyJh+boak49tFCao2LP40T061t8MU
vWetRGQ9lR8O+6gH6oXor3BauGFAoEfDw/oEkGFqUJINdKvqFfQRZ28wWFCHkU8g
7KDKbnLMDee1zmHNPtx0YV/VRy2NT81oo8kmwYEiTbSuMFStKvSmSFcVUD5DLk/Q
S29df/IwNfiDJCaNE+GQakG5O5zsnWe3RlWrRCZs2WJMVk9ygHUikUFJPeF767va
qU115hcMk4sJrIle+AX+DgX9dEjQMo/6DAVPHPAQHMpNViokh8eT30rUouKK+CdS
C8SbwbFMTxvfD/dTNqhmij4ImVSYMwUUnm0R3ktOSbBUVQww/3g/CRScXYSGaRP5
ACzB02lcQf3A9RPBicMmKq6GMYMFsecdtIlTdbtt55hDeBNOarbQBlt1sVkfD46m
65NnzxjV2y71aT0B2WgRzHAIN1RPn+hYB1rpdhY3rmwV3n9ndLYNm5T6ltiYjMzd
etDTz+fFpS0EAugGuMA2GFtjTnZdwByrDUoC5IO+CdaEwI0zkG6nD9SSVEmJOkpv
DAs2jgC35rMf9uqACI73WFbzgUDwx6mRsODFzwlC+6x5/WLhByG1OpO+WJeE0g3m
Rpc1J1zjg4AHPEAOvZGmmbdTbv1whGVLaFDYYnpOriwYALzgQNGgSnDa7dS3a8i5
KUPLzIKaSxR2VJlmnbhynPjhhGNAIKN3PrH8g+vecogbNQwS/3B40AUilvmHfM7j
xMQ8OxFLyCkW0fjMYD/Xyv5kvzX8eihd8RVkjyr6Z1U1qWCZ+f7TG4DpPPY/V4ZT
oMsxbcDAUxLVxPNDVLCNguRJD04SOPgaZIzpZxpZ2wasFG96JhjFqlonBuCIail6
QIUI2JP9L2cEe6D5sVMtXXcIaagQd4n5si5yVLW9uEw6Zjerqqx85W0yBtSKswMP
UhJLMZXUM/Tf3f0c8Bv7HAJzdYzjsRk876w8Mt0lYu82NDhuEBizD2HfHhv9rtFT
o3Y73e/LLY1c/uX8SMIjxhsUG4vSlurlDSwHyBg/kYEvF5i0xvaKAOzf2H7fOQyM
Gh+7k0O74xVF69jL+KI6hsgnfGxwSHI+JNAgCboanWgufsW3dIaLOonQx/JoXjLl
FrjYjmIPT46IpOWx9zqoO18omtBUxoRfyVZTxSPYgzFmuKlrp807681t6x+HG88/
grMiH603woLOMqIggVF7Tp6/RpYMfdAI08voiWKGQMYAwk0efnvYpB31zi9zV44L
sqk4CxCdHkKxzJQlKvJFUPhzL4+VsKDNmy6Rsm2quSm7buDvBSecrsO8jrgH2inw
MulCsVDkuSZEKhqjNV49b1COgk7N5KsoD+H7A6/RRQQOfVqCuQ6pAX6aMZkZXkPt
zdCBL8IvVz+ft+rHB9PKrX7kfdTRnl2W9vQ8NUo3gkvTM42BCGOf9JVUjUFr3U97
1g9Q01w8axZBTUe/XC+dk17DHqN6b2h3yIOfA48Do2Mw/sXlxC46PawpuTRII3OC
qfDBHZ7wiFlrtP0axsNhJH9TU8VjP68OJGp9/Up43M6zCKUIeVrMikv7MPvciY+t
vdQnQjyicoMzzxdo4W0fMw/gp+1ljxYNZ1r/6iOzSzvlklqYEaBn0qA9xtAEZaFf
2va9R0EtJ3ryBcivZAnzH8IMMj7F11Qvns3vNOUGoqtDZRa2K+deMkFXeO6AgECt
DeAjsXKTnm/CuDKukyR81wQqC1uuZWLnxj2t+63j9of9LVNUF3Gtf+src5dtakGT
srT+s7u+HKQ/yHD0LDmKg0XDoXDIPrOK2tI+AQY/ywH/huhXIR1f9zhFcFG7pVZw
okKkiVXr3pWEMtTi1Ew/R6kLuxfkKR+CFVmq5YSl8arJnnz88B78GHk9SXr1rsVA
5waSDzTa47SPjM7tinQPFM8mSoaBIv+cgHAcSA90q3yAcZCbvrtSktWbIyWOSevf
DTosVgM3DzomC8PH5yV+ecj1Y9+BHZMWm9lDygZlfDQS7ALOnYvQdnf60Nwpzgp+
UknBGISQtVtKgrqc5kp6zTKfdcngFEyILQcoLsmISJzdoj6SLNzgS2mTrQl010a3
EOYcHhKzQqXSdzjBZhJasrtFMzLnKJHPJJCuPOQzwj8/OLHGlUgK9yYHPZHHKENf
E98A8GJvVpgxpt00TIERspLwVdi+aB66QSGZpaDbHOCIbLLHbH+fKFSxk+B3D5jj
LVNTdmEmHYPoO6nL/RZFOK/8rvul7L5QzUvN5pJHr0vvjuQB+rkrznXhxdu2ZvKI
f2YTDE0rgX/VzhZ1g/VTF9v6tbsGKCzNNawlNUuYYzcy6R9FqwkihE1ZED5w9KZv
n34RicCnsHO3Fkx3zStDB3jc6+sWjzaLDRd2+7f2yPySimWTCjDHPoI19P3Su1/9
+4u8nWCOoYs2Gh0Ye6nAOVzofWR639MDZaerzOWchYALIOiaksmn87EhSLp9oMbg
tFIOyxR+v1BExEFXZXsxD1+OiAd174rjgQtKhTwTvALdRSi7vgSmKA8s00dXqosG
E35pwKSMRmfbQdo7MW3kN4RSboMelXfNp+36qO9Zgjk3oXytWbrehKJFvPT1Ev1H
mvXjZstTYGQQfswS5cJwPywVHXb8bLCfl5u7r0mdBOexyhDuWwq+XpZ9ZPuCeAWF
1CwCpK+BEBHRJZvuBj0LhqQZ8nDonU85f8cY76xRQjMtiYAY+aIfDE/80WucorIi
7xhUJUpZEq96MImCX5hCrtykJ0+RxUjYdH+XTe5ueRl67e8wBczZ+3vByUgPLDsV
TJciZnsXm6kINKyF3rNcHoGu/eu1YiXAlPJlGAgADDwXZ7ZHh9CaUbrh2QvjSt5R
TqYj4D6MNrM6V/Bf6MOlRD4i5EpMFHoKcOKPRUeXS74GdrgCQIJdk0/Mpysy9Coo
9+8A9iv7rjQZQ5RevGzgAaNTQZD0+5SQRHheg2EbsWBWM8o6C7CqmQWoIqm5LILq
f96RMkThrepAScI/iTu6KFrTsDQfLmbZRnzcGeg+6Qkajqk7WznfDU1uHDZwHXkA
g1oP6XAMGSvhhi/NSekFj1bWbPhiJnRcXnQX2pa8kI+R5MVlsniyqdkHk3565FIF
BL7fglpGG0gYLN3NYAKWF+Ysk5aOPQd15kes/sWKXbpXDZL0BUb0kIbUOV1CNKns
hPV/uNMJLQJLB/AVSCrt6pnIs/ZfBHep5+aPNqgEQgDBTUF1BK/MuFa2wOVVRg0D
lbNN97ayFaXR21KKiwKy9tCdrPvI0QRBEydr712q3OxGOUjJOZ9DIaOx6dM8ksHD
HvP7PktHAF7+5sddFgQKdIdsxrB55nRbIZG9WhC5ZzEHzgguU3vMzxkm3uCp7eMZ
Yuf4D0hjhoQoO/uu20jYloOTanukZoRxJ8LGSif4hmW9Hg2WDr1TOrA659BRD6IR
SVzoiGzRBvwCq4c6xzZxD3ZG5RNJb69NMmV27Fea0Z6GjYSLe6ikPJYNu1LMd5BI
qOQQQRaYZnhs1xubTrR6S5xVvPcJ94Wv++hW2lt5xeJjscH1VjIiurR8g6kggyly
CUSXyI2Wl60yXI/iIX+P1tvWq1myo7VpLgiDj2YQlGAb5+/CfrZiZVrxpOgQAdPG
GX8G29oBCoOKiIPRfjLNXvWaTJdU7FTctGFWw9j8i31APuCogjmn9BYGpztB0X2W
KcUpwBGtlebQbg+4xOpi57LAPY2Doicrpr/QNia7slHB1GCvSZG8VZxsI0BhaDrc
qJ2rUNm3Q0w3n+IkBJ+lMCJALQBmmZ0pisz/Cm61cxxqECQ/N3APzz7qvcBRKdLs
dqwwwsoaCpGkzPpUIuuoRerboC1cCYUXeIiLcSb5bdZPM9h1N13yJQxejGlzwj/W
gNU5DStzr5SImtfTkYhnTSQNsDkpNeWwDEdURlEgQJpxK6CKgXC1Y+hP4JlORB17
iiOJA4FmeCEWn1hWeXMHdH06QRrK6AHQ1wfBVa3g3oBMRlMFqMgl/4PUqeeAERs8
ZRd9l7scKhxRoenDMHb2oGK37S5g7FfJfxjDqxkT/tlGLVArZMnnwbx1n2rNGwku
YGixSSvl0CKQW868ROlRqPFWv48wQ3WEQejomaosQBu3G4EnWdqK/p+4UrFPaG2y
nUxUYu5pv1TSQB2gfruDrIzFNOMbyHksW/4mK+DFO8t2srhO1I7F3+9PkAzXdP2M
WK0AHnQas3rQH85+HZntaiYMjjulHI5dIy4RMCHmRWmzGVqBRc6cDnDMCkZrNcJL
u2Ws8wv18mkBctnvPRwzXXj6NEtZcjXVxHThK+Ws2Z33DPAxIV3CMpmD5WOQ8seb
/CwA8p4UltWdHPxq2zb7Tslfa9/oUe+FRBtWJ+ms65KKO6mY68UTDKLfBNWPJMRI
l6Z+lyUC3lxI+STdyoPV6csn26rrCbT5VVI0JeLgHHBVIScM8Fy2q5pvQ4/91go6
o3XcrIYfjdfRXKpuXZdaGtq7GMDvUcHhED3qPDkfrNOQlVwXiLvfOFgHdPC+f3Hl
goSaZpkBP9UHDVL/4Us4l8+KMBR7GI0MVJgYTGjNS9NpgqFHNG7Yhbn94FDgtVLo
MsAmKM/v8ynwOcR5PJH8qUt8PXqzWS7F/a3y2RRwttW4aHMxL4NbjbQfMTBBKrey
5zwmPPbaC13mE4GcgSHaf75jTtNTR2EPV6gbSkZlse8w58H2iIjfmwq5hwEnZXW2
l1PHmxgmT93pdgxP+9NalKBR92bi5ijJgv2Dksp2mjavQHd53+y4hEyVflXQxMYh
HC3Ij6NPIXY6a+FvzwstijONzUTHe7A4/Y1aJn7cHwomAhfGqd9h7WBqxNJFDLu0
StDQ6qyqiT42C6J29x5BE6+aonhCgcmM3TxY5YLQHp1o2hAvkQRXYjfeRyqBzdsy
oofnpnof18dp2Ik3S0TazOmthouGF/uvUtdzMGvm012a2+x5Acd9lLnnc66TdKM6
FykOh8MpATh+bm7TLkbpPFkeU0jyDk6YQQpyzX12VL3WR32CWx5xxadHJJcw9bV3
yTPUi6E+cMH+SOeLUoDlT2tyWA+KT4CaPDWBo6LJnjzrFhZ3XiAribxyVFgxzr/U
ngaj+LG3imm0+NgzgN6Y6O9RuECMBKXpIa3H1lGgw+v9Xphg1XVM/Z/PIBSFxXED
+ORodpqJ9DL247Yx46OayZc4XfJoXZJNXHMI1HhhUnCzYpyBhfNxKu1ehmR69r22
4kvGP3gEtebBrRUaMmL84wblnFmfhkEueqmQ/XCR3Il//vOfQy3QOAo3Sqz6KDc1
bDFlteP6HHVC2LooxzExFlDMtZdlO6hRr8+RiADEFiSzlnJGKR1opZ6/8N1EjvWd
b4xX1TFxFP2JbT/aPSv8M6QkdDKfriKb/XayE0jmMwnLJ9XIiuDImdXD1YMC/Ijv
WpmvgVytlvkdJtX0FM2PXJ0J5LqGNPkT56OQ60zaBLPYHzm5KIbiZ1DyWyDX+/qt
8QVG8HtapalKhqz1W4TpCZbQKs/buzjsh9hzlWI61+Yom2NhCdMbT/+gYR10iDJm
zUT2pqYuH4AFDM3OGHtjFxUj2lkGx7JD5C2sb/eFjDaCmDqh+StNy5bGxPDnmaso
nTgQS1th70sUBZoZ5HhD6uH/QGsGyqwCJTw01TE1wvtCSqVC8QDv8+drdb/7YJ49
uihzgH/FNmhVo/hIia7PV69w59b7toD5ZcuOs+HpDgAEY6TMJXBeGIVfWmGRBlx3
J92xImEhKgqPqeuSPL8c2Q9ifV9IkH3F7gMqG1sv2VK8KmupUsbusgk6KdJN8bWn
JKqT4y+LBklUr2Y4z/OfmCQqTD5u/yTmEqjRDqTutzFM0ED/D6jPuZboV2mXmkpx
4JOeRgu7dwf7GklJsWBlMlTqGSXRK69PW9BvqUWm+5FeKm424zoUdSwTUJG7/KUe
I6h+0dO3c3NhVV1BvyWMPA84YSlz2hlxzfxaIXUc2WI9fsXP9G0qBMeeCZE/NC2V
YBuFvqqywSEi4dbMICTDfdH8urz75eJiaRePWP0k6cFbBWrTClw/ic8os1APM8qj
iwKkMbRnIi/LlVHhH7Y7TLepkuedGM05ic+LcK0GZ8xYhrLV63FBJ8lQNyB5LNgs
2F7XvBabdxyxOE6Avy/zaDg+uUUehItrCP/O3cOLgAnTcCzqbcXzl4/K93L9tW+P
mEAGfqPXusQ2wi0Dgb5imZRNy20Ikei1DMIuR5W7ZQoW6qrf63A6RkMnqdDe4ISK
rbrmOjaUG15mIwBkfzfEP6hsxLr2+7RKfS63FW8Q5LPCoJpjAwWAJ9XnnnzPiJPg
kZc+k9yqJeM13n9sE31tzK5ExAu13DiEPqJJKrOu6jsIF4AZj2VDXJGGBhHh49qk
Hk6DKnMh7yJk0inac9UqWXSuI3boN3E8x5kTBL7FX/z9ssCSPTz/5OHJnZhIGLdZ
7SsmciXBoShFXMk3wNDD3DZOlYbcFNEH3CBt6/kG8Uwb2FbzrNihWtk+YBI9ub+l
iunDnDGP6YWyp2hYt8kr5OdQ0RuBcCgjzaqSxxXA8lgVMF+3w0xpm86Tvi+73fUp
a9d1jq8cOubnmcZMPGQEJnKz3cK5HHO2JdGL/mhPKtjIGJI4EnrN+OBJDxFpupQ7
rR6KWWNXL1ZXBz3h7fiolxTS21CHAra+j3SOymSZteZJQyvtCbtdBTl94gi68kXO
EFVBGg2hXtkkhULqt8b/w20C9CcFs82y4v3PEqE8o89D0nfBRg3PChigL5sVGqXp
OQUFa36P07/2anHrwAWI+jBzJn8JbOfLPEuj0e5Pu4yxhzu7rTZaPX11HyJrguuF
ZfSU7Ry2oDBHmf6QPese4Krx9+NN743Alsj/IAWaE8KbVe8ECt2ZK4nOPccTk88I
ZL14iDiuPPp8bedrOmTxyy2HfvvwBRAPMCpVNvdHVOJwNMS22itaPhXPPOZ55nXv
2lqu4YsKyMFevSL3HM02IY17qRxNmzQTgFCD5pok3gR/sdRgDmYzcxj6wAaDJLXZ
ni8wMaH7DtX2YOFiPBgcZ6roeRHC4sh/950Jx/EIoj0eT4o+lgTuHJ7pwYTDlWZF
M3n06hHBy5DtfSH7nR0Vv9ZxwXnPngJi0M3hdBTrrugOCEq5KMGTugyhoeCmsEjb
S+CJnZyZluoyfTz67rfs3FOHvew14pJryIsVC8En2e4aZADNFK31zDZHev9nuPWD
xFRpyWLNFEo5G0R6okjT9XgPOemyEokT5VW9p4JB+Sn+bXRcgYKrRpBbLjhr61Ff
ffzTEUTQ5Rng9+TzGKStLyMsz18K+92SkXG3SS48XjTx+NL1fxXZuQ/S0BocKfsp
fQv11A5ljzR0D/kCUib5a+LWVTUo58JCXYiJmLYl7Vwpl0LMynN0TWAJ7pXukpIW
AJ97wdPd/ChQ+M00RXFrC8NrN36XI1UIislFxZkfWHayMAMASAuygGIulIuSeNtz
AFQIPtkDgl16EyRrG9NCpg6sTLCoMUJCEzgDCx2H1EfvHQep0BUB/pum8TWw+hAU
yolZpEgNc3P+WH5a5w5Bqmp/e+sEuQZO5yzUelKY9NCc3OX25J3BHvHZfIH3ar2g
bxDNlg+kDsZ+2ZWdbjUNie2+/nDTZhunbR5x9Nr1NxSIw3Sk4059lxutG1+7cux1
73+hRj0DDAC3oeZMGtv0Vh0H1ymBnm536u3dYm6er131II5WvB5xlHdQ+SPZzrwq
aaD7cSQ6NOJsLw/D2+/gId8OcVceDnh8iawQxifSaoEK7vHnI1Fhombr3F8/l8N/
gWt4YK1/TQx1R2zn2m0UTTv9c+9IcueyImOSyJTJBt9StKyZgRRsxjd8TW9x6wDE
EQAfI2m88IHPKxlSE1gQiaTGpoPfTPZMXFAlgxsTivN1q/z893hI01u5ldq0kmIH
5S/8GCoS4bwXdv7lZAIyKue9uePdnlNBTCoQsi8Z8KxHovxHI0Iy98U232lDtE/O
Nutq9CtRxLQOLuil+ns2G0qFqm5v4Q4kPq+9HqgjVrPwHJY0Wem1YYS/BwgbiIHK
FEVLLuciHS6J4/3jrQWRMrVTGMyj0jAaMcmHgQimsATUDDe3S7kHndz/mjBEGG2B
d88QsoEW7+DLswqqBm/nS3xAakf2lRdc28yjJyq2dnelP1MNUuk1u0epemGT4Als
kd81l+Z9nxqfwKDhI2f2s+KGr/oRQigOtzAb42Um2OYrKg29I49rg5ZmE3wmBbmv
N2VtI87u9BlrXs14Z1lna3NqfxdmDOfdaqDZEgOl5uNglD01wTXRbM4nBEzD9P+2
f8SOA3Z02Thso5EICu2W8KaNMO3mS4HWmPuZPiPBzZSvsVA41ZYxo8OktYm3Tety
NSputUjr+YfDXiUPDkS4nbxtGJK7KSMBeirEvzv9d6AKUsXX9NAzlryEExHlIk+e
4fHqqIlAr/HzJlI9XnWCZNJFsSM0Obqao+PZ+Crd5PqpTI3laoMIuuuuxb5pcx5O
CmgLNi3Fsuftu7/qsOOot80eQRW+hHGtS/xEz43SEWCMGkRNMTZxOUCmWErCsbH2
tefO7gLy9w++vF5gJFH1w2ywovUvG4XRPOUrdFK7kmC9DLPvinyjUduxIrOxtcrv
RaQLv5NPNCtLDqicXnNTUeUdOuv2eo/k19+LWQDk6C0y0ooKIAgQL+7GjqxK/k1N
wQqUjDA4DPWXWLZjXkJl7c5gar/+2YAOxu4m4VYrz5kiIEXc/Mra6z+GHSUwVoco
vj14VVdqgB615JVNdEXOzpEXTG8tcWsnGX+Bpa8XA7OvUUSX1W76yw4b6eAMNDVT
O3nalThycoAy/v9w0ZmsOQNqU+vmh5cXwANScyUnW9jhTZgTNC3tYQUWq9u9M3qJ
TK4ToFhp3qASEF9y7+757X/TOJa1jPqYgmhmzC6icTmWDLEJGS1Orj7v1hoFeABv
l9jeKl/OTF24zCskQ43NtVSdmiB9htHB9PbtwYJ62H/MurfH4tm/drU5GelWsLuV
n3T07CLM6FSA10KH1kwdfJ8t62UziwLmBLiYLR1wCjc8du/e5+RNc1msxT3I9Nx2
xaky99Dgr382naaBAOG9xs2hZmKmwF2ZyaGssp4wW0xPz50Gdx9YH5LbCgGF5vJ9
F2DcdN3n6qj/ZEYd6BRAjNJrVKpEgs0pdQmKodqdhtAHL/ijzwHwYND38mtErCcL
Ve9r+euJz/+zxywYX+1cwuRC/3CxlsuK769JfSEwtHz7JLwshgR5psJ1DfpOVoJW
1M2ZW7BaWtj25bxRTq1zqKfy8W5PloTTk1j8NrhKWyjheoecNcgj3hBPVxC5HVIC
AjRkqwjFjgqEHvuVlc+/Km8ZNmq/YjtP5mWWQuojp1E2wsA1L3+9Zti1epfepLFG
h6Xmyhj9NiRxKNc7lR64THD4ZDw01E4WMbOovSJ1ZmiTs/aRtEYR+UmeezVZx2JW
gLAMVgPmpCunuBqDDNFxOy+RcbofRHPYzfHdRdV3/vbuRaNsUWix+dxBdeGAULwp
Qeyveuhwqn3uT98GRaU6A0HnDVCcxJX1n+YOQofSwCLkcsr1z0Tm45Np+dUeAngQ
mzCeBLHL8F6m6OYw01eLGig+mV6wrRUG7vAirW694QTNLtou3G//oeaOlHpX5Y2+
ztznyZ1zo/XuCzTLyycuSoYeZ3q7x+fewi8VpF077jlMFfJaxF5T4BANbW01MCoG
v1HAWomRd942zmbq3hroZRaQqQUZ+6jtBPUfkAAJhISRLUfV6hK1a/nJ574fSlIQ
D03ZmjkDC0ESwcGpcCrnkTCddeIyFMLDITosqvOBVGueECZuYltj+TrysMdOzsYc
e91FOo8yQzaQ0DDhO/hwMZZWxFnxSmzPVpAx/5j4Efky3x5B9MClS/GWbrbMZL/Y
Y2fAb7aNOUXlWpWUz9KhryhiHF3iHLAmfF2JWcSJCq6hBIEInlriBG222gWtz82b
wczbH4OKvLsTTkoJkqvPykMgfLr9ReSa9Yh61+KOxbJeKTIkta9T98vdDPgOJPTg
HBuy6mnL/L4EJCgY1+GKlv0ypcT7q1OPWZF+kIoWfKbXk1xdKeCh841oiPd9+41S
woKnZrfvVDtDFaPqDObMF+HIRcfdXsPKFvhmfxqFJYnVIuOoFyQb405m3GOonre5
N+/vhuoGhRlx5Nyd6vsasTGnC6tYu9yMLYCP4f/dtfXwy++gYQZdYeQGELohCdTY
H9VRilxrZEpuMiHz88NEo3s04SxZQhqteQQLtqVO51FNDzoZDIyY3PWBhCJ1hN4y
w+hYajY/0Titin5GegPholS+ERGLOvGNmux9X3JYBzAiGUjbS7igvkJicDEotSpK
mJKOmHVjy6BIx9WOU6Pq0u8Yf7yiQ9HDtqPfvI+2EiGGbqQFro2Ne+Z8STujSV//
DtoUEZCdF9uQQ2qP+loTtIXDTD6QAcg4XMuo8ua+TBtdbWZEiX3+0VRiXi3R8/BX
RMPUCQawydoWczzAqKr7ch+RaN8WvYdvfyUGCja8qXgARmr5d5478+IuK7lGTbI1
QyEd8tQwjlkKHX+XvkzqGhvA4/+AJ0lim0ate3eYwhlXSwu3948MiuUKxU0cDkyy
2eczgxcmAf5B4Eki+NxptmvxsMoiLSK5RG7EDuWFhOa2DQ8F5SBomAf6KV+emf5S
Z11c/C4tzSdqKw2ExlOpu+5ZsHV/Bbpq9WjlgJovZvoSzh0wf1r7wNeoE3D4g00K
eFEzXiZ6x26xuSbLOmpIVhBoBZ5xbqoaHBGYgrf/OHNacPiz/hX9zEbas7lX+vZb
iIdWnrrUZfuhq1+97UVe0pLyWFNEKLl+DGf/pZoxtdgtoUo9nufQ60JLC/9qQUGE
/cCdBZnDK3j6jLhbUdr53iu2LEue+/OI8uF+arlNZs5URd1qB6Bb1Fwgzfu9tNni
2M7qkfnJi+tDnIox6Yn2IeztxUTLAfRTZl5vhESyMXgdQZNS6f9sMQPEZZirKWVm
C+/nHmhrv5t+8dosjxwdASgH5mu+hrKk5Lp92EUPatX0+rqR2MAAhzkeAQ7noA74
4vKKlSXk+UGrxtkOcbHLQwtXCs/SI4iT3IUckEkPHNTtkfDXiluaQDnAKbqpuVcc
Ei/x7OtvKJtfZv3i5+cvNF54kEnQ4vnRPjZuLe5mJYGL/5285UxpulokDAAYsW4T
DcUVdggM5AHZqrACzSjPmTno3mS8mZ5RXWVuz6TJD3M0/Cahm8dkjVAiBPHLnDRW
Wjbx57f1przB4UTLskK6NfjD7z44zxSMQ3B4MxwAKldKXhbHtjsapDfphAyplaLE
GC35C2Bi/eIyJoW3moVUgIYK+gWbKoglCopzEOmVNBCAPUK7oiVYJoKJR+zu6SjM
eg3MXlqxsRWhTJ+KaHPNSWJZZsQKrS9u8c8ujN1Oq6leM7XptBmbu/JoMyYhepaN
mpPrvPYOIxvix0qsXXG8OSxcblKRXGURsncw/7M9p9BNWczBPq0zh2Ukwg1XawVo
V7rXZTxPo8GMoLZ5JhuZsdMLAsXPEA2hQ8s4LpoUuarjr7KjN4/2j3r+pQ7ZCitt
8ffdU3T3hwIPwzLYBqhncWwM8VSyJOGwAO1BECxg896YsoCo8An2686CgtCSoWAF
pmYOdeOm+jqGHh1z36bsA+K7Hep/a/adJc7RL7xhAEOetiAxMBd+QId0kKF/lhrO
hI+dD1MqSK0UU6afEummGPLMGlAAKE8lQVgPQ7zBIcqiIsB98GRBbHpH0GWgdylX
4Ewtcf9MXSHsv7UK+HrWp76EH18E5uC8bFjeBksUIHzd4zNjQaRC2cvAgvM7p+i6
nNvxtfTGw8IzcGfIG6i2yn+0rehKs4zpw3CmRo0zOKHGagNgjeL4Of945wtADzqw
XDwKwq4vMklHFSfrzuO/JJvARgtjnSjfFLYmuN0BG5JGslyaY8IU3BCnZnRHqsaY
rFYjoWIM2Yud0Bi9IdS0fvJUshUl3+NvX82yT4Mwfg4gVQACLCXb7Fl3mUi/uEmH
nUoBlCLk8k5VQfUpWbO+09VjmG2ls+pI65HP8OvkebN4OjIo2Ym4LJHA/KjG0O0l
3Jt5yy2cufmUPC6ho0Gpec6jWCU+saxFdomwIJyRtaw2KVx/u8aX0pd4rclpD1zr
LDro+qyY1eBug/2QsYTYrrfXkBkDQQev7LZCMkVRxpBGX+S8WphbqGWywAQBrsGh
mVVYintCG3OiaOx9+faRAgmYT6KnD7U4k6Z50HmBHy2LuFw/OPnWpfoCH6Rg4Nc8
frMpAvAW2O3Ru55eXhpXUS+ZGKBOqEi7LPi9KjacD2s8ml8q8eWmn5xK4eVcDzoP
N71VewpmbcOAtRtQ9p/yYXjNFNs87jjmq9Iev54EI04LcUrZTQdgpE1VbxaRSf1s
aPnC6isIv7un5Egb3htO9yMUGh5A13sd01B5WDbBiA0SEYrFZgPgHElwq13WCtSz
llNkSKa9ha/xAVRbELJVcoUAzBgXoGnyrpnx65vr6VFaUg4b/sMm/HfopJPCB5Jh
JuF8JIySwWciQ/9Pdc8ykzgaLS7vxBWNb2FRXIjHdEj0UirTIt8TKqY2oki7Aw/a
n9NJWVo3Ku7GEL5xQ3DRhZtmD67GHRv3Wf840az9+G9hK8yDpY1Fjs+wNASHiaDE
ZgHOXOfhaefaDSIdBCkU5HhUkIKrYq1lJMPw3Pcufude4ilcPzCQEV4i/PE/nA0a
dW40xds2TfxvSPcpZLoSDiomPUhpCwl022YPEe2PQQFVU4wZo/ZhOrDAuSJSU2S9
5g0zuQORhAS887AGlPoSIlLZW27ANmrBygxRnjId6xy4ltU1/5ahxQWQwsaQ+Hju
wTDU52lPp3Ay9JFLluOGxzkuGJTkCrmK6ZA9Tjf/Ydq0/9ChvFABkP9uOy3YiMty
zTAUVGRAZoqx/qtl8XLw18flRzWQ3hFsIBS2GDnSTc205Zx3+NHHz7drroRihkmB
4Xi/X3LvIKCw6odaPf1TyjZBC/9jNjPEXqZB08GoNDLgt8Gtx/9tF2BoHLfQna6e
uzvvR4QXTJKkOwmW926/opef4rbz3bPGRLSC0p7NJgYPWvHKgNqpQZUpIytb4lIE
/TpbPeFTNQYBMvzqg0KoBL7Zq2Tpwxi0x9V+74+nwkTYCVuC01TFvG8RoyX9ZXoR
UNwBrrCojjd3YulZWMFCPBqTvkcZ1TTIObtpiBqA5VxrKNC29BW0p/H1I3Ft9XcP
AVXlwBVhFma7i1bewu+kEEyhkm+yNUlgs/6uwiAGNuAMyBJtabOwp9bliP5rSImr
wc3p6TmIek44H5AxcZBfM9byHtryG4F4qwoQJ/Eik4+CZoXhE+pXtNPxUpgLQWOA
pF7G7wu8wPVIatify+ZIiHe6W6KdZyxMtC7hSUdE0J33py/OYXoXRs/33we1j6hI
+SSEpU1NAbUX83SdjIU2S2OVHYHO2OvJ1oUp70fgpEftxyv0LQ6OSPbVInNX4Vqp
IX4YorA3slMuYGkLVfh53K+pQVceSxKxwly7cOVMu+GGOypPwqsDf/XKB1K8kZwc
cGvNvrMNjOBf5peH2McizHlte/kc0gs/tLMAxHV+gx16mzUQUAHQ6L7jZPFTF7ce
n+iGDYaaVVLxh+xsjegoI2QNnIC1XXmTIxTDaC8zU64r4XE8Q0+tZLYmH2Kh/96Q
U5aON6cw7nQLisHEM6xVxiTIDGkMyq5jKD/TO9GvKS/rxBtlZmd+54CgX7c76TRY
Dp6pl+aOr7pfzYGkbos9+elV3n1TIiMqI2m3x1BjLhbhlwHLhjXC11FO/tQ6Un+c
opE7dcw3CT1cb7Gt+GnLzMRatQWZRRg+qotx4m4HtwdmwaeMCKnVju8taATzN5uq
LENv+yl6qYZuYNDQ8nMNYmlWPZn2ujP20HjoZjok850lxcZWV/ew42ov+oTVP6XM
G9S7xm0Ukn7WSGhZoUaIlKHr+1yrH3NFWx28dzlliW6bYxSLWpgec0dXHPRVhG3l
CvLWg/e8JSD2U+yhl0s46HfAAFvWfY7wup9foacYGRTGShGzRGM7Bp9+xFbZgPwa
kZwE13t5mQN3+zRMFhGATB6aq+vPFpLAFilCH6H4C0XIFlv1NI6rnab2nzhko2hs
TDMw2VZOp5y1emULcTS2gX+KNkucypjaM1uIs1jRdD80AJdWHvVREn3SJpnq79Of
cot8EU7N0sD30DOMP4rd9dDwL7bHEuZVn0Ge5CPU8H0OovQ1XWzsMtiGaadgldCP
4zyNTWQAQrhpI0Y2nCvDLlOtoZiyfpX3hzaXpjdLYe5qqLK8+XRRWQ3xIIVvNzqM
uloroSfKzjkzqgKOjGzDmULUuwMlNjqp0E7iN0JdAiPsFjt7sYVFX1RaQ7Se03vM
oLp6Zo9ou5aKbb1rGwUyxiEkKFOd6xrajm17i9ya8MZPB2jnSocjXOcL3w6agSyW
YYjTw2MnF7MOGau6A7sQlkUWqRYfDvHSc1tzQ6qbnS22wbSBXC1xeXxrlchmnUIZ
XS8w3Sg8m4X067+MZDfRXldQpSCdkh03IOhTSTSGL7snkz8BXgUMPTxItsr/WNOk
31IgrO0q5vJYoZG7JTeE4ZTUrwovINyLV/683MVk3GCua0/Su3NT866XwPq2IiX2
p6TCjs0JfpBt8rvTw923b7jZuyzBaalV4GTMBXt5UC/BzxMR21B2bQFU0HcTHJ4G
ERxHsTf7tOCU6Nigr8Df4KSi3YUXT9PdaYNEoV9AhBd1fJDF+UEHuFdQERaGCEwB
HnHZxXhJUopHluKMRMx5tMWQeBM/nEurgIf6w+3x8llwUoMay5f/uynqLuJUYBLx
Ua/KXVkxYL+XB4KE4Yn7PdxhSHW7jkkMDQr0L6CwC7TBJGgNL1WsSH8aCPBYL8RB
DuEE/mKNkxOV8ZhP2iMo/UNFmC7+L6N2P1rzFOURKPH/1Hd2hwfQyyn22IXlnTQ4
4H42hc4JJnDgRQ/aIfnO/520K/IYj9IKBdJfR4T5ymwuCT+Vrxy/EfjL0Iv4TCWc
JaMyHD3OUhSx0A4iPLQ50PZEbqZNYZepdF1Cyo4VFJuxDFMJsSF/k1LQ6Q6sSuY/
B+B3EoRrZneqFNzDMKvEBK45Kob1cT/zwrbshEDqm7PIrhcanLPexfGubr4nxJiD
clO9og+5oOpVNr1fIP3YmsU5WOjVsoWUoqwLD9gpZBfCPVToZFH0PHfjARMEk6i+
eumvZ0odQ0A88RdFH747xZIi762Zh1T2TOW/ArvtD+8CksV76ahH8szqLVu5olmJ
LcHJe5NJ+KnE+GruIgM11JPcd8dhFRc8PLhyggKNqNVCvlUfc6nYU+5/yGbRzPbX
WKggkv10YNU0bnTKNnPqLUFlk7GWKVxZLiOFYvuA2CAGlWt+nMmNEameuYmYHb+v
8zJDAb2dTItor3hgk0Ibe92EGWrY0yhY9eKPUREIsWCOwlGv7rab6hyA3IVjbgHQ
jOhZ67iUlChHSsWwwdHcjLSJG5VifGi4GlOc+fcukmsjUEWPdDf1N5QKV30OlrGd
FevRuh7IHxSSbR8QABaMGvtc+jqn0sBaKA9Oso7USAKiA9OsFQfRwtJTbnbdWQT4
vdkuyXoatT+Q+KM1Qr9zSBr6PXtolqw4giutN10V1pCQcSumATxrKBGXoDYlaoDu
O066YCaqDbccL1NsTS7EftYyvTeZcb10rrj72mmyusy8Q4+3Bh+A8M0ieFiXItqy
Uxis5JeFKfvpQjHX/kkUTBOtvk69qA0dYQ74wqOONHUkz/2ln7G5rFkIeh/4Z2pC
jGgC4Z05Kce0dS/cyTxQDceC542Lf+QiwknY9UE8JZ6mn4pNKOmxbryYU9n0dEVC
3o+ry0J0kzuYT5nRQRhsSMKJLORUcTWXbU3JbY/E6qinJ6Gf8YOZ4J0pYkCBU3S5
EOYznY9vPE2U40KDARb/zc8mV4JPdxexgb816B73PHxb2Dn9FTl0vJ3/asrj2xwZ
8xOtj+THSo9hOWoOrYwgksW1pk/m9jgED2+p7xwwgbwszldU8xasBbJxdJ1ze9pk
ThsmFeo17n11EV+OeaQ9KKOMAubZgzIwve+Ih4y1YpXqF+Eztyu06I0KggqkxiT+
ISTgPQrGMKFSfOrolXy2z92RTaC6wz0YiCMdyIfC1FUgRo0xUmpvD03MmTgTiDAi
jP37AjjRFd0OzX/uoDgqqMlcAyFCoa3HiQuWb8NUzvdCqlFnYMkTQz8xCIK/kvC8
vvmsxZXq5O2tELmzenG/kafm+c4uWUNDPZk8aEGz/zg4GsABm/7653s6e29EdaVQ
W5di/okVg42ZP8TYuaQvGMCi5+NV6qktd7i+undcKvAtJT1yEt/7is5lXttNpk4Q
tMGtN/+B8y75lvhMgYWSJAp2p9PloaO2yTKXVcSjGhtNyCu6mjagohtqQIgVrpXP
22wAI0aRMr0Yobpm9W4M6lwcxFFJ6HRSC5OXlOVZHMC4C+m94rNV4QumJ+7HfA2L
RGC4VOwdvBk7NNejYwMse30VIbtE0APaZmRA+XKxVxBfaTLSoRklsl6IXdyVz+/Q
Lbtcn316MiWIDDacuodRLTSGdyHXt8xW0yZjKwgRBCtLE8gSuejkasAJ9dgvbVQs
1Dsh3F1GF84kNxDYI1vKTc1S7InQOPAmYz6Zpq6qAe+1g3+0TpvLwrF1Qk3I2/WC
jW2wUFSGIxD3PxZGoMx9a/nH8XhJo3yWNIQ42UKe/NJ7zuxdOjZiLiiv8gNwMUZI
o9HW2nqJF26zyHkk1gLMtqOfoQn2cYKnohr948JP44H0uj5mRXgiD7gXZMsimT08
XDiWPWIIrw3f53pb04LT31W+x0BfiETk/bW5IA8iyXob02mUG+f0DZGhRkOmPVyr
71XKjX9zvM3aaQHCfXLddHy3f/ZPaUXvrgj6lRxokSL/McWct1a+Yt2wfQdWloOc
RxMBCg/tqrguKndDj1GtOu0oGwLm+64BMG91RCLJhVx6/gcRUaUE1dv5s2kK8dH7
joz8oMEhUa0CtDYCELPjLmnae/eT0Cp6mVpDQIMQWDPDd+cOizQTo2t+ii/aRFyn
0wTYyrHCRJNIIgOglpeJJYw6Ov5ioOjzFAX+7wOLMpDzYxnT8dA//VbtY3TsBWku
6Gc76iRB6Xvu5/qLWIp51gJEsp14xZ6Z/bxT4OMl0+rJj2N+58Xluas1BnfazkSk
3jWA4pVp+u1IVVm7kvQJ9RaSeCi8UL9x0IoAbAHmFGrSiF+qTyL49pOd5sV3063l
xLFKxNwh3Gx4SLr3liJrUaQ0nFAuGKh43iqCeV1RgBJryuth4rdceDEjXEmMU+LD
ZTW6R8xhIQlGaW2JNbEA5OPziWXLkrAgVZ0iR1GEOH2SxjabDh2vdU4gGoYk8LIR
bthadb5DRadS8GpDLz2SsI6wOxa+SOw3BMp+KdBr2h2A3Qk0d+H+g1lOvGkO0pIq
+pnVacSYw95sWMOu40xF30Ra7jtqcLArAfn6FmkAqsRWnBvU8tmtQLvlpVz3l50Z
jftFOPsU5H09gERqlabV1cE/56tfYle7qlWBcSfbmLBVs2eNTeUD5PpofnKRjMxp
mRHhacHRJ6VCKZTq4hvhAcW4wXtIm9AhVBoWObf0Ey50Hfjw8vHII9zPA1WQNmHi
joqlkr9kEVbvoxHsQWY39rLGdProwKhCM0dYLxxIk2h4WIWaJWA7riELImZw9Bls
zZOzIYwn3aGC3k9K/8ph9c6/adpMmG94cTxAROsy2JQZdFZPG0TXzTC6rW2qf+wL
kfWN/TwtkdErD5atOfEf8VQ8fa3Mh/CO1oQMCag2Up+Q49zPDlxzs5UYM1AUJv9X
ZD/85lR5laad+fdCnAAuCrfE+dQl/SgmozT0yLGuaXfOQapMGVfYqumKH0C3e1o5
PBxvTbhbKeMCpxb83AfLZ8O/yiLumdG7dR0z/AaJZdeO3VipZl1KRiV2z3F+nyXL
LDfRuLtkTcDl5L+jZnMuuueLMqq1Vv+SUHNLW9utMk8iy3lHfPlrtd2KWlTkDbSG
56c8FHiTfCN+wNZKBumq1oYWpEdgJz8V//VddtqdiSpMeLcg0MNGvwoMM6DR1Qzf
0d9SxxGV21b0ERjOum18LNf9G0aPN4MyxcTkE9ITyxKaDQcGdV4xZhw+/tzQ1P5t
hp2wnxsBbafQ1qLIUQ7Aie3ZcVlSKsWU7OwY5IdMSR/JzmbhW374WZ29UxgszdMI
oOcTeWIY4yzoXd6SWr2N2aSyNpbgZX/dgDheQ1TR/FHX0ltdcIqJ+P3Eotl0Iz2+
JVVH75KehYelYYzmTUzkzs3nG6ywCofylvTua/bpel/iV4vyVGyWehQonOD1wqb/
h1vVpS4bAKlbSsp5RMyGzx9zJDg8rqtkYz2VDWSA0awQw/afkmBmWH+VMsvEie5/
WTOXiqhBb0+tTc0XnXU3uGCw63Frq97mazwO8I+CT1uyJrHPMAzjX6nnI4j9bH2S
MGVMH/x8ZnsmU+Z6uzYeAuZOAUVR5i9GairYTNBKMchMVSMzriuWxorG7eNJx2Of
QudqWUL0tas/onRD0271ll3SJDjHv0J68r/COx3GD5vbDxNnEuRwV5n61X4tt0Os
CkFmjOHgLQ9ypylDhCW+sfIYAmUsANsX7bD672u3kCf/MtJ8SF+zwYMi4y2/AlZx
1iyMdRsaQd3KqUpwdELe/addfHGAvTib/qLUkKkyd3uBjcYjlWxUwKdD/QRVvpF+
D0QGWmTibBVZdmNpJctgu0gsnBf01ZsL5PYhP/ORkgg+PtH+ulmBxSdoqxFHXwOr
5LYz97YZYHvqIPL4iMAdWXqPuIpor2n4RqKiw/+Md5toEHyY3XHmF14Wo1FSDtLb
NKftp5ySvlKP/v9dNGx6k3SwKUC72H/36bM/ZON7oDlT75YHj6QmTFE/1q/Ixmox
EiAl1bbbYaAl6Ei/IhjKTpm95eMfoARnv7bprgxRPmiFaEYZhmSMw1v1yh0YnS0J
5RPIkr+4AAGojJZ+YngN4hKhenmHVnQ+AIxW/cAbqgOsj9VAhDGyH5VFsSb4Fkp3
IwXjbEhUIMduXFljAz9VCHNkp1N/G6sQNVqE561M3rHDGbp6q7+AAk1Dhc+m2iLx
xKk4XXFz5ihqSyRGD19xngBSi6A2oM+XdemIlm97fOiJpCjDhEWIcXKk366PGyO7
7A0MKwnXNJvdmUfOOpUUiutwJEufK7U9q+7+QMFEYclRU0QWLOs93b0QTT5vURiW
76Kg35fo5SfL9jAzFTp2SCSCPUO/PSfGPS8DfKfWiiQiQNqNsl+MFx0Th5ofKFRO
XYSy9luPIf0UquESPSWgmccj6bKKg9dET9k/XzbJNK4QGaS4XjtR7hMyZGG+KE76
zxTdLMX5Yc/jQ4WC2mqMQC6jL3YL4/fmwrEFdQHgqVO2+sWKrsXSfl6eYNgTbm4Y
gBJr4sXx9qDKkUV9J+T1XNbk3oBdUL4F14a7I/skXW9lwe7Vs+37W8/6YuBGn3eX
wxN2VFYTH1hymCtTIsqr1YtWfPk/xWghuKL1XfMxoyNxaKkyOyr4ovnBmVNGIQ7e
EI+ycHdSPzZ/WobmVYSGTXUZHQzqiINC1cXKagEzoyfWJBWw5QQrQOWPKWhUopI7
8ld35oRlnpplSXKckvnR4o6n75K8GRLgRqlfSY7sOHo+JZF9k/Je8wNx5ogV9F1O
iDiH5vHGFADFohkPrWIS8eLyxrXfIaoULfKxnURO7DpOfolV2spHy+xSdeFrwkgD
NsH0N8RHqehN9aGHr64wNrmmZzsXO7Pu22icAGJnk3BjHQ4Hj4cbUTme6DKmWiyy
8/fKRp6LbJP3QzOHGsZMlWPEMizKzhnFxHulQg475wZsnnhwuY9Ww59/XQphv66/
5CLcRE3AqA6WanCYb1kk+gEegRlbu41S9Gceo5GY0hrn0wgBMNgRUKnH+X/DvI//
jY57ahjRHsp8KqxGGWuNFXplyoP+moMDtHUZVzoKJgwH2UKVv005RKP79BOjKoE/
W4EidbIAj18lTfBj2lqMnPXH/w/UJ9/APpXU+GFxusrfvXFQiNA9E2mbbTiUuTt3
SToDULeyUdJ6DnHuphyYrP4V1VkqRElcx23j/ZR6d7BbwLG58mKt40XsmY+7QiKg
dPEjS5zVq9TwJ6r8H0ymprt57f8+Wm4oZCypmGydwtT/VIeg33fejHdAYZ0c4l65
DplQDYOlqZr8aIf2khAIP6atV+Jf3IV7HdiIeeV0PDv1it8ZupUmvYfmFnCR2lTH
YwsmQSYG3gYw6NnfhrL6R1b+XvY2WlLXd5sS/IjDf5tnaqTJ0OjjORGbws8nz714
jAVR5/YSaeStD5qHYdAz5iF2MdYD9usmsb+oDpkd4/2e3/sxo68ecduGpBAGeaOJ
+tFC5M0WU1JcA89qa4wIf/C+SUpyDMtGsugQFPl0ZkxQsOow0RqKiIK1aykZIiye
7oxohYbrLNAcIlEKzcVTjO0QxpY459a9J+wpHugmvMsNjDM5etx7vBfyzOR64A5i
7phzgI5DSimNMLYV6ckw9H0HB9X1/uoAArsGReC0fEKS+MfD9nFZtPZ41fPSPEDa
4o/cCjVBll+k6EVxAo/kBCAXrFfRC3nhn7E3H1/zfIW+hm4fcxxHpVRTRD4ana4E
GDLSWH575MUI/336BH0gVhcEyswC8aCk6KqVP67NlF1seJgnyIYz+iaCb+RgY074
OkwOeowB/LEbjkdUcC0aOFjNfeashZqGKcOkDt9DULyqEkpobPqCPnKtRTCX54AW
J4hP8jgmqdcjcDr9L22TxuCIiqNy6mye5BMCopqGAqtiTeZpxtNGVkv66m8Hgn2j
ooaPH31bK0kp35O0Yr1DTrHLODbHPle+oJ/m8cPYLpLn9zq3IOXWgdJmLixfauOJ
OZO0euF2VJZf8oVfXIh4sWZUtloki4pIhPTeLAmxpW1gpZg8Z96pm94shaX+54+O
VgFRMa8nzFKY5fWu820+2FC6V87v9ztLLJrmQ1mwbjQv1rcIyKe6NTttARhVPbMt
9t+SL93TMwL8ujBDDqL6oHFt5aJHJQyS+gY0kUFA8h/+mxxi69gZwQ0sdErYNmkr
3MmqqEhS+RemTyFWnavAYQag9All06o8zG4nKSQk2uO9/+JVu5dkP9lvgp3KfGdb
irlqOcSG5uSB33l6ph19kmFyJqkOFglLJUxQvHWdP4K8HzYETsqndkziln5WAoXc
ChN/yH9r2G/Tc41VIhf7m608L29iPMr7chfbiGEdDOH4+H7u3kTjjYWpZZWhmfJH
MIjceEZPxu9tu9bQxRzjGr437thv8qPznaX1qoqHstAL4lCMf4j7yRBlXdkDhIXU
8YEygME+t39NoeF9ugVa0ULmD/NLBHAQk7fhMfsAPdD8Ny35D01MaOLypvDtFRQW
Gn/Wnw8tn2fRo2HXb3o3X1TZAaOVyfIby+aChqQLb7uohHpHCiyB22+SWj1fLZIP
Nep/6bztxB0RpCjohVjDaA9xa+g0AuY6pXvdHJqwm8pFkyrBH96zWB9/hNV5N74M
M5B6WJZM4ge33FXx1nHag0bajn4Pw0yQ7Wa6S7HXfIKgL6y7oL3/mt84Rcn1nUOT
KCNxhmpTgw3Eiyq7I80BodSEDu/LgD+C5aSj57R1d1N9agjqh1KcQijaX05q3lQ2
CnNfmBorq3BEMK8fS9I2ZW3AsoKL+alUybfS4B5/Jipuu0Zm/LSDrcLeqFXhXSlq
JyUOLr15MxmBAhFqgjpTtHGeEoFxHwJy75gaAPOwyVhHohMc+lVga1zjSMnbkKxb
mOvPXnqB5QhQU1YGDRG14IfkUSfLZ7r/rUPuyqXgtytz7ZyY5L7uoPTbozZo1FXC
GIPCGgIuq65Fp18vop+YVESAmpDx85rDFVCbjoqjXc/sWPelI05mS/gjGaUUKJg0
mQbcIRdD+ym4QH0ogSwUfDnyJ8twL2AEGnk0AseE0hAfowpZjSr1x0zHnIOPc9rk
sm5tgVjpkCYDV1SSNktubdIIU98CUnm9u9cOXW+TRgfFp8qI4DfU/6LEDXEF/eO0
xTEaeVt14cJLPST5xRdfT/ZnP8Cb76h71dtOuFZwgyepwAtvan6VtwOpXgXu6mUX
f+jfs0u0EMPdgF58VVVnEW1ERQBSyMyifB19fTTn/p2ZDIbtWQ+urvYefVyO9GUO
OpTJoyS2U0r1d6Orfo4DvGgcGWiXYdbjjtcTde9a5xGVcJyHA4mGdgk26xKZ7w+n
5mWMpR+Xu8pGT3pIJtmM/o/aMzvU/q+8eXV9WuKsS4Tt7bNShQZJ/8y8G4nsB2KH
l9+cx4a021xIBgrn/szzzB5/QOkTubm0VYN22S75Tmb63SZNe6G0FvOumMnxE9jL
T+sbZaR682dTDijcdKGG+X3pRb/aw66jdmJuAHGh2IaNFKqUAt/uJupzgYAri87P
cQEoSbeTme4JguYs+WpIInhzRK4+OG7JghJnHP7JFR3tAzeTwmgroLcHbghAGclM
mDqz+hVWoPiZTQVrOiMvhmhFWr5xEWrEuXWUj/zR1EYTGdNCTNzfUQCls58tHr5u
H9U2ZvC37iMktOYT+M4oRiUpRZAu11RzmJ3wsmSkBIPATfxF4TUAa8p46CKbVVk9
PDYu72z6pxITFbG7oa1+elWCFImgBqmO+KxrVCbR31FTE9jO/AoTArHG7PU1jLCE
li3NOL2tDbectoPXv3PEVbCx3LXE9cFiIX5g8Y2zH0G3n2//Pdl0Bsz+7GzJcoK3
TjquDyb20ACPVuxiKE1d4txLzdI9021JQ1YNF/hhPJScfgxbdXGERigPFQ/UKH6J
lw61pUYKNXrAhdWrM+GZ/FnWqmrDIkdDND96qhvCBHzcaJgcOa8+E4pZJHP7VVkF
58NJBPyrZ00W9tU1Di6t30wWVhsc2GvnwHHPBryAX/v3JpmmnZraZh1gHz6MTwJx
YgLzV0zttP6cFj0LCmLqwv1OGZw3gm2D6OFut0z5AlZnolnzjFmsxJpF7c0sjd3I
ssRpOuS9eCJN31ZG2GKiyT4fT7KzFGnV4I3mVVajk6Z26EDdFDyVuX/Lw7UlOnJ2
7RifvNk8uO/TM8ZsxicdO4nJYEbJF6DhnmKGCBsgNtt6qMjNuirBmaMlEW6a28ls
/z7qADFLc8zt30ekyvsF/yq6FDRK+Ox84BUKnEs3SvixT7O9Du5em7pZj0b4xgzZ
c+hYiN+XC/4UF8+0qNictWH2ZgQB4Siqx4I29MThUzy+M/8QiUwA/MjodYhch3r2
ZEACSnh+ifdwk5rlAf+gaQYTkBMGuZli8UmYG63XIkc6+0YcqI9oh/S9LHSdbBC8
bKYbmTxtxAQE+eJrMrxE9KQX+QLHKxss400WunV8yUQNJ4sueE6EhwbyYYTkD3XV
7qKimu0NlnJSfYjPk3u2QhFWol+o4piZqVU3NY8CDdOKqDJ32vwPME8tisKrMh2l
9K3RihKLE8j0wqkI2ohFUhcVaHyIZllPitSWe/o6a8dWS1F7cWAuy36JVl1ytwdn
EvCJy9sqOAUCcMkFkn5vAVxi+JFDhqReuj35gn0+YjNKp0eArrwQI5lo5FMs2id/
PFWowb+0quZy97BpuMQVRATUBQShpsm6IYcYVWku2fCmlf3S8NouU696TGoeFSZ1
XXC3Ul0l2JUhutzlsktKH851Ifu01UPBICWY+8ndxZWEAwMMV6IW2Bco9lSuijqT
NCL1J2CVXGsauXleIVx5l3x71B+R4Enng2zj1YSCdGotjHxWTrqz9Gg7bidpC/5x
TVVI9VssBmJ1RgY9wf4DwG9dqBhfYr/xTd5oLo+v0D5v7H/mcYu1FjxgMUDZl68a
yYeE243BUCDPW9IbXwucxVUs2ZBInni9nXhNNt8S3kPGWbgajzce4eZln8aDc6AV
AYNGT/tymO/hGys4jXSxkpqN8nMz2bempVn0NoV8bA0XSeTzmos+HJaiHOx5VB5c
5EJZp2xgeWbCiAmgTHvUuODBP+pbY0fkUk/ZVDw7drAa3e8OSCdAN3awgOlkm/Ji
Xzzz/17nmq+E9SSTeF61veZxSQn8QsNdSRB+raFLQM8sRWcZSXroE+EbJ3lV3FvB
AjRFVKnIePLusBYRWG9cBiv9XXw1HjhHMr9xxqeK0BldJ3zc68mLRCCm5jRfY1Zt
Nubyd7QhgE7G9Hwj6IGWbVNPWsoDno2QoE+xICVho6SZ8X8jNmxobo1fs2Ez6/Eq
TU1RYnzMdF7hVzn/0I6M6Y7JFu6TWCrw6np0trpsVXRo8shIrHXkNACTwcikiMmk
OctQDGRGbbquFU7DTMyYwNm2OSCrgtQYo+woBHmgK1T7HyOQiy7DjzfTANzVC51o
5sU8fXe/P4R0/GnUTqGx207jUTK1YJFERKFtHwsKgf1vHpPRgOodglfHr19gu9X5
YAG+E+tQ2VgwNiwlUXEG6dqutM2JGwlDv9asYQa+u2F2MDq4OnIANqoJjpurDN2R
3T8ufHxfHDgVqR8YWES4zOPdHQLVSietxaHkhcfMHcdqAs7GZ5PhXHFmcEVgk1Px
DakTDAuy323FDuAkY+eit9SpyXDN0o9aAUiUY0Q9BJWDK2OJjv2gEUYRuvp2ZERF
LRmXxpoEQTg6aLNgkjPVRs7n9z1vRV80uvGjr6yNg4+YyneACmtvww1Wq4ZqNUmR
lUIo4n68JplSTs+Fy2kw2QCUFJ0teintnTt+jJ913uZ74Dhr6GNPypQ44NhVFRK0
qdHIgkPFSusrmUvPo8/r7JQGQKcb7M0Y1GwNpStKQEFRWV8L60VTxM0HRhbPvix8
kc+yvHG4t4EjQ77kB918aahzCR0b40SsHm6cajkgki3kfdLRHOZO7YNF0T5dCd8Z
58oUcaBVEu4bkQmGktg5n+Z/1CZ/V6b5YkIQ9yrpsyutY4SWp0g0+ceI23ZmANdd
5+2nxz2MlJXBorBdw2uOT0o15QtEC/apzIs74/qPbG0dRE3OUDBeDl33Zhq2nDZR
+0C0FsqcyJ8P6quomNlp13uVmN32MjrVFsO4J9xqsQq4vYbrgDuBDfzEoV8X2g26
1Hg5EKESgJGb3BLEE6Q+dgJTc0QwlRiCcUaYpo294WS3sj6qa6uYxmNj+SSURzYm
JGTTvJaOKE5wClYH3pO1mzsDnjO0oxsOiqnqiSXuVrkpIot6iHS67xLyi6b7HhvA
oQ/+21CRKA9304K2yTPJxSrAgecTzqeJ41G9AM7F0VHk+RZFLLxSOvkp0Gx+7Pcv
aKrQFvLJI6psF6v2cSHkmxrlHlU46Yvo7exknag9deJE0xl6c8E+qr6HdW87C3zr
tSxUgAmoVLy03kj6hrthBOvmseETwR3AfrO+Ah1k+dgDXChh0Wv3vntYqMalzQ8o
PtU+lc66IxSInfHWDa5yr4Td4fTrGaEHAIGfx1/8iIptY0Jy5yb5QwYwiMeH/pUg
StqHHOt+BDXJmx0035wql1qayhhAr3AcTOdcklwTwMNYLGysGA4MoVuPYamwzMO1
FnH4E061WfM939gWpZbSMSmsA4StZbehfA67RSrPxpL5SE6r907mskG5nA1lF6To
sDO+VBtpgPP0MkB+erCKyfJi/J2WAR/reiKpbj31mXzQbe8wvUy8ZOudghTklIzo
HUo+tRv9QDHZBALDytZAWLSbgCKvZdkAb21fTRde1ilJhsQob9/xn4SlYQ6n7o7y
SxS3uMY7EY1aTW0vXZqNF79PbweoPBQyG/8P+TxgklemQh8cagCzMSSuMvuwyDLj
R8pbFg6amwlKMRTEjvOUDpNubtbdcIganKAO6/7cAdSr6jUozSQvJywsfSXdhEfd
iArbhLQF5i3Hp0ueFgHhQjiR5HOmaGoG9w5rwUX2MHSHZtZwcrft6RD9IqhVbY7p
CnvGMkd0eLM/wAFzyENTDrn6zkO/BIvDn39kiNUvmyFqry7f1arwK+yRyKF4ni0P
Cih8qZnWB18+uMirYZUO9KHOmnugW+DfNgVOUUl3kKWiFjxoXsfbpZXa3T0GLEWk
voDAh1qzuZPVNwOxBaXPdo/V8fyPcaSEIgpRCcZYIdTWIB8fOVArFzU5j2fnFSTb
ysqQ2z6EbkmIfnlsUcEN88psIg52kF5Nf0fP4pxQ7r/WYmv4N5akbyOmeUgJzGip
g6/NCfPRCta9m+kiA0sLlnr67MOHq1cSlEs6CZL8V5buP8hzOg0xcBoWUYrwtWdu
+vB0RJejjFPl/75fY9qilygzc/D0yEiL5XnQmLzxNwPQg/deuaU6VvDFy/MFZeD5
IUn5bwx1jLV5BlpmePSyncuiFNDUxLOusX/rDPzbP0rx6tED9WnKkYSsjVa0sx5W
hBWXmpZppC5cp+OgjzbZxX8VbJKUiEnEEN4q7q5rhSjSvrh15CUZaB7So0uUAlb4
o3NGjr5WUMlT3M6ceQJiTm5cnURszHSRX8p62DzW7RmvVJogQViltksUwfqL4Tex
Qfp9fJ9DbMySxtSWSTbB18bNbgChLAfpnTJzAN7gtCzBv0cziFJIPmHBFl8d9JdE
JMGrkmaT8Y8NoC8MkSHdJbrya5dlKNK9Fydd6Heg+5FhUEu3IYXNM+XWayqQdEHE
41aZO+1R8HO9Aifgy1I6zq82+RbZ7YZ3z2kgL4eR+2KUXrCB8j2Qqm0BzOngp6V0
mDyBNyd8jSTjYD/aqDyJTbQFJ6kiqSZhMbB3dIdFp1ii10EPqQ7oibFim5AHohdp
B0tC5fKKPSY4A3JiV/arOtKLsJk5WEM3FxmDkIpjH2CqyBmlgE65Iv5LIuXQPfS4
gLx2Jz6KteyHq+g30drcfTzQJELhNjsMMDnd7k+WHRiaO9YROCWo0qSAmIAioQVx
B8nMW5m1M9ldkDPUUcN2RG3NckXZYjMSwN6Sccew2Srxapu1gGan6rViulldH5a0
lPkJf06ph34rYKsIFDzv4tUV6inxuuQd9wp4M91+eUAR30lQ+CyuwGyHbbeIJi5D
ZOOk21JqAKVKthrv43SJlSkSSnSoZpkUIUlBYUxXNfCUz9sOZQIl1WyZE2uHFS2j
ffvlx+fLI0zlfqeS6GWzoXpYqZYL3Yee+4pB9vdAC2Z/B6HanV6moP4WNXHWURuz
9RarbWGMJ59+Jc7QJ1Di/2+NNEban4uvLC8UbBBYjPwt4VvDdjjVKyzLUAXNYnBR
up2XsdBNI9uww3Nfftt/uQD2FifkY+K98Yg4JT07yFuKAFJrSjOtdpUWkN9ZPJf9
UDQHhhx0AsxVsYHhQNxVbx32f3Uw2JaX2seFKNCPIF3Gh5JYWoHv4aX4WZn/yZ0v
leuhmkVEirYbFbyOlLNI4xJfeJcWdJEC8tRMSb1tPqj84r0kC/AG2xu6327h7MN4
xzAfbComvdilyAnIhioO6CDtf1ZJYltbb5YEbeli8h2dTY0y1Nz4MbYspiuAHC1z
QexEAoNq/VAXo2XPaOXjjZyVGlUUuqPl1Hw4agFK1AyOnfQgjIL4kbH2MeHbgJNX
DhtZZp++2G8YqI2uni3w02jbFwI1U8ft8Zvj2Jrdg7nIKYC3IFYTvg5lKr+wV5nu
H5r5NUcD8ORKowOCrSrf9ZibYd8PDM3q9eATFTzu0oRXDOkh83y9hm+qiVrn7Tx0
DT359LqrKSEe1G2Dpn4/OBbUm7G2ydTr5FQxiIS0vux6WKCJW4g0VVeOpzpv//8r
9aiJiLysUm3moTY/z4jvzDcwZQievU0E0ntdSInGJtDOA5jL5qYrrwS+bjKxbZSQ
gLvm5Dyd4mkfOVNqOgCWufmXxnKX2/lKcTV4Pav3ea/3P/2eE/ZvRshcW/9V9r8m
T/XjqxVqZeRGVRRXFPfk34y4yrqDVqW4AdncI1YktoyEnZfZXfVtVFLh0m01Past
fj0fqzEwB2T0EQJMnz6UiBivoosNeicHlLBOi63uNZnJykYeXEC6lUoQx3Fgzb5J
5xvViS8UNgpwe2nynn4HPx2wWISNO1n5dQquxEJfhqAF1H+l0B6wp8oiRib4ygFy
+KJsziTsx5ghGtW+YM3YE55o9+O9+iTGW6vWEFL6K+P5g0YMD+fKanmPn2vjmSay
La36iDO6Mp8XYnK7haNuDMdZYy+3GLYDHhsiCqbyI7pKk9tC181OW5XTYkAtGigl
0w+NRcD6ROo2naCw6wpwl5FKjopgfrYrHZfMf6hDiLeeOYDOuwBpzuLHp9VG9hg5
2Ju9tQ/vy3fJtaLsPner9ioiAmS6KOifhZN3YwSHbQuS3BR47gWCW6ok4zxQGiIB
Jdve/OHuBG5DhbgMxcPlVGlttLQxtXE6F0ijCSkQQIDM+DGEbdiKcF/ItV9gYk08
uEox3mC7VyYR+jXnLA86tf16XuYRMp5WsbnuV7jEN2ecnuVuTsLxQ6fxqC1HoPS9
2Z1ddK0bnQgyZ+66MhaWzep+zrNtdwJKCZ9D7O7CBBKuWwss7rfw3htd0vVM1mHA
6OFeoQcuAKNJRJnpng7V/WhcTqeHNp8QMWHCoaPNITKkYSIXMzRye1GogMxQ9/9j
9aAHxSwnKoDWEjR/WVocNzkyhIsUNsE4jnHWTky+0NYqdvfnH+eviOxCO7Za3gMC
NZ0bhOD6feR+dRl85iNcDVgwl10dSoBUsL5A5L6yG6w3/QvYSxZxQIgI0mpS6lQv
tkUZDCTN1AY+uh2dY2Jm08Ciyh3MgTnD7AwmhHjHAJiqlpNofQC0q95CCq3BgqA2
r6V74WVGeoZma7NSbiIH9uPps7DOPTJm0qCv0Q+5Ata6diuNd1g7zt3WVb3SGBDm
GqNkH1VYMmuH/L8RBWKudWlgPLHJ/CBQfkg83btjsWSWI60lmzE6LzEgS1qx/uDS
+3bnk7kJwKl5Fm+hOWYZk4qK/HfOXF3PjucbSx7ubcq2H66/zjw5wov1D0jUldyB
mrB01XOBqXrVEzZaHZJhONIMC/8kfJaw21KB1tpJ2bsaCd2c7mbgeo5nrIRZCktC
7Aci0b9TGWA0/nQle77cDqj+RwF7TW2j9vdf/Fn5HvK0caiw94pKGQCQ4kjNAuqn
p8Jh0xqdY/j6hACv9qT6dqy+B6Qit525e2Bk3irYKfuRjxnWWdFHIqMuJTMfmM8/
MysiVT7S/6jCxocODTYdRx3dpY5ldYBpPhnBpeqblizGwXSXlD0paOoTJVIubn9F
SY8vgqvaZrL8jpFJJD3lXx7iQ+obUsU0z4pYqNVX1v3/bz0Qi2JtFYhV82Y0RbRJ
s5hSIfxjc/NVhpm+/BxTA6G6Rm9zJfHB16Q5fYSqr7KO6eBP1WTjbseYY6LGYm+K
PqeLklSCGyCi//4RF9mhrQP3IhcqJk3mqLdCpej7usYYaqlRxfcmoUPYF5bYRv2C
zcYgT4N+xpMF7US5vZpKQLftidOVl/85eea/Sujv+9kAbUF2nynDXgMPDq3VUtgi
fQr+6xWXJU78IV9CHFQJ45GOOHYfDJ8iVsDPzP2wONXikDms9lPDTbBRJuKXd3Tp
Uu/Fs2YqN3sB1HsaQdoEFlEhwnuPS4CpuZmsiiDhvBFO1/riOrETQo1jyK4TMHOS
2PG6cSKe05lYypbxgCdfn52WfM9Si2xEKeX4jKYjZJVO18SUHVJgE2hguDVll35g
Cdk6neBLcqTcSaD2VbqZrZmNfksflcQy7vwlDuky1ZS5A1LNtsCgwriN+XiUzwT2
jYtPlqegQbhirnd2zol7O5tMwRSQsf61eiqBYQKMfPmIYkDDKn4gepZFURV+E2V7
ogOP3saUNrl3WclxDLGbPAcpIV6d4f4koDfVK0Yv4Jx5ouf4FAbO++JLfKsgNCfU
Y+4go11fAfjGqK16U5nFwG1v5Vo9bqUwbntIBtNUf52ZgnmpXxT9eyY/dEAAAWDy
wFov0E/GrR1OWph1L7TJJK7nSzrQS4uc3vTGK4Q8RExJnel6aR9N4wROS843PIiO
kyRcfdmUhATNw1HGpc3Mw5aS6MXhe2QrszwOZcEmLqsHDKWVk3f7yplTlM9LDPFK
rBR1pbP0AHzJj5Gcxah84znfh02xL+WK5egelRlFSm4iGC4YWO9IpdKww0VTuar8
v/xwyy2KxoANLF2dxzAt20xT2NC33oQvRRoJpP+tIE8=
`pragma protect end_protected
