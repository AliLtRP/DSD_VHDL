// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:16 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NmR7XHi/PSScMQ7KXt5pbe/0w1kdZ/vObh7yS682W98rsijVwl32QiE5KB7upaCs
3DmUpFUhwJJYwzBqDq3CnWhSVMYBUmlAc5QJdkJYUBnqfGRfYSqlNzfemALX9ScD
IFEmi+hakI1YbjHYne5EchGP8lqyvgrLvByaDMF95ec=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12832)
ARQC10OsrtmKdhkmCFEfzCygtt/lSlFQ2VDVF4fjASqrFcoq16UqlDnpLIUwnGhe
06L62iIJ8rhrYig6Oex5izhEg52iZ97S+akWM6qu5GL9sjxvUILFXr+I1xmrazZv
jN57y5NSeQw4UDS9C/GPQCJVSxWTUhHU17WgLlVegTHi3HLNElS58SN4bcvRn+GO
4DS2c4JE1q1I60acI17yIW5+9yAjF67iUgAL2jH8vPSzEZAEpbK7hNbp8Pn0lk7O
+OJkdPP3FfKZUwIBR1sW9sQFGkiho7NBc/a0fpGH8u/f+FToxKUPryveshc9gtyD
k5u6yMx5eAgBmvF+jV9PoPJBbdzBNJWGStcF5G0zFHHWm5oValqZvfFMuf5gdBR/
zXR5FdxsNChueywgL1P8Q6nRWrg0nAjFjBT6GQjK/B1GW9akTUyNeUvWNkhb9FbO
yFtE4iDWPxjo3wYQCm2pOFBV24v1CTkppUJzQ8pfe0bfa0Pug45KfLQJE593dhH2
lkY3Cz6TOikAjuseGwN9D0EwnPxfZpqWAT0ycrGdaS3RTRUJF44hRShwFNona7On
Du6BJ44gKBQmIGOFWRL86Z4NG19LScde/F60qEDCdZTjvWD9DpRY4slJ3purvREt
PQp6NWM6Gb1CT+8vGHx2CmIW73w6UFwjg7F4ckye03ZoFiNHDRN2KrLrKhzSQ4oi
QuApqujBoUkyHOkzMRYJ5hNt0gJrRvhK2JH5SxBDFe8L2/nYQchmqa2wd0dICPLs
g/jNGOYo+Vf3aGSDW3LqABLu8KEwG293fHsTLnpuSxQuDRbiN9FubmatnDXK6h9W
eZa9sw/U/lz8wVgszpr2kCFrHruEUmmrIjM2XTO87QlK//RFNshQOooXSf0UQsqg
VNRHBoKyHD2ZOc+pqS2HLRf3hik4TQjXnTcLV5DTdLIK8jKXiNGRgO+EaGQZgLup
6rysHoeiFRSdBb/gr4PcPx/im6XImpQBYS6KhV2XWT8TFFIOvNYOEXU8OGFxJgbC
F0uIZ18DgAIqO35EJWuyUqXMwz0ACe34xaOgt0qLub4dhoA97LAoEVZhzHA4Esdw
TpAHFbJ7CwNTsjpwiX67jKG9JKJ0/hgljj6lywVtrtvPGia+pCjWC9VQe7WACMHp
D3UNhsb9VQ61rXsTO7yWLMaw3gKssfGdGAeIscXh2N5iabqUF57po6y0gjqNyLKP
wqASstKgc30NhF4+SikbiMSo0r7q4vpP7PWYa/5rhZf7/zCJO1dOYsh0zjlbMp89
a9QvN6A554kxH2zH/z4552QR3/TUQ7aITdIEJnCa4bf0T1tcbWmkOj6wTlSFTO8b
IlvUr1mFsDlTGDt/VLr85tLs6M11HWcsLKcZdiAgnW6yTabdF9EpfWbqZa+J9cd1
f7imKtqsBcvWw8yCYhB3ZtgDbBF3CRP6169726YipKOP24jSmcn1s2DspG5YOIoJ
9z68PFKaIIl6enkLOqFJaiDv5+es+TCV7yBbXOC2Lzws1oH36DJd/sinBiliN09C
hV8miXVUwx361lr6YAyEm+8958UzFEbX7gB7lCTbWTSgvkWJb+lU8LWo78/n5a2y
YpTohDSLvj1E6M8UuJ9KgQKV/72n9QFMFnDLq5oNk8mJVzJU8V/Nit0Ozp31WOG9
6SB+tulNYx6Vf2uCY+12Bn6zPXrf1Q8SY/sl379qE7BA5wpxT6nIGaIxMQ1dWLy4
TZ7H7c8cdi9zp18EeotpEk02sFrGGVjNKDn5hObaXDAGNChKIxO2ebr3hhYhR/ja
vwuauyJLIjpCgyv9NVAwBWri6hDedNCDFV6gxUCVX2R4DU4kVu/p83PohG9c9F2Y
SXfDqm49yWtNO0i+5GYwrDAdnEO/WEEkCITl18vNOAMs0rL2lZXOxcPRd8kI4DAz
9otDsXWL+86WND3YWQemwWUyzG/L3MxOY8DdZYNIKV5QCQammhiH4PHGD+Q8HpSt
flmsNmqTbrrmH4zy7/7cp2pdRT7aMikGSLLmacoie7EApBRLGbr9NQnwHM+BLkAF
3+tfmytXLBsEm0+uSifjpEigTb/QB7K7MfwfxzhlDHCjhOKvL1QPhmAEbavSFMKm
3j6aoYylpbnIhtFQSvDsC9CsOoc0JVossk7ZCFpkSTLOhVvbMqy9qkunkD/RozVr
XCLbb1t0VrIPByiHsXczxOJu0HYoFf3zeen/tlrxiTXMZgXXSVSNAk5lKPuHjOcE
7INhnF+RqeZIblmWjaZO2BTaAWfUi8QRgMPGTQm4Nej6JnnoEEAmuvq3M42ijxxR
MXiRCqDoUWvkGx8nwwGHHUYgtVRJzvwoZJURtpNV78NSqwXyQLX70Y84w7apfTbP
P19lTKTeOKZZxPph74j0dYVW9v7o77Jp/4dXe3AeWdeux2ItVau75RqNmLCgcnqz
EdjdgP615uNkxF1njZd7H1YQN5X7gCaGWtp92ASQnpUdozC+C6Cte9izct/uJjho
u30N+i9EOMbw0zG6Si5WeXGxp2eACoJCNKmsaaOejPmDxtsJCuaJtg3jyKUNrAQQ
zaYNHyT1TXp1YPLdxcWBklegmmtZN5a0ql7svcc2LvRSQJXZpu8Ooc5/yU5Eew4w
J7VAIPXIaqbmgFb/LAJbPMeqJFzWZeRC6tVcDLpskor2nf1qW4LwIqV7qlJfG68B
Th3KP1ZgFzN1K0paxdtCaihcgZ8cf1kyufNg/n+B5z5k3yDc8KZra6PbbHV5uzIE
0wuDEdMDQpR0qtG1m7LfFoABNz6+fAEaEC07BUxyHDyh066C9geS+/1SRZPeekbW
Yex04HBOsgk/IBdG0mdFohYKqf/o8eNPU+Z7/zVyqsC3y17NuDtqaWTHTFRW/Mck
OrOUk3Z5nP1Hv+8Ba9Wwbepw9NbmisAVrhlRsMZEWV66/d8pEjLfrc9WMmfL8FNk
nF14+iKmvnxWGkcJ6aHlh+Y7PxPijlBSgGt4DRZxSSPSAgzaC3OfzeHzIIefxqcE
sD7f4pJsmUSPNiDnWuUSrA+i0o4CGynPeoQEs3YfBS61l7TlfV5+5IZtvWfeIvxU
0WEunJhH6h+AyDOuQwm1E0xu+0CAYZOVezPeyUzG9mxtB3jmhrBhQduS3ophyEXq
Hl11PVuuW+faFigjhnsDMDhbOZ3GuUlRk5fdyGlge18WaiZVbGa6vt5NyEioSAGq
6BWQcxTT+BVR9Euv1EFyzXRh6UaRrPi1KNX7DcM+AIrN7bjanQzW2HnWDOZ/pAPs
9Brm35xXRBPeYmYYdqWShmcb94T7um8hOgWaFUOLaQEpw7ESJ2pydZ36Z7jCJUhn
eQhvPnyDjulrnz+WWhhF35/iug4DY4lfb8qe4gU4B6QLnVq1i8PUNxLNDrg51BT/
pgI6iJgM4AY+HIrYpA2wmO3dGf+XMYxw7Nf5rkFc2dXPGJiXBvqTUdqqudBOaq7d
8PMUb7Cai12sEhVLWpZhfYmoq7hVKAslUE8cqjhi8YsIUjEZyRKhej8Yxpdbh+At
5B/aSbhCOaYN7JhdSTlbSyfAnvVSEdCaiHr8bep9k+Sx/2UY/Ruq3q5EZEvLR82A
XPDQib3vLcMKmVI7y5A4UC+py4fwHZ0NQqrfY+ova/9qleaLB4uJqDTX7NuL7D2y
xJvGTzxnK3mGsAtyRZQEmufhxeVLQhUHzOv1AiTgxmzIiDtCXAomq9bg4V1gNkEL
aUNYWZhSe3s2JdMYljDcs50xx8efGYfPxfnnOaLX9jqsBQJtDFHOYpGqAewRabYN
jVww62Xa42cSIBNtRGiDSz1QK6Xfy4fbt7n8XnJjBpCKmVP23fab5mQsi2Q2gAaf
TRIsA0RiN5VXs+Z15MbuHLlNB/Z5+WrnAPdaaLe7ajnDiaR9iQjNNzv3d0uir3VE
I48g2w4YZIEu9uAzT71Mq4ioF0MrAbPG4IBVKIpoN0uj5p2o55TV4ZHauXi6YfI3
bZt8ssS2UVzAzPuNCzF9DagMXkKMy0oz4hpNeSvsF66n0iIvp28RvEjFzagWAll2
1BKcxrUFtMpYmgoz9NzNA+yKWGLAWseeLP9q6mrzwy1ML6fPbzJ0VvLGGTFBR92T
JtfxAcZ2nP9lbRyIfPMTlofMvCe3X0YJQ12Y+EwxMlWCqMyMCd71tlbAhvvS6na1
0fAkAzt1OFLo706F1t0tZhij2vlsEzmGuMMMITg6KhDHTyqkoMcLtO0gd/44iVxw
AqZaL3NQz/iQvM9HMV5+hW3v8iehBf5qXSGjVk9RgoZOYicMwwmU85QQ8+8dS6Uz
VmQq2///S8vqjsEPHpLbFvsrIAPdY3nFkZXg3BudK8zXQQw5RlcEyHzvnvPPLPcH
SoweQa/d3LjX1R3A8MZgrWlY6tnwXKqc6U7FO/8HTbPpLyehiR08EGawPY9/Xuo9
1GnWVpc0VVwgKxjNYH4DVkaBSfOxMb05Mb7fh7GHZhYrtPcSqZKEiwKWwJut1Sxe
g22yqmFf3YfqivFaDOAzNhNz7Lsd5kg4V5bnd4fCYS67TQFqP6lJ3fLvp56wZ6Xx
Ch3dCvcmvTVIip1UMrxD6WFNv0tJcV83RyjWalFoZ9ozD0NwtRAP/iB6P5/1v5FG
41/uQsckgTZNsLgRydnycWDapmehU1DAQr40E5LuopH1tqAXIsrXvSMUFk6Mp97L
oo294YFqLMIhlDhTy9wJC7p+FLnHXdKeC7VcK73SUg9n5a8MNK0bLjsRrThS1joB
/IXlhVtVJILUi2LF5iuErg57tYdc+3MjmbCkXBLpgkistJc3Y4hx6+TNUTqSMh3s
KpDJZtUNXlwC9Q75oK0cRlAeXkqgEhOQDjQ7NzCdVl3d2vZzsrMABgD3ekJXWYKU
XcGvLAc9hjc0gbAPPKlazLqqV4bPeFxg56z0TrFHeKc9rGM529F+sXAPO21qj3kZ
j8zSiKFKwC4vdTfFgNZbi+q4Moxqd9lAasyRUEq1lNoiWfh3jdz5lg02F1raMFR3
30/O4sq5H9HyyGJQISlCrT8vZsolfXmGsvmUkFXbZsd1SDXyoYoIxsSpZzilM5K3
kijN+rIPRghvMO5NH87I3BYrV9W2LOrE022F1WbwkmUNuUWImFBCQKiSIsnxsYAc
W7NhH+irpxhd9TiJx8fPSDdXpBUsCNkrWSliRro0TIwLgZmIo1YDwuuEIM8XCK3a
st/Q/f6lXuE/MPAaxkee/poYi062YX/EJ6MqJRvWGS88DsKo1XBOKe0a1eXBVGLO
teZtzCLzcDtPOnjWJRzrWX72IoSyKp5/LDwyRCU8Xap4vTVIx4s8d29l0X5Odv/w
LMiPWVGTum/OTMgG4d3Jhq9BKYExMlRsu11Q7cM3BPzLA59jrAff8Af3fOFm8BMY
Y3tLbwM8iQCr5od3JvFLCJN9atEsY1HdKSC7ndwNwmeMSi5YKT7oBHVXrOHQUZOm
61NKoNK6TuXfc3GruYL/RuTMOZyCZTZrXyaCrNr2QBAiGBmWTzkSdNceTfkbtr9B
KJWyONYFjmLUx9vh9YBYXJplawM/pcQjEXteY1O5aoFaxrWwznBHQHfy+PhSO29Q
pT3M7wZ9D0xRdN+1bnJ8U6AGYybJmDAYIOjIRS2je3MEYzgU+rqSpLVqXnhZ+1ry
LPLYSSEH0jEfkyaGVGMOUPGRSOsBnrxHbqjAq6NxQHY5O6J+4/CPLf1SMbgTgaKL
vtVmqf5NHK1wxwqewk8/2IOSOPEV2Po7mgDobsig4B2rtPfPGhpQA8Pw7CXfBi+3
QVZVY2Asu1eAMSALrU7eViKXAqaGieyZ8EzkEAHzCK0nSpsE3IrX8YRLrsydvnN0
pLzdDBhLUqzVZnrmIr8jSiey6fLFtm5evcqH8O3wbnn0FM07wiROivwqrA6gLHvV
hWf3vprDKDYzoxMshDcnuDrKj3EWBXC3CqKWxjeDsdcwWdIRQ9PNS6gGm3+71FwA
jxw0db6OMM5NsfFCbemzDhjNbTv8RPPFTrJjUEZns6UutlEUam+m45uemNzwdCdW
cQCwksEydOsbzNnRv1YKqCzMklpoiUx4BFtvTauPiPt4NFxjnYtAL1Co5kcVRfd/
7GPmykOlv2BU99aMyHx4Uvg74FxJuEWPjAku7R0Dj7HWbgNNhLHzCMGHEEcnbQTr
B0SeZ6xdM/BdYfs3OMngvFYBsVuhAZ/PhKhI1KkANC4Nf+DywsNx+QZmdxb0AQrn
L85qNuj/R0JHksB2ZgWDjZ2ioc7akvN7gPRq79Cw6Q6tTTDB36gBLyFEI7cw++1v
EINBcQil065TeVP623TsIIQaTULemFhyuoW2WBkw5nZqFpd2dwvraEFfhW4tuz99
psgDZdwSuNFj9dyvw05uo34fS/XGmbs15d2hLV0bOfarqwm0Ht6nKBAaa6A0/6RI
4xaR5IGmOu7VGg0iNoJxA6DctZbvPBsXhgrCwCR4AFniHRIO5lbUD5eh/9y/H3t4
Bov9L+m/krs+O7JyF7yOIMPNQtQcwRHbU8hZX6rwSuRFTJUsz+SQbsvzcFWbIBsd
WnKnXaAERVpc+XuSG2xtHdoFvMghdl4hs8K1Vy2YIXroCkXbPLDGCnn2+L/mYz7s
bFbERxShSm4RjGsweuY8V14Z/Od5E7p1F42c5cLfR99e3kOFOVVBNGummxsc2ciJ
ZTBLnTEx2llpGKFZFKdHrKSq0h3rSwTVyTkxzwyWuWV5jbsrp4pCttGOqXOHbVSq
i3gBMnGCDscli5p77NNAag46vrQ3qPv7rt4DH93NUI6qFKCeeA0kkDdchgIdV4fY
RraxiZ+sgIYagDaRb7NAlA5gnyR/dksirraR07zdrzQKdAk3vQNYFZAt+1Gu5buh
SCtL8eqw272djajEhTwUQUp+wmtbG0OuCQup8RzKqpY5SgmlGj0nqPUVWAF1aOaw
PS5Q3eStLDjsPPtsQ8eeh0MqtIz5fvOvR6DIYpPlyQxuPFZrTV/raK5oElJaihlE
h9JaV2LDXddKfCvO8xrujE9+svl7WFNxekeIbiqKdZ5DE1OA6AvuIS3EN4raNSNZ
RjWNdPpWDLzlxMvEOjbErqfEa8JrgI+Lk0F/Sky6o/xcobPCoXuY8pG3dfZTDbYM
bnmtnV8xTxaokG1uEy6J0B4kX1PLPeIFS5lzdfGUIRRCVDXIENKwpECzHiwIeAwp
zIdhwsaxkHQVvis7BBVKKxTLYBgtBgSbF4JJkVrfpUAXeCL3ARj51uYNOqCCFcN9
nt/SmS5ZD3BTrm5iscFQmbipBozvejb2jO8i0XV+bReWHqETTvyOf9JGAtUr+CM2
vNwpN0ygHqE0cZPc9IbybvF+HsdGs1Dav5uUjm8NKbA3nrdzLFHgfkxN8I78RrUN
G6k3YqfReBslgpVQUCzYvPLbpRAOn10yKKhxEdO7WrpTLhjeBmOkzNWYCKOgLcaE
0rUPO380jwX+ziRcnhN44tMKr+aDXPQ/Vxpu8niRYIP/jhhb3zgpp5SQn95o0dvH
KvZ1mz0OKpE0gBkBiK4QD1u2GTM8HTRosuCcT3jTplX7E/TB0ZkdXKZhK0UsL7QT
ankDqdeu2SDqsOoaPtfgN5FEolICvmUKkD5o8lZQkA464GWtdE3anIOlsk6MUCAm
iJbv0tASlpk8bHgXG7pZNVbOBSEhmg1h0zpskbZgDMIUDYgAIlPg0loEI6gRSktd
8VpjPX5LWR6DvE3F08V9Ucen0okoraVAif6H5z5sBBOVKvB4Udm3HeySH3kv5olf
6Alf8zXiy1ftWnFiTlgMHCv+tBcsmKTMyMk+RUsskx7QWh6DHDMsDUtYk8lPA+nZ
juD6e1OR2i3R9jPhmH8OnToyMY5N6Nlhc/1bl6+R1uJZ+k1dpz/psZ2BbIK6MEJ5
SuV9/EsOkxKEw1D1KdCpQ83C07qubC9ii+L1aK8rUjTqFbU/0bk2Sgc6RKX08IfA
4Bo2KTUIaEMhsjwL5mK83JmX+Unwz466erbSHImZ9WJLgBbKClhcAeMsYNtUwz8M
bi7u1Hv28qQWQ+NrzgrA0TeDFvtsdnDmeJwVDIOU/ASnp1+ctT3icZEAew/Y69Ep
BaS3mADyQGXgkgwopJLH7WfCFwyMiO8o4xdRgAeHtflczbKqGMCLJ97wiHNlVlPI
Jz6ifIpDP+WQ8HAyeCN0vEsKpYbfJqDw6IxPip3YiysPYoLbhBW1PxaZCjbvJXrT
fAH92iRBRSE3tnDFB0sstGadXzqXzjqrbpYFUrpo47/dp3m24mnP3St9EWSIevjr
Q+hjF68ial/Qk8nga5PwNMHGEWiLmFR02oFbXMN25dGtZUVvavDMquHxVVbf4H+K
dtq85SKqYhPULZ142UOJJVRig76JxQBcpWo3s3oz7Y+eBtoKAVwfCym5UEqWrjQY
VLd7nIBjqjncsEXJmDGvgyzE8Dl7YEsx/TYIKlYHzyORiZoi9QtLQ/FTl+WY5zGp
GMIiStP/lnLYx/D75cCTHqXM8N1TMb0XwqSbIcG87zGrfuJU76t6ciq7+to+0tIm
4ZBlK9G89fqW9LUcL5QJpuZzE8/maTle4hc3ZS1q8FWJmGbivmmcHS9/mAGqFFCG
tQIiSJcQWcFtzZfMk36F9Ef4e05VJ1WQd6F/9aqlqWKL6I7qgaHau/GvH3VT3mWX
fKqsz8ZY2Gcj0mdct0ThJ2S37eFqHhEAZyejBCOLeU685esvXnfw8FtEShxkL61O
SynPecbO70Nyrkdsgi/53sEFZaZukPU2gZFsbs7fjpW/ua+3SNZNk69Ze1jRgzfU
jd/m9+INQUm8sQRAmvYl1jWqtdIrb7atrm+zuWEkEKWiqhgcBflL1gpJa7F3VofV
E1bNOFX1BWP9ngewQjihkBy2179uU6klcyT9lXLsS4R40oW6jcC45NILUXqtH1cs
QYLjazCW6GuMMNd/7INelNgY5BiwCIkbgiRyERHS+BzeKI8cPFy/YbeT4mMFcPfL
b+sDZp8aM0nFpZ5ulB71xKqo4bVBfSa+IUq9jJyMKgrH2k3ppCflf5KB/o8ClDU4
Clt6RgjViP3nUgJmaKhKL/Zo4tJPCorYd4cez5DTyWJLPTVxQ7ejCLV5jObPzMKL
hI+VtTfQODg3Uf9eecjsyVxZuCSohshtb1AFJQTUNiYrTF8liRSbcxAzQTLejzjK
Ihy8pYAxLM3Q+QuM6e5TF+/nyNHdvR4Ky26PEsBW4IGAscJJfmUBK+0g85MeoZTI
dQbxmPR0FYiF0CnpY0inG6KXiD/dLYVB0AXnG/8mhn1f3FZdG6lHx97nNIaJqZg3
KA9jAHwsM+BZexl32KubcU3GKML0g68zTZwEMJoUodZwn3g59gqh0IEMPil5iYYm
c2UrFCUdj67EWPNdqRUAX0xqF1QF72I4ouaCwOwRS3WhftjUsAkWugLOsrQVjbYm
15fbpRZSD+l4V0KgDqWKYiaqxGIfsaHpEGW9BJVofzqPdCIh63fk1l3EWmuIGAMc
u4GCOwGc5FPTd5HPcYBTbvz9gNqxzwbjPr/HbWxfXGFfGDUD27IihC5aEzy64m3p
+gCebjqeRzf763PHPYR/CndjIU2nWHF1ZoAS3M31ikIHwJtk1uIN6wL5HYaMpZAr
vcRPMOKYIta4rucGVfS6NUhqYtYRb2A1kASl/SXuneQfj4sB9arwBJVnjV4MBnBr
lX6H5EjRC5GVNamAFNmE9NdMDk/f8lFwXjjZe0bexA/Uww8qfJDxJrYjrH8g2cQo
4E3ME9nj37FKmM/UQThZ+43LtorKTLHfroIZ/7WDqGFnP2PqWHdOyFNbtTKxuLG1
jtQsdRKVfQcEZK/mhuuOCLog7NLiug8A5VtZVc76xol11ubSr17XfE5xPoxIdo5e
SAxIl3QYSImm0AEbRul6yD/sECc3Cx4iJTCAGgH6UyVg3IOm6rM3AXxL3s31mcbc
24wzjFmp61qQ9OoeSd56aj/NIRr0lWDGMYqywmURoAdtz2UUSLe3WAzRgG/cHmFf
cIqwCT2RaIOBThCQ3Nx5FhItZsx6T9mYCldlAqLBw1P/4QUvKdgYCYSa03Z0lTxI
1sKtf9sNpwZvza7uYNXg7QgJGrVff53/tBuF8JMaD/l7uaF5UOtFzpy8hsAgXOF7
4bExxvJTTNSKc6/kuIWnk/w01yuDKO8U/MVXhe8aP0RpaHcHIKoAxpzPglz7Td4P
qf3G/hHDP/rPxD8hPcpfqwhBj5RAujq3qr/jFncfuuA+7si+II1TEXk4hYoqG7mH
ebmEh7vmf8DQxaWUlCW+5lOs2M7LpXpG6Mv4j/nFD2XmVd+LGhASjLyzZXKyAtTn
KbH0IsY2qa+dmm/BYi7z7EUKet81XvDj5rsRAToPEw4nNITRzfpbaLwjMzW5Xkqm
zvDUm0FU0n1rLCuqjbVN3s9MFdunC/N5GMIY8kM7KdLIgnfZFZgPL+Ya/GrwEcLy
C2vyO+FzJh3jIjjs6T8zH+5vJDqUAzzGrweaS1xGTF97TOhXvuPS9fzR9Vf0rSyV
7tpTqWPiFuLQflJeaZ6FZwGWcy+7IxL/397YVklc0Azqf0zrxDnJknBn76Ky+VXL
XeWs/Oib4ordz2z7zE3QbWhN4Jj2ILC6ZXiOvg5Fk2O8/jqUTRAMHyoldcS2Z2K+
ZLOs0vmgJ3lWm5PO+Dr/jtgcfPX1olWK5KsIe5+ExQFxiMGFp8o3rhm7Qon83bpi
X7d3j48lAuCODdcg8AbMqzuJEJnsDqSa9gQ9jY5xFvjMZEXGkIjFlgqFxb0v2B3t
a7OxNC/TBKd1INkME4gRobK7zpSrAG6nXcPzPMDF4avvnsLJ7RXPKb8XnK+/QMQ4
FVRkBZOb83yFZLEtk1tjaWBjvvtna1biUsLnWKv5ve9v7Az+BwgZrkzZSgKlI5Q4
2L2hJhasrAaqWxlLRSwnGKjBbbxC/yLqq3DuYly28Beo2/KEkCPshDUsXWmx+wrt
LpnmV1JaYROl95YqNFYHMMa9D7Ak6U2YsyL0XC2Fmb+JRvxZlAxxQQEaxfY0ymzb
QE1FfALLybDPtU8EygFlv9DwCaKKRQTdyuurCSpL9eNA/mgzXUNRglyxX6iZeRAa
CETcDebCADGgl7c5ktbvlcYRD/N0fEkUVRIOfBh9+mc9os5lHsFRAuZyS1mOcdYD
KuNzxlsoT/5VgYOeRbgTl82eJXd8gY6wKqBQ8jUOayELmfhJK5aoZDi1UL/W2S0u
fiBmZe5CNZq2kHqvWnyXuOBEdtdzMfP5ewThyO1BmHdN0esqGmk5CupFyGW0LNXi
Vcb7zsIXNzaEE5aaEemxd9mSbDQUi1xKTNSqYa6h7qB5KoYkdT8jUTlijjC80J5n
S8dLWGqWpHGtOsZKSyx93098K2t67mOTPe2FB6p35UpJmTi8QBsvxAyc64IjJeZZ
56x+wkySou8gjmpDTSckNb2xHQ0CirQwTcqXJB8itYGgOvlRaaHQ8iMQotB1BQuv
x5EzPmb14PRQMXDKLnbe/3X995I5kLvadw/zLG7gYredno8CWT0odLNWrdPEj8/d
FxeYcFEeNwe79kGsVwvZAFpJluAPj1m7lqe627L+2BmPnrDH93cb0WJYU6IHsmTl
4yPS15uodSIiTXm1jJQkTWyGK/74jyB1hADMusfAh5HAuErLyn+S2MbGBXbHHhF3
ExpnLX4/gmKPgqsjK88GtjPGrRV7Al9rjZ23wJwtXC9mq4eHAtp1RF3rGKT1nJqp
nqKwp9wZ29ep/n4HQXo2X/bVV8AdRDt8pnAkItAlcGMHiin/UkRmGE4BAjPL0mwm
fJqyRUr3B6orYQjf4aVTjvn9eQB8wzto0MSUM2w/yblZalTSGNhkpFZOiDBvtKux
0VGlpF7bBlz4nonDwAnywYcqJZACOKi5tSmoBfytGm8z/B23oybpM9W23p+Xnz12
2Gvl35pkXKSJeO7PWAnfQAZsgCBf7IQ8TYvmonZUSTCWjSvDGyxLZBhNicWpq63E
LLRJUcrYX+rTtVA0Q3Z76CDcT6Eb0aeogCOmUYVbWQcGyeQrqSFWaqNUxxlrqyWc
Dj7KGX1YINeF8hpsSSWqwowqV2sC9TYNod/TfgXYOynXL4dzaDY8mM3PKDRW0zg4
HHjNG7pAiJK4GHa2YlFBdBCYUvKzDfOLqhbfNC+dwlEZKpum9Cx+W61rSSNC/aKZ
JbJmgn8jTGRHkgwMu3olnMPqVMBMO+F9hb6fAoX7cHNXhJ6CfCTg7vdBArYGZVP+
OeNlUkRgYEGdI9W7CW9uEHkOwignrlKyKDOA41mgXn4K5KQYXf3AjGNwJO6JKoFi
hMLEVtVLg5a5BainbZvHSbCOS/dvyAOfIzTqboKO2kYaL61v6RxyNchlOmDC+fL/
Y3RKF2ETahwou6uZep9fTkQwEfOBWlT5pgkoFvu5TUZE7eNeqTGrc7RdpqD8uZc4
ZikhmQqPqrB0Sn0WdbdykGkJmuw/Iqk9/14+dPFK+IPRkYTcX63ZH76ZcQaJlzNq
jmdx3VgLACGC+1O9JciUQLf17ziFNbultyUCU/NgWNprA2XPlej9mSJ/MT+7yxwU
ZYLlSvhacQvLAAQs8tQwcE8NbpyCr4t92CYbJu61aL9k3aCq4oRauAYpo3SLZfvd
mHpkkG9PZwumyh1eb2hiznFBh/jLSmrgEeqRnyEsX6jxmBZv8qrjzkL/QAwgzmfO
d2e67wDmfmEafMIprTZXiegcnGbwqv5dlq7owAdvPeCs2eeSdDeGacz0eHjOgb0s
+5FEuwRgeP2erQzibTyqSGbG1hkZcQOxVHNtCfLAXjYxyBNW/dZGZv7eDmpw3UBc
pPFt1GwyOoJT/sOJZKxgeHjAdk4zEwjPjWXVSk0SkFTzaNzcElXlAtiWR9ZgiMvo
AMwnrMKc+i7EYDXJC6k7qF8+EB8vSDHy2N6vA2e7H7dqZhmI8uvqxyjJ7ki1kUkl
/XqX1hLJ/2/Gvm4YUqpAQ7HQTKfCqgljNScT/6gH1za7f3CbiPSBzSAZm7p4M8SD
4sR5Y3tpWbpdYvGWbCcHbUwBsObx6fwvZOu2cDd7cQSfvid+LiNky05r9AXe3jik
KVby1SevW10tXby8AXWKKACbOpXitREFBS1eEzfmSNH+mukS45Ny7bFoClkxzFa+
NnmfIWYrD14rkMfpyGUzpycj2YWgTvXNm7pNdvRa3Pn0+pCoY1ySM+rLYEI0mn07
vD5Ja7FllPgcEVarip8j6MgRuvceUOJ0xnOIdldVO/ljC/uwglurStZscfa5qhRK
Wuk+/909tKTidMFxg7A5IurjimZoybSbL2C63VD/zV8zSbWzFPCJU0Ul7rAoFu4Z
EeWXxlvsBPh228NxldPzFC+AjVI1EcCDjw8nLPy/+5ollanX9qQaN0Fgjf0N4423
Jdj1AoGjZLcdkFz3GJZFSLMX1JSME4ltVg7P/0Pcz4CFmEKzfSP1AwUm5SU06EoX
Qc+fjqZbWa7dlKxSX83NTjK2E3qy7u3tq2sO+TINk4vsr1zBB6uun2QI0kMuJRc7
NBH1qgAoZzHLkvhPqGptuQHVXIQO8kI28Y13KSocw7nTtga8ryV1/cPO6zdzRWce
ZAMyHC4mgtnQjByaTOYCGIUaBVBgVKShjpFHFVGOEBmLxCJUKJbozGhcVjGM94qi
fZJLhKTneKBJ929qIuNxpHCQ4mtP4l8QXPyKMfss5oQ7xKYY3vCvRbvGy44SktPt
+ouER0GfnMkgguy+Z4CblB/1Q0/dNRx/rP4RBbBYyWIpPfogQHJSNIXsv0JG/hAC
XD8HmGMZtONOLGA/2YrlAxLjk3FHprK0xlK/chaYSiE8Qx6dN3y+w/mevgk1UyvQ
7AURbjvxa0IBira3FKKW3S/on8oRpXnzam7QgYEYG/dbJcTtKGaV18+wkLOb0gYh
n1Vt1ixtEk0e8QFPy9FfQSCqFm9GQhn2ezNWZUiGahCaeftOk4N4J6FVfok/RLXT
poDCSEUwcv5keFnRnZJ6eAazCUYhRCxLLgbbfdlsZjW+E1YG9roeNDEQyUzX3bhC
SqOA+xwyG2l8Z6dlyCKK4Ejqer/ecMeOh91QlDCj3GQozQ0umHcZYgY2SVFEiYaL
9ApowER93cSu8h7egWSzwxlDUYsqBM0gtCv8r6E7nJIOP6Mp39X/EblObAjARGzG
G1BQKGiVZ+pR7SQQl1OVORYSLObmcZeHMRdgDf7Dp0kD53e8L9i01XmjjRTRjvkt
yxF9AFuVvEi4ri0u3Mh1mGNUX4G4FLPww3gOjn+vucg/GwGxJgE+L4BPJgpYQQIa
A6/1cHozTy+JvYPUYNgkuqI/2DcO230RwTI30pqz/M1Mr/I02dHvLbO92fZ7cix2
fble9koX0xlyYuc9M541E+/QNRh8qBPWPV9G5khSSJ7P/t4faeNmK2B1ScWrfPen
MbrhqrVjKFoQFuykRk7MFRx/Vnm2PKP6sDNIaBu9s2JY/2Dfcvki8yrjSM5cPTxY
UY22yOvQe5NxsUgf9decZdsmcpDGbzEfNoR6L9esWsCo7bHx/+RU9gWVT1lkALIY
BrDnf4gvjM5deP/5+wSiMlZaGVHpcQGiIfAYBM5Fwz9HSnhP4EdBZUmU1B1d/OTP
rYagdj39S0kLDFpLcAndIMlyPOnQXPsMd1f5iRqnKi+6oCXpOdEHCVAXFWQ9qaSn
gLgpAlFqwJ7lonsQ1cDKLxlPKHZeVxj7lg+sjk3GoDEZoL5zBqJ775OQU4OGVsr1
KsX4VNpnH7MbBmSm6i3L6FidCBtCpw19/6e4nFGNmXHbqgc0Ei0Z4Bnmy9jMPCFB
M8chZ3/Lc0sZ/z6+fevq5HF/FuuiUGBoAwE7pZcm6vhHIlSZI9BbxPsaqnKhjErF
B2mb78SYZbRpI/SOBRNuv2VH34ZjAAOwztxX3JRiHS3+74vvLwDu0eCfV3Tuei3C
K7DUDwHPTvfe6Dw9u1yGVizLRXz45kPIQkH2Wm4mb9SXb5GTxkvRQ7x9m6kTUESC
d3wFakPGS/E6GyWBSwGVIDk1jYEWAsDve/jswoSWJPWA7CLmiKaOsxGjoCeW6ici
rR9O7Ktd6Itp+8DKb0Pk5zLecBWYhCYTPJfSxt4LGkcNMJlljgVZFrQFfdmrvSJ2
E70CZO32DtrwCKy8gX08khPxBvLWZZXYpr6OaBZJpL53b0tIN/wAGRtLGlbbYVo1
oxnIUX2DtCIm7AgtZPbUXeJxwHrhA87gasFF+rODs59TSgs9UUzSXQH8zED/x/Yl
CDFl7h4HcJMarzslIWqDysgfODoRGAXJ+972gDz9NuBdkwKh8s5kCpxoORmb1s+8
7sCCl72NXOL/v1pSB/oZfQtwwISGjdYRGNGcbteDof6dIsLg18Zrrt6i41/9yr3Z
SK+gi8M8EctF5quZw0bKE4fGgf6fNNfpjWZ58Ows6Uj5+89AcI5rxGX3LYmkVww2
J9VuAzROcC5M7d6DV20aWy9PWJQU7leuMlJxLDCIBp/S/Ew08NMHb628R1Otc3bQ
s0PMlL3UpTA9wu0ZUlmrUvCvKOO3b8ymx2OUQygo/ziiTxAfXDaX/UuNHDyyJJO0
T23LmvchqoNCe/0TP6295zhPPMBos0IGubfQm2HBmw+O9JG42WhElTTtgGn+4+Xv
O8sZYulsBwqdJcKB2hUEiPrERdzIspTiR5ITFUe1HfU2cSywiGSmaBvHh6TbR7fa
M9WNZGobMd4cQN4wtC8ujypV7KHUhrlscpbzygf9xasVydSf/uRIlsAJhUd2xhyh
5gF22PNa28o2LoAH/p45mWmN7PmglKjKeYJGiEz3UckPBSq2UY96Id4KxU6eacKd
uVmtErCOl3dqo+Fd36KdrZsQg1lNdMjKQ38CvdFBQvR3/h6XfharKVsLUWabAXQn
X2q8XmXOhl3LYDEBFtg3TEkikZVG+2DaQoae2f2HjvCKKpzGKUSzdhOeV98/lZ2i
HEC4/6hVb66fdWIhsV1RbCxmN8qh+fvBTi68p+TtGCCsJIPtMVpMhaae+LF/J/8S
D6skpCART8sEjKo4UhzG9WEybCKmtCsp6gaFu/mRtRVT9ntOWtERzbRnefscvM+Q
r0DfOg5fru0YSFtflzYYRj+98N1LOqRF+mL/8Purr3/34Vsz/Vf0a4Oo+hiV3DLM
QsJjra6eUNqIhJvpGCmLFCxBQO6KTPL7KX8BEGCJ4Rc2mz/UNXcYa27WkSNztz1k
aXxxXf/1QJ8KWF9ny9UtMhwRotogJ8SWpWLCCy4asGzCWeabKzuGDBpKIqqxp3hY
H8rawwSJBpOuVYGyABozj1PQv9V607culFuXYpe+NHp4fesD3FYHDOuGWnav0m/e
8NPGkrYBqleobDqbPZCyVQNXxRGVOcontWJVmderzzYxrWhBd7OPF1/lqyaz3kLn
kHNtFiyTxP3erXviFt/St1ci9xcxkJeSEoZuHQiabPFQX5+HnxB2ZAIqCEN9inul
BQhTGBQ09+W6j84E+OMfPz0grXTb0AKbL5RjkdUvVQ/f9VUMb0+lTyUlc8arohfQ
U+et4czW66EX3K8h4G/ZRLtNgbxAhCPjQdahHeb1mYfHoc4dz0sDIdHl4Dh4mmzY
33q9KmVfkVVBuS2fbZmDS6kCnE0C3S56yoA7Fu/c+Y0Dqyg89JQ/nwirS8/+i2z8
eX7uAp9FSXzGe3rNB8M20/7EX17WT7tvrXRwIQvlYrvMyrJe4tDL/+1ez56MOapx
fraXm476kBIdbpDc3srdLPagA7BsBWLMeyIJJAzNP1RifszWhGlV/v+AFK6Jq25/
UQG6EoTwPtg2iCF0PzcOLjnRRd6BhfnGDozvO+05xpzzJeLPG5tP3ClLiYuP56qU
zaKJI22TSAnU5hc+ofEUP6BRN6euCf2OVlv8nnwtVfkJtX0FEN/StJPuL9jXQC8H
aqDrHhoZth5tFXDgT/909Vx6ofXdldZkhw6wdEx9Iibr6yy1tMojg6/irtf6NFkf
lkYIYoFrlfaeXaAt6Bn2fCipxChoOAcohoWC1B4Lo/db3d1juT/2XSO+JHg9/dBR
D0JWjo7DC/LQ+NMrsvizFsftbVD0NTFfHQglo9BMBuH0EXvJ2j7GEu1YFEgIpWk3
FDnRioBmMd4yB6d4lXfQ3w==
`pragma protect end_protected
