// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VbrTjcbHapGhMGkPFx5aVVq2kt6Hp7Z2HG/OdViNHhNbIVl9IZskgbIm19QjK6Ez
ij2Zi+sjMYsbNZNCTwRkC+DA+/ihxMJe9ASoNOjVLCGYLInGFttci33TA9kqOo6D
yHEMUbxzwes09XMUXJaYUMu8Wl8cxRSSCBbM0pY1Kog=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20816)
C3NxLt8G43CKvaCim5/G0cybgHQblFKcofEnc3mvoYOnzW5YF9uICV8+RqdqOGbW
nvtOmkMjlnj/sADsrCsuQK5U2VfJvhQoQ3Hg42vyDv0Z3vwpX0ZVKjymsZLLmG60
1+HSamV7YiRVoP1ZQ8ILYrhi8qwMJlqP9sREFEguxn2OIS7OCq756jcmIM/SCqTi
9lABUDz/cZCdsxWLNzMW7xknaCeU5tA31Y6XNY6rbOF6QzANYo7BgFt+ZmNNw+qY
RP07nOk5Kj8YrYeZOONeHNHDoRHeCGKYzaRYH+xJ6UOpJT9DEOADZCXqLtKEVMzB
x0+CHn2tG5a7VcgVjWUbJ0JFhj1bIk+8uM33eqd3THJOIBE8lDTkgoR9Tgs7AoXu
PShJ9fIzIn+ZGBHW5c+AVZ5I3yHdo5cJRd9ruJnKSj6OXdRODfvBh+VgoQw09bZe
UhUpTyyaWUk/OovFXuInPhdY4TbkydQa9lo8rV5Lx9oJY9wEjfl1Uyig5Isd3rNb
YVCuzMrbIoYQ2Gx+EJv/mTFwF6Srq77/PJyZHQeE6lWp+eRPuqysALBDeip4ATuT
4aw0fk8/sppM9f+PNG3TG2BC3NAahlJGg6cBDhBROFNzBcYWxPZ7PHVUshgCQdPw
beI4jd5yDRTbv8hz5gGSB2mlJ0Tr7h4k7BcwtCHSzr10rKyS52S/Exo4IoF0bJ0L
npglBuRtJfCd6iUlknWXAvIli3n0w2HFckEui1oBtlctIzvTz4HQQJz8qfmaRD7f
c946UvOnbhvs1MhV2P2Ds9QO5n5bMoSQ+K4nZ0IrVFLfzc+hSzER75lCTyZAILtn
gFT8UIj133ioGzr7O8cv+OaTT4ABYK3pSofpVgcxF+aZ91dH2bD93xSy3znbkEAM
Jbrkzoo3apXGebxA3kp/IA/7pw07LBZcfFSkJ0GaI2z42kvcpyWUktG/tOxMerdY
kh+vVk69Rb/1AjmPOQHvIFMlGHodX6+IKZGRLyIlko3vdNi67SCx1w9MNWUrLhgM
gG6FFyMFGYWHtFL+ghSt09DnXhYoDBZcp7dlkKWG2+Hfc6sBd0SZnMayaXbVGTPD
F7+PFGqHlobWzAUW3EzL8927lJ3Cme85UWnGcTG4W645zfVF6XxH2skZvQVUv/rF
dMOCyuMNQ/ShqpUZrqBN5NB/LQI9C1Z62uwvd4brGB0qghRs36Avx+GtQazfkCRQ
bIERMtmNTE+2vZ+5FB+TVnA5AKhipc5/w6nFmI7dWnyioYP5LrDlxLwXsIq4wEWS
+3rlMo4g/LrHRFXzwglWPWcrNKAYU+hhwoZHmMW64WlpgPP2sewKu6y5Q3v+oRUN
BDjXoSf8WMvfJz2tXkK5Ve44/MnQ1v5Pu2QeE9WfZFisY2RrMK6uZAXkzfEE8720
fh6nPSJLsK8g4qWOA35DQg/5ZnM/oCH/pwxEfrGR/U1feRPuI1VBuIKfSfBbsaL2
WxKvJlIDOvC1WdlDKye5JQHRWGKfyee0yIZ/AzZEqNASvyXPnLZ/72k433EmpC6E
DBmijrDqdryWmr1nJR8iJKWuAZXO6ECRyNNXh0a3hqiv+b/ObNRn2+DSLVJy2zkR
hKFCq+sAHeUm1OdRJ08FaXW4tsi6oCmI+lv80s+9pbHGj4rNB86pSGG0Jfp7WJfF
Yov0NJB6iBpsLvg2tr5LGl8Mxapv/t0axZEB1a9BH50UFw+9Kv64Ja9ygCRTG9ZU
mbai7QfRDQhSux/QGuyDhF9pTw6VKLY2cjY8DmsGy5EdKBmcMfHf6hnNrKxYUhim
d0jIpOVELLkUdVvthu3a3CLtotDHz1pye0h8Cq0vx1sB2kPc7dOo5g0yhyb5k5Xq
CKgeKT9mqyHpLNIs8PhhtrIhTmZfR7M6tBjvI0kuPEwIHGkdnnMp4s5vyUzB070J
84V0KcKPpQD/k2vlBCBr/EFg3x4JpdgY/JFCkqXrco/l1AzYRztSUlXVyoom2HK4
ORST0jc/74T2VPmCmP7UQAO/3MGTh7YAq6JRLAvW/xPVJAW4Q2lKTnPO/TTEVZFV
PR6MjH6FYwTlUX85T6B8QWRg8clnb8bEKfZR5FwEIa20Vp+TrV8it0NbIocB2iQ3
ys+GwjJ8hUmgJmHV+OKi2bgt6yighxbZjh/tC7Y1Vwmdgv1moH8m4DinxO9Q1HqF
x+3fNNsfmRBnHIo92eckUacSKiDhPV6jFfinrX/aB/muHdBaZK+NskQv0pWL7gUK
OX0Vy0iXUpC6Uut6GiorChy/WojrWPf6fnFvhyNfJ/GT4+2zWFnzk9BwZ5DfB6FB
i8SHOP+8LrHGYQnIPk4YOQ4/cyuopiDNU6Tq4jXvYltzkbEfWSYBPyWplLt4awSf
6YRdbO/bQJog1c/MSBxV3RXSfLu4kSWHaE/7UiBzlLvR2YeqI0qAT21I2eAVl2Eq
gSF1lb+3gCPeB0vHzk0FT6y9wsKFkBWo8c8PAZE1j+z5Y2grndMut5h11ufKGbJN
pGkQI/u9dMRn/33vxMnbpMFvbMEqMiTV1SUh23UCW7R4+R2XCvfLltHBMdOCkzya
YmPedc9VpG43ncWBCH2pJkRWB+WtH9sdDO8+t4SxUD30vZeaA7std8HwWlyxG2Ri
oJhLAvv+B1H50A4eoBWCxgrg/JIGulbdPl5Lz38Oj3NCPp0Hd5UumqZu7rnP1hy+
kkJJbEL/ed6bv2e5hFqUuTs7PRqq6aH5mL3Ej6rQa33Z6UK3PFzfmvrbtgr8ddu6
8t2Y36pGOMnYpu/mPOzyKqJzEUbwmyuZeFh9yb1wU64vnhc+339rz6aExJE5ffUz
5vKWwtfcfyTMgb7fy+egA7fAn+HFCzTKa2OFx8/uNg6nDmdoBfNhuj82YUkdewW1
7NuFBeh+Eo4gdsTgU60OWdetwduG+Qk3u6s1FENNcW6zCgZKLL09ruKDzIoIJ3DP
tBIrq9txa2hlBX4X0vKcjaU/pFIHRDasozLAbUAchxTQYH/Bevex9JS37EheaA9e
K7guUpl/JCgrxXoHmVkMHpdl6r6aBGW1EMtNuCkNtoeW9xAPz1npZj6yZ7HuMETx
tLtFmbLQGxm7SgM9FRI/OrZXX1KJLMhP+Clftp5okRUPTt0iVNZBHJEkiZahk9kj
4qifMjpTQpl6ZN42qpnQ6LnPdhAve6Ug07vh5WkItPEm+w8BejcBFLrgK/3uCLWP
mzM2dJQ7G+TSGpmt9uVEzu+AiTEtBM/tzXxhkekCx3P/MI8VvMnEwo8QBjyAX7cg
666dmGnfeAlSFFHJTq7kzUx2WvEeTHYFn4yDPZeTCP6rKe+dx3juTgSlNflf8IxG
h0f5U3dBNiFrgJSI81GFoJmTtzofb6PO5iNLo2BNDixQluSO/zxin9ML77F5Mnne
K8QwkzfXwEVQoC7Kx+DhGpHHgF3S26AUBkh2qpDgcAvH2GJ/je2SM5etg38ByMWD
XFklL2Ec+9w0/ziQrCzNCelmgFXqqAkXvbW8RpO4FHMNi7LDGLkOwfgbUJ86r4Q1
E+Zt3vXhgSUis8RIk74I7LQnX2E28T+Q4SCVsfJ4qu8D9vxoccLR3vyfy/fzNWjO
KJRAfYgFKymdVFpfit3q1cZNj37Cb3APvAd+vvBHtdANfQvFMdOITty+UBGLYLnG
G3nXzJGoqE9YYahqnwmbP8OxBYMBNGUThcyfaCu1IVOksYKbkgs0CzFZ8NN/o+wG
9LUbRXI2/Y+TvUK+EHjDNb/4H86PXSPSc2iGjhIAKTdgAVZC2ideJ8uYKrg1qjaJ
26w3ug+U/7TfqtrdqLpGRXOqDknUFv5S2laEDK/KkwrKKIae++ouIsO/R8QVLVi4
OR/xvywF8cAEY81Qr8gTfvkFWCZ0JhJGWxoThut2LHqACStUFiIGE2IIOHUY+veT
NcYmtbZDULx1B4+y1AYUfmHffvjEbVPSEveY+WxlQ2a210RoOCWP/NhtrCTW0Vhv
6nk6vFSVvdbSlH5jnufJ8cy4yS02ddsf8ghy1MdeYaGLoDsWXQW2I6LTNd+PyNDP
z+iWUjcknMQS5O5hlso+Nl4Gdgr7SaRChEvdrwN7Gs/wCGW3I/mV7aWCAx1qsH+U
fvsqDN/30gv1dbXXMshXGSNz0Ur9z6SFQ+QkcJzuclFge95/y/HvJqNsqSa3vZ1w
y6ifqnCTA2N4Qi95NoTu/KlngzHIvKpQWtm/A/RWdLg5TMRbfwb22K4pDpw+8QV5
XfIUllzh6NE9J2gcZg3lTDLgsr5uY0oGnZobhVfwMFbWQIN4dzRS94JgPO+gSCNt
w2CPGVIlsy/9JVVVmkPO1rYUAK9rICsK3Ghr/fKMXzRvwZgw3HEl8Eu1OqFagjJv
tREq5FDwQ4Yva8X4LKu4CChOEP2UvXxolpIulBi7oYgsCogyaS3upoYZF220zAeD
hGSlZ/OsXW3GfpcShS5dzHKrP2U7+rcXfGBg0O2tZyFEzQRJ87ALhqf4acR+31NG
RcQTgagmmhxFGIQhIQljlMs12JOSKP+Vu87PEDySomAcP+oiHt4fHyq00eG6wU5H
2O8e7w7BFJyAP0YDQxLNiaLkXSmIbuatCJJP2aKfHSBPHIrm1di5yWIT2A6epP+5
f3G9FSPW8NF7nFoqbjIec59nRxwcuXe8Eq7Urnh6QrVTIer7L1sgL/muAv0L8Gap
+7jAEn7cZ/swbvAIbLeKt19U6mRItwDy2b8UM7cqFy2JGffF/7MmPK0jlCxcn9z5
qX8TCoG6rQ0D4uDyFwMIKRPGtq0TAqOb8ATeZcCCeLwBeO9kAlKK8cpNAcuqMkOO
sCtvDfwBOv5RHAm8bpu+ZJDcMJFw40XIA0ebm+s2k+0BMg35nRpMllRJQhRHr43W
RZalMEUnJ6i8BeH0/PF5kWrbdXSCJ9eEpeqX3khv3n3jvvcPaQ/iEH9IZ4VCRctw
6jlEVSRP3x1DXG1jNLlvjZ4fGlTTTIZL/Izztfq2GAH4wvwk1ajGiuQBZeoVLVx7
lJKb9CQlcb4ZrvbgjOHASw7BoNJEBJ5eAQMN2hkO6BTRtmTkXekObc6DYVuTyOFS
Ei1hTC+1w4mCmR483u2EgI7LgQ/5szkEZ64xK03wsN+GPkoOdztB+6imN1eTXhcR
gfBna2WbzQmyquqUo7nHETB8wBnCGvUmvpQeLeoRFnh7/ObO10JTHW91etJJXVx+
5p4WPN76xzI8rPmu/kJPVs6e+RFq6L4s0CdzU7cPUZDog9SwE6cc7l9qeONPuoLu
J2ChZpq3JyfhW8jLBw5ZGTkBQzrdz4GnfyBNkogPpX2+AWe6EikZ0fim3g1FvFzk
EpcAqR8dtmAj2zao41xYE2SCGUXjVKxJ9EQ03UEyNdr9JfMJuFjLOsySZCjFdm+n
YTaeyrEHI5wlSPo4ynd/83tsKTibrqC4H2f/s2esIUBbh0AK1pEcU1axcnLqcLPh
xfBOBsH+JvB5hQ3RGhxw6FHyGBIr+2cFVrxqh5JOHWWCHbv49dnrDAggzNL45err
xl/YYH8cfOFJwd4MLuVtiYT1Aqg+N/DKj2cC0rkrF8KtuFVCAwrh1qIh78ppPFse
OlaYqkjkYH258NfIAM5b+G7XhoIErZL3PHpJj74yDhkoMzvep3/WwwV1AmQdq/LW
/Grn6ZLGliGC9UIijG5i6MhHv9Q1g+6ctAyDl+QK+6x8VtUlcgB69WdMDwGQSw0b
UZMai1i2PSNDDyck4GsEZSwDAF+EKeX59aMvBr+oGxpM8URQYDyY+0dZWkC6kZbq
daAcKi+d0nhswO2RV6H393ijgR3QlOU9+ouKUqtTx8OvBxh8+3kZagKSkX2aU1sE
CLGHuBzF+dSrKuqIpgkq+3pksjH+vZhrLVkqKbNnAxtDa1t+oZP0nsw1mH7F4VDW
9MuMZDIOpwdqE7V36ZeyLenL7d8I/gu6ERsS63x7d03bo/45aWIo93pvGGyghP7P
Rb9JHNxXq2EFHW2MQQMCpyQoDQj7e69Gb675ZjecjjLeXrqsLhrND61R64ohQF4k
WmWiCkiNIkuat+kUNCUs3nIv4VDvrU/KPIYKrq4SkRZHisFf5KsYw/7tGyc0E7a/
ogtrhmPwVS3dAKOWFLTfKuG/+UcqqFs8g+tkIH0V0xAyUBSm5ne9l4B9BcEH+RnT
XrP5swv8m1fqaLhblNzR3l9IT5bzUwwdOKBTSLLpiQmr+xyqIpleorDYGVoZcY5o
Y83cLlCT1S1oM7i2PWeRuhWYJ/vya7uaTu4lIUBsuaHfz9+/aYd0i3IyXKJoR8/d
8M+PkpqVBA7koB2SuqiCP5pq+TmHcM0iNOuR0UPsxtGwvXh9Z4rlph4f5CtcMs6O
6Gu+4UWv+QyJetfaDhEMV0HFLXBFY9VTD8pvMvVw7pMadSyB1fim7+YHPbpXKOss
OXzRMky8JwRcdPsFPZkS8oRpN5FErJYVsrEckIFtpdLNvET7L82R377rDIn2tXmN
yDdhDerDoJ90M6BmVZUx4bJfRz4GFpwbZFhmH0Lq7CBT7CxKZRi62Lr6w6qUVIrj
+y0zjp1BYTurv7RoTvDw0blDeP2Dee0oijUviMnpgPQ+Yg7jwZd0ccP2uz1lrrXW
+nkVsh0O4OY029JyhgEeH1puioG0ahXd4587yb2MqVhr4GdK9QRT3+QNAfc0SFyU
3K42O9+HS4xS7tU/YvwAgGctOMg+uzRFnFzDOdIyyi/dAphnQlQSkwJrU9QpLpjD
NbzDFTdFIkzyha8GNlxbwN6fd3BexR3db9uvaa1/C6OqRkNcuIlIOQDQmd0vv2M1
UVrtmuT/zF0IxLpTqmnUTpsEqNTDiPJPFnRSk5ScBkQ+7V4qtM8bYbdQxOnSMv49
JbnXUfiX53r3xinl6X77p/50pzx1F4Y5q4UXV8F+TCakOezfO5GyYrvpFKJWmeA8
Ie08NgHcIJRaXSJaUjHVEd6wsyAJU/gu/6ejs0vkl+OTGypLzRzE5brvDPujWVbs
vUb5MsB/8crJB08JzBkK5wmXAJa6+zHTsCU4uxm/oQbXXI3/Kg6Mwn7Aan8ZBn2q
oGFz0NoCcuOoGbmgQPymglCy4qk7zIEjWbwp9rJvVNcAEGyeGWyzxYqgpQSR9/71
sePvo6dBWpGF4Vr/2i94Cy9/G9raEKOQxPee5SAPz8tafyEzwdHhrIPt3Fmf0niy
n8o5KWeDPfy+ifauukPZki6+LCzkLks7PxEuNQGiBHaRMLAUSDUf6NK39fAKYoC1
RRca1fBIwOCGzNjQa1eXmfKn9gIZFEuIHhUw34ITYioE/lK+PDp5P0aZdlfT69lm
4Grt79hC2iRS25RRy5DOW8mrDT4n2f+9Xz1laEeg4tiOVN0R6VkorkWaCQMybsLP
yec28AnVTu/ABGM4voYY3GaW40lBemcZl2ha2OBktuq9mYspvCw9O7G1QZyNBDGS
/3OrTCDmspRXn0O/1dvdM60ogV5y9NjxPGfuJe1CVfmrIij704E/WxiO9MiC9aQQ
MNkrYQDXoBHBRzyIFhqEF7NlCaXoS20EpFg8BBLT2vX1rL/JsadZ5MDZbxzcMTF0
7sym6MZBnjDOhPcJae55vIkuh0tPorPA93EY8MtHUoNqTR7FZDJ4Oa+325tX+RIu
Q+HsIY7PCZF+h2qNoG5Gi+erc69e22cZSVCO9vHcwKOh79FzpJ/RYOuLsORVbgXz
rvkMNOKsF/5XTN63eEOTIy4utVY7CGEh5CdiFM5Np97kZm1/mH6E1zIHlr43jj48
ZRhs4GIT4qCDyjyfsE3i4p53QRjSVrrixu5xOqp56I+M2b21ftNuwxlY2fdOJy8I
dRF0r49BYKR/4Lq6waewMaAoX21S34jZCBCs/D2XsAyyhptfTC2lOTarnf1dOKv6
WHv9kO9F/SPRF7jqQx5leNNOBWMrKi4laVBwLSufjY0fnOshsGG7/JNvn36JFie3
dvoLUF7GRfiM9d2AXXZgNmJv9OKoZFyFYfv71k/dTE84HlUcftPPD09isZKXLFW2
I/iQmhPGdn+m6MJqzOlNhyueojtyn6+S3T+n8otYkTn+noQwpIkHpM47y4aRkjbh
p7DNs1kR76ASxOp4Gic9dqHmgoV40I53DA9zoP8JXQYMoYPfx59e24kHuACBVdFF
8nqBxIQWcJ2NiVxIJwldlOK8AnpmX3ER+a7yUEFHblzB3PbcZinCPAf9777uHFZr
0T1Vp5GZezLdLUr8lpfefbVO2hhIzWXD6ajKiWWp52JXv+zBAtIgxOaW4UtItnbc
41u5PgEoB8Gp9uSlN2vtU+ShQvIz9/azhG9YnWR7XQtEQ6DqbTc8tmWkTgMq0rTZ
UVFYlJw209qOGLUmWE4XI0xDUpbtSFWf7O6WgqXr51zhtC8Z7yXFY7flvMMXntZZ
DKP2cE2CA3Q42LqtKord31pd/yfY3qC0Ui7kcjYpp2AVwfeZOoFa5pKHhX37HQEa
uyXl1WFcS4VUX/KEwX62lD8im6pZHzs0uO86JED8a7j6iW4sInANDKSjY/1CPFJ3
+/16MoShjP64KnyXY3YfM9tsnL+IiTNFguOMGatnWJmZ6vCUprE/V3V4QP/Xtsyy
bJOXbXXnBtAJ1BzXx1ALcg3nOE7h/cz8zSornG1Mo8f1eIYuAEnWdAdBQdXF3LTG
qutoZ4vfdMlEiIvI6bU5uMilQcW4WgMbzCOCvxJlU5KK3uuJfurncULvFvEG5LAM
8Pu0HaWD3IZNObPX5nRYLbiGSvZoEvxlCjFM6oI77p8nPwiEj+5GNxTuiEg5IN9Z
rilAFlH0ka73GzpiVhWF6NJxBE+p1U4BdobHQC2D7ihWs+h42MykMbaVs459Y0HA
v7Md+2vpkY/lumfp8MP8uhWR6RQVbXARQkpKcO3AxXctZ2qnXZQGnG65l/0qEhMz
hLSjtlqKdc8B3sMBcpCTD8g/CypADEeoM3i2ZZZuzAgtmLYmyPjtRJhgNCfbQoTH
a+Fu/7JYaQdnywmy5Bh4Y/Czgu4vT3xu9HWhFMD9fHa4MixQJs2QceZVpeGrxuyL
CYIZvjHFX2yMf+sB7x8Zb82N86h8pA7JZebyRpTOo6kM9jWwYmbIWYuicsslobVx
8Dm6B7d5Doc4+Np+2f3VQkpqgcfel8jg5ddWSRVG2eCT0qtkoJWBcBAMEg2dIWak
ch2Va93GhR9bzpFNM3k3Upcu/w7JsiOdfxPsQfTPokNZ0xw+Igg6J2AmIx10T8zw
5HyQCJ+8K98waJZnjBnAGJsZPhm9q6CeTEE4aKo3K+nUohX0SsN60j9aimtLbQ01
gfuhw2p3BlKrUOdr9kjzF00n/14O8xUaaOa7wjE6qmaxns5YaWIQJRuxEH5/jIyt
Oww83J1XmuCEoqkUUmR/PObmhRbwpjGE1YyGB3qiQMywHP/myqX1sFpL4l6n40rW
PrfgLwmSC5KkFDVo1qGSZVx2jqXTnd8t5AlnZPJMcA01Wx/OmoVsanMm2k0vKbTX
GaQMw3eLCzCrPsu4EQ5NUAeEIrX02RQS6IfDK5tR1L2wjhcGswUfqMZ30PyLepXb
6fdXvA/VuKmeyehqaRRLoyUQXHmkFUKTLR5+0NZDf4VPxfl6UlLwBi81LU8k/mVh
1caKtHvwJjvV3IqTxgvcuZloyjGqi54HfV25alMWaL8xTU4uoh7oASzf5ifBfinh
R4gNBZoFg1u1VumlAG2tCYr2iiF1j/gaKFAklUwgIc2AaRhRUA0V5LFN3G54F05P
Lpel08PN8NZgGOHyERRXiHCcHrh8mdnw7S4r1thKmKMiMUPrX873n7jDCcVoJ3t2
mwi8MkVRheZudNpQ5T/WoVFlddIiGswSp7/QN324wcApb0sv7riJdhn8mdWeLMZd
JzWeRGcNML91R/AFDF5w6dD09PT7czpGd1yRG6tCufjXjnJBI2ENWKIrZnZzQTez
+m4OM3knjbQNUp1f6D807hvzEXr1JBGtohC4bR+8C5JB/bvhedG1JGffY/elJ4YQ
fmRfvCMxjxFt5Qq9ERxcYAXu4/WvLMpuAtjvL4tkH2fTcWYrbca/QPyL0hSNYWDB
Up4uZ7WnhUN2/8r1OfnCoNmUof2PZTg9Huakg4xCqtU4kE85iKDGHLO3tThy6fjD
05QjUl1CiXXxc9ZnWESo2IgpIpSx2wBQsU+0mtCRlOWWuoVfd2y/ZuYh8Pi6wYUw
6xZwUOnEzpxLy7KgTSXdhcdxK8E7f+h/ZYwJ0bhhxEiyNQKp9aeOHmo6eOiZNz3c
SYXHqGktfYHfNuAkO6HWz9DDPg3kFQ/E/mZ5IZg3+WxZj516csgxp0boqpQuS5pC
0ffYZOD/IGvniSlU5X9XzmqEDK0kg/lNg8093Iu0D60DmwrXuGQ97ZOY4cbZueVo
CjYeT8Ved0f9U2uZxBAq4gYbmF83CEE3p9XxubtdIN/QWs13wQw/YCEtuMTkaTBx
WUmsUJ4IyUELOPbTj+LFRzCdIrL0Xp85ZceMfvb2ZVGNmoPWNw7RE155BvdZpQLm
bqYqlJjleGs7cm96O7Lx3+BXrAPe0neEFdSoqRI6hFWu1diQ80k1KndOX4WPOVVX
HpGbInju6Cmxac3lhoJoszBKZlcdw0wD687r/Q0EUAzK9xbnoYel3JJvB5q0Yqm4
2UCafNqPyxogXaQI/lwxpZp/UJRo5hhUgq9Z/oHIhYe4K9Rpcg9XMFFX9yTExbOi
a/DrmxrpoM2LWpkmAUMaWqftHs+2dLhdRWaCjaH9UZ9RtV/fve2IV2WIHLAfCW3F
upFxUd+OHVHWRElZ0KymZ9Q4zZPqEECrc+G77YHZMaBftahpfjj9jGqfXGpF4/Dj
FqBH7wYbzB65uY9fjUaze5i3XD6om5KSveLpx+S5Bg03fLilKbk6qJr0N/Mv4PcZ
EXyoFB80cB6ima0MDeDkfa45J7Sl09m8XK+8owd9dNWVVKY3oQ0CDF2aNCbax4FA
I9YM4fSIdgyJ7Bz99emqaS06BTFFcE8Xy9kg4XPGFzPDVwCb4XY4307MOQ0ytLr1
ua4ZYeYhfFAqP8TQmGsogptXjmFpyDF+fhWaebUmpFD/Jrq0xteMyyyo9CaDkS6S
JqcqFYVK15r2Pl7GoA36qev69Nii2C3ENghSdtHgrtnrpjkWAWMmW1qsXBcml8Ni
xTTydtC04BmUbW4MX6Uccib2jYNFWQtcMQX4j7DpZCAJm19Ai9gTAJzQMJouFim8
LCIsY9WFM1OvO+aNDxfuiDes1rMbHX/EDenCNrFQN4+VwBkI3EWS5i1UHFqvb8vw
qYYSuInZ5JiHwk6CxnSGPwYVQoHGssNvkB676U6QIbn5InzY/N1PaNPsbWX0aWz6
DID0tUDPuk6LSD4pPsKj6wa/CYJD22ThbMrfuuYjAEvAKjyOchmUd/PmJUSbYhFX
O4Fhc/aup1RFM/e7ExqfPido3E12rME5D556BwgA/C1etHH7URJdkkocTbHExR3x
7twNcwNja8lbLQocfPuC+hmPAiiKmZR+JrELhOs9O3qTgPo0Yuk86rcu0lcJzxno
7VAB3XcZfdVhsVs7Oxm5UOSYvvOv/WRr9hMPUSqsTLNUgCe9t3LaSC28PFPYy3xv
+aFC+0j7xFaby0xThLXAVQnQQud4i/MGFVLDm3MIkjIJhs1tTyq5muHOXnc8ginm
R1TcHBjZRAnWIMJ/UHBcWfKXBemGrw4UPzqFVbdVZZOZNVTvWtFB/LafnqjDm5/L
KixGDt4OUdLD74bQjfbkvrSgFs9hAQkPXqZCwyccYVzflEyCbsC79Mzw1rAqB7US
HwIqoX1H0/qkEtL3nZ03HCDXA4WWMUTi4MlLVE1bbchsG9v0pEHYlxOxHEREQnXi
R7SxOqPOEqgsBreAb1Zwu4jblta90d7Co5Qj+6JwjMS8zk7w7qqXzLwHQ0+yYFbf
RxA3K9gs0qS1ZEPCWyo1Hi7mLNZeHmzad/A+L9Fawd1K3dpfLksLyQm+8oO+d8DS
mUBIuvk9UEU0pvLwtBb2xrkPPz4JAeM+08kTC86xI9VQyNxvnnytiGsbDeaagNED
RoJ820yVDoRNKDUJuaiEVniARzqWM//jlh1vOaHUlpv/mgKsTmHZgdFvvgxUmJv5
rnZannEAexssQVqERdBomC0p0vFHQSeQZ+Yp3OU8y8vv6yLZK5DgJhbOpssT3Gdm
yFD4yrORjob7d+YUGkb0FH5dgdiM1GVXg1iRJhlbMzXiAZTFXP+VdEP0p2SdR98l
pAFEj/fDI2sesVWKzxjXxuvgX3OTe8GxNLX3cl4whKauYZro6N7EPye4Zwi6QTSN
oyI157HuA12zle+FJJl4GznHjm5gsgXP6ZZ5cPhIOK6nmaOvb+as1K7FGRNVheS1
Goz0aUOl50cQl8xOB9czLTn2IT+9VKktk1tKn5h4Zj+NEl73EbFUAliU/JnKiIZY
5f0BJ+6ryUd4xP5FoApzJ0NWNZ+EelYjhI6IJnETRZvW9JodFECs2Wtd3knea6lP
3WLYkJzrw2CEhDOaHk8Sblyc9Wckd0rqA3FjuhmBdmKmcC7O0Opxk/v/qC5h+hEF
HjXGHXaX96IqjKcslzYpLvBYtFJcrXou0/R7/g8roeXHsT1oDCK7Fyuyd9uiNWU6
24ljklvMNgF6L/eYy7VbGJX4ARt8Dog4atiHKaFoz+bJ1QwnuZwaojeSIZ+gXj+P
MHXpoGxlln+rFIDThuqAUA4XdAEAFAl2NgH+jrVCUpYWmDy0jn55rwjWv98OUthN
m2WCRunh/TJ4O7+vSVK9mzAhGx3JbtFnIZ8UXPN7aqiN5/t/yS9JzUle0qU8Mp5f
boGPE8V+Lzej0Ke8r4vPz1Vqbi5wTn1FpccZXutAAfyyKEmbVgn9K0p4raU5w5lp
C+962HD+fgaQN40ppv/l1t8qEvMz4Tb4QcbiNvAWDhJMDkaAn8NPu4RSgj7mVPVG
MVVQoZ1ojcVhznGX/764maWCwZohLdJUeRpZ1udo37xG/zYfPH8vDNGviIsFzJQt
VTxDPR1Omwq73sCEaRUk19sj/qgvQ+5h9L3FZMwGC2jpuIsW61Qe+i1sbpGY2h7d
jqV+NK0hpQtK+n1KQzLVg5d8FP079MXhPth5ueOvTpWbgF3eRcusBydmx48aP2Ao
MqNs27c0XVdJqdCPLVrfhdqkTwZSQ0Qb5Hp8zCUh3iTHxjA3C3vz1+1eMubPDxQM
pt2hTO2AJ7cfD2SVQh5hOxWi1x0vZ+qIFDLc2koyPM5emRApD/OB+zmcy9QhE3bd
F+qb3BiUyYr6VHT9feDtjRufcuW66SqxRechqBNwwSDI8lQH1GyaRkEljtUlzNHb
pmL7uIfQjWbwqof96Wp/w8T6iMg+7ScwGZ0Gw+uRK4UTE1rPR0Xq8riZMKeVrWBU
UFTP55Lz1lYOpRx/ZNsI2mTATL/yJHfcDQ4k1iE1K8fQB6LgKI9gwCoXnBh8j9ZS
vcnyUtOUFNTdMwPOXr492mxDKalh+rbLEXdtMVxacHAZoiGaiGzs6+ewTbP4Mgd2
kmuB/rKG41fh9LFUtZ18QcMIQv8TvaVJReHeRvsL4OnZ4aqyOqlBMWxG1hUC5t7u
mGCLVg/TYuPnR7/1FYDRMuxfffL7jlH8cOX5JEtQzjlcEXiqMzEqX2uT0OCSRbZS
JoZ/DN2jFZqzj4Z/PVOyikwBS3OerhdOYIGxym/Nyefqdpld4eeYrgXX8WmDHnZH
WvVu9LdQT2jEwcBObL+rF8BwXmWXt4LgOTTQ/q7+UK+OfI9QcDD7eily+Y0NJNLe
xmFZbV8EGpfITCCg1ZODRFzRbErttv9eQWjdpaegCHG6tWnSTpVL3ipNCmTmqxL8
cnlnZurhzO+ub2v0B5pFr2KIZXI02r3HZzIqGBJx2BC0zqhAad3QUFc7VXbzXxCF
3L8qZoYQwgfjngjQS6E/0iMhBO0ZdN75vBtt7Ozh0FMaNJZqlcZAAOCIjGxF0eFa
eUvwlGDF29+kV0CIlwDvMmvSUmnZWk6tgLvDR9y8Z8GdCgPhV+Chieb256Bxcigi
toYrr3EdSm3BULgdRQbJYq8mMxaMBEGQUQz4ZMqBlWq2foBLILPzyTe/S1kAqc6P
7m1LqNAORoycrjMak03yjSdw4jYgsh41ZUzRhKvumf5jav5XJGW+1eDyk0dH8pmW
ZCfu6rMxKF0oCB84R+0VH8oGmWq8VA14rvWP9JZavtuO+DZJqNVLFRBYYlQhcgNU
eWUqy9nm3kgVNxpEruqELtOMya+pAy2EIoViy0cs8FXVWxaSiTSi0/H/lxdPGcJ1
PTVeavcnJdKQZ04QaZQDByuBHBoff9/XVs+tgMIFswsGxxoGXc+UUtM9v2QiFcga
AvlAzvwHeTrktwOCeCF7qnCTHPFc1/f3BQnSUQeDiBo+c4ycD0wVK4N3tGhhh5oK
NqGzBZi6oE4svmCyqokcBzfOmezU8OEOguNhkOuvrRutcaczIYHpz4owIYklyIL7
+qi5F/7UXGHy4vpDo1cn0QK3C7ihIpPL/DUIri135IRBOW1eVfcs8BxBocfAfVBR
FskHqtGmdgn0Qo3upPdAn27u/AggJxA8S7CsK5VTDGNDlBFntUOkVzHB5lFOhpPY
xX5xjMSTR/aa715pNXB1hJm+8Vv4tAVF0VuEHxsHSVbduyFOxkBR2v2d8e51aDjJ
fUKEcdrVrS3UUjSPROSaQP5oeU9ozTooVrFeTxNqHoSU5hF+6baEojBGDGOZ8wvT
p85AX/396zOb/6YKcuHyMNKDP7MFX/KbxV0JjhM4Ze3wdQ7hVvlNgjzQwx210bqt
Isou7qRbGyYkSYsq3UCUdYxFx38FwUSPJTYlNwfWTeb0U7NA/tmx+1nTuX4AHgjt
9NIYdeWsS/Gixlp1dEVKL5ug176J8JzTIEZ24EsrtamtPgVhtbJ95QyP1GFbCRD3
tfrD7MLN2YFO3lwtAPQgSWws0HBq0adLJCFKQljqCe6P5XdGYHD0iDmpEFIbXNmD
JGcwNmSBtNp1fydsG9FWyfGM+D4Ky4fx91E6DQunfZM0ZSaufUJqAFgiTOliz2PQ
bFDyDrFw6YXNP9e+NMs0jGR12oHFdDdqeqyWNLlb3KOpSrSjror4NJFRcZRY7rzm
jc+Iu9/rBN9nQO2Fo4Z+NMK8/r+JLYxNDz1h56gUnI5RLjzkTGp/phXNCbXRKfJ8
D8fcuODsRiAuKelG1BB8w9fPxU+UpPYwFAu3GL6qQ2t4BEvJDSIsKfNN+X9KnxB3
4kArNE467XUwtYhTfFkwb6m813MKypJcd9SY+dauc5Zud9CHphj5zEJkYUedL1bw
8vH9OxmPx5TMuwV60w4ZNaGtdKmkcWnm4GticUP5Ahn1NOsJhvNv5fDKfSJp0Z93
wmhrXZ8bYT+Htq6KUBARlh6knxSYpg86jn+MLPKJDkK9nSNxjZIshYLwvbyexF3f
94V5NHnx+sRGfcuUQUkrBkBAnwkBsl1XeOa9X7pI/ezdczkdvWDVW21z7Rtv6N+8
x14a4pEbJ5wSkRalMAqebKtEIPG4K1MWb0XwTvPJiI+BY5R2T5MqvmOyjNYtkQlb
5m1znAc4PG0HeAzIUmkwVzpLL+KfotLqmURK2U0Puso7XUYls/Mx5N16YxVaT9uY
q0dOfck+D1XjsV1um7isyv25FDWNkjYSelQx+096Cng8FeWEe0yAtVu2vqZ+UQkL
I4mgT24QI+50cHG6XN3NrGXWW5oVr+wJcKirPVfxs6VhSgKJLKyIbenMBqOqxqJZ
qR/YgzjVOsOr23mHFIDalYpjsmi7EJy62rWEOeX3DPRyakeL5tsSM2wxlJHPtGjT
leaXTo9/iIKzQkVDYkcykl6/Z7QUdZibYq4NTBoMcG2zx5smApg5p8RkznP0dOfU
W7DIoT5BdUNfn74ZmeeYFSUE+/jF0ouB9+L9/WJy7nwsLvv7q37dI+EtGKEiNMXC
gBuRZwW17JIQ4PnhEY9pqSVkW7jpxwW33+mBpJLy0f+mx/gtUyPhAHKSm3oKfs5y
QtNht9tbNeJHcWaKPVdDhgb4EKxxowYHwZIfFpfcw85OZGPNohkczW5CQV7xBObP
ymKA9DxSmconhTf7AZXOqrs95yjEbKCl+vUsFnxAtKRvaKwRggmjOYvEboskfpR8
SR5hTplIBzKQABHXc61MnioRo3/DzoiL0NnPyPkIbg1cFDjNYwIwUT0jWorcru/A
J3CrJm+uQ04EzqdhondfNtCOuT62TTeSWLnHyVFQTOApfVrSq81ItxAZuOqD/qMY
YkXDxRiA2a16TebB0WJz1qESBEhDvWCB2qovTGEStUADNmrxBPVaTHF+zkeU/s0z
0J1x20lylChWPu7+CdXYGWKlCFjr0v8bf0kZnYvN0uDabTYX9+VtjOW1y5Bzjk7h
jkqmtb52vZTAxbpmiqx0X0K2TKUz/pNjwQndiVatYSIT4OwUvb48kAkl337wVIHr
iIpSovVHtRbaA0rsbh5N/V3GDIkSFF00ApptBNm4DjIszTMidbf/EdZ1Fji7Rb8y
ov0nqMGvfDjMUUVnKDhXj8EK/jCeO3DXVQGp+ErFBjWZehaJSaDnPTA7nH9jMgzS
oUBtLm8D2iW6wd42XE5xLvZG0b4mtKEW8NI6Kr2VX+8qg/gQDjCi64Sh6V9qC0Js
7gdshNAXDYmGYuFlcUsVG2r727mrRl3JjU9GorkiOGHh7JWN79rx0kpGkcuHKW3d
iC9e9i0JAx2kI5sC8PHnbwOtUW7thB+EOiHS6QL3zgY+GzGGpbYUrt8jvAd12Lpb
cBAzzRLupxOtIoRE3OBwzCH5Q14rdON2P3jpwsXehclyrsAZxrj5Hj2BtLO9zY0i
VlXcLy2YoavRQl5PeA1VKAoTASfRLOIzlKiVXO60uKUgDA6U0yfvk9yHp/BcJifL
06P0JzM78jxfCyJmLeRhkiUW61zdDrNppRyjLZ5V2DbbhJ6UMrsjvYUC+xf3EhsT
qctPNex9zyboHa9733b2khuGRqVZNlmAOlKx8TaT/d71V37TWSf8dwSQeM8IhZLa
D1JDu9qkmqbFuPuNRNNmcgmd0LRJBBx46Hio8AUw3lA9GvICN7WahCAkPAC4+Uio
QXvVLA1W+EUwRWogZmdJrNzcLTGS6GtgNECgs6TJrol4RVeQ8GXyqTyedw/2MbWD
hcBsAQhNAhM4CJ211iu68ZnJj5LJ15vnqBgAU7HgVN3WhDQYQ9RHhiilJxFFUCNL
u8g/iEjY7dlWUzvmy83clt3gdd70UJhOviSrqGbF9lH0UWq9HMgCdtOq2sVWMW1j
JFyyF/AMHVAPrQYmwfJHATgAiqQCUzcKN735lcr/jP4XGrUy7VvjuTtGXYK0nkkX
K69dJALS6czu8TYyT/KFPyP+RGKwfsyoPDc1z1/MAmmdPxxoPC00QCdDeumpjcVm
E2AxFMi4HbspGj5K4fURLoWrp4exSnQD6FZRX3RBNp/fosywWePd1rgWfcWyBmnG
bUUTTW45MNVwbPk+WyYy9OvAbQDuJvCCw7FggQL7BVxppJd0J781LORe2frl3X8J
dtTdZ9dPcJtdMlvtxN/1zOgEAM/2ivpQUXiEgTgdecdUBilHzCGeW3KUEAvI4fsp
sSeO857P8IZvFLnIsCG4fGMZ6K6by0msRiUTyww5tRQh9T4O/wP3fD1cvbLfCATS
+Nu+Tqr37Qh1kBGAoAN4BC0gY056jrhefK79KjsKYTYntplU0yF03dDOoKNZdF+u
Z++PqAFp4D/qdbFQx72EUZEtGXVmaGehv3bnyOzLDG3cTYSEFP8Jv2dpibFn44dh
cK7vcLA6c8YhRyqfFhAtBe+CYVGEBXGScBB4kKaPTfavKCuYH1ybo8z9DhGZIv8G
lpckjWzTdZIO7i7ua7O06bJf3m52RxSKUPdFFONWijRDpm//EFi0EkeOz5leMqgD
PPO3OVmqAAF944VH0nT4BlTIN2K94kmRiMwkrjNy4uFuoigGJYdQkU+6HBOrNCDs
rE3+byXBQzu91j1AtYDKKosNXpP3Piw9xFqOaCgqCADPSzsFdPVJ4J3P4Ru+SPWJ
syPAwi7Crv1VxVtF26ehkzYcu/Hql8A0zvCJjfL4yvoCLKlWYQ9OD6L61yd5uCvM
F3u6S/Wg1wlq6tEpuVTXEB0ki+VtObi2zwHplS1UQhrxOSpVQ+Unqy/pwK6C22lo
H9A2KZRek7wV2FgjdlCdjdbYh7wIiwZ6fcqjS7SAzKWRhkLhFVHOc1L/HlW10y7I
3t0/DUarJ7UI2+Npotmd7m/9X5WJ4XG4DRlQWU4Hr//ZocpHfKx0K6AyXtS88sCV
4TwaBGJfyqQGG26FIP5psNV+WsI+n/90jXDwxzj84u1FyZvlg08iXNqtU30M4G3U
oAaFX5wokuacRlKZ9myEH+S6uFb2mCl24RHrALlE9YOxm+rvYzW5FrTCrQVxLccn
Ktw5rzPXQrjFQq48eqRbENZNZGwcaxrBfvPFB/us2w3/Bd3w09Jl8J78oVwmz6GA
krvmz6e6sy8LedRFnOYOT9qSUYwjGrrmCHm4RS2PmKP7EOljQE0CjjxksXH6Fft6
5INIcEu3Mirs4nqTYrywEkguMXotIIJEsNXS4YXMK3SUfzs4wmW420/Py5qtqUOK
E5t/NfFSaPk+kTz0LHY7NuQ05guTqFjgTGCeOg3ve4/GPM6JcBjiB8tqpYNp2mfL
5kN4MY7HfOpsjhSodmNp+TBOuK8ldMNLlPTzESNDVoB1wp5LmdcUIirKAnAmb/Eq
D7gKKqJ4oWQtytk2ka44jzoKiiOg19nFeJkcN6m1tz33L8lyiNN1kjdYElc8Xlxj
DSo2ezJEWVqhd37f+ZId4uEzwDu0CWO1L9cP229n7s+VNtVbMgQLiyPFgplhH5+L
OU7uX8z9IzpsZRTOaLo4e8JMQOYTb5BF4Y0Bo6d2MAArHPZoBnU9lvHSg31vtJgU
G6FI/AGkKFF6as8o/L+fWEi/ftSNKeM7W3y0mLblouoSYpwWjTdVkTw/lMg8sKVM
E+CBdF+mbleIy56CRlegiww+ovNdNooILPiO+ykFyqhaNI2AH9DoLcWqBIcoK2ax
n0Ph7gvv4/a+0FHTGle2WvNzaubEt8McDZe8yiOX/ENvmBn8itMf5N+CYByMGJ+E
J6l5TTqjoB747CzkYbeRSO9pIBkLyCcM2eHiWpfOuuZR2EoLQmwmwMMoMhiVIvoZ
VUAo5AdgEDXQeoZFe4gDDBn8yLmd072C1CnkYkkS4YsXyg9w3Hw+05F4NJpEd5sW
ZYiRWrw985K/kQjrf8jSwlwR5Tqm0GmxRfnp6GiVAoIP4bSmhvsL5u+28svPWQdh
32nfhtqL4aB8NmZ0U/RvjLItYy1LSIRbXHyXrtNovpXUHrivcCqXnvwgeCNdkP+0
1G+EN8uNFYrzPL/2mbjIltOlLvZRJ8mjRS2al6zbpOxz9+Ix3Bsr0+vZ3Tk/S+QM
uR0O4FfVaUSKPWgG6/O6C18B55E5IJmE10AAyRWcGWT57D2gmeL3/41Zc3D+PrTc
1bQzyZ50d6PrcQrBZVl9YUEbjAZciZP4G0xu/lXZgCQhc3naW/grNUro2KgRPvLC
OsNH81GqgYOrapoHJr0TbEhVUcBG0LjxI5vrIgwyQ2liKHx+pQt5I8ckxzgXjDft
4WMeRryPzpS+WDkIMWTjnMLubrlkM+3qNge0dFvtUbzbrhDQH5p2ItMawqJlWlU2
JTl/6ip5+Trm8V8zcKxEkZ4xyynbC/gS8wBCEiygObz7LA9FGCtM93LpjpHxgbCC
ZD+Zyuxdcw6Ln/7zK0EFAWZll5SbmKTpXrBTGpZ7zSgaFfnKJGevSiZuci6Q2Mqu
KilzhMlq2w4UTPaym03bfbjXeU7mEFgLJj2eank1iM2Z1roj9FjWuA1QtBN+IgM5
juY1a9/fPkaLuzilb7f0gDbc1ptjbfJXg7UjfqJigP2VfLIpNScM3AkHcNcfXRoC
VQ4znoK+Jy36t+x9kImw23VLclbCghJQlh5oKpnLZBvlWwOPzmJmg14HP1xlRUlO
qRd+yc9mf1YkX6HbCH5FLh8deMAkeKetPKbWJfHPTHqzJUZaJzzy74cxajHwq9tD
61FT7mSfJ7fsnyQEbx6c6XPqOzt8VSX+60+7Ie3aV1D7SSDMHFOM+HTk+ZCvMPaa
gvSUuBeGP/zyaOweYvyZo61Mc5g6Cwank2bsYjxrStgSiXpWLUanG1mO3RH/qB5d
t692B9LHc2J4Z5sFIxMDFKv/2/CKuktQVAtR1ilArcgwkbT5hJ1fnezNEoQU9Vsa
tbCiE246Wx9YADf5+waZkmcjlwUkUuSr8SRfc2zY19Wa9NYS+tkY1LBSmiPQO6/u
Y0294qRISSXkI0u1mhLbjDdwj1r9P67acTsg4BuXALUgdHIZpeEViAs8aGHNFkSk
3FVvzinz+9PnfEjv9umNWAS7J8pxcDfeVmL7Cbk42ILlB400z3snokz2LB4t9vVx
e7JQC2BHbYlfOteF3u3WXPqcwrUIvzP4GzUfS8rhWAGhFqKfqpxe9X/JxABmNdVL
dfGp6qm4qi8sTeDygAQ82pdzsKQtCNKtBqDvIgEirDCiqxb5IWgLFcwGUKgpQhY/
mGdbRato7lVfFWy9lvKdVA1ZzcF67swalqJLcWTHks+5hCOFdRfUOn8CVJ6RJ3PQ
M2B/9CYI7wcpSXI31hZQyHM6DG5bSmAAly58S19mmk6qAk72KgdMTx1Pfq8jMkFG
s3irpP9lvzkg/oC3OaLpaNIf2hqLyBDOO5w2yMLL2o3XXHrNc1+ieuzFTOQvYYtI
rYFPR6Fqn8c8HJxhtiI4PT6PgJFCTUigQJdFfJolmJjf0wCIRKr+ngpfdgQUpDkg
W66N203dw0U4TBAFAwa9poPsvna0Sqh3DcKpOd1vVIc039xlsV/1ZBS3u0StC3Kq
9C3/zoxtuaGuDnS07gLdUXvGAqjDkffNM2mGrVR8dhWQ40FjQ6i8KUsHg4FY1Z/C
Jj7087+uLDEyj0gUS782FY3h61t94vKT02u4vsT9PlqMAMI0P6eVdAcBfNKBeJp5
M4AaKWZFEk+UaGk4FlZ8c8sjSHsjWNlfncYQ1Oh00m9zXUJ0kdpFmLeemZCMVxcT
EKjH5NUmGlaPE9eQiA2X9i3GjFD6HVnqDMPD8NTi/tnw188FHYxCO1d2L4Su+euV
UDcgPNVgTimEipzl83ioO9G24eHlPAp+KGMpa1/lg9D3+woY7DKJBKhVT9R4RZQ+
XUM+g55p1TF++h1bfXpfn/9FV0qOLj2zYeu/VjSdB3hVjcgO9kdC3/PByyKc1Qvx
FaM0W9xOK6CzJUyh8jUx7rwQcX8SaBDwn+IBEttR1z6yZzlMj7QWevF4H38JM3ee
0e7eNUrPeIN4F0fsgyCHnk8+G0x3kKcFPFZGsH91l4FR+h9mQJn6NLtN3Bb1Qe3w
MqfnCSiYHVgZ9XxgB2WsV3DmFxw6wcBgO7p8ir7hBH14fAuyAtZkOfPfUAUTrNm/
eMLbFK7AqbEXz1PCQ85+DEpjSCmMS2PV5e1lHJbIXRcmaLxusEOiEuEi6CX/k1bf
XqOy5YYVADNlQbAL3Q/6Xrlrnuz+JZ6PiJzjzkEPAOR1fe+0cdJf8/AzNuIr+xNf
VMB9F05wxYpPsaUFCDEx2UiqNDfszCTBzvtHGryNsjT2ZGlIflcFzUxEVwh2Pul+
E4ak3PWQ+1FuvMOg8mQIqTVodHciOVDPCd7unAdq1PPBcINUOvZ5cU5bLRSemPvv
0ODqsXQdfYi6tXYtdvuDxCURq0RbHfpn0LEIVmVLuO8zxUJ310FPANDaRbmW30Aa
MMdElM3odoMCsQYchs9VAPd5TUhpKayaxjn9mwreC4nMiuSF2YsmrxeDGiST3mTN
k6JTKMORR64LPF0D8uzX/DFMOD8BgiQ/4uldpJeZM9wQbEYvxl8uNDpjcp/Nwg2Q
VJp79xDLkseMKVt78OR4gW1E/3Uq3uzW1kMF6WYIzG5wBLOJItsg87elAWt2PuMJ
k1+HSFMboMBb27deXClQlqWHV3JHvDtrDaxXyFVJP+lD/NZmA17jnoXmbjSkxDTI
rGau5i6U8u6C5lQYqDNNYkIZAW06hSgb5o/mNig8M5yCjHsjRs/ZVMV/qtzDoxgf
RzFU11i4CatgXy5yB5ENxdEGIfTTsnsH0MhXCFv11+k6UZAnj4BJtJ+qItOj/nrG
btr3pgrhYmzZzwfvNUA3yZz24MSC9m9dgAzcIj8rmBBpkMXF1uF5K7Gcybymyl6j
ztL4cP/2tGtE8bVLckf4yzrj85gPzNoC+0WV5iP7g8kO4laGKuXn4QB9u3rhuh0X
UO3mLbm22XKKnK0OxDRLVZU7wPwxGRKUGE0UQjBjIVcNbMX9mOWSRPUz7FEHE0vL
fRKuhXSGqmwUOIRwnvX9vGKUF5T/Ima79z0Zd1ogQbmzLTmkwgKtgtIu54ChRJnA
kto3XGQYz49rsNWkk7liIOBt3x4dymgzm6yJBRCrXXNrSY2M+th7sVhVFYAsz7gd
kSU/GWSVzsal1J0vSW7Wct96U14aUWMwTiuiw/1iwWs8cKanba7ECaPKsNjNTdb3
EDAzXHSQqtvRP9ALOvGR4I2fgrByBfIi5dUDAqHYVNtLfYyjvjBINBh7iZk3fV0/
WVycCL107eeRmmq8gqAUvyioItqtSg8+iFnUG3kIc4bHtKIejMlsUqAL1TnzXNMs
og3M5Hdh8954QIHyFN5dpVyJg/ymlaM2J4f9y28Jwi2cooKRSjO/nIp4iiLSvGKk
n1PGYqlKS99zSLGjNNwwnL43VRs6pCXdW6k1OYi/tiLgtQOi64Wn7+Is0iUdCUXc
qskbCVjycagGDSZ4mcx9TVZo9AnQEaNSX5QOFLZMG6Fnu/Xv5uxCMDwyQp0oVIJt
wNcQDJTRiqi8DZJnsPAKuH60M3CVug3NlhUu+RZlWpXg6Uo1Fdi3ngyI7PIFFooo
56gT8suLI8Z0TiHNb2jdx/9UVZv8G/wq/HZbFNNHeoSB97Jf45/WoxX2Gr0wGTYT
2miX01dL0cM7Ba6GlOKLB6DXk3RB6WnWFqI2Uy6jqhTshyP6vy9+xQQReTduUIz9
00qKl5beIpcP1wwhPtyW2ZlNuN73+Y4TddgYxWKwfkL/WX1RHKKdJU5Z5n4Gbt7m
O9ZhQc2ZOEXEaCLpeYeYgDFq2tMY+Sp3HMRUhP087FK+lwrCELb+GLoejytQ+SEj
u9p+Da3tN2ym/gXzsVE0yACFrHQRlHkzmsX47xzq5+FlJJradbEjeb/nPbBRD/LN
+Ay6/PQuIgjHHFV9xtgQwz8Svq+FvbBmmy1BtHqhKtnX7ARqIv1bAvtmrmuCJEJL
VwNhSbvG3XVZ8rxEH6e63KVBZdPgcv4dfCXTrZPBu63ZDf3DKrZJq3OPIi2Ek7wU
qN3j+mbSf/7nRZVKmbJxvyJXRpddXH2KcuLpqaWG4kQVVPEvkvVo76pp6kVgNa9O
u8enwlyE/q/Vwf4qhvhWXV0RnBu/ogUZ7TJA+39xLp6vBqFMvniDei6AsJEcpo3F
AY8krTryTwsiK89+mFa1KtJoDwnVcjp1IZKpKQxCnoaQDcpmBx092FwV/6bxcBY4
zQbkVhwhta6lxfk/w7q2EatGrQEuW+k17UTBWStFPFQTekcLwX/oRqxiHkX4vb1I
F2GbemlTT6THv2za1DlZFea5igsI9QhVNVcC6TGKxZraRTYeafVnGsqKSRQL8FLT
v2kNfWo95ARxU8+qY7621bi2sHIQjcb+03gQBMsFm/eHhCqyfYPsQkO+0cyTDCKC
ZtPKo258oeQiJ/7hBf5iU7MvRgyd3jwFEGpLaz860HYF7Nql2e61UMzk3M3KrEqz
wONd1bgGH/mkNfqLDeE3K+Qf7pKTHxyc86sIOko2b6qnBPz/tP3MfgM3BN2LMmMh
gYXinM1fQma3DmBRPPCuoyk9POdzB0tWKOT1VfZ7kEjWBwRrYxnkDz5ppnMpckU4
o7Ib9unR8naozgt0VnJJv+PnpG3oMNHPZXfI4fyUPD3Ne4J7ntS/850jjTZeCb4l
i7hY5mtIyRNewphWsfQlbfUbe3SwUnhV17eFhtxsxD4/otMCc4DwC3X05W2jXfOW
z0k8ws2+4fZR0bSdtFuLQQWVbE4hHTrumTOm60+SAuDW0Tu0mvqoNRXjO1uvyhMX
xj91Fslp9JaiSxAJUTMpiOCLVpogSNXLqNLIt4lzn67izXgl+ry1r2ZM4HePrvgy
l2alMe+RocOGboXVkRlOtzdiUa3MRQG98eGs3bDUEG5Ha70fwT8DtUDgwyWXnwPs
NZZ8KTkfXU5gPp5J4/Dq/NtNnogQ5bj0i9uAs31rJ+DwUx48R0yZ8FjUrTgQlCAc
y8JWotRymga7aBhfzUcyJqRv1uesCd4pOi+RYKNMsYyHW5zx7yBNDMM/D5oo9Kmr
qtJkLyC/DMZeJ39YNxLEqEMhYHC6/RrXhLYvcSvFI4e5ruY7MABZVdsJCU8QrUAQ
DnibnvuwuDTGhVKOiB2UHdz3cJ8/3mDzNywaGSQQXM38LiDf0uWj1wA/rhYb4zbs
CcINX6qszy7qO8X+MxgnDpu6zOfe8cy//7PghnQ1DzpgxQ8BCoUJR0PbtfZxRP1X
UCG9zmedMyU2JHniEZXBntAL2kUDbw8ruAR+QJTY+gCZjnSFu9iyLovGopxyUSAm
vc3SzBAOXRsXcmiYluqQHsWdHl0gQg5l/PLEeYhCsiExqSFjtYwV7M4a8CLHhTvN
WS0+4en5oBd7hSeSACeR2ubCXTKJ8v/OWxTt9/AjSR7k09km+zYkhIkdaQPrMEd7
0kDQXT8TlxH5e6MjsbYYoH5ijoPW5OrQ372KfdpUAQP++b+55NIZbETbBqh78yIL
rRHS/2gdGelvf2H+G93y9iPODIS9ACIDJ3+2jAB5uL81LNQCddPEtvtDI1GvG61S
iRTUie389uNqTseQs/WRJtMHh/HA08DCjCTjSoreEL7dbUt06Gs1ApJe+26E3TVQ
FJMNwxZNoTz6hTPdI2zmGcSbt0aKS4VR44GVJWyvqYQyKlzttrtlxyvdkuh34unj
ItlEQ5kPH4+aNKq8Wz23IE13Ss9cl2/xz9OEzDn7ZYdVx8Wey5pnnOkTjlzgNRW5
15zGM7BPTJBbr+FMyUrAtoDYI0pD0b1QWeKPwjct5w382yBVIcLqI/u674Tzimhs
+z1DLAd7yIJEQ372c0FovuzXAdKx+8TUzllVvmn1r73ip3/9Iy/ADpDw6ZsT/XVS
SXU7+FnaqJGKlqJIBJ4utEY/O/QTaCglxv60Z0DeuWeIezJSRNczwL7JKNKlu9ru
clkQazTSqMtFijJKBX4+P83JluF6JvwNou+SJpH903Db8ufAN0gzPbmNLirw69rn
NidPjmXEGds0kCnIdayp29s8ITXGYsbx4zmbXtQZUtGiPu4hJdl8qSyE/hft1ypH
WbhVOvo2GYQF+48ngjPfjRdR/WgOMGuijwfGVHRvBFNyAQez35kTuV9LWTgbaXtS
BTL6KMhn1psUZYgcZ53G9XMh7JdFZlIdc+Aiwt4w1e2UhnYqPAV33bEwKP+NYI+C
Hly2i8QicWnH8yMqb7sSr538STlbInAZQyhQwdeCtIzQSKZZABacE2rB6zmFbAFA
7g5xIE9Dyo2uSiZsnzmBcLD5kd0jlpK6gVYBaPlyQJ78FV1korZdaEMWuLwIOUio
d6hHRx0Yy6N2di/OqAL1rcxri8+ZKmgQu6twxzZ6rIIwavB4jf66PAaELEF15g4Y
8XIHojVVx7rSMbJ/mntybqC93bVwqtfSyE/qNx19F0B4dpKbqvrbJw9isGo4NQWq
M/UZEuJlrnJBI/8MGQz9ZZLzy4iRuL7Okog70sw/kDtUES3cyDy2fzWy/sTWJj21
uG+D09WRjG83xlwTRcc67P5nhz/eVpBColyNxCFLNkhsQmbba+fvQ2tbmeP1tafY
gZBAV5hycTLLYPAA4IVN5+xfE2v+7+4TlRjY/6vy+mjixqyBKmE4ITUVfvMqsbYb
Naw4/X1ldvDOBdcnC9H9gN4PTR7KjdF100SQXI4rd9z3yZ94DbQ6kolOOIesQAdj
lu8j20FJ1xhP6CazV+IkkxdCmtA+h2XO+EzK8wmuDMFWdjIzPQDKFQqxQSaL2X3c
Ew6vDQwDGrE1zlgXivLwqyrjUhTL6vlY9Kt0MdvGVJ0MlbOp3v4UcynWH58FvZOI
8CqG90qVUeArBQ575CiDT0BIwWTmYzAGc8IsLaTxnKYFlPL4K2vygiBv0kq1lQ7A
MLkyZ0Ds8IF0hNfHyvk7bOGxFbYr8zp/gpMHmRNSWX3/SoG0LRjHwbn4kns4IYGa
+iqMhEFoSRBg1umqPf5avlqqejOLU98xjEyuC87QF6vt3miWBkxy94F8U4iPkvio
Gcc7cPCXWhqQtEnM4Xmf1qqlE2LXqc1ExLuOktTRMvZ2vjeig4ndyR5xwwT3Wm3l
7fx3XZbgAFP5HGeCIZSjmytHj0iizPzq29zSw2nOQE2GS7WQodd5tjdj8qgaPWT1
hc6r2LPLkPee7S4cSaimT6/YtFTkyOxMBUuLnFHNKAo754tWNeDQRoGYg3tYr4ko
hTOfrPxmulWtV9XuM3sUp/aFaZKhFFrvJaX+k/+bq/ulLUGPIP3v9rxHtSRjE5y/
Z5SKai0jpLDuk6lVxwwdf0NNZuEmOwchXNZIpNPFXDxLDuQM9bjHnS7hwu6cPZAT
Q8KpbnBfUxivFsSDZOrZDrh7zzwpAaesZcSsny/GinR3eYAicKxpdNZ+xBnjaBRA
V5eyYi69zLB4/9glH4NONblGhj2QLH0o1aosjE5+KsHYXGzGly0koqnd/eQR41Q3
DjzqJqWbIcVNjH0NmV5nnLedvFYyw3KdeyHG9OxugysYC+Usw6z1df/API02u75Z
Yw5ZJKxP4+kBR+1tjdIzsc1N3Cc4TZlKQJry/pcIzyecONPZPdV2JqclCVCEnmSY
S6nW1qD8euVLoBDMGtriDuiyhrAaPq3fQ4WhcQ4m8c9ZUuAo0r1Kv9qCwO3nH5/3
bJmPzkcS/kzoBwCzoo4QdVVFdC3+4pF35U+OYAOetpy5RFK15nxxWKkX0cVUE7+I
dNwWxg8wQgJ+cw5XUlxz/OW38HD/WqpbwPjgdSA5L6eNxMpQCN/S+GvEXTMEE8CE
vUvggNpm301Ent5u1Yqj2QVV/M+oHeHLkrHd3MB9rLj76MezMcrLcBH6Dt+BwJI6
gkoNYqRzEF1SN6dYWxqgnWhNvAJ7q9VuPx13BSJz/DGIrra3KmKLUyvX1KR+ahgo
+ukotOHnfGb1UqM5O2DsgSE54juWKN3JO/SfTRKRpkKXIsr2k2z2Hh1DBrokYvHV
EfBqAeAVW9ZS4xW7uvyWiNl5LLlOg0YB+ggbO7l1X6wyLOnP8NuPrOqPaHXqmM5k
uuHCfPsPmrx6nRtuKgn20Kw3uNgGfGPdxm1BOKp39cAC6wCArppPEft/Hl2CpV40
Vs9/6Bk8+aq1KMyKE1KbjcngcdavFVEzuPTFDGGi0bGxradaR8OwKUhwi/r3JISy
7dUlD8sbb+lXFmUxFmXUWnr+BuAQukUnLunBaxE1S2A+KTJuMrov4LPEMBGM7dTZ
BK7qhWKIrQpeh7TzmSLUGruOePyAJLl425/nHDlZkFwTsT3CX3R2SV6auLFMPUtC
L5t4SnG3T6th+o2luN34R9jmMoHv5budbMLBXOI4J8s=
`pragma protect end_protected
