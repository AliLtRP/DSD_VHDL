// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:28 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jB7DeG5NfQTTGZWCFewVJQ3GP0gHnonFoZ55ri1tQLeNjclE0SM2YQ1Tnci6wjry
wMGiurFFXDlhFAEycg6Z2fFS80IOPPRW4XVinH7KdOrjgmyePx4AMxCNVeYpwmEY
kQaNqj7Ao2/+fnxE/GBbJE1oHz9vx9VKlc75tBJhMso=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10272)
IgiHeT+G5z1pgqgHZ7su9UE9HgZZsuzvl6Csqb4MyTungV0ZJq+J+SqigL5iuIyD
2yGYFCR4oUepa/75VVR+/pv2b3KFtNa+e3n1BRtld2L6a6WZxfLAvtR6Op712z+c
iWJThCw6yVYwvrtQgWxkVYVSGmQE5JoYcl3kfl1LkVp/dlmLx1EfPHn/mZqGo5WY
dBfBMLEzmO2xr/KCTWMB0LS87CxUJAutEfAeRK/ElC/CiDX/CDFlG1wI/bcl/8aA
Sj/xylk/QyK9LL8b/SrDxlkxYRP6bIu6jA5io0VZuRF5BCc8wKs1vq5qT3UkMq50
Y0B2Rkccamz514PuEsW5rgqKWkWxkaA8aaQn4lknYS/Ea1GDR7uCJwsiwL55l6sc
j6Th2erizdOJ+Wt4KN3i0CgG7Iz75IazEQKMWZ+9gbBOjEAd9oio1i7bniZQ+lhw
bmDVb2UNgW63k6AuEJGbM4VeJdTiwHpUquEbjMe38veeAiytwIvS7HnyTnDIAizU
2ACcYRE6dlfuovnvoyGaAwjZf/mqLl1eFKewf5Uf24yrGN5xA40z886sMFk0l/OP
Mwh1nNHraq7qlIHB5vSrjGQuwPf/6/6+u/MfFpCnQdH8Gw6XMkRb0AiOsSSm6M4Z
yLZV6291g92eIH+4kmZrb6ilYJDZslzy6ccTvkCzeEF0DRupVNZ+btytaa4paWiY
falgSaVG/9pD5r/I3r+BqbmDJ9wIP7GRFIKS9umE/xoX6Usi2SSdIoBS84w/u4eU
C6R4JeMGiIJMB8tv8mtd9VFCmZzAsiun8mfTV5ouXYOcFtsqZjH14aTBuDVxQwKm
GUTFR9snZGlLHv/p4q96Qa9Xp7tmDV5iGUkOalWJHJ3EGSWO+oE9ly22G3WTwrRG
ml5pQBiUOSo6VKrtmSRC269H2hSH2sDoLzTS/LqsVe6f+DBHF5LEJUKDtj4KT8C+
1LXADSRrHL6LVgjegunTAw+9Y2QmCEgTkrCGEEoq8TpryBchJHzePFHwOmDSFm1I
8rraEOKwTP8afs1UOPBIgqjXQSsY4H8k4egWgminfUt5CC2ll0Ss3fT7GHxVqdtB
s+yHNFds2nm13lyhrfgOBVAJ4Jv6wAPjk21C7DnzI6s29JdAN8ZcSEnc+w5ujeBe
xw0KbAcryI/8l41vjkycOz17MeHqWDln2VEMx7ePdzTQUHknszbEFYIdiqav78q3
ugmIXwKY+FUolahnDGMyk0SHu2vuleDOaSGZiV3YQo5RHgYuuPr7ZtjK3lHQfjhu
WnaamsyKEDVyi+4mj4ELoE5JIuqVz+EyVsOAyVTIhkBy3FgzcEOFBzzNZjz9S0zC
nOWXJf4uQRi0lmz7+L1oBbZXRoKkU1vHRUKkXfC3kmd4p4HRpEcO1wLIgNYxem0Y
hiEdAYVAgk1GswvOtRde7oQDwsub7FbobNJk1pSHR8HLptKJoIlNtxl/iweks0P3
Ws1o5KQL0TljC5BmUEYbdlT82KW6nQ1xO/aY/oYPmIrE0lRKU+vazG2iQIzTVIbY
oizfZDe9tctRYFOWpIu3Pg5KfYH65rStkZbGSdApAs8gT1h1+NuW5a0cg5YbKUua
DV/FG6e+SZxlnVeUS5PQauAnVxQJakKOp1VkW2Zn/IB+OL1xOkD/xmcGe+kn0Axg
CrfKiqaBMNYX3q93cwuL9WVvoSpfBsQyTqVABePKWetXBG5vqWyOR/kqptiB7nko
XrOFiSCHJk5D0VYrqO4aguS1gXKCBlYPFz7jQV3/X1FAkYuLd8vQO9KvIOK4Fd1c
VIfW4HmXiUQj9npClwD+MxOHyvINW/WEVih68B0mpETItLSWvq680UikmSWQ8UEe
I37KdCLUaMmwOKeDSIw2avlzqrrdaV2s2q/rZx/N4C0O6mI/d5HrAE39efFGGiYL
0R8qSv+DluTyk7ReI6zx2BRUB1lHuEkzxPfW8kIPaGAUktMaXY4FyEUnpRr8hOqH
9mssJ1i0mN4pRkp9mLSXRzsEgOzEa3ucX2qb8jcklu2nBL25UPZvJgnP87tcODQo
5OGOKHpIFXmHv/h+I7LmSkbC7TtyHaneUwfKvspsjQf/uyy0x7avLwVn+NEWHoHV
lzRWNW9h15morubos71aiMhmLCIRLryoziqpRISVAKxoyXuhiKTqd8x06zkNVuMW
ue+Sn/JcqWiyEa4Ijw+/xZKO4VFnckXMJXz9ClsyyRKyqosfT97cpwesxvPZIVfx
K8GiEbEM/nrRVyYk+FfcT7mBU6KfGSG3Ukyc0w2mqiT8QxkZxjDwpaEKdOFQVJV4
D6kNrQLS/x5DleyDhZNEOr5PMM16WT+dEYboFVTC1bDsFAW0c8ey378C3bWbJOMD
6AwmDnrPRb7ejdT01zSHBNbGkvbzVK9zIA4gf2A17ExM5N+5g54npLr6mbekaDkG
mYJ1WlPFWZCTULOhts5tnNVOk2ZR7v6lqIDsbJMcyB1fxqgw0ZED8JaiOJM63pVp
gXun2JfErUEsGqeNcoMcFbfQQ398O7wMqDNDz/XO+RrecQcoqC2y7g5+yuLZS7cm
JHQqmNw4/cR83ulv05GS16Ssl+kCmGSMR40X36HfzbEgnCvSMLn2hUJzq+Q54i7Q
SViD9Ro+NZteeHqokCept6PleDRnoGE5R74J5N1LiSfHXQXpdgeH/x1cAJzBzFxB
ZR5ukAg72ydWX+CmkOUQegOAQ8IornlYE6e2VsITUVtmTIMDTXoeFCvH8c30CX0a
cWgDLp5+4x6n9dnGK00kiwokKvpHnGRvD7q91zqsYxa8tKmglyqElviq+y4plhXa
1NydjE7XaT15IzdThuZ/VNPlQ38Q1Er59vlp/zcDrAZmY3JpGem40eNvB5caiqbj
FCIPbubkW4knBUJwatwaqt4XqkVuW2J7p6X7SfgFHYD/b/fRin8lHK04s8UGkqMn
v79SCgR/q0bTZhLQOm8D45pG/SgGQvGoednL+zYvI6GWGKifpP+RYbDbez9pD4IQ
EPQyaM1jXHyRPgE3O9U2yyp1M/G5ACgFXo/DuWoIxUudBB5uXUPzIS6becFbHkGZ
lAkSMawGmPx6kjACMk7YE6P5EX2P8wO8P+9MJvHbq2/TxFgxFkyMdzL7glgN2KiF
OVRR2iKTwdwUszjan3VcEqXPf4AMcEMeGh+RdfToUoMtMfijo4hsX2mVm18dD5h9
tHoDAiFenJaa6Ey039zlfYuODeEoQ2niIbBOsw7IL/gnFlPUBbmns+cXqDYPe48g
dE/kNDBcpbSGedW33Bp+yymFU03XbHNh0UBxHAJdzkCpt/B/lwEFFXggUZQFVprN
iV3hh0tYRgDO7Jl2XTaqfgjxTANP9ARhk8KRUtTbI5vF0di5HJhBX8rb5vgMB38f
L8/GJzsCLOi8+aq2iMA4LMqDUUMakrHHJoXJuXVfsiP3A8JgNuF/dB3xF6O9TpGI
kI+KclpZ7lXbrE134YpMF6QS3gxrlFJ9g1ncvytg0qYbr6BxO99RedmIcYJ9gsHI
/UnU4Qv88gBnpPBrScjLKcSzigtILsE4yYpLF7xaQ1r2M5JPOteYpOdSAddRWFRI
eDGBy3xsNV11AlvqIv/98rda0vGajg7EtRaPThTCUhJOsnc2J9xW7v5chWxmts8q
3rCFQdIouyB9VXTYseC5c94/pOtHl+XVByp03JqEyTPK5rL5EDGsMJTv7ulbOyjY
1s+mpJq/GyuRklL48qLVxPi8ov3JBE00HuDAAqTrIuP/5u8+/xb4bDNpEPGruVob
PJnk3tqAcSvSI3pNcIVuo1LY++kKQDRAGycY6RHyi0oAv34FvPX7PwVZ7vnfnk3v
IdZjqFlpITAeeJoNbB6g3UyretSZPmeHrkKw7axFR/zZw27tEXwhEiXQv9hiIgXV
eiQIn+6b6Mxm6JpPqQuywoHak2ZFqzx8JUW7PE6tii2VjvhelTqY0pA6lIZXfelY
AEp1eVJGnYOkQb1XQKBg7CuNNOqREkooQ60NThacQIiBbDIgLBl3ytYGK41TbCDM
7l03M+mjk6c0hiM/EXfm2ebyFleGPc10jOPH57NLZaR1bk3ENVLLQU5xT5rxHNeC
GcYL9y+aCrABukOu3XZgeJOY3H3Wtd+8mD7rCFRypuGWtH3JtbeIL1RE+ZzpXoQ5
emGBqjym2dN0CID/HhKbm9ws3zcFKFuTr1tufdzV5zOcR+lfatRwAxhBLXzemAyz
EciOAKS2hkrl9qJTkPeNWwKZWDgVpwJj+Q9aVeJDOJJQxRBs7Lrp0HMswH8w7f1D
3fJ3L9bXWqL/UHIAt0ooSzBhOlA1uwdIJCOYiGkgsNSag10H+ZIx3vc2X5U7cLBH
HTsAG7kUtyXz/K+4/r+miwB3L93HAi+NtbYlSZd0TMiP7D48ky0Z5US5O8OwQuvr
hsu/J0aQSIw+nfGTW7M1KSzZ513aVEUffU3veH9yO8/inLITrmOMQhWkZBwmsQom
WYXAgvqDB8N8RPfEpihwmRGHF6lQyhPMWKQDUSyWIZo3yV+IGdlJ/87BO2Xf+KHy
DHD1WjINNL8WWeOCuZVKB6vOGgsVnderpjCwudiIq7IpD7v4R7i/wvOpY3X6L0wf
ht01T5VUyvBIzIuolq5OkoIYWhyjqfvyiJNQQbuFJ9KF6/PqnkMayhB4XsRfGPOn
H2E3SaikyRqiRiTKioCYRHyOJMo5IvVsjoa0QXLuBgb1CaVigy74cDUA/fvUU0M7
iQ4qksevP7JafxPMR7diP0cpKd/cj/M+f8huTYIh/iCesC+ZId/eixQcSrB3Y4kw
gRZxRyzKLFJcbor/gCWPTq8ADSO4GhGLDVXMXUNsDWjWqrSH2+6zhQWdVmxcQUAJ
t9jiathVjIq29neF+S/vDElcouNvSoy+izr3Xd6xm3Z1cTVqKqCnVjobhM37jXID
7Se0M131EhoCklJqpovYeRk+tDTRmL0wS/KSUVZfb5Fw5JlyGSCYsw8rcsKL6XYa
JQ8WsjLaPCcxD3nZmhfpNPjI4q0R8U2D2Iac4l0erUMMzGs0Lhh3xkb2dNuR5RQm
D5HQuKSaOtGli+JiTrgda8IhnffRcAzF9kjzDR0T9GOm1MUaS/0+FMkdGml20wRJ
p9y54GIG5x1K5jAP3jg5HH+qCS5rF62YvkXEx1sIf6xnvYZUYQekvOEg147Glnrh
a1Ga8vgusWjcW238CckmKidk9Y9sB2i1o0qv0bFtUJv1eOJCcTNfQwQwVYk6v+33
n5FbcJgwdqZUGiKnZ7iJPaIMTimdWYeA+CbWGXPlIgSe16Ly+bZlbZrO9YSbNZGC
gZ+Xf2NwnYIGZF3IoHAWq2v6mD83m+DMmNxUz3LZDXRCaErDVEmPlYuWKQXiNnP9
Go18EoAbzaAhIbFWSmEYUxa20pz9TH4MCCX0Tl4H3DI1KuV6gdu7+mpWLyqVN6rt
kNgHgDd31yX4G0kiyhtr7oMZ08SP7Y/9DypJkQF1yAbYCs6iEEtvQo8Nfpnk4uXr
OcHy8b05wNezD27A6a45/sIdTt11EBXovCmTCF7GacoFbJAkv/McREb2I6ozKrj/
aOAitfXdvfCyst08ZzqIBT6Q3OlwQz7n7aOewRbW9BDa6/vUezG1yP+sAbPNcaEe
CTE3O1AQjTGy7yMJcMLuRK7iYmAQvGY0FVP5ZHNifAC+QTzoeXjCFiClPzKXFUZU
2tk+waWE3nQjg1BS6/uLdkGWm/IhGvvEsjaIxDk+44ut7dAs/952BsJCoRMWggEU
iBBNnHX7rei9f230onZHzkXP9RZ/xcFdPZ7OdJyxmSLHZ0SwqxK5/hkZe2t9kHTz
VrZYEAlV14XQHJvdoSfXg/CuPV9cCMP0QLBEL4BktcGEFECRiV/XHTyOO2mDVr73
9VoKOqmwmycC9O8cBCapKUQzAckJKYuwCfQgMtrHssOxIO9GHaA9Rjc/r03PXWfp
2wsdWEM6TmhhXgSYo6B8AUwF2bcCdFhKMvQRsN8Uhomnd4rpVX7LOzhK4OWrvUcW
BuKCGE/OPdPfzxToi+HCKDm+CePoaptYbqPJh8WMbeNXg260k98vu/Tk936VkNVQ
zFTHxUUGjs/MZ8ysC5auCj2iC7qvGz9Y8gWvYdKYzi0VXEzCd26/ucxSANRJwa4D
3n+famQJmhVAN7y5xdBdIhaJeYB5HQ8f4RGwMrChAXLbROOZVQmWO0Q8Epz6dhmE
Ye2io0NPcQJJ3oqoU8lDjtZYolS4KytjAtwBQhSbMBm6VU5121+NuakkiuOTeSam
/FrLSJCpIkKU0xojRWM+7UQxlbPfABKqc1BVmaiDIBsPx74c2ztk4Rz/OtKNHx5m
+JqcTb+o28QXm/VM+x3jKIr+tjfRMXOOwL3DblDJcAlMrxn1FIb/Mkfq5Vk/jPl3
8Tc/pGNFUV0/bqkVksp5Q2i7rPwIDcuu8KDe4S5fqYMhJ8ltfN920kSe5zajs7JL
td5RuowKj/vDICM1gOyjMdXqSGxO7wpmAHEqoDZ2N0arVlUDljV/zuA8n7cqzdSO
bGtZNeVUXeVygYvBpP0Kj1VKnu8+Y8pCVy0rW7LMOLPHDErYwEIStM1d6ZvG03Is
5iLrNracR7BilGsv3KxQldjOrhBYdS8qN9B8hIj0ZkSpGYsA/uH6FnNMclZCKslu
n2tGC1vsmb4/E+qJ3bjfyUCnxhQR/Nf8XoIYJv/dzh4L7RQkin45MhhFu7GH0cFI
M4tUA3oUvF7OlfQt25kTARK+xErMYu9zRrI7ff/LZ3ozNmLMxS+RoeG5KbtnT8B8
mbnuilRT3gS5IYJZ0dRmQlLkCIUcMz3KovQJfX18W24KDlxbgKRYF7k26nnBz0b1
5RxPQfFv7aEIzAFNUjeejua/122gwgHyedM57+9sHjwMtOMdmJQvSya426qygMgh
qrmYhwelS2tUkGs9IuZqRE/P1cdUh1IAB5r0GqW0NZpHM5W7476k9GZc1PiYkRFR
e3hux+dLgwmkmrKvbDoMcBRP+SdqtYBXwYlQnlncvJRxPGsSgNVfy3dEUheDpotT
rV+ND4nwepcgJIqxPAOEB6vH5lMw6X6xILzpIiavMwCIP1w55hBM55kKTjoFXi4s
ObgSz4jchSDBwQv7QDZ0vzR2Bo+/f60ozjczm9fTUFbqvsYarRa30/U4gxz8j0ec
zL6qyPM5AvFoLEXWPa59AHak9MaSFAuWMx5+C4fXNYkSPi5Tuq68os61+/KLZbGz
34saNvcH+lvWHG1Hr5342S9pKaO4vQWDLRFQ6LFTjEuNXwRjQRkBn3eIGg3qtIAF
gwzJkrVeOPJ8Kw/PYwMy5EytMMW+MfnKin2NT1meN3ELyyHcVt3CtFcnJJeUphej
tgIcmb48pvHyY5J0+PkOSYxnE67RK84SjfgWcWP4WD5x/IelYYRHoI1uNxsVfiZM
Gx2ksFfuI3tVrX9mwXtP1CXOyM2dAiLp2nCNwECCxvy9X0SGo7/HFKtamI5U4Tmq
qdBkGOAFOkGGbUZVgtoVCNYLheqe8KxPIkzlq7pDz5peQRrA3ej6vNGJxvmt+GdA
Je2BpieK0zkFv001sV6Cb1BJusnHJCZhhLhjoCts7JFlmkmP2YLTdRZruGiNEqXb
jW0HordJInwhZbHHIn3EQz199b4QoJ15X4cJjWLVyUKP4DuJjcTQieKFErDSOF6Z
KlzpdgTiUawrd0oIo9VIPMeNvc3YtfAguTN+VXXRtFcy5fCR2Q1FQgRLmc7831aL
KJ8qCR7VLL3x5H3C62cg/LZg9USSBPkRufrfFkD+9dqqSeNvkKw/QkbwghNQmWPw
1GJIWEAxisBKqYDH7JLiBFKT9lcT6h0vs7PoErfBZgZsGHUPSPpeD3FWgeejmSVK
Ay9Bm1A9zbl8QKNAp+Ma1unrq9+jQ9HNX5LZbAwxvH9PxU2+vxN51ffkEwtEq4O6
3kAy+OiHS+mfLOv07uDXXxm6EmoOzUJ7m63SPqUUC9kSddl5V/Q1tvZG4QSwjH50
IjAABbSg3pqqG/wiz7h3fyEg8LurvWtnirBGkkcAMg0WmXGYxfxa546IYXuKss/7
2xNz8CjjgUQNiXRUxNOqNx2uwIS30U3ta5kB7Gwc2iIR2Hk7Q7zRg544I6eYrpB/
mWKWvN6jUjO+/sTIlPcFI0ctl2d1+wkqvjABZ9z4lIOMdphJkpeX5MGFpxUYsQRm
mL63M66twvxfMq5tnQlWMhXNiIMijhQ9Lplf2OgJn6pqQ0cBLO2SDxCsAqXOlaFs
ij5El2hnunP8oFUU0A/Hc/zxvGeagOOdG3Me9r7V4q/8tpdXhD+Dt8a1PKJW4d9/
nyrilfLZZ5KwYN+zGH4tgClieguvjLqiK1ecFhjn1CxqTttts/EPtUuIbxCOLj/j
HS87iLh/6AxmdnC/DmxTE6lEhIidI/wj00frLUScecXTVDIsQME25Gysl6F1KnRV
25J/jhcKFwA4g6cH2DsZgkeNaB2bK+7HkwFffN5kpktvWHdqm5u6kxXiMInQlAuS
Dz3zki/gfZYcUQd3WBRfiL+JRkHihVHqXQ0oiVf7Pdw6m1yFMwRC8isY4kzxiROl
oTOK86Bh+6oKa0tAwTKt4E8x05znOL3jwRKgRYVe+6gEy8HG3L/LyefkL6BJ3drV
ThXnKUGiwzbMKwMgCVPXynPT0l3+2mPU8+rysqJb9fNxGxf6yXLVHf+q0mvcrM2n
BdJ2j5Ql4261QFjHmoQYOhd0zuEEMjDdrkioXvhZd8rHVEceiA70c7ZzxOOh2MZ7
W6KtnUh8CyODxKyjmj31Gg7jahikz+lQZVdvnX2SXMYg8IcDHV69+Ions57NuEim
Nvm+Xe/sVXO+obVVYoKCpe3qfCUoLySttHFme/gHZ3G7FG+1xv+5JBt6hT6luuMU
urU+2EscBpseJVZVGmtKGrYmSehUFy7LbXweN6gCFB4ehxa+TABASarbQG3UPbST
hafXbK6m/JrUKDE9jaXZQtZF+fRflXBkAUCU7W7LRa7Naf3ZY1YXhUMYK59wqeZG
UibAz4GBCT69vZGNuVNkx5gLJlJry9i30EECkByYlW4Xs7k13sz9WOYa/bn+wwLg
HaPtmSpwZPDzmjNAKCQi2OZglLncUZUImIm6Q2HzjmHWtnYbI3fictg9Zkj0hk0x
sYfJoOm8AkhK0h2J3ljd5wZ4SRi6cV5N3BBJogZv5kuYyLERI+LD0XRV8bWUWrMv
N2LyqnN/Tc2Y73RS2lTnD17M0ZM/Edre1gxuP52HyOtYxD0hF/MbCSl0X8g5/RuB
F0KpBKaYoOGX5mnIRBxci/4Ru1YnNl99B340nkvV0D1kfLxF9WuUTZ8LyhVF88OQ
OAt9qM1ah2gdh/a2N/DcEAeB6y7la5vmrRZFXtju0JZkAtvvVWE1Ss6PkrF3I+Bo
kZTbQi3npJk6m8KIjbhwq9++vVhz3ZTox4HoVSW5dlsJ2PbAqzQwvmCGpyMZVeGU
QgPx8zcw8ol9B4Qm/JD9+fYXyti3CWFiUNruAnD/uNTv6guGzkgK0uYjy6XQH3Z4
umcVrt0JXv+wi5D0iY/4ZooSeuzJftDwzQ/UhagH090HFi05gQfTaAcaiQWLpsso
Eez9HMcX0/584+0+52Up2hwG0rtL2VENilIbadh/g1AxzmEr30hz4b7UWXbG7grV
K+fc39lL8Z4+od4us5+kPGkbeIvtBB/ggsand+23Dd2UbS00SDq3A2ovP4IyAYjP
liTjaGs19UGMY06OEsHSTZpJpkY1qXvVo+/xTzONQHmQXnHFhgHOpBSl6ORiUGlL
7zape6YUrg02MP6X2Nvrjw5ImO/LT10j0o8dWaxR1HKK9bEIhoXgyhnRkSCwFAFD
tXUIvEomb5FHj9xoVcF4bPqU0JKLctAbWPua6xjZyxHT1wvZL0fVPCYqhiiQOuWx
FwLm415L7inpXSwME+d/hjwBnHhQ3yXvpbKCn27A24QhWdvPha5h9GDrJ/n0hlyX
VNy+ZAEr9HfTD6F8c3KCHjppEykUxqdAIG9bbXQlhLqIlMdNKIOHXFVHU0PKvxV0
3usMhbZ8ubxKjN+ZnGWi5Gp/mT89jolc3kMA958JMyzAh0a7fae7+9KSQ8fQ2Sj8
M70KJi5+rdt2480UGNQOskNurKZ+YJRmg+PTrdOnPf3p0A27r//u5uc7EcGYit3C
FuN/1gLxMz5U4ezqJgP0hKl4VC85o66rgT+bt7rlYOZjmju+kC9BjeqSlNTghu0b
/KhdJG09kWKWdQZP1VKeIJDJML8yb65YRnZR93BDjtjEPhWsD8wq0FVfgddWxeWm
CrsNcyxD9cTTG+DHPgX3MEoBLmQTgW3gDdyik0OTIjgPaMP3F+Ip+6CYNzxAaXPB
euy+Pt6APEHZ4h5HCzvFh4dwftwlnOxuD/TBDuuRn834S2lCOgHFG7xFQf4Cfp1E
9LnBS/YBBIOQRm4ou7B7qbxYpgL6VzAnte8zPLhFnqw0IJfS3K/83g31E2pWVG/9
ugoR7PiVa2O3M0eyD9H5jw8EGozkoQmQQ+mLnv1Zw7IQGgOxF3Lo4Mfx+7Md9Cdz
40poN+KUQDrjIK2UXzBSrIjjDCPXBkJHso4bBmp/uHGELvNTDSVbnlIwjQP1HOsP
0MdQX33ezLZalYLs7iz0V/bQ0oh9mz4mojlzC62Ix9Gz50mPSw5kiYzkPNoxHl54
hycGGXJ4iPhC1UuN8vszFblDv0d9mwWEyawpBAEyuVmPnMa+aTDI8Fh3cz/SSm/D
a5aeTa7WE/w2OsdH/OnrJWHWa+BGZWjrVLtTwPXjf7DckgaHJdGLZFXOdmXWADwP
Ys2GEhhBo8L+TocGW/8R+sBn/rLeQzN89asPxtTgTDQAPWhqSOhJdab2NBtsAohs
kBKjFNglJuKlPZR0yem+RN8dRx/z+L5q/0iqqUS4LjHXCSH/gIjQLUi1U4nnT+Ui
Iw1l3Hp98KjE4VzXx81bLvf3ulkvew9mwWbVZYn5VzAkQXbXUh8P/hme0mFlLSYV
F6AsY6Zslq3PjxpR9eV811yYdOOUz18VnYCZGq8ASBNDIquJFJ4BxvlSqm74Zx+V
qrhJ8VbjDeOSxdSERwewQTYCf0EBN9WJCFm7KKVH72SMkg1+XEGeXz44GdymCzGk
tAVTKsOTjZZ0W1OtkHrc+6GkaE9ioJYaNsRZK77xw6s99ZE+WDbMY81CV2s5JGHq
BF9nt9ZjBmBhCwlFyyZwT17WGskyRAZfzhinoz6jLLgLl/GfPhzEpaucipxDm2Ms
7LgpSkKddL8bPCpOCpSQZEcBYQJPyPkF9A0lkZIEfN8RNhR3vRCNeymnvP+0W71h
i+hbmT5fjFUDW58xeiDIMxGDOtY9M7pgPul36nkPx0l4V/qRkv4pdDQw7gG0NZDB
X7LjnYcdC9OJAbJQctGFu2mp2IFb6ctecpDq1LDV6SXbC495fMwmB4jHk9pEM90w
pdiLuGubPFKWn7UOGVDj63AoYfXb9bw5SzS7hgUeSPcKkC33JoIFd9y/mV43bVBA
h7es9+s7a8r6M7zRi35HbjuEXCg3ms9gLyLEIU4Gy3TvVOKaxqMKsMrLDFpmChea
ijZLj6YDXlYustXuHNzGqyh/WaG7WbXAKAB0o54+NuaSoNK5gDg6CuLcHjbysiZH
vaL02vp0aawEUqJBoj0auSZrJtjk/f+4tbLGi5vAvOTWI84osxiFxdBcgn9rBISt
t4bhjZxKu3w09fHDFGh1VCz0WN2piLmPON6WUAbLtDKA/PcD7UQdabnyQFGaCIt/
f87D3h+nmmxFf/vZhA3tQEm6RJS0TzU/icIpcZJT+X7BalY1ljIR307xbVmKrb83
4wfImMzgChsxMrjH1OEckQRaXsxIb8ce40c9IAUfCHlnNbPc+oYygoIbSL2BUNku
esiwcwwk4qsDlLhLAHJWecCe24OOhOYJTrB9bubMkzR0MccgYRdinCSQch8ZPeyg
EAXryv0Lr8HvVJulsqQ322ijlRCM/UzGVciNcc3tAfKsHoJ1BKdeAuTHASxGS2G4
QYp9WUqIpvVdb9RalmC9WHqX2xZfy5gP625eLpDV7bCLVQjYZYzh58Osd3pPVSkd
x4D+nFNmVrXemPnuMQht2ZG5J3ZGCoMDMQ3HntgyLTeCd+VYIbP1GSSkmvmD2iPU
86c3Ubvk4DtiGPklx88yRArSTZLWP3XFMhyNQxmmm+1uABESyWDy/cYcVyPF5EjF
OjG9iYuoBtTDEHFK/yvTK0jnqZkljmcYBVzB1/r2Os45Tdhor+O7M7W5bzxflgKB
m7RD42baQl0a531zFXBpyLWbJMlAeFn4O4CtUwqqf0FMjbxjeuzChSfNvek5BwbE
Lri7BhQ5KU/jaR2qWKaLgE5CWY1p8WrLOXkin8uAmCRrzfKznfHJASOvtTgCD/GS
zvIBl4pZGJqJ8elRIJ5PkhGvxvq2A3J8CRkV2DnfVbLyf+BErSLSptFxk343Sh0z
hO9VsQvtZXLZNNHLcF/GYtF9pm9PFuG49IMmrqk44eJWTtJ2tnxxESjhwEwvnfdl
2WD0FsaTlwKMj2XmNzrKtKprWgQaa1mNimZulQBJy4Ur7IzQ6QnlWXJgXXTudvLJ
dlo3+uNNwfmyWI7GT5qYFVCa75GuieHGFDPTKgRTJFrqVnfirHPWOU/nwHaAy/UA
tk7bkqX3738UAIbLiO84QB94ahKDuAAojXQ22tLTlzy7H8qQqVOUTWCYiSrXoRlt
5xmg55D/nJpuZw5Jbx9EPm1/+5N9yYsDkKeicmxrjxFzqZNjMXPGcnA0fuFdImr8
8g2xP2DkisdTlQCGCWDHQaQC8shw/l1MsLJ8epO0L5yrn5EoiL9q8jvy7P0woa9J
/wKXaNfOkNMTew/ngdPRhsrrxDtHa1lXyKHHTnwTcHkcm2mEi9C5C2+1Jo37BOcA
2nH9WJxrQA5gtzJzypKPdtwkcp5bGlbXnHosMKszWruDqnsaPlzYkC2Lf8+gxtrO
xoPZ0vbPdHtx8XMe0mkZPoDjRkzFdttlpIjEzfO//65lqWFXYswqcEIAV4KykIlm
zz/gHn+r9o6t45cXDO3RW41t7DxEVrM+J9Op2mWRKmHl3qCDjNVWSaWIMDOaw1xl
yPtUngS6XfvgZQR2L0BT+kLQTft69G04t82PGixgyUVRylxuBL+06B0bDDYmokE3
7mEpboHMC94eQlue73GwH+mdchpNxs6mlwsdRO9aBhqP7ylrNK+NiXqnnthElZE5
x/6eChUj91QdOND+iGl3OQdBHil8rIFWoqEzzqJe8Kwj37exPb5ZldSBOyuRajp2
VrvdlejKpWmwacHhR0L9CzNXZyqKj1BGaxMTQat8hhcZGQml50zeuPxrGGvTmcbN
pTNVCdWAknzQ5grnV2ffW73P+djRmf0ClYbsfTHfX2eIrB6w35sODjnwTL/Wizq1
5nQhFLw5SNc0F7+ix1Vymw04Fhoqy8F6R6dyZMC/NO6MBfdNfDH+to1+etlVc9ZW
YvHhdS/ymrh2o+zWi5jgNARuU93igwuqVdc6+r0wsSbFpaEiuXMPaBiER1s3vH7v
oKljev7+3869c0R/GsVEBVui19Qx2l6rUODSAsYhX/y7uCJvJJ/OIXa/BD0qF618
su8VUm/LdlOtHjdTDg63mfgWp1TuNLNl7X7NBrgsOyfO23bms0I1h7w4TgBSXOkj
`pragma protect end_protected
