// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
SbxHvBvCY3MTJdWdY0fO/C56yDmlhGu42Um1S+kMVTxAcG/jZ05Rg4irUwz52n1G/2djFQe4AtHY
wvyhF7PxqT0RGcDCNSUM15MB0oGA8FeMiHrLtosubie02NIoLRNL2XX8MUS28052QSkDNF6vyy/n
5aB/clRV+9KJnXEuCq1xsbMOkZZk326VZgNs+JTE3L9rAo6L+pHAFW1vlBU/g8p+i8PYA2Aw4IB+
nIYfIhMnLD/e5Qp31IUYlzoFOdBCdnjJKMB0Brrsyn3APV4EdlLlS3eMIXKAYf7ZVpuZKba/sGy7
phoeeghuHJbQm6KtC0kn7qRXo3hiSYCj5nikpg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
t8Z9pIZOYXYnbBm3DCQ1phE0GS721Fe2ABoI1C8nwH7PD1cP51QQnDrpoQn1l1msf9WrED1nxJqI
xcaZtPnlMLsUF5dfhDL/LXcKe61nZqy2DZKIQBd46m/ARve18QNRwJzbqzbkBN8B+XDCgfH4ztzs
AZsYjZMAUEC5gP2qvWICWbX3Yp17WzN/s7P4z6239NdSKnDHeCxY1ofzw33u/MYzc7STqdBg/Klt
vtovhV51yf5SYlfzwXelZN6LZhAEL8H9php42LnrZINAfJCoHejonmwdRZjohBML8dZCWm4MfKQN
LeTCVDWmfkXySqR/xKkm+kefK0eeLHRNVXOCrBOqC809RjfU1ETJlFWYpnpt01A3Pq3XrGSpNLJ3
bXBCoDdmXOv8Qc8hU7mG+fWiw6hfvNA6CbhcNBHbVxJx7MoDowoIQ/S3OI9GitrjCLfNZ+Y4it5y
rRZBK1RgMp7ObvaOD4QKZEMKhRLvLtIk8HIlZA62nUQEUzU6D1l6P6gW9qXwxUPg7BDe7kn8pEBG
BHbWS1tMnThsv7sOCsHLHFgpZGNlBUdbz3wGGthblj9rcea8k9K3aX/EN9gv9+amQC8D8BY437ur
X5Q6RQLoglDS+JGxBenRWLrBH3WAemWU+T1c0Arxl4M2aBVmcsS2BfCzUr90SiFoqQCi6+aJoSig
BmyiITPetY4zy9/MKtv1qCx1ePkalwu0RPoOIsB+B9n2WGH+QwYN1SZhRWIEOfkRNoGdBPdE8Xut
Z03RqzNQ5eNuN9UG1usMPYNcX0hqv+Yz2eRjc12qrf0ZMXEl6Jk0ARzAaA+LnqKbh+ayTuVSLgWv
FSPsqq+uRhlDF7n77LOSM5GAbv9oFQ2gWrj5zjIyR/0BFiiaOJyIAJa4gG8GQ84lGMYVIEmKaOtk
saxZ6PxUXylw1Os6pTEjeLpZ3xY/cLDqPs1snvcFuRCGyQLzUSRLiD3IT8WGpLNrCfmZ49A/8TCZ
z2fJjNfXsL1TpvNLNsrLjv6CQphMXhMlUUnORCLmiLBJ9wk0nbxJBtVcG8p2d5iUIG70Qk6DmFm4
OpARKDGipG6sY3Bc3RuXynRmREjtsUz1Y+3YwRafNLo4sIRBlGyb2nLBZAnNKZaWbBKiYYBJC+MO
Nvj5boRn0ZUjwAGHua7yVzc4F5M0o3tbcKTwge+/PuytZI+FUYdBn6Tnymt2yaQvvvCzD3dWjPXq
Ul9W1D6p6C+D6pLkwAFbOSoyVWiBpGpg6zjkMW5QdjKqudMkQ6mUo0vRkUuxNaFSF+U8x1CF0upv
UcUfSAWhXAyKdOYvaE16yRN3MXYf4KRwfUJwJd5wBZx9olvHeBAbdpJXr/1txHUXlr99oH+C5vlQ
xPjb1bIP9CZE13XiQJ8Xcmx7ue4oiDi5ueJAWMkR1Ce4SNs3PRUbUQTspJ9xqPHDMCq+oxPfVfoO
9Q5IjlB45HBmdZSwRxm60bTGaFg6hcVVglNYLlvQAVFUMvKqleGS5g2nTsYSapDQa/8aIpPoHn/y
ia2TZ5t+hF0YyGgLZ4ni/TsjIQEZhQEt2p5JNp0FgV/BL94aFJiYDsflUf4LpBxk3H71ORyI3Ws5
w1UeqF9h5mKPZ+5tX60vLq7n/ltHiOSsUe72lkAPrhtg4A20ltJO+VtKvv0Q503EXMvrOqXuXN9p
g2J0mTki0NaT/5+YMJWY4rWUm0VhhVv+TrGMzRoQIFw+uAeV26PHec6OcCxZPM43Vv/2dWVSQXDq
QxaabvYty5kdHgAME3lqqwICJ+pNQ7XvmKqJrJDE/6SlXB84kQeje1YDXt5v30L7+HVWpNjYwtYi
4D6zlQpF83Tfnv8Z9d3tp896QhbpVKK9+qTpIlqivpUoZLod2VHUWkDsMK9JkpqANpycBUR0ITNb
gxpxAwrUW8vXQpG6kiUuvog3K/vhlX4dszKUE5Ze40b7TV2N23UZiNUK1qW6i8207TlCx/wtPHm6
ewZKGn03zvp66TW3OehGtGtVz+K1PhSShG/wrI/qDbymtDHdfaBeSNh3WOJqYQb7Ec4MyfAMFENB
AofZVgo6/P7anOBggRhwFWockWFbZJT+lVyll7uLWFFkZSRKLtVQRx9oCWWDdpfp95jwtH3AnK+x
PMzmugADvn+0Aw1vhOknrEuXeicDr82qcx0SWnWs2j54LSOCXBWpFei8d8HtFG5StysL1lLMIfM/
SPQtQJtTAuyvyvKCsTQHshV7znlJy6gZW06MlzPcOVzQHjJhKYjZ7lWee+zC7EgUgYMelqLgC7rf
WQdgAq8ErUELgaO3eXc2S31f7j/qoZefyQvSBkAaS9tbnU7crCATtcLjVW0K6mpih0BXiHAmuLUZ
g8bPzmImfL/dg/uvAWdYDUaGVUfO9Az/feuYNV2zwW5TxkBiI2/4kiQ2YyD4DiG155FJZEkpUY+c
XiVbrw+gYSdyRoHxOLEVy+w7/Me4MMY2XOhnozvou5obKqx4So35MDrNOYzNXtlBi9mLLSOm33ax
55T3QYyBcKqLg+PyFSSiSw8I1052P/R0z9YT136rudtIhW7vHBgyR9H0xO7LuAMMtXSpHaGq1qZZ
Ot+Lwd8rpQuPb0fffKGgA7eYYzpyhnn5R9lwlV6oZljjeRY7BlCuRaBopSDM7Qh9Jaj/0/dF5j/v
3CmOcG9sw/SmnIn7O0SuSqB1a6bgi3IlLLUrPmw9+874yVB7KT1PA09OlT0s8Cb2jjYcU1ohkj0j
lGiYu2tG49DlHif7qw0Ch5jrFym1c+xsJO1uGcrKVuJuyUAAhXk3Y+B431jROAkcN3wo/aJ+D99o
26j5Q5LB2+pA3Cl7jQ51Kmtvwhjm4h6K2gUssz6euLH4Hk+jr2/I/WfIFyZ6BtcDscKcXhvVN3YT
EHFLL6jBRPh4rTYFo9eYWl4Uy0l8fSZrocB59Crtgg1o/IUlOemJV8qRieY3xAQLnnQtzMZskGNg
DQCSvtIi3NUcaoeVi2zUlYtW0tQIyMsdWFDLClEoWA4P0l04q6gonMjL9CvBaFyhYoyaqdUficNj
lEDoY1jnOIYZHbZauNWWTsOa0rZkT8ogxBrCMhZa4F46j6MuPQOyAA11WxFomRrzWd2Sb5g3rlUY
W4yCAMt4tBEjD8VhPmOvRw0hZTSs+vlmnJcxgQUj3yn4czcyGkxvaHn/2BQHy4l78WeKsmkl7L2C
MVQy4FE/0pJl5dSLlL7/GVCIro/TvwTcBH8zcey9cvUnHedA3N/AkITmwBmVKp05PMv7oK43n9mj
+6K2+gH8CjWIphBlwlAdw75Sl6/nEZPmNJ02oqvXDAup+8wYZ+wAKHnuXZN6hl7XUnKvPAgs91SX
B7iw+bdU7OGa7o7RYUJLGJBbqklO2y0wFluZQC8QF1UdHb4DyF3K95tSZULjjUSWgSDmtsIL0IGc
jY6hek63EGWu0c4CXBm90fUSZjAo6emJDFE0EzTCiXjukudO+GsVtcqkX1FVdwMK/tQV+4BQmRFu
AfFHkyfWueX1xQqqtHFMmytwM8f9BRSU5aOttAqwVR4xiQayEK+JiixxqKNyBFbxBaKjL2dX83dp
4/fGQmEdQCGzq4ZRG3hkSwobHU0uoCOu27b1tlmygN+WasEE4YYBGIcjt5jgAisackELkDklyTJv
EjjL+6zHKJtek4WQ96WxeyCrVirxN+gq1/w5XzmiTqJXq1gDV/rvmRmrS7OBTgDoEfbdD491YRyo
gYuPu3iuqZYueIYtgYYsv1A6QGfNj/UVAitFiGCmdWWDHsMHJjG+258Ps38ZpT/oXqAeH3e8KL37
tpmlMTzuu4esFZwXV+m4g7ySJXbZ48vhGzRCjAxY/eRhS11MqJ3JUGGhr0dHrxAFdlFxeWwjHiGr
ZI7cmQHhudYFst6mF/BWSzd/ZSG9Jz98sT12QwStf3vnA5Cb9nY0iqVkixbEIHvNk3CIm3epvby3
hPdf/sy6ddUH/SxZZEwVsAry/j7MGeYzwh9MRTacIyQkAxCV4qGrVzkNJejlw7sgl8k1paskyQzN
7cYlU+N8NkQ6bcHHRzMUEKsZq0frz09+RXitb+fIdxRWjlpF22LTlzRjaL68i3cKM26xw+tK7RG6
m39meiD2tQRkkgcXIoQDH2gAsaBX9NBHLDfbDC3his8eg4LMos/4kOmeHHhyL17+loH8r/RouMLX
/z3lWF12TbCW+nUSrnqmWdTW76Jnj/WhQ9dL29sjUEJXTPsDrEmidGdu3AXINUlSAFvC+z6E2uox
ml4fsSJNasuy0Jxb0mdSPbbidSnoqffn2yazpsI1QwRCaRGpS8i4Pm3MZM7yl3GLLdFgx2rVaizl
RShlBCjlarLbO4AaKVLIh7N26KjNqFpkjWlpx1KeJgtyNsH5aZZM/1Jtas6UV8ov33s44ImjvmJa
3le3TCCyoCOWJYKn2WgVeMv7WZ154IfB42CnrSeV6FQMlgfSUhryDeLOPfDIVSneSdBzVOQpb7Db
EYijGpf8G5SJfhS+bpbc5CRoKLirGe/WL/IhEoeILgX8UJA/cRK6I66F1NOEhevr6NIZQsacdQPU
cu4eqpyVK3l7lvFjFpvq/FI4lyKLFWKT45aAryQ9OL1SxHbxEwRTd8/XTzxsYhAt7aFvMdxXhw8J
FrMI2ArCVUCWdkNzl8aAhuqmGBxrIFkoOMjo8A6BvODPIBRbPuU96muOFsG1y/99Qn/4c14Ku7GS
pF1usm9aFas5Ai3p+tT75JGB9Z5tk3XI0k+DVfwBE4Gl38xHAbQzeyJ+m5BaRiVjzN/X3swlEWtt
fUbUHWM++HigUyVVHvw5pE8D5p8AwY6CSPjdvjOOM45QrNVvt6BiMZzHQ0hNvxeo99eySd5/cDjp
wsN3AZDQHR8c1XaQHAnRKVFRTKBIDoBdTFqQAAXwMVEsv21hB7v8nYQ0v1MrIhzfkLvMwAmNK63Z
mKRSO1ZAYqdljbjo9o1sx1i6KlNYz8O2D5JVj80JrhHYir9qiBHnoNgkb7nl7j+02JZ25V8LbdQx
72lYrZ2tEdBw30HFO7aeTPKCm0h52PkMlGKf+t2+gONo+8b8BXOeCZPn9a/M1sE5slKhuwX4Ol4o
fYkHe4YkCkO/8p8YXDjs3F3xfgTLWlsTU2K/puzCKp7Gwvy+IgVBK0Vqmak1PAEV04t8dMtPAsxl
5zNl1GV/CSqQX8tVzvZU1R1StOymZ1rHFscEIvVSbemnu/tFyvDvJBOz0LfgxCANdPHnlF0KYFhm
dH2tYPCxNB48mmXtfumM0LYjCLdZMQc67/bCDhxjsXPKpJcMS64YyZu2I1IiPJJlK0OUDFwfwxrO
Vr2T9A4ZGbAqfOUHrfxKR97ivH+MVIsXfp9cMwUBOmkfj3Tz4LxTDxqiGWFF4YPRtb2OR+Bq+jq0
VJXLMzhrWtvF5kfVFNoFQ1UlYXfr09gzQNYraXd1YyaR/zQzOOuhAgRD06ToU5oyVcnukrDFMjPM
pcm5N4mxVNyaz8WJY7ZujtIaa8qnKNdTpS+E9Ci1Rhx8Q1/sqRYw6AsWYnIl7B9bA5OvzHjCWFzM
1Qrq/+xkgTRl1Gd3IwNVA7ScK9bsUHJWWeArQ1cGcOVW8ovQo7lv2Y+H6ClkuZlkn3D7kPx9doaK
3+JzyHMk1XPwRoWS2fj+C/fe41xsnBB+h/ixpChtQyPqeVSgRWdS5PkJeFVDuJ9yWmGqD20a+0fR
5Sx7viaPe3Y1ePCOn1UvYvrSOd7SQBpBbAekNkT3/6t/2hTJR3iNrNWGJcWlzq2LvO7YZalfkHWt
fjE8c/Q/MAl83Va9K5Uq+5KxR0PwnNX4h2vzWNnhTlCK0VJEnDbFyEKIC5liKjPEFpFwINpkEmLh
WGyIF9/mSmSFQkV2BTdkhGe24vAE7DZY0LkxOHqTXuUnOe3FMLW2ASmOYCV70e90fhJtvHLI+wN8
s+S2vX2c3L+3HoIEhRtHE+7ccYCE9avhH08H52SU0dkBxWft/mSUHSchLlOH/DTsgthfky4d64QB
TJJek98q2kElk0MA+Ol5NdhigNii1Skj+3QhpkARAHMMXSrE2kUPp3uZgvoy26bRGbA6f1ghkzXZ
/asTDvMLFgkWFwrV9/jgcE0zQITiRnqog8ArVFE24M5lTfPDkztCJEBjfBEztCIccKYABlK3V65D
rzfi2gVAKle1vRqt7lnZhb+s8uqXm5jl74akkzRU5RGhANrQTg0v2UTHo0bhsXlWi0z5ntnO0+Lm
jWcHkZLMJC5D+W9BW6wL334LtQnLqp/la7HchvWv6gqu5+o5J/Sv/vRdNSzEXrFbEy9fFXASbDQz
aVk31PWijvL6NFqPXhLtoqnQga3q+8M1wdX9MEc8bXTomxu7m71eDCJGpwLezjZB6SgsQPBF8IlL
hrRCbgphjOWVhgBGvC7MPW8K2mlkz70nMsxGG1QxQM2te866ZLwLaQuCKIrHu6uBoY6cpi1YyUqZ
UyLv4JLNdk3DPVsQ1oZz22ZTW1yF0CfzE4P/jzaQ8i5BxYBZR/JEBIAHaWAfsXziWK6uhIakuHFY
o7BcqEysviX2wAKQmFkbBTRFQLd6amDAgG+7ciWEpY3Q0Qq4KQlhbQGIiSpGEewHggVrt8kXRB4T
tk7WVKa7pDMxcQ1rSnwS6xJ3hVbtpt8YnbQmDZoC6pCVxXPNfv8uTeqSUGxDGcQnBY00hmy8kFFu
5Lfia7UaiRcHaDyxqCgh68FTwRrHtzuWnowCIK6X4Zb5OkV8BQ9JtmYSh7oycpOJ6VeozGWuQ1+I
/lFMJ4ddPBW6F4APzQinYeNxSda0+dg+I9ixSQmUt16ekHDG/duBiftAlJABDyz9HYjLVLg1YSUS
Zz2iBjaa1bgN5OT/91MFpeglLPyGYeg324vjiIRnihazmhVt6M015B79QraJgGmrnFSv+lvDn46e
7+WmLVzndiKk4792z31/S74zUud4oZQY/Qv7IpXSCr2G3X70iH3vPPlZYR+2L6PH+fQNuyZVTQq/
HZH8pknrdDkr5wcUXziZBxqbx06R88WWyIhb7eXS4KgvTV42+9LapHVpSWTBfDWU4gbZaFfsu3QA
9syXsBX/H75TcNTktx7jxR3I6MfV9wJyUKXzVvryvSSeXvBZT1oofyH2JrqmXCOgiZ0+2DjEq7L+
pePdC0LjHHMkweuHupMtJ+aVFPrEyUEqLzohZvM0+QzR70XYcvp9Tx3TzdlYL24wX+KiacJnYlDC
XiVZ7tmyX2xJQPOGLCsg94vfBSWl8Uug0MA2EftQHVMkHMkOqHW8iZJQMERy1O47ddhJ8sTZnbxZ
B/JYYm8MsXgOrt6RFDDh1LFvjAtVpaZ6t6Y1Eru9feq2MHhBRCuQ13LmCmH2STkFRfeuT5KVBw/P
TslHtYsTD8gNj4TD38ZuU7peyoDgsFkc/h00a+dTYlwkVoeYwz6jf+25iP+3I0u0SupVXa+W2wNz
fmzczsRIKQ0ZpT0JC/oKpcl5HUxIjrrPJn2s831FmyhKexPUuvfbmpu0YcsDYnscX+II6Rd610DX
gKG0UNqGZ78JPRehrhz1Py+uvYGIOpVXoPDnaJHId8LbsbmR2ouM2iTZT2setcAcEe+uAnvATTTV
0Vx/uIV5UQJ34SpxHMXM7K9x0wz0lAXKcl2gOe15skkxaDyihtRf8rDxMlXm3Iq6vSuUqpf+Nj/6
jMR84ysX+GpWoeWHS7kDGnfUDvPc2M8POAE3HdJvM/moxiN64C3jju/ct1v1VVjOZg7gmrTKXM5r
6D9hEpqxuhcLhxxa1MoMjH2oBLg6oi8yUnN8KOaS2hpmr2QChFFKp4r/iCLT2YHq3vUZG7/v9E+l
SFfGjY4yubM8yciEsxTDIhYzVQyq/xhT0SsJIy/5zD+c52fLOHzl9ycs84eQwLh9BAKkpYXHsxY8
5fRJKM/qaHqqV2PQ9hQvJ1qZYb6iCHorbcGx6mwqx2hoHU2Q6OA/cSQgT5xgrBLedwerzDkScWoM
fmP5TO7To6/mMd0GCoT08SgiOuoVKdw9fKnmUJTNRa8vyLbiH5lWaID2kZCOXc68FTt6FH8LuDIb
q5HE2Xi1ifV+GMWjqG0pdtjzwmPUy2myQvN5tCZJkUApkPerU3k/bPu9RRHyu2bfNJ+0WwvELIV1
oU5nWqjN0q1hsigpD7owQCYlgaCLT2a+X8Nao9dbs4BLBcI3RvOTG1B86SxeuKOSqeH4yN1QClDh
zjpORUu3xO/+3vg+jI3oDH1C1b4NnCUALVkvJt15llcyUEf7IgpEzY2Z+eYFEELwvmFwqatm+9L+
Gqktai/TJp97HyNYL+sjWVEMUh1Ss0CJhxy9UE27fMdFBtwXf+J1076z2AHZNJZqXIGKjZv/kHzy
0qOpE+5Aeup2zplVCVcUfUUzmnjA2eI217uM3BOYj9wsvmbBCTAHCm7ecv3iceiTJO0ytuUwC0Nf
IzruSbfmN2ZjEkb8JYn9BtceVWW7IfywbTMQ+PGFMIzQac88SGNkqTFO8gZQ9XlfJ2cXNnSpVihU
l1m/LiYkK04h9Ak15GqXjLX6JWzn4wxp5UPcJ7cWE55uDgUnyxNaDj/iKwcSp+EcwV3Mbz9pwRuE
vp7JCwEB3ye7aGoHzWokpj7uIvQHJtual3wbmPa1aDij2/JIzqj8d7qQOkKgJHZBxBcW95YPt76e
+kzixBi9JPnFfRPF+dlSoBWc01slyoaodo9a4OIPjAW+o0dzq0H8nTur/nqRq41SVGMJf+X4aK7g
atfNk0AK9HF6omKvetPDYza0GlrXZsh+GAKh6/YyQwElbqe7vCz/iDviH+8fCUA8Oo1/F1FGTrtj
jWbQFyq0/y19yZsrjxy8nrthzIv2YH4FHdohEsFqmtvEColRjM4JNeDMAf0gQz/iOH7RDVQmUJBn
8Ke4riBtzgBCP80U7nj2YMedH7NPn7P9D2/Hnt1+4dvrIeClUufb5wyAbAiQwDCTqHqaZYGNmaxy
Vp4adXg/NWB4CXRLKS58f55hOCfO8EU46VNxFWLb52Rk8hDJAeXakw5V7/q+vErjP7uiX0ymtOgR
yhvO/sThYD0okEpMHY8oIixNJAf8J2DExD0EOlDb4/lpDV5avR83ymkP697bkD8GSCudAJdsm0A6
5QN8qVRL/poEob6uTzJQXaLeIVkQXFlIUe7PHO6d1225znF5gwUHpnWzIqyarSoaM/5hmU0P9rHq
81obTMYF4K4nT5w+uxi1Iz2mL1pFFHEWVhuokNfC9Q10t/Y0u2l4OP4sNRp1MyoGddplV9X00/eg
ZI7J96Q1Q3w+uwXCTBYQ0oUU/FLAaswcJFWVDxjlPYVq7MVhFSptaBBsX24ttZwxkYozQCRQlRsS
duc0iI65NBf5E0WU1GTTPGVkhQEW0B4JS3D8dzHEJIA+AX7cHR1sIeLAHq05IDinnPLnmA/kx/mj
Pae7Ld4b1Y/wocMxBZDx3h/Nftvq6VEBCvoJxK4/cZZqAkYjGbhcHxunVlKucQAg89fJtmdFgA1p
HjjJtnmmLcZFEb6WIfdQ1AiU20FyobJB3KRPqMSABzUFw2Be/YmwzPtpD+5pyyGD54VIOzb/dna0
uvFurTbVEKMwWXE7h+e/jFPQoX8OBHagNTixfr8jIpCuNIEKFrKBbmdM9sRj5pvVj7luUdoH9ifd
2i+ku8g9Nt2eCwz9ATHghP+OZiH8l5H1IZyCQg4SE2wM/i7Q80wGrBhmbvNS76qjpxyxLpTMBzAI
pSzFYtLpuFt/SofNqRRyzzlr002956gibA4rMeJb5GW9erwClLPCTCvElMZycz+04/sXXpoV+n5W
O0Vi8AibjQ3HgTiljPlSySTdVQ2HRH+z0RUb+0WCwn1oPbT1CDBa0dViXf1sjSteTMpRxjVxwD1H
817g9FPMmW8kt5+VpezTS4Xzbm2h6zlL9qRnI2Xz05PXggw71NgQNZb1jPhkIue8muZZtsdEH5cN
bP1tBEM+WP15OL99N7DEDHV1zOgiuFrCsiGLNWrtRSduxlrR3h1c6vHyKMWds5JGWoB+LXIjj6ne
4b/jnX4XV5kNuXGJVSezrQuVhpevphOqcRATHpjDiKOy5HSTrFS4SEBD4LV5L8ehwD/oZpZYFb9I
DJTX60/Gtd5dCyX04/UpWvt25S76rgnkplkRfeKswjUp+JzaefyBPg/Z+0OoszqmThi4MLbLJeMX
oYBSLESs0T+3verpg3gN6Hwd+rysn4EcYtt9t1cuAw69J3yCkRIU5A6+exlENgYnfr+RiMSCScxV
huuk/sr28lgatTr0FZYFLKrBnw6Ytzdc4/d3YlDyROs/y34TOWlA088qtTkyr6PKQs1FXw5b7vtf
LMhfznooleeQxV5ZEJ0/wYMxiP35VMOLDcYvqSLMA0LxExH1vmt+M987gYwH9LSGCZt6qvJUvAw7
of553W8eXqrMmhOG2Fwyz/SMvoFvfGnYgWOVy0NJCNK9jJ9XAnvz3vEtOX+WiQpgjisxDvd/nWmV
ff5l/c1NDNW+byEuWCaDG9auti1yPB5IwsrPITZEi8FobgcqzvKTEBNhfPxd400Nkqcd1G/KCDeI
RiPhclwW+f0Jhfj26XDAPiqW4PxflDhUoj2lPP6fvQ4IvjsX8K9RYLnD5kO05TY9l31PRbUO7+cZ
kA7nwZyFZRIxcJLPy8b43S2uUU7kdLWcXAqy8Z7tNYdAkVOCM9i6vix+Qp5d6+6pgEeQ2ik0zE2g
2+n8mvn0O+6N7H4Bmc0O0AtxoQrniP62VgXG3YXyA9ETo4FFs6mWtVR0FNMnHE278fAEatHDFkSX
LEIFcKaj5wmC+cvOw3bU/VqyPl8ilA2SmozcDtdArbywWvWz01JeuS/MTAf3Z8YmD3WkkEt2H3cR
BEUA0ojtqmYwT/KJ+kbH8RRkpT0WFO/t0wXlvewM2ABYgelCEx2Orb42aPHIPbrSxYxBjsHkSNVL
tSBnu5THAuFgrtkRFgPYkQpQqbtjLNuB7AUtsjUw51MgKoNlUsHYO0vb+0MMojaVcnoTf7BSHlQR
LRvzl0w6i/65Jl9ZR0w2VySBmbxtdbEG7F3qcFIUyCLokNYdA2+X42wf3oqSnf0ZGQm7CUmqU4e8
LLkyY28FlVKKUe/GzP1MxuFJzfzivFD1YBwwwGLbfA1j3CDhd7XxMp/VwSprrdeXNhMEjmIpO24I
88GQey6CgNGhGTbCV/ctf29cRwtAoxjcr6hVMP3CDMY365F7ZQ/ouzqKliW+lNf01uMFJlEdpggi
06RTBeSZwTE9Fp9MtHiFKt3j43UmNae5SrZ2af/7QGTNG1qo4GBDCZa5/9YmYApdw8FgyX6Q+7E4
aOsNBL5Niqflj0WfYl/ZKVmuXwp2hNMAN2l9m4BXFSssVZN5evHQoqVLaICpLlebVoxCH3Pc2crO
5INMgpRzRcbnGrNVPBPvy32dyrIdhf3xTfxLoLdIFKwNNMssoE2fRjP7AUzsJ5JNJFnOC80qhVE7
hvd39sECDc8Ya0w7cAa38DsAphPyhVfqf9FotVRnUfcK8BgRmBDgKuUwLU6VtcPfWEVgzUEhIYvU
+qzTxpL4103L/7g/gMnXeOFzKzngMJ1W8aLdvf+GAmvExBht0tR7Nc54x/26b1ATEmX9WZu/UtZD
TQATKX6qGHdhUUOGxS7E3VJDs7ERv8LifQcGu9OFruSi6qSndqzpux0QzCb8dip0AEYpKpLOsrvM
rKbcOHy3Z6H9F3uqdRrwUkBEBKVbuzKcYSySFjWMn9D4LACzWOPICV/8t1vN4br5VBwZVgul8etc
1UhA62cy+7F9z31mrvFQ3Bg+TOkgehg8IwD1Kfzh9B9/xnA+yXraoQyirknK2Ec5ydKP7nTnwoLd
6Do5WghFDPgMq9EytMKARMKI51/bKcu1WSHWcYFKe1Bt8chGQpMpwMqdx9Ol3YzosBuRoq94jVTB
LCTDjyldQCxTUkHHxcl1ULzy2isCav5qLSncW3fRViZu8tP//77u9SwXL0Balj4+UqeSegCqWq0W
Qe56gXq/HdM5cTPditRQIZSjrlh3V1mTZoGcq0we4JgXTw0fjCALo5dEdgrXHHJ0vo3miSZOZ1JI
oYfkWIvSl5GOe2ml+BJ0jVtX4crKDJ3ctWrFNME5UWnbXzIkE/dSNCLjz0UNeqbRgy/W/OpuYSxY
782dfxymhemj0R+jJs++y3s7YP2WFrTC2+WJJUcCKqQqc1LxsLnoo3C9fiT+asDxAoKVK6lEUB1t
dzso/2lIwKRHVvsEovec91CTnAGqy71T4z/KK5E/9WlajbM2Sq4o4qP21xVSoi0PCXM2QTliXonT
iwf/4puaRTB0i78/77WOzHNDbTobBNvFkbo1s6xfQZGOjajh+MOGHMdzoeJkxx1QqJk3YagHMHnL
NEGAYRxK7XyD4juj7sEfDr7zEDVh22+4r3SDvcn4UtxPwTc+s04Q3cP9KR1DoiLZIPOPnMh/SlY8
xIscdZpstJfsEOZFPW2BHd/rFisrH3KvKrhVgjaNzgjoYoAireDegv7YpIut5KaM647SxwJ8OhQm
LJw+ddjowQDinpNvzrE2wvAeab88Q9gjwL4b9kqMWOFmKsYJE+GlAM4Puk4P+hpezIx/eJt1ya/G
Pd9LbRLXO8Tr6CJT/DF+C/rXXO2c301784KJpMfIREyhP44i1B4nwbXHdTCVi6SIbU9VtzVGqfSy
TFc27bJXdymAGJhuFlnXRcf5JBENTCpv8A/9ocL+gUZsmDYP55+wxe28y71xGGUlkeIc2zaDXbk7
5/zxPSqSuBces5kBJ603UjylRvdd6peBtxzySJWADoAVh833lr0jgn742GCjLkLmL8Htp2sG+xtz
UcEW8OZu8MjcnrQpNG4ftdwX6yMLlHteIONrQy92UZWcd84RWSsNoyG3BgarEk3blFWzJ1D8hEUJ
vXIo8Kkbb2+pYJ8a/TLFIm0z13NAE1uZmeuqOxyzLmBfM5tQ5Qw7HvH2W4LT4kYjZW5l0dQ2G3q/
nvz95CPqIqmHa38e6B/rvNuOVyP07TkaWS414issykpCa/enyzwt79FPyOzKIEZeXhPPQRD7PMIG
DvbQ/SNqMf4XLTqZ3pDAU29fcnED9QS0UicK/mKjPqgyeuCMtQvp6TBuWLkGwzJi+nsrtYzhxpMx
ms65pkNAdZdJUNBwx7GUqGa0h+PeeT6vpvJ3st0W+x1bk9o4e70lC6EatIwsfT6DlGjz9eUTlsyc
NIaD6X4VgmHSKJvmuU7kRaMNb4PDXXmQtcN/EnU4mjjvKaMsvQVNoM3YDuoxDMcZ9whbwl1dfCzh
4gPF6i84VcqTESbo615ouOLyElqHC3/euPGNRVVCeOItfQVCsoTeG9zbhlWUr0Psb7jWg9RcvlTM
G06+cyqzKxZGwSidIWY1V6K13pFbbcXlnPDPbM5jmfGD3rZnw0PEEhIZz1qmFQUlVuVnTlScwwL3
UE9zcxVtqTxR7QF8HoeS78qwNVvoJkzmUrjF8nLh50M32gdcUyxe3w8aEfQzzx10eeswrxKsAaGj
2snBn73ALtH6KusO1bjSmb6WqmEr4/JbMUKf827UjedmkvUoiXugnHigk+Ji+B6i8ApwPlln7pv/
JKAlOm3MSo/xFU4LqXWydDdnWBlUQXtBbs3JvTZ7XvM5et7TvsriChqEljU54AsfbOypFs/IP+IN
UWtR7wVPO/OLx/TSuHWwkFM/sdrHuoZQjNrb9aC6qjSUW2u4QAYcDnFb5MZXO4Ij4ydnvUlUNt8b
y9EYZSfEgUJib/EblushYkc2u0dXCQNfrOG+rLxsNvdjkNrDjC5g8Y7sNCQniGKLYTIxGB5/tZxA
tcSRMjDpx9x02Z/tnlUqihoVf3ElsRo49DJF0xwbdfcVpb6+8MrL+6l3cuT68+QQ1eVU57UTJuYo
OCvpIg/cwBl24Y9G1W7KatPBn5OAW1xuTfSYl6SNkoocaB+8PGzoTh4mug3ukRHMa6K9FVixoTFN
L0X9U2LIy5y0fo50YntLknIeQggiEvLiwGMkaPrTQLG7uoPVEn7wg3P2F6B4R0TEZ3nykE/JOXX2
n+dpTnWxU0BGscaKRAGjcEx0a+B5ljuoBKR9dsJO39e6iMvqVTeUmFrzCdyMd/Yj+tMYGcxiIvZn
Q3IbPIlRPpviQW+rmRJa35pScJb1nEnn7G+pp/XWgecE1oQETc522l0SfH4oNtY2yjkykITqPm2Q
trpv5WRwpSob4o/euRxqS57prqfFoIaNurJ8PEHUvDXFmDvedmWbZttbjPXRQo2C12oOaqiaEMOP
1UBvLvOFDcYULCrn9/S75DnpWksAyOsthpupzugKVG5roE3dZihfOKVU93iSSQCNunQSsS6SmCDt
DTbZOXxogSsX67dz+18cTfHCqr/bFpvt9TiYJZW0K1AwxdVQkoJcAiSsqGwJ9fV/D/SSbuV0Qh7+
Jbq9J8PPN0a2UWYAdARKh9jn/6r0UdfXhhiyMIezNEinfNFXYF0x7ArE7OVPgbCUrXUvNykYrCYD
40x79TeqN75TzLZWWo/lkaBITjz9GRzWRbn6pI67nucgwtAIIVvzrorjOn+VdSEBvqmqvCoy65Do
IBoKMUxuAodIM3YLtyBAX4j/a7TyFV23UfDslSLMyCk46Eu8VwVzdjvFJCUnAN2TLTI+n0zPCoNt
1xnDR2xpJvcgR7ps9WZfRh6PAzqR1UvSTxuuFK6jBV7v8J4c1px2PmpTJmWSW0/mQzM1XyYJ5a2X
hCvwUzvNIWiJUMHLgXLl4ZSNrlBABzMXDfRfIdDhb28s4zya+ds8Z9UOjdecJC6a90xkFM/SqU45
r03lLZndu5kkP/0LbQFP50CcBt4RPeUdJbeNj7wLa/gNWN8JoBdx12saLpeXBBOQOYMmMS9JBCK5
Ry9/KmSEzhjB1sFtjQpC+J8Ln9KlWm+je3H6WtqHJ0fFhl/JwVZUbgqLtgYdHmky87DaRPD+ub49
b0iaGwENWhzgFzxxsik2IPrQOx82a9Um2SDvFYQDNhZYrLnCOUItN747TwvIHt31pDIpYUJNMjWV
euqSl+vP4WODkNYr/xqN50SgQPmzqQtvq9bJsfVtXuCV+F5kxo+HAWMkj2F7EkmCWsxihVWr/wKp
5kJvQNeNvqEvE4R8lKEuIeW+GzQrfHzgcWJB9yVHZdQVzaS8j0uQJLitBLxb6Lg/VK2CJ3AEJ1oE
oyD8LPHX1I8E0VicImoJJn73gKyLJVy33rQpb6wKR5smlK+Z3tbrjQ0oh3L41bXhKgczgJHXSuWa
ReVlmM5QLUycj/sGck8lPszKfr+P6bNStoFg24q79URSk/jfIuWXJLE8+eC6mELPfmKSv3Cpbyck
16j9zkCgzdx1tPaI8PbYqy9I2uQYZN/26opiwK9ZzJSWSG8A8KR0sryddTsyHO2oXEfEb3wSeMDi
D3o6tSWkG2rTQSB4bpUkpMqva+bbwPdZ+P3Bw8ffZEPiU0I/tOR35tQv+rN04tGb0JmkTwnsMkqp
pHNKq8bhV2axTUo2AqCA/S3xHV7UlRpebUSjx94b9PZxXYe+hKctTlC4QJGo/rfVg6rplE7N17SI
QKZJBp4mXE6Y6QxLk1ubHgi1ZspwPKKCJ9S7VoCORw1ISuA0m/tMzWkQoqVJqBl3SC3hqicxs51u
m9WZmr+CrNMUsmCWb+JEe+3gyafflQ5p/yWO8Zxm+ueuVDR8Ii99U03P9QEI26pBgy2Ge4qUo4xr
hCnMd950ecyAK7kwEzm1gdnTNs7B/OODA37pNim+0E71uspIEK0uDlCnxFIIUIm1Vwd6oL5+3Vst
DCqlsCmkQ0ahju++6jWuihPnzFYBIENKlnsTAtASuJF58NT8vtvZs2Kwhix6ElOb4YbLeHK/imMu
fsbiN9I8y9294fv9rMQglomLBSJ5OoS1Shp4aPBWYOxHNJxWx845urALYfcbb2Ax3f5Nrw41kkV2
xfdSeGTzHrRbut/nO4CLt/San5DXAuYZYeWAEWbZ4AZ32SZWRxSGWBS6eCzUuaZ7bPtnHIMWnSMa
01T/mAN1USEFds6EUupNkQXnqeYmWG+pHktvpuAhIPANEBHJMgY3qKPoOtTY0t5sjMu0iO45IZM7
swFblO7ejJO8KdpRxCuF0tP0gBzd7wDp3D7ki5O9sOtsvIJn6G1qU1wLwlsc92wPeA0Wz4NdanOR
nHJHsvAU/WbI/YeA0Y0ECW7Lq8DDrDZfQAzskz0c9Esiy8waj15grkNjtkik7mnNE/WLUekglWtm
Y9PMTC2MwwgkqsGa6DaPUqqwzuyJ1tXBiSfGxO6w+tEJwap08e6bwiL4P6wMLuKV4Qq2jz3skD5B
9kKvMGqe85MfsHpeXjxY4P/RsUy9VuwNrlwHAZfDXi7ckroUDszMRM5Ho3wN/BcNuRPfw7Ai1xcX
7iBARclJN11ygeaIDRTz4pSeXtAkmtx3KpjpVqQx2P3zTTmRFcV9basSDUluF+scr9CBzwcGRWyz
3R3MtlRv4xEOg+K41jk1tSnvTw7bKB6V0Rcclx56U7M6i0e9kvAqNuVZ2T/58+4dxC4+mCg1DO9z
AvU5kJX+yvbfE4t49W8meSWZeji5ornz33mxVLIJmJy7/GrHwwSeQpYNxv/1vTM6OWRcDl3zYat2
j59Dki76546PmkQ0DhEnHchsA43et1XQX7euPZvxGiU7Vi8OpAYnGc/+1b9IslUi4Qt3oZWYAgbJ
DCmXJoIEOHuveNEigTpVyDmM9HCtb2eu3HEpBoMV0/8YFhsuc7It6p2/VkztWwy5nkzvnrVkniGD
k1K3ETAUe44qPAW6EOeRnU/fPcKVve42NGUJEI1fYCQtNNgi9WsZbnrKax+ecEaGa4zcqoLdWXTt
FzNvH/dbZJPdOAR6giElq+hIXAnYq3Jknrn+3otOsBymwoUQqWZ32sfoNzm+PPIW28rx//Bu6uaP
seqv3pvtuU//EdKhBXP+bOTCKhv8k9qh1Bg4BFnnG5nGPgRcj137PrkcsPv/lYWvxck9QQO2nz2Q
5MVOiDfvqtcOXceGW8tlAbVx88TWApG2Nfu4jdaHQiTzHSO3SgqGJjI1E/s8ep/0bDL74sIr+iVn
dk0jsEP6xH2Kd0OLL8KbqABZofMawdCVBIqW7Gc2HJ1TPcN1TneDW2DSHlzjSMibVjr9SL1C9Xzs
SsibduaOg8idv0a20jXNS+F7wHmV4bDV/DccNJ1GL+LInprSUHumS8rQBw/f6vtVxis55uu2tMdu
unnSn0WGO1D4phxBVc4F5wJkOyh2JwTgd5+IdXD08I4NVqB3+UxpcmcIsy8Kdc0Geukk3Sb793hx
xTnoMo72wWvsMLhAwMQII3RiILO8zX/OW25vT3A1+dga5E85KKLX72JtTIL8iX1IZT/BO/JL/DUn
Pku4aHxLsY3SQzp/O01S5g9az5BXq6hBaV2b02ONucaIJVaMD4lqVJSxNXsHnCp3QWxyGomxUQR1
noStZHTieVN5/s2sv50+1b0aOHSmIVm37rmficUnfwB5jiDCF26kcD430LBITNmKb/Q16/iahF62
Qu1uoCnP63AcXtiFdLliz8Bl+xJsMGZ7TOLcVGnirnZlrDgYJLsAzzqCyT+MEIfpg3BOvVSqpXnV
y5ZFplbh2P5mGFrz260w5mih6pTkBPAbhs8cYYwyhOFHWxbxI15VkUrt+dv6OsSh9SqIM8Qmi1M+
eHFydm2nUBDxDPh71E4EdDBWWLNKp9YT88o2jJ+6fItqnxsIxKgNXy73i/D8vZ5nvPXvpSuM7Wva
SeUICwxxLwe9CtcFmfYLg+5mVJ9B3hAFchUm++MVrz3og3LSU3HX6J6WbcyW6ppJYgpGhO8UgYft
kbRD2tjI+iGeybjvEPF9eR+n+mR4RFaMUKt4mJENWpHXSxTXAHWnIKwK3PL82CS7Hd2FMX+9AVlx
COGm94V3XZJg8K7iiOI3JDtuBPUK9v/B9DFdv+WNIybvpDL3k6a8lOwtfLNLTyEkLe30yihE0kGV
qkmpQgoRBycn/c/kLPGkRwhGw4PxFty9P+b+REauYw8DIEsIU2g3kCYrfQbqithRGH5f4qHspc91
TyDD0mAaQQbWw/u0kdSpWWlDnAE/ZSvedE4AySACHySbR5W7517IgUW8k0SS/NpuPdejOEKmebQI
7lwfv+svUIQuGzRVlH0QfRr2B/hy+Pk47rZPTm5IwMcF/LX8Km4RTXkLKiQd+skkLs5yf3hhCwcO
SfJCvhsLQPIx+RieUT17YWNU0GQjDJuSdNNfg3+gYSFoSxjT0Cs5NalIZgAn0AiYRpH3pWjLUrTt
oQzgItG9knei05lpbvOp9lF2AuOFZ70Oqe2qKs10sSEilrxT5qizkpiMbNIW2k0x102dtBVyZXss
89Ly1kYJ8+teCAH3EDimT++ifnWmo0C4uhEXlz8C8j6WaSwOWX5i3hUh3lw/rRqRKg7FdCqhcJQe
vopu+gV5d4msgH1LOBmUY/MPLDcwKvmziJYycojPMgMG1gxPqa618GLoFfhxlXrSGhfdNxHqIPT7
b4eEKLtE983y0/NFeMhPDdpYBEtHsq2avw8TjAx1CajrJP5aLwClJZ6i/VYEKBcCI3sXgYxl3CHL
AC5JBnpw7Y34B26Hv4Tw9vfDXDGTmzDBtiDelc+SeTopaX7a1VrtDpF8ZBXPHkv0XxI6oMjvM+ZS
OPJNyO3t7oTjFqIj7tHS5R8TAqeiMZOLkn/Mp7qA5zHMRQKkKNVLNOtVeQvlrlMndH0RmEFDbfiL
ZQzu3Yuk0UhvVz+6SoOWpRXBCTshqiSJqClM96ysCo9jb9Ck+rgfHIEabRYYleV+ErFdaO7j4D1I
qvtAxkhhfTh7el+GFz8WQvviCEL2F+4hgUq0bFFRL+oxqj1pow4+AW/9kK20D+iWQAk350NSd9cL
7r/ols/tpGsfykfVYl/a+n3mylaivGiMd44JBqxum7NwlmPIp/XXNOcDaryYo/yNhsZUAKRZVEAW
5ktYR/glTwEksyATy6+nJ/Yxr9QPzOlg2BfTW1OaH8keRnh0C1OaQfqraaYzytKGBkTsueBwWfNa
go4dG3PN8GWebkG1z9arByiTHnkzsvp/46dvwVGRp3Wace5FGQGxpmTU3VYrywIHhnphhPwYVg+M
nDTJMGnFBuCDVXtuCkTEqauZb2GMKOlELxQOYrKOBPqmiRbLiJpmXpMVYQIQRofiYBAagTE4RuSH
2AlMBWYg66WXLiXuak5OMwG9SvIUAeabpJITPn9w6zwazrMsu2nhSdU8HjI6UDHKkCYzix8Zh0Xv
LRijYIULzZH9MR7po9qRk3EfiG3dnBsz9VuNEKi8/uMf8aeSLWu1b2ypH1BX7D2JtEbP4zBaffYE
PirAGm91zseaRitAKlvBQ9pVeDADeTqN3nEYyHqvEUWbAPPVOfwHsZtQ+bhKYz7P8j9xZzpXGNfX
qz/XvrIwUFwxaOT9nwKPrm8ssii6GADizgr1E6+Qz8ooJtHwoat0IkghtM6qs8xDQxfyBLveGbYC
ILtTcFPZFWVBIQfABDgxFgOL+HRVnvS7QU3b4jZyKohNHz4xwiUQmYQ4E5Z/Hee+gQFuTDeQCejP
qmK8d40yOUsw1JXNEuB8E4pcDS7tq1lBO5pu4fnXZUX72J19kK5Fb03Yh4IWDuiqeA8bChAxWSRI
E2JUGzI4Rva9cFbcjOE1f3SrbtVKMGLT6KBpLDGE5OzTmkPnVx5vfjOjVmVYp/OUtB1/268RJll7
4JSzL6ijn7DXvd9QMneWFxpdme4W+wPK5Q5L0FnTfImh2ZgFQVPOa27NCFOnvQfIogz4BCYN+MuP
CJs0pneW3TVtU7on+t1H1ynGnyOsI8Gjrlb9oyNty78T+gsffHVjnBgcb2qYxYpCHj/rqcFLjjGg
JO6b+LKMDqbOs9j+oJJLZfdIDbV0EyAyzkYSHTmzsxFGZVXUgcVX5Js6qA21KPe/lAkpayZmQkR1
V8rZ2f6mojebjofy5koQ3uEpr5y+BUZmmWNKMxhOAnt9mlZMpgjFa+DYgIWNfj8XRAVhyjZwYypU
hrUrc91ReWdOn8YVFngolf9VJzvUQjA5D6zuqdJKgQG6k9Lf7/hmDoJabwy1Dxr74/B9n20CODsg
vXwEJ3fVGSv4tTx2PcGKNGKOZUztk1Z4UUfG9am/oxXNEsSiqdFCy/T6Xbe5OkfSJL6SDjMgbkCI
lD405rp2jDKHaSqOIrpQ8P3lgw4+zaCKdNeiQVl/WC50J3sNRa4L9odGdFrPEJNpWQ3CQGjvMyF/
jDYrUB1kBfjrKDrLnstLoOC7nmfYr/BNgEkWsPhdHUonvMsOhzOCxkmWU1C02uaj8FFQAM2eIbZs
r0R5MkdFFZc1iVJIxufUt2JhsZ3pEK12l9tF6+I+uShaN7Dpcoh/kHB9KDlNdk4VV4b7+vRNZI5i
GjScHhp/vNHStHOGhtopOFw0U9TAG6NGG3Z815iOHa4Z6zrrUOT+4CjkYF/SUk6QaEm8eVkKGEUa
Y9Yt996x8CnrMJxVAFfd0lzrVZemzXDZ/JFmG8+MpMr33jT0o1Q/T5nNBQxk2b+qaHmoQg4kzw1a
kSSCRUzSJTiNyWqnVAP8q/Lbi67izz/R/d2BsQ1LrzpmKROAJlCK8NG0UxozmMRn/H3nkERBKXRk
8hJVFdeTYV8INs9BGeMapljj2UfijP7pnVtQsrMUbr6cqaJGlwDZg++nkixXPYDbgjenojBAcwPS
4qyyxyg7L1Gu6gtjAaaTng/g4PQk1df1DUDZrQBXmQ+wgorUIkNGzj5MboOEiDUBKcoEorc8E527
B+8p3m2yH07bc4SGdjBdnHlAf98nX5VlVyWBMPQqmFTLcQqu1OeVJ4B3uZ8MgwqTnIXW45+goWfN
6Yu3hhb2znr5xgI3rdiDhjQVYzgJXSTuH49phQT0PxfWQN3U3riUuPMHSP+L4dW3NIXI44acjhHf
FuED/9aYTYhNI1WrFAOeYEjRRiymICCX+U0KfL94v+tpdYht521JSjaOLQwMXM6C/bC/p0PGSQQ7
oU2PxCKl32WjXqmj7iib6j44u/7gU4FTn9Jma3FErWed1xkoiRSg+s54K+Bu0I0FXZ6Evw+pe5Mk
LCvPuEq3jmS5zCZ6GirsEhbwhO8a0RPnR8hFOqNdjlgASmcA60L8gQ9JsiIxoh2m48MA+3FIpdT0
GB0DKWTIDB9mSohZeTWXC7JQ8Kx2Ku2Pj8NR3WBYW754XxIpgNmYkSoP2IopPyfzOHFEbTUiiKBb
sdShtoymjSKqZPUo7EUhn9RwrjJMX5qATKxHY2X+oAtmw4bWXlot8pae9SDWtsTFCE6dP61n27HB
1s+22nyJ9f62Y3nrE0LGr1Y8mkQoELGTi9cbBuLjfnzH09VUQDb7zTl6nfss75wG0iL+pp6Qkw4L
ESF/fmw4q+p9UfVl4b4YnaXkh4P6W1+he8poGe4M/kCRVa7i6pgxFVa9g67/GEobX2KYhAVgOCT3
J+1iBMuLu9YqIoJzlHr3WQAR7wVMaPmya9ah+Zjrt8EeMellBqsrakr90WbOWTKtKJpW0paUDPgg
cN4D7y+XRdoUJm4ybpQ5J4CqMTYRyB35shfILSANOvGa5K4Hu6QB2QKRrerjyMOkoPcktfVx5gRL
0xGZ1p0d4c1i+5W/F9wRC5T0w6d5SM8nasIM71mPUtuCEiu+uOR+jzdekx66e3m4+grN7Tg83ask
8v47HCNsOuYyYEMKOdzrvaBu5BjRVuwXKUjSnJlrKVxYxiB/hYyixgCM7pAsuoppn2Kh4P7MXNL4
BX0xcOWi+3OwR8DXfKXk2IBAdBJ8PsYMdPwrzmCdJyiBVdOB29Y7Rv97hD2zdcp8/7kPatLQR4cw
5ppdX3SSaT5DbHg1iNkUo4GFacy5Q2oiPssYKR7uQxz2wCA1gvphLHT7R7crzhUnRtxQVrd8fAOy
xaj/PADffPfYChg6X8TgJ/QE/YO3L8jlCTldT1DY0OeTfkMBuNObKzqkEDxAcOCZmLav3kl82znw
HzBydG4z9aEkmMaD8ANDEoq32etHpD5UafAgsfddybvu0SJVNZULXenJ1ro/akLToLtnNx5djuHl
DeLBhw0EQp5Grbcle0PUuPqTxHmgFWvn15TBjad9dU67HV46ojdL8iwyXNapdTKB2KjKMQq/lA1L
cHPCk0wdbOYD2PTvu9jtA26xOKziJZ0DGmn0T+T5hwnhHDUjBCyAj3H8pPzptqlSGo7U0joPV6aM
zg4cQii1KYgtGjsvVQTAHeTj/ZkJqw83CTF6ks/p9uWSwwczdlkhduQjP2qH17njthz/qOsUU2xN
mjOQeLe5rPqFpUHSdshVBBeCFXnOnHuQVMfo8yy0t6IF8Cv+4pjsj5UkQIVGuMKGuxL93faFOvf6
GpehXFaoDmyMKkEJoypqbzBZnwdnER+inLUkSBYHV2wKBpzWppchBAHWcpNsoMq4Uw9MlxWwfcRJ
DTHBr0EM28iARuU50soyOgwdWelzyXBoueV/hJJSD/mq82s+F3hExoyOEE6eOdVDXz3kKBIAFG8C
ql1IOcnRE4XWIoTA8ti+gtxshFn6zHpZnFmyy6WLqA9Erh/YBY6hHDNhooXrwA3zqZwmfqw6P0Dh
5XWt3YFN9svozPIPAcjqTfqhXlzrwbla3IIMsc0pW5oOdylAx2faUCIAJqmvQHWOQrJm8YRrZyfF
sF7a4WKaK1VTf+reULhAGiat7ls7+n6Kptky3ox+PGzjINagyBEJL5j3HFThnfxEDQY+icpqqA72
x0SS4CL0RdHbcXkKnNmXFxRwPZSIShb57DgoP5TOoGw136zZQPFa/YfCcQ+oL1ewC1iypLTTnWYZ
fwCm/PaXgbgZkvPKunSqzrZmibB9ei21ZwWlkrlCPDls2kewJp0nAhCDP+cBHG0WfFpTSYKQbXz4
3Fbb9SIt5X7/CWvIYczs1KJMZ5ESLW124bB03R0m/AMG+wuzUQ4t2VmdktkjBjxFm5xKoljafk6q
PCvRuMNUjhjHFUfn3O9SX+WOQKReSbZHe21NSj6idXIQX0qk3CpPI13Cs7bk/NopR3KOlstHlF6A
p1hpkGd85n3HzHj1t3JpbBecK7WAb/dRS2FkbcWOD58T/OrwrKifzaXwhbT7hsT4Uqr45JnFZHRL
9fHe7wUgj09jnFMTvf4jylUDVLUfuTTohur9FqpZl7gZzwauHYYwpLbxQ9pd3pe9EOOgaXxLAlbC
Xvs9XbTCody+qAyWabUy/9pys/yHZfy2vzU6ipyV20SiJTXfRkibp9rFX2uSFYk0vQFoaTbEIujp
vQ0pnW8nxSUG3PTPrcRKnQ3d+sN3wpkkMu0ffK8a9RkE2zqIem0YyaINvFNwyZeviGctOC6XNe22
4h5V9/mYHQB1brD+3oQLMvNYhVTX9NYmVgPSEy9Es1gNB2molJ5Mx0z7FPknJvThLkxHNbZxg0/G
uj+dz/FzU2dtAD0JnjkSGs8iBdXmSr8jgPLKT+irFdsSvv3v6lzEdndLRTfNKMoCDYrqYCS4ZkdK
q+8nRzBXzMTwoN1YsbSnvZa5qIfY3cGW6Y0YE9UQnjop/qxpF8qcLeIRbHJycoLfJmhK+rhlp1Xt
bG5eK0aB/2vI70nU8O0QQpsC8uWh22IXlmjga5bHhrgAJjSw3kJ+aFTe/c2iepRzsq9Kx5CwXf6N
TNGGZ5F84lwunDGejCiYUjKabiNzKnA76oWNayo0UabsWhfKCPF3OZ24+Sn021Bcdh6LIAhBZucZ
+FEvZoyYHKy9ifzwL2r8DPLIJqDDEtlFGDhiHtPIMGGcijsVV8ChGWdK8zSdnlolDP33yO9xBB9T
/O7eW9nlZluKu6UT9Q5fDgD4zTJG05qIbAk8AlfSgxBdlsShjFi1eyjOR3Ml5Sq3UqqWJ131bTIy
vQMg1KpeWGUeS5lOeLpx7Y0NAYstctC7fXkCx7dNDQUFsKLvzw6fjx+47w7epEELBfokNacoVUZT
H0XRqlT1j5y0ozzXpMss4Nw0n0NcM+aPnksIdWMExVJ0FK2hCZCJ1YSJtdqdAoAlvvIu9HzvBLHf
KuntHWN9fm4rqfosm570n9xRrY/FymVM4t5xKW3ElSqhgfR2/Cn4gmlHAuZE0Xr0EJhz/qapIQ9k
KczFv7JRmmbqtQcuiGYXY9AalLBa5miNcdfd9cZL0qnsgffTJDKl+5Qjo/G2rwVVCXidejpXEWxh
nCpxv8JJYN42vTpkTuuxQkBzJj6z7IcQf1oibCl2ywJR/4V66o4vdTk/9dZqCFPmxrfHY1BUGQbL
edK+tx7K3BgdCo+6VhEZamrFptkmdh+cD5rLNHPWriOVpSbNsPuyuxtFJJNKptW6AbEsKGp8sg2A
ScxaObB2xIDnttXSebnoGWe9JhqWHVrtYwlRN4vgyy6QkJfWN4Qoh/CMAlh+s88mAbqOllMh94l8
4hE5tof+7hRKMhEqJj7oEGa4S5xeJNRXMQdYgSIRgcky/em+Tct4NRGHOi39NXfkt3NmevPYNOSd
Wn/ae8F79JG33CKN1tyjz1gkQHB84IIcBPOXLoFCEZXg+EX7WmalXsT3zw6tGsgE5cA0IovzG29l
vuNwLdqR6PL7keSbCCMYhiLfV1Nh5TU/IcOL8MyGvt4hCI/J2DnUF1G1tjM5V2QaEPOe/zKRN13f
S2No9foyXadEt2Xn7KTJWFH90OevgAtnsp90U5BfYb7uoNvEb7mPq8GNbu7/OCvB3GL0Z2+ZNJ9M
LwW9yTfyIPWCLy3cLlaSRSN0WgSJpKn/I2OcHkATnSIc6wNYh/8Dc5F88Ci/l/UEz8rm+6cAuxfi
RZvILNYn711xRv4AbraevykV4N3xrd1L53AyeF+MfadLw7EK/JjX4gP25b5zFlIckcTFHfnvIOXL
HBtXRv90o2sS3JR6a8IPzWqznqTmfQTPVpTvyphii/P6YRxnIeIxojqEcnliWyR3szySkmtgVoC8
vnVLfvAh1sY7b5p0zlZcd6HFGq9aJKOPNrD70agejWU1xHs3W54F3IskOZ1QcLRNEOWzAwFr0shn
nREHQpAaC0ocGc7xtObZ4o77HAiilAb4NcMCRDjSUlJZEXdHEaf4OzW7iOo4ApefBTVoxODqnN93
Y1IxbZistCUiXroO8mwN7Kjv9a9A3MnLFs3JwzoG14y6OKqZ5hppkANuNHMSCzNjXblcXZcMKACq
3klEC+04CA4WjJ7eEnmzzpNrPR5kzmeUwZP4Bkajym1++wa2wvMvf7MR1D/hZcfS4M3kuJYH1XWK
1eEkKk36qDXWRWEC19g9iye8oHPHIAP/akUn50FDa/7o6zLFlhW6f6EaSav/IU8jn+QFImwamvNl
V7E6sc+F/eUywABjQc7hhcKRxz6c8jhn/+rfWoAwz9VS6uSnIu6cy2tHPOuBR74mWnAVdgK3F4uK
7bvFoGw9IqZ84Y1h4LJcmSHpx5GznSFEL0suSvckOKFpZU6zFVVcqP1Y59ZBkj9yoImwIrLrEQMx
VuvvOA4fpOYNkG2z8UDMblghEvH3QSTrW7W2xbZ67QVw5at9Rf47broPvuBoB+gk8JP2mT6VzQ0B
nImEkB6zkBFwJLHNTgOeaM4BlEFOFQkVx+MrEC3fOYaQwtFVOg+DfOzBZUqmljiRxgmQ1Uvk+KjO
Cdaci9E2FmAy3T2XSX6uKuXHCq3H6iBmDBGrp1rqVYBlotu+mY/x81fD7EHGVz7a8kDkakkTFAWr
PDVOWpg4GTwroyhHlPTEiZW5lroyuLrA3Difun/xFJO0pcVqUutM1XH4DpBD/RmTDSBxKtWH2yEC
QG8EFea78XN5dUqVBmQaL/ry6QQsHGENpCU51FrqmaqPLZDvL76EoOi5x80NvFIG3FJWdjVDh+1d
5Mhxls7u3U8HHlTDlw9t8HUpTAOEorDCRcSvT+CPJop3z5YfgUSqjS3/RCyuFwgkB7T0ELI4mnjb
cbNArZJhZMu/bjHjW5pAHwyXqy3kA/UIKg9bJVjPQt6Vl0zGfemTY4vr0BDlL6pNTKisOuFuWmrk
Ug1pA6vsKA9kFj8FBFUedQphtu/h4l8Snr1S3sa0GNDol+tsmUk3NpYWis0QivX5urdVbuixnT6U
iesh6DMOmFCICEzAGVmFcyBsB+DpiJtkgqsgssGlUFFr/AxU+jdvysKFrhC7cQ1tNV/4dsiuXVus
sgC8w5hwb2qr8iLYDt8ndF4yZMOvoiARn8BJId5Zsi0EfGk9zW3YmwINkuI2xBktxZhLMNhIVrMi
3uZX9+AUhgN4GNYRqCz1H94yi3bRqDneMw1lq/LZn/2rhSmCoPlITp2oM1EzuhONv8hqGJDmyhke
FaeydhHIvIsiuYGB9CmIxeX7SnrlooXKu6LC5lzcl5jFtTQtFfbc4rL5TDz4YXSHCU5slO1Xwl7I
FJhEsIAwL2Or7fT+mF4veaDceVXVN8w5f2GEIrAnfpEboRtZb1iYUmfTqmSeH6Jg/xdReV4CJoO4
btqZ5AzinJcOdaIF8rd/ChT6lHHxYm3tV99M3B3x5g3fwfQZMlrF3FIdXOKe9TZbSz1RGxj89TsX
poHsOETHmukfj7/Ck/3GPHD7bS8sx9H9O1R44EBjXOTZzZn9sgCklotX/dECDNKFPNZATtqJ2fi6
eHoCOx/eTQmWBxRApNRO4+day5JesAtjBaVTgkvLdoaNWkSnE0ZK+G3G65AX8CRlg/W/YP3zd0OV
LTKhn/hP1GYjTpnH27awjTF12KorXNgK9iVBVDQo4YSBlXw0q1K1NWhLN7t9Li/KBggDlI+kecbh
2gxmRlATgaFNmWVP74WYq6k51uISUYM0bDpKWfr9tmp3/r7Vcj0uIllmu6d2vIzUGf4AKqcUDqhL
h+R8Qv+oCncpIPsJkKpY/Wp//Jjf0tEA+0REYFSwSOKJHgim2npuaPBFRMIwsNmsOSWZOt1EDyDc
5wW5/oeQGY5DswVW3xIhwY6WG65u+VJek7MHquBRhRfXgcP8rbmngf79kRNjeHwxo+PXPRvAqPOf
mw7cH/Ow01S/OojJ7BaQdD7EIYWG2lAfj5+sd+T3QEoDA4g0j2hPt6e4XI/i8k5/STSFZk5dll9w
GSUaXRYxt2YjKX+WqVFqyJzbeH8AGRQ8l2tcseRTef12kSGRnZsYqMdGHSrJ55aBaNRwsEoIcTcq
IQuCBvLtUE9fscWCGzUyq+JCmMysIFsU6USuZYuqacrAsBX030Pkx+n1hPs2f8P1vDyfK/cJJrGJ
XKG/F5mXGy1NPDhjgcPf93SXrErJhnJWRH/kOLaKvQyZBafyxtfh8/I814qhbb9z3IigVRbbvm34
xD6m+D8Vv5nU8BQFpBQLhlzs3gIGWhvoLVfkLEaYmKHetkaJ7vnyiLYoQ4GCm3TDs1lh8UhOYH7F
AFP94cKOGCKn1ZLMB0X1n82J+c0g9Gz+CM4bUntEbeQEX03JvP+k230QuqJsaFAMOV6WPO1oP7yP
M9e6lsy5gDZsuo+EIL/v8DpvcrXepYqmPuLIcUkCOnLhr41ghCI8P6RQzg/Y3NUFJ+w/NJEQNaGw
NGuOXVxuIZ2NI1YeGyDa+gtRiPp53E5fDCYb/TyhUyHUUHZediP+QszPr3rdFzrRIQlOZqTqaKHM
yUx59JkS5UKiQqZ4xyB9UpjPxC+RY/qBN70rOdwxZZIpJ8/EyrFAWTA8VPHd9FmBJouRu3n1ldxs
An1W6ilcw3OGxgefrfA35zoBzKPo2sMSs/5lavqNnSJJNx9tt0T9DOsLHEOcTvm3ZO6nyvFS7Tmu
8UtQyyX0t7l2bX/A4d/9Iw2mUjNCVAtHjKEXkRCzdyORO6cUGEkQk3PW2aIZLbONAleVf/0Kftxz
PaWxO43LGLDOKAu6olMfYataPNC0KIZOLLfrT/sr5+TXRTpNd9/B/Bvs4uFo+zK9wHzhFVe0p3wa
5yIGf8pfZkjBb9Vt1VxgIuU0hkTi5v1lr3HNKWpetsQypPYvzM3LzeohMmV2rNSyvpcX2VVOpvwe
ifFf5DPSSh8Ywn9y6NKPTnI4yNrhstg9Zitq17P/fssAmDG1IMxt0e3+sZHC2f4v8wtv5yggI4Az
49umeSipxddZA0PzDzIoyTGUQpXbhSGthOgODQVsypWucV8aiPBvbdUsUUEytJL+Qrkio7oV/UnQ
268MRr65caOX2vSHNlHVC5psot4lU5KGk361y7EnwMrr7UEkui2ZkPRndbm9wwHMc5SgHuQjP+MX
QSJ0e5IGXD/M1TTlr2HTJ/oUU6qE7z6TgQCcMT+1wYXAavvxTsc64LGqk4OH97XIGpEFlnpPvgeh
aTtLnSmKC4rQgNL5A+r2S3EtNOkPegbAC7bMp5AxrAyUk8z8Z//DMDuD/3fyj5zBLVO2qX6TTSu1
UAjePWlaOxihlzsf1YDFnfEs/ObCpWunNKQy/JJNICB0/apE+VLQGok9zcVMBBNUcRkoNoDFyeZo
g0ECGh8r9nCfsX0EkBphW0ROWQhTN0puKScni2tL2xBfl229SWjoABwUHGyWRfvRXSmT3gi/vnHx
C7kY71Mmo0HZJHOztymApBhoJ1fu9fkcNhubGQ+Xg7fdOTd6LPAfcVGTHk0jATBjb37+ImvvgfhY
7SVHj2RCVUMa48VpxOr3qmrXaNX24FYC+TQVtXt3IgR9LvX3+ymlC61mSeQizZ6pKi/DnFm8wT9B
hBXIMJi9cGL1OAuhQLa/EtkDKpXmgLmX03wu8qhyOTPE0PkQZZix+D0/yWGSzAWiLuyHZEAXkwe7
4bl+SmE1qOiP6vgF678k+4puVKZlmpA/xg2upydaKefKRUf/LcG8I5/cJbdYGazMCz5AV/Y9TrRm
zT/CyCY8yUlefCP0WLQohms1PDNo4KK2D3qYrYKDJjv4WyxoJHBgIG7wlV2b1ZaC5QNL3JwQPFe5
WsI17i2fyOOkUddi5zPXZmhHmfWWXdndiBHPAI3ZWgzR51X255bYmz6IsUYlQmeyAvZ+6+yI3+K8
Y+Zj/htXz4x9H1cGtGMrqQMciVY/MUzKXdWV0AYim1U80Oz2h2alzSvb53nfm5uutJx4M68pXqkF
CVj21rpCy3D6gqeHsrqtBh0fM0mQ/QqSjVeo6pFwCleiDGpbASdcXxZ+SNhjtjtp4EZNG2ksxZhf
gFZb3dg1WYASTcoBUpRdqyarR1pgShmWs8VOY/cETW+rM6X2qzFQ/KCC8GUzb5T6S6SE31XGkPyY
Y9Xi+Qy5Qaiuf5xQjLnuf2N+WLMxzhvlWH+8bkvchv4KDlHlheZRk4n8DXYIxWe04r1fvkIcMtPZ
/Eru8i71pjitv4H8GxjmIPmELBcvWbMFz6LmJRXTURF4SZ736BzMJRmzcnOjIamDfMfYcnxhVR1Y
6nN4E9z2/0E0IhOARyOfL6cuBfbqXAH3BaRQQ9UePSe5TZ8FDq+tvYNPC4twRZBa1KLdcQ1q9dIq
gRxU18vfUh9qit+8Zgd+9xD/4eaWflKMXZyK+vm4pljNJ/aTrOz82vi7AWqmXmVUXQLDS6Qr9n4p
gyZZPHWypDszjuOwDGsuY3fY7Ffto9wkSDbd1yp1kvB582xPdZHRiHWixo79KSTqcnf5A0QWsebU
fKgvDFotF6J9Tk91FxT7sIy1wH8Hpg/8afc3+5c3lF1bw7w0gaCeia+u6Iq283IBufHD5nvtNrs1
XpQeZMoY4U4TyUuDwxHckWMfop6g0tkLsBmIBaHYgNJIPJUZrzFm3dqABXF26KqO6+k3TqRbuV+2
ZyMqKziY0Lx9sJm2yeE0LnunYrnI6GEINHtNyt3Uaa+YwSy1BpwoM3E6LtP9Ezw8G+WVPmkSVGOz
UYC4IS9YUGi9EL5q91GrbC1YT6w6j5vronTg2CfsUg7Yj6fmkitxnlDLPki7BQgle8r01WWpADue
XiP1aekF9fXnBKmqezR45BYuS5jvkP/TAJ0CACowI3lWdt0e7paBwyImmE1U3pMgRR26xaNPs8Ub
OxuTHRiAtJKC3ceu6TpgyNTQdDNWOwOtE/jXrrH6rKqSyPYe/iUMHGp7T80OsIQRNJjh6bLhNTO+
ErBIj7KiVaq44oFd3BShcNLqelHCFp8Lp+hCmxLTvQgCEJriinjVED2S2lRGCJokwB+tZ/Tpc0+R
gA5j9I1htFtJicxoifoxQSTfIOpFX3hyVtmSkZ4Q/TjmnfBDS1TmxsFptqomRSY66MK8SMnS/E2L
zo2hOzwQHReXG/eWCAO7t95F9hul7YOwL6b2ran47LbBIXT2ztYNSyHOlS5AgzjZiZgDKQWwiX0p
TqdSioLDFGJVp4OU8nsxED/8wxbn3HSEL5DhEpDwepXkMq12mMjORF4J9y8+uTYK3n2/ddUit5ve
sg3mTtXLv5SW6xCRKwPxq+6iokUvQF94t0TO2lnNhRQ0q49PZtBeId8Apgz5sHIs3DOYRzW2gJ0i
aRc2rfN+EWxXm5wuNzkTcNq+6pZDzI/NPaO+67jOkTgHaSTiemOHbnjebYhblaFN4BTJLQTLeZnu
p7tEfcVWGMeoxivpPSYBpKpUQvND5gaTOddWhhrqwD/H80iKSEGo4lNwDGz26kfNHG25OdXx9rDu
vCe6AS341BJLZl1ACCfhy5vA42+0NN4lLnJNcEUW2krTwp7uQGfkFip4pMe0i1t+8Non+j4AT2EG
srGDxH9L2prLY1PGFO6jU9KF7eoMhPAhlGVs7T9UV32Y0BaVfp3rOxw+HU/pHBbA4HMCsq4oC8UY
zTIeHZIN7/cfcSoX9FT5pevCyE3gxMSAJ9XVSnNd5OEmSB4iY5qCRMHhrQ1zYHlZ5yVj4smvljKA
iyUAKOCPsMR5Wo4/uKW15vUlw0vv9q0M9T4jNwYi00YKKMpNuT4DCa64okOP6sfPSxvOh8PYYhba
flrOje/VqF5B+25btAhF3QgQxwY45lUoKgb3xBXejr6hN0eenB6nKa9Q09WRshfIWwUCJBwDljuB
uJi86UZ4rSJmaICuhoKvMTUPdTR4vCJO95uBHtCe4AT6ghAoH0QYDDUxuTnG7xPs++gSuD6WtGGG
LqxKPNE5aHc2YYrV3q+tYbPy1aIn6SaF/WYEkRqnn3YohONjuCgXVfL0P9uPHFRFzlPEEz/mCL2G
auhxlpromndVkdtPD3whf+RzwZlscCDfTVkcs7yLTcgrXdcEgWwMY8OmmTwOrHVquhq3BT3hqMUk
1fAQvxUYoV7KIMD8BloEnqXZ/9BRNsT5FomJQTdweO2jf+hPSqL0PoRkox9fS92x1YnibI4XqUeL
ph8Qvci0Zu5Nny0b+Z75brjMMsveurHbg6sa96VdS6jC1xCLbB3UH5YTZkG+R48ZX5bhrqdC54Mj
mC+CITGD/wbL/SrYPTnkMsyCCTb2QwYohiqDloJHZAz8eSEe4QNVosP6xWdg3yKpWgdyoqGUdXhM
8hItZDhfuDcT/ElUuE/PW3N8Jr2QrJd/iJOUD5gZ3LQ84urD4+YYpKtoOy3iAO5/3yL9yZnL5jdi
xxpSW3wScjmG6EE2bSE8iL2qHj4NrtghbFcXd+QCEzkwV9SnTBW1z8GRdvUC+xdq+TvnKLAoL2hg
WOdqMuK5Kg0wbCuLUNJ4qkdsHrI23xJD21wcCTLrKBAgykUviesarYuIzWxw3/me9LCM7UQUlOGp
SLOUZwRAJn3VG6XxfxVkPKIqMNG0s9W/QDO+YJCfb6qwEJFLedhtbBfShurACPypedHsa4UASpeH
OuH0KB8+rPiP1i77CeBDKrRpq/3Q82VA/a9/LKpJ3C5xFZdWVUUL+1EXvrzW0N5EU9fOBALumRAC
rIzWgP12KsdtodrZz3rHll1mmspZqKvIYokAwWn5t4O5w4qxD3UysohKUKTr8uoeZt7X/hnVLYlE
JPQmtazuRA1+vgNdPMJA0e3zLP8uKCQbGW2iNyAh4tYGj1nLExDPc9mQ3Bnd6sz6lnDPVDdGLs0r
wCacu03r2cAz6ZadXtLM77dXt/cWffsBvWwwxjuxFnEDCGGZlxUvjYMqoxZLdgr0vR90uyczwBXD
lKY6d4reqqV5ddRGjDsNXN4xMG0/RqeCjWOqV9VFdA1Z1qDXYsALJMrqNVG2br/+usfvdHqIMGeQ
RegNyiHsRSBT40BPWkGqJ57wbFhDTntYj8pcjv5/K/4A+Ihz6ryElaUH7gjMR4uGUZLiYk/Hqn4Q
7yx6L+JPaupzr5rJquCX0r2GK+9Cr9IsAwxoGdy3gJfPTVEWEmeU6+PmYRrtrFsNTiU3lOnCW4UG
S+TkQq3+7+Wg8XkXKyDEGi54eUo+fEyxSLAf1p5ml9kVGKm605VaeaoLfOIxEWGIVu8jP15LEZAB
6uemDU1Ls4yMrsAnO7ga23Tf34Z3vzQkbtx8GogSb7JuD+1P3LN13+9SCLa9yjfjru9jdjQ4Nvgd
3bNs4pwcqG2wiWxQfida3WZR0zevMirx3E+E4hs2XGUgjMa3w00ODpEA8fuZhjXKz/clYZUyB0Z7
R7Mk9yWRTPDALVPIzLuNcHt6uk8cGO/7oiC3woL2uzxonlZxssDhtZy+H6xfoJzrgyNfgCl/s6zj
TL1+lY/6YN8QmcxCzCuqbyAF3QQ8F2qsHVsyck0YWmGvcjJKnAxV6gFXdXggPtojTtIQlG4NyDBr
n9P4qhXNhL57Tt3HJ7yKvN5555mQzNU2OO7jxxkPBoP8rubwqBK034vIa8YL1qa+bAYba02oMLxe
V3UcYY0+bNT1QuiztH8+EqPe+Wbdkqlp67PNNofM4GRAtZJmchjWWilUkiE4lzGXA0cQjCqujiw6
dVQEvRzsUthsyMEH//5/AnjfsVNGYAEQ1l9Ct0Txmlf4LxCnTR8yPlFQ8VjF6q9+npjG8d8MpgNS
grsg2bYL72h0e5w3HhFVS1NvJoYme6Na7/YTcpXuLZrMde0aSDIjTS3qPHoiaEcAOQoq3IcXXw91
i7kI5rJgQWkZVVnVNwViiUIp4y8WR6flEBhApL94oIzOR/cZeASZza4JOXEUpb0lXjwRqob9zvIp
yT+qMpI0REDWVox40NPfY/rmQ0f7gWRmnPL85/BHwXYyfzqLxoiWE0IfTto4w51e+n/K7sdAIKQ9
d5XM3//Cz3f8XKKe4ja+uBdJfiYP059AbceOC+f597iki/vezIwxhiboZMa+SqJu1Q7hxozeOfor
w+D0dln6UPCl1IrrdorpjavYlQxBvKPUUFVZV8Ef9FSNWSVY2nm9h79cqruMmdl7dnAEf0lcCrof
AoYbDVCOxCWP7hkR2mgmsB3lqMMr6oaiTw2CE4A/KsMfojj9CF3Uf4Z3YuMkSuOioqr3IylY4DPZ
uICBc5DnKgooYokvK1QFGfiQNsWyNV/CoNDPAy3eTYA4CFIcXFEqVDMCpfS/D4vFgFGxNYVOxd3k
myA4ISlLAQFAGqTgaqn/fxBOJiAU8XzqfykAx43bdQVx8jEACIfxG/Rj/1u8ktPT6vOJOY5bkCST
GqT87VlFnS5NDfzN/AweBg9wNqL1i3DpxSBYiUErDsMkugxEJrN8itYEFxpteIghreYlOxdsKtMc
AOK/3b8urc3RvMUlV9MVEApBKGU5szUEa3v/QsFqBp6cLtXmr9zmjSUYDrtiXXSWXv8U/dhfGhJR
HE0Yc4e69KbrlwtVVZwNz0xUxALw5UAswLLe11aYn1FwHsiNTnoszv5aPseFSEqSkVATX61FwWUt
1+kNh3VadJK5l8Xwnpfo8x0P+AVSMuMnc2ab1BL1tCyE7Z3es0lpP7VTMe3/xdBGI4+wR9Cuph3i
dtmBPw1PEv1bdMespdTYvNUX1D56Mz+wk4liQgvNVKAJNd/6JpJaZewSqLx5iTYSKwQkmXwlRNfm
nZcZm8MqrH8hziC0slyyBEjnDvB2ulRjdBVo8GlG1I09ldjDMd5wwPE0ISIrcGddgmfomRPV4pac
NIRkkc1aTIlZIrJdsSLCCm6wcSuE+diZ07v+kxowheSB4YfP2kHay6Ok0yiTMphNZgJTL8BRbk6y
/HgsgHw/BS+8kSiwhKnJWz/97ZlP8aE05VQJB00oKIKCeOkiBUnElfIZaJ+ew+YynjDaiPlClWkq
iWA8VjYC0wlJvif9pX5AwrzikYyvpHHT5OBBOFP/CRJtrB/jqgCFF5QKU1EF41hiaUQN1DBaD4fb
RWJhX8ucUcEMI/4ziiZj2eyvmSm4zsWtbQhIs+RveZ7D1LNaf3FoY/MFfryaECKxnWiaWnVRMhVb
QtsfSC+3QiciFynOYwQ5ZJJvYT5NFD0MtEdyJ8WblH+jVz2NxKR8dZS5XKZ9ePKIKHPrIINFVtB6
HGpWfXiAl4kIkoZf/ozTH+Ya4LRZnBRkJJUSx+AysskXhdVwWkwHQbXcx7malk09rVMjGDv9J2RM
Pg3meOZuRzKcnkCF+ITW0wFszwboES1+uW5YgRdZC4i54LpRyVXHV82onwMiNckggcK0k2s3ay7J
PIkTZOWZfilG3zyXux+9b8WxO8uvagLW0XOyj6OW+fbqREGDoaJC3QPnD4Pw/LQWkbSWcMntjbbt
n5VgIJVxigS0rwXAAm6Zb6jCqwdPesSv2hYR9LPJV6i8DXPrDnJVlyv6iYSG9miIK+0pFQOi9zXi
wSRjnF85e9QVJ1LvvM6aRfT71onIRFdbamg4vQHrCyd4gF6vIFnnrTMBkb1pvO2j9+xzyRCwNEzQ
YvEEgCmN2H7I21UvOz/Od604MzsQwFOSPcFo6isRs9YldtIGsl/bvh4zZUGdDbJZ71NAsp/z9J+U
c37xgtmKnqONsIwW8RXDCD8VeH6fzlqNb0RduOMQLj2SLUAMtCCkOwWF/QQ2b6WaLC5HhVY8s0xK
7PHG/Kf1C6YSkwk7eVUbvNnKh59ktHnEd0dTxRDhuZP5ttC/IXsBl+yyLtsunhosB/rj5Ko9193P
58L9RA0/cxn62XSHoNkRUoGpHKlQ/oHe9XwyLnccSdjlvbMmf5V3Jug8dc7ABXpFoYp1BbprCEpg
3F5QaYUe/lACkLYrXLvTGAuiA+cJ6ewXByoNV5M8n2V7g/2zpthHAIPfIbMhXL2bfnoEbLF5su1y
DijaZUqaCjzuy/4XC+jeehPYUQ/6OD5VcVNHQU90FkjVGMqdz68xo2HSGs+AU4zNe626siJVPYRg
DO+khzwal3GbwKtb1fZ/6pFJTj17zUOz0YSI0nLtAhApcls6szlyiZboGABpKea8hkb6cIJHesUT
SO654ixGv5ETQhQKsIp2W1ayKmzml46ld7zBXpoCJE83UL4ODMRk2oSMWPNOl45TScXfEEc63q93
hNbIeRJXTP6WQMOFcLg0+CdN2ZWEDWq6FcNc6skPHLaphSMilDoo88BRvhxc/uso8l1dvpptSwbM
gN7UVUk/TsHIWtssAR50A+7LGfk+QiRA+Q3G4vJK57fC8vYSjEYyoGSA/Re0pyvzMSaeyxOpWFvn
T4mesvKurcccNIQVffJI4r6NDPnbFToFixi0il6ER6BdwilDBAgZ//i3JWlDR3H5lo1UF/jdFGuA
3CaUhxHA2nmqH84MW4e0iAc9K0rKTAkgrt+/nMSqaG8s0O1IIJsa/9apn95NW80GmGwRUq5JiWxd
tlQppWHOQNyteq2CqDaiEzdC8EeGp2GXQm0E5J54AyM5BFgyN8G2HqfqJJZRQHblVSasv/T7ix3+
wvYX/qpIBxRo+cvQRrdEh26xbRty66tD4zxHFD2GIyV1KXjOWUVMuMnt8i1Bdl75g2prWo2Wz+gU
2Oxeb1VUGspoMbMMIcr7TbiMhETqcZ48G+3jVhW5ty/WoPAssQAVixPPnJXZQrAZ6SfDo4j+d0Tc
/3zU4cjGE3Kp/t3/aV+pmMZjnnqjynFA88TGHqHou6C5oRVghdVvXLx69trtSwP0sVRAWFhvwxFB
0jv/msW3atStvHLGdQYXzcIHeslc8liaIT3UbYbQEEq5waDPqKww+gu7SLAGvJhEFXEyJyIdKR+7
0cIpjIQ8o6hdl8m/pecsX8TCMhdvQu0qUIEz1HMvj93hpeGSIPN4xkJUvafnWiAwA8s2HvUlEvPf
5W04fSSWt9Ff+LvObQHhsCuYEkiFi1UBCIKnO2nxBNpu+czcrHuWErtspR+i+q4VFqVCyuHBk1Ln
4axeQsoe16WMzZ27Rm62v37/LLWCgFHM2C5IBuUZFC0oB/1wUVTkfB8dIUD0A3/gtLBAQSblAWBN
F9/aukphxU8nap9Pi0S4g4YPaR/Hz/G/21KIfrj8TA56NRajzamQq9oZhng211+J2aM5YYLyXRyG
YqR7Vv6j6z2ZxRQRZKmztRV6yZm7dlTyVhQcsXlK97U5eEOgrAuL8X0UvDIjDrMnqVSmgzquAsGe
+xQCeb7XT9lmngWRf4IWs6QfZniPcjr48sM4olebwHhWma5A0YkZVxmlpXycDZvYxLcaRpmlUVWM
0JsY8EMWsAoGSEFrJxHeMTE8ZxGTraefklaytQ2yhXB+sumCdi0OveXgC2P59LgvMJxPkRauDDgd
jkSOjkNMOfaeVhdf9jazp47VCN5jIvC1ipNdKcgjkct/7ajQFOGA2VputlrKYPUqc4fPBf8MT6bH
g9VLFkRc8P1XlhDe287WgPBiex1jkSgrrA0rNmX6Ki0PZZAs2Z8gJdrgphuur5cR1j7359sEk0WK
DfVycaSLnObJ7ySz852N3c1QoWB6NSvZM3Nihpm5Sh0wWNPBQudcQXvvkmCgU9ldBsm4wmkPzxiP
Dy8IR6xsNX2lviIU6XOnimmjLr7sv1516byLvG/yrA8SLq2XR0RkXJGrteifbnxT7UOz72qWraHV
D2YXU29fywV8CxW27v3GGd/vxqhT5xCUMExjRpUv3QX09p0bNE6mrOX8FBT/lF4rAk/kJym3jfui
L9jK+h3VxSPc1LrT/eqZWThi3VGgwhEBYVYDJFc8k7G8PkrYRflYKyDwN2eyDAmw1/9cD70vhXM/
yDezP0nXGDmupvT/gljAqBcdsUMc/XSbC1siiJRA4774i9A16F9DqTzXNtuekBQgc+uFIXJSAHJ8
QxMCeUC0fow8XrdQJH0qCfSK6yJqMNn6TnuHTLWFZmA+hmk2sbNASEy0zcLjVvuPoh3kgGm/a1fx
c42beXcdV36/hKJwPAKtd74VqKJ1QNRB9oSfEjROqDvwEA+XyQYPpjUIWtR8nAvVjlQ1eU1P7SFi
7VG5ErsnW3blTjIOJW/3kSMVigCj+ZuyNQuEXIoPuyBhSvA9JwvkgQit8FqMb0AFZxZRJOCuqNQ9
wAQGyoEuXo1mxFZLEXvkRqKGLZ6XBf+BiQnqQYUULq1JHO392KBMlr7APikHqjF6Ktp/esa0lxDy
DtBAfMXIRlM5AYYAePGZKSCniJkU6BbBTyV4WBOwskb48Sx4V/bCSOAPurjyhGqsUUwtqThxdk1Q
wDvfJqysknEHw7ZiToD/fKdvG8L+lS1Si3u/sTCWKM/5TI3dt38ih8a1coMjul4sXDECt0JxwRsb
Gwr/XO0asuEW30NNPmBzmIBHsigiNcTx+eT5Ghu18/rxhw666Zttyr/r7pAHzfk55v/YSnZ9fU3C
M3e1QuhNehnQAPh6xzPkQwpjXQsNFKvL8rGf/EGyYCBuggUMsUsjEqiQsfiLPSdsjPMLgGbnO72c
LukEhpnPag3a7NtrLYdKIw6QIM3maopbboil5B8AN83ztsCEx3fYgzhdZYjlX4TV4OBnIYEIKsr+
Pb44cpQDyMMb6ZJBMy3oczEaumnsFtcXmxsuA1iihmQXuR7uaZWo/nLIkZCPmK7IGT7NAQjNcOJk
CF6tznbP266wcaxiCU4xhQOAXaiVveZnegbxhXhMHDYRplQcG94sX3RQsCRGXp4bOJHwxmeShuXB
LW4zpAMpmH1QzbnY27Ar+g9jzKmYEIpakDmqtJnpw8GLDbSHs3QzBQvfBKRyFlPbxNaBeZ/WQa4B
1QqK4Y2qGLQv+4eHSBoXLGQXK4U58xnggPOja6Wfay/syZftwJpR52Rp0xssck3wGcpeO6J9MnSw
4KUxcJ0F6nyd3mSDb9/nWOAuvAp818a/dufZznvj17ONo980KXO4uj85yHfho3KS44FkXdafEAPi
CCR0vED2mGeJssWOwYfj7CwcASo+YaTNXGvwJ1IrZj0e4XJHWWb4ypeeQdfH7l9MOS1Z0mI0a8B3
M4CooQsS7Y+/qJGzJBXCjtO9jrSXgBv7vZwwXt7Fn5K4IqReIr2vylbnW1k5gkWU8w5LEyBJXuor
gP6R760MTyI5s/jS7O6mIwdlMh3C+MfGczqCqtpGa2q9N/zYQbQ/SmsjXiAUC+CAkSF6UkdKTACd
q4DUL+K71FN7dNKpedi/DWe5BCFEOIJEJlYGqH+FQsJA25zzPpl0Ai1vPlB1c55Z/M/3XKXFKhAj
dwnDFgLqSh/JOGgY0zpJ5xHnEBAUF5c156y7i5lWdxqEa+9P+uR+Twe/9TVWIeIPv4QtgN+b088a
mfS23BluviXiAD7n8oHQcfRm7DDqFiDWQOPpC/nNI9KdVdEn0uEF6ECQ02m9InyQiARnJWjmkSrm
WONQftvsAM9a8eYxnkVU3rnEx1ZL14uAyK6HnS7xri3PBNn+K1wQJj3VOPGCbGMJhcMVluHGuxlJ
0cmhMBZ8Pvi4T4PnYYdbb3ITJXTdoP9viOlW9FU6ZODJZAj5mga8+LKst8S78rFMla1s8yA0Z6Hs
0umwgFy7iP6MkPtH7DyId5d58fpSvlp0HgmW+JhyiFjic7q7OKnJYUwn95Nire2tDdnU4qtqAbjP
rBY9IPvLQa+CkMgpOJesmZg4y0le1v0yoHGahk4He4ST1q9Z4FgHzOONj0u3I8trwT8DuFMg1J/E
6hplq67ZoJQMobWJ/IYRNUBaQik4mszVnqdTb3XJnhy6iD786qqB1J9jZy+keoOqVojdOfOyOxrf
/J8S1Tu7ulI/Ao6ZsyhbbHxHqsUX4OQ6O/TdZSPNuntKDVCCEznJmlUN2Zlw0PNVjNTqIIf72Aic
EJJUAvnNYOvZ/14rh6TH8n03RRgcWS4JPVNAvClPtNivrRX+dBHo/pYfvrhRldhrmLOTpUmvzKTt
BnnDDBThOjsuY7LKiH1eRjDu3d5fW+942vENCPMi2vFdStT+Ykkt0B/Ku3TuL0qN1haAePZTxOpt
D0dv4W0vBx4Umry7DL9Fqs6tYX3DRxysvfBIa4/Gyd/9D5PeWuqA49KtYvfm/XnrA2zKq3lgBUof
KnqQZZWy6B+yMeDVXQdptMnbQTXwTyxv4BgQ1hzR3It4VpY1nRJpNHUkng7wbh8IilPMp310DdNq
mw6reeQ+3b7aihd8cd3r4T3yji294L5q6uilGMhaH6/kDZERclYC2PHm+kWoVuETJfuydXoW/g5W
1EnT0/XnhJj4JLeerHHMmBRcDQVOQV4OZVpq1wFDA6SFj8xwknb/yUwLNBZDklOcBMx20SpoR464
FW6IP5+TdVJLiHIaSy1vkeeAmDk1DiSYYpKGLm6ej8fjl19AvOGVBWvaQ6/wC93ZDsJj1JwjA2yi
nD/X4DdFuGKMNpHIu18DhxXweOhvL3uynTcbY2giKXlWarJd1TD97ycotAdcqbPEi/ikFUsHNU+O
cWeULp4SslQFc4qMgkLHuIbfhKhRyeA80X7177pOAIeb4rM8UWdZaA8YTRC89FDJHZ1nyULhbvJC
gF+ZPh9fPONOKCijQjKD6q2Me8D4MW74Mu5wQNEuuLvX3izTCGAMnVUOB3IcjCb221bg4HlT5Vdm
S8z26BsMJCqi1XPnJ2sbLi82LE7a7k3jG3wUZ/TzPHKqsERj/g6SgdUrN9IZGsUggxfFR9wJOzIw
g0aWFLEt1wD6V7EumUytbuQuAJX1VCpI5rklE3QQyYGAZxvev/4113F7I21WWcA/X9vcE7evUIrh
cNsfUpqbpjFu2U+ivLOhm2wDLqdBUb1YuGv5+kQIvnVjMXsPy+zFqoHVa9YxPVypAkApE9T8h2XJ
ch8nz/kaVUs7D08ffK85HlOpFHNGx6qd0u1DPbqha4akEPgiQzlkJs8sUwPe7xH4s7KKKs0vTV/Q
HKlkI326UeU5v4N7GSIJ7RPio2tkK9lFZYIbOmdE1jrs6MylCiDUxM42UQ16tRQiMhQDDc/ZnTTp
6fD85tgoJ7h+kHvrayJCFyZYx+McBxiesfRk4kjAE57A2eN0vMCEhddAUQ8+GEvil1ZOtna+8jXV
8xd9r6dmnAj004txWQUJJA9KNnsYMovmuv0N+RFcuWt+gm9+X4iwETo6+h/q2dvfYH905u5uhUTM
Bl0PhnfmOdxzED8TzNinrvnXIbzR1/9n9sDNSe/cDRzPOzMXhWR/spXOPIAj+Efqi7iHl7jgbMLE
ksBHBjbPbCG4Nj+IH+B0rRGnwaFUGErQh01bx3MdyqNAbO+zo5BNSQhz/tiduWeHlnxv0ezVjTUC
rkOrrxUy9A757STb5sIeYwBhNr2Zg13wRLcud9TRKuh6QlRrMFGVhtIsnnp9hVm0nUObOnoTZQTf
5rJTv3nC733BgkITspRD5bYxr5iM3jc8U1vnsKwBWhioS+KpPsT+k1MZFdeqt1lHFYUuxSqeyiqe
PqifNQRPJfIh5B7pdFvGrt8=
`pragma protect end_protected
