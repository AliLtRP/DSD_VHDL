// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:00 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TD/lRkYFFhJ/r+S2W9G3Z6N7FkO9pPASeN0606177XsNroRhrez0JWBspAbkrT7P
lUrOFoH4ojtaMynBIjU8yo4dfgBUqz6zMPVSSBU0GLH4CNkmqeV11+s9aQzKRNyE
D4R9YRJz4tSb6/2QAioMxBQLSoBQ5/naSd/XCqupIN8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25408)
Sok2meRs/eb7HEelA9I9wvIoCS+IqFhiLcKcWXgq8efladroRcIu9H3HwQmEMcBf
QkRQSxJNksBfxz9vmK6PC4eqprtv34BKSB8KmmQ9uxx4fnKbnCD2yv/KwhkznIe7
fi7hN/Q4f/NiZCDY8YFul5K4+jp2hyfOwBHVCnZfdq1Pjl+aHHkCjvUi325qPCec
HDB3ONFcQu9Cmh0SXacRTsYP6E58uBXSgqBLBx4HyeAPqmzPjVKwz9tpYW/+5dHV
vvhZmtQEuOtBJqF3nM2h4hC0EO3JFvBWhoioGw30QIg7Jdb46UqbV3tIL6cxRfVn
UH2x6k+tZ9zhL/88dqksDBGrKLh59NAZHnHXhSaTaCTrUtdUGsO4usJJ8xX0U0QA
Ram8f12xw1SChOup8nOMstdT7vKiD1YvKclXkNWbZCo9PvCbVt3nT0W3Y8DaWZ8S
sz4kYxEWa5GpYcUIzxVZtBj4AqDwehf9pEVVF2aRy8eVe5v5zdrX3zFmyCXEcz4I
/h26oDyDUC1z6DrkVXUZfyVlY14ccFW83+Aw2Wly5G9pzJ5K2zDN40sqtpK7AbY7
1x/VkoL3sg/k3AIhT9OTLEAQQZIXdF3lwb90A5UP6nZRq8IMU7wcPC+C2ghjDuZv
9aPhoczKUh/rCpzCRm5A5elYgvPZ8hIN9l7QimT6HtmgmpICGvkAU45tcnElYHD/
YK7aZe5vq6cE1p4upqihwg+20F/aTmTcD0qcx+MEWMszd822e5hisZPNsuwt+tWX
h4mYKGF1EhtBByGWChKEN6vBBlc6gm8/TnUr81MZtlzWQS21NDNHRY7l1/x7+kQv
hlj1dRC5NNarwMGA/vx+Xk9pKcqfrcuq/Rj4hJprd7mKxjFp9JCQ91S8NpI0EymN
SdC4uKpz2nZ3Y2oAJwnHGafJLzD0bV1QxI8ZxcOUV4BHq3U7w66k+c2n5Mte4jBw
7DEAK1nzwEzkpJ1mGGg1cNsbbUPxqVkw8RTVMC9aS/rVLtdbD8E0XMVfXlk5iNtR
EhkYpTYP0LHKhXWENA8ERqTPaTKiaa0+eeFfynccgOUNY3PDzbxlPb62SWnjBEet
0SMZPet8YjWjizc6E65qRKgAtvDfCfXCyeqIroAwQpSetKvdogWk6WyPq24sWUbC
2/lv7exWN6cCCCsB/PuXd0guPnqvZXBJNN/BFo0Hkz960cyRfSAiypnxF6TWfUxg
nx14oW5P2xYx32HuzuTJvaWeIqrTXtUkgkZkkSXhOE8w5S6co9MfSTXLQ0VcVRhK
yteQlQHqv48Bvn7TdmVHZTHc+obuA6WG/vNsz5aGMtc+X63j/OIEGKKkPtmmmV3t
z5WnQr6kdMmCF+di764Emz2+KNeIEh8ogcog4KhqnRVbbj4htjJrs2f1K0aI5LrS
8ltRyZK4uy7fvqNuVI7KAnxYls6jY6mHpB+Ozu52I0c7NiQkSVDG5+jnykMnQZVf
py9J8lhegLPbQhMKxjWQSid+GBm/m2ZeRDDb1jSH6/TZ2OXldgX3brHpU8Cl/OB8
0d4Q16iywYD1eF4CsAQSSmJpPI9DUIp4oO6bkMe/nWxP68b7wgkTtuHp9pGLlw1C
IGSyciXpMsJsekzgOfaB3kM3ggA7xJoSAQxntsd2JASXkzKtN/5OP89Ipc+DmVUd
q8XAmAbn1PHuKYQNsaO9kydASoLenRc5V0YE/MU4E3D/of9ZxEVu21NPS2x/sCz2
qn7s/RbUGHcV2TnvyqshN4uVK3NzN6Wi5Ju60p/AMQjii03KSwLJy532/XfIZHb0
a1dmF+FNzGUVhjYiU/zJDPQxLzKwvdDLdDxvweEKRvQjZ0pzzqwyHSLNlhCdkWCz
N8mxV9KrkGiieZRR5Yzo8vfA2FgLZfc+OXgDruMW0MmHkG5IOA+vC7a7c9yJeGNd
12tYMkw7BGemm47F+hovM8u//Pm2SV0m3RutlgplTPzmU70NA1F07SURgsIMEE0D
pIwplpaBM+cjK6l/dMErvcM9eCM6mqzYFLgobJGnBDRkiO9UpG/KfspnhDey2Ss2
HkYXHoo4kz1GDkpEu8w9WEq8s5UJEMrD5PAzZHtGpdwnp8CRE5xrk/dzCbDsxCxs
VIlGJvRhPSF5sIcHI3pXz67O1Wp/axiFHKReXuHDq7OSmln4glJEqE9tSZWC4G8p
7hngys5Rd7wKcCLVR4Ff+wCMN6vAHrDgCfDUGbjrzP6Ts0gvQqRmYFpFwN7YZoYT
GKWNfKGMzn5NYcPvNjiSy2Z6qCTZVzFpBsA3EleR18BQ0s49ObrVZS949S+mB3QD
91i6pZrs4f1juDnBHKSSpkFxU7M0czCVspwrrjqR5NkrHnaZma3X9OXP/xeHQ48+
4kuqPXQ2i/ugAQpyvoU3z72gCFWR1H0iFoq6Ngkyh01Ank0cvpSAdOpZ0wl9f7zb
uih++F8cE66WCXym70j8PqPHm2m3dZB8+g3ZJVx04BXtQ7eHtw5/P2a+cAaKFCGz
jmI1trHdvItPBXJGCpCv0QSl64Xawr0eY2NCby4DvZeMvKe/v/D1+LJC4On3eX2C
RNgGBmdq3vFn8BLis7uKaxAuyspP7makCN8LV6ccV8LXZASznQE5umGfSuq9We23
4FpILT3Zhr4bbyo6zCtNTPnmNL5KQxVkF0uxnAV3+FuHb/Sa3L+u9HfXl+z2kkT+
Qylkr+BpDldDWj02u2GlyaRDIb7ZnJPiEwvSzsQf3amO3PWUppyGbNi4IhoMQy+v
bYrvIyPtZrIukj9yyBoQAZXFwEizMSIh9A2R2ikde7C4Nu5FBMDoOxWxxwOcWke4
yL+ctccMbLCAMbjRiGUAi4t/ZQsAipa3CyBo4r6xWARJjXvIo36j8KifmzyzSHC0
hr/3zLib0N5K+S9xanQqUIPUu5mWOiWs6e1vhQ1ceCLwcM/V3XdgsHn5NjZEV1nJ
XKCOWYOR8MovZm/NP/SB969AhdbZD9TNsYXukeGeXbtTNjW5q7didLVvlXQD+2hO
QCFm7p9wUaMiOu1ndtZOe217joC04Eyu0GhisjAhXxoehLuadzSZUFHGiyTDu3R/
OpLwK8NLXWL52YiiKKltdYkYR2hfksF4N0auO7TN5GYW4O+8WANw6g3xn+KD7IKX
mkwN8lXzz2VicPDGoP2+LVTHF11CGjZh/yNKd0CrUUuj7nfNP88Rl10Wg67ZgRwR
Bndn0Qj8C35PPFYMj7RCuAqcixDJbjXdHEAxcVTAELB9oSXLs/KKDUTnFYTl+64B
6yJzXSmE5W+Dzrewqy1eCBkR1W6PQ0XdmwG9hik1W49srsHhjsAowoz6PZvFWWWN
BOKW8LKvqmvgmTuRFkbwYK5EzUnjyYGutKVRPpuzAoxc3FSCvCjvdh3VfqaTDrvd
1XnDXGbxkaZlO2v4hyl4gvwRzXTvDCORxcchRoAV6VHTJcjh5iR2vnOzFzTN4Ecm
QU2nk5rLhmQaHCl9G27U9ybJpdYwL4yriRlU86tnT+idHtxkHNqZKILDPkEjD8AY
x31RpFfWIesv17A1VrvU0hXR9DCgDTZP6pn98cw78RH3LCzJ1gr0WoVwgWtcJ9ey
7zhni64RwiDyXCwWNCkpePa712w0nPS9vtTxfK03IBQUSXI3d5i2FuzB1QCHqXUL
K/gt2aEs3kmxxiPXyAu49Jmfip315H668nz5tmNlQM531GB4NbTzCdzBLq06j9Wn
zwo/zQMrc5zCBw5JSox4hdFv8W7t42SyxNpA8+gby/Lr8cesWjZT/w7M2goH8zDW
+y2O5OFizilaAoc2Xw4pNNUkJ2sV/z9kdsrt28tEMNYjbVI4A4J1GFQTTtAwDLZG
VIreMDWPgWRNT/h/xa7+e4kb5hmi74hyT9+cQaNOJym+4sf+CxGRurGgYAkMKEk3
xdQqqUIN7WOILCSS14VoGEIEarxQWojWqiAuyzgmCOgSgznjTsqj7ekQ1xNVYjAs
cq34ZsJrmWy0MUaUO4REVm5PZIPJm/tP558Myp4HVDeDgCr5x9MKR+AmEQwPObzp
IZg4ojpaDNApsUiMiEypOIjtwJncVImDtt7uwhM+U09YrOI+HEnYtqoh+qbnfsat
btOFAAqO62jdxnfBlJZROx+wlqq1piWOP0ZvpuhGl/fZ+9YfSFcRQOooBaBzTPkb
pEvGkCwQaA8Ll3K+6Vepclu2HE750RrmQqTcNFCcRX5lUHV00cqp4UZ9Je9q+gTd
kgR1WFVKP7dFpN8swcMEzBWQN9ZV8j19IAEwxXzXhAoaWDaXxiuIZfmADTXQDC8X
ajUsrthCcFjvAAPEaiiO4WSDnIfdzVlwO12JqsP/hz6lDJtqnM1wDjMwwlbCeyZK
Mw8llB4JGT6np3B46PTncw1Z+CG1bQutwuu+swJ+qCj7Y38/LH/VheCr+Wo2dCT8
RifmbqCcMakeWEn66rcahFZE8VJQF569E2o4TPiDKDLxJA6ZR47X/WpBiBF7ojt7
+o5GhQW4IeP8m+piuEXn4I07YWOaVZhQwZX7n5HuFzI8rE3MZ2SrKt+W7hBannCl
hKaXgztcLLOIWr/tzleYk9eJgviRJyTnVtn9oMpVG3P2w3yJoI/NLmf9rkh/fg2O
YMBg2iiqjYQ5EdaqCprSZYxLfovfms/dgBkIKfEu2aaB23Wl2fb460CLLCajE9bU
1vOi1x4kkgXx7seqBLHa5OZcPDSF+72JXi58HvfMce3M+oBNf+BTGqO+c+KkwnIn
NNWWG3eKtmfxJwkZTaP6yKSSgh1W9cgqnhoFhoQ0anaYTP4Ho2M+LaJsBJtkzSxF
pD+0pQKp+qaTwgh7dHmrcwLvc3usVVhF01Xwa8wysM4Wnyv20xnJrX/cimHN3sYo
RZDDBxLra+TgpKV92hfS2ivQdbRFvUNp+WgEJc6SpbB5uPNaZqAjWKmbTHjucJ9p
5Tu0WZ5e3AtnuT2RXq87TKAxLecG/w/JY//hiVfRPDVEsWOl4hNXxJl+UhsEjxDZ
SaJIFiap6WJ5J7k0bZbfxDFXwTf2uOW9vmYaGbBmkNXoXCoOQQI33hiTK32TIASg
AmCkoqQsZyt+FZdv3FMCPRZ3dpP4uUE7Reu6JI36XYsyUmFUM1llBN9qm1EdqHab
F6ahGTnifKo7BdMZaXjEMmjgaNC/g3YbA5kRz8lh8XnitDcBz1b9eUYApxSCvYr4
JQvdBLa4NYDj47DT3V1GmGxArixbYqsP/gqCcohRSXJJtPzbG1UGOntLgafFW0I6
XXWURDnCP0PFQwTiCYGOD/IT/75kARdUBFR3A8qtcp/tCQVXRrUU3jANyeuHVdKw
BsjbPfBvdRjACxEwenK3Tl1boe5UqE1JHpZON8knjFZkNu+wnk7sbyA3QdWOFINp
d3oLy8pC8g4h9NoZ7U3VsUdxpcjr66G4io+vo3/nNCOPG0hC1ToVAA+4nLFS1vgD
53E29B3lZGkMqxRcoGcj8k+JM+oDbazeAc/X2Onb4iiOFWspunQSEk4X8US+AaZa
Uf2WDukJPpNk36e+3g1E6TMG65vdYdhg2bFDw9iOMaFq42obKb7iwVN7AbANEuyC
21HPxmM7BXVeyeo3R2AP1YldyGLaJsz8let4n26h6uSmNjTWZD5WH1Rq+al303Ih
ICK95bPaTI8s6e28NO64IVNG6VxHitxt2RuhRtUzFr+j4dHM7ge/w5s7UczHlnP6
ziy1kxLgMUxqJIx+NnJlP+piG3ZtdccULShhk7D8sMs/6n0G7Lq+FjucgkbiNREo
YvB3msBpiCsTbfzRNZmCe4ECkwIXFj6YympyO62sTjiqlx/gLK1X7qmo/o3tWqjG
vvQ0H4j8SUzJCf5tHkR2Pw6O5xE2mtU0Q6EP22p1nvP+K7jYuCtefx1H+RSXUe5A
7ByzkUKj2wtbCJbEYZD6tCMUbIv0fseKqKIrVklHUMhrOivPQxtSJLapSfs4IRRJ
O6p0gFOSp0Cm4bMJPUzcbpSpXRvlg2eVIsIvrLKLhNzwWNS2y24115Nxj9g+jWcr
v9JCWbETLdHcD2+HZqz97XKyXwa8kOKAl/qMjzHfAPWexNH0rtxllCpuCe2TBQ6M
kvRC6yD1JKVTQs1CV7EYK+ilx5fIaSIiTNp6OOlzjfLFGyaMxcdJEHqLlO7SbxtJ
D+9WJkK6YvU2Sz8UnVdIN9Ptxn0884Sxpksh6fGhfqZyNNRpAjSEt17J98Cnp0bI
Acrtsf+tOwNOInqbaDhoAeQ1MzujyNc97FXgV72KdvmMqM7bVpEHk3aN7LVM73ak
rrX+SMnAkTAojTHI4M80+oWmeh/N/6ML0KuVq7DoHy4D9p5WmLDCM3yT2j8CI5wP
bBGdD27n9WF1QRrXUoOWeW9Y2EgHVw6AB9Y1zf2hKQDSQAIQCt5csBE6nN8p/m54
Rc5IfrtVJfB4BN0QrpG1/8TIorQiJyqIjE+YccDNFVoa7t0ppGvWRIUpkvgLV0kt
HhMGhTT6dkGedeXo/Afnmch4eBMhkFOtwh/1xXOrYsZxEHaOGmS/TrPtWK3VgVQo
anoXP9UNzJZDYjX9bF0q26I8vJJDoCTZjU1HixxNBo8sksBN2Pw2+fdQZZ7ccmpo
mSCepwW/PPZfyo5aNm4H1MRGzCwqCKIqrAqPJw6TPJfM9E0uJblQZSdu8WIAirf1
MTI/phxDQ2H62K8YQztZ9+sDwspVIg+bN+GJ4jgFXUQLFMwP/LHCYzHHbDL5Orlt
9nKqq5ZffN+w06LT4ZCI6sbqnzUwUhbsMlavGVElzVk5BqzHrjP8MWe3KlQzcSp0
2tvWwWcuPEoDuA2lcf7FMvw2w1ZvAIi4Z1+9to7gYMBGxj2fAA/+P5nnkYtp33rT
z0k2pAePqxhNUEBTxTlTQGr/KDi16FL1/IFVd7ggCoY8ajRjzE+OnFKJb1y1w/Qg
XMuOUT+UytZADwC1bwmDDz9yQhJcW5NT1ybiwCrewdK+gG+jgXTK++EJ3tan3Rqg
nODqNnXSVSPfIbEwmJuNC6GCICsXwPYVgD4V4Gc1KtQwNU0kzoNW1KtjtIlsyovS
+zjMYJrjvscaLYQY7uecS/WX94lG2TYref1ic+5PG4CaEZZR5p75sGy4ooeHEgl2
ELU2P/iEkP+JJJjNu1Co+lZ57ZPGviD1Um/0SsptZ2c0o0Z7WT99dD4q0D/QAhOH
7m2BgV3rOuKB+RXlcoHRkhP2Uw7eQM8l6HxQ7icjARbB4cabC4wKjPBpf4JakvRK
K8I2+7HKix0K5QDdfJgtRLUUJM9Nq60KqNuGqC8UlFc8hCtuHrLLRJq6cDSDq/FJ
BXLnjYJJeeDUJ1w/wVYtkfL66AG2qiBRs2lLtTtRaceAYwaT777BukvLRRc0yxhm
MNJDgT/uJlCmAQrFz/GGKGJG+89pYJ09f5BYGmxYi1LNjC1+aSzJIu/R7Gjnj0RT
WVz9yBTYRhOcMxEWiogXYCJLJcyy3V/J2aAvctil9C1tcxnHJnxDrjfTOP4KOX5M
wSd2AFZgDPs8RQ6ijeznpxF2H/nFmpbHPWPgM39NBUKLiIy2SbisMVpb0DuWUx1T
wfsOGvBvz3tIiL/9MxIt+I6fTSJF6pKiaG3deqFC7J9vjwpNQ6YvmgBreZZocwbZ
NrSbmq8AL4Ka+KgjzFvpic/r80P2uw7hrZIUPk5l6wKRVN0u6Y3VXg3YLZ1SiySx
nxuwm4cVjOV9zxb0HFlSMDnG904R2P1eXonjrVDHT7O82WlXC5doctnSydI9UGFC
Vr4ZpEJ3syi5yEsInXqDlOYUWSH2Fo/4m9yrvb+jN9LdYQ9tdHrdLy5BnUPBuguV
XbT+6NDZDu+tdQBDm+NofSqr/71oNgKiHgc1JLvFHs9U3325SbIwTB1b+Iajb1kh
Llz2g3R9PScfyrfFzogtHFl5oEO10ntX3V/3wgL48yadN8iKNIFKNH2g6UT2gVlE
NIhonNlmZ9O6bnGWissbciyN1Dd2brMOtwQQ1M/PSTiSZP1d30/Du0WVv9DZWMfY
ZV55E9yFueZiyG420ioT9T5PyT96DlrGHCYHiZjpPVbS1zdFYjWc/lMRbvWyh3FF
rhoSQB6eBVnZwIpNTd6Ut+JO0vd6iI4Lmqq/46Cm6TcUuOBYWODHbKCOrGWzNaDn
3b3brgc8BjETzEapaEJEe093uI4yeCBdGG0M6kAatPI50wxl0rxG5kHkMQDxUZVR
0gtbrjH4cx0fK6SSodT9fKDocnivK088VIYH+Bd5IAuciXA6/cKFYKNrNWdgXcbM
Vj/Bhe9K5EjUGGjRVg9JyZC7VDoxvxynGJmG1UO1EbadHtnmHoYrpTlFaDBaZrM1
lK1eCzOxIhleC2onKQ5IQvQZZA9hkJZVtKXJPNXVGnK97fLlkbK4PTQ2V8vq4FSM
NPcv7FuIbHLNU6/unbQMUfkC4RrExf5Qcbu3SCMlXeN9WfULuZ93FgVj5lwpEe1L
cjj0bUnwZeZ1pmnvcFPNMGqmlrTPjcg+NG9OTQiOwulQi3iyJE/4sEWtcfjPSdX0
p9o9iCmS041wVE+lUfMr3cJcbfQhkrhE0RMozN4CfnEEgBKU2UYejNCcV7yI3Zst
JXDm6H/NaPWdvvW3wzPyvcDuU+lDky+Cm0g3qUy5Wz988J+GDuChQz9NMEt/MSxO
YOnZ76LCGEQFOCa1n/gzO0EyYXnwloIZEqfwoQO81lsKwHoNgDUOk9/183VAwE6W
hFhS60uCvJY4Wq9hPw8nZX9mT0LexJSYM6yov+XYDXcHlg93Z1w8pFK4ImDqHhYP
AKFqQJ8IAxopJHFm+rYZAddGHt3zXu/4jqR1hW83kYzlsuDH1COSPj8n50+ywbVN
hVkrlR1OIP7t9H03yfpFY3jFiBew82yhNCtNSUP6vw0c5zNtnigHS+T6wYywt0TT
jLX65lb0CHYbn3f2du4Qkoy5cyW+lUmj2TTWOB1GZ6/vuLVblmAdXl/eZ1DnPtRE
QM2ZNTiij7rw/m5+5C90Xq5R677iAI/fZQklUc9gYgpAkgugrY4Vq71caiwSS2fv
WgpY1OWIZzm3YRjdETLlgJYHoxmFM7fmS9u6m8nbwxXYE9sf0Ms4nUA6qKD+kZIi
NHbLUnuRJGrHKUgcQBQU/Gd+f8/j0GAszQiBcp5V/Og0IkAMu3hfxAKN6a+ndBNx
lN92aEcmqpHMi6XCkvJ9CbWuZ1GnkluISq1CRYpry96aYHU+Z1rVw0tNDsm2sxda
Qjcuyf1ciyw3fgKKHc7yxBnEChSTqBujbruaQ5nkts3WUfzdGaZp/zynnQJYicoR
484OR8DzPC546CMbEFX1WonYljfWP+faO5HVpkCEQbvqCEnudV7faU/mpgSFS+9o
dFeR7tLAqfWSYc7l4NjJWI9VFq9U0dOplCED3CIijNvKK0IToDgLfBqxzVpAHN7Q
bjP6KdU5iHccNuaY1MEDQx9s7b4HkI71ieBwnodKiYJiGskQJlLgX+N2FRIR+W4/
k8t5gxxxGhVx6JmT19cbKY1yhGIMHG+AG23phZHKEAH59oyg1Ujw/o6rSB4tYsGh
7u51RuOUnI3ACLebRE7EnX8oLRmZ13ztkBXDNJbizex+aFS6PSMonulhLDKfTL2M
eMOhXn5PoAmdCjEPd4uk7UTRCYgL5m9fLNWxYRl3bwe+TOon+i0kyhJldMX+VPN6
yU4/qxF16H7wePZHTXzJFhpizhwAcP1jPK2zTp7gwKcpPqpOT28QPn1GdPyg+1tL
Wa8BY8R/FfNkcxK545dgMwNR1MOvCjL9dEoG6v/J5gF7uN8wNNCOaxYA/w5yR4mj
7xhqR9Tr44aKXMkqgYEi2lfOiQRtJKhpy3hCzrekwCPxP/rIDOvofO1cmjdACfrf
nWOGuyHQqWyD5J2I2z7zb4SJiHD8W/BL4MvjRE6Ozl6dTkNTd7PkgSBZBfJdIuG+
DTOS8cOqvn0rDV1GSxtV2y3p43xp/mquWswLr2eXY0GkpA1YfS0Idh3OWDGx36dR
dRPkpGo852s8BKnqIUcvEPmKt7XoZgOuPaHdQqbamsBD9OnN5WMrwiOi57Dd/J1r
H/tTxkYriiVr6mdthviG2UHEKUD1PzDaxpywHVitEWhabEJstctAzlbOMnsIQVZy
VL3BfGmJ+7gyUnNxM3f7TRPCN527C8edE7/bNSC/XnvaBDMAoVNfpzAlpZME6Tfq
ow+YsdMu9EztbpIg+AlVB0bYjnIJO0T2hzbOdNH1fepixq2IGu2AvIddoKMDXi0v
89dX+9+QEznxHRbplSaj7Z7vaS0mLuHkhU8bJue4eTxJXiziLOjdDRLA8g13WDPE
vpR0PAue5KRux1uh4dYJTcHSKJDZ5ruAQ4yCFryg/VJZMcjWVs7V2pmqYp1lnB7P
IuSd0TxqmGEsf38n3bcnSs2ZveCY+8wE6uEdnsuVYtKT+BZYz23D29HXiRLesY0N
tr0MF7Q5T+YBycQ1IInUdpybmby7/y1DlJYw0hUz8w5YOV5AIUtXkb1luUyxikSD
eyIzVmqLZifOQolJQQ0fdoPBDhJsbEKZaB7yTFn2DgVLbmNXYYQF1PfUw66WGHM8
3BY1GYO0kgWAWvgsJAzexmguds2iEBoBPn7gFLIeIybFrmO6eLJjarjZaq1UjrWP
7o7XiHPGnpahIUR+JErlL+5HrOgACQ7A7YruZwnTK+N1Mcbj1bTugnvi2vNaSXNV
BuSe3rfwUz79A6jZQ+zL/I6ijilNEt0k7iFOMEQEGBo6oRj1Vt5PCk20j1f1UdUk
20lpIlHFO+8IxRi3j3ZGkKLWlM7F85EJdofdmuKfPz5pnopTND/pLNk1/1hARC5u
1bB05mlq/SsFEHeFeCF28PrbXvQh385s0U/g4WxQhoNrPyiKLLDvGKKao8DHNUYR
mObHCYUrmRzWIJUWDYw7WdFcj+bmZzA+hq2oUUx+8X5ipyIeZzFkzMCDl7nbCZQd
SlylnwRlo3UrsAplsWx6SwCU5sKzEX2sDs0giwU+bDmbuAx4FDham19BNPe+mUyc
jlgiWujVBr/ajFZytuPoGA2uc0CIWokRaPzeEZm/9ajMERZGGxBcV7h6BU1HmUqj
4rPKfEg+28j1ZfASi41ipIYwQUiuZ/g0B2pGM9zvXQn3GmbCxhWGajerWJSS05zq
aB7j4VoMVGzO57rNYjkIi+wYV2oIlGSfpslTnOEHkylPHEbjYwar9DU5YrJnZ+jF
kxlhgzsq0nVmO+tg/aVfU4dmtjACtKBerlEdDerzKB2ZqwsYXabb8brytQ86P7El
JFYQWdkLG2/W4UipjtDbZhBIWf+HlG3uNAenccztysOOaHT8B/eMe6pAhuU/BmAw
YzccYNmnsL2eZVwbXZY9DmAVIl9iYerjL6ETSB5qGdl/BYzjUeIZkF/plu3Iwp7u
z2Z9BmwM/zDgk/KCSGqBnJgcKknTveO+Tm6j29Qw9f8dIwKJhDpmi54/XoRTK3TI
BbDVQyOdwdDmoTdu51j5CpVsfVfT9HkuppEux1WAKDs7Eb8MBsHjsRUN5fviRGaU
nsf7R+GVfvMhM4dfYd5PqiONKQfDxYqJMktsc9h1tS4rYogfDfrn7jbI2KhCrlPv
xVeSAhWQQSgxs2sLgQ3X+d5zxtT6cH7Ilci1jAe77HrgGqEGFU8nuNbEfksZOkPP
Pjg3Be0znOjjh13ftWCtFO1S+4Cq8M/VJLj0SJumORLvrY/OQFkZBp/XfTS0RH4D
JkXn5iR1NN+7vk1mfHhcZXiMGhfXQlFYrE3XsBnuMg7M4dFasg9/sPVYol4cFob1
onQfI0c2UT/fkfemRVEc3Z2p4VE3ba88yjleoiH2DKkRoj3TwkQReUdjI+jMXOVH
KuB4hluBhiF95SjssNHrjK/yPhNi4Zpe9X0Uob6caOnxkCe11AsL/EcydnSPOEr9
XoyNFbhq68EmToanLKSpjLLPZHehxqld8yyKfnykwJMx9/wXYziKREbt25Z87zix
vvv+PgbmnMFmwCdaUYSfI1YHTEJY5Opclk4g9uFd7vNZkQtf1NcBLYJM9MZEBTTJ
s7ulwNi4Wx0BwyngTXcLoHYasL4+pYCQJ1ERDyS3VSVs9jMHqfZTY5h+lv+2KKZY
kDhpIIVlycSpJtDh9oBtohZJT7ewKjjMCXxCNLek+KXT+SFK+pjOGG1O44M1EDGD
5Rl1QoGtoxk8fzu0K77ER9q99Z7ReynoZ49eyuqHSCMTubr4hyDN6+98Dos/3E6S
oWUnxjTQzUTT3Jau89Bj3dS6ac1Mp7bknFDcwHLOb6Op+8BK1TeZZQwTmFR285k9
kd0qMhKyE5twWuCq38od0ZtOjKHEtcUWQgdcIVd0UaFumNaSnbbuQbOz/4xzNGBf
jfjix4iAUy3kb8hvIljy1PVmr7b3TiKs1F4IfG1cPvmQ2rhqKWeb3s7pwmUdC2Yz
yiKe8YDPhDOa5auvwymImVdDjt7ny99DSvo8q3weubgc+sHrFupbRejPE/eDL23C
jy+Jsl8PIAQeE5560Sr8WrakwBNo+TBJYE4lkjzNfd1+8Lg8WYRhW+/ErGvywJkQ
vmVN7HdwCnS1F/MJs1x9MUzBU4GOmJ+z6FNSsp9VD4X8Qm13snwc1py/Brt8FjeG
LjWphTwJQl22V4aygMHAG32BlGpMp9frdYzpR/ybcP6pw3lg//IrNEgwVRPDHU5w
GalTqOJIRJHSRDqtet7Q2wGAqq6SADeIMLSgtrAKAgBhWYgQyGBuRzmhPh+dgy98
ZW8aAS+5xS1kO/4MOpq9WRlEk8/6b4nf1O1skXZs2m7ziCNZ8DoWzoA8XRuZVDA5
4m1Yj1qf0Ktz/L0h0ESS1Z0J8n6+Mb6OI5RXdvt7q81BjDt5rR4Ieh8y2j1xTiHr
7lAqx5Q8WAxrU4uEH+4NFI9ncqL4xcIyrlKwUSm7QR3tIKS0jxZgWyUxem6Jwn52
Ehi/Otz0Ve4m63v7p7MxjGv1tZoEnhQYwUKlafa52oit2gBArRyoWuGKi4r1Lz7n
po0xDhvQ8RYzbi7zNQjmUAXbWY0tBuv6J1IC0wvSB2uC4xdik4FjTOlH6XYPbPer
amz1oeVwb07hk5bIi8066qsuX5DVns+ak5vh/EbeLbtyPPHxvDaHFyHEVUQfsFis
mFGY6EqQAYi/+dKNleHIH1N+a+Om3JACvRCkLrAz+RalF0XPJ/vZCSvTU8bYunYG
59L77r7Cyby32CNiSAiDm9raMg7iiSIdOSkPVYnyIPq0XG1RrEfYgs1pcxrJLV47
Z4mL/LJoGEX6Cqd5W7/YhgQ7yUDQjW59kyFYrkthwa2ZKVjt0NYPenc6qmsZH7Ix
jYLtKG51cmUSxuvgAbtOBd8YILi7rPPxqOZaQmjC6J23NE4mMTqYDonBlLkzKpUV
1isKv7KjXWR5FEiyjwgCL7qc9XMj9jsDxa0sDc0cjWjD7zWVCm1xO6CNoQIbPUyb
/mT2bQRNHv9BNx15g8YsQZ9UvCU95orn9OYOjh99P9ZqHm2/VToVtWntkrEj0YCg
LMGD6bDjgbI5nxU1zIp5bWCmug7SiwJgfnYCNLeK9+0KitEKax0x9FX+2O34PpVg
mzJo7y7HIg137f7YH5N7sDvjmKc0OSWyKXZZsYUMtm4CsBY4gfItEVp/uHx568tm
OoxmqqmC0QS9Ek1DvZ3GUEp5qLTY7YBxmK3ASN1l8DGZmi2dWxYkjN+grsL/1zVa
PGy7kGw+7LlCnh5XcRVXbaa3Fb+ZAI5ffnslwkPamOI6UIE0EZG07YcLXYD81h/P
Ne/x5Dj6F7cJy30cbmytzKrYAjdJv2GHapsO3yvku67IzFvdotyzjj8uuHMKWGim
W4BBXo0Ugu+WYNUmb4caGUV0ewleePhpxcJ1U3tFeMrvvFvDmrnNpCdQxuzAMU6v
bFGaA/g1CfXAXBw1R/wK7Dx0TVdol5g32zaArb/e4MoqczSPKPD4xyLLUm0xG4O/
eEDyuMS5aQX7EDUtWdTzlYnJF+gYQldrsnLAAE4cUgy8oXi+5owCJja+IKPHadkU
i51SAsAPZ4vUdFU5Tf/vUyjprIGgooXBq4paK2QoqO9DoZ6KsodN9sma6r33TPTM
tLMjdfezKW8OkOHUnkXmUp4458Bml3TMOANMD0q9BcGYxV+Yjp2t2Beewc6t9Grp
9uVRttDp5hgUGvmOOm08FcvmhpmwYAsOcbaesbvfm1xMBD4bf6N7FUIG8I1odRpk
NdccDIQEakmhc2ZpC/6UNE6KEuZ49xoGc21/7QydQ86KVap8ixiGRfLVfJPfU218
if5jYihnBISyDQWZWJQZ6Azt1VyO1lEe7hkOyv5WCTeQbfr0s+3p8hleM2Xu0/NC
+0Ys8LxD/+edUcl5tk9mY4pyJ5uDqB/+Bl2YW0r2ORqXUKGeisHewCr9QFnsefI7
hXSh47ik1A4PKBPKpcRW53rjqYttaUbY+bzPiQUf+aIO593xqpm5A7//kEuj4vSY
8TScZMc8XJbYhoeH9MxW+IqAzQvQQKOP+UagyXxsTRFPHKhIBlVkRDF+GcJ8XZml
kYz9a/JfIldGJ7bs2CjwC9BL56zJSP0LlBsKkhjqhxLqg53MIsc7cf7U8xu+mJtt
L4cqqMplsJPeRaB16wS4ked7GDhgnPIBTg6Nu8CF/hDD72vAQe+JRuJFAacHuuUI
/XzGniZpytUfyraAqLAsCNGPWKpapw2TTE4km4cjT3iiwrLw6uGxu6uyvcsUBDnC
FwcImB4MulVah4wvuZuOQOW7YHfJqBbpm8CLMuo+ZI/gMUOd/vpeQA+9BRom7fUx
eVAlHSJCd0FtgcGPcnyQ8f9GJfLxvOnmBNf9simPsvtX+DUrnhRfA0zkchkL7BFH
7sO7APTUwUqMNS8GGmvNmMDn35TyIZnD13gugo3h6A3FzqmW79xPj/D8SzsLARkL
2Bvr6GvnLZ6sxr2ou0ty67T2LoxADnYHMbMuTa2680wW0QLBDK7fobU5RWSezLQo
MgKXVh0OY/PxZSTccU8XL/Glo3I7dwC4vI/O1VbW/eq4idWOKoLLXW5ydaQF1B+G
PrG3E2lagM2PP7gtTUaL+KsLaXjrqoFQj8krpjSCoA0P/iqyKqBuaku1FYXR+8TO
rJToa1awzcR3uxFh1LOcuZVki/fqWg6gqYYlxDNBFndK9fZu03BJZ9TeEjvVn8yj
7kIzGtpwVBuKskLjO6TVFygb2pJr4DpyhWMRXgDJPCQhFbgYaZGiOgM0NCINhbF3
1y44tVIm24CtpeKaQwuhyjWVE8ka4EwGm/PtBEjUz7Ok8s2qy5lj7Hh09gEBzf9D
7z6OHrV6qRImPCM66VbEjtHkHwD7DJD2kv+n7KNnjazd5KJY6r5JPx5t3fl7rdpp
efuiaXi4bBDNGdXRtZSzKqjo/IoLqgKhUpOIwzljwHup7Ph0mgjKJv96mBRQNflX
JDCdeaxfS2a0bjPxpjgkTrT8h9CbwJ4/fq/+7OYE5GjtBF8zHv2rdwN3QTQrHGge
PQaNKVNjI9TySK/UKZcazCQgsZNh8eBjrrwzvKWQO90KfN+HZeYMX9NQbZWPksdm
3fU4qFAkYEgV0baOFYwm4V2YDZQY1cWMKlLXvzj3JN1ZGAZUsrlXarycgwqW3Hxc
5YdYUj9tdKCY8fc1TxmHDtnDc3Be+1g7Lpdlz6xmh8iD16x2+QVZkKNirJYiPD6J
vowjXWdOHj4Ub/Shi/Md97zaMs8hNQR5oAMbwUfpZDNi8TA9RDsGaF4NzB8ExZsD
o82Hx4YnU54Zrjzq4s0JMy5CT4G4kndYgVNx2tZceV8wscAdlhsZEjvJG5nGKYWG
OgmjGPX1WYy0TWYumx9CND8enhOylVHcinfC8n60COt9NoAQLn+pFEE+8otw40yc
79A83rKaYMjG0O0rKe1r/yYKwFIFC8HPAtajAZ59ez7Hv10wDoJCxtHBLW3Hy5Xz
+RSHtSZaRoYqy/J0ml4rd3CQEUI1nwxNjX42OOSnTDXt/JmcH7F55haow1NcOb+k
YlRDW2877yry8WCJ76xDh4nFRJX6/75Vgs2eP2ZP5vK169CRODR+Ih+eCcyRdHJD
+m3XgL1EOjApnqWZbG+gckS03OP87fJP+1cbZEYUCtwvI+Omc8XG4ChXpkFlbf2B
9t2pSfW3BF3BWeVjrZDeGOKkJwrFFUTenSRoL5Gt5leivkC3tuR1eX5b4EF36V1M
aO046XUHLMZfb4YJdj5Kg3Ax/jwryWEKeUhQm4wkwUbQg8h0BpqvrIJwG5RguY8G
oV9VtKd+ZrtjNAjTehYuIiw7djgqrAlGWahPRzgipbkLhZmbEAE7oFPX8It+Au9w
k+VUK8SnUtbZiWwnadlDpY4i1dxj9ILMBwdWHPRw1SkV8JBlCGAfWh7Jt+mWFaxr
Mevehz149YgBSfUQB3uq1BCCTGQ37LWPYKlJJ6nVL/lpgvW9QHPGLyPKFt4lDogx
FKWMrXW0B6CW1Ep91/8HULZbkL9ZPEyUvvspsCVqLWM4Jy9LuGz6z6XSOhoQYfCx
/OUCAg/UKOg5aj+kfN6pzWEnrap/JkSImRlgzei/ZP9pokfEBi7bI/ofS3KJqVjx
ycHzRHzgYR0NP5ck5SjlzqikN38WvC0gh6KY1TQ1nzT9gbGC7bcDZc7nYV6YUTgr
LOjiQnSlL7VqUQ87KkSBCofjJ4whTTS2/f0bwoY+dUYBizrYWtSFalgEptKowTxg
f7YbZcHZVlpUzQfsMASkBoP0EBdSh6WWrEgxBYHfLe3pJgU5aOBj9+LazsecRk0e
KxLouXHLqZWhkQgtVEhd7bNlfdYHZCcuO9vhTHEFerIYtDWKX3+uN/pBWtdbq2FH
GDuJfKtLF0JP3fhROP3pQU7uI/KmJP/5AqZhSXGE4hbZvJF/wgRRs+obnEcJGsb4
pOUsDXQdDHu3Bg0yY8T8S7d8mS0H+LDGVQQ16mwjSwYixh0eGstQyDmK+XuAzJ8R
pyBoM+CTzJXq+Vo0bixpw0SVHSwvNPR6CdXrwhoC1k8Ya2RqUHfRqSmyAiWU9QnT
Hx3/gVBmWhL5H3/H6OZHFjDOBHHcedIIWvCh7JoTlesjS+o9aAtNY6XyF5upJLwJ
FshJ5viqK++e8dKFt0AS1u6xZKhnQrZPcl8daeBPIQPDhW4vu7pEMv7jdqD0isrK
544EZuM1FJ0vwwOg9j2Voy6YOUbBnGFrJyGqskTwzOnPxpScjgBBMfeZvE5ygDb/
283yMfVuLPcui/fMOfYPOpq6TgnlhPAayRpqVhLREaXrV6FgneNViEjO3v3uVWwv
enYCEJsVqvDO+t8uPD1Q/HlFr7VokMAkZM7yrkahpwkwJD/geZaZ6+D9033CJ75w
fj/LpTcAyC8SLQPJxNLYEldm0ekIEx6Tx4FjT5tTWyNYDpWhqzwMA6mDtD6nVKSf
DaMlIywAeq2J+M3r4Y/AV9JntVHdnFtDNEcyB/ueWk9//ZRdJdfPMweosTIbiCWO
QqWznu1yOyRURSYXLujxlfINYXL3v8yYHQEsfNx8xyhn2RhrlYw0Bz+SzKWVmSi4
EDriPD33e9sV41GkOH3Mf9qmC7l6AHbHtBAnGfXsZavWlN12hWNZgv1pCztWk2Ji
OnZn4HIJfGVo2JXOzVuTbQqhJ593KW2XOfQCCV9G8nQDblJWyDnLvTS4vDNAZ+Sv
Hit+IwotzeJr4wumhEixtBmCCeJjrCYuWoR63l1qguF3kKh+37m1uEPhmS7wlQLQ
2JfGtudE/SJCfLeO1S8y9RMFCfV+EWx7hH5Kw4+WEbQ++JWDvAheMu0cZ3uOl5+m
S/JY9q+5aitwu4vbfhTyO8v4EQz2iTly5gqazlYHqtD3rzgkFkj5A9hL/D57Q+C8
GIRmbr/kHMCzW0xhERX9AcYZo3bYuvdD6sUsNqZlukMzyLYV5jbxUHsm4C3r/xRu
ciJMA6lJekRAwibMqYPie8sNHyyALXwfqqBXPKmADin4a9mdHxkoPDYxpunTHf71
iw3RdhxOuh7i0SbALhQhJs8hB9w66h4rt3Xt4etW1o4S/xaZxuiFdDlj/TYoFkxU
fSKuiFdO66+f6yQAaEVhlItEHXFhPCFvcufXwZFWMMx2+7D6yVqSnWkS3MLCSGmF
zwPCZ7dxXNrBDkczXoVIjwmRjGRaKW1ErYB5thGOCTHBLPpxvF/7uN5PDb0ZFA9t
oycm0pzyThs/ZnxHx2kpmdEvW9NqXyGctB1woqqcYT1M2CqdI8cz5gioXT0QF0T5
yBugDY6TkdtDVFkgoXLoyTbKxdmXa1naZCZ0a0XoSCR2P9uaoEUeookUel5NoDTc
R3pQiKVdpC4U355APrXxdy14tu2Sg8jRhjWFcup+oLyl137KIuXSX3+2Az8Iznjq
ZaY/FMC9D48NjR3g+JRv1YK79zb1+5fsPx8/KkXHPaEBwxlMgjEiTY/aRkJTuiYg
iR1hDuoI2uKVsSwnDJ2MFu3cBHcDyBdwQEN6Z0SdhkGfqobOkMdNCFKrjZHcsNmg
3mQw53hr3wbwGepxmAdU8C5J59y6L9W09LHzO20aVQxgKFtUIH8o9yF6JLHNCNFX
1R8HeP9srZAbZtSYJj+8CMan8uF5oH6qHYO7Z+qRC+l0stEmHu23FlLE80Ladd15
IYrGWSR2y6x2HuCSLgao+cZUU5AdDIHqVSw5CidROyp1YRS9+QdFvQThtWWvMLZn
YNfPmfkT/S8qxceM60HWQv7Gx3xHGm92ZHT+h9Y7xnbfIwhbkmGgTPlnM87gbDe/
leX3MNAxiBZ6nfbErqaRSFPTqabH9hhFBDsURrHQr2bWlhihNIvISprH2chRLd0z
wCJR56NMx+HAvGh4wyXm2JWyJFTPTgoPbJ3sNC4N17pzTjooOMOfn8nsW5GtI62b
m+KsusvNhbQwXTi0CBBet3Am2R/d/3Lnmg9SD7h071rvaIfd2/8lxjudTMQaC16m
NLAF33sKU9GwA9C7uiIrJQVXmdO9sTK8fbClLKMvXqP2JfugK8eNqusfbyXJ8pAZ
TY4yyvn7SHddLfPW772JllG+V46MPBOF99acdNUaLzItZfXj1K+0SpHB/A56Nrdb
d9QVEQmZyUeKAbktlHgqjQGq2jDYHLIW9OGJd1JV837vDBjKXz0IwG0aeafLQQLm
5xgMYkmVINAIJNZ0QOe768R/ZNKyzk1C7wPIz29h95bEdF5A2UhHcMdrU+IpZmD5
/SCrkZmlPpsKeEfLJ7kZJ0e0PviBBi3XOvhhA46pGsRqI78TuIaIexpzN08lksDz
9/ThB+Mkb5xZGiBBvf2P6Ls+1i5atb+Mh4fLPJpLLGL6uWq4wqnSScHDomAYbVMn
QH4d6osnMuhV7gSJ0cny3gVhYFIFo7ngWjtEM1YeV2StVZMS7wQH/1iWqgXtI9i1
6rRMNnaJLUUah/3/BlO2qFTxVuakBmcBpGa5bzumo8cCrh1zRuhF5SjtyuGrgTim
8l9VT81P/vYdIOLnfRYfDqZjzkYovnP/k7fBN3UW9NsWCp7KEGRbIcQwaOIyteYN
3H3gDHJKQQ4VIBQZmdX9CfH1+4CzaXP3Qrn+97977WxZUHsoF59wRE12yzllTgAr
lrZRLYgzuwZ/IU1KcLasr3p/HLQ5ueQL0zBbyyA3qMvA7yMDMDDgzUd4GGcuZZ1j
lPeor7g7mm08bbdog5pIGJiMByPRXJxTpiQQy4P+mrrOwVzoRMLkgFCm0CPXzDKw
a9cOOFcv8aziUVePjMoCcLed7zR+dqdHXZ7NLL3P/VwU3Nx02B8bXHVi3wieW7e5
hrFmoAEdFuWsmRBJwTiNO+hgHpoCI+WCBAznKON3Xcgrfu8kFRnZ7LoXckOSS2CN
eZsZaPSanYfBx0JSA5n+R19AdZ6WaqaMsDxoGcXEkU03nlL8ezrm9ZoRsxHA6Tdi
EscE9fdfDgwUEbsq9k4/YpPCgO8hD+ZIFDu7/HWOOeAzta+eac6oSVzCsGJ1LGo3
Efm4DY5NF5TlwLkyt8BSwQDuRW4ui6xLU2RmBJ1Z+YqHbqA7IxUbqeS0+jYa4Bi2
KGYVZ5p7M86OtCLQHFdKzodYSpmJLc9K8+6VdsZM3/CnKiUljjrsyQINz8k36DeV
g/3h7LMjIOLprO7lBrqi8ExBCZhwj/Chhqmnz8kuorcbNYRLDzaYks0QHm2fgz1k
lFvAZA2PPE0kQsqt4BoWZMf6fCtbFd8u6qD8wVPoXZzTgV81FTOgODVGLMSVXyS8
L/1xxPDNXz0in2juAcqLy8avKm+A5yZZ3u81TPgovrFeCMy3dIMvjxO8ujBg25YQ
zQRV+AD3ZIn2v4iARVUYmsUrnSe2Tt15/L1DHM+tyghYTz9LrHgNJg9eqBffQ/d1
XcCC+/YZWxHbL+haMAdJsEYqq7aMfzrx/Ya9mPt9w55JG+koGY6VX+VyoVbGOPSt
+Wql/W0okllq5fRsK0vRoY+rNBi6qSFRLErj8PMwOuFYpfenCia7pZSdT+j/KAmg
8egPu8CWsfLElGAMIBy4YoUdQUmYDtZMFanMyHeJORMafuNbycwgPnFXUWLnNqBM
92WlVA6dGUfRaFo0xFdjF/L/ZY5y45rVt2r2AC3KcH4faEdPHwBxUunpVvo4JS+N
oqEj+zo5Glu9IcjK3t2jYHSq+G7SxY74KuPO7LmswgSJWZRlGlBWhDQ1mU0ZQWi/
wtbUGJdvAmah2cxsp5q2pj/7LXuoSg2WQqvvKyW5+O6s++ViMhC2csCfiScJNg6z
NP/yEeYXJQ9ocBGatcIEDR9bu4v97J4JXocdIMmLlP8OEUeUOzMDg/9tPH8AhHem
DGp4EU+oeJS6+eVduYx/8bZm71V+svbh6bhuhEfrZZUoqlm0THa3ibmZdSnQEqxS
RxUvhtVR4hVZz7iDVtH92HZS7OpNyGuZppxS4NvxGJrtzXxIONoAhwGVo93fIs5O
aK/SbJoK0vQ5BrF0bNVhVT6NpiKCR76MRK4Kvc3QiEL83yIazDvoVI3pr1VQtzMh
9thvSXx1E1VhPyZ01n9kFAZYRZZs8QZoCG1eDf/MFJ1cSVQrDAEqZtCarjwFMDbg
JHm8VP7+EScWwSY6YOxomC18Bm+OQdGtbXFutwWcXT1EnLa+A6SX0D6bSr7HeWaQ
2tlbLuf9f9UsLScSG+g79odjtISYRQ1xWeO9IvkavjIv6X1zU8Hw3vLpjFiLFknD
ELMfbkRnKLbqkNA3iwUR6SLRgO/Sa4c5w77Twfv1mH9Vp5m4R6cdLdd2tLwawP6a
8M3/kfNXr6p2C6fSzECgbjSwbsFnkU2kfZ9M0cT5vs6Au6y6RNnBSuMOY8VY8vgI
O9NU9l7JR+AK14OOp8L70gn0V6Jq5nX4cWdNMn3H+EYbrLxo+iDQxni+SLJ2zIJQ
Fe1MgJDvE/IP2PO56lACWcXw7SSUWqcVYlDuCPx7MPNxfKbOTIDhYeOEhTOXPDt7
YJ7zIXqs4GPY8B+2oyykfTpmRObt/3W2u7DgswOcGnDuOIZcPl6fzcpgnsVjMeYv
IILE230VLfWCabaiHtupOTue1Zja2/9fpUJMpV4Uyk+0IjZ5mO0bERS/YXavvQ4l
vy2znc/vfDlsMbm21C/cTSnMOIZp8Wxk7kwf4VzNov7SlkcFx2xiiuROePWsymQL
PZ45xGo3qavLTaRIs8zVAFF14xu++ztsoN2QAG+Ov02/9Sy4ZbIIEvlZ9oLqXxKz
Zx5s1yVyHTUwy/reXO6bIZs42p4QN93m3pSTVAbWFJdk+l/Zg1xJlOXnfCjL6ce6
LTfCV+ZBeJG7PqdXZMRjdOEgjKj0+dPoV/oST11rPEujv89JOgtabzC57xDbkRpL
mRyqUujtxxeHVJjTGdM9BlJs7EJh5lwHnSBEiTnCjdzKIx+xvMc4SKka0r080du4
ddE2jTpRMXCPM2BxA6CIJQ7JpmYO6M5vju7nZoxDCsKUFv6fudSaS8WmCQ5MKu/0
AjPofwisztpe1XXRiofI2AyMD0Bk13ng2q4RKuWpDyesrgWxYv1P5vzOvnZ7VKTF
zW+sqL5u+vzx8wuZHJtzoQk92QUUda42223tMbBKMcyAnAw5Y6ecQ040vVg0EUic
YdJMI/0Jk6MfrMRoA8mNyywwU6MbcpwsXhYuuq7mAeWgxrl3F6Sw0JdAsPCFkU28
482H11nF7Xei2ATUmQlqe8qQdlIranY1gaerCvawtbz9VoFpCYqAteEJcTn09CBJ
Ip4Lih8faXIi2xCKdjAdPasLq3YJp+J74cfjDSZGeEcd7FZnwsoKdPFdMU9dd/2X
vxLXUUfGqlDqspXrEI6kclx7ktCy3s2YsbdStA02PbbA8GFaa82pf/P7nr5xWyaH
+v5mirBgeeNxCclQQI8ZWHpLMzyfhurHQa/YqBFt8xvRGdXfOnhMk6EGaJK4UizN
dIkHJ2UL2g0dLlSOXjvQ3yeNQNAwLpGJcKLm5HtgmHid7pLjNq3UeQvLgmHWSMVf
Z0NPt0KQnm9rSrfHUWvwLiev1DpOqRAi8s+UE/lqnBG/QdJWkDItmA1bGNl/5Cuo
3jbfbbkJGxdFvJu6uhWVcBz+ly56Jg0TJHO1HvIDDo+larKKR8K3PCrodoavqYI7
vXF9d+x7kpSqgQG+dGZNGU+Os8lRVw5cjyUleUj+CKWfYMJ+IfBrjtJuyRa5ZC7E
JgWDUIAPZST2zJJ3ZJnXVsO0r0cv+WxNkTveN0yzTnwkhsFYF5vFJb09wGmYsuJ6
hFgHqHhywpmzeuCxer/IX0n/2mVyq9AdPimSHquf04o6gzMTc63LJkrDueXtvZZV
VtzTUQAYiTwGIsNlVl458+YK80b+iJsXg3Cum9jRTp/9h76IaoPscisdoROYF1yL
leJVgcFHOJHP2wvTSTA8XriMvFghrh494LzSlWLGDRF3Hy3ulvQPlPnMkxbiltV/
Dj1IP1+K5QqepYDP7dDUh7oD0QXGUsItBx4X5K5nwlhGr1Q2xl5o/6mpSqSzUWM8
JaPj2M9oUaJwOu/p0exEbySYIYLGJFNG7/SnjHF8xDMthHWZSfERi1EDqZq9Lwi0
6eyncD7QAeyjrB4fUecpLw8KX8idZDeDpwnkl5vsYmXsG4euWwn7jzQeINcpoq30
xkRZcJAttdUQwNmx7BcbB8uGoM6/uoXEqGJwkK+GdmkvcSQUv3edfuQcbvW/gpJg
2EWKSj6gqzBN1izQA/f9CEcx93t4x3JNsU76QPmgTFIMRqrWcoH5Ub8yucEqsGtk
5g8p7ijA8llO+doCRqvLXFKdImJ7ug/G9uw6fGkM9JL3fWpJHuLPv6SC2I2Sivdb
CAsHDmlqrK5XAPAKeyTcxCoB3aWWZDHJumEnKRKY+5g9EQT8zJVdfvImRGQ3RgPc
tm2SggkFawmL0/zN+NrSyMMA/ZyitYun6zRn9wTbdcAsZmGRmUoIIy+EMdWGvBM8
Xya5loaiH78p7KswnMG56MszWN6zxKk9uW3Z4mv4N70vjyNlAwBf3l6M8LwNXV2m
wDVBaDnw2sO2KPpISQI5Gr3XwhVMux8/X17oQ2xC2BPmkHpJ4yN7agjvthVwNB+4
wxnHMDONlXAN8z7ugIcuQiIFMxKriSWfDycdS4UBWLozy/XT1YuZ01ETxh+Yb5A1
v6WQiELUvEQQyAMzMHZGFu0kcBvfnC/odZqXi/lIxQIeYLroGktSXp/duWgrMdGz
v+wjkf880Q71LijgxMBClh+vuDXAAbA2s7Y/LO6eK1fw0LecoEa4EG1sIDyaeArj
zj/k5MvbYwqKjLD3wY0VM4D8bbZTFxWRNEUg7a2Wi+ZDZdJlyKtShp2qB9SgiFVg
SQRyjy4NdyAKbITtzm5D47fL4fkI/hOtzEtl4cvL7vF3COUIhcwWOweGr/5dFsJg
QhPc6KMPoVrDhHLgrJff1Pts92cGPOPCc7MxUSiAykb2hIQn2GP60Q+gaMzw6zlc
BfIuEyphcgbvXt3P8u/nPyz4dU+w/bvcwb+MaI9VY4WoZNNGq40aIkTcyrMAiWiE
SCCw7HSo0uBIAPomgaLkeXM3Ug3gAxtDPEd84F+qVFIQZU4jz7TfIbwQyKrVNodU
MvHaSToXBAygWnn19kjOYM2lymm7Uibl35w/K7P+TCjVHne8zEodDg32RQVdt1ZA
ygXoRTHN2zK1KaZIIRaSiQZGxm0h4kDuwVaJpQ9tVIUiDebrijDVPhxR4CO3269i
eJItn9+dV3JO/t7iU1PwVi4i+E5VXAKL87r7gre/u28WdecIBTafnpjOc1JGuDnC
izsp4pxjxge/PldbikvXEzq3EexfUAZGfsOtKP1Z+moxFAIv239r5mgryUcXR5GP
iBk2gb5e+QmTxNbFSaT95Ac5MYtCnjHEQjvMrAH9jIBOlyYxeCF9M/IbWD22XIpU
aaBC020PvZnlNyDQYGuVGSSbgT8QIELzPo99Bmnas9rxaU5pM6CiDqaTTjCKqq0s
Diuq55Fmx11XlMG/bTYdPcQg1COhyKiEK3MFpJpJet8jQB5nG3Qqgi3Fd5N4P0Mj
Zp3WCIzegV3JJCflZn8ahCWLs9bFafCQNnMQZeAVLGQtkNHFB3T2Y8h9S0Ru29vc
SHs9+VAWzisbuwMj65bo7YDBxaGYSfu0VI0GN1U+DColA2a5QhygO6oPDoLOCZ0U
hxl9zQMz8RbSiYNxsVp6TkwERCRd84++RwyTFfE/a0PTm1aLgq8VGWTlWcEPCaQx
TUGFRvkzsj/ZyCttXc23TgYmHDfP/J8gs5S156UrGuXqrexeGGj3AFp75YxfkNXO
oq09V5kwiU9Yrnu7MOQ2EPL9o5bO4Wk/YozUNHef8lZ+1PGDbyWvXaHNUjzBsbyR
lgNyOxNCY/ry98qwdwLAx3oPCjuSzVSLqkBHjI7ulEBx29QKdrcKXtzAsJ5VraVL
1OzDA9tUhDIotaSrzGc8Rl4IgOFdwxjT5j8J8BHC5DxNSaghn8G6z4E8Y6/9x014
bIQ5DjSQYAG3yPZ7d6bckPDlyFegZWe7lFWdLM9WQcDNkpFlpEqg3s8FFAIxnqWo
1lcWEfM4fQvKUghouOrNg4whGb5Tboy84uQV5ysG/aOA0NMVlSYQkWXL1zz2LeqV
zSzByxHfUXdw6klBWefxqgRKpYgFVkEbwSNWcjfcPw5UN7NWAKegJ+DeL6c/7sPt
HdyG45HnuPLUntBPBDz5VW0FZrK1twON5PULOGpJvVdgDgCIXD/tHO2uMCjaNTOx
YqVKFDl5KVB+k5XlA0ijrJKoVLeLMQ/AKxtPkFYBOgtTOrKwOMIsDqJb4wPyFYPq
B99QdkCHHiU6Rybzm2HsQXbZtt6FjMoNZ/d21KpFVjLSpYognYPyOIzwkVWMHZBe
cfvQB7RUKxEz0SnS5Y/m34O+M21zqDiBcOZiMbl0DLKWDi7czWWULtYSRhPsc/Lz
7ireDKCJ9iYxssu3cIwqmajBBr9RM2dMoqdGTHF7Pf6GpEfI8l0YsfcwgHQQ52lr
gl2+fna+cIGOHm8gLO5rg4qS8f4Cqlc7fhpHs5h2euv0Gk0PFrhi7+lQdUR4Q3O/
4OrLvCifkui2vKsE48TnapBFduWAq7KjJATzEqZ27ASCZcw8iRHPFNcOsR52CdZW
RV7x+Lz6rnAqeTQwH55CUTZiAR4FXVUR70kQtWBI/So60HgTcJTPDoedn9ZOUOiH
1epXip2uoJ0GlNHp+h3b+9Zpv73nG7cUM0o2vSy9lqobLvJKq9Yi3bxh3Re3b04O
5hPSft5BX6LH/Yybnm+MAMJkyMcFTND4YEkGw9/8VWOsz+HhS0ukeGj76Swt+Iyd
N0XuWgoqtaQUqld4DIfoGsPWypfaoSfYSVJfDClcRM2MGIixopfUJXLn3YIideAJ
S8Nw0uXB5Arp+uiDmjY5pGuZBlXLZfm7Iz/62u0ig502ZT2uhZ+KokqtuvOmnJui
EsDxfxqQ59c3Bzi9WIoKUyrivXvvcC9+cMB9NpyuGC+o78huRRnG6lhkvODrFd7r
zltEFgyee23QNSSEk7w3WEUi+nxhoXI+81hDM8E860EIUxHyvrBV2sdW3wBcC4aN
7Uuu87B+L699P5kvUFa7BJ3pecj0IDivhETmzDijPTdOcvr6nyVroQOc84ocvd0s
mlrccCOS3OfBQlhnit19rWCOOBUq7Xw/fSSyWpGxFwfG85QJxklOsN5jrldFSDdR
zLn5pPiHu5oCuG0NaHfO29BgLW+YpsgBwiM+So0VrtE91O322GnXu07G6Cxj0TbT
iNXkZ7CKn7JA8DCocRLMEK6iaX/D4IH/6RQYwSDWRNuKMyJS1g4dPiUU+tRDBNJa
m0El4yqo/Ul99KskJHQLfSJBVOlXQZMQvTViTJq3dv6+znA3S2Qtt0YX61ReIyLq
aARQERYQ0+aeVD0RBrR5IInTGZksQJctcH5hOpU0MYReFdiE2iVjGTO2pu8J06Bb
PQpt0z6PspQQnA17VHoz63jK7Lmnf7uv/VDxRXgFkeEN+mXbmFX3G3RCe189tkTY
koeJvMPtXc3oFgug/AAxW7zslemg2Fl6qkp5unp2j8So0jP5Ad+Ha7zi6Lzc0+PA
xmB+Yit6JnFCs1X+Kx5mpA4X6C7NRTlswXpQaPwiQ5WVFRtu2/ixdeEbM6+mFnTC
jVA9oHjD45phx1ecjLESu7x+X5VCxBk95MfFwnSEkv+1lUSffgVIKoUxVMaxhxwb
BERh9kjpHpjkq+8exu0G8CbfPP+A+ukri8XsQFoFVz3uxJjRcVsJfqV/grmCB68b
V2jTAjzoAg+MRnCwjOL7j6Y8Ybsyv71fLbAxIjIJ77dFNKK8XZye0q2bmdy9h97S
9fjKOX2Vvmsj3ClkNJrRmfrLAWoK7ag51XElV9hMlG+aH/fY1ySK6uh1P1tPB+kD
YmB+Q46K67x86t9c6j8kuqWPwGrROyHYfSfOeLel78ZbKjhGAm9DHWmqHP/Tbc0Y
lKlmUE6yIPRUNie2T5sted1u2eKGNs0x+FxtBJjG8oY9hODfn1PljPI1i7Bm/nbV
imPSs/Ums+G0/P8xIUbG37LpTR5cDwavfpOqJNh44Ypc41HlqP0qVP5TbxQxHEEE
z4gl+5jmtdqLrzrcBotuAaONUr2viNgTjTvPDpYQoV+XmTsRMQjrzYngTifAIXNx
ypovCRzjFAiqefJqBJShZPT1TmgA8Injxzk1eBA+zFZruKAv3wVD5XvYZi+wVZcE
Lu15XIzyDmpg5XSxKL38mC9baANu7Sc3TTP6YCbclJLXIWW0sf267iu4VfohhkgC
A+P5xWsLTDHnB3Vs75wKfWLdaPjnkHI2fE6mEuRtUNGf4IiCsOd1AcAYxZ+Cebgn
NZqJaKiexCeGCJiWR1lfPHm23eB3iAMU3+INNrJCbNSMVKQYcFe6VJPmVsMdj8h5
IJLXe3tHMrrp76gmM+S0+APwKB8BFeXMalUE/vUecP4b8JpF+/0N/9OyHH4ok/Jk
AGPWVIAyltrzj/Ioj84oK+6vf38t1AH+mDagx/FBIUjA4WY8Ov6wXo1sGnnQ9Nqi
hpewYSysVonQneRVmTzoy4Jr4KdIz9My2FnKFzylULRNrgYkwAFeZcOLpMaSpqyw
tQP31ssWewHvK9Fo4iirwegbcUyGMN9VkNq+/LVmt0eVmS0cW0GSZRPPtASfEyOF
ASLYtPzfRA4OnJ7xQBqVM4reWdNoEQ7MeDB3QTLFUyS5onFmMx+fgShb73eFF/Is
kx5zAObR30E/mfEx8AF5Bm8t3epXL1C15V+pQtHZsNMWYEHjUaSC1QEV3GQy2DML
NpvPh+7Lb4ZHG10+If+InyyhKk+ltAtPTSBNljMFf7m98L04qyYC8bC7Hwi5lDlR
IKtzf7hEOW4MLN4i6L54Jd51XkjFSCKqHdEo7QuxWiyNX3QbFG9+PLSn86dF7Il6
0rAw5gTlLNLGCJ8LyBu5Bgw54TzmFn9myXu2wL86XXQiGN1hUu4K4RTRjOr9EjN/
i5CUItJbdaTw5WSzxk3AlmqWXZHIBYsWiO4u/DUieIY5R1mGDU3Ns8EYAuANOql7
Hux8inJOWM5vHe02uvDMvN4U4p8+IO5MAAG4dbT2MX6gTm0rncfpxrOV846bSeWa
n8s9EGpy37a7RMcVdUU8g22lFjtos+pqvHukECPxOFfISClEhY+hwMawCnl7J35N
QQcAASSBJoc0EDEDdNoAwGJoPlW+ZEtbU5YkumMsBlonIeuKaQJNg4HQsqyPi1AU
QUvv+aSrxorxw1lIWWYSrIjiXqGi4vDX49b3E3PKnKUn0j6IPHESw2GjOtT2u7Bh
JhmvMa3XSDCCCKl8MSJA6CHT8lD7zYGN+iWkc0jtJNgOzHPsYP9L6ncA88+MvOBI
iiQqkkjlruD2AZeOEHdswggoM7uUV0NRuRSCs0l0wz3TnM19p7wqw96YW8lxiGJ6
3EjZHNldQkROwGLRVpWEA3xMTgk/2s73tUKq73uUVy7Y97N8Dz+B3IpH8C/YdGfJ
maLWl+oqGQgQ1K4sG1Xzh2sck8RTwJe0EYWmJxcYGPXWoE+oatZ9bl8+tnUPXaBQ
cZEsYrXPOO7M/nNDCLoqI43YZNtvQZj99fR1QM4xxgNADQIe4DC/Azi5JdPMuxof
omxItKKZW739fCgcqHXPn+UW3CUEZXjaRrwL75esLobFcq8MCc4gZaffx+ooa+Bf
3Grr5QLRxdAiS6s5AHM06GHbgh6h66IHKd7l3mpabOvzQ/HgL2yX3qqfaYMR05cF
F+MVc4+rx/txSVTnyq/bDsLRZh1tBhFe+rBFMrzPdcDFz+aqT2Itxv1Nt7rd4Ia7
7iF39AojVGzDDvGusdzIrpxcOTEWVnO44NYkVU5D936RnsQGWtBjHWBdYbRLB3Uf
D5WrDJkgd9F/ypC3zpw0wO60AMxx5RT57xI+/RK4O1j8n2OqbEsjmqaxP9NEQtHF
vkzhD9ZcoAj+HTofAj79aeN1YC8qUopWGWCcnaAZDXW8UX7wrCvW69Lk70zL3+Qd
bkJb/P/QI5DrGN05121+pPRsoxp3G3uC+K3NXE9gOVBTTVIdfXCZrA+wjdSi/DWK
RK0I2mFr8IyBCdWcJAKrCXpyWcMMR3BHh40MXA6Sh9K6qUCtAwq7UWfl0gZfLubd
6+Wtnd/0MXoPtnvQRt/tjBzZU2l9V08/ZIL558ZmMQvbWquhTxiMma6PzhB4Gi8n
dIFL4F1aBK7F27jgu1w0sNG1MR0DUgqDhG4tgIjhkecXaOTstC1J1YJQozNcZqXA
psCv97GRRwHHpn3RA8lROO6rm/2lIYSY/p07OLwxuG9clNOpjxdFy1jWmlzwq1ya
xfupaFrAgPOWvtqmzGv100aYuLQSGPhzs3RM1d2roXDuPBuUoYu4JpK77btYhIvC
Z4PzgRJ1Yp5nT+81kq7XtnwwUk0R9Iqr4paUiGiZU6lTL6yDy+Xajl2zdxO+0w5G
R0FruCM34wTYhJal8n/XXwOgxXy3O6ZRbuwMU+/nc3nUPur6xUcvaJ02bY9eaIGW
zm1EFmtM33WLt4jDvSeoYXN+eNysLr7ynMqNFwOI6rHX0RI/nfSXpBv+68xOLv8c
VvkGNlEiC7e3P2WxNI/Yd8+aYe6vHMjG1HrXiVGGCbwQ9CfYuipcO6X8+pESa/6G
wOWoE2DWogvlJaWOvm5yZ+60Iv5AfHkxVsvPm/33+pRq+zf5sWlYMH6FpfFyz+et
rd10TY9xsuJeolP7y2pFbfQSZPQQjxiFQOgr4pj7U0Y92PhKEpiGm9zzr86h7LBT
73HmKZkSI0VWR+5p9DW/Im/Dleqbse7DLvi7/1g76y7M7B/pKFP1Bh5mn5eLZD3L
WYex6fUSVYq+q00Ih6MkMNTGUyrG4sUX+ZlA3KKJbuBTnKQQ3LhYJkk5j7n2w/VN
BS5yztpzjScewg4yRft74DXXgouUtAjdDAFfO0cSsR+WIG6qIOLHpIM1jBEnrOiR
zTDfrkMdPtNtC5b7MmUj55a+a15o++7UCRbAuaqQsQrtXWhMDIswgk2UUrI78RcG
jWEeZjfG4DWgYA9ZWwy+3BQ8o/qc4hImPa6L7Y6LH9uhGubP6Z/bVXb6V70liXkL
J2BAmwviPe613ciWkHmz615DgCIx//Mh1Nf60P5IBdOAQpiC1R2GNJJzm6o7fagq
23lDIf5CrywVAlQS1eZoFofALAOWYDcpEMpfgDw/3/ll92o2QctzozWIn7lTNCc1
10N/yyxNJqFLf9DgK7FoZdHYSsu4qxscySyxFjSWMhpUo6UFPAIOU0pJgwKPg4rk
hSUoPmQ3hM/eg+y+gzO+nrq+2MJYlS9zv7it7Ri6CI07LpQNGGDCqZgHu6YGD3ta
4qCMKPQfiLdxJFYIVFhNqV2bFOnOeW2+MBqorItrsR4goS4Lg2ryJ5DPBZWMq09N
ACbDJ9PCduwKQ9lKyvoW5svvZhE7+9zbC0MKJ3oRhjOqXxQqeqPHaFNf07NDu6hT
ekKXlwtB8esaryLKgz7qP7CfvLLqJTPIb3LNIDB3h3tSFDBPku0VUIHASCkORF52
fTdwbRwkkSeD25nFDGi9S3UUigAKeHXCDc7UrmcWEUaC4+9mMRPREfhnLNJzCBsX
DoPRFk3PJ/B/dEXVn8/FrxV8mbtre2HKy3ga/tYA4Z/zXeUx/sY41X0Jdkewr/C9
Gb8WNWqHcwaGhqHijyRv8uKx7rGvQYgxffoBIabDS+RSSrjES3uN9x+gxZYEmyjk
Tjooi8wtr6xHoRLZK6IVaNkFK0wuTlQrP1JV54PaU6rhwSldilMFQBQcSk2ARst7
3ZlEW3NlnQFgpZ6mmX1RVpK50hVsM9/yytd8tkOGMmTCQ3g5dqH8PXXPCevbYxsK
zduKKOo8ia/qbV9bSiyu2nVQosUwBAGf3UeHvUr2wRk9qVwSoT7TMvkTXLZt/re0
13SZndKEgwEgODfvGTxaPaGaRNA0y0tGqeoM6Q736lDI5rpSbmuxmQKZSvzc/oUL
FxbJPo4EHlt50Zb/K/VH7fLQfSeq5KhdpMd8ivD6cP6r6VxwUTR3liw5fwMFm7Db
V9IW0DNil0//YKb9l6Phlogvviz2OXrs9TuFRsquG/41G2bNCkhkV7F3Pgzpyvo4
7zI39MyfOxs0uoeksM9MSJ30r5yj9kpn8t05d5FhlFPoYVPzQ5K1nLjEfSSyDVB8
VS4fO5qB64imzHip250G23dqg6YJhBZiDzpi0Sv7PqM15W3nTxabaz44Ajmk+JE0
3f1mvkRIaUZqbQ7IqX0zfnRLkO96mb2FqgCcPLDZ73ho3Och2z0PTTrigoGP1Xb/
5WiTw2tWwdIDZD0wUnc+3Wtd8CZCTkcQJPwsXWWQmJjgUIOnYnCLJxGql18jOtkU
XOtfYXPEtL2lDpNZp+hXubQNwaUI0UhVXVm/CcKYV9OCRLzOIr6HZ66Wu12nfqP2
4Vm6HBEs+TrruunR5asxfnekv3qWB5lzL8M3Xftos0uOCnHMv4N+Z8kDtC972y2Q
TQcF/fdvlr66Q69XSeEcelW5UY7jYOHdUQQ/W2gz6+qqhHl2xwctx57IuQbQu1JJ
aWNL6VGSiA6NKK4TX9jaCurJXlTxZfbIJImmiytH4vxDldBXD9h2/U4I5f8vKOft
OBWVGycg3l3Gfk9YRm6RHNpQNH1tvy+kPY7Q7eS0JVGqWyjeCTC/SBpfkklQ8RW6
iSLn8GwcwsJoPw9sYbLtCWQ8pT9B+uKYyaFtzp6J054yHm6UbWYpbH89nkqe+kg0
4oIBQpI4Xcie7r5OWxxEWbf+E/HB5Jsl++tyAsDJdpDteyxVN6DPgHDwHuxLZYA4
B55zxeGOI5XgGLl2BIhElhsV0SbXw/tio/YKK1ndHMf0fVB8sLi8PsKWuikVoSio
i/9MeaKlxYHC12x/C9huLyWPcjwujpflEl6+GfsZGQnDO7FvQnF6fOU4BsFgOgi0
vlHfpx9RevMXZVLooWyTqsLpSmc+a/GsPeExcqmqP78B6x3eQNLjqnO65HOlC3ly
GLtOuVfPf70vtg8y+/gdf5UgxUwaXT2UgKDdo+aWvIkpwfJOiJnqTmJv+8qLLfQM
xUFSBLTXv1BCEl4QCi3+oTTAr27AiAl5fapnzA0rgd+Q7WAg97zciTZowBypTB5l
2yxy0fmPBPknNahEd5f0uoAnopqExJjjWMiKGpvaQfhYcCJyv2w87xpopdcpu0A9
wVxgS2AvdAHeKQ5l1M+BcrRHzOkvYv3zWEFQVVlPCrs6sJXqhwfRBcKUut9TDbL0
Zh+39oB5sQ35vJ/I6AZxUxdjU46t1NaxBx9z8Bc8RrH8qoQgS8QcVqTzDzPkbSfB
XY7nZgywhStWs0lTRmFHk5K7avdLX5PJlkbW9f0cYvIXMQGrdaOYrlWp18krVRlE
uIbIQQlms1vu047gPP+mYDKQoGB3ZtpKPo5AEdz2CXZcwPOzvSVkIRFsbC9vCG2d
9QWlF2ucXvzlHiv4m7xamHBb+WrQmgB5Yg+8jCanujNDfqax8TxQF3g/KHVABR5s
Nvd/I4pRJ3Yqg8OtX6+R52Yr/aA3+ZxmY6ZvOIL+c5wEHGzG8kukGKVRQ3C1zV4Y
8UhGe1C4TogB+s5pXlalpRluCTSAslTJ95YWigSBawP8KXzlooHJL16xaaq/r3Nj
d7IN+jqFz/nkTboNCnIRylQ0FoTU7k1/CNuG1dKtiX69CnRazgS652weGn0GuiNn
7fHFN5i8JBid1hVHdLJI3dknFd3pD+oYSd+OfpFH2DrG343mDgkPCESTVF1IICMM
ZgvfxRmdxOiPC46DMci6swxVu1esoENwCwnRd50V83Yzfch+TBur0oacocxvTkz8
+MKHBvkD7NAVbJJ/CYp2NsEcwRujEz/Q8WZ9WrKWKdXh2/7rA39DSXDYSKuOeiBG
gZaMvrQ/nM3QEbICXk3qx45tRn+1fptGdEvt3bT2hZ2pVds9lrAoUGjRtUjeldNz
DX80z9vYD6rEdaF+L7zefZRumyfsM4MUFmCa3BL6Ww8vEQ7SW6I53yABCQCOpUNh
CEWJ+keYqEeoo2c/3/hjaADm2eUi3ayFcNTigSEJdIFqmd162fjIBsS2FILXsdf3
uQLruQORl6PV3poE7Wgq1LsDiMmSl1r+vCKDVuxPemcylW92VQIGaKHUsvr0R4Lq
Pz4QGMrAiG46+5XtSmEUdVXI3e58EWxojV9GCEAlt9DbXa3RYfHrRlA2+QVTRCfR
sFkDZZQf+IYs3u33gNnKyi5xlu/UvUGTPb9UCWVFiu3d5F8JvLTWK6eE8L13ZC8v
Ww8umJdIxyG3c5YXoMfKP0yL1tidNuatce7powOhO56uRjQrzFTSx5OPzk+jS0gM
7ZE4wihQxzUBwKdh09FYNgLSfYJoZyRmOk30KqxRL3+ih1zl7iwOq4eNRAP0Fday
/hfo660M64sRMg7claCvqtPAPTp9U1qU3CdTqcJFQC9e5mAYzSjX9FyC79OId8oh
NGtyV8xUxPLAPdjBxvhjJvdyRLVmWZ39YvGyZy05YWZVRdrq7orlU3UDwYyy1Tcg
lhFU8EsJEmo37uyLwE7wXKV7HgUM+sHmXe+t0TrVjl4fnBkPOdIy3ASddgtBcGtG
/IoYNtoEX7G+r0JT0g969Pwbw/u6NtVDRX/ZSHF258xqCrK7YRof2kJXEIBWaOsT
7wD3W3tTU/6xBBVpYsj+H2pz5Y3Nhi5EHzIKSgSiOvrHvzSCUdMnOIMqlWz/dMHA
ml1Nu5XzwUuV0MFW5oX3/nPBtOOchS3kkcNQwbOaRLMgzK8LdFzGiIkNLYWnpVir
tMKheSmKIOhGaMHyALbgoMyAMwydJ8y19kOiUmeFI4frgBLzckVuWti+a0xNuJGK
QQMIEE9SIjHrvGz9w9vZRQ==
`pragma protect end_protected
