// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
TdoukM02lY0vNZgRrxgnQ9xmYgz4pIvHyPeqqlR1DG/g1BJqg8LjpjKvrOP5+r3XtfeO8+k6ybux
Fez8Jxyn8Vk01SW/1jgyO3l6WnttsNAZRe8jTzZ8QzeLDx7cUPFajTv0XElsUEmzk2sCY5QzbxmJ
aADPaFVlhF0fT3/kUktlnx1BOxAGGLftKvuNenqCfQSPq3Ykgf6Girmuyh6Hae2rXG3t5ajzGt+z
boBeMwYaKzK1NTr7MsvznokqNaH2DYdQkeoqTjqnuWU5V0XshBZ5pd8X5cjamrCKyPIEhq2WGltw
zviHvYG3/JKmJCBZDduodwxHbIOT4pp7+OX1RQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
4uCdpenIeQQ14uk0/EtY2W4ngtk1WpJzUv3e7HM9RSMxUeLeZ4jCy+lBpsB6IcIp/fPzwZqIfdvi
ZvbEEasGeFWTZPxt9IyqiSwJkCmkmZhxlNJNAmnTVlyFDKZX9sNuuaXdHRSf+vMIKj5c25QqIc2W
H8Q1WP5LyS+SFvEJSJ6dfPbIEGVz0C8C7py/eQMjcAcXgv1Z/lQPY2cXda8PSp0r66dpFIfeMuAA
OKHDSOpaiiVQV3PdMJu1xVTMmxS706qZkhlevydiY2GzW9oWI5OJ8I3dbntAvMq3DbkAINhRBj4m
7CUf9OY8WjKMTLbj+FYeQC7qBOp7cEChPHswFnLrqPjcYxcBekYQ904FHAqe5jToanSOFO69/Ntw
d2fx8KpED8goCjAchvJmUK+XSnX8sn9Bq552b6hZAPkVWSh32MH3pcC3pOsjoZ+PqqSVf0YIlG+Y
YsyDPfSpXy0ZzLPwR4QrIMUYyIdDE7EJD31zGC7PX4YMcSKZYG7CaY0jkTm5MI3iUHjAqOIuAmQ7
MiYdcu9LJMwJx31u87fSv4yq7kmQTuRySvloSUCk38NVrmEjZM4xU3qOeVtqwY/c8mwznYLIc3oQ
HdQkPUU7+yO5EjzG5ry2Ky5jAtCmuV0O/3RfuULpVxKJ6chqhM1pmU9CtUgtLJF25wbW4rick/sT
FmlfjQQKRl6wD/xmQDBGHJ295qZxzc/aHnT/NHPyXRLYexA2kqmKNsC4ozq1ZHyhFo10A0KCcEL7
CcIjol6Aob7N9oY6a9bQFnlvOFv+9Mm3Nvkwt9fFK12oxY+g0dyBZesGljuWVogbmaKAO9lb48b1
KOeQu/ynhKvB1WkWmXv893x3/Q/HqzvRS4SuE+ynJUovjJazcX9UIV7XY89GKeVMBBfjE2TRahl1
CahF2iU1p2bEF2VRFZ7AOgO5rrsqpQHEQsZXQi2tzZm0iTYB/O/kfbmU+EvZDyaq5+e86V6Ti3Sx
5keRdW/C2hyf2FLaqbiQbn5S/rpmYID+Y/0AI23MdWYNRxT2nRz/buJwq6jLTpCVUbZmv8Z/wog5
eix9Zfr3NIatOFc0omFhJNZc8QhZgFvTFsiVPHS6lk9pzW5VDUkd8YQ0J1QpcXdXRSIWsP+UdIQu
3JoweLGUBBzYwiUU3n9c80a/kF9NAriBHx9n2xEDRnZTPViojeam6LH364LfwmBqqxOXeETC8lse
HAFL6njm1Ma4NIGNXb1+wWh4F+0fi7M9Im2K0N8SQGwqUXMOhIHobYZptN+a5ZsS8z1I6MjtPcYh
2Q7InObL3y33j0EiSzcMy7dYazEUWCMzuLNYikyrlTWJeo+yJuI+fY1dss23cM9ZUVOWoGmuMWmf
jD3AVf95lJYaRCEm/grbYlOYKkLeiYgmPJT4HrJjt3r21HTVVRrGqNNT6WwEQYt2n9Eiq6KW0/0V
4J2wVDld2CSbwVyPvh/PXGwmCvBshLV9uFwhPmQeo+jtTdc0xYYjBEgK/mZdodeM587hk/iZpFuq
pnkl5Y8iZnPpb5nfknl/xN2T/SJL5apP1Csy4ACFTfSjbMDUk558b8sSzcwPw3AhblcJJ1jbozbN
HREn3+YUhyptvq8gNXdzQEjYrk79vkAeWzBPl5Ph1Fmx1JAB2s0fRWV4Dpbyhuvd3Xn8d04sXV90
AhQ1v8docs/Kf0y6D7/6G3Tv/PW8vkwEbBlCjO8K98PtYe+s7VJlVohhBHysDUktXs2RG9rDtl69
op2ruwRWemJrZczUvNvAoUdupEdE+Rnm97dXrm9sDIFp6UWP3woS0Qu9wmjqwBpywdmyaaJaUhxK
j6TwK/JV8C0jctM64i100BDKU0qkEW2xYTd7hh9CYXRWDTvqFnmmR7jqSfcXiSYiLI7RgBxYj81G
gAQLzzMaJKSoPeYO+wnNKO4p7y8JUrocirvjgzOTjcPhFDAgc/HkjG7DPzA1KtPsTTQKWd4li1+f
3mIkPudTjfbHC15GtKcCjUiawS8xctcrIl0z8OAM2z6a6EwjlKokG99pRwi9N+wURvxoqrRTd/kE
bIGScEfDPhUg9iDo89rqLYH9lSHv7Y7rdDVyVtgRLJ59PyGke9lAf+naAZwLFNkJ6bQ8VU82x0AI
7CyIp/i+NVQuSJkwnzsGJcGyGU7SXuWC9fUJwJg1MNkCD1iG36oCI74RzfOc57+EKynTNdHM3KCZ
iAIFfGLJYzpPuIbmI4Ky7mbIGypi8yr+lAqwi9eeo7QijY8eUvzMSPwqHiMbx7uhSoI1oo2mItJk
LcDGf9eh04NjYzVVf3q5+/AV6hXlfO1neGUv0dHv/xglcYjKB+GJbEVjKY+0l3isQ0igRVay9aC2
Tv0bL4dipjALpeXNsk7xsWRnE6rXgcjQT+a7a91RHLO9Al8HlR5Ov63OAVDdclbtmob5PXSDELjI
zJlDDgXwOcY9JLCGlaVe5QWF92j0CLifOQaK9xzFFpf/zNshOknk7oZoskcFFjlM2NvV6GTqiaU1
VQEu4q4bzH5UmKcQuROXthcWIWZeO+qeDFXMbZfs9nwLowOHQOC+wzTW1SsXgVUpJijcqyK0N49n
4u0JP30aE8oKomGmyxZhnUt3eSCV6FU5fMeUYSjMXnXmyRiYx3zuE1wUsX3pjudXhU+pyeJfEQQV
bplBpINfbbzGARftpx6xWpjbly+xpxFV3dhTAzQATKAcElQc4HISviIG9K9WG4Vh9RQjC+X7i28F
+jEDnFEeCOL4ytexqw+Tq82CtmPYydqCWBG7fo8nQ0ii0Ic9z5iN8R8KZtzvNBHmD4zcKGmIcjmx
POGRtdXeutdxRMfEyRWEOdtWLkvzyCstcD0y1Iz5qNWjs4oeEi8MCZ42BxScMpg+hVOJ4ZkA3cv0
BsbDYgo5IpM4Jn5u9wXioiHMcBfwbkYNC32mSKp1h/Q0jlNl41rIafUXxO0e7n5uNGcHAIXvTb1j
HrFUqGaRpa41sR/EdyxfZsCLsa7j+g1NV1HleifafX8aEDLNyx1eCH/puG3Tmzu8HYA8zMM8lsia
+R4vR4VFtXrmsX98GGMoQNKBOpcyNFNbU3pVAmLxg2HgTb+YT66cpaJaoWFZOVsWS65EKSdhtyWO
6uRYnBGZvFSQTUy0N5MZh+aiv6zJZ+lA38IOG9JaYjrl/2QBdumBoWWEeos7mWWl1Y8da6+5mo+4
FxxYyo68u3SNE3C0qeRt9isxtVGS2AhzAi0+urk4BGtcct/RCQSo/MR31Y9nX/wq9LqW26tapZZN
LXtJxf7Xrqlh//u4/ynnSVg8FCS8L93waXlKqtaHUlFWlrk9WuYH6JDrk06n2Zn5XAu3JihtYcm4
QMgghxLr691s15GpcwioLkAdkYJ68kdMvWYOoByTLeDzKBgErN/1SzH5+Xv6JQKW+huGKlQ2QJTV
nHbjOgzbmVWdelMzf1/P0cSzeRZOymR9ltkPMpQBMQSAR4Joq2QW97eEbdcuTY81EeURop+enOmI
ebuAKaHGhwvfd23Zp+42Mk1cpy/9ZMEI34xmYJcpOOTPGpuwlhldMzJTyTPDs2R0zv4INExuSfJY
EzPGCAKYy2tIFLJvxHGRqDaI6sJyQaeZH7zg+s+FCoxn91tYtg7fnCBReiVYuK+K6Ot1ji2LaH1V
goVXoWe8VtzFkbdDgHwnJ2GWKqml1QcUMJSy4+4a6utuXhQSMuyFHpokCCVhNmjnz8o4hQ/afNL0
RTF3HgM/XrVgIlqOjTqji1apOgqpAo3MRwBl835rK5jm31dtzJJsX+y4p5Qow8aHxnHVuPmexcfh
REf4Q/5XbzaSNUuir6Wlps9Lfxje7emXGNfHJCjfu/BRWVH5f399WBJLXQwxwzzyumBW742cheaZ
+Rx32uZVkTLWsMpK6TRX37d1I68bJBnyhlM0afB7ihhkbQRM14ABDH7gjE8EARvURhIwCVc1dN/n
C4fcaqNdsV3ueNsGM983zLW48/LkzOYDdlFYMrLtIztIel8I1Z2YOVkFAKJ1rKw60mwVvTzxTVia
hRhp/pxJaUb+IOiYeV34uzTMA2Sg+JA8Zseh3oHD89PIazCs5TKac1SSIwvzln4WgzauUiv+XeYV
XvjlQuPPie58DsPD5pCKFo1mSPbXy7sEz45XeeuyIYYwoWtfn7Vmrw7DUHLlBtU4KbPnIJnN6Pqa
EKOsgGI0YqsbiIXdEgfTOlhGVr+mj4hTAPN3Xt/FUnioOMjQj5/j4uMwG5sU3rpVQlYfAir5Oxgj
dygpIhtMuWyxpZ9PUMor/0bVDq1zaw1I6M5G006dB0ovsJMqi4IL/wHn7vf+ZbPoLe3C9wvYrjIY
NPpEHGNWQkZul3DF1c1KzZtt7wr84rNOfk2vRYSDSaNmkVldkwHA70EXLDP0QV5IL6dU4iqq7cR6
apCw1V2teqPRK+eGMkYBI5xktoDFUJPwFC8k3+ddETAyfQupZthUOKxQtPHR3jZ9Sc8ua8H+upHw
S+yJ+JxSBlr8QFSiIUlv+vYwa+3R3tQZmBZ0GLKcBDOhY/AO4Uc9GqNVycLIceJ1PRMTN1XmYvDL
sybsc8VFJrLFIZaubIK0E7DRJY67YAF8/xm9KOOI2XHqLPh5y9ci5hSOn46EP+1JSk1XDFf+NfLD
5pZAENUz8FXDcxkHcmOV5Pqw2o+Yl1w7jGTbZm6oNZxXvhO4uRB8IZBWxF7C/eDH23EYrzzObe86
oXvB+Ap/pkBTn5mQVD5a+UdOh3jmwEYXiDhsG2MFgpXB6wIIa7QdUKgAyzOhqtqpIFAZL9hLhKEO
WP0v1DHljqPMCiK5yMJjpZyJQgGzYsLpGH4sudR/0oc7ebHZ5qLWwWVhkkLfHNUPadjpJnpvCkD7
YYqaNUUnjkcPprN/rhUecwXO5i404YylQYNT4Ke6tnOINhVooq98vB/Fx7DjWpWb0aCmIurUKmA+
7sOnqC4w0B5DvcvdpRC161D4QqHocNOD7SJnHHgUaT8voUCOl2lG7eonktxXtJBzEjmGcHpq+ZBu
YfsW6DlrUpDyfe0vym53VzhzCz6gbO3xppgsiTPA9uHoBpoNOlnItmDox6ywHG/01DdazG3PJ86L
awVLIRa/alJzGhKDJzLDHGutSnOTQEBh9ab0Vywyx5jkNFFwmrBFvrEyxrOo7OxaqUuXh+B2fanq
3jvDLgo+rSv0eD3FUQm5e0XhSbPwXIT9dNKgJpUgifFd70svDG/HulExNAO3BhjAUtctSIIv/OA1
ksrs+aqEbD28mv0Xn1ikwYJz0XKKCisReIGrkqKFdNh8+wWVc3btdFGjqhVC2FGD2bIUCNctU/VW
1aES3LvTGtPOS9GclUU3/FFZI34u0THSldW5rfWwN58wnbLY/0D0pVYEOL8QcvFy3KddS3XpCaJz
Ki5Yn0tqMMOK9FZgwJATI4sHjLRHLRTqCUKMie5+IRWB5q0k5CvQxHu4xGBwWp4eFxsoSGSlMsKG
4Vz7q4XPmjhaxglwktkM9Hptd0AOdGPP6fZsAeiGZCZ8Uu7eXo1cVbCOQ5kJlHbLiSaZmMVkTWvt
/+0AETtrfIiXc8xquSCkksWP42L996+iEP4gs27kT9gFgApWP69pxWG1h0NGY20mb7M2DwinMtC9
GTlwySQfMVPWXTC3bwOyMqzF5g5jWPFVrzY4rRC/7teWKHKXGLKgbbEsAmLnMEzfAC5mw0kiyyxd
6rCzdDfiZBfPKGRLA67Fmhif/zvIFvWR9vIse4vVQIz4CNJgSZjI39hjLCVM/5OOWNGCqH//avA5
oUH8Pr86WGsyoLpPXPypEEwj/4p3k1pu78Sd3zPyR/l3BQLs+VB1486SH5kei35l5lCf8Ssxsqj9
dJU5sSapIj2QuWAEWS2uym47F4mcKfFSc+LgoUfbDVzGl35inegzoOpjOobd2JCiwDqDFqdr7VIQ
6IIaUA0N5q5WLJRNzj+Gsoq+DXPdrrD9y5VcZbVouaioFTmt9SFyjVrU5xqsmatG6LqeQWmGpK0L
GzL0hooCSBlTh7vp4XUHe/jnLfHJa7tOwIjgj9vaKaZ34EBk4uadM8PiYPKJYZJ5MPNYDz3xqLaF
U957t31UsVw/EiA2yuYDOSZ4dxO/+P/XZcehiZQlmYBJZRxbbEHoPe1zfNgjoYoLw40O2xT9Vm9K
/WXLofUpJOewJcBkb4XanORFxmNFXPujFrM1mY621QJUej/NDAL0IV4xUhw9hc2NeA6Yt/j1byV0
3DIQYsNMesWc42bd1+mUOnRNSHfKXbonPu3d59D/P9B+yEjxwvjxWHtzz9uj5pdBSQHZAAd/xCfr
sNYWD9wTa/G7ZY0hpfQretBcrgSopK0QEzf7BBQlUQrKdhcjbuX1viz5F7/XwERhJF7qJwncIK4l
V7OjNvf8UWVj21O0WSS6z1GnmWRZ0xG6u5trX98Iqe762MH9GnaiMGt4DWdaa17Nw/fc5p4BwhCN
yGhIS8gIgH3XXLLVuqRAZ493R+sMb7DUlWKTi96pkIDHIQfGUJQzgPlu3xDYDKPVI+YDHT9vTiDN
a+JlXYg3XqeJq6IcPz/5DSlFnTcacF0JGI+9edFk5I9fL801zcEs8tJC5/PJ7g7mYFS8R+p7ANE8
9y4nr/Yr5IPHPJRGtczpat0KREnB9yCocMr54+eO8TNBtqsYQK2fLOmT6bQ448bpIB3D/g7RAbo6
oAOws0gUZTmgWr/zbegSzr8bDVHtiTqEd/SPiOODUiguMQPmqlFXWmtXWBNXzR/NWZZVfv9eU/gp
f6rPUdaHFq92+SXSBwc9lbIoTeHJmXHwljwvevsNiCmE/CxzbRffTgZYvLLPf0SicTokmHL44WVR
6AHBv7fbyftgezipxejayQFNJLboaGnm9eU/W1AruvJcgKXFcjkwIgX+k/eEcNjRsUnvwoHBwCiX
cCRaXXFZRj7Mq0/C4rqczH4EAKmLNOuyytzku0/StsiE8//YQ6TDlfwHVMms46ECEVi2fP1IP+Ji
gR5aNwqjeynRn5tW0oUvFhjdUm9wV3p7kNLauaSNO+w61Q0BuaC/P2lhoz+2m7hQSjh92AXhYZP+
4n4mrCvhFvJssh+1+nCcY1s9A9krHBL8sdW9D1t2y/McIwNOTSnaqmbwm/HVX4A+ge3/J0KIOtDJ
tbCWFXnVrZs5sLzl697PuSWgrFWWrHHwd3sETPQ6+DuEVyV+SY/dGYtWockrR8fYBvI08xA+CLN4
9p1Yl2ocy+JZ9XNcMGRSoWO/rIflB37fl6pZeb+deJJ+CmJ5dfDTuiRe6/czhgqP4T7Fy+UB470z
GMRTWuQbxWPptuWmgds/hX9RepNe7qW4IMNDD0eaXVdPhP6fkFOkuZFiml0LiJW+i88BfEfqC4ax
xsuKwJHf8YSLWHscKbK6naDMT2G34+yLnYfgdV45xPe7lv3p+dOMXk8QdC+j8rBmERk/JIF/pZfj
v8Z1QA0nVkkuIwkmjVPgyiOrZqbknqeKLNw/zH5QBV87gN15H+aMKck9SBEk4EvD/wLRo19Dudaa
04N8Cy/ss/VciITXeSRp2SISSNn3ANsjiVKVN1uN7VV2OqIrDOSZAJ/aIWmSvA2lIflOU0vhqiYs
z5/6d0xDwr9UzdvCZHEX//88A/9I7mMv2Z2jC240cpWt0w27ycWOEl7rqgvGPbMNgUBs91s61NuI
/IycRUeE8RZdDHXug40+3fTv0HjtsCnI1ja2s/kXaB1aC37jl/ol8CREhNtOmxyANHhqh/hm937o
eu15Pn3WBVynvEL8EcmudZH/p14rc57w3dOWdBle6/3ToHDb+ATSgRh7uDWp2YzyR9bSPfxHt5FY
3cuHo+lhWJpWrZ29Ew6H/O3Glmgyzp3YWUMJFET59diDk3g4KWzC1ziAGx5IrI8v+7pviePh6ny9
U4ngb/NA5h8A/XfhnzLDRNTrJ8fDWuaM+0ibOJg4oqBwKpQ1+TtvkM64NAhjiKaXkpS35cfA30WD
/CRyxC0ef+ADkedyO4YLI+MqWQFMHc5XL9Rn3r18ol2buKlTW29FvR1TPgiIIGKhSzNLa2W+b3Vx
FYl/BGEIjJPIdBzYqXRF5S7LxbATAe0LWkBwG7ewTxO/YO3ZFyH10sE92+SZzkjPqYxSscRjYQ8e
q21JA6uRdzU4Sx0FwbicKGoLPHP2z3J27IDQyK72DComE4PrQuk3aUcSXW0esQBJppatsWQeiBlc
t58tTPyfT2SWfQJ5TazXoo0uh38VeWuGS3hgg5+sIWkVZ2j6UmyYsJDLuNGm4SRsrKhNqKp0LPs0
ZN2ZSwR7+kB2j/SwoOmlAb9om6zED/HUgDFMKwlJvKBoKFS+xjfpEjIpCxecMf5dIu8/OQ10mNkN
hLo4g11YEn1FPXwGKis3KFfCEKDCMWaxZrUnOo3iHe4Q8V8o6e7MDuJw1rPnnHz8glkcbgi1RTfY
fnUaAh7XHEAP0Oa3C9zIKOOTm+ltNw/DTGt5X73dymllzeet33sLKAyzBp3k4OE7BREwfTvE7OdH
QEnB+QqhMGgUICne+AZXJZXRArqb+yPFWuE1Y3M173yiSGqVHqDcS1LSIQtbaTL7FQ16o3mJ5nyS
/C/eGnvoqVYNp9mj9Dx4LmvOaoQgX3kMWeyjxB7ict15tj/omfvxxG7mFpLljX5veVY87O31w38C
43mMceF3aFO5udRi3hK5DmpKOMCQ/FtXb7M4TNIQe2HCqnfcWRd/BUy5yg2ihkqiQcYLcwuS21J9
lrc3GenCBf848Dm/EU1MW2NtnC1S2sbzheUuYTrZI8S/bos0FOkevKI5QF8zjVVLOcKyvwT1rJu8
wq7wyQzpc2nhN/v01lwnu7e6vs2id+q33oZ3JGd4ndpXfp8cNnsmOCAIKxGZJQ2hTDIS3jDiK8Fh
iwf00qaNJeZEk3L+U8+Kq/0zvTAZSKorK24nmv02a2o5d+oECHOdFHVTe8cblPyKaiB3YTr1j46G
CjlSVvUgfXD/nt5GUQ76nINt7L4W1XeEM6xoI7y07M8TmAuSVaHB8iXcGyJUoBhjMBXYy2023yyJ
iaIsxiV2zMA405QOsUvJP5lVmWpZugzdcnI4mF+F3VMLiB3f4tqXmBdfO6oJx8kffJ1R6YOTR2ba
QJ505tpLxNqiJNhdygVS4mQ39thOJh+KgMHa25FhaaMqIRTQxC0QwlIgkD3p1JjhNMNsQ+8ChZvR
jEiK3gP7ZqTcoe6NNJso5YGclCI6pPgZgHjC9IM8H5Yu3PgxdAfBECQUMcJLdPNPG6/lfN9QSJuP
BTUo+bI9zUO8Nvdrq2lOxptl2CoV1DCVLEplL34meqjaCccfwRHo8EVZewbhvGGUTVTqMu0jbfrG
ulmX0kcQ8g5DroYi/fiRCMsi1aCoEGM8Cox4IUmxkzheogjKRUkD0e+u9DL3ILuQawHpV2YBNL1g
8v9jmGCmvcoH+B/3m9QMujcnLGq/xui2bJezrwMxzhQouczWV7GRCsLBN7PQAuvJ78BjVKYDP7DG
WHtW0UqC9oh+BbhR82xhQ02M/eyWFLh4T9lvsiJLY3y4pXVOMaisR5ldXFWgSp/mjtELn1wYcdtr
s864oS1BlgUqGbYXakfaYgf4ubTmej1IzhYZqsfdB5yYUSgR+XnMi+uCjzKKpxYdATomwLXlRVtV
R3F0kzU+N5Z9FJKhNrwnrZJOFX2LsDbpP9G+pjf9Sm3UFB04DWzLWdmx11Z4H63BsZKKpHU9J1J8
pKcK6WXNDRRxUjUpdgLxGHlwSi9DmSeP+mNdicvJLKNgSYHZKJpo4qDftXrfU2DjcoyDeNrsrHWU
VyJCquPoZNBg5hb7WC8XfsX7O2q+1WVq7Y/psgqtINr+JM8zgtyGvxIgwzDXuvoHev+tHhdE8hjh
Kn/jfJyD/0sWqVCeG69kirHeoWuhVKeyCOcfaWNpC8lWpltHp6yCnetCmRvzfoGy6kJ9pR0NgYHo
MwsS68Yifg1djMehJw8PxktWVoy2k80Eg+Swu8m0x+uyo8FlH6eThjamwWLJroPoAOyfG6D7KYWW
bXgIUQQqgIGtWHO9/mSuNj5zE4o2hp9u9q02Yt4z7VnuG3w5HqPNXXSraLu6gjUn4LPq4qpIbNq7
pgHbuJ3sgkku/JmZtgWBDmbpvW12t8uzTVX7SIhrMP1mv7rBvOx2liGgcMpjxSCsIo95NhuoC9LS
wdAN0lDj3EgWJYZdRUAscZwCLLAy6zFxCxXLzNNMg6CG9q69pZNRDb38dScONmIF5PM8e2ZfxUg6
niKFIunIXV+Kob2hUCdDYKbYzmFY54aE8HtaJcPg5j0cgy9L5whtRR4yByth1HRFXHjirx/cQiR+
J7ELQaP9PHvFhZP8rrckm2CBY17vRxWYRtaafncEUsqup2+sTR01Ho3pe0pDCD1U7wpQdZ+FRdr0
wqf6EAB9oc0iOMlH2MY1xmJ+KKxIASBr0x8wx3jbczSSQPMkeg+bEGv3VAfUklE0BV3SlszIttLA
LgdR7uBJFeeNdu8iOirGQJqiI9e1PJpA4gZPImY9q1qjHJTrEs2GH4IPMJJBhclJXzr6dSTq1z2g
NJWGwE+4syDCOvIy2zwtBNmNx8HybhRxzVkPefO3EMKSpBBGGGIppVdKmUEt6pxlotORWEhdtaKf
7Mawq8IvYkKXOX6RN2VN0NMmGEgh8Owzag4LPCQIWtKId+BEE7smnM0lLVqeuLPb3xlMDAjqlEjt
r668bJNJMNuFYdpMuYnXqWuD7tRo9kcwYvDkr+hewYkRbBaW7vhze1B5nm+5VnfakbAThJZdT2Ig
NzQDCU4eHMzOBYmAgoqn4NCDnWDOTNSMhCYAyRpteVq9dL3gIP9MCqU/+BTVk0sHxe3ReWxp9vby
AxFDpUn3A/rSOzKhRywF2KunFc025bpusE1SJ33CbbypOaPJbaqNOqOH7exQvcV8XoSqLrVPJywt
D7i2RxnV87aoH1rslgNq473U2jMA3M/r5tlWRUfevyqDmjWp9gJeAMKYCuhxgTO+lrSo7fM+rYdH
37Gv4D7SNObTXUH1IF0o4WI/6LSHeivwXZybYkhgGa5/fzJ5uJVUo+wAP69F38PuaZEn0I6NhdJN
vXKYvsNJCwVYZZrLtRX2NQVUkaT9C30AfWriAFDAnsxGxNnEXArRr1NinWH/1MSLNyTE94GeM3WX
0WOM+RhR7qrRurbRXqBs0Q6M4NkWIOIC42CN31MC5jo5gigeOvv5FcSpSiTpFZ9JLXbVV1vkNkdM
bJ/WG7pkPv0jMrmA6SgQ/9llsrSGfATwnR7tTUFd8dFmPoIQ3QHre2UjACMSVBtsOyVfxJd7ikMq
JvNNSbr4nVyOzco7htbSCdtzd1Jj6AISyU0t/2sEwEOZC1orvcpiB7sfnyOqrzbDv9a1U3m2uSoB
3FJulIRbzMvtHAof74nObZhwKbt4XIACNLvPR7izZwp8sqc2G9+g5QsKs3P951xLh1Z3hCQxF7ll
P/j+w2dd7Sm2VG/DjpAwTHVLpe6LxCczP5VT5iFrixle2d4JTHWlq1MnxZ0RVpDMVaw0iK8xljpY
EMDRATt6UJC6u5+bYswAMXch2muJ9qltLVHltja9iCYqIXENGBrwJA2z6D96dNi8nBGQghUZWgAt
SWEepPzeJhCcH/jzxqNW0N9yD2oIoqfA2ZVmVg7OXxW0bubfWdA30hjR2V6uOGwe+E0gbfJqRw2y
4nsBAmqXYvQQYpJ0nTOY8v0szyrO18pP0Fp3zyfcH/SRzhEQJOWzZQ/TV/34a+a85TFpG5CYo+TQ
GbFCiK5gMuVkO+agfTXtV4+/Izi8pB5a3STZ+bu3ExV4hsOH84xltIxjX5jnCTSS6xvNlZwy+3yZ
IYT8tZbZ77osRJ6Uj/h/pgNT3RB/D3vdDZ592g+zYChbeCLDJqVjT44Oj4GFF6iTUuKcYbYAc0Kp
ZznW03SbVXSkmZCvgQsu714l412ZBMtWwT7RjSzs380T2kzluWz+tMdtdgGu8xQskbSWSucpcHmY
TsBV6KPHhqBg0S7Zs+gcZGXYsJF9CRLEstHgib3hxfdj9gu0eJLjslbqKKuHq1h+J1+jTa3zBBa9
yHUP9lUKapsIS9PZzB3RtWA78m6NpEMWkW+GJ3kpYhhTJnf3mbFcvQ3lGeJPV9yl2fMh/kCgr1ff
U/DOiP9dO+Zeyk2DUMu23uX2rPnbppmsiENWhT6/MSz4hePfbaTabxFfRujDt/9ndaAz602n4gPn
ozaO35gAXp2jTildHj5hqnBEn18WxTb74l2c8Em7ty+allEv11eeH+sX2hsIuH+G9OUxHrvEId3J
M8GySZPwe8qnH22Lfh62renVGXuG9xTTb4V2K3qPVeiOo7ga4MS7jgYYC9rXlSwtthuhuUKSUQ6C
vzTZ0qWjL/nqi6VV01ocqN9oE9NhlKkCf7S+9niaBmL2dnsYrM/cIhlRgXwwaAUd2ecSCzMczUKw
u8IWf9vFN/Y1/CxpLtTITi8R1x5IvWuzITW4S3VE2+FOfXMtKSJswVWXCZRhuCFhQAztyN2dMU1V
2v7ejnK0b3Mt1IGZkPptdE0idhi2nhEEhHyPQB9H1wBzIRXisX0xabyzbuvMXDSLwb4HFa0eEpuK
CutR08PWku8y8heTfR8gFm1LPwjPsnp7yC7kvVG6oXcrfdQMPVSl76RgOHSiCQaDOk+d5kaRJj5G
3u968w3li5Bpby2kleeF6GaM3F9Qi4h8z0b13VKANT98CoF4o8TNfkKaL8UaKuVd+xYD+2Lz4SKg
iDntRTNZ/jekdmDkanlD86X1XfjVALMVDzMg3dg+yuYZMC8lhznaf83AXY0+EJUcJctEaaUw/eAc
ZIW60WF3k6HFbivQkPFNRlsdXBQvgzwVe7iZ3JU7jlis9QTrM0Dt7b8H347fzqWSyvJ3+UoID2EK
BiKYz7ux2IxZ5tGS9nL51GhAGm3mRmSH2tLqWWPLS2FPX3I1brVNzbDS30IzKM0pZYzKN6KQ/JZx
DhK51UrPAvddkKyKhtEpf0hfXyfMeL9kdQzkAGg090DuyWvumXJ5PxGmOHVdqLBE5mJLLG2/gWoC
GIeIawGgKwwae3Vba7w9X9RZz3gbmdodsRcYkLYfln0Wf/RD9YfiW/INNsTDeoifVaTlk/hgtWst
bq/4rdKEXA34SbUkcs5fyo48QP6juzFupnin4vFzIOXoSnvDZ9Rx7GM1IoM6jbWwUzsJtm3xwfrd
yVI5ZCXRcOmnJ3+slAYtFJvPCl0s2ztwAAvfGGbiqdwhye0xdFZuJyQVeuWRCUTkyhZY1Kfopk+B
UI8MX6ZnH8xH2ZGLRka1USO9Uj58viDgS/yYaRl1hLHvdzeONTAvja5NX7A3haPp/pl2+2EuZsa/
NqhT3uay6pYAmvq2HNFn5FHvoqRqSN3Zm8VftWkqtmFzXHD8ogr7Pd9Pc3JPBZA08XCCVJUK0lPS
jo9VSKzCvU+foY/RgfdDqZ9Te6MLWyh4d5lqrq7RSanC2I8s8W4S4HvB8mewMEBLpPT+7+BsohKi
qbMwFWP4EvAwA8wPkT8DCtcCVAEmCd/NeMybh9FDkTGKiMcuZs3G8ZBlISHLzJbyUIKM+rDac0zI
kycuWc7dvM//MX/8/68S/4I5/noxakuXAUjZgbkuK4RsrRVcgZb8S1GoG6f/lPSdt9U658Lzguvq
UrpeD6iyrpNXsNpygro4Db+xj3ueNAeo3SnYFO+m8vPFquE71NW9nHVfVj+sqvKFKgQnOsT2oaMA
yY3kNAg2gw9BjtqBVXK12bU/oKwL3z35ct/jYoASu7E3Bg5XBrvOTVsDhIhDzeHDxfd5ZvDOLiGe
4jvx83fekKWYqkA8DqAg50MVpzzcYbOfxnOnWrdO2VnC7eWi0OcMIkCjUCVAE0dl7IZVZ8KsSIMt
+bZEZMaoVV9CWpcIZdiL+HT+bf2MXnqf0o6wyu0XHS0GNgn+yV1gxvUWDwmuHfUq8B6+dclKWew+
bBJHOaxW4BKxfG2BkTVEaQQRnlWkvS/ODEf0qmzghbwrrLsn0w6pUeej9nlsUfOiw4FqeMmIYU2q
QuQNSeqbFx7Xuqop7x23qvOZcpyF/m104hHZF37TRKaDvl3SnbLk0iR1AUo3TIn01Iyv/hmfcg8G
TdOAzZoVDWSXPdP/jhIN0j5Dxz2pEQ0pY6YZcspMt+Kuh0/4rcZ5a0hmAulBrFIcPwZaD/X4NOMi
0LffCYAQ9PDjv6KtpgqJQY7IMYgjzEndIn56/sC2szdCoUl5cgDX+/jJExwESyu6fXawEy26CVvw
D/oTB/YcAeUXutjjOqbtLx7/XXITyR1b+gWsIqIPQu/p+pzWknr1UMYIqMZo1P+5TPoMJ82c6FVm
K/MAD+zoDDBBc2CvENh+AN9ChYelP+mxuwYymMJEi/+zjE3quk1nCYnawYX6QTtuSn1JpUpodkoW
vWpSUOL5drxZ7kF2lwW5nmxQw0O87MM0YAlAP2Q6isWFI++q0gsfKrwSdrjmXY8XWrjqJGKdIM9j
X+EIbC4kCFSYH61VJiDEIXPfUc4+o5sF+kjgC27mFHiUGBZ9DX9T0bzudOaVJIX6UZFOAJ69b0tB
vg8HT3k5DdEPPMlUKWurJZZ+eLqp1Yed/Q3LRq9+FQwPlQR3cdY2zRwHserc4gj/
`pragma protect end_protected
