// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:35 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JYqiviHHiQ2Hc7DuWlOLAf8/m+lcuLJE4HEVY3smtaToIc+joM1jFt9ifCsLE8Um
lPi7hWh2h87yZGvbJNXiGGl1xM/vN6jZuj366351XrSn5I5LtFDCkkvWcLgoVCNm
nrHXuqEhjzP+niL++XsScqib7Xlu6Q4oqRqCvM9Ke8A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12432)
XBHef33N82DhT70g6cq4g7cUtxmhKSuG5JLYJvlg3mazTbWhNlsUYu7XxeQxoP2S
mRdD1KK3Fl9O88+tZ5M7RGap+QQnvA1z59Jpdq0QwudYLuitK4+HIY1X/z17p7Bu
kxxG2+4TXO25H6VP8dU+tOYqTCT/aTbFvmRHhrs20wdmtnySdPeebyluHWb/XNx6
pQcdnhadX4MXcL8mKwLYYX0gLHLKV37XTYrZ0kg3nhjVAw4ApgG/zktPnftTYp8s
KSDkhPGiNkaZDcS9Y+7LNubB+diC1sdLEbdsYWsp77ZFkzJ8JfAFatsYmSS9TETl
sfIejmZsacEflkxltQ5hhubSZPIuFXi0L7lxwHmlDzG4c4btmoD7wFk73y8nUBeh
vi8xgxqJ3S6rGHgrHy0TDb/wBY+nbEErgcbJww0kEFyLdXmZazPPkIy6Pk/1WmoI
X7Q6r5sjlyEbg4IGGnLTTa7g3qTfJMRv2XWW3NxHCJ7qxl7kmYjPzno5NeGp7Vwu
bRztgKKR7eUxF8VTbb6rQMWeuisfPCdta0d7Cl4O+qIdjwJPEBVeHUfflvJ+WB9W
6Rl2N4u/J+1vcAqcHs9v/ygSbeHCdzNahzRAFSZ4MB7wy5Ev7hRFwBoYeTLHbxIO
eUJfg2s37BsHo3BLjqtr06F4Uk01Zh/hKZ2gogXNSyj2Yb1llg3mZCSnGhlMSGZQ
n3MRMER8lTC97M9dcW/X0HsnnbpimCpo0C4XSCMwYxOhz8gSJuYd6STyRsNDGbb4
4icWIPyjlQ+skW40panCkPkkQHzfkJ76ZP3NVYNVYf6+oNBD733B5hmhxqcJJAmh
+aqhJMOY568yBqoLhgvWLX7sNtz8pLRxF4q2JqTEn19wsspZOpRv1Y3aLG9Z/67j
p3XJ7vAPKWt8DguxK+TmtOsTLfFyk/3847voaGE3g7dtX4+r3WM+PSzEClwHiroE
9jdbHpkSNpkSq8gYuUqMJmGGDjV6AXYizElBBIs8yKBFY8W7/zPpoWo/DXQ8n0TO
Nkdab9DpBCgcccB1fGnD0vyAe+73aqieG8RLz5b12XH5Z8yLWO6sIb5VdUumRqRu
nYKst4KtxVzN22ySeD6IYArnDK4mWCk+sx8H+h3eL9VX3BZdZGk365XvLEs0Y9Di
UMUeuEiTsaeSMmIraA+Hv/bcyfa8i4TbkK7vZqi+kfAO3LW0gFMVXjxR0rbDCkrh
Y0LcEP9TCRbEvE/OqlbUhCoppD5GuSL94lqWbayb5zMfRoo5HYT32ERZ8iSsSRrt
anEmCpcdn7WU/d6cqRcFhd/yNgP0VYPj8bW0DlEEfmSHYP50ampCt3jTv6XPuoEO
DupMRZOgKuN8ML5J7oN1WR2Z0MCi4Sap5GM1M2C0rZ6Z0B4nb3uQSb/lmxIverr8
m0ktBqq5jdYsMN6i3icQUg1dJK2hWm6IneM6o49NCJmDNTI7ImF+b6eTUXvnPQSo
xYJ0llIS/WrIyIZsBw1xd8BuOJU1WID9StvG2TeGFjpL3jPHDPQvvcUKWjJ7DRtA
IhsWHW42+xgZxIe5D7dnN7UPoha+R1kKIKaeDdOEGCs/D/32B4hn2KKVfHfYBhsq
yDEkQUT77fSprzCbEUNsFDhR3U1HhzkLZdJJ7zxdwhQ1MRhSNzF76QTrxyFj5cMw
PF6hrc5aYwV2cd4S4VrVSyMEzneDh2HzwMe7Pmv0ThZvq99qYazq1SMX/OXDAgCQ
mrUGbX+iFOge8bqD3pe0LI8dDT1y1UX2/De8LxQSmRpaQ9Tj0dP2SaEexSJ1buHj
fMTokgUjbra6i3povdza72nLSWrfXnLJfobzAxoTOEXv8KIEDWC63VSAa6AWWZvj
Wa8May+9m4edBMUZ/jUAVqEcrQsOFpqC1/+mTtXLNNtPL9MM/QMQ32ytKiofZooG
pws1t39oXjYB/m+fHNtJsHHavhHbRD9teSSmyy/f/tL9jJphJt6oCLaE5tPWArwb
eajjTFFHNDbhpQ+rlL4NVyyC8p+NVcNmOd1CLoMTEjMSXYk1n79/gH+c8ZywK+EF
EOOwc+wJ8NVXMVQBQzTQLTU73F7ZnStUEJ9D9uP1k+uP9wSeWKaiFlbdDpOW/4vi
VLHWUOi+nszUPha+7OyG3eazcpRoyeG8FYqIxfRSWmgeLjGM+793F3pqQXJ1we8n
UdtJlQeK4bniYOcQaHd24tjGlka57KxP/Idhf+d94MpmoDcg+kyzkTZC/VoZA0BQ
3f8Su+zNon0w0a7ZuBZj1bUl5C4ar6J/raUfPs+chVGDJ/TZLkdRkMIl9V6sWP4g
jBtCcu8o79i+2fuYp1Rt8RbVz9uipEjIkSt2zNCMwhFcpGtZpzFWvirFavse06MA
Q9ujzrY/Lhrj8ZmtjQWB/fsHy50GEMFSrZMY34ABw7C9n6sn69Yr823ivMOQOkwu
TQK7jsTHbYd3p/KgNHcHqwZ6yVb2zcGoQ0pmLUOUbXH7D9hQUL50T/FBeY/UYu2+
gmYQa5igw86akXwUkHcyhrFMvKLyHqTMnfg41Cln8zWNM8ZWdXSr88OJywbfBpw9
zE8yAtn/wAonrgr8Vsi21LyuEmalrtUxQTi5u+Q0MeGrzDmefnoCgjiF3Nqg16to
rmxpzrPXBIYNvtnXhtw3Vx0uoQZuAnL/uGuG4dPwhSFoJbotTGiUkpOmskVa6ep5
ypeFToRlSfhWp60lKbIr7EeVtyzm0iitKjraDHyzI6XX85PmScB2J0K7BxRR6R55
M/dXkR9FPuChBm1WGVk82JW2RMn4jUeP36uItASsendlRpoI2XszovG1qZ7KZsnB
Tv7qtQEfPKsTogrZ4dxgIvF3F5yL5+4qm39ch4dUbIxugy7GPllO8YWW8H3M1LMU
QNVZpkgpvaQSU0XVfXeCb0Hwce/hmjpU7gLFEgWzOyLP+8GMUfK0xU242WidfjkM
o0PQ2ECgIbzwVomWBFAezm6NrP9mW97EjV/jLeU+bdMNlvQjORJGGU5WdQA1TPuN
ptM1oAI+C/PwdopgcqqbJ39hxeZQUa3Cln/8y+oF3ESQ7g1jp2V1yvA3nBLFcJJI
i0a0BuZpZGnpqch+y1XWrUT3RrmyysIVNcHGzxLNjBdw9ETVDRMJfkMzQBy8BS4y
Lrlhd0LkJMeYXQ4QrNHfSB5cX5mq//6do9iomxxbYA1t330Zh2FPDeH3NqoGdx1o
zQ4ihk5lDRCEAX5fbBO3bbQ7sSW3Vg7/i5mng7Q+MUYqHPJTvclGqmRMrcKDDUeY
CvIdpiAhcNF+wqx2EMD6LGdBissKB1pLRTI+Ci8fvoll2751aFqoZBNmCJ22cLBI
C4PzbUTtK/eUtxurnH/HTXAd12p2rVaXT6sXNejSsclgK7ZbD2MWu3kOQBdDG+v2
AocwBBnRbtptDgs9rRQHEc5CNTbRI3ZwvT/aNNCvYmpI0+vfAJsGsC4IyKjIFurk
NuG+YUUQaxH3EIIjzDmxyG06cuV9r0ffLTEvZAB8cX+DZxMu/KUPEgN4uLOP6o0b
JGZF4I6OtpVBETJu5WBqpm1tV+1MSBu/PD+jam4YXrScfkIkpOP/sw/8DvNazUQ9
Age7kAgkOwhuPQzSg3Bly38OHEbsUFObgtsjNF78U4/GTohVo6tjsXIiorc+1t9D
8iL7xe7JHmWr5R7kcTPc9HvIXtwoYbrn7yYDohGuX40U20QRfFyawZ4wjH6h72NI
5zdAg/JNyAyShdAKz/18OXNrzs4VY3dd1e2z8gW/ou0PILXIc2/kYNlq54zYLHB+
PH7utGYuq7lIdjExVM0TrPdlRcl9XwJzGqTHXADLFOmE8L+v7cy9TC1VYhxRj3Bo
zE7n8PLL3rWzi7Im15OHMFWUv0lVRJPtqy1cLjTxMTRO7LTXCJEAmLUSmIe8LwqI
//jwQFnsrcRBrRD3DpqQrM3Tfv7xdIA4h5HPwDQ84Q1z8tgUZBSZ7pxn25xuMZx8
tVWjY04Hz/N4LWyAQY9nizv9YuSKkjU31jCdnsxLXEAbEkplfZO14AG56yyr/KDU
KHx4GWb69ItIAyRLI2nZKWBiGtVHpneg84s8TQ1NcNBsAwON+2OTy3oP3EoGU2hR
kKL8/g5f9WP/8hyVLkKRGFFB9dYLrmoECh+RdJT47O7ALrZiKHhsQuq89bSGwTRB
lYpneppmPgsqYVWGE4DRpsfWwJCCE5Ho513znEAgx2o6KLcsdiEqTVAnYo8hhiRR
woZ0c0HfoX1bA9XV7OJt6/j8dqW3GLfPPyBOcYRU73mUsuaUGPX+6WDXjOM8M2Gx
FMv5DzyP0psG/jsrcPZ/8u9yLINhp2N/6Eo0wg7H1DPWlwWqmelSTefskeN1QJFb
1Yuc3HpljzlVXqF+dJs/TDAFl+T5WYDYgFpGJ3xcLWEPpyIXjjY1/3eZBIpnL2pg
OtpuUBGGWz6jmR6Ygl61Nz6xXQMQWJrECtv62nIF4y4ydJ+WfqyHB+GBwcMGTmTN
YBMsecMCmZyYer0CPQkuSb7GlPdc1IqxBJ95UXctM/tbK/0cj9WlqF0BFJDsHquz
kvN1YhtEvAgppHBnR6NJeybge8RFjkJfvQCU3mzP+zy8AfRmFGh/krjSK/yZ2UNh
YIern3T+QmxjQG+UuJQxtJuvPfvr8NmMoeB4XwG9nF4xiCueknam37V/pO95+QIe
oGsCLsRG4BbdMCupHkT7uBs6hQHMnHvWlgLrgxKXjvJoergP/l4tY49NvY0dAsTK
W1D1vsotwUNQqUwi3f0NBre+WBwMiBvRS/lQxOKVpkjGIhPNDV/UuRXQ7xq1438n
VhAyWstEw9cmCq8DI9uKQg4FBqhozVdZANBz7E2p9gy5pD7B5wMo9Gg8xk9pAUht
TH72hqH7QE1Y+jmht+kUoWnp9tC1HxG6SDmjbvs8rbLRDTwGoUJLf4LxuZ2KlKDG
YFxDLgVGbmppSs6fF1U71vdWTDOf20DIsm8O5uD41c8lFkQQkf7g95sGsUl8fDJx
4Vwax7246j0ZNfBKLrUMAeGTh/oJGyu/m4VxoTqOTr7GkOiIv7e+t5WYAipedMwh
QYVRQRW/9z4kCQWNxQ7iRrN9KcKYpYvMjtP5OhsiI9RChiEmiEBlKY0rbfBQSLhK
SSU9arTeo7BwLzyluCocOFXvYznnz58wmdk7X8cMt9cBG+qca3NOjMcWWFZagAam
0Z/vlNCUh1HztliSZHrZIR63b9WZcdnK7WO0BOGRH9AQVz58hwz54syyYY3qLJkK
/KdaWryPugCJKZ42WUfJeQbicHJ+Oua7nsc6+VxGZARFVFqBan9KuTsKFZxxJaHY
XnKqUJmskZgejNq9r+X4MGf2DfVD47mzD+sZinIDTYNxbtKNJJmUkkPx+Iw/6q3k
+dBECpzp8GJZGthtKFk/68a74s5nFIHS6d+eaQr7lamXVmcWfWU0Xd41EfA9KiBP
E69NVH9STzJHEFqdOfIAjR/QZdSN9ES7PtipnuPrYONIJgOrCQo0Wrt77QdGn1KK
qAcC4ZkW0plIn7DIT2SpBHXiwJ0PEv16JGd381rZMtlVQNWoD+0JRU8o28IxGAAR
qLd7l6EeMLXzRPIHaoeJ1HNOFsMmDZE4L0YCQRyz8IckfFHTeeeT3qMAfNjQTAqM
t5sV4tHeFygTerEHkEfQ+S/Bya7g/PiiqUZ20HBG80COioGAyw/PBhgzbXY8AKqv
G/8Wqa0StTHv+B+apJeXgDs5ULnqDWKhFG2Tnw7NhYPiQYDeiltp8vZAPIa6DShB
jBTcwQBZ55xcnmL3rHHCvCd1XGV39Pi9mGzAzCB0HyuoiRUWzazhq/XHKPIk7GaR
wBjqYzFw6FLTBlbuIiDYQBcdNxVhERCWpxbm6qGft6SIh0iSifb9G9xFGOQuzA76
oGIpPHydgETHjFDhMC1JpJDFl3Z7qAbzyl51GOJK+NJQOZrw0ZbWx6DUj537dUZ1
OsARdHxSJNRf+bXFHaaqCTc/DLwibXXYmvUMy4e2WSNVWYAoDX8w/AcBXIB+0GqP
BntaQHSMIGAj9yj24+nfKP7uSN4YoFuawxvNdS1Py2mM0hFnushHxGhx9MI/OL5h
tcEQJvj2Z29o2VmE11lR8Z8TUw+Vxc9puhPQSeuyoMpVrTmp+e5gjuVVr1FdFG0w
WHBFnIWcwTWuU2GGrkI6icHgZ2UWaOrQpJCQdHOq29d5bULTLOQTDWFBjG1dS/mB
xIyu8HaozKOJxIWEPwA4BVQybaZr056X00COZy4WT5HCNvWTermmt8Z+dt8D6CG7
Hdvd94CnjuDij9yiRORR6PXzEELXIgZLshiADimF/OXJAY3Wap05IWsMaX6azj8J
xLBgiuKMYAEgSoTMjdrIOtoIgf+ZMFKLUYz48iUgCrXfk+cTyUFj6hBC0GMaXqZA
nkjTDWv282wyLAuISir1kFBkeFucBgQR7axMZNMZT7eKhuvKNAu/fThu8CFP7fc0
c96hLSu4folVoBQBfW5585lTe4xs3vEqJQomkwtctORHAqKh3XEg8W7vAMysKIAL
wArtqZjP53mdJxTbz44Lu6Jx4dFrYp3jloDnurFU/wp0+k/eK+F+WfD6iJp2jR7i
tJcWuqb3yY5FgS4l1Mcz0EHStqMusOM1vj29/5Jmk6GWAnXXO6mnGEF6EG+dUfPX
16tiPIT5cdD9tcuXmy7yjn4qU2x//mzCNdmIHW/m/TqXS5Md4MjLjOlkp7nb4hbG
MyQIHgBOMlaiefSmFEDhID+ZiW33fr2XQ7AZAnAe3HHsvNDLLKovItAflQiI4SgU
7YZeLLsbatmkERB3sxccbz+TYja1GsV8bT5n/bf9PTZ5lsLBcHHLhbWJFE6cZ2qL
CaP8h1Im2b5smQZg+kaNWnE8eE9x49P2hQ28O4Hzd6wAqd4QFeRL5MrcMUgUo2ay
6LYcA32Il+QM5rZuvXqyZrvUmtZvs3aq3dAqVhq4Z0FRXt4i24u+/eZxpZGnVCNZ
o4yMDFMOI6m4BrbUsGGK2ZvJNTJ9fMwZiMC0onSCoNvKDk/T0naCLYqoECiVxM5Z
1mJdsjeJ2b0TXiP3fPlcgiAMfT5PIXk11HLCJkS2WEVF84uPqF4Dx8qX7adm1R3W
h3LWtbR2UmJoB1ajTjHJvUtQtWJp2Y+dJfwzXA6crDdv5ygmLtT/idJq9cMg62Db
UrSddEH1hgby7M0yDo8p25pcidNeQv12RPEgrWd8vwf3l0ivfZw8+PIPuw9/kk3I
XWQYd7wDJ1QpQqE17nJ/UYAVkrHVH/G/sNwGWmJ1OrZoSAm81oyHesnzqGLle6DF
cUtoA4nb4af8NHNZDj7aSLjm7OsKPrYkDR+OM4PTuUA0GQNgGa86510O3NvqmVfE
dBqMdYYJvWyOTLjUJ+onyoQOT/ngmXNK7Q/IKDtg6tQlaGIF0hJWiVdh/s224CGR
R18WSzEnfqKGAScDAjvC2XHIPd34QKdU2PWQAEZXGPdCCzicjvEqtHgrDbYkXTwV
Zpc6w7rYviCz2TJr94tKKuEayJp44FlM/E+rtW5ZvJAKnay3UWF3dLizbRKgYuKZ
pHnuKJ5fSRFmWT1VW1U50x+1JmtGRJJxHGHQ1Onxm3RqSmLPnx538fK1L9CHAasG
wcQsW2wX9wYQkQs+sSB8W+iCaeYQH2Gndv+f4i+XRPRPIoubWnO+7eLPvHQppGBA
FMfrENZVo9WJu0AvSebVBcSfZeXvc9eAT2FzGj9ochyi+jq2olXzrz6Qdpf3smkn
3ZjGtmFCjm24pMq8HUcIg6/cAHqymDLxMKtL/SWeY4WmUCwM9Flr1e8rGYR4Sb41
frqZaJGD1mVzg/SBWHqndZRi9r5qi+jMlhQ3Z/7yHakcRRRyOfydyfsbv1xHBBwU
KeqTNW75vQOT+hqdQI01SJxqKiZxIkIADhvRJqKWh50OC3L5Ff8FNbTwBS4lKtWR
D/iXnb2WQBHyUnccHIzVScMpoMB6K3gzz/1Jo0QvS1mBHBFUEKAp0FHfewLmbYfd
z73ebQ8YE7J3ES0ZWtetAcD9eVN5ay9r4V7BDbNnqQWH7satlgHNYfixmoPTph6P
cq2EeLTZ26XrMU2W8/GMM9Y/qDYgAFNVXlEXjCyNRsn7nduPIZnRmWXnTJecFK2O
LZEnqcetvFVIg/rgb4CWar9SzlOBq5s/oY1O73GsvYHpKF+EUdto7eKJT/SdBvkC
pBbkjuCsSTTcsVv4Y5yOO3TKhKn7dGwtOm3HRf4/Oi7851fZYyT1j+GrByd30Q4S
TcSxVfCDK0vqYJACiQXU1bbTatLQ21bXWrXn3qqmkJUVainQTs0wD/ib4UVJJqEp
QD9mC1V43SsxpkS6KsPMiS8hA+jlmR/E2N0tACayRviPMas8wmwfLCrsLMQGYr71
PO4ep/IUWCj1YgAM6U6m51D1s+lcTXr4XbrgOhkL15q2iHCPNMTUOXMTzrWTmih/
Fms5+ndfwZ3dckW2V/w7CzfTEjJGAAZGDplz/qHCrJCyyOvW6M7IULvLPAf5pf0R
QVRpBwGSUehHRgIV/9YW5HYXDRnQH4OPON4Wb7bqJHvlB8IG343PvyiEg+VCJlz2
bmbXJH5PNaGY7Z+NrG/n1Zj660g3MipWZKnnQ+xwOnjLtU7sO2uKTEOxeA3gJrvf
rrt+GH8Vq8G3qFU0dqwBz9lxKWbMorKdGpGf2hcsHNzR08BWVFzgn8EzdNJiMmVi
4yNbCHmm/UgUnWZK/v92lBSr3C1F9qBA0qMc6wwWxB/Vu/sYk3SeaPg7CsYBOsul
Wvb4rlzf8urDS9xrgV+lff8jnXXTlMJumpSm5mMivyYu5TGIm/wXQC+TTP5yukfq
Uy0EF3LPZ4KfiS0VCUNrlx1pFcYVVYnZTqoNLjzIt2TMDbCBFygbSgl/7bWLsP5s
CYR2/Joz8Nh4bTlEyfKXFYwP4N3DZgORuTInVE2Og2MATedWvfZ8XSii567SSu3E
g/c3+D61f9Sd7ebFlLb0RGKMfj9yPAaE7FLuWQYWkLmZ1g2tTRqbqnmLNCVj0uFG
/Z7DWe5jj1nNDLGSyX88nHElyLAfiTvCbiGO0MFGjRlbl3kFWv3Hnbc3IYy1SlBH
FAnZT5MNHUGksnSBudXQ7XMDt1RVwDE1izFMI1bJTkgACBberWStuO65YMceHEaq
MDE1H6YDC5c3zN8dQTcpXool07SxHB3n3PyYi/4uhrhjWIr+PlWkmPmOVxn6UrAl
nGNojt83VxidjqiOeHaox8c3CiBIvzdvjTNFh9zGat8IK4BVRQ0mmoAidWswur1x
XAOI3bNOjtLtC9sk2y1nXuaemY43o6UJxaK7Lkvmt67fsVysAMAllMk2/hZXpqOY
H7PDTUwOWcANOuUPHpqfrhalXwGJURTMRkroWsnYFftO/+GeDbrKk3hpTN9xrD9e
htsggT8zZGh/AU+qRlmZGEyFeFG630Az4HP8a4RJJf01LxkDJHr+tRzQW0OuNg5l
NUTjGXkLzlQqTOpSkSqFQukPtb96RptSiJZq72u8lBcrP1jBGBH4F5vyNSp7sNgN
uEUXU0ZbUX4MMNb15Ra83+sRIdqIz0xD2NypJxnQdOkfnf02taCRKkIMa+lPRqHF
uaBsK4+ZVH7DyKWRXRLmuJOFWZNx6dXjVJWVUYFjQiEdRU3A/YqztIxd5Ehceelv
g/jPw60Kxfud6ESg8DZiXqUN3bGgi3AqCOVZf4vjcbSGIV7rVB5saaugnVIrO2a6
fg+ViWAkYauKouYMcFSEwYektFLmu7tTpI1Q7bbTnhXPn3N+WGf72NDZEITVD6t8
PvEx+askjdA/aQeRf18Oi+Zy8oA0Ycz/tHXtG+/Y9dBBVcmCRM9SX+bv1sZ57ACU
8Y69GjYqw6Yzm1e3kV/7QUJaPlQRUOxr+IRsHg0Fo+u2KcGT5K04pAwyYCySStRd
x6YVvyvMjbUC3d6MuFYxRhmggrZs3KdeF5OarMYlZL0iQvPw42MqhtS5O/ht9RKJ
/Foal8jc4EDsmOqCJrvUnQ34nqwjAiZLxKa4/NNY4Fp4pXVkDl8U+nuQPGdabecC
mAewkySlkBhihXgm0oMhgFYfScspsIFzr4/mBfffxziw8kOOY1D24KvmkxK+kpdq
k+gbiq9xcblSyqzVP5EKI1anuM0V9MulHCFPcbeLYRbF0ZAqZoLlac0/MvrA0Nqt
WkTXazkFDRmYHGAaZ55gbReI+4VkxdqCFtf1xQo7gt7tjbU88Rphh7do5tP5vrqv
SeVz3x/9pkwWQk6XHESGp0LghhgCwBRZDDc22XiALihk/rF551hcJRH1Q0vsh3QA
z9FlUB2q6mZHMR5LIzn62hh0uOLi8yC1CDDW8qeXWwaNyzO/UETF11x3ZOy1+eF3
2lCszGpNqL5rgb5PGJMsvKetZWs70wGuFjB2Kf1LoEzdJpfEeTeJpDCHByZ8m4Uw
bJD6YCJ8BQaFFuFSINBPhNTjsBoNsNccTUOWUDZPkz1SMstfS9BN1ElG7DH+RPLE
OjeoLK2FqwBRZ9/RRU9k2vLW1cfrU5/r2Ln8MmJAs9ouPCCZzIXrCdAWlqUxUHWJ
iDC3AHKm9FEy6bT5Wv/c2SpazQ4fRip3kcdgrpzj7tb9ogq/srYZe5fb1jI/s7da
Ig5O/YBSjUP0C5WXMy/B5hNP2Pn6T+k5jNJuS/302f2BcNSwYipqPirqkWPjOLQR
gTu64IdSncX2IOjc6TLkxqdWJ9SfdLvh0V6BJupYcldud1dKj/5N73xH+7C/bmVQ
L1xsHQOxqkB89m0aQpxu2MpdoRizzZEuP1xKu0k2IGs92pKwQ4V/lxCqIMLfO4jn
9v/vAm8oyMzUl3z06T/DF7+yidZv11BMDJRu3dUXG/yQinHCOyMOS29BVh/o1JKn
2CoMHf1Pom9opnhq/Px4J3RvlN+aozd/awbDkAWBi0f8JA4gSubB4Q/iMiTVsJL/
4Nni+DwSd9cynmg3QTy30MYNmVpfNGLxItiHr+5j8PYR4K5TbIciFlPyzeTpAiCd
+2nmpgVWo8miTsvPDk//8kCHaH5dP1B3VFXOCQaiofHkEXUXA9txSI7qtg97Us+u
kqdHtKwRr6H20nLkvmXYiGHwuASoaVNN6DEZZNtIHY4aXH9uOOlLI1DBu9hongez
nYtGv4wOIzsek6BDE408x20iPVTBUaQ8d6CckCJOaLjSTYCYCqikH1ROAIZHk6pB
Nee7IVn+95sA9DRUNm+m6nANTKzRDY5na+kcnrxKLPA7dNLrvdq/aD5d16nAgTxC
q8Vl8MjFiBCUByMdleOw5Ax/BpsWi1yBNAe9PcBacLsivaIlyNZzx93/+Kv6q1X6
pfFcOdJmFvyXFfBEyGHC5Vp42r368rmZz+xqAQqliC3AzQa39a8T0yQG4qjphlBh
xctK0nWEvK0FrXokNzG65YuKt1/kI3Dqeas0WuWfSMSww+NB96L/prSuhySZW75d
uHOcfeRvaPk373IW0gDZF6zeppknGW5XLfojj7YOwyEpn/+T2do7YrDrQixugEgg
jA1oPM38k8ZTweFB8DkQZOduDkb9oxONEVOV3ZyMH+71GlYwyvoMqvmS5qPb+hKI
VaujknpRIuNMXqpWSKW1wS3UiTbDqA3Bi+162VjnpIkoOmcq5T0KVUszStYZcuZ+
QVBXt43veJMBBmxJuvxAcDy0m0zEH4Ok/IAX6mxvQfx8tn9dW0K3teaXo883RVSp
GomQRcXEEdhJGy1ey7Rk/cCw9rilL6/Czgi2vasAu1t9ACDxyuFl4ej2D0o21d30
MA3Sic5ZwYKofcE5XlZ9c0QWGgZDe+XMy3oy4inBIRGPPK0OfPpEZMrzYSDFfXUv
pz0qgwiamz5ldy4gbK1RXYpd2FM7i8eSe+DEFltVMk/yqPeEbBzGTVHNXzlg8fed
2DofyHPIod6OmwiAyQCpRxiklZ79dYwTNSqV8O1nUC6ZEjtIV2D0xkMFKT2TM/Rb
QvYTjkeORrFpKDgWnxNQh3MiY4X678O39D1Dd6J0tlaiOHbeAnVVWzG5D41VN4o2
GHBtrAQXed4E9BndNEyvNo+ipsXyBVL8PVk06a4Ie0gJLyMyqqQ8/OYiUSOYN4hB
DDlxO+bT3sWpKDaGlM0KwGeMM/ypCGR5AhM/4uf+pv5sOsp0LwysMpf8e04vDsRX
n7gyCCUw2fqEHyOdxNqloR52hMBGoNEg4g1+mudct/qC8c2mRblZ89V4UapiH+ak
lrbEREyAMqqfU6QXiGQYoEbe8/2gqvS3gWs+JGYxggwMhomjcO4+5K4ydxiiM3bk
Ec38AFjbkFJQvlNIU03PfUu/s3++ks2zl/PX9YTZIbUEaw3Tw55fLKPKdRugdddj
Hb/y2o8e+uKmykRintdvs/uEfI5pWyv69W2VpkhWhh9qYKIGaxJE/IzzGsNZnnKA
1memKtPTYvjoUE3T+1avgL6ykmjDBtWQjrbb8+FZAf1NMgmNy1K29WX+f50YTroS
y0U3wpv7jZkCVivfcO1oj+Zq/EyIRsVdubngoOcShP/4xs1krS65Wf6ryxax3SWY
SFVELCsrKLLT835qYw58wcK25pVKXpfK/GHbcKLHvjyky8DXyRFbzWT0gswPfb0o
e/8Vqcvgw2fVce4MixBc93oR/hRuxuiX0AQ9h7GGTv+3beR1b1fX+D7ibiRjHD8s
xIeDtpm8FQEd/MiSvrNRC0R3pPCcHVtXGbNReICYGW/B1lvcphOFwdTPSDoVNWDg
gUF2viqH7CrjCI2djXnpWiY4f33IjUzJpi3tr4jrBw0H+HvKdUGiO0+CdEAs9o0R
zLXcSzDD1Us3oAjTs3OjOSR1afXAn1s16PJyRmT4GvnHHX0nTVIMITrddGoLTzfN
3pESCbD+RfmlkY77VBO8ZHwJfpInm/JW4eLhqTfSnY+t1+OeHbKW/8kgMF7cjPnc
XUBKTncYYboPIaVyPR1/q+6x5VuD0YDPqGRL3Pr3lx4s0sdMxJ4tvadghRMuoohl
CccRl71Yoa9VSdNw/RIOiSXbIpe5hRirUUTRoTS3xNF0ZSWaLeEPDvgpdupE7T4u
Sux4NHPYvm/YpkH0uiSdqMdRlbxwrdR+e2xLTPISyaMxOrLSaHRIJVGSSypgKaiH
XKxnsw1iNliswXTq7MG87eK394WQXwUKgJZYvOzzJzfpqyyyIZR3esPQmtgFnpAe
sHZlHyeZVG24kDOIBnR8Dt6Jy8FMtpFt81OpkGuoPQv2fWDOcVLcrhZqeWcS1zdx
tyRBOCEdUBLMJ4nrkKu2W2Veyd3/LDY2ZJDEH8USgYlYJ6/Kv+9NzT1hU7aw3Tze
WraiskQjhwkSOs03XY3gRzwiB2tr/3nDL7FGPIaHHXiYli7FF+MObD9sXH6WDcq2
JxftFePkjMtXTmubfjz8SK54ARFGwKjpvpg8lqpUIMYA+2gi43TUNQNvQtuNLKbj
XAFwZLwXiDLniSlFKnEcNJfRj1HBqReyC2mI8VaeJIXm+Ub59oU2xXZSfX9cWmH8
AtatU1tFZhceIL/QSpStj2ZlQpmOlUhhZauuMLLpnb5Ozi54UBOlYxUO/dO49lil
7dwZ+Ox4LyrUQb2v6EL7t6fZjRvwMJKpGgcncm8hxuLrd2RCQX9Yv6ntpjZZwSf0
pSc84uxqStoloH1M56Wkmup+0CczUPWFvz+Z3rcz8ZKGR1a0euPi+QGKiFcJjEkI
8WIMORd1N8HMhqwPyyZ784l5bSWJvT75Mun+e+QdYLmncnLQAD3D+IY6+EkdKW5O
EutFMWg3ITWQeObhkmMu9hVLQaYfUInV1pD/BzH2yzgEa2pfOvn+e8TZOtZ+DvJ8
4a130OaVjuA46V6/TsCHHWm4uKR52dXKa5Oe0+3GsFqpIaCYLroNtmcpC1x597Ms
iW1TshCptPSh8fByLbMsi+0YhBzVvAJJbmX+OT1Mh2tqFA9gKO6KtUYP54/iePya
Y8j1G1lD8Q+ZqxriVdbQyP4EzcFifW9E+uMxutPcdnwXSEkX8CyiJ2pkCByhU0T/
KKIxE3XLmYwaEV/I2WrY4joCqpJsatGEPtsoIPdi0r3DSziToLGU3fczWYO9QBSV
A2SE4lXdFUgQh6y2MoBMFF4vRRvyfGuvYpc2gyotYoW3GXrnYl5MRL1p3ta7J364
aUx/x6pNhYRu400+QUq+qbd+O0hOawOkZjxfGEhgWxJpaNbC9SMIKfA1LP/v1zPr
6UOqIPFi6XsBWbthtLlWXZiC0gLCttTMLdHdGMuA+zBlpgwXEAKct4uKpo5sI9Dp
snmZtYEE/aiEtJy5+t6mE3IoK+9HdxWkwiuwQe9praNz04slQztEnrFLYGgG3aqi
qOryFyjJ1Bg3YPxjT1Iqw8846PtNo1YkV1ED7M3mdEAI5neMQTEsr6KmB36ap0tn
YCq7nCexycLbeAIoKYnSCOvxgZTb9Bhdr+xYFj1R2n4/70pL/THXtefAxLpdlvrt
xGv8bGnYFjuNAZLU/F4w1DCRibtd050gBL3EgFp87eRoG94kT3Tuhakp8kCZVnnt
neDDTeplgbVv/lcvwW1hhzPfs2qsCyaqFEt1F0MMRSsaOsIvyDQ443UcapbNcsPO
pWJltdFe2Oij+i/bm4X/imDSRz68hbJrJnw8ZzA6dPHIsTTaPPq91i8GR8dyxvfg
WiovK6d1nKqQGAOS8cilhlKDuSJOPyDeEAUe/37Z2xqJkKrjyFl0erUPtOqMGsVJ
vp2pkQfKH7XZECmAwhnOJNcEBIB+nxDU198EQiXaahQpTwx+HuNNY8MGCukIubA8
UhPFel+s4LOip9EnqxYQxK7XZp76+BXgWnqcOQ2HT1MPR07Si0kDSqvRpUm54VNy
ohhI9qs1ig5IALJzY38gDtAUSi1v0Yfuc9b+X5SqHqoUWQznN5nvgz5ms5C3DYt3
3L5KVzo/nsYylIdM1ZXux+3rwsAOhqwdGDeKTPRvxBDNSbWmHvaObaTL0mF21cmp
PDpB3Uoxza32Q6byJQ7YYuRbMPLP2uLQp8G8wThhPUhKqhIckk/OP4vMoM3+tzU1
gY7c4ja/FVx/228fyIt4fIhv/gPd+jRRiGTON+i5juK5oYLm7MYpXPc3fkcEqX/D
lmDEwfCT2SruqxT+/SjUvuY1Ibt5/4mXv+/sLK4zO9bbANJdN91+1V5LNDWj2EtA
FcHOODx5m1T6L31X2gVeUK/fZk+gny5+RfoXdrMvLZWzZpqfX4UMjwKfDjewNscd
tWKwaQ4fGI/OCPlzWPrC8T4qmorJdoaQbXLRPUI8k0Sx+E/GXSyD6risVwjfRzsx
uyGjiqXrNnQB7LDcX28E9w/YBO0S3H1A1ODyvC0Zy+FkWoUx6v160KtwPcl6YOOi
x6hSI4i3uX/evfjznb+Jt2Q7NRYujx58WAw8kuZJdojE8jkiyEwkucBuH9QvVjhe
hhVR6ATn7IEq2yJkR7/3/+6Mmju39dnBYz9SkA38lRF2SQr2UivGvnQb+6SgTjrC
I/iLYFdBSXSwL5Ob6aEcfyEDdXsY/m7BAhG+X4oB6EQprBfXYM2MHsEnX1ZBlJG1
rB1hiP7YUThhXP+k0zs3cNtnAjx1dKpomRUD7UlziLLOrZd9qkZ9muusYTIQfP69
nSo851GYMnRPkE3RofKpaXrqqnap4L4SuMJcAFfamHxZ+Jyp7/EGFN45Fr9mdZyt
fWyI0OHltJHMELBmWUQ5pLbuhvr5zT8BhSuBGdJampWeO5yM2QL+ypoXHHTkIXTs
s/SoHvsZIMnhrCRMMPRjGQwsNAzuF7KRMv92rSKOfG7cc+mYD4geLaJPbWfKZ38C
aROhu8m4C/HtKU6lsdwXsfCdvr/lwiSJ1XhdLn3Qhz/ovWNSnw4Mdp7YtM+INdsE
HXofT/nlHiPmA3UXSkQ8c8hdvZAVT08HMZgfAGpsaV3toohAvwnHZsbEWtqX7Z4j
Y7WUnSdk2akvOz7EZ5TioQVuvjKtgEWemVSb7CrBNBw/r4UGUUw2tgegnozjgeDa
x/hgb7c+v/ivg9pa7JTxAgbneHgxhFnzKRMGf8qryXdvlkqjj/lBAEx6II2gsebr
E3485NmqL25BjS1zGymN3r13LmUA3Um5ohO8s/Ll/VzgXlNXLXVh2+MpeJjhXd9I
/KpOiri6xhnLiAKprBDpjqU45BhabWxOiy5GlPuflGVCEhhIxuKGxamD3jKETZ0l
cYKiOU3IXc5q/Ua4aSVmevq3x4BoUgT7LtR5pYQR2X5Lijid9iXYIdf2OT/e11fi
lJSCBFpQTC5+vsOkO4bS8CeU/JN1q88+6NebCPZH7B8ZDHAAJh2w2RJdO999bhcA
ippLYLIJWV4TqO1Fk7iBwkW4x/xLDKFgJzsSi6WRnhB7kg5ZbpHamw/C84o4c/bK
KaXR03ALHorZdvu2OegIhtpWQGJ2uCoObWBYQnlnGhedKCtWyW5cmPmUjWyfOtA9
7zCr8iYdKkWZug6j1WFZFGCwNcDiQkYLiaazv9PnDiPwzMAMNpIXPL7GqYdb1w/+
Horokw8W5362Tdkcvh7saDyz9sOeBx9tipJNsXZE2NFa8RzsSkl+c4zhI7oK5RD7
`pragma protect end_protected
