// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:03 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GVLy4UYw4s1+Hb30+yGl2bKtUuoXrZI6sH4kDbnnYFUejHmvF8Qs5mZmpoy35wkP
4yADF8jy9+VxsKxIz9l1F06MbM5Bo39c5fEGNh9e6cuCSQ7xK94qUMCPZPvdzWMn
ry8T4O8iHRyOipu3SKzUFH2o1AwZ3zgvkUPnC1ydEKE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12928)
n/eYg0XKC6xWfu1o0N2sax9ps0y2p1jKHPSYKy5IKYJGmQq+06Wbr57dkztrsKrI
Gfygi07nIIrumiMJLRhEdcAHIKgpyVthun6ocKqfwrZUXYsEVmbKCpTXdfIcsTh6
XTgqa7WTuNJMSEBVqB3kmoTIUs4ADwjxYnu3c59320/dab5tHk+wckj2eDOBfI7W
Q6zR9dhxYE0tfnRmweFl2yRCwv9sTzBrEi/15xoRD6f4fdyLsTQM5Y8pj0ZP6Hjb
pwIi3QYi0vgQ2h5bgcaj1VUxefmy1BYT16uRB+iLw0o5mgnVJ/C90HF0A8ujZEbA
waTeYzHuG8WqVVrnTVOtqOoiw2qigAOFZOchrMC8Ujc/204am0jIFJv1wf4k+7Jb
Bzslm8x5UHIqPAHk1XlmLgFAnYtBDMBm2823Lb4O4eeovnMvcUeMJlwIcWVttzqG
kiTGoBazbGCJD+ARhvGke97U1uIn896QA/Vtgx32r4R6MtwWytC36L/ev4JGV4dc
D9HgBL7/4yQVEv/2XTQBjMfGZgggKU3EsPeiJIYy5QyZ2R1Iq0bPd9BOY3xAWzs7
Nl9CXfOerRsl2l+PmQX97gPWAanl2I4CyUQT01Mh6eldeg1Rlw8TQSZv1/IfFMeH
8y5OETAi0dGtXVGXb3weSj8DcAYRCw3p91ADyyneXpnV+USKxuUMlCICFCeoQGZG
kd7/feF99XE5ZhHlgJGEnB6ZSNLU7ty9KiTJIqs1Gl4CNghf6G1iTnDTSMhJ9otW
11wiuwfC8C1+enycY6ckGjzbqHv0E3PPrwleS9aNorpQX+GTF8vmqVo6Fx/1/S0m
R8+cebjj1YlOm2pZp2bNxUhn/o4a/A47MpPkxyxDQF6f33NVYZZSiUTmk8WAMu+u
EmjSur0Zdh1GWyMuF68SucDgqPPzBvdi7Iv3sZqIE/64ImO1bXygEqSy2TwUqKfi
wfQlxjs0VTeIk3oDG6xdB39OvH/odI0klOthOqjTAN6wPU4BD57KBk3QeSnjYfGs
bzRS3BHiYTiUPNNFzqjz81I5oMhOUYgCCMJWLldFbTYZw0fJrWiyxS7eBMWpXFpG
a8bBBo26FgO6tigOr/Q8QFIvrh1HNZBrBA8e8y210KbpUFB0qanMacd+eZY10L5F
nnkhvr8TVrvDD4hFdwaUUSCEM+VEbzDLVwvk4r0qdWU7+9QulVOlQvYgnpmNtiHf
SSfu4C0s/6oC/iTB4wZkDqAGeCdKVzrocqv++b+hUICw5nMs255a/SRvgx5EZNMr
PNh1arLNRJNheSh5yM2x+H/Ynw1t+4pBl+vFaDe2vohiRoJIJrFMfvRswPzdwqze
rEAN5NFsAkKbvg2Cso7gzglzHgB4vn3uTlti0sBz7vTl0pwOgvkKyEPR6JkNH1cU
6weZ0F2j0+gi1jVMS/BYGkrFgwJCM54xtdoGQ613TQZbhRY00LsZUHCDXvAmjKir
ZjTKvcv+GE4U5D0SiKLYcuFoEuWmUJrZKlsPGR+uS+vWVnRDIv6Pz576cUn681kM
psvK261oMw1Zy3Fz4Wkfvs7HFB7Q9faJD1ymYt0V/yRuu2/ByhKD8cOUUS3dWzUA
4RGq4WWh0V4Atb8JGMymiUwbL1tHF1qRBaD2xhyHBZj/q+IpC+mk+fT3xeqbNek/
rG9JK3mPv6JmNjRknIya6aUz3HP69zjGEcs2n0BnECHiSJyFZfQ3JBnldPBCeY5N
Vh4mzZgb4qsGqQGuFVxHUDnWF4rJc91Mhk6tp1ncaU2EhBxuu74BSS+LlqMU+71R
4DQgryoDtFtIRlQaGLt8BAFYE1pJiYGIKff+26z4j/45W2HizXhB34BRksvV2yWF
Pg0Vu9n5y2J3m7jMRMtxGVTIM+fuVrbAKaR6tBPuApWTe5ct7UrmOWZUk/8mWxgB
Zupy1xe/plMvlb8t6069sOF/u51gmNfaKWI+lDsFu2u4YytA/ZMH/HnTA4+mHVXt
3rrTesfov9iruPeNaBqoC6GB2/s/gxtriGEa5zPXDljycPYHxveccGNM3K0X9HjK
qtqnAzTO6NJ+YrlleZJry11QAAzb+PupU2XeS93InY0kfxwlvMnG14AZN7WhQ/QB
v7omQbXRAJrDP3thklSKPoVFZWX5Hg1bvEIi9Mg6x/GCr7WZtJ66FTAAtdWCqQ2e
VipRV6hm+vtCAxbb0YTLL7MVl9KgJFPGxelsKiHC9OGsjfMaBsSFanh2GUDhutZ5
2ye5PrOR7bbqO8+FB3g8k8pRwfRiDg+Woc6d3+C0kbRZV7HccYmVVnqV5k/96iCI
bGdoX2XsluajNW9tvODfgGDR09pMihJz+PELsBEhrWahu6vf05hg66bH+2K7CX2C
bR6sUcHm8JoqVSlexR7P1GkfB5rbJ2IFJ8kKd7pcrAzlSvlkEvvmJdkX/KQudFwW
cpHmG0zLpIlP6wnqhTMZE8zSHPi1FLyOpm/s36qRxGoPYX8DKTZ8+9J0nVX8myVU
Fu7yPwEF1A9XaNaP2IUhUNXLDZ/+h6v1OmcE67dwi0ew7XlA55zRkoJILnv2W/AT
U4bKxCjj7GjjEKOylbweeHpHVUpPHWm0W6AigrdnBF2QKZ4N6hk2U9dToojKb+Oq
U3tItz1Phtk032cNDAQ8+eyuSyLY6in1oOwVJQs4oq53Pc/B+bmFAdJQz4fU5WzW
whJSry06+Cr07oOGKTgahQc0PtsZRQAo1it+cqNGLgpDFrGxdgFi1435zErDpLVl
3Evl6QbBKqeLdOZ5EJJZb7Mlvnr+f7xPkO+XpRruNWWMggog+GK/6dtL0DeDDrdz
YfmoEG8kV0Ab3L8UtBF7mNUGWw8nUoRAJrXlwqZxJlOTC6y/Du8vC8BleUV/N/IP
b7zxTtJirSrAc8heVaKPxxABUJQwGLWwtLY43pcmiWs0AC9gHvyQbAPp1qW5/1yz
hNJSgdhSL1k5MLHgIrI2G6c4ShTLwFDL/NWkau868EnfzBIrdBW3sWtH2JriC/ZQ
/x4GT2I3vy2l/DGI2V1pKPCsNBPPJV+5MVG1IYdmxYAfxg6JLc/5Ak/XlI/09tK0
QtEeXb7X+Yg7cqEYw/cjYyGntq1YIgyqFEJdB93ERXJRpT3uttN+872MFiEXA4ib
SY1Q4DxhnUQeMdMjwdU66tgbWxosocxIRrtqNwy/7D08ItE74KJRBUXS/KwkJegI
RY4qynn6/HXkpm68cVQUn1iELhjknJQ19otrnRYBhn4NK9RnNgv7CRXikEhJrBFK
WeizkOeWOSU0GWuO6MCBPUGhAeSgvP74HcYVWsyjmkqvkCxiQekSa+GlOecSMye6
xdSicN2GMNqmpT5pnlGUFy8QtyUs7Ii+SgkNaaezGqltJAb+bSHA03PFzFqEDFQP
KWEGJl0Tj6qV3Q4NgtqifVfOiAQTkMtD4UBT4pvRJ0l8qkcyO/SLVdbbPGO2qR5i
B3qZdtaHLagWTVZjQfbuRSJ4rnSusH5Ss7uoRyJGK/p6l+POgoirZzL3yiO9uWN5
MjzvKzzie64oUES2kpjFFeGKPztlWgb4NEUWzu8po2pSE/Z0vzuPJJe6FfXNIbRE
bH1VmvV/BlR7MzclTYhk81L62ANzU8oEIPWppaFONvWFfyFRD6u7GYLhzpuOTbGX
41+blGlXNOMJ7mv+KUm6mctFxhmZHele6XR+J4W7zaVIejLuLtYBnxItFSeLrk9D
HN/almTu5phnC/usJjVdarkD180K01a6CerlEZZjd5fnOGTGzNqcPlRGmf8PTcUG
IHq2Cy6qSPkqqKQUNqofsMnUZOcvnAFCvj08fihV2hzAkyk4OyG5CEmbPASVxzyX
rEDDbOdBSryIoh1XQD3EN/TwffoOTZqWeJWFziG22v4ejaeesbNK5MHPNMxdu3Sv
OudJoJz61mnD/LgQiex3ZSg2rMgPNQ18/I//3zXLfPaGzydvB2ovRAZSbpSTgJ8I
8i7FOVZdtcBmIenb+PHmDBQBJTouPAmvMBJ31gMn5iJW5qcTgNwg+z93pH4JSxO8
j17G69VwD1XvrphIzvlHKyr5MizxkHkpFQr3f1poztNiL0lgbPCru4eUI7/F393s
FMrZwPq1LuNbF+pcjkSQ1wTXkc8ONb3YrHJvGkW8nS2Z/M/pUPI/sxWrHpbariRI
io2kDuFgF+uz6FW5X1eTei0ZBryItwdU2QEI5//oDxYiWSNQ9zZXRH9z8pNuZjf8
8cydJJpWJY3QxASzRCD8DD3aZB2DZXW7EgfkYK3pWBP/g+jdaLj06d1UUwNmPrjx
X/Ut6zeCq5K5z7O23oCgWTpTlki8miaU/yyRZj7s1He2uYKR2KLZdeJjZiC7Ei3F
xDJY4iJiTyJeh4dMssh0lIg8pCWWqUqWoE8S38xP5j2Go+Tf/6zddtFtJTXf3p+Q
uTw7PRByYBpt6tbPU7bVSYKeOrQdGK9I4N8Ed21s+gtopJaOUsrwvd3sHbshiE6A
cBLsyoHxmcE+fdelnjBrvYbEzcRyvrb5/ApDjjsYRsqQdrhll2zmX3SWD4ZpDs0c
FB8zw2CbvooN4VlrUH3Pg7Qs6KQJ6krAZNAwOeJJwh2rdRUwrTFWJ3pjWjGas30T
DQquYysgFFOTbt7+KYYYzIP59VV1OEWiVBcZS7N16I2LDj9eG/Q9wpCx+SE54ghr
04ZpJiSBEW8PtPKaFhe4y5KCAp0su55Oz8JDfsLGk8N0giEau+bWaN7m0Nf2puxm
/J2ZuaavnwhHAr3pCpMDTzzNsI5ePh20ykBq8CxdtTN5GUmRYWW4lZH04FkgYO97
0N/rNkz57UyHMnYTJgzk+ulPWxhatSJBUQCpCPIZ45pYUz+H9Y+PJxFr4ulXKOu/
oo4HToC4cO8FQnMRMcy8RAatNzNIsS6zQ5INHauLHnQqGiD8vkkDwj6DPHGIJhIL
uVDPNDD3AeZ/NkD7hC5m0MmjEkcwB20kZagkmupRl5kffzDqcVWTFUIqDFgcNsfT
TnjHgDAyW2vQG45ZztB7qpTc2Kf8YBYW0p/QXlZ7LaTNzUaLVqPYjKLExGjRQT9n
PzpI+B/rjJMUnf+sFXK4W6eGzo/chrh7m82Jka6ilMTcIN3K7oKWEP9+Kqlx3D4n
/pF0oUBLpXlDhXzAK0VKPVp2o/3qN8ArLXtj+nXX1WybjsQoSezeS1vB7nS9Q9Pr
Jvm+xQCD/3c09eQwnlN94d3UA7HqYpanSSrc1WBDxjztiBCVGzEKf1s4eQV62XrE
siZxyKjHcqHVOzwRov/1e5IR2Sz2wEF4UXH1264qx0EPktEEfmfpeoWP1kC3rTms
K5+QbKMM87t2tVwsQD4fn089lpoFBYXnSboZhydh5JBS4H6RL72zBhn+NNSNvLPt
JbY9B+W6vqnfeqy3LJIXH/OSXYctBwMByJmnqWcGpwzgnMKi/YQwvCC9wF7ubiBD
h2FG5b4OjTWMTPYk1Ab6dcqR1Qp+xJ4KRJue3ESnMwYA6YaPr5MzDvebZVwZ5q9F
K5dkHueL+/Qa6ch9EnKUOHnWwXp1bYVuqlJ1IfEKqdA7m6G8ah2c+wFrsD5AOQk4
WvsvXr5ei5wPpc2CgH5C9xsbGrGtL4KWZuKC9hVJW50qGVNfSXpNjBhDTQ0aYlf6
hhNNufqY/JDcgE7FEB+1Img24Jl6+Q5NMQX/WCglMsZCQ9ZCdO5wDapA6MzzvO8/
sNv4pDoH+JnWm5OSI9ElckU2vx2MVtxOO9hvcZqjunIlalsr4pjGraj/jsZSGfeQ
eMBQPfdQLqvfHgs1zKaqnOY0A0xO3BQkTPiogjq9Iel8mahfAULByHxz1r3Z8592
Zk6vu4n72zOuUNq7n7wBj0vy4ziHbFyfI5wBkeFOYIhP/GneyVKihTBxg+Jcg1LS
555976lzvtcifJsHtvK/iBVlFIKVkCIQZ3A6UXQgb6sXW+LDOffPXLVHpTu612Hi
t9paHqQZrD3k3uY+8Cy+KFMJH8w+UpVbXVh/vvpnsx6Cr2ZhyF/9gnbpBrpw7y9L
fQW10JdMuiL8Uw3myoHXBfJ0BwSq3Vjyq66TejpwbXiRvXMzDQQ5/+J0lCeoh7Y0
J9l1BKFYDFliBWKIGoPwTU7HyNzgbMB8D0r8hc/a+qdCjP+PMiBxf+erCEqPI6LT
DUbuuRChXxwoSCkTwsdGhPwzGY1irPrh9tN9gFFoc20McRg2uz4GFMe884i8IhzQ
oeQfh7dGGN6mSzqw7tTnW0IdzaZ8w8TBLQgLcydWS4htUzvrD8k9PPvQobsRWgvH
J1mA6y9y4/4b+WmNQZz/tARcgBStptykxUrtGORO6sOrTVPPMhlunzV+xovabIx0
jOqeyethTlgC7lry6AcIc2i8QBFefh9SirVNZ7tCNiA9bmDjECAs96aDcJVqfMaS
Cg4cQgHJihqDiCJ8LPTv1TTXFg8HgVnk53tonVQOwoJbPZLl0ui7S/yqpoUfevgj
BNwtz3Gj5yh7/a33ctkxojZ1KvxDLy0jirI4CR5kbagouRD/kkB9YXYlfoIpMcys
gBDzRxnxK6ar4UqP2TZf4VkFH+nRyLFWMktwZcGEYtzI28PUP0IIwcd/mRkefbPW
N6DSHLORgiS6RjZjx15Wgl8W20kI7AvvSKPz9X5Rp5PzfJABLagJyz3Rh6/hZuGN
1qbtMd43xEOhTPuEM7KL5qJOMPziRbDk3LaOLCl+HkpX0QimFmbxC8xG9E9GpgH5
ANbfWL4wcKxhySKNR50HfiX9uisjEuWYaM8c+4TUyeLh/a75OfYnrsP80E/SXF54
awk+azLWO6YlATf6e5zi0Vyo6srE9AWBo2A/i4T2avdTcWQ+lr0iubxLH15GbMrm
f+zXDcYE4IPvSIw679nriPDvIfqHz6Lcy44VJACf3atv8E7wON+Bm/Mtmrwdc+7D
lURsOcQXDbOXSsb5UPK9FB0bfuur3X7ZqYnW30vZpITyzKm0nkIZsl1nOjJ4U5Bc
JwJo+Q5da8+2pwdjTSrfFW040wV6fXDXbiXV5BIaqig0/6KQEFVvy5R9/chH0hqL
LtTB6gDjCwhRR7I7BY8PSCgWit+OVASs8vpFJiFOSxgLRRe6Pj2rWizavnADTv4i
aOarnev+qx+dFINIWJRyF6LO0PE4jDkdLgkpjExHPTIFEvY/cDrzsrrdxj8WkUvL
bxrsJ7HoaP/diiFNaWccpscyWBpFEQRuctK4j+ZTVaXw7OOwyIN8lOh/HyBsUm2O
PvldZpxvwx/kI+Qn9juNIp3gr2QHsFVX1C/KcuMKajb4lrLKOyzaQZIDqfPWlrDQ
ak4pQ/648MP0HV9unHapU5BOc12EvpeoK5xkIz7bpk+8iHXzFk5gb0SPROw1WM30
o/FoTpDzAvDgpRNdxvFGnjKZyFZDgH2DIh1SZ2Efs2ISTEGb1+BqevATq4H4ZSdP
exM4DFAcK/kTth07CAEp2wlmDb4evy6NmUWPE+W6zUxVXxcgqaiVy7qcZPuCn+bD
P1liY/X0FPNSlTUz5wxEhXrXx8EkaR2DrHA6Xd8eWSYCNCpMbxQ13Yt6sWRNmfn2
sKODKt00Pt8PHkcuQRJhYdLTG8GUAhRQkbtsS4PMHWTCHJ3Gw0NkFMwEXQXXTH6v
O6T8i7oY3sz7ozn0IkRvrEi7bxFlUBEmL4mRJCLCTYlEsDexdZwkVft6hM3/na9E
DbKKFuAT9KooKApLNr8uuLLhaI4+lK+Fo/rb5Czkx1HcR4K+5r4wSmnfSYhts1ga
KKIjUk5VOgZt0YAq4jemnK5YEaxxzn4t5rdpvMd3i2ySq9nvq4cmj0eveQRM9qlK
DrhTUSAqw1Q8xushVin/GeOXIkvrCD4dNQdXU4opeMzeP4N/wTLNW/F+st5mkgth
i2IAkEA1K4ioEW/CEumslljrvLgnO1HXBV/E2ssm0a18rF2VTYiijgKHt9roLlNe
6n32dzg3iVBHThnr5lnkmZToYEaa88yuGri/7BXdfs6SEaXKLIfpnDxvGDuTFMJv
EdqUP8ouxQtRskwLthxlwEG21NumsS6feOpYlB6Gqb7BvTnC/4tFZqw7v9NA+gSg
P4Ggl8qUHyXzmYpqrBGFIa4g/AIcZhq31G/9kyLu7cd8NhNqU5g8zA7uWoiX1jl4
aOFf3rkD0IQ+a+tsAFdf8Fl58WtDrRt5Y3b+wNWtPYQI24jpyAyv2Da60hyYm6e3
feeZ5dTo+942FypWLC9VFzXmdw0gM7UV6397cQNDsltrZr9bcaq0rnvrdJKO6Nf7
VExsmDqom/mPo0sz/Di5rvZIKsYD1X0JHDhHl4qbTLMCgRi7EtwKbxHJB+Pc8mV8
q7jjUYmz+07V36gvhlcKBOBm4dyZ1t9lEzgmffYXgzFo14JBHn80JFZSc41ZSioK
CEfSPBlluiWoybKFVKG4Ba6P4ZwIA1Fp4bbYSgu8+jB9O2mnX8kMj/gc+WJOgGoY
tlwepPQdeSmwfPPBX3GZSyFqYmSJLATSatBHnN3v1BlEkYZ+7EDQKSFUKF5giNB3
XvIWbBQtCDcTKgN3Syix/PCnEWfQJcCgqrboLzq3FfTEJZ6O09Vpey2Uy30/GqCw
S3EDjrFexiRx+vb1HEjKCe9fERQrIM8mANJbGdlctUopI6Jqp/F317W0hRQTXkKi
gDGfBlbrlYCmNnqaRK1mhXuQbmIsxa5sRmjv3BrT0FG9+J85/VrE0V9cuANyANr3
luBwQl6Nl6Q4ZxMrvHIfC4FRSwrwl28Rw5hiJvRAJ46M481+2r7aocGckqtsuRn4
HGzGgwu/swdwtFJtnlKBmAtoIg+S2vQFzB9Sag1/4CJPaRKwJgAVRSorOj5ucLDt
bPZsG+AXeQdIgv+PaRcFjkABzuiCaQd3xNCw6vBOzgJjlZalCEYed8ePAJ4XQp7U
D6u47QktgGyxL+sPJZaXiiPzreGF4cCCgzzyO0ZoM+JetkrPQHpi1HBT8oDWCMBv
6rzIMezBDUOXbBkoRETtI+lc7bOaqaJLhSg3pxgoKEXdUf1LUaZxhI8qP6Y8G7u3
IWuuNed+GBxwupO3p8uFZO32eUGzEwRBas8FUvhHqO2ZvqThVVGYuiCbx5IFLZzU
axcUQ0082QhW0jeWvlsNCJ3GYeLxy9+QAfjQSfi/nzm1GgeZQwHG2dHsOILxNWE9
fqPPeKo6M9ZS/UG+vdrn9SvojtDKoehh7eIscV+mpfr1R8UNuIjC5dVyuk+5affd
Ig7FkpKeReI5EikGbpt3K4Sza2SomhMf8JRrA4Nqqqkee2uVNp2Hju15qElaBx1C
tdB2QqNTWY8xk4bmKt6wa6hx32RRVfjplA4MkyFQP5G9lxSUxRFyOrQnyfU5NGT0
NLB+j80CwXTYBhXHMbpd81Plxo7zFE/PibWPDgv8FMwU1vYSpIi6PoAiTJ0sYEmG
h1qoSuTSkRScyhW3q+HdV1zEqxWHTqEPq7SAOZPtrPxotDvdoVC90PPnAeJ/VeYs
gPn/ma/92zT1aTv11SkVnfnaphRnKZbWskTGugjFafAaPxMUrdrZ+QQQUG/BUNvm
O5kDzxZIspOmupyzfL2NAtvH1naXTjFHTZhuRpQ/095Ji4qqwNvIYVBV2tMg6zRZ
RdpiIleUIx25B8Yy8MFXiTtJunxnBTbZTgLliVUaehZFWr//1k/bknzChWyHOjL+
Q7ohdzqpxsl0Z4AOLRYep+xHFxn908S0jdThj/DuxDHNgFUIFg1UnmGu5TOrtkKc
X4TlZvFadovGWeMVj5aiLvkYlG6pTLOY8OdbRdG/Mi7NXJSTBsjxYACxtK+tALRp
jNKjH46Tby2b1WM5SqAI80o6V0PFNBolyC3fxHa9zXpi2R2asw7AMp8gBb8GNr5V
NodSTgJKbXKosKdLwhaf6iK6Nm6JXbz0ri4busvdntpl2MVkBeekXDKl5tLMeWxS
MwcKvVaYM0V57qX2FWCfg5/nGfGonLVW7gFfaUmqihdgl/jYbGuoQlshSygJhxkC
ga/ZBFRHOoFDgvRUrmUNfz22PVtLgw0SrtnIjwM29iaIXoOcIUTsFQ65CrDcz5KX
1H+CkQuS4CsATMeIqLBk+cqmAEXEtdV/MaYFT5mDnBJot11KOdbTsaFIs86R+4tj
WFPtZlMKsqAdxT76w1EKYwqcQNmMEZFNRgy2xyWTi9DUd/OiFpaNFyklIvZ48zac
zdHiiUUvncDSDfulUEtNMzOjIudcd+GcQWJfUuhAOOrZ4hgxO7tQ2GoQl128xVaH
/JUI0JVxTFEihb4k3JZMq4fGmENLv5kahcAwuN30AGz44ZhA23oFtk3FMNusT0wu
YPtW0D+IAdMw/uZFamnHUbTYVNE9R2zUwcpNM4T2VPPnwAzkUHK2I90KeiTOhoDp
wITcEtEhvj7FFvE4AQRuZk6gwl0SwGO92pcT9lemEHYT/jdC+Vo9luKKJpwirHhQ
u+aBOu6AYumVaTUt+q+Tn1KCduw7eM80/fBVdtqlzBIVwxg5cJkwFSDLJoxCOM+u
B5GLwIg20TpW1WKXQJOEYZNLFyxPjXhZfVZnudvmZxUagqf5L4f1ZYOepqe+VdMF
MWaIiOJme/ayc0gFwcALEgtQJNqdJS/v54hAUPeZBWkyO0fn1NlhcustLooRPfT6
ICp/Cx/yZ73EGX2ZVhv5oONLmtdOlCh3IahU2g2VSmvS0LYwWDgKSC56VdejM6V5
FC0OWWmXSNSVgE6MtVehpUG8gqSfN4wa1GbDiaQC++yfIDXH3gAXSrL+tWQrJD4m
XTsppiQs810V39QwpbV+/G2iSgiN+4RI9grkzjlCZIct3TCmUu13APVpgnNb73eH
klMN0JceAQve7EHtMaeLoz5S8WcuazYkWaEfg+UctzUK7aeOYs6GGQOSnGfU5W7Y
3Nnr1r6hYOkvFiF6w/iyZJSa9P72JPkMNk+okcVCE1X84qRcRnIaxymatTCx72+n
WgjOPGgEYTwYsNA36YSy7YGIX6OKpUsgy8p/xCjarXsWH/THhFdxYXFQx1jo2q7N
9prLtD6R7jTcrEEBjErzABbyeu0F1RjplAaCQz7ektXfASvamURpsESekLS1F+5t
7PszAazp9jWTGpwity4krkjFJDqoGLfuKkf9yPAh0kpBbwmJkBelZGjeaYVIC5Qq
dk13OSk7B/y0u4GbCfmC0MA4QDumOHvSVd5cZ62STGgNzCII0iC/+RnIoBLlLPzv
GNUH5fBKAXW8824M4Y2THtgPaN3yig2Vzo5/CHy7/h+m6fSVUBkjl4LMloEQ6tAZ
bY32G/7TCKBzjI3e8h34ddCAV7I51ApnNJceAodtn3p/mzavm7JT7sb/T5bqlQUm
NZxW9Xpn/nlRI506xgHbnsuZ8DesmW0rTC4yI4KvHv+Z8aVb8rHc/oUC8a6e8EEL
nABXzcf8xi85v8ExcD7nRT372gX3I/RmOMtUXIxR2JVtD4h4hOfEFu36C05sQfXl
ysFcespYaaxSW3clZkZhLyreVZzqilYuzXm+QKqe/ybHMHY/Ei3UdUk1XR4kxPz1
XSVRoQ1FshUzreGBXZZlX6vMeFGJa6RsJfDuJ4cnZL8uPCe4i6aDI62phhbpj54f
IQCxlzLE35qW0c92+As06/p0SDZaOxyiKEs5ltI3a+wKvLMc8CHmDdsHu2LkPb1q
WRwVHJIo9kIBnWcZjAaJDv2xCM+9jCGYy4oeCm4aRFHfZcp901Az+JPemoOQORc5
Ff9AHubRb+5j+f9Ywe1VfAXfio3t2gFDEZ+2U+o4+ktKRGkVUPp3fU+xg3/92C8A
ZTYRXytzpU3MTZc9F6sNZW2IEkhuNwEUb2FWOiGnklLDtPCGNn2kBk+Pkj+xxfka
yCKquTXerjSAtOeEfwC+8nqVLz77VPRQ8u6xoJyO7q8GWo30AqhAl1PDWq6Gw7Qa
ZKkdrQBNSNomXoO8rKDgR4tiFTKbkEFgB2T/6/bZyOu+p9iEpuIkUHAJEO0hidqw
hkQGB2EIRGAUNNWRxEakAgD9QRHJXGOQF0IAL/8tbY1rk47Kp23lPw1ELojAysqi
Hmh2sRvUjZm9aflN+oiKU+FmxnVov9Tu0y1RlAsgrlt/j20uoizYpPAmC5MAGz8M
yuS6MS1sUttOpIq6AaMkB26Nd+WaJT/mFBqv3MHCidu7n3+DPizAnhijLHqbpaSX
qdGZYZaxRBPfCtjBxHwnA7dk4X8CaxXNccR9hqJ47aLR8KuzXK78D7v6aMWFdr12
JzlJuDutWonccE5CKSHtRB7NUOAHD4pfr12JQOB0Jq0e7Sovw3Ov5fRuHCeykdKQ
TZ+ojDs3+i2o82/i2O+LwYFWRV8yJ8IH3rx4PoCKyHV2zJ2ZA1cmyre9qfc+GZUb
lGjhvD7xQOiYLHENnmLhovDDbIpfw4fyeQmdOqF9lw9XSVEO2mAanga1bVU/RjA3
TLfPVQZrl1+vkoqkgXDS/iGjT5uYzMktAQGcrgob6dyaHv/UObMmnZSl/NpTTRfd
sGu6TQ68PgS6vVCW1ae7EnSALM2fYwURrIi7lk2YKhcQUHoJqJFFy5dUMM2aJhd+
0yuyGDB7cQno/BC+5fCEK/xGLJV+du2X16OO394vYPOA2l3Qv05WYaTro+odmIGX
hrAVpHFR1/K4R44MqKjfOQIY+HyyMbpEdRB/ZYLL1Gdca3ZUl15RDpp63W+QM8p/
c5HDQ05HzoVJ/O+yktGMwPfTG5sKDjtypgdOkJilwl68ybGQ77PQH4WtUadFp+lP
O067rAYR0hC1KmfagAo9xAQf/Fzd0A1jV666y4KovZLrpiOA0LnSL1DAqQxkGh31
sEzHu0lf9RARGMlMmD5uMeuSDVPAe1xk/4mVLiCwpBKKVf1+D28tdklaOD6JXSUE
Zej4yx3MKUxLI/7enEMKTpd9TU33oHIb4cCqBF3E5461Yq5xdM6HSCq5oCFgSRVN
dg+Kd/aj6CByPzvNnA69qZIqeC0O7IunZZk6K4BmHGLFyQ1HrHFunUuBFjV7bra6
Q2qkwxdXKMA0f0z/6PbIJX+96xiuwHmB8rwi0SQDk0daH4slNST5EWGjcEn4ypEj
aTIADUBMlcJ2tniGewubhgn6TbMAsw+8+hKeveyPZcZ4QD2wn4E4lRiz1anPSqXO
zjrcMD19LE9ar0dlGZ7vH6GA+1ROdQpJD1pGjnqwapglX+BN/HdhfD2hLcYgpyhZ
pDxO+WA1rX8E+Rks55oX3+/yaay+Z8LAjUau5HwZzcBpI5zmxHyQFeOeuLOslFcz
yzG9rFQHn4x2W0fVIV1Y6+Sm9ttDF3NM8LXFZLJIC0Cg/z5S83p/P3okjLUENlGZ
YV6zFZE1JqyxOmfdgYINMYARZs5pfJ71Zq34/U46lPN+VOrNQFqbFo8z8uZIYB1l
OVtaDtRkEs2bgi1GrA1vZ5ZHGZbVQrRo9kdGnrExHl3luBSw2g3gRZLFWi3wDHhB
nzwXeUdIgHXBW4aLXjPsCcwEAtXpq8UaczjSk7doyc6U7QOG/ZGZ9fZmJXq8d8pP
U8R5bvOTrLmqEu5Sqv1tli1L428uBHFhPpqRmDqUE+/rKkvsuaIArI9ts/L+WfpR
pzlPXQKLWEhVzwWl7julK791v5Upw8RNamW4fKgZsUJW9sL2NAVKwkdKVepdcDdH
M0+ZCU+bpF9M59okcMVxaUefdzeJ5MSBE6wB3KuecIe9+mTPoAsTgBBO/E6/pM/o
4eOilAy/rRXoytTKm/ccpAP/A87DbKLp8bX1LbxQp5EfKVa3+duyBMuQOwPoihvX
y0Ad03hEohl5hslbo96+iN8pyo0fbhRC+0JDFDcg6D8R9hdiBUzCForompYPITYs
BQ4IiaktOyrLtYqFlvmSWhBk8bGOwRjNE+AhyGK8qtIWTM8Xk6niU4tHPYEYbaz0
FbvUCKd3WV36c+qz5hcfSpPq5E/NMwQcbKAoHkcqbZOo7AKzn3vs/jNeix3wEDuD
IUFGHu/VOKUj/EUJJUYxKDmNzVfRIvfRjwhB6Z7I71PYRNJOs3qQj8Yk0qcCdiF6
F9AURUEAnacP9gvtpymWvP8g6qEAPSwEHhxv4V9axkjIZwURauubIuquTrNLrYOv
Bttv/egP2KEu5MmvLND12xJodLXtdOzRjn9Ap/zD0Wp9ZOARQIVOnRKZJfotZVaO
HryM1FQtl8W/xH23/FVnDozFS1lCsMEuH2o+SO2gMxIWGbKjGnD3ULWOIHiNwsUQ
AJH+v20f30eo4MLd2PbM1NGzD36gD15f8wQ8FiPDZ1d13YW48+adSQ+pDeoEKjck
Ut1ROp1ZtEMQ0hqpSnPfN0Cb37N7V+DV8F84pjG9rseuE7EKY+Gzidg8V15fwS0D
9DPOiPbVDzp7SNl6aWMnZ07lNdUepDcFNyig5ZocuJS2EZ3+ovgH5OVx0DiJvd9/
nJ28/3p5CFUOJoMXrMUA9rwfHgCitgAaXjCEdTHTtoKWTVnHQSCHvRnPudncg7Kh
w5pOUCw5s8h1wnZ+Telrc7UNXQGf2SJuoSGo9hNB1HfNMcx7g/fKy7bQHLdb/i5d
FrtjnyuBLEBm18b4V/DA99XfFJf82A5/R4zzO3r7OpabtXDkmDDxK02q9ad6Qnxd
FqCd/fTqtszg2bQzfpx7LF9nXJE0m1GJ7B80wsQfl1ixe7LJz4ZZSa1WyClNko/N
00j/4JIbLVMLEZoW4IWgD28yZdlEXnvVa5+JfYM9BDS1x2eL7pzrGOoxcNe9dTsX
/78rS7QRJDN0kmCCrAyQNAGIC+n1U69Ewbr5T46ukvSwyKN/sgCm0bhcTxEZyZ/g
TuY58FxMlmCrg4Mz9DQ8FqQv7q5DJbqOpjkWPtCqOCcrq+N9Pdql8yJp2FYIwoTC
l5K61Td9WNUevIju2br00ZYpFPVAlF4E1GD9FtfJjQdOyc5Mj6J86AUZBTmILLVW
D4bLkzMIHrXFvNwJpd3Oap92jqiJS1ASdB8OJCLbHyogYlB1M2Wsw7LmcnaXTe+0
cax7pCcjkovgIxQINiBbEU68MWz5E80EiNu62Yi1YMIqvb+Hw3k6NZGF61KfoisP
Wztm0MUq5S1CJNRnwjnC2WKFzn1AwK+Ce7qAKu31wGp/JuQab3aHygz+hAvVJ3c0
w1e+ViCSgs8ceZOsK260rBebDRcIPvmvTIJuKBlf492B6Q5ezmLp1M8pXNdieYPn
rLFohnQDI5Fp2kfAM9D/bvW6NeYKGo5xVklTnISL6XFy3b7xLbQ8MDOWlK0WWQvV
0RkhOJoXoclXd0ka2YifHZmEYeW6XP03eZ+nR9WbSJCgjPaLBqHxyFG+e9KITsHL
nFirhqsK+Fkha50LnBFi4y3LP+x8pB/P4pjkZ3KkHYMK70SINsyTG6H4HJSkXdIa
MY0LVKYfrTVXYCNOPBHV3R6wm9UHRSb95GejFvAQcYeUGy9EzoE9WvW3OrFbFB9j
HH4lUoFS6IifgfRbTBdQpcGJqVN15wLfrGyQUWA4EER1GVAI5ehsxrptkl+mivN1
Dvg1Ldb2F6/O/8X9JZ5Wwt4gehoAm1dMakhNnPqU+TL7TBlefNxYNy4jctckFlQW
INguRREhyjI0piSHmh3YwTogZoX+gzqnF26s+yVTf27gF/9La8koiisCZK/aKeuh
GYHYWT49cCSNr+otjyJFF3LnK/Jt/9GDa2TNdyruFsXSlZzZdF5C9NwItQup/MkN
NQaYFH+BTHH/dyLKWwu09+tiEgr9o+uNMvGq2v9dyB+fML0Z+xOYGyZtWmoF2z81
4HLrWl7XHPh7IKo10BG1leTyOcQIblYNpBDFuauwWjAD3yisPdi4hZvir12hpb9W
jtDuX+jYfa50R1pSlGrVd1jpATSSlJ/6w4hVMCZ40TbtZ8q3K5yuhrxTnLAZn07B
616Xk8LFjgWHyF3WC7xrIc1BJQs2b4iETpTxVzh5FbUQJEO8f+EkKFkrs2FuA8KP
Of05IHGNX4xDUxI/4INwJiNwbh8eDy42MWN/gh5jLT7PaDWGXvlW4LqMAVP9gAa3
yIyYzj96+k/B6EKAro5hJxGqOEuwES3CqOyVYSbUOiU5SaEYcl2nIHFCrQttbXX+
0d3Sc7rVggy+wBdG/FKuIS/aexNSLvqhDMIFdgrnC083/3t4EWhfth5w/YSW3Xwc
icrtrjf1v7iiipXwIpKHplkU2x4fVkxzAfeTgN67ob+43aqkS5rohMiWM4j/iY4N
ohUCk868MsBIBZr+afhJFyxbuFiHeMxWrIsvLtHXmpdJN+1jmyCjU6f7a5Pk6hSc
r+C3WllbMrWOr9YU6SpbUixdNo5adT6QIRv3fD3KXEEA+gW/7Y7T0Guu64QP17KJ
7UXeSNobJbPJBdIFT/REWh4j6ixLGtrtecN9lCLPPs7tXWn1sYLw4V0eK5hMocDK
67hWdos+qqWq9e+SBql/WojdIptz0FZ9t/wbij9k/jEMtduvkjWyGndMivp+keZo
MdY1S/gX+8KwRwoCUixNFnGTPX1436Xl8vgJYMPP93pl4ESEzBtSL1LvkoRjmsiu
NXzmVj2WvgfiVvNiR2YoRjf/oCUzKSggNaySfxqnDutWLaRtzOZvoWKf1DxUxwV9
ZPImP/2yJ0dOxwMj3zsarpB+0zKYKRyz6Vu6WL79kygb9LATsyyzxP+XdFF/UuAH
cAqwzt/D4C/R4lmSeyKFiEqR0mwfyT4CMD1pduidWFPrpCBSumu6P0vwlYM9mrWA
CfZzvolMNlVVnTohqREJLTVB6MI7cAkNLR9FcuvkP2QHYdaIotaK65bogNFz7EY7
AGhy9P/AxJPcVw20NW/r+JkYTHgU5pjGpnmPKXyjFBuxaab7ndTbj5Gv6rs7WaaW
FtRevRQo1tMs77OjoeQ09qzn/ILIcBY6tt3ypTjJNNzQXhPZDk8yk9lNiVKBMD+t
OUxz057WY6pBJo3zNbtUYPQRJrnc+0iMhcQZCcExegJxQOgc1om6zo+yfoxkSqTM
i/cP4Do2mku02sEhz2Bxr27Q5QG3tUUTtVHKl/n+c93Zgh6JNTx+Zd7pdzKyvdSz
luSy8UiKxxt0zVxBqrx7rW7GTJDP0Zar5yNJ42V9JFEH5ildHlmrLoTaO0TZjTa/
vz2boAeWuiq8B/8s5AKB29O7Sw5jU1d66TP/41oFbUH6/Ln0ge6MB6ocXA1+KaHc
c2vKwTFB1teg1hQemHzarE4rKHN8gFJ3qiypAmw1L6rMbkJo59dViuHGH1W6sKTx
nlwXlMwbdlmbT2AlBRA1GQ==
`pragma protect end_protected
