// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
VQB7uzaa5wIsyBak2JV8o4Ph+Qo4BuJejZ+uQ2QFmQ1Yi1LoacQ+z8WwdNYkBGmLra8eszEgJipr
CRurXGjAuZDq+eiddEhFV6rDVo5DLNPdHwjk60FAveegvuFlBZMfW8Alv7lQo9VxjXiC82Pj2zns
R7rRwSjnKcGKkenmWknI7ehaS0jvZddheFKRUSQdLuLzwM7TrbZkMrXKVOiooeOaNuZwI5Ot/5FH
E91rH2ML5OHR8SaoLDBzk3IzPCJssg9Kn7voNdt8YmUwfa5MdrwMmzGrF9AIBx/qsjEJOHptn6jX
8Mynqzci/kyUob3QT/xL83FN3d3AeyCx7gxlGQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
/z4iUXeYmD14A6L3UAZ4J2nT5EE/fb+uSRDu29MFG/FzYBx9x3T+z1mXp6ZUXfFKh91pznQeqKZV
uI/ytcqgKOJnx1SIBZNcdP2WfgaDpydORPYHdqI4ftwHsKH8GRvwJ5uSkPaXCsKHEzF/9MEIZk7A
oegWwVLGlkfmU/3X6K4y2LzBdaWMrxnhDin4fFWIjMQTv7Ab9OrA0c4KK/l3ovKjwSQgGEN5lvQG
w1wDJxQnZ4oLUsZqjjB8gzAqo4YimxRJUjMUTFE/8V42H8tcwzBjkm0wC2NakIuKi5Ov46A5nvAD
s0aTVqKbDLpqPwOQIklqQCRwZmfnehT/4ipvrEUVohuk0v+/4HLF9ujOL1WxTwFKgPYpksrWvQzB
c1a4Jo8lqSG+mGIF5uG10iPfDsv/6/8+Algn5JB4/ConWwI5JrGV+8Chx4n/FI6Y1R18c+aGyper
s1Uogig35jujnfgUEm5oopDDAh3bzWugXdtu09ykx5NwbArWKs7Q09mACR6MLcOBdAvYDRSP6oMQ
VHwipqboGcg7zat830PrRg+DfZ14NCAsG2DurSrMp+TWE+QFPVgRtih42p5sug16cXh/rDHOFy4N
COuytsetnL/Sre4mhIxIt+2vUxvd9AVPvU4jZXzgw/vdWTg6rXp/8aT2JAPIpUBZaPkxypZfd5Rr
vedxrL+Cg84CsInfcnOD3zolEyAdNIWzg8LmivKXV/8zlKICFp7KJ837Eeg5b2eraMFOsv2GHCUI
JpCKhu3xZ0ZLFjLNwomQrSrDd92vKkEJgjwOpex02mncfpS+IBV39cmgH7rYRnxvfrJL6JVMotht
HQjfdW+XT9GCCUTVOmyNowaHvU1Ha0NBlZDUsWKHoAyo1k6Z6DZOHX1aELdgvU5HtoFOIqF6QiKt
115u6UsCk81bZ+itmDTi8ta1BZKW038z+uxAAqALKb3LFBvhJT/Pu9okp9KMpGgGcvSjSQBOmxfW
Sfaxy5oTILpI5L/8e3VbBmN8mV0AN/KXNV7jbV4Jqu1Jl2alDy1J+aqLZXirrWTqxB1mYIIB9T0B
BKOqVvRzBhwjXfEiHpy6H6Uu0ZkFeUUH2vgI4QO9c5DLrdyDLnmhcZi7vRNJd6kr+inFWfkeUTuS
Ev5p8Cyny+q87oWUDzOcLhygucNfvxJae1owPwwLMIPVIiHz48jwIs+8fIJz5vBStAgwea+Rfhjr
92yBQZMb/lZq1p9DekVySFKM5jLkqFwedfHVbL8WF65wEn0aLeq1t6R4rkA0DCqo6rUrxAkoENCb
E7X5XVw8VjYC3u0c5SUy6rTcMNRP20WEJk/7MLK+luvMt23U0tgTPbAkZryLmCJqxfALRcYdiCq5
64JBVVr2RVX9lAbQRiDIk8V0CaLVvY6y2R/nrR2BjxxMYRpfEpsKwNGw35mKKBjdgvsyo5T9vzB7
w+aAEYbZxhRVmYaeNczRcXpEm3RdwxJW8uDdEJxy4SC7DXgiJdqbg1GEo31EFtjU3T2Y2kfQw+h6
P+luId1OjH8zsDenNptIwGpa4Ll+g0psDY4V0Cl65+o3Pl3Fz/l9sHgvlXMLuUkBhSweM7sqgzei
FGatG7/sN/KgU7VZo8ffCmHV0pwbEFhf41939mQLLFRHR4n9V272inqpFcC7p9uZ8enxWRz4wR1w
kgF4edanBrvPl/6xxGIRB/xFl8pLmxLfeRAVycWYslJusCLnhljbGWISB2tJCcTs8LDvMTpHhE5S
aamxes0gXvjB1URhwMVjmRqCQn2ECEsWSuvO8haU9qgrid3eIQt1P8wjUde7UbeJrk0OPWtPWHBu
PxGCYwHqcpZVYSj3BblJ2H0wOPKhLrMty8YHuSD6wipIaZUqME2u7wjNIOwN3K0HAI3O3aQmjpwH
eIe7TsqVH9NaO+mclfihIJoJofDx4+KFpDrSJsZPZJaedFx0GWNXadYxj9PSmw1V71maJL6WwUFz
OjqgA+GhMrFmX1IPVJJFNJExvp4tQ734jRtZI5wDcL7k9+M0epynKiwMB+wbPbiP9h0wHGXOXoFD
J0IvbLF+2MlIT+KE5LV44LygeYqS4Y6FQHVcPX/aTrNVnp4/BH+7sEIUIPH8aRjCJeG3KQTdTeNx
8w1IUY9r6GwpFomxQVy9/SLTDXjDnnR/WcJXRkXNes0FVTzLld8I4PGR+kuFnK93WQWroH1upDLs
iCLmhiRlL4xRr4X6tnooqMc55Aql4U4XJN7kfyaO9gCVLSH1zxzVYTu+rq9YVhX5TUobDTESG7wb
214zMms9cT7iH6JqCvlNL3G2Zumf2o2RMXkjXhsBCFZprMqlCmWO/kS2rCi6RHsHhJbjMu3s5ku9
u74LcGnfy58oSl639W4OyF/j1XQiYt8F/P8QWRIw0UDN9HI2+BI/GWn9IOEtgH7urK+wCWByfykl
LedkBtQeR4eAWpQmRFxCGt8XVXmAOa29hoFZOw96R4g7oQmsIVWE9XLGJlfriQ1YRmDnyFXabo1x
vpgUl0nNg6i95OI0pTk5Guo1NDDjZWISGKbwMWFUptQemGsdTc/UPetO7yOTJQLvxKuwelKfbqWx
5yeMYxQpDNaJL86QM0IX2xcP89IneUS2YV/LjQ0gU5Od+WWAKPyNOd8XiOLMoXvFT5W0WltcU6SY
cx+2WdD28VL0I3yhz2ryUlKaXowNE9AjiFEzEwICln+DClC7v2Rs0fN1aduY8PjapAzkmxBsUzrQ
g1bZsLE1AR4a2u0fwqeGSCrChbIBxp7dtdORZsFGT8fxf1pHYm0bYeVKO/g11oI9INJjuh04c+GZ
/po1xP338e37ydVuC7mW8iZoXEZ+fhXs8xLSwrpHLnby7vI/CguKCiTCMYD4KSzwfM7jtcH0tsym
RUdQknWPHqFbcKD7/RXsZUcZmUf9APBSodF9es/+2v0476Y0A99Cgp8CdEuUICH1v6bmXNd/7Cr+
dWlq7g2cLSOhCHLOPUkDfMF3js0Iet0o12wvPcHnKREaF/0FG51zk1P+C/1GDFoAGawqH7sxzgHD
VWTV+i5MIzx0jjy0MHwITl6SgJkkqSTdeGtfDQ3NLXcgtDxIJF2zGqh71OHGOI7eDRznP+xnrrfb
lRA4sUmoAGX4CFz0GG6iuu6VoH/aA8XyA+gzCjXSvoQmfv49GGzXPxWQzeo5/VtopDHT6dj5v4+y
A3VFZaDBNmIYBMritJ9vgweDww/5YZxQANPLIKIO0q29aatrue/DtBw96pPtZa2jMhlqyATjQ9NU
bcb5DoKPps1sEQTWD0V+4AI7/aWW4aXlydtruxye0dSMA8JTkMnzcE2FnQsutMFdQOQKVJc/Eylr
kJzU6cI8UYpdyJpIbsaE1Zv0fJy5foyIQLOvD8KBWl0hhIrwFcOafr4AFqa6ldZZMY7msh+EjQF7
vCmEIF+XMJG8COteyc0thYumrX2H/sk0TOEkit+WADeNxvsPdJP1urQ0SJQsvJF351/uGaHWgUgD
HqTMpcW3OY4YTBvIY7eLUikooe4Hd0Syo1mkki5eNV/bd8ArqxwhSIB9dBnuFo/HxbgJTlzoyNN1
ibfD8Y7kzSOtS97OJKlqLupruYzDS5W8zfNXbT/LI/weqeTDBLoPc3CdTO6CsDZebmM5TAHfrO23
g4Xv4Zxebs5HQxPVYrSIauRKJXuPlBh5IVXxYBIOjCbLuJFkkcOZ5rvHAhBm7k0RRlE8tA0Pr900
iCqkutA1qDZFM9K3kxoJR1kyfUVvbVgz43FHWuEhG4OAT94fSkRnKgkWuSzc4JcCiHv2PuA3Yhsz
CtAVScONHvI2qH2TZs3WUXJkROCbNgQY5c9MqtihIxRMPcZLiZR2LCQBCa5ClxXxqrURVzgXcma/
2ljhRy+x8rnDl1H2Q+6o7z4zHLclYloiKTl0iy7EyyKV6Dvbo24fYWTouULDOhM0F2GmE4tbRJKz
kfoiQGYcAf+uERe9UIOdjiYltqTDnZHueUY6cJUb0FuiGVq1xRaxAdM98WFj94hEIpPh4gPFcqcW
4B0WorA6vlde1cVk43Xq8m7XCSZqBQwXwc7fBrD3p2HH4m2I9iX8jcijqxBq/QoHBhvy1KtvUvz2
s4e1AdVL4zt/dumiW5KfkhmcUtRbdJ3/pt2eaCvvMwMN0eifQbBCA33I7CFi4xSa+5kU7YJH2x8R
ecjjzyhwrNt4An7xWSmWd+DwvHmeltNK8kI0538QZReRjzilVL+oMHSIO4jMGfKQc0ElQovU3p8i
KsTIlZPzrerHpeObcNcODvRWReEy4QIYxE+JusvfbWY6PFLQJqlBfYw037QHdRNOq3axXuPNEPME
rjmU9ouRkCUoMfU5V5b1aQt1qNgnXClKIJ9MdorReCvgHpNdfCJ8qfhqoxDsjxQF920VZa9xdXQv
GrpDYy2035eibS25WHzMHlsnRKkeddlXpdT1o6qDRcHbUyFf79G0qYCcjVwePU4yKCUyEtfuJTMM
uv7vNtRvLTCbYf6RTdXgJ72rqdKSrY4ihCGRwGv9QkY2/y30xq58CU2Of3AVcSarWuqK6QG/Mfsh
X4Imo9a7I2JfxMsoelhVKCzRcGCet56Wvsol6Z/i/MxSvNuCL03sVZ0nW8dvZvI+xNM3N9mpzHdH
QLDNcxp2OSR3lLCGrK/djUnMkVE0Pjj69c5HtJeV0vVU8b83j6y1mmXnRZg99eMxwIoDYFpw+2p+
4Qxy4IOK8ef661yhmb+qSGIsreHiZldTehwpvxFpzu0+Q7T1jWEZh6DldTcJbMCfufBp/vyO4LR9
Ohmflg/QwXOS2WJde1RM8btHygkHCrq5YqqSJQGLAfxhM4NrTUPoCuG2EzdoSu9zdhOzqvMmjIWs
ouD0dmbUr3zo2OFiqfEzeJ56HM7ebCmEsBQ6SBq4COXOzmOoU4/BmVlm27rNaL9skbnMT5xLTbg1
FSmqqc2MZZToO+kC6ls57xhsmU2TGlQRcPMl31K/cAjEWF1uW/UmYtxyKXC/CrBLo9TUnejXYVJ+
uWByTOHn1xUsGZYIe7E+MnwvlPvzP1TKdG0G1Ra1ylVPoXFDLGY2a3miE3mk5Jsc3C8AuxR+5Jpk
/OtDu5TFyRvm+Lo0wWpNxy5r/oxPJUbnVwi1ba+SRGym0e/dn5KRxlC7m21RSJIF1U9yahsgLceo
+D7p9B2vM67ihrkhnjW7UGiZsZsxVllVyFGmZMdS5IbIJ8atAjpVaCeOszXslikrK5yX5r4YvvkN
mXKl64I/H1u5DxozoVdv7QuNho6ChCD0nd8CUjq4/4SHOKXa4EkT07WObg76k7QBNhVffavGbMCs
2igAd7XFb1JmmFt/v+jB6KXCl2ry67Q7lsQ54K1UVFXthjPRvaDxm5N5+RzC74TFxnoHCnWQsj42
L4I2rS21pzH50GzGWG+bhjSOtqT/Ri9NDISZAyigYDAs5OOG6sajae18/ro4S7RuN/x+Tt9SaQZc
ehtLRYgcwwQOlxhKwnl1DR07m+AkzlhhapGbBFaa/cJZJGMRRttg4DIqG//I/NjLaVx9Pca1c/S2
MUqDYM/tg+Kh1YzdInAuGaukH4kbObOrY5kHga8b2yaR+EDMVAfwk1nX6gbaSXl6fsfC5SGquEyW
5n4D6EUPMsQsFsYkO4x9E33T0QA+xYuE9LZdDzSqZ9UblJZc1GYta3PgNy6xwLajn96AgXc6+CGv
JkQTtNJK4DRwtsoIevj0boCpkIA7BxVuz6fPaszQOHPGRfEDaISdXZkyRztl9rB1ucvlV2Dbx/Fq
qNnHngrgdgs9fS2/EBwjtXTXTtIAmA8Lk+AGjMwES+B+xp/2iRzgyewMmki3k18jZ2FhIJfvhEit
GqGTSmnXxDwt/+ttMiy6cBujvyC5qcbvlFpGa+rxtPLaw9z/IHcrA+gfgPl6xduDs4icx4eH+47W
nXSyqm/67Xp364VLvqa00Nnz3eL+9bD2h6IsgGPYRzlHDh3CkR76aJcpKLXfAsEXwOPOMr6doCm+
6qrURVmA9j4ON8Z5Pk6fRBak9iDcab51WF+dKheb1LaWoFKe741rfpRyBx8r1LNPZ9Ow9RA/49OO
3dvPt3uCy+xzXLfF3C4IdJZO4D++eGDBRU1//slFeCqB7zhViYG5yvALt4+ZyR5wDbt1ONQmzOqt
nGscu5OfMq0Eq60oeAhsb89fQ92uDH164QloQU2FiecRjMvqbCLJrb4k6wNh6n+zFyZ0W0vhARP7
6sbnwFRQU+gTdpl79163k6edIsKG9UPAtqAzJwue2QnTMbihXMT/bGIpBPNP7j1gizIasqqZ4aWy
8l+l6LIapAgfnh9NJ1tmxyw1MCYAJcvGdRfDjv2qfGZofw/q4LtjVHMeZDYhaIOEmWbnukFAZxW7
UUqcplq4W23CA/Xx23LL2I4HbdgrJ7utLT/xWlilvgzSTjjIVxDFQsiIkc0MzHEzlhmTs4Yo5k1Y
iDP6A9LZ6zbHRXyokVEgKe6KpHQNIE9aFdqFBr5bs6jHSpEFhCXNfVtmPrx0vjQkPJ5hN7cMucOG
GZnNP7Dpnloi83tyaBq1SRxZznWfqCljrzJEqHB+vgl/KkBE4Va2Fk51asXSUdX/lPeZK3U/L1DO
lZfjCALLT/6f77U4zJe502rHEXyZiwmHQapk5mAvxCrBgNKPlq09wUjtYxUe6ErqcZN9WaOyOCad
cLm92kZtZKdyGZhprsUQcImkNJyg5xBsAhCXGk4Vl7nnBEStJgIFjke2R4YHzPAnpq2xcP86d4E5
qyCPHkG5wPND04VwtIku/8d49aQsPJNkQ7pxsdhVPvFDH1kF5of/EN6OEBLbmY5h+xwu1+d6F0M0
Ljtc0GI9SRCVUcYevrdiqQb8DfU6A2xyw47wIrSgNcsVibR8BsUFts/xSrmgMLU+MF6FdnoV+NeI
khtL8UsCKuU0XuqIX381DqGiUcUBxC67IYe0sNVB+6mzFh3OyqYH82D7BZ6JPLHqyYaGsRsl1I8q
DdCl9Pj+NH3p+cYcuQLdOBd/BJbBJXq7sEnaznrUqxDX5VPwh9imkVeI2DnomXgRiohG9fCDwlrN
E/tXIqIucf+0ncTFL20MBvFL0UJbSeK3tjHr0Vkcwu6di8bEhaX6YMOi8hqnY0Ua6j7XoabveUd4
GgprYwZYGoSKGmHDqIziKX9THZZ5cs+DmOvRTWZtHDRI6mLsEizn1IAJCDbpt36Ioc+UBjNzV8cn
+7PZlS03khGcpmICmolMjewKqXRIaIyxarv+jphqoW3Ga+y/uQHcZPp5LenCSZ22MZju7An2G/hN
lDEinEElpNpZLaFvrdplz/iyQAbrvHotS9CzqngHw+L9b6GW6DKBHTJ1TGF5/6zsAaPgseO+Exkf
PQL6MFqd/YgU3Yvnst+DZCaz+iatQksgcDpC+3P3Uxl3NpHg+oGPjCp9L8Eh2/DLBfmIcsIqChtG
lOYSSSW6HYJcwnyWhs+8bSolwugGrCyXfOeRrZEiwClO4+e0m3UWAG4FPGSupVna0M/BRCMgjZ5D
RChUCmlTBhZGQORSbFS0f3dwCgUysUGyMZKgfT3u3z89UoAyyJBXdOhA+h1SsY/BDN+q9FQGf3lU
AZYKjQGVaRdxtLv+g+2Jmy1FPREXgWBbyJUz1B/iRSg3jPdFAR0FInBpUiyEmh9yPSgVEUZ3YS1Z
7Ioy6JZE5sD4hSRTUOzDTRtXWWbL3+zk5U8oRta5wf2p06SoMjPY7ysBoq6gOs4geX/OPPx8AjAP
airqRIF8g8mKcp/FvNABj2WL7n+OQYGX0zgEjdCKK4deO59o4vHpuLWU70OtiNv1vQQ6hWjJUyFf
TUkxYhLbUfW6eCKOz7eJ1zlS1YtBWrFYD9vn/xogTWvuc2bTnjhGuQlJwIovaM44QQPsvEthOD7/
kRQiEdkScJG68yv2e6XP0inOHSagkiz93mUKompD7tTwC+05B/DT0PtU2uoNA7kkeHpVYr8PxaAt
0a0IjZaxdemzci4/ZWGjp7xBROJykWhPkEbTVITVft4mGuKxBRjW2PCjKRqkw+KXPnNqolJJ6MJA
rfxhkHaohpFDdCaIiFB8XhL/TjUsY5VGWq1ynvAbETEAcRbTSXLfirvdvTp+Ynx5tcyuvsvIy4+d
BchBeS2bxR4bwZBJj4rIts/W6gmkrNrxJYlpkbwEMNMShC+qWUg0gJqF7KhwfOZxr1syIwhzS/Db
StfDNnjjGR6SVanoY6iT4OyD7jNDrL6Npzv1HCdhAQu1KL3EwGlQZ3AiR73VT2kyh53anf2iGF+A
cSExvsuD0/No3k69HozlSoQL3tENJkE5/iOeV0GFqgLf7ZVak0XAxXaAHXAn8cCO1ZJEUQkNQdfJ
kzdMJuQA3T/JvODN2qHzzVV3bHinZEG96EVxVHgCgBsshXq5IyneBo1VkeE6x030n/e7hltmytdE
AftNHOSVqhe+tV4YKYhD8Byi5OBmG08DqvQpjEQXd4bzd3Q6FBzIT27kSO3vpCQl9hvik+NdJw74
aoiPVrueFZVRp9xdWJgIbeLnX8uPzBv9gD9DNlGFJU+Xdqh6sCmv9LslRxdeL7VnDYFOVu038ZM1
dGAtAtFmPLO42+OsnrgxRo4ZV/MQ/KtFBDE2xoAjVCsTCSTmUfTtvK7IhwHlTOiZW3E1r4xPUHAR
gDQLHQYQvkhh4gBRGoadNYkqpz9P3QhNtsromqjUjszt7d/kbpjs5HctB6geuWVhhUEiovU+j5wY
ZL7Wprqe6xo5vZKAK2bgy3BZHDZWYnJ7qKjhIt+aS95lMmOHU+LPYP7IFGdBRI0yVByEWGDWwJr8
tm2t09zCpg+3vuvJNMS6EzDZxw2jnpdHg5WQz/1FVYX5lDscnQfyKDlgaLZyaGZ8Y7XFnx7I5Jpb
3Q95n3mQsVmUj7Q0dSDWQjnJufWFMxnnMvxkgWkRtq9J/uiGjuvFxClpABeUI2dh9xhSO3TihE+y
vL/KP2f5TduYWXt0suYR6uP/1Otk2oU0Ukhf6nbDG/jGCBE9Ab1B1vyRjJuOfZp15t/WHaI5XX7p
pNWUf6gczY3/JQoQO7N8vGE/51t1JnGR7LNa1prSDX4sodvA0ztzFn8aB9p/4yyAm5yNuhHqqpZ9
yhBbqXxLVrloC1148x+xv7kyvwzs3ain6FOqaQTaNgikFxEaP7rp9ORaziM8cFt/RprHRHSG+eKn
hmy0+nQeJbJ+GvDojeFyIozedXIRDSkQPGLGM8asaMECm0zlGZms8mvFWQ0Bah8/tVr9PQudx8Hf
8SebS0WygeNnLMFbUz9wzXVcgTRJfm2BU+ZT8ut8rooYL3ZtCjfJiFoCcW3S7oGRBrdXoj4gNWeL
Romi4I4wkiMk1q7rg5XmbtTuznRKfDB8FVLK3z8bSht9WKAzPF4U3ZHZhIXBlAGREGEIs0Cezhy1
+h/MWzqU4m1wO0jD7JuIwhG7LQjsmPghXVnNZ5zN/XbSfIUmgGeIVcFUBdUtoM7+pWWvCeCkyidI
GhytEyjKnGn09RJaURJTSTJZUfacU8FxSYeNKB9q/o+P2Vsw14fF2WwlcrBk+Lac0i/XqdGyFP0J
M0WRm3+TxaCmuWtn0BDHC0iwNnW6EYJum9Fx40KPiZr5x+96w6v/nHVH80h0lWlpKjlvETGmZnG3
nTVw0MfrQAW+151gbH3gWO/mz5gWTn7/cM0dXY2r04s0mjMUxksA6mgBW8QONSke1GhavNMJu77T
qHaT/oAi0Ng5uH7HfPJb0pHR3FEmGuBkMqprfijoLbs2fvqqJqrm1POxsGurIVDwmH/92gMzzZIT
hub16hPSv4zcknNnYuBcFA0mC6CTKFCDPe7ybsLdMvTc1hW8G/E5IlrbP9Zo8a//Tt/PrNcsdye6
q0+QzL3YrAEpQJM4pO63lxr6M71hPudeoScLv8BVEX0PR1Rt529WopkUWuFfEFdM+vE6pUJ5VxZM
7qYPqqDaDA1DsKCcSGRP/zfFyS4gCM67YyS9Xfo+oUU8NiUbwaUYBF678Z82p+xGT7VelMQpv9f5
M2T4KB6ZlYHWgZyK5jzk3/8J7cRNh9DMBfxATIjVu+TAsK50vXhf41YjbxETyxF9pREKcqN2UpMM
b0BH53mwEihEwP0WbsxfgjelFALDR3J60EImnMwgQnFZA+NTyOMI50M2fDyI2r1lkKzyvgQXqLHT
McE1MiLoOct5KBq5DHEsQjH9mFzqUFin5YJ1yG3qm/+zIQhEcclDDON7gd9oSZescIw1Pq2YSw6J
2vLEYXz6ISHhGHpgIhF60+QlI/c/KQITzlaMHGj/OGdvpBHipWKNx0hz3jaN1NIz78de1GU7+x1N
xa/qa3AgI81kyoVAi05G/TuPkIFSgRsAsg15CJ03QirS6woDyqyQ0dQhknqu0h6ysy4+Q3XqxsIc
tE9Rm4HjAs34+bKb7lvO7OeXrnz+waBjWcblPC408psk+YL8kcQWTwWJSXWRnx4azVK1qp7BLtYh
UHjAmIckNWGtfVWsI9ZScWR8AVA0WWuCMozYnjMlX/rNzgCzurgO1UOpIXdy4FtNr8QCm+ZQI90m
i4HQgEkK7a5Vmh085a252PzH8eUXn7EES1N2mHyE8rOrM4zigswClTCFKbh1SxVwgVNGbO7Hs1Lp
6cACWKgDt9Q/e934vD43J4KKxXSohTeSPlSMnIgdN6mwjHzaIO+4L/CpmCP0xz+ZcfcJxCPUVfP0
1pUii6g7KlBrr24VbJqpD60zapzbemxXySPikNZ6Y1KAPUTinlq4kED0B4HqaT4IOLvpt8SWInu4
1OwUR7UOeRUvdBhZFOS1EGSKH3kb4dt8PSKQcsusNEs0TcXYGWsiMOl4NSIhwPc6gsO+q+zU40Ph
PFNlH86l1wWHN3XMbjLl+1a/bCaKjiu0wY94R1+fnBoKImfnrvuUXGLvQ90sEkYodtBEafKOj6OL
4HDm9/s4+u2DFbjWAf3ZX9RR0KMJBUzqrgLs6jhUbX76vTIIQHQVkjLxQev54F7VnoVLX5/PS9Ic
feoVng3EyiUoFVyXbP5X4zxffQA1k0959tKIaJmIli1IXd0MWHb+UBbfOuTNjsy8+zlwg4dT5eT/
+ysARPkvxPjFB20J4MpF+HxeijrWEO4U/8OO4TGU33hgpG6xvxqQZ1vjdl9djxHC8nJl1BOEM8HO
L8JAS3YIX9PkvRT2xBsaWE4tB7kz+qowHeXWPZDksueY5GKyM/8Z1wh96Qzd5D+6ZJLFgxtz2zX3
nD6Shia8JiyH2Cp1+OpOE3qexkg/OmIpW2yBe9/eIe1/WEr5RsZqFGyGVltGLmwGI8wkgilr5WnV
I1NVFBXU5veDf+wrW3+INgI8G5a0ljlaIullPRz83+84kuKkFM+dPE1iz55h+z3+vi80l+guxARS
PQ8Bjdd0Efnn1M29+FUxeATyCBmus62B0eWXNH/L7UJ9iO0ET0x0Z9HL+Fx7rSfbnwG2DPqurWzz
I2goi5xbOzOQc5DpRopPkcO50TUn/+m0usC8M96OC2oeAmR4c5OJ+7F8WwXA+PaOld1zaOQmHTLs
a0Fna5MSEv2AVCLIHLfKISTnXbV2WjKTGkDv4W8onhuTISQf4w7r0Au9JDGODan9eY16q90YwA8c
iQlmko0VpuxSVPGtP73H4l7Px7EXOybHpyTZabL7oA5fZvLf+24dNotsRD0ym7PmWKdF4M6HGLsw
fwvv3wQezme7YqXMDpcu9T07sc2xE1sN2Zs/dA67saSBceASGE6nlqBIUZwp1Wp4VprnOVbLiVj4
fyBEB7Ox6tmzTOpQguPAtzq9XldD241mXWSKQaEvbYw+Skomv0dR3QzsvDH0P9fBj+xfbc46L7sV
sdvxaDPlevnqBPMfEjP8Xv95BNdYkoYuTSVnfZtOE0hh7JyTwQ4VL9SrBOm73wqxTGtwNJzSVSAG
WCJyDOaJPlEpAv9F8cjnOJr2PF2HGU1oMtm49Hv5gWzHbN1rTZMWJ/B1PbeuEfAbPzKsXDj2NgO6
QdbJ30YujF/PTc+7C7sjy16N11zK7vQKMh4IAm4al7cjckAyAgntP/ooTfnI14OtlhbaMmUEDLCd
5g5IX6RnUA9e2Q1AKXEMHtbFxEe4naNdrCCjPV9mAPwoBfCfIAbkWXh2qZU7qHvPNbSjmZSBVeki
AiVzRozkv2D1q1+MEeG5U3Re0c7yN5J/1390JB1ZdSLGfcCmh36frsuVcu377+IFEsfHxWi+J1/Z
Ll7jn3f+c39JwLA41M6FN6d7pQZH9YfUE5wbCMZtAwuOau5t1xww8JqRqx8GvIEMASyzfIrOqzqm
Sf7+JdrEsGZHP/EX0A3a68xhPSyUryGjwYtAQvPJPEyfjw2lBAHDarT1em9UeYKcrNQSbwsHGKad
tf+rwc1D5fOI5piP99pC39wtlVRLgIvUQzwyj4M2CZy3OW4CN0OlgT3qfbkbo07XPC9C5c8QXuWU
qIuUV7XP7tGr0ot1qMLwzReMp2Zf6WjnUk9PloF8sgwXxEMgoBSd8p1OoyFIhN3j2an9gslrPpvL
y6kOjN9fDloZcVRCshkUigNnq609G+hH+Ht1nXQBY2fDJD1jtoGKalHfTYaqG49M/Q6oW4eUQk9m
vxOuM7KHngKDKWrxk7AE5pWsc8bjffIlzO0j0O5uULQtuoC/+t9koO3qmYm9Wni3+S5yiIhskQHu
2YVNxa9c64hqua2UEHUKPG07OWjHcfL8OXnBS/YtrTQw5U23AT/Zwy7HfLfPkR2RkWekcl4l784z
Gd4ZZ38zavVb9Xxy4PjpsbY5olNsvfr1Pug0N+uS3FGutY6aZnVf9gw4++HCEuet0Y2PBVobTWWP
01OeAge6SyHo5ztv9z/lMS6rSUw6cw7NnqhVMzKhbWtgTYMmzxTIg3bo7jofFM7fVLdB0T4acTH9
P9hD2t1KDBqVieR34iIfy4pFxrbpKFvMtm+As3CHu95YCLytCi/zjx9VkyljVdU8Pdfps/V26cW7
+8RfoSv/zUE2fNEhY0E4Ty8L4DCDE9mu9PkX9nJXJ9/52HtUcdO9ZDSYrrIXTkJqsjEf1rPVXqua
toFd4H24g5Pz3kf11Bl2RYVxsrHbnLGDqyuP7DwrH+aCHjncuZFVL92DgxZElIG2DVRlZ8daKD7E
JswjpPv9NGjkiPgBv9qn4LhO+4LwvGdNFkH3HFw4iW2qJrQ92r9rqFodLtnFfTx615eUpIeyOkpW
3zBosDIzD0Rcxu2fYWzC6cSqt9wJhDu1POZggoWi7dkqpkwY7akaUkKwI5nBwTEKerRZJ4Cgbu/V
PtnhwaI/iopAZLAEWRq0a8NAVXtER5NXqyUA5s0J04NqUzS/5TXvKII7UX8pfjjUYmM48Fv1SL7J
g6iegcn+NtjYuhBJDebZ8FIlsglaIs+1/4+J1Hlfi+fdvE460tr74j1EJtLIJHcoZbri69MbgNTU
z+ekFt7b2v35X/CO+dmCLAIJZn4V8odIA/HcEP9JB9vmeuONgQhjyuj0A+uJ+JJ+N0KXgX3Vdy6I
YB63PmCmefTI3AyFo0WNQU9HghX5I6irkbdbHdAJkgAlSdoS40E6T3QI6ZJTUSkJCwCbFfZTN1xZ
v4xj9n3OI6hWbZfxVKFPkNPF0Yp+GtkO6YW1/w23N8HvTm+qX6+sPO3l34pspOryp2EMk6Kkewjq
v3e63TbzxaLatAI98gW9Wth6t7yq/t7GH/kumkngYr2INtO6A9mYtKLMB17sUB6PIWTFvtCsuKvk
Yc73EHaAMZumrL1ox+8/9ls2INwcHiBnBnxwX83IuYhz7anUffDZGSllgrE2XU5wTYij8PTtLCip
VHgcMmdOBXu3Jmci5qkZhNgSFz0ZDV3s4L8aTeBwsDxCCgLTAuVpXCl3VIyeNjgtZGqRDI9g3Jg8
GSZumOru30fPgDKtAoEcpV0VBXmWtTzYZScDpaJdSPkLdqfkOwXym0LlLihk4HGJ9VSV4OE+FljH
ZZKDswJIVk1wLw7+spX1OYXOmJ0nzT13QxeC7zz7Xl3LS3y6g+Prr4ppsr8QuJKPOuiU03yOjX6I
qfnaQcv/6wDMHzZLK9jGFU7tXAV8TeVRx0jAlvfy6bep2WDTfosoUqoAseukLjVgdR5GEH2JYyN2
QLwX9die9aa83mZnhaoYAS75OjzO4K9ESsZFDVv3b8PRmlWLOLKtliT5XHZqVX9IOp4B6SNvVmVD
VQnPOdfdLWiJXg+J366CAnaktvu6mh/PAV/jeVv/MjgViYwZsESAOZJqMFX4/+6bQfNrV1udhcwd
vYW3GcxF8zh/Ul+Az0hxE/hxJNy9OSpbLJjak7jtFjpGBxcHwZ3pL+Dz2Euf5Ccne5PLEmT3Y5i3
/DrXKHPk0rzWhJ3seu0gu3/rTpS52QxaeuLnnZcZR5UjEOT1lstXu+647nFO2LCG8XiT3xeqj445
Hn5iBcTfBqFuc827E5eE+NIuNLzmJXRcwQy9K3DCAzJheW6DnevRNziBVT6CO0Y3kU7MewXUX72y
UJuMYYMTTmKEXq0xZSuzokldSAe8wgKJzsI5ZrYSZSB9AmIW4cByBpvLl28CkOW29s5iyQQe2kfQ
e/h5YF+PnZMtiNmXU/c5FwZCjoXfjvO55r533bb+fTggRZ7zssMjVrh0eeWlEbrE+UVmCtvRPydt
IR4hCejWRbgTaKU4w6lWegbIXtEjoMTeewgO0hpYSH0VgElJfg2pk+qVPnTFL22/C+shtbf9sCxd
1BM8rVCVvNveVddDBk8Va/QpH/wzLjzFN9NeWxlK3reX/wG8VNDxF+ZE+wrEV5Y7TGSkYC0E5V+d
7iOgOfikV9m9sqBidu/kbc8nA5WI96iw0iHtjXhGJsQzzAshS339KkUwoV+FxdUMi+RWelNvdEcQ
zjURUrhRmTCy5rTr0pcJ6soISXf4tZniBnJpjmMSeM4J3QdswPqPdpa1osApg4B59Gg9ARotivr9
WVF6czQGoNm15q81+ckgnrHMID26CD1CTSbKX2W9Cw0o3/QQzOMW0HHxWS0YV02ACPlHE9DGfIAw
Dju9AOL41XGWeDA3Xw6VMnRe3Bifc0wT6muB0+wl29cQ68z/416CEsb6lJ8R5BTtIB43a2gtNS7v
V/iRvhbSs+VJaM86LHKcHWHVRmhqFDE75WYPcGoispma0QqI4tTvPBssOWZM194h8VjkoHX3K7SA
BRItWKRHlGX9Jcwu0YfDwiBiZ4hG2qP/RCDNOKy0J0x6yfNaAsgyN1f6uyR/iMsZd88HiZNljJbJ
equp7BVReC5WpD7norn3/GYyk17f1qAp2ZWXfDDQQorwi9Bm+dN76SRF3RMq43ARVlZ2JkLjlxHb
RO+0y9QdL7U3Eh7KBGWhB9BdcKtRpsDcT39X/c8+tXPnrCldYyZdJyWomQmRFMkUiLuEGZ77j8a2
RQfQiR01KwXw7oM4TRCT8fi1FgEvhW8Mx3HSbuNudeyADZ6QRu0BASEuq0TU/7l6tS/VTIfBEFJe
c5LtIjLq6Hp3xR8tJJx8B9dsZYVnkwzBnVMaRwaAvZrZAmZ6y16G3hYNDqRHvLKuOzocQYcqctY3
pTZ6FhNXXP9SIxmUY1RWPn0Cjr6xD2tKTaUuvZpaLXp3rySjYxdS8uOXYiOKZhiT06B7IP+3Cyju
VSkINud4brS5VPscQ6/pnUrdr1Iv1VVBN3zT/mPXgHZoVNhnVpWNKKLVh/lUHZnAIMeS0C/KvTU9
bhHnzizXuA1wfLsUnKVb8bogX17kHVSl1GQlBZoXr56tQf+Jl25230FMt0GlWdg6WccuUVht5y/o
YHDHC/z+0RHC0JZYYT+9nYVO+/Hn8PJ41RXHAIy9fEFF6rpH0/smj5fCNBKvdYWwu+TEQB3Y00FM
jjM/zsW6G5tnJ58xYxI8WMimfKB2LCBzjC8oW2pmmLLGYXH/vxO76ywkNe8louAf7H6EoG7nZTl7
Xs95uKJ3vKccGcPeqSENZoQGZE9sXQmUF2vYEXhZaDGfFjngHTPi3m/uBrwaoOxZ3uN8D/jS7aD8
gg8U7vIZ5QCvLSwqB9GQhCtuxwYOyhTssMJFOipPrXBQaZnYQqQJfmnlDhhB32cQZEx3wEzYBJt0
+sKclF2FgUsp2Ksx2jg2iRa/qhTMesDKGgDpofHxoDqmWbq1qpW4wZ2YljvRfpwAn7zvIMRJPesw
qbpzp5JAcRVWBZYrPKQWEvyfZn1kl6Rb6tahndGvQv8jLImv9lI3uK0a9RZS3d5E2tmCHsnHtPtQ
8a2IQ5jqi80mD4GjHovyRrg2KSwsgCgLIE/8d0UNqmgkE5Pv6NZF7rVDhZeN1mKvLbq3RwZq8tXn
YQTz1gH5gpweVFPlIbFEp2Mz/o29ySkVv+3qcHH0591DO8NfxtkCP5mUXwlqF1PNkumGR9FoII6J
5EV6YBWcN3OukcXzBxitH6V+RddfUkIHGJdDWoZXLVFGOlg1P6I49Uee1YlkiSj4LfUzMN6mKkbn
lPuV8uy+vPnXKraCoXlkvM2cqc1nNqkDs+R9wcOt8ZkguRSdujnyZRqhapL22GOf+o2UG01Gp1rp
kmE09Z86t+DnC3svu3DmZzPZMW01Yq7xMge58xNUqC6e2pZMndo8S/XKOQyeSYE781KMTUtblpE5
0dMM/lMypdXEe7mLoDC8KmWLur1HQRNT1pPa+YzmIcRYnTCW1S1kpDQW8iTgLDirWf934qvkcdsw
SNhuRQ2o5NhupSetlB/iowp/mwsKFML+EUQAek8WIQbPYeOX3vCMJ/04JNve9v0jMA0u4DQXb15U
e8XPI5AedyrltZoiDpb+BDitkshAVMwVURkXSugYCI+VAlW0DKLiHEKDaUHpCHcJ3Yuc12+blXL/
yU4e+JzkEjUnxIXW/roSys08HYoDf4BvHy8VW3j7+O6JFZF9qhDgyr1dzfPbFgyV0czQBJBcZnxP
i4tf1fktY6UU4k1zCGB8fiiLvhQW/SELE+tRh5EzYsBjCLdFSMvs1TnEe2/00TiZ9piRywG1nrUa
F6AebZZxVy0SPM9ozTWM8jb73kpA58dI5em0hJaA7IJAh7Uti78QwYtSzJ3k7L+KOq/0DemrOqRG
fxikJ7iPAKLwonPMQ67SaMSubwmCGAgjd23EvZe/m6ZEScKHx5phiaH7qFo6p431SNNXOKX6usMo
q6+8NUYPdNeTzgJyaDfPuydHTdv7ng/I9wY2etOq4BHf9nePIq14f3zp841VQhAtZTrn0R/D1xGc
LL8WPMnbTLlwf1kKOuAHtulBY/ls4W7CdRXyAMavyJhRjfVY3h7m7kFQ3weXTTiFlI0VGAMG7o2G
Oj6pors+A7DvAmA9vJyScsb/IRrLRY3TJ5K4+9htcWeFzPU2WiGA6/hF8RqwJKFlWeBKVsv0Slkz
D7YwnCeSwiX01dK8dn6uoG6nIpTbkW1FYT5ghuWlWZ4yrW4et5oTkbvF5pFKu3xYMdosa6FqLK/L
bFJyNenIWuX7oioPo9eBnTN8RxA3W4IKkf1d6XgkFYQX2/d3LaqbJZlJ3G5TleFbWTu64etC4klo
aReHwCCXm00V9epFtuAjYYL0YVMaNM3nqK37PVGmSkOYH3bsJ8b1J/c4fXnRzkvwYXK59o4retd3
ICGCGhC+or0KlrfNFl9io+1wjlVotPxxagQFvSBmPRKDGOnY5NmZoWYGeITR3zCvInfyNsnNDKoT
MGtfbZAIn5O0JzFGtAlNQ+YLCG+qaTen+Hqa6TBUqNuCwr1J8jUWhjrlEs3TYzPddUR1UVDggHbU
YCtJYwnb+MLQh52WSOkEkLsifvsvJjx9rIatEFJyvrUGOKR/QhRRoyrRTl+/r7/CpxXrLCdRW7/K
XBxcL86PZOY+hbOBPfuaCu1tLUsx7Xd5l0T2FHuTVFQTOiai80+yC3DP7wa2AQXGcJ/Es8WpslNK
tlwxLBX4tHXwpBjWfI5WpBab8bYivP20fcC+a6eysddUudYVDhCI9Gyr1thjIay6D24fC/UR7Nz/
JgvJkwyA9DHVxgASCTBnlfKUh/K2T5skjRnn2xI9PcYPwkox58QcI8yev5qbwwyLrEPRLUoxI/0g
0P3aWzkascXkpktp6qEAbGiz1RICYU1ERCJoX2/XvdFvI9yPm8nVdSMtpx2bHw6LwaHs5ju68uKt
tkRq8fnPlRwB7H8qOHL4jOTrnDM8SCD3y9he3nAJi8CmFhkZVU6mZWXdg22DNnHk09mqRT87DHKP
d1hC2Dhx53c5zQojUS8jXluhoxxylgHjAHjWFiv3DX3GPA4bm2R9RCOf/koXx7RC2okF8lQqxP6D
1Eo1/x8qR2JAC/SD3+5ZNHngyvXOUuN+JaCSXqmnjF8BO60cel6YacYKr2rKA9O1hbf0DL4CBlFO
0LEY8hfLtJtxxtl6CoUrnb0KJJAgkuHfsEFW1nqMCUtkYiHvJafACvhB/cgo12zVxVjyk8YwaYjj
ykjMlhYJTThZOYa25lVB+FbIjGKNThYneVaoTspjByaUCcO1D2utxxj/UsAz4MCWQg4vk4/iWj1u
4P9MhsqStNxuR4myRXXHCkKlkdk14tUOJrhlLh3sauQR7i/kXVE0FVHVe6xV+vtO9TJ6dqtx1BM0
NSvNE9qaElg7ydDDkOYFWzFCNomemAMmzo9Kbt/uAQp8Nm37J1p2SCmg6Cgf1IIe5pwcvD8oiVIK
0O1Ok1uVwoPoaGwGBeL7r5htUpkhlGsU/e9zYn0Hi1W/s7hQSRTFwf7yxkO0j7iRP2cdAx5XO/V1
qwwM5Kg7BDwodOTwTzTp9++EYVEgs3k8YeJqs6l5WXlpGhP6WjnRUdmnApjj8jKqNACYSKzxpOK5
0AiOFVvIE1q3MYHKLq8k2ffsTvQMv5sDdh7t+SN2FcUyrcU+NtaeMdsUlS/xOB8o+H3yLMO87Eu7
rl8PufqVBDFHSbx1cHevrab8Mzisb/btlCEWrgLgzpE8Y+ss7j35hztlrXcajP0SQXwXiZF0rpvd
pN+DLq9MwxxtX4085iu1zn9fvX+iRN8Y8K23gD9rwRf569SLporGyMM5EzhRzTqG9+1+xaQcS2jA
9tuisj9xsvzNVbukB2qGqchJ5rH7YbBaJ5tCXVxVmTHmLVhXaI2Ko5a8EXw9OguBawVLv3ctDgWM
fHk/wsH/E3sPuD7q9ZCqEDinE/yM5Mh1ftZImQZGvNG4dJ+jr4oe+f4Yd8fhRuRxl0pq3Zggn3Mz
6mQHmODW9jotJ2QPqkGZFAIXjS0Y4Voc8udW1mf/YOEJe+ghXxy+yvowmE4CPe7bof0e7N7xNXrB
CDFTwSJxkWauXDZyFi4hFPFHS7y/ERZFRleo9E398X0vU+PEXT7lK2OjOvBQoHuUaVpNusyxcNLV
wLPIfmkmjbv7qVjyQVPZqlxJ++Jwgp/hfJ214ifsW7L0NycuduW19BnDrhAgSMAFbMRY27rmaoym
X/OGUtWMOYlQQapEHQ6kJp6y350OMgmV/tC7h6fVdqjeX/jQ8F10bjid0mdiF46cuMd8yNfqymA4
1sr8xdWh7FXATbIL4YG8Y9OeVkPzXNRzrIrw2vURuHcGawAKXef539/Ok0a3sBn2pgcpMS0r7/tv
qUwgsUo/dzqwvyRgg4Z6/swA92esZMZacSpmO8ObtYrUw9fMzbDbvQt1RshFELlQoP9oEnhcPgRK
GPUwclRI0kD1gQ0cmN+ivYVxqqtg3I+56k1HevTQ1+GD6ealHUnAjPWcEAH1maP/AyGjbIsZRHco
m4oPYmoKxZm5T4yZcN57I6uCplXBbem5/d9EXRpohTplyCM2NFdifQS891SV5sJx9aiifTUf7mcI
5ijthziD9cSHuzK01EvQBiOeBCsMCe65LCNYdRfkSfJ6qFmcm6fcO+oRgzNfcQgCJYBds8gAGPtm
8NpFaI+T4TOOqzrvZIG46Kkk8Nko79KuHu7zwJ6UAg8Pod7VR1c/scVZtUTzjnyyaMkY4eqz/1Ed
WFqVjKS5xFv24uXZL0a+2DlfpbYGFhMjicVBlafiVN9XxNFmSqRVxKjgmkTP5n9We5Hdn+Yw0GL/
vo2CZOpxtcOXKOFY6R3Gtf4/1jZsuficCnyXRrle4POmQkXXGgnRU1mVqytgwQE2nv7YvWGIzM83
ZYwqHRdeQoumc11rIen7rPphjmRttN7Z90KhMD6ZlafV6E+Rbwh474qBg4JQRWc8Ed3B6eaM3Cti
vpfaL+2K7evoq8WImxnTlEjf7IuoVIdQ/6rvEp7aRUBFSHIKpnMUVFHQ/xiAoJFsjXQz9hDEfeQq
wQDHWIv7nzatQTRNGZ6dgOkjlJ6OlrYxsMUSnfPq/dXYWiGnT1CE+cSq6jwTMPrB5kH7i0z+49TH
A7eUC9djphXiLD/l2B4hoLMSYm0o9zDhx2CV07PbUGx14d7hFtksS/9CZqtvRdSAjJ3/utt+5Xnc
9IlJPXu0yJ0YZFpckGRodMygXh+J3bvrDf/AzWO7AqT/L/NoHL4SiRawvJnMGlmVDQB2fUIsjVGb
Pkipf4udRAqL2wQj6KQJOdVVPKECDaWmKlEcULhGft2K5Vf9dh7zq95lVGpwwAZne2BMPkKr1NMV
iRq9L6m8JQ2avCZ6DBGQFF9EyIP4aPO6NFIXcdITYuihWV/d5kJtcpcURMrW5ZNNOarRxLVpE8NY
yYcdCmpL91/M65Bvg+dkqGASdT8mKSzc3GpZ2l1Fo2oqpz5QPku0PVIcUzFw+7ordrJa6VliFmJo
uG63rvCEj3EYMMXKoQS6St5ZLh9qLbYM0qMs3mv1enZtcs0bG5+GYqo1cv3sxdcmSYAzzeIGYtYm
2fWAEMGglG4FODaQKhjCdINudX5Tav4d4iAqbCDhiiBso4FK/1p5up0/GrRfVnVYC3sIKsZ6lUGK
CTRsochE1pSNBP05lpppnQK6m1aiCtQ+YFOcQO3YGpqVKe4est6JOZFoEIEZ9UWLB5UUwBsD5DSP
9R/2lCJgxRswXSWxW03t8+FW4y1xwhO3iUKKXztD2A51c03+mYJ27Nv9dimxXzOPhvfqOwPRIE2q
uyNC53HN/E6cpmk4c4IYzY5zlBTgZ25xRZLSXVIBAKu3aVYz9rMzWwt76nN6DPEev9hYn6J92sw0
6AoLn9IRit8F/F1DLLtEJHeMiJ5dg4vlpdQMAdXsK7oa40aZaG5AN4vcwyhD6vAo/ObcMQgBWfC+
x63SGd3mnWJylG6U+c3uV5QOSh49+x5WF6YnQJ5axJxprdfwrvIe9PcIjV4I56JiPRSvGcJoQgfX
nwNoBWX0HMvoOiUs2bD8mYsnm2TeyQX7u7xtSmeu0SNzTiNU0ozL48WffwTGMjneC6yOoWrHD9GY
0xRI1gMTOGSydc648Owb7KJIBMSfwre0iypCNANW/0IZM5qjApDjMor4wCdXb5FGCAk5U1xmjpwQ
uM39519jw4qamgbzhlPv5en884DbYjyrkuDlVhyrF5WN//EkPW+2bIj5SoxZzlLaa6ZtWYLe+8xK
u3RPHteUzNuvYrr8/hc/Lj8e3DyMcmuPqJgtZXmZ3LfEESn7eNo3nnSr/br30fFOH9hhK0hcWJvz
3ubkpipmt8Ro7icU1pGUQTOxq6T6z2DOCPEYKuHJMCY1h4axLCzKIQEVLFSDJYW+HYUCM8AwXJbo
o37pQLKeu83XRJUpNLzC0JpfafurGdH1YYxuiM8X2OnEbSx4LAU0pHximmtuSFpJJ/EE1g79rQPF
fwlOwOlGlwWL7Z/+iylQ70joWo0OctCYmoFJzRVjxNBU41+NmD0f+mmHjOQ9NNA+gruxjZoyJHQ5
Fob4aA2p5/6hmmzSPcD3UoFj7KEcydZ/OOGOWrFZojnrR8NCRPJo5dCviNdxcRoyfzLovqVPVUMj
t92jqifqM+6TNVQxBOfd6YnZcJXrFRHqpcqXjQUnnJLdA2aedH0mC7eIdSE6vQpPD6j90/2CAYWY
Y6IKs1xHuuRlY2vZEqpaUNMtjny9GxJaJ7MSnvae2Tc/R4gyzjfFgPWMM7GLJ3pc+sA4pFiuNwuj
ZpnbX3G67T/MMQxpjyaiyF7G8k55JYuPCfC6+n86FgqjpedplcE3DldTikJ3td6bc3jhDhqQlFJT
mw+n1V9k3WHw+HrEqO+rPDpbwNhKVJJTgmy/TG3kOuB4S7ITsLlZCdcufgGUK4YsSC1fEHlFnADt
Sjbb1YzLLDrrWJHw7RcdZ/kSOM9mYlb2YCGtAIe4cpZkDzVqruGG90kYNyjU1ZAESKmbyfY1M2i8
VGUrpNW5QU/bMFfW24IvLqBq3oI9QbSmck1LvtfCIzkRTcHzArMo0kXu1fUj+14G0WPfC4Abm+4s
BWrgpd9r8JVL9c82Rs9TmwWFIfqF6tiMP4Aj6TlFdEpcOqYQ69vbNkZpYK18hB3sHj8ZN8LyAhu9
GRTfYDuDKukZgWyonZCPJMtehOl/6hgoNcZ6I2A7PgzhqESm1mb0WAldEdgveFgNcLXwbuzs2ct/
kT5JoszTeLyEzC8GAjswJSdL8TiUi7hgeQqPaKQlWPb48O/yH2Xaw4tKXeiR8PyTNyoO0vcWI0SN
STmG6/A/Yr+XWknAl4V5cFByteEiDsP/tkcw03STWxAnMup/7KSajHLoECjkYzEY9u97w4QsdzeE
Z2K/vcCOrTc8dyyxQtkJN2j+JvwysQ2xbH6ZuRhqoW12DAq+YXUR3XsmuWxetlwBj42hF0OCXZfN
2EMt+Gk91HmrJD8NV8fZxKhjRptOGswNaYQZD2I8eiwGHcd+pMaavEN/AOUYdZkLkSTEvFQsRCdK
ekNL3KOFd66LDDn1Li7rfRgapp7sirmvlZ6on+zrvuDLHYw5YzEEeOjWM6b2egfE4yhhLlktw5MZ
/3/81DSUYp9SIUyNmuv5l83WerZxWCS4BKgtKHvYXzmkR1DR44CniVdmyGbDvn30RDvooBBSuabJ
5fgb7ThBCVaO3OhLdo75Rgp7jDn9ZNc0wBs36CQhgWJbSJndX7UlGJJ6eaLpNO+e3JaGGw0GeCTu
WGbltr2KSYzhyTF27NjrFbvNefq/fr6dn9/kntWejflK9Lh6LbCBeU0r5iJGKfb85CjQNP3ErIdT
tz0qk1TCr4VMwMgRZaknPLK83dEDYIUQwmjZvtLa+jctFA8YIT7pbFf7xFQiPfToycQO3rBuhv4N
bcC7RJrGWTgHlalQSGGp8MFrUaxSKzpWKq+eBtuFHWIhYygJ0V/x04Xn50KqOeqYVANWRnhsrmwd
wprgZ87k3RS4HXDKaGM5QAGt/eo1BYa7sFqzos1rtrpHYtxbpMen1aEXZ69atv6672rWc3EH2JJR
bc7GGNivw0kkUpKQbWz9h9NZ0pHUAMtAxETa6wiBNyptzNOUBYDw7nUTjfa4947WAZLsEeXcolxO
dSK9bk9M7kPx7/s5/4mLRJSO8K3OG5q3qMqFMLLcmvPls+16z8nbZwUm1Lh5iZh8UkicREJ8/Dxj
FQH6bYuI+rqP/owtcO3Yw7YG6f0YIUFLwf/CIhFcZmRpn81CvoL7xrJ1GxeUMZDAZm+YB53xRlRq
iAElcxvKl2tFiBCbe1I9OL4rp2iHHQEv36doNV/ewOW/YvL17zIiCLRZWUGDHAj3zAFZsatQSjuA
JFPjqxAq8t6BBZjLTxrxMAa/3DpIYujZiPJvvGZIFl+IsLHNyRx6rWhj74FZMqfnSaNKxcd9QogG
weNni/cswaMvVw0oIENrsEyf6vxFWQxy5koq9rPLdBOzbtGEJDpEnfd2+uhoL4EjBocO3frl8BXq
XMkiyvO5Q3pj6K+/3zf00xHHJBWn8yAW7nZGcCT7Aaadwn0bCldfQhW89pOFOcegBednfCm1Y/+S
+Spq9uJdAS+0SE5Jilir3Frqq8ekt9AAAxLrlA0qYkrsCquTPGvJMxinhmBK9Ua0Ndyen9RDXsiC
B3gy7l6byX9t8P/HZZHjgTTB9iSUhp6VTdogWQjGCRcWuGFyulSButS9mxJ742r0AdGD9QfI7sCf
ymH+04WteG7yVktqyGAK+FhNeu3e95YF16msV1uY1VvQx0U2yhq/R7eCDto+M1MJ0u4wofJaWbPy
eLezTCZV1TN8KIfEIunjP3e4XGL5pv8kPjIk0AKSoX9oeY06tdBgEEIGwABNaWMfyd9nqygRyB8l
bNCr/D3HJjkvqHthVLlTkxzGyhJfYLHoIqNMTR7P3iHsiOVoNvwWTdyjILexyIkToXYuZM6ayD2w
qLeRXDGGK/9ihAZYSSx1JSY6OPPaEuWhFEmSg7b8FgPX2AMN2Yeb45+kbtTAWBCKfQNUJ6jTxL0f
4HVG1yPB65Ml73fXcupGR8TAi2iXZzXvTZ6gGo+IBZh6IDSh3GZaZLFb64J9JjH1isLxxOGg2gRB
cfkKFro7ry1lRii7NFJxNq30CGLxl0vt7GnAFtqqOYYfWBhqy5Ro3N+ejWh59Lm+/wxm+M1boUXo
ZWu9fxeMtpqAVmUWaUDO+403itstCZKAd4tOUMG6hxTWX2AgYlhM9reUvkgbqPmI+jR69Q6Bl02M
liEkgTZ4BCiy7dNUBoT9A1v0eXjTI4Zurk4N2DELHVR8eL3M5YayCfrIjBsMuvO+O+b6Wc98gAaO
i7C7Nflsg7ZR9z++s+O5p5yvQKbtNcPqk95QrRYA5AFqMwWv19+w9jyay3hcggRPc4eD5PD6G06y
PB42k2vbfg949dx7cu935zjS6Ukquhopm68lu0+xnmQCzz/pU/Dg5zHik98xGlZ61REKPCMk4Pz6
KcdNBdo2iMcXacQhD9RGzQgmcaDNnvaUWnKyHXr2mch3nGbCvHJNGCe2CJONJx2jtTvF3b84T34P
3jC6I3ytk9QLzwrOZEoeuxa61cFyYp1MoVgtXtMpaJSrsUSf7105rRCW+vUDHTqZZ046KmgD2JA3
Nt0HTaTqT1hlRcTfwdLhSN7ArGX5kpFqYN4KWGhzvYMnrMffuOmJe4qo3crqt1ByVSXmAU9z527b
OQ6dSkkYS8h3BN9jHYTcTXZ4E7FlIPe1A5XzdmPrX334YXr4+etDL1UtWAJ6FEo3a9wBMOB8yfRo
Q/H3mHXLyOQRvzwNb36LGpo7XitnGotiXjIqQRtTQ/TymW5WSlXTx4cEy0CdT6+jgEcm0t5y0lmR
4mMlIW5cNp2FiioKI4quc5HtZDd+5wAYlbA56bUrU+vUyD0B9xWHbK8w9S+HyRF/zy54mQPpgp6h
v9IOBQG6d5riViEBWXdqggJvsPtUyvlR+uBLtCl6u2ZUXkcCTGFU/WF6O156/KsZBgI4M0+wop/f
xqChSHzCjDyxsKIH+ScgfW9zNZqYNXZdFyuj1Jfi8nJOSJNhd5NbIXe6vKerhyu6YJD4BKYbZMew
ngIrxcfUJ4McKKWFeEQD7mW2rUIlW3kLQt9DZITgYid44gIKdm5WDDps48x8f+RNcp2BUv4LAKeu
yRHr6u8U4J3Y67BrVQWSQq0H0KwrQYGDFe0QZf4x4xGZVvzKmjVljWuF3zbxoSBFkJYL9pBkVK9j
Aocz8Wu+B7niLklEdniWhsLizFeW+bgDhXEif1bjj6s4b/wjVu+MPLf6h2g6Lj03LdE1xQwk558b
K6RezpV4Pt+usBZEELj9xvH5+/lgniKl+eEFYXs+fT46EyQR2KnwztGra3oqI83/zRYzS0gGjl5m
uDBPlYtkG0UGj5nuGTfFmZx4319GPb5LOYKz+KvfClWnh+jo8RfFdzPWkgY34gXCdNm3BNMcq1dd
e4M/xiRre695Ht7Wku7r05921FUb+Od9kBw+Ik9DuRKzRXsWqpSsCrbJtuXqWHup8qMFnZMNXxSS
DebFB1JIKQhrYQdyyzToWz5qBzpy1tkmh01XYyNq8etjhadjrSO3xse0IUJnrzXIUiVew0QFH7S9
GJAGg/5fP08hjwtHpGW16RwgCVZTibKaRx3upc/O9F5hmyxFk4LFUhptWKm53KlwqUDTijb5FAZ6
nyiQw3ymiig2Zv7OP0PbhjY5ka7dKszedUk7t1WZFAYgB1EEsoqM2y72khyoUMcl/QeBKV9AiB8H
a+IKKbpRso/4yetJAw2uLIS4HeqxUIJOOq1VDBGKramImeoQlXL6REaAwOXUavBJ9anW0Z7ubRB5
poGd7zBjKTYr64WHvqht2wp3Sdyd6ySycXHRM3n8mfRxpB/Iv6+lyGN4pF608MBnjMdfPx5jqVk/
BMqFvxvUjfnXpIUNdkD6cmglKozKdqN5xn1s1hM8RK9RMdonuIrptff1JwnSRNKVEZBM2aw9IY7R
TgOzaODyhmbamTF7EfasbszCYHtVHEPrHSihK8cCLXdBM1JBYiTjcEhQyXPj8hVfK6nhZTnEWiFj
EvIEcrwtwyutck6U9GvEjkEJrVtHWzd3KI/bVY/Tn+ZOrcHmhKbTcd8N9pYYOmdjlB0POUxzNtV3
wB7bhZp6GuY7cvqLAtpn6HiFZLMpeeMs/BiydW2DeEKy0h5/+qdYOlwqOMSVtAp+e5IoZjDfry/b
/BN5gmDNNbJ3YHseL2X5y1JhDcAFWO4Cpr35Tzm1fcVDMaPhP529B2OkkYLwLG7x9KF+kNq2ELiz
/iGRBIT+8L/CLUW1zOK9nGveIBp7Sh8v9NLO4Dsaqq5n25tPXFeVFlerwul/kx6yant8U6iNGQOg
ZasSLGFYvunHa2o5Ncz82GBt13aiA+hBTEpznthg8BTDqLVVhxiOTNBFybH10aWwkQfMXO3mebMA
XPUQEX5E5G3vLjDVJcgLTuGxdW29A+3zA1/mls+dYxN9ayYnAXw0dX8XidEpnDJ6NQdYQ/V3YoCp
zoLHwFR6e63idCKAAzUzJl5ILhPGLq76Jc8a/ZtAzNDO7iA06xBbVqL0iK1nMa7k8wNB73BUuNYl
QhgMnEB3PWv+HCIGsd9410apacbk44wC3yqTCGgYzHurh+MsMa8l4tg/QbYB//UlDllRDd9lSETL
ttfI+Bnt5Ri4HJtpM98CfWa6cbTL2dgLJJt0XaE37uAcp0RI3QEzAyU1w0PAUvNE3s02fSzp9N9j
pjNvwUYOtxR7kWs6XyH8eENSvrTTyTm9sIfXKZn31o72Mk00m3Yk3xZeFHcJZlTqfFkAkyBGbV6E
NEiNFkCTtHLo0sDxJXi0686fvjMGNRGPohbHUfrnQs70V35fPuqLCEciovvvMGL+wqJNjgsKsmnt
ICQ6TkJEHe/O878tNxQwM/PdijfMi6OpLNOY06Tz1wZ+9aE8c9Z6I1arTohpvKRvxQ1QTnVZxq4g
HCBq6tDeWwNhfSEOXGFz1LdhThcRG486U0gxKMYxQuoMozDfNTmYX/ovMWEITIRA9WNPL0OrOUuW
NbskUQbBUI65MjiVO8eZqjrZZ559vifCEQbiAJVXlchKEMSpPkkNCc3N8z6OQAwpX156sQIn7LJI
8JyWUJxYueDOZXHfxN1Wn7XwcmPsXzvGgtBqoWJkDSHFaN2R/J8jPjL3kiSswTHXf1cvDNlPcfxG
mHhgkLkfN4ru6fz38Kg+oM7iMG9Jp4Lzc3wQFcAxUpXI5PW45ffUJbYrChCVnMI3WGuW8gzcBgH8
iDiKQvBXhzdwZ1f1qmR4d28LlRN2jMdlA9MQNpdQnZEzQyCFJfxPJJWeVPfg9W3ixx+7mK56RPVE
oYPnv4/n2bssmP3rBhKCIhEdumxEjnqha+b6k5U5ISZ0ylAQ3LfjSnaAkPlMK8O6fYu/vN6BZsxV
WDIzs8oqDks5e5md7rlS+3ww+wMkaTyotAvxBTSewAqj4vL84ZtDiEoxq7lvtr2jUfNm5qrFMzgF
rEDkZ1gDlNpPDF04Lz07p04qhY1l4LZNetIZyv4N+hq8DvpGrYbJIiZyL76o43U5XGuEnOTQCWi/
ErFte1vq23JflGG2VSOFLHuWqSfae5pv6d8jzWFxe3u1Uko1ayOjmLeriacG27DYedENYDkg4Zjb
ziXKqPMyrI4I5ql5OhzTD+wciWCGV6sgaf7rEkMwbe8GB1YSgQKQANps66vn8YLZUmHN6tqunQPi
NbAoyOrRstH/otqbx5mXT5EPSnVdKioy49d0GYzTSyVC2rN6ycvn1aqgK/b9rjLeBmgRlna+OsUD
Ki0aUB5SFoLtERwGipeFo7Ko8V4ikXpgjKJ42ZH3lVqGYBiGHmSYwYwFS1SHchtxwQkVn1QOCVfz
3KCqgN2IiRiFSzVPjgZSn3XvszdAAxWHdxFgbaEZrxbGmNWe9Izo3HOgDIo5cDr6xHzvWZFq3YK8
wcDmT3/n2hIGsQ0AGrViJDDvcLwwZIGuWKpFUS1Z9mbT/19fj2kODSDELDUEtHysC2ie4ClQC3Ic
ckAF/Vt6vzVZ2C+LdIvHCBY9ZvOvqK9b9rV8MsoQ7rT7MSfTc33GUcVOc0jMqfH4Z3dU7AOg+Q3M
OXeXD6V+Qxa9zoV/GrnqDVPTbuQmW7L1IjHg0dh2G3vsScO0Rt4cnel7qjt9GYZCs9mqawnWCmfp
5isG3xpghGSus/VkTYHgeVtKP0cqZl2CbNJkVB7k4sPIP9UhO2fkgxmji4kBkJkhGc6aozbFY670
NSdOTnOU0fjMkI5AT7Fa+hCaiCG4kI1+5uTgZlWVg5xkQeeK+NKX5wkSAiv68msqmy4X9Dt6NrRy
CG03jpJWI4WFhQmjL5aNNQxFbICVKwh8h6oN8jgR3f/alxW8/YdNTjQtqNv54Zz4e8snfTqavnNw
sC+bLccuew8kwBu6ET/YjMTbAwsRSZ2fExfnW7Vqn+smeFaP3yKeor0g6IH3jDVJ77McWarziFhT
PTVEGKD2BOhEC1ms5Qv24WIPDW5EfKh97AH9yB/C5Tt5algSG8kMhBOE7Vr0PBI/tD0u4/V+iMOH
G4oJ1NdQKpGgS5cHtlqEi1WAbnnngzvQJWH7rajwLee29hkw7b8//l2p56GSniYjRxjUiaF4qPZR
93N88dZLAI/IE01Rewh4d/PCZii4B//Wfbe/AVzbpKPCeYiABRHNzkwudrJpuYAqyI/ICqJubZ6T
K/NpUMVsihdvJWtBAWlzZXO84SDIVdW5oHapYhegn1x8su+VetcubTey8xHLE+8vaBRMZgaAHewC
rJOc9LOVyFv/ZgSrtne0MW5vhQkNnyF4yB0ocpJtgedHWO9SM4vyl/9E2o+z/RufTgJ1BWVuPu1U
dB68MM3fooqQC7l9uccw+k0OjOjJAJuiH5b10zhV/HVOtHKy9w5qn0T+jh49ILk7Fa9AZd56jSC3
C5DaZn8B0/2dzeGFNk9Tya0TsPcRcndggjZKA/wHQSX1KwhGKiglY70ZgjYUYChH9rsPcG3y1VuS
rCWMcrZvjAUbAOXlrGeZYEaMcTC9x33h5r6s/soSPFA5mNdsci8AhlueX/hH/GlUhqlQI5QrTM5a
8hOJvqYy+fkdZNs6IiGoPyFar38nr2lixhucQH2VsYoigAKYD8urLvubNr3MJ9MLLIKIgmGGzh0g
uF+ObcISy2mGF3lK75uKLix/zk/8HY3RgdKyEYr8AhtgJBJW/pAvHXRELyiS6Wv38ZThd7zs4jkp
8ILmVUJfoN/Cuwc1vc/kVql0fUP532+i1IpiGK/GqEzSbPEJwDYIvqe8HFRD9fxJpttKKFSwNf6z
6yMmcGvEK7Hcy6H+LnfRBQa0FgO6KM1bxTRTtO8XXNkHI9SvW8yk/E3o4P8nx5vngOA5vT2vUIFv
+CPt24qIx9JXjTAz8b+YyocdYk3bH4PbL3/ovcfi8awshbNHQ4FHZneF/y1KTU23AHmoPZ+BryYn
VFS7aG5XCZFVihw9ftjbS2v9BcGYkau2vRqAE2fGK9BICyoc06wGTg0M7S6JmtwdJHnfWYdF8XpZ
gvIgVntVkpeTvwD+rKcM6gqpJydr9jC76cIL4FMulD+PhGgBA4RAphmf17tJcsZ8dnLgdmxKEPO2
gpaBNhGQDyxFIgNqudhSIwRlkvRCBy3ZVsk3LdtwAO3HoAjJoB+CETWMyCYq0nmY2Js24Ue+8kjO
uYtUVE4u7fS6Zf6wyw7JF4uvL/4GNvzaUHgawi//mbaGzWJVBrL6R41au37+1dN4ohqme3Gnq66l
CVAfmfx5jrMdVARipJCN9T0JbABeiiYVFQlR3Zsu1/yJ+dPg0nSCivj0K8SMODc6Nn+Jf0UbXWYt
FUYM1usTSUtJ5tWviIQPBS7ed2BgD66cLyNblQEd59PWSNkEZGjMNhofeFINAGDW1KArfSsqcnAa
CuImv2EvmipagocCbCxRjnMvjOGMNT0XtA0DbOh1Qg1hK3Z9pN7qvhnoiR5PJuVEyQfUtykYLAPT
ZF2q8tVNuKzpvJoI/0VMUOB04FoZj0nPQ1HTKQ6bfLG/OlP/kD/Rrw974pWfOOPkvo2ooJxB7oC+
6S9QlO3YF9eyx31djo6LfzKSyt2MtSO35O0OGNhxbePEFG6byf7r4YIrG/4PKqsktlapV+V/MxXV
Sf/6QXtxQmx3I/rbUw5LTieQhCvsZyNNr2A8YUnrPfvxBIqB3KfozLIe1X3V5MbUmYbmMlDtkY1C
bshkKDiRZWCpRwRh024tfBI2HzRCPgFeF4mgRrZ7phwKopDRDBEKawWEFfvTCV2fkK2hf4K+r4bo
VTYnLpu4vLFS9y+5F/U06ONp91WIiJJrlwe2hOULz5unZICLNOK1HCQUuMOzaUaFugdwMmvIEeWq
Gz5PgbPQUO5gzEWAcwWkVd119CgbiRIRed2URqnDiUExxRQhaSamReQe8S8BgdQUn3wSdNRCblO3
pnDUFMDnhqdn/MzpYTwSIr46teoCxfIS8Iu9Ihwv1+xyzmpj+6G2jxh044ADe6AwroZDckjn2Pgc
70PNUxD3sJcfC/aP+Iu0+EqJiD89aTT3zjsJmHnz71PJ50gq5H9s7C4CETjPaGiu+vbVnZxyWFd1
Zf4wHHp5X8GTGY4I0/R3yWYjlUcqaOXlQLe2PwHqaOBkDRKb1zVLk+9iZXIw17I1Ka0eLWDMEybw
ixssbdgLwQumr1pQkvu9m6ENt9gjuyEo3GDMviYAntUEIaGWPNgOEangVB17PkQqXj3TeIEk26Dg
Xmx/f7H1zhGTDZ3x/Bp7Uj3x+8FLG7ClWBhjzJvWcwLdTy9jA8Pejs7vyg0tftPVJR/OHoAsj/Mr
KjUxH33i5ZH3WFeaHC/40rmje7k5mPDs304yrXLoDBeu/GaAK5dacqhu3uH2X8K01gtRvxUKxFcZ
HBQUFUR7UTXe6ZjD6al7SZID0UmmNVtI4KuQmcWtAMKHxJWNq+ZsPO0ZfzF0VuewGaD/jXUwGuMq
61QeUP2kqEDVYtrt+uwYr5YNDO3qY2y211J1V+yuY+Oau6Oz2ZfbG4JCYHb5ARmzS+1J8erxIxZ5
thjS6hw1H5WydiRxBv4nTv8m1E+4w24ohQ2jFn54j3+AKbjp+fgZ40Kh/8tNVlJNAMt/uUH7aTvt
XGcmamnKjB4W1ec43LeB5nnquvdDMfNOEpMkNymlvdpw10y71XxKmfpZxV37Hsbg/fMam/gqq8SK
0331Pd9zkxuMN5oJ8OuK5H+fzUMckKvBbzS/c6gRaTJadAT0NQx2q6C1+O0ah9WV6HkHBWG7kHuu
8ZfF6zjA/0J8irTtNZz+QKHKVegdoPmpAVxfZA7WDjzTAPckjfbg93hPM5FloSCU72fI2a4F9yfA
+UXRcYZU59WNpYgk0Ky5hk504MJD0aNtjJ5JLCGKlqvMJ73G+IUL4tNSOHZmApNdJX894hKaE6+f
QKAbd4heQDcSP41yCiOacyDsP9mRHkS5iwOiqIfRnZugzhb3yBBrCHo9yBeoAyD+hfDiXHvJqpq1
6HuC3fUMOJgpmrngTNyCdF7Ckcv434FcQdODNkGOz2LfvbB/b/a7oolNmoiksExYQGwl6VzR4Skm
lJ9EL6j0hFlFL9kGHc/lM4UxuYTCh7/OYn4Iyn/8IXqRZfNDt5tk8rvzMge/45qE6GR7g3EpvLik
5NeyAgcEDbJpau22aA5XNnAnJy5cIRars8NOzwjsTdMTPvy1d1f3BCWzkW1BA5/FGtvLcz29S4rw
Qf/6mZaeMrTA4hya69IvlBXkVtN4b7HUtzkhy5TDjS0IhY9quj6ZlF/a/Zdtl4nVYSXBDX/2eCxB
a1LYenWJi3eTr0EGnDibCAU6ru8OHKpeh0DaLlPut1s7+w5uFLWG2IYW6e3BjxseA2XlyRjl0Kmm
I7Z94HdYuhAHE+9VMP8G9awnUju4W3PE1wDc3WWgsy+iP47kqaz97xUA68iA4YBQS2jlcfNyu7oJ
lAbblfItsyvdgwDAFQOwG6Tr8/Z4lwFV2A+YetXy2935/InZE5rjjup3GmrGTnmVZYmdoYer4NM6
MrXMNiKNOBiYFB1vDbafTFC5qHxfBHcWpV+d0h4OCYVVGqQkkJuAwh9MRjtTkQiM+tDYj2MqgVOM
cMmM+hxH5TAKEImg2VJlOS+V5d14ZC6Wk/JW+nsKDFfMoztK5UAyTAxCExOFZ+7BgKejP7OwpA+p
SKFybyVc/rQO+Lag89cahp+GY+OdDD4ypChO3qy4OyY4hIFIqA+l5d+tk//YGdr0JTc1BpfB7RCM
DP+8HdloGezPNUqX3ywA1pVTQV6LNsau3JmKbj4vK/FOSytIgd3xcRPSgAMQPMjzLXwkWlucfei1
5WNVybE6G4rVNVdU3CUwYl0Fn05NZ8DkqVazvtsyJ5c6uZ5S6noRkCCppIEzFdi4xzaPmugLMHdQ
MacC86dY/AOKZg1WLQeKoHu6MO8Svho3iXza/VnpI/cgiwYJ2n0au/EbzSK16rC1JRyNgSqdtxmp
uGxojqiaB1qmUeypEwM57MBzdxACm6+AO9c1h6xGEEaFWWid/ZndruhiZQP818egL745isWPLqix
M8qnEaL+OkN7aiXjIRfUdFLqfsRRm19Mbs8CiphXgoO9REl3MnScuVIAWyYe7NjcHX4kTwQg9uGE
opUnaoeedLsqDY2Eq/vCsJQLMfhyDDLWoW02Fy2g1fd+tG4AcTehxHk0V8nD5mtr9PppZkhlBUr+
TuWm9V8JistUGiKs6psV5Tr0Gc/GDyP0X0jgZFJB4DRktqcgBuGicGLGBZT5j+93UZenK+aCXj2g
zhMmfwSs3yQcQ8inMkG7649PheeqmF8zUFdBoCqzWHMns/iGcRYJgnF781Ku5xGxYopF7/leUrFT
obmt+hjggQtRiR7vkjEkyMO8EFjHsVIgrZMnNDUOWrnmwfTo3pQ2WxRoKTUzuHzICz619iRhgXKA
puqX3MNqmIykQlkUtQLVvzkZ+oLa8roe2ov7vjpRsuVDnoCD7j6tY2ku/90003cOEhAUqGVZ6qDs
+zaOJyhMuumyFRoRhGZnZ+YwJBpe+n00UxworX8VzugJ4k5eyFRqgONvxGTbgnR/vtN/gnnGxCO8
jtOjstfm/wLiFK5B2d7jdCPGW1n3SI6fEaFoSOA25V/Md3V5eUBv8eo9Z5RJDxQ+wFYvJP/yKAUj
3QE23lAu58ttFyChv1ooqHkqU2jkc97ndyO4xZvFWMgS0KTB1hotzUy6JXelYmN71JYUYDT9ghlU
yAPmXldP0F2qVtLo965Ra3TK8BmOM0wReME93uM61KmTERBPmmpGsb+aSvWYZgKlHnt+6ZM4Z9Zk
Rx5nN+zL08eZZgPaYUi9MP07o8Ww5OXeN15hqWVX2fM/dHi2xXCS2bzKroRGpoysAn2TEhWc1BMS
e6a8W8kkHncSy57B5V1DFY08421H4Fj3sdmEx8JeM0ZGAAJR5WQhABLktGBa58R6d5TJsRGcwMgN
eNNqgP9tQeIiBTrGEzT3RXmqJhAh/oXdu6Dzv5eROjE9R5iIi/G6EeUrsMl7D/uazlhF4mBmFVwr
UAisQ/9/arXtGG1e2RqZhxKwbp4PQGWOTlFOLpU+dWdgaTbf3GbKfcl6g08d7bP4UNFDn4K8wizb
bgpiGJ6t/+FO70awu7F4H8eD13Fjj5DsN/DxtVGrJNaHLBd3Uin05CETliqEBVlbj20p5oDiS9Iw
vYLDBNSoS8drPV4AbXiIw2eGUeooP6usvkKByS2YRSYMjFVpNFV6JvFTsSU4yQf1t8As3d8rYYM2
cIV8GLG40M2FPqe99Pm2AY8qGL4mm5qnySKW/GI6ixaTYgimzO36Uwy0F1FMVUj9Chb/ktrp5qcQ
TmysWI7mMzbLCX2mpYvfhx5xZcFqZFzR9jJWfXzm4HRJUD4et4YYLbLfnAAfCZ1hRcteTCX/zNqA
WNrY0N4xsABHgjKq6spn5ek61t3e1TZQFrN7CagptpJm0K+tP/A2X0Dt+sNHG0/LOum/ZW9hduKO
9y28Ri/J2sVt34WxocJia5UFiidEUKfNrxxKNMQusqiqOGbIS4hNuHuWB+KpgMLVRb7AAiJEWZBR
ClPCeuKS6hofNRQ/RmVfAHERLT82ZN/0TWF744oCdkjnlingi82L8YzajMwOBWwwF3Y1kFKMivbz
UDRdZLJ3YMGKK4OQkikNouK2wGNPOWak9sg71+KQiP3MJTHF3CsxVt6fH+xgvxG6lEhOGAXbQsd4
KYrrStfphwsQhtw+BCtG6lWyAZRzyH9FZr+uzslUqELpcUdWDxIGyl4EDz7JvVnXuKA5sSTYcdfx
fiKX58YX6BXyvwZ3XHkCLNUWn9SYE5GVwbMxhN5U7vZRMUwG2QQ6VVMn2hKKANKKpqZi6w7Dhu3L
EuK6CfeebTIqmUXgY6gwsjqIqBwNeqrVjDI4l0fjvU9DCW3Lk3YQtmBNtU7iMByr+7HfFNUyjKw4
QGBzbzx2Y9fH+dTwoqt6XhZq3/TTy3QRr3/g7XWAv4UyTFko9S2xAHKfqjwz0mtUoOpGd0zU05W8
xaNPwHn8efGZzKQ3w9PJFgZqj10pTtHVa4RD1EB5HDmCRlTIPMPdiEpUablHxJvcO2hpB2Vms3hT
fmyvVFzLdKUaRmjiVNef1c11NL2xPxd9MQImNYFE77PUIPino6yIFsCRaSopWZbn9eO6k14f/d2c
vpaUgvAbCrG7pVMgsejL+4chuowAlPPuqjgCn8c5SZeFu0L8VKiwHWb6Y6hJld4dwXx+vMN80CwH
lwFTfwHSGgxr683JiFfC7Nh7RvsUq9HnC3BOBWd2LYtNgxXjSaE3hJJGd53ShX3XqXtweW5EsJWr
lo7LcwXHD27LfIQGGnTcmvnK/JiF79zyWq931UKme2UvSzRX3ICh4mOyz1vX+6vepHiTNXZsNrry
JhW94bBKm7LJ72lcnrJXM9aD7o1tNuvUTlWJSoLRHTSZk+8hTGufXgfBfIFh0iKB7XNFb5GpNph0
wWHvKOhihufei+GXhCN8s1I3Fx7LUlc1sjXS4t3KK68jTa25s7lCy6LLv4qahK/ys+rdfQwOoWO6
uJEsiSfVXMu/gptfzQdnVE+8ZUsnZkxQgzv79ZBUAPNsOZx5+rZ/+ch8631SaMofQ7Ub2PCs9zhB
2bPM/Gvo6wwtzFIZl3tiUXq/HN6YVFdGu6RKG2irnmbck07s1dAqDCaPUmD7tfwtiJVKp7sxL440
ZMNUbkGjz/WzVKKP/KzHJa9Bxc3AVeOYhyrmgZTxaLVvOWuiMClCy83lhfF79rtRN5j8TNesPEav
ruFXE11DbV3sVB+adoRTEjL2rBnRfOdPj4Uj1BIbJ3mgtns1zmk9zDn17LebFuF2JF6Dw1gDaRYy
Vf07taeSwRFmxcZq+op5N58QWsyVgds66OY2ldSSPMJWw+cZ6coHs6ycwkFuu3qWfNdDbcfCQTPf
DnSl8UYNoK7KjyS9xyKKiOCZ4FW8VIxK2KDS4OIFW+VqVGR4yf7fkAYMJCYffbOJI76wHzKRmehQ
2B1xUoVxZcQ3vRTOsl04yqbzoJyFlAiA344WiBRsdWk8C8AWIozGbkCeaKpeiYCd9nSLOQggNMC1
fC3tjcjyRSBsI0NiKBCMEr5Dh0tZC+hDhAmiESqStSYpuSPz/1pXca860lJBP1s9C0lNxhO7tKbI
kRHX073NSMa/t/tAA6JNsy2xbsEzvQPfO41vkdQZ6yF0iZvkvs/bnzjWnK1nUFAFFlfv9mFCF30f
lThlsepXyUoDHY8l808WIZCsvz3r8gG9AgDa9VYiSP4ye2SyOYQ6NxQQOZDSfIYz5skLrzpS/h/l
RXtPNoyWoG7iQnxp2+M6wUN7uAhaWFpZxtqM++e0Stlc96XJ5OF+6btp5F25qz9W0EU5Ysm3acdy
RZZ0n5Bbfad/xOuLUKLhdNvQx+MkZVkNX+0fs1bGuhWXBOEGZap8WrZsrWI1fJEcG4jmIWaHFVUd
W1j9uVX58jYwlkWFXYlpY1ZPvQ65NLR/+SahNBj5MtWTQEMpTJP4oRT/hUiF5OzMC2hndrZajs/3
mydWWIyV0x4eNh4IBuXGQL1E7spItvsUdXyOgqmSsowPQbqtSa4jt2yVUgV4qOrMff2RutgW0rS0
u82TrNeXTqgEU2tDS5dNbZPAuPLSvkMYcrz2PRLRi+sdXI5ymd8+d4N2RDCO+PUTmVNts4j8NCV2
6UOzKHmiodTgRAIoeRLROuSKdnGyjpGtOuy5sqFRcLXpcgjZaBQ/43WQL5kTeTO7lHFqGzoMIovc
xYRF1X0pvjsfMGdwb90yJxLM1H3IOSAhaf7Os+cDTUvX8ueNrxdoe0UvwlGSrd6REtHtym/4dNV4
Br6hQqki4pi6I74/LRMuNxlwDY2vktRQuP5psvMjoPyxttIWq7WmdLP8FJ14O/hdOL0odrX18UyY
CdLa+ch9FPVbP645Zn/avYnkYytDD7dQq6d208XetgfWKUIq30BjDAr+cMgPhBcePMH9XmLx/P9N
+oeMQs/xXA4dv90TtT0SYBDLslBhlqNa7hkoysw1Apz5/Q7j+SXZMiEGgfjzRAYvhVGj1R3MjDIa
9iVEkNcAQCl1RT+NC8IbX3yWUT6qtgA053meUL6vgn3Eo8ry2XeP4DWmphSIKq/wCUCKj0MSwkam
/3b3bHCX+Qn/kfHY+WFgzpIrOQ6rUplscA5DaP+vkHmqexABETvQz8WevcVzph3lXaXvnUN+E6/Y
W6NKZ+o63dYxWWwlX9DJlbsvza/Y3KhguUwbhR8E1l1H7wi9Rvm5D0kl+GFkK2O95kUHyfYysAEr
mzNd8kh6y9hSF2MqEgSlyi0/UaP7J0mavv10ZMAeS+Sec3MgYtkBrmIg6I1F92JEDn5M1Nj3VM1z
5S3urhMbAOJ7X86mJc7gjt9rGclrjobwCheLhR0076VaJBKXiMSXeWtOjjOV1gt9FJSo3yRcbAca
nVY6eZKDQoTjAAfOj+mf7KEjnEQH2OSHlkHKPZRoVCRI0Yj9Co7SUZwBi314p5a0+lLGjJLzpoEh
THz/HMUikhwP345McLokumq9oPscZqC6fgjXSeO+HQlZlQCcuKHY/UjNRgQQ7zaolgwdrnbChyXc
gi+3J7Q/v/KQrJGkvwt2oECg/YaqdZK+HKHOuDe7zZNEJoHpoqpeLPTkKRiTAhjOwronfX03jorD
ijqwao+mucSaiS4OkLZa37PFRoaHUwOcdq36OpUBUCqsZAvFmrdzA3ZX7bEz6iPfBejeI32R/4be
z3SMqw0uxzGx
`pragma protect end_protected
