// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JruShHsaqd6j4gmeRMwQ+aj9fo8xOcBqLnutulE8f0RfF6/Mw6xL9jW/VLquYE4b
m4RS70j9lBM1yvD+DFYF2JTkn2yFqmusn4Nfqia4udNaPcbTGNeC/DzF/FAA9AAb
aEl1YPa0ZXmqrZLNrCVOiRgg6M+gsiB0gBaG3Ut5xOc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11728)
a1uwf+lj+VzukXYU7m4ZeOV7CwdsndNUln6FYB0pae6AeTTyNCf5S5v4lThSfnZ9
4w89JGIQYO2qrxEXiCUBAM5YvrzkCfycGPxoJ/a9Y6tK+DfesOXyoUXxaQwGo654
aWsVSKt1krzHU5ji7Ec1/XF+yHp6CdH/iP67oFY5qadOSS560+vp3qJcQuYZy3vu
D/gvo1t07q92h4IEVBD5hhPo7/8u6ZYb5w/WxZ1nNqWcUb7PIinfKl3N3mzntqeY
7TTrKEVoKvNTO5pOsAWMoNW3a7efz68HgtUp5o4mZlp7/aX9diRmDQDm6ah52wet
KqY2O0XUlB/TNIo5lCTdkz/THFXbNGJZcvOGT8g+5F4Cugit/iTYR5gpT9MzpBEl
9ZZTmix3ddMQk+X9VIeJltPyUVdIvPKA28lBAtJ1mae70AUfkeYHpg8weDdVE0PR
MYtYIamthYBnNEG4TmszA6AfonqgrvOMdMnukc11BW6yjEhmbLE9d8+dl+npFb0M
2Q8LdAgH6LXRFbEHfuenGnAMqxD2aSPl3ZHOTl+evsZLTBP3/qP2woRohGLq+Pbz
pz9YYS+zaGuSxwJIobJuoCCAlsnIVvR9uN/9xXe6Xl2fZV1pKmvUBnIczMiHb6s4
7buGRSswPhqKWrCh0+OOeKzOwHg0hpWsPUF2SnxWIsArrYJRfXU9MJC02qmH+ScE
oR/VIDVRtXqYo0uGjNAonBwbaRRi02/6kLiZPPNPju7nGwL/ARhx8gIoaWw2w8nP
EHEdroV24+qQEozKxcAgBF/T7dvdp8qrBFtgoFeJ6P4uCXkZ6H3WhLZHmYcH8fwF
bGQ9PN3UXD2UGcSOxR3b7q5ZC3G1Oaox4mvLMxSckpReK/I+kUEs1K46G7/jlcrM
QC+HKnsy5Ev3hZDYUSnIWmBJONfL8kUNxbaQS0TNH1iUZ02pvwa8XueCezBgMpLd
VwWiHXwaUlwSkssrz2chIVIghT/L7efH5nb2uuoU1IoUs1wNF0RdzgsRk5BeyAB8
d33+uHNJktReO+O4ExSsbXjgZc8/YyF0zpgiTJkaUFINS3I8qxtgrZADIkXQroIL
oGU+y2TeS4+Uzn4NZA675Zfp2Pyf+lvpb2ueFsaTAqEMw2mGyj5reS+2guT+r3yV
v0+SkkkPYCOBtR9Bl4A2cIc/OgKqhNp4dSp+l+8J92GNUuWy+uu1eDpsUi5E2EQ7
+NHPaN5iwynE/tB56sEMpjCFQriC6jbOkxIHmnA4qkQsjXK8dp/B3zEqevYOKay1
GMdbCx02beSZGtMIChbm9H+AY62hQYQEc7O3qGOpBqlHh9shtZT4ut7FiDe5PHmF
qEoOOhlm7gU9ddT5v56hPQa3SFK1ffjNR/jLpNgVTvNoDlBqDBMLgUt9SxVitofO
2L/hfZ/kEYpu7tpB2oJQS8WXftO5sfba4HkGE1a6nToQSax/KF3AUoc7oWAproRY
S8sZabdRWc+lY/Sn8B56HrzMoFEgyimQY7QD4q4lejNAwfw+52Cpy4xIrUIIDg4S
OjtpDw+VPa2P9JsgvTq4ckPn4SXoL4YHPRk6OpRKfh/1tr4lCh3OELglmW2AnAEb
3yVfHwN6814+Qh/FtVb+i6pWi3ItjEcz+a2+3yIj0+0jtVw8KBHWqihUcB4+RTn7
kfhCFmjT8uiwy4XDAN+izYJ/OnqJrFrG3FXcwAbeHyHm0zGiun4rbTWWHHBLfEeH
CxTcFAG6dAKSDyVJzKPXjkjQMPfoqGlSHf9WVrz4JfAOHCAs8D36sLG/afAclKob
Y54Q3CV2SSIjpjoJ2gfMGyfty3y1gSRgSqAdKXLLSBUqsogsvGW4R+V4psk8jcV9
IcwyUCFEC6EZmf8RjyvWFnZzQ5RHtB437xqRtmfSfr7MNqdi4fgg6Fm3spBvWu1s
DFSDLmmjkxs42DXbO7WUwaVD9ypJ7husGujAAtLpyGq4Uq1svNPONDLjeD3f9hAZ
bQj8V+a1VKcht0CG0/eUXfrN92ghTfG3nevtofHGxiEs2uSwqzXuuBLFCyK30g1r
oIDn1bupuxJ5G+j5tXIIbKuXBoBPovh0zofJN7lju5y2SKHqxuw8nhBLEM147ZLF
u5zOrA1/CuAbYmnQ5uwCjq0BBrhmVTrSck2U293NEQEJUNQ/2eQorOgfzvXAdyqz
KsCyKLxM0oDOJnyqwW7mZqODoAgMiR6XCS9Mx9GT8gVZ0IAUaU9USIIasbipycdH
/VJTikMwXd2QsKP8FzaLCpHiVe+ca9RpWvhKG67hikV6Xk/nb4OTwPfvADXJchnp
cq/gjac5ld4RHIB/g03KPkWSleNFCyJKtWO98DO2O2W0fO5JNhceg7mzKKa1yp6T
Ci96DgU/0n791SIB8IAL/D4hC0siarF6ZDd8ze7YwY/TiuD88W4eT8833F2/AsdA
GXsOV5JAT6oxo9FDp+Ql7hsarTKYoZBors3oH2W+iyJdgnPlB8A41mXA3V6TStRg
lT6mN1eTb+Qvhk6FKnnDPuPsDq+GPe9WVgVEbYTVBysnHmLQ2nfX3Eq77hnrEGcd
xoA16iXxtrQhjM1rhq2xZgb6bUWeBbn6KRT+g7m66W6TvU5u7QjY++f+nYNB6QPj
UIJUJz1y50cpPgSTq6m1NbgS81tOO770tlW/ZC3Gfl+cLlE7AE2Ps1p3spZZuLLR
INGpPoL1cC10R3GujW/vbcmoVZltH3wSjSppETasVwFz+l6XoGJANgaTeH441wip
HwLf8dYFWbrLcrO9dnrSEBeLUVZ7bbJ/po4lF64NowqhD2odOjKEe9U2YdLjMVOA
c38xLTLdtUQUwwNDflSWAxo+ANsCxNcTUHVThpJ1Qu5xX8cHhXpgLdlxbWQ2bwtI
WSQz7TeJXRfitbmFKAOgJnrlIozGAu9LeHt93BqnJnT/Y7wcHvMW9RiQeO9fP/NM
almq5AVnX8CAONMYj8mSGStkpAOMoOz5Ud/osMc5CxtOiogwui2FKf0TQfKoPhMt
LQyj1sREUr0qcAmZPV2G4sBUXXf3kQft0kWIhUcseaEbdEuCyGUhei9w+36T7D6V
vA4BA/MRO3P/1BuqHVnwg0wogEXeWo+6aofwfAI/4yPsG3CMsnYpuqdZNp5iVFsy
Se3foRD7DwPyR4eg2BY2SoLRkCdqMuW2QYkwpzKGSTIr496229NllgFovvq8BlA2
TDLVjBa4GsHMToJo0b9OC8JVa5f7KEgXNPSImcWFLM+CCA+h8kaM5AYDFLEflE/X
tJkJcqL7ssizPQptKsOr/yzSFBz5cX3Pi6rQEBpUQiQ5OYIY8noVA9BcvbKhzkEx
jd0Le1Nn1UAKO/y2FF/6cHl0KOxu0GRy8VvPnjc1/wsal0CenmpbIKTMhW/NznGS
0a8fdIdrMlPnRH/IfPhByuB49GOXt8QSyYHOgKUu811T50AblH6A7XU0xy596wIM
PdgWAOhEpFEUTBYqfh1AXstDm9qAOGHU3V13wQ6t+2vVMOhHjtOR92JFFalvKZrQ
BkMvtauM6Ox8BoLEA9IyxNWl57HiAI2jZxcIChqw5xUKdclJ7Cakk+BjqX/aZISQ
b7085GWAY+V4sdfhKkCKm72wIOIVXdhJjqexCea5NNzBUa/WRYom40kkgg4UkTb3
PElqFJU4VAPaDYSA72/eATBrQkFtPGALk9bVV4xTw4irxuVR1wuDYFf7+65du0KL
xF5UldbYvPOl0Ok4dqSaS2Sc8S8MeJc6NrnkdjQgiEC0VHGDmVBBcQRBBJojXqkG
MA8fsJTGoy9e+IfG7lVauidEbr1kmP+1/tkAlOb2WYe7DP/QiHZjA5AQdS26Jevj
RwoX5BbF7g60IRs6WjBM7y30gjyo8qMNAijmwOfxGnEhei4jKWGAh0l5HpRcqayZ
onwrvyDq5V4lQaZZ0VeB2UDvCBohqQ1XEdNnT/N2az5Qayt0QcLXpPSpdFjxE5We
rJcaala01ur8Z0YwHqFsxTVZgMwcuu8eyPOgNgmwfRkqxFiWhZ/jnkTeL2ttwYAt
kA6ZiODkPGwWVnkJEgWbsyi5b/P55IkQ8y1rOeNWVIporofbt3/opH/kmXLq+zDY
1nl/wEZACRJGXV0XakLyVd28h+BY8qON0eamCLZrmV5qaNgGHr+wVDzOHPUa/Qms
lXFK9uvpKw0dqt4fvWUCbROEyIFD5mB2vVe7DVMItNEvimHmHwPOVWxDgC5GKf9h
RFW1/ofK2DZJodcHIBaNPY9UfTHJpoGPvbVF8kcfe3QbLaUyWsO/Rc2Hm3xQywHd
Vl2rm1bXUcR5AP92LwkFekD1n1fllrSbsedjMCP6EGaJ+2qnNvf5cImQeAj7SYL4
E4C7hBy2n4lr33qRk9SxDshNgqKR0HD9J9gLfxmfSBaEWUcieoAGKr7y3ROswYvR
o6Fo+Eic1OFWjfeB2kQiQmh5CLVEe3OquXf+FMgRsQsBvxAbLnjoSJPzOgP7Yp0x
i7nFi2VctQlLI4f1UvX2LMeizmFqT0J619bx+3XrfFonUN1c9BJfRch4gTkt7ji8
9wABDtWnI204B7VkQr4I3V7kHh1wUcTtwVIVzchzSS+taNcyF/snaV/kyKV7uL+M
M6cb+BoPtemZ5XJudxfozPemm2OlN0blvSu7Ie9iKKFBP7rpHJwCeP/KR6ZOM+z5
3srauDVrYmBiHVf8hTzWRK74I7p/K6mx06hxg/0+v/akN+wdk7B6pxPo+5VtC3v3
PtRFXtu+022p808f03xwlohotwQa1eKt37xb32I/SQuyKVoIpUARopYWCTKxaWCJ
K1VCl9bibjG83AIXpT+DuxKc1qZ/mYyT5OxgQJltoEAg+rBSQgM7uvix4FE/kGy+
wI2T0PrNUnLB7nYkilpVIA7thBn3Z+O/NPb5WzusmoJsDjteq2sPgMLKbTe/uozq
dZ0mOe9WWSRe7fP1Fcudvto8ELbLyhIlekvLOpYpbm1HH9yNQROf00MQiE9YCsM4
lJqXCStFNzSgsSA6j8RnpMWg0ULkhyaozw5rqDOaVtrAHv9oLkgMduDT5B/WU74d
UiZID/tFHd4rb4H1TfgDnOA3mhMSt0enJp2T1D9yCBjspk2hBHSAqX0UdyjVgCds
hKhc+NrGbTbLh/fbRCbnevQCRsU+3ceOyYy1JBh9zCZPgZvkzib2lQRPxzPE4Trf
56MFelVbUvBU5e1epZ+Rx2/vKtFhdH/q9120vOw2rXexNhTFlf/OIUH76V2gDhgi
bA3DXMJEjcyZstUTfQZzq7oPXDpfyEIm75Lj+Z/+s7wqBPhTaF7Y0CH6UqForLfM
Tr4Nmgg8Pmi9S8CS/M4cOnLHTL7Sf1Ncd2BgPH9jfENjgJ+W69GPO8g68TiIC/LM
mXSFVw4CoodKyexAWqcEk8Mtnhhxq4SqcBvp4NN3MnZOZsIUw6py9KCwpSjN54Zv
E+uZI20wliwJXxmbAUcvi3ei4A9v6pcjGF/ROJJfgpt5vIGzAi1MWp0L+lLky+K+
vuFg81jfCLxDI4yvScMrI8QZyRroFWyqdbPRs7ef2F+sHiVlhAziWMfHJctRM/zy
jpxGtaMhY0G53Sg7QJsWNXXHxKXlZjYcLQivH/WSAubVLuMvaBl8iL9MjH5na//4
FALA2VjYsynJE6WQj0wfUhByECDVAhAUUCKUaixefK+OWBIxac/LMg9/yEoEYiHm
YCFifkiGWKMybjcqWmhNSYTZuJmWLGOf7CTnhmg/EVgubbsZVozyxQ5haLgoZadE
pZ61rF+jYFGM6vDxkq3h7zMbk6871tLZTmiSuMhwOvCRa48D9esfK6E/nuTDGfLa
Z1k+tqspmaObn4fXN/WRN8SETeQGuqI5rF5SmjDRgZbo5x2IFqdVjrlFP6CPxEbB
kFWdVQOrezz12gC1nvTWnhOsq0ohudV+7C1p2lsGH/h3vJ4qhSWZrvTFmnUgqRu6
EpZbD3U71XUwR9FZiQlXHkBqFee+VheVlz6ulqhqJdx5rolgXIq5jKX4TswkF4rz
iu//TrsarAwwKkndlm7b4kudwab35D8fZ6JYsiZai9+7IDK34Iiwy6R/9IB0n2NK
tlHVyq1qxMOffgjEEeof6Yd9cqk/cEkZveE5UKruImgYGkOkoJHhxk05lVH7S7gb
VomUOmcmkbdjaKYtihcJl6Vg0Qidae2+n1cDkiSVX1iQko3NoAVTOB8Xs5o91kvi
zez4z4GAJ4oyk/Tvq9JPzfo4JmOaOcj+vKTsi5o+N+ycvGcKIGv7LhLjsyZ2Oeci
RtYRQ0JIft5T439ZNRMNAw2Ypew12C7nKM4wqQC4fVuyNzoAdxbyZD5zxN8GrT74
qQf1ea3t2jCOdJip1HE5Tw9Y1El6I2CneN8qxMovtFw1G24eXnqwwKUJObV7zOUr
N1fs6RSNykxrSbW+ONs6VbF1mQIHsUGCQ50fRge1k4e90Msr7UoQC1HJQNdvDqCd
AUrqT8lFaVySDDEQJ1XCdBQ+QYGhiy5hOZ1OtMDv5rbjGEO7sUSwhG1Vv8Hm4aWD
1ntffnMQ37PimuYv4F1aeMB44jOL2USW/EvaMXskugdoVBVB3hfyCtn8o/DIefXT
AN3zP14ec0wNlLtv6foHZYQWt05QBU7qx+zCfFQZ7mtfYllpAuQSRAk27qt7XcSA
jIYwzoOynvuXC/zuhXdBYgxxxDCJvd1IySBek1ot1mAWTCUJF25At6nfIL4KTw8w
ksCZwiRKyhqfqe5plhYvcXqKbpg3kVshlZU11HIeCxSO412jkNfqXEybMavbNj+e
5oZFq1Az7VtEkF+IhW0Xz1z/Vn5I3/VKyABX3rMdRC9IjpOJjIt60XJ8nNTSBhJa
f+c7bW3DKHPxyulQic+2aKDKmHrVZ/jso+jCtcQu2bzkJ7nWkETwbg6TqfXoFGv1
2yFnHNU/yBH6OtGiFXKGidpLZTwA0HAFPq1zEtd6kYQyeVmLo05uCzpaejXbWsbr
90BX2ju62R2VgxHoCNnIvWqVNAXjntmqota0BCeNxpKTbQ3kTWAoZc8pke4ByESs
AJvVzogWwk3R9VJC83UYvxLa9aISeWG9vOMy/MbOTZYVGtV8xRWNZ9SLFu9dXZcm
mziDIlKqcv4dX6K1RWbVC6UhpORQawmF/W3pkjI9vglnUj8awetoO8kNkyju5J+T
Qek6fpYUx5iAzLJSonTjrzWB/KtKysPOA1M3xp4rsNT997J+CCR8ycytNhh+rDXT
WywjRLTwJyO0HJE3MxhWHsdYXDJTMXx/CpPCmxx27cJaJD9bxFBd2hqjDQ3G3KvP
h/aTavnjKIOYDKeewDDbuxs3nL1ioU+1zVaTNtChGSVFY792fn/IN3bgB76mbQrj
GGlkz9Zzl79nYsXXS7eXLuRZmA80abUjJNJsLG7sAmZb9AwDk0oF1MYWCR08Eali
8MMbbjFyaJrTZbzz1eNaDTe2KP2wWSCNYT8R30t7XbHz32BS6LWh5/UIIOstVVdK
PrWCXZbcSuGmAfY4DrnNen2vr3E9ttL5SBgAwUJwXzPgJWaLF93COW94yI1Irwz0
yzu3dMeJM9mfZ5JjKPBv0iZrDuQU+ZF7gyNUhPf/WVoXhrQMsqjbly48MrTlwmA8
SZXYPh89u3V1JPTqMle+Ci9AD5JCPOw7QIdntj2pWYlT9ogIgrsGaOGCEufJpxQA
uIgoc6jLwP/a2UQBODwnU2whlehc0GSnmQp49ercz1Pwk/gb6/OZFhA9AYTHZSVp
F/nlLVS/Yb7Y1u0Hr5em4Oa3ZHgleZbP/XJsxsfyTLUjTOhvNTj/5wZayND3TRsM
WsLesvXVvmn2Mlt3iNQOJsuksyPKa6rbSDTgoTKjPQup//Zv526Droyp7T3Hb2D+
OVm8YkRTrLp4HeachiEk2+/RDOuLgreZBcrZ5y+sRtbFSOrKCJ59TIXbPQhGnWJg
ARvC4M2EiSe2/qFu3O+pBu2LeBVhhnRwDNt/7O/PmUOAlqroRChe3qWOkiBLVa9g
G85pu9SLbJ8FhNtt/1gLhBKmsARJ05Ei1i1J7DRm5U7GZEX0Q3GfoKiu5rB1OB55
yAaH0x9OckVH8aJo+4WmYh8Zdwvg8dUhc8sgQ5FUuhlhCNBgkAHckTV27L0D/5PI
jqtpwjBLpqA32PD1NZdrhmQlKBKvYUHTNZ5/X7K8sP6zzS4uQN0WX0h0MzGf7wd6
+xNxJZH2wSLv/7mHXxb/YLcQuxLZelrwNv/hONufOP1szvqnwngnvhMlHiUSVJEM
ZXpW9Tk0vdzg9l5R4t3A04pBp5fFr4KcvtM/MwQ+EyudJ+h35pLHw1vWKNrbj8fK
5fgDRybtL3FZS/nRzLWEIGp7oH63eCKQqzWMCxvusYeLeVxNioZngZM3al0thqPV
YA+3fHbqKcteZEwYKXBjcmiz/MKDFFvlxblu9xnW2MM782TkNoqTOINqXGZZw8TQ
Cmgevrfb8wPHPwjLQN7hnAfuEFWRE2aKk9+171SgTy4cUkFPwL1sE0AwhbyQUO09
cUTlTplmwtaMlo20GO4juYS3y1ynGRrteQ7AQJKtVFXY3IyLyUOsvHe8lmqgOo3E
VF/VSoNdmDPCZvlU6O1fvL1itBpYn4xSf0DRhxKeuQDVTkvf1RElIdbiw0OW2+mQ
v0qw/2/XyLB52i66+KxoAXOxByohhkWOIoOmX8WRJxotAJiOjSd0lLuO5iiI/mVW
UJ/X6FuulFAmliVT7TKZh9/vJbpQNm8RaBbnbDPiia3Fl3reUlR2cfeDWU24FBHm
6OCOS+xDE5/FZIK9ylNUa1LAMbchy1UtBA6n7q+Il8EXaS3qA31LmAAfKxok8Q7I
LSfDgs6XvAsC0l8dJdxSfaMUt+sWsXUFHephmnX1/pmZtcaiY0+V4B+ldPkdXsim
oxd9OpuQl7YbaiVV1ijZPCmvWRdfbCtVmmapAD4wCGpfb3x275ZlVjp6UCItNz8L
13yXGm4QwUuZ9EwPXfV+7qQ1S+j1DTBaqs8X4I2/cNO5kWPmnQblLcJ69WlMShqg
hMs+1ySIjXtSb7mY3/GpZq1VJbQk3y+VlSleKC5gV7Y1TJSB7aOZ6XWb+5Ko0vZs
NphkMFzQWKc2c5ecJ40y6qPAx9KJJe3cwW4FpqfPVfmlNsL4Y2G1IjBCtzlDqk7z
sw/v7X4C4XulhzMHO7ouugDuibbB6C84Am/FYd/GOWrfJQyqrMTY/S0MUnnCJlyF
YamTRsbQI8jy7WKXgm3LcVa0xfNcXXXNuwLXX5VKMkeBtUS9ZaMBiRTyXa5TbHRH
mwH9LqcyXzQgz2kQSMNDQFD/GlU2e5If2WtG8rG9ufCHnMUJEJWJJHDTKNSLCVLT
HqJSCnyimnha9ijsPozQklk4tKe4fJLOl8tteu7yNzizrXB8PvOUpOrtem+OzFc6
16fdYYKnn9RL9exLGeTuiJXclW/DOsfvx06CbHSQCfBTepB/2NbdYGGkyAg4td/z
2tnlchqML/qPbayYRqCIki1j/rD0c6T7texR1ewFnt3OSmyr/66npIp3slR0anUf
uHtvrLcemgNt4JUYRsTNdWQkmr7Mjsh2L4om/kFOjRYTzPZPQjA7u881ojzfz1at
v5wXdoX+AWLfNhaviri1YLmhzbaXvTwY+9KKqVn0VEB+GSf95KDuJAU0P2/kVYMI
12OC23Db8DGGP3r74EwnrSIlaJ1cTZYhwqNhCB7uTWMFhF+EN/1ZkekXBylimeDM
8Lx4bm3P4PmLjkNkunBI2YLulRs6xNnMo9z40f5FspjDGyAgA60sxwLZwcXaFMns
plgP0CpzNB6H9AaaZsTWGz9Do5T7lQ7Jr8CFkVwfpMEnpqEiH+anod+wB5LX+AgR
LzKaen+5XUOgRQiF/fIpvT9iy3yBc4gUfhnGqb7P2pt5DvGcxHamsmaoZyHs5j9z
sTGuPLiuXZ4vXMZDSjEC1OazUyVZofagl2S5cN80WgfAOF3IvZ1UmrXQCQr3xn+4
pyWuFLmFSHl3sS9aYZ9Sg2DX28aTgOFbOSHNPdkCLzng+vPCjlMH+TyPGkCoeshJ
ByJ6SFv5bGUfNkfuvosrBbAocVBEMksWF+enOF+X0kaTleaLSuMkqt+YFNte6BPI
CjSfF0uo2kujAG4wc+yVWys8+GRGbZXrTa87MOjOv5nTRHGxq5y63hsT1G/nnnv9
kiyHrZeign/G/pDbyFD777QojdZxuReZ85GyPn1K2j8tWmFpArWbWLe7/pPpaTeu
ghyrej4Vqv6AnhFKT1NUvbSiQdcwOIKKv3fqO1WYDckocCvLkYmjGI9RDxpK5UxV
jtU9xKGLjTLfiCTUnfmsu9cNKh4DvDl1VBMgaMWCFA4QX9SRpZmoh4mb1f4xkiqS
fSI018S9I/9if7Zvdbv1YWDBFwAz3c3TzSEkGhXCXewpsu9PJVA8TR92Hp+2ZNWF
4k2MoUDeQ19IN+QBV3l/eCrwv/TGL9thcyu4H/ZAMxo+vpnXx6QzrTmFsQEYIjQ+
tjAKnKTOTjlC7ix2/JfkbhCCwlG67KlsARqbyBwYiO6VDiMXhkK7yY8Pv4KvWHdQ
XpPZtYy+CB81MD287Pvxw2Yk0nmS9PhE/1NG+LaATFt033SqASLfLIhhC6UDSK5x
U2xpcwjCMjp+1IRZtFHMdpycs6Ii7Oy6xnM05oDDeyEat+Yi+9ABRYEyjCiGb7zu
Czy0UGx7xZimbpcIBF9IMYiIegT6XSe7SaUW8FeGMJIeWO8/3oG4N0Roj4O0bcbr
7YnVXOlPBKpdc5lZ6iVsffEH2Yo1vGRs5hUYEVEwcf2XInKIuUqUPeZiCbg+vOsa
kUGxWfiMQ8CZniyzJzZ84YdmN8geoJCfYH7/u2vZaZWnyUBFVKDYubJpPsUKRn3a
8kJsVoGsrltg2HZYwkoYyxJkmGVEDZcEXSDH20j1Vj78feHbVBuHUAoecanUxYgR
krQKaUK67uElLeKa/mWOC3xZYdv6MKefdhA9xJRZeOwg2DwnlSNu8ZtT7YYT7Wdm
HWChY3dj4JkS4DfvkpORX5mkOUW46qnrUI09j0RzcC9uEF3iEpZwCGa6eTYWmCn9
RIH0cFlHvcq9NNE5a+vzwTj2xf6soZjfpaz5UL6HP0gEEHpp3nFKSBzkPZbfb1mN
uPJO1/lfGPw6yXEOgjLSkS3BbqBPJjdjXFhFyhlSuKBBINT/sf+RZWS5vXsdAfzT
LvSJxO0bOyjqNdrOsv2C1tBpM+t9sNNfgP2BkL08y+L9eEKCLQZgKVd6gY/RxzGx
GeXa6yinCdz2n+V6lXATr7Sa7b9odC2JlCodKu/MED6ZJyzp0eLqxS8K9MeqY4Ms
yNCESxb09LW0uICpUYsXbKQFqUYQVVR8+uHbHE2AkBJn7kThTUbPgtkVngaZ/02z
ivttqkrR29+YknpTjvl2hxqWvqMWSqOC/3Y/V7QrBTVGINenKCYttT00HXoL15Ny
5ntTV/F6FsqywuR0Fmlvuu3cHhYu/oxAElAMtUUk+FSXG+JmZ9mwKiNv1JHmuyzK
1AjXc6ZvNBLxGNJ+/gYw5ybwn/kNd+eGlBnEMZwRlg0LqBM7TNHA6IOXeXF3SYun
C+FWRT1EvKDDJSS1XOS1CU1nEty5U1QtbAc7bOmbhbUliPNwwSYgPK8y+UoMR0Id
mtsdqStaI7UdivXAy/WTKDKoPoft1icfl27ZLPvLmeG0q1T6++h1LQK+Mslt7LX/
PlEaz6Sefz1vlwcbJ/WZclxn7LRwRQM1Kx0FqwJW8WwBPRzJsAwe5+UBsBIMi0N8
m7mBO59gurru4a5PBzT+r3RDQkQEEDsR++Uh8ahkNTQ601LryfeuJ6FPE4byPEKm
PljPYRNvYsoZT8qqQaWJk9sWcyEFOeDyVN/gOUOeyWZaaHdH85ynos1X6QHVDf04
G/i6CJ/inqwPTuanp8ni4wIgjj9fIwkugP1mPxgihH5G8amT51W3tmFUDZlNuk7k
5n2tFHL1H1OZXeleZkyYyvqxZYUYToRfOa5qqYfn68xsO/NmrPm+m7JMev9gHoBq
2Ha3xHEkMZCdZgs8Nu0i8WHonuDtxyy6qBr5MTFBx3HfBi/ZITr8sdULTcYobCLB
MgvCAB7od7UxbU+Eh4Lx5l2Yxf6IJII+F3S9UzOEhtgYhC+oKTP5K15oUJLHExP2
C7CCFyId6YxbTT1DtWF1k37GeTNp44+el4qWVAMg+CfSluh21QQAfKl0TMw0zS/V
y7gzG/G0ck/JSa+c3SJ+LZKpW6PtxhNAFjTJJ2orPQuQLkC6tSAuiibCxBlcjoEw
TOudUlJfcUH3reouC7DvNguOhLExNdz/UyK9vjiWuXwjau2Z0rZeiTebb82SBP7C
+U4pECcKpRrbdEpn1HhoF8aoa5tPl7PMAGnVqGIY8My+eqyXeVnESgC6/JMOn16i
wZQRXIzqhvSeuPDRHYr6FC61JRCMFzAb0gaif1SaH9LtJxYe8hnEw//K1v13MRp4
9ldxoY6L2tdeqVtFwiVRtxZ1t4YMwNd6zqAegP5V/00kcXpObHigM/wg6e3JvsBF
95o7Em+z0D0YyejH1ENS40Neq0qTYS36fNEtEDWUhrB3pxRA6eWW4y6HcwF/YUrb
eHgFl8RCo7RRzDU8GTOseCrOZaeHCQHNT40ipy/GlkqMqhVXCmW/w43BBWtyWKVQ
kwCHsZP8SjpKVo9Uwywv0b1cthNMPZiZsQnh611w719HlDZ/eoQbpiuNkOZObYDf
1nXyyQs/1BV1qlU3mMy5iWsyyBjpwQN5wXUEQinGCfwULPyqjp4xBZOGQbKPdKF7
2boXSRiRSFNYZzgBErgfJ9hU0qVTXZul3yxEiSsF5Iq2N7NQ/rYSCzXY9oRbInmP
W8udm7pdRMmMbH4yXK2eKK6gEK11TsVUSnqXFxBb7xkQZZtz03YYE4/1nHQBmuHC
V6Rdhr/3aGOIw290cx9fEATfJuGl1DKP+H+UUVuYETP/pEcF6boeNJGwWh/b1GnB
LLTR/ZcKa0Nc8LkfS6wAwrWKq94A8UkA/euaKdHhCHjb/VJBP3JEKat/+XbCcnIM
Nhclqtj6WhMQefhr+o9CxZeVE43uNk2bb4yrZJYZZsE8tUld9PFv4UJIUq3L8z0J
eaDxK1wS9xtkRAYTS53FJcj7F8ptAfp9A+7MkhN+0h8BtcgI5u9GGoVRPLTrOsmT
3A0vOuQEjp0klZEyaOO8lCjeX197jbtb70d4tXIQvPiUQgKN5//1r2GXDk3gsP3B
kIukl3Nsng1DY9nA9CWU0x0nyNtqDkGKUCRT7nQWCkbJPXulgSx9OosYtCke/+hG
sX8OmxnONXXOoRulNLTG/iFO38AKfmb7wju3UM7ze2pNzTEDAZZi80twaIfynilZ
7k/8DO4y9wDn7hOdUt1DZTnQo9P5ap4ObQ63pIyzTeTg1Vm/A3/Iyb9oTl/zCVAN
9zZuQBQbvyGXrJS9qfqQC3D+GJwMZz4XCrRPKLrhJxxaHjuerY3LiM0A6OpzZ8dU
+OuR3Q3fhllhNufTSE/V4sGnauJh5l/YAxDjDEaRETlZvZvAeIibLqLiMZDOL4GT
K27Kl0hwE3pjySOVzRKlWuXKyktGWxjb5IA7pxtSdWJWuN+ZLRAkB4T9BqKar8ar
sByyE9uX4TCbnNqeVJTtivrgvg0NRLNVj1JsRb1efRUpWIgmFFmgg1u2LE4aoKqS
nLt3SJp934TRluc7iDnHH5440NfqoHW1WeXCZbAfh1odh5AddaHYeADM8azCCxN3
nzZ0ti1IEgKNtnwkD5fVFwwXGG8IuPKclbcLxQTjwmuFcQ7wgGMkiNPcmFA0BK69
D/Ox2VaSMtfAqAF+L+lpGfxB2ijlmI/56Md31yrIEOn2Qg0wmcYyBHIqLfWvLv7U
yRPh9ikVDaA0nMQJ7tttArh4Nn0lTpNkllC9F8w0MxLKk5FChjMi59272QicabGZ
LPIY+kcDIsJPGY+C6zD0jxlxy6xwk1V6LH+vgIeRa6I1qdQ1ekLJd6aug8rvGwue
5QfXg0xz2MSRb+6X/oNsGGDt0Z5gmYaflPDSu1qrEBYb08F2pweAct6nHdalIrbW
XvOtGt92/dDsl61+XZuphCsWflF22x6Xoi1J2YBuKix9lsNkK7W+Ty+92R6ALdNY
Y37hy1o6LC3Z4g6KOrV70EcBt1dOQOqv6ZWd/jq4aTlAZid+qw74kJ6rpuoD8htO
SAgA4dTA7JF96vuLNILdnMIBtqddciNj0HK+CXoWw8O7Q4SccuKASltI80wp5UYy
x3E6Mn11h+7j0z+EW/bkeYMLrv7zaZGfYI8gmFHeHj4ICtG8Xj1fM/y5Twt8/WD0
Hop2i9Ajr0CBxUTNMCJNoFud/ZILNZwDiPzIKEMcO3XWqktqqsTWABXXNz6gC86r
oOr7jCQbu5degGjQ508hJOa+xnfAJRIw8uq8JuJKC2Rx/NDZGuEqZtB8v36ukx+B
2eGULnRS5GoltQXObwmrA7mnNFcJ/cJ2HikKHoX8zqraPCNta64SZICuFCS+Uesl
aecDECqt7orWMkgvfYuZ6xC5vxAqI1TEG/xrpWWD5f5xpSzFU6Pe2TW6RKSzsMVk
t/0L005xSqLbY8qFgxwS2Qyp3H3RmKoJFc76rXCcMhsCAIuXGAe0ImyNcmjoONJc
gmD6iZ9Jvf/z8jM+HweXQ0k5FHNqImLgrC/kcCWUowRGdauTSrImwi62n15mb8RA
p0dEZ/kJ8yEYbbRjjMQZFihiBFKieqV2epfvqPB7KHcDWH7RNpSsQ4yaU3QrQPyI
9LSe7lQBuTzuj8gm+hFIpqyIx3trRRhsFea8gqTJdy+TZSqp6gv+nbXfa6D4nrRV
3fulUOm42lNZNSq91KNLeXxua96ToGqxznp0sbv2qRuLToe9koiAUzNdpJN+MXHF
N9qT9+vxDEXfGbdC3bb9Gjih387N3lwKA35jHSoINw6GF1bND/5/+ksuc1Xdp0Dd
WurR/pim+mmkHH3KuMEz6sGfHtRfvOJLe2vuG9YN7mLceJd8pDnZNr2jQcnf2xGA
SeKtEGXHoymHuz+L3hu3/VHf7TzA6ubHaQ+RprA4f27i5iU852tXhDgwKIlteOPH
VYejxYgGw7BjurNOGWL/HLgUuY+beM9ZDizT+3Y0wC2d6bEl+px/azia2oslVjdb
/nYJN+Dp1a6nbYGiGK+0vLSF/oIrlC5HPqb61h5Z4YduVkf35+0Kq5NZJNRXVyvt
3KbYJwIo1rim7NQQUJVkVOF4akPRKMk5OpBX4CNuAmOyKgJnpCTYC12js+2Afezm
uD9a2R1IAarn4SlePCeF078E53tFLr8pkU6mfAThyOAnYJctw0YrIEbakZvnHUXb
0COysZ8WoMt9LMxxAa2zj+A4E6G5Zi0N9wlWpjTt00gVkV/dm6M9kVuTwszw3hvf
AsxYQKHCPscEAozeLM7HQb1L9w6YEkgbJKGICCxkyhX1FOx9QGnEkVawQ3BJf43j
Nh2lyI7mq6pZDYL37GLF+ZCxwN2T5SGNuFr2NgbpUpoHPd9RC6uG7rOiQd/H841K
tGFHDKoZDQDvI78arhV8/IF0k1ApkipqDKDdufEaEHlPcBSvE8lVVWW1bYHvGphl
8x+0QGDt3VyUEfEA3eMxJg==
`pragma protect end_protected
