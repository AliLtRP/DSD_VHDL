// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nkLVXcQXaxwc8SFZYQodICkn/nmbE11wWbwLkdxDdm6MY2jQWtMvzRA5Q3et6mAp
6gJxgCDCuLq104S5BxOc28q56q/Wvcng354zU4+vUrmohMToFmj9z6whc6morFju
Ya43uUo0C86okNp9MP12fcpthyuLGu6KXU+8mEk4AOU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19344)
Wk7CBu9JXQYEomhfCBaL75eUIPFL+tjfGeEifq8kp7m7DJcGp/4J0EGUk/kedV9W
85zdOyajlBnEaxE4j4pdEyd/qsqcT3nLgHAB2MAqGdrxbDsSC7Tdo8BgUXqY500e
tVDQ1LfIjL7Gt9U1FLs3/I0KWj9IDKl4/PlMOWLW9/3cJTiVpiolSEg4/kprmU6T
4HGXJUkzG8UIa7tCsANdIMsZNBocqv+QnLrsFgQnNZLF4e64VM1VGFni3z4tn+6E
zD7cpMA4sLnKLcDro6Abt8/+XDX6b1Go55PghewBqfjqutNDCwjlAxP2ollx0TBB
MWH9RicnvdvpdCFp+Ajv2mXTAXXx0DVP0ol3gZPOFsXY7gZQYlGlFL5SIucIOElk
JorQY60uXgcUfvX8AGiKvUSzvDmxoMO8SCR9Uuf4a/kUOBgK+5QysX9B/if1+EPR
CXA/rgmmVG5Ph2HVsRNEE6WsWaIwpE3CtTigvcjc2hjck+cUnXHoKle/HlszOiO5
uRcaQc4I+2wBDbUeZ9fcyLDoww0OfkyOMauZ9PhDEltdywhUucYFXb1Fy13r+lWn
g5/UXFl/VBnKWtKb0s6XQcdJV+PdFqFKcNaYqOw/6miznThoDqadMCiLo4oKSTEL
V8OlALWSt/gFRRuVYCyi0nE0nXQBKMJCQU5fMMdwVStG+8MV+8oQwAQD7x9mvR54
zKpVQY4g9pjOpxnB5eAkfrwhjM88gm/441vlpDEgFsXGSL+WXxXINPq+DRu3yI3B
fdHQHDrsrIU9owBONmi5LOzKAycgZKPAgcLze5lZXmDJdiRqJgv5UpuSWcQxQGDs
QEK7WOAsqvk/ee00bbQrec0aFFdi1HxhSK3SJBP/yvehwnDZQN1+UCfM5fG4H7s/
UoGvWBtVaQu9Y3YHQfVLBDEbdtSr8bMUFDt003w29ZxFrbYbGl+BE5nYDWITBUvp
J+Qt3DyfyNydlAAGCD6S1yjIDOhz4lD5vwZ056nAc2EccxyM8CmMley6mL2iE+4N
1NWmCbYeZzvflXTmEzsRADRf/sQdoXEtWG2Oz6LS090JhEInUeoJn2ikiqw4ez+G
tTIsu9xZpGF/ROczBBEdrEbb3Hb9DHlHYz9dBn1Exaozm2f2bI+J3j2ttKaPydKQ
PnfH2F0f1Fcwq4ZyJP6b8RekdmKjOOshPQOrRfAoeTn5swM9yzmSRGT+Nog2kDbb
TzcvIAkm+koIEh2F90YedUxS5u7NmmjLFjWFAfb2mZf72xFNAVa68eulVaZeJHNG
UHY3mhfUzh9ebvOfHMo63tJt6bUuBGIK3Jo8JhCZtveDSwt+6nkn2NhnCHFsFJ2t
ko4mzRbNcrhJKW7neIu2prkL+3NG9Ti5zMaqbhIUTr0cUu6XS7y8lbAjo+cLEX7j
xe3yhSJ7j4vER8K2IQ733Fo8UiKP8D1apDQBEPsSv9bypgV7uKfzt74KOUBz6Pun
cgb7uPqX82C3CG1ZGC8O8yqAFtdstiUoVa86nPF7Jsbq87Zl0RzRu6B/Dfrg1wP6
E2Xn9z8YmtXP2OX3v4D8/QBA4HuayLEQJUXWE9A6oifIaYaMN13H/sI/8fw8ieFd
LiDJZlkFIyvz94fukHH0e3RT1Z4W9tMO0JoXE5J7KYfVRnWTimXJ9lnosnSQ5Lmz
y9hubyRRkUUQP98+HgclBT+w1YEAvpr/aO+shcCRFAkGJ8GfVv8hm491pEa3SKrD
uU3SM7kUIs5NQrXJ8dKyiqKkiB/RZc9NdcpgizE92rI2IolwBRKsYKp7AEoc02WP
2i+hhhiaObfTCWmotJRC345Rso6cqqCXvdPM4thzTWZNQUHY9oCtAt1WQJ4UuVrY
OMU3+wGQHpcieIA8YjxlqrLllFq7OwuGyehXfJ7ALYWtttk/3D0MzktON4EsSpw4
OhmUzJnKiAmB9VY3qHeuYPzqM1ZUPv6YL87eVx4338gtacNUgJeEYckHpR7wpfNf
mewH1rVxpV44MgJf6ha0ZqK+icA4rvC7NTHvKQzazEXmvgYIPK4JKKNuMCr6utQP
Uy7bAiunNG1K/r4lJmoYscNFM5ua46B9qpRtSKNT7AZzB1zfVokVc2onT1o92pl3
uzUhH2zWWxlNvCYZ8+RK4WukPd107WK6hzZfqVbw0dBxFfbOo9MgIPVgVCAuMr/H
NHIZd8o9v98eViiQQX9VO6XZDBiXhb6whqHLSWh5zMRFCqrdL2sGTSuSGq+NqTAR
Oqpo8UuN7rEKtXa44d5Fn+9DKrQOWXk825aqJJTfvwWYCBPtZhYU17dPI/uJXvuh
+EV3T8/YbPW0wjhe0b2Kj2X5E2OAMgB8MA3cQGRg755IRJIjUpr+JPVly0fRuvU2
BYb3oF4p0jltSbmT+e7c4dLTZ4u9MOXrKscCvfYaGRlfTgGHcV4CEPGRjwB01Eeo
2ED59EqmKyTd+oBhqKWjpudqJa2NUH2q/kYSkAzVa+X1I7vQ5L6NWtFkn3IQSsrx
hM4CGP0QnlhNY6Ng7NxxyIS6oVMAuOdkQwYcFE8VheKt+mI8eiNDmsU7Ehh/nNrD
daYv1eV7UZgwT4uZT2zUqulocobvZQQwJQ1TAXO7yTQ6JWiihTEfasBouoc5pLBX
ROpyS/VHpH5Dewg3IG1WNCBTEhFTxFPT5bdqdfWAWVt77V7xaVSrkEPltlJ/5+9i
BlWMeXGd8ktm5rjYk03Bzo/dVKetC1vFQuUf3topC5q/0b0VruS5rpDZrpmjxjnN
F6PsJUB8V88G3PYh5cZZ9Wzk9NrEc2iE1IC2XGwArtmUx4x67d948iAkpG27BeeH
DjCxIXQXBfEMBnu5W1nVLi1yAM9HRBj0ZcgeWKQr1L9HuE1EFjsgbE+yi2hAG8w4
CXFm80BFtzMOsZS1uOeMKs1U8pLOTJFkEEDrSCHhjzUru20sTh87/fTU6mNA29oP
pn6gzy1PzfuNX+YrYYXb/0Nj+b6gl7QuFmi9Azc0prptl1ll5ajf2BhcFKS+Xnri
VQ4AbkVUJwMzlb19apKiUHURHrdQgRTQvOVsEWB0Lok3vx+UA3RWwx9YKndABLWu
ihpS9EklyWv5P3UOv5nkusZZ4lOFEQfmGwn02cfT0JHhLG6LHR7F2FoAdzAZDmnP
93kosk6fz/U6VfJtF1wKe9V2Yb1GlYm4Z4VqWb4w9wF/DCLzWl/4DajJiY3Nz5nb
dXRMmjY+51LOuaKZiG2jCHh/G10pf9SyhUaY/XZmoaBhtodptTJwi1WWAxTrgalJ
3DJ1hXCXoaWvT/RdB9OFiRKTic/CCUCyeRMpPcB1I8YoMQIPDYLcJLfrGUbeUmWd
dFnS0mRC+0pZDu3i7q6LV2neQQfYgWSV/iGUKdgcqeqzIfFKDIVSLvoB16CYChZd
1JeFkgy2pqzwcokNBx56aNGT0YBVba0jy+NiddGFDwxkfzXgGCnWx8XBxjbp9Ve2
ybshiSg72lZ69uw/yMld2KQCZaAE8lAi6XxTNdw9zpXWnP+dX62jOXfpx4+qHkw3
Rv+tu9RIX+zl4XHm2VPVzQRDpvEpOFbfZv/eqRhE4Vyjzk7x2NvjkYSZmVFKjLhp
UZTYVsjz/KIcRcR4IBXmcHWYSkZKE7fUJloHdgA9AsPfgF8J2xf+ez5mbDq7Dgsn
ANT7yrGxLh98qlLn1e/6bpVHXxVAwLj2bN+cmlenvjBRP59fk8afwaYbyQGdvT/0
XW9HSmX68kBVjelSSGd6TDGCL/WJYa+/gqTrtoHkkGOTwpU1Y7OPH2t+5FIOw+En
JQSYGz++vOWYECsTG/RHXrTZXt7TWUbARwsEm9qKCm2tk2j14SDn+HDU7DwOn1OE
JpeKDibHPvvMkM6R6HxGE08n7AeKrhf+iVpSMeciJoyjwKngWdx+tzrE19fNdhUZ
CP5DQbw7udQ8Ex2wIvCu3DFwGaTulh4qdiQX3r41H3jSv+yeMH+lNel2kBpc6xJ7
3nzn4eOSGFKeNNPHujIKHAOaEGVj0Js4i56YSEnNct9XT7ZgLVuXenojoTZyaG0W
X7+YKjz2p+vAXOabanxSMwxsQ1PhPhi3UnRxwZzWNuEhQwmPiloxMKl0xOh0UNqx
mHT0eRlPFZLbOypFxjTvCjZM/YNQRVTKMiApuNUN5SbAQJBL6luWAi5bKw6959W5
YbAGpJqvZQvO+8gIP0qaEcS5RXPXLO8RT/O7vfqn0QoyRG2VTazbwoc7dpj1W+Zo
cQhsLBpX156B11ot6v/fqmI0uLsCbMC0N/Su2d4m4MyVeDlKJQneCdaJ6qJWrfSs
ffBpzUc5/IwkMoPowqCTTKc3QKvsqhsbaJHXPJtHDOwpzkuwohQ4OB7T05sK9v0H
R94d0YsOJzs1nffSpRrCAV4sojDMk3XBoLLrfVPk1SSpVYg2LFTPUFDw1FjkoBts
THxQ9xWxZurnaekwJU+TrDXiDN/bSrnRczo4D4MRMFziuTukTEqhARnWP5XWPkha
F9uuV0Mj2m/EZ7u9bT5blC30YH1F8+PyJ9oe4drTAAPVdUZ5eRxCHj4kC6WcJFU/
/OgRe00EEEAHAjgcrMq3vek310SurhAxCXGGwT8tZRPglhkGRtfNWNSuXd5tobHq
NJQmSvSjD9PO5U+tJD+CtL9I9HtfP/xSyEhz7BZ8MWo16AOoeTokZGk1FK3SqGig
S8Qu5NQrLyTUktcRJ0RkDyXwUZnelbzZdXvMSsfz4t7IKhOCqB0V3jN2mUUpKkk/
/kT1fBeMSUGezRgHmLT+jxx9CFkzlLXnQwRg4gcsz6U9mf+tR+mpFMc1RYUBpN3z
55RLQXtaHKZV1wASlUZMw3ba9EVjLV6yLavoJT3xhkH++HfyYlcI1SOe+l4nLK3S
ViOiKdahmwdK6hUexdUCTcYbc3RXTzGRRHReqENKpP71+Y7LNNxjQrIBA8yqnn88
5Nqy9Jlhu/6YVZ307W7ZqTq7OFNtp/63LI3OL5e+bTp01AaymAE5vbj2WJUZfTYQ
dAoCawVfM0YPr7BOk4LZb12yUpb8KOvg9Y+wjDKPVFIa/idgE6eNGQx7nGrwX28J
pv4g725KTcarDB61kXxZnJjWs8ea8o07QvAveUSmeCT25XysgDaDAuhrPHQbdOqk
4Fyed+mBODJJ9TI9WOlE1O9u9gREGObWGd2T/w11YxuC7VNEcsX3BnhcvpmJzrh5
LUHWcJ0r0IBxQ0dVk5MoH86QDFK1lxT7i+MaPgbYEwFXJ5SNYpxVnrCgMxGIm9fP
JzOfioftV7EYv8Lv7FkaDYb7wA32DSfpMTotlpEb7OSPyug8SoH+9dU7ZtB4U5Db
XtZFrmv0D6aNo5m+Tqkm+MvGF752lMV6t95iWkVZfHRMLGoyCHxl1C267U9Jcz3c
lJggQ3nnum6Odn0lUGW9JzlJ1q10TghOc441rMBKCspuu4isuPGVl93KF1/VRVVy
yZaHMiu77f07C8rJHOrSm/ItQ7fLZO47WjXj2MZ5eQSFAHsOpP9Pv+uFdTIM2tlX
cJizIN9ckhegyGD9sUa/cdZV6B9coc7ChaIOO1BRFP+t6asuEPw7c2iCWZPibtPB
rwkR9prcuUi5hjYDgRb0YDmo0tw5VL9sWV1PFikAu+7yFQu0GNXaSATpcGU1UFws
jhXkjsupitXRYB41iFrRiNQjQd1342pWanT3YrjmWFVh5bPjbBzBAnQYbnqQBNsd
fOTwq1IIkXFmmvz7Z+GMHNECKdAa+bhUbzt/1JTH8Z37Ix9RDJ13Vf89hJU5SnWl
D3bypdOO/iNLRYpBaLIhHDt/yflJMg8JiLM2fmIBncgPME4CixFkZF3kOouKtHLh
CrlOELehydICmyE1bHaH9/QVk4GeXyifNXx5K7C1MWCXmhtRbW0IQLmX4hGFTRem
bz58Loa1MYTYABm1xB6XUHahY7v6gOVCTYndc3hdNY0Ub1fy6pHQGpnf76qndAlG
IoUQfpgGcQwYhpdM0IYreG2tBnr4YatF+gD6VKisMgxUKKLucQKuZUksMfqMT1Ri
2iK8WhB10NMjzsLWYvRhYWNRWB/GUCWvE4IT6EQp8oN1CXnrleUjKKyYOHCCTzFR
tvJlD7V2YbGA9mNug0OV47wUXyTmVRX3csWett4yBO1/pineAVadRFGkDjvx3fyd
HXHv9+4iLOhD5es5qBYZFRpPqVBFHoE4e8RoHHiFVvvdkAHb40y8055UjWmExU6P
evkZ5HJdFknF2oUoZRmseFkJStuX3kKKAaHGrZcY1SBFy3IBkzs3QqP1eNx56aCN
h2UVQiPZIo/KcqXcgIn2dAqmNmmbfO+dSOvxJ3+uZMsAiTplE/ba31HQg9iRXk/R
B0NpId+fS5RLEVyYpS68yA5hAFmLGf/wsKLEcaRMRdUNQO6dbQvpwSPA2ad36kBh
Zo919EvrEPvG7/iuMjmnfGeYWZG4pxsFkaXLcZbuDfik0EC0Qo2NKUhn5V228G0P
O+fa5Vo9QNNKDqjEe1iBjgq6pMMWoey1C7U4+vf6wOF3xdDws6PY4oGQGuhYKiN9
D1froIP6oCcCmr/r7d1fjTbPT0fnl/c9lidbhWkppvJgrgiiypC++UNliOkvftK2
UlG84VxJ3rCQfTXZriNODCM+vngTYMwfQhCdzcw6X9GvTBLebTyI1uiriwGyy59O
7XdNTv+WtGwHnEkcpsX5mZg8I92zYdo8gDETa/pVx4CGbOlYWNMIetRWPsm3vuCT
ZNTU8GOEFMn9Yl7UtPpOqRBfdtmBb+PHcSZJOZvQf98r7UWkwxWh8klm79/7tITf
n4XTM94QsLzgWctVWxGcXNFgxfLbhQdNazTpXNpJvzv75m3y0oUO9P9OFPOfYetL
51H7lVJ4yq/BoLPld/G7m/HFZSkhT6n99UJxVNu7LWqT/JNe4tIy1fBKGCONnmqR
e0OGMv9nXq8n7E8HES/POwObdfofpMB06uK0piuhylTjcXCS0g8qk888d03Q8K9f
BeYuLmy6By3v3JWxMIGHeBMsIwEDPeiUxUY4sratcnkwk5JagR0nrTFZpgRJXf7f
L8RwfkjFKHrFZZTeAbYO+h/XHHGnayXEQCSZU6+TqpmGn8HaSA5dk4bfimGuGfJI
eowSNVjyymBLMyCbAsZM/JuKGzkrXF7VqB8dwBQoEsxdfQ+7mf/ctaK/HCYaDC0A
qHoWH1iy8iq+6GC/e+SfLqrbW2fdVAdRwkrKF8MCmavn3C94gmm3Cyrqq5Y96W1b
nzjjY/+6csqJuNaziOi/i5GkpRyeEgznK/OtH1fjUYBNqMVHD2QY2xsXqe25KbRL
XUA+GetKw+rmMu/vqlcyzeX3Dr/vJNvoN05+FAGjgH1upHlosqjIS+NCSX5IlJv6
ex/ojQpuw+bMBzkOVLZ132yofPxYURWJsKMiacQ7WjjPbeDaSL4kvjAxv4q/jOSQ
4uWnIkpYyb/kSZh9PbxPpPApwf2NrseCrdXHJvLcXy2ucBsQ4te7oy699k0xSteM
x2m6vlXHewJH5zagMefjq3qSpavOREfUy7u6UnONK04W84ufSspeOryXntExbHaE
QTmPBrmJyDxdu7n6+lsW01wOxhaWTm7Y3VvpWQH18oO1U5Sqz9M8d3I/qVFhjwY5
ZuPkArRu9AxOggMmzjxHdUTfJioPsbVIlHKdOE/eP24cOAJirFcFnEmFrPkYF658
6bsH1H7y90AguVqbrCXjUBVr24v1Lp/IFBSpjVTqXIZSpOKaCqVfidbAzynIpjht
y5ZhDped0mjbzUZpS73mFmApMuS9+tlsGNILnBjrdunnqFnR/ZmCJewrSnwgja+l
rnmfLibLEDe6n2mP0T8wz091HUanEUrk4bn8LfuMCPz/tC9aHwHU6Gn6ZKAz29AU
KfXgtGo3k3TQsRaG+zbOgEiAUukoPurzKiiQQ0MRbtGi8drBdrxHHoJ2UIOmoekX
kW4b1DYmFFEaFUX6qIdsEgz4hJD4v0pwXuNoHRUud+dseWhwhsKxra5il8dG/Lp/
tHZGvLQQHJVgl1RAck3IOaeskjuY+AjYhfjOIKGPZIZ3BKmjuzadDmrTbtqOzegs
A0y9Oq2WvHhkw9fYzeWRV7uK9ilg7ncWvTQqhN0POY7Iyf54DqpmktT+yzabq9T5
NWvG+gK6RmTHSKpjAkLmMRVBZXTiWsZZzC5xdHoN18pN0U/znwJ/fALry2NnUlAt
VdpZap8dkKv1xzjGxJqmn2DmnZ4mV6EhZ8OYEhO9eBA2ow6Z5jfSy0dcu8s9LuWP
C2/gPY7QnEnNP6WoIQ9JxLPenrgpoV3Uj/RLFBJhSa4RwinC30P/iJTiNxcNSU2m
KIphGm7hmQpHcvLbpMvPViCBXwHQMBN1LZl7zOn0ULCk/lo/yb7PCCESk0MV+SlB
n/PDg8EHpg4WrXzG4+Lq3A3Zbb1YJD6LfAzrxpdZ65kcF4S/oNcScHoD4TK29EmZ
gGme7H4973+VLp/VrXjvMKSLZ8cF42aiofNpQZRt7WwRj7OODgYap9KGI3izMD7m
lpTykVmfHbMAhFUiSGuE2GHyYJPMcNykyhoZHL6ZvYVqAjr3kRVuhtyuQ53i0URH
qkAz9qJWcr/PTDEVunGXXhnwilmxvF1rOIwCdffZ1URAoTO/2MiLu2ZG3q11cY7p
LIeDmtuD+0BFJkDrburfp54G1DHbE+QKp+Brk0ZdKu45Rxi19VJwqkMMR37XIZw0
B07cz40Fyi212WD0o2+VWzeSPRwQPj504UgHuFQrMeldoksiq36X5j9RJIYWVK6v
K7dj4yO+uuQ5dpZpwXO5aA90n74elemzopmNKdhpJa4G0KTkB7yGzbSn4x1un7Mt
kcpSQ8myBwj1l3hTqPDdFfosfDjYIweEbynhtU/yu8Gnoy7oY63tIa1TSAgl0PZu
CeSWa2OBLGiFwpJDkM9YYrC5Y/NbdC0Hy1/bTp5Ayop0VJtRLlAhjZ8g4rEknWR8
l11uXi1cp2TzZ1yLUAAMPHROkkRcGPIVOJUnbHIpnqGYyT1dYv9KAdw1EPVUrSC0
voU4uftSRzVLthrZ0gRcsVycGuXZEZXKssyJOQjdG477Cw66KuCIdNI6O/iQZxV+
3e+N3NGqI4WvpgjHMEL/pe9N9tTLbQFiIOlrRtKxP+wr78FpUqq+UfA5eXnIg0F5
Eh7gETP1nEmGh9Hmnq8mtFOjyN8Y35VP68DSE0LhpiASPae+WwBp7aACyBptTy3n
4CKZITIDC3I42efXK44CcvBg4TXF6YcScEE/nHH7TsVRZbUswWN2p9a51GCQmIvH
SvZHYoNz0cosBKy9sym27UpD1XkBw+EcF54qYm1NeysrtPoQrlnRg2E8H1Xegdea
DWPd2Aa3jKXqG1Mu+Lf1NuB3kQnswBGJAHiVKiaSMTbeyCHzp5h+Eoxqxm6Xj3bG
OjvBKu5GVCZvIbbO2k5OYe1aSWN0Q3Sx98u9PYSPvqzTgYrPULE7yGdux51ykFl0
+I8YKZWc6udMHu79TklBWus5Gu1W66nzkrRyR5RRW3ZhhCTC3OMhHguYfShPcS4J
6nwNAO245ZgJFb6CKCGx5H4BV1DO6lKI3n3P5x8rIcu/qFhvy3BAxWKw913xpJbJ
8SQFBJayxViSEw2GktzvvIfK1fbsbUlNRmc2HJzjZe+8OFSeey+ptDsCFAow/Fl7
cNZVr1JY18Yn3RUp9L0jATnNqm1WR4ysIXX5plUjB0Zpfey63g0ScnpH53Jm4vu3
FbyrzEI1EnBYJI8MoqAXEyZkb3TGKn9VQCQjOaJH1VgjG/Mp9zJ8E/FTI5+Uvl3t
zJrtkAU35MHm4M63joQuUmWWvxbiUSacqdFYqiD7d+1oEfert2eLp6LYDLrfuODr
IF6++191aYV97jvzrslnQKiCQvhl3PstiFEFb62tayo132UZY2GwxzAZcuWNT5Cj
i3RsDNsY3BsVPwPMMhnoRSTIdETDvL4qPQQ/7886kwD71F/q8jXdZoGOXCQywpGF
+zsW/uTbNX/yis8jkC/CbqCDb6Jd5Jelv9YPFO5MlLsqZ2B65STC8Kmjhm676/kp
dj+ONjrrVae5E9WEwftaauxvn/BlGfYilII5ohOtDd/mpKlZkQjgoFFRzOv12w6+
M0hnCL7W6voXJfNj989KZ5bpATZ/6BcZff3tBuKGqDUu+6YExUk1BPKOn1/TceOW
RSSXsdui7o7n0k37v3JpXRkDz0nj/AIEL3lwdO4Mwuikv9k3ItRHEGgj2ZmMcpAR
GUan0RFcuEIRfn+91VAfRLTVraDLT+VrTypsVm4rxz2jTD6sKfIVhnu7mJPCqb+u
phzZLXDR1nCBM4rEXaRkF0cIfW7CLKXXbeEaFZ72bivcSBJcXOM5eNAAQtcTQzaX
fgsCfU4Xbo6Sgr4NslfThZXbh/xTt+yeEGb34TWdgYVdXZkbapsmYHQ1nFYv8zw2
LKZPERcEY/kVT8SWowDZNMvslc+1Q6NvWPkBAFEpMvKYTmmv/f5AlVlgoItrho/X
GHcQJVSLQPMIdKjXQpJxF8lXWAMjyBiex00Z1012hX7H7QjhN/jC5AESZF2n17bq
zbYVGNdrqGXIe0rCa9434f88CTtY08Rzwr1kHXA52OA9a/SMNo4F+vVPvCXj9NF2
aCTUNk5lCTsvabVmE33H03t/yN5eqo8W/79vZFo2Dk1tc5oO4s96XxDXNLAD0lKz
Q8NdAsNrmFyO2iGlKW8/QzN1CMgWcfSVivvoBUCCwxVnHAB8gQHPS56QT+cM1KEX
YKcm/hgrUQbMYP7TLBaKJvvTV5uVUreCjz3tdM4Q5fUV3DCNEtmPuiT8Ar5HG+eT
L+hkQNsVSgXf2JUp3vIkwDEL9JAey1QTQVugOxaiCOfBqL6VbT3DyQZ4cQqEFq6Z
U93260EzWfImbqm4Nfzw9EXFHfQF1JB97Z6aVyUtVkF1ThG89B0MdjMOLD6eJp5I
XqJjeROhSN7LjIvPYWlkJ+sUdSuapBnPW//PeYww30HdXZD+lsK5l+6QiuhvH/O3
hDIwDNuAIqzIQXY2NHgbff6nqzC8E0Fxcj2dwG0H2seaVYVS2w9Xc1upPs5SZuJs
QCv++e6lZFtUDoldmB0n5eAr3vK40r2KtbxcpD8/RC6QZcKwxWLz5Saagq+2s+45
TGNnJ6c9eK8K4h5QOYx7aVec+uzAuW3NSGvMvEuePt69mPbk0LHl30lCse59cktH
sxaE8hZnK/pNJ1BxT9h2d+/mRBNfZyze2drBVOVouEH02yYvKC33afu0lNpyD1Ui
FWpgUAcz7c9TWOUtkvTpgI+K6LjtlPbJ37ipTiIAfe0dGoXlhxjT9T0sd724N1A8
Zd8bC2dvjzI0XuLYk/kaaR7frsWSkuE/y+JO+DN9VCla4WP1VIiZoBPxPqpAeNXc
B1IFRKd4GsUuMT/gdpycofz67/79zXGs3CAp5uv3KCIy13iOVPYMgmC6+VrtDeKZ
Y9Z5DJvuw6+lTuSLj0d85rhDrKpfPFGH0K9BJ29zxu3KZBD39kMRHwPjVrmx5ZzM
uWH5PBkYBUSmaqQQRNZwX1p7oFJf/A8JExkwtlbunFgSICA7qQdB0lnkRl67Q4DV
D26S6Abb8XiInAsD3PtfFpgivq+WIRoIRfwYhDO7hCr6plKsJo9teSIv9t5bB4In
sZBWuAVhSXv3op8z0dJoRARHNISwo/0RQmmQdhCBSlbuGuG2k9JxuDV3CscUXf+o
LS68GEtFq4VNuv+xWh0p1OmDV6lX7n6jH2VJ+gd5OmrCukRSf/cxIWoe/6Rphumm
dgGcFkvAe+WCudXoSnBmw3U546Mf6tzjP2EwjIgWlWzDjoCbWJQJVNi1XLyZiXK4
2V6RQVHLwZ7N27i5rYiuvQiGNzW7Yi1/nIZMm+6rxTMYDmk1Ny7DTsjsG8zh4UR6
6G4bgVT6IYM0Iuy0a14ZhNamzgUS78NZnzXsoktSaJYxlnYCNkG1AzbVeLhDsa9v
prs+CRF8r6HNn4BhwsVX7BxKkCh89ipOnJHah1g9Zizt3UMVzQP5VVKfQ0WziWXp
O63v6fJF4GzKjT9LsP63x0OSc7sEgflzv22Ig4Oce9dQ2mQph70T31r58wOvRP4+
sp3d901XMnmcUdgGvN/NkLUPwNJnNfBlHRFcVDvpqFmrrtRKJYuqdkt4gXyrb5q9
B/juOLl/ulDAT1FwK0fL9kQvXEuufPL0InTt+zyNfbiyTPUfEr5ztkisUZyQYJYa
qvSyv9QPXQnUrQcAQkO4xX+8+SnWV6zmbczdjSa5K4PxTcwKrdsAal9Bm3VaTbxe
ifxHh9H/GsAVRzzp7UChj/VgmMjvNFBNjdGq1pzP9LNJbPa+YL7U/Pqy7E4VBYBG
B1jZyzov82IKs8xwBQsK8IJHCjISMPDQgkHO00NfmR87ce8RhUs1Q1UvQZUpjCp3
b3PLOTdmGYgdsvQVBr4RRcRCuZznLhv5RCeZJQkfnRJXTt5IV+RqYezfpehVUoyx
+/g4xtTaLrioR8MtUCj9oNy0EuOkWIOF57aA565vZ0AvRZYuV0xOIryDdZjtCDYg
Y5WJIj/exS3InziSfNE9ApifFpBv3hCFagWl1ps/0EBSiGfGwFe867qEQbPEC4K3
h7VN2ZzhpIHXfI/8YTz89ONNLuSPA7SDD+m/+qSSe+LiDwhwkg6l3BCADuldr32J
O85809C47MNuoHWekG8x+4XQyfbsTDtTDqyeGO1RgcYFWPmslv7Ro+DBfX2w5VtZ
hDV0d6YrFqPkkqg0YjmXpCjTEiOQCE365yuR6AhYHQxd1IWD5MlngQGLoqV2W3I6
hvwi9N51SdMP4l0RVfvhQME/WkJlIqXG0+m289LynntnCDA8b3BoGfjiIkE6jw6z
bgQFz6Si/JR7ZH9ek5iaf+Flk0Wk+zchTyJChg+TVMuYa4bKoHizD6kF31fo7++p
ghhUw9VtGc3hpHwS6C1EDAp3/Y6jsc3KJLn6MaLu+DKj23iNbhQnk6q/3MbPyLbC
yAa9Q0EZoV79oF3tdSzXR51MKYzXRZd7HBNuFxh1ptkL3DBKikEbFPJO4kSOat4o
ts8zw/TEbhrLVdimhhSf/tq0ACah9aGEjmaMzAaPZofin2jVplnrPG9gAsRAUujn
aXSbXtoR+wAJeiiprvDyhBJlqI0RsrTqcu5aQWssvAp9ahbodsQf6+Ux93vpxZSu
jdZfbBB+M4NuvbtS9oCZhBuXc9fQYTOo3/3sv+S7Wq0ZACoH+L3uov4HjUMmfQ61
Vm+BTrMRGnEy/KrKl4GYmHne8LeOxzysyhwMNjGbmsXChy2L0/tmfuKaOnCxwiri
WqFBfjpSVamZM1w6KP1KS30Pi7d8YUrW8KwPrme4nWKUoCks5RdKZYZakyVzPZNJ
JN7FMvhmKakEAQB4skZGMtttT90iRY5kGGCFRFRscxhvNdUPr4dAvQ7GwoDZcG6p
3A0knW5CyM5X1k99NrDbylEs+i/80o9RSG+19nnGy1fJMM5rrMD0QjR6M7kC3pdn
1NAAcvgvKSiRzXK9lI55yEEfKx/0xlv5v2gcfwlNF4doGtsSp104a1xQGJoK7oGV
JRW99wtiWmLUS6eVzAST6+0qqv53wXWnfVwliygQKO+WoXTAtvZn3HWyE430+DYO
vgfTAphYP6HL9ABNpGzI+Z8FhYekcW6kN+0hGfuQq8zvTpMwWiUrI7aZRHVgwHz7
rJzB0dEXKJnb0Bf3EWjJyA8CWz8gHH2jBJPTGmroUMUUJdPexEbqyODxEdSMwo3Z
Ei2jMj7oVf1oWnKQaT33LOJKJPf8xkJJQINQyUPhWjVuMaSMRCxdFMVgdl8ENRPv
UAfKu9NAwcNXUXK866XtsQvJ/8VfnmGqJ6i+bqVPxO/EyOxjYssQ6t3AD+FnedOQ
1bj96z8BhtqvDijbJ/IjyuJGZtv9D/9LRRZ7wiNOBJA90Kvd68+oKsefWz1vmAeJ
1/3wtOlUoS3EGfSQcnM6qEouJjr4h+zCkoji3T5kOvyYoTAAf6GsPnxaXwMLFJZr
dyCoRduWElgk/b0AHIKuS3bFd2FlngsEriaodUo3/7gXov9CaMPFZ49er4V5QagG
S2eRFdD9+LrUdeXLPs73J9kFkTKobap5y7OskabEUXOIuaJ/Dtdiw3bZD6vk8k9n
587zMHr9Dexb50XrGmSTgWKFm5h0Fua1f9Z8vECYEGyhzywDDkpAShCd/pNu903k
YCZsV/pCAcuTf1qsWW8WHWyfXqfsaTa6J4Htw7OK+ucQHWHmmmdcpBhGQMU2/5Z7
e25IEN18IRtKpPZjVICH6LNWxXgwYrtLr5l/CPsewl/m0PDbsIVyLUP4kMzrUY4A
rzklqXIuMGtxcWqlW+ZDtj8AoDmv+waG8TWiL3Ebc6wEoA+Kj2kXSAiNIpfZ9Q05
mPllz7FMLko5qwwIyf8mtQ+ZVCOni7/kLbSsP+lsE+/r7RQWBgGYPw7YWhV+t76m
mcWshlVsr5W/Zk7E1vioCJoRAsmebBA6waatKzQZp1mZnEu41YGvrL1j1xFXCjeL
8AM+BmJ6iVdLuiqymbv2T9QsqjXMbKag9k/UB29VGMjoAtMjb+NnSR8OPf+51EH7
vWS06AlxQJxNGQanqGDYkM/4Q6+VVEsT0/m8xwEGUJbtIU3nJ3FhhEWDzMH1oCFp
skm9KCPdpmQXfMezsFiuEbJ2TeqPqC8usEz+dmwjjeVOFLlz6m5UEHx8TOpNyYOm
H2zLbwgXldjNpCERld6YoZvRLT0JOA8dMyFdFa8Lsa0UaFQn3m7XHESra/7Pbfqc
teOUPhQwDULOHO1ePJgKiWEY9/2yVDGGH0vxITLNbbRPS/AxdjXJiuRmd2F+8XTS
Z2WW/Kfvh0jymaiefdbWYX2x/WHAkEFGRaP06B+ar5ICxcX3U/gBL4udX+svVX6n
P1Cvmpy5RsfIV9a8xPey9YlWXU69Wi7q7TMZjE8HVYIeR+P/HWIdYyLdHRu6eZk1
H7fTV8qiPXPOmYAsqJT4+z2lY3/bjhQCuGN/75z8KYnqf8gujAa7GiY6hPEXwvqT
anLhTqdun0iaQjRSMhR1DN88zDD1gnabAFZxMnE/3OghYrmkm6nnLTo1kgLJUzTn
AyodAccCEAy2cLfmGpyRZ4smmn5XVQHmfRd4610wTXaOasUxQf3mQW93Na5CY67R
Dh1S1QNBEySjpQuiX2dRoujD2Ed1luUVrCpavt9WJ42yiQ/aMA3dPvhoou6DaaY0
ukdW9pqs/4kxwGgzZ54dwFY6HJJcOqktE/dQPOikEk67HDU1wB9LtC+ltQU3eEiP
iM28RQqoAVuEf3Ni+Eq6p+H6dNfuTnbzqLIK8Z99Gse7pOd1PCQ9/ZdYqxx2XyIW
Yu/C41iLsN3TwC4QIu3U/v7E1KO4480fCM7z+gAdOm2Jgaqub46biwfukhYu7wln
sCu9R7H7NVWG5sHk8McSNEwuqin8nQ+T7FIytnlz3hZp3fooJ3kRLWHmqHD5JTzD
ORuQswpikBYyHtKOB9O4uZPoHjQ2FxvojTydQNcNKOAt1jXeME1QbOt1UIDlfL19
tkgrY6IOG9coT+PJR3B5kZPoh7qcNbcIsg2QRtMzf1Q5Jdx+VgrGpQqMLX8R8zgO
nj4Qrci/TUk54pw7vBN3vKrqPk+goL2L9h2+vwhxGVcArykqMaxgmgiwyY0Ds8ey
mOPXR4DCbVnrjyICpsMBXvHm67kx4dvM1LnR1pAB24IiJKyaiiSD8Xd6guAltzGs
GBlcmcBorJ07sD8dXmgfXzg2vgKMcXo/jK12F32B0s0F/iUoQ/VWLQpWzGAoShH+
BopB3hnurI1BorV4jBYrFtSaCsne7rPIInXNl0uly9EiGZa2zQrRAM0/D5igkQcR
m3pWFRXhRLZ9+5G4bJIjEXzcxd2lg34G4L+Hwmixbrjvoa3K1gERIdmJMz37yTXc
VJs1DCSHQtqcqBrewIPKZaa8pEfbs6PPYE3C6JcbQV4JbfThT6i+R2uzZFUferCv
BICdZitJVz3izByk2ecnDpMRLDfDVvPG4/zE2q7gKmyIAdQ2eDF1FhJU63e6RWp9
bSlLuk9nOHtciUpHTXvM4UWs+t9ZixU7IhIPu9Ct8bIhIXatFP6N8lj85J6LZGxM
AW/4/HdfxqxcqJLP7qF/hx+qDRq3fAL6qTzQRi/PzFW5GfZn56ZAhRj8q1/4J6l3
tIbj2oH2Djc9ddrj9xgjhMuHUASWrnlNNhB6AXvSoQrk4NWkf0vmT7uQLI5KWUbn
qq3w7aJ6ib37O+f8g7EfOJ3eGYVhE3O3yYjqpU8aoYcZM7Eg5qn/HNwXu8e6YLBM
x00yi9iEaxV1+3AIIUGVbpeXAeVeNCwIH3kbKl2zDZq5Xfv6M69jt/ZJl7axqjTH
MXBaAWXwpqhne3PLh4vyF/johPB01zdSrYsJKq6bgLwYiT5oZo4Lpvp1kn+EsYe5
uvJw5Czo2cWrVivYpOc+PwvBQM6uoNmmbD6umfsnpyIK/h0kxrazxNTRzWeFzTa4
XeepXDstqltW4qwQgcBypOJWJjM8ix2ip6kBWhf8K7CJiRb971Jux4260aEPmfch
RWsMp0UtEmXX4HIh8CWWKg8SpDh1+grmUj8nx8XWCGvaT1LT5NKuB/tYh0KWpD4u
d9m0oR9s0CsdRI42wBCrS7s5iKWhIN0iGx45/QXPwLYvn38Tr85qXZvWO3b6BCVn
OwmdwvqLRfAOdaSBYgkrjMukFItwuUTmESkaAB9RpwliO744hhHbD7BzMBfYq0kE
AOzqzn2OH+H1SjYemWsBQCmEXbF5ecrlBT0/iBdvbvRsqs4ntlisITbaJsXRKeKJ
/3yzT0cAPxlGth9gGOMpE54b2XQPzF4LzIKWTUni31VUwxwC0OxJQ1pLvkvduqGe
WZyAL5Mv/0SxM42oHJrERnUMQWTOboMyPpsgBSbvGZCILOgx9h6RbTTQSNJqd8OW
f3+nY8ZQNKUrnhvqqAsxhW3BFcnhImi931yvcba8tbiVAL3ZaBiBG6tHU1uHuh4n
XkrH0IN7ZxHR0RStE7qnWtXyA9cSVBELAj/bCqBqTzFYVOIzx+D3xDENR1YfhRoV
W1q7N0hrjZqOWMCl2NTKr+H6mhWHetazB1bJI1R0p2PI7QjeNwq82rPIuDoqzWpk
MUQmBymp8zwp0WvySgFPsD3Rq2oOX6Mbfm2y6yQLUgp2DlhcECMFlrcdXN4m2Iw0
UA/xBshGXk20bEC/5dRUwt9NNZgk2AehkXagM/B9c4jkH/uK9UDLz0SfF9xAb01C
VBk/865UO7aeZJ6jy2vR2ZU7aJGCmIq4Jatblv22C5c61Xut3OOwHqQLs5ty0/mz
kazltT7zKv4vrwAmmehy6EWaNRiaTcReol4jxb33QJyqWi0DjqZN2L8VSTYtX2kp
dGithdhaZZnb4JD1M/eIQGSsxNZA4xZXOpHE4jpETaDsJu5CMutCrSWi2yJl5IGu
zIbifEOW30MvVsctdksYgqbGmH3FYMciCu/yrvbfk5OIADJXdrtm7dMo14oW8CpS
Lc9be9Nu3BTAMbfENI5UVcaejqWpuJbxrRFZiqsxEL7JTat5oi0u0aNhUtvQG6yL
W6vRngwQ+Z57P+dbRdyKUYtozdZlfnjU25iAp/xtE2Z8UwI944V+5tCnoLGikp0a
9sW+UBgdT2CXJi26n95w8e9RZCUfU6vtBzjwgAVJ4y7+3RAIayeJKlfPA7K9oKIw
NLbSl1fCOQk1DATto9w2A2SRSsmAeGzcID5gpH9DG/KOCTBKeBfpBVmvyXemFgEd
IDmWjN5KyaWNmoF1oUm6FTtviEHFDQNbyHn5TXajqL33E5S4hKNXH5/6xxkjs7EP
5gk3HRiXmCYzphdhKLUVdAhpqLxBOjlztSt0iUC4aa2czM00MpxfVgkfzSmd5MEt
Pi4FtigtNYBheMJplxwi3PeGhq2yfra5vZ4VW3YigggA4EFjLHe1r/hy/1JjmVYx
bLaVZQnf0LiVq1EbgNl5EwasbJnqJNFqA/39z3VM8zIeQs4CJcDj4lcV5XEb19CB
WcQjDTsRdU84UjoTRvCiM/X5/Yd1xb3oqCfAn6Se8Q22xij0/BlryyYbJHXrjfCC
mGpLfSgMsc1/tYrF8PfsRS/7mNPd/G9O2ECO3jEFk/SP/P2lwgXe+VSw1dH+xyjJ
tHmjPbLWeMT5u02MmOUoUvizS4UTGRhU1xH1gJUsC2dWU2/6AzgyKk/0QiBVGh+6
RR6waEIBzPDOgtpKO72HwEi87qluw5umb5gGlT+mjGObqyP+rVrrEpL9gUL6Y7HC
9w9flWC7hBoIRWMUDIJWf+XI8vDDtchf85UIUV8txq6vckur5V7TTk1ALQU+FkPD
oKy1yBqM+Ynb9Z6rRDwdP7v2Y/Dapf5o77qx3BQEQ4v11wdz6ud7Ek5zFKrB8jgM
JQbJKfyH8+GDJuJGDL5Sc/V7u1nJ+UdT+r1r1MFhIh8xYHonAf4+T/gn8Z4o1gFW
vtIrQM/lYFnSrP1IHBMygzJE19mjlKoarSzXKzbACHaF+BS+LNnWmDY5OQAySQIO
1oqxFDX2QuKQa44f/IigJBxxWjcR/F6euveeh4DDHXAPSc6LWYc5O/OUOe1Im7Rs
vTg9nlzMzuptTLOMyLHXE5k5rdACdkRogh69tw0K1Ig/oMVB00XOivvyvH+HqB58
4PnW3/82R77AKAV5wr+NBL/fIyRWru3Ce4teN+mhLPgHrh/7z25s7UmXEe0CNRQ/
hNZOj3vbr6m7GzR2fWYRhlXB6/hScWeMErC089E0jN4F2cuLM9EiC3IBV2z1Ze6H
f1eMMNZD6JzHUFyw6zOgMAEU7tEnt9005cqgCK6ADQXbqa46e4enChtnZkAT2r3w
Ff0sFnGFGvX1L0FWdWIO32lBZWPyf+WwEhBGSPsk+72QVLr6AL/2HPSmZ4L/x1u2
lD/aRFHEmt8H3cJ3j7wY2D+i643FdD/DDQhCW6wzbdPRoyp4kP9Um83okD4ncBTk
U/N8LFkJunB2GKsAE1p3Njlrf3G/ekO0iAj6za/QQgCj4GCYI/LZclsWeM6f+5oH
mypTJ5jX2eJIWdnc8KrzTjkY7gasEIMysqV1xFRjmbBEmHGn2vIn9HVWD95LH073
FJBhWxWdqRWJMyWoAfKCg/p6l4Ec5KliTxwHtkbYrfFYAVj/Wyp+vT5dyMS4hx1e
Doj+9/IvVKg6smQPLh49zR9xkbCmPhv64Q+8jUHAo22YdqkEpBWA1FgARio9QLBW
rZPH2VcsYmZcXmZyjpbCW/y9VwCO42YQILqKEwcbt6z6zjtotbqe+dy3Fbnz0jgR
Dr4wleKqFZp2AOi4SFeNgLPxnFi3REHHtEX2mAi80vUU2wrsbIaM1r3n120gtd2w
TLKJ0PawRfxP7DE5vT8oyIDgryNRvkCX4zXugl4FKHIaYFEnL1sqpjj4o8pRhaNN
H44JcpbF1qNXgS2OTNuevcOg2uZAT62MCZ16ULLee990Zv5YdKW2iP0EtfMkPs6k
2Dh98fX0garOJHPYt2bz/VaTgEm52m13ZDMxQwTPXgHTgmDZllnXX+m3/H9WCgTp
8b0x3s4kSJl49vyb5wdCVq8Sg5nqfgOpTWsMsRaBNIeuXvpAwe5/Io2v0pSEYevC
iT7pOtPU2w4LekyNI2U9GHwNfJTgFRqDmcvDT33kiwMfuaQ1JVNPaMdFLUe3UZq1
5144YVk4+QAAtDqDVzH7gNifczP6kpC17rbgn0Qf0JUX62xMilJt4T5unk3QlMLS
Xq2Rmo8jL6nr659/ookAHzvqio3z5i8hGa5kMVMlN/dnu2q+V4ReWWt31njL9vJG
4NKkWpGr8Nd5ZuYDkgUTE3Rzd+EpwblN4Fas9W6qde6Nysnv3xx+psHBhp5ZRg/z
YVJ2vnesg146o4tLg0mITdIEXSWF/VSPBazECpTvfdocOzJ7wiYBGbzFku1G5kIC
l5kXeg0BpATcp7/EB3WOSddTpEHOEUBUrwFVAEiJ7ee8Izr/GiMDjgDWDP3KrnD9
BkARxQ4yaO/r5wWRyfqibYdx6VrL0ZFUmD94qa9TbGk7uDR3hUbEC9l/F4YIbjhC
GphYQNHen+wExJZBj6nZEOhJqUgeF+aBgqiNn2oC9svHT2HYMcFRwMK7Hhf3CWDH
yFEr3UD9wAS7IA+/AyfkQLiQ1vZfBOLthhUSekq2hG97FdDi89L73syHi3Au5CKF
nWAkwPytAJWR02ifnOzpXUZ80NenHfocG8dHh5CRAlXVsI3hV59eYuO5Sqtz9hjw
w/c8h0XIPDzWDWLL0rXOTJpeXQ/CFR1iQQehGrF4p57yyt/8ibutGMbWwGrISUux
FfCezV6a0M7BEtz1x7XFtul/O+om66mLWua/OfczgQ1OO9TGSHuN13tSUDmxzMkz
MOwcazxnrox6m5humbZFL+1qUugoF/c6Vsb0nBh0nfjCPM7uebDgO8QvOog4xoJ8
x1k4ML5LgW+b+rTfyXe/lJgbJmGDDab/YspHjDaOOPyBByuxsSXf2RbafmQKp/ua
yQyprJjVzTUcSMcw6SmoDHiaJnfqvaKcONfPyDK6Hn8evtmMQhiYubPrHEw2zhKX
MByc4ZxzSRXGNrCwxuxalrJbHdW1TXqCCOOixcls0WShBxdjGo3YrODA9wnIOjXU
mRULxsTVm1NcNrCg7oAViznw8rmkFYSK7/lvRCN9RFAZCNFkM+Aiq0FCiMWvlHgQ
my7fqDBP528WOhxeJUazbpXw+xMCzxFG4iDuy0G5bvNNZ19hprj2to+lVl2NKQ/B
6U/t+XMGVIB61RKrJG8InHTf7RsUEir5nGwMXSr3treEiv7y9ybbs0iaI7979VeQ
W+8Qjb/p3jjsqfnUzlaNsNUkwRd2+YM6/axlqhRARTTlPxLOWibuuA9os0spFVOW
jE2Zy48BTogC6IVSc9aCgmky2mBIJCj0r2MhUpf6gfzdKpwt0zjleAojvfX4aUJ3
zsuEwJUqIJ9YGw+EyszKxwXqBRFKAg/wIoOmlxqRX8hy/Ey8qLFdQoPNP/FU0EbB
ci+37r//Zh7w8aQLOat2ynp/6ZXL9yRWF9G0EaHbsETPVyl+YNUF3kV7NiulU1O6
F9SHSCl+rApCBPKr04ULF5AQyiGDSHnSBIvr3zsRMPmLMj1UgwSyW7y7Wv3qnzMT
uKQqEj9SreuH+e01KPWb8TPP0Xz3fukpmlMpHqKaOdjVmiZjGZIPM4ssZt0yLR8g
Tv4joTNwoOGsbxdolcBFPzwHxIWaKpcNeHyO7vt4f8nxDoQ69vNrlAoggTgVT6KB
aUH9kWcD4nDTHqi3lmX9Ruwdk8Z32n3Cj+dYGZtEAvDi0qq3aMNwWuqFgvAqqM+3
KfFzOScChKPKZ+Gi1shKQnVCWnNNSar25SAyp7IGtZ3MtiqD5kNBnk3EGvTAJBGF
frvXFGgnl8KHjr4XJaSHh/tUx03Wi5q53kcnjBB19+nHTotCX9bphftEhmlgwWVN
3XM4yY+csA11T6FV3cMqyAZWTDLCdYKCzXcKLc2YE/hFDg3FDOM15464ceQSWG9z
4lXym4IJUPccEIN+31jOnZERCwyMCcBe112kx96SwxYuHu0vX+jnOgvtVCLqke5m
hVWsIjewmUYyZC/npyPMNSBYB7lP9ssotfYLtXg8EAvbkjWBH8W0yF80OvJ13WEY
flZBO7yClltRb1fxckeYSDqFBzbuRf4K4EyRAa9T1JRix86RQIMBp5dBRpLLSM1z
Wc6zZoxLApY9zuUIhMwt7wn6VtbyT6nqjvFHewzTQJn2CiF3xugtmvu79HfM4wve
OlQSEcDfy1/2570JPsWok0jMFwmCZqrBx75u1bN9wHpUIxe1QFKubghzmNnTho6B
BXgDeSce6ijopfyoxTA8gDNH7/y+6Eh09VzGN8SBkcNQ7/ib6K6YxCpkbJ2Rl3vQ
gafi/8eigVtCmp7V+NZ0L5yWxv+8Me1W6Zv707YaDI2MxQ7xZANz6wE7wb8rSyVz
I4lGDT1fZ+C4QGbUYS0DnJ3rS8krdvTM7Pv6hrJvWymGkdxIpIWoFqqtQyFOCzyJ
4LZMAGVXsV37XKqgUsWxk/ZII/as4ZJ1VhlFd4+VL7ddcS6wGXbhOPHtFvwt1+H7
42fP5mIDJLkT9ZWPWTSGRk5LinULes/1XHcZW9eS66XluFp6Q/+JVuhj1sMZys1O
WS+jgnyh0CG7Uo3vzFgRroRolaFZMsEH8bGoz9EH3TywRJMFcva9zr8vxkjB/4bm
PkIQu7CsWn+OV45o5iSGFzdNUy4Rt9fNjDLdKb4fwN2tfIxgjMP1JSziEBEI3GJp
JKK0J7ZUZjurn+BUDM2dDu66gMyUxEk2axYX2dRDJTF2LHgwDqYZHkCyV6a/ETjp
sMh2kGqn+uT3RUfeQzg2tyaJNsYrK5RMrensdLhX4vemXyAJnThKR919FQoqWUtw
sGgYhlq1ehdc4oadxtNrCUBSI96PtSlqmS3/mweThcasdzVus4x76uHQm5Bemkri
oYIsO/vK/N+GPUzYpaHeuyHw+Rf3aKmQsYBvX9dhDxrIoUHkGnp1y6iPZ85csiZV
IA2VUf8IUVCHL/8JyCG7tVNh5sTDiVEKxgAYiCqdPeFz74GdDsyd8Dx5Tew7chm8
VX8bzlAmfK/lXC6OsYuEV7SCdNBiAtej4sZzG7lOsXhvZRhNyABtkHY4HdRYShbq
FzEjgxyVPNyWtesSwa1DOFdrtB6GHk8cIbeWRxjlmzDCrTz5AOVDcnrbR2C+lkch
+kyVmnqIJA6mIMcVjnnTA/vizBU0CM7ozG/7u5Z3IWtt4V/iDa4aNm5pzMX2OjfB
1LOlvjOI0+kPxswhcXoJ/yu/2Ucmq2CUf23j+Wojjxh2HInRkf+3fx2dxKnLJxkf
yL1aKrbok2LVtPiP8alI4nc2kilGs1PIYDOXLycqeF9j3rmpmzsNQUaRvinaWd+u
NLv6H460pdgT1aKuArqfElJps4xitqaGPYidcFfpXVD1d/E05Q5KxgEn7/3L8bxZ
WbWBnk314+4kxkDrq3cjVu67WQjM/ZUsWY9q5Cxd9QEOagq0uD9VmPxWnd1jHHc2
NfnQWLxBymwynBs51uq5jX5YX1Kas5IWO/xk0YfKPigbaurXAlz2bpSYysAaFDWC
G/acCRsgSBawKpkF7J1QnAOGllfAPNWur0ABjf/P3YoHMPxwgNvZYHVGw7iNEb2g
7McOP0B4bD9BuKpHRccXjlacJCm1GGJlIkbo/xePWleWVVMmRWUO4Woy7bVBVl1A
ZLKwCo4eDXmuUIE30o9nea4mnGccKyq4i0S/fuCDLnc+Eh6wrLx8cb3nBSAfIGLe
JD77RLEZoIN9+cNWBvEzbyQ9lBn/kePsX418rbm1SkUIA4m0m1KOzXd+8fJ1TCoe
6ljvQbZVIJdudGpFmjvjmfInm8ZZRIeOQDzZ15gi1T2ncKYHkuQNGwXoPQjSo2cN
WaW4oXc7F1A6H8Cer/r0W7K8/ZTR61l/cbl1g3risUzjHk3uFukyFu6DSUJXW8Sx
kBLqLzHgoK6IOZiQXMut64lmKbpSqbDVC2dLanpTvjqMFc9WYrUhxzGa86IeQjkW
NOhPR3qp2NqFxbvSqFISYOPJCKBcKBHMbyxVt9jAUbwIhT9n7KcGbhX1c8nU6f6r
+g6X+tP6Q1il6YArZlaN31egIa9OigmL7m45KzKZm0qwnxeogGg6VHej8QjA8qyO
+wKyUJEpX0IQLXlpAAsJNLPRDaTBZjkdwHZM6pcFppKoP6kLlNw5DDE+1NH7qGMf
k05E4e/wE/Sh9CwCNjpJUAl2/3Z4Zym+0sOtaT7xYx4rw0Em/PNA/KJlhsLDwkbJ
KIf/7fnTb9wh7HYPLr+wwcJUS1yJBLqkSmSVi5LMz4+C2FBdLZgtxk0VohJc+9IG
SCp+mChy6XqXTWY0Mnf5H8S4YneNwkJE/i0ts+XnTj1XFP7o9Ibp+jLccTIlvbGF
HAgGHlO177iVAfr9MLTp6tlobavfSjynPzB3ABcAyPNTX3SYWmletWnZhwtRy8dc
k6caUhZ3KYjRQ7igDYsnPBuVHoaCncZXfrvwJybLGEoqxD4AuaGTloGyh3UyblsR
SJjV9c9sgk83NHzHbN13LQm6zj/QnOaumYvTRLQC0HpK8Xflo7SfeLbetkq7uSf+
i636qkzzy1nQyXVF9jrMgwRgiQQ9B5f5rA0LnVjvrPXNQ8wseCRMRvVC3qlpm+hG
nogb21GYH3ZhSRXQtg6Xu2IFZUWCxOI+YOY5L3z+8xALTEDYucr4u2pfOQZG+eI+
1MaUuV+LAdgXAEBu0RCzyY6kDXdB/nD1ZdsSwQem3ihZ2ZQCRUm1aG2zoOOT39B0
zlYCMuqXtlcVtLxCz0Uug2Ulj7wB9QNJ9KVsw69LzzLrxWl5jarfgVCI5pyPUo8O
jTGM9VLLRVeSzrdNVjcDOPbPbyl5GC4LLRPqNHzeLqaFdCLTgj3itBdpfG4NbUk6
AS7iEEVPcxKfD/abGASF9VDkY/2Blklnvo5fGiC4gEDnYjqd7T4dP+T9pbUdN2+5
nIYSAAq6EUF1r9cbCxFVh2HMXoPKOIX79Een08j6G+dLBcSGMM652ka09oTo9pE0
WZmUx30OYwg3MZJa/n7/yrwXEC73Lw933zpLYumUzt96y8rwhd4k4/q87d7qg3xQ
bwbdJCY2Vle3faYNSyDXEoP4Vy0kbgKIViy9R8t6B/UNJyQOPDKaALFNXajbHCwb
Xjf1PiGIbpw+egIemYNNA6mYHvk4wOQsSp+XFsCD+5p06+pc81DRmIxNeOhCq70F
AJhE2i787ZLhinKSEFSXs1cYRE74KIqFOXTqr4pcucNzkIDTIeJ7xHm+RtWkcT3Y
A7X+HqZfnNyuwQ133OMDtwvCDqFw1AfsEG+MzV4/NIwnmdu0IdkRBMwVfxWESNCB
rj9z+z1L7+3vdSl9Ogp85Vkg4yiNjo2rpUJ+/Fuzuqqiu/G9wUPA/6U6ll/212Ze
cZXiiYKKJQt5O8PsxNK41uUBf88XzKlKfL7A39feslGs0STsbLzSJNKFUo2zSmTD
LThkiKeQGZykyU32x4mhu5jAwI6nCyQFVhIGlMD041vuZIhE0jB1aebfGKqgV+qC
lJqtHD45Y+fD1Qafj9nNBMjB+fPRPBlIJOZRbcT5iH2y/GaKuajZYzMVUORw78y3
uHGfwgavKhDNV4H60iB0hhNP/4mikA8kE4aG1V/Nt9tHbFrbrE8N7po4/N2/rGTG
1we0f93G38dXhfAOkGLZxAmu+FEO7K70xEcccVscezzKrbBJf1EyZPHZJgJfX+Ws
uY4ihdzlumHFIbN936QiA+9ocvDz9UX2yRZnOCDSLX53r1u3T5WFS+RHQ7U7G0LN
qL6hWCT0CbsJ7ga004T0IMQaJcwgMO3vaMkXiQeV6J9K7YSJxRMy785UTl3+iiEt
nDS8NctzKFrM8fQv15qjqQx8L76rzuBk1OQYLQFmXp+I1iDufOVeZ2cqIUpCGlTL
W6WMqDt+Ih8+g+YzlReQ83hJ7P98C51ltTtkedtQ2eoxRz2qY4ShhX5UpYftbVfU
qBrhLGynWW8lz73XZ3CndDWKeIj18NsdvC+Kdgk9vgdKv7IB3K/YUfbtN0j0GQTA
ySOYeE9tKhbNknowzqsbARtFjNAqFBe/QgR+kwA9Ssh2xb2gVtNguMk6PrOqPuNn
aieRSgNPqnruyAdF4w40Xf+rpothxd+QE5b/UmUFwMraemF/wQUyPEs9StVEEDJe
`pragma protect end_protected
