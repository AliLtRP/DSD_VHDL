// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:25 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WsCkGbNrtnmGs+ZFPj0r2m+mtpFf2nfqA/L/7och6vEf/8x0YLRsMLtngAxnoKvm
MPBos6QqOLKxM3lACA+9ZGKICjKgAXrJBIaSP09003Y3gBPhbpobtTVdp8Z/rI53
tXlASKZ2Hp8anbhpXZ/ItiN/UAzoXH/vXzoBIAtHcHY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10624)
6nLEktAZVnpXUdD8275TadCU/rYxREpHQTVKay5tTD6IJx1VMqbvtEzUNwgg6KYr
L1gXwRJIqAT+QgkO3rn+k03JGav3d5/9pkbizoI/eem1FhldWzk8JX91z0j9NkG9
P3NTSnhKWOoGj2lGeeZuH3dvkE/8GMf3zBY+WVeso6P+7VclNnApWzCdfPmopSpK
cLxICp1PJ4UWWr25Luh2IvweJY+ya9ogNsHEQO81hK0aMN81Vb15svzuYIx02XTh
7COiFMxX0MkgRo/x3IqaGfaKab7GLsN1FcQnQJMs1Xz+E2iBZ/y24Ofu0oEv+w1l
tlPhsz7fuJDXSqrrKthECoRjnGRVYJ/iWaE+2M/RucCMLgTIJubiYK+sC+vtDfyW
+B1X/zsrKeNgACQuRbLdFoOR8or0/Q73vZ/uDkxCTSpR7Xie22sEAJYVdyFab18R
+oAPlpGJ6/jLxn1CSZaTHDnrk+f5fMe8Ssfnxpr8LymHPldvhdEeDPQKA57hga+b
uK3MNuhtpRtDeBBj0s/940hc71xpD/h3wyWDNHEDfvMSAVkdc4CXPhVbXCqCRZ/+
BavsZlsYCeOh9+y6XHgpe25ZcLD/L+aot2Jurdb2N7Znt0A7JuxfI+6LX6nuhiI5
PeRu3FCb6CjcaaLq9/+DhOVDADKSGNYXQsQEnUw24YGvymLGvxACvnZpRHmUDymT
eWluUhHq4H9A+a/bOa0Z09ooouDitVXNhYAbIMpeDims5GV+pllOZ3uh70exYWw9
qtG4ZnJ5SZSW7z7Y0Jx4J0hzGOA1GvmQbEYW0ttLcuGWi0A34gtTuSYU92HL9H8x
WDTXxbvQlBTHQ3uKBl4yaCc1XQvI5qT1Wt6nh/LwgINSM6+OTaxCoy3lbFb95fh7
4q5CpNp1vLu7gGICGfbRs7ZzeiT+NMSvSBjftd35ejyBG5LQke6/1Dnz7tqAQA5A
+kxWbEPa6ApXr5k2Xl5k0qJ+dHCJV7QSMKgsDv8wAaHGzH7btKsEii97gCql2OyS
ojR1b0BisyCMIickvYRa/b0DPpa8YLkATi+zwQp/JYgOwvhB2EULThQ7ccXC3iSe
bbWYlqiunkr+1SYRfAZg94TTUGoAnzhgNiEjjGNZQeqtFDqD554L7uspR/+Y3G/g
leKkuINdQGfgRe+9iGWeYWfrpmfhd4wCZvjV6cXAVRGtpLjlvewMbH5AipjtOypd
VLvatjuESoO7BVq0rp4q52AzBxsP5Q4hYl7dp6IwHF8c07HOQjr2pgmqhmS8Gnwa
p1UOoZ+b/Gd4EisjFho1hd880/YEXbVrhp1R1TDjsIO3XdsMgHwuneb+UeCm5g0o
5g9i9Efy7fTg67kAHtSSrPjaZxai5RN3HZyoaGSsM2VxGRL8vZt8ksQl2Octyvxl
VgK4obxgbrohUGneJAv9uaAdMaR5a37Tq9gVZvh8wLNJ59pHT5d1Yyj1R2Cjv8eA
ttI7JbwqV2+nftABR1Rack3FOe0XcOVjRBRUBkxgpAAPYNwnTOovgoPkGyownhLh
LsLyeQAJIWrsO95xcWKY6J7ghv9VT0cuHSG+2xXAAsnZyqhBGDY7vLXLA7upf9dG
FnE5IjtsEL0hDUqpl4HrdBq/QL875gslbsKUpu066dxwY1k6Kymq6guI7zOXniDc
wnuDpP8vmrYmE/vj0d5xGc35+swRZwdYzSoAtf6OF4i6def/d7q/iTLNPw165NCi
56Lprj/z0WjVAXwoCnYHnD0lXDXH6rdbwE1ICvUSu6x/kdXsl5eZcX75oOMVDtHI
xl4d9QsEAb5shSWKwMvLcqBBwf5DGbtpNZitkbbg6JvAJpYN8aTNnDxNYLfIfi7V
jZ64oxhXCfxYxYceU6qUEyMNM0k5Rp80HwI1m1KIw3AI84XdkIkCbDd0kZ5EZXYG
TF2UheC1jhkYkZWArdsb9XlI7L8nLVqrm/jLQuzsxXVr4psA4wDXUu8vP3/HpJVt
ZgA5COkF3VKsxOuNnQkFTe2Ec2fQy0SZAQGGStBqgkktk+eiwpGl1x7jNJcy23/W
tL8OKo6CC3IWUiRZ2tDqKjLM2zLWWnqrj36UHWsddyGDbEnUefRIgI8sFHVCRUL0
kTNqNSZwGaBf5gYNb7OVQ9CEhIAys/oxD/L4RIN/cofVBGXyJGhGC1E7BgPYEFoB
Tac2dzGBe3XD5aQ+SgsA/PZ9k2CFTa98WYL7FbePdbIru7XN+XndKiaVu0V/41wQ
kRfipP7mrKU6EHhYHV4to+Y962YbC/Ml+hGH4wnIshEAw0uMg6+Z/Yqj4AWw4rtd
3AV1NGDF54PU938F3jwQ1D82X33i3bC5x6LpLXvDemX2wqvYIkRqzfLGnjVZ4YrK
8IGaEO+qlzXF0/bKlQvXYD3+p+O4aG1rmq3EYUyDH1KXXDcgTu681Bi6j2ulWvms
Uy6jqRsvFwSNAOwyaEzEkIbiveXLKwmGpw1t3OcibPC0J53/b7eiUFk2NU96FTMM
9co9k2i+oUl6zMjaXitreo6w/Jj/TePF0BkMcNtkwRSqnXzccy59IIlJS/JrxyuV
7yK8Bd/ZepdBUFxErlgf6sgFj1FJU0vof0tHqDohMFXibecNCbx3KiLoH0IpHjkX
ZKW9qPIKc8pqP3uIoYAstOIJ1DzYNtUrLg24Q/CGXyP+ntud5gSJgRv2ZiPKeaMw
plhHehoXpcJDtPR6wAukvCBM0GkvBDSfUOACQvq44CG/inj03Nmec4OPITmfOa9B
olDvk2mDE6wq/3CiALpUoG0iU7DjSRZ1vccWTBf9/vaXMfizilKv4DgXP/VomKIZ
PffnWJvVpIoee0KvTtW9ikPYam5teCUkSryfnufGElaa94P0f/Sg2SNp+tv15hYA
UUc84Y6OUwEuCSDCO5laSmJ6NAked3VAG2XGJYRL185CWtjf1SrEgmwBoilmEFAg
hctvXbz412o6DdDqm74wjyikn8DgLG8BzvFDUTfNUPOja+e0vbp0vvQOk2TIKE8l
mXhGfUdii9uKy7WjNhKEnFGy1gnG3EYv3VFfPqqJnJVKPzhZQoZNpILuF1ZASNfU
SG0nzG1x5La2hwkCQ2PBtwzd0E5nsvNwZ//bvzAyK7yMxhdg4wFHVD2X/bxCShhf
qghJyoExWLUArq2RzDkOxwR8by/N24CU9HbbkhGClob33h1LbZ1ozfaYF98CbJpS
Z2O+pz/i3ZCxTCKj9RFWFEpC7qsByy9P+ir7ZZwSuSxDKfJjf3z0y90GtB220NYz
fX2D98Ppn5Pu+ojSqi1/slWYlMdgVt9dU3Q4xQiKpd7p1gM0v6mUmZkSnmtgZ6Ma
jh5tsmkaRElahMqIubFoMU4shwFGMvyV7cw2O3a5g60/fHkZz2/dVOyy4C8e6tQs
ILOMGqp7163MAzj4WEDB20U0HDXiRFZB5Y9wE7UhsDU4jpO0UorF8SZ0CDcKOH9F
VuFqNiVqFXiGg4TaWiAkLOf/s1M2snhyO7L4/P3ezqYZVgTAMkFe4/FXKRAlY9c4
VuJN8pIkecvX42RxJ7yOMTpNchDdQjeqJxztNXdH/GUfYSgepOhvryXvHUNbIkc1
IYAEbjrmj3Y6hdiUi2N9dPYcl6jsKbrEvRofhrE6db6NXQdnGbD9Joc3k+jmval4
Wr2W6dfsjGILM17rK7dE2NNjIlpWUOoqFAGc4VGEwAnuCLNvR1RfXS5SM6tcpOSa
oOcR4l3nGLZ10Kd7AUuCcan6+oZ0OW412zLg3tERDJpLI+4iAWkG8KhJUtb3vIEP
wI1Q8nTUztBxxv97ezzVSn2BudTGOSLgxlUurqLABg8AS+M5u0Fjoi8newegBMaO
7UT9xCyy87HWKWDsP/Cz/4HqfPHP5GIysmoucyTf6dh9Yj5eLZCDlMMVB1FPL30t
HgG4feRfKqN+w+kPDgTBOO61bWOBB3ozDE68vM4HZt52DoGHsZl5hGOwJONYBVkQ
rxbb9/EB0MIy0m+6pbp+V+4Il2nNajjQsEl3gWNKXq/b2NxGNPcitx9TQtSAiEwe
n1TczmA/cEAQaOEZpM3SSoWdf5LUs/f7ENQuR6nkY/9jKjMdVlBqvMUilM7hYLkG
kDG0Pf/LMu3CHo/8m0pnmtxVSGXo6dzXiTXDW/DtoQw9vj4vZM9pvLTqvhZ/YeYI
ob+tT5PBoThk2imeMgTHeFtVvN6UXlVrfEUMt6c0w+fcojXgEaDf303wtovg1eAq
MubVeiCxjOpbGa4+zRx5uvtFJU2P0Aknhv5B5OXeKF7azCvXa70/QA4gddGmViuA
D35O84Z6I7urUjrmPx3rqyFjEVYG1fro0IoTQKvkCJXxeoG5lOjo9NeGSqRZPsYb
681MBCnaAgeKxI2KeU7eM06MWwcuWhgnRSsnFgMzwj3H0vEyfUC6l2bOpc2fScE5
cfPBGam4nnS/5bIP4guKwRN0yGGXJS12ciGq9ycdw8QO9xaQ+WVFPeci0+sS2vA7
rIkbflFrUU6JzBWds/OSZ8HX6sCl4xsYvkUvBXetwCfXopdLtYKYtS9BLR6FQ8HX
r6vHqPCq/Rs0XV4UAiDQ+OwHZSE2xb8MN+hSAnH+q0N1gXN0pOwSwcFXoEdzU8/A
61mmpJVC8DU2Fhhzt46KxmAe/WMCTjMmPHEsLuT3B0r+IaoV0bAmBA+h9Anl+KdN
KCYJxpP/riuvAKcPflitHTa0TtAxeERXrmTNHgapWRpL7c0f7zBwFLMYZSf1h1le
y4VhcOxLUZTUdttrrA3Ph194YE/6/z1jCu6xA44cC/so2tcGj9BWnhAjoWb+PoZl
T9EJRdt6ITv5aS7x9YtnFeBJ+qVcuQYRsT8Ynvwi0ry1GNgYgypWeXWnvAV9+N97
ukh/U7Vme9PtJJl2hAVCzlfS7bReLFQDc28/+AbbQWYqk7tZRQ90Az2UELaPShBx
UwzTDkcGtjUe92EjuXmljhrw6IjjsRH3Y7xtx+XLztCfSJcSE7CNDhryO77mkxZt
kmipTIJxl7EZ7IJJBW3+7CDgOlBhDas92/+qVWJrmUQ8qyRMWQEJotqUJbCDUFf6
rJ6Sc0Whm4wcqD8i6buIIkXdRS8uf4PwTQkbsF/qfw646IzL/5DxACzL51zeQSJb
rAJY3/teR6K5vFYEsoAjV2RwLvd79xF/irBWtEIFqPExtHNT7MqBiHmOFe9vzeyb
Zj5VYWAFB3kvG6s0wDxhoCgE/EqDks/RCAHBzYStlIyzI2fmN2nnFfdFf2Di/Fb9
9D9P7tizlIk4bOi5ootkiTAcCHuv8klUdDy5zZpHoLTka4PgrsAGwNXqpDlhPGA/
A6HuJ442cdPtAtY7QNm4uQAfU82goNvx7EGjqEvOLfzdRjEexsg/+L+i2y7Ww0wF
XeBRJnBzAWit8dDQohE7icIPPFFk39u9g30c5+h23zTmpmnOPOVVqrqSYldFuT1k
Jwi5QW1dMfLumnjDrGyKEXozM0BFq5WpDokeQwi7fMlmmDFDC29ccony3oFzAV5M
tPle7W/ztCkf6dL7IITcQWvoqZHMeQiRrQd2pxKEN4eXeTQLQdWbzgkjOIKhHtm7
xgLH5HzGimRFgAnwZrc+/wg/7N7LHL6N8nWz+L4IbAtlKmz4Y4YCh4NqLZvOhotL
EvkWvSbub8AeBGBUe27Dpyg+bOsXNKd1oATvQ4ZBIBGtj5EU5mM4Q1rlbEt1VORR
6yXhg/UdgH6r+NeF8n+EzCCIwiimgrUvcvFT95JJ/7AA/KP/0QpxiKURW4nYdpeZ
1kCumEptpnmwgqtMLI+VQe2Ngf1bpAP17cWNWOI/U9XpjbQhh7IhTR27RFZe7uEO
drFwyn+KXXtLwxU4JcycGBNtfnyaueXZlr1H52CbHSAGc8DsD/SCzaQryYHX2QXP
eMriYYS47tpcTsdxGBNBkHuBl/xb7QQ5deevKRdjFCXII+X83jVh2iE/dIYuFuQQ
TJljZwAnniQUGKqzGqWOhm4GL2373EvHPAsUuW9mSGg0/PdKdpPLF+t0N0ILeJ7c
ePa51hTMQds//mthHUR26yxzM23HeiQak2gBFbtJjxvv47IFWaK45u3PgP+X96wk
hQMibIuvSjDBV9x33yCE6u4XHLm4/ZEsTJWJQ2Rx4Vjf5pm2zwzn/LtxcNuZriWZ
xqLZM42DP+reVo4EnTVV7Mx5Lhx4OrAcskv2NfLVUW8uk9BeaYsU6nmZXrCL25WU
ukbbIiGDOLpS1sfQyLyonXJLRhlLuAvB3wDvQyg8XkNVeAFGjcjC22VrLuAZjdS+
24RThiJqiAdc+BQU2Yga17Viu6bDkpBTKLO9mUo8AzP0lCJPSz7jzxTKfbALA5Ck
Xp7ugJ+5hEmt0j+ZBCfw3LcOmPCUqWUmPD0qiAi2H8UDHwuO+ql1KXK8X0wxqZaB
zJtXQd7CWliv+HUvivZtE2qBc7goRuOp3XljUA7E5sfoyi2So/n93GP/d08atON9
emPr5hs3nDduFXoCN++r+BS87wtj42eLfTho8ZFiOw5vY2aY4GkUXpJO+16VuV/Q
qhazBOOe7LOFpiG04ip2bG4LQfUcnaY6b2CX5UBsEcEBuLO9PorzwJ2/uzkpp19K
LsdbmKO8/tSfUaUFnidUUMWC6wNLIrzw8HsVcxRa3MecfoHdEj3ilfCivnYx0u6V
dbLa0YGq9lfy3zySPfYA9QeUTso9ED32EHtW217PIlTPW7uaBQUYW8v/oIlOQCFE
sHB8wC9O1CXcFAuAZunWwHZtZPIakfbp/D2hKt7AtCZ+rixUv0LJXqpznMphfEwy
5iz33ZZL/p9YJ4ashkpWlwZLw4I3FzC1TMN5M2QDmvKakYsupAxUPplO4JwBS/ZP
+YMuj64Uv/LM3dEey4DtLN26mhq3ChPRWellz3fxlpg+Hk4VoU7PTKG68ZkHvXM1
/Ojg2GVYaZyrgGKTcBwF0HU0Jz8ZAHcdG9nJ15cfAex3fwyVNajb3906bPzfE1rM
wL+XngL+iCryJKFNTP5XeTtbXBXM/bwTL42MNuXvDB2hPk54XQ5BJIhKvuBn6EYT
rE1c5tp2MUgE5PPdCnDp++DOSAmz71raY8VJNxD51049fGhBQDSy9ZB/kYeCFhk9
4eBAsdBF023O3wFdSZmWpVSunsCghLI5PoZIumvf+WwAZwf5Zdqy1UCC6f/9X/D4
MfMIWNolvBVNZ1o9SuYjP/sIvdWclGonXeX78i5BlFE817wf0iTR3DF5fJNXoAxN
httYKChOP1UDrbL4lZYjLi11R8X1097uHz2W/fBjK7Ro5/o/nwiSODp72R5h9ZcJ
XLMtWvljHYJx2IYlY1gOOqzXFMHI4UUsgtF3MIokFhuoOvVR2xuC3QuJFW3pXd0B
yYkNo5xFxNIrsja9D46pQh9zMe9swKS/+exSxQe4dHio6TdsgGwyFNisRQ5cqFFW
4L9MHHQqQWWMs5DqvBiEScNfV+X4n9sX1VxAjcMdvyrmNrsD4rQbcZnZkopIJ3Sx
0eQP+6M8cTvmin0u6Wb4PMS+v9CkWYON+5lAz1mfwisMgA8BJuvtPWKzFWGVTzgb
h66p4KdI4INsW8TPcwZX35YS4C1uS1RoIrq7snlZ1bVBs3nYGI6awnD23yWVpfDH
LlqoytKiN5FvJnej3NR0JtYatOIBiUjV/9cgLZszVK1lZE6mrLXuhyzHJoZpdixp
ta+oShDi7igMTTXI4O4tEkv5mMst/r8WAB0JYBi8vdTuofyDsZpu/ClqJClNfzKl
1PULWbeDVB6BRO4w9YdGmXztQiMtr9ADNgkD+l72zRLjH5hr7ALszXTI7d6zZhWK
+WW+ssoSXkyFfjHQWohXcntLfiWllZjcA+H1P52Bupiims6WQ7FZdsOrdkCznNFw
THBkh3GnbIjd4oYJHK4womomJ6L2H/5Syk/XyxfEM1B7GR3+hZtsoR+2N/Nzaugy
yKrzobpOQteXGdKTfkeBQrH2ezU5B4e7v3kbbg6xCR/uH7mEjGT0IJy2+n+pRg9m
RBN6zNcioqmgZM5LmMbtfw9VvgtxiucTRiD3ZwBIWZU4q+dXx8m+Yd7MnXBqNMyV
3VU/ePV1d4ywrBsg7XusFWMAcNwKlMEEpS51NY6L4xCXK2759giJL4Zw01EGNhHH
TQtniHfnR1BO98VgCVFnlzHxlVkV1zM7jIz23411Hh+MuadzksHxEvVK5zvFF8CT
0VYaWDdxaHLzRHB8IDjU6yxx6GicRMuajt+xddpb7XaE5yAi3sUK+b6EVVHzRviu
WEMtm1rq9KQ10OfllGO1q8PAy2bgjtPLc5wseTbZ/SuFOeicDAtIqsY31lYaRVSE
RMyp4MNd1/1BagHzZ3WhyAnFF93P7fJ81wOKOf4JmcNhaS3sPlg+zF5bDXgksGno
m2wiuvvAfb2sR8sIJq4KS4p2OURrRxHCpizUoEdyk3pvdf678i/Cfu3Fw8/5YDW4
e/Pkytfdzk3ohEit+ecW1nIguZJ0jnFY5vt1PBqQ/NtEJfQZUcZy1UtfXQYQ3rMH
VUEGhhHDYxJVmbSJTwrvhAgwbtYrxj2+Kax/oVLIfwVCCbVH+Fk6v4SJRw3342XX
7fLNjTr+c6TqLaC7glNxJnaPa+jWJsUBSbcWv1ttUUtC4aN0x6fEtVEBChAFRby/
Od7SBDxES8f8gD/5SDb6dNQQj5aPwWPmyh9Rr59i7XphC81NBcqCUVkSpya88v6o
enxzZuEqisE/YLAQhViq3etFpMJkSne6VDHY2bVuA6eLlEm9JSmRdK8lVndNUh2g
jwk6tDlcbtb4DKNdvhCzMz78SALc0t/A6UYEnJJ/bhM47O1XH+owhfn2NEBGcscO
QZz6X7yn698N3spM6uVFPngC4DMbnYb8zogm+dFYFtRHqDmWJBnyO6D0L83rqQ/W
020ZRt/1YSWZDFIhWC3cd7BdoXm/y6/NYfMsYP7pVbm5jl2CBKkeRWFst/pUgr7k
VUJms3kCeUmF9Xi/73pUbQe1zzOxAhbuSqBh9r/87JX6KZu0zrd7KplkZHhBvlVs
3Ii5aLo8ukHIXmycPrdyDBlbCgyu0sw5JteutrKy/SlGAqTJBH8pd6ti4ZUOdDxm
ZCmNt0n8k3P39Hp+e+VCaeOWZYXBuaF/Y1WCDYMQLSaIeWNjuZIUT7tiXc1wCRbj
ZxDpruOVKKA86w47Ko9lRjSn4lfp1RU3u+lo7nErtm1PEl+ktAQ3ZuhfhjQu3YAk
hcsnRK/+09sXl4y/NfjkDegsobqGWWUlei90hPdruoWRc2yzcog+nnq1Dx6SBZDg
aUlk56LfoF+Iw6K8bXaSl2OmIajsl3X/B0/tZBniO4H18GkV1ixphctPMmBFBDdR
hvzrM/0FG/mEqsIUJEB2f00tSZ7rfJOFW6eEIZzsmHylmeNNrGq59xaNbATGbxjt
hTb5MwyDEZ0k1WJRO3U3mrMsal3IW03+pmv+u0eT2zA1WRd75hZr0EyFwensFjKl
M6iOGfKs0BDkPGt9Cqaf0xQeVL9FlaHLxlhOXSszyaOlnwzBnZGGrkm3ZWc6PEMP
tZlqjayeWoN46LnwclFhD96lrR8HyxA6y6Ux1/CFAW8ZnrJGCDM47ojBQ74712JP
bHyrTETnyFptBfUVihE0dRXY081rNml3XZDJkq53HitUOW+VlhBKr3UREeqFIcx4
4HiwDd+AWmWbTbWL4Mut0mPEaeNk/q+OjU8ZL1uG19yjsXe59wTYmtrv8b+z/f+B
WchJkMVj090RDTk+Nc5H72Lq8ntPrMUSxgxObVTucNMD0/ARbDxIgImyfQkNwu4h
SrXQTELe7/MTky2DSpIA5b9fJBRs+XZqOtQ0pboe15cW+7A0EOuKryk2hIbzTtMr
C8H1/t72NtTx0k2pcsdhpn+I1oUdyQtKvaWu9+4jtP7m6aM43K9071DtSElwIiiT
34z8fMs+1PElU6xtdDcvLmV5qiw6GV/jyaTN2vgzatkFJLSzTLplAKajpnNSrLGF
i+THT55Z42wSPOuZ4wXDLjjo5vmquc+DqG9U38wD504cfieMs7lH94R0X3cEcS/I
JB1BsAIG0B9I2gMGGEDQqZvqnFzC0q8ofwTHJhcUD3oIuX14uN45/SGnMbcJ8f7B
oPKJXKQvQUhzlbfIHvlC4PxJpRV4v+rzTaZ2TEUNnqCdpX5X6s8dSgaZ0qFp7mV3
b7PGtKkYG+k5NDiTd1cTSbyRq9kMudYaxOry0vzg3tRyZLowhvdENIsstKNaCbD9
t3cjXcYrmKCbaTXRt1QWxT4+2fn7kA50/86nupVskRhQ2pxbLMhxvOSerkfUe5om
dkYW2y63RpRwRNmHEtGPpq8g13tuqsqzp3U8Oy+UXVG+QgKCS7MvuIe9qLAr83tQ
AsK1jLX7T+zXs/ZyHWQidadOBKu+xWEpz7ShLOU267qq6bGLJgLOUEq6S2lNoppP
FMWg3Vb6xAdVGsHepufvGFBXkLUPmCH45r2sY/wv3DfhE5fnt9qQgHuveXsNc0pu
GepmLMyef52zAYWOG/h5KlDYHnhAZ8PfdR9XyVS9ByFoqPklsefG2q2dkxlS54Mj
y0EYZ5D0K8RlbBkWf9y1iyjVhIybEs+SyuX97iAFXyY2VmyoOWgy4SVp1EpXUBHD
QCEAgypzOMvYYtTUL5LroFM3YQpIBQ8LI5640cscowmvXLJfBZiHbNvUMYlBhnhk
/cYXn1NH5QYuT9ksOw7KfQnLA1yFw4PPVNxOYMp0bmmmV2B0apFdfLsArvR3CYOi
XW8vzy1584dWQc/M1U/TRyx5VArfWCkIwB60R1BLFaXo28SNgMkwXW7q0DJ0OmdM
C4bnR2PdsZQr/XAb6X/V1+XGCCXKzwaBDLFnQsCYOQEBaURcG4+Qy/idxuqBGGCN
cW+jm7OsXof8ZpsQFVmklzzuLBgnczNlrfrBzIx/bClJE+wXhcZPSVB1yePJfgu/
Xrw97QJm6C8LCZIKAplqvQ5cuAOhufan/JMu+5TrR3lIPYk0/YCuoeqWFa0dsfXy
ivHDgBVFk+xQGcQGL0plwGgqqzhGuif6Gg3xFtkquvSbzO76HRmK5j/7/JMsVcaa
TWhgVeSr+vzzMOtTJGW1zxqz77ADXCeXxJwX8Q8ANI2kfE2QYHReONWmFW0auC8e
vOjZPYYy7RbyZxuhNXIwPL6ujRCnfKz3J7sxSEqZCJ6+i8iR01EJeLO3jrF8gPZZ
ocjkfnVeMWq1++0y63j0s01cNSPsmXHJBC1nap++bLPV4xkkE89sP4YG18HmoLRP
e+Kjqm1tl/ix6hLqQ+W9haMSstKRD9R9/hB8f1S8n46kDMwhxzuwAuXfEtCG5/Fl
MDA1sXYv0gJ0f1I222z3TwKzaMnyItAH9Ra1NchzB/FTaZBIHsW2UxeaV9Jd/bE8
0+md4dhdBdsgo8i3O0tiwROuLT6F06GpGvHK7s8joVzadkTAqTV+9KbI3c4slGIj
GG/KkP4B+sq3MjZpxyUTUnaQnAXmM+z+lEDrNRq7VxdFZQ17dePCOchv0VuIbnuM
K7h8zYqOM6NdK6OdUeHWlq7nXt0yyDc1JzIsdJU/tMlD+mIvWT3r1AdTIQ7N4z5z
FINrE5I+DIx7T6tj/ulfUNyjo5jsib4Nq+zmqmFsFiSark38WlT84BfRfxu4oL3N
0ya1S2cYjfF0rDOgXn/v3aOWhc9IYZpwaPOKCMG8wXm6JwKS1Wr8hLRYBVTI3gAk
hXnVWLb4uR3vqGITDGrduWVJNJxsp7Bk+cPEesunadIAOqgNJY0zlHp0Hyimip7K
mTxTxD3SduIK2C2Gxco0qRPRCf22V2JkVR9u1Tt7hPh7ogQOIkSNHQ9za57tAFrx
T0iQ/pk9mtvMlMNpQtpg2H3Tc7vpZYUhC7mSAx1QiD4WJAQYGWtMxlCqva9oiFAq
5oJxRxssUjMoiShm4gTyxKR5GwYn49K/7/4wl6ohddzI8kpzeMlUr+1/bXUObr3G
3Eay8rUW0Juq/U+dllHmR3kvTMxjw7HhC5FyLQjnELosMnb9aFEMczqSZJRi1nK7
yPWQG1HXqBSwgjBAZiiO14DWp8hVhbW6YYMlbLLOzXagzILN5fLpSmIRLgTf391Y
gqIXaNY2YybDghGrURFuA9IjBpaDK5J7b5HJsIB2FswoP5qzb20pVqkn/mom9NfW
gKDzLqMX3GzcH8GLrjwGk6aceSZduDtN41DP22iPkWpokuY36zvWUURedPjuugEL
fHnpEAzrOS59oj35pJOb3Iy33n7WFhR7HsXfCb4TBWGriWE3B2lsxPdN6MHxbuFX
UqEobNEDj9PEyx2DDQUnC1EVN9KBGE0dqW6L5olYcbb34B+tRbfa3C1iQT6jMuxD
TsNgN+HMkQXufSNZpDZk/E0PGqM2sRBnTeIhtVf2AxESyYXJbIZzgmA59zS9Mbav
xHr70Rs7UieXKXsgnDpoAlwqUvq+nIrhP8hpLIB15aETQi/c8nQZzku5kS765TF+
Fimn9TKW2KaNnpVg0KoW+vMIQb0SDtb6v7YzOxuDQqTSSZDEL0qnukAzka/YRW4A
gXCtQBN69C+yNv34Fia0qer3u1ZYQOXa1J/x6c7XUYvH5Y/AhAQObvz70sUIOT3p
ApIu0V6Fx8MQc/fxYfHyrup4SamBlzbzvulOP8vUedeEzmCiBGRTYv2H4rfMG049
7JRRETTabIctIfJGlyEkc4vb2gt51NKeqYdOuW8rNRqDjbPcOjTJ5oqE8QvST/fS
GvsjE/YD9aYzF/1SW0/HT4CYXAwzbA2PWTlA/G72WYDvWqhf1DJGZj/QmywJcnWh
KBfhim2+Iq1DSwk/GH+vbbsuK5NmAHqj19Im7wEln/LjueENuQ2DYeSvPdOBCYAo
xpHL68F1pA8KMCCkDxRGCuSpr8pzRVLLT8q9ssZ9Vf/yBKPprzIUNtAHX1fXRWKQ
QZsXkDp/txobTke55diMOuWbeMLG659hU/IPILlWMEAQY4jiGhiw05uhd+3UGLlw
MiQ/Ff+t1HBPbkrjB1AICuXCnUQvFGL48lh7zPtVjzinHKDn6yqLfx4UGHDVBQV6
va+9cv8tz6XWIQAGwHRkk+KEtRoox7QeBics1vTC1EgPJ+bcMaY+KHWatfLQNJLx
fAhHi/WnudLUPCrPpciABhHwXCkCW8tN9+1zgtEUSlQlBDOfFfAErpVqkljdKIuK
BnojeHQM/pywsECCfOIT/ZbUuyPgMWtubMSiyQEZFdIvaL15CO9BOUS7/wLiQ3uA
PF9qhI7xfIl8N2Xk6RCaUki52S1q1RswKp4UbTififNjIRX6hIAxKaPhGMF3gJp6
Bmx1OZT8Vwf0lzOoskfoDXkQeNAHwbtq9lJRN2udtl1k9m5hKNKwtiSm9d6DolDO
Sq1/6DfaEyCfVRdpVlqwukof1F1i+JkbJ0j4IFxrDafJuj49Xeoikl54H43rbY5W
XLPKbz+83d5i/nflHfiu6O5awnVTbcEzcSMH47zP/ze5MKzQQaVdDJFKmZRJW1Dv
mYmfKkL7CO3Djvq4LTyFcGz4fDqNDnRqaLtGl5vgwStkzijPL5lGtqxApeMnDHLl
vl2MmgNyAjR9XBgcaA3V7kbTTWj+oM9FUtZmkytYX8ifE8vN5ezsevJRGyTsvB8J
s9v5Ehm/4DMG350mENjZAR842dmPqE7VAA0tHT8Z0AL6jdX2ZuBibBLbfbc7d/1L
Pp6yj4cFh/Y5c4DrJQPP6pTy/e4xWlf8jXuIrWUXC8VUgKxcqi8Rs+Tb9jSOyQbI
1SFNeBh7Q9EJBqFwn7MfVu/UNU92DfboMLFtuu7kjHJGxSPvrp7lB7/A9Of4d7NV
O/O3W8Bqegyp1epK4g4wakiGA277/8lvFq+FMNCJVndMa8ppkDIMtsp+dk7vShKg
NhGnEmKJWPzHoDPmzCIpvVOjhx33SmQqS3HxvQFc/1RkRpUT/0Fz/faJtuXVYL0J
VSxkG2Q+JRDvoT6tNd74sH/SZPHF6muD9p5wBG3wcltoIb1AJBhqRIanlICxeLq2
QyPd3VatvGdcrNcaEKuWL1rYcPuHWdsZ2Tlismo/K6OOwpU67B385ynu8nEWXx1U
N7F8XEeTN1wtbfAd1XNgiJs0AixVV76wFlzg/IgfwAdgm2bsF+6IXH1VDHagazRJ
1EBfTGjH+Of8vF4dFhdbtA==
`pragma protect end_protected
