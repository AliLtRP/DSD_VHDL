// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:46 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AvY98GMoOUK23OKfRCkwZo4qyR1+Eeiz26M6+Q3VyDxUWuj859RLnTqKXOt4EiBb
e7b7aQsLp3x82ooaXSMLAvDc9dZs8Q5b1TvecrWwNJdnpKzo6BrpQFKXROT/ekcN
f/AAApvZ0Ors0Ebmnok66F/anohf1kv/POWiLPDqGHc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 43552)
SE7qIv149UYxQkijBGXBvdwF0s0SCl8WXAOGUZYZcA53PVYGs3TDJtVItL/LkB8U
bN4BUAg4jl7LhHg93IOui+UBBCvURFieDbGN1657hA77zXtaU3GzHWJqadLShfyh
1mesfwvV9Wy/+giv7o8LRtWgVfmYzDrq2T70lnTEmtbU9GO35DKYWVU/j/vn9Muc
DUIV32Z8DHG+YckX1xD5wlkEla1rtMD2Y9VtCcHUAEyBBf4f4nPBxgM3VAQBYAg5
O19ReM3XRwmFLLvuekXmfRgyVCge678Zg9JQnRvs5yn7+SQsxeG86ZW0YEsW2qqm
ni6Cwj88srx14vfQRxe4A1tUuLE8/utzlYDpQbLy3OFGGx+hKhIaHOnXdxDWyR/R
6WqKoQ0jGZEPlwK3anRe8IP6MrBb2a0gmyuwcgqW446CIBkC29d0IgVwuN6GXyka
MEYbjp0K0DiPAGoG/xL1XFcYAIHtEBVOrd7KV11RJrnl4x+N9V8RfLA5b/l61jt8
7QzYx75CEbZDvDZnVHfl+4Q43CCkeMh/TN8jYKNweaM/xDLunIyyPQfcFjWbw4u3
yX828k9LcLKQekBBjAzdPWfUpigNnugRvlxmsMM1UEgjzAfabwWengPPohDrwbd/
JrFyRsOF/FNbBTe2fWxjymfiO0OHolWe7vgxpW5XYAn/xV7naHEB8xrB2vYGMhmF
QotVyS18g8kmodMtdsGSJsGdpjVLiTvuf8DXT7jPSeCz3Ii400Hc//hq0Ozi9z+R
LWkWh4zL/UiI0r875Q3XWvWWr6TdzobxFxHKrTZDcWE7MhcgbqtswPNVj2uRn7RC
v2dehmOwOpKwxbIFWk7IaTAGP1qMbBXUie/exQoPUjVBpGs+f97OpqTWa6CIfS6g
LFJ/ywh72hWaH0SZqx9K2EgJBCaZG7UYXH+yjl5V3686t011stdFjRkh/FN68h/8
qinK27NRF3YFyi9eIFs2/7mPoy1oRKeWg/h9Mv/n1iSQGGly0bx7eIoGR1BeXzFO
Ra8R1oRPT2k3dwmGs24WGWg6DiBT8Xn8YQfn4ZrlZ6+jYLTNW6CXVR5Oqp9Boghn
GubjGGJ8z03fmHN8E9rlTMAaGCp+hvW62gvJUOPTRaCLK4mQEbjlTfS9YPiXVDOX
VIN9JYWxbLTFjvFfke5eZQ+uixtI6sxwNrVtvARMbuh3h3YkZ1Wp0WKZgtds16/U
5+anhxIOrINw2G35qj8Xxjq5FEh5bvNF0ByiU9luUEDsCbP/5bNdNiwax4pbJwI8
B6rKo34wfRNKGikeaNGz5kHlVau0Sg8xSsLlCxVFowpDHKEmWK7+yPm9khFG9BUR
+ppOP/UYOxdiMF9tdQ2dU4RqfIPgQR2ZW4QMfpqAKuPiWgMBqHTdpyTVJi7910hS
udUPj7Jl1A+90LIvWdlHxTAwqBNowzcnY2rpnc72ExbMEP2ILSW16+S58z3DJYDz
0hUzBoU5a9+5gi82DXEYuSR7CpltzCK0EKRFihqQ0OaxZbw+ilMfo3iIkTIVx1nl
24atDHN/Cv2Z1W8o2ZqtsWdE9/UBZrasxuz1PvcpVuhbi8f7R1wuw+bXU2MLoM8L
Slt0fFZL+SGefG1s/f4gtM81EvJTOU79s8oXDaOc6Dd9RYO8KgTLonMc1KLgqXRO
tEeIqGbugWrcXljGsjXn8pbC59IDCdXiLAhN43Wxlzn5o+m2j27wJyUN2BAQ4CcA
Bu8eof+satp9KK4ewsU2mT5FIcFXigJ4zvcAcuLM4EgMVAG4y7YVN3iq0TInm9K6
u6iKxP1O2ULna5z1mc9c/GjoRy4wG/vDn28sqTBrFYr8A84JSlk13kBT2SVhCPfz
bojCjm5W5G36rDr/HIdZeujA2PRavVRtmeKmZA6oFoxAH0FjpPBUq5LK2tP/Sqka
Lb2z84IF6MKEPfD+Q3elL6sdwVPLjFVYNSDF6KIzqjSOEakLudmhI7eDwJL1K53B
0hF11rwoDb0FqmoVVp+SqtAOPaWQ6Kq+qgMKYeMnZKP4cOehNkJoa12ru/jOSZ68
PiA8/LJja2Yhuvlc9JKR0PSpASp2NojBNVoIdOHJgM6SrdnD9vUbQ/a1GJVHBXpQ
3uTuyUUDtFfHoO/8g3Tux8GPPptXq4Lus7QwV/I7qk/9fz/7YOkUQ/CnBOMghJ2Z
a9yy5f3Q/dq8ai7FZVIjccq/qY5R9nYJVja8X2rck0j3mzkHIiQc8IZEY8PnQQ2e
bZMDElZTDN3wd+bhChQmatoQY9csZNokzgVQ9+wZkYSfuJiBGLRh3b6AltGumFDC
5dUU048h7B5wpMOKn7slXF3u/2fZ3+fYoXdbACkzvqoWkejNlK8AdeHlxZEfhGX0
5kN5TV2YPF9/3DRA/NKka7j0AQQtiyYgjh6q7JLBeRiti48uglfGOheGZ17BmP20
JDRhxZjEpbJlCxKq/MOlKWcRwKRd7iBLUE3oe/JKwmF7PtfGzFjK2OP0oA038k9x
u5B1EcoJd2newIEOM9LnEoafFL7FDX4b7BfR/UuG93I5y/qP8X3ABiPbz5rwIRjm
zAlbwGZ/0/FrCPAma/9yOirU+pHk6mHuL1rSHF9Zo4qWL8u1fK1yvnxX2O6D9BPo
EoXv6pWnVJaq31HqChO57f8DQoCop+hOPQtYS5zbXl8nMFL/aJPbljno/BTqAeaT
Wmr4IW/S8QWmPaNFu7p4bRxdQDp8ECmAqQENCkRga6bE2sSXAs/6AqyHgF3fDm7e
rrKcqQLwcIFZ9EeZKBlxtDxDf8roPOaN+9PNzQ09Y2D6UvneJPcBje0gWVhH9gFs
2jqQCwYeNM3yAZI4XJWkzNQFyCdwpVf6XkwNELXFAOd0oqYlEzT8CaQ177t/Gxuq
98BbtZlycxf2PGlCJPvi+EeheewwWZKi6EFUVIAwwfEaxLHTLfieos7wqcPyqrSw
ix7JuKwKD9hgfne9ZUGoy3DBH43cCnZA6/CmB1Zy30i9HGGiA8fSmD+DZDsgR+A2
Oq2Ohzp0LgNqZjVBx/09U331CwwKI4nGLEpnzyd9j6HTYNcrhDc+jCvTY4Yc9qBW
WYugfDQ9Ya6f+WPNaZVC1irWa47x4+0mYjlI1MzuPRibINUZ9QGZLfdJBESVuAdN
6UhRgEnU22UiZ+q/i2Ky4KT3NWregt5zadtfXU9YB4WD2ae3DtAlLWzh5qzQIFXr
zcamz9+A2D/kT4pZwiKyM9PH5Z3OD7m9Cu9AETSoPlRaaOM5RvOnw+XrrsfmTBHB
eFzEs+y5Q4zbf5LZ7tZT177B8qH4vOubJat6EYRCUC2e/vLqvBCTH/lz1LSdV0Qd
uRrL03P7djdmqb4ydGSE8B3OnFHgeSAejXVDtxzu/vdA8TxAc7GTZro0SGKsmxX+
dYXhot4L2Hr5I9h3WG6WZt7rVV1jEMYOHpfh/PC4KCatg20V6zhgQIPtXeSt5VJo
oYu1xuReeABDaeSfgdvOTqx8rd35fustApXpT18M21AmqP6KFxPovKi/+gXZoZel
hLFrzkHWi7qCIKibZyHTavKjTLUA/FlF4eSy8KCNsqAsItzAtCAg1dOmQ0gG2cfJ
CbL7tgmihQZRyGms0B6XR8YvD79NTSOKpqD65hBGE0LoaastvgdNduCDuG1ArOEM
rC7Oiiame4qqTWyu2gBwPR3cVBf5W3q7gJPSJxyU9t2KJqIV7pGPS+M6FP3+c+5b
DrQFZ9R+mQ3u0YPu/zMkYmfxYOoO1QL7awBNO3Ylnj8JiPQDr7QfS565FL1EEtZh
/HbBWXKZMx4dj97c1JMPTo+I5uWCpozoAofpPNm816qLtlitanMu6s9yP+rlgg5e
1ZfmhyTmD3mYhty8EGvZQLlVeCD3yaohJcbULqAHbek6PABMJyXfb75DOoqQKRqC
eyuH87cMAcGXAOGEqEp6uIfIFFVa63M/Uuyr7itT5RP/vPaw6RcWDdsYFnjsSaU7
/shsk48iPJ89dgl+0ImFmtbewWERo+F9FtDA/IrXeG66iGRvnN+a93TxjXcVUKjI
yz4PfdzCwv0LWr0d+tj45LyJtbE8e1Jys54L0y4RODjhro0OzAm1Pvsjcp9cJW1+
S8vqMpNmMG0kOKVXr/+oadmFzOJbkSCegw75pKJnKPWXzIeN/I/F5uGvrHsI7pQ/
YTm9mMAFNe9cZFsHzu8C1o4mWbw+H3Q6RMwqKE+VZ5C71qR+vyA38JAVsphlUWgu
TVS1A2XjzTnxzngdusL1uhgx2Tj13Z7snYJqaH8KxuuVUek1FvPwAipPyxnZLeQF
RLzxZz5eQa6lzokF4TlO6Lu8hX0+I+FKcr2CQl689DgDaf2u9F5WvHFu6X1egLB8
3LO5LIuTtDDk7+fDJ2hd8btrFmP4LCjsrKXsLcP5vBAGZCzCCWDmIaW7g9mbvVTw
cE9ZP0yrlo/RaPH4GdPmIRB39R3uhUkO/U42bRhTuvuDFmVDKlNDKnJscaSbDD7+
voVVdsKLY10Q2WE7M2iT9we3qud2ltReQVerjIaAoVsfPX75O5KFKOBEZ8KY8n+Y
PJQqvA7qje1t8AIsXt5sg2vph6Ds79AjJhOCIP4nidIFwGldH3SXaCDyKhI2stTk
vjd+xm3DK7CqmOBTa8Scvrlv5oO7DJiN3eAKWovuFrByfsq0M44qGiCBdO0CTOnc
j76j+dNH2J71ASNjEbVizr2ETa15Bi/2BQFesdoAosLdZVaCSrtFWxkAYzyy3dzn
V3fsClZIJWmY158e6ryB3VwhwoXstno4VLW+W/uPNKp8ocOqs5qwaQRpTHQvFlsB
XqFqkIA+5c/y5PihIw1wPkOE74EBzXr2fh0dKEiREDY8DzLWBAUCYynCkAPP30yF
18XXynLkGXAimIzcYyG23G4WaZS5P0rPiWBVzJLNokw08n2/dGz/cHkDr5sNeEFu
iA/Xe6+IFwT2G7yQpwlL2JGWhdBWbq4L5jSiCRpaVvO4EQgrUoh0TSNA5Fgm4pI4
r+6iL553+fnzvWzUDDQUlEt8/xzcLRv7bok+Mq1wqWwFcX8V+xynH5muu8Ij2Wlj
RBjll/ollgewB0Xm6MZXfXuVj+lE9CGWJM7qZAR4+zTtGKg4gHKW9QIGCOeUgbHR
elJZONcMopPy9rAD7IJ4CVceMg4DAOFB4glfFRwFyD4ltGJuDnqyQNbb/jFOuB6H
Uh828oAvcLNT1HZ6nvy4GcLiXFPuKl7yZHcg4+xqYpEXw8OWm7k1RsWwKsMbLSx4
7PSXXDHB9ktt2ccpc4ciZZZg/EaWzZv4/sD5WYXovLq36s81zd7HWBRUdE06s+7s
6C9c6MEEmbGThdfMFK8y2IshcExbpC/Ppcg1UYDhUrC2/snRmSNWVL4sgpnBh/Mu
lPyH4iTT0qxhK/4tq5KCzSUq9fhtiofYyOaU1MHcDpfmfamOeFVEFw4DQUdybNdc
ans8ehWspyYjc1W0Y800ehXN9tYsQlNK5zsJn75FP+yClLbJ80ZbLt/bL8L0vAD9
jkTiq9Ekw0Ci1pF29Axhy3WQYsEU9DOpy+eBAgwXgAKXFBxP+6+i0NbgvtqTUZCs
zHDHhc8oV0+NxWmkUm61136GYhDDEVXIxRM09AvRwdnjSTLaCYzVD7aNo5YU1N7I
CXX/4d1lpb5qBeIbT342GWFbBHhM/zlPRTbutWo0O1pMzRYHaEhPlFv0N+FZYMyJ
YhrtifyioeDeGWDheU+9ToWfa+/lDbZ4HbAsCyw5suxjjGyotUjltwu5SqKZ4lOr
HfoiEGJ6MqyTMXw/jTRixQcMrfpcqLre/Oa4VKoMohAG6wx4JH2MNdCYwpifqhfA
EdZt5RKT+q3EVuAJL3PTjVQjkNcm0rwbngeqoQsfD+LkCelFnA3WlByvM/YUE7ll
sQWepyjtzm18uD9Aj9s8lF9sCHYkkDw8d5IK4FdLgyU852mKVe/QuF9Wj/wmnfRz
9qgfb2zpJFJyyvWQoWuT7o44IcOjy7njSj7Fgz0yc0ZvQtd9wrV6ramP6/rYLgSP
x/eNfeV74NJJk++COR9mtU1bP8+KfsSJ8YKN9YWC+TiqvWRG1mPB1RpxTsVtkiKJ
obXMalc93ZYvKcOc5Kcj+5J/4MOPIGJL/yyYNc+UimK9ByPX++xooZq34Ryss5/y
OYkWZWz2on1x+e9TNpjCY3FlpKYhj4edD7P6oBupeVFGMZjYN5dxbU7GGWH5Ih63
WYeitut13N0cNdZYX0idgjWeJHkqM/sM8/Gt8F/yF+2zwKQ3IM8qx4O7RhJNGuMA
/rfH2cz8400TEaMsvWc9rSyR52S8fPmm4n2SEFahy0gK4s2glQrborfFBilW6kin
PB6DRmaRNNap3CuwaMKG5p1judfd3Cc76y6j/GDWzKFcSAk1H7p72yfmc0ey+Z2d
5YSqn7sLX5aTk/BB/6nB8ujQDckFEwPAVBLKLB951xonU+2QT6r76DLLT7xfy3p5
8/BbYNrop4nu25BhDgG+gXa+tyClftjjZsd43q/WCisV5KN1b6wbfgzOL7c1Ugaq
KnI1FOPjO9+HRoFCA92o/tQ9Dd4dW5eqdOlAL3b6epjf5Q96jM7CrppM7TPfwelX
tPuLd6AtgVeXaDK+jz/KR0UDWbE+WeVNDOG/fV/MNCzxGN4MLO9OYanZsV1HhuTH
4bbMgnxZFCBEnq/bCZIpA/B/CFNLFFIF6SC37O+PEOryLEvnugAbvkfBwS8mtjOP
7za0m6EJROPIfk0ED8gpOVB+2pyuNLcHbcCqIfisDzKYSW8NZs3Qq+zKw9OKtLTP
iGBXfZI7bcZw5ferwcnvD0BtlxF531hvqtYBuOPazMwvuRK7MusjWKvN+daOwy/O
pZP6YFFgRqQLVk9x1znzS/nn6k4uzpmCQXoh4RtQmOs/UjMLECwQfq5VOqQ572+Y
xsz4ZIMRgW6uFQ+o/PAR0BjWZOtFbWSfVjQ066k7olCiuN10eFz3RqqqdIdxpP1o
p6loRsv0uhEmIFB8JD0UXVwEKqf1hTupAApSwkm5IHsSFsUaybohb9xZNI69seQH
YckkbxoHQVzd4ObFboYxb44qTxNu4CTw90i3g8kkkFlyWRSq4mb+VMn9732uY34r
SG9ooFR3Oyc9Mj4u/2JwhZ4Wvm+n3NFGU57Mv/VcgLY5pyzIu0pKKiL9itEKUv31
wmQBBjWfdV7JyPqtJohNAwO2BGF+HBlrld0P6wZufXaerPHrjcbL8zL1lj+XGUbf
QXx1g9aT38rzFlCyCKWPNn4nJLsAY3nPQEAJspseypDZY5mbwtBeCkMYYuaI44Jd
8kUs+k/qq99wZePj3tZ2k2k1crL/KxN7qUBK4SuULNFQO5GVxWtvucHy+AR2SsRJ
/QV08Dg16Ak6y79OfK3NckcfX4X8yRRfH9Q38jcHPbNHFHk+wzl815uRe9rLYQJR
7EklS6mOTmvXwhmtlG7s8Ho9EgxZZQyfehRwQgeVGvkjxsX6SO0Rs4bdTa9Vfl3a
T5VGamBAOA83jUmFRM2psrjBs4UNOvyaI2nMaUc17RXJJnAF5L9sdqO8MBp6OqBa
de83bYaUEXmUz3ENloZGjRE84SkPpBxZqg4OUySf4X4ZPVRBTSlo+X9oh9gLg6gH
SaFK2ZjoEyoXEvVki2HNw9DwB6uzijuRuuvJ+MDsrk2dSYYD2Q1OBIJS+U8sSsC6
ntzJFAVl4ErQJgxzu6ZUkSL59e1SNev8prXGAJatmDuQuTqg9058+6fOxy6o+ut1
dzVssPkxeDBiTo+dePNK6ENO/Dqeym38dJBMknwxklW8HCk4WGMHwhJpRiRs3iTU
7SMW7y4Jh+vK63Idu7jZNyAHvEwCPF9fwEw0kdNmJEQzC3MYP4LB/9hQrutZus65
h1OJ0+O999czkUsRbADd71s7XcBuZV+SxOTo02igcbDLsONGgHPgPyW5MeVuHk9s
RnVQWsUs9Oa57O68+6eAc+rwOZKgmqcQbtidm9H/DW2mMsLON/xG2KGiVX/Hu33w
xk9GMcqGgFE3hB8SoiPpRhQyr9it2R4f3NAqNrAH+ql2RMbT33ibP59eDtgGRcra
HzaDQ6MsKtCXU6n/y0RaoLUsJAAukdLWX7oTIbeQmD5OCpl1Bq8ydmvaCaokqzBF
ADyq7SbUWwZnpXKNwYEuFcP3mAwLE/0XvPsGra5GHpEw2xdQIKmwwGrNfJNk4HSI
h9Q8l1gKr+/gZOL9Q7Je0s+p5BDbmf1WQKYo0En/TG3sFo4OGOeFcqX+IryAVHMZ
+l8aeAxb3JuOpGF+4R+84vemUEEUkDIDipTy9je6XumgDrNuSdAJpZr13EIlFtGo
Id9/EvrEmb3F4Ry6tnKqA6Vst6GAf9zKbrFXz3ancoxO6j8Rdn3Tc0Gg4K0PXVHp
ucanMlEnyzKKdwrR++gbHpR/wIWI2NF6qj6z8vPdaZSnFi6fC4Cx6EQENolQxDkF
NHXiJGlwwzqTDwP+2guxcS975pJmuxjL12e9PCQCNBeyi21klOFeOn+5NS8hAqYJ
s3jRWZ2DpGKbmvwlKGzyAIX1Y4IGBAal/W2TZ6Qps5XBJWtrmk8g0xJEDefpn7R4
cIXbqdiSjXX/8IPu2aPJrxQIGH/wq+BdHx4Jc23NO0KO1XGHxm2FMIZRPGBoJPKC
Nz0PKWz2WboPhuLxXRFOF56ECo6DerloVDo6OL+L7qR23cwVcvd0/XN0/JrD4ffp
sJ3Ma35nFfHRblQJY5Br7Ebs5MhoGzcUQ5nOrWJwsQWmlK01DOwmKiGMXxFrrnXp
Ej/oFb1yTecg0yGk5qzTFFAgfzrdjQZLhQaqRbhjRDCCOfkRO2SFxZJAI1+cYHvj
aeZpNHZIsjElOCIA4Nw1IRUHDVe0XMRy+fFl6JbJRasdcJoFZMQbOFH21kO4wou0
00dTHSJ2NnDXCy9PY8LTjfO77G+oIPWiIajk/cPBfitGP5p/U0JSwIuI2Cf/nVYB
nQPyfHUO8jP2OGANtRQMeLT4S+Wv2NCHCJ8PU8kORNFQkCtxborj1XNxxjpV6ZgA
1aZugFo9C/XL0XkxU7LO5skiks7egEkf5UTR2djps8P/ff2aeVuGcr2CBVFGTBTb
O3dR1X3oc0a9VdV1Jle98+8JfCl/bhFnQph5ysGGPNQmWNIqJkriVEYPkQRgw0Ev
xDSZLSwerfVGm/VuyH62I2qfNmUIgStfY+lSNGD8sAnl39f+ofx9r1TMw4VTR1GB
DfAySWXsbK6r7s6YdxiMmG4IxRnJPvashMgrQ+kVIhgqLIF8C7gkwXEV6nY6dkwE
FZIhqk+VSAzzJTa4ywQZA7NCEPTftsF8ffSDlsK9FGPQKVCOZHISEaEr5ZP4ijGc
xYE/k3Hpylsqqrgl/DUxUUvM+i8ohaQ49L3G/2ucNML6w6DvjmDUqP9ptm7KEyGm
yyQYCRL/9/goz2bYtUT+oyyiU8AcxAHrTOW0oXYO5Ccmqf9WaBLPNTUqDoWDfjaX
RK6qy4vmaTYVs5qTzqpe8dgrKp/FGQDfUUVncH/JEJqfxxLts3FF3GinswHzwaAJ
dwvfixFP9HVnZc0pNQBsGSslHVIeK4/Ezzq5QABX2FQwIuppbOVukCyX6Bzya2rH
+UrBZKuDHxT5+Cq5oAa6nnRbwSJXSp98VtsZ4PIUsZp3P95w2Ra8Wa/X38LpiimA
rUnB7FPtIK1odEt+nFRgya9dmFv+OKOq9b0idZmNi2X9ZZk7FSLvtPK2RrDuUA7O
lRoTZciVItyWkt6R6wCObJsRBSbtRbcYA2fZyc9uNyB82tqweLA7i+DzICnzkmoN
bekeaXApKiCj0vxIEc1a+u9rl/dtUF2M48ghu7XNlD0DVrXcdy3CXxoOoynJd3Bp
Xj8k+QC9fsXAZwYqTAjAcMrEGlL/DthsVW5esqScQfAPGVy4TKa0Aq2b2silcPl5
+RwAo3pIUIW5AGEIZEzTDnVRWtGj24AwgN8qZdKChqnaLYmrxfdHhqa+cMowlZ/2
QhoDwbiyr8lhnsp814XDljeHYPggBY392aq137o49m3xsL7UeMy+QWdwGt5VIVdj
j4dBVjLX7LnILXFnn1KKjKqlkkg/EKy+2aJDJGhRrzkAvPD3FJ4CWU8ojVveQaKE
zcpaJbbnvANanfJIa78FYqN8tBbkNBDCoIyN+oaRQ50i9AKqxdCI2i2i+AmYSLEh
rgIM+P0nO/AaCjk7+D27hHsQui8NUbW/YooZoMulJiFzVmheZI9G6sF0KoIgMbht
+vnYxz5fo0LVTFTkuZuZ28gCxxCDxvpTMafQo75QQW1ttfEoUf+1JL7oroflWcc4
xVGTK5iJHWVkS5zQqdXb+8CGeRCPs7H0/UP3elS8hLNWUUFM56ydfSQWIjNQ4Tqz
/wYrwOGqRrIOKDJ69qUovF8azib8V6ob6tkWQRky9Lh4W1sQQdI2e3xclsA7zlqH
r03lzm+vxw0H9KhqBtPoJOwTwijHU/d8T5IlXSNHx0r/nQbg/HxTkRza0U0wF6WH
c8xBy6vuJCi1ckKoQ6wHzzJPJJAtMKdnE9Ox8kD+9zRombvu+oBGeIZ4hvFnWBBU
V4gMffx471D98Wb2KY7HI3DnwS6qKtAsLK0yKcqCEc5lKvsMCsELnegibfyjgR9R
ncilnjuZDNnW1blZIQ4VHDvUykaU5dEDkNUgzLmgxppF+5PRu/lH8Lh3I+csWOge
sLZm+DLVHtZRrU/gAcWK/3nLqODkyiPsGPHFPkE32AztZDadHxuP6/a6+V6QNVmQ
HrcjPj1IcHtkYw9S8nYqrwsU7WwM4JSUq+tPoIQLjInHORzJW1091kBdPsJanzsc
W9Pq9sy5Bx5h6XLovmX/66faDiNI1pRT7rcuy0kKJRU8DpHt1lhLv/pbZ/WPW771
7Y5lmSeUBEsSRrELlZNNxk27wblWKj89QTsFmmdR77XrEePE+QTMct0KOBFithXo
gc7XV58ebzQDiaVSSDC0PBg5Mq2xbVyYfl2UouiQxl1gJEhh2ojm6Z4iVk8Wn7mq
JEKuUhbSAFCHMAVQdqfwb2KergpUMeao+zQdP5SoMg+X3v4vQjJoM3ykvte3tY60
EOv3Q+qtNL/PulIcc6bVqvrVts3+cS9jIMszC/0/xGWw4eRyZ+zS2pVbg2iXJB2b
Uum/ofROlQLA3CE5Mq0VjyX6ApMBnJuGCpYnLJWseXI4gQGvktgNAodnIcjuJEeG
8v0Fyr0wnQ3E3EUCxRVkY/9BYOcRRWlgkIYdGtjL3zEKMytL2gvDykSUMNzrg+EE
PKfobjHZjSSi9Qdhni7r74JzKkvg2gVEP4h7crWERjJU6LeEPPjgQOwhoqgKf8IG
H67bqV0cYAAnfHcRAgpUuj8DAEnCgzTBs60wrKVIOkS3TMnwBtzc+lYG1aLNNsUH
GgVWs3O5K6g+PcwnoOL8dxocnUdokbtBsDoTeqnAEaaCqAk3YkYP4Ju5/uCnQhFb
UNNc1pes9jGkLwAaDO7LAeQ9oH689MAGBPUraHMTEytGvtyuftM02TJSOt8IrqpF
ZQ3J6a3uWoGGS7rOlypKamkv3n0hxVpHrlqTXLQkZzIlQ49swVZCHq02oNFzWVxb
7QyOdC+wuJnoyoi0nEJLNuRhO3XPsEDIIwmY7jil6VFhzGCpwCd+m4cjJWwM19JR
LMZpCc970QVf+nmd6cSCs/fLytj8nFjCGEDKE4fmePpUo3++PqVBZy0SqMqGdcv1
gP3+HQ1QAoTPxD9KsoxwSEs+JiarL388kayiW9waMDzovcBLQu6mZ+4gof54wu3s
QhC8bkAdMb70lwMSEe/S1GPmt3ErZSkYwiNhFvRqI3PWQZZVFhDy3ko7jXeP73t+
faezCUFah4ZZGZOYoB5Dt3VxPJ2bXzCXc3HKlLoEXS6xhwDtNwg/0r3yhWrutKjj
DQI25KX5nly6PILqFFktBp8bbA/R8ZAl2HK/B4vh0Jb+UnQ8/6bfLaHOlJqaKSkI
gR0I481wYcm+qrG7Fu+x8llNCpXRIfi09wf8FMZcvoT69Uv/Ek4gD4mGEJcRdKBE
OQVvPyEvRLeo/ceVKSHxHM4+Kh+qfJTmpFHUDyPER0TGeagOJbnPxn0WA0PNcdeS
Z7JXF3xqtVaQI9Ipl6ll4dgVCc/T7SxGqj1CKlL8w54jbgwEAX20LYZe42q9XmU+
KV0pg70wnYsYduM4rIuT4yXhmklGVxHuhEn5QlRpXzrVLOGaOh9ZH2Yj4Fh0rTMu
LnQ/est+sIKO22JLQJEmGu4xMlVwHftOWINhvhh810PozT3cIg/EBMQLPAOPPDl1
4nwrEAtIgo8dOT+Ep9TYU4jadHXmg8jmsxzLCnLDDXM4NYkjvDGEZT54SnDFGyow
QOjcqYWiQxsRXSy+Vyl5xmhMrC/RfAHeaOrXz6o7l3Dvd7pVnH3K6reD7IMggJep
oeb1blSIuTsx6PFMJd0/QiAFt8+8k7iAp+Z8brhddPiDu97iZIrUTKt+6cqckLaG
hbWFZ5Ym0iV6J02wHIbf886gmpWGmT9Vtkg/cAvNCTJaIpxciLD8e5OueuvUzwH2
ng6/i1UpNerCzPkg9gh0x1KjTuwcGrHwpO+g0uPPmAGYcpzWEN5pOaj1MkSYF+3N
5NW7n4VqZsKwZN3k9rAfO0t3Al4rIdoPxwNY3IfDF+eQtkCpvCdIoNkyySGisWT0
xC69z0eSdRdVXLj8v2e6K3k/mcOSj6KfbRrYhxE/+CFjHOf5ZA7zIMoK6hcP7+dh
2ZbtLgpHc+zCxGpi0zaIm9TsY+UWpT8TeO+cQoDIpeub2wfwJZWjVienjg8osv8Y
kwxr6GP+tS0D6pzhb3B4SAnU9kp8MktqAl+vLP3epcci/Qac5eKUHkrQqAMb/TrD
2FS0A16XFmr4MT9wvU9FvBpmZ4AKj/olev5/LBl4I2CH2X0PC9ajPn5c/nKVulcQ
CQdKP14e7+qZ78sRmMFAwhH5HQZyEv5l//X3f2Si+jBVGoKhCPlM4kbXkR7/cVD2
OCiV76sv4EmPibAT1HmPcB9btTaxJObzzq65ElgJgW3GtU6HFoIAAmazUsMrjLSe
IHZblwH1F5MTg/sNXQwZrkmW6oVUgb2ii8QIdxL1MGWpSpT0BDwpJSn/3/+fFfl5
tHlNhjs5iR+krK8PWa21IbjiA5eGGnq3KzfXCTypv0QTOr512bGyQ/DEkjAwpVU7
DNdZj7tkUHfvuXZBGmjyteAZoNOxgppY5ELmSl7smoCuLHfcjLA+Ks9shqQPLsKQ
LS+U2QYaKyB3u/zX48OsCdAhvlJooYr2P7YKjqS17g11efBP+5DuScqoVcRDRTjr
GYEAL9jFvyo6607kZPdfIfTDGROWUYZOYOwXM+KVUfiYuis8AfIh8/F1zLkz447H
nbsH98y2IiUJc9unjr2B1NnwoHMlCIuwliZ1UqKIaEa1A7g85XhIa7PzlC5rGNYX
VEsV/+LtP+nIgD5iqRSn81gZAw0BOX+Tp4c/ZJNqW3pTR2SxnkQbKYj+mXpzVCSr
51WF8vGx66PJQ0FsxpZzQ0jj3nw+4DQ1+KaTIKvZUty4DrhFjy7fcqzGttNPfUJX
+82rknKgXOy2Tw3pBr8w4H/jyj2UtSdy8e2FMlM893Rtddm8MvI7d6xhEZU+zlzj
nrZdhgXGsL32cYvKPgpbg4CJ19azRxE8GcROPOfGtvj9WKQDpQyEKrogpRmUg0K+
69G8CKEoHUD3gNlKJbo0SZ+iFaYkJSvs37FolP8hyKhlbI+Uqiw5gYKkABmzXAtP
nPuAnRfA3EIE9UpNaKkPhKWEWY+UHus4Wc4ON70xbQ/Dr77b3va63deekqK+bztx
ERkOZquKwfPNKBmq0ikbbNrILb59L2WKOpjJxhRYsTTYk731uBsLdLy2md9NxR0p
i6eWOIxpRAxNzph9YnABDZt5B8i70dL5OgWtyjYjFgOImGzM33qFhrlXgc9xj/SJ
Mtw7cSbWwu6X5bI2qBIyhQIRRGufGW3K3x8HJvy2GM0FE/HHqLN1dtsZuxI91tqJ
w4mwr4eeo62GvRnatiKjOuKEdn5owoaTdohIfBQ7M5twgaPq0r6g3TRQcC9kFr7e
PveBgyACMjvV3qtB/18/qbHk97hTaSo5VJ0xwXalSdBeWGGjD4ijE3kqAJqzHGIS
Now52cUMJesGLCHaaYoHzzOuhtLdNWzwaz2fkF529opa1swEdOU3O+C/ArEdTlwx
1mNdQCB7CWf1DpF4CfzNsRfNejWLzVOZT08m+b6vU+OTNT6WVcmBtBiWrCzskhp7
qPPM9DWtdqWVluaxUoIig0HPS8LqrwhdRp18dOVVixqTYQ5blpc85exrwEYXgxdR
rRsNj6DgxQsIo7B7z3xDx5zWeLy/u53VRlLi2KD041VwE8JO6NvfclZ3QBdpI6uR
qmxyTO93jk5lluwWI0sCdirnkfDqWKy3+y2cH4FXsV44qJ4cDOaecW8RezQcVOhR
WOp5H2qEnPotB/47YlYAE7UWk+0kW8UI5Mg5/w1viFvTGcbjeruFJDsv/IKW+zTu
yzevK8g0zTnjPgIbyco/2NNPnKNPMujvylYlEgMqLa/Jnr0Wr546TWEvFhXv8HNY
Bw0Ucd/lYGuqwETbs0yXxHX/jw25j3I0bik3l0SeVAK/lXPZipCek1fpfwfR58+N
W4Yd42OP/e3v5VFxtmFEhCPX6mSnH0vorIudzSZG2ErcuTBt4pY19Owqe/Q2g/0u
7pN59lo8s/A6vsmemE2RaGe+FP0u5Ka0tyNpS0qwLPuRwm0pmr22t/Eu45hrZGow
mLvTq1n10cipGoA6184/Cy2K003Uba9DdLURqPsHeFLqaNNZ3YOZR3GzaB7y4Tby
TUBoG+o9GcSGPUaJoryVOKYUZ83VMnTgmGIBq/CW7N0SZixtfzhPQ5wE2MU4dBzo
g7T36lZ587MPrI2g1YN8FlqOeTcnoPkoyrNET/BKQab6MDfucWCwseFheZ68Otnr
a2aVeoNFfQCH+FWjW9GQn73hDhNZsX5FLT0yN15pUwzRrwubYpJCKwqpSlGhte/e
qBhwvmEMVG8mr+J4Q8EFE6achy1iS1pNK9qg68LgSO66d681id8ynV8SJoDqQOEe
XNdrp8E+9Thb9tXMsJ47COOgd+jxgXL7IwBNBUNqIbZ0M0Gr6WGv6ps7CIOh5H/W
/m/s1O0ys2H3pWxPkNevBLJY1RIYcwHrMBVFxFjliELfZRY2IjhDJisJaFP/low+
DZ/lJCKNIc5LmqMAVU7d2iwGfIFwFH5CapKl/p5wwW82yk1do2twxJxePvpVT9Tp
xKbcMlIrRZVUoGr737ociwWpAoNAIlsZEkpWNSIH0AWOrjXtzLpZKzjMbqK5EIuP
SE9LR6LkHu7MVbYXHb+CHpSCF/Uz7YxnOS4BMtEMBX9yUkz8deAsnSMUIfujojYe
eUxzwWi+I/USxdXgSvOQc31GSoroXkwanIQ21qvitbHHEgzbUHxvXAV+6vEOJVtA
m5wlH/hCMQ6zQzZLUK3gMX9SP3VfYJMPIdrdTp5D2Ix39NOMY21pjiEyieLG1F++
cnHwcnQqUIJ1adiN1DygAWonKhCzqHpzK0vKCY3sR787WiQe/GJmNkmudihnEkNl
gSADCmOHEOJJLMjge6pT1U0746NQTCALUVFW/DZEdJr/XKuB+S8Ir8kgrnHmYqGJ
DWNDL7dgVT1XUlZaQPgz2dTnJ0vBJEzl8jsRDLaFzV/N5b7pWLqhWcKttp5vF1mP
hcHUOjdxiWWwBfPmR/dlH+pK8T/WNWHsS+M8XgtHb4TEjLA87tJlP8He8KU7vrSI
1GsSHF/IxKiFExir48ZfiV3qDI98Q7xdbw1DA8bB11FvbTh6MsdaI5Gb7J1TKB+c
jPZPrik5OKKyPkUGZDXT37kd2x/ZKxioetCtUTOQFfOE7B80H+9CGbOocIG2w/+i
5l96ln/MYWDu/RmeL0eVlzS3jjITd59Y8DmjPphkOH7yehXbwMrLJnUoqd0hGaKP
jC6bu5JqDt+Qfvw3hOwgJYxU/FCJVk1HaWgZJPknSz2bJhUJlmI/pMwd1w9HZkVm
fI4t14dEbIk5IsNslwtR0gw1KbWbiZaPOjkQj4SW3fO9kYAnk6P/dUdnWhy2I+m+
xSQU+dLmfgBH4SR+QplAp790RvNYRLNfYZEeWoRFe217SUW43x6zsEAJDoZlNN7T
RUrGIXU6hWDNlPeuuqZY1Uyj3uRN1ushd8CKVGS2EM1DjjojdSbiTPJRfy9Ooi9w
CWvr2ghKkFIXD1kAQqpPdFZtsnq6rpwpv3OqvgZxnei3jkx2qQbMBnXWt4LdNqxj
+Bjb/gO+3S0pGV3DCsJKYz6zROohN9gVDcE4eTR9zKqcLHDO+f+WD3Z9jMnHy5Wr
3f/JF0PQcAe6DQPL+gn6T1dfpoJrcmnuil/WIYSzwktC9kzgQJANgoPvPbXh4O53
zkuxhcqmpXAKS3TWBkpo/BjfBQwKNqbzIMbQvejsfdT38FYaGRb+KOgX6lmzeeOJ
Pjc7bPtSLi8NW2Lp4Sgm+pFLFc7XYSijwaSow1L/ppBn0P8uBv2pezeUfbcx6YVa
E6Q9vGCb37fY+fQZdG/+U9RkCzYXgZL0vSuBtbqIgSdDS5sSyIbRALK0pgaT33+u
NkJd5kUzVxBMu4wVWjpE2DrovOyyqbDaQr/DpJ4fF4vn/k2EyzdprFJTsn3GDbwb
LZWeny49MmWh2oJVBJ2pCs3XWeKpNtJskdahnMkIw35EaRyRfCB88PRfOeliadAN
v3UZECSv1korXZBdgcQ3+pEsrl5sT7rxFH7NRHA6AkHUHjNCMp8Lsg99PuLXdEWB
pUvfOPqjycu0izlU2hec4sAwU8dEsmfZrnfdLoop2Ucf+SyEELioLX5DLjPGoWHY
9SqN77SOJOIS7dA+ds9Ou47364wFeFcObcazHeoludhLVTVnhIqupYiADKTveY/h
qbifxSumxO79Ds9bLYKtMoH4wE/m05j4rdSWZUfA9guECzxvS/H36TW51ItZU4Pv
MFk1PbuIOGqsIwz2XrU34RtLcZvHXT4buzHL/2y1sgv8iBhcKJlSHFC7Y8dGMGoe
2PuIwdX10z+KsASPA3t2tjGSKKjRQZnAdN9bw6GgfgQLpZ2A8JqhspTFHBz659XA
UtgFHMjiFWWqyhVqO7c+8AG+b9hFbO2RyO3c57qWXV+30I1QZ4tWbVrQTD9KvvtY
0b539vXwgu2o+AE+rMiAke4AWZwipDqrLxh/tUwKciJYqva2N1yrjPN6XzIBOKPa
wom5BjpC6791h9pNXDd0nsHjTuz3MV7JSBfxyShnGNqarZ4I698ufWYQ4er3tmHT
ibSHLuRQXdtjyuR7Ax0yIE690u6EbsmkB040UyELy5gG3h71ofurLGYEaN8C3NC3
ida2rVqTbmX8iXbc78feY17HITh1MKtLFEKwfTbkgVQfGe4M7mlJiHeqVL+I3DHE
XgCV+fgHszwF4XKQQ+Zj1mwan9bjuDZIzExguxuB2nRezGgnsS4a/2Vg9pLZ7GTb
eS8gbHHhHcJDA5+y6yEQal6FV3nzOd3pZINwageJm1XEKNNf3uYfh9aPwwCZ6Dku
r6qaFcZ99TPPp2PnOBA0NLTjeVDx9npV7CwJm48krwUIc8SYnlVxzCb4KUijlbdY
wYRCcxcPHGoXVcRftARKqFXV5CWJszrllxw5aNMh0M6qFQPqDK+H+tNhP8JqKLFL
UccIJgld5tzIUguOO50ThWGYzlCFoD5O17N+4QwAFi499yE3SQT9OfifoBhuQzYh
uVbBsNgV5lMw4mKlbi0JjgbIi5cfn6+3XWnCSM0rUedgfaI0XbNEl7kdPNybiPX/
LILF5t0mw7oRuNz7Z8We5doykpJeyuUiEV3MjlAx2WxJ9lG1TdDBUsf7PnjTA46G
WTtUdYJG139Ewg4JH1nP9bjwoFYl0GrD393jSFE5QEQC2q/mEsi2gc/E1v2MhHY+
uwu1aSM7nG001mxwKHbLpSIM01yqlxvciqBawLTjhM+42EqAiFXKaZeUAUCLg9Hw
c7IZlJjAQdchweDtl1UIxofFHQ3b7tG/AcO3kLvROZYD1te9xvFgXRisaLy2Goi1
HUM1hq3tqOKH+n3T+Lupc6T8IpiceApOrOqmfL9jMw3qxyR4BwFNQ6U4xPs+poFt
2dRAakRe+cYTPgixuzI2asjpFJ3JYfkdsLxL2YKDFhexIrCbjVMp8lCqyzbHjrah
Hi3bX5ZteBeizCOzaLT4sOwAM8RJmvKdQPjE6U/U0ADnyYhaRs6zaACheRCmRE4d
nxsEOoi4ztMJMKmD0nPBwag4Nf0vNYIaPHjxpszDwjj9nch7Fhpex8IZ7+/5EnAw
Ll2LkMfTpK9YyPTQ7JNIU7icqvjZnAqLVVRIEa1mMm048K9m4i++aseHG/NyiDI+
ov90nY7cx1iUdfR1g7io1O4UdlBoDeUtT3ZElNWVsZ5Av6OuINwTx3TqBsQuzys9
+5NeSq1dTWZzuM6yv0w1zfCSBmQDmuESIkmXMh72jeTtp9wYPKDJBtpwSkIjqLeS
SyQpa+uvSfguu86HS8VdJJs/EWUi25B1leo0qnZwcXDncmbcDI1o5jz50txu+HpX
Xb2HxXXRXdErIHLXeeH75dOs0HBxyCHLjBk7p9qhIb76AXILYeo94oOsBBCby+e8
veL2O5tG4AjslAg879np4mvW5lglQDj/vC3EZ9g/oXiEzDxtiCiqrZdn/G3JH4WH
HeAtxlfRR4/rHzMRpFindR4u+BWJh8XM6l8QZRBDcFAZn52CNoc/6V2O5E4N+Dpj
tJu/SttGgrB5yuoOqig9mC16gvSNtevIxkh7vPy6Xlx3A3x7WLxPxNTlGFFg8ODs
MTrLHrFc2DwpFHlS/f2pU5leBLjOzfTH/78k4Gdoadm6PYaQCyqCBemHQq7OdlG8
qQFq8++8vOOFVzkm6zngH3eo+HXSd9zlvS21BdAUtHJqXgYr4Zl6BGpPCvV7P/H7
rRKM93+JTcmVkcVxzPwM8a6nSra8nAW5/XBVGDDpE66IUOl4Dh1GyxuSISf3D1W9
Wn1XbzcQ/WscftjYi5gNtCoTOgtXOUuFL47ex/guwAIck79RB+e1d1p6QrHbXups
4st18b9hHWoQLwmbqZwkM8iLrAFrEir51y0H9dk9nVblR1o0uTF4+W9yqVJast3z
E93mDgaoelBpFDTc23SyIql2QyvdXe5G699UqMF1/TDXI0WwUl/inKDcl/p1i2BD
GQUXcWUkJVphaYbK6Vtb0h3JoQaojMBzAXvSzzpWYHWXBlYz3qqRxgIu1bMpMai6
Bmj01kySRNa59kL1YXlJ6TrlxMkD3MUNSEMA1ANQEFpSDcmcM2vVHQcUWO0F9wtU
NeuDtjHPUFIWPlfKdy1JyN3pilX5iHGdVDzd335t2cY1CDjENFgE58jw4EejDZSs
iRazHgFcgHP5GT6vo3zXi4qGguj6X3I1YIaDXYqISaR7NUIDphQOFQolZUbLE7S1
zYvUcWlhnUnliRmwMh49J25n3R8qYNsCDZ7o+L36jmr1c1A/zxKQobLR+o99lULd
S+e+C8v7NqZlS0eQIAl6uINg6kh3fWoffWpuoPeev0IVNDSTdB0ybINaFGmNyOvN
7mbAGr14UMZuPCgC+J2kW3yl4QHIVLqGOg/p7UzHUEp+NKrLxaj5PDOxdhSlIrvh
eQdENn46J3wizWsjzstoMECQtP0RoMInXAzNpHPfIk3Yp1YbOVirhsFGgjeLTRpx
Jz9yylDusdF16WYhHU/+/LaNBIWR2JrkFuP1+9QuiCfLWcp4txGd4x3os17CLhlp
p/el/HBsC+DLKf5Oy2eH30qpPRWcr9yfGTzCT4T+mkhOL84/Uog00IVVvhhDdZKN
TOkE3thxRB4+CvjLcpZmblLqXqkW9O8sXuR4gXGszgS/6lIhkn8jxZi4tawSDNRh
StBYjALl25t2A83y8Sror492jBCzQtP7srYFIApjUkoJoZHjzBvQB34WabxqCgvf
bTUkMuhbH5zqVzUCohkAATwkilrJjryOj50gC7b1ZYMLvut78d/lebb2nw/25kwg
+bMIOcvYwCL+4hFp6zFKqsBYatO3Ebg6ntDLCICKBGcjw3CnKjR2JOM/8rRM+2FD
fvt5Bg9JzXYz9Pk80XnboaNMvGnFqFTMGUzbFotd2gpU0tzZXalU4T7g5DvG77iJ
n22Dnangx+NqrsI75NuCjdBawV6l5IKg8FkhL/2yLZFFSnc2KSjEScsMPP3usYFa
cWnCZ6LqlEJVNW4v8OfvuPATUNBIZMmpi+lfWojEDiooCYUrYebDEzB+U8yRmiHP
ECmfMaFLUjFuyI+EIMiymmUXqO9SAcH1C1bJNdP6UahpfMi+OvXTATtlyBptlpEg
OV59AgC/5ZDAV64XvFuef/GyhEsKrut5O8n7N8ivVqGtekJYdFXN0YShUGEALJLL
f1S9ZkSgDTqHLXqkXwuG6VZGLgRhY0SRZheXsalgoSb8GDHOWAqDHOm1LEGkEZN4
pxWXPSXWbSIX0tC3TU42TLOVKgovwABo47jkrzeTxZrSFBoxIDIVIuo2fcONgXyC
8+A0zOp2MFq7a8RuWEbtiO6p9IHmBvLcYixiAwwTOke3tnf+FJiKwj+t1T7iMPWc
ZuhA/evn8R7sg8bcVkte1jeUeDNAl60FWbsGfYvvVE1etJwxfCac4Wq6i1GhM4yu
oM3C9qG/hjOyOs8pR8dhwA6IuwfB+Hr3AXJ/EhZHjtlzpK3/kBdfdDrv7PAqksWB
w/eU/wGOLRb/s/rooqbAY0X/Dx7y7J18oCEH0GlEiMQ8iJJDbLJDKmMhRn7gXa0N
uVGMKbRcby3zoThJGWWPm0y1sS6RN5KGuWGaS1Dz3FIwr8iWAXeDzAtsBgyxQJpS
mWZGfL4ZOfKGUkqkmOd4pl7uZUg1bq2IpYw1dxyv36d5h7Ok33rQZlqQn1Hn9iLg
K9xnH3u/bN/zNyY415D4b6g2KOPK+q71CZYyu265h459xPXgPYCdjsUUrm9Pi3Ob
zv1GSBnVh0atox3j7fjy6sm9PeJHxqgvMfwlry5T6pJMITowcM3fEKZ9LNbvqNYy
tEoWq652FarbI9Nr8TMZcaVTMIbkMvkH43FA4N8Tw3GqP6f44UdXUVKXzlXKopDV
Mqpayi4eh5Ggyc8h5qvpJPDNViS7RdVpydjeSz5FmeRsTXJ1jY+GlrwarTraEOEW
OYSPKRVlpwpvozNNDqINYXsvNRxNnYvAxHIFL6GbgFJs0LyCMu5gM+4OEib1oGWi
QjqppAbWTtwW2yOZkwuKXDlvla3shoxHTZHYt0bhZIfbLe7TTAgXjlIpJdtcoNWG
d5eO/n0n/FHCtMZ4Hqh37V6Qrs9BmM4FzKOzjSCcpP5Ip3K5qpLwge0zOMZqb7Ck
I3wEXq/mCpTPSyc5nJPfsOWDN3Xf6VvI0v+Mc1RZFuMTY2NXXjxoPywptI4CE9uE
RiRyKVMFu+kLiEvxnO6m0nVMDmOGr3h9z9PpPQ2hvkP/UTPZHpDhiPWpDDZIDzpg
ezjmxEhzWMKhK02X6BgK+ok13O48erMWvt3sNkoez45Xq+iPHKcfU/0I6g5g0kcK
AGpGcVKAOQrDiwUJ0MD6ZXmO+Hc0yf+pwA/K4FrDpwoT+laQqUwv6Fg+lh2rPbSd
DF3A3t2v7RePKvjVxX0pDl3k/QyJ2GBXwgRXMt/7UhZvZQ6Ov3TEJlKPW2Z0wzXn
ufWLBUdLS/saUYY2a4Nja9DRjn57+g8rhK7W6Ng9AgJrtNK02HqhTK5C7aCinl/R
AV9XndUOpigZ82HHOKa1RDDJkwWtaYZobUXWWPFZzbTLkQBS68enyhAg8vX0vYqK
eJwEg4Xl3gXkW9y5HzWOGqNDZPKkIwy819DW09/FQUky4gvmJPPQJB+XtCEYjYhC
kS4KJdIcWzl14XKMZIF8CE32V0MGpa3qGVtz276cAz8J/k9aw/5VK5ygrBjr1ilX
NS/iGk+yRVjZDkJ+pyXnLjMsXgHgtbCAj4QtUTG1tUPmb1CLzEa5ZFDGEyySJb7V
UOghiyYdoQzTXEJP/xI+R6zjLeg7PC00oEFzTcxDK5BK6dBITkizsal44hes9V3G
vl6KWJXMdMHbNWBMWbOVji9W2A3zUxGqtaAoqhjZYTC3Vn/xi+EN3a3Cs1uV1Bcu
iCfWy59n8dmG8yY1rvdUOCLG3gtXw5Z1YcqX3AnpeNs1RUyRKFcQeVVAsnArWbHP
RPZAhEVl38waPcStw32klxvucfXaLTC1/YLnaZITWp5OVXJJkB2sFqGZl4I5ro1C
7+Y8rgsboVV9rYpBK2lmlrjVIr+0bxjRCqLFf51pxB4NvAfRS/Hp3+yGOkQqRVNL
MNA/SeL1IEjGX8l4qE3jkFDJBNls0gQXE9VUOpm9K8+IL0mJ1IwS6B2E95Mlh3ZX
oKpfJaLiuaLd88nKrqm5L+PjOe7G8G5VVhKJzr9ZwK9MeV8PQgUs8oan9JaO0dPO
1g1/pBRzGJ94DPHEEgw36F721QEsWhootunqOxq0JLY/2d2aszDsuOopqnul27II
h5of622UhRTj8D1qFkzgH/dGnVtVBRDcBGwL9SK+VnrYOk4yN20czuufQ345MMwg
WY2IjCeSNBMpf22eB7UkLNploz5/bwzuguAAjLqrcA+3uZ6jT4air8Qy9nc2GxqY
NLrE59cM+chbgkueWAzdFnuKV2mj1jzHNebRfeRo41d3/7vPDVZTnEgsaDs2xljL
ps9y8PjxTRRWPPhJp9Btmu4zWMwzGTZWWfgv7zM7oSBSpYTCilQeYeGaB9ftk3D1
SdSLXl27KbI9vJjAf93Nx67V/wKlSoEK4n4wQFmKnbKHev4YTWaHmgo7MZu6vWOr
7tYQR1loVEFiwrUiex3ktHnKtS57odQqdwUTj8qhXrDdRLFxLxGmKQQkJQF5lJqx
4cIeewwAIvkw8xVwzVYQ9eLdoCbBp4EYoa3w1dDGqFH93pN2RFp88iLiK8+xv7On
0mp1yWX8/RzdBkL3HwLd21DuaVv6s7HAICXGZNOB4LyFpo6Lpl63GEo4ZOgmz6G3
fRGfIUFyUMy2Icqh/ybAlXMxKSSbZNAZpNzRqvkdf4qhHw70TPccLcXzxpFXjTwV
Sknwq/t9e2z+MxsoQvA8gcWZnnnWibXnSBvwC/bO/fU7jlR1Vvyx8Qkzss2d08Hb
/wPpsbo/ryi+P7GEahw/8OjHqjVW6RJR+jfSdIIS3eT1VZGRiYxUgvBDn4Ain7QD
RD840bzfRugvzQc9pj+xNhn6PdDGOy2I8fuyHhoTLqECvPSK2drp4f8JjEouNs9s
2yP8Xv0l0ABIQm5OtDdGRa3IWh+ajdtw0Ag5cKzdgat6aj7hMbVwNVvxxbVOYpAs
2bB3BxCTPQparanNsbWEKsV45obqFdkxmiseO4bYpmRojliL5zy7vGB9NpCA5uct
7puSornCV/HqC29i1bQUrl1kg7kS+vPD3DMTXv9OwifElI/ymmvdxGs0zH6GHD7a
eG2MrOn7tge2l9tCyZVt/fFiDCVRefg/at1il23FkV2e6OO2FZuzuNTlL+u92J7B
h/2LixdmY205nVbJ4TpqsI/0YDuj/SocBNQdnmvjOlWnLsMesOZNBY0OJCKZEEXb
zy+hB2kOqa4YHldyUJa8JCx+ZYTEvJyfDec3iXFuEoyhOfmcHpXPUeUMXx2+tbLx
55rE7fseu/viECIDslyxfcjT9jeIA3dCTC6/Pk0NRrGlxqBWrVBaj+cjhg423Zys
cuBVE/ROT3eV58mjwYGESR27GVQvVe8/WJWnJK78S2SAk5ypcCvAHrQt3Svw0/C+
hExNeRZQKp7y6hm75zFgyIi+mjR2GlZVBzX9pZ+saG5kp6rb/8WaaUNrLSu0QGCc
rxINeqq72krQTNzK7iXpw+Iky94v6Gmr07aCIMSbqCs6100eDFTxIOkzsCqBfSl2
Pvhx3OOrhE4TjxcCbEHR8YBRwPbJfQMnee2Hsx+1HN2Ke6xgkslPRJg2gV/vpTO3
vJuCRqQ5wFOou3glPnjw0xfSyiU4VEaad62TWSMKmOUAhFRLZXhUIYJI8GqsMZqE
a7uiED55la+uPihRW6pztdjNv6JSLpCQcGGEq5+eY3ybgO8L9R+WMeMvHqmaQfGL
tk0NhJUsLZakXSPYu9cd6UaYV4D331mQxytWunLXQuqMb31LSR2FAoaYPbHWRjQo
VetEtLQ0PTNQZi0Aj88z08Gj+eY2rYRUqy6puHptoCQKwplLc8iXflaW8SrLJrzl
DyZZRnfP2y9mLbirUvbWzu85r3V6oP55UGApJ4OXgepS/VOjYshq4qpzu/9IO3R8
VS1tL5xDD6SSzAzyNCZ28GVo+VUcaYm+Nhuq/cn4W5CECY92HvZCbYwez/zXm21i
a7/gYEQcX/J1cSSMlVjbrexsml9L4DRlKc+WInOMlpBh4N6+VL/GRrt1gnTrNZL2
QtgD1drPnLNWWfTaumTivRNICbnbQCxK1HUQNwOwR8hEBuUOUWlkeoLac7SlAaAh
bNL9ZymRpF3qDRHDQo5jjvR3ttnRF5boR6Fpp340sSXchT9lJVjQZhA5sNwFzLfi
rTvf9YCb/KWaKZ3oi++NQ7P7ccNtxUg94NaeW50m/vATU/RsbA/N1KHAPZSwyjBh
3zm8N8i6E+4vCoZSjuVBhUXiPqPuZjw3bCOePK1/gcXsR7bNe9TN6/S3hYKJdnSs
6nDqFidrN1aFukvmjxn0Q+5iT7twJ0bj08ThPlXdRiwc22IpQX3cAi9zcpKQMl+2
C6kaeO9nxb97CPT4uQ2tWrIJb/ORWX1hnFPECO12AB7WHFQ7PNxKBFkw5iBEQZJb
hVSsmqTEgzaBz2hyhNpVTP4toH+iC4s2CryiD9MEZ251Wd0KSQrNp1DU1rQYqXIZ
oxiToQQJuMIrTvDqd2/TzTXik2k0b53b3opOkGE/Ky/dEeptEx2lwG6W33cvXEcY
eobH1lyMfMhlClkS+wK0MukUK50hJHZWtRlOVLQtQiNtuo4l7yNCvuLODSuq78uL
0EHzZ6btHTgxorO1k2RWE9q0MIx+VqVakv1KiUo7sE3Gis7ai/AA2swYEezGqKII
R041v93O/WsnvzuzNP023zXO7vE8zMIuRqnoELW1N8IdyALUV0U1qMwq5//JL5dw
8QuVPLaFk4yBdQ3QG2aN3HfJBTXtfDf81H1qHQLlZhsa80cQ/mahUwxdkIdJemoh
buNRgIv84NopA65tEK3RfZDfzJvu35Uo9JPVAChEACqQY3V/RZfVCCqyT0r7UW0b
WgZVQzKDk6Bsgm74v1f4B9tmq7xF8mm94k4SqklD/ihQ12ED0iNgHPa8ZiTeiE1D
xzgyytiuR9Wt6eVCqUL82tzuy6S10gYmwIIChE+RlAlK43A1rFynnofZKitmuF+K
nRP49LFqgDser76foMSg33IG5rwng0i9ZCH1a3aIn/Cf+SyRHc0y47X3ptPC7V7L
P1A9gEAMfu4ucCE1gQL3VdI5zD7TIGlM1TqoOytPS4VafK5oDSDHDv2lR9X6RjNT
VMSWr+EIAZaAxX6AVCRVqWgVK/FQS1Bb1alHMOl7DNRBadzAR0kyupHKOEPZr3mS
/LwWZ33TQ9+iOvjb8heb6bttCgeky5p7bV/UKS7KU5K1jYpAf7jcC/d8Rht4NxMZ
466E57GX6bg08S0WozqUUNhKsZC3KTJY51cLaYJidsTOYG4cjouSJLHe0w4xK5M4
V3L7bAH5S/K1uszaz/hdu3CQlBgDPg2cpbSVLDf9RCGxBWFdVL3P+9wAj3KtJ2Of
4J6Vr5cRbxAjM+Vt9IQUxZiK1WZtI68YXeZV9aJPPBetpJoJZ1I5fcDMGf8gLFwr
88tjtpER211ksQq9VPZf+maRXnLqLIU0kb7MipXADHYfjcHoJjL3r6+yWx0U2Ocd
sVV5WmafErNv+1iXP23kVpXrnNh9sTH0jb4wfosffwnhW3i0orhuYTYobP3exDah
C3Ai6eNZTw4cXBXJt0YgIKMHAlYCxHY+jPCIPkOYZCK/Wts3LXxnu4e0DklF/1Pd
22l+CxGfDyWjy9ngoi0MHGaITNkFlHRb/kp1pFzI8yFAGHCtaueplc1ytHGXdYa5
uM824GnHZU+TQx9AZxD/LNZ8fGyPd1FjJQUmsGtkMJ96ClGOP1WDZUGyOus6g5mO
4EReOGH9t039ZCDrD4vRUkkyPh/DbyazZ9g9JSNjSOvhov8BOAck4u/nYNHlpit2
/v5JdwKZKucONRbowZzDM0AJtuNj98BeliXUJGxL4Y8uSPvbhY6Zb7XmgJLp5lY4
C1J7klR5Cf4Vs6u8S3BFRNXWvmdrZYVX+boU4z6to6T5bK4gYIglJeVtDIlCoEID
0daOH0j4w7qS5nq1NLFKJkFe+oclhaZsYBdXg7Zw0eMgtDWuPboppv9CDBI94YoP
oJOAL0snkzJqc3tqwmL947M8PFGxIG3LuWstN39nzXn9uEMsSeRueXasgWf1K7yx
o6NcoSsGvz/KVSq0aGXrNAEKqI0bv5DOqKIooLHnV9jcRxFhgcsWPeY9hXT1qPBV
3w7H0a0ivjznkW4z3JB2ZejS20PwBCGWbcNhCfcQCL4iOtJBgccRS4Xs4d0lAM8z
UYeBLEZXyVxDh3sFAJdRskzrGxrvhOo8onAY6YaT7HoZiCzMUPZ+U9LY0OKSXlmO
HnbLC0okI3LuLp0fgJBzjkwMWfAHNnq+cBuajWQfD58Q/5lwV9bkj5j0zaoOjnxl
iDRldIICMNiMEQe5dFi+wq8GwO3EJeISzv73rR7ABxlubgsOiJL/YCMRQXAXMgpx
0GkgqzrD+V3tiHhy6HgCN5PwfQOb/aApABWWOSiczZCtgzqeYL+A3V5recYlaVEC
s5RJYXQe7qBwLKKd8WEh/58oz0Q4oBYRf6PoInys9GObQ5/GVWh8kJ+DcfYjqsVl
hEqNO1KQM+E7ybZlyXwkgHasiFwZP5wlskqwE0J0zt9RSOzMgzVZWqa+l83vWo9r
5jKnMxJYjSnwizEDnsdi5HoOZxjA98QN7czZ9CtBlfKLBSmXGps1mab+qAbmUEut
ej5oEEp9fjjgEIep6S2AgN/mYyby2De45DJoIuqWWYr3Lc3pw5haewLuwlSBrlUk
+fDr3MSXsmmHILCxJCV7QsuwZSaJdga8+3x6aiGvD6CAXxzEihLCySNJYO66C3ga
DV/3s/ogeqWaxbM5g7hEgjcZftFu6G5AsJl2tvGrVoW52b/F+wpR0CIMGWb0Ko9T
cGad1vKKXGJCFQ57uun/jomcFamTpsSUiqrj+DpsTHH24SZnAXbDKA3OmyXyU6Ag
+GPKiQn+q8B3wmiPITouBjOVPx5I5UCLTaldZrdj3Y9HWPUVSrftecbHJoSxJTGo
FYkO5YHGk46LB55Z5P8QuXXjkzzUdQyxw11EXR4gJJ28BMqeatG3mDumYoFAI54K
319UryHxeau8IrZXiESMGAyqf5Ii7ZeUuch72GbzTiC+bWNuwHnuqyjMdm0Zp00s
KFMebx9GgSFNBv9yD0GDb2CoYrMROxXBDEDEArkfJIGTGjnmr2kh73nKg34mGdEx
Qu1ZccwR/x4ov9FY2M0Xk9HKNxlOdjJvV5BqOyFVWEPkfSqtWO4OkE96y7BsZN67
2a8ZVODyu5gRXIPOXAiSct0MzaRggIGVn9voJfQnom06Pa9qiKqoIhPHHz/JPdDP
XWlVr1LycjxJ5uPwMQVd/mVukpVN6WiUWe+JqcqQgSrms3olGTgtjnIAq1Ix918A
W3FlwFDvQD9pHvxnKt8Pb1SB95u8ePZDkPbZW4SRdAE3AE+8a1KHpQfEUr94lP+L
B+R66A9h3tGevTFxImwOiVpVZwTxglb0U2r935it5Xlm3K9SNzwyGdqsOqz9wTeu
NRL4d+rpE+eHgRp+1DLCTeqi7pkRekhPtEANJ5cH/45yngjzdbWWNH4Edi7DjdLT
hJG7MblgYvP/5L/+ozV7JIGFgYyaGnm1yCz6qcrZn6Ya8cowHs8PUKVph0HFk+q3
HtwBeKb4X8Ff5rq5FJpZQHUepj0XLtSZq5sNIJo5sOzCf9PlZIAEkEJzOSxGnpF5
aYfzUP2aipcRHjCuMfzKTuokBqDzJSnQXPXkz1Eu93ZiOjW96FMb3OZRjVXrKxjj
W+Gshi+8F4SmLlRO8xc8S7/XrYMnxn+eih2zihmBNaitNf7OxiTaehvvLYooRIU3
7AAJUspw4w02rUhQ7voB4NKBGQGdceAOF1o2D+r/KygjNUxpzUp1IZZ+41xFRjYU
+ORi1O2n9FCz7m8urdPwxRrIz1pMb7NWN3maIOW6lQkY31fupjIT1gPKtQRpmv9I
8jJGWeVrMtmuH6/i9liVG2OpHPRvA2jTuG7X0FvfDTmPwVoj2gYsoisXeeVk22Wp
C8iulFqmoJNbuofUAfbt0O4jI/EipelhMGOJ5J4iN4p81BG0Ui5gKHDLqNcf8aX3
c/JNm3D6RVESWYZWPMcwIEjZ4AS9UNJ9GNKgCe/Iq691LYS0hmXdgqAAefBs5Jwm
qY5XweTdQKWEL5XwamaZIwyCAe3SLRYOi92OiAGJc3AYanEnkHzo2MMD0KUPGHzh
ZJiHm/uSMNx1B2DKKCZMtV1BDEyMEzyHG7FC9ad3DScbMjJq4zNgIhDOJ/JK+Ix7
jcy125tjS8i12GCbbPmtEoXh4KBZGcxXgi1z/TBSimSNkXgY3kU277PdBsArfAD+
WFbMnmYSjaa4OerB/nP/LjGeNfRQ+pUvW2SdMwpLIX5wKng/OaR5GRuqvWRqf0Ec
siZsTzdRLpmkCAZWxG9fgYCgQ0XhYy+XKI0WoKCRJ2b2zukFciFGLBXGbJsWQ2v0
nmBnM6AjUd+JHaKZ0MZ5PRdZnPoPvbwlrV1nMzIzMIdXgtNZXyXBXNjR5lqQnuJW
+d0j9oIAj6Ar88uE5iO/gHQxvjh1F+WdlbFEysy1J7t4dS+zjw63iFed2/FgUTxH
SRG9WdvmVO5vseeS+SfjNg4c5o0rXrJwBYk/vY0feFLv/lYahwjqXM+HPnLfeg+V
7xYwEcTuzboyvodZ0u+9ZGrf5F0B4KWhG55UJd2PLbYfWAjavBaAtWZ0AcTftJco
MA3IvYWph9CZGg6RDu+ApnbnGv1xiBDLS0SqNAG3qswef6dnhIMN3W4kiFEJR3xX
YnYgdR7w/6+Gj6QPJWQA+rF4jjo3K3LUe+TDeLdH/KGVj+fZzEX7zveY+X8DxInv
T5rUQfT28baMjJARB8f/+MIJEN8IjOpBsrWtd2Tho/z8y32MnyiEYXUG6780VtlN
wOUSiqB0bwmwKEvQiS8Ztom5fTt6OEnMdk3abKce9QtN8kcG38sB86qNam9OZ86W
EPdtJCuYXMa31q+1OI+lJP+UtU+yXfrYfqaaew1Cn+dsndokwVq2m+TOtem2LR8d
MkVOFddk2QhAP3uPVkxo9hZ4UEYgeuVpEFc/Ia1bqugQ3EXbEK+JxcN9llszhdOQ
VtFYolOAYRm3emBjPptJLRBqZDCrgR9R1rxzvoWhYn8O/RTcHvohDT1B4RBdU0v9
3R54wEcRhhIo5k3UyHn9AknZdcIQm/bIJl60ZIYuNaLoiMGZJIF55Bvkk/IIX0TD
ktY6Y+DSF4FbPCGSsGWCtsgPP6HuzrphD0sZK8lkXpgumOT9XmKep2XVZjOt8HfW
PSP6NEY+kQq84KaS1Fsuwb8VfYBneiYF/rVBXSWry1exHTpPu93Aq1nngYUT77RO
8sKvCPEm2R62+xlrzNaDidpiIfhacorqqqxluZBwBkAidjVmiRQ7cvcoiacqlQKE
PpsEMEwN2GR6YYlEoeXKvMhsSvCiLoNt79r0qzkehyD74ASHecaxKneL9yXrD4aI
jC3SFotfTrmc+LlEofXWr122Mr+1/10nJZ2s0qse/NkFXwipMXOsRXjuW5C/wcpE
rogDYgFfAHpwXYqIkJ0ehGb0nMESLxuiWfcJnbPB7Uvwl/G5mOerCydTVWgXa5O7
KR+eFlw5+EXUaJZc1BBWUuPNiATgTthubKfvD4ujWQOUNU9iXAr1e1Ku4/el6LDh
XU+YdZsHicBrHVO5wCz1UNT3KlOVleH+r995nRahOs9g1bHvZ65Lk+03h5xdviKn
BwFAMVSkronlc4hri/2XDDJ+1WuBWqWZ6GpFod/o9CehqFS+O5mOQ21gq33YPJxF
NaIj/to4lK7qWiC2ot2dapggZ6U+WOfE2KRIA/pDJu8hoebquOcZoTY0ddv0H7T3
8vSmGnc9o8OxiTm+vTmA6LOYjo4b1oG5Gjc+GDA/FqQvsbt38ELe07bnUhK2gYui
b8tpBak0v8DloHaEnqViFJsTwty+ja8ylawA/c5+w85OgcpYxHiuXDrNWnRZ6+Cy
h6GnA2S/fdTBQ18myh9H4ggk/clBNZ1osi/VAa4J7Y3eeS5GBxnoR9yGtnyIdSlC
BLxjH0WbDfdaRUk8+tNehulf1Rb8vJ2n5cQw9OW1oZIBX8z3jAQ8aMRlQthZ5N4E
HMWojF34Jicl2j5dGSsbCVIoJXFa0TDYZQjGLHzJXv2/SmzWbVc/xd4OUn/u2jdk
nkFu2HEG/uUncPs9aKzMIVRO6H0ZfA4xrj6XTFXGDC8QGcWjswTnuT5AMIHqqxSQ
k5528GbIlTjd6tHGF6sJIjozrClBwtwJrnLTFjGhN0DeSHeZw0LbaRkwrWI/1NFw
pm5qVW4NRlRW3PSCAYVyky41TAiOVu55mApoYeb7mcT47OIyChVCTel8J3lMj4Hu
D+7XfpeX/qjRYSxXVagE0/MO36B1JNxkoKSMZgpBD5s7rDlEI+RXlj8R3KYPXoUD
MWl4ncl8Y8PyNOVd/wEZ+IgK6PWRc5NM8exRvyTYU2RZYp/mfwxfciBW1EzjH5os
XgsYpS0KPGN6ikqZP17LqD9Dv8mo4OWMk+lHxygO+8dzJpexZuXHbMpgcHEb483P
tFS7hIx2letnTO5cC+EOJWhaql/Dp97B9ebwEp+J7RH33mWJvQ+Lj96Tx/Y6pUjL
fG9uLVReC/yTxzfo9FosLK0XT5/uU+jNbwswUCj/2o/C3aLmRlQQTh4GvRhL042o
VKBgMIXMC37A5alAq8KvNcPlR8DKtYTgU12Or7+AUvb5faGX3d1jcbX/qFlh04zs
qBtcyPU+gAu1cjY5jw1TLcpgLPoJpticsNW/INDlniIx7bprEVP+oSeUMGo+xZ+W
WJ5F3P2M/4IINHEf6/kSdZfisgjRBvmyMwYOn0zQELjAnMokxWscpp8EEo/ve8cV
lKOK3xTEd6OtYIP7pGhIzVwlemFwlM73vbiLYbg+0Tr3MmAgJjI1N1aud4DLj7w9
2+KXvvArg7R6guj9QsyCCJgFD/CfHfR/AJdNBdRa4KMTzji0WJ34MTbnyUPQ7tC3
Pf07haec1CMlgbDIGoDLKKGgwrqWcTgoi3IFzjTCKfJ7mmXPy7vD8kQk30UnOX9t
Kf9hwAKC960Ba0ocg1ewhMdYYqvNBwHkhJULV9DyTq3ZkZaDFbtSHB0zWWlywLZJ
wRBHGzzbXJpFDyWx7IQM5/fqGGY0mvS11wVwnZvBiW+EXtpcThIegADoy2J5xOvZ
olBagwuixRNUEPUhodJvMR5HZ/FiGLhSFYQh7ZN8RJyOgISHLKPnhXm5q7oYg9yn
NbiItAH0lHkFKcMw/6KzjcX0UuQMooD0sPjL4cu6JoS5gchuGhlM+/RoGvHgbKn8
QXGlI+smKc7NDALWw7CGGxUujes3wKQyRn5+m8JtWUh8l2hTZKnHsYLtSI9lNYP7
m3a12cURrAYUk0IblLmX4BBBV0gRPcYmC+O4+xY+UebfCEqIgE9yg0uK4ObluG3s
RovmVsUeE+/NNCLLLRAFfYqbe5wEdGW8FZnpBu5QB/ppruQCCfHDStvi40istn8p
JArB7JkKhFqot7WwRKZz7WEpd3OcCXor5K2Y/srNSMOE/o/Eyil1zCwLsFGb1ytt
x/h7jCYPEAsdqa0v9TK9E0WE1f53PC+5upjHNbZwlTHfgo+7dyCMeEfPDOj3Auaq
mh/QPoQsqUe1CAofg/yE6Cj6wBbQxxbMQ7MStHk2NdwHGMXqOzjEmkd3S36airzO
y1CuU7C+goEFaAEaKvgigiSa9K44Smdj38YsEz9Wxq9WhV59StItbebhT3YvwkJe
j6WMQ0qVS9uXiqEax4HVmUVMAzuHm3cEh5vBSTCJKMrsD3A+RQSAo1yvjVmUWrAw
NUQLK9mshvBQsN+vdPTE6pnee91ec5cSZV5uZxb9jVddLOAm/JRSUlVKXQhDF00E
ZXiYy57S+WKxF3LIHFnOob7O8RBljS/XmygYhq36DLy5ENHJbFxzBI+WXPFO8IeD
XSGLM8dIDzaPUT33IqOuVmjeoPptFWKUWoCLyM2L+A6wJdTvrXudXA/YExXrfDoL
6V2oWdngeW+1NxB5Y8H4I7y1owKOhbWzJ3PziOW2zOuFBmUtks3OuhmuN5A9tjac
RJQHie278BvLuZUGoN8iwL6X0hJi4lEjolO80McZWiWDhr72jYgzqgomSBRReuUb
ralecKhJoL/Q34LcLkTFysmXyoMv4B14AOdIelIVC01TT8t1OZv7ty6hTc4U7Xl7
mAozRdW3l5e7a9ykOBoDP2lmihXf+NX0PH377QQaYtdSGsFjv+4Z2BkIZkQytn/H
PI/FkzwDlEuicc5nryaXpBChfccJ7f+wrcxbeP71AD7nv91NzJPuGttzp/NbCt+q
BnOEuyrofiS4aTYpQyZfIVV06Vqzu9CDuFnIKbTbqP9GIMY5cmX6v88M0cX4I61w
jFR7QW9LhauVjNIJ0Q3aLPDoh/4OfyTJbt3mCVZfqn6SHsvHvh0rcAErN7UtMabe
GNrDJfebMw7shEMbYx8V4mVzPS/1PKKY9tEu6UhN6ORfd4kaFnXY5IK8u3KkPzOe
7Cai37g6j5h3Goo/JSiOJxx00CtvbiLPhwD/W9YSRPpZ6VERIkxv0USNEJSnty6u
d2N9KG7IMy+7uRSwyXrtQO9JpQbZYlrvgt7Yuz9s7BTIk4q6cVzOl6FoonywQGJu
2+esp2vMO0hlR1dG8e1LGL0QVlvIAShq2AYfl2WrkuIt3PmV8IOG92gjCnYQQUpd
pT1z12L5NKbVPo7NyH5O8vfNIJIxwHjae00bWHAAm4qD8m/SEBNS5SK67ffi8IS+
9kROvIDx43GCzvcMtIqJSW6W98p+BQS+co8ZmIIUVhg8nuZnhuWD+CLdNbrvwU8o
nsr+RkSWL4QeCLE8zhxo3XSLzhiOBVKZfF/RS1Mhvz8eNCPnLhZNzZJG4bzyIQk4
IjKwh/XDwDiNctRlKaAnsOxF/FqNAa7G26RekMjwe6DnRX3goRD2+6Z2Lfu9jUqH
aFK/5nZLADYUaIeneDdDbe4YszFFbZLtJvuMWekJeWbwvaIocTI2iURvGUAkcHsQ
vdkxpLE/LVBGceIyscOE2Csb7xW1EtASdGfJcZw+Jc543Yi5jGJxvZu7v/JrxjHK
W1kqmLWVAUdieIfW8VDmNI8E2YiuY6UfOrJ7jyPEA9M31X4bvIXdA9nDMV0e+8DC
Qnjslmy8JVwQnC/AnjdkM2ePevmJ+1sMZYZoIdPp1hxzkg3iN3RdawM3u3wnrpzF
lCcqod57k9Xmb/f4+qvdEyiBfGSxEvAzEqxkRG0RHq0IVsxeMpEVXncaChtZnNfJ
V2czcwC7EWSVLYbnzi1Epg9g2ZSvPVyHaSAN2Q3PkzbVIUwXfpIRuCiKZAa2f5pJ
wZr2p6Vm42jpYfOQtfxRr0Ez0C1fZ0JdLQIzvrFy1SmsKnegwMMduDFAoMejYw01
E2ydYR/PdP3KQAbKJdQ5Nl6Re99ag5NgaqZxRUXZXPnYECGYuQ5/VKN/onZoO2W3
0lkpDlrd0fE/3pPHvAKpAjfTU4X8EOSgFb62flT8woWSFrhLVoj5zX+ZUtE5A+6o
kxGtuiXbexBKsvZ8Rb/nCjVhR9iYxOW6Zp+6tYFTgFmvmW9fml8C2sczfms7U8mQ
/zqwR7bdkO0J2rUMH2ciOQvk9CgBbFVFkuW0Dv16kdRgp+dHG/2fqK5+Y0iokIjQ
Zo3w3tnzS3NeOU+EfeBM1k++MM5SuBm77xkjGK24XkbfSI4bTscALP9be2H1uNf3
XxlK5+xL7SSARjC0eq7fK0VOGqah1Na5OACDECFyJ8j7m3BGcYz4Hz6iamsCL4N7
nDFvVmhyVSueDd00wpdeP7R7F65x1Q0WSp2/3BSU5MaqPrSqIHqIbqhYGX0LgshC
k6nBRHHz6ifwCiR0ao5wqeEDleeHXg43isqqFZz96NBtqlnc5yHJRjtuDvo6pqy7
/9c2gJaPwSc16OVFxd9RnnZMG5tRoxVnrgMjBsC8/TXZBLF518L/U+hmqwMgldM7
rbqRMzq6aKJ+zC7EFqWeLCZ8hBITCLlLNbeANW3DoNC3BoX3MHal9MG+8RG1mXRg
Nci86y3Jxn5Zp9QBgWHHM+2JUI81BcatpGgGBpByZ3PcDAIN03og43OIRQeidc5U
d3ElPqszWObRKOiv3v3dXXjll2FmkgbIqYP5Mcq7Bim9V4KQhBqak80XnXGHJs7g
etLzyUTmvGsD2YRKBRYy/UoF/gwaWmc/qUnu6GTrVHl0IJLpV9N9V0X8zzVcOMc7
FeYp7SVAWOtWSzFCp2/QBJX8EGvMIzgpdRU03ble9MPnlwUVOnLbfulsWeuQXsLm
1CNrdodnv1+hbmyWOEvFvun3onq7VV7dREOcCHzZYt5BgvdKuHMtpteIblckRdUw
GeUrncPGjwAlSKQQLW9PjZijMpOn/3b4jPBNTIG6hCAihd7d6Vu6Tuph+8kfdTBk
pAgE8GgY8X1b6GdtVGtPLZEWqa+PTepOwZahSP28O6n5DPhD8Nk6k3JFgQ6hW9GR
KJpdKwXd740a5Tn6SWBoBrSa9wmslQJumxy6tLbCNfNQ+ZrR13NyuUBE9o497dDk
MUJP9cHihvqWebln73we45i3y5Bb3mmzTkFfEnKLE126hdONNi2OlZ9S6Fz8X/E8
FQSl1/I91lC63Vtc5+IWklyO8W/E7z4ojsnCXJLHKm9Z1u/I3WwRGF5wRUzwwAWg
Ek0PWYQQDoZlRBs927eGa3tUba+Fz6pB8PqQh5uFbwasAxMl4VvtqKe60SgqVqjp
E2Gnjcnfs9e28arjIPTbyTFWFFZXJBGWCn/gxA08PD4EZflK+lJKOvfVrvnSdgn2
1EHxihBRTWutMeTI0KpJ5VR0h3jOU1B2Ys19zxHPdw3eXrTGRJITgMie2a1f7TSl
2Ib4YFPJnRZ9Hp5mcLDzPh9/0Lgq6VAYiGN27g3D6168TiWZ/j9vSq4eUNW1qkff
6Kib/4XdFfHmLSWlKbcyF0IDtMP9wJPrcrA0bBWqiZTM7k+u+HaCRqlyoRfGB8sD
x8Z+9/dhEfu6PdAgl6Jl/2nUvIWsgPnMevzekdIxX0j/s57AQgcsYogGePd8vxQU
CNZdgNiuVcSD2s1IcmRIQA6UJit37lYZCxfoix0C/+/QDBDupvAbxjyXinWPZ1I/
njEjBp+K08oM3m4pa4tcfUuoBKwxYJ9l8y666JTc5K10iKAd9RSNGBlk3gF6ESJF
/rVDOSZnl1MGz/rRMh4+uOeBmj9ZNDEZ2PrfTcNG/iIoBvqpow0roOQP3nc3bkxI
PsuzZByvpS8+auJywnd3GbHaOAdgG7E8KvjOfF18T47uwnCSqAqOoCoYYsAl//BE
r52C4CjrO+puuCw7NIZbkGuYZfeAP0W5/C/PXoHn9vHb7ODjKgIcBuTq+Hjyz83e
EoDui78TY7WTePKxkZea+Vp3UralGIBwt4mPyTwmn/S8iIwnUmNOkAGJMcJ5y/WQ
8cSkqcwV49/MiOx+alqXrZ6I31deGRSd00jPL487nEDrP2c7T0mKsKI2ItJw8pow
p0E9fC8970926osXmBI+zIpwlFA3V3uvuX0Gt4HG5d0JFfB0Ge4luu1PYL9VT7R6
xyOeOyJlYc141Xv8J188Y5422rRHqhDjgMYB2UBLgsjF+/fQ2XZ8sZ4L4ns0tUOd
cYlVRnn6qvTCBZiN8vv6uM5x1eIbWBz43bGrwE0OXB6/nig5xy/Ws0u1h55k8V9F
AiZwSd0lpNeXuy/akomo2A9dsd2AmEgvviDAKqlUW9yalZhywHuR306fT3tlFuw6
whlVI2GFkFmqVNpZSbtEun6pY8h8kPXPPfs8R4I9e3cxMP5GRwGKZKtPR8hBii/t
9IcCYLUhkDgIpRyRPStoiNdM37l3U+z31F6B+1BpvxrChQdf8mqN15Iai0DHquI6
NmLt7CAcSJvDOH9f+Ie3kj/+fxU4pr7AoNykZLcay3Niq+PrdD40C8Q72oO+/wgb
epiFzDgA5OqGZvbO62Ty45DxW8fkbMJOVJ0/K8coD1iWa4NuI/7GjvS3/n72vhLv
2UGrBkMUi7exDzTaiFjlCO35G+rczo5PQpzTtEx/EVAeLuvFuSA85/w9sKSRgmlJ
UWPUvwqag2npD69NvxpaUcpMcZtNM6HZokGCb7dDIivGHbfwSQYK8Xsh30t+dfXI
Beua7CPd+6+fzuo5zhWNu2rsPQeImV52mrZEGCzu/8W4yHj1gbBDkRILAs+sZZmM
38u8/qmuic5OAP7/lAMNnZ3NNNVcESSOEF9oyjElLnAWGrauBOJbfTW4CREkdqAC
g8SwkZyi+Bd4gCe6BSZjWNCYk+QaKDTrWeqRWT/dfWxC4WpUDqDnx6GLSyIpG0Hh
v4gXEy+uPKlUM/eupMHcN7nXXTGGKv2zz2SjOMMuXMRFtfMLTqOActXfcLf0ejOg
DSKXzVGA2yg/YoLtoUDJm5UlxmWGIoUg60/j+quiZRxr3viIf8jBuVZByf99PaNF
Q859IXk/kv4GY2gxARzTtWqRH8kipowNLV9+mJHvhEBLKGYWdmrEAdsjiNzLBxUQ
j6Fp/cEg8Xz44r6nNuCIoONpwRXSQxdamYK1PCS4uCQoS6Bz/m8Qr/TpMDNQ5V00
fWZ9ikL0BKsiLoLMeqU2mzALCE5WN8hUgqBqHp4MUu54TdVUjExPDNzopJdQKqKv
a1LDNdsocatZ7inMY+AeyvtjV6wEgfFiXyFlXM4PqV1m6/dXJ3558d/zbk78/s7k
hhjOFde7QPsu3/bo5+NPRMu9vgCzdYDrBWT34X1ma/JYdWkXBqhi3R2PD5DY7xxg
QDKrsP0lN8Hynupu+pb24tKPizdja7q+emeUOC3yLjTCBmEAuMF65zghydDlkVQn
eNnufIBCxdPZ04uMG/d3rB25SnGXlwE2yGKVY55OmgSkUeZpgGd4aXS6NC/y5WHs
6ZTqwt50+JBJDeya4J6Cw8cFu8Kq6B92J5XXWYJvXH3RI5M8CijeC5LOjhX4xCEW
1rs6va6cgJlbbYFnlHtHlWgH5LrAC7/5P2rM9D18WTAWmCteTJIh7zVeivJOQB+s
oRSx4dZkXbozxr9NLIfRWjlg3cWRVAvDn7VPc8x6MpCuzUwDyoDrJl9x4ZppyQdo
y+pbQhsTZgOt2ifkH0DJANPmVTDQYSQ2M8aeiDisxHMXHrymW+WLYCDpjvdO9E2V
Qg4qqCVOOm18zxxvh7KGVR9uVBnW7VqEo2lAUiPf5wZrHnOdiHRKTsutJJ6MgoOs
UqfduI9I399H0JwQ0qmbLFmCePqEZszKRMdpIAki3gJlvNNvuWGIbTCOcjsmzAMi
DAw+Mr3CQSD3ubXIw015ug/UZwaXU2qWXlMVgqvrBiA3MP/a6Tp5DwaQKqz69JN8
TWortrX7+u/VpX2buFe8ITroPMcjcjD6MStte19zJVupCKHc3uEMf0V//nS3Y8O9
D1JC0Je6WeK7d6Peams08V5ClQOGDKjxfrJiDmy9ZUmUBCf8A/jxT2YwudMQafgT
+TkSG4XsTEwt5Nrf+qLvfZSPwtP9UaqeJW7m1WTSjnwN+IX+Et7gikhweW7Co0av
VGI3QtRGVJdNwH9aarFlYKxL0V2zQSjkgnQFHP7HsYkQ4PayA/0mBascJyOFZ98o
FR/hYKRBYQlI3SQ1Cii7hHj38AH8Nt1feC1TXIlD49HJP8Xj8g0Adz62KxSTstT9
nzvITeq5LRAdiiHa9KVEinHyMNBSOoKpjB2dTvEDJfm9mzzEjNrtSJXEpdkttmdq
iek7Wz5cZezc/3zflZy50YCiNN5PmtL953EqWuUT08YwDv78vNgPYqT57KSfbiXB
5SliJQVvl0nmNKMfZ/t0y7etQFd8RChaXQioJV/oh1Ab89UY1jVF1+OcmhIrVpIB
K4WjeSHkwEXZ8ihunCWBdWYg8co6KTZ5ZzLiLKvsv7EM/8z+DrmYCv4I30wAWfz9
DIQcS3pAFEyN75/MfO7FJ9n3HQ/bd17Sv/BOcHZt78PbyKyFeNemZKrcz8EhuzTK
1/kq9/WLohKr0c75F85Fk2zcYx8TuLDdNwHQu5DFwQjj3X0zxFP05/7NKC3d70cK
vznpvY/Gc04lHLSpQaS+1K53kRJ4OtKxW8kt/ialgXhcQTcRDDZAasyKa32sMjku
xlkeZAEDdDmgNUZc3wnrDMbC4QkdPDdSia6b1/AJJ/1VYx/92B4U09qypICL4F0L
r6jQJaFUxjbbHNH+EPCouEs3tGiFxUojWEDbu+sRQR5Az23pSAszEB1E7ko0psBs
Dm8fANhTatY7lBOjMdUimWqK686IWNz8hb8XerBRapyolxyx1bl1xatVH2OLAw51
BTborZbH+Qui1yjNktgngkAtE17TeKDFgPBC+qJ1eLgPlLHbu+5Vdqtceh10eNux
MbGFSXhZx4VFyXaxxkEYW4KxCLJ3ttTq2Li2Sf7xTGLGtPLKQM5Vh+zJDc9VqgwS
hx5rpkWxhao2g7sy4VLDV1zZP3Lzk7mKnr8db4ADyIxp1rXbF9rcWXys/l5dmDT0
pFjO++ZCbCDO/r+jmsJaP/pGZlsr4+U+m/1x4LMsaZ9FuQMUcb/vQsR63dkYdHi0
Si7UcHeatQIGRq9T+HDc724JfQFag/KNo1cdwKd13ZxwXDJRY61JYCIUggtlaHTn
yZHMeuBMdU0dpPpVa9mcTI4tp7VNRs9Jt8dGHlhrqt55sO3hFLzDI5MD3/qoUm9x
SD1paqODccRj5It2tiuHzu5r9NkX23ADQb5z4SwN1W5dtjKuQOVrmL8wsJWivAZ9
RPYuoIEYm+NgjHahcQWx4ay6toPVMz6lFpOGoCtI85xzh0gQnpdm5k5NEGpseEUe
8RT9r319VWO2+/UWmc4pvqCxbCqtW1jLXEgce2RvY1uXXztW4lf/HMfxpPkAoVX1
uM0/XPOp8D0cyTnEDyGk19wQxqdPGdLnPuaQGD6c/YvumASiuCLEopgkKgkgpUwS
MhBb7abTrrkcczTrAdv2LUwUSALTzbiUC+F4tTrT1PoYzWg1lUzMDIat/0Se8svV
A3mdAA1LuAl9/IBBBEsNHoF4P0wc+kJ4gQBRzFom0Zad5b0p9pef0TvngrxKH0SP
UyT1jHxpiES2Xjr9WhnHdSrwiNR9vwnzNBK19/AYRN6/hYFplF3aLSeNg9lLROps
kL8Q4glyJ+rz6qV6ZZK/+GtejprmDQqcpfZiiBMWCUSfVbdxZGmPcdMXi1qQphkf
QoLIFKlCPMiswExMJx64SG9Y1d3ld14eRx6LPWwUa4bZZ78/2J1B0kVvVpZYZMgV
OTA1yNn5Cc4uIPSZfibiCG54t2zmza/Ec0lmZf1lqTS8jgkNcm6FuAwCQcq7fizS
l3r6Mq+1ozhiSK+lAQjwRdvrPt21rUra2c9+SkzGgi0TaEBgI8N8wEvQgzbUxe5O
pfld733A75HPJ7NBAy6DcBtPslB302IQhBRx087pRM/4DKZoWup9S+oG9Epl/A7s
xfHNsvdxlbIkfi/GlqPVKL2caIT9jsbOvQUmrIle3T/IzcnEd7Yog4P1g34MlJUN
f4FiL8LUG9tQSeOnptA42b5mBO55BWU+Ek6C+4YaGzpBSDAe/K6QtZQYxA4CObpf
UDHc9R4AzJzq4v0JhH9yhNo/BMex4CIaU/uaZ6joAi/I43gcJ9rXDBw3IhFPrUYt
GRDDVnE75WpfKmfQPB5exvfw8osHOPd1V2vy3KCBgxPQohR2LVMXiFkIs9wfqQQX
kjocpi6T2GE7HJLRGj7MsjUontE7idHsVhPH08/G8eNHLUEMpCDRww+wkGII0xYc
TgsF4mtFgOuFFoAYuPiDreb0suvQ0zLYUiftKDG6fyFPXMsXA8lcKmBVobwCMtUF
zKV/xmHL3vF0LRx1eii7ruckCqkMxECDQMRE1zOw1O/XfWICsmGBn+JQ8IyyvBbx
dD9SxuNx1foPNF7luICrnP1kpc6LpgcJTU+VMdJl69JAom4gPaZE1JFXjgmhOiSV
dhQXtQ7IKBjUDg70NogsLiXOTKQT/9Uqozo5IVOmsFerTTAC9YD/ru6UpbcjoqMO
kK03pOSePodLAvJYDwl7evhpDHtI38R97/iVGDfC3HRNzmhuEB4etXC5MX6DnDu1
e9YU6En1L85/3KbSHKl/2oZeuLY7sO4IMKJU73HgixUnnVAivWC35ovDlUmDgFVq
p0nc+gH9GsCVeqjpR+VqePkkJ5C8rjzD0jkTN2zfr2axfR1VX8XPHtt07rCeFYMH
nNoi6cd9YXXnTPpEw6dLqf5sBbcNtKW7BRXn/tAlTr2l5+uX0IQKxC2xmDprUsq+
jEY8mJ9jcBr+Es3VfQlNbqsLDEg8XU36JS2dVxEG5vCWVHjf7BhLhgXEvZiNSAhE
21C/MbTQugCmBH100gokGSTW0YRH64B+LR3XhxQmGhYnAeUSM82Zl2656lNeRz0I
S0tNsJMRj/bwzywyCCLkJffew+jSMNIXZnBn+v4azpyQZEfNie7pohHD6Ewi8UpC
myyfDtVGdZr5ebiLw7EP+BuevNbaIWNCbChWiMYVdx+RRwqcnUYb0uN8rQEQs4Im
UH94X9qoyCJ8Wsazjjyvn0ywmFR30qJ0EtZOtnSKZuvuF0KwuWSHg9EQsV5fqpAt
Gi6pm3eojp88v7CkubcubJPCS/gjuLfw00lDd73IdJlRzPWa4Pk+6Zf1KSAMl3vn
gjXG7HmDNMnpZFgKOM7R09DCiAntHtAPVnnBoUQxEeG/mo2MhWV0PGm4UPLBOd3n
60s9EIf292nsRerntqSqpMf5akqsZ2pcn1DF996pGYDV3aCJ7Qa8fm4VBKlopcQ2
yXGNdiRnjb/qqV6BITeUWH3miVZG5qJG/U9LUbUU+Heb5bUBUDf506Zx46sbOGrS
mGy7INjc3iL6BLdQ7pwk2RN9AcFZghx2vzrpVXAd5y5Blo8aLePKRYs4drk3dfYQ
0pL6XP8snSHxmxIh6Icw42NuO5y93Vv4KspCfcD2TKwSwx9wn6iltaS5h1Shq70o
iLpvQMos4+iLMsxk4AyzP3NUY5ej9fMazvkMxzc1C5KbKtCSlvcQBLvTeppEMDtT
6zO83V3BgoHVMzHMpyC+rXGiRqZvLu8ZJaOWGkj6kEO74RqL0L+oq66O4i+ziyZk
8LC/Sa6ZpDImmdyapU4qSTNETEjfo68269TE888RbiyicbTPDuogyZQWcD61psLq
KwDOjJPb/4N6yoIHodNw3kXzrJy2LiRJ3yu7aOD1Titup+75r4j+fDPUqTIIvPhQ
HTaKwccD2ED4Gk53lE5S44xWVjNXAyH2f211061WTZq40vYHZ0IPyEBuMBLD/w2g
jBJgd8VqefGp0hMyhsQgiFa9x/Gqg/I2BBB7r//X/X8hA68qBdwy4GJC0v5Xy74e
S4N/ug/ZvDxlcMAFGbPwkw6HbbasY7QvsCOajErE2/XVhBy7dOWrvILBdg29SI0m
uY5x+2gEPaOMrljibBV5uth35AnShFiWRBmIUIci5bxNQWa64hbVl9uCpBYGrB1F
aoTh9/vxwpYaodKLrKXbFOPnC9M/cNHz4BRYqsnoL37TSxIoraZjKXotljmnHO3J
SSkUb01hYByZTlGhATMC7JVEUpZxz/doXevN6QlxyikYA3IBYBKhLO+JgAiCkxxF
XkwfeRLx/u1XdH+1waem9PAHxgBuizbE3kywGB73+kB4yzOTBd/pe8hfZA4e+lga
kfKmNqU4rgxq6bbBTbPtoPw49Zhfg2yH/uOK/Z+sVh5oD2/vt/OugZzlljYeQxiU
kE/zJlLZuiYOssMYMSdkj7f6JK162mCzp+DoLfezv33ZV/0xmQnnjhbgBprblqnr
7ql+nWS91j8uaeI+bA6v5vcQ06W9oE5ydJKPlY3tJpGoVQ4kR9QrfVMPW8JQzYgK
+AvJ1INAoo3u5/M195dQqkUXidtc97HO09yKwqAZEqzUExotXWSM2/srQEgUCtvU
GxfwzzkOOY3tE23jAuc1o4WaAYNOsTdw/4P6XfkR17MKWIVVDBNY1b1dDW77vDK6
R3iX/LppIxMEhm57gz4yHV4ZaHC9A5SS5W3GsgAqLF4fb54rByQEBkX/9O//HA20
tAC8yi2+n0/0Pte7RUBk4GT4TTIr3htWUN6DgAQYzxcfBvY9QiNd7bZ3jsyCHsCF
4szWVYnU6U/EGB+bbDodrmnrH/SOtHGApxwl42EPapySebtrcz8E5xrKXBaffPYh
QHc4xLAlR9qaF/jCZYKKTFcNAELTuOQn62HCqKxOCfrDWPRWdtlS4RjPBN+EiP0k
7stqIT3ATZh23Mtc0Zm2O4hchjiFaNTUJBPpWH5jS7KdeEdGZBQL2uVvoNFu8IRf
P9BS7OqK9ggdJBqBuY8dAEwIH/8cBXJKVcZE8GGu5gSH28ui+goaMgwMv8HUXaUj
GTw3zQ6L8V1t7NCIMNYNq4EtbzEZ49BarRW47Fh8bEZQ+t8VTP19RQi8r5Cy33Jz
E48o5iXAYunX75dbqpjnRmFPt05earJMg7cAmaek4WXTb+Fx05WhfU54C/xTInqk
FYBhkTQbTQInNywPSZo+OlADS/c9stOhIKx0mOwpXH87ZuEJAxULvfafSmuzsAh7
cysnSgO+7FkzXHP33KWM/tCV8+HM8P3aTm1KiiRBcuH8Xb9VWw2sKyEPNpGSOu5/
iN4OQ4dSfp4jooOfrSXMoKZYTWMOheRNo5c8+haV1m7/MtiOGwupB4sdExwOsXFC
qUBwtYqyEssz+45anWxIwa8t/ElRoxXK87sm0U7sk7yVJ4r5blPB0qEFkjTPINP9
94ykVARV6xsx+OvzPywujnspj76qy9xJKqL+wV5tVk93cejx92XvmEiezbk9BiAv
1dS6paY7TyCT+Ri+StsOEOToLXtX5/dBc8wZajCJn8a27Wb7elbMrNX5bvM2wz0/
4hWqu5iWIr/gmnV1GxLgZUAImirPc7xn+exLBrgD0YeZQznHRUFVCBqIp8E99fPo
IUSdPk6PAYupHKFms14g58MMPQNxMxWMJLENdJ0XgdcdpfQsYnZL2NA1SOd+2ivY
mQksk8LTcNPzryrewOBs2D8v1uovxAInUerzTwQjaMXRn9F9AQ9xIJYc7VfAN+wl
5HJ5hJFYwEpyeL+wm/JxVX36mP9zSYwE5teQFMSOPcCyv7jkhGLCF1jTGz8UQ5sd
im5O0PwRs/dKEJi7qOHtq3w4YvE0DNs2YSTGTjbVgjanTZezs+AVCan/lqV+DFTi
LyMzr3Ll4x9UZY6AWwd9NWXfmKqpFWa0cOPvsifNiDGY7IzznUSkhvse0FMAruTj
ne+owY8n9V+j+BVKwifwRTymUdToJ6DHdTkNbkfbGU7HaQFOuvsK6CyJyrLD8Ewu
Qs0JP7ndTePWhWsfhmkj/bTgLbXz9ia66uKhnrl4ctaA5UPGdFRPbo9WkOlf8XnT
9BkkXQjYmiIQJ630sA6dG2E/Ohp8dD35dhVeSw5h4ghiI3mxQhnTgPCWIiAuWh6d
ww9jLKHWozbm+Rufo3dujkSeUgFMl6Xtx9QnKwBia+9zkNG65mT9u1PyOl1yaX4L
HKggSR8ufyYj04djhChd4KQPGKvvGUyd4SWtVgYHy91T4rISFKc9WawhBGD9dal0
ct/zu6IgDCCduZzo0C2O8xhwYTQgkHIeij0rC5whjpVJFWmFBJ8DTPYhtBXMy1cJ
jnsmhTjnsFp2swNr0+24tgqHkHRZfSAe7oAjNq8vTPu0JhfvpcJe15o3RWBuhSu4
AgYfc7Wmw5d9vc6ioeYfARwmDwy7BmeQd2uVLiba2M5DcdS9GP6GASKu1sEmMiSE
YmAcedHF7+BdpMV0zKVGJO6z9qjbPG77/qinDpxoUZimyxGmfw/90aMaFO/p8jwD
Z2HWxNwqml4SE9qJs/+MGBdRwLB2veLew8nD8u3Now0Eg9kFrL9frJDsZI/jCwOp
mokpQnCs0NRdCaYlIWxKNTOIO2gAq86ICfMogQ00F2gWGYPMKZet8TZbif2wCmwl
q9CAQXGivX8+V5tt624Z9C69WkvvUXJRJpiLlnyJLIxTaaZO1fmPfwQ7cYHECzlX
WTktbJRJ/jK2VGWG4yzrtlYWeOKnvxS5EA/qco7efKbkOC+sXhbe7PEe5BdCHPQS
gi3tQYdwqeRNMlW43C74BxI3rGiRg6+NjhQ2eOfBdT1zSeqmAWNvxQ8SGKI2N6Q4
CFlp+6M1lrIJXVE1kR+WJOykw6Brygq9j2eE6xH3ztS4YCGn4IYMgpYW2pNgLc7O
0nUgi8ZABvEFqX9eCM3CEZ2zft7OMhLKmx6jD0A5SRXcLmKp75HGszdOOERdShEd
kd3rRxGau69OX5YG6nyBAhcg9dtmhh8QekKAAHw9wbueWuj5SncZA8FIB/7zNdlH
8h1PZNAroP/NHSfe3E8QXf1oJhXBaNTmh8RrqvheMOMga41/wdI7M7WSnEtV4Dxb
L5GiED15QLothNBH3ozkvia9bWegTbTRksRfGCuiecryx6OtYMr2ZCH7zjYhbM9D
mMHajQGQX9Eb8Cf4fvXdZZBuCp0JHBWYeqJACvaDzFpU6ydOlDS2yIhk6/kVsUd1
XNeuq9fl829CyIUotBbLvd5HdH24oArcQ87fL8paV7tPjTLQ1R0kiz8sCPLVgm9M
YUf7XgCFbBjrX1anDf0SkbMeCqaikOYq172N46W8+ScZHkbxVLPm6AswwOQivbQ9
LNOXcvVv1GLe6Dzy2O8RLGBt5081GTTf2NmkSBiLKRRt5h1S5Q6FEf3caX61DoIw
z+W0e+Rro+/od+nuQ52X+HGGXXK3iW8BDPrRQMCa+6bIiG6srmUFERNDN6LfgIj5
Lrb8NyAkDZX2xukwWklehVSAnFLQEGWWM1BqI+7SXxmmJ086EuIFJoa72ekWj95s
L+shOA8iGpRPd9O+zroCqNTCAOszN30w25yX5aUqF6UPrpLM/oHn1Udm/e4GN+hm
rXa9YMs8sDhqPFub5r5lHBajO/p7H9+E8iDyACpNc1JATp6WLzLk+spWkGpNtzYH
j55pBjlwgeNO9gTFyMqCG+tTmq+nKcdF0Cv2dTqaYO+j4XMTNmLbcnkQfpB2FTw6
3Ohs412KrX3lBUY16Zr+T5vfs9hjFpKYwHPQ+euXG5Z8ng3CXxqx02XkMQm4UntV
WXsr27PH9zDHf4dWif14R42GGUJSu31gmGZIxDsRYgpgpwZkDR8MOR0RHWkbDlYA
wL9KoZxqXlmcP+kd3jMbY0HXjIoN/m4Hf0ay6J8KBP5eLJTxNhGw1Zk+2cUbB08k
gQvrhVFkW0rMu3s1wqVfjFBuKLiZVdaXnxp0Rmo7KFtHFICdYqFxZkdYWaBwn4AK
bLprrkNvPtEvGYkmWLFhYl1pfHPzUFPVdcS968NVjr2O+C6lwYGBMThjUbMvtdBs
Dasw6ChQdkyI+jRKcfJz/wl4DpmDyB9cqsLa4lZOm2CnJ1PT8lumdPlTvqUqfJAl
YYiu+DuRzpGemHYKFf5ftA5Oz5CFGkq+beQ8CHAR9GMBJHQSR4amWy81miAfTcE6
P6uxAEaKrW5RRBipOTwgDianrnbJyc6a09CcuHMAKqiqIH6XXnpW79Luph2NPQNf
Nj0k5KyPbn2I0tiRbFOV4VXo81S7J+E2qFC7wWQM8bgtW1Q36TEYAoe0+XYLBOH4
t9WNXCOaouYevdkXwfdQ8TQr3zCxQQslg8a5fX5cp2vyj8yybnk9T3K7Tcpv0EfK
7fzl2rj39fXPC6CUs6b+0WTOaWhCL/JMiQjzG2PxWT8VMe4AYe2OyklqaXqb2GdT
dZmmxvZiAYi2w6YAprrWTtpkYOmojM7e8wksQa9Snq7QjHz8VdVeSMuue7n2PXDO
KT5gHwdl8JaD7BpYY6Z9GUyAOxm6258X/xAgn3WDO1KoGoJ8pkqOjIxGX6nXwave
DT+U32UcKnJleJSZhk3CFoIqfMjx5/H1q5yUXz3AD9U8HgN7ObJxTsG+FK3qDQZA
Wg0QE8U+/Eyf/BfK2dvVsV2ARNS+Bf1qrpxBYdgQigvQsk4/FA4lPMMyj3zQa8mF
9MAPhy+5n+sXWtYBBp31Hs7eSvF76h6OxEIOC1QUGE1faCnut4A/ZnVTOEmBN9Q2
frD8ggLctcZrOCfhIIBTLLf4/QLVNo1VXO2GHafRwfvSTliYQLxZWyLdnQBrav16
1Ali0wV6sjW8wQABEpv+E8F/MXNHQ/DQxsWbU1QnpWK0cGo/IgVnHPzPwadG1Gcu
Azx2w6yqgu4AiyHnoEdKdvwdUaqWjhqsAUZYg184yDWALPzKFX3AxS6xrVsPUs48
Kw3yMTpJ8AEu+rJCERxoH6x4E8MUHuxZ5DbeB9Mg3aOBNVlj08ZJJbUySHdbneXw
e/hNMbp7CrwIQ4Oc3FtB2yA5SBssp3VHojxrgEQLxMXDWiHUl0y5yH7fNBGOlG28
EtTRIEVze9b+zsSWvZONOKmXeHauqX2Y/iJCHwY5DXu8MjRjRe9/n+leo0E3r4tQ
RXCEh7aoMw8rU7ClCfJ7ZNHcqbTPgQmQTiw5V1XI5Lg+vdmMZG4kNy9kF6nqdvBB
14/pGSId33d7iEArf69RxmcVEvY1IkkQdt65tr3MolW5N4mhAcZiq1+2Yw1HS9py
B+w2zRRYBeXZz/XWV6sRN8mjNyxEx5ourIBiw/Atbd8pUpi8N7vjwaNqeZeH/n/e
50+cw2QU4jj/4d+rr4bVP8ebC6NYB4UBflOKWJE3xYmFIqf88YrXJIELb/x/hvu8
HvEmJbhtQnm7M82zbhekMAy8PZeh5Zgu4ZdVVvXnPpT6zCdaUVopLGxgRiRy3w2m
wjLhI1nWFEOcF9CVToBmgnQGYr+6YevtQHDJQ5vgtaP/G53mnz7+q3HurN2VgZud
akClJZoFb3R8OO31nX/oOLP4U1aYtK/JDnepoIK4REtjyUwUuZr652GxGuhK7kqY
Qv99zRCqQ9/Em0bUYkBJpHeIcKJrhqnzGVpsEyCilgyoT/be1oDRuhAgKCZcA2hB
VdZtIiHH9T/Uho+kEXYUPB2SDy2C6SYkFcvcXBfHQuaAVCLiPM0qx06ZDyFc4pEe
KT2F80BkVKU1vgi1hnLnazSRf+WpZXZ5qkyiQW9PazRGTdRBYVjOjUuC1IP5l4Cb
/tyKih7h+1JnCYK0NHaDumTYQrYN4rn+5itufr3C6b649uzaKdXe48vVhRXX1VF9
NBWLfKCVCejK8JDrVyCPEk5AbRv7IBsa5ksVieddToqmkqcIJfM9mwMGwMMSQHU+
8ca5stJkNSU14UjIUFvRMqcxvwxIghdHNjdla1MExGuXh1EOTYxW8gilFbn8um8F
2mZX2pVskebG7Dc37C9upCRprFVIC+/AdekfhEMzQe8U9UH6/vnVSyel9SM75ocd
rmUBUCj3MwQWYZ+xDYOsG+bamLhIJYgl99B+0ivXkovyiBHMjCskpZkFCUh1gwf3
CYv4bIzjNPZcsWUfkyFyrsiONkYOuZ4wUFiABzZfoiMVyakmNDeI2noMCDrBHER/
P9wDJFBnfPPUSyTgXpUSR8Q573NxOiTCtLTyeBqzij3yR0Nt/2mvb6u2fUqi1IB3
rVBww9VRiqjvooLoPWbvqokT35TxadJ+EV5UCVbHQ0PaQBfYlLLlap1AB+GvoM5X
51wn7ZvUT++l65kZzuqvLdPjeALDFEieOJFIhIH8/37k3Ah27gzNBqh7cHJgXNOL
uA1q6NXXQd7IPSnDfU5INeQ69b3xRoqZ7PAk2WuyoQiKLl17Fvnc0M+wmzg9DztW
8v+fg/kU/sGGi6Icdpk2SpxRCdKaCW93esXKM1HGwxSReTk0Y/kXcP5aY+NFWpQc
Qru0cPhokI1brGH3azFr1Pr3zjXoyZV3F1bxTMpfpLSS3eob3b3FoP7kl24Rmber
tNYTz5M50JBEKOr0Xn29RMq6ceniYlckflK1nm8XCnaBwZYNSy190a/6XmZCnKZA
oYFpMrc2nVQWhMGp5cMUlcEcNE9NKlpwbHqaD+dmUp4sP4O9VHwQG5/sugdARLZ7
RdN7BnbWqiMGK8E20HSguS8lhMrja0dy5MekB2Om2oN0J1h8cVBsOQSD1TxoPHIk
rz70jdP7PS32oShksMsJxhzQ71wfraF9QA6oiHXQOKXHjgmnVSnW4wkLWXew7c09
eEwIp8FysMGqFtWJNgM4wiGsruN30XinD4aVHXklXngA9DcPJodKHNJDySsCMsFx
zWh/P5zJxnwtoP1fJbdVdjP2vdqkxihRtyfYmQXtzjELc3fQDYXC/eAyrpVlHvcp
OG3cnOTmVQRi13qagNovSF7PxcuwdDXg5yj0IrAf3gwvfb0g6vb1chRChoM6PxUG
WBZhwTojHX/8JNvPQgRMbpsYGswmdscbx52Q+Pg3yfsfXJFwJ1LQaqnNniYy34rs
iXGC+O678Bky61ilC9pagX4zNpmNXy4nP8ncI09y/Ao+xrbG12z4zKMPicO4gqwP
UE0mBW6Knegag/wTSQeBc4Hf3P7IEt5eAU+2yhjx/I8BmQq0StKQNndkztVcNpaW
vX7tx7b6A2vYQG0dhrxmNYgzt3iE5SfJ/+6v9YtkRY+qjOzL7dzdMaH6T7Xv35R9
E9aLs5sHqgvi9AxsNKTiQNLxXr+bKgK0KCW8PJo/YeFOPsbjUlcpR2w3cP4dwGDD
X3qU1cAXusXFPmNVWvMa1Bn7CPL8jQDHMThcPRtZuOaAtt528EZQJoMW4NMz5snn
+fMpETS3BrdrDd/Gk7e5vG/4ECi2LmSUjQlfBRBVb+JYhLW5CS5TUDF/0IvMdikL
s9VG0DpXtc6wJb0J7w+NVCOkGKHx5k5jMRmag+xYzMT0IaatkYqlLd4v4nQC2P3l
fZLPvZE7nOv52C9zXBJtzfjMjktYiZ0SGtxGqGpApVUFqJe6xErJa4BjLnrCTZv2
HLAR9VT2+ElkzcwqsBJeEzSK3ORD7XYcEPIE7lxtrgyij8smjeDGgf76ymUiuoxe
pQx68sbyNnEH5QzEk7S8DyC21MymZgYxkaKpjlOiinlo2J26Y70DsuPRoDvD8lj+
bQsmv+bwqeNHyll2kHzWLxFwXfWfcXFmQu1zomV14+pvljWdwp4C3A7EaN+XnBzp
D6P56CONddDca62TCyA+bKB7k4vgdgy0zo47MqPbpQWhZlrF2VMSKVeZCvVNckY9
e/tP9j4opvG93vVf4EUXTUDPdrQMfq7QQ5k2C6I+6dQpZs2S4YS6hCWJU/JD1XJX
89mseJb3bbmF4dQlNhOG9LI0roL6MADai6W9YaKh8xtsoeKuCXIEFutN6Js5xLsT
MIBspYINRJo1oRiJE8e8BLYF6G9/sn4AAai7NFcLahJEvfqP7hU8VvIWuaH9V7hb
HYC+TPo+qKmbzuq6nkaUsN3a4/f02cyaPbj7dzBIB1yLW3xLDGRYgvWLhSABr8Ji
jo6x+FJimiOjGcyUt8m2m7i+r5Sg41UDwszGxe+hnPAIJGLsxIWFwkCs4PuElhqc
HSSrdGW94ZD5eb1wmwljgNgdP+Q9A6+kAiDSiBAw0jhYoEERkXclHGNLdPPLNPJB
ilt2LQ4L6tDpFdIFI8IRk+OPKyR5RefzFfeByWFRu/9NdQ3GibKCMqaLZ1Q+GiEK
mJQM7v8dJBEnObY8OXSxtTt1MnwrVPTuE5u1pSfcT9Z0pJ99WE57Obt3eqMeJv8X
shtlAyRV+ERNxSCeV0szuIn6oBlo4wcVuBBDhxv1L07Jr1am21iXZ8nr5Xx8ozsP
XljdBvHoM5KXLRK8jVOC0Zy4wNxsDT9YHszcFrEhnitntwXxMaXcUKLYx86BL3Dz
kcoFdD6z1ftuwXCpTjpsLVsJV8RVIoaL9wW6IcDNI3wzUIPgitA2kyU8EC7w+DGM
WrzcpQbitdV6SxTAHmY9ec3/KIxDaLTitIHsmUcrBbskH1qe++DO4WZI8F6Glaky
IZGoTAmrgmnZZNvsOiJO+FuYMcFr2dgDAKmkx5eY6o8Uzi80UCv1eAWZwiX+o8tX
C3AVbPsBUk3axv1fz1f9ebFEKAmAtqT10EWpxkXYkdbS8+juMJKPmz/5vSpgrjPn
nK2gMuRE7c6ZMiHZu60Bk0q0jaqCfZIHOlEsB/qACKnlyRsCuRINdxrKWI/+VdJE
USH+BRh6wf1xKV8xQoYHGzbWLqilhAoUXNBBuqZuefvmUnhSVyRgiUDckRQauD0O
r9B/sGjEDSYAGOd0fG9A47hoGqtPRSjyIpYAsph/6YaKXukHCOJ4upVzaRrBOZFl
vrzkvj62aLl6/X5+NYm9eJpFJgVw4oFdr4Pg69G6skLfUXaqFbXe9p3irrqbnFRV
JJnchFoM+fU2tisGbx0YLFBHK6mzmkI/k/m2hfINhf2LqlBBasnA+T0U9M7neAVn
5gadDT9vldBfs9SWRkxumtFm0Ry+hONmQoYFTOyxa8BmpNEcarG3f2hMw+rJWYPs
TarRftHzg1DLe2pglM+uCTfOZFQe6CC6WuVdtd83XLegD2Sug5U3H8jnSIC2swwI
Kj2bgq7VhmHUekJuSJDqDVV19OGqMlADCe1oE4YSUQK9O3P3tQGa9R2Lkhv1Mwbu
wkut5IBAk0nNXAFI1YigsFkjkoPWYx6M/Y+GHb9VdjxmimOg1S8Z47me2KeQTHhd
a/IJlwziuD7/+Jh8B9PmcXORq07rJ62bzTlsWBspQJQNINn6b96/BmGAvOqsUSFp
zJIesxuZLKCBqyU6J9Ud9dBy/uo13UDnF0Eb/upfKNjyO0M0uP95isqQUE2J5nTH
cpdQvPGW2qJUW0qR/ha2ZQ0wvgY6X8PodCs2eUhEptMLvYYsYhCmTiHpyR7kSa40
AjslZiTsBPP682fFzYEcOC+M0QNqqX0hWZJecHifaFed+8KSge776+hvnpyUjE4k
9asnF/gxS1sHT4V8Dd36ujT7EhcJiTqGx+au6HLYLf3N5/W1pNUlr33ELTGIXXjP
E0+8JN1NgFHlmads2dvxBPhIEzFXZp6OiO19p8tp+HFIGyt0Jx/9FyJEdndK7+1K
7s8KfTuBd218tozQXonz+z8dHoEdasFDL4gkBsw47reI/ogryIraJrr72bUx3+mg
PB88wxEBj6Sbi/qIVR2pyQeJ9Fb4vwVfT0EDFVzeRwn/WEeRka38UWJlZKvfmlYz
CG1fF8dZtL9/nUefNSlKuW5uvwNo1TmQw2szXW+GCfyzV5DsDVL7YAPNiQZDQQNl
SHPh3dCvgfMrpN3FzuOgL6vAE7o6HwNBkeywSkHydzj67/S51QYR3ZN0m0h9rJ7f
+lYfArj3YaF3wvvqqtFSKqiblHWLKNoOq9Y93sRdcuBGpWdprJOtGQGZeHSVbkvt
L1JxHa4Mlu6A01/uCyTBWwz/f5YssxqclOQiB8m6OoZZW42zouSK5IY0ln5Nh551
vaKvJt7MEamVYeafaAl8G4rbTPOF6cnpj8l50WVry2apmBopWyQpOECFbwP2Ts25
eiXKiRLO822o4WfQ6nhPSscmTzXG4SLxeHqMdYQaXTrqLPDITkv8WUpgQ224GxbW
ro1Qq3n/ocX9Qtv9yPEexZYsKh+5mfiq9m7X2G5sLZup9NOivesdEfsWWRV7gyk/
YxiSPCRebjw/afMx3hJck+DH6uGk6d56N2EgURfjL1GKnKW5d9kH09YaG5u8AwDU
5Sali1loKrZRy2GNbeXF2/CH6nmNv7JHQFGPT0tbot/sWE83Tzd82TFtIre/XDGp
x+qBUw3wCC3qUGcdBwa0sQlqBoevHhnsUN3LgwqM71vQtw3eLJse4IzZG25MDBfE
pFDf5ZkrMONnohhD73A0KIBFyjPnJ8othhT1dfaAJ849gldArSXmBnMemvt+5KXP
K9kzd3RW+et+FGDUCi5ugS0y8Ps0kXBLuY6V4RXbdyg/NSDytYVKDbnmG+RJAg9s
fzysbckkuCkZ/TrYsedtoT9OrdE43GyZkyYJioeUOQ9rV/fVKPj17BtT7f1q8ZLK
fy24MefkFEvjWJVynfdlmiV0wlL05WwnsdTcU8cfEsoqawDq9hEce/UIjHIlLW88
wIyzMkyj1MvRIjWxNx1KWiwJIoB9hgxT25fp/G2nD5jF3+Qi+cXYx8QEQKhGVDve
KB4BS+NbQQp5GYPzTIag7vLIXca+zAN9xskTwnn/0uvyQqLyJ8pg+p9jNwvkCadh
RaEEH/+HeVNyrSP0iLPs3qmhwVGhKJda1cuNLkd8v1SUhT4Kg2eqODXYmoOZ1TVc
2qPrzXQlI8THpk2WltwpL+wDhlQo07BXzFl9g9HUPVhIlwsfHubXB7ckWcIP49gR
/AesUiC9qnbcB6Cu312Eq4kkbamf55MJqm7P1FEHjArrbV/C7a1Km/MoFFVLbf5M
ESCw3+c57S3KqCXdMWuG5w7fzoE2gF5c/s5GJve6qnzv4Q/9QhmNMOHGxDfg5D5t
gQxyQ2gkGilh5Qf11bXfa/pPHASuo5FkhOgMQz8O36yn6Q1I3+ED6ikv4KNBL/U2
XBCLT0HRs1vT3PuYP8BDkFYGG0R7/NjlcOEFoGMpkpWwgHEWyRXs1btZUzUoEABb
HlPBS6qPPiS34VxO4Y4xkH2o5YCYJfPtBoM4f3ympHIHbLaS1ZbeYJd9UkiEa0bz
cQmZaZ4y7IJ6SCfeyvCIFiaarHcUUzc+YFq1uE1/DHHYE8n7tStKLLpE/HFAYYD3
Akdcu04854QV6J85SU+VrwxitPcNfphiZX/YutcAMsPRxpWnwKBfMV5Xh2soE7sp
IG2qcc25x+AHV9TuUHQJ8fG/rA8vAoJbpajVhlutkiYDUMPmnyPtOPAc1XwDLbUo
8RlBUtCo1aJ4U6qsOE66VFBNz2YEBOoniLY8PEs7HA7XR7atKCPkhdXvP433akCN
gl9fWiwe9DNV5B9YqSLRluCNDEkqa5+0AN4Egx+mfGl3WrAt4cTYI7Ldzk7XWByZ
ISc7b7OsRX1+ZzxSHV5dh1AxeoMUM9qBxs/EK4jrYh7Fmj4zgor6lV40hR7foSNo
D6qTVymUlJWgbk3h+Xlemr1qzz7X4sB4l8IXj+uTNe8XQdFIncFHe0Eg4wWTI7lf
u8rLeGzXrYZNpVJwELssYcXyAukRiUvSMbKuaYsWWQcVSKCB7nq0JnbOUnKq8FCx
hjwGa5l9PjWJhHwINxF/6u4wieBiReNp3ZLyrUDyXzeSUCGiwlTiEDvEXPRABUrb
8dHDqMGABlfJlkWYEc6apwKx10t4BlSTKaNwC32Fj6WzB8l7a0JpiOK7I2iPYqvL
jjaDXV2NMuoFBX2BSIh4sX9me5ZgD0lq1zqDB2FBFw1quG6pPFOn/TpWrrC3AkGn
wCmZwk0GCPsBwxSuQL4lBr5UKRfBtua/fDArTJxOYy5dZHvX4Sd00nTbv84HJHjl
IC/v+CA9UlfK1gB7k5f2E3XCm/ddUOz9evKKgGU6LcCUt2tKW4TaaRSPRoylPmAj
FvLNU0/rbUmbJmPUhaHQ3uR/QcPO8nsMJ0j/GaNNIh+Updry1AyfbvbZv/2vaL2b
+aJ6wn/W1Nhm8lBuabujFhfEWM2Fz8/Uwrivr/jO9aZ38pKIsaDPcUq1I1QkTq+b
8HPApmFia92wLJiIlz6OYQ7APUnxiU0q3IwtoggD9ezEXAnYVTnoHJAoLm3oDXcV
NMEMgykZ2Mb2Hx7oiCSIFnrDu2ORUE+Ubl/RgvyiYYhsjPKWBPbXz1Lwitw7GGfd
arIxJqcNW+4xpM6bEtsxY09aA33hTy1JA6LR/7tXOrQBce3mEFDARG4ahZnP0OAS
E0MlMVR4FpB2wFye/V8znuNvDNHzn36HKSTRNkb7F7oMaM//a1Z+wglAaRIgDySN
YKZrCT3awjJAA2L3hLxsr/LeabRVZX6JC046WvsYfBhVC0K+gBbdrBpcE6Gp8/4H
mwUR89C6a0gq/KeKnAvhfV8FNZC65QX/6UtsmTpd2r8c4+0WzkGkaztrlXoEfdgZ
hcCXvpnQo4nqa9HAwDVRoAtERxKYLJojlk9lHqPyZJ+6S6cTfz0F0Z5LYC1/nY5U
hZRKOTNZQOGFKxqnHW3NXFK/PrjfZHYRkuo2xXzoAbJa8aRIT6a4T7wjetCwI8lr
jUtPtVOMsR3Z8Okz6BDlctYU/Niox0TwZ+cxoAslFgxpqixMflSthiM4nJwifHDH
FSQv+V3I/eUZv3gqRQ2B/ZQQL1o3rzkWqIGjvEQW+htgg362Zqf7+HiE3gkn6//A
Zlym3XUs+7iiPH+PqOh0/dHBoJEkXq7Rv9w+LmT67wWaOq6m66Q3mc9cFZl4W+G5
4hiOSKkeu3mY9rspAb7EWWkat/54v9xC8umtVNG4vzpt/14imeGzA45Ws0LW4qV9
R1pTZmmknOMZs+X71OnMyG3LU+hDG1xF4mubKi3aj4okL4olN7emmzaETa+xGjcL
2kglCYsm+MONd/NRZgU/up1qzMCdoFbl609XBUiknwiOpieB3iPms6zzfzs1poSQ
aQf1ZqofuK6ZtxEujqPyvtDwHbFfHE02oLnAWSYxFNkE9x6vrTdUndlO+k5b2IOF
Xqqt/U/1UCewHXyTNtkFXVh9i3sCfSBSq3QRLZRl5jtxtseKXrW27XinNkb8EYMw
HSPQRTynrud9Jf3uOgz5CNLu1hpA2xJglllxbDxg1K1jbHhZLhLAzMAX/2tmE0d4
gJDpRjcKhyDXh3IaQIui6/a4hUMRD4DxX1ie+BEhkARYiZSjjzcswkJgmjDVD5Kx
eu/8XHTI+KlcFzCHF6Ezy5ajCVDt2DYYESoc3C0X0v6z6Q3/3kjQ8XaZ368OORcz
yvGDHWQcINhPIvCYGxONk1hK001cHIjivfN7YjOfPgJtavRyJXbVsBu9qUczGHHn
1DVp0iw87tX7t4t7jxY2JPk6WdO1wEHVaguC+FNewkRwaFibbctyGEUSmu4xD9Qi
g2qLXcnVPyRYJxuWcaqTddLhsas0eUPWftpZ0DZktp0Im7kLat3r8jKNV2K1J4Ah
76cLKYV4ImFFn6pwc+ZZLoTQilSWnNHLlckoCmUxbO3+B1mU7ABs1nNRmne1dq67
V0ekgwLPEZi7B1iy8SUxxNwwZjVYblSfUoMQp9Mszb/g3z+/LH7daqspp23l6UDu
P+6HrwpUvHqpa7VgmM0E+p1Wcuuz81hQ323+5kYzHdju/IaEhF3/3LD9rpYq0A3k
6dAbs1ZBhoUrzsSYDZC1+3ATeoqWxiVGqvTPejQKEQyrZZFtOoThwsCMAK7lu4K4
QVTYK9D/HxyY1Cwg7+QnqgLRCqx6UaxF8lbSLnvd8V+PD/QNtMPOolaxbS1Gc52u
RoMBS2yVkd24hszAsdj28PoPI+/enBrLv8o/n8Qwrs3nQ7LIC44k+prBEpPhGeZj
ZNG6QjgfD+hq8xgVTpmgHmDMGzIjZuNhah1Nr4sp36GRVYFORC/Uko5CHiplSv8X
Ot0hOTc2psCtA+LkW3bFEEIgjKMph1P8FrariC1t87wroIEl/xP+2HyxzA3r+d6I
JLiWt3n5kijHrvH4h2L8JQANb/WMgx3np9XqVc3tyQH2zjkLfXGVIpZQBQr9FSJG
PHvP2kXNlpMzFRdlrZqGpoHaTzI/R3aZocTIyzGA8CjCsBVtkyWEEXXYXzguWWcs
OL9V/etuCVaFkNI/254+EXFDsbjzRt3NgfZUjYx0Yw9Idf2eFo+SCtJdWxPV/jeF
BLPO9NVHoHuZ66XCIOMWKZ1Ch8RegpeBf847y7CwF3jRsvBdQHA9FkfNmRQIdgOJ
FB9LicWb+n79b/FRaavih6pcv6b1GkTv8QUDiSut3/NktObsR4eB7MAXaT9l4W3Z
gFnNgPpLVOJMvOpYfhhGP1PCKS8rebxoTtPBn+7DH6yo2rlxl+Kkh7WLm0c15991
QL8Op3IrotHh7iYfk/Q8DT9Pai6iBtt0PFsxj2dnwF52Fyaj5/VoAibCEr0ARvtE
mxhT/K8PnYP3jC86JwQZQOAJz0eVvRumPqYCtN1hgINlC5il+IkBjULM8fcYon8O
1WTk+puiL4hCSBDUV+tk33D2xR0A6VR29WHyTUyBFFiD0jvmLSlH6sGX2eo7o9Oa
myVb/gyNbY5xjsZnxKMACVBEo57K/m40SamzfL9Rp3aJsA54kI5u7WBXx4cj2xrG
oL2dnAgIChHXgAvvNK18ujOBlo1Qbog68TA9IWUhxDO+rx9uld2qbR+MVDYVTj1F
GHP5HfiaVJxa7n2lsPcM3ibt+h1WgRKfgmkt7zyAKsRnHzGuRwp6jUg23D8d+Fe6
E6TnuRggaCZjM101bWc8k+6SeYN/k6SsOJRKwgVnjGSU5cC8yiaTtNRlu7KHjuQN
10opakehD9Fj6Ktn4UNp5lkQcno+lU9hgviDLBLrw2fqt93L5EzI2NovY/m2XxWF
z8zw/w2W+Y91/+FAslsaUwfIEp4NvGICfgVQiQQmDJF2TvZUHsopQXdh+0uooN7f
vadsnZJXKGgcXQER+/Kd5F6+I05E8WqNzuoy0/f1PLw7tyNhPplPFavWqtbdNEdm
3UfFGbKFIm/ovG30h3sAkN5sN4CDv2WZ2lI+l4paQe+paBeikeCJh0qXwZRx3EH3
QNcvDdyq25UhsTxgw7BIxtc/33KPls2HiaI5HYncqivGCHAAmeeB34QajcD+jl0K
U18s4Uvg1acDzuToN+pYe4K1ma2uscwW9TOU/KKYJvFfQGrLU5CqHaUTHaH2nlhs
MYC4vTovJCFvYcoIJXJo27r4n7GUyh6PHZci3YG46iCJgOd1NvbR097ZqcAuRtKS
ucnUQFIW5oRUkVhclRpGr579/jj+ttPv+URRccfWQtq6QNgNI0l9fC8QOtWIRfLA
FBwdqaamAQp+CUHYGf/2hDYpYjJwPvOneGUIPwJ+TEEH4hbRLjV+Naopj9TNPMnv
ZJAkjRsOAYSGqNiy9FU0JanViyygjF+jXtHViu2n4RHjmRRGYZeejVy6ZkYzDHy8
qKVU9r5I9YMnxgGkd80+yfxb+1tEk0voUpxKeGADeGVhJFqB7VkbnvLVmLgvWhaM
37mCCS0FoJSOpFEGuQCSleDlLmhviAWryQ/EEzEsWwsaJdRTomD0bQj5ECXZFNMq
OuNu7D0S5oWzpBRDk/Hbx4eYvqUC+VAZ1vQ3YUI6VD7d4GVKaGbNjUmQAcbF5bmp
vToewu470ZY9COLWG+PiWqMh53s09lL6Uzv3XEGKh39tBN+MUcOKySa11ClzTJ8n
YwmyAlTad16HOpJkTiD5G3S07WpZD4o57f+T2hJ00QMPobv5e7YKe52tsVibQo5e
cWB/E72K2mqXgbkanwWpQO5oY3Hy9m1gn7RqSRD3owiW76RKqxLWHfB8v6WcZspg
gl0ZsTKot12qzso+gCoRiSFaVfJXO1J51S1RsRKuJ/oI0v0F1UFDGPNSGFvsZ3iq
PK2nKJ32I368I+TCdSPpyzt0TtBJ+/zE/BxWYXuGsHvCTlMe46l6ASQOdaovCOZq
kyBm1ZA+5h5S7h8R8WmtYA==
`pragma protect end_protected
