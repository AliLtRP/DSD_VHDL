// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:01 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WkUXQmEhl6rQe54diDV2rFGyuQz3G8sYrhU83NnE1KHYDt4eIA7xXxkzRtwC2UpE
/t/gksySu4kzo6Bx4hWG2Gi3aJYyGtTkFcZuTfkLnBLO01S4znZwO9vCScNP3BOQ
Ek07BduBZ0dT92+o8s7BG93gyIlKpfNuKd+qTrWeJbY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17840)
iGWvqoloEFJptfRNQ77++0WXWCuC+3VJsfzqKv5//yfFC1b35g0MdFSRVSEtpdYP
DWCgsD62byKDNO3+8godhlEPcgcwTR8CJ+9PORHzTsIzhVvmydTOC3JsP9xyyGzG
c4zfCmjifTriJpZMEpIDr/XSiTahhzivS/VhmvKBlF9ppj4Y1s1xDu4MbXGTYIXA
9th2ghoVMQvU29sxJr6UyRUpD8lCT19cX4soMVT5EciP0KEOSJTO3UP9b82t4M2w
ohp0kNuDF3ray1UxeTGz5Kb8TWNWJ7RLLmbj2aMpXl/ABT9NlfjJbQAYSTxni4qJ
GzZ+Y+BF7YkO/v8DyHM86fxCOsyRdANlIFaAuvxPwTDqr4HYn3f7M8uzaJnvZjFu
8eLc8CUfY2rfJSRQRJNVy3n4iLQf9yQGxKOfoJgxWrdQayt1AZVjnpedY+7keptm
iIY6FKkM5h51RgLeBA28NTIpVFHXbzulZqplqKiMTTnGWPWBBco/NL0ZJuYyzHBO
ElxtFNea6IqXeX1WRneYe7d04WvKROTW8/tzs+33YlkVEGkNFnEfMYrjCgFJKsyx
gpovyvwCH7kWNb6TcalndHJgyXiJOS+aY1JKnVAUQ8ODgL8H8jgM7vcpH4Fb7Nz0
OJvO6ky6tVEQRgWpVCVe9pwHflUXYkyrvZucfew3M3wW1zrMBdVbr39RFmmd3PNR
S+3eEl5uoVwEWWExxkF9eSqrzXbwVCVAEeqlfz4ylprlRpPz0dzyion41Y5AylLN
Eeq4T56qS52TpNl0hwMvngk8dB/iMj0YGvkwjMyerj9D/x6lDZB+nkShODJITECP
NIRbXfGV4buCdugAMO7zlqRYsKRqavfX7csy6Mf/HT8xZH1c27YSr+iyIIR4hEO2
iOD7Xfc6t7wS9R9cxnFxklurubYjDczPMb363Mkr/fG/2KgoXCpdK9pIxd6B5DM5
9v8tReU7tLVJIFrLqGEivq8JKLYcmFTthJUq0Z8gLsLpiLnnc679mbvRfLugpARP
EOjKKn27t4tTcVbiJm5eIVjUcuqp7vg4njD2ZmlJJ+N+AwdLBwcnEotWjfhdE0fw
i+yYrNfVICSToIPe1G9qapfaXHafEEMBl/LNHXslbhqcNC34uWbWfQnZtYau404d
JDJNmscXI7SGt7ZtQ40lcb254KOYjtZHe+lIpRDZLxFXVEM/wSQJRFis+uMIYpYC
t9Fdab6t0bRZd6Pwz1lyYHf5Sp4xeEBL9VEuZ0e6ZienqzzzGQqlR4De6jag3Xpf
RZirJcOrfSyIwqWfK/8ttmrq6v/6cLE0w3C7iJDUZdepdsQPcj3wvMAlKeuZd98q
dle6silbKPm1OL0aCEq1U+9zS4oOQw0Zfvu1pjFfDfh+HQMkhVkwBmvjCYj6n5OI
UDDioBYf2MINLrbFfeAdhIarCeIDug97EIquxuiKrF2y6rXFODSYcCQmPtIE1cDO
Ws8BKXCADVuavKhhKK5VdvQ8Ag6vPXmd7L2X8FMHNpMMKtjtTCja+rQorTjgLF8V
gQH1VkvNNbgn1R+lHnIQXeV36tuniK0LpsJIiJk1IdkITNQw4et2cqOQ2k11MVLi
M6rLWaBSp1dbV6Y3bq4rxvdd6iORAZ+QhWObyio2IdgO3QSch94QsjAHDfwrX1mi
tqJu3jLm7F6SwqSJfjupOcoz5lPupsYrOpZnULKOEuBjqwWJ9VF37k1pqnply85o
pVx6ZfjNbope5MBfwcUIXEuY2g+Wyhij9uyHYX90y23iOVHz2tugroP/A2uNvr9L
snRX9tY3phD8gijYaS2qtubLx7wf9fhnZQq3c9ey3qeWoPA5JSsdanE0nzHQpYlH
cevYJ08jiezASl5gBXqSbzSQ0mLzyoR9fXMmMlB65DfTTSptSOblIvoM+y9q0nIc
fDViQk6+J5QrC90P3+vN70+8p+BsV1PGHbLTIeJ4a5AGogbbp92gKJPKEKQm9oim
CT5bLHBBHnTSqSDRmnKiucYJF4Tc+UerRqaiktKu6jEyJZw4Owe4jccFNObZ6kpn
f3tDbIMn2jocznNDyxmMraYPE+8D9QiamF/D5U9wUH7cM2BJc7YVLZoaknXqeNgO
wXMyTOeiercnCxSF/e+HWkLhpuoMHQn+jarLDn2nV3ZkPB7BCCtavQAxpHku+Cvt
J9bUC3GxDX/mFVs0mBqGMHZtNc2oB0ATO/e5Vb1YRKK1Vk+W9pIXVxRLS4VHCL+t
sXT4gaszT0VGxfjeHZJFSFdxZSDfv3HTIAlnNTHzp0c0SlVpE+bEBKp7r76xP61c
jv9lF/fR5Yd2wg0LHyal1GcJLChYPUzJIudnchSrYlUu7mwFI/UN7TV0eHbSprdn
AY86W4QdIcOeurhaBRZb3GurT9at5rvISNg3AISpLG7/N/4s6tdY/W0miSSuJ4lq
rEHWaA+KHgk/TA79fXtyMmPd3DnDLCCkrrjcWkihFGUJxCLKaFUyGV7gg8pFdpkA
npJYcC7S8HX1jSnlAvvB2j1YPJmosJXT0xmFNAc1Cckw5/yZxp7HLu79Frl1eGcj
SAzba86l0c77LEQzAnuCaflgQZbkJqj0NYv0/Em9brN9+uPrD3xp41NOhhURIeyn
mqcAy4N9WdLor7rNk4XNzn4hg4KQk/3xiIJ7kDQx5ZYiJsuJjYmWCCVgn1TSN3Vw
cCzFW1qG9eOzVWlEYY51cVroSyXy4/31jSyyaWOpJ79z+1X7XjdV7EcT/MATMUZZ
kV0FfInHD0ZgaWqWSQV7XLZ+rXLWUdzaiTDo4n1kM8p16KXkXVrIoeDFv/MZdvd3
Y8RFGTdYtWuUNUuDa2HEtqf4rqihbaerFTpHWMjnkGSWQ3ePwWG3ZcLVKpMMj5yZ
hPvPzRZZqN3Zkm7K7wpvYy7g6VZ3kfEt12lW/pbSCeY+ZxwiYp/VnJRjezAKKEYi
LgZVwh5+op1uZkZoBwhy5SZvbm9UKP+7tzgiyNzAkDwcsiDfsOxzwyDWDbIDPcpt
fuqppo90t3AmY0pXRl3bJFJ9M2mf66PV9AFWupuyYsneXTw6PaJ2Rd5R/Lw9Y/5S
yE6sePnHExE/JJOg16kZK7tpnIkRlwFmB1sYfoCGc4wnreIT3z5nUq1JsT+4xUpx
DCi7xHoxqHdDJM7HMd0HOrpgmKO6e0ONF/za+npTnLzc/diSU8xfKg4nNpEu0dna
SlUN1up0x7bv16pPA7fZbj2HCkt55Mpemh/xlpVJ/WkAN8GCNu87a09qOjSMQZ+s
KBk6JrB+TJQnAzMB2JBuwp7Qo6MOkKMlc8TfRj93fQlbooFr6ParfmWwpKBfVGJG
ATFT9rMsYwHKWkHYQFT869QrTVApQak8N44168Jhi6YrKFdtpClC3i74gBBfdMSB
pcejIiCE7G3KKMPFOHeifFhdO1zleXKu73KBQtDIv8/p18WtClUkkCNA4OjETiIq
Bn9POwBophjf16wfERzt0SAneL0Toqx8gQ0cJL0j945gTQSo1VyMQ7xxvd/MpB7S
DF8OvD3HUKnFS8lxwevzuDKUNK0cp15KPQ/gzBBk/HWuW8dM9zCS+kbVe6w4aTmW
hNNyDIuwE+RBjLq33XkZpSiMI/LmXpJIgZeOhOfYjGiG+pu0Cmd18EXTv8cytvH9
H4WK3qRh75z/KoA2wBXrtOhXGoISlosOqKUmdoE+Lb+yblcdNPcqy5igMx7FuMcz
q2WXJH3TK+hyutivLEmcpjpTYIysZM6Q7GE8X/3+APditT5mjqQ6MZFAQyYBftis
vcN+GRUo7vvPnT1OuOvqF0sUvYEB9v4HHPn6hgQYMhvpq/K6FRYX85I1lkop77R+
/Zy2w1DQOzcCscKB5YW2lXWrgy1Xnvbe7V5HneS/CBxW5pnralqolNDkHe+4gWRq
hh8KuGDXPRjacDprM3PZX5et4jNnKdJMpVGV3kUqR9oziwllgLh1eOufjh7UGC9R
3MbjUtjIb1d9yAvmVJTWc7nCvgaZswEp1EhXTHuWTAiOBUlocOEfwYKrc1m0qgyl
cGCmEEcAbQUcunIelyokTD+V4J+qxrTJz83K0IoBf07S7lB3EB7yuQVOHZpvC1nb
C3JkEXRozPzGCtgWYDIP8duudFz1LRN0IF1tDHzdyfmON0e2Z93pzW9XwHnSaVEQ
A/fQzcaOrmymAnZdU9Wj/WG2Vf3G9N+KjO1UYwGhfKY6kwQTzmAXbvEbOduCului
0mMOuObz0PqLG2C5H1p2RebeiLE19f97eJfOrO5zBR/cTjwQN0ij+6trkDfhCD2r
yD9Zq19naHX3baHUSM/B0YZLsoF1Es45DSo+K5XXHect74JrRnGSXKwzrGUoDYOl
N+oUuMef25q738LdonJ60fRhcg+sfQYWeIFw9GhcrMJbQ7pwXErfQPuzlE/LQigT
UiM1rULVaJLTiWKsQFWhBimN3/PmiHB57B3V55rezcTqoYBwFHy60bbraFhEGGmB
JBGoXrBwHmUdYf4+orMHYMgS/jhCkt6lkRvdNgv6Qgk9EgnR/0Imf4pUn/eIbKWi
g0ApakS1f0h5toYl8qzhW9in86MtgNjKFxGjlcfBijs7wLGobvu2EI0kq8qUhxHq
7L+lmwM1m2YpYc25Mh/rPXUq5+mAzGuGNw4fnpOKf/jYm8glzq2XYO2LTHQWMLPs
k2MdGuMZpnRCxDRNZpHreoMjruNj7RwIxFVmLLYjI/qOtisqDA2ZCDwXBbEMYcwS
//urHC+97aIC/aeg9LoIfyx5sjnRJi0y6w/0+bXsoswNMYsTp8tYhIBeVBg4Mg48
f1NMws0l0CA2ax5EI0zPQk5evLqtbJrojIddZH14N0pOOIWbWr8Cht0mhmlhzDVT
Nk9mB/dx12bF2Ipi8fN2WuTqqyHLQiNjVXqoqBYcqZnyql4r2qq6JthiTvYNrcCC
IpgAi5Q1V2i0ZuBiq9ul7Fei5VEbLPQ1ILtPlSwm2YPFqQpf2KR8xz8qVzFnZMkX
rh5v4d1yS91Dfxf0S9N0r8qENs7K13PSimCWFZVBWRAF1fiXcPKLk4whkgq/7w27
Nhb3IvkzIeJqp1ccOBHO0OHj65Xj993SVz6EdEnl4Em8xILxmfkUddEguIP4/bQD
E5ueQqD7r5yohsYD8KLcJmXiM1k/I629vxIyDZQ07ZYPapjRuLWzE4jIiE3KhOW+
9cnTExNnPT1N1m8zQx6zvwCTaHiw8EcKWYbgjE9R1LZEz2wPNlDe6swrbDAvp8hG
QebQeG9fA1PqrT/M3J4/ZmI79776nXRkjLjIJUPZC6F99vRuhqC5wQU2qF1jMl82
sGQE7sf4yFse1eP8CCTyKDWg5BLuv3jafi7jsdYf+tDyaPy93lLUC4P89XEwhBLG
AzEVh4MaZT7meqibB17W9DicvaiAiX1LegVVbWsxZHeTNsKlXYl4n+CtY/qUAeEP
10nlfkzS1unioTBGoC8T4k8rX/hLRE+9ckfh5dCXHQvxYjEZ4OD1LhaD7tVMo5dz
Ro+k4M74LAS7NIMt2Rovo2ICn26q57NKrvUP7eGUXwkdhKAGVGWcgh7Ukix/qq0u
eBrSIglUF09Vpg3r/76nHtx8dbWs9E96LW1GVCbsFWyuOpO1R2UANj3UDiHsoQe8
pVQH/1oKZLA8pTFkUX5crJtwiYjyvqzfQqCCdqhtCdVyZC37BeKVXxrwQh9Tuac/
4xYaamMBANbV9KmACrBO3pR5MVRTONZE3nSDKyyoRXvOb8YjSeTMwEP5H0XftKNv
zFkQYoocOQIo0F2/N/W71QIB7Q161xkh/YmTxuynEDdncmYZALXb0LbVojAzjzqr
Uex/+xhbvY2fKNQzFHmv6v6AyiRgdawEOpXwfNDBhikYdWqI1bVNUKRAK8mUDxSb
UFVCh879yz2yb8luUODCy3ch6O97R+iQWKq45zsTIEQRdxx54xqq9cHOWxqkpTA3
L8k60Mi9NyhMHUirdaYEO+Ix9RX2EPsHnzYXJBVlXXoPdBa6zan3CfZ2wo+uvtrg
1sheM7H2efAbopsZsgTQOE0YQxeedsHzQb480ceUgplFOzncO1bUf0StEBACES+k
hul7j3l0XG9SEwhGfi4g3T2424MB04eKyJSliQYjISLmYAxN0A16CiCyiIBMWsxS
tMCr2FsGugIXJL2usCnS+GP+4rxHqyIGOCUhEYy0KDgjK1satDtNAQiaZi/j6cQA
Pq+hW6906+xa/Nh8S9VrsSe/jJdBXTf2qkbJXoG+k1ae3z2xIrx2ElSTgsWGmvte
gqh8hE86GznEq8QqNs/7kNfVBluNb+zMVTW77WYW07Y9jExyhhiieSR/NW9yXoxt
fYbv2stsHt0U9VmZLZVO+Ig3T258av+dW4OK9FupGliYSxNNTH0mI0exGHrkZEiZ
Zy5LqADQDC1dyMeylH+rg6mGQIilOrTb4dEqreiHflCd8oPbcD96FLRAyriJQuPN
oAfB2sqIgYL3j480f4MPY8esHrhMo8j5auRwJclK5MFRaxMpo+UGXkcPGhjiPi7c
vavil5AQZD7DbN4NJt6lbNxT5Ur6B60BmYsWlVLrs2uqUp46/DO0f/AsAN/gab8u
AS+YDOtD+RYutZu2f8ogEeAXmi0+zvQ6mKm5YKE7nHX6QhFIOgQnYnBA+AFLqcbA
tZUyLzcj2Jps4t3Im/oBNTfW6rpr/aEh5bmPCGJ5NZB0HhVm0K9m3K+ib0ob0C7I
rYQATBUyrAvnSMk+Z2TiBv207C8CZ+m+isqhhwkhaTnpBrmoQ3xRW41TYUOzPaRU
CFjofk+yMYlD9imCD5lJ2qUVmtJyKHM17ccg0DsAdVnw/h7nq1kxxorUtlAjpMD8
QrgY+AJTt42QsBVruVpHFhpfCK58Bug5yYztzk9CsfK/185QZz4TTUN4PImBBBGv
rAEuiicQyvIJinrXDX/FsjxGqB6o5qqkgx7xLPaNeMJaO440+I94mU125u1rasVC
jVNS/VLWy3+PZ9SATTP8980CevAc7dcIYISZgvZ0EDU1zMMhWhQ99AnjRuSwVW7R
zTPK0esIZs0m4HWgFjWbimNMIy3nC/CALGFuy5PsUzPAZHC1dK+rbuQ2Z+uhyz0U
u2ticIiIKy++C5PFjpngGuC2c+tgQbtIc2nZxs3udA2wrcdqh3jnoNmx5S03Zmvi
qkORyDbeYlUpoggpHxp5pMlu7pJdpVyObIpz9CWLu0KegpwL2ZR84eVAuh8K+XPV
BK9Jj7v26jLY7IBISaU7HgrO6wQsjQVcRlJhdookynYb9jRdXWIFW9D53Y4idO56
4jkcRUzjQT/aO1MEgNQHCEFTXqK9WQwooevw1xx3e47UBQBUaC1vtYdu+vD6rzAU
YrRrTJS5C2rgVAR2WrAtsPGDv7sPj2cnCLSnFXnAOWyd5JZNn/CGA4T1gt5gOYvz
R3G8wIs/y/GNhZY4Y4wAJBAz6GEU5I9/E7w73WdESR4oknuEGfcoM36dOXN0o/z6
aj9z2t9DOduJ/u0iTKlVPFV/n99b7Sreo06cHyk/qLmrYx2TmIXrUyD6/OGFPycA
cEtrl8xmyCGzVs+7Vt8kd6mU8ItrNorQBsyGb0bIq4rn5dCi/DBWVDv1fn2S1LtQ
IK4Woe0Xc2zgW27qwDL59X2PdN7Epzr5DGOn3kKE6ljcfxwhz4fTgGq98yqYqzcY
IAij3KdizlXIwGgLy5bzN1UQCOzwMDf7ko6Sl8WR+xwwyOxDkV+akEgyosO1Jt1p
mFTJseT/gv8m5duZN2T2W43ClbUPsybKhKyhYZdP/3C/Ev/uGUJcKZfFrPA+rZOz
qiyD2qI0bqxUCHWcZvNT4DavppaduAd+kKXFk/dafdxOU8UScyXhwS8Jo87XQOpH
jNL39ISrHPpwC1M1MqFJhZMUnOMya3lj86jRwNjrEXsyY24vwgizhrcDuoFspflB
t9oHlWNL6GLLmfM0SA42U8jcPk2DtKC+Y4QyLIBzkxxCWvptGbBs37UYY8OGQH4Y
pCFctxCV1tiM/JvaT/CdX286Dr17b0XP3SATtG9jA3NIIkF/pCiqSF0W3XKMXsaC
bgCT3mQXqVFSlOeH6thn7IiEnSfhHTfVtD85GBLxUZEWJU6AN9C9h2OS5uivyTOU
mgMV0Dcfd0Tlb8O0j3G/TvtIzydwznX0Tnh+dheef3t2nmbp3sBUlGH4LTRVfg9s
iFCuV6SqOdt3IcsmvcMgJFNL6GlgDq7FNSg+R7mieJk4FVdBRaZrldi7RAqJRW1W
d/0aTJeb8rTIjULQlG+oTvRT1Lhyxnm4kuSIFwu5qWgk4MpelZo7PO7jzIxs7AZO
MX73MnDEOVoOk59YsgndmIaOQIXvNB+8D+mU+fgXIAOQv27ZQhGANWMfnidPIap+
Y0TUwjTUjEP1ipGiTQCf/TCRGlzHqX2kTvnbY51rdYlXZNRO9LOAH4JbVLkvtbfO
f+m5qLfAhiTdOlM72F/qrsim3mIln82RkD2gn+5WlDB5jk3UXtEPQx4UF4ldAWkj
EbbwhjKfvXU08vCB+0oeVir70RakHUTH3vTfFTyPVTaPjbPaJR+85/A16x1/Z8j/
4aqDg4cApUVVC/UhwKjkBaHIjNJ7MxwjbM5OTLgMzybNn2CvTccf1idpwtXfkRes
zZdpyJ8xa3ecov3UWgZ+HNMMB33iIIL4+59Dh8Oy+KWEuPUeXFWIPuXBhoo54s4Q
in6Zm9tAegM27TYeww3MgQ5qM3d30bkm2LYjJCauPMf0TdLqq9EHje0ciU4wHCq1
ibCAE+nZMiXUfnXp2iRtjVMDC60R8ITQwWwwDe5ktnZXsMxs7z+LZVcApmgvDSND
FDCmuQqZAwo/LgPDvUsV73BuCA5nRraudvrIL7ejuOGOZ+ncnKyMCcnQBwsLNV15
4yKSgmpopswbSuXCt2sJvuQRxs9U3tSTJA9UWqdyLj24bAxhTbJKZ6+M8LQgZdW+
8m50vnicKRjozKDybgDyqQEswKCge+vycip1Bimxt/2mg8tkqVpMVcI1cuoiOdNA
Am9EmG5+5S1wOHzREUBudtdq4ku5SPbgKHu7m9raqqzBB2fYOebuDejALmZxktVL
aXFiQCM4X09NmxYv2/7dNUhK0F/vxbsM0UcBcFCadvfV8CgqLe4UxlKg0J/wQQbK
a/ZZTU8pouHFKt7XMdlrGy908s72UV03vlL25mjTV+C3HgxtOixosAPe2RTwxPjE
9MGplqYKvYYyoixLT6BB7bfDX8h6KPJn8M73rCsZx+LnxaMuDAsAyLSVSpfV/Mj3
P4qG3h4iLIFgThQjBt4iKUYSAFB/d4spERmzUgUB1rnm4oB9/Wy6cj3KJ6FFuw7C
GiYtwUrwJfAKEh5cXDf6cOZJcFCKfw/oxxCcTTu6TGWD8KRO48zlzoP5UEofzmVg
ZyuIMDv4H8aPK9YtkHgA8dsNyByfP3JwrtghdjH4lvbBXLFaDmqJuDGuVOMDFLTB
tC/ybSphZShZbhj6B88Wb4WP08JN5xISoNAVnaN8BbDmDqRn2aXynQF7Kulr5L3E
TU4yuDBZY1/o0qTzzDl/zRjdteAnX86Rp9E6Cg3EWzQRse7OLb7bWf3EZKAkzFbR
9kuI/PTxhTCSqPHZdyxfPnoR0+iWvcvgLGXKbFkqgozdFnhQkDO63YBOdxu/9caF
fCxBHSpufobtOaTP/kc0miuJ44LSqXdFX1v3bVbiUvMQlzupxCy8q2ErSqy8pfs0
khOtmeqLqm/ITiFOkqbXbAXMOUb4Ufqq/r5ayZ/WdWTHGXAeC3Ja8PC1CEjhBcSI
AFX7ZSUx6FDOj+qmDTpaRVeqU2BQKEVMWNQM47wDFzcEdTorfYC/low50AJoBqai
/EZtG2vpLeYjHOdjeInq14tUP4mR2QJaJo1Tx5zb9pws+ABCUFAvr1+8fPDswe6g
vOv2rfcmm0521t7KVZU+79GnPZ1K1aqb51ITLP+VU0KdfxoNn5Be4cbzRGwZdB0Y
BzENuxVPOOkpspPaMeyLizjmOkGgt7T/JAuXm10PeVl772sqJXmeJy7uHt9SHuKR
jJ8X92gKU64KJWbRYEoKN4XDFzkK0hN85Ps6cbqT4vxDEbnyYCrFRz/mzMv6Vdai
wYmA6FizBSPPxwhT2rB+3CI5TLoeelx523u1AGUZ2Z/rjsCzwOO7Heg2RYKN09gW
hoBhtNt+C42Yqw8jtkuOrzLyXzXtGXLEAGjoJS/wEbMZCIsHbYZ75JvFvjaE8DiB
gniNQcilEgdnBub3AS98NXcCNdzafqlLcJ6e6zRsD19K0Foa6UW1D8R05Rp5FYcE
vnnpeAaPGA4SJpExUvURgFJp7YqQ5sIgv+E1XduPOp0eGKvUBmvBdnBLd1i/udHN
xZVod/Gu90EK63nDcv0cR2Cd6L6XF/95Ad8BnbhEc9uqxztcGfHmWUdcwxw6CeQG
1+OGKvSiRB3tKRh6ZykOGkGQwHSSZO0XE73WQpfOZMY3mjAG0ghWqsZHwIvNrJDr
rkzQEJyFTIQyh+0n8NsSp1ziRSbI09yht07Uq4fUIIUm/3rbFT9iOMm2cCB6wMlN
4sJMp6sqcfUHT/AuBDB4vxIdR3+NjRTHm6dMHhiJ7Qs7azIvkYaHyB4Eljvrm7MR
BRkSOOkpRljLuOckBg2WVENXXxyVdIDl8c8tRsMoKEq06KeYexer6egVmtCOXPnu
vpRk4Dt7YDVxeAG4qVO53YOorbXkMtdwRNfMfbB8xDFLALLwDdlYIGpkFeid2bTI
BTcwkZYGP3siCQp25dYv4bJN5fyQd0izurqtbMAQ+ZWGhPxaZsMo8fwPF+fT1Qqq
t0OHmCUhvjUS/7LaOjhYnmZktUb8FqRjP+iCgwVn4/u3RQe3Msvx/P8icnb8q6jc
8RBpTq8GpDF3jEBl6Ql/X/TgezEZToesRNDcVoSzSiL2TXrPp1maib9OkMARBQC6
b6RkOwD7s9RTHJxadbsi8fQ/ZtzrAqrHivuVTF5GpEpumkvDzO60iIclqkfv6u7v
2LKvWsYkygU4G/RPwAwWJ+I5JoL655yYlezQFLxHn/HoX/f/WLrfqqq/OpJKpfON
WXsCVDhBh7IeK0RFMR8dGvJT0HZw0THKvxEi3Llz01eVLU68Zkrzw8ps88/oROnw
8sG2isI9dwQbv3zWxuwlKicGh/1pPx7ztI76SwwtHYQdBwjgq2Mn3dx92IbMApcn
Udm86THnMofZunBf6yktQcYCt9e/jk0cVABcSlxVtuadPiUtinY48CM1Pdn/Bb9+
PhliQBgnua3Nwv2qxQiRjR6t6Pk7A61Gdx7+Jfzg+8TJq1N/BEgVbXpSl67VawdS
c+6z17jNVWIxmqL7wdmxRe5HNj85It0GsoDOK2vjDLOyQdGqoT9RmBeY6ApCaYF+
NtQ2FoG68sp3S16d3pqpaHfvjR74cTWpSXLPWnqxQziBtw4Z7+Is3ES8DmHq0T15
LD+4Ks5gT5xx9923dCBcw8bpoZtdL7X5Ti5t0xdvPGcIsussIElFtuswFw/Zfsc6
FKM8rJJQU9i5yDbutjU9YUB6yfaC3rAMHrDo18gEuctfxFoo/qhwcV12VNUh8mA0
R5qW5Puh1LgvqV6gnk3EHTyYre8SaoRFH84BgZO1OWg1T+G0yh501zizz0Acw5m+
44f6e9jxGtDVbni90gAPyCzzrI1NFCT8rJtrM0UI0AQtniXSKg5f7Hp+VsM/LCDh
JKto7dE9csYYhJ4WJPqKlsNBVmeVk+wl85rGAKvJDLqAB+OkS7COxpVi55eHM0RR
8Q45atfMoU5b3hnfaX2Y0K6T7uSLguIuteCwFK4L2EUPiGqy1dktPcxRZO5N3zc1
fLkP2dqgK2Dz7IohdLR6CU5CnNH9Iv3FE2Lq8F5nBj6gItWF/pluoVf2lvCCZxzS
273SDoTZEZPamRrbE2+UMLcOgAzTGaR1P+4Jqg4t8ThsnLZHldcECheKfWavl3vN
RcIY+mwHfr/8CYxRjXTMrM6yyZOlU4kLmkjMoeRUWSTsM/zOhzAyWYNWiT6J6UAo
L7yev8/z6wiBD/flvkr6AzNQTEfS2TDmTfvFPy3lHIHSOROQIV8uXwOYGpEV5hLh
z6wdQk5bQxzvB3I4AMAFfpsv019xyDMl5wBcz6CHSFh1E7+SzX5fB40Z4KgAON5A
eZiDfjuntPlFGyP6MQtQXCC6tCSM4RWZr8+v3NheF/KheH/wGkYt8+Ew0dIRsgRJ
7Xcyj7grQ5Ui0bbteoMG6kxB8SU9PBlAr8rd2DA/VK1i0ENCQ8zdFfXyMwWrFOUg
NCKzjM9ipYHW3sZXkXE30So0uK0Lv+UdDm4x/6XY1oF0++fAHv0H2c87hYiWzwyE
9GkACoHq+5ziiqD8RH+TCgZusdj9scqVZuC1UmB9MRApG/+vFyts0PMeck3nnXuh
MOzzWKMRtrMCClkUEAXi0Jxb8M0uxr4PaMJBMPNjQImVwPH2HVUr8Wzf7pUg5wL2
F1BKFDAV9oj5BQ6+fY78IFboyCbBrrXKOHuQfIUj+oXy9XwWbqFSlvXdXvAt/V3P
IlimUOmoKhqrBrO8/a9/rGYocMGx5A8UB0gVoKwOWdRkpfxqwt8brd86w7Tar6se
QlELp/YzYFA1I/I/zLv5okmuN3m+sCf6GW9x1NigXz8oN8XgaNFvNUFZ8ksQlCPk
PNgfplNVW0D2NJtOIs2Y5g5bZhcAgQK2neGNXMgfEiIZPj2tBQ59mMpFzm/HtLkU
bCbnoekRG/MMsuLuUw8kPDFMh8Nsz2PeNN63q1wBmlzsstdZ3C+UfJxauNuwOSqV
0RRLqPxcR7jDmJJ9+EBvPx39GK0wvt7qdYFng5fnoWu/Cux3K+4qwD2beOqe0MEW
qmoJK5HbFhBIDw5rr5dNvl3eqEO1fw6tww+CYcyqqF/qZNfzM92D9fbpHvtc1s30
k6FJVH1Ydh0tQf3Vd66a1Og4eGiMJ/mJAhUSOhsxszjvYft5asjCKmkQX2pNjvVO
Hv/NIAEUpbpgi10JAsjJqmAYwTvAfsLYiMTPNAy+CQZ9uOTOMdwpmaY155P8zxlq
u108jY91XLkgbWECPAjZduXEnYJC0NKkaZZOp4zHHIYlFcaNxKP5SxbwYNIAsQ3j
o2F16dO2cUsFmLy65cxsgQ7EF4Gt+PA5MyDzf+g9wv7q8l+mYH29vtC8U5CQnIeA
qaIKNRbftBrJtLloJhL/E7mNjGmNA+tIsj2wxyFpeQ1whqw2x5ZpCcaicpsu7jSU
HtOy/EeRwsD4zQJHoK3bYrYnaMDGdkcb/jsPZXRaDfvWnrh33t0gD2DcKAbfdbjO
RERcIo9hJWNWK1sLKZBVWu7LY/BZjAtr2LvBQvCFiPoDtfJbWg62me3nEbY9+gk/
qqsAcxmtRSEn55oRVXEuZRuvs2QkXk8FOFlk26WhPsf/9HBt4tJTVWTQOpV5+7RW
rTZNY2A7YPRj7rCtHXjEpA/bOHYCCmQ+rS1cys4iie0nceSQgVzMBfBeN2GGPleI
MFVH2GgxzlmBYVvyjGEtLIynp9xdQ1/dyDPoz0SAQ3JZD/8H9oEP/wyMODrQExe9
1vURQpYd5KbJaeteiFy9hbOiVP7rS9l7d+0oBkdfefnVOg0hUTx3q2aELFoGXn0S
Yyxkgcy/ELbtVjRCijcqBWroXeFX160wgQ09FNs0PtkBs0avx1J+oOd/FrEb6oam
UdnDyj7P5Dr5D7UoKH6QF9h4QBse9hWvBV8djcB6hvJ7J0Fc2BuZKjMtM/Z8R8yE
fBqZZQVtQbs6PhMf5/kVdrE/+pJNUpqYI8r1+WHREXEDO5/xjU0WSh2Jn5DzuCmw
QnxGjpNX0vranIURQEIXtwr7GaqV+M52ERSIDcpJ45xunXzzTS0G6ZBDGRs0yhut
/14dWugKW/M+ZIgst14xbNqP1QhMxsy5o1CLFTP0D0iIMvTVuWGNftyvDbyoU2M5
fExx+e01E6tBViEzDEzlaZD8EvEE6AzsWpG56jvs17d7yak5dV9NEp+Fw5ogzXmZ
r1gjVhESyS2dFPdwRIgTHGFHXbywRJpALm6oWrW6i1Q12q6JzMH8JzVLioyqaJVp
bhT0JTsFiAJxeyBxyLoPn/E58OT2B42RpNajveEpfvrK7/FuZUMzTeiT5qdCn/GN
deOvjKL0x8LLboneom2t3tdsUef/bcsjjAcoCZYTmaxMwOEPBcSOstkNLs87zM7V
GQ6n/VC2mPxdfbzQ49UuXMhNPBpe4arkFrKKDmCr5Wh8rZk2firFs1CrnJE3AUue
eVpjPN7dZ7ZNz9v+p992lhP81G7M+Wo/QWnDf/vSYmKSUnc6kaZWxgUcHNaY5Dqh
Du2jEu3fiJMgLILeRT7qJdz95uqpRlArH8xVrWMY0KT+q3/+OTZq/jY1L4nEcKeH
l/3JBJ31J1R8WBfK/ou9J4J71V8OKDmO36V+seRVMptAlLRuPKiCx3MBe2BIifUh
DM9+rSEiEuF2Tbdv5mKhEBYjDSeaYM+Q/D1oey+fjsMd9dQMqewe8ygcP4BszuGj
z6YE63T+3Jx0FvluvN9/ppXLB0ryMph7Lq9o1qGkcH2Rrcls3YEacGZMe8T9tiIO
jRJqH0z8xNYuF8x5XFlqcuUfNLNgfgWlC0ctvzClWrrYJK1uw/ITdPEn8Z6GZVp9
jYLriSnJMAyjanoz8V7JhS9ZHX2nFg0a1G1Wwi/qe6P2RMJwgkCb5pX2EzsuK2wD
IM4P6SZZR126aK/Wuj+4DdzfDrG31LvD8bBLWHBD9XaXKuQAccMh4XMpNcXfR/W6
OUxivnnmkCVM2x9qmJiv6QEOasAHYD399EYRU2AgmcRdjiHifPbysTO4JSrV2C1J
xhI2V0khVMIbTnZszlnNCl7SZEA5yRkzADhY6pxnPSIPhcS47YhjFuqcmf49dIoj
AmC9f+l6VFpqM+evQi/VYsnNlaEw5HxXfkrt44mNRTi9paoMgtHqbFg5qwHCD4Lq
Og2LlsKRwhLO3B93JGXagzH/iXLtCuPl66789sRVq1V0MZjIKnEj0R0/JgQyJEkO
K/5MjGYqlmojxoPThm62GBBAzIoAj/lbQYq/lymGL7KbF5BQCl6DSnEXMCV74hjN
eNKDXmB55IlnJzBcbRm5W+Lbv4qXmY74ptGCa3cRAFoteAzfDKbU3Djsh5QKjW02
uI2hSSDpP5GjcbonQG97IOwmXtoL6d9ubPNmSbXDoPE/M1yTURecZRqfZWYygpnD
O1gUDOMqoPKnfcnC91AxxDzWhvhxIB1qRRGf5do0WsNvye1iNyF2Sl1Q0aOd2n4K
Krbe2YP6TkmT6jsqW4TmeGVIvm8HirIQ3hpow1q4HEzfMlpNisBUI55ledtpUUrP
Rf3P0hjEn+Iun9IrViZHR2QJoFOs/R/UCeCkJtBwYVqRR+rWTn4Za5u9HEUvwgn/
z2fuv4fxjHyhorAtkC26gQlZ0rE4ahqNc7uS+eqGsXAcHkeZwjsQwU41Tl3o1AFe
Nt0JFph7o5bqONCf5qpiKkwOmXDfRRw47412ij5I9l8XccPOjwIdtpPEgnB9XNP8
XF13NkY+v4ZCkTVzD5gXtBsT7jDnaULTgjxMYaZIc7oPN7Q3nIePE+5qg7DvEqKC
Vt/0dJrakL8PQPjjrNaNYg09ML+K6xcW63CXugZ0L66XMOdqsTQ1eB9FJP2/+kmh
m2Sbe4bYGhafKcgCksqN6wiUA9VECrfnYe2Si32Y6n4aQMSfj2yn6kF2RPG0PXNK
sQj7TNkpzLwUn7AyXrwQoDjSyMhgmopyVskdPzZ9XkGwcmm5+udclNCpEtuPhOMh
daYxbUyIHqe9EvJo0CTto3vgv0JwgRNW3SVcgMW1VlRLEW3FLXNZAyRHoEJ5+cEf
GG2J01Sw5PnVP+6Ji2RDazv00eGoQXDFvMWE0JlwFUzokoEZ6cpP1SwA5E9WHZ3Z
3UVoDRoD0tvAH5QAIOF5ORLURxKky04iIVlX24ZnkiwcNTz0VImN8XTCWxj4kBLK
DJfPsIltCGVSRgVAV9VUJSC9eIr7snBf8rJtfP/SXSjb3AF+dwLQx6vb5QAw2Z2f
kJ20PKBQVWc6yuW+lmnEkMSNy7NzA4Nhk51yZN3skv6a4qrqN9sZbGroFBZ6wC37
h/F92ibls1D/KjGDE2t++l6Z9NGTvntHhrb/miEx289pxlBOrSeVjOe48O91y9w0
vK5DdrefIfF8EgFyQknnLUtnAQcW9u8XN5JyFnQEzNzisC4AwCOWekgCmmbV3Fu5
tTeLDLX5qHC6oUx4C1ee6QlRp+qK4zHWNEN7/Csns1ZEBU1L6J6mKNJAFcpK2U55
9TGpKAxTyWGWRUOSM/4vFDAiRQxoZXPo2WjsMc1kelvu3k4GejOFbIKy+VA8p9iL
XoNZgGNpTN0RNiy5mzvka2y8AxY/sGYa4qFFMsok2VR5a3ha9OolZqcAePDgQzFe
LbPN9OXhFZyJ7sBqjmelMwom5jYEC4DtKbVurfCdGtB6OsM0/jFlqQ/9vB6aQ921
nEbfS7nCQ/lR+RcK2oRKIk/KUCZIrFNK7mytH56Up1SebYByfe4rsHY5HuxcZmCc
vrR2Pgtx7D6+Qkht5qJ+EedajMJxUZb319ZLrLEhoeE3FkbPA5QseIltfpgIMxqr
nh5pCFgGdBloFm4X/453GEZ/geV0PW4Q7yNWhFQLw9j2zLJo0LCZSvvbRxABnGg7
pxI+4aAaXUeipRft/6A1hc/nNJziqwK+pqy72MJT1NrLbHILkgLQtM+lnsX+vq4e
fQtnUoqp/Po/A0L74XlFyRwvfBQhq+d60FtyyR+uYI7XLu9+7TPP8t/T2Qn2kPhm
gj1HkjYqxOuf7P2A0NOFj2WkQa7rF0CJLkcgDH83TTC4BgKjansuFouqG/+aaHEA
fc9a+nDmnJIZ7MK/pMNCQwHM4+58HBuI2yD7k57fWIKydcdAineufL4EprFkteoH
/Vr+1W69YNrgT8+CRi2lS6KBnpaz/4+/Y1MwbfmieGnJ+q4JRdTi0R8emRURzGjB
mXH9XRtI0ezG1HphB6bkaNx3lsko3Y0mKp7GNiINFFkwpMFQz2ANeXVIbASdgVbB
pu8suUPT3sHnbTHmIhACqAf5EN6548wFjWTx+lB7oOm1cujrV1Ca3gwYj1GugPYf
B4mwjziHuMjjzW99lEzivmhseyDAJJHV9qzKZ+Ro5vRujZE8PvdWCIpQDPIV9KXF
KzkHsq0aEOU2Hh9F9UoirI3p7QEmfYdIGDz4P8dbyObiGttfaJ7Lee6jCvvVZAfN
tii+r2tL1cvRYC3NPZAYsTMc9kgXZ2yzmdBzLDTHukRKS1heH3JXU7Vg31oTGGxy
t/fvlW6LCwkhKb97/e5JMY+5HAXnVXmHihQWe4R9c/RfvnP9aCECTf3kg+rJoGOK
2bts9xPJmF54F6pE64u2BKA6a90SKVDTkzjzg4eHZnGGvMHwKB/oJr5brTstv2Mj
8HqXNqhTdR9cVsw7Kvc+8LYDDzbXDy2CjpibioOBmKm2c3Xp2um3g3lUYf2lfvKj
oESQTf9cZ3vvNOxOezPbHsmEObrSBzdJsKMhDJjDt5JJhA3FzUdoQPRl/rIIhoFa
2icuPDusuR8ETWv7HKXlcnIcm4fbdT29DPNzLrG5u/Zq4Z6xGefsOM+HoLvSPrH4
CiU0RdkVbWqnpPlNGG3yBPrV/ew5dI1a5oWMGBgIRljj/VU2leu5ymBdzq2CWJHl
QDiptpBAVO3caPDLZ77YMKUgKIWzfVl4y8+g48o6p62YOSP8O0v9D8TvIHsgO6EL
aS2scCmrj6jXkJICklzCjFjTaZhOsqGTHUXNzvVZ6ADpNMZYywd2eedFseuG4ZoC
iUtmV00upvSFinFOqS4pr3clxHY5o0KQ64HsNqKK6/qMxIzuRacso2xvEtRJxKY5
zNan5Y4b3bdDA4MChuuYDRSMim4orwcuSqhw2sxg6+wV9T0GhST/PEsEHbTgL54u
cLTLvMmi5CsEtH9DB5J3nPbCX0BrenlVSxK4QIIyxZzrIhRZtuMAfy+UURGej/le
aOVbWD51/QIaysSxUwlti2w+lDSgVqJgpxkosMkWAeCPDbAUXu2Cfgkxj72Kk7yz
u2VnSQVFyQYAxXUkhqmfXQcCIodeWO0a24d2y7T8xsolZu1z0nkEX//86FNiexTY
EyhCONsz0OULW8TfSA76xNblEr5ECI6nY6X83U7SaWC1sIHoVfQp06cW3KGmtQUJ
m5PqzbipzS6tCWwffLxGZyGkgfuR02LL50s5TPaSoNVuabGfp3j2pyxfwhxBs9N2
iP6R3kHcRjAXaDcO55O7PaGDU7SYjv/8Mhh3syk20xQxhxlKAmQVeOKLG06nwD+b
kpFF1xgLCopmTn/qpmXiDirz9N1DXQEFXaV+rfc+JDLcpQj9Sb/XmvsFnuX+6D54
Uz0QR/WJmBW8VAibFvdK/MeX7E3QRLLlgP7RpqaA0V7b0Dxfv0SWXL0VZ5Y5NRk8
ZHZTqyKT/Gn44TRbGWjPRqvozKcQ3/2tppz2F9OjC5eJPL3kW99+56bWexOTzmdi
vMHLGK6EGazzIiuo8V6gffJZT+86ZxH/DptY1/bjwtdbJR+Lg3hDs3+qXr9zkHaa
EhSp1zEXzCdCkRD4EAuvrlo3pJ5BROCW9YXt9Q/m/CbMG5eV/eaP1/FK6ykRCuyL
ZfZqL0pLUlFp65u8jlJwCXhhUc4bS5kD2FuwBI5AHG1sVsf/AYZgy/HrtexelwbF
t/+CTraqdFC5oF4IVuoZckbswuz8yA8W40AeTXVOtY8iohmHkBcpFJe3oQvWXrnW
HYFNadGXiBNpXHdjnUaEtnnXrfYRlOFmBA/ofe1HSWR5ZSw3oBhee4X8tU/BVYau
7lUIwcfzOhL5ImtC71ugaMi4jmPRaGPNhCgUSgBM8OjehJXoN4Bn7Xp8d6n6oMuM
uMnHW/nH3IMGWb/hrshX5QVCODnBTNHY2TNZllR1m5vu9KVVzqu1ePpYDV/XHOFE
/k+kaXFCpBC70UxmTPTWqwfMIN9+EmyFCqsvk4M14R4YB8Q61fbacelUcxNzvHqD
Z6a1aEKtlY6Kc0gy1d0hBtMv9ByrPly28KbF+k2IVWgh7DsI2R1z9AIOYGgyXAPw
eSzvtnUM7U9nd8AItUMwRsu1JQtBg0bdmOVlrX9rPCDD+QkGT+d4YO4E3xxmaRNP
tsnmgEkIIieqhl6Mpn7V3f0C4cGVQpXx/GWdXGY49KXeOFJiRLwQtBpmdyFTXf/N
sGPCH0ihsuzL00Ub9/WYTPgvLVugHQn+m7pq47xnMvejiGxtEKlytOGjRifS0R2L
QL8ejZufRDdUYNSgnMcW0xcnxYGJZ03h4cT1OERPATwMdVgeHVpFyLCy0yJ0iBId
9rGLMSpBIGX3LgQvT/DftOZf63BpaDdFhjmxtn+ae2H+mIHSx6HEjAcCgSKspwm3
6f33cqTOX4qc0T6ryDJ+Lj/yJlF/SY0ugtvfvmENVOiYrfGB8Yrz8oGp848bj9Wu
8TOBHdw+iH+gEXg5pqyuBxbZFle3KNIaczFqUk6o8lR3ipIj/ZhCVIxF/FHm9uE8
gEKTy4jHMItIuEvFQBm9ux+xm9P+u/tPHhnYokRnrmjfS3apuOxIXE2Zd93UCQfQ
kmZNff/FTeuUiVmTxk5SAHAdUJd/kzgpEZ/+2YOiib4oGRAVijrteghMgfV7QAhE
wijvNQON1xVPw9qT6kSS8bd4HcmK8rrxNdTAl7PE1xM72avKzdlvtMJBNxHWVQBb
6JCL8Vg9rXRj1DmNkwRveY9UlQwEhDSODrC9d3Sy137TpKzu26NZ1VxDkzMoP73f
KFfjtQLPL2GNfAelwfTKWTr3rHWpiWUyi5xqxevV2NjueBjKCBjmmjxdR4HYgs8Y
0l8x0P5rQMBe3jlIg/bc1gWPOnvZ7bGWsoebIvC4GtLjN22XCH2K+qJ9NH7Cml8X
zB+3B8bTIcWT0nWqF7tQYY55d+tgtrMhJTMqqixLWoVQBgXDt15+sEcJGF1yxcro
Rg82tCo14GTwFuqimOo9OuFxv7esLOfoVCrC/LNox+KMogw+Iwv6D9C63mz+eI1x
e4cXi2EY+HoWQclDojyEvjKK2gPRM2zCtR8a0zjaddrBiT5WD2++tr/VFIfad6io
ccdRyYxLAyM2e2fKHM35Py54hLgPxrFlZXwj4pUdOaHNDqWLI1mbAqjbu+sg8out
x+6kbZrpMnoKcWOJM43TvPFR/HU5D/s26QROot1cqIiOzmsFhIIuk0QfzPHxlxZJ
azPPNOfSq/LUiDLX/Hi+OYh4O80IVP6y9aklrtp3OPUy2W8cYygNyaUEmeAlSjIL
WA4hc5tU02u04JsJ8VYTIMmmbMSDC2mpExnOcwiVryEsuuVYGP1j29tk9/cf/KvB
CF0e6CkGIMANotie6scNsGSQOKRwkRTLGXbRLcWMAR9msW1PopRXtsAo1BcGgCSp
myXuLQndP1Ro93e6pp1dZD1uaEn49/xCD2I5pp0PmyNDHAKhqIX++2Lvk6tDhknK
7kon+cpWvk9QtafBi+4DeXNODJuu807AbicKSneFQpwRl8oUEqgVfuowdvLkvj91
NLp5xX/d7Dk43FSiduAhlI+hxM2ZP8P0AkdL3TWGp6vcfJ1LeniPB6qrT4k3LNDZ
kxX4o4Uca4zS4fZcy/ZINnjXbDceVYrO6G1b3qzt2N/6bbqUpJUWHGTD7ZEdmR5A
20vYVEk3OIQP6KzLILKjAg22Hd7cMfQ8BoUUtXDxLGIgcl6n5zA9X+lrMeeeq/5U
qf8BJ5KvlS8IX+oUN/DlnX7hGuveF5NnvXJc2jP46lpCN5OqxyMjqwF+XKTBBuMp
VbQT30ZVMcGrNkCk4xw7AHBdk1j52ZmFXZyEJcQ9Sy1bkMGbj3SMnBiEZlbgDuLo
cbYaj2m8/O7C6f8NITQ3mhraDVO/Y+X4srC26t41bUeQdZlqfzCku/m/LeAcaDBd
gXMrRa4j9hSgnB3/Mzdd94fCHoQZlBSuEXXtbLpLuQtrLMNGHd0G/9dPh34jexhQ
ZhaqPnxv5nVaIExOa4XYufsJmUc5X8cMqdhY2z6CUMeY+CNHZFWPBvpnkXoZxCbd
LEDphrmBjQLnMkkbj2bMxlXlopPN0u7ecybYqKzcJJnWfEtnrQsiZ8KPgVk5lOlO
N0hZcpM1eUvOox/Iomue81cRNhqOwhsProXPMcSetm/uQstJz/T9TlzG4Fw1U7gn
JceQIJxeke1MC7OLP06N/tMfcq1VbWWKS1LQSlKbKmlH4gvADetlUFpi3cuTQIim
VqHH+OxpdUX3paV1BhGEnr/0Ao/2RBY+P7KCV5IO44zo4ONjlSkeHuAyr/pNcKyn
8LY2tVlMkUDxVtkyPusmOcYDxX8LkxQECJ0maps49yVSL8seyJydkJDam4ysM7aD
SJ6QtGdXgC53XIa2TVEu8Rg0Bg22C43u5aFfXk4BWvA3Hpyz9ES2YXObKM9Ultxn
EceQtSkq1pDw/voGxMzH1D3z4SDnxvLL64fCUp/V/2KFdeAZDPX47SbLUDHsWtxO
6V/xFeSVg3RT+72eHgE3bXeliT6eT2THDlXBuCaWV/JCOj1NaV2g2RvAYVNK4Qo3
z+oKjNxYRjgWLQmtSApLsj55kvbbKEcy3KLYfrhcTtMHWq4jPK1Eskp9jCs0Az+i
uOtfA2OVrW0t5jtvI1SWE4gp9Rs2b8WyWdFAvOBJaPxssczgGsc4a4g3WqUvZyFf
ymjI8a3rHaY7SNSZCQw0aquhHYqowX5QS1V7rK/W9f6iQRhirL3cl1VeU6RZcswR
Uimmy8ztywi7nmVeS+qSPwlsY3MXT5bUtwe0PPWzYPbIIUTD1CDxeBv8DAB9g3/G
qIa93hgihqEWqL0PVPJG7utJOJDq1higR5ZxeRNX14LOxWtHsaVgQR43UZ+qRV7b
/guqfZ9uEtfvBJNswFezJZ2n9nYrbq6FBlJ1CntvFv5KjNRZh7EKDP7Sl/vBftA3
m5epb4zsE2mgW557MIDtHUb9boslCwQpmWaYOktUrSLBbtGTvXfsfHpurw1FV6QM
E80zXQA0HMccb1qZj9DOGHZcpYXWisMvPv6Hd1aA+ekr55sbiXd7xYTXcE/rEm4E
05zrC4JSIzuDofjwz79+2s8mXyUx3ZZxCvCkJM2vUlCHVrCJP3REAIOrpHgIkYVt
c6XrQzfJwGL3QtVQi/t7cBDY7wek5yf0l1nLTxGMmuGYAb7Z6wBpsNQa+sD53qpq
uZ5UB4KjN8X/kNkY6X10FMvEhuQVyhTxq+zB32ZyEEZD6INbkTrtk4Sp9BLZCs33
WpOwJsf7Eg2GP+nxur2frCaU7ez4L3avUZKoV9JodOqt2ch5pzJ727RfPJRaCVpi
VICVEXZ0aVkMaBDdCp4d8ZO6qCOyYAnIkKH7YH5B5XmNhBcbw8IP7ZF0wf29Vcbm
rycDVC7FFNS3EnQ6Cis6hsgyJHyOKqjy6j9uUj7nE9ahVM50b+U8x5QQFcnS1hrM
GCYKqWmGavjJvCQH5jKTSzbnsAdJhasMl0zo4xaMjAx+9clzy108gIHsHD6mEsI7
sunNRA+5ILCEgoGxq0s/Q7TNL2W+Vt1pNhvYoStM2/6D5kkkmpaLkPk3qz2svX+Q
sdNMqzFhPDc+ocOxHXPyjCMBzmxxiURz6eUaWBg8drKGcwYR/MyY/IN5JI+4a4Q+
qcCJTZSc4D33dvHfrWaH1TVUcrnDzZA1Jf/SlYtfA15k6zWo4P112U3oLjkk7D0V
Hc5xJkCG4TzlOoXMNiJLTxHRpM8A2pkd3h/LXAqYBu0Ac07h/ws4NTQ1bUGS4Df+
Cn2TqxHZpVuz5N+EdU5q1sdGcohm+Q2/R0iC/VnhelVf/OBHoNmT8TGcHgd5Z+ir
VplCcZ8R0wSks6+Znd+FeOy50bO7lad5xfxl2xZGKU9yeGb6pP1iEQXpdgS8lcti
jsPtiWjx0PkGVaw0+qsKZc9qs+pqwa6cH35u6D+bPZbgxPx1Hv+cKeqjcLGdWoKT
FYsmexOwzln/9c1iDk7n5dnhwgPgwUXMXVRpBG6PQaqWIVm/1bZdON/6Q7+YKXvW
BrpHGCTAoa+xrN12n2zllva+2+DA8E7cfkMHMH59EbJHbaiG0392JRpHeJm6bo3Z
JZSTx2sASf66ZrLVCBHk0/vjybLa+SM3RAXTl/yZU1tJHI1+Tl8j++dRtvs8Pbyc
D/vkt90unWcQI/KqDQi8qlMpdUgCZGUMEhz8lMKH/fS5xHLUp1G1XBY5I50iLZRZ
ANyoz95i6WAvPhGjBLoN1XDRaRTILDcA2qwsWrWNC/EYb7P09AEqK4fzKB5KJ6OB
ibJuPmnsnWs+MOMRTTvsgR7q0d19KFNmvC7Vp6CiXLDc7EyQuaOYMcx4djva6g0Q
elQHDaY0xndrwcQcAxiAHF8J8ma9C8PHNOAtDf6o7P2fixLqrmpJugXqV+AkA7zS
u5QWwfANvEIPszqRxD+0zaDIXwIEriWkQn3Y+nI/jZAMEevWL4tQRH1ZQ8l/m1If
Vy3uTWpBzfGy4hMjVBPLfVXlF8I/r6lszTQ0SJNy4jPw7t6Pg8+3ltmwrVhWqSJo
AaUmylw5YBDSgm8/rRLFePqHi4PBgqPM2moARe7QKY/siyrj3zZVPiAffnxkT7Z2
+EWzRq60KvRS3SDGzLQRZHf/LjbUq6YTNo/tZwgnkD8CnDeA/W7yPp3gOctHhqVs
9PECR0vau1AJ6OTNfxI8u4eXOmVA9zwjkruF9r3qrag=
`pragma protect end_protected
