// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KOV52eu9sW+mZ5b2C+3gPBPLAoFVSB9u5bMAKDRD/UeC6/5of20tmWV0zgI9owRF
yJkD0eNpjjTizREXTpIwTHIUYAzQgphLZcw7t9/qudHa086yDQC2F426OcCDg5Kq
T44VhXc1HLdxqJWXuCbtycxFEEm83PnaXI8zZBHWXEM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2464)
VriubktcAp97RhOx+jPs4sSyfCJGojvpDzRnszFWBTPvcAwJ279xu0wEBTsgQEf0
0cofgn8ytAaWtDs4XBfJNv3eGdeexF4OBr19M0O0cuEexdgOCh8a/F9ObNo1eNmR
+F2QANv6K+Zn9ak9GgtWp4sqRIW7RrekZ3vQ2WS7A1R3yk9InNsYM23a3VIE7+iC
YC84mjN/tS3Kkuhclb+2zqGb++y90Q0uMLOu3iJIJjVxummtHzyl6N8XKXO89sPb
geG9bwtUk4cktwR43iZ+GJ8w041TdEPyLXDzrDLqlNtTMJDTrqbDbwFXPRT1ockh
FCmCKUl9UTqmzLddDXPRebHfv6Dk4fIr79QLkui2uAUF4k3vRix5psYv0ag5Ueaj
NgNbj1yqCOdHJiu1DUxElGdsLDsDVO5zItEqyCeNU4SEzhd0lVnGDYQq6e1yV2eU
ua9N+uVucxYEj1lfZK3/pHIRq854Kem5MbS8tZh13PMi2VAekC4QKI0x3ZS84b4G
RbG2YRcYxKPCx7O8hRsy6KSH6SHkUM/GcFbufUr2zEqiOZYcFGfVEh+HfI9YGvvb
s4CuJuI768AtWucqQu0W5uknHYanJJHqA7gqvfM3QkJDL/fTC215zTrWDhfjtWWn
9+o/4cQ+262a8PetRIGmXd+lX6r8SL4KgUVWudDIw4LjAu7ryDEDcIMlIrohSh2t
iPddSRNHAeZWT8JAd6kJr+wN2u2e7pPlaogAUV29BUJRFSX3SRQKgUWqLzSM3wfz
BRYOWdyyPq2bYuTr22iVIhoUi19YE+OhvThaB8q9D4j2P4J6E4ZSIoXG9zWYCPC6
AlNyfczPXzj6i9FH/j75ZHmQMkamQJZO2LCy6Ca9ssRb4BhxW0PasckB3nb09hcr
nCwxQef4+Ghs4KE+12487o0sgmB0py4yz7rsLYoWfpt+CN0qL81zTn75cWQgufH1
CPuKKUW8Arg4DoH7xvyf0SZLax4BXgp+wvTk1aZbNDYG8S677h7GN7c/bzz3e0h3
/STWo52XjgNdBIHzpVheyWisRVXxZQCeQYe0LeG5A0YXPgWVzQTVsPaOzsPon+4R
mSiBmD982TFBKZ/PXCeP3liBTqaip8Djho6PxBE8iow9kcMCqgfjpYyCRf3H7Ezx
jBCAqk92s7cz9vCi7A6txkwwHfSna048jTBlC0XnnFeDv2TfjHEf6pdgYoy97Izs
XAtWljX53iQ6RTeAQfiHxNNmBdpinLOVBGsn0NMfkVpdA50+a/yTrl+lLPilcoXG
RD3NgKXIg3etYS0Bl5WmwTlOHtJXUn+d7x6Kp4CJbuCC0Xl0A7xX/dRFkYdvx6DY
FTK8OG3wLnS41VAid03aDfWi4Y0NeVo9GO/GrnTt6Y7hCXP821FVgZegIQBcuJu2
2OwOueiqgZ2SPcOb3PxCPngyb4orNFDRAGHuTDTPaxscqV1b5LhML/l/W6PbwPyU
5M/3hgfe6s7gsQa4D3ZOm7m+oDnZ/4pKN07+P5623eEAb4pjdbTh+gmFNT4uUSod
i0OgMlZ6oIHCYxCiMMEPmtla2jNe6Q4ni/xgB4kZrQEtIldH9xOAJL2iznTGiLWH
vPHFm6BjPUgG9mPGD6FSoEEcWobuuD235K4dmlJ2xnbOJYcfydO3zYbOUMaqxei7
Xh5GW31PTTtFQRJLAftr3TfNSJErBA+qsGfMmPClPXYKsiGCKFUz4FWg9sCExynz
PwsWbjPT7aR+OAtGllEOiAZou1Nt85nfLHerjY0JvqTKmL+e7WJr5jcb9BYp4bV1
w2c9Q1K+Uy/5yNrog/YU08MPvuo2s1LqFSw9ZlOh9FUVsA5Mgn0rPp/jMNVw+IVh
ek0a1e5SAyk5ufDwn/iFTV/OUK7Br2HqX8oTdxECrDxQ8EhKaSP/v0ixZyIWoLHb
eGEWhuYDYTIM6x4+uzSxaWlseFLygvmlfK1NYxGcX6y9VAxW02yvnu/u60+31Fr2
fM8e/KiHVyKOaiFQuaS7KXBPc/+/kWkmjigVo1IFwkTbWUOhLhdBqPKW4PSJbPS7
7a4iCKTPo9L3QAi3vPmymYxJcD9WVnFSP+EqwCIual6nAOsuZhsyDeR57ArTNsNa
VOGQVyyvhc3USCmg2GQkslbH3p/rbbnwSv4MCfUjpwBksMF39c1NeCPPI1cYNF3Y
0JZvu2TlReKwhOjYounDdQtKfw5wR5fF+rEx8/CYfxSozbALHSGseqQfw3zi6k6W
vIeX4eciOWm2Iq0JxDxqOajnBGhWdQg3zrA9pTAD8sx8vAQt2/WYRame1tUvr1A0
NKLp8FMSri2+pyrzgzXh+SytW3JKsphKgJo8I2GOk+rCw+uYDZz5ksBJporousyB
gVcd1EPnHU8FAMRy48Ck2G+4C+GRLuupPjtcL6o+8aGI+t8a+0pNaRxawyjKhham
nsfgPheQYgw5d4fJIwMNxpAKD0USf40J/O68NmF72KWhQbnqc02aeaoQAKHiwls/
Ovx8jq6f2/Rped8FD7hNKJ2UhMR/aJWWrlA/BRRjFEdn/PKLvPPljoR/LYjbuBU6
tCM1P4AIMvmpFlRZCVa5c6v0OFDNb+79YCslW4SHdXOzdWbSMzPWzCy41NVnwx1e
8KSiDc76paWMJuqnmMvX/e1v0MJOiTmFTV2CPok89QzmPuScfGZyQtBHTwMeruuU
edli9rKqwX9EGr9Cz1HjtqEcYftzKd+riuo4SaA9rQNhPcpmnOpAimuOnr6e6LcC
gRAq6GkpKY7dMmC4TK1uupeIzXbKDC43U3AprRYR85xdIDfqPCQ32U4cDtA3H/CS
yujdUjKfKXHMzCxRWEoQqp4Fj4hSJqrypaa5TQsGnDgY7SJb2ah86JlMXC9XX8cU
dy2jSgJAGCjIr+4owWYe+8DYeQuxK3da+m5voGDumDLQuPons7pk4XfC0QS+nyzI
7lTXIIlLlPY9TVz0scOtV5pOKdenBrPKJUI7982/+mOaQNmPIQLbrbz4SUFAZl9/
ZDnAjSxi+uq5lKJRcKyATYpe/eB2GNjlUfM+8Iq0Y9+RAObvcdyYKcEhmGShpCW2
mrafu4fGx4TZ/AtPBNUBxJxR9fJ2Df9ZDgL0rvWP+US8yFDp7RwAg1XaXrAYjfyy
xyNQfi83HV2Q/003A4WXp0euC2PB3jHihDpY5k1u7pU6vH+2ngeDrp8u82ntAdDY
zUnysZuwnbZbfOPnBAwM9NEeTOnbPQMcAtSKNGfPYwwFqmA7OUlxpj2oKpl79MJJ
oWN0/R54F8VpOo9RnowMzQ==
`pragma protect end_protected
