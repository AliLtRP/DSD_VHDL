// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:47 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
jRQ+4YPO+KAQ3UetvcKGCrFNtEHiUH/gbCfDe/mQ74NzKMHOPADDaLKkeZOPBs3f
jvMNd2x+1bbqA56v4DyiqDc9JJE/MYfGJSSa9C4VP1SIFjcr4jTppeco126AclUF
b0s3BMPktHSpwzHeYinjTgfXwueOgfzQOZi4SUMI0LM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3136)
qBZK1gAfjmTkpYw7Rr2rb6gvaoyki81GcQod5m4mH4oFMvhd8pyq6uXc6wH4bnIN
hdMpkPnGh5ZCos0yW9G/hjSrT8xAjej8t4OS8mMAE/+vBPzI9NH+KHPvouJw1qYP
vbqaJn8q/Pyi7Te5DR2pqWj6gjzzSt1TT3gJwg4HY33Ebs9bu8pnA7sxz9jb6/uY
kANxb6Kr8wrECsOQVu3goOYhOU2PE9TkRoYWBaU56DJPn7mlPCEZYq5AoR4DvqT+
7KEazppD8blR58vvUyA9tzN0X1ucBbnIcgqgi+ykyVFahxPRplZFfxIyfgCTnCTR
6TQCAj32CSxmtLG8QPZteGVTVnntanykHAcRCS/3B5W1RCk4a5vqGKLz6FYQFeTL
opGZw6+0Z+x5H7ML6O0+QXxkcOWcHD54pGX6kmZ8YgQpLViHoEyUPBtaxDM61ahv
Rs1Y7Xx3PGsQYM0LTD/5musGsnsL7PiGLOIvhepDn9aPPu3k8NjjwexDkOL0FSmy
qofd2XRpm8k7C0et157C5965kOMGWeyXSofgO96bvIEZL4YnRDEassEsSM6mq8S3
vAYr1tfhEOosFvn+GSAla4dY1wicdk28mCzSqi+N5lbzqHogAueCXwlhhw435bfA
+ixsupJHA9ZUPpU5RVr5Z7RRqKIhyfzwKuHRqMQquDsKQriMe8ggVkd/HtotGDmM
lY5u+yoaNU8k9JEBEUo/ZMY2MiJBWy0hLf4p2oXq06bfC+zkyVc8aFNeLwDo84Vp
vH0cGB9Vh4GDoNtgMnEQeeQjTfccyIuovE5iS4ZX62DyDOPkv9EIcYHm5lvKX+Sq
v605xlyI/URuL5CSsnxs4uJFgT5FTd2AMFwedaIE+n8JUwTteWrj7hfnFXDEihhG
Y4jV4oNMrhjMKf8BQNINT+7VUC9AZK7IoyR0v5v/xutW4sQH47BGQq58JMaO74hW
YJyKQu7wyLoP/RtPWhp9w4WiRO/eF8g+AjYbxWegtbFpxAU/tAXxKROyAFI7ewVB
AbNgch0O+hayBZsQJMxr+4b2SW30h1g/kSE7uVlZgMTKLx89dx2k++a4ZU0fpD1U
xd2zeizgA55T72hMWU7dMZxfhgWnLoQ3yFJUTMFtCC5tKeV2K7qlboZQgJ6CNmKu
i/V9h6nshgcL2F3ydjizNl+y0sAHzsfWuC48RhGocihFRkbP4X4M8oEM0pjlCEmC
9McMMQFoDcCUZPzFzA8BdHdRcAXU6dnu1sdt1N8k+T+ZBvPePrYt65EcMVE8AkSn
4Ae+Qd/0+JgFTUKoiXdutuZzhhTqERw5N/8+3p5jKpUpdxM1S5y5NIpoCK0CKo52
JNhqPsbpnHGBz+sDR1GteKPBfLRIHjuRoj8Tt/icKigtc2/2+drntJenezhcAVlq
+0uxYc4lV6VIMPOx5mmLhyjL8RUaAP+R2uC4A0FixH8F4TndnYZOaG/aFwSbNVCz
fhYbNEoDpoBHCs8rJADjjgzKYwvK78jvP6vT8S7pJTQRpEnDtYw+w9YylTQ/lMYC
xQXqpy3cdEVVd1gXRfe2I2IN+WopY8PROp1Il0RMTgkNRXh/rvEQ3iZYDLpgP8x1
eOEP6eIEn3ZlghTmn/D76HaAH0IPgBt1Ksms7Cm9z+17o3BEgDaQ520l++dHFvu4
+ZLjWPL1i0YiiQcusLjRymYzfqeBpqA8ui7waKo2zcdD/3r6aY+e1tJM52I3b99I
/OjSEZ/kNq6kTND1SETn109KRsD6D2vWmbAUd0oquQn4mlHu1Bq+J+HXVg8fyXIn
qDwmUVs23rp/BXIZ7NMnDTUl6wtT0Ql7s1yTCXrlOYn2j/PhcRLAJdwKpmQ7xjOg
CNvrSI+hqAVmiZjWrdiVt1DQ/t/64BthVhqxkjYtMqnj2+uD/kjr9Yz5jutsHwyy
BdNnXXVn7o5zH/dmBe537PAFUJTSsEDMH2yvPMG8OcEi+13A9xSYv0LDQ14voBMy
ufyqiqWaEdlkMO+vspbfS1+5UBDefFnpQW3CwATot5QSkdd4dORttiebyQGom8Pb
/ySefgkfULwQaDbqYMlUuH+/LtRgPkzXEXwR5jmDSQD2zfNkw3WEbf3B6avpxZiR
2NfywYcyejVxpy87qM3a5T9lM8XUdmD1c0pI9efUMljftyOX7a55VDS7LHZkFuL8
4P8U6zL3re/AF1JN/JqOmSYXpGu6FugTgIBuNaJyfVZd5I+tPmPB7Mbeb4DQThx9
ouaqxPFtc4+fLC/z+Oj0cxqEs2amrcfwo7p+DU5Lv+wOcAqUwxqbrN1RpdWu9hAL
bGZe4PPXPQjGxr1XE3o+UZdbd7JbNjX49zOhjXJZZYUcPZrNHxVeHDzWBpe40UxS
tpyZAYPrHMV7yCHca5chsW/kmM+j4R0e5/xSlxuAeupas1MP3nFuN0GgWOLAOk+i
ld8eCC71Xbnful3PcIKJQB1sGfM72rPy2atetAE564nSKoj0r1Dib+80MWE2mzjc
rY4xJIgAsGrQ0dNqJazOrH6zN3diWMWRj7p7CTuydkgSWFUfLaIx/iW+hMJmd5ie
8/HeCaLlVU6kXmlYVKAigfAZd4VIiur9ahrbgRms0Lnr8ZiuzYRGydK10E+fKeyI
nuHEtY6r5oi9/V2/78ePEZFVCcJOktDt00O0G9anUrodNmdq4Ug5OYXMKSsdUT0/
bT1KVoAM8F89j5EdfPx0rGYhfoj0/QqolM2dOag+8YwvnP4xlIU8jrUcFnqFSgqI
GfE6sCkqzT2WWOsNJDKD/jDwD80/3MWAgSyGfDiMmyyd9T5iMzov/aa/Au/W51+B
ECewd88IxERXv1MpsnIdjj28H7N0JDRQGXvKIzvjdxyF6QzbIt193tamjNlQ8FUR
OM0su0QkovgL0GVjoWZaLW2H9wqhC2wWL8xwu6EkqJ+tl8DjsjFm44+SumcJ/1rQ
ZBqoTxIz0vNkHjReZoq12uiMAALF/DOXUmPudIqGYagivOfCx4K5/YBRfQljjyYo
Ko5rvakp65NXYVlauJ/yyLa3yIGyiXCRJBTAJKS9r+iYME/L86AUwp4xJWr7RgaL
7mPGi85sRntJobcbWdAsXAPqAGzVzNqvdiQ7IFvwnDL6maQ50mqHpGzardQjjuhO
BNsItgDedFuh/YGDVOR4b2QZJytrA9Klb/xAu3mIMmUbZr7PZGseWrUuqheFsccK
tkepBiHaAHlRY394e8T/56aldlZ3p+Pl2yp7j2YWdzLxAuEGTEe43aYqS90xXsWQ
/QqDPdsi7w3TDsetkwQhYfbu6JqojHpWY5X4KcGwGZI//w/F3U2huAw2EOn4iM+m
4iWZfwZ/nKeYlENINJQzSocQh1CqUbN+FiNHDmiVDj8Q0h8vSXgW2jsUeVrz+t4e
JAL4DwB6KBzMTH1kGaqBHcEsLPDVgoUxYtiXndd/VX4y+15L1T+KAfaExp/fePLz
DeaaV/eAUkHJ8LpYbmxZGyrVCo6t9LdQg4gatiQJWr8mCTmUGzcKGah4HgIOa8um
DtxFeb9fL2tuCor8J3l2xNat9DRg5FWRMuaMHlyhYZOOTFVY6JQWiuRA9i7ZUBCF
Gc2hMZBEiyODyItj4CoLeXnwoCs1fxwuZohV7pjNDicOXIwhMYwOygAeW4TnpDOO
6udx7AaxnFdjotYhGIM7K/XtGyzc4yn/bPLXOJvndpPdpquiaeRJqLKZA4mMRO9W
d2Aojd4zLoiIYdA5l5wTniCqsM/6Q1stFGgL+8mtb3a5mVFqL/GPkEAKbvoiLYJ0
TTSUZue3i133QlCWBCrA4E+5RKrdyP2c/20IRTKB8SMqnlfbZ3VvxbFQMrrpLYFH
9LzIFwubSBIVt4e+eUi0fGGE2VvgCthavJjD5gQmQreikOWp3TYKUmQ2/4n/c2d8
n5i4U+T5ca0bCjXv6vtcFzusiYgcOFn+GLJ2hP26qsgGNsEOfqqAQqfOgw6Evw89
bGGpLaUX86qkXzL3q2ElhKghr/ZqCUOgI4QKlXpRPMupJSGsV38ttljVHdF7dEcl
fc1xRJmE5npTG82w9O/oWF++wAApcX15lxV1IHHDf2STZCf6GifrcwdD+QDUQiAd
ILPassHv4g8Tav25RoNwz+qX9FxDvcizzngrEjn+ZSfu0b/4L8aMe1kS2eTtPYoO
h2x0EGf/wKYSirsNCaArIQ==
`pragma protect end_protected
