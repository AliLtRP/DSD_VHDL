// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qVY0Sum8YBuluA4wlEYO0OGH76NKUYuROucqKnj2f9eVUkdnWmxtHhzg5VBZUsVA
lQjgZZvcrvIkhmLlnvg/DwUeFFBKzM/tK9PFa1/CFyiP7oOsMlnWtp0YwLhXJe78
ge6gEMBNFarmrnwo93QLtuFt/lCEGr6TCpd2z1WQ9kw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19472)
vCW8GsG+Ko9+GI97Jky82n4xO7ZHacw1ndj8GtAvUWSVZ0Lrd3du6EwwNCF3LEMm
i+uOtg1WL8N8SjAy2IVn7+UtIUg/s/V3SUsbyWP2MUXM0WdvPhi76lViwjs+9YMn
Vsbu8gHNThfQt0rjSuwMGh35oA4YtRiGdepLrZS1E7Vm0M2ALKEhadFWa/hK4O2p
oKTFZGYBmBiT/GzQl5Og/lGXFL743BpWwegl3nkcKHTFenpUPjvmffibyJ/rPTvG
OJiweRE0EZ2NqCPVbzRZ1J7vG4Sb5wfCgBXcarS7YlLOPwS3qvFMoYTMrxgCG6wM
wkoknhiBAc/xbjUuBOozOjMxTSJ/coeLnYt/kbSj8+D10dJgVasQOsTG8jpqYiGd
mDSWc181HCdV5Ty3oQH05mGsOzcLLvg6TaxV2lgoeDxEa7ok8ERptlj5vpJgxu6I
N1wHhgyzQI3jWXV0pQCxFNe4vbcwd8ebcUERYLFXflWQeJ5Q3PditmvvLLsylMuP
T7sPHtN5arVtFpdZRViCKL8nLX7DYScg9c37GG7UIg4hZk8InbfUaoPBAGkoKED8
rRR0/MxO2R+DUfE9oJ78/tHZRlEgvkX2Fqcf1C9o/4ewod2M+77+8yPnAPzLSfR0
48Df5T06VatYBpvrLahqFfZp5iIrFcloaoM1C4ZXZIfGsKjSfVUkd25ChkHI0mC7
b1PWeMWtOWOANO/QmJ9LFNqzIebeFcfiyzkvqlQcZGGcvyIOFU1ZKJQtmxywiCy7
JzZMEvGPfue6Q2dtBwwMbY3qKNbTxX4HvpjfmuhYfitPGYuidSZo3aGVZu24uefI
wta+cD7CgVilEAgXTl189J0hW5ru5SiZ6o9/KiNiaO9A4/eJce+jJzC9M4WM1Fmp
bp627JFj5OuqjjhjnelaPKXoTt0i1pqmpLVSW5WuT81mLw1L+Ynv0YDKU8JVIcLo
N3vBI8a+JKk5SB5fBUDeNK3aNbfe7SxaVDokVyggOa2xsiILlhaH+S7OKxu1770l
qulCNhJQzdv78PbU4koJjvkKOemKe2CDsVEg8pRvT78OSfE3zMAmvIrgIFmuCFKQ
FMj2qq5FuoMulQ5g7YY5i13L3O3Y/f9yNQEkImv/weEmDtUpxuwQrP1RDUdjSElc
rhNeYGfBRJ2vGqC1RVBxQhj94jF9rl4pP0fUJFmK7KmW0Y9BWgt8KN+eblRxAxOS
3hon6EtJxrGlC5icboeXJPihmqCBovc8PO0QZuMqElZpheBsSkvM59ufVMJSb4P/
MwKKjOjfgtN0qVg2par7RsxuwXCv3uZE9eahkgFxTz9uOFJVuqAwjKCcLSYH/u2T
QZC7bY8e5mdrT2WE3eGt/vBMjE7Sg1oVzJe1MEdx0BcI+du37SVshuF+f8Isw9z7
yRpGJDHUdgn1QBWeHMfaMYOpz/lZm0KR1r29vM26WSfZggXKS7Wb2U7yz1MUCqKc
V+8RBRDFR2uWNxgXrh5hi5eHDUbGyXh7HqKJZKrybtMTKJqVJhFJylHgxDbzWeuH
QjfKkSqAAS2Ez1Fhw9bUUQ0mlWarRCsYRXg+Vo14an94ZoPcPKhHjr+kjD+J+t/j
wdF/0Y7riDHvCNVFsO8D984PT+Gkrr4P8tcoTMX4oyVh12yMCWy/ooru3WIkkwU+
68QU8HaT6ZBCuL5CbIOpxXyzgKwVz4dJZ0aEzLERDrWinVPbvy0JdW0IXNJ60dMr
nAvWMDUz1L/pBw1iYx5L5mrbPY0xuPJChkSrbcPGX3KL2vgEKKiPVM2zSIMauB4W
8DdIST/zFZ8TFbq7cuyS24t/bwSdFJ+qfW/WXiB+DouI2eiRmpdxH+RnTpAEprKD
kif7sAkmLyJg5pzVri4GfSEocZLUCjz7Jf9IHkTrtp5HNaVMX9/Whv4IIQDHRBjW
dhbvwXMZUdm7uyZuQcpzQNJT2sjTCpCAkweLoTevKRgU/Yw38WFgu/pjfi4c+fnO
Xw9qgo4NN1QRKWTFMXOGHiYMkYkaR3Xp06g1anNAoAw0cZx/hXNC+Yg4odjefmOU
mad1V9k8YhdVcBOppEELX49YYnHXC2r6jSYkeIXEGkG/JH8R968pZyEIN6zbhpCc
9k388q9DYo7FlVVzvlPzq9Icp+pEPdW3ZAtMrryaRuZsNonNGSv9J+YqPg7UQhgM
q0GAnOw3uHI3tXl7bWvkTiYAzcE0t3V0JbAWsffU53Vc9fdx+EuAP/pfSMS/O/nr
60dZmR3X6mdwzob7NbgJHPI7QSqjQUN1yE95UlFFlSKEHpguj7cHGZOPdylj56mC
azman4mTBXWSoQVnZWX1ho5igEXZ33EYuB7KKESMGDwPK/MNd24pRU8HaiUJiYym
h1t0DztCLbuLE9sfkN1JgROoKxVOKHOj3yej+BNaNXB8PgKr+CTwj0DA2JnKQY83
RYm0ugR0+PXt2RUjFQkLbRexfBtqgsDe3j0lVlu+LGFFzKNwipuInC0sQTvsZz9x
ZBzQpnSq3W4/KOXoiJNA7u3UdKiPcA7ibS70F+Uewk0xKHHlorTXi8O8oavHsSML
h+PMc1RiQy1ugnfZTU0RRXi8gksYG3bQtEf9iCRF+nIijiAp/MbQ1MyU2xwdTatB
7C+UyxHD47qUBp9wNe7yWM8u2IjXynECBoMYQm29wm+o+8Qp6CT8usF9OtAJXlZB
Y3zvEmnPip8Zyfm+sNuiA3YIGmhL/Ixfh0Wk49mWigm1hMs+ED3zUWrUC7OTa/rc
1OtorG0wsmpj15scrxpxss2DuakhUWJn4tX5n8dmBdqaRFKLwM9OOe2S1ZqMejoq
4h4VU8lU0WgW4wralLRNhDfPvyZb+4iFBhQ8wQSz+Geg7NfkXsicBl/ytmAIzWOZ
NvvLv6WiwZp0LQbXizurZjvoduH7qDYrYlmStWtK2qeaxKhlxsBwQQRAeSYJC5+c
KkCjGLm+Hr0nuo8qlspmZ6QbxJ93PQQvN70xLj/KiPC1IhXCazRuSZ58CvSFbLWu
d//t/hS5IovAMFTs7O+qsl43XwgxhXx0RWKKJ/VBRFQ5sPcU7zD30HjPtzs3fQS5
XaoDoSMPWBFsoeaPi0or7ZSlC3zTXIEFeklkb6R0MWNtLOHt16MKidkp5FrlmpKk
te/aj85t9qe/ZeBKMFXy6FQvjuCmbBJqkr+2Sjq2dxorZ9PfaCPdl8lmtPAfaGFN
dm4IkAr/ZNJKRrC9LxWdCaL5KTeporqKbqfHyiUnVSdNi3Tac09GMgm4bFh1pgoX
6eOOEgl9D3xKat+3uhPDHtLjV0r+TOOnTRBY9gCjm+n1vk2vxwd0kLbBZMnCKWaG
fSslaEUendqLklvcQ2CJCn9MZXFiw35lpEpn/Fq8mTgsiJTZ125mkdPfgRGETNYC
4LripiIUS7TM2mVorCHl/OV4e6a0WlzkjgliM+h8JAvChT/ePd2yUWKm3ysRihyJ
l3QKZq4ICgh9BsgfYIjRqPMxQiHt9euw2Z6Eaa3RX1iII2uavDSX8C8DjEmSZqI/
sXdKiNjmq1SLnpYHNmpb1xotAoPoLg89rrbFyhth8JHWxjF+6bXTxYl8jlYUj9Yy
BdmMRKH3Ab9U2k3nEYlpEDNi3Yd7Y1Z2yTJJU0xQ0m6MBv3oq0v5jfO33axLR3DR
Iu4dXxiwZXzHjc7rps+ILpXgR+arIEHWA6xL/dgp09bosRxs86R3Kk4VqOj14k8D
VUGK3/hSYI1T1eDJEd2gn1yTk+Pr1YWe2nM+aTaDjagPzvdsEL8t8TZFDsIRpSGM
PQCCPgyIE6yZhuNfTfrIHe4KGWks8ULYq0/b5IzAw2YTDV2dIvWftZJkFTXe8oVq
ZAj1yD/VbcgwjKRajX5A6+D+mgh+Z3gMNdi1Q/TcVf9ZnWDsw+ViAfaom8UJTdcA
V+PeP/Llh05N5Bd+b3rB2uD62vFWwsk2lfn5pfRpdyranq8sozY37LNqVErtyQVb
PuVF09Qyi9Q7yvlTdWyW4kYg6PZz4y2/00cqoXb1nzrt6SGNpd4rOQKJq7pKAV55
duq+tnoeifw2nZb/Ki7Sal/2RP4gbKLchjqobqXjbBc1mdC7xCjAVhvNDl6rLQ5c
hetSeQKRM4tZUokFZAdI1FOkGfNyZvP1ILkE71BpEES97Xf4qGogY8lU6f7qHPc0
q4S23Lb3EOtJ4RUifxVQuzVPq86ew9SvsSscYDBT/qCuPNg+cveNbe2edKuecedu
Z5ahGQqszfdycKiqIOiuwjsPONqyalHUWDZuSAjLLkehMzqWn9Vo0KRGm8qalZ3Y
wNaLKa+5XpOdSVM9gttnHp8pRXVLYFU3lM67cNfqG+tCdSK7w/8tCRy+JJOTBO2X
owpcVVOsx3J8xoL9uru238qIb2rCnRQMYFfk+yl0i4uYYBMDzeAHeRnsWPXIS7ZK
8EE3vSQRG6NCtWY/EWxvd7As3/Eqqi69fECxpmWQoOebBIOieGOFRw/NKwRkWukF
oT7hcylBZLsvuH0qQjAHjQo96awYQ13jeZWqwSbTRwsdHTTjjCxq4mLnXvWDFt92
n7Bl8mUyPKxlvuqZ+Yx7tixIHcc9jPihjuOxV9gPiGcvcu6HF137j5Gg62uadCkF
aUeF8jJJkXSi1W7bHdttdG6BtnO5fkhclE4Sq/Y0Cd86sOEbKuTzbS4XlVunb3fR
rLeI0dJriqC5XHbtZnl3aF6o6qgtpJz6/9jYVWFfDz1ZUeRISMyt7XRb4QxYwYYv
aVtKB+t0x0kmKfmEstbPZquItllPPYBoNFs9J423vJBlr48tPykVhbjrdrMe2WbM
6L4iOGXgeEKa+nVzDGF1fFqibxdGlSht09cMluyo7nhN67/oyqx6Egplc9YriA+s
0lg6WIkC/lQ7eirSK64H8LWCxiPp3HlejCWwTIT4aD4gZ/giQnV2GFIpbMXPbqlN
ZKWLcXqWgPnZCi5P0UX2lUVpaFSZ7JLzae7TdwLpQ2+8JxiRCEBXAl20m8kc4vtk
4fRCMEhu3RBsrC5HNeJSzx6mzIRRMfc5XtW8yvDyDmg+HY5MYpzGZIkThIEMVPHB
TxXWA5PC2p4gdNnwcMa+79st2vycJJaDV+7XILrNJMkNMwCAGPWSkH1dEqZf+R7X
t9SdQJj4bVtFk2gnbIcTLwxy7m3nndNssv6rK/aRAdWs/j8pM+IoOc0QGM7QCCGZ
o564y/FpUbgtshSqIbY7LzX9cqu/8IXBwvN9Br6aJip6Za79sWyC2nAmwlt+2a51
Qa+JkZVGWvKOPftQ2Is4GfcdGUSrEgGt0fAtqB36Q/zjKkZUUkwWhXvnB1ll/LtF
JJ0gMAp2/HgGpQrmColZiZWA8fTTJNz1ADU1l/7/p/19tB8GIoItn2RxSzmuv1fp
bjyUy4Gw8R0ECuliFdwxuhVNMKH+j/yRGccSblaNtK/sHUuxwCoqnu8o4vkuldl8
eF/L1RJjXIFyQv4F/zMH8Rnm/WnesHu+/yEQoqf6E0u8h9C0aVCkF0msvZ0H9fvV
Pdwk46siBSbkAnIRfZl6zyMjIMfQJnzK8BXTp9AOEeKJcu9XCJZ+D3vQkPRcVG0N
Lua0HwtVcHDfhkmnuf4lfWMOVT+hdwhRR5SgQIWaKNctHS0u1TDMGtCjDePj8km7
LSzq5PSkToxFtHb/mRQYBtJWhE4FTd2ORBH3HtFaQJMZHhhIcnvsZa9cOk+kFZIb
4GxZZNIjT9Fou7/41ktfssyWuDCKyP+wxDI1lltITnsf4kUbNqUyB3lL7Vn4SPfV
lj7XhHkAcJZbjeF2yth9QF8zhtjZygjS7hzzmLcmdPBSbfZi5nnUcnelPTIYR4+P
xVMo1nH3i1si+abZFELDeZFVIP2oRGYaI4yE1We16SoKsDyMhw5vy967wEKMMQbz
7S7AwF2UjTMZd/5f1zyT9y8tzRpFmJO9L2PT/pyJ0UsIQBBXWaPEINxfzSgrLxSf
mY+WlmRNm5zNDsN7+/PPnzB+p0BkpwItJ6Td+ByrEXPTylMhi366LMCdXXvHFueP
QQG2vyybLeUR/RN1TIK6ii2TVPObnujJn0PZXY75SPVuutKWUJ6bWvFMXq/jg96U
1Do953sBNtdoFoSktOqlA5X3wI2yjJYIFbE79CS3qO/ngr0oWaOE/Q9bsL8vTwUk
gJYXHf6l+lvBp6h3MyX/5nd1a54EV+AkR0NTL1CgkKGWaPAv+x5qwVo7O/LWAjjF
pnyeE/m2WBHgr+UijcR/J0k7fGS+ZbmTpSzMQm+LC/xYfw8NC6khyUz2PBHjRTpJ
FV+tcW0PR5WSP5sZB/Ix2MkB7b/OqrEFNxu95dFvi4+ubwBwIUKEUv2xEdh4g19h
GHVQebJACrpdT24EDvAOfVdOVNNNa7xjyC1RxAAYuzQLuQXSsNprw9AKAI2Lg2KX
ruuzo5yveY75exnOUCIf7O9j9zmfjNOUo5YFK3yvZBWLhsgaonosTLrrfphZ1qqL
ZImndYgXCVuSxCaIIp+qLLSHi4+hjPGI4sBB+V6sgUobJNaJFg68Cp4Q61BX8mHt
GLdbG3n1DVkOII4qjBuTWmAcNDh2u4UkU5hrE6gckNVCbsumIxbNtyQhUaTIqPpp
Ww+m46zyf6I793wbpJy0ADPwYZ36VgAvQR0Mjosj8jQv0W/9/x5NOmPqyucoX29H
jC9D3eT60I83T+8TEjCyAqLfC/V2mFJIkGmCajVuSfZw7y3GaBHeAx90lKn2uZpp
nTP4fIP8ZzL3bXDBRytxm3YHr02lkNExy7m6bLDHAm8Lot13MasI8z9eUNcWM1KZ
vf2tMIR1c3R5k5/qqdSihDQOhMhmQBEB9DFzwWUA67pGfheho+LqA5Nq3E0MFTpm
a+Pz+y3xVsr8jXZnQqgWzzw8YVhxCIKBvIXxpTtBLLO/oH4YGgEhLkD70VI0bdNt
hbJDbqes9rY5P6efWnuJip6pRHc0zJ/bMGrWGp3ZW3M+o0ULvwMuRgK2KSHGPuap
bOuuj0TBd0xggsjw5XE15MXCIBIL4xszKg6W2Hvgt2dmU5A7C3heq6a3ME2L6zbS
E0IC2mp6E3p0uW1FDbfs8x/IS4t4COFsWpS2CEuXErphV47N3KLpd9ntBTbwlQQu
0C7wNxATdusmTgQQQ89XhMXuWrU/eLET4tNzRp3oCH/A5WWhHhg6T87BVnjUh6yF
D1bBeDnuUTGorZ8NAjeGfudwiZbXUhjJol9UIrfUHD942wUiFpNd+0LLFjDT8KXh
Wc7S8rTBrjD9aH8NeXURieT6ahIIQeFrvZBGTJccWV35r29pk+vcic/8so2wtCBR
Dq5NHxFDTevQxkEcxhlC4l1J0R2A0Ptbo6/6GWhv+yXdNY8FCexGBjT0+iU/dW4a
MeBA8/Pm7dDsR2339Oc0jXfOdIiZ3oumK1/GcZ8UfG4x6VuY/bEkWLwOCQS7tyom
jZ0GRrjYzMl/hxt4vkBP/tNI/WXUmsC5F3kVIQMKb4cWpKLrAg4Iq5lY73Km+iNh
X3fdPDCdbBEE0LBtdYo6TvqNrciHQjgAmtx3AxV6zSmLjrOCbpTD4jXIWL9kVIm0
g0R5ubmFlpqgv0W5tdFW/Rsx/6DXPgn2Rve+fOEL41zgnkRp4/wI4ZDuVdtejUbX
rTqgpSJpChDC6zGDXQ6X+A5wdTV5FuqThkkNfKPZNrqBuLFcVkwBBiLysEPwNbVn
/HUcIzbs7sAroel92wqZ9D05QMUcjKO415eiK8pMd5wu4Dimimep9ZuBPFVhHYal
w7VVPjLVj3hR8+LqZqiZEvCGto4Q1iX9ikNcsfavIJnloba3NapSMd5Uas/0CGd3
RZzWcppjDSC8JuhqEo8ERhyE8D8DtYjYzwonNExlbMNAGeXSO/nzr4YpfnB2IGfX
Hbv1a719U5IOzEJQjyn/lJj5QYXB4T8cpgWTvzG8PtZmEweBtYC14yNLeOzGjqks
qAyzTqzYWuzRuNlNP5ZDq80nDPadBdxPv3PamY593ExwoMOlBOooh/pEJR8SFCSR
2Pxu6JH8M9d4RyNEsuaAbd+fC7rjlrK6HWr9GqeatGcBHlJAZ6QyX3+p7GsGafvW
nTVe2+4ulqMC0g7+uFp/hI3AZimh1JsPs9xA2VihETjfows1c9iImJwcqMWCemTx
AherCmOqcphyuvN6RMt/eZbkSe6g+w7OYr6rI8/JDl5c4vCJHV6LNrJMKU0yyfSS
8XFFUkBWfZOcpeuzpI0meXUrJI1d+wS7TK8V0CW64BGyQqbtofZgrqbO8uvo4yi5
dNk4OvxEjXqwmv7xXzVVLW58j9x70U5OXefzGRdlE+UFu+4Pcza4JV4Ygz91kYn9
rVHz4zmJRGRCcHo3eKeN/V1erh2YPrVtXUFHCBSsnuXWkCXD8b5EZBeq+gyUPNb5
XfwpfgFm6WkF+66IN7UKqcxs1apWttWVkipMaffrJEf+tf6eINXKjHgDonxBQfbf
+FXDOXeNTKHqIetlobfUIwFvahUwHl21Bcqkyu2BIyBPrzxbcFQ2e06u3lROIkdH
gszhxSpF8Lchbkfe6rgvsbZMqQ9Y6xqkd3cf8tq25+BqRrKzgPGGMrPhpO50dqPs
C+bzcubpRgGQreKkKZY8kAyqS97/EACeKppUdGciMH2nWE5e/nev2Nn+BPpwIulZ
uumOK0xbcjRSnKcxXsueF97kJJNnzh7JY2jnhjob1ZXtD3ln+oL+LcHXbtexkhKM
yt/JQm06jxyseJcAO6JSrO7MvjehhYcnHB9g7zFM2qsCfMw4MMwxnNxwso16DXPD
w+GQLUXMd9YMLXN5la9STM8YJN8RoB2Xz+K0oQBynIeSa9uyt05twj8WdoWHdKju
QpQA6jRIab6wkBv/q0p+i4+EgAqfEezNLzZMoUHNKad8VnF5TI249/781sagr3yE
ec0JQic3TnAxH4AAPz/D58EZ0GghVBFV/hbytQle0T+oyfU0xjLedihqR+fLru6s
/LAzkSTrab4bAgl/uq1kRIplGBkHrkagerhqKcYhsTgdx6CCTglMUqcd85sQRmvk
3Px1t0UVz8z4R9+ea1Wia+updmvL6FVEXa60Wz4DD8w35aackdcwQot45BfU4s22
ldk1Ha8vj1p72oVe+52OqS9iL/Sk8a0t/AjrjxYeQn2/twhRWxZPfJD2axRXKU8o
/NpA3zRBzfAzxDSQRBTADF2kVlbkDk7dAiiM0oVzdv6877JjQHErMp49v4drK4Ah
PZj0X0lyFpLwISXzJoALouAU5cPIVukfxG3b56TStKHMDITQ6qWrODBQReicBxQi
eazAcqU1RY9I/EMNst/AsxPqfEuKdUQ4SwnpyMoEe1kC2Czxnrf3yMm/4mtIZy9D
2HbNANbBMzeivdpcYGEbsgm6FtJwuJTIUzXkDgCtsqjjqNQ2wE2xL4B7tFV0CY0Q
D+oMadmBW5RWkOdgi0qekbxJ0x2Nxe2pJXWzulZiFh905bouVlKU9rf2aA9724Oc
vOgHRRdg+9DJKnCLCN/aROKZT7e4tAQzwdL1DM1X0pavIgckJJaSCXjPv8Z4RqG9
OcUaAzIfg0zSSuRZ++tJ1wkcmvyEydygQD9z1kfdA/LhdrubDFcIOAEx1i6c09fO
LBZu9RJKYJ7mjYVJzaOSQ02rlv1nLuLNNXqs2hok5hgSm0T4memuY35HlJC9vo7p
BqhbcJFkunZOa5G6J9XJ5zScdMT9/kkefuBxADO5KfCCCNQzq+yxVFvSGdK/WBmg
Aql2dqflhNAZ1NZNuxx5+SsGpb0rHxBLapPffqWDvjRzuqH9zSPzMB/a4GjDWYbt
4aUUwSsJ9OtRcOiXX9VfeqV2Pt1ziLvKHXK4R7ag5ag68F0QkUTg/DeWK64f9yPi
cSO+RQwPGbxyOMT7PbIeOCv+mDoCFUUylDTEIQmhbDoBKW8HXLOiIl+N+Iyhs6xe
EV/qQzJSZfvXACvNzaD/w9NkORE90LR+16D9nXC4U0ZQ2B2vdhuoyxeE9xCwBQ4q
JMMVqkw2XjoKFYPe+JmDZLrv0E9fb6fNqW7+QpW7Q/fBTDDN0R2fP8OraOHE1t8M
64WifQAhyzZtxYNEnReqROoJZhkBKJqhztW2RrIf1fiK3DkYZES1G6yU2+GpzspU
+r9+MfgZ88BadesPuyzDawCv4b7hSOIQCcFM2sbzDKlPY0Fj0K4yLdSoHS6yqU/7
dZY76oaZg237kHpJoZr6ISZI4KJujkkyChUDaowkO/FouiWGIE+DvBPhqYbvVh/0
QPzAS/yTj85Kj4FCOi2Jt47Bvh+2/NlTOAKWe89KZtA3J5QzjxF6yV94/NW1Q/zL
SJki5GVQEMgW2gQCXZCO5FqJ4iGdWVKb1i2KhpMwS2CLlJdbiindVia2hZ6F98aw
Jc0JvViI4ENKKzegrVBnJjFuGLzN+GbRTupTEeWw05ELQ5GfR6pcd/Kc/bsKZk9h
1VIVUrWzIgaUj2kmBY9vwG+MJQ+FVOODG23t+C6U9Xmsw12Z9pOQqPs44fGuFc+O
xgfdhHTB1CNKt5+JdTWzLW1XojFF2iquYdT24S8nBxhO8d5iv2by5y19/jHtb6ZH
f/klFgBSTHJ1nRJNe6U4mKrIU7g3kKINf/08xe0vcYTT3KqfBhUh5xA+dwpbBhMo
78c/Ep87uhuSdhl6iORKaw6Q8LKv6lX29msrlOu18GxODJLb44PMD0Gl2x4B1NB4
jULwZnQN9xmkSWTDJFItpGzVohzxQQ3ZfJ06Q07f4tYUwklzAEIR+eB2C5hyYuxH
kN4CHs6qsR0b4iJX2796jlXkHEMk2SHruK4mpWkeB4Nwe2ojLIveg+ZbUIpA1g9Q
BnQOMS0Upfj3Ih/3tQmE+7OvvMzF223ELa7aDio12BYtdwdYYG241cNkqhpEnjWT
apXtEsvpttUIpBoiarknlkG5lOWdvd1RMyj/+2M3bipr8jnbOKEFXnfog27ueTIe
JxVXkRzS8q/zcrhRGsGhJm679DfPDG8/oWERfZUgPqOidaghvyUm14DomgPckQbS
FI1ztMiLxsDIiGeaS1neFQ4gsi59/xj3w/NI+KEC2uI+AaoAjoFxmNqiI6Y0qk+Q
/QyASBNQvgmJNX9tv3+b2rcqafjXwyWIpmmoBullZZ+PXcavV7PvejBhE6Jhvj+3
2+6yxjiIoWGFSQL2LVM5EwyAOOVlSszIC3JUJUxTtu7HuEqjP/95cO+xAoHymOsW
/o+jhnuVzc9tZiLn0o8WzGjxLZ10Xzx6u+jrANuHWt2LnDWM7eqhEu2iH5j9oOn+
FsXIG0KVLaW13GkUB/O15AC86KqmTI95eFoO9q8+R0TnOt4Oc9fuWXKcAvMnaSZ1
VAtBR6hKksop7S06AaBE8nsglyeMJQfvojfd0+9qawD7e2EPnQXLnu1sMwu3VPcX
WZMiScsL8Ulqg1yK49UQfIr7Jqk8p2OdPOIN4J+XEUqvGIHRsK39ikkN1kcza9Z8
QPqEpQtjVxkEfuLmZGF9Nheu9Z8fDZwm7sO8eOmxxsl9g5oi9LrlR4lYxYvUfdsW
E0buZV54F618B77qEmqR/GGKufEUyA40bqi5nZtZA02VB+LDDYPgK/zvliIFySna
fIhpeWQz7MrbxZgsDl3xeCWGT5mI4NiPAnvL/MYlmlu3ni/4h4eBTfgzhKEJn6ae
mpiNgi1WGPQDHxcfLv1wWP+KUHwfR60wFi2LyLjULC5Kn2vXlUOGwIiOvqLUbTeW
Ueb4qsIFKyct/lvq94MDCwiRK+yYEvJa2GyIg234YJuQrliAm+E8ThBFClWWd/Sc
0oHQp7kz2rjhPoFNdzgyl8IQu1BxmBhr4+3VAC8GFnBbQ51fCX5pbicAgl1dalNw
2M7mElLiPP3XrVfP4cNEvHVpxAKtIXBI7kZvxiGW/QaZF+AE5nn0DtzHfuffG159
pPn/pvq+b/d/reOWGzKTDlH6MW1TFnx3Lvy5VmC2IvcXkBuoAcSwDKp+O6LE4dix
7uo5/B7rSGzuRFnMLOQfe31gKBvHHE2Ku5rbqhdwl3NdHJuIgFsfAK6ZJtCnVOdx
2+cVC2FKbl6WatWpW8CRDfNjPiTspomeXA1sqqQIjVZCxl6c/io3tdKE/g2TpcRJ
WYzxrhzJrdDUTQAyTMwCWgw/ZPU9Gh77yiEDWVwO1CIiZaFA+8+AinKPZv68bVAT
O4Zb72VVp5B1g8AMVlGKxwW2jTptOM1l8mmKEK5/Yol0bWWl9nsY+wS2cKICW3mh
S/0jUJ0noIsGaJhiYrSdLyI3NZ6+yNipdy1sgU4xLON+g9oCwAskKtAUE/xN08XL
w2PVNf19Y4zC5KaowTI2zkzUmYEOZGP0YVA2avjp9STZbkeJBJfGosrM+Xi13Epc
fkaTTZSEHQQztC910UGX+uUDhfSS/MLf3h8aFRBbtniaFil8kgY+9Cr8/57FgmAT
VXdGDLdXLRCkIqgekiuxLKHkFWzB6gtmRDfk1vGQM1XQJq6zbdRXCXC8hJXtNY0y
InS0T8Fn+m1mAlhQ9UFiI4woXsQN/ZNgQq/Fpp7Qb9JQD7YCR4rwExWLIUgjMqR0
c5gMDLFuu15ffZMOICv5yrnF0NjSq3kDw57LJ+ywRcCP7+Mehqg0hxSoWDyq1qLK
+8AYfQF1CUV+67S+V6/ZtAALotf+HDVvhR4mjBnt2g8qjnQ1fH3SAw57qt39ODSW
VFXO8ZGIz1Vd7QkKvV7ovK/2dkd6KWSWJiKSnt0+RaO0fRc6KZ6RYklZ5UAij6XG
8+fKsPqnOSVCG09nNdZCbAyVsPhcOhiUVazsmyyEJGkRxqBh/8Wb+p8FyEZbXFTb
BfyDTHYPABv5WHsh2MYciFK5EZ+WEWGNW5aa9pTzK2RZ2JzeIKea0lfSPlGQ2ZTb
Thoj/e2K2hhUtMDtw8M/x6Ng+RBH/HENhfaLJl83MDKr7YyetqTlatfnYBpzH0Pt
1Mt5DUAFEfsOX8tfWP30daWvoW7PSbhMznHo3ru2KD3WorcDoi9wTxo8Ei45GIAN
OjiCMIYmIk8T4QKq4/ZJpn9OYvL0PCJhGlrkfJZWqlGylwq0mg+kz60Rcj8fX6nF
PhTFnpUeN1u6m8j4GV3rlTZFmqUvHEjxtC1F20B6vTSGUXtjyUq26JicVN8G/s6s
qGGlgq/czCgNSoSg1DYp6dJ7K6PgK+D3qTWrmnRZ0NigVwBvTx/d0W7Xg5GsMeDk
CfRb1nE8EYxqMHkLORcroAdv1icyA39utH+N9CAX6jNcchUW0QmjpyJI1TjdRX5G
MLM/jiHs3N6O/3ercva4lyqvteOMJtdItMzpm8YnnsNdhVobfugNznUExZynDP30
QdEDCdD9/1VAzRSPvEKvY61cGGkfW08t2loVmLOVsY+kONNnqE9n4FraKrpLDFdT
/JXT2hEmD64mArzYTr4ZLSj0BrOxjYam7YL1zqW4FnQRHTv0Nr7+v7IqGmA66B0L
6Egarghpe76Egv7C/GcO++FhpnsWNpj2M9gYQzyFcqYU3BBss/8EF+PZhUeS0+Xx
5r6PyNd62Xy3B8R7CGN2a/D0O0pPeRvvMlIiYePVlsPi7amuwKyLVSRCQvdCLTjK
Z8f9HtWq6hKOyvs6PvdVtW9SDXMv+DaPJ6K0VEmnW37rwTIMnUpBR+xN+bHwL6pm
zgJyR1yzcsJQhax1a60Tm8ad/0olimyTfgcl19gOYYY65FbSqVKHiXxe9XgGpB9D
g2krQ25SxJeurc9X2W2YosbtXosyEKKgLudKlBgrQH0m/JX3wmj8IzJGtPCY5HOi
mIWcIJKg0uuHqFrPgwLfLsn6hqDKGM1QQmfWw+EJHalyppinWYmi40rH/pCGdzZL
3mycmiAbjViLQXJn4S355q6j0mJzdKY+vYr3y4EP4GkJyXJomrW8W/5Bo6I3g/+n
I4H+Lcomn6zAwp5kyoRUqT9mBpiXygXEW3FFwd14xq7zOyvrtw/xmvWnd+EAkorY
aq3fbZE13MeNx6pJreJrNPmeDlVWlVou4vc+up6tKj4hEEVXxkhshNj5lTW69Cx6
Eh2tQRqrf9HR/g5PELOi0VYHdqXeLzxbfHxZFz1q8iDwGoBb80DhN0ylAGivZdZr
LaufKjPNvu/VoI9ESTaHGm2CUlmKhH1pLsrYm/fAH0Kf5dBzINlQIJu3ow0/2WJb
DP8wNVN8ExOOo3lKC1gtwgbHzafKv2t79NllVS7+khs2pBLPW4tsETXgDS1o8YoI
pMi56m/SONra6SWRkP7MDxG3+T08WbRrheXcK5LU8yQRJx+jmOn1ZXFEx+p4Tpkb
dt+P8wEDs/UaQVnjel+PDFrdpnh8W3ykRQ3om7xuorv8HZMhb/WJWjQ9hWEOjRyK
rLv4HENIRkJsHTZEXirwPmHJDsX1V4Eoxk6zEJSpvNpzzvVNUdcetfDGDwDsmunH
0srUR2QWSjk+oBOJpw6POjoTfulQZecbu4tggPL0kIWI4+WEe7fq3Ohksp05nzhk
bumiikl1yhhF2XjBhOnPiPjY9owCyM/4aygzqODmilCWsJthD/NbBq2VTuhO9aTc
xd8VU1gkSkcJrMjz5g3qeXS0t4F9CjfGL+HbIg9goWsPHM1P1BmE4UmyAX0mXKut
mGX3ZREoXO4akdTkuiNWmmlPwkP3uNTd9zGKwVbf6erNlmUAdRY5Z3/bb7X9x6WA
isal5DzOpf9igvDe/f26S2PQ5C8wB3unv8p+7Mt3F6nDiHgXXxNq+jqSosr7s2zf
zNvv7rg7MHy5+i6fATe9090YfQQq5x6HUpYKYig57AwGQ+YfL7oYM2T/Z2bwFlgE
c/ny3sS4Ar9G6mMWGetkw0olXO0ugFvIOcZipTb08Z7/zcWFRw9wpmhJ4Ljk/pnS
jQ2peP8+pdRsSrkr4zpjVWuAd6i/wiA0J9UJeVRxScBqVscGBx0Idru7laIGETXt
beUI4r5OhwG1pEeoiKIeN/sFqf7YC7t6/joHGkAivBbHwCYo5Ey6wC9oVtPP9VB+
sei86TkrD1N1xKgh67tOJa6v2nW/PEIj2QQdPo4AZ6QAlqJUrbjeHjecFCAmwxIN
/RBr/7NryK7NvBCEgjepbKC5nADnMRHyhbbcC8UgGLI1IyJmntTL2SjOhZyqZ/Zm
oBHBHAZddm1/1LFS6gAVgrfKXUBqr+nl7McCC+GznafJH7T8rDf6kIwJEdR51RBt
Y33Gk2s8Wk9joyYtQ7yZ2Eh4SzXl+z5LY30QgW46LK0RKz9RbTbXC4PvnjjHckPv
7+CFjDnY0xXzsFloJmVt86k2zqNyw1gNHy2KDywo+zwC7aO8vXxGXcNyUdzvhK1N
R9XvoA/9LSDTnwy5j09/DVPGgW9UT3+FVNSlpp3474wFRfy7IAdBAvRvWvs3dbHt
DefILjkv1x9I3fW9PRjOpsuiAPohoAyOWquBNMFk4tAE5tzvfImDrOfl3V1ypdpS
FFHL7inM9n6P8H2fNO49xU23BOX5bnQRbgywnUj5HLUeKwNT+ZUyY2BfPEiLDRDf
0ViSP3+su1AdNxW1ygQ8BqaQqqp3FmpF8tQwSj07v29q0Jby2pfH7K9XWLGKVywA
EzQT/PkQ+7huDiTaBO8qCKTVBX4CA7ELF1mg97ZMXP3/U1k8vcG2WYxyI1WP9sK1
31ALxrTcBNpDB7pfo6He6MJGQ8Ng+EqTHr8womGtR9v4velS09+WCukThnG1GLsS
ze/nqK1Z1Vf01dm6awu/Hie/P3Ztsn1C+tZk9xovbMeYcm+f1U00Zt8Wlubj0wnJ
u+f3E4rlpvNoRJvSI+xVLwZ+k18CjX6xgvi6vVdQMtlPQhhPqePw+pF4/uPWfV+4
d/unOMLbDWisceGbU8OTZXcM7D0RE9UuqPDGssTQD0d8bJABM0pEW+4Faguip5Q/
bGNdIbUZgzTszmhcBTYCF/kvXMTYOFFLl63KRorO1+aUNNNPJJUROSYM1FT7oVIf
SsEEYj3EcFmt14gTUkt2d+0OyyDGJ8RBlanCnAsKrpOAWXw8lnoGbfVdvAP4gPGr
XCZTpSZcZ2ZZvYO3njbT+Yx5qGr852NudCZ3WCuRvl9IvU1U0Nnm/e3YJzZF0J0z
scAG8Y7yUQ2nIUlUXgMOadW2i/0TtX++xgKmluVmATbcSVKS8Fw8h+GzV5uKfgkH
iIMyZdug4u4uVory8GBJUrxGbbh5bYF9JHj8Zgw//eBt6/X9SAQSHPqg8xuVvJyI
xKTQP2W+ajtvZ5HyaP4nW1Tw18u2oaW1ycNSzYMAFbsd3/17hCeAEGVCwMisgl2q
pbqHT52QBiMAU2mJvnuD7lr0QwSXO9NXw795pWzdWSs5bk+LJVHqJBhRxkt2ZBl1
JS/UXeMFpsr+MD6UVB/+vgtS53rgmX00caqV+BEIAVgnCJE5mcnfNMjUcftiXLEZ
3xm7a4suEN+sCwH7DxQd8TKPQVM2UzuEHB1eSOe3VThPgIw84Oaz5VLRaewYShQ2
yt4DMAxSdghxIyUTu+Bbk+LXmcHHVjPK6f48VtPw/dxdqd4a0GbtYVgmmUlgkTqe
pOb+l4V2+HWqAMG0VM16H7OZvUCb9fR6OO7HPRx96ngtdg7EkOKfApozwslDWfnB
PQy0IfDqOvpmaVxj/ps3nvEtbr4HXZFDDs0CvN7NEEoHcPmGXr1AXbtg8ygn3uu5
Nl+Tm9e23MdS7mGjFgR0XE/DMYOlxTU365qqhd2gfPgQ5eT7fCRO/vzMju034TSh
yt+OPivGZ5IPQhPLH3glNhhOhjS0LZnso//nWZ2FpD5zCUmYjDLD8j6txlO2oIlH
EPDIK+jsC5Lg1YewsexWIE5CXDc0ewxrdp/T+QrLJfz9dDv+wi810bMYoWG7hiph
yaEmFU1EAD5ToLZiHYcXqlWMPSFjNbUiAu/onNXj8fFMkDQ4Dyk2JrDUzCdHckGB
pnho0GdgIx8K8bCjK04Gy+z+uQU6WgcYfIupQqeRDAQkrw39tofrXaokne+JJdxy
C3Anwefi6sOu4iZRXJvPulYv5Quj/OXIOuFpTNGfUsCoR7r1XGmrhFyMlIBEShG8
wo/DEPiggDQFwJF3QwcZNLmaamEtcMvIzNHT5M79Xksb9J/nBhK36+tdpCo7wy4L
UsDh3JsiVeuuuw+RpoQ+C8An+2ZC7rm10dYHzJAWJvkcZiSBpmOOO0xaO7cstTIE
YBUarplH/CDurRR4KvsioGwBSQq9S1adB7+9ZKOCLDLDDju73vOlpXZ22wXvvGyc
jbedhqIeetXuE3mVOlHubjbDoLClqy7L3n/q3zsO8rUnMdZsUA+JM+asIXfkTEX6
r3Y/VeP5jAfJtOHSnsi9dbPp6y13cFofF1jbVETppToNu+zWnTuBjEw9/4rX1hkH
JNzEDDLBy3ryJfay/vT8SDXpw6SfEw9pp4KD+qIMVbVktZDA4e+F9v+3D+BZKqU4
Dlr+ElI26XD7D3342bX7Qn0BXR5HsussI0RWCCikUGWvl2u/q3Ry445fLVjuTgND
zz6ApsU1R740foC6dXI/ocphT2JYdg9tHYMBAiaYunRBFKKnwfI0klmSrPKzoJah
DTzjUFzv6e5CMaKpLtijXOSaixkn/SpRMaDnijKveOALbZg8InTKfdFVSHxcUhKl
RSGg08sSHvDizDdytkJJmle9cMo9aM/okWXH8F/uesFjpEJ2AxM8qM1VxyI0Ntw6
Penx8YbDoUqe2noJUmGH9gaND1+fNpUUWP7MWSRw50Z9/iNR8O7f9YoNw4+/fUsA
dWezsVfvZ9qzFyl7LnMsrxtiw0NjblYVEu/+1WDYUZDV4CeM1UFhDfV4ol8PhG+M
c3oX8V7yFjLKa4RdK1usRiz0JwkawWRjFqusDKsJUootsJaiPXclUz8XID/Vi1Ao
Inu/vlGRzrvEBEcggshF26s3VkDgLhYiY0HqMV6+qKRIZXI9Pz/u9lBmEekaxQLu
TZUcDz0TBTJ0N5BMky2CodvCrmvpnJR5hXc7g75p1wphsnuYpvtyLSkpfQzvDKmQ
L7leQzxv5TomuNZTPbiAh2ACZzHCJIwq1Rf3WYiO3NW2x946hbggNW3QoVvfgRWx
30fwD/J9CqYCGGGdZQ/8hA1Wgy+ecOH96QSN0nuQAD3idt1jyXKNCUoidOeYsr39
HnXHBYk4BNLJG/uirn15ALtHr4+VGb0IMF1pj9SXv9MfQ7//fekt2Qnms6KRjXMp
OqbERnsD8ttgi+fwk+DXljM0+r8x1glbRqlPnXrqoCaypla0FtNTxKHEEnX6FTeI
+kcqdY7DQAKRUNWBIDESiZ556YM8+nHaqh1EIv2b2VHVN3QFIdrXMbs3TficxKZT
CP98OpyP4jGpQQEZn0Z8UMWzmzi9IaBB3sCSYVCs2gDR0egGlcuNdOyEl22LpoAt
3odG9CWoaBw3DXA8TLl2w9UQyHcxIExMHIM5FfALupkigWLzICTimDIO80V+XmwH
zl3YVNWNHWNsDs0QyCGmoHcQTKhkp6+WLwvdOu7lV62xV/py7X3ZOVGynBFw4a5K
/l+UGEuIsyK+PCbWpz+f9JyPfZS4BQK5Ox+peM6vqWPwD+0Df6oKUU9BfVFwg/7h
tqWEW3Ddz2FIHaJ616I0dlxWBsMeFCVqzbgfhQuYBVTygJnzkUbNcgrAPE0F5kxo
cOOUgwJsTQz9eWf0P1409SF11+dgyd4gmr6BIhM6hKax6244YnXfBj7V5zo2DTyB
hLEuCInfi5GZ5ZVSII1WBfgOUczzvGpPH5cIwUEcJX2ogM8HnvB3r9rYL7pvkUbf
Ct1NIZcTjwjVvBmXgaF512afuyQvcdrcZd4lmTqAWFrthSqc/A3OABUqMlgtvTue
UGVoM+ev4B0xiy9NR+kQqPIlSaWx255nf7EsvukxdYCBJe0blq0hCysq/zE8HyXF
LtuuaCM3U6bIW1zCIG/RsE/2hINixFf+Hb8F9YyP/D3q14Hnj/3/5QOKLrSFfLby
+GUH3i6lIKrPlM+1tDLBQ7wT0ML4FAQkd/WV7rW+O/zDzHWiZC4YH29wxbG6sXX1
8ACROcuNZXyd/qRWzkFiOgHwwNJRutzVdZo2kyR+owZsIZMbKpeMQwq2VegZWSzn
U6VVusWybjzz+woszBFE1CzVUHqYfKohWKuy1qq6s2bDxt2B8sSantWVEHLSr/Ot
M5MYAG4ky/XsPbChIph5cj5WbllMUW75LtV8knOv0BNYlS8YFTfXTGvCma1r5qWL
dOiM7XRv+SYshz1gE6YOULs7tHZS5uWMJjBzEngnvjWtGlmqo6axGTP8yKrTaby9
voBUBXyHjY8bYtetJknhgLo0VkXL0Yn561lK5+C6PWTj71uVVyFbMwzQKI1eaKFy
M+rHPE4Ll/y2OUbf6LQEMxBw+3jCB2awb/q7c+RGvr+Uqd5NM8U8qvilimv2FMlY
upIN/sUJ+dwB0wvhuafXWjqZf8WZyYytpeyA3F12XAY9GcMbhPhLmbG1qCqfmIS2
MM46jMVJ4NfSqTBmbddnhCWvg33zi9NayVL5GoWVk0dBIGNswvrNH14NXtzVoKIP
CL3j8DpE2Kyjev4ZdmR4mD14Rc7OxrH5GAcF2ljKMv8ZOba9qdw9sUdW78XYezby
g3m6HrWvl6V9NZuEHZ4mRKi7Nz+eF+B17F+BYOxhwV0ZDjYAWdZFd81g6ztIBj3d
OMLlxTyZVB94lBIUDtK6K819mH17Ef08uFwrxIynEwyRtPanzaTp39MmiY0YBLjE
Fi40fUmJ4ZZVoy5hCCEA/IAsE481xs+29FuyFkD29NCgQxr/QpaQkWBqSogtosWN
MjVHbXLa4Jj4UF1wg9fL1dGZlRPLEq/vdFuZNqfNq7FHmUPCtAcTxF0tGhCwEzE7
bOPaVadC8SExgJLI4F/ta85ua6o3jGBqfgsEA5EOuGkxmBkU1NSXTjSVaLLNx9AY
OuFZt5MFyA/FC6CtqxPaWTNwWE2aSgQnx3dzZx3UvzyzJbspCp+HCw5Q67i9Lw4I
znFtqKTNwf9tozAFYwP/OPmiS8eM3fTmGDo7RbV571PBjN3B3TQIVCeElUCgkvzA
f0nWAV7Ox6EcRBWhOGjBnJbmAWSqvUntAmDfqk2y8QeU4U4q85d4y+N3KdramP9n
K4LvE/cuKBzdc6EDSZivbW9qMCWHKF6U/W6ofXr0D+RzTWPAQu1rW7JK7MILZXtv
5WgsZfOayvuQ7PM8+v//6a4h6YXTWA4NwajvKpIgBfrEzD+b9SDVHcpGb7M9zrpn
m9l+njKwoNZEL7nc7AFqDqvg1r/Vf8Sa11R3j+O+qjYQV/Abn7+qMM1//E+5esyM
aN0U8kovAuyG2xNAxRAKQATheF6rfmauQoi55RdAtGlHRWGVoWDFHzizGr1bsnEx
KTBGW5jQFENwsw2TvvKOmpuOmdBv/Hzt+Y+qatKP0hve7rDp5Mf+ZeEgrLNlnBTM
QfDyOAgMKb40hRM3GiyKY65tYj2UFa5OkACvlNcuukIyPVhI/TCHGuSfBz3M3wv1
T+90WKPdTP/7LIVv26JDHuRv8Vnd5Isf52T4LJgk4z6DtDIuh3p69yZKpuvynuSq
4aiNORRrN/2185mZWtYCshlhnoRwuCmNflhI267vDmVTvbkz8CRTLQAhnAjoYE26
ekscokDwwbKeZaYGq+C+lVpj/b78Q5fINr2DLNF2pKDmP2Nl800//166F7ZyllGa
jCCRB3IKtRqNW61rs0XSS5sUISs+f9pU5kXb4iCd93NyBo7AWbhuWS28wpHLRrPK
ulME+X4+tooHTIWGvhC08tdLdDIp4BBpoM1WTzEbAtju4vAwa4AtrwbDN/XvvGPs
vNLLUs30VW0I5eQkzYSFdSt1H2a0Sh3g+AOP/b+4cCaP9W2co5UekWmPOmukT7vO
pMDjc//wjYft4i7OZ4Z7gld3sGafWiWEAAzfo9zHooKIFO3Q5wynwJqe512w6KZx
KCcFB4EG+ylF3E0A6rj0XHhsidJjgYt4wQrzhwk5mjoiQdck4qXLB8yDbgH3+6PW
bDMvkhAokGaM76MA0DgYYlgrfoTea7aops8WWkOo5N1tPY6ISHCa0437IUdirdqT
gC9MlpZ3DesudlwfPE3d2iGyVlpF8R3PSo/VjjmfCCctikeuvjUeYUouYyKH863O
rUOf3R2Dfmcr+CxT62JmZRDp6H69LiH1zXO0uDamUdlqTjNIFoVAQqlA+UCKil3u
qahqTIzdzsA3ustHWw4CEZ7/2Rds5lxq0iActt9H2XvcDBzIDxutfmj4AUq4U9+V
0yD0V8FSC9aQJoLIT+0fxvzDRjf+5Vl2/WBmUV3cvTgaQPcMdBb3FmDwW3noVYcN
uJNvdPESxF7OBK7z7ewy+tliO+ZBSAUu5eo8A9Glaq4Y4Xv4ep/vni4oXH90voLA
OCc7Kswq7Zb7iAsIf1mZzAY6ra56jAK2EtJzFxC2AtX6GN9IUrGsCWFOu1eLRJQe
VLuDlKXvcvk+ekjri7ZJP5S+PiE/eaDXcwdGG7VGT9VJ0I4dYSYj/vXygRTdapcU
VgKcQ1djEEv30Zs7y6xsAYJekuweRoNCaqaZV/BZ0ihLZOtJQBPkHud8aVRQOAjK
T5zloE1CQJv+9FeXov7+U4B6jmz48gKRzqyVPWPvCj3VcvWsGJ+LgubZBTV3Wf8q
8OoRpQk9VOdiXy+6MgrlnBYGTC/dw0Xz1vUo2erXKh774ooTfInuMWeUm91BCMeA
xwarJYoZEpXwoMGKRhCBYyjGSjPhlr+fLqXwTh2wHnTy8IN91fEojfwQ/TR7URfU
71DubIGl/X4agEa6v5JjI+tbnQdTS7Ia27hoSfPsiOXpCXStSL00Pd3TPVQYn5ql
01LHgFeKK1AHrQjNxggWR9tMH9AACMkKtKfcxykotcDlZNMy1Lt1Xy9gR7DXe/wL
9iEqHfrJpNArUcJ/dkaRNOuacKh4yb7mmEE3k2UYD56ZPXi1Hy2W2c7sATDcBu6r
uAnJEa8H2msElGIB0ueL0AGOXAr1moWsODMcoEkJ8bZfVvwfh+pfqT/kI36gL0E7
HgljZJSuaSRLEsqyWByhc/W3DhGV2i/WW/gdpt/a/FuegYVqeGkiKx4AulOh0caH
MbxK4H5l3e+EDHm3EDfT0EKNR5O6VofFkp724fv0zYTCBw/Yet8LHgAqxKfV++rf
uwRJgAC4H/bw9jLF9MH/1GvnziVf2VZeMeBfJlKRILkG/eDTnQPTJZUCXdaGw9d9
S1Vhb8YGPbaaFuaLlftaVYym7AE8OIAOgjeAnQ4+PaqyvMDv8luYh5Tgdb0djPSx
mIpzGHRu9rxQ95vrmLtj0WWmvdmqyvae+1iW0YESBs3dw8ooxLpbGNITAVD//U0n
g75sm+d1GZ+aE2CIe0tinic92esdM6l4qq49Da+UfTDVVlOt1HJxyQ+60ZFwp6sd
4NWt1vkBpaak6dD9bZQ6eBB37dGUf4OrCcc/UgAKT5lS4bzotj4lsJpjUrQqYdcs
5oDUTDI3OBV84IS4TSZx4XImQTnfMnTsqKXfLpFN0a0shYh8L3ZPSgHRw/xg5b4s
XnbE9rK1Vika6538y1lcb3EdrHhlIua2PpwZy9In4f109xyjk1kIuGzvevMXIxtm
DkXxG+a3nQCVrFsnYDymYIQ/LFexNunuua3w1f+a0BuS3Zd5hFCpdQJGZam9MKtj
dE6H0vj33HsvL10O0gRr4CchSd8Co+rbR9Y36IUy5wACy28ahLVncBdfYYewONX9
nmT6bpq5mFoXOJ3lCksUGVE4SJxx3rNq4NzZTE8TvaPW0YpClSG+3U7XVan+Z6Y5
GIDtXQxHa5dG4I3BSdKU9xS4gxV81IFI3Muo05IlbqPHtVHqlCrR0m6MhhdggYOU
kgRXBX61CsWBAC72qF3uh7NtlUss/c/XIokByxwGMRtCUELY+Oi1rmrv30zOPH/+
FSdqqtHcoe9pODDa15nmQkgl6LPSgGinCppEhXnAFIgZ4s7+7P1JdUoCjiawovzx
FuBMCdk6ka5BYdQvb7TbIn201yVXyKs2S2nx1+eV7wQrUWWCZ/r/20QDW15jZlm1
EM0fJGlEUD8vcXNclqYEKUbJiF/jVGg1hDKnqRK4pag8wA9ZhYBs/G25tDvhXzGB
XmGTRUpgQVsnNXDa2rtOSy+G/P4iPQtrBQP1MbcI9NJ6j/7U9jBHzI5KZcsG/HWq
0p4mwzP45c77YMB5Pfuf1HflnH7aNR6yDhKebhIWRv6c//rypBt7wtfHCt360FQQ
4ibL4al0AvUD0RJItEEwXk71uhZvx36XliMWWzFh6M3ZlXDg8Gd6EpVI1XBVkwdn
aiWzbOKWZcSHt+ugmNoDYFtK7rYejM3LUIGiwDhf154BJ2IZRdztYzSLrdaQAnHB
y5saz3mFHmn3YlapO659brChwvOvHbJcpZIuM8JmT8lpECFxoVf/rAqXq3SZ7XK7
Ag3lstx/GbLApsAZ+w8ozyKCck/RG+A7K8qz+5RbV2hb05zfxe1xJqUMZUah14jK
9d0U719iFvOzXfyJcHqX/LSUiZW9VCkKjmQ4Zl8eZLr6Rc7sxIbhT1qZVcbSqQaO
rsnnZSk27hmo2KMzyurKaxUk0Wtxh2ASr5PVJCzNwU2vvpct7OC9LUEHo3wY3d6X
RRxL1zlj6r3FMSzD7lH6fk4geLpc73hssxsifcTeNjkQxIaH5NtDjdp/5o9htLu2
UbbqanGCm2PtHU85gFNdHPYUqrKbtZXBR/Ya2zBr6WbXOsLTIwydIFU+oRtX6XlO
i1fWb4O0YBaa5yyvne9NqvjuRK74V2BCNyMxp7ZTSeJP5jQl/TFhVF3Koizv+joz
43PVsQ+Kq4Ek5uHvbQdFwlWTmPmsIjhSGAK00bllBD+cnIxJy9hOS1UataIKpMYm
57HVOSUXF6doynWJnVIhqhXokwZwdnqK59apKpY+8FCwjsXivM0XO3UsFJ755/E3
vfNBNn4o2b1lm1hM7+Z1zA9BLjp9aoz31zM1+ckQAhvDje/i3ayo980zmQ6JYrZ3
POzpvJahvrhfj4ZvyV0HYwIh5s8hr3kZ4tbXwYZ/+zXNQXUP7En2fxxMk1uSFmJr
M+MfiszIxCWJAWGlXO5kIOeNqlgFXmYlkreu7Dhjw8GkjmnBBk34/d7xyNsyChSO
cc0fgX1BMVUtqML4kWKntwmt7+WYCiVFKaLQUcTwlAndNSQrnPdfQgk/g+sDC8H2
bev1yro16xZ0ahSRvjWWJXYptoTBHCt+OrZ2Bembh0wUeGpTRL1YV+HIEpfC8hkx
zHvU6v+82I9i+7mTs9BdwH3nqNk4p6KuSKwZRhzkere+YLzplIR+ChaWp4pjZTEj
JtPRmr2ydPFY+LKcnz/nMpJXnhR811EC+QX0f79Io0NcWlK3oFxO35VRd28wZbpA
FpyzWvrhxvmLJew76lJ58N33ZfYalX2qzMY5xAvPadA5BtQuini0VPzJMyl7NrcP
BMfHqbylBQ79odLHu9t+axZsxQ26IlzCQbGn6W3cTk/3D0kZAr8LpO5oKnzAVhBa
q84CamPGInt7V5muRZbQqSRLKjaWSd8QzTRARWJDl53/otj68hTVUUJ4BEjCMUTj
TrXGuVldzmTAfoO7DsZkNMTmDjUYG/vG6ucPto0CRmsAdly7n1pQwS/oyXaKz5YT
J+EYiFoMq3yOtUNZwGHOyPWnlrqz4y8XSuB8oEUMS70PTA9Kq8BphKoDoCCSNkDE
tUNyagHqZ8HfXc4xF0QHlxuLUg/BGU4JOWXCh25BfdsNIYLWCiTqwyHD60Vkttgb
JCmxxArIy/svq5gUJ7D3HTJeGlM/TnxGQKWOovqjvBlkubmXUHkvgE6yIjcDTppQ
PgawwTT2UeyW5+XIMSy7ndWZl4aR+KjUwCNV38OtoIZmLBuZFLVffDqJCE1qwy1b
OvHAR25lbUIywzQCFDKBSiLwkMviiTzWnilKLj0VdIXviQmZlLhTAQT0b67dqJK1
LMN7UlC83EpbNW1vt9p+rXWNiqpKoy8tSPafgNMwfeYNa+8anZeo943oGX58Hkfu
DRVlokrRHntWYlQ7kA+Bnfxacv5DOjn+M37p6wNLTw2jPkEV40p9YYcVVU15OcR0
apVRiJRxBQI/mVkFM/tqchMCSRsmoM1tigFutW9RY34YW9U2xoa9etHLQHtldRey
+k4OJ/TMXZN3FedAPFzZJe+IbPd14dWwTY0XfqkjdTu1jZGAMTkV1FMo+/pml60T
19BdO9wck8G3GDH7hjB89a6mr7FRVY32cmkX6gmaPOd39twrbBFMWGBAgSDk3nbI
YQGqbbtEe5hEpaFya6EASiwgWxz/s48sUyDkiz/6PamNar1l4J7MQEWZC5H7A8WJ
pb0M1sSgpochdws72ul4Kum0BXS98yY4CTza94KyRlcQKhG9H/VlrFgAbLM0D054
vInuieEv98AV001t7e/LhmZuWtfVCdIYCJl+55AnscaRoClEGVg7k3W6B6V3Y8ti
LE65dXrKUpol0hzL7GTKPJvh7OLqXuJ5V3qnLMEzr8UQ3icBHgHfhVZUOnsJyjaP
wqJDQFsIwtwxaecURlLHYwoyeycLgjEiBoBPU5FoWsmJXCgzqTKVQTErOf3UGTt4
xqkJAwpbf0PUdEDUR2OK+RtCIVp3mxlX1TsyXtQE/TfLj3cpB8zKVv6fmbFzQTIQ
+U8gs4Qxr8SQteXjF5J4UtTaOKDN5+i+7LuQCU5FKCNW0QSnefpgwirnFKoqlJgE
YO9lPNnRvEFU0RM28ct9YbCh2mIMXCGTzpfV1/XPLMNaCi4sdJoKHWFI015LAVrF
K/0NgwK1o//6iMp+QbQhwZPeCXhCO8tLTrV/kXYemjG+1fCa1wBQnPfZPZEhx76N
K65guBT7eblGVAYHtmXqmP97M0bt4Lnv4Zjoxg7YB1viVDm/BVWQzPaQy6j8QsPW
iYKGiBCEVqjmJ35txJbb5V+AxFir8hAOns6b366cSvc=
`pragma protect end_protected
