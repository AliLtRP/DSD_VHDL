// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
sCYs7jrq7En8zYz2yj5QWR/DtML5bXMfL7XlMnvavjNfzKcUWqmt2KcQhSLqcd7iYiSWUss3CjcL
sDnSIuyp35cuZBq86wuO8mePS/qjQvvbnG/7laQ/vTFf7EonpG4BUu7c+CzQlS0+m/jY4MPlF5hj
HWphPfIbUNtAd7muNO6zuYBLcxKDHTedYPk5h+juiBA0e2Scbbtzf4yojF4kW99A5foysyNMrGXK
spUaBJOvVGdqBZRObO9lBlZwRRNlALwfTrc7T6Hpflkoa+eIAnLm16bmeBAbWANfXP0UtYaCif0s
wxFYJTUcfxvgp9swKxGk/g26pnM4zxVCjEHDIw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
74LOgXz6xQf01ESLRdmyjjzFrasmwM0zbOXon1WG46CtqIWHV0Y0eGcArFNjWeorKey9m2UnF0gu
BKdai50XAuDQmzhSd9dkRBu0dzfn5BNYErnWk6El7BdSkcG6uh8lA16hARS51+HHOjgJn77oyqjp
5eHQ4E0JYf2qQYv7jXsi6SVC2frqD+zraZ/C/PPCZaXxw5jDRPurkqTZ7KUw9rQ8aeYbZHYW4gdA
7zCfpVqSsJiMInufO6efONOzl2eifaKdgaAHJp9y89u9Gka1Md3w3fa8dR/uS4i+e2AmTYRyl6ar
no2s7zBMAocCuKdD/PKygLTXimjvc9I7h8DXMwnaazOkay/OdUbyyVo2ZlYygnkxGGHBWSls4KHb
4JfE6/NJbkvukI25EXZlzaQDc47sjQsx5eTEjqyCAzelphGgLMRiKT53uuRB/v1kge6YGFm+aLht
f4C6f6zYgJM8I6NkdykHfNrNYvA/F1xGLQycJoWJ2emAcEjmT2eoISfr8F+wcOFgBEITgYDgxgO4
TTXha7XMhr6cprnXHgPjubgjvE4XpWqUM1P2sLehsZc2xor7bOzYo3FOr29POwe7iXTWh/SmwZ8t
CF7ZEZFRK77b5r/rhI0AEaQtXxIoN7lLIud3AH2G9XLbXhUbGa5UwH0lq1/8QQi5LO4wSTIJs/A0
KbfwrgCmZsv/XRgRcuT40QGrYaVngU9CNSwOHlrkL9DyOtjaZTApV3OeGpk41gBsIlpN0ZNmp80h
5405K/AumkLJh24IAjXCLdfeISrVG/4FUcAFWbO0Yv2qoS0qDlnMQrbG55U+zf5GvJDuH2wH4Axh
mNAcuSE3yJaghGDHMFQgwmEX6J/+GGLneuxVCis2OcI01noT5fUGvr8h5LAJjDBv/BArENOrXSTK
axLKOdyYviA+1RryI4OC1K12wIPBJk1yM7th/QqOBPygzRO+aa9CvfcFzd2oDSqd5uC9/EjdGrOh
JuDDvISdqMMExLeXaS77oaMuLzyXHMrcp+dbyIaQRqCsf079dHg5p+RFBaTFhOHikeuKJGXiibfj
SGx6wOzuMYRFvC7xbX3/4z2v9R+tKVjrhH8C1ORD5fgviuk78Lj3hMYLmzjfrPsiPSR/zlTYyjNd
Sp7RR9YTLZcE91fr77epZMYsaQgWw117d02D1/NuZRRwME77Ai7EKgdNk8u1bPK7TX/vamyAyKiy
HD2QR/qZG5ZpMX2yvwPpbVhqnhDW8wPTbFhL5dyNmVDd2Z37HBLJbtiRUOi+91klST+RpMeLiuNv
xwJiyTtVwtP3bKAQ4OvtKbQuCv5/ZuqkuzAUd8hdD+ziHMK+f0eY9cXEIb0Koqy9FuFHocG/83s1
LfD0loPcO0vcTq3RqVLtYeKER6VTRFkcvI61WFgVo4KcMcNbWz5SXtSFXFCSNeBCC91/nBmRUQkH
UaHGicdmX8/HukIrgsRntAydGA9CHpPcKbwcAPnslPW1w+9yT7R9GPqvc0tHn10aUqKt5Q6+KcqO
bkVRWECPzQIj4Fzn8MBEE9s1twTnJKl/P1+K41/uPnbtO26ThGGJZGLLWpdPZfIwL3qtNpfVJujU
o/e2LJpLcOxrpZ5C88lSU2lYR50aqL3fF6//7Nvn78rKvtAfJn3GyU5l9FqfQEMEjjHGHd+23/05
tuh1lAvsqsEBaHLPtfI2G+0Ft5oLErpjmhpzOsaa50kfmiFq5C8BjxKM9wRygsO1yvvYdwvG0UFb
3ndTSfQit6R+in+lr0Hffe0gV4i77cJz371lIhsyd9xJH42/piqVqRFAzb4+vdYDwKIVmbcj1r2T
D+Gd+rbDw687pFb3OxiB/OC2HRP22jfXW8jY70Uk+PcRj6zyIeIrgvCeBmuO4b/ME+JSCulTXMjT
WbI2JOeB4ij9ucC3+t2RTutCk6KaRLxf4Nxd0XnYVpgWiVFpmhWsTMti1Mo2a6KLwSpAd9OMaZgF
iDg4lrU+INnDU7TkFf7bzSrj5JOWnGXBbEhdPEkEBGuhPmqPTbMIQeKPa5smkBZA2nCqCdgMWdbh
QuLTkyi+K82jhBkks0wqIZshJielQHYJzIMzijTbIm5hDQEk0mVDp1AMG3rKkiYXOjOjtvPQfcKP
/JTsZxf4hV0dW6A9nN+9ubOjZxSvK9MgavFyhjIAKQSD0aDoWjl4qnmnzBn4Qrh7Bek6vHqcAKkb
tqCUaYka+MP//ng0TXQauMvxajwmrfkko+qWUoyJkc9I3T+5l9geIxy8uKrKtt5q0AhvgoNjB5ja
Ta+4pPGsr1SrF8zm9wBtXbbRlZUdq803NHZ/GP7qRZ/WjjAcsCnpuQLWIQK8Mycm9bJl9VdUuztM
6DzlJneOtV/NmCLVtUiJGWqKNTlZPh+QCiAKrcY8vJdcJeQaBg3DZRNCgOn5wik2Ze4kIjJsTNQL
HvpGCIvE4Gx46fCljA2+O8HZjxI3X61GEDqqHPatIPjk7CxvsTu1DorP2ieO0pS1iu/s5Lk3S1jd
sUn16cV70D9tG3KsFYp0Bly2LFNPYpbVFFRE8OBqC0G09smXtMKKSkRL05y0Pu7VJyBT7NpBSxPM
dYybLsFBE1/c0FA+GH/GjeEetQ/VuHjuNmYnTfrdUR5PmqNO2F2gZ07tMyOMBqeDzjiclSL+Q/xK
/rLQtQ6fVbuJQeRC7Siq9ER8y+x3A7IshU9tHAnHxAyDpQuqrXtVahNz+ArvoOww47h/21hn5gRy
oZKocg8dZT8UPnFwKKFAIt2zwUbCsi6bcvJ/ertVmzVRe+/GPXvtIpvKMOQ5uXZ2xSpW/J1ArvTR
cuXVepTYH4T1BK7iE0amYplOlvH2mhujYEO1J1azQnItAnQlrNkXnoidhUAbxEDBMWYXhncl3e1S
ap9HkfqUoYp4ZJAo8FYHyAIhhnvEWeCP+IaoIp1qzAeMs3c3B4isbeo9jmRAErT1lhqNK0YIQi3u
2CYw8taaHakM+LvYCYd0OD7Z3aO4cebVxI4XkwO8isjfwbDZ4tXnSH/GpNzfX2zbJzHBJPWxoFt+
HZ0ZEk9haHJgglWHp3vvFYcQS7pmdQTaHB6mWOm8aOV2e/2X7U9qul8uO7g5nEPg8XKqMLu6T0hI
9H7C2ZGli9WGFHJDs4iBOBeTWIg//RJ4ldlJ1NQRshVKCwJisTg80ukGhSHBvlYxjzREMacz5MmY
xWa+1G36uegJ7DXtqVk0IjQHk+i/zZgYfhanZ1hiYS+gJ1oUlrW3lFVE04XaQ4LsWshyyft6ggke
eSCPLgK/Mx9QyZh+ZG8liPrqmTXkmnMkLUNMaDPoGEKVBgN4w2ufcjTufE4TZz2mD5COb8YgmWJS
ZVNy5P+prIkRVnpciAq4n2IfrIDNTB86imFaVBZbAW8XRgNiTJK/6s+c1UHZhu5oHA894Es+5h3g
h2tUXFpn7uWOzNp7l2c+rsxAXp8dKfX2mYcNj6SFH0SCp6Izq/PaYYHoRP2HvgiKpMMy1wTi3iEZ
P0jkX/fFdzyzfjcqRh4YreJfjUgdOWlYYa02BeaCHgcp/IJ2jqp9DbJT1yvLBzvyzcuweTU/Wixl
n6BPZNVO5UzL0HHzG+j9EyrPlqNSYx1gyR8kBNW6i8H1BHHEY+iC7Ukad8cvd8RciFoGqofBtFaV
Ku5Furmtymi1QNWsuxlcSZ467RwB3yzHXqkDuQcQbC9zyG5SO8mzcC8z90eOo3vLLBzQq3+psXGg
787kxCwYZAq+XXA4/RSsgomw8+2+g4RwkvpsSdgTH3mUun5abVBl9j6slevU5l3tQD0zTbakfdxQ
PgzNLhLXTHqOKa5Qhfjg6FNHJweqxjVem+M0u+dVfaTiq6DwPrPD4JjiNk+C7zRGu+sQvl9QvKvZ
OOA01I+yZdhoTX47C0j3DJqxmrFcuIoLYkEE+17MFT2zi/h0MfFGqpi/5+g+jEjKrX461WlQ1at0
q7Grl5W3jG9kpxxbTyebJZLBnYM70Lyv3QG65G7LnDDPRz7aQfuc+9U3m6/6glpymfEJf9MEYd3l
eIWQxduP3H1GTcY56s0wm7J0aHCFepvGCKThwT6ba4cRK8O9590tmfgtUnpZ+yzgcFB+am9hni9a
ZtLOsJBlfuYktV7ryTDGWS6ipZ9CmTQkqaIFNIg9uZAZOZ7Byc5ThyBrZHfj76dDWjApct2TuBn5
CTJwEjNt7+j6TPqw6PBuTr/ujc6O5YJFXWeq5oKEQAexnP/nwFcS+8D+/9LyVuu6+Fl61XAB9KE/
H2+GPRwTcsxrkQwW5ua8uIVSRVrUyBsbE01dn9yIFf3sV/HX7mECPU6wUlarZR/LV1wt+63Wiqw3
LCgjYWnBfpGGbj/7YtPmOMOdNDcsqkvJCRy4A1hFAKlbNeiT3NUh9dvEEMtmdKsBmi/zzrYwOL6v
VH1meXzZp3TsiIeIfI75AoQY1eMkw11euWn152vk8whBjtnL28BbEBJl9uYSfDG0LRRrX3MrA5gS
VxKEaSC5CD+DlPUDjByqe8TzuDN+TgVJP3+Nhx53ppfVjPc0a+ZENDuFsABlKPxRBhWNe1ZrzGRk
0Km9LRcmckbhvblHy+Mt/yu0SyK8QvuK7KDtTUKsrSkdmMB0536f6FptnxzOkJC3pVpI+fcIPDas
6jymh59C8rMwD+nLQNqEtBZswsvdk5WWxm5eOadJxHdiqJ9G1He43WZmexaz2xh2B92S+u6iiJ+b
89JmJS6BVFVL7uZMqfpf8c4sCajorciXda1/V2Td5Gd8+KNj6klHjm3MRs1b6eC1w15EtUff13qT
97jTwwv4UdArrVATN/+RNpN1MRaF1svxqoJk8G2v6JS/YpTAqsG2IaX1EyOPcki99g4B2yoVLB8o
Pfp+vZ9wfiRCCctMaUpIh3FCKtw2eBXyLZO59yXlFdUSvQa0M4Z1BnoGKsWdWDM3GkxlAMp+A34m
r2GMH4b9lQU2CVoaNMpojyqJUgXwZU4yAUY/WvJfiqcWb+9S+SW+1SkP7bnM7WG9edHPtE0k0KJF
JoOM8ludMbloVOlL6diFU08SSEHs4EcIeSxlb/QHBJTgCr+L6hpRUXey9b57V37ByriaeVWeyY3q
K9DyrmAO3REXZUrEL56ilsWsAGtj27/GNtdvfkKle98EXmdKuntvsXbFUkolgotgzPpzWIpaDYR0
L0ZqtxYjh6C55toR+JGo7I+QrXYglmprrK/93dfALmhtTZYgUOkL6ubaQpYPK+FYrisCzRf7dIyp
RhKceQ6+VG8EDyARcOpcFJbNWleDnEXG9X2aGV7TOSTxgYz0Br/REmckwtmR3QOEuVxpGITq6lFN
GAaYaGhEhJoM/y3+mkuD/v4GKV5c86K3Nz/K6WpnI7Cb3NK2HBaTW/DZhQi/alBakzTWZjauBmn1
/O+RTUx6gwPCjOxOTe700Zs8wkS7U9ygOrjVIvDlbtUSnTErrOF4vY2E4AwZ4vsYiOHWZvCs3NdE
m8P+3webdXlPrj67o1qDvdIOzggdEvCui5xcpHhvlbf3zJRjpCtV+kE6OuRHXNog+tUpa2J7vj1M
UlyMMI+ZTPMVd7oeF4deiAEBMfFAp4qJgW53NclG3/0WGMnpdCIeq5o7Li6MG7tiU43/gfZvjIdU
WED33lnEXjkdjiX6akr27KOV/4zJsLt7u/4iwb2flU3CiFHr2G7bV3FC0dPOw6trLOKqwLeY/kio
mirK3rVyEWH8XNlZcAjd3piU5JyKKYqHA8doEzyuFtY11Sz9puDg6mXBsgK0aEtjQNq6PUJeXLn6
1fzROz3CXXfsVo5QS6Blfw8L21fpplqXyvnzF1FnS+o27csC3uPS8eyf9C/b309+69x57vjSigY+
U9s2EihjNbAjRJmwic56yHvpKpRlOzoY2nWBLJy1SHfIoZPhDLFOQuGaq9ZYhJJp0Seot3LkvVZw
fPiLNG/4JY8AqUb3DmuTFv5LC0Epw7wrrG0YaGsjAxhNGz3Pe4+8iCvh2NtC9RxBFk3emLaK4rMs
iYTprTBBDGKl/mcTiOxHkvxF8W4Ey0HfAMmG+9XK6hWVF4pfLTsAMy5Oq4HngY8A8NstDUJa9YDg
4jrwu2+BSlV0Wl28uqR2Y8vlmPhfw+hedNlqRsjNxgE16DRToojS3QT6Px6dftYgsy9oePiUytDp
pTcGp4ibqTFX36K2b1daxbYQx+9T87HzUQZCUjRqnkmar4NvmyKd3sgfV80i4aM9ZOwi/9/hx/a8
1drazyKSYnUgnXxdX4ARjVpO2GZp1fPJLPJ+yhygGRWaaCQWcjW07j1JfEZ2gWwlicKYJbGjILBl
7K6yfr+mYNIzX/TOtMPVWYOiRqO9UQQDtrtykqJ4d8sd7uXjW1RPAc5NwgmBnZBGoNx/d9oIJu2H
C3ig4wv8SzAkfjEt8oiS9Ohnp3PYFCRxY/ZjrWHqJfdNwPBTPpS3CTp45+ud4AX+dniwozJbwNH8
xOUcMwdPh4gquhnLMmBW9JtW8fHrpit9RG68s7N1nUMmWuurj4xbCVtEG1jdpjlaVvNszar+hRU2
g+UYpqfdVKMPmpp27cYlyFJcLknsclReD3jd2pGo1OoDJoZS8Qc4QpQSSg82/xHlOC6QzRPCOPMO
kx9vGXmI5wJeeQ8mFTK4VenXL4yThzrX2q5aa/O21vdRf323zJ2+IDwC9Csl/D1pum1Wl3tvtAXM
5Ya94xwwiDXY2TEV8yIAVy9Go9uFTvvKLaN5iElB5liXil7YuXFcHiviJ4vAWrVL4LPdXHvZGEuM
guiqXFK5VT/KX4IxYI5ri61qCgYIPxE+jiXDuyLOC/H8DHkaL4nZUQU54wkxlAWVRacGYIum4pVQ
8iUnuqxlJQmxCJay9JJYB3Kmg9GrDFeA+FhibpTEv1dXG0PE6xLvsV7VMWuhhLFWn4IOLrzptTqp
AhBzjmFtkx/o+lLw77oOxAiONWUsr0AEgfaQuL/mLcecV4zCvzQfm0MmvzXLCEBYdyZkei031Mlx
fZcH3ykDdn9ZBoZNt/aUHmDAJqYN7Vscdh1bALnpnxFV7NdkhpTqZDsBNERWiOJvELBzH2jDUbB2
GH0q+2tVCc4GIWTOobrjjE/1vfevq7qfA694mkWYBhdb7L3Z3i0Gzd+ODXwWHcom6h3kDI8e/c7Z
8X7Pe6VsCkPvkvHqUqlaQGmEAudkPbqkAl7e3hSWkDvx581tBlTaUQZs4pL03DgYDwaexQ9g+AKy
F4lnzY9G5fhaIfvWw2vFK9z3qGoU2AeBohA9cYfBl5gcmBqRPjukm4lZypvmU5i4rGvmlTtLXMnx
inEbZouJ26cs+TmKFx65pJbhAVNOUpNSGp8Hmq4HkVSxoyj3nWSKqP9U2uemzZLmywpdGxXZzoE6
xcLNb70pCCVUWs/TctFGmPgqhOMhQrIlp7AgWdsjUlwgzz5j1VhziZXH8DJxR/S+8RUcT9VidE4I
f39vZoY+jxh4+cz1cNSYbKevbQQBWjP2APIcYfMMwM4i6RysL6lRyqzmHML0+XeLvsADsOb6eMJM
3x7iwNsm5tw3bt0W7XnnIJblt+LYgR0+AqJpEl3Y8fl4Kz6BfJtznPddPflJLdLo6QlcEXOsALs9
RY4kVqnusbLEfhb/MA+IiH3y0MLbjns5RkLrQg0qJALpnyudL3XwqymXhJnxq1iKM8Mhaf9oO6i3
GU/dqEBX+MFFIGzzOGf9kBkf+L0bQOneSxzruLr/G9sYFp7/+qMb6Gh2hTXL5szMtxY5LTErFhjc
DdU1wdqto93FDoXAnMLNO7tIQ33FWWs7om+uTE0lx4IbdC0KDWTOPZ/9rzOOcgp1ywhxlIlCBvqW
R3UwfMbAVn9JpUQ5rxCsziJ5QRk4602K/6fTFWXtMJIM5Dh9pQrzV+xQHDblzhhOP484XChKsDqk
WlQ7kbPfJw/a0OfDea+VMc4wDnAU6rqmPjhMt2Pe/xpDtgwpac4g8AI1FDSeLPIKOZID2TWN8ylz
8SK/uyVwDi9tp9xD4KrxS0JhOJIRmeZoEDb29/kv/uU1F4VX9KD4XkZ5uLSAGf2atZ+Ozs1eY208
3O5EY/trAIFNxS4AhHM/VrfDhg4PtOgEad7y2V+FdeQ54LqDko2gRivTKa5vFt27gE/56Ol5F247
sE67QS9tsLaLTe4MWHo4xaipMti8FqNoNln4nwVvrCuGtrvsDGJTgAQuTPOP+exIFI/GmVdcpAV2
VyN65AKBwlDN2/7KeGI6/9urMroTo+6jFWJvJ7zW+90/ba++wetLNq/6bI2gbUA8cBvHP9nKzutw
REqG0KYgXzCx4+9ocYjpA6we8A0xAMr2jPtqTklBiLZRJZl6nH4MEnOMf0R6YdJk2gokIpII4RTI
I0HjwIw5kJKsGxp1fS5ExQxjdMQApI4N/B5aytpY88T2+Sg2ys80nOYWF63YoTuG5NCRltOHyXAF
0rq/iJkWyyql5INdO8KLylRAE5Jnoolsa6VQg9+jwglOwllqelvajNAzYDow8c6CEsEPjTvWNdfg
I+//72jF83l2L0nfHNQFz6Tkkpast7znsF9Zjtv8tJYNAU241ZLZJEWFA9Yvm5AWFYwy8Q79n8hT
KYD0ErSDCcRkXJ41FF+G5tItn/7NfCDA4nnxIceC004AIY+71uLJFLNZCBYuUzEn3V0PFnGiYODF
jJgSEjPSwX0zo7pXUEzXfp0F9jQX+bZ22WUeQciL+9nuTFir9VtrnzOZ5OLlcJVhIpqGR36WRdLk
VbCtdbWaPkbj7R7t6K386hzTqjKoONu3xjVveyVFRpCwzOuylnGOwkuJkrKXEhW1hS4vqkK0jhHG
dljwBGVI+trJZdDxru1UNcg9m6JcMUCZM15welpzPrbql/8ZI9uC31ZaaErgZ7E9S9Hl/c3DvhCI
UXyVhZ+6IDNeu1mirkmPXSIDATH063oycyzFn+Q98wHcyPDb20t4jdkBsGg7s3OlbS5KDY7sydrs
6ZHcYD2LKhxHSSZdVQBLi/YDPsGvitqfQRQ8XIyI1rcN2wMltvy+LB1vO/TqOIBLlAyZPfTA1iS+
+3Lb/nqx+83XdsTqSvcJ7teWAxF6B5xEXmEStLI2thhnUA1bzFqVEKRbWZCFtSlOCL0R27pNyQ1x
RvW1bkPukfbwt/xO679YtpJTWJZ8WzXflCegXU0OzWcazg6EF8+A4vat1pJ4vpU6HMqSsMDrrGYe
5awulffzUxTv1RydHWSu7IyY+X+EAp9jfBNuNbIp1mwMWEzL4CMH3MZMwx1U97kjFUo/I6UERsg9
ILtKail7cQ1e4oa8K+MZTh4smLLSygL/lk2y922zyzFzzWFWVS1nR7a/KQKS2Gd6r/4H0driFZ6c
jf4zO8IOTSks+mS2CfGeiqMiyT1mWos7M6R3phBkTRM9872NKy6gIvaWrczZsHE3nL/6jn40lE/t
cPvjbCLs3yQy0aBlGPGkRQBu+7dBMm1b8HFPD7E8FBD12Icw8S5MycPQetDfH7fYAHHeHY9WFbwq
LJgtjvyI7TmivK+zYKSVr/vm9GFBYCyOUdjeNvvOpmwzLmEctZhEIHYLJtTurd1CFUIqJzPEXDgP
GMR2+DieZEB8o27vFm5kobUKBMI7GsRczky3fpf6HS033drbp2svTeS60PoT4h3EtiL2Skdb78os
nn3JX363um8TnfK1M29rsWaTinvlzsjF171VS3ynvkMIfv0Uvi44kMq6QaD2UsB+Wl4Qt5WtTtjW
Z86yT+oQ0R5HmlDIf5WAqMZ1zdHTkJOFhSHuO+QaxcS+jaqm5SRdV2lhL63KCbOa5o/oXMFrMt7s
dmIGMLxR4wT9JWp6K1iiGhfeHsy29uPaR9/a4yweR6o7J1NU1gKQwJmnacQ7bn14XwsKyJUlxSQl
weioQNUKfS7ccOQvBogUM9ePFYI44+Im3HJOBoliedRXqvqn5DU32u91/iUbheLe8L+ESXdcZYV+
h1BhU2XQvv0+0+/BqQKBhGGo2Wend/JKGmmkqZrzjB9mF9xUDhbVH3tELggjkEHoJHAtIRGPdl0+
rBaTjY1sYcN+2aCubfI1YlpALJb0+v8w+wGKjcgAkxFrNnbSvs1oDF/8zd2JFCh42ZWXovDFLarB
0+Ane+wV9GRVDiVou/g5OZU9WQDsXIUvlBvEGCe/fJib03pXj/HkOlis5QF9CH9P7VQTftM/LY5M
R7ZN4K/xB9mYB4vOwYlAg9Znlxt6s2w+UKgXLr2hXVsaGhZ61ZphYZYqvi1e44I2TJL4IL3tJGEI
WPfdxYIVq1jnV7XRWZQndDjXojqCP5af8Is4xO3PDOnM0LV7IcQagnVxTraHpfZa3oNzlI0+s/cP
cI8eUxhykNvFsdpr1fgIMP+XVFN9a4MWD5gGWw0+dTBxVzFKNSVFfxvtaQiM7dKATj4sl9GNPWLb
/hyclaSsSyD/ASOFXXtqc56ymn44OhzfQYw/l+O1iKntStGt4oX/gyAGwpnlvqhiql9nMSvVyeJ2
SkgFrvbcoTSXnA3UFoB4Tnn2OPkcw0aM0NJkKm/MmJtcJ5wL0KshZw8UlIGX1zCxJOwViHrJAgvo
hg+AoQrsH1MfgWxPLM7qHDBCZQe1Y5WFuAMN/71nSb+YOry8wiGUxY4AJRhRT2nY6fCIseenHlcH
Q3rWnpuhbpsT3E3h33qrtzTsvYZcH1F38A0OyLixLmiVisMR2kkWY9FV9LTuK5hBfnVk6cBLtRDJ
ofXq8SruMqBjWRv7jIqSwNcBo9TfW69NSwS9EfFVHk8uqoGb8L/Ba8+uMaKEYCQXiTvhlc33AaJ+
G09a/9QdVpD62Nx84eqN/9mELbq21RN38uEeOFFdNqQb19XNW9Cx3fKvppYG+CTcsaUyyeoup2ih
6ZhTPGtFuR0ncw0zwcfc8eUfgUKLxXWSiUh/4RV9KmLv/pWskS57Q+P640ClZkWnDSRSuUA+uI1h
H9+fCtQrSzglVruAm1BdsqoTG6fZU8QQI23y0DEHiAbaliQAoNnO5EhtCj9C+IcvRlO0ZIHbY7zv
t2VmvQ02+WqTrvCZjqCodUHqCgu9I2OsTqkAuKVfcXF61sPaRP4XQjpdhB3SXW9gMKivosVV8W7A
xa6G4N0zRAKExFnk33Ojm92JGBI6Dv/d8Z2U30VE8kfmuP51jFtC/rHmKCFLnH1xZIZg1VmnlvWt
VXgpFbI/ALIf9a66+m/OyLfPA3C/6XBIDxMCZ9lVl8KBWSRvbie5tn+8e+knxGBfTWihqoWlulV+
2EH/vol6OnBmPadzL3d3q1uLzElVwY5/AXcTzvj6pEMnq1kKyTZkS7z3GLRZDp8WRdvaOvP3Fw/F
yp4ZG1IiDGPEwpbwcd+TBMA4xlexjHA2PsRX3IQ+e8JP1CjeO9oa2Jrifu7dIfx80nBFhTgpaK/2
QTlX+r4b3vUQVizKyp7nkVqYrC39FBmfs369kL8CUL8d1NTveOdnzWhDb/sZvuS9hXw9Q/Ugr5C1
iGlo2HEBYpjM5AfPT2dDdWsvV7T9qFEc1zqOZCEqqGZVDijRG4IWwUTWXb680HJPolmhpJEJI3U/
ATSKD9Rnbla2FwsVkZS3z765cai+pk62qZ9+B5II21iR+bwfoa6eubDotyGEhrbmgb/1gqTJ9Hk+
8QyBnBvjsfz/2F5jBe3koAnWtZVmKr9YIphiZnCGHDp157bp0oxnnZDqh3lfwjtmfFsHC3pCTTCh
/qxZEeedtKE/ppV4xxsEjnMeCEA2wubV2Cw4GBHtmGA3fz18elgzyHUK1QpTByv54iRh/+BFj7bk
AQ22jXsCRjfc48LtqwO5nzd8YEj4cDdmIC1DfXCi5XUSuWrr0aT9r/t6wxYftJp1g3MK2ZOKvAUC
FoWQ6YVdRyZbtKPC3kjIT6+StlFd5hBNvJHvJ7hBdHrTObPXMvoR6qhQHv0eOV25AMwaj4lHomuO
eNETY3URdHDwJUcrtQxXda+Dduor06CDZ/E255XFlEBT9aZ8oUcZT8hrqpC6ioMj+uyUeyjMJcZO
iBHfiLr3f+4T2LZ8paByQ6SD5/w8GH2EpYj1/8WhAa8hXxKetGEdG2GDVnb1yeB5WTwJtGCAheDf
ZJGgsEvNo0dA4ZvsFAXHMrnScsIam/ZKDCNFClNnD73b3oiBs5q4Gp+EtofJoSVfMJ0ioBEdRpRJ
nfqGITVO1URd7eMjb4tiyjOEaaTEC7jbCaXL1TnB5YSKI+3d/0wcb79eLOzDQgus+FAvVwoJi5kv
krKvytqITv4xOY8m0I2swNDZUhFcJyCiiDnfimLq6gbyJt5rvRY5ETX8CO+Hav4EV4DeEGeRa70H
n9wMStYJ2bRmF69tPYJ/rQCmdWz7JrJomylw32bg/kjdIPpektlbgDqwXXUFmb7I9jM3SUswh00M
c+RThnqpmgzlQIXtPwRHsQvQjSShiQcD7epKhoHEBzti58F8Uh28cBmB6ICsP8dYZdqk0g36FCQ4
SXNm2Z1vkxDDW2X/gRsb1URVGgxPSzI/GzUfvwCd94KLJtkd6Jelpf5/I4gu4Qeo4i12B60xBszn
R/jwpU0X56lVes4vxGuDKVX8Y+RLUDkEPZic8916pX4lDxN4/8dFbNF0g4JHMepoXXxJYD+7Vjfa
a5dqPTg1U4dLl3i8rbTlgI6Q0Q+PeEKLo/uXMdlyTHcYGGsvPn+0lLIxQNo7f+6XDjgVhjlztec+
P1tKoAZgGqIyFQ7BOdHxLU/HzOkFwaPTG+Nomgh1SzvT7sdU3xqXa5eJyuWQ7S84wBC2QC7Hq0ne
fx0m6jZqqb3W6F0duTeU+1Zu565sYqlMgpl4qJ28B6uebyva460vpEz9X3zDbcztahf2RFGmH7Kk
iR4Iggr2Fsq+ktpTnzvCZ+bCfZFt5dwvUiUcMoOejzUtNqD5HU6zlXRVjWLvu5mijE5nGLky2uha
ztxsh2lBgm33fbNsdRSb+4CdsH3CmugowBZcgKh/xC+fXtIjKO8L7ZvDHL+yE2gLk2HuTDPI43KO
wZ+QRKramejQ7Kw1x4VTlabb+OdVp8pZVJm14egyhLkrbBE6F7oXEqYlmDV1K367klrvxJp4JXkG
60cmwL0XrWE28AsrYC5KxC2X9tn/fMuUXQzaZbE5GzhGhb/bR4f4dQhUwjnCvwUJinVHj4ZsFgU0
EDNE6M3IgStzlXRPqPvSJZ/H/NRoX0cQlIz2AGaytjcorVUvjCmPQ2honyBW410B+8yC0qWJIfan
JZ+6y975Kc8T9jz5hTctpHTfp0pqVKgfiIFNILM/ssTVM2PlF6YYwDJWTvRo5yLSNFhHgGQS0z0g
4pdgm44A3Uyl0QCBXtaFvhUOvlb4yK85EeQA22VTH7d5a+CP3EDBIucs/qae9mQGfe1XQEniVv+e
qwgGYfrW8Zs/dLCFXmeVNYpfwJAJyCa/0sGZItMWTsGW3R+GzU/SJFWRHHBZsBE4Cd99OazkKXFr
rFaaBWeCPuPsbbF+EKZblXf12gjKOG+ujdkJE+gsbAwKUCBz98hYAP3Z0oWMwLQk2nvslDgFDJFu
81DIEzeOmqmN09ssCUEd4dym1WjBLuYHhP+u9f9e5ABUBi6frpZqMzCl679ZzqfvV91+lIx80MhN
JCEqIabl8ohULnzV+BX+u2PQSoTeiEtMxHVJHg4PPcajPRgL1IiQHiiEDRYYIfB0FNgWAOWUoU/A
rwkGdkHeWn9Ql/Wc9poa+I4hiI7pXbbhRtGapisWyB/BgeY3tUJSWwmkQlyUTiNGXbhqB7FctDLB
71lfydOtD1QbNAuGGPE5fSULE4ER92Ciqf5esM77jlfgaHSVVPvswJNe5TLr91JRusy7VcaD1mrF
wL5zEcWjqnWo9p8/fJmE7uDK2pmFZbTPwE6YUODvgcM4imLqQJemcjLikpNizjZIhwl1OulZ6HQF
JopHzACPhsGYxi98FVQ/oFOKzUZb3PUXQdbRH2cXkxqF+DML+wg0vdxFcMNavay/E0aPar91SeN+
Yh4aYRCDgmitf8BZVsmbKAjgfiL1LgzRtQBY6OT5xULjWhjjw+77d5ObdJGCH32JCgCWfaKRYtus
Zbbbt3uUAK00EncpK7Qp45Amh7O5jFd18MP6MVnY7GpXhMu9lnXlJUopzEYwebdJZuLF967L3rn5
CRlOZOGgGumc4/Hg8vNg8L5g3x6DTRvDOWm2TUCaTXM7VxjddgaUe9XVzjG+u4+7/dOBusqLvLpI
Pxe6ggglD5G9oYeBnh3u1sY3X77PRmpjFS+ENlYtzJg8SlHn/Dwe0K1fS3/t55kBab80qRTwDgnW
G6rurqqUjJqfwBgDVMEEL2Gq1+lUM4AY8WrgTCUu0mK28eSCi+WMK9CLU7nTW4GA7WWjipPyomKQ
rDKPdZpu7HIfKRcDng2ATNX0jzWpYvYdObl41D8CfY7tFErsUnB8bmRiOu0FEb7VFReZEPkbym0M
MMmGEtFkPiNp6bJBRe3K1tDWMxcgNkMnBAFw4+i49/925YFayT14c6J55mfDXbzxIGdxg9ULcX8F
rEorDtzikcfcQuJLEdh/GszBqPDfWPvK0lUPqKft5D/x1Xk+wtSemU9g02KVKVATk0QqU32sMyCQ
GWPCVCSQtOhJB2uYwA2GjDd7PBM9q9ypf1NTsXMG2HNMIaZTtulzh85RsXe+PmiLIjOFd0TUxXyf
WT2GFcALUslJYrQprw2rjxmmwdC/8PtlaFFMV2B9xx8oYgct3VY8MrnpYG6+Eo65qod+HBe03UeW
JySqyUOdO/9h1KPh3irP5/8D1WtiOef71OaEfcDhLqKTo7uwP0iWwSLsa3q227ira4yNdHXKAKwJ
8pVxjhvb+/sPtD+H0pdUdwLDMm0eUTDNWius933fEpoe2gUmYldZF+gTeUD+ye3PHy3QQBK0E5j3
ZfRgWNeZHubkoebCGc5FbgIBw307G2ovIfaasHKVyC8R6PkkWrk6BHMVqQjtBHRuf4D96cegq7nl
2NbQbrkDVxIPwz97y3vFlT0gZYYQE9vFFrXdlwF49wDTeT2UjEBSDSPxsmo+y/VmRzqWI+uBqg/h
5mLBd2ERlgSxArJKs+8M3Ll8FOZhxOQk/d4fdANlrvwYkllcBcuuCURmQw8EmN2YyXUVzkIC2Iof
DS3NIOpkpM7v8xCy5Ufur/VDovsUWGTZDclJo1u4VmhapXwHhm5x2f6F8HlDaCz0GCXWcWXrp/Kt
Lau3clhRSo2w9dDqG6ocyIAaVwcyf9aMOsVY+HAJJTc8d+AlSui1A7jnhv8EdMMuBXra6AY1WEA8
cOqcKCy9uMC4OKdeVUv/WgnVzVAmukne6GjhCvwMom4KAiV0gmmknvqHGJGhrBxHRAqD4p0fh33A
XMqendBVPIMYsTaLnKpJfam9su9IdzFH0MrpMrNeySHJd4eR8kjRCh8yRS2S1U1K8CuRc3n0SemO
MZddY3hSIgXcbHLD4n24UXQ/7sjqMcteFpZH78M7rxvPMfetAMLYpzoOfnFESgDiK8oPtqb5zkUJ
tfiv1lNODR4qoHU4u4XH2XSd4WdQah+JHNB7r3bFa8mzDDUm+oVtYvF/cTVi2yS+34FTBU+RdLNY
JAZ73UoSzb2BooF5g8chaKJ3p5Rtni3NwQlCjKet1bf0rYQp5HuZ3TM/Z5/i6qGHJYoaeamWCMiI
37E4Te4u70mQxY4NX6X1zjfxpVhr+okesqptlvZn2XCN6IoJ9Kx0X7lhQuQKnGCZVpq8xGAaFwMf
b6Pqsv5MFsXB1Ng6Z/SP5klG/OETI7Ev35ahbr2m2eJNHXoMiD8T3kTOGk65bP5TPxv2PVSvUrFs
8TsCKfBFmU/+Heax2Vb4hvjNWQn78VyJpv3e7rY24A19iChy2CkkIgqG/7JuRxY6/TmoozLOgxrY
0+BLTo099jve7r8N7IhQIaUvOMCV4pndahEgqZ9IxUEZIQoy3rtDzpqkSSyfvBnfe/v/FF0gEjUO
0MmBGPtBljXERh9IC/cXFiS3E6xKI2DNjmbM5fFXwbiJbrZ2+u1l6PNao1D6DP+76qWYRH0To/Z4
BCimJJzYdKPuZLJcotsNjeqRvc5bj7JYjLYbP5gFvp7SYOAcSRqqN8L8jBSiZ13PhM8UwyKqBMJC
YQoO1vmqLYXNZsoqZNYHGJ0HkQhzkevwXDUsRz8dLnY4T3fB6HvXmRRCdQTt/Op1uDJPDIMoys0C
t6dbv0WB/uVWiU/j0pwfBfHGHQwVYMxrQFzBjJ5phrwZmeGufeynNNGR0+NjIb7sWKmy0LohhMrR
wkCrGQWfqJ6wGPWCkOFxvV5ELq1UrwlPpoPFvY2Kxe7nr42k75b2PrQN89uBHeZFXpr92h76vRrP
ibV2zNctGPwnTbN4OnsuB8zUj4399ZIHN69jJGeKppgngHdE4GoPeQxe+YC/2JrauGhMapFR4vi1
qxyzAmzyPUmwCjvWPwIcbtH1RBnJgJdiBA7BE2zBSGnaZCwnPMm5riLMgSfg/6jDwUECTl23yaX/
208lMsjWHRK43AG/4bOyDtLbslLjXpwmOcQM9/L+MADGdVUux5hMnoi7Is9SZhiCFduUyORyOlv5
gciSqLN9AkcHDEHcHiaeiLKtIzHHgPVSQlC2aSEMVIyhemrytZ8iLMc8LisgqaGwMxZT2Q9jSWRS
zu9UkoknkfingujpLKn6EnQClLAQpWjhWU1+pcq4KW4VHYBEGj8cx+LgMUJP5KgR7cB03pXOv+FU
haFFgyyxfP2RGKG8ELw4/C9WhAk4RN/eWDLG3BiaVnKaL23gjPnc9zejpWHW+h24q3VBGprbSjAO
00A3JE+uunwkSxHccyfmcQ48s7AW6I8WPmarfjK4HJ9oTroIWN/KghWelZwsPQEAFTgIbLKvpkAa
O7AA2+XbfWtBSqutQ+UEMgnGv25pusACWK7ujFI6BFZkrjn5cATpDBxYak6TkWMJsKV691ztfWjL
1WgqCv33R+j/pvgtXrzKRt1s1XI4FZBWHUnaaGMvR4UFoIoLoMFTW7lGMERUcsaoOisBzYq7EF+8
TzoCqEeLEjamkgrLpmw2cE1LpMWitr3kp3fYfH4Cgbi4vz3knN2pnAswB5jHfQeggg/S5k6BN2ZR
pi+lcjUubv88r0ykhSL9vaOlYeM4UmOLadXwb366eT2K3UpA3sKgTFf2DKGzLEA4bOQmuQwHXH0l
KYT/hn/F2mapoJR5aBseBjogRT0MKNiK+JKky4wBddlvVv+MMRbO4MoE1GCC7ghpazvp8Sk3zjIs
cX2f0whHBw3kaFcIaRzzXVthzDxGCpC3p5DiCTUUbmiWo+20fW/VVDvewT+vuhiSuRgwhgh7j4s+
ArudG5fRvOIrt2h6PnxdlWuUkFgyyaMbPRb4p7aAJ72ojvcZMaGkOshxoNVLS+6KYYqGUjZyHIcF
/GEN/ZuN2+MlodT1tbCZ0pTUOmIe5yVVBc6PNk3mrdgSFKvAfR+OY89mFz+hKOiYScAIWj8HcTGw
WUIZEwY6sZaqd8UBc+ySz9hcRwcmd5nQNn/opeM4lhumvzZEqZiWZyEY8pxmn8y9/QDlqg1FszwK
iD49B1bew7fqVotHX1evVjFmGB/ux+IopPVhkNGxGcFvpizbUXcNS2q/F0W3eRH9FBtxtbQFNrZk
S3AwWoCh99uuOWClif6HLHXm13dIxBppLmpCdaLrZWOY3Mhw2NghfAP38OTjC3KUJsW829W9WDbs
F4yuLCEl/fI2v2RTjb/pTph4YrRkFa3svoI6wvZKqJL9CJo7NdNuGoUwyvFGKSDkPCHpbF16z0+h
eVIXFvnqA3WOxz+Ha1LB92n8PBiucE7jAM1qVruGj8vciLA2n/sr5LZeaO9GOy8H577a9fFU+G9f
Mpg2hF/DG/EpznfDgjZTn1pF1rDECb231zpFKOoFtP2Q4B9vFv2QkbXBs2FA02fbGCCPuCQ+oA88
m9PeFsOBYf7ojUVAmjKCXzlTXivZ7JwqZqo6xdf0F5fVxii+uRhEBH2Ufs0T4+IFmJHksbtG6QY9
qxtZdova2KaS19Dzvp9wCC2lvRIpbr2WMR1FnxPdeoHnL+prjoRzen9VQW30uW6rRKiNvwmiQj+a
OFnoUePyDtZJajv2pbOR/yuWIDutVAx5M7NeHFjEpp2ccShz/N7FveX8x5v58xEi+iFGe7vlsD1c
xvNwPiu/ggDCkXy28xA/ifEtvX8Me0bPI//jN/ohzvCMeMv3nVpCHWWnAJmybKc0Hm/vqjdMJT6O
6d31cGYnbQrru6KQr0ORxa+v9abwkFoRTpXIgvF96ofKoXRPJL7rKUHMK3SaJuKgEVuQiPi400Fh
c8jsVl6v7KH3qUH8uPOEMhJsXNSR7pziqATjL3Ch4Ns3AKjQzA3vfg8K5WbX4Ihk3tDEIvED5R+U
jhEUApz///GGZSkaHqpNoys4uWEHGvSc15FMUQTePwQT/NNmwOT/Q79HUGVgwLS55c83/PEIP6w7
iFjaeJR5mqnA3SYqAEbenEtLysfoNLAaTJSZkCWt6IyztqikyCfylEjgdfsIuiK6lrWFXIWhzkoX
w39TGyx6/ZGXXSCiTL+nKzEeqkG83ltVuuhPPasSHKFEU9/TR7wt2GxBFSMjAY1VoedDYtV+Nq5Q
wX7SMiUyZGKSENTP72o5qN28SxhqgePmDNszolLTtGEMwyWYCGnbkehlHc1NDWJJWhPE2nXClakO
CmLtu4uu1ej5HVbZWzumBvAngPDTnusDUBtU33K0YTQ1paPutfrYtosoNQslTI2R6HzpRwoJREtp
MCzYFe0a44OW1MoyA+BGcKdk/AssYxldw2DEFnnl1F/rgLxbgj/Kv9rE58ahdhyFTV/MHZu3uS/H
mxpeoCAijSmAhwTmJORT0JSVGGWk3iktxev7gpht7nntUt8vbp+4B72+0vaH+tHKRKt3dLYLgaSN
sl5k9pzg2wVrqaVG94a4SOO+kd0PqIo7BZWk5pWl0PmftRT6ClgDy7OegnqXdCMq238UaFo+t3rm
LNQ0aknVxYN5AgcMZ4xZE+YsDI1J/TOZpD0IWN8VDRfqTR6eUr6ah+6OvXcOofssev9s1Kb8SpU/
csNCFIxzDXW7d9F1CHYFBnUVSc608DM6HqF7JeDBqfh3E5BGPAkWdlrzYcIrJ3prTnDKexo9UQm6
eVefJXUNBzSzkrIUaO2FXuva4oOF+kG0qmYZWoWF+0+Kf1Ot7U3Xz0zbhqxmoZ67J+SKnw8gIIoc
MdDJQcKE+/ITALFHjdlFrNvZ/DY4kc+pM/wObkDJZ7KsLj1tGE8KwvSDswrxsxbAwXNtcw9xkzof
BzimYjNoSOBHYfF2lkiLey990rgR+L53ZzqbFCF29odP0K5eSQLJH+Tgh8l2vjLk4nUpCzXoDaWM
ULU8FT6UxYbeoyV6ahF434RM0mf3N4w4RGr2qV2SsJ2Cj9HHOXnXJO8S0AsDNdJwK4XQWsgTXBXg
JSpLMxLgkA82Xp0gypxU3nwTLs23+EKG8TJ24SsYWeIPkSCXEysrnQzP6PpqyDXRbyzmLgUeMUTE
jaj5GKZvXE24rcyQq9gsNJszoFfAQz+XezqCNN2a38nTIG0jlpqqT/5U0fWBZrYow3P21YMgV70P
T13cKX6euP9yZwm4vJmwg0kReh8VbzD8f+7uOSLhG8vDH0uQMZAf/3JS8nlUd7DtSJbpwN9huq7e
hezMTSmBcbAjyNxSrKIY4ZpWxHW8FvORXg+Zy6xPgGkQk1Stv5tuY2XFjYNrLhzycBzQdHVdCNkE
9rDPwTFv/esHNWwNODdX1lBX6ir7TBOjS3UcyRXLmy4ouVczeTKlZfmPlqzhyC7PdQHQxOtgWsgQ
Tu151wiEnhv/hJrw3z/J80747CltZmd8zYhRCKiBMSbcs+vWy6/CXSVzg1VOVcEOZwKYbdJO9SCK
/rtl3R6rXW5BNUPHymjhP6qxkiI6HrMIyvjUcrCdrFspMLccrM5j0wEyulmvjVnx8ifXOaGJ514H
lvzL8vwNIUaDZFOmgWbeV8HY8hJF0PxBxiKvXdN/3FXhsybWZAq4l0YUXTfreT3D75S9OKpT0hfv
wARVpJOH7ZJD7fSjLlEUORm8IbZsP0PdcQ7//i/JROtt1sPquPVoYh066UwBOF6GRO8a3Qk4R/LE
FsZrgQxsqId20vHMcW3Rwo7WknUaqtNJTCQxedzpDL3Ng+LtecTVxaxTO5lhre8+nUoU9Io85zN/
38tpxZvdDpoP8+fQbJz1IQ0v4dxL80ttnR6hIvzkPQpqHpBo0tAOziTgzJHrD3EtINlRY1NtHESx
u6Nn92ZkDDPtxKM4rW8KhoMEmNooW2IAi+vsNBYWdpcNcxrrT6+HnSHcA5Y7Go3f+C6Gcwkerw52
mpfOyvoLVKGbeCb1djiQmUQQQKyHTqqkxKd8asgi+5a5nnvOa+VrsGKq5MRIqn6myo5aU2Rpevgy
kPIRCWP3qgPkz/F/YtMRAG5b36LJs9hGwQHDS1LHVqifapEbB9cAEaDz+yVvGXTi+qpOQt0QgK5P
4Zoy6PDGUPXEAWYJkJhPj74xPY9+Ri7YDIzLGlx+ACGpT5fGCb57w7xUzkw+h2gWynCsDb/HRtqr
i16s2AnZ1tW3uhgvkms3IEo/f55yUb73eo1aU3s7ndgky8ERk07jxKJc07wTmmpeqhvZW8lM7n2h
YvdUtg+9ms2gwgfQctaXwJ3ksM19DIWYCBi2iFuuZspx+xViYPj2abAk9Alx8ALGih4tqIRMEYiB
vAqWm1OkrL1ON5vS2i2mvQl6O972gZw306XVSFDdayJfp8XDbGlLM91CqKkC3PmHamLLD/ct8r7r
IMhNIoNbYVikjkyvSMHJHvWemlkmfJwyidh6G+AZmTz4bExRV/LgnEbjCkfT3xrH9Ho2SninsA+G
/jxY8eBXIXCSsUhqlpAQRQyyCjBf6lqHxXtHZ/t48KSSuBCPI79noS3YMQ+AdIAumvI+Q5tRV8V+
mhqX44FcMWZQan/9HJ3e/HXIvk4N/4KSvT/MMpmDDw/0oHpsbqbCLU7I9drFz4AxZ0iFZhiiUh2h
OID0t0wjk5FdgYIOHwNVOgIDEfMRlcWl5j48yl4G8g5O+SJ/goOI1cc6rBJIN4q8BnJ5/xYZvMc3
+HQpR5x6jGFq2w3qyuV5EvbW3K9uchBRdDe9NyzGJGinqu3ODiAg0nFaZCflULPfCCKo3asauc7t
Wa2irTMf6SflJ8x0oLEtO8CVDp+S3OBU5IAZsiVFPMJom/Z1iddQcrUZ/oOjmQt/Nh6au9bSvxN8
8MpDxXRNU6VmuYsosN1j4+dNm7zdEn9YvSxzBoHujo1B5HQLhzTDiAti7H40xi9FyXDGZ3McdtHd
ZgJaumYvjwAGjT63VE2xNIzYcxbCtMJHGOZjQFb+JU7VQxd4lGP4B+MFmi3AOSAh4MkwJf+pi6cY
LGaqjarBlr+lnj049fg3s9Pu3oTP5HrW/uBkmRMQ7NLvdnxDtpxEM3Y6pFPcYABs4WJhZeCMyMSQ
p+BiolK+Pj6mFeCFKLPjvM1xaTvSww7dVitRkEvRPLhFBCWMdXd9Bm4bUnEl7801RdhxdqqtVnGR
YkgqtW9e+QqcpD/FgMRVxGpxREu9Onx3X+j38aoQ+w/WD+7sEmsa0JbQLWUFWi8pUcM/mmRybOKK
JM8PZ1FLCe/+Ox5QXGZLoOEhDajSwFwUHebeuX87FrqXJu9xQcC+I9+ksUlDkCxhJQgyw/wytkwN
B86Y1mjEXpLVFX5JQZQzZrAbwFaJoRaXnmhnLbIwkzoSt3ANypzpShnaKoqZzCS9sGYC0TvhEKG+
1dZz/va6mB7Iz8ShBWTaVAB4YUOJHRg5f4Y7I6bwSZHkQwaPYoP5nPrRSg/S2evz2cw3fTOC88Zb
lFhZAA9QFS/5K6Kp1SE6vNEJhdjTSb82vFxaXcSoGQz+JUCoWKeWNjkBaOKOr8oG4nnHkF05CCYs
OIw8P4wifxhfWQcbkBPklBodZOrzOWKG4lEPff24f7K2fFBPFQDnMG4PbLNjZ6qzVpYf+27kOkqo
ZKlwTYyRLnxb8Yni/zpD24Qn5BgVQXWxUr62hmLeWwTXiY5UJzl6tEjQjwD2/U2j3nP5/1rZqDIH
n97OR3/MY2mOpC2qO/VHGl86gNJrKeJhdSEC+d1wImDv/xS91ziPYAU58CeXhU27el+1kHiZuDv7
lzUcfNADwBKFAFtgr8Mq4RspRDgwtixIQG6z2QsX0UjbVXCT9whdCed/34q6ffKdrYVo1xYeG4Df
43mRwOBK7ad/rB9xX/uVX6kpdraWlTJytlEXDOG9pHMgrxv14WevzCjwI5+fqi5OlueO6W+U93a5
7/AAAadtyEZJNph2DsUxdwWFiGgzybSwz/CGMlvR4QOLZmAYW1NIs00dnwKWfl4mo3HZfEEtt75d
HhKGvUwdQmWQ1R8WEsgnQ2cfj0GK8rcc24w4wGifDQHL02LTBsyARuXeYv74b0lNdULmmfljxkOo
gJEf0Ry+O4cQ1G9kBojnVMa319sp8V6uY0alK+hChUhNfLvGKdMIed4sdqnVVBxYcbls6GOFZSBx
vjtJrs1V6lnAmK0nnoZ9/1nDZyJesYrwRqJ70shW3ctrrqitmp2uRKWkaY5EN4xIvo8fY82yEcNG
6E71tTYxQLY5+j1Blqb29cxa8oAT1GBD0m7qaUzCfuzBrt474CidCZnQfq79MEjedRY3SssRqRHQ
7UegoKz1aS3nHx4T3Y4t06ombn6tXsRB0ThabfO5HBUs/za/db7+Mz9dF8IAwe8tODldWTGLuH2F
J8kfo3hvW86qqhXpu4uc0j4IREN7Z9TUrCEdv7u6NIK6aeJayr0J7vZ3iguoRUJKJavXmNqCTVu2
s7YzRVNeilX/ft87bBePFucLoJqV/gL1DbENCsMftbezDYoM992xriKgGNfOi97CWHwmtvpok6EH
VLvL9ITXF8OPRPP/zA2qUXFaHjomYvPyX0P159wI9khxqtTkmE20cw70aWdGi9WAi3EPzhJVsqUS
hprretvjsTSVAOi6SNQP0fA46K+3nQAyMkg7pKPTpTGXv+2n6vLXA13TlqHeFBAMgjg3jOlOBQw5
OY1Totys+RFHKo8DyL/YWQGbMkDaQM5hRzIz1QySusqxalTi2tlvioNJrYrFS6m8affuAknifc3y
03g+UHZhKj2xeqrSDjckByMCXEh+IK1UZHA2qFk04VK10g89g5yf02PzSHfwSyMrqEhTrkh4up/5
FjeGKD3OzwwtdTKb3b/4jMXLeblra98HDEWOpR+HQO/FYlaAY9AzD7AMjabnoldgqMscYsKreqa9
NXN10Zs3xdbWKNH6XeLLsfplNyEugCi9iJSMyCjvvePYElFM20DU+H4DB2HmkmOBxRQ/65ZQ7qiB
Y1BHOLVHGgGBx1a8JrtQ+/3+STrRqbiOTEBr4o5HMQkeE2RjjdVg0fFTaenYM6G1p5nm1yUeTqwH
/T6pKrB4A4Y+XHQAjFBO7tVWm+pjQFU+rL+lgG2LcaIpSWvtUPzQ1UAYz/Rml7/ybjlN62ETgGxi
vjbbRbWlVV5/y8S579cFJ1EKiu6k4UpUpCGVDE2jrpYtUJZiXDwGn8NBhLT/wG2VI1Shad+7OeI1
iJYX7RWeKYX0Jnh/QS8kVaLX+s1BfTp5sdInOHw7kpWCMcoqGmkcf/BRmDvrnxOLH7F1z/xZPSeK
pTa1ijEt91HreUmp8lHRm9pX10D7b3RJG46skR/An+liTCtsHBK9idaWpTMSXyi1SGctg4A24nJS
3ncIoqT6GYPlzmIScEA9WriX+MY9lKeUnGMULmAtig9WuZIlAhCFfWJLxq3+cniCU6N9jx4YDPs3
0+jdZhntX6SrBCKzaTRmZlylG+JXoq+pDL8ifeO9zlAzeZq2Lm3ra74afFE6m2mY26hhXrNBqaBq
ymPufO+aLzpgJ6m9cI7MMvJFNFI3MvWg+94H9sCvV9mtHr32D3MRQsYEGMaDfnR1Fnsmcn+jeKV1
c8Tl6Wzcoi8pfw5zdcK9+0FR1ZSiwHrOe/Y2g01pSHKc4dj9L+1ra60KDC42Z4pOQQdKXV9qufjS
2/oodGVlxdMfwPJeU/z7zjeKTxrGe4yuJsXhnA49QCl3W6jIQEDIesWyG2IllOUEEW/p4DnyO/9k
cz3iYk9CaDGsU43hwrq3z1Ely8UyrqDfE5xliEaDYhZycB//Z0bkpkTFGs/UahrCZ4v/upEsIAMF
PDTcjheGwsWRuZ+GoLGHdIReIHEWE2jSVWzmZN+D0uYe+5mPQw9X2xlxfMqhSN/ta1qObyqLEst9
HpB4AU+++sn0doLC79BFpJmGyejDb5LTEnErKJ3KUpoa7yOwMcJwifIQS7Q5/yzMtYtfLuwG8uIM
PKeSWFVX5YyIkR+9I4vKUFt5qQH+RLrl1fCoHy1xkvS96MCawAlHTukIEW0Vsuf4uzz4O5IKsJsm
2OSE1+42Iq0SZUQly4YfD+Iw+k/dlCFBaK6vUADpP9NiDeNG8YeAQysCmXALoS72w++M6fmBdhmZ
/YexRp7ka5Qzsxg4x0WW55SwSou1T+A6yTob5y78e14JCbKs8Ckfgie67q8PzYyeNp+URInPUduv
2e3FwDcyTjkcwPEMKiH6sTlPgaBFt36fh6Janctq7e7Bz0MaUSnOAhqS1aeyZs998LX2I8YjnpFF
sPjrHZ4LWqDib/lUYJQRGVVrHhl/goR7BeO2AbUz1hZiUW0X/5C630IHgqB4239kbKZuCs3oBF+C
xwDEfzGFbNKFhdLNrdGRAqWRk9Dcq1IokVeYgpTwaiUi9+kNdOIWNY+SBiM70eKiO8YgSOeS+6Nz
Ozq8TnDvtN7xvnEjSm+Z+K9SM5SjAn6hGvkt4+0+gN3pgTrAFmAk3eGlQkd4FLa9F5y9Ih/o9m7f
qjtA7Jj2DiWbEA0VkkWzjrpsLMHy1tDbAxdghXvffLY8k47yUXB2W9qYglRy1mjCexQwKMFdv7Eg
an8fGPnwaZWcvAinYqQvsGQLVZenWa3PivGus5mrYAcLAYKANfzm5Y6gfBLA5koUWBvUdtfVgqEV
DEURVW9oL4z3KCLIdOCzNOnuVQERHnksrxpbcIlppP8efrMQIGOLxLxPG3N235xhlV5VN5aKKMmv
mafsfFv76nOG4pSlUtxTU3zRVolQdyTJEvf8PSqFWtTWGndsW6TnuiAm4JiZfXcCz25r1mKEKkLi
t+I6V3eEYzl0lx7zos5vvy5WJc3MIv60bTUfyxygU02EeT/J1i9VebYQ43hOlxHUnl05exBcGsjq
K5eWIBLL+1eu4j/DUvhyIIBOrkb5gr2W9TeXl63BcWyBPhX5/58b5v/OZo4qR/X6H0IWdkdNyH5r
Ivhf+M28joNnv6qcSa18wFoLF7lv5W/UMZnTeA7ytk3s6G8CvqV9sW7A7Vi63HuezZjlTWKshAcL
HWTpSiBfIEku/8YDQ/k62bH3DGYGgC3tj7sEBBADmAX62lnilFtaQFOykNZ7Ypg8x9hrz6+R3M9+
rqLQvpuQxA/kMUuP31fSyLniRKcpnoVAHh96q2CufggSYrOwKWdAn+SkyXgu/PwjO8n6cL/4pgS0
Q1MJ/oGrkptkClyqxZpcMeE/3AvDBuWMUoYbJgkviem9SilPdFl4cpytzqX2aMx6p1CD7UX6saym
Ovd+JWVuzsx3GiKeC3PehcFlTIbB2AqEBCheaIyL7BpWGJWbta3KYSKZeoM1wVMjApamdoLTPHDt
H/isDeqXzI/R1KcdNm12OTc/LFzYf2YAX+YdxAsVjFN6gBBAVH00UnL1BMLhXWULNLZLOUs/DyyD
2KMljiYOPxgFQ/AmPSdafbNrTJ5eXU9fTlu7PAuzdGSpZiL28+fgqCggrOuoC9nHag5XM4iteoBG
iFwvznEc7s2y2WnR2JVdJ6sPyHXIqh3RVAChbvk06OsqvFFq0/xNuLdP7AkY+kOQOnN1bBqZODpu
dbi6UU0FLWkBsy0P8vI3Gk7DCGeZMgVzMZRkkK2AGWXX9c9HjabZ+7aWl0kul8IfH9DpvkFmO5kF
4+ug4HT7zldp4yXZkGOCRooUuWkwgzp4SqwtDPjDct3pdCAK2nyArDL6fC/v6kEY+KtaalGauwW4
b5V3wuN1g2KFvJR4wCIv6gnDMxGOB/7FofPjb75IhP9CFKBCCt+G7O58pMzlsv/+QQrdxvNdEKLz
aW0SXzQX+LCScTZpC7tTWZpCnwFlPFQ2pchGm0hre6kulzPJH69UzawiAeInVUpuVIccSy3m9DEd
HSk6fbFwCwi4pHCKvRO17AAquvKTXXZBteKsU/CPTzxXxSzTJ2v7USyN431DIW9CPtsqN2ZWo0rj
uN/L4upgbZSrpC47n7EA2s4FhtIh+PoR+gDu7XNlZJoBiBXtsudWBXbsNIcaO9DBOl4DLhhqHNt9
nCBIVgP4AbQQDML+4dj/SLt7Grnuip6l6/B+bXCeHPAPG8aIKrKlG0UvQ7u0t/wIK62g4AgzCb6a
xghliMq+cih0Z8b+TEaOxmWo8WnnYENZVYkyfMvJLh5Moxzd0Vd6DEIk6ogMPAovlr6UH8EOX/xh
ZugNnbgYXYv9QWX+HMlwRs5HOti2VW7zhyfqIYMP3gPYRXgDrw/w4E0PcdfQ3/hy147sZM5i+MrO
Efgs9KJpO+UsUb9WDvLbh+DXIAJJ6P+t8jp6gPukLuM2smqANbncNxcwcQ64Z9ip1+1r5irTuuQo
7GCcjyw8TLNetGmty10MKoR7WB8GP6u25YZ6tfoP6bfPxi1jDzcUK5h3ia2pRrtXCYWwltYtzw/k
oDnaWjUKcRK2KNvMB+g5sfFfe8nwhmXNz6UfDcyIV+Ufx5R69UymzWXRPSYQxNzg5+wSpWwLKjki
U/Txf2TgdSIDUfFWJByRvAbGxJucQDCvLLcv1spkYOA2ONr59bmRIzmBP48nuUnDrFhTF8+mAvAb
lEhWWTKldxLqYPeQFLOLkjt83aSyScZwPQCaGp2kiUXNlxszeIZkQqGiPAHQae3tL5zPaSX5lMqY
CjUx918SKgw770AHcgFWS6fDCigaVzs/aDBInxGCUdHd/vqqACXYKh/IhQlJ+7O7lNEkUqpupnY6
4mnHmvVCd9WQFRQBnixVBjAXBoyDHHd37oaBOpRLdot6g9fnDNN0hV8zH41mjvc52Za5Bnuqvd11
FyiLstOTTfJlTYRX7eE/rVNC85inhDLqgx0NJmRQI1wiHXhA9+6Ha6T2EuRqgE+4vldLQNYE8ERZ
ZLu41kgWGxWliKNp5aMxjVgKPrEbYxsO5YWP5yd/l/yXXe7HOFxvgAtNL9kpNnaZY5/MVZSA738S
dokG9yTM/naa5oCouX9RkNx8cMjiWsYV5JzRddTi8gIyjep0ddE0qTNdErcu7Eeb9/t0ri5Vd36i
KzbdtoWb70pcv78niE4jMnDM0SOSi9Po7TWVPdIB1LtGHFSZKlxIuZfh0M4q2vuMmFi2yE0luDc4
j8AfmA2wdAkntkiYqEGbXgYoEo0gK3s1MZajuoetAA8m055NiI3IB/LGZgjH4O/EDpi+EJaMNJjG
K+G+2tVrr++SJiqWGpbsNvzP9a1hPuVgRYMV0eKg4TxC288IATakL+O4xHCpwXPEKCpuCZ9Z/EBB
FqxfE8LwQtn8iIa8AuIroQTMNG2KfiPSDJJsByOTry9rhJqwCBPxfMLS49aO3tQUbOzvU07C48tJ
4fv0jh99rCCOLfnadNYmZ5qFQGf6dAEhh8Pc0PQuYRHDqdOEAWLMQrKwPv2c7RgbQoLp6H6tkXxs
ARMjT/dCFb/U5I/P4y7KMzK6UwZDJo2w3o7anGHJAt9VGOHKAGtpt6hAkXrXJC5YGLCBQ894zM4E
YoDhrEylukmnM65paBP9cqQTFnmzmE/UqjwcOthdr7GrVXzkU5kq7j1z31v8+loXbZoD310OsOpF
qE/+QNqq0cdvr3tybXWxdSn+JvTvkLDAV7QLWB8pK3oclNPPEYfGXoT+Tuxfumvdwrfzasvd/yIF
hpvQ1QaeNv1cC8hhd6bTyZrqt3leHtuzwd0SmH3G+5kOUGNR6nDqtnNOCSmanJTXBSC9lLl0FZOI
Agk5+LloxPtrNg8AdSn/Nk+Io9qOtkiDqEP0iyyvYI4UD17rJjwxeEohdZJDMbBaomeWUyzIIvml
Jnu5xjJwZATTGgg1aB+O80j+lEdBre3RWNMl8XxLjSV3bKLSW/mjLvOciolJ1QqOUu/lPJ6xqiLv
g/eOemZJjIeLjLm8t1fqF8BSeeck5iuUYdbAXHBXFlwP6wiv7dMknD1XOTKqfBVg7n7P3n+jZ3va
msQI9QPJdYvVDlyfLX3l/9V+nZEuhoBGxWwBewWCNSKuqaIzFQI9pZu4+/adBVjnOLcru1iRFcfP
g7FWd3LAO3dYnFa+d2mDUWd9zR1UCkPe6Yh6en9XhvYmg08Qvok/80t2pIvA3eI2gGSTGoMn1OPS
xebUOAk8Rwco/yKlZ9ifHbzLmjUNYbLCgtfZF5HL2SEaTesYAxHoov7vIcRvVdm+Jqp3LnNRsSXh
027cH+a3zV9YJ3V8ZNhSTAjFAGk6rSrkXo8LBFbJMlilaoPaevQSf9Rxks1YrA1XR8jXjJDrTvI3
Wvj8f55d4HRheBsyrQV6icqZqlGKkDdI05+85qz53+9z9cBzfrmM6wcp4+BZkW/3HeDMOtwBWEMh
8d/XrTr3/7gVlWsYJbp+ufl8CQkw1mU9XeHRQVrJU2pNJ/VbbDIYNdYFdTFvC6Szo4hY8cUZKDfi
wS3nCtmbiYxEzDI/CWa/1HOziGxHxTYMf2c5lDol3YPliRJWEbm5O2FRsGvPTcAb8b1M7AlAmhwZ
8XNlz7VbPfDDnA8+vturKQ9y1B+GfqxRI7UML0XTQ0IezozFtnvtzPtNvbsmk5rTw2MncPotl58N
EVWOi5BCc3ZSKP7eZbgAbHNWagVVVHv1bD4Elp/0jE7rD8Yd5jJiIlDSDoNdjrl3/peuNbl3mv8t
9ikFRYbKBA7VEIhHJdR1oGlhNUOMTD8Vrl9m63cYSQzh39S92XVNGLbOzvAj4l5M9zKYiSucCU1C
Bt3X5RQBxqDOHX4pwYgdY1KCCSJtWOIzEKdMbnpNcD9r5CP0L3tsC7WAWNBFkjQmH1bywLxbWo4v
1Hkbv2F7CUOWnk4NItcim8kitsqL0IHOOq+zorhQgIEmcVsBgKC6KhJNMi5N0iVdPoQ5ljpVXT7J
yi7U1I5knr6VZC3FCGpf4b2wqs2qSLZlDnp68KFVC2IJj1ZKjYDDrRAV2p7+FgTJHGG+zwjMI9PM
ThVKMm/KmTFa66+tfPjayUaYWiTIKLO1EmJ9RLxfsLk1f2i9D5fjXphrUEV7Gl3hXuO59GbuC6Ut
66OuDPR0sfl4r7epO+wrChjT3GVa27WC57JzVq8H60Qr6/j5tSk3z6yJd17oSZiTfYlfrvH4c4Pq
47x4YwEbeJYqeEL+tLIahAilicqiyNcMemlR8uthpP5rJ7BgnEZ5Vq4zkQpSb7kt58pvUkvlHAjO
iIzkZEJN6/CEichpwK4a9TCY3dFL7CiXMNNB0lO1C54qfYLex3oxRJ7EvD0Ap07sOuAfDx5e3xN4
qkQ2lj5Jb9rF5aaJBxFpVs7cNtQ/0t/Z+drdulhtHRL33bQekWR2vahWMOVY57oybN9QnVwWlt/S
fu89G+zO+QlmN1qGi6NaVFL9FWthU/lSLOsLJbbvjdlJZuFN5azZn+bZoshr+RqDm2Pw32iFWiEP
iO4IXj5soI3Kh8qzCdH9tGTCSvyKlhzURurqG8iwT3Jx8sqSth3ILuB2pHOWYbBtsRIon7BefP6a
VBVHqZmLZGahR1BjLbO2NNJ7U3oDcANXR3aEJuFPxbarI0+OneQiSXW4s/2iC5l2TitYuB1BsT/j
+GVGTt73eIq+VmfRfNmsP+/WKXNkbA2IwFKBLuuN89sj0XFWKLrQlg1V2r4v6bQMX/DXjgY/xD9G
Sff2ygqbnjxABIIJNhCKTVqRP4AS1bAXgoT6VQ6B5+iBrlji1yKrKGhZ4BsbYLa2ky6nprr3Y62h
MSHkYtNBYkH7GahHxdgWbpGZDvIpLUGpD+ytgFWp8rsJ1LGZBoWF6Ky01Lo6RNmuaOaS0ssd0Gja
0u97AGTa2wNG68pD//fOC2qDD3BmmYPOvsZA3EAvWtf4KlBLgQ05h/q4B6ivo0/ESI5vqdtaNkXj
DZpzIx2sD4aORg8p0i6p9Sap9Q/RFXmSwhhyEvcp1pzMXAhglbH9PexIwHXJAULwlaIRHUtDpQaj
w++OXuwIhTrNEKwkDNzVYqDvs168Yiypgm/k1N8aei7VnURPlcNXXAc4HV7DuoBmr9mMgzGizb7J
tl/PmYzfVQrPClBKFuiN6uyl3bwMrkp8RXq8iEAOJ3qzVD39CMN2oOmy4One6YbAJK5ZBDc9dxZ3
DNatP6Jc5nJQ4bQweWsjKTGyAzdFSNPpwO3sV3utRBOQ6T5GDpNgf0mfJESj2kO3sz6WeQgYoGoh
JZLsxzBtULxpjK0pccGbRJbtBI3mMGWFbFyf8kYs22lkFvEHrfmhyXFMerMY57ABp4alEpgX5J+0
RJYxP98rqoDqHtJUZnQGnZ14RYUsph0z3Fwa/8DvE06Dp4YUWf/THBmqDC8yI+ez/U2y/tynDxxL
aLRrSONYLjwrNrUWFtFinYhnUg8RSdS9K+pcQskEQ99VcrTaYdeaUBb6VkCQhUsfBi2WyD4laSvM
x69QR4t/ntjD6y+H3as1j9aF68QiNG8uhPXBg57aINBxdEhkJJd9rCGh73TCnRTSI8VOwsR4r5cj
B4Wonk+7j4//IAjvW96gcz7VN68irzy8WWqkvlbGYqhARGxF/va9Qzk93uJH9DokbD897p5bKbsI
WcHDK+tVrI7ECC5bz3XupeqokqJWKr5ll4plwQjxjv0Y1VXXof312y8v/UMVLCeVq3Fj7cNrswww
blm8BZ8SVAkomeCIP3RJBZrB438v75yHAanr/fJs97soGlRukowk7kOKvsPQsM6AV2wZRK2QV/oh
PGSaCyWeIK4nOygzitefc4R8H0pyCsrkvF073Jg/l3N/SjuScau+jp7AJnygsEWeD4vI8yqExEim
DxjgfcMXQcTPYAg2jBMNf+HMyApezSuXHXOFQWWNR2ZVOy132k/Em9dRiIbVYvkdEQLmePeeCpPF
TiqYiXz+J4AhoN4nb4KPw4ETMqkhPkQVd+aTlfnPF/BSpWbtQSGOj1qPtT+0GKNhtvytaDwYk74S
ogDi9h53g1BPSPOGYFCxecLwZTZPkvtGR5TtTHmytcc28NJW0AZpviDVJEJWDrz8xr++Kb56+OG4
SBsDjSVz+H7ddP+zd9C21rBbheOvQo0Ldmz7OFQfrI9XoLsTihvP0DtYM2R53bdLUUgCTlPmGAqj
3ui3nFC4s9liWvJjFEgCInvQV/qkHojRs4nWCpeha1gZLxm8CuswGAstQpGoUMU926cBQPO2u0i8
c5l0hAlBFn74kPhVl6jSr2ce9KjQFMp4tF7A41w9EZwigwTCNgDYifOqzwXnoME1KYpx/jYVhqaW
Z2ucgZaFIobP94CfcM1HbkLQCAMWpWNonr+nSUiQ7GCpODVD2hVyISv8xgr6OG6ZerLVATPBy1Ut
dp1PGsKtsAHntrfdeD4+SDHQ5oxh5uVL6A1o6HXAhD5jHtxGkIQChS56j5qWNxVSMb092jdFl/39
KnExJQC896M4j2K6rwVYFoq7Kp/twpAoDh/J8gk+K0yz3yb4yGdYf+XanqFTgxGsQTlpn7Xw/GDd
w/TlHU6Q6Oiqr6mpVBLun0Os4FlDT0jOYSq1CfQCtEgat6x8CcrDl2nOlFaD26TxX8ux3jOY93GA
WBXk1ReYJJtHKO2jF1IAkQNCN3hIWk7Nm4xxy9/4fL2vm3yP+KlWlPOptxAIHcU/xej3+i+XXMSG
XdxJOssUDiM9I+0ikWo89sQbzZcCoqDqw7Oz+BK593lYYYT6IGnaTbgewjkAxcP3J/EdBss9n9gA
wAeN245mHKGhvZBlC8ZRz3/jNAAgfuH77Y4Cl11wLbR/D5aIw6hVMzehP0BVoJCiYQKYgUPKlzhP
+a5Fsh9mxzl7pDsxsY8vpP7baFdrtfcJ9Zjbu/Y8gRvSTWElVtAHe3P/5O6wjsxFRykoPiUtFVxg
jlKKtmigMOZJe45RFTSyzx31a8cmTTtMU6MF8Vjwp4n3k0+WP7vhdu5Lw4FKeo6JseLDYHM4eQ2Z
cYMX6qd3vb92SeAbgOjfcGm8T5SJoJUkmLK5D0FCXSTam8vqLfshJzeE/lwwl7gtg5xxE+7ZdZty
YYJZQK+7eXW9YzUUdqX8nDoyP27OAgjifvbiNSeWCRox5UMysI8vxW1r6O32AEOtA+MMO3bDgUqM
oBpp/ZIhK1VuQz1cYY0P36YzXyTHXveqdUD2/udLBAE7XKEdBtVH8WywdsIH7z9iXZJmW5KVX2G4
bEruIrH+TIws3Ou8IySlSQmgZadRQELUVQfrhQ/XHjMt2TUUHVQCxf3+u6yGydvmQdaQvhx+KaxI
PaeU/zJrUkekabqqmnuDXhtUKSUMVANEyMuPp33Owr26CmTWuMae97MBbqvhn+e2OcYguevaFawY
VyFHNA2tz6i7dSjG4ZFwdkSlmPRpo1OgDUSRq95JJm+F+LF8lHGhsxgtQpsZG+4HmyG8XNqNeI+/
3mCAw3OTZZX59/lVSzN0gLRtI/Q8DtwExnAoNYQsPglSETFce8IVcGxVPxoJTJv9wR1fFTQKmbtF
wzKvZJs664chTgdF2kh2d/q/UvC2ApL2lpLFRQoObC6cT4rFT0uDEctLq6fG2RuiND3rxRvqf6Ff
ngWVGLbduiGK8PAjnI5cyfjc/yS0o6OioDV9uVenlE3kne9a0+pv11U46Ab8U1iGN9eToeMk/Ejn
mCt+paWzZEDGFQINyt0PKVK8t1GP569QGdS4toKJb/YFJ5h/4CxiS0oJIXpruBWsjxSOVQA7l3B9
qSyShY6vXP0E0UVUccT2RINuZ/6u6z+bE7g6bTKLx4QvRpehWkp09r0Gpu3ZYoVg+LWdDNSlkFnl
vJqOR2jKfn6yLA2VJUEwXw/13AFZE4V9AQVQrAeBhbV0hPrFJiP/fi3/Z32DacmjAWhysthjBBlY
4MVemDhtEqvNRBWTkOCTJVPQNVEq3gbAy33r+agMLJSBJJ7X9ii6N48ufIHmMbs032KHTO/qpz2B
6ck7FeQ1O1N1WRqiLtdZiaA1OMSJlT8tAPioFmcnFj4qcRmV7MHjYZz5sgymuut09gNykUSfkM35
3XZO2MNEvHOA/MMUnye6aBm/8AUTxaGtAYdK6jOL76O7FutrSxA3crOULxSlJpyUGGqu/GFhihB6
rgCTaIzPU70HewMLr9M2ql0GPPgvzRankBMdTSFjvEXMRdZyHK7L2tDBzCO9WaiGvz92XoyYE+U3
NoQ2Q0CfgbRy/f4G+2dQnntr58JVXP6XBNZGmUGrw+OF12NZcK5hLaY7tpklMH2taupG8TKJ8dEJ
Ye5rBIGfQneMo/jcH4VYLipzP1WNY0ZkkqmZM2943likY7tWBOVJtbtEepjwjk4rOECe+5Fz/f+5
+QOTmVfNW1iNCsjXVAAtQVjtt62Ax2pSPwyoD+/eK0v//YXeSrl2Oupio/Re7h5IwlnvEmDj+hgF
aZZzMzu1oCScu/dh8s71MUFn57lkF7His1HYkWRJrFC8nlYzWXH+PU2XKDUj5jK5W56JhTFTsYrB
xzDbiehPSiz9IWgn5G9TXtp8jCFZQrUUax+paKlW4XSE9PeckttBkc4o1gh+eP9y3AinqJQAKLCu
RkpEe6GCG6Yja1evN5i9CmGw/s+TIoyPofuGEXm5h5fesH6RcxzRVMtcFq1flt4QPK55GOumMliX
zxS4ZJvWsnB3RwhYdzb0ZEi25rcpzwGHI43xtwc8K2aLKYmeRfBge96SjqPgf3ZZrV6z+wEih41w
zv3WDLt5ZzljdUdcvJ9xkSuHBf7YMsHQXaDK4fIr7P9d1kg+f34tyxfgfYGArQiCOke0Jgq0sXGe
aDzXvCyhFDQ9hfFq1/JiXMZQwQf4eEHtIgFVSu4KgbwVSiAm94kSM+Bqk+yj8J+DDDPHgM6ZPmaz
hCMSjLChcrVBSXy+4UkLgdM8OyIOiF8iEFOgYNSfZz0KKzNvD/HKUPtKLbphAUqoDD7CG4p43LMk
u37g9lZoc9rmZiI4fG6tCKez+nhxKqf4qQmXJqOBcRhzHNgXFUfmte2Ap7j+uUtqSsZovguEzwMh
U2itjmeUjrJtNegkVIo+b9T6Nb2PHWKDU0+i1Ta8srUzZcFSFOVeRfjAqpNQrSAc6m2DUc/emovk
yPyEP3A2trgnS4xBtOnjFJZYzVS1rhlrHEhF6JTUfHG7dQXAwreMIyyjP/rkl6dogrQG5g5OYeNh
ZkAuIdqnWJEFOmyvr6Qo2eTaMd3oXMNp05CAppJrEfNHAD40m1jMfqZ8EaEgp69YoYPhsk7qcNWt
gqFVbyQjPFgWiuU/eDDvjUx9YGpeDtfRpD8C1JKmx/cUHA8CteVshjtQWTTh8Jp+AHQ3EYDqz8h+
iYRyFa5KGf8g6hsNFNzVWBasVcF+stdMg0TwJBm+LosLV2VtLlf4Ft3FHSQFqDSLiCpDJhjjeLAb
cP2qRO7Fq3G87nEG1rt9K1a06j2qKMGds6JcQUYT2DStFSSpt7qhVlgJx+1GhvYbznp5uYdouRaM
whd1iUfgYqkIFPFVGRjm2I6E5RLtfreEXn/ZnrHQm70Ci2P6jmERxRe8NZ9q3HTC1qsUXsgp9ys+
cPmcNoXV/5lM2W4SRyRihG0WZb96zbPmD5pHep9bOUQ2O6Fa+mNwKN/yaSThlfqgtK9tAiaAty2n
ovkbRCL6fhfb/3r/VRBczkM0evJfForJptoNUl3Z6SyevjllVg4FyeKbRG5vXdHcD9YTPmuUc0oL
s671QWZILPT0R6tpc/5EUxLOqSNvdoYPNR4RcQsFEdMA1rTWtojUNDm6+ZGZr/X/ryN/txYb3EKZ
RvMcybUEUcvR2/26Q4GIR0hurZHMoTvtEC8abTgBkhw90ptR0NsPxLRqhT7SRKPXoDwe38y778WL
wY6/Wud0t6UIpZhV2auae0mkI5j0zBh+721ra3qLn8aazZ664yVSfciRH4fMYZj3OBDThW2KpPda
pmEahzQeHCPafpB2fRku0AQMTDfbQ9ds1uTS67ARIxSfPXxzI4A/KNTYZlN4Bbf36mxKSBE85ZWS
pokD7L2Tj0bvUCQoPI0yXm6U56QK3+ImUDCYwlU7yR2U22UAxoKUEPWuheI0X5qZYiy90/uAlklb
827xK4t/lhEjqJRc1Ta1tdUH2u1eSyYEQyZ8U5RD16ZQ31R8uuwSU73cos22hNRlWSpeqTfyRYCY
Z8VR9GY99G50yNf2C1lR2/fcJohZVoviU5NnZVnYiJM6JzcBLFPT4E7YUQGFygbi44Nw/Xz8XZqe
/269KSd9dE3wofZQg1QOtDmbW2nO/Kfh55bNdeh0i4q5chebV1dKNc5lcCrQE1LrzTGMaopPMnfz
B+RVbuBpqkqKov4ujE3/Ninav3n2TEfbCsilWW6awJnA0lBShLIjREQwtrYDsnAM/d4iNC9WMNWq
9Q+kc9XA8IxMYeCCTRKJlFKtRA4EzthapOO9LRtP4XfGaqTb5WUd3/q841a6fMw7PF/LfrjPPW6h
zIIGUR+DEmuAOLf5r4qEWCUb1OwBNnDGckWE27V72dNQFdS7IJcycqy2q4xRWeizffWlNxqM5ioT
fUrcIpUtGrryFrZ80kNriTqBlU5HbzEah6goOztTg2pnTb5yCPwysruFP61luuUOzYnUWprNlADr
gzdNcw9qz8FlxdhXYfrXFxYatFhKylkEzLTToJJPLpkupJsTVgn/TpoOl2nxFu1E+yaOjf2bEjOB
FhDPjxK7P7gkevpBWFbEUb4iD20nt2rFtCkH0H827eo9boOemc4IK7irPZBZt1QnKJcWNz3Qs46R
17PATiA9BuDdhK8a8JYFr/zGqx/WNMseO85UudKCGqenvbTVsI0VanIl7JVeE6oO9lqUscC6pt7D
F4hSdv/EFSExaGl9mfYHZbo9Ua2skeGAYfP4Em+wnhq8tpst2X+lDgsTR8TuWSHAe3vtGPKQvOck
bAvNGnECsZEp7TLjCPprQXSiV6vWvvU+ztrwnsZsu0d1Uolm2Lx0LNC8BBHB4dTyh/QfLdycw/vo
3OmgBo9AatOuB3SlAw+fgb/UQBlWLgHWq7TOoHN57FWlF25e729NOmkRCz3E/oqhladD/LdKPOgA
m4Q/tnY9uOq0Vnzzr7VjNciZowkZZodZWSetZJOH9Qe2189uBH68/XHTDgHpaWszvvVIkgRTmIA5
f2FnIuUjMIb+yhlBgzvoXbANGUd53PXxOoE/p1ZiiWmWn0pkOyOct74PrJVOu/75VfkQJfgX7Lc6
xgOE/K7Hf6Gzbk3wjyVLwPuPkrRBlyNO0CrXz4ebkrxSQCfRVS/tT9y9drhRWmtt2RAG4L6lmiQI
XYp7ktng5hVcLbpbc4zSScwR2l66z6zFb0g6J2qWlooCaq1iY4b8OiK//H+xw9d3EkkXSrm9I8vD
wlUp8qSF9CzO4kRLP21YHagaY4XnF+rtBYtl12O/q2/0dQer1I/t0pdrcc9XFW9WZXCokpnaDW5h
EE05D0gMzGX8+0BI3F6B8iliu40gX29BD6ongjBhRcOXI9Pvgi6KTwM+ROUNtI3rMytcgZ6eRXoz
DCYDRA6y4gm2NeiBT9zQ2I8ECOsrDzg48pMI2izA5kERoXoyOfKmKX+fnTncHWhM7WRCd7cYSurU
thKQnTlCnW4MUKm97C6Js4tId0TTgLLmr+NSfyz+2avaQYcQsCT4QdHNWa/ulzfeA4Llx0p5+Pgd
20Wu3IGHP4AHG6l9l4FFe+MSek+a0q3DahJOdWB8klka8s59YAF0Hfi9O6pkiviLRihrnjCCQFNb
pTc/dfgUu+5HytRbuHZISacaeSuCFr8MEM9ZUrlJblcYderACCNBqkjkJDIQ6WekHRoWs526NSGO
cIM8e97fcS3ayXMgu8DFAtc/COBznY7lM1+aroow73uy+N2hXhMKYuKD8JCX3ZQYQw2v64WdF6SB
uN2rb1TqellEdgWlcqOVPAU9jOMBCkM6Ro0cPhxZ6lImG9t1dwNC+RwriaOgXutJk039JHWy0t2s
GryIxBzwfZGYbqQQSfv9F0DPDOyr6w3DCwvTIPoKUh9lsaA2G8viCF9LxhXwao5Vzod4BL2k41U8
vYCFrjOfhJBeYXkFB2397LO8/NpGwIANRwrl2u0lHIGc2pN0H+nRFoLa3WNYevfmOoPpwKLLi8nm
NBs/RBRhUfcxG1WerSDEuthavN+p2LfNbzH3flYyrBaTA+e7PQTk6GpXbnr06pWDCL8iFrYrFXKr
BvsPwQMCyTDW0NAiepQA0kdm9bQ7gH+fbT9vFytkR4xkOwPNztwNsbh1sm2cLR6PFEKn4mwq0MDA
w8Wld+Yp1UYOnyPmfyxlzwpl8eMfXoNNPZtJdFlIz9DtlZ6H6X2xRBPUL5KedHOe7lvBqmYINXwQ
X7SY+Lm4mKrG45tiIUdFRg56NUlJAGELrJ/xKHIyyfmis1fYFjvuEEgu99kY8oHVuyfWVAdo3GX8
uagsttxSVp1ro06p4zOWgSpkeeuM4zHRdGzveiznzIIzwFGJ8EIbPQ5f9inpg2bv76GVi/DSeMub
a3g7mtVj2t1N2rqyuRW/AK4adYH94ZRgOcl514EJ/U57Wmg2FT/+I5FIPvi8TkOliky819J2A+mL
Etcp/DSojlbY5frjXDayqbitEJk+HLse6xSR7ouL0xet6opkNKxxGr9l2ILuV2nGpUP8v0wiY6hB
II8lj6GvdFHVsjbiBBxa+V/9xiIQ2tJfRJGTt3uyYNwpLFE9oRhRh6ORWobtHvL+gJoadotGZcCN
4sVQVaTC1quXqNr+2jaLJpKkFKjbNxDU14I9OyI0/4Ihx3AzRmSd9IHUbcfSpofvvdeerwzBY7Fm
RFMYep7t9Nqy48PJAXCcY75kxk/yL7/EGDblNsCn1UBAc6Q4QQdFD25joJet9MKvomxH6bqORwRx
PaEDBwQqGKlyRX/qteKuDiox/4yWDv8fbEauHzAOxi0QXhVK3KCWlAL/ixJIaL0lm/DgMX92AOcS
vGfyfhLHyNX8O9xelbxOLoqZNlQKWJH3hSLb/H3AXX1r8gRGQLWLL+rw3OhaBvgneGgLnxkJZjhR
WGUVOZGIshT5/J8GNbjC6Shg+neQq5tvBb/KJowat3PY+azM4zBwkq7Jp/ZfnPMSkwq49M+4Fygx
IBvM8dyO0kOHwlZXcxB9RVYff3Oi0YcPgX1Yd+xppoPLLpWP/y45n224bexuhXYXYGXFXNMf+QEG
B4BE153pdg9rLdzr5M+zNB07Etczj5Xm0NIFKvBq58IYj+rNbhq+nd91J4Iarfq26m7zSJgQ5E7Q
/1UUorHMPo0NlOaZ6Os+AEGJwOBdHLmjm7yihKxP+bjJbX+Q7+A9UbhtuYrlzoJGVajDd9h9/Xii
mMFik74nNzGyI6ISAJOKyf8aY8OTJYySMxmpEwHUL3scgFKMCsUVg2DkwaHkQDFMfJO4ip/Yg/vI
VG0VFwDUlNCJmpHD+Pnng0MfvJHCEOyJcwm7/d/9o0jDBjELMzpa0Qxd4365wJlUst+kJ0elt15y
ewrhaI68iALfuO33qyhmMaiecdVGD9MgzviYcq09rELajPWSI9TVVlTeiZR6HFt1qs2mdjIJHBMP
tPKzNNjdJpylDIo7Wj/dZ2GyFXQiKFxAcRPaephPpG52gcnenE7Vr8WIt6wHI8JOLGsXDrRCFlrf
F7r+kIkMiiZbEwF5EyURh8t5S/G/eYH7uoVEYv4PjbwerJedy4mcLuozFrb84I5mgaqZr3FlBFjh
AF/w7wBdruBB9n4leklLMM+aZQR5V/gGqoL5A89y/k2q4AIoDzYwZsx9J0hcIx1qHTc4yE6iNvMn
zF0YBRe5aJ0KP4sXB8q5NwCAqxc85AtpnqBkmLahPKzlmmfSejRnweeRpz/oZIxM4+gzxvgTBCrg
pee0tPMu9zOWQrGRuzumozTna8EN79A1IXEZ2KiDh40zWUTWZTlJulXHFyrD6wRRCy/Qf899MKuz
4kHIX2g/RlX43lQMaAuosnd+q8rjqI0536n4Epf9fHiG0VNuG2kWRmMlSImTWLHEA2Dpt7PLVzZh
lGi1haSneA3HH5tv8SMON0ZQoSWKOZtw9IeqdV2JAbtNlrYYE5szHan0SxMmzDvDaK7YgI120hnF
QCfISFwkCMMaTTrlL2b9xsRoyfW6S2LxEUp5NoyFTBDxwgv80FZh08TTyFxLZWS6UfCDKAcgrGG3
HkTdQfeWax0A3nLzMqUlP/3fQ9XwZ7iPP4h2rDhSNrsPqaDcJ77GzbPD7NXeV0TxXVmXbOcSwsXV
PU929AIn8756lTkonAzTGf+pgPTgTeZC3i21dIL999Fabz8uojfeTg6fnq/OjCmx1DKzZJsyPffj
1WWtV6UT9FJv/ntDu5xYZS7psB75diytdziCCA3Y9DTDxTWf4ZwCKN1tVMthBhKs7e0IhaB1Vjux
+XzNxn7Wvpo91tEacJoLbnHC5RB231rm5y3OYpQAZOZhH0VvChk5/GTIGYsxoYZuKVFMOsRaDe/q
DDqrpc3/Q4xV7FLIfuWVKG+x35ADyYHC3F6iNlRjAhkCFXXBOfuPQQZYtRkYu5k3eZVoSDCHXoXr
ex7Afozd8p4int5CNmx4K2UAvR35FAc+bIRJypO9fFucgOR08ofjJSVTIeucM2RcHwcXzyKd034x
KPGewKlE64OPdYyeUPFtzdGqZIUvTNosn3Jv0ccQaCs7w6Jq7V466uOPZDPHYIsDdTBRKzOtSJIR
jPQpErX6KChdUklCgseFGvje53B3lE0Iv6khy3OoLWfOznJf2PgeZ+BjkqqAEeaGXcwZH6Y6jPSa
dK/TQs0BsHkglgWLkSAVTqfAmemS7Y4zlnNM8xe2Jdd4JwrLoIONZ/XGCB+bxl5IxkLuYGcFT6Su
dmaHJ5Q41MIc2omlzvUcn8rEUH2u+PUjwm1udQLmIPTnGmsuISnlq9ro0fhYjX+6JJ42vC1P8xT+
RbJW1EQ+CCtz3S5m9YbEmn0R5oN55tTxY2jqmdT6lLFtdTOtnETXHkev/s7r7feyJEAcYzOlm8n4
y0ZEwTdXbGB0vA1S6txmSRovnLc6rl+k6essqMxzO/2PGK6yzlDKpYvZG+r6d+6FUT/Yv01SpdPx
FLw9KqjFQQ1kw/ZWiGJIDC0jT7jzuD90Pc2UX6HETIngGN/kjyKHaxU/xVwrWhnd5lFE92sT37a0
a7+siDrLPGmplat7UPKlW36gXFfO83SWpXdwyDZYYfKdvGyDOCMykkGN7k6j/E1i6edcS7jLsd66
yOu4VF+41CFZmge/g6/jcROhD020TcI4ke0A1nlJLgn801PlbS74ZNTX8ISzqnBsoKJae2SfVTmS
m/quNJXQ9v3bJ9DNcv/m3PIU2Ws37yns3GO4nUcDeVb5c9IZ9gbBRQ6/kd4j3t+j12wI8VZBW2ob
kLvI/6DV+CDJQJM0klmKUTJTou9JIOZbJ49RWQG6uw5FOK+uihaHCkNjyoT378/+mX80KHk/y7g1
6AZJYJBBxdeejFVWy1aVQwVaHhv/diTTlEwFLyvgb4LHeZz64xzZ2WRjg4oll1qWkKTPzVxyXUXa
swGCqE0e10uvcw9uPwpxcCTvQqOS8QU8KRE26XVP9yDVuvhXxclUyQERbr9kdT3KklK4VnceExdx
AYhrqrJDywpwXzx4xYHLwcKQBXHDUd3t1tWIpB8Dnfiz/p0wOpKlWoB1QiX3O2fBkt99P4C9rgqv
6jaqdC7Fl+xGAd+nTSLp7pcWFuDmDfrXsOELq3/VdaY2KMpdldUdHDCsrVNFynKytPG5G9R6v+Tv
9Hl7qvDmWD/KuYB2XmyKA5AlJ+D648lKxf3iq3AUxD+mLlyxOZKc/AApc/BKD3DihXthugM6FuWx
5HTSgKDlgFViXSWAlrN7RNrStWBKxGecXPzgkYqKeieihzuQUa01GtEvUE35WrTXwnxcaGF/5KVs
RvP8nLNmD/A64KVEJkzxatQyDBzhQ4eBxCwkUdSFYkovIuLajoXutsUExw2VmyKIb1BjWmdbOULf
bDDkn8H5LvADG6kJM21jEgQe0F5dWPe0QRV0OanT3nJmP9vJ6rv+lSlCDd3x8PjMFJJmiB1qMZxW
2x1qoSSQG2OawCwbOWUJGwVvdC0Nva45OHejGXQ2jy1+bf1nbz9hbxwxRv4mdn9dhLEl6TNoz3aC
jNANLYk6IUDeJS7fpyG1xDa5OMg1jap7j3Tx1Z8HOlDZRwUEVRqUBvStgbAcHr6FT7IHsMwN3MRl
dRing1Pg/tKbF2/54Q3lH5j9Op/keL7pT2N5antPgxV0O02R/muOq4bb/RDXUTYzzQ7ZtQQe4L/a
vApT+gz6YYwQ+PmgJ5CRCLoLla0vIHqWEbJtWWz1zqkaIymB2rYnygqolg8qTSLSU6HiHmq+Gm05
n4/szBluLRAtCmaKkvVtt6e68tZlmr8fHHEXs8gRWjmhHWSoOWxYQB/QZ8pi5QL7vbXY1b4E2LSk
F+W4GOcLIpbKqV6OLKbYD8ohjg2/e4IW7lLdIjen48q0BvwUDo9T5XYAJrc7f1S/3szr5MxzFipC
kuEhddJuivB5mUf213oI7bUFYJDbWX8AC/rgxRGJPrsNwYl6djgd2QnzuEZcOq03cmvkrhZMDhue
th+S8fTmCsd8MUM4SbFKDo4GRgvu00HhrJQFyA8FkW9Xae67epOhNMOaqY2o9EMi8BvbLx2KEMla
WeIOxvgk2Zhhf6WUXLrYG4g3iy3l5Nb8XOB9al1C0ENyF96D+R0cGehBbf5z7JUmf2UWhk4TNjyd
XezlUtADdQ42Stvhds1V52D43Tm+p73YtsSBNUZ+6s6sdGZJlAysVeHXQZCkEsD3BH/ht7ecabN7
f1+SFCEfnMWO99cJhvRVw7dnGMEaZMi5IrC3KHgP5I7S8gV9WdpblLGytPlGo/2XFIx697VUUxOd
1MWQoResl+CM8g7fjzz4H6BdQ46qbW0MWE4AfGsxQ0Zpl/QxIi/YeZBXWKQjnRwn9vfTQlx6q0Q8
PdqVHJ0yD+HrBSOcMe33w+LJKg8J99fNFhD6B9uv5TptJeQeMJas94Id46GcJnadyX2l73cUkpEh
gidmgkjwGS0zpmCRP3BC8ptXrohIBBF9XFu5XnOW5chXr3aF4y2GvZvht3GiXDYhRqpe0VGGDEs/
DaYFS/jcTkpP4c3VlHdcWotgUi+tCI739/wA9TBZBehpGo5TQOcghqEs6qpRNrxeh29MTMwQ1f3Z
J6Y3CYlCGKz4ox/eDoWvpC4MxqTdhEqvyDL/NWMy3rit0p+3o+qI3geNOlIgmzy6JOttOXGy2F2T
K+kLr1/QFWaTsv93B7Hque38n9Sbj/HTg3FSM4BZZZR05cXXocXajrTQc9JEYZ0l7SWrYtZj1B34
fXkxAelt36KstjkARuswHKCY+diATEVFc4UmlmITcyKz7bKUMNqVbKQrbEx7B3e+1LzuvK/9fwvX
kshq3kvmgo26kpJhAPOz8CLp/Kg24vk22rQg3+hwywBbgQNKZwnQ+CsXqazAeJs+GGYy0ocJopsX
ILxouH63Ajk4g025xRr7B0Zl6/3Vz5vNjbi35li/pK6Eg9tNMqf6l27LxCc24V6CZpDeBh7EFsXK
ls1acFBMnOlTGTQDI8dCFHITdlbRGL9TFsicHvcLbL0xtJxNtKAv/WLe6ZfRS3sjYAzmhssjUeeT
N615BIrQB68XAa4HmTZm0ZTdziiKFblgdnfMTxYcf6ZrSJGFXLBpCfS0VGFRzk+tFpPA7bQ4NkZe
0orMsmi/rE7HYcHsaTS0j6fKalvFeDXdSHmZZCA6R7hu0HVzebBMheAyfkWYC4v96IAawwFzHEld
ooUTrII8WgF6zXIbvQtKl4pVDby1aStXXQXkihRuSSAUpbapCQszOQVn4MwWdz710xmS8EDQpVSq
xHZMw3zAtrhYuLc/ew5ARiu43PHnSb5k73hETXjRTKns+wGiifx2alTzkU3/zj8A6+fbQ5VYTrA6
akki1Ang1ExodPAWyVe+lC3d6PC9ZrG/pV8N/ww5fkahjgufLtRm9vgTZ/1CXkuMgShkYRhM7wks
r45BY+Duk00hXuxXAHoO9ireIGoiFJiv02G2FemzrIYFPPn0Y96DBjoDP2A8+zRmS30QafuwDS79
Z7zO7rUzs54QcWloUejkpDHjH6TzlSnf76zxpGMKEP8WTHmtykg0S7hW0DyovUUASPvhsAuZ2Y/9
j2qE8qTTm0rL1Vbc7KTiew+T5VN7jwxvk0rK8c9EjgmyodOzMeY0HH5JGyKd25Tz3WSix9TouOwu
QYY3QXQL2dVpE/fE04kZVhPOKA8UJh7sCl03R3fgA9eNGylx7JutxnA0xEgWACmQN3UULOLxUC36
qDtn5TnUFhtHWfl/ZMK7Zc6Bzw/RRwR6mA8hQPyErjN56CLwWKfcskDcCGfuhEUU8unAYIgdreS7
qti774nLf3xPN8yHhHBwng5mcNUt516/UFbEgMps18ahDJ0dSFZMDy4kJcrmLiOXktRJ+hp7Oqzj
qafSouj0X7PNqbFREMmm5Te5vIo4cJDV7E5of3t/jDyQN5TDsf+UMFJpa082Bk299FczOBaAXCgh
FkYKqIPqsTaHIpWVHksCXwvpAK0DoKmiIdQfPGn7LiQa2Ffz7fg/A/KZBdPmMC7qzDXSkYT1ddbR
pW9y8GjkiijTF9GD6FLJcS8bPb4Jm+dgNZdZczx6DFFpPuDDgPeo6nAOTnlvB6lyLC3klQoXldf1
OCoVShuL9NVjnZeyi9dbR1wpERA8CKBIP0Weu5niVo8ZkEhP4LDNSPn8A3LzLoDbKwQ1zdsI+0xL
RS94rsmUziiA1LZ2yMy5Q/YPIHziMH5lAy3BI8DNABBphAWphb5S4kTM/0h5yLI0lSTGoA9tx0qj
BhSWfLHVRqBYG77ItvGtafyyaDk1hDsTtzEXIpA2Bm8dcCwBVZd8Rrv0dYylEct+QUsCY5LGjLOe
siu64SDuktwIOhLXB/mu2Jm4sY0JWB+05/UDHRwTGued6ZpU2ZRNas9qTXjwwTdmCOPGtfeerVrv
Ybmf+kTULI1V/VK0yb4h6CvNekjsqCQ9v+w5xTTwFl4EhyhCfXn+ZXEpuv7BSfE/dxBw370l1+f8
1ucbFnHZNDYC+W83Vi2Vx8vp1AJaTBk0GZ8dZbOb/6EOTfwp9dd85r9BJL2EUw23SKeZn59Py1py
ciGX9/s01pQ37cDExpIjWr/3H241rz8AsIqCSofRen63GvpgyeVh3J4eyp4ONHpOlmV7yPWzEtxX
r69076Y47j/ot+A6M1qlTxaSOAtWm/OiLIECjzMMUhKh76siMnOuYPp/C9oga1ZV+8po6/egkiiO
Ulb36maHrmCLo481toSq2LHMZstOssbpNwx0K/e8IFByfV6XTvbJjpjinn2IXG676UfCCkY3p3Sb
c0zRfdv9+6DeokloKPPFxUbYDTG+ZoSzfPvsTv9dsiNdW9PJfy+oR/K/oxw1ruZKe0OfinBcapL0
cT8+G6nqHIKyS5ME2yXMWDCtP1vStvLbe/vjVSJlonDJL2crpEB8bN46XRQhPtXhkBOJfPRQFGEK
7rE7lSK24NEw734UMzXYH8NrZcOA+0sENy5ObK9Ois5AMZsEZi93dXEMksdwCMZ4AurVIQLhC9ya
L5PpyNU2+gdkclXJcCVgjP9i1J9VEOhL8WdJs2IAGX71gvroTwmIl6z2afZ4lKOiZKDuOJa8Vi0B
sKK5AvReKJ5nnFpwSWREHh5ukzNCBNAmf6OZrsxUBRpzfXo2Edar1Xgchek2t2u+BYnm7xZQlQec
xxwmdxYUI/tXpMRxNOAoJfBkbMY4cTKMFK2XQepzS1PxXYX+oEdzKmxy8B/eqdmgm++s6//TGEJp
DQL6q+erw3AzFJSIvb7RE8Xe6xXTVNcOOMUVr2dzGjGWWcucHiW4cpvnJUuC6m3qs9RsQijf3GKg
OD6rNGKzdNhscGaRDxnUkrZepRCVlD9StPdFqiQbPcS6IQK1EjFbDypTP4CFqESZA52xR6JzQC07
+iW0EYRWRZmB+CGVCwplthPDeOU1/rA38MVjKtQfO137PuA3uZl5gjSTmfls2LhZJKWAhYTqerKq
/IrNfoDj2GN6rdv5Mu7ElwGGximoxfItAYloAQ1FY5aMaA71muJwrEXhzp/4kkBMAf9JvmCGhI4J
A5FObhR8ZVus8ZsybknAGMPlPHqt9gmNpUWJBeeGZ/f0zmYoqTOB7GB2S5RdQKKzyTOl3YGllRvJ
njhzmz8mgjFAB8upJI1fY2IH6y7SqtM5z56bh36u1QJFgWQtPj/v+ynsCMgUnrs0rgWl0IVyB9eo
OJqQHX9r+0Iy2SvB4Np8wk0E+RvIDxABysZ94RY6T5jRINZNI52QUNCkrhBZyTAmPx6EnD//lOLy
aN9hwXNfhSc/9A/DaFvqoHqOHGXPmTny9LoMRMdH44o4uKkxnnhtxNWSag1z1dhvHWGbM/PFXqHV
7+JA3G7RYvAw2tkuBUYEiYzDfWsw+D3BQ1NedXQCGTI9x6tTsV0Xequ5ON9Rwh6tQVF24DmjKuFP
yHDCecbb/zb7d0ep0DKRZLPQKYxdXc1qdVtVNckSS/7xrBU64wpPAz1tGN9ALBEGS3ILkKj9R+IR
ghGpZMwV8W5cfX7GEgtAj87WfDiix/dr8r9vY60zlyDdiCDjjf+2i31aT1JE3W8owleqcwP/9Htd
8+RqJJK6AmjSOLc+ic+FCfToM6nq64CPTKJ+iVSlSfMRKjyBwUIYjkef5hq8T+yOPnWWZOXXK5qN
uFyJvcoBOgjIDw3kmBUDHaxHojlv95sOT2cp7UYcgn3GoqDEnqQnHcG6CeSz2jZiR9RBt/J3Gc7d
cw3fChAVCU/hhl+TJMe1P+NfCNeFnSqoVN7XJetbtY/Fm8s2C+qEBIoyYIBIQzseN+tDZFZtwyrw
hRXwAfc/Q0sgj+TOC4JCas+VYcycMIN5O0e0mMu3sgCvAXgv2oODNJ7hlAJRf2nfhjRh6tucnCu0
0uiFlgNSvXRTDjvJssP2b3Pk0l9qa4TY2JaM5WSvyTobNt9VWP5ANdhxKcz57+FUW0p8GLDikpXg
I4Bsqd07AH6fDKTYkVQ92iIfxNGD+FrXoCIhTJ/CBAYT/SOCqlRmBkHiUk+Om53FHV3gc7/Ia/vX
ZxM9dOOxjndC5Tud80hNM9JpfGuI+bi0G0GLsO8L0vubO6fdp4a0HlkWwW8CB5o1iIg7z5vhJHdy
U06+WHXYXETcIis1of2j62ePNWe1LGIr0IFtyVAbipsAO410ksP73ppT60XtP9ab1vJGpxX/zQ8t
WeKTTjs8lqgeJDzYWeKQvnjYI1DyHXP/0TYf0pDbCTtYFHJBxljNFqNQmAojo9J2f1LTMgbcz+G1
4pF8fsw/tEo5uD3MS2CpG90iz6INzhds86i2Yq2E9z37sR1AXcapFeaczxc8J5cyUJfwikDqZvtr
BsEVZCZMFNlvYGdVnN7+VNB9LMXLo5Ae6rqHud3a07N8UbsLGMZmHZR6HIaPmuJ1WiohVnTvVwAD
Bqlx0w3408z1LX1fkRkN1ewAqpIRKayX3svFWN7qc3PMsTe+GahhW6SQa8jrMHSoMnjLm7uZgffa
DjxdZHRM7ta39trElvkYpuM8gW7uofKCNxMa0237qyUPVrDjLY8Cp6V6gmzAIrY9seiMUAzVs23H
ut3GENUdiMhQIuYU4jcGsvv4v35IjiDOtjov+W7YY3VTX+DqzQgdF6BBn4vWosLzNv+cfNkL8/qM
WWis88waInB35ViJTLt7qFQW+6wAiMmJF/oHxdp1goTGyrbL142ROxcpgljywxqahoNwCWFJpe68
1H99TS9CTF3Ph9jwONwdUS+eMyV2ecHV050tWscdIET8y8wUqoCrtVnmKQ7ukEyWtpHOQUDaiGy2
UI0J6e5heRLc6yUoSDIgGAlR4bDNIOxr+F82wSEjv82sgsmRqc3QrKfA1OIxROJTHTPnKIWO1lqU
UOvqVfFZyfisZU7iLVnAkPnMSy5zNg3VjeWvDcX7XeYcl+ih4nbSPxEuHqmzda5JPWXdMEQBZWi4
NOCfr2jak/mR33qm5xT34VeEHQZPwI0rA/NNIWsLH5PgtTJR3kd/kxx98NbjcFum8yQQqGmtLqID
HdnGjXKD5PU+xKT6+xHeBVuyV96jb3rXCklJgEfNviO5siSLcoTnsAwxFje2mrwRFIxu+ciFE6kO
BufB0zPUNv7a5gEKCJKn0nTxBH/Qdz2Ae5CmKFeiXLOEkDtCnv1UY5xSZwLUS1YRdQ0nOevMGCP+
Ckn50oTTwc+AlfLQ0v8xCilutsdwJDD4Bu4N6oVYmVLJFP/E+Hk0EL9+I4RM8oyZLzUPs9f38BNO
n/mnXJZVL48Zsgj+ElsDTzaOAZwjrIG2tRqyM7h42lIzF3nN9TsIz+ckZZYgGhjImQ1Lax29krqt
2gBcwRRynWvsb/SS+WvEsXCzLqh41+tSrhEt1/TBwnvR6Qyap943U9FB18z4GDBXh5f6bcaOmWXk
0pFtQ6+UxVAfcnJyks0o0LLg9XI+NqCqJlygBRF7kSevnw8oXo+yujBpVRZP7whxtTqatB0nojfc
2FIRwCiPXCBlksYjb/x/TVgOcdDs2YrrAw49IbrOFQVF5pXOTWYzg2k3scxT6vf0QEEOUTHr2H52
jZvwzka/nO53NEQmMc46h4qK+EGrRiKzjmWcl8XOP07XAsShsXJab2VYkc9VgcC5scCSdTIJEI4Q
UU5+282raAaf2WFoePvnDvM69eG50oCpBpGwiEKpbovW4C4bwUeVe6KJjRqJJMblC8JPUXcI3hLx
se8ZpeUyrIQ+9d0BtCvjihZ08hZ5QuuDM7tUKXV87tYp64Mx+TEqSLWPU22HM/NA2VNIdpC+h+0b
kmScrvO3FUN2DnCY4MoGc37OQpEI8A9PQyoTW7IorezYOEHxTnGhMmqa1cxTcxhJwOOxn/rmGyqx
IXx4j+EZFEMdQpjz14WeHIybqrWxELfjk5yHrVcZWlbWnhUtA9DjfpdfdpO0yXhmLLfSMRdnci9C
uT72C67BLqKJN3iPyrBeALqMyKkFj3l4tgtRy6MPo/lY3ij1dVlW6suHtDdez86kNCEJDps8cQZs
JK2JvcnTX4wbRMi+NMbqU4z/eLz/THoagF0wkoxh4X/ahx3QIi96a+DrqtBGJWcE8trZV3/3kEZf
I98jWHP3U9LyK4RtJoJhhfwEzb9Kd97ed0JW0sNnbVk1N3Naf46ZCCMU7Fhbumoq7jYlHMQGy/v0
uT1u9MoXvkLlsNoFSU/CjAb0lUTjyR6b07WJH6bPMkAvZwq2zL2NHEiA2tpFEFU2c1bICMyznbX4
qfNYz0sGDNcQ1IjKrT9tC076Kxal/vrRSRWSxKp3a0uzIB0EqI8vG/5j08KdnAYlSS5DkvzUmFY2
yueD9b/G40zGAVptekiSUwWd+44AOmo3FHCibcrJ0rnf3aTcgrpozGJwf7oKcmDqXORp7Lsx2owP
2+uosOkdQS73GlOOF4Q72Zx958FHBZOgOsHBh3O9aY6LaXph6aUjdssA1EUH2WEapBe+0lwXZeOS
cqdC8YLYcZ3lZaNWJv3WQ3A5QD9SZr+agRqg3b5CIr+6R5lToYlRgtsIvE/hv4c+BeNBjTZoA9oB
t1v/ifDgezRC2bQpBs/MjtBMQ9thH/AYRB+ZudJ5LOhOFUIuf16V+aVgEKEiH4ScMgo/kdRPe01Z
6RZIhzOtuId9VOJmXDOge4Bm2Oy+e3gn16VyGVcKK/J3sAJ43KURxxKyltfGXq3i8HUdILYFEGn7
0pNBY06GrNvu/Sza0SO86SWYaZLdvi6vbxnckwWmKfzxTXVYuhwCvHTzTHQ0vAMcLuY1nqGYGquc
4ZsqL/hRKPtNfdyDmw8NsIEJ0o/x0IVXgKDfmosSkCb0bPtOgENnbzBK4Hg7w/2RfM4blG+XuQ0u
d8716tAnss3DWXgCsxd+TwEQ33ZrxUK0uoMwyrTDnzKicZHq1rRUjcKDISNL9ZHejj7cYLvLw/6a
b5xYl/TIJtqG9fx2N8Xe1JASW0isAxjke1U7ucu9/OfyuM0tj4wzbUean9ksfmnYNPHtG109hvAC
A9kwMqDqSgkCiuKvwnNy89esD7LwOyNKBwmp64LFUSvmjJBf4dUz0wcMXXTH+8LDIJxC13r4SsOJ
YFXWD74KT4g3gmQFElyZnIdnEaew5xKfmRmFO3MO43XAcmvNR9d3B/GUHbBq5JoJkTqEGvgn3saN
5IyEUQ6X8waXd3igdx6jnhfxPz2xRXUHcTV/OPsP+1V54bFfWS495yvsLamNO2qBhi5N3EfazWfj
g7lDLkfLfA43J680M0frSt6f3PKdPMrcXhC8N+P4BG5hQ+JIrgXieSg2f8pyOMwnMqCFK5WZbxww
xMTmq+2HoiBx5tzsXZw3iWM6RzXS7Y+hNdhjtKQqg8B4hsnfVRkM5Ijc0P1/BRUfccvCtk0TkExl
A7zhQMuo6BVB/L3h4uVir/ONvh6Q/SuRyRs/tqwx71Z3zeuc2BuqrfitoSEUxquF4T+QYJ8/sRNh
3UDVmDM//dadm2/lz586NnK82nhbHB/v+VzSplYqsWFKAPdFGf3kEfceLdAOekamZ2hOmap8GQcc
A7B+jwfCYdNZVW4u7GN8jgc/SBG5yyH2nHdIgk4cATotdC70yc+wXesl1UnkFWSVeKdvtkd4PtE4
axtjuHLNCA7CBYk7xkyQzDAuWYdZkWoBL8JfnBre/p1chfH2wvfqgc1WcqZxpucEK6L4vGDY9+b2
IoWpIeeN+fMV4Qg97c0PvWqrPvFr+n1Lo6HD47HUe7jTL7tmos555iQ2Az/RatiEN5tr3dG3uKjO
NWIwDZaE3faMTAkTwj7J71wZreHxJknF9nZFmaLVeJKGmoL/gGs+aAHBpPfFm2yAab1wNM45bvm3
4Z0Nt3lGI5q8XKDlQt6LhHT+K7afbir/rMrV0c4I7vxqS9E/mnErCrHAZea475hl5WMP0S9aFezE
95hYKACepwWoI0HSHb7JzPW0muvfcNE6tf4qUlxlklPrALUc9isq7aITozVmphUqOrAK//jghtqv
d1GfMEj5bUu+nhLqSagQ8KWJFUBQTQi+h6YlvaNpKCIyw+3LuZx27WtuPsG4q0w1Ax5fuzwdW07u
6f19rmyUQ3Ye9JmQqAlPm+dyR7YXgUTNFtnzG8Y1wyIiv6tAfsPCW8ZJo8HYiUz0IxfuuZ7VjOae
lCjaxMz/C8OJ48r42i0QJY5smfon5RPw+6X6hhhlzbb5to/RFL2ipGwpLhirBlD0frjZnVGw6i57
5ZNmmSX4F/sAwUeDAmhVTjaGa8vZ6sXSWJJVZZlWlyacd7rz2FhVJyMadktDrd6Ix9/TeSbWGiiW
Azx6jUxLOXQJ45ned1A+G/69667CZh2p51cbPzLTJhCFGc/SxIzpHQ0b5cM6xlr3K7a4wl3zIS7C
VCR14Yem7q+ilkvGabHZ0jIcCafrLKOvuERt6TjkGk3Dta/wpGo+EqjVR/ATAyvV9nOhqsfsvOzz
S46zbSgTnUBDQCrThvoREnTrRwzfTRZYFKAyR/dj9GVoHM05x7xnhDhwV/JJafN4j3RxQJ6Z4kBa
L/et8dA36mNcIC8lM/uyQyq9AN9dH/e/2wTmIvo3Rc2pYdbdnXvHrFnlZKYNrP0e6U/OkB2oNlnX
AmfL+qRRmDVIzJc4hyoT1oOJAxfceECZ/4/Kim8O4AdawsOlp1mz52DW3l/r2y0aknU6PF0iAeh5
XzRsONW4qjZqO0l7j+634KcILKLQ1QDOZ5O7OAMPjJodkaguyfgciWIfFLIm/lx3Mi8gWbVdJ/5f
mBbJ8gaNHAIAHkHyLR+PqXoXctZ6eFA1cLWqnds4OiynnT7Ac9vGo/S/D3L90Y7VvWAUTXG8KJpw
lynj5jTZnB3nsURpVmrinoCuhbrSvA8XWBJuRyrBRudo9TkqAefq1IwGFIzPXesiiXxj3PHdxyBP
VIcgRvN7b7xO+cPscG3YLegJMObfLVGadv9WMa1UApgDkH3WxRCda5BnWh9lCDC+hoS4HgpVDlVq
2488t3x74QJGrr0UG9Ecgm63CPvAAqL2rGlzWf4QAXbywXSe8bhSANFXhFhjCxKC5DQM32Cw22za
rh5ti1FMWb0S2CMTa1tHMOuUuY74HmSSpdomD02M7hpeLuARCwySUQnOr4JF53jgM0BDWRLcLrtT
cuDqLolbhTe4zDAmVvIEEN/HCUsFD/nEZ4WZpZ/4oaoRtRbA9Wc2rmbCiYCREUZl4Xal87k7TCQ5
BQrB0FCry3NpBy5wjEIj25G7P4O37v5uEmLljmaNWX4sFrEi10BVWzgf5ueyQvpIenEgw3y5buST
jwqwPdphnq8/0XwDWwU4NcfI8ze1z9WsUxnOg9o+3y1TByuhLvvDD27LDQ9wtS/cYRJgFhOPP6/9
iktGAS+tUmTWeZwRo5z1kmxqdh04M2F+c5vF++ASRLKDGRBtFIBp8GbOgPyyPRi8ayGFZN9x8WLE
7W+qXyrtqay/ytAR7SSvSPtzTzXZMuYVGshYrBLCTID4aISCdqJgG1BADo7RB0fGyDV/VqL0/3qj
0pe5sMwLabLPhiI0OZXpFwweOXRA5IvMvm9is8HG+xPggZxfiCS4cKUQwhsrfz1xc4+Ylznktu3J
4nDGkupppwHdy2d3YicOE5b/VVGjIjze35eztPIgcMlpU2/783xvnq4tgBeXzcMR9I/fUsl0RrbB
PUZSujgIjxT2kaegNKqe/ST+QdRPH2a4+uU3rsnLjf150Jlv4Zqc3wy4ZYSEKyJ0KDJhgbTMidwu
sZIrAXt5ly8i86OQ+UHnEWlNE8eOLVB4ELDtX32i/1PM6lHlevgwCosGfBez8y2FplZfU45jDCRk
+EmFHAHbBxs+pxIJirxLeT0XggFDtNzL2EXzOfZMFf/9x5jj7WF49aEoxuoQjl5cmkcodY/8am+W
iM6QiNLOuiZVMpFIqh3EX1ZFGYcDbJkRbiaPClSHhumRvkjnGWmg8IuRbVYCghcMS1W42HAyCTWM
ufQkSee2+2ycrDdRjcQx/aEUQDGcALpIZv6o+NQFAt4WDRka7N5hJiN1aFOw2jGVHdWxzd56rYu6
CsQEgasNbJLNM7FQ9Olasic1KyyyXT/BzCt6UuwpJ5ravStIdsU37Lst3/ASixmfvNIcsOHZRg7F
UwAYxMHsVTOn2+YmaMEkboqaBd+ABrvNNT+KqCKzc1YTOpdUn8wK3yNnI9L/PVEj99uLzQMHwY9e
C6VYMCHKuYwLdoZJwjPwVnVph8sG6mS+ncuyYH08/3Wvt1tmiWFR9RjIMAmHVsokbv1Yk9lNiA4v
x6hO5aaDDpbrPitHXfb8Q+LZrJvxSdXa++vM4bHrUYmN3jd2Jy+uz/luFbqyOYLmASndNmUAZ6Fh
QJ1yigE3MsSKrzmHbVVqnr6XmE9/NI/Kd4fh/9RInPfirFLCXrips5s3nk3IPQ6ROASnQHUYxZBc
ZHyyQtxgYl6jXuwhnQQVvDK9ZfEzD0l921BMTkfh0Oyc/qdNPud2wGnyV12oOUJDD4Ak8LPxOeND
iFR4eqFlBUr7cpdFO3mmg+LC0AjtFfNLGoZbLslYsydINURNiJ+st5/l4XhsUTlU6y7En6SVo1C+
dRm4h1mT/OwFp6o+AFHQkhgVFme/WO2L5CKeT2VPx0jlQDZUerw1VlPhzGpspXThgV1NyFCOSLAp
RlZ3USWmLneX1+BiACMnzCTCxcMHd1xXDeONUNC9FlaS3e3u6OSg4VgEeFKqqP6dfDRyMs8ZZGJ4
jzP0Joa/wik9FtohYppYeCgAtQX4GAleo1HLYmFBauyuPU5RoGQozpp0YUNgjzW7ucUswQBWRX1H
JYb+/pF1fXv5YtOkGB2PwgQdacm1nZ7aPg8zVuzCUkG3AmEausWFjUOitgCekzZMjCpDk22CT76E
SjyPDWh9lnueg1eptxYFEv9aJC/FO90ODvDAl83Jt3XmQ8t6ZQlLvvzvJCwacRxusKBPpICTDGSl
cJyl+2CztVYmLXtuy1lD46BCziJYWKcbps3XBWCfve8uqKBfGdAZnm/z8rcN47k4s+Wozlu0ExHI
Rx8pjU+EttL1huYkNuINTxjz1rHfJPQlHv73p3eI2dCEWFWSURbaVhBQKOmLY4/unTagxE4yzDDP
H43dlAu0wfY4LFvtlkXI9zid93Q3YSFB2j8ZJdIDU7EzI8CQbHmu8cCTuLxz/IphgYNkkW3G8JwK
3q4X4YodtpglHaNcs0QbuncIl9i8G5I0TUHpDgN0INcIqByr8IrgsV/L60oESDRh202g/zBGg2D/
kb7v+PYl7HyVEcaPRUvh7WsY5CxtZl1Jpue3hjIerl+ViGJXdWz6mu88rKtSDb1P4hV/MSMt0UXz
YTiByiHVoSX/CJyESMcVA+N4Qap+SfXYikNyAnENd/5Xn0PkK2IG4fL5IPi6WEsny9D7Qn0l+iTO
+ZXMRPTympoQaPN8RFXgfNQCaO89rn+/lv3zqp6SLOOiR2Ihh8UowY6suIOBHnDUoc47gB3aoJ24
JRxe9hNisvVbaNjPUhbADiR6bS0Jdin0jI50BVPT9J3S1eNqbTepH50l04RRKNNFR5oOtxvyisob
3tiaFElwzc3RWYlsaXqRQBbPBe7XNpCgxC2kesT5mIXOube3LgGgcRMGqqfnFrAyq3NaZ0reALNL
usYTtiU+/dskRVWRMG5+BZ69VICv+MXQmj9Wt69Dl2jey5iTTPO6tgTrY1IUCy9IaESxEolpRdDn
NeY8M0GhfuF0/u5efvhCLSQ2YdPNWnrArlvLG9zaDLjFbB4s19X/YOxQ6pYpgvO+NphbEZPk1QG3
5SKReo+uQGNbRKza7wRaLIfLzwBvv2hrgSjc/g8jfz0tqpI9boR3jeX2OSbQsqgLMGB8lzC5JKC4
ziHg5T6IVsZkDY4UgR9Exh5a1b/J5kxGJrRD15gvPSvto0AKweFv3wx5k4oJMXLy9HQcI7ZjyFtk
U678fcWQ5wcGxYMwSoV3tLaFVctbxAbNV7LS5BdPtVJ9kt10K4fIZf9KvSPmfZSZ/4O9Iblmr429
8Bx6XP7KItRcWmpU0gvxMHURwIDyo3YlUWr5kvbod6Vp8Phq7K8Gu8A5x5piu9BYh8BpouK/W+zB
H0hwxU5c+oXF16eu64L13RUaxTxuiUcMLnMlbH40PGUEKe4IF6hJ9ycKHmJCgRpIH0hqG9EbqgaS
9CLHByVwbsD1yOPksS58VUC9MKw4uodzO/vGJMGNapZxie/vmUFFP4BN46tkXgaroWXUIwE+r6zL
Uoz5r82UUmlI0wtZlGR/6cs1/8BGr6mWgkTwU8NhmB1dBhAkJt+6rZI/BmIUfR6ZBcKx3fSGzOz6
WjeIgy4Ap+csgu0pd2xxD2Wqb7ZQm4Ec45Q4wEgZZIi9QeaNSmwRoqX7noQ+EhUotTEL1hqen6WM
FC00/bRxzJ/Pq55Kolecyq0nhEfNZ2KWzn618XiD6VzapDmnZ5FXvKLbq300mLw6beG/RfqLsCAs
B1TGjHp3i2RU1PSQDWVU0g62Fv48l2KNYqZ72F+lyt3+mI1YxsmndBy+Wb06yWSH4B4Jt93B5zGP
hym6KZZ+9ukCialN6482BtLqJf0GQvK4k6jf5fz/l+FxQuPBalRXfw7kd7N0JNOcIsvCxa6Ngqbo
1jh5s2HGeUwj9l5b0nGtDACvEt6h7My/O5y0lHj96a1bptSY9iZpJSW70ZvdP7rFBB+DqQi4RB95
YbQrQuI2AN/2kqySBWwMy/x+HZcoOVj710PTW7qbqbBMl5v5+LFVT0Pjbn/nP6/O9uHRE1PBGu7N
zsgLrnwQIzU7hG9gwDjB2g1ScNbY/JKq6+tPuX394lYtYlfuXC3Ft93GvSrhOQZrMOYqby8UiWA/
8vRF2IirTvaqwzi/XPsfNIbnfgX/9SuaSxU14MD+bZnX2AQxrbBiYbY42zCCr29+EtNP6l5kxRRc
73UrKLC7++BIESXWWC2OqvC7ogyKv6j6c+7uk+TO1D5stDZhYbCisAOo1zB3AxN4czPTVvh5o4k7
ds1xRjhPKt5nFFxX5JCJHLVUW7qeARB/uTvthvQln7ZECXe+m15O8QU2yy/T+N/EeVIyMK9JrpwL
YWKW/Ue+roUIZmK+05ZOf/ysrwgMsyOrjT2EiACfUR5XcBrn9oeAso8qgXnO6Lw/EGhTIjR/6Zw9
s2/0x4FPsTDXwc8+y0iv/+vaslEeFRUatRs8h/Hge2tWLldKCWLWKwKUd3pV3dE79Y0XOC1FJdGO
6pVj0DdaFVvXSGIba/BiKmTG4W4j6IMkwLaTumaBoj5i26zcPDG3jVkoPZATlSX6BgabZwzEI3GA
aouLm3gKRkuFMneQcA2uIKwWCjshP3ToXWB6/rcZWteYrKP0j89dOSn4H3ycJFRqGaUBYOTLyeOA
D2rG2ESnpnWO+kRclPLgjrko2XOO1Pw3IriFxZ8SmfswOggeV3ZIBgNyLLYd/8rX9Cxze17FaUtZ
HY3YVdFfjNZdyRScrmTeDDMhja2KUj4CnRwL4ZBBkjWDFTIrhxnZK01WZaWMG7T6UE9RsGeXkr8G
2sZb3yoSMad1NEnFYnZ52qk8P1mZVVTkoINem1ArD9x2Lgz3YWpfmnEvpRkFeswGX2gjgVS+LUNV
pcvqyFcn9yFlVNrGQ7FEvusx/Cx7As5vUmC93U7W9RAnglk6kJL0HH9RqJ0kxrNMr+i+OG4n5eYz
AklnO1Z7aWV4HitKH+gYx8RF9lLDhgjEreq/mDC7Ui7Qup1h21AGzI4M3+MMKG9AAWmT0tdL32C6
TRxorJkUODUv5csdNQ1H5k2m7GjQAnJXZmIEr2UrhXr3HKDexo+d9Y80ti1/qVQEzjnZ3lZNQy3w
7tuuX7wz3u6V31qcSSeACKTQ8LgKN70sksv5BVMWqjPY3buy14sFpMZC7rEHXDSv5Ozd1Do+cyTe
fQFhPA9B1tiPGKpsjqtJuGYebnZvU4PaAUvumRpsScne/NvrwrzWOCn8JmOsa+XFtILXgXAvclJV
30a6nqGE9v93mm52ehIkzjMUIrALfYXhY7nIpajLLvltSg/T9qUmQFJkI81Ksgdj8PqJpXTfFCEU
aMlGSl2XItqN0q0WY0u2QVVHRmB80i6fSfBUiVjw3yol9dmUtMhU+mLYj8T9wJXleanvi2zssQJW
zyfWFazRN/03iNYhTNJ2E3BkZsMaP8317UTyMY9X55wCYVj6MAz7QY1WvwDPyQQp67jfuFuL+K+N
giOFJzHmR90T1HzpwnP7lql2HgqBNp90515Hd7alkPKVCk1DVVnLtRihLq7fegHiecyMqv58kW7g
oEYNNine8FaocqhSADQVBDpbIHIaH6HqY57wrbUuUc2RZIMosAP6GlsWMgiRbcspyrvHhhEnPQ38
AzlBSNDbE+eKgQ2YcdluF8D49fH4yCUryvf9Futzcd/ldmHZfsgJFbw+T6eaO7MROMruz6AOtj1K
AqNTr6oy1GoPv7/bShefyU5ATMujx+Fh5I3kbRodVO7ZSJfmfS7UlL6AzdV6EarO8Zwb/L3/kMQI
hZboyNNKxXimudi4lqgTaMmmGfiXJZsU3YNtdFFOl+MUV9bTGXRbZ/2wBTd9emyF5ebRbVOtiwXq
gpbm9/5v7g3ZiLVzsMuPpQFrWl+prxWWtfdGouzERf6iquPegrRXK8zFqRUn/WGS2DIPx8mdQsY0
CdIouwcFowDCmmLwmEvSgXYQ79R77OTWIAM7OeGhPqZ2IavRsKY2bdUGnxXEEbqM7J7WftqEGikI
CUnjot6/Um4mCMFbLSPjKNmQlvN36YmphihxJrbDkFrxtIRc6ttXDDCa/WOHzopjZNojzjAOu0SK
AlP8jkvwenWhazFdwRy5ItQ7h3HrVILuWafjw5+jFQW30GFciemXo2Cct5tWGimk0htKHSRz7a+1
rjr2/kMBww/owiFElV4iRBB0kQFFh/X0B1Wov37V9lUXVcl4/KdDyLcf0/f6RcA7yaWk2e4M/mJy
7zfii66Czq+H57/W6peK3WvdwQ22qffpSyDDMw8U/CulhUesGubeuF1O1mdpfzYXq3rYo8jKCH1u
l6xij82KKj/y3YbAhuDh+32soQgeRJ9wfqoJQ17o1XmrXVmE1R9mrTl2oD+KgFr82QGYwkPB9mpL
9LCzIYWtZJbIttCPjHjZjNDcpOGDII68wEaE7iilLyzGyqYhhd55utJeZq79ojg+cj+XQHE2uu+z
LDVwGlpWSBaHaC9xHI+2Up6CPCVEsF7sYaAhiJlBBMZr2ovLF9duMqrTZfqJwdMjevIRI8aJ2yIG
DO70fXLtQ2N5DTamYsOnC80Aw4NBMzhTmysex+rN1dggwbPSAKZNKpmYUOTOXJ7eFPFa6Suyuxb1
lJI/ifejOsikOd2gJzKGjR9bl0JHTB1aoD2wziI9Va6FIrtytP1QWQMDU45Alfeo4rZBiVpizwNg
1dCj/njfE7wM/Q0JyWzYtkWoLTO3IeuzILBRo4SAMKAL3QotCOHMO8x9bR+iNJqb5QoQTZcjqVxG
xDRBFfvqD1QwIGPcYQklhH2TfHgPV9un4qjghxtEChMI8dI0zsw3n7xSttJ4a5L9WUD2UdYmKYgW
AbKrDX2i9h7I69ru4QsRpAwfHhKEbKPuE+hanRMxLyN4416mXKWv81D4xXtk91YSBZGuZv2izqgT
xy1LgikH/7RkvzeMr4LD/VAz4yRYAgxUBLAOY1vCSosHNZNCKKvvKEJ4NqOMImQxp5fjtBgo70n9
15JCbWLyh6N/7jXaKAYS37Pz+yn3+upjuipHwHPnK3zt3g6bfAVnzqdZhrnYgt1r2905F6BsbSVV
GL2OgO9U7kxizRpBqxT+OcXZVG+NCEZg+080gNV0c2n+f3IIA/OU0vsUcSkDaSq9Ajs7g5bwVxv3
E+8FE0EcVAaxQmFx3vqSJ8vcyiv0YMulpuPVK69SW1jmCB+L4/KYhTg3RuOrdAkLoJMcEHmCQocv
Un++Ma5J/J9qYvJnPd3O+s9rmpQa8PdNXeh+gdtydG18ZZ4md7U2vNdhb2CHgQW8r8IZmAGtCRVS
SQ/w2ZxE9HRic+/88q6XHavqaFZHHSjFDua9MadScUql2Qq6FbwT+/dVVT5o9K5ckt++rjpJn3x/
SnirkFPHeGDYL6J1Cj0JfPZM9B65RBLI6/5nlivGJ6LUQbgoNrSNEW05p677QxAbsxhCHJsU05AQ
t2xMkXA3JnKqTBXEqGElf11kAAm5/rQlu0Uuu6ZcSCVSJsEcNdVvzClDNbUDmPArOLvLPxJlWZpA
yHUExj7HrqT9UCfoQ8FP65QcDtuFEMkMO1xSO5VlkCMotDnNcQnvXtgiFYbqsEGhdf1IuYjSSPpO
nsJ2UoLoql5VjPIZJJfZelJCREaNTC23BSO/JkjdiXiLPZ9U1aOpAfXPwnfENO5M02EmVl1b08gr
arUZG4BC2bTZPcTDR7T/6WqWBXXf4EdtVv5Ml5WDO/UXXrsTCY9mA9M3RJudTBwGtCypaJ3igsgm
mQmIPyhj+VxEjDpNLqiw5GKsaUCgoEAOgCAh+2Cnb+Wspyt3YcaHef2G2N4/tfiGDy4YlKQgYJN8
TsnproDs3xim23by57PzszJuKWO2Io2z0tSsu2h128o7Rey89f6oepBN+KzYhThb64HK55y9SzJe
0fXQBVsUUZFQbEKEIV+HHW9gy6GURhP/JgYOJnp0J792BW/fYAW9eSle9pquumt4oMPMpkEBP/n3
4WdL3+QgNxLXsyaFwKCF10vqiGWrVds+iberhmkK87rcGzJrDg9JcEg51Ua0xD/+P8KbVFuJ5UHC
fQ6fxTjr8S68SoYom0vdBrY+kiVnnor8uGMw640Xo5b99uBnxSAkUTx0J/MpvnWR6kQgAKP97VSH
R+rPWjeKDWLXOIMwCWpjJqY7YPEmwAzdZbykZbrDf/D2csX2LeP0eGj54EdSr4vvPAOTYGrT94zS
JUa0p+HYzthI3R4lBFsJBRAsBaP9eahhZx1HGsT+9EQI1w6cWJ0XiSCEXSH4LVovC0TGxNAebr+d
fqFCgL50773SICKjmJniwA+4K+zA/euT6EXz3TIFLaJSo+mcnJGeEyRf0q5VvGASrdKJnsqLLgKc
wBC7bZdOQ7yGHJ/pLDeFnuqzZwMIiIKmeN/AcrrY4ChqXv6SjmSEAAeSnUMxAZNUvJop7ZEmxrlO
iSmNRIzeCNxA8aDeeDDlYmcgEwrG5+QtHW2n9I7B/RnCZVY8025ZBvaR0c3fEiwCyCNI1eEkF3zj
J1nhxdviZ6b7buBWWM5cWwLxR8PY/CIK/OPsfcHWcfBKY89lxErU4keVHKxolfwxCt8AfhfjLqQP
58zwnfkgK4yAl0sLdvyt7rUoFv98rEjsx4zaXkWHSJO9A/fRrpfouFkxUMDNy9uZdl3WARmpQrY8
eFG1nkNYhKOqZuzdZR4wcO88nK09+oFotdZP28HdduOV1452udnWVr0EfdWgEi5Li4mkHY7JENLh
lI0wzbwwpAZCUEab1scQ3tpPmueeEk5HMXqEaqg9zfudu5AectfYUWKWeNjDf/JyzeIMcpuBFgCf
fEaslClTl5IAUU+3F6aUt9XxkkpMUhEwEv6lE5D0+YVAozpLB77/KthmyFS0sIBoyC7LGi0N3H8x
bSITXT2OBUNbow6huZpLLLwC+UWP8sjBvJQ98/+fZfliWkaEC/IRaA40FWVIe9Fd/QpPd0wMjiYg
8Iz2WWdMwbLRTBphEaIuOvWI8VsqVV7CSOskacJrCS+ZI8vZmKSEP6HcM+WAoJJmT8luQzYBFHMM
hmFrm/lVh/bd85ziFgMKoqYnSdfpa7of9Y8uvcKuXsDBxX4gJbLZGcZEE5+hS3yJJgsHgiwCRTP9
+bXYampcrDZ4AOWaAmHhuwYfbcCw2XEk2FTUz7ZzZsXxcc+k/i0UVPvJ8xsrguyCY3LXe0sueYl8
jI9YLWCSinrU3mliOCUWFXla7G7I0l9bnq8gllvRA4Xcy8gF2eW2ue8eoqBxYl51zdaRR2dBzi/h
2+j0gykAOtIQdug7FA3uWrWrlS59WvLqKheQmnizeTMK46xf2H3F1/dd6ITkywhNATDVjLYVoKJh
+zFu5BXfDE85LT+A2zgGUWRn1hgYipF/dn7UJASZhZN2yur7v32hvVppOPHmRXdG4tlD9jkugRuj
czIj8v4MzvHd7ZkNwvQ1dwombHzhfZGOiV4rEFh6OUcvMWMAPVFtgYKeynzLPAxjbO0BswvSRtCO
dpeRbUn3+A6m+oUBEOzdEqYDhGnD73Q43U0MCi0w+vGyyUQMYtO1o2y+NFM9zC+NIALKlVC8/59i
+6bOm3OFSYvxkotlXyLGXX1r1u7kxQmQOsoc2HCD1Sliqmd31tG01IL69LTszaGvay7NnFMUClAY
IAD8gKCvet9wGoDo1UVsAVl8eaPLb34iHvmTcE+aRwHaCYhob1BeiM2TfFIvupeM1sPAgct737I4
2yZruN/X121B9r5mCUZ7pJAaCcmiAzmCEd3w/fiUxQLRdhI8RnCs5M86msMJK3nNJZcscwWzqVWh
+5znthMCUo3Jc3aTZW6J3uUK5tl22YVfg/bagN8d04Vt3zURT2rFcp0XoDwdBtR+Af9lHM4WmfBF
BpnvC0FJyu2zvhe0zzWv1/Gfe2RP2cwcf0F4EAVEfM9bQPtZjPyII6hepbs31cpnUrjxopaNUesb
kJs6TLsj/yhc6xnQmC+VvozgJ9LmJf5KFxoluuJst/lh9R/wOg7Zef8aAfDcq0XRPzV7MMLh/FCp
lHNAUaMbKuHAyKuLiD+8UB0pc53b6TQrquu+UjNKNhKq9eHj5AErCMK7KNzjD14pKrQSF1JK4haF
xE5gSgVoTVHvcJEUcCVF4+sRMd3emrzMxBtxYzN6XlsJ/+j6i14eAt3BFlxb0GIpkR4DwIyyWA5o
BZQwEqETjl3GZZ4o4qZI6Fnq0uK4Wm8ZgV+kEIuGWVx5F4uG++WX8YGuoEUupG89/2b36i+v7Hj3
fy58jodZmAj6eBCeG4IE+Y6F1XqKav5/IdsOH+gcaf4cMhkRX+VIASfkGe9cua6NpCfXAn/RuAVw
pcmKglBYryAA4RGh7+uIoRgJJ/hSDGA+hOF6mD7bFf19A+Gx166XVYVnFco2LYBaMlx6IhA1JYz7
Zo4b8cnZjrBb+lJV7vSTyI3ag+Z4uzEOmJOhTWK1KijlsvNNnepvnzBh12ssQnN4MFiW19HGPtJP
35Z8JJDdQ5tgP5MwPqTmYNE+AOnxPrXgfli8lYpzA5JlmmhDz/DV1Rx8mYBLElJjL3MRyrXZb/1w
B8NzSzAp06rM/sgUGQeMuW5mgy0/oRrKKOYRCWMHxbs3vCK5o7O7yai5prbHh14RNqfOKZFSlSca
1Rq47c2V7oc0rQiyOVlI4IlBLGreRVCqobxK0g1Su+fM/OvwMv7GMBHik/nJzhAOjLecom+x20+N
jtDDHQvjIHdgXfSmoMjs5FHLPMBzAkJysWfRTIKQNUbVKRe7LkMijcJzfCn1blNuqXbAqpGzTD+4
9KPMlTfZsLkJ31pAAITiX96cjQZ2eU4YxHJbHAM5q3C/pmMLYFfxs4JzNSM4kN2ss/Uv2PA00K+R
Rb7Uk+IiGu9zCV4KUXFVG69TAxk6k+3Qm8ku1ePhprs6g/TG1lAVCSUFFfHCTugP3c+S5s8KbD3t
UPAUQQ5+b5xk2xHXMrjvW/UrKYGLzHRX0y1qEtZA90snC5pgowXKw6HP8zUZOpxfByWcbcQkefIS
ba7V+DHnOISmi5McrbcY4c5xkCf4uTrL/IGr+amb2RkL9mF1+XWIm8d2e5TMVL7tUWIwxr5f8etS
soE4rDnCzAnPmRHfFtAfEQRliypJYJCMGQqGp+tQRbJNXRwX+PaPw7XEvo2eqICV2+2wBvGLUfFn
r46u8dU0ewp9R6boSLAcdjNqjN6xzJAQCX/R5MFLipZBAywjh7m9OnW6NxuoabQYKilmw4sWiBQ/
WR2RcaKAR6q8YrpvBKHCy7iq14C37Trj+UoT3zXP+zRIX+4t9LEtZ3+aoQ5trz0Ayn0jKUiFOztf
cU/ZYOSlG35NmrHUvNbNaQr1JmJ2Qt7b/JWpJS3m8CwepThwz5tgV/WoO83Vl2IRgLmDHLIbNUv4
DER3mnlXaErwoAXbKcmfdqixgiNuXfHAIKMR8vM5w3Si4LG+ws8PWikNdmd+HMenlz1Ime1+Mcod
hoYRPXCNCg3RM/Pdux0uyn1QW5zHKGulL7r8+pmzdFH4wKZuVGnIgxxgyAlkaaC8x7TSabdR39Ia
rGl3W/sVDH6jlPvvE8aCVYLgi9zXqxih7TgRA3w/WzUYIz3eIsMs43oNHRsc2GQI72iFxi4wZuKQ
BYBu41QEnTYmPJcDgjjGTDufDjoa1UzqqgSDbcmUQ8fZiLalC7BSOLMxi5uJj1oyYeUDjQNT7Xyf
+CuPa8UV3bwMGw3Z0UEaQ4wphQo7/L5T80L9aOZvYxD/j/gtUrgA+hBjkro9/bZ/x6kivXSRnXDI
Mbo3M3/mxKcqo19r0ytJr63u/qFAPzF00Ig4/Zfq/ffO4qWd8MJv9HSZEsOaz7XpbDcOA9g9aN6s
wmGS2+yJ57mhOaXKTu1Uu2AZElrJjcfpjeVinrXStu6vDrEuPrtwVeJ3fRqmahpjTeiyQ6D/DMHX
yzM7M29a26qOEPLE4dvl4x9gxf9Pzl4oekEatxY9K2IQpAb2C69iHA3scFi02hM7bywSNVW6ANrO
NlCgbYdgnMNRNLviHtYL0ChLNZNhvsGKnyphiXo6V1w7mDd4KCZC+gk36/GTd2FWUSYdifWSkRHG
+4aaJxvmVolMc8Rjf7Iy4hm1rUMXjfZetnQ22peTFoOQ2eLI887DjpwyG1sM+XVYlbp3iyULtuqI
oJfQnM7JnbpdAuUzJyV4zkLHOUpWyVe1OuNY9oXk/R1WomkwWBTq12aV3TMxeZCI01cIP/kniV8E
dRUe8cDILmhBHQnaFcT/zE9BybRfGigf2cZKz0IQ3i3qU0mnWQc6THgR0fvWK8aA84N4bIgOugyR
QNtjp89cdGFiQLngMTWMbztrSchMXfy8ZUCRrB3iIq9k9GI/CFafqxp9zoZdAKY7irN4wrOIQZt5
46Kt1TXXkEawiM19FTmy+AE/k8KNeMPzxbUS22dinh0IXSVmeNPw5FwWa8qBxl7i+KfqfwWuMY7G
90ZdH3rgH82lgVeZHq7KpiY9tMqxqV8GjqW1Tw5MLpMTPg/Bkup1dUAQ5hP2nBXWU15r/L3eceW8
EggA6AC7Z0uNN5wgTEmeKmSrQP56tf5PPrlbzhXiClb4RqTNnmhYAhpWqC00efpB/YjKc3/TgjFU
esx5ra1/2cQz/GiJT2pYtkuOV/cIJ8NR31C+X+9BSiVASfT7XII4NctoSAHjTAf26sKNlZI5Np5M
6ZQ1y5Sg82ooHNJdYKOGEQTbHCmU3mEAQFamvG2A0bX0dTLB38YTZ5hozBxu3bjBUoVbsgOlVw/e
RquFfkFeBm+Q7FOSFEcUXYNTuiyyqQB9hqSRAchaRZsKPVDfwgf9+eOPjH/163Tly7baTcdy6nnu
JBWgTrOJlGld7eVyhYMU76lbXKx9L/nFu6LYCVbcyNY0hGlDAwZPBy6YwX2UXIhApY0oTZ5LbGdm
CiES14JWhrGF3Bd37hCDLbLcQB7Nl/zzTXf8kCZ6wiBwOb4Y3LuDe/Vtuu2V+KZ3ju3x9X3XC5YR
FfULP/3Wcp7bHq3BZztnMlhRJzKJxkE7WjfnLv+hNnk2UyCKpEIsNEvhoTiTiLhtgzCXEz7nMy/Q
/VAlf7IUInIChgcrZlhsQcPhlXvgWWwbsq2ZBMCxGjKWk8Sd+fwmO49PrdK8hFgG2ulz5/kVS+P9
guuD033RAQT5tkQ/rXXNnmbXp1dIn4DgHXklBrKVDbVNCcxtnBiulZvT2x1G/Lw/tyRtseBEXLE+
Ze8i8hDu3TFd6LCPE/N3xjBCk+8GoTGbUFUTBv2u7swo1kg2Z9wV+G/OA1hPoBLxcmbng/fCaumd
sOAEM5B4KXFkfdJEm7zfJeP+h3eXMwuWOhjhrPO+24lzvMO6vcKEu+U1KluJqYSfksXqRppNzOXF
awxInQLCWF0n5F2n3yyOrFGwA6v7iwJwhZKQY8bGD2xj4JCmfzC8xvVbESbav2hvf1hHlcPYFjIO
g79gyMpIiVN5RyMHmkrTKl2ZXFKTU1q/My5gL9JGyhqSH+y5V8N7xut00gwY8EsYNpxzM9ZsReXC
hitWIPIbdf26g58hF4DJeII9xLQFtpNbi4gy4xt+y0rUyIC87M4qrzZTFF4preoeIwN4PUTzkdwl
t3e65oOp/SAQPxPD5spxz86lNs/fJhWVepNvjSeMbkBy9WXiFvydBRfGiB14AxE/m470toNsINA3
lE6/UmTyJN1/Qr79HTcmTrNp+30SvIQaxQ9HJYz/E5R3pSW4EhWrOoTymn2hxXABky9pemx0f+W0
AvIbT9GG8io2baXXJYtbiK37b7JHqVL9Eazel0P8AVcIvX4ureTkfNnSJuqjfkHZFPY21hganI+X
IL95oJ1tlaTwsS3JV4pJBI49WgD7r7BB1GXRPo5NN1zkFDeYFLF+KO23ot8ih6+2BlO4WWRDwX9M
UDG1ZBfd35ePQn9+YI7rQVm/QaTMiJD5h2TdCM47SIKKHCbkcE0uBkYRppbEW8AXHCM/YXppBrN/
l7ZsWwaXHt2JGAMvIctNvMQGe2WnrjPhh0Zd+syWVNwVBsXpXQTXTN4iI29UOboWNhqzoZQzsu1I
oMrDXamjBT5OzRC+7PKsmi8+STFk2HNTTKwOlqeWXFIHn5EVm+1lmLCM695IC87OM+OeN6Ecfkra
SNruJ8mt0oVH+z3AZAhzGsk40rDWS8AcUekL94kuhDk1eRVVImPmsE76SersczOkhdB7zjVqMQg5
d3M4MS2dm2MkZ7aYz0SXCfyGXLCaJ/hcVJR0icywz/lnfqxzBi0iFf+MmE1CQHkdAAiskcMq8ofk
hwHjs785ezfQOZBeIOR5pfLwP7K/m7wbfASXd7qMCM4284pAiQgVmJfo36j5Y9dUfyIeUA2pTLaD
068WuLSmfZsazCDu1S+xUNee2tCV9d2a1Ff98JiSuNvOQzhv3iibSNXEdnr+IGOqyBCGKQNdVKi6
QgMbVwWuKC4M+G+SWhqh57x3cX8C1pOS8P+IQK9QjcIm7qaAvaFa5gRC+LyFHZiFCgK5gxW8y9gM
B8xiFtFrHqantO0aEwSFCm8urK2B/VwNSCLsvyB+RdGfbrMSFDQuFdW/FV4956f8Edql2OZCdtM/
2qWBID2VxC1Yjv07ak3W7Y7UsLIyYugc89Ru9SWgbVgVeGgFG/rN8ZJpuo2tvvbPcUWM8lTFsvSd
eY/2iPGVW5RCRa8kcfzw2uK74VWazzq0YyIgGtwJeR1BGOMXkQ3p4DN4JyH2CI3eta5slvhhxjE3
cK0aD9w3ypHkoImq+S7OhRXuA7cFedC1x0rppjTC1/b5NzzlxjHE4P8wATtnL3wiL2eKFHlh31Qf
5Sxgmh17vo9X9EneNUxrekIW/cruR3krvIw7uLNxvhBWkxXly/VMRNTDessakdJoisdgLoXHnysV
N2u2Pvi3HFg+phSIZxelxjZ9ok923CKMd8OD4fn2/uFtBlFipv0O1rQieIP/FgZVI7TKR7W4UJdp
N7WXM74AB+qBwTvrVdnN5HEBMAglYriPVLd9U7I7GNfMI8dOKXVn/sCutmXauuk9NphsmcS6lHOg
dKKP6cIyQ3a0NhSzIpkEPQ8u6JT946rYAsfjnYWsop9fmZs+JClA7ZZ+qocOh2SruSrNNgIdlBiv
uuYwZmnuO9iHcIqxP5dDU8fNvOHHmboapO2/VVplA6NudOIOxhhCh0Z9aR/osGdbtshI5x3zu5h5
mMnyhwO9mVxzY3k8InipMpln4UNdLKd+vyX8ZcBEJdigQwKkrnlyPfvT3MVC+uhRnqdrXeO9nYAt
RWFg0N4o33wm4EJcQaeqva/0ZAmHzni60cYf3W4AzoPsSSxVNdAWI5AyiXWty6kLkSt3qpUBKImq
Oc6rfLunzCe4BNJSfeACdzHIz7EB8IqufpHwP75dqwPITh/ok/U38anoTKrOnQH97XyiG45yMGy0
l2c8HJLNRvET7uZGd/QwjSMIdX3WAVeDYCf4hCml/oWXBjNylSzQoO3tqvmq4MlFWIC5MSk0QT5d
w8KXH/N1tatfdA+FK+AFzPY1DCaHeNFBi/duNO7AgKrGSI8QoREQpaKnoaVdcrRdN2/ef7YQlqw+
NATqmZ76Ba/ED8bsJgUKNBE6Ufw3eIGMRa9TJrpNT6sfXBZ159P4RAgy7Hwx0laz21OZyoYL8+gy
umqJwFVdby1/vFWfe0gE1AeS0UFRaSiD6X/HTQsUYjgS5gLxvoXnNmG7mfcCUeaOx6wYeCCaagxz
/V1sUHksAXqGN2bGORbwtdlH436DsTm+479B5r/tWPC2GoH1DFviYXa/fkki2llB+Lqd2qPfWUWo
JiLn/sV+rnQoy1qbyQe8bfqjutZ4GxPo0kpARP3scpGDoWtozRWIpWf8jGmO2pII298tcCuqcutU
5XOlhbhpx8XOVwuZh0SD9BzorvapSE+UG95T6eCZv6eXYoUQti9y7Ad/J6/PH1r+6xwrGRahpD7q
cS664DKJ4+/sErkwxQR4ws0NqBPhl03nIbeVaHj287bp7cr9L0AdfLfehg9BcEwvfot9+bfSF8Z4
r6tXDLOwCxV4tfGawP91mVieB/RI3m3HnVQ2LqeJTQL9TKcIeWh6tjUNnJFzMlUJCU94Pw6gTOur
BSSsqmy4sYsZcL3lTQfudpziyoNZW2rcyQ/IbnutyLmoG0T2LUBfUbedYS/LOnZEztLU3qKazxA+
eFA/wNsB5an0tn6IzsdQqEOl0KJh/JvXSvDGI5kmVYVzwEdYLFg8Z2t4yos1wlj8vbRR+jagrFSO
bjO5FFY0UDd7g/P3TluN5Xh21Z2TtpoQEsQIyOW3N5wf3fv9W89gco4pAkbPhTiGY7nVmrSnO+7Z
koRFHa6WkONZKSXcNuiaWYzeyg9R8580f6XVmiivHIV+eZqTJAvSbesby3LImqgBA9Fa5i/i0xUq
UGuBFlrLSWy9tOG+fnVzrOH+GwrctJuUhMLwNZsUrdMziNAgKH3Q9pZWD2yHt4njKEeExcRzZPDm
NfJLvaZw68PjRM18HpXsoHEgFtUwlD8xGvcGb4BXylS1V+mUPasUL3p69CVpeeTsCJf13DIYV909
2gTpWjESLgXOOb/dZiP7QZRRLHh+4M10+mtm7u4sEGaNaowx03AVdRLIASRir4CH2M119uiwvPM4
Ai+A/1MrCXWjxADMP/X3VH2a8cC8DJEQZx12NIqjNqNYSZ6Dp0lqa8KSJz8QuTPYw9FUvfk2gEze
+mOaCtemCdkrI5CxAqRq20m/Z2CYxbNCkrOW0WqfxTNgxQioSZBWyNOS6WEwLVbsXipIHZzlVFtq
Kt/0nIrHiBazhex23RUueiCWUqdyk6TAOV4+c+miuQ1ep/V7gV96Q1XrjWb0CQG4iq4Cnd/Tq30+
4tg6tJuDRUo1sJSa4kWBErBL9nOwkF/2OFKK0Miukbg3PP1xokE2o3gKmdwinfp7tN4eAkodNqKW
o9R+GSiQneZXSgDZqNMUGRuKurhe7n7EywmJ1JInxZ2u1ZcUIMyahczp69cbPN4w2pnNOBFZo/CP
JnQ1ZRyXV2pwbqlRytJCKZzrRI7xBSCReFtqDO7H3WtPDbNmjTHXu0COGB0zq2SnhJXKFOVF8R38
t0Eu06ymgiIUD+fF6pPtgxXrAeditNOAbjGZpWh2pMggx1B6dcO/KJ7FckVbGCg/gs7ut/fyGU6H
nUVS9bfXTNTzl5sv4XNJl1/3oMRO4Tj1Liq5W+ZXzhz0r0S+WTbY0UPWYzmrcLvgokhrP9NKbNvk
MmODF6x56S8fd3+Hr+U8ZcwPYqlwHBr6nedUWAOeSl+Xr/awICk7fy/2tM2Ut6CfMZbh7D3I6BI6
vBujxG9hwVOHRRaMe9D3AWC+CcLS/3DaUfRzr4luHXgsxfaNI78iMBwOfRPdkAe0S+LUtmvWzfMd
h1s9t8jfbgQC66cWdVc+ROy41C/yszZgUZNiQCw22olMmhe2uTHLGDstCt8dbAf/g7tmkcwgO723
lZVKH2VPV/X1ZjBVuVTtS2eftBBQ1Doit07AzX4cUCtGyt7mzxUHaE5De/4E3jELG5SpA+UXARLQ
xTy8Ja8b/9EOt6QQSIPuHexu59GVCVNRVfonyv7ASRE0zR8iCacU8v5bHwRSgNVIv8lnOpai56EE
LPKyHcS8l/D0jA8CoS8kk5ZKX3I1J5SHSL3YnYLWVa4VrgZtYe6XlLReYsxIlBwTtLeuN10QisJp
jyue0BiUSwMkOax7SOGVlJ/BuTRTxKnJ4RtnLMpSZdnQQFHOVQSISiDcWpFXyZZkGdW2LOJnJyR9
dOFlq/7S1bM77VmKscK+rkRs/zDfmPeTl33i38qvkclv1s0N0au2uMsPKmKT8J7JUA4gEk2Hne3U
sjolnwahsbBBncY7yoSbbevq35+OAA7+siprGPSEemvgP96RSKXFH38Xzgm5icBTyEHf3pXJNIj6
uoYPLxEGlWrH9q5P/WsKnCLmZGfTgEaWLb+YKYkHmI3tyJo4aBoxPJ903rQ6eL1E00eHZdW5rOBq
la6xRzkcnIeQ7iYohxbJcnCPbbC8Hk0rty4KzXHLX0q1t2943VJeeXEM5hWWz3jdZFVupMhOHnm4
eDCsAWB3l/pZ0+fHFnLl79qfHuIMlpwhjVknMPUGDq6PxbE0sEPqHBmofV9Htl0pf1VSI8hywbO3
1Blfl05IbqFlW8mEMV9l5W1HeELAbhj5mOXwZKe94pFKFG60paoBoE6gAqBVMfot6+0jaFP+hTtl
KlU2a2U5JMHCwfZcNf6jTCZUPzCL2BBhUFsjkCimztXjy5Rq3ua4uwjFUVRwanGQyNJ2k2fHv/cu
zXlq94W1Ril5xHtdOjJgH2dSZYzOxGx6wODxMsTiAfjHfY/HHOklG0gqFAXYlQsU8MjqY4FcnBQo
EAS/qYUHRgt3o4TvZdkebTDFyJlRPaaE/K1a+1cOok6/xj1oMKa08bR0ifPjOuannVz1hF8c8Vn8
lVRGdDP2tom9m2qmxdrIKr0/5SvrCII8Pc9Fg8QgP9oS4aa9fzo37YaSU4Ansdh1VqhZ1WKVpIy0
/uTUw8/SE4ON9hqHwxLEFjWfezy5q35fa1PdJPGKgcpdaxSdQgo6wCfM2UUGF/vaNxajKG1N8PNw
MxEjg7mtIkxI8Jsj/Y2zIyI8PwV8WO5pZHob6oIvI1eUQjZcqphjnR9pMSpso7/kYcoXunssWsjp
tkknr/HdaFGJWQluv/n95ltt3cqkfLNnWb/rHRvZBfnaqcXiw5vCpz9MO3jv8uBRU8NEManHUZVp
rORpGt1kEwSchtef7atzzPO/VyyCKxpARKRiNj0LcfMn+I7WzQiMQ8kWicNsBcTFPezr92yp25c6
N46IwNyRSDSZU4NQMn+KxofVBS2zF9dr6uXlQr8mWIVhmEs8uuTwDEPCI2ndCqVNUkElNtXTmB+L
A+9vVSwIaub2STq2vr7fwZiNjeDmnOtLiBsKC5aAtEG9XopNFlRpSP9jCGFa6aRcUpLkkd12LBvr
zFE/6+vpwOTU+CyRlc0d/IOjcPjPGgGUEalRoYC2ggiJWgIstbBgN2XTLoWdqI1I9mtz8wRZgFMw
M/OHx3TSCRV/ruFWYMBTfe157xlS0TQXmxf6fZw4nizXZBtz6sXEEmskXPiFhOymqWXsYRwjJu7q
DoV07PKK/Y5reD04sbw6rB0pjpwfxdVbLe+6OGAITZQH8ZK84bRF8PLbbr2jw0jwFeHnv6p9tux/
IAQBL/CMWPPi1DMzeNWXiT6J2wPhvElTHGYVE/k1MWhkYUjwXSprd+72r4zO3NncFsmOLjiWoNAy
tYIiG8mBoY2JnIgp9dLH6wGg6nsYknhqDhz2ItU+eqAv9AJ9wjmFq0MjRmYlS3Prp7QWiuM2GFaN
4Cj2R2TTcpdO6usDccCMac9+BBsJ0rYA7OQhQ0rDdyX9Yo5jMeCEwMcituRP+i9o32aDOdxATwcH
AoypwdBh6R6LLLw0EEPs38my/al1qljohicwPdmd2TsnjWDx9x8HvBxA0WUswFcNFj6kIJcWeRdL
x7DDxYEZwHKYhKeHQgN3H2Ss742kthvu9mZ2cNfjDZvZFsG9sOVbz1/80eUbX7HvbWJ6Pw+2UCXX
nVS+x6nxIf9Pji3BHNSeDn8VlxVY4e01G4Sp771mEbHXedx76WAyUzcT47ToqYRVNMPF4czP07UH
oeJidQM7AeLjArwlMynLF7jlHJY6KtNuDNzvaaq0mhYuiXMpQ4tefclIk7b6iJ5MtAENee1C+6Yf
bE4RRfHQn9j8w21sF4a0lqusz4fSpzFwXFuYgxuoUlaHBwELVvh0F/zF7Y1HmTUVbO/RYh0ejPfh
THZ12jc4e+eHLMIWsSut43uIYZozvCP6cVFiauWB3HmHCKdKJ+DOWgLJCsfzJalP710YMSZWYpKm
KWyyQcjuzEZPacwqPH9VkZeMsCBbgvsGffssYIrcn1b8grrUk2Y0VxZQXlyvFr/WZEwd+++08KY1
F2RXBsu9Uk/siVYC9EeIMOhOXj2C0iXkDd7ynfctg3qRcI4B8gVKuBtWZVLfflPMROpHf4aPgixZ
oHnk8Qwj+qc5MfcWiIzo43GJVZ4qSXgMwb3kxgFU5yCUkckg7ZTL6TgJknrr/BKZJad6aZ0yL1T1
34RLeLLF/q4K51fXvRAIOH5Q8JMxCsB8Z7vw0os9v8u2oRYus89LXAzbpEMHiNnqtisYJXh3x/S5
fjQoW3V4mAFwcJO+mN7HXDNhI/jYqVVePenqWQNt7TAU+tHwEnHtM324rCeoZhVSuyJrGBK6ZTNj
Ug2crpAxUWV8BzYhMMaXmccutFSU5GKZc03/Hqz4i2jGsWOPUvmQCnTNVqjcCfu2lCNBa3P7kweT
qnTt7YzV/xGalzB7pmQvYULNYvzQhZMMfRUH/gFUeBzxpmxioODmKTtv/JZqi/8CgMRVk5vQCVYA
0dHIm5RBov16f1y50VL6cmcIlNYsxdwjC0gKHnkSAxOKk4H9BGgAheuGt5wNW1wBCvgd0XUfD91J
jFqpdSApbfhqewEqwLGfMSAeqVzApubuam0AhOzaY0kUEy/u+MmYmWjkn46nGC7vFfT+uwJ3CWAz
dX1yEL2ElW/D8M0bBL12uKzRrx2pHB6SWGjZ0APPP5hQUDF4ZvfD5ch/DIlf0QafXnJXRcruX4q7
YQ+E1JzSUPhz0y30d+UqnjRsYY9XplkUB21X6UVMX3IAL7PfeWyZCHs6X5ROv2QrqH0ynA1tY6GR
uXhpDPw21zphUTlIfRNQRIzIQ3eZ5Bh5V3xSWbnfCmKO9vI5uC672j9GO9RkdTJmSerTV+7o7eTk
4Koj3MEmLF6tcTNfBZuUiaWndrV7bmDe0z+/rSxJPhtZuZ9LhHzkgqvfDANhFHriYYA+aYmutprc
AmGvyzQfolZHFpbphzXt9tNyAE4cOUiW0oOdQEfxWB6fQpGyadd59XM7IUOnetchWagu/zRT7qxv
Ucr53tYN0N80FkjSzUcU5pRTBeYKfQYADd7FuHGn7PrBE2dEKMMq3dVJdaV21uvGMnqooc2aJaI4
5cgpgNYM8Ko6koumvU0lO40YApojQgggDB1BOAcPbI/gbZySf7R5PTHVBbEB3YdK20lpaJcA9/S5
2+J2aj6wZCgz5vh/af1UDuoetmv84y48nxJwxq7kZocLeOuL7QI0VWkINXym1tA1NczjEpNStrvL
Hp3ExfKEYJ9yMqzCq59cDegpNndB7wS2m8dxtqBCZQAZ7IV+pgs8Ad6i0ZW8RMY5NZSwieS49x+X
Fh8qtDrRYjKGvruQjeVZGuj1yMYCdvMS9xORb4Vzj0m4dwLr6k/4WlDwsywtiYMp82se80yqzdYg
/Nu1A9jya3tlJopajMk05DF+Lseps814/EoV/TGndrt0JvllJtxh3kV1na4nlHzvY+OsX7FIEGnI
sIe++GfdU8rqiC3VXaYnGQHGkSnp4KIl+3JoyieVRzY0LNdS8mvQagn35xZEYV1pQYyMViBuwLCg
4Osg/GA3bC6NOOCqtTFdIR2NxVstygL7jZLBAKELbFyDMPopor1PyGJ4K+rvwaaY5Vy0309LzI8B
K6kE+bq+GStMQteBvcqu6TFyG3zNIhIBItu+uuNlysk18sbb7EQC6Iijc1Te3FSoY3numDbJjvnQ
lkGYcyhlqye0o2YahZc23eMbqVoHq3rYu3CtodfOx4FYFZoTKGzEabFQ7d7LRLC3TlDMirGrgwKS
ghYUp4kZtEZge7BLbjuUKcdCtFq2gL74deOifTOS5COyw7aMJyAcaXSJUlki5M93FFR7qL4adLF5
66q8cs714cppSJ0q1rpXPxnMAobjm2q4gv+kqXDdCxyPAdjXE4Humw32dr1C3qu5tPPPvLEp9W0g
gIISz+GjQJ1g+rvo7f2EQJTyqZiynQTD3GtDBSCEKibqfshIvmnLhtixv3gwv7IVh8aNjOanBAHL
lmnU/UJIznkCuTluOJnnUmCAFzqT+lHQDLHL2cx5j9JQxnPMWhOiSOdCs6MW1qDS6ezpwk5J01bn
LJrdY+FTl4mHa7ofIQyIXx7aPnAs4GwL5/Ll1IkwSiXqz4nvr04jjnEabH/+M3LDGDr48MB7JGEu
SseAwQXMiv8DgK1KdVUkbTjd47VXlwaacRZx7hjtrCa5VLHksZtTmCZIqgsD2jFjzCEOvGD44F7x
cMVZ79cZsoCv3tcFnizNrBsTngxSLN1m1/CqtrJzAw6nM+c82N3pUTlM+oCwI1J/XPPAdHlIZ/jq
y3Fz4drkfhSiwr+ISfSZQ3VkvC1JBX5dcsd5Kurwwvd/+sEJOo0JEOa/W60MP8+PRiSReU7YmUXK
Q+Ucw5Z7bZ6XbtGSdmks97IKnJkgqGP+nCUDW+yDNh2jAAxiNl/Fq+RGj4QCf5AFYnMxoy0hytTi
gfTn36kSVBYLKv2umFYN5C6clWilczSxXJ2RTfLuq8Llroke7e7+kj/VM1DRwhZBb1OfbbxvaVX1
aFsig/rc5ovkHt5sRkNbp594D7rU0eBC2DP4KjTBpJvoAe3ANVijA5ehfEa0YTMFowLpL3qt+XxV
Butq9GrB7Lvqz0W6QToaSXjU4d7N15BjbiPytDAuIlXIjf4P0F+L6j9lPB0e4q9VVUXA20IOqPo8
W2H6TYh0C9hKMgEXlY1/CPNaCafSL7HNldLhWI8jnQSP57rCPwsGZ1LWW9IKYJ3yggZF2mNSPEr0
Cqheg4vKt3yhFGewga6ecvC58f/gFJco8zONe88QS2Nd5tQr5d+opnEiBRcaTfBZbHoffYUxBj6M
7JhhJLPJ0LTq+jUhqaGj/uaQDcxTc7Q4+g85OVzPPqTH2UNirwNblRixvshka7xmmtFRGjgNNmpj
qVPIur+v2pTDLqpCLRf3BtNGejqo9Z9b1BEwPmoCcdxomDU9zaUi92TTDxjdlrZ8U/6w1Kk8CMsp
893okMzCQPPNc/d4HcNqUC2mxhpa7XqtkhoqBz1i+mJxNBVyYc17JedWLLkia6QPQ+U76wrXCCZJ
pIOPhd7lvl67If9MIic25iAI7PfAmA5BjgfBUXPSAhRQ8HvRvvyE0aYFzdsgMdFuhUSezg/mupqp
LH8ZqVbvK5lLlaqw6dSoEklGWU3TPMf4JOJdr45hkyUgiEybqpSPxNYFXyqu+RjJMtZkL0fD4lqM
ZXjSD3l+kALWhLj5Xk2Hlb9wkCdn8OkymlDsEXdWmOsNBzb0SVgQzZLBeFrTAqKL+wOTTrAgpbY9
XX9ZrdjMAWEZm3AkpRv5DztxNESXaLVw1dP1DhPQW2k0elh8U0yZ+Hbd25RKOGHeF4YDBqtWwWFk
5MclOqDmndfMMMLge7PaQOmAvy+q/pmtNXlZ1fCgWcH4et4C0E7kMrH8Lm5pBo67CsSv+6RD23qt
dFjKE8Gtjc5LMIFW0CWZKSJ0JNBvupjyC2L9VmNpi45Hm4CMsa08nZNrPZkMCj2QNch9WvubrTt8
+iRXSliAiYwSM5sg8ZbsIyGnExBiv0Hzozzle8H1JcE6YjwkVoBziYyOpq/AOQw63xj/e9ly9/QQ
04v2TRiw/5AnsJINv42LxUIED6XDAfJ7zXiyhZOq2hrpF7awjHiI3qgpCJTImEhMp7+MwMN5auH1
b+xM9vdIg9dyw5urU3WtB7VGxmCUK04ShPBfe8oKA+aSmZ75cQQeTebP/KielBGlmjCx2G5xLTe+
UQw0i23LcjGoek9Nbh9OzT1fvAx2F1+mZZ8mPfeUAZWYBSrpkvkD58FhY91SG4NFozX6FlzCMYLq
NLmkRmbyvBrsoYafuf04/OO5TcMKkSIxKLS53ST27sKaA3yw1xs1pZrZiIt4lfUBWcSolOqw81gC
bjSH9T5SHE9P9tUc7WvNmLWBNIvo8xIzoz0ZkR2Rs+0iPyOciGTcL8dAHa9EvAlOA16fHRFOJj9F
7Ae0hOcrQB1tk0vPY4anG6Ff7b7lbR44HkHlYc548OOfXJCOLYWo9Q9IizVv2sUt58qWPA4gMVhg
InG5294uGAb4IAiD2vJgOGp9PQVWJIhiKL2lTfromy0GNyvfV6es4xgLWED6D7LWq88Yd5Wrl6hy
vIzQQPovfOXUWzg6HWnwCwc50r1+ewxb4CEEqA//7HWS1Yyl6ZMmRF5seDSArmdzRjysndUUqZ5Z
MWnWf9B5WzX8UCWO7YxDjqwZPd1ZqCfDvIDgZILLSwfwrm4hRG7hmUG/5JSmQRUChXr90ewpYX8I
nwl/+yiRb/kOTIFexg2ZKVu18vhi8gerD7kcSGD0mWsTHWNOmNmBaMM97sq2crSNJ9R6zy4BuqXK
Yzs73Y1JCyDJMvkRrTI91IW5RDzn7p/34NTGHUJHyyhh6PSw5S1Qq2WpW4AV2OzwlKjVA3Mp8+Dv
i+Ct4EPQG24Zv7pPEa6KINhCe+JiJtthFkbqGrZZN4pACVb0jrMMqEfBXPJaio7hNHeL2qmIMl1q
8CLCYImopuc8TSZ1jIm/dkDtP6ASNLLb4kyN/7R9OeNNQyHrzAmLocr113+1arqXrxU8JO7BMCG7
l6GKs1J0lQK+z7NBiP4jkI1pVi7Biv8CIVmhuKT3RGZdAem/2CjzhidnoRnZlj1W8KNKft/0gghu
p7Z2CIzHqZlhF02sH/0/5c65XT/amU+mOFxpmH34c1ApuDsfGb9LL4wfomUQkIG1JBWTxIzlxXbj
R9yr80xX+cgoF48bDUvuYiOmonhvmn1b19Q/Wxzz9Q2OfMcIMzdIp3oMcsHhabuR+R2jDtE/OwAg
SAU4OVJEFQ83X7avYLVHfVrt3NJw2T5cWTzFyuGpuHcDCuIdf3cj5gAwDwrzDviQNbHt4O93TFOU
OYgFOTcpdLnLFq4RMkSIYAFo2mBt5r9OYZwn4UDDiSjXzeKjrXTP1XmwqjJ9xNVXqSLsereg6+QC
eKSikmMFg7dwBhqm8Bu1S/2I0Zuo9uDaOZRrK2Sr1PVpr4iIKaV3YrVR4W9mTwzKeOR2rptyKJeu
hv1xRRwgL+sVMM0kcE0t2Isqv/+XzPf6jbOoKhqo0RXHOBokL+rJnddnZ+sMThLasERPRimmiwvw
PFMDDB5yIA+0cD/PzbHoM0N8Wou9sMKR+dIotc1PexqAyQik6bJ6/mGd24Jio6e0+nilTDTbT9CQ
tvm0xhhZvg9KKnzjcvFP8IXbvbwjYMzaxkifxM/U5hUKsdjJD86V4RV0Dvg9aYwMrWXWqH9D6GKu
jqCf2IggwbxX/R9ObUCF2hZbHp6ZJbSWp/Or+99wAoxgXhZ/v2Eo7gFEG6J/ua7jPmf8MRMThtZy
2ezNArsg+zxNfklgKGyT9cBsS5NAF4FqsBx5BxCpGbcIqB407NKkvUjinE3iIW5RQzxrnVkoJjAm
il0iV7p1EhXkm1fJUuesRV+OSOeAlwd82gec2lXu7J2gPUsufk8tPO0KLqj5ctqvvfbvwrEsZBZw
mbbSfDfdD1djJNhSQlg1O/e3VaE76pJt4fpmUB3Fo1pr1hzsLRCZOf4jqGD1szXhOmusm+WApGcm
faWVSfg+l6q19cLQeiWaBLDxRLnAsY98SrhQ9vDa3TNM9n0phBuyf+58ydhStI8+vYBk/vy0+4jf
BJZEtM6fUPGua3KT1+MLIaLqTmWB5p+g/2Qh9gnt9dJ7Kon1ALkWEQVOP4tgFy3PJcD6L3T2IJak
WU9kv70zezXPFnXMspmx2D7jFaXbYhbuX/2zB/FPZiynTejpoyJ8pWEX4LUNZLKuoTYObn/zIuHF
D+CN5GPv1IOeOvp9qQJR+/8K8msgRE0cmsr3MAkVkmvN5CqshJ4j9NeyJnH1s5R2IRfa8uoPhO9E
0x5AcpL1YsCoKjxaMDjMt0RVyBZ5ZTEv2LuVN0mTDeMYk+5Wx8bqNJn1679pyK8UHWzxFJxQQs9w
CllR+QiTEPwRqwrSBESj2+bw9vqXsNIg0/mZSaaTI93ZQlOZWtNf/n2SZYi185Wrq/K3e41p0ZK1
AndWuBh+fI2MzG3N8njTJmmcMPL3HT26lko4aJx8CeL07HJKb6b4YT3RpeH4htDQ1FiFzoPeD1Ci
NKxpfSrtyZJU7IKrWjJ2zWQVxbJS5TPF22jOzoWSaw==
`pragma protect end_protected
