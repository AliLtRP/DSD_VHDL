// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ey3QD/hJ8aKLqkCzBe680+FvTTkKwY4c1nmBJZCanRwo5SvHvKaypdUBTHpymv24
XQodNHyxDCa8IghT2m0PcsmplTtZ064yO9ZNoegJyrbOc5qSLrNkZWodnukIFE/7
CastDY7GI4llQO6siYnPz92F4UrppeBMchbNygg870o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 42576)
gVc7794BEt3EFIYiAVSMUirTl0cNC+Ys30pI+zKOCg8rLoIgw4WjU2Q3PIdg/7Cl
8P8LJzR/ohUPOIxfu3sJUiOomLF+HgUNbVIboLkUA2bFdLtA7IXLRjn2+zR8SXs9
aAqyY/oEA0epqZ6LAWe4fQmcqR72z7doOfO7KCwGJbl1jUV6IGi8bStNeG9vVxkv
VCMoQq9feeqs/oIsDbaGp+7mehpXb3IbDLG33T6AzRJuEO9OJa24OXnDT2KkLeTd
KSPagdKKMOPpjWWdLkrNm3+rjv8e19xMmW5fthpqqw0LlQbVcDtElnA59Ecn8MY0
1m/0dTvujtwH3MM9fr+oCG7+VdxtsWmzEz4vLSuzO8eaBWu/XglcxbBraxUq0A0k
sain1do8T0iBxo6DL7puwxArBbcTDjOxNKyJO1ubjK/fAs7MTZ/g/OkuKPzbzWJg
NniAy0H4ixgLqSNu+a7EwOHRw2ZchZEN4MCNg5setVZxKEqjczPQGv/f4lLPCWzk
a6p3Jp25G1D0yySjpQzBkN9QdQr/wNoFMscQadc1gRByag6aCr3nz0kG9tJ6mpKx
GdmNKFj+xav8Sms5q6ewLB1t08uFuS5rMX/tcYcpZYTYWimC9lgukIC8UY7SpesR
SjEmr7TOMQK8exclJ7CNDOzBT+IvClEcGpM6atBaORmKTW8agDwSoEc9qh7fn1jP
vMx7Ppjfkjr3Cq1UbLT0cjKwfPns8PIde7p1bvYEKf1pJCPY225lYGKFwPaoZ5O+
EUo98JZL2ew3CLqXkvYH1uymbqbsMZZ1pN+78J7U8jKd7p5YXOTdV8OP7f+fDDAM
uhDpBhgYeb6olUHMb4RGGO06I9eLbO51Ik4DseiK1qfr9h0hHJILr8YIljh7AP1e
a1b8Cv9PrqB+sKpBCLPLy6RYzdWf8ZQ1O7oF3ypYAmXLDF2rFZIKdDgJJN7D9pTQ
jVR4zlgxmq77B2uvU/YteqhDPF0pJkCpI8aXAnFWbkM1ghcq3yP6wUOo5OUX5vEs
GVmmBqx0/O8UHUSz8xD32YGdfZ5P6iZk8/HpXeYNyA8IuzgO75NzQXIHiAksA/8w
HnuZQ2AANjzOlo+Hp64F/wrvo06cLid6h0QvJC9kdPXAK1mNZLN9mCyvy/lejF2I
tAIyTfFGSmaXPaEGsw8vpcYFWfhMJFxumEuneOEuzLhwIndSn7lisL9S8FqNIZ5Z
Jr/SJDJm/ZdN7X6nMBusGOisRYUDZMchlAVgewFcO7fKP521Dp6OBTYveRcJEhwa
ipxdMIeE4cNgxAc6z9IfrSThLe21ewWrnWfVezk+zh1tvegqILrnzd97XGwp/fhv
ID6gHGNFYssfwkmPGyhraXRxvqQIZ20Dy5YF93O68/WWkdVtJweMhd8HQyX3FGiI
2lEVsMmHhoFypg68UtL/l97ojPk+AJHaj5r+L7ASQcijKCc8MQ5mSNW/H4zJYLKH
58LAOeQs9mzPFk+JTSf6ZJ2JgHiHoPwUwExz4DBIG7LpwynBeme0dnj98dWRwSbY
+LWjT6vPhU9ku2DiNpdcKDjbShHNv5yiIBNe9gFQI04E5R4bD6VUo6hqX7lF6szJ
0L5RFFeEY4gEn+q1GiFiwaPXWrx+Fhkl6vc5XpfNLdDJsfULc5RzMOd9o3GnqMcc
vvKUXUAJJnRYtl9eQaUuOhM4qnmJoE8P/IgzQyuExVjwayuw38lLmZKnDQWUI8Ow
uwWRG3oLrf3sNbPQ2zy4RY0UD3wotbbM22gvBkvc6ksgnCS24EKHLE+l/LKWfPCn
7tIbSPblv1JaElMg7E8Zf4kBgl/4PYcWNIBAeSMINvfp6z5n5DHAAi34c3pztj5y
/R1pLmeVGa1dGFtqaT2RK5w9BKqu/e4bFhV5RZJTU6qNEScUXq98SxOWrBCFM6jl
KYAseEP38jDYJkj5CUM1lZMBehB4Jx9gmmCS9p6cnLL4mfak79//rCQRfjaDJHu8
cFLyTvuWegjKyHrgHz8QOqEKxcb0ZlVWXiPDSTihEGcEWAPlZbintf65xc6TzvmT
Bb+JORKEhnjZBqAQ/3WbqKKV+8ON7p4EeNr9CSB81lu1xIoHBeEdIViBWb1RUMzy
gG9DqhLgucHv3JYnQxGL5eeQY/t0DQXXIddKtn9qdhz1wS+czVQP/t4F1+FEHhkA
oiFif6YgXbM1sUfIfQcK6cpllc6pZYZQi0lY8Lv3VACHsr0a6HX5xNPPMgiQIATR
B6BX/E5P07lq0m9rejQL8ABJX9PRfsVcUdX92gT+yiv0GXHBUxgKe3KB6E9uaOI+
6kFQw3dQf3yO4tMzFMdfGVdF4jgJ5fXcPVGURWUUL5pU+Rc5d7YTyAxM7xpvB+fD
LWjtbtfxLJqBU5nVe9xRnsdRTPPKfcRFZB2ZTZ92tLtqxEPzRL20DYnc31IFEE0u
DYBCku9T/fA7K/Y3tsQseOGizj5XweSk1pGsCUX23Nf5s4FHoIV2Vaantq0vdEpH
scfreLfawDD0lkbcgKmynw6gy4cI0iEreSn8CyV40f9TtFWPhRjGr4uI5Plu2TSN
2eBx6gr65eL3RJH3r7HFnrxmVfIzL/BjFpphNlPWrSbXbLOzLz/5KIHCdGAxv2PC
PAztXxezjdEH+IDm6CxJLSDoR7sacwq5Jc5DSxDQbiZCZfenknTG2M5IoGTnHOqz
sEtMlhs7NYKB98z0cQR2JKdyJjfL6vGquJSgfKfvaFqFYKPM4EV6KqZK7xqDwzS9
LJIUg8+G8ZF2LAWi4jRCpcWzlgXrlUGzd3n/sRh+HqXQ+iEW0lOZftX6D4iCZn80
+b4yfaGhRSG+DYKX2JRx5TG5QyiL0owni8Zw3XdLwDia1Ki+BFVJ99w7jhDTB9Lq
ZESpvUgNt2VSqy9WeVzmlGP3w6PdUxtyuEx7OTn4lKR/bx5upTF/VVJzsyES+FqQ
DLmqCElFVR7vgsYCySgq1v+DoEgL1ME+yRokVK722HncgR9nJbgGag4EsRsdYLZF
5jFpsu9NwFGpgj7HXVtN4WRCEUnuNKByGqgIkSsLUOUOXNVbsXu0mjC+UkdxvtCz
HJbaQPhNHcmrWsZaGi4TI0H9/faGNMIaTMPiNWwGWtGQKS4J/Ld4MLGUjgeyNFTq
AK2mBaaF51pNZCK/jDE/jOdJdhCYZPkX4kY6hchablJbweVKiqMYkt4LKPvX5z4x
1lz2H9F8ZxdDBlZApj8V+9kAJLPt8w7isnAnDURUFbRgr0gPoG4yATJf7E0/EU5a
64TcwtD7FuZEH7onyrIVJc95Wm7Mh1LTTmIjcjFcwK4ZCzhLxCLxALNFMv/TaTFN
Em3eUJkoRfDmNpM0ApOoBA627ZJPMiVjcfKQejikIWd5ADqUeSP4iYtcmHxEjflN
dYwUePd8ahuM1RpGtSNyE9VOPUNDY6wOJZ2+BY4rP3OnO0J5I+RoYgaZIm0FTx2l
iHkj3zEtGy3C/qq+MzZjcr+J++WrTH7mj4heEvWnbi5WhbPAWr9SPl/MSVc6bU3f
4MzNRmMmI1ItyCgqiSvF08y2PT1FxBBcd/XV+dyPTd9HlXqJ/GSDeNtjueyGavf4
pLBqqlX75k2a4pJ9PzBVhXZwO63JjZmOc2kJeBK8jA0kLCtyhqKr5eVqTndIVFVs
jhlb5gjmVfk0n83Luu75WO5nuj+dq0z56QC5gOJ7fiC9a73eBUI/BXPkJF0KFROs
25ViyVVdAx0RjFtma0VUK3H+Z3+ZeQd/3241iQgbGzuiXJXzGi7sFGlw6Qc1b6JP
UXBZ7Ifwtb+700kLElLV3FGUW7bCL09j7N+2/W5T46qAIg5wdNm2vmQ+sO2dbZro
z862flrXUJbe9k8yWhkU79YpyNXDh79nG2Q27Cek5q1yPZG1IzKVk0MapY/xmKyi
luHygy3KB+MPgbdasKdGWjnjdYsB7msT5kRtmisHbYj3xZJPRERnCcGU9QHutRS3
8sLIYATPBmpzT2DQu1s/FkWVadhRvSJoRT0fiLK/Ir4tJCweOpeA3xUaXn/7O37f
hir0WeZptalW2Ont033iuOg7YiUt7XR0CXF1Dedm4mfGyKiTxsiWC2bCHeiAT0ih
7gP6QWC3rOW9Njrdo4E7DrGEQcY4OzIG/gckOm5Ya81wQ8ovhdrDatzynfyvTNz8
O4ylcVgG5kveAKiRhi22YtTyQEtTHH3lrfcucnGJasP6k3b4TPM7BVH3ax/mMrL4
ylCuDvTI3LKm4TxDT5hz4p2sQQnO8ShuCwAaNWigGBSZMyYqcmBKkN66QaloszEv
qOI/XdRu0p4g9jfWqK8FzfwC/JIHjtdA2zUPcJZK5sARvgXJd1dXN0YNZPK2FvKB
zzqCCrZlmytRptEwAZH/O/WvcfoYi4Q88j//Wbzqdt1iXKeQaIDrVtWJL77aSyKG
uLybdgPIoIaJrOGGJ24laKl2U8XBvSZ6PYl9iMIdjG1ypf3eg/2ncNkg2/hfe8Pp
B2pkHbkFAtr7s4q7eXEKuMaKcI4sX2kDyuvrW1TExmFARV+ir07mGco+nNqZJ5kX
EZIwICRKiboxYyF+YTLajBFJ+mAHW3w5027gIiEGpQCfBXMNUCm0g1OvDyT9U+kc
QwcN8yvBsJHx22Ofxt/HBClNh6x4c+UghmsLCP1NMlHvDo43mrrIM4O1wmF8AKE0
muzXM7nCgqGtymik5MROPFjkmjbJdXE7CUnhlt+ejSkgv0WlOlAT2J6/xQMHcctb
Y+z0vvkLLOZOXnDsQlqRt1CQZufvf4M58OOleRCJH+XSvCDdZPjdTNbp2QfLaT36
wbQMlusCIfT8v1k6RERGZyCa+lD6m/7qLrkTN5RtDT43AZF50SXLPp79TFogGoVK
MzSYCQ4CpVYLkNJtWyFyAY6YgUriBmFOIGo3WMxtKVwBZlIh57TLL0D7bkcpGDJe
8ZhGZqXt9Ja5FF5e8ogeIJeIuPxc3EZBxkvQTtADyC1HtLh+6g3De7hkDLE8FwCR
TA4OsmJVeDupPuYrJZKbAkHdZdnrwEo7T1rXJimvKtZVqehW1TwcpxjSmNWKHqxt
7Ei+anyexsRgfEXvvnwh1jGXLhKmEfbttcOzKmiZQHBAoeg09vyvlaPSOIgGKN23
l7rtWeH0qDRtPyIoA4BxumfeDIvetKmBD5+fiDue0idm3uRFr6FJwlBdjq1aZTp9
F8IDwBF0l4TbgdCrG+OQsTsKiDyMJpSkatGuOF4k3Y9/JhBgY5u9DtWT+cOr6pNE
5IfReua4g03RknU180/a0lsfTsW8AgGQknMpkXF7iw04OuCPyhpa/WOx9BXqvyEn
jaVjF2ckpyEsSu76ZBHN4fAxur4hX2F+ZGvhjIkGmu/aJI6+uI5J3eAdQoZmUcTM
kwh297f/yHwUyx4NKcRoe8dRY8Bd5xkggDajvwkyt7PJCqmBZZX54zdugIG1hfWz
/tHWlxZ23EtTejpewEonqM+Ey6uotTerGcbYARoULTXH2CtwypT8nyQk7twzXofr
noyYV5KccAOEN6U0PWPiJoDVS4LlM2IbbxqOUruKTQqQ991kz169XdOPMIpySBOG
z9x1IxnqM72azRj/E1fLp9UV9C0ydTao507uEUcOoF3eMKcRj4cZkIp/jflK/b4Z
C9r64+Tc4wtRp6z3Dw8UPFUj5tEQJa3g1vpNz+9nvCmkz4tjv2dVdRkCmN/OA9v4
kiDeBwJrXEoZ3MERUwSqR9EnHGzv0Ao+emtj3GdGKKDket9Xg5ldfbIvE3Xzv6Ge
x0pvokyvtQr26ImTrln7CIRTrw2kgjc/9vWIIF+/jNJbSYhOUBu9qVbSBf9zM4f9
VxVOuBH9DOvwfyCeFD8aP6qA6ayI5fhcq8DCCnVUtY7Zory8l5kEuhfF6unaOMYe
L2YuaKaxrRcD3Cf+biFdlYt64nbL+F7zNq8PPyxZU2sz5uBKhey21bIQj0OlyJz0
Y4X1s2Fk5EFjP2pHrryO11d1T/sTjEDZMnCa288t19KCvQBfKDhn2YkPH9xoTAzf
IX1ha31EwKuQpFp/kzU47BEPQDNhzx7/4PRIf4yMiFHlCiexquGsToKuPUMyv6UA
UqFX0Ju/ewkQSAPlAFk7UPMK/hPhgka+NvlDxkiQGmeyUSebEUJ04SZhrhLAuD5W
lpinCcMJUeHmrZbk97nSiTiWhH9QnObrOYu/k8iJGg3bJD7A7m69HNpgf3QLUKh8
ENwUo7KbITLQSThStzfRlg0SZ/x5cHg8MeQgcfbrfIGFZDN5z+dwX3i4gKeV3xsW
AYWGBcx5UeSkxG5WkZZ6evm6RrRQSnmwUHB5Jj3EkdfzpGnUfXIMJ97wQktW7+xx
qVEucgtPX/FiLXmX08IAS+B64Bh5WFtb/5LwwV0mBcfY6q/eWEo4GFu0SbEjR62Z
tue7ufTPiHkOJf7+PnmV8loHui0In10yHyJA4hUNNCu6KFZg2RFsaORZfEMSVl5X
80Ymjl0+Aex8lJx5JgbvqaDDlRifmw99lnfOqy3kBewbElevYE8lj3qcNL4PI954
Hk161bHMfa/qSaZYaNbkPJx6AJ+m1Dc06GcwHTieprvOirII8m8LJMNdOx9tNp62
MbZG1HNk9gvJk/V8yc6z3YJZDWizDGLRehtKQVbJO2JYgY5oJUlph0keBz0hlsgc
apUi92aHHE/jvHSFjrwKNrOvj+VUw4X3ZcRzeRayIs+M91R8dI+4vWXRo4QaxsVX
G+kV230zAx4SfoZI+LGjAzj0kAbqsjcbRuVruOUFJeZ5iUVSUzohrksTf5HMU9MP
f9sToxeeE55ksEzv/tZ6eXItLH2iLGu+iKajj/ZDnJ4UCE2yL3GDkTnmqlYzF42C
AuPCZhboqOAbACCO45kidi8eWRQv1GBz6eK2SZvxR1dD+w4K+fhVOPxjP7vXC3AR
H26GhwuWhJM75/u8s4We3vOvLW5NX0pQJYvaq1uH8VHNC//TEvWq39+tw+Rhtdk7
APYiXTIjjUwHzhm+EAqVptOGSi++oIts68ILlxMvwW6eT7jyW9tHvgmzk0HQU3ll
MKXqqIppLNBhLRFMeYTT36IV/G3Q0AQB4DO2MPuGrei0CiM4wp5KUtDdnEBpIX+z
yKoqJCXCpjgNWNFEvIkY74Y6Hp2rjAYBbP1n8sx58P3n7AtRC5ep3YSyZLxWVJDz
IJV6acWXY+stnVOyhpa2E858vTNLENMKIPRHW9u/OX2SXbtSfPgX7wAnIURJhOd4
613YC3tcEcnCsyt/hVFnp0y6XeBOAknrsXraXWlYkfT71vaBdG9NOST8rlYA9Rqo
k2W9CXDsxlQmo7ZnJTQJW06w2iTFf37E3BwE1Y19hbKcHOfMMW7X2a5i9GzS5JkO
kJD03PtxOe7n0m9jMmVFPRX0wlzxJrBYNu9KiDdKQWsBmISLUl30hu0bqIFG9ZNN
WT7SB40eMtBSj6+ojOlfhyUPu0nCJaphYjulFn+FtVPlV8T/10be/IcBokuHLt9z
V5UfOm0H7zshJUaiHbUWydh7H6SI3cibT+6iLdAHGsqyKbANMIjFKxlYd7KL+zKn
SS1jsJdNub5Fbkyy7X0/AV/O2FSkj87+c3BOf66qKhG3xhlu922nI6aB4jN2k6Cu
skR+JppmVfGEYxeJDWirULc66afgSM8WMPLqC1GEylfw+Jj+B69RswKxxwtq7S21
i770WnFJ8FNxNVQeD51C01HzSQ2896KRp+IYwt3bBftqb4HU+T1yrGKF+MknR16G
sVd6DXUzN/5t9KCncX1f+NSNwvPDF339EQ4e0c5fZtFdLEKc4vrXOauljwX4W6SI
I1+IhX8GiRineLGOo9dih2CEaoEfvbbVBcHpiaprDAOG1A6oEcR3a4NUixfnkZaY
RG71NFK+ehqscgT0uVqyIU655BSDhcD6riX8XQ3wvj4KcvsrrcCKnBEd0gp0heEA
sBpScklrr0R2ts+6yS3QWXXQOFMdgDR7+KEPRLWFa/vj/zcIfFwaJg4qhGlzLqlE
ZWckYG9/eK5EfTuz2JOqTmP+I5GKXOBAdC4fBrzhj6go1A8xDN3gP8tm3m/qOMhb
3HZdCclXxOG/fQMfe+6pCP6uNNSODFcoek4WMvPPYAcaRxXa6m/N9h96NI5o6YFp
g7DjK39unH1RRtbXEbHM2V6Ck9JZO/vrtmOe+gOPf4rI4prRjQZ+BoH/QX27DYUm
sgJzhaKsxc9qopaF7b0iy+s6Vaa8ZeBt+QAc/rKp2r/qynQ4mDV7DmRE5gDR6R7b
/OzJpFkPZUrOsgMa+jxspYvcTVaDxaIOX/dFxSJEMlUbBXxlFUCRgUu+wL9BALaz
2coh/F/r+NJwQ+dOvIbVhnh1v9c/cwiQ/bSTCO7ZlBZpRDX4bPVhjJqNJ1xgWHcC
pIBpB7N1RkUkT/78ezPCw4j4qSxm60QbQf0TJc/98KOAXtj8vw/kjuFxcmz1qD83
K0RYyzff9aCwiIbW2ytg+BoWFB1L8o4ked4XCbrRxxf62iiTHuRZ9uHhc8EZOj6x
nkxUpmT3yFXE2GACcZ0Z40u7D21XeGeBcoPBSZEwjzjIHfw+IlOt+kSpLFgfodcZ
hjk1l86qtUIvJMWzVy1ipdmTe1q13hwM9QSfCFOELEnC02eRGCKPRfDMZhUS+QZ0
PfLOUbkg1tn19tIUbDYJPXp8/8EkZKoq9pWyzLNbIzfBeiq8cDug+jeckEVad0CD
zU5UP2BklnuOU7bwfrvjGC7NSY7jtmBF7iUd7yUhulupLPlsYLzmXzzv8eiKOKwj
FlIxovBtiLqskRZVxqY8YNwSt/XnZwi06EDSyqnI+jm/UksG0tE5fxsrwz76qHDC
l21XMSGa+jBI2TR3E9D37YrBrZMSKntgDKw14tfKNGi4ywW0C8VwnBq9ciIVAwab
tS6JxhHQNvSGqfqB5uih0LcBL1exkqnidK6ax6NO1OlbmGtuwt3GDpvbrRePm1hr
lETr+WzhwF/CzzjquKpcUevVbeyxmsAliNRxY5H6q7gamtgpwNv/7jZqKdukbzbZ
1V6LVvJmFOFulvzzjtb63m6HRld2IM/3A4NocYAjfnDuSUALYTKkAamKPbNVlVPb
P2A5j51pUeBYbh1a/2zrsJVnMZBbtm9MpJBA+nhh5GrUfbLicpPXM5y2TU4rs2aU
3HLfJgQ4sDPkcvrtWD1Qf8rt32nFG0wjjhcnSXOb1mEbOMOvHTdVvL4egdx7n4mo
go/fPUvLVHlTjL7XF5ZnYL6v/9CLnHX31A40r9B0FOTDWLLK5kxmiiR2H3OceQPC
EWWKMqYXGT+66gv24RWYvefJ/jBEo6Jr/SjNEJbAkRvDdBWzNWXRTxxJ8sFdjuib
fCTvJgFNJIKgyb+3uQYaT592A0Oq0Ah34V1TlKHh4FGbqkpNO5TOomh54Np4+LWh
jfuG1wh/BeDqD6BEjo6OJu6Tw2qvu5rnlhjRUuf39HdtsgAS0F4TAbfpD3TsUF4E
eNlybeHjIML0rRtnBPvvh0h8UdeNexzyevgVxVsoReK5ZQQ2/z3lg4TCnXVbLaqe
EsMdEjeJ0OGrIjWHpqs7C4QRfaraJpsX0Niv+NZeG3S5VqNC6B0fAiHmsbozsJdX
baO+QRqkdEQ9exhwQ4lFStdnO4IxuSomUrabv3bh+zVeXOhsdoBgM1NyImgxtNSX
la9U8M3i1ydMrtLhi6umeJtACwh/ov5vje6BAMlssqN8LV0hdKSBylS7fihScHOX
SmehUoTm+e9N/Hs5JH2pIk/fmE/u78KVAXTVEyuhKY3nIPgDYSzsOzplDx5ZhsQo
6nYn6tXRx6fYHnZD0ozjjgzUETj5fj+lNQROfhaBwXj2Eez/7kjLBYxAhJ4g3goW
XhCyCDOozIsvnvjpTNY9TGWOw/dxz0WtthCEBM9X0VIFoF6UIXiuObIV7G/Cih5s
bEmWXB6wYiZdOYQyl3PLudhRYW/sK52QsF6xW/NKWvkjoGH81KNdbs1MXntDrnlv
qVOSy4QCikiM+Q2xSKCh+IZ7hQSl11LP9EJ/755zuUcrKXvg2jyH1bKXb0IIz0Vj
jykmlwvuEfWf77dbvnn/Qtsa4xJ5r6dR2E/L+MtnPe/5UsbeQbS9XoO4Fi1Sg9V+
Olb/uJ3+8yP+hkIPMp3JvVDmY89Qhbp1hWIw1MbBtSqlD0oW9K/Bcp+TC0cBlgo8
+6jaKBo7jPn4L+kzAxeBOGP0Z5ZaqGzYgs4n8ldnl+B8HfasxI/+enn0FSlpq+wN
oiFiL+IuwcelBkKlUnDj0ckj/lL1nxWDmayVUY3U0gjuKNmEqk86qqxzcciFH3EC
SLx7s9TbtfT+S9nI7Zwhp/5cgfwFuzE+eFy0yxPE6l8r1sNniSbb8lhkt6lohY3m
OTbg+AKKCGXfYNR49/tmFV5Kui2tGNVPqm7O7AwAslBkmAKs5m1c5iYpXMncG68y
PE+BpIAwBwerGnyElbYtJfZqD62YKQXLQkpX6DXsK7uLDRyn4ZaPhVji0aHilKMO
bxMpD5U/nQOZ+Xukyuadk4os+nL2yr4HuPwFHB0lbdpThwr/Aoi6afe/LJld1HeQ
f1xEH9vbtYCbo66tFJeNVFS6CSyvksD7bpkJlsYGTBDA9tDNvtThWRLbgb3E1Bqe
1RY7RDBTUJscMs6XGEdy2vKZookxStvxsSBvsjfDpCDKNqCYjQ/UahDGbJW7vjqD
XfbktZr4lVsKwiwWuqS5S+egF6u9U44zO/PCOv71SilbkX12FzSenstwdcnr1HhY
AHSKlBxMmZWTuSe1nGQ4ay9acwMRywzpS21aSz6ECEybzHKNzNJsi3unviAw5iTj
nlx8KXLqrkwHrBb0+sF0hL3x7yL4dW8XkL+1fttUHCT3vQVdlPox6r8X0RThHpYL
txAFs4bUgPl5FLVoIQ8qa3MDJbt5fM9a+KRZ8BYtDJYusy2/j/LovgGKCGldVImm
gtcUSL1gSooV5Ro70Yn+Jq6NLZ1GdPCjzrETFhSOeBh8V6+1HCvkTQlDkvqUkua4
xdoVsc6g6+jlgHBh/O1ORtylskrRfYMGSMqA65nl79lsZo1GQG6Qgt3+zKe42qt1
hONeUzaBSBB8dhYfdFWXjBXl3lBjGSOnISQ6pgHHl76PyucQ7wQYkKDoHW90ctIv
wbkp1rUcSqW0xp7bfSB30ybJgZxFvE6RBCvHeWjy+rNBtkTNizxsPGl4oyF2HynK
XRDy6Sq4kgV4Qo0djVTd0TVJ9zjfMe0dO+SRRfW51tZ5Kx7PhlncOnlXeGjCd8y6
7+tjMfkLT/DnIpgY6cKsU1WZy6Vs3gR3zLlvf8K73qASZxb6f01fWVRYadPDF9LP
26Vt1KRTCmPPLKXJNFnMTtkzpBC/6E4mLH+dYGlsb6EaOAp0MHyZz9syiq1DY55/
QoNVdYBVjbGPopde0725oLIhtZ8O1pne/zEQ8VCRE4XXWtoI0HOyKwkUPooxvOZm
pFZ9oxDoqz8lJUhbQ4YvwnB4oDbW5nACg7h/4cCtL1VV8XxF1HQZ9GEUCoW7E+Rj
kDxCtdGpyZGe++2dhV9pcPJixMZSnZvI9LcNaTvUhCCrP3F0GatIMVY1FhWpuUib
unZTI2V24HRFd5nVdakSaSBhrarRgODFi8lCrOnt+RjjslVMziOOT6UEvF4uLbCq
vOImNGXUkwp3jxEQ9EDzjOUT6z26Gg+FIcuHJvEJOju8TrxoI346eOpyzIcFUjzZ
3AFCk4Zvw+iUG73CbDmzOb/q/eXTX9mlzYEtHwjdWsHxtCTS7gFcRN5mb54IbUkl
Z1b2Fg6Rmv1EAYRG4ipD4Kxi2vfCWdpLrTh5Fys8lX+QoVyUZYCHvQ0/zvOEJXtT
SUfinb/38DyBbiEUYjbyLgGMjomQnr8wlggBujTRt0MmJnNCSnDzSzginNjGnwNu
hjTTPourPTqFzm/W1Mj02Ee8ypavIWAK3nDPoZ0yIW7dhYjaMCzelMZrfzIdETIZ
2hILHoYvbW5EZC7I3jKSrP9l9o5Cl+ZqeKO02txD2zffzIlkEoPLYl/Y/b+/R7Ux
JSjGlLQRKQwkIC1MRW2dZDqrQHcq3zOMb6LW590uRsgiEa0M9AiF0I2MLgI6WEvd
YgJVItnnD2cn1V7xO6AHu8CW1pbmHJiNNXpXvcHqaJkoWuJdxQ+jLkAu4Fc17NVc
BLEIAeKoU38YdSWGaLjQkKpUnaYWOzeosuKbO2ThC+lwJ0SoG8ZC9SDDrRsT9ANq
w/N6VOA3dQKpFmXZPuRy1yjdTvplX2pmsaJ4rjfOgrOqAsXkrX2yPDIEnC9H386i
JJIhIQhz4Ct1DP+IVlXICfpB7HCe6qJFFr7+b3mlK0Z97zgjvZgf7qk1oP6PrWge
Sdn9UL87tnbbuJDq8pIcGF2dQuv7u5itjuGJBYyZEKQ23sjK7+tso6PJf1Z5T/er
ndyKfylEWUlHeUaDBdgGHFkmtjaU6X/67CGg+jLTeT8L+VJcswxVmrxnaekQszTM
/CPs8V7ZY+GNG4UYP10oZ/OmgReZp9FN0QqBpFx/qpa/VjISrcmGxRCCveAJ/2PS
qDDYnaoXaSlMz/fAu37B1xq0Uy4Vwz1TCRdZBvOEJGm/3gmgvD3EP9iIuGgiGUQa
TVVdwjf1Kaf2bfRWeaZWPE70Q4pJXOYNOs2f14oCH1vahE5/wsjvdMC9PlfFQPz/
tZCuDNSdoivoVsv5t+SZMhSPYAotdaNIVjdXHcDAFgusxRKgA84nnLqEhx4MFStJ
5Xbdf543Njfcg37qz6Q2ItG4ragDumjJOjTek1QNDmupLUVJSn6rwX/xomN9Ihc5
ZfUUmR8E/hufcffBjhPXgPVkTi/1VQwc2O1NbEn14hgKFjZonvT6IfUFItcvuVbn
rL+pgKlLcC7AgxmW5mrKPSABcL6DV8vwyyDmZaXnAh8LVhsY1ogxBNInA0NKKZp7
fadspJRPokG1JRl9P7S91TXuzQpJXeRD4yfQQLaF+H1pGdM9AOa3bUDcnR85CJTU
wBOQd7NftxSVW/CFbNsIzTUeU93u34n8zpUSsPv3gwL1csqcjzwMIQ5BN0Yhq4wl
bcdQROVuZznUxB1x+2OgVQbS4yIP4k29blZLL2/glKerOh8ukya6or4pBkw+iR8G
v+w2WhKw2Eaeqb7hzwteDqVh2p9cNJldnAhwJ6JuGb/NeJ9MQuZbE6C4MBnRFcPM
CUfi2HCCRp5mSoC4wnt2FVFk0xf+dJJqWW0V/SS2nEm/Ml+LqA8Gfa/VjSbkm8F+
zPlzfZQ8EzzTr9ByxSAsAXz62JWmE3eU8Nnfi5Mff9T9Sg+4dXGKPxTrFM3wTenv
4yNM3B2avxA7yd2L6yEMaQjt0eXKrqC+M5cdHfUUn6uPp0yIRowB6A0u+Cu9gM6Z
61Y3+GZD5A0BvtSqMA8YwvT4CZ+M1WHbwcyduVUBmhTSzw3MPPB0xmbqhTlfPuSP
SjIKezK3vZg7FHNLeSrUFQDWYZDUpd65Xpl4JTij/Nxq0C1kVoJUZE7XyGjyNhCx
AwGRIgH4zyAwRVNcObcf0vI4/5fR5PTWzb39a7nLIY3/ihxXDrx1306j8otH08tF
PVVd7+eGpKmPr3HcJKa9+zvfvszYqwbJk+gwhpY0QlJMQ9zazYoLceaYNvH2xeXv
lN8hWsm+mwC0knTAd2C9DKoSf1x2LKty9Z5HBxqHSbB35uq3zjWtQ/NfkiOeJdad
+6+ww9nOpEHKhN66WtxDUi8BnFguFNQ4sWELU681J6NECcKghSpiSJA2horseYF4
olWUp4aD1t3o28I7w3IvLxB57KeWpYfxcIJcOt/GjMYWD60Jv3h0k5QkgN22EpaB
LvngauHP6Eb66yr5/sHmKeJnXdvv2zEhuHWsmI8OyWSBER6gmQHRH1j5dezhvanH
kEXPfhd5mfVTYwLgepVIMgjuasO1HfJmUEpcENBfQkm1SYo4TxXSQXD94+WHWPvN
KwhUd5d0Ym/aoRYK0+unHYpMctUf+t7CnUMFK5XNNvN3GDfEAnfLmRYgcEwWlRHd
3bsMiCb+Pslg0Q+RwmkTYrCHP0t+4AiIj0JvJwUlIUnfnYTbkyJOTIk5Cq4pY1oV
k7ybZsM5zrevD8Zd+izYnaS7tc7G85GXA/NlNWrp2UseVAoOWc6AAU7QvLAmeqdE
3R5EflnHZxjmHvoabh9CO16X4oAkY5TEjUYlYSc7Tj2vAbC5Knnenr0aHzeiRHKI
cxt8vXwAHVi+TNfLnh3AOserPFUi1Aazh3KxbijF7fu4cFPv1mrxeCVIVeS/Fy2X
vAmDubYUvD51kUQdNadENvpd67Xe7V9+HoIzG3xKiOI5/wzGhokXRfR3nIx/gZuS
zUJJi0PpURvX1YH53pCK5ICgbMQkt035SyED3wamgp1wmX5NFlBmZtCCHoyO7IRn
Tjt0rUxWqzOOz5/6iPaG2hUd7nwjbkEeyGtcT7tJsL5Dg6AvZUkgmcj/am0WU56B
y8MuYGTUmdAETdr0p31D/rhO+FQ89tRFvZswD8bDyEjx1vhIh2bUYwevS/ixw8ey
CZ2c02kf4RcN8JSa5EkmW3qLKiEyReAKD/N8LkQQRhoNmnScC87WOrdqnRPxjy2d
XuugaOtyEUkkg3H+vaCiydf1DJsTBD7TePnQCFdTlSlVTvFcDYhcZQr7lWPSdI89
sy1L0fMzZkWknYXkY9h70a4b2W9AK4kRo/Jez2fV0Zx9EljBGqdvz/bcIKsdmo/9
sCp9ctynS1LHs4Y0R4D98e/UnCZR1fZys/sOklVeaMoGxSvC60JJpeDNLWg+fij1
h0/uCd6z4JZUW42UwAdmmHUKOyE0fcwGonDDDiDaOjwMlGbDtIkqm1mVZBOwDi24
Y3ppGDZClkrSoQgiQqm1hH54192gw/80a52PcjzHsrBOi4gsuo5Kh00tAiOm+OI6
hraLmm15js6e0WjPNG+DN3j2yXXvyAtyowHw8PRnbRPOSr6QbTe3KRIgmoQNz7dp
hPeE7jY2bq4Zy+H5bF92MyX2WIkXqjuUFmdO86AID2tOiuk4PcsNZoTOzXYQ2i+7
2X+gYxWoD94iNPTMBV9pmrAmq1nwrur3i1uW8Lr3LUAAnE0gxwGeyD42hH21E1b0
LIq/dFWjBGrmqdmx0pvCHF7tkku1/nlblgxY12yUtDexTmfcECME+qZGkSMXDL7o
BAZwG5Q6k5uMMX4EvKccvmBmSs/+Vvf9xd81Z6LlCMfTnfHKam3GOxIgs2xIVFPB
D+5pykjSL/WNFO5wFeqgOt8XFvwmVIddsWrcavX/c7qobDsiVH6u+DVDN94brhp+
+1yCQVRHzLwEeV7RcBc967gy9cu8FxKHTbtL83hzXDoxHH5CW/quXd4Blk8TU7Ri
sf747/U/NoSf4Zr0ors3g72zafV13qy0+pOWd00l83FTCRMd6z3SXdWvbuhV/Ibq
dNPo8ZPTjuhoJLA7pHJtYRYIw/COu6a1YyS65rQufeJclIYQwxyl+JZ9OFDVwxO9
weYGPE+s8ylZM2v/SXlCoDJ1DVYpsCDreeVh4FNM8g/OFu/y1LuIf2lD1hRp3Ea7
TEpGXY4XYmKI/fQwCcA649wtTgt2+5ecjfIZswLT5qnw0lqC4zh7lTcqvIopRRr8
RwjbsfiaQc1GUQNoeRUOKmxbd0M5GAufnkETwy5XpsIGFo8zCywAlwxzuB1Updbp
ty7/181gN2gQnS4nMTzZGm7Ycd6WmNNttvfG9cdifLCT4tXTnIFgdyGbRVptAtRZ
CZxxRCF0bTtb8i6ta0yP7qjymnB1Ntwk/BJlVYmrqTE6u/uQ7q/HKrQHSKYLWQ4E
+T3ktVtWWuCmTN/XeOYO0Xso4VGD+SN0T9FaorM8+xowN0AaVEwg02MI7mv9/Nsg
GxLhQdjBCawTFpwtwPBrEexx7RM9LqsYS1BMGy5dGDAcVEeW3fAwamE3jhs2IKZB
5rrQ0q5CaIGNbLQ0wLd3A+RrEm1nqItyr+vtcqFGG+8aIwFid6JE6hY59wUqMFf6
NGoZRU6ueKY7K7nOjdBWldrFjWvOjtqEf5YGillt1S/HMiVWHkx0CROufSFaaFFk
N43A5Aqa9A/RRe+lqWarwYyBr0dYS31AEM5rUK+OgGzDACub+f/9nEtZV1oGWIUp
wnReCe0zGdqvf38G/GUfapcRAjFn9wiTfimHd4PP+HXLucKgH09fXU0NeEWG4KyV
cNEDE0YnjMfaEQKmnQbeASVRR7YXAZAK7FE80Jr2hhMGr8rhIr/LlvS46netF6Vw
GhqPt3fsxG2aiH+591j5cQYh7KkU7KnsEs/S8jBTE+KxlUQcpnXEGDpuvBwY6VbM
F+LVRJ8wwtztZkMGJcg5hpJuIjmdUlXWRKGRJfi3SHA6tTw5ftR2KdWfGveCV3Nu
HtmFctSkofQ0RsV+2j9xQwzwA1+zrx1VSunHedrj1d5wmPgo/xwnufC28ZpcO4gi
8zdrxJV/WWFhe2Bqz4xmwNIhYkoYTuHgVTKlXZ0tq0O1J9d7MkHR/6Xbp5bPnS4O
znFvQysfNDLqQ2LHYN13Yr+PoHSvlY0avpuBSUQTZ02GFrs5URBtnMsUjkI/OpMu
sxvmfDI/ququZCM0SNG/LGTnDsasVYwaex8Zxr48uHccsu2X7ZXIQoj44d0/c3Y+
FLJ80zOGBnJBv/25CX9RCkqMbqeYhP8Nv5Y1S8VsTlZtryuNS2+Qd6/1VCzuAfij
aRw5nnHxQdnKEMEKRvliua77CArVUEENe/2DiHPHanXSdM3TPgYE4hcFemKYlCno
gL7knmbJEgUFxpIM3FfdGBuItiG8ffhZAPrK+PPiXHYCo0uTp2tg/VVfCzOwXi4F
n4EUou0SVqRnjUw2nyuKaRPUHDBB46lna0PvZJj4R4T4xB+wIOxhOX//FZhV7Z8s
eQoVn8ykQNiSC398Jm4RIdPTMks4qkr6kfnY124OE2wRZjd8CgSnI0NPw8RPBKYd
BcGOK4aQXdGUFBw9uyGozmT2sf0Tij/t46vmcOicw/FPI80DLT/r6wFlj1dz/GeE
WGaz5NvlQnmG1K8M0sUp4RjT6HJNuPb4tSMjHaqEF2eg/0ETZxFqxhcCey+mfwpk
gPDOgDyrdsaEzdgfmNNoLxD8KFDYNxexFC6Fvtv687hDoZsy9M8S6HTQDby/kRsd
iZ2SHJfZ95Jb9KKxsGcQAn6SDbJdFmsJU3PCzt3urKBkCq6HRtdhrYJ6VJLKmqH8
l/WOAfP9tCAwFU+COqmjtRng4ufDCICzh+Wez/y+sunLSWQv1JHtCCa443rF2Z7N
UsZEKko0UJkEUh2MheMAOc6dZjgv+v8cB3ZKc1GDO0Ct8tUz3fL9Y8kvwQqsaWpO
Jgq4c7nM/O7zXm3mlDdRSWOhIfw7lY7zFDHJudVuCqJWqc3MiAKGRCMSGcSYRLOv
8ZNENUIQtRBX84J+gItUSAuNZJQzWILIlqzL129O+x4D/m20p5gq+f8JLbAzaFQ7
7wDf49ApQfCQ32JwW1rIpefOj7NCGeUC4LSKYl4kFFqI4R2nfBVcC7K6WiLoo0vc
wlZAXBEkNQNI0B/UNTH6nkeFEFAxKhBp4HZTwdHtrgmImqrHj/Q6zq+hNgN9CPMz
t0JgYzyWaVDI0qkCfgKVi9n9O3g0nZFia5knznH4Firzy/ZbYO0EtvMFJTgIWLpg
YSS0mpcW/TNWPJ6/WnnywZvq8fdtPs7+KKnuGiyWdvl/1xy6kOtnCExe8fpxUfXb
NW8etJb1EczQMUFeDZrTFsYR1Rund1ZjScCA637PbUQ2/9x6JWd16REUjgUcFDBy
30VsjTm8nCKC//vETtieLbFnUB83aSOBWKxfeIV7CKK5KIE0O99MrR1SVkDEZSDY
QRRU/SlLo+BDXDNf8PrhKgiD9eOy3Zr2q5+/y1nNyXwABNEwKZwUJ9YCNpTaCXsf
R2mHxFVrY5YmVmUOiy093xbxO3FGR/KKHyMjLdvfbPkVnx/uA8ZUT2YiUbxbe2l2
keRTwRXmXpp2KknB1j7JnYLvzj+6huzc8p2ZLOLLkpA8oMqrTy7Nj9eEsnVB/axS
j1zUlYnWcjzxxx9k6wG6MDMYawJyJvC1m8qdJhaNPMtLsgOtvLyyMAV6uAr2boz6
UIhtIbTcSoeZjdkGtgizmFUt+Da8XkTwclUOeYHTKJdPq2c4Mbjlzk0wpD3+G+e7
dwD4YcaEJxPTrsu4ET8SI+ymM+5+ZDnTHbSp5AZaU0CbPVJMfapgEcHIg/4+imYL
UYtEfiWfpvkjhEDWebEKR9CVOmVcUbX5ML9Eerd8mAJTIlwrhtyqAQ/0D0jWpVpU
VBqFgBwytRho+R6dq6rRa2Cn++4hd6HsZ74gvnQGZX4Le7ZKd2RsNGB8L5loYAtF
xC7c7NvjerDOC+CjJtGdA6B5pUyYLL3QiZ695tAg1pW5amdREd7Hdk5waI8TZxQs
8ZN0nscmcZ5GIe8zhK4nB9ywLwuTRI3rOhAC9D9LipvTyR7XZHfsIfWFrLYlMCAd
DKZem1zNgkfUViE6BIkVft/DS/PJvQQiYzNOdKWncQqbX3FxL9z2LvbpQzuFWcJp
ghqI9WXIDpKpDtgHWLrKZY96B6zmCT2paYc7T3Oe9LipXNPVNMSvIOvaaWSDCdCJ
NPoEf5vIxdr0jZwmGOnhfJgQrZBG2pV8pIY9+6qa3oSYRVKLRb77UMC9pRI8lwQD
Y9yfxyjKqIcjlCei3q22lag2Sa5XqUgqQEjZWl2TnJTji9UnCCyyY6RTWbHsN90r
oOetRBB9pfMDz0OjFVGnVrI/sHyNEgVWwgFjbYnCphSmRad0/jvAcEv+34Fqnw6J
oT6O8NnwcT6FzgJdyWLi70yqi4qmMgynI6j+P3NTDlNQhIQI2zrdamvEdjOuTmIm
Y9vuJik8pU/gbZAc1Dofe0wAPIjJhF3b2sXVZ5+OGHUrOxDKBL2qksfLz2SmEiXS
VTvOzpkW9t18CtJbc+GHAg3Inaa4rKoRyL22w9fjjAa+1UkALLA/ulpEglzkwWcF
mWLBwPAXkoVErUG06GrXupmvjSk/6uWdSc/QRTjH/UmAEgQck+/NsKZiWOxvzJ3F
ajxyX3nA/Oj7XXroeVSlm3Hq0nf67rQP6YeezlzesshFNe1csGPzUbQwvv5UTFr8
61PcvN9pYJ7/zLH3o/PXfWdrE1KLIq2kLLpVQQTtm6q8hQSDF30hVssTY5aUjOh7
yzSqhwLySZUZTxO6uZc3gWemMliRq8j5LHvx7TiNNSDR0NuXbCQOF6S6DlzPIsE+
/mb7WvEDDJM+OB+Y8DpCBRL9Wc+ZjBffxmQBMZKfoXioczW/f0c20OwW0cz0kzRM
TL2HNM96UnsDvKZby7TXIeD6ojwGp+ZL4tKYmYUA190qcqnwHuAPsA+NPgp58Lp/
+jx/+sOC8oLxu8apkcBSI/cM6ohFRCgUDGauU7vsIQNB3jC37vNd96UbYhioVEk7
PTl/mkpGpcED3eIJWm3tKQfU3emwaps/mLw3UGg7Y/ePVYBIte8ZBSidLHSbzHxJ
T6KY+QLrlpLgqkbz+fbjf+W4tFbkhwqg3A+vEUAfG0xzMhl1/Cbh7F5dmlPgk47v
If71jvzG/NQM56xKKxKffmhv613D4p8/Rdj8HKo9UWb2mDL4S1I3xDcuz+DF+min
zeEMqK5IPggmMmpeWB28wvasgEbnxVPLPkAyoKM9eekixUflIXE23WfvFl2qd6Oc
Ncp40ECe/zGljZexoihjBn5bhUTcrMLrwByDFhOWS1prgvRsVl2PoSGwICRGA3PM
5XOXkA2Gayyrv81zK9/zwjFHWXwsZ7eVxVhT3prZNRphM9EzMjJ2sulCYS34ekhB
JYPu4AtMzJOZ9yXiutJsyFlh6TATmRbykURcuUThjDx4L8gMOi9UdiqCdMSJw4CD
N8odMezeaiiQF/f6NVQGIZy9ADcOOw2sn8bNYoa5NpVyYveI7MoNGWyIvAO0pWIS
1d97HHwE2nIowmdzE5Vnslk1l8AuS4Z/97J/duaFXuuxi3oQhg3YNBUiOivcaiWv
b1jf5ubnBboY7kGD0u4sq5nA8eHmc8AiPuGajOL6C95zaP27tyrRL1Rv3TV+GiWh
I3vMLBU4d8d8RtixSLlsmmFW7Bzlo3ZFXSm/u1x4Xt55Mr+FR4HHwCTeINtX5WIQ
8b82FnK4ZWTAkJxhUpK0O5T5uUoNocpxYikeWMKuRwjAqJO6HBx6BEpTg7GgoC7f
t7b5hKS5W8FSEtyWcpo/NmW4B/Sw66h17zyPgHA99nb20vYTX3QSdewr1ngKJ5S5
kFMKNxi5hnwOKk6TcpEpBvOnCLetzjZbUOwTnBnr2ShFT4Ah8VFtDgU/EtKfVfOA
ah4mkFBfiAz/ZUOzSnO+qG4kbILPlnsRkYxDG0zz6yiG6MNmHIVNQMl++t5o9/4H
q4IkCLNn4KrgwwPSDcxAydVjAvR7aq7Gveq2jKJXxu8b1XKoflcBW2S8h6KZnRzF
inHG2oENTtvNtJT+qvrKrphiTzD7KD6AACvRkbkhptZdaj6GBIDnY9qkbY7kbxur
98zY6tTWU70m6fDjnIwjSUdkTdGPHvJBnSQfKNcY+9pO8/oD8d+LvJ6ZTGT317CQ
zmC1GR1dALHKuh+DnBagP1HJw/14TIo7p09D7u61fQBRkgssViGyjPCxWcPohTRn
ScKBbC0mDcIQHrEEWmwOk795Jy+nR/c0ALAG8Mkq3dzfWyDbS6z+m+eHd+hXYJ5A
7KVp+QQY95fmxmIx0BBW7BSJYLNBBua1b+O6ENRM7yu79I2gZZMJAN9uxfvkdJeW
mOk+BYC2rMl1AKJj1FQYAXmuFEfWx7UYKS1cO684hV3RFZyjup+GgRUDSM/F4/k1
rNyneO89FUYmOS9u99W8NIuW6VIFWS0DLRdS6lmz8D12iXBeTVR2aeetReE2tk0h
GCOvHvf+uonADnQTB3xwaOs4aP++n/F6rWcRfC2jFU61u7JzdQjpqTnjYyQnAZjw
7tOmJ+h5iIPRIl03MjgJ4OlECzHF4WebGoGvJhYslMqFs59hG4nbtVKWPee2otH6
2uklX9rQgVI95wmNSiDJeuHbkfHaWcmylsDFVMipWvWHVq+9jnxs/B3vnrxHD4Oh
UABZg/1LVnIFzaIO/c+E5ZxrMU4ZHn+R+2GikgfSCJZXwe2cRwUvYR+0mQdPB7EV
39IGjQbmeeJYb1CIVoWkgYTEK6h3HMUGuuPHDuDnBXnMM1e8XL5Su54JY6R2aFvL
V7xPfT6zMh5Y11GpfONNKn3SDxD6rFMiDyiefo/NoCZMxa4Ma/otl/dUQLyqu/Mg
2UsyjJdhuY268q9bLzpQhLRltjQ28YLZbl2y1zwA9qaJdjAse7DUWj42JL1s2Sk1
c6gU5s0Me2uszsm3kspHCYKe076CjEU7VdFiVqG52qWw9umIA0jqd8FqCW3oobFq
kZc9a8OeL4ratKVDJ2muHJTf/nMgyl1XwbRFTHXYtGaePuzRL+kJ3PA/WirKQtEt
uCK94ZK/GTrewk3f0tjNR5YlY1yQCsM4gSgbXEgtKgBQhU7ATn18v5b7MGQ4+NCf
DEJyP4vCwWyUtSRr5oPcS+tiC6qD1O+GWruZZYXf/AwJbcT75QR5xVxm74qp6Ll8
RuoIyyQOix9DSblq4EwT3OLFeef+y5mZKZmAHAKorwPAtiXG0+9Zymj6eVtlBNKI
8+2euTOXauINeMW9XieggFxhVPAUhGdBYssyTvhN/6j6fHrq7ANZ4SdSzcEaEXLP
RuoRbGljVb+W8OLpudOb7WSGedz802XHuBRWTwAWWJ9MIXR613Idy/N1wCwdYjso
LRlL9G5llls9yLUF7Air1HiV6eLK+YmxBMI5nKINa5BJQbpYFx3VGd2nCATdWaju
a0zYW5TA7bMjTqK+X3m9qOLgAdkMKWHUAkmvgy8NYS9KHHpSeSblPvvg4bRp474r
0AIs4qL4Q8K9iAnoT1lu5oWcez0P42+crDtNSv+3AR1D0dKjqSEkI8OaE7SgkqJl
A8fm4DzO1MTCuo8s/97nVOjPQSeE8PBahX/aXfW+96bLNigMy2GKlRLHbgtdhJ3O
B5YvdmjjF4/Wt8ONot8LFz3Ptpv9BXgMur06U6ZEUoBeFihnGlV6CWtu0lvvnu9s
ryVAXYVtOTEbRT2a9ZNWQGpRj+Z0v+fvhf4pVApe/PvC6TBaxqopXCWtO1ywVUh5
40yIuEOrLt61qoepEQdnqqwFnHHJjs2nRQQX+sHlz+ZYOxMQtoeDTsQLdfXfFdMF
4pUhu2Uh1XMwvINJY54YoOOlx3gaB03O0cxV+4Od4ULC75xy/XrYA3vQ/8mUOf4G
FN6rTgx6klwTXTpItssdRndnlag1/S4KyxFEa8ULZ8QYoWOhdumMMZPgBO0hUtEB
+CL8sISmlGXXXT07UibJCSTeM5cvqTdGlPa6n/q5k6O66NMOEx7fb/ZkJWe5XMzD
YqCxT34c7o9gWzSm2xutWmesr7tEXRPAVe6wDAboiQAfVZeybJ45hv8y08R6awNa
7Ql7yerFY/1VsyyoqjQHUwJ3tQWfFXkmK0j/vVdiNvpZcRIYFCBaJ10Ou+6DG+L/
N/bPKBz897Lx+uxO1v/7mZfYJ7t7ig3Kvbf6XQjiQsQVpZkf5+HJEITANbcbZIDZ
V5VmyoRMV5MuNooFh1LwoQtJapfJKHsxIMyD6Vmrl3woIbtzAO1twPH3NTtyl87q
lkGGLBuBbKkX32VRBYwuly6WOGzJUCiVTsX7t8rJ66gjDm6X6luXRyafkwCNUpc6
uXvbQmG2WRMOPmhXc7J8ZhpQ8U0pAemrXiFUPI/7OD4al5QuB9XeJMqFDDx1J5bM
aF3hDx1BZHL4lAcZ6UqS0j047sv/hwSQRqjpo8b09ciJfocvZDjAohAgAlXoHIQQ
wU4LbdVl3N47Lxsppa5Na8jlkzvm7XIeSCq5UfdFyz+6APxSY8efi8o0dOlX2zZ5
+o3cysCzVbLz/JsZadm0Cr3KI6U7ncZ0Dvn3nxtt9bUUOWswSmTMHqy9UeBdDQ7a
xD+roAswNWj1YTHoQCB5ir/vP96M8iOgotfSWDiw3C7ug26Kf6gcV0CkWE963e7O
ReC02MJUs0B8cqdM1bWu7WT6QuJBLM3DaMMbXpiM6o8bK7UZJUIHpJKDEcCkZuHZ
4qggqx55JeVuUftkGufgMvERo2WEdV/87lf2UE37PFw1punwfrQEue0znu5yExPl
smpElcXNsc7DMbE3gIqh9c+jh5VRB8pDMNSATPYxLuHBqmDmCfNpxKKsVBbsTV5R
oLQ7fB3xzub9ZIg/+6UCYnwjv3+ElrtMGucyK7hn77+uJnJ+w+bW/RQ/Acm0s80/
uw7LwGsiga/Ow1goZs/8Q+mRjPMz3F5kgrPq4wfmywegpo/67Z/+M4tYx+rA/Kl8
8PimuyZ68V0DZOz/WynZ4CWLMqvOWQGrXETJi4GsYokA/rHyMMV8Bl5Z06byTsEi
Jl+63xFMG84x0OvHN6z7GT8ROAc9KX19vPOaFBBJrPa0g2T4tOFN7E8KII5lSM2y
1EDFf6on2DVefYG0YzJhmhk+I4fCRYCewytgQyWe8Guq7eFM04YLI88qj1UAn+T7
sDu1J0MZebNyCNcaV+xfDZjDdmm+E6vzGCMw3nuAtzNAi8OdTzStC0pf0x1yQKJS
LK/qloYKIxxtjJm7rsdqFPSrAjPnv0T/yyL5Znv9f3Z39TxPM0wmbAidp4ua8VRW
B0dRrfA18f/NB+MFNbN2+hf46852g5Ks7r3j/HphX6ESepjhw+RPG0OmUMX6cszz
MXBuPViSYo1HTq+OEGCPGi+E5KMk8SHd9N0RHYAX1Hha/l7lZHcRFzPt7dhszu9L
aj3cCR+aNGBVUU/f2KK3xX9VXDTVAGK1oorMo4o3SfjoBzmvd6MvOAY201OM8+48
cWcIEOTc9bYuNFb5hT6GsGbw6InXHJKROjicfl5MNv3z9IegBOE3p1oUQbQzBHaE
+i6yJfZBHeyRZ6JTFVqU2VWz2lgmpP2CULuHUPixwJF9snyRRy/y8ld4m9MVplYC
zHdsWWBDo6mCAvxZKt3IXTLCLPAA0N1I9/1mJh7mjeFvXr3nQ+YnSJR77MGRZBbA
1BnhUiBf03zEZeNKyKXtw73Fbg1a17Ahsng8oG1WMs6FenVxnMlbZTooYll0f95O
9yhxnWsAGplERa8cSfliYp2Y6ZsKxxWTvZfuli4EYpTaQhR/lfSQw6HfOHZZ4RP6
1pctLaXYJYGH2QCwOTDc1XYYZD8XDpyseqOCU7FdMBUIiceOK4nsZqeovyOakEOZ
xjY0wfVjaYjQ9nJAuMycjtyhI9KikvZzHq1xrmfPagQow+5b2dNNsJGaZIcfMgO5
fCSZY10FYRDrV/7eINor8Et4+gzwMjVV9HQp2o9+lixv6Tz/HwBA4tNZaOz1BQvr
QAgC88MXyUwsYs+u3gOVzF5ieOtp9KUMvuW3IfMqF3rdGL94ldApOBUoFnPTYePB
bwcxurfd+N7JCIFQb8qpw59ihyahPD+C5k4vGtjoyBCf3LpzvnphiL3/9VIhTWhu
TPrkS0ngWSulfFoVQrBBEaP6mmjHJvqSz8FsVwpqYvuS+xnLR9rrhtYS5O3r+7+T
8PT4OOdjlKJPNOBwJzWKN65+H9B4B0DpKrMMu6lkqgdnhHEjQlPJrW5y0tpVJIqQ
31UEBg2EyK8KCG5F7HLDWeJKOJwSiKxlA+IgCogOyWPjAB2XZYqXmwnT5ioVTLtl
39BZt66ccaFjgD7FnGqY113cbaC5eQ03pbpmWdLKKIWcqNswH2gFVw8hrcP0zTFD
8Y9AAYpxslPQCeAM/sDtYbvTmKp8qoXfrJrAeyIToP7nb3b0/XDN6nD/665cbJ5v
lW6cKW10ZZrg+sdeGT0aYUywUoG9VB3DY/NjP0VjA3utjCN+mQnfDQdJhRpAmsS/
AwHzgKyNKYQlUhQ4iM/M1zwUv6ZxtJDBjVC0zpTYz3YrdUDkRMEapvWaiZqQOTdT
hVLnOm+erd6sRCoRZbDbGBMIVTWjPUOAkOUvbGgaSxhACHXczQaLz27LW/t4xvXT
s9Zm09akp+xbBNewhe6EdSkNAK/WB/azxDdI3UZh3+xuntdXn2aQSsASiWQz5cX0
qpkKuaKqv0nBqE0Jwxerqy9Cati/Art0rNV8iJJyeSL29q0wZ63lFlnZRYFcsHzt
smzQgBcdPHJZG7Iw9EytOsbIuAdlE2+GkuLYf11nfL1y79Rf8ck3RaNbPJ9wDJ5/
nhKNpmbAxLJJIJY2h40TU/vqPT02mYYGFeMPmArp/z1rbbKfMje6enKZOA9V5mbI
U4k5paT6K4HU/WKDeGqjGwZeok0fwh2c6siwVkEy1387dLQJ61tmvRpjix+6w1Py
q7rX8lhIsAGWTpIqoHrvQtwp3O9/9T9a1MWzSxyVPT/bU7G5J8x+lLchimYhbyDG
WM1r5r4jwmyq57Vw3sPjLGD9iVxgKSOvaiMXNExxC5YqOYBLaAlN8V01JedxjsSB
nciPqVQYKcLKSASb+i6b0sgjDzMcgBtY1ge8qvczf+nZrZP0MXHJeyOXC9HvNfgN
iqqzl98nRjeNJpFJ+iZlt6EfXozu06ZxZyce+rSa99HkSHO6rjqnMLeK28ErEV36
ekQDCFj6opZAg4GPK/6aZhWM3tYu7JD7BLweqXcjVqIj0frjb7LL92CIEOjDoweS
Qm3DdqmMctksBQc77kRdFEsbXriO/JGeaqzgA+h7l0m2k83h8LcrTC25TLv/Xn/W
pRQ7MTYwwWvZ6RDh/ku7Rh50nh0S50lB6uPcDrJeHHGonv5OGb1SQtmzxHvnSmyn
sCpjzNdXYRa5Q8A6ZaID2tllTjOwwvYHYyq17Oel9kgITQXruaOd9+6vIXG1/pxY
H80vGebrzGX6om42OR7xq8buSOPw++djzk/R5wNk4Dc/6daJLh1weg6LZLp4RLBO
TCDrmlGk4KKTwVoqjinZmpwwS+zMuSI0JPMelCL0tg2EB7ck4SGECL/2Io2cayre
SGYC3KFGHfMhw1IdHgILwB+j30zFwgUDFjhHQlwx8rpqd64FOlb1hv+3HUbBxA83
FZjUz+faVjXrCiMCHa8/rJ0l0j7RS4TZXNBRbVokyZBWEFWD34Iit5RJZ8kYFNFl
xt4yL6lAK5VPrAyE2BlMw6zRT6U/6A3V0IJd6VR7kyUt9Yazlt39+5Pc3hIumAf5
MHDtWcVmhRd8vqal+uC3G9ZZ6U47lLJSXS62vBgYObYaYViKIjPo+Qh2S0KDOEYY
5G5JyeaZ3iev3t3y+bPKF6+4nZaBVt3bArsrWYTb58JjzEIZlj2p7lBPOkHkkPfp
HD9nuY6MgtGz5uqmj8ROPrmSKYTP8wkgO2E2nfWZ5HMlTpsG9ynCtGudqfEb+NCJ
Hu0JzrTv5HDVy7iHIWbwaTrikzH+MScefGHSmYrN+RCGqm0t16o5Uc9q9BOczLTs
3ZCotBuv/e70D8AfifjCkFBuKozPI9BDGXZxBdt7z127IxZvY38tgVkP37z0z72C
bLzCBuqqk9gvWpz+w8t0tJRPP4fv3DrH6giqGlnISisaNhTP6OKa4uVKx2myESBC
MCgMK2VWIfxyORCP+R1knKodAAUbi+BM7OiBwPIpu3uolwFOr84d0URMMQMIecCS
ubz5R5WZhmnGZOrUWXGpKikiNXhLPUBbewSIowORSULrOR89BSFOn1+UrPzRk6Cl
LwxCH3uQZpLl0LoObwvg/JmsE/naIX3ORcuT+BHEpMz5+yg54rE3nLFLA5TPE6SL
BQKosIzmzKsx1ogbctPjsJ1ANNrRtdal6rQyCFEDM3rV2FNPQaOwGxtoBJXOrF80
P0Mw4J165YMQlZikYllwQxdyHYNco0m0YE5A0f56YxIsPW1Bk5Tgx2trtSUeiCaE
2uXNtMcy40MzdzyKtLfq+zYEzPJ8Ijut+wunaOxCX2WAlFP4Iio0JnyAIpiNMeWU
ci9QFGL+3d6av0lqFt80VJukBA4O5bHyjkzZ5ghWqUPGTQWQeG8JmOSljvzv1egC
/lEV50xwyBZFdb2UA/yfXrPwywTwwtPwHDch5x/o7B6Gh/OObTKb0+j04NTip03x
Fd5CH1dIZ1OI0ylfLTSxLb4aWOGkQzzuj4YtmHFz7chW4MeMMxHaPyWIUSRQHnU3
vq+DoOB5aKsIRcO1YohrtUQIShQK1a2FVSlWd28jFK8PbINkHzrSXKtcuNYm2nqr
rIxSo9jgGrC3urFn7Jj3CKmVIO/6SuOklkPns56S4FQSScdAZEbx9QIspqMAU61k
ApKXK/tPaKNF/4Bit1gZIffjZ/187EyfO46WTaMPv/P0T3ZWmGBixjC2ycsDS7C+
oN50AWicW9m4up4ETOoAHz0a0qKzh1wZBVXCQRsppRLtt6fuLZTR6kzDBnscn+Ue
gFEYXycCgYXEZhEEE5JYEatVtnIkdnSjp5RUSzUz2ToWwACfHW3h2oY5nOv+WGRD
NmxF0jm/RNC9SQ/VKERDHtlI8hNSOkNg/3ZPFy9c1yd0DKNAPZQvf/s8CUtxaKLg
rJGjrLMpgCFcoWVjy51GXY5EdbRnfjA7iFISdestKEGIuVATGL7ecqei5lxbE85F
SvPeQqmYGEXvX4gNJqonQ5Z5ZJQdVt6AmTgX8z9UZifPXpZo3KtjsHTbEH5rer6p
v34PrWMhxR334Di/2+97bBQOSpOfhYlFJBycPRkwADw7Vp4TzQya75JNJP6MWk2Y
fhg3dX8mO7sMjmt7iIPGFtCfOjqPGGWKtygv/jWK/x2wVp7f3F1LjAWJP8rvuU7t
sxiiuVn9oPyZb018ezxbHa++7Yxu8MYfW0EnauOGhm18j10QCtWHdZ6g96IItG4a
T3pQEqiOU0EkqQPmo/SRRTQsJNhYo6h7rloAXDFCYf1O54loe1sTrdmwhFhs/Q4v
KhG26jjlPYeaAJoaMZfY3+RtIZ5INciPG9VxW+UpboF2ZJISdhtYIX6XlEmreSey
UVTqxrRdamObhq9ZZ9rG4e2rz4gJJnvi/TKT0w8cyIPYXPdOVjbbQRuvE28iWQi9
I0M+dtVw/YgTSh/PZPOLDcmoViurv60+KAGb1d2Yel6UEYSRqCT+/QzSVIwp+Kno
PVFV9+YpSsvKhvAPIJi81Nqz66/KoHvOe4S/Vm3SQxOMQrqJZ6nGt1yacPhRO2Rc
/GjCsihpDM7UupErUR0p36KKZn7hZRI+CDYujTGGIeyzsZmyTwDSeHmHyrmW3S/6
yT2a6XOZCBaRHWo9CGOOb+KJ4+cUxXdQsj4TSoXovlX7v0Te0HBcsuB5UI1oRSW0
Mh2v2K7nPErvRYT299IXih420i/QxS31OcvPNRodVYcbZGd77rjxbZy4DbVW9lR7
4e6l1OkrvRNurr9TrxSgzKtYGCl8B0xd2O2BTUbDvepUSr0nPmZGtvV2bF4lQkHW
lY1BIzj/MiPZqtOBPBubNoi0BnL0aA2X623zgkRh2roqDAaL7nHDuJn+qTXH5xOq
M455bGiznRWemv5A05nFQFmmxqOu7QGhe76yo7InlN6qO82w0sQI/Pn3VjJaBfkd
XvYHINP8ThMySazP8rHMRPBxEsl7qVPHXAkNiYtD5/ORB7t8dXZadhifysCtlhDN
DRNRd7SfaMPol2k4amAV7V+RZYCg3AizbGP0PwvyBjZsQ1w1blza5UaAWK1E2LS6
7ru6EicVRbll8FlamymtTxtOWyzVFx8bE9upUU2Xa7Nh/bIcsZVsKeUOqDsVQ/jF
B2qHk7ez5LshDTY68evyptx5eadJA0TPaJYQ8RYjPw7L0cAV3kI+nd7qzNh/yT6s
O7270ScizzmehIPUXR8HrGXop+i7bHukEL3jHWJPieRRJ5XVqh+ybPPBzFbAgJts
0/1tx11z9AcERMbk0+Q7jJMkFtrCzPL+oWnbHPyljdVNSzH4Cp6YXKqgGwNFF6XX
y61OmApceoRFJb7s0M+22PNUxNnvpajfz7+hksPjgjl6jwSjKibsZ7k5wjeD0GX0
/3vSP5R70wB1Uu1dRg14i0u6bpZJ9+aLjxCW0/wqHBkPjmRZfChcJR2wL8q1DF2h
Y21CQfsbxS7HAVrdCxd7r/h8VhfF4pHrmLAth8HkEAn2A1Uup56nNDudzyDNhNwr
ulXnVTUOniajz2pQ19SdtOSwJY3do6JbEvEQGMSYfEWF2Egtv9Uh0oZKEvtdOd0Y
4cfLkmaiFPfub6fIqOpMY/T/hdx56bEXG8gSDvQGTWiIKDvk7nTaKsrJx84kMNSd
AnN9JOHC1I5n41nQhaF9pG2AfIq5pVNKraV4zSODbZqaPViC4NnuTXEnnF8gyBHm
Nz5PD+7HkJSTgyN4RZ4OYI1uUVagx9FXUQ/StzgGHxgXfu0hta5G19ctkXkGr6hK
HLrr27NGMVlzzVkRAAWNaptTkIWYpGXkbTfGRYnPcadMM+cFgs+8SS0dgwXg+boN
H3Walr/MGBs8DLu+mshQkyG2xk0g5eY/MYMUKWk38m9W8coOYnXgQeTL2GxNbFie
3XwMP0iuN/XMfsoQ8+wzGfI55r/wxtH2BphL/AouvktuemAhyd/yfnDnVwQlxvyV
toRjYy4Mick6wkIhLbk2WDzlye0CjtD7rSW8L8hK4zEg7cWYM0X7T1DkwxVmYGwP
Lhk/lV7868i58lEPxceLXUuGEXZZMX8FNU/DSsoTgnhxCeV3toUVSE4SbeQOO6yE
45h0Q10Vy/PptgZoN4MiSpNyyG4YEAiImcq2h1hIA/FmcRT5/2CmPysg72aDUn9Y
VvcR6UG1RPZEdY+zH18C0ilsqrLL7TfPmfMSFMs3J8qbL0merauHGB7vphxUvQru
CHblwMbMfH33KmVDDOzg/qlWd2eo8akpyxNHZwFEqisrSkghOxlgKNP3S2HTZGMK
zr/CE7YsyLN9robGoroG/0GwLnx2QqlUR34exw5JM47pHwJSVU/bmkEfXI9VuhYt
BmrM3+HAYycYzDMq0H2ovd8nRTUd4PGwCr/MefCzZBvlH8W4bW8IWZHTkLMTaEbh
cxkFF5amMDgLdbwNdqwZJajStnT7gZkfyBmC1e+wTDRWTr7kNVtrgv1FJLFN6ld8
pvP328chwoIDU52tDGKhZ2MxhNtIpJ9oFxoKY8pIxG0bBjp70IqwJPnAoTYID2oF
wffh8I2eP0Q1U+fSIW9Vj1rtZUoxjKQgb0HIo+1HTexG4OFtn5FNK4ShanlZGLQB
J206dlRiTsjRfyc2MBT92nKPOS5MdLGRqL0N4Hd62TtwpNcPh1qIMPH7EXTX8t15
8XHV8sOq4B8eI2ZHXS0ObvALjsbZnfqyG4ido6Ff5BvJVPZHSev/SCSdbZgoSGFF
5zxfLAhcxKDDmZCkTBqMoM7VElNxKqhbahfqDmzABbXbeShuKZU7RZ/FKTrtPpdY
PXTIU40nG5Qr6TflwkHPUsYY/Cm+oAm5dmiN/PKHq2ebXUkLEqMGx888iXvoMWmW
cZ/20vyK+aZAx89tYWj5nEE0C7LJ/rP8exq8W83S9EsR5y89o+fbkXFXXyTp/OiS
ks16QG00pPviqkcUNm59NWYCxB1q1Hf6fT0wPAe6GFRDWskSH41kTI30eB5MB6Fp
otHPA9ycNa0bLvkmpshB/b4wJW6zwcyITqlcYJmQ++z9bqQJcS+Pc1zZr6pMbMh9
YFwTPyXnVf4p7Bcq6u9X5dL1yPaxP9qFGg1Y6VYmaHVNa45Gueq1iyUrJioTBvdV
6GzbnJNM9NsAndLU1MCXPy56FPgoHimxAvFDP7uy6UIbHbcAjuZm1IlIVTB+ZLv0
napRX1HTYMD7gZzI+VlX9oDdDhi08SP5fcuQty1Hx0cgzurrbdmY27n08lGMdaYG
C4tIYROy9QkS2E7pJd99qGpIzaUj9jn52KoEATkKwaRvKHcwATddhNUo3JPL4qcn
Rop4TcjxcRK4BLRqJz+ldYq03ZSxenhiOLGyAY48gIlts5UKn3k7ggFLFEXy/BP1
/aKTuRqfhXehPMpkpapTog6L4oSQD1my0hnw2WSLkXjK1ANT5zRGLtP3fDajbBFw
pzhaIazDqViNd7qBO2Muyh/OuBitdCQvp2MSDxSYFqvw8A9uGSCg1INKeiL97BUt
Vqwss42mszZVyQFMIQkilIzP3wHZtQ9Sr78Rs0aXxn5Hdjgci91jxf8e9H8aDQi7
u/WVcKbPum+YuNr+jONNRR0rMSRVAQ7dp2/kXDBy723Xlr/Mzj824PC1JoTnAYpa
uWtB9yin2gPfCouByyM1BcmTPKUVLvT9lL6H36LJRTgiwWftzHS40k0ekh8QEosI
EkxdnbIXS3v95PyrYaTpdeKM4BoU2BebD5OVzpzAaJuk4qjcnuaY6bbMao8OaFi5
teo8EZExWZYWwSIWEUIQC4wUurSAl5VAG10nCxrqk4rvwGaN+jQEWboiCaY2sV+6
JHAMb6AY34y/UkzDmwbydLWqT5IR5yb7wiFHmgXFYFIQlrjyigjDcxr9m24Yo+7V
Ywp/rOjXG6WB++V6dqyFR6osQWNsHFNQ+MFYEfsiLoMhhopeIBBlaem6ustDUGvW
YeE8ufWbhVrGsxYuaFy26/SvDPGESnwflNYtq3h+JQApvrp8pnxkF3hxcv0yVD30
7ZrLAYzZ3NsS/qLQeIiyc/Mef5lN+h4KkoISCh6Df47CPiu0QgFRkWKaJudZL4eW
4FPbeM7OR/rnft9k7cEghGL3FZfABb6vF4wDYc2O8v1v2tgdGilds+1ZVoDgTJ1M
D+2V5Ry3oyyl/DOzVNEAPdTTvqBXRtNDy8x9Uvc8c5ujXWlCQMvtafxHJQjUrMdC
dl173xk4nEGxPDrVKEJBkRXEu7D6BxK/wR7EYr8fj9KJf/yWNCOXF5zBCnSUC6Xe
I+nWOMC4wGIjIOpk28Yj4OJJTnmMpqaBvgxHMyjyk25MXcQIpDe40fi9/A0GnieN
JJSBOe/8GSmEJjHo8AMg5PmKR5AMKrb/8S3xsQhE/j24PWVBK5ro/EZIHxfmC1vS
wP8lKUy49YHINjFTNsqu9BvR8+l0djeXM3TTDrfjWvGujbCUqaF21aLdAKwVdBlS
DkBwu7lO6f5y3P5N2woRfp8gTnEbKjVyDqhmEAYmAHRNRYS9+WpRcpNqxmNKJzur
WOww94YvPNwMUVlnSZfWXBMVoQu8OTUSqlFlA5qSuDYgWQREgwbx5hpkUNsbH8a9
gS0v5GoAOV8o/ovubOTfF7ahG9vgw+8luPI9oabrvBlsfRAW+nwTOtRnSapRQDe7
isWopyJaRm43l174pVGExYFxww3eVhhPogj5DFYztpHy54lM3guXntEp8Iv3YuQq
wH1QPdhaN6Z8SEV6lXi0SMJAd7cfd47yDxaNQYpkLSNoGRC55qkl4XZoaYfLRQBT
86qcgvGNMtqw83kERQc74yGCP562HZwGPEMkvffdK/u7h/OCP9i8IE3/ibDH9+Rt
9zqO+VyUA99nm49wh+7zU5Jk2WWlWXZRQhGWFSELzNkAk0h1/DG/J74ykCjGDkqB
j7bQCcucKBwiXM2d1zxU9vzBZSHQTpRneB/wFMNnV469wdt+jk1OQbg/mUQHDsgX
k9IWEaJXhEPajdHWfxJbswLLn7Fj2uer8kfTqia4KaDGkq4gbCyuloMuHutHCdig
hlve0OvNqij7FdZb74JLhNiJiHadMRo30NVHlcbNXTanrGOEi6zVqKkpqosBInkI
3ZO3g7o8m0oHctTIec7yBIOwXCrEHeLEhYeJv1k8e7Z5+0N7EJF4CvM7+kUGf/X3
6J/ukiO0yP6lq290GeIV+cVsHo8iKshMDdoByhZsTI1XUb3U970uwLJtSevASsI8
nw8jQ4SDY6PelmNKZQ7+5gpTsE7dZibDH75s/QMhfS6rJMEOoWktCD8cc6H4nQ1q
s/g83N2kLZVHcJYWJrDzYghsWUpMMAQ49t2MW202etLzAejROQ+qvbDEYmbEUXke
uh+lhJmPQumGMabS+kLXjvZQZxvvO5qY87rRVXn8JDGzNTlNlPqNbxXi+9ucsZIU
QjslSH7bC7TYFWoqzYrv57xfFqhfzwivJMtMVLNbySMGKduGse1Onw1nwnaiGH9k
BA/os8AiprK+qUwKTW2SPY+y5yz0pyYDsESm2JqbxXGR969PCjKqjKwkYQ+4IkcZ
o/bJ6LVHfNbPd5I11oKd+izrTDVvU7X2LwQru5mkQcEe48UW+MtFg3LZ5CB6Vtwa
UNlzJZWYFuQOC+84JJioR3erxaI4q/85ZlSteaETJBdkglRw3rx/vYryhqiXezyk
TSNDaZGpPi7CUrUIwqpHIM7LEfmPikfLQ4tgrNhFrbOjiH/tg3Phm0vC35pYJ81w
cQLKrxHV2dzqsHb+T6+wPARrNvfC2mjO4eYT7iYj6Mowfh8YSddD6TgSb0kvDQk4
ZW4dC6TwyBZtqAdUy2+rQukuLeQzKgFKjzcLlkwOZvLOaqQvxL4b3gNi7TBuHEVn
YHBjdrWRyU+oik/6VwAADhid4dpbu63cC48jPVeyxiJFfzvHlcnI+Tp+r2iUAMv9
xg6uULtocoGkDnxVYW2zC8Gb46FoaRHWf4ylLN6McWNccGLnecf3s14imFvYvUc/
YeyB9J8dEaKu0f8FM8gfdOGKBtsl6+5C9MZPGpSwrbg92sEQgJJuahYKPdc1Z/x0
zchiDyAV475hx4E3qYYjd/JGPANQygrYWmBRM0us40kJQgaUbEbLrgxchfzq3wrv
HnZ8dz+aeUqDL4c8CzcogyrViA4Bt303XjnjDWFAWJi+AoZwoBS4YMn9NZlNjtvb
efX7p8buG54bfuqkYzlQBsLS3hhQ99Wcfp3FlBh4aeYDmWyC44VEAZ/qhur1JGGn
/anAHJdyDtQ5UK/TSjv0tpY8m0jNn9WPZsF5b43mUfwKP9mWzsoGN+I4pDYdva/z
KwlLGsJG7VwQ4SKVWhH9yl7Fkh3WP8cp+kDCjs6besYYPuwVONsu8991lHGf5EiJ
nhKpeuTS+0jAG1xNDCMmEh5U4ADl6t4Jlc3wUS3bEUEoRGBn0D/7F3DLfQ5NNd1S
qAtUP1muGuct5sAhbxhsK2Qzk4DWcVQf1wJL4Cxl5auO23GrwEMOMgFy1B3c/gy/
IMHO3a/ppsrtcOHgxAVIBLm4C6n91Q7hx3ho0jtexfkloWUoxxzxVfn8kG6YoQF+
tpzhP/Jn2wRQ4h4WxM8EHoobfwCndeAOTKsYKcICk4McbIQn8lzBLdiXL3BDLvb6
/JBMqQeuOUV8sfiohyJHR+CK2pOXYYsxLUNjczCwK9xgntTx0uHZ0XXRUbWfQDWX
sGMp1uPbw3G+b9II1fLtqi4PIE1KWR6632bpYg65GX8R7WNCYMwKZdLwo5UfwhRq
j4RBmUSosP6RgE1+OdkAoGuY+CSiCel5oLSIMe5i/5ajYgnuLQ4RUNFf+hABDXOJ
0sCwPODiw7uuMw8ezCsriHuYcYLdSRtAdRiDaieeEnCXv08bGE+4O0oIL+kz6zrS
tHzLCps+yz7HPHQUtUnT+M9wRywf3ALp0+fti8pUlCOQ/DNptHph4dV/tX58D693
oX3N03dXrIriAm+KuOuGuQ0zepuk26wA0WmTXZdrx6lcpZyPnsqrFR7VdL0kPMl3
dRSG58/RXOHk0NtATt3r0cSx2veJ0OwvX1xHNURHSEXuRYyCg7na876STeM+s9N7
Zq+AIaj7zNI94OOK3xCBqU+kY8Cns9tEMbJGojK4cA9Djx0Smfc9YkXrovW+s+Mg
ihOVuzs0PTYgF/ffz74y3wuvFuro91MvKAIeEq2LR9TldOSJHddR3RsmPmx1GaGN
WAcgFYpWhqw+g8rjiidkViorh5edBD5Yi5uDisfgYsdA9VitZ9Vtjgbrg05GjgGc
vh5JCse3QmolkB5w0apOL39CoaNb30LPXBep5gM+a2FGNiCKZCiyUS+Qda82aVMV
Lp/1gyqsxaPrIbv5pAov1/lM6YoUrB19Xdczac+DcuxIYhngHhmr10ZSigMwMETD
pwaUbZhEooOXXcweT444KvHJuWbdvHoTctH+ctUG6gThrVl0+GoDJMCujD915u2n
svm8fcAlW3vbei0Iu9XFIkcKnYhNDD0ozIEzczEKaUeYHuf835qz2P5PRkXYIde4
0iloKi6ELro9HzkwqnvwKyhqbnfIJuBY2NWYkMAZGtHACN4EqeyvjPTjkJERl8qu
Me+lO4Y6M/5otS6tG6tinfNSM0c7y8YPPxKCuUtdcfGay8nImLbbXXwUOuZpZHwZ
o4eB7aRmV5qzAPlK3r7wSkPqPgI5QjmBP7/v50vs8EYInJIPYf11xTTnS94oRfmC
EUNPUyaJJM0wAdjYDsex17KpOWe6A5L0JEQlj0LygCLDjQHdL7P4sd0mgCEwwz0e
BGp0iACWAonOcSM7L/1anuABsi0M/DM6La0+OAWo3h/CAHBX7ZyyVkY1rTjyluyM
Y61bk1XebbQAZglMI19Blky40Mwa7WFgYo/ThOWoiiD9JpkpHCYwQ0dGpTdheq+y
UWHbaGbQBXCGdZpPZuAkmSc9+/FUHiyEHgJPKC+nG9gkIBvnYBwlqQ3EPvJNii61
92d8Zqh4gdlvKghQd9bNmivb6oJ9HBFZoTygGN7Sjy9PD05bRwHiqkGA13B+H35y
9zGZJT8VpVLuq1NjsqONE5SKAld9uTkWqsQK0+HODzy5nTSjT6PNeE9dOkmMyPIE
EsKIKYmlWHN06wiP0huNIxaOMhreLZL14RL3TEXNYfaN37/GTigq+VuhxH8p599q
9kUfnS9Gtua9ALsA6ER2dC3kno94pX2cBaSLnnamnQ/+Yo5KOmif6e4lBdXN+7MT
EImS9WWqQ6014DHjanMiXarwR+P9ozlkwXpNpSdrvV2pmEEAiO9p2aSaaq5VmQAX
/qc2l23JJ4JLbYELdrt9xo6qPTb4/Ulgwu1Nd33wJT+YMuNc4/RDj4iHhz31i5Xz
qgRQL398bTKiwrQ9TVmsq2x9+chcNSWJN8j9e4G5uZKg3Bvvfm74Ar3MoP/K5Oyy
TRuczYE7747tyEoEiEtrFdC83QV2Opm8SGnyNhTc/InNa8AgS+JxxA97NcrGQ8Y7
pnHd/s5qi0ZNvtMjjh5EbySfIKwadI1f40TCVY0UI6MoWI+z2UYPGWguP/R8KmYF
NY3IjSQe5/zyttsSvbzPYpRV28KKkxWUpF3nI8cP3J2QuYt4kVBf3rU7Ycv1v1HD
cX/hY0O/3maO3cgewpi4XtyGrUrj4MozW+MXRh+Gvzj9n3sOD50rzy8p7b5/QVeI
xIo4wVJxl7HhtSVerdttAzOpYkMWINMBSL1Mi26XuPj5QSpZVMdkCJQAjGQriSnk
q1ssk0gh3fWIUwSxO6CKJVPYSK6nkS+lDEoSFbUmhrKx8xyLmfVxY7Qulbw1ZDO2
0YeKm1l/4S3Q0NOCtPIbYF70doxM53Jq5yAiXzLeS6KfjxqOtERSonDec5oZWchK
r2OyJZm/S7CMs8x657bK18KCxU8Lq27oir6sFsg492RvyU5U78NoXXs9DFuVeOeN
Uz9eQgXG+SArkEfgcRdFbl4vV4boQGSvJgNZ3BCWEEPtUQlm+uig1nTUNArSg6lA
KB86YrBlkWirXeNmQPFpy5rlz66dNXebabpM88z7lrxEm1CA190UfDsSAPfBC1o5
EJUNoObQY5fbZimZLXNW26qCU29qZgcA3ANfBSeBrCAWO7kAySQWIRccgzN7f7Bc
CU4OUGQ2I5KtZw/4SAhfELezLqtIIrTE0Ndov6VBvK3IiOQEML15FhgpLHL8gFtN
U/HfsmdUZwaYT2KbIgaqV3cE+GRjKa2ItZ4KlzTaGWviDpr7+epfCm/dJAlICI/4
PAuFe+bJgPL+sR6hSXsDePVCjvbyUGUuO0PIjQ6JwKhlOUDIrUCKMsbw54m8tblf
9GeYd9GSnoIzAD3E2TRezDvMjmX3W7cJRNm8VLBWvxWHIQ90LGmehVVsdR4VeLRU
poIybKSbj3HhdhHYMlgIFMxOek5ESHODjmQ/XYhGcgf6w7bN9kHlMI88pj39J2CO
94zs1IktvOj47gQMfLDcGDeguTo2GIVNq9QDzn1IwyznubUkQrfvD+YxY8PRg6D2
S/oohYZhDQoMF09gKWx5CuGM5CYRysc3T8/z2pgphp+1nSiA0ejInqYNDDdAWeXF
fAeLk/Wqp99bazXlXEzx5LZJnJoanq9W+M0y1i3N+zUzAsik+2lMEw8Vz+/jk6jI
y5drVCvTzqVRXMakyW1sghnEvcoLH0y8fRjBnT+SnWw4HgU1gVD+EId+j53lY3H1
hbhCIfKCAhlJtekgsxU+ZNRK5NFavQDoym80J7d/qob+R6h/bIa73Z7pFtUvuNF/
Nv8q5iyMYKB8yK/7o3dN8txNvb59kBoruzL7knjzEbFCGP3prj8QI927MKZV/LrL
8wJIDwidxRL+s3mmE4sPVzTYecur4YbF4NE7y4Flafo7TRXGtsLCzmiujp91iD+K
Z9pV/qjj1NYi2W3Kie8V9Q8zRIVlqNs0MdLTFH6a4GzyZuj5gLaXkYmE3ThFS7NM
oWIfSCpnD2sSzmY8xcCxObCz2FHdAfeaJgQNeLZmx/Gt1hi4Q4ttqBjtrshd3LO8
0vcuBQg9nGKaPEbnCWBqxR8dj9KAGv1nKq8pOH+zEC3x8M1/QNi4P9/Vpwwypt6b
CKjS4eeRLuA2E5ozU4CJJDybTCOddddOI7et4Qt2/MlDgYrAsuIJxSCP7waRbUC6
AUtJOVLj3AshHMChHakkPVAe/QyGTpxEiZ86Mlye0m+uS2s/AOM4+jn0/IgnwGBx
SRPoSSSchCOmM9NnjRwHLOwu5ukvpROnKyLeEDe27x6a400hBtZqWRGJfwgDUyuJ
AX82AyPCujqpZ9S2E3XOSPD9sLoPLgtD7rDJOHgHmk2/o7EfRnYr7JIYCF2dIlbh
Y7q+SRqTYTCQaXwCbhclwCAaAWUtODWHpbVyp0jNvWNDFmIKKjK5HeclyCD5pKvO
QORBXIcV5ZTTnLyjWJeJMoHbRX29dwubrZpa2XY1Z+4yvMmmBuxwfU1wS1plYukF
LtnQLJJcmiS+z9OAi4TRsqHj+cRAwq2CNDbKj/BCuVUYl67p7eejqzds8Cy4j9Pe
deQRl0NEET3S5VsIroi6zyvWjhfCP4R4XuA9SIdm811a/U2T53K8L9/nMXSzRBfT
UTohsj60d3tipBAO/Nlb5mzUALPjXEcIgi5P+d1sSRG9WlHvgR5+HoiqOE9QF+DG
9pxaSjksyAnQL/LrqBoIYbuTJkiTqZBO4sUGBKfAKE5blY+2QJeJiDI8FmmQ8e6X
w6ENocUhyOfgUf9neNlwqS+u54B3zqYDlfse+G8g6d4UvqxjbBRsAuYW2rCtyj9/
vMhJMbmQkn2KsxOG7XtfZRcw5j1pCnwLTNCZKH5ZqndFJ7otRGOKMVlaAESBqt7C
H8js1La0AB2VLUGnh1jny8+H+W7Ta9qVShWjp805voyFhAtuKIEtxMGH8nLdmyvw
+p9Dp9YzWviS/n6CnQADgVJGH/q07azYLyqZtMOIXxVZY1rlwqEk3KL+ZGXuGOa1
LEFY20C0oN3r92lQzcadCGuI/4CQ00v/QvsWfII3qVvpPnQC0K3N290Oa2Yq0jtC
SAadulbsGwuHsNWM8Skkry7SS4qaCvWaxvZgOGNGfZxwwqvA2F2kx8VMPNnxombh
xCoyQ1Dh2ZDfVJhaYm8B9MQgr9DMhkzqS0G7d2BtXWMWLED8ey9pYZXq+xwc3ZMx
8FtxQ8Z7anQ4XyBIEsp2heHKH29Yk9OyyaMUL6Mkql92+kpTiIgyZEdAJIM47cyH
mwqziphlAncWgvLjK/vuG+tYhvlSWI+aVz9Bkir3WGC2Qzq6+E6ULW7RBqU0YkMD
zY+I0xmT0M5VgxVxi9CDANoVcjurrckcZSy5KDBbiTdBLQuRMYzeyNrQot7UAZWx
6LmsBGMS340BHae79jV/N3z3PVE2Mmjb8343m+xkdVbwCqWlW/z36q5/BZHdwA66
Iwh9pOWEJainUjDm1SJwWq/snU+FHm4Z9EtE2w6HJDuTY/eSTBJ3pD73uBCN1Dc7
4j5g1dw1mGJpMszNlwsr2kO7ZIlHSmI86hDepms8qefN05U59N4iXs/2CZEDxGi5
ioKWEqO+1J2dCcyaKAa3S0rDDrE8G3NUGmgzebtknwEZN9v6LTiVJeXFvuBSMmnx
CaS6nzP40SDBl6xqnlFslQ0d74TwJCELECCL4MJyBgsn6l0dPf5c+z94Ndk8LXRE
h2RdIDPxFf8YJoIc3YO+6hbwjc5oVSKGSWdd4EPAXLnvvP+weVFiAQuTTp9BXvWt
3N1MwTort/+rofYJ/4S+k8zXp/A03XJrBCrpZU64lBMA8eXK1QsjgARe2f2Bv2rx
XZNTHx9clFuHhW16vDF5GtaKBnK2dhxEz2g2Hup0BzKtpzXRI8KdrJ0E0rpQf1hf
mQ0hU4SKzZF0hrxIGeaTt7vmwqRcZtxDy9FocFlWwG4WGuJuDbYUn3LYK7uQnSKT
tZUiEP5OIaD1qOUUVy9j/Tm4JIZ2zfdLy94hhDJPjQVQyKV+n1JvCkMz57Ezy44X
0T0Xq2qTxAij5EyYZJei2zr0Fqkus7NcDdVQm8x4S5BxQVmMXxpZfa3jejDGKuJU
XTR3YScbgQ4Ovsc1q+WsXnFMJTtx2pZN4yvQCQ4SpCk6YyZju2StSx4anTcWbMPh
MfK2H0qdxfJNYD8tJ0FeF5xXo1WkIaSaroO/7a17Ngm9JDvWBdA4T7DgNJUZvEEn
xpkl27jLPPUQ1aSSflQoGG4DmUgsT3zPTSnm07uYwILk0eW3VxXMfOZzX3sgw+gg
MTmCY0sh2PE+HOFSwJJN7QOpAmwpamHPvF2JVKiuX0YiRWxiSkw2+PiOcKRZuPMs
lzsiRY+Y5pxlyDeYbL+U015rwqFOYYHSH1wYFmewXIBfFz62pDLNw8L+q+Adexe4
lqb12cSorevIJTfOxsv77OGzPZsA1OyNmXLrSa9tWGbh0PrlvY3V9TJBDSQSFvML
wnycy1GLuo23qJaOa2m0VckmzOcNTtg8DgJH1anBY7mF6gdmnuUTlswAgKKDuub1
2F2o6UIrSfki2lhPLFgCgoXULHDOVURfk8T0mSfB8tPfi4BaWAZomXmzqLSGhY2g
vrVytrvXIonQ8JqRrzGDe2+KXU6fx5kQfBw5w0+dVYZ+XpOSvZ2AFpmxgDoQP9P5
C/EpOw7JW8pzXvqxykT8ateFzX/CUTpQqzSu+lPqWsJIs0lSmeDQyyS/2lMghWqJ
yrpIEUgvbUioSd3znOz5PM/Iazq1PD5G68ce/CLQfJFZqogabhcc3ha2uBxGYYFd
n/p67PeBBa/7dCfZI0CIi19URoisM1wjlSTbke35LnhDoEiM0KKrPX38Wl9Q1Tc7
8QUEo6PzcwFSjd3Yd2U8VZu2Or4cjwA1mkeKDS36CrOpD5djyOvHnV19Nj445Jp4
LEapnRRpv6VITiGz2ZpVt1RcrXY1kXv9xP4WgNDuPXRv2xHtxrfrszanAtE4iNty
w3W+XwcAcuvKeM/xh7220SJoIm3ALB1907pz3BIUBA3rMHv0KR/8D1D1UvvI84ry
X2DhGntGQgLrXqPTMTCvk9/oNHf5e1U7I3Twh/TqTYPiKBHR225Uv9d4ZSkJIYZY
X1aQuw0ra/3HxX/+Wmh4RAgexyju2js2b+JuEN0wfni16kBB9gi97AJPXi0v91wX
Qd/rIEjLwgHNKzTrzOSlzwbKmYPnhZC0fBq8YxsaQtkWF+gFxC6EcmgdbD0gM2AO
lou4EsQMb1OSJifgtUskPAzSvkUYAcLfCCxOUWc2UEoeJYoU+CLqInFK+Em2SyCg
46ryHJPqIVH/EpteA8C92D0KNjTW8SkkM++LHcmGZ7lh3wldM4v+Eq2gyzQf9TzH
EATOnbrIp2fJEsZ6Tt9Jx+/fWQAU9OvLPEJCqHn14knV5+oAHHCODlyYE+9hVy/7
sonO96dftU5esyOe5sYjlyCCqvA3TeOFmKc2lsaDV2TmYnPBlYG89csaj4BSeXoX
4LlPH5Y1tXycx11hMAPUh6P7/46Z25e5bCsivXN5/OqIlUaoVbSz4xVqS7tfSu/d
yuaOXvIjMGeBfMj93wP95HRixU5+Mea2pav9pnAOpTxl35Iio8MeCL9f1rcomxy/
NshLGqPINUhIVpM6PiD+LODS3MgCCvtVXSzZxQ/ZaCSRFG8UXKzv5jLCMKeOYEHp
s9OrSEu733Gi6+O9QEFKxPp01IWRMcc3IzKrelJS3h2vGlhIXEVhzxTCMV4BInaq
b1XPp0ful/Jpws5tUZiN9/7RUpnM3731jDkmSyuU30HHsNNk8BVaLAvdkfhA1MVr
98kz/UMK2hmYYSJiq//msvLC7EmmblO5iYC3fmTomRAWQMYm2m2bGstF7SnHvlk0
hwOm0uoDregeQ2/mbt3E5MgqXmrP14I6LFBRek3vncIuimJsnHp+51zyxm5WxE9S
skIm6DlLCfyVWDBUL26lZHfzZleEx1F6HoplkRVVdt3q+tZHeGjF+0E5QYYJfECi
JGkKqoBbx0xNyc2xX40x50ScDDqFbTDOEkrJC2GZyAUlgIFpAvB/g71tGene3c3N
vN3GyFRUx4JExuW4bp0ukc7/OUGAVXj7h+J9ulusEYvFNufgbHyAX+dDostVjj/2
ZvSk4m+dyzlr9r0YFs0Sb4YK+EP4yVY62/BS2Bvm4HItQtGzZAHvkqNRwUPOvDpm
CI4BbgqsCn16iVBwd8n0hi61O53Odgu9RB6P4blRwbw8vtfHyythjGXrSz+5apjC
rFD7wQ/2LIqylsNvdIM/zL7fNCnidD512YnF9fjNsnBQqKWpm5Q2rE9t+WSconJ7
04hxDgAnWhnpWLyu+eToIMM9NF1VykchTYQ8JAA1OHx29hE/aNmvJeEp8wdZkGxc
M3e42Qu1ubiM7HHogXNhgoZsKF2SobtbZDfsEDKxa3MMlJ86lULrJVAz4fizatxb
NLUG5J0ZXPiA4N9NZZa6GDIdC/2wVQDfM3XQ4r/mcvWLRc+BPmo/vXUgQ/DTdEHj
1fp2Bq5kbfvAiGONWVUkoR8YIQPKtGfsrpLxXKNM7cCLAHEBBvFgUc4IyIA6Xw5Y
2EZw3vJbR8bIYzVUrmzXLs787ws9gjdUn9sXItZaTKN6ukdfDmHYJe3JZh/KXPU4
2fPU/AY8FQtzXYxptC5XHyvPSh8ed5NAJ97FtyyJTQLOntTbd9pj11bXfFou3LQR
BH7xeqCFdM06zlmpaVMPyA6mEIMKul5ftWpDf4lRxXcTiXOkb7gVCtVqbDR0j8Nw
6EZ7CARTTllt+hrga3csB3eUfTr1LW4mUrc+3XYkpVxgpQxBOBGxmACkhzMClnv8
yNolnOul5Ps2+2p6LFWSwiZX66odin0QfQ1JTuZVJ49BFL3x+IQg8GHFRJtg3RRU
V+nopGa23J5BI348KmgFEF6AWns4+peyMeU8Ju6FIvMI9HoKa6MiDffDUA2HeaPu
bW4CeKWScw6zRijtf5f+fycQ5MBiw8ZLOtiES99aPIrshT2WSllwjFl8MOivMHT2
jueQn7b/pst/JtF0jKLQ8RkBYmdw9ey37D6QJuv3kRJp+2UmQV2KIrc1OTuQiggh
5LuTNK80l2NsijXEuEqYkIC8WY1gz7A0bSaKtpmj590e+KISHbTXV5RwRaTkwLSU
o8i4KqSdTaoh9ADP4L12oSbKAH2al9+3nhIuaSEcpvBToNl/1Y7UX4aEupKaf5a5
+/kxqSt9GVdK+WbqL2VUo0MNaaUQjUr5f4GSlpj8D4WwrPmd0rYpcsLEBobvnxej
T0rW9mYbiujO6oRGWEPKK5jIpuPzGvm4zkL3gxmNctnVkUK9L6TXikv+fVFaiK3a
5W2sDPt/s4SAB6cTrDNa6OUb1ZhkinzPj7yBqgc22oiiZ2j+d0jM/t/TVhavsrN9
W9OcobJGmldLBPvB2fs20QpxSQyNZiK6zncjj32S7G3NNxhSBsdAISGL7RQneY3N
E+YUwPYrnkf9ecGH8QgJtFwOUopnkex6xTQOFo1kUKQT5LmU5rZiD/yYTM583Gam
+rlXcbnwEZJF969f1Z99OrWKFX9CrwO0wIDx+ODxpUl6eRF21THasIV0MVNKF6JJ
xi77s0ONNmiAfLh7ABXNd+/MgtdDvrMd0zUFVHcz3o6XpnXxAyoAdns03zINQz/k
TPPAYOMVZSM43Abn3wA7zJIUYxL7h5mA1boP2T4qiwCVCG7DdQbBqbLjq9eEdUSg
3aY+fNN87TJIplcBbDgoIJYqJ1pfD20H9/FRQrHE70JLUsfEh39Kgo3As5d299xO
mGF1YVGOt05ZZDy+3q2pCjh1RwwS3eg0zmt5az05eMlb3LOrZM8z1GAN//fiWhKF
Fdb9OPDzjtd+sy5GzZ0XQa6he9+yOTKaLDwPhAreICtt3luafZxhvRY1CpEl5o5N
K5zTYGbxkmWrVA64AFleceiroZ4X4AKbajkKfgsoLePDfbJMR2yMFrPgwdiSUqjn
KTD8G7h13RZ4B38bhvOYaRTTQQlbRKmTWwh7KtqxbY9yBA1zaFc0Vh6/4W7jjdc6
ibVSTQxOfPJcfy9EYWJlArbjEkrq9WHfadkTxCoOnE8S/yV0b+XyPnEBLAdohHAg
zyjg7LYKII33TZp5Xb8HE2B92GBliXGDxVGkBK+Qt00V2lCvkPGKdIkE7GgKBrA4
bRdgNjac/NMa1ZRJAwQsw4sAJgI38GVV8j625R/a5HOXooPHNvtOdH1jiV4i8j33
esfp4zDx2ukugR5Fgf6yB+d5Dz4xRWSbd8kt4ckOx6oWzYhpr31nVNaB4PdtRXhN
tfOgqyZ/sOI8JFz5Aeyw7QAYOf3SnRzir07DGvVIvZOwyodK8DUR8SkKZk5zQxtS
i6JKxM4SH7t/4p/IK5RUh1kNU55kmaosoA0dEUh6873zohJQRgagtdHqkUMu0b/I
+1rAbp7Imtcd3X4fdIuUrnm4PQ2uzT47vawc+EGO0F0MHDw1pmSZwaQyGDVCPIVH
nVruK4H36i5+EUQObp3z/BsnennznpNVKW7Qvw9ftXJmYJHu7w4zgiS/vQG7+kSf
75jpmyC5aHV+f2AEYjZi2DFJr9lQ5LND1Qkv//QilSgF/cqfAQQA/nMBUk06dhHp
1AQgaCpGWHJo3g+wI4rKg4le5nvCgna/zkVls0L3IGanUcIm55Q6T1f2I2mJewpv
qYcndCXA3DextNv8T4SAC/gr2/jo9xfNgM5G7Wb2LCWNDTtkaY606dgdQp88wl0h
yfEhYBSHsBRwOtuAYfenF14AMAfgpvjoew/Nu1/hbQGjESEffG0+8dIZtoCvMlM9
+Bo2BXc0pKW6iKc+1T8nuQ7Wa4saerzms60I7xH6juD87BmS+ye4gUg6x15NZcjP
gdM2WYTNecSaBlDqD4pMj+I5LHDUYCT91uGyHWQe7mxy8HsXnI2nOLel1kn86/O2
dpKpKuoHOW69GE2OgiLVoF6rj7tYwXYCtfvowPqyIbxzP5JbX35WG/7ZuNrtpt2D
oEYANFZg3oeBPPbDV3DclFrdPjoQUlgOda3PGqOsLB/XRGBPDuiKEDZfgsDeQT4z
2s02kKSED952/PcIii8BcYWeEeDWYGK8LHo1rXf5A+0kzpO0h5yFfebVOU6PlLYf
Q9uFgJhJLRkuRQ2ZKbemZUhc4mQ4M3xKMV5vaVQDYLhU4oIKVqbopG7B+55Y4rNK
PbsoaqhuWTc2TlHeIBsA024LGtOQrfz3VkEzbtaXg0O1zN5xD2kl+9jVbnnqU0a3
/vw0u+Fij2P6MZlFlM23y5mpjGIqG2jJKwpVJAsTzcAC3Xf8IY0niGneeZMLqf8p
jCk/3NxY+ORsf2cMg+RVuZSv3qDchgoDAC7qXqXd/dQ6+5HQ0QXdq6Twe6oO/4I0
vPh80KD3Y/nZA4vAUkgW5W0c/aLZZTXtOG2MjobJ+RdCX/qgQz5nMImmUJaHgImL
D0ukHBvPkbOsTmMhE9KX3igiDJzL0NTCTqcmx8cj2t3Ldy3R31Y0tg7jE/GaeS7f
Ezb0KUHJE+hbS9tWu6WkhMd9RbmIZYIif4urAPh9KfmNCGbGyChr7byvB3hqL17D
PUAair/uq0vGo4zkIHNt7Sp/+hPY1Bla5p2QZtlu2yPpReSYIyymOW9k7UKvE4YR
rKFnjzrl/1W8cGWQl9E5KSpzJ0M6vwycjuQmKo/60DpoX+rYuUHGKEEP799F8+bP
Fy6WQ6Qvkd25skWcMEJKE4Ov2/vm4j87tnTAc8fUdoNeatPVm9ka6Y5uq8Vg009p
aPphVL2/J/3d+rawGaitjiGkncH/376s2b9f5XE/K2dLrmjQ804C8PEp07LiM1Gn
Ew1HNpwDtk77KQ31ZE+rAVZFPLZGJvwUXSTnetAdl+qPyQ9+5Gxd8TUdXEcx069d
ti+vFMhxZEZjCSK/oCL5dOYjZSR3E0Ayl+eTEG6k4UxJmXN7/lLpOtV8xyZw9Kpp
QX6VsereoKeQw281sRh/jQGhMfUN6zYjcuJOyXz6v3y3APUvM+HPwLEEfEF/1GV5
0jQc2ENGg/GzgLsoDHa1nRBHSB52r0JBQg6Q0gnVQfxIWEGZ3sTUAQz9tzbL9X04
QdsQya4sbn6qg7udOvzek0X2dMJdxjKi4gEDwbWTNK5DaxmWRIlT/hkRpvVnGcs5
ZR13EckK5tQHH+oOhjWFAF8j1rmuNRKF/NVgKjYytYqOk/mYCwuBqoLc56lC4ylZ
Cs9TTvPoPOmH9b4mkFiA74JX7CjydIghMWCSWAtKYr+K/k1SHifXJR7HZWe495BU
lY98QEVVp5YYJzjtJyX6d2SlXkWKzhWbzilIFmZzNqACLCdhAvTAA6cC4lJRPbSb
qiU8fdHVXuKOkpuXK74PcUBnC4P4OPhpH6QPw5Y7g9nW+EDdWZRQOVvECVlN84ld
MBppts7ciJlpOTjlRty0En98yO5mems4qfuQuVSv/Dzzqku/YR+6jO7I/cwuafMF
yRdnaE18WBkq+ZG9hI5s8W43/FQMluWw9hUNK2w+MyMbV0Kw/UMNRjRh9Jt+VFnT
aJZM7Has9pkXLerz49vVJm3yRqB+2rwCsmIeT4EJT2rZf9NCjp4V0qGCrucPnBch
G/TvAx8iCbpre2rrnJL1uz9PnsFI3PToc1g32WcOprSy0Vuc5U6vrdRDuRvr/3jC
2FjW99eSt6+wCMCA8rDI+mcUWP+mAcwq7rWPCgcNhJDRLDUryla4q3yKeYwR5+eX
6QcknbXyJXvBLrhmMcqKYBanB6B7YCK3w6s5xGEQH8E/GIqdOCktjWzbBxCNwCFx
cMWsFQMH7YLSVvZVrHvUa7hB4GDR/3vUxRYqiwdF01W04bnDdqit1fv/qIq3sTlx
aU82m2Cvha9jH4LsyOoB16sT1YZG8OQzhXpo14BTMM0UQOGlfS5mJNTuLa6VVGyG
45/8IBzVdK1zkYQHSMG1XJ2LScvrf3Pt3jE6UW1l4ATmhrqxbEYWsZH00gVlPiZi
uTXJ9u7gTXm7b0oYZeNopAPn6+TYrjlYiPFGvLn2BtiU8bB7e7hyzSa7ch1oNEjW
8zShJpsSVTnVHQ8hU6Yyp5eHw/2vCUs2EOOGRfue22MSRMNdvuouaPD1RtvlfpdG
GTuwGREXPbGH4jGDU+O8yFMrOBMHhnmu3qx3Ynf+nCoIBF3fJ5wr0sm13NIXnp6v
TF+bSIomgjC5HEzBb/UK+dN6SoVQoaVSW+AvPbOjE7CSaMcPoZSieOxsfobJJN+H
qx1fLkpN+vjHLIicZ7yCJYKA55ME1MRyb4GWpltua3hkqesBHjERvFfQCha3hBZQ
z/fdA2YMcNTul/inil6tS67A/JGFgfyT0snfE+T1j8oUs0gIdneLlAL9mBt8NIem
3bKjFCFjqaHufybd9WBS3xIXc/K/Bws/FYSggIe6xGNF6+bb6Stub87pEoAIkHhD
M1WGVJkMo3qJdv9y69CuA8bhxnCF/i22cFz7z+DPexnIMxM5Q43CY4tMPu0mLYRt
LGAf1bO4CLMR6WSnmkjoYI5m8v8B+2rt0Z2ANC/6qksYoqQQ/uGYROMhXlwHKrjG
8El66Ezmpi1iqMPIKK/eLPJcy2lWGZhsJvZeOUd8vcefWVIuzI7ieXrEVeceJ3/L
YT9D171QnALKARvvPlZu+OJbXR+Bff+HAjmVI/QOCH1iR7RwYUt9MVv2j586le85
RinY1LacmsWd6aPW8W55jWj7bDhI6ljnua4124e+SPNAX6MeRruDr4QGNTjz+xqh
5VeHVydo/QgKf+Vba3ukHdrk9+lLrr2kUj9u1ah69xkKJn6cVE5OxYx44XCBZ2ti
jxsrSb0+z5RHuR5NRF2me1XqDYoFyjZ3qS2OCywWB9TnTifM1wlVy6D+I03qZVJ6
kGW0+0x/4WhFZGbiRNZ7gMiX9tCR1IOcQqHgpPHW386jknciEtYyy2yrkWG8t6YX
sq7IilRcyjWTlhyCNJvkfovF4lj19lhfi6nrdLGWReZCv6lFOC3MsNr8O0NmNU5e
w3D05OswX3oEFvz2ScqiParlwEQE7QbIG66zv0aQmeBc20eFfnmpaXfXtMrk/xnw
EImlIh526w6b8MfYJd789lJaycl7vJxp6qzBs37jdBN2lcEkF0rloeZ1idTaDnK4
XVPblTj3pqJR3d+LPFhAKZo3azFBB9mDfBUNns4pTp+33yPv9Q48cG17JbMkhTS5
TI+vsX0HRcAlGI/QGEwfDQo2nEsrYR2zdG06hNp0u5JRhvZE4NAuY9e+UG7um7dn
kdErlugGYd+tWx3NrtgbuVzK1j9qctflOAqwLZ9S1ub8I+atA7av6S3nNf9cyZGD
eoUhIpV3jqDJFEQ9VP/1fX2w+LMZnDNI9sLiSUAP12dWemT6K7pFghH4e56vasJU
U2m7FhvCie1pkqHi4BWWU+tjM3rU9BoNL2z+1PmHoZvpGDLmpkNxV7joKQS0NSl2
L4dKZklzaBCe+PaxzecvQG+E7fCFFnDkmz/1MOSPskCAvADVAL3qeoUaHg5//vCb
h066Cd3Ii4VKtwaGRyAMcrkVKc4KelCRha1HrluTcK4lf63P6qqHU9QRb/2z1MBz
ovuHtZgmr6MzHRj3PvAc8U/cJRdh7wOtBiMXG2fKmLHSEPR/ohyP0TcXxh40H724
x0e2GiJDwblCs9zS6j4SO78AjkurAeZxZNtJoNJyD6efdoIjl6jo7k7qLhx2yz1A
5vPasbOy1W2LNPxq1cQMJr77GNhNLs2SqXZnKrDBzkCABKzlUHRnWcah7RTa+i8Q
3RlbS9oGtZjiRg5D5oqv7as2/OTywbnVTFPG4WC/lqtD9KNon+xoNlu9ZMOaV8Ql
V0+UIGkNN1+GpvzEDsRz5rZr5r/xaGzcdGyneiGvPhl7naHKK0Tt1m4b2CaAKQSa
PWdXNIzPe3TVucdGOiBzf4J9g5BURr4VXxXAOzvBu71r9dIHIrqkSaXmd0R0JYH2
feLE8Gj5AaEirb8R46/fNhIP/hti/F0py1dMUgjgLvPNq2IcQK9ew77vcNvp7WfF
doxG7zgxalFAaRIOK1J66/bvywbDu0mCsxc7jWKkhB5GN9nfbMoNHIP3hFttSzNj
rQVOYc9KMMBkUi6q2OEMyR7I78Ni4odjoaQk0JgrZh3FHIeyAvCoCDaQbz9raPw1
QTW2jJ3kJfAKBkUp1GfIxefA2mb+b1xA4R9pri5xxIz/s3OwY3lzl6lR3bOhJbZ2
FFEYnRt52AfaxJZT/i1Z+yvBwIxkUsYmAzpQCjRpHsAo202x+HX8NcJYWRb0jzqO
GieotaSOrw4sxC7GoKygJ1gbccPx6euHXdmG8TW1Bf6Pn6Z6HQB15BwXBsQqqJ0j
l4PoTq78HOwjPWVLOcRyYQwYpu1lk9c9bzrR3MCepSAf1wOQVAGyqzz8sfJ0cTYw
SP5517aIV15eGVg6vpLwMVnncE+3NEnysFPMyxav8Iqz0vSrf7PTI9BXnDgGF8BG
gqfQO346Ix1ajEXCs4nuJD91aGv+UtlLRgSKhbdkbKS9CKhfdcD90RE8uLCuwTE1
sF93wEq9LsrTuXu8zhxtbvcjxdz3JbXN3nu5cwRNOxUgWWr2dZwh5WbSbhP7LtOo
cViuq9k6X6B0wz5ADRJD8AHMBLy4JgmnA+Bq6bRDd6mY8lXflJPshOmYMAnNfM3o
IBzMnvjtHiuyVJpxHcF3D8u9XNx9wCMII3WZIZvHvhfcLugW/66or9iX9JKNCdet
twLypI6FAX/ypod/k4OTbuA1miJdOWtqb7Fu0tGFzsN4pakUNZvMRKOJTyz1AAuC
1A3Mu37UsfgoN9peAkEHpDDzrPY/cCX2a04ER19COG5a3rAf/wwO1JQ4RVvCXRjT
PhYltReD+5kAQEhwOmW8aenAjyJX6TXQbJNZrvAJv/6u3SSCQm+AETf7sxWIBW6g
vSqz6VLiG0VgFM4saoUu/pT25H6alVYhlOBsh/aM5dOPa5ZChTrgojb1RDZBgps8
gtBWaYr67epL9pSipOCVpVVg/lYM8JRzrFgsaFsKjaviR6dY9uyKIQave8JdjF0S
kjd1vs0SOILBjwVGjaPHujHHaFipgR7eVV5sLhQ4+vVep5Iw5cKxpOGhM6B5iugw
KIPosGdz1Tsyp/A7DO8xoDXC2y/4INO+2X9uJUfj8uNetCgzQ5/k25HQv9QREPx4
UURwE5K2PP3B3Z+He3LR5urWzwk+0Ifh1Pml70mP0F53yShDbLHlZtqzk898hz6y
MxrCehxl+23+7Ce/CqhjZSW2r3BN1hxo975bhc+0dYOolF6Uc/bl34Eap+Kq8rQk
L0ctHvqvPyef2nJLYV4dUY2ZuNDEGxgv3ZrMzNmxaCD5TkkwfQA8aWqjV2HtuaIN
rNH+OiyDhUTnqfVQQHCOkj+AYXzzD1HSIWFjgW+jiost5Z3TTO8Qt5s0gAib0WAe
zLA99/LI2FWbIM8+Aw0Ydl+jWOKDZ68RmxLSxu7yIU2tQsMIT0U1bFH2wcG3Q0Ae
7c/CuGvJ/Fn2lhNORBgN9dnbmO1JWZdivTsNGAfULiimwg4C6nonwrOIBrBS86tI
K2qgxCWMG+/dnq18YMhQsb1z9LyuhSvGiTDCROJAlbWVPHqhGzeWevsTpKHK23vq
GoBrQ4eBQqzHWVb7b6JDyuLYLEP8p4jnI4Xam6a4R98QU+3aNm6Yf5Ny0nhyvSfD
hQT4S7LRkp/hzBf2ycSfrGrX2b4nUQr6il+lYTDOXB28XdqIMLqzEhFjjmdlrJZ+
tDZnX7RPgg0vtNeJD/TJD+CKcKhRKfvLnXhjc6kgESdSZbh4UM1g9lhLTVs+eBYr
eqcBEeh4/0cD3y3+TE1656tckr88qOKIEri1RNJoxJMEIoDvALuOaA6WzRdE0/8Q
AN4i+Xt05GOyLpHwCwB9X9xk6tcypU6CQCQPZlIk4CKI7MYI3Vnvhc4Z0ucWbF7u
O8ExSCP7FoHmvvrRYguRYNzroeDfm8dM1iCx3IOR0Hldfb4S0HiWXz8qNoO1oqzh
LicO/5N8wMgq1FvboVR+YhVKyJiSJVMBpML3MEmfPBIxrqAEbp5hGW2ZxvjELFEQ
h032IurFrKdGm3KVWJ0XRQFJHWlqtX0SMT4vddIlXsKsRaIBDZwZzk2bVgw/+gr5
MWCpXt55N1/5iFGlzaOUrxyaOf5Mo4iGINqpMa8rYTNp81Li1NTnEoicKxvGA9qJ
tadwvS2fF/A/TSBNN78T8SAjIxd872tw/cVhEI+sELWueoxPUJEM+b8gcW6nk+a1
DwyRkMz3iHc0xlcvsC6Pq8qCkj8uKdwoXWp//rrQ3ll7kRc+nno38jVMco/hciWR
hKuKNW0/hRsIOm6lAKxaeTWS4w/2huTWb8+7ElyrLSnL2ozpPP5OGmMv9zzV5lYF
t3T9SL+PeqbnzDVtH0x9cp6DDQv5R2ZydoVsaI2jr1BAq829EGzWcTbOtRGW1fR/
/J/4BHQux9HVIsuLEy1sSqMZZwd03B1QDV1N28M1AtLYHXRTPLNa0XANVPwAZHJZ
hFvyidvDzHVKOLw0sE7P2K+r11uck4Dh+ym82/07VLTRos9MOgSnKgPFF9iC2UUe
Dde9BnFhhJhMfog76VPbSpnzX/b3PoUEQfpZbGCrlZ6ZmUfuC6SnWYZBiYvjGWM8
5p0Q5i4dDfDDLfMYh6Wk9uI7ue+l8ePkDJ2V6ly4TbSDdnWh8yCNyKA8zWH6SLUP
yGjSN2/sXtPyWpXOxzaO1sJDrxVygnCtDBpSUsBrB2YYxh/SCB/GihLkCRaR0ofh
BGQZZMcr0pjT35sMwu9d7BIz6m5gh8bGIohbctU2Qp1Gw6RhgfCRLer9WfpxgcSh
MuZ6HOeCrZO79PNZRPf8E9feCn5Yaw3zBQkTDNvzWGWoauMhr+TaO96OgQysPdLf
rfvhjRY/WTDrR1IrzQEQ4J/Xh1F4QoNKPgE4AVQqFG2ay0w45806GQ2SHumMACm2
jnKymH7LtUmOUTrAqOIBzJgyLCWek+g3UzuFAR/ZYoHClOirh+P5667cW41WuoEb
BUtHtRX2cja4IAkCxCb0kMcvsBeNLPR8iWqK1mEaa4Tdo9gSXanj1UcWsu23lYV0
e3kH+WTrA+cUws5PWapl9+PPiHIOWtoqtFS4fT6d1CxcYu+9IFCyTQP/DcBfH/MU
VUQL7wx9J0xYx+aPpdZJfzEruFdfvyyZ5LI8nn2oE5j8jsAFtBAWwcNeNN1lHnxV
Ia0IC2x/ajIyDUy4syKvnXFCT+4e4qmK824oOSkiNzbulo4PxzhCXR8dZYQz4hwE
zVp5/b7cNkQJLzJ/9lsEP4ltvLrXAJrON8Cui/c+T43cMr6stNejxfoli8cg2hae
av3BSDALYSGPeg7ar+JJcgtJn9zcn0AByR+2s0fQQ0NB0O4ZbDwJdeP1W5r8Kyf9
t5QSEzertoWtpq0alzvkamu6e+aWbGYgXEth5UWX6kdC22zXWaQMBI5QS0lKaMix
cwRNm88uLddHJhfcS0HF1qK7wgrl8hR+NuOjseDqQhYQzNC57ftmSGMUo6sL3rdL
tljcVzdFssCZCW41aLAstf8YCITYoS4woz+/dbSDFQD84O6uhdskejIim8gPz1ul
6S+t8ov03i80jID0l+VwYIvNjlF0nWAjSVqbwTp6xf+GnWTxS/o3e250+zAIjv8o
DUOhg3FuLCFB+RtliymKpitGogbLybCw4rf7Bckqc+OsD9POSGps3NiSzWhgbLDo
tjZ60SSDM83z1t+J+YCQ8NaYrSInieT6M2w1fIgWfeMHAasVCFB9sD9BV4lIKAco
M3zDZ6cXLJo+VOQZPVNGrBEfxwbS4YlxKe3OBjH1kojkJt4hqlIahT9l59Jw157C
6CjzVDLSyj3vB5MwTJ/YWooB288xT3WaGRIzsGsjK9/1byHYSfN7aI9Tud2+sVXK
Znm06bsRBE0pUdjwoChj4fhb/5YgfruKzC+VDaU9MeDuw7G7+wjxwSIGIyGH0rK7
eiX2KO9wIblOHG25lJmk5S2p7nidmiKAi4JGaVPx468NX/L21NH6ubN5lFviNIrV
TdiwbZKsW9fyXETdsoubc4b+k7i0fgvRBVNdip+3CcceqHZJlu5LewD9NqC4XIgp
iZ81ak8+zxGMW5dB8VQob7PgtjjuXje1OWSL0veFHhbLl23TiMSu+wj2yOVGgBlA
r0ImKhcKNcbCWsm9ilhmP/fhYPfQx08b6k9RwuuOzMRD/WLIEx+aI9W9ioh2aWAH
ycHzY9ExiMfIjNzWZdC8JCuF3iMAa6kDOQ0Eob4sfqUfH7cA1FyjqTtfLV6t/nz6
ASSKMWDFxvAdUaf848tXngwb5qKGLzBAtSxccEQlHColiut+UtpKWpKuo8gzPhtO
jWkVvBMMhbMStcj7w79MsKgLF9g24umR3+lHSS5rksLU/Hs+OoMQgFzdPpUDd+l8
uT1Cmwrk0eVUvNoV8TwihDWOc7tyQReWV8bmNcs6XOjrsU1FRZVvBTIIVAjX61AU
QnrUCBpLnzvToxIoqY42rcFZfnXtu3bQ0kktrqvCnBR5rYc/9dTwSngh9FcOKBda
/dfbBPukOG/OC1T98XkSVk3x+Wq8vb0ZHz1zU5qetlocT2guRnZgNeqwfm2/zxzI
E4QIxhbS71p+yWmW6wDEeWpjb9ZJd72AFad4DSvQ3paxj8jbEJ+tUzsxFIXdLZ/d
X2AQkdYAwzFeHDjJLJA6HODlkZsLK9kpVtFSGXCICut9WsqlDt5YVpw3DYsIEOb2
YZxX2RXaiZf1QKJyL8vm45gJYjOjA39cBlQhwJBYCruErThG6OViEjTjxajuo7H5
U26zLML/zjJyLhEspHf3lGPHvMHI7xY/8VzG0EOWijdOOYVF7VUFfO7jy4O5hIqX
CZ9dOU1k2FFPiZMpulNwf8AQnQ2nUFZ1uSN73Y6UvdbeFBEkCA3J2OlDrP1ZNHF3
xZynaIbMwWZsuA4t/ZEFkDD+6ohWg2hbMTrn3NoV3C5uI5baP81Vkirub4xLdn5V
GkZXG0TeetL8ylqGs+jVKA/UxdlXamYipeCOreOKIFMA/4H4c8wOQKj17999A3Nm
+y61l5yCz706cz+/KfF4DQUap1IkqFhbsvVUPCdBR5dGN6/W8ick68FrqfwZwl/+
3RymwAX09eFuQ5fhQh+8SxSOFQ7s9o1elDIcFpWI7W6QRsqrK1flvGL6KqBC9Tjn
VnYejusjj0pRXdqNN07nWogjuS42kJ7GfL5bTqWkENZRxd1dBuVK1c2A2774OvwF
d2Z6hr1KGlxl7Klvenfff5pEEomIDyPpd0xOC/oJf0gFGARLMxRIGX0+edIq2Lkx
elUGkTpqky/IrpuEuLPYx+/CF6lYlChYFA6RIahWCnkF7jghgrSSgFmq9s5KXvP1
wH8o7imgOoJsU6cbeIGItOEZtO6Tm+aktcrlJcB0NYnqslk1sVLx1gMBhSXbA6TL
W2h8hfVYXYUOYqZS6SGT1JZMrHBd90Y3n+xfAv6zbNK0+rKlRxj2cIt7s8OkGI8W
BsnbuSA5Dss91ajWFRYfAxzcMwzpWgdh9Qev+rwf3VBn1phxaagrwCziUE2kSsUf
JFsouU10ODE/LtCFpE5n43zvtiDZ77+PvUdcWJykNrPPb5Tjfabqqigmmjm3bpSD
ugfbANk+jROZ/0k4WrR5Gt7tmvuEY+5HjLkSzW04MA95z9jOUxrDNXbww76wfi5b
YQr7vFt6ogpwM428ecaiUVqDVcexOH12KWCQbEPkk14UOp4jFl98MXA6bhbA2/iN
oojKtdNiqlv3DI/DezpZFBCCA5RHvZz5HsDAq+BTWfzbrx+dji0AsaIxj/DiaFF5
6fAH+p8ViPozuv2Is5nTAvlQvR0RrS8xfMyej960h4XCTd3KXEvIJuvV7hKDXl0m
KFmhpylh721vRXgq3s19rQuTch8/PAx9rKqVU5P3IRLztBTzN38ncllyB0xds2Nt
t+Dfr65CjRGGtyqW6xmsAbVp6NiJMkGf2Qnr76lRNQyN0Fij4+nMkoI93S0x8UBp
yhyPpt9t83AnFyUSxtatMzLQRR5EucJADfvRFtbkzVeo6QZmcY5xnrDTFGa4N8iL
XjzTPi5tyc6fO7Lz72FYZrDgnN6naRQsVeet/zecbjHDAhkEoUpnjo9gopHDwBxF
FzYQeN96ofcZ3jZd7OD3jI5yNGus5gHw5tbY9n6jf0MrTuFp1IYC8kxEA3+HtiJF
SXNmmz+FQnyrL78MLEMYjLm1vfET9c3BmNVdVTcCjA7mt2LE8t/ycg+kWt15hUVK
v55LLA28KqPZPKnojQbdec39rj/mTvuqgBvu1SHQynnbllvCzdvLE+E2kyer6cOI
3xDACfBDcGlKvJ1CSgWlsbWIAIq8PYtnhn9EzuMppLjW3CPA5khi/cSyUv6sUAAn
iGcjt8k43jKBYAzR7KjPuf32ZcJdzY+WOsVD2Wzs/VY+F+v91HK7XQHgN5gltUSi
XhBNU/9vlQWhvoaHXVHTWOXVUqyAfBK3R+WRn+a/+9ZjTOhXjh5xJIUn5jwWQ69+
hmegmoPbrgkLRjcqsEmNfeqlFI/9r8XlkPlXGVPP75MrwTTvOF889YhY5PG7CZLS
shI4V6DDhGhXQfIimJxO6fbbO6CwEPzf+qsyJwflAqCkoyDcWeX9Jhkem81xqDBf
5J2smSl8glKkAZ8BO4+smXcVudYv1MvhvZRWEdamWGz66W5tSIqrsJ0Bd3x+VCez
tt2JhXZwYcp/H1gfPpWjpJ63cQnvrPgZu3zhN25MOCdi1sruJjj3PRRXJiQZy5I0
Y24L72qIwTdTJXy5PtleprSWepTL6T82IV3b5+CN5uOBcLLkjzl0agdMgPRw3mYh
aSw1iD5LBGRQYD/20jc0hgo3O7GMBGhuFL1sHVACKaPL0dJ/Cg7u3yBigsTwLdsH
4SEC0o64dYF+x3C/OF4ltLwPcT4QWUFKGMelzgdmbr1n0xHlvyO+Y8NogSg3v/6e
SIZ0Hz23cWMctqDIky0CMAvCM7LJjSwZ4YhyZNmmqJOvmoXXLHq872+fLHk/N7xE
2cljWcMllJWliwobIj62WbMGU2/TWeLlFTDpSlXtqTzTS44sC5uQ6u3CZDI/r9Iy
E2ct8Ha9E5I5cil1pY9N2FdVyGinZiTsZjIJoz54Byvk4Cir57ObTpUooYSYprTr
JSElCFjGQvgdvuEQlKUSs5nf4stSO7vxSskubLzKhjEhJMJ32ETTe55Ktr1RNJvN
8G7UAVxbnXanzFU2Wpdabm01Z1u/cZNZFxDbcy9+9BL9kw/sW89VmVaur5OV4qIb
WsaVb6py5XzJhb3R0iH+xnzrVCb1uOU8gqXX9a9K917aQWQkggINHm1wwR0SBFt5
cizrmP8o5EVYvOabRFOBd/TQV9IXQxXuD7Wu1iPtapsaXCoIEaGTNgk8turpRKYq
7OjWvGN1jIeGXNPBtLQOhn1Oh2ysXlGnA7Z6ok8i1dxd5QTfiU4z6U3AfMfeAKU6
iQrnr9fgtUPq1gL8kaifCuAL3naIlBbl+W0awkkTt6Ezs1++dxK8b0JFIy5qvZrT
qyoqgZ4VMmlykXbQgT2IYJUDZ7DhrqA4Vz57JrakK36yypXqRvL8qQPwUCv9exlG
3wGAey3osYEGpVP3ZaAEHdXSy5SQ5wcIKyXbOPTc0dnVBjVz2h/oU1vutaCWs1kv
q/bPHrUlN4A3WUG7jvLhO5Y7J4VBLzZ3msOrRxR4S/D0Cz5PuKOSla2/UJVV+/pl
caKuuNrMFqgkfjZ2VyGgsqnOLEzV+ofaF+DOBWcwbnODEIqRmWc1oeG0b54tsLIa
GrDID4pNjekL9UACD9dV2+bOHi+CNdMOGhsE4UlojKsGrWu0tQjT90QCmR+tWypM
fL3cAn6tZErAdehCXHzIzSRV/Ljleg3g9q16GEjBLxEHRJmxmAvtcckP+eu1X/EW
IQk3946zfZpGiKohIdAXAyBm0Hq8hQSEotGr8dBY9KPzdGFC9rMwQj9CkNYJMd+O
C1QFvGFozZiGx4ot9hcDU3YOdMAa57/a9+q9s7QbAcMsfX0AitJJllwpkiadXdKZ
`pragma protect end_protected
