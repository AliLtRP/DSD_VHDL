// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
L3I/R9FQ2EDjrYZKcHA7FG86diXCaM0usg+mlZgUXlwCsllRUc4Rku4zv83JNcfuYgsNyflEo5Sv
v66WXhhoK7W4pDKInV8AnqxsYs0Ofke34gt5bFFPwVs7U3t62r5pFumqvnETMhPazBKPor2iv9QZ
+NaX4Jx0HVXYsxIul7U30EfTb7iMjlhvW02sedXPf8HQ/SwkIfTt67dS4Dh7Bj9ix/jGkZwZ4EAD
vJ0zlVP+HyzbjxVvCBWKm8Esyv6WWK91oFvSfY6tT0CG+/KI0RGxgrx6rO3alnzPryeIBMxU3DAL
fiYvtzUHH3x7ZNQrmYrBLFUo7Xl5gAJMxp7qCQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
tYrilGShghrwg9h1zk7UFOrnqEEz+jwhURB1wxs9R22Kw/OAjcwK6tqw8jNcBYwhrYgECvFKl/x5
LrnvUtJIhswlxaFlg1X1hPXxL3pzjBrpcsq3j4fwK6AhTWPiYMP5HOASCpo2aK4x2DBFEV2mlclk
MOXfSq5mKZUBIfaMsPULNbYy+Zv1pB4xvTdUlhZCuYcGiLGvfgmNcoye4H78Zuz8SKiv4M+u22Fv
ch7V5O8BeXXz5MsPX7ppklzUzCPPT7srWjUeShTpSlleNInlNUbCBcCF7ng/jNyBV26jC2uIzlVH
kGJN/3kwd3/EXHR+eJJLZhtppong6L90MN5JQH+TpS5/EuukIOUeW6XLhUa/dAMCuIy6dXodzvSM
AThJn9Ezng2irbsjuyJ4pcR8zJb73caHXtfuYpTemiTsTwz1zF0v5ziWufL817hb7+zWqoJdbu1M
7npcibFE23AMNYUOhQreByfmTlQyZJkNfTyykiTltyTPBwoM2w/nQ9+/7pobuhpvaD7Auj09ZpT2
zu/MucA5rpkOO80gT0dZmSZl2w1HmVTKESV1rN0gmdORHLNmlQTIeoJvOebEQ20oMSAUipCAj3Tj
7467k+C4sG/TbariepoazD7W012FZrzRBSIsVW2VbxSdsijKLXSy4l88o/bs1UWx/imrD6eGg9kd
AakhhrcVqf2m/3pSXuLKnz6O5kIYXeb9BSjm1miHbQfF9I4g9C2cjcwDNkFF0K+duetAELEyjm6F
3KbcuqgoJHKO5PQwXWOumWQg/Oq2YaWZoS3hFwqvBhDWIfskKwViJB0xx6rRnUr0uHCFGwy9pZbS
6sUApF1R/CEyoMldq4KAvgFWX7JRYfxIEqUbiogvjA3i8/pNNAoztqsNtzpJxaWyvk1OAh/C0LUS
rh9UPhQO5pvV9o81mpgCv2zQg58a/jwRFnQwjPYPe+ve9BD6irv87Unrf+A1keijA+Ra73e5t4P0
5vcizYc4ErOC/MRQYlFXZkFm/WJPSZtehhZyhTpSC42cSk5yYa6EUWs4tBhi3+BOR9ddfev7wYqa
eyIskN3F8J++slJd6//aWRtn8j/e5P1l4YjX5XbDz/re5VmQU0Or0BmSnXw2WZEU4tA/ngd8c2Kj
jW6Xdktqfr47DMaDS0prkgp68LIvzGggdevDLhi8Q4CAX08NhuYtArOI5EjYwowZANbW2yreqHJA
Q+T846iIdlQtbuVUlSNAO7gV7GL/gof9naaqXP4zyxCMwkocmvQIgQtRPOPA3YabMDBYfJVvQE0L
rLzeEhbiRBMiCXNIA/WSYkDVxys36f1NDKgNvJvaoGoDZCjPi0r/IYOnQjCwLdVtwGfv3l3C1+6W
N7ZjCm+v49N9f7DBi/+uCINRokdgpC/3LkIAqYVjISMjSu+oeHtOM3nXk0NZ6aov23lwcP9flWfm
PHcHJ9hwgCm16MNIjlaW5aH6LFL/+awXEXZAyZjhrLHclIikAT2d0JUPha+SIQf2oFYeqBI2eskS
srImAOPusls+eBGruhKJdRL11yXdjTk49CIqddD60/TlzPwG1+Us/lRxs6BIXb+zd3IvXNgOMZvU
qWeu3wnbgLE5+XpIfswySTNQZeuY6vdnIWndTmp5fbHEg2t8OoAlnkd7PPXtYlhyLSQ8xYWEGDFT
10Fov7wbLSlo3EEyfZJa4UyVJOKR4L8WpMplrHJ2QGKEHBzZHziGuNX8736pYp9s9veyRjEJlwlv
IoPFg4OfmzXxJ4T4ch7DDf/VD4BANJHAFdNNG8QKFNctUvUwItDeBo7nbIu7jDqG9EXdOktvkWYt
CPTdCCOVNn0w6US8t/fRQLDqibIavMG4qDk8ipyycs0CLdO0RYDo1WNluAT3dW4R+u/uOF7iEv0Z
O24IcK+hYjJKYMMH5Tq21/FYr3KwIcvs01iJDl1AptBUioSy9O9bmDtYKsK0MmsT0b7nUcroPbju
veIko7k25gGbQNwHm9W5qLEmzCx6nxET6W/jwGFay/MVplBI6MnTDuONmfyamv/694SRr2XyTI6x
qk79DdSFUtWpNIaD8odRu100xikCViqUZxNncVWl44oD09IGD5MN1VJbHgH1s3xPen13addpRHqu
jvxQ/Yys5YMgEyOboMBjWf9MPm0CUGmQ4FKBNfbiHSGPvThugJZQrlD2NXz0AnkWZ8XcrkIUcSLh
DQ9d0BLj7bpEggj9zw7wlgdnLe3ytztpxCJ3z/8O0U4SJmX/eFZ+Kslt+/wfC5OQK0vr5ujmL01N
MNtAOB9r6otc2Fy3E1I9p/U/qeS8nf8xaz3nWtKKR9Nq8SUhI9GSTjEU2TrmYURYbh5FDOWbVbZM
KypFYY7GwpJzHCNP/aNP1lA78V3XB9mlJ6FOumHhX2mI38tkFORjGZjPcqRz9XQpEb/QfeS8udIu
TC/GEqTfXwduIloRmc6gG5idxLodREK7H1uvAWJgxdbqAJQbkRuIDsIwEYwPqZLEo6c0tjgCNtPb
TXOGfjHToPdboCTPNrIV8n0BwTqiWoIdY+0CFO2tUSu59ZRQEUKjcAWi2lJWQt37wlQAQv+Svy7v
ML/bcb/KP11xkD8H4eIBx2LG9nkB9uvVXJ6jwG564ylmPXBD5LTfcfh32YS7nnVN8L9+uf5sow1P
owXZtbzCSJPbKDPT0rDUcn82LPHp7xecRd/kyWNkC9+EOiZpunGpy55O6KraRTSI0/vdpmiLFkSn
Mcao5ZKP58GUYyGq3GXvmF9yZMh6wT92Mx6KvnbBeQbYth8fMvzLArlhune0+5A/LPJyD6dVlvL/
T/C3/piIDQw6Fnmoe7inqGvH3mXYOu1kHAyyhoYbFQXvRmfWkUwLQ+BCfhfAp+N7x3h2P3Y2TIPc
11pwTN9iBkcQZXcm//gcz9jTyzo1L887uAEHKNhu247vMZZn8SRV3nmguscawqiKNaXtr4JomY+k
N6GUZrWkORhMnqayayReJkFd46o6/az/AU9ICHZL6TbQJSh7S0jlDJDYGkci3ZTdpHDGnaqfbrOM
i1oVApvjnyUMd97cPqubnyOTE3uhuMTU3pzqbqDAmysPm2/cADHWAT8RlHJwJi+nc/nJusrTKgTw
CpStkimDPjPoDn4nc9kLBnTCaAQcvmPa3ddB/l+coXNiUBqsuhgILLUh1R/z0zhrb411zPCbLZC4
1dNrPK/ffu48wn/F53ol6IKI/PSJHf6rVsad61Ou2IkYMGp1SGwsgmyyJfXMEacmLl/odMCs4hbm
/NtElcvJX+8hfHklNcfPL7rZPvWErSM8+F2ReTD8mNwV7y4cnxfORrxm7Q1mn+XpPQWbCA8nakw7
SjGA04kWMzI+JIGoYd5uhVUve1+uGUL9LdQYyrsv9ViXiYUJXEc/MA6DCHcWjQK4/eycGCog0kvJ
6UZP127yM/MQNbEqTOfQdiyEl/5EB6kI1coYpGRcM4MwcjAr58qgl5EvOsBcZCjiElxSmEgzSAkv
bVcQsoorguKsQ8We/K7wA8DObYXtg7hcOPQnKSCcEp6hOxZxP2u5xY9BTKYcV0nSohlOJXwvQvym
mT60t9JlbA+W/yPABl7FclewqsRmui/2vIqtMB9n5sbzJt/ze64wtz90OzHCGho3NENvRRr27wTO
FbFGGald24/hWHb7Oeep6XwfzTCuVzARazZyHnZtXwkRGIdHBEyZZebHuPbIE7piprebngK1yPN9
GvSKR0sC9vHY/I9KT4cv42PGEfP0AGi9lYU+JygdTj3sgmoEdH3WpMKtpbgs027gcji52mkcxQ2k
DVbh7XL5i5AajnxyZsozBVS+9AQRfa2uQjfhz7lZb7AYNebAq4atorpYSPxE8N8Witw54TjPTSYT
q5C/WVXF4G5pnqebC00sdg97B4cb6Vu1outeQ9iazAuLH90OAt+VzE/W8sZcko+NA9gupThsqbqD
x6kVxSasiLh0P81guzQwoGbMuyt464ryAc0Qgfi9TQLHDaiuiop/1XLQSlk8U8ScsdaHccvm+rnW
cs7yzGoFrN/+qc8ojmuyDrAD24KSWlPjX3kGG6NSMA5+k8LqIsC/TfgCfupMG77fyXKmh0AAh9HP
FrxbmOT/9Dygfd8TOtd2SRVehapovRgMdaNHpk9v8LPgHaPBzKi3dkhM9C6817I9lpimj29nYlSy
pJ0VXz/Gg75caDpbskYEpEHTVU2ieYD1kZoY6vX6znoMaeJA2eyivi7kC9rLCe8MW5RJ/mrpjGl1
9+jTln1oG76rhDxxaT/OdQ2mjiFjgoaejuawX7DkqH7Ucw15fRVyR9XfXbpMHrJYJiz+el+wF6H2
RCe/PsG/ZRcS14lTKr58e+OoP6bal9Oo7DuTOY7cZlVnRe1PXRWgwgQy2F59Zdb+0rWZlEVMZpoT
N6FWPEQN/GchMN+6GHvI9B+Iy2nxgxvmMGeue3Ly3Aq6QHmAT/7Fj5atGPgbx/DAUFqo9wUQiNcb
CznlUHd8iX00+w9Bh4VPBj+ZLIQqdlqKlkuLmPYBc8iMX5ojB8B+gAENd+CCdAphsgdD6Fk8q/eR
lXT/LjCKrCnp45u9zLIuSDuq/NfPKY7FlqdNVJx9qLbV/chJJggxQFlv8CBu9QqoYzv9k3LxGrGQ
mHNAngMkXMkFh5Ht57TJUp6NGWR7eIwrTeBKpXg4HEwvcrtc2bFAzoL6tA3E52BX0X3fdZglG9i4
S3f28T0LJmDsOnru1Z0avXAQxV0EXqJDtYwT7D0jrBz+eNTcyyiOEVh6zOiO3x/L5fLNQDG0B/9N
UxVa5HH8z15iTh421dPkqqeTHYaS6579vCfB7xtqVcSkBGO98J9WwON+oY2QRz1crrUj5baHStqy
15ok/OewfdhnmLsBb5tdfYgq/wL5XLm5fvHolVtZJn384pxUiw1q0oD9jEkPSB80JCICEBkaht1g
X20UPVg0htSiVhqm++8FWqE4sk49cYq1hu6/4nnxMHL5lv1sljVjUQNbjrd1hrr50UPJLCB7zt2I
BXSlKLPqA5B/phZ2dDN0sMkQysRH0xA97W8lqhmMbz63pmOjjbRoLjkKWn2wb5aL2D+fPENkcdYn
czmEgJKAHAP3DujtZ8pcKN3MNilQH1zQAjdOn3LDsopV6DmfvndEm5dQ40JGsRVliHdf2T1n/+gk
Q4v2Up++g7BZVnwExXdwkqUseR89ZyoLxQAreItjdljj5ETmPjyFBwW4JMsrH6G89m+b0XO2q/zA
SBPNEicYYuCd+jB9x6zGgJqLoIlGB85a1uGKDTW/vQYZk6ZvPDChKmewW03g7Q89bCC9hpsKvWC/
J5SoxsPYeb9jlSoWPRBNobuKMDML83Wn5dmhk1cOpFnuAKAmVzDqAxEd2rVFd7JDlgNtzaXKgfn6
H3GvVdj3J2pdbSz7CdznJPN/lDzEV0Oa1DFxM1m3qcEUAYl4jXEyEkrOcyTFva+0dvxZkaCAFNRR
Y66vQouTEts/z9aQNPmCbUXdcJNVmXQAKOJ2s9wPZI9s0mNtsiqe1sUnwpVAr4MDdSawlj4YWXGC
1NRIAnVhInVoCiTQFU2djFDg0Ortk9QmKyumy4pnt7xLk2auRP3ueTuyetw11UTHDiv0xsTiB7rC
KrndgKbyf6ElaVCR81NL+sSckfyiTzVVhQlvy0XXhoQlacqL2H7gZIcg4K8rxU18okAi7or0dKY2
V7/Z6z++AlGZeHi7Kqhq+Q1YxfV0E5oVfh1q7a0IoyITJVSwY4K7txbVeAE1wOjszgOHfGE1AvMp
KMcYxey5xHyBzPKq3lmHoiGjl+hNxhgTLTkSsqx6T2USpVDYb+pDE74D/TqOTfHwQYsaTHZCMnTX
vSjjDwYB0K5dGUhxrRsQ+1igEpSnfehK2BiQOaVUtv0HYYq43FbhFhtpsJi5rXFldn+mY3w3834/
iQOY00iRsMfklNviH2zyEsUhJ00y2kNhegkFR+Sf3lCISYY+9uE2VLSqdR2WmwQY+xIofJ8KfRHi
iEBDhVmWV3DMOAYJZe+jFaM2geM8pn/GGXbB47uTyJ7KjgGsoo8o85XgCNP4MN5ijkFUcPQmu1/s
eZe0J4l9mVg7LQ4sxG57toMBzMG/CmgPDHdqLyznultsOmt7eCJB8UC7B90HhLnEU2cQldMhC3wv
Br1iqvKovIDK9XhyYieyrkgh2BUe+4IdKJ0qv1KllTOvAsA97+r1i6EqTjdZdzNTtDTrp1zDnriN
Ab9esn/LJ3k7feJj+2wuO9qfdHy82TQaGB85AnTAsbiRpWRsbnDGndau4m6KyBLuT1Pd4wQbTQMd
y8uyaGEz9XLNc0UQ9H4m4Xdl/8zIs9MoVu6qazLwDBMP7+BOC+gY1fLwwgFIzaJu/zhemNXhukQm
XEb5v67YB4h00pvuwVSHPGJxWn6LED8J2MFP7eTfBElPUffbLkYvrEqQhZZJj85lDV8CvTxgooKO
RpAQeGiD+CRAViJg3yQmW8qfpGSY7/Mwh9sYRatJ3Qd7eHjV64pIB4ZXKersDR2OWIlWoKoMOI0x
VPjvEIK67Yi9CGOtdwyUc+dh/jX3s49AFLjaJRXhV6e90O35nawlN29jE4Pp1qmWuhKi7a/j2On8
qaPMfi4cRzJiHox0xkULL67lGfjZWEjAkgjcSrV2wSRUYGvR3XP5P9rczO2VZ8+mCjOsILaa6S87
3hbt7q+c421qJ6GJdMOFxRUR3ig505CvlYrOudVqcmOpXyieFFR3Z8FkAqZUXubklBO9MjC8+2MD
LhmwS1Nuif4AaPpjWDBHwP7zO1hTMPkBOEIg6QD1DiSU+Err7Iz3CPn055N4xCDXycgtfra6j6um
KPGG8Ugrr2wFjcp/5hSmIm1fxmtQzJpeqjFydqFLOwyxL3cUVbohZuxDlJHLmQXqvLc+5229gabM
i5A1CbM+Y4lowNCqEzriM4ufAGL0MAfSKwstmR/37gT5k2WNBLnuqxKovwYCYlzplXf9aPvlRi+H
8s+CF9zcUh5Gv91Nk0a8GvMtbsn4IgiqgOjsKppFVPgkstiujd+J/ZozHTGVKwPBLKQijw9BmJ0O
gXfrA87zW4RHbx7YzkYe5oTFZVE9rLLteGTAnZRsL3BjXC8qoOwKtP6aiZ17VE7ARSdrgPVKrIcF
EtMn0BglxoJIiRYiuXSASkUkNe9WHxkLJOvX0uak0QWHa5aOFha4Opn5IHtm+e2M/b27AESUMgjb
A8+tUvO3Ok8GWbONfQdnV6F7DCIgBVEb+n0aO8r9z0CqNxSp92k2KjJ6Oqx5FtKJT9NjgkInEdqZ
8u5QJO1dtC5lo8il3hitgC1OA8Ax2rcsGQ5zS2EroZGn7ZXZ1zl0/U7xgzFR4aXbOyze/sYLd0Fi
+tEv338AoEQWUK8xTTG/ZgR1wd8cGoqGwHYp6Flzht+BNeFKdSf61c7gksXeLADcAgbcgK26i//V
uCSCNQidafiW7pCCILDYa6gareTU3XN31ekUXLv5IJZvuobTukWkEIMmcEp1A4UFJFdmrew72DAT
sfe4LUfzvDohKEPH9u17pLLCYSaPzkHs48Lezc8L/1FDUMbv/LA6i/IUqNRlXi5eIGFl9XVUlpAJ
FyG/8nIBiu65oF8F2sOzVC2Yi0QgFXk3xoLFN9NVuTkLoY0DNJ+s3ai79rgLTRGYhWIRR6NMyFVv
1UO764ikoc6+wO2wLka52OLo3Kaj1YFphI13UWbVszt3HjWKLp+3xb8L43oyCkDxqWiViyqMTWOq
BZuOwj0/cz2y+2y/LDy1YDdyTENJQsz8oMoaZamAoqpTTdCQ2nTRUjasSlsKqxPyZKpVvFJvHVVm
ibONoWePHL5QlNyvSuWaWdTGymBp03u1UNnG8P07od6cwlNOt7vmS1CPeiDx6lMbavlnd+Y+n6FI
nGzE09HTnGj9SjOaro6wKYQ3E8wYRi8nBUzKBfMdQ9KJmpr6WcmB4lN/kMvnBBD5wyLFPE6tXBx5
iOTGiwUamDnIdL8UZx5Fv1pmQnZC3T/t5CqFl5xoMxKIdRJ5O/r799/aZLG1FZbY5hxRi8WONTBA
Q4YsbPNIlyWfXJsZbUXac9fQ8QUIr8++HWN++ffxlivXrNAk4C5egnQqlNSTiA6boMa9u3Cg/msO
9ZYanOUsAp1v4I91jfhWV5/9E9Z33U3cpYlYWAe6txRvrLjSDGQ5X4iwyBJjvskGO/p7e7HT3EEZ
Q1y5DlCyYqe5bYuFSP+6T9zJotLrs4Gf98qTasB8+Olptjt03G1IzqeoMkBa/hf4VOfGfEzAqkpa
ownP0eVfnHS/mPdXlL66o12oeaJ8/SbHHSLxODaEtZHXXRkZVuYylKtAAidp/lVfn8nvARs6Z9uN
Ug9cwIssM5ytQuQc6W9+v7vDoZYsMORftT4cByPuiqtqvcuGk+ZQ0jVJkX9BY9dajf9pTGQ56rTT
dLDk+rLADmpB+nUoUakzfaWKtOnjEkyzaM65OgvLlufkF9Xx/shKzAY1RSprZzpOJg1GXcXF0YjU
oLPb6q5tRZdOHh8OMG9+GIoSIAyd7MdPdSbqlPFvigjZ+/PRDuZCC/VnLhFHc3gcP7pZN1I+1ui1
FUT72bRc+VzuUgZqd9Mu5PtgRgepAd9wpQioM/NN0lRgpagB7zYnqV0EjLpAfTaCO+BdtD6e1dqa
5YNCGRXZ69UkPX1sqH2zeLAOgwFgFYmAx5NdAPJzeoj/8QKXsZRslL7vPJSfW9BJJuuEtn20b+OU
YXQrt6Vn6UP64s95OllBIsyIM4AJMMWmEKtYR9PK4yMCw18uS0Y6p8B9SZjetUoOj7bNZlv0P9Ss
mUzIZNGtmdh5rogUEh5JsIWMZsU8XDKuJQTeBM6njl631zZDGtCioYwItF2+1rGrTPOwZ1KvYUZG
tMvvQuAVPzKe1+fQpOfQ32YdX3gqh+163cruu6K2UvNwZwUVojrtzxfOxwFN8s9xOGziMfpPYCw9
8bvEt+iwooUNFI6nFQ/KMGkatzF/xaIvDMlOMPrtJfY2WGoIv9jbBERwxjOXsWXEbQrKXqTh22zH
jW76wJxEmrCrkLFeRsUujMAYhTWsX2hjB4n9hoRSYOqrXEYcYJQoG30jaFehhUJ2CxvR/RX2OMK8
LaZtg4IGTMq/yK4lHuuDY4VQQO8pk0xHpHRa3zUNqURoyONnQRzSZw4gTMixfP/xu2TYsbfi7V99
lEDx40i/p/QVzNYvahlJ7Ohly21iql9pZgy5klLHq50Zf05YY0lrj+soP/FYZuySF3ern1ZBC/jO
+zeO4u8KypgBQ86GXkbSE+RwLH8AYiB4oe8RHV7Akvz5Nf1wRUz7HXvLcAMZMu3Duvrw1z2eVsCv
795+BSV4SM9wrZRueFUG5i8OfuHxxFHGI0hfY5JYS4H8QvGTBpTbM700eM34pKcKq6XXwuqtne/P
dJWS5JnX0mwiT047G+mxDQaTE4nWwVSMj+afiv6jAnfVh/cU6PBN0RKmW3MVvRjnB1kwHu7y+HJ6
g14DoBmajSY0+0PHFRQmCl5ijcJ4gXHVJZRcUOTkFq+oap56HhYLmOVY/a1JmIMiuEzoRKPhBIDj
cbNu1yZM+QDDwJExWO6AzYTIafDi69LDSJ2W1q3wsCvLW1o7EI6nN738YWCOdg6a7Zzju8DTIhW7
r6ELbPwA7tYYsfTu6irTIsTWMCdgo3LlT5xvZunzyEtI5afz7Hd3grmBvvYyHGyQ7gmTEXiaq5lx
R84JRxZkQtE89C3HYpAoBrYe64T0kY6tiQAYiqhKzgXXTqx2y6yzMQQZfIx3X9aoaEmKpsKikjTo
nbGs3xCRVelcdzjzjNqeWzfRcfVaXIGrh15ePlZYC+Ht5JJGwpAh/DB2UC2GGpAOCFPxOrz2jYV3
ZEVPa5ZL+1bfKgZnzsDU2LrdAvyA3kyLRPnGz5kvB+8rspOQLoT/YLo6gb/dqHRI3iAjL/6p9RQH
7URYoEVgQc6HEd90ReFazV3r5MOwtYbtcyCWZpyTsJWm79KHjDZFDeFuSgfdwazq+3hQRr+Jajpq
jiPyKEowcf6Z48JBTNOfBIkyz2SjG2kxebKXXK8p3YGWteZicKVB5rYWpUB/eUywRsS3a+UJ5Dcu
ngqbKLXBzSVqnWE57z3syzRfro1MpqR4h0KZBYEXAYSKasYYjnn4+glqFSj3kirxnDvQgJf1EgmY
DR1RqNQbgdXyR3WRm6py6SpyPbIbP6SPg9+45lww+zvACKseA9SquJaSeSTQ0zoDfip16qPMW6SR
I+liAQsAi7zZef74dnt+EwxzLG6ARQ8qIM6/SIa9sJWR2FParpOoM0fvEAb6r8kZeWofM3YqEnxR
K8ThkgTxT2S/04PGTu/eRzlL/f6CSsKWmRSraC0rFStBFVMGGkY+Fn2yKLbh1x6Kr32QY2JbKzJJ
K2oHAI8DbZW4jDKpd0ulWBNqNlpQEbwPc+hRgPhu3h0NBLL6eQv6lSne0pv9sHZzNT/zesM0VjHI
olyHMsNXpqRPERsoBS6p/8xqeOZ5cJ15cINPNLzDe+Xpt+p1sm6Q5fVx9yPvIMBM8XSfFeSJIq67
ptZ7cGAX9AFUYsYTnaXTao72FNwDmhbIjeYloyRg758fZG3/4KIIWnE3ShzbAHl2OCDAxKzAhsRa
GR4kQ0PPGCapK+AF1qiWCzy6YoNM/G3n90DB6ui/kC28ccRJIrrG8EsHq1vKLSRMiYd2SOy2jIQ4
1dyv/ReNDrjDTY3KQZmfgta/D03StnT3+cR3p0soY2Guz+Y2OS1tgC1rxGwsjabYuzfClLiEvbNx
7EZwD9lihxkK1U4M54fOH+t4iqWf0FFl8fxRFvEfqGd4LaO7OqDNDqrrjfbLChRHpTuvgTH17aLN
v/w2XS8FEciEbd//B2D7P3xLItq5xO9OZm+J0fdBHvUfagQFj0Szsh3wCw+xczMfes+hDxh1PDI9
51gyUHBzB1afPsfnqq2HwYZk0AEgYeuTpqG90yos+bwn7XpwULlF6toHsjmB7iRMtdgBuwq0QXgJ
fgPTcZVKNgfQ+O3befLtuznx+X3EfdYnc/LXGFdIuXzCU6uprrVqwnY6vYC+FDLoXQJtefaySruA
O20EXS9PbzFjnFAXaBi48m+U3EgnoRZONwmGHpSudSyLyBz1PtLg7hUKi9UgWqx+UU6DIyYrYtTI
0wDpkGH9/gu00scOQhu1eYWMLJkMdp25vYpnackJowl+oZG/vi2rWUGkoFtpE2T0n00l4m8jwcm5
h9LqU4wx8RP8dEwqXkWaFbRAdcImJi3bPvZ2oLXK4fP0EKEUzS1HqOzyCvNRSxbmNgphwYACjlWv
0K8zaDZjK7ru0hVIGiNRokDDwTISM9zQ1Yi2oi35XiPxq2/iYp3SCLz+MXw756VGMeJC2zVMXNxy
3J+7IxK6Dp/+whVmeDEB7L5KF+k+RX5ITesKJmxCWQL0JXLF4ryW6jGtWSsDtkjf64y2qkkhHCTq
fH1kNMVD9HNOv/l79xzaZ2XqtIniR4tLn6y1QU5unC2+YUU6+xUindVgKgK08mryzXErxwqQscqz
V4ACt3QTlmxyCoWJkilufkFWJtYBrkQ/SmigYws1LGlTD+Yl4moDmgBliUk4Q8offAYUN1y0nWaQ
1w5y/OBX0c2y+qcGhP/J4a5z7dd+baDNEYDJV2h9htQFnhL63I54m8/X5oOJQM7GmppU37QQKKSX
NFimlMlFPclncOjISPI8zE8BW4lC6rjta01pkyx7ZrGhD67fc/KxbbWxpxPUePKNkLz1D7ZK5okl
rQj5jIg2R7+uJaHLFboWh1BtxMruch4vGNUhXfsGSuxKpMv34w+NTLMcWppSevt5Xb+QF5gFtuoy
hdgX8207VI++s8GgB/9olPNxfhyf8EXaRaoiU5JxXJS17vJSvICBRrT5/RYeUkfemC8Gm/iCfglb
huDjMBXLVN8yOYJt2f/2bPZ00e/7654xd9/AuFa+dV3BGTsmdO/pEY43CN/ISoF7IwA5uFeqjjQJ
yEwsQ6LIdRAs+7lYeMN83jhjZbUnjrswnEF1ATwMZj8hlgvfO5vdLfgIeo2yhnt1xhuKY4hmteNL
KCFc6EGmfo05b/Idzx50umS8Ui+dhLvVTJwuT+bUsSlhlt4i/00MTk9YTUeZCYqzlH0g/PYGegmw
Jq5WPunOqirTK5RO1uV9ckxHZPujuwSY2DptIMHhypNkmQtirorJEw0/RWN7ZC194nIBaPXy9RnF
0NlQVxcV8lVuiViJh3PrBcdXl6eMuzR+rXSUPUBH5MWOo6qwbYkHkjTPYqgYn7wAXX5ss+vc4oYf
/apjqWbVPX0uUeeEC9KXdB3ChcPb6zU/kbrIQ2SaQj5yrhczSfEcE4myLncxyp1uZC5pW+9Jafg+
2GUH22C0vfF8ToYQUM4qmEmSXZE0h8tWTSFGgXW6mhOjSVdSZppAeBkY3qwiWBRVbn9MX3PWQ+Dn
q5FVAJWDgC3ZNHaJG7CcCsaT+TWcZejOq9gbg8F4Pusl/WyartsEJRpbqFuVrPpr6aH9DVLoS6C9
3vfSH1A14zUF8yJDQUTp4QuNlXtH2nkxCGQ7HmqUi422F9uOKHWo1I5VD/zsFyaAGJXOReEpMmeq
tIdlOGGYvB0OK81pIqGUD4RBiRVpUMXZgCIWTm0g0WWFSStyMM+uSBEZoUdxp2UhZ6nGuL3LrvZR
LCA+xbrwuOSnJFQRIn/VWKLvhvLOw5TV3hvX6SaTTtVXH2t7NogWBb7Zq37hJO8XdECxv8+8tSz8
bz45V9ZOG8Wmr/322T2++m0Qckjltz7kuY2rVU2mbXv2cPIPgh/3s/yLM6gcNXyil8YF2HL34aeI
TQ2+OdrV4YUwU3kU7/S6F7HaqCSKeidvGkDiWxh93NJi6itzRizGqBqiV2ih6J3edY+2pnRV3DeE
KpPmR6wX5hoWJjjcy0x7dqy3fwNWkexomhfwlOT5ZTvJcTGL+JKqZPyamT6Xeypb2UViOGy+hExv
LNjYANxn8EiLEaEp7lu6Hrgg/N21gve7LGk8hHqqIli39fJw+spg/LHH5Dmjdn0vLOsV7FtmC5SN
4kyQhKMhRDq6jdUkdQjD/R5F6IXAj/CZWvXr/Wzod4ufCjbeuTJCrxPv+Ov0M8TDF2gz3vj47NIN
f74Vr5J6EOIcAdaqPLvpaHnW9B62cXBe3hvN+oPS/IKpGqyZfZP/8t8esKZWdVsqE4Xf8d0iB/tf
+CsZVVJwgpzBfsSCNB2Y0XBVshjMnKTuyxFUCuNVqPtnM5JJUvpwd/rOe1WUoBYQNek63ZAfcNti
PWAkr+LsQehtcJm5hjEUsBhyUGD2l3GKekHYocPqm/5HyXbmwIidJqjgtbyaJUzdnpeIVny9QymW
fbpMPw9CBsSX7oxhDuaEcLhDAmIwUs5U3pD2RTd7k/WABIIpIaQgICdb+E52nKnn/Z7QhNxOjWSG
8rRgvhGW6alhuk/r5P7b2F/h3cU/iIgHo4HhYLo1MCdGPuTN8xMYIUOgYyNOG3ep4lOz5tZvvXxo
O4lOEGd1Uqucw6Htuo4CNGgJ/N6agsIglW5V7qWzactocHtorsDRcwoTYaSiwXwEPT0sjPzdyA4C
dHdYTLI=
`pragma protect end_protected
