// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
t248lPuLZ5e/h/v/wYhNdM33OiXeC1LHvEnQ4Xqr1vjfhiERN6z2Ssh7l3qednrz
48nj0GwBJGmY1I6nHhFOsaSwjktYmQyipPcFC7XCB7DV/nYaSvsYXSQdHFQHyv45
c3snyxXrbyG/gRozE+OcWZnaKqOTIWLtUwoOf+2NEcw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7280)
sIa1EKeykEt0wUmWEANogaA4y38h3fiIgv2VqT996B+G2h4DtxvLvstPkRAx/cPH
7SKBPB1S5hIHlPNCauVCV0KN8DnLttIU7qECREUOjuJDwnsTIAkleuIuRIHrrCky
VoUuRLHEH6/23Zazw8b3O6msDyYuBXlbM5O6d/GjxDKDpyRhR8lo9zJK+Eq/6pgv
2XXaSXP8ct1Uplane3uEkFIRGnC7UUdGX1imXIfWLx+WFUlzhedXzLNotrvjuXVz
T748FxF/yMTajU3qioOAOLvm1F7h2CXJn4mLIf8bTUpju3N5pmGTD4mqlM6Ye6CY
S1mrx4a/+mItTLwbWW3PkrLEZOQoWiBHZpfB+ZuUj2o64U98iFKw/QpISCDkffZB
Cg9t9A+abFdNSXrGTHQ/tfhdriubC8pkqMqX2UnpglfdbFfFQNxugqk/Rat2zI/2
YwNNB4iF7A5wFogoBK2t0H35I8cJdYVURF/lE9N+64YBeS30/6IxT97u2UPZxdc1
IzTf67RjFQRt6Zg9AxW4pg8QvEkHUvQBtLfeHC67Jtc/TQPGQSCpkMwDR9RJ/4HR
vtebzJMFf0w/PGBJoaBkUU54njH2P5Tgzg2FLA8W7cy1DXkBXNMj1BErDr18c+pW
pLxneZhouTm1Lq743xqM6LAmktpD8iaJzvLU7EvDoKVZdLS3tmHdxYa0xETBdIDz
ur3l7BD8Hagcxyi/lQ9vhpqzOP4yH+Vo0WVLFLZONp8xzFet0EhpTycETbHk9xz3
U1V6VLsqBwxu8zBDSKBBoYrHTzY1kjcywcYuXOeEYF8kW5Nxj08Ja4WAB8p4kJdM
UNTyCjCTq9Rhnl/+v1K0ELlfeC0eTEtXzB11Xe1O5BjWnIvxu6/R/AcABXCFHX5h
IMnvVdnhw7Ul29fJEX252cnWNON2COikUuYLyczP21dxNCdY4Ih/rlTy/6yzWzEk
xirMccX1yP2FLtueQCuYemmmQ8qTXdO40oBpXUQZ+h0tO4AAKIvJD/VWSaEl0Byp
5+dRtsBgSywdOxUbJe1VMutQpdIWC+0t2RypD75qOu0ZClmgh5uxogn3id1BgTwo
l/hy8IjZy+e1cdANKOBID8QTdTnb6mO7Ih7qIQz+quwrvSh3I1U/7gPMZ0qA7qZM
nd+OIpTP8uAFbi6tioZw9gTSbbF74PhwYjDk253s+tbv5vsll0jKtZ9XlSmMYZrs
AvmxVw7CyyDKeUPPbR3aBWEihALSnzCw2YXotcQnCMVqzUGgTLu67SToMFyHEjaU
M5z0khAPznnZsTCgeiibz6OZN/ozGCH3EhoU4zfYAvgDwVuuszeO6kZ0vFYlUlRX
U6kcya4lym0dw0P2VmVHi9YOmnOhccnI1px3yB16MNdXa4wXRLb+rLEETJ5sfANv
4PudblapJTGywID0zRCR/Xcbaa1VOg2A2YC7ub4WbI/bMQC75+eKlpwvOpREIUuM
en+q4KSN7Hwuk7EajxngGZWlId01q3k0yee/P/66bqbDSd15+8z+3cmV1l/yfdKo
6XIix99exWX7R2xtumfzu2UKMXuPE9JRA9Fn07vyZ9Mu46iofsLGn79RnVjWdmLS
r+jPkmcFJeQSupnnEH1pX4/jATYA6G0fnLXevEfAqi1HIu3OPEy3By+jXVZvPgOt
fluBkzZwua9kMkFuRvg3PWh4+xX5pxACHhKWI+lu8XAqPDecx7VRoC++OLt6EaFN
wtpqj+FxWgJv37WosRfixBsZ6rgXFxjQh6OGO7a4nl6KbYaILbnT4qouKJgcjBCZ
kPyNVQqAMWEGJu91/knhaOm3jRQNSbrNGsJU0owLSPaS8AK5xdTLI8vejDkbVF3Z
hwnGkCmXYTu/OaX2VO/ngu1rhrIrQha+Y2KaNTu5gcsNPQIZhKHzQv1A4PJUAj3K
J8ej2SmgzA3cxzWF+VCpttwOMk+eMjCpDAFokhPnui2CkfKLwOQOAIwq8XzO8Ic4
9+YnycvCJcrJEWfvLItJ4ofv7Tmj458pxqeJx7sYmDagZ90As1ZseWHvZYVDmbJp
Jdq40YJXOxTGq3Ow4iICjZLTJX6WAs+wDYPOEMDTGVSMRdDE3Am7YKUvnmafIXLr
lXTup6EOf6Ggb6HVT41h0zzI+E7+toJuU25B6epBusgKzZ3lm8LH3dCIBOAieZLh
y8xufSF8JZkOJbyg+tWf1wqay5RZaU3XRWFrS6fbzjEULQh/X695htl04M/LKY+I
dEA2Y38ofRbBJ95qd9vgI8pmBZiOxWaqwwt30eKirAQsew6JUXq/nUieFF1mSRvW
SgF2gykOOYJrd53f/3tAXE1towEQfSkm7d5JXxljh+lqwFr2Bz1YeUUONhGTrtJe
GVut/EV5b8UqpipA62Hi9io0ZsW+WXaxiYIXMLVW4uu6vnRSTE1F12LC383Kch1c
WYiFgkWOR14nScFqhz132dM2p+aOCwWOR1BBoa0tgLX/e4/IAM6JT79CxBPiEhnd
8kAbWWHhOH/7AB7+JYtYiq7cF0e6q83Vr/BX265AnIq+5QRqK2A3aFE1kyTATFYO
xpB9AX9Qqy6xS1IoXVp3FJgt+HTNwM0Bqn49a6d1qDdiCX4UJBXhTQXq4GJe/uZb
pJ+k5IslB6jdj3n3rA2agCWgx17KbaUJNCgUdCBefwhKojWDblRFLxlZadfP1STU
KUM307oCU+fUDsoyZ+QzBgkyyd9dDzY3yP+uq05ai6rMD+5b/FZtcGewGC0hHyKn
W7ck/mP/Lk9IwUQnGT0cbojcxFbnJJsXz9SOSkiyMMh8+Af8kH3A5UU3oAFWkjpK
P8bQ2ZUqQdSi8a0jWenLsLSr6BXFmPgnxxq4a/bwo6lfXihqlPBAUUln/7/L+aLR
y9CV/Pq/ScjsNbwqJiwY/VQBIb11SqglDzSUBZQmYREFsuvMfkSKjHO9Vl2X9cUZ
K55Qi8k7gYgUn4J7+mAhWxfiA3x57EmZvFeDzsqfLbYHU1tDCvmjtsghQNPrD/+z
RyIFFIXZav7RRojQCWi5LI+wiT7b1HFpL4u5Ub7Ly5j3W9tQWGh/UQoYu77Mzuu9
AVbiNEHY4W8zgot5Hzlp0p1W7LU2xo0IBC2lZXa7Vz22huQvnWRei1PvTdPF99eh
xXlf3vPRXBvoNCU9qu5uO+lBmmqtSoOPGvZ5EWqqTMN6CB1Nyd704n2lMFXqi/iD
GzIm7DyLCOl148xSZ2OZFILY4oVWV9SlZtUmH6Z9t943RuMitotbjqfb/+zaVMGP
vD3wOQPMtS855nVWi4wJQUMgSv/yVGuXbIupA1P5CooA4vz53TZKEX+jhBMHJPrc
xJl/HYKqXQmUfYAK3n3Ad2r2yySUeIHfONZ7vsUbw6eEuDwd4ABvmQ3SMrW+RSf+
JWNgoW6aIcR6ai2DpfTk9XuD+8TagbquXdWZhbTbXvnB5Jf0PyowvcloX/DUO/dc
DwUJU4p2RhDLr0MKkA4SEcf1JBfiLSFUndTwtmHEu/t6TCIJje9RgWcoUuiwXWLl
xooZJR4v40Ddx1aSB0c27oVozhwRYVYzdHxH+ljY9u6x9kzLE6kh9ZmWwFzXnhM7
XyikFJuxQpTCPx3zUdK0YqZJv6Ibdto7hu3i1JufnR12RPyd9W9OF9IGvKpM0zJV
uf24ZgKay8A3bbm387OHi45Gx6p2GIaJu4KOX9iD8ZyeBAV3eXLv6vIiYipltUNx
k6QLJv20idxpa11BDeW4l5lHep0ZqH3eMstBHEUrCGm26gvMVzoCPk0QzBRy0Sat
U4QFAblV7+kn3JtP1766jtzYn9ux9xLOjiS0mAug7X5h9h2tu58sLP4thIjMTSp9
fW0rA9yxHjNMtwl7R6O3Vc+quV/roJR9LyVTFpTwJ2bO4naeWAMuSTznZklB3GG0
fAodtXRx+sS0u4Gb6YxPIbSEHtSWcFa+P9mVNxK38GsDE0tLcXY/J16MlHkFXP/i
uFMNHKNuE8zmlbf1FxTaAfV5tFiLPHVPFmujnclVIKZVL+gIyTuDurm7Wk814gES
awjEE+ZUT0lM14flb9shHPi3dowWn9QZra2c6azCEksjeutE2xFjiPnQDT88KpMv
iZk1QklgZyWHZVmdLIzJNzigZeKFtJOCE+GxdPwbzXd7VGadWeihz/loNOJNvz1S
dJZFieSJz23eu2yxUYl5YfADsTZIlMdPdz0C+2lo2a9RTgqj/yQ0bIA9MxzNkyLz
Z3mr656A1Naj6wwCPXCfFuqGbiniKntRvxWip/uSRnaDDT/LIuzqhFE9SGdKW8F4
bsT9v425dm6uVBtM5knDxtQZGBFn/SpxVGQob3DPLqRowSkXw2hKJU45ahfCsXXS
2neKeCYGG7U7SzZIMssOyr0Jq0haV1B+KSGEOddUmuxvmfORRSuO2YcO1KcW1c2/
pjZ4AJD8eGz/xGJKusQ3rfo/BblbVyDDXFj4wCk9CZPwh7rht3M6HMvE/sZPQGjR
jWrq3dNMD0qsH6J5WCLC7f0WHcwiwzOSiHWA+9r6JCP4AWmXyvbQEmp0NybSXZcv
SEoyqUL9ewLObUXcKqeeVExOVdiUVYgYqreYaEmISDOj3wU7ft1YCqiJwNCwPefO
rWYEzRRQPagBk4sSj8fvQmKJ6NzBeZk/txY0V23M90gN5eNcZ2WVLMdGMGnnP2a9
PzCROYnSE8ybOpMCSsK4aJ+CQITuMSH59K+LF57kAQ8XIPKrxJIWLoDWlHgwqmVW
2fMbhADfXfTh/Tt7UmjE7SBRxHzocudFAeyoAolZ1yvy+mThFQzNkOItVg27v9kK
mlPmZgOcpjSyEp2cSOh+lBKTE8eIXhosb/v/IjwIb1yCNZ9qVgHZUGRTRCtO66hE
x/AaLj6TKJS1nm/Hc7FNMmoVWD4RYkW3zTxWhz4m9fAmElxY7TKF9B6tMrub2Dzh
YvCtS+bBJ+YxgQ7+EK6OlAYPqcu/mFIaT+4Rl/QRO2cT7zyDyTPft8F7siCtfglI
rQlfb6egpLJLg0+mL2bVFMFef8uj8nL+Od7aT7ZKQMfCbGyDtvkOElqGt1V4msZg
LvitHWtqm/OaIQn/je81FbIIS/2d4GvWopQv17o7kD305D9QkDr5KKZBkwO13/NZ
bKIPP07PY2oLOJueOSSfnLaawuQiTx+mDtVvxWWOKVbkZsMJCPYuwusPqoJX32rQ
Og/sIzc/1+tTAPWALMor9G7kIo152eNzjajAAZl19O1vUgZe7I8OofkeZW9uLqs/
nfRiOg3dl16uxRLVJ4bnraku4Va4oCnzcMaAZKo4l3YW8ge+FsDOz2Z6hthyjUVB
gxW4MSJ1u/1uo9tYedVGYeflVqNIOiaqg6Ey9SMTtyW5cQNsTOcJ2yaHvw2HO4y8
YysdBfd3UmAidqMH86schIzbaQDOq0rml+4V8MFssy1LPdev18brQHlEUeP5Lry8
KVErOhfr6+sWqsERaes8S5Gtectek64Vd1bV6AJeNAEDsId0UF6l4wArLXPFI0Mb
GHeIy5mgYBbkjN4GR8thSsOaN77ySAl4Cs5o+c71Wp7a3/QQ7yuZF7FP2hLZTzkR
KF1U8iCue/3rC5PfiO5T+YE4Sv7AbH/XPu53UYoXeLZDaGgUAtoEflIOO0VHfxjp
cgdthvjps6TpXQmeYHvmmeCt8jtb5sg6sAi4F3kYjcWv+5DncMOApcQ3qV5qRdnU
OKFf6KwuokcYQWARGuBsDFluTDsoPaEzSZrmIj0d4Vr8jlQCcfExCM3a4vIupSLM
4/RB0dK2nphd6rtV0kUokRRta5mQBwiRzfhEYbwbEF66rYRT9KBUfeGB6x3efdm8
Dh65IifTfq0jl3ds0kQFuupDVrWN6AH2o23rMItfVDZmW+eclMaF8D2yRMFAj4Jr
zIvNzb7TgDHdlu/QgaICqvetXrA1CJQKm3kOKO/Ulok0dN99hHyYC3zi+zFoRXC6
hzgPf3RR4SG9Tni8BwfErcRG4eV4fxDRgaHgzJpf7oTLkyks5oheyKVV+9sHL2AC
sIFJyeQ96tEuNz0AqMW4+fdrTuIjsQCcISNGoCAQ+NeOvlKJTuotXC7889UdOThg
LgDkzyqZb/jha4KGXa4aGwwfTXuWFbyb1/UWl3KbHQ3VVzir5wInh3jidQJ/8tvT
+FTeCoQrLaRz4nB5P/9DV+gbK+7MK3aiHWqLUKjkVc1E8WGl6j13EC3dK09Ic7BM
etjmcJw+wQHCN/EbJes6UzUz6shW2yP6fE9ne8XSXGPzsiv/Bs+IP6TmkLTAxFgA
y8WzA+X5wiTNd5+E4NuE/eNIXM3pUfiiHyqKcIQxuxrt3ilHj0eqlLd9+rqgXR3+
NHQfjlpi+XyO/ep2DxUjLuLi1Qg+P8xdPLMdOGefhokrCo4ITzS6JR9c97JGmKEb
FZ5hFfWjIR95p+qOq/wzLJLj9DxsQfpBnlW9mXkZ3Adr8k2A1jdF7NBkPwJYMqP4
cJ1FRSQLDMzXI4MjKmH1sw+cWGVBUsTYkmFBkXngPSRLRmcFV6ACBBXxdT64E7Uk
NmfW1t4amM7Ee/lkOZwvh4cs97D6s4J+TMPN+4rGdXfh+v+nzYL9FduxlO4hrGKj
tdXRdar0JJtxYubOI8JbBfz1tY46sxxfsOeCKyW9hWZid3pSfcpcddvKNXcfUHr2
MAW7TWIFtFQzl62K9Kau6gmAnXYxduEUu8QCl3nSu2WqoiDl3ZAiSyUJoiFvLMig
WiiyJGH6ztSTUHuxA6QYR0QmttFAwjJp/rD5Q3zZp61/BXSGUdwLh4yah82aCOqV
mSanT+nZTUsDHiD+GxBvqSqjrRhdiSWdKW7OkCdYkhC4K/Ksmfqcp+5rd2MAHazc
AFqUffwLD1WokUHPnlk5UoSqntnxTEPRA96+BwmZYapbZbvdEfiWD/ta8jq8/OhJ
wAJOqpZNrXUfBbZCIZfeBz9+E0I6cxqw9GMGWHPSKlCU5k9TdImcaDOEHKQOYp4r
mYSaoZdu204Q6QlriNpz10YX4G40hD/90gyvMxX3AO1yy1IIyH/+yFAZIqVuwkNr
9gsio2oQLIWQ0pvH58r+spQ4knUAqkOBRmKzwPHkdfOKSd+6Sv/voC/IViz/J36+
iMFnqPHcd2iwEKYrjuN2saKb/zCEnL0CzB96fAPUNWnYoRh0XnXoSc0S4sn84BMK
Wm2Lg5LAFb/bRoa8/rRavD4T153RuUT3/DnEsI2sufbmLhiY3U6RgZGnWwevk+O1
rwHVioPsgKpCdpO6gbpLi0hZpZ2v5uJxEdUFfG7ggOAJJ7idAXf0NEsaCji4kb2U
9Gk80G0DptEIBgzeUJwGttRrV3oxZ6MgZK+AoVUKAEzDfcQ/GTak8GhKewIpQplk
w0NKHnDhKWmVdieS8OnmyjxZrJBa/1JMO3NDbw1fm3C8RTNyc68Ap4gfvl+9tlPx
SrpXVzAtcHiqRS64xx//1F6K2kOTGE0lxh6MYXSDN+5181oNSQlaZ0b7gIEfWIeu
DTlOfzP0IygtcZLrKl05RNHoQoPy0CgH6tcvfK9cTX9wV6jJ3vo5WOZuoaLpCijp
J3DNRNd+d+ELfuIZC1Paf3i3rL9/vz7tfnzp78ZL8ZHljsNW+GdsukZv9iJxa4HH
uRIWeKVis6S7fRPQtoHw/E/t6YkQQkmp25rPqM3wuBhk/dVYq8jF9hGBwMTXUN9r
RN+XzrzkW4DU85WODV2ZWAaXoGOTzsyILd3hepbRcE4T/BhUXBLPhWNUToZ3jKNg
zAxx8h7hz2+3jOU7ut5nx/iayzsQAsNsKdW/2UcSal9DIZnhrT5hJ3ixJQ7Ku89H
xKK1u0bwatnrQ+E8QFYezSJ3JX4eX5ECgxFk+tkF1rqtjQGHWm9C1vcOIGJUjAeD
ZVyww72KRjFUS0mlCZ1ZMbGlc2BraKIHnpFecm/EySZtZsIHs2OAryBbMyfCRoaN
P4lBlL2qFs5zEBrDjleo638U3T4Wg6ZErA+rywUSrLu83f6lGwgfkKtKHNDO59wl
jL/OdCuFoqU8X0622T8hGTuDzcUE7yfOItZkrB5f61Pm3cyhgsLNFDjMFkvPCKhd
yAIr5eiIFSuhybUoBKkkZCMxeMvo1HcM7DaOFg+9PnYlq+olEt3OiJQpR95ImNBh
bjM+roJUw21M8c9uuwDCgX6KOZugtkxmGpgkZnBNhP5+wuiFxVUZWpEy3mU/rGyz
1nT98OyNlrpwxIUAy1qpgDXqHDmTn4FryofX5WxySqI0s2B2Uf9jY92M5f+6/nIC
qN9onVwSjL3XbOk6WeeXa9PASdQ/x7xTKr1SNwDNngGTqAkFaX4622wSQ81q/PHK
KtDS6XQ9ZW2zHUSMnAuCLMtCkDjPtDKuvyfoPE8ameEYeX2QtC0J+UOs/8id5Es/
DHuQT3mGwX4ERJ7iR6tIeeO0G+fTX5NHfDBOBgC+hSL7xewidebiAYXRH2jtf21c
BoIHSM5c5eUQteJ8nzOnRi06sAEvIMAUAmixDWmajJqkVD2/sKoO4r/RJJZ8nhgK
EQOkDR5ds9eb6qzqZFWMHGSbhtzep13T/dMzrtWwPYL4C4T7Hf8/d30N/DcPhcmP
adGg82EodmV/3qq73I81GqeOobl4udEZOt9Mavs8B6ua3z/L8lqakoCUmrlV7LWh
Rx2Y5nCfjKsDgAtTm4qkg14Muy1XzEs9Rb9AupGhyNREkD1Tf/Qp+UTfUYWujyvB
GEOg5YZpVvH3SprK5YcfjWBsFS0xxBToirEoci6CxwAw4VAL6RYxaV2C8O/m5zyW
fRxz29ZWd0cp8PbxJJ9z6PuJQ522smXh8eoDCwQbANV4tAWKBk2fYhmtxhC7Li25
ljebzCYBe93Cit7IjQBcxK10zYfKWrNOEFTTEEmsdETgtyyXhbZONeEE6pkE3XNF
sfsjaQQDd+r7Gt2KqjOPwDIEzWJhRCxAs2s2UWkUmLe7KyNaYt//WwDTCsI5FYvC
ti96PqhMKIqKP2MieuuFbRsOMaNlh3I9y+2tRtEbOFreaiQd4/tebFVFFWqGkKr6
XSDAjYmbA8i5fAJo6m4YuBsJUpEqav43FTl13Fb+12i7WuculZ9MF4QEneJXdnFv
H8XxsNTBZZbpr1ciyrmqIKj4Jx2n418GdkWLUSKeppZfUy5AiQ4fFq1VXJrTXnQ/
YnoK08V6BoBFCpEaEoCmCAadl1CLEGSW/A1YQl16uSu1km3XzIFjLQ/oKo1zePOE
2wjFzrVYkEvMLmusM6YhKGha/ld0cBWyWo18L8ey5SYEtLxZYaE3pkhdqq0/hmf6
0igiRSAaL7RAn+rc00na3MdT3eLqHrlxpzP9mMGTZ9rJuJ37tlZK3vUvkXXykyLh
y6J8KVXFyDCRWFwYJ12FFrpMqWwyOsDDcNSsVbKqmNMKgVfHsyKDxCT5zV8fKnUo
J/Pv8EBI7l6qKflfUFeQh9PQbUsBOytEbem22oMFHgcgmSqM8+5KXyPhpuLTMqia
x9pCtexeDTY+j9eBwnfSQXLVKgftD6VeWJplEGsbdlLwFzoffK/rRVVLMletmqi6
nYWpkML58a0lbvCkHuWcVBR5ejwWKrylVPnSoNqxJBb0jeANM2qvFEnBNx6ZUBQp
WlHgqyg0LAhGunB/FjRzVBdxGqdINzvg3OIHIy89Vv4WvoM1fW6fbLQ2G7BoSOhM
wrO/tG2IV13I9xbvVEbR6bjxlLEoUlKyQNbdP3EGD4Y=
`pragma protect end_protected
