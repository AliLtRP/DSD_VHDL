// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OuS1HapFhf3/jwVUwrSg7uS9ncPkkn1UxyJhztJUcTzaAgvTH3aJfEcg2y3kZCNf
dmWpZy/qM2ZbypnJvPmST+h4o7dnTg1JFSQ1fLn5NsDZM6S+0qaCEBWyXHG8aFZe
8DFYs7mPUzFwK5N4XM+CNSGjur7krUVl8jPrdovfcA8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29040)
JsAGiFq8cixAXIT+R93HHv0/DI+8IX95Fm2o/H8VBUwt5TZvSy5KCw5WazpWqUI0
ItydfLjUatmj1dxE9ZzkFrgTDwqpEBAJ+GvCXlme/udCpPe9o+S2K+cax3MRaA75
OfcvwsVjEn5wFKcMK+qibuz+v3Zjcq35kweMKtYs836BQsHidTNQYjDE9gUTE2Ov
qJXwsYuQsKnHUT2PKNj7tCY2ncnI5O97Mzrxf/tN6cBryzvnujaxeBIjuQrbgzAd
l7GYuK3/uj+24ydY0SbsUbxbuauXjOd29PVQ0DxKOlPJ4oD13lwPmjGFiP7LPKEN
Em7WOngvFm0noFKK4y4/SG7ono96GL0ZtMF9Xv+Sr6trGrpiKUEa4ltk3AbJKdHe
esCH++NqDL/AaG6aOFhnJmZVOq1s9x1UffXAF58fOUHYk+zeZ9w44M/vtuPCE7YP
P1a9sQZ3JMMudemKt6XcAdGwxP2yK208QFqx+rNLsFB1Cx9owfDIsc0ju6L6Vj2U
wh5jTcuW5B2kSuZiyKJnnl6FvkpffLLl5ione7IAZQMVxcLLqIClFbFykfz2IvB7
5T5dfNJdzEjWOknkqFVBRRxxBlXg+r8K3QuYK6mKpwTnBDk/UyUuv/m2emxsDUGF
rsmYnLROpSlblCZ1ojIytVDlJkiLbxf/oc/aDrL28u9FwObsNrXwVsxQ5HbqGb5e
CINoG55VHsc6KBTDC7YJXATTZoDCJfpsa4xIIt+0EVOaDyc12H6dSnUfOh7iZD3u
O5DrC+eV5mcUKPsHx01PPRMIIjtBd56eq+UinJlRFxzbHX23K5BSI6iXQ5kx1oDV
JS+trxeJWkCMZOd+LQFL4dd1oRRTvB+kZSqLTbdY6ZdBDL4O9VTEf2yWzjED++c/
TfD1pJJkp8NtfRF239J3iUh6LHn1S9u0D/2hZlyOkG1hANTLqDz7Dc5yuSxuBxnG
PBwunh/OecfBqa+7bBxZ/wmIdy5QF3hqWbLB+PqQZFSLjtPs1XHILPPjg64oRG3u
0Ls0l189zHMVlevmklhFa+9SyxChX/1BtqsTYBe+eDJDIbLO56tNDVrTYNqABTxT
Tj3n4636yEw4asF5rU8XopsUNwzOFyy7TaQzb4i1ERrRLFMQwUMxv6BH4isuklUm
sZ/0Sff6gN9IGRMq3/25rmxyVnaXn2wWgwQtYZ1AChyIXb+GP+/0Fnu3P9c2jqWS
pIJkE75hNyK78E0k2/ySY3FSQT1ja9k50D/AsBNVpEr9IJHAnQW3a+IzmD7ROkrA
JurAk8xSvCs78vOQqdEXrw7RuTrL7KuwdsgPGkta4Jpn4htOVrasBYbuCOk6n9lU
lVCY/Fyqiv4xu5n8LlvyfGOqOT/LaP2lKu7Aw66wPGOntd0eN3r7wvgYbcDZ65Tb
oGYIX4auwpNYZbSsYsh3tHgvEB0XaemUhZokrJNAdw37YpHr4tEZOfFq/QCXRVf6
2wO56CP7VuNKRI39kpwHU7AjOBuVnwjEE1mWXFb7Fj2JWHE5kie+1oYqvKqkLjIp
kvng+Lkc3EvaGnU2y0Bffm0S316M6w997Wl/FgFvJxDiwIjVHfamldipBL25DIdo
Wx+Qkg423M7dK+Rs3S6nj/NE+ENIqftISGlI82Z0eYdC1R+ED+y1F10SkPjwqvva
8l3mPMWG8ttMzS4eb+xU3rx0npnqtIcmiVE+LpKHELueMOFwbFiNhobkOzxxvKJj
Lu5vb20FA0K8oP9f7JmzEX2Kelw6ydaNMaqFkOI/08M/Q+fgsPgUNRfKPOUX5Gsm
giP/CLCXrhi4rFbJCDUHAS0IdhSfDTsC5gRzag5qY/j+ChD8s4fyUCcvrB5L6bsy
qa1uvItRXMXBf7zoz5w0dtHWxEuVu6KSihSc4D9NuRdUsfbG889kF1FiviKsQv1o
jqkzKKfnqvzu/z+xaT9yu4ChyNDaX+nrBkPRaXdr5o4J6kETcher9Eo4GAaIytVc
CRjLXLJuIrJ/nheVVTpEEGT0c3iPwoVe2qONfbSPArStFHLVnzrn/RXQ0XKRTDXi
3X+13FOnczxGrtd2wUZy7fXm1/yRIJqFdBlaOZuLc8BVDc6Nwv0FeE2GG51qLJ8h
eRJMcd+nDrOGP7olI61pA07NMMRPQFYP30afW5I5etwbUYGDCayeLIYlw2lb0hek
G+1uINKAMflGlTt7NZCyArymCccvc5WO35smsTBuhb2lpASK6T/Fs5YUPJw7oPpe
mlcDZcpW26JvY9wdzlsv3bB2TjumtzfXBAWusY/0/1r2cWJ3qaKNVwuQ9apS5Cl3
THlltyY0G6volVtqe5sQ6aE8I97CyKbKXW7uHUyGN3MLps5Q5GuqgGEC4Y6si8I4
u+giJ5aZB0bx2ekJasyCVGlo4jT36WSVScPBsc8EEO1HHaXwmUWgOQpL+wJCXSuS
9lv1QncecyFT6btHHnvxmNE/ozTRsK5hPYaeM399hvoNp6J4/tkt6YEg/TminnLI
ARWlVzai6wk2sz1DtOx+uWE9ucRtK0hmyI5HqHNhVazfBUErRTEZRxCcQJn9XdIz
5lQ0kiSQDzvJXYLJFEZzQQU4FzV/FzKDYdrqNnagmb1PpWIKwmVadqbegEpkAzox
8/iuhnM81A7aLFF+pqTAo5eOH/4o/beGbWRvSOwNfK0bBnwTc/iOAGz61Tm8Vn7e
2Kuj1IqqsbZfXorvBZdBNzyBaqDggJSO2OiplVZcD30BsdYIDEVHfJ/ujK3OtjcT
Kf6ubEsYaTo9V72ArMVuS7TPCuGi8PJX8q9BybQpirJrCtLuvRwlH7A08WQ84slZ
+tdFCpgU9o1Zl187ZBOf3yoC4XLtzV1eJy1thq6LCgf47TrwYIFxxkolOUOqYPY0
eT0ss6L8wSsDOMmZFnrr27guWIwSobVfexF4cSCaR7lUPjD9hSyJTB2hoxxj6/Yo
rQkYOhW3mIHSSFzisRvxh0TuOjtfzCvm89TkZ6xk1D8QWyVixrs1SgMpGg7px4Xi
rPSdSORvcnT2+wcf+Im2StXpnIkTuhh4dRUFd9UtCtqUeqBW6lb7AlKdCmwdEFl1
5EU4ln947WAYLUkztoxZ4Uq1quxQaAtK8bawPsSoMeec8A0wtnoizj4QiR1j10Lr
a6yTgZZD/ngmqQDZOoryjo4/mgeJFAWJ1GHZnPk6OelT1ihOXroON7DkXWuNdDUK
8frZLT68C8GCdCg782OPWKD9W7lj0DdoxKfvIjTVPqFzk8rXiOE84FZigjOQKqKz
QhR0KfnM9tTkvkhzXih5eNpKSR3KlH1gAhrL0LAciEQJsVKboLAHuvr3vmISv/hI
Tha1kiAfjGit0hWB6TuvY+CvtkHfLlgwcPr8K+DvGp9FH5d/R0ZX8U/id86qfVTz
dST8lyqY5mtgyr5Z3QIUmlMiMgKzmOVZsC8uUdcm5+RlGGhn/Hyov6B0eCBfHKAt
qyReh5yJSA12cUjUKOZqw1zsDijMU2u5qYbF415C6nd03+xfuDQs6WuOx/Yxdbpn
fL+rXQmQjff7P2q8zdY2Bp4t8ff/LuB+5Gs/HCFlLPM0KA4vFmb8va8Ubk22dbj0
XvKPaO4xu7vdFal0DmuPZF4jzgOO/aqpRZQT0RubTY4UabrAMnJ+bM1Pgpdt1sPM
Hqb3P0IJ5+d27Dvce70bOipJ8DxaxAdc2xYugOGFm9IFxvGnrOJCLOKmrJ1xSJZC
rTK8gea5eogQHzs1RAamPiyEKEtWTEQm36OsrV19zPidFizQqIJXA9D2wodcLDP+
Z3ruDgPtQwqEDHiTsLJFfidZ6cJXI9QEbtPciHJWzIrL2m7aQAq1QTAUk/7WaGOP
MyWAv49jzuWG4X7b/Ccf6EPxESU0O7Qgr44P0t2bsb0tiHK4dTiVrY3UF8kvWjPn
/tplxp2Ke/zIJeSD2dhaaBQ/gdgBFtmWaRCXDrXQ4ikTSMjq1wnGfoy0h65ttaKx
WQCGXfyBPoOQlTEVT6cF87/uFR0vP7kx6kIKmlDaxbcdAbjFecUwPNVD6jrjKBrl
rAz2aXvLyxqLu2FvUx1qVYS5/R+b8b0H6U6VlRSdhrNqSEzKvlmGuu16e791x4rU
FRMCyz3aJvCkgamD0TnZNLf34nj0nw00LSUHX4xW9qzxI1RFj635Ldum5A/u6NvJ
a6RFovRvcinM0Hc/F/2AAqOMoZOjXD69mgWBjR5jNaY0pabZ7lefmie69y4RbseA
9NdTVZN5uR67esYW56USWKhvaTw/BIh8l5QywREzBH8N3Yx3bZzYRNxXo9L8MoQU
d63CzGY/ex/3QU4YtSNlAVvDE++3ai72Jw+yXNFG7f4ZcdCtjL+BjA6h1gr51sgf
ESKLDx0p4C7A41IPDxlKR/qjgkTr9EoFixVD9Be9TVNVLpcOwb/ow1kbgTV/asMZ
WvBiCn/MAeNVZUv1+6kBQFq+BrPswx1DdQBWJ7n/4X3KHj7EG+jzpFzJk3fmMOsN
St7P/lhJR3JwloZa9vf99lo4JNAinruTqbr8ar0xCRJDlbjxnR3XSc86praWixYw
QiFywWXwsWP0lunSmupnogIOtwGH8cbvWpIkm4xX5Ft+nMQIrrnMmCHe5IYL2+3I
SPRJ1NQNUtfLSdWaxTYHTM+wHX0BVF9QfCme+wGaijmXFVOWgxGgQwrBz7Jr52oT
WmFwJaTKCdbVjK2hnvvoWOLb1iDt19cyrdrG65fU53DUY0IIgYLQe6vBLDFV3sbW
bSS7HYu31WT4QCExuciMDh+Lumkj2hoQprL8Djl1KDWIYsHw7Ruv4VIdn3bMTsne
m9rRZzJf9JcgY2PLYVEHiSvZ+b+m4Gd4L6R3ETdRnr1Rh+JvISbkY2HdpSN4d6+8
bnIDV2iHfCObxINt/efPtkcOFlNx7QdMv9zRACzvFCKE8/LhlbN9b4oVZdq6sn/X
uUdrFs4J92J0PEcFzP35GMF1MVXNpKGQ1BmE4zW3R3nqOkw3HWDUmX54aE13s3hv
3qibY5UDana36OOpY4DLJeHsOXZ6l9HWUzEfIme28yIQh2Tx1Bvn3Gw4MwZlUUXB
SbnJNMZh/xapreefaksA5s5QB6PUuvizAf6CBxdDQHuvADxncpwFak5hjBiqufaE
4PoBmdqxOElgsiVuWxYSeT7aF9SCfxyZRLQmDhw7Qm7ii+Y1Z59BJrHlAhEawRJS
CrDtojOYgqd9Rv5dMP878H4dCbj8Xha6axuTFsWiYNzutxtpegPZAi1AlfDg45Rt
8mH3g2YiS5u0CSkqyF7XmpYnStmtuAW9ODtE9ApPy45jPN4W7pO8DU2WDiVW3+le
uSv+muFKXfnckACE1NLPMvDi1L4/38ii21FBLR9uhU+YoQV+F3JbCIXTrdVgY6C8
tKedjVeJ3o5XGkdJtOedInctnRu4taoA1r9w83eiwh2BPgn3B5tzg1I9UCOVwlMc
1Ywq50e2w+c8Odm8IEeNn2BF35oSOf2quoEO2Bwn2IiEmT6NTxEQvPlYxpwZmYnG
FoAMUa1ARnwxRjGM9roCWiYYE9lSlVp9zwnXVCkgjSMKmUonmhe9JKCuZEIihXlv
cIrZ7qvat2gN32erhAievd5A5sqg45UM0Mzb3nZKufXTt1G9ulOnPLm5HSAvKsq/
qiX7Hv4yCpxTcTg8rFRXOcRE7AtAJUnOCjy9B4D/R9PbEXDKRYkbYIjNnRniN5D2
OeQMVzMDQh72ZEK7Ag7qfVOouCvnI48f5f8wzXEGknLrlYY6+eN4TmEVYB7FSlLK
wm310qSQDSyNdL5c4TWjpuK6yc7HhCo8ncG5cORSaaxS3l5mRGBV87ydSS5PpTNU
L5MFVPIRDhfZAQi2ZwPhXe9xX2Zb7inlBuGZ1jW8BwD2GAmCB6O7xT1wmbozJFDX
Sj57oBVsUoO7OUYW4hrHn9/7PkjccIL5CxY9zPttMFP/je2qShiHiPCkSAGIhATa
mrk3UnzWwSbdoidCxWcZC2l6ih4r39PIWMLAo/U0AgA3aitt/r1nj0aAC5AYapme
BhjyzdDhvsekc1DAR1HRQsntZGWPRnBvz6mVBxQgw44HLcG//KIkbFExZIQkYr/E
7oDG0K7KL9VVww4eMnQ6gggZ5MXeLicr4r9Q0xpMLxTmqz5jWgAJEjmalkbXmZNh
P/qxkQ/e7SLYMmwcKVGt1sMV3rU2XTFvT18m7NArdoQMKhTyKyyOzALr51W1gGUI
+G667QXhjgzR8OnDiWs/Ymal6+YLnFoJqJ+4f1GfJawnh5TB2Nwx4KKtxsgE6hoI
CXdrvxBjNdyY8HeBjg+DJiVYTrc6Mn7K+wcFiNYqadtisR4tkSYh/0hPLkZPaALg
cf/80BxwAorkUHW5HnLmMCG71459LcDbtS0WrHaIFUWepQKtPS1SkSuV6e46ZWxE
NU/myuuChgTVeogYS2jTLxLZeosZdaV5e1Tm/GjpGDKH3GejM1geeYaMxuxnd7qu
UK0irVBkrg9iVOAtmgBQ5ntYGc2t+HLALkIgepN51JQgzVK4n28eV4rqfhD1TyGe
YzbeRFK64PUQVmmBPgVjjbvRx62kir/KB4wlNTiRnDP9j8u1MbGIo+UkRzNogtzx
viuhUAriGVEmfQlsw7vVYJii6BGcnB4wKUG7F2Yl5lwHaui9epALuuhmpCWVJyXE
sMS1Ia6F/tXLmKK3Bah4B2ng7HI5fmuBqExZT86bIUgqF3AoGFarC5xu0sHY6r0p
fsSPWjyeMByKautZuxyWjiysY/836nz69UL6JbJh/r1YUIKudlyAzf253MZtbiEd
V/PW8naedc/vj8E5edUF0ysQQzLv7Iinq6kGDWWCVjvrPgi6weORM6OOKpVXoRGQ
c/soTR25fBwQ4maww3ffsVM3kJTAI9obqIWPnRCV/fq5HwwKGDEWPX6HJtw11lGS
GokbGOK+frh0qLsBvG3wlQNYCt9vwD5UUeqRGPdFMRynd4f6g+B2ngjnkuJkQYE2
v2PDvuhSahFzpVJcz1ziJ0CZvBhgcgGvb5Acot7YcUnXa6rjWvcoIos838oIOIjR
OUQf0JFFtKWTHQZfpnWzZ86QWai2Am0e9So565fRVKeO+UKKNjoBCaRYmuMpJVem
GnA43IwsOJste5/Ku/8XonQameMZYzDOh+7dELSdz27tlWGNxaY0QfuCQaglesmC
/Rn5Ldx9QXh3RCOzorOg89tHFFnY54RJHFKkU0CrE6Ol+IduQyfDyelUqvxTq20F
yLYmkzOCcmdXKo6acATfx8VX5NxuCiOEO92juJhKWOFV6U15EHcDWnJ9fgl4kTXD
H2M7YaPsc8FN+5l6KR/nG0XbrKhOrPsbhiSyvktRiTSs5+XkQhOMEMlEgSDMxLKB
13iYCRESMZbez94cwHEVEk5iwdpd4pfv5d8mm/BB0X/CT0EzNmOeWExEPNBxkf04
UvtdI50MWWqlPcZISsgISoscAi1GSI4LaW2S7quM/SmqjdyOOjY/AbbagudtB+nd
6t2my0LoPTdh0lNv61cynt32lcFpqcnT2O29Uj8dt3w3ltrrYg0zZHJSDHjq6rlR
/4Prh4pAkbqiKwaOG+5OZQKvxL6u/CFeG3zoEzs7+J5+rZEbLyt8n79RERxkQT5M
4gxgSDYJsoDqLFyGOaL5rVDEDkIbI41wBfy7+TRj7E5aLKUtFyqXMCuDa4a7mCum
H1iH0HyCZX6z4Uc1zIBwXNxEGb9mHFLk116+zwnOPFKXU/d5vgGPbxcBxMPOO7F7
L9aF2N/3zx5oq+3RI4XKiVcKLIUnk3nmvw/Rt4k4noOvim/NJj5ujT/h7CpjJLjF
pr+Fl0d2GoSLcHfF3x/vPyRFRlklzXfk+1D288CPNw1BdBWzqEAZUBmX/mvXZC7X
WIEyT/0vqcA924l5XaSvu8ApHueQiu5cFV35TbGdz2vVx8Rm5j8XTq9jUJ/08TFr
lO2H1ybg0/x5whmtaEpvs8cpd20g6BaoufW3PT5nFx0KW1KFr6yTMTMDIvrp8j4z
ZZ+X+dz3W9IliH/M0c4KLDu0Ed9grHKviZWTc23Vp1KsM5rc/t/TXVcmHKBYglCm
VXn9klYZ8so15nJbmJcE2PAfFGnKdN0RLIDhQVdnZ9S0hpp3WCprjNyj7RE2ck4E
Q2Tpx1s+jSL6fPzikSA0Xsa4KAoSXlJ7Qt9vykE8oa6rSSOXgW7JuDEaEn78E99s
QcFXpo5QqxyrEb0MbggAZ+mjsR/6ZFrS7TfovBmTTS6f/Z9PqacwCD4jpEJzQL+r
Xms1QH2f1C6fzXprKoKiRYv/qxcryV75LS0rtaeDSGR+84zRP3QZzrohePATSrtQ
Rtahg3m5bqP6pEC1qPj+v1F2Y5g+RYZr/knZS+Qb1wLAe3c7WLBkZLZp+H9N8Pbs
eWwZtRiRUtU7thGNRZ4DyeYaMuZpIdXcHypdqWuwGuwn6o0mQdSVwvCX7eqWAbnT
HqZmNrl925saC72pgxbYcpG62LdGosBezqghdDnLnjJnH13R1OKA2VuOmHwamOSb
IJikz1uivIVtA4fxgj7WDT95lFgeO0F2eGRacEKVMQUg8InLnLInyM9yWfhgK+OU
OP/6vzVQ0TVjFeV2k+byA5Lpq8UD1v6FO0bDKimHjNBLZz4icllTXqChdvEl+HTH
EKRVcPKg36Jc9RpKAwUaUokrQgcNUZ+1kdRe0x0B6x0VqNjIdAjbjENbDUNH1RF7
0d98gifyf5/ydmL3sf1ipZyMCeQWdI1qDzpJrblU0sqfNMvF+PX6YgIYb/eEPy5H
y6gzLHJ89QNXDFy7ydywH9C3l7aVDst1rvzvlvtyROagrg3VgfIhUgT0TkVZZ3Ze
/UfeLYdWmxn69tRO3am8B1Lmkawr8a+hmB5iEF5HIcwhW8aMlrWefjavuL4dFnhS
49Y8Z69Rh26McMgXQXh1+PNlhOvaon3GJXkUnhivVVacreGPQSiRAO4uC1yPlbsv
Smfm2RblYtU81cdfloPAh6L71EZHDpgQYIdzpdViMTt0cTHP1QHtQAiGOBxVMnsh
440DaBjpGJ/4pEuAlPGeufo4bxu/lSQFRK0MSjMByOyU8Uppc0bNCKYb83dQ2lXY
sGqyaJuDipKRLkNdBDcwdNSGIqQDu9izZdX3zuT6y/22XvPVVc9QRePxhl9ws5RF
OXOtx81cBPov92MtxqNt2iVIKMLk8mjAxXdsvnz7Z/pYLJILFD301UosIDemp6AZ
2ybLKcgqgjfBcJ3anm7YO88sb/Kx95BhUUS6EEY5I/ZXNrXymZsXyxK0bGKkmq+M
MH/E5BuqZloSSr1t8Gae2Hi4ZZXypnebp4ha9sL6xf6ndA/UkBNqf6sc6Z7H9pXW
kM/C9ItjXHuugrffRAq0uAyzVjFcrE+GGyUpUgB7L72Qu9pq3jESj57hznOgiD2+
Akhcjx1fWJTJGvYnD1YfdiTetSq0/QwAqOEp6kaAy9xl6qGpbqrkva85a/+VlH+q
BR4fgN6xlt4QfalwEbgUb2DMwnDAmEr758AF0O9lLQPcEq7oZ5WVLvtjgHre4idB
Y7qf8rZBwTntJtXdISEOch8Y8KwxEhbFLifRLq1vGZq7J3Hy5xELT9nDhuaIzM0Z
sC2eagU1UlE38FDk+ca8HIYLmhyRbT6Hrj039didZwVjr6xHepsf20yoXLV5p3Vb
x10RYrkzWwlDsyzWyTWmd4r3zbu9qT5H34TjDBZGST/JrdUdSejWOy/YQytPWJvx
yvJEwSjFBfgI5u3vxDzJRYlhQdSI8OPk4F/RPgEKjZLL1DeSK9aQFnazWvyCF0xH
PxAC6RuTzoMQ9xrbzC2zsyyQzdRtE5ejrvaTsynhcvAL7KvJ5StYOmqNJ6fE9AVx
3bL96LmrKgH3Htmf/964fjATTXfb2MEz5h+Df7cvs42kNrDxO8gzpE3vgFm0xnbU
bwawllg0XSFT58yQX81AgtuBcCcctyJDYN3t0bLVAfqr5l0q4Li0TrhxO8ZlpNoI
HxRASYULvxJJ3xqQrUS3n/XwUNWm4b+8ZOsdRytRe34ZyH1elJtbyyFdIeBWGWLp
Qczsuu2TotMo5w2icC4pMGMidro7/zaooHeq4KkdrIIfOQ5SgjTWiGvF9eqxzNEu
QOy9IWxtB9RqlCpXipTuBnmo92+2480BRcaHwPF+kkYJHny/QhVF5Y8RJsWuypQt
pEwTVwHUutRuqn0fIDKQnbBiT7dsMwTpHsAM5COvlPG/oeNDmOXXdRjsKp7D4chv
3NwsDTI/Dk7Wpmbuz+Zz4pcLHnf0elfy8wqit8XNI6jmIqxNMyG9QK04QEdBBTcj
NvMiJCXaA6xdKp3y5kdiYNZzlUIQsNPi0ha/yItrE+vxRd0fJi4PjSqIs4qivYSb
P6GQBpQB7ZV7qtVxd2ZULUqKWNz+IGg/0zuUPQoNEpROK0tkI8HHCDQpYCXbgLpV
DyjHLUupQrk8vUApqWNnP1DNVfERoW/hic2mTc5aqoJy/s7SkHcaMl0/LooS0zYj
MCFFkF9+kDAIZiCtanBmU7NZvQpYStPLnMWiU3leHZNYIxITzjSca3/TVMpfqKya
rE0W6rL5dB52d691VSOg4Bg7vtiY5RKm6bxyKTrbffGSJAmiQFZVwnTUXDNVO/He
AhSNDXgczzbBczkNlXhIlSV+LlgFe3ggfj9suGW3HQ5J+pGxSsm9moRdEc10vdi4
QOWq9W9M/mlshMB8mEQesZS3w1ylbdpbsBNE0fYojaKOQl4DbeItlA6WstS8qS6w
7U9tD9kuF8Ovp9EN6z9tTK6U0Z7q7X6ikj2BZy3JgBux9YDuKyrQXjrNe1XCR2zf
BK3DVH09CeI8oiL9FxD3iOlDAbQgdNh9kdOfOS2+5JTkPYNQPiUUYhRomtX/HbPb
tnCFxqq+1Mld6HXKknE8yCkXwZiodFTZppP6dJIzXDGufQNn2RW4ObVnp/pcxnYL
KbTpnyy8vJafcw2NIOdOJ2BnbjfrjkNFr3VI56wrqlsyNlnD3wWgd56TWQtOo7p/
erhILYjxcsnP52k2sq2KfMK8wbSR8rbQAsnCPUY9V7SBZg1NhAKONVXlT807nhRX
NldZajCtdniiCUwMc6XeOHFys7YNA5XC5bd2m0kxPrBvCKsDtg2N72fjMG619Sk4
s7mSlI30nMoos+wXXUxWRwbKIg677JbiTm5HKPZ7dkbDBl/Bp6N7y8HEKLt45tcW
bqoLOSaYmTxJ/Cx1hWPid2u6XGB3dQUKhFbuhxtPgOzecu/ZC+oUeWovhkPXZHw5
bnvzAAPqQNIRRMcTj+eEZKvOH3ypcZJJLyko94hL3Q+QGxjgeVPJOwch4Tt6fX7S
w/GJrdrXwwWlW2CMC9C+0JUtCDqhSnqfumk5834qfL4bl+peHqQckcaWrdItFyDU
nyzAeaIyXr/i3XEdI6pAti/QlxydSndPWsHPuEhh6uqsQ9IVPEGVGz/ccWDAtoO/
uf0SIM5+6eaLVsxaGI00qmfMvxmTFXDzmTVqHBOTbUIlDGyINBGn2ZclwB4Db38N
r7lh99Si10sCybYhp5oE8g8A5LM00eePXUJ8hz3Xso7PXz2+0J4vrmuuj3MTe6/3
b+tI02Nov0je4mBH5eZeXB9BwT2q2PTJW8ysjGkd1R6/d5uxbjgNNBA4VHkCxzng
50F/PbvN4dcWNMM7rBnGXzGI0tb9rlO1HtpeV/+LZmO5jcerV1xKaFoRi4RHUzwC
eRNZ9Fm+uEyMLWji6hyFx8vo313s/wi7KlEQzdk9yWvLskx49GpsGqeFBc9Zxc2m
qvY4nj7gEOROi661+/WJr/2YYafJB8RVO269bWjj66Xon91m2llrAO8IngKV6l2f
EGreX7RRwGPQgisCS35oUXMNFFN5XEWNwppPvrt5sLNLA94qaPaJ9dAzzhv9x8rp
E9vtWvwvxtla1B2TYGdHpJJ5HCoiII/OPR9EA6l8HxQMmIHr9euR80crReOkJstf
3NrT2zQLgvdkbOd3Feu/+hOTDPFqRcRsy1OxSfLM65Uy4Ns7imzHrLgXakcf1huv
g+RhUyvjodwTAQIk62ewfn4Fc6GVIHNQS5jt8H9HDl16Y2CbZP14tmFIrYhtJeNe
ugdnRmSozELYf/H9ECGI1sh9KO7y6rGaHo+JzMHQdN5v6F4lT5SfaRvg0L2gL+PN
YN4cu2ujRVrlL9vTUK1Oa1CR7tMnT9RT6AqiWa8ZFiX8oQaJdWyh2h9ELmPCUP7T
6qBxeoZ7SJEuKLdO+lW1Fg9jYDOwM4D4Ftad7mZ0GvrsNOuZ+w3BA0e6qn9D92I9
08BhR2TVn+hpEKpMkBtg43fhczflksXLyW14Tk/a0jdremOcgvLtBQAY2NJd5VTW
wr71kveRCTEiZ35wAMHKKWXnqdreQ1iWfsv1GKMK5HUE/mWGaYwqWppDfpYUfAZc
0xC6ZAtEhVRJWHUvIlYNOI+GLlM0RK99JX9iKWNSTxC66JO1LmLREvdV8CR5uucT
/sVAXKr/4EqIqC+w4aCtyksmMIaaEH3JAHmWXPTI8ztQ/qjsUlvgzkgq657opErf
qNYFXME6oM/mg94Xl4rAzAUk0Ba3T5cws30RlJBalJ/LGeozC2dZyDMFW15/DvED
7e7u5jz+ggVQs4qhLxaqSDWFNQc5Y7O+Cem1ImDg6LApFH3l2bnnRxeNXbzrDb89
8B2XiAbtDi8ABJv9QANLV5aE/gVIO/QY6RhG8F94Xg018HcMprKmJvfk/GOSQR0u
JiVoGh+VvMSRUIOHqSr6JkupOlKs9Hy863+gLKEJQdsunjN2/fHdFGZdnpvPyBvg
JZCB0LDzeDce/P54+kPI1RmbtkbuDJqeH38+kKK/WrHHRbL5pHTwUCnHNIIKMatT
U0uRMAdDul6P9jxKmMeodgN/z8AW88176ZEMqDPT4jFrJ/Gj1G83l4pmtdcwLF//
vm2330KdcMsv7p0aaW+gMIax/NnotQ+Cz8VxdbseRM4ajfmrigkrMSBvvWXGv0GP
mI8m4KquuPK8vJxX0a+EfM14sQ/d/ugQBV7s+v2CqApilfTG1GEhs2lLEXAITzPn
cELyXeMrP73ziTdbkUWVXgDF/0ZhqkFJc9CfPdKywv7THpI4YiuO5CUCygDgGm8h
wLccYIhqEyTkejpGgP/dlTZkwt5DTNbF2bxGK3XX4AJ5qdIdaAjEgXnDfo6DgU9P
tWkFTUo/KLAwuJPAT0eKxWALnJZMar5s+1MXeg+b3KQ4mlJxGUa6bjEm5CeZ51Pe
jXRjyTPioLBNJKZi0wZJlXblKH8IRjEVrEIivxRqmhWSrZvManjYjsAkr6RiGZAh
YKCor29f6GdLc2+v5jCzoFBcaPVEx4FRSptUENfUwSPC40fFtmXX4zwf+FfLtHeL
v0hATWa2CvpwiyqG7v7dGRZgtXjTyHNWgm0qFykKhiTm0YHZ8LDnNyo578kKuECR
+DbVO6hwID7XP/sSYdprxxlIeGRraEDq0kD3vncyIxfj0w3DoTEm8uUMsBhiDLMp
09F1IRlQ5jtAS1jAbScdgjAKIGiKYDQxeBXta9h5TlRvX354m0c6kd3HK9ztmF6/
NEamVhxKjmuYijGR/ku6BmiNyPgcZEBcet8URnBiSWXvy/J60axYyv64lQ+WoF7E
44BAHmqVjuVeFebT7SL2VwDDfFuiVZRt7nQjeZf5y+PFeWZVc4S1Iq12o07aTr1J
QMDm5vR/9Jhctzo6nvlfpJIQAioD0DecA0Q/drMJUQiuPraTEBlkORRaQmG0diqf
rPUJOX5J69dFmQS09ji6rLCYfaoxTWbuxtfw63Q5bTBGkR9aydtbUGoYzDP6+AjG
CxlZ97tgA2tbcHJHeXNiwXA4NS9F/0Qdl9DnFNsr9NPVNLu6iHNA8PIPAriaa7qm
ABdnAoBgCN4dcRzEUK4Lwf8qM1Dki2lxrk1KQqNszEyhmTawwS06/anj8C/KQ1ak
y9TM8MoN3AnugjSb/nZss4Fhwtrw3infpyw0KCYPec++SGXpiG4TEMDDBbnq+27H
HlERuG5OPjWzHIOvHFCeg7xA/+wZBcY0Tf4/hrJzsHn6/3vk8G7cP+joxG3t1EVt
LHwr/z6MUy+HwI+RM6HqOzlX3dK/2e2894KbZCI2i9/AZ1OdclFb+xD1xvXlp8Bl
m9Xavbuv/ABLdeLndDEu2VJca/2O+7e3AvlCpZnCv7ewiJcKAaD+RkIyjWiyh9Dk
g7Yi9jvW3dNMnGUgsqK0/+R4x0HKXHql24Ur8eKbh1M8kwIp7IzCHYsahsoQhAIp
Sj35kHkzhnORKVnkb2SpV4ZnXCTSSmG7D9dq1Kc4LKqctoJ0OpSeiu94iZQX+DeY
qx2T4Nxg4zlHt+32fGUgRGfNbiytYdQjhfiNsWC+4DG+WpDugSYQNSzRFhQZyvgA
uu3KAa6PlpUKFuS3Tetl4tpXCpzfBdmL8zKo9pQGNc33jfX60yQPLSijKMhaeOzT
PYHDCfdsd2f/xFmY/cyfmURXJFDz8nt3iswXZewmAU7Ue5FMEDapjjVyFxE9qmYF
nT4ah0mMsODcYmjaa4cjVeDQYj3axUMyXnlSYeX5AtNEuQzHyw8anRdmxD8PX2Fz
/NjKb3DbzQ59NPGHBu0CpDXsgOndZ8y5G+Ho877M3lv9ElMxcDvO+50WH+SxeP4r
zgbvUHE4ij7xY2733DUdK+WDWyUuY71lFCeIT7zZQi/WZVJ6w3EM+fefa/RBEb+j
Qk+nK3EN6dlRWj00Odd3YGBHkDbTF4QevZ7rQJgzPbDXJeiZ/kXZzYiNthv7Am8r
ek0CbGtk+CEc+CVzxmDIu0/DCStP33aUhcw+PRZH6EBNmUyFyRUxsDSVT1fbxsmi
t+dMOmlxMiWTy5HwU60kMXeC/A/QNqIBvvTu8aMaRx7aA2Hwdc72xd7Vl7vAvMQm
fjCQwVbco+8/et7Ird0XC3EyOAMumqUmN0z0AXpfHtaxjZjUtxdybBn/wV7tPJJU
p2c6g4dDX7bOdOi1IwIyyTlUoGzBWoJtb6VDrmVnRcRwkRi0E+IxorK6cZyCWVRf
vhSNEWFgpdEyPVXyn6kqkUtBOs/o4ZnM/2GHLo8EOjR0na57cQHZo6nYXxw/Qk8c
BPTSiLvX8wa/PBFQ7FfEfUgpgIELXormmf2KH5Q1hv3o0Nq2zy0YjxlWFX9viUHL
PKTx4YNfhCLqgSU0L0KOZgsurBSUxRZCZpWtMUZHlEEUh3SnM0Dm5RR19AxxI0V8
yvZrQbvo6Pra5aqqYrpJPPa803u7wTjY8doDE+tnADGToky24qJlpQyOfiF0BfiK
vlNiolqtnLIjBeMmVe6uGtta6k2v7JQ1Ha3nppO61tw186Sqj2GuRT06ILD9lSyO
wifwUTI3rd6qUlADtn1x9nWxRCxoaL9DP6VkNX6GT17xAaNTr6JaDwazm/JYR7wZ
63JU933+8NY3cz0wDA7LRrZgCoLLz6TyAdEylWWH5HoBLMIJ29X9x1/uCjMu/ayw
OUg+/1L3bQVp3694qhK+jdch+d1FgOCAc+Y//gzVKsvMbL1vs7EEpnIce07xogcS
7KfqGgYPF+/jan00TrUlLMaaFXsVF79DDRL8HnEAvvpf5zg8wG/A3y1nin1/WpMP
ZKp9ICntG+GZ30lCz2xXN/I/yVk6hiVfv9ICkGUVyT5XcJ2dq7GMerlAVrSk8KPe
qvUe7sVxcDMoRV94y8aGvY5S52VSUUQITRBdUHmtV+ZaYcu9kcYTegu4m2Gwl0NY
o9IRGXlM1NQnEQv3NmTz9s54/9f/D3cbfZbbV6ciKNL3P6M0ytSTEx8GV97UnxHX
ERLXgMwDZCZPniY2RSva/qjWMkRyDm1H9Tzthgy1Oz3J3foY0/Pk4CVHDKA3sVLM
1iTXZmIQ+EXE8+yfCJoxl3xmF29GfAJWUM4dM72ADTDjkp61EXJTGwbPBz/fdkzc
qo/Bv/VSyBVx+5tkCIcn2JmslSCjymMP/HBQWqvT/5g8569r9csRMrA1nkNSEyOU
A9qs9WJAdanUEFpafSAfKSnQlRd7c2cVvD9mX1/WvQmjIGrCf4LVsNCLWmvn3ami
mddin1hChLktDYcV3H/bZLr0Z4lcXkcei1U008kFpfIMzDQjAkrXQpd0bqUM+FRo
f8lNbtRMRQhN+UttS59wW8He9Bjtftejc1uDXubUN69WpMVBnCqrT8BQmPLNYwTJ
oJ6nNat9QP8aaD75sPEEvMfWJ0dIowDt58wF2naMf4pHnU6QVIkz39yuGRBy6VsB
CKrNiweqgizcAoKlkYQ+PUbLiiVfs3i1SVXP2EALPpsSgwnQXNpRSxxl7mM+3uTK
VTh6KFsv0j8Sliv304A6tSHsHkrcPuMcuIlBlkCW9lE4hdqtqk4GXSXB1UHgleMq
goAOL2iHRjPVVmTRD2sMJUl2Tf1os26R1sZl2E2KnuVtcdy3w4v09hhKgm7wnKjS
sgt6sv2L5Ho3B94qDH8RHaXLG3bZtXLsC5WIuvXadxFJuO64nobeiGUxOQLsWPCv
Uo/mRY3A8sHk3FICC8Co9PIOemmtgvoOxUP0QNteUkkHi5CEDPsD0vnVcofXI12C
faDlO/cuSWY5M8oLI3mlywO6gRW55i6ui/Zmb3sGzvt4uENhW7ulVErxyIkV4PKs
PMZmKJg/Dx2hyI2IiLRkU9ccpd1REp4lakahk0VBQd6E6zw3iHkJjyevn4JRrzv0
/brpZ+fn6YjakMVmQlgGVbMAormQlG8KyR9eGtlc4foatg/CAC2wT4uK7G2LNe7G
oLkVgmJGJfDS78D0ocESmHugrrZbWm++ZPVJN6Rqe6ot2wixS25G6295/NsCr++8
uZDiIn2vMCAgGF0kb0KOgKg1E20qcpwShUwOfQ8j9VEsIWjsArs+iHAgbldBF5aa
G1EP/142M56+Mo+7nVzOsA1viAPJnKEhrH9eIb2xIB6TBxrxHq/osmtKOENxcphf
zFlI9mbgp6zJUUmnmvlOpNg4rbPfQJb5krZZX+FEQ9AOGzzDEzAzrWkRatYtkkLL
wchJbZVe6F8wTQyvWlIrqFkTvke9/ciAswkx/bN2q77jlBCvjrni9z3LmU/sTyJt
+J/FzwyRXQOqupTTnbKHgLAFdLDnsNxc1KAH7W9t2G5sjvNLd1mzjZK+p0YTS3v4
uh+TJ0X7bmLkZH6dBMX4rz7o14U2eLgcXUMQOzaCy2o/JJMK+O/d3A8b1i7qkQKe
BPfaL7BepyJTecAWlbbOT4ASrY5lqmPYbxyp8MlP98TntMcQuwa5iPTbh4MGFbKG
kUHtUryMSjnhdgh79zppM0WPhtejXVkz1KODS9e1JIpkiNKA1AgvXGbszPClF2E/
Vo0W+M/ZaKMmB1epOjJp8FMt84FHpWNH3UC39NAcbKed7qxHo8xfjpshxrK8ya38
4EpoWZtve+dhyJQsiJG+Y3XXPyoZlZSll6Bqf1kSOhjCUGmoJzuRx6GLp5mB3e8O
ELh6Xa8FG7e6KM344AQxQ4h1cX6pSVQqEF9cBN9ldKjL8k6LyeyoWCvL3prLwsgy
b1f4c9uGh3FPhDyWzU8rgH1paycFt9ue8nvLuLQa9E8jLNprbH5bdtb7EUGwUQ1L
UaNXXgSB+aV+aj62LGwZLFTlZ4wOaw/ZiC5MsYXVKx10d2SLz7mH+82iwavAyNrQ
G7n9id4i+q9nMMCvOUy93DyIHPtcv5FSF8juqviUXD1NnVsyN5hBZDY1Cxd9R2ED
dbWJkpKJbtjGUWBLj36oViBq71mKxNN2dH6DWHmPZ0KNMtwgW64NtGhTD5h4JDXn
9kWlquTOHlcxY/6VoMq9dWJS2IJcg6AUmC3lwCka880q8uCLqn9ALLZfBlWYsRDO
Y2w0379D9O1oXHHqmPHcjNLqsqoMOK4uQO8fekz05Bjtz3Ep124sqEUj8v1Sc+IA
QzKNOOEeRQc2i+l7xjsBIS+pDk3ffbQMaxAD56EAp7QtWA2OhnGoa62B1kP1B+Cs
qfY0MeV59kgeANRUowm6vn/F8c48VyirPzKDWF6oJmbxNDg/oFmFgcWoExDNFlx/
fTbasInXtMqSTCOu0zIbl8dvf0ihfkvOS0/EjxgzXSgh6LxvISijOVlvIwWEpXY7
EUafWiBv7Yw2xgr+BRsp8CMumifPcShFOMVtE0e4QDoQvJmLzXEo/kc5sIbBF3zQ
lSTG+KsEB0RJHEBs+muTYrAH7Mh5qvZ6Gjs3wEzWD7Tdsq4zRho2WmiUkdqPhz66
z5h95IUqt2wKICxkExBS8N/r4MfRVQlwnBwAMKejAnovTKrVQmh6s2PBb/6RFoV+
ym/7A0g8ZUAyJUmF2NsqmdSVq8FucESCP4OBB6iSV3DYOoE8ZG9UjQNDXcJgUro+
5/lQB/FSx200rehZA//a7DlQaJqlT7M4f6ZpGxihUuzkrKnDLKgYwCHqtWCYjRcI
JKTpQpaUDktWpY+mzc4/u7ShLJ0UYGO+M3axWYt6h98GZACizj6wC+6KQHrl0yLf
EFtZMMrZr9S6OsJYf4BAZPy7+7flDERB85tNuihaAsF51NYnDk666W8bb6Y8sZsJ
/2xO0OuFeF2PImmoeIzu3KxxbHVTU4bzFR3YbWgGxlzIZWpwCy6gPEhLn8GUz/Pb
5B/M0EfO+H2QGQ3FgB2xOCRvAsdIFjht+kg6drUiTeoK/F5mZTsj8P1GBVJ90d+N
TG1zMRaOKaQvJs2AMW1UbBeI6eCV1c55OFgv3m0X4N6fad6YSoaue+hD9mG97GTy
avDfsqxA65dm8sUflOYrFE609hVxHUkz/88HxqKl3KGeSynvf/NvVfJWewjA6Map
BjZAhrC3Zol9M5uYeVuhdoy60pznShHLVBaOrkOa8fw89iSQG2HZVA4zswpIayUg
UX8e63rAD01NWGfKdCPcEiTpveOVwjdpap8kZ4i6G07MmiCbq3BO+8wHiGk3X3x9
8cSz1fMSdmoK497ueymoBqk888vm9nXUqf3VYrAP6YRjJhvfvdM2NV9ykNjss1/j
TPt+3kwXD1+NOdUe49bM8TVmOcyQ2JR4K7kPL7rz2wmrQWU91UVQO99VTowCZyTL
AD6cgBAQjEgV6A5udaKrzs2c5walkmBAV3EhDJ9nidsYFK2bzvQgNgNiEQuOMn0u
vH7Q/qZ1t4rdpP8x45JC6sc1ipAXYMw4SM6mqE44w4Z7OVSjxVI3205Is5yV3HiC
7RMLUnNtdoEMW5XHN04g8Dap+1nBQyMPtHNBsgomxntu+SsqgenqWjo+jRWg5Vws
SoeqphaPbfRIYK/p634N1+stkVQV4AdJxoT+WDT6X6YCEGAKCPa+tOUBW1VGI07L
kN2f4x1/zBZYyB0X6Y6PJE9skQ+TVHcdL/yWD5uRK6KQEw3eK7jx3CEBmIO18Fm1
Y9/0NURKykqfCZvu7y+oKW4jcThohr3o/OH6QN7ctSjEaF4h+VNaguq2Mv3UyxZ8
+SpUVubb+v1PKJOL4bHunpVevobpcZXNagDSjFNhamlNJxnsiaYcXY6p6iaijUjU
kLPIUP7Pnvd3gfJvQi+MNyxrrpFjL9D2vrCMt6V5YFQPF1zpCHQLQEYeTcziCd+a
5Z7FAWWlfsx+/685QjbaRSk3Mo4WMTIjpdqiUCpfShP6eXDayw8CX7cbH5n1h5ox
YLYBfDWykKSvq4ZWXZ2C9MkRBd77hkOYufIvZapljL6UD9T/K4c02GlZtMUvWfpk
kgez51Rk5O0aP6N98G/OWK79Td+0pTc6udcmTbhpdM/DGHOXVR5vlTcxk2Oz5z65
k5rXdfI03rEYh6ZHkG0Q4JKy8G54/TkQdyNJIEXwNP3UaR/yB4TidAXraJiqZeI8
boZFLjU2tZ7H4+CYCxzMuYwHWW1YXIln1Pr5qIV24KXeihZAYKfrY4tmc7hI5CkA
7GQw8QauK/5AVrq/o1tJzcspEsD9fliVWseCjCQODyTum8Ppn+5Yhd3J9ZlPfzS8
7cGqJZFnv1OsjaThuV6DO0lRzB3jTYXkGENLbG/9CJKJ3egYgn7tXRI5lmerYl0+
s3RwDRPLjspP3ms4mjX8OzgBohVP1tj2aJVKgLi8TbsykjKshtsaYQU+4JTkmLMS
axP6Ub4P7460bClRDuUQwC/v+laDF8yzcSGlO0hgRz81fbwlpW+oyZB2LL2zfkrL
PIffxLuUQXx/9byf3vDpjuJH4767YVGwxopoLmMvOy+GVEZp1l4OdCDqjQloT1gB
HyOWrErV5EcQFt1oDu84v2SLOJtGPGF39zqvBXV0PLxoXtDemeX3duTJF9OY43vY
8iKmvPlt2RA6o9d9o7OYhTKBZZAR1iutyMbF6UUXXclvu4s65FihG8DxjzqZSt5A
2QRx2Tr04JyDMK0eCpHQe5psKQrgeL0Eu1Cd4DWoOA2d+ks0C5rEEOzxHuNscrT+
7Va9tamBAL4giKt+KGoCJWgHHPE9h6yPZ4isqEsaxjQMMFYT/uBhd/rT62OLTXm/
r5GmwGbv9ctPoIE78IW5o0DxCYkQHJL0q7eBA40lmN+OuD0CjRjkqpOwVOIc/HQh
Cz5FVWVU7LnYNXS7HNcEaxPbOQjADZgDpmm0ZnJtJdxhM1BmCdj5F8bNCdmT76Y/
qCmKMxim/lIvAoUX7OxrPnsOIq+0ZX5b96ZmrQGBlm+Og1UZ2BMx1pSYB+gDhse7
5S71XwQI/i28fc/bgEkYQ4geU9o7uV/7fo+XERhZeszJcxvP/bRL5+2uRYDF2NgH
Yn8fw5JgdLoC0xHk4lpzIHew2cwPoVlHk2ukuZKYtX4SAVrRfaeR67hh21XV8vRC
pRx/G+5lWKtGiP7hXOu0Zp9fcx0dRLkxDGx7nLDeEh0tGhbi7xBpkpyAjWy6y1te
J8GyDOTWyZcF+ihtjJi8j1aBz5aDoD4KQEDn0dg854muW7C4hdrUUdcMEKlX2L58
EuPmcX5i4Ndn8C0JNtXR52eKAoWxDwN14GpxWM7L5vu519hBdtpeCX8jvEZ6SBG4
5zmY9RVEMrcKu8pmVWodTroanhOiAgNM8pGs/T+bOD6rIEk1aKd/v4zxfg6gmhgL
8/0FoECNUsBhBlu8UQHkjlRzl5EPZF/vuzHQdYQ3YMMzwHvJIWsFjSBWoHJsas6D
wCZxyV8/iiFNWxe6r1SLNQcTFVKZq3vloVWK/EE8INE1mBXJIB4YZX4z4n2GqyUm
OFCOdU2mq3d/cvjyMh//9EyiXoJBGQ7bDS3DtYBqI5EzKWYWmDS1opfYQfy9E7ra
JSAnBw1GGNghinjNLAMHkFHCpZZVb5krhchPT/EPp+Nl7QUF2yinQDbriwvjD794
i94GekvPj6tt3MiM0vExPDT5KEm8iB+VPn7uCJ0VEVYSZO+iXLWPjzjavQ9aP+jO
Xhj2nY3ox8Hi1cg+uBcCSJ0e/9e4dsuTVpwrnGshqcNhN0R0j48p9oltgccih8mR
jQgDuZUdZ/Y8igcXL0xtug/3EbhRefkuLnZnW20ETBOIPMLmzPe3VPuDBXrk+LMe
w1EPa6apRi/eWRenn+oU998dCWI8jZcGJvvGcfrYa8WDaT6jezZ5qaAQYNa4fD3W
gAVk/KXXWnoWryB/rLcdN2Oy8/XTM19nB6m1jek3VEDRFORVTtJiWV1Ts9HfbXzf
zo2tvRQPud5yLBL4KCF/freoXvnIXrZ2M4vVy17NxGexgi2IXtN5b1L5eU4zjH6P
xiCNUQ/34p6cYJv/eSoR3aiEopVxkfN4GaH9bThCIIpSk0sSWGTuLHmOC2RIezpe
1DqbY69LdylPrTLb2Akn0JQJsYbSIdkJlKwX6gy6sZzJYuIRAmr991DyjH4ZHk9N
so/D+JmNNomXDTlVoQs+cAQe2N3snSShA3juLJTbX0P/6RseJ9G59aQ+NY7eYIzw
ctAbrENLAk0tOMTGWUhgVTkVAK+x2lfVy7/iMYRpMJsJPQczWe4lApHZw+Tl6xK/
tewpZj4+BOIJc84AEAXdtKNbwlm5ramBbdvx0CYUAuzxPin5jGqO7fFsZeS5tDSV
Qd+8og2HGDe8y8Az2OFQDsMoXlXj2S8LZi9aFbpoKxSSJtXuGiT9sCvKl9cCms4X
10En8pHkWfJ16bME6wtj78Q/544vYDmYYu6XecgumI0rQ+YHha8JP2KICluEcdRL
MLtyXd3gVGd2BqNkcpzHNSW5Zln///qDZPyghIHrqFOgD4PfYkZknH7WI8qBWjJg
DZQi9UemrQPYHRGZlhjGGfPhQeY0KI70f/A5C+4qG5swDhxcLozsh1ymbQJob1Qf
crvc6c6bhk6xlmQBKA+kMflzQpd3JkzkfBRbn9+kNbheZdpCZ827Sgt+O1DXNvWk
qkLtVZ4KeJSsOiw1Ao1q6DJefMSmE6pIl4oSlUDaRjzxbOWh16mLuz4IjSZRPmmn
xQ0aB8ILptJYSCy+qNJAHHK5SAm2X+tm1Hp+EMExJakVqqn7j0Fc3fLWVidM0KfJ
jFFBwLp+hl8s5ua9vI+P03/ws84ctPmgbA7zjHeH/jTJJ+eMoUozhcLaYGh9W3va
1VHjd8hKgDIpL5ckXtairCS3rdK9bVaaAZWsGsVuhw6WYYYSfwKrGSfb038wzlyO
VYZN+9dXUMm+ODUqkwg9qaIQAXQR+vuCs/bcZ//mnoJQCQGcj43BKHGHJDDeXjcT
2QVW/VbMWxcjZ36cQG2hgvr62CmIvKVaTf8TqZKnVrXRR8DOCxWevUt0z4TJpBqH
VPxpD/RAyMaCG+c6ltrOHC0LK0ehchgMqiywpM/MIP/v6vcLxvCzzyoxVUW5uX4a
RlXtac04DndlUEBOBQd/O8MTuhz3rDlcKpX+/yWd36lKc1Prv8S1G+OFUBD2qpEi
4T03Y3qB+GB/5ivngW1jqZV4q5LscFHyp8oGiZKDpZfYWeya5FZx3k4KFE1Er9tp
O1yEn9UgUvDnLoO7e/IQLrN/UhGVl6ggC0n/ny/sgKit+f/YGnTp89SOtuDZlGXU
PUZTLzurFnCfKCTHNtEIxQOZsptpm0AU2f2aXIBn0gekxeIgL6jn6YPsbmJuUhvG
i6FZiWQZQbznpQGggljaFwVcKK+DIYERMvpYc8zPeb09zTuF/KfpAvpHv7yJLozH
ok6iWrvGGdahFwfbj2BjyOD+/L2aZTTU2RFt5PPbNBK6nJ2p9SgAvC7q5vMoqNYF
edeHCQUfzm3MbLYbJb+eypl3/t+338rXK4k5hK9hKsSrc0DVcu6A4y/HzT2QO7Zi
T7M5QIvCUCpM7cg3M9vExbCX/LgjsDfITjgfPSZW7gVEmnMnHU/7ht6sEfxgu1dS
9nqCXnbnXTO8cIWc6e7QhvM3+A9lLD0FPE7M/rFgZvvcqX+/ytNRdxwu+VkWJKqB
/zA+ppmQilUBU77aBwF47AUy+t98CZ4Cuzmd1uQweRLAI4O0VMdo0Sdm/7g8sz4d
zWtRQKGT4AawXTdXfcIjzW6YW2Tbjt3qFZG7Bw6mEg0mu+aCqaRZeYUsE1XguRml
Q2j4m47tSs3AlSWz/D+9kQeNAS2rzNSn6+sHacygn4UEmzeyhyA2WIZaPf0h7tg0
tEEzUkQGUhOU3dDqVXe2xFWpjueHhVfMO773I64evs1GKtlOtZFzLT6J0UVRP/9P
DFy3gLMbeS3aragSKdqaDrbIORycn11qwWYu0M3BnwXVcpBb69TgNcngOud+E+2h
QaxTG4dlBkLuvy/MTnZX61EreX0GgTDxX86iRAmLAJQd9e/eEsW8U2nbOCry/y6X
yvL6JQcQx5iDS8GZRf/gFS24vrX7zHFeqNU1vyQTDIW6W9O0cZX5ktJBE8yret3l
fnaQJGSn/3VcFTj9+Zh9g3sPNAneTJwhOklx98UXP2TtEJyHg+62TZKFEq3vFZmI
cW/qyVo2KE5DMD90vSB2YcgRWRH/mciILsXnp8ExyNiP5E4IAtUusMx5S+c6Znup
ycDgO4fy6rorelS8uRGnLxsB+JR4W9gIzBjnctuf5v77dG4AmUNytx8zUcU3S6wY
PAiICzmHSSTMNtpFCrWup4Yya4spyeMkJXm2kNP2Nk+c27mypVnJ4tM2ZeoMGTwv
qHNR5HzCc66z/zLsULN0PmQ3iXQehy6mZMqarG752mwJhKHVsqIv1uoWCULzW+2Q
RuREPXYB5n2v+/EDdkDqUgfyN6+BHh+/qkOWTLpQF462o9kqzFIqauBM2qgdcrsh
FTyOfVkgLgZyAC1LksjaWY5K2fa6R4UPBhDwEEmeIuEUj/M4ofYeJmQ6yXCJOsMh
6mcUgzoaX+VhCAP9zxmw4mNepte8JcFGJ6xsgunrSW5BmCPOEfpcLgVoEQbGIG/S
4hMM5EsvbV6cyxrcc1KhKPtGqcHFFe+XB0iMdrYTcrbHPqvojMtQHj/FlJ5g+sWc
nbPswsTVpL3n5LCI64a9PzPRKMewsK31bbjFk4oTPk8fTEWfEviEEtuBEZ8xuO1b
7TgSNpEfkURvQpYd1LAhHXpZcAvEqKcylprgCZrkX1ys2mmI0AgD8Mxe6aFIovNr
zX4VryQGxKkI8haoAyPDxVeBmGm9+REgetO9R73/HQZatcWZqbOmB1RPa9SqlFL+
5rky3UTfq0l/tbGVxRNorIyxms1hImQEcoHUC+BObwTGxPAbTemPcSHF1pBhgDW/
v5IPLg6pwC85K35DkwWT0bmjXOfBqj8PlcT+chw0/xfVZqoz50v37xoA6o0mNr/x
cYDfVilwxL6ZA2gp2z0L/uQauFliq81TYMDTWmPFsiHCwGHdcJJiwg5hctf3u7oO
AFO6P/rAYqss2W/RePcJlr2nWZ9PhXy8WTLzAFXb+DBYyXmdYCNUcQNrHFRIpcv7
H5tD7hiegzQWtYvH2OXJGGfkgswSVfvAD+JFk9MUl3pcoTWuNro9k5Cprd+CJ2/r
JRnkga/yJE6ZZAQYVYHh53yDogks++WzccJaLtTadd4Mp9Pdcfg3XFQhmTupuNWd
Kj9DstFhFwB6sr29h3hnG7JRr7BdkE4Gl9wzfBnq9WfHGwZQKKYNsVijdAM+2osJ
6xnWffMWOElDoNeziy0zNySh52EbnLMw79GwvQ8bJmm/E7wO1xrzcTkM6bw2ZWbO
bWnntsOsGNaIFdRZZUJrquUp4ybvR7DLEwL0NTs3DHE9jeA4xlqVMM6wWmfhK3Tf
yA+b6IKTjdqP7bArCuKOiWYxkNqPEYqyefzev8pFYBOq4STHCTqJLrJcqc+gUnMe
WPlp39CBOGAIyJ1bWlxB5yIO9tAPCab8tpyxZ9E36qf58od6wSyV+mUJMjpCxAhP
hDNdk8A/ThbEhpt6Ydv3WdXcJzQwZfc3MypChKROSEpWLJErTVK9dp+YbgVO05vB
XUfomdd01ecxkjoCzqTVHRTu5tgjcbrQ04HTWql/LRvE8H68tQy7odGPTRTUbPy5
S6zH1h+z9VjNw3wUyJ4VCp7jdBQYL/Iqml7SNgVEU0OfJd9muaxp0yMH9JRhg/K9
wCdae2Ab5hUXeYB5Je8ptZLwiDh0RDIdWrp6WO3Bfj0EQIYsyA4PFK0q8qZG5YSQ
gmlj7vf7RyCwcfBO6a+YPvP9Puzoiz5oUHk/PkkDAAvutQ93L+Oun9kX5W/XHgQJ
iG7HY5Q1sKpQjRB/qmp5jVqBVFv7iB7Uih/9haRYKLrpDMzZAIFxEjW1kuBB06Zq
pSEg74YJGGJQ8HHgyMzOOs1pN0LREkz11u1bgIfOe7DPZsEOHD17A2xTjEbMWTnW
O9XJvHDx+kOCd5UZI6wlPqZR7Nk8Zo6dXNPtzUHASKxQayni9JXOaQ9KiRcMliYQ
Y4QbqR66e/qbsvtDsaRbtF0JtcnJtZMLTjBojnzNA0+q2jEjR/6eMbEPOTjNxfzO
LU+Ticnop7hmfxzsy10+GkfSe17HQSZ+TI/nP41bvJCXXVKK1S73UhkMxverNt4/
WE7pJ2a3CPmY7JD7apkHsX44PpkKqnmjjIq/AqqCvUq+8vsj98Kgqtg1YAxRC4/A
hqsza3SMhjgJPzPf7uCHWVo2oXScdWp7MMT6uVA0EAmj4HmNl76zt5tFWuBqFXKt
wRklJFRgwJ/41IGHQHzhj1U9iWQ6Y2c/IvNVW1YOOss8/Xcpyse3hR50lbTLQjBV
eVT6imp6dzg/Ywq4z7ZHX6i9lDJ6jR1okS8vSnTpMIA+yeacSoZP+etz4jht4Rxz
vwTWJr3fzjKi9QJoN+VtlQ1wDCxE2rYsl/cmCRw0Km3oFrVAoUlZ5UYJJkEhHo+W
49z4Tq85/d0mxOvrdkBdNa//O75dUIvX2oJ5YE+dX7BXYisVyBV8q2hEylZXiruu
/BkG5dkQlRM32Xpot4fIyFGZqb0UjtDVEJj1y2667rlfuzhAYi3sVkycKaIRnodP
lCnVgfwaOKWV6GONukSbfMwZv0vT7osDpU5nRGDEANN1S5wYgTCCeXr1wgj6c5oX
NvlRO0KfGC6B1P+Yt6+TKFgJGi2Bm5z1/CqEwBC3jRLY2Hs2TxzdAw6sqn3s6ppY
5IPEAvUeeWgw1zuSiv3ZScFB8MNdOSnrA6rBDRPpLPDtTbW5bHBmwAoDoULVYUxV
QpTeaSE30NOxzBwZI9x9iXbNzdsXjbFIs52hu2ad9N1kXwxmLhUYBCzwvuIErO66
FsZylINU5sFTd01wTMN66/eyZUQDrn72QZM7/85g/FNl4tsMeUYvqieLlgWmYogC
gHGNwnAwdE3QbZ80qmI2b+o2DV2/8sTIWiVEoX28eUDAzHFjbK9LwhfCIojuMytm
h/Y5a+9ROr/b0vX+rNVn4dsF3JPr2n5lQ3wexKWarPdlHlYqcmMR5N7zMiOwH1Hl
yZmhq7gkzGVUFI9tZ9Wgt+Dm3dx60s9kdn2oCdyV7v8Cz7uGQ5KQNJ8nKUSTn7mj
4uxj4aWGkACZVKIK7XFgIP/6o9OUlXYUzvaC8o3SouxaSBbrdAY/+HmrTx/PuNui
l5IyfnVK+r9GSbrm7/ZVRfvHadbaQ8FpmyjPLMx+RUqrtujcjgDDYLmrEdt3kDb0
i7cfJmMAB4T84lbqyvauGD2D0dcPYbVkmynvevy78Ghs6UtmIC3dUOkaDPxOZVaa
M3HFiKSRoXJgsTwnmwcJgH4GTadlmkrmnfPwGOsXr2UVqjew19sleG3TGXaD0COp
+Yq4te9w3yXq/wbNEX3tqz7mGtKvP7OvIZ5+py1tdSQMwzukrHhokErzWwzVLsnj
Ggyki2Xiif3JokgwoDWPa7jLoyaZcz1QzLUVg078wqoEpGohgug6PR9sgH3sWvDQ
zUBJz8Wzc9Au7JQO8iJaW1MFC+s5GCSMUhtDqTYMGDB6f1QxN+CQYWP9XyP7pDvQ
iOzXcvsdat0vraAvWw/zZDcyBdnMPaVwHy/hS1hk692QSVrDAumIc/jZQuhFjp9S
DLV+J7AaqknbAYJdBBxicuGE+ltjzKMwfdUxn+wjyzhIkPTypHk07Uv7J3mWXM83
s/1kY/22c2CHdG5+ZpnmyggYDm0g6scijap0N5Lerc1DwubVmohxL1oi02bc8Jmn
SNfFWTQ+8JPEBt3R8POPm5/BdOtrkDFd16JAPpjMdO/SWUB29RDs5kVAkZc528g2
3wl/AmPkBFKh/7xZV2/8Q1wqHNlKEFloxThrT75YuXZ9ejfkTzsgXXYvTPryOLGs
dy/QCStnkaiUFSPEEFvsmJKplXaYqSy58aNPVxP+7dgeb61O3GhCmYwaC1EtOnVI
JvqHlCZ/MhApdYroEWqKJsPiIVPL3lN2NTCQmrwT/1/0rxuiG4NIGtDSsuhG0U3F
2/LOLPpnqP2O0a1ST2y1FkZslfRVrsy81c7jxsDNEExfXBmo+kd1JABOLwEG7sn9
P4r5wMpsBNxxBTp5IwsGvGvZUhQ1+4xdUpIK1rpYC4VheD9bAyQP0sk8VrhY1ewb
TqUOMQTRvNbutEtkK6N/jhN1kLzTD5Zbn4D6s4mLJwjJCjmN/vxZSu44aqwzXNYR
UPTzWDsBFNS5T+habtEP5O8Ewkm6Fvi/Ro2/fnNJJT3R7KEjKetxG+reyXGqrFGy
LuRB6KrbVmSJ8d+Nzq23yKOpWm0andRs6CHI521Ft4O9FN/rJfU9ZV8dHZegl5vC
OD+JZR+kWzMEVL+Xox7sqcf0jk+1Q920uwAGjIWr6artxTjmOC8yJI/l5odReG2r
0J+jzqEOGN3ovtjLTP1E5ywjqh1diJkS6ujHR+I358Mcm3Wpq71ZBdkczsSHt4PH
nB0baWxBIFa5Oq9uRsfdRY/E/QufekGM7SPRYOx/2bGQN4ORoukPD9HeuCT/PxkH
Jdo0W6QWJEVwsp/zRR2hy6wDS2WpsK0299OkaYOWqI+W/5m9G6Qt7CYW0BzO9c+v
t2fL/yN7OAUkJiN506EIxEvssQ23YYdI5hAH54NgBxrPasQXc9BZWNHCyfx3w85s
owl4EB0HbdZMTZeU16i41w20H/dLedNrFLvd/zBD3Lu2Ap1NqNmgZ64ka1cGnEd1
Kobf8tJ57+PIoY7gs1Y74y66Y8wk+Bs2VEWCnm4nWiyLhSb2GAGbaR1zVkVTOG5C
yuhqstxa6MTkF0Fa60tx4/uiZoHsgZrUYVG7aav6o3HNQavMDna37Vkjbe/Ae6r5
FcUikBSgCf1QThm501zfiHc3rBCHEje8j3D1/odNXJZ9NFyDQkPCBiSwqrgXoJ/v
GhqjaxWmTsUb0vfqFfsA/3lLh09SKEPAqccVAUMIoPi4R82hrrAYZ3ZBvHZAdtwf
JxqilLu53YGPZqo5RMpWBh7Ue8oJT4F3o7yJX9ujVHFvbnfV02A+d7uOIwn7F3gB
batAj8W4yk2UUUnZtsuLpnWM+DZfXVMiAPyew+ovsNl15edlR9k0EnWLJKPdhQyK
q1NalByfZwWKU9ZMplhCehzeEOsU3pimdMCbGjPcEQB3W4qR1bVDUhIX0bfFwAbp
mfBokULeesQ6fUAb3FfGVc/voznRpUxSNdEwsYttVppFAmIpvSx42B+ZkeIfDFdb
79mAWd38SHishP232XLu6Mk80dIRHrc9DoMT8Id/LFZzZje/IckZivLdXTXX0siz
pxwHP1bOj35pYWbl14M5luyshC0FyFYClV5zerXWzg+mPeS8t4NOJUJn7ciHcaUd
NC8LisvtRtf1+FKr3u5Mo8qjkAS9RkLup+ufQ6CIRETfcu1fIEkWIeRB5BUusyTM
o1QH9n2XVTuu61Tph+n90HHp2NAlGZSkK38T6FuodEAzVNql+Ln6OXmdHLu8g7vP
P7ijDyrXXf4NlgEVMtVEw7EKi2Qa719e4idGF5MercBYNpCq9RapDQOWJf/4URU+
+laEmK9dp8o8L3FlmnGlRW+E1J6f9Tp1avYgKSt42io9BwttcJkPHZRPBuXk/huV
mX6Rvh9Zoxs1yHYhjDET6xz8KDHl3HQPHQrV8gVYRh/GQoLqxGBHMFqU+76j/Lu9
YqwB2BhsbkOl6lIHlwu6IcS3lwDUkf97KozqBJZ+16dsqcL3PvtvNWiIi/bvnp/V
DbOTkXT8GAMAUS3t9YM7qi7lJLmh4fqu0DGb0zIqDlQ9rVP3iC/rWX4jWcaovTX2
ABTpz0fGJO/LT9kxDY0YciCeajXYtwUms1A4BZKnx/m3Hhl1+fwLNMfXyI/DiKX6
7CklyyoNbv8iv9JCncdKx3gFSyK4J3Xdz13bHXsy8gBs8sCzJYsKogldFbZw5tBP
4YDSaJVvEhiIxmFc14tR59r5dU4IHaEEC+tQgyFjzfOj5b/UDicrGIkDgVrBb78H
AzMBk0K1S8Z7pkFK8oyVQzz76StucAZRyjSB9V1vUfwR9S1Wbjs7WjYABPVbM3mi
FE0xjIjlNMmQ2LoUg5UjObLIEUt8/3PyW7KV1uowMugqUcSnd9dswRaLNzeAYZu/
vIOICuuJy+b2B3DwN3skSFsL87qAiJ4hCtabJYQTVANRhUX29Uk8rT/+cOn8YcLO
IhfrTBp4/S/yY0dAxTw6sEzMRz3iFi2EBgjT9QjjGGATW7Skq7zqeb0S1Fdqhvgg
MAC8IpE2rgg+ZG2M6oQa2c6pu5aj9hQ3NSKBGHulimKA2YhMaT9bOaQjwsRlVKeW
NHcxXKZ5IhaivKYkDwRoqKXP85O8EC4TwF13h5b8iXCzucb84W4uw0s3JoO45py3
CUPGkmr1HKQeMhtL/BSF0IVFMDcIfRvYwuTbqPZlHb6rjJo0SLqhjC51SsvUd/k5
sisvjNGnlfc3MY7X1gfC8ev+AnESW9S/s1Y+G0vJllw6xaKbBUMYLDAn5UyWdwgs
35At406ybRxE+xwVZAD59pELMlNugWyjJbimDdh0p7wdw49hbsqJgs2EX5Wu2A5c
aw3oaGd6ADhJdMApv0wG0OVRHZfglL2UotE/PkZ6LZS9ysoQxo5jZEnLU1P7qHwJ
G8pKjZDDSab/HCU58J1zc+RvMT4na00fxh78yg7oVkfmyneMtxdWEoszNrXubQsa
tCtwpKeFnMyfT9RQUUH4tHlXY+OLs+k3vzo488WJFSdvpAmtSJIVoFYms9GHstfL
EGAbwTfrR+KGmlPZsBFeBB44LSqPux60Dm9LWPGEKiFmSk033BbeHu9Fo4zU8atm
JikmXI+EpPEV8zg0/PsH98y22fNj69EYEYLTrP/VWl4sSNjDI/KaOfn6Zrr12zBv
UxsoMlJinZG4fmpcBMKYc3sq+aG8KBkVQx9AZAcyPEjfi5NxPyMPwKP8ObtsBkG8
K5WeKit/WRDyl40ACrsbR/BuKg+p6IResTIS6Jj5Jl20smVJXdeZb/z1Kr3YvzQ2
egBPR6kIXBtoYnGX7hBvr3Co0ee7f11L5yqsRP4hJ02IMajrh6zJgDEQ2ttNNj04
EVGPbxQxxMKhyil5uXhBu9VRl6a8SXYO0lBYCDQuoVshRlLwS6yQ4B9XgNMGa/AL
dx9Lzq5pxPDkqPdqX0XbYHXRieEzy47MpPT4h/uyJOm2K4ATSA7k7QsWE0mCzM5/
gSpIS+R/HqI1ECf/mbSZWAG6Bi2Gshguy2mR3Nkea6WGdTvikqFsHl1FolNyAxR7
bQTF+plU2XYLwEfJkdkbArJiz424CPv0qvQVo0zDIgFt1mhkfA+Hje6LdMIwMRl0
k63K4aLnlypQ4RWsoZ+IKNkxusKLuSUgpzUUIxjgAjDhRnO/hqVS2ztwAX8VEYZI
0rVN9VtvhE2VKjsMuUfIMMD26XlrYn14WEX5zhPODfx/lC88mgw80Vgi1Bjf/HFR
gyO45jMWrSAK48caKhcOw7buGjRkr7Huq5Betp2xLeUZ/t7sdWuP0iw8N7vVkL2m
o3ovys6Mo3+p4JN4cFbCa4DI/NvKcc0jPZJpxsbd7mUEMVOk/ASJl1TPO/CXmPSe
TorrytmmIrU+Dft/5B9Gr3mlw1xHSIkkJ0zt4d4cjO40V0qibfIUpPncrjF/WeWu
DLPk4gD133DqFnQOYpfCHie2Jl7pSduh5Rdn3NMm5gBlf9RVqx7ocr9xKrnplsco
IgzSpwJfoDzm0dIRrBbME/ElW/nQ9F/31Rhz7EglRSJ79jtvPg1lzOff8cMGMQ0M
MlqlTX++YMyaIwnmZRi0b33edbwfrn4QwyWOfcWrEUy13EiQ0HBRtXFqqG5I5b/j
+P0L5w8r6Z87GMrKQuLt44kfrMU3nIMdTzUr/mMoz4+8IUp166WmHgq0ltFI6lwe
tB3vtFUaVae8pOpchN9bRbUw0JnK+ZCwj+9chUiB0lXF8f0NyrqxjxcvPrPjks6f
1zKrceP+0ESwtFbIIze/WAlrtc1dgVw6bIDCtNMR/CfHgXU1K28WANRSdIYs7mSi
15teLB++qEr8ICCxTtFc8O8eMjARFKJ23q6UXRs59UlufVGBGXg7yS/8+e8ir6Lk
uPkL6xLm76Xshn60hw9vakeR0oYXVqLItc6kg+/dCL0G3joK6ge6JuSto/wKSAKF
p/4+mEsfgVkrSBx3T+YJGgIP0NgNar3F8OI7LFosfsY4IgspQdRtzw+H3i0D3f02
ct89rR3f/FU4SDVD6o4rDx3yaWEKIpNiJAphIw8Gpgu6lMcQne6Lvbh8AkD+CA4z
va4xXTYcqmJxI1gCaRUab5mSz+oColkg5Ifk1MJGf8u2CKlhzAnMZASAQin9ALsu
aVx2e4q0H2jgECp5Bs1kaoS4EFJKW892mibDNlXbF0rReLpuoWGqC/vb67Lgm3dF
g+djHHZ+ZP4pkMyG/JSwJ26rrrQOZfqZ5rmaPWkAfpYcZ0L0qt0V5qDJ2Mu0RPRo
bh1juhIN9Z6VwZ4KgwadUSHdR5McUcWkNyD/6sIEHehNp64Hm5E09sadJJdqJmnz
1FHLEDMBeY5Kg4FJLoh5l3cjLQ+4ImHtW++d6SLFjU0kxxFQsGe7PPnC9U2cH9cW
YirNrscjUHo3ngFX3/7g0Xx5arZMGBKY49e75IRVRN/IoFQsXKmlsSkmtscaCtwr
I2ee8AbqNat3uyhq+U79ybbolxUyD1cpkcAzodK00BDWvShkUJsGNjCI7F8p2A/P
zIaY4lPvVSfD661WS/SZQ2/2b4C7Ah3N7nqRY3fM6YZfpuH0p5+SgHqpKmRETRJq
9nT6oxw37eNkQAP6hdHh5RfhDGnRZBQ7aQyzgqW8NpDL8stgqy0aM0YIUZVx5Ay5
QU3ZlJufhZXSLYhVqgXBBDvn/MVeAuNfRwb6eN9PADylkgVqsm9wwitxmqr/oyvJ
1yvAnLi+uX624tZBgt5gXYQRdeBphAC1YYbjQOMMHGdTDN38B2R8/nANqjC2rTRi
MQvicPHMw2u/WiNozsbkjyEhiamU/IUw2IfeuL1yQw7zXNg5LrjGCaK9H+0W528+
YX96eU8NLXLr9dBkc+jkT/+yArT56cr2S3b93eO9PJpg9HkjJtj2EAGOShMwafup
oZKfFeeDbYkqoYk41pr69H8uKZA1woZFetigl9gpR+lph38EaASahv2EcWExvuPj
zWba0yIikNZGrW4ELDlT1cChGY4Zi7so1p7IQJ0VjJJmvocoDkyzPnXIFk34OLRt
aNcHxLoO+5FOFF35mbt17wNRrtdyvdO4U7ENaTiG2Mictwth2b+vstYaiOZIHGTr
wG4iNThCLyygw13EDPv+MtEiJzqKeIZTiBS9Ex4jKApdrqK8hQQBjAuXp0EPJmFn
zoC3yp5B7ky7bqTnF89GiuUc+5IPVMZKairICAaLF1E6jN8vO3s/hub7Tt0EmPI2
TBsrHSydP48SHblTYtztpq+e4ZQ3iST42/1ReihiuL50QUHeOFOA3Ft1QUTtqI0i
bP6Fwp+maM5bI7dBYM5YXVkbkYMsfhF42sgKKoegjhAAvOSQlwWReoyCgz9Q+aAm
Nie/oN3s3/fSXgwhVW0iMCFekccnZtaz987ve7A5eFb0eNfDAX/jovOb2fUAD15V
6AYrgvPvQT998erZonFdteXFTKdD58a2CSB8YTzYNCAYXTWSTeYxqdrrkeY52JN+
G1ShRM0JVjLh3s580S9mSCan1GaQNwog9GGvyI79JgZfI8W9IjPtUYOgGLDSiNDp
s6WJ/HoWkSC4wXN7sy6QRFcdO1sUigF+F8+e35eRKHRX4J1xg2idcrDocszna4ow
cJ7zwiBrnOIXvw1HOIItgl1CFKRRQyU+u6jXgwfk+IKaRoxCh1Froxu4nttwr46f
kM+kOmo3UN8yDaOvU2mQQsIQJ/3z8xDDxHiTIA28ifvEY5PnJgdP8jexC/iCV+q0
h0m5XURk65PlMVw99oxf/Q5+eiSRtp2KMP6rs4JogWAIOJO2E73+ahgZOoQytFj7
/0i6Ewt1PnhViz0Gcbg6lqUSWkuB9k/iTv9juZsJvD08SZPKZ5wycnxsgcBJqsFh
Glk96uRqEZvKqO0E3c7mBXqSUfKmbkQGmm82U6DEF/6RPZ0WxqkeYojR+5AXlb5p
5oqGau3+u3nbDK0tayROqRRTmJ5JqVIznax3uniD4lZ1qqv1SAlj27KlJfzQ6Isn
HRcCCqwFo+bnLZwnPGxki1RRI42jZ22SqlgzwrcZWxKxvLial8NlFLC6z/Nb4OqL
QT/D6fUgJp8IXEnL0rza7j4hihSW1SmPAdY+34J2wOeYESBhwYaAmE1c6tLWh2Z+
0cL3FQQx/C7xvWqHe5ejWUoFLY4VCRhGLEtFWrTWDt8G+rL/tQkQb3+1bhE+epgU
6PyH6C9ZCczTQ2dHsMYnZY6WLzD1rWzLvuGX8Dblvbj9mW1udyetARFSm7Yukw0N
hNT65L6m918hJbHHrm03NFBCK6oXVskmaeDNnY9ZN7Grn3hFXIcPEO9StUPFU9s0
CcF0x/nu26SdXnvbheUlGmQUWPGaEJ22Z8gxFwF7PQ2Vr6953AaZW4AR4vm9GmUq
V7Ub3JTuo99fBxb/hYhJJWhvbeWupJMD2j4oT/RUROWW0pQT2Cv2GCkyc3XEN/W9
FTywX3/wx0V4VVEPqD9p2IH7vjCZt58D3UCygg5ai4MEaqasqxeLW5VGHZY6Ro2l
rcXsjokdIsx6jH+QnqiOJZwqE8Jtd/L0DIyGjQydi+cd83TkY31KkREEPtNjtJ0j
jXkmWZQQfHDNLU26C4qPSjDrSaGvRi67GhYPi6cbGKNw3/7PcdOyLv96/ToASr3u
89VVjwyCAsm02yRN9kU7lUu7yYAgmBAdetm/00bc2UCV9qUFdY1WqwPFVuXyEDOg
YLPtN006CMndKRSWAK4zfmSRpWHIWFXVSadsYHlJruGU6LfUt3T+FIfitVHnrsaH
AhAz/aeqebTfgBWlWabiU0ZEIDG5KS7jtEkCEKqnJk43hJT0useqYir7db/oRkZm
juoKnnviZXs6GyH5/LDz28KB6GwbZcRUDxnqunDq2D9uwwuqG+uQwWSh+HmWgWEh
/mKzWLjvWIGAqkTjJeIYIkT8GGarustxV4X2PvB5GMXWZ9HqGxjYXhcDlfyva/mq
9KHeWcp+kQ84GiiC5lYtPhWpzf2Te5/JkS8IWPWAWfWm1WXoBwhpJiPFJU18//m0
YqJrEteRCMvdq3Q718jNHg7NWK8oCmCYPfK6xArE3dlG91f1mHpNYCGec97ctPkr
5fdwR+ehMS7ovqbY2pUxV0XQ3TvbnepzJYIsuA+vEBDbX0x2AxavL0zF78orjFcV
Kkn7zdr78V2rYOL3iSoeSyT1y0vDzAnwLAkWPWwI7dTqEGl1YJx1gzbNpQRSQsnz
wUsq6s7NalpnOZPijIYdaQLkCkRZ1fLQ0agMye6kRFgTCePDMCCpPbEwk5zwHhhn
SVeeNv6B3M08J8hQ9BVCI9vSXVUe3wY3w/6EMK4xA0uF3i4YImutxeawSTDRMX3V
rMVkr9i4FMYVUiPDk81kE7K/2RnfnJdRmPwMyi58yNyPz1z8vlVkAP+LolNqQWpD
TmgnaSS5OU+V8wpJY7FRM4DUSWho/fidGx9LGGHdpQeli1GqwkElt8mpDFE5NPhK
BD+GASX0/d6TrwjVL4n4cMb55Uds5m1zWYS2M3UQS4/lU33k5cxuQWAnnYq3XBGE
FZ54lmKBgcKGY9CC7pdVQcpeVBCxs33dJx4WNbm48wn/FBWC1j/Q5ZXyHmZkfrzk
aqlP5FOup+/+0I+4hBa2xy6sn28D75Uwekku9fnTTkPr+wemrc8aN+K1BgpXRM/r
R86p0XvoUWqXFQOjvLUqKKpGoZAwGsC10VL1Gic50JxtYMPynqoBjvOXQhUuIyiK
rmEg756GF+47FKaof8LIRmXArfoTtC3sFHHOf7J7Wt3Z2huer9Fyuq1F1HBxDaMM
ym5VgLSU5wGAivEWewLCvSvHSHMNWq3tgZUx8YDssbTIA//BleqBVrVUKR1eUXxS
c2yGXI8a9eOPaEahhCNe4JmuAcI6BVPTUQo/OIEwds//TauNueF5OsvQ5c5JiRJA
Orw8yOnWvB8KtrUgYoedTLc6bmuJnUlxl2hd2DoVFzbMvZNn3eGV14jTH5S7iZNe
JXuRSgHD4m2umAJ5EPNBYCOL3g1KDFqC1ewJZRnxRtsCGgf8Mu2b38a1gytnLyxP
mKGThKggje2KEiQOER+m66iZf6OD8J8VD6SNyjAzyW6J/aLfOCjcq+3wTCBkVCWd
p+WZjF9wqg/KwbDPx2eM+dJfi90hdecGzWhQ42aZl0TXrNwowlw7D/iS6XJgAbXL
HJk1orDrHPryVXXCSLcotffdHEXwwmWIv3Odf2T6AGFxmoh0GnpZCWh+K8rI3Hxw
MTW0NY/9YMVxCuK131PVxm4mudrxrTgF49zFkqHO2Bo20HnDMVkLeTUCllP8Qa+3
uVSiMwz584gaSFs6Gd0IFpo4IY5cTO/Q/jcrGF2LvHeffW7GXE95H/CJoLsDZSGP
/vmstNkW/Y8dI8iPeCXho9VJnmoqVeeGBVk5k2YAPNjG+1FOCXC0il1Ga2XjcbQ6
IdLtN4rTbm0HdJI3TtMldxYuVAVnkTDJmCnb7UEdDlkY90wjKrVMjgBTeIXZShlS
wB45J5lGNxi0kaQdbaBbIHHJzx8YSjmj1xKMebLqbSzESBcCcp9jzxhZlsTKN2yg
ZBHpLuYnDBusCvcE9kWfcAtBSp0G0tdExN9qlg1cv9iRAQUhZ2mCoIqMsaAIPpQl
tWVhxiF2jglQXa9XlZMTPtd9Nm3REsElMXBVis78ay/j08EuncmZKEg64adlCxHj
DW/Z6fW/Iobr72dYM51jMzJiKfjs6Dqv31z5efH/1NdjKu48zO397doCB2/8Il1o
ipbKxY8kaZkJWQ0zlp+AB6ga5yzjPU6plTCZ1VFjm0uvOQDboaw4VVQTXf9naF/L
9Yk+GsxnahvecvoACkIKxZnkWYk7OWuGZvPSj50uGM6H6i8nt18LZ59Amfs/MwtM
JzJdkFm58qxXqyz12BtcU4+vA/YGeOwGEItVp1fP/9DWBBVdoRAiD2bTYZGwDHw0
v2vok+DaBXu7fGo7F5w5ptdvBwY8IF4bbk+JGc82I/qjllXz6wbNHlkM9OIMexsn
6DLDmx5ENZKh5qSF8zUkXNmvBJpay1usqv6BeB0WRY4qNPPxC76BfqtTKorR23Fe
LTVeegXITQrvmsc9WWwn7As4J+zWnEdr/3CGqI2pfeTSRzDhYztuMyBxKKOKrL06
T26DBNxAhZePNmOP/4UEiXxNqsxrHP0iiDkhLmIIYIue6qBUYqNBl6R+52MtLo3o
ebRbsaz2XfMNDhqjKkWVB3Jt0xFRD/XdGTm79LtySB7k/75YLyzwqPddi9GTZNp8
efNuM80ReXEg7iePlJzaPcF0Og83QyjXHHfAXuBYOBEyvDJWqKFS6ynaXOkgQKFZ
v5VnPwZ5wrJ7ZpNiiVdyyXv6l4SJVXL59xa7yZDZN+wnYJz2YpOmflnWa89QY/TX
7JSyd6HmA/ov+D77y4PTOI+F9xq+aa7VN4D/XBRskdXzhbguyvh/sppD+jMn0Ikx
BP9rtVvDCmMcZjL7BJBieME4fTYJynfzmDS/ZEGdClEXoRnjQkyPXMCdcnbBcKDf
om40bosCaPNSLm+5CR3GlTKHoqau8jpxI102KCi/URb6tzoXlByAjgEkZhqvu9sE
IaBaUFzRspegAxSZoBFxy2YLAffS+wK/Qm8kzomv+my5pGeNik4mWiLUpABqfBpq
48fSPJp+v+tCPEiMdv6vnFai/SJ+We4La/OxhFZ557gS2GCZj5rk4uhMGJKvV/yH
GpuGgkU3j7P0dyIiChStzaPOT9bCcdR5dl51UecPUElR5yjzUmF/JKYGZR23EEDq
yjojdF/NH/qjJY57cmEmds+nr5T0N9THuVZX4XN5gZ+FuT28tHAzBcTU+kFsgBRz
N/7TGsPEbAhJc1OiULPDVdBTbhalDD6M9te0jXu3qOfOUAIWLTfHsmpY+bo28HTK
NoogFQDXpSQqJ6TzLFaNvfOrDg7kUMuGijZnKOT78TLSLrAvWH/CTZcCiOaGL3vM
McPuojKCNS5fJmERdP0xQQORuuHglPlYdHMmQ9Str8LSP2ErDZ6zl3C7GDcVcfS0
wJ6C7f4hcffdYHFJ8iVxjbAHhP2/Z+iQ+g9PX/8QgcmJ5ELd0PYuHdTKdcgoFUJF
ODkfE5vborrZZfUyRj/YQG/L7twDh9l4VIXHiD1cJ5HPnzyU4zmWiO07JOMkZLmm
d+wGod/hC6U/jsArBCb2XnPDrt6BaUmi9JW/8nEj44xbT0wF5aaLvLCpXXEFWwuC
TUJ08y5ZcRuRPRBxr/OapmvdXnY0ATSxMxYZ7UXD/Q+XYBH5bi++HYlH8iuyN0CL
6+d02y0jbdLPagK1xPRmx+6cBWgO9b6/5EoeqFtX23DQ+kbHPM4rbDvWV37m8Dm6
/9vOd7ZVBvhUoRtWMuJ8ul9/YdH5xYy9MzbIRTRXN2p2Z+InStF9E5akbnMgauzg
14hEfLTSQ4EoUCDPnAPVH5hfMQiFW0GUAB5zJKBIBhciqVl5+Ki+B5Mplta2vQHD
Ydenza+sTqG9sAkzIRpXayFynnt5pDAWCJqHufNr7oqNNQ09BkQeqEHr4BkWil8S
FOGdLLA6w+RmDIJi9/MwI/985izbxPnhVYRsW+pn5mxcdHHDJOyuKDqP3PleufbR
R8IlJGXQBRS8j8cKs2+Rt8xxxKMuZEjfrW27hsx5tsHjbebNRabUE8E6Wm2jHkGm
woBcA2PH3jujq7mO10AUjPfz9/pobQDfRcD57d3Rbys0KVSJ3FLPkQPXIB0J2Atv
`pragma protect end_protected
