// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gweVPExFcdwuFEL+/LW3JHQNm+M6xuuAEuHsbHXQa9LaTAe5/FpjG/xfYCd4j4/1
hwfqfhl1o+g0Mjtw74JErLUoWeEMrS6wCJpISxRMz/H8MLJn06OIBzURG4jVhJ95
J24bX3PEcBAIIBOWk5dRUwmuZm60IMQwWSycqM/vWtc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9040)
gszT9iqyXl/FcxL12wV9zegF0/HYBfz4uG3wZ2LkOmt8VoEOjzts/cbDbVfp+b8d
s+9FuU9jSCQ2zTMT6kmB98P/0AzHRhz/qfBioZkh3Ah0WfFxFmK1ENPi+Mk6Cs9w
J0yljhWXyCXWYX8VH1KZE6zx50U6AugPts5E1zsWEohXhbqdHNM/2DYblI/pJ6PY
QDkQvSV98nQrscs6jZc8dsVh1JHwohpr+Ej0Amp0lTwj0qvBS+kDc65I+KyPyk5j
4eB/lPEkVjONq1TkH7ZPaOw1B/W6Ag/0DEC91afxbHyW24jCMZZlBAgTC8W8DAMt
gIt9U3xymNXPAgAg4wHnC21gXpTbnMZA+tWbBzIzLkUqKwB3W4X+VTmTs1e+Nd7+
6hOlFs8+1hhXkCtt9wlbfnpKJB8mstj1bpejulG0oGXw3tuVt51nvjD4BbERfCcN
DyV/6sFi2wXT3mrwQOOmBoNXMzTAhrUj49BsBbeU3oLHu5xxBnXYzvjZkk9VQaVD
6Sow2KDagbZOKe1+HL66aHDcP3NcIGFIAaiCB7qQjA3F2CStURO+plt9eATN3ZxW
IaUQB246mfWN39nJFTA6J2YSFhSZf/2bZRQ5lByMd2bO5R2BAVQSPLHl2jp9p1Bl
xZC9FfM7G9A1UTvIUPvfoK3ewHsrSLGsqneC47SpU+0yHofPZjs4/6pZ4q1CErNo
b9hv2moea6K0sV8NAIsg0cNALSqB2SupAa355D0fYsYUTDNOp21AUqjiUoO+BZq1
SMCyrbH9fLm9q7AJ/jxvMAiJuyf1Z0Y4tyraE37fUzfiC/5ApApNkvbb+be5aIyu
2XeTqk0Qg+4v9g+jxoEIW+vG2PfjLAzAb3jveRtJ4NNOvILk1rT92xUEAeEwGnuF
j7xYIeZIll7MTzj2G1kvom0RZjX8sCDGe5yiiu5Ep+rGx+KZ20e36i2bEnatVrD+
FLqh7t0qLTuNcDQ2jlRoASlpHVt1wxxkuG444NOAV9CoRsTwJKcfSvwGh+pDA5CD
4wuGqVERpZEPMFHjDCnM0SmzNmCIaP7CNlJ9zdYhxIUq6GvH/w0yPCOOxUYozgam
DVw+UpRxszD4+xL6FPsxqdnDJs+kO2Utcvhtg594cZOGa4GuKCLts15plWCCL8QA
+VI+gnpm9dfeYeiJglSm+2LxfUEVdecBMonrJBrQJUiK61blTALHoYdeA68kzkkJ
Bh/g3VZKztTiSU4VlbA10rlabWcNENUhgf4uq7zsuB5IVgzL4re01qI1dsVoa52c
MNqC4aHNXrnRbEALs72PyaXTO7dtHGmdQ+nJuiKfY/sO442dsa4WaWLWrsG3oz4E
0LAkR2tGIm/TEw8Y2d0bF7H+Ba0hI5TeMzyG1462SapxxqDa5XqzasXoA/BueMzK
L/tVNX6lCHbMp/N4/NumvpbBVtOkAYXY98qA2KOv1bTbAMg6buEgCYVltHzS3m4G
EZEgdnHokm3nfMXnbzEY13Vp+MjJZLno3nJ/78qMVCg7iIw6Cmq8obeS2KRUy4AZ
vItY8NEJcw39OdA3zDRm3G9BHqG9ElEL9Cry8BdBDp2RSLuHydunCDreIzqJ7ciV
RpUN7esJeOapxyjhx1CY2kxuVitrszwL4hAjskPHv4WJmcpFP88ckgeWMpqLSaUd
JMS8ySB6dqau3gSDih5FUw+yl9I1QQVD/zBO+13T5LTqojR/uRLtmN4iJA32QFER
dGwFrpAOjv2yIWxhHrq/VVazA9AAutIz7JEXGI58RslACb3SWIAemktc6QHrpsUU
mhmfUMI/wanPoDgsf7KcZ+gpgA/wvaQ8duWA01KB/7Rw9ztsg+Icwe65jIRJJA8b
tzVBjZj9RCC1DoGhHJoyB1rs28J8MwaGU/Jtl23MlElSohY063PufsgxcsrvWvs2
uhjmnz2Yq4ZnMIkfhigxOjA/4jqlK65/+4FdNHrgJq4YBgcC0SSfrFAUAqGaFobm
mm3q7tqL8yb31TlBroC6HzsgXwwNUq8q8RWF+oFxKmcmiwbvK1j/O5U6fS2ueRYz
CzgePl9fWo3p1rQ6Pih+j47XWE59U8skv8CTYTt3xUO5s58M3QfWaXTW+R14ihDC
qjIMNq0SPj5sgOD1TVVuywci+AmurfGMPIAi2tcUoPT+qYWAVM85e3wFr0/P81wF
lCzgKfy4Ls/2p3c4pcZ+LS9FwQW6x++wqg5mCYrT94nKqRdNWtOP8EOzVg6freiD
u4JmWSsehOnJdmu/vrrEDb6i+bOTBLCYutg11oUO0DMgVNmm8XzlQFe+HzZ+wnKK
SWe9djF/4E374dM9fLle1NoevnEj94mvGXna/3leSAk/ar88bWnCMAApW2n2XLDE
fdLtR+XWxC90qmI9BC29ideE3lPxyndM51RqzEcqM02xRDvZZfJXEXgNJDcZZRhh
btdTLyK7n6Pdmwkx2TYC/0YOV/3Zerpenq5Q7U51XAKv4aJLpXKzeRVaIdGdGNGn
Iz8/WYNu/ZI38GeEB1uegz9ilelrxPfOP1j4ZGmqP43l4rb2zoE9n/9G36lbEuTA
6rM64hSlECCg9hABDYnM/+6RlccBw1ATJaHipyqV+C9hFnUGQIA8MZukUi73Yf6j
MmpHv10kxA31ed1ZJB9LjyZ48IGAYLONMAqBENb/Hxtblo+L9vFCM2U4qjySuL4r
kVmuSeWVgCk3FkqyA5diiZSAIUI46sduLqcYlC4IyXXvAFQ5ru9Jeqf1rboIOH3w
uQ1+AqWvgNPSypG9hsGj2ZWKRtfG2vrmGdUIdD/upVaMKO/AZCLrHJI+/Ox5EW9n
3jpfd5LERtIUF9lCqURRqA+b0gh6/GG6hjEpL92pYTKbFwW9fRwny12YbiWIOLpI
/ICeBkb4MtmzgAgYTXoTidVC3wZe1Q2jMOpC2qFBMeZ6PRUSc4c91XaASPb4VMwF
f0SQDzIdLuMHO8BwQPriKuisNH/U5KlZyBeE68k3KaUNfQUKK7QWoQ2T3Bc13Gun
Q1ZcueThlyEc1vFy4tpxkaUJLrW9VIvHQcx5Ak/hOmTZStC6N+MW1Pvfy788sJ2A
EqcgfLhT2Q2YFg/wq3lwjhDigM7JJMk+1cEFi1/+7Pb7ibzzLsNJEmueRvFGVzk8
Abcve4xgExKIyHWzR0znBo3BqHThDLjt9rsG6ydOapwzTSuIvdAM8O3sRLJ6Wd5S
XY6FLR2Hiy2xZ5bJ2PjO5s6TupQ8VlWnVYBtZmZgRJTjdV+5oM678gWrtOY4XUCh
so0q9HkoElyeq2OWsRM5I2U5UEMR0e93LhJvD5eTium1lawZ9Xwnmw+oO4qTBVp9
wDQqgPGF9sY83gziZbX1uSm8WMqnT9aC83AdrBKYArm9NULXj+ft9RESSt7b4yJ6
dPrLwwR5rc6Jrr4cS5m0N6LwTbnkqfZeE0CdYYLp8FJVsT4dseebtz1rcL26jRmr
ukB5N8ee+986DkRQY4UJ35WYGepK+5UbCHzhoIckT+LqwnT9m9kP5/Nwowd6XMTl
e9Mzje7wf2gVtz9sHgvwJEx5MXN37WQ98sQvMnrA6qi0VS1oHL/z9gmlJlm8bm0K
bKYvpvuqd5d4A9rn1hByzDUZ/hSudFghPWdCCgzvKFyT9XBXZ2/COIuOWJ+lM3tG
gR0hfZO/7P/WySfX3x/dJfh07TlUEJX56AjTPdnYslPFPBrN2IPaT7qUk5r48HL9
lt+B34wa/R/b73Jt0jaG08+b4o4GH7Uf0FHYV1l7ybNhvdw5n8Fqc6YF8m/scK9t
2LybcWjUelS7tBUmYqhRmZscKWcY+iDvwRLE67zUnhCyMSaIHxvW9lv0LXimMbUZ
7GLfcS7/cOAlHDvohqTo9/FzfM98VD6wottKivC2X+D5KmpXGYLXsvi3pgtI1RaH
P1/XEup6WdNBLQIMo+d2Oy0G9WtUr52QuTmDXN0Om8PwhMyDwY6eZL0277nAYo7F
RpcuXDqbKTXOXuqx4q/dTLCSdoMkqqBjBYbx2v2Asc7TY6n/7XsI2Co4a1e35NKn
bzxFHpa37r0I9/UKfx9vuR699urEa8OxR4ywocRcJnw0jeiqOInLxmntdSMQWOyu
jriO8yGIcLaC9yKkg/xzi6rC8LO575Pvhu67G4J7idtXI6imdBRaGlmzQRDyj8mn
XSKi7RguBbhsoJ8lzfE8SlJKrLem6zDgz4vPSPn1c0o+76lykXDdenUsKnQwE5u4
Io0yasXsv71zEvNJvInbXBqnccHIb46yqwN2/C0y2M5jJ7/xCx0CL0YNeyG/CJmI
5qBUFj7NBJEH9luBzaNf/YUR4sWkDmd57QJahlDwM1tLQVEqPSpRJrwZqkq3Lr03
ubZwJe9wbhXGaKhYKFMzCggok6e81sxRV+49govmnHYNzMFltKkBfgQ0rGsfKdO7
xa7Ky1ZMCvMU6GCTfSumjE3rO0DZg3YQFT5++VxmM3j2VH027OgrrWLT+jvORORp
ezI6nl7kRsMGqbOaFQnlD3NUmHHwEnnr2Ryf8F3bjkI46hPVjUxo2aFaGaiyBEyf
Fp0yAwSHlIZSa2uDHQQzKelTSdyoiONuKXM62o8sKp+O9Rqp/UhhfYMuWEu+bTKD
fZJL0xvAsbDDUTysN1P2RAGd7kCxFuHavskuR2oJWmTv0WOYemr2xa1EGU4LJQ2E
jeqPFuAlc2ulRBleSTQ2TXS3SdBbLIejKG9TxrCDHifNFW6qetYBXhzpyjXPscNd
sK7AB2JoWcXqMNlXjqLu/x70r+tx7gJnzPtAGVKqkx3vlOtEUzv1wB0PkkQVEcBo
haX5ev1M85a+V6ffbsNRjH2hweKHSGC2tAz3MzD+IRS3ajoYZYhw57BMlztfCUPf
mUdZdIs5ubVUt1l5Sp3ToSD+mkp8Ys1+85rFDXGydLtTbEtx5EWus/z6u48b8kYm
rqEeS37ZyGfL+MHhtWMEGIuXngEuU2ENUd1K82j9ygk5qkpPbT+1yA1wmgam7N9y
eoEx2MVzXQBMC7+S9m6fjkQK0UtrnnWa7ktoBLZrPueYOKn5geXgc72JyO4EbBf3
Floe6z0Py60ANPkYJgQYuIulOUJULmUmcsdVnKecucXYVj+WDQCULOUorIMFHIeN
+kKcAImq3ipTOS2Z6TtqhcA9NLbANHsrVXhhtkOZJ05W14iv4IjNw1X8VlQCq7U5
JWTDMCEZ4PA0mMzaUN7983uge5LZvcFuJQ6oGPIA759jHTqG5n8gtubBMwDR6Pm3
JocsFXlRMA1fs62QqAJkEFHgTSYQmPCIBdexMPQvcYbOFCkYgIx450kUyEy1O24X
DJ6ftw+APRkU1L85RZZAy1icphpmwF9rlfBQLiQ0IqBxZmpg4B02oPkcOqkhIysN
yLtr50DvGWNAffZdND5S3CeX9g4C2SwWU8kO31wbh7BAnFe3Z2ucbaUDKrGLnjhX
VnkECxMRY/gduoAR7kivRV57C3WjTBd6c1YXljRwJPAJOKiTXp3pV+aQCnowVaOM
9gWxEVqXDB+MlMmhUKDPmaOM3crDh8yl/GHZB4rXzble1aCnRo/OUwri0WZyD+hV
j1ZGnORCpdcBEnYbf8nuo6JaS68KO0hOUD2+aiKt0+3Ry+iM09baPt1/0sBClY5F
d7ppw6DIRk1Yd1DF60o/5WkdZz1tUsObe71a7M/yXZI482NI2S5VNoq4I3qu+PtD
/DJ+/srlt41vwjAW5dKLA/ZNgtZaYoMVvqXlQFO2tNByiAeW76CbVlX9FNRQMMgf
fvNajxJT2HiWDwK3YNdBJVsvvI7oIhPJkQEGfvdhgw9SyncTh8Yhp3qtL3z8F3ga
uH/5G2BvFLHrghJwb2DlUVLm4wr3136o6ubJIKmjbskYZkHRDW9eGQGfAWZjVkib
am5G5ywz3h80hexoMMsuex7uaH7XDfV2DfWe8LXWe0lasTucQ7i++vlLY0xLC/va
FvE3HUK3Etb/6La5TFI9DinT11uc/rj1BwGFnsfY+2k+I0dBv0o4nI6OKja9H3HB
OKphwOUXNLTNVoSiCnd8vfD96eA7lsl3bBAq4o3krHzh3pE+GxWGjezP+uoc8vD+
4TNfrxhAno+azQFNCjXY8JH9y4gahAkFwpbLidZG6J7FNr21goeAH1wRCeacGylD
FKSJLKwGnnzwyqp1LkZoFztBwfaUD4Osfp2iJheMKoPKzqL91ndLe8mGIFjmBHZv
a8M6Ctf8B1rV8XmlU2DtJ5Jl4tMxLNDlx8boB97yTLG+BP6Tup8ySj0Pjijcn7so
uWVqvEc9pEqXMpC33DjTOQC5ICQfRJgSdPSIx0jF0CvL+InnFp+UmN5wi4r4GkZM
lOEYzexZjAViCkb9z8DMrpRajkqu6ijOqqTGzPFVE9iMkW+h2PF5XTqQzjr+xnLF
4Kds6fM1nUhN8hrFWc7Jn6BuPfgwkw51oIz3KS9JOvPZCknBvrhztOyMwmWhXB0y
oS2udE7ktj7N0Loh1DHGETDiX1olthTSHigiwX9DPF0E9HQy7PLjZ4q7G+a4MBtZ
EoXXmtmxxobWQ50HuLZN0sJR+BuQxUjK/kren9IlQwmwPQ2dr1TlRltyyzTLxJy0
wk1sokr2ZOQKl80GjcxZn7Ad8EPFCnEi1uALhO7o0LYPwGe788x6yZMGOVi0o0CD
OBMZ3bck82wICpbusX9sHOd82kuZfTFTvmPefh++5W5hjTte5myKXB1XaOL5B+47
G2IybEuQX1h8KSt6ptFlAtJvA8Fiu8XgT0Jn9JpyKoYTyV50DmXALzhOLmgL0xdC
/O7VFgy/mcTNvCHenrNrbJpar9bNaT/ukDZKNQ81d6GgpY0NfJ/Am0BhTHuEuisf
l5VMQyqr4gQy7f1rnYwNpPs7qdqVCrDmwWVdfNz9m8fT4DdBfGbhjJi/21M1qlbZ
enzkhSw372vBM5GwsLvgWUIGvOKgFLTz6REFHwgyHXWhb36ELFB97SRiCCGXEI3Q
rntHNynNkMVEi1sf56lodoqR23fYOEg1HnxeNKmLpVIlexFvatya1LQw51qTcA52
Kp56olI8BaYU1vrDEbR7U74KzZuDjclIh843vFEAegfdLITTc8JcF8mHXj06idgY
r1Fow58J3AdkXH4Zn4OUlvNJpIvhxNn76FpXbCo1eFJ0sTxLXn01m+Aw2xb6hdn8
Pu0GPtYCdkTtuZHSyUn+2ns/1wjHOzevQfj4FFpQL5lMymRXk+M4QF6rJd2nxZsx
+85oYDJfWiTvmmu1R8hFcSRH1ftumtn4o3gV/1xULEeZ5nm+ag23FV028sfgr0D6
w6UlkducxxN2QX+qzEEBOgnjvI/YZax6B/Uigm73fv0TdhZpq9aAEIgUXeYv2I/D
Y9vmN24YlTFx3HZtRaKMWooQe6VxE/PREGt8VqyID5KLQ2sQF0D6MiZ3QFmgG62W
6CUqt5qqXkj5a6L/fx+0RuccUwkHAwXb0Zjk6H9y3jlBUrdB8KsugS2SpniexFbu
MjFNlA868CK07VhIzh4u46I9OQq2IqCMaQPd+V5nfCVe4lYlYadk+9I/yyJzQNl8
mFroqU0dfofPJectakxauZZth79QCKsTX8PYgW2n1X3h4tVBgVSkt6aaQtpjcI+C
QWOxHCYLIBY9WI5mpsti1akF/4SNjS12bDb+R59pUAz+u2yGsJHz7X/oTxL3gb/i
ZnNREhNPboePLppJYqclIfcF54iByuJD4tvYwpa0+JmpuXXg60JHXzePuiBQi44K
wG8Sqhhy/p0BnmmHd2bzypy9AuvCtE9KAmv5biAzLV385YBkHJ3czeKbUYrIfs7Y
F7et/z09i3SLDsVGBLa07hoZYuikeUk8RPuMm3ZtovVWHcTuit2kjLXZVgZ3Nd5+
iYMEzSh8SG24hiOuF49eENXEYDt2Wn+UWIzzLuvHqIH4e1ImCRlDKtSbpJFIJTu+
2ilDLNGw6h0vKdQjMZ89DsBGIDe5gALWeiyJlBx6Ha2X/M7DhLJ600bZzzfS/Pvw
AdODW6TSeQEy7YfPeCzC4hHTdvtvCbph9InFTAUtX5bDy00XHCYUYBaeOGRQJo1j
N78tNJWZKBKMhte/A1an4GLp8Qf6Ehn6iWVNYZtquugoIhHD2BerRFr0OMG9lvhl
hJgSY5M335ZxQru9d5AGJ4ymnw9BPOOm2lClQ5411mk6VJbPmd33cVnRpyOl4R7l
S7uch5AD0UvK0TWiPXcxUf105x1FF/hOFgrs+R/pj7hhvmMg4Z6neuQn4Jp6wOUC
0XoL2M+3umeah9TTs3uEZCy+hv6n0uhVniTYqxbDm2c1+kCOjx6GARVoUl2MToFm
KTLWQNkMrlLg5Iuo7ECRoyCspDSYpiulYJK5+/YsOD6D5VV1AN7gXEidXJB2xVGN
DLcNQcjqWxxkUYy0+vUkdjI9N7c4Scb1qeWIvROKbXO/M1tHw/2Y5ifyggMgQD3y
EHLcafFJaEMj6AePZrrF63HrKlETetJRSRJW7430/s0d6geL0+sHFZ3ATtwMwkEZ
LMfnKU8g9QjWl4REsLvTp/5Bt6Yp6KCzIMipwZy/mlPHY2RkIGBhqLrtzZMgV6lx
PzSUo6TmAkSWZymLm3gmdRmqR++tpqO+UCW7OkF7jnC4OIkc5vnc1jUGkJzenuZY
CwfS0YE0R0ybuj6dZHfhVh2QRAtAuqtUS1Uncjdx8P1hIyKr98MKtUvZjrK0btak
g7XALCr49WuB3toy8i6P5H2S6edBdB4ZUgJZIbtCrQG8Ypjmmp8WGUhI7bO0GpH0
OKz58fxoVOJdUnvWtl6MUUQYI0KLYQJDKbnry4jB84kvxMEHHgS9rYvpATmJhufZ
w/OdXqtVWjkhrkcSZS6v+r6LCk5I6Trewcp0rkTL/VvcMjtc8fAnQYPuUJMMwc1c
19QmmrvCO9nz4elLkvS+Hn9JS+j+AxS+9Okd7JEj9EFhDKKSKetRy7LolXcVvXmg
4X/BzPt6V251+4z4ZOA8MKf5QBCZ87uzTK26UoOaZgEfCxT8Z/U81YCfYEJ8orTI
GZtxZn4usQ8PV6Qyy7pnJOBiX3a3h6J47EBITIRObg2cDjhNTdI9XNgsuOeg0J+K
3XyH8y6rDhg1lyYnXyqP0PpSGVwrMF0RIEgNccd4/PD1ZKZnxdOWP4nxVcfdpyom
YVEwIMWB1NvFHyjMNdxYwKif5s5XSAAp8/Rf1ggWDkcPmHIokUYRBbKdQpTCbjp4
zA+yb6p/Vs6ewZGQ1WOjlUsAgcZDcFC+bWYh8ca4e+ciiHESWHhhO1QLaUYpS/8/
hu5RGrWNoMQ000v0ZXwpxGLnzcQRy1VRdBomXFShjEsPboy+7XelFQ9uhAeaJB+A
LxSADqv58hNZDKnk0klpVejKiLAnNFmDu9Ca8H4DlgzRvPPIRbl3oqSUYOws3l5s
G3/GTjtqKXIO02Cc7fCbkobb8zl7EGPbTw98II0SWKuc6lRpaoebZDu+shr6klHU
hADH1TLGQD/K5itkKK5XnyxEDx8n0qdPyws2yoyr0gTZJYqwuxIzSOQrJQdV60mB
V+3N1N/oXycCPdqagLIQBLuOISW3XB5BwkD9ekBOhBc0zmeMrsT2o3gWUbSV8ln3
r+TUOnCJ7MpAR/67mtXu/inP/qFmeojcg7rtMJkSdmt57mktleJNSlrlaSEQfN1M
crWR7PvG3kqYXq4j/6TNIWaoIJkB0e5YdNcSa4ZP1V7ap2h/ICuuwReCbmlGFare
hh86zxbQUnA5FIOKTi76sTuMA2KsapSdhR3V2hN6IfUZyUq6uzZ8x4/N69US5hMb
L8VYclCHWJwmZ5Dbx604lYrLMRvV3N7VBKBjtjs26mQ/fE5mCfkWwFHN384Bqq6p
XTXJQt8I2IjHOExLPZoShnY0lOkyMb8LU3s2Dm7ahQH6bcDDlDmPU3fOub8R/zvQ
CoG/teNgO3WdAJu/96sy1mqjOr++Msv8xYOn7htGOGj6r5HY0KPH1gBj7GRFpSYY
mdGtruOUrRAdQX7qD0w9txwAoYFT8dZNR/suSi5TIqaMVjMVNS04fs6Xmk03zaHB
QVdE+YwX0Ltc0XJxe2k+fzMNQKFWNDMi9WWMb75K5kv89KHjSy7Gg6+IjlM348ko
8463rm10WPnJalKc4GcJqUu7pfTquq+0cK+M3o7G+SQPcTDM7ec6WQLsDbI3THB2
jN0C2iij3ytRKjuqFnf3TVT4Z55WiV+/Tc7hSlFqZqp6eoqgKQhVlSjReA8EiHon
iDNkL08PuaBQEk6JOTSFnQ6UrZHqanuBcdhWMO0O3No8PZmwlBYShp1L0jvLODe3
RMySRJm31pSj/jkHPlLI0UR23Mr8/qeAZ5zVqm+9FhBicC3Xi84y5/gxAySo/ave
kG7/ySJ15vqn7LqAP4KjcuQdBpefhodzUn3yk9dojkFo50/B437qgHQo06f6JMvp
1nEBHJnl5Awa0M6gwawic4CaPA0lWSEa9FCie/63GNmSpCk9dhkpQV4KfGhp7DeU
QTAUD3TV6C/J2dfZipIlVCkqFNOFLf0LymR7PDzZaI8Iuxt5glzfVVSq3GKiflD2
Yw0GI4YqY5B9uEpzuIiKrfoQ+Irzk8iJGNnSezTSBBbbiGLt3aGytaRVLr4E0xHr
l8lkF1rqu82my9ZS8+wRX5UXzjPY65cw4TBbII1WWB2SgAm8Tk2VzLankB2ph0Ut
Ox8ePZTaZAVD5sijibs2vvjI66TrsaBsP4MCw9Dt+vUnMEcLMH7iaIdqanmzEUCx
OXzXhbNVtPVfZaDr8W7RkkGviZx/MxBPUneoFyDRNhAeqfvWZJT4IZOvqJ+gf6gL
WbnXVR6lqsYQRu6yHcFolPvK0xhJ7bmGYP6GrAeX1Y4Tlwv8207bdiWvoaUPa+kc
fKu4casAEHrG6q0rtcemL+xarX8CfQZQBFyNDcMZCcqd8CLxthCU76vTr4PmAGg2
Bxd+NQ6ODDVX+NG4QVs69PHRVwzKbX103Q9SlzXtsUoGbTTJtG5S1UU2q8jHzUxB
Dm31uU5L1qZ3iGXOugpgyodhmvu4Bp29N++MXTphMjF+qNj0ilEy4Qx9r7c5cKAm
o06EvqzAx4/q58+0cqsap1HOPPH9wJKYr3md0nI5SCs/UToMGJbzwC0EPJ+zec1N
g5PQuS8uk7jiBeqoQBAYBDLcFs+FMtpGKeKgI1gKEmCgmYUQPbRpxkMq558blWNT
hSvsUklRf7Laiw6G67AAnxNu1E0ZVvD4Ik1z0A3nnJOtfC+7wRi0H22IVGCyce4C
CUY7cgyHBk4E87/psX3pf7YWUZiG9ty1baECcXNoYv+u28WQOzJM3DvM6L4zlxg8
kkTur5VloB9S1+OZyaggTBbIvmMsBHiS6ksCwwHT/fMyUH5Wy2CmLlQ9zlU72jRX
zHfr3HuLIQ4yVgFlvKfzuJViPUIPo16W2YqN7kar/RuBdrxL9Qu7cRBj9rWOzWqy
nC3TQHIXANtmzAxDloa80ITgR0upvF79dZumR/NheBiBZ6+kfPZULo+1Nu7/y3Ev
2MGWezqNn0MQ4KoIzsgn1oJ0QKahjzwthju085JcFlfBmO/BBgNj1e2B3+kmMVSg
7QuWXyyCPX17n44vBqCcH3OP2WYjMzb8qG9qmFhRwghElKjqti5lqpgm431IHhxB
+Y2gI0Q24eTiTPeun+gzWjrWSd4zaFoHpTNLQtmjj1ZXmHPv8afChi663/O+1QAN
GH16s+PkzYd+/Nmci4kG2msXsTnmPQfNwIpiQSi0dIG6UcYiRPXzen18BAqjcA7S
EaJzTsbKmk3ZyAx+Gr96QL+rIg/JAmih7fClQbT/nawLjkN4eEUxNfyOSI+/Rux4
vNe5pf8dYl1fUz6BQdgdjIqtvy5UWBdgsfWnExcRjaKSNvX5GXsos5eXkR+QcnGS
/myGJNbRFZASveiCSIOw/1F0gdLaioaqw9OFRKx9zxboidYDFXtOMJSRX3/yFVZ+
nxaVfdZIL4zMESZYFIYkBtEUYAh2kuAyVT787ZwV2hDxFHcOIf16L1IeGl8mEJN3
iIejHc8do+K6XzqDIaMDDQ==
`pragma protect end_protected
