// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ThHA33O83EM99fB0nVoTixlLgJbWn3UJbroOEDdVCZqvIYJOHDNfj4XayE3UdlYz
dDzwUDKdtFBgWaB7A3sAQ4mFWMgoL/SnL0BxBK2XOn4wicn+Lsv91DKF8UDgedOS
QMhamBvwP0nQjXGdrAjCIo0ZI0VwmJuvt7COj33WkK8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6704)
bMWAIsKe8oJNw4wTeQjNogqcEVezbzZEiUbVvhcz1C4M0R2CVf5/3Mhd9kaB53oj
LWLmL3/B/gCmveUH2+kZNjuK+JebwqtHXvP5MPEXaBY1OfGTfDNDBpLHxxx5cNUH
R4WfR16RQ8Wk/FcTNExAy3Ki7j0BtXDwwbo+ewcPVOhk0gFAAHtYmLxnSmZKppKs
87rGIn+OIa7BquYwr4KTmqXuZb74cUJl8PWoBrpsPjyYw1BxFb2MHg7qr1WGE2UH
bpdULmItbgQVar9RTaffmt5QnZ6KMAcwfelLR99y5opEYOxsFg40KNZ/G2vA8aCk
WHxnyNIZC4EOOunZEQW7+j3MzHyWYAFihgtCVd0uRsFT5CIHlJnR696JU5NchONS
MnoMNc943BHaoHFA7lqqCCZaJbt1gsNl8YDEnjYjM/XlMLGZuuS+QHybDvFkwSfU
8sqI1/Sp2AFZfKIj6sGOtbtVNqNLwOgus2YrNiGm+8fYdA0O109EzKRLzRGGve1a
cg1zFytPAKMp5velT/oZsYH9Usgnip1zDurYYMMPqtGyBncgZTntlyMlyLJn/uM+
fL0e9WRkw+O7HaSvZu6AysyWJB5NPXVaJmB8yvQh/PRa4VUMCZWno7JmsmhvoDdF
nPdAni1/OSqhrlv/xCq6KPBZkGCyA3oRvsGdwRE4kf3ERciM+Uy8wy8d2XIeJfFN
aKx8HXPAKnO/d6Wp9+x04cAobZIMAcZurA5kIO6Xk8kFdw9xOOejb4i5eBQS7jP8
Mny3glEL6RhhIve4140t1o5+FDNiPMPBq/A+JmBr1sNA7yv2wUNyYICpwnuZDZaz
6QSQ7Bje7l1CJP4twMVf7dTduDmB2SA4L0+LJLjhnWYs8M7gok8T/XEkyouXMWce
Qxhvqo7f/aH4VPy8fsjSh93/moPfaVueKLkIGyExriy1VmhmiWbAWCJ31KTrcN6w
/slMRdxlvzovyJ/+XPEnVwe/eBu6Fps/mmR0picc84XD9IljPw1cea9HuJ5tqgmd
BwV7Kd1mANxMI2D6Q5ow/YDQWC4OgS4i8SyqamIrPl/EwS0Zdr/CJU+RVngBlaIX
1Z/J35+lcaSH71YrPXA3leb1f+zoBHVuMf0A6EhIGHQjvxcwDNfWO0wIRt7YociF
QYCl4Yb2yTagNAE85vL3xBXyd0TGeXs5RLi0SMJAVHxrdyXUBfh6ryPh+4NMDO1z
ocOhmd0PwJ6v3r4/zltnU1tr8H1jlpyXMOI89TV5vWBQ9J5L5U+xPfiVbpjyONzJ
nOnaZh0R7USTuTG4u9dEP9Scuh0rQoAsa/psTz1EXn9tResTgC6U60yNcNjn1hI5
Gzq4h3aH3pjnOLEpbUEK/KVi6NBd/Dm6rAPDlf3Ud2yNNWka1m087pVCJam2F3fi
LW3YmMcU8wzUppobjZbBEktkcosKHMTLymL0EtG58aYbsGQnVf+MSS5DBRk6fgv+
hrNbX7+CtoXuf6cMdbzw+7qJMKMdJQ4+iW+NWjfIsaNhZeZ9NTT5tn8D9jlCIG/j
cI4LzS91hjdP/n0/IPmOkcabssmQdY7CojUJ/KBGkMJiSeeNF8rVXPFUyYF3Q4NE
KWAjfYDWjnsPs3sjdBBYsWOaMCM3jZaS9f+DEGd1JUfjEvrRDSJb62CmL4RGLepn
zGt0FSbFl2pV2ACRFSa9EnuinqRH5TBBjsq0VpPY7JQMDI//iE9kcN57u1WzqMIq
SLcyyQ8wIIxPt9fK/nvwt+EDSDkfsG6bnDZj019DwbVOV9zPU34qqiyQuRvYS0iD
2mzvz0BHvKtc+RnVjE/u6H1S7u24v1srJypP85ZFydhVE9bGnmZW+JA3FcgSZl3+
Kl7dLxJyrQOBDuBQtVgZ88TPgPtD/Qe/NHDyBjo0AK4aJwqznnbxafg7c4ip45G0
liFTqKmITq0z56N3KJbxaW7NwDc+xRVPaR2NCNtpi1xUcW4VWIMQmefsUHTbgVEv
1qffRfaX2E3qt5rKDsRtQu0yvHbCxCxqdqaRWgV7q2xoc29O2tJc+xja3/jckmjC
CEgFlW5E8e7ENwQy+zfOIEGDm/+QN2NcmAhfIXr4QAZF+HnHomAttojlrElyAh+7
rwJz3JJeD6RRKW5JzNREwA+hR3CiQBVcUje49zLdp+iLo1wKiyeQJlZmqvIBUePf
PDE6kV4cYNtV9Tad2JliUkKFQS5lZyBqCSN3zcK56CUOm3CjhzigFfTM6sFTdqwG
Zo1/zeTotu5u4vJjXPj/EFNnpDfjCIbyTQcw+Tipjp7zH876islzyNj4XwhICsnH
zxccLtKqJNa2zxh9YSbAnBT4nhQimR1Vk3u2s6TLn/5c1GcsRPi7+rMBXP/0sRG7
Ozr5pzhxRaBcjbKHQp55vUcHC/7rPg083/w6jUQR/RsNvNp2NwtfXMZ7zFJBkHMU
OAqmeO9a9tTWvGXesH60DjHjqvencyS+B7+Yv7xhypwlXgwfrBaqFUmnyNSZDv9/
2MbZr3iNuQmgjVwlY2X0ckKTfUh31+djolcCfwHU5lzjGyyDeM5NiyhNwviC4qYv
2azoNEQ6z+22NprTwSjk9IknL/psb5UWU1RvG6QkbPmYwJERGaP1kgipgWiy8VL6
ji7X9Yt2SLEzTaXQ96XzVpSTu9blhRvxRERYquhQ7GycoF7Z3klwkGkNQyddPzyy
jMoiHVNkXSX7EmBBhtvA2He4Y7h49J8Sxs1g50L9rNFAVvL4WCWLfruI23u7CGy/
x/gEaubw9LXQthLLQvQEeD2d+wt3+9Jd+SiDNP++ObQEWP/Y/BiLdwok2GnD8HxG
1LlQ43w7HiNcBoDfrT80zTm41w+lYdmC3Fj/l4ZNCLiiLzh0SEPsjif9oMJQhUny
VkJcb1JK6zSHsM0Mznh9+E1uSvtyrrFDomRy+0jNJHddHFSKoBtv04M0urvGcgNE
xSAePB6kG2urnE6AUH2VFvbBCq8q0F0CM/nzTUHoSt7NhTUW6a5WGFyF8IQA9jBX
ZNbZByRoJtg4uMD2Lw1qR44ZmysbYiEuazmsBUI770Ozi29fpnANhxkocsTz6exG
ff6ibmwnd3Pp2t/GCWWEbc29+HcK9VHXK61oiNwNMuhUXY5gSnPQaYDoav22NwcD
HAkQvK4YmpSprZKG9qDeXDtWURIS9kwGykpzr1dxBGfFNFiF1KXr7AERh1IZksrn
eof6/qVLXVfDynhn3vELVt5jcM+pO5OIYDVzyUwUPCTe7zyrkSHRDY7oNCak5oFY
asm6jEfGk8XbduSrzdb++XYTcX0IB59ZrbIa3qfYKynfPd1Alc09lBAl/GWjX8xf
5cYxj83UV1zV0G//h/+lnmMMBHdlmoM0pOe2d9cuU48s5ItyjQf7KluXKKWgoqxy
JKJrLN4y2dGlecUWRSYZmMqGfo5iQEnFci4/7VJ2lJaEoGO9De2kCAzIeap16jJJ
Zt9QzJ2jdbcAqWYFcLfW2fAkA++hdzMCzpatsrtAT5PCcUTpiSKnoQqxhK15vrq2
0+p44B/z1AS/iTc/WpdMAvNUf1Ln/T5OG7tkOUWORVTUbbMUp023KjRddWRxbbw9
fAVCe4AuChaZTU1lPMop0BDECxeHCAW9ExiNmql52VD+0Os79pNLoOoeP1z7BYq0
I+Q9KK1Kt3LCEB7IXoKQze7QD6QkOP6wK10NNo/cxP7e7OSL/eIm/ZzQTLzORbJN
7zfR4j4dUY3xvVa5knNB8IkrV6WwIIyEwFeuyE36kSPEIsgMxxE6CUU35dC8Lh3F
fb+8Z7OfbOOvos2S0nBLpxBQ4edz0YGuthY/rA9Rw3vPqBTeyxlA4273fn6lMr3N
YVSAB2qsm2uPDD7I5k1uv+MFU1xEdSdqTTZMitb/uz+mV+tEnIltJY5NvgvtlRog
FILBwe7lxpCeUf628AnXyTj915jzLPPVICM4fa9K10Eep1aiAXnAvJzhXCaaXmRe
ABBipLJhPZUDCGQXIorEeKmbTSDQeLMDSf+nYmL0cflrb5HEAELSjx8i3Y8xoUus
OGXow/wj8eWuPNpbKxYrDGTKmgUrUxpO2Xz0oPYge4kIsr2hfeXXv3RRy1BLMGDi
HFzOfzQU0hf2pPyWHIwM0ghDmDTKWL3P1w0gjcueTVSgVuN34NMlDoKcEDtQhBy9
gFPmqzCEQUVr8786H1DSunUuomhIZLymNsMuJWBoscHuXVUC3mcOE6q2js9soAu3
RooWsdU34gV6jX8OlcglgxMsTIcuHlTf1GB60DAr2BLXSTTA+5U7nQBzEQJOEWMz
Qoc7vlk3+O+OHOjChHhygI/k329cb/WclkjsS4h3465eehNqIojKTKHUlJsydDSQ
dEcUfPyuQDBbJ1zXak6rb4Si9v16R/DMmRhqQ9al+8wu+KUEfRHn4t10qsM4i56f
G5YuxYNgU64or2MBa7aQjw9HBoLKTvT8xA/u5jfx3Djdc3gxBWM244VFDjZhYVdy
+Ako41Hb6PAq/1M9O5LPULaBuYrWQxWg2IuJHvu9lK4rTPfE0kfrf1YGBbBZa8Xm
i7KM8rwbTMPs0ghVyOBmjLNt3qzpCiRC2rKgNyTA9TtAGhkTgWmfEKFFucMWEK5a
Htw9nMew8/oh/wwo+TybU+24BqMuapO6x+SmBCrNb8N+nSs8jeN5mUCreExG7955
ooON+aeQTw5Ehsf2ZhA46+Y+XeAVIyREOiXVXEObpt2sA1OckZygFU0SF+1ZfooS
/aCqiRxSLwF0MZLXrVzCW9sQ3C2k0PQfcBynj60V7GDkaqjr9XKsbkDolG0iGGgF
06E3m8IsjpGj5QMuvUET7Eoj94pkJ+UUXIARRYhKey+VlVBWicwVSgUr9cQD4z6T
Y0lju7itL0TZT/AXWJLcmZ9sjUBIf3pft3Zg32cP3QfNzgyKPrJiMQWl0V2fLk/e
kfn6mMn04xc1vqt4a1GCqe0b86mwzvuItaDsF8LtsBhNTcmMDGawZHgB8w39oAKm
YUmElinHznRTsXJmQskiAs2PPewph9DMt6DoSKdR3hnBxj5Aozr9OT+tlXLUGNKJ
RNiaPlB0fex5Xeom934T3aZVHrh2tZTJpr15tFlkmTsCg595aWuYFug3fbhiVkfW
zWCYVHWICNxI0OrNDFsKvLj+CDadWhTQbimV6L6PYKu+n8updwzZv1FgJIzKWr16
mRN96V02XW9AzmrEMKbE0xOf78tgzgpEeM3baZaJhgNUWbV8u1a3Oq/Ikn7SK5Xo
4VPrqehVJi0I2lEtoJiGNnuxrUL5OObH2HBiI8YPUrfNyRELlxSHb2AMCu7Sq3VM
QibHBK/Rhg7yseiMMW30kztn+xNHUNmedP7+svnSpWiG6D7vd7Xk42u9Xkdq8BX4
e5b7XFWxcsOuIyWSSQKI1IsJdndr6s/7D787wcJEQeIomteAdai0kOUpPP7stqPP
7EZolYLAp0jyA8HHnZBshHMzy/AzlMrPn1gYy498FPy8JovrReUPbVsiwGfQv0fr
n0g/fom+8HC/yeKw49IxIPD/AM+Iyg3PoXCwkdkhwqW+YgnVU7UbBEswsA3s2/lR
XjZlV/PTESWBsr/aop5/ZKdwTaoh2zi+UpPKCcwIGSDdPpBhkScEhpR1wRcEYHZE
uZy3vwI0Il1lLsMqprLT3bV0F20o1SmRpO4medYYSB4Q+Uhgz0pFPqFJYSizYwb6
yU1jrPP+MOonJZFY8gG5JgNisFIrYHvpMT5NKQ37fTGqxsaHTd2vIpAlCQLnEpQs
yaZDTnt8r/Yv6K6pfYK0Y+4ZH0HPr4VKzMx0So5wfW76YXKjcGBPLOah936Wbhwz
slsMp7GEL4HMtysO6v0ygbfj1ICj9tpHO13qTy7292I1UlWW6xPsQ/872a4KCt84
LytMOiOZW49wjJjVZF0ojIZQZVE+lDbaYPl7FFMyyVpnEndOZ+RoKuBBH3VMzXKK
VQGpiADur9FRXnKpWXBYcHNE/bzipI2wXgjTYHkQb7EjZKM01aAYDVaX1DRJguJn
K5xK47PR3q8YPX/4yA2Z4T+Im2EvFlHxMRdFactTRqrNgUJnFqi1JCxaQ31FTM4F
NwpUqYt589Mx0JbqiqY/0VqjR7fq8WQ8zE2mVeXuIBunpLF5/nB9hySHgtNNZnu6
Cgy+YRU8QVrXlxxs8aWtSGi316mDv/mzy2zXMeVE59nYvp5ZzrG8OMkRKoc/WOP+
B44KHWu55REIQAGERTXJsJ0/jAsOq8bJPJ3SwKVE0I0wHhnZ8q8Mu6v/Qad7gtsA
A0sBqvfgEgJ3ADWTZnY+RKayobaMqXzZmtQMbMQ66AiHdqPjS+7JSAfoevvJuAPZ
DwPvVH1fB2Mzxd8XPfP2z6CayJKtw+LwMWAzYuyOCVJCVMHAd9yqUH3aDPWXGll7
tO+aZzXKKDPpMjgW0irxSilw2hrslcPW2Hg1USKNDFXjECwbAXKWHd2EJSvVblBQ
/8x1y/kAuW89ytnZtD/82BGqWbf/kbq/0RbTXT5IfvIpMBul0FUWs86g2nxnGwqO
1ZgGd0eIIkiLxghbKq11HD3x5b9sYem2bjjB7Z17FMDOpMQfwiM0yQE2gLOkXGcS
BvUH6jz2XGNyfHeuv1qKxFuu1M3gUb0TRpQYjaWjq5qy4bW9kZECsD3cSbJZ0HIJ
skrX8hwGq0MsH8QA9JvCsVbH7mHoiCRZXIZsvuSy0p7Y5xudZVXGAgjeEkbURCG8
e3leIB3ouWA2xQkQ4yBELtzEvh7+wbZiPCARiDQH/AElT6n2lyzMvUG8sdnX0Ee9
/+upSoJ/8nLfnXwtGKx5fe+6VZsl3bHg06s0j9mxnk/ue5qqLLrK7YybBTQD58bw
WxZLAy+I64R22euoPi7Kp5ELmwmSJMTMOjJv32ZpUl+8Hlc0iyfvgKC/SOCYARu5
KD7mDtFLr5Mx4bG04g1dITTITnEhD3yu27EcXak3MaTU/7TE2TnzNHJOn85CPY1h
vh321GTTE3QlCyR2MG4iyA86AyYrd0ob6eBy3DrnS3OfFfuT5izVjJGEiall+O9H
5gPWy0fPVkgl+OI3buwyrfTjWxsJsIkQzwmHrAaiYqXAb6TPgV3fqD6xWOJW7Zjr
TylptiAAbWRl3p3g2TT5d9UoVlcx1BboMGuSPpzdplYkp+S0m+HGBFaWyQaZpEeb
a3xMEBb0TQkXf/0vWbgLZK4zv+7i3soCT9HXrjuwu6nPa27j1w77W7PRIySTPfvn
EUbkOrwYjUqQ5F6yNlKhY57T6r6gCJjBjhQxfd3GhT4JYRnyzUyS5X1MU+iMjiim
j9OCCm/Ps0Kgdhg4KsZzPi1CQyI+MCswjCkhaBsAt8LDm3b9U6U6BMtrWGIqKXFs
FuJFHxgbavhrsP0MZGolgGcTNOcVZ2hp3JGEQCAjUgs9MbGIibw0C/uRSUeUic+e
K9Zbz0MZpEQ3hYIsyFAE/fnZCl/QundPCPVhZIVGX07vn9x65XJ079Nza0a9QRB0
/a5ebfoOprNbM/5hWcCkInv75bVNRnPg4ckR9W+cROCpindoLn0y3Q1o4RLS+Uji
0PH1s+MuLPoDvaiSnX0BqiG8fdjCFb1qpgRvlPPS401i+KJ3/oxNWY3RUG7zNC7i
/Df6OYweVGwoNyZ/Uk3rCenT/nb/2dy3al41Elitw3zDhmhD1QYuNT2x2m7ZVGEF
EOEySv1lpbQKWVFq1Rsu8yVtcT+C+HPXc3qrMx5eiClUSEkH4l7NJ2afoLj8+zRn
eXcpDSCGll66s611F5XFZoor1pE7ZkYmSBNAdml+h8LJCjpKNqv9kie/tfW65GNc
Tv53xcNgmg64go7+wbzn4jZMf7EqL3y/yhJY/5LQCVQrmV05j9j0JDTOmdwt2AXn
jyiyvyE2A19dkb73Hb3K84Gf3lO+fFNR889jYQz7TpoDUMaJF91G3fYOCC726RhV
9zjI3PISrnDSrXZ51L2xBxVPx7boCJrozpW51x2jGJfIA6VScbCIiIExmKRneQzM
vWXq33rV1Q6gnT9o8aDXCUymKhapSltRtAl0I8kFOyEwPXlcsf/RI3KeW95T49LC
tM3zn2Hh1zLuaL887q34I6v7S6AohCa318BZB73ksoxore7cciDksl859Qrc1dS0
KLXy34QE2lqN7pNYvu5lhgpXDEFSgimPDYHPsRtOL6F5dKtsX8XOyQmfx1kZiIMV
nZUtQP31xcbJE1JL/l1TtPCuHVn03i+UxZkrSAXU8GpQYKD/8nnbfIvrhkZpWsno
OSnsg7+sZzdOAOHP28L+6CmJ/nRDz+f0IPjgiPm4hL52ggrzzjwMK/f8nm1N4vtb
+tY5m+zZSF305T3DgY3uRixdux/4c0OI/iepuAHHI1Zj+d/meRaWjCH6QwyX/r3P
ON9SKNuK4KDEiSldUucLJ0xF8V2+PJLTtDuYpszbbnZ7DoWaV6c7bHJ3DJ7rQAAg
V7yMcSITabNlcCiwfNH5UwiI1Bb8WPRdhKen37F1JaSagF3uLFqaUx3dDhtJPpNV
7H0j4OVReCi17wsC8dCEi3/CdB2tpIvPXJO1jU3LBcPmyY8ov9pzRFBNTITuNYMC
uGv4UMCxEZt/FDqAultHtc9cc/id1CPW4s8dROtESLqS8Ucehh+vacjbHmtcwxnX
1uIqp1fZ2XmqkCz853SkI9e2KgScHn2h3rpzVH7N/fVF0kycAhuYQWE5bkbSTznW
GyYUFxsHB/y8sRdH4fzfiLcJG+OcdJsWP30VzAhOt7IVKW6d4fQarOhbTjDAg21M
e3phH7qI24+jtCrZrP0iz1jWZN0MvASMpZ2yv+n2u7rWCBe835yG3khGobDGUL2y
0XKM+WSJJ1mPRSeVY3hxN0eXgs7ntDL8gkTf9ZzcJNg96orVPuFq25BkOf1Smaxt
b5QwoQCNCzuxqsuac1VCwQ7heGbBlMkaZEkHU8SMiGk=
`pragma protect end_protected
