// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UQF80dpHuOSQrt2u1vDqdN2sgIx77VIZvPV2EHPqz0ZNf5SUclXXwnclbNsTFDbO
Ulhcfi4HGHCmccRTKVegEF+LuwKtkZZRqB5UYxVb1l5AsIU2Rk7h3P4NuGyngUDD
tDgKbh9EgvHTqBsCnurScZdZO+OEJO8kKYSXWydhkGs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6352)
r+FsuJUPVBgiQ9iZEAAXKVkZwseCIpZ99N1GOUmoiwdN5Q3LAi0vA6c3bt/J/boP
rasSMWad87j/UtqxVn2WcH/yMhDx/4e+7ODqyhB7FQ1doziUuvD10d1NdOZuvbif
Sdf4XhfWX+qnIHoqiito6lrj/ZgsGUpLHMV3nJRxUG6frpR7JFgdmgQs716+i42V
yVPkNFk1oi7o8LnySrG2VKyH5Uv3mk1Y1lnuL4fokI8+/EJiyNkBvI9wd3b+RyzM
vNOAgsLk0OWJcmLU9ETdt0qjxAbQCxXf6BFFpbnbWGMamltBuRhkgLqHAPcKq3rr
bZfeoORN947CJo+cohWEuSXWcB+0I+xJMZpXLfHB9u9MmiVHylipqHIlXgHfCC/+
Rr7FWcs16otA0YiHxhLyiyZqr8gcLScgjdSSIYxQGNxJU3/PCXJEcY1DgVYaz5q3
KG5VRzaMfn+O+YHNkrn99ytcGctS5w6JYyOzx8sdaT2fxIEP4XaI75L1C/H+ulZL
CnPO723+CrfXxW/x96C3rwYuyl54B8G8fmm2nshhu8QVlwUu+O2rzuwyVX9uZm/o
TBzaH/0GMiSpRhjn2J4UvphoqjApkk/KxuTCUYgPvlf2IXx5mDD55om6bqCHJLUR
mZJJQl+QgZVsRq4iPKRcb7VtoNQXnLqS0kabhl2Tv4ABjxLDFaL3yJn3lDvM3x0e
SiGDVb7NQc7xJ0STL/UuaA9hno0RGQv5mLfPxW/G//kddAVbpifP+vp7aASRdGbh
O3dZqKyPhutXbYMupQ5dZ3TBkvwIZiqrRUhYwFqjY0mK2ILAfSsGYYhGhamMPNWB
8x3nuH7BKBxPm2jkfnsM3p17drh9uxd8UwRVZzCUNo4ozQYhS9JbEyPvkZUlM08k
AxkXjxNH2ePyJBgsuLQFYWgWBeW+41UdBEklxtyj0suB1O49AgnQV8/8IcXn1R/l
IBB0V8vovFXad34UYlzDKFXAcHiFpu/X2CTwikkYYlr3QGQlcvJlXeLDZ5mfBRNv
x4y9wgE9cxTqZY41neF8MrvTyfFADCDAvvztcUZi+1usG5CrniQwtRm9/v9uDKwK
5oprKyX2qJSSGxs1VoGALD6e/+hXL6U0PZFZ701j6rvh1IzHtIIqyllDXE+Eb/y4
Kz5cY3SmQ9jSTq5mAr/0u59buQzLLYhimQUk+bnz+e8tJZGHwgljaX4Xv/nnTWVZ
UC6UhXGc4fMcEU+Xwqxide7T56iprm/ynwJ503MuGMN4QThbUK1iamtuix2WKWjX
aejHgRqDN819WKDw7Jh5hv7waOq2OlIkkEqFSKXlhzx5rE/No5qxBRTllmrP/PKl
oKZkwV224nE1pre+Sejy4RUDePbx4vz2HfE/2z8+BVa4mHR0WaEcWBiV+ee5WSDg
jo2xtD6VEpXA0HWOuVJo5o59hOkPLQKpa66zFrLQx8JCi+XHAtaEks2l3Yz1QD9d
7oAmHEt8I3ijLEIq9h22HHzm+mBt331eM+ptUPQZjG0P5DXn1NjOAbDhPx4eOSoF
fQ+EprlMkKVEunHBhT+G+8yXzKiXJKylqR2cfMz2YOuutekc3dbLIYgEuhPZ1PMa
n76I5bD57DT+rSkBnPGMMqBZBN8Z5ATVVHPrD0lKYGLIQDG+gi0+0olTyN76Oboj
vvigRJU6zbGZABY5o9XD7ylHH/PSSzVLvnqvmNYgkaRBB4EX+qrcn2sKcTtkHahY
zqkTitcxqTJiE5vA0DUQgoa3id/px2514uojTlkv1OWmRVt99KdjPdTrptmQNKFS
ThyAfJ9Cy6r6ksaDVI/p78ub+Ekn+05AVPjbsivGQrk6KH0QiCngnsgJVlg9kEhs
+bRmuWaTReiA06wxQFrMzmYBjBaeArug5NdL3tTv/4wd+10lBcdbizu1P8wIf+f1
xX4T6Z7+ZNF0qdF6ExoDqPRm/D4Qc4CQSkGhPxMQ3D0EYRFjpQJ9xKAmmFSTVyxP
hCnzc85clp46savMbRZO6c6OVdktiDu88XfwoPGaeJQvLh499nA0SslpoxP2ICfb
r1epG/t8pSs/6et1lfUb3DnAexyLAib1CiYzAZh7BNNuXODi5zMGVVibda4HZtK5
tMlI4xaOcnJzyo01eqJBEeR+OsyA7KeUDOoR8HtVbB1uTFcLeyIg62rBWgboibQ5
mhTRjwVYHGBfzbD0YX4l17bp/8EwpqeXiBE3eVSA6+UG1mdniL1OvXQ07X8j2C85
ZZCTPpSt7l4yAPeLS2nqXcOmpxCypBb18NXzqpc5GEz9AHXIK6izDjZQUTyV+tzG
ApdQH9PU6yXfzjnVSOkNWzNkLkydn2mXqT3rzhTFp/iW/jQAlFbQxhLO2HoCoEBi
zZPWQ2KdQWnwSwoNBe5N65oCm8TNFGReUgfaFPqfWrW3xlmRqQG3uxs5qmIXzou/
fWGpqx/D9Av7MZm10f9DHTW+n28DiJqwqO22WKXMqhTv+4w5O1SJihlQLKBiTqj+
XhswoS9vvTBVd7BHpxWJgulpr2HgwMoEzyJC/ZKVk+QSWL4Ni5/9Z9naeYHGTHaL
gv8UbNABPI5NQtoBqdkzXNqI6rghEzXNQkdNhuOCxU7uR6N7lrIWOZM5Ygb4CrzC
8waoUTXfuiyaluFfYBYfNp3+dZeOHebeaBL/+XAFDSx4dVcTFIDNGUtSYEfLYsfv
E4CtE7Bkp8vdGdV2OGZ2jkl498PIIMvVyr0hD5MsF3mQZZoRZzcO8RdsMxImTruJ
KRFz/mCSqPBlozsFPX1E2RwYMFCf9cWA/Ym3pc8WNCOALtdXU3d8ZYXQUoz2ADxy
YKFQNGEKvg54a+KMRX12iJX3yKCFSsmGHhCVz1VBbz0lVtObA5GloYOs8iGBS12n
GjQS0xpCYy+dMZb7bagmfRlvv+8reuBqGH+OBOBmTbuvKlODl072Th5/ajHmGS/t
9BsrIoAJhyNagWdgLPGqgefdXd8s4tcxYUFM+elU3UzveXGmaTyMlyPTSzdOwjd4
Z5YQnq8KZ89Grv7IPmF771ZArvbynZQYsTKgzj82gQZggyawOETyLfDPIMvVgp31
inaJ29kJ0sipIHphR1wHiLzrsw9sdBgwtYd1Uqu0x6ECEWffSg1vzmU2Xj4+XRqm
+O58mluI1GElzG+c9AKrhkjHNKNPOwe+CqabOaB6+S679EEJiJ3i4BaXTyWgZeCU
tIAS2X3RWE1hpCrAf1ZzpXR6onHkxdz5EhRwDLp3O/YkYEIQ1T2e1MW/oizgbuyx
0Dg6szb7Imk8DN/Uih3XE6HZS+TZqsVybWBzQ2lXA5fEhjKSzaJdZC59GqdpNhUG
iLO8h9UZNXkhxJixUeWFFdRgnUT3q9V7Gj1qZOjCfTDpVaYdGnnI0c5wN+afofQ5
kYchdk9vUdHaE+Ox2RofQsy/RMuhOOd3Bper3jemzl8y3w7JuMWLVi1kqMe9GUUU
H5klqFrSLRD+h1PB1jj9tk37J5AUrEu3JyRvQey7Toq6u+Jr82JPvFPtpCpyOeql
GtIJ5JywzhRNQRP1brteeO0N+Q6Es22QADAa2FX6MyhqyLSa0aHawbDO8RM5PKcm
8EHqSTCauOFyTJFWxsVNGJjGgS8a8gYLHcmHTFnhRmaKT1zP7bqHzWoS0Y8ECpRl
xpMMovT7gNCaT/2QqLd3IPT4R5qh2UtZHqgWVJg4cH2sPH7iW2arDljk1/Jl24nr
hc0FrJCpyg6bwTCqlnJm1hsKZy6gEhKuckwqs6GSmxAX/hzs1Kg28lwdUIGAE7sV
UX70WlUvhPJXBgaLfC+e3uW4QF1aNnXqMgwRlu2lz4zBqxEkDCFNCJh3xjR1cnfG
qDlPcJO/phWLfizqi11NPapdH2yiAO6tp5LiZIrZdxU6sEAQRUyqCfPU0VLbHtYa
ezyhpLy21xQwL/3eu0KCORyMsGb174lJTV7OGZ4PrDASyiq+oN3wUTZvjEMLRxt7
tIitVwOFfWDsoXkLJ5zqNy8zIpCsfhFTC2uvLZ7Xftef8AFzJ/bvLpJsOOR7jeGV
ov8TTU3Koc9Euxn/2pJItOWCJFD/iAAlrBQDj/X28W07PtsyID627Id1gTvSCgRg
gs4dzmLuSdHny5RAzlvWMTUf30r/bOp9GAk1pRfwEow9+2jfYhOTc3auDFfWegWc
0F+Kb5NNY8QzgP6az5QXSCr18EkE8whvA2kFv3DGSa5GI0wV5cFvayYzzJfSUUJu
XQDh/ZJzEsnf8iN1JEAN5rN0UOI+M3mJ5dA89UiZK/lgiTtP47//OC2i8WQJStvt
ax2HtTIytqLnJYmg3ul86PgReYdP7Ao9Rlr3J3Tw0HxlBAGvI89UmxRB9m6D74h1
b8zVUNVy0VfF9cdEfo1R/hJQBqvg0p8Cjkzm9KCHrZyrJ1vxa1cv7w1Dvnx1E/MP
zsD5CTUaB8CnO5D/FB19ySCKZK+OEjR5tNAEWubAzPE24OLfvxVIRtOFZg4No1kd
+sAWi8jITn/6KZSWjbrNrrx5ukXBJ8BkfgJVkRNNi72rPfAXjGz9xSYzjAVgjgJO
A+mkXPYx8sm194FWDBk4duYwUQCFVhzwGVjQI/QfVa0M/tFJxYapUo1XtBS6CaWp
dztE0a/uLfp8b1PV/2Q15KhlCHokEePZOgV8YCed97pDuYvhAG22YdP8BJrW5G/6
HrjHJdVhUG4eZnz94wBLprqKHocaa05LBDE245CEz/ignafmx/PYtic6iiobAOqR
diqIXpbIbOpxTKLjk/HjhVFqyUpqJINz4VA9i2IIW9cDSaM0ILFGSKxpYIqdzOB+
BpL2Eh+8EkR0v+n5XbRjNyTeioXG0Dp7l0BYWEt2oQcfTyCSDihqTquNLdy/anST
4Ju3dOpXt8AAmbsJS3namiKmOvxlHOBlgqOBXOB1AVYo1oNAUI47EXmxkl0s0afd
jwY45bUg2vFZWQm/l7DT/99o6WOkttUR/Ij8NIxbMqhJ93UBKgFavZW9Tp26k9lE
/EYhGpnl29COJqXSBJHlMPWJrr/VV+xIqJe7UbFHBmMJtqexc9HtvkLPG8v9LlLk
79EyVoz4ZHIzAXN0OcHF3jEHwzphHHvQDAsfXAkMkCqI5E527VOty2l5fgN6VgQR
BvAzcK2IaF/GZHicMRfnu71wG5bILuuIpHceWLh8k9/Bu/xlVrCBDy/eeBTImfL/
220ST0pTBohEkBpPy8Q3oNQo4TwZvQbJ/G5GMpgeDMJhnYC8hGX6muanUuKX86FC
MNsfRsQX4oXu5tq9m4gcuoiDpXyciF2c8eRWlWQ0r4qtweBGSxCFSdq3Nk8jZfod
VOtvNd9UrvloZucVHau4XeIQE4+V18IVIBDa/BBSj8jnqZujMESgUma8JAzlQTnq
pIlxO4NHYWUjrXU/f7wzKtERj7KFamyl6TyMtyBPI9vHdFX05oLGrNOcD6C640GJ
1V4sAnaViPgRmbGJ6NU4iisE0wgoVYd6P6DJyVatEqmv4NNy1pMTtyNTpi42qhxl
dE41Ie8Rd+X0kkw0cD02SGvpGkHhdep1NdgVk1RHDK8CBq+Tdz/pJuKH5Esq3sbX
9bcyHQLPf4pT/PR7hCAQY7QO+qOlJddLeqBHx02Qp/lf818JYdXaELt3mRzITwdG
vnRpdqWUd33HsWE4epXfdNX1BqeY9E0NEM78A8wRWJF3cBYHlY+AeoLle9Aq6xOZ
jK5aSrScTrJWN9a9UJJ/Dp/0VXDE58D5AonbSLwqycA3WK9C7S8qZetwK4lHAUta
fbdYa/9/E6BccicVNp2DcKL/w4dcpc0MHTOr+JRh9bvOmfAv8HTt+MDWX9DeM9l0
AOm11YAn4hyYdJtOI8wPiA0myndf9OxW0N5iQfR/5u0ckn7N7qBj1KDG05qxtmUt
dLx4BkS+6talj4asnTIy9m1b1FDDKtz1fn9or7a9G2OlFIsdR9gtSfo4Z7fyiDaZ
WBNr1O8tn2pC6cevVTFyNvjmSErbaQzyLWrr4wPZnwcsMuiJRmkGyyrXW+AdhdXM
fHcxmSkIrSVDs2x2FFO4UzCQsRpKxdpWIALSNaL9j/EhXiSAbdfBAmbNAOMWgVNl
LAsyZ4B1yFHF2uBdaKT7V+MooFVtNdR5S0NS50yodnKgfn1ua8yzmA2JQ7MrCraU
skVYhn7NK10uRUJEiH+KHhay1Gg8XFEE7XjGmQx510MiptXLkxEmCHB5ijzgIVzq
IMrvXtGR1wO+mO/fSdmhbZx1ZrmeBnyBiWlnZMAI0g2UX/Uqv1KQeu2Eh5Z04vR9
ByHitoAMiKiaEeztADwspzBB6DU9K8WebX27tvvo2h2GIziSzqzT8DTKYR0eBqlE
GW8j1H6W9y1iUBZWZlls1Zgs0NeA1puk30Wulyqzq/1HU2GP7EyLeR8MLQE1Sg8I
+2jtia9ewTqLKtCbLKbdnkrJBUSgWGqitLigsVAsrzgZYvFQu5nLDewI/sFFsFqB
jcNaZvmWTJAcUrEnfqEzYUw8CRYlbVVVNCl7ZhxCDHOHfo7+KeCjYNEGdtyN5HL1
krhVeK9ObvqgG1/rfFF8GsbyxpKlMUVosIv13f4f+hg8z8XRHoyRfz1zN+Cf5IEt
47bsZ0/nRGn8c2naq2fyW6Rq1dkPzipgVtPYH1+AoN5zuBUoqP7gCOK9a9dseUfq
d1LLOKjsS+qiy0ty/uvWiJNvXglBIy5TX25EsNkodsTEW0L2W31YCMR/6spH84HS
S7Z5HhxDcqBUfgmETQiZTI4sxmGzPY7NnD0hc+xLcnqXKYjc6ljaAzWEpxaMWBAK
xec/uIrURuUNeHBm54WvRC8gdS9esmIv4LOpUWSnxyFtc/UJ7GkFldqDeCOdoCSr
9VGejOXbPqXnZMo9A8iXscWAd5vAFqNR1iSofuE0lmssGBkgsvBityxE4plNCKHD
JtpGMU7d/34Htc5h1h0DkRTApSTIAU9G6l8k8FNzU3wYRtSnLbnPSAu6JhZGGqWv
rmilBBaHHn+oCQpSwHrI4eh+Mm4ChzCcHpHI9wHO2FPIfKTt1UnhU92Vnu1SnQuv
lpSDFYTOjrYwjlMouCuLdfy4ST1CwNtRxKkSwTQaUu7soIlNwHBCYfo2szjd+dgU
JZrXo14xmCYqrZbye6rwRuMW0jEG10nViAdjp7qNCsAesRKW1f/7Nzzzr8E4ACgG
cXL/jJ+QP3Oe2yI8QKdkMHWSgEfNHh9waphqeS2HeDQgaXcjcZNsrsyBID45zIsm
j64/ljNBHTSGCNse+zjXwFTDP1YkPexWAMb9IQe0YdDUtFWlbrT9AikOdkiU3k/m
SNUBpXgeNMvDJTCVrJe2wQUOG1VkaYjlI0gKNr34ZrvKHR6VUbiD+rYj8n/VK2PU
V8+C+KYrVZ11ve3Qvvl9veggXfmP3mf8fizwrgbRKRJtb5KtVuCWiGSHiXd2bicV
KmAQg4UXRtsiVggHvICqqFtNp3s+bjWlT5BVv7KwhdA39nfbjKowC5XMz8Sb9gFk
xul10PkjSdj9Rer2p/+hS3iIIuOpyzGTYMW37XVwXWiMl0XwiNE4ZcZEJ/vLgERB
PdxXAeLg3zC3NQggAKxQu/Qea0gi/FvoQ47ZaZVrG6T9l83kQP4K6ZgG0n6QuLn+
hdHxB9Qd2XuMeesVbTH17ZHrkS7Xhft2g1BNXi+zc5GD2aPp0L3MeexOFtL72lw9
T4c4DLQ2FK9E1wdpkoT4aQwm6YARJ+TGGu8pvQM62avBqNoGuM/qu4I6Pe7971W9
yPZfWhsCn2VP6L/TVl4RGbSC+9gsWSpIX/ffLtP8WfstEy+5ghpqXq+wsOUeHoAp
QhWTrBrRRMhPUCZO8dYnBbPvtUPRnYgWbI90fxr53A+hMLaTi2M5in7myBpHYMt/
UDiXXBgxmRZwtcHf2sCHmyUFt2IwN60evF3BBLVMBvusJwcedMop6rZgedTLlSEG
vSwNClGYkrT6gpHYn/EeBE1CZjZ6wR6FV6vzXbCyoXMYdKJ6yfDyaL3EYPgMYMFe
2LAKGPArkD49yo7m8izZzftdVu1Utcd43VTy/QKvoWAPbAzQtTh12skWRWDuELV0
pG8a8B3RWaP5JOMttcl3Lmswxjrx+lHliZzc/VrJu37Q3BeAZN6Nu79jDFY+7w8/
mF/cHyjmH7blbwLfnOua54w2BvNgdnlF9AHGb/OqxIIPNf8IphwIlaFeBmiS6x4b
ZXROdYbjkIuV1ls+oIBRSFyti3wGJTiiPmSxcquLks0MV7NLRZADxldaB6HCgnvm
s8guuzBcYy8zJ3Xlecu62PLvs2i4WNpG7H2uNyJyHWGzOg954jq5E9SLyEuK6FTU
+kBOL5s2NJnGHBxyj4L5G+vuNujCAM43eTeIQN8WoS12Ni/WW9hQvAHhFD1dlKCW
nzlz/1/9MRPASjKU1z1VtDjJGsuEF+Ya9rZLB+GU/It+AHIpX0V6LItMubZKffUs
6H0iBEcI3xEdTG4CrzgKiA==
`pragma protect end_protected
