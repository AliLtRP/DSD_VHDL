// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
q3HIytKCn2foDet5WJqcYzCL4AXRAUTqj72NJo4pScjKzWZp5Lavc2M1/RQBjTAn/JiDxsPqixWa
A8o0RmmRQLF5XcojME6wTgCxB6lNax3ZzcX2//NmNTEm4QL2tnWNL+vMxMSIqeACfDNCFOspvGmI
KU8ct8LR6/4bAWAl4PjCdd09s9SMIbqaE4UZ4Bqbdb5ra9o1nl37uV5SCSC/4omlhjNiVPL2AsW2
8hHbVJfU7qzPUjKQmuqcvRJuIrsyc7PW0dy41wSLI6RtUa+DVXqXN+lpxywBZL3LYi2JduaRZh+2
rlHQS2jc9Hc0FDD16XA7INFCeACQKFS4J/o+JQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
6H86P3QHcfhKNU9ZYj2EGGAbM1OMOxKn2obNEoD9omvb1rZCQx0a6mF9EQEhH/qiwx7H8yfeJyQ+
RaLBobOtMPlDmnCldEhY0SCXJzRPbVKeq73eAjln7V6naLnCIz1OnhuS2/DJsAYbNBtQoDHwIEv/
wim6RN2kPmA5qxL8XS1di5aotNoW0cQcJ8TUzqT+kDzCFdrNq9RaoCYVU18afwqFKcQNKYUlXXeF
3d65JuCF8loCQEHyDSdT5ySUaAd6ZterpnUoI605vW0AC+Cf8zv34uoJDhhdTVP8Qc8UVdTB83n1
Gvamo4QPyVsSqoR1WDOmT9j/18J+/1FY/PIBB7ma8YGPprV1V9cKL/hsbBkuA8PBbh8bUHlQD8EO
Pwhx/BIvINmpTRwpqdodXKqfCLyfJ0Cb+hLrJDkcWr+89MEd22WeW/ieVrXTtHPzarWMlI7WG6m5
gtBFxUWqPkuqEnqHpl6RFM02FNBeoR5sTRdkdL3gJuiBFWQ7HkoRPRofkBbEkKSVjfg9MTcwB1bQ
6Sg7DlN6BDKuz09NpLk//Dm8W5KohzUZ3uLB1SIefrXkJ2l+Be4tPfvX1EvDYOm32gJA3i5gNbpb
1P3cm4zxGl83daUvOmABT1qN5/oM3ZqYETmm99+cMObEfsM2tnxao/9Yga8bjVxaKBWjPn2uHWMu
hWS4sh73IhFn0vemJytCyRdqGQGASPUfiwuvu7rWhmkOBNIanZxr1PR58YkELrsnUFvqrskYfmsd
ybx6W6Ktu6OOuXszs/fzAPSthuAFOHyeUS7w6VoNspXAslO6dr3wyXsnDFU+TJ4V08S5o8+NGigv
Q269hzV0FAYPX4eoFXFtxuOS1sWPphBHkPveir3GUHo/Qs9SDnS/2PFlAuSf3aXWmcGt9XDcEBHe
f9vykMLvRTCI4wvhc9hhpi4HZ9XYevi2KACaEP4aUuFvsD1H7rY8cBc3zPVtc2fO/GIxNlPmGqj7
XoxHMkPW3hEqKKKyLFHO2q7OpL8kG+W3Sndgy1+i0Rk3Aa3KJKL2kzl9L20DGbdjvIES9NRVpTcH
Bpt0QC/8yoghoBn+BPTYcEqja5OLKLmqCEnC0KSaSYRMYfhYskhhWyrmfNn31UQBB/39ElP7yVVB
S0VTX3rd5Vb9hVeAvIyzWdRlEJJ4aRkNm/hO7zactGcjGqjwmUbrCx0Q2UN/YsrSD8OsS6jSe83E
dPuHTp/u/F3EiQr0OezSozXogla1GXnwPI9Uy7Dmb/eRc+wkzeII8ZRYYLcgCatZzsWXKHfvomwK
huCt+3WIZO7iezbwuY7JKLYip/MeR0DtONsXYghDTE4W/efz6613SsYmzE25W2+cWoR4aUljjT8w
57+6NvOGTnRupsXQEo4Os7qX2gSDlnTpLkTTf1ymX88rk6kYZQTKOGOaue7DZMkIiVqQgJtd6aSu
r8wGGaz18/H+AZjXLGwb9J24uWNov8OKRS4j6YTmgdJxzrsnSOIQiUzG72r9yWVgnlp87qRizZp8
R83vC6Wqp/lRoNuXP20Belp0qTlock0B93X9Gy2wsR2bGLtJJJLr5fwN+U1ISyr4pMHF+/RYMQJ0
6Y48KTavgeGyau20aIgFon/I9MmAvyhlWIeuwMSP2J2DD9qikiRy2ufC8V5WLL2tcESeZgMqJ78a
sG5cdc49Y/1h86MOZ096hAYgvcGmnihMOv1Zie0TkJmT8Ttf3jd9StS06OSnoM5AQUhilkXFACa5
NspkWPdXQJOGyhaUCPBEtfmeHrGrpFzZQ08+8TEld5JPBSug07KNHtJBus+LLU4pqgsSkzMeOOIO
N/HuzqBc2vWgRKJ2tbIrSnOpYfv1S6V0wcNhUgiJlPr2Y27BpiV5dIA2u83ta+c583ZvWRrB22jR
VupAuvDL19WcMmMXn315xLbeGBXMTmg5ZUQr1O3w5qPN7eazAS+VdC7eom0vldm6soIx9Vjz3Ef7
lbKLMKkBZxN8ps+ZmoX1FHKHvmZVqvBQePcxUcdSUWQN+iM6ijX/Y3ryHkzgpWm4u2XNhoaysixL
dicw8VXZc2EcvKUSdi55vZlnLhzzzBVCnc7vxQdhVrn62M2e029D40Iwq04PR7Gu1LtYH6UpxDq4
YwusdyLS9bkVOU16Ljy5NN/kHabpP5obeTXPwVB0Ew4EmHZymI1Z4ydhGA1RrFER8t9nU25BT0oX
pPD7OajDbySBUqPpYocG6PAEq/9c+1RMoeZzNsgXc9vxAwnDYFlEVtn5m1/6+PrbfjpKI2C6B7oP
73V4iEVBKVOzfP0Ch8Ipngd6atbRyIJYBS7+9C1GZyYEnIJN+8XsbK9d46AdJQlBTZfNaEMpklQy
ineo1gYKFsb/OTNDsgTn0FNbhhzwnujWNE3LZcYjLWyj9NA9XHhX6/wmJF38AjA7+La98l1Zu0vp
VLFQRqtuAFayAdx6bk1tyaBTrIC2ioJqSgqTY/6+6v1HRVBKCMw86F6SAuw9ysJ6CT4VaBkesY5R
dGP/DghKvmff6G9uIoGCWYrqeuskF1Gtz6FVu4H1vVegPVQljHql/pWYa7AmF0KyTCwk55vfk/SP
C4h3ywxdEQ/2GTd7EiJ4vA7bgP3ZvhiRWjur/4mymnPEiRHJRWdCOYJao3dX8j9vK7r7UZEg7mfE
8uCDKLoda/anwfo6AZ8Xuk6Pt6w0WCOmbdPpYP25eaOtOfVnftunDN3tv558bJCQt2Mq3HLMVvGy
ZEoCGUNBg4eH+ctw/HwMf96eFX+tOKPyi6zHtH4k/sbrwHOoBSoa7KJ/FpchrHCIISgjkQPObFcg
8PWL2PYTkP7aC1IZY/dj3VDgDSOBP6Tjk9eFNoVaiq9LbB182kGajqjE0OOEuWD1+UL9DDRcriSS
29pvSwSPwfaqEM4xCrfvICodDPH6SXtIEx7pWxTnAI6EibXht21XF9wkjNVMH1hViQHS0HxGqvR5
0xHZYZuRPv9OHYzm07zAqpd5/z0GxLF8bhHwUZIAwjYwU057I4SSCByUz2pXNY1R1K6jTONyUMk0
T41bZ8/WiNNonB8u9SCoLR1e6pdl2xr4BzGBlVMDc5RLZbl140hCpW6sQc/Fdz4ehErgPzy4hnV4
tka/ptY/oixD8beWe3l2Tyj5QdsDAQl7DOenrznCyQLC5nAIDqq2SQkCrdRHNq1oEY8fNByWXTK3
PwPREOy9mp7QAQg1nVaoyt4pVC5N4WWNk0KHUb9uxLdOvDeXaPoH4VA8IGd9Iatm873dmf8oNIfD
2V2RkOnH68enU05g/FhEob9VEsrXkYC0s8SYveywsf4swwKuTPFVZTwQyRHR5Em3cF+JWXmyhv3r
2km3StFrD5jvdaJJ2JI4QbbZrZ4agEzWJ/lJ/4C4PauNAwXsQEoorZK6+5bWLk14FP35XFHGV+FK
A7oR3V369MR6rn8vCfv9QfTN5+VUxFkwCTHrIfarA5qjHWyVhM5YD0YWP+f7naHSog5lYty1nQNR
/rPpU0ePROVvB+nHn7a/9qHUGlVyUDEwYw3CUWwfYWLCOSkJDqOMUw0+W2JzvsgH+TNCohe4rU8B
e9t4rmxDa/bOwDcRVoZNo3TvvQ2nm1tGo1Sv+KlU35bUpQ3FYnxfksuhTRpTxGzqNlNxVAGnS7Yz
qReUgrmIwaIk3aPBfzmBDedL3wiwIIiKThHKhwYy/0N0QkhARUyihvcZC8x/VIZ8HBfFfjmpOZs1
6DvPKpDYeHb8qTRuepqPzQboqqWnUcrI5GdfW8NE+igzD+Rc36Gltk0w+NwsGJ63r+n5fNq73RQW
/gk4CttB3xt8F/JFx0pWbOFayZPGcEmo/oh9F4bt5Y15DZfni+ZB9njfNej7aMH6fj9Bu2AWp+J6
SZ/brzyFAehSKR6iw3qz4elr7G3g1SXnFUCqavdz16RMYyVIqgwoFd67ZRuEHFe0LPub/DOlrtiN
zB4IQc1BLu1tKU4yJvmUzLL89IRZm8ZuORZfiGKwZkW/VKwkolP3ncJOJuZ+nKPOlA4Da5DIlilo
+XNurfnoZjqplVSuDfCJtk4s2AIjm+CPy9cr6dDCsUawk1WQ7kqmvvDb5+Cbo3PSqQD19YSGcaBu
VywjVF99r5J5uaU6TJGOgReFC+Cu/srBh174X/LhiAbat2du+coA/PvpQdO3JXxpcVKHYF1OoVvt
0sbPPxZYCKrmrz59hPLerYR2g27slKmHlOqkmPIOS1Ij6zUynYh87E54DGRFn2Hli6IYhqqDb0Aa
nKSdmQdZlLeta277Cvxm1pYhRwTXKlDqbtBsbjaMBGZmPTD4wx7r7DCyskaJXE5Hbtn/esVJK7p2
OMG71GPNpTnvrH01noGQBvorFcU9ypIrK5JMZhOywGorpWwabLDLLjCigB+awRlwWzWa/xxu9k/W
EUOLg0PeyXP7XVSF0FhiaRcKnEwpiXIv+PFBfnwbrHIEv8hJzrLQjoWpcm1TgP49InBUrZld6+VS
Hshtz1lk8g6AdPTKtOibACT7BeNgOyBCr2fZQDj31RQbSnc6ePiylOUxB0H7SjHDuD+E1qO6qui7
dPRrVL2l8RcdtcXtddhypWojWdYdNXsMoVxJnNHmW7LEKW11ffVW7XNt1kI4SXJqeHimtsyiOSE8
DB+554Y4HQqrRAaso1G+oNof03DV+cxX6n5X2mXHqq5u69R5IKZWtIab3su5beI+BpxF2Czu6MOH
ow5lXNOhHs9P4W0XcEd7fLJWaRgZpEDxPFJT30zaHFtOy5OKLInZdQzpvIYlKWpErWv8riv6MYTl
xdyNKDmSOnLSZ6NjvMrl1fwW2rb6JEVlHF1flUqAejGQ/yhRezt4RBhI4jDR3hfgKDhl0ixSxcQd
uMHZ6CLYK7SrzZqW5rAzT3MpopPWOHxuq6e4Czwm9DBbk37L7O7Py7l+EYyDaQBYQTFvaamhcg/q
dwNNsv/xsrcKpyA6LVIhRQDHa8Hy40PGY4qx6QGhXgMXygzS5JROtL7XCqIb58Ib87RZXFLaNtz+
Q4182xO6zzm27y9gKj99z+um9yr1g9sXj1WhuL5ihp+S6/noQ4W35W2KnV/CikK//Tb4LTPamsoo
XV4RGJiVgDWh7xAG3Myyr87dyOOJHVH+tPiGT9Zyeoxkwwf4/O8S6XRCZ7HuBYzb0h6v8/BG5/P1
7blpMujBeUoWbVaFYjkx6ybcqiib8zqQPTaxygXyyFXcz36CAAxZQhIfiWMuL+hkOIib7XxK9pX3
uGoDSsiKqaY/0uiQRHEdoVQkyYuzADNwm/cGdbQ7p05vyKXrWZwSf3l8BmBT8v2YjCvoSvPo806F
UoOdMuHtFzaRg+IcMlH0ygNAM3bzFp6Uqr8HFCPAtJP7q9X+jDdRNFE85igJbUcpLfeOQ7qIUqyN
/wxc9tmyOQBj2ap0Zr1wo2y+aF7ayKuhwjTrCFZvl3SGVduF7vA0fj/NOKb5/kuLJsJomDsKrXhm
QnyrfhScwaZbN7QpGW4SMT5DiB9SRDxrB6yMPOR3lN5+xurU7aqeLz5xSSleuDHMe0ljuSdEtPDy
t70AT6QL7rdxG0wCP3Aci68SLFFx2Y0EUAYfYV0uKfkfRZHeI2q8Yu5qaV7Qn07CYFA4s1Y2TTDC
wBcdsUYnAW5QQXTj8PJW+WIbYptjNRp88a7m7K4KZF4F9Ov+l2RgQsBI9YIfAboHA8bCWT3ObxyV
5hdb1r7sRyNEPJjhsjN1BB9uWOwqK/lAMp9BUhLSjgOjVl/x/VgOmHSu1Vvi6Wt2HojtsQAMRenP
ooskjeV5AKe4aRLVRzTt7vYYz8XmXvqrDz11NarwfAlEp6Dei7Li+BcJBX7My1Y5pdx6g945DStk
OowrDOFDyu9yLE4uq1SvlSNrtm2IOwS5awQUYR0gjt/GymTpOTyuTFTwSX1aEbIUah+FMK2hQm46
1ZFftmCpUWd/hXkHWL0jWPjHtYPd+BuZ31R+PqVySs+9/LRh6pI8yRrhkVWuEwHLI2hRZJziCWnw
wd1/LE6qiKHDOqSSpucTZJsm67GA4uw3V1KjZA3cMQQgvt0jw/pzt+h+gx4lcgcP/pAeE0vS2ge4
F8dk61nTUQltLjdFdumQD3ucNsEt4Ywm5KaJK9a7UHxEcQdprHrAxi/r/8uabjtpd67alYH1wOLQ
Ki9RatI62VS+W8Zhi1vdUQ34WPlaUGRqWQIRAs0SWh5yY3jYTWAfYDVOxiMieM8JO4sST9NEm8m/
m9YDOwgbEvcoywUgcTXpZrCzLJu621giN4xlz7nN2lysRNabj7SvPceClbtFq8rG667XvGfaTzzC
k+oxIiseVnt81SCkeId5qW+mCULfMDl+Pg8gT9/alUWXpTDdR+gEQsHvJLiRjVaVrAHAZvYoh7xi
mJXtyWHXK/38IRjisDgEZfv1Uj+JHPllPEeDRjxvCVXN16QbpMEup8Pf/NxLNBVvWD4RrIDm3OQX
/wBOeBA0WZIklQMdFXLVgPrw0ONp3R1EMaECaa8ZOe1ElwTN0SKhZF0zw5HN1D041cYILmLefgur
XSGs8KWu10J5CNe4XOiCbu0k70wlV5jjUkC1/B+aFQZzYHS/VtCnmc4IF3PdWjGurRDO4l8JpPb4
0jS9a0enh5TnUZ9HhmOdoWWB6BQgMJFmQnJLVqle6x6Irss57C5JaDI6MPNG8Lelf6vrqiuu0qV+
KjkCZUXyY978HT/rrrOJYUFyiU9vDAFUk8vOIG72kwBwHhUBO7QjIp/J/Nup8i231nkVxGF+FkAr
iAuqIqsw5WjFbWz995u2+c13YW+NzUUmjq3zVNIdUNMWw99CqMpc/FblgjJOkHorntuUBHNXouRq
HXLSNcyySTpg65w7YqeoH8BLtXqNRxXqtXaBhQvN2syiyMhVls1b6RNoHdvcggfKJ6W6h5o4EEwT
MIQNBqUPKc5yEadgfbnBND4GLmkTblOZObmXryojEt7rsZc+kQBPYnYdygMxNaDWXKsrP8DzADHr
aFMuSlARoT/GYCJpj3Nxd2N2/OuzFO8NUC570LXh3GVZFMm8Zvud2/LN47XUN865Xww86eh0tv88
9eqz8zxhy6mNJHJZj1+0ytJnaEGJhWehq5jKRevgb4aHQOocm5Nhy9j8y9tFYJpn86qGOozz0ux/
bTogIviwf3e344fYGW3B2aDrKDXSxGaMZ4XDVt8iZbvLwTShquzZmBNEXnxg9wFFYUeCjrwMPp1M
P22K6T1OI72e5jEEO23wJT4wgvZaVe7Kay6ACD0W45KVSlq0i/DH7Ec4y2STMr2nnAbhWkOp55rz
fDlF/62BFGkwcm2qs/aIQrxmFwJbnriBm1RMPj2kzyYviorx4Vnl5p756wXdQ1WABgr5/WNzW96a
VdQL7J3r3776SABL9WUUKq/J6g0V/aWNFE3vBf36DXUwJ67Fu9e1zNLVRBpUJgeKzpU+u67MsmCU
4kIJXahFf2ytce+F4u71tzIlU1O6tSr1UVk97XvnnmD74b/1vnRr7/ao0LA4qVLBucwLSq/Fwg/5
yTYx0iK6XRgKu8737XQGB52VSep1ZM8tUUc/Bwj+KxSJEeFJJYe5Z8Kc9Kls780R/XrUEHovuxDy
ZEW8mJXLOkJFmJ9FOpd8432qajqdoiyL3dod+TtDo5XGysgabEfzQen1znyOEbF7qWDcschLymMB
rkmGfDniyXjG8oTB/3TSo0NIfZC2tm08WQi/hBQXwmmsQflXhpz4AR/TK0XsYy26DTbemdjEJIXv
XNCCtMdd7K85O+BMxBqdTPulPdTrvffy1ohXo9nQfb/DUbCEaxOJr4YlWgFEMWy9a6Jt6cZG5LZM
/CR4UzMhoSuUlMs50YtOb33Xz12WrrfUeyIGAuGVL2cHcybclzN9YholAk3B5xbyoioV5OD2FlRX
Yk4zJd+QIzglHQvjF3p7B/d5XDbofM23j8Ptfmb98Go+YW/5QVCSlutp7uEJCj/R1n8DCYMj/xI/
+ObH3Q/ZoxGeBrqlUR6y5Fv0PRLgJWY2j61IWSJ7/wiNdkv9CNQx5RB7TtYur6IC9B83ywjXSZw8
aLkcC0jPbSOFYXo7+UoXKfOFjJiN2g7M0DlCevuRl640YrLQgFpPFKyXAr24ctRKBbonlqNZJcsv
5xz48DlZeydnYHy9e/nP+b4R14wgHOpPU3s1lJWw4MI6iZwhsk5WfvYy5AESoaMoVTQy+/hLd+97
lPLf3WBf4vVPgd9vDsSjuFDv2wYh9kaUR14TViyjkk4QfdYru425oGHSUFnmghKwyYWPu10HmL/O
iUPgBxozA34AEamDMXoYq+C7kpNAa9X1of85m9H5e3Bq5VpRoi+OxhwGgsGb5HgAMmZgYg0ZY08H
BKG7LCI8HXanqlEodXNf+iM7IHJX2wVe4n5CQ3SZTUJF2nKHE6d0RMMZ1T4q+L4jTmGAnmVJ6YKI
CEPKZkWCPDmgo9BJ5xR7ZClLfi4/jegVJxNWKGHC8iedsJfiJWCmzI+Tw7lFDm4hK7tg6PO/6L4/
CG9X3ZsTwAIKM1VSXAz7I3TpWxrd4MTsfMr4dWvDQNmVVcl0cHuWtvlCd60i2yWzIs8lSCi9m8eW
G9MHrjxrAXJWpl7E3gX8q3y+Za0+ciu+cm7ClvVyQ9SRmez3HrWNWb18nBQOhKYUiYOKq9yAGu8I
I4JhNCtACAntzCK9rqdVQA7Goxp9kf695XPi1UnUwVRT4fTp6eiM96PCEwVBdNHY9VKBsRNd+EbX
Ux/PEOieRhQAhQhzcPksbDQ6snn3WLWM1ZpkicktnoQ8dypzwzW1tPXPkgyvasDhbEOYzceRIUj5
84L1BHaDhqRAIig4o7c353vUg+BGe++tobyzEm+xdzskzhWJ8NRyF222EnS5eV3DiS5xC0SEkY1/
dSH2N8GDn4tDuQwnMjs0mFa8PSuVu+18Rg/K2DP+C04C5dpS9EbUg6Kdpe+OI5JUCor+2ePo9ZW0
e337P/Xf1zsHJQezZwQX2Xik6zzLgDmj5nLIT6gh9+gz5B3bYBJEJHflFYAqadYSngwhqFy2Eg0P
LMb/PPpLIqbWuPpouemTNPNdd81by3kwNsBcHf0Zx6jONKZ1MD1J9J5vVf1Dvw/jEstjO3yQumtv
MO+8+lO2pqn9q2tE33RfjCkx+n+eE9Zqt6cd2IBt2YEpH28rZKYNIWa/WSjsHPwgrcJNrWzcUx37
dXqi9qZB3KTorCvK5umcYaJNnE50eMPbk/gRrPMGBknLGYy5lYSl8n/p5XLvnL2kbh3rwRa+JrwF
fhuWlQWG+MzJrZ/4/RvFaVOYloOTDhlvG+8bntu0AvH45icrNXGj8SDpd7uz+uUpA2Lk6bf71+IF
Tlh5AO6rDMqHCpjJIq8uNyhqSUw/HpMWaFWl03RkXXOMKPqqG7P4lSrS8m2s7mKTd/qxjOkVxvjx
7J2DtCTqoTCtU41n19c3NQXRLJ3S8i4f0S+L1WXzEFZp78JKCEliLiouzhYGJhsEdHvwS8/pcLwB
QiPiRKwYGQc8+NdHFdeRl5ijl7G940IhnopeT4AeJbvZFrajgq5C7wzWWQP4rGea2GP+STY7CDlI
H6vBj1V7Imdfh95f65AQ7QDrHvV4BccbMrs97pWfNpQBWPq/u0qdomfviIEq01qfwoIoe/Wl7JmQ
2DWWfHAvOLIbbja57qvwToLqeH16fWCsqbOOLVQI3U2sbQkxIMV/NCTpFbLVRmz3047KFX9mZmIF
/vTDjLs6IPPpJlg3JfJAJ0hw4asYivg/EK+vverwDbEvVNwfs323Ce5W/HZ91DF01VXmjb/I82Ga
zsh/yJ5XYKz3y1kI8ioV03ysY/jTawNpnkKpK0St/rrDiM8deD8N+YEbScSNgjouo7fTJmjzaiKX
sUZts6u412r4oRGrOf2ig+dnt1h1TeDp4EcSKwQXcrUnYe6E1tx5ebbIBfHQrw549u2alU7Dts6w
zCBbKv/LBSh5HeI9Sd4F9s30oRRYkENR0Axwtd94n6dkx9up/TD8/aYcCSQ//dMxUR7CrF4KbWxN
j3zKJOXMOoUTl5rIREhQ1oshbPSoC1OcmNEe6Evp3Wd0nTtBkM7L1rdJ5ftNUpyaHqvC0gARwOOY
AuFAzNYW3OsT4xfNXgx0M8t0xe5nc6hEI1YdgUPgEw9UrQEZm/cs3pBYqrJw7lzFPBAnn4ApOOFy
MsBBw+l5L2dGvEAPCQi1cbQhtGNUsU58NOUaZBMr1dfsGw9viY9SWa+4YWkpTPKxj2EAHKEvZaxg
e41gig1vJkA3uqU6zMszJIBfZ/7dsjT502hhcE35ZiXeHnrDFrgf2a4Nfp4KDuoioEA4Gy1NIEhT
g49H5e+OvpGY5NFx+mRFOqGbnxxws5CEAtfrsTQipawrFcQ99bnqYEXHjonjuL4OrW872jJakmGn
ZIZKRlLBuvrQUqIhS6WLKaKeiSY3884aiGzox6ncOyqVVCz0Ej5BsanSdxlbpamC07W1LoZopK66
wejeKTw49BZE2yBuoRV4xcGzgrwmqcwa0wO+KZUduE1PKZrIltvgogqvYj+19iLHAY7x2cBjFTP5
LATMKTpnVR0WINdikH4zveIdnz96R0RoVZhXTxnsLCu1t66kfavrHPmjDPLiqjdNNtLmXBZ0ag3Z
1O5JXk/ZKu0WDTWKzK+VUt3Sx9lGSELUAmOFAzuNrIeY+xOHT0Xqeb/+v9YMpjmWWDR/yKOFECBT
1c3tTifHPrpQysvNad6gZxi9FMjavuuGY/fbF8O9zE1dW/Hv5+vlncCvnZfvDccZjMJNbAKi9vyM
/t/MzY8EWaH9EvjH6l3nKlhktEg1+pjAHwwnH5rvoO7Z/CitV9yC7wgag9BoVHo9VWIIjgcaAbgy
yYD5ZuaAKmW1eDBc4wj1rIm1QGaPHAAIoSEAqBo3yayLsl6Dx2Iy/+XKFG+/k/W5ii7wYKiMRIKi
DkqFgK++jZ9ZmKETsnQWQIM3xqP9YT8DDvDPDV4PPRUpn0gApuuHm1EqrRc/M4mxzRPxMf5D7oPB
wQwvDzwGJmnBMUtSu0pRbREL6qsJImOVv+cqozbN3GrCzDolI9cONmkyqpXxmdwgwIX4y5WOD7ow
RnUaKmmdBtn6aGUBeyPpmi+paJOIl02GRfQWumOY5VekrVhTZJVZt+a6/44UGUv38jHKZG7iMcJw
wicjciNGNAfQLx4SExYlC1ebdBD5seX5ApAhdEcdmWTOlLVStmMkZ/pPa6Ex31hfe/iPKFvWJNtK
PxysWjQKfK/Wwh+3+OV321w5/HSFqlXKd1aPuQ5Z61yi/XKh+u9I2pnf0MP9fOtLq+tO1A6l28zZ
8vb0XvI1pI3q3LeiUvINa9d55AHnIICJv6g+KRm3Ra6Cbt+L0wZM8cEZim5rD8+lIDuRi4oQu98/
IIdsaazDuj5mUrkcxb70rIZNKGxi/ni1mQPkQjEot9x7f739pCdNwg+OYe8ZTuJihYWy0dm9YwiB
/YpwUc3jYdzKzyrnlEQqf7C8+9PYc6+JWNTbd+BuR5wLnbyn/PtnpNWTgcx8X9Sapm+MHrkzSvLh
7ZEUJJKlLd1s97Cx7BrVL7ViiE5cPoRW/Ur1cpaWtl+JoZsS0pei2uEqZnwzFew/aU3qrDnIHE9/
Q/MljSK68YLhBE8Bmkx1cA63apYfSjYYFj2nCyv+XYkumPxr/bVVUdCZATuBreQkV+o8Zf4KrSDZ
CGMTA3VlLoO5asZL1Pb4oD4sOrDIv9z03h6iVEDotmJ4+7ob2MfyxFeSgwglt38ra8FuM3kyMLpo
DdwxA2FY132LJT4Rsw78OAu72kcd3T/MaAa8huSv0pjObX1MpsqYzmBk7NCQE2/MgBwjLmzInyzQ
PvZFJXN1W81hPqeActXzrsqY5fH5o6zB0o5N1+EFCJHhM8xmniFAm4zTxxRljzcgNZlftsEwF4Ff
812cVnh05KQY6Cw9089YcdrcFvSaaZdiAMJCkigToq+uiSGPQUaS8SuOdF6JulSbO/8yygLCemlQ
uXI2TpQ3PHdKgX7RxEx6TCKAxYDLBP5HV/lRfenuAyAqj05VKjAtw44b8hftVLS/SfG/Rwt7DeeD
Bzm2phqG928vwxGVG+WEw1CuPY59dHc2dFHjDFvwkmUZUFsd115sqfbTbZjhbgz7KeqFATvrb4a1
LWzdvx1N8TKYcDwHo/ctDdm2LfEcMfnpqbR+cZN+nq2Yz2YSi9e1MTj7PvsL7tRzDHevnqoVesGl
KdQBdLI7f5RaH5U2QIorKF8VfIwPHJfCczHlCjCk+5dRMi6Hf2ywb2xI9yOlSUbGT4YQHOKJGwGZ
FXv8IakpEnXoHAJMshoSDgR14ILOylzGm3CwS1QcBcDT/OFsC9dqBLjB6ApRefDGheoGczPM++oH
QOHakTB4c7wI1m53toa770N01/HCrlQYg5vC53V9sQCHaN7AXHlhH2f1Fad0m/qnYd7oKh9E3RwH
ZHArzTf3LX7XwnPYw/v9OYlOK6F/VWIPBQH1cBkSg+if097jRkwfOu7baHaCAiE+rlCdwKGrbR9w
vnyiXXBYr2XRHtPcCsQLOu7lzF7WnzFMR9XCXJejHZZbe33KNa73plHTMiwxOOCwGlzS/q1pSxet
8AgIkDTHUqABariMRiLNsXwZNFGd76Hpi0PzRykDDyZt4Bd3DzPN+ZPCDS5RYP1vto2RTyCdTZsR
LDa8SEhhB3IeuZ/ZiRBW/7zuPbiuP7KUxlD+eJappmD0IxwatmdnReMYokasgqLQZlHrN0YfZ5Af
x3bv4inRvym0WAOWmaie+PgJxRfKOUjiXLR7O78K17rVdXq1AkV8fYcq13bAefYAT/D5neS0+ZY3
BhsKzupJuXNP7bZyet43OiGrQzMBxhH5Qktou8bL/LsTd+cKdTlc74eupbCdDh6//2g0zhdvz1FH
5kw5R5OraIG5NWr5m6TReYMViAEWpg==
`pragma protect end_protected
