// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
N06eVVOXgRJ3LPHsYYk1z6oujPLwRGXNGaC0BlDAaI3xX21MVVFka7rTb4xtVTr4
72rM6ncw51WY/lyZ0hTnWUyLvFZmuuUndDzSt4smwrUOOS0LcvSxxIS97BwKnulu
ViqfERkh1WQZ4sJUzneXx/HQsZiFqnSNr4tRV7Dnnuw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29040)
Vg0oTD1CCSSArUl2+9elU7Ar8Z+fVZSmCP+X7V85OJkKvze6l3inV03zK063lVFB
WuQYV3NEv/ptheFbFvWPkp4C0Y1SDeUjFuM+SB4FWIrqknvuGBCX4X5e+eEcOrmx
CAjJdD/gT+l/KI5DIRdTmyWO+nAKg164v7d7hmVI912MrhYL39JHJyJN8Wp9OwZY
bTzGKpA971jMIm7JHRsLcSZYggT6ybu7aklFr7ekLt3K+pQC/5hzSUzrdrEiydqg
T23pXDwycK+m2RPTOGaqpjpK/Ex8G0lRvxOZlcdhmtYkhlUaH39K2Qn3Q5PEQLhN
0wp+0PPEKLlwQvrUVQ6KLYntHsBQHw6EOGjE1MyPQMOWu3e09Pmqb4rnkS75cuFP
iB2B7cc/7nzpdxuFZ6U/tJnhUL31NiMuDUJi8/ZPJlCj2eKK+yrpFtZ2nxMF0sSo
aRJburIw5Pc7O71gl/R3JOLEu+IPrYCclXK5iDKssF7dUxdspG86xSZLhkxbeocG
fHcPQAqGWTXe7yExbEkqH+WlJn2zvkPtn1rohEH+OjcFu2YxY+b4P8Melcoaa1ZL
jSIx93laBNA4LDWyfIxzMKGQPjLi3kXRmlTt+csVQUJojCU3gKAwG/YGAq5ITmLv
Qfm8GBdAHtKllMPXtXzsOdBIUxOvbxlMMA7k982PG9khI2jg4GcAE9LkDER9b7Zk
9ghqnmiAek2YK1taCzmwgkqXq4Mm0KK7xWunozz6G2uAOoya7jezH7qkxrUXPt8m
QbihIa7wCxmJ8WEFP4bRkj2vqzl3VOLu/ogB5ajzDBJHgbAlMPbeWhmZW3DbTa1g
KcdxEKi+/clA0fDpRKcFhbqGNVlxycU21qfl8e0KGUGEfNUxZZiRcNvHNFNKchfp
UzZNLwO53gxNYt5JjKr6ux/4AXOMFezu2/KimX79zf1oXp5WPlp3MKbVTLygWT17
21/Kr/mAXKIE+RSjdJyUTKTDWIEvUp/OOrivet6ya0GX8d8kzqCEJOn6MNHqFWAE
L8I7Z4iiJSfxq30QgcGLOj7HCbyLMegGvYOTV8J2cRSJaFp+d9u0rH+Ch04YJ0/b
sDwY2KwgfNszCnWWQ1aHSFNaHvowYD3K/fErkcN/zQGp1iG5Ng/9+NnSjBq7kjHI
gVDsTpjBwvpmXHbF3JUHAU2aZ7xpLEVOZ55X/Lx5oRDqkh30VPe+WYGJxliTcdoZ
R/GFGPyx0ZfqshvJYy6xUkFn1r4oLEl8tPxpQy+UrRk4wugxNnipWFR00pPafz6n
NH0GpcuoSLdGPk7c2gDQRE9mWUSKgiR3VUW9j4+8lUbWsU9yqMHekFrwqPQrehe7
WjENLUZUcu06NzwIk+GV8yXBeYLrBog1xA3/iQNHyFhzcNQm2bQwGxUk1Oc1TtWW
oxcNPaeH1Z4tAzUBy9NAvK6U5nzLUIwDyCafikSSSk6lX8A1iCwpv+gmTgEND0CF
vflJZ++8p0KBEyYFFFQhoN5bRBhbU6+/UMzGLbVJXVX5ZZ8NcFlGJpR3DYwMAZYV
O4c0eNpf/cw0KPqEx5wT0u8y7yhhmiAa9d0Fz9OjV3x+aw0oWHatakpGXugAitEW
Uf/xuy74lq8gbP+/+sNxbgInbqNZOsTBEIm0a2y6ENV2PiIc50u7iBBzakAAW6QN
JFxnMPNTDReYkEewioXmZAsKeeYpq867XyLaNwvXiWlbKgSR+3cZysSO2/f+mrCE
UfXDOkdfhnFu9R7Zr2wqOIIzNwJMfmqtE5MtXpyZUR4yZhdzCrFy4RHdjPXWfkEC
Wm5SrmAEXBPgQQG44qy8dtQ7iqxWXUYD5WG32EpYqihenLEmn/TJmL9UCjVhgcwU
y8vKshPzZt9kMCry1W5aXJpgaVEBpiZxQbCKSvNvb1SN57s2KMEJXAv1HeTa0MSg
yMddV66s5qfEMau4cPA+ZApZXb4KU1qWVDBf5YnB3IeYW0gp5ZZTlRZd63/ov6l2
oWMtvaYtkjNkObXOw95tZ2zh0fDRgcMo88+D0YwRsR5HFqrBjlr7sAV0O7QWJcP9
k2j4SyNTxoVUscJCDqQm9moZdscfEOWq4HzIitsDbh6FecYQAH9M8ZhbK9vFAFXL
l9hnimIeOYZQBCuwPo6ZQYHIrbX4S02AgCRgWbbD6zfVgeDnZbCbfayZlfYfE1hw
t3djmiHwLcLOx38x9Hw8bMhBkTidAUS7QlwqAwzPypP7gcsJWohCAEMHydhnJhJF
KMeBkgI5JM2cS7RvrWQqss24qFrJmXjvX4cs1U7fsFO82gj+WGDCZvnwsPjK+M24
Scr6oTmEQmek31Wx1nuWUqBRBW+sYXFJbc08+EVxWNcHSCTU9HXoaiDlXY41rhym
krMqk/Y7yrC9oDXysolnZQziXgms+IiQ34uqwAvN+1P6HjtgVe0y8MxpLWS9/tTd
SGxNVEpgdVj4NrfoV9yA/4tcGiied1L/OJzIZlQfCfrD8cSG0bpmLFsmhtrgaK8k
pY8No5vShYfNU12qwW7kZ1sbR+5OQzRCRjGt2iQ7v52mwpxtqfbhxxiz/L23c6hm
RKeFah3E+2DUK0s3VXG+rOEWfojZZ1qXXFc7kvqKMejVZTJVcPiaXboDeDbJXAYa
Oy5xx6euPwk8+NQTKtCMntc8ycoDnkXBaOQw3Twm8y8fsK59gvMEdfb5B8j8YedN
3mbaseVQohCeZ2s0UnYPkmDSS5tAGOBxXOGLNYYsOV+T693mTcvaSyWqPXIUExkq
wXBabSl6phfsGi2PkCTwVeqymZ3qwT7EawhKdD+Qedi3dNjYP3akPujA5shXMdWK
I9VHgUisCeH9RCghkh2ZvpHUSzAfXIguxlDYrnxAFeSWq4dorpfXFR7W5YvCLwGx
Hmx7C00sX8eieGRyoxpyUtLHC2cMm+HWwGDePYACZUrku5ausGjxAPWEnLXPUmZV
oOW1Ef67YoZ6ZCsO14l95pSZbw1FIiylFpLggRQRy0rwFQC52Siy1JYk32AobvmY
pkCQU+2VtrlDek/UbDLbskho2g5ja8PSBvFFfOF0C/GBhkeF+yeKT1Ki0Z21sfZN
IOO9iFE2IbFltBWyXSP9XPv/awPk5o2voGzlO2TL6gdMZvD9psHN3Un9XkXk7GSt
A9JD3LsCmEeg1UbXRAuuGuKL6FtZQ6MEcxMnvF+w0OolnmxzViQ7P/tfn08z/B78
+76cqPJC83wXXbhRO1WnPPI4QO1EdRFfV3Rw+jouBdPX0jPX1Sx+AfLdUvrRDx7v
+kvZcBU4T01cWFLWdeKhy7Ic+PfDkTo+ElH0ON2cNzg0j4SxmUfrA58BDtfahThd
vDxRbFWTuKbdI+m5tmImG9qn+fN8RIXftW+MLAeDHlpTBJimBpA8DzBHHuYWm92O
ruQDKEW4e2E/+KP8qq99yw1ZETwH1pxMMtUHPfCqoMoAh65gn394RjZN8DLanMid
jiqYw2gXWE1LIpg+v8C/h0AG6Se7s188pVIv9lAu39jK2mPZtuuP+jq5yFnRKLNb
2RhigC8gbBDpWCxiaop8as8wWGhx1YTyxeCH2QxD1fS1Q0DYhweC7id7N3WM4eu2
KyghHreQzCT8DMtnVp7xyqsyKBpXL3SG8BE/KIByiDSNIvEwy8RX1NkjKw0gKL1Y
2Q/2pTiqvfv+Yn6egGb3yHpmYkWxZw7QrbhHjVWTGx8qQ3E4YtUMTmbV8d/REssP
1SHSS6ROl/mAhlkVDRYh6af+b/mzSB78mlZo4K62UF6MIcKoRaSmYMNmhwpnYvfx
W0ehAtgungMUX9TTcjN+TnFv6y4D+J9A1n+NLRxGP/wiotK00RsOyagk8Xjkb0wg
1HIlGSTLg9K9hiV5z0+cJwg/1LxKm/YX6/8eFxw8FTShbYDjUbSyF3bg3qOPkWaI
1Nm6PlVlsqauiQS6J3WucOY+ZwMNpvE1rb0tLBV92N5ESew10jnuUEVHsLRapjgh
Os/RUQOAiZyFZMAj7wT1XkAyyHNpsW11CqI6htjyyYVrd4otFRGDRLCI6AAiU25d
lqsWEvT1NlyNii7oxVhCEy+fxCZ7TKYjPha35QSY0J48EDRfnVttoT2Rge46SAqJ
NIwN9pvHntEtv4JHzbxuekU0scJKH7lHFEFbVZGhcgRB39fb5RfVd3MhihBP/TcZ
Wbnx1D3PYmBS4qDBRY2VOnpyBCqeEJLtFRd5W+zXam+vPu5fkUjq0TNVR8Kh3sUR
zeAEJlLilBvbkVF4wur4L+Fz3F4y9OqiU+VZBE1JUck18MNcFm6BRevnUeHm8hMu
FCKBlDQdkKrxqpnb0VHu1iw1YHk98osVIiZGJFF681jikc+Mp3vK5utCKBxgOvAp
J80JvVU4yX8ikGGjjcfDxkS9IpujUTAKpRv+SXZ85G/0ie5ktTmOuxoKLcaDdKTY
q+BLI2oeryKPvWO/ZXCsKUP+bKAuM9znJPSrtq7Y64t4Z+s45E4fdR0590xlvBqA
BWk8ekYqNM1b5GO4UqG4o49fY7rb5lttSSYKJlV1HjZ/xdcM7x734FkGgxHNB9VD
D+//qiSFRCWgL6/13LDSNttTd/VmTzR7rKVZ6tnNs3fyXNUj+0LEFJIhsY4eCcII
ZiZRaKf05nd+zE+73ZasQkWIFWupNgY+BdZZFg7u5Tab7H18dLDg69oIjZk9HD9a
ep5cCNVrIA0ZDfwiipOYoEBb/dGaknnGmlODQcXJjgodOYxYY2p2SoWBO93KeuaG
xfRrhRfBLWUpRp+A1prBlQHu1d5hXtbEHV1FZ0KEihtTrgbBreQ/jvYKvHu3hUCI
7OJy8QTDoZ9WZ3pM20yjblzYQWosevkgW/VxT30N2qzG/zBiD0YLmNYEBQ69cUzT
OQGi8/4NDj+7sxe/gQscfuEJvucUSKWJIr3Eor2nWo80kDkq2u4RGvXMb9luRsZC
9JhuE44BDdwM42+WIHJNtQgF/M7AEfxOe7NyDLpN1P/a3h8MW+0UCBK3dUvdxs4p
P2VpqCDiJ/xksWk76kc27DEiX/+uYCI7ezFKb+/p0hc4UJZ6O2eYZvhghp2AmbIP
NaOT5jz0X8hhCIgN+8CEAZrIvDzHtQ9T3WmbQbffs0HceV3i6umTxllbXANfZpDh
SKXZy6y085tX9LOvoNdYUJcr5x3T7KoKsA2sjDcHbJUpLC/21pCmnMJjPAXqdkSU
yxk3kOopyXvxOEa3/rqMSHVRlxKdnuyTPs+91WC29DDy783pCopyr1J95R9iGsob
O5eSwC/XDAA399eMrM/1e1Txa/D8Ik4FDaoPt+3E3ygcWB+z0UdVY1JQD8VwvRfF
1M3B/6YSWc8tMkR0UISckmcjza22Jf2/SPPbBKXbfHuc3KaVj3KutRTLC1r1YUPe
8gSWesi2zemmMDepv/lbAg/CPu3MTStLWoRPaFaZe1C1CxZQsyTzL8HSW550trc/
l1ragqb+1JOxNv/ve81B29wj8BgL0GEyebLeeIrIcJCfhC4RLxRQWld90m9GU1Yu
jskB6dyTgL3S6XaZZY2A4zCFn98Csz+NN8qKzptw+VeMWuDtJpAOJ4E+06I4/6Nj
WiLTOb12VZigx0/dT3Ha/2h5emT6U32Wl6FIjpRLMkO2/QVSlrhZvISKBmDhh9Wf
mehechTdDWIM2NVjvP1f2Zttxp+6DMUCL2Oq434RY86wYlSbWw6jqPPwDixrDW6y
12qTpSD0u+2l0PPHP68ZAm8YXqjhoohIzn7P/V9TD/nqvzWDMz04YRrybRaJQBhC
5N1Nz129UORHuL8Em8Leo7TIumewlqOOfzU8tcXRzJ58RNSGMLIKRSQqbGDE2YzH
jc0YswmyVQybi6bXTyFvEejOD/Z1BJRQSGGh3HSDBxpd/eLV+tL/CCoPjV8xeZXp
tCxTyTQLCpS0yE9NRh5HF3HDLrNcdTtys4nJDzafvDMgeYZLY412+z8pIwIR4mPx
66Tpc7xmwUvyJ6iArBvko0cZiDTNZYhI4PRzSloKsWnf+yUXt3JvkHUnW1s9vSrK
oWybiE43yqvTe0ifXWnjAJb/iuqclHMAr7z8bbJrfoX2vqsfL0DCDyNw8nBSvMI/
OMKzI0WxJdRVP121DJRECIt4ut8UNolFuoEMX8a5NaH0rgwnQ8Ga+Xl+SVNQVnBh
Z9JMFpzAnN/UjoHVlZV8Taxs6baId4o8FwfjIqeYluoyuBZU4LlswaB5Exxdcea0
gjd5K78PvwVFB7BQ24OTIlfNHfndFR2YAr6UZ04LgljGMzOUb/FZRf3vzL8+bBkX
NddoW8BUivhJhJd63K5hMGDwnMyl8vBXta2K5MHjzZwy3PCxvObv20XwulWqHRWL
VsLWfnCmTPK+6ifFKLvWl87gBVZgODEYktTpcGMLfguoxa/uLEY5qD/sK3jgH9KP
FikV9pIM7pg3V+FK8NgNbYUsEKNoyOjumiXGvpeq0wrgm7xl9iwg+V1u4Wo0y7Ke
ZKsc8AGqDU8asMr6P8aqc7XsxtjDlMgDB14jDPKfkp/V9FC5woxxjHjNAH4jcCSP
hp5nQG7QreQ4wqGSw1+UpwzAL2hKQEL95FxcJGlWdbS20cW1laVFiGynAzMd77l2
sak+8bqUjBPOWqHsSiKzA25NK01xPe4iUQXXQqNxcI8MdSLUSyanx/7HkJbBquwU
hkqQmkKdjGZRmMhcBB1aPg47xTCaqbW8rtWH5E58smnUa8dfVatEZoy5yH3ljzIK
n8DJlfD0yCry6y7kgmwNHLh0vuGxAZclN7KYr01KnEeI9wfbG3K1Hy0+J9Myppbo
GaBcHyqxa1xaSKvVYvW0U1BoWVl4KIgP3D12x4LBw/1E0AWKvXyJAre7uS+s3/dK
1hDBsSweF/x61Hllk5O0A6WImAOCxeLl1dPKRkYu66nJjp79lcn/Gn+Zui43q8t3
TM/x/gSeeJUuyqo+/TkENR/BDiVyqaoLE23fcmSdgCqge5eqz5bfpftcQimzJpxd
lzwsehxTdbLmm3QsqXqqFVFIrZ1CoT1hwscw9FcGKdr7/wn50nI/0iUNriWmlrS2
VmdaGA5SJvyjchQLrVGh3ZeRWgZWuSTXsYEsTYjPpjooesKztw1ibfIZlceInyy5
U4v0mDUvU8+neFh5whkN2+l6P6m5ZoLaufkFA+n3WxDh6umLCzBadrJ7WZDX+Xbf
0BXqrIW0FXI7HgEoTewu5ke4rIivXjXzt6m31zqRFbuE5docuHyTkfP5VgbSiJO+
FCnU339fsAh57s4iXDMJBy/LpZmvSeO/mJVg3loVwJ4jB50h4UNw0NPl5rrxV/06
9vqkZNXoGpNxkgo9zghCPXA33Tnt6B5loBiU0a5jGhISlVPD+EEjUca+7Z2SY768
tfm2+p7KIqUphSeAdO4CUc7JjFYqm4k+XB3G/UrXxEqg1W7FQdsfUpnf5DQt3Hnw
2APu+jva8SiczJ5kCV95GUu4XPhnI8yIPOEF6HC8J/CJa90YgPKvak/8xGxseBFi
QK6kAweWnzBTXXlvjol5rEk537SY8Ny1lobzSzVklHrCJZ17kzNRmIfBi2GqDh1u
Tm8I66y581Ylywr9KW3LM34W+FnBkTQDzcgCM6linjjPACHE5ISO2iJV6zN3Wh5A
B9lfR8TZsKMdv+1FOgADhe2kDrfzLjTwRYRb/TRlAwZlEKDOom7J4FDaQL8Lakdr
gY5TE2VmFH6gtMXIDGzeYfrEU0k3huCl91Rr5//nn6RyUsZLVgBVLG71VXlkxdat
N21VWwIRREZmxFWtvnvCDdHPBzXTWrurfYSWrjzHZNB9Yddfr5zHqppGwsrEeyNb
JPW9zBG0QQB3pfj5cfPMI7XB6lfvjgJWqApdVA3QDoCLSKL5IUWhrRIbCS/ikPoA
rirsDq1lG77H7TwQ8Ba7d8m9MfD7MktL2jn4tcAGkPggbfvqcH+xgkeTFEgqjoup
IUJfNAQM6nE3sTYmNgRh/RhDgg+KbTKI4Brde+5O7nId80Qg/M3ZqJZqDH9YNKUx
4WkDMcTDq6IEU/lMUCI94ZOoNy5sjJH7wvMhiuyGNzHDKpHbkRlosY/2J32VBtzJ
N06Ze0N/0BzH+6tPt6rbvuqo708eo2DpKTdMtIZrwH1f5Tofj3u41F6ino8xVKP3
MppBd8WOA0vsGv5r+cf+TdFLca7Tp9KKppYOCxSqwkVoQ6lVZYKPKYeDPHVRYfmx
Hm1kfVzaEPIl6/PnJHoopCwLh88Ezq19LOvv54lC78X5pNEdufq695Tq2vorG0WU
3+2WTIXMnRLHcbsXl4398QBAbqecvRAlA/rdDvV+rq9ns3gJWPtsfw1gRXGCdoeK
fNtnH9CqtoUOVhr3GiXvtU0Y/63oHLBOA/I3bh0wE+nrLnSH5csLfY+wWj68VrJJ
VdEEhIffWeiyk6JPdwC4rVt5eGWFy9r8WOjC0/jJ9VV85+LWJza1qB6mS6/QUlsc
bwWR/E35PUgJPwJ9WfZpPD8ya4OTNtd0n4JOOS2XB+WiKX8pzmvsmBDxhLTCASpb
XdrZGYTtiM0IP+A4IWcki70NvXgRdjsfdTbeFPdK/ybxYMrm9LoYoPbz9mUAa5M8
fTXclbVJhmWW506FtC/utfhF6jAu3p/jQycg4QzyPqvr5UVHSgttn06uuplMIq66
OnwOwxRLE4HMYb+h89QPMkKsaF1tiG1Ij+kl0qXUOlxUo7LjXIs6ukRTE66j/qan
Zvhuicvo8RepqGZ0m0uScUjo7fs0S3l1lDA6z3n8b0Bk7Huu3iz8oCK3KPJBYa/Q
Y8nqnDVxav0WjKS5Y5LFyodNqBWeEsZEFLt3tqWisijWveYMrLwKsNuoxqQT8Vgi
UgpdJqdVCx37XN2+cc9c9hUvq0/zoPYVAGL9LyhZpcTGyVyqUExOZFcID+rBaXPl
MQWLIjeyw4ZLXLwzmLKyXOxpMf6jVtclTNash9ZzjzACAZA3VbcNSKbvc4g3abb4
sHMz1x23gg0gB3jouP388omROu+dB2hCNRwXGYS/ziouhEhhtkEKbXx4qqaFyHIc
y8K2Lf6+eOwPx4yciRVt5crgWWB+tHvFhYqCwSm4b3iYnam2SesdCFlXUe26eDPM
YPn07w6FGklxOhxAqIy1bqMNIDW/n78EgHlAvt1yqwzXu78PV7wQzwoNkAPDFcCi
e+DexmKUVv1BXes02JIqvN6BXZFcz9HfDWA1zhG22lRoDo0E9hH3WqCcJR3dzY4Q
YH6YNWmbrCLvtL6JArlNxHradcITrVzlnAEh26iUFW9F6ZE2v6yxEmJiUsVBS/ar
1nOCpZj47jqKk1MZRPaYxGcsNGefy+TPnFVr0lc7vvXQJ0Eizo81aJBQwKkNjqGP
U8oTPMKdaj/GWNXsaWtZEXZ7z1ObjZ1hIXP1ZhiTtLTqMijl6JHHtzKeNB7Ya8pn
OmZOUObKRaA76JUPesu2WpfHz3XLqA/FZya4zQlXJcCv57pE6PHEdH+YKpwGf+nq
nsSugqeixKn7gz0MbeKTSROnI80Vh+S6TYd/ebfb+gksqutd7p7FQdX73hjmpLtE
r57nLmXeuMCttOvxDMeNpckEIsZm21dLMH8YgbL6Zq037nLSDOOb+A9YcP8yBw6b
gypd4kbbD9DAvO1TbXSsgDt6pZdLCNb5VpHSxWhx70UOxgTTJ196MMHz3ZqNGspp
W+48WUW9aoTkF+CjOcogmWW2Iul2g6R+xYLx6+34KikmppyLvfBmUB4z6ZSDsZph
ch9dk8tJIkSSO5WT+ehWyxEo1TDstIPcHOYi5ior3Z1qSgLoKWwhzrmMJ5HEhJi/
uxb4/bd/0ss/kCOMkaoMY/QtvEwal6RmhwCDivdSAalGRcHOehJLWTN4ybX9+VSi
uweH475EWMslQ27uN/ZGxwqEaHjO5eH19aTleoiWQYsyUNdFLVIcMlIUXDGCwV+C
v5i35j/rQ5XT3Fl0lZYxpsuWww2U7qE66Ev7Y4xEWQTmzotQjyqMSjdewaejBGzJ
tLQY8J7p2X7evwp4nWWu8DNZJybKYwrYv+IrBHNyy2IH/nuVKqRY/wNvlEkI63bu
vd6IdLaMPKhXrvJAlqyS8twiPFfmW9hmOQGiP+LD4oJr27LOrSba5fGO8R0SfZqd
9BT+6w3xwmmPA5mvtsCbTbiEPNCaAwngdltnpznq3IewC6FF5tgzzUq4coOAysaj
0xpdJ2bSqS+BP0Td51/JLn96TjaIQYAUrfDJ1JIinbGKUcDrCheXM9SVBIXS75gp
bgfQfHICdA3+ZaKphIxkL3JOiCaXyct5PsiMCG7DEYZFaNYkkxW7E1z7q6xQeKTX
K29g9pGS7icYO6+lx7e3fRuhpIU6c1XhguB9YLwOt9bd47zYcAsoBmqK7BHQivlS
rzHx4OZPIl1KTa//sHkp2z4ZfPDzve/tqv5J8p2vNbIvF77vXAah71Qx7al/NFNl
2/2XzWzUiWuldikwsrinVBd2IOHlkQtNBGbZAWzkXAIkgVUTXNOonIFzM7Pam/kA
OBn2jN2bbJIjqVh1of81bDfJVUiOC/ROL5W7F63c+8LCMSNJPZvfFsUwLUQ1Yle0
derQiDFiRNI9NroO2TMl6ibbIFx0H/E3izltQiIhRW6KSUNjixpzN33u01Z3lf2Z
ZTqWmt+IVqg3g44Wql/0Ngs8OFz5TMcXz//EljGMupscd9fdFdXX6Kp5Zwe8gI7G
wRh+opuPd+or/ig/tB4ZtnBcLzoIKHkNtHqvi7HxRkpycUin7wConCE0tjjnoHne
/caVkFJ1vR2J9UWz/adGCsGQ+pH5MNSE+vjyMCgGN0+BkU/lP/Fwaul0uy0jRsGL
KJ7T5E8ThPjqqOg5PNO243LBWNholhfCKTzNdXxSXf2xaXS1JqHddnp9XsLo4/KM
grnlwfBNgKVGJt7080zumcbkDs+kvhDK8CXD3pzcy/gkyO6F5RbxzkcaurJdEh19
vUlX9uX856yw5fT+vHE+A4XGCYF8b9oScmdDZQshrjJL8Nle9LYAIKAHccHhDMTs
XlCTP90tnp8P2AqbN+XY3NkSNXObpadsaKywc6iPVZ6tTdIhPOAGv2EEsjYJwO2l
/DPeioyDBdMeASiKbHi4pVG7KzoOSyM4LcYbZ25trfkGFWjBNmzTGv+c3rMXgiHI
CbUH55RUPY+/p9ojFZPj7EctI7b7P6Nglv40gjaRLpUBdlr8HF7tFT7s6QG0IKiy
Vsu4jRVlV2K+FYPSRH7IYTqAHkDPtmr+JYLt9L7q3gndM8NUDHgPC3Lf7zcbG+Pi
XFDMi3HnT3HHtzLiugsYHsA+SsnWLY2YB7XJtQvc4Dn4MgUzOtGT7RMj+SSxIfSu
WjGCmi4SqrVtpAJRtr9VQo1+navtD46S0sI0TVZrNAOMdlLwh63TtbZqvtixOoql
hbM+ARG1zFNajQtsz87vQoNjfYevOFjXRxEnJHfWgWBCU1jUMC1T3z63adazNLq4
dKq0iof8uZD0IwNWSVYw9PSlSkw9n9nx5HzGRLwaQ2Fvlbuh7vvOgr9NYKRHf97m
27rsdecEJznbwW3IwAnrQmtg4Hs5EJAirMJ+pW6jCgPYV+ASj5vuuOCm1HnhX/vY
y8EJ+E6qlYpt4pzdQo5S5jmQ47AlO6E2AugWFJTT8PzJYBq6OtJW+oUf2Sc41a0F
FACjbGJcc0nLmvw0K6CbFnlIVS05gZ0PIZqJgVOMUdusB1V3JzawZhh/cYPoIX4f
gGb3y6BpRPU4iLhDn2rl2PZclOXCfXktj4c5BhVH7nZ1ef6r0NiBK56IdRQHrLbz
OTotb0AuZmrovWDcN7P8uWVy0UBC+bEeyb62zcWuOX01vHcNMU/sIDVMXjZBg7UL
9quyjbCBJ84uhugmvNzPFTrjHZDD+IcEDqLP3bFPLFspZa+pQIdbUNRccIYqlHFx
YJPNQo6Dv3le4MkZmb3rIgSql2QAAiCWWeTyFKH8WhnDnoKVVL241qNOXyZe7itt
szmbPLHJ7//u8e9V2K++Jlc0/me49L2tczG8UVLjgluoEumG9fDmuRBQSOdIECSc
wdzHj844jTHAP7957vvYR6VpX+mo2jzgA1J6Uh8MeemI0WcoIJ+8IRvmdfBlP6gY
E0+a8AQFPdrokdS2v7gImmxP9cmr5pYMUjfzYxV1Y5JmOz3cf/H+JdQjfEVuerR1
wyYGbNutLCfLX/1gdXYvxrm8kDgMyfNJX0xcAeQ3DnsiPmmY+ecHD9yKRNHu3sKu
yMM44o15/QX4+XC6JJ46skhurb/rwYZSVT690wuUbRHAvqOlFVUxHzClP2yFUrPl
QA76cY7mUPgkIgGwmnfLczcz+Cw4YQv6SIDnXxKQBxjCgfcHgePvzYij99LV3SNV
kRYtogFwGohiqxQduPMWv/Yc3NsWoGsrr1YmPK0WB5/KmF6P4Tx3FkikM3UkVq6P
gltETFDYsj1wZbdfaDtuNnnLCk7PuWxrYa809lHv4iKa80CB7BLrbs4Q/0d2BeSP
RSX8a/lye10t+oQjuTQTNS4MoYZDaxmQxeANAoa62OdNYp6PNWt+rw1Ujq7UixnF
Vs6igrIbCH3UGw1+fvuORFk2RcQ5DwLaAMmNFoNh5kgWJhotH96ckzQ3b8qysFvM
y4QLCyx9iPBlOHiC+it/HHAL5MHLkl+EquQRw7VsTEkIGarOY9sqJIhcjxOJO1RR
KF9W/0rsj1n/AnQ/L270iUpiT+bgKskv1CySRAb+vttLQvhGElAvE6bNZIMOAyVp
pRhhxcM+clFz7ok/tGvgBhrnxn+oL1vmUDhQI8z8F6QWo/Mz9mcfPuZpsXvgX8ES
YRSF7yCdJ0rRxF7HoicoOK8YcJvrsLkX0AJ9auwO4fB8LqCyQXaofD3yKQPJ0cAs
B7+t7xLdrF4Dzp7GJH59oKQbRynyANQDI4agSZdnyF8+SCQmv0eBq1NkMqiFWY3H
jQ9SIzxDMHcUAPV4gSDZKtoDjjjuOZ9bdpbCDqmHwT6brlTtL0tumr+7LEy/YunG
Ra7x2vCFtcYgtNPx20G6xwzhvBR624NK2kc7YDx8mYfQPX3JEeg9cp2evx+vRzzt
X/Eu3dufUa7UL/41rr5GEMrYMyK6rueHl5Sipb1gEtM3eauztaFXAz7qH2sjjohR
ZnsyenLDXQD68GUJLnyZFO+d7oSALkh3bHgNEF9rSPcFRpJwUnbk8I8EKP7jrPG9
Kf8Mefz7mJalmqwkx+ZHDx9XVb/a5+Clzy0kSkpx2qn41wzIhqvX8MgDHZujgCpd
VhvgW0rl061LcjilpVPGGLeZDUxJ8U5PNATA80QvYo/i//oiQ7qlRcaBi5AOBCrW
rX5cFGwSlTldIOINEbW/i6GpMVN1dEhDZ+bYNJqLfoqa37TJ5T2CHIA4UFlimrn0
OnyMHiJ9oBc+q9dbZUSvXkXubxsPRQYmyLM0TzOkCoVk60Oa4bKehGwa3rq4YQ3j
Mlqk+KQMsUOWsIQIPEbEmbXa+oRqVoHSXGf92+fN81lR7mf4WYynDuce6P3POdec
4l1jqL/RSxetp9+1bwP0tcq1m2YhZHExyb4QpTSQUmIgXHEfVWmdiXWFhEHDOesC
qE2sfzTsp+rYBq9APFquWjZuBVbbVoWGjBBDAPb68febWJf47pqki1Ea/P97ggtm
WoImxM7MazwGIMVR7MTAOKlKV2FKgpJ/66JmJ9ciyVAaH2Vyqbo7IN2NBpwW0OmU
4p+FzB5k79jpM/oBXFZyOWNb4nl9/K12901jQC1nTs6I4qurGE3v2+3O3R0ETpYq
Y6y3P8Bj4olGBXEk/JYa8TIm42MuDEtclmT/3YFn6cSZ1qUehz06zXlR0E8tgWzs
xKcANbV2ukX/RQQsfjtBSIsSscb4BrpsS0X7qazAcprQcZuqj38WVsKOsea/gY6U
mUvXdxUCDiyN1wxTiaN+4oi6kC804ho/dyduozuxquGj6IROx6haOOegn7qqvquI
LQBpiLgpfhbk4g1fpFSJ6dZ5oRIVMaxUaTt8z7zE6/pM9/88AJ6dkDUG6HbLfbLV
N0L2qp5lWhivTyxTuEtJtQXq3DwNZfvSeBWKV9UNmMjfnQt5HHeYHGg8dxGWP3IE
xt1A6Vv4tpM5iffk8bYc29MDk6hRWVYLNWOE4i1XHoQBjCQ2T6++DDLwO15CVcnp
XwT0NHXJr1VvycSLSRBvGhy+JVmB+mrJ9UPN/OXtJZ1DXzWkUaLUPi8ejjcHrBCA
+vSYi9MPjcphXDqa3OUjo2dyihf4Jw/E/n8JFlCJWIa2IV2+g+N33B+vb5YKt8PA
ns2395mwTfLnd1CxYzxvJphX53e6RNwe1iiyZWtKsngHLvpgcw/KifvJPxUrdBor
aBMSM08HgxwzS/OkRWeVnCdzxRW8Ae8njrj3lQgIR1LSHVpkzsUMSC/K+TEetonV
K2v/x/QOQDx6+E1PgAX/eWN2ky78Czr7zKlN72wt4htlSCihC+sC06kzb1enA/Nx
G0F6eMpwu1C4RuVJ+LWV1B/c0LgBUsRZ+dhBX5xvEgSyctkh4FMZOvx+hZx8uHBK
8rgRel8KJEdQrcrlmxbQFwUiLqAd2vvmNIoJ1rDdCb1VleC88Ih9h+UA1B9/7UWw
3Z9JoPkO7+JdcI9cuDwjd/lXwe242MBsovhamxgjRj+0AGWouK9I2iEVp7kgcPPu
fv4ASRzvqCA6XIqTp9rtWw2Mwqy6/EsbbtUCjOeLEZ7cM3AH29XRHSn1Eav5+Xe9
z+HY4Ol1qwQ7uI6PXaqtDU0iUnIA7Dzjq36IVH7jw4mLlzU2gMkvPoqTYjp2FIGc
MlW0sRaimihMQGeeKwMOIwAJxb2+qE1W3tJKsk/PCkMGmMmBKra4W1Bn6JUTf/4D
EhL+1ndojW2aNEbrX3KHlkkCHWBRU2SKVUIT/zjV/wXrRnhSCkk/G/kjCByE6xY7
wEN9WcvwGLc0UVQSee2vFCxX6Sb6Ci5yGhKmqlp1OqoJH7gVF+U5C2O7aGkFMt+U
2qxf9hBdDOJl0VsUQ9S57L2O7WzrDSNiAev45Ptn0zhD7sFYyj5KpG2w24ms7H62
74iWrU1WZqP3KMxPzurU2B/Ey/Pfwpu6PhpJ/L5+2yQopLoay/mjjlpFXzDnkAMA
GTGHJ0S3RbgqHLl0TtbVriD0yRqOGgnT8hoRM2jQYyWeH/M/oXt6EeF07AInmDpJ
BtIW85LWcpN+HVeiwOEHu7pI/6If5RIy1PQVbSilMALiNiDrHiFcPKLBfUIfkA61
SIkte2uNtZfV06fD05Xq0bqLmnDYFvc2moXvZfpCdogqbT42tAXQ6/hO7ajN2k+z
o5wYdfak2E6zxQhAgr7jr3NyPcmb395IcAMuIjFY9pVYlDB43YLi3BhREBzLkbVD
uo9bKhNgoY21ryECH5yiQ8Pi4EMbtJ+34qNXpk48tBO8C/NWKY08TSlGKAClXFVA
3AH2Sfu7KcpQLYiePNsXOJ9hCRdSlioKRHK4QJg4T4qci9Y9OQOyf2spqhmKcjyR
LDgzxiSzzObOnoA/tR6ID4BhfaWWaMZDlXlmE6VypE7UXtTo2KyDWErGMdO04hXR
xBtlc/ochUMfixAeye9khGZgrhuPxz7IE+K8pLTo2qAj+a4Aju4GkEDrX9w7I/oS
QolLrjgddadwWS+5hp7ZT/tSSnYucWSjhuSF9XYq7u8mZzz86KWYgwI2hLODXNRo
nv4r4OwmvWad/wPGJZb0pINCIfmL8H0NdOMF9CBuykXudI9Wq5JpyMrFZzwp671v
BBCiGWBW5W8bHm38ofsCezm/Jnzo/cbptOuFtGF0OENgcm4p+V4g9a0Tu1eR0zEQ
BKhYS74ITRn42AQhJ36QWmvbvQFOted3+IDacsXvmJXUFD7vKNqFPpuIdtS0dDyB
M22yA0FyFKgfaWGdbksVgqm1NGkSoV+OUhLVlgdKfYP3gBpFI4683WOgSYYcswOJ
G+M+M90tXJxdwAM7ZI8L7IQdIXiv1advXJ+U634jpM6b0xY+QD2MAlEGOE+cVG+B
rkq3WrskK2hlVHurmKtm3ue9Bqn0b90J8EITGHLrgy+OznQbp02tl0tVPhLxBBwz
ZXCu66cgPp6tOI+ij1F7GPAn7uG0mFOGt4FLTC0I7eVqxhM8G1QvzycZ3A+99B48
y7LdIe/k4lTT/7clu38ARhMv2AbaZrec8a0zFIfGN9qxyn6vdKjdDtBKSIc5B0dC
9WX/FkmTag3qG6aA4CL8EcWJ0IziBEJuIZbFl3v1nx8Bxmve1yfZ+Li74Wr1OlaJ
tj4joJyqUsTEFdMamfZuUkpIYrKyJQY8pOYxu5PQPrmoBPqSqpdK0bhhTWMwoaK/
3Mi9nEVZrMLzOMDMn7ormH7rrVerMDT4pyEIsaoxzO+CZumjacxqsQlA8PuZbrrt
rzWsWhtAcvvkNmOFVQ2ibu1zC4DxKii9oE0hQoYE2oMHrSYYH9W3xTMjmFxkk9yW
NETEELEigHC3+wDVsKaXDL1h4Z33RD/YivogPGCZtwuyMyksASCb664FEgli8RKl
FWrJ3RitHEZHtKVeRp+lhu23imJIXrjADD5igH9KXg6DHeT5mjzSLEoMQQfedv9l
tgaOO852T9GfJIidGAnJj1wFDNEQDTCCGZG9C6p9wf1RWM+qPn+skRzhRjrpMU7b
UfJs4JO6GEUUci60pgd0oSxSfyc51q8u0l6xv/u7ez/PcIDWjgH/7+l7To4tCqo8
9r1ImypyK6XcWw1GQMZimlBSQA9DJfiZ05GugGfOhCKkY2C7nHWwL9PadUkzkx+f
enX8CpkaPlAOk0l65CyQZXJLbzKwptUzERTPeJgIxF8zBktEU/hHrDQHZL63OlMv
rbQnghgjdA+cesferNcTlNLR7kOCqFbNtynhspyVJdVbtaPvM4WZdjaqAB+nfVyu
EeErjy0doqB16bGT3nnd/vWE9Qff1jjqt0cuwvfZ1su8AUw/JWdphWrldkdNRso2
9UBW4G8sLxZ3PvX7i8Xp3bOfHQWpjCa8nau3hfcEV1HFnj6rNY5JkIM0qKjajvfV
ZmFu3Un9+9z46quQ+2O8Ew9VvpsR0MPI32weYM68bTzD4m9pzeLnWuNH/yAggyhT
LOzweefB/eeVo4+ESBmVVoxe+bZe3wkG4IyeySf319oQBJDU1uxotk+X8DcPazGi
y5L++J6iYNrGoyaLJlh5K670kkGeT1FKyxxk5iaQQO7vhUiX1+H3s5DASGljoG4l
8rSfiE1hiPL9OUunwkCOriNa9QEyhYdj0bduvguFYEMZYfKJrBVUyzKUcyX6lptI
/lUcDs9KIkZyzQBhbJ374rrzuj3bxyZ1k4jP6BYATjX3Ho1NFAWaiGbOj0lkxbs+
CZLw4t7bU2jt7FiLKlt+amjeOjM/v5UmnyTsKBmnvqli9MhuIF7qpqwzqVjPAKZC
rV0zoMcLa3t/+epC9zGndlrz5+Dz/FHRdE6uFrrWZIQE5WFd69KmW0JlGGN3D9Jt
E775IHvUNivzrdhVeBV2CkrGnHR+FlvESpd7CkGPGMqMMcYc3N0j53kuxrmldkZb
jS5ZbjXqJW1uSWvXjdiHX0fdmU1Gi/Q5hPhqIQyfcGRHC5h8XZF0Z/lP5Uc0xRI9
PJlGCKSNHL6x6PltPH1E5RgMMoXlLpMdkhsZ+Lz59ZSYBvkOWKmZmkkjBQFk5Dah
0mUGszH1cSTJ2vOkjFXyZdui4biy68mU7XdZPaYjcF2y9L34iTk3Cu9rJcRHjARq
5Zl5ka9aBlWI160Jjmoo2+ajiC6oTRyXX7SZnaCK8wlQhcZdHEkuV1RDN80wWPIF
WWA5VzdMj1qjk7qv4W+ZUNGn9B03VjZ8IsNPS3cuHTylh5WH7nnUq7/RKBD2r5gN
E4y6B9KZFWXKFIhgfjuBZ55QCromdAdPUBrPriEZZjTzwTj1M8kHnL4ewUnc1MMv
imRugn7AxaSgRlyRsPyWsgSqdyHWGlC95f3oGqiIJHdPuLRLoaBSbhyO+fo2fGhQ
ANso9kbfp7Es+cvOEQvM3reU3hHVSuxolPnZA/8q7HTYQbNy+QGmCuKg9QYuGFUe
qmQZnUAV69hYHII1pcFjjAAidIgc4cJKdkcu1hvQZbv/vhPMBEb7zXGJJkRMnFjS
tK7R6BuOsUqb4vdlF8SDmvKCkUd6adb0F8wCcV0GDo78xQTQZp7YdojNPfqlf0lw
b/9/PlXfC7VVtkGYa7Imv9dHVkgvWHiPmSkbbqXPW/LPdiPmz2hHXSjQoUV+VB2H
Ub6AdruWVVNAebVCLNvx5tZ5J2gwMgIdCxq7umk4wBfSzxVQhH58H6/DXOlc8VWn
BLzw1/9Us3KE5snMEx03uMdfAUxLWvXhNHtOScfUBj3VR3mKyGvlNYJsp924D7oH
niLbEj7Y2ApGX0BDpOFaPkRSOYHMXL7wWMsd/e74PAOy9R5l32aa5BcGb5CnTgzo
6lQKj9V0T/MNyZizsvW3aIvsJwTpK5MQCLCUl1hXjXSJimaSTyOZe4fElN1GCskt
LhV5R3Jit/rywhUEOPEHBGy6cKoh+n4cx6qqUNE7veEm3Q5fClrC7GpEvIg+sZrh
sK00b94y/m2qNlb2no8PCoV6/Tr4um0zs6OMsx9AeHaq3fX3XJsNQfB+ql+xHmp7
o+7xKLKUzyWuPhf5tJYfxi/2E9FUaaT6WfLSPzCtVOgP/sSeQN0zbu1TasBcGn7U
GkNUy+0uvr672TaUWqodOnQ17n4KVHtF6m5EJSo/j7FRYnzMNiSB35kXrKhnGzqb
XuSURO7iSEAePvNXnml43vY9miFhjy4BMQo9J81IZD02oPtmM5Zuy/5TqeYhR9/l
F48fTPD/6xwuBU9+0/CRdQ7mYsFTtTBMJb+3i4gwZF6oA383nuKyGRYE+vlW0GMW
+ZQJdhb2KCWzfLOBK3zlxhNWvHTuh1VaS5GHM5OA3j8OBHH/AxZNBW8pMD/Zap0L
P/db6M7GUacyf1+1x/5LiAmEidwDsIrH3GZ0eDrxteh8JmeNbzIODm5NREc5cqaB
uBfxHG6d1IDfcFW3jcMOUrQFWzdHPenR9JchZUdRgAcap90ab8mz6x3+W8qLFaLi
rvCl6DdmdrvxDDTJ6aClu66xGvjVkEJGxFGPVy4IyTzny9H1I46IJ5RvebK/Awq1
pOBSn6tSvCpz1RRifuyMdttr47Q16g45gCUHknBf4/rsQsBRVHP7wGlqt2bxRFk5
mpNj+TR0Ri5y9+X7suQvm0v7xWI8gstRYziQXCtSnUJhpnTdyMXq8oMHgAEJnJuF
Y9H6OxZ4wAKIh9GcBwtRNY0ESNUrChTBJmyMtFpCiTo93dgwGEpf3/jM6YRBf8GY
MP7cGIA5RPxtuwdryudMaIj7ql4A8gd0DduaZcqDP9yImo08OLfvBz1kPIAee39C
Ghw2v4y1XnafOmDtx/Y9n/DrWzh55aiwH9kdtxtHVHzGDvA8djhbwC8Ni6PyCS9a
JqZ01ItfdXKsRAUyK9AK90tO1cb3usBYUYJYVINHPPYcJXzU7ykf0GG82ehZ/Nlu
gFb8IBPZImOVJ/+LupIJ3JmIo7K8zYmDxvQM+iNyslvxEtkkswSFpIPthqApixB3
4PrI9JBy0PQIqs23v8JeBx8VRtZX1dZo6fv0o/+4UBrCZqNMKV19FbsaWW6mwH8Y
+T5hw13u3GoF1ff0EGzvgpark7k+5ZagHJQDUeLUquY6VVSRyrgubEEFVt84zh93
Iup/PXB6h+erDlGErrz0w+ZxdPAv3kV67C7hQODHY3qD+iHbF2QaU+NOUlNN54Qt
DhzdNfgbOFFIdFyUdy3KjVVvA0lc7a67rJB4MC/hseesiLsIeZNTJsa5piun4djZ
YtnH7+BYgQRrjer/obASXLkA+kiC+8eD0ReNDEgMQN6wGzraKpWQukd3DCM0UUkc
EBDLXdAyug7kH8ZuGYQL4Fhz+7dvEZnRI5DCItoROnr3+l7DHgF2AlQ81gMZjtI5
LBcWWMRElfF3YWTk0qXijoYp7ScPtfADnocUpvh4l45dhnXl8oTWBI6xrEp3t7eb
WYHqFvPg/79hszsPuU54Vao5ZuYlicjyQbElteFZ+CxLZkBUFXWuROzxLbpTmwmP
3k1dMdjaPfK9OqDhuxsmJYaE2GX9iQV0waDgx/BtksMBlU8DvdQ6NQsx4rFJP+p7
6+6HsC1lTiulcIezvMlRikVoWcgpmMFYz/S3KxeFAZuv9L8XgfUGP/u/eABPuyXp
P2Kq6qFqa0YasXgenIpjafL/Pw4JueyeXVjONx3ujYf7Pv3EwyiYjIxPnPetYDck
G47G8y5EFdXyFkrtq9E5kR1QS0J6mkUZ4oRvYQ7IR72jnaJhRKjt9s3aMCEUZaTj
ts0SmTa5g1Uv0lxW1PqU2qN5v77rGoCkStUNmKUfWNU4n8a4CZ6iWRqPKuKoCHWX
D2YFbJshcCfhqevt1VAnqOMb11HO0H9yhJJ7Bu8sEpVeVZfAGWcvaIhSiOW3OUf8
3vrfC1Gf3jBKtmd8wHTuF7ZN0ZikigltP2Sx4e+BWX4/0Ea6eL1si+GIYJToQdBP
ynOahpVz7HOkZ/2nyYv4W2XQeXxYTzDMGT02xIX3PW9rFvftEs22EUV6tt0ArA+1
VKKyQphJwFcogsxM0NN63ri5Am02YptKacn4q0JMreIj4SlCONE0jc32YgNd6doN
dl0teOC/GDi2lX7ZMBet9bWorxHVJIHpJ2SFs4XSjvj4CxE4/r/gdR9xMkNhhqqv
eBkyfqUGXf+zt9CeRfAKlv/sAa7YfRGBJgqjrvgU0EoV+Ys1sRQHrBoZEKVowLJn
Rclg2M7bPQZnCA96+1Fp8ZdtO2qWCY8lvP/9MbLuWJAEgSrFrFp4EKQWnKai6Xs6
2eLkCvmhVAv0QHmXDo1OnsN0tD1iW19n+qJGMmAljdpKcYSt5mS38iYNl5UYSY6z
lGsYr2X2JRMV80OYuVmNSe7HTCKTGzIARZYoZ7V+oT+hjN3KeRy7xyXhkLx58wyp
gwtwG3nCNpqOxxmYzJ1aAFMZajykwWuxxcuHtw1C82DWIul2FB1BdNm30bxMucWy
ORyqGc1pjM3bDzjLv5hEDKrYIiW9tm3UfMB/tStGd2eIStAcUhxYS8EPiBauYFFw
RltVYns4TL+AM6SZkFRFNEP50gW7AJ5g32ksn5xbVjJWfmeaEGwQzytbdB8BU6ti
jGETnW9leR3LMyI0OJb1bh71qr/gxVepUCoNEOd2o/3FEHi+8EArp+GM5cLinu5K
Ww5dg+dbr8Pu7St/MNj1gujyiPFtKPYEfDFH6jRiTpqkNEUo1EGzClrDmkdfRZ/V
CtxJ81L9rqS6yClXw5/4CwNscbilUzrmvtui/meM2x9XR6Z/pZWTC/B2Bxgr1Emn
wzvRfHHEnV6Y0HKjtcnkVLqH3uMOl/IddKmF3ADfwgH+Tb0xZ5+iCMaLsrFqBeBA
Va2xV/DQuUukR/mjTFDuXE3BAP7rFfLQKwJaZWdEkjRscG6RIAwc00wMX2UhrPVG
e/BWu9kXOyIXh+zcsZBGFhEX7Cd+sdUrfRKHKYenXCvCOyaa1fJ2g7ThW1lwugS2
OoRad63FdMI3hWF7GHh7XAjzbbfYi2g/iR6X22ngfSjMmhvsVAV7eCmQ+09EaxYY
2NfTp9NEat9gyUukyOxMWJ7Oi3OJ5nTValC57ucifk0x5nTJZfTrxy2CxH45EGNi
Z/izTVrBzalIDBmIL1xrd1xwL+7koTqINChZ1aYOBGUrL5Frv2PwIzoxYyZ9ymg5
NW+87zaCp4HfXmcQQU+e00o40SXw3hxZo0df0BxV+OS+qIKFYeT8Db84edVnvwho
p6w33h4muwl7zHIiPkHxFO5R1ud9OmhtGkzF9Ymk0cZFprFnPbTGg8o3VBYbwOyQ
GOQPBWRpRLzatSW/vucLFqr31/E4GETU1b9HUj7OTNM6a1qDTZf8q6O4B+sajRE5
SVGzV9DjaNra+RiZXtN8gykfB9e8c4X78pUy4EGKWia+14qUeXrOhTPQF2Y1Vv74
qjcgaee4VoygUWdY9G+TCJZJU52usD0ToXjYSW0HeRLvbU+O8ZHCozE5HSm9baA6
mSleO8jOTR8jvTvQ6v6j9hTHJKACd0YrftC3gn0x8/KwNhmJakY4FX3g887opGjw
2pXfAWGnS5eGSeqE1TJ1c60/GNbi9iesBvMHsLG55ioeKjfqJfyP2o2WFQeT8S8i
cfUhDISWcHgr1BnVjHIhzdlNPilqIDZS6Z5RNzgMWnwNuhNhlnjCLoJRRqZgbBzO
0izh+YOuiRkqtf4SgFAu3/ftopIg5ErBNGxmB3G4k3v8FjA3RmJyeX9nKvSe4xjH
quhCeIP2XY3DioI/FbMCpifrlpDxseeWGmV4goqCHk+4Y+eZJ4ozeMhT7aXxjTEn
SoeZ42lE8PnMJXDLel1cKx/HBoiBMSqpnyY+hoPzBMEepriV2btl6Y+Sh7c5o06e
6p0oGylDpbK7/dhTuRhf3GCmnjwJlDqd7qRYkKbkzwSnnmeHyz0iO1BwW4dI6xaM
wOyWWq68bs9kICqp6KxiVkjRYA1NEkuU+0K8TGrLPNmFcoFVecmjXICAQjamdsWK
xWvasu2W3IO/eVgGD8NhQejIH+Zm1N60Vzws31OI/KviSJGYchYLypFGfY2ZUk7r
I/iPczC1H3weHhXQqkMngPM/jn6nT1YQgsaU8ergoM/NmFsvu6bgGlW12UMMjEbl
fYn4rvn4JMlVIzLRr9S0+awJkxnvVidKGHY0/fpFtpl8YApy+J0mrtcHndGGuXWx
PdS2B1kpSTFAXFSjBEi55QnG/1SQxB07b6d1NLnnGSgH9i0//BCF5kGd9fKoaWJA
nWWQ4Ahkr+ayKyoLH2Q/bioj0G5mLhDdggsx1MZbEItN15kJQj9p1bf1s8xrK59V
/gSladPku5VhSsCh/LUz3txPPiX8LLmTSQaK/vbkXGM8BIgloe6xHhyWz4j02EgW
r2VH3Mh4d/USrzWW8tqLGirOu/OxbPMPyl5eeAcLhAlyG5umOWDjNOrFXtVfWowe
7O4Igwda7jXj6cKgB95McT9ulQbj4hjm0ubM17EGrOm/cUq3nCkg+jSXzm4csJAa
v5cs73jHFDY5cOG3tkG4iTqm/9fc+4BxUPHqisbp6SCQuiXAqgcFGCXpt+/BttAy
PSEvUadNKfSCvCME7OdAPDIg1n3Hf9sMJENnSKZECMO0hUwNMUeXlYE70PzrjB5l
3vcKYCeD4DAY0pkiAjcYLqSOoCHHwn7lcGfpns9YelDN78a/MLo4OwYi5ZQjLIE3
oyHtAMEQKPS/kRE2OlBbRqKBPFXJO6873GMQN304qQaXD4f4e8Ej5wV1DafOP2OI
aONqp6xnkHSAUuOSHQRx+60046rlEJzxWFTW4Oonl4+PqHmape7TdNSSz8ynSv9E
LU8ceaU7fKmeGEJYecyz1suFngWqciZl/whFibVj9as2hKy+euPnoph6UK/cEmZY
i88KY8R4PfUn1mKp2aUjwAuRZwdp6cUGz8RtfObfdXj/i4DxGqxKKDZ+7FNtHe3F
jb6sAfg+n1VbueJktY77h/2hNnUGPbPMwwprGfsPBfL7g+lsGSqTkR2TXikXG0Rj
u8dAWCcNiJ7V/vfBCX1pPlT1714TIPS0LVcHZCInHIUo1YrrXCXe2LqStvBLBjoO
bkyU8agBalX8PUtxaQgAV2HzGWUBtO15BmzHtTGxrRrhryo7+rc6LR5wT0kBCH8Y
cgsbdi5QTrNTSx+VfIllxFsC5aSlXX+IzzCuOFhL6a26DyA8WDq+Lmz3rr+KAhMY
RpV6HnYX7ZoMEfTmZaZ0ILCzV3JVS4DLkZ69Fyugn71k1ytyIRFl9f1A1+1ePH1Y
NMN43+auh+1xPbVUWDQKg/F1JMuyV/1Zw3Y2VJf3i7dIG6w3QpOZz9mEJ6VwAtCB
3ENfgYrQD2qRPp45ayDTAURa8/rrN4asiUfIJjI93LC6jL1uGKoOMHgaj0EpI9/a
lVcsu8zTpUiUqFQM7jrBjOwGZewFMP3kn4cewEte6zRLPdovNZzjDe7RNi8b5e1Z
3BrYZFmIXUtEd0ZlbXcwStfwnfDXSb7DpeUTHwd0T5pUqYN5/7p1UeMG9Bcl2WDM
36AcSjYXmIIOqOLz17pDAN1wPCF9Mz/F+jkuW4M1AWH2Q7t5LCyYGkZ09z6f0yEJ
J8bvaqp+SEiVYTuylguxuyNToz1kIaEbp/kNrnWs4vhEKWy3vNggJMbRm9PJbwSi
h/hFeszgziwMsyyHjosxjVQR8/q7h9iIrF96x4xbL78jQy4iOm/J8uhOuJsnxRIr
Vw07tgquBa66SuOSOg/Hb77c4MHOf7ezZG+cAEyX7UjLkkB87Tjr2RteiK/F09zm
94Ue0EScNuCpm6v26nBr3pToH/Cv8Q4V+GsgU6t5kdarj7KcOOd4a4vHmg1ndBkn
6uKNIsezOoO6JKaspy6ggFksftCknZ6RHPDGx+16+IiLlfn06hRjm9d9cvZ24w6w
GlVtH/yfymwR4xRUc4yK+IfIkfImaQO0Qxly1OGKxgWfOGy+XZmzu/c1Ky8EsphU
mW3UfG7fIVAv0ZaKZhq+j/ZpLR07KR1J/XUqr0dIGCArgsmteo2CxHCCG9NqQ3Rz
8M1PHxjAQ25Hn6lZ+d04qztuZUUiVwZZ8bFBqpnrEc7ovwZt1n14A+shofVn54Cv
zBt/ANpnQ7d02DBpiUdSz3pWEid5mg0sDRe5VTV/hhvMnZKDyyFNBwsLyMF6RsSx
nDDUWC6mpcuf8QdbftE/a8pwZ7QQUMQce35MtXfw1zevIT2bvhzJsDugdB5VTE31
5LNySmew8C50ydXhdVJcD2jcFg5NWHgHQqrpP2WdbieI/FqHp26bb5ZWl4DFrZK0
48+xPpy0XPVW3sNDTeV+GJFF8N1xm/kq7os5RK7KYvgWEUKxvN9Ib+Tvb7QMh96R
qNPXFwaQxgGtOEljC2R9UfzQ5xj1QkfrNqth8lHcEVMho9VHCQ7B4VngrNij55gg
drAM6vLuH4cgkxkFc9OvtrPlPSFD60SwKLueNyV8nEBuD1+GR8yWEluar0DyHQN4
9RrJ4i6G1ya9cxUZH2yCCBscRMcOuoSnm18epz8vV+2SVwiiE8GD3drJsxdd9ymi
NUkpo5z3GVXVD5y3xQbHwSTqR8NWWhC/MqZQkMnPqDQnwwom0xm4PjSWS/g1ji06
KPEVNXisY45/mZvEu60qVWo91xF9JCbQHXmmZbKjQfnoAT01mgQC9B21q/uev2UT
Xob6q7kp6N7S86RUWIqq4yJcbsrmvaY3il9XD17imINDUB9xJnZgrsNidkrTqrWy
HKXxQBcWwjFPdkcbpiCM4lKwVUnRek+7LONjYkIjwEmBgNYpI2ntvbuTCI0qS2eQ
eu86n0H5l+uNUN1tFZn5H8NKZIhXjHVNiVUigxFKitDXvH9cYAP4g+D2Lcb7/wtl
SZ0GvCh6Bb8jB+dJwJN29w485edXQKX5QLJ27NjKN+tM1y8B8iDLFOD+V3iBKUwq
bz6VanV+uyULB6/0fgKYPb8ppse+vBw+/UyT9M3FL8o8eWd7m9otvui/+5PpW33Q
dvaupMvsC49Ve499cGR94Ft7DSV+BBGIs9Xb+f0d6JyuGgYCs3tKaMiEwB+pEa8J
9MXADhXJxN1Dy/HCglGlgqU9Eqxq+qwhEOsbYfIMCgUezpMCVB5u6CqLwgu33p0H
T6iNW5GFKmFPMz9I9GgE4tRc92qLs9rU7VxSaifUxQPG4poPkPtA45RZvUo0nzjw
75LiLYCJ5y47MnhU3nb2skoYH0HCVlB1YOwWu8dbmSM0BPmiLeZVDdMHYi2HuQAF
WpleIK7wdsTPO8K2kFXovvCApTwKQ2o6qLHg/FQfSjZqpRo0vEkhzn2UudcyByWy
hui1rEYaF7qi/QikQw4qzXVfi/dTvLVa11cZYgZT1ipFzcLoY+WuryYFtMSmpRF9
Vv26JHQBUvMizuGHXq6BwTF1r3W7d9HM3KKZmOhgMsC1IugFN5t0UbtDi268nQOP
OMm91Y9SaEBxebURB8NDcDuEkj+iFsUCC+BBstOujSgPmkOoM5uFrDtnD/vcpYnM
5SwEuq7HA0R5jCcbk0XQm969G/RyOuBi8rG8HpoAY+c2FIQRUQu3MTnT8P5TuHK9
C7avwDZ707bM0xLfeeriYKDgGJUNl0RnQab0ApUlIutwV/4l2fLeq/euD8N9VNtW
AgrKHGUc6DjYkFbbM8BBXVbivyJ2NMmdT643z4CkH1SI27RlXusnhoDmuqLM0WVE
jAZKhHXFVUEeKyeUrzGM9La3+CsDu+K/lkz+pVlMV3fj+X0fFfguiKiGYqiFgYbm
OWwivhan+WdDlNiRMGHFqInR7aDKQAEaPp9uOIOm28b8/nMSieHwWPD3/LYniZcP
vNepe+3sxRLaq7gmS29kKDVkKKR5VsaGgcFpQllngUFRpkt8BP5I0So6Z41tvN8R
do3cLMgLVZiBkOrh9eywKigJdRcmNC+aIBx6NDE2xM+HskZMCPEl3rPlqGV6H7y7
IBrDKapTwLusXL4/XgLb9x2tsKABIAWCetnMydyUp5bcnBFhNHJCi0rPiyaWa5dr
BrY+BuczsGYnMIG5WI/0GBEdVNXCJ58Ds9uBNYwemNVfdgNcg3fhTiJ7E0bE04Xf
IuI7WdYslXYwk+WPk/E8pM7e6iQY+KKW29Vm7C0oEtwuRdod/w2O4Kf8lsyaVnEc
EMbm4YEs9jBSYiN/o8ffq30PMg8V1blj5VPWFOKguhhghaHes94HbfZyZ2Wq19jN
lViWSuRXy2h7GXGpf+Se8gf6Qm2fVqfNCubq05Pe9IkzwEa98z3xQsodPbVlQrLP
4TRSAjJe2GIT2PAG+/GJIoaUhYK9fTTtmLFKPsPsi7Fv3KXQ0P8t+EFGBcOPKKtI
+aY3RRd63iLyY0fuargUY6OuidMwRXMnFGxPeOfOO7dWrhuuGJk4ebdUhe4jpwY1
8ToY3qj72Pe5wwHY7iAK9RHiThLxV/LtwnCCDVXWzJVCXVUFu2g66RKGA5iOXtVZ
oj/yIiESxqJZywJR7/Yv7TurLOhkWg7itYkQzHq+QCWHb2pHrBLWS727v2vzOFEz
FegWN/D4Uh/TQ1xLPE4kvJOpxURWBrsgpIOt9qoYDYD3EllLLh6DjUvYP/LlCPUS
5jdsX6X6AwYwwIXURwOID8A2+acqufbxwmAMN/86w/Z7Z+aH1zC6sXsolLVyv9u4
zzqaipBGBSaMHzYvhnjm9cw3fwb53Xs6V8HcISj0797xY32gceyvGBSP2/xQuADB
Lq9i2XHr5eFGNj0Avrag5KzpFfcVrb5NCqGB0WYW0zOnnJRZ2rl8EyyI+lH/ydyk
W9nyEZZHf3YmXq9ugxH9kZU0sRQxdo9NvWumLinCy4JvKmGmMm50qwprjgPLFbU/
Iz9kmKUZBcJOQ9Nxg8SYP5wtFvSHe84zXDn4rotI0r3Wko8P+wi8hTRiDawzLB7u
/O+4EJV7+W9Z4/MY5QtGRP1dlWGYRe9xHGsbp0AuYc1SV607PZkr+J6dK+icEH0o
c1hK5wvorWYtbW2e2+E0zcVVhWbxkVTIIC/xE9dmrtxsHJTtIyYu7Odl9aWA+/w4
8LnctNKHDvi+ZevYLirCsuCIaIYEMAP1ZZXm89dn9yBxw9L/9E/GjY3nspzUk/iF
2yN7m7h5V73ERx8HRUvyHqd77t1/rhjNT4JNQMiQEB/t6n8h9K0NuHHM5QYgwcR0
oX9eawJ1EgsYtXBcvBEVZf5VCVY/B2vzK8n9nnZzxVIttPCQoBBOKBNlzLYtNW9o
q7VquzPXdsak2lBTyqxl0XOMqg/KpWD0p9t+3bH9St3c1a4PW2PYAMJau28u3IFA
DmHIBcH+CCLVep1aNsmdqojxPPZy9nqb0KxiZzO4SiljdMhMbB3WDSEC2rUXFerV
cjQOgMRUb41PBIec2h3sRec1q6YlXPTCbg61eiAPRAKbWofwMwgE84ido6ucubeg
tYCSRdLSHqXm73KLyczApEjCKQ0m/bZDPjssgJPvu6/5XZ9qK5CYMfcMMvxcVsJ9
vrTSFsMMH1lKNB/iFWKgpv1CWRhBJOl4Jx4JbFIofJQ78GCiA6q+q4LJUake5h3s
/opkduJiaNYTYy0z0GeQb+XBxlF2a5Si7W11nNdBxVm1nKuPr/0shZ5QqxAK2FTJ
Ln4x5OdrtdxjlSr+bXgO3iNv+/7qHRRn44jQjq60e+yV+MC3aEVfMxqNUCmMLVe0
d4LPwFtNgxbB/fBVuden1bI8CRyTK3QYNEWYGWqQvW/p/PKxeasKPwzH/LFrxkhL
LJb8J1G7GlkUW9n4CrsBsCOgxoSXLOcxDT9u8+QmKO+BJ+IEu3Lgt7H0hQQs2zse
DoD8YvHCsLChlslyoTS0JaDruKx4MVeoNHCf+2MPNgg7+btC0FmgYJAmWs5FYmuf
R6+BXca/28Z8WQ3aVW3K0ZQgQIeTfi4sQpAi5xWLJjyxRBR/WDCfpb4Fvgen2EZk
IQ7mNxD4KJRUrd564Sm2VeKJxViYDcL1A/lGd4tf7PdXi0UOPJQ+lkEKleTe52jx
1d+affVQ4rFrbXPOasKP9i8vcfD8S/vh0ELgZ39GD9PTQgQyHF1e+OtbnYjH7lVB
Indw+wG58OlVTetU7JRm4SVTrM/Dgna2AQZOXTxnsd7sQwl007YZ8lqDHh7W5NFP
DUj/pRMsiIvdx4ZLkvRG7YJ/izl3PpzkTXUHgcU4RKoFqtLA8dJdMD+d8adhI9sV
YMPNta9aQ2cW6xM5CNAb8+NCIS/4HAiHj0P9tyy3U4hNJJn0rt0aRjuyJHGqb7rs
pZ/u6hJjjL33dE3gPxWbj+QQX/Om3/AVlTgfqMhiOR3rFrbZYX/PlfYEHWJa/R79
UCyBsP56Jm8VI0VTWX+UnnyFZQY7QNTRY09OEHXIY/4wySQqrYiLgiorRLX5D1E5
L49fXUe+gc+7cOTa3WMk8o8H1bzEs6LaoEJxooYozqT7t9Fd2oPa9Mzz4Zg+VNq3
f3WvPECMgd1XT1Y2S/Dy7mU0Ha57K3FygsmtjdEAWRXo9SEtz4anZajx+Jt9eBED
DH4lriyUIrdWwuXowl3QXqoPtLumJrzgd3TLqeo9KL+cyReqFrxguHjfYTFsCtIs
R8QzVgujloT3H9DFukd2YbMuavBrAJ95iliQuRtfDzw84xWa+O8pwzjYbYt0NvST
E38Rf8ry7jnE+3zSUa3hLDUBdC5mCiN7K6Gqz5WU4h6MJO0fYxY38Jq/4zfIUu+K
n6s9A8ZoaximMKKQYV2h/pvQLkg/g88QUG9tDIQiD/t0ChIrE8lxhOl4V7C3zwqU
yFpHByOsq2M0CGtnUB2a6MxeV+xLWJT3rm3aoiglsB6rlF/zKL9/6Edtqf2bPmV0
Z5xKSgfFWZ+9o3jqT+zWzkFHPfltVRFqgHYJ/57p3jrLecGEBBJLRKywc/BwR42R
9EFh08eVeajEfSo1pYNlgLF0wPw+1WKGAT6QOtm+cffF3mVIEikCQJ9P2wtpt1cN
kv67M3pcfVttO/0AbUri1RplQ/pOP+giAbsiqr9PIEHpue9sZE7hMySJ7JTb5Zm4
KRqmsja9aEZHNmX8ZvT/SMbVJX3pUJwZAuFeBxZaNKUgB1iT0p9ja5ZGppgiyrsC
zloBHb1753TmXBzdBbPNZTyeM9TqcqHBEy9N+XmCuexQsh1MD1SK6/XmWSm1bPpF
YjV/crDx04x5jErbXg2BtUkDVvSnhYgTefw7gZ8f3uB9mQxJw2u5SgrQZaR3V5FO
VrfOBe2DqtiqFJjZpdcblPO/Ub6Ng36sV8OQnxbqStIPg5gOYYnBsHZAnMGNYfeS
KRn0s2tRkmSIV023+lSWYYv4Snb8byuqMqD+HLMxjCERmH3teZvDEPdZWPT/QvFk
nbuf41CL9uU0biCevWtyd6G+gSMGwEQH6Py2FAu9rkwrjwVYtOxXuZWk3xmf0YC9
qxXqzzQd0TkwF2y1Z3jZaUkEMzYhopjMchTlNawqLBHdl/wcWOc6Ux8zwaxwhIVn
SUHrkcEt/sU5c+wSxWZuW6PeizXZFdBrkEkusy2W2SmE74VTBPp3UoOj24Tqwctc
hTpJiAu4EHvgXl7g6M6yxsigx3a1comCLZrTHSX5PTkFWvJj9kBRftYE23mV9vuE
Shjor6Tnx+QZXRAVYJENKUyFwM6kLkjx6ozlUfJiJdgNR10WkD6X4QNhldSkXBsv
qdwHrh1nkIIyAxk7M9dMT2VMCUImMRZf2uJOfG9nAB28WJcBQMkWpaLnakcsGeCj
P51TU8mRlgQECC3Z5rAApmKNuV81IpZ9ZNDcR3U4+MTkRViWfBJuc/Sr9cqZVtSq
LpNVtKdHjokJgEN0JjBkJ2GD4VqK57E9g94ldgKq2NnviP0hguDzJZ7XjrSNI4r9
lfEdaHH4Ss3PlJ3snrcaLlGHLKdGaFPfI/SU79D9Z6WfYSjCU0e15JXi/6uVsRcB
VZ+BJMaaP3dDcbWqfXOboV82iiR7S/vy4m3teE9TM2OeId80U8DbwT5M9917h1uP
cNFk++uSFKe0k1mY+kwWrONlj1f+M64CfzTJLbGmYENnvBFsPVhpAuJTaiLADDjm
b1k5FKl1K4r5aMvB0MJ3FAa2U0rC76gB5PpH6NULQInI8DJip+L4GgG8pW1dmjG2
Rn4But4zecQvJh6iH4K53GoY6eD+Msiy0Gdg5z7efFanVIHXNvwT78eym4WNshSK
YsGwyGJ20zYuUVLYlNKUrl4b37TOM4GYUJIYGCV5gxzVVA3Bfacyx8lGu3RdXJEU
dRtFkERB3l5l5sTj2wR9e46v+vtTlFGiI4IaSFSqosJHVvMbmbk8dfns6iS/yIXR
BUDNPyOIEq2gKZ2CsCluuFdMuzKwB1ZhlfNIIRjLPJGO1Jb5cIMIvV4yLJqiHv7C
Erm6RSMLB8+4vMTVp+m/NiIZ6b6Eyy4UvSiQVZTL1VhQDEI0fqSf0VNOOBmKDg0B
fuIxOmgigIm3E240nEnE4Vc3VM0Vsky8sftfIExILwwvxqFV5s/tmsvxJu/yD9lm
aC0Nx/zXuYyL9FnX7gpHf/ZJKP5FRhP6wEhjjHIuX2BZ3eyOz6pVIJr/VcRHayrW
iXzfoFhNmY3LviGMy8ymaSjpeLiBb4wptOGKHJmtj5+t8O0E7ZN1Xqi56WSbGzJp
fJg0fgCBUyIoOaznKXOqqx9T2JwRff45CgUhAozUk4ecencMazqVvNZQ8LQoVgP3
Y9xctVLIVrpTryPk7dum/9kKBD1pDzyXAaegInb3njyQwl98s5/L4EiTP4uhCYr2
/qVw1ktRKcMTnnKuqBpZYD75SaXfLWu6wCN7YsCw+z7GGqNIWAnCjqo0PmQzKe+F
K3++po8St2Vz2cGDQVixZEh8kh1ZWv4zUyQk8KMBXZDIpT6K1NagH9OWjba74fyS
Rp35g0opJP/IeA5tB8lNr1g+BbVpLJbLkrdGb8dkbKU0sjw41l7n3jUIuCOAShM+
h26kBtvYqhufavcJTrA+/jhvp9gNdlWTiq2HUJjY4ae+r1QmQJQL/Ch2ybYPxzD+
vqab4QxKFsFglP2Ks9adB/cXvUf9NHAm54u0GWlrAo5ItupbEkNI/fwsqXRMeey1
pdTPRP3ajasE3Xvfz+doD6/ZsaPbOitfYWCESvLs7xxpRxzk9a7iAFPyReRfHbuU
ERy9gWA8V9Ey+89Os0pIcMrKsHQVH4nV+RCymSu75yUXF71cmYRNHQ3rv+ng910e
PaKR506MrwNOXgqta3U8rnNzT85gwP6HkwoWXmc+4bDKTYSsGHKRp3/t9ghnDC5k
HbQ/bUKU9M5Rmvt9ty1wJfEN0CK9zuEotgn5SwTei8xJ+Sk9V171clEpZLZXnyf4
jYY80a5/wpp4ogK3A8ODHVW8dZI2Lg+r21fNxrpWMV6WoYoVLOzL9YMSnRnj8ywP
IQUPstxBxda0liOoyArfMn0gkGcSQbjiV3q/H0CRv1/u19BMGIKgQgSJQCNm6ymY
WG1XV6nGAI77gfAkE+A60aTppZWdR5y3gag3iYdA7N4SaVkJwgKdskaTySjnLAb5
35itwSFumdlQvbDCP1NkUHu32kOaVzDQnBxL9Rl3bYxFKXRY5AkwrxJPAMiB/zfn
LgdgiFm/s2IiTEku5xTFFM7hHGRj1R1njT/3lyDpJ8/MNBJw7E1eokI37pcHry+6
m2omfvq0wXDEBSCBJO7bsTGaMwJWEgpAANWnvRMgGyTFdwmTFU1HdEcCHgtFeiwl
KLeO/jADxR51mY7C+lIQYYeVmDryQeee5mvHDLkBEhlEY85hXgEG+04xGAgz5o4S
T8I+HepRfc50WDaFaY2WvYln+e8fDtBBA526zyvb15R6XJncbTdL4xrdwd0bQVv4
u3JuiUCNuohXX2gdwWjP2scWTXGf7y1ZpzOfW8Y3IVdo0lEftp7xb7Jyfsn8dlZy
tOifT5QA+FFDSwloCpHebzOjbQEnR+1M5rMB0DDUMKtsVar/auHr7UzeQXXsGSQB
sC6tqyH32KGr6Lu2vJ8SWjDMISPxuaVwdP/cSbUzIZETCNzkgO6eSJYdpBI82u/m
HUVv79/zZMSYySVuvw6WUEAwQWzt6KoTvAxcciUb53J+GVA+1H8P2ilWDEz8aplP
XITen7l4vPg5c8PnxKd0alDdUXJkoeM4Gj+Y22qkm5jMJrQdat/td+/J6gkOIvTg
JMEKaIElq8l5FYkH5sQiE+YSJwckROM7YAmNtdFiDqbmuZKaoqqFWHtI9B5XXH6K
ab8OAhNw9wUwHOgXt8jN7HnUnmAyWBckEGeciJDBvCt7l6frgPQ0u+zbEADPolyw
x9UVZlr+RonD6C8lHi1NwPKJOI81XXk5oAKXrGUs2ZOjcttMLldnP/8Wwm03pUJQ
5GeCO7/QXnn8tgfa10Ig32GClI/SFmtuU7GWUAEGTAKEzSTevldWllcUlg5P/SG2
8Wz48cdRU1OvOpdQuwjYP+FRLJjXGZ80GNH4IcUe6IUJxQdm06qbHLXNZr5xcGp4
cfZXNajTu/QaXH82E4KjwZEmEIykNt0/BE5uDlHLaFecXN72IMiLa9WqZCwX3WlX
B34JQksdOBlkMvsT0vMy+nPDy7UGJhZU5mnXuxqhJ1l9bfaXtCXkZy95JdXjQkRX
zrHvbw3M9l7xHdmL2zaQI+fww2EPFPauD8LzwQQv48CZU8d8G8Kj9D4wAH6BqaHE
QrTeOKZKxhqpkuZ/kBmZTHyksQPySIZXZDEpsFACR/akdCuxEjtVVqDY/UUyI4Fu
CaEsbUZGn/u3uVOZDhNLO93/8yyQ+etHS4iS0QYAR2pBslbLt6vkkZlAYYpzhMJw
ZynfAWO2k/Ztfqc1KcX6Qc1Q94Dl0Mt19lFUxoiCxcgbQ+GxZbKqjmKiodytdhhD
lLWITQ5MYQ2LIJyQ+I8r0Wbfv9Zf5jcQ03C6WrVsav5ZEzZsjjUQUWbq13H+1yf+
xwDw86kGE/d/qYpqWDS3+WPnfRrb/Q0Pe5Pcn66QrBzd+ktkLBeooaEgPIVecHg0
D7SnsupYcTkK4lxR2gTQSv9lGLir+eegaM2N3k1LflLHYI1BbT0YSGLo9VZS6a/p
OPYGuWj5+aNDSolcWICLv+RQT05uQ3xeGilAT0xWBIFV46MKCF2L+OS+a73F5B9D
1Hv+CMVC3x1PxW5gmHzDqHdz1o2WfWQNrkZlnCq9ev4JknG92dNmvMTJqZ3eLqvy
9VvGgcjJIUNcktQapS2+Unxps43rx+EmHDaaEOW7BghdJCYTwBe37I7PvDBxlqeH
aXJ8JtjeCOKUbIpU8ERwMPH2SBYNT5ic8GgxbLAKOZ7ksKjSMy+iG8ESh80LGgqA
iV+wEbt6hfwFzwJfrw26YEhaxcj5o/zbyYDPw2x2eUXhak7idJfvigS63UK1K4pY
EzmXX2nf3yOgbwWXfRf/i9uyCaqT9/W74IATyqxGfzuz1qliPonn5j197HX1nAh+
fCKRsosylgDMgIvbu4XUylqEfkE9bu6ADeQfpkefYi1tV+5P3OzqDgpaXFGhCsr9
sPcjzPGUF1waO83EDqYenk7Bh9UWm0AXMuqBxuO1lUk5qTePd4IziT14/R3NFcBC
EJ3FyrPBESeDnOxvta7GJqXdw03ABihtWlwId58xUI/MAfXPwibGMP8b3DH9XNS9
AokaELyK7s4bDHNbFWffH8pukB0NNTee8/2xQdEvhPC+Va4qTZr5AHs5zHnPwsOq
PwyJ55wM3ew7stwFK0fW3nYJdZzx64sMvyRkvL7sFl+ORShA1KKX6rU5aqvB4k57
iAns2BSWQZahcij4rJA/qyvkiEZccey2G7asF/1MCzntn4/qjhdtTKP2dAHHNgvn
v7/+hmkrXwZPO68DKfkw9NOdhL9mYKuQ8gHEslkUns18PIsV45vlCghKEZpsEHcv
gBULjtOc1XP2Im2PQ3RpZOaNlEJCTLD+kObXS81hc9qeIZY0/FOq7Mg1zLQraYZp
UqyNfDgOvg6TE6vDlQE492p6Oz+uXuls13BRALSoK1Er0gHsx18qgSnKN1efDWe0
1jfOmkxODwRCguym6c12g3bRa2nBZcRzsEz9dqNhZL/c7PRgg4ZDqkrNbZZzhHQr
D9rcB4bXSGIfkqJGjFRwkCLKlXeCe2wBW/+dw7l7teBWHuFzmRW4/LMtjSPW2qvl
toDiTon8hXBE1k3R/8m+U35gr2Bcytnvs+bwpG9EScWbpGKx/oJgF+jG0yh83E1V
/34K5nbw7TiViX6/wTuYlyVLTzbp1PhWqLZHUd4+q0c7i5FbQmYsHtfxUCS+cns3
grFoZdNSEQMaIKgiL+CuEO+qyR8SvzX4Fprl2XXnXjZQugqOf1EDpXXJ2SP8r4FW
rnUeFezYx6VThKaM4hwysGbps2IDSqf6AzZbWIC5GclMek28oe/UrtGc4o79APMf
XYiGA3BKKmCW5fYQIPP5YlqKOkt5n+5KrZNF0d3/eK2FGkhaxwHyh7369BBGX6Jh
gyI/YF0tLAENlcfgkgPziYh6jj79W4mvy2kL6p5j3m8SH/LoIPtSRhuCiT+kBcHv
1ULP8Nq2AwkaWWCEC/q8mFgJSGC93AEHwSxpGgtbpsnjZj+be3vpw98F6me53KCA
OD2x6qIQpW3F/0Npd0sdAOTmUEcP0imNdoHW7fa+31QrCsgXvikCNZhjJD1OOKkw
4i2vjyW1YjvPcYPlOCiwTu+TG7e7egYtLZcikRixLPowharBnoemaVDGG2qpto82
GXNbTo57IG7hJ/mTuLqBV8h1COOJR7BkGYugX9DO0FOTytqzvZa9V7gqtL2P+njF
rctjZhv+EAfqXNfTtaQaKjp/YvVRWWBBFoFrhQIxKjUGOPAKvGhp7NrPXmguLhLk
9wF/Y7lR0NptlQj5sQ69hxSc9LEPEd5sX9mgKq/TQMahEXzsvfuafXz6LSIqmYtl
d6m0t3uIiS6w9fivyEY8CUhjwV+ZurExcbP/QAOMXdeRV09ztapu9VbiI9RhD5Y7
3SKUrBfaDaVZBTf65t+E7Y5hlv+SKSoGIuHQhaQkiMJiYHh38ZNKYj8HPzGaWhIy
Ply96RddyiCaiUQJ0yRvJZYTdNWDhLbO8IQj3dzABwVxBH6omy27/VdhIrJVsbNZ
OszzJxJIVD3esc7QwcSgRl1PyD21Oiovr7zHbBKT2Nzdt68YcyhdKSk5UhsFlIdy
H0udBfJnr/UeEjpqBLkZbBf46lxwYerEN7bsnVLFt+D+zSWpaQIbwjPFzJzrW/rt
HaSzRFpmhE9jbzoTWb2c+gGRREwK72hyr333SxbiKyFIvF3eDMDWYRY0y8sR1nHd
zfDi7/mNHlBW3eCSqQhjS8s9YN5uh2LsAqtBKHu5x7zv2BUblhxZetZqtoWR0vai
IYGgkp3U2v6xy12/y3tfNmzcQ4YmzittiTnk/pv41u5sG8V0hSStRUpyAlIS9Wo0
4NXQAwKRfi0TwvDp0Wo+Wdu9bU1jPp7iq6QoIPOJHWjHCeB9LG0H8/oGl86WBqP0
BTKZYIYmvf1kOWpzP75Z2jXGZRo2eoKL8Ers7vNb/qSHM8u5nL4dz2d7cRhYxdk+
pcveaL3J/s/Unrrfsj1wZTfWHUV1LzGeIcqRwE4+ppHjEpiFpkCDdDcbdk7NETvX
+ASfx9uTM8M5u/RAn6UDgkg9pf9e8oju230QRV2EPqssXeij8bDP2MY28W+TODSa
xEhmbHWaWDWJYqSCrrNjzOkyMDqXVyTOsqDCUVzG8EJWe1Bpz2W6a139VFm6jokN
Nxw/u/vdUp+E4GQRHrbaGfwU8jjcvtHdyliVgnslCULU+WAHfUZQxmo1/2lUY73r
lh5Z86HxYdwmPahRikV6xZihKa/KyyP7hAA65KcqnTKqtnlhZUmC8La64LQ0wGdU
NYiVNKMGt+gR8TlRaSgKHzd9LrY0G53cNraMSx8sG4cWcC61M0mpJ7RZM/YY0duC
3Zw2w4qg0oOIgfirnDq/4jj9t4ET9i7qhwzx5BaguvGGLXCIdZFEqwpf+gh4hQCT
+obZe/l8yKvgz1MzQTbEVTh3IzY9J0vz5fSjw+V6RIsHdPGOqJ7YmOJpO9fvTZGe
JL+gSVh/EzVafCUPGonxmIz8XUtUIDDXTINl+wDrye4cUC7dqRyM3SOoD545G70U
BIvSgsrRyMJnlGRw065UIUNeNJQWzJarEsVMBg/23zVATSLfMLFZEzUBJEU+wCnV
7skfMrxai+QqfJHwQpUgWTSaU9d4QqAh3UW0xoCC1aItgHACEM1ZYCzza5Y16OLe
5nmEa0/pLu3Ll6qIE9jveMwCQgomAsfWFylrxjn7FCqOMyAMpW4xNr57p24Jjfg7
S9+Qt90yqr5yArJiZ8pYyfO6UyqeLmBimen5LQwroVk8Lh8Vmz1jgqSet6yXLwxq
Tfl7FPZhgsDyip9FKiryPt69AbZCzzWtd1nZxyqdFxuwAAQtYQ2pzFnuEVR0BYve
ppHAE0VJjMV1swT5YARo0Mup+36VA+I5zaoAJnUy1QK8KsFO3cgNoea6Px5A5lfN
StZhqn4ZTR/DgIU+OHf/zFXuMd/c7a+pTQRDqkoACg8lzwgvs96gSLe4LYjGdSbk
2LK+peXeT/qdK1VG5vUXTXCfUbeCoCgsJC9q9CIEjeAoLaD+TqI642EboKEdIP7E
ZRBCbgld7k3565ADfkE9Xkw3ih9if055eVg38n2AkKmQ2vaqWgT51LIox7huJm4l
BT0aJEEjn6Q3m5tgnTM2+OxIUny0Vx1oQSykgYpzfkXexnjQnPDDOpUirvkROdmb
cxGoaRU/p4uRAz64fdrRf526tj6YHextPTdfCGP4MgpjicJXabpkatQqIjT2/Hbz
duWJGRRfLYc59xpA6O96Gz5u/Y/IMeD6CpYAncXc2VOeBQVIONUAWkMhYtah0r/M
TBy48JQIhYYO6YCebaUy89TTy5wvhHwtczeEdelay40bOpPoCTGaW57qk/WRa7HY
OSE78N4OOW4H5mhXmva3BbOCm2Me/mKa/zM5OkMoPD2ky40kpOREa+3AR9let2zt
wBYSxSV7fyo8s2lymz7anyRFDsZKDE42JigHAi226xj7J7uECmQdRKTFOIjq48HF
sBL4N9qZp55VYKql4qZQ90sXR//aXOaUnBDQXmBSBQIAaFWVPvdbHyZY8//vXEaZ
pMIeGjAWCYiSyuignvcs6ptVnvx9guXxjcuwTrt2vfmAt0J15o6CMB/VkZcM1iSW
N6N7C+1TzLyg6ep/70fe+bcuGJ3pSybvRmVPLueXBRvyj0BKzc4jiubSlOiXen0f
UtWyzRAUtqSwl7/VbD4OObHkKjXnHZvrRouewIuWi5OPsCD49cMghnoP0RuoR9s1
bNpU3C7N4pbCvUiva2gMFWDxC/73yNjhtCV+noCJ/JPRTNvqTzlGV4g8XQuej6bK
rvmB4QMKuDDUd9jL0bYoTIqjk9X3Ti2kqgF4zdf6FXxkzzV9JSDPH2YssvSWKK2R
nVtg4eHqasycyPOUkp1DRzOH3FjyOyVotCs4+/Ust15EOdVY3UuqesRLlJo1SrMd
Ea1RKnLIzLutXIcLzQK+gdy1myJuUtdNv+DeZZvTrvlulEjSewYB17yb4NcPGMqR
zy1zYocVvXeWh/js9fb24C5YaNnXO3MdHlOK1NHIavZGy6SFYYkZbSgLUC4yvH4L
JAWTRu3rzwvabacBbAwOk5WeTAllEaUkiib00v9l05osi2toSED7dyPwIs7+Ihcp
hIkFS1Dw5x8GkP8kqF+1wZVZJ1mETRIlEsGFFz12cG0qfsEWEzSkI5yumfnRWUCI
A8/WElWwqz2EXUxdmIeGVCNBd5t273U+WicpJgpXCcRFHJYuNxem++voww1Ed5Yy
dqR6GECYUNUNte0Ht+73mTzfKkCKwkZOuaqD3gRaJfqb2UB4T92VlK4hTen7qt3L
A+SukWx+C8FvkVjy23PtkofHqxdAQ0aULe15ZuJ5lJQ5CxGKPMM8AZ67RIpZ3BcZ
BBmW8tjQ4j8PxVftLPHmwBDWT0AMZgd9qajjspXkKsyveRHxgnlhyWB1Lwc2Al3g
GZ99JWwQ7jtNituss+OZF4gOUg6DHHidddnrC46t40pjq+dZL/rrcx7EQpvkudXq
`pragma protect end_protected
