// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Mr4N4hTT8VRrmXV6SaQ8MhYOMvO/RolzfpxFCsqr9vARDFLaYWREXljvr2nS7fFLrrTcDa28U6Nj
/I5m6cGglzjYMtvD3gzumhMy9S+fkn/yz7Bw6rJaLXS2Ivpgr6XD/ah4nuCVxpEpVcDzPr3A4Qfw
6flQlynv2ymvTiBFT543SpNysXJuhMUmEjtCLEjtg1JtuSFy0UW89IL+DEZ1wZ6ET+RPNlSfXimL
t0tfN7NY9VapIWSahWfywCrnWEHId/1uRVtogoJ9EKlqoMfG9YFamGyORS+LCzAJUBODDTL+ZAOV
mYvTdHto8BI6JjmHHuIXKdwQfKz6KBHvRvRjHg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
TpKA3OswwBr8MpA/Z0glFe0zeWOOOp8bavEM0wRJatw8motlrJPahR5sBX7mG7TdxiJfItffMO9J
lJY8HC+T+DUkrzAbYv1LjvFFaQC0kVRFFm42DSFK9NLUmAbTm86MLXPeR+RUNWs0Geus2humXSRn
wRFQEX/ere3OGRiOothGeYvDRNBqFMTOvNSE+PHzQjTjMfjG/5X8LIUYQMuIZAvTxLnvsmpCoR+B
CrYsowd5vjUYke+9YPH4CQhjwc4NeP3vZ/0ZoKB7FoLWNTR/fU57U4Sjx24BvKLzW4/zXlBiBoSS
Pg/NWwNfexDUMsT07NJK+0e7VMjvJOuKPM3taCnkBKWU1KNDNfCCdcm6yvpt0AAnPsmNLobtKiBd
w2Ryn7xA3/CSrDRUpqPj+Roch8Mtf8RHo9HozUX/3LgxJa+pRI+uTRa/YW/i32wbwKJJZh2MwfEI
K3qqriXaBKauTE09549gPT8U3d7eo8gNI8MYmQrgJoJNCatqxmvtYySlFeHjf3BCSJVtlxOz5/CJ
btjkhHgk+22lXlMb10cw6etIbn7NCklU1IQO/Mz20tdO/VsyveeefBNJOithcrh6yrhQqLtGiiov
InMyCLqJsC6Q2zsl8of4iyzpNxY/vfcj1UGBzWjzzNPBftQ53visKs32lXsHA1gf4GWB3/3C8ADI
b7z0SkNFZjZR7gJdx9vQjS3PSB3WisTmN1u6g+A9ESjL7rU6DJOjOpq5M1SAbFc4cB4DfcIJGTID
qHC45cB5SwQS+k9E0epzYumLI17Sf1I82z+MjABeQNQ39t+hZ/RYeUzBGeoN5jpCk1fwHxsDOH5U
gD/VmvZncQyfM4VLm+R3sxji4TCxY48xCI+8b6t1Vk3V6gJT9rrhx+IF034lIF2K5uHO0UGFriTH
Dy1gQkbcJO3JE5dYo0sE2cnZqA2YY1L2KZcknwkZTRIKEjdP6npm3fBDlLZhy+a5XTVqORcOsNB8
5uDDZ3xLuRP4TykrwYV5ToBKSlO7/UpmBCUrJFt2N/ZMU07PW1jhzu8EVUmTl4/YZ/dVpaMUzQ5P
x+9cTThG+Yn0C2U6I4NjhLHleCNNlcSHcVThBHkNs1X1ViykfL1hpnvnLcVcPvW8c8xDJnD70j3u
ucx5b+BVcDMtuQQnP1Ob3kGVPIGiZaUorc7wuZr56yPyWNnKGekCxMkCoZXYgJt2iwMgCii6bu4Z
WteU3AXBMwXT4kiFfNQRB9E9w+iF2WkzioaW6BcsuhRIV7q+W9RucCLxAs+l/xBQn4EG1dJ3BV2V
kdEjW1V5dm+1qoxTbR3PqgAgOmZPHwHlLQaYLXFFqslyNgDOtLZ3uYlKvRfGkVQkhH/N0EuzP7OM
POatpGXmbTdXHs29MZG2ouC5OmIpQQsW2oJaUdknfUKJScN1kdlqsiS13Tzqdhjj4nKrfVVMDquo
sJeLASQJZGkIQ9KAspK/1T79v4gkdurtyWO0skMGdpbfv18/lm5C6d3Ame3a3/0RhHWE/5HqI62H
1Kx9uPJreuaSZGVbz7kBtSO6kI4mTHqFcSTdKGnkLA3SnU0SiaV2Lj4jQXGFkJPorefN4GYEfjKs
1SNmI0JfX8XFK6ysTDQ1G36L2oFlAOyWOnEeMlqJidMdjiiGsStyW9vfMiIEjj0BDYlMHBI5dUvQ
/Ejcaor3DwapZJK6gJFrjR07D/WVG0zr+o2OljrdXSev3l5QUWh3smSfRpggCRWQQcI4iedvUrT7
zxRADmtlcNX+oUN6ejZt9W7QjKNvAHLWPgXzL5KgdzSgpGt9X9XQQE/+DF/Psr1H0iHATGtERHL9
6esHBKqKSizN/A4cfOAJOHXkgSM13wGxc5cOEaYD2SXqNb2UmcfsV6UDd7kdAImS37/OmecCOu4c
sYXrvoTkgunZdRXIAzUYV6D7WXKd7avyxStbD+V4h0l2pTfT6uI5R5QobhELg5vRenxcMSh/r6y+
vxiQTYKnSpZVWICIWVKNASzKFeazKLS9D9Ruud57sbpmfS7Us93Jl9x2IRV4Ag3K7OmdMrF2lSuL
3rl3ZMydO1PExhh/mVQ1pWrOGs2T69bP+eMsDkPFT/4f+7+h+zMZ3G7FzIWg/sbRpB02w/FLAvCw
Yqko16xky6sX0kshSbzvhzu5hYdCG0soRit9THrMjhCYU5eJOeBHgzmkuEBJ/DNnWgxLUJPtooqC
ORsxg7arzFhB/NdjU4loP8ksMPWZyjRL1H80ZYdniKG/x9JlloOEQaYM0cD8cFaaM8QDyz9OdD4d
t7BaMUMsRfTIYgyuy/CHTiVk/5cRztryetQJA1jz3dPsy9M1DkgX1DxPbq/1PQQ+qztXukyTEmwD
IRLaiiDNGMgsa9/4aRRRIN9QkiB5ONATXDUZ3IWKZuoqNd7ekT/EmDHao65daph62gVJqDHCvVvG
KTXfY37bKigKZbE4sSZTnG86/5bqOGHpE0fLv2+Vm2g7FXwh5gQPDYUyybfMwV+pV3kTjhIWjKGv
gAEeSZD11Q1H4Z/UZgDGdb4ZBqpQLSct+rbVsG6ryknMqtPV1ZAirQqLPu9/VToW1IG8+MomEOUW
12ummSYCH5y5gCKysnNNF3WzSd8frB07S5OtZCBAGN+9hUrUshS932ciIQUNCcZJhyVO6bjwxgC+
NDluOCBsK7L1KeJ7wm38MHuCh1B8x5D25ivSinvUFeIDdnUUt0iZGN3dKKA7NnT6mZcGCN47G7sI
LKa+bRUMCUacgEIV914VhoahhmWVxQh6bCFACJOG4PoWcMA5eLOW8S7p+DqFrQpMrNDwbLxrbobw
dpRMpFtc0qsv8f1F5BSwxh0DWJ5eUmD+SyYvRZ1zBNTvmSwfX9VIXHZjWxVPurhPRukQgMYwfpRs
qABnUn6eLRgnZ0wrwrdX1nkXmeyDXRCD3TeMz5kwo6fF3nKjFz9ATYBOmxJKkoOr0uRRqRp+DoMm
XNEYHDOtcGDApT0KXx7hMmcuMJ7uT1V0JsD0mi0+QTAPAFHTewLn6P0HASwKmG1kl4u67R9bTRjR
Xicx1Xfx9HQuJ6vA44+TywVxYMFnMMXaDN2DupG8Hk0xLZWcZdHD3Pe1hWL+XArvih7zbLn13h+n
bT+9vaLve0nZQtU3xj8QBjMq5WB1JTc6sn9tK0uNzlvso0H0jJR8rhQcYn8W9XwSjQ6itphYpslS
2AtfbLZz9TO9aJJj/ZwsgYpwuwJzJibFqq3d3xlmfnlCx2Mfi1L5cJUARTnFz//wQmrSofHyMUHs
7i+RpVk+sv9Fr0ED1ppr9g6iTEgkIzamm4e4prT+w8n4U2+wfkQk6vy+UGNPKYu4xd6jexIuIAaC
jAXcZSm4NJ9ne4D6u3Na7yNiclYcPRVKR71BUl3l4H21eUOptmGDzDiC92GHGVbgNYP+jgUnRyKW
QkymVcOECBosqrcl/bhiPgFRjjs6J4EDLX7MMKCiajzsgbcK3UXP9ZwT/tv8D2wXMDvwPfxcEkcG
poiUi2oAUfIksV6A8MRU93lx/0gg8eOeYfTfD0iuEYuGy/FBe57ovHVv6AxD9rRQPD80rq7vToqC
H7X5Qv28korrAO1V1i87xRadQtLcfJRjXGjpyUY38tsDHeJm1QA42JvFv/L9RR14ugwYTMBrxZNu
gmbdjGscsg53Idhy1JOTxW6mLm+JZo0InKU8WehUQ+whaE3bOOzejKiofcYqr+CVQ0G/Cb59F6/P
NdCR/Vcm5ChfwMySR0MZ2Y8iTWG4gnsuW6R2fQkKB9y0+Knwak0AaZPnE8Z/Xnibu+xtFrq3UrOX
3pwsg6fkhqwOwn0F9sGLC4yL37jchXqrqlDLA451XIdSDJ0uKt2A5FLgyhoWNEa6NSyLrv1CPT8b
7FB3x61gGpiD1SdM7pw+jQ0bzsf3DNJqvq8b02DqjIBY84ksda9asZKsC4LQLR6sae3vhg4j/Rlm
wQ1il9RT5YqZNR6cb8FjiOcszasUMrMHGRNlxM6jseHcs/emjlxMMBFAwF1WEpjgDBubwsJLXa82
OMjLVki5cxh/GvK7RdMjQCsTxxaqG7kHArBkQ+p/F+uIyFS24GllLwhSJYqZ9dxo/LWXnrHBWN0o
lmOGC74213Z4tGm8+o+ZfAViqbN/BfPKRMLoYK4JwpgaLZVy2Ho157emuLKkrmSMt3YHluN9ZssP
o8hBXtwkzH+FvU4BqQhi4Si2oBk5NbiTNlSvSIis6ul6Hqj1mjZynY3aM0idbH9iR47OQLTsGeZb
NnvC9Nu8b/HtHEy6bwzLpFdrSZ933cxZPOEcDfryN9sft/HC4WKijPovP5HBuRFzJq3ugg8ClvhK
EV4c46owIT1o25CqaXUCG5ymwvICLt0Jp+6oSr8VaEoFnFCMT2YWkwuYpOyFJBtFVwWbbxqYd+ZP
g8oq36Qzrbaivu5NqjtKQv+Sm3O0c0vERuf8tsQX6dWnzyd0pTF25VwAAgNasGuHueiKvuCjYupt
r3x82LlzxBIRJQ1zuNTC9Hl5sZq7b+Cn5ItAnwH/SEUL4tJwiPNrGumykSvmxtmlfS3cRyrWEDPu
oV0Qu0lmuX2iPtkzttGQWmNZtUcFDCVHmmO4y0+oELOE8kj+A7RXchJvMjPS4/5m37BaZIYE3lNX
+SHCLwtJEoJ5CbTHbWaAVTrir6vmk8BhJvXbUNc1rwX/lO36UrllRURcBFlkTMDyktVDHeaYNlhv
ITJf6ImSpM1W7KEq8rzSQaR9LoYgCW/hNaRddK0nuej8FqzHgBQKcWQH7ZdiJ/KfDWuvVZkTWV+Q
FQ8BBQAulBQ562ma9AugTrwAaJZV0B6e+lcET+8l1Cz9sjeImkQMmzdV1pZQ194OSCFaBrZqy3N2
1tG4OTASyookZZqVT3b2YDKv3PFa9iYFbDeaT7RosNTPeV7YX+nzT1VvxOXdj/ydo/JzbiLnEQv2
CdUKzZAiAyvWjNxYaQ3UeiGiI9VSD/G89GbVAlBjKh1cB7HLjnsnwco9d5P8OnKF5RWwOxJ6a4J9
wgOxEiF/4Rg/HxoPH9EJM0UpUF2H6VhssHo7WxdCzXq9hqbzFICEgmE3tmQFLmIgmrcG899H+4Yn
wTFPKb3isE/1zGRJsHw8DVg0AqOLuN7Y08jFk8lLKTbZnvkTKeuq5ZD7vSApAunomgbo0u1poFnB
v2vyRMtCDFn33E6WddM/zv4UnrwDxVSir90dWMvkXh3yT3T9eS3Satwg81yksQtDRsujxNs7fCmH
dvyRsybW8dlfaQjaER/ttT2/Ov317hslwTvYrgSkrBNHUkoORucR9iNfgU5g5dQDns+p8GN8w2Fh
S7bremjl0Od2/Ly3sEBAM3TFeHTnKnbtu5FC44M6BOQtvvgN3wn/QkLY5H4nqjx6yHFZWEk4D8Rg
pxOIksQYUNQG/du5LZaH1EPFWI33Nd/VDx3K3y/uMoZI/EHoYxW0TxBL/v/oSLUKxB/sGsbO5CHa
tCDOyIhk6wckflcyLQdrWUJ7TqfGKsVxXGkZfTR+cxq8k9g57YxG/HcOkwsCrIFn2znZHJufT1jG
F4lD9PKxRgVUKkctX4VXpAGfVmLgJ0zl5qYFpj272lWwhYkqDPzd15zNHy4WvsLr6G5APe23KDau
488tHcTauSfbDLwAoVfu44TqLnigw4RqmkB3htPuRzBzbQeLRY9soZVW7zuLaK2r8M1xe0YJojDk
+FcsCLy6MMU6QO/VkypqDi6iJ1xoa00FkN4o9jY5M2TVpRRexHVx8Eh4hZ2kpZinygFLF5gCL8Qa
HQYnPxEEDLLklKY4HXGZBgaU3oQMmQsJ2ZPK7oyFdoHpXI6PCjKQn4bjX8zCLw4R1ta20yssX8pD
3e7Kt8tZC7I/RRnQKNtTmKEsGwb7WOewivLAcco25DiQfhWwI4+5bbw7WikIxKsbqNk640Se9LsF
L5fMSITuOz7suIW6bF5FPgtuL22TnRWQw+QgJJM/+XcF9nLCz3mGuP4j+0Uzh0JQI0J1ei1YmLSc
lcB3KunOTQQL2N5GjfZygMWdbM6B81ceEXpOYAgP0RuaRs2CqZyt4BPE6gWpskVpHb8ydnRiqg3r
PA2HJRnYauOh32AcS8bZnzxXpriPWVtTKYEwiP8B5OCagSjGqNTo+0qtL5FPvHkUHy7RyfemoQ3Z
bX/BQelSp1zCKJIg9zeUsuSNmI8SWBErD6Ru/ZOmVcGofQyD0zPvD3r2DBgdqoe6KChWfhOvknnd
6582UA3MoiFghN8CPXYgnjG8wv8iEwhwB7JXzBuYOICfJ28njzTKvvPR6MrrUljj7MIs1dRFqmSW
U91ow4ORjbmTlXlgOVNknfuR+iBzLRNCz5R8zz1EeK977wLimZF0Xytm7tUUb+TtM3NLTW97MkDZ
t+9OBzwz8mUseFcMWUzNMwkLOLvBu2GAnjxBDYHloFx16JHVxv8LYuRPbgzTPL9arkgzrGuj+mMw
ZgsELdAB0511x294JWXql9cdheqiJg4aqunydngq2jS8lkY0EfR8FEinPj115Cc8Wr0HeiJXO7sW
R98cDoKJhtq3m8ZY2lnTa0dgYaN0BfhMcy5C58ozvCrziZakPmQt5lTkr3H7XFvmK1BMlpCqPajk
gRJRMlfyQ9F+Bm2igYSNdZrVKOAaoSaR6H0/ihPyc2F/s6AzPND15Jmmwplrm6Rfxnvhw1t2HN2t
35x6x3Y8/jiDXAkXmsPtjc7p2GGPKse7wtNc26rDtZI+jYHVvU0nVwUb6HAmMNuO/jDSgJJtbKSH
zKIM2iHlzbwIet4AVapXtVFHzWOQpZM6SHmFEbYa/oU/8reUAoj9YaSZNRj4AtVnb7VxSmWbwyrZ
Nn12bwF0HBlvE+jBNqLdQhKvMaSUe/ThX/BIGGTkH8Zn4DbJH+cF7dByHpFWBK27xevJeG7ppO4T
DpgzYHoaXZ6F43D9G3YqegGniXwZm22CBYPrwQjd6clvIb2eYWIWJf+1fgnPl4hBQqb5Y9RhJCmX
QtCisSjA+Dp/BqI3xS9hr2HZfiwjo1333XgafPXPKFLpSAyYUBChd7XNbBaMRnCCFdlVsjPO8ur1
oS0PRaAo6N1eDJ/0FSmynvULaXway0vrZtBxuGERCOATgwfwFDJgLWKawiWSR7UD9Z9P9NdMEC2H
foE+F+YuRCy496xrG+FsbgNlYXy3S1QZKTTJNAPbY4JXEW3+v0KCeY767fZSuYVLqqYwrAVqg2p0
hxnnHRAIXmYbXZD1WLlApua65xkOrLREFKvkB8+mPiRxX9McHqo0O1JVpoSQJYIluC9TSyYllvct
zLmmNJqwjDWndBbZDO98HqB2dtQgW7zA0mFkJLRdXs1m+cHRQS9g6P1ct8FPp9A6lVgoExGi7iVi
0vlYGBM64NJXexPVxKx/i2iEZo36vB9/1ipV2dLxRc/kFq0SPi/odulilQogne14e1OhdPv0Hxec
k1ZQwriIGxdVkJ4zejwfUzlvt69mmayuaKSDmqglFGmM7YilkrBTlS9GcZzQjayumJtGAPwDmtl/
zy/IaN5kLauUS4IFj2FgGqPetGpDTM7jyKqVDgyGObk3YgRBhpcbNp12egvG2KvUMrGaoyKQzu6q
I/v5EP8AXKwOEf23A/SD0CWisxugCcHpwmlK4yLTqwJ0RdV+U0e+1okDB9dXOSvSwBrMfi8jMPXR
lr/p6W+kfCdYWd3qfH+czKCd2U/qzyPx97Lem8vp/fInZ439Jn8//uMQ3jY//5DXcYQZuvF1eplE
DLQXdIcr71c0bf3BwKM/Mqekiz7UsW3fnEuWxfZp4M2DK+fy/HtQTfo32Ru2YW4cEkXczJZMEIgW
yLjpofcfljXxJ5p9K1XpY6j3209kqK4GJ3rsVbQZEbUDHhK9oiRSRX2fFg1YI3gUOy0jYZGLlp5k
eYhOWMlXnJ0vDdzCztOuam2awNjthZAL1/AEwjOd5ZnT+yscWDmXg0hOsplytgxEBXjMltLNl1y4
x+83qG2FDIv5AYB78ftci/0wEeXLjidodWBb/sn2MSQZSZRv3GVuGzCaCmbEp5wVHRMQKpyZf0yX
XiBdZPu+iiZkYewHtITCGcKh4OZ5amoSHxIx1h1J23m912vpSIU2SXRgZzQ1VwSmjXAgE4h1x74N
hyM8dt3B2CC6WQF+lG56Z1E0VjHgdRob43FgvV6sgATMhDCOdEx/AdmNcIPFO4njezsxixOh15GB
Ok1zBq9iGg05GcC3O2EMx7hIYTeBC9oB1+wPNaFl3nLU+VFFXLXy+WJtvuNOcCVzAlXWT8PUJIP1
HvhfUZdlMuQq1RU4AJhuECVymyH/dZC7Eonbj6Ci2JBlmHAAKwV9FAivR9lv4Suc1b6jo+Y54Gjt
7qW62QGmvjlUe989oPHPRuvfyIsUwpW93JOdYqWovBZAqD59iY7kwi7mmeI8c7OvkXTdkKIOx6Rp
5ruQFHIp28QkcmNHB+iosBebnNyEy8tg8yOEx8q5pBghIVfzQNxtZVgLJa9xlJJ5mq/rMJZHi+vb
0ECpzC6gFB9y9D7aM7fxBI7zD9Mvy0XUcwOHcNa020yu3I3OZ5F5RH+hf7chEb/OFEwO9ZQUTYb4
yNNEajufErbDIq33DquZDKVCYFfgEqR18ACdFmwUhLngv6G4NgnwaUyC/J22eGdox5Lkflx7G05T
dKqRpV5tj4+fDGTutW5g4diz57yIn9+jDOJeeRiSbqB0qeO7W6iCTc3UgBMt12yZyWp1WNTZrc+W
GNXNdAMNqy3lvyVJ0lk3W4TYAAzNgwZsT4Lxpqvkm32biCwHST0XCqlX4alAdahXFOR/3jvE10SP
eTP4GeoBsg7XqdRsXZj5EmxbkMAaxXBLVHoYUM0XHZ6KoniH2NTIKDv5ZOqax8mnxy8LN/+ilewr
+GUOyplJV3q9Z0tsaeI8bxRYXk3om7hz/bhJjhNDkyKHV0Nty4zgpkWkP8bIwslUh1JOo0OLxY8f
qxSr5KT6SPyqAUDmyeNjheTZCsUb5GbgG0sRJmVRTzG6ROsjmBTqkxN6x4JAc4M72Uexs3X8pdQl
7Tlm3BZjnyNBfembi4UZM1HA4ERopQhWQ2fUCrfx0zBYMH4jEXXMD+ffurC+9BetqwLhWu/hKw2p
rhhZYoBk4zA9y1UVsjR6hsGJinAHmiPIp2IcLSj/4cYk0acfxn2ihGTER58jjIcH8LISDsD01dtW
t29WM9sPGSowCqqZmkWF+BtHbdF/llYfZzXszzX7FHgVSufaa4+APY0cTwzo7E1ylQzueK/ahzja
hQjoRhZ5T1JmRMzloaSmr3jBWItrXlXQJwdNd6g+cyeSDpHKhY4u2/wH6PKSpGfT/bwpJzu2RI/U
16IPZ+Vj0zx7lStRLjwfchAWza+5GJmwMRwIuwsvxHRvFDzSRDMzzRIRMAUAmlIUb34iSvpOgfIw
OFOw+9urw0bbmoT1qooZq74XDQuHUgKL6qOKnK0D6oclTXpjn90OdgLE/cAv0zVJICZstxw6RPbo
8eqV0jIcqIjmaOMtUuA1etr4iP8es1LJWrE0DsIPsVbxaHktlKfC8tB2CGnmgTAasSzc0iZ8N9D4
hCjgNpVPmMHMBwHfAGCM9nrxq9QQ1XC/4PvUtXpQmmZ0DoQsNWm6ZkTl4U0RidpZdy3nl8/2Qxak
bEVLFaQPLpeqzbZUilhyOMBWyshu6ss1Ku53qIyrfIBCrUmpNhWETsT/ztAn1wE4oOeV7ThU3z5+
/uWhCmkktDdB1iH8dFZtpSgipEj1V0R8ZtrIWmWR9Iw/GUHL2hyRXLjh1lo7KlMmJl8FXJ0bLRXV
qjrfBlivyjS+BqgwXTOcKC2rXUolCQHXXpHZiX+AQE8ZwX2yxNgjFG25HFucht0/C1y5HFzlWcL2
g8D/gkFimyQC8AkMqgHvGlqBwFd6o+iZRFtEyDgPzBlBfdtLt8DYynFDkKJTtdKXsS3X6rMbfHZS
Yh67Py9NsCPrib8DOm1dJV1NkxK7FX9x9HqU6yOAQnoHN/y1la/u+MvSwuSqB/FPS29VnUwzYZN+
KzB+5Lxuh5UdNOxAQQL7nRQ7xo2BL4AfLtiCu0l/FyekI3qX+vCN7XSCf2np08/YNu7+7jvXAvyT
yoZ65L4RmWrHiUgBa9jvkfUo6yYtddXnEzvV/mlfU1865+VLWDXkKOkZsGZxWSjnT3NwLlmGGmaN
burybMyWo2HNK/10dzy1IO8m2JL3EnoOrlXiISJwP+uEtgOO7flkEWgCSUMOcyNEpbV9ExeBhhog
eAWeYizHckVReZpeACYmGXQ+LoSrxi/OFgmsOCPsuT/QBEoRFOpd08zEvWgykDEwVXGsLWO/GUuY
KRudiy5UTXgbThXEJhOtoX8RN+8y5iSg5f0cIiUeT8k4MKga9z/RbdQ5xCLfeT/AeI4R8tfbMiIG
NJnQAuG+lXIexgiFdvs7IoN12XV93B73LHOJ1eLSsoChloKUKQAPOMxhRhTpoqbslm8PxUK+2Qgc
3a4/wTqz4MeUmFHDavcrEHrH2mXKx7rJ+m5D629B8GI8vDke5fMMfA1rboWKNJBXVvsDHrWdNOPr
tnFw8EkHkUl21M2B4jDhiqKq5GYlySnuRObbrQrnspijBc13zt/3zdVXiLb+M42jzABY/6uhp1Ay
B1Gg8i4E0e5/oJdYeFi9wIm47qJVXiQAP8gTfxqK+HB23yZf6Epkl5lnZX9YuI84V7qN6dKF5+V0
Ow6JWgVLv7uFZgiySmF917jOZ4FNGHpnnlu5fRRtU/0DRkkKTNhj5PYItiQ9nPydwnMM8kVEwhgX
Ap0GZ3P9dXP/zTjyOJt8hEL6ffmGeFNmvtO7Y+vHlO6c5FKMlm108A+VJvmtn12M/l1iIw/PFNjy
2zCepYMXMCoPXT8suZ1iZh3crz9Bd8x3bRZXa6ojobKpcsB3LRp7SOjuT+Ri3kigfI4MM/kfmugQ
cMjdMqrxZLmsjGQNIlLaV7Tdq0fVJzDsDSr4CA/18fUjRhw9o9bXaqYg8PqyLgDBIAfjSouqQvgk
bVWYeQS2du6ltSPtbw/3f/U1StvnjKEc1qJQfP8VRvjXBTKwKkCTCUqUzFDklnikSWk7LQ6JffI2
TGI2r9KhpCs3BLVZm1crJVaSIlRvlA1+Yy1lYiJZ2o5OpU+PgVQ5awEEVKLepY+G4VrAiirNtDAi
PmBwo5+kXsrfhW2JJlb0iUbNPwaiphEsajiLbJsGSC7xLHdXH772IN9KtSuiFXnBLCVK3eskhsEu
kwz6Kc192ZEFaaJKTHSXXQZONVMDZyi21XxiMOb2FbbJstAgzIXPsCpAK8e5F7wbGKjWeVzywKMY
5z7O5V7Tjy9QH9Bm9EVOjrS+O+1sHwUGSEng01FQELAXmloL4cwWAyNZ30rI70mlZo3DYlYC3fBd
yXXjpmAq9KGd37c8bkxNzEYjaiw3ry2WU9QBXSkSzi87Zy5AHUs3aEFb6C/xk9szg1OqQxwkFVj5
zyOUHcTS40Ns6x4XwxzDTpkB+9rSTvnEe43vCVDgRkoyaUL+dkDaJaXyKh0xdfM0Xwv82w0HTKL/
JsC1QC1DTVojS6J+V2CPR0Y3QWl7f0NoPPUJtON2LvzOmevqxqQg7rewFlv8BaF0ax3CFZt35Rj4
B9t6vUFznL09c8Tjl4VvTpQn4NzlzM0lz39GrLi2GfpLIdGrSLQVf9mkYqXycXWIx5PT8bwu7ZCi
+aDvffzixkRKGm8m3DFmUQVAZR0n9nT6N1vG6tNz8jf1s1T6t32wZBeKfByRNsP8sfzYF9GjOgBm
mAa6gu/vyp1Tf9xcinq2+HEzAVwkfI9KbLuAlheWB13JGlKMWKJVA78C4tT84AsZQgqm1eytJKh8
1wDdFDuyV6RNxoYvk7/2jzFLiFS1dFNWhsw+4l4EX0C7hNqy76DgbYy711CvY5EhO7KK/bMnXVq8
XKqeqLP/4PORqPrKzlgURPT7JL9+WpnZwCk4SGR11Nh/YndvZnGo1cVmd05J/js+D8Y9Q2rQmZd/
1qASJkhAbThQXM85a+egOjjNeZZrpXkK9zSVqWvOFgpBsYnusYXbhMHDUSSX1tAc4Gv3y1sxHAto
Qrga8zzTuI0luUd2EQI18fTKH7uO4TG4iIF1BGriq3gH5yOpk0viKvn8hFxi9o6k7lRVbI83JoZl
D1dWmgvsbXuZri4oghiuc3DDL1AOSEK+DMXniTF4uQIVQf++mOdpupugTqxbXwD3+wRk1DkRgxqN
jZ/pvxxUGDag6dOg/D6AWzpiNF8+sbufINOgaMXbAZAflICb0UYgsDuusFMFp05QwV+4Cl9CvRh+
AYQ/p1UCzZ92FoOmfDnSrwGDGMPAyUN56MX9A8QMeSl5ZawnPir7Zrgz44KiFbVMO0lVntfALK2m
IB9c5E2MvwMruRgqlxQKwLGiyHwTTSkqiP2EvRVYxDlluRDwKWl1OUqYXmkC91+TailPqG48iDh/
KC++GOmrxzzrJLUl02M3As305cBnqo9jHesiJusgXpjSLmh0uyWlAE0KmvH2EHNsIY9moLu7PM2Z
5YbkhdrCaQYF6itYhnyacx5ENJ0UpK2Ns3WMdydPydLoa8vtELxBaQrJ6+yrjHBduWGDhR1KMlcM
zzMKimuCxsT1qDBbADny/OizMu6fsHyaxSPfjSfeuRpBdExPJ3JWO622zAfJWEEp1HN4EZ1wP/Tn
mMIjDt7qoqvodtkn7lNZFfdlH1hDCFpGA6aoSb7N75z03tPX/cEGz+hnl+KHnOzvRJAEDIarMJyN
6zgHZHj12p8wBLoIY2rAzp1pNUbNrPxU6wZvT8eIv4tvmK1l0OLfaQzsbvhUr+Q8DgTwc47HkYQ=
`pragma protect end_protected
