// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:13 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sqqKKM7/vigH0TA9qqaeMKtJVUHIMVvQi3JwsLWV1kRNXDVe57hJJKX68CRCjeHW
C4kmLiycVNpbmdrnR6GuS9IA731DBsl0orakYLQU98aEL/DtsuBHQx+LHgEnE2N9
vKLA4qgX0JFG/7FPg66sWGXE/yQ9QUFIMgh9IoAZ7Nk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20368)
u06jq3J3IvtjM4WHLwJYheG0C5GYIGj4eiLoRr3l2Fv8q3ZlL1CDl+x8DARD580R
q/RtG/CNgxBKoR68w+ysPSrW2uP1C60ryOWyj2Hx01w9cUfNYBH9yoAizFTdBQHs
z/qMeXnb2bQUEL2Z4zatnqQNwxdJWVXLRTPXwyIb9tXRZQsvK31u/yYDWkfACDNm
v2OOliSpI/PbByKfA+a3FiXQbHvBYW1P/+F/CvU2DLVkRk+sGH6Ni0K6c6J2f7j/
+wO2Pd/Yv6keVzMcpIfpP2HuQcsOqZcrGVXT3CrfRaOWGdwRpV4RX/UYP0hxTKC6
U/nBvx2n+LY+vhtKdkzqz2GPMRSAdirCiQww1rVWLfqcJ93OZYvtLjgIZGxwpbEZ
2VEpZDc9AvpIzOoFLIla8MrmJQuP5Fyoys0vPJHcGJQbGIp2iNC0CcBzyA9eQUlp
oEf/MZZffIc1F58ZVboBN6hwpKB+wk+0a3ALrD0Y7kTyBwnky/IXHu82/jrh02bs
NbvtkEs5dOqP1M5j8+c8mRbzQesAuWSCZC2jF4EBjykkPSLNl9h47EjSObui/0WX
/717Tz21KhKRvbLFP1+Km1Bdgp8kthBU83f3hXSeZU77A+2jkz3plNCIVpbs0eOC
ZFf0DTYKCYVot7q4vRK8OR4RmMDIhveb3oYHvICMGztsO92J+XuocC8Pi/ogRyg1
8MExxJYbJDNBz40mXD1ZMgO+R6gosZkLrMp0FfmMJz6UlKkw4uQ4GjCWfRo/5mXW
EhOCLrmBxCMF9OMHLyg9OBcZ0uKxcXzT1bh5Z7KFx1AKXblfTErymr4o3WX/t89m
gtuZ9CH2a/5w5ZC+pM8uLKtuX3eRwK//9DOSpRMLMzFkVad971cYVWWOBxrzKq+U
N43r1ljpQ/h9vnsmUssE7ST9f7TkM1FTCGhOOzVs2LfjvWA/wtfiO+5rC6ClLnmZ
SWDkrHMJtKKNNHOWjGDcra/M/8JndNmWrZTRe786iwcdJku8Tglqyl8Y350fsNaR
tQH9ev11A0+V0YTVnwzxFNYzA4bYsiyqdp1O0LCc1JafnICAPPYGRwxHNjNctptH
dLhjePsxw8t/3IqXYTlTvOFbkSKhEmdS9moxoAX35mZhB08CMrxiQRuYDSFj1uPM
oijjuP5nnxRmOfIx0CgtfiMlW5fqZ+fSuArn8TX4dppYsIgbPlAePfLGg9DIBTNX
kLCbT6Tb3I9V9ZNTWV1oEiTYioswCZXZYVLo5IjN8wtu0nY5RZiXlrEY8S4Eua2g
ghHGBMedpvQA5d3P8YUPgBxTKJzLkx6wLmFtAVhAM77kbUPYpsYT7m6zgB+DRdtE
aXjtr90Zy8RH63TB4cBh/5D+cYVAg1m90mpM6ioGSWVkSdrDEwmc+m9hVG5NWuS+
glv1WHxtj99bIkqT/XMjgDdtF9e+bmIcxhgIBNGVym5TbW4Pa3E3okR5kuAtCF85
u31dtya9d7/KZhhpfjPMBsy0SRFlLAgb2NL4UmXYJrAwqV8045wUgak6LWs6M+bR
eqyqmV2Su9dB7FFRtW/GNe8Z0zGD6MtA1slhRXpfgUMj3W2nTXPuiTuwA8UL89KM
a/bEWrVX3UZFkoGuIyrT48KFyhNN4p1TTjTWl47P3tsJMlV8oinH66QxV5Uq7IDn
8M1pyPcF3dUYcHpc716gau/A/Ch2KiU13bd5BjCcPpbqM6GCh7WmwmCK6bGy909x
GfphgwveV0ZEgTG9TvOEDT8rBlZiSq4xCNYVyOgo2vDdHWOfwgE1UmBGN/NA6L27
81O+QHxmCAPuDGlhfwywh7rAk8qoW0w8C3JuoqBlyZvnmElJEHddTea29wntXNtz
BP7BbJh+Em0jJWEfcgY6vk6N48Hiiy+P42WHyZB8CXjGbC3AM3P32koXNeQ2dfv0
qRxd6kordz5CKtjKko8xWJ3CViuEGkt+pm/eB+CM1XoAeXqNEGfZ+XhDAeFtTX4N
DWosDxCd7smLknuw5z3/dkzIivunqCh3UYNWn1LonSHx729uW9KCuWrSJEbNbJ0S
A3HRoUEp1iMG8W5ozBX3SiApPmkZnYtaFOAevc91YCr6Qmk8DYYfCzmSUWuxQYKO
e6Xu0Qan722kIfOuBf7CbLC4AAgDHttWqUBYEGtD7D3TsUbhbpdUbR8K6uwJZAkH
fa6rEzG+gIxoX+iJTw9WKuNDfT0BgLjvJjHGRNzGgrjeRnROmEYH0iJEMEqLLZD+
b8WbRpPAa9JspRYn+1m8NXpSfUKXxeFyCG7WcKNRfDulyl90zJBVtz8D5t3VtG1U
9J72SzousDe3iLONqg37EKKWSoM9WCu/g+Y3HqgUy3MgunrzHDKFlUvZ1N3+XRv0
YDlavi5Hn/C18znkbpw4gxd3RpylQ81fQWDP7RLpjwvmXyH/xebsYJlxr4hh/AlU
jsmwQgYojpyyS0k9KNPNBoArafahgjOrV2N6Hq8bPUSA2TES/Y7IHcKxCjrdrm0c
iSjIphCZw+qBVvRcvR+rCPoMvQBwzp1A119y2yNB66Mutj+FHEPUFkybJa9XYdaN
XWgJP0/sySJ62unfg1gkMvUhikAd1q+traS2WEwpxPM78XKrTgL2GPsxhZDx1Usc
KeIx66Fadk3IDSc/A2h2T7rPqFh0Aq5I6Lk/K/TL5JL+LDD/XPZHBZmnqLnVLJuW
toXwIqsAYZsYRBeKvgyi1CubcKngMXsXqpgkHjd1ztHGuCmi/iufafDfD9lX/ryr
PnV3jYgJDtfiJmLzamTgrY4AHky4jWjvcojAPMBpLGp18uQXS0TvBc55HXPsAA4O
HGGyK9cs4Ua7tFrs/e+7g3rZdkW2gLGYQg28HDotpjqi9Nw4bkxxLVEA9Teteo32
ObSfDapIM4SoyOTM4Y222r+pDDElAGol0zspLQv56rpwfb5+124UDaxQ85b1wYaz
/5hZUyk71vWhQ7d/e2T5GHucrI/MP3g/oK/zMTLxrm+HDnoxGr7kH6GvPyDHC0to
0o9UN5zYG8uBdPikYR7nyup+mvYQhn9mpai+uMMFsZuSWlIa/dDi2yNmx/IkNa+2
yQeJKUh/mU46i+tXKD7KOIfNJLRo/3gqpGBtG7yoAWjK11Y6nVkf1wNWJBVaJbaH
8cpmQUmxI2/80dpfg330xQ6tL2Xiqa8Tf1S9G+SW/NIxFi8/kuUhtJPxnbFpWml0
XQ+xNa1Fgvd7t+UtYh4tAdJgEzhC4dG9ORkfOcSWM8tG9ZH8xoDrREkwK71Yfx56
3xxZK5ZrIBGbkj8xWfXBqj4EL+FJxOPXNApoagl7OUIfwr3Pphd/hqg8TzW2xhSI
qKk56lXPyGeOrCq8i6z36FOLCUn+NCI35yZPsgN+91BOxrk2mTNkhljSDaPf0rBQ
gvYGWZ4JM6YjJ7wJZMW7Pk+KkDkpt7tbij+VQ0/wv7baWrXMmPdMs1ww+vKPVzMQ
QE89+q2d2ypznMYEasiZAsNJmleTXbuKwo2kn0C+Z7iqPG4Jxo1jBReYjzqcILQ8
mQc4nGrAIMD1RuONoFPjchaG4h+3gAvG2sdiKeP09ES3fVfmxP2sAauvPrvX0GuH
+RlbhD6sfyI5bBoJ2VQIzpPtop3fDFBL65mHCe3enhMXF8C0eOMJf+54PVf3Cy6w
8FBpuelrWp4MxXQycV2cxvRC6HLSunuRMVNWhyErCxiWLBMQIAbnz/Sh6rbZzoxn
21ptQiR2dMCNl58jHLUjHZkJOJ3zfPcW0BLF1rKbItrWjJw3Eiattf4poMD816pk
Xj0HmednZT3Y9cAfw9X9LtcM+JaIJ1thFwnxIPPBZeCkXKw0OanMoRqt8dMMULMx
lWOzPiCuD+OZ8t/zizXpL3VPSJQFWof94AsFIsQq2sX8e0jt1YxHtmmQR4hrXUXH
MbSaFX9MyRRsEJ5QeJhYfK7/IKrZUCddXC8KRbPV9UHObDJ9ue25m27pmwVCGatE
xJlyLTn7WNLx1xw+Na22R1LIMBo92WLYhcauZzz1L9+NfHqgXuBqnA45Mraw/UNd
KtnAZi94WikuAwj8pHhVd+qcAtPLAA0X3dKzQVMs+inL0oaEvh9ox1opr/sA62Dy
kFhodDjQN/VR7rh+bhijMtfrrr8LKcYLrgDr8sQCNEWAK3/E7fNglWQ0SbZyeCiZ
HepfzFwhB/Eq2R+PoECowtcf0wZ3W7+vfvAhKNv8X/94CNaIu9AK1/LI63tJAU3N
13jxeArbld78Ne/XlVTnf+7DGrtxSkCbUy4vE/YoiTwrvQXhGVlD3EH8/6e1wAts
IA/Ou6THiKGdTdcJmsNGJOUxmH7/L/6BqzBKRRxF6YhA99nNo041M2ZonC/F+VRh
ALkv99mIKGP+ro9zp5Zn2STqUh4WNaO/bnYW1mQBR7QHRdAGymFzJia+w8DLBPwo
SR1Anik3jrnN9IFoGcDDl1dzfuveBxx7QdoquhkHCxZdwbha7zuCCGC1+T9Hd4N0
B6sD4U975uUs7q1YfI2VmxRIVN+6vbHFiJs5+z3n8iI6s9m3+LaLpEowhGKxre9V
grHppQ47iNUI9wZWMMV506zzT/3EucsH21m+8Qgm3HmS+cBI756IUA/jB4HXvQlX
SqH8rArHYJbLtPJWIPlbJHzPu7o4E5x7QjgiCGzq6iEHWocmBLkvSrjvdVKHf2qx
hgwXIGfxR0SN6qX2UZePL4N9zrSWZfXKqRPAF0R4woF25KEPfsjkijC+VdQ5kxka
o9fxLndsBV8jUB9k4VDmHGKZNIc11o+06SqaNWjYUh9iRc41qbrzdVqBs+kUrjbt
ReRosXXi16pWkCMgfCxFfle/ciiFCxH2lC/wXXTkGg33E8hdvW2WAUucd3N7x8y2
yZZR8aV63cxHCXkRtRg3mg/BnIHo23xrJfqOVsvNaC0A+1BeCRs9gSZMe6QZ2Srn
+gmawwvdOQqdz3g4VTiXC+VzRZATrfQFw7pb9HBhdrxYvAoV2zenqs3u13f1XsOA
ElnLfXuWvU/bx9zl6BsKcQw5dxh/yROCeu5qbxQXPSjT61LdfWxdOd3qpp8zjgmw
4R/Wk7qjT14+jO6EOL7b/5mJnil7rRgZBMpgEP05Nc7ZFPdew5o/ihVgWCuaXb5d
y4ZHbNzCGppZzf6H6yMGu8gEzhg9sgRWpi40Ch6rXhOF9oZha1nrS5AH4TPWHDbn
fg91MbmhXXPu1jh/joZi25Oa/z+ICmTsQsh84t3pTF98UGrRFMwvRuJq4551SfAG
rGx4Icfm6qQsWOYxgtmwZ6yIGt6KtTPkDI7x9rhfc0CRO6LLglsPUUFf5uSgkB3w
NgSkx+np4/B+WQ9RqRoptCo42rL/aUvGmXmRRGG48lVvhuj/Ku5LVF6Z58Z7Ak4h
SPoqY7G5PFxYcsFvNfBCzA2sXfbrJtQNLW5dcJRZYZQNVi8wMYvuBnwO7ZksswdY
TzgeG/gq7HjOQzYS2OWEyA3SrTnSrjZamblA/88Y7nh/EDrPMUVjWzWB0CBhPiwG
HWMPfv13UuNqEjNdBhzpyfaRx9X/wJYUAs24fb5unHeUOGeKw9RbRqPyK41O2ot1
+Lfn6zBXPLHtBmaXlvy5Q4MmULN+Ak+w2davx9EmiE0a4Wv1MD1UQ4sUGbLhma5U
jfja6hG8z8DvdEvOEP90dygdg0OqPRJbCuAKqao7z62mWLByrNUytEhDzkWKYk0H
UJT132sf9eJXZy93pV3rQOkAcGHgbX+CuAGNyR4yFsVJJGY1RvcfXkSg3IvrL8em
SwcEdSq1lizC1Xe3Sd4kIPe9oapu6dMY9l4Of6lFxlRCQercfqA/x9/LntcfKEr1
XZnmkqG6AJVUMVfArNHLbadL2+bYugRrkHTFESHAXiAvb0RmTUyOgYOzF6t+jx6H
TOe83aM8E0dfPaaQV9BWoq3B4kIVaA9nmJ3goFWbaDbKJ3FWyByZGPGraWaHFGC2
GqJnkXfetOW0NUcyD9L0Nwi5Lxg06Nd43BsMYtXUapRtsR0E0yeCjTUvCFgDtnDB
xKffjny3BvUxRpjs6HhAT6Fm8jgFEXtXmWLwYAHkxrQ21SIk575hsRVKcZn9APHu
0ru1j1XcRmHmHCohDp/X8MUWy4UPGY9OAqU9Re64IlEWHEhW3v08eio40WQlUeTm
7Vcm1F0UdHIC0lImPojXrZ3Ebd03e3QKKpprd3S0/i1/nE3JM25kq/3VCQNHDMnL
UAQ+JEX6oq8R+h8QBWSMequsA7wQxIVxdCZJZrkNLOlCfIMD7u2cZSaSxPNrLrGi
lL6nsdFQdzu4Z/1SYVFxrFMGip8zKdRfhvtc8RSOdvkraoh5lgQvHRgvIAHceqS/
jaZxeC4kqSPSh6Y9mtr3sm1J860jFTvo7d5ZJ7IwPPmlUDjjnWTTM5MEoYIEj2pV
lSbOj6EjKXYKTrblSFMOaGIoVpuxZx9/Ad0iJcmqXhNtal8btXPsx+svWd5CeP8u
2WACU5fxwaqklwrMq8RdpwykbKSxgoMQAyq6Ka+0QWq+vwIorSkRV+k6RACCujqv
1UD0exSpGgvTRbga2XtLM3h3ZaHkSn+6tQdkSRjfqUWcO8XytdP+ldN6VK30xyoC
y7CDOL1+mvP6q0bh58GjTg4LBQ12/nsuPTL3by00Uuzxb5K/deBTGO5dVbCozkO8
w3Okk1mkc/O/A3Ozu06w7lCCY/Xd8pZpgs08AsmYWQ8Bw6C4lwJt2WXWe/gDR25+
syrKT2LOUbgq3T4iCSLhefEkaxDUxUupu0WD5ALlvm73lv4yx59wx5JltWctRfsJ
eqLalIFtQrRZNkr7vmreGx3REvfGJ2clVTqYchT6fRqBaJBBjnspnyBqaJXm2i7q
0hNWHxmpYQ5A1jJye7+qtOD6haXL/zk7SeiHNK3f0RAKuP7rkhZRQnMv6nvbh5XD
uidUcYzXu6Q5BC7zm2pjRyHJC29P8FGPDnRBti2RtqF3ybtWq9cVcvCwQf4xUTWE
bW9SQDOsQbLaDf95sP8bYI71AD2l0BVbBYR9Uz85DKWfv66I1TpfMC8z4xFuoWxV
cUm+o6ur5pqphJK9IVI7eJXhxBz6QwG3Af0uRFHlFBCmCySHuiCzrYLEU+yTpGgu
jx96NfAuCw5lMupZe9oOkrx8FA3rBrPtBfjM72xOBYl5vxqP9cqAPNNcrl614jYG
tsSdrXg3ed5LriOAPqcJMi9wgQeLCfMY1EY2CelPE9fs/R3g5wMUfYXuBNRpYOvc
rermMMTusZCT0o+K7sjNh2Zx28Sn8RwOBK3kQJmHah90j3FaJyUPZ09PXJWxe5vF
Fu0J20DdkalaKTBfomPno2gknFSkTMpwMmsV3gnaxSs8w2pxa3HbQ0J4wgVSUZXz
pYvei22yNLLQUAXnotC9jBX7A2XZzu4SU40sOVZmoYoW5AB+d+qXYlhwqbFyIvQ1
/KdJyWaHTC9iIUdfL+fdgea81Ao2FuFsNNRGb1hSiXgCLVgsgEXGrQWLuv4yTvjg
2XsvVVlVp/Y1SEvMN1O9KwgnKisgpKleeD4b25G0d0EmEhMH+0mS5ThoXriaqwdu
9f9wYeRCZrGnBATjPVYuAWnz0Ns3cVoqtVTyKtXTlAR9lcJ9eWMSYIerd8eH98Zv
ndhl0izSXyE0FraTS0zvIdPUJ7iPGqupoPf5T1SJ5bEoeS1hNTGBXRUW9gm0VTdT
oiBRP7ditbH7C+b10NBcWU63vaOJjdVoib72mXcYiM4QUKLT7Z/lDgMqMprAbVEe
kPYyJQRAzxKoBzI0+7ypsNAXFJ3PIijtsM9oTNV2k0tIXRWrR353SF+CkokGYWEG
y8Orr4rFJs12XmzG1J1o6FR6fsUCkmq+H/fnjUZGANntw32ie6SkUXzVWcASoGef
CxJohYQLVufZYgTP9OZ/mG5TQUaMVE1Ui1BK8NmEiC+I0LlU2+ZueYQTaeLqOdYK
ngCTOIvjY8fiVMegaZp2xmzshBHWGAU2+MeT2v03nrhKm8f7zVmC2Ft/TpFTjExE
mSiqmW5YxzRkxUb9GQ5YmHL8dnv+QTDMhl6KeW3iCVMiw+X9LyhR/wuXokWCqLMK
rRvvEApIxP73SdGvZuZAzQrr2zu3clQKt/Qpf/eHpfJtnULvxsxJPPcjOMV+KDBz
8IQbqIVDG17anXL+UHtTBBmy6e/bmocLwBE1xmiwHx5fJ+7PgYU3219ieNPadu/W
5WXskEdrsZJnZh/HuMkgStWCiWy3QXRmZvRy1FDcCEhyBVRl+rHR7y0rqYreODae
OzSLSqUZsY4mFgHIa64+UhtLNW8GxzmK4ZwjhJjuaIBV/C99ZU7Hh5q6gdUjd48c
t5T4r1Y0EoEgR5F9tfB6+ssIIGHednY5c8cPMUptUucGr51VVy8A2efejsaR2WDb
NEFOL94LmYHgpuP3hSqINaFqpfRCcFGn+0oZZ9KGrsGWyY56FrVVOr1VeT5qgm7v
MRC8pcHCSKzZq16jZUbAnm8ddx5BAFpLP8GBxjGuZ8i0lE0R7Y33D3IEWSJVz95j
dkFiP1Ss3GUErZyjefiU/rGtfzhhntwt0FsQ09I1Wn46mDxQfSkpusSAfwGuNNhH
EkaxazP+QolTkRxdKb+3zpxUKF1Zooq7DZlfTDURw685qtmmAs58f41eIBwo+XZE
ROKW2oXo12/Okc9Mm+JNenu+MC5h4egE0rizM2o87cK3Koj8Ii48OHvkPwCVTB2x
yaUYiNVThTxXAlbTGgYAta6gb22XXyoy4Azf416wLf/XrEHf2HgzD6KxKoc3RYSP
48Zc/I93YDC+B2k5z3neDfoOAXvhTcgcmqfvST90c7o6NCZ+Hgry6QZxtp8+U8pV
fmftDgEM/f7zsEmIR5Ib1664pBXx4RQYj+IlGKGtro+MKGnBe9apFZqYP9bh3gWR
yhc5E25NscFwUm6TfjXLskDKpqpCOXSSO4PbWn1I9I7QFj4bNANLkkbdwkjvn2f7
i36ecTjaOWvHt1T6wiXFUezhj0flXaS+Wr2NTOONucservE4dpAxAsBiATxt5+T7
MwI+KIrIUFhZSr4z/wTw3BGcYtIFHLL2fqfVnw+TacgcdOjNxOTtWfiaEU92YN+0
uxIvbG9MuQo4pYQdNFUHXTpI4ucADnY4kBYRseXX9kUpqsmOLtMB5pEMssxq9ww6
CxeYkSx6bdvh4s3OnqoCc0x2nUNvQF1TTo7Ajr8Pjr8m++DCdO15Tv8iOUFyM+Qo
2rkIFSag/+oWNGHMC1xktKMIgV+zllzbtI7Qhhv/+iOFtu21QzJuBKvud4hpQxGm
AZ7VK+3j3pwH5dDVjgKZaZYoh9PFma6IKT3SGhzdu8nl1bjLEF3zVpDK0nKtHICP
2T5dAOytfnf+l1HNiZaVAzvkLSMKPoJeAuNbm6nWsZbZHOm6Wph/xCU8KtY6EDGi
eZoGgiAGn7teZbNOkxPb/Hq2g3HJygWbCbi7cfgInfCSkmqlRCYAQsbsDRHwbNUc
CmmvvMUz3mZcQWpjm3nPiF3epzNHSXNkcY15yg+33LOiL34naYLLHrcpx5kjcYgW
2T+sG5r72/PvBvKfFGpOSV5hk+Sa39HuUyh/mMTW/X3Q6H3Bed5O/W9mCcWTVYuK
JbCpLBAX6+UaN2ort42PX+vmXKcjWFbJ9sV5u8rE+YtRS1q3VTB5O2qH8eRpnA2q
Ue7Qf8wHt+0iZlH3hWo7KbxCJBIOWMQUE7T0E72ItMeMX9laUJBfu1m3SVZPZkiM
HUhVedX1Ff7tApP4Yj2ILb7W1GWdeR3m6fjuR2n5C+n26yzbduReoDkdqPlsSpnc
J13KkuzXDK+9sXkpG0t6rW8jAGcpTMQWP64bKuUSUneW4BrP8WxpcoZB9OTx1Q4E
JJWfFKHY33q7+CLzJFzTzJT1xS98lqLlXx4JTLI/FGQRO9NWXPwTG8cfeFcbfUEj
RJNXMFhry178wFKIUhrj3W8dZgdlfmrKdEtt7M6RxNNludVphOdmSy1GZcjPQi8Y
D4u8lXtFtqqHxwozrTRLkj6Z7JvB3du1yE8t8YNOF9lLq2H2mzeJfnzA026HJgNN
yzp0+DoCoOH21JZ/PYEVDpmsW0jZ/AvUhVgA4GbM4LKvhzCEFPTZpcqw+ueSBHXu
hf9WI72xox9Fn/VgR4zx7/PC+J+yaSjZcwCAhVfbqdSeR/ggKZ+QjNsIEssA0fwz
f6ywor1HRq5aJbcbgL/jogJkIUa8X/JOeYy834uscQvTETYOaL+54nYqiYQV26iS
xYBObxfvsEjeYjFuaagcvzrLQh9ZnbJNhal7loi9f+oNQJGP/xKW9y6eHBs4c6AH
yk65KdpR6qW61s0OylKd9eK7uBqzF7RI7zYP6e6HRXaKXq11iiP4wZ2XHpECu2Y/
3R3ToXjeyIJBz8aeojzg/nNNNmpgTYiynd+I5vAo17oQgexOqUNJNJoZ0vpqkday
rbKB1LAoqwdNu0Udm8eOlQI3ZTyyAU0HT3wVe3zYY1vP3VZQIHCeQmvaSRNyKQ8D
VDSCEXWd6xNGc6jLbCaEM/5GNz/WmaPXS/nnQRgHsc/4YdEMBcz1jIb75fS6N2xk
P8Hs3xTcqBju7GJMpom1YolWY8F0vwmBIrUmBI6nafB05imIqVZoGQKhZ11m8GcL
ugVCTLEyaLJxSZkyo5UXw0DVKsBTVAYSkQXSnzCoqjfVrErMkFNJYHEgmM1Le3Kf
Lx2XmBLrQ5gCjndFR8b/mF4qH7cxTVtlTS015Ksfay+lCFwhAfGXtQ0N03HTtV5C
RfXSLxLr8TvLmgeheAh9REx+neDKRLUwgKSWC8Gpn8BsYui3vl3gWkAJ7TR1Sd2v
STOGUcsDnTIa3uzNgWMvZ6/9MOAiS53CN+MnQtGVWRNc+vAtiMGLTLq6f8QYa5nX
uEnyadgPuxQ0TKNgCgFvNxjWl1W0CuIAyvSwKxhIn2uNpL9misEwmSm60JYFnA1v
4g4UTYKvNXDx7LJDZpMGAeKuptUzPXH7aO9bKNRGlgeZYjObMFym2mTlYcfjZTDr
j3lvffV+PmkE3qkJdGQZ//7aUuDV61evmWL5jyLDp9QKw8UIwx0f/7GYRgEcsPHC
v0KVDiFkdcsCpOhXSNG67I6mZbjQJHlpJc/JUO7k9kq0FXQPxtTtuJoVbs1Z5E5p
NMHBa2gILrHPsVoSGT/1dzyumBaw9yOw9FtGqD+pwyf9CRrIHKyJ2jsxx6+So6TE
3+6c5v8I5olsgiAlbuSQqjM/85+PWGCvUcgV/z6MJCrQBINZeA1p0VugoUyD0RRQ
GgkT/z6wmPb0B/DJhv/XNKvBvOliPeVxo3n0lmTOBV2cgOMj5ucIbel/Nxo4T3Bx
j+EJGrZFbWl3p5I3kAUMuT0KZMRwVlId0wIvu2qFkA+ZhPYaPSQMwE7sRVRjofxP
Of3G4sjeUtxXo1fyRmRZQuTBhbbopG810chMQY0sDG6hhfinDfqgmeqF7UcfH31E
Y8Ll6oyu87nMQ7N/r8w88IVf8KytMWGxD3CrZYPgo0L81+/QoSshMm7cpnZoyR6h
XL3kK8QBEpManmcg9wO57rF/APhHVtK4mBFF2QzD7EErr6Yc3jfxoc4cWgLvVJ8w
xwTg/Y7DbE86PG9Kk1KNgewBBJ0LPTuvFEZlJL870yB6jqwDJ4D4Yk/6KGklP05L
zc6TVSw1/gXDcQgP3k2c8+kCG7IYJnJQHxaNevlWE2MQMelCZcMVnnU00G1kO11s
TrDIDb55I763lcdlyVfq6UREiMdvmPzuRD9wD/2rtacVYqWLGZEC9kpY6An+6P2J
wue8eBsrii9JOG3TvzgQIx4WhzBzEx180r/eASMtWLs0vTcaQjnPB020NE/x7m18
0c5rsSi2auPWzfGuderdewtzJAb0Glm1cYL6cCR8NX4mrhQzseFjWWey5+5hM9Rw
6JYcfPKV5KYn0V2tNBQmXkZLWx1hfup9A4xqYWDic5sAXHVCpuoDmDtmhuwM4eS3
N3+vyhAFl3jZ+Ynj2cpAcWjkTeQRTsFCZ5J8zLfzlEt6T8rp5UZQ0+4Vrjd9AP6Y
yfmzEWD3sL2XHWH/iA2GZy16WaOg8atg9uQaITV+iXkFvQjjmNrz49Grp0M0uRB7
x0O9Ez+LLCju3WYvIBlcz/gFR0pmIS1NmdSDRcf712+jeA67N04mLVRkUClnkEis
v5mlCgjjyFgkKoLQgcrRNvCRfPTsolo3hBr2YnLQiQh7d5eHND4Ve23gXmfTa74w
IY4toqlhibzmBk2Dwj/yC2uQZcjhtnjKlKK8rq1xM2l3fpjF1WF4py0xcExWcb+a
w5W4tMI1a6RolMNl2yWdwLTQwmM7BK2Are0agTce1phxruOAngaV6kOPHRII+vgA
f/tzq6B8KseftBQO3GKoZD8l38vvUcYe1zt7Sr15AK0gKiPATV+ImLdM99CO+Ng/
dHrcKqsO34WAPBLkByvOczQm4oSS0aA0tf44qYikWNBqcsWut+czRIKJQybQZijB
XRHWeryENRLehnYpe1EZfTgHipGdvGuUDJ+mJFqZyTQ8KRLPP5/RxZiJ0NdHravy
zgP/LHzWpq/KYfze9aEzvAK6bFNFCjJUO/mQ55miLjQLQA7wAFJZJ7YiJ9odacu8
gbPB4VIP0FLU91gI30TLvWebj2XObJ3cjIsC1bbUapZiQGHgCm/JgtEp5Whz+L2x
alfVYAgj84kdHfGjFb2jFlmpPQmflwS0E7K87t2v52lefL9b6wYbVOJLoxQZx2rl
IQwCUJkTaXWFAiM3ZLnRROuCsaj+8XM0vvSMNaYq1uCel3ABqbRCENVJAHfGOIH7
TebBW4enUfVu7wplYznV7v2SmILcY0+5D26XaiGnXNTL73uYtCQC7P9iI+1Cyxl+
MtuomcePO2SVZ86zvzVFiFHEJNddGa9WxwAbbAlT2ZqKr/W5idCrYEOmgtYwDnkx
YyIgSdOjei7UsmNq2EhcVPl3D6bmQcAKFhJA8NuHEVDwWl/E1PjncBmmUJYfrtK5
xtKWy4OyP8uKsF7DS0oyglq/V9Hl1w6WKMhYvuWAF6VCT/STzGjyxFXGMmzoKA2j
56OJI6q6hSbTy7wo4IFo2FRdqfxULpZmaANY0XKBwyKalKJ5D3oZk7SZIbnBHyOx
XVdvDJtEIXHZLs3j3B1Q5wkwS+2o0v1DF++VlLSPE24n+5lBOr4xh/YOmnnS2goP
aJIXKxOvz2zNCJXQ4v7cLPgCZ+F69AyV9dtRgUVzaIPOlWfihnMEUEIxjV+J9Ivc
7mQLub7VDjQCpd4OT6SZrlkyxrgmH7tZSZfuIQA12FXIVbL1GsqmEUlX5lszrnCs
5cifcUbHLQZ5Y8GcOQBpXVJcovxJbLckFjO79j52Y4mUSvXchuUdUZFKaobP3i+D
M6tVBblM5+ocDsUCoBDMVqbZ8LhUe+ldkV7RE7gAWnI4RMdeljXmybPyaPJl62Sg
Bf448aM+YfrZZd0LR0JxOWJdRzxr/n58oKFS/1kBpUQgzN1mUsHDjYqLPoYyHmzZ
2QB65Xz/nDgPSg1cdfODzIGB9magAnh9lvKeQIaoJBAo9i7BCaRi98dkFfTlO2Dv
xfrGEkXGAnXU6+jpBepDW98ZkmsuziIaMIFdUL6UJVlhE6zBR804gosBJwy7YXxq
DizgiJf9PiXpAMR47IiynQLXA9nXfH1pAVLS8nfRF3B84AlkeC3w2kEgBLAPBSL6
m7dkVXSVIgnjXbnCEoTCwP6htrZvx2q7cVGja9iIO/apXFnuYO25HKLHBnUpmHbi
GmnhNLlXSPrZsDNcMzxuaJS+8EFGjuT6MS0ZubCXQgzJbBcAU+FyCw4HivT53wQt
exG+HloyZ1+fzY/hyaSFyO9KW4yVwOeBaCzmXgNAEosjkToGVB3ZqSwIVTo7dBVo
/Jg8D6RhgZH24ePGuyKztDPRTPnirjJkyhcx3C+P7oaCnwygoUNEEjTSgUrztY7f
CEwvXTZN4OjGBxlaDs1+34HnTvoxLSc5DxH869UordzEiGL5yW46yEDc+c0UQrBB
we1RtnPeE1iRhlCg3ZXsQQTFCa2dGn+b9nRrg0laBeWKaLgOzxB6UE06yiB11gPT
jZ+3t71mbzuyk0TbRIWVbiOMxRtmPeTIY1VjJmfPk+UFH0bBbj0gNOtGOtS/xNaO
isMx3BvijW85D8+cObVlrNz1TrU89WAmApLlSvD3CNH+ZXKgrzwMK+oF/lc7mdY9
gzfIji2bmUrZYJjlhGZfeK6eSMAXXuDFOjdEK8oN9sCPxmuuGDsqB99XbB5eCrH0
aMtl+lzbQgPTgOo+DAgslfWS8+yIO0YBBksachmUdXW1nFGLrt4lpclHpA+jDvvd
VF7cS68lYptPJvedw55mEYcKsoNlPAuiHJVwNwIbXlvEiSQp7K0yMqJ+FEvpLH8j
R/mSIWZ8vKGhghAL1cOAn/yN4wIw/RjXRIRjLDKGRTygYzsMuWiiksecwsVk9Hs4
w4HnyJBAAerrStDI9+wO08Oyhp8BNvKY5KNMYdQf6ZYvIKZGC4ksiIGOx83afakp
oWfyGrCZXUy6KduKVdMChWVHoybTZzGXkcP/IQPySj4m6TFDYZPDoimsWjXZwbDz
dY4lRpJyN6FyD63QTaQP7GTz6wzOhMwNbx6VLV6mytka5uwBI5GxnOa/ixiIcxgF
9kThpyciqi9YMPCSxA5uSF2AqKqzwTA9LDHJ8LLHxZeDBI7rMNiaTH1hjczgislG
6valONP9jCdXzqM4Ze+Y5uVEyfBZI7CmXHN2kMUuzV0OK/xnO3W8oDMJOsnLKj1+
HAbZUmoOC6HvlrDlfznF7IN+5HQtKlzci1GKXw361az6LqhCGGYtDcon8m5UT1sW
PT/G0EKfFEx/s0iEVrgXhYNQ8d8M+eNx10VwJIRk8nObCjWPl7uOlnNqbOoG05fp
cWzaAm8VobZRwciCfS+cWBFpwr69lq0JXr8HvVxH02zfxINoOjIW/NEXmC2xoL4/
Toh2+As+kRDjedk4DDX26q01IPwR8nT8aUVI8O9zUo+nqffhhtoH4akESA9TCU1c
rUdeZlT9xUMN9HsyQ8MmTDOihmSJiYmBlR122IQSytTNHAXQgPWOgFVxinGi5gvc
fZXQ644Rd8MejfbmArRtY/xCaAashOnU1iw/TGTFIjPraaeZPcOGIQvuLaE40ZtY
9C1wBYM9NaojhRuz2OAKS8g8pWEAZZPrkEFfazJs7AXDH9gYTbNNJN0yl+ZKI0Rg
PxJ7mcnfRkLuLCbUp/AtOI66qqfhNhKnrbjfIqG2HQfQ4X7SywF0pDIj7kr5kWab
BtaHeEavu9EyYdi6DzSXiN15s7rKOWHEcF+voSiEzeGw/iFwe+ximuL03qQtAk5R
eCfbkktsFOlI83DX/2iNFb77DL93dcfm7Q+QvLTk69/E2Esg4KGmL+vL4lN32CbL
MWsTJ+tQvoqtVYUARdIxA8deRFczFLOjTeEbKzxvpMTcKc+z1OFplzD7sYfPamX+
CwS2tUejzpiowDr8tjt+fdB2L15Xo4M2O/Gb1rIRz+IP/riDnCRz7yMohRC+qgQb
IKSEAS7nG0ROjNfouSN1a7ik1Hdzc/YuQ4fhDFE5CXqFMUQ8umOYASRFDSzlUr0s
zQoAdsKZ6k7isJhirSYNtbSDoZrDfq5qSOExinK97+XNQqUHGskRbaYy5Yfb2Kwv
64JmpqhMSeQ+rmhAxLtIXIXk3QppkB96z7AYQbP4Mwy0xKaXmj6Pw6S5Z1SJiXKV
woJGS1DsR4wDnmU1vAROzUcow11lHzBS4v2YEnMOUcGOJxf+PAxdCByWA7UTaDaK
PMsnSYd3LTGO2DqfJ0d1VFbsvQU34QmCxR3CifxBbsHYvygKkgXAfId6foQrr3Aj
PbecxiihzICG4WMfixJKC1gfbYHGxbDRz5+Z036aHhRPWWzsuNCnCTKLVPgkRNtf
nt2IAoM8lQ/ew7Bay+WA0vAG2SomFIdZyM0KyyoKntwPcQi3R+VhmnRPQsNg02RZ
YTO/YFA54yIFFdAJLSI66l8XACpDlUgdlnNCthb0dCGUEAZy3NkFqA4clioEvoT4
x6iFbJLq7m/vR2psnts0gXi0zh0DAK9q3zXpEB+benj0i6l0YTWJHzfVFM6Tj4Wm
J2n6R3cBTMZxmOGTNaIyCrSSG6/HX0ydJqtq6I74X6BgJHlQRME4GGCESt3m8Wwi
kLB4G7GYCLeuR/mNMUVRrvertStC4OQnR9YXjdduoJwymxDNuX8YkHUcV1WLBCgS
lm+zpsndirxJ0wL85ZEca8BnFeAam5S/7pYICTPfWBxWe2TN1Sn89x51NzeXfY81
4Rhmv4bIO/0gOCqlYitSXg4pJChdoHAMBSdR5FnarbFTX94WIscBk/0fkmT3JidW
/OeEUiFmA1UuaJcxJw2kBvS4zjlFvWB/cV8TfSF/oF7kp1H0+ZRzK1L4ZZT+fMrR
w0MSfwKzsNKspqpt+bVPTncpzWoZw02FzQINnGV6b3M3JAMWRp4+C7mbbpWXVn9o
pvnosXWG5kUWAOK3Ge/gAjp0DrwfHhtP/bthXERWLT5noyMEW/1gsUetbWlax2c8
AWL+6nkI8aVGvEFCKwwFLtRZJ1+ORIfRrJ1YaiStA2G9NkHfrBDEmaLW8VvJABbX
r40Xd9nBU4WDFuU37+vM1t1m4/vRMzoCj9IYR7jyv4YAvUtxYxqqkxLPVzLcv+6b
qW4WXr2tlMJdt9UtzLN2TNd29V1wTU08nO2Li2Sh+97IEVkfiTbzyIiWrpMNd93X
znT9ozfURIAHR6mQHyHTfjdPUn/VdAYIGNP6QSTrJWIDixqOLLlOJZvK3dHj2/ZQ
4Q0+ipv3YS1KCORusJF5XIUA07wzyK0EbHOESEfx3r824OUhJ6szWeDoCNIQ6N7P
46IZh6PRKIhHJ8X0NaRpklds1VNPtU2EbUSVdvOtGJ+hGYzE9bMv+MyWiyDyLVw8
nKWWZiWlS2FfP5wi0+7RcBbR2WbWe8SkxTa8sO2//1oP9rftrijVQJssWsf7+07Q
Su5c3Bw7zz4NhGieXwkqlXwHbUkVyPz98SRT2Wr+QFMokYQVSVcA+es9/cULJBHk
fHoFJ9723AMUUMnI9W/mHSIP49wy72je84iW/uLQafrXVSr+LxuQQOHhG64aB0Ei
G778TbT/de0jUQ9sY3yqD2w/bCeoLmgnAnSfCXfhkWeIlMTc1wyqFn3HJ2oPQv5v
KJ7uKpahR5A4r7EfboPN8IbZxzSdE/AnZkJKVWFqeKDgUY/3Wz08b1h1SSaNg0pK
dV6IlI6dOkGNtQfawJm8MJYa+aFRKkT6Igocc742ZAFFJPXr6zT7EfuPPgEloyKk
GGTAStR/t9GYlBNkSFFrxUrrhJ+t+trBDBx1OROTuvndOC1tZG99Wh4xpckZy9RC
Km5cKm6K7YIE7CT67+GTfEtX0ankYleffLl42PfnIToGBtOl5xdabqdX+ZHtYPNb
eLUTIL//2nvbf3Qa+osL5D4TtO1OhQyRjQUPxc64qdWh4OtIvesad7N7RJo60Hei
Wi9fqLfGZUR5e4JANQgFlX4bA9UssAw8sTvc0kJ2ERseF/jWdM//60GqY/zoFkiv
1zmFFTvSUAP/hG8+hVi8Nyul+1OtQjyHpIuRkYXfxHp9jHtei1deQdxSm30AOauh
nM7Tss8j64+Ti95u5l8G1VQg1uBKUpht1xX0DAyQ38ZKUnB0MDfvHBteGE8zBr4W
kjUFP9wJyUX2gWHQQIIu7WvV0r8sfoEP7JZPLoI/xt84jtj/12JvDR10uE+ySA3U
0koDDM5wyoCDnF6a3WkC5ffsF11d0FcWv1H8eP81WXRiiB1tv3vpNmAZrymSBwZY
28peO2LdSUMtZ3Tucg5CgmipgxNQlXFD501K1Lq/AJkv+oDdYDjQuq8h1QCPs/iX
F7eEX4zHy1LsgjDJb5vw7gIV9YVc+zRxrRpgk3iuUlYgWA5hnrZ+aedlOAJu75Tj
AuBqFkgxbHSFLd0a0yFbKgbySbSEejzRV7TsuWLIi76Xl6UnZqn9MQce7QW+JxAD
tsGcYaVrvRFeTvmL2sxeo29kgSNO68SdJSMYQAs3Sc8unosE/GSJC+RIOM4IgYhH
TpSB54SR4DWB2BPi1YWonU+8oix+z+9K6dhw3axB+4V+iS4g3e26O/sfo/5OhqTP
c2nHS0eEXOVCg1Xv0NI9U2LHBuqHEszeYIk7zF33tp0NEVVX/9i45TYLJvMV4bVr
fbfWxkU1Cgdzeo77057ajH3hnA0H+wzjKRGJSDL+kpNTHHvbSCqCxAdS3bNu6dvw
VhgtJKz8ljXvvlR4rmTQehc+/Hu5E7Vpp0woIx1q3B/JVtKlWFfUbd1iDe+iF6SL
qlQPxsakm90ofe0l2Pz2RrJOJ35/DkIdkU79cRJEVr2DDGr6+rALHcari5yh1aXm
aRTBLqzX/V6OHxUZcNbimXTjDC9k7Arg/t2DuTDUvUdg09maWNsvEZWm6F5yPDzq
oGLAVA6Y0CaV03uwTAdpNPRj3XV5YEEIhcroDlx9kP3rlRhwWH4LYotF4LMl6F8N
N0QHhYqsPSJFKTjM8JHYUbSR1coS9rSRXlZRfO0cz4RiU3SvJkMl8CvV24DbkBqr
GwDDn+SjWMdIsvKQgjeXx56pkj42DwOe8zW31+ZvRvrOJ7IaI3jO5GMS6R+W7xFE
l8Sb7TytqNdi118a/292E0s3qQ8Y+WCn6bX46fxLolBlvfq8oWvnB/TW6GZPEUjU
92Djl6K0UYgONfBfWoqYyHX8tPlF2j3B1hh66soQpC6ZdtZWqprOSpXUQEqkATd3
mGJX8ujLIDTlk1F7qDzpZomQJ5CnYILJKi45NGkwKf6zYjJ+2SERmWRVO3z8UQjM
1TVFTNvJNZ/EdSLLwG/HWuung+dJMG3WEIjsJLLDpTAKBgq7FPxBx7fQDCj0xyEb
6bFbBHNulWPS8RAsm2PhGgrs7e6LxKKP0Qpl1Ob84FZBhBQjn7XoM7JkBR5uBPbA
OJsMkU9+gz9iwAye1j3HsaBcq2+HKAjhLkSkz/VrDJ6eYGhN17zGvT1eitiI8kYa
lXK7Jfx2fppkTyhwYWjrp+HesIkvwcz9gf827zRZwWGu5wg13kjCVdvX+YtHQdSg
JrF2GJFnXXab92zuh1qvnySBm7lxnf/A3nWDrKbkxCK027dJMV4iVdZpXPbZczMC
UtSTS7EacyodWly2V/CsMTgxW1V1wqT1cFFH30hZNpMGJPM12dCuiiQQ/P1rPF4f
+YBdWLLiz1McYof97FXrfRjf48QJnPq3LInB82IxZlQobDvk7x2gZvFtxQ5xPaZ3
AGForqAOYiaHEOHUhFHk9bE+hJkCjdcoZFNmbMJLCXkArRjRSDhLIMoWpLhdMYJS
197qLdWhUr2V7zOgwXzFWYSQ3v+4XlxaR4Qqk+I9VtmwiaCElPtqKOxfwmgrHqdI
MojcMYGWCMcuCzrmwfE6Cq9Rre3vP4wdYEGdZ01qp7Lde4rabHzXzRtLqzwgqx3h
67CJnPDORXMPzb9KQm0PFIDBU/9Xz42WdB0wqDizNreUF0iehEqS0jQ5kAOTsWTH
y5BJigElW0DVxxexPuvH6muv2gF7qiOOc8ZFSRxq3XnMrWdXnW9a9irJtckwL2YW
pO+UvDHmlfi0t+1AYJp8pso/8DQo6u2W7WPa4yDaVIof3lBxg15ya5JhjGLLY0zC
Ep4zBTVMMUxCgFcOPXrb55BQLAcuEG+s1q6eehR1WShZLfksZvDofmVVIN1RNtdp
LmIE+XixMThlwM6ANX1n+aiV/LgU2M/cVCyiEJ+yLHD0L+T8gXDv1aIpsFl6OWhr
jvaKMJhb/g+8od7Ey7MN29C9LKUwGMCr8sTSRUrr7RbakaBBmWynOPWCBltiTg3o
peSIoiCovVmwyv0kfD3C1evFJMP0CXJR9K8xH05V7OOgKf0bkDWb9LMstMMNqbMN
RvvfkkZztP3EVAgJlD8f91u9jTDCHezmLPz6dFwp/VKqCj1AbcfqXIuGWCAl8V/3
R4eFbsNTkGUnEzlom8JmDwDtkpdl5bFHSSWYQtxxNjz+7OgIckTCfa4ZgDUSzPM1
CV+rIU+X7xX460xHXEA2+v0isF3KPjYnXzk1ljhd1NzqOp1T/Q7fIeWFXNdbh8nL
BvbruF1Won0aKV0jdfYMq9Yki7UxGIESjzcedYoR3spxZuOHTFhhphcz9OkDz1P/
GuyNNvu1nbR23zLCThsRMhB3soNkEYT5tJxKuZqdF7iNHQAYyxreIfTYSUrZaTPB
xVP3ZGJkCULIjmutai8yVB7UL3r9VYzhRXCIFJFX/v1AC3+VsfSnxFqfSDfkKfR2
mk86nofO+xjw5V0sQHE0Tgry1tjVxNQqIPw/w2577RZuXfaItR+TdyIYYKxwxJvk
Mob9+q/LPHNNJEc/mBwskveehKzdEE5yATuqB0vf6xifCSy8kHuPdrsyic9/2co/
VAz9gv4kcb4yTnGpkzIpCC05cAqQtJ9z571c+DOzIC7Lbu3Hs1iJ+lRFl/UyaxWX
YNg9JvyREN4QCD1IKMrrA2MxAn2o9hfXMhD9J8dRlUHCCuAgFs90zeny51fZjfKw
KjW9KXEbLfYhB8fBJQk9oDeazCJVA+aBoaYxrggs6Gxr0FWHtimADAqCIO27G7jJ
H/SZnXr2pxj9irA3r7M0ELZWO2112Tj4Izzwla8bSr/kPHa1KMxsNWH2DjnzVI0F
jCuy2abYxr9A/p0bHV+4Is/imCul1d/MuZv1IuevGIq18J5GSwcFKCf4Y7xXvzwe
uGUlVX58RgSG9knjxios7pXnV23uwJqp8bWgqX3Cs+I/e1RMvSgAlKUkXeem+Yj+
O9uv9U75lQJoBUqS9qFdS3tn7k61uchcxPwkG5KhliI2lf1vo/ps/XFcK/+yHPqQ
kvx7Dwv2RIELYHSG2YyMBJ3FyPbBZQlaDiA3W/pZyqfQ39RMvWpSzKruQFERt+oV
q0qWBeR+IvspxyWtpcEW47E5y+kjc2x5dajAf6m+o049BbfdpJ6C1QE7VjgN8vyx
zbjVq9YM1GyzecraxknnVJ1FneEE9aaMzBeVd+7sTR+n7PH7nMRGiXTwEGXLR6UB
gMa0xCrxDV+4GpVqUCRoaMHDCEEykrokn5Rbz+sU8CPfb5/Db4LDjP10odGkXSdd
q7KJZjhC+2Obt8eoJU6YraRA8uJyY3RNKTeevaMSI1obHhqfwkUQ6PyCh+Ed0wqF
ZzzBVYRkW0SBS7crpreK+L6JyqtHTVJYFzENIleqE7DyyJu/M/vJURDKcS73SvEG
1ulqw7yHkNTgTEacgZZBEcQbnCrrjZQyR36Xzhc2jRH256MT/BsbRqZF5JMKCHD4
p+klUZF7NZheiz+999UoHEyhYqBey4OpymjgErVweerXmmlyTVYPHV/QA5uhKzN5
E14sUoIywMHIYk9PSm/unt8S5bdxbXQaSZco0N6r9cSJcpDip4tdXGPhkk1IpNLo
9sFou5qNR24gg7/D8PbE1TaKQgTn3HFTxRRUC2/Wvk9VYxymfLab5Men/QbKPvSn
j8JgZFftuUhhVmJRBIzX9XDGWA2oZJLVoh8vwJIQeH5TwAcH35R7Dl7gOmZGMqai
GnLCLKV8TNl0878aUdoS6FhP6fZxRJOKsTVTK5GUdeTN1TixM53YcT4sYrS6ZaNF
i/WMNokU7sw9bNbdFR0E49MfiQGXls+E+hVs8U3q/FT8rU3HXfaycUl7kb5SFNio
cFu5fby+2HDPWs6ebfSzk9sJ3A13txlTPlubZ6cfYzjCJN6d2nvsBIEkg6VKnIZH
gNe6OLxVGW0QaFGmRBXHH2OOZiVQIVtwGgcT2NQKII1XQISVLxUdV2lWWyPySPjB
eCdClux6HND+skV8xxl/62CqAvCiD1J0q8g/wduvsVkZ41CrhnIFBaGBp/v069+L
h7TtnPKlYWsOCsWexzQs9p51ZnTcUcFjTCtYtQDSfg0W+22oWjuBgtQAUSzj331u
dJbyzhU2bWKpScwtqIvncqwdtf8SX1PMmgnq2hvUwY+xiSrTbc+wHaZrIMIL1r1N
ZxEeB1WQePwdc5mfgjMgXcUBw5t9zGsUu+4iJMLYsV13mM/XCm2p4EkizvZHYmgW
rvGjznMm0OAJDgQbu5HdAVj3Pr7O8ijR+0DxWSJyz6wsHONbz+yUdX5ftWM1qeS9
w2tqAOzKyERlu0+d0ZPvFWlg+mYvTwnnxNBEI8J/rAmIP1zO5Lh0s3PS5wJBqC9x
CAhRXHkLq/TND3v7sY0mQly+84crAdhVP2Ut5/6rkNTVZHZ7iSixqYnStLJdUwG1
mwOt4ouHWzca7krlZ8azlCJ6Kfc+yZGvIxFTqAxBKfzIKlPiXjm00V/E73uM14Vh
oNfN/Oj9cPO21tgU1UzhkTafDB91EyFxi1/ETZ0uJ6MHwZ9ufcRu4q0IAVo/WcsM
yMwWNm+tBW6BQDDyLEuM74Uw383hpPJB9q5f0RdAEo+oeIHnGbexHS7b8YvQniFX
rjfzAgf1zaPH64YPmhX0pw13IbnOXKG1CMd6kkJWWR9SFafxEQuvEoJdyPSvzB6N
XvMPDJuecyPqnt23+eSE/MqYUKbD5/OrbjpC1bQeOygKGvLgOtTs/IXGmWZoH71J
gh7ALA3IWc+OkQwdwbO1jT4HVW21ZSNNJWmwDDxvkao8n9WoQBm9lVfkBo5GxdaD
qoxI46sslsawIsxt8FQsCRjgvX11GY31IdqLgLiXi/1yA7HKQkU1Kw+3RRTo+ZQg
owHCR0eJFw7EO9yJ9wDP5TivMla9+h8NzzM0Jmmi2mDvgrCurFR8FbmaiLRR1HpM
OaDBn63HpNg6lsv0pPhNKbg2b+10lhndPgcejK5o+hiaUKZ0x9GZ4zKPJBXaMu9y
oT09dYwM5nVpvhJQA4tkNR8DrXRTP5W8gZpo1kCitILjL2QQiDdUPJQGCT4KdOcv
UUKMONspDs8CILA9TiohyLM0BAU8ELSTuM9gaRM5KAiHe4+pDGKMpnX3C4J9tgWu
10TslrhWkFOfnyljBR1hVsQQY6gaic6oO6xptLhI7EusjdGfGnPRm1oQ4U/4L8jv
uYNRKp7tnhT1FDeNkmHLy7KqgyJ8PY9peX/6ag/GWn5HugFln21cXTaLDGNDkX32
zK1cBMaBpUpgCjU6RY1nfxIZ7ErkkyX894VwojGBfrHIPi3f1V1DOnEAsBUrz41e
yMVpk0NrTHWneoE5ch1DtE9QcY8jhc85zKASju3hItNxxwV/TWch6+2etwNwCDDQ
7LtlKzeMg1F8DQ8/vro/nFcCUNYlBj3BHRALtd5jWnyNKp/a5QLuosAMuv/ez4e2
AMnoGIdlQvXYBgXxNuNNmfOFtnwNX1VkSZxaOnjS1h9bjZYnPTpTdPa/6beSQuxO
HgxYR31JAphH0ZngmhgsmVSJkXzxG8p1orMN8e4HuGg/AinvVLv/1L/dcSQ8OXxX
lAMHLQ091u3NCSP0set0Sg3tRBAm0v8+oRk2D6Zj6+iKSnsyr3Go4mcJkn1NhAfS
lcrS+JLca1J25YuWfE46lugkolVO+fPEu0WSrPwxU/aa86bM44y10yYR7irkANi9
CrnlSoUIcKz1qoLEmF/9G/020ZaeY9WMlFgl4uRPYKfyS+rd79OfRyO7GxO9Ri+l
h+anRfIFIL+WP7ZwtED5WwuIi90Q9HcdHULbnFnhZQovl5cgYVHIZvvUz51Q9/hv
LFAgmTEAtkQD//GQA4K/7bCLOacNul2OgL701drVlZQBx4pB5fY1ATM/0yFNNphb
OM9ci22VfPILJSLs5oNOLmKwnBFAKR7E0Mp0e+Aq78L5WsZ5d1qYmkCT4LTerwM5
Qha4NtYCo8F34QJgzNE89/zPu7A57YBmqKew4x6Nmy4iXRmYfd7TX9D0siNd9D8j
pT8r8Zg4bLdfU1fSD3g04ZFNSw4ZxFqW+y77n+jzZsreIqnE7IFpQD7ELf8Qih6s
asMKaG9hlHr2YQS82HUvilh48Sf+6cXz6E0n7nYfJ+4Gut/oLO6YkuFFWblUmX4i
CheJ2eh4yV9NevaMAr1BYMYlhg9BnMjISr3k8a3eylNdxOAfQsN1oOKHSwwZL69s
Py8lfzxNTzPmSJZYL1wScKjL/yD1JMFKiSoG9cNrMzodJ1uqi9OoXZanROYabyEw
eXU1xaPqXnQxf/nG7qn33xl20UJLedsrPoTiL5MIGre5dm0XmAjPJ7CWtCiiJFFg
tiWHPdzpDt9JkRuUFaQrl3lUIz+A5yoyN7vWyzukouKwhKPSZ880j/L4A4FxvEsB
e3EyvuBRy3gwod1nSW/Rl48sHJ3F/BbUN4/UeobqiQiyGKf1PDHdx+8k8vxVSies
w1pb+smZB/smaw1J3CagfjHQD1NsUqhFkKwpCafoJu/Kh0o8Va6CuyR6aiQbdUZb
aR9hOmrF0n1cXmTi2G7rEqnoQSeBcvur2BescIH1iIYTbS2AadSPc6VvMmXUVaAo
F6fGtr6MKG8tZ79WzmkEFkbc69037eX84qSXT5a6or1su9PwXO7WgywjIGiFjY1j
mZkeJc2t1S0m/SW8i6o17QrHtYDtUKpfR2Qm1cbmBVTjphm4YC2pn5yldRpqsVB5
3Ja09tTwOCenn/UqXchhYhyJYw9EOhPOOCyRnz+GOJb6u0IX7b/wa68q9qpUKWFj
u4GsC8hOZHWU/YWm2BGVbF/07GCQj0iD99DJXEkwaC29ejQT6JfwfkVrTe0E7Miu
20HeuEb1RUFA0YKX1dJCp1YRsIlTuvOtJRTRlFFRk1EqZri1kkhjbCZE1+c69uDU
MaB2NcU8KCZ3EIKyQeOICTVcbiOm7sD1bEvozUsyZ33EMsuer1pfU4jf3kvhEWcB
M6C4jiNA6EcfqIpKoc/sUVy795akiE4Ht1rPMovRjtIWdem0fODDkekvYKJOLojR
ne6HhCzrrorIb8eFS6nrN4WhDD3UZEe9HuNe1tt8untbcJMCMp1hhKp5zTHZ7ABh
gh1vFjhWYlx2E0d+CKV6TFonPCjBSAZNr4abX3+UKcZqVOqyCGlJE6ZoiydbVY1f
mLtUVPykdZgzgf7FQH7cI1S50gHbmigTTKPiLCOY89jtFbVv973U/7m8JLDklEAc
RaQ103qJN0Oulilk1QmDLsnAhNJywLIBMeNPOFNdVwVCTXWhkMEURcQfafcpJA7X
k6/dXAvU4Fq2to4uCjV4dFLwS0U1qTozSfJu0Z87Ack1LcjeBK8ZNjDVU1EtmhKh
kEiKGH3q5c+J8yy7cNqek99uLCKVw4DzPQVZGKzmqxEKPFdspUp4/od0pjQJYB0X
FnsskVt9gWKCC4Y8k9EymKm9Q7lmKHKnsUaSuP8VtTLRcU9haIEIVCPwbJx6+yZN
NzMM2dLvrpN6X+4V89norUzaTGwAryejHuscrc7QkGhWNXUYJi+lGoh2+XaNrvRO
tmicMUx5C/X+kU8gTvaTwZUGaAeJQh3orJqxHGJr4sZekqw7sH/GGuqc282Hf26a
0EPwUZNkmYt0J57D3hLAP2q0vUeogQGNdrJ+8Q+oB4/ulBxolpPpzcheEv1aXPug
ijKtfWwaTnewo4dxGtfZpm3TrkLsPxnX0V+0WFqi0JMOkh6fXHIwxb+AW5TRgylf
vimQqpS8rC2bTn08kfuehe97d/10L6BZcONdeuZEIYeAAH2J9thyARYbizn+yVAQ
+IlD85ocnCX1p8h9iKDqA1mP28O3lclU/M2ZChy2bAZY41A1sqa7PKl5vWtYnBxV
eUFu5KE8Ih85WYdBjbVBphvlHmFGB1yBL1Lp8oxU9o0Zpbj6nVvznqKFH28stIfX
TZdaZO4Q2GRWIlDN71mQxNbPaM1l2F0Ma8G36hi5A3nsaRsIjll9xuW6aV28/JPG
jpImCxf/oV8gRSEMmlCzHvqBOIUXvS8QM1eznUzVt+Mtc3NuXbNavGZrny8RlsUO
n7dLLCLhx25zjSYrL2wQgQEsBYTuyd/tah+eyV5K+8hy7LwGsdnssmiX8+f15iGN
qCHxTPD/OCA8bTk3E2N7wwTEIwLTAq6PRTiM4JhG/hh3qBCtFptIzTbJ4yADMpku
m/MpQueb9v810fUrop0VkqEtSSHkhYCpNrTtvpH3BAsWMDNlmSv9RmbpcW2dz1Dw
XzcGQxLrsbqOvm3UyBpwQHSCazfJ6xfZDfcyTeqkrIRuAvG3wzx0OeL0HQiAtXeN
z3n5OxY4ZX0sAcB+oczZEBks+8dyFirMt40qFOvcGk4wvR1yJHzWgVuy9Xi9zcNx
YFdN/EDtllUr1M0DPjso/nGeLh4Mw+D7qjZBSxiY131c9ZfgaaUv9cWuP4TxjLL2
9mQcI4jtcGEeKv3ipBAg2+5V0JwNUBgAu7Xl9NVMc/VxhbHJmC/9yPDj73nizvXs
x+AplXTFm2/+1F22xvZ0qj5xcmQgp1kERZ/a+jhPGTHLb+zdGgz/8k8XuwRC1XUH
JZTCHF+VbaQt3H54hZPLeeZ850w5en/fyo0+3N6fZ1VA8I03bSiE+yDVwHmCFaG1
/ksSq2ujyyg4BxD+I2NLVYJXQpD2GyrANJXGkwUYgljE0Ndq3sexdP+3Veo7EqDe
kvgnacPh9qPPW/8wzlv8bfLHUIpyLY+nZbDRxajyaUMzYAE2R1wd1BdcPi1bNw+S
fsTmg8T+Z037NBH++5BuOmDirug4v17bIMEGiPOPZud11au1RNk9XWMNnrqAy/5Y
v4+bBeGDE5j8TFmx2rx98Y6XcGAbq44woPVD7h8uCWcA7u15KekB+iAnBzoLzVo8
O5a3+nNzl6NwnNX/f+0mUEnWQQH2RX0kG5IrFAUNvnh6uLkZO6QdI8g6Xodd3NLY
F0Sd0NYLWxAujJX0JfoCrDWMWe6sL+Gpr6qEukldxyAjk+LqXgw7as27bf5iVOmQ
OWXwzCYI3WXrPhMTB4qpZjmfjpghA1ByI8zZxpJG0EycOfN4xfeP5BVuWo5sFlKm
bkBbcHAjvI7XF86N5a+zC5VWysCAyWpnpbayRMCVr8TP8sRlkxswKtWpZosPEEGd
Z3wzBY97uy98P47UczWaGBeZd8ZAdqS+amGpNCyeHp9zB+Yp+FrzwMVYDPug0Bbo
Z0+z8qm1WrLgDrz9eR1+fQ==
`pragma protect end_protected
