// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Z0OH1N8BjVmS6xihUY4N3WQ6F4V1o0tmJOIXsdt0e8jZxauiR/xZhOeBGsmbTync
K3SYMq7A4UjYPRqc8DQDHCtImufOx4ZSeqMjfoYSB4nHAelCA4+aH9Xm5VpOnEAE
Fvf4mUM8hvS7ywc7IRKnG1UsvGhOQeGbDbSe3y+cEQs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17456)
orRIV7TOQBFtfHeKSOnJz1/ADgLbiS5z+sJQ8tIJth0z/mspiEdOhFSTRitJfJTX
Be10QTVzmlxv3+Ovat4F2jMjrOjk01KB0FExTBhPbId9vggk4VpzptJJDSWc9Z/F
BahDQCMxeivB58c0jNdec0K0oW+rc46FIqnIsnlrDh8mMZS5feidsCWsFfz232mG
jxdTC3j8BgAZDacmJKv+fmANBxtjZ0MCkyZinsuCdPtpMWogRd+6lk9zzhaPvNiD
T4gwM4JLmRgKVJXcqMnayyFYB2vWWBSC6+IsNNnnNqqwjN9NC225bOWIkurZUN1o
WW18MGrjP1H4+mBoVOgZudzJh4mlwIiUp7Md98642h7/eYjlrv8q75n8LJlijcXe
tYVyKrGe5f3PWvF7QIgQHv0mNUix3tnKdzjWfqJ+QqZYreu/ch0A6vFmqvOCdJ10
QXzZV7ZVgWYXBxoE5ktYaedQW19CpP1peuLVOXkLCBTliGq7K2inIgZdT/qXoJ27
VjL41J+09cYk7Y1Vgxzv4r+yE6ikDo156D2jDI8xv6kyY4atcD4nM7Bsg9y3tH2u
dMlOvpy5/SIpHFRoMgpnvJlGGq/WjgreVwrWTcxO+AKCr4O76iWFSdTyNMN1dHCB
sxvX3p/eYGPnGtfw9JYuEitPazGMxero1LArgkj1Ad+QNfHg7u68Hg5JR8DpokYq
w9zh2dcXs/Fw45swXxF5C7EzIOkxUMeRQhLrNidKQpt9a/HtOns/OkMCoEJVyr4I
6PvQtL/m43DTuzRsiCaEh9+IM5RpKACUhIo4ba8T7e985M/3y+bbpUrFDPkeyjyZ
RTj7mJqDw33EHS/O6IFFMLqzGM76Vscth0oQgdIJVWXSFbGMHOZJczkzZGykifeJ
4Hf3Itbb5FzpkkDo757WNqgYxmWcybzlw84aRvPSflEv4r30qp24Qqv18Qtc9mos
XhRThWn/FLbG5UvbSJaehIL6/myZlC9HE37+4J+3dC2bfSFNw/lm/DU0CZ7hlYoG
oEbO1Gj/Rq7awQJKNLg0cx1OXN+omQNIaIMHSEubTpNPqdiAdxcqVej3v+bfElNB
bIFby+Pj+jiuS6ann3ifxmh0rRy0gwaQwSAP8P4eup4n7Ry9H+X8jMtboyHBG2IG
1NPcQPYRncfcxVMWy0PTTnl8KCMqAcbao8BFFIukJAqQTujuN//qrQocsNU+yHmx
QLBTrCLu7kk4w+xFuYIXFfDx4dclkDPUwedry1OozPvycKE9YLQoqlDs7EMpuH3K
cZ8Q5RVEUvP26mOEUJa9IOVl2Jj0bisREZBcZT9Awuq6CJ08jVijThY4u/V2wTZj
hVQOpd2Dxb4GwrwdVd/P34qcB259WIUIWbO4viV7/yYzEZTqFHLFHSte4gxLHTEZ
B3YLtv/wsk44uwHiXKkOWntPLfXIrR3unCmK1KUacohYaUxB9pKSWV9OoFYuskVm
0mO5+HS4gzRb/rZgQ3ghhlqdplB2YlDaLUH9WkR8sL8Y7TEQZt3MW5hQJJYdueZ5
/BpPwTrGMavcaHd7ZLzZ47DguiZE1zzWK821g4zwtqe0+t5/TA/Ii99Cr0N5HaEc
FIAhkJzyY9hs6XrualrE/8kXjKb7zxFf1n2LtUmkWdqgDy5hUuO3GzCesowuSO0T
/QDgrLHJJp22KxLLLE5G1wtNLaD4rnoWXTrzN/mpS5sNybrc/e8U/+U+n3IG8hcF
wsuxrvAq6RjTf0JIIcTiwh7DzPEDMz25VgGOx9LqH9M6n2XEhah2RWk86UongvJu
MH7jR+Kc3cfym2/nPTjPwvlzMFV802gUvNKLfOUD1kB9b1kStRINnXmS49O+HE+R
W5/dtC1NRS2s4mL6/zgceI+Y4V8nP197BtK07RZKoiynSWJk3DWhdYRA0ZpxFEm4
Eaea9kRkP1N+8cFUEuKJxdIE3sXhKFkBLAyudEt27ZNN9kpEcOQ3uMPjCZhhzMEx
wRoYdN3qhgiSiDIk+LYIgJED6zA+QM6BFjNRPTolUxafsB2KCkFP3hBrvscKYvHC
XFD6jy39eesDNIBQxJ4GnIWjOg5mbn/KuFEQ0fRfCkgpCN3xMcmFC5Ldxq7LgCn6
q3mFF8DbedxvpOz9mU0ovnA7gAwNm5CRfAop08qw5kot8/CKWH5k0W2tFxkApwFl
IAUU10tkvcBuJLqfJxZqIHaBXOv9WeFyx4IjTNBI4oiXQ6UVitSTgbHW9vhp0Q58
h9EMN6SWIphYaEwp37feABm7qPlCkERb69o2IJZ9BHSOfa5HcF10FMaSLam4vm1B
kOQqUVjZKqLI14Pk1/tbogitSmslgLRWjZYoowag9vBIJMy/er8fhkSrh3q3rV76
FSBdHiL9aRMY7c69UPutNT1twmmD1UZ/myhR/pNzMaBa3JDOIy6/ottdsBmD00Ms
K9tsSJvg3WCAb1ESORDIL7osWbrFyfwjsLsBylWM1ONtEy8GoYQuDGAIB7QeRTpK
AoP8wI8bt+olMaLrxjkrLOekR3awcd0pN/SEIB/XgY+Nr0V107T2UYDpcyt3xQMf
QvIsadIr+kh5qvoWNLdllONR+NuEdQqwcMjzT3uuCN/G69ppV9ntFU7iBvG0usPZ
GMkDcpkohjBfj36A2SuQmtb8WGm/DBVeK7DHd+3p0nwJTKD9pPT73SbvUfnko/Eu
OldHwXx4vIloqMmETaR8GQeThVDDvVXYKXJmplNCax1u1PJnZQHTPktlRiS4HBaw
iN1/7fWc3HMhfYKqs5dPij0+IwhwNrlYwagZzmkkurd2DYUYKelrsjZOkwGdG2Oh
c5Xd0duLEzccV4/BTVYuuuEvw7nBRh413C0uQC0TU6MB+f4tFBTcLxdXZO+/kL5k
+dhLP0k7qKMBt8Gv8ZMaYb2mqCzvPkc7LSgSR6HPNFduzZErK3iQHpLvLsyPW+iw
oF5HF82N0jaagQ5xrtyNp/JahuFOopsidzy+hHJkGOJ6jYUq7FOPf7gydqDuoE5x
Eb+RUTzePEW3cOOv+Jf4wh6+BKrZh9yTScAH2TJhFY0nOj6yH91aW+p3jG26N2ri
/fUZv2yKNKitasuycRUPr9iQdJNfUOgO3bnMkesLQgqiychsO3NZ3yByBh/JQFhm
40xLtkFj7jWOita/F5MN5lM1XmyDEMEg581cQZfV4MuiIVxxB9vjc11OV4ElmPYZ
Jy04Gwv2z4QykLuWEqyhU/9zOvNxjU7Uk4ScZqm9GdH8nsugD4GJA2rBcBzt3duj
DXcgVE6jmHeHB60UgM5F/ETtXfBgyDkJ89Z3wK81dQM0d2tfy3qYKNVrTBd91hoG
hGoJKgkScOJQ3Wr4AJEiTJFx/+LNqIp7fqi9D2LInW5j+rbL2z6nt83UdvJ9SiVu
kSXSzupqpSjq2EwPem6WjHJ+typ4Bzk+/vfK+3uu0SjQj/cUKG4R/09eATApvWKq
/zAAJUe3PwOMXpPhZ+VvOJmjgoI+qlsfEEVUFMXW2gDQVuLtqi1D1gsTO+X5v0G9
dSTv5GNM9XEnuCq2loBh3dEjHDIWcxerIyxf+sjmfcpXU7dONGvvEY2JIBDAIX5m
EBlym3cZQT0uW/39L7jSAiq0K74rrpqQfgD9695zC8cycToWu6johI4hEb51+4mi
B+XuuCuw5stEsAifXqhNi2wYw0EYo9hhpZFW6B6FlZuhzLRDKj8YFM0N9aV2M5j9
sdZbkxv409lG6wWJxAdgGbtK2yMxyD8UnJC9c/xnatEw4++fWvNGAI5Cf0RFozM9
xgSqHkFocqR2fdX11TpVnpSgxabzYSDt2XR0ck87TCBMoy+j3SIQU/0x5PEsvcLh
0IYALENz3BMYA67zh6yrUWRtn4uuSaufX0+rKTfL8Exa8BkzQiY8k/wlWpJ9caiR
PXGy1nm+zOw0nzWQtx6WXD234/e/1toxwAVdu1aGsSFePo/ExViummdVpGd8a772
28Kvf63H/kpQr7ZwiXWsA6E81zzPOm0wjBjzhbV7H7e2vdEX0jXXIgaYM07kcN5t
kETrciOl1ROOpADDYMBy8/FxY5dwEGGLy/SKusMj9NRgLYoQiM/Xaio8di1zSj3H
dISeDjJaZLiuEq6CkZHbWP0TRqMYM9N3+O+/vGg9VDovK39EA+3p2k4rS3djqbe8
GOFF5cKpJayhEcQU8ejbRR9oLqw/lvnrAyGMDi3hm71crm2Db4LcM0b8/k/HueKK
NqV+3n4UeT48LJEkPzJt5jKPnZUZSMQfvFGLO+91NKj2tcmKYbLDC/v/+VwegZgU
M6s11Z2bSOLCb2o4o8j0pfFeHUkx1VHjULNHdE6a2O5F3QZd4SRorBvpdyvOaxM5
pARcGXMXZg+6glPYUlL2N8LmGNQndjgkRBZxcTPyxXna0ZfTuF1wDVhf3KqGmIFb
iYScMMrXoSj3owOxoOQrKVHbTKV7UQgFdivoqtA+FNny316UkWA8MnBDWDGTy1Ia
0g/PpPLVmnunBYjkEtRBVoi/dW0qYN84lxuqsSZXBHAHSoZL7p7lsE449VxioHrs
vdWf9s89wbzy4/GQShp0LJxMSOQezyIniFrdmKvtXoHeiSq7i/SVvwmc/bft6mnM
PVubmIJiyrxE4o3mkLpOtykc2FRjQ08gtpxBG2V3bNQvt4fThaC9t1AmgfvFPmjb
IIDzz1EiSY39xRLfnt/fg7RHkKjOuRBUaqtXHDikPhf4qGpW41hOp+RAtRITKT+n
2jcYaBkkOueDlcUado5uN1pxsDFQaiGurDr4bbKy9UVAGOXB0K+X8XEqfYIxwU58
dT2L3HhzMQQnt6gsYgRqAU7xjxFc4oTcbGRdxD/m3cj/zD+pHUwiy6xi/xW3yEit
egg0ms6BW5smFTYHcAp5bq7kVKa9jtAogQsYl61L9DR7Cb+QIF2yzCxmrBROj7z6
KXbVhkNlH0jvkMkcb2KZkvS3+Gd8GS0R3SrBRJSdJss89xWwYHM6f29Uzqxgqtgw
q4KlE1DWZWoZWy+tAzS9DidWc8Q0AKGDgvhbUC0fF2+hqsG1j81jV+EaVWR/1+uz
EBIE3AZchHuSWV+5l6VZSgszPCIzeWr4zo98PKnbPhiy125BVJgyDeI8to0gIVxR
KXsojvZgQtrkvShUMesXMrnM/Rh9FWxb5omQZmmxnM/ANHHpSymbvlfgVRPx38dJ
d88mhBv2dVLdXJ6NdD8dzwV8ovtY3NzVz+9TaRTEQuqjr65VoUZXMpqAPwJtZo9z
DGv27y3ErI7lMZvu7+uu9ArD+ynJngCHcjU9jEiCwEz1t9c8vQujbN5FIhHhsKZH
nTkliVxbGaUJEyc6VJCLON9yL7k7p435HkYUXVxLfzLynz4ixUOxyi5es2+f9pJn
4z0Ehn6FjHJckchTMkTPRZn5YJel9sOPlMJOj9t4+ldbCGEILGGlbCNHF72JyUPb
/ax9IQtUD4MkohQwPERcvlT2Fe0BUOgKFfegimg/LBGODI1Z6t4NxaQmud+y/TCB
6kTRcZiuAlUPnHL4E/gYyjw07OsstbIKkzDVn0CzcuUfD/lA1+/d59FejjDxjm7R
P+yoBxPmiZw0/C0YE9UUV9IcYGjlIci5uLRWWHCdnlyozPxwXQiYIt4OkU9QJubr
fMJIMJ4QXgdxPtma07B8yrx9wV/PlFCfwuuxNKzBQkqvZ+pCeDRoYisN4gaTyo8V
ilQCFZQQrqB4FKwxG9JN8KJhMbhQXHQ1wUxShl/2QR5azBqHPFCvck9swou5SZs1
XAhEicDtNRpWitfhOr66Iw+qubmnE9NJFeaL9zqt9YnKeUvmv2kPcGmNGauH1imd
VdOM5ll+B7xoStxojkWxZiATpkoKaNjp/Xhmg0+dF5H7OdGyRRvw7CTKcuAq4C67
P/gNc4oKbB+Fs66mrBjMgP/YZBxeD5euSdijZW6AhkOlO5cxbDW7OFkQsTdpY4rS
I28U+mYxxCpiz8MudNJDM2bNtreXNv+FdDpXbNQqP5I86CehTtr1hz9ZVOD2IWmd
YMEWtGgviNXlpyyonpV2rZd5HKPAz7iiTVy3e2zo6Npv/RwJYYEwwkHU81VZ3+9o
7p6RRPMwnU21ASeWX8YUEMLXI1l9jLGq0Eqf1rFrJcD2gE7trROS7SIZIM4K/wnv
1z7ikx/fVCFr+Hxs6em77u1KSIMiOofYcRIHB2lC20MFfxtSrhGY9fzSPV52Olok
nlxW6jWShzjXfYXyOY4oA9JZUW9FUyf7FUAWUMTgi90LzTi0w0mNWQRmTBZ31IJF
ztW/rwj5+r0fr/gEePt6ZE7V9JOzG3fT7Y07R0wDwPspwbGHFH9sJiuSwJkRTBkY
po0W24UgcsJAbSEFhCNp6x63tXJhUDJCwmJ/Og8Am+5OtjLIebNEabFQAAymlzn+
NRCoQj8X6hdqAsUPysEWWwFbGB3KKuUp3CqALwu744vPMJBrClkvNWaFW4qVaE17
YXqdlLkuvDNbAM7dVMIp5gTCz7HdHn6wGNZe4yo2YZVLZ7wlsg9AAilg0RrXZfH0
DfKV2eli5jgtuHMVrycN0kiKwTCzsmIlGJcyTeXr1tA6k1RaQJ91GsVojqj2Jbli
RWdh+O9wfPj/skjuk1UHy/aSY3khtROqdWVDC++EgGN6R1IfgDS1KoBoS+p8HFAG
n6oelsIX/fdc2VuWmeUYBIZQPBL7VzUkL27HAVQSvBVr48AQ16zTrvoM9gbkDNT1
mor1B7OaGRwEJRM3YpJE7C+KczpRLFWrTy3cAKqkYHoZPGD5kPIRvksfUNPjZx1U
shhTuPVYMYmCOhkEzVGdT7Xecylicu4ebx5jQd3LmvLVkRXkm1PlLqxoFgwOf7Bm
uvCp+2QJKW9lzjydv4B/PRcn2+MEs4vZ5naJ0SNGnNJKQOOnsaZx/YyjTYObK/QZ
FtVybc3h2zw9Y1dHckJ2M3R7GT2N2ePyjHhAxDG/cIGQzyzm7jixR3VfuwmaYMI8
5f3uPX+CyI8PXGCoM6cMNLOQDqGPgIojVXuJFgKwyEcdQi0Sef8LV4VHGhIqwX2+
zNBzQ/2pgDYRAnPtFiFJrL1WQu2QegUPu4wcOZ3KvF2Ctpimkf+o+gSyx8QsFHSa
ytLk+XXk026urHOGyRbUXyR0CUSepKL5BETVUU68YOBK/PhesTbz+KvImZVZZdzK
hzRK66AnxOjh63loqxVHIpmLPZx5wUNzmMKkZyCtZmOexF9b00BZJB+VWHTPOSjD
gkOsBZW2Ru0OtzEmWSnnA8RC6PMHTZKbzpI+APyhOv/5dQ2NdDxxs0LZY6EGJ2Lm
sdsXz+MBwFbjZV41GnWSujbv1szGhJdTnz1XlSsJC+G/24TD79Ul8NwDmSbCKoid
LIlGkc5CpBa4HDJUUYSid4tACFtPu4PVtoPdH3CUAl4UgqgPGV4BjPdSyuBEGXpL
Bk4zcs0q2BL+J4FpB7Scj7vbtMCm+cX+oMU/9PAbowXZ9mRC2KUOGuqFhwE71zGe
fgrJaoSlAr5lQVHsMSHI/+CP3na+pyHDz6JKWS8IZnxOzJ9WGblFz97syxGAJ77/
YkuvI2KjiEDWk93mRsYFFJ1snoKK5ZHGmmT0sjOr4WbVrgU31DJS9PEmJwsK0/bp
XvraJVU+DPZ4w0kAKnPRgnC2MygQueA7RiIllsbDjwlJQR5irBIMu2H/xtLwfRQP
SUnTE+HGYfRv7PKDCIg9Hu2+jcYZ0XEATTgyHyQsDr4i9STceZq0Z9xOtd6ncagx
a4aSrWtEQ/7QHc3W40sp7OGPuXbeKAYxfevjmCjEbyW4Y6nnag2N+fCXQSxE949x
qRy4jFb95qi0MsJOiTogPlWeJIg2wF4b2lpovJ5z7zXmqzz6Zduo6ga2vV4YKtbB
uAKD5EOdR2q6EmCnQ7UwrLXXXz49zK5EuJATyY3mEMnr7yG16iJRZr3yYpdgk+mk
t5bWJG4l+6bl97BFTOAQNpZXLDUZ1vwBhWXe2jj36jgrWNQcxCiqZMWN7JE0+IqK
cbAICWFRScCPewF0wLR50eoGfDV4j6VCtQWuebWrEyh0Krz8c3U+fa8CoPP5X/by
3tOL8jg04YLWRKpXs8PQ57ycexsIGOL5zkQ87R+e+E36F/drYIaULh3CCzo68beG
93+yEVJJBFKwYnl91z6O6JWALOvSLRGaw2HuITnKtytahLlch2ApdrQ0JZyroWkk
tSf6JUuLw8ohIWbLwD7N9GrxgecCZXhpInZu6vk7b21PeHReRicJC92uq2o1W/RB
/XNyGxuilylJLtl3n5M3k0vkjpBWpamj1Mw+qhA5sy4eCKvdY0mEWHF9/uLNOe3j
jCUN8d2MPktqM5lTQpQoSgKCgGzKe8NPtEbbFt+gfCAE9j7b9c+p7fD6KIg2/yub
4lclZWycPyToXUaT5u6w1UKIlCPW6lLTJA7xjvk89sv+MaYKyjdt53viRk3nnJlg
5xMSZHP+5agsVYJfIxz2DK9LsF+HQkuN2Yr4aEQFDs3rsyw10inAYQaakweY6uBk
wbe20HM77wCnaqmaaFDQYhd9NMZj4vg8QV9Na6fiVzVC3A8SvT9ZrlxJsO3Nuk9Z
2acUMFSEiQJeaYCywBLZeJQqkjUx+rtBwp2iSu5zFs+r28Y724UHzvyVHlCoOMyX
UBC1x3KED1Ivwwb9sPEbbA9vGwNfWzL/0KyqmJsnKfupn4YlH/8XTkfTnh7Hnlze
U24P36/pqx94MwBL8HLc3QrUvN7tBLzXeh/8lNnB8vEKeBKqKzF6uSLG+sj4uou2
DtMIxgdWZnoCQGRzmTyii27nIeDIb6vMd4I7d+LPmUj3xRB2TmBzMpMbtbSMbvx4
IalvBiRX1wgFFH1uk7y48XJdPTvfLeHWmm639jit70gIrDSJR3YQoZ6Gm6PVLdPD
ArMtjXiZNm3vE79IKd5+FSW6EPAgy8SAMYu9PtVvRNaYul37PsnqthHMxC0fZSka
zUZZU/qPXqMbagf0KU88TqQi9ZAfkZq5bu43lrTOhAeqJUHszZ9agFnbaYt21CSu
Z1i3TEChHHPH0N9a6dWuCeM3h8fqM6L+7l8qm9WoSv9iURgYsEbXNWnMMmfnSANq
16SLLBQND1o8U2PY0aFr8MA+8QlJxhL9oZ2J6/yoHRxHZjRFvGunEDW7ch98nG7W
MNbyaFdKFLnrt8nf/ih1ymGwI9y2WyTATf5bsidtac7HSXNklNNIeh34/7SZRheT
N01a7MkJIj9337HpuV0qPzLpNZDqH9rO7w2VmxSjQLKDfVUqqRXhzPrYt0gKVBjJ
kkT3je53TDRfdBU9GVXW7QrKDAnrHHFSKLD/AXPuHTB7AJUDYfjdSHwSr7tTotoA
oEsOJdBE35/pZa21msb5kDZzwnE1T85kQKvpxOXlkFdOr/jpiJblYQTenNLnUGq1
NexHXCT0C+Yw4RzvPF6YDupR9QJ8F+MCxAW3Xfot8GfG3imzVH45xSlO2LX1xMIz
+iBbRWH1TShvvMG9PmxTW/5edC+23jiGEz2AGGjsv9aV9aj99GP+kcl17o+KeSvv
Kjz/q8RNq02luOUxfMsKPMsB80piPMd3v9iusS8H/BLYft66nzlyDRXuP2mT1Os4
4mg1FDT+hdlB8sHuRwIgEVRXwpYWuvoVzbYbkGTeHM4GnAvDmdLhOD4rxw6J0X8X
3EzugbkJyxldRdp1ECuMvK3ylbolRZanY4safdktJcl1ZXriATeXWjSjTn3Xj4xz
+vS/nAWKReZyBUNr+4TjT2HWdVWxBEazaTu3MVmMgEQE1+JpgEfHnhT/idEzpsYM
UJlB7S221eVdYA9/2otFgIFCgfy5StQtR7Pmbv0MSA6SG/w3IMu5/E5fgo+l1bcm
bhEwqcJ5NC9tNioqdTNC4bTmiFCsB1JPPWaEHK0Ai9r4NyY+RvM46HcCeSl9LeTe
2LO+UH8vdLkP22vBtJJS8rUthWJdvpmDNt8OeMtAt8tTm13m6+8sDeKmvLoA3Fve
wf/rAD68MkqhxYJNrAhjE11eNlA0a6m6g125HOGYb6r1rz1m0HdgzwLDaKWiaPen
Y0HvyXB82+pAfOrW/9hK9n3NRZ3/xnM/EBHa91l/9+t5W/xZy4vGwQLjokRFTb3u
eRNUFi2Ld0zm49634Tg3F9KYjRxFlsri+i7JEWIHrQ+tgWOjmJawp5HV82S9a9oP
RMD3+f4/XWvIJ2j1kFrMZWcNBIcmia4q8pEVy/o3LeYSDXZTwWVFouuHnXbAoRNF
RPypGSx3E0oLCs7iLYU7CrZr7qe4Gtn9cvmxQKCwVabGWGRIOXxszDUkFSL8VMuM
unKiqI1c1rP12gmZ1ZwP7HK3BKRfw1xXe8WQwJp+Vn0ywV/sVbGTR0G0M0C418MP
sEUsSzxrrRWR3gwiJbC61+3KS7P/HJv2WeUeRaCtObEsWJmgvoRsBbOgz42Uzbli
1xd1SXPVu4CTvIBs7m56+dHJeQyv4ptBEOCSPonhmF+JP7vPQXfuuZ1bgq288lYo
uB71vZX/sSUv6CMJ12qvbWmOEIHZ7Yqfs4vnMQ77FM/E+x3wDfL9dj9DRUq6fvgZ
pIfjlzdP1tS8HZl3//0GX13PxrFqNtJl5DgW1+psdQnpvYGw2tOQeRE9m7BhUhf+
xR3TvVbwbW8prK6oQ0+iDix0EgNyH1AJNeQ9tGmtyhDkn3qgp1/PIFpYugMezFe7
5L2wbiB9ew6YX//XlI62XtVRdVF3D4Z/CzYq2GpFTGy2wNkfnJT0uPvhTLeOFTz6
wZL4Q9cogbIOpHeuwFRuL2ou0+fuKzIOp3fijBApPgyOVA2XopPheTCX7WpHV4YG
gYhFlis0eE5EaYOqvGA9tcHxLPvLwKCNvn2pMd8KxkpaG142tF/db8hzStYlvgEM
fXRzr9n80hmeGn47/FQ+D0aNdLul2UE7r1npvD1DyWnuDKg/XgCd3Y+GMzNLz8Pm
038qaUojH3DfYVyiQspfJQ8jABmJKvU6p3Vj6ct05ekTAPD3ZGfdGCrDRSE+pyQN
ajwPaKiY85VABInI22ncfB4d6y6o468rS/w4RHQ+F+4sAEHq+/NDElBN2u0ygN1P
dmLR34kWwUQioTj5230RhAUPaEWq+Oqna9oyiEKmQQUt44UN0LCdRG/0VU2R+k9h
Mr95moAhTEUZIKC82rJQt1kbwIXrM+C5/S4nR2HD+h8pvvaQ6drw1GnBpzA52RAI
paGwP865sAom4RaNJZrmzeVSbnFpG9g9RTnH/mCPxESJRAegvqeJS1s7v8bB5PWs
z48Ze1LBj9vY/ZzttU8ShVd+6zqEKrNGYKBbmy7S/zAKMbFFQDRTiGUDaaBMR/MY
MceVCKUT6rFGsIei1h4Y0gZiGyeRD5c4RKpT5SDS6MGozB6MXS5e2Uc8IkICG0ga
PoYdHtdtw/iYp1Z4NOjunpTSRw6y8KU4eO3iQuYn8PhQWV43SJoJVylJCJ/cqDMP
bPOE/ScIgPKXeIFAV1eHExeQqnejb9xE6Ah6Q1GZPe/gmNPW4qBmVELUWT9AxXgf
JEyMk8wjZouX0ATKrmxktLbuhhmYVgKJ920uG3udgrUi0Azrtks7KuTvtFu0E+Ti
YjYOdq/13IEWXvtsVgYhjy4lk/6K4JNXpg7SlIQp5sKR6Sf8ODAUqvMqPXAb/re2
fd3psAN6X3z2ExBXf91U39waoaq0P+h0jKEBwDyC4KqA+3uOXibK5fLsC/AJDFKO
Z2ESpWGBZS9tEd2b5z31IBIJooqgXQxPHrLPXb0qII0B33GT4dWsNBEe4qKJPYVt
6kwAhTRm63ppLiM/t9kudgAeKoJ+1cbt9qdyvQF6uS+79RsbgZjREfCis5Cs6nIK
VQcofe6sHbjOpFrKEGaEsrrsQAn2nchxxM4wxXU7AO7wtdJNLf2H6zBCyL50chBe
sHgCstqZJNCan4IKUPH1e72ZJHWwFqkKS5sx+27IWdW3WOFOR1Jax67SHMLIOkit
jLyHNTNZR7DKr0EMMxDSs3IdJTckzrfRpSOgjgC4d0kLWhL8WJAo+FdFMxd0T9m6
ukaqGpBCE69MPwpHFHLXIKjzSbzzSBg9jcDbmauuEdjT7U4E6h/KrIgGt2j6DI1Q
cb6b/w2/7yf7nO6TxFvQ/Zz/AtmQ2gBwFLtyonvvdovQkwBsZXmK0vHow35zFdJS
BLjK7u7hnWGaR2sg7YLFFnRBEE67ieqgOAgcn4iNtE34JuBlocFTBTlZVSt4NJ5Q
NR6GQwRtFhpt/uRXrG4/7nhXe8UP70dgw6heIK+2G5+iBTMU5ZarT6JV2uhJXv4T
YH6R9Lr8TLphK6X48tXWqMOCucvHNVAAG0kInZRy6xfRRHM1orbfTDpD2i6SM6Gh
MFuebWOYGfMkVDqkZxxomL4lfH3hsOrSi5E5BVZ+A+EaHqkW5YFqH3WpxppwtFq7
RO1IzETXR55/Qg2VtxCB+dSjd59v/N6V4E7qm7t6qtraBC6C9nxXSrSc1NBRDddI
blKjuF2iaY6n0MfAg+NTYqsDZg0MGb3CjEe+HOYC+sARtNm9k5SkzJ1BUYNrguby
u8lufQl0XF8+X8jJexpCwNOAzkQ8jB88JDVxiWo+cXEue8bEguL0Hi9zc8uA6iUF
tAO49diGJQXCcKR9kH6cNPN/mJleEqzU3bKZdiixS80jmKIaFG33NMhtBwZUY3Vb
dFhVeq0SuOyN2jM6xvWq4ThHWyIXqShKHKwxZDgLtF6/ffh0n+W3XI9lgATzmvwO
VOtwyXlJjN8HASAcR1K8IE6+nwdI3GahQ5S+vgetVnlx3i/v6CK7j8dYujwnFwIV
2qvYrHh25TPLbkYWqYzcKxyvqxXaonJAuWHzKogYOAjypNqum7KsDLSPjo6MRhh9
UYTTa+MLDXLCUkQfzWlGbxzDXix+qH8Yopr+ZSviouw4+xh+kxRqS0NaBCBUpvGl
b1y+D+AdIoHSC3PWW7JiePBx0hmNm3/zqW/Mo8kv3I28kZsmad3XwqYvCQSl8gRC
GtGOtafx7rx8N9ikFsElGKexaYqD2fOWQYCOg7fRK6kgW7+4Piug3fTc0MUacUlS
4eh/HIW/apUMkU1AfZTRjdq9/nI45KsDAlQU+J9g+A+cBGsd9nF02UhavhrXKYiZ
tbR4KlgIzwl58DE0P8l2iyWSH695IJSgjHdFubN7Mf8sFlK+/GoGxYhXQE0kO4qh
/VNc6e/IPr5JkTIOYWwph0swmS7PTWIqRF70QqZs7UxWkthQHwQu4g2pzv80ZaYV
AYzBkXKhpDj0Neu4AX7c1g5XOxPVjdjBi7WDKhLzU28tHgz4cHkxraOE1Zr29k5U
OZ0GuBImrt7DwxEoLPEP2VhplkaMjr5Ka2QG8m390WpVfGy/O9yUnKeUVZJHCY6a
sJtZX+ZAPa4AXlBpmCqjSJP32P6zUsq0+fKsiJ4VF+pKwIMDA6wu9hEjCUOfBt8e
r3j+Kr7Y8XM5SVmWtMQA5CZygJdXU5O2wxURPA5RLhXkml6jqVdx3mjnjPCrmu+1
FAgrSRR3NoJbxxgDanDrtTIN5yMn5Ky2C0q6KYILDzBSS1YPx7xejcygWmZTnw6c
OZbID/oA7Fj0EqUN7QMiZIRZRIovdyfAUsCXAKCUMmi60ljEiO6IzsPYAWdb9V+a
LAC71S3niB76N54PXzH9DL2tVF8BURtXfLRIp1gXwgR7eyVe2IAyOVSE7UHhPr33
FJCu9JpcGFJRhw7pxtWg55qxm/KCuW3KhGk+5ZUwrDFbzL/QRjSnbLiAV1KSczo/
IUTyk8Vlz203qoYhD16modb8du3u1fN4qmkdgUskX+iPW9GeDNZROpNSC8yY6uLs
0mhrsJqP41j6Lyi4u8H23Qi1oIRZF/Pxs4M/E8661GU6nF2WMF7ulU7q37ylrR7c
ljTykPPvGrVboNXMAbsrFRcB4a5Q+ZoZDzoPw4IjbwKpxhOaODbdnx+ctkMpxcRN
JGHuy+XSav6Y9t1ezOQ4+kUeJ2O3DqO4tLbLaD16xQclKdVYmrf/BXg/tOCfzeqW
LDy7dUkegzNDJ9hoHENtdcThj+ax/Fa1NrDjYl9nQ9gO9uQPPiawEdth5Kadg5HY
UcrI+8bGE1ZzeHE9zwdY5kU77c3MXNyLrR/zxat6Tsq7vWuI/HfozgCHjb28j9PR
3AHzy7y+L2U7zuJSGTcuNj70MKibJcj/yg23oTXpYY0mGNryO1S3f3Ff6y1DRoHZ
uOM9hGNGN9qf3bg3Y9GDldYi65NyP+yu5czFycFDHiJG+aaZRIqtc+4gxETRhft8
zE4B+PfzRexUSaJg/fjFyRjGt+kQMjWYXgKVs8QeFV9+YxVt8CWYzYZJ0yj7o++z
KFJDWuleLTeALagwUr8H2wYptDNgAl3SyKZR4YXXekJhq0Ysb1pV5bT+YnIdvPcN
336XkNma6Z1HFqHTWxWM2yp9poe5hZHT+8BaSytKWYB3dAC3wz1N4yOefac7yDJ5
OQq6hYqliWU29tslMWNp/T5xSfvs/UIFBbck5yYH0MvsRTZ1tewRlFnFG8rK/S7X
4gC/NSmDE9Ue7aTPYaXoqJ267X0HQqfndWicFgwScf07RImT3oEC6hJtnaxPkifB
vm8PFmPVr9QvCrW2UXqv6wqeiliHsRxAXShpGoPksDOzdCLUycMnK+upMVH9RsRF
0Fin6WXxS9BVk2SiwZ4Q7CqWrA4u6sOCVluirwN+h7IzjUs+h2LhvQ4aI63sZIco
sIPpTaDBt1Ldw1GGUaFagVWTR7b1rt0YwgmqpS40tUdtmQO92xAkSoaLoVhgwqZc
JhbGBafpf+Fv4iqrH34xwrsmQEVLmoE1lavj6uKXjUZNGF8CpBrMtSB1EZkZHgPU
V1MvT7AvNUStpW38dTQAYgZhz9kMUXoGz2uWZtH5oIf7rS6GYEyiAK8Q0jiuM6wv
/utYoAOd6kAblmBVvbbfAPxu0vD78MV9DCeGg0LbA9Y84Xs8LpttSAt3GfdYbSIo
gsJMSj/wNNPS4z+74RkI8FsaG3Gcmvkf20jumO1snLcf/DX9giytQVm962o/z0Du
3Qax5LHTo9wVkdWZjfo4HBV06zz+JGS66OmpmphyD+KOoZJRjVzZTD0hVeAEGcSW
hUojTG57LPQ7NPiINbkdkZg6DYSYYsvVkqd/gNxxVuHb6nVUs+ZMev3IWnhfg/CS
j301+ikYXyaiwMjyYAZd4fGogg8tRVFjsuVd88q8PyGpdoMYquw+lIhAVRZFYbhi
Xdvpy4fZouhs1HiOupsS6/fBKMKOu4MrETSbs+doL+QoCZhZU0jov3y+d/i/f+3X
2y8scOrjnWih0/MD5mXXfSvUvVBpl2Tsv5q8CN77PUkNUVbk1zIt/yvF4wwAXQED
Dcb3TVcn9AY1jEApDbQLGo/pccHoNn/7NXQsOUDq6OBoAStGUOmt9LH3cSC9Iely
0YlspDfoXEdjmvpZGjrn8numU+9ZYnobrMNPlRIheLfmgJd+i1fF5i0pDpCeoq2N
SfPBJtNqX64kS5WU6LtQTmL7A+GVuihxqlAmjsOPHVF/gjcZPrW8QHxhtHR7rT/8
TT3SOj9d1+1eUbT3bg40X1N9iH8i5f1PW6M3O8cOOpttNAeehfe936Uvu+B0s3Lb
nSdWA5zGeW0FVTAKUz4YyulxvRVptOM7vdpePNldaTH00St0Rz+/cATjFYxX5Swv
ljGm10I47r6sNATwwdQcj968IviQT3+Da5roYqqNBaua6O/kuAgz3tg6gACYzwrZ
tYhvX258wbkoZAS2vX3PsiRWwdaV9H2vLjpI6K2FHIUiH28xH++IgLWeRXTnUlqp
yCRC6nDI33rkZeOsZpUoRE8XEkGzYW6RaNIYCrF5eSSb1SkAK716oWChiCTCiAm7
LKPHLErXFzOmw8/vqrOvngEL30xJ2eNUA2A9w7hxUMWVhrO7lZYYA7BTXNRTqGwk
Fe6Uvy/QUNgJB9DCKwjyV5rHrQcB//aCad8F3SQqvLNzeExnpcd55NqIXdKI8S0w
DZDmhGYt3oDR0oowgd6rmpXNql5RvgxE5iHbT+5Gm+CdLm+wEVk1KWEesiyqFrfo
bC1ec0mK46hbrVcE3BqFGckKhwVT9mg+8qwl9VyhN985/u+K/9CVFcTzhNvEuXCj
BXzAZIzriXEhMzM+mxtvejmE3PKSnko6BoyQncaBcmJOX1RlFZYu+8WmRsCPNCLb
1wUFVY5tYOm/rAU6271diRWdu0d2+gDG+S90wM83TwYqjIM4aUVo+uSF+rjg+6UN
m0GaDy8dkDF6+yhrFfQv24qWM+zJoJiYfa2Tu6BpZryswDUescfEAlo6vY3+u0a3
9DRjYlD5MEm54Tu9cRRQbeg3TRnVug+o+HouJvmjieB0O7JieoGtAZY0ZxcZup/g
BLhJQuAUIU1IHeGLxagQFJXBu+6UIluRy6wwy3GF4Mz8x7S711h2NMWme2Xwahpz
+vSer2++zrkX8t8brozV6YpwHh0JHU5IWq27PDopfguPplywILTkCJulrA0+MCiu
GxK2WhAdOpE4mOl1JpiwFkubNNCVacup3ghdn4eMXomMTXHOT9klWyjtZhFgBCz1
x1Cqc8TC/n62YzP2c0QQ2QXrcMAjouA0OZ3RXvnVoKvw0rzHDnHLOgY53Yor2a2B
utzxoBrcjID9yyQnvToNaafsYsPKTWwQgtElt0/Ez7v10SsA0x8liY/jNgQFFV2z
lCwMtcRI6A0in+v9B8KzZ8hBWs537x3mP/El/96yB/G8G1erIMa/CeL+iCIE+z55
O2jxgBd3t43Z6yA78AbBEhr+STqpGIAHgWq7yFgFIW27s5UNOaIn/RIy95aApK93
wTWcySRz+06u4oOtngbpaPBhE3lIfS/lvgPEtvjsv5IxM8/yuu650rik5PzAgZPv
HNNjCUyCiNsrwZnOESGj9W8KqsgyZ7Ptb/p9eD2CGPMq3Q6BS/9ph3TNRjWiK2ZE
khzonppK7FzcnPY8yN1QUhcRG0cSZFJ93QTGoq6LrsGRmi5R9tsyynuS/UEj0EFU
AqA9LWL5PjKYtG/G9t097ywSkgvxj/4g4HWrZHCx+bOFEq4URc765L8WwrSYojUo
sqmDi02PXMVChcPXlCj1kYxyFDDVS+BrIPkTwVdS/V+QBUSSDcfIEubuB1sdSrao
5ojAd23pE+ObbWGiKRQGEFNeUWNyw6ZEwVmhX0yiYiNX8ucgLiQvkEKJK10vWa9S
9EPrEkNNy5XXJLrACICZa3GXIo3c5hwrVhDxf54L6akaWywSLKeY0mpx5y1uMJHR
fpZo4EzsDFsY01rN/zYk3p1AVRu3Fw/w9Ao50Gayq0wOnvh8a16eEfnwTNaH92Qc
T+DQBiALUScSV1acu+eTV9I9aEZb1x3cahp2k2nqwNqg/E7xo8WOZBQFEwaKXQUX
/ezixjjodVtdmD05vlJSTD3A3XFhn0+z2m2N/+i9hsxcGvBPDcnk/lJtW8Ej2Cp3
FppKtc3Gg3vre03r9yafloY+n7IldRbaDkegmujVRchWOJoH6kB46p17LZAkKGc9
qcZ2FPEtQjrBGBq9eN1sGBlN7RrqH41eagK5tM6KydqFGN0BK8Vj1QE/n5yqB2+r
Hz+2pzV15g+AjQeSmlvA+lu0/ZGo4tAfdh5QybpOVSvLVL7x53ShItM749jMBGnb
CGNVz7z3adTFOFx4L382XvnFGKOSVn4DVbhPdDkoC9pwboGDXK5aT/HU6D4hwd/3
mmQeeUUIDHtWa6qF6DvYx3KxtMAXx6t+ZvLo/8v09a4xDw/W19q+UtKFIClNhdtW
2jvlMqQEia34itE/Aeclvks1uUT3GqshRc9l6TCMIgh2HhqHs9uPN+BybjMzVgtM
5KE0QkPiphHOFyv4xkzXT4eqwCsiJB7hRGvYD06eq92un5a/JJQ0XrWtoNz7Bp9O
MnHuEETcDWDmk8JfhWVNA90hEwj7ZGUGwt2dvZWrOfSBOjc3rvmmHgq9rWh9/Y98
4AHIEAITEzDxJl8osybtVAVrN+mXuVR0mxZQXRSdnzJYVVncqwXdCW6qCKLJ8wA0
uJSzPN98eJBGG7ZGriE2Cc/VK4tnPI1GzNSpbpL6NGUcSa6eHVbuoX8bXKPQ6DQC
C3XWCbwjFfZhX5xCGYQ9vd2oXWa6fm5WHJhYwgNdoKAxVJJWqeyLt5x4WIxFpAws
TFunAMay7SCwsYdPzAIBjbarlVK2KNqNJRWzl8BxTn5KgNQUOJNUuKY6shKTLLew
Xx/M9qRf8IHNfxTjJ3IyjOaZEc4jTh6zmZHrhq6Dc/NOAHULFXWv/0ALJOR1pXmR
brNtkRNVV1vz7axI4TGb0pKxrQ2UEmEAKu0puQbDeqC51u6+9xDkpPTLV8+nhEGd
zly2a/IN8uxVThw66VxBXLvzhKNr1zdfm1Ok2BflO8S+D30cZm7GDAYSAcYn/GKc
svez42uPBiqAs7NFrRS6//PsAA2C/6k39EBjl7rNodup6b41YvxUnb6QzUfK6qMs
LxBQ1uq237cj/1cRvei/fxZS4xnOGBULZEQ/bv1y7+MrJbnfnASgC1HZaBJx734T
/1Z5fUZFJA3J1bMY8famWkXlxDYrx1x27HmTo7SlwkM+XnU9kc2DKvYS2mXeHIfb
m7bwmm3tdEkwCF0dygzCGPUMKAMMzcyj1U4dO00+G/07+OwarsItU0C/+v02Y+20
Xogcd/U8LZrteLCqSGg2J+axqiujjlgnPG29YXQXX8cHezrPKKaz8uqctR1pn8Jz
bbW34K/FHhDHxKUYhEDH8ao26Ug62Xk9UGOTAP+GpnsmN1r8x+gRyFmGQDRxqqnq
WvP0TSYgZTERPaeJ38Z02zm0c3F1hXWKz23IZzkdCDD3H9KX7MysLVow2DbnyBGm
nvhlv0A9GvDmRntjc28V0zCauKt+PavUmE8Khq7OLBvXAiMgL/VfyAebhHOojIyE
fE17B0dY6zfh5wIspVgwRXmStiQCtFk7w/01SWSeuG85FVN1kKtolle6GTKeK4xS
0bl0a5Gzup7RpXO1smV4f2mcNVf39/h2E3fb+1SjY4TCAGlzXqNTnBg/sIJlqHRD
BVuKKGh6UGr/dkQRKih5pYAn/FR0uf447IW+DxVdeP8iyxU3rjrEKxLoKaLCBQ/5
3gAR/2acpx6NZG8IPwGJM20VHNdnitIV6woPZUSqHdoVK6bMooPfWOpbnUyptwaZ
ZUG6KmX0GmwzV0bv4bEz20ElHppdleltDMO8p63aRbsWDZryBmmCZiGVoCHHwBYb
sQE2W1DTkRCZZA9/UygG8wXDSdJBh0FosNjsrq+whvUtEDTe93CsfUm9LcqnmaJ4
1zxY8fuEgLHATOuWNzRqh58AIjnzoFkJXcNrr9RQOOhCC431p8I6YlM61m5WuF0e
9Dhe/t9MkXVuMBiRNof0D4HG/aQt3T8WirliEeeLmArewB0NG6Nprc2wF/oqAgHb
u8pFdPwVZt17lwM17vfnxoFzmH7TY9PayMVOCXxjYzHO0RAdKRqUAycWa2Me/LOo
omZ/CE70/m5Enbbw7pNDkKcAKyvFYfpB8CdzO0D9mB4MQSVgmR6mEcXPlC3H0zJN
CX2E6B9uhf8rGzmn5axm8Qn512puOPokiRIicJE92supy55/m/YD6wQ5+pLwA9dI
7JZuhgYn27qaOjLLVJqzgxQWmPtHhtiPE7a8qmMVFOODr2m24EZTVJMtS9SZNR5/
oow2qvmcsyhJ1Qbfvlrh7L9iyqxBq2Mm1myhFkOJUVJxlJzziLqfGY9cXPjLG/zL
KWy+QMhEm3TJrrtYm1qK13gMmNz5EqpEjVqPn2YMLYJLR+Qb2yO/xiVan/aNUzFF
HYytEkWFRjPKr73nbyu5XHpZYOihjdilPTMJxA+FzUFFStkEM2IUq8Tclio1MqED
hJEehYF/+2i4FmWMqVR5GReOrLOxVusQUhTAZOe+beXIDoQ704G1p5xdKnpeiZWY
y8CGoU4eSwv7zhRuMYHzaGyAFe18QxH9lCkEXvI1FpPFWQXET9xOKou14ApQvbl5
1e+NPHnoJe+3EKwV6EEgZ9vUdsUHDsXmcWrrDLemUAUYyBzNx1V5hzWPGK4Z+dP2
xENwigYTbiEnZbEJc7MEqStoMMgPPrsILGAyYiSXsCowvvCPuAICRguazdWy4ltc
h6CFcILQs+UjuUqaE/QWTa5fHv7mCxhYzKD0ZXvkKT4txoNK35Ib8XrQZ5GoX+Nn
As703mEsYqD1jYMAMGWhZcUqVFlEj9gPk5S0ficx8Oy3ABAY6YaTnYZfyiW5IZnB
pEW4/GXFJABfTp4IIrocbvj9WwNvXO2Q4jMoxQLPv79wr28VPEawa7akWbc6cf0R
mVVK/ejCL9CW7bmIckKeuS2f7j9kyWCpUGAaZLvcCFOFDLSis4U6ECqhYYJt9w92
1rV7QBOq/U3GKLPS6Gzimqq5kiEMD9dyMHLSOXEXnfS8GfaJwxnwYQgLvXfSFWHp
RGxDHm8My1c3sY9y3YZC/n0/912nYxut2bEyvUxDB33gy2ZUDLzRZ0gV9NEYVqas
aUBSI5I+7amCKIV9LAJecptnKrmBX5Jk4G+AAijJRsK5xcD6sSf8x0zptNaWILf6
T62rpDaTLEnXOIwDXFj7TbhPAGq1BkBVPu1d0pTC/bSy0WjxNxaHes6xBLufjhxW
ivKYFVgqpUZp/8aukD4POuNHrT78qJqHNA9DdXZVqe3PnI6MVcttbahgAqiO30Yd
syrFJYc1Vvi/z1RA1C0glWYc6A9Rysqtf+MsqPxhmtBUT55dfRy4eZU+SLSELIQZ
WXeZGTZOmIfSM1zvsWQ1Z1E/NtNrbJCGrGAb1ArXY8wS/HVgtgZU+8GiKHs8OsX5
PBfKM094IVnB3T5weUdVn3wUirVLp/jyJptLuATJimHwF7CIXmLv4c/I1gFtBzPQ
YJY1aAfcmap392TZ0HiZmV8pSE+1xaqFTpt4ryFK8tB7ge8zV/2PSz5mwWEdFsMQ
fEcS57Djyy2v7gFhpONEUkZTn5SWOB2MclUi4dJSuQojfktp1nYIRpyt7CrJ6y4M
tEZmkymMuH7hzzku8CVgdYmr6PkY8s3IT+JpbaWrjNXXlAqgd5stNzJ2f9+DjYQP
lzovKeqYjDiU7sq1TOHh3f+VaQr3mQ1E7/jh0dqha5CsISCHWtwfZghkM2wlRKT5
q+9ykmnYoSYrssvzen2ZbbJ0RQnj4IQW3VK9IesFHRRoI49BFkTb1NXBEWmEziSQ
N0rkp/atxyi6JehNKLc4H8fMPTa1v2Qdt0Wb4oQq26KgOIB2q0BONJnQoOV5nKQ3
D5typdMzMx/FZ7MUroPuPrXXB7LH9Hlswl0zhwwQK2AWfSzbWTAiD/ldLsVr/JU6
fjuqPFsHYxmgLfPCB3Jm2lNJLsnEWC9cOkhmZsBPyXE9l4JkPR3/XqG1yf/bHFzb
mz/eQqZXuoCF5YM0nOaSCt3FKdtcww2Q/atn0b2ghxP5aLNUI6D2G4+5ZpL1A/be
P9EN5FlGiPR1EZYZcwYp1WHzuGKA8JvFY/2Cea/aShW6pOGoj4Dw04Ju+0zUF1S3
6q0H+hykLoExmiDQbGA6ekr++DUTbZO0bKp4XhP7sG1I1h7jmrQZ5Ka1shG3Sfot
Awdn/43mSDnttC+ONqS7iU1dKyGzo2mkzOdJNORHHDrGPOH/8epzpcOBNtz+tB0G
wTNCl6VMDPCK/ZWNGFXNT+UHJbK6CnLm3R6G1YSGPOJJOXWM5mX+pen6h06zXFlU
dr+/A/GOX4GWenuw7+FnpUG5nqrMPOqrFJl7H5SiFdrkl2Jv/3nDJQBWpUzZNbj/
93RQPkFXqveQD4v2inHUKGHSW8J99Pah3AcIh1QadOdR/9Xi3k7R06x9zoR9TQIn
cEyBPpsGNd9JvDH/VBBy6YAAz1Yn9jTx1kuv3MGV5q8Dyw60bS/zu66QgLP5zwpa
N6L69obiCnTz62y5UgPcZ7wwWDD8IgXcczgbqBcDl8T8mXVMSxxZjID+giaVFGOE
uci9DuEMu1Y4mzeWdx5KRFtBmwL8Hyp9uKlRgGimiQSSDYOc4Qm+LkqbY0glxQgy
4z9mTDNRHMVetwEeNyHjDFGsT6GEPWw4RjSP6biDNi7tdYD2BO9AaIGiYANeX7FZ
4gZtDuT+RMvb+dg8TxhY/VgD6nvjMTeaXylUfS7mDHjQb2qbIvMIFMDiFN0r3VAI
nd1BhN2mhyeUpwftbrXeq9Se79JzNvz2XcHmPgIfHmIKKsQJI/WWVveCEQwyGOuy
snGJhWvcqvQUo8MgQNrkkn++nyCbOJnng41ZmJg4lw/2yKiu20uRZGgjBbe7vMvx
jW/lSXE+hMQphrMroTWndHUJNuuVN4ZHz659TH6ddI9ZI5XgN/G9VdnykurCtzWO
BrZLQaWnstq/9MBbDlZ9dnGZpwOJ8N2BIuxtM1toA3IjnMsYwCFmeFWQfjrmD43L
i49RV6AVOAWwfp0dq+D/TDvNvOCbPOWtFpMoSW2qw/O8Pgq+o4wkSN9ZBaVZKiWy
e3eT5Sq/Ra693gjJ2o0a3dBtNtvVm7Fq+0rjiEG6USXc45GI08WeIYf20p10gDMt
89mwPpQ5keN/VvYkViJz8ie3Taf8cq1WBzs1/3YK/KDBREvxTEVV0PSuAeDEWw45
6GAmqB0YE5rDFGsqEaQ59qNrtHz9QgW1RKBLIAIH+5bhatXDS8v3YovxcKonPxJx
rpEWn/faFnT0IOI0Y5PnyYowSGFD7JitJTInuFAKGxLAIzwgGU/ouLe9DZwC9bMT
TV0DLVkNOuOlhDW6ubH0FabblADQlRJ5rP+mBmtIaqEqnRbqWvGecB1Q8foTidqO
jA+3sqUBS/jwDpLuoZ1aNpa6WpxxjmEAxZ+/QHbknQABRGexYkqZE8FKU2clLQIh
CvOQe6xaIC3XBWY+A8+tfsaoHNDg9pf+JKw5GMcOIhWCikVu4+ze7W4whKm0YdCQ
+tzpGPWbqlBpDvypGNxf0glp6szU6RmMERIoKinOiRcDagLKbZ5y1l+xAzzRPz/0
2OHWxXi5U2OQ6qcwMsZbdCuciEs2aXaKyFS3BIbLDLxhhc7tKGSmLJQLaV0V5s3n
PYau7WIw2kSF5KZuINs3lBxECm64ugCpp/yiRVPGokBOPdJpqv8+/w3ZHz1mJYAJ
KHOCZc8ItN8A55iKrA82T17JjAstQuGXap5qoR9BpKhZRo6AxOjmDFlaqlydeOAi
zxYMA+azAvFd+qWvbSg86Xp2PX4/mA6m1u2uSVe+HbM=
`pragma protect end_protected
