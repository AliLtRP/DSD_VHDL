// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MiquLJ+Q7maRvTo5efKmh7OfHo94ori+PX1Co1VRABXhJWhj1GAkWnnbIypdaS5D
nlJnj9gLlQVmkseJkiJZbVe7+A5kMtq9bJv5BPpXE6NeYFF2iSGqNv9u6taXLeI5
835j1MWND+1edgLt1BCpMBIFluMa+d2hSaReTKC8guk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 41792)
ssUnfBgl47Qnon7Kk+IYP4udvDX+DKaIeSk9Q96Oqea4CCwcAUwpfy4XRPEwhnBL
6KnWXteFJh6wqBsOeg2K5uh5bwNRxtnyFIW2CByQM1BdA+rV57DSp8Iln0/B+BXI
o043OgQPxMCN0TpkMOTEBjJj7m0bUbH/nLZoXVDs2Pf3PHJjaqt9OVAKyElJHetC
L9u76JHz9AGtQotaojNhewH82mzEH0jbe397ZpaoZ/Y513eaQKEPmaNAoNDXcz5i
B2Q4lYJ83cpKbVpk9k7Wkp5yj85y4YpezoVcFkRxVnqmukfR8eUaAvlRjfQfGAu+
vLsI79V+6Uv9hAvPIXZXshn4YB8EZIs8Kx69FsKvpa2Dr9cOPt+ZpmTBFXrTOCvs
ArIKFAH9xMRfruxrYu6k7NR4GiIXi5vzVkDIMjvRzfR27D7YBPRCLsmEQBwtx0k8
cUV8ZtPy9uy0STdYuAfOAcNYzadoXK48ds+DJdfYlPJkrrMNV90d0TBCNCkxBCbj
PZVINV2u55j5cJO/pnA/+8FJLbjsNRQSTiO9NIIaVkIeh6dHzmzXQR8EDieeIUXJ
i87fAfPRO8BkijGu4cFohaSyNCJJTis8lS8WI29JdR5F6lEXVGpDsP+fZLjl4Pb0
J1sXLXZbvGM5lHc7Yd4Rz7eTELoE6V4pF6qTgEmWCHeKTm3M2iWhaAmRxNuy7sF0
gLihoC2uJXNzd74+A2wZn7LAR60+et7/Ea2eF9gSjFxCwXL7uIUEBnXt1CHL3TIM
aFFGKtoLiWJpwczr8C9wAoR7t09ZzCfZACZ9h2zccBl1s8ga2OgZXeLX/+UMK0aP
/KJfLEvCaWcmsHI7i3SH0E++I4zBLbBldgf1R9br/EyDlDbDOuftBmFi5BDByBDq
6V0RCShP/xJTG3pxyI2AV7MN8OPAV/XnV0LowbmHzt63XPTb2JBKuBPyw1p+4h9S
1apLwQlamXRvG7iRAOGD/9iMIG/uMCtHtOLuCaZHlbwNUeBUlnfIfe9qadyX7AA4
ayH0GvQBBSFEcMOvrv6uybJ62W/U0EDfLIW6lm9QVme1vcEECtWHq2Zu9UAQ+Yn3
1HvJBb281wfqmDFhRiq3E5FZdqcfQw7SwyIO0eoYtqCba3iBlGcjCIj6Im4Q3xb6
OHUeHAiHPt4uaggVUmAKLYD+W7AlYjj7UoH2Uv/2AODFKBVzcSaHzwiJjgwS7kZf
xQ5+ubbPfAw2ufGpJsS9yChYU3yEpUUIkZL6VxqNnknC/X7Wv1dH0HUb4DQ7BRIc
0IRC70f+8dZYDdI8jff4/w49mckmJFlok6So7KYhAhlSrl0Vq2g2LaJawVRbfD+K
wEMSQwv7cfFpca/pqleBvGzw5MmUdk5sc8bVynylF66+BX1VFN6Xyl3uJGADYH9j
Vv90gfAiUjvbSG8gx6VYI8Ft6g5Xqzwr/ZunBsU8HGb9hh5lxDaAXdAcvWNa9w84
egHM+Cg3ap2NjaNB1Xa5kj6Vh51UE56XwG6Fi/LacoCO6gBw1sFu8d47/wb7CYlQ
zRWQP85bZPbjxhaKMVas4YNmDjkA4LQjJ0ZdeF1LZUaZ1vdPUIRrA8DiUYJxif2E
VQtiWL3aHlcHw9JtCOCact9NFindM5at3GnFr/aWVBy+nu3fD9PxTtlc8SActtFo
9UZI0xZzsxOnT/qSxKF7iiO1sefYXTAMC+1sq4NgsWDzI3TPU217KLM9xbMrVKN+
KhiVoqKi4cXrbASF0g9h9Gd+SejeH1DqMfrI0tyVrIGSMICS4vpQYhc3hwyep1Ye
ti9us5LJ33ySPpmCBhkqri5rrMO7wkJhiJqgeqf/dM3oWO8tKW+5kV6CByNO5bHg
Wu+VP5KG4VQYDfp48DQQF+U4Eq1+EziEw1fawU9EiPY/YU2QacxCovwYWyh8zrZc
ZY+0tmSCIYqWxEZz86oqAD5hbZod7OxvQYGv3l5B0SD2o4NhyofU+DIDCfl6k4ge
xGj/HG/iMl+8pUPgxy+zT9gga7wyaMbr8NdYHUdFWD2eL0rn3Q6JZhQFUFehoxb3
m6X+uJpY3cLAB0TEpoqD+jMBEMGuPpwDqyx7UFdCzoRI7dBGaEFGQFLWjq9KMsY4
dOfUv1dwzVS0lUm3ZVjsZND4cSfS3Ms/L0B/L54Q6YUE0tvhB/qxrOd0d6fLG1Ny
CJxgNdcj5ya0NjHVUb4fQfPQYA59fUXIziuj66CGSUbGJdXCm9uQ+vCW53rywZEw
zhfBQ3HqbJMvw9cF9YskEMXG1K4iO6gyMR5kcuI/m2D6TM3ZXLrutQ0xqtLpDDQb
+BU6cP5kru39ZIZJWyciRll07T0+GGHhNpB7IZMfLty1kz7D9XbuEmziKaNGjzCG
slD/U6c1uzRfI9AAyC0Is+6UIrDs/sYdWJfysOvRV73mpIWIGEzL2VRJEaNJZiD9
yGLay/rTlC6vG1nUiCDaMxPHLzClTS362WDu/rGHJjxlpSWQSCbxKwY+d+oqYPhA
fdjI1QJK6GPIW5dEWavpDq5N+73L84jyZ2fwjHqyldjisXkbBH7bGSk6hobernSk
BJmVVk1aRwd/fKIYKIgJtjCw0xBMIJXwWyWf5QoSGjZJiBBqPFjjHbNwizMFrv+u
yS19QYHxAZEtHPQtMM1D67bodi58nCHJerDyOqfA4FPu9dPX5tdZw3FmxxZkMVrt
FqofehFV2GRVnTss9hhyjI80o9u2/xBNQR31Oelq63ftfeISysJs9STXeZ3GE+wS
zcOQTdwSuM6/u4nRQmjJnsc2OOLHpcm+w0nV87CZneSQoiqTplqnHX/Y0tLaBJsH
mID85m0XQK1DI3uJRsKpGm5XxnB+ZHXLzFqPycZyn1r+QsCs2XBIMbQoqsGqeiu0
swt39iRzVQnK/YqnwVyK8FhLxTHOYO/FmhjIcVdPI2bN7NMbuhiSUQqcsOqAy8rG
J1IbdU7cLhXYdj3wZd1gzOV+blijs9BGebquCFHTKPJDUEteS0RJycn/k8dWSMHd
6RkfwEPrA3w+6blak0bpeSiaZ1pSRi0NX5B7UvLXW+egYOCi8tP15LDzOEFktUUJ
1X+ThT8Ix9tMQiaKWhcfA+X8n/Vlo/zAPD7rwb+r55TdP1MN+3RJIL9vx1mkc6Eq
7lnDSzcT4FFu1UrHF7WKfCl7NpDmvkG8AQ6q1q/D4QYNqVE+FL7LlS/YlxfSm1Yi
Suea2jAkMwg1mMWBbU5ycYa0AeELBStYFkpOnxqWGb5n2MLGgIP3jA6oGvBLXK9g
97rQ0lIwp59AABhmi/X4DFPkz8koOvpjDZ4Bd6cfUrgha4YU+fv8U0vP9PfCAueY
5Yy/sRxe8Vb0feVutl0DMlztaSWHcMVH8iyuvqPAtIsaOEREk4eid57EUOqjeGJr
lAjoGvnb+LdEyOFflgpbQWBG+2i51r/hzWe54wS117ma9I3eIc723/Mad1RDsv1l
4Z2LTh+YZT3/zIcN7AiSp2PTgwtreGqSz/gV1aa6BmJFx5X+PlXNf58zwcK0lbYz
om5jD9nkOdPZXw+S3cfcNidsucV7f6NhGtinNe5K3Yv/CGcFMEsDFNEiS/9xwRdw
q+j4voCOF2tVIdPafmvw0mhSH7jhoT0jOnoGssJlCTT5qqMH7Thr0IuzlnkEVb8w
9m5/Ln8a33rd3gebzmngU9AR5opNfmfUe7nchInumehlCTvdPzaeyGu0yx2PbneX
zn/BqpQoBDd8wQzdhJ8hDecOMIpnZq6ellixsVAY77XZbUutlhCu3kxkbEvWFASL
fZ5SkTe56qGg8BWPZe8mum736UGRemEVjsNOaky8ydmIvMRonJ9HqA35UuyESUzv
P0E/KNGJrNyVYU7IfRvIb7FPuSz5vfIcmTuspsc6xAGaxBiCd9hb3zfXQUHstpgN
I2tvU7AX9g9LpUWRhnkcWIpxF1rkR8u+hAH2q1NqvP3a2HhIYCYlod1Cvb4WCwje
usK6r8j5bnlPGKW+TqloRZi7S5BAMvXeFpdd0z6Q4S/SsluwguYMxgEW7TTf1y9v
BIAXlfr7JK6pRqazCnou1tbGfJCo1jH5kUb1wBHP6E/whHL8w+sDnx8pr746weoc
AJZSVM2Lwx/PJQ5eP/PXoyWkkamFZh1fWzF3lspx70BrQv1xzLs3cbqyNI9YYV7Z
HZv52XGXDdM5Dx3KnmWN5+1naLDHPagedOCFA4DkCoOdOrBlz7G/kpNXNJz6MpnS
adqD/8418Npbkuz9z+88M9eWBmz6z+RJpPR1IzZ64vwkXK4mT7puovkmg9X/aprq
M60hiDAd6olCn8ZywGUxwLYTQ4cUveFBpZq8ml0HL3Aslr5PQFqpbSFDNYIYpkIs
Dt9DRiQjbS+Uhg+eSQyFqDUgk92l+t474law0kHyBIvG6047R4/p0pOlGtGV/N5k
MGYKoqYezbcHvDZFC+V04zTENN5xH4X8AhPn8VRX6YnSqueMntK431HVrSjXgTVq
UZIVQ0nq+yULyHy0X37SZfIA2tcRXz4mx9R9Y2sFj69PX9wzG4eYf27jlr/NfQCs
EEsWxArTVzD8XEIBcm++qFv7QBsCT7PqTpTqWjCRI7Zt0eGxuVpgO2fi0/FNXZxG
oIlvVWuMqKT1mVjivW0O+b3hKX3gU1mheeli5QXrPiGujWIDWo4b+JEjmVuDhXGz
uHDfjm3o+h8wa5RdGuptbPjGQIawnCCxh9hT/7GBX8QOEPwXVBPBg7wU7ysNVAXo
1m5c3l0bESAvAkQgivxkAfWXBwDdLyPKuKo+HljYnF6kWEOONxB/vQgopOLNtKbJ
Hf8P462CE4htlba7sZDm/05HUOD19vDbSg6LJQafFu54G8hTJ+4Xkw2M5vrpR19I
L41Q/a8X6RM320VfH1E1XxXuvc0aujq2m9jsJB2ZEVm1XH2tN9H6LY2bjj/lQmuf
rhLXGxnWRUeZtOGpmaJvCsPmjJKlD7bVa3W6bpvul65ICimXhXKFBWzcYx3R09Mu
0FOhMIcTFRiWK2RZLFGMy7CkzuA4iG7gKEsCTIf5wujpBovRuvpS45lIlP5gV20j
S9PutOfBcFyjqaMIn5k8E9iQv6mdnmgfCNqEodbT0seR/bGpymE5KprsGzBtYfkK
nu62PqmhZXDQ++ezJjvs5tjf8d2lCB0KvtA+0MCtz+KsdT6Gy/vjadWx8Chkr2vZ
CDkUpMGvi4RM5gQA+avv91zPr71SxbWQ0pC5wCe3wnDwDWPpoBCEbm/fxOQUvbq8
dJE+COPAfr3j+IJegDdhxzZhHvP9Q4Zn1NxRczbJRm75GNSXERM5kj+T2GKUxHKH
CIX9V937M8jJ7QXyd7/y4inqU/nlrMyFMVeMBui7DWL1PP8b3abocvSybSp0aJZA
pW0gjhP5a3h58UypBWTQHehiuXDHbJv3LXdXIwTTLJV3o5YKTm8asfdyHLBwHygm
H0ljNCuyosEL7J1fURI5Ipyfe8LRD7LG95jkVo9bpG8QA8XHgqIC4X4tt2OQLvvJ
BglsxIeLRdWP5zo1g4VDqOOsqnfPBYbUhiTt76Eoc9RzRXNajevJOTM/9Ms4bSvb
ehhGBOje+R5SqrIKJD6yY1rz6PQnsJUv8mFPYkvYJ7jClIgBwdSajIsXSbFTVqWk
pDvYNJHXMuhPqkJE8lo8FMb6ZEiGWL/U1qOWI6uWOWp8uilGfDtlvyniYEf5rwr2
a8lTmkbIHe1k1M+6tqQyzs12mk6SGX+uqaqTEqwPF+VcuqZ10ni5oeL1YORI+h4O
gvx3wgxGtIkCKngZvSkBGAkrP/Io2KJF7quuVl5amQfUWA8HHf3TG74y6FPMkSkx
Qon7fT3aQWtln71hraXwALMUZQ/yoGRMPe5xYQs0D9cGR1qkA4nbDDSRSfK71pVt
n91Nt2SPXvZeGUXlbONiOQuPaGsC8hjrqKGvqmz1gsFFBhQLLhZZgWYGRoGu3usT
lbuzAXk8DsGswvdJP8AWpClQN4WyMsMs2tcAZs8JuoRKwO22BQRprrSOF/zuHJ8V
BEIYJ5w1SC3w/eKvjVpCcIlgXSZ3Y/+gK1qDJfpcjdCJnPEbx8g7K5OfO45EsVMk
kZQb6aNM+09g+EjSr8nqIiOcE6Dc2rrvirFJrmq1+mt47bBtww8BeworciJXZBht
HNzlOZdzHcghyBNrBrlcI64GN0Dubf/Z0X3kbZiauCeATbxbaLfWjrwRSdeXhcU2
4t/EgTuxRRzKOgyWj9Leb0Xi55sbpPgAbd8DReLg5NJ7S2uSma/I7MqiWSeIN1Bh
5+LL2/Gp30W5aprPV+RUM92xRgbb2+LwFGE+krDWJliaCVuXy1pwg76IqNj2FEGu
rbiuLuVtlsk1Ov8Ip39GYbJqAFfq4Vz2eaYooreYGz5qXADEdFebjh81cOCIDlA7
2QKXOenasnyLV8cfi8wQK3yV96aQLpZK8GVXxWiD6ghhGrOvnMzgOgae87eZP7zK
bI0Bvk6H+dVxAtZrUZVj9dp2PkvaJY3UBnsnfabKJ+UswQKZpd/jK4z/7w+XV2Yp
jXA1x2NcArW+omaF4hBeSsVTakSa1ZOcXY5YNJA+yTCte2dHJqVN3lSScYHpqWWG
hwLRIua0deQFvtFFXXSVNBAqXScdD/5vdmn/S2O7qHp9jwSal8Lzia1KNlIhYyDl
NWIHardq8dop5e+yVCKeyclWu0M4l0HaGEQbWSC5qFCqUAzLHlRCOcHQHme9mjN1
YqLQGeIXL0r+kCjrqQLr9Bmee2qSq9zvzCEBJT92XTbJ5xdnWbCLim/MRtUnZpV1
Z3Rvbi4IAySvc62rdBKzxhiJY4MgCKx5BbDXi6MnycN9QZyw1qsd5a+CShIveCwP
3GR5BROVwV6VUl8BZcK6+nWHKXdkBw9H3FHRUeX1k91xqzhkWoV3pnLizbkXdTT2
6mnCdpOUNO/2SynFxXQvSTmCw1yBVIj4TiGdnoWsogPr/FtUo8Q5bCq6eHTlr1S3
u0xTKyYJDzhO2zvCyavLXO3S0jSnj7KiRDMhPNMUxjNyIAHMq10nmzeL/ahV6dUV
HOK26cQ0QeOQHQxocFha8L2+dI8V+9eyP2trlDNQOdBcck1MkDC232PNDfTub5un
oLVAvmAutBPjkDbs8iupSlG3yUrfFrzSZXcw0RFDhywKsmJ2FHn7IiArrmuZgcB5
5taPdmmyJdiQdjdC8nIhWg0kn0hzDEkzHOaMClaao5EQy8FvBdCTaLDd4ifaS4kt
HJjW7cAPyn7KN9fHa022ltX5WDOEWh2ko7eVfLxRFq6Dg7cSBby3nmT75OQwU2Rr
okpi3wfNlhjIV/xbV6+iYMA2flqx0IoLkJ2ZTdIcP7iFzadxjAVFy+wu4Zunhf47
YoK+NeJY+XTxPDYmyBYA5llUJhQKLcI/L9TRlXo4bfKWUcDwGoHoe5Qc2fKL9S/g
2V86trVNs7iR0jYonEtUbImWhVirTMkucgs1vt5bEhKrESfDzp2JvaW0HC9NJIVL
/5KCt5nplRo3LJqj4A/AcnFuSBMuPbZ8++nhQ4rlQYALilU8XhgQd9UoLq0t+ukd
D6MCXg9IodB9cgkpoya9X87b7/apnPxkUUMHblG8fjz3hVR0uF2lXQ3DH4lSxcDZ
eD+aljUtkJVwg373u0AwILiIOf+snVMyqKxBneLkC3rLaAiu/iAAHIbPoX3rYNSu
LObJz1PtFaR7wBcIwwgqWSqfKTmiWaLDzalXZj5kZucCYD3W2Lrd5nvR+0jikaKI
4q4jdONsRsWf/rfmBQsT0Yc3XrYAMW+1YYfqGKWD32a96a8ncjQgWXCS/wb4PcBj
zrpjctO23CbKleCd/rbaVWr0oxSwFqhMWp2MIVRTIzyAvGc8mQDRVX3RiNPQjK6/
V2lQOpmmDiP99FmSYSN0m3WR9qfhMKeTHbhvcEfJ8A3wAwuWsxjCzz3003R0l3FK
jkba18HfT9BNf52NyRBJqi+zo8TxMOoHNdKqWzlvgpLzal7kG5JMMqhHUVwQyPSF
yyEXWYPEmhaWRkWMy+UbpZcw3FpbSLNuQp8HJA5CojvK7bz1mYpHa/lqXPWm4Ny+
Cr+gxfK0OGpxgeemLJglDjPibMimD0CDh5H3CA8Vkn7Uze8tvFE5aFFbmGv6qh97
rL74UO2P788bRb2gR1T0jPil36bKw4/tGhFV54UbEBzzz02g9V159DTiLFs2pQJd
dgliZaxAaMCiZDCkfLgSW9CONJAEaVB/zSGbB4M8cSoPlPNt2lr6zeSZDa2Vpm0u
ETAGzD9/h1SOtX6te54upBLoHDD4Zly6IMOkKLe7UMPzmBc66zR+RIyTQ9Af68Wg
ilx7DIMiEP4DFWwTky/mDDxClX4EbNWIETTwbkjgkTzjEWrccwn8u7tz2ikob+Vm
78NzGfxxPeB5T8V7xzIQeG36vCSulxomY1YumtVuVH/K1ng0aOJKBSheluB4OxNR
6tkc7GFBl8tq1w9GrtNi31puUItcGU0yFbctTvoHQ/qcfWZU0nCxqYrShcY+preG
kHEAMNbyprJMQ+nty+r7rKh9bAliMH7Qu+0na8wKrKe1P4ydLyvHaxpcnK43bS1E
S39Z9OfNJPdaseu9rUYq1urd6rongL3F7LDga+43Gka69LiRPs99hFUj2VdreAHF
PLP62gZNt93lxxsZTEuGHpa17W5EXf2ULSZwSg9k7vr0A8siJX6EKTcUR+XHBMks
DyQbWG/xf5aSODNpWFYVx1EaWbuSUENVpm2PeK/ZBVjSMh50f/9D4XP6U+EMCh1H
cO+YZ/Dh4DOAYmc/ybRgamGvi5vq/Hd7l5PUtAHvJnbWrOErMeJF1P+yomgIS2jy
U1FDSF9mX2t7pj6Y0fa/oNA1Jyz9co/ipuIZ62k2mvNGCUzboL+E2ui4MixwL63k
eWntQq8LFdHzMJanMrkzOwflyGLKyReZMoC1uTKU85XGWuRGmgD2ogui8MXQUv/f
EU+GAwhz4AKYNlUz3sg5+/39bXNpDF0tHasnU1OfSewAJPvHsdwkpTKAQCQiqKaZ
o0q1sI27fh3ui4gK3lpkF+Bta5VpSuUIQEriqE46wYSHixdERDXdx5kUEU2LaqKS
O19nc3T4KTCUVErum2otrLFLBi4DclQMnzRahKilDcS6rXZ0nA/f5kuMkd3EyeD+
RDiVA06k0jD16ACGceHqsgGrEHZAcyZ/SFdgrALMyDQs817ZJXUJVKskIkty/Yfb
PQA7OFx9hc00SoM2fwPUS+3STJevWzt2V3e1xCYNJGAT6OyPcS1mK5a7QEBE5VqN
5CFrknt49Vtf98bz318gvRFlNFX+4X1QZi1p5NJpo/nC8CaoGhELVCNmQkBEWaEh
/aZsdSs/pcImlrsZBAV7vyxVXsArSszO0oGW7DDkSiZiTzfqD6BJ0Rs1jmCYRwd0
VmkWWVeXcequn30/LsSB5Wyqv9okscMbm6lfNVPNHbQH09Msqe1YsHfJOr/ipnZo
t3PBzXiykQlzeMgeVoWhKQ7/jLV7XfUn2oRsGVtoYfESJqz3PZ31qzmByHJ+9mtn
aFwGqMHGPVxHDMscYSUWdrLyHbDxkM/T2dpjPGuFT952C0C7LXOk+chFkyVdUJ8g
sZDX8JE+ApJkQpYe66+OuImc2UrOAL58Aq2MKdUVopQslM5wirCLYiW0HrKUIevd
oEjg7rbSzcJkj93nfPgUonUa3uZbyiGF6mhuY/KMqPb6uhO5OS8YUmIxOhtlL0HB
MRl3+QkZoOM3Kb80ul60Q+iVjEONlJR+hEEbEsFvVtHYdARm8ooaNHH1vh8HOeyb
d4pVYP3Xr7PciOMDRvx3FhVXoUqjazi6ocN4N3EVXYKxosOesiCNO4EdpdZUcN9d
4hKpTKCcxdhECgP++rZ3N1JCyHQyIXBurNKTQoY8FI8pTyffZZYHLytsP2esGx7L
ag2ImRTLlwmvZmktRgWM+/fWqJHDYsvrtoGlqsIi0NLgVwafHkP3sWqJFGwoaydJ
Mo7cUFVve+CJCj3BMvPLUseX5/2BLQor/oe5u+cu81gv5YWQB2nXqvfgA7IcZfZ7
F0mglhf5SLNeUs6GDDZzsxtx5qslzydajbXsUX4vPGV77YKEeO3UgSMljb4sS6sI
cbIGDFxi6Ew6zhGH/fVsXKs1DvBboBz22IEcJDqcYDO9HUL+1kspGhiE+8pI0J4d
TSQfxvYTchoTkOIIgyzXoK9b+BIUG5T7+8bbwoiA6Os7WBoHoug6RSjerzWvPF8u
WpvSwOv0kEqnvNNF8YvYpBBxuJKSp32tR9HzphhI+4XLgVm00lJFqCzvw2xGGRY8
2C6mEfblstQWP/07UoPd8jPYN+1cF4QBapUjlCzPA57hwjlDASnaWMAxkaWahN3M
usBXImfY49F+o7fjvrckH0wNBxayc7Kfj5qj/3mZncNBTWBGBR1zD1izkoOgPNBR
ex8d0LP+2sJy4p1IBT4HTSiuU4dJhPbcBvfcjSUFxOpqnt84PxWGCHNAgZxhF5sI
0zv5g0IUyBRyChRjLySImttL4L8Pjb3h9lv1XjXEZ4EPfJUi/Ror/PBlJWmEwchw
LBSS+uKa+X1ksQX43O538XvJ9Jdg1UErghAVoYPKhgRggs1uAxjM1WIVQrOaysLf
tkBtQPnVl4WTaVHS8CluQ81m7Z3W4K8/YpsQh3ubEMkfzQznT+ZQMyjD5mVgNwf+
me6B0r0qjozTuPo99PAzLIH2MK30j4jRePCgcnBEeC/bjahs+fJmEX961CNbMP0L
eO0oJRxT7MuCa3gZXUGSAwJHoppN08qetjzeNxtXL5XbvftWtjI11JxHHCeDTIAC
pbXD5T49NyneTFz2Dg7FcGWVVeOnMwDAIupBEi2y4Q+0O9YFg69/7zRSYMgl1ns2
y2DapTiyuFwVE0c1vD3qLeDfDbcPBU4mtEQDz8W1Cknb4u8HrWvENnmEKocPw6Ih
soXuNRPK2njJ3zItXySmwVnEK/LUf/OGufjwMDMmI/A+45sRfNdpik2P6Nf6SkbL
/7N/3Tf+fcX/iS2Z5SxDFMvG1zsgzpMdj9ADSoWVEd6kOpZ0PoQ07WEhGIBRtD5K
VaY4lz8nqNqLwYnqFBarqx6qGK1cuAabVam8zebWroJhbXPNnCj3dMvUcMz80Bhl
ymVFOJcS6priERe6WrWMpgKvMiPo27gOjVn3Tz7B+2J2/P04C6bU4p2bq9vU3xRH
k2r+6gqENJthsrlS5iFnraLuWSmGyWOJfmj6VKyoxMhGWsVZZkA+/7IPtAoyXAia
TdHpOmVWOmKx297AZzWS41u1SGZCrXHHN+ka8yIW08N22lHcOoaSX16QXbYX2FuX
+zLcTTLgG6WSHZolArFS2pIkWedMiike6X4s9GfSPPT9jLzRdJCvGEgru+xG0BcI
f/YJP8q+JkuwRlbA/m3wsvJiL8geYylsEEcDOqMCxoee1Zf8n/8XpSyt5lznNxpz
YJ2VehqGduBDxY2wIvyxl9PjsFfj/y5LsIdeNax5HcsFTQwect6VaYb1PXWaj9Rm
c23iw7lxubSZuKtTnC4rv53o3Yxe6E9mouTXJjJZcnjVCaelarbABSv6E4wBCDSc
NCvJeP50JfXgKNj8ZeBhjGiwNlTKR7ht/tae6q/tFaSUyJFs98y3qRDXD1TGCT2R
bERWUZssPSVBo1lWNCN5b74aM18ETrC+BcPU1ra4P+ukfagUJBt+1N68vrK4zvjq
26GGrCvVLIrGzXrOTh+VQzvCZbsM8WxR6wM8YCxuE5P7UDg+tSpuuQAHm0T04h/y
iu2XcKRpNmSP1HEXlJ51M5HTyLbMe3Jen7IyadCfjnKObccPEtMr6eHpqU41a3m6
Ls9k9R40aNROp38Z4RHq12LA/GTV4oIUbWDsC1N7jNkj29AFhVndvMIXAKLpCis5
IblEFUDH+M5Ik2ECTHAB7OneC6KyFLgGS2hj8pXGZbg2Pbkpa3P/tV7Dv53YLod0
LSi/BN0oOl/yzdsSh2PoMw6Dzk7vtT7V34PD2NGvfWf1NZjm6v5MC4Rq8GS/25rt
h3XQWyXTrXiJ0laMYzgOQPllFOc5hY/2Thun9DPWKTwXvl6frHD8/CoOjDBMAKOX
UoROj6fEbsWs0R0w0BxUTsUwqo3W8oZsFzBMS/WvZT0DWkt97F/LGlLOPFje1Nfr
uLqfOZKxg9iZF/8r1KIJAsL7x54YXS2rms7qpY565OHCmuMwU27//2+JhxyhSscx
tpj0ZB1Pu6blcRhSY1h+gU0SE+AVmB7ToLvOva4Z00ueP+pUSiR3RhzR4AoKCGKL
DqgNedP3uULoyGeBnKw1sDGw2kcH6mLAX0aKfDNTyuYgEUP3aM/QbBqAzNp3VK9K
4Qhewi9wC0hSuhslmyFj9vH4mVykSOfLd94US6NNjsVtGBv7AmiwC+fc+IV3Q34j
APgIFmXULq4GE+Fplk3+g6ZEIienSyExHN7zgksauDmqBITZRCgdEh+rNUR23KXX
IyPVtf+EBDfXpTAgX4hEQgnpbWe40Y5nDc77obovNMlbnRbgc0rtUq5galyF1Sb8
NH2KD66bz+dIseDlhizwOYhiSQkAl33oSHwBW5Hi2He1XbjciDPxHIUXvcQ/Gf53
pJ5oF4vmmpaVVuY2q5Dzyi1U5DZ7wnfqzR8tV3TNcmwf8UEhSaW09guMBSY6HGlv
KS5lFIv4jXojBoL+QBaRZUbV2wkKo/0yVV7jjAnv3Ts/BbxwRkAuR0DQWUXGdTc1
ORCXxSSennJG/4VOMohS1E12kKd7f7Am37GHaskMHiAWnJJrb1qZ4pkIaA5l6M0w
yvGZXD27hAB+WoIqTDUFMnzYUagkKqmU6Glc1HkNxg5/kCza2+Ca+Hag8/kQjNG5
unjtVnI5hMsuHRbKxXnKAWxGeBRC4S096PgC8DibNYWi2TaKo36/Tgp2BZdoUZuQ
6NmH3VmosOUrEWL1IHd1/FiDMtNantoghGmBktPEYrD+IFKubE8+FKZz1ZTuI5fb
yoLa6KW0t5pb+7BnL2VKtgoTqf+YZkAfUF/SSDJepF1ZXYiHP1tRgBwN7OY6HBvu
ALqA5Dmt/1paep+rFYL9d/67sOaynPD52LSIPJbNzvkOwylwVb2V0Rtkyyp0M8jZ
qtJnKbTRS03+zoD9nO7Y+TUUJZjhIUs7DoyLZ3xPjnJKdv4ppSvtdl6SVDl5QFbC
kBfcDB3MfBZgHLPtKAev/affTFQnAgxNXMYrnq1WuX9p/h1tAOMg3Xjd8MMfV9ee
A9He+SxQHCSpLzx7jDl+3yl/UZmzF1RMSLD+5Ldfj4z3o2SpbtIhN9vL51mm2FFa
hqSJ47IOByyB2339rCXNSIv6DT/p4i3EPkuzgtbgR6leUi9zVHJ8RUezZUqOERhS
Y95Qqk14zA9URKHP+fJ+GTKKxZhOVEU2SpC/LvSn52Kd/Ybl/jA+zs9ifSLhqJF4
tbhcYDePmrxdtt+IUS0gWuAY4hrD4T00joYU5YyGPxgATIS77eIowzq+xXmET1w4
zwSPM0eZSsMNI5nRVJn6hxH3KsxpHkHYsKikBK+sO8nBosMHeO9B5URkSK/z6Gfk
hIjGq7UdH2WUxiGvNeU4HUEWXfmzfw1/6am6ek/nkEDdDipf8R1u73rY3WjBO8Qp
L4tkHTFEZOytIjnRpV/7/MigLftUYvjJM/zgOsyGiWZ5qP5Pz7kaeLmUA8Ut0+kb
7LbWiP5VmFt7spUQpn7QWuu6qgzO/6mcYxVbW+SplS9vjlzvPgglUiDwyDqJSTwV
PRKJ4EXLamDEqbaNmENx+ilh1ucph7kmlhdwVQB8J6g7FTaCniXq2CIQsLlw3DJD
8Jbdrq0vJJTjKpbl+SWuJbRUcjB3yqTr7Oi7crm/MtekX6dcoFqXF/LcpeGto3/M
IaGtUol1xudnuT1Oxz26y+EpicJAGKlPAjcg5ZwuIo57TqhydC7ZYlFAIoWvj+9S
eYB03osEfy13Rz74bopue4dHYVMoEMar0NSO9SQtY755gH95N2aK+dxDNy4pPoGR
0M9ScuGZGNuCRNCHYqF0xAQYwPtsMnML0mQFi2/OoA6Yb+nsI9HfsuOhohczKClz
jkR3c4NSbC3bFCyHGL4cKvsbsAiUlTJyPNdJVEwLLGnW+Z6oFbwcKIoszXTQuma6
f0iEeQ/3xLKk9LkFU9JmLTjqn8MNMSweVp2Vxq7anf+qa24xq7YKQpqyhslmH5rm
KrXQ5qcMDTBcWvb04DtP4FNpRNNyY/aAoKM4TWLeRtXvyJZHe+spL3grwiEEQmBg
KgBaWe/5Cic3AXFeSsz94tQq8CzsJdD6MxcIkX0f0sQF7Hcw38dc8yf4pf9bWec0
OTC4Vaj3Y7B1DcorsstMVmgth9A094uYtWvQY0AjLHkQ4U5OFLLjp/ilTItrwWd4
9/P3DOginoNzgRD1gtz7VJ+R//eRrQAliMr+rMUUmNHfgmFdAcU9DIVVCOIoBpQO
jXSZcKybxzJXdnvCZfGUY3MGMZwrReyX+7nzoP+cJruKExKxDFrswwj3pB+in7rX
X3zmTidPStMrcrzIt+W9WNkipN6TLaqjJgo6VMNHVyYYFZu/G3BddLUPRnLyDFEp
f+4WC8ZW/fjcRmLrwyb2ygnChb1CE+zxKfL6FhgxX6KQ6sZJXiHh3UMtRa4FQo56
rZegEGPjZrEtuWGuGy2R5C02/x95rwWbjbakhdOo1D1xrgf8PYn44s5m4U+hedkr
y04b1d5e3y6mdOpVGbYVCEkzovkNrZ0XB3CrGpaL2RByGbTAprQ1CkGanCqeepM+
FnoEfuyKqFgQ7W0fYfHhd1YJ40V0zh+ql0OYyYZVZy6uPvOv43O4HHnBgCuhYaws
4iSdBx+1CFeBevVzTeVxSuzLAzXBUyX26wh3pQ6fb3r/0q4ID9lE1bEAVsTcnfsA
t6rjf4QPKryEMoCgMXRWN0UzcKHJDxDo7EHtofHkyHPg9j8kPONxNIhA1uLiJeAB
fi27t30DKPGU6QqZWZyeq59FtFzvgBo2kT5Ow6GvOlahf5yBNvZ8epM7x9QTRTzN
Hy8PYr6+Q8fwNL83bQHrBf8K/aFv9pLVk/xBNeBUttW/p8Z+txudmH+bx0U5aXPV
wKElhUGkMWmK0eQ95anJNWdFjvBrHv7dSH1T6aWGA9YUG/uIRE8TpljpKspqdjhF
bZazAdvZyWbPqyU9l630KlrGjRLe7/f9UKA2DXp1cJIxH07qDKl0G3/UxS1YZvQK
QWUohHviXN77f1EnjNrnbHxUKmWB3ZpF47uXHn+EpBF19y47+NAvAgCPMI8VkxSr
HBQ7N65fdzZr5HaWcsuyOboojTZG9rKGrp16ikBMu1C0O96Jy7PGMqSuuZ4LGZXN
33rgFvQ3Ke4n2DraMl6XogWha8JzjzvPZqrqNqoYc0lWq/JpxpUeoHiS+aP/AJ2g
IeN+frjEnS742cHJGPNgl6KcZI7CilRJcbPzhtf87ndcWXpbS/2Ug2v6p0z/ktpG
YV+F4MaLFDwISnnpLi0lMvyrvXCMe0iuuCg5mSVLC5ruM7qQzNYqv9hk+d/d+MdH
ja5IGNCyB1NaR4xG8FWtxd5cVS2L3yvx79Ov7DBRIqWa02kEyHfd2ejGDP8ke2NZ
dQaf/9azmsUx3h4fAVvAMRmBJcmki00cOThHX737W2jK0uRcrX3V58jyzpu8JzMN
cZ0cWiD1JfoHlLGwElHuxL/+a8Mtpzfzi+gfHxge4mdnFnfz1/krNVS31z3Q7LfS
9/vtH1L1oaSQvIe5vUntZB+7neD0Len4KWp3bybXiPl/6LZWLA4DIeXo9Cu/Qtti
2yTOHtwqx/h586DU3iFDdnDl+GsAUoFhwPHmTqHfO+Y22dOrdYRXJ+xh8VryyNej
HsUuAalRHJzz92R7St+11MpP3GYxzdfynWhWspO+yVzGgHQBxVSNTtypzPgX2UWW
Jcz7msxkdZe1FrBpk/gKNeGPqoaRn6sIM2YvA9eLQv1iflCqQKZBroyJAuB9wsBd
yzgQw4zOwBgbkkMzUfSl7O5csvHWjm0HOhqQbqg8ADDfvR+ngSKJxJcY1jvpNyLr
0pXGcJLabUm7i90A2Zh/wcEry0CpGZ6IhDg7mo+bercWSrpU3IbU8wAuaS/cXQYN
HaZ/U3KsE2HZneP1t91JgmvuxBLVsyFUKxijARVsi9ZREVxia1sylOwaBJtcehVu
LklmUsHVVdWLXErVqVW/VEoqywedmQLe89SjKJ0XKwG3FgT807qfzX9Mkjz7JWbz
gjIqQzJ2cXf/mly5LuCXTHPIFu9Jsl7hyCgjtq8CPV0CSX4YBSsNapx0hNsnULPq
27ezjvArRqGmkAkVEjnbS384Y/RnUcs7q5QQEbeJsYuDfPu2V4gFGW7gsFBqr2Gb
aRkYY5VwVqNkm/pWuAcPh9Nno4YhCz6Ws5iBXNYXUPZPCQ2nacfNsBempYi8hkFA
HP67e6lLxOLIwJsh+Wg7SQiseS+Vi9J+yOGYBybDBhdYLTJSioqVLUPjod+d4tLo
uVsa1UpV9wXhLTQJXclp1B9XU6PXdfefUJltTryYza6ztXr2o3aDqvvWymf/9YhE
UOGTttSAlglNB/IedAnzmiLRs63FoQF8kVMdEq1L8eGsRKHRGvSLCjQEBU88hk4s
PHXq4dFp6Od69D3yFU/bpY4EUFb+g0oB3zQ+qQ2AqEzJq+vkk1xbE+DPKSFlT5t1
BbrSgzMMM9K9PpnAMiS4eYxyUBXVJLNMSw0cfak2IZ7bTJiBxSqDTWV4nNRQS2V9
yt+J3qy75WRuAak4+2Sk0L34q6YKjvPl9BJjwy0Vn3q41oche8fyVUKbdz3pHmJw
nfC22ViUfzpi4h0NpIKe7dUG9YI9TI5CWEEOs4U9yvy/mhq1b+lyI2Z+Fvza27uo
Rxf0TzPp9IwC+vlv1iG5SwJ+3yz8J6XDLvgWbp7m1QTB8r086omwoVNvfZPmUmBX
V2yWMrI+SkO28voXaYnPtGD2EBVnv4cZNo35YsJrY6ObFeVY3QrpgZ++vVnD5tIj
7ShM4PtaD6ANxRPwL5oWm+HajdOk7PEYkI1UN+cbkuTWzzuFx0B9M6qerEXIxZ5a
y+TB2dG3iW9Vn0o5IOVu+3mnfxixmDAMKZG3lJh/lqJoh6/K+yivhYnsuqW16h0O
YYlm79nTtOsFZkRUjB1gv/BBx3Y4gDOTw7GuR7XxZTt62VtCu/sUWlK2Tc30jwSK
lC+/xfglWjeMZ6vIGJV1vhxpfpOzR4HLkY2KqRwGGM5PsqfEAZSTRQ2l8oBTROaP
p2vCdaV8qEyllmZwPyfmcbrXFojWW57LaFFrHQ/WoRVFUxC+ot5GpeLb/oj+mU0v
DwR9aOvkz8CWMkU9OC2bVTdbLF6+wpHruz9Vb7N3Ln3kabdDTNYKSCM7J8l6+QZ7
yVNYoqcG2y+JXobZQCEh8hAM3fQmAmDEFa/986+kRonF6LL/z8fFzGM5WlT8wak/
vXNdXLK9GHg3OIjFmziT8YUpuqEogy+SpNN972RORQ8JDQPHNpMHjlRm2jJ6gf0A
EXN+DtOsAWSEIVMUqrvjI2p4xrBj9ZWfwbJRlR0P2eM0V62URyv4/EiL80NSfZ/9
jlJBExhdI9Cyw9KHcj9g8HXdJ078h0BfvLli3CC04QvZzKhSIMMkx6o/JdXLuUwf
SML6g5RfmbKC0FlFTUkTCuJyChwaw8canfRZNGu1+jNoavczIZXVJC3hWQvRibFC
0UYDRpMPK3BBpACAVSpAS6mrWQPQpJTWAb/LuGGGNEUsEXJAbGJD7493OXeXWCmq
gz5G3veGkW+JKDc53XTVgl0vFH2mzYZdsndA+Q2Hw08ZKhwAGEcJNXwj7kQHK0mf
MOlGzsw/USNk7NINtyzyMG8rryhZHFPwditXatG8BKHWkasl5vSSP1O/fuRthKhy
Pxr2waDWjB/gExrpg3RjrVx3H8uAsLVEe3weDe6fNgaQTDOqv/DuLK3kox+WqMli
mseAdgMrpEYNNQhHyRcn8v8C63ysQPOozds1j+tCJMt1KWE7r0991+QfrZQKG2Bp
8d3e3oQ0V9GR2cqFy0kyW9w9iksyTfqdsZiTYKVcC/h6PtluY0bKn4Gli01BOplV
n0QxjdnP680dYe26ISvapdqXuJUIvgEaSLh8chF9SP4dXySqf4NYgvlw8ncUJRU9
ZN06NBQT+vV3gPTpZXTYKd9tyP/V24IB6zKwWSnfDABVbeWBtVqfmiwqcAMgXoNh
8vv7gEUg0rewtTFU7ROCru7k+8Q+f+I97oQ5FU5Ih8tLDqr5tlOvxVm4ywp27D5Y
YHxt5mMs7P9QKOH/rT8Chjvx9Y0abFJ2ja2902nlUcaUIJXl9Qc0qRuSoVwhK0aC
plW9pZwhVaah/qQrz3HnaKvof00N39l8kQwshMSrNQlgvL+AcsZKPxnsUtfoSpWQ
j8wfX1bD8TgALiv/YEy+CkhgaIv8/fLlG88L7MfFGC9xDmzF7bBiG1pqjK5LOu6J
l1/7x2bcWEDgoydGJ4VwNmiZeCjCI8rkdXI8ev0B/l9tPWxC2iH/DARXsQZyQ2nX
LGv9b3QtuLKG1rJesf5SXjmjUva9Ooctgj7uqgTWFAzzNgmOkQA6nYVt/7zkX7za
NWFRZw2Dw278C8tnzT+0R5m7BLUBZoOT0dx6avmamyvXHk83Oep5gEIRX1mMfiv3
Xc9agc5oE6rBDEZosqa2ORF18IJ4N6E3MpxpHQn8xFmVFzFX94qt3kn1JA0xCH1T
68M2Oue+NvyB/8UaQtDt3aHhaAYtFGX5Xc42RljXkHx5EjzKBGMkGhH52Qzir/bB
cQfJEpX7ytu56nuN1u6LTn0x/ypT7GTP6/c8L2un6wz5WFZMV0fgnFJN2x0l7pBS
T2ZAMucZE5EOTiuT+6XgNOC885WQqkFQVFY1aVjgqIyMV6rFq5YPx2TKqR3lw8yV
iezORykX/IJg/Ux2gsP6mWHIwrsjRcI9A8hOzFBxmJM+r6LzBCon58iG1s6dwMEz
LVCz10lGBsrFdeqoDKPMhz1tSN6IdeUMTvGu9ErHWeGE2Dwm1ZIq2iG+/RPuaZRM
PeWLloA5gjrZEieyXr/oq0JRItn7kGLftdDIESzjZDvw230VgzOJ5O93TtTfpOPo
JI7D/j3T3MYE/cLNOB4WiJEZ1w140hsjshqgExS/mqyP+I6JQ1QkU0MLU6NpMkWj
3ZonXyUDISAjR9H8yieOmLMmkE+TkHPMCKOEORFrbVIg4Je+wVCHPgelAAmzUl6B
kB0lO5rroUNpRcAHASRU2pTIr71/73UpRLicRWc1/D0s79NhBERXseHYXyTsPE2G
JQ84M4qT3am3RrMFU4+BQuUzgTH4iYc4qdDJvF2AKNrxoPkCAnVnoAxnXX+ejVo6
Ycwkc3frYoNtUDUsQq95hNJGvfFmWnK+XmRYtOUMrZuu6P1QVAH6pkNGicbxy8PK
pDJL257tuG0y2zdRUo+o0iy0qJdF3qNEYhd1RPsXcAxeFv5W+rZgpvo5+PVq/nIm
6Ouk7a8sJl99IEngrBUCDiXfRO6qmO1Agc1EtwyU4jVOSP0LxwJkLLP51DjNwoC0
75d1bq56mefjmPB5fWFh22VCfvX78Pxv/xVnskfpMKOcUKw7Ck92QDforbvtHfM2
tjUAWv2U6aa3pmIhq/w4tKCJh56itFIaQ2m5WGMOBIaSQcrmmUV/XcHKlkXXcyI8
olaWNWjvm2JSYdz98Hb44kK8FFOP3rXlrz65ejDbdrFi/MvAIFTa9DHA462qglNs
Y63RTKNn8gqFPgMe9zbeoA7nrVu50vX7AQfGGN6q2mTIAmX84QRmeP8ZCp2gQ4/x
aJlFA4P3BzLMoicoRdANyEvdhwHLxQYEK2hESqYFD9mdHHCw8Uio6PToCQwmv02R
nk1lMJKZhKGwYNE2Se0z3/QRtrvQNwH5LVGIcv5q7335WuIQu4QEya+ZgVAHXyGp
QRlMwO+H2Zr1qWtR7DS5ITNkE7BEMIvqYtkT5JbsjbpDz5UaXER7Pafo8oDfS91t
3BZiQ8y/sVnJsDsQeUT3GxbE7+JpOgoiDS+JyJ/gv0vZmtT4mzxRWjVmw0HRyO/V
k6MMVf6sHQ546qbo+apezfnNTOOUDRs0sPn7MvagbqhhiwaDHL74aoKF/xKbGx+W
4E8OlHZbRZ3J2RN5mCVuWmVuNSVv3o8NYNCb+6ZzkfRMnOqx6nr9VANgs30NRzoc
HwAcipOcGHAiU+anNnB2Zup18w+f3ujHsSXVF5RbdFHAFHQDo+QwnRkYO779lNGs
YDd4VA52BH4y72iMw262TZPlzW2BDyhi0IJ1RUIk6d4uZLV0Z7mb2XBdaA9z8W9y
XgPsBTo1BXm/yiAWTNzkRHkHC+rwqW5df4Nm7rHOesCQZv1+NydN9sKeNdBTWwV/
WQTrukOflZd0myvXs08R9wt7BfQn+w2oHz56/JAlLchl3bw5XzQ7oTCruCsqguh2
I9LPrxW0SV5sb+ldZENgIcTXNfOOHdOxgX0YfXsCpCvJYQIH60YBsP7L9PPKDha6
4h3S5Axf7Gy2b2eApras8Bu5TAKin1L2r+ffEJz2ESrUnvqfgV4e8SnU7qnOk/yd
Ej/RFf43qKDGav6T3SVqaQSgqKga4i18Rf9LSKI4n8dnBk2KwixH3p4IJiNuVVtI
2Z0kbW903xv+WNJDo/Fx8OOFETEi7cDnvWRspxjifyjuzt+q7Olyt7MqazD9NsRF
EiV5Uc48sfxMh6hqK+EjbLc4VgrSjTSeM2Wp1WbvtzQYdgfRoDGo3+2by3Y+GucO
1rcFak0RW+LrqVWyR4u3B1/WGY59Ml+n5XmVyKZDDzFMXIjvX5EuYYwQW6wnzgYF
lGlz01G4IRPZqi0i2fu7/mMUj4kmT+kGD6PkH+uE3G+s05bz/EVvUFPmI8xWc5co
4bcdh5y5Em8CFGyL7x3L6a0YFpy9HkvMlNFIfK7loINv+WuHi6EHVtw0y2FZfPyW
DLs42upg9yDc1nBHs53FcPkMro6xO32jFRDGXqZD5Vj5QKeYvQEftrYOYFXHQ+ki
YeSeUcWd1bcGv6bTdwTLxXMTErKhTx3QqCYNCtaAnGlwv2M9ReTypkhpmDt6KDfD
MfCQj05NYjjUnEt7hcGmeo6HbMTFSOMO4bhas4qPfTvXfygNhN2Cxw88/yeOZf7f
wBjCjgqVrZgYZcBDWkplTCctsEPsVoBKzvkn5zM/gdP4Zm3gxwUX2w4Os72Pltrx
KHfR/dKPGt+rTyRIKmjkjUns2RvjPHd4BhWLIaScWkGpsrZbkxOs8F1AdGyaF/ew
Bb6jn4ieUK3kSHAfTKa8pYvTJ5ctQWZ14WdtIt49OsvElqr5VpCrYc6DvIwRPU3l
0aO314uZVxfZFsjdbXaL0/bhd3BT72xqfrdFP0oHKWxXMiUbkTKhAjJVghciYble
/GNOQ8BpS8M9ALL6CqTSklm6OEmJEEcz2kX8erz3ReP6cobUiVcFQk1sQCk1X3Ye
T99x4Gn+SGnfiIWERsBIiiWAnvoJlzenV8nMR+T/wK8XsUT8ozMP345Tjg5oBh0D
mdai6rFzEXOyh4MSv8r4CnM1iJIA+R/ygKTD4BYHvJAYr0zunaH3TGrtsb4exvrz
/hXWBKODfIJI4hk5C+J3uwLv6IgG6wYVq95l34XBgrckM+K8epa+9VcH+g/dpXLw
qgE7tgQQuSAcAwGVb+9BPbQmfzhKlwfClGeaKqXValDdWgSF5OkEzVSxWayr6G8a
Bsbliym7F//LPjAQlc1vwIbYSCdRWkUMpZIhxjnSWUZkxWRzS51ob3TjSvUzPIvR
rPqufgQlRapBakBpxniju59ZHc+0Z8ybLIxjgNT7MNOlxazXRSH8TUmr/xc+uHhO
/XfVLkVqHJaN3fPWC4+RldnqCVmOfpe0vN+bC5xCVXMF9dfeJ92+QJunur3K2Tu8
gR2R7bU87dYeJtNGCKyZyzbI8kP6s57IKF6B/GvlPI1hc7f+NcaNnOKhl2E8uUVt
52rlkJrfLo3hiZSxHCe5Hdr0ZOAGNg4a5dzPZfx4ZjP0lHAy+bpI8/v590+p/2HK
TGDUDDuLSN3Xq0zFVFvbH7n8VZIVULbAyy4COoGesZqzojLpDW0MKLkB1aYpiWNn
XrLw1ldnqC29MIEv2JsYjr1l9b3/ptuZjyst2wphXB517nuPuMuCDv231cxh9RRs
fZ0MhKW3oKv1RdS0Aj8p64gXRbV0oFAWWb/smRmOlVxRv1VQKWq2huedbnD/uaX+
v7bqjm7GK8owRx6AmNJrqJuYQfBZnJNSaahYXUm8DBZLspfG9xw7y9Mrlxvp/qrq
qITI90LHqh7u/wiJh0iR9Zwz8ffH8bIZXoMmxfxqcOhaqCtjFSTaX4VuMZZ5aTSH
zNu6hsmoCYB7V9Gl73dSXsWHaIVZPs9Z7Fq9zVqwguQo1HCmU1Hm0YfGty2UHwg/
dTe0kxaBEd7/TojaPzpwjuq5LlsueUEWuDu+hny8m9Uvy1guV0x2Gxva2RfYvbw/
yFR9ePob7HCrTdmKftHdztDMGELZ58v6DfVPbh8eqnPKMuxfjLB0YeHXgpGrfOiz
7HLzl5K+097gotpS5pVU1Ibabo58msWgQwblsji857fk2n9bUKa/bTJrZ2iuyTSK
cwZ2i4NAncP9td2cyF3H7cIwSCVWe33k8yPVF41picxMobppVMYTdf9Y4HxKk1aR
fCQI40Z2823VfM6RXRH/79EQT0oC5qJORZ4KNC/qTs+nEsdG4BOufoJCv8ra6MSW
Q4PPF/HvuvgpPNARHzi1bTWQkU3uCyNrim/6oX9BQ0wQL8UPM2OJl+ocFvY1CePY
E+x6EdCVEK9PL03mqb2qcsuq77zGkud4VOZAGfgcQZOjvO62x7tiY1zh9s/6n6H8
wDckWBGhQ1DYYnA2Eg24GH49TiSGcTMgFiOm8C4fLxF3yH4sKMUO4goMCqv4JaJ/
GMxz0SlsFQblmD2kI1DrbCVFQOfXjSpw++1r0z3wEkUTK4iL/15aPawMCxCgVtEl
F1l5K0S1Ykkqevu4CC5kCwlQjssXFy8a0P/2TnDOxyPEXLzIJZA0AsWUxnHE0TGf
SAW43c2PHMJYgPeyv9HKs163jP0ni1314diLEwYf9230I5qC1w2PoaBhvqAuX+LH
SpG1YN+iRSauJGLhCq5pc2+YUaL33IHEbDq4MfKYsPfKoyC1vps0KP8VQsT39x1N
0QvP1xON+1HUUITr1lhFaWz+ULUZGhqU51ZtM9jPD88bbqFi3Gey9NF3nDLFHQkX
Bcz2F+Tau+3+aFwM/+S84JApDLgjovMXgfGDmWE3qlbbSVFxbQ1h1fcDuLYFwaiW
/uktPam3dGbfEZu2zBHlBAUgUUIgp5ocK9MbgcGPQ9MWJ1/b3oL1d4zxzt4wBcUm
q0jcSuwVv79F63VhrVFBJJDPjPYOnY2ah6igc/tnywgdJEUj+N3U+3RLtbmsx7jU
xECeb5LMvFGsd/9a7YuPbg++3Xqs8gHsw29CcZxgFJrKE8gVc7db7ryXSf+ev2PL
JK4mAg6POXywr39Bel7hhBi9PIMNG/mTGa+QZ1NIypieX7QNFrCydPd5T8FtDe9T
NgJVRvCt/qHj3ol+Nodgeri+9OPkU6h8GSPRdASKo/kBOvpCx8q4yEXx5kv6ZWcv
vJS12qreA4B7CRSec2sCJkQrXZSCbwmtE05HjtVJFSu9/LP0qXEq/eZ9rbpX1IAE
gXZc2DrmUfT85skNDPD8qTNAfaujLkBSGsF/aNcW6+gXY5n4GqqQ1kuADXLgYblG
TWj/Ui1qTjJdn9IsKRAgrqDheVM95m0OwmyYISoh92zJk988tVXLtNF98ur/yX6J
kPVKrOiXxYh1MG3DyXwhdIY7dBVy/sJrvjHXXgnk4gVJLII7xlgOBQxKS9RYCBPr
ek9D6S90QmhJDkwbSYUfuNIHqR1i7fenEJinOZFKNPP6bTijPywx/F2OMiy8rmuO
reIF8hXnYED84xCjfndAk4xTrtEpCw8NLehHhvX4D1GPmniapMmAJy7XjMqWdhmz
MXoWv+eGCWhgfXmeM/06k6n0yW2p4++mYQW8K75rh6qkttDog+md1sDNNyRqRfYL
lmu4PBtF48sl/wsAJgBeQ4EfCrrqPc2fWb8mpi4z8dt/8z2JhFiVIZiAZke4UcWR
XYHtWIIxMY561ZKy40VKv8V/Wrq2WBvnC5YQzjBn2pwE/YRGVCw7CyJ/GjstLeBF
O+U+LeLur9YUNt8noBpc79qxpn973ySunm/M1S42hhJZcO0zpd4GEnQal4Oz06ie
P7u/qOqVURoEIfGIWFGkIJg/WMMOz1Iq2WwjQzh0NYG8XuS2KBEX8THJUDMgXEgq
ihKRtmKwGxAcoKBr1p618+4Bp5aYZ49/OhEd/RlyGUi/Mkmw6xsw+GvsWsXey+NQ
/AxEaVgZ2k2Q5MQxMNfXeNQiMIh6kKglYR+LmBULVwQr/iSeBckQd0X8lMvim7a0
E1SS5ntRjrS6TZT7+Gnh9nT7hsdekPO1HKRmZa8krcAfuLe8r5wYN6IrFj5/QBtN
H0u0hKz1J3t7WXXp4WJ7drnshccS2brStJHQiMw4pw/NeAIwS+NLANGYAbFtgHkY
9rUBqjjG+pUMRteif+S/W000IuMMrOPnAzPsh8HOQpt2LSGBITbekw5wwy02IPOw
zDSdAjGcthN+PGgDbKdtegVm3kdDrJtJsYjAHoDjMeZk3gQ4xzdhu6KQG4V1n8Zi
M9sks9Q+9qq+pG3q6AWp+jjM0D6wRisymeXNTKJnr1A5gyyLerhilYM4Mzbi5m69
D4lOMt/a0x9dNhRhF0ohfSOpMf4S+Fb6/edsqGMAqI1vVswP9eMYXudxgiGTTgU+
2dfqYtgi7KZ0w+BkOpYsxNZtFwL0Gc3AtVc1pQETFR29B+sA45wyYVgLpOKosVUL
NyObSTUllZwZWtLXaVUdjl1AHUzw82CmJQY6+eVE0jOpzeP2OlUPvX28BmNSnuNd
G5rz3OnEDdcaxwCoNyfdHM727e3d0LkmNZf56/nhL9CcHiLvyTZqsojxt6SLThvd
E3yD22c7Hh82KNW7DSOkQ91QJE2gKdeJF1qQQUxAdnyXxwJxZzBxGrbefkSPYjsg
xYYNR/4MW5VC3Nb+p/qHClz9qFibx/fwAoc1mv+hqnzHv3Fdp/009zXAvuU+nE35
Z+dUKkJfUqGatpjp7A1rYitPGJGKq/7p/d1Qq1Q5IJ53FyI6tiKxhSCfTverxNWY
HYiOHg5HJkus82BgBmLZRePH+bGA5vXUvXswXN0TjBKw1H5C4ONGGO4loogl8B3g
8qcOuSSIRCcZP4S5qJ8vCLoP48k13RHcUV1mi1jclT9CryRFAmZfsOVaxkFJEjCa
FFdCpBX6h+6satPiSteC7D0saVKGgj2vyukll1JANYCtCnSC59xZq2Aj7GyWWfgV
xtYySP+r8Tx/yrUY7qkcfPJagH+X4ymBSdUITPmbp8X/TF16h5Lrl/P3PqSBJvlx
YUS+xqgd2SnT097rHbEhoD+BpmWRWelr9YBX0Y7lnIJdYnQi+ih9buDEXuEfdpjU
iBKMK2P2+/DJEnpQIXcAi+f6Bvh5JIXNXGUrDTMc3GKoz3OJHSmYAAlq4OqD25E7
ZXQEaUW7TskeJRwtZi49iKz2UoMoxZnPuyt3C8ysn8fHnem1bFj5jV8ceXH/kyrL
DhVkERuyizjrFGofUB5ePAscbG4sAURs6Zto9gQwxxNnVCdANSbw+CbZGENLl7+L
Sey6XxdRjSO/SnL54DZkjD3GyTwF72RAGYkiCjI066LlP9Ww3VFmOVpexs8CDp5c
xNshrLikYc1RBVlCdAP4mPQhly0lgS6lPawge2taGkfKkDUPX8u+0wLKcl2G6dOX
dQoa4P6jbTtUdeFgnGBEbvw0iWPlLEoLBuhkFUWAhl8+Y4ZJQmUctPYhEyKbhuj9
EE+FsnMkbs2fDawiCjoCM1IZH3oiQeSZ5xf/+RH//ed0b06BbMdFd2eqdxoRa3Ub
dt2wPPTGIcOA7K4wu8WTXRC6ktUIXe27xIfiTUzs7gA/sL+1CitvtBsapLeBSaww
ud7L8hjTlZmKa6k0fC5uaK7myeZQeh2NVUvtlIWyPQoqYI/KYkTu+9b5o93txShl
YuwHkm1Kaj89wpZCmzKyBpqFzfMO1XgZLsre5/AQxENb14wG/SETger1Xs2LZZ1s
dUGfzCFzHQVZ4zhPZKq8tsl4nD+jLEPsYWN8j7vI0rjfhXhX8TllagqMzvMzktW+
qTHO6SI9uNhyzR4ZIt/VQq39wc2SwxdTE4OfEHz7unw7fbj6tFzQzBYNdeuQ5wdL
Nv0PG6fRdV5mZvNR1q9v0XcKGsSVJqRdjS3GVcO/NTOJp3BnwzF92R+w6xcu8yon
0ZJqz22RLm3D4ON/OFGq/886Bb7vktxTzsDTC7zdJYDDsAOvgCIIfkrUCYVPsln3
BDFr3phABl3UfOkbKrTA5BiwQZ+yoLbcUdGVERA+r5yrH5QeDm37ECgJIjN/56Xx
9xWLW/82gkzzvsWl7R4DgH4t87ajR26x1Gx1iRJeOlu7axObz7KjqDsZglKgMVG8
jmGNaQYWADRy/7df+M+pmMDIHci+09IQNxttMNnf4fQU/9KkRODsN7evca8LtGAD
JYN+WKRtHfwbZrMg6Rmw7gs/1HVPdcTrIvfykiUBI6l0otFj5JkpkWEymyVXt3rE
CVI3Nted6q6j/bs4psrkzMgcZupew/ZrSZv06L5urbDuFiGhVhdk1aVApH82y5Ka
Ck/73opE3dio/SlnEcyG9PpBSxnpU5XO3p06z2DFkB6r/i59r9BXN7mXcWIbnQU4
Di1WrBoentS9RPBvvUAG+d/+mEtw22qSMMvGSMS1FD1L8DxHbRGyn18mwiWJX+T0
W+ZoFZpdhHMfCxJIutmP4IdQMZSnH4VkxdhWVYkFBavLGyuuOR/lHLMJGCXSQ275
1wjV5KB/n/tAjFZ3DTiVoz3XU2Ps7XUYIB5/Qo4ZL/TBcC15/XMIGksrGVb+KvcJ
3H7EbASKDvrsByGyn6OK+EChzEfCAH0vJPEmiqLK+RLVlaxdSkrzA76XAceSZxte
Dk6P4BmvcOFVpOqXCRgGURkGZ43oT466hMC286+jxIS6TzBttU76fjaryk92ZU/R
1rCtjw0/LJGQ0RvVR8RorNnAzp2yLoY78WyxJqi2yw3w64KziWkY+phvUa2PRvep
kINd2OVjsbRw97lpxi0tmYxmU0Q9+MMOoyxtNhV/UCYaRWVLPHltQeuK/TjfWJ1k
fLs80GmwbWeXEj8HKD515DD/uc16VXFHnK3y8C5KnDFSuD9GKwXSmIXugy6AAiHI
0Y9VSRYtyf2lwkMY7icywIIThoQuSvBHvRDI85r0T4eBI1zuQup2+Calpsnudoct
ZjTtGfMv1hctG2+osHQCJxfe+arxalIpekctYLtKt8RHjwtm0gyl5vnGOMv8KdPz
GgHF0Cd6rDxzZRuctE5xJaqvMMHoHQ4iCRn9ZfE58cG9otOZOYT5ZVN2UAwpPweW
06zJiG/xsfc9q/B7GK/gtD68NjC88nw3V1oe31BlykBYCp7hBciLfxwTIBrpI6GN
t3tCy+3kqC46w0bSDOQe8lY3Xqj5I77OrpQrgWIFz39djQaUCSidqnRf/JflvkJh
yRUtSZes6/N70SP0x625YjzlnPP8lVGhmicsZRjDpBkSJUJqx1WjvvNt6TREpDhF
EstAbgFJRIrXnaw/q7uTVOto0C4v9dCop5MRJbO+Bp+1t3m/k/1LHYaAOH8oGa0G
X3tMC+tMEjJnI+/rT32/pbuA+UOs3ZsBPbdIt2a4vsAe6GRnoXLRarto226D4cs/
etWtxBqvjLH7WgvF89Yu7r6lwWR6smKcO/WqnVbmsMGt1RJBxLreA2nZMKCBOHzO
y0jVGtd/bfyNyXv3nkAlmO+9lkej/UiwtyJ85dGD34p9bExKoPSY9MVpaNY/NMMB
ogndwnbFPAznpuU93X9MZA+LdZF8aetgD2wzY/BXsD25FanrhDM/JNu04wJXDz2f
qZ1WKdiC9NVk3MAm0j8bgdARPjJRuZm4JaTyhs47NL03syJv01Opfz1/LRMH9pOb
ZZuC60QP/cXyLFmibyTsEdMsPajEVnDTyIvYwG5AtEZjIcReSntTzglDrQ4uKmnm
8oXwfKmqln/bF5TmVIxIT7WI1aQvphX9gq5VeIxx5xKSw/+Gey9RslWFiQTO63bj
/6sL/j1XvwWN4wPX6PTNGwda0TMAjA+gXvIbMKsn65OUqUhExCYH362YUQXTPHYP
flXfRMfAVVAfRTo0YLSZ8KHzHrFcIU8KBTP4i0tQgVGEHMkxrxQ2qWEuV1vkZrvu
hvqB/EeFqCrTci/g6FuIILmayaoO2z/XpQKKQEdH/aB3k7kXxle5+hrJk69fXyMh
QytVbtFhHAIDrqBN66dY8Tj80CeANfrEC1I/wkpBR41ZSChxXMpQKKdoksKK3lx1
ASZt+nuG+a0NnmjbC1DUH6gnm4yQBo8Q+ZozNwhzXy+QIJilL9QCknL5VuL/WXdc
6vkByWG7IJtFyYj1Xg8QGRhY/ng35lsrvdCrzvCYpAFLyophHnW261Eb9cpNRQ7r
I7TuoQaCNjll9nfu8KpgVl2orRixTaA1TMEEzYW/obWuhhs6OxfHu7GdGVUd/XH3
pCzYPc3BOytE/Aayr6cym+iZiZkh/uaRlaPT6bc4AzCSN+u5qITmi89ELjTXQoXG
TylXj1SeRHT+bT8efir9GuaEmzIIrZEUaohB2xPNtRQk2dCaej/f/jw8g1YMpZfc
h+98TjhR98rQKKT+FUFECKyqbsUKWtwKeWWk0lz1fkQPS4Zc56jfb+/8sx6LjTKF
R64rRrM17KTuLw8Ibf5lmgaaF54fN5aLun0ynz5UiDY8m794/QHDt3TcnQvYAD/a
yWdsRCL/5dThVQ3Hc8SPhMguAhstbArQ1n0WLbR0aHQsJiOf2scjHEXGsCSSWmUx
l2cQEYdKjBRe+McuvRNkb8sSqmUrVBNpIy6kUhZuEqkSYPj7vf1pirh9rKJMdv9r
u/sT8Qrf6V/RGX2rYMePauoheNubMQQROk3S+fHf/Vc9iDgpGrgOA2EouN1oEJ6c
7A92mAJBFfjmYWnRGmuehDn1Exd3+B+B6iKc/KAmLV2SYnWIkggxPPKj4pjVHVim
wv9X2ygdJxbnH3TIWtBRg6hiED8ahp+vGRIxHzz9jM1zq1NjBttoHZnI2OlV9uI1
+65PhlJcLjZKjSuYaxqOGM1n96I6B8EVCh/JrsPh+H0XqS7TI3AbdyHRoedFq/BM
pMRZBHXBp8/Ci0Xg7iYUx1wNwU1dpH20CVOAVAlOXAMCpsDobVE9S1nTXUBCQudj
xEAgbhyjYUzT7exhCvmGofnyXWdUCTnpBuDhyO5jAlZIe3ODG/JpHkKKlpKxDcpt
xEn6ZUfcev+i4nOq5ShNdJCXEet1xx5qBMYdsBFroBi018axcvmzNhIP/SS6qi4e
R2xhdjKEdHAqbYvUapFCMiHZ2eBi7vfWloVythLTZMjYmU7CemGypQxJ4Arn9EVj
KbYDKwmjHTCEx93IOvIYDvNcElnTne+A5mYodY2L4fN5tXVEVaSFS+YaCtltSE72
p8PD8twn2Y6n43X6Yg5LLSzG2h2fxmJhoEGTE8KR8oA6w/MPnw/hx4/Tsnow4R4Y
VtEYjB4cuhihOa6DRi3cshJRX1heN1C7jo1eAIRHjUXf3hjI4DPL3NfXKHunUwhZ
+snpIXhrJxFDWAoy0IlK8amoXOSRrO6GnzM7/wkMT+M7qBQSyQnJJdXVHY8eiMoL
eG7Aw2+VhSGgujKX57pJTvZgRrt6gkZ7uZZJ/OwdiZvDKJuzKiadlnZMX6bCaXM3
Q4dvWYRJzHxKbU60t5pINl+rkjlX5VFuv1GJO5G79YvHb5npoCa5PW2RujKCVAxT
DHhiAfd6KetZjf7RZS7IjIUUc5NtZlKHjvbLcXUi8I44KBq8473TMVo/oC8YrKX+
jb3Ja1D3UQwwzmHmQuldzvBfOmMuH+8VuYNXQkbuR08MI4q2JGlJt8rN24BWLqLM
9KQZBj3X2ZYz6BncQJPX7ac4HfyW3xmnh3femV9JAuS5bzHWBKqqIOsxLgT72/SC
yHaxP1//TM47NRDmTazbwWMchahdr5dnJXV3ye2sTVLzwik7Wfznrblde09tI8x6
sPEwKDdnG+avQRwo9qjNFqmwbVxlKXrsHpOG0Ui8Tj5jq+SrQzlmqBoj/V0V4jTT
kcRxOnZ9hJ3JVUsIOizFTbJa7FXZLudDSzdt/AKFmBipdkYG6lg7HDWa6LXSJ1Vb
qZ8UEnee3dhbjR/hS7bw5ANMwH4lsLYzIEIoVqFkjCmQiv20t5IcZR/Ru3UHBNzW
d+iii6CLNwIe8use9Ts0PFdHqFYhLm35/RWUD/f8Az6Y7e48n2YycXAK8xhFaOVL
EoAllurWuLcJIAHRyTOkrHo5NJoFH9DMCq7WYBGehuO/TWFvTC4GYUA+D8s+0L01
vyY8dOmZGfzDBg7mHn6mkE5MsZmdVFBi8Xb5Pi8NnKiQq7Vs0N+DqFcugnR0tWGc
rQqOUdW4eqA7ZM2Ae44OzJeJ8b53Fr2jyVOFNi+wE0HKtiu0HwiETgRbT2ms+hJz
A9Wb8AzCmgVfPugX3sJnKmLnmwcFg2pLMWnAlOC5n45Vr57cxc+DjDN/179VrL8u
JJrV/uMSVvy+pMhMOdO+s0VTnq/mwGr16ATHbxrKCxX3vLgR6HsQz8NCmHIAcRsB
N8SBFaI3w3WSzzW5PM/y4ToT78oQ4H8MOB+SjkrmvwZ3zekrca44/305ggLP5/j6
5aLDCr1+qjffUlccGsoGDhEJKFwgMBcjLIPnRRYtw3CR0Uq5pxR+KgVouEyi14kS
+Je4iNfw+U3G/+Xf+wO8mAUMSma8RJ+uh8qIyp3FYxQ3RbyupkNVzMNDeM68A3Sl
oUnHo2/oHlLZrGuHhiHWBMytMVQkIFA7deZsMl8BDPaa5uRW1Cq+K211CLjfXJ2K
iYz/X/pigZEiXT6ONATOVuBWsAPnfTtKky7ewTZiovaMcXku+wnvi4OkIKZ6hXLk
XLAQRKml9nl9Oz0lg9MezfJzUMfC4XWS+9ZQPCdD7rhaPy9bhTcFC9V1sxmtMbuB
ZXKplDzX0GqOdGvcdc5okMsRMEcOeFQ3P5uezZl1+TkkjkLhag400aripyPVKC0E
Nz7Jdv6gkA5w3ZnoNWpPYm9Hlr0s3DZAJQ2O2MXMnfmyW7OM2qKtMc25yOCuRFqJ
I+Luu70DMWZno4pvmDt/m+gbxGbKYOGChc96FoOUJiR3wHNcFuXqhVN1B3mBJrzB
vf742Ys/hdE4wV5MZu+Y23XIkV9xK7KiqBpac+vGd/QAYPyavuOs0IF9G2hoZQQf
GR9+6v4qmLKr9uP2kcfaFQCi5JM+fZN6ZbwY/znMXfzxGBLq1z0u24P/BTguvf+K
+WBnF0av83bPmEVCVirZGlwUtCf4aCZ1UqWDkcON6CYE1koZ4RMubt1UDUeBXP6Y
K1sCeuNn9WC5fsYI9DTDQflIy/sCWitwTB17NLqxXP1Yn9P8NjIT/m5TvuMFfenu
Vpquyjvpe06aXPZfTK6KEvGcYi95umy9tksJ8/axessxouuarw6DM8tJgA1S2fDr
D2ruleO6gUHQHwA4y2clMQsz4GpMU8t1PGU+cIiKEFh47lc6WlrObwkEPRRb1bpF
eWZ1lP/qX5t4qGNTM3m7KGCfL57+rvxtIfLUYbWFp99YRSgIrK0hNbxKbJXV8HbD
iGYuU7/lk9JIqrBZUlzUC4/1NpRSqtK3Ltzn2f3JbF+5nip9hn7Meo1C0RG6HiOO
h812o3nO90hagcn0bKkFzOphJMVhS0qdC1VlMRwpiTZnYw011MAkMgGo5KJf+MQy
OJPtt7O5L0yR7RC55BheqVX8qpqZBUUEhXGe4T+XzKQBtFcvato8gdXrFMrzEzDo
q7f9Gj4PUGREAIpsrQT6BNkRX68/BFiGPSCRgHl4M+sCZfuE3ioaEOBrrLzvvmT+
tb5aAIBPoRQhXT8TDK4CMnvEB3ukwoIz8B2Nq/rfG6hq8fsnc014cr9lQ84bEp2m
0/zcFirIaVcZXETmB+MF+Ck1sdNxi2JcLVZcXsu05tGcMIZaSv7kT+jZqkGP8I46
flZi58anJPEycH6xqYxSHGGPCiCLZyGMwWO1g52Yf+sdtZ2euJqVUpj+jAS2dH8P
35Q2UFPqXbHoOAintIDEtf4+NA+g55+Vj2MAjFs0OvyzY0KOQd1RHARuThnHcX7G
NqmRtd7jN1bA1kAU3uys6WOFSZfCtKntFnU/uUuevweamR3lUukdpA6V9ogaywih
gqWPkrfvyY6jnkofUJUdqdYZj2XM+kjRP8z93k51aEebQBn6ir+SUy6imHQStU40
WU5raMQqXIF5AG+xgttFUUq1UyBwL02DtDTysoBl95INP7ganGfqbEGG2po/NJwt
j5GXse++VJ0ff6nej7N+rya3ECGmGUtR5+1o/hCQK0c98UU+bslfsh0v7VAGn1yu
5CT8sN5JpZRtT1bnrIFdHbqDzujyi0N6QQl1Z8jGlIQ3/eToOLvd2zUCljDGvSLc
onujOfWvVXW1be3TKZnEgtbQ1LM536ckAnC9xZDbqbmxeos0sL0KheCbf6olPZ8P
0jvJnbFrZdI5x1hNnEj0jSwKx7zqHRjvQc2LIHU10/IYY8cNrwrUcgnwA/L+YJW2
VsbcQTXKlJ/ijzmnvJcS2Pza44UbtTHdefx6TNFABnoRo5MDKfbDF7+CkEATktJf
EqUMJkczVmJbuilD3JAJ9B3alVJ3nv4N7YoP80qVQ19RblWv8NBGyE9OYRU74EN2
dHXSmL/H6lgiheffheb07bs8MBbvZv1fpoe8z7+1iNVY2Ba0/WE8I70JlWjyXuWR
vCNj9D3xSLNTsbVEUmQwcxeEERlK4v9rcMRx6Oyk4bu8iLTPJPub2OJjvwdgEbwn
ina2kDcNpSpjgPoLroVQhmWcerA998L0CmLfwLYU5Fow1+LJgpEkELqKFApGS8Mz
+PzJUfyNp5Tix5YQwSIaKz8PEZ4LE7L5gIBOBjjF83CpSnMaxBQ9yALzGbbpCamA
5qHS/Z6pQxvccymzlu5tgi0KYA6tErZtS6ly1KlLWuPh+nye0s2b+hVVApIPacQ7
4ZDekNx1G96nZR2Q6gwQYn8Uy6cByfe+D8eSsCXnqkDmr0/b+QHwpRWKvjz6heQe
1z3rMeq46m88avbP9LTbarjCsYviR+nE+yu5vd1HLBxSP/fLd3WL2XEeA0L7KrGi
FNF0GpoweMF5X2EubNh6hAeqPBpwjMHioAV2kmT+017buLeHNcs7LCVC/zxICA5V
MvS/1hUTXW0iONsbJ4isGC3+KXwI0FOL4hX+lNSOVgisO4eODtVBdJAVWL/Oy2gQ
rBlKsNqH3sS9g36KeOxJwDNwMfLMAEg22NQVjOboVb6ZkWEn477uSbaOxUyZUBY0
KdzCVA3vj3aXnGEwVSvR9XPfWNFGjMNajAnYOAI2rqgtNTGxVoZooHGFPMC74smQ
SBUEt+qlIqVzbZflW4jhLQchN6SE8mDOiJkhssNEpPcEUHG9fIORjr/hbngOekAH
XozbAC2GZCE5sfVuZx25Uhr/x3XqDJBp4Rpbf89xHkQVxFmfEyR9X7Ua70pn0aDL
e5MScS2tu39XnDudDjH6IFzKDjrTIsigigkaWSsxuDHaNOmsPGR9po/ersgjSAZr
nloPp6CrND4uZTRA9BXuKz0F1rCwxkNLb18a8tdz9GgSgBhh6hhKKPDW7vBcUn4y
lzEVn81wiTyHTGGuYDiZezXsEaShbOsml5ka8sk6qcn0IpMyZaLiyO6ky7hc1Edy
oH+iNuoNpImbryGT3iBi9uZ7LDaykCAkUORADuebNL49d4nr4Oiqp+3oqe9IyVtN
cubj5+2/KTL+uky1g2SlIPwF6oqI3CS4ypQV37Tfe1jMYTUtrLvtaieJ9gLC8XaD
XleWW+WofYj13uxDkG7CtKRTXUN3BIwbyIu9ZREhE8MZIfAerxKk04TAfJUwno0m
v73nbF84mo9dzci1BfVK41NLf79/Q3BZUD2VjqO04YspFnufFcYJak2kPn0XzEEU
ZVrdIUhe5WoRE1DNJy74ZQtr4wsoYe0ZUArvut3jb+D+Vxry4RHOnpArWFOxMHz3
Q3LXZlpwXgIXwiT7vRiPc99++/xP6Jv8nTjFEg2YsLCoHIss8A1Jh9RAxsMj3x/L
Cxz0c6fJXPQPhL9ztXg236KLx4+cFg8eKdMWf7Ik35jLwfbLao1fz2WKGtWQKbLB
1ZtZpD66awnPYbzGlNvsh873jjCd9g/R4TLhrcRwAL9fR1uQTWgMhcAqRCU1UBU/
E/tyXR40DYbYayEtdOkBUP9V+35DA2++5fyBr8iWX+gnloteN9fHgxkHSJFwX/Wt
nhlMg45go/+46CAYAVhFVMQIMyzZ/mya4kAEelQ9BjkVFiG6Ka2Q4BnbfVFhasxm
Q0u5a9MRQ9e4HwOQUVMyatJL54XOIcMTKFQfGd1v9SshHT6Cg6BmU0qFxH9x6ko9
wbcXpbXveCYGX2KhsfK96w56YZP/fxCiHggxFwGWbRqph272LmO5fXI6ev76erH4
q59Q0L1PvMpEWR27sq+uI8i3+5/8pQTPEqTdYcW5sGblwh/sxqhAA9B2rqyzivIY
XB31TPfKXlIjMi1EOVD6JZLplnjzorxuXzVdHBzehQHTx1hWrfY/fuqv2FJsQipw
GHz33V09HNhEUb83aVhHxSp6ZGpx3onB9Du4H4FPljp+rWnNJxmPf8Y52VY1ZHr0
q3r+vEU989/FdQZA51aAqJdwOSzOMotcb9COmSAxPfO+Ppd9CZD1894oCukOl11C
PUE1oOKhPgHK4O366UanG8wKLB/7NIpoV1w5WGyVcSAP0fCA8lgVvKbaPBqengQa
uf+PEGLEDS4T//4wU8UAXJX+Iray4t/RthAkn36YJ4SNNdfzytgExbPzV9jGiY/b
b33xNZJIr/hLc5/PfmOJ4pEqy69CXiHZyScGZS9fNu8LesVM1/vtQXPxqLop0v3d
x5d2t3ShjT/837YgOVZCTLKbiQj+liz8tjFzb6TC4kcy/vnA57rKwFz5YcOMLcGk
JrLVbXnK0OWabpmexgOjGzgOIVAOoZKnfEypiX6hb6wHEIdlnAT00mjsZbQZov7T
n8xuLjUydL8sRbnrHuoZznf5Rs0pCKzWD3o12SUZF+b/98ig6El5bCi6uKLw8RGR
vMnA7DxTUpROdEaezEoVxG3vvCr9uqjlPK6RUbltIXMAhErmiWd3pMuNr/qDVTtn
mtXm1Y0T6kqCb3x5SUZ3DawzFNCQU5d0byF4sYrGWLU4T21tY9jXrvfMr1ypSCzO
r5dubou2qnIXcEtQn6OCO/dbZq1ADIurS2bWyJ89uMoKgM35NJRbWuW+EtYT7mcy
K+VwrhRE4mj4wNXLYrXNoXX7hHvXLtf6rfkojV/ep+T7S/BnN9lq8CfbElpt8M17
hNboOQJu4VKFyOb+jh8PF3mvUN80nF4rjYLcLz0K9QiCc/giHiBnvr6wh1e7iV8v
3dyjK5taLJ+lcdTvoKBKhYSQNJb4ar2jwxPrpkR9a2toC6BVf//tCuh1CjIF6H0w
kKekI8FduOtfwKDgKYzj+n2jOaJLa9BgN0dwJOZQJUfNUCuEPOMxJta2c7EbROJ5
AhZF7Zic1R2rkH+4I+U5CZiZI7VGOCoQCryzmlN8lxX35dyW1P6f++eztiAbO3Sz
Z1U3oaxUdVOph545UsTGpwTNJRhrIefsQzBP7eGJam2sGE16QeZpPhKhWyti2HSh
RvGBajfV+L+Q1WiD3cCESqSZOtjaDwiQ4PJOyGZZ+VmJ2lSYE6tA1ryEx4egFOHI
I4KyueCtLTb4vrqtxpSnQJf48z/58pfSijUR4M9/huwuz23jQVl6uxkAvgYlkCxD
1PpY+GkOEPYUAkHby9UdcI5WXmHr8bNvSnC/EG5YxzEN3Xp8hLcJrSRmn+zo/0ML
OaB1bsii3ZctNTkLjhpl4LVF3sV83XVdIe/56yzlz3p+gWlwA6G9YPMvczIBjOWB
sEDp2dhtT+qcGHWAHKCwaJWsqVComgc5RzF6PYCMVIbZRAK7jlF2XS4M9pEnwMrn
D19c8Grr1BoAtK2vuuo//nX9JX1gRkzdouDw6fq7sKUxfRLi6ycrg8VBJHgdImCB
NbMhjm6LG8RsJFscZiZ6fCFxKxAywNkB3EmSsH2KyTwRzdMhnKiqIjJEvLEzOtRj
xX3IFB/9JNTwj/aMPU8ggBpAADMsrTNYPJLFjW8RMEOOwxPrvx3Ku2oW3cih3TCC
ggQADJVKMjAzN/EaO5mSfClK6EELhm9r8aSL2mspGBbTB45AJiDOu+l/gdi0xiG8
04XfAOsLYyrIxVAxhTm/TJ8263iUkpiSoYI4lTfVfcGVzkOFT+KaAM2A0/kNw5/c
CWyVpZ5c1DFaJEOCFSrGJR5bXpJvzdLfxjsf7BNPcYFsfhroCTrvtRqcObwiPkbd
XOury33NvKg9IlFq6VC1MLOywHfnE4+PzoxZTOflxI3/VipjHJU6HiX/WXvUw663
TjOsEw6mDrCsCJR6UjsmG2yJU679O9vPdsjxayKQ66akzgG0snAvpL0lUDELUlvF
LYtcSCzRuqJqbDDB5MQ/Fv4lRM24xSikzI0MVeZniNNTc7JNYNIFZb9ZSPwpoBet
uShJR0obgvQnG48XafOT1igxtobQcYxu3KDtAZxzYMsmiie2vPCYRJ3y9Vj3T4Tv
9XBdb2X4dgO5r8IIsQ3WKqkhI+0J2BtuNsIxfW2GFrDaaeS0OBJu/06lIhfvNOXo
A7W6pm+U7VWBza/xGi31fnuLwY2OBlPg8eXYElTyKH4g6bGDoeCSEaK2PV+Wl7SC
XmaZ+s46pEEjfJMNiudzJQfObNswgwzl7laLbJTZQv2bbhLFEeGqC7336Tw4wKfX
rIXCHoYfuTnTJQ9reK4ZVIDEK1AjsIe0m6opXnhIEIay6ll1PvvdzjxNokRz4Kwl
BbonDT7qEn7DMk1JWfM3lKNrpobnr/AeWgWtUF2fAqD38JdCAPbz/dmjcyIJ/Lfx
Sui9wMuneKIIAsufYDjQC2e8Z6RNCO/NhBASZoTGJVWk+Y6t5wJIFO1braorCKi9
eYnt4Vy8oejUA8Po3zDfw3osLMeaYDXyxh2M9ncMC6UAf7T8Qvkx58l+bs1/Dm7A
QlSdzD1tkaahUm71rIIIJRTjohQd/TpBSprMBYtvVPmvp+JggxBRd4gCZ3NE63gn
CYlsYlBQsvjQ5MW0/j9dLz741ClgKVGgzN0KHHZ1soosRMR+kwQ0lkn9cLVCC2wx
EJykSWGV3YpnfBc/aP8vaGeMtT0zGWecRLawwpwzLbN3DmN6BjHmrACoOZd8XFJZ
vpLqwXNlCN11IAmvGAGZ9B12XbcoCFAX5S0tI4+m3nQMBM7wnUxjPQpe/bKjU9V5
8rAZMb2z22ru9Wnb+b0J5PVuDH5BZarTXxnbpp1hRRSNC7fd8H1kQ50Lq5zpNOeA
+lmvVG7FOFCgoK2aOrGoSr2JOdRsplU2FYf6zjuJgxuJ/2noWUlH8SY8zfOdTVSG
VV0bsrg3fS1+OouFMnpTnw7WptmhcTV9r8j4CHjTwkf9TXmInfF04DNUH4u8Ajks
WuJp/KZtjlU5PBrrjMejc1SCQNbHsiyP0jw9esKiDERaW0oehZpX+NHxktWUWYmn
YcjaMWXyesrtOZ4i938qns3te+3aomuNJoEKymn9iUt7gOLD/5U7H98FKE2hVTq+
CTanEPpkk7WeHcQ+qw9BF6QNk+ouN/vOwDZBPN8PssHeRy5kop1hVPrmSYrD7ghA
pqAoDAxXX4oJ9IhWOin4rr99NcZnFKD1w/XUJIx3ZSE8cAGtB6sgRBhnKgFBUXYS
MswG5AXgUIOJcFSItLubhGDzRgqQjk4uyLT5Nl9GDErFRUzFrxA2gL8QV5bfLkh1
/MqghkzzXwzBOWmeZR9S52fS3yaR8xR6OwpHDsGmc5meKYaswJPs1bDYXSOjFL5y
v9SibjVB7Cz2hsHapnXPkJM3Iu2czh8PGQim8xkoVPXkBAxGT0AeRsIRtWiwPvAH
av7HBYR2h7mo7dHOmHUOmY8J5YspxIRqjmxEJlMbOoHeQUGny0SOdci7LnafeSrc
efHwGgK85xM6H9rSi3yQ+NA2lZ3yd5VyWvMRVFXmyun0ktgIcDwTzCFKk6W2rvKu
mmcIeiJ4wzzc2f2ZnEvEG9kt+VaTiwqWQk/q4kd4yLOAZRd3o5vpA5F6syFLdFy7
ZYzm5qEpISXiE6neuGsXJMxoI0Q9ADKI68nxd79VQ1yIVQCK+sEWFdPKgQkjAiDm
J1E8J6ojtwZ3G1Tb7OiuHiU1TlX91/fUn5jTsPmdN5t8BWPOQ4c/pxEkeOXdjzQQ
sI/vEwty558sgHXpOK5DYCHb2Uqign0VOqKKYRRtgsdHXBSzi4JWDxXj5tpN/MeT
G6L2IwwJtuqLs6+NRjv1ji9yk601Uer4PaSsRE7VvpyjgVFXZZ6s774ViPaKf8PO
ayMpxGVH/wiYU+u/Yxy8nOhoQvVsrEzymyf53mAod+bH/zxJaTm/QGiOz730LCVu
EDzfTIbudjxerTbJ2th06TV74QT04qa9a7fk6lsrqCL7z7/gqGKWeivXLlFHj3nZ
RvALpIMH50TVg2Kvo0dN1gTf3b9Pq7Vkgyob89KsqzFTkxsa9flFoApCSvj8Q+7v
6OvuNvGLSy+ZdZuDsszTtLwWHHhSVHj9Ekrtz0VzIsZLtde1rO2FVRsDY/qVKeI7
UoT28AqvKmvPNMAyuFEd9q17ki5Wn+vPouYMI4THaQAAPeu8cEEXa7eIh0FEvlee
6szzENGcKL3Atv6NXhmAIiRouQaWez1JMngGygWBiv5CXdxk3mHa6RbqiE+/K69C
ZXvHcqXzBbcZbjz58sOQBNxGFwRXk1xlGzFIxsqLgkKSUTqS2vICNXvHtuBZ8qXT
7IUgaOU/pmsBVVes12AWsVCpFQnTNxlxYjZOeIn/repMZJrvrAxbUnD+Vt7H62OD
RblMtMjPaWWsjR6EWbY6Nd1QAql9ix3QOXM2/NGaFsTxK8OQWOB3oZik26kocyaj
1p1fL69R/dfkOqyBYva669277YITIWmHwwc7hnHDn48ZLgpNYniBGf1FVcXXyCLx
H6otAgKPbBanUAu39oSog3uZE8WE35+cUQYj1sbqPZ4BCV4xNFGv1nirHOQHhUMk
PBl3rPNY5zgv6d0Cn5fprOrE8TI6Or4YKz0K1b4A9KRzNpLd8DwbOh0Zz7N+lYrD
nyd40bV2h3iDycl6g3jtV9aLGTblo70wcU6qa4nFOPc0slWDIMBDgkBV0roZYXfH
H/mUNRZj9oqbIwno+XIS7PXp/qlymGFHXLZGc0e2QJJQ8xv//BO2lOMWYY6+jCC0
VGLUjL2Z09W7tL/9u86nszH3PEdfgbdchsxBzGNTBKlw3DTs0vy+2szYUEah1NpG
gn75T6GKkwwctde4We/5MbDPbeexMQHBDGgH5OPrlG5kDzivAzIu9fh7QM3wt3Me
pp+1ShlTiG9y5CjWoAeOZOLKfYVygSOtcfQuFVochDm2BL5OfjJ5Q+t+ZPUSRx+P
p6C8v4KyfPLiRLIQzJGQWBmm8u+IJN5vh5Tyn07CA3k7syufwq3DCl84uzxU6NRl
gjWpltSPc9bK/b73HzDv21nMdSlaHtfkCjd79wS9rOabUQ+0cQdcyPYCTuQerb1w
i2XiPlcV98fmDVOKBS73oNb9bALtM3fECbKQimo1shlKahOb/0mvYC2f0W1SXYKX
+5b0stOhSb3dANuEORAkRJLcKVNLPAY33spWJtZtXmr9qHWlxDWwX6L2dXxthP7p
kxZBqil9/MGXH0WNt1GOFqXBaIIXH+0mpFs/3K5QmfAtoMsHOzPNuKkT49dLxRI9
WC9Pv3PMyqWqyX+rlEGTHVSn+MTup1eOU3yiQHGqJGc24UUMgdDGswkJfDsWtqRk
JnYmonrKRiL2FHrxEVNFuL+u8uP9tBHiknmZ8WAjGV+Bhx/umwWB826SmjRuYgoQ
InJP2UnI1OpiDdlNsfEfzhKh9SuMdR/kR0QQ5QXvhTCdv+m9HPvC48JsZYtyAtPQ
ZfVS8ZRJhxmyxw7UPEFb/DRvDMc+5BmpoSPgOgZD5pCnoHxiKgptJ0ppGYdVrCaq
K9eOZOEeYplTKgkLG2ymPbYtjA9AMfBx0Myv6QWhtRMSTCi/dRnMcbHnNLDgXp8c
46lCMtL+QbUq1IzXFvJKT0EEGkxD3qiTaRcTHsogZVnq0tEdtGO83uXB6P/N/z0q
kKsLsbVkfWs7EOPdvm31NOa/RgJCx0YPrTDSyTjl5YbwpJJ+HE7wKgt1V43tk4gl
poEYdLh8lAs7l9iTzyYxkryeU15sPckFkxhidoSIX57tu0xEvrVlPeCE7KJ8uqgp
4PB4zyHeEf9nstNdliiPRwzociKrcL29Oqcvs0ThgZQBTq9AH/b84OIoRZNTH/DW
E8/x3eFdCvuciJmmrpyA1yJ8Rw1QnZwmcl1tvVY9czTBcL15XIzEnBp3buT9uhr2
YJ1k9kt3K7oJxxQu1qUQRrsP/a8zh6KGr7wgVsm56EQBJdwJWT32EsXO5bhBVOko
e1gsD7VPz6Kq7ii/qcelrhGPU956nlgQzW+6kabqtnbDVmrg2/5ByzSP1e1NhUrq
LR+KJ1AuPJE06Nq+4/0U8o1cn/4PumDUflBQ8q8/7u2g/46OY6/CYTxmGt9XxyyG
Dz7WihwMgkx8PzZgWTJySJCIGg3S/d8W0jKB9bwuhSvs5tjk0pExrojiObqd6+Iv
EOo9RZM6gLFwtOU1oZ2qVEc7kczda1FB4+e2tA9I6s9nlLN4IQ/T+Z8gII+VrCRv
h/8vtNGYVxRQYQCJzgGLae5NRN6uDl9OSkZX7xLh+f2iaMom96HR/fpVlXC8qoWX
PXtmxzUkGtJkfjpOpvb7thGwd3RO1ZOuPnThjAH/rjD/3sTv2Wplqu/fK6Kbrgnd
qmAZcfWVUJAAbbLS423G9dvnODOo0ckwLw3cvOvmxCWXhb1jaPuGE8Z73UtEsIYo
bZWPl/ZlIImDSV6fORtCnYCZI3B654PGGDO8chtsXyphfAkOoSjzRmSeDoNLqtKu
Lj7CP8DgbAzHqsiCWxXWfldVebyzKKG5x299lN0cU03jg2lrLvG3btzEnk/4JmeY
BHPrbTQu074M5E5eOK4Da5+IZ45ar4akW291DgbnAYamxjYaqAIxUg0AP36Uh/ly
I4CWOZ+oH3X55O3VeAoWQvq9mz3yHKS5J0ElR9RPbsYhLgdkZf4AaHmhekaxBB2e
kPavwuQ0ZjXMnQ/z/7YzGgJfuuYdEonEUgYfYXEt4QtuZTyDrlUC98SvEo1RQdTB
PrzYiAGJL8kao/ic79H3aH5vCDxvfwabvThvZpBFrSKZOzSm2bCjmKvwcQB/3sXn
AS2wgavRsbYBYcEht8LbyJr9ptM4lng+zlRocgxAlM1Io0oc9tWEAoSVwaK8/HR+
mPGr7t6FjzuuE3NiwLdR+hFKuZDirmmEbTo4FgNwBbAxOGuwsJE3i0xxUy5Q68FT
SN+oNhP7p1VL/I1O+o6a1WgRuSB6WxNcbVbFBNeH1Az+mnIg+LEvBROTmep9ePbC
wMBjAuadCr4EBAQDWkz3/S6lsMKJ88qroIKL/Ak2NlLqAqGVjTxiFP2HHD/+10qg
rYJtH9W317d4hUVpBX1i+YY8Df/FrSDOKuAPWYT2qEoktvNcjmQABqiAsoob4NTF
hXY4711nu01456MOPxCBswu8nE3FMu2/Gq7/ib+OJI0Tx5JrGt/fOvnVuHTbr9Ef
brtUswmlfP6jdIcUZOi/TumjLy+wJYB7AsrrG7QkZNDIZUKihY/bRzy/zQEO2M0y
SDvQrZOMhq/ISUCmVDXYhw6cXrBcv55k9UTS7xHEq2lzq5vRxpL+KWdDvYhKpefZ
DPRO1PnG7Pi4vQ9PlrdvD50YmcSc4azCspAch03gpwjHEfiybQgFr5CG9C62f9dK
Y1P3va0eVwxIwLKxJrC8UkhndUQBkpJlpWONWCMIrlv+47NzTeErhUz7fJCj8sYh
34YMNT2F5xNrgIcBUHTbE6i5Rg2YV3zvsgq4dV2EMl9MtgBci0bhjQgWWZv70WMs
I98yNeCef5OcHik6w4WdiCwL6RNeDBBZ6QSbsjb0i/IoWchSPjzbT6/6004SCJr+
AzkJKEtpMGoE3+/FjMbx4rK/7A/5RJX0Q+wgssFCVW2C/pf5/gCnoBKeNMtSagcb
ZzGVRpZO5dB2zMfFoQkFVq2j9Wrtp1vMUhH59px2qU2Tg2od1UK8nnr7Gp6vT7Rt
TJ7TY5DJDQJc8H9MT96MJ7JX0dfCTyg78NUzAmVdmVorBL9IjLWxU9fdjrEKRSY/
NJSnQMnPwJqlnk+aUBHc72rnwAnp06kf+1lfyqAVevS3BQBsDzxUWEKOVpU6bLtP
jEAQaU5QBf6mv5vvyjZrvb4LVo+cwjZtdkc5mvTo1wIwEYNCzPfMVUTNXEckkgpr
hOOp/+LN4wWYFukFBraIVkgs00x0xdj3atNE0SAUvsHFwv42msvzMfYjXj7r8QGD
2n1JGjVTgSuSZGUJumO7D9d6m5oCsktdX9WjmiHyn0BpeWE8Drxf9UbhYBLDLwlZ
j0wUmecKQi26UsNtdkR19JJxxnRkhX/CCtAUPWA05wGGkA6mgRhpSOq4FxfvBP9n
TedenA84qYZEGjL+1R8IRm8Q2/ZfRtZi9fSXQ7LhEq8IvjubQULWuddIri4HbehS
V6JFTAQRXmgdxXbiEJVqDtLQNDU10FPLPhq4XNwNEDeufI8PbECBIREJ8iboarBk
i1SakIjkkSROdpavXxX3+fHGZiRTHaZT2cLy9cA8Pe+OtiABCqSvqtqslPIPa6UE
yMn8XjpnPMYgR4uzM5/2zEzxG+JxQ5xCOCP/5iHReRMGjaKox757P7KoXjaVz7lZ
X8kLaX2+kYBZLWwzR03RcY7Ld2jS63Tm7rnPL8SgPvipLKOqkL/RO+uOa9WQraqj
HDhMzGIICGS+UpuxiSWw6jaEbh93YsBatTztN+AVTxDLK0aDaEvFEgut8eRDEp4k
klYR2PCOD7i4GbgFd8zRmYkImQ5uPGZz2x5tbUV+K7833tByRAsLTMNsJeZoQg91
lA27ulrpPPcR7Axxvhubd4CWitN7WTXSSHJiain1V95G+gmdsN932g+uIWxmDqIZ
wQ5GDVXHQX3F4/S1fNmbP1Aneu5iF+fVbTPmxF8JVIRsEy8Qy8iWskqnfeTPt9y1
bvKsdOp/RlzVD5MaSB//8JRG/+uwyo3C1DN/U7h+qJYTc0yHgLwGGaoncVBVB819
E3h1gSORBT7pT/zHq+beMsFcgJPJrSOcO2DRBgmDbKW1bHqaG4N8GzRSSSCDGg90
0vC99lf8jIvcSF3f49ST8m2GtJhmvIb6Dh6IQB5x5HDO4e3rFjWqNYzHunNT7x1H
7dzRAHpTdqhYxdylH2sOBaskFJ/tjkneOMPp0Uw+gkTNcOW/sTiDusI27Izu5cfe
LjTDfKGRd4PpYCPS0byqjcrjLUqxiGKSYScNblf+wdiAiAzLVNHUinPxmnYa5O+T
lkSBTFre4xJaGT71/edqjgIbsZ+I3F5wzZwxR5tpmZmFVp31Yt6DRvtpcNdWwCWs
0LrSSqVvd9yi4mQkavOVe2c91LeDBXNiCFJAhOHQNf7Eb6tu84bZY4dIoL8Y6WmP
0VWrtcFk1jzsSYsSnJ1awSEcBQ7WnPWdwnRldti5vAJ8BkFxxKxMJqrtWQBEQq26
b7+OjGi74uv+KmXx1y5c0qwccprp6nFkluSYNjAUZXedyAkeDjyNUAUULFPLBMTY
6ODnb3syBth2FXRE4NFzV+QLKwMWjvGlJTsXOKHr60dz4qyNSLY+A8wjOULWSt2S
Kyhwa6pGbd+ChfMlUbr/gBbUODhWI0f+xq5IS1fWWCWYXdk86GglXyfn/7Dqoxzc
DBERUHSe6cdeKl8Wf59xquRagKgFcjFCeq4p/WST4q0eIM3rkS0aIZ7UWn0HdnwO
EDlnVF8kwzDpIo/s32YyRal3sZqLyhXc9rz3PnNOF7kp7mjKFfJYhdvmyNk313xq
U10tJvEEvWpHe7AyIBYlucZ1i2dIyozq4eDOMAn6bXLaHG0CdogDXwjirmcfOBPk
SafDNgzfDXCtLJz0XLgDSPvyf2WGwqfnM3zVjNMbuTDVhLWPJfMiiQGe7qJgcWi9
VMvzXRT1eeuPGBSxyjVM/6nVteR487bc9efRM2Rn0ct65j1d0uweqQ5EsCXecHhe
T5YVp/a9BtKunBwfRJlCDUVdoWVRM4ouOzTSVYeUfLdohp/jhebWpCXsFwJPb7Fm
5fNm4HwxqEGr+HWkCLFq9eL2/GtcUrQMh312WHRT89feRNIaN/6U4k4GG+2BDN3P
KMze8rDr05YjMhdiFPf8NgXf6u3n/+tYwNymHphKnYyeTMuAdVCBmGi+B2DRIihV
U3VqXcO7RJCvyU/6FpL/bk5QeniiqmGPkdYlLdynjPO2kFDbWGcbZUZb4AzFywMM
tVjgkOGp8futy6P7FZqzIo3+1FBrovuU5rf65nkLIn2fgVG8nAyarPKfyNzvBdbO
nE1K1jKRguuRm4gr7P3PvoP2UJWUMdr16OL//nTDSKS9OBNztIKu+3OXcDsYy88Y
pTefsqborweWL3EqXYpZ/MgK7nFKtguu3ZOUxLe2KX6JiJFwqWrmkoukBvJhZEo6
va4hl8IQkFTQYuvBaMAOfLm9Bp9qc4yc6SLUwJ2EYA6Es9qsSehIKnuTjK6duDNw
lxkKhcOfb7SgESAmNaNgRYxbFq2wMSVhIqLQa1qDlYiwwPvTXjD+M/szyd8Mc4DG
L4itPy0RJmSMzEa6WW/Rt44SVzHXbdNssIhMsPX99zvdvqUejOgMVkBJ2PMUbACi
KRGoAMKjbKnNTjB5ABCDMvKRMsOG6zUJ84kqokpo21QoT7Ya5NdOSZ3b6Z0fkApm
WwiM8N3zibXc4nRUuuGAuZ/Eji9Pn0ElvFA7zvOROeHFIAtBz5H+atV1pvh58Hjt
boyMcjKKU+OFP/fi2vFdVzIrcljdm9a7c28cLHo7oDsfM+VhFHxZeziv9LP/m49k
hzlc+71xZ9Mmz1HoKdeX0ZQm3F6Wh8K90/DzdxRk1w1/sKWutf0pvFz879hBYmtq
K/q73t9s423Zl8IEI4GoWQFgCiRjDgAt33OuRTeFyUPkhAn5lpDX2w4XyCH5bXwu
/PBVZtThEeU/9uF9NByNKm9x3C4mF5CmvxIG2oc1+YNXwpmehGLfz453qhaoM4Rh
jxEnwP2kx4pQMVFn2T15oEyY9rd5RuUc5nHFn35AzzrCmQiMsVJ4cmQ1o/6RWyNl
NgxwBOjy8AO6pKUknLVgj+MJrxm5iOH6wIVBtyAOb1OBKPWxyBnMd54kVi65+HgQ
m/qGHcMYcFlJMkYOx1Ec+OwCdTT3qTPvAnMeNpm21MqllqAxRiMzDQrTR2xPUSKJ
By3XCKTAjL6aAhzlP5gK1okhppRBKILtI8LRx0OaBfdZvORd56gjpL/G82TnbZzR
sTluuk2WRoM2sK0byxWjgYTfQKJvrKayQk24bPKZm3KNvk1G5tb6nKLV7LZw90Pv
GoGAt6TuY5uMlf+HTmCNdvL3Z45Xj/wGIX0aA9CJx9RcjNmTj/YSs0vk/HiXiTLh
IWZiJp5QKKmXkYg/yRkOl74wM1W/spnt7xGGQanjNolKo5pDzmaGwqIaoQhnbaLO
cq6pk8Q1/OWXeYQ7g7GaiYpkKc8ZveaGhIyQ4nlNoWaCN8wbaUFLveZXeHpm5INZ
syv4ZYw6PqiALxv9wm2zGNq4pywfK2n8HquT4AlOLAZ7ZSKqqqXMSCn9lqIDYc+d
l0kI4k6v45yc1rguUM40Am4a5Bi8ldJjTw+oQ/ry6WCrj6UbG4E9M3St6pAfVsd2
/ZJPV5VcMp90D6KWo1cgwpLtEn5IxeK7qzK5HrTD/J9mvqVFIpjYOjsByvKvuw13
gicwMAhoDBURX1Be7KB6HO6CM76xKv01OZ2vMOjSMIXZZV1d1+Sfje5EjPVRaEbP
UBXmXKl3rO6V8jN0wmnCunpDJuzSYeTzYA0f+LaMbTNBX2sT4XlIjHAfCWhxW5JY
wviuk7lSf6L3CiEtsF1lm4HRhqxLE63a8RhLtdjxjKk3lv/z/a5lUSVbVtTBf65g
Mz8eIu+A7D9ywhnPRAR+68ew5fTcu2glXoBm+JDP9hHz4t3kaNc8Z6YiGRrUHF0+
SgWETNIgTMzJ8FboO+wHxvVwjPbco0i03wSWuDP+TxNS66KIMZOXq8F0CO8vJjy4
E/oZyuEY6SVZQebPvQzPD4ntDXkz+L5rzNgcp4phVAoTl8yILKDBdl/5q5VVmmms
LJazBsWL+d+/ZmTPSyw+APkMZCbH3+3tZc3RGHiVzc4lBP5LKcWLfDW+ck4V0dZ6
CAhs8WMa2DXXKocP9YKyk6zA1dOHQ3PuVVnW+mccNODtFfyFimv3MV60JninQcIL
afEdQpoWLEDUv92ROlX5JNOV3dCGaz3HEGroMVBQQuILqIi2EiOXNbeWK0Gocid9
GoU2Hn6SfkCY+DlulvA/FzMxyrmMwDy1NNbaYuT/kYZ9ZC5BKlayN1zipbmcZ3Mf
h0lgHzhBXqCpNLlVQXfPZV66bpNr4QGUd5VPIeoZeG7bgSw5oCRjUB/sM3yHJHHp
Itel//19NRBZgV7dWAfoa95yXRnvwP4+JRh1VdEknds0F1QOufrK+GJNhaRqeOwH
RQwxehGStCz1l0L4SykBZo3h3uvffHtnpshClMhiX90Geu4x1UaQZPf0ZywXtnJO
vBPF8T22QNWMSY/ZVJX41jQ0n6KcdQqRYpYxHz1VHXTyPHQ056/m3RKDmz9JQGwv
LYp6Tq2WD17YcmCtioJ7W+Od82d80IwFzfkb4HdhHJOKjGClNRXFCV2emQYR4ulU
/DEFo18e694BXvV89WpgCm35Zw4lGLx92JLPYg52fFMmjecbUpxQYSgFyIZg+rtG
edeavGxAJq5hr7c+c/yLYC2eAQCgCJNuBHnQA943emos+pLGcItqmQl1W7KWCHsU
wNDD8q1achIdvWYfHsgEhPGzTHRVMLTYwookObOzqo4i6/utbvN84PPNxlokUKfl
624rNS+JA20qmOPqH6Qq9ytGct4xveb9kKrS1vcpqdo6l2u5F6zG6jckTw3Q2m4U
pl3Fyv6Eca2Fj+VjBB7PbgYVZlCuo4CybZfbUA64TMxtbsPAN/s2OIrhSddhJoF/
sNcCzfT2OERkNwHRC1O4B4CXdSxe3FQyn7OwqEUI6eXaZghoCJlrivzkgzZ824o7
cMCGG4IDzjferF+n71ONBRb84HrCDM2Wu5FNRTW1606PhZmle9lYw4CFV4WsQpYz
atjrBScbh+W9a9R5ePrFSjz5TVmmltotXQxY7LPNXRomrvye5qYYAYvJpIxS9OKJ
ArwTtL5XHNZP3h7j60tkB1Hx9KrC70+6w7sK2rDplbosE5J2qgTJC0o/lPyxKxCo
+YQNVXXXzz8CgjgMN9hzkczClphjnxiuH4TxRHvrlLenDCGxA0Ft0GT2Jlf+ZMAc
yIVpwbuidw2fdqn846sasX++xLCFGrRmxVxL6J2q26gmqYHbDrlrW4lfRoYc+1lD
rccL18S8eUrNx0H3an7ObB2o/mw2AlJQjBd4InfZe/+FXrItpkw0rI/hitPREwYS
MUa2FGEqAOxCu3SZTSB4lpoYvpQ9wcYGengI1BZ8SWE3C4tXXS+bF50Dttkv7DaU
qaaDG568ENHcaPwnNtuFqciewE8eHhuJTGZFnegJEddC0r/znQRFJ3EYvu4JABz/
9geBhbv3dWBU7o1tvZVMZ7NAcYZxGHxTuzU+4lJHta24w7nVZJgcGHx5zLeIsiFw
NaCtuwVEsuM14HZn9w22uaayHtYEDpXtcC+4d/lvLYHZSQjDba/0JkrAJuOibvbP
QYy5v0Bkn1tUDtMuo/PFUpys/hL6WNghOpmYnBawEYDnM5Y24JL7mf75iofRcJ3H
YQlEFQPa+5uQCbsCSati3ghFmUtqEJKwyMULTPRDYAEt7nxzUVrVP7KqTOI5miOg
TFoETDJ0t54xGWjqs+75uEkiPpBqWQ9eMiqlTp7ODEs9peB15tHAMxa6kKKJ4+pB
2GtutQUJbcCElBtGxtBW6t1VIEwzDEUS0clXplIpAZjrzrANodmHnPzvnm7C8/f7
W8egjIeiKmARkJrrqyXD89buJ16YMp6iGa5CYESxjF5PELpF2TDpUDSFvkrOkp2i
S3EsMTVsizKAXXKGlhp1hsMKaiBZd7Wku5WaaqxOudHkSxH0lzApBdr0n1Te84Jp
0Kd00wmUdADkDKUWroHJGXA/3OzN3n0JLwVltF4Bq1y0tWE5qy9Fy80ZAV1Jhjcx
4Wf48AjPTgRc2Vf63O3Qmg8EA7ssRxr8yD6hhcGYytFYBJGHYepL0Ll9ETZVVVQI
zeENHLklSMcMQzi/i6O8meY663egZdxpMIKkrXkCD6gq7lxMpGDoZOBYi7mpBfoR
9MVw69eBmXP0bKFLKkA8g9Ig9IhpLJReznYabxPraCA3ftyodjjvGUh0RqzXXVmF
4BQb9feg8rwxxVxp8Kdda9GMoo8KzJK6h3BRqiLhpi7lS6cgjfzXeFijqtkUlthk
nRKJr0NMOwChzksPA7/8832fPiwo8i3D+U/sM6mWj4c9bV8mKuwBaqj6CWgYh3/W
midjvjBQceBTSk0/uzaLU+zxltV4b5FTskim1Mqu/FhOK5gjImiJk/OvPhF3Ldh+
OqX5/m4fK55ocg3bpsfuJPzZYEHmHxJHkGdoMK0qktxO1CqFe1f/EcpQm5QnDncW
yL90qxVUZ0M4g8oMR5l9vzz8qVQiHVpELLjpqLk2i3InFGl8B/1QbHevchsYe1oq
okqCoP1doBVpX/j/VSKRYLR2E/MP5AoHEqHU3nNli7grQUu3zZyTlCBwHhp7pw2f
pEbcjQokVkn1e/tSkH48sqOUH1FO2W8PznSAmSmVCLHmhFN5BKtnTfW/V6aK4I+g
Y9UYZM84bmJJB4CS8BTqLp3/djMVP+rrsyBJrkKiYWyfz06pbijsdPa+fDFalDyw
eycAP5MtTJFmmLbCBqEruezoXhzlbs86HBB1f6bPXWqXjgFhod/YWz5hUaKVEvSa
zHBq0fEKYqwffXQVaKW1AEHJxu5X7H35AHEz1ONNPW1BKgt9hvQHRlJaTRXhsFkn
vM6U8sJYqrU+W9J9szXdSkXZcb/DD+YDwTb4Hf/LVQuRBk0rGiDbh/J1uQZNUYQ8
UZUDkiXA5DGnE0L2ZKabuymJAs3DdzlN57I7nYYZZLr851Ns+evTx6NGHDI3qBU1
bf5QbUMspXg5tY7kYCmfWVBawojcYKLFcCtoweTqC3L7fGjyRT6Da2EbBdyvXnfV
b4mfMq6oWU/glibBH1I0VRLlQlMh7FiPWJ0tAhXgCY9Ld85oKa1pj0BwzA38tnXu
Xlx2i+KAnc7WUrlNsUPfiIB2qFCH6sRKPtf7uRQYys8xQ98461XTWPIyPj2Ius0w
E8sTqaduRe41xSG/bJREaHFycAtflWpSaUYTvZhchvrImk/gbqgRM0jdSI8juNct
ygUt+rJzNchyOnTr3fBay1cP9GNnB1ACOIiTrcR4W8zgTbMf/pSfc9/EmsivFKC/
0OzlC+KfeLgR00fOVRtulIG0Kutge/cQw/lXmg0SOHbaH3qzcYj7LI9S9+j/OAn7
u7taKcdZI3avW5AYDguLiAayA2++2MSLus3gW05LG5jbEyowjtzSh9I2j3fz3juP
34hr61wiTPRjdaJ/d06ErDw+3xUc/tx3mQNlr5vs+Tix5wNhuR4xvZLAAsNYBKW6
iJ5RC5zvYGPMYXhDGFb6C5yUoAB6JDaKigQ5U5xgaRVrT3Y8yPc0Gfz5jeWJoXqI
LGZxqO16JU8+nRbK+VqSopkVuXz+XO6CxdWyJ51K62SFtLRlpcAKVhdY4gwSWxVo
gbEqxJzQq07K5W/BT6I8PriiiiHfrNlhfWKAEKPjAx9Buo+E8jz4ysJYa2aNAvyf
hkD+AMYAPm63mS1I4h0tg5xkoRPqcuJVYAJp2dSE8x2Z153axxwTd2gKl34wdnII
psPsyesNdHeP5TfLh6MmDzhOPwUEzU1mEZ/3BztHtUs6pDxMp0dIAs5bmdtuYsOe
P6ZEr5pxvSMBtnt5IP1v6/UfFBKPv8fG7atyLJ1Vu6M/u+inYU1d3tq+T7S5hfug
hGdeAQiTjrVoT8RKRr4ZntRI9Q9yjeaXqlM4QVSNad++Ohggdb9USnjDOBtA4z23
dHCtJro5q2fBuoSxtQUrjmi8cswb556gsm2M28Iwk3gmZxXfNW00lrqJdJvCPsb4
jcu1LLxtH6AdcpXFEpHqD3Azyjgv/UXitUJFl7zUqgDz0PlOHloioJAdBXbAhfoZ
oHfXO/PGsQl2TlBS5Do4OvyTRu2VgK3k9IchiUlCX54Ik4WBOuP+b4k0b90vsz70
GSviwUxPbOCpr4nDLqabwZC65MyqUrj22vTMHWe6/gNqOU4lpgLPuaRUIPlqSX9q
yEHXuEzR0HJS4NWrCEChQL9tnXI3qYjTyNirxLX80yoIq1wFbeM3xXlwCqhRBXAW
KOPUDbZGVZ0ZHGUf810pIqQJC25Yj5yCYCMyvr7pgSw62iq7g4BLpq5wsHgzU+gl
VjHVRkyIuPFflPhHlihtQzAE2M3aAApHMgxfpR6LilayCpO6lXZ5WHd1ynkNAQd3
Xr0GR7qpJt5CB3ooMMWy02RNpO9NuVlbeUD4Da6qiGEsE8D+/IYvKNOaYtPxAzwy
jUad2pjcldIcb/DnOwNiEd81WwpB9km9GBh3e4HYc5w75iNnA5U0YHxtsXLOuVmD
IRV1AEpKkIXLRDTqkCFGfgcRZ9A+7hxcTopEes52QB82Gk61D0B2UqU9RRqYhPoi
CENZlhZZNICQypTD8qb/WeINRIfyKBdjtyMBmJWNR0jIVGfqStv0jFgAeglapiya
aHu52mpMQBpVICzi48c9EkkZyr1kSd9RTxu1R7mkhHkLOU//tIBgM8/EWYlPIdMd
ACXbH7OQ0x3xYpgiPeuSHz3VpUYeDPIvNFpMOQDBnul2jfaTcdwRRbEI7FpNaP3k
kEUvyuxlXB7ojGWSJQ2kzXuOUkFD4gaDIqSa5/JNks81Y97Nh9VHU4JSMMJVk9wl
A748on8KMPSCQ0pLlSVX/sn0tEawpglmRQ3R4x9hRaPWy7Kne6kVZFkHUSNb8zA3
/louZ60bl0ti6EmzvwItrBu8UmNgPH8fAndqvpjDfdykn206GkY97QziQE/4cIi4
VxxjiULfYcRrKQw+YGK7qFtHZY4g7BH1S/CT6sSS4tUblku6iMKGt+nKd/stGmbl
tiDLC7tMEoZVOUpvkxthedmTUJUC31duHTTIcUSzTKVc61O5HTJZYtIQ0ZIP5e8W
0cuJ0xW0br/vhAOU4gfxYZ6ozj0WWZ6/QUumrjwPjyBY1goIo2wmmKW899h1Xs7F
0wl3F7nSZPFpkMjpBuo5Z3gocbT/5sqKi290g/I0hLZYwNei3t8NvefeKE54UZ6o
8WUIL3EAMiZiycShJ52H691lP9KRcs4v1B2U98NRf5lnrxA2lJoRimFof4rsnwYQ
j4C6OK6fBR9DqqNp7Tem53v8nYNLbyWttDZUu2faAfgx5b2jau0KcRJXbtXgFvS2
q7gKxaEA3BSVN7h3Nmuv2ghWIsTNfu/cG1J6c7W+f4PYSGg3Bc2npNM3Lj/ml6yH
btLmini95pU9Gh1AHbu+5ZX1nl6ighUjC8BTKRwgrdrCi+MvUd6Cm2vIcMGYHaUm
FtUevm9aC9qhCi2rMw2vefwuBxlpzi0TmF7u6rYqZr77BdOJT3v2RJJozziaV/XK
e98opiamD/XxmwkR+ovxylbqE1Qz5sKY8y1UU6N/Xn4ed++NQkHrJt9bc034nxNz
SGy+L+P7coHYamKgPMEQY1VBDj4B6xSQ+jYfJwfidXHLc0FhIbgT2KwDFISpJZJQ
QMSfYkBpi5b0iqNEhS1wRsV2SBJ4v0g4gJLqaYwlls4wH5OwVggLYWqhvv3DjISQ
MCu7EfiezTQKKVy0LVQEjfcxJuXAF9E5lsLrhqsGWl/pYW9teKvsHCXAD2oWQmCZ
U4EzeqjWUS8ni4Sc8tL68Vu75JZzaovGdTWQWZh6SvVmhKVgCWmutUMWSDJX/Mag
1jw5MXP6uIwGds2RHtKjDysGmp2HmrGYOSamk9hOaGCRcQ9cZOytRmpteGI72r2r
W0knY36NEMdTWscdLNa7UOmbbhr3wNgvW6Z0wD01OelcBF0AAqzhbHVRiV0jGY3X
ns7fzeBMjtYbWhxQI+HS5jDjMh9igfBT1n/f6pMqJvcz7eyMO3bek7cS28h6VYGX
3FpsqvA+6u0lHr3UgTlbFcPEf1Fe35JCN1wLWEnhlPzpw6IhhzWd94t6gVD9meSA
ErrxORr7Rb1mU6bOy8yxZFWTxEXiX8TffKEseqAyzQFFUc3gFxkEdc2c5ps9KrqT
vMc/1K/w4IjnkS5GgvVQ7yblLToFkRwmTAemLTo9wmufNvMI/Wjrve5h4pvqoS+n
OQ+X4086upOy2pxcuIZ8jfg+y4zpkcm7okKty24nQoGgL6p/UoeiWrKXcLnkeyFK
XgQAngJq3JAE6VzMc+dK79pKFALY0eWnNdoqnLopNykypxklYq9XZBLpKxmJ8avG
hGG20qCYbCP3ux+bCDMnt26J1P/V3Me8qaqPWH0asVmZwsM4tGJuWtQlusx/OHnM
UhofeouA16LadZru3OJQbDxqDNTRa1nzaFiMVQZl4EoCBUr/oFbA+oHHoMCUbu2E
8yqzz6KF/5ystHBuEMyWi/pnACFmzGnMmf23uAsWp2MOSJzrXnjKxNZg+eM3y2sI
m+Ah8oRGye5wKTrN+Oi9Y0UMlUelaiKbOBb2V2u4tofV44i+3hR88Ek/OrmwAHgm
7g9f5C01m9pWivPbDJMPSrPfZNA1uhIq1lZzR4bDpF9CdPwb5I/mu4YewNcgHiW6
Lpp+qoBDlaxDyx75J+004eqLUNDQ+uF96031x00VRuq+cqyJt+3pMaNbZgKEQWPM
eeMUHBjz0HhIKZfd/AS8lUbAXRdmaSQOiDR/9IAzF1daaR/Db1j/fPX3o1G1XyvQ
tBWQ65q09NNd/0CLmuSSXcDEfntJ9LWHEh0OkmxKuaD4mwjg/VV32I89wkdnMrqU
EhxMtsGGCJlZ2uZyCcrDLlcO5jT16WRunEPHaZQtlTB8x8umpqT2aEYVvDYSXE9a
orA4OT/gMGL8akm6K/PW6WcIiu56fSEn8xrJvu37uFAIk2ydDU1BMZBOM0ze1Fz3
9DDnWCRxZpGaenBYrpy3K6IDVY6UWfav46Da9eTWa3+2hhnW44JYc8V0+LpgRem7
88WP6SvTQS1zr4HPOCMEJUh4n0+vIm4o4P8BEZwYWze2Ifj6bTP8dlJqQr4O5Hlm
6q5pWMNNvh1Xv3zE2eRDK5mwGpzNxmuuoFoMg81mWxK5bmtXF5USvnQEd02pc2SX
i/5ZhmFF4AbzhI3bHdeAy04KTrNtQacqk1u+6b5rVpERO6/UDQPZdYEgKfTXJ8da
97IXpwIMjONEfyaEaMcdRB+z2k2DMwTQhhtO3gCfaIrGQOE4Dhivg6Ww7VTjhGls
Yf8R6IR6DfOv61vf9dvk64YVz7I32YsEHVVN3k0eRR+pWw/7Bcqpyiinekzc9IoH
MjquwEh9sw46ElJXxqy2FhThZKnqlcgBPLaKIhfqeWz2npufBxdG/E+Eer6zg+VN
2tk5qEVmD9U4fhTol2LV9utDYuh06uzIt4hb/mGc4leXAyVWFFRvJseON74t5JWQ
U5C/X2EjAVVHx3ZDoJ3ABFSg9kZ0AH6Y3cOAIdykwY7qE5GfVyRlZ9yjnBM3Rz5E
BNAU/UMOCCdFIScS3UV+yBaGpSSijxsSKCzsJkIe8xIWXa62ZVxDijM+VVfiUzsA
ayGab/D8BMJvpBbc1JYT6ozZgQvS2nH55iilM3PF09yzKmrZVCAhcVB3ZanUCXku
SkvM96oJhzBZyPkJANdJ+6k8TZ5WXlAq+htu1bmplYV+OeJBQYPJSaIUVkudwIOS
hxArsMdyrB2RKUnlBsUE3Y4YDoVWoamN6NDp+U1qTUK04BKLokVpBGK8q7AW51vt
xEzmTpEI4PsC+8sMZEi+LVhJgNv8ICnDYZHi1FsuIkqhUOaeWU1naXyEQ0CNSOTU
uEQE3BIuDAQ5YOv2huH8DqmA3zl/7xaT4sqd6+GFs6JxH0qX1gpjeX07zApLZ5Wz
mc9kIfXR/MaOVTDGeyemWXJcXRl2NTYfdCdEcny/dHnQvreAzBgScReQDyn/IAFE
PCNcapocualgSbT/11TprpCuFGnTU7Fn/TgWgpvj6X+HtRCoakuRMk4Rm+80pIsP
jKygDnJxVVw2IHNKmwfXRHK/S3WX/3U72F+uT5FJDdY+nZe7uGwpZ9i2mtwB51/0
Yhig4F6oJ7NBOWsWrwrReZrerH4kckF/gtVGXfh6QW33FUXHhp80f7ygXvIRoQhs
Ngjkx8SHcqLsXewPBRjAemvMWAwhIn/C4VDw+KsYKnOonR24HenDdurIFOnb4kDZ
63NfxjLDC50ZhSW8p8PF1Z4SqXvJNtQ0kO0PtPwlw69svT7niUH8bgYNZeMQUAJK
P5rCfHlw/nHtKBQFADpv1zevhBzy2JMFPF3Y7P3H9yriDUwATV/rRgZeocIPe37T
JU92Q6z6WAPdLCYwssVIdCUdSZDegleb5KAcAnM9JkgDK0lTlJa31lTW+a9XOogZ
q5uX5QGhG8ANryp9G0PNQRo9PBN3YubhBfWoW78Nf8Kbzia0Wj65IM4meq4yAK19
SFmnqGI/WuClc/4nexOGq6zAiM5seZnEiDV8DwaJ8N9QPsPzzI1U0CDAh9LjsaFO
X3qIeG269tORX2ki7xJgEBngpm8fq5WMfhaUpCesByOrA/PMt0fX3BcXbccCmNBH
rAdlFfetU0UT99ckJkqZ51GHEbAs2ikrWdhjOCasDSUQBnLbtvcmFW6kHY6DuMnN
LIvcCIV/Xp4lmPEuuHVtVCGYr7IrS+6CCNJI1qJ3gY1PhZiLMg+4TJQTu1DpQCJN
SfuHyVbt+TIIuNi1UHRFh4vfxZHylF67QfqISdE5UZvCZwAEh6tll8Bhp53XDifp
EnFCOf1fONEKIXaylNl87EsRKqrqLkM8H9kwDwLbn8OPw8Aho31jiRVlm7tuEyr2
FRKWbYuFcF/rWcwrqLWel09FxdW63NDKlv7Z0ccRp+eLymSUjOQ6cQ7IhRzWAP+F
2ho98QH6sSGGyo2wXwsFxc7A6sh30fGPUFF9omBErlA=
`pragma protect end_protected
