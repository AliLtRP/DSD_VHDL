// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
tUcn997Nnda03YRp3qmJ9iW+UMnwNlN3CNRyji9KXYvjo79/ZEUNuofX2wgwg5l4DEnnZxV802q3
ERJxX9miSZJUHMK7NfCMY5f9mexjUbueEUaNGFCCjB6xPRV03uU0gzIeF+pOtHHsUoGkPKlD4Kfw
MjbhKCXuY8U7fb9IpUTiKahndTlqt66qr/DXWToh9hotXlqNbDRJ4z7k3Kx2lZcYb/Uh2GMRqDtm
ssl/rzrW5vfmaB/Un6je5HNvE6wHa12atsSf0GcXTqv2kGmHJm3P1epQGQhDKxLFfYk/uv2h9eI2
EawfqsSVC5n0TtbLssKjpxIqzOaClHRWC5Ax7g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
qnFG2o/OhZRRyIf289VHIMvQDuZYTd1Xqg/TFJrdE2jBQPIn0/BcQPmJo5Wc8rivne8JjVTg3hxA
9vkYu/WqazQ/gbU5u49Kx2aayAQjQW+Fd5P66EVwcQ9f0QoQhEkHM5xM5cNYC0FlyXXBF52l1yqd
IFt4tuHxrxEY5R8OW2pwdSXJbv9Aj85wsZ5q1ukhx4b2q4330JS1m9uRR3/Q18a/gB6Hmj5v2W9U
Oxsxst+3Or7a2W9MHFC1QXK5efgnAMXDXrDfB9lJV6uwVIduP0NstGmfOkwlv+N9aSzom5ANFayt
FVaiRirVNFPRxSk6/tnQYSHs/O+F26F/3vbHCgwoIeDzIJBDheMI73fmvARZgeLmQK32aE3QoVyv
tfhQ7Mw50PMib1OlBh0ca4S7RyJHZ7FK6sc+37TkJ/VwPzl7crMJOCxbJ4NrbxL9PUZit5NLmuS/
wsQ6gfDg41aYt3opyGA32++5BwytGzyZNmf2aCl+7KqpH49oDpqoD/LGdLWPEy3oNLUbaixR+mPI
gByqSS6q8ki4QZR90Rs5bq82wbJhDfLwKZhC08lPZOrtXvC+hTIAOPvOOOU7eaDyQZus4dgwMDW1
4AvTjkjnvXzJ3JSPdre9pPJb6LvyumcmKDJgyBigJuus3X8m9shQpoAoJmcuVTTMxlOIk3bGe2S7
gc4tjMd52f+Jzw2oLQwNc1+pjdquJ9QRRBdRpS5YRKxpIluRGc8f/WjTSXOj8LOk+ZWXBLG94+v4
WtW7ItyjIxC/BjqTujGStm1cyCe5v2jf33O9NB0Zkv1n5JaYjClsw1AhwqGfSb7w8PoiqUnhFbMl
5CfSg7OOJ4sNcFyTWpp265W036DxPrJtGusmHdUmjedEPoxQAy5mmC9AS94QqTz52nOwUY+kZRbN
KZ9U9ovVV4AylN9Qz3Ij76ovEr1j0u0in9P4MOXyq/h69tjA4Oa1J55Y7u1KkLrOxAeIf5XMt/Kv
FbSRl2TkJT0RfJPRf846qUQoEUse2oxqSoEGsb1epE/u5I3GWXvMnWFMRxRXkgl9tJiehAM6hMlA
cJGO+bOYDGjD4GyvudpB/vxxDvAlS4k8o3NTyca9Q6jRcYtlm0TDI/ctvJB/31EjSnIdRDwvnCfw
OrrlEUiJdveIiwNcHY+cAy4WY2+YOwIkLpLZ1b2jgkOabL6B6mnVqiMGB+eEeOyChrmIYcd1ewcG
Iht9hpMZkxhJlY6feFuVc1PwOi3jeQgriZIrC/ScJ0lSvJ+ylZ5U0L1p8aaUHhl0AdO8+cAV0CYq
9lG7LiWCQ1wM5ty2q0dLJ0iMU9eSruK4D1wT3dZ3FBPbzO8HbED/Opx+aGNy53qcyY5lbdqzVX8X
daHff66Rwrqpg6ubYJaoMWHx+WtRAbanCh9oRLrPihk3zMC43ugC9M0+1a5TQ9ce4KlwrZtVhYS5
cHjA05sAEDVslvch0JIG/nBLSXLSV7114xEiH9fcsO9nvR/XR2tILoFG/HRyqM5g92rbZw4wJbsa
FqW9JBTfP+miaSARGA8wqdMAyG/OuxeV5sVgTxeWpDLrJjQ526g5G2B51qeIYRekM4087p2rqLdp
tqrdxgvYTVi3w3vN6o1F3CtGIlCJkwgob6km5ejLgktu5BLqfvBv8JXQj8eYeRr8kDl2JXI1Fjde
OiN6SD5NAHpi5cK9gtJ0cBCxeFoolVwGJO0bqEc5gjjFwH6kgMqvQswJQVC/MKHSwmTRPL2vKdn/
XPI9ckQwj+rabEJ1bRlgJvm4EyB4J4XhANdKqZPFLf8f2RpVSaAvIXItdypOPbukccZ+xYLsqORS
SvM7JwMhPdAVTfxrqPjrldupEKAoFpse7hau2sVFu/mL9OEDLElRtRaZkKRx+mPZfANe5/+sQ1J+
q0acjnUAHj7iU6OyzndM8fTzKfylUcdgjk6wmLMvW1gMbEq1oS8I0aMCpdN8NniH9XWzvyDDc6Ez
aeLkxWmDQB7ycD6MOnawZQ/lSV+eRJIV1npr5F+yg6Av9IDgZfPFtKefJ8CvJLxI73fQFNV1WJlv
nHoE8icf36O3fF/HjB93Kqroc9MkCLtaGonPg6XSkHXyxi7iU/MmDNfufKML10jrhrVs7xXsgY9q
t3c0HBasJYz1hvmcxnb6IGdnTOg+JIg6kFGtKVfQ4lkLgjKaNWdouydz34LVZHqV4R4GyxzBTibo
ESOkm/TEn35YdM/OVf0pOTAOZTPT5EsSty1ipB4GN453zBylnq0oG/LSpY55rEYg4XMtnEjL2uNw
W2KzMjidqcJgBft2iUAx0f1FvWDaDkafpmcF5rJrRwTz2H/3vptyB/LQcSABI/qOpqzy8UcYc3EN
EbJZQr1xRWAiwq8k1RtFYtP7ipab6EZBe8z9D0COxLakQHp2J2gqpU/xwiUN80LXGA0Pevkzjw+6
apV66JRhk4iPwSGfmjHcmXwLS32uwVwnf6o6mDP6Gb2XI1SdgF6pAe7LKHTZYqEGjaujfSPLsB4X
xKH2jPPsd+7+m9mGXJ460411/DlbOC8W6hS/7oMg4XGvm/Sbj+q4asPX/IDtSBY0eSy+jeOJ3omE
OW1hyAymjfdyCY7u0iZdh8H32MJQItMYjeJPdi+jHR29fQ9r0HkdPuZ6893Vl1lcHkFrHTjKeYNJ
kyGG3ddiPqRqz9ubCUULRwSHvGriDD/eMCQ6c5GcExRYCG14iY8zVD6OiWnSxlpObgnlqEA5ScrR
VtIA9jMSHagdNvbYa6EpFxuevVqCu2UdR/S1xQ/67Ojgjp9u6UOzR19C6u979vAbZ6wcr43zP6dv
+Yptyj3fsn2k2GbN6H5vqofngef/kruyhGjBDbJ6NIkhT78abjYlcmQ7SyLLP+hnkwYKGnxNqkWM
Xh04Jr+sd0qdA6NH7i3tkVOSnIm4rqPKVNQTjw71YW0NqUxREOjWhDuetlLMqpSJuzmEG4eYm4oJ
E5D4yDj/YH30b3PCTxkBzPCEmhTfUYt4KMhJRkiWy2eL+OS0/+XzQBJwTLSB3nwB7JuYP5gKw0Uu
hWlUCb60WExnhqME65VeRoKLj2rUhSJJe9lHrPy7NY9HraCCOHJVDsvjUbDDKmbSL8hpAr0hbjKF
kdJHTkNcasDNtjVQihg8pK/UDS422/KzU82zZDEGx62YqR+BB4RfasVhvahSBKXlz8pI7Wabq3F5
2z0r82p/m0mqmDClrUAb783Sa42XZLgFdo6fKGqLts3e3kPkc+ucYjk9BKfU3UFJ5sFcELca7nVv
w+/tb8rI7suG8HgHlzQIOMWs5ffBGc1+CE5eNpr5+myntKVXoaRKo63YSTwqeAf1rFCjPOE87qI/
EahJmsB3m5iITpLR2BeMzI+QLuy3Ya9h8kBf+cRaJ2c45XHtvh2/ZudV9BEAJI/mDGmXUSypeVw/
PQ5+bxnnfTX4iPFRn6VeLgAjcy1pNeaDaFE6RDf4Rr+hBcJdM6DFE/HTqihUCYYPTnpzDYNFANzK
7DAj2DEX8e89MfVzaX1tKzmFN+5oAcctNJMFOBW+8zodv09ELOtJ7bsQXvVGB3jZaWzDq4p+79b2
CHmJLPr4KLzAWtLekHIimgRyfMIDs3onLWlKilnrmLkv150pfn0l+6WJ/tix+A4eT24pfsPVj9vi
E6g7BYBipEBXBLJn998VqB+ezEviFY/Rhyd7k858uEPVYgaeauwjiwiOB3fn47pSpB38LgGlpjuw
5mOrnfldthhhxbrpxkGB8jPij1Ue64wgnxLYOKub8nhWueFBOcVlXx9wnWWkB3FOSUK38SXNOY9G
aeBIBiyaRoBz/ls58vuLwvd04memfmYO3TMAzmi0zHHIx7zoWmNF63aPM+HMmord/VrYbLMAA4P/
TcATOLz1RFvG8COeZSP8VlQzJ97DYdg60q4T/3aC99UL2lwnfLXPiggXusrVDwYL3IGHtpslNfCY
C/3Gk1jd7CR4P3opkJSAfYVGTBx/nedsNiyofH3G0V7OOdSQPXoBDXoLUshAyGUXlO0tu0Lb0FxL
L4KAAEw3P1MMVga+D7yyOhl7Fv8RsJwHhrHk+a55IYIEnQZe7WGgxwVmCMZsLVtShYObIw2zJTTu
Bvr80KWDaFA8goAJi8SaXi2gJxmhkhyX3aJfvUWUckns2ZW5jOSk8sneu+WtL29NEgS0As7t/krJ
Bic/JswhyPF69Hdk8F2ZFac1n0nyO3E1Iy1dDn1z2N+Y6u3J6eSx5no5zcTSiNDGAOK8OG3plU6+
cwON1gC924eHxyUZRWFFTnk3pxMQFPTihHL9hl3iydHsade/N8QomoTw5dN7tS3nfge+CkjJmV9z
pX3MVJ4FyMjLXHY3VMtgWw6RaiHooNacJ/V65uwKxzHt/t1jnCgL21KvLBEp+zNcKWYVxO8i1xVD
fRePkJ7QwmrZkEWzNnE4gxvJG6kxT0i2HL3Nx5tLNJjm9yiW69WOSLifK/mequlyVrmOIAEWYJAH
9D5PVPnEtwTgnbgNz7VCZoyiQfi7sLra2nCGKiO8cBDtjVeJBT7j3Jiw4bTQBTdHQDYUmY335HNh
yMT8vzRI37Iut6fn+2UjPKEcju/KSoXxjkfrVepoFRTgGt/7orDwzFg6hjRHrPKINJVM5azptiyT
gSBzGJNtLTPigZmSwkxvY7XNdHiLAOZ9mm13lcIUhodaQ9AfKMQn7qrhRLn2o2cNRu5ml6OgEFnB
rQUs3xGzAIJoWVPMQ3rl3TbiEwagA0oIfH4RAevI/l2ovTyRNlcf7PQHZtzfK2VL8C1bLrtXCS+N
Qdoe8Y5PdxdpvEmZdfHV5Ehnmi4jL1r/32h8gbk/Z+wnnL+dljzsC4OdxZzdUGsGXsoKTVusSHwi
YKVwHL/PY/xG42avViUobGy1rn1IOuO8PNWL6uERX/UMBVyfAaxDVeS6GR8NnHmN5Li28fzV7L/V
n2isFKd137Fftt3UkEOkbNKDrL6zKqXEZ7/dvIGmCOlBeB0pYj8+tC/o6ydU9EAJTWELbFpFewZD
hxZmabuZ5HlTpz4ffvQlPFfuLB6b0QYY+AumIiM1vrUfyCiJ0rMJU69LmSP+P9TYzDlS1Yc9ou+q
a9Sjgg9a38p0piBeQO4mv3WFdg0V1A3HC0zOPauLNfhm8iZF6ELQ0u2aGHqdmuUp6Q07zPv5A5+I
t66P24NX0o0Q6n6c7wMNX6AvPYcI9E1m4l7HQdneUUgCRzXGFBPvpBrvM+a5ce1hurf7RBrX7lqA
YyUAneO+TsJoyJeZcmTdPmrwpbU/GJ01jwgMCYpDOG4He/5TbL5v6k3HUgmHp7rkvIzqpd9tsZUi
tUFDDPV8FN7MJXetxQnn/sSDe+/o9Rn7BNM4aBxw2475AgFIBhi/aYAvBNewU5Yfdv1FDpDT/R41
Z4nD84w2k+QhcCZ9pD1E4xfEnBDEfF5844NnHjZeW7dYBTX/Tc5gbsNed75QpVh3q+obPfgwKsQr
kah+BY2ZAlrQ3i43PcwyG11Cel7rfWKUFuEzwtvkN8IsOU7+J2fzwb6/2/cu7MIiIjINyvL/Axl1
qy6f/fqyS0DfOeR8hJo+Z3al8Hh6OgY4R79sGdtCEhJ+RSfSwKhEPFHXIKXOO9VOi7Y8r1o1YLFA
niiah8b1hnmO+T2sZ1GSbgmGa4xB7mAxZoYRsQd+aU6MpytKaWNRMGUKESMiriEyc811XNEvdXg9
HmnTEW71mu1hEwgwZkAsFPuDPzj2cFZoLYQGBYyYtX09hR33oRW3WZqgc0YOOiqChIyjNmpQTK1D
YgacQsdsiPN5/rMW93G3vp+RUOzzSWWj37QLsuLYM+PIQY4Kor3Hez+21HMFdaKuFvRs1P+eXt7p
OxHynkNfHE2CSyBjIC0T56d/QT0RYIHIqJ5ICssTjMs4usI66zPv9lcdAF1kAkMYE0GgqEvqwnrt
BgZdIKPCrCL4FxftguaY0QfzzWTIFDXmillIhGR46BtZUT+69J91NI/kpby+saKWrmlDeZkuuoM2
3S4KuJ1rDs/pXhCRWWSPalmhu7kchnmNGBl8DdRbNjnYVorVYIMT7Nm17aXRzXFgZ6IzskqplZqZ
sjdx7GsTEn0guChddiH+SwmH+cYXouQ/IDq3y4SreHFy+RiLW2ViCk3PxqvxmDsZ1nRlU92OZpze
7qBNAqOSSStIFNTcnshXL5EzySPdq1Crp3cTVCM8KwcNjHA82HJnrg+NodJtvfDLzMyDnUVsAOnm
tf6GAcUhtarjlHdtlgPvrw1fjWgmfSiAGR8Z4e6oIk5T5KlAOgixcQ0BZ0j7Yu8Fn+9AwsaCMiZR
Oc7co6+lKf36w2bIiT7hnCyM9tDS+iRrJL9Yg47WOndDM0ZHTuDOPPEtCTyV8ONnUlNNGg3+nggE
oRVBD+n9elX2Tb5OlPnwNo4O2s1od33zS4YntPefcU9B1Y3ljRu/BsYq+zLKLLff0ONXPT4IW5W4
Qx7TcsAG/hoIiVL9NurusubGFrNQZGNnNfHLAQqhIVut0AF/0OciE507yDe34NjF9siSUYN9gOuN
YWxrshX9UeiuVVPWclWnILujksKxUqs/dZ7+mCijUqYQxjrpbSyabO2txqeENUBlLhpf3cLKItYV
Kc5rqbJDZtXngQ2VymEueNhUa4FoM56RRjOgppUI2F90Nqc7i7h7Og7ymaiRVBzUiHO/ZiO83s4K
TJqnkaQq4iKebU0UbbEzPtOKPVuIrkcg/PiZqbRfQWgkrxvrgYP5wFV9Y1hprvO7lC2UO/WlAbAN
pSNDpNTYQ72fXPZKTRe2mAYImAH+ra8snGWBhF6WddFkh2k2EJoHqotbodD3DEufOeOHH/hIIqiT
9G5N9mWr7ZpJnBX/SyoSVWZuhEsQ7dC4v+Qd+ibCUB5kXGce7Rcw6rpuvTrEEoyhFhXam31expSJ
Pcbd+lXSgiYjdKDsYIAHnEGTrPLsHr4/wUXQwlRwo+WW6jd+74cAjOQiGu7W4KAMzGsTustiuVc0
sDOccHLWLJuIV4/LkgNVWeYER7YM+4gz4Dkf8v4ddK8ChgcWbdHEYTGmFGvueqeB/2ZYpV81Ku0e
mu1yYwA9satc0X1QyVdQpEuWKvu788s3IYPbAeks4y2Qrs/GwAKLu8LTeqMNlsJwULqh0/F/w8lk
2ueacSqZhQiDiAu+HDtQPXyuTankXJQ85+LeOCd6FoEgPyiR3EGwqkYCM5CRWDurVJ3JBBzE1SUS
n5t01ZtZCeYDXUZ+x2ikIjJqzOrNsUEvjlufhDb167KBGOVJ+ltj75prgwefqFsxEW1DA0cGF8np
CdUwiUCQIRz9eCxf+V4CaTu3qxc5AvsrrWsvYWimsT+vQh+l72x5mbhVmKzi5nNr3P9o9W9puMrn
g2a/YugwwHxArieuRrpXpeIb/qq+0BL1iTD+sp0mYcRaqqEI0psIi5GaXxcj8+mWL12ArHkemglE
o4Ll0hGfXmaqykWMtRRqXx1B6Lp9xTeUzufUIwDX9qkOzDAf7SQANrTzAEhekI0IVbx7jIuzEWCd
Vzlb6UimlOobmTFivryzbtpA89kjCgY8sc5+pvqXPzNKUbKVhaE66sy4XBAFs4bM5Ii6iqy6FYjU
vD/tvEmLhWc2B9izKGIv9R+O+57rLLmiN5qPEQJ4dulnOkEsdeM61ubTH403kis6eq5T09VxC4ND
s9w6Zi8zeZVg5WDrx2fS9jdt0IEzO6vfeVyLjnnJvh7UKC9WqzJdyHdkGhp0nXg2aW2jLy62iHeX
N3Kv7+asE30MsJTyttzlavtEyeqWOb7Io+C4rxtdrvtJXbeo9BT07FH+zleT2KrbmEQEaSv0+ScK
VdS3clAYjvyvRMIIzcfq8Nr8f1RpmWQ5CZXRKtxXREzXMLRSeyq4gikwOZqjE2mP/OxHZalIeaXb
nX+zwEgyNWVfM7d8Vwzu150tNavBflFBpAGpXsASGAxdeL/g2RfVUuyMQ77iY7OZv2i9brGK/04M
hVjwq7BZ6bEOVu7+KVMIKT08xJD5GE83720V0zo2X/E7htMV+NJ9GAsj2DOOo2dSjXu84faXl3Qb
vszs/G6gk7i4w/9aRKzBrd9aRnES/sfbP1IbhlvPDCY7I/nBipnb1zFLF1PnG+EhUMlCsTs+481V
+ZWdLFl7hmMxeBxpTyHzN+ltuu++4ow1zqiN/7SNQM6Ezr8r2dlsMrT448nsIXkQOd7NeQougvLq
g/8TryJ2vBssIBqCnpr9anqKnv1WXS8uUXKwR2Xt/YYK/Be4mL3YiATAB59ZnINvWvFbBdCCT067
57UJE3Mx575I9+SQJRzCxLgtLERc3q6fvQBzNyndZAPl1ddW5iHOAW+Ae0Kpa8QLraypHyfvxUOj
gUGqYCLYtX+oYQL6gjJKYTxRu+NOH+yfif1ab8botPKW7PVpeqvE4WL7VOwc7kj0MstQwwW1jijq
SPC7a8dnrxIQ0s/crnivRbKv4v5jepqnlw2dGxmFxNJhD+UUgCOotDXsZF6eQY95zIFIdBl+YCGI
GGBOXZeTK4GBYdRCwOip4dvPmR5dNkCpI27U5W46smGIFKfHsLH5TYQOy/lQ4YHrD9QKxkZ84ZJs
5UDz/wU7BBOaZ7yAnoKE6nEa6AelBnf+GckthKB14Bi99HipRtRiiqu5iSw66AYouGrqgC592L5g
A9eoPFI/Qd7Y95C80Dsx0MDITXhv6fEIRCDg0hpYUky50FDw1+FEAWr8qomebV7nywHw+gcxeGdL
mi12r/l/2QGO2eg7cMPwAJlcuGQm9YLIt3P2Aao/pMY0H1pN+MveXGOqcrb2DuRafr5NNse20WMn
i0SU31950q4clAqFywb5yxnFEQaWODEeZ8dVlfEvsl7oupjhNbqMS/0NAOGZPKOE4eT5aLBNixuL
JcxpX0C+LX2MMRfdN4ywYmohOR1AYKX2W9AFPWlEu+6fQBlR70TZgahpVvtESaK+AS11FQEXsuiW
TSJ6vQBUa2bnZwIRzUiZuNf8dfbEzQtgQJ7ZNZMku7p41wH+m2USh4fDPx9nw3pM96+L/i2lhqQp
g62AhlTKKQLCZ8EjxXehFSPPG0nKhAFII8KMgIvs48eDQ7AsYYfHSBXAgCZCvheUnO24Mcwxz+8o
MtjYe5OK73VMN6fsmyT6O7bP6mFGQYKn6q11OvaSn9EaPrYprjsV0Q92x5ySCzwL7yjpTqaPg0l+
ue7f95UNbxWAxw59Zdb3RaR8OQXd85BG/r7euonWDzI9rj2s50zt/wGJPGnnFRWcq5uoEEuyF8bX
+T1fCpchiJP+ETGcuHmHeRuAYw6EWXhCrZmh4+jVXUgZLTSJ9lB8098uFq85rMbU3byBYDQX3BuD
gnziHj88jgzE/2w7vCYGViooyBUzB1xrTD0NmeGfSIwSvBQHkr7c+UgaP7Rx7ymnA2O1qYk7lm3f
FMqWLxngzfzfs43ipg4GSeByjyrS3eOSBYvNkhzmSSqeD3R6SwO05QWvo0EYPpUbXufH4msMXDdT
+RVal9odyv0Qr23i2h6vp4b6gqaF/BL7EuL42RbH7JXKVWZYMrIxyGfd+wxx3tKhbJZ5BkttAD1B
dbAoLSM2ImDwbc8h23+iB2ygnyu+BIZ0y/1bfNzQUgM/tsYmjRtfW+bNoUTZo7TIeyFzaXmTapFN
D9nW0Y7sgH2IYbEVOSEQry29l/JRnNVlumxQgRg/lyfAraoaJ/Xwz1D+gPaOB9GM6SyEHxleOf2i
n4NxSznLlA2w+X0uHgyH1I9rDSpO08PX5PyzmmP5LJelQImxh/Y9xxmyKY57JwB/zbNesEP9Xqs2
sHEclcxnUEY5o+TGXzfsu2+rrRAc6tcxfzNlUJcFUGJ2zFXantihISt0Xrh/uX/VT0EDBARUtdZN
nHET00EuZUrjdeekjFj68zcPUQLs2iTDh+92Yi2Io/2vILUaHY+31wBRwttHk0UoU5kukNqA4xZ/
d0hd3MEbjudib81Sekrf4LnUFKnnMBbo6Mogr90Py7/Ms1Jni9n6LylhANSEuO5zq1mYrsXYc7wA
uoKIBiYNlvicL1/4E62SfT08SUZ/2l77PC3NDfSrUwabPqOeSybPJ343bcByW1WTdx0oodBp7mi3
EYkHaucvETksaaoYmf6P/7o02AnwAWgMi7pBxih7Zd1t1KPz9E9vjquv/GxGDUySz/dJYlGwDMWZ
ghbST7h4jnZ3AYalJTmN3N+y2r/aM3RGZ/LjXBcH+ot5zgQhyN2xLGUBnV8z2DnsprLcMxh6rC6f
1y+PheH94sT6iTfdp1QnmsbywNaxwiTEFV/4VRoqzZ0tHB81QmZUh5A/ti424reTJ1wygjClkf8R
IuKCYJ7b1B7SWKPso3by5QA5sy3Vs0oyju0rER6Qfmsn83gSReNIKdq0cYpe4Ww4gsgL2m+bClst
rlEv020+nffap8f2wEax9dbAnJcMkZsBMfsrDGMSrVA6C7pF2ge6fI6VgjrBD6hRhTlg0VEICDJU
jiP1P+CWAhjCW5LdZySS3TwhY8sBY9xXV6M4t1PEfnFFe1nlf5nZfrxvlBpEBduUcHZYUu2O48nO
dbaJdQObncvOiokSWeTxUl0wTmt5rizsko4PXB7J9gl1T79UZneAjfj19rAI2VwUhn420AAHHqXx
F5a0oVSJNtlvmIrR/E76t7qOCgq+Px9A82J49uvLDZvAEqIYGT9RgLmiTxndE0X3LsSI3QxAJvSy
9eYAjVodjj5FOfU5UmLc0EeqWP/34QCpsSjlqNU8e1KGh7vlDQ3p67BBUaPcmb29x23Ph4ld6bNn
/C/P7rz3WsitUsMe0Lnz4xiE6yBaFS/FYWTc01bRcQSoeM6tOgHFhrP3llidWsgXRuhJ/B+uXLnO
kd4yjsI5x2MxUtjB/eP2BEpf/5ICyr1HKxaQ07u6KKULlk0jbMD3MxWwFiSBluj5QEJ+ZmpMkawR
xzQgY+tsT3q2I2+ioUhY1I0R/JQtD8OI6GTZ9N22kA07VbbvfA0SPnAI8SWkRBybl+aqWUWTqelb
ixdpG9NaA4iq4y1bidVJ5op55Im3CunkKkTQgiJOJM9BVcP/4j2qvPViiXTFB55nzihcG1hKggly
oTWZFaOM1r8MmwgvhvIHAA3eAGr5HuioJ8tqbCsZvWxmnHOqcYTdTZjaazDu5sb1kfrGdY9ZCPqE
/le4GoCfP0AkWFmWblqYe2OC9PTlJhAnJ+0Vd3roIk+zKpimJIOA1RxnXoLsiwIJ+SsQwOUL4ced
kvbfq3Lo6xyGfbqDsnl11p4E4paOV36IoIW4CZ3sLf6fr+PkBiaWvztdOZWooVL8PttoJUKlMYgs
SrMKeRQl4OlpnGo3wnufmMxsvs2tYXKHPWpzeN/koMO2799dCvreUcor4bZjtXtjtkmj7+CRQ5IL
o92YjMPHG8GsvophesDv9c+PZhdP7AOxcmHCU7PKRPzXKsi8LU2Dij9gze/rFSF4bJx67ArTxOzL
cIWu8653+4hvFlWALp1JR1FJq6d/Rw9SwZu67gIvPrJDhQMYtqHy32LmiQ+DGVzsuh/84F3fANCg
gQKYNuAl+n13qNQDs3AkRYznuDOBNjXFivyZ1NPyVgOdkH+fMQuYQD2uRy47jsGWFX7ZS9jAtZlo
AIKudnF1TZsZnJ+joJmJCp70k4lnRcipDgsgsik85xzaMKQo57ZT1PBNQbUVl3yajbAiJWX8GoxQ
lb4iD+bcgyRjwn7mYkZthUJtgLk/JUoYeWC06GgZM0LFyeFWMpZRb69b8C3QYKVBHD64leijF8ya
yMwGmmn284bebw0fJqeapkC7Ag9wt0y3jteTTOs4iDaMDbDj8wtHgRMcGTd95jnNg10Pqq/CcHh0
fZ5jmX/pa6hU04bYaYrE2IIjjF+tzAZCUEYtlev+NTKeijwEp2AZS2rIBIhY138Hb4BIkXQDHjVq
lLl2aBavGT7kIoGxFDrx1qeG+B9RlJgDEMVJJJed6gNMHrBadNzGuK1uGkZ1Fz21SvZ8HxCJQDow
IkuEze+UelV4sh6aUBz+iz4C671i5LBclYnERAhXeJb13rsx43vsGVHT6NL6B7a2FWjfGQh7QrY5
EQQ+OzRq3DO1R4OeblWnHa6+ZnbUlkzXut9OQyMf0serHWJYsZA+atagqJA2IoFmuWlxX7qWjirw
cWuVhB3usmOJQH4vbCkX0Ll17Sm60GV6Giadea0qiFpHRVq/wObuS4WXO9/L4YR0OEHlHhY0+DZI
YEJxnXMWmd8yzOHU8X5ATe5HcmVLJYGYYl3HPX8dRstKMoeJ90QmtsDYNuf9WBSw12Tl7hVExumq
XDmdzbZYpwbWjbFKqDsSdhR5Fnzziz2Uswz9UPRvBwKgD0sQ1Mzw/i/7Ev7to/chyfp0xgDFBhcB
5cM+wttQuIMkMHTXA78RKupGmCt0bPJtHHTfY6iJWRZELdm4QU8aRA60PQuWBdlMkCzP8ZZ1OSGt
OIOb1kazKansBKtKjM+6MQDgmwsu2tz8NL9q4KqObN4iAqod/AtSxWMaIigrsC4fLCJAWPY3BiDM
0G+EuNf7bta83yd1vpedYm9xuKYe7POK1Glzd9t4JTCNUe9wP2o5BdPpZB++f2MWATXv+KaYEW5V
3t7wbWk7/q2akTH8ejyYv3snSaDR6o2jZylehQ8v6nleXucmQIbKzu2AwVTKdbwoXyf1vJCBBKUJ
2/+dZwsRXj6fafOAXf/xGp23WAUSGUCodhtEhhGTVwvOblea/PsWq+sVdHMPKgElAD5z9BofCZm+
ov7IOimhFxqjBhUmpfUbk8imrIjYxW/Yam2db/+u1QcSZ4MaqY3KqWLZs22kWZ7eS6MUk6wUtWDs
ILeLV7peCodSDJM0m2gjx61yNsv/oM9zBw4vP6xRpgY+eEa+g3Y40l//tMNYooZNtltL5jR7Id/x
CM9HrjSZ9eLBVi9hfbzRHK4F/+gmLEnOzVYfzDXm8ktoMYz4D44JkE/L5J5CcSIGAxf9JTArIkNu
WK8oQmwMwUcNIAirstYVo8e9vDyESxB3Kgy/WFmPwjHLYuv3cB/5otQ9vBzB+besn7xWyjDp5aKJ
7s+eY+EHr9V/4qydu8LOyQA1DYClPrdTIsTVL3jX1IVGldnLCdzRn0Y4UQXVwrjrlFmscWULXPHX
sPFI9RuaVhPLJc6uiz1vCBjoTq8ozxHTupXndUnP1kS4xpGtdBjkAokHqbDY9LEebSgIfPd481rM
xMuZS0RkSTGqy79oA1dyqu+4xO0qmA0E1/M9gU6kTYIyVBzr8KFI2do1Jq80tP0iI9KCkfhICiqR
/smSSIgu5yjUw2aUv5CF4fhbLKvAKlMeFymFDMpts9uA7tFyxGlCg9JVMhEK4m/kM6loUGuDlngr
b6yZh1Z2654VmU/b2NFjSV1/aaaIapj2NIvM5JpYxzBGoFhnmOqa6LAra/cYuC3C8fKm4sITZLLX
A2pAMqq2JQOCby/wPW9fQtEDiqY5H67jHP9u10VfPt+QDbXtYzi4S0Ynf4fI5/O9Oku6TJdCN88c
CsPhA8fafk4lBHm+AjA6h/q+RmHTbZrUIiJGrUJXXcpzOfcHV9KhOXtn6U2d+dBJE9vO4a/I8tSx
5OtaBxy6ZUN38/9l4rZ4NrG4jX9DQOisQvgfTRsUHoh0CNnvDHATPs+NJv5m/BlxvkLnumwkXsc0
COjq8mS5w2z+dFfFYdtA7wl1497KSFI5xEvuh6MDAZdBrs0G9tYL9npb5S+aV+zrR4xfokR8SbjD
tapvphfNbvvNOI5nOPDy1FjmGcGNlpmt00mmHmSD8k91q2vQ+bm9UEN3vCrA4ilaE+UT50tj4B9v
eUNT60BUmLQ39+a38NBJvpISoAVltu50pUmVtKf3bzaAzLIe1LY4Sp5JtS/pU7TCmooPGiH7syPV
h6ZxMOjL4b2Uu22QrjxEAtWsIq5xrNuhtR3DMMI/XzV3cbYoY/0NLdGD1+HK6uEkDz8Ez4/TGWyg
WxhrD6YvOUqrMZmg3I6VgSjxEAHEb1jfaxwrvUrx9bn0XnJAvK6aEK/bfhExQW/O5E7PMyCbnvc4
/lXcqd73nwvgjNbUbE5NIj31Botpjs/+VG0KQwxOdYUFQB3tfBI+4AR44uDsGekrVrn/OgoJXTEP
zuT7a56T40+pED9weecNOST20t8eMz1o8bPYUfYEy+ogVBTRECvBdbMVGSSYW+ALtoS3VXYG/CUl
jFhnxHnZUl0FB2EAwH+PJx1w99k2C6UvMp66wu15zONZ8hUMDlOdi9WHd0+x1yNGuGkodi2G5EN2
UAYQDYMbXBCMVPQBhQZPuz2s0d3zWx+xpBVK8fGpMPJ+OtEq7x7jTgZn3sKF2MVUs3Gj//nZy/a4
rCYo2S7IzMUoj9ZxTVj8IrYwcvlKP4RonQXt490+dtuXnq9hMOfrLVJDYetNFp0PvzQa8BYuFhWt
TF6v6X6Ua8WGQrdWxjZyoaHJUEikL9HSx7/EFhp9cf/h/r13166pe6o7Flj+DYmFrNYumoWm+R6U
IMzakQtdyncJizZzNNfqq0RLYhwbmCGajYdMuYCdXHaJKVOsNEjNS/5SJ8QU6Q97Oq9HqA41tbQL
PpsvThPNQUjN4QDXIyfE3xwjiTB6QLtuaIwjH5P48jp0aSMtYBaJb/ptvAoU8EGnymax+dgQd/0X
2D4zbkM/7zJ/KN4/JpfB8Oy6MDjmVMMBqOvR8TkjA9I88yJNJIcIdVKWZdZ+U7HajPZjXmIxYHKD
FfblTJJteuir1FhEtX10pfiEWpP6Rqy8RmLmC1gnAXX1m3VloPLno3FZRTxEIuZyQdkx450zpGfF
hat91wD3xdxG2CEhgLo7iODruceIs8248KambrfZ6zFamU3cuN2vZw3Ei/GuCX7IH/Cl1hAc5MF4
6cEdCOv0pGONztYflJjAemNe2vzxvoDXCj4534BF8SUasp21fUR6aFaSlAENgDcFlByN+eUYL59T
o6LVR9m14FZ9DIvGqUbvV8bwQK7yNRP3An+hj0AeQvJllDstVd8YW4sCrclgXUfFOc5jRzC5BTZW
kwTR3ZBwMNfmIAXV+mbp/AB0cWfNZgXnVCR5q/7tFTreU3vU5YsniLX+9SEeen5/ybH1yfUgK80n
fgSVF/8x8pocai11IFtsZI0WFPIekh7TpcHDGsOMZ8+HBZVqz7Z2mW7+OIzbJBxD+B3Y9OYRTXAn
b+ML7rpKGnZ6X/51j6G/8/X9oQTSwclBk1ffv33hAcdplZ9v5uLjLXIYd/5OxEpqG8bFxAaf1NMp
yYuSWNHgGfZ3qZLSgJUW51UXRtcyaYAFSrBi215bY9ayyjqlvqGpagBp5Dx9bc9xwwFotQakSxbL
xDBnE0XYxDI3XiNpZay44RLCBDrw6SyqoF5WBpHnhRcQkojCAIkuUO+zfZlBg/K6kbXu+E9etoEE
vStVs5B/+gndL2gselApLudaFybounYmrnsiq9+T24cj29LdwN+eLv2JJj7KFif5SEVoagyGHQY8
dqZK2Apk2xJx2zNI/BXrawA5C+XR9gTIqH94ZaVSWImRH+K6SdqRukQWzQhSo1fUod5MHJDak4hV
8DfqJWsWCu6WnbaC7TWrz1khamleb6SD9DZ333tfXPL5qz1mjkFeLwf31YZpRWpp2yhSO0vDEGLo
glOYXNEd3De9eVw7pvOOB7hqK8ddKpHNJy+hSWc37rzNdrm/vLzH15asSoeMyf145gD1O6VLWu86
kVdjRnHVqIkGXbrdOkVmJDtZocEQtSQVr14QiU3TjURat9U70x9JUe/kz9cbLDYNHI7a/S/NqopI
7hLZQ1FOAdrZ8rkcVtwHGCch/UZle/8AHoyiygkhn2vIB1I1jO6IZ30IBu1VO4+Gtwg9/3JopxP6
Iz0aeHhtNVVhDvRC/aQZ9O1Hqw0quGSUCYQdtHpzvzhvA6DdPou8eIDJTYJaSDgcEMcgwpzXMme+
Hgf3HwU+AVDFysKpx+68ZSgozd6J/R/aDpnkSwB46J6BFIxlQLIkB09PvYwvrP4G8zI+6ACcABTX
ewtOKwRclBhAF7k7iade66ZDMuZDlzLfeaouGxRhUvfv3AtRo39HZvNBJ98XCEnHsEOQ5PSm+3GJ
C6fpUE1Haae3pqPBTtxZu2CndTeUtxZFun5ojAmUrS6IP7OXDXdSqb/yopERmrlB3O23xuhDOewy
d4bWJGQMk6YbhYrcmc+8cbEVQLN4YV3Vus51057Dbc8DQeEf7Pw9FUk5rLMsQDaKNnH3OnG1WuQ9
GximjUeUROIiVoml2tamYHHJ9bW70BwL6a5ifj221GvObSpdaHmg+RycmuMfmNEpg6xUIXWIiNOg
qsqEXRWzQkCQthQSKcpsttvg1jn7/uPmI9B2Rd9n90+4v5Ry4vuCANpJZgiEamRP6mMX3hAwLrOb
cEDxJEevQdLe3gYwZI3D+Rxxeh+5yvU8QstU20t4PPqsVqsGRlAmJE9qiAOvgkqxUHcREZNr2jW+
alNIGb83vy/0PMe0jVIqg80iV+D7aim8QChwNC0Ucwn2WM1X5NvUBuxVBsEymvLkQ8Exeijs8Hkq
1d3sgiXwzIWt6kv5/ziAQiWL7SYRJQCICocm4D5I3lXekp0fGZNlQA1I5GIfFk5lJUbFubLKu0E4
0KlzWJR7LMxpJeAcYFSyXI6kEGTjb0YEFnHwrcC5i/ttQccWJyS9xjFXnJo5SXXDNH1H9RXtmUeg
2X3W89YKKO70Tg/3HGwHetSs7ywWYnSvSTmI/vehuZKm50lCVurRbz+uy8pqqr9orh10MJMrzaYG
bQrzOxjh5K/NWyUx53EqFhnkfr9WVxREkiwQLQYY88ei+MYqL72apUBx5yrgP/uxqw8gTVCKnGXO
his/6AJhU21UgiLrbC1i4icw/qry9RS8MSPiy3C/aod2rDCdT/aK/lRYXZYS3eqi0VlpHDma/xgn
DbbS5t410V+tLAe2y+jxY466Tws37KT1CzNBJXL6W3QxLdA8s457Hi6cJHlwb8LoB+BoFoIcFdq1
5DlFR+dNSV5NUiWdYRYbpa/UnvyhJ1OdULmurt8oEF+gywnvvnqF0mNhLzLoXp2WYPbc3B6BrmCl
75ugNancLnQp4QvP3Gc3TjWYLDRgk4JHe1HIflsWf1EnMP5f/eIuL/hOOuTmxrTndeRaA33aMXBB
Nacggh6cHsr7FLwtJu+538b7Fdqfy+NnOvZ+QszX+fBAgDSaSS+3Dtl/GU/SixHpqKlvDS4sazVo
2NQy2gzcsQ3/1ax0fWpZlqw4eibD22I4WyBdsx9it/Okbb4Iip2mrzaU4JMPpLaZmAl6lE559CTW
YEv9ZgVuby4PkvFC+4GPTrTK2K4kdk5+mB9aHhmzBy85eFvKEnJ7XkpmoUtZf25zW0u7zc5sc1O6
mQrmGt9JReuYtxeMkO2mDbP0p40ODAi4tZuOFFJbio1nn8YMaFWvj/QE51AevXxZWPK0LmHXpT4c
0OjHzt/N1c3RWPIaAiZBpi/sfXWvRVnrSLpBWDWXs2qVMDR+zUJku+8WfwmY0dxvXgMrQmEmwV/J
kfIuVLc95STfKt0OpEpHEXTM6udCrAJgU52Kk7ZHqg163imOHwbFGhY2q0BJxWchbCYMQ7mTWFs5
1HanFI5GhyQ88Oc0C/5ihN0HEtuHzXvWdaC9LNLPTc3sHjcG00aCG6dLaiCh1hZ6+82/7ECwqnXK
mFYoIsHFLj+ekeDik7aR/lEHx6/kOXqwx/gOId3lD3hbrTlesQw/NMl7GlGousi+Mc2uo2j7sMoG
4MddHytkgW6e3tqnDLdtdEbfDR7FvsSIWGBSzBf0QE6lqOiWhaYdpuN/AmPLw3Kz1/491dFaHjzD
e6MK0cq0aYPkIV89fyzgy2b53N+4pA06k/4jLyI9kWm5vf9KtXvm5toegs7OwBY01JyCWzsIO2Hj
CwEDnpcy3uhLBN/54QI9sNiet9OYUIYnSfhEp/J+T6vgF/8DIlFqhPvbVqIxjmoBJ3kN+UA9gva2
Wv4/S3qQlNN2MlbW9mPjdTs2t/tui+I7npjIqKv79BTiClBxH4mmKlmNbNei85LlbqFIJTuOL6J2
G8Hc/EbgDS2U57c3s1Pte18lUW1ioGmBvJo0JilQVFIU8NUENXEcKffO82+hO6NPj+nb/QbCrbA2
Ltu37S9mlx0kTWY9myfq3xYvolZfkFI1aSrn3HOlnoZPO237ZuLgx88SOC20gCO2yOWlT7Stcfz4
zNWEMiJl+OnsM0KA3At4V/43d397ZLacZ5UuxdPbWy6b907BdJRy3/SJY4HHSkAne/gAHpM00C77
Yab0HI5bmEGO5iUhFDu0HynzWQcTWLeW6g9cWs4Fnm0nWK7OjPYVaDuhA0HcTpIhS5zP2LgHNTOz
7+QUweBw01/qzTUMQnrln118h0lQGs3HldfwscnIWXPoplWlIASdi/mhZDL5M3qHl025c11Uf3Zq
A1cO/ZvhGatmy/17zKQDIQoQhTkJfqqOShiiRADllTlA0frs3q7X0citdmveRJ0ntTS2MBPZjSjq
ueuFxQ7TBd3Tn1bOsA2ERoquBnsc9ZGd6VLoFmP7LD1oKWdcyasBBaMTEVSyxsvrKo09zFyk7pjf
zvp4PISJ7oFTiwdRaEUdhwnEqixUTBUL83Crq/JtFMKiqP5ftILlNYi0d1Q8hUcdV8JxhFKW7u3f
vNDN4thxtNQfhlGCHHOAHCKggKzuHJ4jZGAv4q8B+EO5yZMmvWH7jacWW4jGEja/JGl/13Tg7nkK
8b7dQX5P8l770+255m5HE5vwUzO+Ue8ZxJQg08A11wopJoEkOUm0WtB2C0vaY8DNj+kBLlebtCOh
qV3yS7ek+67+Vp4sTzCbor0pT6xjTlOTFmdfCxekO/wPFPWRTg3x6QbyMhVkL7+puzQWGa8jbNc8
8Hm2XlyPezzjoLIoXpR4ncUxhPQoRPsuF1sZaAJ3IYZdiqUhN8F63Wn3I3WjX0f4WyWQSN/AKJ0f
0sfAtTj7piOkRIC8O/7mPKeBCe//FYXFcDz91DqSXR7hm9O+/Tn3hDTllaZmhqAW04hA7MA3v7qy
L3gJxs+lJimTXK31VWvhPsqVwdGIR8Ied22wBndn8CztSgb4wo0lLczBLSi6WiReY0QeuSVPQhOx
RbHyyr8Of64x+mICrDjBUvMFefRVopWvSVUbssPkD3UBxKK3vFDZtalsPOYSmEISQM3u9dMGkoVb
d9zcoziFvEB8Q3PRa//gp9HGdOTn1F9g2XhP8eERMKZoLWOL5Pg8aicoXCES1xPjCTalO1djGTRe
uWENo4Kgpx9fOgaV9yl/XA+KA8UtsbuHBvD9wy0ueLMTW+3YNIiWjAZ74mM3Cdx53liY/SheN6ff
J8MkNEAYBRiQSkEZfMdeOZtFAbY3n6wUgal+FGhuGbuNZeA+/YBZbkjNFvFL54dDfcmvXEME60aR
56cza28HEfi1r2Jjqr7mqe8BfTNZD4ic0vIdfEkNp8Qfg0nDh78/PtgK96Wyqo/Qko99C6NtX+/t
cvZ5MnHjh7q2v2xr1bYtEsuT3+iL2y9tVHzNMDmBX+jZgE4FpVC6Aniu21NbqXtMdkV0OXWYTRd/
k4jotC4JPjzWjA7ecKW3rfq8b4Oj3Dz3qThYaz3hQ1z/IiQDvpXvT66oVuklT5Ls2x3G3ESbm4Mi
y2QEZsmTlGSJjGhj/D6yjiZpshZRwIS7EshtPK19s9IDyK6Q2cmPqzhgcXFuSTvCIODFx78uRHMv
/eYIdNJ+QqlM4snv/gJPBMU1ZMn02tEe8qPmMoWNqdK2jNUOYIMbwI4O4gxt5oJX3B41Zfj5yyPp
U+DFcO26qhWnVKqQaQaJTJkgoyYCCvFjxhKU/XLAq734xOn0NH261MRweAOB3gJiOzzy63WPTZx+
4Jk8VZ5CqWJd6z2HZWwAmkYqggfO63gaheEnHZOv7vr99qKggi4QKQoP8tjI3aXekmG65LziOJWp
ZbFtP1B7jWmw4uEKwfkFbgw5DZY8LBfv8MgQ+PMfY5Fbqmg37z1hpGoZnCLwCf+l3IE0BeXPKbbn
qGKf/gSOpK2UzDcRlzAspC9kKDTRtcaxUknthJ2LUv+nX8Yi4XbsWAys8TX4dNFoRYG6gK5TtIEp
prWJyH7qOAQiYi54C2xXX3e3YWSaH8umL5qVGqi50Dt8uhFsOYWVPrQfjoa3T9W2uiVLfzoJRgru
9G0iqawtu5xJncPCGmo/dLSs7wSJiht8T8EDjAFK1+5jZVxpfHtESvn/3FmXYH+5+xCPKiAHpIqV
Y2iEnCaYAfTvor3sD9D+8J+XGr58nmKVpLfMFRLvIWnWrkR+DkgDczYnh3pZwL1YOsya8UdOIeFS
jFDHR0E4hAtaVyp+R1B9cjsiXEMREkJ/EhgtLtaqQwbxHrlk9RZhXGrW6c9ya03nYd9DIE17I+xM
Y6/b0CXw/IuWubRaJz6Gyys2bCGDLEdkfAg8NM4500//WNr4EbbRLA2EbIDLuzvvunHOkQhdgjeR
GC4l65dQMBtj/FeKwCOr5iKFHeSPl+zQGvE0cdJxJl2DG1Ln4KzYT/CqXAHG5lrqMS/PI9ckhqOT
W5buDYRo6Yl6+q6w2iWGW7SsSSclmTOSdyHy0cPW0BMYMMIA2OvG+17zbXszYBN9PCUyierCJk+Q
kpIYPJWV0krhOHttxQBuv9MUS0K2EfRCP2MYH0rrGFDNgWs7bNpTiWowCzFfx/9WWDllvAGK/Ian
VUop3JwxcdSL5QMgLJakPXLh8OE+wi+cDjTwA1VkrQdSfHZUAc+gi3wo883SBSO3Tqggi3yxFjBK
ReFSLOtxf50q4iT5shSo/sJ8rARFJ5lUy52IBPDX/p1BasWfs5P9Y44shLOPSWwS0DvglNFJj8NE
Iq7WdbsilGY/LkG7JWey7+k4eIRqXNySD99c++GSE5w3Gb5l5+oNqokbjjtaBT82x9LsUDP4dlN5
Rm0Zm7VrBXy2zAjJW0GX35SeE1CJSC3v01xafafqCxQM/B3gMyC4B7lzKEYjl5FZGGJBFBq79i6P
qjYGsFLKb4MV1yLHuImdjGmapUIsuhExa0CaRvuXdjJ9tLOreCW9bP/aAGz+5k+NvTZHuc22YFG2
+KnpzR+UbuvJSixO5Ywyn+Kvdx0TtOJYULBDNpjDe7h8j5cgD9QCIBaMM5pM30v5FsSP+HCJj+fF
Ygephbji4KLWYXk/Xy/QS+ctKEuRZK892VMBfdzmJccqHRuozYM0Oxl9m4XXDzuyRQdmi4pJn//3
IoNkBYFWHmS0/vw3HIkccP7mWSyJDXWvYtfGqhdvY2IS1IYWuQbgPrt2nKeqFS+IyudrVuIfaPG5
o7+Q4GNvmEDnBis9YRb/VStizTaRFgD+Qr0QsJqgvlE9Sw+hvmnu6R6alU9vdth/FvWf3KvG3Vtw
dwrr55VF9SWMoAeEEtBLQtbypfw5O5RTWpfl62haKDJHzMtA30sL5j7C1mwzFmvvIxjjov7bN/cj
uXbXI3L55ajVdY0gKNs2a8lvRua1YVFPPiCRW0Nz4X3Tcl0KHkA46IW4whGyItXzBd1OirVrefBK
Ow19Y74YJC1WrAe5reW48k+V+qwAnw9bbUG/96ru/0aPrE17lckILsJzmbpcNNffMYPFgwk5RO9/
3eAuwZGRhDAltO4TIi9bcWXBgBLlv3NYD0mlviLIGVhjWciQ+W/GRJfg44c84Xj3doLT3OpMD9eh
9f6b7zYgp0cmlbe/M38uMWWP1LaAYZZ6Cz6aYug3PXdbh4xnnAtT5onRMXYwzd8xstwYqYBhsQww
Piu9vqupxIXDLSJzC3eOWVLY8KhnVPNUkSeKDYMigAgagCdM9GnqwXoB9632b69fx01GIElrt0au
oJ57TOPuu2Dx/aMMVsH+abvlRStPrSicaSfmaoqmDN67NVX2CAtkwQPhTzjJC/P5Xf306XPLy3zY
MkLbtyldlfZW126xZ4WGs+AGgDvQeZSJvm5CX2Mz6/3vv1sJ+5ecTHsSQv0epIYkilx0xkU0tuhA
23AeCspkNnGD5Cq0e/3P1X3e6/2U44hQ1XD++it8V8q0fC+Cyf6ZWhFilHUKzXkr5k08BnBpmVIb
ZqcwQx7nfk0Ir510lCanTxfQwQMRmxh2nU1pmXS7NBw/lad0AawgK12ZaoiecpKXukCr+Bv5HilX
VdWLbcLpbXjLRRv+3bdhEm9ll/dfdetUuqOdLVZaJ9CIa3793Ce6CM4umkY+toq9nSj/s83MetRc
PjJFnWJcp1eEBkSl7ORt41o483R7VDkuCNLAGa4q1XSzwR11Gi79t/Z6PxCYqZiATiVarTvvWc+y
20qQOsNZkd6ghxoFy9xtEo9q74vOjYXIa9thoSG6sP/8odNjLMqSzDS+FK7WfVQMLIlIoFy2Ftrt
46jQweRrw7RzXmhobgb69ogxqVYWQJldmMiI0nKpqNyTi8US+EtKIstXpZ0J4Z+RT5TLwRY5zPbK
EEFE+lf3ee17K8D+JvUFWACByFiSdz2uaulgYlLDDbMjrsbv/oZ5vD4ElAIk2ViSBfLswJrTuhAl
UUXOfUyM+8UaKOjlq6Ul1xdxqNroIvnK1Q3HiEOQRPtomM1+aI2of+xtqFI/egBTPRKgk43RmynG
7kMgt+7pAFOj0pWs0TsQ5y9GGzrKtJbQ6S47crQCMywFszZCdY46qek6CQPBS4OJWGoGKKirzW0T
vjONtIC3JMKyPieZWBQIvQY/Y2Z4FHMxN0Pdp9tCPPotyj+XSl/eqL37LKcBWAXOdxaLXWthBAEa
BnUr4cBbRXAr4QfU1thlwAJmaGiI4esHHOOAJpBCtWiVN+SjobhbLXaQH1vQMu530ioWXbw/TAxT
5DiVn2ctfh3RDOjbPaZmg2vwodSF8DVul74snVYYlIi9kNUdvoDDbXP7LVuXt6EFPf84j2iqcLeh
Pfzml0wDblaL8M/E6Stnnv0qnP3xUBL6RJBI4RM6GxaLj/RL4rL05KwJc+qFAvpi+B8yX/lteORJ
wEC0YU0WAXDuA0WGxGgIt3r5qrn4BDLyUu/tlj0R+46GLL3yoKDIfrNgF8kKAYPrpc8uDpyQjZuW
rF9he4d55Qi6FkPtA3HM6Z7GiL8b1P0uUvcoA2Tq2hbEM/IXymrB6dSmwo2hXSUkXOzwAKH6J0cg
V91fkLUz8RU3NjRtk/Gs6OuOnP9CMB/YCaERP9ABuywHBzy5iSeqaEMKSdEt/cEzO6GRRMkDGEyg
6rf1dTZL1Kw0i5P8LeFX0fNXoicNoEEtVhFU6KNuOcdpUS7BEn7xYrRDJaKIXtpRUJmsYmAfnOIS
gemyqQ7mQ4kbBRhmkvDdgC6Ak+AlK8lnt0Yezdt5bV2G/qHRdhVPSZglgljZnL1V+wDC+yLW5Ojr
yFgyfHDIlpxbu5X7Xj591zC0t5xxnS98CwR2fhr7mFgxK9IQbQXvTCfRqxMIW2J6emSTMgn5mrV1
0L0VFs0jWxnYQU3tox9P01R8OwAWLJXO6M7qfsCLWXdMqEt61zCxzxJtKPD6NDLasf/6mn51QzQs
pPOyvnl3nggQgw2mqzrfO1i9yx70dx4bfVXG1bkquEJ3qJe/plpRC3vC2990YmscINsBXigNnGrr
GDtV5pcWu4oAqea2QQ58KnMLTl/BBRXvzMXM8c7AsJlRKUO6gFPP2V86mKLVYqwcuX5fOjgqIOMG
Rw55QPGN2x1eLzuzMLodOxjfkqtQ886oWPaOa/AAdVBwAtsvMCZQ3/UIptJEg2X+mQtpqXXp2I2V
evkU1CurHOvRzhvmtTmaRcHeqHHUJN4eFjC8UZ653S7Ws5bf5Kf12dZqmNxnT3VehGCWA8h6Ce/9
HzNHuFkis/0VY+SFc0II4Di65pG4UDvxrrDDTgCc7aFmhQRBJu1lNNI4n7nSt5E8bE/MbB1+d7vk
9VmV6ED3GfrsnynIQj4XBnyt/uo9miBKrb5p7H2/5kuAjlYnGqvek6eHiL6LZfpbHw2TLXlyFYWo
chcCzo8o3PYkrziNY4eXDTyw0OzuXkThNTkXhrTrShn0Xe3OHCgLOWuaPEPoDIvdU2UCzqbPYun8
WsmzlwvkOZE/g6tusK2lpogSaX0Q/CHiK9fsawErm9FJNwI7zorfnOFjQCY41uIV5JjkXwdQ52z3
K2uS+vJ1XOMAnW2xao1hwufZbRgwZUbZyaNdCxpxX8BImU5Z3P6h4eABtK3Pib6O1oNLrnFSGX/B
ibnYVxXXyHuCu3Dav5kahKMnxJOQ6AwkqX4wNv2zm1m1rkpZ6CiCWEGFzwpVRFZoeMx8Thiv0rhj
eHCQFn6Y3uKgrH5j/B6gLPvu544Wnlsf+/1FiwK2AhcLJx2BPrr0Cd3z7J24ApsO4xvtsPHgbpEZ
4aPZ0qiDj3Of+9lmE1QSMvVFRszq4CdFD725MOEoIAG80gNtXRohaR6y4DgUxJVWk8+UuZGo2cSS
QLD2s02ls3ixgYAt++KuUrxKkcJHsH4+9BPF0F8NxLoECi0O7R3s2Rjl3CyxOBZeG/8Tvw3R86Wq
N/cR0k6T7Ojlx5AUrOi6lpCi179Wdvnel/DmS5OoyvqLZ8TrRVlub2qsL7+8zRyITUbhA28HH6gK
DRmTLW2Q5N78KnaUIm/kEZtconFDLohSFv07wMKAUVPkCIbQMvNtuGjVeFmgGz7Ca46l5WdjUT5n
fJavGdAiWg9IGlyeHeTy/7C8xW6gWQ1HVTZWtUOq3F5SFIUDQW4vZymkoRKTPaG0ZMthSA/CbCZ2
ttWckimIMo6Xd33btKay4pZD+yEYce1+VcdmgB++GoKdNaoLU7TQuLavYo/+f6d7M/3KxRiXxDnA
HdsEHHXJxHh/3g19/Wj1vZlSIlicOZt5YU9whr0j7dqPRuzyMm0zCID+bcdie9O4NzdboewBvSMN
KKy45oc/yoTIIXP3YG0bTcKZziNNraHWoCT3U+ViRrkde7n95lOZXOfjC5pVELN1IEBlQ5CRMFgI
vIAqIfNWpfkKn/uOoI+6ZiGs5H1MExIADnqJjVmAiF0OTe4n4zjU+t3VQ48qdXZZ2K1GMbWS90OC
2E6hqH2M1qnSVODfO2VFfDBEkGvaD1HBbBrTsFUZ0D6chsvrYMLeZ+qyJoOjHlj1XS9+VwBWeIQt
0kblj/AKeK270kSI4i4nfFE4YU3vUQXHdbKnUpDbOVysXV8u5nheQRDLU5w9NT6tjbzW8fZ3KUQt
8++FkdeOYb8pqHpe5Sn+zEzg7IHEpw/GegPVLgPYXWMU0Ii5JxwwUYjGihyvNwwl9tqDBte+0W2b
DdU/XtcCKMAPP+YYnqvXdopgA3bZ6/gQMJjd5xOB+8W/YZk+5NWrJRb3dwS9u8UX2z2EpZY4N8Tn
rkA0yZHuoGASNK+8+LbNo1gBXdP5JufHvA5eM2QW5mQREa7gT5jm+iANUT9E0nCXIo8Ys0ufHnWd
HiPLCBTYFLM9CQnKnuNez2x2Y8uSSorEzqQGX3GA2oSqrsa1GUKW0Nu9d/ceYZIu0dnEqRlD62hs
hkPyJxOVH2FlHvIevg3MRzHuPtOxL/zVyLmk4Dv/lVIaYa0Lyhe8exb3QRvYPtedbOk7369S50wS
+r8Vk6JRQZi5mgQ0lkP2XVADvqaHQizQ6sTdpDkQz+ZB2ysMwUjW5sdEgA0fcerUtFR978526qr9
NkjgI1EizM53zAA+5ycZMERIUBs5jF6+HpVjyO7zOCoNSEa3A5WZAUPM+xdUZcRsQEzFDrCJl9pD
TvzwgrXN8VBn3O/F8MLAyi2gFDAF41vpm7jw1l1wPemdWX7xd9N28pINpteKVP+gEhnXabzJnJGc
mN8T2ZhGfm2cWnfVYn79E69G1tAErn3BgW09UhKhjh8DwAkhrDImlyhhvEtcwWO3O5yLVd7QSCH1
afxmLxs7C/UH+5GyFjfP2CYGWTr6xL9UCpm+3O4ilWJoyB/Yjjy5YIq3I5S3/1d+Xq304UqJbAU6
n1MVo7GKnrW1+dgrc8/oG5za1npmvxCNpO3dR5wk17z59HboQMmoaAzyWUT7+y2Fzfrm54reKi6O
H5a0Ddyk/dFfCkCu5n2ngPCWutjvPtjb+UHEBGOYC8WAjnrBYfp5xSOjHNhMBogvSwXwN1WeCxLZ
t2fvXzROmTxnYJxkp/y3Paj740RfheopBQOlkq67GfyAsdC4ZbMarNpro03Vm9GW+PBzGByiXOgK
L4I0kqhwac6z3XLedo93WZMLlPyn5GCLz4l6A52F7Uj2ngZlISNhY8PfLIyQ8Bgu/zLWoPMfu4An
YMhBz0DYgPXAXIpM175JQX02Kk83vxzDs/Rw2xY8OXfpp2/kvtdXLrE3yUQLNj9zDB4QM2q4xnNv
vf++U9DjFFHiLc4muykRjiqNJmcky8k4si/WY8Z94zLyZu81KmMxOeEy+tOcxAASoKPHeKgNHomr
dUU3AquAHSMYVp7YhIlCmjZCLBJBmTcpc7G7NNa2Hk0E1Gsp8NWIHP1fr8t04yckK8cRey51zGfv
awhWXxov2Yiy0wWz10nfTeTmAYu7AVKe2gHKHgUIaw48Kp/WrVQCwV04Esw7kYkjD+belEaav+eJ
RFrJifkan4VtEBQHMci4sBVDeHj4vOBi7NcAOrFKdPQ/qsM8K/FhaDyXoWKWiHsuDNBRQojDY1Gi
GszbZNp5Un1npw00ME1C+mkiuwLy9ojAdnBrCCMHpLCSybSqNel8H8o2n68x2z4/wY0GtADJtC8n
R8Eeu2ZYq4L9s9LlQ+syfqmToZXGYPVNDRD+IPv8TsqgLqrSirHiPqrPSb1hfKRUL2jXPrgHnG+W
2wd5G6mSF0ThNgAZ5widre6wV78kIdrzkGpL5jGS3v8EjpOV20wiZUsvEKGhu4Q1ZTvHqxopk0Dd
P3hcHFqTm+1WbnA6GaBUn518JYlUIOhf98sRVcIuKeUzvg978iusApXz4oBLqccdKPzf36u43Y7/
9ntDYkmM6pDpxbRWWTyTdJO4i2R0T8+UPpdHg3jAQemw7oQz64vNETRblNnxfgq0QbtOpu67A7pl
rWbtVHUO66LRhkNXlgUobIczJfrMiyauMDMaTrnDS2MJ3UvCZA+DAt42uw+aotpKTEYEgauvL3xP
r3xqwWMfNN1S2pZizhivX5nmB/YGuvVOI+us9YKZctB0A5ZvEaEZFBqalaorl4OYbL5yMXljR9s3
gNtd8NZuMDIGrSu/M5URWsV1l7oRGIaz+bKWuFHsa26/vAWDotK7Hzz9ATgWxQtGiTCSWULVCX/T
oivcZ1gs0JhGq9FqF0w9QminJ6+oQgwH5nQtDiTelDfVFwJ+ucIsIu6XNdrvYvBdaVRiycU6REeB
WqHh7VpRjV9LYwNr1gJU/2FsAynFM/c2kGOU/eT8viVszv1LK5X1ctBwz2hmUy0TAVY+EPDv1Mff
5JxgWrrZitpqsms6eUlf+1jUGXjR1JOFneTP5FS1yjox3XhdwiJJV8hgkefnU1gRimau7umRgJRH
eaaI8ln6bYc9Hb1ExSwcSQa4eEZO+jOJDQZK2eC1nDofO22Vs/wYrFOtLbUx0pY/OXUzgQ/Scz4m
E8x9t3mqDkzcJL5gHKzHaCmKORHwsFTp7suQnY0rzq8P+zFLmZR+QF2K/AkPb+Z0QRvKcUXaA9kn
Wacc304AVg2kUR3YDGoA9ygpukuvHSz+eK9xP/yFjQ+wMwrY4vc1+l1U/msYRpVX/lyzltI+i68n
3pfWkEHRCDr4SBOfsiZWQQp9zFD7lKiq6SZCenQ/E7kkZ1yyIPWOPAc8K8Fk84FxJeBArEENMAeB
+Br2k2lx0wem5WerEWbKSUmTSxvJh7LZMDIqfLYfZOIrcJIpa/TqGxRF5SYCGDQgvo2ylZx32fdR
NulCVN+Szg3GszTI5E8i1Ea2M+WBHyxu8z99KsSVuBRswjHLUc+mP6Hrk4uL8PPz6fOQxpuBNo7k
x9VsYOz5hUWx0N/E2BjoqEv4bBEnJC9AiZNNlf8PfVTrRJPRvcO470SRqNRK8Tyfi//5nEYi3mNL
g+BYhGd61wKoJCwrGEoNpiXEoHZcWY7HBk1z/lj2lk6+hg1auqYP6Hs9XTbBjkLbZNN+fBfE9B7n
aBSVU1rL8ZTJ/O8n3FHSp6YmU/lEz2pRRPH35b+WibgSUOfcwi0Myuhaq6E4ZQs5DBqKvnMvegNt
GxOcmXWMxexo8tjb/TZJtgqOr6ZjHrQmFXVjHbY/zWbKrgNxknvS34zpwybgQvggXdqBEPxKUpgM
pGvyoidYDqmXix84pC9OEuNhjjCDbTr0bSFTZr/bRVcjXIcajh3Wdhwcgj0oXoGUkLru6qxUVg/l
lNuCR/cmDisr5JxqAtuIhnYqmbtdi+gL3MxS85qf9ZDmkwtwq1q1iyUQM6p3Vv6YHLBH3HXSodBe
GUxAgUGYLJrLsOlunvF/kDuF5Oj9ncPvl4chvE2yuvyDanG4M66EGg9jx/gfXgIKmek6yYCJN6pj
cwM+qkOYyoVnUnta9XbKfk7twvF9FskNoHeztJJE3+tS65yf6vqgrernetbblS3xe1Rf9rrh9f/S
e5jC2M7UvX15znvIquvoyUXy02xcNx8k3p0z9jDL3IRkE+9iNu7D0HXduD1qID1ySKAowyOZgmui
fJ9dAFv4xorJdg6FdNmcTCr2yu9HS/bulCzdqz7PpYDWpjMx5BgEB0AgJyebXYKo+6NrkyWEG+x0
kYLcQUdacPXIrTlwYJhYgCG7bUzFvuuKcU7yY47BqfabTpQoKIeWzzCMEJM+S9Hr0Oi4o16UfsOY
oulO5Qd8SoglNn52Ky0wWnb7oVgVOd0O+j+eRp08yX3YCseoT7YfRXyn5JrV0mSqbUs7w1M4YSBj
lKOo8yAzUUCce8o0/w0bmDPbjNqewzf/fS4R5hgeHdvRyY5IJelT4Ioz1H6RDP4HWMQX0eba7Vr+
DEMKvIb68oFDZjG/2Ihm/V24iK2sWHFnoJ7oNHbWm5ySLxzgIJJvl7s7cDnIKKXHWowpfaBbj6s8
Rsrq/SrLDoO1BbcRdb190grlFTpy7phD2nF+qpiiYX8W/NvxisOSw84ihXKs4VZVgZl5dDinEPSz
MzvRzAJDN/m2v+FMslc2lBU0yHCYEYGysbC+9Dun6IXbsDWO+3oUF6/RPkw1UjYeMKNc9xZFWtBP
cPjLnbRFCRz+1F/tHHpuo0L/CjBpyftSMaFXPPHNqDx3yYbsl507v/mGMV+8JK0kVgMoF45hkJy6
pcCvJE/jc1e9vfntuymIrWb45pKsq46XWeIZmCOdn267RwmRgAOGY3HEfa0UYT4f+eMdV+mv51XC
PQqlxQ7+t5wNPPQmUPUyrUFIoGiRoUwHfd1AMV+vV4tyv7+/OOqIEqz5rg9cmt3+b5ESbymu/FBY
ngf2U96q1o23JGK3YzlQB0BBAWTUNQD7Nap98arws+iEZDNWNpsP9HJLUENH5zvWpKpGgDUsr68Y
7D542sIBZ6AmIkltGQ/BoCl9t8ynU2LmbCL7zpsuXbCeYM/ZmJflRuj53u1e5gDUK8te87AVFv4z
g2cGAPdZZ6NQCpf22NXq55epcpfvsYJ23ELN+tb0cioSbGzbJQNBaMqXsoirhjBfPUzV3jeMRxZZ
WTorqXdalIjNaOz1jQnG2a5QL4EkhwWUL3Va6n00XXhaBWJBRWKpn57mjgZzbozwJYglO2XstfO+
ytNpkiV6zmtQucqMJ6zhAiXsuqUk32Npxj0QxZpz9w4HcHi01//zIiZrghqUhRgtG1puYYsH+AVq
pv1qjNma1vIr4vBkoBMEFUUvS8NBkLKF1xCc5Y2zFbEj+8QeXIf51ORdxBTaH17PaKIiRVqOQXEQ
EB+kX1e/3zgJJzeb+5kAiE3GFeprUa/J3PvprV/rMcQKw8o6JwGNDfaNKfIAi/x6C9/5p0GrvSpV
vN51AVHKhnHqfiSnqD4eKy9h9pwqpIsjOClQCqBBjiUoppaCP+Zct9HbsT2G+WMDxz1iYjkSirEB
uzKg+lmcg2V9zcY6/y3Z/ZYdTG5BrRT8GQeuY/KjX9epaCvRsi1gtZiZiiYenJUDsdoTJtl0RNBm
/hhRyQfHQyOWyzCTAI2QATsvWU7TFD7mRCQT+VaDlLiu5Pq3i0UPejSMzOvXh5WYwDFvhS5b0f01
OqFJ+tYFxfDzoVuW7zGH68MJnIFk8vkZ9xPKQFlipGhoFkW4RWQg4205uyWRRDQGYhlmmX5YtGvF
o5ZNvmW6R8ggQ5tIgK52Qj/sh8VoBZ4PrCoAMRJvhLVacJLplWlEMCcg+pG4aw6l9hW+wU7GpLEg
oIPQuSlsjNhbq30c9JAzAMYpNSvsR8P3Y4BMcepHEodB2Tr0W/WCtHhnNc2OAyJ6OVFweobM2H9y
XlIhSDYP7bxp4qzyb8J6PsAjf8JZmvWWyJZfboEh7ArkOdqlL7uMGJW0k+dgOUfujsVNDWvClJoT
Qj7btXVI+slJy55ajg9TFJyjMMS/wJKVsM+bxS76hCF24kjjxROBVdx2QxA3rZXBAxEyGzVuYYjH
aPRYmuGybDbVUgR0xcBW2beXHYWvikY0h09BwxlHe3PYE+s1RZKJTRLrotDWcOnXgbWq356O/tfS
1u7fSSt/IqOYFfoQNLBYBMz9pc+Iv57rnuSfJx1EgbmkEQGxDIB/cSpLMi6IXGWZPn4hR/fpjSqu
B7Pl7C+NbIRL+Ia0aGgUKzDuCpZzyZ+pesXncBd8KI0U3Tne1M2tvX1VAIAZErdYxn5/bqm3ax+k
0h0y5OB5gOfevb2JtqNrx+4dXcHiETXPp2FKfaZdvSusJMCWAkJS2dJoUPWtrvk1bo93Oi9Ixx8Q
1+an52IznkXtTyjybohLw7lUCaq+/HnVPTNrZPvL0YLywa8hhCnfvuKZiVSVQ4E6UdE5n6lMOoEa
E+jhbY9bpm2TXGKKR41VHtCqL50GVmdtRerCbzTkVNHEfVtUI4IlPos0QsveMY7wmeUg/5rotuaZ
mJUjRb72rAKfAoicGyaGDAkJNY8lRtmQ/3YyeMaxYK+kH/i6ePBWXBIurUsOHTiFwXR/NwKsZSdp
IvQj3nq9a9wj3kYstMN729NLOozo9keRf7fVmWky4xuF8cFuiquj95RUhcb8MRVh1ntYGdNdHN/m
1e2Gltsb+wXL1yRwrDqlJmTgBWSKS1ggUlKPTK1EZMte6iESf/0xF5Ha/IQalGBN2PO+tbgjl0U6
EIotJ2swujTeGxauRQnx5iAbEITPVc/ntcfa+keyWxsRpuIknVqpPcuyVOVDXxePxHzgOF62MpGW
vst8oEIUFe2VSjxb6VByQlfo3sejnJ1v7cevdexrYmcFNTOF1qFnSsOpqm42m6/zmHl8TrlgH5s6
2CJ70PH13pCK3EdsJN5I4SjvE1/Ds/EvLS7jxgIlVy0GYV/ESdhBvkRLeoYDIroi/TZtoqywqAxl
wz47Opvfg19cavU7nuXQO/gzh2wX4hqt6gLt45TDqdXQRR2YYpzPp1hm8vV29iQoXsUSXLUFNrt4
5CeVJPGCFuvTEy1YJyLhLA3/b6urokLmfKfMNn7JbvkFyFvYEDP8gEAexHUm87gSGqyfJT2ZQPp/
cSjlC2c53Nq25oXZYoTrB482Uvj6ghbojrXhXQBXBObiedZVWzR7yK9rw2WmO6OkiiYnvyXeUhMg
TIanjgj4+WfkSJ4UleNDQ3r1dY0IFdiY2rE9BtVXlJzmcxGNDL0hGmy88fZcBsJG6WO4sr6N41dG
FLBDylq8wdrxeCsOl0eEeuTFZIhglQa4UokDHYD5P2fEiNl2mfBQGGRvYtuVlDlFxiD9wmYcnT/l
HNvb2iUm7bWUI1rBDXLOBgaz0fqxR/mBts7NcpCflhj3v0MSpyApSgoGhdcJHB60il7hi4bGm62r
qSNyy4zEZRgIemaG4BIFUMAWZbyA4fb1EHRLKDIDxrJXO+SNmeZ8OGr7Mnh4K+e/gRAaUSt4EopO
gDRlCUNe4QhAKBWCdXDWSiQaeI0Hxrhkqhmjx8kQ/Y8wtBQTy0UvpQfdfJR3zC8Z1KOas14NOs5g
86k3dL8rpE0A8NbbAKXYjiIxSiEcepz6HRoetaz2Y4fu/ZB1gOY51JycnRu5FSCJqpBV0RiOaI14
xfJFznu//2ReUCPZ+O5Fnb2EcPycHY8MmzTY86E/+oO9gHBjJb7FzHC6DwjgYopUwGmZv5LCLhLp
lDStE2qTNb8ffl2AU+NXg4LqEKwfpVRhglBEH3+ttVo8ZOBdF0tIbh8s7wHAnXr3rOtHiilKHmbs
j9vKuqMbxu1BxACf/fZZVKl00FOR+r0+FLPGni/ZjhxZjMeKzGecg0ZyGuYKzQ9StKFjgUYSSl0u
wr5UVTh1hHEG5/g3C/8leo9NOzhZNtgV4WvSdM5xxFBNEn6v3/FiR34MbYF+2H3MHSgK9BCB/xv4
TudmPbLqnyz96SbWeGTaERpEst7B8QTkOS5sCVres4I5U1zubyiqOirzIhcDHjmk77xzyPJVDzDS
Az0dDKhleY35Ji0cby4lEOmTAao70yait2xm6F5yfGqcPWUp8mDY3hsljyY0HgPyJZ/ZQeCSkcWt
xt7UkzGGqng5twVbqOu91VWDWEkBNGR0Z8VfHV1P8MJDBPMnzc7HjMqDuJ7JRQ0RHDEVf202BZOi
LrSFg2bg/h0GHn2RK+B7Dmzuu89PZbp4UNciwMRfRDIGKr8KKDIF5uKAm0JNiRU0mSAc0It8dOa7
2EjkCME+sWov5RaunD/xLpOJTj7iWYPw/vWimSLk4dsIV8v9ihkj8dN+Hu5MrV43GCBLS1kyolau
eZfsJsx20GrIsjary2OSQEsZSg0596pbXiB6leXek7yukPI4faQnrfxlTTtvPi61TmrjtEcflV1m
+vrpRgJBLfuHkwiCpZeDAyezJ14zG3+7PlmsEwXBMlOv9QJlcAbu9BsdrTtvUeCfM7s1vuKwIPNz
m5JZyXTcAk/rHdqxQKmWg4EXj+O7Z5KP1X9wWbEMrh90+L2YzL8gD8ShfLv3nR13z6sTSEABiEe7
Of8ZdyZRKtGWj3uIEragPUrfo4nuhFxiRp5+wlG7gaKEp03sVXRzrjdeUlZ7NeiTXti1hfo5J9xV
su99KP2o0REpFyMudtTq3aFNKf0so86g2T1w+2bnAqP+2ZpGW/wLwXh1+f4jzy18QBcHYnKl4sfP
8g5bPV1Zw/kS/Low8Ys2lZ2eUDHWEWsF1ZFObb2TRjEnLOLTN3yEBRMs3Koyzr0gD4ceCTtLTG3v
A/ioxP7qFEI1IUZaLZKEwnzyHyvY5FRAxUKKkERRyrBeLkon20P18lmqpIeWrpD+d/4e7PSF6sfQ
IN9ld0bapxu6jzSV7TwijICpdmxkcoDrqo48OYwTHfz/GvkKUdRK8JSSK+NJVhwlRRG02/WnMnXB
/lg6ugKgbmwcjrSQJgphpBeZcZzRvSeieCd+3tBjMer4GFfsVcfKM6Lb53RIXSdkP7RHyuIHlppY
IrCRzhmFwdozUiyIguyoaTxhz05RymcKnPF2rZoOts1HMbE0O1vbUAhZOsMktU0+W4czLq1Wg9fD
H6FPoT3ESDmhx8w27dROosgLUhQDlavTE4P08j8HHjI03jcy5ppW5F77KTReSpiu8itVQHGplsaI
4a3evz6oD8EU3m9+K26an6yJpcxa5fEkNXTOwfesfYyzvXf4MYPDhPFi/3JM/diPt0HA0n+5ZkIO
lNbnMpGfDuwDUplVQfVHrbPuzAwe58JG5QI5wMsdo82Lc3nQWdYyLNGlS3uQCfvdHuG9qmZNPmHf
rouO2YtGcXL+5prm+hKS8cLWTKvpwFz+CvxLzHBMgeGWIGGdB6CouimYzITlJsL6eZp7ZQo4oWis
p3wz2ApcqwL2i8LDaCHnkDJ1JTQ+wR5b30pqTI4WbRMFRYyc1HWnhtx2Xzi7xyKpmmDudisiHVrE
pc1zTxfONS3GzO2GN/fS9c0l3Ka1fkFzeM8HxsEkNfn6HnjXMAy36MBz7beeYKV1AYKDLl2v3nQz
HsD7GF7ZJ+I4/km0pdB61xOzD96VylacMlxZgrDqHFyWs4uOi/5aJA79ZbwKMU5fiPMRCAabROQ4
swiVxX1Fvd6XeAJPakS6RS++xysxE8pWZ92w3MT+etP0StWMWkOnghkZtLGAKwPPaQdKLfQqxc3d
7lfjg7ISF6ZN+nDCjYgiXm4Whw8Oq3kDlfxjaO7vi2G4RVR3B+VGzUyCan6PN6b+pw/klnhgPGRR
XT+9eFNwngsZzTiXD1DIisyVVAMKzx/YHsJ1RQYZwXJqb9omo+yVJjB7QIt7fnMcQGA/2UN3DnOK
NKJtFPi9i/yB08T6Dn7Ts1D5D1jIhokeNzH9HM8FehhpdY732msdIOYW6kptFjTW6veSDeV7CRgb
YDbwnvI5+JCwpi1rY/YifykB+vNVa/pZ015Ox8YCyFIGvaTgPOvi//CJzAXWPcd60aKlus0ForFx
SzbxF1Ea9IWWNO3O0VSutCEVbjH/9lT/b/iCq2J+q/2iJ3cpzEp1A40nJoK9vs9rbUTDC+P7Z1VC
JnTLgZazYZEpnGLU54tq2wzYqHSSsN3vx474xnN37qSw04eZhPxzTfXW33iIYyNYlznm2+BHtt+X
YQjmHXEtKcaU379bx/eyWPZtOHEQsf8h/xrJ8qPw4Q0L5y75z3EB/6fhjbKYjztLMROCeBqKJO4I
RwCMi1alRr1rChVdNACHtyl+gQQFqrCWaTCYtPZwsOdOyTbAoLaFdA6y+AW1YgWZE8QDk7P+MX+1
GJo8f0NcOjRiMWg8cM4u9UfQcM5QAsZZJMKwYJ8VhVIsl+z++TAbRsRPSchqFZ8TJObcxqzsXWPj
h0RsMz6nefFHn6Mfmg+3uvfXyc9sLf5E2QBjZwghcJU8wm4TmqhRZtmRr937fz/+MfeumISBwpX2
plC6070oQyKjaO02z6DLbakT1WUVkvDsa1YwD2eBaFIj33NXEqCHvrJuI0T+RN6NGR9fYTBY+XVF
s0Bb7tfpct7m2f3jVsIFCkJX5JIQv0OEzKEdTonDcalD4hTE3fV4w/ey9th1ng8kkFo9EPskAIDa
OZellU9nZyFkXG5Zu9GGhgo+9PuaLZMwEj+dZxsyzb7+f63Pqf5CHOjqw48l/K8aIvDecEDRT2HS
/HWqhWVnra8GkbrFl0QCL8gjkeEIE9eQ/eNc+rCZujBno8xy78wkHZIAcCJMWwWfA8rSNNmVWiv/
89eWWnDNj8Kpco+rYRbYDgujwBEmUBYJACs5bD1Hbg/sRbUTdFMYTTWUCvvHve81ERbdnsaxI0Gg
aaDfMkzpmnJedGcQVRNknSyws3BQTwFo9baKSed+shdtV8kUFA64SB3dACJ4rV66XEV5fkXbw71M
5cpDiyDUIv7OZd4j0mEn0PSj/bN6v2nL9dgESYV2qVV57q8coyyERKSJsNuFrOVuPxOsO476/gdP
Sv7HEU8StChkK1PWfCoe3dqHM+t6El9dW7v10JdrmqkbAd7Lk9Ic4eJw2c6M8PKbkIleMi2kgAPO
CRdPgWy1omecFWoYT4JDJsBhrOU+S+yC545igDRaMk+kcgYr7bLiQDMHSsIj4PDtSptHmN0oMRjl
eKd/EwchwX57TWLxpj435Af5LpqhjjLDlOlTLdm50UKfx2ztJMp4eC/ZkRlkxjflH/UjNx4b4452
RIg+PcEz7JdBYkORMjTEoX8MJ8qeGGXs37qPVH9UvzSJCH4ZtwkkQYoHhJp1cSplbqcJC+4GJ26w
rV3bnILssALjt5++RKIF93dwfPxdsNeugRDGgXOGO+ewQRc1yApKyGKgEsvUZvmcNe6458YxziUu
sVRF4eWpjTvadvczaYrv9aty4oz7NReuaez21YQ6vI2iCvyozlDjJX5hZTB9w2cz+wLEta5AOB78
Awi7V73DW3qVd6PvEopWCsQFGlNtMOXWrKx+TxbeK26j+oV91sTyigphPV+pV+xyZ/uBHSZXnJFL
/YS8xgKLXyAbdD13lrSwL/s+nyJCBUt2P+JNrktTHf9BrryiuAxIjGvJXiEhZdWLVfqoQspgpBlp
4vsnsn2kQy24/C58FbXqkon+H2IECFn+eXKsfuE5dN8RpQFz+9DF010Xn1ejv1fLrWV35Xgl1J1N
JS/rjhcjfvjjN32ROeAfQdKq+oocK7xHx1WTL/yXE53amfG90HnidkU1NqpMNXH1vMMr2zsV6eDT
voWuuqK9HlmfNiHJOCLesPOkEnM8O82/hS+RyYTyjc1rGvkq9SVsaLN3q5VGQ8yBaKKoOR5Rehml
0x6qEMsSzqJ3S0YOtCjjVyYao3RuQfN7sqy3pyW3WiDqBtgc5cWXdft/z2ySWEA0MZyxeRpa/bJr
RWQdBi1vQmrWHpbTboOIO/S9XZT1uQVglI/HJfA3YselwBpfxVKpZ0uJDVK/vh0RqhvBrIEMoqFh
XTUP/RDd42wUSK9GDFyGYTKogMtGkPwxQj1J0RKipr94UqZ4Kd/6fuYaa5YXkjrKe/+JWqgaaguP
aZuZhbwIsN9RuNovBWKFPrtAbkw+tNzQZnSg8ZbRr4EMTOACufI73yQgvLkx6CKsGuiykUvYroh5
XO2kZcDfPsjGKZMbbRkALd75iUYoIMApZincryJbooTMYv73TF3ozMibpYpN9KII+Scc431z3fFY
w/8P4QoL9Ej7zee8qCt0nuVNtfmAqqF2Swpq6TLDQGcJYjiAFXkWZHv4fGOWAKWxcAYLdUnFaWWV
a9s8uZwWJ7PR1MXVPODPkswMWhyIjVrMG06XeOeDGchOfcTKH+l+QTVW7+KQKVCC3h1nJcn815ox
ZQzT5PzdyR61NF90r+VJa3IhCZhBh9Yep++hz0xTjkdS6nuAL03sijANAELZ5+v63nCSCqKYtm3D
ULFLs+UXNW/u7UKRPguab6NDPbYgwOFHWuC9232yeAvb4zBUYR2yD67aIW7IVv3+CEdSR2RgkRhh
K23zHFJqk0lEiwWNoKomkDncZik6u4bYezB1nINdF2eaPAUe2MAAii1xRkeC2G8FWHEhE+Bi8/oN
uWHAN2UQ3wjDFJz76IFBw9KeEEiC+STocEqqCQNpGgYTw0AthPtK2UttNWgTuatdHXioalodhck3
ja1iR81WhBt6plGd1ArljOy3y5HlqDLN2A4G8mMCgjEcmGoBP/vnBHJWRDfFUCDIFYb8u+76+iIg
L6BMQHsiWCvOfmGeKY8HshNxhbKn0LoCpzLuizP04tMOXpNdDPC7Wyo3NCC7Pz96ce3hIWzzoOl+
A7TdCtKsyXd04hjzDwM8fjhZWZ6ZkQEKWPyRQpgXH/wf8XqFSX6+AneSFIuTvTPc6fSB0Qyq4AI/
Xi7mHRIitc9uCaQKmDlC/HwggX9F2SJttbFAju6nIAlhwBftFzU2fc77HeethFYEHXX+e3B0cEZg
lu2LITNBjRY6+eAB5SmCC6XkqUlmHCCIsHQxOm0egrMxulLP5Oty6atFIv7/0jz13nq5hLXcUnZ5
/NhMrfdLXeOqx9827tpINSbfFezFPZzttf9wphsTgx9w6MV3JJwhUzt/6H/I2a0ati/vK8PVrkNu
mpz7msh6ZJinv9Q0KHReC1OuHxsV2SzHNZgTncZ7i48cXzt6IxTdja7kO0KyUYv3c4e4z3LCrOyf
JBf9tJl5mycP5WOW8KtY+LdGayjaBmDtTungbhSWhFuTAk2n50q1Kl369dZXN5ljOVXpPsdfRuYi
pv+cVp9KxVQe8MGNwaPZ2CkD5J3yNHaSZkDmEocitwR2EwiViW+KD1Yj0dB9KSQGxRek708VrUoJ
DXI7M6abPc/ajWMbX1n2aAY4iWHv/fJbr6phnF2y9bW2e/t32tsPfSkfPL2TB0JOv6haJhxua+hd
izfRP5d669OBRFtz8sM8DCE5D84+gIn9+qFGlo/waWgCRlR/iegCCO75krYCG6A2WxfbFTQrw5od
A+t1HJ9Jptx4Ve4ShDmkyb/kK6RhXzTSTntm1nD88SH0DzBXF5aFyUBRO6ta/CtSWPqnGv6c46G1
f0eW9rsGNXnXBFIuCHiYr0qSFL2yM1rkhKQO1uZZ5TVjGkU6bUsbAhKS3lQLXw1Bq3/vwngEycO+
rDuTLAwwy7NVFQvJqPMT+yJGvVFzVIpRN+T0OXUgt3EeYkMNYTIeZCil0oJyHkwU2Zm8ulyDTQ91
xW6MPmH9psyugR3xUWe8ZKvUhZVKF/9pnFamlv5mxjfeqC5Myn3g10X4OFUpAkClpryuQ1IksC+l
3ZyT23eGeLgFWC4ff/S9GoBHiFDLeH147RJiyLu90w3rc0GGMDTRTlYTpFqS6vIY74ltBnFRD6DL
YQGyOfLFRSw0hKK1jFSEgg7RzK83poh3snKqg31Zeu1jy8R/wfaGL4kLBo6u8WN1Zx1s3pgMn1Jn
LK6RevyFM+IPRW+xJYQXFn1dcLv6ffH/DYT/SeouzQyEeoagjVWM5rCjh2VHbWruPggAR4ilMdCM
Qq7v28vTRLyAk9oDsmglzpxvK1NKkV9mtmCod9jmHthK6y4AeY++fvjjWguk+mB4lzP9IhkEW5nv
0VNE9LVVz487QX+YvcJEbsP2EnOlfqP0J1gL+JM5cLYJVYIBXX5H2ExXYIsxrgCVCefH7MiyUYnr
IPDkC6/C2N29Ar+JMqz1JAj3m1y8n/XPtg9H1w0Ligs+8r+6RomqwX1r8W0ym4/w/JdTDYqfltKJ
tNsR9JVniCD7Opvm6HIL9uaeuZyxLEd+PbetCjGe9S/P7icKhnllOOGBorIjxp924A75Q0GhOhIA
iNrVc6A22N2JpZdcQsmJ/uyDyUHFi4yhf+ZiPFlSBnWEWjFcTdLHz+5e59cTk269i0EO1FnaxkFK
EbBChUslLbpYbM8NmYhme0ToICAGk2HFb5Rhx0d0AbI/c8NqxXbaQeA32S0X7eqN1XrB8rxquNpA
4Fe+q8txS648XRjP7W63YLaSaBIBnwshpxevD9nI6y53tuhweixwcw9nDq/qbfZ1kpWUT0aGLrTd
AbKy15VegiEQUvfScaRttBKYCGtj+/2i6mMwMw0fEG/inUgb1o+mdBEve3mTSnLWwWwq8JLzBbJM
ckGvX6szzXOuhyTyTzZDJnRmzPep0B1SEPyGSo0awI8X8NiNf5Cy1dcM6cZK3kyTlUBOxvn4UTLF
FnnU0S/y4Xcu8U0s1g/4+R/vib4je4Mupb7tXPk+z/D5/MCIpLWVm6L5Sncw5j2xjSpH0nJpcY/5
PxBF7KazmMw2xZdqf/4LARdgfssgxQ99O2YU6vjWXzjGQvM8JPssVQ10TbZRnBcsGfRzn9VaBwjc
o7ixvK+f4qj0FAB+vd+gPb3NipWgJaC4Us1jyjVir0O/9hkBUqFRWH2y6yymLMCZNFWij1thoJPK
lsNeY9OPZ+4cKG2bmurbpTbfGBaAhnhuiFPgzFG1S+xjlQ+ocL7oaZoPlz72s8xzptah5Cv1jxSX
pT6Ok4qdktAiFdwEOglxp1yo28yKfI2JKuUA+6yk74JS75Vmm+5ZsbFPHSiIewOxGulYVbMVLEdf
oVJlKmkF3XGJ48QKdL6X/SH/0WFe7iubvl+FVSYU+xu5IF8M3O7lFo4N0G3fkkVum6fc/I08E35c
zRHDtlvQoQ126WSvkelYWFisop/YhR6IOd/3bOYIT5y0ww3xCE8tMPSv+YCOv5hOVMFcBYtS6StN
21jOCVrwzIAZMMR1gasNlSgMn9fe15ZirsGPTZQ+5k7Z6SHKdqfVgbaM9zKveMJDHb+g9BY2H+SP
PSpSlsSCEJI4bM1YFRokPbE3HK/zt9XmJTdEy2lhd919WotZXGf+YeLYNO/N+o7kxqSPR+DpbLtx
gxfEp3CLjjgJW9xmCSsw7iXqZmGNBP2Ya3paKdgiSCZNkw6paob5w8J7p04Rgwvyz37ddn4jcXSZ
Nf7595DFjQWnoYYAfg90LY24Mnj41uQz8p1xGq7MiZPbUxiwzEsUcjTpPeJ45nXUe0HfkxDGh3vV
46fjOqZzQAtfcCxxwOijjuh77KkqxtNhB+m5qPKQI5jX7WvLfrSf84jaM7tfVA6nTXUS04bodSSw
AUr5LP6LvwmQCfnidpLb0YOFk4UnKKqi3xarhl5IgNwchErBaaVqeaCXrAqZMFH0XBJVR93BWc6u
wokSlcfS2CLQ2oJfFHCRH8dJZOEdNW4sA3ud5gIj3/HP+LU7iPOjxYr3Gw99vA9/kqFru+USpa/t
O2lrOb0Nl7UpiH4D2QufgzwQsxagWpPNvQKaq+TaBq4gRy9IEYnVu3wKJ6U0i57o+jSuAKqh5DER
ftNC1lyIVKQpbnIGkDe7MCOM1jSWVTgHw+G0GUV0fyw+UknoVxNUdniUtMwwsszNNAataW5Q8409
hEB4LsqSqYv0ZdJsqIm3bBiloI3S1ezuelyS4nKAYOIZhghvLkqP09RUFnQ2ISTybCrKLilSfkdf
n98nfszb9MfVyXfDVJExcsvLk7PDS2IFk2NJoMxmbHwSWF/F1HThaL/dZ6fpYv/LprLj5FfTQsXL
zB4sgPfV6RnuZEhPLP3prG++t4ckImR/ZBCXNUmRHTIr/rEi9cDhbxUhP6vKB3wF2GMO2X9boMZa
j/82E9fnXObgV3k5pK+cv69qqCiiLotp2X4gshapf5Q+YHhLV7Orb/8o36VeqW/Sejg4rwmYykle
Ot+S8aXZG5MgedKxxMWDHr/gl96MYljRWSUoScKukI9BC68vKzE4K4GFuqoPw3+WGXLssRjsTjkS
MBfQHbRxuutyvoRFinFMAKRGrt5f4XHOexi/e9YYugRBCSA47FIBLWBeyhlXcupNZWUbDpWmh0ZJ
PzJuRG6bKsawU8bNyQhCWWewRAMZIS8d/iwkeEifEzm1MlTsAQiZbACZvT3O99KvHXxFg3moeoDL
nbhTEiEE6sjrSzfllRi0kxONta/kSFH8IR64UcI2qJsjK56eRDEX2Cme/bgtIBsKPGtYD5kz3DS9
M0InSQ2Qh6jCmXAE5RVQ8iwi3SnM55cm0T7gugfmX2zoF0js5lqdIxgt+nujIMlig9CK37zZETDD
n6tDfc+HFDeswyyIFPv0z3Td5LLlx65gB2cpFtEDnDAlFyXuo2srIw86vZv+VxKJOFlKjnlSKa9o
9NQxoLGahO7PzVohug4Tk9FtH98caKP+A5tNeEU2jjDplB4rYRKFOy6oj+2qqVNxm5/S70YRN7gD
t4OpekBola9ysLfc3yEMEAzBhjHFjnQJ0KMgo33wKhGnZRuyRBmp+YrBYxPUXrFgO4gz8q7Ja71/
bnDIwhL3E+6IERWRrp5H00GN4UeIqJ3NnnJwMLL/O4/0piX998FGJ3etswlFt75fY6qY0CbgPtoE
RJd6lJ0bGfTNhR0Y8R9lFut78d0f7dDGCL7F0rHZ5UoryG8bRzlZOtHLiIC6OrVvu4uCuOwideFC
4bzMoYtyJAS8KkJdQbOv/5ssyGmlGDh59YwCcEQdurKg/qFxuUcgkiALg9HYuNG6WEnlnvbtQiri
NIe6pLClljBuOM2dUj3nLIgrHmZqqudA4D1P3UJympjuAGZIOsRWmftqT0wezXONSjtDGqqPP3fp
dsFUC+ECZXx+7MZCL2qmD9VqiRfb50xsbyU7rKV8Vds1ALEz1C9fcuAPEDWA/8a7TQgVsv8nviqG
5iO1FT+VMWLnNf1Tgezoe/r3Adlo9nJeERqYHW6WuhbdAD3n9l7F4hrmYPMEGWSeJxlDzWxB1kdj
MMB0si4J1VxGyWV51gCvojfMaCRWXMP376Z2QcwVvxhyjg9QcpN5QX0+fxQvSE9eiggVkbOEuRCP
ciJimu7xOG3bgq2t1pJK48PG45aLJiHMaL7cbolOFW4SgzrbHSSikx/0NZq0UD43Hpj22/9mXR4H
VAbEM+4c35bnEId+sN/O9wojFx9hpFyRwFYQZkcrK3wcdQKZvufxQrZDOiVrFoe777nHNM72XbLt
N/NH477bd3RAmd3qw+rMXeOXiJQji92R6Zbyz/vkfZeCz49WnsT64zaF2mgBgeBnqwCaznMlyR0u
dlzknRwg68K96ny3Dx6J8iwBeVhVOEHx90+iLMf1Pn6xn3G8WET3dfa10wy4SVQ+D+XDJ6wlBM7V
7GQJpCahFL5lZqM2+4kpG1TvgUY/RtyYSgj0XE7SBzMgZsYwacTHDfsK29T0lWDWwhG2mkt86IGs
EVEDI/nl06N7mZ0cjpk6GQuX7ByPTvcgGk7b8i7lNOvz0RkGwdAuFKjQ4ZWlP3sVo9Z9efBRWQRf
p1Few37X4Ltaunktq3N2eVbdv4yaxRdE1mWheKQRfXmMVhzrb7sRzzXsS46RQAk5sP8mvDTIN+en
khlbV4LTLJpBhuFBDrTZ9Sk3QXCjaNT9mmeUP7ostlLXzjYdsjGcI4DZUvgM1FkDVMsTpEQwTRno
Rwi112PhC0DcUgjuuVcVU+2xGjbGL7cYbC2g2yAcjvea6iXhXhSO3hitLZWa6zYsUuFglVvheXba
e/92wum7MrB6Y8PjI6cUYdTsgWvnwcb5Zkj/EqpNpLLk0/mUP3hSJZoes2onx4fhw6DCgL381X4b
4Nar6fuLDpePF/7manaW8ApJabdTFw9PdARRYWTii2BfxlbdnoSJ4B8INNC8Rc85Ou3cnGomSSuY
r5d24QQhZMO2ZZ4sLb03DT15DNBsMZpqwFj/awcBdw7HhWqQU1zZVIwTEUp/9x6bPIGWEYGumBaB
zKZkA8sfniX6neo10U0PQp90QMrwrEwDSql1YO/JRFaKfQY622PnHWDe2T9iDTShn0ZkD40/vHZD
de+ChUJL9mQawxfi03wDUTScBoTXTMO9ZEM5RiPM6HS4j3LnOrsZ/v97IYnwMPv2UWF1hbDOuFCd
tvlmkwuvRJ2lZASfUAdnfKs5PdHq6kb6HyXZ6wldv1McFR8YLGe3S3GszOCxdaqz/XmEAjSkkTqA
bNwej2920QHkfylkKdNh9maQEZVHgOt/xWPz+xXOLNJhL+z5DxqvmgIdes/Y2uqpVITUmXeNr092
dfuZud7TCANLQbGMb1WceiiScjdscynRZgcs2j1Jn1mQm/XqtONtuevmnzD6jJC4E+75ej19YEnw
ea9s/bzQ14O8UY0ZIzBSrRa7a7PH/fmy4gUT9+HhfdX6MXGkAJxQ65CA4PglplQjF790Ur3bbIvV
AO8CH0nCFZwzXLRPz/x5oukf1Zhn0GPnTqLajk2SKxau1WsvPnr2S2JwnAu5GOzjgftmE6KxW4sN
Au1cLI/JG5hZ7h5eFuZV6UCOU71rbUnkR7JHXArjtr5/ac2PW+pZ+I8qvJ09JV48/Kw+MZcBPz94
V/u5O42nQghZjOoTm8oCCMEa41w6jsevK4jm3D9NxhSofQUGNG3jYYDVO7rVwzt7bvzNyjI33azp
BSSAXqOpvgio8uUQ0Fz5sM0nsO/C/R8vivSZIFBnDzdVkRE2R8r95P8+zP3nmpDwErE7N2jjkQVt
QzobSGMJtNtEBjjZe2RX1V6nfyVWUT6MF4vjRHcIFU2rdfJRZW12x/46gT2d2E+GzyCax6ATNSn1
vGHa+PHeOkFRwE+H7NvoNafWgCAMfSUnhRoy7Hu10DCl+GOCVtiXhWI/SKML4v7U8Iqzgv+WUl6h
6NPBb859d/LYkmmRPWcFXeqjaMGsewmXmWwvzYvWnhhxT3EWQuu+K427KcRW+BBRHLOt70W0PoXh
6IIzwWJlxFewqQJiosGJtto63LvAfT2snSD22eQ1IrsYy3I9+pyZhQqRQFniXeXr3Pn5YBSolu8Z
qiUnlHp6AHMDW389gO2HLgcFy4b97y5L0dZRtLUgscsuGEqBI/lmpSL9r1vKaliqZO+3IfYtMrES
j923mlrZiKXP4FuxRgtL0kbIm7KyDPP/9jw1/K+S6FPKhy5xNNKdIovh8at+K4trwDdtpz99y7ba
CMO4al3wwxqXcD5ZFBWfnQCgVXV/wfCOBGM4RAiH+8hlIwlW2BkELML7cVOg39TswJ7QObxaWJHe
WSC2heswsySNSiulqNVPX7tC9HxiIImB2K0Q2tr7JAQ/5iBblRU6UMhw5MsjRC13bjnChk2m84I9
1/oj3TJaFnfvZGFVM+9WkkJXEbE62iAw7kp0ckBXDn6Mq0h6uYvZ3nHWnBCbGnhBwA16clh9D8Kh
R2bWofnTBT8dXGpiCCTGcQyxVT8E0c9QES0CPGlFSMRcWP/cfxcMWKpR8Spdd27yBtsZmi0+CfsH
ZMwjjaZDX6AHiViYUjzKYBSFs19/bRxr+roEYkMLTl175XjDw1rBmVrNoVU2W+5t1ALpUlfrD5su
1iPQPOiRrHp8ZzVktkKDkKsqfgdP2IkBdu1Nmet0ZApXR/z0k9eB69VplWK5eWe1SVPJUBvub07v
5CARmEY8oGLT5iC/pujDP+BNx0i7ILoE+aVhnksPn2juiBHhQews2n8H9/fI14XJgS9VeU7N4faM
724/xW8ETZoyOrlGD615zeJrOB7Yt5VpCW/B4BSOY3Ix7ZEVMLQItn+rbom3EMR3HFkQ0fgIJpeZ
ScTLkHLaevpyFus71O6S1w4UTq56RyoSSLCITq1Lzze2neJiWQW0Hq/R+5Ou+9lnSqlzyVZ9fV/2
u5tzoZWoaQQNxjJw5qXsASAzXRsj3sqzAq8oOp+Yc1xDh+jpZtYByLK9PZXfpNkq/eFlmPJhnqnX
LY71Rai4gwionReN1OZNQiIFjxC9MlykTPgmKpt+gBq7mAwiyliMbuUxgvSLRY0JsbQvqfi2bse2
WTM3YZGvpooDmTfwHvpjI2CrxY+OzCGL327rnSgyWwR4xsidridJkTDG1AFU1D2ObgEK18s13SvF
kj1OEjZ1AyfvQ8ZvKIkRd47DzmUAzA5BzyH90OMHRGYlW3yp5pzUZT/oPVPqTEnq5poJRF4n06qE
0/1JMJ46CD/xhEZ872h89j9x1RgM5uIFla1rzRSmYwb2Fo3nfL1cZun+kye+9CjhM+t/GiQ4YRwg
20jaR1zL0w8FjtRWtfAWUFi2dwXwlEacJdOTz9Ktea916zPdmHrDhMmimdJMfzBwyK5Jq+KlV/Jk
O+2ovho6ns+xU3zRdULrM0VU1Bnu7/IQUSREG9N0b7j6H5ocjk5Qoc+jH3afMapP5BuT0e3KZU7o
gFgSNA+HyK3GqLfxV/YOkCLjR2Mo5Xb18WzbRtUC1QIw73prbSDz6mi3vzaqGbl2mFap03XFn0wP
xyqaqYv1bOSTlCT86V70X/SdbLjH/knSYKKfWr8HaH/lveTeUoK5FbbZOPBiAjVRLLoTVlK3Nn94
+8k+i53y5KTyTyX+WCNyin5TM6ogtHvGoBpMkmoiCq//2b9C03cJLPo6GZY+VI6OOVntMfdqtvsa
DZcftXzK4/rOL7fPzEr2xY5Betxeb32equWO91OO8oeBj1yiM551cI6jdwi+xnvLF452+3ynIIhH
sLhTRowQEeTZUCtxOIQnalG7CQQDus3I0Dnwk7aZdKIw1BohTZDAcFHb4TlEPZrkTm+61fUaRG+X
ktsxPUVJeDVCbTQHisa0eaaT3n2H993PGtV3L4xHCrtYvUO14zk9KADwVMsinnD8tODnul1NvdK2
Jj8dPqt7t/KMYDpX0VYJ
`pragma protect end_protected
