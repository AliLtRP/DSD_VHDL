// (C) 2001-2013 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License Subscription 
// Agreement, Altera MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


// megafunction wizard: %FIFO%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: scfifo

// ============================================================
// File Name: altpcierd_tx_ecrc_ctl_fifo.v
// Megafunction Name(s):
//          scfifo
//
// Simulation Library Files(s):
//          altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 7.2 Internal Build 134 08/15/2007 SJ Web Edition
// ************************************************************



// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altpcierd_tx_ecrc_ctl_fifo (
    aclr,
    clock,
    data,
    rdreq,
    wrreq,
    almost_full,
    empty,
    full,
    q);

    input     aclr;
    input     clock;
    input   [0:0]  data;
    input     rdreq;
    input     wrreq;
    output    almost_full;
    output    empty;
    output    full;
    output  [0:0]  q;

    wire  sub_wire0;
    wire  sub_wire1;
    wire [0:0] sub_wire2;
    wire  sub_wire3;
    wire  almost_full = sub_wire0;
    wire  empty = sub_wire1;
    wire [0:0] q = sub_wire2[0:0];
    wire  full = sub_wire3;

    scfifo  scfifo_component (
                .rdreq (rdreq),
                .aclr (aclr),
                .clock (clock),
                .wrreq (wrreq),
                .data (data),
                .almost_full (sub_wire0),
                .empty (sub_wire1),
                .q (sub_wire2),
                .full (sub_wire3)
                // synopsys translate_off
                ,
                .almost_empty (),
                .sclr (),
                .usedw ()
                // synopsys translate_on
                );
    defparam
        scfifo_component.add_ram_output_register = "ON",
        scfifo_component.almost_full_value = 16,
        scfifo_component.intended_device_family = "Stratix II GX",
        scfifo_component.lpm_numwords = 32,
        scfifo_component.lpm_showahead = "ON",
        scfifo_component.lpm_type = "scfifo",
        scfifo_component.lpm_width = 1,
        scfifo_component.lpm_widthu = 5,
        scfifo_component.overflow_checking = "ON",
        scfifo_component.underflow_checking = "ON",
        scfifo_component.use_eab = "ON";


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: AlmostEmpty NUMERIC "0"
// Retrieval info: PRIVATE: AlmostEmptyThr NUMERIC "-1"
// Retrieval info: PRIVATE: AlmostFull NUMERIC "1"
// Retrieval info: PRIVATE: AlmostFullThr NUMERIC "16"
// Retrieval info: PRIVATE: CLOCKS_ARE_SYNCHRONIZED NUMERIC "1"
// Retrieval info: PRIVATE: Clock NUMERIC "0"
// Retrieval info: PRIVATE: Depth NUMERIC "32"
// Retrieval info: PRIVATE: Empty NUMERIC "1"
// Retrieval info: PRIVATE: Full NUMERIC "1"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix II GX"
// Retrieval info: PRIVATE: LE_BasedFIFO NUMERIC "0"
// Retrieval info: PRIVATE: LegacyRREQ NUMERIC "0"
// Retrieval info: PRIVATE: MAX_DEPTH_BY_9 NUMERIC "0"
// Retrieval info: PRIVATE: OVERFLOW_CHECKING NUMERIC "0"
// Retrieval info: PRIVATE: Optimize NUMERIC "1"
// Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "0"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: UNDERFLOW_CHECKING NUMERIC "0"
// Retrieval info: PRIVATE: UsedW NUMERIC "0"
// Retrieval info: PRIVATE: Width NUMERIC "1"
// Retrieval info: PRIVATE: dc_aclr NUMERIC "0"
// Retrieval info: PRIVATE: diff_widths NUMERIC "0"
// Retrieval info: PRIVATE: msb_usedw NUMERIC "0"
// Retrieval info: PRIVATE: output_width NUMERIC "1"
// Retrieval info: PRIVATE: rsEmpty NUMERIC "1"
// Retrieval info: PRIVATE: rsFull NUMERIC "0"
// Retrieval info: PRIVATE: rsUsedW NUMERIC "0"
// Retrieval info: PRIVATE: sc_aclr NUMERIC "1"
// Retrieval info: PRIVATE: sc_sclr NUMERIC "0"
// Retrieval info: PRIVATE: wsEmpty NUMERIC "0"
// Retrieval info: PRIVATE: wsFull NUMERIC "1"
// Retrieval info: PRIVATE: wsUsedW NUMERIC "0"
// Retrieval info: CONSTANT: ADD_RAM_OUTPUT_REGISTER STRING "ON"
// Retrieval info: CONSTANT: ALMOST_FULL_VALUE NUMERIC "16"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix II GX"
// Retrieval info: CONSTANT: LPM_NUMWORDS NUMERIC "32"
// Retrieval info: CONSTANT: LPM_SHOWAHEAD STRING "ON"
// Retrieval info: CONSTANT: LPM_TYPE STRING "scfifo"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "1"
// Retrieval info: CONSTANT: LPM_WIDTHU NUMERIC "5"
// Retrieval info: CONSTANT: OVERFLOW_CHECKING STRING "ON"
// Retrieval info: CONSTANT: UNDERFLOW_CHECKING STRING "ON"
// Retrieval info: CONSTANT: USE_EAB STRING "ON"
// Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT NODEFVAL aclr
// Retrieval info: USED_PORT: almost_full 0 0 0 0 OUTPUT NODEFVAL almost_full
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL clock
// Retrieval info: USED_PORT: data 0 0 1 0 INPUT NODEFVAL data[0..0]
// Retrieval info: USED_PORT: empty 0 0 0 0 OUTPUT NODEFVAL empty
// Retrieval info: USED_PORT: full 0 0 0 0 OUTPUT NODEFVAL full
// Retrieval info: USED_PORT: q 0 0 1 0 OUTPUT NODEFVAL q[0..0]
// Retrieval info: USED_PORT: rdreq 0 0 0 0 INPUT NODEFVAL rdreq
// Retrieval info: USED_PORT: wrreq 0 0 0 0 INPUT NODEFVAL wrreq
// Retrieval info: CONNECT: @data 0 0 1 0 data 0 0 1 0
// Retrieval info: CONNECT: q 0 0 1 0 @q 0 0 1 0
// Retrieval info: CONNECT: @wrreq 0 0 0 0 wrreq 0 0 0 0
// Retrieval info: CONNECT: @rdreq 0 0 0 0 rdreq 0 0 0 0
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: full 0 0 0 0 @full 0 0 0 0
// Retrieval info: CONNECT: empty 0 0 0 0 @empty 0 0 0 0
// Retrieval info: CONNECT: almost_full 0 0 0 0 @almost_full 0 0 0 0
// Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_ctl_fifo.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_ctl_fifo.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_ctl_fifo.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_ctl_fifo.bsf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_ctl_fifo_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_ctl_fifo_bb.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_ctl_fifo_waveforms.html TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altpcierd_tx_ecrc_ctl_fifo_wave*.jpg FALSE
// Retrieval info: LIB_FILE: altera_mf

