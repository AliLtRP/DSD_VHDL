// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:52 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
U77vwYvnAXoh2NT0OOvj9Z5MAf95zZwZJaRUjI/K83lP2ilVahIKgegscjUV6N10
wVaVFXhO0FqcOOSo6BeXYLdOKslAzd+Q+GfT6yG1cQ/g6F+zf4W1buFMy53yQWK+
qrh6URkWBZAidTm52vGJh1dtEdBWrpoQYa7sbb2xPEU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 39584)
zrIC+cUwF2Me32H3VHdNxNLbzKFwjc83a0xCkwCUQbLDL2HgyCTHH4vC4eIbwZ/o
LjeC2LidkRTDIsY4cgdY5sDbx1V80HYuMgpzS9BG00/N6YuzOQWOKV2w//0+IhYb
crl4VCzALVqGsLLRwxlqyT6vI1f3Z4a4ZpjFjefszlE9/uaXskUOHhDVEWeMxfIW
zx2/kvMI2OpLU2dkgUPyq59/MZvLyEFWX9r+OE+UJTwCK34rVPxre5S2cpySSasd
SpaYMnnCV59brY/4qo7OrWQrGEaYGYzQczYdgDxTX6xhlkMZ2yJkmJDFj2UdTZs4
2zmYR/A8oLq2ooQFdyH9YyEzxZhTGmGl9+nJHW/Gzp2F9vuJYBbwre+ybjE0Tnao
D/nS5JRX3U4wBKuE+Dr3p7yX5LekDR4m8denBePCzbuu+wc/7Dx3246+ZWriXCje
x1k9CVRZtp0jWm2Y+tB/kzqFeUT7x+kZ8D8784q0CgWyE+OG5QG1P8vsX93BnwjJ
Qt2a3lH/G2IQGEJMcn4609Z0HRhFyJS/8rkjl+tCPmuaY5DkIs7JiV6Y/PgI33NV
S5NEBJrpLt7LI9sfkRCoueHR4r7QDXReRjBAySFs3BFwuVlMJPUP+hRwYI84le/b
NYaKcTwYajqwGGv1Zqa7Vx4v2bNGkr5SqVmWCzojgOUCdRNGAbHatj+Nc8V+ahJo
TYSjSxr4YVajhhOpt5XznEKJ7UbPxoFi8OLc/JGhldeNILO1kbpcmWa8XVpMLs/i
yDl8YyNEDBTAwkze5tDLLQGPSaF3fOprmvfb8jCSXZs7UMaf80tS6vLzCYblP74Y
c7P1CgYCtJHi/VwGLQfMRO2llxvDO7KUsyiRpC3Q1VXQd+mMIBKZMzEN4zSVaSj1
22NJzTkV3rWZTjXhOR0RnBXPbKXPHU8zrg/GpMJDHHLTdIrXqQY750gj3W9CsdiK
vB7JGJvXYaWMLa0XhXLL8B1TSYj69WOjI1lc1Il6rfwMbVgO2vcIMOI5WE663NrM
z5aDAFj/KG4iC/KFy1KuXCLOoRcMCFzuEkRRRgbeGO4425q+vDhoS472kCOW5846
imU8juCPNfc4uTQTTGe+LRFryhTob+4y7+hLqYzOaPix6AuXX+AAZ9bYIliBJwPS
R2y9otyTcwIYnWdw/PxRY6RhQI5n0BoQJwZo2V2HLdvlWFKNkEqaPnr8Ov2XO+Bo
4kmOnp1qaGZRBmrxywDyORLrS5mNvVw4tvPzxrcJ4+I667GDQzCT8FWa+KcgXfja
q7FqenozfeVnOk4BaxejK9x0lQTxlxb1X4s2m2O5Va9QfN+HS2rAsQPPqKgaNGCD
YcFP0tcbHGH7QvveE6zTitAAMTQZv4K/npTlbuMfx4rovIWmwt0lQAcvmOT4dC0x
fI3+Mn9sRz0h4bWl+1JHgRN21IifFTWCTRatcyTHvFDXqO0UAtJ5Bnyk8Ghd0EyL
CtqqAVOKPxradfYvl6ssgCLJn3rL4x2OLBr245mjvxPNbq36PpFoeBEq2xc2/OT7
hrmVsiZKeeBPp8I5lfQ0B8bm2gIf07I9ccV0BI0AvGeMMw2h8bHhh/IPli11qNBG
CWFWmUmPP87QUasyeApsfKSv73yhWAs/4orp/frkaID93qtJ8e7IPjvf5FQGxvaK
3jV6kw9VOjA5Z6yacjpaVPW7RIRfCdHz4h8CAU+SBMG8LsvkY8+aXE2FoLNvISzZ
FT9uQWqGFRih8BiFBLPYI3YNnjzd24wqg2zwj8Web0ONPoRaFr22RhC5uqiPSd9/
ORyAlH0jSbwddDsHg1s7LgRKMoJxvMBsyAE66zuApuH5LLbPYxP2EBNaKxM61TXr
NKmim3yMs5+FLnpfBGzAIPtWdX7+qWC+CdJ6hAG3NZGQDtBxPKMimAnsm/ZUAtFX
WwiXnEQptDgmPbZDt1UqAaEIDhWme7RZpONh9CTEOQ6xYxscLu4UFqLYmAargogX
0z50lvvOpcGpInjDf01OVYYNtFApnMXnHcvKKq6gbmT76kmYZoTem8tIBoDRrwDT
o1rgxZiiywnC7uxZLy9vdL98zpxHM9jEVKrXH7N3kPcPERxQVI17mbPCfMLiG3zM
dtswC5tam1cOFYigREgyKXB51GjbdJdBdfR5B71u/RZEur6UduxIm+MyayoCkpqQ
lzoEb558ciMXBnug3vCAFumUSc46CNQPc6GTlulqefCIX4qACg3XG6vuAmcQeF0C
lCOBkF8SV5p+7jCoK35E672GV0bGqM5bzm6TSb/lzI4mZJEPPCpOhTiVoLZS9MS3
QdjMWY0L/haJG6N83Zk0eYSUuC1SbUWr2RS852WAYjP7to4WWns9ua1jiBT0boHF
Bgmpw8UVQycDbCf3x9KEjrbvABH/Chbwnm+uOEzYPDKIFjYVwrYvSySFHYttUfpM
OvGRXdVJn4inJXh8TIHkhrY9u+HhpoG+hiUCJ5GZT7HgQD9oyK1qmFEj4/fvD6Af
VDV53I3yEnS0lL40/axP4egHosBqNoUOYv/wbbSJyQBqqw/6Z4XZiLCblbruxtVB
exsaSzFoBkPm1ajZGVNMBHbBQxZIR1drq0Yz417iiehZMJzES7T1sX904SRAE2KD
SvWsMuU67QmtcA3DYoWpHC7mqFA8okIQAzfoCEffSYhvko9ZE4rP7KaDSS50mXc7
Wp93hhhR3Ivtj/MZHKKl1AS56+vxKzaEW8sYPy/gRjENhLZFjEHoR+nT/zSv1sMw
hVgJmGWzaeZxv442U6rvVYZ/IHNXvXLWiTPz5q7N4Gma5R46BiHGNEtpW6C1MK2a
vjuymmvCQ9Eg479QSl5OvlDN6Ax0nnXT6orpWmMKuGArjBu6dCF7GkaghwhTrB3A
YLkzms+vdSPtrRDveOYk11xPTHS0MgfR4X/yoi4KULl0vwPletWnZzLDcngbmP16
+r/DgpHS6tHHvL+82HyqNUrV8dbP+FhwKIZV0l2n53e06moXdNL59etGyrNDRxBx
+lYsUe81DI9eOp3qXLNd43EaQ/WZNc3BCQ2sRPbO1DhBtl7tHvo6PI07karOm7jD
8VLDy/Yrp5uFu3zaC2BzeNjHNH7DlzmhrJvK5CEb3utyhYh9Zz8OiQmUf+TJb0sQ
qUKAfeL8bxVuAKY+ufpnZeT+eeW9aTjcHJtB0XVs+H59uCn71nPBxpRS59pmc+R8
0BAWnEaCE8qGO3aeRRzG/AGpE6vh5Ekf00+40rBZLllHYPRBupC8BEhd4OcRGjls
QDWDQjOAE/nx/o1GPuDOUF/7Y9/fNM1QBbpeOtLWxClSG31zhTcSOtSUBIhMAshV
6vaekz45NqH+wXmqG/Id6EWmvyHMOVSg9eB9YONU7LOVPqZ1IfUsG60oBL/LaqEk
gdK+fZNvHAULksrYR+RJX1Xexu+oqoUKDp2Q1E5hFhkSCm1fLZ4Vu1ucadFX1qhz
PgcxkxpmdXKo9Nt3gaSQH57fG1P1mFZaY+kAnkeJvY3kHrWoR2VfYu6PZjxqOvP4
Z+HdDu0W4RduoU9SgPTwAHKuKkxfYdCUeHTmlftZC5bofaiH/H95jny2Ut2eH5dC
+/A2nojePrQfjAKpG5Ug61g2B6KauDwoIYebmEdUZmSrLFncsgAdyOYyfX28xwXf
Jhy9fP/pwThnSOGL2bWrCp8yrWXKm8TCb+qRm9Spr6uZC3boAb2xgOuRB0R2j5im
eKTW+OSJhq/+mpOfwWL+0Z9LkbX469dJFvIZZFc5I5WomgfADUZyxoaz3cgVVsKr
+0tsXhtkTqCzMkhDsmwsVKJ7qmpGOYDaQ+1BkbhDmoxVxWX5+m8Am1dcdlmGjpAD
FvQtV64CR8FCQe+nr3dYaaSuNYpnsnKKX7+dwJ/bClWPJyBcLoTuzP+Qfqpxa/T/
0xOdXeCVCCQM4xwJGqJVElwlPQ+6sTbrox2wb9CE5VGHOi4Mn5A8HwsW01P4Q1wU
fB9+xLnoTFqjADXuFUGzSxZmaw7G46H6PIjXTdETp4AmRenw0pbhKIp+coIX3scx
ksjkxcVePxl3XU39HEjlA6i/ftLWlyck6Yw4CmFjd8GKGIuxeAb2Tslg61NJxnDo
5L1krIBC6zhYALhFNgM6XfFRw7HN+jJxVJh+Ly90RKJcSH7SpI3Yqaf2iGwvDp2M
Q6lSJXqpSNprlACA2qghn/Hm27aBU0DpRn6wAUvxLv+x4gV1Lzhs4VDRyh0iLIBf
qKN+Q/FIh4TaI/CkWe62skxP/FjEd7pxiDRr6oxeUY9YufKw4tQoDst5R/wAWeGS
xtl84D/xkazHSXb8CBz1hspuH599eergBna1Iq9U9JK584TtyC77E5uowZgSRZA0
QpbBCS/FP9B2+T2Ur5MSJ8nxJSSEARMTvNPpDPNg+2vF1JHxlf64YtbqY33ru2mP
4jW6fIYI9Bh6cOxDFTtG6IkeE32b8b77CUUu4+VdEYjmX0RwKvZuQOkYvQ7m3SGA
SO3d6D/Cw+0Qw/M+RvcUJiVzVMQFSOdxhA4GbANUvkbMCSpVj73EbP7Ooj8tRy74
5z9oFnkAZw28mJpMCPGCGnYOekjvsJGf84BF3Y9ViAgGrrnk3gn/2dT19cFzqygx
5r/3PNyhDQuHDrAUBxchDsRp10WVePGJ5gq6/koJp+K0lmTs/MgoX5XY4yjczJMq
DaiNdMqmWi1ED3M3K4Uj4rsmnERZtH6OmNeiyoIljVsLhgd3yjHLn2ugTVOHAK8Q
bEhqcw5fbQjgLHzPQVa94yMonY5s0uqDe6c11jjpq1xgDIg+7hkte087umzFvaOD
R3IcBe6Z6WduFXBiBnBL5MZI/1MKSyKUDWtIiG7jkdlnRVDt9fKRGPdcaRMx/Yr+
enVtuLyqJ9Aqh/DXQ7NBzEF5eRp8W8H+4WeSWiryJzX+qoJ9wWpNsDGsi3EaWvXe
J19efG0eYlBIMbN6tVZART397AnVdsdbXK0aNcBHAoA4ACp9jBtnWC2udFbxaUEY
nDoajlD3GT2C+4mkPNn9Biuf2my6Qlevd+Je6bm5jiGxcJ25yxCMInyJfeauyUVz
VPdRyZHYada4TFIZ7XIw8h7U1bZEy9Q3CfVbbbJRTpThfEgbA43/r3i5661PGmG+
mkUp24nDFd7I5ghq3h6M9S9zpwvqRSSpglScPfzUve23mDSfgt9LZ8rmwyqkqkH1
HbVmNd1Xs/tg75IXUPluU/vUgAez2mvOCAdHGKksx198zqqMrQr0baXDC5izbM3v
XdMmOEZbrc14qHg9cqz09cnjgZYiLundrymXfVji+CBXYa7TZSL6xb6AFZZ0UBzr
GAkhv48CXQDIjixvfV/ADorPn1c/ux+X8/Jm5tTCf10rBoF8AGeKtAbgLfnRoOFw
RiEW3bzjXlljYqYLGN5FX5O6mC2UCuSe62whnfHPoboSqIkNEDPi0l3stWuEzYx1
zn7gRU31X6q4W0qdNkxfw/osneZTfVfKNKtIJXQjZqrJqQbYbzosQthw38l0oInR
8ZDDed/JuQnpkYwt1ZH/r1oNfJJZdusubgYS8nAx+PdyBLzCv+06YipAKdFjvLtu
XpY99+zZx3py5JKEJKK3TRS6Jka0GpEjZZ+whSqT2bM2lC2NUA302YkMEKoYWVZN
sSg9wPkv6uLfUoGZcR/1rSSa2faV1aAKXsONpEF+AIVsiJC80BT1Irho7ZvDY1jP
lJLPWKD0jkaoJ9FlI+vsmVPQRaxMea34zHDIfz3vv9N8QmNQn73tAgtqJyd8NmKW
URYXEv0sIO5FrFE4L4RM3YTnt+eBPKoDFyrLo7WqNclOa4bmPxiwvtxFeEgnteoF
6MPRiIFUWvn/UZqjrRA5PckqVXzdSFfFnBelCK34IBZLUaoiu8IfI8xFT0FozUfX
60A5KOJWiAx1QKriDItoJ7C4h13p+aRAAM4OcPPzGALPAeFrU7ILM0d164lK1SoW
RVuPx7I3dcOe06ABA1/XiNch/mF8jvXVcuKpJUPlj9hU9pCJL8T22sLj59+Od2Pu
/rzPVI28PpMkYTedvVDCF4TLPlfXCtxRdC7LfC6sq14NIjcDCHO2yX0W+D5TmBms
uV3mz/bec1wFfzReNdcKyYE5gT4ZZvkZ7AhY/dfuYlIRWio4SgdtPAMMo+Ga6H3k
N8sVyviP0aoVKphi4Vw+0HQFulQZ/LEM7eqwp4coFTrghmOE86/Dp7WbZcIOYwR8
L/r7O9RwppSrO2TsR2KM5DxkAB5qUch3QFP354RDAS0VpVFWYZFTJX7sdQ2w5xdw
wv5F5NzCEcnrNy8iAZ8UDd8BJRxkOby7Y4jnKrbN5mAVfFPtOlF+5s4KB8D0KM+5
8WFqfYLKBCoBhM4RwoIJrw2dng5759bV1I08mTCW6OIp8iVKDA1hFiPVzk3qKF/F
GBC6YluUzweCCVl/XJWRTXfB0CBriR0hNTZdN5N5pPXBhwv3xVf5Th9liLmIM2fH
iUzAZ0nuLP3d1cSQLE6CBFiVHdAgWyxQOUFbwhoMYMLt0MEcqGnNA6OJUgJV8Kjb
9YQjh18mDkZ3OvVLYbT2oUSDShKlwgxo93KUMOObLi6l2JfpGtZtKwrzWwgc21qE
kpEckkLwnfMUhr0Gh8YNsSdAsM6doRPChr03xSFgM6xAkczRGsIyIw5SQcbrhjYD
m9VDcSHsHjAnzCHPhtaoZGGhiGENnucMC+gQjagTtl9bDKFqhsnSnQPFGVs2HYmo
/RLlas0Z1LCLsHljvI4HI/C/Cgfx+FwBidm9k+JtqEQdvUpv5DLr4yb9GemFte2k
ftkG3kagU0A+X70CZdKqANi4mARqmcFXgOxoGQrQms77QGTWZDHL5jAeEcWzpTLO
aPSzaHsHvCH8Hr+KYA80ToJG71PknjsatLIijlwLmuxHC0X8hmivoeC19yAou/2b
Yb6kONjjk6YJPODlSY7HeHXuI+9OXfNjpcPY7i16F6jnBFvBZi3GXcb0FrK1/fYD
S/dojFLMRQC9PDBcmK3E+jf0oFMOHivldc31cj0ofQisE/9LBm5cXagMmFaQR14z
gEC3bKvmouVDsiUutnFnoaLTjaUIamimujPW8zzrTEpr836DQflLWE/mVCxLvoHy
xFJrNHn+4ILOE7mb1Ph7dUmpwv25L9CH9ZZVcotVptiEdriunBp0AcNnKGNNM/CH
CfIKGNP4p+tz9ywEzAedtF5AKUqdtCuMLaiYoXFxxcnDqKq6e2P5s0HGkQQ54wcb
C+4lZtV7EmSJ4HZCa+WcfmrG0iOV9Gy5ubkmjMpayTbgs7t+JxANjcFueOiWpZ9u
8Ofwu+lCqcbHLptj5I6jSspknXQeaPzPO7LYRFugRDuPNP2DUSp0szTwZy3Zc0wg
TRWkEvwqxnTjHzAWdRAm0+bNBHlH/GLiWa6UT83n/6RkZGXYaU8t2mCl/YpNlY4C
jK3rLeE+mTa7V7r4bmvqKzmJSIQmh1Mzlpb1NvB2Auoqtr8exyAZxnp88312nn/9
3OSVJN5xDlru/ge12qh2uibBj6Qf3knOpxWa+dy2D6ElyYI/tA+WEWb4a7lu6Ktw
DN6cQY8x/X5OGTDSUucVWX5FgnYrkkbPvZI6KTyf4vOr6DUu0Yr2epwltlQxCPv1
Xs7LsYUJxSy5P2qr3tg0/ZBVHoWpZQnH+a/wkzwp8co0GzmChMnkEqGmj+D9xURv
LXer5DMmz+617YCVqNJH3lLl1yYZsNqkSAB0tUqhPYcODNbWGU2wnoua56HGCWvj
g5hChDLfV4ANlEC6TMzyyjsCyRwBZnIZHLoVxE2uXqsUj/SK6utHbIT+oJwF5h9/
CaV2ogsICJ4FRuFVXNaRJMa7wXJrEcT6jJE3P9sSfPUruUVyO3+nX8h7XHWD1ZpK
UPvEJOOFDrj7e0N/IzzZbYewG+sbkK7nWLH1l2Op0KPI8Xn4jwJrbxZVJ2Wv2D3Y
RVyhXzxugWjVNh7TbPI53Ai+Fft3orgMqBQqhPTJdoHkch+Tovyix25fQdUqxHJp
tHT7fCfMNjh+rCF4+azSy8PqRckXKMTQgcdmvMXuQbt7cjbMTdSyEhHpqmWcz01l
usYNy7x8rAmedvym8QmkuPPOHxNXetQxHnTSCdrBW3AlQk6XKQH/9nX4U6/KZBnG
RI9z+/9tuKC8B6i+hzjrJ0NRRaV7cHKG7g1T5tCphfpltfvK630foUioKXog1rU6
nq1M0CWZBwErlIjWmeZUYGacyvl2K/AbRMnRSTr+6Z2cycu1Mueppxw1HGifUdZS
Q01ky6btx+I4hudJTqLO0Mz1Jx5RA9hrosTlS2dAYR+zxfuVEoCyPHLljluPpD93
WTekfYTTJqyd+matHJjFW/AvGIQ0EnKFR2Vc11cC+3EGtNOaOM/T6WZtbu4LdvYK
ezQL6CpEVm27JShrJAcjMXptF1yuoyc+khFMdUZLJe5kZnRHeAQ9SfyWCX75mZC7
9TbUsBmYDZ2VBg0jeD2VxfzHit5EoMjSkhVR3s3RztU8bl4dexPgiFkqRzvbnIKR
vB9jlY7Z74tTsCGbVEzp1nHIWCGbmteYYtp88C/SHa44MsOhvn7fh67nrnb+U/U+
9Bpd3v+sGOv69LOFetwa0vjLJmWonyx5UoVtLUKMzsbEgjz54yps6YiLeSpQrp2i
GjnklwojYU7VChvG7x6xFjiYf2EtDNTt88/+J80R+pNzS6wjaNFE2HYOGftT5HTT
ESL/Lu0yTyCPGfBaJNWXq2aiijXB2qKTSYAhnCgclT2ca4Dkq9Lm0w2VorsBeNed
5j00tl3Hu1y8M+P6YJgFk4UrePu6n6lNN6DqlLvl8UBULx357hHlEjFzE5DHugDv
G1Zvk5JO9IiPef+H5e+FoIuibriiP6m8uMb7eJwa07d82L621ku6YBIGVPbN/3AK
1/I87JTt7g7SmiK/lQwBBE+NO2SBb5kHGX32z9yze6oHXUgu7c+xfJjToiP8AOVy
H4/sb7l/T/98mzV9b8HgyJM17OG0SpkspDoRZ27Wau39v1uwsBIzT22ErgtTuDgr
DwHQEDm6NgvRWLtXsyf8uAmL4ldJUff9q7+wcuFxjHX8r0Qb9CyPyTyNNvK/V8xA
TNnA68ysIHHehU4qJOEMCxR9QFjfmvWYFSKnaTZs2yDvu6kGMxMo+DT9ZWb+qn5h
WLqmXHrXsnPQ5YWa8nkJY4s0XXeCNN42QF7oPdd3sXKzDE5QStKGK4e3zTEyGHfk
rUO52666ML448Vrj0AmgttyMytHlWxMHqMbjNrQwJjDCzeMOSJzlekvCz76iSALk
ZIGtOehb4oACyOgGFXJvRzlK1rvNtBr4TW8JtCxnSkYPOx9DuJV0NKgT2YU0PHsD
Id67/TcQwAVOOM+xEom264vessQbNXiO3gPrKqtdmF9020Dr5MUnVUtR7wZnBTci
jAOUnUTT1onU+rULu/R55/ul1g73IdAz+0bLHM3MkeO8+EuhtSPjWHOAbmB1r61a
Ydi3tOadmiSeVC7yGk1moZFk1178odaZX63ezfaVi0wM2E1nuQVdX0fPn/7OJxC5
FKlfbftkRJtWJsMQRpW1XHTXbeKZ+7ZZY+sTOXsCvkEfOHHtJeWNQnCxwwB8RU/L
/v2yokmwojCwxC3i2dDaVdKRGk3mi6p3yQpBqINGxUlrtxF/BWQkRkhuQzwNJsdK
iDRn9k40DDO3DnXwozBbLLaRKEe0pkRbNSgmxE31giR5iycHMk8KfnbQfzbzkHaA
0DtNUaaDuIvq4iOVeiDo7P0w8MPUeRwmwGOrxVwSvJXYFRTwwi0629RcndH9Opms
EqSSagopbjuQ6rUPwvA5TR5C7fL3s4R/Bh80nxoAjPkhQlPUtl78i2bb1+eavDUn
Or00MbYm7cBoqHnBbU8kEwHPGC8xNtazi4pd5OFksWWqUM/x5EcCBCXqRWC64FTr
BSF/yPGYvwpSUsgg7BNxzoX1jDtAa5epeLZYUIafV3T9thEibKLIAsd6QrECrFJ5
G/aKK15Wx14LP6Ecf9P7oUEYxzwkmqxswNfEo7KU/z9/0pYKEYulgK34Mh/3RN+g
9dcwuwUe+3fwF8QaQ1Th4XW7y37BJVtnqkHhgyI+ZE1rRd3Fhck84iZJCaFNh8bD
8rm/iRvYY5+qR8PNY7Bgz85GIF/wFtmJecn954ppcogVIl5cCuad6iLvR9musA0i
2NDsKqTZMZRhgA8dIH6tdvpHq4bx7kFzLQUMwVZKJooHBh8RNPyNcDRlaa7LO7xt
EGNa2yjd8YOaHht7LHUCHgNLbHOcFkRRET6RNKZoVN3CHUpRVVaCbYJVzKmTHs9L
3OE7HmJcQ922+Qqyy0FWYNTj7ANncbOaq08/Nw58lSKLBEZhFXHGNysZivxzstjQ
OxS5x33d/p8wdfG9O6+BEW9n9RaZdir0PdYKBfFOS46SaBxc+3O7pIRvWAWRQ9zL
MxCpzc+KDWPLhsiFav501aOSO++Mt0lBfAQ3++tlGNoThudYMZ7efdz1TftNp/VW
gly6TpAWZMGeUhtNoUrE8Pw+sT1XGA48lrecmpuoR6RxuUCiko5bfUpDnIxW8vRz
iruwVR3b9hPZ4ni4566eD4bJmlRCHWtEy/+dNpuDP2+leH2yLT2r/RYaidMliSBM
GVbu26g6Pfux94/0LN4u4lds0ElrCz26yW14ls0nKHCuD9gZI+Z8OqGCCxS+ZELV
mEHhhiMJCfuk3RCV84P84nU5qiepLz3B5bFByRMTmipqf4OHjDntmK1ledh0lJS7
e9cSYQsUlg9xR0mgDm4jmqqa60/53BfOtzjN1ooxeATor/1wLhXUkkOK3wH33DyK
yFAYfLgYsQtW2/eMbEbtsA4+zw36VFg09URLt0Ids+Gn6bGK7km+B1TeR6cuh97U
k0PVWIpkvYpQzbTT1yvEhnUYscMq1rO3uzKZUJyrigYPyMT1KJJSLEIXGQ4fqvsi
R13lwXO+FeUY8AsHPCFf19uNoohf8sZHF1YlmTDdF6hTmWByhRJYfmddcM9O4F1m
gJmOVFXmOAbh+33ffTmiJ/7ZPeknlEf/fTiuO/qtfsKAq2Gt596wj2Udf0AALKq3
SeK9Hi3IVIOJZrdhApvUteroU1eQx+SwVzqTAt1bxmKBIzcMPbloB2HpcshiiBPj
PSE/qqA/QciQ6nIPuUhxZsdpvr7rCn2pl6Z5OlViK9bh3nQcVrMbBGIE+PsDnXut
KuK4RLEjkKt2nKBRjeIAdacMg8Ms1dXuBhAiDkfIG7TXTpdBuuVHhIMvBLnRvGHv
PYikidTf/mVvQ0rH8yiuFrHUtVQ+mX3rN6Em8mFmXyeF3YaJfFzmMmEr0QS9wfFA
18jkmdIaMo1JTNJ6IOftuAcB9Tr/RrDvw5QL+OaNaS9pK6OgwsuQ2yWotsgdkGVv
Jqb1k4w/HJSWEdNNE1tR5FyEm6MOjfbGDOaKNaubLLXZIQWsVQxu39TYRI3LBa4Y
O83Dgk8i+O6H7QLm316Ay6cttmy06AOLiBABbK16Y03vJExeDKBCYgroLz9PBfVu
ZArAP3lvzPTwPVHzXX3kBSJvORhcyroKWsrkmkXxUhr+Fe3+BjqMBnITC2di2aPf
g5Kps3JmOaAcS5+NHKXAQEFgujjfcJlpmVdxPf4hYWSNoZ0HAikU0LdIm4NrTDMy
uiopMPgUFAjSfR79a1UiXaz/oDb03W6Q8u2S5yMQ+96MgGH3QaUTCJe3tXHkWuVh
15XDyWwTqlPvl/SqF0QJOU9d+wvYfZWqtHMPt+ylPy7XZNh3re2WBhyj7m7peZpA
ZKE9ZlFzVUCLgOYUVodEe5P7x70RoL3lNhAmssMw+Q09Xr4hYt/DaOUmV4ZD+XW0
FOUSU9nkMNm4GoiLu4NloLf0yQ2a1vtZJBPT6rXRbBb+B8RVvfC23NMuL0K3gvXC
xCpP1XFZ6QM4MXjF4IsIvQ0dI6/tmiGbYfATWNktDNsOlZSjheK8Rpe3ne7/eOzl
VgP+v26VHBoTi3Nh+4obD0LQlttM7o/Z8uXk5U2RJPQmRL+x6xCQeoySTqrYgMTB
j1YmykW62xK3Vwk/+5WbTc4lzBrbph/6YZxj6fBNd7rQ3mhhloxPFh2Dc5cpUaXl
CYhMsyFxCyBeTV+GtT7roj51wmFMcsx9vDQ0EG/xz+dfcYJyN39ZAWo3kxoNnNN2
+SyT2+Bj1bENtcHjHupFvnBuCKTySqZWye4jXNVmv/TIChlOI3pJ9V2HFMTPphfx
44pbXAht4bfOCLHzyTEJR3fzxykYIxdvkeD7bjxVaxvRXhHYVxIG8hKT/icxI1PB
UdVjXo2vt3FCs/J+BA2HQyXwVBRVbnj8pYU1mwG234NB9AE3TToGTYd3K8/GUGeJ
a4RixMHQnjBUqU8oxRWDNvejs+/jot9vz+dPlm6rBVL+ivVrJFEmL3ntcwRpcz3O
oqAY/IniKX56Qt5vTXiFDvTZZphPLPLds4G3HDEouod1NujQlxVrbDbYYwQKGxeF
y8CndvIt7EOesO/DW21lYLAIo1iBpqNlqiaeskavAc/PHgHp5//AeEq8wpjRUBD4
SOpDgVwNejxDA4w84JxdnuwDm6xELbCYjl6O1Jy9GMX01w2hfdJfJ0n8Y6iCbX3s
6CXYV55cJQmapdj/kA34Xg0ehCLAxX8SOuQkZanYg5k2l+8ylnycOoSTIqg0pi37
P51kqJGo9t+had0/IHozBB3Kv41CHtArpzSy3ZEWKXPK8cnVjaE+1bxmEEGG4IpH
lKJVGmm8vvetQY6aavVtSaBCuGQE1/Wy/2auAnjKB2kOQJGsaimnJyB9bWQKu8ht
D5v20y8EibcJYGwLmGmov8JY0lBvqF/mHG6vKKi8YFyGtfoPVRCtHKwhyPM8cois
zoDVNoETPEWGGDOAFVeEkbE8L3GhnAvHzGSoJluXVd2ufw4jABLnD7sqeL4VuGmo
9pnV5X1SCZfJsD/6E10Fa7HjcuVLQ50Y7eHJk+JSiA5FaaBO/DhEhRBtvbHfDLO6
RwSo6fv/XlpC6YWISPEIOSt4soq1j+q/BlRfoCBEyaYn+7NTW0NDNJywFLyQsAwN
brlOYyhFcrYm7WWW2NouRj8Ct9X/mtFhmQ8EMKjKjXF2TTm1t6l6xYI7m9L/6aEk
VwjVhEzUdel9RR9PwrZ9fuDLSfYjaGdSLfR7XHUNECaFIk6VQMLStqrMRHDl3hPN
eyf6kqFMeKpliPKnurHQQ2Xi84U2Ms6JXqY6TgpS+v0zrupo2bsg2pk8MTANipxp
RWS1UHAx594EY+eCbWG7C66V+8PUA+ovAdV/ALQ8Jy8saS/wfxhWxL5sqP6/PpPT
mIP8vac7gF0mvvaIWFZLzOR02WqCCm56wDeye55EhF1pxU/MbokND406G/yIznJi
ZNEZbeDsQ+D+LBnrW0lReh9k68RVdEgYBBLLo/jYnKvXCth/WVnTHAGCdgFZMKRU
oyyxj8VY8vpQaJ9Pm4LuOPOYZQ3t2i6fgbWVrkWOSxu3QR0nMbMTNhntyeligDz+
j+nAQoLXCGP5pjB3+CPtvt0Eq8exCCg6INDv4ZkPrRYw2iXEvhSqtR4AYMzcodjL
qOwd+A3xAHJF+x8jaPLN/ysl5WVox5oy99GP0xRBXF6ElgBPMRoAjFgxEcSTdblI
sQD1nI9WIwUV016Bgp3nQxDqiDOaEs8/DiFvkvAwKUKAwqY1K1hfeqqw3avhEAuO
p0f09SnMGX46lIPGHZDnNF2ft0hSAxGOH2x0fDwxQEVMcRIgVM4CrAYotcefAVRt
wo+PFTob/1k/g1uF6VirTMIcCzL5zRul7qOOzNa/7N8i1fGhx0uNyPSQT/K3OjYU
pXtjCorlFjyFF5qgsSAr8S3fDVTupGxeKOsGB3nK1UvmI4vXLZ9y7m7fb5sH5JTZ
6a1eJZGKVAT4Uhn5MQcv+9w59P1UFnaDbwWNLZ9KfNskcOEN963ApRsCapKBvee+
hsGHqhnJkwPRq/ChCvJVzZcmfTULXoXbRIigJ3Vx000yKxJyUymT2s8m2WNUFHlq
EmKs4M3d3Av3qu4zIU4LzWILjgM/WjZZKvPrV2C5WK0HGVHNncFrICE0jQXWqiS+
LAT+w69bABGpdRQhzo5XdhzYo3SAZ/Ra5dfWW4S/RtllANcx/KoxajHLtGKW6DzI
T4T+GPMdhFLO3+a0Xljk9oKiYMDhqJ/Jco0b5iuFTy7Xs6o/hGwctnr53EywE4JC
vx2sw/Pa3efsXqfwJ8g+K7Ix08dM99FpsXaDXlBQoZvleQpiIhkZa2SQfNZSsIEA
12z+dJlaFD5FFKEnuf4/XHyyFNJl8Xsqhb1chMOsHERvPftttPmZqkfOmQChd81X
no89BiuauIxXrTgeU+D373QwdCDqU67hMsjnquNP5+WDSHGwq3CcmUE3ureJos02
HUDhojYl7MViq+5fSg7uykiTZSvvW/CYI1iucRyCXBZbcZrJTVm6TiOGOhF+XEag
dKlQbOCWnMppn/n55m72GmF9DWnI31GQP5q0WL0o6QLd2p1qRhzOtQUOhdocPhjH
j4jzIB2sd2pA2gsefGeYl5PVOAjTrStZZmpP8oZJ/3GAKLFEQw0jxQetnRC7rj9m
slSjwNnyp6KahV70CqS8avJ3submb8rQVkiRIb55IlG/Jj7rYu1IZxR0dtHE55Wg
xA+0B258SnaqKpEAtjs9TVWNZrBKz5pzMdm1+bwRFnP18QFksr02Jc/UgY+ZGCfI
nV1l1dnFOHGGSG8ff+Pn1Kp77MyzDdlTv0W51PP7NCJZv6Ko+EzwfIOqa4XIXhKv
GymJsrKLNBW6b1Re4cyrl1zpHmI722ml1Xr2V8d7Fslrtp/ayBB+h+3GDQYv1w+9
TxNQHSeu3RKef6ifqFCXZ15u9pR85ApVVZoiTk/kZ0dD0WMy0ub/HTNl8hdqieJq
dQOu87kaAnP8BXT+57CqIQycGCMuD05ws5B9utw7eZ9o6YLZ6wRHG8iFglDir6mF
YZONFK3hCnh2YgwaV9HuTiaiidWURUv72n/144lHA+zDEJGdlstUAMrRcIKxJNuw
r4YPcaZv2nAg3pAKWx7OnLKaW6Do5n9J+8JjNYXk4YaWqc9arSyIGTNQ9Wc5C7KZ
YyeUbRZKR1R4mrE8HV4ByBODZ4amTfQvSrHztGxsUung/8ShYScMGDcATXnTGbF4
h19HG9Kj5My6bEvnJDpeegrhLD9ERwjdN2aJ2lxxRQm28GsePtbOdndj6S+V5BXa
dFRTa6p6bTXwpZ1Ozcbxu/UeT3oNPwZ6ijxIBIC+pVziuYmnYSVxiOaDEXiFAnWG
Oz01XzgoQKU3uoGm5IfzZ7OM9QBX7jj6pI6435gBX8TiAM5mVzlAoQDoYpt00kxp
7YKCOJFUMoyteQmmsxc0lGd9WrbplSAjlhaYjXBLaH4b39owluRF7C+ZgYRKjfdH
7yvqRJ21BvYWrIXpgoJhLI6T3Nc0es+qXiJlPfJxqJLtAPzsVJ6zi29hAYeVqWJH
Nlg7jDrK/fLhcmH5p67pt85ssEBSy4Lb+TY4CRGwMmaXXPsWnT5z40J5pFfDbUpw
R//J/Q4shmouRfXEjA/uvaUvm3/9afOVwBrK4j6g59eS79VGEhOhuHyVtzYnyeFn
DFm4/Ja2W0QpR5LCei4up5XtB4MJu2sLKiCVfbaWqJE4ua2Qw+JnQPsgWmEkPiib
BUlvbUiG/bcLkxDgVsdpIXWW984Y6EjwM+RDAJIsXd+tJh6867rrNeg9xcp2kyN8
IJgaXuakqwzHNkZSO3pZuTGzpsNPr7RD92gNVNCnxv8KcvwFG6GKwd0t36JM+L01
h9aRvyCz42JF6kmQf1e5p1e3HmURERhuZ0RwVecECs6wgD8+w3ZRJwoYQaD8aVUo
5KfvOn4bDHXqDkiFMyexfT+fxvSkuC05T8fQYIQhTxBDp9xpG9Nq965hTrC41b0f
rSv3HFF/u9r8MndYZFr3MvXw9hvl3C+ct+vadm3oUnryt6NP3dwlSeV5b1frcRN9
/qrTBd0vaYfvKj3BT9crLGlsQS6JKrOGbO5WJkGCqJUKHurh2qVhk+PgTv4op/fT
4MveKA4Y/haRTe4fFkFpHx0PlSKVwgpU+qt3cg67AtWR7kAgdncBal2yWFKAcsBL
iJMlwHKn2bTaxbB3hvceg8WNNiCrBpGa8eaOYG0ssUPxMgimlT2V5OcR+0gegihs
8ghVtaD4ZntGLx+4ugUvJZDpTEGsoJHk++3GHEB5N2UK4M25xUVUccGopNsRZWi3
g6L3RYm9dZ94ayUGXKH11pCpnuzBC3D3TSCnCiblp9ScBVfprP4HS0EXtIw4Qv2J
XbDgTsxs7aNQ84f4sYsIhHR+YNWUdGN57yC4BvI70E7CAL4nE/6AUob/c4527VAU
AfFoLSWNQdbBwwAEcbOIkf+8oDFTXwtIc8MAtq4m9uMlpWTl5kVXleRBx9W0/PTB
7Zn4IVrEPwyPFHnpVzfZ5Dp9l7I/DDK2PJLi0pr9H1QF2E5Rgfd5McpCpHYAIXbp
zfKqQmIceg/RrLcJmQLiC8ZxIALtlTl2HX5jsqBUwSUmNoW+4fvGsN1gSZYGM7J8
HJTaSH0fh28uhDHHZq/YSItkYdP+kYX7tSFmtwJkoA5/lffLjHruV6A9pE32FXSO
4DVqNnHpIp9Q1Yuu0iR4lDixJMd1I21yX8XiyG7/J5X6eaoVozYmGkIW87VV23QV
ZsOiLfhuF5ZXR1QTyZOJcVy/9VgtVQ2po7IDznD6DqU874kgbB/uGO2eq8jmjtCn
bvcr36goOP40jYxk//KrXHp9xhSPA+qbiV6ozpfQuIpBWItCpYyUoM4JwYXzpsOC
DfYcHySv3CkoVtqRV+9SgB5P3DNAOo0QIWAIIyGmN0Y/MolI+JKLz8XqCp/KnjAw
ODcv56+SO801o0IJRoWFLwezbjompL0oIRaOvspyKx8sXUpMrTspRry9071tbRX1
yrI3YuPb9hPlkoWvSDLVWnWcmwee0qOU7BlqX+TTD1IcOi3tSZXaZRSZsZ2mYiIF
f3U9uhzgwlWac7SildqRhd7Z0X9b1VtLIpD8zujn3F+G6AenD4mM4+zzboHEEoeb
JDNVi+cIORFeITWOi/PCfK7sXUBvoj7KYb0FviqiI0OPBVRn0yIOIyDCM2WaW1rZ
wgP6QVGCwAATE4NzUizyEMECP9oAoxjHe5LV9q0LAn3ruxJ1xjmMlJAmwSwKoSBh
C/K+OItT6mbPPsesmzrcnV3IKjIqjvkAOZuwqkCj+Za75AhHKw9iDaAx5xL/eCD0
oabybUOq8ad6D+hj1ZTUN6ld0Ss5Pgcmx0QUltjaba/iDEwH12nkn8v1ylk1Fqi3
/0Q5SjdgB6ykCpuiy92V+3CG+VqLYBkhAaeBkTYUGENKEMQF+pO9y6CePjfs06cP
Y+upZtNUwbBj51HZ/WzhgiU2ROX1AUyVcetRYrXu1yAiMAv2qZWAzPT0vs+HGMNw
KyNdblknb4GyVy5giXEKHs0sArT4cTXmWyTxUoGEGUurNu2U+Bmb6FdwTO8rJOCN
FOqXNAzEVjz0u2wkQdSlFwi4oWRFLv5fYZqRHUYXwj/dr4AImRFS06O6nK5ldQnD
MS6kBVyCp5K0F2YSXGyJXojEW9TTLiyCm8V/L7Ev/Koka4nJ7v12B3J9zSqN5jup
Fn5YeYS7iiemeMMkygHpQ04uAjEN9S2U+azQJIR5gl88I2iQDKRWJicLP2c9Iww2
rXXPnlkAy1GR60/rUdidGfpqtSWRuTvYVt76TEZpOushHYoa/cAlnLGNzJZgW51E
6aPcVaPUgfPOOve7jsVaCdlVmVZQI9EmTzv8n6gq/JBWt6h5Pd6QlmWLadn4OmEh
nxCmfyz12d4EvqFAnyqM92Fg3ruho0JmswS+eA+BQOY999wPOgXbGabY01UQFGZ2
Jj8jcwyjVu3gFAPOUJ7mqvGiRQQbeTlhDJD5itSpCvCU0q/s8myCA2lQPwM2XfLg
iuNnM0oeqBafNolU+FUD6DTwuDiqP8R1ejJ17vZS8ohvTn3OTOuen4n5LOYWzm+R
xhMVcgYPTAw/mGUaFdDMqo8gBL9ptfiSMXbD4vpS/6/BSh4IsQJaP8Ak/a0kjvBc
B2Ao89ZyMoVNwcCNKJCxio3Ae84E/U57j76jSc9Nankw2Kv9stLwmCq0e6GK93o3
emaBbEdrky5Itl4mHl45ci0kaqkbV+CYvUp2+RhW6Lxb7b268zyzqaPnDQwkEA0r
/WtbA9t1vozOjdxE+FAwqOE6rE4Yl1faWP9t93CxqoiqG5RyDHtUTSFQR6QqRgaE
Yg8IucLcyV0GCZP1zWZas+PXAc6UJwgif815uSfjprFqTqDRdu8CyNcm8xgChiq3
RYkwmKHBL7dqgw8o8QcUiVz/fH4+WZhradK1R6rzLAHBoZkVNQcjgrmVc5RdNDw7
RJNSoTjU9j/uI8q7E4mdFcPDuk7qmkMA3WbS+Kf9iNQPnOFY3NaNfklOfrwnHLqk
Ssen1t6CBgk/4htbRQprklZsGqKiIGHan4sBT9GnHG7Tdjf6y3QGbM0h5M+r3Qgh
BYL4drOJ2FvIK3gQBPkIbLXSktD2CRoxoP2GQNdQVslt/E+1FrCTN3AuDFdOMlv7
tW8Ib7zzskpY+3PYMrzgfaN8hZHneMzJW4RLc5COdQZO93n8Zlg9tEZlnJQofE86
oULINfLWL4vOw9OcZSHwRMw+tN0pJoOQO4a1T/CLVJnPgITt0q+84jRsNBp/65Ce
Tcxr8K/fMV7+ZKbU7m2yU5mV3VdAhkHo8kYtPPp8ULYbWUCf8HnoxpqjDNKVz7nm
y+Jbt8DL9Z/YJoU46M76FF8NFHwilgBO5QCW83Na5fxRyBosKB75TDOELK5XsKvc
veHH0cjlVKmFUNYEXCn+s5ghoBFX6Jwyo3x158MFsFvxCmubqFoOxHIgv5wht+r9
3YlsjET0x3iS7oSQnaD8PWUfn9qxgwzzptDZSIGxZltAtLHlJTATjw+f1wqsFlUf
lvxTEIpmfRgkKnTXj3Dn4SeZ1gYjehsoe9g1krhXlh9Qkoko3bWQRsJGhf4DETxr
jkboC4wyU8I/Pj10JvPsynqssw9XSDCqbJXjWtUHv0UPSDtPM8yzV0PyrMzPesjs
qpurSudoM8I1rmT0xnzhIJfbAKzJN7A5xxG2gnkZY0AgyRPp+XSuVkata6qpWaPw
CE333MOyE7yzTsSpUks9FGMkOMzIarZ4DtgM4dvdoqyE3vPc2KseNzvdSSd/oKNs
ydUyPbYvBAQqTwd4oEwP2d4jFZUQe7ZEpqQEYILyJ+d2Guuod65HoFQEkw6BpPEF
dHAK5Li7dHF/AxgtOw8iDqNM4ITtXrtZ0qc7LZ2Cj5tR9fiPxe9G/91OPJA7pmop
y7CPZnvSqkXodHIAbfIjTp24cDbXMxJn6duKe1qy5b9pnDJ+FVgfzeXo7xgZhKME
ja358ejJsoxA3ngqWRLRx3/AeK6GsCuX8ZRSxvGqrA+BpiiUeg6srmLv/WqX5mys
NqfFmeF+7jvNPnIJM/dmCnfRKsyzV7AXPeXfLMUDuoJeWnnaAgfJOKGayGKGLvip
nr1a47lVrQFnDKDHZYDDCrPTAJcHFu3kp2jkgMGIuzvCoRKOau4teU3fZATF6Fjg
qr40/DAC+L/Tg3iZQBwVRv3gfVQR/HOq2nR30gYkLsIHcAtDrlQSV6FXgq29BUQ4
cmp0NoYnL3yXcwrLVjuQNGRVgc10QRdE7SC0qo9B/qnQGd17kJYTwZDZH/4qvutf
EbWz763CFJwnpOxShUM4S+q7EXsVWHN65O7w20NySrEvwAscHZzdXLNZJbqSZqH3
mT1SVYM+Hk0FSt7wAwDreOhen15FQCzrEJU4yjv3WerfLQQURjYVkpd1gztJpwow
oKi4xgP4j67GdhbYoK+xXUUM/HA4AqyNtUghGhdn2LvrAvh5P8LTsxuLVAlql4bl
9yId4AQvIf8PR9oz0OLLGCwqRp89Gw8iTZSVAnnQQ+upiUNFYwgzcox5RhDKbIls
JqrrijMmxxcdi1/mOosfW07w1RfrA+pd8GMcJU8W5vtZWL+tz5UFPIMgz7y9Rh19
kTQT5ReqvHlkaxb7mofF0EzJpFU5cp6SJXcySV5ZkY5V+IrbmHMTOyvR/tZQJksI
1Sb/D0a9Mq7T6NL9ISGeb8IpDQk23GxTQopWS+06KXm0FHAVc4nn1LtJATQEBwZ+
cuUtoIT0aEfdosl1PjAIVxhVptg4CrdC9+NigM2NDltc/a3i21AwwXUuK1ouk/wv
7DG02Hd2A6R2ZaAxy0Nx6wCCZ2poOL1zza70eUt0mzqaQTrQDrQocXu7F3/XkX9G
KIuBKRblIDhd610b1NvCDMr/S1QBinIYJXpFKfrM7KuBj8Ua+QK64f9EZ0Z3rswV
7UIchYneOy3CmcTPCI01xzmUyz3hVsKjDqmgptXyNFTkqBIb7AiYy8Px7m/Fx2Lk
dVDXPVtcI6CHMlNQ7khb0XGYySzjmH8TjXuZZwocfLF33tJeHV5ZkKLsj7Ic9YMq
fMQbvvjsTnE5y7mPzZwe2lC/s58llKunc02tiGdoGq1GXgVFNX/FXIWGIK2nt/oj
sRC/8pyB4hDVPE2EconY8If/X7IuBjFImulweJb5zlTRyWa8Zgkv+SXE6gIg2vao
SE+KR1ZaboBfpBV9LUKEEfmeAnntpS1DjVvDvGPb+bzI7hJ5zhEV/fngB5tgAc4U
FFTypCsiqNqU5dysvefOgCwD0RNmSE66PMmbMfMuUYEn0Cr8893tzgNG6E+KBwwj
fVFzp9hl57xqTmJeGbbcZJE/Qr7U7oJuTPi+cP+eqMm6kFqYoq2lx6j4iBrXop9M
YP7+3EGLAvwX0bcivUgRsP3oohs9XYmYDqaBBtZH1uKdH82RuZbEzCRyQY7IeL6z
G4tAVQzUqvP7tVPS8c7pgyxmoSGbTJXwT2lYmO7z16cDRo1IWXc9iRGw7scbGU6b
r3pD0MLWVrvPqb2RmE8IUt1uwtmt2Tjftr3vBEs2/IgggVibEbqa4cmompKN2nPI
qSEXmjkRYAjwt/EvI01QS5oo4x4dqpFSli5aJjjMpgCckwTK68jr12a9nInz7vnd
/glvMOFE3sk0GowRwjQ+fXD+g4HGCKG2Llh0k5swNioWERuINdj1cfxv6sfalKwb
a2bofsI7atvvtXefBbfyJhTs6kHBkt+MezaxNCsRvEcytqbQA2w5ul3na2OGHzOC
chhgq/GwNqPZnkCCpI3K+PwPEJo5NIeq0eHdM7Ptv9bmt3yriwQNOUzbdkUgmFix
MO7j5zir4Q27haewtLgt0YrrBGAb5W4Q+4/Lu/4HXs4zp/Nx38BfXJaRQABMAZCu
fEyfhTVyVJt27mT9ol8d2c4Q6CeO+oofe2H/R9VPY2PPAZt4e3CLNmNHZlXbsmgw
qdYcOQVx4m7caWrgZJY5i8IM0kTkC8OPoFnRdCkg3Ct7FXO7VKZLcDIOj07sPUZs
Og0idD01dbVVeeBTpzfzfDhWT8OlKYq33cTg0s4nD/+ZcfGaCJHGr7J70vKXWcUh
Hs1673sDjG0JnJ6carUZZZHLfJLyxEF6zDJZ5Y5s0Nm4ZTN46F/GkuCKWD46d/MS
b/2hjkw78s3EofOXQ3T7D7Bq9rblI/DDvoIAYVESNwND3DotV8G7jlCcv4VmFY7B
H05mS7Vdy1TfaF7ke1ZKpg09Sd34f0nsVEB42JJDdp3xnJ/918tk4CduJ4Wwjleq
Ka+LNWH7NwTKEl49yDas2sXn34ciwvnDY4kFmNaxwVWoQ416wkii5cTaZU62jK4a
mZXZgBZdAllgjSVp3RdfNVa16/PSr3f6V8BSTukhYTxBbgIkv3ryctuZdg2yP8Z2
9NuCRpKsQogGP7I60D/zLDYfXazauip9im2uL8OqfVNn3JewFkDsvk22tOJhwY8P
mO13N3XOEQNBxCgTvQydvEQeFPS7TP1lrgl08nBgjaaAPa1McT2ahLvTtpBkej6F
6ZCKZneSUSwmhb4g4WtlXCAUs5udXW9HpFTUi0pa5JLhb/goaJc564+aqJkBx/ne
JMhftaAuPNYKU5ib7NaXuw2lfcRMWjZMGZWUzj6G1xWGfhN0xiWS6162WNkT+Yck
PnAP32gBonhnGoaGqgkDPF1rWksg33Z78mIW4m68BoLgsuH1voBPZMckRmbVeYpq
c40kKuFTHxcOQquw7V1T7VFyeAauDoDhyP4Ax6XlV9coBvOwkyuwDTmcL4dk891j
qf9NKLcV88RD6cfGcFFpJ1jrG64bCtQ1EpoA4jQu6MVnw2INtin41eRkcbEqZAEV
5Z1VV4abzd0Tothh4BxaVonrFedWQmDZE/h4EFKGKSUKnejtXhOpJtD4JzYuf1nn
rW3UYSzkZH6l3uoSL56QobSuYjalk1gUiIHwj8Xw2tYoFkR9sCvU3YbxEqAYXskX
EjBXG6z+IhXtXRYs+ZD2BMcp7lvN4wUCGlfFdL8tQXOIcEr9dP0zaiCKCNHDixk3
viGIkhHtZqfyqJXccEIsM7cC/AIc54QaDX1/3NN92or+jxsQ5tnATVxR/vyOVkuE
kvDDXlTCDjq6RvEvPYdzEohS59a4zHtGbE1hrRATAiLmNwJHl472szssxhk1n/rn
yo5+ljM2fiZ+vSyHDzHY9ZdS4Bgk3ngrj/GRR/waC9IQdRl7av48Ww4NFwZI6PKJ
wHK9SaSdArwzqOSvw+MglOo4jSRYqJ1MUSmQSwc3Qvn/ucBCADt1fTE2Ho0YJQUQ
ryOa/vHSaLSamyd2OvJcwl4EKXmgiuU3douWRjSfzaMeMH4O3Z0BeXkR/96HhMW9
B8pm5MWhDVOT3PQ6pRpsdA5CAuDIYkp2fTY7a136+aGNmxn5mYkvm/7VKaJMLYLe
N61AHgsseg49IxZvX91H1O4Zq+QxbatNjj/bmls/1TGrNIE9boAYs2oMUlGw7Yha
ggeortb1UBmCAN2vqdhgdbLarKd5JnLYocLWspZpfU8mQ19SYWWW4I/ER5WxAKR8
bs11Mvr/4CGOp3kvKlEScLw3U2Xov/zfQIBRwxQoz722xYLzfZz6LdTdPfFsdPpO
zElXosxP2KsCl+UwR0sE3fA4DexUijNNFpQhDjr8nezSA/QSmU5y+2pbb65b1PL6
f5H8miBvgO1VBgsgmFF7cP2a6fnKg1phvplf/UNpI5pQ9WQeUe5Ncn8BB++obZCS
bq/D7X0oGBR3yacM5F7AjSm2/yVhYfiUmOw1IV4QIaoj/EogpY6GinSrJCygDlBB
SrE4xsIJWVZzxorJs8IihcXFN8nYYxFgffha0RHAL21uzWqelCNeOYtRQ825p4rR
nru8KB6DkmJ8oZIzX3XrxuvzyWElygM4XBWt+9yblj4tJgURc0UtDpn9uqjUEKUD
NFKha+zLRlV0btrgSVhDvr47/SwOZbw8Ar1QgTFXJ3C2LUmLL4g5YYE1X7yd20kf
LSAF4WRsvAhuoUYQsMBJRg5yz1WXriNUVUyN8yT0EfSYAt6Wa8jQ1GhwFZE2Vghb
dejgQ7xQsnA5zK29gdZFu++rkg/UebrklgeV+/ZJ0B81dFhSLKavpvHUKdtjjF81
i1HLq8j0BE4WsL2c7gqEq49b70ATvxcUNA+BWYmLpSQVGvd2RHCDBNbp7BolMSiF
XTaE6emPXSqP24NflIHPKnrsFygSdj779vrw4F4wIm99R5RP66JYmK3zeuMUZ9pE
QWY+YUT8LbrPdJqi2E3OLNPbYI8O4LJdnusBJC6QBunNVHoaFnNcktZDY4OfSv4x
rMWQaJu/vn23pT8OFYY5jZaM26+75DBpgdD8OrrxfKM99tGwRi0grmASFxATaWKo
7yoEXiDp8a1tm2XgwRMKKcM8ojsvcyrdFfZpr9y3HSbLlEtvLIX3USmAbhRLj8OF
cwiav1n9k8EUEzJ9IvDo+IsMddfn24qSYKo21UD39ipMGAVQwlc0nHHZBZ0HGc27
BFy2F9uADb0+ZjZFJxtfHhR/VmBdOhTHoPPE9x7+5UnVL+/7VKrxJHZiuzA42ALZ
IyCY/qaA+EdhWKCqlly3EJvbXDwhf+0k2Y+R7u9CDCv8KzaWC/t75YBveUHegK2e
CiPur1Nx9HU1iUuey0TDkhgMZAfC1eo4/1Dphh06rmB9PK1dOzcvvJK8BusTJaCn
99Dq7x3Xd4RH9qkkiyVBqWAFaJYxBs/R8MncH5zVESWHZ4pFxIsc9GQ+dT3QyMLA
zOT6n2svrYYM7Y+yPU0hWeh/1SAULaRDFmzMIYzcKRRW/XeXIyNUJKU8Kb4bRV8E
oORhOMQ5Nj3z6VZO++6fQd04ZAov6VYhedBQrwT9G5B1TB9yWjjTIGMzDYdTlVaJ
LTdAB5vw/2ULcp/rtJGqqiVw8k8wGclYQXXRLQg+eNBgukXgxz3VfbFPBtnQ+3IR
82xaj6lQFwyA0ZtumjBUkk7Xo4k4777cSiuQCLucdoeQlWKMNxqJiKZgcKpJlF5+
1jHW+8wq2UFzEzS2OgwwinfsVZbVPiLzIe8lrCC9PmNQmrdaNHYh1+4FKllH82c3
k5bQTx8MqBTNfAm3+clNx2fBeqKDz6As6MG/aJFdpNMvSLP1hYPuSFohpXIuo4q/
Hf4jsVF2ueMaqELYg+n+xKkne9ZLyRg4M2pq7TfsBQCXLHTVzJPJ0+JhCRn0Mz2J
9yg4peZm/TuKNkwFKZOgr+Q/CTCqnfLIOqUBKnNUAiKqMwCEPpxOD25XRAEe/E9d
cPlE98pafV049xNC7ghn4rYAe3kZV3qKOgCRpOyF6CZxZkjJBoBqfopHR37BXijc
6Pyu9B6nQEFJ29LbPB/05v67nZ7ElRljC23X+G9PVV8c6ieEZsl/90T1DTQ32dJC
xgI2EQ9/rFY/siI0mctrua7JoQ/or7OmJCp30VkW0L38XMHk3zcNtvnu9U73WWAH
9ntw1yQ8rkg1vLXvgxmcvfKkRG+by+wyqII8KMvyTN348W4B4yan+LQOl3ijB2Hn
IwcV2gYyJXu1Ic2UQBArSHJOrJ7N5tUcXQQW+nsUMOm6ovqwzB9KscxjVo1xWx/I
nmFFDqOl81ishJsTrcNgiOvRL//laqZkC7GBADUC5rRpQJ07rk5QukuoPu28mzsL
/IpxXtilkLPufnKDbo+0NaUQ9trVle12JrqK0NjTWuVGmzb9/cLkQPLn3c1bM8Bu
xopAg23S0PkCayZ3Lajoj9RqCudkroizX7F1kRmTaTOWsq0CSi1K2fulsAovVYYb
DM4PwnGDIM14Nb8lt2mqso2y/EsIq57SHCL5epEPd0a0yJwR8LAZMtSW5vuEyZdx
NKOuI+yXyP55LJyVXe0FExzRxP25nuBsImlqSJ3VfdqTyyEPjl81aKldgLbwU2lg
IPq7SXk7R9jHEguYIrQxQ7l/ebMLyogoXC474zSYgmHp1nvY7e1h9FBvxkHRlhQe
eJQl03fQADbtmVCPfwaZgOIUWoVKXWu0TDQZXe65/xy8Qx6MC90Sbu/uKzNeN7jw
NXfqx4K17on5zQp3OiZRG0fDkqsQbuWe46XLPV1IdVzZcuOmUBuP/Kxe9kNRcPa0
VsPjJW8+aQ7pft7fuI8U/42tfJJ6GT0QFFBGNxEaBcXRbL5e9mYvTwlEwyczDFQ1
osF+nexjsPfEkyLCc+I1xJET9IFEX5jyE7POVvRCo2eziN1W0FhH+wdomQt/ggt6
TzAWmVGFzz9XsvS+VDhO0FCvN0HysmeHHCgw75YFXT+/gcMoGKsg4ObnSO70IYza
/2DlpF1oGgYBh60tmhneXh/fqhaWF0P6QwgQhWFnND0h/4sCUUagZY1f7AEpFFaC
oAbnao80Og73aAvU2NO+gx9fALtYFhk510HsOIhJ36cC60V4PSaWVqVOx1VoifFc
W+Z/riWEgnJ/3Nous6JRu6mAw1lLLLBUHlmovUD8m7O1o+bPXzehoR1fP7LIUNP5
N7o/Xv/x1hCU7J+sG0DoUoH7KrFoQpw9taJ7KHtHqsiTZW3IAVnojHsfUWCpgHu7
vw/Tmi+qIW5TJB+tXmW8/skAgKP+j/tiMMDKXh4Wk4i+kCCI9uhSc7k45QRH0LtB
ttCQqelKlK+df46Yp02J6PGkt3bCKCUv2mIAQ63hqs6MS7spKi8ct5+B5foSV+hJ
dok3XdyFeRYUn07Vq0TQvz7Cr9bZSmbFLoGkvwfHPpm3G4jftPyS8COGcwqhGiSE
dkp1FJs3lrV3+49NRIFTe7mjaf7w6FvZOKhxvPojgNBB60OK7CBqzzHGxFsCzRia
4BMbdxa/cWuNwDOJ2627kaEav1m5XXdw3mj4O0TRcmxPpwNvuBT80inDxaahHsyH
W4jcLDtwF/64uvUrpP/5vSut9Tu77L3Oe8GGwQvY6B566v4WrklCdwSyMpStNFS+
jn9VcVQt0MNSpJsQdqmBTQBpAF/TE88e+oV+jqDkoiPZ+42jgHUr0oBlnSvdc15W
c2Xep1L/OHBmrFigm3VEofUD6qrZf9/kDE+z8h5knSN5y44RLdg6BHJnjgxprJ8w
OaH8SIZLOy48N3MQoPIT+wkhOC8IJRx2VpYd+mOtAcnL4k0eW1wom3h55i+PNVhZ
oX+T0q2gDbqIbyJ1FmWt/oviWHwXbU0dEDT0mlPUvHcGBR0Skse0w56rJew4C756
sNuluOHP7Frv+vRTTCA7j15Uk2xfUnQzOL4DXQB/xLggTCXKPcw+5vgKzt8XekmX
QpqhJ7fG3bmDlOCXt/mAGwnolvK1CFayTzv87pFe2fZ9lwUV5u6o1UjUIpJEcxOw
0otlYudyqy4BjECiJd+FTRuIUSI1QCc+0XY3QM+s2w5q2BOqsMuo2tkofZoPGy6p
snkuazvLDwkfd7iPA3fyRq5+ESDmDb48BnfRc1mdtZmCYdzs1iNsRvf8xOWaB2aA
a8C9WVtOd+TNWpo8dU0z6SniRQeURneH4PbwrByG/Lhy1mA1uBdtZf5awee9Uc9Y
WHLKJILEvyqyt89HDTcRvQTC4CGIL7mEFb20NZ45/eF54isuHEGPR0x9hfAVa01r
ZpqJCiMl7Rl1KKnIYD48/aVkPu5Y3Z5XdHKkBeE1zDBvm9UZXgKeMIfaA87rEkRt
g3KPAgIcmFIdrKt+2Np9T4EqykwfdeX6OZ/2lDBjPNr8QKSQgnY7t+GdAvu5VMQ6
dBBXBdjPpxcpdIhOlotCmL/jEDHCVRxIG1K+3rObkF8cyVa7PCgxl3G8MFpDVNaS
Q9cInATilIcXQ8Husz04OQuGL8kUtT3XyRz08VXKpK9HMYuwxI5btnVGrsU/crZ0
r62HYK9OQTShf06L6PeqXilx7mgJcJVfT3IlbYnCpHZDn5DGPEDQq3rlD2Bbhk1Z
GdaIuKIPSLBLMkcS6A27QyxM7DVQW55yTksbvq3Dm1gyBFnl8mZ6tCEzM2jol/Zr
J1cv8nUhtFJ6wrSbexMuNJgmxqfWcwkOHuIii71j14ViSDl+7KsbDAW1lyXQN8SG
5RZqC8jIjqvsZBFp+3KGa9nPum/C27UbfT017ucWOu3KWvej2SU1x+xfogiuEg5K
8M0DHPGkKedMb0+co/xpx6EdeEEUtIpQvVkNqqR6P935C7A62qIDnQpSYJserrLa
+L3ywopjlPl6CX0H126iDp/DJ6VcFr0jNP2mdkE33fxZ1L4QX4xlmgvaiTm9wJL6
a4u8TfhvES9DPQ6BTMRwAKVBV6l0gqK+FwHl4T6HCZ3VJzLswJMx4l33Ln6eQlR9
UFiw4dDW08euINswl97/CBHDxlxwwCKNPxOAeC+1vpEYASyCwB708xSdrLFyy4rB
RUEwW+gG7wMO2MFD+JKJzbY8ASD5n3TvtgBK+K33DlgNGz0U4ynUBRq4Mj9EKwxP
Ekb3priTHC0BkMMDRkzuBGmVilNwSrBUT0WhIF3x5dlbLfMhN4SyoPM6bLIgZIWE
lv9dVS3b6/VDhw+obWsmUi6oNSY/O4b1XMlqdZAXQ+pcV8RVOIN6oE7YhpFYvvi+
akH81zP0HQzFkfluu1yfam0rvYuD9CEuKZ45WLl3bv3Rru2xRq2DZkP1lFPxb2vt
Dm8EwCDYPqd9ixQLV0QJufTvK/cpnnrYYpXlQDfj1mhXmRiBS3uflxrjuUaghSQ0
hmH2Y2Jk0iu+h+uiRUvrvDbNzlwDpUZgulkipAXBhcm5yh37Idtcnry1lJzTyqzw
1GplskPH97aank802cQDpSUofzInebspVyRW3mTQ6NqkJvrW1c/fKI0/s7OMaAHk
j8pMeuDpHMWfuYGyeW62gQDpq4ciGU3j0TMYQFhMwXf6rcIVLBgkE9EkjEqsJ471
WZh+jTsU8VohThK2QzfjUD/AxOf5GCXCIJqZ2e7hCVAVBMlGxPc/LgHThgZM1usW
xW/z9cOfx59y1whAnImk/5TX+FRR0B0dYh5lTuoIen5TLCCV676lDGGR4O+NPcMW
qSxTJgUHTtiktcX5BA97LYAMJQEKxZ9ve56OXPJECu3KKBqORHBoeUZ6ezMsXnl9
B5KpeHvIvxkBn2HaStOP0k0j5dqOjCe91+Lx3K+y+eyBcfEzOwBCE+TjPHkN0SCQ
U8d4N4qBzvIk2lf+VZ9PcEtVYOWVojN+0Zb4v6sdDE5l7Mp2UnVepZkfLLX55Yzp
M+CNw36g7en+GfxTTqEY1myT4heJUo9ckg4uTD6QbN6kH2CUv/VRGyUEroh8MYC8
+kgMOphJaetEtZvSEkZEAvjx4lWICnpnXivObA3zNiZ0wFz/OcOiJs38jafuQUxO
QnLbXLya6b/C8jQV/LrKSXmmYkCrdFlmqLO8dSbvT5lXRVo/i/O8hYnBStsObVc7
AtS/khrt4XyutQsNJhW/WcjuO48jpJKTa31Il5aBtEL3ngzho8Inn17EkzEFeEcn
xgNdKiHSFp9Hy6Ezfgs9Fp8wk/3kbe/muiJuJqpboy0H6TkQ/VCnGJzkmwZdNov4
xJLlwoXgbDo40fI/bRcuA5fxNVv3rUaWvFM78u/p+01ClrVI2e/sfs4ErfgxSbei
qF4LMwvx7TnIohVftv/bft2xci/9JzozRrGVWOkd2tCs0071Z05B6TkYGHBA7Unu
5kwXAjVE1XpMSzg6BKCutW+1hRGvl9YkpO2mC3d8DVFzNTjEYvKipiHJFKctpxEz
S75H/WSautgL83M/M/VNq7LIVtZ12wXymZ319TGoRoaRHw8yirke4rZjbDFmTdGI
wWVkAPpRpCj0fLxnZteEGY5pf7Fokq6xOYaG0rHiH9kgyGvGldTF9D1P+9uhPZZq
Jr9bSflWQHtHRSjc4sTbY3PXVBB+iNrMJOyK05wWA9aI5+JmlEPPsA3ZDonPicoT
LE1lMGxloybtbIPmxg5WHVbTq7xNyvC0x98LuCeR/ZWHoX2IUS2+ajfP1jSV1ILl
hc9CqHU/pVb+hALwJPwETxfuw5ibvSBmbdRYQ63k7+dHr9n7/bOcpdT0lkTYLEUP
lReBpUmr8jVrgCw7+WakQ2Bz1ciqtN9V6RgAGgPmpaOqab75Y6qPZZ5eyFY2a1g3
k8M5cwXaUVk+7rg1HWNU0SvbfAsu6Ez0ofilsAjc85g8us+BMdwoinJ9MfQV8lHf
iTDs2fjK44Bi/9mTANLHZSs0l0WjzqnQJUP0amT3qXFfWGTMj+mrBJLHXlGjDC39
epo6o8vBt9wMcKwB37fiTJoREqUsjYSsYFoznGswA7UEXgNy6gIcc5tuymueCHhv
NnIPGjTlMDsKstlc9h8xoBcFr6KYreEYvMGxiCWAw1Jx5cpyA2MsZfHA/WCriAQG
S1GQihjwh8wEAWnBqPCWnpI1kpLNG4xmdvGIoDZl7LOj0EGhCO6hvNzCmSAPGEn3
lBr22K93D9BokQt627Bt/T43vFVzSoctKkOnmyNdRcdu9DfpkqU56UD2TFaPGrIp
rs8fPY2b9j2PAYkpUc3Dh5tkHIs7uV04IqDK9rDJJnwFpvOSdMQiSrX6/Wqsa11G
Q/JLrYuQJKODRQNOZ4D5fPFxOb6+ft7tsCJcZt921GMWghVv3SI/swUQUZ4r2v88
79K+9f+fCs2KX+Q9oAlSBk2dlJSykwFcdQY7+oDO8i4IrgDDPRAVIABViE0yGseR
pj3+wN/8ZXDqaeAgUkwQMP2GV844AbZcq6MA+kK589/XcOrs8oeM1p2mNiV62v/D
zZe4Z2zFrEonvXIFxquQ1GI1/vkkrI89PScI4cxVkcD93bBySXAvM1HenWU0Z4Q7
Ys/jeUEzQRtHcMyHH6uYVrW+qZ1qjeAWV8Ls9TdYDVwrhDxubPCiRLoZqarXn/i8
GJLzDPczMd2V6IpAD+CTyq3Iop+4PyLEIlsA3eEJ00h5gr+EeLAkXm7w4PS+mlAA
2fbSWw4cOsIvdTy4XZPPLAb1BpQgfNTehw8Dvt7PDzcyWqXvk972SF7HSUB9LvW/
5BrtuAkFpes15C2xNEfhtpTYFJ4vfpvrFAgOm6ik9rXCVOCVqm7D+euz8dXuzEbz
autk0rya+29wWTk63ZhI4bF9bmwFbbv8BeQ493fsPUunsE8ym5mwaHZ5yzJ0nmN+
eYhYx+ARwOHRSaOjsYnPNwGXqWvNKHBKqEXPjRPD7LOxlNTPYwqe54yGLth07ZAI
5PlGJ2y27Y1rHsWkCPOyuXYtq2YGPHPdDjNNFUjhdvwnqIjLZP0MSIssEhR8VwKU
a8Gl+m97B0zqcApKBEdmuphZBVnNinD2CjiKRUeB/honSCmk4dyBTuguk66y7zUU
bjBadl3XC8CiQcCmlNIWSuHBl5M/oqRXm2ijVrAdPCOaOiHXvIOZLkGIforaxuzg
7+0tw3itFV3TpEEufIkO8WQ0E9eCA3nk/Sy1uKhMg+gpoCNVvkKPuuE6yJ38if1e
knfWhgMoXYb8iiEd3CYxyyFUDmLTjpk+vMA2dFoWG+F4hdYUwu3ZvZUodY+aiNuA
1feQjbXd9tY941tQ1iuz9EHwURKUTvQl0mHXb7vcwXVCYZgpTdK3T6Fhw+zQcPqh
S9wcW3JwZrGA55d7PqM0YJCogopvHwUihe+ZC6Y451ilSV3TiMIGAUbDMWdMUznk
8z7XnBqH0zxeUBS3nB0rTZOxkHkr0sQUgAFy9w9OEe/cWuDWEGtEIQFgqPGmBUfM
z6O4F9jmGyFe68zh9SIuOMYwMD0xUeI6MGANTPyIhGOR5D0T4Y9NjRKHtC81W1nq
J3Fhm06vNUHffo6DS0mv+81gTNTUmjFQiE0+GcqjJSYUVqY+q0gk0/sKy8/7zTgl
6elSfkv3bS7NdAA6WfTchp4C/cD9vIY5S+h81/58f3nN+NPpDe+nwOeSDdOqStXm
xw4tKg77QCVUwzjC4+967D26p8fB/kRyHwmyIwcAL30AA7sZEJBk5E9FZsj9+2rg
JvdhAhFOOkASmugQMU+OOJwbtQX0m+wjSrI9pUIEV3K/neWsHsNs3eEudCGKR37+
4C1YuK71XiKiWRYOjAm+V+aC7bk18mmFire5Yn+oQso8GFBjhE2JTfxQsm+z811z
vMycC0BYQUvwjYNdQQnE2SqylfrdKY8WxfoLtbqkdqm5pV9DU34hJcn9FQo4m5b4
q168QfFsZXbqE20pzc7YLaO8viNCxgjete3Y1hArKr8E0nBciZIaCGEYQ1bWX2Ft
TkNB859d71Ah5aMt1CJGwGOPTZyrNSJ5wkvrm2mkdbahO0XEarPAqePLhP3j+PP6
OqppG+34rEGV5n+0LcjSIiMT1z8DoWuuHT6jex3Wjbn3dKC61wkqfnyae44LObtO
X1q+GZBJaiAkkFOT4GJTleFLIr+a9CeIV1zcwXwmNEfkWB6yhj2HF9vBlMszycvV
gOoKarZGQDQuHA5+QOs6ml68ObOp132wkxDgXcszWeDH9DxnQXrV7Q+J1dEtJnwD
wYdH6ltbH6ISKHNU8djF/aj1gCk/OptBEgSgQpOfDOhwQKs/TnOS648Wi69D0qrA
o/GdImkyJjjYEUTXfcJwHJtlqjWWxf/o1tTpaz7xkhn18M/EanbHG6JR27Z6mihi
VETDu9igdKMiX6iBaAXIqehSmT+3RSmF1Ij1zSJhstEO8z1rEUcXWEyIHxh8i97Y
cvPANgj3JvyWI8SNjk09Dl9E5zHnLI5Zh9epwhReF0NNFyMCZ5brbzA4mYZpz89h
Cj8vdIBbjM1RGsSPLvWnS6CRVUbxLqK69CAB2EKTNWRa66DJD4uI1EuWG83kqCyo
TI9CuP9IAml1pdJXmpHdk9pY6DUa4dH6thLtMqTOiCRe9zhYd8uHtYuDuWV6Fghw
K1WOnRzVJG2mbvNVTpJhyhdrJfLrSR9g6M5zfA+dQD5f1He+vdI5P8V4NLe9H14M
YF79jJuH439WgybkdvLx8u/6xzbY0wuh10ixzAWtgCj2pXWun83JhOJVYEXlHsBs
fxuslAObMtTv9A/x8tHvR2vJXGRQRr8qNwH3r1j92A9Xb5tt0DqWhZ59Vzai1icy
bTKJaaDsmUkIqH8BTx0Vsf/DkViM5lq9hPywMHZlPYEagESzljtHCJKcGx11xTF0
ZB+aj5B+u9iKpzVe+NS1e4sp7jVaZSeUYkNIH6w0ILAmjwzFZBVv7zCdoV0IOwBJ
ywQetOVF9EPBkAWkvNusxIsI7GT/nsZKbQESfjP9TMLDyhy4em33SGZfG2LMo4v2
bJczm+h6x7Vq9d15mWoReGJb5cF+01SRUA5aHFkdlgNoxTeP/iQkgj1JuEUeeCdg
U32ijBvx1R+VHkncsRokmoUoRH+l6b1uZZEni+dv3EWQuwjO/Z3qHIqen80poeM0
sgWMPuUlDRIujXWZ4uNPLaThpoXekzMrN8nn64lgLqtM1S0ta+qO3bahr4ml+9zu
v8Wpa1VZcHJ250Q0fLOppBmyJ6r36dWogslzr9bmEs+zzh2V4YR4yk51EK1+3ue3
Gscp3oZqSJ2txIlXkWnXhgpS/ctXMPgVKdFUA4/cBsgKpzWwyNIs7F33cqYpFWgf
MdsuOfv1aecCwUWPHffkm2OaKbqux/Ue4i1KAInKgAJZGQcqbvNEs12203D3g18Z
eTAF2dyaPDft3g7ni25tN30TRhNheJ9h+cXOCxdTG8oOub1Z4thAOua9y6I69lue
Wmgvchzc/kJ6NMHdd5O5bgD69Oq+RH8OMb7oER8fzEcXmjM4gfTnwXw/oQ3Zvf5t
F1tUTh+iwjQ2lmphxpDfwzxrV2Iz7GVN3Gl1X0HjjMdczuOOyPA0feKYjo4FJXP4
BVf7+0+ubHuqtLUTNxod6gGwJRQWVk9MfAF3Hvs6YkSItNEHmR5g+B27sx13bDzI
hv1VJ+7aM/6QgUXUvxLbzYGl196q5pTtnN3ZdI+ziKPSOWmdc0v65MkPgrd6lSSP
PpxrpjN4d5ncbVRyhr/cM6fr1MWVVN8zC6gnPEPsVvcuZmoqQuFJs8IFL+8FZaW6
zB9+b7w3wb9emfXE3sARElR71gQWPYGnrS76meE1W+BP7dtu/JXrgoaKHBQxe7Ha
DOZZuWEQ/MTQSjDQQfdD7uYh0HjE/wEsBk2FUS26wHboXb5+QcCbOjN/BASBmGz6
VIm7Jd9Ju12cJ7xcMCj20VmQIuzab91EKHGw91C6mHeGjYFHjL0XmlnpmD0ja5v9
D78Nf2EsVuNXHRFzkf6Y5dwsFPqEPMOXIawjfmWHd/lx/El8FwCMQi0nXuaZZCFP
TIBLKZVQY9s+JTitSK/+rCciDw3iuV69nKCWtqV4Y1s6ymFp1Bs/W8Hk3MTocxLx
FAHsW07lSK9OpUVYhesXSWXXIC8hK46HUEnLTPpAiTS9n/YPX0lG/5VUDPze/fu7
wRxY9KLp6e7UxItlfTwoOB/5g/DPpvkMl8BGdmauMvk8wYZ9UJV0dUvz2g61ciUA
nsCpK3nVQuuEZoN/ZQC4AEFhsTWD9e19sSNIIGpXdyDZe6i2IqV1kjE5raIzkjpk
SRn0f4PNhabAaAwfsfl6iXXW3slmXzcFCEWDU23aFERGl6/r1z37mze8TJs8V78Q
7AOWPhu98oq3zl7iHmL0sgKJeU0SPGNoLPi66jibqDdGT8SXJYujuVOXX5fRl5mu
N+S9nhNROCtMDJIZgSM37ATTfJCHjP0LNgvrrU8dMW3PxxUpz8e9TgKZ8199qGHo
5jEjBSAsyMUc7CsfcA3yFg2V7J6i+A5xwS15Y1AgKdVnxmW2u2usyM/N/C4++7/K
U1U64vBD/9d5+6y1LGU0CnfYsMyYLVq7au1O0vfn+XnxxCliKv+QL6q5cW4ctby2
ykaP7gkDg+C6h81LAmciyvpO7yPOCudi1GWHpXZ00zYHusv4d/muoFg23cstPmGI
KGRLkdav65Bc7nQkDEuMZgahMpGTsC0LZL8QuJx+nyRL5rh8piDvYt3WLDqiP3We
JjePWwoTQXceSG1hwHAW+Q+3sfjobNa323+wmRzlzKo/27Vn4sbWhveVmXiEungJ
pLLJFRQPDwtIoS3x2RJyrCdxonuBvw0g1PFceBfWMBkxj7QrC/YIj+YVt0lB0UyL
iQ2UYtVTDaQcA3v9AEx67DNBS7uJV33ebDvC0cNroK1OUyDeb0qKt5v6q8kJMvLl
DrOvKDVHlCmBMk2DlkuhgVIXCdnO1q+eTkF1GuAOrHMaSgCSE0vIsWDR1dqx3HYc
S7I2RAMYi4CrzOQYresQHo0drRXe4jxcN6AFVdfYyAYKJwewYc48UU16scw4/LSf
sw7RgdTyzXAbC4++ptk/7rlCgUHo9hh6jkenuPV7dyKz4NQREmZbF4aubj8wCy5j
0qOZ3aYy9cgzflnaOO1HhmVGLs7kmR/yYcic3YknZ5OGEkETeXVRSU1YtqcGcf0N
G8i4+lBp/5ePWownYJGLDlJdOyObQyLQCRuASNv/HGXPXAaNvCvdVhjTqFxIjEGX
XvHspRA6zlfacCdMXZ2XG6YVK7nGGyEtHTDN/n3GmV/YEKTVtdJmiW+YIDJDfiO0
uN9H9q1xyHFPfLLTuyHbLKfJtD33nbhvOL6cqOHuW16AvDaf6ayhh4u7pq4rOERc
gsDKCjfNxxyF7RFEuw/kJNc+D7PPTzVO7Ts95bqx2HErlh8LmItttWiQBjRGxsns
u0GD0r5+s/VBSK0bS7hrEk18SMkog+saqIKPvivJiPSnIuOPwVBIG1wZEjWAhMxL
c2qsl/IN1dWPgNjSU5e+FRnT1z9H3sACoFV93tW1JqSLwJkEccvE+PXyMnetNpGN
30vYcdBw+mdpA4dmtEviLgdq/CidS4MEGCBK+M6BEcBgLUyjL7Ed5w4QI/qNyJiH
Qk5rqq2hE0OD8I6uJ7w/wWDOzPpmIrszWdyT7GLSNB8+MbI46cSNYRhUs+GO5ljD
yBFfbwekDuLotmuLiCVRbQ+IU/gTcXsBA15V/8lu2ji9J++SjTnbruOHh1IiDuNU
bswPFbZvOEUa+QLW3jZBnyZRNj6QDPgO3fryiu95+VBR/oRhQhNpASaD+0UDPaA3
2oupt43JTZW3Jvdes9b6IZ14sOPshDERC4IokygK0x/JcVx9bpc/iX4U5Au0hdll
7vN/apJXHICclU9KMpCubOdXiXoZPAdDFQI1XHdcUeWfKLI/QHzwzGTeXMFj7Szp
PpxnIZVXXktfj81mgNOdlXfrUUNlLJwMZ2OvzBFVqbsMQzm9cxmoYDK7WIxZBgoy
eR+YvksIPMwnWTsBLWNmS05B8sgs7lrIo1rrtIH2Fev/s4w+MZrJyWaY66wHD+Ys
nXdD2YFxisDC0Xd7R1C8Tg1ewhA4FWYsgWigP1S2boHft3js05vMD+GR6kudIOSi
/6kZh7NG1o/6eckctlzBjLAmqErWAIfdz/LRjS1GKQNCl2RM4AEsYnugGa9QIMUY
w3rHGxKO3rE2AXzzcIcLIhm6XpeF4q/4wai+KBAbVxEU7DhuNJoSqCvCGAFOT9cF
4aZiMKid1hnUjPe/jTDuTM50fz2vXLbOZLmAGImNGn8C46WlyoOcfztok9J/b1zx
kCPFShUHxj8P9zF/bSvu5YaEBx5kCItAPGqXcApkCEcs3Po4+BnpT58qPTEqlz6z
XcmCNZLHwIb5pIIn+285IxHIo6j63MSFLaiaYfNgP/1ufzn7PM79FIyxxQfRP3OF
f7zIcEM8ywtVaTkAbnomiTAxcoFTCu7brkaslS1CAwPE+nh0MNxRP/Zpga8bV4EO
CI7vpXZ72HPz/E8xXk5lRWMlU2zWh4PL79ozvTer0Zr6/tfIV+/U6vqviqhDWRy0
jDupTv5AR//QSFUXoVHjDGlPK4pwfkDUK75j/zsoPc9N3Rms12HvyEIzY+quEqqr
SyD9Ya4XpTdqx2tOz7JVcZjxfc16WkQkfrAY52WhCLxGvx2SmlJrDut+lN3PC8jG
iEi8FmNU8SB3Uxs9R8L94Mfd9piHF12OSdm3hPU2UiQl1Qj9QIHN9FKqeV5h33VB
fVQg2w7bSg2okU+JOSWfXsF9WtbWuXylH/G/1+k6XL2s1wS7lOQ706YgAbaj4LLH
lpmAgO2iCn0O+t6ePTxVlr3W285m01E6a2APk/WNeDuQdvMocK9ELv9UHwmL91wX
B5prNflhQj7UsWGgR8LS9HfLaQk3w933y1b+MQnqDzJfiiRoA2zVsCcL0nOkzTu5
4w82eTx3MRP2p1mTbU95u3Un15KUsIvzqfwnYN5hjSQ9/6x1d5S0jY5GzSMhnU/O
6uefC9bkx60zrj0HCw8Cmx+91BFEfujvBCYxnVkSWbxKHTPHXBj5qbkim18NfFS7
UXbeqBj0Yv+TB7eEFWXt00y81dCKG0eKSMujEiIS8bp39LiKZVRmQshICx+v+gOw
o8cd+7AHxwFz1YIDespl1hAQEZzzQAHYLzgaFwi8tnc4unxYi4oBndoP2tnkJwJw
zVsslqUZ6XZRHRjTU5TpzGHoDr9cc0Munz+4SPBC1eF38pSZV8Fsz00VS+VuFwd1
5oFwluLJUHfgIfcrWnSMXK/jW6Fe0CQ4c4m5sB6G5zG5LD5EfSrmPq+caRi1IDEg
TgEiylkjJY0L9wcja/W+8iv4yOf+tudMD7jfc+AJzeRsuKV0HHHZ5DULZA9AIT07
5oG6IwwSh21CLl0rPBhFcLBatSqAl/BGdMbgHBFb1+NvRLCPi9/JcfYAVcmLt5kJ
6h6zQsE8H//EJ6yScVsnbKCrrmQ7GelLkLzw18OMjzBc+v19teu8olAIVunVgAqU
wmB4kpnUuFtS4A7WQrMB+hwc6T5VlYJsecwAWr/3/bnoC7dfTEcbJMr48p6b5vSs
YDy/SY8qijYiV3hZnH3n1aVPTk5AZIwM4Ip9VPT7i8l7DoZFK6FhmaBEJC1L96x7
olqGCcSpu7lriknzVmpTs+SQngRxpQHiVranzfzeOK0aTDXDGZ7Q+QgYu9bNU6zE
DvCeJ+F2Vwr2rkfvtGy3Thde225LU9nai/tSXgtT9qaK+HmNjup38IqT5uTob6I5
8mTPnefKB2OiH1VqQwj5oKRnqNWIW+ndl9WQ2vL/8wHbUFzpEwHrq4YTHcH09cjF
F04s7QG/zgDkdGeGNdFBvvpzpPGdza4g7wMWAnPqfkw6C3TVM3CEP3+cw9YnNJY2
Grc0LLk0o+WQXNwmGXwJUl19sVbxMAj/iaqVEENKnjFXr+Ve9bCdTclwXfBfvLcW
94rPiIesd0yRUxMUJ7Jahugw6REHH7rjxmza5Li3B3FMzbagazwqrqXs2xKOpyou
2NiWPcoPM70sCFue0irIOkOshxjmfXskcAK8MUytzZShrUu0F8p7H1x5i3tuUtVF
DpFP+6RfvQ/vNswIkAr6WU8K8lMryzxvycPgNCGu1GARbx/nR+qXm9K6fodvfvVZ
mTGOKUFKyV2n17rrbtPK1Rc6DepfZ31bN/apL8FjTUSgy1UHVyTwPiGoH/Krx9rB
/NzYshhHF1Bss0/jt5IyD5NhFslk3G72b+9Gdf8zhr4XGFaqPYyeB66W7pNgRI63
778Pd+JpOdWOp7T5FrRBo3Hce3YNSC0zI31c370b42KeitkTXsaIw6OL4v/lea+t
R46ey9C6Jkav9TCyooQzo9pTH6rZEq063AXxJyMWpGAwGGzkBCKEdmnO+5wDg9OT
f1+RfQgNF7JL7vngKDjPQcm6nmiJKpEsH9gIMjZk3/ZjadsG4h7mmoq9hGzC75Mw
lg9oWXd99LX4MeI17WplH/guvEquk3LBDwwrYOxcEwQR62ivL3744FNHjvg5jBmL
Poq/ud3ULk4+tc5bwfph4D2ZK/kL/iZXevPUbSUoWHovB20v2jK7EB9ggBXv+ilI
TuEh/T51Zvi3+4R/RUV4ew22b4qhHmVBNe07dWI20qL4xd13NUvZ6KIwNkardb4J
05ZgDVShpISplgQIK0pfJ6T3zj8e5u8EPwl8Us6+LyP0ZA5HU7eSXnH/pPIdmUZv
PIzU5H8spl1BeRlnA1UIrp0lLiekOu1J2UjwdcdLqNqR7pDpjIrO/Ryx7CepPQIU
vU3bv3D92degpM7mEdR3WNkcC6Hc/msmVAdQEJkIFo7FkwPfFtKf0/Gi+5Mm7tyC
WE8vD5RMsEIpR03UbBn1jZjZorlc8Hx9STyW3xCPYG4EAS1jPX9EPFWJceuVgER+
vLGpf9fEwSBF5TGBnIxmn+ZXrUXFW9wh3wTd8y7IDyNGGzunLJ2JfinxhqGf9yxw
XIw3FanWJ5dwwIuRMFLB2qgC6m8vgl62/qBfjhh6ggOJM3o4OHhrKHeB9hzSZbqw
jNF0bIUSUboNkPmaF2P6A1BqG4iLW7/3SD8IgJnCj6zuL3SeVVnOH9IbEtbMoQEl
GFqDOhc4ps2k/o6KDIS0mhSmKhHEcvxtepY191z7qmujKRQI5mOYOynyDpiKo3TM
Ss0GaaYmm3/uIdTy3ex+xztJlYSE8Cpl9akWSVHUl9AZBX6+kftggJmoQa2vW1S/
X6TZ7EmPqhVawIVi/wELuC8LquSGXpqj7c1IOWM4+Xac+kRJcyBH6UzrhsEx3GoJ
LgjCyEoFamM/AVO1quWRjZKeYY0WJBWa+ErV6selcgXirJVfhlLbR2V/f/3GXydA
Uj8bFXyM6YT62H3vH2WL1IMYmpWl+zGc5wcnreZnyu+5jViRgqAenEVLcGGbeUe3
kWRdfNSl8V1QVpFow0AAM7sBgEBQFqzaXulaQ2ow2Qy/1fL3xLLHfrijn+Ptln2h
ReYUymjSQJnRFqTyq65bSO7se3XWhOABGrSaIhvdADKFNlqs7OhOwPtcuL+G5I4X
+ie52eFrZAloeJuWQIrS5LQUIxMq0JFpl7Mxso1aLi31k9TiIAyzbhvDBSSm7oBZ
A+SfqGeTe0Vz00ZZ9YhgOLnkrEGuS1BTPJzXrQXfPx8ZwDjhpJXvF0w9QknQnMtW
ihqowEx3/3+TLVhgAWHEcrCVdg2+4ymvy2Y1w8RaTJUd0nQWjKTTbO7pi9iCBROQ
dPtarhDhW0J2qs1Ay0xS18SWbn4ujwAygA1NOKgWUJ7Z2hb47l2Uqifp266IqPY9
3MLKct3ijAfs35+6zMT8J1bQu3RsHa8qZNKc8IDJen4Wto9mul+qAcXfgQK7mWqx
NG8yCjjGh3sx44owjz3SzzYS7fwCuJmeGnpJB6l5EAc/sUIBvb18j03RG54ETtm2
Fl1UELPuJjIlVFfgPKzsol5OVkSytKLqMzRcSdeteIZOyXpTFD1J1ePMNOQTW/16
BxlsY6iEO7fCNfRFRdopTr1LMHyO/dJnZKscInDCMXNURSv6lH6A2g0k7KmydlGc
fxBmk7FiyL7PjNCJTMPIrJZRd1K7w2eSqwvhZuiTElUHOnUywVr+41Bl2xlLEfLp
f5jUrFGvwKNCe9LvJrbSzi5cQiLrwM6pN33fUUKdboBbnhf9WOucwOhrkNEOpDDz
un4AuD6StITtllFMYDC1grSmM7zSzcPixLpCQqy/846MZ0zsFArUymtaz5c78qyi
fUG11dLwCte6EW3S4gNBCinU6/mC7z7EoU8pXr5cGp0DnQ0+4y51YmFw/6RhR5TJ
xgFuPpZYST6vyJg4k2vuFHm6sHU/lXbi2m/1jWHWdcA8Zc2K6/IJooPBFHGdvJcx
E50w20/jAqLlU64SRdFdWG43J0C2kO0UzdjmGnysb6Ww53Zu49pSrpQ3jmSiMO9J
6VBf0n8duQV7qMcdLqb0L/VlsFKql2af8myUws1MRH5IA1wU3DT1PqhVydNgqloe
qn47bVcSI+O4vg0K32BxXcRWMHNn61SQCu4kiArjuIZZzlX0M2rtQFp37cGQ23vP
b9bM0mdWwM/uR1LOhrO1TRUZwoKRBW0jfkr5dDivP98utUpPAYF17ykMxZ3/3HUA
eTvakhJeoGTrAiWc1zgrneOO3kKpEiIEKYAPaSA/oubfybv4STG040einhANBMJS
vH6XJARYhfiDAaCgKB9BLz1P+JtZDmAbZ3Q5gBTx5tkPSv6xnUGTAXJTkSHoHIqh
yZaIDUpCn0acs0CajBq64rTzc6BaOtsJMhzkuWorRYRAf3ldkRXPEMN1xCbuQL4Y
LyPj3wpKlYANrFyTFGWCgHXnbgN8ZFfHPIrF9izDEk3OH5y+LXsqPCrfrAKYp8yf
NmkGGi+tiYIFmWOsv8UtJGIPGk27EsZZnESZyZ5efpAkJ3VUHjV3J5MVa4x/SpkG
peaC1mnIJCnMqAjQbGjrkH7bGQREVXLt6veNNPaJgprfBHv+uPyDqmpYgnDDmBlj
xxD5yZ96WWIau7qkTWLLCiiqaMWHFRDaytBRx8xyVMV20aMuB7z0TGZF4ft/0AOb
+nJk/OK00ErqNcgRuBAF28KX7m15ZLKKn37RPdQhH3n80N1l46f+e7Qxydpxdt8j
hR4/d72dqePfHwaYMhdErB7GegDISRPuWM6PIxITidtd0NWB723rQQn/RjiQTsfE
BYvbZusMs45jXt6+TZwAARAwd+26r/ndx+ZZAsz3+F4cLEzpvtEJLhUU8vcOD1cO
mjyAnrwhuufkRkvpBMv2yyrTRca6p0AfJz7AqLSbN2yjcACKPdxbDYnvW+rmY+4g
Vw8cIHOudb1kZLPs6hShxaWPvgg/8apFFZFaoNycwExe38g7OOCf66Y4oE5blkOl
2rwk7TOfh3gXb0Grtc2JGF3UbkKn4PsqEHcc6Cin2Xk+B7yd02paNEyOpau5AJXf
xMjWPBHB5LGX11IsIoJcgiCb6AS773eT+NbCtsbIfrA0ESCqGGoMXaGfSHx2O2g9
2W1QaXlJoaJhB5Um97BCLkF3SWjCIuE3bVFcbVBlemdJH3ebVQ4cF5DHK8z4bXuk
3G+OsGz9Tzz2kC1xEf4rd1+q+8+s6KPYU2evGYgbQDd+Z2BMNDJ17Mv92+MnAnv3
dY8ZN/90Fdg1Kr1tHLTIOpHcFzH/Xk9VOKqOmkS0kCSXSIwIWLPujvHkewWzAYm0
VdRW2Z8/TNoyRgkvSp4xTzLg05YmQq9x/jmhXAyGF6q8x7HJJNzxBjte0VmbQig6
AzFh/hCEQ8eMUxD1T/dWDUBm/dw7zEfgdqT/U6DWdktFQC3v189/nQFHpIPB8LI4
JyZg7cs7a2uzsc7VDWdQ4aLajxvv7/b+fwn+7eqIgxj/1gZqzj9OSyv6JkShQ0OI
ZKoENprwz3O5jq4VBZHJROl5qkp46kg2k51WucyRX7jWODLmBKt4bypVrIO+wolg
eMeSDxrU9CnlmtBoE2jWaVvBQibeNB+GMNzxfMZ5j7L6WLCVnDjVnqOWagb0yjN1
8/OEgQfDQE2t6AYOG0LuZAwZHlKJDIY7FPjOGRYioIhNzCNBxKwKalN6FJe223IM
guu24AbnAsrbB0qJdObaYaKMjZkbxjo3AveWi9I0RplVSAVfya5hUZ9E07aOmufT
kMM0933CAV7+by3uHcH/zfTSRQ4TYwRisfDGfUzjQWyCxSXttDUHNbDL8PTy14uO
h8rAAb9X47IDzb/syM0IQVpp6a9wSIozCysvhqRfhTumQ8WUaXNlQgrV74KEHuNF
rx1pNgW+1Wt9TklOT2qeq7vVEKRzNl6+O3wZckqvMFAzCgu6dDIBhOQxFDG/9NO0
M0Y7PZfDWd0119kiHQZvVu2Hypah+g0NpN9Q2u04kvgeXhN1wnICpcwwgwbtnHux
jD6fOa+KfinGOlMSA8cZ6jkCQ5pG5NNtRmcqmQblN3nmD/tv3pgPLktsSOeuYImT
7nygHKLQIaFfJu06I93vM/bfDOI3xaHuJzMXCZdQjSmYoJgEoqqz3jA+6sjmMePR
ItWrDx+XpDOHAbPs0anGz4kuLap8WP4QN3tILX2GXTxkR/0jH8Dt12QglNCKG9Su
lZUlsqMh/e8c5H9UMsbazenw2kcJO5wm0G2Htif0I3UxEYq7ZADNFq28Xb1IsCRC
Q8P6mc2S/ynEpMWpggJPOgEXQFZtIqEdBEVMOYMJ4qbV0LQPSzDtqRnKXdcWM6J9
JcPmCLwNtXQARsuYAViKlAlk0GlYJrIEtIS5iyWTP+Q1c+82X0B4XEjVczYnjXfZ
QjTrE3wF9lc4uCu8KVH87+c1gqhOmlpLHwTjrGRT8ySKd7GWYG7ZC6Z2Qbxv2FYl
LcujadA7yhqjUp+WjBfBxPO8Gv5Wuari5vA70itBWm2opfoGVdguUiwp92QE/ZKa
Q6pn9cNGfR2FaXCckXB0TMRDeAKvjJ594GaFWri2Yczl4PwhhZbXccxXIpyx2Hrh
6XIRPWcjFUw3bz0weYij/xmmvz3JCPXBOikIgSP03rLU+pzoU27vhX98ltcEH8Ae
N7c5bRdIJZL7UAJU1R32PIB5sf136niq9Lk98Bk7SZA0knO0978KCa0YWqJHys2d
cxA7zoThlo6r1gds+V+YjqXizKvbu7gaU60ZE3L9ZufaGNsE9xZOLVJ7tcFoybjj
FRYKa7iTXFtLIzA9VPuhwq0wzjr5fWSg0iA78gLc/QhFDFsXXi6p0bzq42Zekp7D
LpK7YVj24v2vlgnlwz4XRU2x74evRsIuNGttreuOy18jC9MkAfNBoP+2A1xwWtbF
SwEBltJ+8YkqkzSeUtawhpitZ3so0XpAJ2obQShSK7Atm+jCeuu9BRHrCnp+/VLf
7nmkXjOSRG8b2Sfv/Q2GrI/PA4FdKateXEzSxBvpzFs8mqz9y/jEN/nGWRfCS0+P
UPwKGWIupnCRIUJD8ZhwJLvEtf2fEp1D0C2P+lJnCAtm3UBMPzRp5D6WHIycFB9F
dDisBx0mPy23FPrXMPIm2ezjgU8j2Pvi+Z02o/OlUP9IhKqiOYQbGwBkD/j2H+Ev
YvIZBd+PO1jgsFzJ2TNIIJMzQP0C/+ZWxQbSDqDLgAbD91dh/zzcIeBNerxXKGra
X2gHKYP2xMda7nZ7hfHkfw44W8hgcpdq7fceGq0c4ShCWZJ/RMxLcGquUibOkPIQ
vJi67rn+GtUk/RaaY8tOXjbJvhMKulLLSn9munZA+e8YjxcWn0Jr2p9LL/o8PkfN
F+uR0Lo07mDH+Vgovl6n69Fhj+kxsOCNLLuF2FfKe8sve9Fity/8jRS5YEgV6Y4n
PrjyJ6hI+uLIbNneDbdHTaPpypzI7fN9V9q+KGrPnGN6AByebfR9mFEu6foUOJ2P
RP4sz6lEjoQqkMFdlfYZ9JQPrVx8uTX2XHqhTMzi9SLj87JBuLz2eaeZvNK3ncHJ
gMfLYQ+ZrREvXQSXTqsPklaUMuMqljhVFHnX0sCsIcaRIRBz6Exlqs0ittCoecYA
atoMwLq7LfM5O65a1JkFC44Pg8CBeSOrgtIfZ+r6m3/8QVWZZ6crSsrqm1CsDYGF
WULVpP6t4IPsR4K76/fpKvHNhaR+6CnuicDVqztn+ETSuCdJsO4ruLJIKTBpPfzf
NaZuLbt7w5fJwaWOSYUyP0xZ8Zp6ZNUwrXluIX3TvVYfRaDuq80SsD1qAmLhKjqh
up/3jHnPjvQ5QpS0E99XeMYzO4JAsMoqZ2DWOpD+gvuvVacaMtAKGbtTZviXwTJd
CHEAg30j65rA8w/4fhR/uXLaXiF+zylLWaTHWw7gv40gsPxkGG0L1EZu4bnaRwdd
M1/lYPLMbfT0Fa+cXjOEILI+eoHGxYjUt5t7c0KOSuSkuk0ddT4GUg1Mc7/tEoBO
F8sT9eUeQ0q6o2zAZSJmE2wUdrj+CEhs2pjbvh+fmF4s1hO+YoO7NxYlB1+s9XTb
Wm+LRBCFEXw+rUX3w+51MrHxlF7RONzIMdmsi2PNMa7FElCJ3X7PgfVbeRxgZtTL
/cDHoHdie009LbkfvJlHwB3WXDnbuqtOOXBK/D1psrQONSDwZnk+ojg3TRsTw9Kz
OusEh3wxv+lEbIxaKuXD8esaiMc+xGA8qb0XEBgC5C7PwU//GIW82QCdnihK+O+9
+r9kxKUeWMxlNLgtci3olqwa7S6+3s6H7/gcMuwWo/PUVzVo1Q8m8Rb8gB+8kMmh
0XarusnqaiGGvtHlYDFc5G4N1QbvZN9Jp05npy35lc9g85kTaPFuK4owMHejOP+j
R1wCXi5ElHUa6BpNdeYEEQbAEkB4Rc7cu3AWGUr7xkc8k9CAh1YxrNT/0Ol+ng6B
6zMzU4nWqo3crEjMPRFP9hI3hQN/kwHsoD7f7UZUEeWE7vPXtuz02KjuuudrI/Qa
UtyiRPssOW/HCIrqk6oJquu147rB4VTb8k/9+7RE3srCYeCxqywFQlM/aVO6Zlfw
C2y79MmtZyk7bsGueSanU9xvEs7t5OAGFnO2cFbMS0wxx+NnjLzyq4WvIdDOe+SG
iIez7ne1t7nljuyDcV8iBQyUTihD2ff+9mOWaI1x0ZGbEcInRK/05fMRu+cQseJd
bPWScbiMWCrS7gjVe+BJ/3vjH1k4uR2YAcVmaCI55b/nBz1gX6ijo0kKHb/uYKCW
Xh1pKl8xOOXze6UbFz6y/7AkDocwQ4xYb7zbfD8txeAyB69fZ73btV2rzbH6l1xF
kQ7J1/LOmPnS7vGbkZxNTwzLmTtiQqwMvG3v1kMODPJm/wHTx7V0ly6l9SElrgJO
U1sg96gWlYbAdo2ZaecYTOrBkPcadEZnacqUxVsjDbYEafdU2GB4iV/IOZDUDt0I
od9ZskJc5tkb3covl/dudcENsEIcBEF/jo02zFvZTfJyOrZgnmsDac3t1tAxmxLf
nfte8Zwy6QiQnewc6Lh2jxSTszN7B/CDyiVn3c4Qv/6NdeFvSsY44MA/DtmGyAQ6
SbWCzXdE8sL45kjnXnDCJblAgXiVrwVsDGAjT6B3PMqPPPbK1UgSCzl4c51soMk7
cn+ptKRUb8x0KNctv2amnfX+AuK0/4knh07jAFtrbYdipKwNvv/OEYfmCyOGInZb
qS5iwTk6D/Q9mY4yOGWEx0z0Q89mKg0ETZL3WV0TfZJ6HcHC2xNRCTxkZhlMt8YK
knyPoEStwXp4rg1PgFw5FiMYuBMwIDfQ9K8bawrOlVQoC1+74mTtmgze2r1PS8dv
jKmEZ5j+BPfhIFqMf6DPkbDookNtWXitJJT3s1cKRemu8Jk/FzF3DOxJRmTbnEP/
Dlb62iWwlt3NZPPagBnBMTkmF2NYa6uueNb05R2lcu2tLnsmcsfKslgbMc03Nlz8
sFE08SNNWHrtsYh26rJ0FdUcQ+Fs73H6+cyZTB9X8mp9U3WiseYidDBk4Nz4TMCe
zxuqwJjt2zXiAkKwECr1FCq7Uwy0DHpJZ7tBpij63VpUgXQriScWgHHDS00Asq1j
vDj96GknUfZEtl5iXP/Xwj9CbqYwv7ddYJO/Gd2a0VfohFbjzfm+thSJCy6+j5Iv
vTclGOcRJGxKMENiH8kCDlQiBFKJC79msKcVnjo/vMDibb2mjbH1zQknZQGhNMSd
8jihVy+jbXuXdRPO3NO6jLP2cybpJREHQxNy4HenlxsXGS0rWVFOReL+KIOXG1NW
+k47XIapfhZhz+9f96A9XI6Ww+nL5grEHsn3t1CSKQVRNUS1aaMXw8jIC2+Z7/5J
Sw4w9hN0+9qAkZPOdbXUUCXab22xNL/EL1y9RQ+L/0Xe05O6Ps82e34AVQqo1/Uk
uGgskM2qx4yqsGyNx1pmU8hTd0v4av3KUjAV60KLZ+FJNj4BpWNGluD9PbuKLAIJ
7DX+323V6XRzD1amLq51q3zbVTB40ZfMzWaDxBXeTl0repAaKRLkCgJVdJjtRNQX
rwrgpy7Pm8s2ARCIx0c0QiwHhUAgaVNGhVNK7wWeOHA8EkJqV2Pgx0OmjTycamov
sgXydyYMt2vl13QJyPwLlCzLXFkr1ObsRu90+OhrUjG3nGS9v8xN8/lravptBBho
YAHVqVuaMAQ5zugzbOpGTZUXFgVnGeiNHUfLv9XAaPLmxOaxxXBfs4rlziMwzxH1
ZgHALcd9WYCG1NDN2JrUOZkXjNQ5+HQbDHFqzaM5tWZ5mz1Cw/8Sl+spRwh/5ND+
7eOgNQ6xqUN9i1xB16TRyN9MceoelIvr1SCCORNNLdGb4wWRZmFEEmW4PQuIEG2m
legXjNBTvKAp0SLjPpUqFvOytnP7kwSJZ+vSqaW01irujslqd8I1IR8naJdLXfMJ
U8m1BIkl47w22EU7vWQsuoHdydMyfjQd+ZfdEu14znXHGe6U6C4D5Qxl1RbRG1I9
KYhmH/Kl+kYtOX7p/Dugs8sEKwl/pRUY+fS+en+tzFMMwQdCoZLtO08+36KqgVxK
iIY9q3ripapjKPRKZlTvd9bJI2ElzG2EhHblWVspGyCGy2OHQaDGI9e9pRX5PAxp
y+SYW+jut1FaWD+3gDSgBbkP8RnGZYx++IybkZwIGzlLxBZpb87viuYwzz6inRMI
GlXVIEfNB87AopFlt04IfUx1IKzE5Fjz1aI+XqsyqbDQZcgtO5BwEXGmMGPSMMXS
9BZtn1lmx3iBzceUz+CtgY4G6ohXrWs2LzSPeYuN7uJccaa0LV5RaYU/NFJcNk/8
z9AOSrmj3adZWdN3igjuJe7AO/iLp+l4bsoVPEhHUEhVHLM9AQ24HaVdL1z86YKz
uwcIuLNHIF7E2HE2yYGP55FJKIx1nxxicG2lKsrhgIFyiYlPWXy31xrJojghlraY
Yn0/Vgqm7TmGKodDFrOcxSMBuowZvoURWTfJapuTUNK0ukBejORkdlzKK98cPdGI
Hyq0zZOHGcz4owStvwrUGSXSUIvXUhQeT6QpYAItMmy+JGZUT1yDoAhD6DVU+VuZ
YOifTjNyrD63AhcSF96zGNBjWe5smBSWTykhKcOx6iwGuo+CMoufDRqP6L5uRKmc
Y+gDbgP9llx3fondnP1sPCp3gafzLbFB1IRBPnpiaigtNumRTH5M6uZUeIojVJp9
g+ZRYP4ZxdF2sC9kJOtxjIwDXsLKGg6RnAul2yApI3yA8fqWw8VkvJi9Ovhf0bcA
R3KoaQ9zbTFoHcB2zJS9KiF6lsm/Gp6k4AJhWhDSHOPNQVIAwLmWOhxd0THVEn7I
one/30W9IgtiDx3Mr6j8iMOm6e/tRO1oGdQODrZbMKDNpA5RZ83jucfqLaqi75Oq
w0NdaEY6RPL3cRC1bcfECqDZKUumoRrJ5rx2PW3Ih8fxbqxYVJN3VBnE+p48UXWN
8os9ZBYl28wuyjImiJpYuKqnNC0ewPsWhmSkBqVLZbK+nicjWtz+ICFOuLfeW2Vi
TsuW2QZs0EzBzAqYfHlD7VqpiyAuOf+/465v6P1CsvfOHmlMy5sEai9K2d3GAYVt
GcoZV7wxt3xIWALAfKiPl6SL2lmgFPllwxe9SCMhrjTjkgbnvhmlKlzfxRYhWqxK
oQnwQZtMlqCmoO+Umcoo7Xr61ZCkW598FUd8cpmKCOaV9+e+JBsme0o51cTDuLKD
oVoi1q0SuvDue7DQq6Gue0LyDg2mPbpgTMsxBJ8M/OmLyoXqGjVv+JsFJD4bpX0N
fghyfRaIcJxILjuDDVMs/LKV7hPSQxGSM7sw4cebkKYiSCFDGrqjEKRCNuzDXQir
RvqWkhM9NcuTQVnYMXZGGTM4Xh6bn+suVMCpy+qfjT6fMOQ5/MbEyFTcJN6tUd7+
gSdwsvVHzruK9ZYmi138p8TAwc1uir/sQt5nISP3FYGrb+SMMAwaEp+HeMid2P3+
9k3J4amR4vePp82AbnPbVQOMbqb6qZvjRjlnPL+mI+JHLpgiLlgItzMLQRYIYzY1
c2fJLmKISzPjAc17yP7wgmBtVGnJZZjPCKMh2/i/DfJYFy5mNc8ep2fGvDTTGpLR
qx9+9c1WXKsILepC4Aivm1p5MbPA4l6UqGzvgEiEPHY4qYHbHhJCYieyBmmjTLyq
GYwrDDBf8kwrzFoR9U05qRxCmSTAYJGB60cUe2TeqfMl0AEWHqu98hWUtN14LoYe
/MAMKtZCdDlAT4zKVYSj3dA9mx0cwMyqECt+OGJUWMokJZUTQ18AjmmDnrSZe812
rpbOUezUqzCqvRB7lS2ChTG/H4Veau/6aBzpI8aPWXOOwMddaLo1rRdsfgWehpG6
SCGb3M4sTd9RTeBj0yaY9zCNt3xkWSoAZjIN2jf65Kt7AgyaFaW4pSbrKfCUZVUk
I5d6ILnwxnhgE6bJhmr55y1NnsZjY854L9Sa/0SUFaikzRC/l42s28LhaL4QUOSQ
9bEioDXe2BAr1YTGmNw/n8gHFQgy3fizsJAarbbLQGilNet/yrDs0cHt8eZ5rv7D
tFGdo4XE4U1T9WmglMyHrSNXFpMPHMIZKtxGtNtw35FJWdHti7awsdKrs95KXGNq
L6/LP12XrT4+kC4T/qIgXlIkicnv+hi2gUz67XuldYaNHnz9rNy3E2rrYLQ1mXFB
IuRT1Bh71KCm5TNf1FpBvGvwgVI5fI6uhCj1ShZIKCcMAA68hJ8h4KujjHmFEPUR
8FFHjvlfNk+EZk+JjVW9oGUbsusvVlo6a9KH/bTUA8ZqHq6JA4+T1DCjc83OsKDz
Adh3JpIzD6ZOurkk4KmoaR3P/dT265ids/OhtbV918ET8lF16dTdITNKtR3R/VLS
NK52vDxw2O/IJ5mUE9sk9XZsNKQuwUGy8qcj5kZJoFbFmefAJzH0SgkNI6BJ3PzI
WzlL24e3aJBKiCpqBKfO8AvXzcMnOUaMjwTLjCqOfsmytaNRvTHZ2BaLp7Ml6e33
WuFWnaHJ8+kwjzNsZrd0OyVrhmTqZQlEq805Kco8NA/9SIXN87wwzS9FYlDl3Xtl
1tVyktsJ4bHMPPMrUzYQfRMaOypfzlqpN4AD5ydU2Qt4v4rLzxzxdIq4ij9DYdrb
BM7d8Mshg80y2LEUvRe5ArH3kYv7pq64JfYQetltct8SFe6IHIP71+z6AdaRNToA
1rQgWz53s9lrxb7SmviKGhuCfGzgfmhpUyJd892RKzBVVAVbgv4J4HIYQZK8hEOA
Phe3iloGjOO5vCCNAajhuWo7kOb/3X1IRN16vHcrV/KvcirENgTu1durphyM2MEW
NmSpRS0vzwjy9MDc/SlNKvGqVovGIaNuaV9mHy2kiSfFi/u30K1GiOSlBgSt3m0+
zZOvbxOyKIINjBEp50/mBfBSQ0qJWj7wkpboEuFAJN4wlFFuVjv2WtlzCqt2lJwO
QXCs5cWofi1ioVf/IN20WRWX1z83mLuqjA2pVfGjjSsnPK9VUCG6WcVgGUY7Czl/
qHX3ClxpyqpEVHSJG7r3AzyScdKNPBwYZMJQ+PomogMKGs8VeqJb+PKqIEgXe2rA
OhGHx2NnPofEZTlupQD2eE8KfH540uQZC+BkA4wx2ka4FYkdexJBjUCWZNUnb87t
+7uAqlnCZ9U2l/PvPNsqil7mSNT9VCXZvpCxbYPy/FSRJSO6g+sWumHKl77vNLea
fwM0NsHf6Gppz60F9rLrtoxskMLONp0Fq+r+lyBBPO5ZC6whaxljqB8nM7evRLKr
pIragekQFMC3EQN/Q6uPU8Hg1n6ehsN7PuckvnXqUf3IFN0xtP3u3lVbNbbfG49Y
zyCCz7QgJ/X6WfStFXQozu8isa75uuZMqVt99aOF8Jrf34Pv3wa3/v4HEOelxUX9
OHk3+imLNTML3vcxfxsPPfYySAUFt9cfp63jgFssG0KE1ilys0QwpZKxM1aCU/7G
tA+M0RjEX6ZMrOGQZ3S1uGSSgWqEDXyk5WJwPZIPqFioCNhcsU2PVe8OBJTmG6Ht
KQUL1yxwthlcRP4yOgb12kOYQmjwxlBzoCl+OEWJKtoT/PAEOWHD9xHvBHc7sQet
/396lDsVNL+4D6j+pYogNz4W8Pj0lowhxafsbWXT6ECmcmC1qDH9EbAn9NbnCbLa
51RQ6qMYbByHUwEfQau8BpJEYWg8e2KyQH8fY7xk5WGv/tc4dFQO3PsNlH20k22x
Uw/22XvhkTgEq0czvFr7Xsa/OEvMaawL7qSWeLwXAjo4+/k4GKu8UgvcIKDrh45f
c2lVFnvvM/WewQAW2zskqdK+e4cyzq/3qPG3Bd0tuKvY/FuSGh1f1peQ4IHV1yPI
SYMfDJ/beYTJz9czrt0GySxmMtMsxsC9n2x5eyMiVstPAeRlYMHVvekdQe7DK2Au
tX4ImbCr5Ut5d6xRYn7rA/eA2SivXsipvYpQMTiRKdGTYA8O/M15QXr1UlX35gz7
1ffSZ2abkLrjSUpxaUoDAiwhZ1a5UF85w9I2uGz8NIwHdiEVI9hdN3Js9Xt9g7rn
Xe1Zd3rDgbNOGw1kY0W3cc5FikPyy3lJ1FMb4G07K7xvjtwI8u9Qf6knD5yKjYmd
ddTCJIW3E6KBIGYSTULhUVsC+9yqOVEgEqMGgtpzHFG8/bcM8MAD9cmlrhD8XN0a
3LiCEpfiGQdCcJrkoLfKQJrib3sBvbDGaXYvV3ixEoPnNJ+1cuwPS9i6JpKtW1Gu
Yws/Qsi/v/9sH9zp7qOlXtS45YiMv5+QXR87ziUloM5D6zpgNteTboIQSMMFC++L
hDKe194wato1P4pRkZ5ts5L5jZNR9/lTCFr+G+Cs8hdAkKfB6Ibd0/CO+QGrZRf8
nte8EpOBTaGGoY0fJRDLT1D4YLOO/1E1DTcjFph9ha4p9hDoQuNljTpYvgPOR6un
b5YQcLTiCkF6rxzKD+5mTzplNuRATZkUDN65ao+aU25Ras46tEr4aD3DQgeH7aVQ
DA9ShLnp1vOx3YS1JeZxwRbBQZEB3x27HuKXOTz1JLixheJw4IFrJUKaSIalgAS/
R5Hgu9pEzFsq5Cr3XhsiQZp8WctK9E+7dmNOzljQNQxEFMqpj67DR/x4/6uPNi6p
9Cn8JZlvhw+9sAxnlKErOwio3BJ92LZ2lSTcenRR1JQtwP+4qIdXn2nw8wD3IFdY
xMnP2PmL25kC43iTt+djrPWADw7flPjHWXnI3Llfurj9JtYyEbQSromWhOGhv2SO
lUj9IyoSsOcHA03ZvlWfrTiEsVT/XeTG47Rl0o+eQLyatYCuv6Xm0ejBFxiRoDZ8
lwBwQcFbenEd36FKrpR13I2SYrf2IEMguJPIln/uU5ahmQfZijEOkkUXnGkErl3u
AcN/gbPmoclBNvrxK3O/mayj7IUYhcZBIQuScNNGeF/jHXpMiuuwD81AmV9pC5v3
eZ3l/V3kH22tw0sk33s/pgroDMgiXkd2VPbLz2VU1aqfAVP0grK8aLVZEP02ohtk
XZuZitoEXMvAl5E+K2c49YclGP1Fh+rNGUcoogBtiAB2goXiXSP6Hkw/FuVKGDYh
lMzJgmV7VPLG4yo2KRgPwzdcI8zXbYgQ0lJHKIshqTf5VutZoLYcAgK56Gt6fTGU
ht0mAO9ddf6tF1AEK8YAMxjDvIyPHVONHpXhfYXgAWQ8Ze4ch9vgvyumLHTXmIUL
KKDuKg9r8d12kBwU7BCL8XkbFzs+dQMYeOECW2cNZeffMmqggFHQAZtsQ0jEBx3q
niYZkkQbejVl1ovvsdjUevy0V6EhUgkCgyI03hWg1vW7dP5Olk1i/1tMQ34oC9lE
A+K6WK1B4jNEI+4PvIxrAOCHrr5mMANvWyd1uuE7BUEbqUSMqianmyJ1hsvAlovY
29xtQAHaVl6AsyMaRW9KnE3zj9bhXrCnpMq6C0rn7PVgaDqM61lWKBe/2Y0Nb2N4
43rB0qrqh3EpvbjwYmV6f/Kv0cNzyS2zikFpkKd4S/a4H3TxAdVNNjZdiWgcMaZu
qu5ymgA+lPb3BncBk0tlfjsLV2JjQap0iemcbRWeM74rJ3n4w77a0yhhkNZ4+vvC
6B1eay0JEyUi6OXCwwT8YcNLAWm4oUXFWggpxgzBOwdPLY5ueDsbY/p4AADw1sdO
xyZTZEcBFw0P0R1oa2fS93myL+BC1GC74a6aTiAK32V7VWL4yI00AWH04a7o31P6
izw96Oc5VF41WtutPl6WmHmEP0RMESy780EpXhv8xanGJVnPsZl2aFTwSozRi68y
SXMBQ2heL/0Jwh6TE9fbERV6KHncgJf8WJvjtBFOQUTEYRTIV3bPdc7YcPdKPbrk
CFH5tbnzA+0xG1VZx8fScV/5TzMsQQMAdtMfWAUf2gC/fHxi7+C1HLzvXYYMmxeY
lWBmFYfrL5ks5DmUAqypaXgFPHmu/0fSlpOrG7DtlFOcZTZJnRDLnmUtnq7hjwEY
72ccot89gETpyKuhQMr0EOdY34j0mEutx5N08w45+GivT+l03OYSWt6s8fHk4Jfx
QPXf0IoYRjMFhNRC964KRscQlGFJp3zTkELeDJXCfBpXjK7w9GWPNpJc6mcOvvAx
TcPpzWvh24nY7SSt+3aOgrCutDsDB+RU0V64xR4KZKY=
`pragma protect end_protected
