// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
K071R+3XbYy0vR6bRepgNxoIDn5BpsMxPqiHOo1CIRKOLzTBgMLDbXtiuFmr27/6
Qod+oefnAtZltXgHGvawPKTn8BdI6suF4RsddUJt5MXMZnUG5pxV7rrXgZX6QZq5
bc1plRwxwtiJXZRXJ98xIT1UBXsObUzOoPb3J+2z/f0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7552)
f75q/1mw/n+0F76j20ZPrgLGhZtHixIXubnIfgAF/jo/tWzJgxViRZ/trRfYrE4a
xfZrYzW6QSWix0dlf8cU2qVi7p72MXL64okPVU2NjvA5mrOC/OjsnIqF+AJkB2I0
XalbI5JINkLPcw9rbT2fk8CHSw0seRK5bLRzjhiENmFh1hOY3aWPTa9E4f/2H8AI
Nx+BAqEgiMO4tjgiL5yv1nRz4rcUTTLhYaiU/EklyFktnZGfHbRlApWedQSqYyH8
p2Ikp4VGUfQOej93YUavhYk0Hm6O2AwD8OBNDU8f6J2fdrMiGpw1d269ngyavxYi
8y2ydB+eaem4BBSEVDRGZql2jAX0WTF8nB/1oEOT+m0+yAn2kSslcl5IjI9yx6Ss
9F91dy+BvifGA3IH38sfzwSZ1C5ca7yKIT29haafhs1YBc+amuM+3StVy7e6baZx
+MrzbI2VpHxhJFLr4k+rt/D4eSMr8x4lKMUzKzuNpSd1ZKbcrnbZgZx/qZHHnVbz
qhkzaYmrBOcox/ZGB+lxLglIZgRFwfF6ejS64gDMhUOXOtiZ812QljuA8E7ZQeWS
IxSCR8kOsQLq273bz/+JdHr+1OHScXqjvc2AufTXre7msG9GnFPIDtdjH/Z8/Se9
9RYf+KT2HQ1LS1IazFrebhUFS0OD3Wa7WqfMX4x8Fa3f0lBTXlaS66u/FzyMsh9B
t2entKuVvP5GrS6Vv0SzLPDTHAz34Zijnq9Pv19aJdyc3MAr+KCuXcVMOZV8zMWU
HA7BKwRUpWXeAxInqo/a+OvsX4/ZHK915BEy0fzI8o+J3Pz/IdklO3YRF06MWGpm
GpATV9scIDCLv+rvZcfYYbgT1J2s7/fQIvMkm0GXIHgxf1rKLsKAEzEFXhcZzIK5
KtsahT8M+DtOd4JYpmOEq56UmG10pQdm44s6fglAbal4DJndOCsRczWLS3J/NW++
aKYrMpABePwCj4VX98txgbH3RVlhUjVFN5rIns0Bdq7cPvKipRXquBOu0gsSn0l/
oUI4Abu34MaEPeG/q1pW1uGAzsTDbx7ZWLL/1ud/0pvoAVScOwkJz1AiRrJBzAtA
8foYHyEnXTObgEP8elFj3lWtiMdXTc8SbXcptwQwWK90mZ9Xsa83nbeicdExbIzl
2BvH/23bMnRZiSKi7N098tBUUbkfNaxja2zfwubC5kF7n//3FMGTi4HhI4g0ZDBt
2Gyc7XXQbN6rlynr3RC+3MkRpazrnyQ8hJw6jaEWRyjsIEH6Bd8KoEx6hvyVapPK
oZeUphPGKr6idHq9KKTwLe1BOLefKc4j1sAZg1X0PBFiy4eUsBRhzw+bFnZwwnXw
NiAaJwDJsX9MFs/FzumSL6LTiBi1CwfaYVL0l3EkDPmW4qxX8EOqCtwWQaw2sqaU
Oqdxh5wan/Iisfqsa3njQ3x3Sj7QrnmgDPY2Va2fHj9K7PuVAk4dUYkT/zeFstP4
DckTdE58MqoTDS9fA978skf45BlI8YpXk6D9bO+GuF5ZvrVViQ20+YxFsX9MkzAW
RaIPDYODtAUJs1EO0NPbx+8PtHYqvD/I1hR8chLaFnUS5N7+dhSSg+1zJZyv20EG
tRNyBkUJqfrUCLqQnsX166Lw2ICFMRUtaTz6TIbfNLZc5XppaX8Z8EdCzmcrK+WT
dFHk7aCz0woh5vHI59URGVNgELLjbYJYxtF/pxo643qZCCFrFbADOlI8Vrd2hXyx
n2S+h1VD7uI2yVmgnpanX2h0uPPvF1kV6+05y6bQysNIFe1V1A/J9BZnMosxaaVI
WPLeVDfxQD0JT99O+KQI+13vXF533N6/35d6zbpxO8HXxzPKHDrsWMXPDQ6YgVBA
TNWp3x/tsUP+wXZ7//1/kF8dnvYtJBgE31PTHsdwxtDKBEhxKxBE5fZ0iTVdWR69
TpKV8maQgcRKZwbY1PdxFEOa1AzWcyK5sWbpRjoKFTD6dPdRRpY8VI7w2WA0Xsrm
DPhq228mO1aOmy051yjxQ4p5rdBFrEsSM26UUzOLtJv+hEikEW1xACfMYoSQQRni
Of2Ze3Ivw/xePCCiiAd3D1hD8zvsuSJhdf+3PJN3JD8uRIsaQKTAus08Fp1X396R
MP+TwtdqNPGMtrGaszG8/3pPr0XWtKNzRzWhofxYzwruyE/c1RKcQZU5D3g01IKB
dUH3TPpXXYuqKW5JvzYiAgZgNM4YbVVKzi9uj+l7ffk+UEJp4Cil54TsgGzVVyzZ
4ViT1BqrNjscU1l1aiLXvXBEswEkAzDO7BuCjzopPdgJrqM8ZLytOna40t4uNWb3
SYDZdkPwBSS0KobPTN6dQg4YQbupZKlzM2oxxEF7p5YYNlh3yNStOWKmozcrEJx8
xKM755DKIq3s8Xbt7tFY/FfjdP7LQ3+m3iYFAYF0oc0ObJgYnFVGyQ5RBCw+MEKn
pscdDuKQjG8QdCiCDrLxeQmVFmluejT0DNtf5jjC8mAEAifAmfzfp0SFpEE5im8c
veu1LvmPqfTx2TiCTQoxbktzj82NbVtpXnlC62/vAgEds7x0Fzx1d2kuvB1gG/Y+
QVYTSc+zU1JBtdkI9Yx8sZTACYIJYGZyN46Eq6l72LK9jQGqyQaBcUJBnDsllDEA
6EIxg1xPG+2CfO2vjKyPRinNC4C+y51PGpHqfPKNAyH3Sfk52esAaTsH/bW8NNns
8NazPeLaBZay72YAzzy8SbZanDnQq6UrDjKWQKEIsJiw3a0vsaur+E4wg7ls44mW
G2s8aZ1xJASu5TUL+KwwhOsuIpPENr2dtc7lPwlVWcwKcZEA9JHvlXnByTSMUKnI
wQrSyu2FPLJ7Wq7Jlb6yNkFl5Xr+Vm+p4PemkDjLevH4KYDpbr5f4o5OElGVw9qy
MEIu/tT9VGykEuS+NJXV/Ir1nGX27+t10Adb621q2DZBjxdT+dfYlGgL7uBrWjCf
EOv6WkgRO36L3vG4OVz/3In5nidWeDgUtMEvPePPibm9278psHgMfcjIjXV/eIlL
W+YMLwAKddNLd4/oeLbN7khOJmfl4Be6bCxkxsdseva9xKN50R+OW4Pi1N46cNaG
PxiELWEgVBzmkW2s2yX+lIhsXfjXjtGWexFQco8JuasFxgY+Z/x+CZNoUv9BvEuZ
xRacexSuHNqAeNqU6bwdyVGy7Ziieo6Omt5g0FfARIFBKKTEXet8u3P9FaeaQg11
h9+6OcoMaFC2ntmfS+3vcfpMp0ALo2+FMfgH0nt9wx15H8LUkUmWsyLjPSph820g
E1GYl7cxWOdVFt5Gm6GeRhWf60O8YkTdQUij9nsnd+wwheTZ6511NqmiRH7vSv6l
OYpb/Z9tsQh8+Mz5KrtGz56JLJomOwNMzFXJ1WZMqKozurAQEOjS8/uJWJhA7FV6
Dafzw/CtVJq4sHLvpTV8BsHruCdzwxT90Oe3Bd85Oy6NMlrmDvhe7FtMsbkGqNsG
GHllRLGDgsO9oIW76keKLGswImDkYnq6ltT4k+RkscRdy4iH3JFCeTB9Dp1HEK48
zi4Z4xKLkjDgn1nfoEejHVYaS2s+e1BYX45LX6ebhA9gwMfonPPB/1Lq6rb6/G7N
FpJH6lt7hABg51h/9mEtRlilC8rSpDi19GlALS1A5pOHQltCHM+v1qt3tJRuRB3L
Y2TlCWQhyZUIyNO9loNk5B0t5DWxqqvUqSFlAdSQzp1c3OslXbR1qaC/wFL+14dk
m8nAjVdrFFuUnJpLCIkYHQT688TRNBHjO+7sB0Iw9rbMoulS6FLwoadSTOnf+XKW
zCKa6cbv2up4nCplseMtRN6JmZWFtOEsi52NURH1Du2ExELpnBpxQVAEDkC3PnNv
5xj/A4/mwQxD324PmAqY8VWdgT8EPqERmcyRox3C3Dl+0fInv497pMKPUeb6W7wt
rccrYZ8LtuC1M0WLT/5gc/4XaX+6JLmI1xcntjXeHj1EfF710c2m1LyjLE6st899
v20Bt+Q3me7sWm+6A95Lt4Obw5jasIxwpO2nrBzi3zvATWHiHad+WBu0jjhP60iP
wafMF4XjXxEXaRK3wGrlCLpHcdB+mtGnALkjA6weFgBsqmEiIO8gq7BOuRye2BhT
uJQyoaXwv9VI6winfPq3t6/88/cA6rCaSC6EzoR7YbVuSqoDBkjph7lEviPrxDSE
XqVPigmm6uvMA89kBZyp633Q6oIWAPC0/WbSnnlKIHEG4w8gGJZ3s1rAaAx3Q82q
vlc/iAMDaSwepGjhMtwopWSCJgCqkWuhaezENw8OXU7w/R80ceHv1K2sVKW5Pr9/
zXgJYIT/hjsGWQaD0O8SqqizdEwSs6tUpGJ1kDpSeK720yQ+BKGg0lX6e+21XjFn
+PlF/cVQ0HTL1Aty3MfmD6p2rgHgpywRaeIsy7EPIO4eCuVc9psz+x+g8ntMaE55
6WhvjTqKGoMmYVyjgjrLQHS/wwSz/7xt4TMZKGdMuxH83C+Lud4T5OEHSAfj5v4R
e1R03iXKBsDwomc7E2TMPVKLHrHkIturwCQxEBc+zbsXpnKwHguLW/zlWOMxFf1C
J2NJ6eYeZMttalJYVd1aMX2Rhfkb9Xg6rGR1yMZPy9ua/NEzXMKGDuBAuGtGk8cI
bQLjU6lsPOdC7eSXPZqMshksV03DJbqwsxTgmimxpRZIAhTY8Vg+0fMqzy7y/fia
yVVy1luBKkXTcBuhc/lpCtWVMoI7zeq+1O9MOFgPUIBTFVdLObxdCMsFzsVWUlkn
slcu1QeabmfIQ7uPj10mLp2VO09uJAITW7qQIKk9639UbNz9ScFaRvmNMR3YsA8N
3aD5rpO+txZ8a/xQZK/tpAg8mA1Ey8wUD39Vsz92DFpmDN5zI8nawB8d5RKinuMt
4N6FTC0jB51YFMcLvGErfjNC8NBmZeQvfL8yTauK7WuEM0v94SqFdTZTTnGc1ztx
ZZpfVIKG3bL88yb/qzEsNLh1La/0TQvknI07mvFL+DeJW7mUCVXsWy/ORhxw3xy+
xNuOjljDlZlBGHY1df7LGYFXAEsK72GMVhnd7KjMYjy65Wc4F6p+wXY282T4WIh0
1Y663YdDntmhLSFbo3/RS7v06uSpQ3Cl9+GP5M51/z6FOA2BwBne9U/BSFanR83A
jiYtzMXgomyJI+pc7TfFggC/llmlV2u94sv8QUDVK3SxqRfrYMHoG8LcyFglq1Qe
R8HmHBj1qTzhLnVVw0C1EFyB1yaf0+pheuHlnmpU5hk+8h9hDGSGRJr4pfcxbP8b
0l8pFQh0tBT2FvpdlorsQphvVngxEi45GgC0vTkLmuVuDjaMPwh+NNxq9cWtONvT
41CmOY8+NdgiAR48TAvdcvlD4wKOJCpWQsoJLRfjMzf9Abq0uvbFhn2fINEilM6K
nq9hNtd8ILI9WPobIvC1CbbjnJDlnWADdVpKOOKfcNZbiTYgUEVlRmOKegqV+bLW
xdpDGmgtx9VxTJxhQvdNwUTV5ZfrTOyx1QI6EfAl+UWSzPbUWmD4dWre1Hk+BIUF
4o0+gABpuFrVsMxXgTEAjnclumIoNc6Npv3Nk6kz8f4omK/its1J3muUxr4sjGUR
dgj7D25IpT7wpPtc4KBMIxjMESpcOFNV54h9379cQLtFBZmv+K+s5W3QZA85oufB
V1bqo28OfG/I3Vgrg24OR+xmV24x+XXwhAfywHuu937cqWbsqsFJf09CZdqp4Tux
uPlFjfvMBUvKWM40ZfGUk7XhXtty0jr47jSNKZd8ifypLc/4teDNJZLMvG1TBtbZ
16t3vQa6k+Ej4f6/C0yHPiOMj2LgJ/QKvm2865Yd6TNgbORN4cOPYDuHo7uyRqak
wGx+uSUCU5aeNmLvAsgG0X1v1ftoqAm3E8PJNIMjPgoaeSa4KbZtWwk7pO6RlVGv
ssOSax1DqrbDN4QKsoSHu4DGqa5CPaCo40gXHYGsOt8kpAFHho8QoT3Ys2OCUGJf
bgFx571uvRMpf6kZuyPOG+Bd01ddmjvMyV/rUQ9pLu0P0IUOBr7TDyWw6fUzIXN9
SjfyGE+svyg2xQfJLHSmUT9tey/9yhG2T+w9JgCxieYmbX7dEVjWywb0BDTARM6p
qC37etl26Wn1v2VmHL1qzwwFlo6U88bRemIIOBcpyE4uYPGo64VwkfIzdgK8vFHi
Q2caq4sMHTI39tYfP5KlRW4u4sVDlzimio4NHPgeWZaIUvW13KSAayBm3BIyqrSn
fmieVsOhA2MKV5rksA+OafHwj2ZcHH7F9LnEcEvFf9KirxlP2kmyeG+pNgTwC8zg
rkufT2holp4866P6fZhv0KOYebXrLAmD3vvU7ROiohivHAuaExdoO7ldD0ilLJkp
E2B5lEPq88Z7yyCfun0ppLGWDDa1tBk/YI9W/iS2fBeL+cxuNuG7m4R0MMChm+p/
iYjjJZ+o9BLp4tlgovy5aGQ1IInBHUmgP9I3spO0hH6KtGWk2Dk/ybVbmGJbAqzZ
1H2nLBWgPmm/NIhPGpJU9EYReNoKGQlLhPmVUHmBZybX2Sz/HxeztYAzaX9vpy1L
Wp2ooRgbf+SMjDe0nIY1pqiJVA56cVMlTGK2z8An0LjrlbADcd7D5+EL4Btjnkr+
9wSq/TpETGrAq3yvGX7kdsmNKsNH9BEw7dmnQWNRU2fFt3ofKUzw5x55/IRtj1fm
h6thJtNjNLJW/z9psDx4d2BSTd4AVLruBbk1Xxq1JpLVltTClSsKKtWvtodBg6T4
cr7vIQ5MwPQzCbXhBsme/F7oG9orkIS0wzAi30BWhkRzTPLJrkq0sDd7Msiqq+hG
6tRUs/38vlOviO065nrfdws6wym9TTjc9tzNafxhozhaSny7ubDAYBUkTI7W3yyR
exSt01nzk/u+l3zttB/zmf9T4QeiGvFzBpljpWCIwTxpKPIFOaHyp7omoyXcoWOH
KZoWC34HMsEb0eMQULXOgZyVDTQ0y7Txh7sElGK+78hu3D8DbO/7UNnWwD6R6+hV
wipPk1AkudI62irnvo0DbWYXTEJ+QKRfBtryZLoJdzX3gc4n/bu6hnRmgrRElyVO
HkFeUL1FgVfpm2vV9nf5W49TbkSEKeLCSHPwHXqCKmDnz7/K7J2RMLxRYJPF2ETl
bG2SKTxmOArW59imoUQC327gba/gVtvAW2I1QusVfuUHkHcCfGGJSSF6UMjNAyhX
JqO2Kq/14/w9PnM+J5n6l5K4XD5zYiSjSaI5DPGVGIjuuGVPQHNeAeNE59He7a5U
rPqigwf/P9KgJP87/iRu8BKB7WtMxRc//r9slb88BjHt76UNb5QxUY5h9JkqQzft
XHzGEhU0KpGw9ymb3FbH4GX4Ess6gTxGsf+ISsguw5nHFcJ72FrITUw1w4icbkB/
OePcpQk6oVPgnKjL+n8jPH8GtjbIRcng7s/Fg9vkBHAku6Y4X/sT5kVydHLfNwJ6
ej+q1BnhW15gL6iOHPm5ORrd8MNDDbxiy9uiHDez3efHBipNN6TrZtEvhlKPeYiD
Tm0McpbwY1655cJhr8TpGAi2ARDWXege+hg4oQ7UmSF4XZBa8HqZszbaZH2+kw8T
fVUnMxHXiZv9tIZoRvDHEcdgWMiNaQvmzxNAbCvycbwqEaLIHP8JO0lVjWqlA8f4
yLNGAT076wKBv3XYEX34rnsAjFpFpzF+B7AoeG/H+n8MUaPJIqRMf1b4jZnAGVBN
gdk+G88zFFEK5U9Mm2XbnO1CYZo9HnvUe5KumJmUCIs+cWyAmwqXi5Bq26OKvQAG
+kl+T2ke4Xx1HzU7u5/ZbmULeh2cbV5xhvxxdAvo1/3IcMrHvTiaEEK8h8F48mo3
6epTqI7hIJFJBGtbAAX2fnhtcEJ4fKTOD9R3445Aa1jtakN9CCftvIShONfv7llg
997w34IcQOGvkkgn3o8qJsfk9FXGuzWqQ5TtEm7sdG32ajVPKmZ8L7AEuREYZWva
T/l36PEMc2MzHQQJMFF5/hTGmgtzZPW+ri9IQgHgP3uYwgPJ7xKu7cjmmueHXAb2
BmhGZlrLEMb7l5WNuIMuifP5+FGpxQSQ7PeFqim+Tl9cTIF1UD0jOpKQugFyKTF1
E+4hg0aeOb6oxhrJwsuM6CmALAbz+57vWYoi0iYJAPDoNmFyCBx6iWYEDFwg5eDD
xGo6xeZEe/tARtkhc6F72E+Ht24Z3w3QfxrjCq7WPg7JyXfaAYIorLcUd0mDeKqh
0d8qbaoqSH4BGSEVSS8thtes9pRBHzsHjQQRUcwi2wrGyMxSvQhpkQyHaX/h5f2L
SHkFEbdMs3qiUQJMzRG/A6A9txPlpNC34z08R7NMMBfQ5oLQofcsu/dRWtgpqO3v
WbRHwiY1au/5jVLbr2XTGYRTNnp/BHqO92bYvGQv73lHKDUWIv9iWrJHWs1s1rcv
nQfSyGaHHGCFrhwgKvZZfKnbsZDcRXTlvFXcx0CHGn5rLh1L+G1wPTbEDgvZVIE6
GbCyxUMRvVtSUIUBfhRveEZKTCnyThCGzWI7zpMGbpYNkBFDW1n+kcmMtTwSAwzl
SO9dKqd64L0Gttpr0V+E5NXpOCsLPfvg7ZRwyYiu5Jwu7ps0bjSQavfDw474bFXK
d7kKDtSCgW4Jok7Jti9ExjMb2Ke6VOx3gJB181/qhUXROBnK89as4Fw1EAVIgsQX
0pvwdAzLznbQEkVA3jVkwaO9i+mau7Id/nVgkRAOHy5Lhu1BAe1qfBi3Gckh0k/4
tQXsqtaOAnDTcpmJKxfBccUxqwNEqf7ECyDO0WHEQrHCbrEZ3yCP3F724MOgjIWy
PCOa8lyJOqI1YAd5hq1h4eDmUL1mHz5e7ZOBTyEVybJbKT9ZamoyoDu9qs6Ziq3a
zljUuwlchkLuiJlDUxshSfgrOkEpl77rM4FDTcOXMH+SdmEgHvTYMwFlrJ9zf6xj
GJrCijQLkpcJ2GY2OYG5KKvS7ts3eSTFkFJI3296vc2T1H8mx9g40JmV71eIQ+Vw
cpil/uUJQqvglZMiOusgT42nVK3+CSigXJ7qJYYL7MqZH5qMpNWqDEodOHBmz5hB
2UTRY8N8JDbF3uDztlH5uZMPJbB3qoUfbMUxXjP9kymKykhhbV68rYqn2jUeOId4
UivC59CPzAqrsefC0+XHWVHxJJGXWRub0StQ47+SiMBTazYTZlUF+SSCPOKs+p/g
E6oO003/FHKBAVc5ETgwxmYuhMMAiTThDVprwKurCUVo1e4GnmIib0pG7nRfoDlY
6BIRHBNtGWQxWWlzd8SMVCpeaYHsw/siGVS9cNLnmrePYAJwrRHWhfm578P4cbnP
F2WRa3rEFBvFbjK/AuScTwpOXg8lqBaOROB1huHfaESss5XdOPx4MVWLJEcxSh3T
VZ1g/jnTH2HnWO6FNeRlgszq1pb+N2hKWiQqaayibpOEUFxcD8ObsQ1PjlRUJ7g1
EQWnyuBPxnAkm7KDFxKnSLhAPWHAHrX/kXu7lE1iIThIBrvwVh7t6xtZCilVFga/
Di0cfV5c3Q2VtgTSbUyhkhZwhSA0NlDmCVO1Q0Q7URhopt77pBow6nZ9WNvZ6/gy
d4B6PCkwKeKhyNkiaUoXpDr/NTIabkFSp2xemLurBk1wr502idzWgkR6mbSyzCVV
8TvvlKLGX7fAHuyB9iThp4rULYTZQ6o21+B5GDV47B/w+IHV4x4N3vcMBzd+cZsb
IYzNf2W46QvyNVqpPyZeuoMndQzVwp1MEXpMjbzcfMFP+TPm4Bj1jW1dF8vxLwZH
F3vX4Rh7q/iXjTQbujw8+0hzG4qcYxZ0Xy+qRN1EJCge4fTY1szcl5t6wGViSytu
LOG8ByvWyT7MY1bikR1IqjmzwcC2uyLv137oAWelmzX2Hx1tFiOGH08e3I+e908d
6sA4eRBpHvis/e8Jh2/pJWYHbZppwt+kIwKBQVirsxej33qSFGkMXLkd+GjuWIBB
k18wbac1z8CAaT4LF8GOs+kz2Ksw61B0DH7vNFGJGEJq/QJ+4JU18SL2EICWtD8I
igXkb0BOEAfiHbx21qK0gLVdm+MCzTsabXJGeJmS0Fhy4q1ZKl3sue9vqFv4XvxN
m0l3AgYVK/0mh1RvOfZ28A==
`pragma protect end_protected
