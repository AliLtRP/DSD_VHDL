// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ICy0qdaixShlFyLvVOfD69xf8hxvURxzM1qrLJcvtecYp07mJDEN41FTWadbEnmO
8olCkxcGOwoSHXsZRhUfmEZ4T+Xb47oJkm6F0265kVbpGg10Z4CWhhYvvFQiUzUk
xg5EYrir7KJPHbNXJadgTXqjszGlaPpy+DPTQarMymQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19520)
+VtNOHo/in1aWsTXgCKPfYTcmsHVj5tBmXu/3FEmDqKJIhWxoo6/3nrm0LSWlGR/
pR6C7cdqfNaPlaky5Xs+FrALeJbjQAKkYxNIJXrOJ7cpBbSNyEcfflhqGTwuql55
Wpc1dzALbUttedyhn/FI6a/ZA6gw8ig/M3kiGFU0kn2vJojctrGFiz4HDwvgkFKz
HieT7VmCaFaNgoxKyNQJzT1gPeFkxCt0OLrwMY6HtflSP/ssw2RLRchSxiCiLMMB
FDB14Izi0MF5By/C7S6Aabz0XDEERGEXTxb498e6bhn5ADJ9WeaJj1P6qVw0PaDe
w7/wsGBJHPKxUULthz/koDIDt6+FPgps6vkLicVbkWVn+smHY4OVcSRNjBJ0pcil
oraNLF+yGJE0tOxoZK0kYtbyfdeaUNsJaalgOmqXdtBdALzNLIRvg27y/fRHPCfF
jzxlsQZhbgdlFAJ51sxyd6YLaLxOM/tC8uhSNEvHTeaJMGIHX0NLZJfxxAS2HeEq
rku35QCwMjqhuuE+hVnVPHY2N8VPDU3y5vFnC32CaN+kfq3xwKEICCMH+ypqTAIA
tO7Bla6cCNBBqI1SJ53PodQT3TXNu97fn/Q1ZHNIIS0AXfiMQaPuFqt0KKWyKh8M
rTIeo4ZdXjA914n+2/wk99hxaYoJZmSM40unHWVva0MuZGIFHVlElBVeI8hnJfTJ
Wy6pkRS+BQM6i0P232YIoXdJcoHG7mLrilqAS0w9vsmS6Qa706yFa6jPjVRbj8SR
E/C7cy1fwCbeBUiI/M2jJop3P9rQaWK6Sv3GxOjM2cjJ4IdTpwY7Ty1uzxFe2HMe
GaQWSLwGG6owb81RKoWY0D0/fld9JbmbnGI2U7QULggwau0gnPF01t/bNafFMyR6
96UcAX90kgwpwsjyCiQwt2xeSQl2S4H/MbF7qxZf5riEjbab7hMt9cFNgoS43g6V
hdTiaBLyV9z52PGXqEpSZDm7hDjgN0h6iA4thF2mXNqqk0AfkOgHlnIvf/CQ/Fkk
opd3wyP1Y84zMX50uuoo4XWz+G8I+QfdUEYn0cW+SCirWWlTP0diuFqPZ5YshmcM
1r84P4Mdr1Npt+LTttSqNGm5DAfYFZYB/qeceUCKE3ivh2sVBpF+9GLs5+SUhg97
qB7B4mR9CqmYeBdpw5NbIhDDXynwYk1bDpYZecTItXfeXLOsFKVImEwlMdrNejsi
QY+vawMerx6CBkjHJLvg4BJh9z1qnsdR6YR33AfHT4vuFN5w6NH5kkwzQBWTgGYe
RBW8pLKofOaQsAoZU5i8fogAEdnJ5LoF1rzzSHr2ZVXhV9PHIIKAnTLqza0g9MfA
U/YRSlTMTKnlCZjwT2Y7DeJTH5rW8EGonCPOCFV3tppyrWjfqZnaGWFM/Y4JeFN0
4eZUGqoe2eVt1u79y/E9eGz6kFJzFyrzPQjXkHLZlQwD5U6kmeouNjhrnJru5LnC
XBjiNlMDbSsZ2G6fGkeBbslXBV8y+hNm8nSjfj6y2+BWdyPFjFN0nIuGtUNcT5o7
+xi5t2bF+1bGTESOr9IvC8fat6ODUebS4RMmutCH7n7ZKKKafSnN3ndv8OvIEBG4
RMwDRtunCr/vekRsJ0hvE9I365lIiEHYquq2KFelZu64Fw+JV8VytyzDuyQB7SSA
Vf++ssgXOpUaJHTIGZ9aZB4liEwFsmwagsu0e5F38UjIwYpLaXWGbJDovt1Ea1aX
LidJ367OaXf1rZ11JNIZ0kBcDsnFq9ySQz50rHQbbEVbFx6Pim/X6dG/CTpWcD/t
0JcTG2O8JtlemXrWsq5edaKlxsB7/fr7f4MlKIHvBHlii4WonjQ0lv9idjRKSgI7
mqC/4PDmthVZNpFMVK0iLsZfYWtvn4/CmjBJQ4eUT3a3GPaaT14YjHpx5VAsJMKw
Qr+hPve6WB++uR0vUSIXR+A+KdwPD2BrzBJHdehYtNxIVqVmSgdToQ9ty/MEy+AZ
ChuMSU2K3N+Ww0/pG32zCvX6brsUNFGYuLYfnd0WKvHO2Bao9d5XZorFKOgpLVkh
QLQDGEivmCrvgNYQKxh4SD0Kyi3NDVzqq1T6bePkOFlprQh+Z5WB4Rye1Ee1F3sC
ulQShNoB/As7VwK7TQenWL7OeZaHcyJtpfZmrTq9my/v0F1T6/MIPPBHaBAT/sK+
Smhk34Fvzo1e16d8LqERDzrn8ezveN9/QJg6aKIjcZUldLBBPGqCD0sgVwlCiV2M
q+vNPHzam6WHDYKXHdm6DkBeUgVSlJ8mtKv1aq9lzX9b/by/zgYYCDSNXViMm7eJ
XHaaA+DXCenbovJiTo2Qv3neR88NYfVlach0yRxQOjTdpJtWQ+mhUz1QBx+vLkIX
Mhpnc6Xhlzf6LgzeBs1VY78HIhI4G9LeRllshtTOQBCTj4vinrs0x4hQN+5eEb2a
N46psnwLkiIwKqCxapM60s/cIi7r6An0jiy4sDXjgHuTa5nLbZZapuAqrGswYy9j
EhHKBYwGPDMrm5kFMjiRwbbuDynufyuw+AIroYenwdtk91ZlTu7unT4pPUCJeILO
A+HR1ke1DLKweqVpAVP5Ie1Vzw7YPgeQPV3RGB/SAF1CUsNMN0xaPYRDJle2VyQC
ycL58e0He8BIryohSCBjbLJqMYyJA4XFOL6ZOZ8p2FzTAmwlJqbeQgqWdwCwjYJV
w1mCJU/iMRO1X0Z14UqKfT8MRREJwxFssORkZRW3fKJmTaAta8eXRUHQ0o47ktrq
vonO8UH407w2ZAnpOufnUlRIUqRThBAnqHvIx1KMsZ4aGKpy1qFElxgbLmUMC5F+
eBbOzvwrVx4GcMZmTxmgfm11pSllzR8mN3R2qf/uPPH41TxXWUgD8b3FTbqtPfmj
j0KFxAJbJ4a7zJVzeWbtDMRA4adIOH2RD+wGbifIXLSRb57y5SW/BVxhQR0R+5Q3
OW3YpBjCyYW3i3lFFOWc8gPzoNxJwKjQbEAcjUVYRU7T3IKtG29SqjDH03DIuZW+
beq5sUVpZiw6+XPztY063WpGzlc6qngziZQXZrSsXU/R21EmRybRS9/tGiNTpI7T
48kz8+ESaHdfhChaXmJ0/ybnNtMiv5bz2b5NaFNfrMPed3N5CXIatN9i8XUvAIuB
2jl4ADqr3nkaR+i9BQ96umRlM3LysYTfEVtUVwyarYAWangogldnOPqgUeZrdjpH
nUHOmuWo0DGqSvQ+ixsbk2MOosL7GKfYjbUskVCoOYDJCb21IJKuNfbVUviq/tor
ZmSYC+6NEMGXBC1J/eVbylc2mNuFSDnfVLmmCCT5VwgFPP2ArniyTLaneo6tfhr6
J6N9w3TQkERLsnvS1MPdqjDZa37RVwFltApbllAdDlEJUEU9QfIlrR0QM0uvY8bK
WdzN/FPbEWqt9KZg3wMbW2U5B3WjGWPA5NWF5zYzkb1bAsIeJLhG3Nc9eldhLzVC
cvmYV+A2w26QcM15fwQrHn9E1mwcAAgIwTwkZ90qeQqHixF4TvrsnaIuUzEzVcpf
fXtOfKgewR8M3pKwcuv3QMwZJPxPQoYtd0QXdaIVRr2c+m4/SSEK6uXpnmS/Gg7u
rYgOOtlIWgdZZCrjt5BvCyO/2URkyC5O7hq4y/XTlyWMN9oDnEVKK4FFgONGeBUf
4kh99GNSSHlJJHtnfnckpH8GtLtquE2m2tQRavJSgcCE4c+69WH533vFIY49GwOS
bsldrsCHgoEMeoT3ljgTuJHf0fNeIau471cOv+xf77/sXLQ6I3muQW6uVHTQi2jK
ZpmU3nXWS6GG3xp1IU9vq61loUnl3xRorFRbuqReg2zeHW2pdvlTN6f3r9/Y7Se1
7Djeu0YMrHeQ7bhCJgnUg+tQYt4yLdlVKu3EJ7TjHsZxskUQpIRwtdwUnvx3p1cm
O0Ox0H9dfeNuNfMPzbyDgwVDn2cqOIM9plkQiyoNFuN/0UGv7HXNltsM6/6BgwdL
oKLliGB0TGlxutxcyxIs0domVvJ3dkFnRPREijN94rJIpnrGIVxq+lDlRyDK4pzV
vxk8kjoxy2YjjucxkTFIK43c/FIjiiEYXs484Fe2WheA1DgZaV3/xrV8QahZfsJQ
JeOB4izcYBvunAXBF9kPaiTTl8XB2leX8sA6PGUiYWndb6T+inAScUA+Pc9eux9r
8ZkRtG7AvNhrny3tvKT2RlAOU39VgQwDAd99rH2+zw7kEppxjobvpmq9svxj5ctG
3onvws40rntyUDN5X4gm6rvptR/ZuDFijl5pzpODT+8HbP0zG1aBWqzgZTKz43l1
atBx02acct/8SE2l8Z5oF4g+hkclESWdAQt61t/WmZDIUamY5dezzZhDMO7b//+X
9tVD+iSJNvWzPuZ4eypVX1H3tp9MWGT2pqZhQT4vOv5EmaKuljxiHnubLnOz1EO1
V6lHpAmY6x/YZ32q9ltc7/zyn1iCTAD6i6h58evAtiG/bNjhFIQcEOfqbiP3iLKT
6HWQx/63FrExE7VAa0SKPHvDm8y+915FOK8Ev8NSdgT+L7uMdVAm6UDml0pMs9y3
p9kyARgJ/kMtW4QNrKXLY9yH9H8feEnmWqg2msmP8GOH+qwlTw5g9AnbaWcQZahi
iiFTTe7uRLa53ZTwGKqsmlOa9bykSkO6AVIziIxc0NeuajhTtNGyJMUIxKrriiRn
fUynT8cDR2PY87BsO5eYlC9/zBBWO83QCkEszvLbR4Cpj2/7lP8Ia+vDbOmhCNkm
PKobPFv/mpE5K5IV2ujWl6b23v/58ZUkfEpLiQNLKst4SXIlS0pBXFTRDy/cG1ut
QQxD8Qs2pVOjpJyyJb7k6yjgjuKvb+LZMTY7iLOtgkENvCJa3bpVQwlyG4Ndx0n9
jAc2D/nTsh/C0SdxmOxkwiXEhfthZ/cOELHj+xlkVDd2sU/ogvHu21HNWO/BQ0bC
iDt8ptaZMdUlXbdQ6go4ZQ5JSYZ+3JXqpQk3X5XJq/HJPKNxKnWh4VgxkUKNd/kg
VX3btJJKz14V3Vw2hT2K7mOsNMpi+0Pu1bLIst63TyoJxhADPtw97Y/l/X73gsFO
zOtBcloddZ9hPrsNIeL0xObShXnpEA57sWKVd9IzL46Tcn4VmdOawJhQgqmI5jFP
9uIZx7KDuD025iIGkf7f8HmGZ4gMYxrlPj9kBRV8ePfYiffd3W8pgc6jgc3bWgY/
JSZgtyJO6qpslx6KpAtm0GxJV4awktX9hYk/8r+HHdKn6qoSuvEEzBmTvBf0vS0H
ijzZCl5XncRfLagJTddWnJ1eY6BmpSuJGzk1m5K2+myJGA1NCsQ4PT2qlhJLQQ1+
YvwW7OYkhyYqsCpj2eod5oQn2iDFge8b3aHLCf+9NrmO9nNQypBMzSIqivn5Yh0U
HEKRWIl+UYz+mVKZxY50P5ewSNy7GorEuU1FGeaUnYdphklZdMRJJ/I0tjeGxyaU
cSYTYldHJ4sM5SUb3JE0fSMIfdTYUvFjzWEJQLEly/zvIWTzW2ZTNFa7qp66k8nn
iGjcvQh1OSISySR/BcIJ2AeJHl4hKh6rNt24iJRUitwz0246/x2gRymNPPKuFS/Y
DF3G27oROeBiuZawVs+qs1LMJb/rPzEroziHwRwXEgc7HV5nRudoyqnpKcIj2ffO
26aXCyKmxjhbCJPH1fj3jAO8qvubrZjkU0KndI51CXOHRaMTJCUlYliS8CvScB7p
B5TFbMI27xExZuwo9BZ5pNsGpSUlsTeV+G83kRgaKPjFl/zhtlxsW1nugrmYDwhT
zWKa5b/gf2mHNV2/r9F5ZKGXhj7WLPcAkJamMV1VOh7F1bFjREZb/swXvHIOxYKE
GHiSwCiI61ZQuTbF1BJ2+bIzr1cTgIbD1T9IqKR1S5i4gHLpStg/v79Q2zI3IZNj
qcBcPUiaBXdWV3IKuFqo4lsUCxHHcQonUqo61CZcJ2eyrwe8m4Mb8WWzNuQ+j2sC
5Oex6HAEu93Z2avLhkLKPKkZPNkl2rAPqxDGJJdb7yvTQbXFLP9Lrim0p12N3+bi
kAC4NMS5bMGmYbgBqgltAbDXl6a4YZ/STVAQH/hfHfKXbMbCHf0hScHkdWM0J84G
Ka0/uWigboRgjxpnlFdJYHFc2OmrdLMwxRDSj3rqzLioivLeEyG3aYuvQvGW6lqO
mE+0RbsZxgX2A8ultvkGHK1YiDlTLg0PtSThnpDXo4pUBursASAd0U57+aBcL5Nb
xKmzZkM4B1lFhfRaAwkJujrmTVRoV4MOtfyo5MpPfXltk4oT411Bu8D7JuZqrQCC
qfOGkOYTBmn090SxuxCY7Kks3/hZ7NUdtY5JACXLMHtPPUwgu5kT3ijzlCYmw+wf
YTOeGiiPDDH3gVih52KFYVimgGPLEtoVwlzScWJFEfFcimhVHS3SnUs1F/smCOf9
6cf0AIXOShBFOzhBvboqtVNFBlG2TD29L10ndSjwHUWic4plf1GXXoG2V1U5xfH6
JSRg6TeVa5HSNmZlVbNMdKX1aZW8Ea6y7YqpGspq8IaDIOKWbBN4Y7gxY47E62UI
wWDjDA3AfCJX72iwIn5eUU6XGREe+FGekE+a4mEwQ/cQqAKCz83DPSEgOWrFqidt
TcVta0TbBt1P1zrCOW0tDeCn2jYfajJJWEHwJQdTohFVzmeZrwuNTS6X6lTLlvHH
wmhBn7FjsG77X5I7ZPGuNYgNNp2C8vgkHFPuvFhjM9+q9LIYl2sJkecQggqILzbi
eTEEPtI55tjwcMYIw8HHbMqP6SLhC17mIi3tTzNUWxt/+E/I3Uf0ceunNkJuKBNM
s3sfphMBBVbJIonbEhyJuzhZrW0QhDgXbZ8xOS7S8m0F/ceUGW9El4cNVoHiKHC+
9Ey6VHPhxsnd7PN95PrtFzPUIYo6Pv/v7abxQ3P6Iu23bHvoruFn7JWeg/VGK4pq
jqZD9T43AvUt9VbQKSBs9YhL5DL5M5YZ20iPamke5bUxU23BplR7s2Q4x/yomS/r
7445RKysiQiusy3Db8ND1BZVrDnesfm1sJflEfAvzu4AgX+7PmzqOrNgysd0efLR
i+NzryGItwaJotdKaahCoQjql/oqay+3RUOAVdmVLkVYLMOvAne4krpsMCkKe2ek
OqO9Qb2nVLRhz51CB06vYRj4oulf2tgWcDu0lLv9DcAv7CAE3Ks4z2oQsbphP5yW
aB6YP68Q/c8+J56XVJjG6bOby9c36EXt/3r5JtNZeV7+lw9hJ7h9WUNASCDat6Lu
XLzkn+/Piv0xsvGX0RUaXmelKrZ5KCv6jOXXfLkBth7OKhhSH3dw3V2vbe8fG4fO
3xX21khHkGmNojT2Hhee8uP/2rTrkiUZtC4/QHlqh9GhNIPbKJ6hKnkZQL5Q0kYb
OF2jyjY52lOUGNBskAcrdkb39l/ABKBk70uIkwePEqu9HaJsXpNbw2A+cbSWG4cU
gin6ZZnmetMTTklzvRP6JzyY/V8xEZ0BxGQ8y4T8OdVlPJJk7zJXYEqDmzGJfJHh
tQDuUAETfTg9CLcBB/5LPkm2p/FqFMRnowswR3FHtAfTI7b3ziDB4TXC9aBycWhL
3tC4PthcrGD714sZt8LLcyIf9lPXzDGRrdA+eYLO6QL9RBSb4qgqBfolMTdr3Xzv
pv+fFaTo6GtVYeWUosxM4B9YVSRPoUmTC7k8hnfNPayIEnxTIk3n+Qgs/YP5QlyI
HdvvZwLLv5uMviP19pNMbzP7VbdRjAk9UhQeyQHEykSNf3x4AH4wh2ZC2ocMfXh7
CI8blpCRC/95Mn33BJj4NMnPHZqZBcfIZonigKfk6NHEyPK0QIIJ2FiMkoIXv2+0
+7iEBusi2cF5Hcj9MqpkVSWnPzUmRKjWJ6/OLuupw+gwkZSnL3HL4TYTPYCegqF0
fjaROY9SIjZvEr+/S0l0zHOFKaXIPaKkFxDAfnv3CnTi20rHYqwrCHAwRvaP5K9H
+nVxj4R4SDv1Z5F1TA1kCmCk531lugM9wccktAwJbXiQr4aXWKb6dpU/gQ6RH5da
TJ/d8v3i9ydW5Kqzvxk4A9E4l+KZW/H+5SuA2UUJOtV2LwOiQv+6XtGvuLvNIFzO
7zBT/ve/AxR1MONEGp8JpVjK+rwgVhSadRYDj9th5Jq8GqywiAPVOO9rCKlFvsJF
t+6kPDXm4QbmdVu8xZfJJZBE6OXZkKRM1ORNDmHtqWZi/it1FKXNmQ14Fi/xTlP7
MCozFoI7GpPIxUfkUNnHxqj5b8zy5jvbbx/NCuubvDUf6dwNUgqeO7y4YeWM9B2w
yJs9mslo+7mwPnnrsntUQOF5iWjoRpFU0cUR9Id2PEQlBnWypy9fvZAGQegiFR1r
dnsiyg/S7Zr6QnPwXxl3EIFeO0SPuy/3k5jVql/F5zRmYbZsHCschkVsdKvNGgIM
GxJ9djxJO3wyKeRFQtCYioJzhFM0bGLd4zOOTid2B/fVUjWZS7QwAsPK9fhgDMgQ
6sebEbEr8ZSw4tRza9kuNKMtzAQyxFixSqXAi2twWUXpn/JyBt+VV+WeEYsgzdjE
cizVLy9Bz0T85tXD/GqxrCYQ3/Wrkddd/vGZ47dm+3WY94JcdeRCk84vXrH4szOu
QVjjFkuVJCpY9iV7KGN6jzE2EqFz3MJrfWncnV8sq7GJu822H6QMeQ0sPC48qa2b
RLaPZbcjs5xZAvowgMcFaKVezchLunI54fq98pryEAPEEm5DhiKUbRl+aKSbH8/L
9F8S9WZK7ohnXWxBgdkMyHD4cokthFNqvWNy9g+Og4jYLuqHif8kVxnJPdIqzA15
WmcYEc11uwoElfaFBze5ahnNMCDS4UI05OMa1PLFKY0OQjg9YDS7HSC4gHbgQQkL
pAczFgy2C0GTh8No3UHpwrNUqRCdTVdNThSsWnnAOAPvo39gFPPNtCqVZPwkAlmK
E7QwQh3/w9qedGZ25/S3w6PKsvaAQop4vFIMjnxTAfuxC5Nq7KpAUGbLlq4BcYyi
VH6hjMnKUAIW6+Og4F2Opgp9G08hZFuSqROo/aXkFy8uuB+qX0TQfTP7FQcIR3Vi
np1gDwXZq/VxscKXAKCoxfVhA1pFMWR/McBjl5kiCHRi42SItfkSewzgYGfkOh7M
4A+3F5ZFApsVYXjG9I/HGHjWwHgJ2lMy1yzetYsS/bLcFLiseGnGp0wIUzaPnNDN
sR/rHPRMxsCM0s0mBsl8RoiqzN/lBbH75DIq5YxBahqP+YjwPKCaIPf+yHgzFJty
KrxZtXQkxR57DDEWr1WI7fgdLO8qUFzdfdneOtvQOhqP9uvfrPWkyHlt8LaX97/Y
C6UAmW+4nMcUBYHS/1fxGTy0s/jbKwmuXZE0JvrTcirBcJNFHZ0NJXZiMQgxEyqE
HzOaoqSOv/dy3GI+JMnBRrZUlpwjWcz5TVXzTd8DdQJto3THKtSOgJ5CvjWf5cJz
9eoV2109ulJP4pSdv8w0zrWXHZsy1vRGc/SBCmOl+fVQr3YMOz3aH6H+KqWrHvl4
htxKZBTK0WXGfwQMizAZ8PwXj1PnjQdmybjZLEuoB+DQpD4mrKbfp/02MPWGyjfp
FhCF+f9xR6g5YZmAdnnaKvja2kojoiewi4yEu1MEgs53bdPJqfcj3/AsUvHBENK8
UMF3glVpnQbMfcpqAKYMARM5B1Nd/nm00u9Y5touC5njg8CRlsDRWazE5QAQf5cq
hNDtrvtRna0tFaIO1UN3MRvaAj5acfQYpErrU6CSrldCx6Dbn7pN/hK05py0YQtE
AcaAZYH/42sz68SD6G680te6rWl5FbMgJoZq5Mk07EXdIHzV20PEhWgex+Qt0+pv
3EifRlWtAInVbZwjc02W6r2YGUzwEedaitaG9PVo8CIAD7nsMwuhNpmLsnHDgPDF
TOD8ptDS/VGcaHvLnvhWufZbUwcATjCAluVCaR2JjCzT3SJoK5PNcjAElkMvoQjl
1xSTrzYifPNRWAIaFhih37C5CqGFG4n3Vn0QVZOpIJWw4TqNonfmE69Er/HtPUfv
Muhi+yCaS8lhgNSd8hJaWSZf922aA4nyzoHjTOOefc7c5y1npvo0uV7HFjPnFEVe
VZXGtTnRiPKsjXdfO8bNvA7uvmH2JMvkAzo26y2wX32KWcjOm0QtJ/IiSVkxQj7v
Z3GycJ3nuztJjD6pU4k0J9GEEgzHMdpZhjrNBdTMxOM1330YN9uSTCjDUZ6PVz+r
RUEqLn0ViKh5p9jXNs62uZSHVlLQ4jJ3Hrd/amcal3aOMO1T54e2BP/lVK5TL87d
yOrFGCfq/mpX7u+LvfTAShGv6EowSdpiaMEizhtviRPW1O/dStDGwBOC6qxMfBHt
1Kjg56YDIV8vgaoY/bDwqTHnLdV0JPbbOm2zNpNTQQ97wyStNcRwsEekPh95oKr3
/gp0EKRwG7GgJQWF2T5oxQp2a2udNOM1kn5E8WxYZx8gyqITGiXBWUUyGFfwNaOg
AFottB8cf8PQgj442AfNVfm7kl9lEVifB5tQr5bKIg7b2PpeBSPS3M36X2V4sYfq
HegFB7Cv27cdf5uRN2AvdIi0GqgnZdGItVwlO9hclP0CNoNxXhGfTCfKEHRcjofK
mM6+L1/rlej9ddPPD+imlb5pBw5kVf9wwHFZWSqdh20lBIAWwb2nrwjxYfvWqvN6
xkr1o6BAdHI2q6m65kVwGgxvWv1d92DXhBwAN8aFD1gfzFCm9MRYW8GaKcOme5rX
fUX/YvKmsMdibagZ6AOI/VZDpXVjk8BmjJ1SYqdG31BED+GzNcC3UKReETFfbELN
3lTqwORr/yFD+NdKMq6d8JhiHln86BJIbOskRjTzEdTqtdv6ho48XlmYo8SB+6PJ
AhFJDuVD1eDOQ5OYnR4reH4z6pFbjUNJfrvAhKBp3Las7KWXiQIH4RM6xI52275R
CCrUXCYzrYif5tX4cEskjsJJ9/fYwO/UTlbzeaXpqyA2v/85/hBthLqZFboFfQvu
YBKUdM9CldFpYnv4RLO/zESSxhz0cQ2wuEn87/6ZHgrQva1iZalESsNEso8DiuRJ
NbLjUOmTTDoOz6qTu/c6P0WccyKwU5yzMAw4Ud+5td8T+5cKhr1J3jywjfj4BRFN
DOr4JXcwB/0tggk/1wEsV4XUiTGdUdLhnvem5rBJnqTRXGFuXKbNo9rplY2QzT6t
xKQ7snZEEW8KtykY4q8VeeSz9U0lO4+FXdkZ0arBYUJGQjaEXO8ZnTcxAJWnMKJQ
DrEQDJY+s8dPt3gwJLY2JgmJqjDM6DWuksF/8QecDwsPPhiFz8Nb9gVlWStWzoYs
/01zC7Fq/7/bpBm0tndCNhOTdgXcm/jdmnASwKMK6pgaWkw1ntyi6gGTZDSFI30P
k6bmq7edv2sO8K6ghbvCqOqvx8Vvm8scQ10gy1nYEjLUlFTwq+ALrph8WzFQJ7JJ
67ot+3SrnqcR8Wwcp3i8tspLUt/g4wflrrFe0w50SCNNSZd3w7ahwfZkbEDC8avi
un5+9611GIFH+ujxmIqvSr5BsXczi/kYSOn+cAMhZD+59KzDIzj23zXtxgoxVSsU
IDFJPw+IOkm70A/Dm2cH7O+W63i9OjARoOIqxlKc6D8sGWw8ixENL1MyTAs3UEy3
V7embUNRmRVM0xT/VrDjtUtq2YXg5uiU9rlT1FUc41nxaB4bsigvID5YUgT9LzEG
IEAsX/40WtoqxOa+F6IuJgkoo9pXLp0UGDAuRMyv4q2PD1Jjh4gF/wXaY84vYN5g
hJkjTH6s4OYhtUx1ZI4LVuZ/gQa1hve+EfyYC0dkY8Zof8g4z01h9gvKVlFbD+cP
jNg4dD8FWddmXElo981h6NWbLDfjPdlde2mXAem4tMe2B0YeLK6UlYJ0CfehVoUx
Vc1gNI/vyN+4ge3BjH50caRP8kDxDahDcpD9EM2IHDcvjsRyToqIJqoA2QFm6Hrh
7yVlz637kDAGsMZac8uR/wGVMYcjxd8gKvj+U32HTOcFFY2ELPzMVRl1c7Cac+Db
RmI9l0korQj0Egdbwicfq4vTiYDoX3x1FDR7g6EVhppjTNR9XU+350+m/InXGUwy
xFSHHbYNQLcoWhg7bTZUWVBL9biTEscpxYz0PatHN4Q2rgYu6rg5Smvm0D7nBA90
/PkCnRzGq37oOEqPxC169NBZmVpE9DX/m2kWbXyQskU3kLEi+yvmvu6ZlZXKZ3kB
Y+TOOUHKx2UnXUEcuDiOeToASWmYj0b0mPT9desbm0ypmV2/ODA7YS62G0sUVj3I
cVndiH+ENrI8oqxhmrY2PU5WJ2GKtEjslw6HskxYoCFHXgt6lZUDq7RmJ8gVJ1q0
BsC37pwPCQB0b3TroNzKI8Hz13KesPSd6g5a5Br4KkHygKm6kz3Y4J+dU3VRn6HX
v3NuB/0ulaB3oQiij8hnPVl+zn76xe5lMPQVIXPr7nJhIXqgqUJbc1ktO9dCy5aG
fh5H/x6v7bWBgTTXOmNDp8UN4BRz+dhmXYSoF4eyow6YR8TrkvqwErcHlifdiuQY
+q8qMl0I6TvXsqcWsN4CVoQyx+cx4YWshnGVZrLgYr6fzAowxbY66buBjkZHqG3G
csjyZN2Mi72b2QmPXPqTK3ACXQyddPExgj+PbxVqlcr4/8B7YAa5teZJOTog7jD4
bZtWIvxnVOZeFwF9Bh5oX4PKCUV1DqDgSesqsvA60DY/Zhj3OoOZptuwDJa/9pZT
Y89E+0cq7fiNk7dlQt8Yi5+CkSSCRZKj1seYLv73vZQC7g34HPo4wYcvjoAbndP/
zZ5K0EAmQ7CSkgMHosdHCGd8ABp0eAH8ED69qJI5VWy9h1r79MQgfXSTXfrUoNNR
3sSd1r1t2AnSbp2Nq4jzFHClIEltNXgW1/tk27SnfDCVigIyRik7I3DXt7xQBMXy
IU8JfqQLjorw9ukmbmOXwKfozJNXsmsYGFUt9i64DJBAV5X3OIG+2SJV/SOAuC7D
UTA7FgmIBwLDh+x/py4wgjjx0nZ7DDKjXaEp3G4HbMFGry74aPA/Jnf5gaHKh0UE
nC9jTmJimyp7G3RDnSNXtn3tWSxADf3utXXP1Eam4sd1TS0xrbrqFlgiXosaHmVL
AycsyebtdYI+RbQvhRxvEYJFthOpjSfEglixHR8BwLy62If57No5bwvVPCKpPH6z
giwzshrHZyMgdBwQyARudWVVnkFt5PoLZt50aXIO6sXoXiu2Yd6BK9YxFQBUS6sy
XBZ094Q4Xp7C31opyMbXuYq2Dc1yT/JhbpNkVwuq/coLxA2tw5mDGYwslCCbqfcC
QyHIYemuWYgeuR8gtTbXQcKTLAbEfSuQck4WQ6eJ3ZPfw8W1/rMG2jaL8nvCJkOG
PP1ZDERwpoAAzeja0fwF97aLKzOl/RoG2PQ7ZSaaNaHZpRzFU/hWjuVl+ovUlyXY
LicNcvnNozVGSnuKzQiuBDuOEjalpwKexsbasiAOwIXJnCIwGA7sj3HlAHJgBmQy
NvEsdjCzKINxFhg+7Wbm+F8ko8nUQkqcoUpX6hCFHLUfbnZRC06/KPbw+wzTJ0w1
HG+esYrEzcwfxaiDppCP27eX2cEhlV+7DV+Dpr5FuJse/te+NAwMVD32QgENo+6r
bN9YZtQFNkbpQUpiU/NTKn7XPOTj5Y7/lNDB1ZJtgwthl+9uToitc7NAjugakWdo
kBDPW/x8toV8ZgDD/GaypwH4sTv+jN6u2nYGOK7ihur4uFvCupaXPscvCzIlUyUd
vniUjimlMs4PDhbMvr0xr42ga8mDzRF1dmbfONNejCnCr+OhBXYBJQRMKKevgeH1
sqX9QdkVohD64MusY47jLswPFHOrnE+o2g6Rwjdvplgfknle1NrZXbOqhZl82FUe
csE6sSQwuZHYTM4QAESZN+SsVQZvkZUWrRF3/AKILbEFl0a+ckukyhmKBoXZDD06
4Oj3DwFbyAPminyhxdEmhAhO2zOPvEo4Y/Nm5WcCeClvVtWNAB77qde3KzjCX4eR
nuGAo0ELx9APgEZvPutupdvwNkGKQAzIQwWIQe4+2AxiXk8ptFg6qkOOk+Voxwcs
xN9KjNDaSXT6pfTdA516V0da+OULWe9jTYEk/EWP3GMx8shEc95KKiTk16hnH7YB
OC/XODnogHG+WqOaeQQm/FNw8mSmVee7CUkAQGjrpEm/s31WWaDxUUTHVLW8hJbR
UQVENkMmSJWp64Liy9OuD7bPsW4rhIgt+HnK6+2KqF+ctEj6lIMJ+St7qvvsuWRF
YWznNIcN9nU8pnk4pfRGvqXoFf33sePPaMjipcH9AL/hwbFNnEPAi1aOux1HkmpL
T/P/FBOEzkGf/2reQfysTRwH4omuzqM9hMeSZZE/V2QVwptxl0rLFBAdvEZXm2ij
C0bQGS35X6S9vp0qg5ic4HOGIZyo3Dpfj/PFCojeptc9kgSnYVryIlSOr8KkYHmm
WksCOw/Ybirmx0+00SXvr7QHDdYNL15CSkbZmqbUELX377qkl0fHxEUxwXnTGXLB
ZbOCtYs9WpyTRD2U0DUWVRJ6w6NXlYlCfceTR6fJY3AQXwejIUjDIejg1/uk1bHH
yyKrGEshj0FLTzk7hMcd2DM6uUAhlxa2B3RNtx7A5oVVCwgeJ1Zl5GvBeV1mz7MH
6z74Vy1Q0jz/sDxqf/WD5dxYYWBJGXfPY/tgpuTJgZ5pkArOVTNlT1Ryu/CW+6HV
Zp1kw7kLt1vVdjTRPn7S/yKHJMj5I2Z2uSiGLugMuT64j7o8NHl1LOJhetiYzBoq
JvNiXr9WTkwJA+i7XAoA2YCtAcstshbOLqgEUTMewSnQdC5BXDZCpKfZ0Lt3ZGob
Hub2UVNHhWfRa6JdU83Hqg6Xqj/mssIt01BF83tS4x8d0AlJl+91Iiq42kn9nJ0W
SqZCaRg4A48meIo0LfVtzv0fwkMg56POYasQQ9q+Mv/Q6yOCEfbYKFA2z4kvtr3Y
PNkb3Wym8AcuS+UM2DgWny+FvMKH19ahO19hm6tLWG7YdxA8E+W+idM0dUFRXcyW
G3kZmuIG0U1C2sVOQNh/01AONzr0poctw6vQlFe9oeJN1R4O7HWTvdWhXIcu3zhh
gkkbzYzhTOmbSlSTURF3P0bugAvbB8Fu0LOezbIQEg1g2iar+sVdENt4l3zMINiw
tNqZ52LE1k8CrM5HvmEGQrdDuTIZSpakz4rkQ3sQb6LU2LThx3nOr57LYoehAPSE
RPzrca19SWzIvU/l32LFu4qVvJxQ1hrjHLd1sQ5Td4Vz4WOAwPSr0su6DR6A5WCZ
zRgMa2cggmMoE5yk419xcXX7UT5EYSndIDOcVweP4WwRsIQZrNJFQ+mbLeMlxNmV
xFr1Uf/vCpUqXnHbtt+ZblfZ40F3Qv3guz+yP7LoAK9/2HWRq22EfeTq8Rs8aVi0
WYTFKaBrR8vM2nw1nS7keM7+tzxYTRWr44IVzoPYf8W6KaGJbDyv96LIxFCkizsC
vcfC8kxcFL/upgJsJ3ggVY2w6fMh4OhY6tNNIo/DjzeffIptAlUYaoB1LjY/W6ci
kTKbWmAMuL2yPsnwxzjqG0dR+VeLOh4D1dTDjVOwb+i6Cz8qPQqNJGGLVVsC14K4
kLOQfvjRIK7UXXK/Gnq30Oj3w2CmmEu5+uyfHaEnt7K4KYiDioCgWKSEWIiFaxhn
CcuOdFnZd4g0x5elWjaRFlow2TVLmjIHFmoUFbQKeZ7TmQZGAza7ZZfncFHLaoGR
7uI5pShJTqAFs2ni1ZYJk2pJZ+fssCJWbWPsuxgaLAWQMxL3MhxTricPFXoBoW8f
/xceC4c1mxSWphW/7TisG7IluuWcjA2AWxMXNMcYtFGCIJL5Obdg5fw4uavuWIk3
vJZBKcyXHj/qtLgb3NLMpwlDvXPWdw+JXI7NL05dzCioBL5aXk3v5wPbSScXIhr/
JQjgZNHnFRvBi1ewRsFvVK25BohGJ8638ERWnINhSggX5LrrOYpxBV7DpD3wpgNO
CGkOD+3Ru1u2UFFDwlbuzXdG9SmruDvRS0rfQ7XGe9s2uk/LVsUhAQuhb5To4QPS
eNBobyePF0S3hIHHB/WYGwWiZRrubQPjkkdVoDhWUJiw0x2YFARShsyC/3HMZWwP
CWdUdOJNueNqkgKMaev90e5ZrOmbH/VkLCKxinYxi8cyjS9cMIj0nApi4PX+YN/U
+aPPcscPIcUNQ2vG6biAkCCEbEVKyFOdw58+84WJQN156s12RZl+auvCtDZlclAg
EdvnREnfZWxlzaeQo/ml1vGrZCi0J8dY1bZHgExC/EbQ+hE/T8sjairZWu/1LYCh
8wHUAT3SMPKHKvPYickfDjjGoYKGxX/7UcEPLDTG1PoyPtaz28SuIydRIA7jqJq7
a1LV57YQFIdGDexdDfvEVyCyMDX0HApkv3rG844EIQwusm3x9Jh2KZ9jSZCQpPfh
/yCaNn/K6s1fTiyp7Pqqu6DZTFX6mUl+x4tQqwkvjF6M+IUR7ZS1MZkDB3xYcTgJ
E9/uKSE10sAER1DQbk4w9wyh2njPQjxmMvT+m3YtFqB10PYP3a5jztMzRdR5gVrW
3iIiS7ICCF5ZU4JCiIZpRWrAn2m8hOb6X3MXfS5ALNlqsFBBE9DhVzDjFIM3upHS
pWG5E6S9wA3laGU9zyAlMX1pLYm+M4i+sSxUuBHcD5w8OQGI8Wnc2rhiv5wADTXB
XYC6++gajDzXqEJNz/SwvianIbzeoNSmPDbxWMcjKH8QM9oiT/lVNBWBrSZI/nVS
I9K+j3a+5ovvvO/dPYCrx4dl52i7DlgT6QP0Obbg8D2XdhfPB+gf6wdSduq1t+2+
ZF2O9LxXbRVIxN0zHD/YcemJyg/WI7a9cdz3u+KLZJRPC1HF6ZxQgOzK51CH7hHI
E9eO6pLMi6M74ty3t6ngASNxYboUSKbdVaI3vyB2Hhxl0Jh6qj3XcAkre4Revhs7
zAkt0WhS5WSmddAnuMNztjXDY6sJuVJ14eZ93pUyxc1RNJFjp3jgEyBMYETCbhS8
hZxnN+nBKDn9bD1QXZN4kSPyouMKT0Ark+I656CKiZXx33S1QzTfhRVwo7vJux+g
PY+HxijpPVpZsn0a9oyiuekWwcXs/ZREfGKdFcDT51sBqG440nTOxpa8D51NU8mb
Yj3MjZuSuUwFeafFzmus/6b+20J9Xp19nKmAkCth8XniGZs2YXjQ8DzSTn034uC2
uqP2rcTJVbVwy2Gscvp4aJdL8cGJjD3WuNfTcQg/TcvBwK1xFLnmRQWokYWRhOwh
BC2yAd9DSSOq9enhcJMCJwNbUZJq4yiqfaQcC7yyZwXVMwZ/sVUqNx1PqHJTSAHD
1PU2zlqUUndPqWtqA/3OlMu6uJWBKVRWfbCc80+j649v+7IweV+2T26sz5tSH0NX
6wyj7dCyXE7RZp1zgArqO/PVv2sETm+vt5uO/Ln+uIV3eoTRy1TZKvMoB5ohzHCs
3gZ5qgJWSeiQ/a+m35bfN1qpqJna0uqKXRPg7Sp70o5d48M5KAyAlt6js6lXA9HG
3JA4M729bM0PVXSQMprtO26HwFjfhxwRzPjvQsCU9quret9HI7Uw5eJKqCNGC4nN
HGWU2z8M7cLeS0479XFjg3d31+BATpw6InorTGthGG1qID/ksTZIM9RD1y0JzCZF
qfl0v7b2YKCmPBCRI+ovppgpPyak98VKavwguo9Z7w0tH3Jaqx26C00Nwykrs0aR
SXhEM8uWCwbzzR4cXWgHJtBgA2QZZ7S8iFZXNwymDfO2lEXPGHfnHvwjCw5fovXI
11Pz8quC6yn4x88HafHDUWqowZdBtqx7VIs2/P83J8URVM/rP+WueeZCzbSkrdnB
TcZUnaosXVmjBlUl7hbHCJbIhkvaCQMKDh3BK+w71BmQgz+HkjnfhzZp3qw9kHqz
V6n0qEsSPyr/7cOfbol4qF8Q/IchFA4ueXZIqKxe94zlujNIVGup3xI2Hf+Zv7OF
lMQ5CkIIsmHDI+hKuf+E+2nLl0F/VtLncaUlntcYLASHoQojKE1dOo8DnfSkYEiz
1n0gyqNJa7ZIryIorvJ1Io+S75OtFMSjQdV1yJJovbd4+xZXJKNiHZ/cOgfkao+j
ljOl9c2MQ3T258d6fwKwlOIp1zLefQdte267TQAuYh4E1FBeLzTkX1Zt1iQ/1v1P
RuITsxEz3pt4UVDMsIb2Adqk9G3uVNGD+Bq6RiK5T0Bt1C39/oLn6g8TYXLL3FhT
/aBcLSd89UMYoMJyQ0M0KZqH3mDfjLmQpzd0vKJ2z1AV9hdbdczyT2nyOmNDluBu
6VUIcHd/zGfYy1CoHG3zIScJXiGBOfo91I5YjqkM5pOIlq+7giTmfToX/8nYK4PT
cfj5Tb/CMoHz6JNnukZFAHbBi421+oddJBRAQfMnOx01KSENi17Ll0tG7JXjxjTv
lc3pLguZmYSU5XkOBO+ThGZ8jztTt2RemZFeo/hu7/E+IBl7NzAZfh5svYqY1AAw
OSAC4KhLmrSFsWzW2qiNi59Q7FpWNTvscKp+y2DGRXrlBr7nyLeNlnI/hEQHEdsC
1XhD5MR2PUbALDn+8hEUMYA+eAw41QQ/+P5uFq8JtdWv2HQLJzYDqX+ONFnqvXxw
JCyD0Q7dhmh1hrWXjwmn1nBCtO6aEY8aBM2BikzjDvyH2R0ha+7WKdLLivmit6gr
B4W4UxPgkdEP7WXTuFk0tbPrVGRTXMIQJR6qsWl4H5rddO9F1nPhh85pyv6XKh/f
o0zwNIRIlGqTYz83ae6ShG9txL1z3OCHQA3rMSa74TydvLfsRmmEleYbUIVJsrDW
emJ95FQlFWBRMkYN97a85IvO3nzyypFKRIvW6vpT7h4OCXuLqy/M5XMJDGTAE23n
fR6ltbOlpQVt8m4DWZLD2LSGC/E3bvuzbTcCyUjtjRRj9i+acZr+6w2pbRzpirN1
2M1J9psvxlAJV5+WVDCdUvGHszAa+7P5ARHroCH95mPCSks+9ayA+jDRm380trU7
ZhWNRElo3fjOfaq1sv2h5VuX+bkgFxDS3DdQ+Al2qITq+Q6NNZ3zTBE8Es3wKgNa
xrB23GAw/+k1HdrhfUBnC1CY1yXKUbjB/d6vMQbMksYKC3h+23moo0zAIqgeBg7+
wW5XkJCES4BaZRqgPTVL7KPuv92v19bPc9XlVXJSGPdEhxECqCkYrwJRIwjUSfwU
NGR8lpm6NkZTlJmf1P7df59fFHpV3I0NDInmfovsEumfn3GiOuExeZk2TUcztNw1
TeR752s40NS4UWEkOzTnWW9t3DY1DslRTn3BzQk9nSEcIMBPNHqbnWCeGMp2fC3F
3zCkS3/QWEL1sxTijYHke1UWnNwOjKfEtv6YwAU9zZy++fMJlD+3VulGPpXtoTTs
CGpnc9MnK9mJNR8x79B3APOI2rjEeXziH9ITC3v3UEPts36aqp+h+A9FJw5PlnjI
PM/epZo5qNuhn4f7gcq+S2F4+yVnoIkHkDTTZXEy87SYla/gyolKTKCA8O/28Qaz
N8tiu5E5H8q8c4hC+u2fsb6NwA63CHS/KQ1L9bLu48wOkF5G1EiIONHu40E78EV9
hGG8gTik6q3G96u6KaDdZaQ9CAZq896cekJ6wLsogSQ6Y7GHe7Ywjh+ta/3qsAzA
XipWTO6zYaa2SEzF8PMxMDq4jcZ7hMrMX2K2nY+dhytWgQ74jsPn0xUKNJwPoQMa
4nqCEdMYn26dXxs6nqeZ7/geCwTJTnWsLJxQsDxyIBDVeaa9Qw3CcIyojZC/QVu0
Xai/j+n/5nWhQdnQUCTykx+11xnWu8WMOtPOXvFsxnW/FmkrEY6GPKe5dX1Qi9EI
l65uNwTJZ9mAqB+tmNHDVcro/WlQcRVX4QQmGFBgqRyw6c6uDNQ/SMl0bEq3zKAB
e9BTiLqMOltWqX6IbbFuFY2wTU0ca5jYRH2i/gZ7mhXCiYgoZFhoy6POanOZ7/eC
HJK78maVA76BIp/IRS4LNONstkBxKdVn/I9r7/k+2cBsm6zj4X1x/NZEDof9KdSM
YkgBqToUucy0QfmVCQ8m3OHNJhb9lTagiNv+NeklEwhA2b9MtCNRwlF2MRMdRFG6
XyyWgOO1/87l5nos9s/wKG73BHWwerNdPruxq2uo1JCEulxNtBE9O+Xfg7kmtENp
e0/CilY0Jrtjsyi0eA80m6USTSK+p5ZiI/AcMMCJLL5vPR1IjgnGHGjVhW6RWJ72
obgHxG9VtcLh0RUk1xJdT7a9AfOHMyCPII+iyHaZFX6B6GNUozCLANZRbBuIrPyk
jb6jlXcI8vkuKpScG2+3guIxpqJq0SuLEcJ7mvTdxUu7bygGs2/agpaKKOpzhlft
eHs7s5Od815TNsSDLfPXxSk118u7JRKQkqhj9AjwRbidqQm+J/mlHkF8gz/BVWgr
I8nWyE549sX2lDjAs3i+f/LlgDgSBA2AMnCri3NHCK0NKRd/nsYOfTBLwAJs8vTC
oT5JK/RrFijTR7UkFuBZA729cK/D89lDm+ziUL6d1mFzxX3otn8fkE+R0VGHaTwx
hkolTAE1y25hl6lBc4vHAx7gXZ059+iSZV0sLKDuVtOl7+dbo38Uzt7/tJ98rA8k
bx752R9s+20BvYH8shKzv3gO+y1AVTE8nOJu7PmInuzyIMMzTX4eggAXAtquYocH
Z3acEh4xdszMKXAdcK5tCHMMsRKwq44LPY+ck1us/zZHZraLu0M3h/g26gDLDkmy
d+WC9fLL/dS3FSDGh+oyLkq9TJVZcWzNQxFZgvV/H+SUE22ijjEnEN5ojJZGRTUa
hlsWesvPSgiREHQz1TJ2pp2vdLBWs3Xo3b+D/7NKODcSxKa21IgRw12l9cHbksyL
sQQTeK9ulAxUVpND4BFclRPBxbsm+ce2u5B6uuJT1ncalLXcemkYxN+50QhBr2Pl
4BXRySiymtzAVP+YM1lPmWUoGsYvZecyd8Xm8GmsqxOTrbXMTCV7fbmc48aUDiD+
tKGRCDupWRf8MzYPfawStcU9Zcv2XUoVG7v4TaQCLmibxYyFghHwFZDx4yD2h5xC
LkMXXb0xZhf/qbYYub1Yew4MGR6V3YnLpUj5IJO5g/eT7Q62PgxQE2zjJWYnFvzf
5ZZWvZuYHaFGEzlXwYq15RRxgcuhBTJZnSC1hYbnOj3qPmkxEbPbTHTptoqmpXum
qoZs3KKyJCEO5WpjU3neYoG97Tg6Ww6rVVDuDAgk7x3Z4bGLEi+fDkqgWRaH/Y/c
glNelZwHOnrAN4G/gAR13BSiYdRS//pbcAsWCAGM06h3OIdbl0QhQr3QIIM8/eL1
Ou/niS8IcdSS7O8ZgbLG/odT7aBcMLoD2AppRtj0j7Ej8NgL9tcVdhe+MY/kv1Az
V3igdAhZVI3we06wK4dQ1QY4z5irThDIWxgD/9LTR7eFprEBE9G2bm8I0YeR1E48
JAlrOq417skJDlGta2iAeGT2lk4/iIaP5XD2LYiHqOu5M2OvYOZbNjjA1hf7EHkf
sRQTXF2rbAzanxBf4wJlKgwEk1vuA7/gvxl8sqOCctJI4iGg1niPfvbsyQ26JH7Q
+d0vZ1t7Qi6H0Vy2DeyYvEqXPmaFvsKDJ7OXujfmGlGNHZpGX5N2okT5tB/xwwcH
VBP/kENeYuFKNhwvL0ZlOXAvgfpwvUjCWp9Cu972VkKPeOZH7k3s/esxOlNTMaAh
IlK9wzh82nFMA+TmQgL7MdDW1pIEXMfsqHrd6K4LFEmjz2SBtyS0gvwwmnalcfDW
NXY992KUPzVuEGzRsU9rcomw0nmoujTNVtc2dIs+j7FJHBCKH/VsxwJtR8rcZj7h
gNWyPAi3BblJ4tpw00qS3YKjfZXA18KVZiNPdr3I+/xLr0E2fRBAs0ENV8/F0q0k
BUd8NxeoyUwqwfnMGjP1ySkJM1WLJS7Hw1gkV6CuhSxttb7Kmnd9vxFqo36xPHP/
UXwY2UzKe7dT3u8axLDLEmQB9rQVHJk0I7R0ZYolOYi//IgUs7TJyMLZQz2SVHoR
N20YWUL8WjKEZ2Zeq+agN+sfWUanqjPixc+Rpp6M5wjsUSnb+boDmUiqccANM1Zn
U+q2slyzm4KxwTBZtFpNzhKMPpM1S2hMCqtX2isJt8+wh0s18HLEfmajXmBoXlmN
MTKGZDIgoM/AWHxaJ/MNmXfpctsItV+QRbFC9+E31PudXMd8ZQtsvexSVZH4X4Ac
lz0rjzGjvxsD3ptJHd7NcZuXCqR9yZC9RM6H8UizKgmu7IMe0V7ROiSAvNqy2zXk
hNfMFQ6YozUTQSgAn/icJbcS4EX7FdELMv5Ooz6O9XGqulUpZQMPorn35nTgAOyJ
ZqAHS2jlgoxAIj0PtbY4EH+7Tli98C7dhq/FXzRSWvvxAJGT2cJnlmQwsbKFPiFz
GpAQpCNds6sp9jqSYkZBolO++EI7OerHnKjDyeqhGd0siYvomlhFjELNDH5OXbZr
7J20dCjPmZruvC2lKoY/NU02896eiozbgQwdkY7bqC2dXNT7qzlD5l6ySIY3pkvT
Q+P4vlEXyyVFKdCdeFOprCYsD6Y8lxEG5WzUT2fFN1j/Mur9h6UQtSFYaqufwgji
0pnrhZmqagLwxEFroJmlC4vcppOzdKUrDbjphCNxY4N9mcici1+uU/W19VCLMez8
/G2BIq70SWr/sr4CAY+2QXxsuKX9WBUFI64St0r34mck+Ue1K9YVCECqbzeJnxq6
OPDGkV51U4b4TKdiSszbCAe0NYFOvKdS+o4/YhnNEFYXiJG5omWUZdb/yr/gnfWD
Ntc8dAGks3Wxa7TFMoZ7NrlEhi0XlI3xDAWVlsWrpHYO74EkwrnclKmsbOUXSmts
pj1OSpKNvT7FlVM017VC3YtTrnrJpdk/WFJ9vXRXNud57hNOWS7TmceRl4iepfad
ihxNrNLmnV4XYmwkp9WTxPCElJugD+ScXihp/nP9OwMwlfb+nDWfdH/C703R+Ke7
1Ge3OJUBNT6vFd46KCwsXN3gCH/dVUQGzEU2MzAHqqPxoj/HA9uakBudlYUAa8W/
+S/ZOVayOHBZ6KF17LDd42PMuepacwjC7/XBzHLJ3CDUxxpMiSi9az2ZgTfH76mf
acFl/BqAlKygXPPIGapK+fK6TjZ59bwFuxEcbtV63WnoFy2c91+rlkX9lNcqd/ti
XY+t7HYqvel7kZknfJjn6FIoIQlMtt3zA/P8XHOLRvaWgST82+2EVMBVF7b3+fsv
YPeHjPPyb0W2mJDci9NXIv+CjiT4zGwxB4BmsqX0nhH7hCb26AhrEla93Gs2YMFu
+tD7oHOUFi2aQp53KdO6txgNn4P2R9oQDTSCdrgSTWUmnFCHg9Fqf7jYBSieaAHe
DCmMB5K48O+a4vRyobm07ml7SLdseBF7jFD0pLu2Mc3KawcrNYMGaSBBYsCI+ZRE
h+EX9xYIdsKGHFzAy0WV2cieyii/OKKZrcl2qj9MO/ZWFjXmLSHNpHZ+uIAqKCs9
kXjyowBSzYuibKymfOyouECeR3zGGTySxm/KoaN5o67449iepTkK0CBxkFlDorl8
meQ+SXZ4gQGXsbdu/91B8R4hEam7ZGPKXYJjzWgkrASSxtsVYxJ7GOmAVj2ocptC
54ZyKfXlaT0UaOQpShkEHks308zKuI35Zrb0yXnZFupHq/fjwAzhKvxdn+kZf/Bx
PCexqe5XcxgePcYFhG2kbE7qjl7Zg9EmiYM2obC/d06vCytipO1fqchpaEmkFxVA
D9RtY1H2IVGfHvwP700VFBhop3ejztjLrTcC/HxUYN73m1L5/9y1hWKLUIu64yHI
7mWB24FT0jB6lH9+ItEuCPhZS6nsuzq/Vq9EQsQQiboOvAE/9cy7VIat8QD+l1Yx
qyz1/mIeZsQrrb1DVha10bgngSjAcjh7x6oyFGBjCVyQNniXUSzA2qExQ3c8obqy
75boVfZByL/8bUHrBQSVVKNN52c34Su0kvCl8sIu6hlfn+R4GAxFfTgatf4qZA0P
RPgq9ZlXBWX6s15NyqVX3PcjJ5HBvzRgeWpV0Sr3c+Ts3gmfMAflu8qoMfAUZaV/
WWd7dNct58aSDwfvTx6E4tJIPJ96wL3HiuTNqb+e4+H5Nchr/Y6hXCabMqiybSL4
qw+mpjOreNGvnJp/kE/+rFRcH7dSRJXuTyg3K8bj7BmaXGBRwYT9XWWgRXHTgcS4
RusNovqWfvOW1ml42/DhvbmCtAUrKMQBKU6mIo+tUARU/Fhcf6kw0wVXMaRS0KuJ
d1J+YgS2lRrVjm6UGrQrTT8WXtiimsdh1X/EXuWfoVcprDxVybQYiviQHf/cRq2x
HEwDuzmYWNYgYNfhMPPwiTJcN04ck/xApf76nGh7vqyy1O8i649R10Nh/iQ6pCdr
CKtxTkXSnMCPCIgmmGmN3SAYboQMbRjC4XWVcN7AyV4ZjH+KLQ2k8TgFisV8Pnn/
y2NTYiodOFNf0iHBTwYmtz3QXuCAOBruQuPK5+HN8x9jlw8wPEzNUqJl7lZegx66
GJK8k8UOBMSdtG/nWgzegCUaa3j/SlaeARNHtBlDBHAr7FMJ5AqLZoLu4MC57hKF
XDYQQWGts62fDNTD7Rmn9q+u8ByW97vnC4/SgW+MqxAilZogRy7eShah1Z9gZdGc
OnO8Ldy5Od1qrtNWlHkAvW71sYqNXXiqasFa/UiLlmvM18egYDjJvcRkZIwzqGV6
kncGxey1fmy/6bQF8Htqg+jG0xD4m6Cc87iuukcL9k08lyrCLwPhvtMd+4Rv+cGR
xijBUCYb7N1v+lMKKnvKlc23N75oliitf2GOLEuQdskfXvicbuqHzRUs6iceWVzc
LRSqDQ7lX9n6RLGA2rpw6CqQ8QW2VmgrB2I+li6dSLMWPhYZ12mvAQMAlQygPhfK
DAvjl4SsEafxY92IsfYXPH88Vq04N064/NP2GmpbQi2zvsVLQW5Jg/oPNgWaSoQu
4MLKJRUIrCW/39GZ+9ua0fN0+/aKSMwmtEpmxu8HXluBCTpl+Ymn1CjVlQlJDUV5
52OqNfVEdzvNj01pTCDozyF+ahTuET3H0f24D/q4BWarPhKdB8w/UjQin2jHlP9m
6D/gVsHxfB7EUWKVyUKlL4O4IHBkRJ1XLoQpU8q2pvE1nwbwhVLhSDeERlVUjcyQ
8YgCtQqAGv9ncKGzaR/7V/MWn+i7DNhxVqV4qHdU5Mrbj6BBGnw85xrTElXP2OkX
tZBURY9FGislnM+owdpfW2Oq7duvtXb0ybB3gaFTr4zn9/g/XLT94mhjI0TWQnne
EP/gTtEgD/5cVqEThJde4N99i8AYG+ZV2zKz1FmIm541XkB6GMPNuGqby8R8pU01
kYeXR8c8MU6gY0vPVK6rD0vWjCTN9hra+A+nOqbsGBUO9wCudF503eeRms96m3LY
/QO6tND9aIqD/80m6L9CqXvb5z+t6gIzW5DqpTXJQX7v/rBEngtvP2A96ZrvA9kk
jXSj4vGqLt0GWRVMshvsO0mOY112wPDncbXrUGUV5We88lE/1G0ijzNzcx/SX3Ou
Beyh+r9tpVpLbh7p7nOXfQNM3PS/dTLpVMh9bqpEUp4GzxFJLpkdhIPxHHBP0q2I
bvwlxYjbWxnZvhbtTytTYeLwdD1pFmDFaRHEzHj8APnv4WdGhoFNfWYlbM5oiWkE
MAUD6Go/RMxOFOonUhxOXYXGVIiSEpDUF3w9dynNpZIBQzR1868myqhPdLbD570D
vHIDvWDaOsi2DwCu4RjWzOpwnW+U7VpVV/hWZO+9fGOKf8xJefsikpet+5zAeD4d
x/Sl1FyosrimLwaAUcVidWKYrrfw/74SiUvHFmZyRNRMIU9guvJ+1jtTCsyFb5ZH
Jy7bI4blDz0Bj17UY41+tOqQGRkqv7x5oEQ3OEC9OsSbdeLZ9Un9JSnw9cMRWzpI
707bYiU+LheHZ79lOYwOYf+PI4SrXuDwnbmNof8NkVzRO95vIP27rjWc1cqUo1DS
H/Yriel7zPxhPC88FN8fTDpseVuKCwNB74ZcLCTmy2X9V2opNTCpKGC+nfenU3Jf
o3vhazqWI5PWrVw/ADqHKqJq+zt/QoL9hbZqdio9eZg=
`pragma protect end_protected
