// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TyTtZSZq6Lca2ZetOYRCCw3mu0BAivuT1H6rBK0R+7enusQZgbLjojjxKYyDWA7E
67NKIHHO5sQeQuYAsHeFp//2HDKr15Pw9y9LbqjG4LUwH2eMLJYqVMSgm6jhMCIC
g8rgxm7ST/euh577g22idyVvJU5n5c+kNYVe5jYk6xY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11472)
XuK2EP/G3cwNazhMImFcIFyyhhuFo35f1oEi7lm1P1qBYJOcWrZ5x7fWjQXOKdHz
beYc81ufleVWytosBcrV5Staelm9rAuhlqMzt7ltcnoe2HrkWj/lkuezRRErsX47
YtGR1cyRpJPaQ1F24HP116+Ym4IUwqIrEhu+TCBbfRcohk15yES2Uklh1VaDf0ey
Cxhmf456Nk5rdetj2OAq+C0QeLAOxA0FmX2YwMKXClJVTiqSXPtyB4LefSmGD7sd
zWQ4RQlKU/US1ObD5f61L7kDzegriuxymbstlGyX7jeH08IM4DWlS+pnQOAS68aZ
z7UQFAiLxm8iIr0IJe3jTj1lpY2Q/xRdk2aiwGYFz+DfdWcXo7cKfkioBsTOpE2C
utMmc7G93xavtGwWVltk0SfTHYoNUQOdej9zY69PN2Y4iuLXdB+lwpI5rS0+qBo8
mV73HAWgkoMVDa658JNIRtdTJfNSCNJjc+mhcrEa6Z9UkR4ojTKWdCFizyE4HCmb
Q8SV8k7TPdAf5Rr2nKWM7E/MUTt7PL4XROuSMfT5ZFDmhEFmmq/TTeUtslcc3C9E
2GYYb/DiNDnEiKu0Q6jGk9BXqIxgJbLaaOiw1R7T/U40uyOHiMIb60MWT+9w8Yar
tdXI8pDgshBOv+EJ66siledyTlVPQ8xF7ne4/yMA53nHbDp6CpXw31fCR93kpTgZ
9WhirIBux1Ri0CoBUIWfddHjaVx80t9qkeCpd4FLwiOMoa/Hu7KNbueS5MsGghjb
j0eTHoYt3AamnxsnJOmRkjfrZOwszhWxavw2bxqDR9ggLF5VsjPJ6Hed+dRXE3yK
bK+4Jrr54op3phdHWiGRfMPeTTRIAwd51iAN5hI3Lcbs6Bbseawtx+goukyjgXad
q3mQvd897bIgvneiLJC0JPSfnp2rrjw1oMIB64BnyBUZKWRDVozATSx6qepDMWs0
IyuhyWntET34WLh4uUqcyugjmZ7P+Q4Z1+aZFsddMxEHEdjwdOpAdo6NOHkkXqLG
dRv1N/cKOSP9/3C+m3m/ABVUdcl6fKLbVg7N9vd4gAAVF4r+aAOnGh9kbg6ttABm
tqr3TjgV5X8pGkkdRzzWoWVi3VovVxVFuI8w0P7D9mw7UsS7nFdDrAj07PJMgyep
g7U2qT8I4JvBtk7KBx1udZlqxQrl3GXD3hyUGPfOXT68sasFHBWK18ycetf3J3zp
mElcLH6Ubt4uNxs5rRb/ijJrhPSSX6om6VeozeZRjQHpDSrT/SsaCxVMyTzyOeDG
PcF0NqctwMYcxAo2QAWxef2amGLCt3CggvXAnd+NR4Bjwedi1vfDFEl9D2P7W6nf
EjU/AkEp3qIfZ5VD60UTsS0ea37kge6rpMqFR0B6NpWATnwP6CtMFRTIquszM5yZ
Kn0jRT5yGh+nU+Myc4r1hQE3lVjYaYFFNaX1bEDCr2PLWAjT3oDX17JjJTCsWAw8
XiuWcv3dk5N4lMostVs29KYx/LnbTupVPmSirM+Uhdr6n+QvHNmJuTP1IDyL/9je
UGYsd0EquQSFZb2C0E0w8EhvIymK2nUi7BNWtlFmVGXCdsTzmDyjilBcxQZb/qCP
pJwWlriB5updmw1FGomscWNSMwhVRbTiYx1WhpoOYQZ2BICi7vRtcM5Re4SPtpkl
tc8CY7/jo6CELEraPt2h5vsUF6sjCCZodIstAOJMDnHU59FDqixa3ex26gS3YDra
njwx7Po7WjNAgjDYA1THmJPUupD0KKp/RJurVCThRcH/byQhyFDKgUt1f7SBoAUz
cH0k8R5xl/RqJeKTfIHuqjLDzFquwpPMz6V/iYyZGYzE3uOh/8/B3L7ir00l1wTE
29Ui8jST//PwRCc6I/YuO1Qg8Ngo50f3mhPJBSgduDrHcmMlUvJJd9PPFfm6Ibi/
0d/uvYosaUeLAXmVgtUiy9+ADEquBq2lUhu1UUlFwWmX4jtpIKnTzm8ViH327B+O
Mj8AeC5yFXmqke1g3fm1EumWjpB8sRhhSgDh8wbV99bF9Vl9qo9WwFAOb0SDKasX
eMrQIyPrz6ibTqWeX7QDRyzYaYXfGj8eHwnsuWoNlE5kNRpUfuHfUqJE/KKydFy0
maaltZ/lF06iUkwaVjc1WJEZwQ3xGSM2M1SP7WWGmcEHryp8+IhJBejDKEpVCRff
6QQHx4R8EnqIWnn+uS4/p4B0NEc9YIRA2i6QS0gJPlE9xdsYPnu3Jh8nmHH+wXGc
MEUAXgnaapU8ZDF5GmGwnQWWU7G1JTemJRbiLxx5Loja6ZlnbaYoEBUmqG0av5MC
gC3EwqFYwzjlHLY05owoI7q44r7dsyuEH3wRu6sZstRekBt5TTJs/ZvS4yxfBKVS
BJs+vKco9bGAFJFxSRb06btruYcKwGV6ziT3r+fOujf6q//1ndtI6oFKrWzrzdQC
9nlQr5ytbVB/aHn/fJteTaeeO23vl3LcgtP6+woCjnxk8Ru09CvGCmw8iKDfOTy/
bNX5e1Ups7z1IpZz7/vYQ1fDUsEmfLsnhQiAmgDspASDBbAizj7YL2WMCJr71b2L
ZOARm/29T2vNMCG8yKCL+ln9eiSc1WO9mHgyMUvjnEIOh6WSCt0JNYNUIBBDxroA
gUC5rlCfr5AW1spgjcnfEMtyhmkLKtZd0gu7IFEAWnSeLNR4DWZGinAWfW7btVH1
CwY22Bn71wUGCYB8WeeGJ5vuZ8QQR9EduKUerA3RNO3ilqxNnHuT2Stz8K+9JXUH
hlZeJBDc9D8aOB0dTHyhVp8VECi8Sfx2reyzNCmw5DopGjX/z5ipCq2+WXvvnPF3
fDGN3mZOApfdRdP8bXTV/v8DhtHnDZk4pQXp+QC66KKjzZkiXdpXwe+sJpgUlDYC
yMtnD7AV8sBzvCtCDiCVZu8XFf0uXsk9kLVVMo4CMxsfgJu2dHq2q1st2GSDCYC2
WZycorR2KMVB6ZB1dGK2ZK27FVSoJRCIuhIrVmb+5Cr5/smcHv+jg2sAX8rVwk0p
md1DutBHW2r8b9kKygMaPO3doVk4+9UyqSQJH21282JssWS7xJlOis6eTn1z4mFZ
yTPcepPcEoSU3pe+KwX8zWqWL7mEWdJ13DTvy74KpQ6Q9559vKWh5bNpfeC1HBC8
1i/UMy5BMle2whNSvIlZiwpJOenDBA0iJYtj6QeLwz8bAxTcayrjbdcI+X9mlcUo
qnucEEKtJU4koq9TvoV6tS1XOkrgv08iNuVPnupaG19/nSpBjlrk84ql7FLwkge4
kKyDLluTIEr7ZhT+QLzKa1C7dAvhd/r62X+uMSQ0fKL9Tnm49PhpVgXYUSYLfxYo
8YhPKZzQuj0XUu3J0Fsp6D8ql03FSpl3VqF5554/sr+4+syX6bLlXq3PFp3NEs2K
vYpUgjwFldl2ROSANitjuBKiHAY5CE3RyLy1Jxqa2uz4irirF3t8gNSwWVLbhOuV
olHVM/PTxWgF4A9bsWMitejg6ar/9Wi+VChZOFiJeck1RWUAKYpifCLqUbkozvYP
PmO1cwTotxhoXSysNLAPXHyhvtv26h5+MYMEYte5xBGQRFkimbls/Jo26ET+/S6e
/SxKUmPJzhAxRzX9mKSxuGAZ6OgFNMW5dqzG/rPClWHRmcHgECIn+vXzOp1W7XtE
SIxSvvOfHE0/0QD/SOzduutGeb1hTZbH7pubO+eOIeWj2wDpK4n3V58RNSwNRVVZ
52iEBeQh4UN6BaNecDx580Lq0jLQH5YoqX8O1x5RUdQW+d5Q8YvGbbwAaJpl1FZ7
S1hogBbVPO2U5QdfJMZBwFkU5dxbAazlrKgAbfFIVL5XohqoNk+4FiQFOTQRtnyS
gNPE56ZOsdfqC2gvgV1/uZcm6T4RJrEzVkZpn4834iZqB7r0LqYC/g4cUrBBA8o3
91lbtt/zAh6Y0K/gnzD0bLZJZnjV6E99dGSyDf/j2GVg1eYKZ/nZhMZvfZUQftVc
DjnEO27yqdz+DQeG2yanPMWvy51SbxhqwMxuJ+EfnOle3HXcNwXiyACLEhVyLK2y
b7W45JyCQZw/Gcd1DCrf4nqec89N1oOynkTV0+n+wK5WjakghpIYfjdQzdPR4V08
SUulJEr3HlnxHQ23OjZXNtgSZUW2jmb5xJXGaPq1sjEdOrvpmkYyBXWC91/fAK74
E52I7MW98uT4gnVm+gHOLCBTWesT9+bEU7Ivzzn/ORqDKCQKdDGhYi9HWEZY339Z
p7m9QKG6MfhFxFUiNsXw3PACelzM5yaaaUNoKlTi+SNsFXlC+oDXMJOpbQlURQny
zyu9BXRwNPjPh6HmFXS4KWPLpQX3Qjr5tFFanUlbb/1W/Q8xV3jdWhqrDC2BuKjz
mQ7z5QpiOPBv6bRGia5p+iqZEmJmk5bZ5EJb5gsM7+ZLcK3K8W7LwGedCZBU27o4
V3BGlp0xzgo7TB3pzdAV6WFHYqeeBiy3forq5UPorIu0gn30GWKKwU3e/xhxuHb0
dP1Wn1mQ/Mz3//5Jm1tVeuy29uvAE0DiT112R9DlJ2QvGNGup/QmC3UmPqyKXLyJ
vm+CX8wt1MlLrtOWDPUerSAJP006Pmx/V1BmiMYBzTAKtr7/yKni9t7Adh0tgiU3
Rvr2vTgG3ae1ftYXF7pwZbIPE1EGiQZbHwIjS+YGVN892fpTE2K2ryld9iFaj4d7
6L8wN8m4d3SmwQTC1JIpsfamH6uBQVoddC8dQLaAHWEpkbFKL0B6q6UUIpyLfVl0
NyNTdaJbjHm11N7p3Iu1SgYhbVoYP6ZcQrglaCaXbBAPGQ6GSU6m3xToNZR0GQ5U
Cw6bXHeqwJA0L2ND7z0dAjFmFuHEzPYzfgEfNCvHe6MQ7ZmTVSkFZPrqiKYhU7Vn
WoXYt/mkkqStF3kxZ4GF5QFLe6IVg1OatjuYmTItNerDSk8flBXBf+ma/ZhM/eQK
XTbNQDRKdMcLnhSTSl61vvN9tFcwl7Q0sfVkrY08LCRsr79fl03PzrePUeSQugES
DE0WxbUdJlKXjkqGLt5sGdOGeVkqWZwGcQsyEI3RqQO/bmGYuKbQKG9r4/Afh+hK
StasTLu+HSEInN+iNPMbjW83EZApQBoaxGNf2fnGWLhAMporS2J4V2F7YkQm80uI
r0vM+DYKNEathVAcdSvEoWdmBoJKQf+rqFVSlDFZVMQ+cBD7C0UjT2OCjfTLB0Ra
fdR2x2N+CqPzSeT4KSFq31ElTL7LgHHjd3MO36CLmpsDcEwIPkI/6sLJj83OsEgS
/OikIGMK/qhCDqSQDBLUyQaH/wbohJ7bjpGrf7uNi7hGpsyy9vm0rj81eI4D5ZRz
l47mt1KJ05AJKvJREXKn2GWXsGBnFtuurvUEjeE+dqW4GsKO2K6Rs2NuPyhfblya
5Jaw+RpwG/E+uLqjJc3s8hrMwsgB61w1fbfYT+rjf6YFwkuTQLZ9f4i2ypOPxgf7
Q7RAMHxlm3uA8DIZAKHwW1bh90kg1um1iWVQtqGoqPgLU5uRqVY8Kt9riQeZki9a
vhyAdZgz8o/DXdx0OOyjSzscfh9wtFcOKQM655/yCj8zVlgosQOOTJlIklAtn55X
5Vl+tcqf/iB2rTpo8Yb3Tzi3sR0xF+jZv5ej7n9hZxF65Ouh5yySCXlvLsA4HDgb
ZYqdbByPkfVuRL21LLL+P7eDNvrRgHcCJjqpFE0bYIVurdFecZufVHHMlWvShLz8
1mFrbC/C8ejQDFezqdS+FF1+1gFtG3+ZZ+Nozd+sMCkNxzXoOcpcw+gKq8wII8PR
NWGKWFsOlovikEZZUofzgKyhIEScGyXgr/sMdGK+qOdFyJza24gkCRh8To7EYXp/
WZSAaNZeBvELxCFr6bvMRN2naNXDS/14N454JiQFKt3J/yXxIORX9qMRHE8KEne2
yARnlYlSC+uD6mGrhEq+5F1ZQmcZpCBbbyX4vS2kq6JuR+JYsR9mGzflp5WPclrr
RY15rOcYYk82W7DTDuC2b51i0qEE0u3Jd8FNK6yoo1dwWQXmWl94uGYbzS3j3GtD
QX3fPqsS4Dm3NlRb728HsS1rfUrsu04+1RRk3zDHyL/I4ROaWVFZFak5/TDfeD1e
y/e9ix/h1IoFuhZGsPw7n3ysCULNcPf7NTypvp3QQt6+M/0nfQ6VLDD9LOoxczfE
SchitFAlqIubZYl0vTRdwC2rPwbipRFNUWiyZvg7jcXrrmwUvMgnrsrqosd6Hv9V
x/MaOA+jUMQurxf37M45DxEPVhZG/U+4hinKMBd4Pw3ixYuZQ1FjY/M3KJXZqibn
bXKTWUJIgzlNNgfs9CyXoBVVzO1BIc+YlnGR40gLflzV1c6ipaimlF9lTfaO2sWl
5OCN/uihkL+64xC0pLCWOP56QRajVTbNo+ji/dtvN4egcF4sfeiI5XVPZCcaYAwm
E2FYq9A4jet61ZkqzYuFIci5/iDoOLWFVydoHb1xmp6i25iK/crMa+hhZIirL5+o
Yc9fw4ERvDVEvTa+T8kztAJDtRS1e68pj68cA3Gc8x4ZPyaei/hTw/13r8w4tQDG
yYun6FOW5orPgIrNfDuzsouR/eNxg0MOiiC4adA16r6Lgs4yO2qnTuSlrpbc5zCl
GW3NbKEWlEK30Uv/fooK9IXDSs6Zq1xfok2hP5ogQ79mreBSv7UklUEYcz96fFdV
QZlWRmNzDb8ypLQyolNkhijEeqq/w1cjLZHHoxZV5/q/AccqRgm29EanUCgcovge
aRYg1nWt1FsM9UbWsCV9FT69Tt/y86jSJ7JoMBvoFS5RqtXTxAbSa4aSRSMsEIyD
MuQCE8JonL4Kq64tJAZJS3JmWvFn7ThDRFB9C9EfGPVZ27tqCS13FpaNR4KtwE6L
oNWkNP0jsi+BudCeug3zthNE7lj6PljIFHs8xiV1HVa4WTS1t/YkwVLex0ztZrB6
3SHMI3oxyseYGQm4fthGWi3v5IxgMFS3fvb9PQaLC8LdD5k+/XymA3FkSrFw6kE/
nNefg70knKoW5oBIG1uZR7f7w8C0vB/cmOWq3xEIHeqVeVWhVXf2QRGL5ZUjvBTb
6YsTeCiRxGW6SL7wIFQNmlIxkhZhQH3fVjEyYmy4HVPL3oXta5eQm/IeolbH1SWC
38X/SBTH/RBLkY0kVOOstNwKm7emZLCm2UBxJ7NNpx7GYndynsUyg/9OSE5O+U7J
a9EOUHzZeZOa3bsCB19Kpz8vTJserY8NOIBZw2FR8Ti9ChIIhRqYYSLO7XrtUoLA
TlN94Jo0L7BlcuTELCr0ibHR18Q5BLWG/h+jvN99AMD9TWRj72xGz/F+uizLDg3K
OapkswmXqku+22MW/yYdL7Cd43FzyenaJMshi+pTMWGaL8ugNbMSzj3ztGRgXwkm
/QYQ0Hw+ek9qysRHwR6F9+PZj2qV0bhmQHfbcM8g3IcaPSwoHff8xdxoKE2KqVuz
wSbXtPtaQzZzHsuQty5IVKft68pTsXbddlnIPfCSJgcR1gTEdB2OrEgT5b27fP0m
YOiuc5gSX7apDawljJF+UO4Zyzs3QBdREH15tGt/w2SN4qONoGrk/rRM4rSbH9Vz
KU8ZE7xMtaMtgmhWJiLlS3wokgeKQROq9xaCoaHgNlOS/ysuzQxv5N9lApoqXiNq
Cw95xmapAs7TKVOuZ9kitukdO1t7a6LAiHw7TZmrW9ZGiwjt43li+dUyB4XZ42Tz
IeZltvj+kt+p/ZDA0O0xX7KqG0311hYY9IpdCa74/hAWh+wRenSWoPo9W3bc9T3A
bef0e2QjfJE03C0f2X8ZGAc4yXmGvV1x/R2XWS75L0aCvBxGdYwazw+P5R9GSmwM
k0WNWMq5BvnYwaTKcEx8UhiTWaI7vITtDZ5J1MkBSyTFliIUHSMq3IVBMb+ruK6H
pBCEyVP74jz10tWUPoyRvS52DVgEvVq7rL4PpwDverdhYshzGpyoRQtu06njgqqp
SCfu8vH+qYMkbncnyUWt3h9w9CjD45KFkJ2a3zyQUJJTFICcNlToiD1psFuKUhhs
vChZu6VmGZimSMkyqtnziAN1U3wzsDVLrHT+5kVtOFkm+awP89N8kd8iIDpagZt/
VuhbEyMn28zByWTUvB4IWecbsKDksfhHwc9/qA5vxkCnrELRuEtdfOc9VTCcPA+5
N+wRILBMwPVmBhWNh+GilhP1wSLs0VETutQjzyUWvo9R45khyeScAkvW7Cte7zSY
6l1Sa7oYPN6l9E20srd3wc8CJwPyLJXiqAdi5DOvITYuThKSnXCyqAiqP8Ny4y+5
lj8iSYgrc4+92/BF7Cp8n39Ds4/fp9lNuXhIQfo9r6X5Q44H8Ul/CueycYKkxOfD
0wMtsOHcCxIBnneDQftWtJ6t9G/HJ0ZdQzz3VqJ18+GIUza/kPFwCC6t0Ic4X7Ue
HiKJ6jZHf9rWFqsDFNgHkNOfJPQovik67VTZ/OAAnZG15b/0wdWp0FhsdUnDcDNc
kFyaB3N4xK5R/cfOtrAQzpbKTiKL2kWm8SxiODZYpgJy5/t0ElhGlUdSNji63Y0H
MfXVV0oW34W+pQUjp1yo26JEJZzUfAOPh9X1mI+/0Ight62mA9gPMrhxcqZ19Z3I
H1Bip7I58jIem53CtqfxoIY3Uv3ICy2p1E7FAP/gmiH9kXK5kM77SetW6+t4bvyT
2+VbI8K+XS155Qa3L2jK5GfP153uJCdgXAYMpqL3W9ADMd4HtefC0kKc2GHbR2YP
DunY7cXwv6rS18gCsDj1cKB95/DPc4mygFWNr6ai/BqVq37QqmRO8Vl00lOxdiSB
qRquA8llBLlc5MHaUuJtHd4HYCnlK4qDzw/YFcp1L4AAJRJe2xzNaR2y7WCZWu6I
FXZXigJWwJUBdoz/obxH//kBrfaK0CIMtdJiCAVRGTNoA83JzseTYknZ9SX2Uei5
T7SdxEBG49aKbpH86mCiz0dF+TzxMy2tjfpm2sm9S4tu8nLfFTjKyF9/Up/KuW8P
NBEYJJV+77//xVbh9DttwAPTg1Lh9R6JuQ8qxcfIwmkUKzWOTkhWiPveePn8YY9g
BBycIyow1GB8esPtRAYUF3lPZ2+Dqv90xO7pdq4Y416UI69zKofEv99Crp0XrlID
tEMbnkVbs/+m2mP2zDwwKqLMDoO7SKgG8T5EuALjyXLA+7U+YsxfrAxLVWUrYI5C
9z0RjZeKH7iqWkIcikOp3Mq6e2Dd//QrngEkDmAEBDFFjpmd8PBDWH/bQBQhHwev
rPLiSDLAECW/yAbPct4AMivTTT4tnx6z2VM9u3HeryOgUypptZVtg4kj812EED4r
9K06DogtgWBrQ2AO4hqsQ0sjYff+XZ4Jj7x6Ks0M7lvPrSCAUYAVjlH+8jrhmRnx
Ompq/4wgKXz2PL8NT2El4+iFq6B2wpR6D3OR7wEfx4FKXx7c4zA5gzijTI49ZV0W
l0xRr96LpYKIsQ3rvX8L62o+/thAh3NWt8lHg4UIRU3bV/dffF1jh6iKTlneg1TA
JnNk+xSfp8re7P+3T64ImXUV39hllyJpxC7xphTxMGiUZ9tXqwf0YlEy76L7Aara
lfkX5fMAOOFawDsnpbEsqv5WoAv6kRcphGeFNERKAh/ByrkudythFec9T2WO8U+R
KUjrxbNYQXRwP4yJVA2++5MCay/nkUlrQjMcU/JaJzQ3yQAJZWlwFcNytMk8eyVD
Uqfu8qrpDWYpw2/y2eO3Bzm5MDXeq2dmsFqqS3CYDCQzxULLAahVgx8NaoRymUlu
xw2CqLytgesxCBUBB+CIywFDA0Z1RYwXVkyvFSBS+5yZ4jukyXJJUU1suhTJqZff
PrYtjCSiy1z9M9PBbtaVOCADGO4UeMCNyWdF2kcAafyae7+rclW42hMOTRFQSjkS
36uph+si+DtI8WrtsgUNciJfnlCGfTldINY6LhYPMNuFh+VOlMId4zbTGZU2op6o
X0YaLeK0xOonkSKRFlm4lsO1JBTlLisu0/FNBnMF9Z9ZXiG2bByMCNS8y4e5Y3N6
spvhVnCuJ0kc0CpNHkntPtK3Nb12kfMIWim5+ATsTgRhcR+vauBgvchhT55tGIO5
kAIrpA2DUqeQ006y/lqG7llhoy6kYM5bMg8YcUqVVdAuFSejipqng5ZiBUN9Pltv
DmZAbyuJRtLqeUBFoTnEPTHd1zYPHht26s/qgdYF+JhD8jCCx8UTKCUrixjQJBWh
dLpEw0ax39WYm5SeZvNPK+sWN3UqQWjTTsKIVAw0hc8alwS4qHBus2CboITHmK/k
PvrihQIzv+WvmnnZsntnFKuQAcO/qhh1Shzq00NfAwoaquOgve3B9lNLwWQwXORo
dY+kbkWsQAOzZ/AFrM8L8QKNYVk+q+6AIUB4BvOOm/iBR6WA58wfEMWGt/rq1xNo
F7cdEmlXDdEAXiTsh3/uftDCfIBlxD0ak129JE6BwNagjjfewC/oW8gQdFx4nGDZ
+lvRkDSugQCK4oQbNAs9N90qxqMgi/Cahn9D09I7JSmNTPO9vbjfQF60m09MuqJK
JZGH2GZnI0c4niOdHWUu3dq3yksKMLsRpaypRmHzWGbl7ZCkBgrz/C3a6tC77Gqk
vq62XPvhA9u2ZeSkXJwPmSCEJaldQ/BKTk7bDyH95LFz8FkLcMRpP4WFCGecOIyb
vne7rHQTPZOVg6ohOlAKsQv9+0ayfarbrT8LbRhSt1GWnY0cOTeWIwndNjY241r0
sthrfQbx0xAuIyrLx3CZFKp4R5Atvw66DwqTtgh5VfzQWcD+G8DSSsuaA6Sqex09
GGgaKL4xCcsPB6gA1kERuJlsDrMDaa/IpU9D7svD5whV1K/p8ozZzOJwaTUasSvW
fp9ito/yt4pzGyPtyt+gT1H/5DFdbm+smq/76twAVCV7sxI/FpKICp7ReI4pvXdM
Aj+HrSu1OsgnC6+ZhdqCNoTS3qJe2aiXTH3BkG0S1/1fwGuRilstb5zM6Sg7DdQn
hErBudh6VcDLXYm6MlRKoCsL/Vurl5lQI7/cVoCCweb3Q6BWsjeiwGv3m0NnJjNz
dDG+OSirSzoD48mqSXuXSbd4ZTCzVIsAbk+45vVj6znfLJERviKjnbTEXXDxAQjJ
uWzogtKudvmmAWzbP+TA2r9fBQCsXqbscGR/PDFpE/jBhv5TJ1bJb9c52uYErpgG
E3UPPS6hbMKwQO9huE75lyE8xiebrzgzj69Vzl0QrtRkCyHXNQZ/YDDhqIFnsItt
fMVPd6yNoQBCvVKIeY3RFFiY/PE3DS3xPc2AbW52XNK0esi1omP6okZGK3lm5y6a
50NVy3vDVCkJXZTKGk8NlGen7CAJVLETcHw+xy4gMWORCAyyCSZl+qGYlL9iWfPX
bn9HpqpzkKOy9x1u0dC7XNtvBnFK4FXsWIu55pcqaK9yxD4jfIl9SJfzgpWO1jbb
Fm4dz/4Fvhb7v1re74EB3oEPTIitvHnuuztE6OHJASNvbc/IeoWv+ILXlHr3AzjE
rqqePgfwC95Fw9SnmJeE0xk83WISsU5PNx6Wu2UlMecB6N7m0CqRlSrtYwMtZDVW
gPYq1ukWCrLOCzmzO6yGfZU0l3qbOZPZRNVJn+no9tKyjx4UUiAwsRmBT0v2q7NY
S/boSJjKoDwjWeQllgClLIJHqHNZshi4hpWgOqAvuaq8VZ2FJeL8v3DVQumJrdH2
f7Y5vefanAyLy5iG1XYnhKMR9OfDPHPRhcFSFMymE4s3KeS5kB1nhOKou8c0/vFv
TrfEF49TQItxBKk0xRhH3OsRyJBzun9OgNXduEOYG1xgceQHCRySmkcMXlr72FkI
D4+rzztlgr59bDWuzDi/ybmsL4Y6+MJTc0K22W8gqFiLfMEJXG+JaPJQSanqz8mr
NoNaI4RvEBZL0ZOy9UkjakJdGsklaIhD9dm/1WmzrKGtpBdBPMN4j3tZBulfIgUo
dhChBEgpLjjvYVm7W2WtBOiXr3uf8DKrjpwLka8wFFwRiqMHxFXpjKzPUhjqiM8k
GHB/71acdPaX5GDcYCaz50tPkLMYnZ6aNqD0U3shHpOimiHtpfZcFpBU+c6RWd2m
YHcTjju5n3irZ0Q2Efi+xym/S6pxqGag75gthIs71fRm7OZ6KOwItsEbU5JGWbpM
5i3hA2bvOQokbJgAzxzQ8RqjRJ4m27/ApF6t9zc1V8UfM5tBIAfhKua5fxFuQEYf
VgsgbOOU1XH0ymnUn45R2E6IPb42GYJ0xhEjhKrVHnSqXzjSvEzg1S9fR/d2QXNW
mph+2JIXWUORmD2oMlIBD+/Gxh0lxS8nGj5gk42L77+qBgAN90lfThjmbg8dLOxw
x3Xti/wV+c1KetVWW6dK6jCeF8FWsI1fj/Bd618+VR5YcUUvo5y/hc7iL9QEUbat
PJ/byOU8pYdwV8W7exeL5nJgNiXs6/ytZDDgB9f5fgQXb8zP3JnvjL4sATQ5LW4q
YRhhiJ7K0nmIiy+dzeQVU5x8axzY3zVNq0kr/nhzFn7ospxM91WJlWJqZnHazULl
9B6GJ1gawIwP3WKwtCwtObJZVGp7UmgobcAmLwALqxKVqlmDhNWU583D0J80H+27
bK+gXYC2pIk/cpKJJ1/Xi7XpBmvkY2g7s/Q7zqGipUtab3RMs4EsAVtzxT125dVh
cX9XKLrAYxjGJrDgyl6RkW9J63XK9X8B1bFo7YmPe3/oyRzaxkN3MVSiLVFrFFJJ
rs8dcEj5OyNNCXVKxMpS2+r1WF7JBdoiXPv+g++U2mbr7N0EwF9rAt4Dlyj3QZXc
ejILpuxFoY09q4gTwhzsJOIzcOrYU5mldkP9owAE8Q+p/fMTCifO6qaGpxyeFeAR
4OmOrm5pTuK0MM28nxXIDdhuZ/MmCfglzNBpC8JBp0HfB7f3Sy/iHqpBuA3Wm523
SrN2kWhye2VcmyXfvWE0ZZLemI1MRl4GnOGpL9YXP24Gr7vpi5x/uJPxFDXGHC0C
1XnABo5V21kZYRR+CGnrMY18mpfGhixIDLW7NZHziacj5wY6JhV5dv4kpjjX6Maw
vcqaK35t/M6Wam6MH6svHUpArmMx0OPZTRbAXWS4Y+GD572bT2J9ddx+SVmr++6Z
Fq3skA53JApwd/UPRGWYAOtaiDeMnLAZEbDGtwzIZXmq+cxk7BwqVdb79PUgJmx5
AKIGphVmUENU3gmgJlOWiRH0OMPLFbc24D1eHsZC+arcq9pf6CJUhB0fQxKT7FrO
BENHNeK2x4odjXyzi6XzU/TAfouHRxmU4vmCu5lUZnUbZZwFm2QGjPlifWA7KCKf
XhLF3wz3lj3ll9rYZw9W/pplVa/L8Vw34dGIlkzY9+3Vpikzsc3pISMY7vawieHF
VqPrBS25+3mChUGP/iMn01wCBRtvdNDgSIdApkavF+sqU0XAWUbHqbDrRE2krWO7
QPw2GgaTsgtpa7q055zSOGyl7fk/OPUiV/Vr7WuFt3Us8CCji1JqwJg1TT01mmyv
kdWNx0bZssXvSl/2q7bxt5z092ZT26wQYcgfWKrrPlc8anvy6Lq30WZK7JIavXKg
3+u4r5G4xA8RLLHtbdZqEaI+wvfEyhu1583lGzge28B7lWbxh83gMxCkgQ121YSR
6uPqZfF1q5NPHBuZlEs3G+9aVeFAfr5P4fNVE4tJ1U28VI2OBNon20r6fYIouhM6
YpfOlD9aFL6ZWpwxGLOMheWLObI1ylmdKk3kkw5Xz1eiIR5YAQYj7yxlGCLHBRX0
3vANYBPNfoqQGnF4/f5UTlhOQK6cgTeBEteSij8+/pTg2iJBQ6DYTp+vVY7tykKq
bnTit23YenWSKpjdnVdT2wUMG2yVrH2BYhMzj6GEO8wAX4NKGeDnbkGDqUQJJAoy
n4iO40imuFHPlqeSHAFVeH8VBH+ZC64CtIXcY3H1i6zbLHjl7JYPjLqvTNw7mWlM
K1WTXzqhVt+n78H+VMgfaTVc9bshaBmQE2VAToDT21Q1fV9WvW+VcNjS4MXuHb6a
u60YM8zJ5rxOFd39aYaC4RG7OlRSzIxdSnNtvtvN1NNl0q3nb8K34SwCVORI/k2T
I+Ukn3IZ2S3gz9ySBVBXvGJi2ctLQh6MClXqlhDhG9AF7+mFiyULS9B/ZT9jRsdG
Vswz6EBWYYB9EChIPfFFf6x5MCIR3UfafDjSBZXXi9ty3KtHHDC0OuuFW+3lXamH
14z+uabBzjbgNt7tW/ly5bM4Z/uNTAXkJkMfmP35ULsuHxYAqxlp/GBhSN7rWnPQ
w/Xr5Am1FWVyKnS+eAi70uPyp9iSmZBEdkcMAiw+6zh4d051Ax0dOlmpaG29qGGs
eNMhIitnXF32BY/Dzh4SfCvY1IEJZSreRKIZl/n7gZQCaCSnuIGaKbFh0rT+GC3e
PQPuo3FkXbmvez4QrEAgB3ygzg59ir0zDtLDvsIC63ajMWo0k8UnwB18aUoIZou9
SXw/DSy+DmxMeZp8MjzTeF+m770t3tyyTFi5W8zUQyr55P/OrgIQ7T+gRCqjUNJ0
d6CTNFZylZ+FKMpvmE6Fld5GjoTy/5xQaYq9V7x1rccBSS4J7e87IkrbHF8N3V8/
Jg3G8GYcHceWznJX1fz84aRAqHQDu6Tm/uc1v2odZVjHAKBfQkCKnlkLsA/nCGo6
yFyp5fUHmC7wg7VVgENk8uT8At7ARnY98e14x5oOXoug5kUNvfs1i5Dt5mUfPDBg
6LWEJ4y9pZX0qguDYEwMdVTGRBDa/5+avJT/w+Waz1VVsyqmxZGykL7Ieq8a41vu
pcMW9ImQLezymEe9tNMQeNhkaWPXO4nNDDMSDsR7kTw/QjXCD+tQWcq7sYcky4NK
J++NniwbyR54r7ttrKst61eKgIv+J5YSd4I2vf5fvuAVb3FWQ0+njEaaJ1SuPbev
mYVYLBDxqQwE5Z4DjKXTaCz7rERRjH/MpvpjSvUOTCE0gFVwwH3mJ5bxvpbflq2X
lg0jJMeN3V1JPKbrvmRAPoOYZeKcss7nKY9m2jOFo+FoWuGUGoV+x7UhbrzP7bF/
X2hUWVXPolgwtbu8bnE8ZK6b2SFGoKwHXNpfXYqLaMZZ5zFHp08lp0qvubARVdml
8TgqSU2s+fYwG8iW6TygC93IO3Ef1l5lyBlY9TCeVGmp7RjfGvyI7k33uFWq3QpR
mAIQwu3eXG6HU7COGQbfT2hQ9pP3VHv3LwwtSO4q+bIP3ZlSdPzltzZ8oXfXu83H
3SW/P+ul+TiiWrvZ+bHjMaaR96rOutd4Ft1MKvmxPXCn6O2jlt7bkTJid7tVgyL9
iSc3Z8uBiu8ZWt0lCwXauVZkiNTUz5bKgwPN+YF9EU+NDkHAkIDiYNKIlc/VCmey
`pragma protect end_protected
