// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pE+uHVJ6GyBm8BGUjLHArkt0z9t1XXrRZF8Cgq7AS3p6XoQvcwtf4y9m029pG7Rq
XUVkiPUx0d6XZSthdBqs7O7wkfVhUoh+wkliFWRFXl+6pxkOkOU5DLVgKO2E1mTH
Wkk6qVa4dyWeyGWDxmi1RK5/SYH2B+ELtF5qPz1G4q8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7808)
dvIBYFPI7SR6/yQXdcnl10NlEss9PlZCJsK05vr/wrpySmn4pSGNtV06l7J/C2yx
J2l5qz5ses2pVbl/0ugBaMRpInW2vmK9H+ALxekEVmgagJMKxbUTj8BTfdoC/cwX
nxhY+7Sjr5lMmXDfuMUypXr8bCPWPwbmo0c56kwbd2Vnh2sFJnpXp1Pq6gsbFwe0
r1UWgnfJvf6127a4pPwAnlx/H8gSU6QqUVTamXw1utpzwuMdfjrnlUt397dT9kgf
Rw07W2GqEzIArZB70teURaWMUaZ2Aqr/6UUF8c+jxUOKHQsBzMiTmswbnf15M1/C
8NCv4I/bsodjWc2bMI/oM87N8Mj2YOkvsyfJCYUXr9mEtnl82B0l6vqAQU31x/S3
zTQW9e4vaVOFxv7V68xyJ9//yB0ImBB6pVs5+hRF4j9rKwKUg/x2tk4FhCcpuwI9
a9A++nDK0s6K6/t9AehBcYJh3EVUv4yRrogoxp+ncSUf1F3cn2G7ca9k7FdGeEX3
GgoOQDN7rplGGSg3BlS669sBCN6bDsZk49cNQmFO03G8F8s84biA8TLINes99i3l
TTfcpJSMzGjCW+RZy5qFJYtg7FTGERJP9Mug8B562vxle9g1QPSN6zdEoeV27Ljs
HDi2L0JDk7xzgtUYt9HscjHneBIQHMY1LexKCoVJ1RK4lTieWtiz1sJK4pqlc03A
yptus334GI7gkscw0/X2nWHy3Mkjprd0BX/+7nqnnvGgHE6e+nHafPDGGBrq21tD
oGLRh9cg8hyFw4onAEj3jLqBCw91SkJdzQsxNnxlbDh52vZE7KXQ7IAO5HLdNF/h
8BoRCocGsyR2o/1PFy9J+PJMLTqDVuEbv2IUsNgKuV5WFDgVpva3LfSueuKIe0zz
BYZsxcyTfX0frkmkuaz+9+Wt2RaPrcWbL0xRcq5uyLTwAWT9g25FtZwbsY0X+IU7
BKW+u+BZS6SluhZ986v/J4UhoGlrSE0B61+KqKir6XMF2dDPAEObqWXVnsg7wMPw
D2jCqvd2vnWn8n3jgT2I7kD55e2k+Ov7cWhQJoZmxtIxsk079mKqKLg0jS40E1Gh
uASUgyW8lZ0dkmFmTqXu8utd1msoZchRD9VhmDEQjOG1RZNz2km+JxvLnRy/ytIL
ShInaM8EtqHIjhY/RKGHaZPtDQU0PF1A++fA1lx1b3JYF4fdWJIxhHxW51fsnsQO
wtvgbkO30D8/RkRvaWA9HxVlmLChbqteTHtq6V5wEzxGKHOrMmSmbDkxz5Gjaa9y
RsiOcWEQBdsMlgo79CccMnupENB0lI8UR6Cg+/uKZjHHKqifX4JGDCVrEjlUStBT
hhPKL0YNn4lET7FkEm9fqz0Ibpho47Qxo5Eua6aLV6SECmy30Qz+IvPhKhfMmJLu
bLfso1C0QAI6jBw7We13IEcAkvK/9XKUyX/a+6KJo6D5yesXwDcNABCwTEuUsRnO
3XRWUvgadc89aCgRHlUuR/itmQIiFi9y6aZa41EoPwi5m968j25PL4bImygPV/iN
Bf9AlZfmX55Y/XFNdxmn656FZ8zsQFpIGnHykukL2ncUl0hf9FDnvIzbx/S+zTg8
OCP3S6+HTAvb0HJdADmf768xG5e0cCl7KdfriQyfKPmNYqRFfCIbKWFdWdezFJny
g48ULyoL/u42Up+O8jNrOG8oqWyC9kikCI+73iGrA6Sa6A3EUbPpddaRH2wvxk51
SjR+h4H0EJle8cfvc8AIGyPRY8jzlwvoKQWTbRGrhf9PJXOn30hIc4goZRJRSaWJ
BkrXjniOI89s57KxMYxO0lSX1fW/qYlLCMtdqcu/dq1NNX0wupm2plCMidUXq4Qm
F08wkYBeQtOrX6L0B8mzHXs/wHc7nKnXr310o6ZxDU0zLcdOXrG+wBE6y9C8GCj1
x6/le2F0CEj4MvrPH2j4SGRMicpgtS9DOmstpn6+IYhsyvimUEmNawNmnsCrl5Sb
aYnEE/1LDFklx12Ck8Us8yZH6x7zvK8AVFXlZM9MKp74U0EBQOPYTNuvU4LkT6DG
fuGoo2k/ULdjiDQgej8Ds4ZKrKMVLmEiIlrznQN5jjuQLHv8T1FN1AdPuoxfEkPa
s75w3UOOCbX3Lb8RoZ7hRe06LM/4GHVmJahRv3bee4vrkByhxzmHnyFFa31f45Oh
ULGsLmxd7k2HPmiK1YfzUXsO8W/mBdapDrDoH/JJNOO4J2+vWYakX+2Au2ACQ6qd
QW0hgkT58TmtrUv1Bg3cwfxW6DokSC1Cq7LU66UYBJqWhVAnVAOZdBx87EB66BS5
S3mQ+vgnlmjN3T1p72KfYZWRUpktyrYIFqOP/e+w7GDrXwfP8L0WyTYy4Rrr26yO
gXWYgszRUkEwzZJ2/i3eksXtp0dFJQEgxH/cV1asiT69WAgRFncnx6pax2ZBCvT5
64khvIZVFODnahNFhjmjGqjfKa+Vgu7PCMMzdsFQd6Kxhbmapt3pYxhcL4Sf/QFV
+6aLE6hQGZFXaTgN9uvKobTdsJ3FesOsWFw1vVs3m0nsFaXB9PQ3O5WfDeHwmgxP
R4N01m4cJr8cer1knGCIn6qZb/sbzv394CiubDaKINXGKq8QfGu6o+ILrVAFr6A0
KOmx4fWxeQ0uECSc357RhjX/IPP8TYPQcabbi1y93efT4xEuk1R46P+nqZbjS6AU
aCqPxHqKjQzkzZY66tiaXvSH9DAFewffcrqcvS3sH2ekeGqyZVgRvy/8BzfDyhbj
oH24Xj4MCL1coneKLuz4JKa8eG4tCqd+DVHhh7JqyYVN2CM1XcNJQVWD6fIC5LXm
AuFXuXDluRuEBP6bLqGKMpEBnLr792nk/fg2Br5Ojw2uwBKRTVJChhGrhT0LfjaX
iJiHgSXdptr5cZ6lzQe8hPhPqaiJAybGzbjDLtLGQEIbz4w1WiJke9JQ1Ky1Lpox
Fgi38J1WfL1KTAI6y6eg0XFNXQp+gBI8WFgGS3tiH/f8hemlN7fz59glNGWAEnB+
0T8SI0C+XUDDaVQ+8Wcp/DJVTx23SiE4Up4EvY/Su0QHT0EFUGxk+SMH5ge/qgE6
3tmoGuSKRY5Ajo0KfvW3R4hVUrcNmlvM8+j+0t4vzce/eHgf4MI8YD20TC8CitWU
Je05/zmCFyT18V7cAIF3KDcudIEXDQ7oNEnUYSsDXhMnmtisTKlU5NkWvD2W/qgZ
ygjrM2V+Dv+H7e4e1Oa0QhIW7Dw0UKmk5hJcl8ALht3jvzAiXTW01CnPZ/opzsxK
NHof/PuqUR7vEkiXGTIsIiJjztdmtjNuG7e59+Y8DeJu7btlcWbH+xGc2gt+pdMc
ilADbBYAwTLIKx6nW9YNegBAfHVP/H+zSFNkO7zr2qz69h1P22o01HHw2uUmvsU2
uZlrtiv1X5sEa/vzNZb9qOmcQ6uqoanxx473qowvMIlWaCGURARYd4XlDxc/BWTP
+N1yBNufBMximWafuVCw1jyPlrUh0L6Gsv+I+tsOwR1GR9PGIwfVCx1AxV7YOEAZ
3D90043NV9vj58Hvv/CZ1f9+K7HuN2LyAVF4OFOZSjkCaO7gcB17ORHyE8ady6bU
lEG7Hdc1IBBtg0D5EyCI/HJxuvFlFFy7zhqEYCN5qKAvzqpv/Cry/69M712GZ228
OFTBsepWssEmz3v19Y090czxqutdn+Cpsfq06AAJAPF6fTHwMIIHxcOO3OeCE6hv
6vK905HMR78E1wS/X4bW6QVwoPPW8QO4uxATixpJ19SZSf/t1wL284dogmPknKTd
1lUyauSF3duEpxQfmSxHsW7U0evQDVuiA3kBEq6oSFMk1sjAFTO+6RHgsrBSHukY
APun/dNRYvzLScaggLQQ5/KxTwpbWahxkieWjy/0JkNFpViKLOO2j9Bu/Clv0bcX
ROLW1+XBkjAQURenLDXFBsh1eeHmWpM1P/MkIUJ4Ar8NDYTvczJgBIQuZvtI55FJ
oB7dQzBfh68dmEWVhP4N+eH/nkU6xS8+jXpy5azK0VrHltkTjEfgTiWiBc28fT1f
107mBkMe3cW6zEMtimfBVQ1Pp6aEjhwPrVUPDdJyP3e64Hzucuxa6t4LrbQPHHCr
qzd49SVaKpOGkqXiu8EIefy7csl5Z+8nt4y05jqjenRIuvJT9YmuKuy66r7diI6M
kubaG6Q4e56ZF85RxsbYFy2erTgRP/x9r/ubnahYNCn7dL8Tz9W6h4fzprO4nc1u
PbhCMX4rvGpTk0/+g75PqX/WQFW4dVuUxh3H4RAzgsXeSH51YvB9Q32xRbL3xSd4
UrJjuGyI7KZQZ8YEoPYbXVLIG3PhAbktN5qfDju2LKHS+/vEV79h722CTevzpkoc
FSAgfvt1Z8Io6lLfVkt+tS/1k7QStxr+SoGEn4EdGBsG5ArwQAnR2AleJAKzBpsP
ptemfiQm8dArukeEF/q/ppedcjG+82RjWqR26FF5lxJGcwcsTX3Xd1/0S2jFWIff
TxOE94VUmsptkRUx+avg4ThheKyfDBeDmEUDLK3wxabKgPnyMfPFo0/5gZcbrwd8
uWiVOMQ7VjjX8qSjnca8INV2cdemDbt65or05xl+lcDhnuRtsY1U4IL6T4kDy7d0
kFcL8TEVNm8OZd0RsOfNz0od7/20T9UHfnJBZMMHsoMErAbr1AaxgR0f18X1suTW
5FBNW4C3T8n7MUpmWaM2r2f6CtrH+vMkJ1P1WNCTskDskUz9Lqieh3qyACVfJZ6p
sUoy65ou9VAoYtUSLRp9l3Yw1V4Abu9RsiGbCh9qs6Yt0DBIsBaayru0CZfwAeXw
fIOiOel2Xf++P/s1uivrqjPKpaMkONxLx4qobSefcYBJpk85BCX++MgboJ94mhed
jWDmaMmrdCftx4ZmTQX9C3/vfy1vtUL4gTxqbZ1vUvPSwYMcSrXD8gP1adxzPOcV
euyFNcC0KLSRBxWzl9VDoPkj1PDhCQd13RtHAYxQRKdvkOnwKBJ0sB70bCMF4ZXP
fYZcER9znhLqZPpzLERFthSsP9QPQGFd9cZSwfgkt7zaSiZMhn9uy891lxaaLHnQ
+mpJfYp6WD2cKPDUSjJK2eou3ljnUmEPl24/I7/vxhAsirW3BI9+bsUd1LFyfR9r
Tkzmm8Ru4k9222FXZeg+IswmM5fvcwuL0suWxaIlaJbw6swt7YSCHHTq1BWPU6fa
YsmH4NIdzoZ0DuNS8w0cTZKQMHDFujb17iOPGtz7pF8tC4U7wGKkWaXoEdXW8cR+
uFAj8oo4Peedjb1kZtfYYgOXUg2EmXUIO3MpPoalgCtemI/zIHv2J2cVgm4cJVoU
ryRCqslHu4PfXMx2FZjL9IgBnPNs2xSIWGBckyXcaXzrQnKTq819wLMH6OBfUgtp
2Kf4MQAgoZZ7cJGjATQXheKV6uPYPqhp9B+lbE1UoH/VCNFefUmqUoYZt2IngDoD
oGRFXFKBijK4TnRJhYy/AoIV2LypIzEt/pCQAYswP6bELFZjZRYjMWTO4QvE9YVd
2XHasWivobZFT19Wnm5ucErjfVEBecEdFFWkFvEGALTXd51am/+deuq0CjeS/3Xu
s219obyEtWniR/0PUxBjc2xwB+WoDhOxu2pvQ+9Z54iG2/f21CVPXqFH+Va/u5yW
x40AqaGkUeE8aYdGXZwECe9KrTTLaz1eDSQxskg/GqM/uZdAb4kMvELkNecm+H+E
rqBXuD+z+LwP18/4FTlx9MQWtiyqoXOS7Tw4N4r2G4Ci8N2drZ0xJOlxJCPi5V7O
2en9BB/V7hoKDtj+bPhQDf6UtAOSp0oBYZP+YLurrJdDseUzM+23aXFr5WpxXPu0
GdNPeKbA84aWYsbItSRFAtDPGEaYrVMNrVDnGJC2xLCqz6OcSoGPYfe85oPShMqu
KsdDzCh2gy/+qOK6UEPNPIPb19ZJvuryoU5sgkpbTltEdiMfkItVxBQNsw8OumCP
CZvLErClKpv1r1JI9Fcjq4oadBPncV8EgetzYjYsEhS11sdK+mIYk2VZTBeVMA1b
1ZE+P2fmiS4zjqchhW7OOIS2gStI16IKIexM+BBoYj28mV8K9mIXehpdil0ue8uA
tVv8cZlep86dpp97uSzCh4JBQ+9uJZYWEF9thPWP06GdxjpcKWTToy1aW/3YweJ7
tGpRrB14rE+QR41mwuyI1Fsn3yvbK68+hKvkFVdsSxbW3WW4Ii1wTWJFQk43dfnE
T5kH7yD9/dME1L0AHRSes6EIKgjnDDzTETiDn/mdRovYdN+MjXUNcAabdhoptUs3
2ahEQZrhwOZK2fWqSf6Qd/SvvvRlzPRkqwEXcr+hXsWmnr0/5tXr9B1gFnFDB5Is
VI4BvTDEJhE1aUMPlUxplRLfJN5egCzbzDiXLshbv4eor3kIshb5CAu0KsklEmvT
crzNumZXxs8pDGiBkyhTALYmkJRvEc/goZxYOzA6FWi/XK/XZ2xVdF8LMNTyAXl7
kb0qIn9B3bnOcyhY/zbSKGbZ0n7J/Ly9+kJEUklpbZyNroXNgWbctXSXnouphP+j
JwIvV/vHCsgMVC1aAEcwarqHIj9cZwquO0MplB9DFYTxSz8iTRq+uW4VzzLF6cgU
uD3hMwPLnM0n5vY8LRwBe8Hn3XL1andXKyMLCvMCE5d5Cw+zb0rYoGjb5z7nGlGx
jbazJDBsFvkBHCwIgOyd2Z8yXnCB/agCCeZoC0Gq3KYH0QSvV56WNxG9K5wJMUob
OspJS21ltmJJEp2FygmQfj4yNtyz5vGUv99GapuaY/6iQrqgQw7atySTQM93eu31
u/OifQVwNSTCjZ27S1D3X+GuZlQuo/968DABdNVFOKRnhoIrMBP2zEyXQWKvfxrp
ghl4lQPRip1fzIRIcGoCnJ11+Pod1PdTo+J32Z25AwttHGmIkpMq/wLQWbkN5a+W
KPNWS2Y7oFe2TWgrBTJNvSgjQzUgWYRHpFtTd48V3gncmCybANsBO3dID7mtSWah
zC8PjrWTK0WHeLSqthD/Sjrwl+AmcwBP0rf8/d4x0SSN90nBi9HpqJfIdKKlHZYq
7mZzYpV5YnZltNufhw7Gee61wMHp6GIXoO7boMzVCkxYFbweO6gx+g+FqyPS6EtA
/ubzZmbW7P2PcYtGrRm/3JIip/Ece88DnUJqa0R0+9d9wK++FO7KjHCP9pVxNLPG
WtMQ3OSDYKTpn4p/r+xu7cLeaLIFhye1kwV8Di8+rqXZq0JgxXVw0+HqX5l+9Lic
x0zyh6rEwjZwiC1QgBRFQDic7YxGqFeMyUH7ywOLxeTphRepQLJvA7Zl5KTk5vXI
XafvCzH31Dl1U3DdOjNUI7L2gwhfUAAjhyFXdiLG5W/4Se61779yf4TY1ZtAAGcv
RhyjqNTnFh5DkNGGJdAZh2DCDJn0ukajB1HfQoszvHobTo8pnGGjgzzJcRXZp/5+
eLtoqXZnhhiLZ1eUp+D2EPSC2C5K5Noi/zWN/y0HHtCzmZbrTvXzbwnM8qwENHxc
q0KJJo7CCJzq52ZFAjJZYtc8g2SNwOG/k6WfpFpjdqh+3TnSyv5qahK6FVugGgRc
SU1m8xc62EjtNpZUk8glyWLr1WuZlODum0V7hJFnHGIWqD9KzgEO8LBPydmcswxt
OmSYVSTBRg2IcRkBptyZ4Kju+d0fbQESkAjVQRGHv5kTkSLJ0vkOyzleh/lCDKE6
6W6vMW/JCVRU9PS6/3g53ozcDXQrvYYzIyj9+dSYmT6k9OH7jINCWVsZF48cN+Zm
wwtztVkBUUYStloP5Y2GO2zqx3jE2e2abXjJq5NjZjtrsKLSuEjTWqHjF72BMX5F
9+6PezeZUdmZUS6WXdi4p4SoeMkoZqhhIzwl8LUCBEftDmmR4kDV9qEJ8tFyIO2e
SJQMstxKQ3GC16WtlsMXVrJTkeJLpNDikMJDMObKsTIlvW7hx1vlP3rCKpAgBJBy
IHntTF4athy6Hn41AYcTfaxAJvpZ3wDls1JK9Sr4BFAM1TRM1VLOvPSMFgXn68OS
Hdp+/Fcg+zawYFRBbkXWmDRFUBwrOSW21ZE3xKYMHzQ5ablMMI/62oUOFOTqkwhw
Ct4TSnwXWVD5LXGyeWPWUCWxehlgCLcykEBOG+v75sRihA/bEvIumQmDwOL/JKTm
cFwTDDTEtTsR/kn1hDWjxGXBneW4Y6TTgiRLO1CaT47Rz5LHguhi/v99gfGpJfhx
JSI9krDb1ZDjYyUkCMgkiQfyblkBCoUJDcBsGbQtNJkUZmTpS3l6IAejT8OcgNaQ
krPnJkQMHKNihLUMVM3dlyOQsPUj+m2zCCiiSHZBUc+rSVDmJsTsQ8iozJNxL4j4
5hwhwV4PKk93quAw3a4+GN671iCmAkLo2W8Ysig+OQMMdDsPp4hvVnS2pomIYpMY
2xezLDuBm3oD7+/VpuNJVQvoXy/dgjM2AKvfjWzlnZ2DqYVU0gpcI+V9vBQwMuaT
Mj/YGGkEmII3ZLASd5iVF1Xgwq5eAbzID5LAfhng95GfcjKZ/2UXVGZSrHciRdFa
6HZ3ExTddfdWy6lBL5x9XtzmGwfSx1MtzhXeuLbI88hXMPkov+WWkt8mbADqsaHJ
gowUelndnW8fOojpdaB3EcD0nIeg5pUoV3Ku2rJfTl7xv6UxOJEuBC+rUf4yCUk9
FikQ3vdr1bXRL60CXT6dcd1N/3fbB26UK58fSKZuaTaWq+pAO4d4GrBo+omsIMHG
+UaYco2sRx7nAIUxGpvtUWrgd0YR20IYNdVoU98ofq4pph4S+GYJ7WCdlGgvmxvN
gDiyT6WPMnMC9IkthTbbSNPjqzeJDGwXn7PgnR1jQ8nnJGxe/msbTOrZaMpMxdVM
CIYgGQc/qNYYtqmndq3kPW0ZGzFCw8Rphv8Y6HPfkakJtBPa6HfrrZNzGUU/8suX
dztaXZf+7tnuQBVHrY/RKL0gc7zSVmjTb4H6xRdE3ndfLCAGS9FJGWb4NEsIJTtr
P4dSHxiUObLmFewnqvjeycdwhfue9AAeR5Aj8HO1+QvycXoeFBa9vWiuagidRqDC
LOvUgbMh5df9oD2V8zmx4JR1u3z34NHdU6skfkvaoTW5S9fy1VK2i6R6Mgl7FjK+
ZDMSqHdA2GxCcia/uZzx//IZNpEkT1y6306iH1IPoINtjENDXJg3brndDapPwgN9
0U+qxNVTDuzO4uTmgRVJnvSnyVnz6ZlpqpLmj7AJ2O15vPfS3i7EvipIRDaf4kUz
VNVCQ4o78+O7WbIXdaNf7WtLC4CVqkaA+qiXQ9LSPdjUITQlcxi/ceRIlMjs2JIs
cO9gAFJOeMrnUcVAGLO+x+BiAKnZxXgsYlKlKVs4cozLdQwuujaGhn3Yxgvhy7Ha
8DhquGbZ4q70l5/aVtxF/jFrujZegtQL8+HAUtzPla/SAN5JewM4/JhOtepTfg9N
AVO6s9B8Z2XCK4Jr9vkJ70v/G+yWiooz8DCK19HbfiRpDrEj7I1wP/6FrmqWo/zp
HJreAcujrKluEB1dGpWZI1i1dZryJQ/NwVS3TfQqUNSHES6Q5FSGtOQ+1PdBa4ls
m7es3KhJYf6aqU46pv3kVfn0eBnjVUcKWi2Xz2zV/MJe7BWzSTghh/7WR/Q0Nyz+
4PoI3RXOGnr8mHCZZPDO0mzL7/G6tobEbvxqOgluVe/5bI+Rri7uVFEHllIdxTMg
qaLsq20kjS6oGaoqq/Rv8CusV8SkFmyLm2/gQhG8U2KwmKQuEf1iYXFhnjfMbS18
PyjCpZDa0/5X91dgzhn91mwJoIjB1FAum68W5B5PK/+vWzkOZwDp1KrBcKEbWHQ4
RDqSgyLiGHVe4bsy5/UcKum+lNhsfFdoQfGnreZPQ0c3p+49JQo1OUKlOq1JLyjD
OP6zeX4P3F+FRY/VdjHb00sWqspVfzQism+QvXKcxyzrvfOGycHUmKyiRQzm1KZK
0Fx6aMU5JWJXwUshZQ1pAcQuKM1RPvFkagJxaMA/14ISLILXhYlzdNfXa5PsPxiM
VoJn25yFaUCRsJu/8k5j73YQMjbTeqIrHmVRrh3Y54/d4L7R8Lum5DpKpaIXbwfd
mddAa0UEwa4JK/T6bHpeML3aJny0muEMtN6OnlUA8q6g8BMZowZoPVng8Ur+lzG0
WnkDlS8RBnFYg6KjutziuoaXC5hi5DFEsqiNqlvEqy1ntNLm47wW5pq8dZUXnp/j
l8d3yA84qW8fJDaNEwOBVL/qGKGKBR8cgMZPETCfjsNyxV18jwOzh8ucZi0LNsdm
I277poup5J1gayCzgAAKFH+6z8N0717Z5nIpG5nG+ohcsajDxiHw0PATK2uaD5Xl
ZLe9bVa3HQ8xd5Fbtufc6cm7jwd0AVMoN4+MMniaX/85CHSw+LW0CT5VUJ8HiFnw
TvMe0djIg8V1OdTs0Wc3injGF0SXwMI66to2B8UKUhY=
`pragma protect end_protected
