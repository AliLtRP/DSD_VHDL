// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
UG5bjEWIsKDQmjTDyp8W0W58fqvnhb9/DmAYKaxjpLVfTEKNCn8e9PaZ2yc+XMMQEAcLG+lDj/gG
OBAmOl957EfMMFQAisVopat6m/iSogbSDR1k4/MVnahddyfCv1MNjL+xyKHzZ7q0AOQyV+/4yMpF
xEYArAmDmGs898DjZpjnkeb7Xpawqt3Phi6atynz3TwD1FQMQLJC24fUAjYzZ5cMZsZ0aYZlNOjU
KLCCROvN756Dc0ZnNeodwfRaWB++xi+0FDdpgfip7SIjqxQsRMhQLGqSP/8kxiwNJn40Lgpm7cXB
CUIu4NcCOgmWSua0K5u+xnG4mV4IE2PsJNIiDQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
V4liLIV1SwFbWI6Hm9b8uXP7JqYr4XR7DNqv90I1jE7MeepYxfLniXJEqrLEIS1GYuiTkqsLHcSi
9SBRx8vPoJwtk35WXmvyJaq6R5MnPBaGRweIUI58Yxc8tt/dXkKCLOKRykkG744l4E2GGAJPthQB
EdYk/Sra+vLnKx9Tp3LSqjnaTOThTCd7G5B7SCGrvXvc9xr8qSYdmQrNDanUY67Eh0cJNfURaDtK
1Y7foD/dlZ8NcjbGgUihEA3/XFVHokrxan3GwSn/S/tD6/DripWTYnK+RSWA3lr2FYT3wB+ilYZv
bf9WKTvoRpzax7R4bYXgvsrA4/mrQJhlUu4yxF0yaNjN9srbHNqYZdW3OqUk/iwt4XVyr09mSLKa
yu4vBTbgEUJkhVjD9DiYIw4iSlCApsssIrbCKzHhXPWiPxlMTXuFzTy9DFRKaj69os3aXB0wC90y
Y5+dO1vrofSFaob9v1v8LB14vxfYniGyIVEgY1MzVzt4XGmbmOrl5kwDTo7Dwvh4TKTwUI0sCEmf
L76SQMQMCF4O++TM4u11Do/UasZqriUyf8D0B1DhMc+4KYGkDN24jW5ri5w3o9MQ64tMN8ba6rXd
nsTWUv9UUxL43Y8Aa8FF2M2TuWrwe9Zv6w17QxgbAVr4VxLbzyWgTfagHadw7N6m8Rs2YCLkG55N
ApNmsO2BXvj8cheoyw8uCDUnhmjlQvUthRIPh/Zfr0fPq4NC6HYnl+0hhx1FFC1kiJ3UN+L1INQf
S1lBh6hyddR3LskA/Z0IexFw65wqoDqDyaYqB7GmHADnmD6ICB7eurr1x015Q8j/BjulIiDjAWAw
LfVoph26BOTSvLdn2l6OMY3pbkzfjLKkRjBIB4R8LcmbrAkrwKwE9JMWzCWqcMzfAsQ61qwxPk3e
oGIZVfnfb/utGS+aG8JeIQ/q74zxXNburcwMPh37y4StDXGzeW9uOYYZtB8hI8MhgI+sBWrnUAjB
N9xEUuZOT5gD98H+ChPxlsRstZcpvBAWeRqvdN5AXHQ8Bc2SmUSUZ/hNO/kIbCAMwpwjRzUasmEY
nN26PuECaXfGsLcmKEdvqlepb8YxSMww3FjjtVgyz8Hbd9R6WVFSQTxH/aHS+uJhA8/lEJqi1HmN
QVNP481LzEsb+DH+pTUyqtaUlm6dLygvxVkWdqqIGP0aNeybziEThxlsej9xqxWmaN+DHL7Yxcc1
jL+ILzBTDj3wYGXwHETsty4B88BW09FXveLNe09efZ3nZckJlohY0WcKho5suG1UqCEbGR//ZyC4
nygPBnapUtUmdC0r19RA6W8uM7vZqfg+gP6X0Z0yLHG6JN31vkAkMVPrC7IAU4DhaqSl7HbiVFP4
jvM6Iq66vl6Ctsh13M1UcdffIaJlyesrt0WHd25mRYLUfidbdhO/ibe9nNpaU66ugYw4GgZ3CH9L
LJDvMqeA1gmcSaXlLQX7YDp8W4ZROuXyVnk0H4fCHHol4afwRMnr0pnMmcxv2eWxE8QdQVLQ0fHL
86Na/2bMD5B/dLvsMLq9iwpCqZ9lT8xUFbdl3wF9XZ84SaefoPaZ+idWMGZ8CpKzuvZJfZ6if6fD
doMgf1xVC5H6OZJLQQb4QTfKH4nzE5lcExWy3IFIo+R462BS73EjW45UcRBaWcoTlq9+OMF++Joj
Y/yoqg43o+3kHSHwy61qY9hkt++1Fc+2CaSv6dw4oHK66wA+EjouvsRIL4GOkhgcjVUK9Mdqwo7a
OU6gIB381iSgzuLyZHbAOw23eEdC/oDnDYdD6qhi7cypo4k4TWNRNop9E48A+DjVI9iwaYZ88A9L
0LNAJUoCBhTkyXaAU1HtdeMdQBsOyqyA8NxySHW4CH1z6RgKfGChEa9Q7Krw5djVB8mh7m3arvAL
RNoNKH0CyczQIwY2cIU9b3HplW/U+jrJ330NOo79rJngcU1YN0OrFD78fp6yh2mqQeeExd1sF7zw
/GUgwe7/VJrD0TeKd7DCJw76nUXUw98D/cMRqqwhlrRr7Ui8nEUlpBsPbh13KWVoKiEQJxQ4yK7f
9sVDD3R25JAVqr6QrzmjoEItaxtplt9rywxYEERN7MytaqzTEaUfv/L7+NY/ffCgpBNCYxghOp7V
HQGFZkUUTAe3l01fN5SKwomzCFZcv5VP6E6Eycyb9M/k3FbEVZhitDSteG/ho3BbxVc1A7MzsxY8
tACzmZwLDQxDHIA1cvRONB09uBs9UoueaH+YWWY4ZW4s0tlUC4m3HEBqPE92g2tXessEYkKNrfLI
JHs0b43xcTV9w/Jl3bSDWEz3st9krintiW6k+0NcJQc9P51e988Qv80xcga5qyQwuoLxoz8CszXa
pmK7ovlFWwx9X/kplPaF4yqADwCmlCQDOI9hEzRXnWkJPmWtXuWYkdKgfw4rhkYdE0YIfPfnS6nT
HP/jd+X7cjE8RSUbLwNh2Sm9XVGag5uq0QfRjtr3aZt8rzcdsgJXqYk8+huZvSQKT34bkr4YKgoY
4xhCCRnciLGJHnDps9NEJwSuvSpqAkpiSppsBjtKOKUZ4c2+I1wLdkLglIVFrv+1YOd2A8J8e0Tu
buiJoDxzXwKdGcBsnr24L8nTZaXCbl77yxhqaUoAVi16tD7ZX4Eo+BGgw0yTCOhUnRGYf6NTHirV
csuNjzsmMsVowpwMKPhbufpfGbUYBopvPo7clL3LnSetHAmg+WtjIbBmuCB5P3d7p2NFbiB04EMN
ya9DBGrc/gXlJBbAShjfnO5kIcL/C1IBVUPZYRv9UmnQ0KnFs/BePkams3oNw4uQp60C63YjFdn9
KEfjt6n/MLQjHwhtvnyCpvTRl6p8ajKA8zbWopF5E7eu3diLnGLt/zax/9WCia38In6uYD3YOpVJ
5cjGQhoU9L1BRkMePqdoJIsA2lyf3cgccy1oqYeWASAjl5Eun5M0AFLDowYD7S06qTKQx/8DJuUq
CfWFO1rWnv5dJntfBkvWDssCBmXH6g9sKDm1xlDEU3jklQKtJFas91bTbSRrPai4QrK62AbL9Rzx
iCyH8LC8lLbguzAEZrZhP0VdCQ2Y/X/DbAZniOV1FKS8vmfzwSFh9IQHU6KVgqR8DGdlNDPza9aS
Ff3RdAzfF04tuN4VeByFcuFrbDvdz51NuV8F4MhFz9rbktgPS+81AXXIIObi9snSQil0tIwFIZF3
JFmtWuogmie0PBFLDlnWMvAXZJCaOBNDUU7VNj7MrLV3DMZD1u4bk1TRFBPmjCK1XXdnOqou4Oeo
Xf5/0l+ohL+WFHchcFTBt7i4u5glua4m/SluM8s1tgD1VejFJy19T5Y8FPpHK7CllTGyAYLxe9dC
yKt1LL5+YP19m8suKEKWbc+Tr6mmwRtfnrwk/L0w9epMzoS+iUjYdmZYwBECxSpe7ChTNSI4zkSR
Jf7Z+uTarXmK2P8AJvtHJeOtbEcOF4zQ8675pjLFT1A4JkZbOT59c9cuSyZcrL2r0F2igHuLKECQ
RArEiIXwhq0dMgli4590U8LMdjRrI4Juv+ixYldlnuUjX7J9xF+p8UYaqq0YbfX6KJhXED3QR4lf
4QkvpUCqSwe4VTm85wry8dCLE8AcysImZKDomXCCpPL8kN/PbUIdtAPXT0VnShgxVeb5YmgezUO3
6H2rw6kZW2HyN9R8aka0zeYHk5jx6MVQSpEDj2gcLwL+cNXw8M/KUYrUtM9Sy3kIxASFIf2yGiyY
hrKjTOv6DG5pDlnFxR1WiPQN+AVWTlmLDDTsd++4DHo8tskpXq7U5DDDcKfzNDFiFgHnCqLmeTib
fVm7TQx8BV92HZSSs+8f5bd2uY9SNZkhuNN2lGsUHGPnpNK//uos9g2XIbCzDdV5/qd+sURc6pUu
J+pnzhmlBc/3Kzwnx2oIsPCIheBdcmmTJ7ewuJUC4K7Wp4gWVxJTHMhZRtJUoQ1MKxFItceajA/u
olt1qP8n003W/lQXx/KXE/W0p8SlMKK2JPUzYsXb36d0fZw10FUO/vEFfamoSQqgEJc/CbU+djEQ
quxvHqxpkPcKHl6D77N6CMasVxRSJtH+vFlzrHZ6I6IGLR24wvPHLXxIA2RwN0QpW35/nYAESXul
t/VtS9xA9O6jRlQn6L4FhlfUKowppL0FM6O+fRTqQa8lAAPWHIO7N1NmETzyQgIyJkzdG2NqmGS6
WzC+JEeEllks3CG1nGT8QmTPb3wSWp+nHNbxVSenrceebcRQJ+VPIGUTWaucHXELY3Uf1qKI28mX
SiROGrUYKPcg+oLG2V/T10KNV/Hlj9sRHS0rrmRA0wr7eG0YbhvinVuOpjBSUJgRb0S1q1yVORwu
ytJljMig8St0GLoDLmerkJFmunQJCujCBlHZ0+4fyotDZa1G68HLaGg1Ay5OTBb6Vcoa5uFOLxdR
HsCEIifRY3neNQJLkHjbNqpYyrYqopvMgdPcDQrazCBdqEEPHQYYX2s06P6TQNiIM6N7GyCcoKif
EwM0N3vdXEc/ExpxupWwq7wuHkKAKaSRaR4mRoxU/FML/sGiV9ee20OU/guc/1ljjfONnyypi073
0CB7nGe4zlhDe8h6Ljc8QNreMt8jku+G7CHgnPgm4sddue+aazXNqTwvXd3boZN57O6Evghu0bnt
Vl3fPiYcU3EQztT68XyTJg4S7LTTUwOukAXNdZJZxoVh3ckw/wrOUz8nKuZ6dFzpduCWAZc0XNBb
7rDxwEsFEaB+UkUcdFESTzGE11ITC4BXSMZ4+/KINsWcdmTQjUlNmk8oZ6HggSsp4HOmvItvzLDP
BRrcQvJkanWj/VTGD1BEUnd5Bn8BoLXOfxw/I5/6Ib9Q9VDwJqjWAnp4eCHUEXQZTKjXTi3fuwGr
6D5Z2BuhY+mF93LIIVF8Cc3yHGI5eXFqDVM/xwvbvV9QE54aW+wcrW1qIHjqMD/NzoAWzLTFg1/0
gQ5b3wFLbuw0k68fX5epBmdueOsPBgTG2m9cXu43DUZ1GVqeNdx9qRuuGKxDoG5DzqRPlLLAvwuh
c3NZvhY/o7+G9kY01KfFQtprj+Demnt2Ujvx+G3XjGW36lbErV/58dLD+R5uad+iA0g3trcgUD0+
qkjkAdnlW9YpF90P8kesTi7ODvsNma+bMDNfC1Lc4cZ+eFy3i4AEjbdUt5TwI30yqVqUCmLOiqiE
EmK7JK7njbhRn7WKFyosZ0Q7Jl/7aDDmafXf8nqmmplWxSdrAAVuRoCIRRzu1EFZVpyzrrl4sJim
mgfq7bCQhgt1SSHMx2Pbou8V6jz6h5p1BUOxNjOI+16mNjZV9SAL2PHhKTqaUez1yJh4TwetNcPf
qw+hTtF9oOw0kUa/MB5TFAsIaThng2Z+boCHHBj87hf5GLwfP125ZiTZXf2HBn0Ka6uejvrvNLyq
fDB8Lmcy5SGIwJ56hYKA1n/DHzld34E5eMNs0QgfPHME+XTo2yZH31kZfELG33piOgRU+g2jngJR
pe+HO9ThHTHTLnQ+R7M0R7CrNKVoPSbj8XLPLUR3zzx4meH5R9Qe6nAlGorLEcOc2RhDVG7aYSye
/H9TC5cWlDbBqbQrO+sFUAaats3jgK5v1wj/EhJgL9znWWoKTzP151TI5Cb7oz2qd3VGZFnKRS6z
Fgat9iYT18Z5+Dhx9ahdjkDtQxfKnCExW/rT6o5TPbnMveLje714WaRXl5e+LPoMGwfo1hxyX5US
Q6bcCFwdGqnyHK1tY0oG80vpm2adeaOGyzs51QWnn59fFPoyXNQAA/IEtvEOBKTqPL56Q/dhX6ZL
ycMpbNnCs90Wjp/QcKWpEawoXVw3wUm7U597OsUeguBZnuiMMBEY8mIBkXTuNCpfWDNXNTtsFdg0
QkuFB4e+vODPzx/dKD5XU+fVb2/gwB5vZMGCZG4tRYi9AQ/0QJenww0CUNqTJOBLKlCVrvVs0B20
RoZ0avQnsAFGrdCF9ZG3HeUpP20u8/Z0b3ntDFnulhEghFXphwo+gOIdPChpy9ww8lvRQymlSkbm
HTjJlj3LABnVm+k5ZBJLIrGh9EVVMn1v0SwQdUEB4f03Rby0NvtR7IIPK6ABTT+HAyZGjmFzPcZH
WWhTZwt8y6WVYA69Dmd+y6n5RAShCQzURrt4GAM7I+q+jnBVRE2rSdaBAB93osYjG5K0nM6CBhXc
Wy7daxzWUexT+pXx4AbakLIKWkIb3HZXT+ov6ZRI1UHpPBbTVHO3VbMiey8/6jKyZV3akjOAObk0
5sYlDnW/B0MnGETwq9jhcv0iM72kq9j23DqWixHR4h4FOxSUDY2Tl3WQpRm/qOVMSCp06fdkeQvk
q+aAsy2cFeHid0KqPJ8rWhQJw9Lr+C1ezko+vM7prmE80YG10afY6Ugw/nwiQ0gxtBCDa1H7APk4
BCUT2zoav4sPnUPVi4bIihbfZJ+PQDIcto4k7ZUX0N4Ogc+7EMPICvT9pgCtyMVUt5NW1bu4hvky
GD6JXgPmZ5dlwtzIM/ErWKPJz6WRKEQbic2wb3Jtq4gSBmhos469yAyKoQIoD1w6nVDZSmkrLKk8
ckcWCfd9Akyy0S4+8H+nbIwBrXT5aBAfO4yu/TQBXVG3YBIn0N6Be5usCVINBzXpiy/8CG/lQ6l6
QY7UhHN+nX845wG7pfoKenrcFHOl28RzWE+b/+XC6Ai8FRWh91RLSUHIYPOjlfdWhHdJoPyZSJEv
5ESHGY/0xXWQElMKxluiqfFeRuHpo8Qpn5nRGyhHxRWH6xeCvRBC+budvUET3D+yz0uXXykzzzZG
JhXzYBJ1DEKws52DCGc33jkT8p1OEjfkN/kcG6y2kSquuXf7mJ/Zom2lyBZLpdoYwz9SSvJeVsr7
P8rgAMncAVcKml66t13jcU+8EDzLReIhCrblEqmCRzhkXSV/1V4Ybk3kJQP0jucNxYzot0jLJtPW
4aMH6NIqvJivRPzjjq6BsY+M9mcSkWiU1q/yond/mf8nHPtTyxo7dWEV03WELSHMYVzTtFXuSHj6
YSb9yLp0EgTbZNOGpRfk5Pc7ez7QWgCGPLkRWHhqkWmJ2EXEIJBfI3jHJAWlODCSf64dPxX6x6Ru
UawR5urLbQvfC111I1jOGyeBjLc89fDrHNUxlasMDxVIIoqt4NGBou5Mj4V5hiy+O76d60Y+Q2NW
s7He8+2fEGfz2mMv5rPzYEFvOjHg8OLh+N9n8iBYNqRiIHKZnfyNlXDf+sa+2PuCpyRJuI90VuyQ
i5J5mUC50S5ChiDCBRfn/kHypFcAzI/JtWm2YQwtIsmaL68++JStpKBrUDvcT0xPnIocNttcChN7
T/Z1AaRI1t9sGgFbYDp+Mz+vQslnIsR/k4nOfhP7p1U6VXcaA0OciNkRZzBH1m+DLHdO7vCnDFeM
r7/Hgp/JIv+TK8x32VS8G3kZyp3Vb37F63p+w0DC92416nm3UHv7s3OlITMqW8rBxFRL+huvhH+t
4f/LvNnlSC3F0fdKlTpUwpdqyrZfNNbxkjy5DA1RzVjrOF3Gbbw9QREc5qY1voBaOGz1SV7GK4j8
KVG5qlJjP71Y1srytJYMm/JnmGExWbDAA1+IXEgYrd/Y5qoS4+GA3gJ1abwecdt2KUWp3q9sLhta
X7N9y66tFDFNI3fZHSBAzbPMZvYb0W3+8RvdR2AUdcSxJoWr49QelEKjhjp8C4cxVhPV3Vm5XFBD
Z5d3L+a0tazJCsQu7M6KvfODY4QbShkrmfebds7AB4Lcg8WFup+Z+O0mj8jKJ0fg2nB1y4yZF3cm
Mm2NK4ACuR23HS8DCmrCyCPDWPtg2Hz40Ytnbsjf547fZ4iByAUzyxQMl42GlaiTDKXCN1nPltqj
MEhH3aYQGKoyjynuq5ZLj4ssWV5jLFUSfUIfWDAB0pqALSGx76sqBQsXgpJky3Fzd4pToxNUHn04
EVghG0I/sJHsN4BVPCWUquWp67+zScVxRi3BLydp1HLRTg/tjKdhZ9Vw0IXGoYnlW0sSkt92bMy1
iYGnApmT4vGBhV1DOmZd6Qo8piXA+jvnT0JasSTixJJGUZQDAKcNNWCneXPS1AQE8kMbe7TS0n0h
fudjjY8NMH9kFqyg+oGkwyoLpcgvo7ArhAYTgx8TcNq9u2bimtUoxe7J23P6azLP5M5S2yv8jN9M
M+QDzCmSS5woVJJihLAzXEBKJVPQlNhus1vw+YkcBZzLBljqmIWGu1IANuuMRgPLU1ZWUO07MT5G
ycjOC6t40PB9ewCM7DExMiptPtFJ697kG7wel4GKUmP9G8hd/OoPqosJq6Rej4UYC70J0m+KTjxp
tB/vLcX9CVUxKhTa4sSsEbGgJbxcOnOKZXTeU3tPlUIdDibLrE2HQlxBZTkITTnvO9O+UnmyVUtM
qInBLcHcix82+1noj6XobmagDPzqO7t6FfhjHEbJoimo4aMJfpt1xVy0b+JFPvLz3QFjEdgDo2Ti
O+bYoFaEcx3KyWmfisH7in/JJa7k9/RXj7aNp/X5ev71MAdOAUdJgGGuIWkgQnTysIxf1AdTSFKv
5imjZ8cefxpXai7IXYKD/GenoAmmujqoRGV7QRXeQOUolWlNidtn/wLmfxvthoAzNMY1xblXVKiq
bG+WiYzSL1puirssFOMOPja7U3ouwvUr2CwNr3Tg8mgLa85RtnGN7cLD0i3CsEeDsX2aGj3QcE7q
ITJ4k5LU67b+XP6b3tK5JoYtUbCq2ODStp4L1XSgnyWo/gV2X1hbClRoUaDLHryKWoMfkfmujxvn
WDrNwN7u/P9KZJNrFTST0EFnj7dKdARMerYuxwMqSLKzJP97UKYKOMmI66lJAapaZXwKYP2L9F4h
5ct/Hgdztha1GoXcGAR4Xh0kNM6jX8IcoySANNItxhg85Mr58Xo6fRUBWdbyUSVnn3F4J0AII9jb
cquigpWuEI2197Z2DPzP9G/tfTCFm5mMDT94cRJQzAGw31nbXsHzJOgWyXzsCR/aixXvF+Suy78L
WOW4H4EvCxwni6yigjX2W9X0mS/FH0gC2emA8pNlp5pvxuYOQhqqBCe4pdVjVCMgs8zpBYnX1EfO
lr9wb90Ecc72iX8HyjNezYoLUACd6J+OUp7yziZ/ypjU5rJ/Y7zfcStX1KMNSVJHJ7F5JtKKBqis
iFVU608FGiIQwOROV1elxoskbBrZuy/KRPMRwhbmMdB81rz2FG/XWFNaX/s50uhAtdlvPnJlI2il
PkEHF19xftD0469jtcrIbpMx9GtUNMIe7DtCg1TCTn2t5PsMExW/HDqZXQZDsmeHrfkOQ2+3qKJ4
EFzjeSsNGHqFdx+sq3zhWaZ2R2FjdwD7UjfuFKDT0D2t6hmSbcoLah70yJqBiN0jp+rbdBFHllu9
zipltlhxCqs7dy/OE4u3bLuG7LjHn9VvB9rkLEfVI0rBWy9Luj9hV/VdpE2tSc5dSUad29Ooh9Tj
2dFlSXbrGnyiEqYfNKTEP3XDF4WbprDptQfdcZECZMM1ifsHkMRRZyj7hQpKyhuXpYGDs2KOVBSR
Fo5a/8T2sLdSJvKkvERp8zO4s5y6H8iU/uiFsujuNYUf8RFGYr+D69QKV/kF9G58NLGQ2fez+Pyu
gsfVwsakcE7yQUYTsL8DjnFoNAiWuykQ4LezijKG+4BQ2W08zc14QxUrHz90++Z5Upu1y0v7dtty
GkaKSNI/DKjYD3ZhmUfIrzZogQV2vNxq2aKhlWVXwDQMSestFK1sMKEjVmA5QCIz5Fg9so1dT7or
YaDMIjMbvF1GjsGpz/L6U3U4bAhN9rPZF7i6BzozbolWhzp/edqxQJ98MUTJo0+dN3xtvPIyoQT/
eGc5DrtrxeCM7HBi24MH20ROJF0h+m8OSMmEhZdTKfDvAK2bMHXzlIFR1dcDd16OZt0MvPrl63hv
iznxX6uSGTLGjdcFze3mdR4Udczza1urBdIvGRwH6fHfWsZ994snspPlsWC99MO4qHYFIoyTG3sE
Stkqeu/hxTfKjNfdM/brC25/+o2SGNZEt+My+PsoCCtGiUZloKHviCZ5HXK55VPKlYFCkg4Qa6hM
5t7pggYeGNvuvngJRXhLL1ZVHzKxGXObQT6dz4OAKJXbXpa6Tvn4XEbzzHjae1SrtqrSK6LnMIXn
vmKSnCkPFQHfdv/m15xcIdKH3RA1USguScVKZJZjca+FQokhwDiKW9CHFjGB9UdDXIk3TsNU8p9F
mY/7ZqDyO/MHBT2fvNr9Pj6XhUjkuoQJ3eExovFcsDlcCXCwzJkqjC2XFy9/xMTqT5WiAipZTvxI
1SxERKTHjm0kMZbeg5uxCfZVJ3NiQ4O1WsCTFL1WlhDWsbGisX+DI1Nw/fLBKAxpy9CYcU3528Ff
NNQHYEXLLEqVLhtxEaXGf4dUtSGgLzMq9g+U/B1MLDLWDxXZDNe1DX9XrMGIq00rGeeBa9nfaIOU
c1ncq0GQS58uCflN40otecdcUjunlyde0yqTR/PMeI7ByI+/5maTaae392cwaGzNmeFuPY9M6Lhx
djLIG6pJoVMS7RwHYF/BZgYWtYu5CueggJ0HXil4KjkQ6LTdXfKEzI6a/13EqHt1z5jorpc1evi+
X7TLHwiHDQWB8AS+5rcgL2+47H+3Zhzbk696bE4oow92vbnO7fu9T2OOqCLYN1CRwEmRYZrSS45I
Vao2ee71U909xBFB/IvBOsoNY+m8lCeGGJ1UKWjvjODUEPa5xW6pbRkW+LX1tuYLbLl4yoEWSsrA
oBn9Vyua2JIQAuyFK8WYs65bjeWvQHmDfe0HQdE4YovRmzFOIZH+3S6Z+Nf0hjYWKCIB8npcxNge
nW4ld5GczF7EmypFq62RX//8emJO19e+lKIfH2tPNQ2R65VOGzQEYY3fwez6ZlkXzQUUp2kD2OU1
PNLVFthh6RV/ExCzFBw66VWxoXv6EJ6vtGw0Q4HVuRBOJyhMjkVolq8b18UW8iu9kpqpaJSDWZ4t
XjIAMvcnET3yw88QM1DpO0SuwhkCbbbTqILgM1oFroFRp1nEyNQTXvePRYgQmlH89w4PjJ+vMIBC
VA4Ffab7acAhWRJ9OjHgZiiqZHUtz+Hk/uDZ+w05X3TspNuASm/xkyHrrp5QnyTUe0C95XnXNeR0
jjGaKWrXg3vwDyXIn6zsPQI7ywzt+/RsCtaNIwO3iwJyGJbQGvSvPwrAYKuv8+6bNXSlKFC0PIa9
yqhnNBc4Pw6oDXYlb6KCaYi5/Wd0d0Yd9hn2B70DFD1HJIxGS9VvhQzwohIPf1G4AR4o9XQvXv+M
a1gPxQTpbPQx9DznoEg6AXqIDtItmSwdNzEC4m9+miwChyl4zHXADQeiEUGI3sL5ij8mAIbqjQIL
3CWpWp5W1TC0swY1lgdpjBG6S7fGVevscaf71WajCjvX5+XSXoCBoKT1tqZYb6mu+4E8L/7+dpv3
kfZMSieuZrm4RvK7gNX4a1HXXCa7Pqff4xfXHeYtDtjlrk3UYLFa3BlB2tlVgRrOhV2b9tNhejB4
/i8TjymsIwOaz5VRi4MX1MjqIPRq1n1YXjPqm6kOsoEKsQsZduw+28eesgTak/M72dd/rsRaau4z
d+FSSqwOUNvof43xdBH7/k04B91POSrtIHgHBAIyKcTqYyCp4psSX7T+2qQh3O6wLOdbVYsv07vj
L1QuRRvOH5mQhQkjyuWp6D4z26QEvknGJcOusgypwQ4NP8EKn4zDZGCxARM7so/l1zj1irfg7zFe
k1NFKsU6WfVG7qFLCrCast9kBUAKxsNlbFIty98xK5GdfsX4SdXuueETdQTk5o+xtd42ieG2Pblu
YzxWK6BPelI0Rzz5qH127thKPweHIqz4yQHJggsiFu2BUUl4ddc11CrKsg66gk13n51Ub8+rxzhA
nAIkWtrhHms92mjpl0b1qbQEhPSihsv9BDGHXREU1fIsAn2BbfvAhO/Tr0LSW9NX1VehutZWdpuy
Dw66qV91ecDdAXKvIHNK9TQS1ATUdJoEOOwGdbTsurVxaMko25KMvLbTo6iEJm8/Q8hsIsJ7ALG5
D9IZBytdUAJNrsDdJfNx4xsXNtJHNP65nv/O21+5/9mZFetVm4hFLAx0suKXpcgabXKj8sTC8jsy
6pCjTqmGoD9F/YPS8ABGSgIIIN665gF0jhhmdsufWBGlqfq/0wnWyrro3PdcNBxKeUxjHZDBfENh
xcVUz/FNr+91uxlxqevtMDt9BXioSv+5UkXOTR5xkgAP2m8WkZoEdWdwaRMjaHTZ8zQFulP2MdG9
l0s7Lu16AHVWwjtiAXLHyEwSiu5ouVfZCHVMgm1QbD1JRsxo5w3JbtgyA8w+TYMB74XDhLCkNSxl
Gafpu5QTRN3fLuhtnknb7YGlCASzXNvUVyUYH2ToNzZ5Vq3+E5OUiKf2yB7OGhhZTYp2nGAzkOSj
2iZaQx2GzEa9v3MdnLq5RgXGbKfBnE6eqQITDKdzRwIQ+6POFfr2EBacYE++EZgx4++8dzcxeasO
MFvKh2i4cHmTX/c/TZ3gbzL0N3uTpai502QSmU0w0wkvs7gIfJxhmjyeicRPx+q/1+R80ou5qnCe
cfzuEQCwvmHSlRpOE3q8cqz2YStPwVn8SXEUCHeTykDAV0ns/XgBYG7AW+I1diBhT5fHDnU8Wlz5
0vzxvN2/3C2GJRSbjZzS4BM4QfFpYlvWB3SzIzsyB7VL01WO9dSUK3VDYNN+D24Nh1XmO/j7biZe
yCNIUdxtsXOfH0s3qmBNu8X4F2Mi5rVpSY1MANsV2aSBjOLA4zDMeMYwKRIbetN0IrP2WRCj9GK2
66F7PqLkapnu/HgIgHGL3u3oIf46xgV7a4a3G09RJlo0NFpFknQdzI6W8iQ7EisB6kUIWY94YKuA
eran7rCGkvu/d8W/GsgTswXRbUffy4YRDHxfvb2JVMOuitZmRSixqmZp43dx6sHMWmhIDS3rNlFg
m347H4Chiy7N66eUQdkEouDlyp7ErrECZoYicPswE0LoMHANmjZAG5Jcm7xIRlBXqGaTu0K3pu03
3hGOwww3gVYWillaCXNERc4Hl/UIjxL37tjxn1ALyPRQHNzWSCaIOdE1WMSXmygvh/VDmy2uZ2R0
89bSdbO81r98OMJf6wYM5wqJSCuaVobY6YaV4hETE96vGAe36BT8NWMOC8dJKu75FF/CYNWQdRhx
B0ZkxZXqqMREKXXf070J1ATZBtA6Ut4Uo725ADyhxIa9uCfiSKAPCO1OJC27T/+OziKSqzecQ57E
KrclviHGL1J5wSyYi5iRnGvdPlP7D94wh5buRESJP3vEPOlCDp4sXJNzaEagwYiJ6fjxBYa+1OR+
JEB2oPzmIOBpiE4RqOp0aC/9wVsu5b4Z89DCXAGQfY+u6xSIZcU8BkKUrCcGZ7Iw5+wMLr14hDAN
vzpPFu0uQ4sr6UCAv3R/2qb5pUIn9NuXp4ddzmDbv0c9ewK8jCV7ZERRur7iC7Tpmo/dLBz0xrEq
F2Qq/7xEc7S4P4BlyFifCH/asz9KcjwjNXm0k2tniIKQAnb/hh+/S6VRYxsdzQjhr431OlkbWuPW
tmT+PzZ0PedyjOAsuXKcrZ3szweW/E1YsMVDhLcm8QFru3AHpT7Z0jDASaU9u7oQ0CQeV/Zd2lor
lb6NaKo851L/QQAGQ/EedSirrMdZ5dVcTJEIusRbTmqI5dJDy2iPU+7LW+cR56yiPGHNJrusumqj
q3WP+UTIRj+bI+S9SdB9x5LBTt1uKUByMJ5y5VfhAPIqUyAve8XfwNqzfCZqf2H2RL2KzO/CvwXM
2vRWbZmDkN3XhnOsYFQ3xVMmN5UgoUQC02adBrxx7qG3QHsDZZnO/fcypuPfVbsUCe9LmAhEUwCl
3iG9N44nP3Sh0NpK8IaSnRN1Fhcga1z9whtFkhxasFVy2bcECYa9wletZaysvXTBdniq35tEN41z
jr8te2VvukEiMQfm51Wvy7f0AyGDsHdK+W4+5kMN7xL8usOW93pdC5ikJ5dEPKtSCq/O4IDgQads
w5lhfcYf9FW42d83FGSYNkcuAZpVNzPx4Z6c8irpXqWqpO6FSce9YACixuYb/CTtNUc5kCFGW1RW
Oqi5mNsZbAxA4thwyksePizlphdy4TeoQ/1GURfF18Ta+8aeI2xucSwUxf98v7p8QxlwUAZW+FCJ
H3HV8CvSqSeqXoO1UXi7sL9XPVdxlDimg6I3jajywelcPr3VKDd9VJr9DF/pihABjhR6FdXVbVti
cUwEo+9a+pS5gctKRbI+FwgBwWNJGdyadDn5dphzSN2syEA1RUk3Y5VBHR2KYkPUo95bDrY3iwMh
Zr/5YzB9po/POG1ShUZ614TpA8Es+mgE/uE6q9S5D5eSkZFbl+XZXXBMlPwkxak5vgStA+5i+TIJ
XkxS6EGYSGZf9tvQfkRiSVNBVfolmPGUOTvdWtcnZMmtuAnn1YNxZB35L2OLDdti4MErVQRW3FtN
nDwRsbLl5K01iHAvJ4nfkOA5ZJ6kvGZWNyuX7cOaLwIY/4lahdXcRrYfgzsOpOxwOP2yea+B9RNa
od03mKgTfYxuyWzSNUc+hIwXx5T3byldK740gO+vn4OTJNvAhetY/7nTCCM7V7+bWG6ft7Dj4SRJ
12MTfQAe9TQO4go6MxbvQZF+jYa2AYN/+6YziTDQGccDixYbKOj4EvbDo4HApAeM17UWLh+I1fre
92+g2KTI5ZGaHV2xyhUR2Gt4za8IUsJr3yrE/y7d1wsp+P/pPckdhEWwLPdItSQDlZGXQJo5b5hm
ZUvydob/940i+S7Jn+iV+MsiyKVXglPqDsiQ882JpP1oOZ4QppB+vtHFd9Qopjc2WdtYOVmnmh13
LEwmyIUofInL8/I6Eo1w12Na00ivqAQ19MXsTL69KGbU/nDNGiMQKbjLwCha4PFn2HUTtKjg2VVM
0K02ogybM98jsvomqniL/Dsz4DCz39CdNQSOlpvbaYyix7W/sjNpt/b2P1wV2J2fiMn1fIVcdzpx
6SUr/1Ycxs80YvZYBAgabDmF3gcYg8tjJYRg90v9XUxvEHvgF+WM/RGswrFPfKb+kPfpuygX5RCf
LqX53ZBiWcdx7tX/hV5wX/m+u1OLGt8Iwo63QsN36wDMfLEwd5coQmtagLfHqycdbMcZWl1h66d2
ZvF+H3RFVUiXB0SYfBV9RuQxfEvzlpf2+72SJiLSaUO0iiBo2fWnUUPcw8AGiHR6rmVXCo05UqU7
iQbZrP+sgRtVfZSgW51P4sPAm8eHRYZVgq2tugCHFgdJh3yXbgh0vKlVRy6k7ZqGwePb9t0qByhK
WMjmkfR2Ge+xmFZX+W7s1HxnYYKcG4afpLwPW/5NHIq2ew4uZHQRCaOmiY5OYYMp27D9rEkKlNlT
CPbtmkvOnbtBxQFgKkyGVURbywh4JfeQTtlzbXuKozTd5GX8NZI7aOq9MCyL/7TXZcSUTuWYghhn
WEzYHWEs7o4bqYOH2f8v/ENEkiV1yoArjHLm1uKSKcmW3SeSWrMcqGLnTHiXbGBAW8I09F+6jR+k
QuU44kpTP8yHgAKRyX6as3mC71Ws73/U9OfYsXMLcHRuwZMeGhWJP1lzXvZgLCXQnhTr4hxz4hbY
eNzrhciFRffo6zhqiKpK662wmAjnPKYxXPbBjSUxlGQuNnJ1SXudx3HL0lJvE+gYPgl5Ntespd5M
sBaqApCT07i4b27IcI5qsKCBj8O2qZyvUqxkxVCixKVUCeJXVhRzAkxJM59+pCMlkhZ7z/Bx+h7U
/7XJHcTUopkiQV6mJrHhwy4TmfM/qjIH781RvNRqv2bZSgLqzUsDK6ScsRE9AiYSgeSMv2kZZH3o
XIqoBh0pNw/PFj9l4kdPnByXbVEr9Ftup+Ixe2I43vaTIphOHrqmNWSoZxAF2xvhiVEkXfDkonUX
wtZTiJk66lC3rtKBtaAWwSk0MDYJ8KVZHDTYx0webQJxUP2PXaalLG1qUkMEPVESRrkqTHIHhm64
i/m9BLpengUbn6TTFOd65DdyYMyMUXyT4YwZBUXlZDi6n0uTSd0tsmop4jOPe+PH527ZNhpFJPOR
W/Ht34oEUEamXXXuMHIlDNsC3mJ71kYYus4puHxVFclu4yO5zWnJ+g30/rQ2KJnWaYR3EyGvf29a
AUuHmLMQDSfVLqlz0kyCb2YlFwit0BHuVHF9SCPZw0WqqlHsX/00JfcT+rKDzx2yD9HFcgxO9vFl
D0cds42hqJu2oVj5/7UzgQycwdSngeas7FPLUQwztdnDt6tTc2ZSkHNKhksPH5lZRmO4/ZlaD0E/
w71le+lEreBVAPuOGYebsrPzU1q22STnBWWD0x8hn5oODHHZ7PbsY7qdiqES0XlDaV9xzN6dCaHW
SWc/sy1y5xnpVtjsRF+2APVZqUV7NTjjXMGEtoCJAm1yDlIg+ndnObzsH+RP8EuDwjF8HeWsooef
ykujHYPmdFINSJY6C61dB16l9RFradEixpZgcQoh1dyLhwEvRz3xwbaGCIx2P6NEg8D12yr4MgbP
L6wvkNyQMPrZybd4OvGMuriUPxp4Uxg7Lut/ROGjqbDYwZk89iV/2e13btbMK+ZRdnz7x3Bm8TIO
0V93ioS7xln9lvkF/itN5ixS8QZZ7fnDhNedZxNZScc4+ozZUHQngn7nIKWygMkZb0mR89TJE4KD
usQqWa2Y/aFeJa9+iBkw67h+xY0uu0c//Lql8xjUOkFlvrOaL23iMZbeV70vZNDmQQ9BBr0sRj9e
QgYre4cSe7MyuC1TQRfJbq2yp4BVzqGGMcAhHvjqfR2USDBkCfp+W9imONbWBBp6LB3yBzPC55+t
Kpr3+tFkyly8VLXM0XsQ920XQMhp9g9kwds8bD8+XkE6JZfW36JrJ4/m8ZGRbfTbW/iIH7KYEfDX
e9OrVa1ks5VW13aavI+o+NV0+wgdISqEQkxImObBPU27dodWGVjkKYvcW6m5JGx1bPKhxkJZipj6
THeaBrbUSO+TUelqnXhJQMRaBbUeFsppnnd+eIPZ/Vgr6A2eW9/E4smLDUvUmihrzRqpYPz6CSAI
kfqyNdmf91spaikcNz/THEU6ZO45EMv2/2DnQ6MX4uzDPg8DCc9BVQtuv6RypDhc36xgWeALLQsr
inQSa0tYlrdWsc+MFQ3PZevQ/qdqc+YaDemJYsESiy5yqfJETtbu06x4z98kmztzYLBZe4m3FM6Y
pc+k6XwivXfsu0v20SazJv6qiTTJI7uVTx9uv4tn0kDnz7sinlf+h3BNB1Q+TPUhGMPGtqjWxZPC
NnElauyVPcMu5XbEw6cuGWyVudAzWUkllNU07R5TqCrKnvvtWyT0mmsiYQlk/nArnuQIlmh7YrAQ
suSvZQdzlAIzs78PenPTYyO7VWiNtwVG5x6pCDvz4bt3wA4focP6MyVmDkEf3poC15JQkPGyg66k
PgfVG6EHA3QSaR+RlwQk6vJ/RhtDpzFHX7Fi7PsQgR5MdSBwJRLN4UeCwXX4x7VFH6Z+eAvNcuVW
4EZ/4efZR6AJlzYiBt65xr0i5y8w520KRHRl+x175Qxt1JGeFUzIgXs9cfurWAs52cFIntXSH98I
x1pcPYrOJ8+kOm2GAONLMh8dTa1oe+e4VpzTPr5lXIbTHgvQIqgtYknBNX3mQh254mdhkhghn6RL
bTp9Y2U7I32U4NeOPRrSa53evZcjTe1Pk89XdUeoPwl+ZYBYokyzNKrEmsKQf1IPFkXj2JjH/9Xa
9UmuWEJEP75SKHTWYY8iIAXOu/LNz3QzJXMHFZdsQ1I77N3zDxWVsRiEFHs0OZ2dmOilGXo8ElDS
IwbKZvaY0Ax58XeYlH0mRVx2EamlCD7x8PoHmM+rfRi2bD/ctIojFBN+OgTouh4177vr/Wh4OyXx
vLZrcAVdw+sp36p1UW68R6ojkS3V+Z/ZDudFiqIhfCKqvhDCpTPLjRBPCgI4EkpsiWZP/QSvb0ec
zbzK5hNtUAsLg1H1UE0o0wpzoutKRroOqChW1M4+Of+ehiBFQ9MKQH6Mbywp95uJtLxq2QhDJMER
kzIpYuCL90NhNnml3Rl6r67QhVSZrBBt6xHU0UdO8x3HbGsBiFONKvIYl5vkZO7TIyEfcRbF4OFi
SZYraVhPWrlL0q4SRGAT+Wn9IrETWWWNHaJJMqR9xugJojWzzpgDcexNUl27GVLONgVCUPyQGHlH
F/QeH9PlXDt/LOZJmmp1n0pTsIGQt1DTIt/u082qJzoNoEyAqS7Qq9X8PPlA1LzfdVd53N4g7smA
cy4K7+ToRm+i9Un/x/F+I60uAUxj04bYgwkkSpUeTkJEV75mQXr1NY3IyRxvLcjTQgE2i6Olof3Y
JG8mJImUlOEDGZpZX3EUWBmAZYuxr1KGtWOXag48elIwZhhnveVbpCklepok18oigSxnzpvFqzV/
5xOym1bDmGZejjYQDUqpeUAgVM5kMUaKZ0TRDySs9A3q4ZCYpw67lEqyspBAQy0E5pQKU9fic9fT
N3XnfS7tZG8HQ4VpsGUhSkuO2eYnc4lAXhtzPRtDU+Uz68b94c9RuU5q+D/Y8sdN565wOPV9EAuQ
3tTNawg7A6Z4r6m+WDIV2xnalKtHQdHXOBo4pHb/lTb1k7Egy7CalyVQ9UYKCqLSew7Foye9LAnj
i4ZHnoJARKLZ0LXxDe3Hu3oQigNX92WRMC6qqsgUkYJFa0x9NT6vjJAMpxbsPkxRnzqVdtK7eafu
5lU4KALhXi80WZPZ3QzG+Rp0thnuA2ASzlD4Qy6DLvVJ9MP0FIZ5RC0cp2mjiJGyDSxuZ5l8JfdJ
pakRUxwPKZaH0TUbY4u+H4RzVbU7pskfGo4zXWVVbn8XAusxZmTfAUnIAzz1Czpx2B4hZsFvKxga
Ifbm13/peLNmzN2uqR6DQTqLIRRT121JiIq/1OQ16EzfPwq4XZa2JTk+OPZw5qujZqFfdeLjNZIE
0TQlJQ4BeG7E/dPdJeVr0RWtHj5iXVT1aReQwEmBGVNlCNNypASn+HgVDIsR5l4XEo50WUPFx0g3
lm7KRqOFcT2wHbNB4OLbWel9conYkjUZ9VN1P0FfWUV1EyqNvn8BFSuRrNRfS8EP+yHSsNAKmT17
W0e8/SdNa7S3maUlrteotm6qlAov3eNpL7cKb2hba839shwwhFv+bVayowka/2jhMfFd13b7cNo9
hG+sHV/rhItdS3sRXp4+EDwPW+5D5NXQJHaS2j/tSE/mTHc4+Knuu5aKWIAyeP+NUzm/pWVVODCt
2j1AxNdpUV+IWcO6pRG8WDGApIQFsR+6VtcpXylvP2xfsMcmcNvTyEedjEpkVbwq1RMRfc0Nsumn
QbnNFw92+jK6hTIxQBwHBQ08qwJwrzc3IHn7pUzxhjTo1oMz5nO8rUYS70niyOR+fU4OyoNuVvcd
QH8Q66I2v551Wnf3Xiem3d4u8CoHtsXDtEz1eODSaYPJa+w2guGEnX48tBvBTT7NUWH+qwZ2mLHH
aN8wIhrqMGhWpkXkERQbTrYtNThyhOoP+Na4An3h5iGuRLVGVywUT2L01HwJYjUKUq+LVyiu47tr
H+mH81Sdk2Tg6OfGIGuVapHjqTYIa2EKznPH5KAOGTTgSlYtLT7kvvH1i8otOKNzU9aBAzIY++3P
pfuE1AN6FHrnjSVP7h2vA4cqs+SdmTnC5pfbsauxo9hJuCdhEFsze72N6WUKndXmeb8axVkOeWgu
8nUSQotYN2kstwRuSaUsiRRVWHLoFpz8lvHfCSgygRiPao2GVUHzVrJEu55/hWgYWxtsRk01tM/h
dk7COjHth3gsdXd7Eu7/qljaTMpyR78xltI+r2LgYPtktOus28GFgx2NZqtnnnrVmf4bp03W1p4A
A46PPtv9FCVUgLFToY6P7wM+RTmkduATVgVTLe88KTPA0HE0EJI6scTXOGTn6dhKeGMO4Wv7d4zr
+Rhop131OgCOgrjypGVxRPTTzWGRrx4IMFoMsKxdgEKm0/9GUAOuvaG0bWDKppN2K7d4isOzdCjK
hzZtZwSz2b0KZijKnAZmL+Dj7R7ULp8w/N5phZNdbCdpWFWQirauQLQIvLHoJ+Cyt5cgPmkaP6fX
yfWnaraNfS2eC54CnE4uUqoG1QCBIxWbAkIVvJiBObtWJzbtZEpDZsMIzMVhmF51TVgbjIVEaKJL
0+FHtGD6/r1fhDPnEelKcJjHNTN680TxACfuqt7IMYOPcVXtn7rR2mRysGI7llKvhmD1nyP9CWH+
05tRLDss0gQk3N6zNhvzQNQ1e9eRxda3Yun4YadNcZCGof7bNX+P9awk3eggFzxYep+13xmH/Obm
gc9GqFy9C8eyate2poCfnH1XzsU7gmWTr2Osxh35yeZ7EGLKZdtGrkANbhm1hMvuOD1B5sL+qE5e
fivH6luTFlOVc1qMvPNFS+aAKOIEgRz3SB4z6sQvwx/+5uZzzGQzy+e+Brm6hvs9LgMjnZ1Tj5zk
Pr/8+906RgGt9Q7K9ccCVYKfJ5VI8J/BPneBl1RSH2mAAW0azypc04FkfYRrZocvOxg3ZPb4poqO
sd5BBXaCS48duLxarhr00m/LUsqCQco4plJay3yMAhYnIA==
`pragma protect end_protected
