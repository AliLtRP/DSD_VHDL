// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:45 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZHPL3DYxDo/ZQltE1oWL+Ph0Fcde4pvCiBl3u1/Oey6gNY5hCdrMFidtTn3pYCiq
wFIs/GeTImvLIuRSW0t9TaL7CirKTU0TyScHGN1uaWAWIz8/FdkXjUkBlGW4sFhu
6W/ZgMRDBgtplbx8Mz/XUvAupxscZ9IHoz8NGkazwt4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6096)
xZju9iLcHzhWUaOxwL75iYIgD+FsulSP6T9cS1nQIXDN8AztLEJXBo/azxoY+40q
abdrYu/DudjxDxQDA83roGluARv5m/NbtAs8PPhJYqdYfEl9AUYU1QcotAxwMsf1
ABIL32ku5zYnYI5GsuXknu3GPjXJah0VIfoNYqG/Pv803z4QbvyziNh6uH9ClgPk
tSlHR3BukdR6z1cfieXCqZoUEGTmQ1kxN6hwzT3qPTswwRQNvGXagSd2xA+LLXwT
lqttfHtOyeNkQvrvRabvWtVXo6wX9yllE32LaGJWW8SxzCr/14vBRIpYZb5ferF/
e/4Qvyz19b8k6BbjAyZmPigEkJIkQ/lBxRbH+IVrvA/v18ygjfM/ylJvRzUn+Gop
LzuXZi91eSfF+UMYgrPr7J+cj/rpe/suXjgU35KMFglFPQvibCirEKYCA5jS53w4
ezOSLZjR88q6SwwpLkzZJ098XEcP6HoiR0191ykt9ByxaBZYHFkC18lyGjCmS7Hs
QbWQFsE6AtXU6BBjiQL0Tiw+0/ajtvft+A57olembxjA+vgzT5lYlsxmdL5qnHod
ZhJycA3NM6IKyyWblXgYJ+cw/vUBj4SyzJsQ2qkO2guE6KxD+dnr7vJ7O2wIXeB7
A3CjTWunDj2c1T/4VNgrn4iAuWPJ5DJX5O2IDzZOGbsxwN3q3UKwVVHY/qwpWyfV
KDEHVG1hn3On6y4UE8mBTbIFhCIFrBYY/g210p5MTmiySosIQl3TxID+J6896UGN
Y8ELZdtvu5YtRlFc76lWrh3Y5QBtUEwAjB3o73D2X/blbmX5ambxNGlqsz8bG7mt
+0+1iMjZV47foF7x5RB/dTtPMPVtuBjJd9cuT3Acb0A6lrTnGpBpnJKd+VcAUj55
KjKw8bvd4h+4oLrBq756J5vLc6j9FWl9SddQ1CcY9xQ7+F3Wp9SiakyfTJtvMe1l
nFS9yq4MLyQTv9jQE4yPWY/RMriI9AbpCB+OUSBnzzQ7DE73541J8Yv2fVw9vNN1
ZrezYAJ0OAjkaz4gpx4zNQyf1Sm1cHs92bn+DSuwla54rCOaNJJP4VToYmI0VQ8M
lXE9aWcvgahBzuEz1frBDoXh70+iK/zx9dmm7j91Mb3snXYY6DP7rbI/tIq3b17G
XAiSK0VaZ+O2BjkLicNJOhbMOgxIhQPtV9gZgjXXahd4AteZtTocSqTsry7FAHXp
w/KoQQZYI5/4058LNLIub78LNXUU2jZtirC5B6ugy9zcDbg70E8Sew8z66hi3ctl
dZVaHkgGupsD1SK6ypJ3f7Y/eH5O3IKdC6PEHZFSA4rA/KdUYzg1r/sKVY+b2YpH
EL4nDQKeHCNYoC00UL+0RNIgmtAqiA8le1eBmoo7Xa57dM0yZup80uYfaQFZ7g73
3zQXUb1/nBFrUAumyfR6k6UUyfmERrgS39GcZeuV8OY2STknvE16W0gplP9qa1jz
NYa6oA3C8iuTnqwU/HFNQr+emIEpR36p2YXRvP6ScbCfAO+LlXfphG/kjb5X87Ms
s9xudK4Ezff9j6Sqt3LZdSQ3bnuSj6d6Kvlwo+2zdebIoHKaZSRnLWVno3YDNW30
wEY0/hiUaLuL0CnU8YNWWjJLsEpofdNtufgkB5uC10u7USjdi9pS/jhPGdVScQ53
HtTOqsLawiF9sTOLR/y/04lh9BPp8yyqr+eNUZqTZ/hn3o8lzPY5LfE9jltRoEU8
DIm71/XgYlaCtIF7untLhJlrUSZVgr+NJ+lNnGLJbI7V7DBl0MKRowzo4gc1Ha+1
EkMssHSQ+kT5oGIhvEc/7JLkjfV51iozEms+zhlcr4pf4VXeqGgKsOWOaUW+TLHN
LiAnGAL+xYm7xxpvwE30q3EIxAbDlY6uMg4CtQe5gyGJKHA07BKsxQlnUO0V9ECf
wimmcRAWhclGguFwRffzghF8aEikFHB5mOwcI0ICt99AzFfe6kbIcdRLneQVAX6n
1cnT30+IT8CiGzOEqUkRwgelrvG9lKWoCe4MNLRbGyVfY12d6igDeQTVjTkwgcJK
GqdhZC+ozaNZbec6q5h6vXV6cB3rHX3m0nEw6IKUs2Z7k1mmBxbOU4dWFGcd7Y86
PxXi+o0mmdObQYVWYw8t5jVQlm5Y2FkbRRHHEt/RWUEm3JqP1EKRFl6GWwZSFlTf
hGvwXzHPtmESeuT8ZeEqjlTycaEHpZgLAhC/UF/O07PgHd245Fu3sfTAxEeDA8iB
7iosHm91KqpYmF7wQPTMVEUeWjSsUh0vmz2qqBKoajntP7lXn8oGEOgXL3U8wbn2
Z5x+LgVw7BM1q2Nr424cwbNzhDkJgY4Sl+/C1AEHHScITYp+qN611LmNJSq1WgrO
9iP+M6nyMj7KUCnJvkNOZmFBZpfIJ1Bk2DXcCRSd24DX2cUvkh0a/i7qSdcff/PX
lpJUvCRcWGhHVuK/bOrdCDXPoR36W2tkuhoVGpGG9uO1AUuOdeRZE5CELxcN5v6f
Kk0baTf8xOFf8f4VWPj57KIekOvnj3cDDAwJfr63DK174bRLvSpbtAfT+CIEfuU9
4qDlL+yGFDJXhAzDqShFyP8JQWnSDM4Hsq2DtyZIXQtzfyOFYq5Sgy2lN/Tts/Xf
wilubZ25Y5j8SMuIP967T/QlsKZCjH/6s2oKpqww3NS5Gx9wlcehfErAKg4W3d95
M6YitH1APOR43hB4pQbzDvuLTCDAgEqKZHI1Qpjc5ATdGLS8O1sHqJ5Oh2pn44UZ
A9RIuVt/OH5XPYj1SrGEajw+c2xV+6/UmNwUnx9EC0WYgqDGsNLXaZ6BFZkYRWXo
bGX9Z2KwP3u0D4uNuc6nR0Wa8wxB+m2yspyhboRHckbQLAxtbIErnYNvLL3bby4c
/0OAyRefW6hCRuADoNE4ajN62JGipPZt7l6rYz43Ac86rMyNwbJy6hTMK60ROaLl
01GtKXBGGKgOqC2tHhPm7qz+H5xdJ3m7qMHxqnApnUrpJ1cBLxFdZPt67iJiPsO0
EllIgqj9QmJiAX+fVqd7npGpAxw/EeC0QQ+lXC2cJKAzH6Rqt48e+iLiWueDJKZW
ogD4FgBWz6se1x+H4v0LKoJRlhhxX9/qx+7cl9RTq2NCgmDgtbjnvPm5XbV8xiUw
EluCZCPROWV+rRiM3ijWOx3kKc8kbLCwD2Ygn33tS9Y43QDtgKvTljyv13fTJaki
PM+QsoN82s1sB+VvuFLVhvyfrRTSz9vC1zrlKS3vgGc3nLF+eLX7ODyVSa/xumDv
K0iCFNjwPPr8zPsGga2lzuLlQVFUzjKV/Q1nVcZ0HnIJuh3e1d4r6T0m3n2htwMU
wYgW+bMV1YOlXEqwnmXiEFs16knnnSfIt4uxfMHuIuw+AQntDyC4OeIkkW3dT4V8
EdrwgGKZBI4JJg9ogouSZonFWPo60GTK7y1f9JAYHdHrT3qGZXi0ETb4SbfoNHC4
7nhr5n7XKIAbbYTToCd0smVpfbpRU/2rE+ZhzDAz+4nOQ/PyxDy2ffPqh31jDWxs
euCJzpyo2yAiSYqmwTDdKsx2BQFac9P3W+KtKN16B+EpRVVwesXC9gDTKU9Jx5W7
GMVq09gQjpJXdvH7vPBimY5mZOU7GYYMJzuUvQvMyZAbix8+QivgzQWIUR3sDl+D
dGILlXrcW5hii11CnFH1noEGLf5gcxe7rCL8IxZu/2r8NhB8ZJ4HYJS3tMSpky3I
anph3DLyWn5LLBxhtT9Fie40qH8ricuG+EgndtGdQDW+DJ6P0OD8358PPA2LJC1A
8ZZ1e/1OS5yD+eCwlcqQ8kC720xfQLgsq/+FkxKzuX7Q5WNDhQTtYUVT+mKQfxKJ
Q290whfHCvQO1Sq6Pf4nhXFCDjrHBs5HcW+L4Z/O9Si0ru0no0xwfu1SSSUNmrbX
Somg494xscY3ymdP6ZDMza2pokvXdGV35N5QKGN78LurTq5XooYmRMYZ15hixZs2
4ipS4Por1v68zXeOt1R4m/hM/yfsl3EzlepMC1tdDxUGxyUBd65ybBYHvD6J/5TU
9T7/CuCCuHa/vX+Pc1jAeiDkcoN1azr9XehuJFwGXkRqG6pUb9izfaTGm8XLS5bs
tdenMyrnkojAg/GGV3JcxmPhjsg5krjsFuLzrMv0B44K/Mb3F05rqhOZSAMzuai7
kwa2H76Q+RzLZm7psY/FIPbQnXMSp/TtHNUEL6LFs7fY9zczsh4jWN4vAv2u5z3b
25UmUSOJ8/TvjB79Q5H9rIJtcOAR73XDvEP8g5Qj0peoOia1/JTWCpRV6gITUIiQ
G5/yvk1q+PYLxGZqDTDrO2Pt6572n5RcE25aeAJzTi9P2zbG08i3wM2YKk1hJLdm
BcuKTcOKnNU/k9Gpu2dSxnQmQftq0LwsBo4HdpugX4Ic8anifq8rWtbhy5CKf5My
+idYivilMxab5NJEsKg3GA0AiqEKK/4OdDqX9sZnTW7cKzLOXJL4BA9qh/3FFhV/
ZQoJJ6Oi6XUZqZxjtNxBo7WQbfmhI0S+eMqUysnK0tYO8CqMfM3imF708DXX78uz
7HkCP64wS3bPjEe6CKCCY2UdJgJp6hjzM50q5hQrxVLgPIw0yV9aVPdmE2dlq0VP
0HdBxf4amZdDfYMs9GL4vTvuCcovgtGV0SLT5+iQLXlz2CKPMi8Sbrb9T9qDYujB
B0P3U8KbUxf8Skz/SVBLaVJSW2QZ+PbLXYF27hUNDfDKrMgKm8VsN6quC4eO21/t
35baE6xlMTGAzKCYNqyuFlfZ58O2Hyh/JushyzWw2x55TBN/K5kYt6pfzhrHilF+
weTVEnNI74ATp7/vIxkodhRC9oPV5tsP0bQ7DcTh/0ENfdINvB/o4G7WeNcWbW05
9+LQYGkFTD8pH52jSxhYGgsTOgnZyWiw5Zq094Lh3f1+wvxjACy9KOqc5WDLYeZr
e3teqY9NU+Pa3vS8jN+/60nzSV8ny/I3YyRZPre/Ru9qkzLSmWQJ+5myPaB0TKRR
U+3BOj8E1z5vU4D22RXFpVeO9WQZbYNFaISPpI93nHNJmOdhErgSnSqfi/iuNTz3
Pr4g9f7aW5j6yrgip1fNsDSof4ezW4s0bMjwBJGClWMKvsc0zVB/vqx5wLhy2b4/
uusCNeUcIeuJDNLIuwqkQObIA5F5pDdzwKrBGu42KhjG7TeblTUTt+yX2GWxBjqU
d/2Rya3XY9lc5srpkHKWhRCL7mNJ38wqXnarcZeHLCTRNqaEB/Ci6fzxx1Jr1UKC
qcDfcWYH/7/bWJ/GtLRonOzwm+5tDANab2v6G+z6wky7geMumxW0l0TuNoagt/WJ
I7DLBXLlkX+QdKcz7KFK4QGWAE47ZiuADdTxtCVRvYeed5RCEq0JqBd/X3mujLww
mJVA7A+IvfNBiaZWcqpTUiG+UqTJzDp38bOEHqsGjnQOkXSh9vnYz7mUa6ddW4cu
htS4yf8ERcSXCUfE06fo1xZFl9XHcsv73ZtDxzgUsu3WZ0nkmuyuBrKLnOl82Kjt
wz2sVGfnOXnoDkMjOpoNZGvgeYF0CT7BxBHpD062zG5f30Lo2Hsm+0aQp0w9/oeo
LgMOP2ZAMg65bCtDFQrbD8KKhL4mI2pw6rylHKze7o7/e5KOpF2pwfFCfcKbCDSE
Rz8YX7cc8uynq4qqtNPy6Sp0wF/v6rknZ4g9rUgbuDdUXtYQxm6C+IEHQ+EWNvTV
+6ZQZAGEJdccxU2gpkyOqdeL6cHSFl8nFhFGV+kNjebRGsJpn+cY7N1K5v3Gutjq
5QSbXnbw6UNiA0sh4VcOktfjzvyd1KdZ0wf9EHJZIPGFnqOUgxafUaZRtSXL6uJS
+FlATcbdGJ+gnv7GKEoEx+usOy+BsX43fiM/mZUT7HcJ6l34npPJaa68NgChFN9V
2R6NB4otMX81Kp6Q+DnSzYa7ijalvy+Ut2bsCjmS5LzBOgEBhC3m8nzP7Aj1zO9h
fr4pDMiZvwOxk80fA47zU23vfAwejez7hD6s+CesxhfBxbMArpqbJOKce2cvKFq9
BW+yHitI/YSue1jLeOjtjpaEwJCxjeo0jafPDtdQG8xJkcS4hMe1c3oubgw9eTm8
VHRp/2LwzdOlH0nE7IkRXMUqvkbNWk1HEiDG6aDytiIEJ0EXoX3+5shwmZQDuQWB
B9PwUddazxkq0bBZ/5YJzLbljcj0sa7AVlG7RwYJvEXSJCqncToj+Gf4FMIUhEBN
H/7/rMhSEs53TdSdTT7Wyhhv7w+o+ivqqqXEI7jL3cCOiVumIA+hkJbQuBWnvgg7
pXY59flmRkiVy2daML3NgnIkG+MEhpndArBHRQbDBxrheZ2Z3mKXl+CN4nRgVh71
4pWC3AkIaD51+2fpo2cS4g1/kZWBYDMOmCH8FBbQ9h1yXiCJleAjqzwNyrcKTf5W
G79OpbKfiewWyIEwJ0F9jukRlOYOMV4u9fCqn/MkgCYJ9daiLNhgiAHln7Ce0fvf
RIH7W5LDicoeYmLclLflWeZZVemqygef9F2ZF+jAXslShTKWLJqEUtQnljizrPH8
CIt5fGCSYFejGmqYL8Fo4MkJeRxkpc1hJNxlf+uWf9mztYnfPmYKX5ZM5sOkUIei
x13f6H/VqmYEqlCYo/fpeHqIQ8KyXT0mEw4WbykaOIgm0viEpbiNNtMBGoXLo4g0
8EjZOrH5338fQhdzeru0BCpmlb3zrmzBmYLsO6uZqdQRstZcOlT8YRAygDrqjoK8
zGxT6YZSzm1UVu1VSvzg77JTan9XkwRgl3/pB8G5F+35qqZf483zUvlKRUMJvLBE
AHPIJmaduISr/TYqZ3DcgLkDFhlc+XA33rrJltcaNIy571iogpVxOylNS5AhhrOn
ArgKBJrI47R1FlGBg9Qg5OrwBDbIWq03XEJoF50nzFdmt7REWjLhZ9QV6PuetgHX
CPThB5dP2ZNOwmgkMBkYGM2UYqdj93ZwA5JXJM5UJRd59BxmjuSpjXbVCtR+jzry
x98K0WNtDeVB1z3aVs+qBZGCHC1U2aWnUUu73jT/V7xG5oZxeJFapH2hnkIq9OKI
4Bjsqw8g3pHjeLbZdoEXwpHaXeRuAWAdIJRqtdZrn8wwa+B/KcKIVY+5UMmsB7ZH
Nt2nFcSZ94TCLQ3pmmRSnFLX6j5xY2rYkx2Z9i+T8jKrweFld5v4qIYEQai9NxEJ
aQU0Uqi45EcpZ+j/SiRYC3JdtLP/FXrjmzxHQuRyc9K4WA+IalkSU2f5nzH2XbLH
O/cmJQTnO5d/oyLtER+DuBdtSOG35WWmkBqtt+e7LvILLC8jcS/kqwssoZCaLbmj
OLrU935ZkxIDpxGKDIdTnMMvDfPemznfAFtaEBn/dPeV1//nonRqDzHX76+0J1bB
wCEpPkFXCi1is/OD1sKBv+WCa+wa7u7TkBZIXQ9dCPYFXgokGGTyxUukgwdHq2Ib
crN0DtSSwkhcmEEdUHT8CUftigkiGHIdhwY2O/lXoX6sqqgwxjDC5BfdYRkmGp2r
rf/gQUAQ/84YX3BuSpjWKN01ZwrBAFn0/IBUUexchmAtmWp8KAPNmZqUyMd6OIXF
x4GhNGFBeTs0vMP0V+EfSZo+w3wxez6QRUNRofdewne27ZS3J8FOAejJSYDFWbRK
KV9h7QBn/AkGQQ8hJka5yjQB1bwvgOGVgAQDn3BiOkeJr8QFHDORkJrseNFuVoiO
ihDM6IxrYTCBS62taCAWTB2b3kXYlKgNsL9fyBT3v9J0xBHoZKPV7UArppoBhYwU
xVAb4Rh0in9cqtirRSyBrMydpq+n4tYMSdr0ZalGJGRpLos3fLmRTAO8smEv8mmn
y153ah8R/RWoUzvR93mpqHF3uIViGdFNNQnRDFhDPqXAGF3iBYMnjxz1L8+9IzRq
ixhsk8V+79oadyLAKxn/tC0tCBbKSYqRR/dNyCEVLQUEyRi7JLfVTSuuuOFTbTlr
RIV7pasaRanLkyXLgimfB3Uxl/F/iGq7+O2pA76mkwkRVqYMQnlcyF8ZleFtIp4x
0DuN5QSHxk97dYcADxyeAkBYqlSALn+SvISpQQAItNLWTpZRArpuAxTH3U5JUGW5
PAitBHTQDX7Iqd3mvL6wql5CRu2MfZ+OD1cIZHkuRoVrWvb1DNwI3dbahL6Uj8xG
`pragma protect end_protected
