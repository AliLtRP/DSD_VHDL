// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
CMHF1TSPXPBkCzNe+Ba2U5KbRCFF1+BC3PYd9GiXCTV8Senix3ar+qlKC+blBcYb/Hc+8QrmQWxE
m16Sa5VoOJD8bNhL0nQhvkSKJfP3R5S73u8tcE5KwSDDCLz2LdCXrLzGqk1uJsZmvQRrhMol3BKu
dRB2K3+nPfA6EMj1BJQ1Krn+eccVwyor0l40+NkpDtTOdF5XduiYz5YDyIpaU9FJLFiYlEGE6IBT
CW7DGdC45nmf8LxtNhpowjgObE5WyZC5x7mW676o4EoOzQW27c4fibCwP1WA+bvfgS/Wg5RI6qLT
izVFKJVIZFAI7zJsdBP1dJit/9GAQYjg8CRr5g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
C43nrJbf+RsOdGac18yg/iaIYu/yKkNPFy1b6a25i5ZyVaI+EOLpR5JQISaThcI+jzR6av8cazo7
8OstqtTCX7T/8P0LjKtr+H5epuI6JmBrGcte0AjXd/kwZ0wW82mJM/cTkhSHhYqLrytHhA/p5+Z5
Hbo/Tne8iCtn5qH1v88ZNuAPQZlXOaQvg/K9zgLq6qLeJHN2iFohmXbsfsyNKn2+gbebr17sEnzS
n7pqdVp1Zc01i+095yLFvsi0G+C8NiezU8sZJ3J9KOCcZWl8YiTNphaHFrHJjXKWWd+BzWlG/tjG
jRlV6/YJCk7CdS8BU05Tpe9mt+AQfe1E31EPWEhs/qKfmlMfHHdNe62A2aikKQ3rTUkHXg3YFBBa
jMqlbh5QbNPBWNjGjWfpONQczFQIaqQsY0wA++/WP1dhL8fO8tL/1uBylPOfUVy1Un0W2tlTHnRM
Rf7CUw6PXq5R/ns/q3NkvW32UWL9OVdtHJBQvW9AbIyZ9Zkpw4yXNVan48en58XEbE20PD2TkDpF
HM5KkdBC9hA1HdUA+uI9ruuMIszzAjO0Wy5NX4gmIlJ8ddsiI2GqBpCknWFZFw0aRIHD+swGneaA
JaJzQQSGfsk1HXEkdsC4cQp+TiGKeVLCRVMc9abOxUa6POBdNqhrxFePD+8+jSlMbr6IpF8rhAXq
D0zNFUhGTPX4rtQF9Ph0IVHhLmSMvaUuE63ZbDTNwfHzljC0ectC+bfjxYXhNANE0Dm/wIXTbI0E
yNd7l/jFpNiXmtO8YHPD8IAnM/Q2Y96z34RisZ5Box1CQNEDjhAfdYxWCN3i9ThbkkEwcar+kCZF
vTR56fW+av6oOi+Ra87jeANXffQCPTGDnFRFuXIxYDDMWOdPehMpZEuZc8jH/sm31qH4ftrFonON
xp/bJlV/3z0/yQBGjj7I9KC2mXFRcA24k+bNM8sjWzBUB/5JCWTvhA1+bVyFA+5/VorBgmIRnWXR
pAKr2fkxdhHv8fcqcm65Zl4jNnBc51e26mcHSIXNXHYztG7zQgxDwsin0i5FBovFwSpi6XX2sStJ
h6KVnrJd9DTbGb6M+SwfIpSEAlhbl/0u70jHI4bDLC0xEdd/3mWUZhWE7rrsgVMVDEfn5OIDjeTw
dUWAg6RP/9QPPVJdlW/QSkLK680800QO8pljkPRourSqichmUXbSCJgJZ8H86F02bDag8BHs9Kep
ur8ALSbrxsRj/xAeCHFV040UPqUUZ5zzzTbLgcAsopMB9gMunA6PfMZevR/2CKsYJw1bOd6lrOkm
A1vyXQziwn3hwtobCybNfblXH9hhWLrsqP4GP1k4SAAyl+9crY029/Htfm2koOI1R4mLzkpxW3id
h+yK66PvLUpObO2QdxIdNDCBcXLBulxkSGNeCPdKudNNNrEmoTNoTcEijQKpl1W1jBEprnRtR6Zk
0LwEfnHm3oTOuOUBl3xPwcoYZ5L4IjhHgnCPCFl5m8fFaPxVxeEQSruzQ8AH1z+VffC0Tjq5qgQj
2lHY6UnwTKSnxp8SLp1acPgo10YEEY2Pwks/VJ40Be+Vh1cU4QholMsAH3eAQ5M+gMoE4Mcc2oUz
lNMs8rQa6tZsamFiIJKPEQv9p+RTzPdCG1Xb3AIVDCybNAgKWhDeiI6C7YPvqQjhsilKYqdJw4rZ
T3vzxUUoZoLyfnrmV16QBWUnuyRTuQ8PCNzHDU2owSIBzjVMNjruzoMPiUJ/FqhIVgCQeTT5238C
iS0UXVhbQdkKDsTp8t4lGEJjLSOMlEl6SMYGanCUYMeet4G0Lv466B//E+uN/GIwXSSuNabj7zvj
j5IybWshhaknPmUhlfRIiFV0MKowPyZytvt5OVykTRDlmoWwo+2TgASVqogmalyhwsDdW1AMZvdT
PZ65HWXl0XO6hJgFdeu6ZeVgUI36ktSgVS4hzyIBuPzi1OkagqvjR+DfNRswefvR0F/mqdM0jKfK
svKHhcMMikov6393jpM7ATuKjjDV2Rkj1QN5sqfS+eXwqLiQpD0mREaRxR9DiDSh9MkIVeuA7B91
Fb2OagMWjXS3qT/yc1pQQuHYYY1bBDfyNKPuJImtLTSHiVwO0mLwYubHCXGaJcxVV9N+UsMPIT+X
BQzQUiDTcKDqfmphSP9buoCy82ZyiR22C1z8y0LMVeZdhAnfc2VLUPLa8QkfrDoVmrZbAqyFoxn6
l/429mxrbDum1IsguSjuxgp3ZbVLb7HbuNGfxPix3M7eWsdn4IfWgU387o5tYTjS+dTrTDs9KHPa
wc1F8TmemvXvnj6S4rN82BfmvNomR0FhmJKeCEHoEH8lKe3JJrO9YIXbrwbwxtD8XdGtr1W5nSv6
tf0b1nP5Ui8EE3omwy2YToOarLuy1Wwupl8Eoy3OhuXWVSK9SCcN4NMsScW/75+rMeicmbe+lOrS
iTI4+IAdyZortxZg1kiUAdcJPfklmsd/EPj4SfuyMHyE9hZFo6Exal3CX8CdXTgzLYrqgdde3rCv
OqbP1MvnBm4okKw+Eupg/LOZFTjwmuF4Pe0uXVERiyO5VzGvBdBmeDu2VTNchzuO1TwfJmbD6g1S
VcbkyRIl61DDcf2bFC9uZWeang/zzeo9PVzOCwOLIohnlmzX0UYXJTDyI7Xynd7CSfBnUKAv5i3e
GsJBlMwepSVPtp8mWJcM+VKwULz5/hWtlTyACEdotliYchhBTl8fqlmgHUcdd8IWtn8eZM7RrOPx
vmpYCPd2eaZKyTbfOfjL7t5S7QXCxc83mabFXNxrj3POXwYVw8mreZUMe0K/TfM8fsAWR/DQZnGA
W3jqGkrTRmq0oQPnr61Yz2cilqtyRLlKQ9VttBbbBElFa0Y1x8e2FNIOlMRuZAqAGe7WEZ3fmtHs
bP9RQAF6I6cvrKcPhvnBziVxq6m+/w18s0iL5rxiYCKu8QUI1Sv81cdmWcCHm6Nm25QCyEUvVUqj
AraD30etELQgbfIfD9kKOxcaxRZZgjM8T377W9BcIocAIl7vXHvECwQmbCLSoOYFCBRFJ6nduOzQ
MNjqfXSx4wG2Kp2AVDm/Dsu1D3kXb7T4fIRqNLuS+xxPO1SJd/EUvEHxJEjBqUm33kP6kckQGJxn
A6ZgRwGsW3n10IEB5CM0BQOwKAHJsuwkF1zvaRrhf90UlHDM5NH4ZWozGbam9HEpF3V4lnbJdXUS
yYRn33u3ldFPDJEpl7fZbWGwb+h5LOo4ZJsQsBQm3JHB13FySQpBJlxgBLjmicBPahi+csgbhZnq
9FoLFXe0I6vsuDzrAnuy92qnolC4+lwdx4wzxdatxtAp3ledbjA1U6BfRPymr+NWVJVAEn1jqWYG
ZxgjrqcNCo6eBh1+G/bCRTC415yBp968JAjHLyWKeVkUaJoG0ELyGspBXoGR5oVchH+eMoLic7Mj
SEuN7J530lZPGAW5ICN7qXANYtsRLuhQFrnL21hEIW8hUUfwB3vH7uPOCM/2+geEENDNJx+8/0il
kUfvAFKsA9XKPwp265OlrTp1UdlDUD59j9rFC9Mbol47FSC2fMIkyGkgNG2lHuSkDnlu14DW6gJV
YM8ws7/9hj7wUY7gdnNAbpkzpZPmafa+xUzukXXlSrnEwG49FRUcEy05hE3mYhdX8xzLxis3nhkR
yGRa9nzstvIOc8qbJ99gxTixwmgFy67Aqk5qX8sK7LIp4InKQoZkgoU3Ku71AiH6sIrK/qVTjIx4
IkeraA1ci9xo7P6WZZ6cAiWLUE6Pu5ceaUhs73HhEfQNEwB05nQ2irOWoCXhtLMvTh1Np3N9RF1l
Im852IuHmi/+8Od0i0Rd3oEY3onbjyp68weFVsf+55cnK0ZPbtiJQDRRvrLEfSJ1gBZ4OwsI2DDl
NFzvCpXHkiLJpXCKUu+Mz0CQf4kLXBhLIZ7HEr+MyKhoEM+o+v/HB4Rke/n+GUUnnZy/JNjAhSaa
1Ye4wC6WZ9h4gdYPpelmIsOPE2rINvTo7ham/x9nP/360etekfbvq9RMC1BKIaDiVkN8iQEJMsae
YgfkOlTDJyRLJF8oorRmEhK7TaSoNdvzt1KXOyR5zDsYQmQZ6hfiLpS38FBt2if05QOjoB4EDg44
9H4bsBF3CX4ZEWNhnciTY9ikFmtZDXGEGBT5yh+O7elO46OHOAQo8TWDXFEzsVuBPE89Riv/3KTa
5PL1dfGnTm4DxRIwf1v/h73iGh/2GTzFJlBLVGAyyr6BpAIdfHn6VqEOvU0U+APM3wOrALMbodvf
NZjQqM2Kuel4QT3fIweHz+Vs8/PABkJRe4/Y05wIjF5Uqae5f5zkpSsDvgrApAYwO8JybBd44qux
GLf9g4vqOUTIBOt+PAvC7L5wNsOfD9UGdMV7/e0SOccn/kySQzFAd3AVOT9LQVgLq7M88Wp2e0gX
JDejskhvbiVbSnqV8gjgy/aVtZnuU6fytHxpi8LMMH8tJVy2mAWtDT1E1qXucM/RKN9SjpYA7hFv
EAuUnbHumtjmGskp9ssq7KKUzNmmkT8wTbkvFwrkxMUJWWbogYpmA6Iwf2fDuDQb4lHAnpYH8lLM
DcY6jHaJGW8yAcD0gE183KYuesZ/0Z35Grc6XogKk+8XwEdwLKQQjChtEAEed4aK8cwQnEnhHHAt
qAFFGhoLWLtB2S98kuUUrsNXLAMxWL13FlsxYAhRNnvT2i7TUHgJNWBPjFcpsb+MSchoc6BLD2h9
G7LFEkSiiHJQG7N/wVJoDOTTy27q2cDh8kdv8Xcti1qozgwYMkK4FbJnyKuLigiG10EnEOd93iEn
1ACKpeRS76l72RJp8W5KFjXzQsaqMltPUPKiLSZhS+2ql/PxATqmO2EgQSwuhUk+661TVTIxWv/B
pTIuLdgGnQwJD0c/WreOolu/xykjZSr44S8i4vNxaS/6kC3kynTstq82q1MMBp/SXsSwvZ9B8mnv
jVPCXyrFz/Dfi6932DZWaXTZdWuevbtgxQLlbFO0LLge9jrZS3TgjjWNORrvqXsVbVtHumLmKfDU
ZNF17hnLI+xCz8Tzjped5xcE1zrQXzTyucbGfwLY38Uml1B6JhG7R1vIp5ANGQssQVxMC9SsrNNV
5skGP6MDuODrjFxk134QQ65DhfjW105s5zIwHzhLUpVcteJmFffr0gxMOpqBhNC4lhNZ5h8QQAnf
JZP2RRBuvoYKJcc0DcmUe9Q1sw8eTAuAn1RG0ZqMAKEq3RYJiJ/KDV1AWaCvRY4FBzBq7hF9wJ9A
9t7duwM/mx2Rnhek2g2qLm+iaWG0vPqF51tHFKZHwZKo+QfhfBfhpuS8ys5Sr54RnApHozBRGGlB
A434lOz53/IFqjRmMCmITS/co4dhm1R4YPWrDftx3SMMfrIoInAAJD9xyJXMehdFioh15/Y6L8aE
GcN+AO2LoRtIeqvd/Hglpg2yARJbs31IzlmBZspUIXawzojuq/67dJeNu0tgGl/lJ2yQsjJe7y9d
bW6bnVCM8cpiCTg5O0pTPbejAFDPR9adsKiHWVpJO/VaCDi2+3CJOSkLsx4umNWt9Mxj+BNXOpJY
070LKgURCzl6X/eF7AoIfjVrTi7XNmpBdsxuQIUvpo7FwcFu0LqtMyyYl5Kke1bMmuRkG7Gd9cvc
cp4pnC66gk82+nMZjk0WZMxQRqW9ircll/QNeKm4zlSDr7UvPv9Uv3eYh3dlY7cyXYAkOTKfiRSE
wh2VXGtfjRDfZzinZEbpKHHt0GjruDs41xBO6rVcV4YtpS0kJ564u3spwc8cPpM2qqg08VNVMINK
ZtzbrtmCtpngBRJXr/jhw3IdZdP0Oqq6HrBTje0OPDmWUP8AFJ3ildgcfJuyxjdHwFidiWvZCqaJ
/vlGZFA0Hg2ZvhQ/Fs6LzOdZrDkRv6EUtrvJRQytBoQRLaJ5R6CjuxSetgux4daALywxfqb61W0I
trWpR0d8QlXrW2388WhT4PnLaPEhgquX71ZmK9+xYMU/f+mfnFTGsGi3Lk8UIODDfkDSBT1keFDH
Jv2Uc0VB3u8htoN2qUDUwfPHqjKqvVputAznirTYIyedlKNlusZGtDXnCVCNkjzf7+pfiIdeWbqA
0PT13ftFXQJEmmvpW5ItNujmodRlLPFP9XV1ZVLm/ItGLgdP/DMvVVP9KWNgWsq88clTOmATW+IT
mM2kskGh727696ME9f2I8QnEGglee50QlUvqyZnCHh5Ul6r6GSdE6MtRKTZ8kqPzBlZokDXn346x
QEDF2TfCrvPo5SSoGjDWiqAkxCuh5VTBMafJSYprORFzM1UfSHbwmLCAV0OpORGUteMJsDIcnKy7
Hon3BDF0b1DRTWA+K6y0QGYYrTUeZE9+KmZVrlaf01JVa3As2q1/70eddaQ2LTwQR5pyCL+B4mjp
W+xuJYi2PqA3N2hJKPSkgyi9rB4it41yWL8+f1MjqApzJv/VSSxTobyK+iiXY12+GEpl1swpDBTR
3uinealf9PaBK5Rg6Avtrg96rsv3B/rXxWBTWgOQYIPEsm+UT1FbrTzUklrHPSznHJZCOh+t1iGe
WHZEomtzQPTyqSYh39eW/c5/7LzSjerf4TGoSndAMrvT+6wigq5zC6oBMIlzjZdux6V7bTRj5XIZ
i+cHy2s/Ktc7mbNTa7iVA0p7D8O9sxqgC+l00SqXeGimx8qdEDbGZF+WvNR4fdQ+TDtEZV91x6XK
a7fFgz8i4O4xEHpBfo7OQAEXwmRCpLJtraBavs1j41OTIRoeH9JG3018/duUGWB8jX6Sft56kTPV
MD7JYgYnWv+Ggh3xY1ZQbb2iIiHICNnTqNPHxvYPrtF8J9qME6EN43nuMj9R2pShABPkEAXI6tun
ndG4e8RI4EJr10OlmCIzFqOZviKVoqiAr2TCR9cEqDmeqOYrU45gkvVT167xLGASfYyTDvqqBJ4y
gw+TP8Ff7sT6iaeCQTZr/Z8i9ddqN+xLPxJ2/zy01IAOBhsGKlhTV7JhAl3SxIkQzHHx5yz5cGmG
Z8vm7izmmtRtHmUX0YUP32zs33HnLhqcGnr6dUKsYZbIuVUVl3Ii8lxBs92sJf6yT2JsldVSVNcc
pgBF6vK+Fay45+s/UpHeso8KsfuXtMWJgKwqkaqJUoNlEBMXxBtJwix4m2jvgTHAdCpg3Pkeeb1l
jSuc/yMpAtydinpjGEXE35/vYULPAPYQRHGOxPQgoaYWI0ZXst0h+1+i0XrtyU6t6z5+ubfiwFN9
JIR+y4pz16bp8b85pl/8ike52g+5la4CoFuIKfS9O7xL3LPTeb2KfVmTbzkpWMAhklnUvIOuH/7j
Kof/i1WR1ix1rm4Sf2b6UT6KlWVjysB9exVzbqqHg3LCF6Fusn2il33IhxUnw9A58kqZGTrJ/DGS
B3IUurrt5DFCF+vd+DZDx+SyYPBipZ7wWB/DvHki0xGP/wkhmQeERQsDXZW5Ba889CaHoLIth41b
ZXfbS/X54dKR6Cvix2KC/aM3n7WH1R+nb7vM15zF8EuODipEvZKvu2zEQ8epkoG7w5xzxmLnWl7X
ERFe378FHLcLHru/W5te+Mk7H+/PeqcPOEeuOSSCUKHpBLpTBR+shhwD9K5wpWCkMyz8L+3tfcng
8vzFsYilt0OebKXAXn8Oho8CyNwBGXty7XSHCC0vyFQtJgzR9+ZeV5Dr0mZIpgSb1wEcSl7Gyf/9
H2NZJwtr/N3KrBGjmR15fNKOJvcNLiIHk/vxhv8OB82dZWsfAO/PDfHmdShx+/GzN0FobDa5PDVP
1loNPoI/cZSjx2Y9yb7Cu21mHqxRgO17srqX2kv+VK95u5OZM4fvl33WXJjBwZBJ9YSLhJ03njPP
KxoCTmN2Dh5w31FwG6yci9nAXKhz4qWigDOI1NmiPoq9wS60Ua1Tj465uKyQfgcf+umzfZHP3Rtg
NL4uTH43MyOmpvvqu/uWnz5zMhFDa8qUWYATXSBwnfYCaooa/qec4ag/8aoLzshzIoNwVPsr5o9b
1EpHaoXsAEHC1ExLOiUfYSdOpeJ+Fvq1ns8mn4RDC38InKbp6uEHDc8jQYlrOJJ/trSXTNC6q/fa
ko7Pt5QDmRZnivP5UcsrRrz8IUKWFXGThZs2NL0h2sb93XjjiUnbuK9YOWhboJ6CZdZj/BYfei2o
xRM1v11N7ki2UTATuz/ZNeM/yeSn+y1fekmn50xlnrYAVBwBo6CTfKLOQZIE5PuP+s0lXN9rp2QF
69kiasoav6MuY6CHw9yId4FynM8TNXf0I7eh+TCbAcIfE+/5PVBUBqe+t98AlqCfKseKFqC3sjt+
1N27+plZJ8F+iZi3x9XO+N75FN57soUfOWIUfsKBuKgUzXhqCSqkdq8dYWPkWow7STbmiefI2bcf
R9oSKoEpwJeWP34ZglitHPKjs+bY9KsWZWUr2lWJetQhZ2GcAoIIVSySaHduooRqrMabsY3lRdMt
Cp5rILi7smFMH63ITtCwiLw94P+lArQgZY7RkItuEK18Tnu+BprzQUr37zuZQzVfJ5t3p2qrbXoP
C8tE1WnUt0qQtCmbrBxsvPNDE6aDs6UcmVrK17qKAAsYHdT3HmjtIpkeZwi3KYA86tp0wsodpCLM
B3a7I6MU4ptoS9R3XSm1zLGEEU+WugKHxV+CJROBfVhEm6P60/kC36jM0IUyUFcg1NvG5LrGrp6Q
M7BlxEcd4H/bMA/gxjpRnYUjdZet5D76f4/nQOxs5ZRHi1yjLGhbTH86RFH5yngk2kzWPwvInQm+
ZF4o8F1KTe1FVMg54cBh+/OFE/9Q+PGPUwx0eVc2VxwEpeCRRZotNcz3bk7xfbuMI1x1PEkQYy/9
yXE8sD1dzw0T149NKCTF1zyHW3UHmJi7q4KroMiZMdi/Y4ul/BEHUTdU1ldtCuGg7xKkxNXMrHBa
6pTVP0AUdW30LCsfi4nzoQKC/Bof4fZ0LwMV631CyBUi6s2Qdj07tU27tkEi6d1h5EQE/eiPLobJ
B9hIpd3q/G+hRpMZ6fhEm/hpjY0fMlOuaIES/xk37Rnl1gOjxOymttTcMZnfN5raG2VnlvPWRiOZ
cA95NpwcLSIpH8ONp7WatiI=
`pragma protect end_protected
