// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DWcIy8ps+FWHhxxnl6ncZR6iWuilp5g02MlkYzryeAu3uEr32bzz998QvYEaEQVr
7iEkWKTSSGAYJVQuT2O74K/UjxxUG+jslyUZISkA/ndR8YsxFigC/lWKLidYPG+R
QawdPH+pOyIGx8LT+B/uyXEz9kEHK4fYNLOYcgovpK4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6400)
ZRcMYgp4ZY2q5rUkmh1WkxiJ7rLCvYwRUIYEZZY50NbOOw5UiGjfpeubQDWaXZNi
5AqvFs9dmGweMrWMHXQX/gpMD3u0vdJR3Mc1RVXDn3p5MO/22Ro42W+MxOSXxYvk
IsxGkL2EqTIYJbLNgQsGe360ll5qJR367WKFiTiDHGQAijJymBuvGk1j2HZhzJP6
9WqBOmMJzOyZCC+gk8jB4GitYsuNbgNhmbUmhQetbxe+TnFD0BwKUoC7TnSzyZzQ
OX/E/uJcU2N7yZqIntkNDslPW4zrtQek6gZXTNTI7nNgGnlakOKY5YSyDV8FjB8n
AzYCvYsxYIXdLFnTG4m3HXKb8MJicFXJlFx0iBeiZXsgQNXjQYLxdXQQiX9m6xkm
amv92Z+kGKf0fOh8rAYqoYLFLe3A7DXtINmzR+AAPaEgTwdfMTkyHuzqEzJ8THxu
Iq1lWcx8KTd6CN4HnTmVtZDdCAWBOlQ3mcHTCz8/AxEDoqj0Y/4XwovzmDk7yedR
ofKmpRaQm0mmVlOTKlmDW/5KXtiKLHRbXJi52nUDwSrtr7sI51Aw7QmaPKsOJMrR
LeCxHpr/RXk3lDG78ER+Ne0EtmkP48oTpCc9LzBdTdCXFtP9m22bJIg5mgv/y6fI
8PmNxGeDbtiLtc7HisSNUXFwDdOqVB6Gu36sC5XOgkp/k1Z6EwpFn+Ca7NbPkshe
WWShUo8MiT1NMH3rIXZh6D3qHUIxcTzEVThpE8k+cML9+Am6pYlSQJLqfpJYoKnc
mGn3SpmtaORmq9qT8XCQCqv5KkJ6qaBm6SbkPBMglVc5toDTe+e38ywEj4XtVjyt
XXdXXat6uV78FjrBF3QJVBtRyU+w8Pz18+AjeXNwx/c89zJajWfCwlCpZsWIgR0h
teQVwzO93VPDVSMoyM4R06EswOYiyg1QRYzEzSXg4BDhTDhWQ9CI7AZEEF91Yw9G
aG778iPeUxcScwIggfgt9KAspAHRD8EEAjuVTNgrGr0vD9pfNzH9JrXQowJ1LmAt
UPAHUTFtAeTR8mxa9Xl6vkV0GhAr8NsVbOcup+oG01Xdsu1i6zH6ZnAWlqAwjQ2o
Y6IK6hAG2Hjas/a5CvgaDBtF+6aeYfrqIXv24s10/eJmIXRmmbcj9MSB57nB/Q3f
hHIFaUyF2m34N1BL5EqL350u/Nom2AW6ueDFAgEt4K2PMPquouEs/KYHTS284pVL
Nd8B3tG/zVd7ZFNQE0sJRDgrIYWiqL5RUZnTl3HJ21Jrb9JJnLRAuF+Di93jTWx3
IAIDSQlvcz/aJ9IrmEcicFdzcNf8Ngw1Hp8LTVnDwtMVI59UJSzjXfV4ih1Z8Pvf
s32xHAX2LdcaT50f4rBTRQz05HRBtAJnZkhkFfD9WkoVtDyYtewACJAbsG2Om7yc
916PxYf/RPJ+ZYYp8qt2CQf5UY3tDVPcJ90404nOg1pwrrF+I0xLwcUR1amFSeVL
nOiNjOLb7bN14tVitjWI6DmdYQgQxJ7s1EkFATpsVfe7bTMVJylMtZNFcyczaLkf
0iBM4x0BGE9eCUg/M3WZ2ImHdyTODWB8QCavI0um4wjbOj9524igb1m2i5mpxYOj
bJfnmh8MiPjnSTHayRMUdBypc+MlCI9+2iZv3QHOnF3wOGoSD08vN51wrbeWJTu+
qRYHw3kAxxS8R+tUo++N946USy2h5M7kzSmsgI8yeqOCrOj8yqYFRydWRUq22nvy
d5EGyKDKLDE3Hl3GIhamNhCqS97QSTy+MV2ulnnNcSDUDBEfcAiFLY98rR9k3DGD
SESzv2Sg5xgKVNdvmlRtzMWOxobU9bsz/fV7/jr2y+vaXyOUL3doMoK6mzebACHh
cUup3w+fQ1sall7gwSpbrKsz5Ka37UmHUf9wap5owCtcWVZVb66p/OrDo9Uiw8Fa
pB9Ytu5VgsghL1wn4/AI/Wn2iUBn9xrxoyNh0Qa1lrJ8ZaCf8UJUHqnJt3OhOMUm
JArvMvPu5bgmEtu9mwldfGMUdpA93E8s7Fh3hv8tz1xdikuTbXybddnMaCmNLTdq
VsDhrqvu/haUnddf1afwerC9nIenJyNN/63tEjlRPY8KJTpHDOwdG+5eTZnZSps3
vhmnKTXh76oHinvQPWCqZvfnvTT22ckvORgnEzCEYRjwy8SCglXPeCXrKU+ErwoA
pmh16Cyp8yMmKjMTG1pxXvL2S3DlCyEQszi/ZG3/mo75a9RxfXUwz3hJlD1pw+bh
PYK1+SDoUpBD4RYa6SodWsj7zUU6rXevQzB9cv8R3IwzIZfYZx+88hJmNVTpT+aG
HdSkBcVoRvXhi0Mb8BDaX580fAINSg15FZxKxFs9YxL8RO/HjcpRfndqF1qaKpIj
Ov7OyV9UoAE9j64gBy2TG6i+obf6jwOQ2K/YRQfDfWocvP0ijRMpEvejE5Ezd2GA
fSZc4II2Aj6N7P8L382x1EVDq4t9sFpyVXr/dJao8uMwfyMvP2n+HoOgzDN6w1EL
gqWA8S/F+GGkc9LSSLKnBiNvwdLJSpLQ+/DKDMoP49WyX3/e9lhPvs7fs/YzVZN+
ZgXlvPfLJdcgMS2wx+kJi38+7IMJIkcGREUU5Api2np1po7yo+JmSugsY1DBYfqJ
njeEfDoDJNAjoVRF5PeXrd1AKK4TET/IsYi75XOGvO/5YzkPlr/HJ7s7qnzmCnND
qONnwfCdyWOpMQCBKOR23oQjhRk6bIn9yXat1EOT8q0uUm9jk/kYn1eIQUYULZIB
T0dJVUjxdeGWuK08At0AP0ETrmvexM2+31DeKR8H8FFglkmTMyecOYhyDKLoan+x
vwffIwydTXTYzR2IedBtyOwep1k986t7UzNdoWrtMBp0hRPLhIsmkN72pRjk41T+
JECbnN5db7ElIZZ6YRD+3QmdgGdNFj6POGax5Yc4epv/1O8IovYYrF3cytcu5xol
WInnISNSmERJ5f3jJR93a4hWf0CrnTbKd0WL0+8VM8Ctn6QgKECkBEJzcYi6j35W
OljxJNW90etKPslUvkXllyUJU8OmcUG/I91Y/PFMXgknXf4ItZvcz//nYUqeUCCU
tb9VICv17O4tLWFQXN6cdIZ5aRlYelTHr4bso1jHcXLYWk4w/r846OGJHn31MUob
srNLuSxJZNXx4iRrxLyfUnoLaqvJIU+4F/YoSKQiWcFEONcotkZdKOslVR0DkZXB
X9V03Qai7UM5D09XdajRQtSMZPQay1L3SHD0VnM+s7SFgcFcY3wBy9j+KO1DCtpE
wkN7mluAwlNXpyHgg0CemyjeX/FoDxUO+mbsh+DBJb61RvF9ezURKBaCIvqohv5F
chtq8+Aq6CZdluaWHy1Nv8ykP3MqbU4p9NsG7GN9Y/1QuT1Im5XtkF0LPDK5gQkA
RwoMFyYZ8GaCU3+eEWW8WRmMjqqfDksDnJ5eNoPNkyBOiEO3aAV/ngR5dyXhg995
SjAMj26jV5MI403ULkPax3wNBCe5O++nDdXmYDlJvZomFonj47NKVXzhZ2aoSu3j
MZYbJx1S+VPtQChi1ULUF2p6BrxRkqWhlcSKTu6asbQsHNhHjm762pWgUYctwolP
H5klbf5jf+VjhLR2gyfuwicuOFOXY//zHCC8+qTIZgkmoJbFMrhQxEAnVPw6qY6d
bvl221rOvCkt/96f5HVzvLGJR/Q442OGLeznaq1HE9ijyMVpKtyD9Mvg58tC2V5q
taa5T/yEt695JKAlHQ7Iq3firau+GeTKZi2zZCJ2fMZNy7VcceNbAozbzb8cPgdz
dIrSzz9j2Y8E2Q5bh2gV9dJW272pdFEL3+NdM13hbZMBd/QJ/wVlHtlTsVVPgKaD
zPTBuXDgiPCg8Gqc19djQkY6ioSTOsQchSJz0pS9NcsFNfeNw/FMeUVlkoI9LCvh
uuRAWVQ6KUFR+LijtR1e5Rk2UdgmPR0aBsq3EEFn7h0OSJEZuxEtXveCXH0X+JVF
atKEORI3NZd95nHipK08awYgXzW6VLeDPbcZUaXIj0gs+hkqt1fK16WQ/4uVXAJO
6LPGFPCh14Ma6JdE/xad0BKJV2vYu241eVS0ElyB4rbk6cHhuJGbj+spFCXfBUZe
KB3yrVP3LASaFLBmV51FC9viUBU49qLVysXxd2YawuUdOal4MVFhuPjOiWvhbC3G
cgQWpKHbUgakcKnHIlTTxa+HHWBEccH++Xkukve+ImxHVNPw7DOqt6P5QdEypaRR
2PGoNPO8/9r0HB1yCin7A3TReJ7JX3CBvweCpOoybnNxDDExM+d5pce0tSX4BWVm
9l4/ULnHu/IoxvyExsFeFZjUVOyPrEoPvovNY834WvGfi9icIDyN5R3V/WD8VSHH
3Y92XHPfpMymhl7GJ/oRn3GsHqTokd9wH5FORMhVHAZLEDc4IuMcbY6q6U3ykiIe
4byTjOfGiLHctpLXQwXg+08B1UUGBipvr1SyYj1V0gAKEg7ZG/wEwzXy9emzYvO1
f2MtPKvqTaNHT9Ld+RKmA+by+UY10aMER0Zwgmehpf8yRpTgb9i0IeEC0Kws0wuo
MP4z0Q2oig6DMhLyhXcJuCU+YwbWxrFPpwmZYToP66kREGNcjtHwrgoRfTaPWgFh
Nu2icAGd1pGZb1ZP5SWlW9iBy8lq2EwYoXnUInu7oNomJdp8Li/zi16mrLkzAqc7
WwMbTWL1ku8/MGEluypzepwZb0jpyM2obokHYZc3ibvKLROTDDn3opxpq3MHiSs6
7dWKMhgJi/NFsjQHy+JCQ5YB84hAZineHU9ZYVJgT1tQNkmjIuUGY2FAmRX6klGl
IMgpCItOrEv1XjGA6M8F988AxDDoAaFZwpCe5tqWVRXyoDU044ZhbBtwrpBBteO5
S5V2ZZ2kW07vZ9NVK6L0vOf2gjWEmvc3mVkzWd+gvpIHwb8syiSl9gY2trKolFrQ
QEndN6m2OsgfC7xcf1WBN0wSJWHV9gsZC7RSq3fSOwzO+uf4uFUM8sPJDw5OCvQu
NxYE94Orh5RCoCqnRvjsyiDnXBGNFVzGTKy3QVJYNrXP4u6ZttoVw2Zm2vULv8rq
m6KkCryvTh8AinhSkb9kPTk6zXQZ5eD2QHv8pHZ99v1kVrKT5Pbmab/et2UE5Fdg
Y6NoL+mOUVyfT0L3WSYLh6oJTi5ptfLEmIoAAW57s1WWHhJvIfD7nWk/At7S3Np8
7K9vF25iR72ayiT9W704oheEI1zjEfQNSQFQkHxxcQ0OFg0/zR7sSKpIqx9A1433
ou4ePIyYpuOusgzO3KX3N2axIE80y+O5u5Zmfj4obVUlVHKLI1GwM7fVSghRS8OA
wFklPyQexNiP62nq2rT/PGWStMAc6ngGqvyu0ONa8TpzyBTLX6HIfJhSXx8b6p/I
qnnP1mPHblgdDdl7GeWbJ2o3gB0Tk3jXU/vJRdIeRFauZIjzhb9ufw91fwcTgitf
cg+Uyv2KLywYTpaUbGOCxGV+L0M4nykyaSoiJWhUQWkm9SYyMg8XVSRPTZUszHw/
CKzy/1JCiZk1/Ak5gZ5HWsTKiyVPJA+0wUhBPUSqCX1xRvZB6lNfHOLIcDoajoX1
PddDYKfxKBlOPDYYBW/DeKbTXVODq/MITbZyUfemfZMAomoJIiJTn11EmtjoMsQB
4weuFLVsnengF3/xNzv6TBb4U2kJVS/qCSvnZOYrwHb/yBae8ORsJIjSzToB/dp4
nGHDgr0dXrdwBis/ia3jDI4NvC7hKz45h7z1YbzH5nCxaLxs9IcPzd47ZI4nv1uH
wtx9t8WVvgARRZ3h7rgKcDRokDAua6yS4ErgS8zyauKDVQV8ib38QwkVCAgNMOYk
us/GhE7thEWFoCOIYmRTu+A736dQ8AkOu8xeBwVUQYeBXi3d5Q4FwS50MA0VQDLa
RalF9SGMtHZehAprjtwwIqFcPNhR+RRmonuYdW/2jzh7bVPMzlWIHAIA+6AZa+5e
Kq0aR9U2ww57mywPtGA3QUr5lWLu7+IXcgY5rQGPBbK5hM4+9ee/z1IaQhKLqSWf
N6kzhQvTjh/U54z2cNSZb4hoIsMfV5mIkQ5IkS/lrhI7q9QchTJkT9KMq5aQdU8x
VLui5uhUyhIJvZ1ZMb0ZOIDpEolG9fEwTj0ERPeZkLDcK+6ID2Roj/vvHTuLPtHi
vL8tJJ/Yofl6CfDP9HzMNGFhRuj3p8Xm0NoD7Afl+LLhmW+/tmh3CoJOJ5m8wciR
157YLW+znQwbZjZMSFVceFjkuPNzBgFNkk9sM3LXuqAaoWslt3pK/1F1m7mCcOqI
/JR51DrYzf19ZC/1tc7pLe8RQ5K1tXyFHO/qaCQqnnfFNjwIanyYRARPXsUWux9I
VvHbsZvaU9Opr3T67Khz2gCK2ZIeBTC7IrvbCjCLd+diyO9m4nxDO+MqxmGyZxob
iljudEubO8WdixxC4TV1URHx87+Pmmw1/fLP0AgSCCUMe9PEwHfoz5qQySINTJp7
DpDj8NkG8m5vdHKt9Jq0pbiYroeOayUlz+5IlemrZR/UnSeIXDdNSlSNiSAQ2WY8
qHTZ/5Sr1R8P1N2Xav95J4b6X1xp2lP+iqheEVB/bRUAgKc008BZSKW0mpDKHSJz
hWZPBb/kFjpUZXClhXlmvbqNU2By4jnoBQ6QWm4fJzkFU9//BPD3zSsRZDtrnsfp
XI2G+I5Yh9/8O5iJvdCNdwGDZtVlXjc6KXeTJVDtO1i/ZqrVz+OwXvVhJdG0RopT
quW2gBw0BFnUCZeOKg6IpIUt1Pzw6ZrXjkUL1dIO9zPYUpzkR7c00jwhsBkAPna/
sOQ4fC83JLqFqZPvEgN3R7nlNHec+H1lLtRO8hekVX18ndC38m3Yre03tL9DXR4h
sYfCDw7pIB8GEcq/8vGIskfQPXcfRv+qCbOMRzE56uNoxEl8TcDgxRXcLxapznWj
yPtsx/i9She3AvM7LuB+NXFkLawYm4vuWUPjqaaLeLw12R87l9pzhznfiLWIHB4y
ehaeabznvLwO+AcQI+nXGM4CIp4R0ipA2O/+sru7RNsjO7tVKIoqhDqB/8Pt/urr
3VnICr/reGseN4Ma7J5aYg55uBdfxHoSOUlfv7vYokmuiAChjziE+t5aeDXBYQS1
PQj3R31i+Q1dLtKeLs767a84rVkDrsxYZxns8BkgSJ9TUlk5gBcK3lhMumLeaAz5
jJNQGn/ckfyIeEL1aQt1Ru6jp9l9y27REYh54BDuIJAQxhCO4r/8+pmvi47cyJPT
6jLG5wWNr+IbFMwTcYXsx+Lrr7tlIRwVJ/HvQ4YnBgN5bpPuFriHnNWIt3fZcIuA
2uy2cAvitsdu+MbX44p5X2sNi1Mvl18ZccTA+PXiLp4KF+KBJ0EFhSn/H3OvxOkz
6OrM6fFcMr39IVn9EzTZJzo9Itqmq9+xsV/g78jzQoTalgtncVUYHJMxYdEpA2Jc
LX+qW2xsa7yGfwkkD05kPhGiWpZrGR4Ejto7huWo+QyUbdvBKYs6vn7lE/jrd87M
o+oy8RDVBXMGkt32602MlGi87bnj9BehtQPY4/kJ/Q2Co/eJmAuEM3spLNo8rLFQ
+faCKWE0F6pT1ZuwxrBcBbwhxlas4j4uTHQOE0clGN/1xb7Two6goxSz+YsL7ZG6
FeMpK81+V1Qh4DUv4FflYPg2fApM1OgWxsfH1LFwK0r6Prpv0jP9yiIJeJ4vElgH
lMwyrNCbfeUaP3Fy3KIEOz4ifyZ1eDfxjTc4hnfVDIy43DYe5EexeZSvfzYJVOOc
NWEK+V2ZRZozsz7ZAGKRjzHTYObIA/wNseAAl5inMwhT+MFlOanvynyGYJk3fM1r
XeBGirO78M+gdFnk1nISvPkbHhWA3ipEEMSOKtpoAZIZgd469/kbwCAGC1uyhcW0
tRuPP6tq552nglBP5WB+cB1R8PkVT3CFI2brmdHcOJ1lb/rmNbTDCoOQXIrO1Iga
kvLDWaCiHj+5HquaeaKD38B/KXcOKqLhGNZlPgWs1rLYG4aZqw8rRf4zOeKF1olP
gF110eldcXIhoHDTRuvaVemNx0q2QE+zzBS/wtxfdOFL19ilO5lfFQjWPkEA9ZC+
aLV+eY74vRJ+S5KG6JWrxwiR0rC4KOTQ73TnAIF87mwdsH9+PgFCkEnhHCxaPOP7
zEQkuXVs7fA8aq8sHJYqeNBMYBei2jCD2/3XAeKWD8ImDeRttTWCeDOygJqprCu9
xSHl4QEAHtbVWMtXkpooLt9VZwTU0Ec80/mySSyl1NH9y78C6NjxH4EksqmvU7Ff
lYVLqYdEIaZcwlDejzga6umNFuV4NY0lc95DvBF66Ev2jeIQiBD4kXhZHifSWW7g
scI/+pnU0jDRJfljSmPYZkHJJpk7vupCDtAs6AchIovUQmkzklMHbfTgy/i0USxy
pLT/UuIuf1VjK1DPc18kHdQvzBlpEKbm/8u1op0kMu/7OwQH9POy0Cdq90IZeKrl
ewZyIe8ti0rDsLfwB3MsiQJgiIFJYFgS2lo0wccKKUkMgWpa6Y91I7WxBNymhEvI
j1Pk1ovO0NoXu7c3EbswUw==
`pragma protect end_protected
