// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:21 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
boPa7ZskO670IPVuGCWYi8lyxWDmJgHzTW8PUGSz+6s+m8iS8wPd5ug5MYTdxKcr
Y+j075l8JVVFU2d4gI7RJ9/wofWfmi2FQNjesSluEThu4+0VCWERp6qysW0Lw3aK
7JveUA+uXjRuTT8i3q6+fVj3oykyhj92XeztiwQePFU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27808)
x/6GlLCNjPqygM1pVgq/aoV9jAo4xpK+ZFDCNuiEYTefWGQ/0iIQb3xXGTTu66IM
77PQ+ztu8J1qTE+mEMAJgL8Ohe0Q7aC8K2X8Uk/rCa4kPzT/RylsOR4mKee8IZ+s
fncdEEGoZJ9pJGPIBeV7Ye7fdgghPq3NmscB92OGQFk5FMbMc9hdN3eiWPIrLyRs
k4++Tb3NIiRpOEWruqg+rToVTW6dFdNvYas842CUFVB5t6kcTo+T05NjV3LIETr0
a2pIDf5+j9c4a/SmjZUXu6ImurFU83K1cP3SncJl+X9gI0LOY8GoJx2Ds6xYPc/4
LuGNF8inpHDXXh33CwnlX58JndQQ2H3w9MMMaE+OMgDEmuA+zZE95vF4jOMo2gkO
LewWKHgDl9CHjZYPLRPN9GYPAksuxol+MnKyPSm1MX39699u8XSclAadoCyPezHz
+39FonCbE9TkabSP5u3oORqujkMCmktWZp/RxqShrfqTvmiOzfqIuNQeze/Xaq7V
zy0h6jCcGzBdOGXhbIWIrWYCAGnITJaSt4VUKGzRz2MnM9vfC1f621suSjkJJTCt
g0fcdqKQX5OdcBZX8na7zfrdIW+ZbEDvgO8bUDugqqhhGVE3es/EnAD3HvDfyj4R
D6Iu20QN0DhQWuE1J7ia3U6uinC4w9AwlzVTrzgMIyFWO0Uogscit40gnGqQa3ew
XeC/+xbUvp7aC8hlpK7uG91MI2dWkE4jQKgSCK9vxI3C1HXPdxdgf0gqRaUhi7AM
R7WPh/1vRxRqFzaf8fHRIKWrme2YlBtk4BDS1KHlSVWzoTfBVZf4t5e5ZYf/brfQ
u7dghAr4KvBsuhXKECzgczjnsY84/sC03rIvFVJ1KtK0ZbHyd3eDHzIJNv9sANis
Xmzax1xwClyTsJlI61cjQMuLXqRmBAhOwy2MficJG4HptdANEsy3c4EQm6Cy03xp
/9bnyoZKhVE6QpvaBinVP+Pjtri2P1VJBeTVT6IY68bui2NfJcA5hIwAAe1hBqsw
gKC6aO+5+RnG/HSKaDEz7UElUxfbuZMt/2CdwCDWAzZMsLz1BxE96WZt8w0Q0xpX
/7V5VM7VhqDYa/golQllO83sN6MS1HdVgzyK4b9NZ0yjK6R0EbVDi82FWXGLhwLD
Z501sEMBORwPyqHxc3PYykS/FXRpFptq6bwarV1KtmSto4PohBzv4grggNVzFLbe
LEEhag3VDccQ34VzLEyLJxZu2B3QTWP1i4lOJnbs/K+Ky13n1cAjDIv4vIXXqiYa
rtoYtapww3xNxtpNoz1vJ3I246TlmoEFtvXtAY4G3EFGaA3xzXgY5GTsZIzrWiVO
SYxogr/0nl9MZVCAZ7YwxNFq6RXK65gQBOmjLdj/u0cUwdaD2bpepamnv8tMATkF
3B3g6QMC+/2vRCvO5wqm//B9dTxQBQqp7vJ74pAcFynpZyWaruBt2QH52FQGPfEo
R1dGDrUCNu3ZjgOlyAeQlkSyUJvpeLwyTKwpwD1fGds+gcUOzxcSsyaZTo/157OY
sYcFNZGMr4Y1x/+9I8CG7SqlWQeOMMAPrKzZv2ZRTDA7bsydE6/CAoV5OT07ObIT
cI/EjAV7GhDtpfx1n/IsKcfdvMsG9uX6fbHjhlWgsskSZlSiCiiZaLByofHcXeqD
zYcGw6RukgH/vvVzqqEJAXn7E2fdRr/WQuA4/f2ENVn01PnV8WPALc/FO0rpAj1W
8PoAp4cJD35IRHsqXdckA/udhZycuWNGQZI0wQr1uIP1nDvOx0/kCfxknexhDoQy
U3hNzxYm8Kck2H37zdfs7/VCXIi4BCWn3XCtJW3ZMCfJEMGvHByj9XEAAEUurZar
qbn3p9z+7g60U20Lnd7VApimpjzU2iC+uIPc+YNNtukljjrV3xlUIfjADhqdB8TW
hcxrUliS4swr4G4GyC7EqmFrbfpcuDWRQdNcStolnMsm6Eoou83/Bt/CzbMkGKky
2ahUcMQpxlwyz647hbLoWjEj1PzOpd59TTZgMB7tsSPiUUF0atZvCKkMo7MQIcbJ
HvCt1SpyN1MoXJT/U5b6fA8S3/KmXYbwmQHq/uUpy19OW58Lmyq05pNBWa98fGP1
J3CBTZgvoa1ILI5m67vmx9zLvWXGthRnOlnKHXAac+B4gOFh2Er00F6EHzyk3lT1
geXLEpm+s+bQazrkDzNYQKV5+oy1P3IXkZp15fYp2KZi0YHaHYBzVhyDbLNNEmrY
w3W2OkbHT3TQFGv2QjL4t5kAs2R22ik35TTWJ6ehZJi9eYO9eUEPXwaYANKlUpl4
DkTIC4xZdLwf+0dBEiKf4wXIvqeEX8aUex2A4KsEzq+519zo4jD0oinFOWtoFghY
8S2lyVLW5EBS1Z6g22wBw7peqN7MbLVUNi+i/LgKBi0ALQ3uNPLSmEXu1CLj/OOr
SleMGMeW9bdDhwC6QoUlg/NGOGuo9kkqiJJ2Gf8GVqgpwb+z3tSDJL6TyDOWuTTA
++DrSFEy4FZDDntrbZOskIarNh3QHYluP7/et03oPP63GIHUc7nyRGbtqi5Zr0nP
ANq2HnFTavhMr+TVVt7Hfxx3D/dbGnNRCjQg+fmx+jOUEhNATnZ8SUl4JA2MkuEp
RyeAablMuM+VDc0fGyDBKVTbhhOGx8w+iX3abjQsFpfDs/Lb+o0XUopboLNBE0sZ
7Y/b3UgNlq690MeMbBUtdeV4S+7ob6WGXW+Xs2tBr5O9ga60gPlQwVsKCRnWZMEE
PRNoIDXY44BQhqBnqMpF6lYxdxS2gigfQRjz9qFK7JevLraAklyyuyqNzT8T/BG8
pW/ZVvxU9/95+a5nO4JFIcuncqN/CDroWg3Do9nqSA02urqGose5Fn4uPOQkQ9Hs
VEqv8Rq1Ndpl+q9nAhUMd5IFTZl+XqJ9RPiGUrSXLhRDjdie29EQEAw/D5zCIQxF
O7zuguQttRaDelEhThbTc0k1YZgzimla91JyhSTegYENhB2JBcZB4QeTxc6lPKCY
S72NgeVc9mPgp53Ow58ptDoSNvQZqaHiVS6q8Y5dqH4igzA7ci9OH5gTejAGT3ha
ssHx8zDliFFbGnDuaQkwLVBPE+lXc/1ye6Esoj7Dt+9mZtpydOxxL2pEB9Db8KGK
1LAUA0u5Uqu7rQlGSw3hSR68vZ88AWpmhjSCNmtbiZz2nan5NicBaWnp9959z303
2GOYTIZdAGjre8TaQYo5TdIp0mgQmNPl+xBHL00xEedkHBdSiR9knK9ywWaymT9S
mXGds3ATnxNhiYQnRZvhYCtMJUQSgz/FcATiGDlnu0eo1H5HD73LJo6Uq0lriIxQ
F+6zilxiDUbopd/caMs82ikl71QEQbfMIbsTfr4X52eK5jUSAkWK/n+rWEce13H1
neIMbdCgAdfjaMvyPCEs1IMUqg18q43VhLsGfLk56GFRn2OB3G+l8n8R6P/wSmUX
BRL85CJJaRX8b88FhI8P8HnQmGgq/OMetZ2ncBK4s0tlwYy/7Iel97ddicLPII6R
xR8vUwsvA0Pbtj5yJ2gJ6xqyA5kXqyc62Q47XgPTdcq4SjPpob36cF/2lQwzx2Ij
fSlQuB5DETeaSCAMdaYbBwHuwdb3pHbAMtxWH8HZu+nqEfQ4OvVrW2dC7UK8SR6C
FKnZe6E6s3TiyX29TNskmN51yLhc0i2iDhhqxfktgiaVqnGQ15ZofqaTKKM20kgU
nVLS4TsJcc9Z8O2s5/8gfYATsB30L4kt520gisNzERHrWNCo8dGZEJfxHgZ5fT1z
CVQclFoEuqOi2AVH7gBAKLzTynfX+D+5fzFc4yrwLFcUkiVB6mORGEwa2ct2Da73
3OnKT3Yjvhlz0Qv1ilMAPM+LIcTWvAeihZw0qx5yVh2nHIfeR9sCkZqOFZwcgdLQ
Irq3RyMDiEeM0tHvWoshAvNqNjjxi0eFxKWFY+oyMMbNHJEjSKHlYxTzFM0B6Cyv
wTCAjLBo6AMDjzzDGeuIR7XrwBTuUxOTFIgSuONN4Fr+hM9jX7XxEMatY6iGruAG
pTyTKKUdChoi3nr/bciQHBu4qJ7+uc9f0EIihHpYXyUTuPZ/ezgbONO13ba8r4wo
i5UWDndpmOYXKt6Ev2qrXNd+VazAjaxVtiKE1siriW43gJX8WIW1OL/80Erc1Igd
ZkivbU7dr2vr2L/YvXVre95XD2A4wV8E2TNvCyI1FqXT12/Z5VImQ0tRESpZExn8
/1unsPzNbWEWT/kJFTqwfxjUm5Ed+e+fAccErnWp8HJR39G0sAK+ORo85S/s4bge
bD0irQ3uLK2PfDX/QhknNVM4cPLwX0bxOTc7X0BNfk++jX1OE1sKTdhK92dEzp6f
9pnh7XGMvh8fRAtkssAtstIV+AWkxCs8i3HewPen3kzN7OUHgid6jhoU5rmfUFA8
nY5/L6989SoNR0VzdJlaZ0yvPiJiC5yEXN+uzMB1XjTF+Rkj82VLf3wNGnhJKEsu
7cZ1a5r4fti/gkvnweCGOL+2///HtpLXsF7/15uh5UeufVu8mlZtxTzmrsSBaYVu
Y9brxUOsdar5w+6Spe3ltK0gtlUWwzfrlKixyL6QfLheWGuY1a/5o7xNrt7Rf1so
FqWmuQ88z70gvTu/cboLpa9AoRX3tDMGlekvka9+SkQ/DFp76vyw3ucNrH8CXjs5
Q8oh3Y0gHImcPEJkWnvqCAOzY8DPR8XiKTW2bfQLRPmKFuwJ7Udm4YJlff6OUybB
X3IKG8pehXbrv9WRj1Hwi35nqj0RILJ8e1BJOFflGwrexqtjOrncaC3dl+pOPnW0
T6C2jGV7ip09M6ddTYS8hWVAohYFp0ttCj1jznMuJX5eXZQ3jvickz1mWaqq5HjD
/tD+9HvXSjbV/hRE3D8DcxB0Q1o6TpMkgl0wWjnTo/bH72g58kQOU5m+g2cUpC93
h6KFJL7H76nWmfWu/wP+R6lZi1GIp4/jiqGOxkg0Rw5wQWipZtge1StbQ2plfdbm
xb8xcTEA+j/aj22VU62jzUFgp6apBTKqJuAbQeoAqst+kIt2ykP8A2aKEYxX8ZYy
nXmHCFZtlQNXd+UI4D1z0GGNTectfioFtFgGCwyPC4hR7BmczIZ8/vesfaMRgyvh
UKFVCOY9Hpvuh8kkBRkH1qBxnac+fNbyDC2L0MxHIKRQ+lvk05lLINVJZblZPCBK
Kb+3nQbkJeSoCIRMlNH9hR+ANsCEVNkaZv72nBbDbHEcdBD0kqB2X2bcoO2N9u98
eau4PcF2s45C0kUgu9UEnVJhP8HnsMuSlAINEsc7RmMTR/SdWNhLmetNgiJKII2L
/RmZcOuX7PQxcnxsNNRBLjmLJkzYSZVBQoctRYhFv2SSg35rn+rWQ9TNOAStpol+
w4YW5EmameX9jJsAZZdD7vlRgxhW+4E+3y1DVRjKqvJJ9cxpTWKs1FIKCp142oF1
Mh/DpCbxy/qYDu9Gyu87gBH0y+ngGv4arrqn5X8AmPHyfPK+I5fZrxDb2MUlVkTb
ZCObBorctUp+7wsVENwUai5siBIf2ZfOSyjFNcnyiydTcKOclEJs0jCGbAKB6rEs
mfRD1fEWSmaiRm0TM8s6AcgBfrlRdYeZLt2I7t8HNcPBnXAu/Gy9WAe0NN8RjMBW
RPKT+HcY7VE6jSU0iFX2fiInUBpEtN2wLfLzlY5bmzpiDgXLueBcWL8mxO29/gkK
URhrBIU6U3OJUABDhh9A8SzHSbHYMU9bFpYnQBDYPqyg1Kx0mwggo7DubzQm0Ed2
TyytWVe4x5GZiXBN9rrvxFpPWpiOboFlbM4X9nXPTmL8VgqJ+2eW0rTSXpDWUUu8
XWInuPBj0hNGN1JHP3BO2LaPdhmTyrbP6Q1eoDMofSvcPm8yJQjDYpxP7fdL/vzX
WRIRejI/8tL+FN3/u4V0YQ2wyWyWZrKD9ejrIQhPJUTecqzR8HOUfM0iCFAAo6hc
Cw4M1c26TtdKrx8oWQPV9BtimwlTAlPip1Mz5hdphS11+SUqDCrxBqpiyz8wx2vw
CYt8jGdZdaPhRcZGMcT+Vzd0lPXuBH15xTgsODY1PmEjS7u/pgylx7sKgEuP1Tfd
r+/qnQvNkOTB63MicnYxk9s4yWg9dKtAZtKrd4Zjnkd+VwlxY9vKf7TJe/Kdww2D
X/8dSSCLhw5QvWzbog2YmBjG09+v/lFkEVlsKTWxzTwhkSVcnoBcb+YMljYaFfSS
CAJ5onbSmZEGoRh2+zXi/N8MNOAQ8eflOSDKrYgg0dGShDrP1qlJ5GSLA8Mq0nY4
MXXkLgYfbF9+LtClih/2WfNimQ2oVp1NSHNvvbL4ky26bdNrsa/LkmwfAJJ+KsD+
+uJPNK91/XC09nwpN5TZ/ltcpk1TAEI3oUYH2//Bzz3dOI4cJPCJEyRyAMi4mA19
0bKpE5Za6rXFbkEm/49910TheuraFBBFKNzzCtTaR5lBKrS9SenqvcIhEn2lzu3O
VsPRoCkT42NHO1kxNazLl+/XTLBfUUJSn3lyf0eka3Iu5Vq+KOEWcOudmpw2AU+E
0pMfirFTWqGwCXoIHYqhQ9Nc+oLp1wa2WLXKikcruJf3VqfaxrRJs/WeUjYrK9+q
J5SMZM1YpqY3B6mb5RFEGeYF6TNmvaed9FJ+0r+mJHo+JNWQx8cXGEIRC6FCx7FC
kLdl8hU3FyFAEKK+vlJKcvZfgnl1Jvj6TjnTL7uEtcxAUSP0ieUMq9ePVO0w1mKn
jQrVL3Lq7myKX61Clnxaq36+D7xAkGJyLKNVSrW3kPJ96FLSRt8KnmLhklBbglWq
GYFcvZtHL+348XHVfw/7623/Ws3oydff9Jg3JUE/2ieJJcu85p1KvgWRcNkDi9gm
ez80W/vyVK848Q6i0Ok++ChfLPQwjRoE7m26bGMvDn0xR/NkzOVS/496YRDGNLo2
uyEUttkrnQ7ZttG2rC3euuHcb3in5x+WkebqZtd5Gw1vvMTNOwpq05EmOUHFM8pG
OSEmMFihkQJf91An/gKdmKrYvGT3qJnyNFW81dI/bBzfbSEU4wQlRcQj63gaw4+6
hNzkRYh0VViXUnE0Lx3WGGDjcOWiuhnnfyhQkEfgyoRFe16rAaw7815oHTZ4BwmJ
yGLtX74Yi0X/PUyAVBbDF2dB+H7WKsvEosXmVbNnYr89U5fKnWuS2m5aueB1vrUF
kD1M6Xcq7S36iwMz4vh03inG/8T2NKqioRcsdl1EFud3/f+KcfOsqj8s0gty2p4H
UBj9PbtDvdnXYeFkeTPdSZZY9buOnFQPg7fLfhcVKhuV3AXhT/TqjQbJcHf0d5AB
FtsMaTEr3hrp4Y5BbtvdB5RhRGW67aNWCIhDXPQNHe58Kwtk719YsblpGBYaAelK
CvHKAOdmoikd8UrHZLrTz7gESB1LoMQwMJl1Ak6fq0VgKV88FpxbrE3lufMmXHZ8
a6SislrhdJeXWrxqN6q4/dCrrBqzkrO4gzNSG9OvW9dpxVvWA7WFH27RDK0godwu
uBeg+LXFY9DxYWde8zfe8clL4txb2ieJYEk8IDVLHO8WFCCEzTjJYTBWGHXjf0mQ
7eTI1xcLKibhtrfuOxAvgszohWR8NKZxzmdZUS3n3OsbAfTX87lGQVmHqNjmpWH7
IG5D0YZ1lfUae4o6B6nREZ0dcZ6ZfGO3JVW+WaD/Vmf89OdLbiqlnmrbU3U2oXb3
4aGp9baAo7p6ktZYTAuR3o/WzWzDC8jdoVFmvszP0OzZ/HsKQDWhOFRfTdCFtWmk
PIG4myfKYaCAU6ak08WfVOp88sE64ymOz/JA6zwgKFDh5R3gnzLh4/HPO6/i6ceL
B3MB6WaOHqOF4GhCKa33of6z9gh436a+mzVGH5YXunEv7eVKgnARWRupKU5LfxFH
JENi6G2bA1H/rZXJIJ7TkD7c5uNMldbNLf10hnE7LuktblQ4sVy+unucASmWCjF7
xHYQ0GVxyTqE4ZN7FGvTeefs5sq3nJP9J6MqjCHjAW3JoqTXnB9HDR4jvsCbIUW1
lHpCeQGj9+0AhCD0Jahovi7J+7VXaIrmmm2wcaaqNEB5mx1jOZAmvvuEAZn/R8ZA
Pz2leUfPt1sPFM+91BLrSHtyAmNmgeVWiTNEoVp76ljy5lBM7BkXJhRVgzk8sElr
8xQ1gBooEgmH0Dt8KkjcbDKSvTPfRKSkNEZou7oyIi9i+KBXrvWw4sRW0ypNCiY6
ztWU1VHvjhzKspIYE/29l+ZGNPmb8FeMAmy0mPlLkPFV0PGitpQciIQXGqIYDlLV
s5L5FNMIE6WqRCXdyDDlLYCUUoqLOSJiNVoTw7FgFPKfdDaN70mNp3JdziJ+yhiE
spXT7smtg5OJRhNmCfdGXbB0Ujuz3P6EKkU81P1GV8MiOPcSE38ICwv83JABCVLC
YdBuhUjlUBaA4uG9IxhIZ1E+tfTUYyqPRH3jIvoMruEAkpll015fs0cJ0PV0R/T8
PuDvWamf8mKJz9mXHqplL3VhVdhHLHDTxTeC6A7w/CyDVJgL6oVpxVDbarkmp5sk
oRcNluFYsy4kqf2xxuvIzkxJoyc9pdCnpR9vjt0UZj7Onbao0aWiIwHEeiK/nRl1
w4wYD9cww9a0EjmOSDKNEMXW7+uqdu87uK2dqflYY6ngFp3NjTpaaSm7FyUtwtG8
bEZPxLeCsc4KrOx4XEEOInYF6SbkAuWpIpSh2qF6q5rB64gnY+N1UBkKtmEX756J
cKnFg+fSuKojvhwGal1wvWKgDhVE7ZhwHGwSR5sqUPxGnsGhU3oXLcux7m9MjC4d
TKGlyzJ5Y7kFbFmwi4QGramAkLMdNUzmhVtFHFi13wUcu/gVdckqVj8Ww8XwdRaV
j6aXVk9FN4ScIzSBUd81+iXfUMLirH91SjWl4fpyZdgz+SID05yqfWjrFCEvxg8d
I9VxG5y6qnwv5kBa885me82tb9hopyKGbBjRiMvTojydhGUktbP2ZrmKr6KUjfZ7
j6mg6f8AuJWGLhOrXe8a5vEghesjd8JdnpCQCgcMrHocPRxKXkMNUOyvzk7mazlW
Hwu+B+bmSS1tHPPZHL2FUm6qrYpQmeayevVEC0wJ8r3kwMqodtb5cg55A8Yx35Mu
CekZ1hWEBPUf5RtLqU3DbnjMCiSnYf4Hls2nEqtcHTElOwxEvRX1x9O10OqFlBkt
yFhZbQHPeS2LRaknGICsx7o+bprE6j3IxzQaboYS3L9sn28LekTpDovNi+ZqHjd1
0+LZDuQgDl5jQL6VJ8Gx8ipmkAc+yR9ODZx4I16TCo13QnIyA5WmViQMm3inA5CM
U7VMJsuU2ylOmfF/Jyh2itLQArNeWg5PpHIZ80iRFs9k8nf2t2kI6Eh3CqFr8AhP
xc/YStboLGchEuS0r+qIMsxY16jXXJXSZEeDBvZMkijsb7JJolqyAbCsPuWPPggC
dW3EJBYXSPwcPcyT2Z3Mvw4cyz52ztAbBXLH1L0tpwQAQL8BK8/spyWxhEKedrm+
vJnVo5k7CZPQgp6L8fQpb7Rqb1YKOOvKxvZaBfcWxsear1T56XlvJBf4hbp2nFMr
8lmaC930AD6I9s9v5D8bKzf4ZwgMCpxgBxu9wTkAVICCWSQCbAlAD1uUtoQP6NGb
wzIChFgS3LWl39yS+HqvEyT/9P5taVMn6vxF6gaCNPCobZPrsMqPFQk3DNCZa+02
/QVp0msWw6oAuRlKkxpK0SMkzFaoaRwGMooYllO9ZRXuuBnrtHJYNaDQfPa0pzPE
9+90sdnx+FsYXBD0LcH9Cu6DlS3Oi2Xnxg4jKZZtHH4b56sFAXEwE/4rKvfK94ad
0Cqcy3cE3thbpUnZ9d6qjyLPr3RJqFdndZpb6Z61ehS8809SsTeJD4UTnUxFn7Ty
7e/IYZHdQ4Xm52SNnRkaDdwz3C+urXHkJ9XEKsgpQqh2R0wtE2G+YW1w5aSlxcuE
h8bprblpGd4n91TnEpDxlnXsJ+XywvlHwu4kzT8GceJgHBloIxo7WV9Mp+ddabcP
9ijI2oG9FcczOvalcmdOsrl6Rylb3SxQL1vSEmuGWoTRbsbgS5CvwFCi8e6HtSlx
0gaDnF2XKuKWbPumCzk1lBAGVvvPoSL3TrpLWo5F4mAXQOYocz5PmIWrkqUICz/N
nVvJWwR1UC7ejV/T2Jgd1JbVhjje6N6VI2pDOd5bh0uWWIpVj3zcY8zPCnXDP1vJ
FCXPqnNCvKQDmHkqbR7iTw4rAoaXQv81C5mGO1fLjTw1Mb/9kbMYnVf1YpI6TTrx
sl0GFsLaqS9THMK5mIvjuZvpVRbhIXXIiuyE+m/kCLatWE0CHrOwe0gRT5V7ar3s
ge99IZH5t6UPX7YOueA2tmeMNswLKjz+mgL7SAmGJnnn1qG/XincLlOGrHjTA2Q5
Cdw/M9W/Td9HbWQxs/hEfTuZZDKA9rbSGrqe275uGeOEt56us3VXE8R9zwKAHsgJ
dRd55aTDhJpxuxtCZdiv6HUlk85/v5uea+NjbQYNz2QFZTmy8ZGJuh1ozlQ+aCSk
pXJ/Tz7BbWoI2RrM3APK7T8b0gCU+p4zsAGODHDzLfNWUZVCvU7FJv8exuSCg7Dj
Xp7GvPEAEIukzlOWPvVD85H+l2qXrwYJGEobXqY8LocxefTsVVHI84Vlipvq6L5P
raRja/1WyO8D/lgnbgEzPJLhPL9HKebgAoOEAQ6czqMd+rfvt0HNn2QfqF3e7WIS
OjcMKH0TkY6jbI9p/IKEJ2cEkc1ZlAD8b4jfLhsBWSKIKTZlPgV4oiWOzH/4km8K
t9IkkOfAXm9/RSdRnKG6BHwOxioGGf5K4jfI/HqXyAOR6L6AHsR6q2TTuXVJ9t3e
XF63ITcx1xTbB23jycDGEJJxWkvcOqDy+45HRfbspGLNbK+oQJuihWd7zsAPc/qn
Opc7hW1aMQCWvu1GGhlUzrbqJk+vpWG18mZ7mDqhJUH4KXLmQ+m3BZZ7Z6Ilupkq
TYahzcUi0/lL2+cDwicMumASq/0g/8JTGwxeDjNqjyXNlSFNJQ8UC31vVH+szmOf
ozuINmOhGQZYQ+gaAdG8qBpL4iDNByvo3mzCV5O2Zv+xMrs7/GTopAcM9SnSKqpR
E0PIE9QSU/4eUht6hKbLEWwDF5nWeOw2B3Macw6yGSRSezTP/hopB3jwkxaedZ6c
hVwk/PvT2iUSeozPBJ3Bjs6YGkzOY4dZuQkxj7I4KmbPwO7YR+C7bizc7Q8QplQW
R6b6C0KEKGUd3jCpKkdJOMcLAjAh2b65gZ1u0jpOBhJdHmj0zmZHe2lYowxZZybG
kCr6+Pe3oRr8Dj58hjlNbZoJXlpdAspvQewVbb4xvuua/tfMIcsByvd5vO3znaQY
uNIAtwx99gcXRzWYCMeWcSxiCN2XA6KtpBhpf/6Ildfis4kuxECjpW0CKiAs2JaO
oKDkaXOiWR4txyr9IZeUT8bWlBhjMZzBrXxEoidu6dZ14QIo4rMN4GuXBPD2oisL
6TzlbT00wmaCeTwJWZPOzx9LrrCUIRH5qO6LM8Vv96tdtu/PcA7NsXfIpXZgOyb+
4DP498q046cdzS5NPpHoXPs69nRsihMN0vcwXggpv+gJOyGHRNb6nIb2m0XfsLp+
avbm6fwUiFxIIi+m3/E6YZEXk6mslWdkZ0468iwvIvFeGmdfMPa0NHPDg81YIk68
WjedEjs24XqhHZ0XnRnT2nkp9FnWnA09YlLnnafYN4hwGan1kkBXw1IsHl+8U7gx
peQAJaD8/HICCV7jQAOb2DlDvb487SDozcjmqJeRokqHfCXR+t8haMRxcsj2QuV3
5JWhSFfwN5eRk8JS0vz/XUlgOHUASbLksuqO7DYm7J4GRzRcwP6d0if7BU1nWwXo
EAeE34lm2Oe/oUvcqorVZiAouq4DuN85NfInjH1GSCW+YO49Oa9wQxxBtBRZym7w
JHBYK7tgtfB4LoK8RxK4aFNWDsbU5aaPYsjjClnlqWvavj231BbI+OQ6GqhDaMQi
4xy8KVGXHOi82q19NmhivdZ3QaalZXnwVWGNSaWpyWcrF+NiCr+fRmNfqNNJ8hbv
htpTPBPJzrgMnKfpJ/yAK+0+WwMirF0DrzKCvECESY9J4ggYVtGnPuLHgQ88NzV7
j7z/dZYnntsQHoUXJv3KD+l2jye7ohKsZVmsbsHc0RhAuRGKSeeixDvnc/CCi9i7
E3t7KED5IztzxZQbcbMOprOj9kNXInErRGNk2QBp5YVI06RHtNX+5RcRry9fb/hq
pGuzNBYxL3rkXA9y/IS8HMahXwJ1ZXBs6s48szhhhAduUyx+a2bvY+gTe/crQYmW
djzSUvrGXqVaI+yIJ+d1HfApqdV+aIl15v7JndfAemrLCKpNC8f28CKce8btWT8z
dfC5U1Q/1701C7zFruNHTwgQ/zCRh6PSohI0Wi+T6didBwylkQYu47sn3rdEeUaY
8ON/RDyRjAgJ0QNnN335ChnPyIHbmPdtX3olawoC7eXdf/FNl3uJGfv9LarxvYKB
QkBe+s27x0xzDPpxjxAeTQTAMVRqdOAhaiKl805543DM+Zq1dvMQcVuAZLm66/7L
zi+wQWyNnXgCbvQaI5KZAU+J4OaoPI6Sg0XotF1Brqvtw5h+lhzGC5uCjGPdhjdg
kfUxcYk2NLphvFK5Uei5GCrACtj3vzwO4tPtZKHDUlnyvvbXnSXvNP7rwin7Jtnm
FQWNrxwBB3eN+QgqvS7bzyv75YNjhtr/abouMPqeaaFzPjPdZDB+tZhrHapMOkX3
TzWQtyPnIScj6eI8w/krU2yLQ7bYZda4C257kJWMKe4s8fBY1uOph6Z+JvMhLpY2
XYU3Z4wAohQr4BiPFuXT4Zm7q+4VrMQmeRVBMH5OIxe4W3IxNdeNAMLQYtylHwFn
fC66xhiCvAFCBSN0Q4mH9FWgIBCAfG/esorAkBmDZynJiEarkBAuhv3k3FHyP6rP
OMoIrkj11ez/HuKDmtHKWI8nO/Xoy2ON243n5LSnQIW+e+AmLs/mXEpSaocmRNNL
9tPsIlQV18D8RZfoHBhEmEPFyavtZqiaFtygqs12dm8Odu20xPUc8e+3SXt+kbRN
5D1IKU9w+Rqut1jgropxNKiceRimlT+m/lqEUOZYe3uS3d36aqddSjPLhC2b22vM
Jmr4zMjIZYYsD7RgYj/E/5yrxdtPASck+EA0Slgnp3d25tIz3Z4yQiLDx48TZ0xi
ADJtc/XWIQjRWKgFhVsPHTAmnzzqzW1LZ2R/KNOQcqDOQUSzHawxU//kllJCMPrx
na4iQjLspgbhIM+Q4YvX9j3XOMt8sY07FbdqC5PkHVV3ZHDUVO379GOX5qArsOPp
pjENFaM/+lNHJuAB8/+2iDHc7iSm/1fK5cvbw5oQR3aYs3s8wNC4EQ5wkBUjqiRS
Nczu9zCGBOSHkEU2lx/grlFfubcnN2y1793yeLpc4sTwokqXyEqPwq83m8+27718
bO7SeYjNn/eT0qAj0wzaT531zI9aaXW7nMQ219MD+7K4dnjUKkDPlTzYal0PoUFO
z4rdfiTVMJZZGO3GdonE1u+K9hcj6QZyBxRMm0NSRSrwCGmUc2oxED5S1WMFzELw
V6rBe/dAwE0RV04nfgz9FY0qNHYIewK4/6uGYIav8V+V0oUVMoTVIAKlYiSWoJDd
AafLhVcVnJZ8t+hUyfmMIqMcMzgEi5cB3BGl2nBdsAyw2P7nUTW6ky+hCklX5XIS
w6BRN451NVwzhVUMRfDzsqFwUd28QIh3s27w239I6LnuKj3KCVFPfBDhLHrTBJ++
I4+SFTXIzaR5VgIu7IrRLx/iFFnYTa8/X4MCz0os1/Zj8WbZEEoGKtlXuRupTGkP
MjVk7f5VmCzUnqsJGPaHm9vCpDKJWBHwamqQnpBHOghcJftKf5Zu1nIdXeleAVnv
GyAfMTmoJ+5Pg8GEvebBu48dCfnx2MoEK8asLYe/IW6MtEf1HYgeogHGEjHE2Ljj
iSyNRtJsKoUtBi0sJ/wjnSrQIOeEqXjlDn8dhqhrJCCpips8VJuKYael8ssR3ClR
yOfeb+cL2WOakdYLTBbywp0IXZthKkcVGcYhFm/VRqWHA1MxXYggubxVJbHBzNTp
lhhveIMxN9Qr1ImlKYf7XAWGUXcQ0M7/hs9cL/MbdxtQG6ZaYLpBjcDIbXYDUjxD
j/+F5E0b6xrRpRotF6oPg9ko3fEzp5a4rD1w+UoLWdy4m84woLj8zmDehOdEF1Lp
6aXHfXCnL7KxcKU5Cc1UkJvExsc6z6DOLLN4dqrHhsCY0LPwhcMdbD3jyjAYEW8H
u8NQATdHi6ZWNT1mDWj5bfjIzzBRsklmz1mVKua3O+/1R2K5bEAYPRGNCUqEOUSj
ijkBZ1A/TvCgW5huP74N0ZER7nqpvPOsi1HqVEOV7vX9cwffqvXfAJm/lbokusn9
JqeF0LpNFc3PN4V9rn2lo5TYNC5LOnWp7M53klLYxh+8vjG8HBfnMAZb8bGZ2kgE
diMXM1rtThyd8XswGtfThTbgHZKMt/hkuAWZ0d8974nXro2Xf19VsMFJYiTprO+F
FE36T/Z0gesxZ8FThn3h+TVI4BWoeA7TZBmh4gdJC10QwCHMT4MO3XaATAKnCdMp
mwqtL9HXTDhefO58zEZ1jyH0YKI0E+awt9SraGUA5iiZ+W2j4IEuhe9cynC7v3Fd
U5SzA1HF193Sgg4WoXeUdf/3rlLr+zMtc5mhDuLFLSmw4xDhWkfiJI+d9yEIipTc
C7U3TcGBMPMH3M3DNchR1Q8jNybm7hLmE+pQ8dgCeQepZrz+S3WBT2xy+Lb8eN4X
KGlYuqj7xeLNnZYvcu/OQuRWCjMZdPGsOTB0gspTd9Gqr/7U8O5YATa7RaSUvyFg
BmS8gQjhcuyTTcIIJR8RquEKI4Q7z21VTDMe1QVsCPWP5fW6bfTjdXKECqFjTMkW
Mmavh9ToA5K55PXYuwPlT7pXzacbBG2WN9VCxe4U1Lkj07sJ3/ImPe3oUglmFNnN
w42nI/KGPWs+oBgQYbbJOR41BjU/OLWSSDxUshZIYZj9duzwoMoz2HPg4/q1TOiU
QK4s1p6Vh38COhW3hM/pRKTr83rHKyruLF5dou3VYUo6dUrpqoGA4wyDY7BDMQYf
hH9jsOpgnIHX0kF2wxrTPiXBrrnjeBIspuiwEQeWQTltlhdCGOQxcqWlaKxd/Vdp
KaZ2k3aC3ATW1sLt0+SRKTsvM26vxKfuzsNwKYbIv6KfLcMATuP5rJ74OLrgjhQ/
GyXvoQQb2Ety7Qx2l/oimjp2eca+dd0SjO7YHOaQYLK/4QDbqbV4USdpE3DZ3OZ2
ExvB1eo4wmXWGYfXD6lfjZY0gzR6hV0NrzTWeEL6Kf91OPwVDbaDwxFycsvCeT9H
GwpmlGeWsXyBr35SwaDey+3eGPkqdRyFdZkj1lrx7MzDsMSSCd77jXwCjlQIDSJM
L2xobIFkZxJbYOoXKaJ6whjp9EgQlpFBmH4Kq5jyKzAovRgEZ0Svutfsby71I2kP
CcROBBxC1SpOb8Kt2XwkAgmRRnSURbKdARAnNduzwImsXMYglG3oxjNBry2rFEIl
0EBKU+2pkWqm0CuI3fZOGm0oaUD2sSwX+oHJIzj9PJTGU7rxFye7JJkLXfiiaPwt
Q5GqnAnJODh2Jbq6TKIld9TvyFHOLxXnx4u6xBDP1DWGqBQpjLLwz/G+RhJj1VSt
q9jleUo7ju0a7VWPJPlBpVel03/4A9PJghFUFt5MdqC+k6JX4NvdlYIQvNrbsIQy
E5/snkFXnNooylKW+1h8xf6i2NY3KTRmvfLCy4OoQUqtD/u8OxmcpRlZxxB6cdIN
sIjnN7WnYZ2Ex216GyqoqJVttrGY1abOar9LFXlbkZxhl+hd8CL8q/nMAe5nObER
dd0llYTbAEa4A+ak3fPe6ui2T/iCc0iwrqaRn5hFnqfDsnWI3B594DFH9NUOi9n2
xWTyMzEmaCStL/5X0U0Yr+uBTrBJWQZ/VCJUVpFpu+cJfpcGP2yxlZJ8InFK10tJ
mPKXym97hcW6TBy9MIA/qe6wtfZbd64pVy4DnNX4sspmNMe+UK7Z99eLqniSpQY3
Go3buuVB4XZoEWNPVSdaZN4dM7SzYWQksVwBXjYfTpXyDDtoPzT8m5uVomjqjA1c
q9nMpwIAmvoQcV80ORcuiZdA8yjdcQ0AZoAx+0zGefRiymQtGntpctrgUekqRy+a
Bp7251m6WAT159aNdaFz8NiMt2uqbRx7MymbXH7IgV+pMKKOT0edADIrPOZ2yyXL
z7i2BZqI1DEdfs1+bxojkXZkMpPvz0xxGS04ez1cFgqFqrF7eECv1oHi20klaD/L
M/OEW32HZT1lpEnyXCjWEdoH+qgX9b0SEWNPHLiLOJIVpsc6SaaY8TSeawLNwasX
uBFuU6qTk4z+NOW1YzBdv+DSfQ+JkJUWCLm5slW8x3/+mDSHpz3768mGtWnNVqio
GeMa8SmUR8VwKhB6DpdBUM0b9ID6TveRwKUqH0GiR4r6ZwQ2TnexMqyKOFC002T8
QL1al4ohS57o7GojlPGGF8kZHK/flciJF6rTbz2hhVezs0vbeSw6BX4v4J2/GtaB
6SyavObcLGeYM7GeA6kzxv/2hNFh/uHV5NCNIUPjAqtczQPjdAmJ7uxOcGO9yAKq
XYWeKBUS8HErIbDfxmk6FlpwFtoYY9Pkep8AmitgsB3cPJNiOfCydLcuOfUHfbEn
UDPKiAJvObQjMfCDMMI1z9xivDZwr6i2Hq8WNBWoi0SD4kki5RefXBhMpkagsgmA
Bqg1+lofEeEhW9DQe2sJ9HFgDS4n5lA4MjR2fpcWtPXwhtRdCE7zoZwzM8Q1/eFJ
l/tYi1m0XFdrfZaHBzIqrKSy1tJk0V9/nqVqt6mn+2AwSyX9l/NicfrpY7Tbhldd
eMLtQi737cFp4DoBVUxQYztNPunYt+np1NhmMRX31RykocT3Buv9dfXroHtwAnQF
z2ygdWVPkOrffmNlrYhVK0d4kEOgVE236LNENkZuVFUNaaWSGoTPHSzfLxIjEXhX
hZvUS2DjiaxWJPpphuyIGIAG8Ror58KNQ6b89SA1vD8l6S+27qcukNsQwc4MnXFd
B6T7IHP5r0qNC9AVu+NvCEUqe4IO9SibWoYZru0/6MRvL9nm+vBm6N66KEDD3AO+
8rcet/MfYL2ZLDERcEZZs34hWJeuXg+viIT9S8bIdMaKnguEq11yxuGcTlk3r9T5
3JZJkJ3XPu70Je1Kd8iWokL4MUNKEEmii8AVeO3hU6i49qlDdyG7dbReK1y/dfeP
HIRO4+GLpuDD3/OJyRfvXusL/0eCiBD+FFmHy+BXUGJx2iOC0A+sIbdJe30WItl9
uVjBcp2xZ9fAwLdsSsSjl1ZYglr2KrBlJmbNmI0PAL8pbJH5k0paVSnLNKknP22J
LHfIy06QEQ+CKm3f6tVs3DEPITO1i86v7SqU4cjfe3y36rq6ENfQi+o5OLlI1D/t
iHhu0x9zPsOSsJMcq/hyHSp8N2REKYFGKmIXsFelFeuIVjhFO0C2teb6E3i2SS6S
VF6U0eyVeyoH6HtsAlKQPfaawvkV/9FlC5J7pojSaTX+0K90NTwp1taAgNvMYYMC
eFd6LqRM7BocyziD10Ew+H3F7XAqPbhYjuj3dJu1OkOJ2XJUPZMeiHbNQOsV6NOR
4v5Wk9yNXG1b4VO+6br4JnZsB7vopPwZ8yE5Ep03AS4kiRF26jMABRSOHHVOQLZi
qkUD9uJcKM/s6WQ6vLU9JN2n/NINlIsr/zk2SsF0ndrpAqPB2fOoj7QYebFoB+yV
duRl8U+OsN9GIB/MYM9mt4eB2gvL3WsKybwlxbMpsxVdv7b9CcBAFaDw4nv+aIRj
enitqdO65tdu3KMDmsBCTifotOJyl6NVZJDiC6UNbdozqh63JRD+eue7EkiCj4W8
l/W4iCQNtwhRqALoVtxfKkwxHtRr05j40VVEM4NrlxzZQWldSFtUw8GjM21Gs7nn
4+bw6CLKwMmuh/k0XZDIGwXbNB/6SlxQSD4cM/yndi81taF2HX+NlWG6RTzCBf1k
zHlIH770gg9R/Vs+fJSemQamcrRdSxZfrhwmvqEXoFuyLbmjcJAOL6MSLKXgXI0U
IadxpKbNT8P8Hs1+6Eka1vdrKAlL/mRQ0iW6HnukOsY1SM5IoJQvk+HjAibaqVYB
ww9H9YZ83RMV/U/fUaOoNknPjSVxDqrVMpRs0pTV9UV+4D7tr7cewAAzi9OkQweB
mevgylxVQdtrkcvywQLbLN+tY0yT+VncH1FbZHBzRBIQ/fZSY5ZQ8K201P5pwcWa
qOz+CYu4RXNLdXllc43S1OgbwSAQq17/y9TaIqo1Xda54Zt2E4z8va1Wv4Xeuw8D
ycfK8Ol2wGhOLCkC4HtrHhFmWwV8wqFoCElhlxYwRVwQEPSvvRg9FUqNnZjwYpll
mS804Lf2FHTF7OY1XgQExoNW8wTF2WAzVGD6453BcYELVQeyZqfU+pKGekYq9tK5
bDz+wjsPzG4S20lYTh3NIOaeXHEybI3g0AV5w/2eDGXcFgbhsrXl5um73WYJWKVn
68vLKyvidviIoE72PZba5LuecjcLAcS3JUYcvTeBQrXcgV/+7JQNnxeZpsFklMt7
zOsWRcITOvN/lXAaJNgz6K9UPREoNJx3fmMpKpol5KODz7yN1KARwieRIBGu3fVN
E72uzBoUeA/2lwOAzkSWksIBc6onBejFHSJ1PqC0+kvQ1wgRuBO3irbcJk4Ify8a
ogYxHx5qrxs6RuI3k+pM7MMapNlCRCdv8D+imA+fyAKFCUo8VrOV8l7uc8JnqjNI
faHok7dO8CLq3nRBI+IKjD2adrsgaMYqtmUtRsYbSbx0W7ADtipKoLannu8FJh62
0et34kJIVBv5OVfNDr61k/7jNSEhhb8207m1nouQ1FuW1RGkMaDepyWv7SNRvyCo
50M7UHTyJMobps05498CMlXdruLal7AL1iEEc1j15Bkqa2rvaiJZRpD78QOJJOUQ
ZVtf5FA6DwAK2A4d0X02CPwdAOrp3k545IdHq6Q8IgQwEKJga97DRaY1KZ/MTian
PepUD2ZTRFJBkK3C4vaEeto1U8wrZbBd66pP4gUzdusk9HILQd665oB97Jvesy01
kKcldFoyu8eYZlz67LzdVec7vglGAoEhMqHnnWJ8P4C84GANfNDuW+eogsoxAmTr
YCLLvK5//CasYHLKWSrLcEZE0QV7erQOzgwL2v/XqoZnkPo9EBRB38Adxe5PrlMz
MKY0QtB4H9AczBZBTVfvKgf21uJc0tHGTsET3P4tqCl26ZyL3xv2vy2d6KlSI914
3UAJYIbn1bmT+tyw4efnivzr0x5+eDHSv5L8KfZtqJmXQ1GKUli4dAoRejEOhNJi
nxLMw/zEy4XVjDX2zN6Rc8VeY5cj24K8jqXwCwj8mrjP7cIRGpVxaifAvn/lEyV4
vPJ3uTZO42byR+e3cW07YguDRGBGT6oQKHCg0rZzB2Ew9yeN1uJualS9VKk8IUCM
zx9gJSZK3IbC0EIBLkGOu7ZQK+1qaBgC7szfzWilZiljcWdFxTpeINXJocvy+Z/b
xmyhuQXu08Rm3SfTYaCOxUZQjbErRbfwaTHwhXmexSD28oV/PeQWmm9le4hRZ8GK
+VLV4DlLogJXW2q8UQ7wLAtJ+ZGw+MeKX9zovb3EhdPvXt8Lzrz6AAL9IxgE2FVt
B4LIqAxQOQagbdl+1I6FrNh7o6a0LXQ0XnF4xCNQZBkBGdGsmWRbJTgiVrD8BSY9
1wYHwupwyNhNBvcQ3ne5pkom59XoLByElzYTYIt7wpP33LoWId2bgNG9dj+YWpLx
ndKppBubHRWS7dDDStdIv2cXqnNxVkL0hWOC7ttkWaYuiBjFqSdAx4Kl5Du9zqBu
o60t9EscxGlK13p5w4mTll9m4UXNpC5Fg9anCy3N8jtVDq+Zm6qJzs1Unfa0lOG2
A4l61f7A5fa9Y9kB0ZaJO3mxY+vn/sOB4rMi453GIpYWPMXgBOcxJ1Cck513XS5V
05h/X+gOqjww1/3iyTvXBrj1gycpyVFlhZwGSuY5lfJN3JUBLN/iEHMnjX9+fPS1
AOgOVXUwzhj71eCw7YtVNGeqgzqdWLdDKygHxjr3r2ctoCFQRkTFI6iPWjA7uhLI
DIzrKm60gfGT83FLdpjJECbP9+nobXnYRpoJ1uSVNzg0PQrEJsw9rkZC+Pvmm9MK
RnEuDZlWHGl1kAGttgJnHPq5NnzGBNYIFIzUaami+SaoEpggLfHlmOs3nPSn9VSu
FZQvn6KfJlf9hvGAcIBdD1hnESLafGreXWz2HT2BiZxUCfw9c+31X5FQWuoc48bB
wCsekAGo89E5F/uEVaQeh6mMMdYN4qs9/cQhZeZt+BUuIhZJDjN52baQYE6CBdyd
1Zk8EQZt1m/ed+lZjHe+0mbEo3xBmmYauCBrBAnkMlCVhJpA0OLVK5GanK9ZtfT2
CWK9qsSYvBMHVgLskCH1Vhmo6amkaOejFUjaW8FVeJh8QA07NVg3yWV+cmJQENwP
Stik6FkF9lsbG7QsTrjK67Bmpw1fPw6vK4zOMDBzmUr8UywFpfopcUq5mi+90Gvz
k7OPd8QsCzb9Fhwa3FJZanT3ABbzS+VC07PQGgtT1yKI1ubiUEXsId8fAhhFlyni
QsGBEc7OcXetPbsvnEkFiuKY2sDek6mbJoq3M8h/dY2d66KEg4dGPmbsEFTFMrIY
PyqH9DPeNcKlsZgwI2GZylACdnWJtHpba3+IeJpiUOfB7uOEMsUHWzg4dIhBJGIh
pnOlouv5EL+MqTuM15Gj+Qk9DUSO3HleociwE4mzyEoDjDo/QyGZxtA4u1pd4GG1
3UfGZTsC9b1pM4fEGMytO2Ed9mgA+QKdP43y8f4ZhA7kNBf1E6173Fwh/qZ/ySbv
/BewjB1o/1GE+ceJByPS/a7EOgw3BmP2TUpXPxt4QG/7X2mAu3TpcxKGKfSiveI0
dPJ2cHbibcN0+iY/Gp4CZNOf9M2qOqkTWWE980ISOhOhyXYsM68VlUvRw4b8kn+d
7T6sHmrlIhGKEpbhqdj8sEtSZE/+py84IdX78TAGUsP9nQq1kKT+2PMuGCg/vRMa
3VSczS7EAE5g9YRFpeJXZ+w5ML4ddevomeUncvbgJZHJ9cwO4LWIzEXGdGLNsmc9
pYgwJHHVLJxzaJ/5aI+J7SsGX7PHU9VT4Dv8S8MfqkwO35y8W7aATaLx2JYhxrM7
NBhaqcjDFr/0aD/qk/UHwtG48ljuS69icse5Q42qHAtQf+hAx7UZbwdVz9Yx5Tib
mEWnRI9kqvXIrnq0dRJJ1rpiwBuTXbFjyU49VNc1i6kKZ7vXzk/UdbX18ZlLdNU3
QEaO+1yORd+t3eCh5O9g2iItOfkzCfkOq3HDH24vtRBYX9/3cE+r09bUfBKyO9yE
Xd/fOUjgOU/ab8Uwjsoj9jp+1P1hM9rwcbmc/Ei3LUf8l2Pw5NzAX24/USNwtcJq
5++wLlOT9cb0NIeuvoQFNyEFm6zgSiAkHJoOfxAGNWZ1WlPxv+8XD3lD58S/0Vob
9PSjyWgppXUWcTHzs9nEYQEeawpSwJBDdt02h1q5qJKyiRHPqTO9k5d1dx83ThcU
OueXp0MyHhC4EjTPR9SjuSZyIg7oyNzcrErD2Cr11y/Jsrw6U0UnDbWO2UawNHLo
nTsmq95/l1SrdIiYSQlP09xlo9fPu63VOD8tZfi4Yweh1hZMYxnp/eX0/jDW+xse
KSGIFDR60hFvmMErfYrbQDvhMmDOqf9NcaGYza+1KHv8OHPXxXN+a1ztJi/ahDTR
C07/Q03YPI0w6YgK51YqQbBPPd5g3e+NQxkeatsULXVlK0+ta6LOzm5xg9Zc2lRL
GazYVOFW5y/sbdkCHw1mEsTAOOomwqP3MiKZ9/lObWr+p9JoVIj3rVlBq9AbwxAL
pkgipXTOAS7qhQAd1GqltnnTW5l/JBgo3Cvc2yQIkD13od1/PqcqayHlHd+e9r76
A2WUDP7/oRHl398w4Bf7U8QkJbur/UukV95bEhcuGc2HkDYS15DnTRS0+vmW8wQI
M9xthE8p89okBuJlkOZlGMS2HsChf80C4PJUFyQWxR9H64yAaSdAFe2sI8HQSR5W
tcT2VYpb/+rWx5sik52KJJiyP2ze/fMlI5oA8yHIsO195XtiOyknOHtA0nfY3V3y
/6VSGNigDxMgJ6woNmOhswf4ieU77esIqpfeo5iXRb1psaN/RknseaTnEACzBdYN
9a+zulGKiD9cvwehX7u50MhB7seT2q3s/o88AyI7HJiIfRBLMq8E9oTaMu4wY6ds
6ASObzedilM5Jen3zZkkDgFBAx3OG88YLFHTuSzvUgd6tddvz8UcvVB9BwJZPqIN
R0wA6aa/besSnJOrkz73sJXsg9Xe8nq0D5MJ26iC7g7w8gdmgM3PrrF39kbAtGth
wxUzCuoKgnhw2niifbNgKxKuR/QKX8FCcin5VJtq6p6GUo52zwXZ2Fyc1ecT0q1K
VRn3zzmANZDIrsHMNw4dF0qjCeD9vL+nnOOdlc7Tsd8VVoL7QMaWpvHz2cWxBcOd
1DyF02MRkzWrj55jAsRtie1eJE/qn/ofluirBSgJCD8DD1OIA76c4zbl1AC/sjHh
4GMnwdwbVHK+FLLBDgjQemjsVTlwDbubcPqh2HgGsmh7ZiE2X9naiqA7kFXByaDL
YTJATpKG6L11LK+3aUXpIJI3LNTsuq8bWNQBnldZ+9YZHxpO+zZ8LkjWy4JbFcB8
AH7TfBjbHV5F7cE3DPgHBlA8SlpYMTW0YCHjUWNEg1DM/dsjbbZLvjFZ6+vm0whb
yRe0jw6xC7c9JV9VNDKSIrkhpOkd1C8H8Y4vc5dOs44tKAUwrQVvsGPt6QPhdZao
8+ifKhnnypvpMU/5GZUrTXnDDZ82/BuAJXBzwBLjiyVIUTe/PFWQMkRWSQuhPt13
htzMDSy0HbzbKKT7p4uYfv7/ecifxxrtf6eOtFiKtEAKU4oY+jdP15kAnMLOF5gs
GWl6ghY/eUCGoKxhV3A0Zry3ezYNlWc6DygzXhVkm8GOzG2NoqJq31CUYW03WPJ7
ftPXCDYxyRNdU09xKowDoohA09SiI1V8CCLVJlaX7EdYs3ExloObrJjGMyT4xzmj
yF+oAdqe5v+mqFoCCa2VZbANUxtGro0CWePbO+blGU3HJfTtIRsVxO9zaoVD84t3
d5lC5qljwhjheQ3qZGv0dJfNKMZ9Lpzae6n9O3VjpUfFPJhcUpqrKDWnBO6XTjk2
7iwKnfnEaD489IaPiN0CzxVouhdibHjDNu4HIocp5/vbDJ1GkIbaMEOIJZogoDjp
wu5LxzuUU5KBVFO9aHlKqfy7imblnSn1I9ReDh3yDODPzND+AchesYexvQvQTFa2
eDAokKRAF+Z2S2WDNVZo5dI7Xqwa2IgV4VKcIjCKisfzAQ1FtykpK+AqO8qSG06U
p1Ua6rEct+TbbUWGoTbahqXho7BCtlWiekcWT0vNHe9b+94f3vV6tuF6xxXVT+Gs
v6YAOFpCoB9bJRl79m62Afqlg2eUUuqsBDGiboeC4RH93y9w2rIX28AZh6GcqsJd
dSucODaKYWEA+HteL7aRTkAflW3+WS+hXPir3PUTI+Xk9t48fBL5hW/gMieigsgk
P0v5T3/qJr0f30cpi/1/cBwKAWL9wT/lYyeFXVG+lf74/JZvJcpMlzR8gQhNWwFL
ZVlNQJT8aE1gAPIi84f6192UWvdgNDpSkyVcSELF1EhBajBOGHLkrbRd8s1/iw1P
xGk9TYPVjAhORZLl3T/paTb7vDxzbig2qtR7B6zk+3Yl+hKwPnJ0+Drwu9Jom23Y
f25y5VRIOo/oZAziWwlLOvpUHdJN7EHRGgYwzsAW9TlmpUC/n/AA6F2yoJUsp50f
saRDKFGoHnl7XmGklcebLSpAFtfDGVBN7QALRuIrh1Vs4kTykaWvTCp+Y3yQlNWv
ibY/Ovi063yO7kU4LAkvBqUKEIE28Kgq7K/WpdpCKQvmCqZRHcdn8QTxc+s+PmbB
rFbx5y4I3xO981jfzI8XO2XZWKgk0SZl1aI7YEXC831tsi/n8Nha/cz+IsaACiwA
fVJn3jWFbYIhq5O6333rMiGYlSpPZHqY5hAV5qPMo6pJrFeW6Gu6KcDhqwREUPxN
Xw+TlWRNOyyeRxYQxtCJD0sgASKj1yrGCq/tnSX3cGofGK6WTO2TteFo/TiV4Pnr
kqLuSw9RYEQzbX/0aCYt2CXhCigP+dvpiZWv1ZJOmCiEaNIZqO1wNFOFt4r3zICp
7RSs5pCpj/i5lyLpHF3yRUiHQrgAVQewP+8JZWT7+nCGkk6UVcSV9wbsmRml+Q89
D0fQK4c4J9ILuFbTpt+V1/u3AxwL/J04R+jePBbBi6dClXYtg2qH2YNaEsjKKIV7
5CSsPnFKlCEBD7g0fDA4WfwgOe0equVHrk59gBWd/v19MzZCEugFKfyni9f/amy+
93lIIe9R3kCWN/MtrgWZBhFInVnZweydNElVkca5Ug3Ru2Iw4yRRqBrX0VweV9xA
XFsd7Ys0qEPcouzpyK3N8WL9AFq6gDy7hvu/SevuP/U5nLGdhScbSo6/zqOPJnTq
XDkx4EEGft6ZT3sGJR9ULmKJtu32taud83wvxS01yF4KiJU8eWCZAv+bmo9QX/du
REd5mJNubpMTdgPkMVJBbORHx4k7lKJDDuo52rOkd0Wpf1lHSF1eAu7kEY1OZJLC
dcKz7S3xVs4KQHor0dSOKzBPqYKpZoAO2Smlt+KyBlE+r2yXLgV/6mmoSUVUvqJj
hP3O0A1vc9Qfy+daKNhl2KHfPtvcMySU9YGDV6SbWUT7ZTz9NIc/0gV9Vwjz59l3
JscVGRsrTQfx4jqecN3o0I0e++Pecr6eJjqtNLaCCwpcAXl3sXpRyGJuEqU6bB5W
8q4KmJgbfr9aEdPs1ZQj+m5RXxk66sPb3oovnnFKZAiLgMbW+55sr4zScZ4vaNKG
qE/WU+phhFvVXgvC6Sz3ZFybid9G1cdblmT6QdtSKt7uUIpW0vs+q4DArkqaNw27
Mf88+5UiducR9eV4Xjre++WdfYNiC1ZG8Eu1F4qDlmHQqTu+dKMjJpppVBZkAgO/
dzq92ErQslUIk92svPv1yD8ZzDYsf6oA+XwSVT6QS69uAtLEKhhyhGNGj5VHHB8v
9hn0zbN0wr6S8+akeMSSZaFSasmrXM0JfhmN1urV6kKqkIwNcpnBn2fijROLURMz
daAm5T31+cBuyoUF0Klytvu7th2khlg2WVUKNLvYLnVHyvF3QVFFv4qkmFmJb1CE
2/pJNztke/RZCln8w5GVUWsFYoiI2UrZ0Bd2O8M1mDX2tIftN9i5PKnH7l9jpBFP
dXfYgnrAGF81gq6a60PG8dlEFu8ZWzArQR3BJcx6XvbnJfSkOTx0x0BE+wIQDyc5
ssWB5E5EBOl01BFTvlS4YlvJdxZ9ZJiQAlA1qDIvJOQ/DopITQEt6kHLX+I+lAe2
veFMqxbttEc6B22PTurRu2MpmhHRr3gT3WzUd8zjkRp8Kj/DgN3/DttjWv0KJayv
o/5IzVTNCvk4qI4iNt/nUIJlc+LSGigP5urpvRUL08yHgqL2fx8w1DU+ZWwfXaxV
N9HQeGDLycAf+jaqgQAHHs6MGWRSNcGfcIN90E9T2UqLZPZA0yWAs5lbRgh/OsRq
24B7wDnHLtS5ZcUzpjzR51+oxWW+Xl36G8Lxzp+1CTf2BNm8uMcVA4zeA2BIVvAU
ApDhtwnFMzG5YzcQShiwPrLEg9tMBAvsY5ieiAKpSlbi/4RKFzvncIBXCOv5/gNP
hJiqT+k7pvnm28tGuBbpGKoTrtoeMJSw5b0bGKxpN57f3Ga90AG6E554HY/5jTpT
AoGSstbBjl9irAHGTEYzZzrw9T22o5DgoXfJxmokL1A3yRg4H5lKGdkE8TgIKy1T
09criTZA2FSr2JTIvibifHn00gZj+KCLdKQCMHI5SMgHbRKqBZDEOPCPQ/tuf03w
E+RAaPGWq1B8GRKVdFFNqmEn7OV9wj9YAzKQtit/qHyLxfwkz2ilfYf+gngSLnzl
iPIgjMSBGZn6KV4kTO4OI92X90GoccZxtI4++RPJrzN3FpEJAhRqY47Kgm9MU3oj
2z9NZG1RQPNWEa2EFL8PKSX3cP00/cXXH4WthpcLyDxYV+Twl+4/ZqW8yBR+Gct1
qaIGydzRUDZAaHUrt0LX7eIZetewUd38dsN99bNpU557vgc3RsMYhlhCQFSRo2uw
OngGR6h1eUw3AfDpCXb+t+HFgmLm3K/K4Fnp4puO26ZLtmwlABukoBOCq6fKc0sO
0grJwSBnFhEO6AxtmVgYuaDSJRBY92CgAlrzVkjkqmIksTBFPLYBiJa+CWaxyNuu
5eXIuu4GODJlxTLqRt1hx6BZbDU2I0l5n5zgFNaBv0rp1eGywGoqaIZjMDyUcX0i
zfw01Rg0NR5k5NTU7R3/sLkONKXRooECKEnZ6jyROaEzaEqp89KjQE4sde59YOVP
af8KRb0ctnOtWuZdwXM11tjCTyLVvOuIuCOCgZD3Ztzymc7mwV7KhKYc8+ZJEY1l
0qpBZJW93aWWEVtzPU0b/L+wSuxxdn4YKbkSQ8SQkxy5rTGj1AKqMMQYn1Ar8nUV
B+hoC3Xcjv6GyksqaF6ZS4GO5NEKCYxGoagK3WiuOKnAiZ9CUghT2QlWJVK6a278
D9uvDS5gA7f39ZyBd+X/XlLvVrdgDv5mBnXQRMPdp9TDGMJ3PCvjfe+eviBfkkj8
X4ye5eq6MI6sJ12+OYdhfcGRYQIYhSIBs6cMrYR9ghA0zeDt3/Kce0U0WIwgnVHu
G5lEs1hcm55NI17XT+IHh8Af6Y6bqOuwP02QJ0Ztl9+g10EEclIGTaii7Rk2Jg+Q
NWQ4RqIC7JsPldtvuQjO9U3ynml8esHlm9YVps/E6qqsGcabu+KE6jQyTiQ1p1Q+
cWP/aFqnGpRI2ItKIZdvD0u1yq//p2qEST2aBHPh2sgNIi4TDLlHj1yVFmfwwbkK
V9YG13vM8QoIb3wAmLLcbQqrb5LOHFtMYA0LCXIpSdIqSJZHnzdPybCXkAu/3T5P
0KnXCxrzhKhhqIYGtirfBwP9FXChFtUG7bMjRSQZBYySCfzV1XsMMLJeBbjZOtEN
E2S+DpIYlhJGh9MaIxGa4JZfh2KCl//96IpuFlwkvWdZEhjbrG5w6EYB7PRg/mNf
EaJJslzKymIn9ascfdwbfSOF9CPXNnjqXmZYzI+46Yp6f/+HTmrAT00Y7H37li7l
2n8m0ldoWnuR/Hj+6RBl2fF97IwQ91kUXwYTSJ4+ZHw7r7Lp2xi6jAEOIm9zBbyc
HvDnDveDiJf4IEusuTbJTTwr1iwVxUyodP6ZZ4fRyOVhnyqVjg3A57Z4OwYthQi+
v8qRL5hE3CzdAjT1XaZenGAHqeLJbLf4KMtcEaWF5EKcLe0VuxCxfzjK+xWPFhh/
FKIfrneaN1H6WoQ6TAwSvf1gmZNI/UDQush+gKXkXP8dko+yrXu8KEsQZJfGldgc
c0eEGrrG68AVYXAtqXLrc3ythPxtbQdAUY+6ErU5Ig+2rWSBUZjLZXXweNn0uySn
HXmEIVtvHLLO4CErTh4zI+NKMTzUepEbNgHcs5lICJDRY/5vUnl9EmmO120bUQCy
KzuBlA46gzkdiw5kC19hFnZ72V2I7+nk1NMg22UoDnheaNF5JVKErdK7IBkfefN1
cp1sbOcKo7Ul9rldBfmgwB78Zz7vu3LXh7PyS3YWw2sFSNB0CqLzwGUH8DFbgA2s
7A9nvKDwiPZ2QRTVbJeG+Ry1HPeNIzhpngUJqfyrUaG4KSMtp05lIwUUQp0gc69O
m0NehQXB0W/rIerjOKDqq0AUqeSfGdUFjSqR6UhobaGH/zoDMRzzYGCtqFwqzR2B
hrg7HWP5KOXGokHWnGP0YB/oYki2ynKHMU0jojlfp9ba4npT69nAh4HKtwwVSQzC
0BKeeDgR5Yg28AcOQRMG1HJv+V06b8Hdz7QN+nnSVLKicEqPgZ5ZwkojCVxVJvWG
mYZBmllnwDCVcqO07HLPwUZnbIuWiGFepa97MjpjzirT3jk5VBphtVdVM8ZRRKUO
Pn2DuOa2pJo95zkl25FVlHcjW67l8fl6ry43bKBuhW61Q4mLzfEd+mBxg7dNoABr
V7j3bpC3coN44L6TIdrWEgZzd6lnWoDDbXRnnRDvp2jwBZlQolDZSItFlTveF+VT
rf8lMoMaGE9FvK/fxwH2vdBtE29uEiuCptfO62w3Wr5U3oieuXfRYpsnH/ND1Mp4
p8tH2IJGgNbBkBzJ+NfosJZGs76I+VXMjd2yHcCAcMEYXK+k7TkE/f58cmlDYHuo
QWsO4/ZYo0apOr4B7fTakny3KekFzR6he7n/zzkEoYraUjEYWQ9BYBoH6DGxwtbE
K2wq7wqVxYsknimfwQn+WSPEAna7qKDGMDuBb41Rtwe/ECtosrRQlj86osuCwlM7
wQBhSecI4GGb7SVIf8PKWeBaPwqA2JTU3S/0S6ANqUdtbzlF5XyBb0guY6UvY5Wo
I7B28UPGmhTWXjp/m9rBzRUAU0cS2fXwLctIKBpVPENLhcQZsUOY1ngChvt+JftI
2kxnRXkgYTte8MPuokgHKGLsOnq/6xvmt2SvWcJx8Wz/qjUKYJDDdf38vMTejsKa
8SVGNtm4VxLVianIBIKlhSmaZJFbYxjIeIUm0Qle+kgmWgX+esWuDfyJboPR1dN/
eQMkco76RZbPyXDMC6wB40fOSMttJJjRlCcyAD4ltzuruA3nyyeFQMRJh+/jwieD
uO2CSpq41Q7xtOd19ObWJpt+HHCefPgrc/P9o7ircQ/PRasiOdc+cSY2q0zMBoOf
UxIpDOFpY/WHFWPb9NuA+fFJKNoIhK36PbhfbV7QvV7c5Urh5qVlnkC0zl3dHBRX
7xmNhtfx3+CT2VN7egAn55UHYORWtdRhxUee/x0gmziYrqtc3HspKZ+AQjgNBKRq
liilZUDfXeiJgEHW85JHtF9nZK+4zqLywHHR9PZeMqcuAEa8dCzl4N/CXBis6H5g
ZIvmn2ZDtcOCzyCHx6VIEjrmGKGAZjvWkk1MXxYh2wMgo5dNw61izGKm8zOVUdIV
W2UiBQA+QIh+q5+z+9wAnuanJi6lWfeMO5CouPpdv9vtgDalVx6XjliJRGECLu6h
yHPYnFilmdcLzZipUHqoGm1PD3XPdA0bun3iR/iscbV8d67TcebaMbVnLA7ZoOW1
d/KRjf2sDhmJMWfC4bHGceWgE1mRWnXLb2LLj0QSNhRt04dPKRKZ37/4TQZrb7JR
y5il+SRWzPtcjXetqppWDiLqOs7Nxv5laSX3qUnue6wiM/DJSbiRj5CaCLOrQwiO
DXVE7BRb9IVvz7XyBCYzUowUfbn3BIO5uh2duiy1/641IR+Fyl90zBJfPw/BVK4q
bDWaJNxlCHSiuDa03immr1tnJf77+FcGYzSo8f59EMoT6pqkMImu9n1t0JGfetuH
tN+4gd2mRgMDTHAY7srjps6tY72h/AoUen1V4D+L7tkWyzmEtXdrsRfaE7C98SDC
Yk0hhhl5KV2X/sbGemLrHp3uMGFhV+gVArzJNer3bxI9iqPXNUmcEu7znvCwfI15
ItTZR0/ONWJ9YMZwtW+OtgbA4CbIpWt4PCPILtxv8wpmJwGbHIp4WtqvEGKIN53z
pgchHyWphQ+75jxsOFZR1pO2a7t0pW/YJDpaXbz7zt+CbV5A+SabGCJIkRvwusAn
22nZ5m1Qxfyt6c5citP/S9OCaYU4rAPfz1EAOqe8uHMTVwopOH/bXh7MUaULFJOp
xqfQrjyLZnGz4xjjuJDn+1/ysA1IyBfp72zYXjqXlsPDHz2bIWjk1jVTzdDD/fdd
1Rv/5u4KoPdKjFg+GA5FyaEOrMx7xttgiocHbtXjDiJo9h1u8VUmRGGRrxj2ih9d
7xslO7bVON1AfuBMszMJr0JDzSz4Ix0vE3+ewzWB4FSlJm+dAyDB9b+MPUc5rOIu
IuemCdwsXjryWmlLI0FwVgbSARe2FYzRjZhHTG8qLB6MBVHfCGfQhtA+qoUwRNmN
PXudDf003I/CQ+KfvrNsstgvltHAtTZIRwmO0XPtA+ob2/DS4zbC08F9IpaiPk73
poq5dWztVls7vQT8cnkQZxNnIVc5j077oecFz58CGR2UkfleDgzLXeO5sMgabGAn
jL35qSjz4nQPHNvQ8j1JJf8DbkHNFF5YhEYBnGwWKR6srX/lapyTmQ1Y4bU3UOSA
v2d0Q9J5ANxGKMk3Mc5rLksdPWi0lhOPgpUlpRX4GheFjw3LQTRanpgnqFLMUI0j
CzDnJifpddUp81tuE0jc7aOMqhpMxjxQjHvMoQuNoL6yt4c70EXywLB57vc1Kiux
BFoCoBIruXhjHC/Wj/wnhWuiSVRqSSlI4FdO28UvuO3749Te6jHBh5p0S7I5lDj7
0Gl9n5HZnMy3+QPhLlx1YssLKDli+H6T5pZNYp/VWe8Y0gdG/QL9+1yBPfZ1DxN8
Q0GH23TwyUsFOoQGsvL9a/F8WwEUAl6cv3Gp6gwuThgalx5qTRi7tePVWVhl2alp
r8xB38ql8m+EaJ1Vfg7nbqZ5994+HOgd8XrSBQfwdvoQydF/nmB8a04s/3e/i+mJ
zKCGNlFx1LT9k2eVYk3FWIqdd6tQh3oVYx1UIVCFheixXEIy4Qa1r0s9RLCYj5Wh
9o6qty3z75ctnzcoUlZF29kT8gJUj6EA9OnHkSk7hRbr+lP1ppXSjFrGdSB1Qyna
IicO4yeUG6ZL6nCKmZKBaQTrq2CzxWEV3+Ujr69ahOqxV8hx87dCabE1DGkwKA+Y
CMgEj7jNInUZBXr6aLxwJmXrOOFj+oSpe++WgkMGvd1GoFEZL5afzs/DID4F4i2g
I1zdCawC433tPhUyxu7PnVYx4PPSFYlSL+AH8C4kIbXSfG4Xi8oOz4WhBXfSmPh6
MzqZTdXVz3dAvNlFtxnBvhzd3sH3M/cSa/mgkmAeeVE6TMBzg4Skg6Scq9YuxSaK
lsok/xA9TrgyGIMSoKf3TApHwnqDGzWtvtCJ4pLxaKqypSBzZXSWvZkMnqTuMIRF
VWw/n77dkZPYsN4/ZGbpN/lPoBS8zvWpFBVwr7g2NdsaMGmcHTW/jRTV2KDFR/c+
GMkwyrnGtr7DJvGiYI+IrY/ylqs7hytPrPDC4k2mOzvY03Kieb1OHexh/BXr3HEy
tJRODqGDwkBNk+DQTYtzlsPx70gY0MpKbiZ0xHWppR3xmQ6bxfM0gLKjvwOyUytP
J9PO8wHNTwlaqgQprdJ6LCbMnN6HcqAqRYYpW2OMtwNUcIOufGS+i72OeGjudkZC
f5xIedmQlsF/gAlBQQPL9r1DvOquF9el78cRLsyHiCgdHqc4Zh31LKUVGs9+Js2k
Snmz8nVXQDHE61tzr4YtXTXunygTSMcdsM7uWhGNJht11ZT0Zypmi47bTWrAhV1t
YEHA0qGVu/9aqyLoY+Xbr/xy6rlQWhZQ+JSrWoJdgrpouL8MpM3qltmMqDePgLPT
92Gz6R0LpUyOp87fxaGhA0FEX0kZqO6Q+5W8vJL7DaI0/MT2hevNjz5e0D34hHF1
UUc+Hfsux2x15nRSwP4aRKX/R4u0KojVblno3n+os/A4RgOLKCGWwcgz0vNIsXuT
+w5rbdqOv5hpt+7buMWZoB3/T1O3I4rmolo9WclAfugdivGmbMj5O5CO5TyhIqmy
HM9lenf/phjNLp2xiKrzGgCo3+ltP38J0SWnX0v6x52OtQbfGADmg0vZuI+JdQ+m
q6pr5HdIxpqME/9Xo0mwUu9pE0CUgIAWHsuXFgtoHzeGINQuYrHV0nf/wtWhi3PC
z5mKG52qPm3OcX58O6HhaVH69wkNRdVRwloqe7Iv4YtbDBeid6tG4aZjNCajg75A
XLxxbdUE4V6PcmS52perWnsdaDDl+1H5svG9hr7fw4dBe5km7zUHSv130Xub7mtF
aRcgph9JWgE2QTswttCbAtTebvQH8QfasoPH+zYTHeJU7ujVlqWjWVcEZEiDSi+M
4wSLnMFdS6c+c5fjehmHexnbo6+ADYEwjOWmH0fNyE2qIJslfiMtp4/PkdE4iVyE
QQ1V8el+C6v9xxoYDGS5NJTjQHzysvJpuhhK9cDNHFWecbXJcKVUFCLApbU360D1
mKtYUgY/LNxpX250kLb1ucoQyvjpCMzsJzDNOjiTkJPq5vCBwatXyuNo8EwVpZu5
SUu41Q21MMOf9M5vzPOBiu/+A6Vqrb3OosPLPDvRqXuPC7ITpAdSRLY/fhc9V61K
ZhhLWbmHmXh0Hl3Fk0RomT4SSP37SZKHSq8qTbDh/tgQussiMqsNlHNrSIpfle+0
iG7RYRr9N4pOUlFawk8Q4bXFd2UamZ0BokRfu8qgx38tQ4wO3fbzssPOEla1ZfEv
iIYlIXwRFAlLj/++8YbPyzu7xXvh6wMezogO6SksJ0arT2zlBrrp6ewkuSH2MwIG
hjAg3F2m869QTW5TnoOXGp7m348fg8WltigEXq8m0+CDc033kJrg8pWM0RCGD7YH
OsurxAiOgdhna47v8FY3NjOfe4UU8I6DbRyeKZLQr/tmlRv/0hmqnaCgV2NloJWC
A6Dkb90y5CLukKusDzALKaqA1rNIVjT6gdRrLAYoSJBtAODle9E/URvdqr3Qa13X
qhsvL/CpURRUAnv5KPHJNCJwVcHHgaoz6yOzM6kwLCs9QiCqR3enaxBtmHfDs87w
LE6P+5qHA70gm+6CAXADwUsSgu1wmkW+r46wCLbfgHeUQuyvUuBgIg8QKlhdDja0
192jO4UraFTJaOHQbGI/gv0Hhbdkzv1toJrxsdTcn7jXwcsQSa7tv3AO7OsLerbh
nKrG/2DkuDnlW8jwslQkuQqGhmkSIqHU8UGTNXnXWFJQ5kVgmlxtT+UpulbmOii7
GeLEJbasSOSwAFIF+r9ATejQn7RqVFb9n7/r3ai4XHSgafkB68BpI/Dp1pRL62Bt
klB+82wsdGFBUVSn81MoKzTCQbGICnDljPv+y62XMZpYox78BspOjP57FWpbysEX
snF7T2AHNAA0Px94p4Diq/W4WJhD7YZcEWhjLUSb5V5T8WDXVogMabg0h40fhmVR
Apl3V1v2/KyV4A4dobsas/SvLpiUIU6GRqb8MuiRKk/gcsWemaz1jZTUikLJp47w
ppPOz+eJhhncLqg94SaILhl82Xjyv6cCq/ks7iCOLG4JjnfFPNQn1jlUl8GL1cL9
seKK7V5W7RCuzu4OCjvXqpMZ3clm4qSAgkNB4gOAgEkFEG9+UJGEaYTW1HNETKng
up4IxcUeY0t1WMbZER0hMjG373/RX0RQkPNSJpKHvX5RQkHEzQ1CAbLnY9Jyto8m
nonRt7UER0RGx5WPC+LmIBUnjyJTS2WT3EGOqKeC0Q05ia43WToSGnFlnhz5BoDU
IrGSUxElUoq6xpzPAtbd6g28aAk4V0CLO7NYhgA3yEwgoOqYkITm2lZ6kIPbaWBI
M/xN4vNr1P6ulzQV2bjXyKxUsRbFRw6wVsx9ZfwcbZJxA1FxtG17rcU3Y33mmS+h
zd7FOcYECCvtEERL2fwAqiN5Gxz1EMBEZUJ1yCJxrmYmKcv2lOJwf/ORE6D7m+im
mQOqhMWaalM5D2M+EJoKYiXoQUzpxUy8ULD2z8y5pmp56ZnSvzvM6LNrot9pMxKz
IobUTPNu2k58irGYgNVUszb7/oWfWbsEYJ8dRo6ebh3MOOS/jugtzrpyzzxdD1Zx
ZhUowqkVFoqKc9588i4062xRc86GkM0Pje5RKCwlgqJQHQaRY40cxsyEDIfEf7Dr
882h+VpNKGdz8F/jdTh2HdZsS1oiAI3bH2i67tQbib+egCdPAmou+nlnDrBsJEPW
udKbeIZ4CSsTsu7p90kiJ02+RfxjlOffLKAtw/nl8uu40j7T+CvICXPu4ldFLIQQ
YGDEQbjCC2/ZHcFBJ1PIPBk6lJYqL+EQJP//QOb/0vCCUXxGQTMN5U0VHYTLD0eC
pFMifmXWbQHSuPfLeTq5KjfXWTG8pjJ444biNnsVtyg72sUIcxD8lvKVe1+LUsSE
XMu1sEmsv1rLE0uj0VCyzNToaDBuTOOT8pl+drJ4tRKj1ztg5V3APSfsVLdfKsn7
58mcaNaD7/iwQtDM0NceHlgiXzsDATcb1kmCOgUaTBBvxHk0fk/LHuaqtMEDXaba
B+ZeI55HYvklDwa6KVT5QRad6INs0q7oMd4uObIrhMigpCzzgK+XFy4QI0vLzLtq
h4QsoLS+jpM6MvP27HB429ZfzvESCn9lCflQ6B6ymK2UlijH7gomd04n1hz1aDUR
tlURp5znxU4lEgWUfzCYQu6WwZxl4PMMdoM6X9XUxL3+6LbclcjJc3jMIonnXDmZ
38yEU+oqq3eO0G99r7QseNUjs9sFDN0M5xpLzL9Ib1bSqiHgniafA+hiys7zOcOd
+sp1fcqZ99mGgUbCvfkS/VHcr1qFo9lylT/y6xW4oQPirw917lp90DuWTNI3OTpA
KxI1oDUYybzAXpGTD3mFCBJDoY0x1lm82fhFqqDl9Cnh9ZOcTKxkkQTjptJV7KDE
dGuCwtP6HAlcjVRSRn4Fxg11r5FZ5ebqVB/eHMu32Gp0yBxcm/7vL8MdZPd1Iu13
OtD3qwdWUGvAzdxvvtmAnvwHwt1uRl8TolxY2l1u+1/hv06+L7dzMRKQPuKkhbXs
sHaUrdwsiKRg9yzBi7sx1ybGOPGc/aajd/l9c3HtlrWbWCu/XWeSVaX9FtgHMhWc
/0teK6iKhwyzGq1PeL7WnCSdyfF+yFoBjpF+QrTy8l5DDC2mXLzkAGa1bTE53+xw
jkRfsXmKifIrx4fN5pC3Tdt79363QOuAkllJoVmgKvzPyPdjT40DFNO/7g4laM99
23tAK1x390503cS6DSMH+2UgsMtnCN6LSPBgsafc2TkbqmI1JNCSFrA2iGaVefHK
MYn09xTR/aN7hsoOgnTaK5WK/BEQklSsBnTKBGptIySsAaLwAfRpdLU9UrGBluAy
5BjYDY/bRlQ/6p806JjX5ZoUf0TepdW+YUSlZEtwLY1gu5o1vWfVe3esVBxcaluO
1pGVd9VCeSNMfXuAE4Zf7fnXA5lDPJM+KB1hAaGIWbc6MIEkjK2CKzsi1/vZ0vvm
s/aJcfG1UzNaYM+ZDo8cvqv78s5pN/1wqeCid7zEeQlZoYMJlHSm7z/n8l3JiPIz
U+uiBGcwqcZKOmT8mBHNi5zy5xTXtsUIVNJX+e/N1U2lTP4a/IVb1XqWZKKzP33r
DrcUrzn1CXHrj40dOeEKLLC7ZOAHwmzBzUPpvhGZ8574dlLZYPEMHX0ayRbv6WaR
CrvzDi3AJRULQ02Vlvnm0JtzqZvq77NiA0nJ1cVLezQpSJf83bzzthsQZr34bSLo
ka46MS7CJSxT6bWdK0R4Wz2foSDHhvJ08KMp5atHfSOCXUQ4dBJ0Nw8gSzWyjS44
05Px5xnWAkuYzuO96r6JrqG+M1mtBFuqiHaoCYTiv5TdLZwGtN1Iy+aN4FJY47fP
ByyiyUfM/Tq6//du6EOW+HRMqCMU9Cq4IlaHIo/YNOQcnikqlYlOMOMvc3p2/2t2
rkpIanGOS7cxOl6Gqh+KE5UxFRTOc4vprxPfV85UY4ATvNQe5w8FN65+GSpKTuXX
FhTr9g4417WDCHUP7sAR20EgR/cc4nHC3f+DFXoabGvKqekk+SzLqjVBpl/5+/JI
KPvqrpISDEXAVgF1ucHYTxJVAUulYSUOLgn2eV2labUITWKN9V3jCEkpKZUuDx8t
gro01q0rhSB+g1q5UUORRKIgJ8cJURMi26lgxo6rGC8uc5nYZV7WYH89WvEiWKhw
QB2fPy83Pvg0IKIxqqRnw0saDYgaufIgnsjmjZq340Y3lXFOrBIWVVbdRDi0iqPc
mfppMpeM8S66ABuAWe9C3PWU5/FjsqSfaLtlRM9/Vb6CyWYLGCayc7VZ39nfOhxC
JktRR2PUaB9Y++pfVyx8POXQ1IupaUK7WgMGg4GzczWjPTDGy8Sb56D3ECAJ3ZVM
+97QrRGaG2Nx0I4o21gX/ubTWAlhCy3T1UTbkIfTecV73zbtdzcMsT/Qis0QzSqd
Tz5VI4YHcHc0W25mLoIT7flivtuLLsnZm95J5MnU7bXQ+qZpspEfscsRJ13Gupb6
RdNe4XzW9mJqgAQfNWsf7znv7WHPKOQWNXqzTSIBT2SnnXvK3V1tsInl+8Yt6hjP
2nwd1OaG6fu5Z+IxqoCCuM8LZt4yVuVPsYHra8KUF6L2/D0t/ZMJJnq4F7WcrlrG
zCkCnCtDo6fv8Q1+QGBjX1e+EWdLWDdi4AIbGTqB6C0iSgg+caWMive5+sjofz1D
2j9+sKkIWxiCCzQ95ghkeIzcf3A7y8Zti9hNEPx8zjigZexJLdUwdZeijHjCYzE5
i7vxBbwBQE0VVXoiZAbeDWN7f0KRRrS9YRgIvmhFsHf1m1tzI1AR3LP2dkDUI6ic
49rrIv+0fct2WtJ96YgvM0OzGb5hrERyx+xRqrRol6jRPAtVyw96ouffDmk0QHYg
QP69cm38sGP11/0bhaY27hQio7ibhNZHYDuUrOBBBq+6mfgH6FEg/LFV/xdIdyFQ
pOm1DcjQfXgm9FT7snkaze/VzwUPxjk2KBNB+QsUaVfZLqmYmaNC2Vej0cV8VDSR
aLHdtMGpAOJUnFigjQpkj4R+TJ04Ys6g6oHTA/T49rzeoADRu3wFZsBktV3TjqF5
rAn5UNMoJ5aU4Lz0Qw3/0Eo3bA6ms+xK6+BKeshuzq5ci2Z6y6ho532MsuaRE53u
HS+olKqak9fGI5NqPIZlIp7Wrb3m71fsf37PFX/Rdc9EEO58V8msxBjwqRsZmckg
X98COObexa2yP9qEzJ/WaAF5K8Q/NQHzkvlk2e9cv93s+hOpR8hQiDD7J7xOLhcc
QNwctJMPMn/SJS4IoVaQog==
`pragma protect end_protected
