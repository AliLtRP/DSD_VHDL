// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:13 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
W1Shel4a+u7p0P8zgEAKORExXBNXysORG3djKh9kO9keY/vuqMkKA3nynwpcQcOe
3XDIDfhCjs8Xz5gLJhejdAKu3bSJ1wHX34VfP6kZmRNQANu+rHA86HX2ybG45oVL
xdPs+E5XYWqABKv1Hr86PqAHrOxEFlqp3KOQoj6malQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3104)
gtHK+ZfyPM/S/uVKb7Yo36dnD09tp6wes7p8eHP9HqIAJYneZ/FwjpNUDDoQAeJ+
rQ9PFPr7s8rkV7CbV+RuafR8QlwvFROjE2b4Lb+zO4fPRgeBnjpHtd7uI1NT4mbQ
F5jFXNBcPx48x5ATrjKFgrYujNv2MQIlgMwXPeloeygT/ctHQsK0gSGU9C1jtksv
hWvaLek1iFvK5wC7Uy8YbCmjxupf2kCId59tniJMb/OGSDcW/Yzs6epzTZZTm5X0
xwOYeBMSAIVFUCfggCV+HNRc0IBRm2f8a9pCY9c1L9suNx95t8f2B8YfvME2J6r+
x5qqR9uSeQbzPxE38AUVWOxWrzc1gxSDW73Yn3UL+1xpUk3IZQCJ56AzrPy5RseY
sGJNv/vYJOjDP8Z+1vuMQL0ZfDMEzUOV4VNa3EFZRuCw4Uqx9JogMfQ/uYuR5P9v
4MLn9TvtHyiv4XW8dq4b30j7N8tztudNhMKxp5KiftJQAWOM/LUayTR8YNXMDyOV
u/6GXTRDQt/mL8j4dviQL8Yzia/hb9hztG/81REzUHjEQ+9t60JgeBb8ptzKasev
UOxjo2p28Wk0/ZrkZcWUHbU5OIv7Qa26ehvH1MlWIuJNt4TRsBY/nYqs7JVgdz4C
7VlPVyDodD+BHbxe+pIhwabq9Hsmu10S2QNKobQsr3Eoss78XzrDPbvLvBvi3YXt
zV0WyKtc+mf7UNSTvZeBidMKRi2MrgBoi/HR8lWsNLyTR1PALxP9KbcTo7wdsiKZ
XomJRmUJVUfWFvJlw54kJZGqoIOk+XHi+x6JwFNuTc9f+s+NuRnn2iJ/3tAj3cKe
MRiUTx/krBN3XcriVzEt/cRaXuTCQ/zdT6OOY8/2tR1MLAiFk6Vo+7yuGV4a+c+s
2kZ0GqboweRffK6BRMa336NBPtShJZYx03IsJSz3LOIbXb5KnMMurTDcxnvFw3GE
qQmMqz16eSttA7vI1sUqx7FfNLMBg1EsPYhRXNAcbCZ9KIibIDYBI9hScubKE0/9
efTIDOUI+h0JpmcqKIHiFpE+I8KWsRqg5U/KfJn6yuPbGvQoECE9iXci6fpSZxse
oFo1WafWQIPJOXGBH0ytix7M2JlTjfpSyWP/ElQCwZG4ZfggUqZpWeM36nI/Z9My
VBFutbgSePmmxfDtDy3rvzjFPkCjxJelipFGsvnEXMT6sSVZS+0DeicsazDMQB5g
3Z73kZfMQOzyY6ZDCU8xcfqJ7D+gSZLaxPBwHL7g/v6PeUlUUmcI/sJGg/ozgqPo
gNwg3H0UXv9ao18u2tUN8NYi8h94tsK2kNVxHEo4mpDswoMQ6p0FLBe5rCByccz+
E1ckokPq7wCibtxd9O1HHbW9sD/6pIRK/3K2ZSsw6z5j3SPX+tP3hfWx3n7nZTgW
jE4LWFTzwBWZd5kcXvNkgrFvCacNNhbYca7v6wWD+MyJDDZXAg3ubcSJnhWtbrl1
zPyPoxxCZB+79B6Sr35DAGgjybYBTZl8MSP8tqnqcKeHOJ+Y7cfSQuTuXCap6OJr
3YUzhglSmmLeIpD/NgdWt240XtFS+RNdm4AfWYkwKminLRDBSdUGuYYWZ8zFBcot
SWxHxK7Qr9V3ovsHLFp3V8ZgrPAMjQPio/3i2UJx/Z+WrpxI/ghwu4DPoqDrxzSR
06HkLjIf+RMoe42a9mu5KEBdmwR0ZG0Swv3NL5Rv1gpEAeyNFVqot/YiGvPgRhWU
iDk75uLJYUX6+2QV/JaCGBtJ3gYcUuJkwEwUV+Zan6Pf6cQQR7BcCdoede+DhfxJ
2fVILJ3NXYRtyNHBod3z8a0/YuBze+DFxWc+a6mvYfEfGFJUXyckztXD3lGMR/Ah
hIv5a/oVnu8k+Bwn+GWy5X9vAEv5HJiC7x2eJ0pF7WKDAN5tNZaxuC4MbQ3axAFG
Ypd2f+B0K2k+eqNLvHdi8G8AHZfj4NFkArPABW1oTY+4DFa/HnFmfKK5NO8gVqkv
3t3AMOQTbEI89/FQwPGcC2BfjlGD8j9Lui+wImQjwmofE96pCD5mqtXijZ2Cptl9
m/Bjj6Ce1MXB4reVwhBYQ2WjVJ4R/WRe7etnvcG0DwG1fNYFa3iD6Jd6Iq2pHimP
0ISgrS4QcWbj8V4Jk8RYVfljKTecHmDLPNYC9o5CbVFxOyW0bSPQMbqeRQxsyV2r
vTNSEODrViE/DPsCdk9x9fmUgDlMp3LaUTOIrFB47RYv+Tx5gLBQl8A80C7+fK41
sXFj8wqwQlRp+gncdMBnMza2i4upCh/MHWE8kycAo1zzMgY2i5umaEPV6CmP+a4j
1d4uor90Ax7wynKMYBQOCb4TCCbwEXMTmkZ0OTIjn0HkiDouTX4qr3T92lZPzJXT
Opo/h5Y6i5o3eTgssTeOzXuuLuKmWvhR45X8bSIay9cjmrz0Ce5G/3CJDzTkA8we
lNDBp+vf1ZpbXRhDoJXhdwe2Kk6CPpSkM0LVMQAvwC3+DmtowafpEE/Y2nmgTx+Z
bbbCnhm79BKF38RiEetHq+mZdgIRO3887VGt42EC2DHKh1IsriRor+9r7za9XlL5
5wZxN8BACb7AVbp6tCld0T6Mo1d1pFCJVsqZVyIcm+2ECqg7O7xZis7wFeKRLdaA
fyUzDLPO+BT4joFkysWSffc8I5YZLCJ3+9iqnIQ25nPpeKENP5nA3V/09y9oBwJZ
nyllWsyZ9TZFcSo7lk6cQHAZznhgy/mr58jMj3ng3sagTVYmku6CAOW/WVKcdxSY
i65S1abU0XmwFXSk89y9pcwC3sOWplG8VpNhAroug7c09TBQRJzPjjXfsyfIr78a
6/YnjdVLAq9Bl3qcbklnKO/PhWAqaj9Mz6GxI8pgJH5+HCYZpdGJJp9sPV02vXwt
kfjBz9HhSelhPXu9/+HYHoYAmyDwCb9/Vp2BB8l8jx0FXr7O96W95VpoqHTqKl8q
Dc/EFW0aE0QLxY0+cTYl6JlRO/sddMANmXnPOiIwACHfVMdZ56espFvNICxj5IeT
C3dLKCf12IIjL564KL95W1c4V9iJ03bu6sdsRewcxXkt6WmdjCyZj7vwooVmjXTL
+GlHMUA2nBr3YEPN2QUBaGaXN5qoh+KZ9E13qNiOmUU1oaUFI4QcB6iy6uOomrA2
X3hqHswQvcxhsoOEdf/mSf7TWZe/mzIRKtCsPHKYSEQ8BPpHAxvWVowcNiT4ItSB
ySI+qFG+qOcRir2RBM2jcT8OjbnbYOFRqg37U0xr6Sdcwjk58o2W6MghIUvIbJRl
1nlMjAVlb2c0jgfeRRrQc5lRQy6/hUR70/dDts934QVypKORk57wEKMYXdyzr3Z3
Qfy36Zev44+DCoD6y6sAKDh9FIpFmJaa9Y2wsqKUOei4zp+JQ41PYq5Tn64j3Ie8
CPgKmlbsN0CYqTBEo2kDoxvra/GQPepUHi2C+gIDg+J0ZjB+bRuz2EcMQgXE+mzi
TUNDODrIE7Z3n4iQx47OBzlLEVMnAgcGoUeHIrMwUBlLKSjafQjvyYoknpvi1Q09
CYY6HhctgDRVI3kEtKIwjAhgykD0m1jrhUxTUEPaO8hqhuHdRnVrCygRiApYgNoI
oXyjvcxKycP8XGwdn8h7ILqy3A9AFDkQpxm+A5Qa5MaFDpimm5mRJryxN29pd2rp
nN8inkRG+TYV6AFgvcMrob9VgYYQjnI/IpbhedjoQm2G1Edffg+Ct0YLyC3oAvtl
ADnFufyVY+VtsxEdIg8u7kY97r3FElj/lu9hTiB+Znup6CDM9rmFhhKElIkwmTXP
u5RjNQ6P5Bjz2gZ4KCxkFxLMGn0/jnN8eMGgmxkCxI80WrFACHSQmsW1/HkbbZkK
UpIM59BaaRi/43a/ImAtJn6ywm0BM5szuepHztRN5c5NcWPKwXvgRbUBCkUZD6NZ
x9i7YiRKWUEuMS3KWB6yDcyL1Kq22FMP7UogyiSwPA0x0YA4ob+Lh0DlAPHCh+R+
FPvQbUEqG91ibN/Dx00Ge+nLWvlsHSWvgfYDGl6xwXvfGNFXletQz0zO2ngQIF6H
USIHt6QjeWpk+9WUtQyJLm38ksrVVIJDvcSmEvzTCuVe2Dc7fB951Gm1JYto5ZuS
XnqJXVwxtfRWlTisdiF81uIt7ZZYvw+L1mKmnt7WysY=
`pragma protect end_protected
