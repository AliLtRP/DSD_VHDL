// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BpDbkhZuG5E8uhCt0LwC3kNJ5FX7h1j7Chz4WLs9oLIqBOVEa5cexsguMM1LaCUO
2k3CAw7dvHhYBPMd6KzFBMPNIMeXrMFFR1c7E1LwXUeVNSsCUKXu76Dzvqn/Mxac
VsktKwUHAUzPQUn8GB6R6Erhy7XhftYgHezeDO4XqFo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5808)
n5Z4G4PDrE0bg6P6Ey59Qe3dF3wqxS/sh55zoV2chIsadJRxU6ty/X56sao2Dmzy
wsGq60jjkQmEOHaPbIsYM8csWmCTk6R1BKU9Xh6cEt9RpAXaQrV1g1B7p94zrM8H
hku8QEQeDjPvZDVYQJgKmZEcE2sE3ZjPIG2PvIH0XxdAbbLS6j8gNz3+WL0X3VJt
wnJAs7vlGy8POY+6UACwE7d4Nr+FeU97nXtQGnM99BnftP7O8ukJN4jXNg0WDs/r
EiurlJXI2L7gR12NodcRazKNMz4VEWG0byU3xh1miEWpfZFZaelkfBCH/wtSibpD
i/LrrTkBuCugw3oDN8n4qk6XJ9wW+TDRtDP8aG58tA/sfOKkjKY27YFoehdQo54Y
49mvMP4/exL0bJYHwn5EPTX7QF6FwkAW3/Ndb8d3UO7cQSbMTwKntUp8g+B749Mu
pzJqoCvcTgLMaSRPsEu2+gdVt1Rjo/7PLHZNC3dl0goU72mqGFP38gfwezU24WZ+
v4HmbUCl3vmqSzgqw+khF3SqG9y9H84d4yrVrN4Dn2rKxrXHB3X3Xv/DpPgnbBzK
2HiZ0zjHDEv+d9Ts5nILguqwyufLH/oOnxkl1KHGs0t5BWgIt84oea1Z+xmD9ANA
y99kZMexe0v/yEhxvtRRw02EWxZAr0z555qMBf+S0nP6WOlNxkNLtsx/COtLNZHE
pRPxg/gzmgn7bRvG8CNAnCv0JQxP0o/mdYTluZfQf+Oyz2mcP6Cp2YLFvo6BbD13
OSFwdhbqGrLV/x4aqDR1LDNE+GU3KDt+cVKC8IQY9O+HmGPfq9lq5d0N/bUM83kw
DD2HbjjIMNxTPqIwi6kvP/QyjNf1oGYMqG4poBun2K19dGJOEXCi5TwWIDooooyI
SxsaNR0uItA+MRFEKbqletjVJ8+cElwKn9+pWtd4VdXz1Jy72wg1h+rfAVV6/jum
2ZRwybRcbgFOrLSE8DBc476T7oxnua7hyk1waQ5sw3+BkrNNQM8kcLvrNs1n6dWI
//TDYb/6f4lkmswMzBYTsUQRKCBRcLGzsR/erQawxB3i2bMVWGY7AKP7YnXbOj7r
g/CJmRMcFexIq0p6y81huRHX5/H01iIUPi5yqrx5hIgtdnEs3V8CrKZNtghOkDe6
uuKUOO77gwn6TfeOkjTJu6YeZodAvdlKxgsgEDs5J7ZqL7Im+Bn67JInuNwmttmV
qgA8lFH/Pila3c59bmXqf+l1oJp5uf9tEVcFMBjIxqwpWqdSPIhiCdvLW9L/JdH6
lNgCFV9DFG55ox2kGp9NLtBFmCT/K73kVNL7FJNxGc5pnKdkttl8F4t/l/lnJqtQ
CrzXckl8Q5OZs8LfXp+4LByEIHYAZHEtRo/sAOcQ4I4SSatWeMizKNY43qgyWB/t
K8A6QwyMmAwN07btbxeNYHSSs0HHEM3OsBfJBhKeqYcgtC+8nnNiOvqfd8Wk28WA
YonfZc2jZvDupOXX/CYiaINTfCwlip7cOLjo5pqz38oiPiyhou9uqHWm6/PqD05h
0nzejQEuq5hSZLd/tgoDCu98WQL5r4lC0gBRGyGsUdoROALODp884UnjGM9ij/u1
nGTpmW0go07oevgZIgA42Iaf24UTnznujp0wEYnvoWumGVwk9Y89u3wa19RSQyEL
ZZGedq9h2Sq5hUXdIf7aoylZ4pjo+8vOY9mUTyu0LZ0PiPKVdjR6bA2qmW7kkkbc
+hsqNnTOvWsbKP39RokfyrNUaXy2IEdt7k0sVDWHdLq2mChfcnWqCVJzUxc8jDIh
aBcvuSNGHle6nGuxktjXiLHs5DssR5rnIZOkQKs9d3RhUwlGxVXsDK58cyjQ/LR9
IeA200f5WiC4f/ygdXVds523zN++gsFBAf4P/qEsqM5a2bIzXRJ/NPhDJ1SZUzH0
flEdGdXbF0aAtPWdSp4F0D1IgV2hdo6iItl2sXWbFul7wHV2GfnpSusrDuHPOgkn
nQk1HbpSbuYKbYh0R3ZAEhWDR9ASDihLSCiBtAmnmOHmrxIis0MuqtKHnNQeqP53
hD50imAB9hntTF91EYh7TQzJOFd1REO/UhP4v9nLm/uRPSkkEKhwUYmzCkK3975B
JCYtH7u4DsUFY9WV8c1SmLaihjARpOGwHHSJ+Hiko9YTiaUbLWS+WEGiCY3VzGBv
5gHZcRVWzAVXy67luKd20WbfSzp8VxtyZYv2LE/jN782gI7OmDNdQsSPiAt/fxDV
nuRXkwRLUWiNKNGybryV254tG639E0ZfnTrLsEKDfuw6IXQCmFuLMFhpksXixpSU
5SPEJtN7NOyDLfvIE5vob7R+t/3FytP3ujlY2mbdFkbT6Pe9iQN7AhUqRssO4GDD
Ba+EoRZeRb6eCsgvH4l4+XZXPHCGUlJzAPIc39m59Vy/UgwNub/+yWNKsPrguXpZ
vIpaFlOmPot3det6ErL6lbzdzarA4Wol6In2ajZV+iPbodcQIzIZ+rTdANwhi67x
SVb6HzmGKBIfoRVbAOdkRCAcySn1DnRi5ruw3Qji1K/9RX1v7ubsRtaq1YQ4RCyp
MJ7rbUqWteGS6jM3PHB/mP5wYPkToyV/5vbuExJDdICGqu4+9R1QHKaPsS0DBUz2
dR+eAniKkcdVZQ2u2CefLORFbMlqth65Gs8FKnSDJ0iQMMwqzzkjNzcNQCTbEPJ7
7ZvhAidNvESLO7BlH7cQD0u7lrPNRXRQaS6QZeOHVtTR9KigOIcsJR7StQOQlgWK
fleyGnXmQZ6JQI/cn5RsQMcZUaohOWIFs4AdSamsAKQlxL4NCrXtPJPTUDzZyF9N
AcVcYHmE+zKZr4mBd1oCELbKBidEn5is/6jx9N/NpyAN3v/y8qNrVZ3mxJ4L/pb4
YNl1Njbk8t/+ZkfpMzaGPNd1AOE+Kov6Rk/0YfSIZmewzL/P4wqWcjSbLLMPiDEP
xS4xvetDlJfKet1xdacy9dBvfmDpQjpSYadD3bZxycbAehEo8XROJSVE7kYsUEYh
TZDB+/OdUHHcdVJdxaMRALxaUS+KHF6mnH7FLwmn0OxwB0UFI2DiVyZbGJCJpqzL
mxLhcW11VK/IYcA5+cP/wQK82hSqkWVN2dKqpAkwD0DPfSbfcqXXyaKWWpAZ9fy1
KVRMcXFykibfKoopLMMQN/uhil+iQWz1wlknWGDlh+gFhjC7fdSDnj+8HUQ7WTo1
BhfFXkC6v1gnvqcVXXPMZPgcwmxMZpZqvQcmnGh8HrEXPJXb24JoYiaIxBLkqH0B
RLqfJI4GCRQWcxUr1PQuPs0ImyxA9Aa7tT3icUZ7vTY79VT7t1SsRoTsAJvDaNix
W/gaGf/lrsqJmdM9w7M1zNvKTf7ZvpB7dfcT1m21HOe7ewv3JoTmsCgqP00dwsGt
eseZgU9X8NKaUI9vwZR57SdVCwGxIKn4tPYzPXUW4ikPOdE8U3v4AUTCr6JFja4I
1o4U5y4MXbP5g5bYuOeX1f/e8fdwGoOXayt8cou94hVjR3nEoUOcSduLKgYHpoNG
A+Sn/GLxX7XxIy/JFOh1PSJ5vSxzYjwTEKEs1OA3ZUXRk2Tm1FjRPI/gf5YCT2PX
HSdaO9z3HFEdq4Z8myLlrM5vwTgCsIvlsnASVjM1gh3wauJTyT0NN6f0yNMqiJXN
CIM6VblHVJgnBIYSiziSQH3TNT5p1TDE9ggSq3pJ6TQk5QwbaYzYDXZ9p13YLu54
kmYC0+x2oN6L3jqcX/cQHoZLTmMqlqhp7uCanAcwF2TfmspjWastN/5pgQP2zhVY
UYIy9NXa3exWYzlkGtrCHjmxImP93ruA3/lMqbEazNni21pkgumA3ybvjGeO2fGy
p1+gnbs0QSdFkXrhrUPQOKkF0ravmS7IdG5sA2FaHfoz8eYW2dT8CkJgm9UVO7bZ
qNEe57e8EOa6caEJ+8Ie/FptATvGWINe1JbvJAP/64XbqQWvnq1iOGsHLJwd5feY
w+n9wdiXLBwI0E9K0I28kZjOEwZWPovuMe5HiHoNZCRnlpdIAcZDkDQ7EMj4GOZO
F+IHYrHZYo7M/6IBb/T3wdI0JZVO/bBIcha612DBgiBXNM/xsBwcozMQ8jyYCKKF
Umm5TO7PNRj7awR3i7D30QcmbalzuoT0dOzj1vzPb+Bdh4236S5zmqlqqw53Vxat
U/U+EhjXx6xh5C1NrnH4qU170mAD1gBnoyMCFFXJEuILYvXuf7gKhUjflHtQE32x
mGY0ldk57jMFVaVtZgUmez40fbo1Pxj5/eRLgahNJ6yFWlH8zs3lgQrUtWALs5AZ
Q2sq5bY98opCMcbiuU4c8/ZhL7fhijpxgEk8Ls57OOuVdL9/Dungs9Y8ZQfyQxlx
OL5C4Ona+eyUpD6uAw0RF64fnRuOD/vQ2DzA4grs66xYi8+lhgY6YKkEYO8J7P/D
LNcYJstT3XQ4zXSGViec314Bqaodqc/DuxTqJt0pmIORX8UAOc13l7r0/LTs0ETx
6pxTQQ4laGBEM/cIXfKNG+ylDpCT+cm6hRMiXl6OAT/3s4LGul2LJNjtOTMIlLQ0
khGihsiyYS8TzPi7w2/EXkXVSMRzN+ptGn9+BjF9e7/FV5+mQoYDcHZG0RhnH9SR
E0mIujCKjbKfJ0AVrYY6KGxEoWFLVI5QaWVHdms9kDl3h+fWL29uMqw4K3mPW/NY
6e5iBGXwEhyGnC8zYLMt9/NJ4ZEtPeK/flZzRNWGNh/tP/segg4BiSBudyEHULCs
CITaqFaUz5FFFG6umdhZYPeDxkCzIVV/mzsBfTQV8aQoUSJjSJ3XlD+Gh2BzcedP
CXoucJrIA6blw+iVwYz29pWXsfyqfDQFtCHOKyrdgGl4pWUVL8b2oepVNJ2BlHi+
lgZXYTE18M+U/t4a0QNUxiV3JbGf5yFhzMhbTA/8DTPu0B5wnNj7OoRC5fa+WQYG
+4SxZ7lexO0S5ytlrgdI/LXE7bwV8Efg/J6/9TGZ9qm1j+0v9M5yYnIrQPZ1eTB0
X10Za1N0rMCT/Zb7zQcuUL/mvzsvX5WOtil0Ji6qONTVQiNhvQJO2Igl2Wbhj9+J
wUoBXhBdoQPndnocOTp0XYHoTbDOgfDKpnU0e4TY1YKueTaLEiNECn0X8nC+nTj4
HN5Vb5m4jrovKdn/56Ou7XSaokDUZyRGwrG/ac7+MeqZW3Yi5hk8kN9XnXGWDB/e
onyax7Vv920+GPpWYj2EB6dSJ9X2kDpqVeCeM1oUr6j8W98/rXq1BggOL7gl81JS
GJkihHNqH0bEtM06Ypha+KsVSNOOajy25RiESqsk/31gSQO1hrwNuoeM8A2UJsyY
GCvq92Unclqr3t7Gj2j4l+H65u+/ArB4C4jXusioDqvAhoYNcywQbaGrnnRBk4rO
5dpkp6C5CjQBgTkOq5MVwHb4rf9lB1Ntb3tMlFe0HIstV89HD3xrSO5brC0KbiI0
6Jz3Qo0cQXtCDJm6UD43LtWHMcK9p0m+W/qWCwZiwAKkT1+41DfSeqI4fArqsDNY
sRKwSO6Ffp4Ehf49Bb7QEncWVefSu3q6oeIyTAJr+hNb+SLs3F5uOjcf6e8vzoil
W/UMqyKuDhqH+f/DGKlsjWrQumZiNqjrlswkaZW9h+nMn2GP2owghe3tQ4aMX3Ex
Un678rueSpuMgwZDLzwH5tUrbe12BVLNm/Py8lsds6qJhkrb+lqZMWJK8vOsKyhi
sY+XrurxAaPJgXfXYgB5VoA8tdAspxTaTBxpcK25QyT/DT+4VRE0sWk9OABChfG2
4YDr6tr/XABKOqYex8FH3CUA2rx/4SWuvHXimP/UImINCJCt20ABo34SXAzXMGaY
/6vcqmwQA0aaPsCLvgxXdnstLlod5ZhUfEaAqWF52GE9TsZ+KvWtdx/iOwCzl3QL
wGmlnucLUKZJeq6lfKcZW3N+kXjnJowg5hSQX02EZy9iw4VzBUkTwnO56QGXjMq+
62jClNAAFMpHlizJENfp+2hSN6Cz8VyA0VfyKOpQiO+KIsr6zBNI39WTsLkbVLs3
r+vK1nghUIEv0ugPncL1DsXfT6uEjMwwgHlpsIhq1NoeqCfMgmxGQ+Hj5XREOko/
iuzrnvKM7oZf8SEgO1sBSiOf8mYPVO4Z3wHM1QuNd4NoPOmHizGkwr+ir1dLmBq9
vUJ4h/MRL7t/PBhJCQlVmKEhdJq1hZlCIVL1JQV8q/nrbQVRMd9MBnBAhTPTbfEw
r3Gg9D4Fz7XuP/tS0Wna8KAmGhxjPOQtR/DJAf3li0BtVSodLevtDlX43Sn4rmG+
gqwdHOQGl9alWO4RDEYOZuHEOC5qrXCrLbpQmzoGxfo0a7gmyHBHRl5Sggjjo/Ec
ogPegXJpfzwNiDaHjtYmzQbpWAYCw2sFclWpgPtVT0W6ifJVGrpIg/hHKNPdUI1B
He6kD5zIAtjd1HWdkqzmomPtUsKFWTuJTmc2fkg3OCxWpWk6dSz3HxR8w4O4AoPJ
n22p7vo/UMAI8VjgYxFepjRRUvQn4xhK4UFhfKS3/OdN+qsjdU85STRZ31D5UwNt
8w+EuvUZoW1z4stnzBeqGL1mtTFQhZKYLl5LSC2pHpa3B8/Skr4UVP2JUXaRxL48
Vo90uyPXfMGG5IfJloqdPqA9U7N7m9Ha0ZtJpGoM9q7i97OKCYWUVbxD+/SxMVKP
IHsvOC/RGtMfa7OvvjkpLu4wC+GjX9pnBcZcmBiOPAtdFxYcmYu/Yd4xaPX0vpji
m3KaoXIR7l++DurYPdVd+Zi0NAEtJJWrNBPNmv/v6rUvZbgAVbZh3aG1MjNu88E5
VlVQAlhRrZt8/E8XxmR0qc79ciZ9DBIyOP4tNbW47BJC+G4oJzDXpZEDTs1+fWNb
GiNEWB/vK5/6ZQZzaL5slo9qKfsaZxmJRPRyz74GgiGLQmUJk8dMEaDa8aj+64oo
Mu8SQK+KZ4415ZhJGwGZKjFSwoY8jlmxlcs3hsvN/fD6ZePDwr7/rjJs0N5nnMhv
oEFVdaj0JHT3sgn3FglUold77cdrjSkeD7P18adS+QouOse6a8vOyTXENmFLMBqN
cBck7axZPhLy23WnbKdIQxG1KhWsc0O59/SSi/rSqH4KCkv2bOr7IIsaYGAZ5Sfh
RwHFbtPoDpdwlFPJ1jo7H44+bLJ5kQXHHPxMyP+RS17JSV/4tJfgPe+aRdvPB4sL
xIrkc0be8aOEgV1S1A/Dz0nZU0THvqHzQwrWVbiNwFkyCK3whc4Ev0lnKtuncxej
PMAZX5zu/mDhkQJB/luEYV/VsM1I6lPK+JlEaf43dCUnjk8glGj0JOcJFNeK1XFX
6w+jb9ScwMkrsbNbq6JCNoIHzGT3xy7GCrMC10N8oJixzljev1Vr3nF4f4C1YLXt
fBMMCTV6FXrrGHV494JOgYJFMPDpjAo54CLJ9EteeogjphPQlHpmw1b/hDeRpdB9
0wRNexmzZH5oKIJR9XieiPX5D8dNp2EwG/CSiLioegL/uO6iFbKS7w9cBfuojHUr
96XkJ2cczOfsYKvfp6EpHUs3qoYUgkCqrjXb0i+qEPtkLBR85fqyOSWSrhD+/z7O
3Ob0/vVsoJh0O5w7Wd+LLx/Ed4ZbGp93pjx8mtWzZdn34cxb1Nmd7rdIU84fZkd+
MMzqhRBcdA4QVl65YhubsOzmqLQu39iUEDzzgDq3CusX/vomhc56ZxOd7YyztlIf
34AWdr+lzZ5wIYIgNbX/R5y7OBH8vYsNLwyIvPdNSVr/g3ld/RotbZg7tS+jMZAX
`pragma protect end_protected
