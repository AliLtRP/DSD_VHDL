// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:45 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nbSFoRL/8Avsu+oYieQjT2IUpzT7O5A4oPm/6p818zl0RzQQUCyRY/7LhGn89Zzk
EGZg4Ib3F5TSCF9n+WOCsUDEqj4yePDgQ3H53XDKPHIlFWV9mseGV9V/QL3WPf5E
7/coNZMC1ctfatEHUyipu8A/CseueL1LjwXiry7Zw04=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6912)
HGqzJqjfqSePBSzebYWfiBbxLAP421ESX7yYQg8oAS3rJHDOknhaCtTWrb94suU5
GAz1Lc0/8NEf9vmsgU+35WUiRKy3Qq90RuL5FyaOtE82tVgvgQGaZmSIwqjqm5i5
HHFjNBd7j9es88nT/m5+aEx2DHxpUT5tQXOdOOLBDT/VG2JRgM8SwehN0kLWn2Ui
+rFe0jPrWT4SFJmB7Mei5LdW8rqgG4y42vnlGNKD1p7B3/a26xiLOgI56fFfs0QH
oQtHZfik5x4VoL01ovGKgZ1SoxsUKia/QxZfRBBnRvGtuLZj/GH6EBcmJ1c6wHd0
2ohWR8aOAUwUlrnf+EaxuEn05RaOurkqc8J67BF7ObTFgChtnorjt/4xVmos0FvF
/BHmQ3LsvTmP8UytnQu+J162Cq0IH37ShYLWjhbQHRh2hk/4Ecf+qWRRXpNbvuD0
aMtPOdd22rcIHgB/fldyKKAbvY7LvYTu8fL+/ZkVGyNjpdihAggTvifcjNpH+7P7
sTXsnBz5a8fcIVdW912FHMvHsKRybKZLVXQ3L6d6u/cJCxrQQQRoRiSfIF+U/bi4
Qbbfigrlc9mtiDwd8v9YsQLW3JS0/Mo7XDQgDkyT66wRVp+jHzgYwI6y0acRUkw7
roR1/jNE0lC2lWWWy0+rFI7PkWpN6O++fPIzuignopv+iPfKLwOmNBO252acRnJw
doFHFS5cB7eMyJhmO6Giwi6/2DRwtN+8zhmrj3iCGsz4s6PMBmesUYxP93pSMl4M
8DPw8HQTeABYWfbk8ouK98fSsXJjpaQj6VKSyLngAd++UywsXdC8DCm0y555xqIm
+azllOrCeNvoFETOL1yu3bhf6XUm2Y3dSwmRCmD7MW8qJy5cb4AwiiU00ItgO6wV
PHrunUkzxMvTUYpEc2cEeWh4KddcS85BPYmeiAiUn2w1UPS2ylb/KVJhNZURB4nq
WmjuFMUkOdz/Bk6zqGh1pZVzfhlExlcEcoFvkkrpr/cmiUYHrWYRd9UeRVnWYuK4
+7qElAmaVKLE0d5dzIXlB9bI1vZ08I37fO9rrTBLM0FGJNTfSH8RFNUiFsc71CfE
NrzewUxfGq7BujRHOXOEq+h3lmXsRtSiczoWhCFbYzFjAfWn5yi3s1eZ3K0axmti
h8V1/n28GtfmYvWvdUtarOfu4WeEvi7Bh7HuemyMt7HlUnW3sc8xwuNx4zsh3cYs
98afblmli/QxINVCvLVIqFQu18i3nAtqKbVL++6BbzOtA/Kpcf6oaEIiti9PmZWj
qwSwnA6M1FgEtFIUEv8BcPf5iuu34wYbZQ6g0OnihLTPX9OvGeMpCb0s26iIT4YM
hfZe4HR7lfr9V+KOti00soNMVR8g233iR+oscPBREHZTsL+Y2+w6U4kqvd2SRgbJ
VATgGT3EiBLKBqAyxHNa3NJnUnVGuJwfvpSJwBfr1rkReTy1hqnQUJIySBoWW6pA
1Ohf/Oc7qIUfdkxVmcgJpPDNRnZ0tA0bEM1WsBJp2ObXnYq84YcoL0bGQvHUv87u
5841Q6WLIUoIUT8QfYGEw9blKhyjQJIPpqy48zLIvEVTss2MP52bebIRH8QbDC51
gIMNumzDErWDm3TF0eTrljbOChxor6XGEeWHr4qDSfvnIEuVOX/5F5Sc8fQPb4V2
AXqtacIg2C2eJyA31gFbKSJ0WuD0izo5VvFkDyK/h6p9rEKbb8QHg1AaflIznV0L
gwKIgtUnz+GU+961kujxdqvzqFJmtF57ndwKafZzk+OAzsTMLrW9oq8hnWmMI5P2
Qpym58/BMV5Bg3dQOo9m9xp9+g0JqIk7yijGpXMG6T3QBw7Tk7xm7IDNNrHPrXxS
f9ZbMqB0BnWYk1llQeBD1zBdWRzXQUqRN1Os/HdATpwZG8tpw9+XdGMM1aUzCQHf
U0SiQQuxXBOWQe5DRkrPnlZ0TAQz5AjN5CGS1KmsB5mqnakk1QRvO8pxG44CheZt
H17Fu6o3jFoqah4ouEWxsaqL3jDtg7hK7bCo7LpoDPPgXHTqO24Rz9SoeJ3MyeyE
1ydKwr8hl+v5qLt4Zta0REDFn38Hd2wKbjgquo0/+urRUsocLUHoXKNc01sFWEjj
ybUtAGGMJz4NU4MMmh9my3ch4vdtFc5jOsEK5nQOuHdZ/en8P8l7ETe+uHbZZVS6
Hg9Hx7fyUbBpTUSCQ6deTYL4LSbwXm9XDCqUn2ASLd9Z/FfmVbCVbuZLb51ppFF8
X27kUOrkoqWBbYv19txC0F1LUXmg2tbEMCsXNFnDyf6v4I0enH5R+V2O1h3ZPuaj
9LhnbBrcI8mj7xdmoR9zVw/2NTqG2lqS5Wf2kNr0CUNifXA0F3Gv4XnFFnDl1ogC
Rxdu9QLKEJ6YNULoR8/VG0MQ6MWaUax2FoGA/cQycHzT8+xDN2Dvqp2oNAfJyN52
a4DNaphFudEvFGYYIuMu+e3nuiCNxAQIyVq78LW0EGgKlechKMXDL+4rBN152xlq
cz1EaXYHjFuW/Bys0NCQnh2BFlvD6CLL44mqA8e2xYb8YuVxzNTkJcz+BtyHj86R
XrR20zLxYyClk28vWqugidFBCR/ysJaGLgs8EK/i20YkavrkBezOxej58eTOuVZw
hPIwnVEO1gYQqiw5w8AkifRfYz+byFodH0dLptL975P+an9qqwe26eNexhVbjFhD
Wohh8wy5PMiyn+BtPLkeh6mtwGCu+sXOGNeHRsSf5S3jpu0QbgojAd7zTXQtKi5t
wGO9GMQjoEmBGAs6QQxX/su4JDxs3vGXs9tyoRhZSgrhZ8AXDOi9F+Nk3K5oJ2tj
LG3P9AtUcvzWHB/PNn54JTXEeNqYKOV2md7UqK5Yc8K6yLDU+O8tJ48yB5+EkvQ/
mKGqFrDz6yNR5PyPWkkOehRBQ2bd1/AmgX79+VBprqGoerSMiOIt6Q50sKYWVYp8
Zr9dMngHUUATvaRxGibGAzuzuF7ppVbddGgilbKchoMmyJnsnW2/12HS/Ziy4vCq
gLzURoYZTz1qk4aO6HDQTwb3A/G9KguUnJRop3ovDghJQ4Y0JlWMWHbOfujNZix7
0OIg84TihGOpvr5DqmMTTZQ6KarVQtA3pDTkqNNWtTXOx3APxNStr0wTSoQRNNSZ
RkRRn3lg/OkOwlv9Vn2TAEwxK+mLSlSx3nWr4wbv00t2Ja5F5wDhpVDBHmHjYbuv
cJvs9cCt+/D6zbFZNYoOOJtQauUUh4OEwt08YkkhO4MUrzucf/fVOwVsGn5r/iEZ
3e7neIux7ixv/0pMAGOtQoOM29eQNPr3Z5Wz8PBACuinbVUD44ITIDlX7D8OkYQM
cpmXX29bbn2Q2iUqDWhD1LQSzHMcbNtB/4bTVC06TxmqP6k/lOO5qsipbAfizw6C
bLIixud1FaNaoMu+cwtOQmGO2az7L/H9roMd+ehPM2Z4OrmM6xjMCS2ZFB9pBgm9
glD/LAjT/fzqMzETHwGRiThkQ/NWdJj6gX53gacXbGxqrIEq2/IbDriVrjNgbCn3
g3Aot6Xnr47BpRcaYd7tFGYIC+Pb/s0at/0OvebQHiDA44cwergf5nHcEiLQNiqs
t5hQ7oqbsiZq7BZ0nSpOmLucLyzURBq/npu4tJcRlVOOyQ+cQz1qXCFPK1cq3B99
TNSPaSP/mAoU/GLfHud+vaS+h4Bi1j3qU7G+DhhNqUTmUqO9cOf/oKKKecdFJJsR
ZVDvcyCy6H/H673k9jNdbjScLeTQdyucTSVv8cb+bh36UoeK+gFe1bge+tdivUtV
ZkfRAa69vXp4n6dWno2Br+M/QLhyGLIAYPvqeW4z5FoNJNt39duasgNrmswBtmpE
7+4UN37pCiQvvw5bGMrq6SGMAeJWyN6cPzQVgAywMHO6LcwU9Fx/P/8t7WWPYCJ8
/Gel6K7ref+44j3G4R9nmVUo5u84HKEPZBKz7rLt1yRSXsArd9CG6o4IlyQyod0B
ATVfawYYposnSw8EF4nz6Oyk7GA4vVcXQF6uaQArU7cOTchCGE/wHIdcaX6AADIa
JO1QlYYUzoUm8qagIxVH9M3m3PY9InGw52MQz7yLNUIjVQ0z4lGFXTJ4py4AjT9B
183QoTveZ1LnVDt7VRh4gP3Pa3hl/pnnayQEwLXioJSSzTu/75AuKMc7GRI/vt4c
sSzcPeiSG8fjTgZm9rECAfgT/5yLu7qj1QUKvELN55QJZEWAKGqrMIBXTGKm2oXY
9K4avGSvddlxwRBt3AbbBzr+g2cCWDTp34zqEY3GaBDs/Xhs8M7Cz+HKqZkbGcwX
DLTPkkWeUh+WClnSZUbIbYErb5lNB+6L3LIWeZ9474zea22dM3OZ6MD8aLn1U5Rd
rw/jeyHdVTPt26PxfIkr8fqROwGBboCYEWlG160KdVJL8B9e75S47W9iqxfJRg9X
X4GoYSZPIJChalcPLOqHF17E3JMeP/CHm21Y9SC/umF/LvPf9XkX1u/7JG7pCcwc
i/4uPuMadMBO6a8suKbohSaZ6cPMwFG4Kl9vWbDbqB1xveVNOdFAKbEjS+i/Q4D7
Fn2Iff7jpaLL3d77leMlwsWt9BEENSp7lW1i0qr6IVnbHFKH5Skt2vC0jrlDMrXm
VKM6AfEqYWRn/n5VaYDkIFsoIxo4NA5FHxnw2UgT4XcWRj8/JkD+b55bK5THXphf
jjRTjq8KrPodFCYmMQy+8dXDLHH2bozLMQ5Y1Aeg5y0NIe81WV7Xw/TZIGBpf+Zo
rPdgGHuOp5QSWtERl88sG+Sc4SaXKzIxZkVljix9LbnBjB3SWLH+rzSYh1nOyqcR
gGQEsj8kMOgmlWqOGDFBg65uBIl0vvtvHokrCm8TGzbZe+aSqfpvzgZ1aNi/n3uU
eW5vGxaVmF+aWzoZeAuo5qcKpuza0bBnjBLCLd8Waf93aUrPmPIlHr23BntQPpeL
zUI/gwsaOX/XbqNJqGKNyGPh5NvYiow4gldjndTTUHazHhDLtftIz9rhYWlT+o9H
oGjxMmC5knxlTxOLJHHi11h2iV05G0/nxR8/h1E0Z6zY1gL2RdBWzHHtUKHQPZwo
bx920Drpl855mDChPwXf/h/p43wLayLh4p1fsQmhTST0Vy7poryyRonJL6BVmq28
QrmBrPQZ1IO/0po/1Iy3Cltp09L54eugUNFD0sVX385A6YjEoSVLTOIysUPwzJJa
LuHCRtJdw5HSpJLupANxA/N3gn/SJRfV5dXwhQr1k2z1TRGqSTqniqW63JGC7xNI
v7OWp0HI/jDTKS4idjiMPehaYwp1nRVCmT5sVKIOisa+mL5FN+qQlPkKbGGaWPDw
f4h5acIcj9B5SxLq97zVucI9v1KWN476GM5YC4dius3J8DOyhwlZlO1eWur4KUUo
8KPKGWIhYkUM/lp5an5jAVMk/BNekp7Hp+eE9cvJUQxZL2m7p6cAK/YW9KMObhn9
LBxyfSV7eVZyiFIKimnCeKFTBQ23it6Lg3bM7oVq/s/HkLS7VM4xCgWBm/9b+Sdj
9ncTNARhz3x4bO9L8x2ggBkHbK5oVtF7xwl2RDDqpKCnKmJE1aXD/4chwl/Oq8x0
GzsscFspCHVZ3uOpSnHKdWAOODT/Qe91q1Bed9rtexfeQz4pFTqK2CMW76fbOjIU
asfaeXFZDd0Tr2O0cWX6XHduDF2wxiOTKegMmq/78AT84o7NCURLBO2JcqrMvel7
wfO5dpp/OHyYIDrMZbZuphSn9fqQTGrt20i8t7V8CXIQdTpy2Gy/aMtK3jB1RzJ0
B9WO5zVqxsSkSaiqPExkgumY0Q1i0Ptc5qi27nPiQK3hbO91Dt3GSLKDFFThbJ70
MIQxCnA7Yq8iWpeDeGVsUfrPVN8HWOYb3AYCoqMt9jenANBVRYu13049dYDwavDN
03HSOrIMWL6I+udq6gwhCUT/03TiblfaEdIouQ7a09JZsFxijdmad/nHvu6QY56V
StF7y7eQCoGjLwVId+XnNa+GccDuvAmUc9ZvwchBGPKGmGZg8xluj0UmEiWud+Hr
9Z+F413vMCV3XHOQd6ruS1OOR5MnvV5FKT2u7y7dMwLlTIuVwl5BZ5jLLUrIMF7d
NYfYUHaep/aJSyBJrgTsfNamr6OLiKKxr+NPVCBdkD7Rl6ksvYDVvWxwHDsWJnC+
hfhHmKOF0hkL98qEBnPDxH9SbUqrFld1IZ7nRIgDarI/2uxgn2MBOqsFRgiQoJ3a
LZ2bIB5SSgTCm7VgFORxqYAXTVFSCiPOcJ4YGUmYudAf8qtw5457nmKaNZBU+jVg
c2d1Ex5+VBI+KLKcBAIYOicukxCOB3Ob1r/93Rjg6Y1x/se8Azv5MabeaTtuWSC5
Qm9Vdcsz8MAhr7o4t6q/W/3b47eunWIelZz/FvU4GS3jUsUlxSSrENcOEmYN/35Z
M87y2mcLWDs2bIIRhMqIQRxRM5e/jRDBuSGyc0Y5VgJ7uoN1p4x6nJN7xdctCGpZ
hJ60HnB4FHsNMIeGQGKVOADzvO3Q0On30Yjml4ZPN4ivvvaXcQvRdjHeahjlh8nW
bbhI0fTZgCGguXomjIBqF7ifkjz+4/3T6SaDW1X6dny1tuVcEjeYYR2ceWWXUmUY
80Ne+SrxGQ/7JIiBUR48gWUkPe9yFBhixP7hv5UrRAyYCZc8dw+VK0xDEdIm+U5L
UiMiJ/VGdWL9f6wTWPQSP/qhtwqonYJanR0RISWzelMYZ7mpId47YQchoaB1SRUU
+88zbFHzRa4tR79b8EaFpYR9K0/H3bj/Rd9dMLyRs6Sub35XuZF33nA8H1ozy94S
rox8B9V7yq0Dqrm4m20mL9O+i5OfhHBi4hZZXNygD+j4+0wgO6TRhp8xS5kxDnHz
rW5AY3cQpc1avuH5f8bm2/CKQge4kfY1xIkCHuM5gOxy8Yncw0ZEjuDD5fyL9NKW
I1vomdfIjHKfIF7Tsftg7JF32u2+IG/l0XlSffbV10pD7RS0vIRJf0lcm+LgOgoK
+h8KE752wcHnZFaElrgWK4JECgTABZkC2aDOgLVLKdfrmzSiG5H+S3LDlZrWKT+B
cCIpFRoUkotg5d9+CrniL43fMa6YS79kn/RWTYrwWG+KJ/D513IQWqGSuVte15on
IrMTSNFAVWJ+mSxvhszr4UqzBEvSiSIXo9EH54Ob3HKhI0A/IC6aQoUjIAsaLbu/
SNkTeABi0YqM6BTiVptzfBd25lpuQt5Mj5XVsd9tDQCZoJiTVcnXuzfE9Fy0mCpP
aLAxtRG4+NO8ioOcykYLc9hafg97zauA97H58kl+yx2NTJyIfppf0szALI1ivjzB
w7U+O4Ygld+tZXgaNUYEFXWVnMxZorlFNRlu1h9QrNDWIU/hwARh9cJG+r12EdX7
eBLtOiIUt+CzcMXXk320ADMvPv9107yiEjy/qr8+U3xl7Yy94NbZ/36SBQdAMFXu
TFD1uFngH5DMATrBd6u77GxIIuRzIfyIPsjpsYtw+3iT3ftcdRNgfm5WiNU50BjA
vbM+Y4aR8a/BsiIxDLvoGe05M4Zm/vIgTgjaBa5wl1GwtYIekvkd7Q+Vtnhs294Q
fSGnyQCSEHCRC8mgUUiJ7GSLHuYqO1442qa3h/IBZl0R2N+ZbCNc4GFk5HbfyIRD
pNTmYdOBVxyTAMfNGln6C074U7A3+ZSCv06SkkM8+U4ORq0is0PyhLgPtKX433VO
Ywiavd3w8T+mukcqp/wF1Jau16Beb+1YdhbYjEp4jvoOf/TlMJmi0Xcn5Vgkrv3k
1h6O/4YVcapN97USz+6fPxkDCBqH9b1Kp8tjIIprZAEFVY6/33IqwRNY4r9cXfv8
FCEA17PLaGnblDVVh1X2KCtcNyvRHdSExA6lsSXwc7pfn7dQ2tJcbSPSphPyS/f7
ahdxbexv1/1/Z8OZAWO8Qowj/Nx7mQ4TOc7EdrMgqeZKSmhQ+uH/aqv8lenDrAUb
q3X71q33cI0IhbPA8Z99niM/gRN8J4rO6FfX1a17UetjiB6WjLSqXTO8IACx6355
t4oyHTCO5Ecrs1X/7bNMLqFaoGEn8NqWkG3q/1mB+dnwkMSxctvZAFj75lZmuIK1
8qj5P4Qv64YrBr48a3oDzwPBjSahq7TGa/MPAJChgFV368NNjHpKmFcHiVRmvX7X
Mn0hLc4GgV0YdwGvoq7Y4PPifyYBMyLPLNiAXpwjNoQwSTi++IinefjuaFz8wMF7
AyX65qmJU03SBon8p8bTw8843llcAPykM2kSfu5ks9kfBmb3sbCaih40JiQ8UE1l
6aXVdxutC8PSXMp2eo2ZXdFHDEudruivKZPxPe/jG/voQBvjc0cW2iiOIvGvRN1D
PHG8oeOPfmRYlXSiw1UV+hzBrY442BKpqnRCZr9GtHocvgrWuhCbGdY564SGuJiS
aE6vrF+NT/XoVOPC2A9vbO71a+cj0w8Po3l2BksRUUQLA+1Le6RDRK+Uabk689YF
FOlj3hX2w9OWmGKduvTs3aiBdin8LcVq9MniikZuxSCQwWZAK3RtPmtoXyxESilp
pF7JaSPLtZDMfqJ+HRQ+46eoLy3qcUNsOeNsA79HE95mp7bE2joGVeXTe4K3czKN
xQSHBTUkX8cvczG61TYCFzM3PrrXh0Fw51gwh0V7CpSi5mkqEw2prLBD029jv58M
YGVNiAImrbN3PMJL7OiaFd1lfpZwShuRX7lS55cY/ctXFHteaY+5he9vRYl0bt2+
7dzbBibyHTD2WgfmRuCJkjwxtoJcOVuRcWcCJwv+TXn9vUpjr+vAzxjnNXlt4oLd
KI6NVD3BCVG7uYxTWH02gy/yNmlVvWl2EI8Ps6tG4NvdGxQwcHQl6Fb/k/j1k33f
/DD1fGgma9vIZl5q8qX5RQ+RWvu+PcM+3QchG4W2In1e2CC8yRILBUYXDWgNWgH4
yUAle2fuRpNvhH34oMJVkLEorPbSnkSQxTVEDDgeZx2n4igYlKgl9x8QCbP8q889
pURHwWUaD/4XALFW+6t5bTsQCFJNoJxG9uqzoJhRHimR+2CEILeboLrkItOuUAOt
XG1X8QyEu2FHgQET9A/CiJelpzxinjYOTe+Fab9IUrDT2EYDQRqkv/OkLiswQAO3
GMB6CND46SH6O/tqwytuuu9Q2F1IBD0xJ731w5UklppwZnBlC5zapWKIrDmAYTp1
dGyUALF5z6optnjjV0IxPbrlCjoTlTWjl9bnN3EaZyngC0H/tQt5d7GNreQ8KxMQ
`pragma protect end_protected
