// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
A6P9JbORAheabkrPrXzRyEbQfyx8Snma4mfbiHJ9CdxjzcIg3+mr2bpDaKUd24Mz
2VOQqXsde7ld/wd3zlg3YWsqfhWixgR7VkxaEks6U4dbsrJEjAxHu660CX+yrTQd
UkH8tQIU3NlaOrqj1RiXBNNzy6B/5Dl1GTWVW5SHRI0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19344)
auaWtR13mWTFX75Z8K54/4cuxkcopRv9fkbj4bOs9ppQkXyYRoDBd05zw1I2y70S
bXCQnjhc7gm9quEE3hHCdx4nNqEhNYPnf12eSrvKzf4pWxzxMy/hY3Ps1DwxPdON
lhnMk44C63uyeLdJ2YkkcZIN3qqsUBtCTv4UODT2nqnvsyFMnytLfS785bxDVKnI
ZVRs3d3KqH+2B/BErh/h7nlEqzMzekxRkAGPIyoiDMNYniSnDtKGiXVrXCRve7+4
vR6gDv0sz8ikb89ur6nRqwU9d9h0ZLeBnszrsGo+TFX6gmwPwRlUj004IGuTxihV
0ZbavvLtNHgtcMWVrQYsceY5aFhYcU6ccjp7jyQrvC+gcGwNqL0BIdy62el671Cc
aS6SRqMwB/5ws13ffZdbIn8g+C7Pzo7/hhxA+XnicARwanDCHxq50wyGEB9aA/PS
UNUeM5clVoR03X3tCiL12b7G+qxeGoFNFlWJ2LLcfjtNbcqsEeSshzpzWvZjqot1
6Ioe7h0IaBFq3dffzLIoEGO2TlgOmq+UrWnhBBAbs2Go9DzM3Mzs4dFeeHFLR8GA
N2i+/Kc3fgmkFfPmE56BXwoNZlwWgSVybxAMbCCbIKHZ5oC1KdoS/QMyA0hLozV1
n3UbZ7/7NT77s3Ih88pp9tiZ93kYZ9k/TUQ7ARLKsMZ5mHNGwvUbE5ng89eAiewH
tzYyHw92mO7guxtqk7gyYAHeRc+hl9rscx0ifas+CULZgzkdlS1TbHKZ4uaV0lHI
m8eLzb3CanNoEXPWYKUiKC2gcmHuld/xtSWJrBuvVrI41/okWr6eSAEE1ZxNR1eo
Cwccyvtffi7kuBNyTehSjtDBccdps8ZSYjhJrol47BaK5PBkbhtoaoIaOBFwVYil
x0SQarKsa51rc4HDwiQ2cgLAJRmIsHe6sErwrBT4j0djiPTyzuOY7NQ4QpywMLEI
dNX7iBH8Y14moTSzv5vExRBGOwPmDn55qcGvdqKgce0xed9A7euMQq0F9TXfpjCH
AUYurnXtK6Q91w8SZldnwyt92TH+gNDYuG0HPKbF+b7o9AqRXcalgBj47ndYOaFu
0k57X0CspfkV+yW0iVtJoTdhcIssES1ZDNj5i8R/3Vvcfyvi4cRLdSba8QFBwJ2f
PUeJRz2t3LQ/pToNMAQmpuaETViwfq+o2/j9DqWEuHhEuT25tMxLg2zCKaA0KEl4
drcYDkqMeK6Ej0djhJbI2ETquQb0jU3XecoFCASoAP0DA64GN2JaAOHpkGuEG+k4
KHFYK/TyDTB2EQ3L2E47PqK2mWjVDOOUANAFNvVf3pBysPI1LLVSR4ZRquhXc0Hn
Q6X79PByn5vXwxL0TFsdkVQJGghPdgCPPdAi3lRq1UcY9OhxOIidfjWyvp0v6uuZ
OovrUAFPVUXSZ33V5ZmzJ2KGH/K1SjXVGZIIZrPlxX0pBj8ueihPiZZmNx7MKSyW
FHtAg26iH2ZvEv0jMefsPeD8y67BySGq8MekPLECOznhREp1SfOSUplzwS0SVUyJ
AVsTjcEPvxPHW+7uIPLJDvIR6ryCeHmZxtipGkuQbpdb8/HGuRULNA+5DdAQ4vX9
ep6SYtYxSCmmDptnVMoTRH2XKgfzzuI2hBA64ABJu78sc4lhw+RAyB73GqToOOsN
FgAehZlFitMrEzUXAMY92eHVVB0lw8plhcM7sC4BmQj82RRp4HkPFQT0DipwaK9x
megyKiT0GvHxtMW8YrZsk6KToUVKXyHhEpH0BH6PoJKxeaqAF8AbrUxux+/Rtm6f
gs2Q+RnItHGJ74kJJ/aHgPLsirZLEmx6u2IMn9/dEQA9ib6XI01wtpO9Kg7Kp/G+
epJLDMXb2gTk7RPheyqULJHMt6oMZFeZZjlgeWBlfsAOs6CYykiGJn2CCEPgNAjN
6Wx3CLnACDxzCME8jV0PEGTM14ofdcfFnBW3m/z42u8EHmXRzWS5yPkcRgrfA/Pk
kUfzyNmP7lzE+H1ksTAYeinkxmxzfjE8wn0jyjDtqy4kRmMYZF73GcgEm8w+kBg/
xJMDXZ8sqWRQiiGqqQFY1KTbzjX8wUPu2gTWLQq8nxVruqUsYRkIMYAkEDbsMlRD
OO9i1yJsgZqo2ibSttD5AGRtpWJuEP+jC2qTP69OqghDPydHvvrPPyjZnocXKbfe
0w+jvVdh/H3LJdp1s8R7YlyTp+q7j2x4pt4f6VcpA11l4SjLDrqEOEpK9T8Kfdcd
zyQWduOCxPM2XVqT+0/bejVymoC/7OxSWLqm2Y8sVcIDa/mK3Cl7+IyhpMA9DLgY
03MMlyv8k1MDeYGtScK5zdpor/MP2hEk6b4v13E22MQoc0rSVWPZPjAGqQ8ZdnoG
pqg/+K6fmsA+9Sbbj/WQFyfbmUaTD85Y9SVVxoQhXJWXybKG7eoU0u1YYJoWzy9h
vuFbQrtini8m+egiVURmyD3UE2ldZIfDvRFmGn+sXmfAnqLm9t2Qigbr7n8Ely91
SKRx4sit1lMomE2CewxBvids1BWyeyx9b6ifLhWTA7Lq+BP6DgnEu2VhGrJxCo7Q
S0UvPbTUGo7TWJFQAqUzHm8ZJLPsaFhD+mLzA0AfzdQE9GXT0gimkC6JgT2/Ra3v
uHRvYgibRX+xEhOP4MUwEnkgkPCbew/MjMRlApTCxu+EgDG+NGI4OQwW8A0IfVrm
KKSegBI6TYiz0aK2aluxfmvx3GJQm7FGzXdjvv+2l35Q2+6hiq1WKcJI14w8++Lp
vswwwHjo+aANWSnz5+MS2Mlr/O4ye1vlypyD8HLC8EFAidFWcPle7LIfQvUvpHwi
F1gcUZ9JTALb5HJaIHG8i1fehJhq0FjYrLWTkenSKmt5aK80hryNCzqgqpbmZ2Yp
rYF171ZZploUzBa2tnkrXWe8iGuJ51vhRCwTBq5uxMijmWo1N25IDV7ddAAySF+r
0tmirJjgwiLw9Y/iyizAXNB7phthA5KpkQiSMjEXBDub39e62ZIeDK1UAJ4E6xCG
tu0FTc+7rS5cHtWDd4hV/l77FsvOK+OLeUukMlul6WTCoTLsWC/DjhINDIQqrY2X
akGd0t/0cKLgzfRfOtMh6i7YDWOL33CVP6SHNcIPhfZIO8593+P3+B2d8JU2axMs
b5X0dfCiCFJFbSAihyP+urg+rmMP7Xg8h1ppbG5aP5Abs0VlJkQzpOBw3iseXfC5
rLTE4yoKcjvDWx5g5tOuwJS5PAHthTmDdgDjPEZ0SfbPLh2b2BchWRX6p+lHjLJg
PONmyqvZb65zjWgvBm89XaoT7rDMscUfNe1kQobZ3xiEVmrHC632JcHzP81jcldS
MbB5DBR/ux0TExoDN2+pDIIw9YN+1TIEO5Q9LvTs1XEm5MxVbZJbZpnKhoFAP+JU
w5bwLOsz/5OCyi2WzBy2APuFFXxGGXDtQXyhP5GWkPEe74XBGE/J4x/vh8IjsJS1
jgPTanZOHrSyiLywnCioo45EuD7GI7T4xHb5k0q3L/MtlrqgV+T08YgkntgvfrLG
Ry9WNesX9r37KAyXQAKXQUKngQLuBSudXDTtzrIE6tYIoFP0inxPApkZBJ2LKzwT
FdVMV5aFN3mrXOQFiI1kcB5cchIvO5fJsAV4b4Cv++ECobUhLDzIs82Ii/RUJrFs
NB0F4n5FYnu889Jvpc5vGSlarvIeQdekvI8tpB2TNUBb/ZmtpK8g7KVdsZ6QlAFf
pKCx7jm/vJ/ZVDFbWDuDpa9QxO3P55DgWQc2dkuq0acRm0LVD5y9QzZMKnnWUMel
RpPPl6fNmWhUUPK+Smk1ACejdnXBUVY71oijLr6lZdEhbN/hmumrjPkHiEMc+8qO
T+AC4QRtFQbmEL/2uCSFik5uITuf1/5nf/R6a4KlB4wCX+Vi8Q8I7HK3BxXn/ZSH
qxGDPdjbia7yLOa6i2D55d/LYIvZFa8Fp5cLW6fjIG5jol1Tz63Y2wO6B1iM13rI
QcnVwZr0m0h1Sp7E7clax+nL/AMPBh7Vd6/CUOVXY1dCOkipTxYP0OmuTPbvaxrN
6a7P3B+CzqJT/ZhWP/PG5PH4ltD8vot/swKucxP1BC4RpJDXkO+qSfGhyN2x5RAA
AKLDbbgWCbFo3uV7hho704Lvpxp++dFt1qLIizuEpqE0Og7BUIxqkq0pZk8dJWJ6
FmLAj5c4ITZ6bZy7St5L4bEDJKnz2jZMiYecZgSI57o7te2pqesmZMwmQ8JeCj/+
gf9s6QbHdUw1NLD8DHTgS8yR1H+nmtRx/QLxkP4gIqagg8haud0Ymj6npDF16J4l
67sQl2DpsaRKvRbWW6kIeRQ7zreQDrAay5wkMjgVldEvt0BUORJIbbIxGP4ax0db
A6CTeZjTShApfxI0DLij9lUjhHiLpjiMF4PfS4x2huvAjKMhlnRV0wHR/jPGlbzJ
zAEIcq4/tlMWdbzdSxqMM1flsW3l2KyAq1Z8XtPjz+gBbyInbo0qngJtMtFacD9/
t53GgyEiF+T5grhOvINn/8UeboyA1hdGHQXSgXArz00X6um+F8F2MbCw0ZiKEdu1
nnpkQ2IJ2qGfEdW5MGrxiQ1zJbxNQy7AqNtPlX/Sa3E06n1q80I1aseQnoyOZhmK
FuGQwiz2MuEZL2o34atin9Ukct06KmBi0JsATM1gEn8TX+PyQ91vCTXCOyzNqSfu
bTl6jnw4eKLwxvKbzz91vH/cIy3QcSzdP6IZby/1LaWw4xSS7j1OVtyBFua24xD+
Nm+XxsafhleYtbp+DM4C4tbaaGI/esAtMumBBQT3T1YKcRGBsej53p8WUEXBHMdx
lIEldPEhTO4aHJp1vJX+IFrlwVDtEGXQ5SS0Tb6W4dJqYFjs7XHSEJEQD7ChPVNl
rUPogYRfYrm+w3MtBmPhjaF1OsPHKnUJ8cj2COAVJCwIKHMz1rrRvQ7owN+ljG0t
ZQuhl1Pa1BaWv806Z9D7Q+LNqVLiNKLumK3AA4t7v99Py3G/PVLhPpnNCd0YrtBg
/k7UBQWfF8Tu7BzA6aH+atyDs2EMNO5KZ1NabndZ4A0vB+b3gzcspSNuzVmpWDAn
paUnEXBDP93V/Tcw+MzTrECgAIXwtMsMqmo6e+/1S/KmxBHia1JuHsrgV8XjKL2P
9nMn4Ls5KMu/OB1hupTDRhoIrTqdYfBoJXUGHc6KVJSUwC+QDnsLNQJwgAng14gZ
hV1jDBGo5/EVoQpODCdI2Q+BEhSSsWzqTyGhsx08Ij+sDxBwcMALVO9CHst7V0E6
jgh+cuGqRLiTZ4SfFcvv5cRWk1UHfnu9oI2SuU2ovVeMkUhcmoMxijZ9Gz7hKQOd
sK1uGMeMVItt35S7PQ+46bam0fELYIGCOGeuKGXJwfwJQfIWPqKLLHrNfDMi05LA
uUmDNuDJBy+2cHkG1EV+3HNvLsuYFcEgWU6smxQLcHpPs7PaZKCAeyWbIgyUzpsn
jv8C5QnrTsAyPuBnKHCtTDP//lLNPkzvhddN8pxcucj3i2WW2xSJW+N9FcVEUP4r
ymV6pg8aV3hOK4cNW5YPrYfiRahIc4+7jOUs+aXd2eML/UV70aSdlLjKnohT2HIG
ma+iHRlGeYhnEfxj4dVUa0DnT9iTgVZQbP7Z6+8ig/Uc7Fy7yhLQpt+21OFwUeFQ
zaR0StBEDI/mGActXicEwvZkinGirQVRfvhwShtKw21XBqQrNjQrEZ9eJMBaCetr
oc4l5TM0su33a7/WmyDoe6XsD9bljalB97un+Tm16tCNOxrHBolLSp6dqk7P5die
xKj10TM7kqrJOlp/Tw0WusnAlmSG2HtczsWU6WXPq6A6m444GrPSh0BKWvT9KsZH
0/eCDBJUwZj6Lh1fQ7Mm5J4aX3xXcrW3TfaFiL4+7wr1D8meP28e4f2ZQQVjTU6U
l/P1XgNFctwclK3fEPicPMBzjOdBTEJFu6ww3aXlz0SlKe00O8ymn+AUdEL/VNfv
P5ufClNZb+BSQpQBniCI3wXqC5j/VsrrmYnkKu0y+ctRTeLZ6f94pdgzDvy0A70A
8g3DMkcVBL7xPKZPBlOnljtwxe2d2A4oe2cJ5HJY+XQvaE/99cUfQZ2QGxWwEMPV
6xxDZ0dlYdTp/Dmhw8JDf6zSm90fWB0oAmB4V8vesB/qPs26xSldMV3ccDOJTAIM
VMcW6+mb/130LbNJCwxEZ7IetMu7qGS5fASQCG7dEAV9KUvy7NAgRBVxxPJT6A9K
N/iRJ7XoI5VrqslpOAqri4sGqOGs4PWioY2S1Qi0Ma1H1lRn5zXJK8VsiAQr47g0
9CXmhr52snKGw0Ur2BObzCMKpB50+sYPs+LnxjbIgrB1anZyx8AwUMZTNX8HsS2O
EUbYrIfQ5uRaZAyIY0ZC77dSq2tGCFGc5Vey8BtoAEuGE5XJBYgphbE6r14BmyXc
bGD+2TDbNjxknmks0/jK6xdTabbKN7v3kwQ1FINnveDwA3mvbC5R+jakEsT87hAf
MJQcoZUfSBcbtL4bRLtf0XJbsYIu06Jpa+CSXtwX6nke68E2WG9pqqA//zojydew
7JpIxjWlvYWEKe6J8Z5nQ4zwYJ8pLMHMCZ0NTPC660/olewgwIwnX/S70C/6fm0P
Ouq0LrDWc7BONay32YwiUOHkdxdUf182/rVHnWvhFJbVa3zWbH5PVIbPH3TiIO7g
dIUJhJ8miA1eJ2sj7qlQF3YSdPzMD6wojAcs5X5eNjtyKfzO6X84/Kd480sgi/hT
OCNMjqKotIUGIhUiT7mIWn10Gao+0fF/PQaWdfMOxM1Rh9d++Eo7b/Lh12FS7blG
v1K3w4LmiNSX/E1N9r7sHHYa6xC97z80P6GU5fxoLWn4SOIvJFawsVRMZlO0smBz
rxXe7WRYfBpYflBVzspAQLZ4wOjeve0JSsPW291NdJy3PQwlgiuxXd8HD2XU2rjH
70LWLB3NBr8uDicvm1sRJWy2yECLAEo69tj3FvT02Va1ZlV6NjMR/iG3q7SIyO5g
Ruo+hTF3vRmPmVkZiJ3f5HrSgkOa677EfrhjGHL6mzXjWUph/A8JLpeUIsTDNZhR
718lFuy4jZpPi7cVirZePi6CWPXfzjbBSzntBpSw5rFrksPxMtnSZSriqS5trb22
sRX+ISTnGIAq1lkcYwnJsSg+WHrRYVAaBk5iS1pvwFVlB1RfQZaNTvnmGZprSyac
oiOr6umW5+2bQKCsCRd0195EMXENHnUcNklRwnczf8lwonost7X1C+Bm9qCC7Rbt
4mIOz3gqAv285pe6imEXha9vVkn/f2SRMnp9QdefD0cBV8tvwBvM/cb51A2YxiCG
LDsaWjv432hwGEmX+Pa+IKDuiF9FVCBmg40vQXBV+01yuhp0QyCKwQJMtlfNjgSw
F+50ggA1VWK4rK+4uKxwJLIHUDKO82jjzLKVf2OdCHihtzBJRp6RPdK7Uo18w/QA
3GWBVqpWnhiRzt4qK3o+QR4bsaMzR6mEV1K/QmLnyoAHN4+szYlWjgnVj9LAwk59
o2kvKiaHuXv30+xa/Wxv/G5zN2FrStn7Au7KVxpPQ+oLG4pLJPugm7sWMXnd+IiU
DFHqDPlhbKnlmXz1r6S4WZ7eCDYKy/qw2LUvsyrJeh1lQld76/sgOV/lq+z8gJWa
QpMDDofBoXOJfONVhgCPcwrJ1RMBV1OEiwOzux0n7bADeoCFAvQ40yfLOjxc/PiL
aVpzdGdbdpjlwgJxSXw7mLV4/C/NL+2Diu2tedH26ptrnMDKMNNM+J2OZgpHlT1m
vuYyxKjnnDmWtfVrMiOukCZrd50F9ebLZQUZJ1cnykeQ9MwZDbJ42dHg+mMInYiu
M3hTlu+Dm5rii2nLWgoZO7UmskuZaOjts0NsBaYPZxmMJO+FxeTbv6tpi0MTpyAL
JAauqzhgzDQRAIiYnPi66yEodz6QPH1+hbi3N1t29g8a5C9+JmKavxBdKwjZJ7r+
rfvoS4TxHj7xCXkRdMBDBHw52EVzNpWLlWJBvO7tyQ5RJ4QHixLbfWYajzBNXoFh
xPadPUPtl175tpsKw9infplZH73PM6/hM5waK6IIxq/kuy0JxrGGc3rHcyLe7FND
4/ofsoSAOk5CuDVGVoeVyPOl6SkfI8fPXYVRkg0ykvm/LuG8KXfWPZEEtM+oCVAU
9y5TFRpdSsc4kqcdLNHSz3QffU0G/mTgIBmSFynZFyTgfRuyRx911iUpUGl6yPXc
HEgoAy2QxAT2l12ryP6KO4oAmzcGK5z9cSkYKZFYm3Es9ZwBtDMkz9rWhKtzsIys
8BOPU8Pm30ONKW8lAh6NQVl7t5X1wG/rZwz1t5+jmBDktPvZmAko1W0aQ/R5yrUc
f0qVSo/u5b59rV+Uc5TLU9bSzPD+sAVtLjzEeLugh3jKdL70dlL3zzf2yd3hk5AQ
akFoVZfYJ7aJaqutA78aP3JCblefP+3ON0VNkqCpUU01iDVZ0nH15NTl+Wa/b7uQ
iKqDZiLLzldZl5XTIiNhJhh86K4cFag1yN8CkLMtPlvy95yA3p3S9r8q80ABSWaI
vvuwHN0JvrGkF3Z5TB4c+bq8eqnZmfPUniTuiL2fkW331jmlZ27naHFCvKdJvq+M
7IipuS2dEpQzW0PcLLI9L4aJg77oL2ZhGJtb0KRXqrRSByBhKYcfdhxOtrAP3hew
wb+MfleT021+z1OBmoy1RCaxJ4spwllUx1fb9g4gtvfToLhhffWxxp5W27jTtKco
be5G0VljQ9L3yr9QBqJpuXOBmv74mc4+U6EcyT6DfzJVcPoysVOj0EEiGVcs+oqt
qvXTGz8ScwiiHmu+q2cRbnZqIdZX5DQ6vNYcWjZsokdqrM5UqirYKkal9nuOD2RP
fkhcqVljgH/u/F/Zo4ntghNfFHCiAUIDsaiVMEtoWBTzPXAzZ3xCtBaEwKCVjzI5
f0yZgPE2RZ+48QAZAP+Vc6FtcQmPxbCkf0uMf+0cxCk7akYrO9C/nXWUlFx8XVd3
UCurkDnm6B3cRbdi+HzEZMYhyUKM1VZKXS3INIuYY5a6HpGswl3KdRrDZxOqGR7L
ZjZ1QgFtCSTGwEUPwW/HumOl8+ecIIVwpgezo/cRclXbPvHpmHzRymXSfxqqrDnB
fjkax4PPVWrLbQwKXSfZlHOl684J9YvO/3w33K1uJcRFrg5aA8Tzzq8FykErPu0k
4cZrsQZVAHWKndPlH8JJ4ROtioZUkMAkZxosYCMG8UwImrn7Oz+N1DBLKR4Jyulo
pmSev3tZ1FYv50rrT+NSbONpOOMYUzGZlPjVYnnZXhFrX+J3VTI6yYvafJr0NWPL
XRbIJb6RVsZah0mQ3t43zSjmMVQn9LCKJ9bXbkJNJtpE+6iBRM8VZjyg6nQOEmT5
edsDEh90TIzmeP/4PFBX7aFQZIXR7o2CTImLMPeuZ5+OK4ORlIjxfC6OMPWpUH/b
V9Vp2m5JH++eqIpQS3NaR1yfgMxtSC09HmRGRHEsewSyLzgXs+u/udjjUoDHGDWw
Ma8bg+X2BFBc1Tw1g17/q9ZAbDJ+Lj5K0bACqRRUY06u5ck6fACm8JKbPBoIno0O
x7kqxsqll5vvt+9aYWUbvr9OIpI+2tAB90Ql/QNhp8zwFxrqJ4mD/mbvDF9TePbl
bkuMyKGeadG1z4AQAUn16loiuE3hdc0fxPhw648ObiuSEDpnqHw6Nd0cfkKIBEfG
cCcASufFZ/2bBpkoPmdgi30O9y786MAo67cvjRKyihi4sw5b3phOAeYeAoA+PgsG
r02gNw8iV3P/5i3t/8rMnhglRixlXdX1gSMoJk3XAeL/NnEvEOW9f5rIDClxN87d
2T/ep1Tm84cpx8IULm9+QiJWjR2z0cWY11UZITWfEamMuxtKJ99Rmu0wDw91mJvr
J85d5/n/DZ2x573bX0AmwX4Ghv6mRqAIcuXcDKhgdXJk72AGvgQUhk9jCwJx8XKB
EmqsqLYbfFsMVWTL0mTutKnQEnFbu9Mw0nbop4V2AfRlC0kwr4vbdovav5X8FgaE
2K6r+71upiOtZ4CeeozaCyokwvYjkiSZDhG3lQ+mqbHwSZVyhnIbCb4TNNtpGfqK
R8wOTJZjenOf2GfjLcy6BOzVTVR1meoOV73C+tsfZfZjmOkxxpEPpy0OqQIjtfPX
3UaeHok6JwsNNVi3v5LNPFY3GGjoe3315HNAJSeCl0F4BIDijn1RkmqM7U5keU6Z
E0Mn/dA41TDAzZHv6apA4GXTfc0DS8yWlmC2PTtg8s0/FbgLJx528M/6efcWadxI
9tNEs78nUO1FBe5ibMDI/I0I2n0pbscMuwmaBUh3UgdouLbXsBqWmb6P4LGYMEI8
wu8rcP9V0jTw9oG5LonKBNVjAVNzUH/elPD3BDSKEU+uY0b9TnoI6T+kIc5tcnr/
JAxw4tNR/f7aMw8CaLBh69mtXmVtfQFJm16k6Dt2LtUIQjSNparYduSgRSFEbqt7
KbzeFqlz6acDQx4YarS42sQokVD63FjKfukMsNLJBu35s4mApHfAmt0Y/jDLxzhZ
sQ6BXNK6YYVNdRjj97ocSuSbzFCfqL17wDMaldtLXAGgdyzMVljLn0iVykyARhUI
hOjokwuSY3DhI5wJmGf1j42skrq/s8kNz3OEEXsq/UJxh5mhoZKnZ3BjoagxQ8ao
Z9Olpf1UCD0FNkZm5Wcm4zmB7DVpgV1IqBrpwaP1YmEJ/WvOnMD3dS0EgwHPmO+o
6NDsP2kw4MuYsPXRK+Y+SLRZglFQACMRVhH6LVmi+/wGcUyC2QJzS6bOB/x2NAzk
B/VS5vScIFcKuTl6Hkfa752fA2He1pcWfr7QFp0CFy+Rqvo7l1HZikwIeMXV3WbN
bLxdJrAd4L3R40X8bMaqLEXpq3SrguJgxGCawrBqLkqdQmInSE6+5aIssZTXJ71p
QAMxy1I0vOX3cA1SAESCZYeCUncuNW5uNoKlopCqG7WqVdVXQpwxUawwenIJqiwY
GVs33xcl4sU8lDIuk+hXHYAIormMyFLqGiPeH5zoSOWIgyRq+t1jrzqaxBjiH6kd
osnr4l5BBzdaeUbtd8/o1tdXN6N9u2IZBu2WKHkEV6dFR1VF0A+BjgLadQhJ9sII
CnNLmosky8xpfEhYqS21bwxqmydoHrhDKemce0OXmrmvs8paYO43w5EOTZ7hwvIZ
Qu6pjoXeiM2j5KS0rum6pPKMBuWEEg9aoJnYZyzvnFcXcyxBr3ZIuqhVWttjFnub
aOcpK6H9cCBMthvSqj9Nt6Bliu0u/6nyuzFDeYASaCygQm5tyR4tISW656VWdXkN
hkfxt+BNf3Bpr2mNP8m9CApb4dv//ofGgYiz8SR0p2RBs7ya4EkRHL+HDWcqOm2H
JHQ/XNbgkbJU3hxJJPmgtzTczthMmePvD7uG7bPm+ECtm/gW2AOvbh0x2WhxICo7
XtHWzy/dK0KQECmjjw8sMUmR7kjJ86xpGWGUIysN98DXsEb7tTyZagWrF9BIcawN
07gqqMZzxVwpIDoAPdT95NfLxSf5iLT9g7LcGJDtNtLTr1Ryi1GSaqINaNLcD+va
O86wuUhh2XXsYmjYGzNWxgOaW9RXw+iwJhizJNVRPA+FhdwKkzlNiKYo51Y5Pd9J
qohCWuZ/SsozIlIcpbCwrBeFMEvJIRms6faA81+HTbguhI+TXe8x5elkNGlgcyI/
MIhmyPlay/AgjVCqQnA1iJsnLZNb4QZK0iusxVZUXS7TBb2DNQIq2UCJ6LX+RUVA
CXefB97EeJ9nu5xnl9uXEljnPnNAJ5unIpM/C1R1+/YgqdUMWVuTdrd6hvExcg1J
mtY8QxnzcV6fh0k3TptMxa7/a9hyBh3WQUT3W6bBEDXR7k18Y3h0CahIdIyRE9Q1
kTB+wSLywGJ52NhHWUYMWN6u8/1QYuzVNW7uURCo1Z29bgWCZRKW78kAL2PM198Z
TsGWplXYOLALSTPfrVB89w1UaWMoxjKBOkmQfhiICX+Ua85paC1873RgI7kpj1UO
peKtfxgD3qyuhqb4q+zy56HioCK//YBA3HxwDx+etb8ztHQrkDdzTFpeWKbIjjCK
WdANszXbaBs9a8UY9Kk3HPG6ba4TrDLewPWNbfp2AtsKQnohZfO6lnm3Co0QLvKx
DAOtdkalZ9ZNnH6yTW3l7oCm/ur2h1O9v7eI9Ns+Rdaimw0jR8xZSQmBUw4viZIh
8LMR7DPIOOkhYRpPISO0BwN0oSo/4141HoCNVv1zk614a8kpXXl5zxcLVRJyNH67
oJ6NYjblEMZj6KMuHmMA43z1ke4nq/CqxwJZkW/Pfk07V7TZPbL8gpVDgEKyw2VC
CQsarCv8A0PAODLpTKv2874ZKJupkrU+wA/+P+gQGatRJ4u+WksNaoXwcqnZCnTE
GCl02k5S5GzQO35lF4SvLphAbNfy8KyBJqgyA7b4cVyYljke53EVgXf+0PPyCrFF
pZp0WC9lNuXQIHS5WbUSVNdfPCz7C8b4vpmVgQshI03JBaa6xmPU8XkSGhB6ndIg
6hxurgYL0HZibmhy866yAMYkKAJQQjBCILuCIBmJV+oYBbtCvPm/uLlvrLnRaJTi
zLNDGr/xU2gQw2wCe/FL9u1gQ4Ycng1JdIMhciNNzk+DLErjWhwutfpm2V9jb0Jq
WcxQ3kFfwSZj8SPxDutgz4yGgp+3fbaZBPuikXr6ezdBa/dVZaD20QxyazYQAlki
Ahit/pAkLwv9bI5ILTpEn6g0bn6THG/vCs67ZCGjAR+wkfCFWhSyBosD6M4Qn2NS
U9ZlYaK5XD3FGCDZ2lozO5cDcQmWcQ2qfUbWucdbjS904FS7gTWVNgAf/5zyBQ/W
TQtUwPCB6XdVyZaojVR8UC/tU6khzDQkgPpnWKtKtY1gOFZc1uL4i9U+6RKfB8uM
A//r3qo03LKkAHFXajctigQKSBRCBvZPAgfUlJ+L8hEZygTm8bp5vAs7QJlFLRkM
iOap5UcYfskgJXRce5HUMX72ls41neuZfQhYuPDGsudUx6weph6uJNoXDui0JdeQ
FrMIYDXTFJhWo9e29mb5Khq8jqJfeLWDC2YzPHe3msWHyeY+yoxoGMO8wJ/1vBsX
1Ui5EhDfK0iSQ6SHtfhnHYg8PTzF2WNfI2O13kG99YH3d9SDx5rRdNY/l37V9Yby
BJCqmA++ho8t7PVVW0PAGbjT4MNVg5xhxit1SGjQNsPRP+CifNt6MzBUEHjWl+SK
2aQLHE1ebaRgKkvK5sS5dQBa5iorPNsABH5y7q4rZnI0cdcYjTShITqvc1sfK7ar
gslVe1Mt3+oFf5efVSHiK83Q9KVikZH8YwydKBw7qZZaUAUCQEQq8dZTq72nbzb1
v5aVd3R6ajUwCb3BqGFXrvIO+tFPlDtVMItMj6EC6/F0MxqOpSq8bTHpQMiOqr7n
JaFdXiwpoxi9cv7zRO+XU65MKx/X7FhDWJblGcIX2I7xXC7++sb+86rIbCeZwd3T
BawVxdEe3fZBOwx+F9iEVmCif2+iTJo2qE/hl/pOF/FH7T3dwNRlr2zxPVl/JGWA
/fYAaKJGGSp8Jl8vdHnHYdX8ENX7He4wTJ95AlYAj5EjUGDfWekLIdFDs/hyu6bL
v1bQotTzfmmU2tnXQZMHjRRPb3q63nDV2fqDJ4I5MnbuQBSWxp6OYYwRaXogaJJ6
U2DzWWQy3nxW8jh/jhBrtsxqpD7ULdB3/xE6ZbkTgglciAjVdRfkeIVn9ECJeUSM
A2e/lKf2eElST6n4VaZX3spgJdfGtmSHQYRBJm0efSDlEzJPnOUeKR9Aaz6BrukV
dihFtTWBFnnaat73OGZZGl95pAQ1Qc6W8TlET5ncMgXRSJzUVFX2fafipWJfmfIQ
cx04XffPe0BzfBOd3W9dn6l748mt4AXQ1gY4bqCSuF/MY2VeHZm7omcCOwTJSg2L
zuooMHpide3SKPII2scWwTAZI/QKe7SAh7LKN0cj+GwhSOIFjjzxp9kfMdxFHqpO
pXM+UNHy3KEcLVQV1STMb1LK+AE4opz2EJwiYuX+6ED19zZSwu736s4uf2c0miGc
embWZUvkeRKgR0RVTjJht9OWGzmSTBiL9mLgzzLxVv1rNbQJ4wBEAdItKBuz9uI4
BjDekqFPDRshDPdsiHjCLURoSD8a8nZdqZ/HIDj+Fsf5o2YINmUhnsoIrqJwTSQk
9o2NcYDWKAUrBaton5FNpSZJ+w1KMKDVBj8e5zv586rqReXdTqQNFyElrKGaHNHg
6XPGF06CAtyhRsZwh8Dd2jaPVWHIrIvczN2NIxglihjoS2BzXygsyLgE3jCNWtm6
cJ8p6K9WcqWT0FZiFgRUAIw64Jtm0yyX/I8n4zFcWOhB9zVJk1w2X9IzojAg2HRh
UBXdVROGal4MxBsiuhiYf1wR6BtjhtyN+2yDs+o/0dLp5lWk2JgGME1QG9T3mUjB
2iQGPIpZBuBv7rGqK8wDTk+cG/b7IM0oS7Q21Tc9F+Xn4SNfk3Gw+jgv+r6EcLV7
d486aXsRNh/EHg6GUAPbCyer+S5d2y1xMZUKH7FqLznFbqO2uhgQ1s01apbB5/jz
QwLLalA3G+CkEToZsCJ+bJkf70cjXM+IzazCaU79Ga5qccc/gqB9fudmx3kLhTQ/
XABPsnmdc2xYKqSsw9g0FZmhHFi87GnjchSUaYAUeRih6nCCekbO3qoLb6fCdDSa
9s4NokK8a3iNBkoOLTQ+gxTc2cNix1ChVCg/yYwgF0tsrq2qThMd0pEiiN0JPOux
w5Y5rIpM6FMhzd5xGCK0ruGDCVe9i2y4U7egbSSaPNH8wGrSuW9Oru9fprQmPs/Q
1/3lgxQkJ+24vxgAo2VQCKIgF8Nrk5dg3w47h2u6Iz9diH8pstSMXMjsLA6W8QYT
mHdqyFkqvqtaINHQBIMbFjO7KH0ngh9P/jGKhhB1F/prW3T6inV9ZA+BDAUdjjXc
+z5KNYLH4itxGo51G4xyjB4GkHqKCOlYBR1UTHv+TQUlDcLxO0/ieYggE1PYL5sg
pIjFM5JAphX4jehnINFp40IusSSIcAjsFo//L9zGwj/yDG4yxa8chUyRXx0bpuLZ
OZWfyEcpA6zxsvzQJ9oGS9f8VoOobtgoVYBe6gXOTV3TFBAlRLCWlGwnhHtEYQTk
lqFxEogpcilgJb6Am6+ZYL17MAsN01f0piKUg1DSg5B47vXkszxPi7I0mQ9p4G61
zXBjm86phZeWKDt/P+Z19OChqW1L2exxGLzIhjMy/WX+mBJaLfWEPLEbhpUQ/DR7
7cbabcxQuh4bXfRPnTF6hqE4T9UxQt5eXMrruN+s4N9LQehhxp1zC2aImMXroVnZ
sTMxhB3XhEg4vNKBFN70K8VrrTi0eoSz68UZ+iHI10vlpeLU25s49z+Dj0IV6eoO
M35RuAB832DRwomY4rOlOEtKvhPXfrhhKy0FnPgx622qapGlwbjcW/4Jaf433wem
y1jEHAarRc5bTKrWG042jncEDbvtvaD/03OFnPo8nS2hmTYicN5h2EWFicE9KU7s
rmDsPnhtIYpvRJTlBcvLthPXcaNg6ziaKISDsdOvCt6ul9j8f020m1I3LljXgtwf
oeyxxsji7gfE5ITYdKKIS5IkzZqUPmE/mcSCcVAnaS0yjqUSAu+rE0E0MZNBEYm6
ePHuvP/kX6I2peo8SsFshOLYiHvnIByqmLlGdUhdXNfs/PhhlXzuXylXPx++x0N8
IPW8y4OQWZAis6iB6m4GsaFfWPUAh/sbjPmW2dn1E1a0GPuMuQ+HJcaY5SHzDh+B
hiasNb99TDY38eq0k8VC7ilWB+P+kzP45uBsfZLF/47IjVzGMNZISvXlXKH4sVMu
/b4hYESK/7LpdHsGicFeiJnnAe0kiMAN2Q63ohVpuWZcjenqJlLDSFl/j2ek7p4S
vy2EHQD4qaTBPSsxdKvmvNeDQDLi+Wuu7+cqbPp9W04d7rNUMU2+2nQ/VTWhJulY
UfCbBEgFt03WHd9V+m/aSz9lLDtpm6nWUbF/laA/q+8IqpdgLLc95XuAxP86TIKL
dOG6YWSCbRMoHCFQr2Pl5VOnOxtqwg5/po3dD3LMO1iYjMb58hkQYeqwUE606/e0
RZmAlPNRqQIZxuWR96JSIhSY5jSOekd4xSezkPEt6Qhxzz8s9TuzcU8x3MaNEEEV
lCtDBbYGLCN+3/mMzFVC3fetHoeqdYswt8dHEaJUJ/nrJ+SRoUyndTJQQMRIC9SX
t0LBVyFqTn/W+gx/5nyc6399c+RTofs8uyX8+CgcufFvHa14Y1GrAV1Rw5bCOxIh
eaCe2JNy2qtT4ktxyD72JeHeRyqZnvCn6SUPAVLJe7d54RMLB/jQspUYdjcjlpJ4
VlNi66RIOircgSaJPVa4CA0tRh71bL/4X+mQvpTe9oR8YI8FNvNYG5VEPkF7LO/i
gxDKw5/2GXII71+d1MUNKm8ferEdqiJRUbVjknY5LkuvNLlWjRadTg30KZ0YLhg2
T1bvaX0ZZPP1dc061eIB2YsxJxh8xYXXlUInD0A881GUdertB+Qn3WewcVFla6qA
fvA/DX+Rejcui91f15OhQBPxWVYt/kUkbNtfNq3c39Nodav9OK2ls6E1rxhM+2OY
IRJvJl281x9lvfRNqQ7aNyIUm62koN/RXIKh9HXzymd11mJjRp8dk4SEC2N1g9T2
/FAGKTDuUQ8Mgk4aUmYvpX5U+MVTWsPixo942qYveEyO9wS+/v/Ui4kwNr0uiOHU
27eD12VmBbTuefWkeqpCTcZElDrbfX0rnnKqrVacLGy1HIhlKPmoKae+xuIKV6/N
2S0AL/NzUXLrSPoJf8R4TM7aWJPcaaIZ3jgbKpKprylqBFCL5pXw5NDZhlTqeg/G
Caf4Mdr7biUrmGvl3b8fLYlsx0KSUsCyZJ+hdryf4oHAS1UnJCCxz9DxnyNEtLu/
zYrH/JFsTsWMPGpmDFVXlZp2LCgSBSM6GI9th64UkKaR7tVfZsK4GTCG2sMzCqBN
AMD/tNseIDCEDYQVTVx0WnIWU5aFfGLm0r9e+pqtpsykmnW4pt+PSfamj+HcysX8
rjtkwNsKlT4ds/doP7uDrkKX4VxNVq3oe1Ov7NSkHAbsSIlQhttQFrZG5AhA4Bm8
DK5R3zP8rzIV1coy4vQH5nhA8N1+RIxgWQOUUqZgRYDyltlfGLj67v86b4KqBbir
0wfbrgX3YW2d0GbTP6riFkKp2s1wC73zyeVeXdussrFiB2LfyXAWMfcSn67JhWsi
w9YpLpER1hKda4LcsHryyESvvyqi9Fz+fmpyu/oCIyhanUsugtH1j8ya5SrJ7Ptr
MAQrmGKhYAdzW7iQmwfXr3ByJdbRtq3V9VZIi+8KDaftX7/5WjOeo2Chvy0FM70+
guwok2MaXMljt6mPBEBBkxQyrMQH9FFdsQYdyAWuGidTFU6tarVASA9CyOoo2E3r
YvmxkB71SbA8M8IvQlKEK4SzZyDRxSI7U3zWUWCX3a8wfSuSxvP2WEhZcPdzbih3
zVnyIDALOu+nUeF7Kav1PCAjmn/Z9sczYevDsGBfBNO+FdQQcURUorLJoaYCktVi
J3WXt4abEOMfVCJS7TdAJfB9Hz42SSmz135vWI8C03/jN4n51JgC0VVX1t7i9rFS
U45/3Pot3w5h9SJ2o103Q9rBcj9bNlt2W/V9R+yZ3kf2O8Q96gEKKd244zmsR+fd
BQPCoL5Ch4BxgUek3EOOWcxyA00xJB4v7vpDtooUFOB7dj7ovgBgPJn/w5G90kHj
gRO4PlIhGpQRWU2tcllyeH6oJxv4Ua7XHYEzlmw+y4SUQdYaDFRIQlg44a+tUfA+
TDfqWkca00u2KFBrM1Qqj4tDMLgb+XdkBZvyW/OCXTCyoETeDIA6B2fPmIq1Zckx
N5jQnsM4dpzMWQ8YdxPugr8lkibVHQwpwADzoFJIxiyrU7aU9SUU/Fx+9ahgBvB7
3kG0t/eGaVRATWa6c4pKERy81yc//1M8wmdqtRu1BcFv6lBnLkJwauSmBE/EdkbF
Eb774dDUB+KY6voIaEWsZmVAHZjPTAq/gJUSb2koHaCruh39Te3hRFl0VyL7lGl7
91rwMvgvT+oXPsqz6eN52rTiIiJXRoi06i61NS5Uq3Oc5N6fQ9tj/3sCWzdFpWtd
bEglb0AuVv4Wz7uiFFWNhYnGlE6UtPYHEOV2lcUcdoflHOQNv+hY/lSnixgBRWzZ
zbBKSxGWgihmXbUa/cx6zK5aLwf0LLjqeG+/uAtaR8b5QxB9XijX3nw1UQ2WSFHA
cpWgeCEn4OmyMiLT+awze0q3ZuEQqX6YFCbwlTIci0lAbg5Qbm1y/BEJ4lcOsXLz
jchkpD5N8ZMb3MVs11vJ++UoqIQ6Ztymlqk/zV6imY9ry1wlP1jVT1qt1dOdcbqK
57N4I/3Od47XphyvyA8MVV6gZc8o/BdkRvh6KIYoEOwuA6EH0sPRllcv9AuWMc2z
G4mo7Gj+Po2BDdv+XkxlME9WnKGiPeMWA/OR5XzZ7SjTCFHzBWhnOJTW01jAfO5U
oR/kf43j9TkaxBKI9Vl+m8/sHFQlVAxld8qs2y2L4gPZ7koYmeW06PGDkrSlo8+y
6HhStIoXq6uEgX92qgBlvK23ugx1B805untZ0d4lrzDM58zGOn7UWpKJNRshf5Gk
+7xFnCFggw/Cn7DsoKWjZ7NgfFi3r+qYcgbHQNqoOpe9k18m3S5UjOVFkwg9GweI
94QwPW7lkshcmj3ndbaK6c+A98VyZLyTf0llTpnY4/WPj8xGUVl+IK0Kyc19ZRuV
+3UYcp+o+/e4ketA/LTGD4F4DutOd0ivS6UrtqzchTXqwr6+NLQOy2dYtldXnvy7
dK+8F3He69CmqvNx+toGGT7DVKDttv8mYGsSecnjuKytcL5thSgCaMWOY63/SNtI
5Ilz4VhxE2J49Gd+Xiu9Xl2cNsj/A8Uk2kBVWX5WGDEX/E3MhLAHLOo7hBMbUt31
j5IWMSeNfJDFo/nzN/J2T6ui2qPne9W2B2G/8P7S1Oi+u5QaKNrMlWaPq9wWYgnF
detVZrI4WBGNqejs3hw48a9s9VwqcHhNl1dw9v+XgTRIAhwtTeDddMF6v7Fi/IXR
gd1tuEH8YXQQRwUkgf/yX4W7buXgrb+pz62S3Q4miFfndyAwA+pHdWDhUEUZud0t
7SavMlULKNL//1hTigvArdgUXYIHEDI7tud3TrhvwdTddqfhaO4ZgwIgVGoRwb8Y
IsKGmFinjjeKdkGaXfwwE9hXp9fmXIGMCdefswUwK15K2wtUzcj/EZyXXP2gOXYw
uyn1g4n7y0z/wU88177rSR0BLRHf4ISY/0OdP6R6LL1z7hQ+OVBVlcD8IkO9HEOK
Mh2GPyD6stfCecLOay0zIDD7AAzjasCmDlSsP59HXcngutRNNQIdGs14Dn6+YbUu
qNUPd7DAIkojK+Fc2LwIjvQ+1N1fuCUGWm9J6fTWjxpOI5EWIDX0oV/ZL1dAW/Ah
GQxUJCgzB3Sdi6uYwzS/TVNlS/ISVViihBTG1x0mQU5h8wrJZPvD1i6JHa/dU9xB
hDErxcRo/23Vus23gQczhIOUpC97sMUTk4ZIkeW8hbyHeihDCIxfwY2yxoOrOn+a
nMHqRk6YZQ2mWGeSLGRjK63slDKoctAk4j4ZL4XOKEW8zFUIMGn1O68xApwysD4D
E548z5c9DcwC+lUaSqtqiXPGUtFa4j6857B1O7rezJdSYL820Uiix+592Q4OLHkm
uTaH2q7Ux0Aqbu5RBlmAMnSSi5xEyvfWfU6CVc0IRNNXmmOxAInGupso1V2Z7zjK
g69QMxteuvc+Vz4uhlhlVYCKoRzvtPNpKsRNC4BpqETZ7FWNAPZK8NNZHPC10Rew
+tRREYRSY+oz6QuFkwQiSR/xlwiYaRo9M2JxAmGSZMsSbSHqcB/1mfIiAhMc9ron
3iDY+QKBeewa7tS/3MY6TWfBDZiLYW0mlS2h8vxoGYVbUloEYnxy4EmJsNvqQySF
CMbaL81VBdK+HR1J4aDctxkoibMKVSMa4tqLvWl4nQky1ll2/TJIpivxuREXep83
Omg8zNx+NAq33C8D/BBUQ7BJp0nzmfF5gZsUJ6W+nkIgYB4KhNyeDtKiHhyug/yy
Ph4brQMcT5MLw7spxULcq4VdoQy8SIAkZdWado/kvKTm4SaiLUC/UCsl5QikefFt
aqVSr3+PHa+udXIjKyYei3PrxqfMSw8HbDFxTSFwJN+DGQ9crn4gIFfVGYpgi/PE
T467w6wwFiZwU8IEkottt1N5sDt6HiisEuXa1JsSeCExciMG93YzA9C9RyjnnYSA
r7bizoeajLilzg+j+gWI/Yblgwa2eEP/z8pX+FuY8xzn217Y/rgpR6hksA4SN0ft
zSPOH77xp3Bh7UBiUpZ5+pLK6tMdFPMbYot3RKjeHjCXzFYXGERmJslyaSBqzt4q
LOHwOCb2e4Ghox24v24o/z4l/omgsccBrM2Y/FLRWAvI1Lkmo79O/Kv9cdBTNi5o
ZWpIslYDavo/CwxyOjVPTvIby8dB1fg4cT9mzyLA0O1FG/7qVilwLtI3eN2y3Wg1
WegbK4cL23i3lqHWgOole9/XOWj82El1r7V3MBN29eLfiDYDw6CwO3HN6RjuidU8
o13RDlq2Or5zsZTEAjbxgx9fntC4y1bEPgHT3iid2ddiFv55beCpERdODZ699M0w
ZOONd00/pGCPgnPHMCwhiqjd/Iqn03OupVuzZ9waPKtcie4GitARNI77ypuqMDrq
HvGBPapAJjkSJOWtqUfpRCCjcaaSAhg9wJA1ZXZ9qdtiXMLGZP60DhhiEDUbwCGa
GHEN2F8z6G9omxtTr5d/yalCEXlryDo9eKwXI1eNNbj4cJewvyjxcsqh+FzGaVtQ
Cgx6NXE4lHK0siz3yMsP5ORW4AlKMEWj52K8h+LB8w+c+HfLm7QnqheQJ6uD2bBC
Zm1D0PFntcHsF/w1xkjXjfz9RVXwuf8wj3AaPHNJtt3W4wtGzO+bsR3vxpmZwJk6
NAzL/e1Ktozzuzd++CpEesKshiD71+9IYKklJhqtUiIwFN6jeo8kjQ4gPJAFXfr7
92fDq/c/iW2CfwfkgrNp9nKmY1xzIy4vEETAOP03p+Se4nkmRIZgrJoE15cbvdBr
+lzi6lKf9985mYrS42GnDuG/IVAhHSQ7YZ1IIh/WN0FtYjEn17CNbXcuVVjEZLjH
r4pYjv4lP0FZJgzx7dwZD73dvspju1WypEnAiv5um3RupJ5rA10slgvjvFoQMjQZ
Dj8iLOaSIAr8GF6Gn7c1f4q94utQgMWbym9C4of4Ii0nVFpfpHO3LxE54iIY8uQG
WYqLb8WZMxLqwjlr6wrWE7mA/K11VHT+5g6SlbCNSDbFyAsxXoHMI3YWSteO3y0F
rWhsqHqw2D3J9cuvtxrsXY1JkpY4lMxBGiab5Rj0LVBPioM/sEOMVL5DQauFld+m
JWuyaA7f7wHx15I+FYiVX00vhGNlg6AoPAH+FFOIWRFA52vhPpK12hoB9JkgrPpj
EKwMBBkXzaGDsY37ifmGfuSfruC7PweRuoakGcuk93ZzdzozRHgTsYnQUB+6zSHa
n2EzwWQyH1ELVPlJ1AeM6NMA1UJQBNwcgDQMguidOP51VKbwgZ7w2lUT+/0TWJRl
N9wbZ6bH0txlY4mbKsyrf5xXfrm9ca8+hbuyoKV3AsdXA3MPUwaIlgvLGpmY41bW
dBtJQWpiMGRmIskc/VF8s2PmnaadUbuli1SpdSwcq0r0aq+0TyCs5415A2/5KpyV
hmFFA1Y/93lEJWeOESlEzHv4rYZnFOeMhDly47BBIt0aHcnK8PuPesBIdCPvVlbG
foe2Iv7iXmqWLO9PNHwNx+zaTJeJ2sQ/imkMveufBDTGpIBrEPVA4wqfJoPQhz07
HtmjjerQPUcnJ9Pne+rjozwx5aH8yfmr6UBGFXl4LaXJs9IOr2Eqq8KlLxN3fnjn
Dt+RiZNhfPIe0/FJ+PZLOQevmDfNrrEEBBjY9X5H2m8fU/76M/L3P4TJmFBZZYJ3
9uoLqgtfSx1N4jYQYzb4RvCxH2I0OCf2PYEZbpUIRy0aAGCS3bwjK1FadzKc1Owq
Wlv1tVlkPxRmB9G5nVfomJVkb8MogLfkn7CNViM8iwOzMMaQXcQ0pnfq7QcUhJtP
0qqMfPmod5doajB+eq5a/MZDaEquqka3kyQK6ZNy3Z1uI2cwuY80M8UI8ixhPsGd
Jkhm0x72BK+5yU4oQr9II3+KNsW8J1fIPn8YHDEmGLVO32qNC7oj++cct1F3HOmH
ZKY1aEo6+ndjY84yO5YLu4rKv1JTUIDMfk5AYBXVV3crQIe3NdQMD/RlC9PXQouv
hZBNS/TJYRFZEaKJj5WTq1C3Aazfau0WXbd/Cekp2GPlkKsIz64FnJw3nEa63L8q
2dDmMTZLkYOLok4IV3ToMnBssY0bNztFW3nlJhMqNtE3Mv005GRiP7dS9w24aPR7
dIh69Tl8EqL96T09tJit5myhGrQoh+9SLO5QC+jui+wqX8DuUOsuow3kpXLtHgt4
rXaPpPWm3OjbqRMaW3+V/wsjrqre+N6yk4wHfGtlxlXMqZWGfj4UsRqplJqx+gRg
UjyOWkBNPg1laBbdjhSX0R9PtudugT69LV+wwc2Lp4yJH2cuO1S92r6cufhhQz45
F6MLKe989bCIs7VmwfOX5aCF+Z6P9FobNvN9zIcNUVul5QHfbFaJL5B3XPEVLoAv
ChR1EY4JMok8XcWe59c1KQktIbQ9x0xaBqYglucnP1BjI9eqH/yTZHtLauSoljgX
K3yN/iJtbdvaBHqIcy2AKSPxaTrxq84rN+BmgkRJKWQ+l9kCQp7S354+2LauBbYg
2RVUvC0ycbNzv+DsW+5HmL26xxTlPFRvsY1DsygSNk1d6G7/L2iukDLLiNMhRnhY
3fu3GbAmP/uzUrn/1b929KIrWX/uCGaQYAQxsiFcQsR71w6lpwmKUPGmDavX7vcD
aRPvymtdulrz8dMKpxT0KkPKnP4yb9TSn76fd7Bnt31LHNnkE15i5S7EZOyF34b3
jDK/eyyP1ZsKNzuOgJ0DQElB66/n4cWhc81Fy1GLN7vgM/59JKOZeIftwG3m6Vpr
KTLriEw8gj5UNqJYXUeSlBtAwd4sA1GDkZ+ZZcCvDR2RvWMRQIBPDtWo9dZfNHwr
T259Gs8jUmKuKOUpMpMrRob47ywkXL+lO9a3gu8EfnSRGXgcwdPRYxWnaasCNHwQ
fpgBYvXr8UgQRXv6l1GZ6niQNZvlvFd/uGYWcZnTW643s9ktgK6HaDZtDmZFqvMM
+Sb+VA4YAhCNdZA9tj9hOoifeSiqXoSfz281YtB4eRjPwxqIO7/e2CQqfiRnZxyV
SdRKEoAx3Q5LGj4E7kx//+x9NkTKz/nauc8QxCkbIAeRnp9vG5Dvv+0Ro33rgI8x
nHyH3uJKdOGP6ZhRc0L7QetXXRpMatM59OJvYL8E/vK6CDdi9PY3gwh55R10NyAQ
5ms632oglQSEExaXINOtWkM7mZJ0sTwCMlExfEainD2gv4Dhe8f/MdfvY+cTIfHE
reb01d45UY9NHB6m0RHvPqo3D3Y2FVpydHIo2ZR2xIEGsXLCSWRq+QP0EyoTJrzJ
m+ZhqV1n+hD5JFSKFsU5hukf7YKFooKt0DS4FBqkj5uSoQ01peBOSlOOUm51OVI1
0ASnvXvb5p9JaotSZwjwFq5y5HSc5u9eej4W7W3ZKC+TbQ/QO4zlUEvKvxE4TiR6
G83rlssStfRVFzO7AEK8njqWeadBhwgyJrtwC8f6KjfmJubFZV5FsjVzdR28j6AW
pugmOMXq7wZPKwidWHQJwfMG2pwc/c6IhQLLd+QxhYmDuwxLh1rsIdE7Om7kLwKm
gv78EDaBPEqsog67DW2fFXmeVxI8bq5K22BR8F2PyUWkQxwXGHiMR85vHQedAuEe
baml5emfUS+A2LktnAIQucEcaKqrnSTjTvF2KgDcpWtJVRLI/4zJh25HY1PtzGH9
cDf94v1AYaHbApJwesCxGR8FglF4JZnhy02U+fnIDJcZn6eh90dlHbwaVr0nkdYo
ydhHDw7RFg1X1+C2J32XCHCdZr4CYUDGWIGGWlbivC1jNMeW6UWjnQ7KnesIMpxn
7PeZ4h6VR1GzpMWzVXaznKaA7VN9QF80vKL80/mbyu2wAnMSWIMP4SjJMcVyjnrx
wmoy6SBV31EPTc9DO32EEEIULmw1w8DqM9CvUoZp1YT7bA5tKUmuWQIHcv4Gtg22
eyXJK1dyKt8KsZgZFSylOy/Rz0+GA3pDMJQ1c4xiQPa078OL+cfa21jx9UN0IZxt
h4p556zP5sglz1V8Oou0SHjeJyJn+CmY+yLr/I8yyU8AZDP+WTYPr3DzvAYsvrHZ
gSAdxSK+W6f+YMEx0HnrMwPaXhwsQ6ry1tBvBDdnNui/3Gu/MJnjiCcILozQ0FYO
dr9Ku1BWnY5f5TC+nAkjwPyeJ01g+3N61JrHJMPg12xhjyMYU19HnXRG3K0lcXBT
WlW8yG3pvPSYViCPtNpZayxpA2ht2z7X5jGNApE3DJ4D6P9wwr3HquSEvKFQPQNM
V2xIKYeQoAhmhQcjTrPPkQDUtF21OpMwgYx/7xANVWTOIi90Tlv+TiQfmwY2861H
36RjQFca4NNJpPMswvIT6JobK0bAWt5ygG5brPSxofyBIz3KUXka3t/8pEPDBfi5
5qkpvg76e+2j8W5YYoL3fJCcbdw6X7Fx35SCfTQeKfm0bomnmMiS3nBZHMMmMdwn
42aFsoZ9Q61N/T/snoofWe4ENQTxwqRG4Lkm+Fdd0NpT2Wj7n7RgkGK0ty4MYYJf
+Ut//sDwFCqzl1UUpvftQWfm7RCjE3fCGz/qHC7hoGMUz5fIiQ5v7oVV9mTasVPg
VpSeiFeWklryvxH4WDfxdPopY4yLIwwj1P1pTD0anV87xQEhen5ALd1impzVnpTI
nQXyjw52Au2lMMbmgbbEjiYFHYbrr2T6SdwalgDPbWSKFoKqgVeuL6S3qLTsVTa6
4AT3bU5CSVv29YURcswR+aOirC/GqIQK11pJeYD+HEgufuvlSTgaiutAuP54CjfU
0114CPoLNdjuq3MLIrRIskxCSObYDTfBAsf7SDytF05IZsNHfTq5NB2n/XSBM667
0Qb/pZ1gyd/g2c/wQII8zyOgJEPqOuz+J5oHRkmJODUa+1uCF4mQ5vql2k9GMJgF
H9GyLIqJGtOVQPtMgdlqeKp7nyHfI0MCY2HniTxdyU/4uXLKG9aCAN3tKz3w41BB
6iHgeE0uEnT6JcUlir1WNQa+I95O3htxXEk2nfq2POrwbj94UZIyX67p6hfwaHeB
299hKlJQNB7hdRPRZ8PekqlAH722gqaRpSdJS5iNY+oJ8seBYHxMF1BCCCYpKNoY
CK1TMzX3/iyhJpxr+2z0NbJS2EKg+GOIEp9eQAy8phe6T/1vCwptKogZPB18MgJH
qSyQIHC6wtkyDmii8eoTNlEFIxKKQfLMbiIRupqVZrv3aHok0OExn7hy++WLbP0w
X4ao3oh93NQj4jXU6/FaUhmZNtWznwEYaprynUqhuTxMW8Bk8xuNmKdYMmNX/ZQg
Y66+Eu3+cc3pAxVms9M2JxyTazP70NkP11zM+cHitFnQMVgYRz1NQJhPcA2PL2P7
CmfM9xaGZHVjXr3TqMMd0Jey7AzqMGYhqQDCypFwSOHdcq8/5n+4jb1POUZc6c4r
JqUrYytqd+zOc3bguNy7yvPMahVK+gK1VHzLNw0JvVRx8NCeoWp25dJDcOUR66Fn
`pragma protect end_protected
