// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bHqLN7uN8nZsKqm3qw116ncmQhJuWA/GLBaFn7aifJHKFC0FmyoGTl1S1nzzxvJc
raam9j+TFXOQVFrq3Rtvjut4MZhVz15V9SKzXhisKvn/sFpAk/J8ZLW6qr9iNZFM
Ye9Pu1kX67/U/qwUftzCijAYqaRF0KEAwArXOUYZ5bY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4832)
+ONzBjlbHRJ4sdjcMCsHpOGOh/0/SGDDffCDe2ZxqptDqRXyuj8yKQUwbTxOmHLf
Ld8SKuvKAuovbEMg5Qldws8xd0T0tfunWZqeN8LCbYUWT/LZXLcO57yPd0wcmM6S
fAU2Y3S7ngZLuGwLLtT7KsGzJHRGndOWSP4HONvw7r/pYkwgprAvWpbYm6j3suEL
YsgmJxTWKGdCuw2mtn9MHVYZe2N7sSiKWrEnos0LEBSJzKdvqhT4zwhrjePpV/0b
TSviVyQoc12XNz7hxUQvKsogH4bdEHQWgjRPER8tG3TtVE+WHibIEs8aEFUrQ4kR
Ohh2zn1RAqbsU5o779XApw0qzBC9HvF77/ZodqaBJsSjnFfIYtyxsP9gTynwj73a
9/2s+jTat3X2umSnMrzp5uP5BuZbGM8VqymMGHloflfiz+qmCCqppU+Gy60AZWH9
RvFhiM23Hb5YosP6bIV7/HHFuvxZzdmYnvafl+jcfho6C2PZAb//0ExRy2WnWeI9
yF1RDpadVBIWdMf4H/fhdJLHMMLcs34ddVbhzkBFfwMBxMl0ZHJCGO4p6ObKsfSW
R0fSA9MoL/b+e6BC4RTdY58p87dwK3zzgsAnhahYEjqXxAn/QmuexARY7MEDrEzM
XYU4ZiGV1H6nUf0dkZLHpm+DAinHx3OPg9nXAKlArqCYBvT8Uf9HCHQVpg4awhQ4
PV2gczF4PXglOXFBoEPzxZrHqsK6HScPLF22CtD7NTLia9vLC/KAC5ig9lhZZtsz
DYXK6wbzcpWTdx20hshE32XwOez1X8upxoj5d5BOHTFu2TinjJSPyymtRiiQyKHE
a1hhjix96oayswRKxNl+8Q6/MsknJEI7Qlq9RYfCJ6Achm0sqg/CM11KQwLvLwMr
pAwEkJbco+31h0z9hl4sdPH/L9OWuG89fcSJbxr/fiyF7ITe+1b0ukMHP4L4G90g
VL07eCMT6KHtmqPjk4akk09nG0FJjDf2woi2LtXV0eQB4H42uTJoJg0CN66Fimes
oSPtVAC4ig7tp+Ol3GZe2eXMP6sZRCxkuLg10+hS+8nh++Bf2DcypqlZRsEcOwlE
1GoF/WTCjFstHYiQ061xg0lH77sYVroeFBdtiXl3EbMgPAc+x6mVuwl0s7KhJd/C
mBYkWYf19NS43z/RXi9zfA7Q7vFPE00inrlmIy1AsO+ahrmosWcOidWZ1JZh/P2a
vHMUC88lc2zQY8FHmKVxsZWopRSzdfaxpq1XLHhiKyQbkYJcNyBFzTsZmsKMEO86
3DdLlRs1J1/fgPf1I0HoVuGIeSyDVWdd12r/1hJjRXpBxT63pGoL9277mmtntAFU
iQ7M4wEqY4ukBiV+5OhXBUpJtKJhyLN9k3RRMs5DmAVvzq6t3iMUnKXYy2CZVtJc
m1Po802bTCCaKCDzHD+HPmWr6A5+IpH6jdsYwYE7zye3kT9vwJ3/ebCZH3uLf1Bv
bgL8X3u6wvOMnbYwNmSS6CjSzQl0tmnqc+iuNUV6UHX4HDoMOxcbPZNFhCVS6C9p
TSJmfWHEDOyhLk0zjGMEDP5geuolftjHMn+A/b891ATZSAWhOpJZpqHrsNj7zXbu
UVupBAy4VNE/ixvoAwbsWIlmFxHattumHhk08S2wzTSNp/E5dZ/CmwNwRdakugr0
CCo7LU70BpL+igMR1rFe9V/0cURF6GvzgX55fNl+zRfnB0n04ut9qXGABHTLbUFt
DOdaNO2mdtUwxZolT4nlEWFuYwNQT0SvVpmFzb0phLe4COU6J6t0YEu8M8hxfBBP
GIGHBvCW2AzHQ78U0f11DXUgD98c1ZCNAPSrJF5B0RnuJf8+vURK9mTok/rsJIoJ
NZsxmvG/t9ytgYtnkw+4PPccp7iE12qHrO/Y6Z2CYITzQ1W8xH1Wz0Mpsks9kMrc
fSjBtt4qsR94+2ZLzpBIWfBQ3yCv/WLhavJJzeE3nOm/cLGajGoLrhF82pc9CYpu
8nadkivFEQG+kbJ4DEgz0wbhXnBc+ZOTYuD6nk8dZfrngma0B+S2+TR3ALTbwTWC
jR0TkgCTKr4XCWYhRNw7QxzOg8IpYC3286/+Vl5Kb+IwYOBGEPI90P3OU3B7TfWr
02JnRGP4Wbc4EMTAtER/PyL/vMdiuS46ysTUJNqjPDdXw13umhnrsKUdVUMTe7xC
2PbfGKSxIejSCQIJWMc+UDHbDcKPjaH9nGsW9bU20HtJEZqM9V0fK84K4GoV/zCv
0XKzZydS+3bVqOdnVzi1k3S3vUlP7rOcCWbAvcDz0FxrhRWXpm6TmQsNZs2qZWX5
2SP7QqXay0BR4MiGh2f4/+2QGcl3Jb9A5JSxBK50O+XhsTa9/woxmimHtksUiFBt
pivvRA9S1OJsuqYx/pf05IS/0uOI4TOIQ81gnSex+LrbRta1H1vgCnuJ3rUv5OJ9
ehSgDFtmpo8XII55awKeeapbbNFgqZjgammQN0Cq7sWrJ6mL/o9l1WvFmkBqxOsW
A7Ff3EmpcjPBXZYbaXgqZZNSfa625cL46jKBJiUY6mLcJBMa0aJID8wV401QvVyd
Y8qxVv0XGgSiB9LFvBaBsuVz3PGUOBxPuLmwJDaSCeQ90XxjCruCHWFCt5of86l0
2vWXeMGYPLvClnD9Qpg+ei+Ca/bd+WomtTc0HEg47cTUCmMPbI025x7nEFjcmBoo
DSGd8PUVcOUljN4/N5DHZh4sXjeWbxDUvkoymjE9ULG6SNlkBh1WgkjJJifNJrmz
YufFIUJnQw5186mq3RoTt1bEyQWgbL9/PDr2gqSBrGp55DU+E3IiM/4stAYgzDRJ
GkWglvxOnfSZG9U4w2rorWeLScgCYhtHtTtQ6jT//4QA3qtU+znyf4qCUtGqmDAA
3M/yVv4MjRsjUkDSG74IfuQbmE7Mnte1v9P0J86JQA2RQvtVUJ3cBy8YAuBd9NpY
U5QMmcbwbPvSy2rc8gt9SXFW9CEzU3JUxp78g2RbwUQKL5KTvrJ0XGPSWIR9E9vj
N9skhphPLsV9Z3MTdLWr0fnphJIQ8v4Nh8ICAaaeAeLC/zP7rTpcshTjdTqyLiU/
OhsFyF2QUtPMYB14NSDRPZp+aNrV5p6PMwrtY4k4aE269IMpwOYgwF1phnPcBSUd
fEmZycv87nhUzQvio1iiKiWAAjB3zJtWAcWela45jkWLP8GyLvHAx3mIAFduRkD3
klZ/50e4PtEv0+QfC/4LmUQa715cuQTLVp2wS2CMm4WtOc45y4WP7PfRLI6MJW+O
es2uzjScQ5JaJWQicQ3tcHty1wyYEfNMvhShDlS07wuXp90NknUrvnQ77qCCLzmd
qAszZGxh4isUGqLkQ289bzcYBJD/dtfXn9n/NmLQAO9bppp10qK0R3C/Wc4e4NSt
d7CJnpK+riu9x3uT7Xih6mhhsZcFjDN0oAHsO6F14ajFHBMxxKXjtGfkpo+ZheRz
bVzOYs1T3N8TFiBDRHvMPITO1GvKvns0/92uTW17A8fJ0wVFQr66jFJPMn7YkWIF
6W0wgssEwt4rCGJ67MaErd6yx14Dli+tem1hqVaxK/oRhaokx/gw9yI6EX+uJ8iq
jkCY9tsxzOCofjADJ2MY1nN26b/uA/Bh7bHBuT7QaCVqpL7neZPCJ9xsf/YJKxKP
zBQBYsearo04nmt+wLq44SFWctUYlMqXOmpMsn23lifhbHT7/rGFt6RebqDxcvKn
1AWt7Cp2+4QGL2xFuFhX2Qjm3qw51irfc04ecHqrjk23SZL+AvYLxwYy/EOT34+L
DxFiaWk7L6D6gTEwP/bHq2S5837Fg0JgpodaUBlsc+ZXHTcuuSddPgnN5JhYPtnT
SC8hAt2dfr4XTEpe234f5EmlLyHzE5P4RWb8niZrAQEorrQtOx6Xr8FthhtrdkJq
4OZmrFthMMzQJRy3D1Q7fhNgTGP4aMmdGKGW/QFv/y0vgdeY5oGgVG9M2gblDaLm
6wpM4BallBlrxGM1nCASd21w6L4QPYtcEFclShsVaLw/hUXTc/ISpL4ZdhVPAUs+
jc4WKNC2WDXekxhl0NxUT1qNXxXoKJMJjWOirrT19lYtZwmu1IlkP8k/RaBw65XS
fEmGRiWd92Ik/5tY20Mfv7WfAYfgZrJOPQMHG5jBpI2Bf10nJu8/LASZY5BUGIvZ
tWCtgm2VbD74KsIYP+iKsDIZTHqXCsEx8Yl9lrFVYqW/ztzYPDVQiYrUq9pA4NTV
7EmVFA3+9NkPVqmkPFHoI0XWPX40cCMrYTy0KqJ6A89IVzcttA4abXKiNCYPc1xn
CDk1bBMtrxpdiSDeWWMOThbfgifcJTwwA8zHeN8doEhJdDOe8i+uB6jXhsF91cdF
uG3BbDzJPG/g230UrUETOyQxm1B1UJT3GV2pGsnd9DCQIf8isk4+J1tyJeapzwdB
pBO3dRBRfzdaDagUyC4Q0+t5YtKpAFlZKgdJcgYr/1Zho/fu8MQ7nqNKELEZmPxI
EyEydOTYHFgeNmll3brATy+eCmG/c3BEw5kdrgniqPpsEAS+PAzPlTvSJLcsA3pO
ITZQgDjvnwgYreqpleY3CHzhcOTft2THF1mMc7p3tPQJPM7RIiUIyX0DFxAebn5c
3WD7dyLe2hm5+swkyBUV5MSCNuOoQe/hdSfU0qaUIcJUgevEhL6wR1YEzbQiUSDj
H3osyPuInntq+Mj6kVdtisHK7LFMXTdZeuIn15fQmyUtQVVkHQxCa448YuNxyTI8
MzC3ZH7X7M/JepDnhseqno4TArcLwfAyVs9RjtzgFJ4UlneCYRrf0e+XwHQcR9u8
x8e9S3fypf0oLAOeQTyLWmQKWQxtwB2lj5hHE0BMpgzka9oZcnU1VhRI4xyeLwfa
OV3aPuShWRPW9JZEqdUbXWslFzRMz/jdcvpJN4UFiU0af6S4eHL31l8XoyL55D6i
vsZPmGYPCpGDXFX82m3R5FmHEsy5SMuxrXE/AcFqV57LrwdsKgF+Ms1YV0vUmjnd
28741jlag6xzdbY4Xzu8AvL7/XT9fPUyDOkl36NbC8d4jMed2JaI6IDrYDq5T7hy
CfzVvL1Lf5SQX6lx8lOYEExXv/zfkUH1hxX219GMCDcy9LBBB8Yzde05+UPP22sq
zD1Ce4BHlxqEblr5GV8tMgOaXVrPBcAeo7aHu/sUkFeUzz1ZAXxAQvJI0dQzKlCB
HKqiOkgiFkCV9q38riWNiZJOTaaD2GMhW8tLr1Ch1gA4qkF/BxVz/Q99gU+Oh/Fv
TQpEZ3fVnF2xh75+vAYbqEbE+2rxpkrYIOZXY/rpAtZoeP1JuK12TP3lWzsMXItn
l3w+87MdlsIYR23oTZPIyxO63FEf+SvOE0N3u3zhnsrlvu9PKN4haLLduNwf4sUR
lPVW2AlbKUdg5fWixxKfzY1llmXvW+jknY7DfQe/GKdUuNARtQCg4OqKQnC46kDq
70hWZNwFBB9AZHY3lvxzYpq23tk06PDXPKvdsPs2Tg5iz/PhxxMJi9ZTIKbBodGW
tpgeFFBvW0c4rjMEUqPvYIPG9vHWorbdVBXpFB5DIkn/xzAtWbEOjY8vOijDGqWk
HatriWt1tzn9DrX1Dca76r311hKZfnrEIMNTMk0a0oQU6k3BeK5ssEhr0laanmwm
5d844JDgqSiu+3i1Z2LgylXroXumz4taYMSU39ztmgSs5VVGF4xGIJLrHFvWBr4d
Y5vQEIJ1dfVBA0xZQPu7heYPhhk1sXOfIuTRmpRv7t0p4AhO9OadIJsBavL+Qyco
NSF9Q6zOY8dcbp5NdotDj+FT/LlII94IXfS3xPwCCjc7N3491rTeuOI2X6YtTuwe
Z29y44OiJ8QJ19tazhXt3aG378j5TvyWePbaY0SjpeZAwAsg7nnV2IjL30UtRCre
a3NoVSWxRWPaebMxGEEwC0YBoA5OftBBmn9pwMpC/w01EYwngw875Ixj1+To6pFd
Qv44fQfnPfTaz63ZitsK8nPc3ZI/NEN3/bo6QegLYGK3YsKdKoBRvQTXTpCbIsRC
tTWHoVNbPVHvyoeoBTDHvFDafLYaCKgQnCGnQvKwpEYg7YzEjkf1yCH5Ff/MzuqB
AaBYznc1LXl+j14NawzyU5iuaAY5hUp0Fc3lkwxpy4q7J6GKfz/6iCiJqz8HQx/+
5pahVvEND7TAOX0lcbPJALm3t+blx1mhPGwQPfeeGmiSACG/v5NX7n6rdu9nvg8k
OEBv1J7HGNALhZU0yybBu5lIw1X4/0K95/oGhfFXYVs/10NR+BIxhcOUSpJTjUTF
Mt/2gFYj53iS2v1AF19yw9URoKLvEOIg/KNx2jKwUQBEkeTYL8+BK5t8LzGROQ/a
zMG1axV4S81nRHNEzzPF4Jz+yCb2ACOh1dKOcHi6ia/oHIszc+R6qmgmKLQLtqiN
CEWVaytyEyUU6CxFTKacoSoSsZYl0zsLqgk6EUGc4l0=
`pragma protect end_protected
