// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:38 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NJJi/Sv+hJ/lEDMInK5BHw8Qu1b5T0trDinaSRQTIf13mEIigyeGDIhRW6VPhm+o
LIde+MslWQ90vjrJCZbaWRu9/mGcewPVQYJE1YZb+dxCwbMBVrZlGewECbKYrL/P
Q9katEP1xHNfb/0QZC4vPWt3TAhhpwm01/wH5Zkdx30=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19056)
BMLx3Uxm0QCGsoJazvo802Xb6Rr1WFbVF9iFnGQOFEnpWbsPA6X5zFOtnRbXSRYO
I/2aGMqMJw/WC50eszOWIuPRJFAxJZcRQcGON19OBxlVZytqiEB8KlD+8vr1g3W5
rchspnWFJZbEq4j0P+cqWqctgcY+yvzQfWNIuAOazNXINNQJgHwn/w6FJxmnajDL
bqhHP5sHub3rRl9JEj4wIWDzoTieFcMDHw7tM88RD0iTcthwbxeAosg4awv697rr
EUx4OYCHxMyds9z7L30AdWzU2R/Uk7BgIXQXgaCBeHbrmct0Oyz2MJVH3HYbisGy
pngaKv2Zas0m4yM9zt/50GRGt/hDzmLpqxUO0IVoTDzQRgwe3gs3H0L3FzUKg0uH
nwGDkvUf9SnqJnZbRTKxL3EIa55/DZMlzY/Hqp6X8rXtlf9YNUIkmfX7byMt4JZ2
JbyNFDZyCSo7ljkyCGxAL/6waysD3e5rn1s0TiqZsddsAyCc55xiM50eE7Lq7qbL
LH/LXwNEA+7SFDNWZqbPydnvGPL9Ubcbj0L3Fh0/AgSwY2GCVPxOUrT/rgAMSdy9
CBMmQtwrS/1irXbU6zHqRZMGQ5f3G1NGx7zRdAP4kD0LImUeRCL48nS7grPsCMJJ
HLpF38Rhp8j5PJ3X+EVXDznaq+BhoI0JhxxiCsFbUKAHp7ey682EGZ7b5UlUI75s
ZQ5ANoJuFsbdUrdyxJZH86JOVdGZ5hG23RGFuEBxOpYFukqarPJD1luKKReYXZhG
J7J6SdghNrrGukV2R9L3ahzFbHNxJf4pjL7UG2wyl/mqs44FjyqPvK5QJOnrYRyI
fKj3IjnLH4qGTbrZZeubCOJNlALeoaiinufdH7uXapWxw76NzCOkvSBoDC/+9w7f
n5DPaWlzmUeRN967KIo06WfBmkw7T1Jnnr5TwpU9AY7zR3mLdrm3Asi26pnuKDty
pgBVBt3Wa8x7303nROWOWQPdrNt2N+4ZrlPArwrJNq/eenKMB/i/Wf3ou2PWNbAY
VkY16vfrxpiEEM8bp80c5DbBRa+OS8pGQqlN95ZFDMxqwyExL4FFjpgv4KrFKKR5
KLIg5f88En6bQPnxl57swWfSMXFGXnEAUccWyu3x91cwo8IQtUeMvflFv3wbcUZR
lVm8fKZMtIeqddWKEOcH8b37KQ/PpChj7TQaFU1ibYJK0On+xFn+SnrptJ46yzSv
bCYQaiyPOD2LnFgCGMbEEI9UL7ACVVuz4C7367maK2esBy81e3HqkuY/6SYpxk/W
vmi8r81PUDLxdehdfmUSkLL+Y8DyAIy0wwHxj/uUs61d2uKm8VQzoBl1TGOeIugF
6V+bD0Ur9//hJllPKM5Qu7JhVAS9FuD859ap0z4sNOQmMFv030XuY6dEggDDXDX5
tcs9Xp5mdLP1AdpbBmYhgSKZr2D8oo3cgEUG+rrYcRPty0l7doSmBGCAwHKY+ByX
bk/gzXIWw77G4y/RpWA7xqH+HoEYq6l4OgStWs89+RR95dF02cLCEHzxrxJ/Z9Nv
ofmNkpBRdAIJqAp2DwmTT7z2Bop8WtZWmrLSZZzGOFBukEVJ+CE2eB1RY8a47gmS
3hGgQl94uiWIHwPk6xHimsoiAVdgbbyU1IgLL1jrjZJeSUoIJPEe2ZZXR4Uc+qpE
QNsJqDZexCo15uvw2MuKruTw/6eQE17VIAsjxfvwdP5prkFwmlJDJnZB87idH98U
qSgg91ytIV45udb6brdNCXnaLyEUPvX/cTneEp2chIQbzpmjwtSimxD/viZYLhnw
SdlzACq5PqqNm6lDNutNwzSsr3KfADZDPrmBplIxnKRSqo9vs/fvXocbkRunfPrC
NPO1Cwke6PvyXHjdW6o12gi5yKlLJO+eX8zeB2EJBY4hnZfybsiQQiCgnJ3/bNPE
JlMP+H3yE1Wv6xznx+JikoidW1gaBssm5sBO2iBykbEXxQULa136FH0esR4YOWwS
Tihqs9b1bd8LIY88xJ1XSaJAEp/rpAGY6y1KpujvAdxT8lYIiqRRpTe5nvCjCvSH
derqMH+XPBYHRJR/ji5WE+WpRmbrtU9Dn7CM3Erah7lN6h6oHlYSof9bK38Ldju/
qTd6yf4OoW1lMCJo7EzxabdTTaBULOQ+HC3CN9j6LLRfhk/7cG+ed/NcTK+sV/dH
9RVwWrecPkO4eszmQ11iZm0EebkDXOb4IIbY6bmSMguybZ500pG+GUU3nHyZTzkA
w0ls/0ExDa0v0vKIVS9y6WdAYz+L7rq+eZRZb9ebP4G2xJf8BFi+ui7vVNQDBitP
ugPlVIxB9gcHj2EDGxPHIXaewNc4CuNCj3hX0aJPi6EaFLvaxMng1dNYz3CgzulK
M1MPFWP/TK612QRfzObkC19aFqbZFYmOOmr9eEj4bHakNdu+qv3/ymQWyhBhtaL/
xXraAkMPkXFKp/KV5N0tdajiK+cHkO2elM80Um84jw1mxXaPBy7HX8tvesat3QGV
gSnb5AkaSo5SyN3Z1e2kjSL4mUV2OMzb69/vF77UNDLOfEi8aUMDwEbm7T8jvPYZ
YlR75z5kbRSuDEgXCw7eKvZRC6T1tn3NZ6xkQexE9cMoAXGtx0DEveA6jNPl8Lke
yW09K33iVDOHk2kwR9QNh6Y19BprTtkg9kQhD8V27pclvIaZv9Scwmo0VM2+WyDE
UVkJuTV171xxBc5Dd3EWtFnwq7OsqPNCyOCMETKH1zZLuqGvT7zGRPJyyuGS6YVR
gGVqHmt5XxC/31vSoKcY83Ui57GbExLcHKbp/xHwGboj5OczlR+f3fGuwlvSU/+Z
adhO4Y9nmVuoz+yx+qHktwH9sRg9x6ZNMkowgT4RbKxtVfWK4AoDnkImi+iAfyUN
ZxGWY+6QyjULoSHtm4WyvQ6Tby7yx9N8zecnHZ+hLFS7n5eizpaFC2BsAEmtq++I
nP63SvPuNAzFvtYQI0uo5Qq5z8BqLGAHSPbj3lQkkyP8VF+D9w3VG9mYGXURJjjB
a+3SNCMA9+EMTQBkfmxAA7ceHbmAfixBiUaFw4owL4d2oMD+JuSFWo3tH+qhHh7X
yAga0b/AfH0D+rLGqdQuPvosh8zI2oCpVcO+kdAiiI20Qxg0n4MYdYS6KadQ2GmR
Zyj3/feG7dlLyQ010fW5M4z74G+UuGWRkyCp+rG3dLSBVAYbuiylqm7nY30sffVw
yHON02DEdHzVvntTw2Z5PSLuoCahmt4tV3K2hEn5PxBVEXmvWTREAZiEDNgXDJXo
OtOMhEQ2+T7T1jE1cIG87YLllkCN/3yRIdStsW2GOyA5o3/I1f63x3U1dDDohd8y
KQvRBBjsS3qTXB9657MehcfeoadodD2/gzcg+p8EFC27e1/ndVZRW4MCyDlRkcsW
fPhMCqhBopvQfj3iTAcyxHPjSkaALl7+LAulExdZVudkqFTuV0g5xvyhYeHHoQJ+
6oDUy625cPPPpnq0JzxftM1794B0AN9Si0OqctHBIbGZBbDYqUKS38lD+NO9fK73
et2qkrzJnDa0vy+dH0JC/Y+L11KtAQHbD5cMq9RKgOBB0x296H1nro/1JC94VZcJ
n4KL91QrWcJ359hrAX71MFruizmU0iI3JHf4/4+NR2hPFjggZ1k4Mt4EYUzFUqrE
TOpGE4QAvuVDJJUgDPBn9bRVX2t7GmouNLRGTwcl3uDKVCWy306+VngWJUP46NVu
AVEfgsXRMOGZF8Oqxhs61vyiOMGPdIavLSK6RoxGeA7NVTNWpy4QnlHbpW1TS9mu
J/OwBE4x+N+dkchjERCE+ycsl5dncHQ9sNqZUGEZRMhu8YLx75tQMA3FUbxxYnVi
iYGy2odBDB1My56ap7TbWqvNi8YbQXmMr9c/ORFFuyZmXAkZmoOk/Jrybw+PR5Nt
Qflh3JGu491ccWSsfi45jO/2DSqYcqEdVMd9glyGO/WIy32T0SWO7bOLJeHKYp/H
Y3kEIWCjmT3V2vIKCnVCw48HRlOGu1a0p3+32WTY1Ns1BEpQ3t2Q1FpyXGMiXGgK
TXObDM63dT3v9CEr7WKOL+evHxyXKlBQMtFG9hoTOc+bH4VKg7y3Cc4NfqKMSmTA
P9xlI6UWjhXFICiUrLD1OTMfzeCFCGAXDVZ7wsPA9E157EmnfcdYEfb8VJ1B+4tj
pJ65X8MtgVNrCzcRiO31msoirifS+5Kzt7RJEFi2bZ24+lGGeBy78laXExzCBl2f
uzB40k3/bX9YmrG51CvMDzpQ0XjBc7CpFkzx4BbiIaqwrhJysBRyz1AgQ7AWfnr5
yyeZWL3sNqNC+J3UzAIIZEx9AgzWxnavs+I776klK5aL3BF+urPA9E+iOKDC7UW1
ilIQzmbH2CxX9CElrzPAHvCBysUvfmS7hhfxGA9XQwtHWpAaPNq2HZ7IurBI0P9Z
j5IbfjGr/SztGvXOBp8dBY/0qaF0nO0Y+sd9/5vpEEHXz1CRot25dMR1/9cCb95n
0cN8emHSWgqh/693hpGWE0eREwcWQ+N7E6XVriWgYz/hv5eZVzwks8S76precK+c
jh7pFCkOsHVRoBoFT5T3dMeI3+TO67MQnNemE/9ylZYR058NK79KV1tpcKtA9/wu
Ks69z2GgfBGIerfjNNA2J5SlzFiI1nm9/df9UNM+WHGiL0eNKnXTYDp59lxFEhms
9+3/uNPl8Hn20y2cjvbzgF9AV6V2pxY8QXIxMiR/UnkUMM+l0gvj/3ch6ta+wA+F
IKgy+Grgiz8Lgxx1s7bDGegLbvro2lSmD8njOzCXgM7AYQel1Q522r9opaq+CFgX
lDU2k2DyXypKfN83oXzL3o02kdPmTFjWIwCXg3qameYGbL25L/eF3L1nGij4hbS5
03T330vIgEoAfg6gtUGnhkNMuADicQ5AaOdrpLS5xLSjj/XqZgPqomkMY9gYu6ot
tw13aSwzJ2I+RP2a0f91Pqo7rUID1xPjvfkxP76OhCRnUOKwKe/AmoBOmaYOU/e4
ryf73aKSlOv9Y1z6bg5Wbygdzn9U6b/av4/8n598xL5tM/NtNMlrq/VZrzFyf/0x
pJp03ip+Yxq/ieGG93Sz1XFCPUBTt3ZbWj067szLTk72RB0GDyR69EpuwvfarzHE
o3RKXJEJuQH2y9T+6KjMJVbrKmPf9pC7wq8fOY3WIZBij3CRNQSgTaGAIfQ7iqS4
gkwr6ZZv9n108b6JX3X/twfAIdmO8wr0GcRy80wTPscTe7bnXzytaZh0ueE1fHU9
wYO6c81T1NnqP3G7f8kSrxB1y/oU4LmV8BmsBSuwyL/wn0XmMuAkhF24ddCpfFok
2m7d8ngUAlB4kwGMzyIrHZyuSYknhyYL9ttZhxjglyJZY9Xv4zRoIXw69QfQ+KY6
DbLVaKwgncq+t3E0Iy8CatmLTepLVM5lkmgPnX5Mr/mG7YA/srFca4v4h8DVKfcm
gCLKqE4r0+PvOJpgM5S4mUU9KC3LOr/uEnQTOGi7pBqjEje6vGFkqeBjT2aB0zLW
Pno9TztAftSuNL0yjn0gf9M7lbO88JQzqPMbTUh0EY5pzN8vj5DuMbg+zEQeLXRC
eVBO//vPJ72si/HC8mGir134DDlYJw77pjTJrjoP5GGRx+193FbyGNA4OV+q9DqL
fli1r7zuM9isYTVjWOalHNX+jCAL3dzVgII7zJUrHOHuGqg0sW5txlfJRm+kBXIP
wsWNzXDBMOiIFqGMYHOyofL6LF1JvWUxF16qIKPcAsdQkJi5cI6351qFVdWdCML0
wKIciAgYnKGA3T+316WhvUskJMxykq5zdE9KcPepce4yL2+Dgx7ewFnU5UOG7lBI
noduW97PH9PIfRz1DAr3/Nvv9kjMJd0S10G18Jm2nA9NMpUkaTNJ71SldmfCu341
YKzM/C6gPD83klTp/pUhmKp6Wl87lkRqPZCnb4+vjtov0EY4wqwQ8g8SRya48TRe
sGkm9XmB6o3fNpdk5Fe1QK2kOFTNbRE5RgdRMXGrmFNCTQ+ZNypVAWJ/AfEHfSkj
/ShpVnThXsV8N7jl8XJVwhlaw1iSKvu6h15DCbW1qDfAz7Q9ITNSvxsRFEIrkv/+
nTLu4dpxuxSm+g2n8xI3waKkl0X3/TBIou59wSDwmAUbVl0EG36zLe/t7VzxihEd
6rcKhzNzXjFGPMPCJH2YgNWjlmNm8uE8rC++sAq8HkzBmF5MAy2y7va72IwouYKj
g6rAlSMc3JG1Akok8bX6jivQUmWN7S42nJnetn5s+8ctCFTyyCtdQUtQoD+g2kWW
GqqYYeSsxeRlcxGKbxl2ELFkc8fx/QQrhHgkyPOjh1zbTU1xc/xJ01PDLU8KjeGS
z93DpHm9295UN4S1TuvUgSMtUnJsx10aOx7tkHVsutrL7KG3NfeHFQiPO5OLwMuY
TwyREt8zT/4ScWT0Z/wvsm/JUnr9b4Pw0arRXi3zpmheSuIHUE5JqCAeSeqyrUVx
VVNFw3+4kneicgl2cuD0JLAltZLUZr9uZEE0Dp89+PAwgkKweYFG9kY3W+6LL49B
+Bb780DKdbNajO5BWe7BmjCLGeYQITG2qL3cBzYU5Nk0SWbz1UaizhnDXz2u4hXA
6Vcui28RexTWrtqFt9+RahJteiGsCOKFyIZHenMZ2TZHOjOIDKFMYpmF+Pqpqi42
XY04uX+vitpExcI7DpPN73GHqT+nUzB+usbmh4hbMaIS9ZR+IdvV/A35LrUmB52p
NsMwrQIsVxsv/gazoCEZ54eyzLg2HL//XnMhCYX5jjivpPxJq1o5hyktcQiv3WX2
Vs4zK1Usd30J2suN26BBA6HvVdxS8yWi3ydF+O1zR5YnMVNXewYjPjSWr+UHJ9PG
kJgz+YVd7fOpYoG9iqE89UzRFbAl/WuQGSIHQS831fIv9XD5fZNxsbj/gcLj8a8y
+cx84VdO9fiHDpdWAONzhzAZzK7thm907t5n/+fj1YppLjAu5wP1IyJspKnvZZPO
YE6vErtlmmgGdd85BFfeYnwYwY1/V/vv7N80BCcvCegAmNkjoiyT1Rytyy/7pZpJ
iNseVEyGe3/j/2TdnSM/RSrZDCpOVUpEBxFfI8tS/krYZsTHWv5qGD9BQD5dwiLQ
z/YufG8wy9XhKeLk1YX6R3N3zR/k9EpjoDQorI9dF5MJD4TIg3qG0GdS+tl2xrPM
JnXIBoISHjlnc6+SXpQAB8EQ71frAf4GThLYf6gTRGacI7Yeg8wCvRLthmKnzbPN
ObRTkhTl1Q0FPcbpmOhowyrinuRNw1c0h4VWqFd7WSpdWLhUmkAAbYcCd92FEZII
ubPbl8mUOAsFQ4XVPkQJw4HTYXN3jshV3dzMzQVohWrRu9XaP1UkcI1K0bRPuVL4
F//6w2ly5ImF9XzYs7nQFyqABPQf4W9rUmC+l8GDHDV4ao2qVvhYSXEUpLwldVb/
kymHsuDnO+KJR5TPX3If29chxsIN3IgNEmQawpVRnIg6FJ55u5oHUN546XSEPvAk
K4b7UbkqaVStjoMepFM8Wvw4VT6Nmfj5MHJUDCpVqxPjBMVn2wl0udnbDcQraJiT
0utvAxUPDnauRv7RtZMI6XfuaBrugT1+CMhFdvPPXkcGWaYHiRANu7eOuloYGvP6
86zmTxDFsCxjE5VoGumDGGAw9EHFrjQxdtTMv+KvtUqwzGLSV7RdCFuWAGlYnK10
AZzJOn99e1gX1l+79RaYdqQTghcRqSYt7UEYIvpo6WXrmkyFryoOMuos3qDvz0af
6XK9i5xSZrIyowqN1WUewADVgcwCqqV4woOO/+UR5yefMBIfP4PlX23TH0hUHci1
bIR+AYLUg5e2GgY/ypWlBwEeE9UkUYD8L+mqiTlaH1HQf6KgYCU6YKSApOSLUUGF
lamwuR6eyhnfHi7a9HXBg+QOBvgTkEnUAf5hPMrXJKhVj1RXRsVCstBwG8TtSeuF
PWUgDnyR7cbofRIQImUKSnEq5SAgxYoZocScE4u3rkwqp2HWz4h4DyTOFvXi6htr
Uz1L/9Z8IO++xyFdjQYzbUI6DyVfaaRV64f9lGPCvGqQDIEExjP1clukPg2zXJan
cd9vfYFmy6weZyG7de+D9mNNWSSAAxu3RvjIbKvhbh0508Zy+ZV8MKh6C5Roev2e
8YzVvnSf/WalOTGAIfPbOoilwZ6aQ7gFGBKuf1JM1JRulixzRWOs9mYEC081/72M
WqxPeT7Og9PV0YheXVbXk5oJkzLdPcvbguUTOyBo9TS6itEFhOfBOBTrApMWgvzd
uhNugHGhTDgN0ht7yHj9btiw2RUCuGp4EVzo1DxgTGitfqb5V70337N5V6XgiKPC
1oVaLvJvKrp8uJpW40hjvxx7CQgx2lU3guOTcvEFDcfNm6anRFn1YaSbxOqQCRWe
ayEiUxgtT8kjVLWvhh8aT0pOE3PrF1MAvN9Jd7ZYIMlxZQ5M56cqfig+jRxTKi6Y
eN8aqNrHp9zW7zNHaKnCQr9DdHVBL/QPZaEtYsiJWfZHJYAWeE/R5vEnDgnRsfng
YDtgvHz90LmtoU8Qz3haoLg2rsvw/GeVBrBkp0LETwdt+9jNXmHuS2fBe7PbcovB
O6ILZPJvT0jhxkuikfZr9aC1Q0af/aDqvTx4C5KTVJV6eU20RU8UdVpAuqnmwbFB
WD2OyMxrARff5qhgJUzerjsFgZGMDR0gaZLPryNnLqBdEKclKdoqq/1y99sv49+M
yP3zBuAW/8gy0BD2oOlScNzcozQYU6ymFR4pRnfcK/TzkAA2Y7BBk7GucKjrqm1v
ajWHtJVVaKob7KgUB7YH+TmryYLHELVXD7ceATdmUIXqiiq4QVyN8odDAAVRi7jH
wE50/oLM+N5E//2A2fAJqlDSaEcDrEPVQ3+gRd7Eoa3PfcaOmbwQEeD1AC+o7erv
nrCMaEQ8MLBsb2h2sFJ4Ph4kCO2t7xw7WYTGUnPRaEGui45nOxC2XGwqNfAXnXVw
4xkKV6QXJaXOUhP8Et3sSAe3XDEFaRBhAd6GpeFUFGFbEp67W/xlKq5voTbms9+v
vBv2mbZ/pL54pYfU0iF62oSHKgkm4jV50wK+Eyp5WLUgjBgd/8Ck1J+pObUh1kU5
zE1G7rsur/yOZsTwpt+mYONSTkc3lzrUpQE5no8VY1Vl9eLxB6qMK/GNNuJCGAjn
zEdRmIGHMIP6Wp5EcFLKRaIDCTIF8CZ6aJBLZSbM1yNm2hrsESkR3A8EEOhWtBVr
/g+9hoFinonz1OJnycMWeavVdUNy6Iz1T2KlyaXXVFQNjSibfWtxwwcx89QBREcw
pwS0MZU/E+vfKGU1cfZ2JLFCv8xzwU74rg1JVAa9jx5a2L6mfGR6+FmWjd+IW+IY
UxlRIh0dfFwFPIbnh5ysmmM0yoDnOCfHKRg3uG/vYxbTL5YSFcm2GAaGfLbl76N1
Xh17fxyKcWB7YufAw/GOAZXJihQMnZTK+ZT2p143HVqhxx3bE2aKhezFtv9yZndP
njEHMsPk518hP3bL/F+6k35eMat+rmQIbtqlNp4b9Bg8y2hsvNTS0sT+qCabFp+H
t2D2wmstkdtLak8czEE0f6k7m/6bNGf5V3xgYq7Bo9Kkjqw4W2ZKykFTM/VpoE1/
gM5aCQc4UTwkptFmJblH13yebiLQLf6Lu3q4qEuV4oAphpruSyorLI5ZlKPTydwj
eYIX74AsSS94X/oPOmROYyoCgpC6Ii9v1+dyclr2XHQn48VluZM+xHU6FZP4zgMy
dEiJ3QdauyQZuMy2GZtpMuN9Be2cHpeJrssQ/G5/rhyhisKr5nHSAvXUR0jogWiV
qxrGPsbzvJKWPn++I/PPFCxPFYGmlTtFSP/1YeSz4HsrLpqR57Y9vLb1VsDhme2Y
ib6kfU1l2JPtN1XWZkWt2oN4C6QSgbJ6dx0erO+3qyXzT6MvSs8cxUclkwEDOBqM
XWNaSracziqKybS314gCTz0qOTO4zNjHO9ZJil1+CathOokoah5PWw2wpe6jzOr1
ZKqkNQ7+/lNZdH/K+3Vi2rsQmOHdZvYlrjcuM8wOsMteW0GWBZVwOnb8qgW8rth9
enbaRYh1XI3yC24WkYDp+HsQsIQ6XDj6Zp9B+IPA0CyhfQtrRuhDScI4VOReTtFk
2RgRrAnzo8HPfr9ZptOoRBc0isTuiSVoTHkshgKYLjev1AYkD42Kb1HWddh3mFqF
D7rd82fltWYR2vsE4pAHj30F+XujqFK7faDHWWD5sm9fEWFaO/xvUr/DwW3BwX90
QE+jqxgiQuTxy3WkqFbpGYfEQ0Vz+nwyPdB3TFKgtCLRerSQ9v+rrfGxaR1UvgCv
8bJ4az6+VZKAwphenD2luXksb5N2hiPD9+4Wlk5UwWO6fZzM6ecBqZa8gEKLC5Nz
yZtJm0SbtGeTeGJwShlFWCOlgFcSzT2WcwOPdgCOyuAPgdzHDqOhspYgQfJL55XJ
vwBas4xMuxO6/rTLa3bAscjTvI/gc4V+8nD+LkH5tj8zYyCLqYKU7ST+L36B54Np
Kjm7ubhGyX9oo/UxzDKk/v3vnl8/QZaP8DRiIuf4Yt0KA2FuWYHPZYoMJnEacXEt
+gIryEoDHRK4tDM/y4e/uVgTIwU9dTk7xn3zsJM+JUBCODp4OG6mkKeLhcmTJjqz
Wwt/FkuvBkUsUMBVTiXqKIHHsOxGweK9CtafU/oMQe97LtH+p30sM+BbR6rx5qXI
XcXj8e/yGHgKGTjT6lb3m/xwlX2o5Q/rzonWt3bTbUNkiwYS6hKCf2SUSXz+/UDF
WiZkVcV14/23MzKW8SQu4A9BuaRcftk4IQmy5DrZ6J9WCbXyGm7Ljy5F26q4hbfO
5gPsHTHMPNbineIrPREpF2PPD/aGdp7nX44pkRrlD4icBu1UacQHslC23XR88/Xt
KxTipWqacu6Jmy7nvx9ZBMmYC+6SVr5qJReZ5MezLhzZXA2rFAAtBR8mS7zR7sQo
bp2SCuU0mbcTyd2Irl8rW7oHmDpOWl+i+BmiQbykmrq/eidA9PA3Kq4TDrpicyvA
9C64VPes/EZzLiCVtFXqtc+Tbq6ar0qcWz2sD3A5iJBEmr5y8LORKODyiRJBqczS
G2ujcI7mF5s9+0O1sKZjVrl6klmxyJzDqJzXH6YkDIDnFl1Rh0e1J/JDE6Ozct7l
oWQU4uu9ztPT22Lj23LUiP1lLy6uMhyT5QEoQ3igk2MrYzO/Qc2Qr31r/MHwA19M
h7bf6XrJbdihFYupLIVGa3cT0PsGP34MSRdwf44CgyL4psZkCGOrdZix7DNaTazy
9LCV1An3QYwKcrST2x8DtQ1HSmJTPFVILSiaWsKhiqG1p9c7auH5/cAFe7yZ53/E
yG4NwaePMIPHI8qHIz1mvfMAWm68r5wgT78cXf1Y1Yb+U8Oh10oBMAMfCf/1WcEe
WUSs49q+sBtQDqHnE0Lenw5VSIBBovu4tq/U6Ofo1CCr3DJ89EpyT2ZBHevAa2tE
x4Z7fF7inprcs25JnCWlb/RKiMUbvMdnnnfeG2esVmS/h5und7Mbcghw5FDyccuM
pds9ghUU1wX608+UDbfgFFRyQVUyDJ5KQ1ObYtjdR7jib+VwsHJnwh3pMsm7abzN
jjnub9tDucSdEgksTg6QJzT5qby2PpcM3cht0h70jve7fhAIbM1wmTXQ04ZdavYH
V1N7RCpu+Uf40D587BjjjiUL81TJ6EW4NBVyXLvFMKpVRFlfxz9nwARcbCSl1HmQ
i3pe4Z1fcHobWu8pw3Qr4aW95B3k8baUPtguU1GH4YIzELWgnyPDwTXwXQUWU/iD
G0uzl0rlV7ophGGPFqBRFm0VYresptRW793gRVFhqMV5oEih/h52yKkMKaSQq9l/
dFaXc/JPy7b0Gc9qCsNuwO8A8Ewt71TcenLPNWG3pWjuBnIK9W/ZrPAaO8FBzbVo
EgQUVGRg9aOC/ouZMKlPIAq324xo0NfElXB/CvqIE3STLgBBM2jVOemZIBm7TAkp
i2qeGlyH5vdzD3jKv6NHVJ0CKYprKtHK7XRTiw2gCvlyLSIiWQR2KUBrz80HzO8x
YUfdkURE0IMAFTg3gb4PABJY9EUideyPhDRiT17kM5YqfYqvnmrWz0FHnXhafHRa
7zAKV7WDHeEbejKRyZq+VaVh84SijNsdVpZxa2TFOx8Z8V6oAHnBG1c+dP7jgIoB
Rf627jYkQmaLxpl946E3n0gopq5ZuudtRYqdpu2wsb04vMvYqDyatxTML6Lcakj0
IrGtuwT4JdfDkRrNFzYgHvWkhTX2KmgJ3P+HmzfU6fgxm85p9a0TWR//s1UXXn+5
HZUSh+RXsBjL2F7aoZmX9xSb1Jc0BpydzuNvhMtQ1rKz3TGAx9cFHsvfO4HURaEU
6eEvxAavfX9tmfkrWOThTLtgeojw/QIzNB2KLXr9MJnVpIbklW28XT++SUbvjUYo
BS2m5cbeXa687RL8y6PWaF7wWglGUsp5kVfLIt3Ne0qjpAdU1+TS2TqpxE/Vuyxy
F2D00k6uGobN+WxsOr5TAW4j19GrQWClbBnlacvydBUTEXSSiGk33JRJvdNwssAe
z9GS78dNViegvhI3fjuTdD1DlWVu+AL9Rms/vdlCMnuYiEtDLl+uX7VSjh+wNJU3
+dyD/hIiFuj65noMvqtKrZKyM47Zc4do5JXCTR3+VQtzsefk9+n5DSyq2xokK+xL
GyhVMYsKKYYRtznupFJ46lMG8sMWry08xLymj+mlxD1VJhA6hUogyiKriNGwqFwG
XyCrZqcsl8l5JKs8iaNkb7STS5teKS5tLph3/8VYmBBIbU6JA+H07xeUQgZAJ6Uv
aoBnawVnj7czDP1e9ZkveOebJDUzIzRrsH2oLIWBo0/ev0hGWndCRE+3zrbqB+ql
FyvylSzDNb2OPD/WPzpxuOcCp6q+7aJ8SBe9VGMJVtqfZrL6scVt/k5b0mFoBy6B
z/bIcu36qKUraYC5J2Xp1ro/2jo6HfEsB4v1rpJiHfnv45r8TrjdxucillEtdhYg
9oZ6NyGXLc6RuTf/icoWOcQm1lrnsgQ1dVDJmI+pAQCoZOuq1n0whPHRQmEICM6y
qUBGSfg0EcAjOz+fm9bE3qQN5T//fVrI399thMMYdzhlLjSvhcu3bzL++QClPhp/
FAwiq6sAlRpWAh92LU6XILoLPda6086EIyDKBzqgEQIsiJikhzgqspKp9nfBzriB
9i8Z3HGU5opyCW01biLebGTgYyyU4CnzGiz9D87YzdFrioQQhLlgVPadfqWQ9Zfw
BFC27RwxlcDtULS8pZX5xOIvrzW8cJBJuW33wM92VHnFcdfpatMA2mK/9dPFxSGV
GKLyrlqh7u5+JEOIUSESUnmaltEBGrNyH8LE+DhjLR7101BzBjajETAcPK8wArhn
u4YGwHlsScRkPwR75WN7nIfVB+/l48nGILdJPlaYJiiSh52euffFEV7gcY/n/5MP
tUYs4KXA+I35RaUXW8vAY5SHDh/5AsN0AwS411V9PJjjpYUZtc4xMMmnVIoo7Xgv
tXKMo0WZ2zfm3RoOtuyNjReGObu9fIAGrKQKUi3BtTc1KqR3pasoTq1QJ883Qhrl
jwbwZSZEpzGbMl9IqIZppwxVQ+roEC6F/h7O3vF63JHSTz0WWGvqXv2YLl2sRlyx
X6yYedPfVvfMKmyjJldq3sUSGEfUZbKYILm0EmT6U/pBsa/Ex5cMa3Pcjw55h8hX
oHSFOOkTsvL4panqVkOfb/TV4heOZ1J2oyTcpPXExG9d7NIVs9Z4CaEs+8s/+hl6
TjJ4nc5vec56Am3sdvcsPbzIyG0T2NRYfL35yxH1fPMS/tfwT2SSIn4LRb0zyVxT
+Zn6FjhcmrsAc5rZcTWkClLI8uah+2YLOIVrcCN5Vm4+Pk4gokgE+K1I0NKGoGeX
HdT/2GNZKFRR65G1pccqFz7MldNhbaqJFEeATxDI1roQZ3j63F0Aj9V1IsRx3+bR
LJ7Cg6PavkAl+FDlwp7RABCKWdLkFOKXslNQ2YeraiwhRfnLXzGTD4YWvzkNhPAR
JGrPV0hUgtfXZLMfCkKfV7RGEpfb0yPeFgLoTxo6kITrxooxRGcbROkjLlJCin0y
RBaLvuWj1/ml71xafF1bX+fFBx4yDyuCJfQ4+AxmKkB2pW3falQEq6DjeqGIDhK3
v3xBqDXdsxsjFvCPn4sYWoea50DdZZPAxJ9KyeUy8jfetxTZ9G43MX7mI+/H3tGa
Tqdn3VEYAfEMoDAxrhxkid6qqYUj/9mEfqytqXp1B8fYsO7FPQIQyIXaJlzJKmTn
Wxu7t67TexObdVlkA4aUcpKa0e4tb2HoiaV0hL13qul/X6MSCCk4UrFiBe3EcZc4
l7Sbb8OV4dvBcCmOJqpkzXJlvhiNNI3Y0gUVbG+aJBYka5CwUm8tT5ijRf2fbpRc
G3qOI6NkaHBwFje/76xyAM8SXavYeleshq/VfDmnNR+hQaSFf8gfmXgeFuJqCehb
rR2SAJDNxYC4V9XkGyJHWxopx4uoLPPBg3LozGkZTgArVn/dqfEPQzLXJ/ovEzuo
mGoOsklfWsyfG2qo+owPfsrAfSwHcUVkc6PL8LstIQHHsACOy3wRze0oMUjweFV/
Ee7SOh9OPSnjFajZXeyJcRBR7nAHqimQwIvgHlqo3wjTB6IWDTc+dw4ie6LSL5c+
iLNOVfRJzVkSuEFOrf6i0Yh0LiPhdCXIKkW1376x9Ef3ez7vosN606ehGh5ho09k
l21ToY7YqZf2kpBZt/I1oRjvWx1brOjH8TNbvreYhni2V0B+rN3fWYcyNFr5Lp8R
jUWpvosJVXgAa+uVEjmhNuWjFxvqpHBH+kwg5MjuhgCl+woxbYaCFQ1iaCS2zs0I
aaKXAiJB9CEER0fe7TZvcEW6Zotn5Z7GSzZKQ1NZLNpcvkIi+c1eWYOTNXRdPTB4
LFM5DQtTukLFaccxVyjmHEu20IdJkqXsnYLMqIg1jn/GPlS8XuhQvYnPIHXqHvkT
YnQT4BSmemQBro1b3sxByZdZhQxOyuKGQ+y1Okccj43TS/8Rl+vc4/Ff8iyjx3yV
wFMtGZsNOIjZKlikAxJOEg5le/BIfw4/mGgUEXhiMgQMH/aDImdBqZ97UkHdV+4a
jwAfrTS/zQGFyIECw8BeSiW3OgZ7f7CdjzbtE9XFT9y8w9ooBO/jm4IE3EsG/RfX
ZxK1EoFkUieWOwufGwnNcT3xV579mKo5EnfQK6qRUqmcMvGZytqXIuH0N2B3E9D3
Lqja+FCj0Du9wKXWPzyGgwVfcdV2A3u3wc1pWxhi6+JBENInn+a6cNUhMOZSfMfs
NLv5LZXGqAXLs5lyECM0IFCCHYEtmBjUpFCCWJy5kPRmdLVZz9crN0T8vQ+XvFa4
pp6RYBuBCfZmLGX5jzGkQHgJNOpqYE5HF77D7oA+y+6kXZ39WU5PJWx8YiL2amVa
1hc1dhvorW7UK8X6GJ0ur1uHpyyoHvubUazq/dcYjfhmbG8AP2CkICxdW29T9Wim
X9H6A4Mgy40M60ar/gTj11BIu5eXWxAAxZvT+D34lW0bjuLzE85t/ut/uRTtsuPE
9NHopEV7q+fJVx4UX92NqYZNcZ82wAdlT/n4L9/l8+x4cs4yrAcbh+a/IVAfJ7Ob
kkfwQmAD1j7q6RlzpohJJOZafxkDKr/gs6skOpOrNhuoB60L53hQnDMB5dcHgXcS
nEX4djEokFcvUbPqbqOInwMVuktxbSzpUz62EcaPAnX9TK41fTE1T/uiqJW5aVsj
4B9gahBtagAZXNVYCR+CzHP+ZP/1DxjZ9bqQzj453R0p49WVklY3Hxc392+Qcb9R
eYEsOmvUCUNOUqPpQ3PfNdKGYrrt/+TZulIaNYoIN9uv3+XctxVO4r1T0xnfEaPd
mSneBru3oGhBwxVOXWyjA7RCC1nMX5GmYWiWLadfVGmze4dqRiv/bKCgtoo8+OFE
UDTkdvbvreXBaGNnkfe1to6gZej+OLo3ivD6kRPvCUjNHFZXzxGJ0KzUciaDz3fs
VhS1q3vZKaWSqD/nAfiVvcogLHaVvmbgqmwLAbfWbW3VDhN03DXRk/+tN+i8IEnL
n1kgNi6X2LlbPhYIB7ncxacNxXabp+fUekh/sGUTeiwsArhcW4bb0c72pN3k6W1v
QWvRUL0L5Ijo4SYgzk5do4Oc2IXzM60ngN/fb5jSGkcKXWMcmQnOEVz3g7+mNZ+1
MVEJ+C6eY1/DS6jPE3B2Zs1UpN/GG3UwDfft85hRM66TCVQget7k80QYrGdQ8aAl
JvGlThD/NeMNjUImrNuytQ+FheX8eXN9KxqitKTwRsUAiATQyVm9FfNMKBhFQx1C
2778y7QeYqcs6p6efceLnfa5RjnQEY0xMjWN1AXK/h21BvEKS+wj3g7qh0ylVH1g
6atDnrVk4XF0PAXHwmfVKJbnuGEGNArIqHVp/M8GReQw1CzebVcuJFiZKBVxF1u2
Kn8K+BoedVCmH8LR7OpI2bxFLlDp0HTehlFrNuPchWlo95L13xynRgpOdnqU/y0Y
c0day1TMbabKUf6qs8CEGCSxAXOk9IBvqKz6MPPs3KAa99fCSKVPZ9ZmEdbUYjDx
a4oiyo1fwnHm5BZgDqYm2QssVW3/Ao6HIccEhHmXbZPHJGO4JiktHm5q0Gc5hscI
uPT/n8GeB4oqnOD92l0NUDeLThNQ9pnyDH2AWR/qWD4bSEj7DrZfmxoxie3y1PoR
YdRg60BV5LX0+zGMBjuU7+jsWwafc3F/RHuKN9UstsXkB1VjXfSL8VYROwl/jYY0
+MHgiHy7ZWhaCehrWF6XXvE6rMT+WOxC+qsjh+zgSLdg+e98e6gh1CmA7gYOPNOx
KyHhraRJvcXa6mzz955GmAe8plsKLMjN+57SEdpfp4+k3nvzVObHD9vtgAl3JPxe
V5z6eF5otXqbPzqLeT+iTSfi0T3nm2bGD9zCsPTsiybEEONAmF/DkQrIvGOhaxCn
XtCSUzByEXqkNMNLVynaL6yX7oWRu2LYUMMiz3mH5W3vQFt+1Ohu9mZz9uTxIjhM
guqrQei1BTIeLT/yMSKP4fxHeQ4uOo1d90hcSipzUxsZqtMoGd6DKE6GiPThBHPn
p61z68raUE5/+pWpUix9Eop4/lleJSgf+lvYyJtaCSKVIeFzqidBnETpeBLKi374
DDZrEeI37ZBg7+G2AD2JP6weVsMJmXuoQsSN1OrHnnbqdrnqRABC0cwcvrF9m7pw
ZQ5Aa/Oxnl47ilTidSVh3hp4e55QlEMwvtzU75nj/6DbAD1XCj8BJx4ASThl2Zgo
ygvYxR8nN/2KyVGrAANUK0yZdLifvUbssdnDEai70BjbXvMhR7JsbT9LgISQbMZD
1mYnLIJXI0woGgHovGsEh7WuMrfPmjjC2rUc4h5JbIny0llGQE3q++o179vhOquE
NIjpDZidKj3tJix+vmaLOBohJtvOuiHlHq4aHn5u4g2NLb90ysPIX7wjRBs75cdW
F1+R8r3wN4fEcWgOSKWLl0q4qiJ1QCm0m1DyDVCTVYbgX0PpTj360IFuzGPstqOb
rztk2hq+ud9be34tqLL/Tz9k0oEwylNYBLVy5UugFvozUTY8pBC8HixJ919EbyDQ
iC369zj/0RO0CMGCHE3T7A9minJ0vb5QU3sFVLWna6pjfBmGHb1aP/w/RWMVBytp
dhrF70eRu6/vva670p4p7Zb2la/VgUcWtAKG/Z2fOag7SjiD572DMgf0V0/MBASp
TSiF5QjmskkS5HPCy5m+9beQI6Tk2wjN/JDHdiuCGRZ01id5XHDWrvpC9+QeHMls
wpl12l23jaXVsSMtpFHBOY7FdGeS+6EPokjHBQG8+zADPALhA/vaPaWze2MplOR1
jp7p6NksIJBt8zCtq0dutnqacJFSDvOTgv5mbjLPiinMi6dR+4g7S3cU+L5PxPRU
getdDbPVX3avxNIsPcwKttakAqWZySO6N/V6akRtEBahkP2DBcOqIxiAkxsnJpZ/
UVuszxZigrqUfeBc2bkMYcgCaRB37c3XwCKhYISGqeeAdf6vLTnIZv9xNzQThTIy
RbeKqE/tfY3PxQ03znATN5h2Sug0azlGGkSk2DA9SyKoiUeAOJQUCiIHByr1PwUc
IvhFZsfS2WYCu78c7gejwXFPUb9ImPlNZR26nSdgd35Q0W/iaeLhmin4qA/dXSbB
/+VU1wN1UBhbt4/U0udRVDk9mauvjRn1JWdMX1QTImU+IRwnqpjRrHlFSGHyb3Db
LKMB7P/Sz35Y561zm3cvUg0bVcIpXLp7JasaEf2D7zSsW0RgBn+HwGLdhf/CfFAQ
0WMYa32jLbg4Q7yoToZyamiIJqo3r4XHMYndYw1MstNTgvRJJ5CUl7zMOHDh1EO/
f5stjb5db5aXG4a8HhSQ7sDTK+Iz4y1vpBNMJlcaK8Ji7Z3g19y1wSDjznVztQXP
diw+RSDlJzlR8qV1OFAupwB7jFZfaCqqrNNxggjkVFjkzqtNnBDGCg0zhzuPkz48
ra4chCQSnea0PAxrFIrV8NFtIJPkKdmetFSSbJCWCGdI8KEPpIqVPvTfMhJV6uqL
sgqrhsstg8AruuklCRcA4SZwLwjO16KwjrSJilXdip+eH7iIQA/iGTo+LlFY6aby
opyGH2ynaFjHFHqNwB/veD7jS/oBgU1fvyAfFSJargF2tBNNFY9GnLm7Wp0aLaEE
TmgdFx2ATawKlECc1xKlmMDwpT5BBya5Ecf800qNce2jZkzR1VSSYHM1nPc7hRnw
fTquLbPoxDKccwm/R9UiJw+wvbWuRZTfV2Iq0XqQrifGTAAJz+DMC76xWsJuylaG
A+iss0v+x3IfB6VdV81XurLaEhhT6up5aGDtBwXA0eSmJQxXN1zRGOQP4gnP4fp4
2egzmVmvEWB5iILc5LcJD/e/tNCNXCbc8vFNvxhwRo4TkEPo2DAJ+RbCfKq3Sa/Z
RrfRld4p63NftoBkEsz65/z+DuCTAuEplT9D29TRMqYnB2c6s+JQQqC4htUIo65w
LlPAMDES5jSDetMb68ja4jo3Tl0Rj1txkaK08v8zFVQYdhakk7lDXRVroOticimP
9QlqjOJL0wY6vEbyzwtfekShZQlRrQPT3hk7ax4VLeYSA1aKFaoMbbY+nwQxY2R0
4PTQHxfd0A6r/I/YiRwmbIGmGHaBVV12g/p1WlO7y+NPOey452WKSDl3MPw4U8Er
cegdKpZiQdsz3OUr+jlbwoOGY5zv7mcRZ6ZQcQkXGfqpaqzz6+bCK1CeOHkLJaaY
Blx0AuJPY2ea/lauv/2KZ+xJJ6NzAkPAlh9u2lz7uowuy2Cj33fDEnehRH0nJmq7
qnMlp5DDC9KQEvxSDc9MhtOo8lCa1q1VtN4EjfBP2GiYE3f1CnNc8bpFuhmP6Cl3
xDWhBlW7HBIvyHZvyd5WjXzkpjNy/NUGiwWIaRlTAg83AUgzw4WOa1yEFt5VHjZR
hG6mxKSRZPUn/JQZks/WB9IBP4OGpf6FnYnrP7k3tJuSKWwXiPCccAOsLy1JIESi
E3mIqyub3foMjhdAGOXYrr9l/AE/9GyF2LVx09WtP57BceA0rkBw6w0SeyO0fuJN
Uy+vUrCIJzxGKoS2Di97TxihI08ACT+Mon9MazoQuhxy5i4oZU9IKEsV/vo1Ugwa
Qfzp2JGjimKuDEuuuE54XvSacPqIpV6eUGM832y3MSprcqCm9l/gEgOQ5rouackz
k6YgGCOaJC+3JASGQ7M+OU5HovGIHL+3gcgUILPrWGD25tzKwDVnvokApxmIcSJn
QzEDwWCfeZzuNRd19D5vVdUnM9TjtnzE+4LkuH31tB+6B9GrgO/8y//C7hex4Spp
YGeE5ByxxA7efWH0kTY7uVkWkhA6nEZsoTBG3JAVzDiaZkDkec0GqM76aFbSqJ5Y
cSASOoH1oNIR6HPUaXn3bMQj1kiB4GfWnHainu/CfhyhgWZdGzShKRFFlmK2MFFY
DxW4YX44WLps7+cYGGJTU8yOIcs1xynLteBeTds/kcxh8gY8/KyqIhQnszsVKDff
3kgia6OLyL99SuAqxbkDVNkgIP0jkDF3GwbqT35jJ1Bv9uFaaFEI24iHd9pKMRmx
99ROvKz1sJqn8UkA4X0JASB1X7wrJuHD2xOOiFNEUX2iKe1mmSKbjaLD7Nqgh0Yt
iUSL8NbUUTMo7nEQ/vSb/zoN20vfylhr/eD3Txu3Pb3Qls1w9Zdf5WP2vL2mSu4M
8wYkyS4hlVlRghCWuQ8knvMntVhtavdnNxHoizcg/f6T0gNVgpi9TRm2RRFagRQM
oWzHt0Orv88MVmgf9CvcBK8vNzFfJzcjIJNJfMJoLlqbEmWLfIfBb+0F5l3L757+
XLWEkLBeD+TNmDsemIsNiZd10tjL8qLuu7V4PzSZ30RFjIhcEEct+KOgOV8pVe2e
lKvXekGu0NMnnbBu5YQjUk1mm5YPfCtfBRVOV4W2P5lK6mDRGntpRPb4iGGClkh/
oJawrq+d6qXJlCDPEmQt/rU3XdYhRGD89855aAI9IJav5RAlQpmnge9l+kyf1LL9
nEc+uJRYHqDGhIDYTzpbD/37SrwjDZgProJtpu9AAWYX7d2gdEhqlpJ1LR0plMSD
tJbqXgKIlVcPL+giNEczCkzIsWw23i9xpm2bMwK1AUcFnQir2S022KvbGWnRpkVo
TBzRqPlcDwPyPDyAqSuecnWAwnWqoRnXIy2xfh9A/FFt6QZPGf5pa3mB69mW/ALG
ogx7vWuXBUs/8L6PrXkr7reZmBOu6z4S2ylOIEEy/cKuoKRCGDCcGbTKxZEJHZ5e
loKK5pc1bmFR01dWyiku3+H9wfmLyDh2FVJoLVQz84gdCVUd0jeZtdlroYITL884
eGHWBnbz9CoqpHgfPmnDtKqY6zjaHLhEtPCEBJFvMJHofSgxokuun3aeOIlrsJTP
Ho+T07VP5ZGLbeM+8X++abMJW5cTAsm/krh6BySRX1of4hksTyZNnFon+ZInDrhL
w54Ttbz9iu6U6xhSVIrjlWjMKl2wB2MhBH97svjPMYxhJV/Lg1WxNbHt6kIwRRXY
tJBO4e/oR3aRHarnv8YOg7r5gZWLZodauK3iJzOtTXH7UNnAhoDGzcqXROaMMG65
0Act/5T/3kHIgrf2SDMdxqqJCaKC8APeELw14XQWhvTxbjV2pxoQ9rluB4/JZ0aU
Eqr7B2Rfy/sMD0aB02NvhpVDYkizbVSWP/tEJk0NQndexmW0JMDSGOrofhlsobZE
U6j9+zKTaDfDnLORbNHKFR7C1+Z/e8X36Ze05gZvGeF2aWSsEevs9NowT7gWjVhG
Q/ATlMvTSNNgLeD5NoWF2z4aBh5CRLUss3X8/tCjv4dTJSYfY4UDih8g2taxcwAb
atyEgVLJX2nnvRHABbqWdu8rRanBj3Jw8UmwfavU7r76oXE6FXG/xRX6KyHyL6uN
XPiIldX79duIwqrnSq+gJGhPGMg+fJ6VrxL4DjNdSCi0q8ngoyQ/+lScLFRhwJVK
rG3GZycUmo4BzB7K/dh9WCawEKVwf40NTe4lv34QINKlzxgYx7NVlNUmSCPHDoC3
81HgwyJvKNvoaf3E+DuDJJkKotBOzOXz9X+6SoVukb8XrbvviffhX9rdd99Wfjuv
3QMbPL1KkIQ21Iv+P1dyIT4B7XaF3c+CopXtr6oLhTaV+JIwTipXejtJpDT3XuRT
UO2VIfD0ckH8OgHZ8EPNKTBuMdwqRCQEJoSW9YY9YJ8KTpanDX21qzCOIUXwpkfo
iHuzhwoifgUfLPJV2bAPBcRTIhbbQd2GLF+Rxr36SPsPB9PhT57YypzHhzt4xqTH
AglluuPCYAb58kkYOaJsTGahauJ2xpnSJsZrz5Hqxm1COj69tj8kL/+MfRwyH57J
f4j5kNrcorpyskO6ADLlivq/2G55cSy9wRwWymdJepG55oZJ5BY/kqY51YZ0vOgh
lDI952zGAhnhWCyb/2CpRqTeyLuJqDUmwrqqTnaAlwRU/xAGTjc5rLJAffSzadr0
mOHrr88OMYPp6M+cF+Rt2TuAbzlj7KS0gUEhJuTK2MFb8MIwLdXtuBQiu7NxsMxY
tc64kxLXObwar8y9eq3tXOsgb7vwnkjh36Izn8snOlB3I4bx6wfO1nJvbx/mgxXo
8EFxwz3y8S/AlR66uLAZGf492h4am7t41etxpUK+hRG3KpK3IYKX3fGPFntkdHjl
wFTyfwMIsC8cjcC085SuzZ/InBb0XSEK7Suuawrf4/PbSjeIz5RPo68YNQJmunp9
iTucVekZpC0eR/G5PzaJS3B6V49xPfA/aIUdVAZqj8l98y2rdAJZiQ0ftNzJtqhh
NoPVzJKPxYQgQeMX7eH09N0g2A1L/rHwt46GWT+P4REbMDLz0Z8XmE6z5HE6KSP8
8VIZezPtp9J7Y9t63QysHuTj5D1+ELVKsxUk5uRYxcMJ2bmsVagiOfpxzqjUXbr6
niWfS8LXeooneFms2V1TbR+5u1P05kQhrM+vaLHkMHY42mMtPxGcCybTxyzpnKhz
jkr2R0MUrIEPA2Anw8mlVppNR68cZ3E0RvRkOJ2XfFiyycj60G0kwqQg2JYqimQS
H9MlwmKdCscHct7Q0rIgGBdTzYr8KJkKk+bD8/2bOZxFxPbsAlsK/F5SY+mLJWtV
Vx5xlGXdJpjyXcG1jTdw6ny9TtYAcVEX5Tm1EC6dRYPzq2aV2tIeXKLZBylqAVaW
KQyTqWci+jA9eRNlnyLK3MGYIJ3ag5rQcRt6B2W8x00bguypZPGVSEJHEylohrdK
o45dE0DJgWYT2LmgmB+oMviFsuGqsbUavkyzpX6WaaZ5088ZMJctdcf1FpAc4ZxG
NN+oNo+l2A5uiQWEcZamIJJwzjf6XbQyY3Hjy0YFXaU3CWKkL3AVAGQsvnAe+j7G
ab/SpCWowQKRV3fhy1Dyt5KGKRCMBCXjontLLR0hY+IIouIh09L+h76cSD6zNigP
z8rRgbhnZJ4U/T/xQIAyH3OA3KBy2jLQtm5vwlqSSgtq1VPJBvcZnmJHsoxiLkti
lD22u3m9339OKB034/W4a2RmK4RCvLlJPJj6ga61wbwZJae9/iGn+B8iRsTVbNqX
jJNKFaVcU9UaPDl67uzfOfHNBtKYdgbtHtfmVBsHvo5xWZNx13mgcKV7xI+St66p
tJDVH2NXoXwMUamX6cAZZLelMrBCczyNZdoBj3kQ2YhfkhxsvKUPSxtUeaHKpGr2
vdLhi5+N3EgSxvb/QLa9fwxKigOOZreGuPBY0drXT/ljdZhiTaXyMhyIwM229LhN
69YCb8WjMgUNdIWFAJcT0uujeCG/U5PLKeHr9EnG2sYnp9o++quTuaaK1P2fVc2V
+BHZEu5aAcnXS3yqzS+GOhnUiJFRmFZ9L4sA9S0GcUb5SHRTv2bImzvx6GfDMP7n
XJV4yim9QE2InqPUNg9wZZyFpBiqLjJGUb7cul6Rs/zwRljrtGuvzGS1AUnxOXQR
r6MDyPK/QGVLmC5/9R0iQkbmTINu+OK2Vqngbcn5wjsmjSRxcpnDUrwx489L/15A
Ec7vb9S+sVz26UcA+5j9st1KttDEcGY8dxN2az/aAVMI9dJhWER02pn2lXSNVfhW
BqMyMw97CDO6FMQ2k8ADEbGa6NLN/YYcngyOGY4MrjhpkK6xLN/lKNISSSSWI9RH
AaJ3OOG7FoRnCrg447UhKhWSLdXeT0bDk1XNmZpiXDGkIw/RBAa2tFUPWyddwGqi
iujOzqxtZHSWcxl3GDYpZT5fkTY7koF5vds/A/vmfRuefGpwBShxVrDnWUVmaHZW
FjeRFruC5dSdHCcTXCPPWKd0Qvh/wf09ZU+Y2jaLLPaC0K90MRRA/i5OOoj4Uu9Z
FbxibfTf+qlqCVIdVetFZbMnzcEWCxXSWMsqFXHscBqB7Ume/OYDwNhGlIteIk4y
GqmtA+gbyRrWD6q68I2UqfBrGJfov3s//gMwkSQKPa0ByoGT52jdA9ffFhe72Fb1
oI4MoXeyVxO8R7q24cyZVoUHpHFlpF02QdvIoAmnUTk57w6wyoGXAbrEdun66vul
yVL5b55t8TY0xB41lz7mnonPTi2lhWFzx3PO/g8RNKC/ANr9fKN/7b0WZLiRPKGF
H6oQmql12Sl0j1RMeRdRBoETs2kQQlpPw5/sKtWmfTbuGgSXBJ9dvSgq8E6l/W8F
DXHtpGx8XZ+mIE92/qrYGMTdV0DZm+9GLBXa3XykQAoa6OqePYw6eaTB5REHBCLG
Sf7ysuPVVaeGtpBTPRMBoWx77oU1Ry3y5fT2rV3Qm+Hb1TaeOS4qsANNp3R/f34G
VepRYXEZ6uAjXHyU1JZgnWR1OM4uY327csqUtI0kJ9sxtsoqcR9bRXjRJ8JontSI
73JCyjZRZd+8sQPjThMr4CLzGeujTs/S+tJLBtypaOvHku8Bk2BXp8B1ygjWIQR/
28c5Ba/YSuMKMcubTailMrFLCNs8/AoWI8km+v52950L85FP5xbiW6rK2KL11NTu
35fnLH38epqsfdAGHZcfzyuwXMpa5yQ+p+lMpC5YyZAv5ueeKZTxPBiDmYbOGNfv
+y8LjnfgRy2/zZqzyCYzAF+Ju9deh58+CoN1G/uMbSYtzOb9RHMUfWJbsCJ7jsUY
em2y2wh18wfgYsLrTpNW8FiGlN4RLVXSjlfiNjz2AqnlZSafuViQVA5dkQxhTF6y
mFK7U6RgZyf2ylDsh6s/MqHPnjb6TyT6JiAhrJO1Vj+2U772UnC6SA+Lcl7mV+Lu
Sd1xHb4lw/9mi4O39yI3+47UHwJVDC2qvcZMZWUNmREFdsH9EUXHXsCfzSOfaY1Z
ZEfghgF2YbwgqCSS2HRb5YeZRECUlpFTiDCIVOhyMqrKZAJpCAf3xakVwfynUc8G
2qurlb0UMRFoyQ+q2JQ1nWJ4lqZWz38YxGJ8seaST3uD+XCOF34K6BA8SptcVTGk
MZWTAL64h7uGFdQhOxXWcSfNXIOxhC74HVI691TqODUemqGpMPBaK4OqU8VpKiJk
kElqMYJxUujEl+2yxb2nlfW05OP/UMNaCkZM1YGE2hGjwJLdA3gQ29h+5labN3Sb
U1Vy4J3ca7J5RvOlGG+No2wuf3icGvMmiePauVtny64b5QkeloG2tj6HDMV5vqNm
xVT1OWgT9nmnmWwqQ2WDhH4sYKQLFXyJXUufzxpJMjM85IRnj11E3FhPTvSGZuSC
Er1Re1sOBbLVtDwy79dQOMjO3pK+65WCu1WLeeeluT8vrUArpB+3hgzYnA+7/Ik6
XPpNVtLci53hcFRVPjJymyasGWtzofsawouJb02f3M7UcXPSfb13qzB4Cdz13LaE
HEreL3MdT/5ciJDTVjmbaMkyIRlpYDI6q8D34QAGPoZQvEV0KcGQ14C5pGNRrQzp
`pragma protect end_protected
