// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:30 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WxzsH+NZ/qxTCPb2DylH+LQPkQRgQzZGFdKSe3aRH+Wp1OZ373VySwy9aujL6jEt
vWW+12bnh28INRC2CAJ9smZxplvOzGWG5WTrgziUkR4A0J1AYb7VADkgXmcPoz7l
dLWVuNybMWRx+bsakEDtu+x0TJXJ64rkyUJ3aFJvco0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 63408)
vNk2+L3RnJ54zJCWy2LxYV/lMEoGI9yZ3FpE7JHjV+8X5ijetpzPBmN0eEQN6ETG
FYKErZBWuabOqXd1UfJRySYk9lGOUZMBxq59QtAiRsfMpPMYO5K1Xs+0hpKhkcOE
n+5N+o/aXD4K5BaEC5RfOrC/mTOJ/LmvKz1hYUTnyQxIq9QUc0ZaZHoSo4PEOnK+
C7WSkthY77PoNi0AAksPvnHmqW/z07lt7yE5fGQA5xhktppW2QI2ytrNaX3NN+El
NuRSUCUoBt2K/RhB3MxJynUuEPKAkLpi4Ee8bIKMEzZqhNgzC7AmFuNyQ6InC7ha
uFtgWZkjrnXrWyqdMso41+z+32b7H95NvxxbuyyWGbHfoSzAt+AUCShiF2qE3sbJ
BLo3GPc95ReBX7mSDOyqFIDL8HZMr9STgOtQkIUJvIxc6E2nUr+deBnTYjRFsZCj
v1hWV5infDVrK3XqQ82xwRWYIA47tL2bcOade9qKavKt0rviC8ovM50U0F/TOCPW
4e8OGsFv+BEkilBgykrutofUVns/xMGUaZOx6zYbvsok4EhFFeRES0N+XQ5/eXTV
YRqHR/TELuFWxt50xBcxvyIKj8GSBTlfek4rRbPWUjWAEXOXzD6T+hqm0OuOvJyi
3O/aeygcDoItI2rQwq+R+cDaWZ7TqKPMech1t8qxYZGR8vNG1yPgHn+nrI7eg2TL
kLZmjCw5YQTaMkIxrdguijTm/SrEA85fpnqaYbkbzSHjU+9EdP0kL8k5zS5z11Lx
tc6X6i4xaUfC9L/KdNspp2SNzOsd+va/jpSdC66dP23BzSdbggc+6c0NFS8QBFNI
70dw1VTB33iB/R+CFFYS2t6VZ6taWWrNLtkxsFN/3oqKtOf3qVO/xRqlsU1E7yzL
mkzLcQa7Z+zhazHuJqbB4UqwDzSGSRpeM1duPVhR8zi9bwD2n8qiWNJ2k5XzV5vS
UoAAd/R5975y27JjtdUM1fED/WAXfJXOKOflRftj0pOQCRmkKk24mKFnXR+QtF9z
M4FsiAsbeh4BT8EmdbAl646LweUA6/qRHgXfS8miFLEEkDyAXXZ3tkz49X5SpkxK
p2eBE454WyttfjtZFwpenKkG+s9IXeRjxwGuSmB0fQjHQED3hlGRLLqPoXNNvRP+
2mOQi90NaVm7ZEwtd2Kl2as7nYoujw6LNq3FOXp5EvAM+nrz+0VnvHPlujxxnHZl
xVdt2Hj74176bR6THwrx/T4GSx06TJPunXhdO6utgg0TcwvTZzclMinDJt0RgUNt
63TMWRmGAQ+4LYPxYLZuj+9OOXCSDaT6uu3+jb5yCzt9itpBz4aqFmRhlplfpdi/
WW4d0KrfxzfCxiLSFaR854pOafzyLdKpsMFU4VBeva0VDV1UPoQeQJ9aFVSJ0RF5
Ep9SNqtHeSOe5HvcPsp3Nj18uby6zdpb2UKhlxt9oXV1coo8m7rbmIW+7eHYLsgD
Zq946vs8k4hRDObbi21PgI7qC/MqOfEHl4glfWPe1HWVIALgrd6sjtK5eQLFL1EN
3awk4k8clw92XEO4rcb9ncHOMklv8aDqpNgnybJJJc6p2A+CMOw8u2oUvEJPPsBu
dSN0eYSEvlSI7+t2HNIASTxDf8hsQsQ/srNQXrGDPal9Lg25dwuB2qJM5KJ11Yq2
ygqEKfNvqQyzHA1tJbknO7Xy85Nk4NU1EvLyeST+dFrav5Kz59AthVNHcaUFxp7+
YMJMNZDssAJuseCJ9JIPBx6w8bixelPWMVQc7K+PGvScgLOf2b1xWq+zprHUwNw4
I7J9YIt6g1xOkVKBd3wykR59R41mWWs0qLYV03l014EtqXrAR6TP23+2yFaELIA+
8OaA1XhJwK/PGlUDLb1rz2P1OSceteNZR5nvNI3NenWRLxczx5RlpinWi7aCGExH
vrMcdHANs2SHMqIxi+Qoqtk3qSS0i6gsXq7tgspzD5024iT2OuatmYLy+sJ8mH/q
mBXdLUk1LlnOPMo0h3j1d1JoqTeBdEZJHMIHwWH0YAJ6jvj7z5ZFBQBOX3jGX4hQ
Urmu1UEyb/NVuJurE/2Mz27an51tAoCHYwsHgMEQKZZ4pYk2PrHdMWbM6s/UtAVv
BiItjIpS8tgBUA94Q6hMEtv+bAaKs7PhS+EJOoUww4d76HFFq43xB0ZymgCd4kZW
5jsHQM1nKST5bfAjqkFZh2/UyvSPz4cUWdj8atlGkFllD/uwbZwPibiX5RtN/QR6
newGTKXRkLeYKZbt3WgQdkfG3PPaHoLr4l4BCtMaL8IsFc7VxkTc7rx9BxXjmM9q
kfe4VK5T9eFmRKZV0D6o9t7p+eO1PGTews4F84LV+BeHUq6weFiFSuMLZyHpC2oL
f+C+edhaM5rAhcTq32X2dB5wXEpGHyFoi3MxK0AMJzIfr0vkyxmszwu6EAtVcFLc
0pkJ193MN57gGo0/oMeV+HN3EVg9cuqzUlBwL4Ohlka+DR7j1vBnORNYRuJMg/fw
w73RiP0CgYvMp1bUHguw50sfTeReZh9lGhNqAbkM//qFBLO0cqy+qVs6I1zS3DNW
4lS3IM0S5JiE0CIk/JV5nzmYHFw9h1nqnF+AfPoSrSn0ElO5zD+U+Pj9o0Q41C9N
7bitAD6yq3093l5DRNoM6bAdeFxaFyKb2AerGmhPxFuIMx18KA2FYhdDyrpjguIh
N0xRUq9UPLdbEvD3a3VvEHHbvtxUXUz6ujCZxiJeKZGnEqmJbJqCKSgfBJ0hTuPb
xvBTlMCOeHDeGFDdOnorCI0eCkit80U85qgETn0q9Sczqht0iDBQFm5x8j8y3M5F
3TEXBVdBAoEkyVcdS44Vhnp1jjBG1pgY140hyXnoTHGF2ryOeIFnhrGyt5KpguzZ
sCgzYHVgddyRf9LI/9t+Oi9BpN6IyXkSIiAu9V07YPLgcOJGrJXQG9balY1CMVgT
QsqGV/KihTitxfy5nLHtY8eWEPi7qADvTTGM2Y+ILaQSCp5gUxf/3LlIpWavwa9L
qpBk9WcoG8dYkMz86SZUw5gQs3N2tDQLmhBFtn6Rn4ZVKb07w0s4saWa3R2eGmo4
4HDG54b58UVEf7cpm5afLzhFg8V83RLAibiazhc2Na/d1+/E3AYbS3guO7eFr6Oe
BLDioZR97J/VXyCi1pKUfKb6OP4QVFN3IU+CkzesU68jmea4BeIYOIEt2W40N9pM
vPTv0BQK3VlSjyzURVItDY35WQrhPUrCjRYkcjJMLV9TETcLFjRugYl9uZEARRPF
Xbe6UXoKwx/vT0izIWoDiNjbaPhaYHFCqe3ZwdROSWKxcWqqTPi2luleoQtZOsAO
JL2DL9zDfH22P30T5EqjR+LzvhcP4WMP2YPZKV5bsQoBEZWpueispLMvcrgFwhGE
Uvh/V8w9uib7Si2pXhnXtsY5f1khCZBWjRbCyQ/ER9zbVHxvzfZ+BDDrkraBiNZn
1j3vGaHevHbi2UgHlKNxvVFu7mY905FOr6I4J/9r9nzqITxESCqd3rCBL0zBuFBF
oxERLGW0BFhYrpd+l0XULK8TKHGbDBK9WQ3lFMBH2ko4dG0GmL2o3rU8dgFANMAm
bKSyQkDy2Q8M8I5XI3iFUGMDg6BKDGjlm/vXhXMW6lpAig2ObH5atH9BtVnP09AJ
mb+TlL9BPOqT1DAaMf1XmoxtR/e09Crw+AcuscQMUJURjV8a+8ahMVe6DtpPZm7U
ZzhF9VenSuntM0yuN1JEkmUWcYbw9sQOVMTAGL/YISlJAeUQYFXc3fSlSmx4El5D
MUyL188UBGvtlRpDuezgB8Sa1UIrqxt3pGDkHILgCpf8yJsya8dmwNuFMXIlL49A
qU9Mt8AibeHjowIrt2JxA7bo7UTvHk4nNP5m01uWv8qcGZYzFJcsEqRIYk7zPDr2
7n9OT7xunbTA8zFXCKjmRiSPUjrc14agl9GYF5+9Br+lxVQus0PizJMoy1zA9oQm
yldr5Bkx/o/4XvRaJCSFhw85EYQaQ+vVlBGKaawQ0tLgLvhnyMiCdS1LFljLs7vs
AlTbXIq1nmTW9I9RNR/TtSepFb4VyRIQqY5Lm0E6aWXYtff9P2mCsYaV62SyphKa
qqsgqtSHWMjNuihgxWBxBAXqP3je7ZZEuO/CYV11NgG3ZMIuP6QTeP+zwmN+Yw+3
QLXolsNU4aQDKE382Af+DCW4CNCv72oVoZ1IAVY2FcJOdOGYYd4biwiD3NZK+Jm/
4buPWW+2W1NAbUwrCoCeEK76KScmw/4Udr0GiKlwOl7BJYMoFe8E5qocI/iQvSvp
QXgAfZo+HuErkbNhzvv6XS7WX0q4ecb7GUr4QAOwmqQdn3yatJBMEAINvRQYp4DL
JG+axFc71dsLq4SkIroDF1sdxGU70PAT0SmePthNrolaZwsh7tgjr2ZoRQAp4Rdc
68SXMJtmhYkNZLfTEwtxqRE33QKWOK2YHrhJjx6IfqQJkYSG0prH9mGWkJRKesHK
3ss2dRDofOcpTpspEjw9i+MQd5KW3khv+d/lzJnAlqi6RL2SG1PiuDckcNErPIY5
JwGcqL+5Calp/SNfOY4MCsGhl8RZBElZhcxBXSNvL+QhVBxRMvDuFnXDNi96XJRn
uakJHiZbZaOkgppkfHuJ9dX11e5ptzo+gpnYmskV75aNoO8BquDn/Pa/Q2RbDDZM
Ybpx+zdu8E1Qcfoi03Pv5By4iwAJyrUvKfeTO8SArCImSDGucdld6G4expQRL5U5
ji08A4kJSFsO2t0W4EqDgth14Cpew0PvV+NZjeXhEVmQcsquOwdTJ8ka5Obmy6k4
uZzUOAIVts8cfEOc6pj1iU936YfX/p0j4FissO33ZCjgKGluOTd1UtscVMFWrPjh
z3+0GIs0lCSbxQMAa1IW4HQxlAdkwt9mOjlyjjNVUhRWNXLwSetSFAu+JDVc5KK/
ekaKHd9IPKrnG5CNKyi0rErQmodckkXA2HHmHIAu1w1ZoynaT7upgfEUj1yHI+xt
egVknNkzPpSsTQLa1C4kxJk4BRcbYeAQjWHgCUQKF73V7iXCy19tcOQGFipb1/eW
DoRCM9vvv9XvKn+Puex4yC1KUikFLe+yuIPpeBwUzfdV28ZFSDxVZkihhOhpZGT4
JijZ54CboPg6MAz3nU1imeEQgxnNrvAUsQoHMOXfM+ah9RiRfyruEaQnzcelXv27
dOJVdJPDZiJqYZjE/boKkrc5WQGdQ0NVYIlTn1C7pym2vDBmlx87qvJnSBE4/q3d
bhubQGRqDVvHCSIG25tmjPixf9dF3Cj4Hw/STckeGU7gsQQUSOKgoy3aE+NxynYu
fXaThZJt9AIOVahyclsmE3jYc2lSY9OPLaVevZBX/IJqXpZjmyhQ0NRcvqmR3BqT
SdaZQH7KF6upj0nDonS76Iu7NTZORjdAPPgJOY8nvkyPMi5jUO4wUIoyxin6S9Tu
JTaLqpqSTTDQqHCNyxcVviJTMDu0RXR2LBXxJzBh0odm5ivi5uUHJM1Aod+MQYx9
kFVMbwzNOq5bm1YGrDOotlf/lAp7h6Qrry+PFWUYlzV4B6KQgq79q8i5fp0M/k/n
gHLetJW6dvMMofI6UCJTilh84lmX+p/o2z+7wUwEurUM88YcKse6FKaTo7Nqpe27
oLl81Vl8NNDcxiaIP6Z6jNiERa2NExnJCmvaFngdp9kc3fM7eaw9EJ4qsXpJEg0Y
gFDlroD6wvGFWSF0PSMgnar6foRb1jN5uPBeQXmDfrJNuf0kZC3JCQ0QpVcDWGf3
LuOkj2lwqWEWbMnaTW+JXZsCa7iKO4ORG92SJP2NN81wi8PlMga9X/OvCPBx2vqN
zk8Jtx7RNsFhxMR13OAkxNg2GeunraiXCxbbAnnLaCfCeQdYnxhnhUiSItBdLr6e
Qrmu8KWKCgYSMEfIpCtwhVwNCj9Wko90qudNbFkXQTo1QaWk4d5m7z6vBsQTCVnv
l51ib2ds6fr2yQ0rbG92ggjICgDUAh7kFVcwkuUDccNRJTJ+uoOcSWNlPPW+U+ti
0B37gzHDdB69MQfDOuG6MoxqxqGtJXuuy+iQu9f1PNkowZsss++8ijAQokI8anNq
IVd/JCY/Yl1+V78/AwLp45Q09w6gLtXQ7D0nF9p4+A39WA+zlo2QI5Axv34acQ6n
OIsF1im4c7M1bN26D/keZB614PGaF724Xw0elY60PQ2VnWRlvVLbQK+98JIVV640
klKfXsg7OgkkTeSqpxbe8pOnZ9m0pLUp3zPHtCvpnhQani+XDbL077WqhBOXg4oY
2z1fByRJvbS0G+6DjSCuqiX/El6X2SLJfgDIPp9Guxvd4POL7EK1S4KRXldAnSIo
alV7zaqkpowgJ5gXGvyp5c/O7ZUdyfVmvfgxARDOJbSq6nAf5wA+a0FC8KRrt4fq
pIdGisekRimRsuEMAi+oQyJKtVjwXC0v0uNe8lryyuP6InJI82AgDjDEGGBnm9bD
LcXEQ5tGL39EZOdJcOHpjh1bfJXRfHu4upRaVNkE2Dy/M2Vwt05XMDPU/AM3dQLJ
vh3qXJ0b+EwMaeQrxMgVlfdiqHYW4QBunYb9hhN2Av/31GM8iI4+Rs6NVCnmHXzX
FecsJewVf53XRW27kaQFaSskz/75ikvnq+9ZmwDa0gBn1TqMeXrczED6/D42GF5d
eg0PcUoN+KdpbjLrFcU8u82I+JoT9+NbTH0vl9us/FxzIz9KGS536RKCASofIiXI
TRK27Ry/d3lAYql/3Wv1sPI3qDOI8HC8GqSYFfDwO1e93iHZ8ktCHugHMgkW9bLZ
hJC+woth7B0UaX7AeZJ1pITjJtuN7dXY9kuRcrPSzGdCM6lxJPMm028vhSy3X0kN
fWgcZOnCk3pnY6OWyXb0oJIWvoR0A0sCzgg6MPxqn7gZXWNvLB2/slln8I2BiJyY
8OXLJusbm56wMVdtHPMJXx0lFBUKT+aZHOfU8aJjJ17F4oSa0oAx1w3SKoVrB9zO
NkTYqpd9Vsj0JGDW/bKymDoRo1g6X4ldzvo3vf44Pf5juS4lNOuxi4/w5DM8enFg
wrITU/Yz5/wGFGWWxpHjxkJcKSraZKhFUWnM5hiMhF2G/LfVvM6ETUMJxH+8vb/a
XBTKmZWwKQpSL/JIq0tz6gBa+igh9OM2CXS36Vs0AOB3kRdCPcEWVrAloKOhxGFU
1P0Q1Sip7mTnSzGFIPugrefmwXN+3XsEih0UpefFlP+hHK5+bNzcHDDIul7VXWlm
W1aXFnftboh25slvFhQBizzRaIQMu2pUNf5RLFf4Wm3RvOW3ZBDoRp3uG5LesEkX
ueGRa3lGAg6YshdsfTMF6Wir9tIu7qZY8yqejUqUUgoSvDOSjcCPI4RIAgR2lb7z
qRsAAR5rcSzNdzJotivaSNa5Ei6uzCLHGqjFspEMd/PFcQy89WBbridxE7+FUY21
GZszNzODnFLMa8EeRCYzv+GUgUaQd+kzUw1phsv01/NrQxxwPD3hU8FaAx9uTwxI
yuIHGmI/WbfJSLxFvMFx6gPbTTYcSXOtx0+RIUexet5Po3z7XOsMWuYJakHHiPHm
QKpkey6b5atHKeMm8uujBvcJDtAoPddTGucqrk4K/qOtifPqC2oJkCMMV/CdmPhO
zI7gKXTTbPcBZ5C8hVF0cGha2XvymQnsT2O87tLRLbyIFT8BqKI5m/PpcyvnoGzb
EL8kbH9G7elhSF9AVWgyvHeVaapKVWxnvGDavxFRGuKwtJfOiaEnX09dYLbgAZpI
zFwVJbf8d49z72eWjXodE65bHwNbMrVjQO/YrrBP2gCmfmsy5VIB0wS1giJmeDHT
9FnydtwsvU1lu5QYqgjftyPr68IHmQwT5+YvwxenE3bgms4c4RybVKW5g6sKC4bm
ne1PhQJN0iC0Zq+1uD5qgKzXoGd589ZvRtRoVXUvO9iYke9ZwE945Y3lMt/KDWyX
x+h8fysGmYvjcGxIlTmOoD+IxdX3bkVsNkjJo3MYXj2dM4BRk0Jr8f3mBO7yNBDY
HMXemJXGf0b+ITv3nTkIFDQiq+X026Ho735tYUogKScmBV8PMx6CNVxMDYQ/Wrql
SxY93YRZqpIQmLnZ+SIpPEaBE2DrUprezeMACLZSNoLhBCXmbT2wAPtiTDnr6IPy
KbzNoF2fC/aFxgYs2CtLSbYC7Ks+pgTbAO+6sXARRZoHUXL3JFeXBYwz9F7I0OA/
4caQ4t5G/uSaFvDsTWUQ6CZjOEzaOaRcNcGpXqk22tmQ2FBFSaEYphVHvFR8Kao/
KK4+KeZ/C5L40lS8FZn8/w+oXj6+xOGGyXH0V2KBr+4E/87/YU9qg1yze+w49Uhh
sY+wc5+ArAic99RTlskWOmQIrEAsqA7xz/cHXG7bJo+SfKPEW0UNsNo9657skZSz
/sqf1SRc1K8q6MaV2/xYQrMa0IsXIRpruY13dnvHHbFyjhFTjUxF3dlqELwn4NQW
gRQZxHEsXWtHRZy4PjQtwAzBjQlYuARdBboSR2H/xexC9QTwa1G5cUMOtbw68PlH
+RwBF0ZFGY+l2+87RBe/I6s+PCt0YttRCkereedrlsMmCydzAwYclk5LfajrLK4L
5OJ8tId3qW9VQRvhchNhCBy1WzpInwb+LNgZNfqSDYG0mfNZnZY7WPUax4kLxwmN
IOVx7KmuRxS9Jza8C5Me37ITU5grzFNhdjLGYo7O987J9b5zW8hpjJzLtDQ5qDkE
Df4RHKgAUJnLZU09yWMnAXmlgSwsmkpbWO40s0yXrVlQZ397BabSeHUbzOoZ0eEy
sPw4EL1g3TQXzqdtPYat8a7kpToFQ2KFM0ENTNgpVYhZMfEC/bsUzRqgHgcbnz9Y
TVlVGXsFbqMz+UgfX/ya6bLxT/r72XER1pbgPFHzNmVfOSQztdZ8G8hST0YN13T0
aEO1sn0KAsYpwpE2Imz8tk+yuqBWN/BgmlUucrefjV2ac+v4DCJQ09n6+48l9Pgb
dD24xwjdwJpjoq/d6Rczq9/vkV315zN9dYOSZgKmdNs88SNJlChD9d/3rlEVjoir
pyfGqK+T2e3q6eyXovU3+/OOGko+tMvCu3OJRG0NotN1H1pyeUjSoeiSSJPeOWdh
Qhwfm5JXPBXwfKCcYG4nqhG0s+5ex+z6eHYq/2GZGbjzx2tHdlEXuaaGGw1aNl5o
c4fXTAUFN/bdLgFkrG4lkwi+IdqxKl41wCxP4Bic72a9ux600T3n5UNQwOSqUfuO
qw4/EPmX/9t8aqpEN4GAWldaw0blM4ZObzPeJQ6xIHKda/XJgmGA8p1vKfIQYNEl
YQIym5VXS/Y7DLUnHcbOU4ogJ19kg60iI0vesann9KcA3tDc3qVcvHAH+EFLH7/K
Lt2E4QKUpHdsPNyh2pPZ3Bg1sZg5zmLo2RylYDnyy+VGc4duwTWNl06OIAp3x0zd
uTupz0zgd3pksHcJf2QWOXIoPhIRpzzpqTdc1rDecL8FO5+SmSIPlZL+M45HI5u9
9134Wu6GRcCCD9Sl2ehlM8GmksWXMsIeIuwYdEmRY0bhG+NAQn9Cx2Wi7qsDdRTk
gcPSXg6N39poupnSEVNEeuYn/1MicPueOuILUmk8ANAB22J08NvV9z/jyu4aYbgU
GsssniWPh5QJysSUsgsw1aKgtlaXK1nysqwI+eDrMXazJoY71bm4x7LyDxoYLMrN
8yuYmd7SmkrZtEewl6pvycWagsUiR6ihC2uf9oc+m6t+2DQr6CTkcx5Bb8qxs2Ce
cFWSE75KH3vLzRkStNJoUZJh5+hYM4wFY5sKyLdPCoKhLSFnB8PzVJyK2lkwTXtE
szsM9fw6wjS9nBrgW7ruSn6GqavDYuwaEoz14YTatrWp4Dpbq0sQi9vxCqkO4FZp
e2w7FjoclBRv/gfOxHOtaXjvUG6D8YFS9l61wG32hEjYfu97T9O7udhQw76BTjRU
IZrZ+E7t5C60tMPZDnfj5y+PnykgeW4VT2B1I6cpfFO42jQycKnKPwArUcVzs2ox
FB4uUON4K0xtDB5gyrk3nmcPNpUqmc9SKW171LfcL0YNHlEmz6YDt5UC6jxd/8KR
HBZzkEazSf97RaZ9ZojAz81uk4P7wWbUrrDzbAUg8YZnA8qSM4KDNVY1dkbFDjEX
qAYqseP5RZjUDOWJT4VypcebOSIRmYk6+AiFPEktu0LRZ3WV8n/pg6uEXCVyipEv
mgIadvTN2wqcTc7m+FnP03xLABf5LJDzv0ez7lLmjR0lIrogMJS4qpcMMq34D4ql
KSPWG76CeiO0sieO4Q5hYUf/YU33yOWVRgjFAHv1rz9NarfHPa6R/GHYdfYZ+jPY
bxhOWJuIOT/Kh2I5rd3EeL+pIneifi1BhQz0oJck6FrpNFTsDQuILisubFl+LY6o
MhcXFiZZ/LQCv2aseilJAPQcTyPsojWEdgqjaxq17NAKK17XR3plmV+rpRKf9Ova
wqHdk1OkA/Sx+3zyk7+uxo2vl1/fhqkQRvLAbykyUXboSvkVt+Vbef7UZ9Sw6xPA
SAKAPg4oeo2b2qNhYuxZxyfbr8q0KYYroIB41WaCjNkFaRu0C2X8sdsogWuQCSvl
QQHL0InBZgYwn8IfHlIahgzHXTGERET872kNCodRNfYqW8qBss+TEkxEK69hUCT0
d39fLyXD307VHHXiUSdXOKyA+XJ10COWbYdI3wX3ICnWUiQ9f5FB29IENm9fNcbo
+E+EWadE+90UV8XhBulCrvnhtfwUf9JETOCLizrR+smzgKCaqZkVw0KpAi+glozq
i4tLXpU/21ifZ+Pf52oQ+TCQ6xiITMhSNgxakiM/nJb2mryBpNKO6Z5Q4kDse821
fRoT7agiilvXaOI+AgSIzwJQ5xB1tjPjITBfIUUGd1S+JJXcel4KpTAb0W1yEfzn
hwlZmxDb8laGHPvDg2KER1ZX1BhPTrRpuke9N/TIqotkS9QsuG/9MTc135OnuPmF
xSlHBW4YdtGY0yrTjMLTV1gnaqMoU408XpLfv+n/m1Vu63Ut/KHxm5xi9+ZDeC/l
QP5komGRAktxNKetJeHZ06nGgQUFpbi3MCjymBlVMa9L1ipshkY9BpdjIU1DGiPQ
ELadBqnc8GK+KlXwWfrqHvIWNqqOF97WjQu4NpBSOXsMR5eK14v10yX76XEczvgr
AkNQ519i3QXfaAmk1xWpn5arJbGTeyLJBtlEOEGgwHTtTu4bzRRVpJMTDoEICNKy
LD6kYGvTe9nilRXkTWrDd7TCNr80stKN8SxOjuX08LcDUmvLXlIYhLZ2iGdaA69u
7U7jFH28h0//8AO+4A6jQmJhfgSFc1IUQvdD1Bb8N4CLCPQNhdgg1IzJM3dDdkW4
jrDWjlXxOgWFFJ5lhU2xtMdOZmrb0z4Z/Ss+YtCboNAQfr+kuqSXrGCUa3GRr63C
6CVaSMQ3lapZuAiMBz0lI7lVxrk+4iCvReBlRZtFGZnpBWM8J/bw2LmJ8FsLMvKk
1/LrWmrcla6IL61fB2yWNwQzx7fFQV36lKjdOqNtu3dl050WA8IgLE+XiibujgzP
01JbpUh9/VKKPjbZzxw+rtFc/SmwVPdUTW4ZH1Kz8VrtOAYYGruOeSe+x4dXIKi4
8FyE0xjYii9kmwCjsom+aou2vOW++njRAzThre+Un1t4VY6SiDpD8OgWp4pUTlIQ
TybFBMGkNy7SWcJNuavxCkHJ/VzhfCIp4sGeqdKpjvlY5ccwkSlLG1ccnvIWhw1i
ZGDYqCyke5SigZdXqZZFri5An7LHpaqdSG7H5FLbXq3jcBiuxi5U0Y9VB0/DWyQ9
pUS3NatNsxZmDv8JR/4F9DHsg7qmM03OP3HhH/bp1IqdgfWuTpDY58WYuVpnMq8J
dnzfYMAvVMSbVCc/fuJFfB6YPb1avLUHJgi1kq7UVazXZA/3yLYgcrllMC/h9YH6
6hrDJ1SUvMQVRv+H+V51xqzQ8KX4AMiIaPWszOQ1SqyLHWY3sbPWoEpY8z54225s
mk6a2MWsEXCqRowKBXiya41Dx1jpMF9wI5Q1nHRlFhXWvJhtLA4dumnXWr46Xjzj
DDZeSVTxew51W75tnNEhVgeuoyYb2Ur8esAvngcr2gteFQUNAR/cBoaSjS+oltYQ
qT6HfqyFjngo+4ii3Gq/wc9oI+IyakenaJ9BXp3/8zXHxpux1H5nnXlL+rRB9QkG
Bs4qlrBOebCoMRfjZRYXBUKp8ogMTLY7B1D8jWjSHqXvk+l0ulkpdAHMA7vmi/Ba
YcTEBOjGvmZ7QLSP75eGTx42GnvHQ3XJZKlmD6dAA0v4ebqfTuElLdCV0R3kFRa1
OdIFRRITTGyT1Ylfml9Vel40QsNSUrm0mT6XDYh1AHnnepLLiVZUsRaG2QwGdxqo
ng61EHHl7Iki+kBkNcSX+iTkCDvS0W62/cAlJQO6nxiS3j9rnQ2fcNNKYCrMPx52
75QUZrA3Zxroi70omQE79doKzLQOHFGpF4M6XKk62ONPt0dj5JveUU2jJGqvE9fc
hHSrfQmyclc7c0MvvkVbbSDoQ3oW4G/IHJ+kcBiKKjVGJko8aljqZy2l0p3fkgX9
o4/xVnL4e/0Gbe+v6T/t3LYFOSLPDI60C3Q5ROIOGWIB54EoyvPEIUE9ppO4kz2R
RvrkdrN/CMs5jP1ktzJi2WYMI+LsTcAsIvI2PYIgTVkV2yMA5xun/FENa4ffBsoJ
LlhtNcudtBxcEVAYFf4bVo+WBDhPOi6oyy0Vm1MwSj3s2Crir6aq6P86ghF8BAsx
nYt7XgK8XdDTGDGBTnDjiapW5MMP5C2NxjcrdRHXEYgznKGB1ASRhO9yfZui2f6t
6x627rdTE5Ba0jsaQkj72wECiZu8KAIWxJwbrvFfnqzObd1cOWgtP70bvQAOK5s3
hHsEJN9BzmUdKFdfgcstX/+jjznmNIQBeHi0c0fpPydH2kHhAcAoIDZsPzh2HIsu
DVB2G2AQKkj+/BgAnDkjibT6uITR06zcyD0hngr4ti53QHWZl1OL0ZE3r3+vHJNC
9S6TjnrxgjNbfO1Pr4cr5cpgMrW+swrUyKPxikJ/3ZptHgg+dtXJ3+y6CWix4ety
ZdJhpeZ+WrXXuBAm8OQN9BWcD3zxgYRBwootcFWGXDxG+PHExIghqIRiEWBG89sh
aTamXP3ZJb/m7t0ax9hnHor22AdKYzDm8SZ7nMYSs7caLoWGr79RDBz12VDRsC6/
W9JT+GdnqWe7AZtOcty0zax5M9KePSD4XCiMomn3GxlDtKITo3nVkTxMNmNWfX1e
xi7JI/SG+Bqq+/YyFQy8kOlHYu2j8RPrk/hSPpGXENtJ52o86GiUTCk2B5y6jE9R
UJwg2BOKUalMWCxDVPAKRyM3flc9FJzxPYX4pMa2PCTeVEvbcgAmE0CWETtgkA0v
COAY3gTKxVF8T7Y7G9tP5G7/5ohTcpHOI+nRgiah9LMA329PAyC1G9vHRtWwovtV
VfCrr/8djvGv2R/2zh76b2DEFYZJclepB5W8mYYQjBNr1DaJqnVUD7TBVoNRZvq+
o918l9sw+fKftoYphSxh3cW28cIAQ7Q7A5w6a3JaErkquGkwJBKhAL1Jto4dRZ7Q
HKn+Z9YT8nmm86rOyZerVbtlNRhCS+RajoyuHFjoC5Xl1s47qwAku/d1QhH7GrJu
Q+PPvSaUDMiqNzDXcg6IZmwJAV9/p/Z7yvFXf7tj5ADTCuj9txtbQSo5Z8ejtt/9
fynBCiY6LhB3LhvpLGnsfZqkhB7vLOOEkv3csgW/FIFvOtSMIk60XAiqpSORpQlB
dSWtpCZgGSzpHWRJrcNnR207OoQrzvolpfjnMQWXnPNRSenX2C12bxBiiPnFR7XX
0KBmTaaXGG+JocenJd2yKHqHn011Ve0gSXKxjW4bsoF/ydP4TFvmTsJEkHJedAJW
IfZqDCbHrIWp1XC8uz66eHaq6BDq4f7skbOpRcqn2fL3ytW0xwsio5G/7xRD+Y4f
G1PEhpuUaW9P8bz38AnhnxQ7jmHkweJu2KlJcL3CJHVfBGrBH6PaNgz/cV74byCf
/eVDBtYrorkYakw8mjcxL8wP55HXIljRNr01vbm+6MF/ipxRoVt6PrjKEc9yqoaB
9OTjeXzendZrVjAHTeHK/+lXesbrg7QTBV8gpvoKowQICsjlPZrtSaZIBD8kESy2
3OizU3sGBTeOjIN+me/Bt5m9BhXIygbhbKW0zMoMwyeNYsLLOCUKbI3nHrX8wMXr
KozQdcS/BFhdlY3s6ijmx787Swx+6BSLs0KHKyJbEtIWXRnpRhB8mYAQK/vF4+Dr
YDOeb1naFLk4qKfU+sZb+uEQeBeNPLPrIFqJZYz8pL9a0Gviqt376RKcmfwrQiW8
AIM1mBnCKxGzoRIbO1FzE8NS6yA5RAjrNV12RBn/WRKK2RIWXqZ6Eh6ZWJ+1Eq3Z
c6l0oB34af6Y1vZ9D1NKuSqSsxPzktvJCJ6K0x5JYlHgOofXYMxSqwH/AGIyQTYT
50NEfBaYboyut2gmDtf3v6wUXnA+iHJTnFjhOG5TE3CGgAyQfC6XKcQKv8Hlupmf
slv/wjMuTocLP/AgAzIXFU9m9SLUYMQpcGr5n7gHXeooTFdo4OLcBAldC8/cLAKh
2549cD0sLBsis7Ne361k42DGwzkX2LxR0JFA3eY2iQAeTiRaE73Br09MMOdgrS9H
947mnUkwr2PAw6YYKMIReKoxNUdLuU+wsYRl/capeaRA5Zhbsu9QCKV8Tqzwlrso
ihzP4yogEn9u0ypE+R10Dk/7/WPxneZTRPrupNE4mF9PS/90IPwXj0laiCkp88d2
/hcZMh4eBWZ8Aahz2xmTdio9iKl6t4N6RdPm+FPxmli740CNUXvyUqI3VVQOcjK8
zOcl73xQ4VR0pnj/Pt2+f7NkqhQV4VcRnnbMq9mUj9WIO7x2HS8A3scIiH1fecHo
k/xyzmYxQR1GisC22gbnYJe8l93R7W+KxU/i8RTvoOpWvhpbrsus/Iv12tO+vRKs
b6Dd7UnW0ivJHV3ilHxyz7URBCsrlPLDxmf0xrvUj42afXsbrsr9r2IYPJg3KF7n
0lZO8769ibDk5AWE5Qpj+x/mhVRZ0TPfzh2OwFLbiHPuqUTGvZP2L+yQEbc+d1Wu
Z9a81mk4SQXSf+IwTFPIMWiGeyVxS3+0MCb4IpO0IifctrXFaKu0aQAwyf9KZLXy
GBH8N0SDkJSEgkWhKQr0R/Zi6IuRgEk0mPSeIUZg+o9gdBPcZnrdTyZGQwJNuJod
ZDZVmTORmVyqvi2AhCZRuoFyZ55XXaoeBA0nfeszj4j1LLqKYTU021Sqlto+B7rA
e4Jef8I1Ie+mbGQp8+YMU/TbmtXeoDMBucFZN/5BXQu5L0d0ymOWW9s9lCnq4unF
RMbKmQF4SaMwWq3DA9+LWHFxBkS+4TEDcHW8C4dfoLEODdzZcwDXGtfJErb62Mzn
VsSOxOo77C470mkidOxpjbIqKAM00Z1NZ7oRsyPmOtKvP9WLrtzB1675kZJjPdeW
HT/8H2Q+Ox7HG126Y01V67Y/zE/cjqBrgC/u+C/6zRDDZvdnePSzQ1qdG61hJ6eM
78nf+//GbG89jRcfJjUXlijqrD1vKzi0kbnlIz3m9xfF/8m89wSnNJGx5wgRB4sh
eH6oeDgvccYiuBsKRNCe+vLZyfNujt4uWuZAvHQ7R/UgEylZ8WAhjxykSF0yXl8A
PAF/gr30V0bWgbee788UtDSnJlX7jxF2/0C9mqbjojrmaL4mRTKHITgAKFW7YRE/
EqQ+BAj6QVYv6uM2oAztMSa0YGDKFolD/6e5QwVTZsOikrJx3Qf8wOWjxqP17t6X
KwPwQYMlFLSsKaoHHbovW9CyedIGQYBKXEnPeXGwoBEIdnHNkTynxaWQIa4NgVXq
44CFJUnD35zKjwq23e/+DMjacz9ig8FwFCk2OmtQJgEI2UduYz0ssyHT+loKBz2A
yYCc5zqrgFUl7bhVA2uIemB+XpXYQmsM3NjXHrS599q3ZLfGWDlAEL5tzXSgGzE8
NwPRG/NlPW/iVXQSPNa/X6eUCsMBTkgbM0Vk0PTd52QLGfu/wSIm2JWs1oSp7l9X
3rOp8O8L0aUSjPWE7evQjjbwMnTYAhlMqKJqZ3s6OnmRykOd01o25Uv0ZKiW6XO3
3I0dir1hNDyNtrzem8tvQnBnwKV73av2S93Tku333diBe+MarTA98rRn36wjq5ht
o9oi3Q9AqC990nmmTm9H5UefgoqD2poT6cONe8J9RD+tAri2kkhkuR2I6RVeZ0Yk
u2LHN6yY7bQ6Hmak8MAP8fTzVivUrd4lzxABSRuak+gTJOPjnJLnR/CoiEtZZAPu
2RtO9M2DYfvZ9E+iFAJLN1YRU2PEgll4+CztiG0JR79ZjjNrLYlM9r+FZHO7Gr55
5I4936ZD9kFx83399f2gAIZYU5AFWv9dsPg4f/gyyaXK/7VbrL8XowmfjXitBEVw
EzmIYCnxmKxEnoR6Jw2cNe4AVVvuRox4BqdqTsazYwZ7VKJ7n+U2XN/z4XQ2z+rK
M/z1KT+3p+zx1MnpdgObrutSyR3eOvcX7OIA+hQFV4ihlv2p+iIq6SWr7cTSq6EN
N61+0b0TlnHNBederXcay/BisNyl8NhZ5mEJwqy7fNYr+NC/aIZDb7D8G/3VK5/z
a4QtPvC0CPBaGva4UdLUXvjfMN6p988ExzwRn/Uwq8aTzKHk/I2pK50bwPq/fJer
IIFXK9iEwEOwuznDVO+xlwox435+2YLrUq1JTM6K+UGo0Y6FyOqJVicidB8BSJuo
1IE4TXoAaDqfctcWV6u2c6KO3Mvop/f5ZzL/lu104acBoeNCRSysPNWPHPFnkuu4
WMiR4ZvdQxeGj1laABbYK/e60FHCbcYwCSpX3upfQfEQun4mr3dwQbuT5Xtd0dXU
myeRUYpanGgFtoVDKOGmQYOKOT7UT10oj2xVcS9GgIQfiZaeIHWQg863Oq+e3jeR
ZLmd3JZxevS9b18Abxdhv28gNvY6dEBz13LIdddyZ/1VF61QGxDgWYE0eErSVPoh
SVWuIT+QAHQ1CdVZjICAoX/Tfj7fyfLZvnh4Z/8+0PC2Sod/e6KRg2fcp735kPjN
fPm7a5XZmSKXQj0uTEYlbgUpaMt+Z457usrYfMisIYRZm3b6j+AR8EpM38H01x9z
3u36AoOqZfMCQNG34luRymMgGud11C5e0t4ZI5ovRgvahNcqPVfNyiaNgn8XNjvn
emiNKlTs8rte0jKy4Db1PW2h++9eOxkZUEov3q5XN7z/CHEr8c1OOlYK8nqrn1H2
1AcmAHdXRQEze8r4WqA2Ws361/q4IBooQ51L3ckzWRTCR9C3KrdnWkcq+dVvYx7G
0bEJHeVKut4Yn+tHdZB80xE1iCebINgOaTORZItZ6c2zbe/x9WBiXYlRdyD23NE9
AE14dpf7FCnlDU3JDwmpGOWDF7G3UzMxlr/gC5xwGBCO/XrjWDLfT4hY7N2exhu3
BfkWQCo1/li/JMqkPxGrQWKoHQxyt6WonNKI7yTQRlqFsMuZdlvbmArPJkiBN+IH
DZVs1dntNd6iQh/mBuT+SlGRb3UtX69EohBkzGRNokZyHrOFqGCeuJs2jmlTWGSg
0js/jEkwRjIuazhBTEpN5itNFIRWHO/R5BiAnqc17+oD1dNlr0e6fgEQ1aVt2YsP
UrI1jUWF3ItKnXiVIoX65e67vf8fw2txB3vyDnjZ663EMpMPRn1nbnUMq91S4hkq
hnIQRavw1jSrWDMjc0830XJy1tdV48Qba6hmLHUD9MJcoZQXc5pTCX4NBDd3lzDN
qSRQa9JBnI+ycHsnriC/5IfIcOy/ZCEtF/2yPVBicmeppxDi5eRMXTHqj3/7ungn
uRaJCybmo9na3X8/34bZRMn5hrFsxq1Fo2eLqPJXfp2A6rXq2wwKLyqB6E2K1Kud
q2CVT7DpOZFXbNgVHZX7VUt+S99oz76mICIEzD4sYtK0qgO7FojBq5v9/UkNiOG1
1SgneIdyJmixqb7YjhF8291egaIWEmv9kV6zvmyh2UcECmUnra8zlMjWRcAeDB+i
iuaiEWPavb18DuOGnHtZwGn4OsJ7bNphuQCCdiAS5zfTVqioifFlMTzEn7u47Iv5
IVtsvJssG4/7wq2Rx6LhqrtKBIATriR/wV418UemulQEclDDI3E/i7c77Ua3qiPF
T3EfON7x9nFYXYIPIhXxO6tFlc4TzaCJ06gWowFPGmv8m3SjsduFKZUMoUxpY2Cd
eI8iuVPNFHVtcqiiqA3YDVxtewRTSQm6P0ZsnVJo55XV9YOCt8mqWzIARSr3Ujcu
AK8dOU8jGK5PfsMKyppuIGal8FXv9+ln5CnlV710+uUQRrvD0Ol66e8IXcDylesD
6/EIq2ilSD1cV2ZdVPVbssqOX3Leni3hl2v6uKzZ5p8rk2mpulnkGcjBlc6KtG0m
CfaYRIMJpNkU2PVw3bjwlr7Fxzq4kx9KgN2S8PPWQr1jTnHi86aCN0izAX9mXeT9
kM4XaNLC7Hb4NsaZbRgFH4U49AtRavqMspvKXKSQQ0cgr4Eej1aAbKDmqPOwS+Z/
ZxKmvJrhTlesvNblSMh+oTW7n8Rem9zs5VelbvUuhPW58H+DWlDSfrlQSKc43T0z
tthij7+M5uJJdUB9F/EOkJK0KFdN09XOTN0gVEcrW2hxS4r6AkzxXMko8Vmbh1l4
sWIJAhreVWNL4PXUr8j4L7oQ9miojhXudsaBHdNxf+SASVnn/5WIN/9/7bpA7tAe
t+CRisD0nF6/5uSHdWwJtZ8WfOd3+xcsNAlPHDSDMvQSdCLeC0LcH8fJawCfbSIh
hj/XuYHhxsapORxOV79UWbywe8wytgSnSXdwXxfy2SnIdDcBU2fZd/iJokUTuMhb
95F7Vuk1F9TjrYxDl13qULDM2g/vAVC+8Og4GLjJ88ZSi5isS/99A3J31zrqI7Ry
wGM7x8T/mkLayjtdAZTg/PXBJd+IGH32M1cSst30zdsLlhxjsquZa3nLYOqKdOsD
y99Z+AUAmITdiLtTBmZ+mpoSmXOrI3ACg3qiSJ8wqUnwnx1ZEWXJ4zoynHggRg+0
gKftuwHl8HOKjltR8KRQZDGFJjUklWdARcJLrEJ7OoDCWaknj7SQMW4kmSn2rrmE
2durJ0d56fRAQZrXHJ5uaDshoTkg9gI7rB91LU+LrQVmwQ7lX748nz04aC9oT1Z4
B2jqywZ7GB3lwLTR3odM9Qd46DqiDO9vXoS1dk6tEFTizaRp3oaXfOF/yckYilBF
KICVmFcjs+4n7d7qdao7nkhcRvxVMzvrIIsLsFMAamyK91KR8kn52hlNfQChxFHX
GYqbdJi8BymxpX89n3URgCo2htDmy/W0KpXzwgcjilkgSQLmGW9uPHqDUtaRCzgW
xXhV+meqKqJnvODkLOei9I0eCg9idmzijOGcu4DxWuzh1OpqDfJMQvAnVC7/vrng
84V8XLWzlC5klbl8r2kBef4CW/z1ZIaimf0ah1Ys1taGKshcel0IapxKm7s/krpX
QrePWm+Au/1Wd9HQIAY09oICayDGKpekQp/7HcfB30baKEpETN6SnCF/mSGeaSsk
V5ETT9n2zs1ixARsLM3EAWED7B1qgbuuT7WBgbz2x0P7TSNFEslQEDr44b6kpLBp
zFHx5c0jsAawOhy1ErSRD/X/d1S5yYk8gYyXuGwI8pmlEGNKTWcbohknpgDgUTF9
gaHDFG7dlfLeMybg9oTldx9JoKgLK69QqAIwfq5BXPOMm55FSgfbtDzpwGWb1f5n
tdxytkQSsZexNfS10diwFx3k0ekSFPiqaNhTzfcDfGCps88QAA+VkFBZlPhPL+3J
R2IdNAvbnU5pQXte1WCrVORnKXQLg58KfzzU4tlWKZHjhb+46eymFWIGm+qv0Xgt
7i1x9g+STzEdpEgOWDZbg8LEUI0hgAHznmVRjT6NnQjVqXLB1xKoWC2E3ZZX68jP
ofbrsnjMR6RYiZT468L7TQ7K61f+E3dczAHzOQXbwx3M2A99ch7+ebV5g+85Xn4k
g1aAZVwHmuhGvRK166EEYOUjLH/lMrG6Vy8pwPUmghkSxXpAmD/KfABRGEGuAyGC
+4DrOIAIMDfXHdx9yrhm3ewmoCUnCJXoNgFHBaU2YyqUoUn3MFA0AWuqVEHhVWaJ
o5vcFaEu/E8XUez8qS0wbGJpi2czQOYyOM56x8W+F2YkwhetAn5UDOZY9Mudwd4T
ob9ibVkkCb46ZE+eMsZ5nEnMrCe54p+eQiFvCethU7r161dbqldblkEq0SqpLwqg
jwuGF7EPAkJLI4ntUT3AY4oO09+Ue95dsRcC7uZaETtSNRxYEGG4kUPtBHrbdvAa
ic0CaGmv07vICNULwYJlsrfK75BOM+G+JGRg8fZx0CtucB7qbIU0mQGwV35wl9WR
jMLoQie7N4UgK5FPrFKsFzcPH+Yh1Gnx0IYKJME6VwIiTlpfoZEY//4G97nOVcG2
UHch6nDvS1ySCEMPtTdsY8uFTPPuMXJ/HlQ27CBvEkKgWsZFlEyuy9apFWdKgVg2
K/qJt1dYpi3J5k/TVzAUrKWHhAf7gCVeCXPl9zh7Lag8aqc+hPDdC3VwcadfYhrR
nfVDPTafv/k2ZriJkq5LJaFMVp3eoY/DqXamOmrHs9Dh4EAWkssYDmA3BuTJxufA
k5nftgzdicm8bgjLtOtzka4/rWzXVKIssSpaV7sz91REVEi9cHHNi66veVOmhrHy
4KNiXq5iM6v9GYCAofaatCrYEAQjGVvpYr51VCXOijh4GcHYvaXODYOzI7K6ECKI
A0K0jqYpWR2GfyEC0X+ECfkowlNsFSF3zfjRb89vO1bdOzu4oT+HEoaQRYk07Psh
DNYwkYBGFWxs7gZDPY8HCOIFmhw7lq9IMJjwMs37aiTpY/fNJLW3VxnuLclPut1H
/wu/3MdXdOUc4vMwBTN9EYl1FVjWDIFSO0gqdMK8wgZc6YFvc1DuHbz2hlNIFwMn
lhs0wLN3drM6JZXLje1vHIUoWXYAf4h6S8oIsZmbT6ZMKibpBHfRMzGnY0ZNiK0k
eLXplbs0JaGa6NsrsPPn0OLVXbEzQPE5zT9mFpoFLv7kCVA8UTQQ2inx1Ya+UTtg
+UjHaJxHhBmAijyUBKsephBh/nR6eREvwjD1hdYwlqjXbZIVJRIL93TJWK3YA7tE
5efWisFLUUV8r5a6UzPYRbbfGn8se9bWLrCaxfgGB4pqU3LI40whFqaWjPNdmtlm
EpvaWxzdGFVX9Kcd8rDVQUbQvh0hgdmx8uZP+5VzpTsW8ZQ2fkl6j03+qpkHc7oW
f/smrJ7Ir0ATpArTtm9TZrYCLBZoyNrD5AYlOkaup9fc85rf/eMD8uzyS9uE+n0f
jSt2S1uxVbn+3GMYgy2MGZBMUfBfk96DiDAY812GT8XJRYg0TDpgOMQlP9EU07Oe
runUBwebmzQ9Ga7AMOo3kgTRPgGambQUA9P3aA10Y0BMLqUJnJceFJ+Sc/mnsCWr
WT1X70jxAfgRTMWu+mSWqETM2p7+ngW9doSCtnNU+Xrq2kVEmsbOmpAly5OY4Ei7
PemDivY/uLZh1e6lsQrr8ezKSiYWnKfkdCgbxJ/sf3I+pkKs9hiYV+a+3YNSUG84
Vip8nrKvG5z1f9bH+38s9wgTcoTzknlFg3MzmSKZLWaIPo+TClyDUVopL0j87NT7
763xcPQ96cgjymb5ed+IVz33ZSspLdEhwsCtC6R5yMcR/RrNcHVTCI7i8tLKjqnx
oYC+Aly3hkOc2Ru8xPrQpH5xvffj9Qu3iiLs+tCPcbuIwPXuatUcCpAcqfakZ3Tj
RxOnwRQE209q0DfO+XkUBWdkl7sNWsqMmgMMlTL57mtdhHfKhjeOuMqWZ7andKPx
y1bFA2yAhLb34SKuFVApUNWXcavAuSykrBXsgK8F8gfo1bQIXRFoXnJWmOe5SQYJ
KJ/jsKleorKjTnJ1/kXQxuKN+ZKfpfKFLYHHdrsGUN9CR6rgj9G0R2ggwEObMk9w
eAwvtx+XzRk0fgbJ50j7uUcoQMqrDGs4WiprEhqfaWQiGK9aekfcpDuBDdanMFwK
WOjZIZmuvl+oLMX4DegtwnDmZVm5yBwMdOVZSiNRBtGnPwTAor1lhp9U9Rx5TF49
Zne7a7+tAwwZvXyqav/y3aQF91gwu4dzYnqqnxWEg1rk8k4Z4je9ggnlYU2KAfGM
xRUI58djEBm2TYPffbI0ZRZ0amtQmGuXs/EOf0u2nL+Ll68IQFsT6QiPZ166/IuY
SbB7NK4y5hIr9wZy4ml2ca2vkrISwjSjsCrcG5z4uorOJEwUxJfBtWxqdgNAJO+y
D2Eqt+SJw12nD8UBBwfAfk/6miVH/dqrdYXN5qX0WLBgAtp+on7CYJn37sIa90Nd
s3zOlcxc/+tuM57nfMN8fZqFZSV9SnGYForkNhhcLwQxoRfNBhmetKllrHCo7RaH
Jg2HG6NilyojpV5XZx3POFQ9GuSCcG2PyUoatindUgAji0730CsoCpF0AYTi12Id
qMQW5k/Y9TsWvI3Z4NrLBMzCijMM8qFTL8wvCtrKZz7+Xk7AXJsbWYlIx0387hos
mnx3Sc3nPEtqqDSMTOfekyFsqM3IRc2taf7fDAhIBIzYLZyzHHOxrAuY+Mv2exos
Hfzwr58V9UrQ0fBuWHPpS8JC3YesBmTWFARRQ6E9DWuOD1A+YX0kh90iAQj36V3z
bx5LIVQ/npgc/BYkiML7zpSMTuuExhEU+qvITO+LqoGc4PoXupcNNza+sUBHUxMG
qab8+4Rj/yn4g98nhzFjRyZvYZMixKbdT3ASxyzNgDjtmyUVaYLoQNYyw0WTGJWP
/3vtxxGnrVZ4oAh+/XhKS+DGGR/yShuUIkoZ63ap7M/j9ho/Y6pxiQneblCEGIfd
hHq9K6detNw9u3jG8PeCYD/09ZmTGp+s5y9zPI3hBkUdFkS5w7ZL7cdrmcBwiXoG
vVxNNDIoSMcv6DHIB6jANhVJUp3gN1F0tiaYGolpTLkjy5uUjv1/m6ui9DbGP+Rc
G//PTYQGGXE5NR1cXFN0nC1nBD+afFDfNb5+3hZ2kcXx6nMoLxYqL8ear67uccbE
EnpML/dpaG1VU5U2S1/HAsohSrTA7yzXHX7StVJUe9cPBt25b7qb7svyyAo3f7lq
i+017vLI+pYHp6e61rXh8n+F5zt4ri2o5Rs5+mbyxzHMRWPmkdkLO1xinu5XOZJI
wMT3D2NQqhStt5wWlMGvhe32EDElmJkz4fhCz6CzlrcOxUMhugNdrev/GbV7Rne/
sWVVDSUB8E0YroxcdtUdmyMsgUHJ+h2TaiqYSP/sXOaxGnKCuZT0wIofF8upDlgY
RcTe0Kn8fVUOn+tcuA0dG7yUVH3RJJjaAmt9W71iR9mS8gg7M5gKHpDTASENBAa0
9mul2EDFpTXRx0g8kZEXsFvOGbB2A1y8RWTZODFL4N4tkY1j1Xm+4XuD3SkMsGPD
ORl2GMgbVUp/JAPa0Lr4fiql8GBhnVRsQ4ol74aTNwBPFi6kRMaA7y8nxZEDY2dY
PX0EEnR7o4oK/eYk94BVabl4TK5e1QnuqDDP1n238zaqehFUqEziTKSHHLax2G9T
XWMIKAYfwFgmrbNoeMG9pUgzItRPOtOc9Tb5SjMKYtM6TzPJHPlrF4L2OD02SaZ4
qdOYIAsJp/whcX7+jgjQM73Yin5jy0EIeGy0jIjsOKU2UM9gCFsYh723k8/oV6mf
SmR6CTwegA8n6fZ7mhcsvOFr4IDhRtfOM6JyoL0+fUjL2ZQMBVi2lP+EcLuKbc1M
WhBUf8EzzWqtRnM/Pts0lksyLgqpalMg90oXIJB282g14cMEyQmT/9B1ogttitPS
ksq2smY/0QcUdWjmMg5hVbWU2XeRt8XynZ1r6SBe7KXEDMJtg4JcQNkpqIZY4QFF
Us8zsON96KzLkt8ZZy3RbwcUGWHiolX7cjQuALwqqYgcBUBr6JA3bOs0NzlBHSGz
1AQpV9ZQMrBD4NJB59kRIzdnXmpeTkZxxrBCUdGq+vrW8WhmvOQF+V4qBq22NT4t
1709F2xZIy9lFQxk8flrL07zhIR3ezPsl37rXtujcPGdWdMbXIrXpDFyV4FbsOec
K617Svu4DWu/C/A6mQexb/Wx3DQ28UXfarkmkxrSUHhYAVy8tAGSWXiE8ekT+A+v
gm/jb+MsomxXlUXsh03dH55Akw4Vsc/mi34jjBLWO8UlLfA8t2qia2SllmXeXZN8
4MQJAIW/o3GaUTxvMo+QqGv9fUZNQA8v3nVN7bqNaA8UKCPnSOQNFDYIWB4x68e0
iSrtM7KJ1MJxWyhxe+8ylWsQVlx1ErgqXLWbXk6fPhXR95jYwscuhw/BbqtITeMv
VtGvPbB8D+IOSZQ+scmfyBf44Q+Bzzshh7BAo94DECqiLpHDooa9O9VcbH91n7Gg
O6puPHscHORURSI/JBytDy9DP2bcJU4fY5GNZqXIM6GpZFhAVBtdyvlEz3KTJDET
b3H/aGhHesa3QedMkeKaeDKn/fe3WM+CJaIIWX40n3P5iNFbzG927aeYyufu0FKV
jw8YmThXQWcwKgTH61VdUCSJGvn3xfdh3e/rWxCtaWvEQiIMQnwlA3eYxSvOBaVf
tqmdw5eEjcjATgEx2MCxUEi8krblO9rhnLZAfdIQldhNXAmMqyBqM76QDN/lwVZz
hGyNxNtRkivRC3xSA6xfvx0nVR6MzVWyE3RiMOWeC63rcpO+5pR6VA97nKHN8GST
+DScoDtAzHtvb4LzplzfKfi4+4AlOKx3hG/UmQuYlUFQ5iDUPaLkcl1bJrtrx0wW
zYwvKlABqR5Nt9HtZw0qJdkDA6R1eeZ6bv3bLqfXHwnJOkk8StpAI5THQJL+njss
qPwayAUSTsfgt1eup8orNDbIr26Gbhd+KVZLUYdyVIwVOWT11SJGFYH216j7DDjF
S8h5IqH5QGXUiBgXp6/acd7qKmhWtqBROpZEJiunTY3Epk6rUjaWrZ2wQPmcorxQ
+RUtaJXczvgaWhQIrhQpoaanvJdgP1WZl2vCU6TcdsPXaFgSLHuylOPqix4m0UGj
n8vwDSkC73bVi34syIEICqr3k53cm8iH0Uq8VvlpltdKMkYvXZGvP0nXwMC9nEYh
+C5DCpDKobZ9jNd/LQtPKdEbr+P7OVrGxi4aD+OimKLKiPitzKiFraDFsY3E7Wlb
I3AO0J8FGEr2Qme7kUdX439eucqv+rJlaqTgJmRWLUhbW4bYQtnQkDthVBHWfvxO
8Ye+NGy7tYlOiiM7gWlHz+Xuzwmw1FBO3+vrbXX3UEBHwlDEQpV7qCUQqs5PctfH
9ZKJ/85EXMU7agjUmIB90Mq0HF4BRYpb7KddQfvOcfkqytpWrYmIyu4kvbNGS1oW
rqb1Mqs02JEZxvEJ9kuxz7p3hVsh7hrWksK8vhb+gvVZAdI91kwS4lfLA/sF9nEx
dMPk8VE5CRdrngwkDkR6JR0pIvV2K5Syc2paQWquFxUeKR7nQpa/HUzwp3faV/lt
SPappbpAmC13KYY3UtLw9998RgVmtLm7BThxXEWzBnannyTd/bSZr24v6+Z4yPO8
dhRdAU3pm5hTu0CWPn0vMVI7G6Jel7Ju60WgCRpaZg/GP8z/uxD6ZRykQMSZRLwu
GM3JzwEheSN4FMUE9II+3sxqVff4sA12ykDAoP5a+3QqjADhA9wS95e+M5P/rZfy
ZRSXqMhsuPO+ZoiHfBqyDF2fkEQywo9cei2mTOd415tfAV0SfoSicEsjaiyGUCy8
vJ3AgPoBGHpFRFM4k1PS7t4n94n2f+WycVrQXmCHRW9VVx4pGh7Xhzcir15qIV5a
07Ee1Ei2IHGwQV65inGEf4+N16lKdiJ+jjsrcZ0g/pOUIDGagLTSVsv6ejpnu8we
6RqriOLC85OqsdLKhYg2CxHMKnRJ+UAe1qA1v1Gf+4LctdKK+RBc9XCh6XGculYA
AR2j2xrmQLxMhyOncYQPiUkIGbGrYtKgIX3lR/Hh/drVYSODHH5sxkCIsBWPKh8t
tXKWd8B/VZiaW0Bf1biuYMVQBpZIesOUsdlaBkjlM0ABD15MMZndUDifYRNnGsBo
jzCoRHdb3vUHR5Dz2EsbfJM0YECXSyI+pjydmZBGIbOwInofWCyW/2sxiz3mho38
xFj6syC5VilyB9+TspDd2N++M1EtVnekMD1QDPiIHTQwMXAHl8oD/0S5ElE6aDnt
rjS/Zsj/Zsyn6Fwzejz/hTTmgq7pp7BMIfg/xvWH4lP8cwKlVmYZw3a4AskOShhH
hADqdxY6B0O0aLIMPyaJsLcsiN/vXRosFboBhmVpbZwq4H3vv3F2FYOy/ZN//aUl
q8SDWTTtMA3c75YnkK437CmItkJzcTfdtkiKSCz1cK+VZYrmjQOa2MidxPOenIn8
aWDW/yOqnJKYYf/AR+RqNvd4deXRdSnmGPpTZb1Ls1Csz/M4vVR/zeLS2mW/36gR
iAGAv9oTT8gLDwcTEJZCh9RkqKKBdOyo6+GA0IaKKsrYWrGILdZb2crAjTjknY3+
kI2/Xh/HX1/M2Z5FS6bgBJm/ds82+MCVIiV5RCzIjJs0Q/gC4j3nkicApHuIzHUF
bM9r1OYhKHraxZI6nF9NupBa9wBe1t7sQAwWKUJU+I70PHimV4uJtpwq0y+5OJXj
NYuzCeDDKXRHjGbFfMHGvE63K4dt/MqAv9T03z9SfNMCTWxaZsSgeDD8l21LtIEw
nqh9B9d+pDzbiTWRUaDfOpyABuFGZBidj9+epmuT7xAGM4JXNfzryqWt+e9ur41H
8t7+ZrVdawRdT9aYdaczLlkQVClF64jO2RUlXMMWLhOoK/eg+cnrXmo35X82tVHC
6CSCLxsUtZ9vsTxs9pZh/qmOG/p65iW0UxQVJo/GP+KbGqJ62SslEDrRXXN6l3jj
SjH69hhpoiiSBfQDYeUDdBk9JhuQx5ubkgPPiMMM9ExRyjffCMgs4S5rrqYBwzeW
5FoQURnSMyi4pfqgBbyMDKvpTraIa5bfqQbm2d8yfEMelAWoLeqiMch6yX32wfGY
+bAPi8ZsQgQBkk5LV7v1NV8ve0uzfk21BWp5ZEu+04utaBVj+lSAuk4Tfy+2fz4D
Gv2kivwEXCCJNaV+0YckMBnNbUsuMAh3MlhHPoBZi0B785hu0z/5JkhRD9Nb0k5z
y45Soj0/B2DWqbdbPo607I4W1Otdd3+kDRQN8ABknFnR3O0rr3qv3IoUd18Q45Qg
1DDhCsu7rIN7p3OGThW0BE38KFVHSjdwSBNbSYH50YfeF1sthrH3pJFJzpoS7hWI
QNyp+Dsd2whYOEZWr0lJFHFVPp5F3NCa0/kwgbmcV2G15NwgVeBzuAW0hWE5nF8A
//thx9t+3keF7V4mrpHCSaXykxNR2yzwUfL4xRUFJzpUbyq8sy0XVRrmWelg9E5p
FxIzdohxpFA2Ex9ijphj20dKJYU7fHp9cD/40P57axu2PGtbaxzvKbPxs/oOxzSU
VEmkSw56eZg63gGyYgbgQQiDHjDMqDd7su8wyj72OGm4B5JeJhqEMO5kC0UMvAIU
8neltkM8ljjkbxahh/lZxIeI463HTLi3XIFXmHurQKa82kal5dgDBiP5jlCEWSjX
YaR52lK7j7i67AZlQXaCuCwd777agX+sN3iL5PLWAiFEspoo1fTUWGOFNFSz376F
WHgtlII+2wa54g5ENUy46CTRJYNXPZEAzfzZu5y2PJx/HkWllh9YrYGkGGA2YU59
dZMWS8o+AFllTlaDHvGU0KP6hkPgBmwgpU1YV94ZKFnCPUY7EHo/MAFL805vQNOd
7nCeRO7Egj4jsv1+BDZ7X638+06dcS+K59cmi+9cHtMnUyBLLUcjel+Z3xf7QLed
8QD2ewvzFOVPPgYFO9yDyBaJjfoGB8EH+1nYQtmLrT5BgFSmbj7nxCls2nQ+u+lb
zlEbcf7tYDxFc2h00Blq6bmA24thNjLKaHvLMzkiSNE99V18LZU5dWqCIeW6vvj7
pCwIbfKSyD9jowZTCVB5cHni6L7rF6o49n9ILQZkEg7C/BU5Zw5yG5ZanbNqAoN1
7bpFvuBNEDI+j9wwOHMgXR5bZ3gYmGTjx0NaQu77H72ipyv/HkC1s5Lbo3Mz70/6
ST/TTOvhBbXTki9ZHtnd8CSJRzS44nSvl87jd0/jmwWd60GobjWlJV/ZCHhA9+VR
zWcnZVrmDgClVgsagu+MZtG1UYN9uknAZVBErICvZhuFDDjqKw40ORxlGeMAmb/A
8wGgIVDq10k5TtaKiZsPGZ/gBGKy2aK8Dl91QXNG7fAY3DhPsaB9ikN6TkgCCZDB
aGhNaZ/6mErKllMPteCPoNwvtYYxhnN4GaRHKTwlZ5l0VmhhbQdTvxs1Sz/fPffm
VDblvBVtpjSdROsZpdUnhU88FGQG0yebFQNbINRt5h3aePzG+VwoCf42JWMAzUpA
H4N8PTJs4Dvqydvj/9u+JQU9Btil9i4q5erRGzDhNuIKZPFk73EyJ1/GLibSoAT2
B9hWK92xLtZUgBv23azh4Zc74AKzFdTfQ96A7E96Hx4/IqU7wt1Xr446EGf8vUJT
eNNtBPREkbLPfDGyQmDdfjLZLlHe83oIaHeguSdW9yb39jjy3w+L46BfKaPi7P0Z
VnZVwAQjDNN/jMsLvjh1Vec3xxfwyAMU2zGIS5rzUAZUCZkBLc+DlaWjxNhTm7LN
XeA9OAbzqu+CLT75jVkBmyBnaEk3aQc2/pI0UU4E5zpf4OgoRp3yP4pjVdW/FAvN
1FESryH3pw7I7pUurIZCUGKpxv+9aajDzGBmAdKjymxcwjXNBWpd2RAVLDZsmdF+
Rb2z1pOh44O3QFTkgqCC+eri/MpJKmsw7lY0CXdSsENvqpzfoDMZD3+5gnEgiIxf
QMxEMYnclTeSghWgtER1jRLHe98Y99gnprDFNNkceuvqDVql7W8l+LTh2OwlY6or
JLIaqvbPbb75CZL/TIluFHiLKiVhr/dPJb0SulK1/KEHDJPhA2s/cKVp6pRIUDFQ
RrTANPduIIcm20jvIwCPBRB76E+yaBmUmEr23hJD8woDjSfn9r/4QpJjmWNjGhxS
boVkjFtfWr23kq7u3gLkj5pfUY4ShnGPWWiU6T0mRmvOeaafa3r+Sbw6hsD4nM7V
GGel6B9w8tp0jQ24Ik39EaST5pa0GWbfw84E5aqY0DGh8G9OE3/ryB6hObRPm6K9
JMmguHPAAmgMXtwm+4YEsQ1si31zg1Xk/4GZ/h0aAoehfjarM7WKthK9ZkAw73xp
efQkEjL/I/ps42bU7VU6p3krUYZ98zFL81BHemIzMq3UKqxNm4tnkPsvHj4XdQQX
juxZjoTP4sno3aM53eNfy6i1BfQfKKz6w5xFVqLMJpJq6j05nrdFPwnH/8SIGFnX
+WTI5ccG0eJxWS8QCozu08HWcxqrQ4rVx0NOUG0zm+Q+R5ncJHXnAcm1w4wiK7EI
LO5PikIlppTIOBm1OkNKtM358sJr9eSuV8sK17eQQUUTwhAASjtRIeXFzeHBW/ME
NFgNw2FGrhNAmZolu/dNt2CHsYvKYQfAwaZpeSCvaYzVQumbWdek+BXK2YUnV7PT
wNKx3s2jf05nVGtE2LRk3TYKz0PlNWcsg3fklRSxt104+A10Qkc7IIk9glG7Vtj3
AGoUirO4ML5Nm3VMHA5MCK00pXw5brrHPhQ+cwaU5On+dIew2JbmgIiYxz7Dltds
PnLsDZACpQZExBzn0kbANLz8whWl/JLEZxzCdTVU6TQ5yjw90alWx9NCyQn8dbjW
o98Mcdy4xW3v6Iv4ClhHBAQuVt/fmSj84S9UeQAxuX/m5eUCUI3oz8n5StZLpzV0
zmMDPakpRP/u4vGhT0oVZXZeCnIgmAQqSCn7fuQRBLI93B2Rj5rmEjdoiECzKHzg
+XMEbPqSQE28j/jo6hX8yFfyWPxQct5OxY3JNnt87pAWxL7OqqY0YzGs9qGClDjO
wS6EZqM0M+ApQXMugIIA90bhtQ0yDFTR8GlEFQo5PtkCwAdsuYrtfWJx/ZShAYyr
+VsIqAchZMeavpmulEz4JIAxIcWjHX9DjakDoLioyU0ekwSQZrZzsmChxfAbvOV7
k7s+hkBPhJOP4agOW4H05sKpJeQHyA3LF14pjocfDFbXqAbX9EwMJXfKIVRmGUDe
TlqzUdwFr5CWVe4qUwKu0iKnUctTJem8kNqxV1t+fmvfUkGvJrh/cGg2fqgQ2hhY
0pFILpH4b1Rps7HSXXa91cRYNkAATLfRNSrTKmIAWApeiEibheC8HTJwSg0Bx1iB
DIXfriXkLWkbGD5FA/XXG0opbJFhvXTKqYJUrhgbBZnwGLMt34+HjZx2QgAprpo5
Hn2VZuEx2B31etTMTApfN1VQ4YaZ/ahj1VOoqguOzl8ma40Vt7zg23jKiyuVWZFy
1ea1lLjBHMNy/7nW7OTw7M2xqwlZWioxu5QBHxBB0CIymiQ4o28ta6kvkBPm0Dpr
5Mofi9XE0z6hEXMRJQUU8kxYWA3VMuNv4wfJTAlO420TL8dv9eUNIPThKH2uJ2xw
D3EfygAz7drlPOeEcpzFuDsqEUiXGFBpr6NK6TpSjeT4Uo6HfNBl2zVI9mepERRS
x8EWIaHI0Swzhz2LPKIXnPtynWKAe3FZnTKY1cuH+bXWn5rJOmppavTFgkhMrHf9
ub91slUOfAun55Tkyq6vkoe16Cpy/1WPT+uDf3Ip0dtPxcpv6CK1QRjDtp6aU6Rg
gmOkq+N0dIBZ3B4oVdkPXpnIMPZ5LfXB2qEfav8wsjzNtT7HeIRQKEJ3grmL+yv/
jmhBC7+NuhZi0f+17PdeHImiPSvjkHowXrKa1Jco7yEAYDwieR+uBDKj92fjjiOm
LkISmvqxp3AQ1WAx9Lg0pJtKmvm3Qryx5Eh0w2gBF09F7pQsWMO5sZFKDma16d0s
FFO2H6ehC0Y8V4dafCsjzN4K19MUlFysS/niT9G5FgjS9reOJhA1pAuAadxnRKBQ
LBOTdVNFkvy6P3kIInBYXVMzADSQE++eoxIkzMjnCUY9vcanTBpv26FH34jvrn2N
llzlwcIAv/z5pzc4609dBvMFNd29sfNojFo/+bEy4+c24KkrtIheB2AU8XPE4XsH
tZHqSRe4qL5HWf2fx5RRk4YjTfOvSseZJpTWZCYg1AHMzCSJw6C8dL+n/rIL3tFL
1CRaJGsoer53vaDXnBkY1vxj57hzKPhRxleLJ+lCpHQobAKCwNAXHNCyNwScYGx8
UyEQYDwhzYKvmrqdt1F3qG7UkmASVfVumYg5SKn277oH8ZW9HWYuFUFK1YIP2SbD
aBoewfBMoYjltAmqB9zRJXeC4SbClO5EDDQKe8P793B2cSK8ru2T+1J2t0Dg1X2g
n1Zo9yYrvOcNS5iNRuINn6X9/KUSm7cxHKqoKdTUHo4HAS86GQ56oCIIUP1CDTml
NMxIBR7NUkIBZt8JFIgN13M974tFIWCjexebz2rebZC1Nz1lKqW79dX37j6hJiKl
8tyXPFyFXt2TKzhPemf2cqdqCVfwETTtTgs40ZXhCC+2gr7tDFVpqcwmU0TVW9u7
OjyfuGUzxfNy7S7XvCNc2HNIJxX948tF1wNbSsbl1twzwiP7TOouqcRXhIdkcAbS
FbC+tTaoRiMVx2PGcaXi/NnnkuBF8cm9cs6BeXspsjCuynLu4y4j/OKi/xbwxrlr
730Ai+S+P00vjxO659WCifnEynastDrtVL8mY5qo5iReToPUngt6Rt4UHiugEHr5
FAXP4TtltiEODN7GclvGDl0P1++8rYX2sTHJ6XTSq6Mgca861U4kNVTGOrZr9cBQ
koeOWx8AlEno316Zcx88MQl8BEXcFxK8nzuiz/9ovXolamNmQ3NOOmBG3nrThyGM
YKcPa/Bq9WHi2rv74lzNejkGzCKaqfOivZ0XMqpdATrQ+WaRERL05s3Tyd1afVc3
ADN801sESoax+J7sNurKDDatQbnuuzQPrTuJgsxKCQhAkiUhCEetioTHwFDISjaZ
sq/yDE1QwXBBo0Q3iUkxln8s/xYQmAvqf/gcmjIpIlosrMOLb6tu2TyIwrQvWNWP
G9A8B+lyEluqlEJcqFs36+Su2PYFu8053VzDYKUw1uqifUksxn7bE4pO7VTUSw/W
A7gjytOHe9NZvpB69nOl8Ic8s730dhiQliSgA8a7PCjkQZAJ/JeXaaMoyZikNQLC
3B48zKAKXS+9WmqXaaVmtT0BHnnZn/Tqnf7D2gVNXKDCfojo53+NiCGrXLqIej8C
Sif7A8J5yyDGBuBSLX0veRS3b/QFot6WKpjlwvjyXAjVyVRv36KKNikNueGjK9oA
RFHbetExcWVvjqt00zxvFvOf12stUAmC/7smUXELqPt8gY4mvaeHmqFJtFtiWD8f
EHcEgjKuRiGCfZ7VLgN6thW1d82GZIKow/G+y7FLNHOP3wX6FLpA1c/kK/TJPyvC
545NJE5wRWaNsqYX7oR11ou4Dl+CqK0nwWI4KLrWG6nRASDiie8POFnJWJmVxsJn
wqvWHzZDws9FuYWhFEWfd8gBiQCOX03EVoRjkJxJfLF7bE26hbdNK5itIvcwG1xP
b9u/EpEo6ReofA1CyYE7IxN/Lx+22ODgdFCInkdU7lqnefapz0qMuAmGV6/FZtKl
6sCsVXN+/ynPy2PCTJVMTp/BRkQfQShzuPBt81YSbdfVKzv/g3VYYtatKpCtVsp2
s9+33gwvHoTTRkdYWVGepZOvmpJDGME5XUg3EnzjN2hGK0tYUk4+B6edm0um/W3A
T83tLfN619JzxsaxVPj/Zkq7nBc4uosvTWU6sEVmh+27CqoISWmEeqk8eRy5AcDW
1UlnNufsMNOM4nNShlbZuQxgcC+xhHNKOHBKIFvDyL4Htw/X57SM2DFIvX3WK8Ur
GTPchC+Dgb33fgS8ZBjbLKJGZCslp2uK9oX916c4TQXHvfaYw83ae35x0wCZpCtY
b29baimYO00m/g40sPt1sqG2cY8M8/260wQ+m/0KHXW5KnfYMoX1kVn3AObejKGn
E5tYOqnWIVedegHBcJnwvt+/g5KvGmpOSmWcpkEFKHb1IOkgjbiBAUYMGTWRJT4+
dYS4phqpi3gegZK/B6ihVsvtDcRYMyieKsh5LOws9esTDU3/VAnE4uWBd3GTCBX2
scHwcM8IdKWVLQK08aqIxJKB9D1L0AyUtkeAjvxDjcUgJozjv3m1JVl4z472U1zP
E+ZdpoieKd0mBPbydEkketzt7D2jB1BZAQDpDEgSexRjfF6Lyb6sH32XMAKvHdCG
e+1r5P0krJPEWaabW6IGJIqc5RW1PCgZRc3gGKhVA956k/o1iJkCdraLU8RRozor
zqp6A4EeZXcvogtK6j2pa195BtugHKWTHv0q+86vas/2GgJkgtjVP3nroiGk0392
Sstq3MLU5H6LnRj82ILWlv6QkE+lXJnJT51Mja2SRJ+EU5O9T6kYBaj95JwXZmzD
2qXM1XpkNT38hRblaZCujti32J7weo86Esz5Hr8+QBW2v6wvTMBIFzWQr/W1/syn
5+u4awz5tIUUU/ZKVGlr6jA+VQWFgZ2HxkrxknjR1qTOXz6DTAN+X/DaFvcNjpPS
Rz55rN0xEV/jgM83g/L4b49u6Kp+fKZM8HP1NCXzeZkx2lRNKflQvno3/JCSEqSe
13//tA20ab/EfYwtrBI/y4CwOQA8D6R875I/yP3i/b0y7/qoQ7kgZb3Z9mWqqQBN
rV13XiKzG7IczfTD2Vc71FhIKKc3Xn06UosU050sA52NFDRlcl09/ieJNFQgwcJP
1eVyNW2QDQ/KXemZ6uMyqVp3x1srYR6CmH5eTxZDAv/7I43bGMXTted/xtGE8gpn
vwFHWqk+T/vCWAxIPmdNogupSQi2vOr5agtHi4NfpYZP092l+q63t+wti4MJF+K9
VQdZzzrlRoTfouquTDS3pADIPiJZDWOQJ7ll887hIoEPiF60bdUF33HB30338CNm
bVPjPR5ThQWsjAlADcO6uZQGwg8GfipeEPezyasYMLlHWQ7PjBWPxfhuee+L6YoM
nk8j0UqsipdfM6qqWBep40ivBJpOiFvncCGA6gq9bYhaaS/cgn3xL4DTXOra4srT
Hyd7TEtBXk0sSQPeMEEzn5cy18iu0/+F6/hRt5nDxr2vyBo9d3RRzO0yqn7ZPNdL
nvQonFuy/k8F+2YBtjbiKfwQ86oXCUt6WH13YWzZSstpT1ZiadKiaLeLK9rneMj/
KmSbD8lZikdTlT8oo10CYdHAa83cnvlBSKQ/EGOaF+XJUFaszktoVDTeNbgWeH5M
FuBV39Ezdq70EQ8WbohcIKkskraEyF0+0eDLRWArpWnM8ZiaIAGjsYYUWgFRB2P1
j75Xi8Emd1mDiOuYRMLUJ9vR0jXNpdds7KwgyNeNDco9Fl7S0aDRk3/VAb9oGA0K
Qet8nIJIdQ6bFfzCF9EomuHrBbCJHMcw8MR7xlGeupfn+0ybBgjci7Zv0FqQnNbj
5pUtmbM2ChdA/SAoB7IhXn663sRL+/JpQ3jrOu+pfFaqpCYEXZiZ6DnvXV2fkzyl
jLDEyBmpwihYMjGpaWXJ4TIW9U6TAqfEvFfY2dHJR1jAfwbzGVCWr2Orw003b9qO
BciDfA0BfwZ7Y626GYx1/Aq75MF26v1vHvsKpX1O3TOECI8zbNKqWaiS6m4yRT9x
4bXFWg88aMTU98HbHF4x38EgGxHph5kj386C0Qkkc5sRyCjNltuAmg8LowBiLG0Q
dByVJPCCw3lMJ9g2dHkQi/8H1iJ4VeTWFCQB7p7cqU5Vgsx3Jps3gn8moyUWpsb5
X3XYzbOLXJeSoJCGs8fApH0so0uqWjv3qWI86joGCqpNp0aqHZjBh0qjhXlmZwtU
dZ2gtYQjhswQzcEAGWzX7sOU6w26dWVcL/izEPhkfgXwl56/0asi/xic7+yA4wHI
0C1oSHRHcTMdSWfgIUmIzFCsmj5h0n4b4EAVF3H/op5OwjDGljiVOdBfDOHeihxQ
2iyecmXO6vjPLzMAQiNZ0g0LJdNKzeSBOfvZiaRd+y85EWOdEnfBfmnyV+xnR+XB
5ze5450/9rokKL2CFPZQCciQ0rMO0gWKgidfSFND7M7rmrtQDplVyzj2nCYo6CNC
M3r0YWnqKmvY4ay+nC5BozS2BAGzbNqPMVEpA0uDaJUHBtEf+1/dghiENFQVpTN+
YSK2GVk4l128RLZ29H411sOJyKdql3S3bSwE7yhwEpHcQm40FGBmU2CqWJyaEfP5
SiCLjHtbMESAojhZHp4aOcuPoKES4XkV4lXdCbuguJtdjIei+0Dddq/5EXYh9eGm
4dstG65Q8kNqSH23KvARKtxBQYs3ln0pAefjQ2N9fpdX5+jm/oPhUc2V/YQ3Syzn
gpMwlJxrP9x8fuoH158P90ISWxfbm/OhxI05mKxCirQ/3OKr+hZbXI+KMliLMFFW
cfQzfU0TYvmc4St7MkGIxCZV/AkIWjut31jPTh4qQdd67Bbl16fnSrJV4hIZksqw
NdJNdw9gJP8Kjw07/p6DaIvuR++M4xmn7C5IzPnQcz6bMIb9spLzXPSZGCm5bC2g
nyjaLckLH1mYMj5hkSn2yVxtKyOzqOh7dZsOMxmyOAgYlnxtPehOpZiE1Zew7X/s
WnSg7rraIjDx2sifMTtQfK5xdsF8z53kDm/yPrdmXwigan1+q5ipHBpbxVnQVH7K
V6U0hFZXeaBGnoh2uQUjkyWE5caiVvnrs5Yt1eY+TRA72qH92OvE/SmmQn06JOWo
DFz/4XFC7aAuQase3rwP9vIxighHk+aQ8m+P8aTD8f4H6VBFPQ6rufc8xnT2twu9
Igj74hms3S2q55ov239HyDR0cjg7m44a1ZxAzjnMHER+4W2Mw55qFnwH1pLKJEyp
rxxykfPjuyT8NDqdNHZxLx4FJ26clu3D2VUtsS6Ltb54KgghHuFG3nkwn9b0hpn7
PubBZ1d1M68UX7vfi0G7BbpYopttIld7jQTgxMGV6dZb/26Oi18lXTmNFIl6Tw/c
VzGZHm7r5c1v8vONpwA3HfCQ/6ehBirAB5j1GSxHf/RJu8A1n07F/6ZpuWr+40N2
g2mVII7RR3ioIA9raWgukMeOd4YNoB3ebNMNxOSA3HTamxS32qAauD6+R/z1/UyP
ZBTokG3B+f4osWPtC+lSgtDn83XEyaPtB5nVUcLVWg820BciJOg9v5GXUhGx+qLO
FryLwb5tWzubPGqU6PHBnH0W+ElB8d1Xv4QzMh40iQMmHUZBSO/imGuPGJXfi2PI
BlJJoMp6imi55CnJNTEMUr0s+V192zuXsdMmZeSfvQSmKhmMBBWRGGofbyVsSdhm
zcxHM+LL63TofIoYtrw6AQghPhg+0gWCp1kTH6wydiM0unMTqmiNEtA0wkjoiKVW
IicEV7jiMjhn+TaeYCPbe0Q5BHCAUWtnX92EiLyrJinKYhGZs2a9wWkT9ysZlogc
sOVdzdw5vnAhRb/USDduQye6ZID/rTn6sQ4jzZ6lQmFyGE+LQmZUM6v4LAAYKyCx
vkbty8tPMv0NehnyCvJLgLPaf2sK1M1bsE70r5Kxz52Z+gMPdsIrbXs9khxCRBm2
yWlRZhJZ8aJK9Xc089h7JUIxn+mjPbDN3eSUPBfRfmqq5/AJWScC73vNE3YejI3g
qfL/djsyQvnqhyAQZQGEF54ZjMjW6DiVhi3FKtbz0Y6KU5bxnNScawKvUwUk9Mmf
wbI0E0OfwjD0U0K7efvWV6lOtBj74bAEN4SxBGRkOcNUhouvPYco7HgmLmagFphD
/wzuoU6Y1ilw3tFOHoK8i40UBuWw3UGzjlqC9ghd3t1AxjcL7NcX2c3DOD+8VntJ
9Agb09yK3AIMwkuNgRtGWFTKBpWO9eoueS6i4ZxARpdj3ZupBSA9CUuADsC2IieF
1vVjoDuDjCGUFg4bLzg/7Vraku5INjRI7bOCJnpz3dzjzfU2Lu+8ddKCVV60wwTc
K4qHfSHTBebNSN/aRmYsVBJqd62H5MNc40tdgYjnuC7OvjncHfQ/qgLF/FPQwLmn
Bw5htU0dU2pG/5RWCsD7A0E80LxVPhjLuZ4bq3K7OARwirumF6t9Z49Dl5Dd79DJ
vlqZsNvFNkYG4gQEpPADcTv3uSZudBRinxtm+CwMEN2r1b4IIiOoeshw451ztmeP
6a8sdevFxOeDYEFzHNmu0Rpfgls2jVlSlDlFpWzDFAk/Da9mbSIaDsgolT3LabFA
BLZIw6ivpWAn1uyQzTGUysbpCoFIffXkFPJj49yOqVA1jjVxDcLNXTLVeV+gJMPu
ltIedubbuwrxUcthiaWBWp6MEvXUsxI7dZj3u5l1PFOAFQ31S061vhkLAdRMhHYZ
yWb9qlKuX/mxONHFP7wZ84pxvI5ApjwyjMh8BCMtNuzna6N09TXMfYx76S2F2ExA
qnxprfsB6+2/j1Q0ClkGZAuN7+4tZKP/69Luemqol+ZzF9xfSxoS3kNHfC+zeLnj
a4mXTXgRccpGapRDPQNOqDAd2PpcCYch8Iquqmim/+zJJakQMrUKrv9xkr7Q62GD
/pzUFnC3BFRirznOyuLmFD+dUMZCNLR7nTBgZ7yB6fGTLdraaMVr00wP9FJ6DXIt
XE50DZNGo6o5XDbnQ4c1Gy7yKFFjL7sK0fUwHYXIVK7qBLhXMcyvE8TzHMP79moV
hbAdt9T3xGao6KtwiBxYAyHwD5ZFobAn6J0R9cH6BcNQ5j4YxYN9sgXQFucDM/Ki
FF3OkfvFMT6yISQWAWPr+sY/FYVElVzodePsT8YF9JWumOM5qBDTWB0XK4lxzD2B
SU6FjbfhdyvGcD5OpUxa416cXd7l7hcHpdIrHnWrG7D/6pqjzYR9DLXCDcaphRXu
V8qijsmdLlF0tJOeRH4+lwHZ4zlFVghj5fkeQRTjbHwIS7zcFQM8dQDpDBn0hJed
l2uSU9wQdcr2a5yboaXEzUAtN/oCG8luJAC4nm9aMmz/1daJi2J8v9DL+yr37adO
AU1i16tATLSmhODZJAdORC02+ntpy4kpsgzQhkgEZ7KxyhJAFLXl2sv/rMXgIJ+h
qymA9VrI8G8sKTUMaC7X1uW5KXghpmXFSCDS7mwlqYBFlT+7eFLdDLeJ+9dHzJQi
ySzQBMy2eHxWaA9c9Dut7WQ2AL90+dnj0Q13mn0796k6KVWjeZCZ0HndROgk0a1a
NQKIcJcIF82NiOQLuU9ACa13Kn+WZ4daut1Vpdf+1SIpg2ZMlSYVIL0G3QQAXsQ7
va80+pvhB/Q8dMqhQbQ3JtfUm5zGshpMyhsiyBGGdFcmiPN4hXOOll/ZrITJMwa+
/IhOx3q7akUEIjVavwvwvz2WcqWkmhiaKhclXQXVIGbIVYRX1EKI6Pj7nUnJeGY5
0Iqz5/AYT5egQYURR/GNNTqcGCbJ5HG3re+U65OokslX3hg9ie4+SwL81vFhn3Ji
q2QAA35EkQQ1X3w9BT0wqrUvepuLk4M1fbggGo2VBSRoWh6oDWIyBhs1Gs7oDvT+
OIdV2TDC7ovkZQPlXSQLsBD8NxRgBI2LebpX636cWPjY02PR40CGSPkDLTKbv58p
MAKwbej6fIitql8XYcc2chkqplqACusnIBWmnFOXA0AQhr5SsFWilErM1g3R8haS
BeYOylv1xMya1BGscr/mUkEhKIPN173RePlCYkgOUpiO1ei9cQND8VEMbv4CyWYR
fkCO4mUvP/eqgeR6O+ARNSHHltP4+/DPccZEWUq//J2aT/aae+giSaP+gBVK/pUK
5dYb/kt1i0kj5UGeiDjoR8C5qCqzhO1u1F373cqKQa7LE+tzjQZL7nZ0GTi1zE9C
h4TD/lPkWXjxdbv5qPePER+l1yUMpNsH0O3ZjAEJd4oL6EHIQKtizVcfjNO7nWsE
mjVUCAfVi5LsRgDGCfwBS9cMLzYzAOAvkFYwKBT9SYaeT+/i5xTaM34dnpknQyxm
0WFEky9l1Jpf0cI4Nnt8br2ynT+RpMrQ/uHnTMhqFSdRLcdvKT8oM4AqXoXYvPc2
NH6sZ7ogPG+pqnwEj1yjKY/FfthtkMPpVtOIkhSTur/pTlonLiWao96CmgyCSrLN
s4zNQ6vTzPldvQ915lPE63UIAMSB7XQG4+BUcjAaojkB1M4zNRLbk9cVq5Je0+En
f4tNyIjwTfq9i3Op0FPontOa89ftcm6O5ymOIj2FMFTxOkDwuQNj7oL+xk4AhDg+
59S8S+fz9xswNkcAp8Fm5yoIchnN9SM57lKtcV+tj9Tr34/AakTe/1+qx7NGmMsY
lRgfPHrJYQeDmAhoPD7lZUGAPa05zSL+q/eQFcUfHAl3v5xTcVWu1JWy7Ew/SCuG
OSGUeqFkpMUa+ltv5pCa9VKvY4j50o0gUvYc6LYhBYOLPzb8159pCjgSm26Nip/i
HS6RK29681V8dvB8TJuX1deDxnN5pss9HKLOdNnrR0mmwfD6L2Pa7XcxiCN6Uzav
MteUY9prjR/62bpXL9CVV30s5E2K33R3jrhKYcsNH7A0HNnEvyCAqG2166MsHHIR
cL2OUJmPKwU5IXJq5KsQfGOOlA5jLN7LMxMEf63wIkzjbSGVS9QjzXBemnZ2gNRF
Xu5WN+UhuYr3+eOmgNDbB8zEIXS2kTDOdFCbxCl4jPtT7u7DKqRfute5ZJGgxxPo
0mdPSyvORyDZyi8I5AYbaeJpU33IUa9/gw1t3ARuzGB97hF+AJxBEDvZAmQjOVP7
LE5Jb6qxxZfGJNDMKJXj+o+J7CtfS4ZWeSLs/D1fog7KD7QumpMzivJLO4O+rBRN
GelB/L3Inw1Fg/7EPPVqIyw0k0EBLWf9puF5E3fGhJrQmKQnPTCDUBY5o+3RAbEx
iz67dTA2epqwHy3uvuyGMH3Tdiqf/rILacpfzTGaVKQ38zBCRN75Yv7he4jTarw9
EvTC1ZDEgZtAFZjWB0YlOwVjp995gwqPmSZRdE+gP1kcZTa1bGk7ofoITBXCiTdi
fS+7u41SljHWjC3Pk35M+mnXi8zJkNkEIv9yZwJctv+goF3CxEMtsEn7/ISjC7Nj
DU/TFB7xGbeYXTJjMRyUZQhtgzBEm4XW1fZhH/adumeWa/oT+joE7iB3Chrk9im+
n9mp++8ZUpf259iVqaPqZ4/hHBj4vYEpC0rNJUZ8gTnuTghnG379yWZTJ6cgp99t
ujD0g3apZ7KtoGBuravdsoAaHTKVP787BJ6LYdebVenpd6eJ/izdv6DvSKc1Wi5X
SyMXU09jKFnEwmSDbLDIi2OLRDxwCUjnw1r9Tf7UMJ41nbAF6yPCx7uSrQfqYs2b
Bt1uj0t7i21m/zGMVKEIOujqvtXoTFBaftEol2lnQKiqUXbkgSxrAGgrpC3i+ABR
RXGGe0OeKnnjkLeuPnRGWVwoiZp0N6yWLJMq2i01s5SEBivmS4DA0STRCoEAo+AE
YoQ3FNhbMfXmF9VigHCtCYiUlgxn0FEiPjUYsd0EzOBBdzf7ehY7CHFVsbeTFeQf
uCSb7vDS1akSwXP9SIrMsTe+MYoobgZ9C4FrqX08znQJzdsRv7B5e90m4PZROAOS
A2QityQUUOU5Xz32pilAMaH+CjYPAoVrrWf1rpD+F3/r+sqYkk4WbaRvhhNdhQnx
roIkcrV2ce93IKAtSzsmjneE5Tx53/sX+NgD9ZkdODdQvdOXWf8TTfUGuhwxz1LJ
ldQ7MJM0j2SPt0XR4TXtQ58rz5yXJHuKFPg2Sp1lXl1iLAL9xPxBbdV2TTRbbDdN
Shvz65q554KoOQHAZ11iYpLiGMHIQ6zOI69hxGBmyjOUh7bn2iP/Oe0hIUkGNjw4
lR0EL9TnfuM0xxpDTMyrquFX71pOhEPpNPdVjWagrhIUSeayR3bqCNO9bzeeZm7U
Cbi6VApOXuGevLq8i3H3BNGi+cLZ30nQOsSOeNtH3dsMHiiohuTw4uBOqntR+XhY
N8oIE/3zin7+afDGrBdaKVPVo4gwLSb4E0IL2tmuY9CtvhWdTXT1Ba9Kbyl2v5Ds
AXOqwYx1ZOEfEfXxOsjb6rvH6XATELg7+xYaug6d5YrrCl4sao2UjJoZ1R1j8iVv
v8oWrKh1P6ra93iTLzelwv6p13IEsaxC2qkavfxw1XZN8Ifn+yDVNnW/Ci5XuD6d
xygSGu1fy2XUYj184k7b+97jROucl6g2JsUC4n1LqYzGehVntMILftZmGvUmctwZ
poxvyopGCIkYy6vMdcVtWG8DIluGkDWrlP/hkcIjFrPBOYTWnbeKqNx4jWi3LIKV
e830qKOLnf9HG/+QeIICfdhs8v2CuRDWtnsr8tCQ1g0ZmSXu/JFP7lPpEZXBMT48
PjjKD0M6NOGvyWCD2e2dZAdLuwWeFgRmzygdhnB340D32sufIqnrVyGDUVuDyeeQ
MtG8pNdgFDJm/O+mqcEIELpaEqv+Lh6d52EUviLyBteYEtk7XZ4GH9MPyWikL8OY
C1iPaXfgdQtkQP7cCHLAQtl/O6iIeZ7ioPyVOZpKC3bXmHdyWEmI2OoWSDRPX1+K
s/3jeqGclUU5ayrA90H93zXHA5AIKKduD2XOurofTOH64uZX36h18i03zFnMwqmY
s8MxIc7kmP6xvvz0bkLnNU8DHKcEInsztlTVnnVQ5wxfivcldvgxhn2Hnn2n2Cmt
Lw/qMaxw5TYKNfZ1rxirjxMNgMSI17DI4UOO6j/KAtIWHGkEC6893nsPLMGR09BH
gpyJYqaohKVM4vazKlQoySTnvd0BfSJGC0luWZ6ie7hdC1pJsN2Iq6zT6D0rtClF
fW0jS9taAXB8VMfmSRHYsMAdzWJzsUiNkpYC1lMhNvskRppFNrg1TQfSsHFpux52
vnADdtB2y4yxswbNL6stbBQDAfMgIK/oawfWQsIknufOTEcAKNCfeYmS2ebWNkmI
ERaSvubgQr3paDMQZW24vo1mMDs0AVE/I0jRcBsB5TEniqIIQzwan3MjRQa5dCSH
CBOzegQA+FK1mfrZvuAO+xQ0UWCiYFh2bT2/BhaXN6za8t1dKOBSyUegGxvMgfGO
8iT1lBp/ckOys/Cq9e98irNPL7ZQQSBVvvfseCpEWVcuZDgXdIQXG8hXtgiQBNmH
sqC0dJoHEL83LNdz/bUltvwYx4dWLn3rp9Ac7/By4U7B0W/3QNvGMAKhqKWKG8zm
OnBrJiDwpD58HoEPhhjDO/35R1onze1cZVPZ1SX78t56yYOlUtwiMRSxl0jlJgWu
63xpl69SXuAn58Km9+MulB5l3Fb00rCPgTdvoTroH+fNPk8U4g9V9KWK5tJ/Edcj
Rk2jHWh/T1EZclxC3MOd3Qx8dx93oOwhSEGEg19DFUM8QXDua3bvw9CFA2rS1Jtd
cUhg0yCIWEwY4aYahMgf5IXK/eVdjstkK/ahEh0QrlhcgdQdJUKXDLmnBBhgEj4Y
TGoOmrn5B8RtiKtob6SS7oZLTOiuT4i67vz8jf2OvhyUoa7bqAlAMQJ4MqhJuqx4
bsifW9WnctPlYo6GPo1anyyTA4O6qGUQyJ2ztXIIU6VlAThLnBL5ttct8HoS3ccC
zYchhsZ+WkPPXzYjxuECFgDGfofKS4PFmZmUXdShG0LXsIpWISfXhf3helrckNIQ
z8SMCpf7RlvtF7dvj/E/pCY1bTPIqjxTrjIYAJjyh7Mu48Cd0tqSVw0/sLDtwh81
SetkILHHKdKG7skPS2GbUQEtVHXkJQtr9wlXJCe/fXAJaB6PW3iXwMY2Riolayrn
sop5J9j4nQHIbQnlRkCjr+fqaa4Nh7wRKTtdu1xcKuf99W2YLobHhPggIPhAkol4
DZiZ6hs1cWBUYHAQ0ahPDy99NGmu3lBMo6oMB5gArEt6f60te7OCLxr/9DKbBrUO
3nIMgPA/Pl2E8slChV13C3LK0y+gTt5ZkI1JsaIubmL3Rn5qnihltEZg6SPNsMd1
pDnJvnV4mi3DYsL1MCfsnGfhuT95J2jCFJT/1kvdWtdDM4dvzom1zPxuG1lfy5Pc
0l8rcix751m/OQpLcnQN/w8V2JT16f6Zzz8w/qDNf60D1a7cS9SQ/XoEQrfVc+JV
uITbTe3K3J+8khhPyPj1zymccsYK9xE6ELmMYmbSMGhc61fenKepTLFghrNcKq9I
SmCrY1E0HAJojRaxPYm61c1QMHPhNbBtOcsDlYt/Kx0p1K+xEALcclfwJ43g42f+
vdkY0Uiv4FGg8nFskSbTM3GHELxaKTV6Im2xnCO//Gf6zSHufK/muA77Q69yXImq
tSfSVoCTnbOh7KYmFJ7ld0ahIc2rgG/Ey3V7BIrmtxbsWT8Y0lN3aDgxFmIs7Moe
Eurqu6471h+75W9/lRl/tTUu369wJHV2KDIHjYgnRZkNr++PQMjgfwRU/iq/pTE7
e5eeACa94QDGxpX72q3T4a8dfQ2AY0E1ycIW4ga93RtghnkwjPjZcAuw1c/BYn5U
2+BhVWG1lGz2B364YnWiBG0/NwPHRmstSkJgA51fR9lGabPgUTR+gJCg3/VrNN9t
f6gCXXBg5Kv8E8TAVODut54Cusbt296YF/W0rb4PKcaI/CEDWh4tDO9cjcAsIbLo
NBH//ZuiJaCVgPjXoqBPjBKRaAEabdFwNkcbKvdVKQ8l2M4xvCQ9q8PRvjigANS3
gG+2s1JqDWYOySPnf9KhBzIVMjCiZzOf5AIih14U/+i8YSU20yI47uCr9cHWmwgT
ifOyQG+aw31pwx9aVkEd2zmpr6P3y40JzGUp7qbIlLhBWz+lMl7pfxu5uPN3fQDM
/JeXSLaa00jUMhcqUIslAX3hCfPxqs2a+DUUOJdceq9htbyrQ8lh//YZtYdBkxkt
mzWWVHykEnBSebNCs/BnTHagYiDHruArTZ7RBgSOg0j0AJhOdCwxrJHH0UDBy7WI
8HZ+w4cUzuWPmbXCcn30UJjbRJ9wkOq8l7+jqHhiPcW9Mee9uwOyfELyKdt/PPF3
fRJQUI7w3N9LYzr1SDLD0YCeOkA1ZhFrMJ0/11YrEWpNkWNAMIFXljvpzS+kwbru
2iA90aK9SnHqoN06trE2NregiHj3z6kz+O1S0c1cNAQdYTo6ouigS6emsET6jNjV
7JeOOjqjTEqpOfZlpYdUiOkmEnuzVS3OweTn7Utdg7OvubyxJaaLoJyf05E4ZQRh
ly5AfNLWZkmYx52lNbixbtHLrvak5SG/KNQ5fYDtE5h42yi0MR05u00mTnlTKnWt
SM0qz5N7Gfglmd4iyhA/FaGUQSEvcpvpipd9VuNJ5BtU1zP10h9mw10T5Kj5d1b0
+2a3KPM3RT8EMFYkTlFaThX33C1eU444P/FUDnoVtqCZ2iPieVxRKU5qbODv+sbu
Cv3h2iCnX2w76L0J+YeHbpXAP5bePrIb08MIX/lxyQolHVi0JurO8sYrDQOiiQge
tpL9klzUveRYBZzBrcaU3mj+WxfTYLCKhrnsk6iOhQzY0ZMe75GUESfAY+DNFY4h
jAiYwcbiCjR5RfetOdwEvJ0PNVbsbCqeUqj9iuyV61a50/+gPbw97tai2RV0RvUN
EqNsz351pEIuYVYkMCG3pRrTVr+AsUZ9T3bSNGAjyf/cW4I4gDdolYhTuh64jLWY
fDcMIU6SCTqHypwxMYtD5KaeCXzpHIl9ukTwbP48PfjnlalIHsucuKzbD/TI6Wj9
cx7B9+gax1sQ4IpPQJtvBVAnpMsID7rbRRc+4IYTyPyRA4GBSz3w5WkKZljB4Nbz
KQQq0eEffT/Y83uSFwrlTkkTNt16/r/h4MuSsnWkm9nzx7GIu0pR2DB7DXmcmQZw
wddDFdHOir3dSNoOWseWjyAHfyU/z9W7yHRp/iD0SFp6Cnq1BMjGJ+n9v2rIO5nX
VFC+pot6Xg7Rpa8jEcrxYCskx6WK3f8+pRyrx63sM4wc5TLz52BhkcjR58KNZmGD
Pn2UwBB9Ga1rOqI5g7MFGbxsVXipOxJxMqDzV1GXHRLdFcEa1162ZY7ejEz0mb1l
tziLfIz1/uuiCXKuyBkY0AhebU4sCn6cotp51423QSDFIsTJRkplG1ksRO1lp936
GgOv8/Q/3NQwmITu+SBCoS7c5eu2yTwzEP3cSHbveLYeWMIAVnmIjWVLsbqm3IO9
rSz/Xf1rpg7Fszls5FwSq0pc3SFbKeUk23UXnlY/XdKHTcwaI7NZmheNuvn/GBh0
t8S1pR59IIuiOhevEOLMf7yIjYvP0yk3+k0/DY48oNVDZCmfpmz1OM+zbyMRLPxu
I1HMgyvg4f84qdfFNEJMetgc3UI2BhcBRXgTx/Nc75Q9YC+E8h9ePi1Pm4bL23xY
XqD78dN+bwPLtprMBVh12DHawl/EUGWKY44S/mJL7MuVmQ9cVdhZ3ezAW94PKIX4
upDw+qZTLaKBvdyHVDeh87nhve38NoK8zZJyDlTFjjYE8CYOo0IOXmr1n2KtKmkV
MrWaG0btxw7zM9JgWDTZh4N8tNDHdW1qJrSG1eGJntAW1ivu3JS2z+/oAQOvUoe0
uPxx0YFmYGPgmA1XWd68l5s79DDJKQ7F2miq6lFrk7SyKS08E+jkgQ7acibQ/+Vn
Flwg47jO1r4MAsBq7GShlIsmslE8VazEUVH//jIULz3Hkeq2EFVdT6EouZvGTNZ7
Fc2yna/ouEhdc/eaZ70n/WsctrbKw0bDThdR+0p7UT2/ssznOIrGp3VUbryzPWll
GOueCR3Ei0lNBtb7guCPrWCzDfq+jwWM9t9ayDyR6c6eJU568t0ctTxopALuoml5
01J3Wbr8cncS2IC4HGt3/mQtSfTS/v2onwzrs68inLzirWwOGHwmzO38eYPMCs+1
Gy8JwbCueFgtL1558wX4ijRMuQJRAypr+SeOjB5JgYdxR6mZLJFZplw5EOHRCcHY
iMK7pBvKOxvq8CqPgKbOmRLcMvlGUU7F93cx1WmD3x4U09u1QCyx0B4+0g/rNTsv
lD0YY1/zT5We+xg/k8GTXT+QeKFmJNwsPhLsBERee1IC9DQZXksOh4xTtpAmQKpQ
1VGjMMqpusu4RGUeaM4AOm2U9IggDWNAERO47VEUULcVdn7H423Akk3FdwHgzIq3
w5oRtcUf+GWeyCatckXP/JIm0OTKXeD+dqR/JYgy1gEggDn1OENGNoG7G1ROJvPx
UZQE/NcZ4I3fXDftwBjKc2jHKdwY/CmWe1sP5hmOfRDT3RtadcG7NhR6eJ4PnJ61
wHHBSpXrOoxFZeTqcH0HaM/bk+YaMDdsyQmwjY30VxgCjEs5kPcwcz2b/a4DLi4A
FCz+w4iIPvlWaFtwGckvFQjM0N46PqM1cmccFlZojN7g/plmxlWYXBTzwbh2LNGv
figtbxgaC/VPzelct8nm/fRj45kwbfuaVd9gmIt4NHNeH5AQyfYwHDAlVrE+eDsw
3LX3mmMFQwEcQxdtOejLqOIRPA0Qu4fllowtxhwVu/JjbodpA4uaD83WbDbd881Z
i7k5axgU/MZeFiCW7agB4b2XDov2XX2pWr02/rxWkXaxy+WCMBxHrehC9L55h/0N
4ipoGr3eEJJZOcjEjE46CxCJFV8B6UNNNpwhKEw/EkFt8bDfsQKozX5vefTE7voQ
GTWK982lbj27K8nUsOjrnHfbAX9zj8Ozj1jtcAiWwy9wy3BgAKpkBPn4rneK0wZD
MOkhDM5EGTVN7AUYqUv3BTDH8XvQCvpqMXND0qj05mR/fSWdoQJ2t63IU/Y5A/xG
mEuGdtj18/Y7Zqpt3CP9JNnBCpji/lZYfse3dHoPHYrLY4NvD7zC84xSkYaP1j7V
TIWfKS/JJfwjKhSdg+VKDLtXZgZl6GDUk9k3ye7ms/e8oGc/S5gPV/tHPq7gfQ3d
N+mzDLW5aCEkReQpbUhJ42z4pibPy09Uep6lCxeDGd556PeEF6AUaToHKb3GcCTD
YnhNV8OdacsDq2Q0IVeBkFOlq0pOKUzJc6xM4NAnzceqFpjhLdoEP2UgClVgl3xO
YpUQI8UhDZmZIgktbLSKDfQoFnwTvqQ7yUdaxEcb17AWvBSLElNwrmED/y61+aU5
1G7Qd7hBMnsOHdgyRkfUJ44izPK7fM+uztc7G6ENQwJVeKIeiqvATb8BDMsBhov7
FBhAKtb1aMRB0t61MmrQm2wNIc8tF9UPZnzSc1mCGsRfTL+GfXBqz5ihFjSBrwHr
Q6TpFEf2HEx0mDal9urH0AKlz4onNBQIdiaI26UYrb0K0agSLyiwukIx27wqx3CW
lltNtGw7WMe8t2u0OxeP60PCHOUH1KBYjAhPjQ0y9RiV15WX5R9m6L+4Ms1IQef9
0X8OWHAtOPWJCS8mrXaJeKCpROZCX2DmKSCe2nNx3oARxh3tlYlK8ChI4uDM0a5v
oySRm1UwJoLOCIVSu9TsGaiWgw0WnC5zKYv2k0cD9D8UalCW5ujRyhFvKADGt/Nr
ugGejyd3mM0lZno2aFgDkAtXt7vKtmnJeXDMjvPxdZ70+3kUuDkA32u/ZPO6JAts
rjFpz//EGGc/kd5nL2q4p12CDHzTZ8GR9r5wkWyv9IK4kNpTEwNvCbgsQgcrggUp
Xgl0ljVr7U/WFutLedxrsNY7vrD271L8Ul+g7aNW6qP8yimj2jPqPuYotvvlKmE9
q96gvb4Aq19iK67WTpsutSwoZE+jEaB59QsYQsx3LLI8C1AOXxLWZlWJ5unKtEId
KbcgnnxD2cPvcwBfKUQyBWCVGPhYCDgNrA8r6juedoXOLWDyObflBrqwP6d4s7aU
rl8IZwD/eVLELvrrYJMaGaHXCWrJVxN9fseVmYm3Ze5+nrKWjp5TD4bDmyywT3HT
xKCijmrbSzRg9LoTYY8ewz79rRCUv5k9qBjLzxxCUSm38JCNixz1bNO6GP6XX3Vl
Lr8wlvZgd6XKc+0FCp6/U2poEcxAn5I+VKw1KwEL3G3yWhd4oH+lHli1dX7MDFtH
eJDFRNNtUgC3D7ohLWBtR/+MC6KXbRZ28hS2HS+sTc3WJZ6nshzzgD8sC9ewqf9z
wL2pj28TOiqqIoP0lS/u7QO/UuxMibEly7T2J5uE/PW3aW+oyzHsCSDllWc98mix
2UarVln5a7aLnFkWpMZvf602n6V9AHlVB773n4bpVN20gSGzgwmpJ6n6F9zQ1IE0
5cEbTcGVG6wGhSe0bzF6fL74ubU9wg3+dw90yUnW47UTfOiH/vP7ALDxUA/HQfUU
29dH0yGEbTVQJrQmHXKCpfvn8UI8o9fC3qhOdvQeG0hx6aQ+q3HLUYZbWXYs+tbt
Cwkjc0bHw95JgVOrpydYsP4MMwXrm/DZukZ/F145sbPivBnGAzMHMXor0PhCwhlR
BLNY3YPbh4o6FmkdT+gBaxah7LJSSdF1gUjnhS6imRtCPw1Ctee6fIKO7g7GyVHB
/E4VzpxuyusM01L1C/a1wjJhTApKCjcSLIYtxGFD9za0JlC5EdFLobEFG1WYsVTQ
BBpuNpYWC9athLV3y20UMIW7JRxYJz1L3rVEGQhPJ+CFjIKZyRKnXbfdJFGhCMUL
U4Vn4ABI4M4NXiw4EWtpKcjFI449F4Rq7x/LRkKVqiYU4d1bIb2QFMvZxZ5hRAXl
6lwW7Re7tXic0iKuKkf+PFYT+nBOTI0DD2NqdNXx+BC4OfpheCYFap32T+2vMI/H
7EHOBpc/wrt4JjbW1lXxC1ciZTQM9kCgasK0Fjq65RtOhBM6Y+Fi4vUIhiPKp8Aq
G+BAeabxib2YoRXeuSqwaTYbI+QFxqZR5xxH3ZXYvNz0S4MESwXVOjYwV4KiBqDj
VV3oAb6JS0IQ+lhZm1yRCxu6c0ruDMp9LhX8pIIpzhXbL41jGnBZwQ7mpMjlFzsv
g5wdMntPTlunCa3pe3krsfAnCg8ZQBz6uf+B/jLcCyAa6BzJKCO5NbgSWWbVQtLc
Vkp8TefyJm3f9niWSxzEMSZKKhJQv/ggY7Gvg9I0uVHhlVVSn77yUGZzOWR8Mrb2
H0joCBVcC6Rkf77lKBvTwzi9cgIc3ZVt07AVQ3qJv22HLfw1sRtflt/v93S1M/CI
+XfTG2bHYZj32FNjyc4Kxn52fDb38dTPNrGnWQo+tildYqsIC4uE947gN7IxqYRS
nhspiOlMK/K+SqcrVJneTg2b+y8DbwaexaJSPwfEnLGvLwCux2Bth7YXiBgo02/5
2nhVd6KUCAVVUZFHn8xpr5QrzCK+Z21jbgeYJTPH/GhXvSm0iPx6VQ2zRE3d6171
s8tPU/vSdVi1LDc01gP4jt4rHFNAwqQRZYQHN0PpxEBBdbhe2jgALrPVc+Z+9c6r
zakg3csnmYO8/KAaw+401ZfY/cYlIbyTylKi1ZBmSeIKE/JAT7syNfTrgd98Lese
lZylpST1Avkohp68m/eQA6S+wyak02dQVnU4+hHnVG1i0FnOJi09PbbW2EDkY/2I
NY7TgXw6cY1OmghZFpPASPcSxosHGp0QLPI4+09n0KDpeUn+WlFlEYSCWt0D3Q0T
ELtwYYztJedWvzxeJjKwxlxNYr9Aex4MEYY5v6OWMzfxOIfgQVzqURWqQbT6N/HV
1+jUR+bmpJNI3aeD/Eld9cJPyoLSo6WvSwnfuzgV6FLIQsw2cUwA7X+dFXfB0YSq
dH14YajD0iwdXuVBeNbjZwk94tetwWB5g3cITWWrvbgH7zbz6wSAqtVHG0fqyUS8
UeM8SUX9ULShN3DzW4o0GiQwU800+a0X0orEgC1/H0gEyAy7M1bT/vGiHf4qqsAH
r9ImoGP6Z6R30twAWjNwjmt7lOQqw+tZ6wU0mWBsCcWJjS1PjzHHdVKfMOJV1gw6
DNRLdIQwXJaRlENDF9RJbXlrvsBvWQJuvk4kEQOiqGxREsccwqYSsU8HMz7fihYM
w+p07oVBLKgDsyqEuVzKVjLXBdMHOuTBAZrqSxizssrKXlSWlbkoad+dTStyoqYf
GjcBIJC8YsDolEgpeVQyJfwDiKXsBf8GZgt2QrfoBU6P9cADT9Sg+3RprbK2LMxw
qxIkAjL5Wf7glwxA3H80eY+8pkh5SQY7DqeSYn9z9E40OaaVReW7LQbammqLicDW
dQJlGGAivqRE9np6GOeD9x0rwmsIBjpudxM7UutQLNtRhbI3i5b5yIZkJtTiI6oc
dIXyd+F+Fp5UhJfUQ+vFsr4YjyE+CzE9TqcIXefh1CuLcqYLiQ8HjAH5InxJ9SdZ
UeV7AEBSZeofQeq5TkCE/ftuylvy4UC7nGMz7EEnbllHVy3q4aSzi0YYkHvTTMAy
D+6iBIMY2IDCwSV79gfRcIdD0SxpHNcnKO/wv/Y4+9+0FiCo15Oz2BrJK6vuG4U8
4C11fdzAbdDVxLa8G+9K0G60JyiSctOyg69FvnU3OOa2dUqA2CpWLmWyC7o1wor/
a8A3/C4ZOITl/BSJxbkFyNJNIVu26GxoQhdmNxKk2ZTL1zRDkIxUof+u9xZLhPXh
aImra8otPdS/fcFK05EBxmqvRjoQFHOOv/okICgFzIOXJMqKSoUnJaR+d/20EEE6
K+WAXaQCnsWy0Fc9Lf2vn2rRagKp33ILAAFRy1ekNrRx1ueoEhaEcC+A8OtJn8Bv
+y0dFsRLMiW2NJiBUP19zyAf9AuVZdee2safVD8Wa2bT4sY6+/+vfyq5gfm4EYem
7AaAL1qPnHvlQkn3SybONG98xW6RHSAPvqRdbTSPn7RFKi0BomsYEKa4HAw33v64
I5g8EtBBcdY3atO5Bx39CuzNauVuSSuPY8iy8HUKhDUJjf3oZ3qwFXsgKUd063gG
wMMb6s70CGFzQasU1Nn77oTo9peL9l/WR6DMvZNkGZKL26Pw39+M88ynA0fWCHnK
2VIEJrJxtpeiu1Zes8n91zAvDUOkYZ/G4eA+Z0Mis7v6TZD+NVNgBrfWs8mgRuRB
9uQjmV4oWafX6a7NG+J4u2xPwrnqI/2INVgK9FzjLWlP5LZjO7aoJ4icP8Ofczbo
T5fKUgVPcOpzxRRzeiCKbFoAsFnMsBvI70nj0qd+6Uu47f424DMqZK8pTBOMkXqu
haaspHXMdHRk2ieA/x5UfFUHoREu1HiIb0RYIpp+W7g6jk6zgATvKM2oEKMhzQad
sgb9VBq7Vk8q455SFJTVdGz6hplQwvz87ljl2l7yfxWBDAaaARsNpweJkC2TqoVA
ol74u0LiQpPpiXuRtiZrSP5OW8EPxcsyiX80g+l3TBCXsYtrFYYxfRHvQOh7nM6B
etxP2iALCLpV5m2XQOgHZHCesXt9596R07jDuMtSZVAWemjIMWDgcn7LVEHhsz4G
fM0EHqvFHdenAN9bvrf6ITGeymZ+X69DCK8effxaF/6h0SsRnKyqjqypXc4Uf9Sh
P4L6KZiLC/3P+hpons8Ba5OAZBes0nKSyfKPR/48QnbPaYPljOdFP0qcj2QFIGYm
rDpBkEwbDBACEYYR8YfRIzkq9LFLjLZ/yzpl09aOkGKAApDbgktdTbPooIrW1nHL
qR//j9Q1ddm2wMi3sTxb7XpslOTR+xmYnCx3pKo7Xr0sqP+n3ri+qAWp4UCjfjUn
g6bVoC5OmK2M7UQy6zjCjx7TXnRc9ncWZcCQWzzF4LooGmALoJ50xyCcN9d/XroC
p1E+5NqNeoGXCMy9exyjb1WTgsJzkGEJgyJIEerCbJkqI8OVbEyHTYgqR0umMKq1
hDFDKVAxMduuELxUBarEhFNvcL2WTQ/uRWxa9zPloMiMvdRBDcKptrID1RhW8gbL
XA8NXi5oF5xf46RPYRz1f8rO+r9g+kvraRsh8WbSCT/XGhLlMxrSscky17aGercD
jjSz5bvmk3ntsnt+0NVuGrLYH4+1tIBe+RNCdK0rntU1FX6cOtzbq31tH74Aa/l0
IkrlmBaGgx9FUyrjfuJC+PHm9kDEsGswGQGg6iQSnoFwFgLLppDP/X7fWaYwDurw
T36yDuYQA1uFQa7GSif7YUZarUJmb1EAmoeYwKKAlC5d4xtukxWkZjE7JWmw77HC
RNphCeoOoZ1vmUfJGt/ysQuT7UoHutxCN4IJHa08JW+2yjPYd7T6X709GMkbldDj
X2ifVL8I14YM/xO03yA3vJ7tMKhfP4pjzb4bp3p4EBv2EFWJKvfkj8Q4RNtretnS
Ky9CTk7wrUY+bZQzhPGocd+fGrjoDuj8XX8lh57DaBWiDi0Ej1GjkKbObm8YREUD
T5AdOSS6mJWCc9YS0cFjm1tNLuV8aVGKpzOniiSN1sQji1jOrsqIF+ZzKu+6+6CU
T07lGzMMIs+01m1GKQLt2LGzSNTYovEeCGhEfL3mZj4XDHDcE0PraJ/0cjbXs8h0
IS4WScN3nlIwi0sCJs8RJNC6DB9d3DGYC6UUR8On+xFFsUrCb4kggtEJoFMqhkzE
/A4xaEZyw/ffiLjIf4NkC4J9fl8LIvdDRt0MvnhpDJfpY/e+AWJNnGYRX66lfWfO
Q9OeKkQ1P4oWInvTnk48qZQtPM1/h9cQ1Qec+zIA5g8sAwUxDb+RnKMwzG3i4CTO
jVSD3LFsKtKfFe1h2lVNFvKW8RsjVLORws7dU7RCyHGVldS4EXQla+iiymAZD4+F
FgKcQ2QoxjAk4trltOC1SaVT6RQ7Adxj9/O/pTEmLEcWSDsfwt8YyJxv9w+VDkqA
HrMbQqKw96P4Kym88C0npFHfwIvp/bDcr+f8ysXTwvlCnTXRinU3tHhQpeLQocC/
Z2AusqMwXiDEdmUgXoo3HE6PrYmzwZeMNg48xJ3+SkxvP0owDmyIguoSfSMRa8Rv
j6DRkGQFgz60ysQtASuduOFoVI0iWBMHNsh46dyrEYxM5zcGHyI2LcLT2lOQsz8+
v/2x++8YY1022C/58DKpqmZNSumwnzu0SJFX2gFKpQEq5m9857ufbvuE9Ploafbe
cOKiYBYEu3AxhDAiUY/4EAndhrKsJy9eKOH53nh7l7Veekb34iO8aL1AnpR51zyj
t4W6RbXArPLxZhW/ILkwunjsEhRJChUqXviv52v93ppM4jgKQC8vxF2k4wZYdpAk
s+nswAIBSF7FlUGyiLsKIN/Lr26mys5lgR1hN1A4b1pnslshj5mMgUWwuvaOl5N0
+qwYkQghwIOqi8QpPHS+0Sq0gFC2n4BHEv7CJEIog3pq/ky1V9VULbZ+o8c7GXVn
A+S3y13ar4UUTlaCu3jC25PRG++JGOxBiSPwLejHcPHbHtYNBAfyQ8ETcQNp/cS/
nCELmZ3LgL0Ozrhmj6Ai2HvIhSUbHM+ajiSJxYEhL2Dw1mtyQQZZ6agac+wS3gu2
FBOgt5mctFg+MZ1A1WNKIcbBThQv55TMxPBgVMPUolUeT5H2Dytg4ml7P5IL/N1y
FtpGdaXvKFct49olW3kXEH2BJleNhSJKk8IO24E3izbNyG5BUm9m+BZNcTbjH7LJ
cBG36zF1DjddNnIz6KYwm/aU3plKf0p7cJeUdJMUPysuNmjkVaIJ8swb8pkVRWME
2QEQ7Y16dZKw9lBy1IgI12Z9Qf+YOLayMzZXa2NxqwDtEya7Mqyeb0GSUq5/PLQC
LCvEK40gzsrZonohPjP+8t/Y0++uJT7WodeZyZewfugrNbqC+YF6Il+Ich1ZOBuc
3FrrsSXrK67nLXKsvYodNj/3EflewUsHLfbOzB9RIn6dDbPdYzTufdatqtGgIqUW
Vem2QpYVh3kFJQRRfRpAcAI9jHrcnMXMKDAwffRthFidvqO7H8qsSJUOLOA55y6D
2KjroK1G5nno4DElgugiXo0Wk/837RUPVkfbRF+JtJQHdqnm6SHxojz75y1URkvB
KuSSDLjnqWiZYZHJmVSk1nX6ucR5rO3X3QfT4+dMe5BtO61qjhtW9tDoRDJ4E8c9
COJcRHi28Shmiskqb1mTwGdpe5yI1Mkgt6VcgHW2fS9ywUOCQAEgo61EIuw/AF2U
mX2j6NVLa5rCxrxV2NaDIveI3sFYUuEM4qN2x64ime/5GCPiPwzk+CKFDjkkyez2
k6HnXOGWtHOWP+haVopOw/bTxjsfAagRPt5y5eJvJPBGg5eWlxjhKT3LXBi/GJ5l
Eqy2KFTFvNQJ6lDkJxCyE869roL+THmepGSja5gJHBzRKlzwz8O9Pi+R/ATR9LPz
nhVPJl9hsofTXZeLHaShrDishQlmWMKMamMBy9f9NdlEW3/N4FbiicTWwiu2A0KJ
TxQUU8QB4km/kujud2M7idghxRRkfMhdMes3QPZsxXs2p1Ju6Y0hBZlO9SBy0h5U
0DVvFAvE2nKdKxePcONMKrmhzMOvSA3MBAdt3DydvY0DlrYFaEZeOA1qtcnK47C+
qpS7ic1UGpfrIRowztwsN7yOheP53qfzRKXbKnYr2G6b+GGv8GFVI8m0+tr+HRY1
inlZsq+hQGTbFQ5E/W2AVi3ZdUmyDyhsM2HGN3DqV2XELNLOwtvyKW4jJ/F08n78
/47Figf9pXz/Jy5rR0g1hGPslgkYrC/O0+pnMgb69GIOgsyd4J8Zwvbi3qtH8trx
h9HvBkfBNn919HPHecop4hf6PKAJNKpt2tP5150kWCL5cFgJtKG1wZ2m2aQr8o+Z
s/T1+nudEita+Q69cbjvvXsR8xpMisERp0IRc6JrHKK6LadF5QG1oQuwIVkb6AxH
j8+2xKwhAgYDbFjolKC4ZwdqBqwmyvthwgDu4SiMrNJGfou7EOgyERWAAuGkRzi3
WSB6T3HsB37oOnqwmcN/gTY6eAoc3l3Eylcb77Z5Rdey7yLu1/qhaQ3ZPXfQiYbu
pE6Jht0I7p7uAlB9vQPINDxAoPtrDrrbstipq2CxM2zNNSj7QLIA/BqMZ0aD1ckD
bKd/B/n7nuAaPt0Gsc0gWTgwXiMhAq15scbi29H9pe+W4dhwNpuof3f6F0F1Zv4i
mvQGkpG9oUCemmLshSsYlMnBsKSFBEQv3AI2Z0ngcM66vppI0BF5tFnC89j27UX8
+dYVlhP3dgpXD9lVSgltFpTZDEqzfFn7f3xNT3X4Csfeg8O29mOpoqH8MokZpcab
UVDtvahcRA4OTHL6Pi+ujp5Xpr4UkuvNsw5rspIwi8/zvd412zCGHekNPmUuIV9J
59Ur5cauzL+nnjIptlF81GvEGbthbdFcBRzi+c5i4ouLnhd6q+7eyIBDfvNA2Dnx
yaxcohJfWwDRuchqw589CVbOTRqs84dbaD0s1jleoWuf6NPCFc1XaiD5cwoh2pL9
cKrhd5FtxUyIkN6O3fcWXVzWE71/a3iBTWNT6Bm52NOKPhLauEce0xFlUpFelp0r
X1xzactmprTq51leuXTQAiPS0PqaiOUp8afa78nJVX8hMNy9LKRZQ5P2bF1x6bII
eVHt295MqhXWk76XPz/rfDIDHKnJsEvZ1vOJ5H/xwoBk5ALFU/9IiPyY0Gm8Iv6c
+PLtYpGRwKmodSVpZr/UTjLknrPZG5PPNmTOJfHIYscXmn8FMeT3c8CSXe8BkPld
1m2RG/Jx1kNlrkCCyN8FPwnIJ71f2pEjcujWt9oTfPNexvaxNKpXLcOy6kXhsJfF
lFVspzRBc1wP4FS5lq8gQYnDdOqxwC63QNIFyA/E09C4M1Emj7YLPi2nVQliGoMl
26s3XMOS1LOi7kF0h2X2eILnHHta2kkXmtggHAT/3AxYLiDUOqmMy2dIJwUavxuI
0ZK0P9LlIbr5/RzZdUqLIu+PXHq1a0bue1UESqfsSEKe6fVOm6HwZd68d7sqqsna
qxgct77zBP0UBl2LjXJE7dOIoyR+FTLo5fibFA+vfhfTwx4+dw89z6GK3VV9RB8z
JwcIS2St7teQFgbhPJzUgCPu/d1EAT794FnWJDub2/5koj4cl+5WM89CAtDcPpFI
jTa9pBe63K6AGsiyTxyqOktdbF7cYiASy3lkVDM0OCZdgD8MT/Xil+xm1lr/LcXz
uv90Wargpk3RCVPjScCLN6hXkd7ToJLhG64klaQM0NJ/4LRqcKfEw+L1hGhylKcQ
rl8Lf4ByYizFZ9pat5zvYNM5KjqeIFc2sJN77bG13H36CcdCcpYohepRjBoKgrbr
KdVhdY7XGnmYHfZ4i3cRwz46zebuZJBUkguJfBnSUBUe5rky0UJxDifrdsWkVhi0
SRKlBRTkxi46zFm3JZd2+lwrrfPgyteVwKe5IehnA0FOTZPQWO56t+iiBwYGf4EQ
LsoYFYlMfx0rvhv3QLHUs0AqWmZM/QrbyG1vLFrgSZMJKuLDN0SRXMar/0GWk47N
GRsEr5DWoaFZo6DiPxpi2tqfUvJr/At4F8eb50BVV2eWzIJi25/jNFRJ0GYrTaEn
AJWXTN+E50Qiux/EFWZ/GcGv3DLIzrDQcPVPhCN8ECYhGKMV/dEkgBzdicqnE4N0
sF6glfAYt2aErVN/agBzJXp9Ti2YY/bDwb+9hnT3/E68WUnmORMiR1pT5nppkXB2
vgYJ1zXFvgMqt36ywayXOK/3nKcHC1WSWzTMkdK8697YJtjZhPaDfMmJ1irfdMeV
QlEhRV4XYwPFJ96LZ8FUrrRzEuJI1uyj+9ai7NjXIVhvVSMEgplY+Rmi3Au1HmdA
anguUmzKHqc3QsrAQad0Cv9Tn1+Cc7ToXcnnuk+xemiw7KFYzO9yVTsuve5ZT1w4
sDiUSFHKxIZbPwruVHU2HBtgKc27HYfU8lcoSGI4KfGnYVRk4hQYrdBIC7irNKme
fjOmKsD5N8/jNMq379ZGKdJDG+h6svhnsRk3fFAqmxKCfN2EStDRrf4hy8cML/o7
LUQSW9sUpNGe3hRqn93Q/olXIuoG1XVyUCJc3O4o/2HhdrQP2iXKJiY/XOoPYki6
YrqrqMzjx58PlhWG6FXGbmkwu+gWVs9rz0p8NKSGGtb09ZAYhqfMVqFSFe3/KLZa
jz+FWECdKbao+Bhc5aBlUeVCqxLWl/30KYv6dLaA8lhiRBrUmtG7LXsKNiQ4HmhW
bzOstjKSZfUFuaX8jqImI/EjII68g2q5+uuisUVkOR/aMIvHhmTqLFCpdkSBWgHa
Yg+TqJ1l6lQAEwDPP16fZwQAEU1eRBIMPHhIfbC+R5HA3kuk3N6SbwnBAA+IYafS
/jUymLvKkEWafPBTZO1Tsa2Lun6ATYwYtzx7TCdna4lJq2XqDfOh8zo10PO+r44X
1ydDFSSB7GFfAOGaNLEaao96KNkF2s/awJLMFi9A8e5HuM/Q6neUfxjSnec5JHqL
RmUM0ptcGsVpP5nvSXNXwqbl0ayJkCCqEGqPz+moeHViUjpOog/gQkkWzhpW4Y9T
W0KqEwrsIvxLxzQ7UtOEK6lJ2Wu79rAiSraQXejYbjkmT0Kf7O7ndW4Ps3mM/LFv
JFnE9sRn3sQz6ZXZyfTdmBPpIaMRYf1WATuTgZ1MNSyWXfz0sMoYXZPNuwQIIjXH
NzYcQxqD7UUjcwaDZg1L1LIccFCtbdjS7O4q7VgQwKHbZCq9rfO1kfCr+ZQxy8J6
OqjydLfh3Uq/+zNQbQYbBTVPg3sTCg2yonGvYmXk2BrI0YVsWW5bVD7S+GweFXb/
P7mV8m+21ws+v/nZXF4Y4uiKfQgAQSuTnQ0LhRJBJ4vtD0FH1b9bYbYDJaOAUn4X
WTeVNNrz3pNe+Pvh2V4E7LFNWGttoJqsjQMIrbGJwfA8Zswg32nESU2jSARM1Him
HvGR5OPQ/PByXLWd0oLKZbHFnfp587Dr5PUEMI4d/SK7kRl2Nu+pTv9iIsOD0tf9
GnrlsZdhvelczMCvpwxGKfEhWqo/ffEMJqV7+Al0BfY/KeP3E294VaP9r/Ezubb4
g6QSiwRSjiI6xwNKlPMNIcQzQqN+7TkMZLXrZOIGoakk4xkheUdZhb/yoMqGlDGJ
neeDPOYm5HB5nlWnsgatGcpbaB7WW3QUwW+CLZC7zdGkeE3g5wjtuFloC+TFfRtD
7kxYL+ApEzzrEBkOUgcBGI7oh5kvdCL7xWvKrKu1R0xEdaRFCCjk+sGcNRX524ip
sCw0FFl5OIBS+jKTtvm/xRYIrl5bI0c7WR/6mH3sKmZ2ZFCrHFTijGU9A+6N7Mmz
Fu1LlruJP5j5TPq2v2tBLDKaFteCHlwd+6g7P2+2HiFs92yWUKCKAoagsELLxrxB
gdE9c4O/wMn8XWUX0nFT0TNBnmLKIXmR68GOLk0ZHfGxJEPzO/7J8GctWXdi4qDm
tRDdmiZqG67jkVLvaX0UloBcOMnmHKepj46Y9Hix3YTx8DHayucXKWa8a+SlTWBB
pHzDACJErjzDCPNDdomDgJjZYCkxYwE4fF2fOy9QdxmuyGZuSD1G1jWg+1ZMWl8F
5yo3h9Hb1f0GsrvZHTqB+QsZoerY+XVT+x87alNSGG0EY+7kmBbUCMhbQyE3X0DG
sIKqyneMGdq3BGImkyqsZ/KYgh3t1NCJTJ+eldhY2WyK0BKzTC9qPFyAKMRTMDiM
Q5XldO5RuRAfXTTeo910zWmEdi4/Xv8UxgsUPO8E4d5+DDDUEMz+fWNYJXIQR/CF
CThoJcZv6ZpvkY3YWIQWNaeuYxokukioo3JKVdw1P9NSIKJKgk9gbxNDKLOjyTxf
Vq+eR9UZLHl0DJqQE247fNc8Vm5rlNqur6oFV6KjqZKrTZyA0cbV77wHEk11wlui
cjJP8exrypfNjGnBxj3S10ilHFGs/Hwih7obsX3pHN4EGSphd2xAE7Aag5jLgrcQ
V1U89mRVaU5HK+N+GllH/h40Q8HzYeaPvKPAPy/G8mNDFmp0vH5Y+Z4VP5RKIfKm
LPu2MjECuJAtqGIbdQVkVcx0SIFu6+pXjOZb6j/ZLL84EbuWn24dq97yHe1GyX1J
fTVBAn4CppOxttod0LDZRiwUTwDnSVXleaEQFjHzU0UA7IvFOaX3FajXZ5HLctjr
4P85uT2Hy+QVz7Ebwz0xrLjx7gFyU5VfIHRyBWcttWUA9rnpkwXVL3gwYZKUkoaW
7pm7lQh98ha8OcnxsWpfvodC7GnlORqhwbX81t1deM6AK5oxnJ4uCmOojqWHS0n1
uqz7xQzAKqm+ewZlWKM/F36xpNdQszytb+OrrpK7ZyqkyaU8q/VJLbiqzyDao6zq
fD+9Yy2HbvRb15rrfb+Olc2wC5WTCirOBmyRmcOjnzioQy9cTxe0OvMshc2hWQ8M
7SJ8vUI7C/GpVxvBeQMMX/hRPFZ2DtzluRhU7BWCACNxd9RfH7dHVATiE9wjDFAS
6SFk0BwEOM3RpykfQKVUCyaC8gpOs1oNOiZWV5DPOMT1/BpdDSzdITqGnmecz+FN
7naTuygB5zmxrYYEnYEVMEon1Y6Gk8Wqczprf0GdlxzjDFJVireqomaWkiz1Jlec
Kx390Ubp2TFFtpwCdVRqPkm3AGaHX5DyyDFDd6bdbXm1Ura8uDfn2idahfVD2eQK
9R6Se2/PILXJEc/m0yQnip/Kgu39eckwrcGvPc3Qr9+Razk2NNWuFPYMZuPIEVm9
SujRM4UoDnHo51n35PyhoEqRukqfA6pnY1BIuKu2XuUe13Ir5twGDAWQ9yo+1II9
xwB4vQK4XSS+URz07d0fsJFm3KYPplWlrMbgUhTsc/j8JntxLjMzVKw0qGrTyu6u
ob5d8FFOaYxqlQDuvtf0fxhqEuDpBZmb4b+lZzRxGkGVUyCUZ1LRHXldqshCQ+IW
oIBzMRLtqyGtm6+/I3JjUPSYDvoz9mdjl+jQEI1LqLz+w2vXeHttFhJSB423IiOs
bSixNYGzivyLgcXzxvw5Lhb5qC7z7DYTbyP6IoXK0MpHUcn65jLyX+nA0yj1vaRF
OyhbW0PS6ruByTjGYs1GB7Un7Arb90EOak7z3HP++tNL0+HOwJ+2uUx4e6+km33e
33RdxNBx98tVvf67UrJZdIYPoT3tZHJP59ivCqfZx9j6rq4KZnqfERxrxBobelVu
djMlEF3QSW2gfpxv4DjJ+A59aljElu3x9S5NZML9Hjw6f9+LifOZCFh3pj5i8T3+
hDopfejDjEURXfzChlKAg+IjplVkxRJ2gZqq+6RMcSCia5G3og8eb+Fpz/9rg5Az
4JjE6sU8QpJlJyySFS54DEe2NjhJAb+j6AeJM9yNNpsdw7jV9tzqEITxnD/CGawH
yKKM1NazqJZVG44nLhj4Pg85aDP6XEUNzBOalyPiP64vQn2/QzDbHEMip+8XM0dY
mCWinLe853U0BK11ZQZ9kj4hIX8cNLLuuYA+f1LxW3h57a8E89J0YTaU5DlT0GwD
093R8XDaEbuxEQCHE3Cq67NRCVslFDxd3I2twwu5+A7gbyPouSqlEl3JHvrqPJYM
l4GAdHEFURMil1qNJ0P6Qbu4RI4ON0cio5Y7G6jgHgJpRGpyO81nDRaaykhLs1h0
YZgvgRjbapqDRtXYxfyVKjr8/BRNfAJlxaAkH4wiMjfjaVWlbMnDjrkq9IWUJFQa
6ZBzszYblhup/Vdi4mAHjGYY5nd1CR6p8C+x2RoItH+g38w/4OOAOYkx2eDL3/ZG
pQv1DrSfYV4gEhOJNpaIR3LawxEvz8ymai22xp8WbnOM4BYSndsF8YTWwriKBA7q
Mt0o/5msc8O5KjVIrP8FQIriUc1mAnVRR3pK+G+mq8Nku2+J/+KuUG4zw2DaOH2Y
NzcZSbDV8HnB8CwXVP1aNKjuVDc39m760XcIYYfs8Shf+rmAsd37HZ9guOVC40OU
2ge9wv3qg/+Ar2ajtZ05eyB6ymfBDWMPbd95hl3pXXcPG4FGHVGo6G7TdtCdTNZy
VB4FNwJDXEc+UUVVF2lKxisk6doFtrZ1j1+E37+an7KFgtFHlsjEpX+dasLNT1U7
Vy0KGGdll64xDBhnE3rYN+lXevCq/Xx4VROD/W6E2X0GAE6EB1aXA/M49x49CpKS
dcSdZKbS6g8ImnJeAidnL77uPkeX34fZPuM/TlcwGHAt60WiVVwIb2ZwLe+YJ+WT
Q5v7OjQu8cC5feAXwVTz7+F64M4r0Se8tEWInwvhI6IcGTKw7OviKZFnw2VG0/N9
IH/jG77PAVHCkIDgFF34o3ip+FCXg21wBFxNMoIQ8ZloTLwe4SqrP+cW7fxV7eJ5
TlgjIq8a7zvoPBnIPmNvhdhWyvNCn4fiyYp+FOgEevjm4C3hhxQF39Aa2itJ7+SD
osRwwjOndaUAqDNtYhoDugNyBsmqc86YiEP7kwkLR2da5QpSfVM+IQvZyiwWm/mQ
Gkc2t7miwIyB11tp9XDglMOUv3FvBx/eSWis1CUI16rj3JK3siswVTpwYCz6OFOw
OcJ6/vVY5+M5jDA+endKFK5B3LQ/L/GPzTbcARZTUmchK3JKK6ZFO8hNmvJk5M28
dSqguxc2xNrgeGqRg1oXhObFQqXYvo0DyS9I+jirvhZJuJMQWFyzXFMB8WWO1Eis
lt/GRADqP6hjAv1JIC1W0xl6piVFDlCi7WcW6R+LD7A8j5LP6HKWolEcrG7ZkMqY
pS56FMInS/nZ94olFDp/SjTT07tpP1jlmWmZrYwOeMekV4eg53N9/sQs3wyKhH6I
tnVPevroj2YhzAEymWbRjrAH7VJiX5gtxOadDzuillTPzl3eEV/9adXMVv0elBWo
kJne+6wnATBahDb5Vswn/e3ZbnSRjHbZf2JPYPkq/wefdgomt91UYME/WjtxmkjC
ggetjQjHF8sQe4+Zkw0Fvhlgwwwk99VF+UlOmRJOzPluseUjjtwtzS+IOkOVFUW0
EdhKyn44+umJWkbIoc1vq1wYbwfI+z3PFdZc3JoCopSvrd9cV/ggQi5HeVdxqF8R
p3Tl4MBSQyKjYij+52EcGcVIFyJnrDKqHla5v9QhBRxJnQObYKf2PZbKq2qPQFqJ
5BdGZBZ124rW2XfFpedpqMz6sMS0BMY1gg/JLfE3/Qh9fV4lVh6/d04cY00QGTBz
64dc3Ujr6hL9HF6FoxT7trGOH2MeKVJ+ILvNvQzU5DZ+RVGad2UCgefDOEXzKn97
1+JWS1CDXWG3kSAxEtCcTolHG/rzhh0m6Fc8uOsPJ8cOLQYi5uGWpfcC0VdCEWP9
3m3uqR8MGJLpuHz9GHtPti32BWFlH3e6ZnZSdJ40WW9eWUoVa0FHVVwYOtWXoK2W
4iA0p81wNKL5JOci5ey3jOqHfhwtUCiMbOdmCB5xm5gF26BlqIAEpi9/xjsy4+yf
Sf22/iBlSi5/qO0u8EzGoUcPhcxoURhleO0CZGQrvChhy5co7WhWMoarnCgxRNUS
1UT9qdZIVz6se3U9Ke7blrxxsAgzAgu1x6NJlnYcPgBmxh5B3a7PV6lTgSqv0ALY
miJYINcEOIVfjMDEuWSBLXg+cZrEMydDo7F28IS3/JP96G6pDP0QMn8QyHmAX5S8
V7plzDSdEIMswYo7MW3hUSKEzvjfQCKanxGyoMMiU6YJ3eK8dHuzDgxFUklnonfZ
kxVutiy43jognCwhoYwrxaRbaV8vfu37ewhCN4QFnD1PGUrOGmJdtz+WtAMFfudp
H+JOesC9TsRag5yOIbbhtQKV0YOgwNiZ92E3sWLwXWJSqwnyDomLaE8qzHI1P4ET
lDPKOzZ6qumldQtjAFx2JZTi9gRT9NP+UL58ypUhIfMkCAycUv0pqcGXl0sd1FpR
JqUnAIActNH2rY/vWaD69nji6pflBSY9aOGiW6K0+T8Vv1rUnRwR2cszbLxbbnpL
XnwgfNDJlbkdtk7zFSe+2opqcSwakNHcD5ERcCRxxg3UfNzMGSqB4E4CREam/fxK
DJrESDyca4BgrZDbeWrbZRZ9PtUjLBeu9Zo12Qg49ZLL4E6M6IHq7fVtRW0gPVfX
OtArILXzZW1Fhxxc7cwOYe8hIx6dwUgaJtbkb9IBkNIkt9PAbdHnr/OERJ1OV2ED
Kkyvx6/k2x4xQqZlvgnA7DHBkt3OdSHGMPoLsJ/ZLS9vGheRZfzIOWqg9VD1/WlD
6KIGkBxQbRUgr9FuPjG+whlWv9MZxveDDmG8QVXnS7Y3hn3Z64F28NTq+57h3oCK
VnMkxK2Kgycq8ahQBgwladZeLd02sgeasLFUlWPBUskMZHzcwOYjw7BzaUuq3DJ4
7S03Eod4N09tb4PIIfBKzafyiZQbkqrx34V/VJYgeEqXfAXufqxQK/NyVoKmGwLq
QS4vNdOBdGELWIxUwpwhFXcdPK6bCldGUeRlEDekYButr/VqF4a3IhtJ46oAWY01
/b7M7AgvnyoVqZIYZzeU62Ac3lAhpqGjrOqP1p79oBxj6RYqBFfbLSFXDF7I1OU2
Uc+Cb4ynyj2M1uhkYYxp2CaLPzggaMiSVNilkx10c9mfY21PW4JGZlBhc03i7ea+
REkq4Nc09OhzYx6VfEdfvtTCbaJv7V+RntgsY5EQ0fJp02y28C50eKtlwHSCSdf7
GtNoFscc5syhR2em81IUt51TsxBl6pRKh10B8n9rtLijVU08Ede7BOwNDaQUr2JT
FTWCyNymB4JHZoQ7AySljn6F7YgO3AmhTwcWhdyo4vxtNR1aZbASriA+3oA/9DE2
KCJPFyifjI//RmxWH8TAxAmVGT9fEl99s14mDklZbPz/9dC0xRdwD7e3naKEhMoZ
A1dfvCFv2mUbE0oXwF6WI5TW3zfFQ6DDyHDopwj2JEdT+4n1N5IerRoiNXYizt5V
twjoLBHuZQbssqDqMOcCGjzhZePWq4Ys5TrSdS7rzrqlSXPztegwQDkSTMxtpWPJ
n47pGe7A9cU/1KWWU8PTeBKWJzac4aV8dP6v4M8bbKokVpU0U2UnGX4ebYLrgHuK
4U88Lwslp/c64+0BL+jH5bL66QwvaqfZXMSH54ooJ3oUk9uJ29bsXkVIe4Xj7Fm6
joOeyYMEc+bnPcBhd+t0rZSBU2y20UaJxftHkSmXE7xMKbN1zkytU4qwkBtUDdLx
iP/qyD+MfhMIoDkiel+kx0gAIo6B/ZrsIzbU9oZYNQHUscjM9Ki/lwfB6YQsr6Uj
HOuoRPbPz9qD8W5+kV66LVOSoarXn/+ksMwca6mXlwSqqGK2a3Z4qyrSSfvefkPd
o4lMx5X+75cnWznK9qAhy3gwWAugAKK9E3piAZu6EZqdJA/+tfK7LUxlKCgk+fv8
lJhu7hKwXenkY6LyGrp0vI3rn+FQlPA2KhfVrEzKWbky0yC8M8G4c3lA1hMo1ZQe
tA8rx8/QPSbO3at/9t7LktIxQOaAYmsbScdOFmP1n+4gqlLHokicr8DwErsOBSjy
7a+PE0a0r/tKlnc4drFHArWObb8w69l1TPAp9oeAnyZOcX9afAsbZGZjJatCmiv6
NtsRL2ub0feIyL5pc3bGWuxHbtW47cHet/LnThDfiJeCyJLYf1f1ZVEQi/KT30Ls
RvR0023Vk9pM2m9gJQB90YT7pYnysaxVhUrIQdJ+7GH8u5PaYH6TiU8WTXQ7awUy
4p5LPpqXyqJ2jqZe9yHKq4bGgE6eO6T0plnPf1gPBScWSJvGacTxyBL4X6frrA3/
xkpLj6VMB6RPXOO3lqOMoKE+6mvMLu4kRO+eXwOO5QjANaW0N3DM94kYoMs6IeqX
IzCNAnu2aPF3lhvjuJOLr+6uEVtlk+HyixulPGn1aR1Q6U6Tbe4oJdhRZJG5AMMd
KiMVSti12sl863iJ6IYPdhOApDXAcz5FkPqpRFzkd8xaBJZCg6bDEvzmfDyVdhZM
SID4v89kdeM9zK23V/a8NAA4YCbE3tXqpPa33D65MRaZiAX6HBhSE6L7TGDXCIdy
M8QUmcwLuhwIgJCIPnAw53FCigyKCEgcbFBu7rQXargMhk6+xpajjmIrczJPbbg0
w6IDU6t2hbjzhKOc+ZEGFc11RUcxEyBgk2wKzhFTHvooNXTWXjOf6FuSmSAJs1U5
GB6DXdQDHZEhxyKBkskvye8pIez8mQoQq4xBdPr76F5bfNLQpGkpkfIQknIwWvCo
gnve0kFCuHpS0dwvegzcnwe9qAwWvgD6ZCgMGbIK0/QE3F3SyCEtHIMeDE1dYnIn
1R3tPfYR9dXq1+hHLbAhAVDmUKHoFqhP/FniQfDoYL4Wr12GjfhBTCXjeb5ezhlR
SAtRzG6sRMvBGpznaoAuwtdg/CMchPIyiGuqwNZQ8eN3Yn/v8F44B9Pha2vvKhdE
pbVeJMO5KSc9NRw8qgvfM7B4wbKYWz8/Zdn+XNir+Kq7fZRtdcxCfUtvDHO5zC7h
tC9g6KHgiZbFbASQgLLFtRQus5ZFFl07ouzip+7SX/uwVpBVfT4QVmoaciFch8Tp
K7T6xxzAC2pcZO4RPKqlXDNiVx+ip2/dQ59S+yizAiV1iSTj2qf0iQxAaSMV/af6
KC5K+LisJl8u28J6SM4J4v5YfKEaJ8jNKwB8M+dljZQ1jAaixdLyoiy4tkAGtLiR
2oDB6iG4Dt4imaHw4ZIsfpZR+GsIcKN8EixAjftuDpVPKWxWXQGDuEOWhhfnumeQ
vzRxaLAOIgzR73Ai+T4br73osaMMjNa2oErq354dAe4RSC6uFB11XKKgfHHE7J3w
5//qb79hE4DsM//Bx2fKeWg+WEw3feh0EJbRpz+7lXbvT3XIheEYAL7uBH6oO0EL
yPtE/mvr/9XrAWfIRzJfsI4NwlYGBnGh3SQR94mVMUrnogyRwGubrsjxlIUFeSzv
mDf3m4kWcltT/9Q2r8aFYAs6sTXPJ1FF8eiHYi72hCZHupmAdqApnRJqzOg+74Om
+nhie4LSF2GMvzzY7X4G2nD0U6l6THyKypVo0eDsAqo6NmquNj5P2XmPJnSX2gTy
Wist2RcuoV7NOiPnt3AjWbFMcJvePhZqF8juukKNTSSbWSFky4E9vUau1eBJLQkt
ksX9LNtlyv2QrqRgxK2bFtAYlvL0XaYUklPcOKsnH1TSRAV48JH8wbOP4Yy689xV
1nOEZugT56Mc3xlaMTL3/YhQYQFvU2lb4Gc0rDmJoesiyLs8cDodFHh99zCEcuhW
rIztHX8Rc91XQJVypDxSwiNAOm4fxI/JoCbjkh8TDMigHYU/54Grv+U4Kf2cf1jJ
i3NC/tn4/n6eT/pwA0pUW/9Axu8wli/9sV1DxRfQmeI6RUwCAyD+BrshTSA8YkVM
Vm80FIoYvFzYSElhxwgNrJj5erZekWv0x2zdouh6c/2PKrZWbRGCBWLh1o5aszdr
eIkucV4ulUuOdXa9Z7Ujc2BEDLccrh3FVyPn/HGUEXFXHHyh25EDo1hewSwEHf30
Iq/7gTSl9Gqd0hwdm11QmDh7W+YGLmh2GNiKFBMmB7g6+jQWXWNjERgDLWk7KT/z
/pJI0CQ6TRNC59Yqy36Ur2DJ2QDt26gvFj5PgquI8tNHEkjRHicss8pkwaUnVw6Q
1aWcqManTCQA98NovXeD3fItJL9YC7Cu/xqjeeOu0ZEzxEh0sPAMTvhOb5IF1k0j
+t1K22yRyA0M2TTo2VSVe3es9Qa7xWUTfmw64ZWGzi+HP5yai6AH/EOtG07dnMJk
2INb8z++CbmLBWHIs4+r4QI8LjnmApu4xFRUOaVnwTiRw6AaOn3pffYs7lQMICgB
tI1RafEDMpEEJk7406vIq2wxswDJAY8HgTPknJZ/RGuDcg/nnKnCREkI0GoJ0eLy
+8a3uafyNBACNdMFo6s9Jxto0entZZ3czYSu7gwvXT3FnFasHOc4lbxHS/xnFdjv
sU+Nv4Zb570dlELdii98Lvk5quk93ZsboZLAnS3OBo3OJhuSL8nRMRB/2+207zRx
GlmmLS4MRWCyOD9WrUWvpSDgp+ZbsErkRYKNCWFVvPXDYcr4L5Vk/1GU8v5sKHq4
QePb3Y6hjJw8AAT8qcOK9Pz5dWzixdsAME8G5AHxbMMdRw4XO+hBsdNhng3v6VE/
BWsLbXpQiLnIsTu8HL6t150joIDC0EisgmKVhzmrd2BhgHZnxJLz9lQa+VnDDxzN
HTw6GliI7M0SrZ8YQAx4hRNzRJ+Li0jCwfvvfKWJa7l+xOb9EUZmcs7SYkyAuFQD
byXZfdgg56MBYFL7HJeHxlCBksT+NqaVofQd9g6PTjFmxB2Ol5KtQVDgZS1jEIVY
fI+PwgmueqjYbmTvcVNtQX97Q6fiI0CgfPqAk3qotYggjkZIXUx8iQ73YJ2yAHby
HyEx+UNYlJ3up0X+lhdElo+XAFggJX1Xypko2Ye6KNov8cNXBnROuoW2Q/f8XBzP
/SpDqpuiW5VjnEslVIACslu5DCMccdjWe4gPmOACTLmQzRnuAKuxAata4lJiO2kS
T+86Z8LSKkL524qQsawfjm2NCvuzUF0FovoLqtGicRuesCjHqCy7RsFSxzkOK4on
uRh7UW/vTu8W1+Sg1LSEc0TLKGdMfArNJDNk4MoGHBbMLJPdVNtbbw/pW7v3kSZu
+Hj2SIB2L+3pP6ljsKqFO2+cfVTTorfAmc7vkmsOeLeGHpDw/hutTnGnukwcTili
eBA0jp6G7hwvIyXMr62z/oL48BZHYuu3pVON+QGK/dJk/4opbUz6hyqClz1pcOXI
FszGLSrpCbYpvstUCoXC7rU4fHqZp5ZkwY8O02qdg0+Ma2z2qrfuWOsLnfJNvtZZ
ZiVvL7b1A3ZtIbxgdrMB4cVYikH5DLJSZObwDH5/esGRXfE9PbRWOc13vCm380UF
9lF2mpyjekMXaCW5EjjMQtU1nkPAKzRMtlX8Iihts8qDnbdDIYAGvDKevoVlhyZZ
UJN8r1MWYY2+obsSj6IBPrmj3WktdAYfxp1a2JsEjAAWfhSAq9bLQEp8d9TQYOkz
Zv/IP9VK4NYhf4YzF0R6PRi5MRE09PXvskdMyx39LP8RjyWSHBK6vzHWl7lqJgfZ
r5vitxZ+O2LZn9FIE3IkTiYL5fGinP9R4LqHDfg89DrmijOX8so9v7M4cPgdVc9H
llnCPBiGeL6rSYDOgwW1pEyy8eEX+8orelCV8NZml7g55My4J73xiws637T2HDi+
xnbQU+uWVzPKQwL68Rwd1MbU7ATSei++K9f5c7Q3c8o0JRBCKsXrAskvYKDTDkXc
gsNuG+sslALykJIRScJrhg+THcP8uC5znxyiLj/WbBY5ivpe8tuSY2z8E76brCa7
/ve3pgJ8opu5LiLO/7fK7lCxLqz7h5m9JSqouxQi4Hbbb16FxG0afO2KjmDdKwgV
SV3OP62/yvzTysia0bhg68soQDFCzng+nNpOjjhJYvDXtW1BiL9ZMEx+WI+A3pgA
QBCxfC4cxoi6/8kpfTFnQh5XtbFWqoXGUYsXcG/GPCeYKd5nHdwLJuoPcyDB6Lb1
XFxBHr7aEM2iDOqvo1w24vM5PGqN1Fl147c57drWhXQBGYd1pxOqeosGwqCkvxVx
9LC77vFLMefWx8Fzf4zbUDuHCGrEo2WayOU72rn8hlTK0Dc4OSc06+NfdfXBr2QU
gkrBFxIxP3Sihw3cH9/drZzPZqwor8iuZazpdBlB3igvYPLNSLgcByMMpd2gON1b
cSq047eP7/xUj70dQlMYAOZg/A1SoQw/v2abavaHJCacTPRMHucaRDhO5e6qomdV
gQfW4g3Xv0Ul+wMdMjiSuxdDnyuJEn40wQ/gd7VU6xm05b9oDbrqhgRhScLP+Eco
QwROo5KzUkP2KfvqvMyLlQ1U2GFWOdDx6AUaMCNL8+MZNzPM2PcQXiv0povO8jqk
M2bDtAp+MPY5MrauQgPH/b6V/IGxFMBy+DMi013qnA0LFN6vFd28Xl/slbco0Zb5
XGZ5QYZ8vkrUFI9FulAlca0xFHk89z6Pl97aZ1O+fJ4sAI0Fnox1z8UEsuhHjgHh
hZloCMYzOd/zpg+tP+SQAAElHWB41HUFN97EICeQ40IuNfGTn+VCfoatZhIn4RvW
XT3zxOMTO+CtiphbduXXmgreG6pF95KdFnENZQykW9woUMTI0wnOE7XFzffL3/sj
ZHekMMQzy5n1MBEIQ/Uc9Z5wZ/wBr2Z4VZNgqArs+zGrjDwJ2L/D/eGcjELHls6p
jIfdCGxWGnVTIYdEIbqb9+7La/bCuP9SLPm6Cbq86jlJvA0qSA7HNTM+l+hQ57Jh
h+3PwFE4K9YvAs5v54OGo5o/KxTNIxsfzIDWRvM1QsGUdMmNXfyY48KDnML9J0cu
phVx+KZNbINtdLg1M2adfxPKH/ukwGWew/lHr+15fC55+98Yb6TFuShfgoqzP+lO
4mEGgORkQyU6/mRHqgUbEb8RJTwXrTNVcd+6xGmEj3gUTXCUCWkGV78+RAsQLbQj
A/4Rgj9TnEeQ99okPW8Jw8K35jitHfosllh3pFX7sRu8Kcx8gKXDf+vnwOneHnx9
TDTJpcFMTx93Ls1bFCP4JWbZKuvhNTouMC+P9zO3mpJ2/m+k3ShzCXOF8e9Gn4Y0
NtwpaZGxyfKWr5LTXRivc/DfgTezt8fZS1wPzLcQRrSP35ELCsS21rqhMlMUE36o
oRvaJxHexhPaEaGuAGaVi/QYrPB2iy6STrOz1pP6MRIHjUOQf4kPCgv+2oxjGBd5
yQVQCLeCE4ggj4ABk8PraIO6E78WZmGvX+686sypjo5NZ8wrNUNOwSbAtAvuITiK
VRIQxSDtzH+mHAhnoNnrXfPMExKwaHrzsCnBZR73vnHV5qzopzGKqP0FLKAe1eeB
4uqV+FJ59xQcdTTnyObbiiL/LzSjzyjkvG5xAzDFgGMhIlmOwLWPQn2w5krbxGNv
uuZQs+Nads9ZT7cYsMWhfMzy/xulcImFYRVEF+zax5VfM2gY54G4NIUZhPUChpZu
tlRysk28cc8wZ0G8rtAKwbAsZf/0/x+7RBUMhKLrNSG+DOBFjOHG7zGw1rr5RUHn
GUM5S46l8SmTCdnL0xvAOEmvnuprcAa2Mal5H4b5ctTALtF0D2ObWjVIuwhooagH
v4Wyjf8DwSN//HWpLoZqi7c+B8uI3eYZ+wE159vhK4eC6x/Y8gYBwLhXkxV0gYmz
V2uIHYj908wdC9Y4PKbKl/0LnstPEJ5kh21GAaHSOoyUGDNjpJeIgbkst0Gu+OIR
QqjzPX6I+EUZpFLSTBg5jmkEFAARBOMPIr/UyotvZwJQX5TD0ItuI8YLFF2Vaq7X
fETgechwyGKn1ybgn2hrGpslS0LyluvUA7Mcv6cYRcl2l7DVOPGCgyQffZWojVKW
Ar9n+oKYJfqeic7KRUk8qZEWkfRTKPvt+dlcPV4J8oLrkI2aNhfW3np8tLEW6tgu
v0uYCjp0v8Ow5ikoNHWOOio1wSLibkYcMll/IpJi7uhqpr1lQuKdwkE80WHfIWLk
5TeeZ3kmu/9foB5p0fjrezUPHdXgQ3lMlfPI/5hpMT4wz2aBiN8np8P+qhOBW/Dj
XZRPN8HuEmBReu/j9AqnnRGe0hU9o8kBkEnads5s7wCxNk/ct99AnC5VoGG1xv1y
PsKB1TTyQBw8IWupv+SUbHCFQTaq2gqWp/Mw2iLPio1+ew9mu8TLpOWCAVCfZGfZ
KXjLhJpdZqR4hQexC/4rDM34I4D2kadXWR+nxPljRHQ58VkPFCF19WIKO7xGS6VR
v1s8YqtAwuNLjebgJJx0bbM0DxWhMVAhQhchLxtMEiTTrKlH+6aKPs3xc0lZY85J
qIHs97tR0pikwqnBN8GN3hKmZDkXkAPczbIrnFev2qqGn1q06FTtrvgSr2Ufv/XQ
QT4n5566Ny7rl4LI0CNXHXJpTBEXxH1uDmyrPgJheMvT9yZgw5jHsJvO+2QQKeXK
myFy0c2n7NBMQzTE+/gd6KW3ASLIl7Gssylw4T5nWO8T0f+V4YNkD5enhQuBBvgo
EixDyUNuc6Ul6myrKbfXvzDO4sG5wUUzIdbr3Cxc+skLze/Exxg36OoQAE7A17Vm
8qbvDQcXqZAdE/t1zYHpwdaPcPvXkcLbHHx2i957W5stoi9EVhSIKJ/0h2llJdnU
+p1O6d1wTFrmdcm0u4thg4/qDc5pA/8V+6+mTdMnnT99chcXDazcJ0hSLBjE2BHM
AU/Gqm20PqDrWol72RyhSCbtW8UEIST438ani/bI4OFa1xPcDkS7Xx3a0wxb0IjC
gpolv3zs7PVQJmAqF1ZoxmJKrWLGUQkgyKJk4wDUX9qcZ2MkaoKqDl+LxG6ZuubE
Wh5v5LpcJe6dVf3zAxW9lnzRw1dbX+rVHX6R1KTg4bWXe+a88XeMpGF6asWJPkLh
w2BzQ6I0BvO/t29zS9VSkG8+a9aoj0jOfiO+R4IpkNvq1ATNEG1HkCBPVQgLRZCE
NwC5kiK4RYqPosD6h2F8UTFYiHEEkManRINSgnh8C8XYAQR7LkQKh0q+6tPDUwlt
GWndxw3KMQx64/ud3vbXwgNcbWOR65biAQObQzsReICUerPKgIcfU9X3bl6Bhd+b
Q0fbxC6wkdp7TUB1AsvEokHB1IGqAV+ous4Ma7AA9flutX37yNZg0x4//4ENbVdp
zNm/meQHsVvfajpY1GpNJxc4lJzYvVoCOJDXxZyNPDxLSEpNCf3ovvYAqGII+LOt
mIv767Fsy9WCBOwj9CEscP9CQ90CUsIAyJNPidy3tJdDhe4pT2BJbZHfqQn3HDFy
XWVTbZBScNQ3CkILgjbOpyVd9hGDj74xek4VacAcq9TmaAKqptl3mf7vEvA3yaeE
goJ9gNefY+Kt3PHNsWbwZLaGduFj7v5BNrSs5zagk+3t+6SzRiqikqndL3ijCGMQ
pqAP6M+oLWKbH/SgnO7eankuBmmAGRaKqjzpYzxV3bFH7f2ZwBnZLVBD+L2TClgD
qPEzalauPtNcKkSe2fNnRrV7yrWgT5e4w05H7QXbLbBGFBQ4w++D66nE+KI9BF0u
L5YA5437YQe6me7xMOTzbQUBSxPV0jmM4ugvT43G6ljztJtOpivRreMuMEut4sHb
OB8rgvk/VIMGytbliSoJ+p2S+HnRTXHHYNtE1RrYZZ936RZ6sObrNqx1jyLK0c07
9LB2v6HqaOwx5hXrUoTUXpeV9W5gBCqmQJ8B3OzNpQPwe2OxfSzFjBwQpQhcCycV
n+z31Hh4PWrGo0uPZWWr9Rud35PQHRpJ7tMOtNaDG3YrFQcUz7oQvzhNxPRATaMC
QK5hxvSmApsqDnoHP1t8gXrb/Cq+wbhtWmUl0DfqtCUrnEsT4LtDqSwvSLk/1z27
U0VxWfEl2MV0m9EOfn6ObDzgPHhsSAdm1ioskO6+o8YtUxIAWYCoZT7lRobk4WHO
lVs5I7MWoTw+cQql+zhPe4MH6N2w3tIKyzyTJVh9h9rF9kqa35XUjoRVxJUgkbhN
B6MR8FBW/bv8oSM37ajTmdghKmalIUbeknsgAqlDaW9ZVfh3b3pK4rRxC0XXGiYX
aEXaglHmn4WVO/a7qBJk1GUB9snPvh6MEK0rfAn0yvoQhN2Eu7zQPFgD6588Gx/b
hOEIT//4nmlkcEQBq+E8PEq0vVq8LD4BosZiV44g89WtrvA6xyzmB/u3Y0y1yYRT
5w83HH6VvZ8m9yIstoUBlpOylt7t2wvlxdfQ2xpn700EEexjrl/mA4SULhF+N9c1
UqqPT5t2g6V7ypiLmSsXehUGYsn0DF5owYjGmhFaOsdn3TRybLV1xvI8wT8GPNQy
j1M3u5UGkoCyFxB+aP8QS823Nx/LsLpidy7gl3Ua4P6KZ92au7jP4UqAXL7qv+Hp
NZ8Ot4IvW3zndVXZnEjwccjACQy8A1CITBdxnuNDwXwmTdQuP4L73NU/1l9I8c2t
qG377cko0kME3Vh92wPOOwPv/mBjrOcdeQAdWz5Y6s2F/0i2UmNq5M0wgvQL4UEf
p+fk83O2NH+d66Xhh7jlcOs25Pe9wNcGRN408j8FUyq+EvgqGBmbwhdS9ttmfmbP
O6/O0wejDeI2l+CT3aRl/VSsk6n4WfHueYdiMFIyv/XKQRt8Nob6pUeE0l4//wW4
Tdll8QJ52strBxngeUGDonYJKdk5+ru44uMqULhmBzOnYCWt/bj9gF/QpJlESPeu
S3pdnqJHJMFX/AvuA50fANfCxs2Zdpn7hKXUP0Vt7GMMnIGPGT8C3PEGwrNddqwx
9CyGlvtFAtPwImkWk/7AEY54af8eOIK7SH1ZZtLdq2+hfIVQHUqJGssx5Tz2pxy4
Fdh6WaeZGUGk6iadWRM1JkcmQcVMgzF+COsuyuX8Vlyfy41/X4YKoy7pFpvai6Un
7CgGtiLyC1DDmtHXDo59QZPVJtPRGmJxBljMcmw/EtBJurC/0eAKxRpJ+DsscIWi
dQJRimlz5zlmK+oEpDu4aKk3o7oaxvirjA1ci43ZrSjrbsgJJwo0JS5QGdy8Ruhn
TuQA/1Ny98MYSpMzLuG3RHPml5XorQinj/ot0hnizRnyUryJ7TBLFSDQJ7FkaUck
ZCZxXBDN2m+Ki8/lvgyLOVmC95EcGMyYHK4IWT9llAkWq6A0ce4pYoIJ9ZJ7gFSw
g2DXTSmHTeb4/ZgT2vY0dqy6HASdVbLtilrtJjWcPEgCwfOHsofobJT2ETgK9uEz
yVqvSES6ACQzV3VTrerq8ZeVtGLU9ukgqrnN5h1+Zo6rRfSGEHKo9tL1DmuAnOMR
/qBBpG3eE7D/1HzGRSdhMnbWV+Mdodecg3Xbn9cO3lDM97T/Ua93MgfX3p0DVm1c
u9KfxLfzibWUKDoiFKM4JwPAuNqsLlA3nHrwBRxjr0wVxhIFVmHgdCZZbAaFGABD
DueO8VZDLycXmIjJybVC+fAuyhmc+PEOTjobFlO59OWZZhnFATLQ4FmsySKHaaT8
UYtNlYBAHpASh1FPXG4ht6DwDHk5Yv3xob3JCHSSuQs/C0yP+byK01hchQqIJrfa
s8ucrTgY48BFSvoq1be6ltg7G9WMSAN/Jn/o7MK+ua7bXNP1uaTs9fbPSdFQgUIF
m1KtsNf/7OEW56CmNijFk/CkNPPOp66y03+3lamKkawTbVlBRC8U5O/mD6l+/BEC
r9oLIHXmHC5xASdk5Kv0hpxvYqoc2TTCdGRTiK5VM2ziKqDKKv6Plzd1tnuUFeUL
cOdIQCaKxtLjSxc97ihIGjjhNJvV1Nc0wsfUnJWbSObNKjoNcWeD9slzx29IXkao
QfNafpT7pFLFlzU3geTsdhNREakSmXawBuVGaxFpXGru9Czm5eZf4WpDxitSE/lH
If/qB9B8R9o4iN0eaarlfGnD2z6DS4zFIA7Cr7w6BGQ4CARDG6uAk3Q/91itwA8T
knpB/yD81AWjDU34hMMC2W9hyPHxUw6Dx9BWdxhOJ/dQ2UQNPuy75p6MG5xV8hPh
0GkWPXFdcKK2Eqz7Tq04QH6+dExTYGRsykdHO/z32+x9AQ9+RRjBWJfkmNdFIJs1
9HCJAT6t3bjsZAopnsy4nkh99ALGWy+22uOlnWNB2SCYJp9kzUsZArLKBBzPFjDn
G1iwrMJ/cZ1MXzCRcLo2pSO44JbUJUpufUSpw7wThNHyprEYYsEGAb/PjJcGEGSU
msA3TDU1MA7T4p3X8oh1xCJljKJsSHG3Ht6hNYd++oPX0VN/ssgbf9FamllN05P/
bJzxepZwYre/6vBHQtkZvL9e2XQguBBzhRIVIpUeeQfpnM/qEDL/Bptw6H4J2gto
XiB7jaYKI9sjofof6fepn1Fkl3moFSpLg1qNQA2BORLrMXmjQQ/fHXNV9vPqpdbI
sZKeedFdBzF8av7W+fhn/6JbcV2K97KUjJNGvi/BTUOTNZ9wtYyohNEJcGBFY6d1
Ke6NiFqYXrJUn+5IbC6l8d/l/Jb4xRva491PHqbTrbbmTMoq+eP5AiE3szLCPS1M
qBims6kprusZsv5x4uJsY86E9HM0QziUWaXeU6Je6sYcHIEGkbcTRhk01JETZlgQ
AA/40g9QlO6DsnN7eVGOOW6BcwDsTzXAvtEnttz0Lo9mE79mIruUC//KODAVRs7/
lmaqZlK5NEN3Ie0a1Vx8NQPBoZIU1OwtP+tqS9gEf+iMNheE/7PKQ6GTVUhsaR7i
UumBYT1gWsS88xAfR7xqwlqNNZnkgBYnmL9W4zDgD0hPp/g/rutjIjeJ66C4ygnO
BvdoPEoxHVYaA+C8OtmaxinTjCkgOXQdhfnGJiAEiMMBwgLP26mWA6cL8DByXumm
0N07SvjNJZlphHbTa3TwNNm/36ApzBMT5PIIjGSjZ30gxB+TFDA4FPi51EPyUDWh
QvakljtuLMHaadmJs7L3LgUC4cLagaAMd4QvbWkkDIYk9y0TkUpXe5X4YJErxz0a
Yue+sRikXS2nSijTy3+u38vH4+fnpcl7sCc5jMW1/5q+Yq3qwGF5bQVWheUPFEB2
KRDqo4VVUJcejAygRYaLyZPwQAGcQ+TQ2kVqnCyvoiuZuIwXOL2ous10x1LQvpEl
15XminjdwAnWsoXILp2KC53d8exFVNNmk4Bj0PUiDNx226Q+If74WHJBkxr6a1H+
OLSqoMnOdDohxXr/VpbV8YqMHEf0BbPW429283LpXF3VRtliEe8u0V8iOgMkw08/
BdQi/zj6oLeup6HP8MplVGwrH4ie3O+sPcYhO9e54wS70e/4amwMAmWU8/nl0z1M
i2hi1wpRrE9ACxWInG7s5YUIKjbXVUXHm7FKpfh5F9NFhCIq8w31e7WnD3sp1M2W
DJE5przKFh+tGMTnbgiSwusdWWT0iPIwwSGeJkJ+BEzoaNXiuzB+hic7V82Vn3W1
qC4FxxXeT8xdDX0ES4v9h2LDOV1IOHT020OLp3Xdp+Ch5SJpUA1PNT1sBEb2bR1J
8WVssurLUX8DB/GltwG2vUB1mmuhww998InqsD6HvP8Vm8cqJISDKDzOHpumS5AR
7YQ7buq4pQMDNyLqnGpZkbUis074aPOJlEXLS8yLyx7i9/HQnZyDGkNO5nl0+8E+
B6IYRImo2N8wpHH1f86w8b3jnaii2aYdwcLV/o/N2dzBJIa7LoS4vAcXonhnl2GJ
zzYgaq0MeMOC87L5abCAXK9yvNn9wK/9wFrPXTr9kg+zHzDG5YHh3rHD0zNHLQ9j
ThoM0fb3w/F1pB3tu7FXXxdSXKXoNC6eHRXLZvNR9gDVBfZDoLnc6hDvvyK3NXvd
jhHn3RH6y1P/G01vqmSRVxBm9vsVWhpvKsVWgTOthxUFaMF8//o6959WGXdIgITS
NkFhHzaD6SrsD4a1gLTxdeoxw2uhKm3K1d8FtcNPINO/5D43ZoweRkqUl+m+E45C
ZNeumNopVSSolgDYtV67GN7jwzvLD/RpmbtDWmbjftdhf0SCUg40zOb4iScmiN3R
3ewEfsHeoqLeEF0iKDjm0x97x3VOEqBBwukihIsNq5EC6lSZmjSbR1/BVlOLgzbd
GpwC9/Ys6CkfgRM4MOwCF0sYZ8H1E6hr1MCaCs8R5WV05KHUtIcbxtji6tl0aWYs
KgMKP+gihMIJEfsPM6gzBlVGoZHqUFHb/l6duPB9ZXN+Fy/3RTEqFvma8QUJ3z+6
OTHpgTdQs0am5j24pH1OaPkw6vgOQN4RSVOwkVTs0FAsI1JxCI0+A4hu5yabgHAz
SeEm00Yogima5N1f4o/N2nMjj2IybznT2yEKUdZ3wjNQnF4KZUOYbed1DURBjROU
edjgagyvrNxDtVWKoNbE8UGJ6xaCXHLkp7mCS2nDaXESV67pVCjAuD623lVc8Hnb
06QjvFrTZnZ2/6lpJdrc2TCWKBuqtqwBlickgs9mty54TgWdt7a5p5mpu0qYKG4p
eF0d+RvlFOvUmp81NIzO3xl8Odbr+AkBa4u32EtYTIouDP62GBbHPtannF3jnu8O
/LBV7kKZvLZZH3VIHuW5VKAtKqOlzwnMlbplsIhcj5FRmeaFbRBemMb+06VSTJdU
GM9+cHVGsTvXjnY4KL5bcfrlWrdF7CyS7o4HtXvlldKDmzzr4s7NeMmcJeTUijsh
rHr4yM8Febe6AGuBSu3t9DWCOLbjnOhVCqtP/oa1Zbs2sie0YX0NQwUp8reTOD++
NfF/NLrcG+W8pmkfypjsITXAQ3JFTVk84nt91mNwlCT4iK0lcjiMIIOL97MDPi4v
XWU9qrP448sjQloBFADKGmIW8VKs0ZM8E8HXZ6yg1pNSzIPnE2G1FwbiLqM/l2sq
SqW6Oq7wrqSYygv4BKjqQrzT+f+8UnV6lnHMMzXiSOHoNCDrKv/r6k1h2VLFCqSW
u67nFap6NMv304isImLVpMU+waZLfkB5B1L7Qu3qJYwdhaebWhwnEmoYHMFnh76r
vMK0grEM6YEuJq/JssAU53bF1JAQsdaWCg5byNNUsa2gT3gSK7nHvbzgNBfQ8NcJ
/yayMKSyvBCiaLR15KWC3JItcWN5EYy5Nj8vZ5DNGP8BQkVaxad7dTgv66fKEviN
PyfrPzeejvjm+S8gACrQ4zi8+LwT4StsbCIZogeKQfFahMjCnZUglrJaEy6jU7qo
8pI1XzV+fYdDHipe1UsHdFVQuhzoFlRrkxXDDM6+EGf+MwyjEXaPVbgtWM8JYhFD
AGyzqGN+ZEtDUfgTjVZXmjWQQIA09VGHq7YJE7rxpThNYPvB1c2FIzpfFRBrNORt
IK4IruNTdHtughpUnUqm5IH72N249hODwB+X0/9SBjIXrtFNaNQYb+NihT8Pw4Pp
h5/BEOaiSJD0Ddv9jmXWDzkjR4IcrU9BF33Iezb/iHxpYBCJJYg+0UULsbrpkmr1
d9bPD6c3M6TdA2wyjgtUJgAOzAVtb+yP+9ltwWiWLMwrTT+JKOi6NMDpdzhHPAC/
cBYxw1cdoIhqOHP8AnZ4R79l+xXZiY83f+XJKTyPt7SYniJe2tDBed9SPYo9f86a
m4BgTWRGK6zX4CWhEuyQJt2l3uPmGVXc8BSAJzACcN18ZFLPmz6551UJqZqpCjNU
cgzbAXvet5KJV1ApXHN4GY9XXibQisFqwi42VgC0klaLXVlC8xszIPVGWIrimEAH
9vmJaSwW96sQtCeu7u6LEkAC0E6nC+XyVUREQQeFzfmiJ8mwaPwh6nBBHNYZl3/Z
VpTQCr1V9yIyjOWlV6QGgwWTG+l4VO4XNuUya798wtCBDVInoR16NfBWYEIjtL3I
aQMyOLY06TLzy0WLkLA3oQM5yaOE0WNm/m+QSXgwoP8FRnJtL64vPq95LXv43Ew4
Z+waHu/C6TS2ZxU4dORYLc6bDK/n+m6h9V2FCR2rgFtSrGKliPeqFT8kZL/N8HHi
eIfnRKws9i1md9jNhjx1Ll15qe4ipoflBaZc18iiVI9hxgTl9xmhQSo+35t/GehV
WuVSYsS6wIQEvnyZLyrYNK5vRsPs55EzcGj6TAeEX3dzq8EOoIEkfUn6HDQDZ7Ub
N2AkMp9MP9759jGmhiX1XtfIF1zZWuipGY2AG+8/Z5KHaiJaAkftKNWVTtexK1vl
W/MTAJpg2P7UKI7wXg/0Y0l7q5oZwkIUx4/el84Kr2b47Lup6rf0cb+UQBXpp66V
8y++RIcn0m2ktmH9CerdHeFx42l+gfD5v4rvA1wKS4pT2ib/mCWyUV60GNnWnhpS
MN3sFM8vp8zPvFCSVJAq0utvZAT1W4TzEB+miHLpE1fgHNb59LfpDeG7Rzmr40DJ
x6VtpZMP73+B0ON6e08JuOx9POF7l+Rf+W2hPt7IHRFMkTXtpKL6Y98k8RF0fWo4
I6sKzkWlS/8etQJn0XYYh250dcILXyW389bhwW3pb7Gkepq0FU2nnp96wDZbWwVv
c8Q9PCoj2L3EF004ZbJ9MbeeD1eIrVCypnYTrZboyOR3qxrmKGUWex6ds90V2bHt
vFvxSL84/aE4ToIK78KasqIcWu8RPcnriarsUT6xbhMNwheGNgq1rDV+B67F3Kwv
xtMU/0tdNLFWhegpkuZfbY5aahCa2uAsD4d74Rz9mVVn8wdlVoWfC1fh1iu7AqQz
qVhFepi5YC3m6h2YRgiiLfElVnRZC6wX2KP4HA7fLNgQLudWGxWy/BHWOWcV2rWN
BKzAVzdpQ3o+qqOeyszlTdIMfmvMR3EAgPC0P3k8u/xNZLNezCCnAnnAjRBAse13
0en5/KWwpA+SqlHYSuqnxPGDFaOzEOVQnzGtEoNhuByRMQpaEtbWtGIbLg6MwZBl
kQ7Xp+jkwk1np8JmhRyYodOXPiWmzdkVoEsK9n0BvLzMgnk1j6Vaddc3J4a5/m2l
LzlBrgWCC76MKu8newD2NjhGV4P4dY2KdIXpQlWAlDFXvynQdF2FBhs+tFWFqOE7
9UrM2i/q6Py4IuW+s80hmYzc4OkyXmHIzp81IIwmhr2Ixw5fTPqjX1E+N3LQyffY
oMt9e0IPKHB2giG4acFnvXUtEdKoHqUhh92fMPeHZAB2z0l22TqqrIYMy45P3C8A
h+8y/IKnBTjy8x0ZDK5vNINyGOmFE/OrS7WfqZaipPsasaSwbe4xGVM59jfjC+Nr
X0K6nFwYY1S2y4c+z/Qze1S0pQNzJiocXxUGiv+ez5cKpxua882/YpJzG2aQbeGX
AoKtF+9H000hAQfuznU9TdGXm2rInPUh0UVuMND/dKouUozpYcyUhrOq0jhXMJd9
pMRZ4LFW5UDKkk99+qplZQngMR6Pfqm//zNPVPXsCkOi0SBA1LFz3tGxFeduAh6o
hCP0unZFAkRAR6uxNcw85L20YEL00M99eZUXX3skndfBPcKfjzOWT/n6FIiztLZ/
OB5FNm/cmoNXzLrkZdCru3jSvmRVpEbZc2pWh6QnRU6OHF1gU/XbhYKvimIBxWVH
7FFGOTBHRTume6ms8vvHt5JLmnLSJE+aGwSioU1gTV2bTrulO8u6JWshV5SGXMTJ
gXkN64o6ers3eGxO/Hon7M18Mo+ryOuOwGw285++Nhwf04lMaVrRo+vmCzsn+Qj3
FmrOAqlaoS57QkcpYrwI8mD+7QF6yJjk5lphiGVQRanSO3s0TrxwRmqw4GSBQVVe
O3WeijXSb41/g3ZlHc1uLnMg+sXwPS6iDyXqrquFiB8xyjXBC80rP9BV9UEvqGCF
WK6AR98O/9zb/r3noplsBlqq2VX2nhdye3zLnedkq127I4AMKDqmvRXchMla0z5B
Fbl0RHVKuCGa6Agm4a/gI7xP4I4EUFlxQl1q1bA5h2dU9JpkCCFNnfeOMaAJKwxM
AyjQOHEExkokxl+DtDHTZKp3t4y5H8vLiWuQBjlb62QvTdRFORTcBx3wKs5tH9r8
FZL/YKnxhgE96MUpJoH2o/a+iBMWKsHhDd4s1JfZJR1y+vP7DqshwyIeMGBERkwG
SyObQcggwtRaWYXSgwKRMeViqerbNHC0y+pbp8Lb645W3Sn2QsrlCye6M4E7aVI1
P/zfvA+iKy7yhX0ZL3ckg1Zb8uQ4ZmR3X8csdl5N0lIpFSH+Pm5q2FSSmwpsPgeU
ridzv4cjlsbzOVTzoZuxROoRopr5JMPR1s8tGRTA0NH6fZXPqzOMeU/S7xTycOal
nDdqxRr+RB2MyokvzN95P6gOKvjWbeDpr9MQwQBLCa9Y4FNJOz4sUxslAWe3b+8c
v27EDrdGhz8D8c5fZtoaU7INS2OuX5LA7JxsO9oH7sBk86PoIoCYv7ypXmpnFdsl
wcDwW9tHPJSxRPf4xoUriR5iSAy38TMWIwilZ4gTCuWPscoVCuoacQMkCdqUmIbv
e5tA8E7hjbkWrxclSfWuXibTro6whfIgJ0kAbE9d0OafKiyDqzLQRxwPr47KRukJ
Qi1mghjv9NDK9ONbYr6gBizlPZeCbswxQtmSVxxnAOzkQNZQ0xk1qzT2ZlmkC2lf
6Wu8GfoSPtS/WtLBgTORGUPZiBl7a/jOoqjO8NsiwFVH6op/sasJmQT3eWsAaGtR
jEsNK8Wv2wCL1kHamCfp7D0mEy8wCj5uqaFyWQSUZb0OGNDJHlaC1Np28ZqOTU4M
r4PqoNi8Z5bGPKRAL3VCJveyCE0Zcn5wgVVzkr+RQKTnYl7msYw57sz5lNjDhuLw
WJgH3/LBXjRxTw8F8PtKYG9a6RUtsWe7VpRxZ5OcKkLTVMVE576rq/1bxdjhenr8
bIk5rYgIboSBj39YBjMn+1EixwxPmQEWe1HdvdcjpQcE0lO4jJUV1o50vly2LePY
UV74OX7AlYJarG7QFqHjbMA2Tx+ab3eE9EsaGHcdkxxiuI6fS4ffHLIWjgr6txMD
oqfWxfKutSrsB9E+bXBTuWPDewBirpKi/+J51+sbVIxbk53wmkOHbwyqQmVfyl4X
yLwWyDwF5YvxZyhIhCLrRBTy38ALeXC5uVs8u11c4u3Glje3gGfCrmI5GDDSlZey
4yXoAkCTopV5CxV3cm7DwP8H0zHn5Czh2/dALH56VE/w5ornAux+22ETV98DbL85
XQRT4+Mqr7ol7EcMhBCcWZq3Dd51gxd0QCBJDth9PToIa4gMMxcm8dHUka4ZvItI
8AzvqKwvuEihskYBge1CDoEK+PPcuvbXKNaj5HoHPJ0KX6SuMrLa5ECi2ZajLWOW
A96IAyJFTeruaE90t594dy5qG4H3gqxnxYGq1/T9qksJoOfY5UbFSXj0J+OFpN+9
B4Y/QQSAbDNrbBpt/N01skP9PONUFrOuQahMBEVrlYdIHpCT5O7vTsPcZXxx+xrY
5rJKe6t7Xp9+SPoOYSrQsrupZp2nWwc6xpBiu6dErpOVX7hsS0s41N5/LPCwiY5F
lSxruPYav1iA3xZs9NPBpLtZtnzJzWBgRqUUPxuw7DvQT53yBuR5XqwHf1HWResq
sl2VaK5ZXEQUUiQIKEmTycVp8tuK2HhKNF8XRS0LknMCn8UygVR23unC7RyuAo/G
JvrN7BxUFT3seawjHbkD7oBUcwemW4V9Nt2wRGNNTcR5BJzDpKMza29j+AEwneA/
ON8TI9enEeePgSu13JtlpP5ToDglE+hCDZF5ubcFN7HB8lEbbONwRb6726hF2oDZ
rKt1tx+45bEm/HJBjFpehQhYEoevBGXa0ICYyQPnAjgDMJIxplvYKL3HgQYTFvsz
MUUjF4m0F3xPxWj7mxgMkJla4p953xT9VtEOjEXBWr8hz2Ly5mErbRCFOzFMQ+H7
8x1cHE/UWWXstZ+fJ54+mVvRsNh6PqcaUp4IMryGQInZxxt9gZQnY0bX7BWVK1K4
qeS9HzqqnQH6Mb9Iot5jcpDEs/3No3+9793Wj2tVVY4MoXWoXQND6LfDrU10RBIL
tMf+W3DG+f3BEqLR83I3ju58Vmhe+I+VqqutBcgR9sI0A5bAPZqyhrLbnuOhGBln
gAVB6tJJGQiTuHBX4+zLzIWvcY0r025RCON5Hy4kIZ96Po4aeuFMnbFDTq/1+0qP
v7pipsWjfG0u7ruUp7dAW4+jWpYgRSJOapWf0stiHWLaocJRXAOpZmA5sSSjslDi
zmVZHjcV4saDjr35GhJyF7d9qb1hJfL99tHvlWVbEeVnxb7BTwHJJJ7tWllp66I2
wNVp2IssBRXJsGnKPksgeyeg1anEOC2Pf3Yl5Jmcr2jlbM4iUpknvq1alUGn5a77
7vPfR7fNPlQR8Qrzr537foizjr/u4dkmOwnh2hY/g+wtOrLQ89o2N49a/j8GlV1j
vf8hsfOqzZy7QFuJDCpiIuukOU+d5nfvf+7oT5ldOPI2QhBwlg2FV7iMlMk8r/W4
50MDPrk3PXPy6ZYaXEL4jM8cqDEZxpXVUmPpfhj6ISsSzYgzMmpWWkLzP/pNId1R
DQOyzBLs/WdnnT9+24nAo9ioz1WjXcb4ur80QknzlhLbhbPw8XVbYpDTY4hG8b7/
q81RfphQ+p5CKTiBGTJHX10Iiu5UbmLbDpoGm6oj0hrFMXX0bqYhhp8vS9UTP6v6
VvKsc0Tn5VR5I6bBJA/Sa4dBnW0yzuWktdhuTZVTUVh8juq7377klwJwdK+dLPnT
3GiT7owjQkN8UWowJd81FRVKsYFjdq6jjXnD+DPfKm0I6xTuilik5WPbfY0KauTb
vKQOoNhJtN6N6JaZzcppG+ce3Vni5IspCLiIVVQHRFRh033BKXMWN4eWjrVdGsu1
d9SDlGlOk/lu5yTxVV8wAlwS60IzMaFp/yCgfnzDcWWtOuuGx6rGul8znmS3x9e+
2UKRz1hEXxXbb7tVpXj50QRuwBByV7EiFcAJljqw3eTUOqVvx4m7+u8BSuSdaZvD
JCfP82+Jqx6Knf2r3UEhzrMKNRH/DR/q7Q0gb5mY4/8amZoeKgzOYfg0CNqtBaYG
VAOEBRhUYoy0gOAL2M3rjuXCdzRCfh0FX1l6r5/ZKHqy2yUhITwdUHxsG1KI0dfI
on6gIROZj3EbvEgbiBfoCWdf0N0cmVidwDDATysVvGkce5/qphp8PSQb0IcwvUuO
AD/1DunWT0J1zpQ32prdYO6midFks/ylnfPUOghrluYsBKXdL671f1kOE3kqrZi5
Io7Zv+9kupd10YphBi/QbdFjvXkjyfsWQg1WSN/fnpMCdW6Sxi/h0HkeJr+9vVbg
+Krq/vT3i68sm0aN4WfH6pZdm5U37T4WCAQP5rya7uIi+ucqHwjDu7yXSChxbpcw
jDtlwQz/ETC7Y89dLiZdQgCQZPQgXTPHdxMRxYC1+k1XnCm37S/ZVh9swHvIf/xd
DfdUiM9Nm2pg6BxpCZGmikUTvHXrRrfq4gMXf6A3mvPX35MRbH364CfUe0kMtvYw
q181PUDYPjnfj2mXJo/kslb0uJ1WpfFDMKipuOlfOLcit/fS5QM8+3Ditsc0cFiD
27WORdgFLpmqsdlET1msN9IM+viutaZfYS7JWXvbjIWLMW7ytv3+VVUkp3B2TIX+
Ey6+19VwSUTRr7Qln79SvhXxRMVfZjDdIHNu0iA0FX10/zL98snETKi4ctvT5vhM
5IhskdW2HWxTNKPEQH40vFW82896JahNLhRbw4M01XsmzBXt206E38BNJocuVGYN
TANa31UxWvQKLJrplN6Rzhpm4H2lxKxJGo38Tyjjshv1wey6WO/3opu/14Outeyo
1yjDlcYzfNSN6OSma1C0U54OyT5yjoNwnzEl+n5N+GuAGbP3H46XmIGPbJTlqbMb
gcH/frXvv2Xhe7qq3BRgkia95dIqW3ilPUz1HAslreQp7ja5R3K//xEM4O8pm/+D
6lLM4oUhYxDL6S6uNZAIvxyAr527KWAanJav8Mnjw/a5HRGQ8ZJswrqWxDo/jola
rAsQqTdkGsx9aDC29zQtmchfaR3yxK9v5GIAWXj/l64i6l+iYMBuhbf4LKaVmpmK
RGTCQzh0Y5bMBGLpmz+AjUheCRrJPTe43ggccLBhb+kjk759O/qEBe+tp9o8bZ5G
2iVmlS4ktc9hdFXXTXC3Mt23TYebM37ScUANeq74Xh0CzKSbhKaxnixYjD/f28xO
edZ521gVsS3aCajTna0PNNnN86+IEbXNha1NQsEuRzD2qNJxB6atNTh/gAtcVVIS
QlVgT/ywEFOt2qWN4bEoGenQjTMAeyI9YZqYZKf56heICx+9DcebkAMKhxdxz2Et
8rNFmuofgUQJ6KlefqIoWAJPupTNEDrOWEJlRuDAz1s8tD9fun23PeNMkD7wLpQm
qApc2KxGBm3X5M3Aobi20Jakb+MBv3BjUgbKWno5Mop5C6lCAO/UnHEIFcaKdadQ
ROvOwRIAMIjlMP20vO5YAyS4Zza/3rl+r8N9c2eC6EzlbDWMqUBdwK3uluKjx5Oc
`pragma protect end_protected
