// megafunction wizard: %Audio Embed v13.0%
// GENERATION: XML
// audio_embed_top.v

// 

module audio_embed_top (
		input  wire        reg_clk,           //       register_clock.clk
		input  wire        reg_reset,         // register_clock_reset.reset
		input  wire        fix_clk,           //        conduit_video.export
		input  wire        vid_clk,           //                     .export
		input  wire [1:0]  vid_std,           //                     .export
		input  wire        vid_datavalid,     //                     .export
		input  wire [19:0] vid_data,          //                     .export
		input  wire        vid_std_rate,      //                     .export
		input  wire        reset,             //                     .export
		output wire        vid_clk48,         //       conduit_output.export
		output wire        vid_out_datavalid, //                     .export
		output wire [19:0] vid_out_data,      //                     .export
		output wire [10:0] vid_out_ln,        //                     .export
		output wire        vid_out_trs,       //                     .export
		input  wire [7:0]  aud_clk,           //        conduit_audio.export
		input  wire [7:0]  aud_de,            //                     .export
		input  wire [7:0]  aud_ws,            //                     .export
		input  wire [7:0]  aud_data,          //                     .export
		input  wire [7:0]  audio_control,     //      conduit_control.export
		input  wire [7:0]  extended_control,  //                     .export
		output wire [7:0]  video_status,      //                     .export
		output wire [7:0]  audio_status,      //                     .export
		input  wire [15:0] cs_control,        //                     .export
		input  wire [7:0]  sine_freq_ch1,     //                     .export
		input  wire [7:0]  sine_freq_ch2,     //                     .export
		input  wire [7:0]  sine_freq_ch3,     //                     .export
		input  wire [7:0]  sine_freq_ch4,     //                     .export
		input  wire [5:0]  csram_addr,        //                     .export
		input  wire        csram_we,          //                     .export
		input  wire [7:0]  csram_data         //                     .export
	);

	audio_embed #(
		.G_AUDEMB_NUM_GROUPS        (4),
		.G_AUDEMB_FREQ_FIXCLK       (50),
		.G_AUDEMB_INCLUDE_CSRAM     (1),
		.G_AUDEMB_INCLUDE_SINE      (1),
		.G_AUDEMB_INCLUDE_CLOCK     (1),
		.G_AUDEMB_INCLUDE_AVALON_ST (0),
		.G_AUDEMB_INCLUDE_CTRL_REG  (0)
	) audio_embed_top_inst (
		.reg_clk           (reg_clk),           //       register_clock.clk
		.reg_reset         (reg_reset),         // register_clock_reset.reset
		.fix_clk           (fix_clk),           //        conduit_video.export
		.vid_clk           (vid_clk),           //                     .export
		.vid_std           (vid_std),           //                     .export
		.vid_datavalid     (vid_datavalid),     //                     .export
		.vid_data          (vid_data),          //                     .export
		.vid_std_rate      (vid_std_rate),      //                     .export
		.reset             (reset),             //                     .export
		.vid_clk48         (vid_clk48),         //       conduit_output.export
		.vid_out_datavalid (vid_out_datavalid), //                     .export
		.vid_out_data      (vid_out_data),      //                     .export
		.vid_out_ln        (vid_out_ln),        //                     .export
		.vid_out_trs       (vid_out_trs),       //                     .export
		.aud_clk           (aud_clk),           //        conduit_audio.export
		.aud_de            (aud_de),            //                     .export
		.aud_ws            (aud_ws),            //                     .export
		.aud_data          (aud_data),          //                     .export
		.audio_control     (audio_control),     //      conduit_control.export
		.extended_control  (extended_control),  //                     .export
		.video_status      (video_status),      //                     .export
		.audio_status      (audio_status),      //                     .export
		.cs_control        (cs_control),        //                     .export
		.sine_freq_ch1     (sine_freq_ch1),     //                     .export
		.sine_freq_ch2     (sine_freq_ch2),     //                     .export
		.sine_freq_ch3     (sine_freq_ch3),     //                     .export
		.sine_freq_ch4     (sine_freq_ch4),     //                     .export
		.csram_addr        (csram_addr),        //                     .export
		.csram_we          (csram_we),          //                     .export
		.csram_data        (csram_data)         //                     .export
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2010 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="audio_embed" version="10.1" >
// Retrieval info: 	<generic name="G_AUDEMB_NUM_GROUPS" value="4" />
// Retrieval info: 	<generic name="G_AUDEMB_FREQ_FIXCLK" value="50" />
// Retrieval info: 	<generic name="G_AUDEMB_INCLUDE_CSRAM" value="1" />
// Retrieval info: 	<generic name="G_AUDEMB_INCLUDE_SINE" value="1" />
// Retrieval info: 	<generic name="G_AUDEMB_INCLUDE_CLOCK" value="1" />
// Retrieval info: 	<generic name="G_AUDEMB_INCLUDE_AVALON_ST" value="0" />
// Retrieval info: 	<generic name="G_AUDEMB_INCLUDE_CTRL_REG" value="0" />
// Retrieval info: 	<generic name="AUTO_REGISTER_CLOCK_CLOCK_RATE" value="-1" />
// Retrieval info: </instance>
// IPFS_FILES : audio_embed_top.vo
// RELATED_FILES: audio_embed_top.v, audio_embed_cs_insert.v, audio_embed_frame_seq.v, audio_embed_sine_clock.v, audio_embed_sine_gen.v, audio_embed_sine_lut.v, audio_embed_sine_ram.v, audio_embed_input_fifo.v, audio_embed_hd_packet.v, audio_embed_sd_packet.v, audio_embed_hd_control_packet.v, audio_embed_video_input.v, audio_embed_core.v, audio_embed_registers.v, altera_reset_synchronizer.v, audio_embed.v, cao_fifo.v, cao_merge.v, cao_avalon.v
