// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
kVfDwDKUrKEJ5BGHH0dyrgrpq4OHSceUEJq++RPqZT65yVlYaoIQ168xru+sD/LmMg8fpFvdq6C2
+6Pka89artAqul3ZHEYsFws+lPTL5aIGovM1dLWrF9Nsi/eHPmQaPSOKbHn0piESjC74dNHolpRz
KlNWh4ZZNTWDU3Ke4tAoirXBkuC/q5NiAU8VEbAJW8boVzR/KnUk0lY56427HlTq+qCVm5utqHhL
Yug9tmmT3QMawrWJ+GAoposFHx2YElVUr9WnzeA/lIN+k4H/QNOrLflOfqpE5wZ2m7WOUeE5ByVL
tjt6RxRlXIuzPZj+EQrHO2zUxgBYchMmPylDjA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
zHh+gCMNG8hy4ohL/sDQqVX+4rML83IqRT0FoLyBa/3+vsXhmCzFbkPrVfwNlu1TH7qM5at6dVS8
vYnpeo4V0xnVMqjNm0f0uI/8/5/GWKNyIEDGhqZ+cJ66CvOcKKdNTscEGikfFuP/ftM335rVw4zc
QZbSurWTNAsfybRCI+b4iZLK2nqtyZZ3hWFiRcIT5TO/XnlPnPddLb3QkZcfymYieQPOIEcrBHjd
rrCUF/8nogtiEKcOxcWwYXfjVJH+h+2BY6Vdd1GRhMEqKP09e18sHst7rmsjmwdUeLt0dfxiDNE+
+RCOfzCVMV5cadvVRaXYlRdffFgZgCFYaRvq3h4RiBJObIKKZ2gKpKOe4vAXTKtXlNcccNtetEMB
VKZn89yeIpeDc/g0LrL4kOp4+ldQAkVCuBVXXmDq46hBaRBv1BRwlwt5Hhw0TF47hnY78AJFrWZC
E5K4rZfLpChpGkULDxEOnQuqs2l6PuVB/7RgktkUx0W/woa89o5ol9DIAGfLSd7MJBpPzUMgFQrk
wibo2gG+vkAMAj94fdQcgJkZaldqn+jm8Xepydt/4TP2e25WV9CWyRDi1YW0GjMXAGeKNZphRlKt
Mtj/qlZ8ZykIJ73VtuasB/znrldUjv8o+1XJ9+3YCXRdE0R02E8e0HAazrTjIrbUp7JYamBvOqwq
3VC4ohPRqdJ1JG9NCnX3741cxr0C5xwldtwOB/ycokRSE5U9wUqiqwpDR7PeJLVMTg9XTgQcSXKG
RVIbpoQGiY6NneVsyNuB1M54KREnu3B04MhamJb6hIXm/Brx46gX8Fwe/BwRKvP3Sa8UvyGA5h8q
TEbbSyVQYNstphIGnz8Ad66VfbV9HtMLnVG2mrv1arifVo3Rsnw2NH/iapHOWnvRc8xKqIo3MEDO
WVlGkIcv2Sy1QfZO7WrQoRZ6OV510uy6pvf+yO0erscUN2tI+vWI7pO+7Kk8cqCwSc/VDDjdZPCe
lJ9Rrxnhj6fzT5Qtb+ACSj1QVqABrJWL73j2fhqfTveGBUAfkqviq0hLGFyM4KMDUKkfL5EGiVAM
eIhtjE4lfoM90f3yvkS8M2SsJO2yhpFM9KvPanHkGAxkutoPolPFFWteYJMa1ocJDQu5pO6CEUD1
0w0unz+OxrOqWUshCOeqVIBilAjfLwHeCL47KL7BIUeVYpiJJvIYnckyUwFwppfjcXPmIZMpLgXn
x6A0T+NXtfJC0Bf95ioGtMe4WkxCKU1DQq/xQsCh562m5VABgr6/h6HxxKnvY/eVEk1JEn6gF+jU
iFZt6nOwvhvU+wJWq1eJLzG0YicXAYE/K8ONFzAx7z3Qm7F9Ou9gQyacBckDFNzvuptG02Ewfd6e
iWu4KlWeCpaEMPMlQcH6jSQxRM9hLZvR+tqEaSPRAPN/rZUFAi/XMhnfbXGf91hF5O+bIJlnvuYh
CrfjcrAFxILow89XztCIILfrmFz0qlMJ5TJW6o218TbuKAJn4bQ2/0A0Yv39SNtAvMThCN0mAcyk
H3IOGpM4CVva8Wgn3U6f5lMievBl0caYu1ao7Ds1P2vnR7WH2KQ4WBfbrbOCCBmCb7Grj23Uk6/j
J0RGER0CwQtYfE+GunokEWUbDQka0SwkuefEIfDm7nVRI8OlZKWOzflMjHqwTnI8Y0ZISCcH6MxV
wkr+LhXkIZXprwdvkQG0OzvoMlMfu1geSbl8xc9VIvvdBW90Yaxp17dveTIXCeC5cMT6CflboKe5
LtKbDFF4Kqjt9p1A3QbRxtOUiKkFeOQDqzurOXdB0wKwFHVtFgQfMPKVNlYWcrwQ//31ast0vzdy
U7iTdqVmppwGJixomHXSu3ZwxbVkbCkICqnx3ZT4Hhlwm/T+iHln0/MDSmlrmot0vq9kIw7Qrao4
tLwF5nIb6AihdpqLv0WIfVlXrHo8mR162Fr0rSNPzGR4NO3Ov3luqzU8671x7PaRPbtW1fuPnd/e
PWxqo57YsxkKcqXy1CuwfZZR+f7FSOwf2VwPOaUcPcdY8ZeaDj1VT8F3GDMUpkWuyi8BYkGYJ/sa
aIxlugK7+3Nuz3RTmJ84fiZ+b50ivT4XKxY6XMprhYjXEL5v2D/5kI9wNIgZzSdFC2hI/sEC8BnO
6qA+V65CYri6dzEoVduZuzVNGoi8dmEIHeowi3eETyod1bjc+qcBBHzfX+47XhOVXLjTSEfsT1Y/
A9TD8J7wwm0Tt4UTgtN8JDx0xe07WGjliNB8T6PwElilmwAqP5eFL7ZsZTY1cT86BnxwRxkAt5XR
CQrH/okbYsmpV1h/TYUrKIDwsASikCcT6OsJamb5XHSADC98AJDV2mLL2s/4OhhMGKbwnvR+EgxI
ueFiMnXiOeFdGbiNay266jPV2GM5Fqu3fAuSbOn7oAFG9NblphHLwYjHStqpZHVTw/+BT3YTwn8F
deAAbkVll01CnPoyL8QMTP9be32pQHEVKavVXQKS0u2ON6//4Ljl1ZZgbAKV1xNiuhu5SIeuf60M
vwGcslgOIEfpsL2t9kIDxN+OyDoVx4oyXS8FmP6dNSVEtV6GPllspMHT0wzKCaejT0I1T75ahJa5
D2N9MjPQYsaHHWkYxAxwkj3+JPHJ15X1Axl6vBVTkCJNw6Jsl7acsfOy14mM9+L9+RnIKh7r5/GE
xntWuAxpPJgOPfT1Gbu4nA6LSaDLmLpnRcYnpLy7a5mHjdqUOgZ5pamtu+/G4afDwPy9kE+yeoiN
NeTbmnnMVjCgxfUkasXjyx6kaZzE/u8D+7Z1Gi4OSHKFxNcWuaJf0EB6BgrKAmUgGelmkwR1n1NF
q3Pyxu16qRxg8KESK5VHkSLFYTzJ/mgfWDFRi2CSG34jonISJfvdP2SIPYEGIaP6M36HQtRXK6+1
xYz5TG8KhSG5pUTZ4sPHypoBhjIHVcKo9UJ85hc8FH8zUZ2+Yf39L/+VJB86wRNnQRxYnR4q83lX
hlbqIQ0VmnA/fBQH1UemEYkjxgk4nPjOws5mrc3byV41UlxSkFuqkfeCl8sETsaIUao8jBieyepM
dGFDl5btgpcz41eqblx5dXylyAVbrNNx0tur9jvgGZOWhOZZNFKO4KA/2vpoJPDCarEF1M6d6bK2
3iOGG+rH6CsPD7mnzwh/x9NlrBw+3Egkx3alSssyP/TBZVs+U3b5BunrQydo1dQ2YfEKE8U28kBD
0fyM1Sx82PflXoZtzvo3RgFc5mQIk4+guhctwDBQeSSsWh4PmAs43dlnaMLCb/23voBFNagdOqQd
a5iu9QueanfuWdxwoUVxWGZ2WpL7WOyHNLi7xdqgQDARsXG629r5AROPbXYCLaAGeGiflMZRur29
aAf/JZi1+WjFLipX2vYWh7iScRSwuPMovcyyfAqtcxyzIu3djUQZUf1uAf5u3HzyTw4bchJE2MJ4
uU1udvtgdXc2++vHoIdrhNtk4xjgDXJDyTR94ZPSHgX0PSC2XBh60/AfRDA41GlZ5m93lAI24NlW
WL1lnJR/hPAjap3gXaqrkORHfWulxCfVBq6IkSxlCQs/6q5znIKpePC2SNnQUZNFqa9p3LvQgivR
2yklai4hsXQJpE7H3Lgx15rwc3HKWDktRlEzWXzd6yMgMZUV0CrE5tBJygUxmQiKbVSuIC2CCqYO
oc0g7lQfvyLWkzGXzPGO7bIA1LBhD//120cEApSRRp7i5RxwCGJj06pgA/SePMjfIAr6VAP7ONSQ
YjyPKxcks3L41OopGKrokQAYjqxaIVuiZ6tONCP/mCSirXhRBu7ZxsU12zYQCuzTsZl9K5ijBpMm
AMwB1BrFvR5v+U08nyU7wYhf/Y6ljJ0bNL+oJWrBaDTxRtfWbJeewDCiqVNxbjversLfzUIChG0s
LBS8x7uvlZHHRlYRwv7MBMcFSmWx5OueeXNTNU9pttz/iRUxPYFZzGJcasaw0tzvZ9KPeqZxqPVl
yR89pvIiA4SBhkMRhhjRGFuaHnsUy/j3SQ2rCFCHSHJiUD798nB6nFY7uJqSGN6yf9GlfjhA1dwt
m591t3sXDxWQXHUzxHvk1o3IQ2mITFStFIyNO6QPiyjQMHS0v58TptwuiO2bTqvMrI5B0sNYHJSM
tN1JseB/lnbQauCcfyzd8wTdM7GOlRi2Kcc2Fg2bt8m+XYHqr4YD4TklxOdQo93ZGVB2xcyUcNu2
EW5L6unVgECd+eqQqfXC5cE+8CbBKxJ6xhgDXHNicjbjcjhjw9CEOSbBI3asRil8r9Ga3tZkyRJ5
i2AQzIQTCN1CX0UaMOeT4XPzSg+zpkq1bPFREcqjSWOodmCPSxwxDwSDLMgjN5a5vjgsLgEOCqhV
oWxfqKN7YvjqS/2986FAwLiUAvjXO+pQqOWs8Ws9Reh0RTOSjltpKvXHRXRSPIMRRDdNbhLI9e5p
XOTTxhBQJqTxkcT9PPxwncLLyfGkskNZfP+juSUOI0efeX0QBiSg+OTy6vDblFXCE7+22kOSk6FU
b7k50LGL/fh/HNyHETAN7Yv3/pJPquxWd+NQAqamR6rTVoaHuCsD55vj2lnMsiNqUBmJKd6Z81ba
0FJjB1sYNf8REy3hBPf/ND6VvzO3tMy+gap/QllmtVfwVDuAEiDLWhpMat+ggXiXUphoqrk2hR+d
EjFx30PhAMXc4zXTY+ZQOn3XNPARWxK/uGOvxTLnsTQ+C/6pJMpiwfPLIq+e2Z3JwkQN2tLVP2DC
YqEtMtyHl5IrwTxk7bqWcYtP26vJK+4xI4+pNhwssBg+bR/RG4b0iSfXROlW6DyypvU607XPBoiG
tcRCaPVe3DlnhSfphVK0pOPYbB578dZHVRod6U0nWw06J5pGrtrPr1cBjTU7FfSWVV6erwss92dz
XzonmhaBEHyZUcvLmzJpwrpzyZ3wPClsvOsMIs9t7g8ubHL4w6P2XoljbTD7g3YsTLeSndAXfSyl
13XZWPPQgfTHImGiIO9JeFjXkhYh98OS3IL+tZFlwNT2D8OeF+DZch1DLDFo/2vCinNnbmogjBLj
pNUWrCkriB1ZHHH++UKvDaPHFCQWxdyzCIQpZnQd3WvAfo7FaoPFvGymQFcXtbRbsEWmsZUkutk9
L1UiWcczYVzQ1Lud13n066E9zxmwMlmVbEG002U3AQTaV8oKjwFpqaufGFPbJhftgU9O6pZZH0yx
A58Iwl7dnYXXlEEA31zTkIIhseNqsMdYA/RIhe9ulUG7e0Kd0M+uW8vX5zMBWSeK6eLNknNqSl8P
kqWxQb8GG1cvPDambr6xYkMlmKv+WNniBrECaMMI6gpK4REyCkQufouIVNBl6vYGrCtOGQXVplLw
yhu266ToYwYWEb/E0pl+AmgQEfpKSrMyfs76zV16F0zmEInJJnlluES1x1B8xwjPp2yLHAOthtNG
+TfbAb1dKaAeo1yErQZLQd+MRxRmwg99PLmxYT1RBRCHPeNbJsX0TolPLTjWhXuoDZy6UlgXfy/C
JDbB0uq7LcGgyiCUQPviAP6O73zVY2O1GtmR2TYt0y+ZAm90CsaF9gXTFC9lWKiMJx7sj61B0uMO
/KAlTfSotFq56Xhl6hmWWtxY+7/w5/L5rxqsHtk9Ac/BxHyGRuJ9KqmVjZgbsFXrjRzwzvc4hZxu
16GY+cYbU3NXU1QTsLRCyO2b6w1ZzKivWJ1vwXMQbFVlIWV4oxpl5laFKb08NQEE6IHHwrIFrMMy
bt35zPxOWZWHxZPJlUCedCh6kpmzuXYY4taRcHfkLztqIeljjmWHOMxv6m1/6w6P94Xcn9mBUgpS
7jvpYN65ldZlirB2F4qEAg3bnCQJcQRwnwLzRVt/pxsupCH1Wa/MyKUOL81GCZtzZ52mTcDPmaiB
yQvtkZ6VcctTeSqQoTSxYJN5kQ/Wb5jnSrzQrBLsGoqpswxefqi8a8XM9X4sJlqyRkIF2DvI2dCe
2B4ZWTl0WXUEnJSUF/Hzyi1ATjNvdtmV6qkXRUFmEINoLCPi+yQDn79961OsaZ8siEOooP/Hacww
bl8mJ+hxxjgBoGQSBYoSkKsMCoNETzyszHS2CcbrXwQkVxncLlP3VlPQ2O7/6htgdEmvqV66ml+z
hv5iTaj8J0joQS6WKWWu8+bziq56cP5LGRl9LjDVp64kiR7LWCe/3zA4DIzzOL/L9Q5T671WkctT
pWl6gly14SAnkwcVtRBwUfGNd3DOAtn1uSyY5rknS8FunRYIyopMTlygq/u5T+FYLxUIyd8Vnpx7
nLFn12VNuQLyEY0G8zj9CUZ4AJDZHbLX790MCOgWgn7iBxTTCCAtE/WjLXbmGPRNrFy8frQD3nyN
Md+gVSVIqjTAH/qqwFvohSFkZlZKpgoFTl02/hFvmHrn93GFqJXQRS4iGACPXhAAe3bL0g7ESmuA
0P+8k6ZHGpILHDdcdIPUi1oOYF4JM2kQnHUrW+PtuGnlJiLA8ANyE4xmLzgIejAfIEBlnzpdg3No
zyhQ5CW3aQ2+DQJNWwOlEqGIcsLO3Nt7O6TRUnJbYC3Vif6HH7hnez7SlLwTFxSLG6dgEi3qgwzL
ELuXyhacJbqql/PjBhP5G/Jp3U5bfbiZ8kVOEAHKyyGzYOKDFTRdfjfmIEqP2hVP839PtrhST3Jd
+0Itwdi6OF+r2TqnkvyPfnZlrcePAIU+JhwycKzIwUDnP4s+XzHsqoK0vezLSGQ1Dln8gwxnkRFt
iZXqhUI6eyYvcyP/fya6oM2aqrCFO+NvrM6TBMQCnMhm7MxamSrTyMr/nMoPIVSwyg+9VMLYClVL
kzHP7B5ajfdzFnx1hu8+IZN1AAOLRzIBOVjEVELfSKuDJv6QBOCYJ6rUQgoi2V9Dkzpnxne5iLvf
1ej4AydbQ8cXAgVc50UOHJyhdh+un/ikUvJHMXM7LvnmoBMOWIpOfz1Zl6p3GkrV6zZPCxISUZJq
24wOD/OZN2IgbCJuj+M+fO8zmtiNApzCZ0f5ind/HzVrde/3RuIIu24x0Lz/PPN1JDEyDviugnpG
Q33nbQwog2vrju6gJitw+7A8CfFIT3tNkmrNeQs09DYV4W3OaZL+on/CX2cyzoOotNMET5o4XYP1
40yr4UHSlNuZpJsT4UD86MevEUBpux0BpRsabiF6k3nL76TvgEK3D+qDo6G7oBZPrQVm5KRhTUYJ
sEC9yLbW7wIewt9l+mYa5fYhm09dn6BWoDNW1+qHEEaT/nPzaApvfmsVEQXU5OKkl6MU6ijz+JIa
7yg+o6kPnOncrOLO1dRqjywES/hFo/nB1451W6UsNk4XtCniA7jd20Gl70ZHeZlWFlTBCKXgeyRA
Ceo6Hh1V7+umH9tYPI2hmaCa2EsRc7lokro8KzMStsHWR0WlM01LTPy7UdsgX9Zq5oxfvKsz48pV
f3FARnRWYntD8qZvqUGyYpmn1qPPXsjdGSnRiM1qvXD3yXGw3oiw99j7nSqpDaRKE9GWXnVI4V66
66hXm1OGCE4x7vNNrPSoXW4kIIEcfj0HaCMAiibQ7kPaBeMMJc+2qL54kHXwdKWFUC72dtLQwmVX
F/7yM5BEcKgV+6JWOlJYsMksQkRpqbo3t3ht6dJaBQ2yQ3wZc4tIWFFP8J/R+Cj1nXU4mQ/BKZYz
Jtn1fuXwXgXJENq9mWCKaZNUBxmJsYVqAfYlLguJFCBkjI55Nikk80IaSJY/HEUvpf/i3lfgL5Tx
5ldypGDdUG0zpkhwG66qxwTxBt6PyY0VIc8IdifI1+SYupXw6+rHOLtucliZhvnz+NSrWzyK2bEs
lVN9ggVsmQdVNU8x43g9Yt6pfQD//qHBPe3K2m5IypnwtUzoavJbyPnrqtuorn3QA5tEoqiDmh9D
oBnLJlQczwPfTE9Fw3Tr+8Q6MXiPwCgDesbyHKxocG+46y3nB0BasrNp2EGXnMi1FskJSwkeot5Y
yYCTYsh3w4QBOobRTmtcsu8NSWZn1CT1al6kT/xxZnPu849h9f9SFRxNnlODwNs8M7OrxEo5pZro
j+VsoaCl+35ll+0lEVnq+SfJzDn4NKPeYMYEpn7lHl0pfN9lME5q9C65xGgOwlR7yuQANxkt4fyc
S3zpzjEFjsUeXs3K/95bX1hScw9G6bypFXXD52bItSzMEZrbHNRqI+eRIL/ZnYifX00Lken0tpjU
x4H+nsJuN1WjfiAFCjB9qWqSZUlFKf0U7hNXkyjxvx3yslCatVhh+gDQxJJ3woTvthbhpa4KQyZ2
aYfKhGF6whFtN0YZuqX3oiimk5bIVyM/FF/kVN1IXLNp8M0m2T+kEhcAbjbvZnFjhc2p86pWhLoM
/RkY8OIM1vWF73ZuyqzXJAG2ULVetZFMWS3x9+j6YxkiZ5CHhQtWnFqnfGBr9pvEMaXjMvi/g/IL
Zu27Wb9RBUtjrWc8VpEWRXY19Rp7Lk9AplEMGSqo4/t5ShztXl+1i+DdyvERYQ82AZyORMVa7ndn
IBbKi6eYwOFMK5uFO2EmKV6DZw0b/V4JFe+ZrquFzKXOVQVZPl+YHOh0dhBiEzP+1wqF5XG3imKZ
CdvWYUGYmvD23cRyeeJ3zUhxbTT692cfLXFwQa2rrCLhGBVGqaaT9fOUJgbDadvV4Zq4Qz9gMKLq
aLYhiWRdhphTJVaEvs4DC0SRKjvoaOzSnVP5nauffH9bJw36yFgrc4CrlcWuWaZubvvdTzzeDH9c
IGCcLbhTgdEp8TeHp661POI+gpUPo+NVj3bwT+Bvrco4JFO8/E0NA5dYOqEBIyMEZKsHD5eJmg2i
CXfBdjOd23XzOtyyJufi077e4ZuiJ315oOo4jNrkhr8ykHSY2E75tXUElk6uoJvrizhR0YGhRXI6
aU6d4RyYvdgq9B+iYgfZBo+tuRKnKSU5PtvxWqc4VUrlw3WsevySFPzlYrK30sYig2hyjIU8HvUt
Mw/W4EP56LxZtTK2KYWKMRi7zh5GuaUNndLzFHJyMK2lFwSa8Nh1AzsTL5iwlXenYHf+nsPKNIBD
X1jI0MMhMB8Cn8Pem0z/8SrhBbxMv1eg4htufiGrd/OZc3n0SNI/A5VVPQ0WTVHVrATr7tYyorvW
VacE3l5XDhK5MnhWQANi45LCWgR+elVJapPXeLoZUhTihM1rHvtoyvU6KxJqP4JDxH3cuMGDAQ8q
RHnTe3kdjelt/MHomBaSQX4XQX6gv06/ncPrrQMwdRv7Ag6vH5S9EYMrvHIvT70t2RUmEkeHh1/9
vN81h9oVWJSPG2BFeiRdcm9qhaEbJ1JttVgyQZ9Yp2sc9BYmjqRRxQ0kL4SY03TUk35q96PTiAsd
rQRDswJyYGRkUCpKI8mVhePYei+3xrFub1l3dQeyydECaTpn6QYC2uze6yHvkbIan7AnCuo9cYcm
vmHY3paC4N4MjED4SCsn+Dsp1lCVroB4uYDh/vTQZnPDvNMf1PmMos2I4rTMOa/Bbm8i83EuOn6A
KTVCExaSTijEykI4VuDw+Mt4YzGpvbcR0K7xK9hLfDDoFWrw4i/hwomyYoYCv5e/ZYu0b0unD0Tq
mkmPWk182FDei5yWXjxK/fcewPqcbF3xFc1TMO09qGhBYMdx8+23jTikeUGNtEgz0fc9lCHkb3yE
sX7d3WyzG6NZiN6UyN8Obs94YT493WhZW9WD6yV3NTzbhjkmPLrbygR7/xFgVMfW1L6YF+/oMogM
7dJuWchaATSaEiTne8fHjMM2xxIHUdKaptmIJZ3Ir3HCBYrCek2KN6jNaU046KY8uV+B7c9/dR9K
IyrqXL1nXYSeJDeyx+AlwtoHYVDBaZCynHyXtACjYaHFsWrSYIcqhLDNukIV1Zs/76luRHFOm5fS
IEBdvtEZ2LTs8DG5swxx7WGM5VvswqAXOTB+B1V4eh9zjW1vCDkhddSuEDW84o+IosmvIUce7BXJ
0uP7zufkSnEYzfHc9NxCGc4ZGdl67Xd4X2c8dmjDJ4+ljvMMokq8LOpCEVKa8Xlao6Eahu1DlJfC
ZsY00jTJqRUR8PPOZNTmFTxqT5Bl6rcOxrH6HBqLpeDf+y9pxvxbtT3wn5rGH5DClnts9msTlyso
DwuSNk4DwYC0D33tHWuSg7Ddke6gqRMFYAkbWU2p4bHCmqb4DtLb8oMbNzNMpDBore0WOrLV5Bnw
VVvLwbIvnlwD/hSPKjHoecXL+ZpNnpbiqR0qJaNOAA9e6/z+L48mHKrcMG2KjvEXwwi44GwV2LKd
lxTA1xHGGPfeetSKWMaSHhG0QZllu8IMCt4H6ODeaJv8VvGSnVWIBMMK6sISwQFghCteVbvgZ5Wp
UpG1uNlfSgHnxawzkppLJfLv5LDD+/ytDIVOfNR0YFVQ5TiC/nub71x7LSwWFgONQO7QoS3UeJGl
fnWQ4JuFTsRw21QCe7Dmg8kzIcEBbIs4LLesuJ69vze5fNTwzvBDfmW6pgm9yhsHykzOkzgD5jux
C/WPSLNd4cWDQKXyZCysHgp4xBbXOLzqJW4i9gFE9XnAki7u4QWeRsU7Iwbj1QkhbbH+2+ZtwuBr
t5QZ1qcmEdxLWp0z7cMTcEoINpaGwy1Ce8LtNnFPvDkuDJjLgq3q2R/kVm9I07r2i/2wVF3X2LN8
oo4UI7PFWrc3/6dxpXvyGjv7Y5YX4/E0nRksyDkHl5siss2YBZFboXrXUs5OVXVmAKm8owGGbOfu
+ShWqSHuOP0YR0h+UErB29guVFbYFjoAndnny/9eq0fD5DJPyN4VMDwby4rDHpHOZBGJqki6pQCy
dIp3CgzxudyzivLNYkNJzIt+6BGFgiZYXqleptYy/lgAfwIhtJ1fXJhglez0sv4zqGsK1ak9Xskr
qYQ78W6li2L1tRSLmaEGi/aRkej6Uj9FS2BUu80qPFIO0vaUOjYdH3JlQsxAQEyoff+WFoae5hZ4
tr6KDPSmJb2nW9I+Uh4dsxEWmuk4vHfIxYZmlykpNu36r/9Q17eM6akWuDK+02O0orfyT6HuGZ4t
AJROwgUkIz1XQrfm+2k3EUpon4PI1VSGqfwcmKQd5mthYTsAEvd7bzCr+ZlWA8Fr42ufzvj8IT2r
Dy00ml7WorYdY8p+ZWeiyBQwvkvsBPgtO27ohxs3fKEs6kxXeLl4XOJqFey5mnDqVkrcUqeI0RLX
4B0bHqO5qXQ+8TJcjjXi22lXXIumh5bejSPOtNnnzi+wOwatBhQ8VEgg3mD349kI6AToyS+E1C45
Lc8TYu1fi4EpBcRk30U2Op1hhanXVELgskbHQiaQkgyw9ae8n4oQfOw7PThntB0OrHNxFzqNbHNu
xJIrJKO0cgB1wzHjTeZnuOqItRt6vawJjdlno+fpXDZ5IcFxg7QkQ0b/y5iGDAimJ44c/ttwLV8s
egkZKVphOkXs70mUOJiW5VaYXYYR0NTqgU82q7vIVBChLjF3CbM7yMuQWrhZgVONljt5nWIVo1jK
SZvnPfS9HUru4s8GoJsvX3n7Sanr7FPf359WH5mOnpF2LChvy0P6Qlkr62GUKxEdjLTYI+xfEFyK
nGbVsj42X3mcQkjQrBYGn7GmCIo1QPVvSAxZgmSN2ZLGTQuz1ZXqJ3qrKbGLa5K0E0NK3KzL68nb
BCEqXyEm8v2Hcln+IS55XPqi/mpSWNgpzF2i3zBo71m2ghGB/DgjJIiWuvIpPj3CSHQvWU3OMo6U
rnAVK6awJ/+yxz6ZvCyebbnvOoWlIoPjY+a92L/NIB5syx/5Jsb67Z6TtLzphoeFq0gi56K6S083
PIOjIfwzemL9BSQAjVUZlqHEfyvmo+8HsuNBD7ztT/LlkPLleSg5/si8biKpb5Y4JwtFmEnVrLxW
FufU6heuwBDidnWa5XQn3c2i7J01qzUtgBlL6AW9QOzR5gRkiXc13AdtYnOQhqLm161ar2h++7fb
3kHw95nKCOse+GfbR2AeCmWR/uUgewF3MsUQWHyOreQUfaZVSWQm07NoAxcvpkAfjD+/C73b+tJP
jGJEWdgay91cAsGnPBDVSiW0z61kD5UImZCZGlBCw5pzJCJXhd9BdkZ+nK+RZn7t9xEhGOgixY6U
J2yZ5XFtimjTGN1fu7t7ntJn8AYbfqyKGLEmM+ziFcKEEoP6+LWsP8/NePekU+Xl71x/uDX8fAXm
hdt30p/RXJtchAJPjVb3Aiise3axebVfotBoBCOwaNRHEnJi0kFQLg3JVDWltBSJXTpI3R5HH0C4
2XyXhvcrhWtHaGMHi+pQ5nJx8TK5t5pWqX8jP0TCb4uMYnpDHW/uFKif9A65gdrEjCKH316FTNvN
eJf2ywj4B3o0fjaZhV0s1vH2XUcsf7ErfQWagrGEiEKyDxIoBjgXthbmEGAVNLg2RWlmTBZRvdNy
GFx49Ny3FLFSB8Nd2t1z7rWPztmoQEeVWYzrd5IWTTpI5huWaXw9iaelFghj76iB+VAHxrvkXXxA
eOKAJE3ArESXitxLvP1HifExpOe+5wtKrQMqdgsP5u6lkpDpRpzc7aMbXc08BUlbsqP7u+FLjVAa
8as8uKdKPap4JFWEFp+uiCw+mePO+c/+P521xX6odd2KnWadrvWb5jVgd0++LYx5NHyyuH6kyOS3
OAiRsMakw+6Jk6FVcheSa28nuWSweJ9zfTnNjdyZoq69/VFFqLSXicKaydXTapdLg0jPMoO+gW9o
do0geRqkBwyVrZT6BTVW1gYALBW3pP2nSsNOsSkWNOE5wdwJcUxWzjzksk+7Qr96UZErb/qbbC9a
Clz+quN1KbMcxo+bGdrpGJkMsP2negv/kuvRsEsSJgDmX7+shr/z71+ritb0e1RLgQkpjmw0fcWV
8sDXB7mVkl/pZiHJxypSEpwYhPAMbzArYhxXxjDQI8E4BhrIw2oKjkdeyt54hm+j966WjuWL63bY
mxm1hCYSKcPlZETeezRfwpb9aZtDa6dbMvzNQhnCrvF4Y9+vy8Bu/yFCZjGJ1vPW60xjo7zjc25p
dRFzoRKhVdgVVg9ThllAQlXRaZGEnRki8SLXhufq0s4ENmy54fgh4/rJZGjoc7Jt1X4deIR3gEUP
ERZwcvU2xMoDiKl8JfaBTFPfuYvZ5tm74kuYu/5z/E7a+f94SbTherCF4ywYkTtWFkcl/DdRe6Qp
uhu0JW2d1j6F90d81UFcr5hVJu1Lpl0Y5d5wuYZcXuNcF0KCAxqc/fw19fIJpwDbxBKwVFbISIPV
m/Lgm3zB99COws2Wzl3YRSPrwoLc/lBTBFfWd4NjKoJlMf5xqkXTk4Q3q1KUnrGNJ+S4HP5cT0CZ
eobAGem3JbWErp8kC9lwRFMXMxg2+Z6nWw5UxR10ghSAXNPVNrdbeyzJH4EMGfm46qY++xMi0nLx
8IOKPEhjfRKuyODZXDSLHE4OhZUcJBQ1663H8vaEm4OXKFOw1X4m5Ok7fD1UfhGopTPoOelPPLFn
XLS6pctxdcT4AfpShPp1MpWaLChzr/+MP8WPXrihT0gQENkNuRUuZezczFZkkfykxjOguftbHT0y
cvjAu1WYqWPjNmXL8vyoCp4t5bTBFfNkbnGY4dSkxnAIx2yL8pY7/mEo/lvg2GUqqolvw+9RebpM
YCXuiDDt5tAh3ptkEYZ9yVvtEwmOwwPtGPWy2fauX822jNO/MC6NNA4Mv6XIrabBw5K5gZa+FG+t
5dOYBNb8iBVbKv/mPKNQyGtxdrpftbhldpRgOa0ZLC3QwWXRiv9RZtcsOqUN6Iv2qAlotB6MsTDy
Dg01heSae/wBYQNwwhRpiuf5S5An9hPw+mGRBJOh/kkicLvByyqBtvJyD2yolvn8XmKmDMQYmfpb
6I+P1FGqxrR7QibHy+RLzcRZHTZ3YvZ9X9rHIaWS8Jq6X9T5aeStlnZzpXIAy37SGcJN+EtQQ4qL
rckK4pYrR8iogzVAyjGUV4yY544gfAm7Wujhjqszpu5iAMGXxfQLf7BQX0ZZNK/o6ByCO6uAQXfX
mncxoN82sbFyi5FsOsDopkaq0Xt3KTuMyjQFA6MuGKA8b7Z1HvDB7NJAjTxWftcCTRaP4KWuGe5A
ZW4pMxeHkGr7fhX67dvh80DS1qxZLSbABMK4pMoUi7NMzqQOY6KlEFAq3HB76Aw8jbCI6gQDZhR0
sqZ7a6V0PMkyWrVd6at2sPJZyEkDMDX7bqTiZORSOEjCgNwnIC4ppkmssCGC6GcFJ1iC8EJfB+If
BZZlro4OvQAbdMsWoiAqqMC8rVnnqQylNXlNq2RlS6P7QLnHUQWAkux/HH7QMAJIVrCgrxN41Utn
imBqqgZjyN5w91nacJGlYri3U27fzRrtsFnpKdjR48chjaF1ev9uCXPUTGY5K+hhg8yM1jHzbqbL
mwiFXh37ZpKtKj2aldbyl9WFAmLLFE+pvh1AqakbhAXd5xuN0/sMpaT9JYGWIbFuTAz1Ktm3mIp5
V1WgNcbXhU0DdpPhLLbj7EBL03iTTzu112RDSXaUW9OqUtnhH0Pq2YBmDXg/JHAk8qbR1PydyagE
g4SZ4JKNYz4Raj0+DnXCPPbRr/vpUZJ33NPscjO7HAf63YnFLYTeSdlWgsNIfKIIYh9utIsXx9W8
wEtm6s8fTuKuGtoP8OMPAB8zsi/yUU3MsIFpQQodv/OFfdryXxtdfGVf2YmUecDuEIcwD06t1Daq
GPIqhFNCZLZhMw6sLE5djVgh3B0hu7tju5YbpXlkgYNA+I7YpzRZOs8a3K+jzFxJ/K/sMhtWkfAv
VYLDFX7ftI9Zft+6+N5i6+C84P9CQYApnOOFI6JmWVSPYC0dljJqc5vYYImBcUtG8HLxJyyvbOvK
UKTGD6A2zKOLrT/valTb5mU7SxvHQoPdGQSIknpTizi/+2ND1VHeOGC6a7YE2bXWCHOj4TXKuG3X
wQjf9/UsLg6TIYXU6xJ0cdVl5AkaUToDfHtza21IyamPNIfycEzvnZZbeexubvR6/tZdIiw9bhM0
6nE7vfDWoTnMIRPaSK/4QNV7sawTYzG19GvbQc12TteJZSVtLOfEcDJwqYqQIG/ibwIPMfC3I+EE
CJvutFKZnAP2mfWEnXZxFLeiEL/Smsl2P53SfYHYLpLa8y/zne3QW9Y7pcXJZc3BSm86xOFlfQEZ
WV82PjiOQUsJZRoXDuky10wdk72Y9++3NIepllALpmLYqn0eiPgEOINRHohVLyPoqrZYslrn2ooz
ssdmrjo2l+g93yl9pt6yh9EWs5We5VPt6nEG+R7jzsx+qqMxkO/CENqlKHwU/LKdRzbNXYe4dJOd
D/f7+2LD1P2pesCY/eFxTiBZJ0T3oA+d9/y8FrpixbTD3q7BpMzQo7K4Z6By/bytFXu4nTrOOOQt
XxSqYfAZ8ls9jnbPHcpBTbGqoh24SXD5VDOnuDTYsn802rxpVsnLThGawiimDjTwKCgq90W3FBzV
aZZ7DNTPxgC9IQMaVk/558EyO1lz8xGzkLBNDf0/wYl+zfxrVLZOuiP2y9caPHN9fYIWpfzpD/0c
5IE15tghIkYgemkGoLGBLEJJ/pMWrEYHa58i90IV4013UFeSDQPVtO2WbPh2X8Jpc5TQuG1/buSk
gijsZI7i7KQt4jo+3w0OtDH3BlgJaEawg5VjnFdzR/puOTgeoPcemCCb/rSCz6BDj8+SAi6hZdgO
ow6tZCbEoKWgcS++eiTqSZnnMo4x5Fzrhghx8CT7DVe0uIn5j1GmLgM3jbli3xAbWCvSHToCREOg
hCcsYRBRQZjE7TNMuRqcXBq8oxuZ7iglJB3UH2pNXxjN2bFsmMQNZCD8F5mwqFFypjBXTSkJdfiY
piT+Nu/a0Rwsv9fRjDTZmSg5ezb3JRjEqliYlio0s31uGdUozoZu16gyAgqFoR1D1XBivHkCpuNH
0i51y8DVggVDmBYonr9IYxTf+FrZiZz/FEl1es0GzYRdO2SIp7DRqvBHgJOPlxi/xFKDi5PxiF+F
jnQdYulXP5wqc0ZF09VkEHA/RgykigIiCui/mhJmw0f5JcxRNJVB78TGnJbm97itAcWdOF+puU1B
+rZNwBhAk2EasuoB2Tc6iiMz5MjB6Vc/liV7pJRNGzNpoal6QPDLgxSxaK6QlmSmWMyRTe1zw51O
rbl/oEMGDeuNOyWXyzv+YCQB3KKsR/He/D/NdK+kdYLLN/Z5YoSUfrlmziLU5amGXy2gFInIZmc5
rs7RNivOfPlfjyEIOhNZPRm/Y5czrRHFqv4ALgw85PS2utQzSC3Fck9IT5qynGY07ksfLnAP7I1g
FLDFkUWVC+rzJnX71Ga/jlZ1Sr6h+T0afbOi4JOYOoh925wV1jJDtWFbm3ctgXPdKO9WgLHD8PaH
9mitR9yyV0CbliGpukMKfRJiYki7Kg2c+ZvD2+oHgeWKRR1ZNAuBz82cZxf7Qc5zgjLFDbjZLe2S
D0ev8M9/4VIcngFv9a9YuyImSZ65TTygXXhqtuDc2s+artFf8mbc6AFaiuMp6eH3PlltJ/OiVbDn
9tvPOoV4Pj6U6cLtrcGa7QAOhtuBal92vKna2iwuyvmgn8nn5bnc8KtgJzndsEOpSdmmcJM6nzAk
H1hlncGThv5hlz9WAub9fW8rTDiHUgBCu002ITpwCI45KSq3cY62ohTPk1VdIv1Qaj4K/SxK1h9y
LZUpNc29+fXstMziKoxQfORZTGYbAZQFB5xujdvJh3xMaEPtwNEBvx2vOgaQSr0b7OxHNp7VLoOI
p4CPQp+4XZjE4s6L+rzk4l3UE56CPiolnSbtsNl7mXuSYYorzNLl6RjGg9Z5P0C4ykdSaik18E3J
qeqjYrjMbWX3zoEEkNTKIFUNzlHNZa19YhIBCVqPFoCamj/d8LsrFqZpWJ9VxOZKIwbnxyj1J5Fd
xSG3ixK2Vhk5qNlev/kw+LfrW7NQ7Bmbx/K1ieNX48qWFcb2RzMv8A+d8FTXiH0KJyUeR7JxxFLE
JmGvRJqGx8cm6iPRwuPWUoDVF/aMXWi5fxQ1SfJMJqSXi7AOBtEpA+mmg759TIavVosRug6NmK2C
Sox2/AiaVdm3PvbcsLHfxjoAWnLZHLi3n92LTWfhLl+ECpwD0/EmHmSdfVOS+yrfUHb0XS6Hf1Jt
igt9Z/340Cw9hP6I+0lY6moRZc0yc6n9ms1tqhcLbt0kCFyL4K8mcogxcoC6+LGVT18/9GebjNn6
aTmYiIeuBY2ysxBEhpxASLS4i9i/Dykr4/68/Q66l4wQcZCKjJ2QZhB0gkIe9T5s8E8o9bJuWbUx
t99YQg58z1P2IPYROjoe+TYSF5b3pR6bpqU4xKBGjvW/vYCi3vJch0RkNoRl2NXvjFASRlzTy/38
rVAPzh03vR1flk8djMJr8USWd9qk7QRHaJQinIzw6SgVDSRTxs/nDa/vmts4PTknLnAbssdMH774
6Dj7vgN3JoVm+EHS6Rv+l5B16vqaQSEOrbRoF6pbS9PAmSuAUhy274LBBDu1gz9wGE1U9uD3EcwT
KZ7KFIKo4jmO2lUPhuiYx5s0p8G44dBeHoFOAM/aw/C/yjEDsddS6XowH/Sb2L3PPmlA66HwKwkR
jPlt7Bk80MVHdPKdSKHPU48qgQ5+AY5yPZwRu8aBTt05hAfItFgYfwWGoIL9a7m60QY/BTrWmjUk
T1JXtROgvIfGqf1sZIvxwuqr2bbpI74D9A6hqNzlCZzD1mOf4p0bsymSpj/uUr95Q/xnjE/N95nj
4ylH2A5vJexFzcag5L+LLKKhAt9m6JUEc9yikPnOjiFpzC1rGUFPJujhaJVx7wXT8ZTZhqACpCQu
dsYuvAvR/fKRZuAK0Dnj86u7vnJpHH49qRaAax8TAcXjnB3eTNl3NToYiGZfztwZlZQz89yk1BM6
5fx5AAE/8rLEJEtsZG6UAE81fLlNkrxLaXRM9fAkLExKPowqn6C5gzAfjPxMl6w5Zak7WZhWEj7z
vrJ3e+S7q/8hEx1Y/R8GIrCP8/IoP2ILuWj8qngUXJSK7BhAm1rRHGeLSsHHdh0C0Rw3NMXWTLAU
TGgvd39TYH0T62wX1OU+PMDDBVjP/t68jb78xCETA1etrF6bHuMOWHJGozao4sHhWAyCT6HBtUJD
iKrPm3rorheAvJewEMcMPJdDiBhPIkM/2FR+rzOfWQn5cKWWuSBV0XdgsDRGmmto66ptuD6uW22n
TkggbhzSdyqn30IKopngb7IEaEn2p0cgK73rzy/p1wi+37EB2FLdaiDL688VTm3mmp4otQDuJWSE
sTsyTk53FEBxDQL7yE1HBBLWmAQ/P5ds+5PDJzRwVAuHM2MUSt2vzqqx5WGrYst2HBTC2wZXZrdp
sQxilrmOjtjCp7NxlDzP41OyH9ZbD7xsdYDVix4lc7yvwLRNgmcZjUBoW6Ssmv+Q1ITAc+SbFNcv
RraM1UYseuc7MqfrmSitzey8VS6mSntc1DKfAdfFg9l8C/uwm1Eyxzn9zadKz6eHZA4GlRad5YpQ
6Ug93Ztv1XyvQkAXGfjHjEayajyNxCyMCiKINn4NX2SDL9O+k7a28dhvasFYSeJLus5Vsk9nYg8/
WAkhVXjw+F1IY8LEAd2puXnbet2CPKs0DlT8FrenQmqMS1vUUGeEKemCVMnfr/iNj2EZ+SPQyLHD
E1b2Cw4pLw2sDjGl3YVQuj9PpICLiqhKT1zRuAV6StHuRbAY5tHjo+jAHSeBYvfdQ9VXQp8itPmg
SMmG2t72mHCD2VGPUuF9U2WU0vw1m+W2zIsU5DRtBJrDtQYilCqWo1ZdyM+8tTVU3aGTb9AeEqht
5V7uAZMQzaLTpSmY6tqJPAb6vZA7aDuSKiCV8BXMqqiaGZRUcTqR6Ai96rzJthilLJkgAj0Dk/BI
/m3bP9OSoHaSkvUIT7iRu8ksBFKPnrSOqlVVavUImaBoVCAGlUeaqKGwLwQt3NGOPG/rgrubAwmp
SRqloY11uOc9dFTmVOQF7JCg5O80Nrk5AruQ1ynu1h2o7cuwKS4oC7lxN+SaztOGnRpDGYzQSl55
hZeKKgXzjSgukgJCz/XmzsmEREyygbIshRRQ0csfhVOGFkpDxNtfrjCNLYdGJplZFRfbziJ2TulM
HQgcQhMyZGSXHYiM5GCnJ2yhR7g1VT4amlrm5kyZxKC+D/UAQccjbAAvHGO10Mx0r0E/v8Ar07uT
ZkefJNiv4nAHBtOMcIr8+EC42WqQ57kFjQLbDs/s2lySzxpHlVCgKV/wGc7rNrMZtDpySEVCIQ9l
gVvlUSjm3ox7+fBcdxpsOMZS26GFnLpPea13VoTvdIsBnwfoFepK/4zDpfIr4aqZ0f97o3j+6JLF
AIQ22irddQFd4WLLsMqpqrRhhNNz7iS2nMORV3rAXqLa8dCBiXuKo6530g3FhvHwl+UCHMiq3r2O
pyuBR0tTOfwUqVnCQctmUrE8ZpfwgrS3jYYaousvDT0HyquVJga0uXJissSL+pSqHrLGbV4bwSdO
1c1/2K+WmoCpOi1O+91CnaIyvQiOmrf8Z3MNQAMJBknprob9PXqjH4QojSlG4pBz0PPPXlPkL9hC
hpZ6RfwdNC8dVR7x5cXZuVCZ6/riJsoq3C85Z/4afAcV//4tggI2MtV+yluPLbYCfhC7maYdBjxb
EnyliyjXpSPm4J6EskDkc/ZcaOeIOh96jFYeHEnqPL8LdFY2KWS2zm3JhgZxP2JpV/GBE3GZe9FV
WEzLQoUMNq6tldSv8eTgd4ldrT6J/5qWWpCRtEYexyCY5XC+F3uT71l5tbNQyJbnlpuMR4ttQISs
fuLb4rZXkd0KaaxSXZUmXUx5U566d/rbJc0h/puGzq83Bwbc7LDK1xW1urNiAqtbBTFOYngjIQlG
ZkJJd1SAU5VfrmomrxeLX5OIWU0ndrTG1oCxheXYhiXQyAXbfzlzUd74h8GpfI/L0+PbGh0Rk3lu
YCVeMC4b7QSDW/KLRpIJ+58OnoQ83yfuEZ5G1H6/aRr/s9eBumIEB74yThMC2/kVbtbv7PrDr8Li
ySm05tdof0WnV54vGxSCZqYXPni6trthFqSec6QDPR/vyj+xeyY6l94nXA82clJEKXR+Xfb3naaA
IQHMsfxkCcEb+3+T4VEDShz3cqzqUHOgHzCjvF0NMp9tmVnK1wesSXJCqdDZiSSAQksf9hIsZNkS
zHIvr8ZcVEzEtQAhqYuyzxYj6XPsomCCj4mJ1wjsq9I7ewRpgZpXKeGQw7y5qrkotoGKI/Wob5tr
Gau6GMlgd8fBJ1MAFh71GILGmaj9Blds9fzI+hTfM4GcwC47DDNntVnw6JuwCkq6m2vmrdwBXNKz
kDK/47TwHbgPDaCbOy13ntKu/3k8+KAHiQE9rJrCiVfabQAHMyLLH87qYewlgOHfuuqrhKcC6J8f
v6uS3TV6ereRWt3TgaJGwEZXZN/YrV06V9UwCe8hPeQArd0VNzcuQYj0eKN/UPxgAfVyowBN0wWs
OAntXCiS4tKCMnUIY7bxtt7rMYmF4WOtspDR4GlltmjDNZ6SkMvwHKQi3ReOHo22gR2kwnzhlF0L
JqZ9n0b/YGcdy49NR+CQiKchfn2d3NQ0HHc7hKl4q70BHojxyvWffaYZfPcUhwQesVlFxxdSkkuH
hkO70gw4JH3ledPA+6yEHrrnmx6lvWSxPTKN2gyYPbxvOMpuVTtAOxbhWYFRY6pw8H5Y54ypib5m
4q81AjYiA6M3RbcOr7nJKoZfMTqLrMkU3gOVUdVi4QcU5Xv40u9E2Xx04FkgjoeCtBOH0FhJN6fN
`pragma protect end_protected
