// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:29 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tK+rdBsmqwmSCppLCSGvu1ilHgqFJWiqCKQ+WlRBi9uxY0WIrap13+BSWDhRWXoY
yeQ3scT+urVm3Ojb3hZop9EmFmJVH88FH91RGzBUgfrobBM9DFFigH9VsPzniO+a
NnYFY19Ne8rptr5yDrIcv1Y5zjg3nJHkr+SpDhYOP4c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5376)
QkpHzmDNCB/fAVOLOmoSpnfKRTAw5gnXTc9IaIM/G0bTVoQ/WXpmG28acKTMM0Yw
dOUmDareGKzM6Z2qUSqGiNDI773sZdMvZBQWBD8Cq1THvKTF1oWPgHkaMQrZ86s9
JiydmkuXbet03SBk9jjauG4rLKtgiVMkFn7KOOt3U0NL0yg7jVhqCKgu7Olugj9y
1zAoY2kFb/+Ow8MUAzEA+FwTMy5Xe1NnbfHeI3eY2d559ae4Z3UYgzX9WYrZQFuN
c0zoC8+jJc/NmNkkC1wzCyezhhcBMAmIGASSmgcm5pW2P8eq2+/y4ZtLwQG/KNME
4znumQ+Z7lTNtFjytfh4d57xlUxv4b1RPG3QEWO0OfiqXpNO3uwJQTsaFFiG9vM4
jKMbvKeOugM+m5T/Qg74PQJf0rxcs/W9bVCz84xsSHg1Rr9r/YseE1PKb13ZekpJ
YxRnJD6cCDGuFaM7fWUSIne+fpT7JcWmSDzdJHpXU/Q8B4Q8/hDwgoloKgTA7Xyr
Xw/JiGS27LJttjoM9iwMxsxs0E8ABix9mCy9wqKBlYE0ohfGoiEMAS4RCA0uU1Lz
zVr2Shd7UlzrAzD+AUNr66Nczvv8RR4u/3mmH1eyYE7DwkP5CYMsxvAX0HIlPP9d
MGYOCjJK5ZIKPdp4oUZyPYfJTjjoBdcDLcIZVufFcckDeMlQjdJO8EYfZC21bvN2
OmhbyJY7kXryAS7QR/JDlUftnrtxZH5YDfqyVKEkllYHjVIdmGx6/n//fMFOe7xD
C3WV7WrYy5OS9E0BUmQDDzl0CIY1jmbmj99QO/YOegnZIrAezbjk0jUB1l8saTZ1
Y943y8gh1//rXdQ1ARAKuuUbnDxuGVrc2VYZUmFgzk3eH966mkuzr3fmUqZN5fWY
H4xvzlJaGBL6l+z95rBMO+yTSZbwGLby/sYqAGvoTnJjboz2uOaI211uFZlZ3YT6
FUZhmEgmN3+gJmJcGIhF1DqOncnUVXGsh0gyDHl2uwK2x/YRz078VenbA71ImixD
pfdDLoNCOwDky8tA85rBk5JmZjLiIUXqN6TV2t+KVm1x1tgJ4VixFQ3ya87/y1qW
wyKukrbcdIlTcrYq8pWiX4dJmIaQx0FowbjKZTLY1I0nPO9kWRKuKmMxxBwaR8yv
x4uxQByZKV0gnVFOUwTmHKO5iA2HVVvOcjMtNpoWVpUXgg8g70qf+N/GlqpZHo3V
W6D5dLx3q0NxIWOg9ZUfXKxwlH0xpxVqxlVdtSSdkSwnPZP3LXkj0CkGjC8j2J7/
5zkFj4jc9KHkJ8xuQRy1LdaNmhYXIQnupvS+RK0CZCjfICmuB0tOeo6LvNdbzVKE
Z+8SxcwieQh3F6VR2VNIT00VOv3L/gHhg9d5OWqcl9zRPWuMmhcOslyW2x/d5G1l
rFNwVXly8Ve/iwP+FJkPHggCUrdsMoEj7s6i0ItcK30JD31cG8kgm+r6nFMcPHk2
75jiHcFMd2umU3ZmAwlfLfbj9j6gBpNi4ac5oA6UQ4+D9IQOPLx1A8VVPqHAsGZQ
Q0rvDAkJJaCCuoXDHaf9ZOV5zAtE9rFz07QpM0zUWVcF0/QVM1LttBR7jsz6E2zP
Puw3qSL6pBMjh3pkdCYobO0VfPLjnEo7mWyZeyHXGWNplYqmqwfBJaQjEovhJnh7
B4Q9z6L0GEu8csBBXlbWoPPl2svT3Vjj28zPVdsRXbOEu316leRCnv1BnXK50XiV
hKMwYabvIn9GlwJ10Hm/1UNKcYsyaF9cHiTUMcncrlx4CN25x4Me0/+fd2juovJW
tx5n7jMh1XZHGZIzPigAfLpXvA2VwfFslfWPO8I3tjZaKVmXe+8Ac3gYzsbSF5WH
MEPT5ACi2SzvbvTuKSbC3sVzTujSntGhMUjKGiq1ERy2p8hgfxdVkXq0jK3Mm8/m
ZqJFtvKjfJ7sFLxe2PB3n5SZvqh9rjXygBY62TBvXmYRMQ4u2POEXMjz9UGp4+z8
w8yNuEuT/T6mI2sSKQSxhA60izJFbRJWbZFYrSdGAivN91b862EWw0noQM/y708+
o7xJOqK38f6vGw+so6w52nSJTYlPUL5XFjYoUbc2I5hC/ZHURFIZ9aRwFpLiiuLx
ml1vIaC5lp/Pzr6nu+AnZXkAqH66Ac/6EnNUsSZF7rlb7WhAMVYTc1yHLMaErwHT
Br+a6Shdr4SJpUYYb+m+z55pjzAJrRrUl7czGJq1IgqguUZ+gvjhJ6sLhzRxqCxA
vSZE5RasKD/5jYs1QdA/We5eBNCo+BWaWS/FIOO7XX2SCP9n0dDBieBwM4mQx76D
6rm0uLC8I7cfCtJzaTchz1ksAwPH+VBbQf3JbPHbBBZDgBvLY0OUZ28udNbtngIG
8MSrdFVDNBFXv6QoaOjF19+YL68Vf7m/JR1KZ/QAJ3i4LIZhxcwyCaounHzw/L7u
UA8irgN7Ay1HNlh/7ob7QRhAYfhbM65BX6yfPbCxbjprEu/PQ6YlaOnXMMlYuM4B
Wod6emPl6yiathtPlQ6lyVyc3wXROKl57oy9BYkAPNy9Urk68ur5MIIJQHO3ir0p
DUcXi1P1UPXVJBBV7Z2pbbImD0IOYP5Nnh5mo8RUkpp8eomwiEVa9pf6K0XeQ4ps
DNqQcK0SFqfY8W9WRaJSurEnaVrB/xRkNszdARBdv6syDamFFBXYooobUFb6kQ7D
hMm7I1mQ7p0tzAOX9sTdY+D3Yo4n9YfcqzbIqWS6qMam/ejs6ykXokQfGIgJf8AD
8mF1vgYD8IE5ZAzjs+1YCo+oeWkALj6ugiVMmtupgusKkol/aBuCN4it+tNkqyg3
b5YOINMqOgRIRJUBb4smInbAbOa3mPJQjXa3q1V5q76LoYDuWmRXZHr4D07+oTXv
bEcpEHJzyWxJIGQzvLzRpuiXr/BHCf8n5Gvyzc9p18/Qc1GwH+R4TDbdoF3/0xaX
XDB1Gb9Oc0cnoMRKQFqwITUpjt/amUf9XLSth0TjzIJfUiXEYIZhRPHZKzyGqKjP
hdsL4SPDAcRDXvSojOso3CHijKsjH6SkdSKRsQ7gmFs8xC59f0dUkf+hCKmu9yNz
CnFsC4DK5ibCpGn6d1gPcL89nLKhAv+Ky3dyALh41qG/2Io7nAc/ss7VodBqmTIr
N6hpF+NHyUI0so8y43f/2D59PvPTTowXA+ufWD3pevEsyDjPKIV2fMsA5aQddmNJ
NdYnk9FBnZ1PjjU9hraZT4Wgt2tWyLQp2gRLMRdBDGL+aSj08ydz8Z31n2vyXt88
WUzLfClWbZE6zdi9bbbTfKE14wz8dIpv6JevBKjsMIYOiQRgB4WsvFZ1z5h//2LM
7NkZwvTQaISg+J4N1nV3DON9rtD68yPnZJHRh8bfvLeZwjAmRi/lhcAtNjmO8RNx
KroKBKZ2Fm9ZtNYSCFB6XHSjv/olSB7xhj0UEjreEk7r0bIDeQfvM/yrkmGgs9CD
mJCzShC1ESlCx9wskUHx4J76ZW4fUDJvfj6QLE9NM6/JPFQVLTLN02zy1G+TG61V
GeLE+L8bPEZT3dpRXxllyzlpLOcn9oh0nns+8sYMPAhjKqENDhs++ffz4i57HxsM
yUFUGpM/pgoOPEBq9dOvAOOKK4zXx+rHPdjd8ytUsgzrHKsj0Fc6JfT6JCbHiqVQ
/13fOhHR77qfDgY+9LmTexvPoyzq1YpDtEcgesAR19dP5L3JW8DoKCR+/c0oOwc+
wNYQGn30BZHCsur04DqiWzc1+HaB8A4Z9fFyuY1s81YznL5INPbl1MvCNXrmQB7y
8h/Y64d+iGB3cBIGQSN7wyNQc9WPUR/NDiX0/gfkBXcESIQ3TyE9QC+dSRw3aqPc
8gT53bWXZFZN35it+GZupOzXSMJWZV64MhSd3RIFT3V/SzGWPbm94KV0OE9IOi/3
LFbFdVzoJsb/mCs47Br2z3ME0rMEcXSkKlGBk09CATZ3is7d70wBEMIfwEf0GNZc
wkf7/+VZBk4cIhC+1HN0riADSPdK5tZ7mMHTxM3x5N5sZyXSbbEhVtxMr4EYy3jQ
lLeeAp/JNbXUKOG3ZoLRy780JZ7hfGZGBHdOQLf72z/UGnBD1zgbziYVHVqLGl8k
ysRnw+fwIc1QDqMSUzIuAiyGcIQ8s4tF+9iLEP+LlRgadu9MWzuWFf1/puUoLqo8
CHdNI2FLaajl5SiE/pL0Q5+R3RxusR7Gpkybz8na+e4iRnV9rXLj0WJoR6pZZaQV
+26Hx9/Bt9MzEomgegFWNyHqugIlch5O+oql7yWaJPSAipIcB9G+j9C+vnUDUsNs
7MAUR9iD86FvoB6KqBKtqoXgoG/pwhaIKqw4JvrIVVrro8r0Kt5c3yzHyOHpvw7s
dubi34EaR8vgY2tAY6VN8heYpVu97vgzQNMsB/kVQG/B7CI947YGgLpDQEnirI0o
KkJh0HwKk6hMunQ+kghlvirevB7uhSSIEACB5pQfmN4+TEczwA9p4jFtSn6jEakR
FLI7qXTTWm+EoRDBnIykzISgUK9YbG9psGLygP9YeSUptZasvyYiKj1FajO4XT3p
jr1aSO5JGPGYika5lXc3LdDf2k7h7Jz5QFtjqtOPTvz1GP2ncsS1bTcPO2U6V5kY
DoS386Vuv6NE31H7oOhvZSGCEeWUn55ANmtLU25XKfa11aGrvYBG2/PQw/rWERbQ
f7L3jEzLdOuZqJDPn6dbTqleT9hfJ8VG6e4Q50wk5FAJHUD+ccLSMRuVazRGYecH
1QosT1LYRQlZA43bsw3YltaTaeyex6pKD5OO74ixmxx/wGFrP7Qf9iMRygNSVNxE
SXhETp74otNAHRnRx/u9/sGPGNFSG3kQ0KXGz6Hpua+VcN6+BRL73PFMRMfzImL4
tXhpESmNHUPJuJbe+oAWx5tKo58kHDalmfjzI/MkPLtIIs6DCx90YyYYlmMudpo2
48abIkQWBgHsQbml4SZMPWyMq+nvdG/5fRn92MmEp4AT8dccS3mgoCI5zviEgRBq
9Ry8bRIel+CBDm2oI4lx+RAHtvU7n545PgN73HK4NPKYURm4U+3a8RLXFAJniA5y
vilHubjpzWcjYQ14tdfTc8D5h54vNg5xwgFwiO9KiaYlYaFcJvaHX90nnUkImRBB
Mo5PMt7nOxNsLIuyY7WLT6zMp4+uD//DXmjqIuznEczQafFlhf3cS4S2i/ipO/2H
ytfNidGhcGb1KWiIarOr9gWK11LXFqDNkfWko0DQ4JWktPEJWdsiJdTUFEjTL4Xd
oTNAaZ4iw2OSfdolMGH18Q9BXBDJs/w1mnWQHUU3kEWP1SR6r3PNbW7AHxUvbeEM
rwtDcDUJRFmVfxmcpu06iDvHSZxAPBGZ0H4aMggkVkdW+qtcnciRAbpdEhy4eqZc
J4M3x4Wqa9vjBOQdhJqcNhigvU4r71frYAFJlzh+z7GARe8RbQmSWaaB4i69tVmT
UWsPncHEN2K9G9PN63AjtQLV5xbZ806D/eZYb/vaptmsUjzvIGJZpiKOvtBd1qoZ
7PupqwtEGyWWX9KhzUdMjmmuvw8Anu3Kt/G0fYRIvb+TZXHm03aobvrqBfkvoITf
2yIPFbM/LYCwFs14woWOWYzLkL/K6JuycZCfJJZ4V7EPdB8gwEX8vGBlcPwlUmh9
4iCKWfdiXuLqXgLPn0VhhxzB9AdkUp4Syu+NMLJbl8Ee69VYsJFQG0h3CMWJApi3
oz2RusFzWvb92vOaoEBy0HP3IfmRT3t4MxYtSiXcKBtOVIfjmOJVaIJ596/0HCkp
+ZMrp+9W53T02nkqSofTfm7WFGog5oCx6x5t/nId2zo+ccyhHZpBxQyDVohaA1TD
uV5pVGJxZEPGD0CbeQT7pxubarBsaUnsvFKBXVuFgZWuKZMXr1T/XJ3LVc0XvwXF
u7WD/ZmqkFsAY/dqKL+Ww6TsTxT9PyL0XfQCLkHHch8JqHNXzZs4uYGTyWeNfS5a
TU4Z/QM3uTYqGR1YSF9kRd0Nqo1JbjEHu/YOa8WFnMjb7RspIc9pkKFbApDs4EvO
2/gqN4Xe5xa35Ha9lINmmj7pTgJwZZicBrBDuPUH/nbNsaza3/Lor5xDrEFrsPTI
Sca2ANQN0k2b50SFQ8v1NyB6WkCx4LB4VAnlENieER/DvjR/dU0jcpQtYpGZxVgc
snp+IzMDSM8bebiWpdN538XcNpe3axPxyCuERuJYLWtGRBG3M8/ZyHlkNPZKBEH4
VfT0ALzGZi3FsgYL5tHeBtg/Mc/a7uw9zS3TNErilNIPLHzntuyUVPPv82wzxg27
8/fxOL9m3MTQRwcgSxf3GLTWHynioByM7bWkaf793SmGg+0w478xfVBxSHWapRbX
X3RgcTIFyuP0TGD8Yp4yGUj2do3qnpO/s8XKNhCh+3oT3KX/3EqcIU7P0ENC7pY9
BuHx6mclNPXY9NJEv/t79p2XqsrQThpLDvhYVnEdtmQoBbg0SFARo1oZlDfC4shI
Zk9qhlhtDNwT9wyVt0fIBoCkOkKo6061NfFVvg8G7h5GAaP51DxPtRyYfMEtKfDQ
tcJWH9VVRdbX3coMnQbzaMsVQoU3Yz9AIPbEeg+HCcaTAGZ4mn/YyMDp3wFKC3ee
pzBwMbOxV50b6N1EYuXtgjDNpYro1CY5X3sY5IiiyqgMIEK48uZ7dPmtnjqAeLl7
pZxoDw72qYZBJFEqSJOj3gDc63RfNBAphODCgLXHc7f6c6fy6AHQ5syZk6bsVlgj
sE4Dugos7m48jvPaYdD/DYzfEozUH7GOooX7wq7tpp3+fL9ip6RyDh6lWN2Rumzg
//Cg2lFMz0x6cuvMcZ3mwW8ndIcYkyonaVbDjJcDoma9xbwjQuq0H7FO299sXIQZ
Dz8TaPHbQp+4K9mOy85OmSxucNblCOtCMtkdQkeGjPSpHDk8wbfyV9Klo+zIjHCJ
2IBzziVc50WiUb9epl4+FNJ0sLv+yi8Ei3iACe6RL9GNWdnebwNNB9Ub6Gg8ka/8
CDb1kPKfKUU+/BHQ/kDpKxjFPYqDm8S7K07f0WtVkziXk82A/y1gsFG4RYiD/B/j
o6/2jpLuY/V9JS6SBOcHDvcN5gmHpOaSK/iYuVCJU0Wt8K7+f89jncN6waagrlBs
AMMnwzrC0s5t09wHf62KzvKvyGaHPWPZpcucX/9Q5d3fK0e9lTn5/p4jo0lZdvok
`pragma protect end_protected
