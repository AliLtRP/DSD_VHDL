// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bITnZ3gQzs6tvMESTRJsLjX3mVktd+uBk6HBdCnuY1lviLyme33lMiSvfqwX5TvY
oalBvzuB7JcJgvvFvHlkfg4Izu6rKDZS8nxYBGRJysGI1RjlEBO/pJcGlmgucIKC
IAwb8WNTopr/v9SrIA87lCsoOxsz2HDRhfIxNs7NzNY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2448)
cVYK/SkQfChRLbtL9Ka0Me6YgOctq3vR1oDL9ssoml+sF4GyuEPZ0SHzO1ZY6O9A
zfwDXt5SJJ5klUtPmZdcyjaDhotkk+LKPh9ztndsW96Xqkuuxq9x9DM23EgaS+Fy
8wD3ZKUTIVyKX6yzh/1QKxcKPIjN6qvkw+TWJj6XDKmQI7tr1Wl4UFfRZAL4gTW+
90/r7+kd5Q6qtmj5YMrW6Xwtu/oyDpi0AnpLgTrwZLlIl7TgKl1nI4GS95Vam2bQ
SPiltPWaa4e2qMFfYKViou7zK8TLPxPp4rvZpn3oeHWSOoxMqPozozsY1TRRz3CU
NMqs7UrHSMkRkA8IkCDr+yWluYLvRb7/e68GqqISQ1pusRApwurwv/08HdJ697rS
kbB2tHh0mTUttixpPS14+9h4abgIyGZgM6FB0x6MdsXRZFe6XGFZO2iULyMKqxSM
jPOFV1QulXKFy6KYvW41ywYzOE3bPzg/oAV0yuN+6i96TQnTbFs7RqKPdC2QgQNS
Lwix7i1QZzDferyCMEzB/8yHR8ixsFZbIOVILo8KNAz7B6Xx4euT+qqaCJIWX+Js
5jGJxlnRqBM47o4AvXIUwiS0nwR+I/5TMRMpFp9IdgVFQjpj/Mz7+dUKj0U60/4U
MmMSc7wGDKkJx+9UwE13slEVqHEtIzLFy3guNWlG2b0pZKJClwRFVWxngYrqbd8j
CpCCOfn8zQZzOh4NmHRy6HhhsOVp4LjqIrc2c0V+UvljrodDAU/yTF8Hwln7uZQT
W/HJGb9ZWOfi/uzLWpz1aOR0zW1/GNMHNmPLPH0su/Kk1X7spyWfdg2gxwnwe1YC
QfFrJZWMmEDPCDPebNOH+gt87ejp0dgbHvgsPqIpXbbOS580jda55812fMXh6Qj0
1wyGCvXSTQonHRRI0DCoFro2cd/gugzK2ju659L0vn6FwVPzRqzm4dYR8aNgSEwa
sr/w1iMHqnLKHDQ1HTyMCjnfl9UVAnOPtCLLttrR9VsbRm6rVm/9F5n+IEGeY82+
Y3diQgyQNxD7KQNOJ/RoLXk9fkh2YOsHD98yacWKfLOUex0I4/a+mWL6JTqsc52H
545ICwkpAOr78wuYI6x+CwEXImjMvYIX0v3u0opbei7uuB6Htj5bKyTGqDJxTOW9
9GRxprNJ2iIh/1D61VkFIr92D2kJsdLCyqyiwOUVKm5lMqJcSmdQd3VOXCRiNl6K
0uLGdVSv35s7tH2WjMzjsEkGFTrKoVDSrUxU1Qkmq6En5cfi8q8SrfhU20+PZhow
++j0sDhpUyEGnX+Drd+RtDBbz/c0Xmp9Wrv4DCo5NWx+49+AJc9Ww4U/WnX2Zpwq
bv1bcL5OxxoqlrC9rhmAYsX20tHkBpzlHnj4vH2AKDyT6d1rxsm3Xjus4IfYrpKX
eHi30QkSlQ9ZHP4G3ZASAGpTEsfVrBrC3VsJlht9CpwPK+j48onyGdM16XaCrnzs
z8+xVU8d9Boyg15pFf0Ix6bkZ5A7cKVgKc9DmcB2610Kk7ZQ2EH06JLFnSil+Dx1
1ZcE0w1zaa7xKmOITkG32qbImybTeeozHEaqF8FX7vJEPGnK0aJD5I3YT0nEypN0
TKGZOmGOwRyy5zgCluK/kw8q43gPbjcMuOE3s3FH6I2CzkUvACNpTGHI0tBwXy26
N4DvR2K/jf24iV+X204ASav6dT1bCLW/KNuenkUeGN9TuTzI8tvSd5Qhl4XGrBbR
9vNkGpeMpD/dAKJ/G2TblKolxZVA2aJeGK6qizdaGsG6x0Zc6rBxm+iDek0+ftzH
EbGeV8fuWYR1U4iL3DZ7wQ6O1nPT1El5fvVUF12+8bQQ5rjfidfhThqyqIokTlGd
YmrppSVoxJBWKQPaJeYRqNFt/KInBRgpkanZDjMH2A5upRrqXzg0W8F/a+8FEzqk
ml1cViZ1lqpnI6U2VDNBH+59ReuSTGb7UkAPurTVPNU+z2NQ2WYTP2A1bSNw+4PW
rFLzl6MwseC+075EHmbQECGos4bVg/kxoQ2hhAaJ+7vvzHJG9W0imq2fJBnozWbp
pKlUUzfUOT8UX4rx16uCEwGPqVv6TL7ftGN2hH7DmRVuAgDuPmRsa89sDhP9/ehq
QNCX5xVSNXXANZ5rbPuNg1OHQohiPWhm+F2RG2ljNekZeh381wTy+Eg3xZCsxtRG
KYLIKFWpojv5pTlaL1U3FEWTVVg5tDqutQwa2AUKPXKgHNKq10Ze5rMPmmhY03Cd
MGeA9vgP13iUk6Bb3DLjf0G5cmrEOnRpqugnsXOW5SpJip+VV7GvLokVF8a9hYJJ
YCklJ+exdJjiASa/xIXQIKjcWAcZ2fQxonvYaCmKZHpRhjOEs+HmOKK/h5X0EDQo
FAPKDp+acyF4ow5HGPAK+ux+aOgkUNy4btIUnznVXJ3LCcTYrf2NOBlPsDMd1Wwy
+/zKhvmj09a40HwhkNXepS8Juow8/LttcEXdHEnBBGNmDwp+7oGJbCaSi61T3H+D
J75Q8hNpPVMK3Af81zhT2WiApFrVlKqrOG2eelc9ALrm1SD6BI+ZIVOPj2r8zU3H
ndg1AFfbWuxyImkj3vq1EWSlbne0/nlXIs0SyM7GAmOnc+rLtHNfKyEe2VE16kxa
hc3I0tEPmWki4ndrRCxgMbdaeMhvMSFwPrBuB21+GKl424XHscKMO+dK6sXnJEQW
bW0voSgaLySTKMeF45IhnekS15ixfXN06CpxIgQdECUnqUKheAAeuZOC6w+xphjI
CQoki/zteqv878C4wKTQhhOnsLnwP2jDzEnmIUHL0K3ds5OawbYTrN0N1tEZRdME
akF1IxwbTH+Q5fq98kXjwZUL/gEP7026IKTjvIDYiTFG0kk/xv3K47s25YWVS+bA
dFPDsdZAfwvhmSuj2mAArMhXJhvz6wwxZC/3NEGUKWS0z/hJIXXWDov6UOZcl3N0
YhF784zNTIBDytYQMtliXI66xGh4GRqbFHyE023bIvGAtPvzUlTWHtPctwvVePp5
hVR92XZqPwfbwZPV5sE40vjz6zWioEit55oqYkuUvNXlMS0wOfV7GclKm2Ag8Y+j
3oiGVbp+XET0vjNZqTP4kI0wV1CBhbm8v2Sb3wgqF4OO5g2tMnW0yhRPu/L2Zttp
ovIRf1o3FjZ6wvluounr8kzHgi06LYuIkDzrtATMAz9yknedG1L2IORfktGvI5P+
FUIAxy/LxotbAp3TA1srLqjGqZTHsar/XQWBx1e8Y5+m6lLC3uEI72xBwU48IiMl
`pragma protect end_protected
