// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nLtQWgxj1SXnLflBtqGczlyrrqQWcSKYh9WpmReFiN9QeK/qhFsws0WLw7MzeJJ4
+xIXW1qlGIE5Lbc7vl87+qqZFI+3qFDIBA5+VVw5m7XneYkXWz0dN4U8gmYgL2jt
6mTNq8CeIq2Hig4CEjRT3ztx1KHml2/VDCw/zxhi80Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6400)
XmToKeSrM+5YA+VRxQOvKNuCMyp6udunRnBSGGKIY4mcDxzBkHAR52Lf/z39Y7js
5CDo1YcuKveBvcoWNl6bpZhnbtNc2RVZleVorHL2SFUsu0FgJ2Ly0HrA6EC5kh8c
DxcHBbfFV5fh7fIGDfh6DmFXLf/ZRQicl78/oyOc60gfY56gMsx85oLo+XUDbUBf
nQZGSBdVpD3QzkPSuyZaSp5nUwVQY3X9t+QVgc3H3+xLSqjSOyUXm4X4Wakg6R7v
Iffd6Iooy4jmv+f0moStC9PSCZ6+VBtqv2mgC2ZXk8EdyYLYg+aixndzsHmJX+GN
8VyshMMh9LJxdjt/27bs3zMtXfGsY5F11UCnOutvnOXCTK6YyPzI5rR2yvE9yzS2
Ys8tmmt7Edx50dSMFicazFrtULshwf75ovjFKJ3w+wNlnGwKPV/c2Oq4i4l6+4ZK
lDHrjMFcNNUa2Nhe+7EKVnlKXI4ALHJzimdHj/N+BYiXNXigRjck5zbrgigDpgKK
rL8MCCuTj3tKKiQFn/oJLO56i4CyrsfPXanxOAGUYANLnnpf45q2PjHlNxG5P4u7
SZaom0eeVSgXdgVGxf68vuap2Hf2O7x2cQm1TgM+aHyxaOfBrM0Ot9jVEvCyyEa4
tufaH4yDKLYZnHOIPa+oYLOH16mByRziHUBX+ckb4/GbC35ONevIZ4y7tUE0uYK0
/DBFZEzghdil1yLhg0NJVPtec3lhqLjvxUE20TX15KCl2xTvT2hAzlo1gpNoIHVE
ivO9Qda8xtGUHLhwIvPagCJebgtWounWBRDkBeZYzLQjzI3x3VUJOYKip5XJA9A+
2Sb6gJacrwsUOeYEVUJYS3jCim4Z1eFHRmPacgPOOf1xWrtbSIStXylmBvjZ0Ufz
PrXAN0weZKlqMoXTthFpYD4TNFaqwxWBtPr4jTXYaHQxBpfaxFQ8SMp/dt9Up9hg
AEnB3SgNiX6FmxCkT9QthkujzjXpXiOxaGbh7HsKrW5gXlD2v/Kb0Ycw/72Xr9C4
IZTs1YwYtno/DMEacofzoxBAPUXAaQj2yMXcj0O/3f9HIsEjV3N4k/S+HlPUe0jn
K2p2vt5sQqltI6f4pMuXURJtAIRmv4XB0w4hDRIZT7THeUD415nSwGGLNjm93qkr
fR8ociEgvC6QyKGYWzMNPwSEjMLd9d5BcvmvAC+bI9qcdxxTeYxm+DAjGpA8TMqJ
HMtTGKPo92pzRdnJYV5eltr/x3LXfG8dc35wn+stvDm2WfsuVtxqhJ5QNuadb0wL
C5aIlGYjnlA12aoStES6G796Asc/5eOKZWZtvlbpwrru7H4OaCMFylGRvwMd7ao6
Jo0H+ykfpNyKeKt+1zcpGnFN8IeH8yp9IztnKCO/EYWna8i5LYLQXM2gZDyYe2Cn
JA8ag7p38nOuLUvnzbf3tMYHMQR/FihbtQdsZS+cg5Mi5Ev4D7Bc+C5NK4kNcKsi
NCln6nXceKVJlujn747tPlOEexyFWyct4rNZm7a7JsrTbA0FsLAc5gdDV/jlv5xb
d0fAMewvmcqGZjXm1/vT0AS37cTiwY8yUkgvnRpBWY5kcCNp8hiJwdlwfctHfXRA
PQtCxKjN8icC/gHbmKak89jMU4dvQk5NwB8mkhphZLW9KaNjf+R7ar8jcBwozewM
aPpkaAzZJP6vqHHRLJLLYCfcfnpNslUtKT4cc005CGAEpmC8T2Ke8LDRS1x0EjOu
UjavemqCmk/Ksflw7/OTSbrGk/1Uj1qHigb1Ud/v9Olfqrb6lEl940SA7TkMsXbh
EP6UCH2H/TZQcVP3SZPgxL4Kr+G52+KWpIx0wuS6giV/H/hoM9yODDhw2sNqk2ag
KKyGMDPmN/ozbF8ACfnwqGRbQeK12CYuLwSBxQqEALhS1wIRXCylTSJU7KqJEzNi
BdrSSDtZwKTzJKjSAyP0FZSfhkHPrP43s8+m5SbHRwGolTJKlG4wl8RzNgg0afrW
vS7smZstNpGV5cW4ka+zLY5qA+mJ57isAALNokFWoXq24lc1xG0zHvvc1hM+oOPP
VLZvJTi/tkkQShVjMjHHuB31KIdoErb6IuukY5lsdWn1Ndn7kgRabib7WGYYpxMB
Vp2hhUQUJk2Rt9KH5wMHuryDboxmAyXxaE4jzmVpyuXRJZKnXbBwHKmHs3UkV/9v
fzI9EKP1/LfPosi93qLqh/Jx3De6BT4HhOqN8pPkh1pG9pO5hFw+GDIcoVPu9Km7
fGCqdug/FGj8H6cPj/zxT7cQOntTwHCNRdEY+MzK9s/J556f0XSc63v3dSMnyTen
vbaM3vK8fLW7GvSTizTYxpNKXa49UEDYKIvbmZxhgOjjahV+iqngDR87B/VnjH5/
JH96yZXDp9EnAmTETjmHrTZ1LrOZAbug7QrFFXvabB3cvPCHow/CVZmonHJrl7BQ
2pr3jnOmxaWlqAnbN3BfCpwXO+OGkKZueoWATGIDKdNfvBYmOgSzRw6WI2BT1hEU
9/zzeKPBWGqMlLkjluAWs7UJvjDv60TX9Qm9Wo/DuxkQZohifIJ2jLdvrmnRIQPk
HuI1YbOJKMQPeZXWFUStj0LQctfNsITiyKfq/X/xu0UQPb8c6rPiWb5rylsFD2J8
stNGdBLg3SvcWG9zbQSqCUj9UDXEhwLYQNojsEHX3Et3XZ1asNbY0ngrd/T8Hb/L
vTyWBWUMyI04yrlMpzXwJHn9rsIT+4h/BTFmWGuEt3ZFfi/u9U4B8itwnzlESdW2
kK05HJZ4FGc2J9A6ASI5gbdAEZr6tC2TWtWPJ76SgVDM7ZgBDXx6H7whpRh+saN4
4BZyBkOqqySHO/mX/Vdk1bNNwK5x+F7xEFyY/OqKoXCrpBxDTuIuxLG85l4qE6qm
EM3RRYPW69a7Ye2Pkn7CpfsrRIWyhf1a1evp0spABkxL/N280a9U83gS3+i0nqp7
tSRcBTKrNxFfifMNyVTK8x33N/TDPPuIudq0o3eSfUw5qR4Yc3cJv0815jkwSMQs
bObTF1hcMgNVYoQghMDJmDX5eBIaMZvoKuENitxFU+UIfPs0QTkPz3aT1lxa+43Z
qwZAP6OrmvIU3Pn/X5wDmwLzpNUveWogUWbf9shj2/Btzp+M7qimQLr7Z8FXrj2l
Qdf1rWTrCSI8kDpNs03sT6E3ag/IO9YORpEMCXbasWJBoucm49zqnRTNEFgOzS0x
yTZuL/JV43kUpzKaeaBL8ZtqVJGTGcIMbznkI1k0fOKrlfoppZp8JXZ0GJE8s4Jm
oyRDKHpprzEiYtoca7rOfFH+mP9HWM3HgNEJHW4K85B3DYKFYN504osQ5EDq8IIK
+7yqQuVwaVm4j3SrCRNw47XY2b67Jgr8nUcAFC2is39RW7miGYW2rN6e2nuaMeBN
TFalpJ/AO4e71w0m9yvf2jxBZWFTTE9SuHT4OGkw3prw4YmgKDOCd7tc5HHsp1bd
aakvgQWOZbELb5tiEwaYp8G/poM6Dlq5+74uY67fxEAZ2prRUkhY9d2fW0/QhZph
8EZAFkbqrahyXF8PRlHtcfxN1EAFpLu6eaysCuFXj2ZNZXHJxd9T/YW8aUlqchvM
AXLgG/g6PdjJeXY21BbvJbva4VPOMTu5vyK6qYC2bxNSbQruxj5nJwXeEQMkN44V
P7e2AuBMyXJJa1UNFvej2UO89OhePajEOykkjg8kki28yLSRT1sGbqVJUOLEPYEr
FOiP6LBl4sZ5brpKIjJ0rE4hmlpamkg6DlE31ruixVGTRl/GrhMnizWueKPLk3yv
a8aT/JQZJK8FTpW8ZUK0z7LUkfRa43InE25Xl+5IMcU93J9IlVUXxFXOrmmOFiY+
UJbj5Udc2MSuOgG52BSP59iNGyuJhqFmz56qfjnebgG0rpjKIaxDDIdgllr3CVbE
abaa8LwEs8BSHpviMy5iov+RBJivbmezo9UOlUMfb5/WogrQFN3O8kIxp3mUFOtR
JOR4qzhJRDBA5NYGTD9HeM2Q+Ze+Qfpz05DTgK6ofCE1W5JSHZW+Ufu54rnQu9ok
OGl26CDDrGMOy8r9klH0h6to9bkNs4Xo2EFLNIuY/8cIo/jTvNb3FZ/O0oqvpkPC
Uf8xlVMeltp0Qx/QYZ3p0gPGVERQKv5xFfY6g+571m5jPZttek1hT+BEtOATGRHE
LZ5UZ1Nl83sZflgl+iGsKRdQHxDjfZ4KZDhmL7IrR6vMoMmk2toqmBuS84D1ssVO
SsbVsDiSo6TCRZ46V3RZvMvICOdLV56chY477sNnGP6THa41ke7Yrz5y0mXezv0v
GV+bNBq93prTwsMIkUcW44wJfGUD4UbVk4UIxtkVRSfq50WbUrmPnU4FPk+kpaLT
tVJ9/oDAE2ngdPQd3lsoFsl33bBZVCiIPCXvacwADoYEwZjYqvutfXQUWeWKF/Q1
4MxLsCWHfclrWYHcdM7KNm+Ve13v7nd4C0rFAEDTayi9OQb5sAMB5qvmcLDuPGMp
+54+/aITFcKjQKnZWc8q9t3MfWppp2j3b3WD/NSsGeuDmEY7TfyaZn22SUTfwuul
w225p2iquzMF4Ba/ddYFXFrPoAdSVbtoje09fFD5TAImubqxgy0OZ3c9t12p0ArA
+HSLoFqQOExyeDxY3FNSxea72RNVDtd2NgHBi2GUNdkxU98KQwvVz4NV8yUUmKYV
OEP+p1z7ZKM7N0Y01nIgHc4wAbchctoH65OzHXYY89Xccm6VwciQFZeIYd1qV9dC
B3rbOtYCzK2i+pvvwUrFQM5lc8mXACuDfTwu3ualeu2z+ORmf0zpd+5V2WZaxAvW
neGmprtvX9xO0dlUXxbxpEG1OlDSvlLtclrxv/0T2BdCPskvvwPUUdHlOBj3Vg1x
pog89vKix4PgRHBAYM2D3FiPwWFu5D8/dAamlUCyQes/fycYQdudmfR8OqUPl8Nz
kHmimhMvQKBBw4pZlLnq1kal/WejqzwotiVPvrgodQF2e1+yqNiU14KGtEnYiHgp
ru/2ObDZM+Rp4dXah5MLpmknMOAADQjkfZR9fQyirwXMtliHcC9DUXS78y8CcxBC
LjtIXeIlNzRHnDHFXYNbRWe+U8JZ0Zqf2Blo6ZV/LL0Zn6nOQsEU6I7JoQ3YjeBE
3r/y+ohWb3mw9oenKMjW2L/nFDewtjmB9R/9pazmNtEKsX6hQsFrUrr6/6lK779L
OEPzMnKnMcPBDrA8avzMKq/9G/yyQGQr5WgMw/64dVnjLQESDeAAoUWJyfpRvf7f
1WaVmAmA6amAYnhMZ/xnvESKEVBaTpQmnuLyOt3GBHL/I1zlqzmzdO9K9EDVblaw
/taRtocMkEo0JhUT0VjzkMIRhN4RnHMsBXXhr+1vM+AFRnKpvxPTjLRNByQmdplG
iWLM/gBrdRs1M80hDV77ncrWn+jjcQwR5vEYPYnZc3FFzZFWCyeh712JgBCHLvq+
IiCW8GVseZ8zrdWNu8/8awWCgBMwtts1Ug6UZNWrX0Lf+BqGqceqx4uZ672zpKbT
BFiQhY1MGoj4LrFpkUv++p8ut+t4S7qNiTlL81jO4Xgwee9yLp6z6csflVFQ/H4w
6VpIc4qkCd/jYBhkoNHEMbFYeustuaVq1KMqzm2lv3t7BGyecaT5JYPMwZaPfNgw
R+29qCHfPnjeeTZSq9ju7XyQrSHDLWN1Si1nZ0+Qf3e0+31WhnDtTazUKFJuoGFk
tltxMV35kEpn1ZX3SgmzEDu8Jcz7J9Gm52E6pJiIX3Cz9B5k8CBacRJPZ4tZ+29l
kN9168qboWBDF7ADSXIrxPZ5QjoAY4AMPl8glFbi8br1sVzCLLQqghGq2YCn31L7
im+ru4XB3SzBaYa0bvMF3RUaPAo2HNw069yEY7BQ8Cj5+wNBRrOZkxGF91UbtOE+
Kk4GlhPuAae+BXlhjWV1r+5W8Ww3sI0f1O3a4myhytJkBPeYXLbx29v/5aVk4QqV
4NnhJTdIjRn8AigFbUV6acBELBr0vCxFjM3FgMiUjcAdz6i1jnAzfvu/lyR3Zsby
s01CMRvHfcAIpGlokqP5XZ9lUylxROheApohUdusranASCy2tdba/OAo/6dCZrDe
fotMDUl5SvWc7xWyD5vfGEk7Co+O6yAToCbL9PZJS9BJ3jHBuRKzPf4cfck9BaXV
j6lDTwcGW429TQ+pBmk094EuP5Obsqh0+wdn3p2ZlcdYIBqJgyTXqpAUlx0OSeMP
yTh2PzBq4so5ejSdHnsWIrIds6D6pFqnY+AM+grkAC0kl5IyaZ+ck+bzZfsUI4r5
MOTKK4EJbtoEepiQM+5sn72DKDdeOgqsZL05DVH0pJ9XOESF4OGvgq2ZnNO/qF7g
Xe/gnJ31jwp7AwcILehJ/c2P4wRRrMaVJVpl9HqZfEJTP54xmchK7X08YqDemMIX
j1SHnj7RCIRpZ4IjJYW3s0OELtalHs2iA2HwnQKevI/5Gu8LpzWy7sFLEZ9Uc1Ve
KCnuaW1qLsZHFYz3Ur/1hx3wpSn3Et3tnsABbMMk99ppaIgWp1u1IUGZg6EeupRx
q0o9vC/U4360l3Z3uesXu6z4kMAQYodctIKLM9odubqeMiNF5LRXty7ctrX0H+no
RYNriX8d6ln2+yeOWAFAEfG9LB3jLqHmHTsO5pF7SMBYYULJvP+QfUrbi8NynHWu
UlnmIcmFKFfOaQLLBAKPg1UkbLHkE6Edv3YxXIcbaLQzS3AiNosXp3OkZ/mnRlMx
Xdp3AtGFJRv/unwY4ka/p9QGoKwGmaUPXGIYqqTWvSxFHYSPrK91CaB8XSqgDK+j
/9aiH0HNtGOYFvmHahSPc1Pcl9FxKI36kp36if1DYJ2ge9lgxCGkYc62r7Piufze
dkykKYPUe+UyHAbZmj6Ly/Kk1pfWFpmTVvmKOxx4eM/TXVLfOYwjF/CL9heAwejR
ChrCn3DTpX7ge06AkC4Nmnn+xjU04v8YiTnXRovTYP5rovisCFSzSxOTSRf5Tbgb
Ti4RKy2GQYPxh6RMFD9Jzs84aANCX4dLYw8BFktV5nZN/xFffvcEbYFWJudXi4wE
P4Ke9cAt8AUUQCKimmloaivmqCjkqH9BAtNvxqFxC1Q23nsdKvnlNqQEAdZULnYH
2QAZhmKloCT14FU6yZ8Ppt556AIAoevyy8OnmuYdhcCSFQG1bCxVLYBV6HQOSrEf
uhwdxVrTB7UShuqwQtZL8RkpeZFSUOAPSMb9CYfbekQCZ1NXW4ertLSeMyikV69d
sIjbIrpG/y9JVaNXu5zKb9BoeKySK6BBFm0TcjlibR+5p9vLTW1Z7dd++U7cYYk2
guf89DvNLB3fPuJaDbF78CBrw8QxwGA4GAesQM9IVrnzeufHErh4z8PGUM2gUslf
7qLdI4+7/eSqq5IMSU7N2jEh9eqhlikXCC5ozWMtdArz8PnWMr3cWjNn3mMLrlHv
H83R7zB1MmkuSovT5NuI9xMEw8fKF7K+W3dkyd+3O3WBCiXM8STJfQ4gSwD1r/XL
e9HdTR4KbT+8q6gmvMKN7Dazr7nuDRfKSwGtIruxz3XoYvwyJNk0te7OLSpg02Rm
PcpMB0ry6DBBrXd8aVL3fvAn0GZgw0VEyMVjgxeeKHWLyoYCzoUZnt9cogk68PnV
bHxDPpJseWrnDYgz6LiDDmUGQ7R8Rsox979Rb5WYJq2U1rln/gi1J5gffz1WAQiK
EawboTD2ckrcA6+pkZeYDg6oppgKmOMKs4AMOC8S06ULmmcyFxHqW+3Jg9lD9pvo
6FGpaqQVjD9PIYz3Xza6fuW0bUzuQOovZoQa97ZmRtk4NhUf214Mi0BVaw60RbFn
0y5yDKtLzebxCtA7FvlHIkmcBksOZ0xCBBlNRJ4DLGYfD/k/cXzaLoyDnME21543
DGwg8YqNB4bx1ThfWlf3or+WwqVt2opbu8sqE4Nh2//KUw7UBw5NXOp/F6c1NC3j
sIRea4U3bP5ydEMm2k9/YsMMEW6TOSs+8aa9kyRLh2DfKdG030Xptl+NbXrBYwMA
8qbMCmnfdu7+NELBtRT2ep4VYBw0PA8PciRflh0rnPu4CHdzbsN38ZPaqkk+Fl3b
NuN4SxlTjcKrySednG95nuEG2G0BG0IgEW88Inf+NaWcXb/yF+mxNO9NTJkFM/ez
59F8H7elJaTuQ6m6p3cDAPC3G1UT6OzAqmxpyfqQDVLbSjIzXN1N2puEiEFfrrOE
VM5l0OjrDnV7J6TCmfzHk0GTePfjeUaRzOTPcQpeObF96X4b2J9HmH0fpEs1gigD
SUpB/T3JrA5yxbJGY+ZCa4kMMVAynqIGRuNKvSZ8s8kBZVTTQIKlnZNq/uRui4Yi
KZDPuGFNOTNd2bhtVnfMi5PrLUiYGxhuZvXoQbyimLCBZCR3Zxk7sX5gzy/WLROh
7ou587ysU7OeCdPmEHVZRN0Gc87IX8IhjCQ3zn68iQyJ77K+4qvyNpL0YFVsYZYO
XjvUZfB0AU9uxOMD4el+nluvCmE39SA8c6jkO0bB4JD8oe+GwcSVjUKKDybgw2zW
Ax1Kfv5meJdrpvNdCSnnbw==
`pragma protect end_protected
