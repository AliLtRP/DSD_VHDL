// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RKFo+EKcR8IFXiJPVlEXh8D+KYkxYO369Woi6p65QvRluum9Pbwv6cwidED5S8l4
BXCAVt8lXLO1ZgasuX0hV1xsAvLAUZW3I3pc5IDw2036UHCRkwkHILyzECbT6y8g
3BToC3dDP6FLk0GCxpI0yjqN6FQ40kIfoBgWP1brFag=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 23488)
Lpk8Lg83a5uktCRLtdBjLpuUnyTfmPGnVDH5q8EvGsio3VRQWeaI2pQKH5PXlgyd
4fR1DGT0FOeuegIIm03iA+OyZzPrC/KUh1gCCbTI1ATc5Muo0/UKkdxU/N99W0pC
tYNFB7X9uGtdGneiqvVS5AA5Y4vpt4ovsGs3c91iLbNWHKZULf4u4Bqu9/hET3PA
hXlwS+tB2IzasaNs8O5tp6zDZmJ5KI2YwTsWLNMGxC5bFsbafXZ3QmJVVMmHjFBn
BEhHrpaK4IIuFQ64FY3QBcQdF89c99e3VkHKp3ZPvZ4/NMydO0429OjN7XDAGjzV
kdZrKZdMFRMutltGtOuGpAGY6+O0zMoMvVI5YJzb8J4fKKA9xJ/yLuajryYpYREd
cXFzeO1ukKBklfAS38WY1dB4f21Qu1TcoI6v2v1c7ceomErNoBYqRUAWjI9goaIC
Ark+9DNxoZeBBHzKbmcj+TWLyWMjFLq5M12vO5pCa2gBxw8sEQHdpvWpu+e/npHY
sKwa0X+m1L2lKeiBpQIjJ2OzRXOVDjijJb0dZJYnTFMtUCI8gybPhyB2iOpg0ah3
8Yx50w8o1OEPWSl2XxHZLwy/P7sq6ej/LkYpYUF++5CyLHayLLmgdGRmgQmvCCFR
TPF7iQrpWf40usCzj08K1yi+S3/Xv/IjTL7JU3AqZdNIYslprEDjmrmGueyR+X8i
3y0cWOXwpte0UGMo6cvCRipkrXhl6nlcPvz+CRz8aLSrwYlvSy1Orf+kWXFDoMhp
M1yNpANjUcDhPJQSU5Q4e6JwXls4I+3YYZW828Z10iYSJYX98jhLDyO3gBrhmZEt
bjjci5xumeeS8OW1iesChpO7P8zWO3ezkKPCiNTOOBEa+3qtQGUDDhI7uwadqOlv
5M8Yf3TifhJaQeyzB5MIvvb9bt75kekeJ458TThGFeJy3psjf+SyztBUoEJWkez9
nfBtSUT6Q3V5pfox1+NTQpb4Bk1lmpCzDnRUFDYZSKWgumpGOTpiYvdhstJnCJoS
32UUczF2l4shCdwRGfBzoPcCtXoBNnGqUXx129Vl6GYNYNsvCerpKVFKrogYDOih
uFGkBcQECm3bj29Y/wZeee9sqxGZ4tCuKnxVTMDdfYp27LRo6y0iW3UA+HjyBZst
Tf1SIwFUn2na6wHKh5cUX8GP24+bYgyivewibEASo1zVpmHLZ3F+YWNq8l9dM071
Hog2vKnAZub06p4DY43wK1Kf6hqgb62FZ1DvzwlzwWRWLWMjS4KYYDgzFxlMy8Pq
9Y3DapfeU34Ui6+QWVTOfIvQrK3ZE2OcWH3wi7phk0SIo4+0uDQgwJh3iI7rVbq0
Wcb9w4snMAsttJog31t38U+iGbI0QE5roU2ez4McWg48FlY7DnD001cSqnL8Q/Bh
Jhtc96hYiq6wW7ibANI4M5zq0Pza+4NiRt7nU3LUUgtUQKWsfNXesWXJSVs1AD56
now7Y9/1vwaGaxVEBFDeCcBwOkcNVnKtS87O/qPoW716pu3CSmvT1FhQtB1P2aza
CfrLF2Usrb9hASY/K2wTkYW0W1Ha3s1tbLD9M4yrnbnLELAybXbHHl8OtHu9Bqdi
l8kCosBY37ltGVLXha7vjSHhtR7F2FZH13vrTyVCJLLed7OTC+gs4SlWD2bUvrVx
z1lDsT5YJpQHDRC1S9wafdU9M2ROKBh9WYUhccfxgbtDXk4M59r6MRDUUKSeyncJ
ws1SVufH03D71WSaXwLerH6neyqOtVWk25Z0okM2c65hY1pA93hgoWSjm9hnECpe
aIWDCe1e3Uyr1LI6ID4SP+nSzgSuQOPqz71k0Gq5q9TpRm0Beb6PKBP64++9z5Hs
ZIkYX2ocQSEzE8VuvK5+GOOs5R4AcqpsvVamWhoiHN9WNaRBsgHnEHyC3Svr/BB9
utzsOexGfFTopoo7IDlgINg3KWti4N2GLdf8te4RtOory9On87PhOYwcfVEcV4xS
kYjgR1JJtcTIsPIGtHgT8HFebFgy9WlKFtOZwIz0NfTET463MSvhU4ab56t559Xh
dcWX6Xpr+4F+XAmnKdcF/tOtyj+CLj4AWZWwcAvdD+y/PDw2KWgwQclbB7l2V3Kz
E0WudEV62cgQGDm5NxbiKNxKmuryDvDU6UHtPNWUULQz3BOWyHyopCWz8Ijz+989
qAjR74oYk3Fm9jQ19fvH5AbFKpJhCDtWPO/Pd3b9+PWeBQmSkVJF1cvcKTWF0izR
1BboF/UhIMvZSQ+t+kwR1l3ZCkl9PVkyJ8Wy88SIQdLRIQNoJJDj25AMFhG9+Lfa
82MH4CSVpr5vdHqaixm3PSkyYs3h2DsVeUtxaVNVsJyg0Cx00Ue5tMHP4GbzeR+b
77hRlsC6ZVQnlA73m33h1D8m+Xbbg63CYV+i6EXFrcaTVEJhwckQTaRNcI0incZl
Cln4u7rm/LeqsjKX/8mUXUnLSNM7+nnHxxuXWrg50syqsEENumGUTVXaV3nA9dZ/
g6klAuGivyGiLoUNC3I6Xrqyklp8VckSc52G1Vd30Nzts3/EvZNRq50Tq0RIUezt
j+X5aUefb7c/8bpW/uVM4Uk5megzBPqSpqrBz/jkBd2tjggvkgQs1HC4T/KKUVdi
Dz8pVLXZDz0bEKD1KpZ9aNZ3WUTz3DQwyodEtCa7AXOf+18QXL1q/2voU6n19L7k
sayV+szOJ8YGY70iAfeK5hH541SJ2axsAyxdVt8vasncA7U6KGrVvYzwyiuOibAz
O88QxWfjhzZEnDmSFoRNg6xHBWDvE4LVQYjUTlGdbe9MI9d5XXsW2PWFhxZVbIuL
lVF/2usu0J4hJnGuAMLh/Ac5uvCiNE18/noGnxvc7AG29piO7/6vggzs6zLdfn92
E9zvDgJYMYIrOzrVSlRDnJRPHoMbyCR+4XjFnhcYnBev5tVGhb0V8svpIIK9NzOC
bMby54x35ffGY9i0v26yy2vZYUyY23FNzIT0oGcoz+yLe8xR4XVFS4Rrxzu/yE7j
DP3QrwKC+BRj3DZEtMt6QrLdS8y31aWLhj2mFqMcpk7whB+AaOq3LTtcuLo02LSC
NH90iSKyae3gqnQNso3CVnIbsJkX4orqieMu3HRX71Ad9k3zE+10zNz3JJKRH1j0
xxyLUrDuPpA/QGjbx7Mr+gLFYPu3yYnDzeS6SO8UntD2/f/b0/fWhCmTg3MimW6I
BMdGwgl/vQeinMo3U2RAP+e4PDqsATiN2LnABZKyAlx6B350JyPHfUbKRvfmpkNw
aV3Pju7z/huDwbSpxfoxRC4zEFYSHu8HnuO/IhdkzUnifw76OnCmvTj7H9Oy3bpk
ZnDTZvS8reub4gJ5hw7/UEnr65wTMaDbgC/9noCldxyqvNJnntlUwBjW7qECjp9R
CZZbaXJDO1PER1aX1vB36EPSJcejryhqQLTHA2qLqDI8CZtZEN/igsGFeJcyXOIt
LV4AW0faQVAqn2bUoiPeu0UQxeNs5FwjApUgmFMHHZz/Y4F+QEhIEKwU+vLmfrMO
hwWL3SISc7/oJfwD9iJL7oqTV/6kn4NAsvu+aCv2RDgDVingNzykiJ2/RvX60ogP
gXC4fM7cRtKfoaJ7pohYQglWhS+KhoqD7yQObOJQ3DNmpoW4BNKIxAVDECUmZlCG
ikP87rgaaRoEEBET2j4B2Lw+i8G2C2n75wIyuOA6wAFy3RB9Lg5Nr9MtPVVrkZDt
4MDUVeji2qHcY0DEPjnpn2M9nGSVeppcoZkRbmw/tIwq/IRbf5sM4dqF9kLKg79j
kBE2R39DTHfu6hbZWNJ5AmDUkZwbNDga+OYc7fYyhHLcXfH2RmtIFCh6yrvHT9DC
Iv0wsM3a400ArnGX0puSLnFNHjMrBYvBXa2+Xj0/uxBmuYenxe8LWWyGFx7/CEvf
fweUXa/9lvSuhkvwuJII72chAU6MpColpiDXgMXeNKbzTKpcoZtXJ1sSXbpcrXSl
/ua5AA4llowHDkSrTFSsTLwm3su6demt8RhVJr/XjygijtrL7aukKwP/x8Q+n9Ic
ixqnUhmqCDTinn2GOu34suYQEp4UKNIuKXYrx3yxTT58KeTEBipO1A9TcrZ6tZfL
uJqBJpzOQJ6FjpzIBqtLjAekc6scXy66ztGRtoXBIQQiAuKHIXkDD4Xgyi8K0T6K
OXCfdXUWWn6Tiz+DmbZWMTyqnnjVyDeYFhQq6B/woOnQ2xJZ6SpLjziQFlmjytVM
afpeulVuLxHKEjaf1TQ8XkdIWOVNvVehap0dBKEy9B2IsjsEdk0e1iaKK8sQIpAB
++WOlJqZMC4L118Gz3zyYyPHH6d4crKgbJyci1TRWIqBOU5jsLfawphod/PKOreX
1GKKGZ2Q8hvp0z4lWlHldYpDT//sTRujnijESEQ5rk+N9rriQlTxJ0sgL3cr3S+p
HOBsmLxd4ETD9ewNP7LtDZl/8t5pQVaIasF9KkDX2+5h/D08GlXk0f6O0h07gPSJ
pC5acQdmHt/tpq05kTR8zSCFBqFi1HG0zRKPZGSeSbhZiYz+yKtffE+eeFR9mHKA
WOGmnxuW1Ym6SyQPLqlSVZUFWnRxbZP6yzI5hyQ0GUxrwxxCUqoZyi11iY2yKMBr
1W0x82ac5Y6Ps8WQl+jyYFhjAfNFY8qTfT/vJwCorb4jGMDFO6+eOmya/szZpE4K
GqX7Qfw+0C1O9q5eKSgfDEwdTaiETX6ZOqb9ldFIzcDivfMDUHPKwX42wvI8fX6w
sA1JLGHccc2RrVDD0MIJ2W/xzasuWEorlrToLFKJTJofNLw6r50xPB///E9mk5lq
C55dIOhG8hjUqsHr7KlF4RWC7kkQ8UwRSO5OMbC1gOLLrrkrYir6nrCXHCR4GfpA
WTuOhRuWjyCM/8HnhrKinSaJG7mzN7ICgxBKHJS9B+6xBQgFR4i5PuXWM++qDwCp
3O2/OS9USQE6kUKIy6AtquP6qsW91kcbBkt9wk+8UHt704XR+xiD19oKQJdHOLHz
CbeBGXav2MFFXigYQnndR65RkBkMiDpJXPgzcMTASgZDseiQu/1S2OXGzK8ARwKI
cZey54CF1ioVWVoK7DW6fZjS/EHdCF7h00eoh3cCdjCFbjanfdda7/hNpqTEAuNb
Sgg8tzHFTl31x8V8Dxm+F5ZeKJ1b59RTCgBWi4LoVPIsBKDUB6xGEUGOXwL7rKC8
Onw+vnljfn+FrgKEc+I/3+qdvOm7eLNP235u9isJz0KrhegJkuu914sm8B74ALZc
oszV+5c+ahoVYkNcZGfqsAGtyGBIcui75jkY3m8psXk/2WjvDN7E3MwGJgtTRskT
VVzIecq5IzVwNpEZGaH1t2sOlBRQ3DkrXMoLt7i7fZfpVVTHrtAfcYdJJbU0lbYV
8YJJAIT7QrU6kw8nBuvKMh0a1Nhvm0Q0SJ8Dt8shfMAjM0I4FOpK3fMZgt2vBx9Z
rQtChaB3CL1xZgyFdVgs+rIGkvIjM/CgPKu4QJ+oXF56yZoVN3sOqkfSpVM25XqK
ePEx6/MGFmX6rfCAo3jym8i38zVNLtqFOyMSEDQB3Pi2MAhEDxTjA+COfA77gk0m
3y5CY7vSk+tHnt0QKClAvdb8w/3vl211O3jOfS+YU7KekxKYF3ckzSPSBfWYiUDq
2q0GRRDyYoSUV/QMtO19BcWoeCOGZh4ea/QCWLqyA9UR6HZxFIH0CMBGjvzV7VU9
bd2n/4YrMkpxCmeJU6mrJsnDLDDwdEip1xg2IIs4XSeiceluvSJDEHjHJhEfUxGg
MZ3vGaxbYc8/dcI05TJeeOVtYM66VYzEtKmGD6JJiVYyNdlVeuUxmIjRgqLxNM5i
/z5xyWb9EiLXKheiVFgyy3gecEfg25Ko6BrdSzlA4A3BIbbIocC603RftvdCasXQ
YjFff21aeB2LosLXISd4CHib9JscKxrysaMNMPDjQarNqeq/ZNxL1Lu4qJreLhmk
eIoRd9k1k7WgaGJ9tbaox6NyAhcTPu9o6eK8MAMrl+411IYLSh/c7Uke+0DyHWRB
KNJAnFp8D7v/h2/zoN/mByXl+hYgOkU8T/yGhBYCce3EOxbpOHU72Rb7a0zHfN94
RHTuzwYXh3881OiknkDW2+tGP67VfPTXabPwuAPnZ13LrQxjyvC1Qz/zEUHG6W7f
W/yvjP0ASKerzLOWvcosSJMqpsMpqyypi2rKZQgYPrnRy1CiAhT/Y2pr2XZACxb/
TMb7Zw4fypkoBIJpbNZemoc+lJ1mDuMG6ycPFIjSZBG96AG6FWvR70s+ksvgEgfi
BcZk1cYqj/RW6GogRkuRWYkO+CnIiuguM9sZwhkPQJtwwlQrDjvc1g8FfI49Hszm
pqUGvPNpdN8Us/fS8mZEnUPeGxa/nMe780BM1WoX4kKpOPH4Q8AvjWdV1neIoqno
EayfQjOJ6XDKAATnIntpcD5VvTMIuQ0EMz5XTgN2Ob1bqVhc4ZWNL9XzWphdNrtK
7geNeegXpr2oCbTEFjW3HZNMmVv6gbTpouyRf6ICCw44r6Ki37COwxZdnPsQ3EYz
L70KizIYq1WFl0HvyeZExBYmI1rqUQd/+7Zutt1LU/vEPZQ7KeGKIAkK8EUNTnNZ
qbgt+q63X8It5pWGaXF2WREdnmqF6krF3YnK8ZsJSjbLLmr1cZIpn8jys5/V2uso
7ZRn1MX8+s/+dDWBzqSL5ans9sZgcYKmZyecT2fbJeGBw4pQG1CtxzEiZt0Tj/vk
BFw2aPsaj/1zJ66+Hd5sQ7PnI+WSXCbfvJ05k9E9LynIvfKaxxfwjnaG/BAruGyr
jOPr65tsvj1FJpZP1oQQE8LixbG9xeqnXmNZf0I2YsYmhgPLxKjaozuo+lv8hyAX
NlQ4EOgsWxqffHCMyXUnan0cAInWO3rhH7YiOCYdcOQybUjfJnMKzjOyxDqiWl20
g/XBAJ/YUpHmGtaHxOHu2+GIYBcNS8LpI1pxVVjzwMCu9ZyydBf6yAC08riNJCMC
hJRsQCIgdk4aD6h9Rz3FThr6CwR3P9PNnfB4fkB7wv6W43Z2fUicGq2KWIOruCPo
VTF5/1ysbyjLVSUa7KYhROita7j7gY6fdIPIp6qYLCjqfwtA19UsD9f2wRwx1wX5
btPSEFNWYxBUUoG1uYKQXqCV/chBodAq3TQNw3J4hiYenAu0EujRBjIw0W/aPZyS
48zmfqRFSXLcGg79bgx+Em/KU1C8Ddy/tscqDOEreJlAMeyYGId21ETciR96rjGS
3hyTKpKp3MI1DMUFIaQS/cQQ6aHmC22sMAFC9uj3h4865U7KBD2MXVsK/s7DD7ZM
TJruO1F1t1JvoEIUKbmU+fuUX9WDfWLr3JrngZxow1a4c4xY+gBFgP9U8UThLOYe
ZqZMk2NnCtQDqH2PsAeBxJCQAM5qCp3Gr3vTax51TjApN7h0Z490WzPf0X86rEou
1LAeMT0TicsaXlBbNNe/STbdFcWNRSU4SlxQfh7BlhkfBV2kSbKjy6M3yvcuFMlI
1gqD8Eg4HTEYDhQYcVBUOqG8QntozN3wl9skpzcQFhrLgya7AzQSMB+B1oCS5CH1
1AJZpyD4I1VruwOC8/bCcbepNJiQ0M4i08j7TgkmEplWtlEA4jg+VanGY1N4PZU5
BjU4vCNwZEDh8q+Dk8JFWGWDEZHlU4n8ksD+c56Rt878DAdZJsbhHv+PNHF3Q2sG
+nb9Tlf4zhmrJ3W6b/jAswz0oLTnViDBRTYlEwJUuI63+ho93aSA8lbLwJE2aIad
a6fDrdgiXFNNo7IZvEUd5kRYf8zSJ0cIpeWMm6MywvKa/+Kgqp5tCcGZEAzpBYOv
JK8RRyPLsflBsZArkVRC8cbNqYGXsz1XRL0Qg2QH9VJk2Es7BpH8zXjI+6wPaXzC
TZxfl7LYu9SXBBbuRTy/KWOhLISi/xOS5new9BgVi1p/O8eSVU+lYc+/Jf/8Xbvw
IgdbnHpFN+um15gQQsPhP20Isa2eHPxPWobEJnXwaZbBBj9Ygea0uxqwN/qVa+If
1N3DzkfxeekJOeBN6I2VnSIo6Q+tP3Fb3+dkR/vPSFn+NRfFGZZQHTkktKHzG+mG
ssvWU+wCumXEcpxaglq+7vaSsoLncjOYrmhQWqfM1oRdfCs1m0MfyHKDeAvZeUAk
Ol24SBo//ov7+1BjcTDU/wTotNi74ubwyK1kWWE7TTIWsBYN0yDUpj4VP6uJrhWp
iG0rjtwjLhqQ51PCeSh8fqzTlepfdzFwNiYJ+zn/ejsTGaSMK05wQyYwKzuraPno
QBHDE7e1uK1+J/BTccpVXtF3mXVZd+ZRNEiKLkQi+T1AeOJaS41BjWG8CWIuMjW/
YRQ1P45Fl+H6DkbvoklG6xdBfcTMRjfWYNhwyGThNiMy2yIq/61ffd8AKM+flxkn
BdrBLGlGHxM8jo16Xv5L20856JZEHArs04dTwV0FPt5m9LVQ2TY2IbhKF5fhBCxi
lHwg8aaF1VzKk1qqeOmuc7YC+mn/PwxMrXJz/5029PPl1LJgQQyhtVOsY4dX+PB0
glD7qSA1EsYN5eqa2UcGrC7Kwz7y5XPUyuxxykxZfvUJPZ/xSD6a+lQkOWqZunBT
cJTjOpHp81Zq1zJyd/QiZYZQrk1FIEXZBhwL+UnUrDpu0Nohy5U5sF9rGwdT/DI7
uflaXnvWxoiTQWfThyJ6ewwWH9nVUv/gKb55pCNxUXefG1ZMI8t+Xw+I70wkqql6
f4WoZ1y82FgESVG7rPoZREGl6tdPe56tKSVqAcAY4fAqoY/yvjfRtDePVvIQ4sQY
lIKqgoM7WKJG8TibjVRNDybhin5su7M389E2w2gdFZ4DiK7ZitYIzmXH55fXbQY2
xEXIAMY2tOHGOXGuRh7w8bwsRaUH947yAuNHzKu/earNnFatLOM9yDiH/7KmQ2gi
DczvAXSNwcxOKtRHtUhAvRTc0PR6lwUmLsk8UIxOgfzEeqnlY0globmFkeP6W4xR
qcHj3wWW+/QzTiwLzZr+5Nv+krYMdZAMmw06iMbeM6GFGHX+xCCsoGxBSN/5XK5h
O9jcuKf2KoXzjyn1ERR7VEgmzFnP744Uc0n4PNSKSN1sFU6ImJzrzHbjVBJa2IY1
ZRVMjcpNQy5BWu0omGyeAubjw37fYNrZC95T2lc2FKixtyDXdRbvsMjTEoEkUyL+
VFMifmdj5pTO1B+QTE1+Ju1m5Ry30dtxlkkjQ6xxDT1MjQ8lxisHu9wB60HbygGt
Ef8IvZN0NDIZ45ZztBJrnypuIymiVowx/iud+EtsTNGe/21vG+OB8rzGcyo/SPW1
uLwT4vcIN5/L6Xd2vWlkZHHtTFc7dIVuwYZrhhgEfikTrcHQ0oQ4eKhe5cJJc1WZ
mVbAq3H4EIIGPzpNt7OosgSE9xbvup9MdiyPBe5ayEVot1UOUa9B/0u0vEhpwYtv
m6BrhsUqO/3fL06mg27A86XNs2UDHhrYxm488Q9OmE7pJ+LTeLRY9a/fM5ohcCUF
QpzPHKa67YV4hM714fOZ+4as38B7RFJqJ+cgII4TOYgBg7/el/fvD3nogSIjMrSl
fjIAJ74+jSn0sqqB912QJmE7Mo0AjOm0cv+ovf9EaLEqJ/TQ8AOS89DZtQy3I4J7
ve7TxYmAT4K3y7YdMCpDjTFKK2wT6ZiVlwBcFIgXROkIebdLy1P+/TphUAD8fXS6
1e7C6onCFA2zkWPX65qRTGJ/WjuzAeqW9ooBJqfrXdodAT7MibAzox9Q+LUHVjum
MP8tM0UD1wqyg7OxYBHuTMAl+y9pfUkoC+oYtPDPlo6+/R/8C//j7rhvyuoKwx3E
pBdJT5Pe3DWdgWxQfcJl+Qwt9NWoqDVm+7s3kBsD8/QQj2XHT6PWBTWx4nIHsTpH
nzzHMhhCaQbfwoe8B8LN4F1umPF6b297Ks5tKVH1Cg/Q/zdWHV+yjG2wICyb4vON
5hF7wX1oeC8+ki8oQIhtkp8LbmCFYbLUR0Y/MqHM05A0A7dI4NKDaL+tpF3H/oZ5
I6+rHCY29wau6kMOl1JJjS+V9Vn8SqLc9hW8zI6WVVGI+AUL7Z++pdth3TbUtwvl
yWfNSdFxggzuFgSHAzN4be3E+ad14mLZWwS1kqWyqw/kAQAx9CYM8vpI1xgAgcVQ
syrdtn+M68ou4RTnRRJP74YXfqqQ4dHp0TfIRvxJNsxg93MT6XX/lBNVbaPlxBhb
PRdAJtjUXj3h24xTNkLHBG8dPy74EHSphIA3t27wmNnAXXJdr6FHwtKXAzX72Zqj
4HJnW5U+L9C6/5PqYIyVtmweRzfuF++jkUzjFMoaMM5/iWcRHfIckbD0yUeGzIMS
ApIXhdqTg3XZfCC9fnDvOMP71kOdJ8SadZ1Urvx4iXcB67GnVRghe8fhupXFKcxM
a4luvebTHouzsL4A8xZQS6Z/NkN0FFVhdcfA4zKKE7F14kOM/ix8ppo/nvzijhAG
bEWChDLQ/B/Dsn0vS22/SFNh1R1Cc7NsSdUB/s0D3IrXa0A5nYYi+WTjQRGLSR+7
9NzQ+y7Qtmwz5KkEnqOEohgQd49Xu1DdqUR9iQ9xOcioNZqunsBUoTxGEhjEFlkJ
tEP0V/3beWqu69QDdkHCRHTb3TExaSIm5WEAHAr3DjYAMIIioVXPIYRalHpcRueu
i/eH0+ZSy5+frc3jiPgYgOSbsUR0ea+AFAuD7GmJ0Qu+uzTz2yM3gEs/xZFSbT/6
g9eEp5pBfyzSQ4qYXEwQ1o3F0IG7Dvuh713LPvkE/1gF42KB7ajs8gOUva/0gmEn
p5vnnoqNv8g7m88G5MrnbHhGl5syrAoop/M5ecoqB9fQcFAITNuCXavHUo3f3eS2
ik3lYESjlEPa2EQOXyQs2af5KvgxHLMF+FnJvr0LvkDlyHpbqhSHqUf3g8UWc1Sg
IDAYe7Fwt1L7dupQMUe878puN9v90xNYs0oMfeU4TfBWwEmYGZQNIgTo4RZcztSw
ftHPgEWwfCgdZmizSGL3bwo7te5C5dOK75CJQyqpailE4/F2GsK6+3lkzrWrDm9z
s6FTdsfmpjESI9/r2txcjdT9OerfjzMXkgk6HT6rFesDxh26tfIqLx509bajdRtD
Fm7eETVvBzYlfxsYeVLki95+/H82+SoNtM3w8BTll1zawKBIkzw8NDS1MpuRHFdo
MQu9N/Ki2Gggneqxm7bWSZjrIAIwbzO1s1qtBNcGt9X3LWZ9UIB4Qn4bUTplKdKw
3Tg/NhorUK6Inu/gL+F8f29X4W17NywtNCPk2RehoklTDLuorjphY30ZysdRvv7k
GWm6xTTlhHEZQaMyqCjFHQA0Vi27xI23ubwG/OaKBf9YpncJ+rQZH9DByDSa9WxX
NhNzboqyoADfq3PZRiquT4t76naYF2mCf8596pnHbon38nC/7WC6/15gMq78++b+
vbvNagH/eI8nHWURraKnmSm/UwS7y2pzMiCjP9GBeDlTAo7YZAlsooTfIyWUQEza
PaUctc61UaDF/hczvmIOa/2STxR1Oz0Gb7X5pcsuWLZ5nFUXH9kPHhCq6sEMMUdY
Zz2GndNm4vC6W6zIirGaCcT4NT4Gk6ZwE70prbXgAa5W1RKPDfAi6AF4/SP9RzjZ
wZU3wkEjsFVSW0glPRlXtx9Tw9GJezSQaEybt6JIZx8wuyaZPy4txkJXyJt9PheB
6SqvsjRDBVHnO3RV3XDLVzxLCHWpPtL+EuyIDSfFwvxtCqVfLamC+k+fD7luttOM
JOCBfF+Vlsm8aeFCArGR3RqY3leOxuKw3zIQMBOXMfx65lREEC9jPs9+EJ43/U3x
RosFCt2VJe24pXDMymnOaDyc0Yi7fBOH7NI/RbDCHacuNIcYxgDHKJGWqIR6ifqB
GHBnz0S/Xk4u+LiVez/6gqxN5sGJ2jgaz8py3xQB2bhiE0fgnUHyE2/zSn6HeDfe
O3xoRJXGwYmcuyWM4a/FbzRe95wjcX+58T27HukNNECISFzX5rxOwGse8cj7bVoI
BubzGmaCbwvs+fZp5WKWmbysdzYMkPS2whfo6t9NCQzaq9LESVW7Y78n1tClZXO6
ZjMeMPRcCMtCkW9PKDFgL7mLz0TdYDOf71ZiE4VNwKI7L47Cc5p293Jv+ny+gWbH
eiMYPuBr1LloPjwdZoAr560qFqJI4b37YiznB4hobsZ8I01vkpt0dEQ6m/7OTaKz
nfwAc8VgrfPWNAAuxfBpEVxHdrP65sZkO588xwza7wPOo+5Rmy/l3HORhczJamAl
NXi+BdcUSq/zBeqTxSNA4DendfzZ6bPBpEylHvDSka1USZvBu8qlekQOGZ0RowvQ
bx/Tc3rHvAsSKZP8fcDEjbbOV3xIimUsMH+El+c0+NL3Rq21tpoHOLWZmmeZY5xO
BVrvlbBzgTLnWMZGbqwQssUFPNChZtO76xEl5FfGeeOC4arahCfd/oq/5h5lmW8e
AX4j6E/UbwYDHgrFpDVGy1JE7MbyKuA8BYAx4qLbyq93sWd+K3S/zVjKb9f5hv1j
MwTZBbo4RXjNNuOqbeFfDAfgkYEkvemPYH1Bm0vmHKatZRBrR/DSqKYpzRMfQpNg
HlsUYXcLD1WzsdOrYTTvtUFRVeTgCPdo1zFdkB3GHzpmYj2iSUaFRJpkxEsoh59+
sdmWjhPBQCd/6xzJ5XA47eEMCdSWzrzTUw9/Qmf1qC5kzfdw5R3AKGiXM4VWsTm5
nmNEZIiJBaIGWjjs09XoCDmKg/J8sZCQNQ3IR7cXkKeiiDo8/3ziKKcLu5SLi6J7
JcTFQT5jRPSjJMUkk+vGc/yGvEt35hzkDpGgUPxR8eZoN3FHWNFRDU/AeLLw6O8Z
o/Thz1B/cqX7ALm9SypdYPC6yCG15qLnzYH8Rbz3lr26I2gLlNgxGwvPn0n8Zy9M
QHBj/UU4D01e4ERt3Ootj+lvdAl+0hucVMZCgZ9QqSpb8l6MLaSJifsFFT2Z+uIc
n0hEXHyXSjCh/4omrpvv7ZdH+upcASLI7tZs6Br63LdIOauEciZ/Hmaaml+p0rgV
81x9agn+oS99nJLJeE8hKD/yaCJJ/2WnhvyhRJ0mv/JtbMhU79he12GrKlWz/YKe
wJBrFQZKrtrX6OQYIHrWQ11mDQZGB43gX7CrC8KuGEY7VCrZ6kb4bk9hhf6XKZaz
WBoIGprYRmmHROn7uKw2WCdLosh7R0VwzcNX048B2R0XfoWVm7PWmBqMdURIOGxa
bwzVAj8h+uefty7iRzuaCoOmRni9RUtwwod1T4Ywc6Yzkw4DocJDfMjGfyNjUX35
BwHJlnc3Z48S5CYBVoKDEZXxOtRMNz/nTQKxMEhi/l5B3a7mfhGDnq0XIuWxM4pg
u4/hFHCRk63afq/zh7h6VRs8lJmbb2uIDWzAtSEmfysURGOiT2hi+y1gJGz9Mnk7
/uEANeACDfG6kcF88s69N5zcEQ1fDpl0xfJ3aXLwxdxGFrTO8mgukfp93UazO+Lv
gZgKh+93EDcuLsxPNQXKll5CjSyjBwG3LDzLWz52gL0ojJl9IGwDkjeozwz7UN3/
gosPBJd7bZpGMW3S8tA2oKnEsS+1peWzKmd1LHcAzdgoo2y9nFFX78V+mGS3RV5E
+Qya12c/y3ZAdM43w066rZpZwx6PRj1UH5niKQJ4ns2AVekoYMhGnPqWLovNVZ5V
lslxxCXIq7J/hcJDL3liPLmoZQ9vvdyQgvCxqH5n3p8QpSZlDucwNzqRKv9L8E5d
HjUBOu0nYHks5iI0uTLtcoqEM/uvf9dR/W/7ztM//ou+Jz7tdndXwWoROXKrjFxF
oIJmJye3iQTacCTCePgeIDbskk5aPiWuiPpf8avgjMJ6YrJom6HtqXxUYY9rYDIM
qclU/zB+tR5w6FsdbweA7nOiUbWKS9IkE1RDu6TryPM+a3FLiKy7TwUY+xE9ho9N
cYLS3ibm2MY97++r+cnjg/PeympcyrOZrIRfOsfqiYvlHQMzk1MZMJ37sCGmqAO+
568cw1uAZI8tunXxnYNn3Oi4M1TeO4onr42TgWvptkHe6WuGozsbXStMqJSi4D8o
JEbJn0AkI+KBdxu9D0yGKT2kZO+Xmr8tqPQrR5mfZJJyzA9uL0xjmdi1qH+F8P5L
Yaslt0SzbbhO3dw004OByS6sxNgK4QVsIG0f1nFtEqipTbXMtpsXuuorvnI+8REu
A1OQgsVfD1XZlZDy5Io5Jx8p9bFYh6j2Bb6hwf2DFGAVckEbJWeM9smm26uOvJNX
BGAIt5kOgw6hDtHun3xmmNUW8Kru5pBbKDUxY7BU15iCl+fVE+C7Gd604nN2TiFG
3sTKScO7/wvsAiwQ+Zw64458EbcltSzYlfPzJIG9sOgybZz7+9Tk8suNdB2aZ573
D4seQMhH6l9pTf1vUo4oWHAn+8u5ORHlDCSkkOiMV3w3ocCHEiXfRseA/FawIu90
FAMGTB+RawBzZVp0jJJ76tLjiqUXtCraf5s+K69QdQvs9EhjDDCHLao1b0tTHPXm
zClvE4uQsEtc3jNE/bwXTuvCcdXejDklkDfV76P+IbFIZzBnrnaT3rzWT+DjwOfH
K5Yb3Mvecf9Xf/o3x2xd49K9S/pdifn9/I//ztknBCiA7+OFpbVfL2yLE5n2MBwl
yzYF2G/7Uuej96jJlAbhdb90jnZFSwSNg4By0T0TS6xmtc/j3usQ57yvE+BmhRTb
YO8hvzBxFtisfxnowiy470EKs6AwzwHCktcvLtaaBwWYMoEYfF0t86b2fIsJKaf4
q23p5WCc02EExdg3yuPQrYxccyHaypn2CB2TqBu8O3KT/7umtlSY/FPj6TOa8Im6
WybyHZ6EYFZODYCqc3n60JSECogR9KzYwypdJGJlQMn74aYUtcIvj2gWeAfPV+mK
KMMqSA/rbdBVwz+G/Q7UkA4DzbRMiBZw3t4dGRY4AEKGkuYhz+Aj+EN5Y1sBba4E
0GWDDBC3vFfDz1OoI3KuwTPiwGbijwKefn74F4MRwu8nQRvSZUePVP8JeY+S/h7X
fOSXWuHhf9u4hY4IlE6K00Pu9lzCRbakeAaIbU7GEoqaMm/rsZozwrLMOvt8MIFT
KTiYZeuypG1qAU0ymN19q/govQN3GG/TfyWSusg0gzSxPwSOQwR5xMhedNbPLiiB
Yp/1TTnYEB3grD6YQqN1HJLeA88ksmjUtJL5hdlnNrDnFAhwhPHjxA+hrWHaBL6S
Ueba88U08EWWx4KPMLm9/x8ElIEyDUb69eJrgSYAkQ3jUUAhUIDH0rZtyLc3a+VV
HvF1qlmPL1bMtCMYUlIUQPjpCMYnljXKOtNcKVnOOK/lCzJmxex+EkopGeUOL/Yq
Dkro2pS9Ugr/UeuF6LZksLRuV7WHq16jqrOBJzMO7PZbw+yitWBRKK9KS9V9ZuOq
u7AIa3kbrQURT89E1XI7dc4tVqrowMkmoHewdY1XBgCNs2vMyarD4eXu82YgTthw
wLHPdo8VgAFaIk87F9mgHQcsZLzU3dNcofGuwIgX2BMtHtFFK6ZFygr2w+7WaeoA
20T3JsEwlpjrLuoOsD8/QbVfBUstLmpiy3kc6f72FDIF75CTEHuxxBWGfY5pGyMO
hxhf6ulZBOehfGkjs92GIQFQCI2J1dArT6K4h23F8bY4NvNsLAu83syvXnwyFYrT
zlc/SxBbhAk7Af6Oi9iIaaVQ0bCcx29U2wYq4dNlfMNfoIxLPdTWmnwRdYE2Ah0f
zGebQ+3rPIpkzmg4cmAcxCdy2ijyh28UBgTtRws3FL7ArBAkmZDvV1HJm4+73rYH
pGTlECt5I2P708uG/po7cLJaSUMpfMUtgJO0VKKnR4LGdgQ75jCwFgdz5P6A6xaf
XXXuo3dZ7JDjuSG1CBUXWbu1mtEnkKeGd7mzoIdqapOAcGypQdYCH/ir1ViiVmcW
gTDUwI9aclOXQlayUzvM0u68Ar14lyz695nSQ8UsnnSGqFeHXPvwlPlDZLJyWypi
K/8BmLStkbfhPqv6LNK2fk6QxjW0oZuhs5Pa/koTtyMV9ENOaDDd/mMF6MvFMyqM
VutsOT3g4UsDdhR9e9K9dl4wTGe0Djno7envfDQa/oDE6LPzE+Z2HfCUZlpwYW/+
H23hZybFB/szRod6C7dI+kg1AWi3iXgkCPGcjQ9SNHTD/vQ39Gr9pbMaFyTrcDIA
j5ryheXPK4TTtBBz2mq7BPMVt0K78/qt0sqTL+lMRLwCljiezodQNSpcfP6Jq+9c
1QjFIKdTOPRbiSdcUK5ahN2UmCFzStr1efkw0pRbImbK7C+ajSCpY4bPT9dPxi0X
vX7Jy6bXrE/rR7r0PC2MFAL0hxp7UJwGqVtzmsDBOdTkYdx3CcDbiLGbTH3psyOg
7aWmJbqHmpI6vohSlVesOHIF+U/X+t4MDKOEdxRklqhP7ueHxMJDniV0mCBSaQ8l
FNN6jwPW8rXW1n3/X4N4mJkBTMwHTJtwo0gXLDduM8T2Aur/FW8s6rengs/KArM6
nhjuwiRgS/9cNh+yTPYBh1JRIaX/VoUaPkV9fvPKKT9fm5TxcI+VOU4hk2gfNAAw
ChK8tQUy6HeVrr738C3FbzUoxOcwPmwe/6OjrDVxn5x7jv9IHZguReKIn3ZpMsn6
ICpMwoqPo5aW6Ks0Gu2x/g3SjEJWYPbA1m8+mpXdr+9+WXwCnjgVfDvfUZAwPqjn
vaQaks+nrU1/4JEQIqlYY97aulS3rMw32ECyTqlakSGcr7J2MzzL0+vNqLzqaCqF
l/Un1XB2ERqKGLCYo/J0Jk/sJkUNkE87Fbt9fKk5mTH+CV+Dnq9WGaeSVg7PZgQt
aiyT9iS5iOEe40QW3DpmW4BGVxItLb0TctvjF3ZWxpAyL1pb3NmMYZMSR2QuNp+m
8dqsdJQ67bbqfFNmP34sIu2TNxXWigaNljWE+cMI8Nbx2/Ylvff9lQCrvHHNsIpg
U6QhiDLsr2pMjAT5aFnQQSAJf63gCpK3PBgwT+ZivIeDUrhNB28RbfCuolJfJoIr
UdKd4I4VrSeBsJd/WlQ/vQDqsQPYFVnfLUjzI59VJ9sSIKmuJ1BBHv7s+0810BD2
lpIrn8vQEUgDx+VxNEUcZn+nZiTUxFHhwlRYRVsteo/bfcj5MV42YCsen3AXccDA
zO7oKjlEY4HJs/BrKNfXoEgZfVohxpg7OeI5tPpjOpenfKlYxPOaUG9sotkXVDkv
RSxdAncUpVDVdDTLbd5UG2mC2eFCsuqEwbLtJ8b2CTSh3HkC63AFnvLySiTsQiK6
oPJxEj6EyZ/PMKC1CByTPc+Albhi7+b2+tqplESYXwa0HjGJSQ+pYjxPR8/bL94W
D01y12dgK0KU/sE0aze0dSXcyrSN4a4Q06AlTFMA+VH6KnagPmbmeEeQlDI7dAR9
iJOPKXV+72hZhmitMyoyhHnIelfRxXa4Hup85EEKm57PUKZNB3X35KHggrOa+hYp
ZRkzwlsyQnPa+LeSqHoo42RzWkvOBYEkPCBIOj9o6wGPqyIoGK2z16guVfLXbSLi
mg5a0nPqQBvddetC2H4edo6XotxG6mRy6jNOdCWF8bkCQl34QpD3DnlZRcE2Ucli
mwQI6gggsqOzUzfAVtTwWHbinQRo0nHYkOB++Ocwxd/mtY8uhg7qalRjhDo2vXbk
Ato8JftTxwXXHvFFdaEP1OAjoYRqNm3VOB2U0e+WPasLGgeYA/TLYM3546ud1n6G
sieZWXwY/KsxjRs2eue64OAiJBrhqsjz/TGwISEUu3z5mR8yI6lJKEUJuokcn21S
1FwTrqGVtUodm7ZQp+fTw0i/XQg3kK3+yj0WI0bTr81onQgUJJhLSwhtGTDTa4m3
48trndwjZC+PMxLd008KidEJG22lJYADE5ar4WDQl+IWU5Uag7r1fJqKGfJ2QXt/
uy4DglVyWN2dxW3fIPj7BnhuIqHLRbv9yrzWy/9jX7TSX56gcrYWdpvBkZ9cwsMz
mlu2CKRjTMa51BrX8/4YDWDw37DDdYj5kM7k0Y4QduygWqBnrJ4o9bJg1ea3kUqh
X/MASMRe684huAjD/YlLDh5pvKuN49JCLKOsy8c+5+1KCZW253VLZ0s7sGY8rCCl
olNdqiLdiTfF+Dbw4Z8h8TzCXjsJGW09lSn/IN+W/+tDps1UmnyWJJKacrnGYPOx
d7IojYLx30CcCjLMZxurbkr//r4Dh/4ha814TsI9lc1Su396+KId0GACwVyeNl/o
vnY1K7fjEy/vz6A38RabHf+HvTt2dFUbL5B4PckMKZiOhOKOgeBiPsY7lhgCNO4/
lJKiodCNNxuG/slNLtTkw3tLgrnBCvHwNyd+LU+xE9DYzk4Oqy/a/vkTC75pgAO4
etxVBKmHqMX3Ybs4yYLmP6GVl8yG1+G0vauWQzi5YGZR6YasyfkUVdjEmNCrg7KN
Nz6098rPuKMHUXZF4hqESz2xQfZBapwQwgGAOnFthRzxHluFY1s1miey+sSOQXaw
PCahQDpz44HwED+ongBw6IpOEQ9O3LaQsVsjYaTmFoYvdk2qkixQYG/TYjzQ/cPC
ov+lGYTvtZnykTdCmaELFMvmlgskYRpExnXaBFEyFK/LUhBwHHmbUH2UT31vyPuV
cvpyjvb7nOFZrYqfO3buvtsWVZsjwSrV1gWs5+F0GG6d/KkrAa1n/KVktxeLfo8H
FXQamWwUTWTBmFmjnSlSBs8WOixMkrLPMcsdpVz7HFFZPtnFoKOh/NwWUSJmckrM
w1qwazWt86EOKz3A3webzHJZgZwau9fs2goOq50D/sMZyacIuiFUE5l1LWuFKPW1
G1th3FyPxmLSzNSyUGGiIeQMUoEIx1i3AybTMFdtwGe/SwRsZQ0p+5YMfdJC0JuB
/yG9HSv664GyVSWHX2eG1Z6yxYWmOS8YUK/IWMJLjhvxolCiNqOFCXQDm3oGcrrn
8/IfPlNXq10A4eSJZ3NQzoB/9Bsf5TxK5vs+7TxKghnQ1Q5T306JKcYoM1pWTOtR
c7yMVgi5AgTWOXG9kcq2zzUPD9R1+JK3QLbN9fmn77cN6boT4S0ws2E1p8ooWS6o
GtMeVKG6oePZisMdx0RrTmZXGCyI0daQ+vHoUhuvymVGlD6vVr4rhMaSiej33bwh
mQozjeZw6O1KN4lxKtAa6rE+iK0kEAQ87Yx/knlUy4CyukGpmn92T0k4MoT8D9gy
yMMMXWApvropGTofgv2OtOjpidXjGsbcC3LOVlxpXBwtnLkNI9cG/A22giDuQv/8
y0Q4BiSZm+jV1SBkNJKz6ZE+QeLAxbBW+CE8cvXCL7E+lwn8rJRoQ++vK4OZfTZl
+D1a3MwN209P1dLBAOBpC923XiSBMG95dY26DGulgUFZ+n7AxoO3tlkDupvP1N5p
GnRivyslTr2RmXK7DMWT14BQqy+C/LcIao6hSl+PX2JhbqKjRjL1BySiG4SvNaPW
SLHbI+UW71mSJ/fX+5LI8cJ4ZHHJLSEa8ZT2mFskOLtVEti6Fmlg+LSs39mn5lSX
nWQMXDbnDw76S3emz0Z5blUC6CBGktxjnvYWmVvJj8yKWy/N6LE5r0XJ1mUA71Vm
BLH4RZTa/3Syo+SRJwbcSAuoQ2hEFURaUAnKnaf9tLUrRZj6ykHkyNHlz1cPUTwp
4JeJ/qivmMXmaPiLZvaPMDnBJ2McGNdpsSvrymKZxJef2aofV1ENMjiVOq/xtEXU
iHMVufB7Yn/c+zhog/FVFsx9c9y4R8aYspJVoSNkHlovcI6/IolOFxxQtKhBPNl/
ZyZZ0QhhMvYE1hELO2TFiwuVH5C3LXsKKn+acmIoRCiTtZbzQ9v9TZzeAF0Lulby
9Pe8yCxhNjupY17Ue8I+4oGU2CXE1mnY7Sm75zt5aIYMUGPSg/ygDo3m0kkitR2K
GYIactJD9CRWRFnNibcjyl9wbuzud+E+763RqMhr55ZZFdubyKkB0wu1K/OvwIQP
24y0+dhwQWQIjd4Bqrwk8mh8pzFuy5OkE+VZzmnjqyAWubH05o5U/ruJ0jdiCWE3
+b7jnajURKxbQnxyJuzUudBGAT8JLnJKPeJCq8d/GTHFvgZypRX5YfE5GUlp91kH
ev+u/OHCQcOi+gleL842wGTUkRrJRNW1j3AOvnP7Oanuyo+7dm/tzEOguKqe5uXD
E+HYnFeAKs3bM36h77b4IfbrUMjdssF9SBIBDgGsNtJux93qZlMtDXS/jpRN3PVd
mVF4/ONOAPqHKcd6Wf8U1fQgher/MjY7Z8hlFElOe3/yusY68DQx7XSGW1qOBXxB
xGbMPiAjYKg787LJX/CeStbOZK47u5CMBvn13rVnXwPJdKejH1yuB8zfoedbTAQz
riVqAFIMIVEqnNNEViUAtjJKy1lMDNfZJNxjMXWqpxveTsVTLuF2hRJxndBGMfcD
Z+qM0A6IMN04+RLMjEtIjmEA3ECBKLIet+NMaYmOWk36oUjjmm8h2CMqT8plDlsi
jZz+1zrK+Wjv2mKmivip3Mk3i3qrLAeeXvOhlyMsS2l04fBA8Fj4L/LFEn6E36EJ
XaB/DKXfXVjOTrIGuQ1oH5zBfMGwQkKFXUq9GdFcrC/y+YZOi+tZsBWomUYVbfi8
eRVNHsBXFZbsxixKYbJJ2EYX/FYjHCjEpYbBwzts+KUpZT9ESJeE5DJNhkXWfXa0
rxoWftaZl2i5AQ691zllccEAVfQwW2Ek2aIenH2hHWfHNGdAWeYzrsGPfAP7mPO8
Kk96bafLWK2zqDsPMzGcYyEgIG4HaRmjBGPF6S39MxyytqhVirlLQOeNAUAQdM2c
tTF+aHBN1dd8C1SL2jmSRosr9AOJCQ+8XLvHev0n3rVKeuTpJA2lZpN2wbwq1QZ0
h4WdkiHJsL4bZLGkPABEPpv7hAPKchz6vgHPTQq6aPEISdDT69BYGWxx5cpS2xh/
N9q9N1hnTybCn1A+TXhEEZ9FJjmGtCBRVV07CNK7Yz5mKRwCefo/VmJ7F4bcpNdy
84spd1sKkf6zbGycsIo7MVlDhSt2bRr+RECcKtElOInd6cajRGtEXmv+An5C9eCM
oU1Dk1b41mfr9P2VVKMmcb5PZPfuRwN2Xm30WT1h67mMZzKADqOh91EQqJO9HiZC
eTBK+wwX+6bNiUu2frPu8lp9GnHn07UeRHDjK3kP4ze9JQvQifm/Gjx9RYFtgy/L
ASw5EE762G3Gg1QympE4B222H3fzjqYu/16TsOdPdQlW+JVxUem0eAwb7VZQNEy9
6NuBofnYbFRskK+QBtuhhMxXWjAdw2v5MWvoQkbMeLHH9zrYr9n80boW9JdQcHuN
EEZjgYiT0AaNBNoylGNgFTyAcRpL6E5WIrEp6Z6fqBgLNFuCFAtWQQf3wD87YHyi
MTFpr+nFWLfeLdkuEVwJ5t3pgWfpynJSHRtuBjwEu3bxejZNfrthWpAZhldtUpBq
ty8BNnag1S+y1r7fwxziaAEb0KOZDaQ264OBbUhR4x0WlUyjdck00ugve6epEwSC
J812myXKBfz+xUrYu65z6xkX0eANxdnf2nGk8h7d8+7nC0CBiAoWtPyDcbqQcpjU
Jbz+X11WoiEIJik7Yc9Agb5b2bWE7uOyE2FDtm3E02ktZ3sraLgamCpaLuh8+ftk
eLVurLcE58VOwivrjRsP1UhLo323pAYZF/0FRbd9dLkHM/5qKbKwiDtzPweKj9BL
DHLR2i/djo/TXSkviWT6ufrNlQnSW3yRiR+OjYh+xeKPcsjxra2qhQe++I/XSLgs
jNOOedYAndZfrbKhsW7BEu+2XOqNf2tmkVMxp2abiBDpuAXWfMnf9s20lkttelVp
ZB2KUG1NiVdOES+jxhDbcuLUmtLZNSI4UL4Qzt4AnYiDlKqoGTWNPaWIFKEHC48O
v6YfVnhodxbQ28m0hZHXG5GuZc7umt6b12ecNoLsM39Z65YVRQoK776RCxTppHCL
WmWI/I9lhhJ4WgaGzzoLg0alg2hN83r0oqv17pWk8EiGnZNGvIvh0j50VMwsINwD
GixgNoFRYnPx2Uw1WPCjQ6dX+QzlpWpM03opT5BFcsLxjog8Bokew3WG54lETRha
T/PwZGYA5iil/2iUpmmJrLTx5Ug8+NLlOBZGveLTa9+GY4kIGa9CHHzfaswzIxj2
eEqyZab+184pmGJrz3QzUiyTDm+UeJD66Xe+sV2vTngNxFfqr3uwIP7AE0CGfmxt
G75kylrxzR+tEvP3yxkkfUtkk685OFRydQYON1+xkzO2HUP0VZYxB0tA/Dim6uLA
36kBPOogqJkVpIBzIs1CRneBg+zhXWWKfkoAzwtDyaTTOLj5df9wl74MBEoHqXVA
4V3+LXiosyx5sblZ7GFBBPuZRnlYZCeruGh9S8MGs/SAM3QGbABCPZqdN6Zkz6AK
J05i8co4lA7enBLgEuty5SKEpig8Bx57cAPlEWhprH8FTWB0+UOsrNbIFemsc04z
+u+2PvF/lk66iNK4F+pZPbN9mmGAp/GhWKd0F2SlkKm6muzrtCSbS+dz9VMsoCR3
LlUXhVAJluL1rEux9YFuzQXeWOcOoZuYgA5vzZDJ2lapnEFH+kcetJaGl44472BK
1emcUI2Ndo350w9ZQeYD7IHkfaGJS7waHzFUUI196Ro8kWexpj2nqjYNiiR+chPo
e2wAToIMIY9eJjqTJqVEqmMfXv3aWjBaDO3o2MmujD+Jzojf5ZG14Rtcd3L4Eu8H
gNS6mIaXNS69b9XFbdZ4WmrdbGsnVXalseUJb3aJIRKNP2se+CgQH6o+44UQXXzk
YZP9FO/ETlle+vd0Zl7+7J6sfJiA1Oz+v6pf2WRkqOoPeRqRvOiYO7KFVZiksd7S
d8dwy6Wj/gRZwKI1yZZkm/DDikolc7MGHAeCNCCA+2Bz+YF1haAkdQYemoSoWTQN
uU1diMruWOqGtB74TJUZgNAyMhyciW8C460HZetEmZKrc/dnLbpDCtZLLkZJiZpp
OhhBgPOiAgU8xbWsa8koQCwNR6yOxAIYFOo1SvArKLLI1z0FTwqtHZHRM1s4INn8
64httXwPjOJLM2vDccOgnTAIqumz0A6e61noEk1Wna9O42sTR73n6o+JyCqwB7hD
OwikvPyXjYWQIsIxszR1US8ZQTxXGF24YBMZG6zi6ddo7SY+LnvN5jbcNEovebHc
xrX7ecv+yeDQyvPNvM+HdSog+9aEPXdrn7HPrt4L91J+r2mxF9BR+jKa8gp9JPaJ
Ng097QJonLD8NCQJVQ99UZIeScyP/a7YFU5998Zde0kOvLFrf5yACJ7qsezLMJc1
gfdzJP781ZOafZSIV0a5BAZpBSZEAjP2WWD9KmSRQTVJP9n9tfxmyXzZnoxh8G4r
lnWUy3chsBbnQp+rKQLMg/hOuBHU5c4zGHKh19SDznBEMKmC7ej7ymjvzKK2epfs
Y5BnTCDB+cGFJf+1qeusCrfDHKyPcaiV4Wm2lBztWi79OIqa1iAU2DQR6KxMhpUm
c/Z0bfCH5clPBPrS0vxG9vcVmCUIC4uNdB4ycqS2OUE8sSh8l89eWv/yxqiAZGRe
jl31RQ68kj08MA+4MgeknwCvFCv3zVZVJTp9zT/qc0s5u9gMHbCdG1M5UKN1VA36
fbJHtiaWKEtzLbTpd42dw3B2bV9MNRf5MB0/4Ikm7aSuhraziCF2J58+mNLdaBi/
zWekvnlIiS2pcNVahAws68YpYk8tFcfI7c4FdXQD4FdjDTiZMdPY+Brt4S1nALbg
z5DU77qDGCF26TILSzYYh3M3WI91tgMbFH/XV6TQgpXhgCeki+29M/nvQ2W9PIOE
InuRwfcgpnR5gZ9eA2gi5506OhVjklluPTmEaNgEYjPrzZ4DEPLd9zS8F0dRkNWk
6GyA0In3DeHWBm2zwaS1M7TU6tMcEVQJagOeOwfUXgYn5f9i19W/RVZr6TSg1jfr
BL5PLjn7ILvOO5GOCa3UHC9PyTaJl9yAzvo4+moWaR31o7ZiJ0H6aNhAx0AxVuUQ
+VA2Znz5Hez4nQtsBLMHS7pGTLS45/c3bJo3UrtsSX/fq8OoHlGayezRwkmw9yZd
CZGrSztXMoNfiCIn3EHdFSm5pHDAkpJ3rd/U3q2xrIQ7gzU2wq45Z1ylIgtnusLj
0/xRkMTACOaMELfTVibnTNG0ARXX7lbx5rw3siA4RqRCvfhaMJZ7LcT7Va/zatK2
WLQpGGus07Mk9GsMfek0wmrVncnCDGUYm5pNwER1NrZ10PK2WsFslCM7992mmIoO
vpwSLBihU8AIhQOYAHJ2hdAHTeSqvt6XPicYsCfJpxqi7/x+tlCvSNYyiHC8MEz4
VitYMpg/OP09XxgxldxA3bu7w4Zt2NemEKf6LpYmhtD+PJfXmwZy4q4TB3qmq/6N
qf3hPwIEUfiX9seVDphyaxfWaTS9mcKl1Temy1cUqQus/t7P57tk8ZKhz/t1Z1VV
n8GLKwUPazRTnDOubcvWulIfXetytYbwMNks/r+nzHoF0sFxpA5E5LZMW8/OpYM8
i3902cwchIFzm6hP4uYl3nLu8kvR9rJrklCJyhdwilcQszV0bSce/Biccp4CqJVI
RR24NCNAIwOGFhojJ9qoxJX1daNg3/raON1ArIGAMB1r/jBJjVJxjOPwC/dCXKdp
lrJ9GsTugCt5p62VvrsvEmJNDi/FQT7H7hoaDiq3z8Spw3DxEdjfLXL1SbBGLjsd
x23jSrLsDCs/wUmv7DMr+RqxpPuq7NtqTnmHsmWZIv1S3GYQ8nOLe+XEzlLyel/j
2QPdBzPOeiqXyjyFhBDkZlVfu2/5CfaGdtLeAWM4nA8wlzPZ2XTQyz+sArSi8xfG
L4Dhx/QXwlqKAsygfxL7jDW9qoShb5syoeLzwLimAA3m/h78yk10Bpey+8YwH33B
Dnutdvyx03Y0MqUJtUBCOvA2mqYdXG8Mh8vj+rjRC3AXUpm4OodQlt0PbqBNx2PH
x9Jo9JHFWaYv0u+HrHi3omIWLr1Mmox3bPksTWPFtGedXaI1vgeBlmCiJhh+UZQ5
Uw+jjFY95JuprNNzgGS1NZL10kICSJ20EzuzzPtOG+DH5D4ScMxJAzAAk/F9UixD
fVYKsWFhENSN/72uHlVL5fX3t/s7s11wxVhcsG/nMPdxMFLirXK6nXmoD69SekDt
7CGR7lumfb/YSQKtps8felLMYQl2rszzx14Tb7xKDIuLSyIEdvh95ak4AcjPSQq5
JJ+bJ3CQTjH+LDLlxQgPxI9lb6FECaof4gBSiB0Mv2HAqi7yhf1PxZjMS3MWMk2J
pxmBkSyups1AkSfBR3fjq7yBzZDeg13tbKxW5yWhCtVjBmOdJO6Ng0o1vERJLOQP
FiP9AiA7vgkKiS0h2u1sa9XIh09FLdr9e9cEljBK0mx8HZG4Wgpy+lByrm7tOpJB
Tv6xhkjsV77lnk5gf7dT7yjd8S59v+K0fc39x5IkmlWSBjrWbPbZmD/vYuOhrDlC
9OD3WFOA0mDNIjjq3YHs5sHRF3Vfp9sezjRiw1DTgTS2WzzAipYlutVLqTCqX0bm
b1Na4Zns/9ux14e/gahzBsildwcPFzCurwYeONptosk1Vjq3w0k44jcQXSgtUolQ
De9VniZ9RotTkHaJiLexSVTrxSjCBeu/zA3UOas/AYeTZAYEVni49REGMlpmTDdB
5z1mQGnXbhe4dg6PWnW/gESikR1N9oY5i9wxQCRubeHX08RzFeYf0zwzC5/V8e2S
OtDHb5iPFK+TAzA4S3oxiWOxO97N7XsIBhkYuQzA11AQ/AnEwNK0MhdkT1H3tfyT
hmwE07i9Ggd3bXSZ2WtyKKYLHYGcIdfjwxfl2xSjZllGlU4RVbTwCrz9XZXcLUp6
u3KAe2LTLYurFmVDOJXmv+/Zxer4VJyVOcv1DAIs6aiAcbeZKZFivGx4xFcG7NkI
4puLtRigfnqxs8Ry5YGYBha/Vl7+Nx/qL5OjeuIAJWQcT5Lu4OF5q0848Z9MFk5P
x26eaD1NeyMToN4BZCs4Ts6dSSyy89RzDarNd1gBw59VOt97p4bkv2VuHepf/tj5
9QAvPT3hopshtcPveVnEMxWgJdr+QHC5Zv116sD7pdy/5glZ+IxmStWj6scb4evS
gpG8Cvi4LfZp0IHR2fyxstzurPAXkXZrWKsFjFdNUl3OeBcAfs2LjbEbJxxwCqjl
+QKqyb06cfv5PgPiTWkxrurmD5YVKktjjHfkr50FE0UFCQ6RhMl1VSbjMBWxJoR3
fVa8CSWMAsJi65UsWq7K9v+ofRlF0dxWmXBv8TQ274PPREC/3iaSMTqNRGO6YpEG
TMidG/JpZ2i401tpeZnmNtW3ekzmiwBCGN1FhGuoCZ8AQTKuKqv30VD8NBvnkIYr
Knam3RuPrYZcSMUpfuT9WnyBxqwIIDSrUPFPeK+FvJuRYot8TFkOl0Vwfjs4Nfei
6kVqWCNRki3DPX2glxdCYQszbFWkyY0lLi7eZ7Q9d81nsJqIrgGs+LH2P/hhXU5z
AQz9yX88Y1a0wwB8wZlIRo2YqRD5fMOOANAVrcZzehnfahm9vGb4/aR9PenJk6em
YF9K0AD55jKwGIgEHq9QpkUOTQZ0KQ4TtEaP+VxgXEMcDN4Tv+8ViNhovJSUV0S8
mi/eDaGTU4MogQvWUKNN2a2ca/6Z6G4p2lHuvX+j+N3SeHxldUn4rZ168slqgzHo
HqDfubciF3iAqERZ07wI8q6fpvmGPrsifeF3AGlJHJAvt+RLVGMGnhxNQvNCGpT6
jQLgvvAOVT+XkPMuUBf7GkkenUPcoGhG3vvDikqhpql9Hpu7MCrWgfAWa7Tis2F6
yaDVmR0Iyo+wQPXkGOP8xR+zfuC6YkdiJfXrBCxp9VuZ/lxjCyseLh2dw9kH/XDv
zxY3AXe2WTTs7KsXeZDVwA5QeZ5KoBCk5sC1pW0uvThqotgumrEVUyzd4tgL9S5D
a1Cz5RH1vSWqJXbPVKNjstUIOYGIXT2alvqO2lGxdyrqzduxIB4ltJLWPgQDQxoL
sDbKeKrR+zKH4MofCt8GQntL0g00Y7akyGMcPpXVgwKhOvb5azWFA1/RKtGDdgWJ
MBWn+qEOXAL1nRyc/jeT4bmr3h4lTrT7dGN2D7lAGPcvb/MnTigL6FL6TjNZ/5ne
CZOGSyx6226ToS6noMnbZsYEo7jpXB9eL/tef4yq6nDkanAwj8cEZyS0GR6lxgwW
aGcw2AX1Jpdklx35ORVLlgABL4vM5i4lidIr8BcIQIlrCK5s22YH3i0TxLkm8Yxh
5/vspmb4Hx1N6D996BgGmTPtRe/+I+wpydhxXKgEwFAFfwjOEoG7uhlLrtwTPpLa
trCzon+lzv7uhh5xkpAZpz6Rf3eryr19NiaFA+GJWnkgdKWCm1GT2ZXePJw3J//M
XVyBDq2x4fOoCsIFtu0lwCcoKXm3XGVEXsYUHGWcpAX9kkF6szaQq0seB9PEVC/o
sGfG89oy2NsEV8AOJ/xJvV/3iSL978Nz0pMxxSRxXmfF3crfTJ4ZF1FLaGi3KvOa
/P2xljUyjnp5z2MdGcc8mwf3eZJJZbXk8951UjF7/66QuumRIgbg5e6ciF5wbsz4
i1Od4dpaYErALFzkA7j6615XLOG6dWQjqU/lBAmzaT0vyrI99BGw5xmQK9WxPDiV
7/4bqoGHFaH44VRsFpIQbawse4ObI/Q1ksDs6DgLyHdET2OUALwasVriMrwBQZtp
/YQMzYOAdHPURE9xNYED1hSU3f0THcdJaKpns9R1KaLntB2n2smjPl5glqYiZ38W
x2kIVr02WnlCkkWXeotue2XsmJfHYVugQfw/lgUolO4eD2PpzfubrKZyDEIR3BU0
Ls/9ddIAUnUfcr6DeLqRjEvyHHf84Z98eXc3e4nDbnzs234x8Vwk+thj4CNE2oGz
GpPsc4r8GMXLYOSwUQjI3IdYy4JL/bsxAnwoMOVttDpPqW1FptbVl4pUB72v7lqc
5gF4aVAoy3CKeBVNExFZ0h591C04mdghhM5rBqQQt6ZOgSdnTNgjkF81adGTWFn1
zIFma46aRiN+hMwpineBscO1WoJumj6Nqhigri+SwGIcYe65JzT0bL6ioyJwi+md
up0MOFBVZS/GdPpme4c7aIRk9fS2FORd/PBhKnK1e6se+eob9Um92vMzVUK3FE3V
N7o6Hk1QA1ST2ejyz9/4k18XRVU1oPbrcu4OqAOl1RW680kbjCL0yEdXbVfspK+C
vS+R+Vmtn0uIcZsxMrmhtzyJn+KQ2xYHr8eZ0/e05oL9BGgc+eZxtpUPkhflZIXh
uC/5H85CHCylmwmi+1NQeG2Cp90HxHtayA2cJuZF0oQjK9bO7Q1t4/gPGEDUk8fO
pXedjjst1Ew2eh6Pn9aIUQfi1SG7URhdIfgZXscotXqLVPQYA1QulBOwd+J2KQli
sN6nKe981TTFjmGTgSx57zZ27M0Ms2SDuv6y1JM/j44aiXMsc+bwtxFPrMjx61hS
Z72CUB5N9Iv2NgNseMnnWgc9JUfse8BGxgI2N2siDeYFtU/FWmHXJxhBcDHYs8qf
a11DfWGGaoMG/SQbELEBYRhDoeyNW9eTBgEH/+Cnk44jbe/oTyUFaMPoW36Eyq1d
m3N0lTi4ODRltycij22D9hSPydtC7L9omGTUim02zQgTCPKVvwMRroZtKBzy7TLq
dp4QHMBfGAZOLoPwwkEIBiUNbeUCo0dbUv6Y6M7p/3z3naiXJMedQ19V8mCneOGM
afHncV2ogy7euf9cAcAoxpZv8tf4X5WNTlM8CBGi7K77aUzBTy8hpUz+FdIaSTtB
4e6HLE9okF29gOXD1W/TuCExiltNR6YVUcs4byWj8UCm8GUe4w88IMkv7LSZf+um
PjUYmj5C0khkHKdR0rY2g2Hskyecuifrfyas8Iuu3uJ7fcTzsn5EZucqxKCWMTuc
aj0KC2JmW1cDOhQdG/g5Jm9HgoHwX8CoArBoUCGopvvGWV33t8QKxBsv/4p86z+j
T9+MbnVyNEjgCO2k6NaeRrV9ftnMZVzrEBJl/iqqWSneSnPYiyRdWyisosnuL+om
otlqWF8UqYVs1VKaGObvf96LqsQengK+3rzUYPFqqx3alPdwcYhz+4yY6/6JbaVy
UIM78yj0dRz1VDYckbr7QpWM+1u5F9T4ZBYJlL6uJuqDKwKWpe9Uda7DPzTb5SlM
3vzQr4udhB/FwXwvO1lbyJWeGZwsodq5en/GhOtPbeajYXCucHABYxTOuV0pYBh2
PK2nVDxAquissyyB2khY7NXR/L8oipm6DSFZuEBFGbNt/0JvPebZnfgofonSi5iO
3iH22KFGOvrb6YLPzx6tJ84Q+0W9oxHyAEnvu40AU/0KMf127MYmONWCXuhGr+Ec
WP54D++ov/uHYefbbBrw7m4EZ6lqEXruyt+TmCFGVZRnBYm+AKs191kmT2Y9UDdx
KiIQ4Rx6CkSOnlJKYIufQnvZVC7KCK2SvLFH3OcZO4A9BqBqXfi9fdoH1ubSG2hv
OTIZQfv+bbr5fFSYup80dS0I0alKK+5Ft1weNf7zsClFDHnPj4rc+ylA/8AkBnQC
CTWTzxo7e5IpLY5vGyeir7Rk/jVpzM0vww1aGawd5Q115VMDHBETBay3owJw4tlO
vQy2diM8VpMDwWLSJyGIvd/Fe/5YGNn4Oej8HeUi9d1S7epfAhJYrOSZ521NGY7N
mr7EPfbsvGrbuDUF6PHxSirjYAvBu6JECG6MfUhHOH2wxw3WnD1Vzv0SV8I8458k
E0yHVDYa/JQpKVZp166KaSqnauv76uE9m1slEWcmEpFSMlh3fpLxf0G3GmEyRHau
eyW0SfYh5n7a1oaW8qVuJ8rcJIrciC/SETGY7R3GuWNFEg/wPopzYdcAfrr4RNSH
4xzbyWwHw4GItVPgEUyTMwef5gWADrwEWc4G8hP5ZmhFDVTHJXQvHivyJ02mVnJO
pUvFsu3g0b/Gtdms+HDtKpl+uNlgvsHqN3w4RciuDHfrmzUgihaPOYDvgb7mtxBD
qzHLo5lv0jNZWk6J8+FXdjQzoPMBmpo1gPm9HGsYGQf03LAXVYoobhorDDzRIOlc
rEIvaVczegGY25OHG8celdJmLqhrjX7xOLFzHumGK6uPAlzSpslKsrbDAPB6BH1e
S6WHemdIzcw0xRXaOg3jcnVDMJM6Kv2pibvoX1gabXPA87x1mo3YaLZQGyEdHSJ9
e0sAh2yFmJO/WzXKRR+TJRQtbhtIpI1StdOKzCqAbMRSXzF8YrYB2TjwrNRi5aZD
qPRxgDkUKEmXURME4NhOMMIQNqcUDpjE8fmjC4TP19uV4NqW4vhFgACsEMYqm2sS
qRbKF6ub3SGAfhUTiS9XNdIFBhWRevrCwrzMGwurXKQB4PU0jOhaHpz3+hy8ekOv
t8A/vTERzxTtBNwBMSCYTphgPZw34EH6xP4TPpgxvebsv1u4ewyO/IT6JgTeHrrM
RajBUA9gbxmJtyEKqu297H2g1bqAzFIo1+EJ/E4U1dDL2HGxOhM22ltYo4sw1Yuq
cRoPrXjcs8jAQrUYFtXSiIZGbIXN0jHNcVa9LCt3Iq+sra3L3SjkfiC2qG0fEKtf
LTw/kKwR+3LzttdyOOYTtyFqlESP+L2LnjJEhxIARYN1YWiRzvLN79C3pukeVb3T
x3LaDZke8vjzSUTzVZtZ4/APJJHDemo+vzy3J+dXwMyOUad+yqdjZRu8nJB2rUq2
bcZqFQDxEAUcqtL4x4gdp9QA1Hn1dsAlNPtwzR3Vf38B7xFHOoSbR1WFQnlKWN4Q
iAFin1b2EYgHxh5Ok/qDjeIasDYUqA1OVw/IqnmbOLJ7657JXUeGNqTI0ZZNLlDx
KKaOq6MPYSqXn6BZAdQCJWtOf01d4hE68QZZ3tA7+4oBvr0mFDDQhjsbcZOWnCMp
22k+jV2iYTxC8aWNvbj9nXATTqMXuj1ISYsxbD8XbYmkkbA0ff1kz+dI/WsmZGWe
7ra5x+LIJ4CMkxlCtLZbDrhVG9YYwqK2dcrlB5nC9nDc3JU548boNOC0zZ+/lAQ9
Qq4ioSoba88rHtlpsosGf3b1DoLnQATErVDddXhwwMOLtOJHLcTiKb7Mol+8l2eV
Wnj/h0I+V4qpnSSVL9oReXhFxgYiBAqFtQ69GTCnyuezBiEw4c4MAq8U+arrUWw/
2758+kRAOcr9aSh4vdD3Qg2/AO0gZKc6P/l2NIt4SFFi3xw2aKmf/iIO4H7bc+C6
TsSMOPccpaTb75VF9YxsQqhQ6AW+cJtupJHzbh97my/YnoxflqHwIgCYLHJOYe6U
JYrN4hgpEReIst/KNUQr+z4ZoJYOhiDwz/HHBpCtFt7A2o3bwswMA/xIOIlEvGoE
q3uC4kBB3wzAdINCKBnNPg==
`pragma protect end_protected
