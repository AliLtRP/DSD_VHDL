// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:11 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
THD/3ivFIGEENNuwt45bSB04k/3blBcJ9MMa+E3mebeFBcPzMbsdWSi3a12lCtIW
LpXwSio7PZ3Ci1w6F1VMEdIek8EbkLsgf9y4uAeFurW1bWGPWT/J08x8/eCl9JPL
UiAf25m/YgMrTObaWfgx0YPkGFMwzWhwje+6AjMrBsQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31136)
fWjSZ8r1eJ6RyVD7TGPUsgdSL7zlil1FY3vLeHvQlGdIHC5OK5nRBplhplekrA5F
+T1emmNLAtMxC/qTB2yp0VGddQTiOUyb5wPjiEz/5QW4/uoRrJnvcK7iAIvBntZZ
TybDVOFo3FD29Vi365ktS9DgG7HkBcOHj/Xd/KUf4w0Rbqx/sWx5pNRGaUsc///i
jo/NoCHIYmMEhIX/unKjajxmO6FCIjylWO+TysXcZckA9xR2X6bYI+JDaKy1WNsB
JoyAsan9rbwDrz5IBwGVbn2bFjbxPSxG2vtBnCbhnhwosjuplzXmz3U0hZovW6Vd
PLSKXLRYB9gf87l+FLsG8JjarAB8yysIfxwDiupMx67Me4NMjDIXFbGPBQ+N35Hn
vq/tR6g2L7psWAuR5ZWn8GMjB7rJuEKAei3vYuY+ni7kYoXIFw6NM3fG7pgOF6CH
8sQ9mA+QXj+gvwWshUUOD8Tt50u1hmigKE1J2x6iVZqZmoiEjvchaEHs4IDJ1IFt
ybwP9xuqzvhW9aZR79wg8oZO3AtcdJoTO5+RNTjaWAFjKioM3HMwszIFmA+EXu7g
ntQCcxjE5wfPiui6b8YNoK1afieQOJE1ylstrKGRMDmb7R2UbOh80CsGr3qDg0RW
biS0H3rLExGVcwkeojUIquBfMONhs7kAMBgWU9KZwHHQuKY6hcWvmMRnN1ywHs9T
Zee7V/4DDtk08osFB+2WPBeKiKZhsO5uXPuSY+7HJmU+IDrnR8qb4lm5nO4KSqbO
sol5Bttl3URJ/GZC3cXkTT1p1zWD2mmbeK1y57VzgO8f3Ci2qQo2HC+JPPuxXXrX
2Y+z5heUxHWJyyRoWg4KEFvsASS/FMC4HSuuycgpphbncBmdIlZ6myCtqr4Z1D2i
2ef7vmaANFrey3XPdLC0nOcZyTIr6Rj5ZiA/tpWxw8DltbHNLtLleBDXAvqP57pm
Psg8U7APvQiT2qWwoSuWye3e0CgUeosdfCxZbfOiunBKf70IfTxF7bGsbKP/KWTF
/R3ihRn3KwAOLPvFeIlQN2Ugu5DLLgwooRnUVHzt4ZR1Kcpj4V1x6Y9K+fm7vtwP
vYaUxki9TudiuBicQRiDnC/mG34RMz52NmyK2zsTFIXbqlQlHtZc0tpgKxQwjLva
OO4dyPCD0fXDRLWy6lTkwz0VST6J4CGPrXyZSrIuuy9xTc659jzuz4uV7lVLeHeX
Wimm6T5qz8YLPvDQkNbm0+7VEW0y8UiKpXrD2pt9lY+2RDXTJETK/gyjXfIHq3x0
cCAKXCWfC95X18/cI2ZxABJktIlk/YdH37JECB2BfgUkD0UkWY6vZXVFs2HtOyjz
MgKVqUc0gOiBkFWdq9NgKVSrVSIuTD+tH2rer0ImHodvzkUB/MOZXQROElre8afB
9QUDnbGbOP15ilZkElOSFoaGkMGU2YSXp+AKy1z68CZLoubPez1DshXsDLximOXQ
dGAuNG36LCwZptpfYW8wqoji6gDMwu56ndV3zJD79caQlsg5zXK46XmY2Ph1TMb5
aXPwBhX1p5reYk2dxOXllIkoU6sR86n1Z3sZj5oSZh9DNUhnYoTFK61DVQ8aJm0z
c7YwfDV3CdrK6ZQuzHx4q8na0sXTdRYn8+mZG2FbRbNAaxf5nKNGAOT23esXHLBv
XPh2g545IZIERXkfR+ifwUJneoDyL5QN9cApXjL28RkVIKUpXSrpWsJbYLCBQ7aZ
n3v1R8jnqTjRBwrVJPtuojMt3HicxRQNRRI/uVgAAPZBh3y4lAYooAYL8FuhnAk1
8sOMJRffxs4e3xycvEFA4jIa/F34nduq2lQesUEj2NSKF6iC4fuEqHrZ+llBQqgQ
YIASC0FOgf1Fz1SEzSCdYVXf+Xk2/UMymUMZgdMeoaw5PA5xtIB4EvQE97VJ2Qcj
hg7BtiXqkLh1AQtKgyYLlOzz+la8E7WRtYy+td/HH40l2fvChpp25hZuKeYcdu94
6tCSrapsG2P8vF2W4mW8PJGqqg1rQy4wCX4X8xMFjWeGBOPYGhZPg8rk/1QWnZ4K
mzBvYiIy1tyBOoJrvniVaxaXYs/18v5K39ydZYbimjY54KYUXrlBhq3++4JFheXE
tkyVMG77X83HF7rKJ9FRr0ed2YbKJvGLUSAjOftKi04Cub9ESpf7QdWjPvtKkTfN
a4idLJ93hOnLa/Ve1l0jUqA3Z8JSpi7KfmU6IUwiq/fwarWPjlC3Pyf4UE5ebbeX
0Hpkt+nD+RMP/pEdN6Ny3BOQ0kiJ0J6ONiXwwn2/k+I7mYtZgRT3mH+09FsUZHbG
cii7BdErqpHAFbuJoo3qXDwQGcXyHoKQHTcMiXFTslI5n0DniL5nkqtCK5wmHPv1
kb6W6mZx2irdZ/sd59A9B5SHYe3PrNCEhgUQ7VUicWrdhcEN7+9YWJsQAHH7C3YI
6Km1fQ3yP8YIMI+PlGPx4a7NyobHlQUy4ScQBmcw0HStSG4y3uY4wxNGoz0oQjnJ
zqJZ9XZRdR0bLioc0k+urMAAkMM42W4OqSjz+O2F7gZIy/uGCMIvackR5sczvfMs
pMfQViY+FZMdXRIdTMtCKKDAh2JM9+usW4AaoksnJc007fw3d8I22pa6ZmQkuOll
2mPEiFSkDNL6BnotjsdD9vXo77aqvWcJnI8Y42OR3bqtGSRl0umFXitIRGrXRFAR
9dJbCMfJsTS9yqozSTDHJ6/OmazqmJ/RVQmfSv2YgYA5Zh8aJje6f5FjRUFtcyvw
Pe7/qtdghLy5zBYVjnlTZWKlVRRTxpVL97oMKtsrxTUOyE6qHgTAoH8PHNRne2iK
WNPmOvXNq57ldzucYyRjOAFOyOqEilhoP2Cby10VVOY/LcZId+9R5oPOOnmhEgf2
wKKFmTSfy3DPtApf5HD96iUEQjQW/I1GC0eFwNsE2hb9e95W8pNqoakftEqsvQWc
OfY5m7t9wuVEzOYMosttdijf14D7G2Yw4cWacDXoWIdFDWJ7H6SDGPPE5+SDj0Li
lcKjXXbK6UG+vR2jPskpIvFd57aU1IahOg2Z3UfvYuQosaNwoU3d8EM+2rchQBXR
QgQsjxU7ThwDXkgdNwimFDVn7pZps0z4+AcAFkgNKv7HXsdKmE5nK9xIHoyzC59n
uROWOjktKC1H65oXe0V3gO3ZrXkJnRixVZHXm2V+NQB7og0Dy1LFbaQ92Q4emUQ7
LHsJfj+MI14n37YysnsgqJyRmIDBKWGuAUxNailz1xDrw1Q6rvO5IUVD8/y1gGrj
9nPDrj9720OThCkt+dm+oDc5+umE1Au4NiAMEhwdgLiqEvX/1RWZI0E9qAKKncFL
Etp8uwJbM+cR+qBQFRyBRfNsqK+z7XDM4Cyk5vEx5VfQu8hPRbigLxou5m4h2lK4
uH4QUnLRV8mjUPyN4JgX3pYof8lHf7w+ONy5KkU+o4jioRioxsB49QoNGDEQ5Nxs
OXiSptpZQA3mH70OOEU+HfNo05hNq+s15EE1ZHe5Ichiu4PuqBdIA3F6DPKkJjMh
e7zaNvRUjgFkLi0uXkqBm+NfOeq27mEKvnU4tFk7bK4EYEDOgEMHRrpChIdrc0cx
fo7vZrLCelpomn550Rnbxy++eGhxsEmC1PCXyJUmcJdDg2hK6wIXrLAQ0JhzWZcp
yNhMbs1/isg//M4WPHSE1BbHs/jkPMh531P4PP6qHGMV+WReFhFUgg5vQdqBJpxq
UAPlOR+Q47oXatp+XEn5wc4Vhsvdv9pTa81104JCGsCQM+3C+fBAZLyVhJtsOX16
Z5H3KaVbLOBxx6fW0J693hoewdNH4MFgPzd8PfvyeMPEzqzyjSYz0KUXUuZ6XKH2
wVpIqDmZ5n/z27JioIjn9bK2fJgcIfnSc+nRh7ZCCgJsPK1Xx8wtZkMZ9gjjgGG7
ZYVacaIMXol5XaukuJ7smjPzLDFbgzMjYgc0XgbgTiTzqTOdzYiEc08giEIyjSla
CCbAY458bAZSG5rr4U5PaPz2IBiA7fYaNWNpnK8Kc6uv+kxnGtdcPKp46dYcliLk
B2Mqzb8++HmcovAuP59L5Y//SczshbRmL8WIzB1SNl54EaM/GRvYqqu/LCLaLw6U
D+k8FVp9JuDS9YNM1TTjG2YwljIKcYBG+lgJn8xaAsPmDcjyZen4lkmVocB8axVs
JvMydCGHY2+RbtlNAB/uytuXq2qKVobgqjke+0sQmUwOpVULUK+QGY4nYBpN/jAo
CGB4eT/PoZgkfpoYRjAlpUUmwD/0OoxSmntyPuplOz/VHurJfvTasSbIp1V3jpQ5
hAWTLPt+ZkPGbwIvgIfm9TXG9DdRRlHXN6qISZuBQeytNnWaye1kwqc07VJUqmRQ
ofzKOE+mUPIvAETt8dAvEkvlPnCLaY0Q4RWKZhhP+Oaif4RLHZCi2NdwHC/8R/YH
yR/YPuYMqIn/frHn06Kl8xegLwRQgb11uoJlsQCtxWk8b5lCu4+OfOBDeNKI7HdM
zu0/kMVwRL2lJRqKL7za/FjHHeR+ChlcdZoHoN3uDSL+eU7wWqTE/ARJ1YlPlO3a
TPN+Rcyn+f8YGUwRL8g8S2YgZ6CiUpr4MhR5i0CtB0RX8rvL+5xIo3HhHFkjpg/i
EMa0fRZy0+i8AXEXCLTDw/i38gvCvL/pZ6igb8bcbUBr0mzdVXmwLRkSt1K08+kp
fhjExa/CNTGgHrXeNkb/oQaSfWU/cCQMtWB/j2VVC06Ojk8ckJGpDBPFyDue4VFa
4sg7vmW1l+rHGb+0qffDuElcPK28U9+9v0HgbPf+Jry8wAnpvffu9NSg7Zer10Ba
qAq5RVNw46hgVH2EqSwVl4UJmnIWG533VUdHvygNr/xfYrYHClgDwq3TjFDI7oBb
ZcpLSWQih7yxcRU+MTZ9WRutbHcUf4BVND9uucouHn/dsz1x5dfZvVdE7a7Mw0QC
pLs5a+a0RjJa7qe5FTJq03fmAQ5Yv3Xu9+XPP50LXqiENHxCaCTUiPJ7nbbXj+Pw
9PRHqZJHq2TFzGq7W4hEFPNjTkcCImXXBgie2eSgFXD+WLyjXQpS0lxkvQv8sb1K
mXHJ7rchkVrvn+niQsdfNfX51gjHRrFZQlJsXyuyHmEtDyFILF4ol1cyp71vG9KH
5rAPcr6nETJllXgrFhi3NoUOnVXQDjScXgWRXx5AeVwTJ2yS4c7//aODxKwQmtUP
nWYFT7QlSfBvaDu6tQ/r09B/V5KUXlmXW9IT2K66XGtwx5hlEyFJvreasHFgOFby
OCYuln/uEUKcHX2Pb0K+HudCnuBQjVBt9/J6qLCVcnNCoBCB5IBgnJ+6Ep3oSLJK
WW5OAFAi3w6+HjD2ctPa+dxBqu/EVgyLdcQvYu6Gtv4c8qjwUELX9uCul8ihbkzd
8XEYz0Nm1tIEjuhC9kXZ86d434ckVGb3yfWH4ghJ+Texf+YaB6C2eF4SEx/xIviF
I1KAm2/pRwnja96YdAFAQIGxekrMNCjcgDQWbhzI/8xXcDRGr0yqNWreb57g0dpZ
uNe0E2GddyJIQSAOnvqixkI0arIUGMcB0T+yBv4wsn/NjMAL5QZgdU80Mz/l6o0t
lam68iG792/teGFlXeKfs1bCZbTLcNbhwHIcBtN9CB3hjfxnK4cxxpo3WovZwTRG
g8uO1wD+l4gYtmU1dm21/lTw9qF/ijw97VEO0nnAE47dvHQdQI9AKp1/c0qB/BPc
y29j+DOKuI7c4ZGH6pY0hrAqQcA/V97yepbDmnl9msQ8PERJrlrEBeqXjYF5oAtJ
dp17Eh28e9AxH9IUvSsnSLH7kOt3D0Xz99oLscu1+28bHcWVW28fho+v1lfNnpsv
8QhVTKCwZHg3yFKNs2ENUa9YyM/rzDsNa+JLdRZmDSLFqKJhA0kIvMbwaddI0prj
mNfe/xgH9kP9cph4NaokE1vde9C9tpCBymu0nNolYS1AXaZfvRe4tPgS7/yr6CkK
rYyXfHGXGKDq4aaaiKoAbrYA92qG0Pw1t9z2Clr/4fHST0rWEJOxGrNtK/R2CX1N
kavuUpYUafWun7kWYvql8jDaLxsdDk8TocV1t8jcTojBqvEf2Tpm03XkautE4UtO
07dySo2xBejD9TJiOw887zZJ2jcU83tW4gNHX3MPoUfocv5wIrXectQ+51OFC61T
diWvGa8UPtAin+eSYcxdRYAsh4ivEtdUNqXKW3mjorYG19g1kVKU1538gyp7Cmyj
g6CFGRFjX9j/CQjzfsc7ixcf24SEGL8orvh3ViuOj18IzvLhNoBypfO+9XVjacfn
Q7OYTEyC6KX6cFeMSbc8JspcAiLFvuDu1zTpnXWK1RA5rI545/7T+kdJ4No6+BjJ
sFTJoXPgFc/9pb/AeCa+naQ5xJhFSvIQr6S/UP4hk6bIo9MPexUD81Xss6gpdAnS
Bvs4bLHtAetORJiPXWeASKyZlfmRvs+h2rKnIJIv6AU6dAjST3vV72teVUeacBIv
M8hLB21Twd9H7cBbFP+g7IIFZwurv3iO7VPFirXS9JiWnMC4+NWrqAZm1s2uWlku
bDw5OIEU6QstNO4jMK6/L4Q+3Mdwer9CNaiqaOtytZqZS7ocI7HQ+xeSOStfcjX0
nAj0z9R5GVQpptetlDEa6/T6kvXhFC0yzTbOFfveqvnGvY/fA6eiI/64DXDAwTtN
2DIH5olEKDcRpmhC+IuCaFUuGHDQx6ZFJse3fUIRdsPDJ6ShDmUaR4TUKvtDEDxR
AZRt9wL8VCVjzT9bLOxXJbDpKIL2xP77UnxENXERK+pPWx69SNB2agcENkATelGx
Px6mVMiqdXyjTt+masmGiqiIZ/fWR1QzIC+yJbHHh+5I92NZwXmsAIWNoDK+H+nu
qsEBZg2meNvAKYQ4G4dSyH0x/ZnvrnxZ7+jXO6knst7f0wJLtaPorUmQDCsIgJlo
Lmp32J2Q2uLn/DChorLNXkrSmUgRY3H37CIZ87XFLpUggSeWbHtZ50MDzlbQ2ix6
v8YxJeHUpCWWTGIwnTzg+Fw0bOTT0uYZFsDhoqTcvgso0sPMsXGbAsn8sGFgfnLP
oS2T7n36ZyVkc+glaLOUVxC4n62Hy4iZ++m3K0BlTTTLB7Nt0lRxq6s4lkfTNe5q
GGWv3fQnWFZR3SnchSGAPz+R7zUpEzak2fqmnDPqZK4kHkiLNq2NWZhngrsSsVyI
wTSUwXYh7eQdLgSX3DfucIuFZRo0ByugwajTpD4svDfUtOgLn8ZvLC7ENgfIYUmW
QxlHvrDXPYpC+fyf4hCavF6cp5Xfe7r7TIiWGngXvst/X21qrAPUYDGcA1ZW+n8M
o4nrs26zOiL5+5u/qlHnN2zyjW8vH/dGttTxtANhCjtNV0ei9Xvltx09rUK3RBEC
K7h5Mkan89LWyNDcs5iJbvSfPxciQprg5gLhZ2zZjDfuXD4d/jJbxdpiatY2X0I0
51bGMXKpJsd6cTjdCR5GKq49q1nCe1ZPGnlY9AAlpYYh7X8O13eAc08DBpIqv0X3
scvtM/G3LsPZ/cHquoM1l4SFLRfRra0zbKJ7E2KociwMdhStXe//sqZQ/yY3xbhX
uGVxOTnd7K0u1gi/KuSisfxvFqFfOXSiPilzWfenwCOQ2mgP5CZQ2dVHe/UoFELA
xFehqd9wwiD/k/HqPyrrlyS8nZtqhsIsgDIi8m7kptNqzFOPFiYzZjnM4WILejK8
EC+YKsK1YObiIXar9tl0HJ4WQCI7ZoQIux0uVQj/UGx7pimkvPs3oUkmRf0hLXGt
vUhrezRKIeLZbZh/DT4uTFuvPNlPF/W6//zdq3T2mSjamzyb/e1SeEZGuivU+eg6
usIn5zj8AmA+qclfnSyNU0yw+5b6TyC/nUsE1UXxxS1SxUKyDnOBQjz6s6MMYJDy
LxLNTt6fxH2syoZX/fDwdIKkoPFwkqtLqTwO60ve66dyn7YLiFkxmCPrQCwGAwVK
kmPPQatv8L/GM5Qke2TdL3iihC6wePGfK6EwGezimevO4kymFM6slKFR1pta5Kj8
ZNYRr0/+GmIFacmQL8nvqz/u5eEEeiFX4oxU+BMSoG58HOWQqUxom8KIvxMw4wfk
gIjdNdG8p+pX9/DqJn8ciMSJybPsIkG3A8D56llJ85bin22NSxYqKbXIgNUphaX/
6jG65Twm0IW+ZQNDvynHU2B55+uS62pTKbvadKxgKmN1T0A11rl1yWznS8oge+LJ
kG/i1VoN1XP7LgAqeJLCKMu7NcVdeuv2Kufc/0UPTbhW7k9iPZR/3rB78lM2MDfr
wdpOMzSZ7iT1ACSLFk4dOmCibk+Q6P+YHDiSHQREdzx+FxBtoOYBfvh8KjII02yy
4rdpyf+th89exK/pGFLGP0AgAWq3HPoJpq14CzmOD6vqTRr6ZG0GzbshjVsL2ivO
EBnS5iwuJWpjjtqDUrUzAVoMESaEw/zbrsjBg5WWVKhSE1sfMLeCj0MDEmW1A43w
FTD699CnhFLMGXh0UieemH1Yjbbp83qkJMVPF+NVSlkxzYQMjExgWOarKmO0AVcs
LEVEj69msTjdS7gSfxCYsuylyblNhLe9hQ1P/hGUi7ig4p0k9kjESTE/1syM1Sa0
QskPi5/bhvVADyfFv5vAmP5/x5OnNWl2S6+9oCeH6wQaNDc7IMzxz88glW8CB9ZJ
iG91J7V9RgOawZqEcSF90sK/SR0Jsq35lmTyasWLG0qb7ysYpIkfV9INueXW+LgE
pAfkGV5uqVE/A++0PhcNmxdpZlwkG/fRY94mVDmDpwM6QgeDVlnqA0d0ZDoa1CzM
yjWiWT8NPvyHNdHywVpf8JkhH9DKs/iAzi1YX3MBL1dvpc+cKegX+M4RUZdoZImq
uBtduABKHqyH7UO6hUPQGQugcjWB+w8gE81M/1tRbCCOlMPVlwP8ZRM4r5x3FPuA
08jmaFKKjKBViucYHfSHGyvqT6GZCl0JyZxw6oBWwS6IxdNCTr+ExYWK6Mp+aieA
pLZUW49lptuD+vQRCoN5Iwv5/R1Eq4oVyd71fKR/TiII29rhLdyWhUpAZoHlTUpj
RDdiVVF0g8DSzSZfg/gFuiXOImN7ah1mxv27Lht4MopafHCW7WkzmS9aRCcJaHQI
gObUq3otYU2z+BB99JIYMcvAqD0g787n8fM44FQrr2XhRXg6O70hSp6DvTPUbcaP
GOanm9qilhhq0Q2qiDLGx0GdR4f1ZRd5gvZG7V3qPyzPJdvuko8dlTMjEHed2DZ3
6OXOoFNyKRDn87S84259uofQcEB3vnsd7kYTFCeGwCTFC70oXz0vAlaIakVX7vTY
IeZfeN0oolxAg92ZUNG6l737x7XQh1gk+ZsET3HSfxaTI6W6Gcs3d+1aW4pc75ig
68VaD+/jZG0/0xOyFUC6Genw3ie3yk/7CARd2G0g9pK3y3PGg95nj4nSE8Gritbt
Y5wEKwudh89gnMzkIvgppCRffeRLo8iuWRIFfghy3HTByF9c7vf8Y8RQmtH1zKAD
S7B94ITg7+sbJS6Vq+FfllhvQhYDr03FKXDGyFMB4IRGUgOI0T8qG7vUlwwT5xcg
1DqtfnRvMuy8L/W4RoOA5fqaycF4+tBlJn7/5hPhWQHGjvaVEr+zHswGbJ9ozIKp
1zCQVwHiXwVe7jdMCm+mD0PRQ540e8Ms87v0r4jDklp/Qow9pvY/LBvDS86m0pg6
OTdAFXorVFURao3hM1UZuNe42Lj5W90RAHrb5JmYIpPxwlXmpxXmke4C9it0rFAe
c9GrkaTIZD4XUac+weCLUvQBNRNDK5+A1KC5eMTDdZl9ttM4VhIbKEE89XINHWYu
HMz0gWLoL6u8yfLAp9S20ab1djFeoHGuOJjOJIJJa2Cap0gCQQakJXvdfdJ2GjmJ
mcNTshib+kvqvDz7ncQB1ClO2/DohdZuC/84btKqAeyjHtputvI/LxlLIKv2sAfv
FcaOK3eTMD/rPEzP0svPsBSMt7eliK37OfFcpP92nVPZTmomkmuOicxuZl9OxBrT
xIuisD4ppxG+EL0FTpQMkUvnpfPyPZGCM1tcw2vxJBnIBXgV5aJlhVz0K/G0OsiJ
Fl6/0XykDppkoqL6x57XB64UJlJVs62ykR3tEFd8HXE8ZiwXvariFH6cNa7rG4r6
Qr3TS4Xf0GIYoskEJvX0R2UzzQHu1Ou8xNXTRbxY9fOx/9KXwGzF9c3urdLRh0do
05JZh5TUbVtOADc57yG3IiZBHzvApv3mAaumVHyrZd+3DFxsahS7pCn6lsvI75Pc
wN2UArDIpL4UDUUtisj7T5dUujMk2TD9FErYArttkExikQq5ALof18NgB49iAJZG
9U3yJgsNRYFRBRLQbMCtqycVQ9bV7Tgigl2zDQHQF4R3Bo2gb/4yo5h2MkS3vXHj
p720+vC5T66/YJnrJdUmMwJ/+S2+fRPVWji4Mft8bZ/kWFG3p8yh4MTyA/zKJ6zs
Fyc1m/Li6DxooGOC4XKF8ZnpZ5yie9y4grNxhJOxH6T543r2CA81QAsioIss310F
T0H1P70rAJ7saT36NMJSKEN4aVaQZL9kCKz4jpZIXWDAcplmWq2CQkUP8BMS0TGQ
odxIPbceKQsul4H2FisRHSq5LKUs/DkN50tyAe6yFkmKSfHDnqlkInKX5R/OCbOl
5G64aia0Z5cDYRqpsGEop6ksK2G71OD1JfgBrAPVEmRUk+ij5OUfe6XYGMuW386J
OAdaZYvTzU8DSSKJ1MbYOobCrqFtAUHnVNyaw0eRklrUl679zjm4atMdq7uK4din
ksZ/gRLxMueacInuqw0es4xEOaAHD4NCjytOgwhTEMaJSLMsXxYfXfDzgbf2Zhjh
diO6x5vR2DIXmiRhzYCGMTW/ygBMxaeen0pIg08bLSMligOsV7LgdTwm8QBSdqbH
9Ffk0yU1Jd2rqakbBNbFYT/phKXEoPmzC5Z4+oEt9gyPe5AuEtsOBxRIp9bT5apJ
Prq9rKIl1RQv/DHPP4nssOAh2obg3UvRFOVLgfKBfI3pyuituLER1w76m+se/UW6
A+JXDgJkJAXkKVDvthVFDvUqMLXdq3IvDhlkMw7HLw6ibQgsVRl10s3Ib0//+aQs
b4FFJ9ipIk674Ltk1fLZ1wPZc3m/jlesUkrHQ/85DIQAUxKqOFT7uuJMeeXzM92e
pft9LNZnzoal11PzsVsO4Z2uDcV5BM3loEpoEOI1PJeyqhw+nSY+BHExMAip5rj6
74mEiUhO0JJdh1o2NTFeI02JUNG3VqGVc5oYXp2SAH2MaDLV9Wh4HFFai9X99bMa
Lu0303TzZHhDSe0AsRyLefWgq5v23V9BAhtDAAyI9eHSvMuV75LR5RclGngD5rtr
86o8lrIp7ZV0sncSg/zuA68dUeiTqD7WK4U7O+T2gxV/Dy+HQNcb8M6cUxMMq6jN
rvz+HDN3y0L6kRuHzzQXQv1er8UttQLhfwFMv0RU3NA55TUdPTp8dAybir8Sclu7
mWBNWxl1XZnzBzhQQxBuVJaG8pkbR3EDTvlxum9lwSKb79Zi0zHFzkNqCrhc0DoP
J8x8FlIzkM4KaGWH9bhYP//Dtt0XkOW8wDBltPj6mpaQ/CVLKd11gad0GxMmB8lw
trdxlq3hxaOBR/+OKN+qsH8YrGCIDvYhmgP0PjF6Q9yuQWFmRwc8t5yWliWJy6D4
OVKfRrg408qnXo7xvMkUe9ZQzMp7LZ50iKvpbLd/V7YzaU2bX9sfTBzK/NWaQpZD
/lF1R+9pskOeNUIQGrHPTtXqp5OPeh8zZ84SabpZUUPA7Uucm1EddA0qfHdzB5wG
m4DNYCH+/RnCKTvi18HZEHoCYo6zXtz5uJ8MVaDVUoqlRTGDZuYduhmg0Nt76PX7
6B3otnE8KIp86rVFfm2v1ChymM9N53BWwKnaAufuI+ZetgNFNm7GFAEnGgyUkyx0
3qwoQx8b6rgUJaNnmNjqS3SI/jZ4zGIwlfkYo7iRgsACIpQ7x9H0yK5YAq93Gp1V
xIUOK1Sts442GiQdp2m9dJTpreX0Eqn7YtnwROXrp5qon6LaxNeB2c1hlX6bDD4u
JWdcv+LGZxecFAjnJNW57nU3fIcsc6+Re6S2K16RU1uUtvNs77sg2XCXS0qgbuQj
WbWtMQ7C80Ntn9drU1g4+X2o2g8PZUl0CkMIcO9BSiteDx8WQ7iSnxpibrarHzyu
bh2ksR2uYvkhKx6W37/fkSzIp7gstJWs9Fpor2VxxRIMo5lPGtkOFsocZEb6AguX
Mdv5Cn6duPLFTPqwNRbl+v44QsodddyfZ6HcDLnhOoMp1/+4BbJEcQemQSMQDzB4
0ANdUNO3rhXUnMUjSLYrbJaPmg4s3mnVCSsRH20s5nSyfn5PstRKAhwsjEWtpdH2
T4MYbzmWlQaOV3BRu/Eup4qzdYW3strVGFHp6o4KNQGKT/tydgxtV1ohLFeoy5ve
ghDyfBpuBpZYgJZvRic9nDlMm0Dfp2a1TgM4zVJul4MVtsglNjXY4ZmqVA2S7w6Y
rvy0CMJDnTkC18sGpPD1/FNSB18byz9Jx+wV4c9S5WfMHb3PXaV+GSL3mHdJxj+W
iAj5wrbqlWGKKykqyb0PlfWoPGAglWEAKp1k8UkBEEPer9kPHpcsRs0SnIAgnmsS
QNpsfypvVFt6S/KWNPbyhVaDKki9qvWiJee2Oo3p2FIWrq1dfeieNSxv9UgPIvM4
OgqslXbwXp6N6dCBcn9FJ+zaegqJE7/BI1DI4DLWPmQ6+yBpuE3KDCu0jvZVyF+5
3eYhvdD1qgSAa2gN+uChxD9tpmWZn4dm0DPIrUOwnB0d2QdvjjQlV6KIF3FBDjRO
4ye3k4VK2UCLqeKu3LA+TeyVzr0Ez3ySK3hEkcVPVLQ0oN4HF5tLdp5lJMhD089I
ObexSppWnlaqO7DDRiemzVfBAPou/24EIFk4JhsdTdIGR0m1/xpl+yizqjpJHOHj
tcT72VshksE7ICv0UakbQWx3ShRDMXjPhk4C4C3Zh1c1b7DcntAjAkKTmQYw9/Ie
da4qgwYftVoAabRi5xsUosy7UU9ClMdD+2SLuqBqf4tHKT03RTXiJcrztFAhek7C
+AhB5jPFUKiqRv3VPNjvZJQwdxM/xGrbJT/ct9WnguoN1k6szmwDlOuUG9spDs5F
7Q++c2RKZLwcHPFrPEiDrFQxuvehRcfLtDEmCPBAJbAobNi/akyxYgPicJRKQQWS
/EDypLxUuGyy6HmOL6brhqRqsFmdFCFjBEh7j5PffAgIr6nRx20g4dEKS83GYVbJ
o033EbNl22ZAovZsMDgiDx8iTJDNrMP2ujKqlx7gi8HVGvmMDP049Qi5NNZSDcgk
fI1ZyHuaiSLziTOgxD603qpiFqXQ3UeZE1vXlD4x9g9bF40wFvITvx+KgamFGzdR
WbIGidHwPOS4dqOWm4eumeyp2oocq3InYny42IUqK7oL7uUmw7k6inX3WMEvQJvw
ja75oETSeJuZ6X2MpyhHMHCtQkl/R52hOrfAHYzSMvurITmk2iCxbi42qTUkf8Jy
kd6ZaXVk6nR1VuI4swIhghD66JG3XhdF7f6jBlt45U6ZRAzcig2alYOhTt77JHu3
gThu8oRNFcV5ilOE9FU6fkN7jop8JRmUZaIO0CP/U2KhfRFlFt7XYXJ/b13ncw9e
8pgNHQc18C2l7nucvtAEu5DVrmoU4g2+8RKr04ffy3blPwBPAYmOc12GCV+nnK0C
fATdcmzLJQATdW8d93mbFvFurbZFHfXC8zcRwka9e3UskjjwqNmcZaAMloTU7U/y
ExtJsZcq+4wp+M4kNP4/K/fzf+2ih3waqAfoRNZfB9QsErBElpTHtspHd+vZsC8p
CynOMUCWszKovcm0sgu3iwlJlp5Pss1aW8ENasbDY+oSNzc7d5PkyEuyZ87FMGkA
Oh1gD9ZB6aie2w63L0WjKK08+LV2xTv6BHt33sNl0CVrmiffAn6VjL3g4Mls/tQ9
FOEOgDiJ9Yx5y9Zt7Nzi0VLLfR+ckinPpLrwbWR7Xzydbmasi7PKVa0awUujaYHQ
7/ChQxYibsYLs6l+Z9LzqA4GPecrp6HDsVPkABSPJ/9zFywNmF1bJCStE9nFZv1d
ETScKVGo35aFsOYH59um6FFFNhSDu/vbhpRTp4wi5DotyWx/iO1Yucwp2DtRIXCS
6zg4rj2celPtR/pT5zEPH9yNGxIEKpC8l51MURx+M2dqz5FQW2ofbq/BNuFMGiPk
bJZxYievKWu62kx/gnwLtELlN7Mq8dEYimI78/+yiw0OLKHA+8LCGDNNgW2XsmpN
qQdau0dFAVo7YJAdD826Xd8ekCm9/b4Jkm0Dx5myBkHlRl71g9VeQjNnQcSuyWtj
a+3vzKYadzSgIoIFcRNe3/5g3jQbFMC9xIAwfWFNt4ddIirE696TP9kBSx3qt8kY
9jc6X9XD8RNtJgUjXd2YgOIMU7y/lbOJJnnhTUe0YbER6BUx7KfRKjP/QvjLErNq
FRCk9vvgINOATKF23XyKFr/uVBbEfPFndQjnNUsbpgE4rnLpFPOnE/gUvnJ8+EVs
6XM/yP8pkTZEbneNeYzfX+G83fQSl+WY7z+5uK2cYA0B3zm+5V4g2uZlw6ffrWXo
1QeG+HtezBJEt5SD2CBFHWygh3QIF5uwT1H9Cxv/rL187i7xctPs22GQ2XNi4K++
4NVoacYStkZF54U2Zj2mlmmkoGWTVmtxkY/8AFF1BUR7mYeNwyWnUuo9NiMvNDns
157Ow7Cn95KLf37H3eqhfBVork6X53rP5ugiPcyy+ITAyFcff6oC6D7+ColWG2he
k97dLU+BGWRRc1Xy4BFEvejTp51vfuChuX7G2cMva1QnBjY6P65qlnUAC4RsJSZg
m3r9+oiH8AiiWoY/W9MJQwlRvpjKkPpYgKFK4Fs+Pp3DMUNgT0K11CMKyjNgPjmk
DWsds0KMVgZySnGmlhp0G7yJqCsPg6AEtE9UhLuOliMfrl9vOR7WHL9oaslZtcUA
IOAMsfMXZfxGHZDNAcI3/Vf7x7tG5+iLupJK24gsDpVAGAsW2SyOBLqeKLAz0Hto
GWJTQZDwaPOyIHoAemv4zmWrRL3lSs/WSeI39K8yP186XwftmGhb2ToEb4nCCZAQ
qHn3TYaQ4JVN52On/L6KANS8fKiVLeLNkpAuyoEqmOhWavtWIEbHfOgrQzKKI7O0
6kYk22nUubbIYxtYremoWn/YdTXhU+nn8Jufzq8ggt7qjS7f0Ua7vtj+QbZkPJqC
LRWhQ4tUVotnHozmrLVCkaSN09YT9odZhlvXVM/o1aMUMlkyM1P+ZOIw3wdU1m6k
VR3WlClHEbwujdXe3Iranpu0anaQkcW0tFkgz7uKglrfdAJdsoksUsSHf9I9DKtD
Hd8n5upPu7Qqq/pPBgUO4MEA56d10F5t4DPD/XL4PuxSloNgwkhovqN2LsR8j2oI
IUCAFm7afENj8MRLrBlxr9JIlIjsMmKKpeKiVJXvW7c3PF6Ss5CEc0UnFkAxove7
EvB5QBes9xwqVRLAB7UoSShWargcjfia6hU758aMIFvOTTLzGL4QOoZ/M2CNoM6x
pPTTr0qR8dzOtDTAteLaDM0FQ0FMY5IH0ZZqtoHMk0PdrahQ/XRuYHkseRIU34FN
OxsOdZWR27JoqUxN1q/qTdtPUJyLRAGsCMEMZXNVTtCnaA1taiI4JI6mM7wV/avA
ENW01Qn6UmKOrd2IYkwkn9nAWO1xmjonNNyHlfzuSkvXd54A19Nb4ziPpbcbWS1o
1Z02rcaZOskrgwoeRXekBOXKGkn6E7gOnJ4BmPuASegXBZ+1I9JniXuQoqf25U82
h/o+6GGQ0+v2CFa3Fmw5FV+EaR2E3K5X3E265dMNEztyfJ2ibJ85A2XXHNMI1BmX
4JGmaUp0VCZ0zzbDju5RxMr6fQH0XV4VdQj6iNpp4L/EJ8TIf33hgPsPeb2LlBn8
z2G8HxLXrLXwf9IV4F5rRNrY/w65/Ne6fEhtYNm3/iJwZdz+w/v5CQqXJ3Jfw1dz
IQ6mKJEioEi0ZiM0q0SUEKr4kq4dWE91EfEeXx06/Uu5cNCcfvFb+n1oYtQCT3lo
uJrpVWpylOH464+H1Rdxu/WIiV0pPoZRJP0W7QG3TiEfiVUQqIdAMzOaWB4WimOq
5suNs9Eg0W6nkXON3ryyKHOz7X3plkH7Kl0iSq3NuWYFuQDSq2HkTlNUScpS6Znu
t3+u+XaigfMKxC5NGgeI/L5QkYzTC7Kr6c2P8kf/hIdiSMcMqN6T1MALzUz3AtFs
Wp+vwJaNqGOR+TSwcY5yQoAc/sbe6WTuBHKtHniYXr7QU93n3N3Yv/MKcdY5O4qz
baZzZrQNZ/OasCIjTzo+7rnUUhLJDAcXNX9XTEijvdtAjuF6n1wSucirbem1Z5iC
dRuR6RVzS8R8AJL3M7UJz7QFVlQsWXhdbf/YFtRo9DtzACHREx+vus2mbp0RpvxC
qFzN00qCZO5rB2SMsIgIUFmvZb67XtjY10n64zsQ6ihMWcAbZQxPYKFADKPCjbSV
4ls4Ph6nPiqApZYQuwOpSbtTdFw5BdO4MJk04TWYQyNUqeuO2aFuLQu4Pt70ZRu5
3K2MQPg1OMWpYg1juWvfb2SZuNEAwZ1YzjOJFo4yyhc4ROyRseiSL19Vg/5Hec4k
SfarM5OjhOqG/077C2DXu4fDpAN8TrSetgSIdn64YMEANO1hgQkAlK15lnBmGQ9T
Bbh1f/qSeybpbxq2VBZPo1skIWrATzB/KJbos/nFdD2aO4AdhnhFJ3+PUco6/Il9
V/MilJdfXdN4xFxZ/rQ76y2hcebEpSFRKVzSdZmRjCI7WjsEtgiDE7AZjN4ExUJ7
VPfCLkJlWg28MfFcdRglmVO96HjKF3iSz4Jv7TfVvqjijPI8F4b4ds2/AwIoYIoP
/QJmXzo4IdpXoIvafjj9wKCBfdImlOeygPTuTh9xrqKlVWPeJUFcPNIh06ZXwyVe
Y43BOUhgfVUY3qEMetotG7YFwn7kMqMLQtHsmkvE73pAzVirpUWdFDY5InZ9S9tj
IkctItmHj28bQk2K4x7U+mTCBvdMn5SuXS3nYjxdjypi0puAiZlDLR2NsBjPfhs2
b3OxAQd3KT/8ubab1Mc0gLQs/y3MpB9LvrRWQ3Rrw4auqESRb/FnX38eGStLL6tB
ORpJKvcRbAkzb5KwM8kfBNEC9yEoNbPXMEh6AjMrJObe99/7k5Xyjt+pyTt2MoGg
X33hxUXfpIVZKU/vNywJCuVgh8nJeM90mlRLdW9z9RXCSK0eMDHKWPEGG9YSBKjP
J/VWk0HsA2Wv+xiOn8sypamXF7OEG7xcwNknyDQDOh7WqBll74p+BCCGOgIrrQC0
giwzIfj0EE9Z6L+pzimsK2XvlN9YhLauGmb3EgpYKilMusUkDWxuXdZj5GLMGj3a
netsJK7qZ/yiVtyehnan1Y45xn7wNd0pNGtOenhHwi6rpnNZRM7m5Fi7lgfAesRr
gRPbNmAQncp/yQEDMuu+ooS8UMshPti7wV9T5CT5MUbR2v7gUr1xVebsaXHrQ9hV
YOKRLaP8r6EqAmoNsa2RYiPXsb7RcaWYxrNwrRCyv4aDqgvqNlRVTFg+bMAwQpcQ
GDIPypkxQhwFaumPyngxLdVfO53E+ejfnFnxSU03AuaSsbgFWvn8tZ7L/aVr28m1
KdYi1UN1HQUb+TyfEaBoC9y8xksM+7do+0gA20/6G1ESays6ZatZp0qq7XxnKNKY
76IsZvdQu8783PkMWGMviAhR2lK507ke81Se1Ji3yHkSdysdphjq27DeCMBJo7GX
jGteems2jNvGtuN8h3fMzNs0CKwlxmkNwahLsSuS1jvhbAzghmdNqWpCENolQgbe
3awxWHbOrp8DwW/mfgqiiYYNUl4Qigov4VS9hA3+sZJtrTbEo+TQyC/t6nvx6+7x
dJ5M9N7udDDY4Or49f2H8WepDkkq7fYHBn6Rr7o26q7g9WY8YN/VlQVJQsXBE/aK
SXxu+7GWVE0KCOIzlwFmtX5m7brY6IJ9AmoVde3yP6O+Dw11s97ozzu1FwjSeuu/
pGAZTma7qZ+8E/UB6wjhU56pFNcRjwoEDmcnqTdVjUFFfTx9WPbnH6Wq9b3Em7Vp
XFR6uD2p+Q0jkqJabqW65/CgL8/MXuGHWB9j4t8z5xlVzqpSLa4QPM3EOx3qJeN/
g6HPqqcb9szdEdN+3M8xZ6I6QMnPUF4GgFzmjhXUMzZ2RozIZx0pYhV+b9sYiwTo
ebPKbg1P4wwsIOFZbT4MaFEEsbKwINjvDEEPVA55QeGL+XjNIR8Rkz3Vb+XdOdBq
GMhHUq/ynp8JLdYtGI+kHR6j82x0n2MqLbf+brUrUB7V89fWfnPg5mPZmlLT6Xs1
xWLHa5Ua2NrD2E5RRRydmqLXBmpdWFKe3uL0Wv6lpguC6MWPW9QLPKKfhZ4K3lPm
K3cWsikl+BCKSUXDD5nPF4e4B0cA2uPUnvZTbYLMnEWH5rGVG6ovIqQqrlC7SSbX
nm0s1HZZnAbKJpB2QMUuC5j8YHubMIKVsnSwpl2VL6VKLI8s8WNzwGWuoyhnpSAy
NupLfXTk6baSeK0bEKbrNgSeqlAovIJz+MlBoX14j4cxPyiJl4Lq5mU5AaB5524I
LE3kkzrNrGyzQXP2w3qeGbwFHlVzmIGwZHOWrfYGLQefzRd5IIsVFHyGmMMR7MuN
DoaYcjQvjCmkm2HLm4Uk/gKYc/9KMrOz77uE3x9+iUQQoUnzySvKqc3AIFhj1waE
4ThrHJaVVdKR7AxCzKTHhv6s5ua/qHFMYDfbbZwQJgZYaxY6XiMLJ0B++hr/p2BM
Q+Ko2fRY/bl0M0GLbufrfNsTTP56YKQH1JA0dtFnvNdYJ04MqfdXsztgHqCNOS+a
IafMqhGYfdIdaV3A1JFxqjX0FoQREOb1jooC7NDYY42lJQJ44/jCzjQiANaV35Pd
IsZfa7MlJCtmyzsRbu7Js1Ib40Pxr7AVosgzz1ISanaC6jUHLL+iaYNipaFGOSsZ
XYsjQvFUqFxS5dcofJnKWbpF7IMn8DISq1Vn6x5wJHrcaRKh4Ek/roFuOnnYI42L
8jaw+EJvB6R7b62cQWuCmJP3IHO0rywEWbjFQnOwR1Bw35/Yjw3vZa4n+xQEMJsB
LJwmzQaOpVC8rSF9xpcvCf3H1mudNyKgjfdr6deJSBHn9hlpWTNpWQKFCHyDBK3L
LtRI3sLAPjt6TERUsC47Cp4NUmWJPSF0IeJ6H8eW3jl9oHExsjAriBLKDBtd3rPw
5UC4TkraRqxTohqvq/5fcYVS3nVSjSe4MbgL1vCAOXxMOl7sYxCAOL5iGdwgmHwk
5qK+nPQ0H9fQOu1DnAj+jl8Xtfmlv6k92JCIVhlCmjpKsMumVzh16YEdsA2klnJK
Xh3tYd4R4vIp+jnjFgCUI2z2NRo9vE4+kblkQK4Vo/JN1PCLGOM7vNEwz8ccQY18
bTsS6EKh/HVHVuadOvV2T9+JLmk8jnaXcMF7qzBlSJM1oFpMNfz7Bxm0cxZdHwuJ
dTF8077ofcT+Ym/MYrUmRUNw9pEScj1xkfDebxr2tKtulcSZSt5+Py8al9rZ7cVa
ZoA7NqP6X9QP5Ryk9MbVLSeFKcKOKkWQwBSdAgQKCQoRLXqlLHbk7VtYBEG6THbP
v1P/JrCTaYe9ONzV+vstfetS4WiidPoDEcLfojD54xCBSr9shG+Ru0cZnP+KdxvQ
vyABP8OR26rwA19cA2C7Qe0OEUcC7iuEp2TC/okoQpnKCIHb5raeLCvYlhpMhCMl
6e041PrmSxqzd/O6Tu2ZUkABGQy7xiPZbsZuWmY+7ofIxn6oID3lPUDan/smUkzB
GB0nIKDZG9A8Cqx8dx+Z7sm6vrCM7EcFhoBPKrEajm64JpYEMtgCEH8iv6bb2d/o
SK5L3S0Pl8zmUATQnwLPso01uB7+XF+8+RKKxWwnQy+mrAb4/6xK9A/CENPtEr3D
qM9zumaoEP6gZiz0uFQ/l8Rteu6vgZf5s25n1F7F0/X8r7AbIAF6GbxS3Iv/VjkU
EIgGWgc5sMwe+XqSeRVZnl7ZWAOz7l6/Lb3JMugYi9KkFYt7i2o8CxTWse7rnCQV
KPjsEye3eKquHhaU24dKBY7cl8ixZ81e2LxzuTFUPpV8A+lcLQuDzJx5SaRkWM5s
huoom3nRcgVe/upJ68TYKF4dguD2yDE9CDSfZ8plP5L/BkyGzZd3Qox2lEPKkfxb
0YcuE95vFSdKkGVpnia9och0tC7YTSWHZxXmP0CWtM8XYoOzaq7LLeZocQNV1l8f
PixgJZARdRZaIyHou1jSfwH7JLYDFfibbO/LjP6qsJVj1DXD9s+Wn4gKhnOM0Qmw
miFMFwODk6fMNAH4qI7tmNUFTyPTzgwsjpzyjRF2rxcXbbf6LG6zCxc+9F+zXqwQ
N5BkSElRQt/x3ciwySuM+9iy2mSCuwqOJLhzrbUphBHrEfPg+6obxHGNaHWyl0uH
x6Vk6LX8F7IYmOIfxkLKQhU8+C7JrXQ2NwgBOXefhNSE5nXIOQDJSGIJwMy7UaiP
D0C7gl05b2actqUdttDe3oX3icLUPPqIEoZURjBgpr4tWkpC//XOcDzndfjzwAPV
F1MmukypBONT8O/x2Oxsj/O67ar9l/8+X0bmov6y0CVoZKjMOYyrWUjluIGUKz/E
Qu02WzC8VoBHA9MVyO7z1+wfg9D1czVUDl8S8Qj8/Xs2/r1Of+Dpoi+RpFASPCnO
Bt7JQiv9yuzCX1zJwV/8K7i1y4ZWEM2uwT2dD4SdDI29xk1LEVOt8MxGap+53y3f
QiL9XL1f6VLs0fcoIl+ON2XIuflRfFJ1Q2ijigKDFfsb9fwo97j0wt5PaNMrlADW
FbfHVL8D/vAbdzSdrN6hFYwa3hyO/idBUoGYY9VgFOl3mF3OjCFLCgbEjRq9KaRN
5SrMBJ35TQPZy3osH9kAHBT759O1aApXitEiw4A/b4XAv8evkLPC+TR8/pYwDqBA
qfPzDq2q7BUJSa1Wl9kCQXErqZ0G6dy1ukcSWi10o+eToj24X+7kGrl31CVJRRgP
X8bZryAOzgGxB/m9msyGwamF1X82zpb+pXzT2kNc+2Gdh2YZ0DVoGypy8ytdGcWT
eCXTq+nMjCBsJTuSaJ9A1KLpLaPkxBGe2NBG55irF8Rf/FuzToOMq2BoY0bIYCqk
caWchL84uLWy1qpFNsSu0I0aTrdd6uz93kb9evvffOLCn+ky0xmJaeeHn0Y7NLkw
VtXJ7JviRIPFePd35gFB82V1C2wbDHMuuOpSux09aBnN9vzUrs47PoAxhu1Ljm40
n2CDznBRJ+VzUC9XxiBQETfK1CEjfDYl4mSdEud0Q8cI8TG0ZsjFJCZIIYzABwgW
B2IYWUVqHSLPFoHgGQSABTiiZkNr//NIR1TFwNtJ6wJiZSnabOsLeiZvwtbDxT/3
J+71szjSJoAGS3z+NOB2N5JJms+Lldl9OIpmwl6RsLtaBwv+WDbBea1oD+QOJ2Si
5xlyG+6KfUT4V971dYORxsHLAAFThRvq9pZm92oh77MPGbsw2zZvGoz5oXq9q2sI
dck3nLq0lRzYCgVKKMnyuEHiUzB66TCRWfKFlK0MAQSJGdCsDecoZmwKOSxsrBmf
0OQd1cl5zcXEPMhq8NTgHpSwMPsbPymKJ8AtyP9sPnorT9GEv16VePpKnT3iCG0t
E/TTh+UGOXzp0bMwrDXP4VoWoR53OoOqHk/23RahthlidAJxCb6TZVmPTbRuj4De
tZGGFh6JlnUSUQYosFuzUWDx77acQk19kKyGTv1oknzBPgt9Pl4jVRMrxNd8F8Qb
WMQiPWIE3LRNcgvtiMnJiVKM+ME8FDACHBreBT2N8zJgwXo9pEo+z/bOfF3d8PAv
u4Fr7ajTWLrT2yKRrVuKzh9GFg2bD5hAiXx9UFeQvnp3GSYCgxvz3H0tLs5tyfd/
1PUR9dFhuyCGucguAMZxKoskHNV3yqn0ubCD73XG/mKx68TJXfuBVqnRU97lArKm
YaDtQ+aImHmU8AL+pwjUXragXEhsu5HcOglTdHNWQoYNuQbDqzuZIfC/N+zw6yxb
DMTtIpMRtMnDMNHs02TveGeB7/do+kIxSs+iz90Q3HqG1pndeosVZFaorW2AQn2G
3mCvv2Z8ncR1WbIQPepwUTY4xnUkHHahAvtk4AWBGbVyyEA/iIUIlR7S3Fo0kTx0
MmkOzdw3BP3wFLCesh+oEcN1TPU7/oaDj2ED6KkpOc8kn9vgfZbwSLxzDPNOQ0V/
uKqs3zArfv2HLwXfDDeFSN1wrZaSySZjvpgFM6Q5MjG6d8rj1K0/e1VN9aYAwC5l
a6osbR+8YONM1Tef6PLj3hxzSJ7sV+B8qnemZCXVmxLGQaS8Z/92jRiDJffFsq83
P00oKszbt2EBAqUea8lWhKdPuMC+Nsk3oPeUvz5RlEZ4GYnRkp7SNU+S2D9aeS5Y
iQezr5tBjlZs5RZJM+HMTntk/2yvEYk1DLvLnsgPTtdbWt48CluqCHMvJs1rJehK
86wUGKYKX8zxhKeufziXqq2eqBMhyuzhNJPDQfOCDmb2/jfMQLh6toi0NUiAYrBa
DOeK5jQZ6x17SkTdl65hHBpK4ZZGPVw2lhgmvTog5laNlHUiR/+q1Yv5TVvLemPy
NikBCjI7MD/FOPSUQpao6g528lI+nXXkr4O8nqXbMWPbdNsgipNoCia9ZprQG9Aw
U1DtQpkUSE0JaIBB47FTnAnsl0Q9A3tfySTS2sbWEqK5Dz/iPWlw4m3AfBnCV+V2
pGepiaiczynurKQrmIldm7dlIAm4Q3FpCTJfSTqBI9adPiOnMin8/laBUhaL3yU6
RBA6tB8i+OErsOzo2ABH6fjT07Bv3+92FioynwBfSxI60y5qTX75QaVi++zpenV4
pvGQt4iWrhP+Sn+h/YJsoWRYXfxUlKWSiVcOt8OoUgYtP4yvE9Q6Y1eHLTsXzDrs
GnmokNyxJXQ/H/ThoiVW4zV60MDhgfBJGetAkJU7heGlMDoxPKOhMFI4Rg/BwpwY
hxREC63ThlTPKTBTnWrFAkgvrmETsLEWbcdgiPPXcadw/9btpUB/wyfCbw3GFMI7
hLOjTZ+CnvWsmN3FNloshZDHR7R98wGom8A2umRt+u01ALohdQB2D6xrpIsn/9Oe
jiCwtT4Ggivj9CpNjYx04FM7g/BiCh9uqMBAiZdzZUaV9O9/j6LLXchhxkUFOZQ5
OUyLJ9owDBPiSI4zb66MUBwkTpFXfP0Y3rrUPRMnC62mAO7cUQL8y61Z/IS2u6i8
O/yeKECAicyaPQG0AHl3hB671yc4rreIMyTS2erZLNfmCFsFVZMqN/5eKmp+E19K
Us7rhmS9EtAb3SbbLrjHI/kBWpWBvUwGyclDCEEr3HeQ61E3afnrMhywMd6MEFEX
rl/fW23m8HkX0m0JtwuL8BRJjN1PrLDQDOKv22+esao/JVawACUah2BQDd9YQiqC
6yc7ugOF6jVQapidHqq6u7q869AA/b4mvLulIyEQlb0iYiUfEvKZ34FptCm8XbDS
KSOASRgQNvis9vWrgMSaOOuAaGhvIMjcCN82YzEn03KOWz2Jj8hVssR6/icV94Qj
txjQlf6GM970BgoCIlIJxfr3FEZ/7sEpmUrMeI/q2Y7xJOcQujf2iYUHAkqlkCy9
8xvigwXC99IjwzqZfQyzXlx4CR9v9YYE/ZLpHGEUVWzdX48YBkU8/My6yrpVaavh
1iC7ywo3jPnMwzmte2Lb3thiIK7hcq8iLpB5U8nV5Q+O+5wKu93g2uOjGJ59b7wR
BdKT2ryLRHop8vwtDxhG2TOE2WZoirIKfBKLWzL1mH0Pf2Wny8Rjh27Gdi9zJ4Vt
xItVjYLQgptOjNsaxEDmTT0YT8rOx6TBaaJVcxlF9e+CvfjdG18IboeNs6PFDiwx
Ku0i90zgVC4YOeCVZlXYoFKUgrhw513unhwKio2bFS0sVbsRWpihqQoIUaZWo8NL
cGflGYhwzEwRerWdQQAg1ty9dNXP3pOR2nx8Amdgpa+TMyrlsAsuHRt6RMpnT87q
ANUAryipk8wyuFrell3JEPCDLgFS8S7G6uTozC6A03yZH+gjsJo8GZ7vZP4wn2N9
TqAj7vJ2LuwZQxJoYV92fGFuIZ2RQ5c692x+MmDlHA/NXCteVxnEtY7trOiGb8uk
6s1RT+aYZYiCiI4Ljfh7Vlj6acA3FcdxvOgPEev3ObiWeTJBi2JhPh/rYRsFm1E5
Uu+2FndL3McmnII/gb85GRXAgCzPWOUs0SeHXDQ6HaQpgEe2DrQ6G8voHjmp0RZI
Yh+9LYm19OGJLbw5CEQknODKaXEgaNzgHLV5O7zOxxGEa9kVGHPmoOPnbDKrHN53
x5T+MsO4DwHty8iEbmZ+WdpEXe/rigOE2yIKN5BU7jG7Eq3N5ql0F5u8eN88UkSG
8PoBH64IEBDQAp52Fk+g+9K4XQUZ/mKly2E3uC2oN53sZcoMQ7+yAOTaSfGX7StE
0xZq60yn2RCXlbl2mlMZyjwj4IpKRl/WmvCBC5U9POlIPVyJ09ogKm3VII6NQGnz
aRZCifvXfEnCDoH776D0HVI2QjNnjxVin/R722ZhT537ACpSe6KFI+3EUMRbWuuy
TCUeO4djsZ5APd218A2kwQ9rHaBiBITiZXVjndu/GfkNetaaBL8bVjMvX2/Kw8zh
VyJQCcqwR10BoihWOkT9mWirZY7eVKmp3xCGaKxcxNNsYs/0C1zybBx3WkXzeplW
X595k24M1Qn3pyohlem2UwJGOuMfS9/30ONAjtlCZg788X06IITWH8vikGrhKYeS
deDfwn8X5nmPvRFUr0OVsQ43tDQ8czqJA2x+XW+pH+SNq55P4lEbP8ZZaXNVDg/A
mgxiwnMElT8w1i265RxeObjT6fLMsZBlEUafcbopMnl0X7QND0Bt2SwGLg0Xv0J/
VJhCN9wTfZLJ/m0BpPYbbnMw2xYhYxanqQCsdB0634dcgNpX/xXIS/DLkF0Frxs4
O05esbjXv2vx8pp5la7+2apNMY8RafKLlcIGSefuatILAlT7Xq6BnGediqnexIjB
Wl3IbcL7lt6EjXdKw/Ht04JVshp7Q08AkK6U/eNE1M3OB6v0s8yWFAo9OE9qCXVq
xl1Y/h1ksWGuCdK0CY4IkK+B02Rhk1Y5AcNezDX8sm5XJpt5Wm3OG7+ORZKwrbAh
iZJ1pGhmeXLYH69Q99wR49yC3eVOVpO8F8eEyF9KtgrM3MhZyddHZv/Y5r8kPuRH
/a2xbuOtWM+c1AGZoAa17Jo0WaNDnTCsjNhjn6CJiYLHo/RSD6M+Ea1pTkBa7Fs/
CxPvdY5A3lb/L0T5BOqkDf5HF0h9xWal/3+jakf5td09S3L9Psj7KXMxB6b0CF6V
g/siGy2QLYkc1fcq+qeiW68VULh5KCrJFqd75o5MaUssZA3DE2THhQSQ9s1ZNqR3
yd43+4i6jvO+2Q+d7HnnlLoRKNZNnhyP/NbeYs/7xR83CtC5axDAMcqkiCUgdaY+
DjOVaOIQ+BT53cglMOSTT+y9tGK3OJb4w/EWM0VGzMH4XuhLLP2KkZhHkdBDoFWa
U9LRSk0aiZ5qZedSjFz7RyI3uWgHzQ6zhTFqoZscC6CCSZo21Abq5B7Sb7LGqTt8
pZ2dJ6b3neKGZ1tM8NWvrIykOpIMzGy1FqxM5PHJ8ebCk2c9G6/aYBB5ld8dAYUU
m3sBLnewVrRvOgT5S1eqoH7Y7f7MagTCyPfPrZ3rUPVeyhhQVxcH314X7VZ/Sneo
fB1KFqzaU0Wkwr70zaCvrX6zMSIsk0KWuoiVtHDc3+sLYsWBSrv9r+sOwTuLG7Ka
xpgXcTSGJVRL9hjWpARYS9w9WxMkPmmJGsYF3N6aDEQTXuYvLcmycOrYHGAh4WxY
USGmzCHvstSCJaNBDYyDvfDpBrmR6SSrDp0g8W2pYTa3E9cVfQA0GgmGFCOaFLBS
Dy7UKMaqhYQsu/xH/U2MS8r3W+yRW9kQknqN13ixm9R6AJ1PXetfgrcPPHF3PF2E
xmoIunJyiRZJXTT/l4dWdGoKeQSLtXvlnzMMwgipgWERQABv9B58H606q4Gc1s1B
FmRp2sMl7W80zPCdo42l3optup5VyjZ14XQeLFLX4xov8qcYn21Qr4CDQBeHAEhR
aeuvxavrR3W8D2W3f5UtFKjqIN17wjW8hQMQxafd/zmEqp6pbcT1dQhroej4+pYD
PLTqdsH1yPaLxMRlRE3V85UKaewkJW68c3J5gqDoH8a2aVBKDWnxtPfpoEwl/DfT
2FUrORp0FU092hGwDPFBTcQdQM850K7L3wSpCxt7PcIij+TXsrawHxzPgWCCRxo5
7bYg4HIKIn+Z/eSRSVEOrZ55BidtUCEVglSGM8uTAaWiZ9XXgEpqKjPGGZcvMumL
20FJfOygDnqMKGNp8Lqk2EesaKfzdG9kugXwCtmUfIXyBkp8xjqGmzR/Sax9OE6g
BgBkEgW+HztOHay1Vx0rDG3BW4faJmF1iuk4KXwc05bY5oCn1MjeloVQ4H1a8B1c
G55DyE3xCt/J4/JYmbTVWvVBHHSdoogD+sRZr9MIWawVcnIRp1dqH6y8yD8u+45m
BjIpNoh48g/X8ZvN1rIjRpvsGKSjyaSi8qQho3m9lcuSnXYPueN+pOi6TYRR0nxV
N7AbrtJoPaS7Iwc5BJ2lvDXd4Eg5/1Pet3raDNYLEanSxiMnzRpBXGV62TV/rqqK
KxCZmCz37amydyjgpnhDjJAtO/nqO6GJ0YH4Q3g5RpM99Oz0/TkgbG6MNViRwz6Z
a5fQ66pDJmlIyRB/POy2h1QlQuOog2gIe7MZLXj+MPhuAjVBgjjs1U5++bs25qUJ
OuadOKq1XyHzVngztwxacjJdDsxVzKbRA1f260B8Vr0pSKZZON3m0Kqgnn4aBh6R
AyPKeiQ4b0JLJZV9ax7SCn0Pz2iIGTXX+jZvqacuTIJT2bJuOGUM+eieqaz+IjXo
ePThYeASX6caqSgdjqfEJ26li2ufIyQD0IE3XGzuNhvJuE94+RFcEMaf5VTOe6/U
zfJilYNTC+3w29REHwRRzRJBy+joda/X8k4rJlQb8MZfrj/KfCvpwpW1ynpXmWSV
0VMkR/YEK6x2bSeP6ye4SSDU486nYe+jrXmyqEhyFRr4Uz3j3mHiulfmQWCn8Pu0
oPscexi8EayoFJc00Oz8HN6Yg+xxk63ZorSSasN7WASorqd0YFtK2jQq4gAJHtTE
ZFPva/aSMFOetukUXVJvCiaXWa1Wy//VewsFd3IKb61vn34YNiMkrm7iYqdT8zQ1
nzzNOaA0RQLjzSpDWFliheeXunSrx6sn9+ygl2vaFyM8sPujPguG5mXIPnBo+wCk
osLxGZhgrIF4AkyaNUvBe0bQMyf2z3C7LhVXuWeBAiwAp9yQgxSKebejh70Tk5+6
XMaGAirf1xbJi0K6VRr7AFKmtcr+s+elfcWo2KCuESK+AthWvuTZ23S1/05oeDSQ
3mOq6kFhOefn99mrG0IDs7qI1f0B34yrgdW5kEY8g7p60V/ODnLW3siMPr2nvReP
DB6xDzFBgmkmw8uFP70aff2Zek/Ex7CMFwAVrRTVlwAvmJ63pkFJkreUwH0TpJMM
o8VWGnWMJ9PyZmPSxw+iidh65/IcL5JnOnLzuH6hjcRxaDKuihq6/sjOg4HOZpgo
rK+H+0V0CbRmTrVWtxn+KGkvfnOSvWMVCmHrLI+ddhkYyBZ/3j9AUI1VZvWBqruq
Zd/IRArD5B8ZhPpuwx6XhJSdBbbKjgxT/EtGh+GUBMSv8ohGVJf4lFA46h+bA/KM
SLtLud1TuPCbOitUqWI4WMA9BA532GqN9JOw9JhD7uhD1aDlxEqyEU+Ujx/EG1nn
qgdC+i+mb59woLSdHvguBbm5+ovXuaqGI12aO2YxMUAbSPVL+u7ZCTguG2TsZbCn
qLHueWHi7BFgp5yGEWaS5cjppA2diJFA6bgQ+KPAoHbLU09lQ8CXQDjaV3GGNuxC
+tkGX06nayTgIPlFJbROWLL/MlscIwUVUWgk+cDfdvJDAPlSU/2PbKR/dg77nc97
uZ1y2GtXakldb8nflBBOindxmclFiKCh7t/q1b30oX30c0GLAciEeTPA0/gKXUtJ
9epoVLTgl4BfBHHEBsO4tmAP53cb4PTvHMl1C9w992ngzZ4dLITvh+QqmXGQXQJz
ye8+zXfYXPoUlSpR5rRiRZMAUOpAUn/if9a4NCfQsTxhwq7G6xpaaoZvjcGV4yO+
D1R+s32FVE66b74RueX+K3nlBdMjWXB5YSx0xMpd+Aqfd0S37K+j0gUfhQZI+wn7
lsk+i/pJaz6NITBBi9kbHiZfbLvbjOKh3UaWO1i2yyYtk9HuCeo2aBVoQcRtM+mX
CI1+HDx150Odd9q7gvo7BQ3W1/LFTlaaoGT3ebQnnl6IB0nTWfpImdDOf707Y9rs
ZUYY14lp2A1N5NxwvuNBVCQNzkcD6OcUp1xQfAvjO4RpcWXKEtrW4f/i3hKwauXE
9iRtq0jt8skTIlB6R1UEJICH/sOY7yiCt+IeazYD9ILvwVDHPVQvdhdmEbZN97PN
Yf34GICljyzSidWZv2hdHa5DN+vH0Iz3txd8GcC992wp5XgcdEIF1C3ex07Qvj61
qUH2Rm1WNRq3/Vd0z8jH63zdzWRW1quEQ8LHyYPpUz5qOVjYWfdPIdnDhZp5tvp4
nqdq8XS1XcDXx2RASU6B+hqKdJJ7+N/45dnx+apwDZAF05D5Fwg39Lp5AI9caEqg
ipMrbzgGp4ZDt4I5E59Q59t/muPe+xtLjlIpz5yuoNzqkDa+VflC346cWjMjrVJQ
GR0GDhfM+eAsFIZFLk7TvbWELdJkrXF4VdJZJw6wdS8c1m5ONV36BY9dSK0rOJos
lf27qKthPWIvB94zmFqeTCXOiqqI+KHRfsXCe2pwDdght7k9LgVmb8Y0+Gr/vyUy
FcVBMmdKSxvvkXeHfe4CXjR/g4kvc5rxrKICzNedX+OZhz+rvN1Qnp8/0mKpEJHk
Ddxf7DqvhN+kCrI74327W5P62Jlj9GmYtcriH1NO2KnC7mpEKWvoMPS35wXfOa96
QltdWco5Cn+9TfgN5sNlM5X26XXUcul7rWSJXfYXtasM8wjGUw752qgT8SkcbjeN
SQ/7zrPxq3NWrhUCg3P6bVFzkqAm7qFogFcCVatp08X4gf2zCYswaYEknbXGmIeC
nesqXQC21SukBCNrTw6UNnzdIbqG/U6a0vU8/qUouo1p2BlUP/KBI2XnTBE3Zf1s
0RWcRN9DW0jfQCpeTMLTi3qByYo6WQrEaMJd2KrmENDJs+k2Gt1jd5n7mkGRWqrm
GGbluxKVR6Bvv1JU9j70x0JrU56MawytKqsweTjpQK6488XUrshoS5MJiej0q1S7
Dz2SUObSMYeiQbQ2e3GnPbjFSAUld3bmNKvOA4ogsLOmK6Ij1vHNVXInDtomrWZf
eZCzQeszez3r/3nlYopgVi/AtJ/MCBT5Bmt1qTB0geSaM4jOC4wOOtIi+li1c80k
V9XcT/ddY5pLcAbs0Ye92rj0Vlg8G+1q2KTp2CJ+mtNBKhlT4MGgLNc+13SA53Oo
eA3b5JMLLJMPYxlrdCMHmlzGwiF77fmZxBeiPO92LabKpR26Jfv6nM7KA+wrBHc8
6sg1paHa2uKGOwk9gq/BqnQh1Ta2r6vw460FgUcMTqcHOeXgGpCUfAwzPD11wOup
v0XX7Yb2/bUph6EfKhuOex/mqYr5kFsqsYuBDoeYQZMTX1hx6oOnIpnoJDjR7Ekl
V1+td5jsKPBHC5k+Yxwkq1q1XAPBK2/lUXZwWz6MGrGJP702yuIVpcHDPNGXhHN+
7AymomduEqFqSHVOBSe4fHez4ngUVTY7jjyjMTFHb5PnZmTDYGM3yHJ+AAu0/Cbv
d3AQXugeQbRyJOcYCDzXc/JSxF9NNEA7GK06Yt2Jm5EarHBE7++Rz0oLxpcYAs2Q
8OLkprY1Px6qNJq6BJfMfpOg1i7V33HbwQ2Xt0HHWfBUhLwB7ilG7R0u4oj5lDbx
jsLAnRV/e0eTizLFlo2Pnk1/EHHfpUCUJozKdksxDes5shF64kQ24B2xnPkWEPpp
y14YEpVHQPP/DGP+Hj53sAJmZCru3ahUfEwIby6fr8/jyCPUOTjdqqHJqG/VylH/
vh3vc2RYqn21YQU0JpfQ8GU5HWZ9hRat9PffaLi5xv5s75En+tf7JbvwnIyEnEMC
dDxCW3IWrSX9tVyaqUE/4Jy9HnVqL1A3g/14ltsdXF2ale3P/4dKjdlht+51celA
5N+FqFcz+VJfNWhiDnCR+oqZn76JB5o6uz/yT8xyYG7yi7LCWTivvZn7pR/SqtKo
jq6IjAjXVWOJhol2yV/JE9XikYW4IoNDrGbqb4zFrKn7d2lIKI2qSQoZNj/rglpk
bKoo27e17h30rXWD+rHf8b3WSgDEuj9Bc2ziqyw/YCxDk7NaFBvxj4g/GlkHcpaU
wcQlYCG0BcRvKQFeGrUH2gdZgUZBSbqDnpJnPQMNNEcDr74vf4Iuku5dhVE5eY8Q
n5MBpVMrQOtPfg1uPh8BiBecBZqKl1lLP97LMEB1F2E/mBqrEszkTiVQHGr4yJBg
xKoPy/4AY7NlsZo1Si+9xfOxC1+HN58ggoa4kRItFnBLfu1pGk6/JEv2Stb+dnlI
RORd2brV0a53gdy+/mfTGwd8wwxCCVV9Xumbkj9swP47Mx4METdrF5XIMpmPN/W0
Lj4hGoBxt9vnjI6QEhrZksf96V0u+T+zi4nbWOQFUHaq5E0yBVe33HlatKlUh3Ia
QRhVl2XjqtnDW1KRv65OvxX+JTl7WghtUYLA91vglzQTTHX6B9coESj+d2OKap2C
+hysYh3GTOfmkfeVaUY29STZxpuyZOCSxoiBk04M3RaAMYE9VTQnIfr6h4I8vNJm
CPE6rTCgHhwgcBNO7z+k2Ew5yMqyk+RNm+AVyQlVR59LnySlrTwaXLMOog1xLPgm
EP3cOGuaYWzbpFtRleAHCdj6j/oz0H5sf0MNK3U36dQw/lzvGTmwfehZNkx9UZ1R
kN9SDyS2J2+k3tITQI0TBD+xfH9T7NmtGW9b0VLa78g2DTw+Da4DwfgMLGcdxxgh
TiVnOa4B06dm+e9jfBLBbkv8mK65k0wMBc888GbzxSWVlUfgEdgOrOXEK6JXI7OX
EzYmkYDCTKwVUcW1tfA2QkbjMdkeK/x/QfXKlOBKp31GAzevaGw1XGNTmro8XqJW
CGGlnczePj1Ng+B3oYjfkSKhHYmCb+gBat9x2FySdF/jbKtwX4fnYR6skf0WSbFB
TGM3gs82AS+9NhwWqdnCopPzh3AkTv8A6J2b8kEDLW5FgzoPPbjgKN2p4jIcpecx
yz8C+CvQpNfYo0Kb+8xWfl1U7N/L3R8HFUEfQMBOxmkHzTFQjXC8vL0X0yhBqg/d
tckL93itwAEe1aUNSloD1cuLCwkpCTKlDi4tmdOXZ69hjG+y6kP/N76r/oWWIct4
y4fbA7a8Vr5Uz4qpWqz9R4kEbhedSmeTINCW2TKpZQfbCrHAjq1NRuvVvqGWR16K
UnL0HsFUDWPFj8r7ZmcYzC+3GX3sHUkli31WWFHiF0ZZ4kwZHu4uPoITqnFQsgTg
5MrW5lm+6j8dvKGwtvXCVpKlR7RhQNtMHrwc0dh70XUzyD+F4ayoT5tXeOLnXUXx
JohWR8gswYdUZ/bUPWShLAwomJBSb81N98kwlR+7ZSXkXHjxKJBTBiZeHj+bllfL
L3I8fpJcI5AaePumjh0L1a8pWciHTMc9+AyBFQpXwgF+M9IJj+BJ37xT5JYFPK/F
lo/W1mno/uDHrn/vpmAXChTkeyaVDxKNp0Y8DjYVZfqQR5gusMl4xIJpydPM99lg
m3OicdKdx+pM7k5ok1MC7VUHHboBe/acjiMKY0ZNpnBKfgLrbTbcnqYfY4QzS8Su
80zvv0wDiz/QFbsodmPVDA0KzSpJGcvf6AgtmXiYrpJyUk83XXX55slkPY5TRu/y
6r1HeIEXtGqIHTYQcDgEE2G6y9SUY17IhZNqa7EW164+T4tHSH2EfPNtFXtxGr05
I3IoNHcUtR/Bw5CnPsiSO5vLrpcwiBGWCqZ/+kSErzCw+3qZJl6iqoMw768nbmkV
m7uwv70kseKYVwyjR0LRLXypouDR32yujBz0Eq/KNj4L9jabwOZpuHvCwXf0vCuh
Ppxa4irTCt5RnE2K4gYCJEzOkm92SMBGdvsKKZQi6R467otEfLWhdbE1MmwnCqeh
ocDmoGSNFnjdAu5jI3k1eWJCcuVPseJrqT3bx86i9rnCbwmBXSx8U6S8W0jAfy/D
aFOR+6wgHqZLM1pgw2ErqV0B4OVKg6JTcihGHVrWw9OdXmfDFYz8tsIgwHyrs/IR
pJ8duPr8+wj3smNZFSZKMBvfi4uITGJZdMQKnIdMxTiW+qGDEAavkALmexbdSRp4
b+wm7GG2Ox4dWsfVtGYTFnRiniK5uNwSNuuiwBHcWFaKdKFbLvlCA0oM5WDHd0Zd
xRs0tZ/nrfUttvE/tBdnzndheXnrwCufI7vH4DeKaFi3DtBE3cCNr1BCQW3C/17P
pVA7OVashOqGrTni3KYe8FON/ETVGO7BK2ZtecxmgZ778HgahUnhvEI6qr5f7FiI
f14ztXsHqIb2+VlcJ4u2ywDD1eWFAPBWx/FzyqKMJh3VcJWyPRjo0xSk01GV+8jz
hqoRyt/lbwf/QzchPyAYn2s4LCDf/kFyrhZrO//e4SV7psxrmZD6QEB21qkCEVc/
qe8FQPuczqkOV0SnnRS+//NRZuiZtWP5YYAKzcnxc/8qAOA7PzMbqcsh2XiGzZ/r
yAe71oW62BhOVKEDClKdlsNLk0tANM3SniMQD9qQtYuAjOswnVm1mxgA3MryhEtw
ieXvlmmWN542Q9GKItmSACLS0VpSh2j6CjcKh2tyOhmnMjIXuG42UtntTSrSEkgp
XgTyWjycqNAa2lGMSMqHrjUNzHUSl4xaC4jhZfm5RJNJzIGg41m3Y5Ykj0Vka1as
ZFII/Gubo5ucE3l677jsBZZYCV6xsG5NOM17k+R+brpnTszzwVam/zGua66drqCC
tvPao0cSYdWTc4UTP4Uoh2m88A4ErEBmET+o4urCrK2jk+xgusEEsPnutCDKJw6Y
Mkl/KuTWN4+KuKbHNi7h87cwL/kwikHXHEqQFCUEklHXn1yOFV7XIJDGULxdRU0E
LlKeuM92faZEpLhtB1y7WMJ2i7nt8rDjw9Fxhyx+S+MPCEHFLvt4y69cMGU2B35i
e+EuT2JLPJE3ObGP3SZPZ98DcqruhV6oYvP4GHNiVWwcZ0DUe19GzrEu6zsmwrjG
FJSTIqp43zLQboVVuY2dv8P6UuckT33s8KvzBMDoW0LEVLLBmgZ4oWpdUjHt8354
m0gn4ie83AKzRrniGgRBknaZchCA3pwqUVLbMW7Z2WIeH3/nDNt8utwKPKG0ljjY
EDKajL43MOdKSJJFCXPOa0J8Gxe+g/zNuOVRZUjvWyxdkOnaiGH0BMOSBUz0ksSS
LvZMZPVZBlQUr3pK/ZCu1rVpB3mB/hEGwNC29gfehzHupr1np5e4O7Znr1j6/p0b
rkguk2orog/uu+Bswqmi/HhGz8Vua+xaq+uAEnUYw14nS7Ih0hhDtLDYwVfEouu0
6WXzT8FGCOSjfGpm441gSrLp8kF1rDEC2/hlF7KKDyKLZrGpeFHTRi2d0yvJrrGe
XDjqcrJVBKOdIlGxzae6kV139Mj54pbhKqxoq6xXIAxZz740Emyfkbrgo1iWRrzj
IF3o1+kDBrgV4ST9lh/Mqr058CAkpAXS8Iq2xkbNafRQD5Tx+Cz7J9Eme6MP206T
heRTg2Aw8wu6DMYddqSPS/gsCH4gpYiiYGoM3FOxJsaoJziazWfmy1LQcoBolaBd
W62QWiltTjDSl/exd96ers2rzUiy1jU/MBP/kgmFjO/dpayB+9fGuSgnLYyaiBZf
gnMjVAPoV1vnq8pvF+45Tgz/yB34r6nxqdSeKnTQ0H3twrwprUvwkv3xFPSxkMEc
kPVojILyH4Qx0ix7IjXQdWpmxaRg4opjS0A4CvBS5TMyJDB3SwiIHpbZtSeLMdkE
KrU5eboHixLtda8KcujuNZtJIhee//60y4qeafYunrtWqtv7ilbfVOF0a1z9aVpT
mcCLlW4DLsBsGtnPAgIeYtXgcXKCIkC1OjhLzmV6DgEdZk1/V4DHljb5+C8XT1GH
cpsc27SFTkzPFHfxLY+mOKTccZfuoBZMDocMrorx9wcKn3tZNpkgCRBRAwkkNsaz
uHd5ssRQ2C+XO3SMwZsTdEWUjP0gug/C4Jb3TDFD8Jm7efcGNeiqxTu/g1XxDzRI
D4UKoa9nDaUuIa1za4JfIGnv3SZ/m+JwuxMtwzPVvHXy27cZxEEWfBHixOSYiTAD
XZZJ9AV8m5JqQejl2JQWl68E/pZFsLCWhwKEJQ8yGwdjbsJfrPskPjetulhreVA1
cqmOI4VvWLD07sUR82hZFVniQTLOwOIschZKTiBb9yHQaqlEkKfLK3cPwjJ3u7d/
Zq4VvHOeUgiSim3wBoZ0I+vVsouzJUbyQow9OqkG2rVRcncG0AmdqbfwO6hkMqgs
fagbPcy+hsQdZjlKG4QI8er7k6EsV/2jhJiJkzGsVMUjpxWFeudKeDoQlJptDiIt
UvjsNzpAEk54w6JYCBidYdu29edtyzTS2fsegE0VE2aJ3MnRH3lb2WUjh99wrW6e
J60YeiXOS9wI9lm1IXwpFVDFYASZB7x3Vcqy6/iVSati4s6vq6YLYAg1R6ESARyC
J80Rt+J2JM6kmNHmzTVcX+IXb+q36GGsjnmhUnjHSsWrgLNNBuWgE+Qgg+eVx5FT
j9Fiua8q8FW4glZQlIu/dIMWXZ1IFkFA6ifkoTILqyYrT0QzQt5dbAXEfeYcQdvY
4ISngyDlgfY3wTfuylxqhCy3yiAoDPukIKOwCbXfJ1TdIhtA3EBQT3KugyqkKvr1
y0G71I835ju01qA2IhIvB+myqlb5o/yY/amCRHfUn20qWr97SfMhk3rTeGl96fBz
ifpTRXDydVt1xbErDyKy6YNOC+XWk5VgAU4OphZlnCJSxL6cHujbap+3ZH8bWOpa
xRNiaAAW6sTgIMUL7ywSDu1ZxmrdWHaywr2G/DZWmE5izDd7VAzpZefSxxhbjIje
QUiLWnlERP0IEsPNKzkx9+GfwRx7OekBlnMnBTXt3mqeXWJNIJaeJCET11mb5X87
qRYXStOmXsEy0/075ING/abLxPEpyIqA/kFhirkPiznfQOe9GEvPkEnsLK0ehRUc
C+Qprk3ubSlZA4DdvfaZM/Nro+fz0ALd3egS7WfaB5eZKuwxyBZAacXR8Br1/7dg
gqM6ydFXR5SKXZ9/09A5HhsmpxMXdBhw//91hrHJ3LC/zWfcfJEAUtQ5EiAorytd
bvg2vY3LUh5EGf5QtcH/0gIUfwT1M/oRcc1JLLpVY4Je9p0UNNOJzdd9ovqIa+cr
e3dDiN59xbJKqIkE193hvXwlLhAw3MkXzFvdfMMnskB9dWnnnnS2TeLzeg1F5vD9
TwnUtj5sa/mYdlTeAzQzKsWqOqXiHsAnVuAYnzmVrZjXGyfJ7v0YSSSA21EdTxYa
z5363vNnTH2pMZEkSlFWuc/9e7KQerR+9orEHhKUc0TuMF69tErl/WYe0tZeUyxA
OI619PDmlcFyUky6W8QSUzs6fJsRqBE9jrqneA22MHcBrLvxc1j8inmNJ08fH6ER
0pIvym9W5/Hj9rmwFNZ6JHsGIzQf2dP6DF+BaSMeYf9hPeZN796bhIcEIdqcjiei
FVAHGy2OVDSjOxN8G/vpPOXWIHDsinUoV+abaLP79bT+/PFBirvV1eSgg59HWa/0
ICxQKqgw4IXLXe210A37BR4znt1h6roLdxFHGt3TItC5qTFu1e8fNyGnGMbH12uc
y6TaeE15A4raDn1WpG+H9uBUTJmQ9rySd89qaACRLz3NNw8ZjzFbfagG1lyE+meb
acDo6wigcOg8awTJlUZ6DWJ9X4diHRyYT7Di2xKU4ijnQsbyqvKsmfcxnVVOBUn5
yzkrodrjOemjAvDxJJCihrfy2Vy/u/6oVWlbaVOW3bR3btfHQLlsQUZBO1r0tQB4
ztIrkFyvlS01gFHs51PqixBxjoCiZDz0758Qo9q2zYeTJ4pjZQHN1yHQx1BVwLsY
f9g1YTkS2QqxcgguC/sdimHim75ENKe1jHA8duZanmqEhxoFQveJ8eT9sHziOpU6
xsTu/S4v4RUEBnimyKGwDSGcAk9uJH4m4Jxqe6IOIhdEfa/OwqCFL8oXzNqTecID
YuWA7YUoVe0cWb79jRPdhZm+FsNAgfvYsW5OedeLYDQAzZS2K3LTrl8WiWb4Yl/E
Oo5oNWiU3FGUd6CYQ1+xUNoibpKRpFwCxV+EUJjTxjggx2Tpt507kxwbtXqEzzgj
Yt/qZdKRXcQLLLg3jqEL7i5GkD5s02GEfeDjmhQEvvwF7V32MBV78cko1xyRwuJM
uGELtnM/pl3fCEzw7ow7r/gKRz6Itrv0SE2v1xenyBaxDaKGehtCqLRLtSRyEnxu
CilD1cZVV1MqYRRHpcwLEfAX+5xCGfjFdHQTPvCsz62sVKCjocP2rbGWcYnu5U5H
JIuJmTFtuZGgm87DkUcg/MCKL5RKdwrxhL5lGY56PSFoz2UBoy4uVkU2gu55w6C9
Z2OWxbMZfP7dvP+P92zH11L6SupC7JywWT37SWwvajgOY3iEpGxuZD44Sagx6DYP
zvalNpTkLzddq6PK0I9CG/qkdCqijMgSFzw/pv4Nl2PWTbeugdGGhbrRceKLJe6/
1IDBE8ontBwG1gfKPrE6LJR07aLB8iX1iF09uu3W9FN3BDocC4Vz6fbVqrQ7zECa
i9QHlOyCBarsTZi/fn4t5qO/MIcGwI+M8ET5zopmnLDWS2aAVKVI9kscVBHdPeFL
W3gu3VIuRL7bC+y6yUxyIRf6fC7CsiZA6OiVtiR8QuWHFoG2UOufH/2kndpwfqAN
aTA7omFVAOhpywa6B5i+P8VcKpGK+SzYxPnZJdzhq00u+kM9wtbxOJvZPNt8m5dU
5lAEpL02pnxhBrKuH3PWf/UERX83MZkpIMRGijIptUzKODz7hCzPzuEx7XRbUZ8r
KGG3W99spDiMZpTjSGRNEwVwoTUsJctg32RqN/DnfVn5DfdrubaeZjuaDuDvI6SI
exmRyNh6qPKgtuzN6/JLL5xGRsU8SNRlL1xNsn08MzpC/ggcEHx6JmVLqalb7sDe
Sa/vxFs+5QmUXduyrDVyxy80Hu1kr9D5gLkwJXLDgqu0RAyDe9jST6ySKnodZarD
SpV7ablyjn6sN1VThOjNLvv7fmrp6lHd9lLFesba0Kah8iI/8Edy7x5vI1F6qsMZ
ZXGcf2+07bkEjx3FoIAho6BnuroCMPsULxbuJV8bZX9Oir7yb41oEhNqCUHecWQ9
4Lc+xrCZ9CNeaTapRr/1TM45SJkE6JHQs2Ro26CvXSpsOHhewyqh++fgN+y9FX+X
Wa3R459AGyozdEVTzCCv7C9i6jZikJFmuO27pvmhu36iGSX5yBMppVl5Qyk4H3b3
wZGfegfdtR+4KVr0/8hl8OUpLxfYK8oxTcJnvCTKQ/ZzT8iQddgGMKuef65CUTnM
FJS8ZZaKSTVHS9gu00EFCyOXhIUi/M07UledERIJk4LFcGhxxYMqMsl1ExlKaNvV
V2l4kcZ66YwEhW8SQEymlElPnUpgymsHwkUIhUatbQCgVnV8YEh2J1QOftLQZQEx
e2DPiGQrR5u5LsaxPW5VJqpxvXLGsTeMRHduuXT9omGzL3XXVPVwj/IoZEQrm2IY
xhYWOAZG+VbVvzOfeuxhxiPnEDe1gAd5pxCKd8AX9aPJXa7jbpEVZCx59Z7FfdZ7
O1C6UNryoFEq4feIEAVmOWWcIEnZTxh+Yo5AExTdEkHekqaJ78LdtpIIY8/1K4GX
f7s5uyfMLAayvCJnEGoNXTp94pWyi9XMfyquoZFPpduHy+ScoH5WG/40oGp4UdKW
IVufzGqBMAyA+e36/ybBNeKbWVjv3mg3PA7FR1OCF1YfgPujjYXsZF5JR2qEVdvQ
UVOIqGnIhPDX211bBS63A43A7/C+PNDh6mPkWykIMGvi94F2Le4yJJzy3J8KBg7M
eRciq44ChCIGGtjLt3jJoo9OmBs+i11u2Bhv2s3xaO0L5VMX/Jr8P8CxA6BcbTc4
sr+xq5uvkzH8VJDGZupF1qpv0uEK2uDIKHtEcYpu1Cv5LrHs0zhyLymY94FW0aMH
bEXZEUwhq/hRbyGLFzNb5avAGs6wNue4yFgAPggnPp+8+EN303SeMbkr3bbKQnqS
KFQiIFP/pA0vVc0Vyx0p02uLOR/WJksRTYizMpnTr4I4RL7gAuQh/utxI80OfQ3v
aCWoEcA+nYSwZuT/q2miayhbh9jWxR1NV2Pi1Yv8M7lPqbAIgg40Re+WNP7gRnvA
aG9YIV3KbSOuBOJE0QMk1qP8nO5f1xsNuX/T/5/pOHka6GKe9ckNXcJ1yZt4stTV
sVxpIdADIGChxlcZzfjo36KQONgbCvkld4OTUoRlz21s5z0IdKWAqb7iuLt2XN0h
iMW0S3I279A4/gPQv+p9roB4Kh4t96Q3w+LRa/l3YN6n4dSlMfUgXQ5piecc982i
kXOCpoPHZhuu7CFLuPkqFhxA+CGFNKTpydPiKn+dJdL2R9VmRilBa/3kOrdy8ABH
VefeuTgJBK3USkGdO3pSIpuPEsPVJgvULAcOlo+gf7E0QzIXOkblfa5iEUr0ENkx
4kvnpqNLeLLt9Oai3xBpieMLXghzG7RZ2rCgDYHct8ZFXJXF0PlsyAHXG30X0EXt
3wluT1Vc2K1dMqm/6u/gZ+DVEdcFLpuwKpLk62MIgCq/jQBDyp/T3cHIRvFeLWDE
M5OpgsndM1mIvShMCek8fnMHmpvcMnxAVMr28kM0T/OD94h+55RjZTBhxTxzlBIZ
FErMXz27daxly7qp3u3uVoak/cWcetZBzaA+rTBXjcHAeYqxtWDLdHkKSl0Yw/et
m4zPE5F5hw+6VE7uR5T2VvG6WFRBeIDFU0Du8kvZ3947C3+vy1gggDXfieFsMw9q
XvsaLyLW6eJff9pieLekv4XfOvKne8nj7xaPXAOjZBf2fj35TUoQxpMdLAiwzxSx
nzlC6ar0Z5E+xr+axx13iiBFStppu0t4ifk4vwTNvA7atI8gAkuui6b0Jq59vDtc
Y4c8ImjjI4FJY9ELSKx0eQGFYbEBSZx4VjGopjlRpQELPDnTxJPMeuIeqX5sgcV9
9764rR3eYgUDHOoECC1V3k1xweOj8GgmHkqF6y1dHWkZHJALGMYXPmKzkzQsdJWc
sANnfWezGjhYyEfnAuLXp//p2yldJjsmTqTyNLCE1l3JPFB175gQxVYPmJbj9mPd
bFu5i+YW+tdTwd8dLY0CNLHgLD1D+xFrj/aF4VMZHxLO7cgCE2pUSzRJCMOLvza3
1p3KrILaWmxQriluyRXRhbrh8bGCHCG1nNvNkWJ/Rl95YGAbV2Li/QKptKxZOL/u
EF4bBqYJoLj1APPzfCFMm9T9IiFr1jR2iuwfmE3s9md+u8oopCFb4O0m8o7HZIzz
/ZHdlkVtzkMkFJuaErhPHo/fbBNDJU/pIE3UuJjHMVCH2QpTKYrn3TqzKSdkiwdJ
mH7AcJltYMgVSJsIucJnM7r+tPq6pZjZ+ut4MSk4PVRTwcMbPWy3jZtW/GTw1x2c
5HJnxdeoiqmNPPAvhhyV09C2QVCGrQLUiveDesh8u0SF86/omzJ6rS7rwmAga1Eg
z/d2rsSZd0sGEwgAkZPv8zf5lRIYFyziogHCXhyYH9IIfBIzn5pSVgnJUir2MM7f
goo6A9kbUnUCdyVc74TX8gc9IKpvuMET9B7c4V18124ugoKwPyODTYYNQ4TsiUPw
56kNr8pRJL3VUdqGYzojj+hvEH+4nI4i+hlnXEZ7jhQHDnoNHk6Fg4ejHQaEr2Gg
2YKvbetNjpIsLBZ5UM5CQxDIunTOwcLS0a332ODTywUDV8pQCpv/2f3z8dmvkaZt
fDMTivjivhvHZQclmAIyuOQ3QVQZ0PgjiXzOwLY3Qy5DZD3KnOoeMCj/vm9jbVGk
npbCz94m6ftjzUWbsz7NWfq3HA3Wk8qvxTTNZrE23ZQaF47qtrQuz8OtnS4Svme6
WMyLSPYcGU+dC/wT1xMSPyxWSHB2PvrFjosGnwW+4SXVNdIgCDZL50mz0yKxbrOi
ytow9xSgjgR98URPKxz+HA2ldCZqK5VU5nXEwbSOsFP1TTY4X0cO9zt8KKOlzpYI
dQOjznrg5sZWOohwaBj4jN9LOjVZtpDJJnqL8sxK3dl8PE1ZeQO/TJ5KpQVrMTcP
ot4csA2iMO8VMS8IBlB2KNsAccBIpAepXW+P7BN4sBWlOppIhPMSL1wfN2dC6Gpm
4zK/bgQ6AKu3u18AD0plG0HusjZYqGI7XylJXV91oPVFcL5qO4oWYsndsXGn5NsE
l+k8/o4VIAcWgjFaLczawzAWVu21SacgUdYoKJH7Iw9Y6jiE6YtTeWdekNfl9mZT
smAMz1jF+EzpNxAUxd6WW88J4T6GzaFI5W1KoDT/QzSe3DinzwUwPdGGDTn7ZyoJ
4N01U73XOjgPNVXH3TX9akSHMMdtMfmskIKf5rnPZ9HKGcNSikXHVcJZRI9fiOu9
3syOa0CMQ3OCI6t5r9recz9p9QmIaF7/TF1a5+BG7+ambqPyblguleVLEvqMrk9O
XaA4ULlWhycdufYCHvD1CBIQAX02Y1H2rfa3f34AXVmrQAU2BgPh8N6cieb9Fsm5
/JuggPQ7dw0jbWbPKpjf7NpEgZwN/8Uxq8g8/ds4MeaLlX06EtGX017+Q/v2bXAw
iAtqgz5voFFLQ4zURGV3i6nbrtgR7AOhtZHZo8L1NT+KUGV7NRBc+KdEwFYo31oT
o42mPM7ljMth9NPhwF/zzKyqggems2xm2X6J0vBBs9dhTSx5J7y7HtMDfdve6vYy
dwLpi+lvdQt861nFsE+3kCTXu6luLxpMk6OXNTOlmpfExOaZ1vbnhK9IPAByJ1IP
UwFeifxwAWXRANglUaUrBbRFa71cshMr910neTys8ryUKyX4q2aKiShQhs0Whydg
JlpVTS25andZd72sdCIHVQnIzuuvWAt9FIk8BCiTjPElyQgVBQPl6YJdzj0ab0lA
WgjIRNc7iprD6trJhrvNjBTrvdkr6Gn4RxslNdVMMk4O48qYJ3pX0HFsuhfGVrsU
QnDCN/ZizkiCOzh37NZrxmuzuCI1w82RO/YaUsDnNvQmRemOe5zHXSDNgsJ1kreG
/NKRy5FfvZ2OKITU92D5tvSID6468oEQ5XBxKKs+RKo=
`pragma protect end_protected
