// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:40 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DdkDnrB0Lbia3+BKdktB6NvEbxnJnY+VxIV/3M1fuUP6gxdHBLqbOTOOLhN3ke8a
5BXwz0vSxev2ZPsDnpAl3O7cbCt8nSBNL/HhivjxdlqbJjiB+g083ykln121+xf3
k52Lf1eDPipZ1nZXRuOLctMuAWmgzJDVqW+W+vA31z4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18912)
MpHTY/BpG6XWdL19C/EcEbI/rcMI0r7ipwfWqy3jst5vXSyB9G/LoFfuCr+TwMzv
/7JMPTNkGg4RtpMwnW1660tvR3h4qDEcSjof2msRQPpc9W/QjPK8hu1hi6rcRIZ8
aABelVt0KBMnPbJv/pYCkW7enLzhejlrxHSqWAoVzw8cFpzCXrAvE0OnH+Dao4y7
N2WfZxH6jcSxrjTUDvWEDsCGImkr+9m7E/UY6I4UFDHTvtqj4ec7waGzlwu+vWEB
bhr99aBnXht8Ex34Xq8BvUpcfJF5Sp3NqvlHTDGjAsuhrTjAoCS+CCwm/i3aD+Fz
T07EQO/mpA/BPIkC/6L0X1DQLtgcUWDlzh7egSulDBUwXwSRB9F3ociI5SGRI85n
hHSZdLB/pPQKyfqywlXBTANmiba68RGUORdf7vAoz5Yliib18hMRhSJ2quZip1Qh
GepQA9vhXlfYRt0qAnKrfQsDOu+EwgQuSiHX+cEyjAgBFNJBO20b7BFRYQijjE9r
gNS9UXgrNmhOoL43c5SBfluRk0FkJxcYsHXYeSwMvrvS0n7b12BDO8miEARUHXqi
hOETUW42mGQTBF9O/FF4NXGr2jIgI6xXM4bTwBbgpGc2RuiSG/Mo3j1vpAj4c+38
oyXKNNY6Wq3ug/q17Z9Daouk7B6Cpm7clpDqrHgZzMntW3VC7Q74q26SCnpKcSiE
qN0vTRlBsAB5pj6Qr41E1dUfihquEWCiphEsADcwz4P0BSBLx9xEbxfRtF4l+PtR
dLiTU5Oyr71RZ3531bggAzZnlgM7Q4I2nf48v/VjN6c/MbPucj2ich3w69TA4EvW
lYFHzg/0WkKh8FKWxUF1dkw28GcNvKhoaAg3uuRA/frriXidM5dAKFsGrzvAgMKi
9M5jz8ylpUzbyw16Io/lrqMdc0vvcoi4GAyYkH9yp6+eerPnBeEo8yIP1+WyhWxp
lhm6jEF2NTnXaWs5nN/I7ZGnKDe+N4kwFlqMGYz9fu5mC8KwaC6H6ULSDGS0AW5J
Go7ZfK0vseRkN6MjshFFwYf1sKWQ5LStHyj2GJfoOjoxTKMhIGjiQ+d4I41mi80t
i/4M3O2baRKJ2iwgsdyUzMvqtSb02p+OCuX1L8O2T0YAp5DMJC+qdjioj7t4DZRn
ibj76oz0Y54kN+WcFXeGSX3NgnHVhhrUSqhV2vU5w3NRYYHsE1UC1VQKbNR+TYxs
LqreMrd0jF/Q9fMZyOjU8LWcTCUsBvmV4FXZ4QSKetyLO/OHZxed4J9ml+lgzmzO
NZZP/fAIMc1ekqAKY245js0Wh9S7rzZ3WRaLgcs5GmU1kQiobKLX+kALUr8WWWbG
RMNrtOkzKFO46SYq86sV00doP7Y0Ubqw5KrmHgZtAv2HrCqMRCP+EyQXT4hIIJ4t
+vmbdyq5TpK7aUsdZWUpnw91qaRBCAcRDKJGFULJVBNhgvyyN7UzqJzypej31sSi
Fkobzln6s5OSXOUeLHuKS2zHq8yAqoQtHwWy8BYWBZ89RxD6mR5lFFTpXZUMRb15
2ESBhpTlaMC8DsMONDgfAyFs3oh/U67P1uT+ZmrZi4PlVqkxlsWuHNgp7iDBvOND
YUTB52+pTJ4FjQw1m9nXjKHIXuHsutk8G0kDaTYqRtx4qkZUJmRtzIK1buV3yhQk
jMCui9RKaXAxKVfjASEUU8Z3XPbEvUFI7RADBKDUFw8zP/7+nn2eszTjzqLCZtdN
hmUxFXtd2gKlld0ETHddSvFMH8pu31NHo7C/OOgtcwfjEVseohlhSvMwCHRD5z2q
Qw8RaHQOW+neKsQd9Z654hDnYuUlfk1WrQCWPx7EhWUT9at1B/gthiFhzF4ACcSY
GUDRcTW0M7eB4o9HaoN5TY8pJ6cGko+c2E8MGaX9MYLJ5VPN8qCGNhqTvXYdo7s+
IItnmsWCHwWTJBFMbLII/z7S9fUYqxI8kjYA1MhiOnTjjwsd1Y9WiSZ2FW13JGGx
dJEK0Fmuln+S87B1luA0S6jUyJb38XxF+0Dp6/OsGOK1MUk5FqOZznFcr4V8Nfv5
Y859L4h3g6d2YLOzHjZUajJbfhrJQY2C8bPZCQfJc6yWyAZIArYWMksGp81RLPDj
GoaVE8DAuYMkdtnECrPMCzCGPPVJmbX06km6VHrWUud7QbIWPtmluB8cfMf0qEXD
YvM2O2HaFS+FggKKaCVDBTnJWBKcPR6c96r3epr11uV4QQwjACOaL7HEGEgIViDz
DRQ3XK+J+Ga7VpI0i54FRVpDtg083OHvmFr4K5icNaCZOoKKXgFNO1YJlYtGJUw0
5Q3PCTvyeyhe6bAyFkBHSQkZNF7ut/OVkpEc+woFChSHXupFGr0zuYb93jLdRDei
slt3SQg4wLKQfuySP7OtbdeVbjeFejT79rFLhhyFYnSeDJevVB7jVWWKaGHE0HxZ
RnvhdfAAObOYOcISaxAeNIK1Mhuf+k74f2Fub8GqASW6XgbSIXi/2PL4rGx2uSsy
0QUt0Q0OoQrLw1qNnJjYsCDuHjfwXjHJUOj+YQNuTMch0gfbtiiGPvIBPBlMkv0z
YbfF4H3dHp14utAK4CMWjHRbSfLR2NclCQUAhaVDcBg0pkcDTpD0bExzrZ1Vwsrk
scxZTzth+hUwKFsVcSmwnxUv816MlE1lVnm8QGPoVyMNZSgnYiUnpgEUhWMeuz5X
wgEurWZLEBJUkt6uVy02/DC6Vd/E2OnFtClZrJuCiD6jUpsrJWVQ+Vwfrmwa64fG
VoyWLAuPUi392Fsvwxirf/xeuy2oKADUkYbEakAD7Ge3L90lP8kBb7mUPaUkNNQS
bfrWTRWpl+nd+/GKsNoyRM9e+IarS5j3u/RW1e5EFK7LHZyxPAX72aqcRKlh4b/S
I2JOefreJ6EIEQrnSDbrHe+c0Y6Kb3eHTyCej9YREVwclu9RJZJnzoxMT9dxgezp
fxzXk8GwIqKz8H1ZMpe2Ld4GhldsAjj9kb3ZF+L89ka109GdFm3JYccpA4qKiEuq
qImZJKpLZn8XrGmwX9hjvPdYJTttFdz6GGfoPwRhDYvaKhUXc8xIdfFo94iECr7u
j/PxjGftjacKpJJ/rB8aOA1A2RBQEENJhUSkl8Ey1mCFFDYVvQjxUs/DXtHjlg77
Gc3/IqUkIn4svDun8V/jDGA9fU0XoAy8daQh4UonqHwY7/cwhWz13EOV4V56U1Zm
poeViDtIDo8S3FPLwNH9gWoG1NQnCfTH4F5l61Y5x+j7bQ+4oidj1IL7ACfohff3
fq4EsSYuMLe0p/8AjuxwPSTnloMhySa3GVMnOr1CvZ3C6dfaPHX1lcfUo8aw9VSn
iw7KTvz58SEqTuFd2oLV3bQkNqaCs69+ksC2MOAyDIvWQM+A5xP8yYULD+GK4BD+
Ty9qapo3VHiXtT9C5fSTh3cN9RDunIYpy79eorIIX29JaiXDZP9FjvtN4O9QmG79
QYTj911U5AmN3HefqHe8PZibLZ2NN7Kx7qsqi0SGW4CnXRNBngGWswvZu0PEWQQT
y27gMvHoma4JqPsHjhdfmUi5mhdBR6ZIgKt25x/D4JKm6rlmHX4NDsc+VUyCxWya
7PN4+B4Cp/Efgw3q7ZcT26n158GjbG4VUmLcmXtvv7c7V8RuH7733Y2aIVjM4Hid
Xzp5pvxaYOfUWkTYTnHP1KGNZtHPZe8xvw7RrX2tYWpWXYvyxMUmil7rzEmbpEmG
h9q4DLxLAe8b7QU54SUqtna7JpRsdmQKzO6/+H5dmMT4JxwsfiWirKHbyHsYONuo
Phu58QMuGWwknsHTH+wFP7l1KOTDKrvqfuXX2n4JXDotNz04T9NmmLgRL6k4pykA
nws5jNRi7+ql+QkkcY3Mbp7+7KfX6dBbxCe9l7M1QP6SOsWayQfweVEkz8vmnIRw
7y7/kYorScZ/YY4TZLxbSU2G2TeSpn54dIe/ilnkCYoK8dGwIHEjTFanqZa0WxQZ
99Vdtkl+JfsL1zZ4EsNctTC7KI3VGOvWUZ2uoOw3MmOz3K4l+oRhpju68aP8Dpgc
YhUg9DkUuNdNmTtqRMCw5OTxmAN4CbB4Z3BRgt9zvWIZPG7JaZ465KmzIQ7u7+Pd
S89CEsP+c7CWpJnwX8ChItbQHCxgnGsJUYTGeLxBGKdbf5Je+ZSz1u+FUU/c6wy+
/gcQRvq7btn5BWe10+XK4IaAE73Ka96ya/iY0lkACGRfflQqxE3wMLHFWLnyskTQ
ypJyAz+U/UrgKE7kMsWgUbvEVI8Q/dEE1j1Rx8lqlZ26c9E1ZVGJP715tdkE/BsX
VpJ04ry32OLvrRIRNinO+/Yv2VMDysjlwCvHOPpRQuOexM42sWNdN+AnROPuV4yG
3tLRWOvWTSrevJVj+gaQOvzDLmoJlB8yMaRt7ODwYh8AqxyTZb6CxJWQGLIj5ikD
EHYtMiznFcI8NpnD0vWPsVXD9ut9xA34PTXJgiBDM6hcYX7UENAm5Vng5VigMC6G
phjo/nU8rooq6HX9RgiUtWFwvTcF+cBAe0/li/b25QONir6ZSpIca2XLscO1V6ME
R69TplIpgM7PxIqoiw+UETXjq4booZijqUoSHq5dSMkcEsynQEAz/2C/zOkMbfRh
1z7zqJZrnol7+p0PQJsBzblmAHtMN+LdpQ0+7gbwPrXcwiODEPi7Dc+iY5hqx5BP
zn3CwlS0Vg7rrWi3Qk904BLhm2wSXoh8kyMYZXu+1zIPwVnfvCsMXIEnEaC1SM2v
IH1Oh1H0H3Zzvdx89b5o8YBpscITco5n8qy4JsaZHqL/DIl91wX9j42oQDrIBkE3
5k2MpODp86QpZi5B4RtPYjkkCE+GKcV41a7RNXaIoSnB5imGDtWl4V9RTyLgVTVp
EWyFDRBlSCfaQMY/W97SND42KUIvzpc3QjliSjLxZmRwiyQoDZ1bOdU8sgGGMpMR
hQHq032j+N9NR8VZhvAKHK4aJkB5v7AXqS/vYhmje4KHgAonpXQ1hQTqZUsNUykS
kWGWs7TN0QId9uhyskIVI7uxNaum0O/Ebm7gMB7y9l2KorraYNs0FeoAsl1tr4hL
rMglyYUiznpr+y7F47qJok514wlHj7uVBwcS82yw68/XFYBDN1dVIwz73LH6tmF+
orTMHMxiSNfznlBQrKwbSMIFHmmFlWiwC19CgcDlzffSOtyuouQfEt94nmcESLE/
R6P5UpfWHFwshMwDN46iu4RpK/Y0fhTOi67q/zWrEZQhUwIKR4P1iNuprkIZ3g2o
D8RLEFadKgPyc+XVXFUT0bieWLVwwV2la/sJZ6vtsTKubssumaEtJFc6OhyIGvIA
Fq1K8YKBEQx80o1BvowuTtdE/76v6apXB/IDi3Zieyl0r8cm05swZpWrI3daoLpr
Gw5D04zDE34i3hEtksYTHPUgS0uYZeAgngKXjdeDekrkrPxZtBzv7zRG3pnHFM9B
+Z5fgpLZJSq+2T6YQzMSSHARKRLva+h2TITTntBHIvw5ZiUF76Bk9B7BGuykPhdE
FbfqM0l+AMw6MsjqMnGjtvc01lacT50fUi0fdI/+nyEQmvExTlohLtTD0uJNB5ru
4MCQS0D6CzWfuXtiytij+J3KjsdCgXc6e84mNyTDZ5hl0E8Ebtp0uimhSoDlacP7
VYAGGWsENEIvIBSkjwUnyPLzOaoPwaTYeG09ujb06vVY70E57+Ue5+S228NK5ge2
Ov0HJPwE7ZLrFT6xh+YRRabjR3wRL4AGb/rWuArIbTC169JKvgZBNZEFnsrYtZeZ
8nHYe0wdZ4D4WS0R9oJFQfJviStn9vv9jgJAV8pD/TNq5/X8bsSARYF1JOJ4nSeu
1PemWeDwhIE/4sGNK4mwfQn9MmnS0RMMraTnU7uwdXFAa5oKy7zg7QkoqArofckU
V0RDFPqlFhz7cDAU3UVrNA3NkT37+aYOZlFNzLGgJboKU9bBzd4PHHmqYKyjl7f4
HHe04oOZcEr7MuFAeBlFqv4xTU0jKClkwtZ7GR4b907ivXU7xZpPahEt706bG7Ua
cLklIxhlWYKBkXtAVkDxsuqMNAgR7eK4Rtw4ekfd7gnEHUL1/kJ3CCDdUDy6dXvC
ORWgPzY0iaXmibCAca7FtREws02l6wxufDW+pRLauJJlFOuU+Ix0WDYPxg8idbBZ
G5MBkKWCxPsi8rN1DBjoUrFWa2+ckCGCh6bvuOXiVjaiQF09cgjfhHqKTJxXXHGX
il3DkG13BuzQo6EaHmQh1jDrygwZgVfs60Rd4DBGlru9JM5xU4JuUZefa6vnjPnv
IVIdNmb3TPsnPlB/Hry++7bBybdm3x+iBd21YJkkrNG0hnBIjClWZSwDgCXUTecc
qrhY9mRLFXMCvgAZHUg7rPZcfC2mg/5m7h6XYNYgRi6tHbFge0ErvuDNa8rIi6Cd
CCVfZ60vQ/sksTmRo/jrCX9wlkrKQoUJ1JMNfZT1HdBgfdN7zy2BarCSC8xEToWo
j2M7nmrIX5NtelqNBi863XNxfLaj3EWexQLu0ZOzz59nuZkop3H0t26EanqulY+1
sV5iau1qPXRbedR61M0Uh0KPqkT7chxKbFEK47i5uRf3cyldr2stxeBqv5P0LYZj
ocZXbdKlKZoNQUg3rC57uuF/mt7g5xwX11dwcGtDvhdlz9EcKOeP/F7lVik7E8zU
T6L7hGb9MQ0vf4XtBTIrxAvBUo2w1Lf+6524PHfONXjixD0W9lgyRfyGemH+gaH/
dfDH1BSlNujzGo9aZD7j0zmuC6ctX0YFhTR251BeNARxYPhY3Q6Z4GENKaXHMs/n
OAbjHKHkStLsE7Y1MJbHgg1DAZDr47SJa1Q9vrGmVLPqmpRBiTpdhbU4i9LD1l4w
dUa8mVrb5tfpghMlaeSJQxP5KOLmqkMRsTjLyjD2mzbJyfGpr4LujDRyzBoY+I2b
orp1BA3DgWkTW5ieYdqojVii/fSjBYAoNnojxZT35wLwKy8ft4Bh3Rd75g9fJvLC
JQPFOlDYOwvdywP+/xumgPWqDxXCsn6p95HVRcdhuBrZAg1RFKsNW/r5M/YcMRAt
iysVQqW8gaMUNt1sFcrtsk8NU/FEKXsVIj+ajTNBMRY2o0LTXi1goE8+oyo2UPOu
LWcsDfTAKrhSBrosjaKW9kndpmg4Et+HcpHh5RiPat0uiy+w4mfRHd8OTaZUXyaA
91CDCZdoqdHGFGyYDa+o9yX/lgbBBeulk+SrwNui4L2wiqC14EMWsNNs5RP2NhBx
t09G6EOGgWlIrIFcD7LFak1LrxgxcHvReeDMaI2WDt6r7vrdkdxl3zFLYjkQP657
ae0JlLXcDWVHPGbpTewbetHldMmFMXTTaoNrpN/Bpjlbe7fGYyELBxGILgZuDEJE
k0jFF3ns7c2wNH6ZSypcYB1akewJcAdMTofXnFjmEZNyg2EkIiETYRTH2Fv+onaF
/U38T4bQCCtjutx5yjsNEUOXEFRn1tTWuD0PmEmng+YnSBGVVWKDtAZXeGbX5Ee7
zO72DA0ktR8SUGxersIQSCksDX1dE50TYOdieopMsiXvHXO2QIR09+Eh28rdW4fR
Ovu8/7ezDRRK8gTnDJzl4J7QUe5OPoB+xcpV8QuyfgQkbH32nq3PeMzs7eDbv4p6
vRZhwcUwog/QqNAZPhfgf1N8tO0s9yKqz10f+Htuz824WgWTNmHzbGhbUUI7YeTl
JvwjFDkrTPTcZdo7gdddjnxn9RLum7EHBvx7MpFijGhG8iOoaO+wUqeKEotc1JkF
R29pKc18fQoFK6qyeeLs6dnLsVOBfdvfjj32F5RQCpbGE9HU3IwKSsryu7FTU9/l
YisUb2VoV02L2b9sxMWMEJ2FNmf86ZqlCBdzCX5vvBFg4m6IRAIlEeO54XAqUKSf
s5PM898Xa9vx7TaRU+JJAP08xeetJoWeu8AH8ZwSFG8rW7nVUoZTGvbeAmrRoQ9W
iUwM1n4FbcD0HMdQnl6jjk4nwyJTJSGEjDk0iVwKDH9KpiDEJRFr4PbiX97BxikC
xX5R7LcVdokuWCIIcj93+Hcu2W9pbGmeZGHmgyXWQGqsaNPptBRN0IPS9hEbkAku
WZZJEX/UTk/STLZkQzQTx6S6ZgnapAgD9keY+3Xr9g42Cx8I7IWDfD5C66E7RVt3
ZvMPDgVakrfRxGYhZU6xv5B53Z+PTClkmBl3xxhfLxVI7q7cIGO8ps//s9fe4rwW
QmW7MYG0JL+Ljb5MD/d5HPBzvH6M9l/u6nzrbbcxNV9nuDs3boBRvv9vGfNVVhiO
zF3x/QMtWgMgUrj0jGR7FDFiKbFTVzM1ZA6lmoWMDdnNE+rzfRBcGjv9s5njQdSO
kN2CcFt98m6QT+Y5OVqEPe7Xiz9gg4/vfdHfYtYIy7FdbDCFiBmxZDOb/+ktz7ls
wlQCqSZz+iHNrlfBQlh1aGL+nZVWVUEyBiKzYyQDhBQz9jovmpIknGPgutVTI7TB
kIZbePUn8UWmjdRr6Bs8j/FHKhWRGTWWIlb4Yu+NCwn5ZguhxGSCjQnf45lu+15J
CSvVUVvTbLNNnl2t4FCXiDtr3OkdxbZwjfnkr72MQ3nSCnbVb9cBxGhq9UOH8Sgm
GWd4K228SfdDSpt9itnxkdeyIDG4z1/jJu2RQp/Y/LOBxdkFP8+9Fs96TBVvwEE1
OAx/X7tVy0tS2zDbFyVmta00WBrpYTk6L+MMC5wkQSwpEpy96xpELxAF3yFDc8st
NHmP5zZtIjSMS8iPi8wMyztFbwZbZY/hihCF5GYDL4KwM+iYN/QB/SafzCf0FtyZ
82VGzVFeI//yXdpePV2sif+O2zPX1+TURfjeA1qEszL5HGTHyWco2owKA9Zryyve
ult/abokdWLcfadmo8VYOsfh4ycdq9+pYSi/IpteT7jYUoeOoEesK/YLAPzGXHz5
LPR0mp79MwObM3xecccaXfqiKlOj3N0mJ4S24CFFSJC+pdrn59nDvC9WF8Cuyi0e
avoSEAdu+AyRoxc9viMlzd9H5UWiDoq0t4uYTa63CJsizz2UxYQeWz5NwAf4591Z
q9YvOzYAJl0JsTVuXacAgUQCQiLOr0AjDV+ekeD7tuFratkMCQAZeprbwzkG8tR0
tb+znXAJso7W4agZZAu5DoBmliopTqdYM8/72a/0oIOZNb3Iqr+LeiRSeFim+lT9
TbW6ur30MClvSQFpdafFG5M8+k9kqx+nR1YorygmJhY1Qtot3tTZ5U9BkwnYvcub
kUFSQEAbrdgwXQiTbAq+TT+bl0M6E05DGjorx85Am4uz2XdCKWqFiU6RfMEWmgPu
eSqlGbk/eODX+7BSZVGS/fuWazNua3qR99KJf2epOD6EbwwU9LKFd3pbsPVPo7ei
FhmWMngziVrq92BvlC6F/sxxsfrBuyTSfPR0DoMKpCRdKrWdBBzMrsKhaiM0lwqi
2iOhrPefH04HZYFpGjMfmO67KN732wMrsInU5mtchAINgBARPpLHClLz82XJIVku
Uz5RS0QIsSu/rCf/Qoqr/WPJvqTC6uoFSjdm+LOTaVSJa/7N9fBRwInNYhkgsgVq
CXhB//MidwOojbbrQFxcxdmN+So5cKWZxAkZ38gBGTGrRI72cnoz17P0LH88mcMc
i9rzVbP+0rl1ooRttkjYec1YQe0UcvoxaL/7j1LtYOxJ3Mbrz7OBkZfC7dTTi+7y
so0Vs9uuxTO2QPHqFXKiS2UnfFw3rauQHTcsbICSN0UOzyh/ptpM2RcKrW/9THEs
aKLbSv0Seq6Fj0z0R7R7bownEADT8wCVzy1GaSn9JkD3vQPPeCbgVPOd0fX2EcA+
VvgKFg+6rM77kOnHQv3drpBCSwMlIeYiJxROhjRF65wPPJqtdUC0DHVpViCHTP0Q
XeI5DKGcWqhpzDP2DlGO8zdT7D8sIkbz9uZvTuIKbVzjjQAfJb3TwlCDjNN9uBBh
D1BnYhzvQyDMloz2CgLeOo7I4dqv30cJxEQNp3fCW1/E/StWvgsXCQrlf088M9h4
HjXNops5FjlDXLN6hHykGWeEEcuQD/JCkqURpaaf4/VTZG9fIlIwq10gRDWUxILQ
GW1HmcwWhwpL8Of/ICzlqO+24n9ObEPhej1WBJICPcwU4FCMFEo0giDVIruGViKp
4qYVfxVZfs8x53x+mA49M90ntxYPPNhqY/b5GlCgeHgYDrrUEn1FHqPpJNmD0dPH
l1jOcXH9Y8JaZd0MRO0EmBZhlW29g7tYKMY/YKWBzvjsEC1SCJfK/Z7RASvx6C+5
OqktWFU9PFnnFkReRnXXjrxKokxmspFsMO2uP624tykt+tPcAG1aa4Qqgt9RAMX8
wDSxd2/6CzKbaIr6+GhMEVhctW/4s41w/e8B/QUbYLX+wFBA0qYru/gBGwDzrHad
d7Y2plCFdVpcFhKQO9ykxp/DOJNgrzRA35JeXB/7VuRYfpNhaKLRyLU7UGHRDTLE
vTubFlZ0n8p4bm1kZVLY8jBulk8mIjrNGE5WE9QE66wGJPX68/T2mnYoQRUIBB1L
Dh1heemr7WcVAzK5PEHLNBi8vWMS4nwhWSBsedy2hU2lOLLMSNLBIYQywZvG2Lhj
zY75xOLkpwTdZ4UkMgILprr2zOn//TDaWgW1aToHOlRVS7cmYO74a3liAIS3o0Qn
CSQnts4XX5HbB12JGQpBZQum6OQ+D4fz62IhcNbHRIhCv0iYdZEn1eVhGEREG7hY
DfmrkQtV68LobSP0pR6Gia3BlbU3D/il5bElcqchSgND8UXDHJeK5bL5TYycDHpT
X2Ifabz5e+J9JxYgk+tED3T8gBzeKBSQUNn5kBC6622FFmdY0NKcsGzGoxr5z++4
ge4PrC5KGHBJZDYLYz8ARyvh/uNGhY4Z+82l+zz8CoVEQIoKzsdJA0GEgznj/9cM
S9ttgHGZmaLo4iLL9JKAt+nKhGo/U3sL66nCP2OkVRFlxvTH8QoVFqOGf2VuwkR1
ZtEdGUKgEULyJfW0lhKVNKmiA7XcIktlkxYcZrb257ON2R6YCLYMtc52ReudMCJQ
vd3Q/vjRTzhuGmohRfgwIqzNRT2VzLYs0POGWQ1h91EzC/hMZWNcM4fH6v1eTwXj
YS/IG3S9/6YyMqcDEqXub9IlSw/hbS/wuY5Ehd3sXhdAz+6UWZpISQ27Cek0aikG
6w9xyY97WBAqTDl9tFft0JMEusQZDW1SS8633K/z67aPoBfBH5C5P1iwnwiYSlDC
7SMwMkS0ZCgQrMKVzqSKxiXcAV4phMd6yot6AXZ2gWOK/6l0c/MAyiXbyL4Jmfce
j4R9NrQ44QMa5iBPOg1RkbZ6STbyuMKO4Wlcw3FbyZTCFmH3PXmJLRdM5iblq2Lu
4Gm2yqEPh/LjedjrQoJEa/bqVaLUb4Ynb2x1aXdaiVvmAsS7AUS3He35cNad/kbM
vU0eCUZJaherAm17PFd3x7Qvbal7FhrXSQXI8KRvk9M4U9axJdbVRi4Fzi790lNn
o7WaOQfLk4pNMQeMJLFK9qoQYvMXy9w708A6sLkalQts2SI3htJqGscB9E+Jbezq
cOXitN7hEpzFILVu0fwp7Z69NYHs4Bd+42R5JgWpUw5zilPYTmPWQYy3x3vS7tMf
V+OzJU/QkTVZ9pczC55JofcY6VoSG9C02fId2/AA1EdlqLsa0mbvGaUyDddfaXAQ
ZhlII9TxlfYNnKTEs09xHhBGRpktVUyDTSFEyC2wRN73wpAv5iUI6T8z/pE+5Le9
aa7dtgnEkh1nhHCxVQdT0tN9TrZfuMjt3hpfEZ4QCrheXipdXuTuKd6Q/ZQKYPSz
ef1oiPqoS8OUMOuNbnsb2/BWoI0JIxt8vm4Y3cz9isfCBSa9h0T+y7fBf+PsMZ19
NvMwZYOEW6pLwXf9Ltc+sYNvSqBT3mYhlmYdvQxE1dZyLCgCkAeKUZT4iLk8V7el
/E0Gi70kjPzVuF4uCyDsLoL/1NMjTWmPKsXG9cCEq+OckkWyLyb/8/+D8Z7tgjj0
a6QUpLrYFUjC2wY3mAb1eVTHS7WEC8MI4AoHDoJatdeH7TiHWs4/Pib8JdFnqMDk
uj1BJBV3Df+lpXO2rcnovMVo2VcK/CcPZTgj8Q5HG9GO3zPmhbdzAi2X0RWMB97Q
F5s5cBObGQNzJPo3ST7SjELqs2HJl0Dhoc25DAJuylOhxVts1dRsLxn61SOUT46D
6MSl3E+7wvfiaDGxLWfJjFI7RHtkx7Sdpuowogp2pI0aLvup09YfxmUPKSoG8SsH
IX/4xxg+O264NKRmFu+oYnH+m4OK4hCOkjkpreo2Fg2SYaI1rmybDcBAo/5EcD5W
g/6NZPC6felBpNdZb2ffMJf34Q602PyJ4bsM4nPULMeb3brPVEjAxiY50ysn6eDi
qCoSdjzLihkhs0liMvy2IdF8jxP3JjFCFkZGJ0os+/bDLpLd3O9lGrR8oAQQhEVk
LdYj1/2F3bw7+0IjRgiYqdgZQTRh0JDk80+K3wyg5wUbYueUxuCScSWpXuYkv2SY
E2484+uhx51Vo0Ol31Uq4fjy36QvS/i/r8a6ei0A2s/t58oxLI6HBqrSvD9GPoaJ
cAKDg9JNBqvmaS/mB3bm0eyPqASK7mCUwHOIZPExxoC5rE6fTTvo7gMOGyqipOLI
qmQkFuzG8pt7yyFDrBb9x0hu+awUYW1sM3aTJW6d80ldDT4iEDkbB9/KvfejAfYT
9R2Q6/W5l38lU/dL/T55s2xJveNDZLnc3cYIo7h1LSGVtf8UacaOQqZIoC6dIK87
AAXCS2NVA1XWtBqrUCswxuEjaIShxxxYaAuxhSd3qFiVSF1DdDk5Bzg7Rsb3+60J
XgfTjgxJnkTZ7zth4MlW9Pe6xjxK4SWxbMsmNdxiMU5WDvP31GgDJ7qycvet4+rm
6nTvMgi/H3VqqD2hsJu3tSvtTO3pT2Zwdt1gNjKIQAT8YANnjju7Al7HEKTHIKUO
425a/sJYqvKVGVMyw/oAgCbvaDz7b0hBB14ocpuoFPgqHW7ZLqVHkYzPiB09BEM4
+2L42W1M6U41G2SkYmdTsKxVyJqKSXlOCjKFSDOBQqMBrMdBYwvbfsSM7lDR5rWj
HWWgIDX+zlgXvTA/4Agl+XfI8pchGyL4ypIU+aCKu+2NiI8NmZkjDx9FK6+X5unL
r6JuR2OFhuV7Xw6Qx0HA3WvtvC2LP+RofFyqBx4pV8TY8hortdtPXvIdJQ9rPlYo
8NtOhnw0dNdeOYfBHhnmDKhPMYoIXtNeZj4OyWqwq2Jzk/MclWFm9ZrD7fcc1lYr
ItsFM5T9r2prdXLJSBGi9Nf7+MI7P7cqnNrHpYlxYendM3Q/dupGxdq+7VV88DaA
7qcDTbWlYMPH00neG/OyK5Hni65LSwAsF8TcLZ6wTiWOX/eRCN7ZUMhcFEj4jkLq
5PitNMhYirlJwKFCMTQybQEiAJzoO1N0OGa46Sdv1J4z3l7VPm7aEWWsI9MwSxsI
/w2I9UL4u9ioI3UuXcYitw3ancX05L0Q2kwjlX3SE8Z8RopfTDN7GKKYEsp+Ak8V
tOQKPK/NbxcY8tUlkL6Rfhatpo3w95P1ncxMOKhP/iMU7wYgRaFF65gwVI6pA/v8
TNLzG2OTAn57uh/n8uedSo0tetEh1licVouwYA8TJtmeFl6kfSpwc0bw8/zRiHYK
cDG70YkWVAq8Eo+ZGHtce7MK4yZ3vpExW3lxT+dEPUR82oeeBl9M0U4pO0CPJJWH
6oHY3dZ9/fCSILjynZtRf0cjEZak5FhhLgryVW0WXZcPDImgq8TDEaV+wuXiaqRM
dSCEuvMZNKARMUBrnO+IlFdjoJvCI4i5U/46Z2fr18aMUiIjKazkkEvghTWveQ8+
jSDP9O0rH1S6EVBYVEEVinLB86LLfsbpVOrrqLtAVr+AUUkIGO3BshFYbMZAGn1R
eHgFmNaaK3tjRwncUJdo1LczfX70GB77rhKMylxdxkK8ThcGdGYQmi3g6+iRY0pl
eAKp5PzpR5gKngaZJdSkkPIW3oP9/D97vQdSuMFnNSb/NPS62iRqPVfcxCjY84ks
73uTEYb4m6g3toAvzlCdnoQf33MBDrr8RYyIMk+YXWG8D6ovKuPQYEqV661bqbk8
ltWp5QKpZNJJbXoszI64CJLUQ8Lth5GKs3qlODJjMKDsW5E33HaAGd4UAyIyJexm
pXt9rRpGiKirwZt8hF7GtHzGcsVICs7qny4ELoR3tlpUf2G0oimKUWmNr2vMpEYa
v1Rr3TE54pQHmxdEHl2ovII7bCbJ1xJf7JG791p37FxwLzAlamfAomfcr2NGW9QE
bobH5B9U1/1+AsSFwR0RWk5XY6sxv+6ua+GNJhMMwtkhUI1xkhM/7bL/ef3LreNi
tTk93GTZ9X9OVvwhiTN9lcH+KzEthMeJDRHURiqKelP4ivasKUfHkovNSD/zKcRR
1pQ5yQ2XewLRpWtpVGHLFxMhTlEfrDAnnrfdQ4leOMa8AS2/aYW7A/eCHhP1MF9B
dlPsiLuxpJpNrH+Dafs4Z4ylTQmYquJFv/Viej3a178e7vP+EJ2X6flInrLRRj5A
PiWGvneVDdqK/W5d27alvbDJuVabNyGoWYGx6ULVmjXzxTwtoY/rbvuJZA1L5lBk
Oos58V08IPltIW7R9zAEw3R76RqvmoH1ondhYLOSWCDsy8LxzZmmFUNLGh6mwg02
vsxXO3ixRHaAoHeJQ/H/AsoushB0ptxacU15h0s+jq/+WEkRjSaaC7JlbAFPQKh2
bKjWn4LEkh2sCUrT+GBP9ahS/YjBDBJPyoALXlADXGFfZOV/TPmu4CVDts8ZVb+u
lTBc02rHXL1HzkEcsNLla4/Gy/Ew+KB0jcTFX+GSO/AN+ak2AKykERzjTwVULc0R
h4TVroh2W1lvG5B+g5m2Tt+93KRSoVzezhcAMxjvNZK8ucWy3CY6v1OKlVxA3X8n
Ah/PsiQfdplELJMh1DRSXuc9Lj+lHWZwp9m3oY26FovLF1GO4Gy19zuDyNTCUyWF
zDxy7g5e5Vq7nbHJ2YwwiznZXImrNbCqyFyP98+xvQO8NRYqKPM1WUPb+6/37GLJ
6BJGiUj1xvGg2mp9VHjrZz/azPZWaoYDVnpgWLZKsEhYezetwy9rwsROGHAW9Vna
kEyTF5Wb8a7MHrIUUgIxVdP1AXh7IKvgaVivQe5heHxooa03h90+s2RsMhvVNwdk
rhhCrWsYz9rwekbiy/AeVXOXAMNEPWeelSIqk8qYGEJpQ4MupgbHsVXBrjec+frx
DxYqzoK0VdBPcvSDZdvyJ+dfOtgnB9lanaON2QEpGoh/AFqdQsm5M41Dn3LvaqRJ
eGZgBouQGNTuWZyCEL05tY9eVeYK9UCnprIWY9F1CWOOfHIROARR5QiFpFXLh3nL
Ml+URziURcEl7AY2blz/+p8KSG9bI3TQdhNaYzlPrrtXxtOdV4JiX/z5g2Qomlb9
Z+sS3FfLpiGsB3nFmrWBTHIQaBwEmsNiivkSKywDZgg1krWKJXNAlAkKUcNKCHs3
wM022vAlcFOReuWfKfk04LOl8jFYTrreiC8KMH2esSlASzMV8tq7dkxi8XnYQ3S+
m+UOpfXhmYVMMM47otRQo83Nbg1iZjNIhv82v2lcv4Czh517OHs1mELAtjOnUTe6
mK/IfVCWhq5Er+nyNOo4IauvXEQdx3bL77UhUTO5K9wZQpECGQq2ukTWqVe6l+Ny
Ld0Wk25tOZ4t07Mqq9tI82NBQa7sAc33BML/+fvpO+QgtRvq4Tz3DH94mScrP55m
ACQIBwvrjfK9L4BvLfAsqOAeAlRoCaoqMjbW+N4HtVcEVo5Dq0dzPbXw5wLYP6zO
EBDSt3ZWcIcN3bbFXDVwk/7eR1Rs9qh8ZygqW3FB0GCTlS6SNrMFKtLjDztO3n0K
Hdw8/Cy4JgXkX9fM1gy38Bk3uISFT9Pux6EFJhYb9w4rs5C2+GN2I/xaqAwNORV9
UxZjXWhihPuSgZeKm8QDZp/gxja5z0cWOa5NG44Eomf1MF8IWZJIqpexVZnmhU3K
dy5t0fnNzyRQzWHxNh9xYYiMda5mPhI+Xoskl1tSTjIFA9nctBzHYLrvfvO5a0qI
JokRI/hhUHMfymgCm+o1Wf2BUeMhziV6MhMwlUQwgNeE5zuMW6ixQSSDciLVQVL6
nAZ5lUSbFbQqY/Md+ORD6wHVCU0h2DJsGH5tbC4fsWIvUQEFLZuSc5h8ARQMnHu2
vAMQclivn7JKoyc/OyVCgsJeLSDYJ674lytGM70wRw002fLG5GyDzE3iHxcgKZD6
cL+yEeql8T3koo/8jM+XeKtS9NSjyQrZD9AjU9aOd6Dnf0L4+ycGbIKkH2KlQktU
HtE9q96gPtoUsTvhXh6UkLUq+rNXMTYn/MlSO4lYOtou4e5Qbkz3njYPqcueu06T
3I0Bx0N5zKiI0yfU6zyh4yewr+ZR2t9Fqxr8H3GuLQ/SMvIUofW3DZz0hN0uf2Be
R9PlDS6SfLbA7mAuBnetuU+QQD12FGHJ8UjCwpqz9xpugY8X+zPWoGRBCAHDCWbq
Szr5+Jwf12nnBHsH7W7Uu3kImQ7o+NOFcCI2v1NaBnA+egI7eZlNEnGY87w5F8z0
a26bBo8cDTvU96OS2JpdnuL/bc0+rBMGpj9BCSidyQL2bpU5ZZy286BQh85T/kc2
AZlTyteWSBkYDyEAKZgDHzICzZSf9B/OOx4EXdqler5UrRvj/m4YRIZkkcrJOhha
WCqKCyhqzOPtuUkjM4pC6sGfTZ0vzNWExkPqBBjHnzDN8PztqZAyErP4Qwl5Xn+s
N+VNKYJ+7um1gwQ3yM6X+fFkHAsKqPAqwpv63rqmTUIJuSCXnvN4V4xumWYTXBi/
VTsGmhiFpjScDCrgRJyXJmuYUnD2gvgMrGQacHc6vMAOX7F8DOqw3qzbXUQCZp3Y
fpEOgS9NUbV6g4UU7OVFR799UAQuM+MCEX7xcWl9L6Mv7H17GF1FJhMddVEP/++G
+fOrLMDxvRqmIom9V3DSh2NcCLSJ43dW2RpwHUiEnoxaDXNny0Ch/Ntrp1F2MuWy
iG4N6PN5bxu3VPnLeaBx8Wy8PkqbdW5CbiAIVVDOPPmdDKgeUiKw8oUTgINEkAaP
U1CTN/eHEa9dL3m+bMNxfNZtHhIqmgAN8vV+SBmQvjBkrVccjwKOU5kteEgYenQN
hgalkTamW5d9yDkL2/nH5Eoxc7aRneYhDpI/J/rsT3ZgcKS2F7VZF80i0YF2YLoh
u0U6iEaJOZbxIFRuLYbPVJguG6xRCJTUaip5cVAQssn8ZW2epDfzZ9SaSzeRFbdI
vuBhbcH4FbPwbg78pMkb2Hb2QNkanlyqQct3jVJi7nM1DAF8DBzF7S8kM1athDzn
ZmQMNqWV4yy8qWHpoeM1Z4VKMePkQqS9AQQMfvyEgyH1TNGKA0HPSPNd/xwTTRML
GherX9ZRcCpDVdfzMNPX00/rh8J+rIBDNMLH9TjdS6QBQJ2ulxGiZ+SjqjWIsqsw
uodhuDqZg6evdIUL+RLK6yfyByUf8IhgCjYUdKhlaydrRq1sZF/ArxmvtgtpNO83
/5pasHtJxWW+N2gH2hCYanjK14TKoJNOnPqDrWMp0J8q4wOEdf9na+0U8lLXUXEN
PjBHPF2qHbC0z52VAS+TRdotQQu4eZVHEvRBqDt54Xg2fLL09sAexjgWITUkvYk+
WCLh12nSaabeYB/swLrNeAVLvSp4b5UrsfUF2q4B9ClRWdp6owbEJSOicD6TE2M8
InDonSJfsP76XfO5CS+8+GUoJWAnb246G8oqMGZq8/1JEYCKqvvgXiOofs9T1G+5
iM7IBtIzf6mHRECm0rW9iao8+FWrqg6JaXcVCRdkoZ/NXi+L08LA5eU+oj8pkKDf
4n38hMyS6bYiAomtwyaX1e62mGgPND4nrePx5RBw26yfCt+qpLuoIojlpvzI0s55
+qldIGwehVvliPLCOe+3UgpGWHnF7uC2DCLnipQdbjZQflmCjArit7gtirqAIzvk
UMarL8mph1j205EQ8wIbY4USDQfyIXy6Zx8dicEfEs05lY00BMKwZ1EIpdI+UTUp
K8Mz/jdv2LQm5ozv9tJJw5Gwrzs8IYQ6Y/RgIXJa0tJiR/wtBnwu2/o5ctOCYf+7
ZabRA3br5TKDJIINjKZgLTK/rxUviYduvRgu1qlfuCJH9ZLa/UygzGMWedBTGgHZ
Rj2tgDq73Hd2BHrj0aBMsAtPK//Cotu0RSTxqml0bxe79cHTIgs9Yd0SmW96Caiv
99iPUyDhr5BSTW7qEO99t/uAnAR0Mobm2q6tVhu9EXe7gMvgZ519J8bnGzd3/DCa
H2BnrxmYHH4JzjPw7EwRuWxHhsTZu+d48hUf878q1SE77T0Z5rt4GF7obrXAyUNu
ijBVadhQ4eVBUHRGkKNe6FXyy1C1tTGVg8UaES7UTFU4U2E7D6YyzQ4uf9Ym5rhw
XZa4UPsSmr4Bff7etVRTqPKEx64ZF4XNcUiN1hjv6HlXNEwj6AKBdYcDm4KhblBx
dLucmABB20EEQKzX4mTlBuvw7EXG1WqHa6KpHWcCuFV/GGNCEEoojBuKgDIB6b/2
Y4WFclf9QUkV/k9q2OiMlgd/wdduwUoEnT434OeTEer6AWj0ZmBEZTqgSKBSnzBW
IdM6ZLGTTlagdtNfOX1D9mm2dBPO4/LVbQ3zLtfkmLGksN2ThOEi8wbTtM5c8LnH
vwpnmq66bslTFrus5V+VoWg5VfgDNOnKzdp48ieNjAl8GszINyuMOKhdu+pSSPJ4
RByKRVcyF37ysLV+cQZ2pI13cd4KUuVcAUvs15sodhIsgxJ9HvZR53qiNpaHBVTr
oCzhTciAp99ny9VhairXLTqVJNKRGlOMD76URNI0CTUoqzlGIqW0RLf5rHQXr/NX
fpWW7WUX4CryosmCzutcr+kH8e6zpNIWJ4FgF+bT5GVeG0D2Oak2OFCgm7XY6F7k
J5fp4STGfGn5Pa6MO8mARhWPGagSlnRHS2A+tJ3+/2aZfuoxSqWK9Hl1QhTTDCOV
0UzNDG2pRWji0VfY1efj2+AecsaMdMlkjCN+OQjNf4GaTrm5Wp70GeWanJ/Pd/I5
FUCtbL0IXDNMQVaMxj6NKiZ5wAqjmDJ2WTPJmSF9XX2xFwH3DkOHHSRpQLyN2TfQ
ANDZe5Hbe7G9TJeIlm8aXkEH2kkB+D3QugYoMGKsuyK/phcQtA77XnoEVyowWUWD
vDs6MjAz5VcNi3KLPr0NQUMTnW+y+w7XGc38B4a+lj5fF4TF9/JiNmkq03ElR0r4
Bu0MfFgL7/Qh+uz+AedYvhUNBkLW18MhH5cMbtuhzWTrbrkVl4EjW/dX80RPgZA7
/accbUU5jtOzMr7l13ecAqwIoDO+VTQG0UrU5O/a7dfUDTVVYxrBnmQG4nN+OlZY
0wjEUujKr+ZkpmxdbKrJDiHuk7aGeiPQclUVJpYUfWEbC3qPrIa3LImprquHjuIm
wS6vcmejEipk3MEcUtJdZFDCpY2SqXiH6xGOpbhRS+kP8z4Q8EvV/V/NiYCccIYV
PbXN0Cwsmjdkmsn9p30UABvN6sWQ/Yaqz5B0lUvgRCwEKvisn802oyPSiTgkj1V0
EIclVd7CzUPcK/3fj+5wTw4/iJrE7FZnzSkaJuSrQkPAO2pDsP7CCu2WSss6eUIL
lz1OjoKXZc4TGmctr5dhXVpimEo8HgAGnvFWT2geGqxzTW5WClE2KU4zjMEZb0rA
biXVq+qQE0msVijw3m2dhPQlaGMuaFaR+WZn270CDWCirJ1UYmfsF37lNe91JH0t
aKiGh7qCsJ2OOMjwNo2GrWYuuph/genOKT4yOb/7VVexS1fTDMxkCfX//oOITVyu
Fv/Vt5Mt2Hoz+yZuvZryyRx+cAa+EmNmfRSYArfYnVUYuowbZDzPBHijC6D9C3Jg
XSF24VsMUT9Um+LIqKAdhPECiJDvtGG0+exuXbJs5cL4eFsDk6wNijT+HgEDaSKO
yUucO7vAeSTo4bZwiNkNpKNsiR/jLhcCgpAKwBZmZYCWY+dNSHmH95JEvvFDnH9K
wx76aaFSFwzALMSXGwceEJiZ7o9v9FqH4UOKAXsQ9cqp+qB6uafBGvmEHpEfukGA
PqMjjlZvIH1QZBSaqy8SYfO0kMXMK7JvRC69g3PaRlzfaAlmE9uif0gtKvM7Hr2y
QIBeCBTlZAZ0yl5zSfnPRjB9gRMSDWJqCR853EZ+hDbl5sLhMQ+wigvqn89TtuF7
wCQHp2u7jbKH+aFUY0EhkyE2aYD4xLb+w8ZygQFlxGt1ngfzp6NWU+xFSXQ/KqC4
qWySbm/P/hi2ZUFljuEivRaOwT4unAMF48KplHKI1C45RrgCXYSkwlGod0djvWfN
NwdwaQK4VPLPV9/KP4Z72tkFZX9HrjqarFSGlvj/nDgMLqGX3wWCj6/y93G19I5W
0aoKwlM2PbJQ6sQWsg0y7X0tzmwDdR4c0U3WinE0q9z+62kBa9ml7oCS2vXo1mYJ
NaxBT4/A7zef2zyt+q1h04ec7eV0mVQ9aHZgAIbYaDt0bNygHVeYxLtqKRztgH3F
Dk5FdNty2we0lPos7OdTJATEqSaYwrvHo95Bx0zIi63mKNUaIkadI8iCx97ftL/L
yb8c82MtCkjd0FYccoD7ilFvuX28+5NXzTNQMbMSgv/VCkmM69CVIOdi3+x76fpz
b4Dfxb1G3UXPfxctOmBcIrV76M0L2cpsnLefYL0aUGz2EnzGSXJoxh0FOPYQ8Axd
MWL0ScNe28o6gk/kpkRT0/Lb1t8vdFz2Q7QbfJ7+LahtVTtUsSJC1EG9CX7S0kLH
SYaZyiLaYK8I6V+A9ofp2dupUeTZLDd56xQ2Z3A0x0cmaAhHtUW+U/4pUQUvmCw9
1RSBNCREUZDlQPdVx/Lgnd6Gjb4xFo4atjBDay78wp3RqBZZWgvwTbmHOBE/Mz0c
3wBkDjS0oQ2jKsilDc4z28j/Ovni53dMZqJy+O4vsjLPvrnJ4FrXRvpOH2SrjcMo
tnadKIZxydZdQe6X2YQ78+TFSPy/C3KI/VmORGFu0imV2N1rQ4x1rAk3Xl65O2tj
RM8RpGvtDiJW9zgJyPZ3YNnhulVtrwn2DHyXuzv2NCnOXaRFRAm2wBUWHwaXTxLz
J6CbUkZojjLKTyNIU/2nhJ4MexDjaarCeKYjvXJB7dgxPwSoJ9rMjllujfHOBqLa
s8VUtyDLzE/+Vc96X2Ad9AHZ6ZXK6wwNGLUs+/grVnuMeu3wjG2X3Zo1Hb3gl3CH
fbwmJ2T9CMTRu++lV2uMfMSAEmEM4Pgw2zm/HRNksk5CdM60UQ2SMfTRMU9/uWdI
VDX+bGDWsEdq5yG9bz+tZBt89+k+I/d2wIwr3uLn/emHp2G3LyNnk8SN05lbZcbN
Kg1da5RVR1Ua6b8iekbUIsNLGr2Brmizkclolf3uLwv8k1IilpUoNHW/aK76u/Tc
AQF+K55tRoz6BWM67GgOysBzjN66FGNzcLdy5xIDxwRpHTecZ2hsQfNg+i8YnwIL
2O1rFZ7CbyOtJyEDoNLW2xtLXG/ynek2eMgCpfioLQ26uG03KaktdGlqqyaJYGya
mMj017MPmj79NnvLxpVj7syurdXzPvlCKAsCrathdfPkSNO8JxDX1rRo8J0wU9sI
qVA7n/geCJrqgx0oAiO9VARpANipKCo3DkPC7s+WTRlqk0oHtlbAADsGw5OXK6aT
Bm0EPs/hIzQR/+H4hdlJ8nJfQSpGUGHZrrt+hyW1dZfpfZ/WFgEkxtpundVy7bf5
HPE7wv0YeWm0TraQ1qSe9ssKRuACe+adlEhD+ffsbvn0OQcafs9kXIpWLmS93t5n
sG4Dj4ev2PAn2NjG81m6QnUGIiwkyJ6MvTk3R5a0o5FuKNwbM2EeCEivqlyU2MxO
2yC7U8eEO/vULnWC3Ut5IxArIHiN52SOWietGXjV6KKfTZzVOXDMFQLEoEs+bdes
GctyYM5PLuj+AcT0Vn8v/8rBMb+wL+MKt9WOQW8klcIqOd4G9GtcV6IRJHoVz3bA
oUYpW5Ia371Kzx6YGfjpLTrlVt/fQxNKqT2dNWLjsifQegFFFm10vOaRjtpj2fYV
5CKBnC34+pI8XDL3MxsW7/RF5L/GwTdUyekWQZ3hctKOGt82pSiOV+FnMO7ske9H
i3DgRAmyuICwgTva0tDZRDI0mIbUmqSn6z7WpveQSvGvYvKH8tAK32XXLuuj6fwq
oCiadhX4dtYckWdnARkSrrAA93OsGsQcJ4sqBStAil8lDXSIKO3QXx2ANnH41p8w
A3PrUjL7yez9yGJAwi0b6p8zJe4S7FHjMG9mQdEwHWtlJPMjXOGsUqxDkEmJcfpo
SbNTwtjW6SFrFgizFzNpLNEaDzsR/cdSGy+2J58evnowd8rT1gFkevCSOLgQ9/aR
ObTGGcpJG2g46HfskkGz7pVR2oGRpl79flLLC3dYZ1PKSMNcyNyIeMj/IxWazvAj
Nfh0G6GPAOrj0UII/8OwwBPCPdfhvokct+nQ0+f2nnvjokSMubONmJpdWY/1SvtF
hwRPy46vmkRGfaZMFo5k2WHUjU1Gw6Et0hluTA/d9qU18FGz8cJz2v5Ne/GmjRud
rqObalSrluy0E5LAaOSFEhkXIoqvXGrBtV+RpdaRPZqdeR/hcQn9lZDjhInOvsXy
21VaPswbO6jE/3X6xQIH/PcVZqHq2/nWEH2MU3rll1noTsLTdCbGjCsL1lVwsS4G
zC5GrSiIcrH5KtKzHFm8UJnAgAeCn2sXBUsi2N3XSW0vsUzWQ8S3K3T2CaOqURE/
WtM7qPys25nHRCPBz9nknkT3Rtkc8bvvDEzpcqhl6HjMReOm3FC65MD8Ln8mA2jd
0vUUAhaPGWD10zUk2amck0zq+r6NQUwSoos3WyHKoE+8ywldXPODpkvLPchGNce0
qcoJuQUDGGH8zeRRQrDuSg8YE0RrJou8+SS+3WjoVD+iKFlMN7GVNFPJCfpXte00
JTEqLKI7Ru9415yYL7OOwnCbASvv57ZAZjTdRNqIOmoR6L852dIjZA/UX1gt1d25
CNBfwBaowc28mzDpC65oHiHLt1SKbsO+FgnOq/4UAWqEYj6n0pw+sw/TZcwCKVC8
pTMn93TjDvRMPBVbskPE9hgyZp0KUr2K41ZutZW/JxBkH4aHi7BwQ5q2LgyKMaxD
7iDlPw2QOFWGahMQ/YLCXuEcMgsqqlUlroOsYnzG0Ilo2jlrqfKybVRlW1hdYQmc
BM+lK8jIURKyMknuLQtMI2TrnpQZWdDSnC7bf2243VFhlo8Oks1R2miUIltPlhux
9IoR9RQJTspQyStU2pKY2IAcmJDt7o0Mlo4GaPMRPOTeOHmauW1V0YbQpBeaQq/W
yfwgBpkh/v0woDB5qx2b82ltyjob4oMw65h2F+sEh3uAxxkN43JzTbP78OmDoGy9
XWtf4WCrFhh+fgrGGr3vwm5GDbBbA85U6YGBV7sVEJqeLRKkQGvQBGiyC3xwSYyZ
qbUev0vKaCwKHU5OoVDOSGeNONkBS8+Q6uWYA67xUDl1GbCg+02KcAhMAkL8TTrn
2O+Cvs8egSVUYi1NgDmnytdedG95PGCexSI/4hNlDEAqeWAJWArcDorlGUDLDKD5
bGzSHoBhXn17FVLnn5te5JMakve4j+GGPkZnsgc8AuyCg/bpFAHRj7EyLLDXwARm
xOFBi9ELvMRSLYHsP+IY9Hfp4nVWLU4i5Vr6TBZX4XqGrw2olxfyAXxv0gR2e2kQ
IT0rqwzGGWcQ8EH+Lund4t/QUHvzgV2h8uFC6dAcduLqmH/djezZ9e2uj/zLnhT8
AbZv8oBHSg9Mn6J/fAjrI6CWG7pqQjqOGghwnbSKVasjqDIsXEz4aZvHSyzd3tGv
VOmd8VYmmnsMAPUPi0EpcKQdfZ9npLIbaMZq0Pk2NU0rn5CWDycuTixeDnUvdF4v
W9tFVzyDXRwBsgK+kWPhQ+R07KmUqimy9n2ZpL0lx9Rsa9Nk55vBFVs+E8fMjIkT
urRv4u5lpVnklc9pxkQpZN3GZ3ttvcqw0hWoTzhe8Pmm+OHX0Mp1f3VHhFF0Ph84
byZ6+wV4vTF75x5kxcwFevgCUiddqdWicnJIyqUdXUZABrynUWw5VxN6vl7QSIR6
UOilYYnQu4iU33hplOeBztSG9+5NNGZ9vRF7vBgsqjYrwcddN9gzc7DC1KhcTrt0
eY3N5+B6fuRXknYs434maDQLqgRqyBOyw1XISd5Uli0MTH6T2E5BFhedaKvseVnv
IDeKMwxP4Lb6fRoQ5Gqwk5cgS3VMw62u3MErOuOkTOQ8/m8FLxZyltzjWeqLKJOw
xKKBo8cKar5cgasPN6Yw3WQsXyHNqqzo9FaKEfsXnMrZ+KpE6MoNuoURZLqmZRta
3lW9xihbBZ3cuRLmuXqFMKsdu1JtrCpY7YI9brxqXEMcGz28GExOjjpXQ3n5MnWK
qUOw0g9W0CWjspUUjK3qC36t0qeszks81ZiXDUiixnWChnia+LAS/K7gyEkAVyL9
OXPt6ivTnTi69BcSzsYWzMgjCNpkuNP6kUkpVYjSfDTWLWApVy7oUqekQ2KlPtdr
Q806MADTdg2zSaEfYw93I6NFnb7ynyBN++JgvZ4ZPKXO+juAG3zeHYMbnLA3pR2t
N3UCJFjEHl7NuaZmgOcR7Yx/8AcZUR62FUjQnCu/+02pkVuAYIILTdNPw1shcKeb
6kegC+xVBkUP7raDqja3TXAQ7ae2l2HTJnHBJwj9svggGmT1HrhoqGsXyV/1FBrN
6eJ3u2FWmlqciuwzb4JjVHFBE4j3aNnHxk5wCyOD7ZKeis31x2ie0C90whCAzaIG
zcSVKVKtcJb4Yo/1DTvr73Hz6O4lzhn20327c9jNSQMQV6eTfKkqugOx+UxHPZja
mhuGthZjckno8RZqz1ffangtR3dy5merGbulz3T0clltmAitvV89XOQcVUva9ZNh
1+/DF89o0SWb3eWpmLoqExBAM1WcdK4T5KZeZd8yzTfSJ8Oe99jPQjH7OVslZJJM
6kIuX14MOsnBit/lNpVcUoZrEZLdL0sItPGv+UOuPy6JnkkUdUzjiCw7Z5ZiNRn5
w0tkR2GLFeuIFpsNq22zMw2AB3WyKavA3ZIaCy0GdHU9fL1RAOX+SeDt6uETf2Xl
e2b/wMkmRqe8QnkTdNyr7QOSnXFB1Z2ogPzTvEVNwNzZxWDWtssD3ib8FvPuXU0s
`pragma protect end_protected
