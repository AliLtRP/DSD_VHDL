// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:18 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dyMHnwPfRXoiG5iFKRTdrA6pF2LWCVZc0+si68HU6c4+lyT5BVNbBCGbCvQkbmJT
so/P+1tP20FlxYTCVs5hpTKG2w3AJdDkkuxJ9KUAZoYKhqEZKk5nTzrNvGQqN2h9
luawFH6nsYkixTQxLysSrATIXJ0uFa5GyCltILmjWiA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3248)
rVcdow5Yey7aGjasp6Os1PS9vIfBCMR/iiLiIRkGduDymVgO6lZCZDOdKtDZcsLp
UCzMCSDNp65ly3fHdMW53yZHi2xMschr6q5dhZ2m37AG+dodQ6jmAvwPdb7jlcuj
CZaC4O27g3GQDLN/HBXe3xM3ZBlDSKH7ZtsLjprn4ZlSxOp359jLLReZTwX0UMhd
4d9oAn8oK4w7DoguIuz/FVkOj9FCjOLk/rJKodt+8HWPybMTQaZeZlDvD1irA+j9
SNK/ofSFUNdAQ/jMML5wos5RSQfhwXD6eP5Zk+UbfxKJlriMTv2ZnRKPqhz9TL3y
F4gHBbyshx8s8jea7iyeWz+XIePpgJcPlDqs5OD4E3tyLYmjm/7ORok1XreT7Cbb
hFPW6NLmkCINzT+3kvir2H2Yz+1fKocHrCS8T3HAE86d/64F1HK0SJEF+4nFtij+
uznMkasOL1fhkeuS/uOLXqiz/qTFijXnIP+4UbsTuGjwk3u2OyrH47+OC2NPhcfl
LUv9bg/h9fIdmDBDYEC4UIrxZtPP179Zx9V8gPIkpbKYMPJIWo+Egg6qKmdvd1gE
68JlGxFyjcz81kujbImmBj5vEOT/goSP0DfqcOJgDHyyAThl6d87tCn5m5azARsl
n/rAXbBKJTO6UUZgQEidHqFUd6uIZmJGby/tewzG1kJkONkoyLKsOLJ7LsDRq3IV
P1kwuS1kRlzPzuRj0f2E/VHhRjb2Hpvg4HwRuFzGf0CqFffkNEKsDhbdz8d8KBsH
iwo37DTRbPLApVJUgShmfojEAptbE6eAGLb85ktv6fdevLMDSjaezbAUvsHIVpkw
rzeusHzXxMBho6xv08Oz0uI8QiocwmrkZ+JDBEi5aK43Jal7CS1InV9Vx8sJOrbt
YnUZH2j2zfCcipBo+5sGLsg5gE0PEL5V3HLtMoyYP3rykkdPU2xoIt6yibTJdNn5
4yF3UzIQoDol10dUM+I4EF249nzIa8ESCOqJwfiKThEkWJPNn0LzCMEkyYsDqTFb
giibybjhuCSOWMnO8CN1P6CRDB2Sl1rA6QGuX4P5D4DBDtiljV9y0O3QrVlHpTju
s72+EXIwW8R+LUeV5NFZA6B2Yw1slw5i+oAbcZPE8BcSMr9Oyjmw54N9IkvznvRB
jHpT0BW6hJ04221swNmwNgkcOFyJN8IXvLg78KtTS8sPDtL19eGDch6y++AmF4VG
bHcec0hltii+JQPLa9+KTFjLt/DiIvrPSIrtCpzCpHWJCpPjru3cmi6n/UFlJWSc
hKf0OGt2E+6vLIvzXEN8ARGygWZYbFSX8rRd3psyxN+8HNt03JDmP17admQVA5Yp
uFDoipDPmuapAChjcKRf0+vdXeRGG+hzHs2+13fnV6v7XSoZfF8rlspckJAPYbud
yRuJI38fvYp3TJ6XTQVMWtwg5d8CSyLCBENj7f3AS6awqj49Iz4pYG3eY9ZBlLh4
rcHXyebNElcGaemby6heb/PYFLePP9bvqRw+g4ttSDhixliAcyyF4q59jEGC/joD
lk8QxwWuS2fi4aFnh8niF+PHIXx5OMJT6ZsN1htQ7kD3nkHuHvEr6DywMegy4yyZ
aeKODCBEtraLzBQiyf+5JD8Tw3mEgQzoNwXdy6VVIfiY3iNIYXpO8cwCTNRct5Ca
ccdUR2jocNpN4uLP9RTU0h1vsdMIW9QSXMt8MeUMEuoy/K/RJ4O53JnmsvqL51qy
E3dQ8vih5DMgDFtd3NFqdM2AoIyQDW9AG+O0yfzXhPKHWcfmpeRjzikWD5FncaRD
1kaIHGZJZA0QwA+fb5YMgJJIliQSzQ/UV3vDE2ZkoXY9XHRv0gYw5W3Iny4sJt4K
xhW4EFaWcaLz1HXiFWWXEPA92/oMicVQnx/ki5N/sbr9Z0HTpdbe/vRHr5xVXwVC
yE9Kn0lGeB81Alrr5DkEgrNG9hUo39dq3EQcGshMCIP8yXtpNojm54e7sOxwvXY+
gLcVzoDykdCAtZihZe9ctIfAEpmnQJ0i89x84r6sESXK8m6HDIWUGayUNDwvuh/W
cieHb4DxZ2YV5t0PWHBs5WVfOO63hTueybr/qtgRr0dVPU5fdTzcyC2fC1CAd0UB
ragKUag44fUd/w/L2oE0Ly6jQnO2BEEUV8ZSGKDoVQXYyANzN5q3ydLXWcFvl1kq
Ryf1Qac5oAiwNjG/Bn7XPgCigHElZsP3bS4M58WoJJTStUgvV8hE3Z3d2eWrY0vf
RQphMhtY2JKrGAbVZuhR5kUm+Tw+68VshiPd4ZoaR69dYVdEwryygHkF/LDbVXXu
y3q2Fb0OCw41cIacq8w0NXGLT646+HJKXx+wB/y5D1g9aaOWzHPsCzwX7/SysurH
jKICsr5c8Jvex2l/iArGZV1vgqc+R1hTVFhiczbY/QCf2Hkw5pZ8bMGWAEJpI2go
VqPb4erCCeItKmlGjGkgnKfHgXpNlyIvc/L1Pr9KitgS7piQkQbNiuJnYiH6n/2E
j4NO7nUxQnhIWfNUNfkifP3H9e1VxpI2QiUqzdfeH6Fo2+QKKt9EmXyHT+u85t6N
S9N8wkY2z44Bmy697Xb/KJFV2QjAbm7Qpby+a0Y14WMd/A4Rmr4fAzg6UdNnPSgB
haW7hir3nZvqQVrV1cB91CFV8BbR7Zsh7fsA4PopbOVIIj5cs//ffp3JEHXpq1id
xA4gLlnSPHxrv3bQ4qGLj45LWRKtMVLjepeQ81unarGFCc0lleQ2p5VOqSc8O50O
KWgAWDJgHVJGePZkkF5+44ZgFS8f52EOle/3KTW/Vw1N3j8mylebyh2hhWibRA8M
DWk+WlmoihBfT/387oAOqy6OO94omP7WWgavfAb0pWiLVokRb/9hXuqRXQmqGszx
ToA9scgsF2pOOHepnQmvgLhKO2uB7Qu1WRETJRWz5bnguj9JJ0A7AgZ+F2jrvOIG
aQxfu/lM9KA3JwaJ2wR+OdjvEirvqJ4XV4/kPCAb7vhmjDrtbY/aAc+pYM7BQzEC
TMV5n+I5ngGSkNRYary+V0/Wz39RJcoranXTGplbXjFt9XfxmLNrbYSBPxb7xMLE
ovsw5ZETx5Fp3bT0e9pfHklY7exaUBEasMylA7E2d26AJXeWg00v4q9yV5oLgBJy
a47oMhvem69DjIWyTjU5HetYKCaub0hf7lsf3CZjftHWh2EsAWLZHIPR/7tH3FU8
P+bDL7DWlGKmhV34KT06/HKj0MZBem9IiroqaVOclgtZ7gtv7VHZpa5dmC7xYSvz
UxqunyQ4/WdS67QBj1jra+8IXBIy1nYLD9ICdd6rp1jlExaMvniW4Cl135CQq6Mq
pzdAssu8fXhHxrF6ot3vwgY5auYlbYSI0Y37w99qSKjVD5Rpo+EonGVVy9h2rJBf
GuLMGSLZ8hifF/IedFz5IVQTCvo2mLwhZAGy9pjD31oB6XGPW3PGBxHoEgyiB7IR
M8097sBbh+XHNpH5P3tNufsI9II/w7Mego44znOhnGEFE292a/p/apwOPLLdFoj2
MgPjkYYKP9SRtIsLHpQG7Md3AfWyMNjioQLQydHLOgvut0PX0CkxklS5PwpB+I69
b9fUu3Ojf6SgLLinYN5ZhtM58fD6GxtEoLi7SXxf2RASVJgtr/KmZNVYoDZgGWj5
2lMK889HJnn84xR8YAVe1XA0NVTwswV+ZagPLGLrhdrMlghCPc/Evw9EhiLRA1iu
iDx5HFjgHNcGexhqVIt2zwcx/oFf4MA2xSmHrb/KodzFDgPoKmrd2m1127XOMM0H
a/p1xoJUaMN/MdvkdZDRq6yPS9UNsnwPIO27oJsHopspGgShsyK+TGw17HyxiHKn
1ES3uJJbs5/K0icQIg44ql5OnfOb/HpeqPH/Fb+dQ2vBqWtBtdilXcf1dqI4WOln
w5BnoIGPAztWelJ9YkEisn6OKVrahTygnTeZMUzix/uzSG80jkxOgAmhN1SxO8af
Dc+upDXbewYtI2v8PNAJHpM68ZpbHuNbbdC/q2ZS+3OhxDN23SWo+jv9Y/sM9uDR
kM/pY7QuHDWm75HV8VDwYL7ibLJHrb6AC6skyqWYDP8ZgijSqbo9lzAcWObxCRfa
OQE8Lz34aoR9Fb6w0Y+nwrED0Lnu8W8ntphrJFDEltzF/VXwGMuxmLM0oYFTZoKJ
LZBBCIoNzB1sCImvXrFoWj68Me3urxSPEBh+CmpVYj6hlWS65CSPvwrFQdKUUWqI
taWHo1KtArD/iXF82LVLJZXfw0Q3J8zFyFef+DHVZKSUw+uAz/cDTTrMLWi81CVW
JfLq9D8avCw5Y/65ro+p0aNGXrOejg5z8JG8PrBdccQ=
`pragma protect end_protected
