// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:10 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cP5Z8rGJaD/yqi4J294cgcILzGL35/lOu77yvNwIPE3WJfml6j5UHkykmsZ5v7Dh
sd+a8UjnAFkNwRzJIz/9iG6Iv+z6D1Uzv25fi++AZ8UKvfJWgMoEcFMK/jNPKOiz
30JzgqJi3wMwxborDN0xLVxubPlYkGDgrqDPJjvoQn4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 41536)
D6GOk/t3KmuSCrzt/oASQ/aNzFBi6vL96nl+CQp7uLA9hJzSs7ltf0GseUqvZVEy
9iA4O+DRyvvaZevJ5CcVlJLKVBn/EbEytz79mHankn5jp5fm5+YV1ePYdPv1BuWr
NAYQGRNHWb92nUuVjZBmiH4sk71GkAaDyYA3d/pjPPHy4yixCECZ23gcHN0EhvOF
tDvNjG8L+ThWEyJRy5C0nJ/whjzJT1kPdVHI/rCyLiiMiTgWp6gLs4lSEk1JMOcY
ZIZXzDfNT4gp0mfOh4dtWFnqX8jAYQ4xQ6iDbfEbWi1Sp9YQntRBuTdS1LWd2TuC
08/BOijnMWgdYmiJDikhcdz7HQXt+ePA0kgRnlnPKaSJEOwTfD+M1CPkLsWpRdLO
ofv+ZUGaYUz0iwOOwSYYHHxZhxVAPqVLeqDxxiuV+AFly5MqOHK5sHCnrbUvNdTJ
iDSn8wAZY8NN3k27r/wcOCMbazKinH0AzbcxGg6olNgVsrvVmuUkF0whkjfu3NCa
E9jl6FUDHKYdfBnHs5px3xXOB4BBg4fG/u9OaJcRgp7dMcqFtLXSF0L4CIlC3tHO
cGIRBt4ZrK8VHksjiF0zVFWCNMP/jY6LejOQ/nR6JYmkM7QTtk1Znx4W6J+Yc7Ts
eLp+0ocOnLrLmuiu6GBr2Yv5YSfIVCpKNCNG6SB9ilI2YC+KWAeA3RwMSXM+14kO
cWklbXY55VbVYXZ7KUCWsVmb3FJ3VdY/T2965X/4OG5p8kT0mKCdhMrhQPs3aaJq
MgSRsLi3CeaB64yko8VKITZqkmXHe6ooR6yaP8rWwC4mjw+aPupBWzczX7gy4gbT
GfnST5hI09wkjE5/tm9ia6TDeWK+zvjb5QGQ3FuXDJFIn0HPfdK5qO10nSkLTxp1
eNUwDisETeqpiFDUREMLW4V9gRphGBlxsyM0Kd0Xj2Mi64jsvR0XlE2IngfRxA5E
2jf41HMd+144ZtAX2qPqc8tP+Nej61yIalDOMnOfG0f8fns+m5Z21B1l12aQi+Lc
vgKI6AuJRCMrAyBK/hXrGHvppIU/KkOZuZRSzeFb2k9Dp8LXelmLN1yq1Z4HRRh8
M7vcUT0fVYE4e00EEu6xR/erXAxuhYdumbHBvlZ6kNLV7B669N8lYaZXG/m4OUH+
BrqOTBY6DvcrzzV/GE2hVME54fk5snmhAsK7PAx+PNdmBvSgYke9eVeqdVLz3g4Z
kHhn73uXrSPVO0KwYiXAJmyFcnBQB1dZWzDvQ6wgSOmYVh0jHdsB8rx1ojS0mg1U
Ve8plo5O98fDVCAGRR3u9/YvHIc+i0mxX3i5cG5eJeyp77i3kMVMbmHqUk3o1BxD
kM+rhIiZucY8d7Wfcf1UJqdvBE/3LU8RYR+zGYs5N1b53+UYjizI/wbiXepyNy1t
YD0OQiicvkQiEJmR9819UcwqgNK4rIyZpHKvUq1Uuf8dW7QiQjMQSqu+iMui3YNA
mCZbogi9Ei617/pPelaSuxBxOvb4KjTGg+4A+Kn+P7G6tvCCAWs7ITNJjzIsrClC
ODnTSUPQ3HEvh+/EIcpjxScaCJ5n5nZ76Z2Wk4Il9ahNeU805X1kiAb4ScTiqrDx
widZ3o5iRlZc0uqJewhBoBzALAQ/7sDhPNWtwrERK4dlZEghla7dX/+pKUSKO2ya
cGP6hqyxyUWmqRJDoXPAi5dBHzE1n1vHMJhA7o7gu1EVevQVXSc5EmDBEM5B/X4k
xaLj4Am3fRwzyst5dB0xPSHEHwrt8wHjSBami1R4ljX4eBRTNhK2c0z4K44IhSiE
6dpXBXR2mRf8q8+keLEansSKm2iqfTf3XiRoRUsc4dPpecsbqrdtd8hML583zeaq
M4EsGzDgJgX+QNvtULzMBexqDf3Jf82laO/DZrCjazEVAgIEk68EQLok5uBE1VIx
UlwBJ+RwWq2vhPGojkKPFQZHXGBr2SnSHCzFk+lDi2mQFHe5hUO8WCMgF4z95k70
JB6jTCK90ytQKN/cx1xvJ9XxT/G5coWkx52cQJLO1PYV0XBPVVTIUwhAR3/4OS/R
DAB6/cNXV7he/SKavwwv28vBUU5Cp4aIrm4tCRVD7Mrc8j+ogID/QCgRRPQJXEj6
Mm+2oem0C3rjKt6AoSv5App9uxvFzt7z6BzCU725dGLXLjEp/bST4tLm2Uyq51ke
2u8zK5iEv8NSggpShUNYV3L6guOn1oqf9ZKc0RNvVoz0wajsGQ5WCD2MziFHUBdh
u7KNe5eTRiGrkMKtq8nA6tFvFpIA5aK9YzrrjgxXDHdA5/YMIjHChsq/PSexRIti
hrlcbG9BMTjHiqtQXhdwTDGu4q+QpamxTp3stlYwuGYXwVqmi+EgaG4BKxMoYFQH
+7e4CIypA8HmW8/8HASZJpWwuYHwtnuYG+be8odKqTXmojGPwv1rEQnPnuSWhPMO
AKYdVCby0RiCt5FKVTV0W5p3llpEnyTlFjnCIABS60tJlmaiy+iVkTZBE2ij4nGa
xlaT54fm5mszuUhqEFeMnxPQwSYrvxpp1AQ1ed4+uG39xa0VZK00G9pjHlZRYEPK
3bAOgAff944/eZJJFwelDgsFp18L5Ewz6XPzePlbxH3eLBb3Qnl7iActxL8rLzYl
+8bx3VHlS8/L62fzhU5TDRHVF4C1Tl2Cg9LxlzQfxTI6Ea8qISvpk6J8qhlm7Hxd
mxA6fgIw33y6/4Sgt445aU4GbKokw3SBFOV+XIrifdEw0sIwkW4NCGG2PV1zjloU
YmIDVbH/fjCn5B/esdJcWnlq93TAPVXPFnGLwSr/DdOv+zEApkrJa3cS3GLxae32
ciOVNl6J3w+t6vFmvZVyrdwPVrcKUSfgZNE6rYegSS0ZXYKvktXDyUgC1Ga+XZCj
/7AFPSnKNCkZvzxc7C7W+gsSE9dxi1sjk9FyL0QBMdkZ1cdLkB2usVIEDcbo1x5p
trk8CWugOXu6EOXAe87zqV9IMz5jdyXs9e5k1fYf8AtSgtabMbGR4t6L5iU559Xq
APU7Jf/HZOAMmzXJ+AQhI8Pt5By10SFH17/yQAErkHlcgUQZ2YqD2S5ZmoS8o/Ef
6LGOkN2TbG1NO4VtsR4HUj+OobkamMhmxTGbnqj1Pan6p70Qnx2fDJ9Nkq1SLAFY
Xx31QQEf60W2L/ZzGNHQMhtvK2FngJpU4n0BOYnbCW+azcoQOume4NLELDBh9vsj
q4jfSeVsp6Vgi5TAHEObzNpyN+6QsmyBA3AbEsuM7al8ATMDXmKP67251JysNVYO
0cqP55HzvlUYHlnr9MacfTKVhXK4ITb+6fcn4qvk7YYxYLRqMBXdmy4hhli7Jyt3
MCOwK82T/6VcnW3mlF1NbqnyhJ6/x/GsXbtFz3UbUtMynH+cotS6Ks32Adl/1YLN
mKStlJs9xGRdO1WToKDN8yg694VDhh24pA9wDTLXVIKPO6fhpDtprwzMCM+NXbTx
URmenU/2zd0F6mX2/sAkLlUxJOy4rNplbZmhLqMqKF3hvXR3OAin0dLWbgAGUhDg
zLDBPkh+hfA4tWz21sSJFXKR8kIpbmDXaJHnHRepgptiAgsZauX9gKw2H1q60Zy7
wvhzcSjz2K8EmvR1t00tBdDwmMkVZQChIVTUAjiETgGAYp8693dIn2qL/Qs3DikW
GpqrJTL9SfY7foFn6AOMuWki/1o6Wreg9bJMjX4pDGYOE7sNeiLS0+Ul2sLTLqIN
CB1hdp0oIPS7VW3QZkEjFMnc18kYwRh6ILcldv+CitULjOi6QbTcnQniMJqjEDDT
grTGuxk+OZ1ezkBaT8oU3qVTbHuWxJosoWMeCsbVCuShZ20Da/9yKDxA3V9zcxNz
XxusOy4yKcQjkd0WSPVEBs+k27Gkh8/VWoP1s5XK+sPKlseVb/slsQqCPfXp7X5L
NgSJ1gsbA+1WDWrzfG4onju3Hmcqrkztc3P1VUwTXKdBJ529lPPO8QMuDmDjOIYa
RRv4jgpfnqP8//ikf6uLu8v3ru4CCA/1aBDFTQSxG6MncB5lVB+qacqHje7td5JV
2oMgVagRgs/FmtDKEpYZJm5fC9J8QgxY4SQouHfGJeblbpn3XicpXPx1IKfLm+li
3+X2kSSV7/TjF/pB3UjpDdl1Gkr7ulNS41fcu9Dy9BKhkPkuvnDVwV9DsQaYbfTx
RIvi95A/0ngKRZ743I6avuTlxSklzcYgtDJhAml8pKfQQhN7FiyNSqwArBoWH9/2
ElB3eWaAjC1fyJlQZVIoGJT/2149YqgZBN/nDbD5IvZbyuOGu3fsgp7Fr40uohhk
v+Ou1ONQoB2AXghwwwbdNAisiknrhQFiq6K5i3g2XxkUgkQVNb73Nl8SvETaW2QA
uIfplI11XjK4Zc5isjaidL7ZPq8K6AITvHez1ulWx7t7Kaf9d4Y1badLXCSR7+Or
2ZMKx+gvZ/ORrnaWM3tnvrNrxsraKDVdmm8wvrOHBmiLMgzmc7zRa06I9xoI8xXg
fgMpGFZWNe6PnxAOII3yDF4F76vZADII2XqNFu64IP3NocdAnXdeXUJqj4iVA4hB
+AdAnPNePmRSWA/N9XYaCDet7cNF818OPPAzpPH08ZRl8KguJzB9PHE1Ck6TYmF5
niPa2eCz94OP7b7e2xt52PDTtsBSCfeDBCc0vQrrPj9/Rn/eeGWOtRETagb1M3KP
y66+frQu2wlzsy160fCQIIpmFPzI6uSneh8koNVPYGQ5pwf9D6qQ0o0dPdVBVj8T
6HgyW72ss/t5xr1ShWSdZyzD0nlKuLQ8MZ7Did+ydbIUazq/y62CSCB9MUnmkDpQ
YWOv2Xrz1Wdc5yHCIwJery823mMYZbXLeVkAvi2EdigUCfVe6vKWJqpqW6mn5WWb
+uLwOHYWWd5vLIgYIOLYnJuvm+qeSNhx5sWFG+fMeD4KbaBjRyEpfUR1uQ/sWdh6
iutTJxlKZV3/YXadeBHjYGCMhGAizraBB7J+ooUpAdrmnQfemkzVyzd0mkbT6jSv
O8So9NU5N10sW5FB/kfc3WKusnOxfAe8c0aBjG6E0MUrWLOl1POim1KKCgUF5J1a
j4I0/WmvUX01MibrFrXSGMfNvCpMdt1LP7i0KdYoMhAVHXN54GAY+6H5mw9uL9A/
yYOcwWz/OPkPzbaTP8zT67rvMONmf0Qf8RCsdAOb9ATB3QhO4T2GJRjJqF4GDTBr
tRnMVbviH7WgvIjhqvQLC0MIx9WGJI9EP595AAB/I/A1FBVZJrr5QlOhPYqAxTLJ
SaGAGNKLMVJinNgV4OabfKN0kn06BCkOPPQpp9D7hbAHbYFA/6vieaX6sG6OIcRp
SvYXyAaeZXbcTOFNYivGiLNzzF42T68zo1nBdcO5ovvrh9sMhTuapkAuGSfJbOkP
0ZUY4gpm0JMUVRZRCZGFZ0ZwQC6daDqoBAMkg6Xz4NPSkB0QXv1Hx2/awAOd2ilf
kECt0LHRt/T7AGh+xqXfcAjxgvABlkVdh8znkVk9skv0BWCNRvQ3cDVnTu/E+SEX
N44BNd7uOAq5gmPvUs9/foS2aBeMiRF6jOu4KqwzO3fM7wvaaA3c6ziVXW2CoS+j
F/zaoItwtDfh+W87dmdp3lc0IDae8cN60MxGF6WMd0IuyonsIHXDpicl8tmP1gQW
pekTg/tO1wLPQyctNWBHT8IXL8lIehrtbtp1w/UkDQ+RfJpHnQNUNq36j5aMUS4o
55fntQvwNwt77psnsGPuWta/Dk3qnOchNEWR4q48SMHBrTw46wjYI1PBoq+zHiJi
ewJSWuCVcktXU2A4BlosmqsmNG+N73ET8pEjbbH38qUYUpHGJnlMBsroAv2d+5Sm
33NBZ72hw7mNGxM3PB6VOmDhcJcoAq5eG/ZdB5FZVn/v2naVgVUzcipj5cVY8kKH
xrXg2Wgbzb9Niu7ML01BKdzb9EQLrYCcGLUdGlobpscTqSdWWEl7G8+vDmBuZSAn
Jh+ZwJQrkZCr0igVuBl9QZc5fSWqKOvxOFi5oR6RZ3R+BRZ/+az2qCn/z0btyWf7
z5HkJe41eScfPyLEyhqteim2UhHlYQUZvleignobT84Aht1VVa0/0XtS86PCsYK5
AXei+0ukrBnJoUv7l1BI0Ojwmlx7ln3yqTNBfNKqdM/gnBHta9kzbgwuVD/bCmQz
Y0rDcNjdTQCc52IvB+8Z1SQ/ZeE5tVn5ajXexWnYp4u9rl1iSn6etzlwsgxSST8i
zmfMbLDCC08wkr1KszY6qvHdI8KebKPGRzR7DA0WjEcAzVIe1xPJjagoHAfroonj
rd0HILyCWYS8Kp1AlMelFpKA39ISvk5uvWGwpMxupNgdE3705p33c5AXF04U1fZ3
f7l6ES2RzY0kxRF6d5qOhdd001nmJK6BfJUeed9K5bJbfd1zA6b1OmntEuOGuna2
XBQwKDo5BTySr5HKlxj2c7dm0fGmbVglhU9huIQTn8mV+xctuQI7UxI5/JZz0RCl
4lj2FhZ22UC8t8aUP2WF8LxSE9WlSrHnNuOP6mz0oX9yw+iUTNxZmIATZkOhCrG+
m7V1JQU4vTQbK90gs8tsfTCQyX0FrmmkZNy+LsYEdykun71BRvL8xBhISlxSMRXZ
LIIhxOxX0qfRZnvCWhO4v1bTL29E0BSXd+N+DgDnQgYCR/bverDk690Z+uJAAGiu
//iXYeV67xs4KV+Yf320LGguF2Uq5WfQLZhxgOyi0BkJIurX/jxEbfDzuwt7ijfh
EqyDX3hPaTp8K6HhBK60E7miyvOgzRBnFAAVE88R8If/9vZh10VFmMu3BX3DPsBq
ReCoXZBXumuXtY/NnSbciUkrtCH7BJMWzZ+CZxvSYYdHarWi8GD4KzHcTog/nc+C
dmhV/ImQo+jwTbTSMAp5kc7GE/1em4Yf7rCXj9Evnm6YYAP0WwLlEnCuVh+SIWqD
bJo+PVdi4EozGaO8V3QGJGIswTFqNtTVQ6/8Z+VLly1ujNv65mEt8ED9eHW+yFhP
BRxL6XU7nZV7Q4Vc0LuApUQ85XXLfKx+jLT1Snl2lDFxv5uU2bP6ODIqJ3cCOyhV
txWgY/koXC7tq2BUGgI9MXBs4VeZRS8JAQ1gMwQ3CwXHszBculI0Oj7zMPdkyH/9
vJif2IX9exnrTcA5jwFRQGvpqv1gWd9jIioZlZe96uWgxn5hb0cSwakBkIZvhHA3
nC9jP8xx62/8y6fL6Lg3GGHawL0Q/E6Fd4XP77RJ8xkl1XXbGVkC1MlsPDQ647KY
T/gQj+vHU0cPUlBiMXE34Tp3/CR9OJBePm1z+uDv/wd88KKiUu4LczrAMcnZbGal
K1TEZ338RuUNGKE3yGY37Jnvq03/zs1hh4NluBPoAPH0N8T4v0tiHkEqvqZXX+Db
hRGjj7x4lSbPcyKYroWoAbg+EZGrHoVIKKylmWxKY6ILERVir3Q9n+yznxVFV4kU
fGrEBr8jwsN6Sxzh6XFpp1GshptOCSgsBsr6SN8nxty8J3SgzfmCxRZ7GhH5TfQC
1dJcD1buxdBKY6GAXfgis+DaBOn4lnzDHrAZkrZsfSX91mc4Dp3hEa0mvoMfOwJD
2l78lQpTx5ID4xOMGpVgerJ11cdXLcRlZ0DjNRFkIpB/h5phtdgG4IQUMsYwPFVV
9WSYp8hcHD8Fbf1pd9Ro838KrthyBnkIy8Ig4qHedaVief/2sx0y0WS+ie85Grun
gip/AaYyhJ0AwmWbbJSnS6cFSICCPelRpHGfaBkyFXV1IKX3/utUGVA4zyH+yOYB
DBrXgue2HbEhcneaPu6CByw6+qBS/Inse8d1e39dWW/g3bqaFPELqq3Z4Veu2Iir
YKUsqTo8sjjm+5U0Rf2ZjFVT/+bcX7hT7tre/k7h08f2lxjaxKvJ+pFP12pOYUpn
My3oQ3PhrGKrpEswXmAoP5RQ/LSqcTZpKoPCUB+FfD4Hy7EwRzJHnEvsWYHL4mrX
qmQQBhkyDP3EZfRVngAX6zocV03F4dia++/DqYu9KeNJ/cr2hCo1wFHQF2cb7uWm
WEiMsO2quYMyqtESI7Z8cT4okBDblbQ3pgIm0ClHn9Aer+uJl5cQ37B6PBknai+D
bi8zvEZRy2pYg1g4T59bUVs60slsbKrWFwckhpJ4XaY8TQel64MbFDBp5Ah2yX0L
ZxqaCa1gfT16wl3GUOTln0PEattZ36X1sLBWcRVZcnZLN6U8ahX0j2zzeAgyzL5q
qGplrqfgjifE/zNYJjeDIdV/bbhsplKjWUXBe/RDHwLnPKSkolrxBQpkrCBtSzls
cq/l4/Tok8W5atPzFKrpMumJfMC6Jce7shBLmtRdaUU6iYIqFeQcLwhofSBPPjhc
tVYrsqgZNzebpOmwZqD/G2QYpp/JBhZoLgQoZVd0lur/1yEuY3PyfLkPEgxIMVAZ
VT2YCIlfHKu9ZmJzh16BoK1sBi5WwWtyyBjPcVtkEzpbbmje6drG3aOXYKKmcfgW
BlCibIC6Z8csSfyLxxfsBCtoAXpwBkXdbxQQUaEmf7paFGU+KmNmAoPHsZN9zms7
0KU3ocUvsNJVNeueHdB9kLDq2E5WCivOPK8WFaVJ/g9ErhqR/XqOFQzU16GFf+Rt
plkQFYaYzg1VzJTXRNawdBdgVySK/5xiAI0zOiJqPnbSnLGDsuq4sMq0bq3GhX/F
wf3Ibs91tcgY6hMcqCXL4fTmx/ugAXV8CbL76p7jW02zkCpFC+3nNgRzNpTRkGPQ
TulMCRbXuRsFq5ViPg5rE2dA1de2GKb6QzrXVs2Rv6n4HPB1xrfS3i6t1OkzOUG6
CcrcCxizvVe2XbbudzXaRX/QpEvux4G1Ide8ryKUtDDloG4WnHYv7WoYecPfU6v7
pvdlw0OH91XSlDl0Xlwg9lFFlqQSIZSkXtIr6DVnHhlOea5Z8ohvbxGNXfagIsYU
MVM5kJPRcxeugsTf7Owa264ZKqvfVmxtY8U5uY/hX3NcQBytsIOlZ8avGslv0R7c
Kmx6FPErG4AoM1WwgHUBDQ6ER+8SiD8IYJYKxVWTEZ+Urd2zY6nf1oTiDnesaBt6
EL1O8vVzrVt26Kfb5N7+yIGzB73RwGovUNiidvgstL/4IO4GlxEUC95h4KmjzwzH
UCd2t5N+aMzNr+lUyOhz5RQ1mHxKqzkbyHPIKyCMYZOXs5v1oMoLq9s9NYYohfAv
YRpdDnRshwFBFqTOtwQx2z2qOU/geHzR/yH3Xb8IxDly1ZYlHCQDH6/9K3bPxHm4
SbaNKU/2U0Yrm8ausPcAEiNjjhntEFMMxKRrT6uKrCnbqgcpMhmayfeZC9ZqSJZm
yg3sHPd8e2PVCrbxe0lq7FyDrvUSLmhzREt+olj8k5Xg00Xj9OQFD3z9r5jhBmvr
JIEybiLyy+mjv5WBAMWyxc1px5W53PjI6iLpMhTdZJUFoivzSGB/eHb/TBaV501e
OHyb2awIsik4Tsp6zotxD5fRHNPL4RwKE62j+Tk7Xo23NQ2Vv+VaOb9AxwYMSoCr
8fkabUgGTeJbqVTg4e0910JdKVbqKmMjdZyoB23WBBAwY2kgPbhEjdtgX6uv9gnk
TORgynHa7NiG6v9xLzHtDzdUdlH1Yr4duCSU5cpQfFnFLxy6jGTveiY4D1rOr0cZ
HiEyXSBdzoVVKM4haLLkSmxTCpFPhbgABTK0V03cmDRslMW8qkIZ2hYr2YwzWq+X
T+bjMn7bDhl9+sbB1Rr2CfdhHPvmbDw7Os3dMCkjWYgsc3LtedcxYXx/g/i7LlM2
bpIYKBPPh5CdfmfLkBz5/I6XNYAgYRLvi6eNl/VWZ/JsJatcOScQiyf+JU/Hrjxc
JWgujxGBNaZzMDXrFWITUDVmpnBhz7xdskw/gQCDvAOO/M5HJJ46jxCsUdhldas8
Ve68rTnooNv1QCsPOWFFP7HfAQvoeQqOk2QVXEcaUfy9TmF4FM6ucYRIlUYAfr+z
8meKgzxxEZQgWSndfnkls5dDPcWHZIn+C8iZxbHQrNrGTj1l/zV6lJUufHvJehlw
hSyxaDoSXrm8UEp5mMKDgAjhtxdTSDh0kNQKOkQ7vz0FlTmh2BUSQwWwFnrDfYLZ
fWyYOKsIhi4BFk64T5Efg54mrpFEoCDsKA3K0fwDQstGbPnaUYDlWnbgVKrqpkb+
VS+/ssW0DqC06Yha0KGBH5TepAY0Ddy6TELnzBmjKjnMCuEkG3ZIG58eUlHdwCMf
gHAs6MKWyMVLYveZvsC+f9OTYQ6Pfb4Gk3brVsl7VcxTEvcUqjxDf9aUj8t3X0bJ
xNwUVzsC83JcSTM1OYgeO//7/KKcYcTue/Ni91dP9WMqGuQNnXoqgF1x88PST5Ip
8XE6ZkDr2l6243SDRTFhfXy+V9JNggydwLcMX12t3xKySJYffHyHzKe5ZChjF8Ca
v6PQHcHUYTRyIJW2p8J7/XSVBl6ITiLTTn+ffP1QK/IZgaxtd0/LwMnAOvL+vMuw
X++1JLGLv94/3WFjE9q0Is558GGodJ0pgNuF2wWtOTuZTd7ecrsWvU6hWYP2Buno
O5lcgmtfeTDKJiDxTBO2Y+90qr3ytlgcPANXPFMPPKJPCcCtQnXHnfX1L9p4DfkD
giVcV03JDN5zstm63/o/JNaHqeeyT63Jx88otIsaDMCYifJF4UItfJoAZly9J4+7
D3qwZGBHTWJkiNTkzRefMnecjPy1ihhjb8dJM5P4E8DTwkOQ/sCaRq5llZPd2vq+
zXcUs9/FiGP/awwTVRvVQ142GBl4Xo8NgeyP+KIRzhJeulGMlJ65nVpJONd7yWfC
1vqzt1+8d8XEaDZuK5sEoomYvGFefN6XjPIZAq5RuMKPn+Zp45+oTbaZBk+d9fLI
P3hY2lfwXKIbFYUpbYydPJ2dzbZ8Eh16BDDh69J12fyVFoQxXiCa39ROG5fTpOnY
KO8NowKgvzjhmR6EIVFBpsZQflVPeuXkpxW8f33PWl0Po8U/12snE/RdoaUf9pDb
3h9jl7Q/jNHEvmgK3/KiAmjP5TobzlQzBmDKtoMCjmrK95nNlBLsMXOfDU1/AsEf
7laMmIqU60q06n8O/4jN83oOqsrb3MsIoxndCW4WiCiqtyl5GE17fD58WfkG0mtN
CGs/av7dC+HcEryCeGIeZWOIV562BMrkwv1woFAUhISOkth0LNcPKNIeh4MmSD5g
kUw6sZ+IeaKxInOPYICN3GkjFSbO7tx5XByr+3WF5SS4ozQnUin0ZnYqakYqfsDB
M6cI+1ohpUUahk1ZCfX8tmWn1G7c/9x4CU6Rq6r73FBrF9Jb98CodN/Dgdxi0nzP
YFknTyWy88Rv1uh4ky/6NeMlB4G2yDI92mnH8QyAQG3bie0qkV+iGDJckYPmfBN6
T14xaz6SWS1bBIXhEQQoOJtrNqzl7TcpxawujGZp9WjwPKsB/+SP2fAhde+sI8z9
prkdQWZ+rp8H5QxW0kRt5m/LjnhaYafb/0jMorbimK6LcEorgznH+Dk0/3WIF7XI
2cWzuSe5J7Zsg4v2KQe5FKyK4ZaoLRbMccgUkL123rs4fUJBpM+FjkXEdYnPfXy4
cV+wlM7uj7baH4lD6KpaDZLOXg6Cw1x7G3Bo+KT0xPMUNK9UYfaermYZgObppf47
vp0PMWOK0Ru01cud/Vjxa84mupmiGZzFGszpe5PqpnzzXGKGNjj9wmr8SH3ZT3Y5
7LgO6GBdP+9j52jdcsziXGF6ZUK9i6HFB5iL9hd3UxlcYgGclZM/WuGSPT7qaeny
ciX03hm1bVYNG3rc3b4ooAnTTI3lmeevu+KtgO9PxWjC8B1gt8lh4YeppCZqkNWq
tCOUPdquwisyWq+yzjvq7kcuDOCes4q/eWWd2lYk+tocOVq6Ayi1Wg7m4w8/9n9K
cuzgdL7cLW65OrKVRDnjc0ogNyOt32dgPsPA20QIUAWRvLSPhZrJKoTT8PvoN2sa
pwnGjBQgVyXV4WFeBCwXdBuYzk/SJUHIaF6kltXPX6492APS11BKPFYQ9TQq93l4
jNvfGVm9VJUqCFcrdjYLkX/XW/ICwJ303V2ewHTdW6KOqJu1SJA+fQRjNlrhzNOP
OmOP58MHU8Ib5Fg0VDdyd4BAgBRUiCim3OUB2IJnS2MiiMV3+zSdHqB+muKYE3iX
t9ypBAR3Q0YlfK0Okkdhw0f99f4PxhRS2RPUsahtcKMAqzpOlHKP+sda3jceUHGC
wMoKkk4vzs8bbUTJHmXgfgdHEdf3gl6rjqu3UafxeVIB5dkbvXf0R5/tDDNBHJvf
BRf/TmqlXBBXXXmwRNolcFYZgHF08vHG6lTnJCJIUye84GiHCBT3H8dEcLINAJf2
Fst5OIN9wzmL2Ut0+Dw4u1kWtGd+zDYhySDQZookXvQ+rZVo34bN8gfmslnkmmiL
MekK1sqri80TN1iRw5w/uTdc6Rp42aJjZW+oJ0CkiuW8jbijDZEob0rNcsjuI8+k
YWlAIkaAfnxY2i1RQ+ocDqsR7XgPzYL/T4abEwb5pZH/QG4BoEc+7kLgOIxFRqZz
zhjUDHNWosThPUR7V8K8sSfVgiFT0U9O9feqbTA3WFMp+w23TPHaUu6GXmJg6DCF
tDT/KTJq6BBWIayQH9lmyZF79MYCiX6g9gvZt0ytndoSIv1dS7KQvHY5wMi5S4mn
PS1Jrfyk7BcfJPX61QwZykeBNHfcRAyV2hwsNCnRL2yoZa2VHuo370HtGTxjjyMS
9HBc/tEpxhivw9jJLwi5iBZnO7QRvFPF3W8MI0k08E3jfLXio5NRpPMp36cry/jx
TDwBUae/NzirVNC7gjH4Iizt4hXq6OpknjAhj69eRwjbi2Shpsl6QaIczzlN9/wk
076GX6NL1xgCpL180VZOZIhMEhJBMT/fQ+pAdwMFOXAm+o7zCvxl6rAu9cEupRCA
M1uCQPj4/bc/C8v9nZ/LZVZrEwSo4b5+TY/PIw5xcctyfHnNbnYqqIKgFK9q7m47
kfR3JpJdhA4o9mL2gTAOkrHWdEneUB4y086kBDxTtpwZqf9HgWH44msEK5XV/jcv
FdVwbKwQM3zT9fSx4XMvOy+VzDq3u60owIwEg21F9N4VwPmJ502UuhiHg87uB/cb
TGoBPxOOVcT3QuIHBSycOhH0EGsITffh9fl1A9ugeQd6tgnJYy1LxvyTPq3nVPL/
mqJAE2jrkDclN/jGaxk8+y4fqFUBvUV0ZNql+BwWxaPypu6ta9pYmAZelKgAc+Ri
kSIh61FYPLC9i9RoFa1fsq9OcFDp5HncSyo0JT52l8nC04nB2oDKy9Sh3yIlgpTS
IbAQ+mNJA75E4EgyCAHBpDe33dtCX9LS/4ESDz3c2tFt2Hoa3AOWAMn3arevyJIJ
O4NeNAry8MMx9qsBDbPf24m0SVE1+ISmgQEqAvIBisAL2RyrqLkEFx/9tEx3Dl81
YiyKHSvBWETJuy48ak9FzHhk4BmPs9LQX7VNDZvNjtPY0GghkQcQkYuHgw6g3Fhe
ChV2hgP+UkDWg7M1i3l2w3llBxfZLv3sBHfZbMHml4qAbjkUqqg+wfJabGZE33eh
r6zOfu9DvCUPXkI5crH0jF+Gl8nduOTNzAp16+DdovVpksVFfjzsOYM2cpt7vLkM
ziSrmUAEkUYQJaRIwHFvwNkDFs3THhghsF92cFFGFcb3pprDW3fnBDTwvOx33o4h
2SKaXbiWrjWuLn6qpVrKwNYKFzUjspl9Yha/VM4mWl6RDvpd6h4/QWM19yIQx/Ih
1odeUbhFMFzjSSroTafT2FPAS4pKGJiOGke8tD1ii4GguI7by/5L85Hg+cAkPN8F
v15E9Mmtpyya5fNhXtwJXB4omSpkJ4bfKCVIQIA8rDXY4p+hYUBhNEw1e3Lpx6Kv
jBh4fDsbsUDVvXEJAOA1gyhsSgBEi/8TPNWaQA3nT7JMpKCwBR81+BrPI/L36WnX
7T95UppgwVeQPC4UT72knLykNjeAysTO4iTDW2Ix8jYpV3jy60Cb1/3X4UzbwnSX
fZJEkTnajVhn09Sa99ofTEFRAT4Q6OGTG6ufTFs1d+LlrUYLVzAuf4XYG81N1KU1
G9nSR4nUYlGfZZHlY1c76+keZCycul1yOjBhRIIuZUeDjvdpzpJa/xIwK+iecxfs
09RBEwXeDiPHYcjonsFC006gFfkBD7THhUWBWc/WHbCdoIgpHBcsCLD7phOqO3hU
lOY1x5oq5Pn5PcD+r2izGC5TiOucCBP01e90OGnXky+rXr3pSH58S9uHNwRYEIcv
TcOeIprX4cogEDGPcXNRrU3gRjYB6pK/LKy6h68huJv9Onrm9ie8KUvlfp/KEjFL
93ZuE8wWBgwlGhnbuNIU+U7/V7HmHQNLEmx7YTnNoz0HpCAV+5Z+ggWhV+a04tLx
xU5KOrI3X5GToknIBanUNzkp/k9kVMJZgt+uqa6ZrjlUl6CLgXyaJCmoJvDnD/kz
4iEq+zgtlvk6TjA7EAwjs+sSU1LQqg2YCp50txME/sFO33wNJe9Z07oJ+2t2ia0p
7i7jvYBF5oC4/6VOs33c2TTLUNNcaX+ZLSFBtjrZBW4TDAHk3TFyi7Xwy0QVE/VF
rEqE4ExHgd3f/WYzbocDiduR+et1fcHeXkMrHOPCCwMkOoC8QhE/ATW3F3f2wCO8
b/xx+w/XtMFgbpkHvkq8ulc6RpbfbER+ixipxJKtDkke5G+oI1RqOech5RqumY2G
y3vF/PMjvIrex0YPzaTJpzp0FHjbIuv3lez0gkkky+WMueXeaj6IeXx+8feiP4fE
T13MLcdflZ7HIzvOh8ArmFd5FiXrtT4z8wcWCFyolRAQMCB2jFTmhECFVWfZsUeQ
++uDbsKwvPabhrQRr18sJSoyHsKh76pJqfNBQ6n1XFDF9+Zbz9+VPPgr85CFf8tA
Nbp3CzMisWNJOJnfAZsvcO/4FGO5+g6NKwEoFi1SxMtTiF9hesfkq/3p1nycNXU8
MOSem09kuBuY8RCRp+h1mhEsxf9nVhWxyfnKDg74qpA7a4ZfEpcpgY1xorLVR/PY
smvE/J/Cx5sweeRIi+ytWKEjwuQK1xCX/ChTD1PDIl1uVxPrAea7gNUmJ+ZG3cn2
SEG6C3rbwyQ8FLl5ThPKccNJYrGkdFEcaSVGWZ1AjptbvpJkyup9ez0vJESteqnO
hx+7O3tBBMcYa+6np6A4zZAsDQEZ2ntETw4c0naeymi87+86jC1ta8fiaA5bIQ7k
LmxwTD57CHXBR+MOQGHdG8dZtp154uRdnwywgrKlOw3qpwyFytHllUjI/3V9XxNq
c0v17zY9HbkicDHCNmRXIgQeWljcKQ2v41YHTHS1kkR8JaGhm6uHH4yC4xtt7ThO
MI3x0EmNfR0kr/hbh49rb+H7k3dsFdM/lf1SZjXGzNzlKaOoQ42O61n54ZN61wss
3hVRax4IwQ6/RkjRwJOmpy8PJuCooySHhaaVB7tVis63aOnLa6xBY9uhY5uv0oRT
yi3Z30zsQVjRfK3IF/qkIjHdIlH9aGTyMYsfdh0fG++HUCRYBcEJQvcF9PC/GH2J
cT8MsHV+31GnyEMG4vrspMw2oboC+jsIACpnAeQROxEw1a2BCj1ykvNDpq3j0GFG
ikdKDweH8bcI98UFkReb8VFOa0laoluvSXlBfBbhlDy2qg4C6wywgiEfVYOndAlq
/ODSlc7iJE9rZfDOHECteaCMXsc+kFj5Jc2c2Gbs1VTSprFOxjGlu2LgNcqwgbvO
GmsnEkT2KUzpkqEAPJjPsWnuQrgIiANPB/JktBCw6ykcEk8x9r7CQjH3pvlY18sX
0nn6S4vGk1nLP8X7c7IYGbOV336YbUJNwQ3xtFOOsPr+0JGnwd5+oY54lm9nbC/n
gGDNAKwkI7opgOIMsaXbeiQT29RgGZcJ7Fm0KtTG44CyrRuyEdd44Vb7OXja8hdE
RPKdGTFympzyFTxjAu4f/mTlL5/XE7ck+XxUHMORZD5IzzuuDzp3ZFE69ngu5lcL
NrqLRwz9xYCRZwm1rxfvCrjkMtSliqzrTJx0IAWx6M6Q+/r9GfYodV0YPn6JcgLB
ooHJlaorPF2Givn9hKIZpG/ydUDWUbGXip/kgECGVH5U0HBVo07gUAmtc+GWfQH0
ECoEEYAWjtwv+vDttnjMPZcUGaBo0OdIaDbcpZSdAxrHrL0QhPiTgg7NshN4d/zg
OEGB6QxK4jxgyaRM1gIWPZYrFVsIiDX37NxGpF8BS/lKOBJzGHED+GErzq/KzHYh
/QxQN9L/Evv+AsQWW4+NI195Pv1uplOGi2hMs6gLU2QGJOk3lCZjjN4/ApKLa6oc
qt0vEewJBXimEHJk/pfW2uBOsKEtfTUIGPRb9qafZE4YgYF/h1tGboDNibxts7u4
2yAqIrP9PB+mPHuVUyMwofz9sgg6R0nnFFTklMtL7MV3d4dyKPCdZhD83lIuY4mi
snI4Wbg9X6q3pPl3Qca8mU4TdlaLCO+Ydcnacyvi2kzrzU+MSUScjHV3Ex1mNdVp
hjo2RA4nFBKdMzRJestGcCoO4cBFTTSbqlkwl3A/UaL/OUwoWeX3Y9J0Mv4mpyHn
mkQz50OcFMWAlfOPMTwtvF6FsCeVVLJJ7AXaWtnEY+XLpw6sjY8Y3jazv0mWRt/E
2VI78s/HPGco+7QAx44OiO2WPx0xSyeErKY+Ug2ANlevF25Np8ifubnr4hFjKxJ7
5b6GulDUUsqxdTYWP/etxkwKDAeVdSwAOVr8qPqb8ZmK1Zcjy6vTVvTQ+Wim239v
4lDbZsQkAdZaj0RjsxTzqTPfNsE6UL0ZHWgF09luxHaKYsryrCpHW/QSI7ArWGpS
4kJkC3BeyG7Kh+FSX8EIcG4BwclDQ5NFidlEpbOezaenJYjJl5pSbg1+Xb4spPvC
zcPnGqBb1EX1pqLb5fMtvIZuRtYL35H6v1epm8X36eFQ16xuL1hUG/aCr491N+IY
ztab2Ds3GFf4vpZVpkcXdUk8QLV6AkQjHyU9F+/ckZi7P2cil0chYp2lhW2opHoy
JJoim+uem5+f2Uw3E6vSGO9zMZye1z5+hhzSiG9JDmqBByX7tUfVQbnnAfpr4qK7
kCMzFs9FhWJ7UJGTnUTk+r0w+RjSC+cWNTilCEGUUaW82R+Ug3WdEQ3hwOVfddXM
qNtMWjkJPMRygjbL6K75whPvjptF3v+vUQq8p1zSL2MRvtwUPwXuWryWn2kCs6Na
39y3lkvcpZIF4zMqbKjtcucCExL6x3bjOtdGSRAI8GxpwW2lfxer8PDNzfiL0M1s
mmexsx6VpKlEnSJB/yKCmVSabMLsHe3HTy0TyLb0qaXim5ui13vkrBmWDz/QIfkY
MQTRXMwdARukEzQpQ0BQuav7VZGyjAmeCvIA50lnLLFU249uqFYtbQkSVWQFNMmR
ClL2kc+nnEtxUA8Wc1IFNms1R1N/E4nQJJTZIQW49yBPzTxY0Y1vJmTTQ70E/yZ5
aBklsIJT5dMB1jY+IZtgro8I51j6lPeTtVlm8UOEoKWwsl6IRITeQelTLiLtm5gT
jpiGKfIegkgui+lZk02Ae0fCALiAJAb9R0ZKqY3LJNcw6uFXzfwsdHKnsQG0+DYP
b0CLfsxZOjg+0fx2236gy82s6QtQi53oEmbBronlGp0j3JvkD8uZQyXMZLplz1tJ
J5EIxh4dEQJNseBYV+hjVIxS0NZppTn05qMLAeAE8nAWu/zCwRzimM5TdOJ7BlWw
Dsd4ObVi4rhMwva5zCgosG4FKx45km2IRVLDv0HnBwS3ndaoXwbU4FMKgXi8tYAq
i6doboxoBA9tjAV5O8dYTF76mKUnSOfJCk/cUGCVqXCSNFuHT8vicdZtNMIHO+M5
40jf6bvP+BB18mOyfPDarlzp7utO/NTSptnM553xvcLKyZTulp2wLiq23QcfLY/I
t4P/i4PKz/7gQAJMPUNu2Dt8X8LGUfwYBCgQDY0pRYLafI3Mcgp9AbDbiEC4tPpL
k2BpGl/mGNPhEI9PkCNswdZAU+oMGmcLzMgoQtGfWQMi9KgPUymzeY+dIRleHNkc
9RFCzKs1+CQpBzvn6VOyy++Ftypjwp/sO8EJyDom/aE2jwJw1ljrO7bu7NXnxPzM
RAsb+izfPwbiCuIcqqk/AAakcnvj6Y2twNp4yWo/mnsgj45ovK46gt2FuUIvEOzr
KiMTcKvIdHEo9meKWXdeYf5Tq7gPSaK79p6zFsiw7Ws+cEgZ4bI1gTNlzAiCZm9O
eB5QW9eF8KR5qn/3fpQrh0UiSmi5beKFXPEh65Et/ZNHVnatA6acje5K+lmIwrsm
Ac9iNjmmvG+74gGaoiMAWQEabPuUk4NMUBuC+Q0TGD5p/a2VsQ2xFWRqOqhdnd3P
+INQ0cklWkZ3kOlkaGNtWEVoQCloPYP4k6LL2K/x274oa9a6x6JqY4fIrLABVaJb
q0ej4NVcA9rT+Yld90SqnSLP9UXSGB/BxH6+nTi+X9sxTsIVau1W6b08AHnyS/0r
LCjsGEL1h/CC0cGPhuAZU918/2wp/uoEkTGkx+7t4BeZkvPSY9kEathpv4sPUvo1
9qmWfu4Qu2GJM7IQXkSvL730hV0CdMpn7cg0rOcXcL90JZ1ceompEQAISeWS/jy6
iV7o7s+u8Or5XffOaOnDZxORqGqKH+EXIH0wMPlojrAM3gEDQVt3mE3Nwq5epqgQ
o2DvhJqe5U77/dD0qIBFdxWfeIpHBcurRJcox3LDNbSGgUSNYD4p6NCBypgE8pBP
dPkTLtfsmN9raB5FV2L0pqpQSr3qFDqyul4i2TFX7Gm1xYLCtRcSV3U0pXVCceZA
FuxSk4dsoIumaayOxQ2bXgOtSaF5S7gZjEC6jkwBMdaHFA35h+1EDjhas1HTj4bt
AvShhnvvOrMWBmCYB9mqNzCc6mETC7IFT5jD4fYFsptehCZ/LmMOJZQSieGIvmqS
JlaLDW6Gx9SGdLK/YaUB+sTbyYj9QQkV9hjvrHL2YgKJC/obYlLuPaiCPWP2pnPb
d7g39bJrxyHkJ8LSwEXHUJgwfJ3x88Z4U8ZynvSMB9pVqhlNi9cHAyvbR/DZy2WL
QTCQ2gLDYohxpcoFIWa/YTejbUmlIEx+QeZiB1dggTPjhdUF0Z2LgZMKyOXI5j+a
PCI3Hcw9WQ91rSf+5Ytqr7pTIAMgap+teL44QqvgB/hlwrx5udpjFkzOKOxaH85B
hDGtziUHv8iQiLxtp5Qt3IWd8IO8irbi2U0pPtAw0ANYj7ylHh7/NLtpwVYYWwIC
mHyrA9LSp2R/EZDZ9ANUKljcPZkMJ/Q2axsbpRnzR2Y7eLHsM0ZNcKKlfcQOLhIv
ch+ZSZZewt46crbs88j9E0a2nn9+IFphSc7J0d+7/KjgPLN+8UX+Dosgik8p4uni
F+oP444GJvGYOvUPWqm7BMSI1RiU/lp2wk+zaS1J7M9qMlnolRWPvH1QGwspTMn6
4FLCk9XQnObAYxkjA7PSgSzgb1eI0ic3pra31fNbIYbEkL6LEN+nzRPgectiOGbI
Z8VLGsTVUjt2h0QXgXjDDs6OwyRErkQsHa5VoWrzVUt+7Gg+hgXKwhFELtihoRKb
lC5k4l6KL/sEQ1FqVNz2WJpbQNihtqEplL07Q8grqm8E9whekft00iurdq1s+M4P
uQE6gi7wd9PAi4qHEcPIjxCHLexoGYpF6rS8bQ/tz4g3HNlWyiYXtnTcJzp+s/Hp
XCLG8tWSUvJfeoWJ6l4GKFMwjQmGO840Qy2qnZ68txfGab1qTAMwolxvCwEtVNN8
PzM/8bsAhWfsGhBZjo+8Cb1/zSGvtmkr96yVwrd6px+zbqVz2PZPK53i9qQ3NQl4
1LbF0SU5npqAhruwAO0VTJyZrYJX9PHGXtJMaOol9dqqbiAOgd8Q8YA+TLmNAXOx
8Wj4DMFwaqP2m1pTyhYsWWPsMpLMzBdxTf9DuJPih13BlqjvcDQaF4SXEDmpeQVF
B69NBe130H56l+e3telTLLTeVLqiX/F1f7tw3xxv7FE8/P8zV40RJFtQs+eWLTu/
RBZNmSWf5zNCAKrloYfexlS7fDfUu5ymt8x7JDQWwcb+/QJC9yPX//iGmV59Qthc
d2BxJxCx2gPwlA2DKSjhVCtjmXtgCRkTJJusfHZTBF0NgTUrxiR0tGuqWjB5ttRj
/CnfBMJ3ibd6XKl9Eb6udnU3gDSowhkJYN/IR7T8PpGectIz7j3WCCY2Qy7Cfpvd
gdtOPTUA5N6CRO4aHBnaL6r8nSDqH8G3GL/95chpu5Wzwb4UfRPkWdEp5UUtwG1k
RCm0uD6SBC1djoMdr46y9tyZcwmB14y446VIMTFGt/rMBxMrz4CNJ9SBgbt5sS1x
dZn6uY087hGctKqVx36KeJp453qit65lc36NlYliOLOZI27ataMmF09/IcATiLYy
aRRCsblqlgL0yLTkZuzqDpexg4HW6fhqPQ+0854KVym6uNljKGuUaEWxeedSy9SM
LeoTm263OOhwXF4eY4HXxj8zeZkPsqDZ6BEY0Q3zVA2PPKLVWxXI8V2kQyLcjl8O
hx8ljfDai5aQN9QviIPqQIeMH2x7WL66a1tEnMxyE8yUSW7g5D2s4Ah702CPUB6R
xOLQaQ8uvydUfM6JZgKT5a5GLq32+97v3ZjPtE4X7ZHP05c6SXeh51/ZPhGX8Ejl
FM6v+eiFnmFD6IbAK4VXW0TdYPz1rxHl2K9TqxP875iHs8gEa2pOisFGslNUe/rZ
p8eWj+tbtpLp0ZaKdM2HtaoG1b0Eix2Q2//BM1X1M9Ulr2bswuO+Orr/04yc17PF
B9+yu3h0LBvOcLScgsyN8Lo7dHtc3a6hsHXM3LIw8qLYO0rD1/bMmq5zVlc8A40n
JsEtB4V0I5/hTMUwsiVohfjqvWBVN+5Ii3BhLNLNzkgtBQkLos1ZKoOSfF13JekP
nN64VZDws8tGvnQhM8jw2dQ4wgIfDskSn2SMt24EO1B8YgNwsinGR1oBJxZ7ZaWo
VUImkVomZwNQnebhBiWZy48uuwIYRAZLx/WN+l1WkFUwzY4SXQRN+GUQovmwXM+9
cYF8RHQLaXn70Qn4rQmDVO/bzwWa3fty3abdlbVTrtqRivvzEt/mkRM2YsNRotZv
zIlOoJ+re7BEdLhX/4N8/6UDOMqLgueJRNOMlAPmb1XgXDPqEaiRCBYQYMdV3IQf
HvtspykBkRy29OpZGsOxKbGYcbcFYNOJl/0HFyqNgOtdYuFAZo6mYw5RvsWVLias
9+lzJ/SK7YgwiBP7fe2tGvfZlegrIuTiuqTYhH+JpY0owrcqxmx0ajrqtn4znC0h
xWyIEr755c1vLjzFTRiAUanleJ4ibvm35Pgv1LmkBLFuqvAvrIj+at2HbAfNvjmn
2YVVyK6gN+dHA+CC2Slrh33o7p0H9luya/LXJ4SkDlNue2eypnMp7EdmIoc7c50u
KG9XX3YElVjZWndBUhMMnumMPxfuAABX1Sd0iCArJMNJkFuVtGV1QR7abE0FyL72
EA1GFvaDY2YiKs9SXDceFLLIEqV8GFqm2zNihBKFsplCj3F2naSop10caqexj2sE
MVpeP0O14S/nGZVJVX3JB04LBuRY8CiP710SnTwWdM0m/Ijz/21zuNpYZsFUS5zQ
Lnh0LVKA57Uw4k/YZi4EwONqCRVIXTYaSVH12uoFSQJvX8MF8cQGOeZE6cgEHBUn
r+zfCaWHgTBJ2IFkab43zmsaeP6W6h9KUO+jpiazdqM1BJHP5ix/h0tY6bd3bXK/
oZzD12Hds2azdjQ2d0/r2ya9rOCstbKuvhvNhPwT0KDFK6XpetIQhq4jUrrVozTm
vvfQR7GPt0l+ZK7mLmbVy2wdcpnewxyqn1vN4d9h2V904+MN2Swv6CvTTCoSxgHL
x/iU/iWtlldOhxQqVmvseH6a0PnwKS7kVtH/Fairo7h8/DzxghUHjsZ9HjBPPg6w
dOPWoZI+nFb+6/QIlq1McgEiwagLUb4ACORp/nCLCp/Vj+abeIBt9LN3bfFIUiN1
hZiW6UnrSM8NSjA6/kZt8snT2eZWGwpIKfZL6TedDIAYKMOCnPc3qqHmt4LqERqR
kMAj73DyZQVqqLnY+3UsLsdY9TLLURT5bInfhfaN+Cd6aPkMt+PYJkPBpYVt5QJw
68uXS0q9RZVlLXeOjF1pOTPlL0rTqRYqnNvUXhSoAt7AablWABkzeV5UEtIUN09N
otTojh+3VJcpbsjsX31VXIlbNmBTli0SMXhv5tJnC81v4dciPwZaKOt85uhKSp7L
vy/l3C+3ymR5xoT4W6J8OEUKhZopxY+nZ02+d1XtLOqinUO0RXFGlTHifuBqe+0H
LaGbl0Uc3TCB4zUMtm7gsSAuVHV0xa2ls2753oiDcRIv4jJ9ej3hUfC59UQ0OgUd
Ox5ydUgNEQymK/d4+8EuVG9IVHpp78RK1lRDSakyYBMJZ5HMYvJQSXoS2YN+PDkv
AE5pdZ4Y6Bz6zQ5J1KGDHxwWKVbTk7bczl8nHK3hXSL21acQYSPfpS1cTtDjsASy
kBuTJXA/nK6UttVkxYpkbEmmQEOFOqBZECjSlXn77+AKIoWHmEqJ5gHswaxelJH2
pEPWyEJzyJbA3Ug60+OD27RgocmjnCtDQ7TtyA52SRm2cW1EN4GKE+IzRzBCRKBR
KeVbdb12Oe5tZP+8Gd2M1s+pQ9Jtjed/wkDB2p0wQ7jcvzPM+F54O89XR3DBJhw8
VDOwHWU7jgMYTPr2Q9roS/uveqNr/vu9EFVUK66nmhAAPUxkkHOAtvIIpwuc1I9J
sayXkGubzZZqvyhyx6x9lnD75LUPMpwxFVRYTlWn8cDm+Xn7Vp70+SmsfY8OJEYc
FNPrFyq89Bif9uvkMRFkODrs7hNVpFdQRoDfdGnLtQGAR0yzDAOQLlyiBNVSOpfH
KurGtsVs5L1KsuexL7plUrRIqJiCJBZDi8AhUaYDNXY7pdKvJyqqCXQ2Ml303L2x
+PYVR6h5PXZxR7di/qoVSAAHDQCLcSRODFCzUeLJ43s5RuR+gQqp9cOyFAyoL7RW
qKJpng9btILy4GTjZTlYn/+7Ztk/9biOM6aKn8aqaQnO913g7+i2eJpFrpE/Lqof
NNfw7QZBqvMwYg4pKOTYhFkESxKcOFIcRoqGVqCBoql7BtiQj4Oic+W19gvLf/8Z
0nr3nkE/G5R0KeJlP2iAT1UxmyCb+sqFC1EzPpASRsd4VzriAto0g0jYyb6m0aDz
S2fKWZf1j8kv9icEnnU2ylpOHEcLqNnKLfyrpfBFjLt5E2/FESFEZGAnalwUnioW
xlOL9P6C2sqluJZvLsz/aLixouSm1EDCuXe0OaIx0tw8YQjmDvvDjfZd9hGzxQQA
c7uMgY88OY28lXoTLs5ZE6Y/3JcAznY0PjmWkLBmNWmXnKahSJxrISbs2GVWfaLD
DLTEoEgJ6qVVcYf67CuGBHyC23rdDYCgjWdCL5aL9nc16qve1YlxmRJtaSY7Ku33
gSdf5gNkc63jlndwWs1tcDcesDIrrCoqoOv08MElxdZEpIRFQHjZjxNQIMuDKQRP
DtBHO/UUWL/AmuhitzA4CVkGnDzpZqso9PyrDHkPPLSScOeWPDFN9n0N6ifH/Mrb
7+OsqDBX7Fj33MEq7a0LD5gqlnkymfYvfnx4L6HEe7ba4iDBuiJ5j0Io8gELFUwY
xJXO4pNd2w2eKGTQnYex+IWpZOpOwe/QDo7WBNrnZ2QDoXb2jaYd1d+H5/q7aZW6
4jC2EHBb/PvHUcgIe1fPx7t0Fncv9YCnCigkAOo4lXUFT9rg973pZeq+eev7a7Up
Y351Uc88JnRoPeJrAtkW1glRVHxBbOvt7BZrjtUohNOimW330Ci0CpYzCsdJRqiD
qHGvFuBYEk4yvNzGaLbX0PZwNz20SVbaWOFhJjsz9vV2ggngR4EDLgsq/EjbEbT5
cW4JBU8F7QH3KNcgwFd+lT3HoCSvAWuhc+gm2ts/EAl/5mhsSQTAhTqwxvnnEBl0
XAZmxCTu+3zEVGjp9/SOnTwr8YzrKUcUHnuGZ1CIFTI+WeGS5x0UKhUbNoizN0Pz
+jk1oN+nzsgKawxoQaaz7mbQHuZ/o0iXtd22QPaNWGNSKcpxCVdZwhfh8hGca7Vy
fKxJvDE/9A7vAb8x8K8DolNU0rzlRiEQ4/Fbng8/zNWd0gZqqxwZ02eSVQ0BzofK
dVw54Asziapgsp/pLEy5UKj+BTE6Ok5ekdgk44C5DKV4K0WTDC4alPuldonBVEEW
22DkSdMqtBehlYK8HlIiFUyzf/veW0BckilRYfUs19r/kKbKTYOKcs27xWxJSQFr
+EmSyUPKQJBJfWppTUQ2Gts6EevWOgNhmjqOT4ybhRXoZFWU9L2wA7Hi7i2iOAwn
F/0Z1Kd7kbl5xOSph7b+mKt2qtpqTYawRaSiL9XRqA57RIC2EPjp0zwNolX+kawb
ZGRPMCY1mzDWhkxp/np9cB9pY9ME63vZLShi2XkHwYvM3oGz4EzzAZBceeR5LpUp
Tetmqq6lWC4C8sIyqrreHyWnOzsAcgrMVg6TX4HFTGMHrtLP1XzteAj9UZLcLW6M
mD9mpWRtqfSwF2XUSpg6BvJfNym86PZffWfFUuep0RFguUudP5ntdlMCCi5SzuHf
GdmTjjbjiZrf5VcH0JgL2/J10pPKvkLwBgFiy/mP0WU1Vqu18DmKcY8ozRLMi/09
Puk79QrUgswE9rricU0j/bPC8dHoU7iASTmMlCPlVrJbdy8qD9nr11JcKt405cUY
841FKcdCyaZ4lGZW6tZaLch/8SSykOyABJJkTy9pKdHEcBu14bP8rHuppWvEJOkc
/yBeXhTXFr9f5UfiKf4lbkH5fubzWAecDqIW5yF96SHkRI8zmplR8jle9xEXSdy4
cApuVhCJYR8XliiO3NJR3yGmhopgjucxLimK53WRNgQ7SB7hangbh0PNcd22vO8U
X82yMMI+qpbGXPq2ISnNa13mrbGxwzVoVQoNWhfGfJP2U01pWBj+umQ8wMxIDgRO
vSgjt61oon3Z/SRUTLSO+94+QuNTdWslZfnsFEO3KoJkZIhCDuJU8VALAnkX9ATT
7nkfQA1ZrKrpuGmCxWkrGJY6qWvTZqeAKvXCm1TF2jOz1kfvlBsuhCoup/76VC4T
epEhXYl2Cp10QRLG5kNChnjeAf1RaM7NaVuWA2TgL6OmXw1BCkN0L78nLq9W8Pza
fT7ZF5W1csjXaswVwG8H5Pl0Y8gh/aWIx3V43SlE0BCJnH/dh3qXyoXezpDXbiMe
ANQYMYHTo1s/AkXMhfoD2X6MsDJsRbRahqFkRk14J5hz3CXUAhd5ezZ/2RYKPon7
o25PC0U6gloj9wjp1ckxH0Bhn4YNeFpCLMyLJvMLYT1y6Q/lLJs5+UEfzIVCaDfp
eESGri3UPRZ7nar55n1kT0jO85TYIm2zzu+jmWA+2PnG45OeYJ9qIiPE0+a9ZGT4
gYJjEzdanbMb+q6lpdM/A3c68k10+e8KwE+UkglftYZ4kBQYAZ3Fg6BCTbUaUnDf
++mHNYKDBqBcF3PCWiFCDj15lJ6TO8Dd063dhAJ1OTtY5JRJbSsX9FqvNZKpfAt6
bliLZzB5NgjmW1+AG68LarzMZ3IE9ApLJN4wPpPCUho8krKh7wZy9Ts00PluVXAI
lt0Ds+MNxRRWuPULCGJCwVdNT21ID2c9CoDmgHbSi3mWQYIMLYnEm2BAEWYUEGOp
B3StKOSUYca2Z/ctDroqzUa8hUqWGkgdNfBkHta//kEA3k9zvz1MjqqU59HO/NnR
8RbadhOhwdjscMosWZSNgs4lygk3Eo4+1tEkQVztq9o2A9YN7Bx4C3Gn3YOFUH1E
pQSRLiCGuB5G7tEs4Fycd7A8ysTL4graIS8U72wolcctiz35bXZTNCJxuJrpYXYp
hrtely6zfFU8VLv1uQ8Tn/Zr2gfG0YvaHCbXafeGU71JVn35AzPtE3r7tTdGWYET
RP/KTqM8UHKQbU1LSOzJk1rsndE/oURXZswoj8Y6XmFiu9NBuvUBPK2pz9vQUsCB
R+EfSIK296GFD0H+U59zQI+HZ4n49ZvYzKdKavczX6IjGCm4ItwBGC8UPn7eokrL
ZSzJrVrVUH4ENymqamJaVbxlt0BADfDb69MXCU358BYcwuqr0huNJGXryV2xuVHo
08JVThfO7Vx3K+aAYiTYo8q/4yaQ91RMDq2c4Erl3cT5f/SNqzHRoUhG1/SlwS0B
ECuZtzv4Yid6T3QftWn2M1uNZfLQu9qYW8+ZfRNyAbpGVZwA3Ffi9FJmaw5GrbcE
EXrlywPT1sdPm5jVNWBPGPvjpmkaR9Z7IB/96UtksSknOqSYXi5nHM64D0/VwRay
RGzcjEUfx8ioIU+6mUAvtLkV4LRwUPAYOWjD65mbNdd1gHfTF4xRzreh6omGh1hU
mXTz8TsVWbBGLtUS0LgKFPBNu8sNgzyw7nSeHkiXE9nLCarnWFn99DrsyGhfvVBo
gdKcQVpSu9gB0bitIUTkfeEXV6YWwsfHw0PsmIb5Ga1Cry1I7nWa0+T8tphi8qaP
/4LClZIeA/iz8AKXYMOxv9oHfp1Q/r6xFUFR9jvbO2dGothJzMtJQnQoFIrU6cT4
FylVIfrwhjVsVyNir5G7WwBva9ECAuTncl4lPi6fQX6SI0HqtWbUV3GqoVpF6vjF
s6nAHpLD6XhU4W4Czmt8YAIZ+TJsKySX8MCOXTJ5CD0o+kNYlteJOGkPj/IYv68g
Lv/fooo33uA772sJthOwpRZHfQ07AfTt8VhsBdWgPtgQPbgMhs2a9DvQ1zMv/vJM
w1ZABEtFz4J2R2qy2sNLlQ2QPmxxEQ+lV+ffNhd1ENZbCbxmoOpIfWAv1Fz6Ol4Y
vxMS8O/b4D17NMdRBESXLaahobqIHo/IA2zqvygB0WUnTUVrw4ODDuKu/VZtROqH
jAW4fH4t6fNOUAhQ1G1xouLSRj82gGrsgNkjRz4nvONizPEPV5+zz1kWxQP7rI7K
UkFgPvMl1/NfSd4CukZwkPeCMiDoEZJ6q9xg2jB9tGEPZ1HtZ2EQYDZHAVBroD1N
CCkLcvVc0j5hTeB6kFVuqWEmZYFKYKZis6jbl1wM6kRC8NG5gjUulEY6xpdDYhVP
hnMV7GqjUcE7eNxidLC7wRGaUxOJZPO4WnYNE5MfOtt2ISwqc5sHeWbGEuAClAgT
EkkA+fomJh3kmyVk8N0aIIB10TIxnXwA0DeZyEuTuhoJOE+UXKdN367jP+GIQT9o
QvhWC2DWyS1RRpLxRceXE23xDn75YFfpVbrNjICgtIo91caULAueNR+mCFBzDBxG
nC7FqRqowiBV4CQVJrlpf5nLFof3kZ5gzw3t3VVqPuAzg6+EseHwHfeYdhKo5pgb
9HAPcN4k8sjUF4P7Hfr7DikCqAJq7kDBQ9YQOHZIna0YOuqqTB89r3jdpqSn9dPm
pMJ4AKzClfA/Ad/sYVvuKJgwxEfcNObtBBmQoJHQP9uGGCO+r5ZKg3IiH+E++PvS
sLXYOvYqkQN1bGCdD0gdqCgtkcXucx0hFeTu4LxDi1q+3Qxgyzc+Td6jfkRXLVpk
1l8+hvvacalsjPsGuxatePryssAKpZ3C285LvVMGm0W6ZNlCcsGc2bh6uN7dTK6w
wNykMVoQA4IgKBFuRALpEl6rJRKyua0ttuAqeR5DEfjDQxI966jA1/EcQJ0RGKmK
Z7ujhCvdiUX9krf933rnFCjWqToDWATOiiPy00i95ghRY700VqIdBxTcfuc2mUfT
mE/7/gPFfDiouuV53O1/pT0e2w0vlXQof53HWzgIdqeX0kDKQ99AlyaIGFzShP+E
2SAA4yfiKOAftzlZNto5MeMh662xQEhNK2Vp7ZCspv6RcDg59HiyIPfEbr0gVi00
wnN1GO5XX9cYFsEGc0luzYbkBCEFlEXpQnweoLTAuIpWQNwYhFAHUaY1RYTU+xxj
P1F4iIRfygvYUa24zRyW+TbFUZeiHBTKXHyY/iDyq/bm6CsXi0b8wlCDslZx5hka
BCAuA2eGWX30ldhmQeC29vXr63URTgJmrlBJZumi/yZv1xLq+pU7aNWMEraJbimJ
e7ZkmIr3qKexgMo9iCyH03WtnaLu1xCcdoc9q4QQVVeCzVsNpSOywVnmDSyLzTbs
YS0SnIUefff6qAVbfr+xIGSpaKzsKCiwvxEr2xHIqjahOaoP6P8zeHaqIoF5VgP0
+O6UlHaZnkO6J2wCz9E7Yp0sbeJKb8awzd5EdcIG92eGy5N1VcFO/h3geG8SMTRu
bua1mzhcBDJldAycBa5KYAhGEk+Q/RW1buAEe2hG2CAIwMBlMpB4fIn1aT7CCDQ4
wFZhdJkloFq1eQkKwK6fld/Ip0ZrGm6ZQgpjhperhkgMqg4ilicnaC3rc/ILxWr2
NOHd897kpl0Hh4I7G1YvBr9Cl4TwB8EOA1JFKhjXYS/wnTn5PAf+cX/CWTacoODP
tJqPJh7JzSsEqjsjjIlaEZnSJCcS0hy4mFjAzkv3e5jwcBttln7ozrju8kB75793
Ji/8H3kzyGjYS1ubajuX3UpsZcl5zTauxdTJxYmZJmuAx/Jce8cdqqZUAq1kPCI3
ybWy3haJ8R6fggPo9lVtPEO/E2iiTatQbNt5BG+qlnSjEauIr705P7tErFMGtoSR
0PiTFKTBK+IhuR9kbnJOjbhNc2A2edTbxT4T3LyDaxpE7qCsfU5EAMDYXqFjRWYx
IPVHzc7lsLchVNI2G7+Oq7G7+eD1+B6UuzI/XlJwSWcSA9zXDkRU5kneH7KRxPtW
+wfaM0W64kcENyc0bNPqGdqVdcM79kt+NpH5E3W9WTsY40j/FUcBSR4JksLFwT6n
pP1oq+KYvG4WS7qJEb+/pTPqbtXUT4BDfHw5p+3bhFRXk9aCFbeI8jug3I/3JX3c
F3bshXdTDa6q6LPUskC1LWvl9ScSz+nZs3esMYFh+LlENZSpWhQNxAD2AshfaAFH
dXCl1cVOIsQUg6keR9cXpzDxpC7DTcDMY9kUJFcMvXylkFejL5Coox5zu5K4X+Qk
xzHn93sJSj22xMTeKyh3m4mmNwKJ0J2ue50uATO2p/N/mN7jUZENfbtZ0HGmo6zN
o+jztrcYvrusfOXAXuWxlZIyipNxJXRuaOqhgCPLaI26vVw3lufh1ZoRSYUMPv70
kS0UxCZbMvnqK1up89MhQ17y664T6uq5maMD1h9mhuwfy0E+ntiW+rrq4+DmG9Z9
R+00huO12Mb8VYLfy63wZeEAH9LFV++xro9YhLsMWFdpzxVfCNRC/uZ/dt/dFoZt
/96pDnZlKzDsx2D6twvRhLSftL8W6VpcnEfputhsVHEzRsCPR+4Tr+nSOSKlvwWx
YSEp9LOT0kdeI80PeuTOLVmCKCKV7TFkDb+n9HHpj/CQzc0+oy5kwIeLq6DptEsx
395jLbC//frU3j7jrTU6kiPTNoN7NodXV7iUiTDrvbK0BrbKYXsVl/WKQwhIfcdA
DLNc/qhg84pHTnW/j6N4EHNwTMVUbStnupVgEsIFn8eieKrTMZTvK2YgTXgBiFwb
j+BTmryNjDy5VKCTMBxddgpCG53RmScls0n1WXAsF69potk8wB5c9VWoP6mmJX1x
kwgq10+4gMe/9aofztVw5HN9591SFNUjOTDOsvHSglSoSUDs/0hK6p/YkgB/x99Y
wSodY+5qgJVoHy5WXqQ+yPP5tG/DFzHTjAIpJXXn4UzSGtQbn/S30A68YbVOA+cG
dY9V2/f4fQ6gViMvVOiOiKfhgWQGTKakG36xSHbyU0pESu2jJMhhtwxcEeH+RXmX
dQJI1vFlBPzWCxPTNCQj3FuMCM/1bxPkqpyiv/k8n7bvseJBjB4j81gjvRZKNcog
mAukd/CpaC2kqXgqbyU3Zl/4H+Rg6myLXY4aL1vQ3gfH2Aiz1b2l6CAWEVlWXE7S
yi1rUIY3VVOu8SUBGDAPR7zNBlKxwl0E18MH6zjZWAEen6Rz0I0Ux9xqkP3dwkVU
+7bNUsOfBUaUH+8QqX+Ngg8BuSBlECB2SWF8UGgpKmdOApvhgSVkQo4rcGup1aPX
mxAc7TEHq/H9rk7O4h7KyxLkUOPxZ8+5sUJ5bzNL5aLVsMX+ejwrr/zw+UEsC/Dq
JbNt8D+z2YP94qq5WaXujBo8+CZmP/KZJ1tvMOAcsoZ4S/N44uPU1TH0z37+Perb
DhpHDpmFxqrTVbnjnUEnYgzFjzC2IJiuHXkomf5/z44fiZ0KCRFylGuEfKPb3kFa
KaB6CCZlFOJu99fqEFaAtIZ98PBxYoBzHL/ya4nz2iRYGqBuzlMwjA/oUztUcs9J
nSPJk8lvbz7Z4xewyWIX0Mw6Otl1neWVD65aZ8UuiTwXH2lhPUg6l700UpEmUptq
KZAacm5Q9GQBNQAoVbVIdxqAvebyhzJFyq7R6BMOSv8/Z/TKz/PuwY2+SoPvE6kd
Dq0IfgwU0DrTG2ST9VnvMoHI7np17EXqtQrGwnCv181HZgGiFV/39HjfqFTZumsj
xWkHXiVK7Jjrn6y8hC7bGa1LmpUGQRUhz23QbupsD6PakPe7j/AUV4aM4HQ7gHDX
zW1QZ3XMLxFrHCwCBtwgs16n1T/0lD+D3f77AlQcAi8CmqU03FS7dCpoY4M5ff6X
+s8r/eqF69YA43N2AWbhCsOTHUM42gGguHK5x7shYEeGyKeHQOvcOb5Lh+NicTw+
BfZ+gF3gT0TxoVnSMLOxAZqQnoOkj0QtFYl+RljECqLmEiPIxdOAhGPX8Q6fWBAO
p2LrqdeUiyj9zu10nDM7vqCc/N1soTyMoQY3IjzTn5/9wt2ogrlFXg02TROXpT2G
HcNMeQ4jwWlH1FWQuEoHp3/5wNyBqhVQz90/7JIC999aSehpGCSzFclyjUCYsw/v
xEN4ve7bsjS6YZY+NGaPUaaR60ps3vHZjdW3zzn6mPqFUz0pzZn093w5RTOY2gnV
R3/57OfrUV5neUmod2L2ym/NFLzpWjwcx7tK8VBXAFtOIaYGv5u9UePOr/JzmTF/
hWrfagu0AsTMvPW08fb/Wt6x47D2u1If27f9fwXjZc2Mz2PGlR74Liy6tjPzaugm
ylv+DHYsF2hryXRzlUIpBUr8jJiOomZzfVmukL1KjYb38qYTvY9nja2+rR7p4Ynx
rpHQa0EuZNMj+061uPjlqet7UI/jdlQdoYC0ahxDiT0VFZ58xmXxQNQFi8rbvTS6
BdIaW1S0R/5wTeB3hSCSGXE80gW7ZtnonP7I7Q41dIBAwr1IY5Q0FsjXPDFmcEVD
2jUeKdv5EDTD9XCE4RgBpY3uWLytTtsbJg2v42rBVHCDIpX95d2k+XkCBZOjPhPG
vj//Z8p+yF4n82bj/vm/uJc06n71lW3hM2pO7KPVAhUJHVjHaKcJVuwxY8LuWeTl
hwVBp/w2lO4sCVCCJwG0hNQmtMQx9B1owzH6FdWwx3gDfEazHgzLHS+jyIN5MhDc
byAJOmf07wefN5KLaf/uZWZQJPIo9puo5PuidX1gyP8fRE8S6WkgxeQfM55LMCpN
JmwlD21CEOgFZO1UAljKeigPNTLA2jiEwoj5dDrWUEJYlEVqx00T0isO8Spbwz2X
t2mQGYDAOWLYEQxl12WsmiC6K49cnj9HqzzPTX6U4VKwnV2+c2Oo4yFLGDSflC6X
VijKIvRLdheR+MU5Ktq78VjSvCJLcn0sQsDt7l8ZVup1JRIeix4wZjYtsOoh+dCr
s+3nF7t/lhH3qM/0eAUJxnkxdXunpDfjZTPGj1Tv9nuOwififDtvhmzt327dzjm1
JDSJpaAnoftKlGvzcIkJQsZ9Vnw945J2nuuHoOX9BzoeQZESAwBdJoXewJA3VDB1
BdcHUZ+yX0WSGSUfd5NoVakLh8BTd8/R2HiONTytldY+3vV+Tab+cwQ0cDzM7JcJ
Nv3AXnB6LDEGHjrq+qu7YxYo0AApyxEJhGfGC9OC6ZYIvmE/tt3wtfnWlOkPSQes
Z85s1SeVv7iKB1NouwkD5ndLyjwf88R6kScdfGXR15nHxeGozABY0e+N7ucpi9sf
aNMtU14IJmrR+Ny5ClcFZ2P0lYYan7E/leh/2OVGjEtapHezRXqGzO848CRBZ6gQ
TRq1OBoevm/04ysSV/zVoRX5QzwudM3+t3tB5CGMRWPDN9YH5STW55+1syat6ePO
pspe5uiB4pya9CkyZVAG0VyF6buKEu/0noo0IOlJ07R6+60/i5bVMkxOaxdtbvHG
/bj+8LVpXFKtWofcQnNM+EEzkPQmwBOitmykGyd30ndX0bFCunq2fzvWFi2gIiTQ
Yzhe436gDhEBt9uIuhdis3oSOSvsW18yrOLKmpQ7AdVWvF2WietfW/SSmFBuPm1O
fHpX4BbeTO8+hVO/yryZ1GNrLTfLa8xsyaF5Bme38IZXt7BpoiSjmxo1U72ue35/
VktcNIxlH7WVxPq/5d/yOyQZbbFbOaHjfpdZUTPzEHnTwYKW8n/0m2jJHhZ2Hb1A
/yH2OFZPgoSLhgSJeBIr9xQ4+AMMnYlQ3iYEFZC7seyhlLf/U31fas7GQNjoQoaI
nytgWOPn21yYUwHX6rFNSSPqsq/D7rf5IPIVA6DwOt+D2G/pkIwlnYSjj9VeTXCA
DVyXvt39ocbppXhtnNU+SJSOPPHDCgl2fKJ3sSPiNP2uc3sC6HRuJ0X+vaggzNQ+
sa3FLLATWjH4P91DKa8cBo7z5ARiimz/z7ujEG52vAO6ZUZAo65dFNCwIAYRMqxq
KKmw+u0vL/64XFcO8JX3T/JH94jv5QrYuvi0P08dgrJE5l9hVkHGwYaKlr7VfdOd
vTOk1EgsxqzHb3TCtOSbezB2DPDGZtNUDU6ptf0ARF+BkBmv1wNGATTzPVE3sDNU
r5QV1MG9O24+uy5k+Sj5khhmCBIGKCPg+/tiQ2ywDgCiSBFqs0G0CHTP4+TLK8O4
lEh3YQxBR3mgm7GwffZex7ik6k0u0Uf0JoTOSDdneb9Z9y8imBWVUEebzKt9HhQm
yuJEJi7wykGWLM1Wp0C2jV+IK3MtsUNi4daUVC0r74CMMdiHDlu1UCCsnVU2Fr16
oKEHEAzZ3AAq9C6VjcM1z1uJtd/SIhRIfoMq11DNjLf3sDxIxbLGiIGkpK5tByax
Y5u6xmCb+8w4l+SCuFbHpEVppAundxXNCj/ahoobCF3S9PVY8KxWMwjk1LnP8b1B
JH6Xfhi4VWfyV+XMBnWwYCUzSOzpfsOhF0a4oQBEZCzAKTR7+ULaXbN3D7zKGdfM
7ccj1fe2n1Z4NbWRT0vGBDGQnRWvVojBBw1W4wXVkP7D1gfI4v0jRZ6Bib+/Qbrr
7N3RVjxgO8MOOTaZlScufqNo/fOF5m1+h+kkVhYhJgNdnXBDbrB7hBwM0OTGhypy
d0H2UwC/vFg5Fh9rFaTfBqkbEZsXiUXd5DIIEXhwHfs8c6wDjWQYOiMV+9jnBTOO
eIhlJ2ZxbURJQU2E0pjJ3Jw6PLYu4eE0QIIYVTTfWZNswcBNBj2MovSbcfBDYfT9
3++XBdrInVzY/QB8/h8wGRvTCW8H84eGaPgmL2L4dYSRGwN0LrSVtOQAwTcdGxAO
vbFZg1oBuYxH5LwOWrXtNXf0smeoIm9mfz7tPJUMzB4oxTmqEZDv5P8r5dgzi95N
zRGcdiFkpahobAS/MzUJEfJFpYlTdof7LNg3lzRUWU2kAGO1dFTOD7KiAOQ1PfF1
OqeetWolb/nkAmE5qlCkO9A/Jxa4exdUMTz7/cD0fwb3y6QHXL7FbPmF6Jq3p9aj
QUnc6kZGJrSljshHbhFMwbrRI7psBLko9FxBJmgbzYdfyH3zeRzjmkuJORoVCP/C
v9oaMc6ZTqUY51+mbJ4eD1jXvPUMwymEcM1yuv9LE1d4okQOjaw81yEFLKkHCZmr
hjKHmWN/pkUm9z1OsT0E63/vJIPDJrvVCOZ383tS6jbdJBSZePQbwFzE4MfKbLd+
VcDJRq/+eRw+dt91v6VrfxbSAX+UmLnin9scpK0LIAgcE555DtMfN93ypp5SCJ5q
8kc1jvr+HNL4Obm1O/Kv5ryps3wHHOPvPtTk8K0Tsh1ALVSit8ArzzEia7A5yYUy
znooIOmEhNq++HWt7kTmx6HvF/AnGXR3M9RBc/zExE3mbAM2miSPZnIOijz4l6P9
OKlGOXa1+Vu5jGz2oyad4/07I3oAwyAM3bIZpD0XD833C12eQ2KBKabA9ddWZ5Ad
5oglhiqY9dTtXH7gPimkPWrtkfMJrzJx0NJ2HJ8B+kkVYKNOj2FkUXt1ZA55kC/U
lZYTV0QlctFvdN/5vVfw2j/TlerWub2025ykeNZEjrh2Zo6Zp+IYvthNARZ210M+
z2l6LbKweY1f1hYGpqqQmLn+gtFYPkx5BcCEXuyeVIIo95lxyPdrh+U0vlObmm1a
EyH9rJi+C4v12UxCDmJlN/NQJCII/LUvc19wtKtXryydYL3IYIZfGdrMQhpotLY4
JzuBDJ8OR7Hem/ujoOVEheVOVdL/Ih6hihC838gMhOOpna2Ll+VefmTEjLsyFRrY
jPXENQ+x4tjVs9AwhNXlcejkjy2wqExHI+zoXxnQcN5hPSEMobB08Bgo6yLP+6p8
o2XFpayY/HAHR7YECq9YFjH3mbP61pMPWsAoLdm77o5r7eg0lDQgZ9xQgaZLagC/
Af/moHUD6EGhV9WdDefW62a3hGd8WfkQjMOG96/tiqMEJOK1gduCebH+0XAUS9zv
WbOHRImk78rjUt2YIOnOt18Xoa/0HM8i8yYraJlt+auYExRZu/kcHDXHV7hhd7M7
o1ni7gxHsrLy7+rrRY67ygHxN5aIJ0Sc9XrZoGlkwjDErRPZPUdvJKd08Q9/60Fj
oVVdizL3qGxSVnZZlggFkYnAW1VZysXEBSckPhyJ/jgdGQIfbAfH0Zly+0SSRuO9
vCd3gKn2KwkkIK07HvSgZBAs/RU+4jNkqq+qSm3rBa48SXfmTaBbn8Tme9nsJv87
KlZu5bJEmPaX29thFQIV49spLT5Xdr0n55Jvny32ivWhh0P7bkAtLlDLuqBOPpVw
wBbucSc85AzpGMFBLnbgR1LGWIXYfP+Ti0wbDTKoMawTKD7/4j+cCjie96CDlsl7
T5wMU9nQGuP9EZPRuu8puuhE2RCi6Vg4EAYbHaDqBwBiXScAF7/ax+LvQvY95mdY
UaqbAewDLsNAcyYIAi9tveVa0NAWQFNt5Ud4Zm9g36dIqW9CVSSlKlO1E/XFYWI4
IVmMhFauxD+5zlcGVKDK43a0CRRdqRepFXtKA0beXiNql8ubEahy2z/zbV/kMxCQ
6hM4Lqu8tP+ToU/6YZqDx61A5C/LWGXrLiuWCXga7ULVvBEnd5vMXqZwBjvkCuk/
xZCZ0OkiCt8cXD6B5Gaul1O8fpWNZ+B9EF5uo+n5fBeSEWsmLmGLvyd4akiKYwwl
U8b1KKvGVXW4cgK/0Ka6t+yEh66bAka+TeOCz2LKeRIZH60YQne7bfp70HEsy2Bu
1TJAMGjev7WLJaWCVIWE6G+kHebnNP+aHxNJaXQy6Ywt8HZ3Yqsqx4QVPpp8DiLl
+o4JER3u12tesD6uAX52EDnwal6egt0EheZnyZ1wYsyhEnDdFlyaoijoDeAyw7lG
idmYUfqomyqWoviXuTd7bGqym2vOUHSq0ELRF/8ea7zc0xpSrduVW2GDLj8hGCAv
0hl2tZdyWrivtiyfhHJi+8qv0Dha9HHW/RkQwR6Ut4fLCbNoNwzAvP1xVtLVV1rY
CICfzeLITOEFPkUa6nFEr/fY/wFld+x5yR74vqEixESYP575nI13nHCwtsWQapaQ
iExxJkVBN4k/ykTwMsv5yFVL4W+QP1lkhxfT9sCtPxfDhE6qF4dTsPES8dC69a2I
x85jUibzq7qWaGZzvDcW2IVqGyP75W9Gw42hwDHxK1NtPLmSqrSpGWsD0fxKJXlG
g23VXnIrq2nQLKml1QaEDoEGx+esHnRxB9vguxGP8UpCqc+1HmKOGIraYKUlpWVe
YUNsN5GUdwdQJfufmB2iAT2fPoPjg6Ab59V33n31eQPLSydpBTQb/HsNRNerOGJn
Q5t8g9oRSq8v8LtE89NpJ36Ikn5F0Z6VgRfBBB4+h9I6yCot2FcKiI5/fueZRYsT
1j1A2xaIkpJAVZUosbNCJVKx7hF9gM0l4FWDrdbH03in9m9LzouLOy75lPyfvrev
PtVZciH1R4+BAvzoVjyueBbElVURTtyknvqq9v7KymMh+EfZQ/sEGpFA89PAm2ny
o50a+AOV+KViGYAbC0O43QHk5cxee47Vx7ek6rhZ8afd+MSL/xd0tiSfaVHGnRCh
d2fb2cniC/vZLzFFXnVALFaI8SOcaDNyhVmPFK6wTlqLKsO6DcybBI01/ywoclp5
Bfjd2n98PAzuQmSpNVPukf8NDejzCXEDzrBXBVrXrHZHL2Z1XieS/x1LN0P1uY6w
mLvitKwxKyJJu8MA73SEu9aiRtV79BtLmjPQUHDmPWKVOU9rHw5HoAtv5+Ok3u5A
YQtVf3S0nEeeGSODb67MbwQ08XESURdTF57zPTVYfdwOOPSCQ5iofsX+AHKXNDpE
0UI+VROf/hI/JWjpqUzra+VYFlm06v7YyEadrcnSSQs7NKdcLFuKGyZfqO9gF7FU
38dt2Ed48G0lisO9224lhQJWbjs0lZqCJOLrjwVfhj3fvi5XMZnUmPGAEuMmH+El
vUZE+roYI1P6/Yf759PUVMmTFTgmvdNgKw1bsvXVUH9WWdDgV8IQ/fdzCEm//4cw
eg6/JDBMe50v/bRoKXBZD/yWAIS4X92x7cPJrQq9VaxlIJf3Wh3wW0OB1kQ+xn2Q
dOFHCbeAOfEVIVJ+sFh3fLmLJGAWlMfp+dwIuqALqlmUXPzZC2/L/eabzHyNSBV4
E5UVsGfVXp1/p+WjzPbqX8kyG4kZqFdLs655NgYZWVrIf0uYD4gC2vhvgXi4fuib
Gc0LObFgbdSLmpefC1hothIgYiICg11LEgtBGTCODbThQt8nv8+k3mAqct+kIaWk
V4PM2sZn+zUN2p5gR/wBMAU8apQKd7hlHKFUTUceCPt69X4KnQEKni20uZGm1A+P
lsq3rwiDmTRNZa6Ha1UEz37g32R5x6c4y4q8C8wFDVCIRFycxbnQM/FWmplLlvF4
4Xr7/sz4TEmF1ifkSGZHetypDz01NlXh+22Pv/CCAGOcpAK8/0aGDl4kKY3XruAB
lP6hlQP5362cW5RPiD9qAIAsm7DOge/lpppv4N/bFLnrrCzgB9PlPWXnExS73mz3
F3d7llB2CqiiiOlrRt5/RrQRnNNBKViaSGRRcfvOqjI8ulrl9M62V36ia/3tJNg6
BIRvm2k7JDi+Q8Yuc9uhWE4qyWav0ta4rP/VO413ysXjVOe1VbgAxUJbIz6gk67h
HqZ/7LnY4Hyb/BI2iZurYZ+WIFPfuuga0TrxR19XYojJjA/N7uWdHgwiZKvwKLeU
NMJJMEKT3vCZVxlOS1gtX3lHhFZZ5dB6gHpRL7wHXUt5X5cvH8oScQ8JedNa7Ids
hAzJEPMzg6QhtoVdhk2b+cJ6AYwY6eAjm95WOyNuxiSpY4KUxQKGAmNdUtmRJUQI
GhsC3HW82q+RzCNZWoiyX20YHbS6BZkjIikTTKbC67PXP4psJimCHoQ0mogkr3ka
lQZ9Zw4pbcy/lz86ugaZ2355S4vsW+noLLkhmpgCl/0nu2bPNLbcDoBA//1f1apA
q/zB37b7zHKtbOiNh4Jsctgx2L+lNQekG+6iVMLev5US3Qc/tV7jMIMDb6sG/Kme
QdK6CCEXfNkCjHl5DfANAr1Q33diwHcuxz534/6Z6syEUVarNLcnyCrLAY/uxGkd
Nugg/uWJDHc5ZinHHyPNNaJZVV8DCmcnGKLuq7/FLm2TwUvbFqBVukwVK74rDFVI
YhX6kY4RRBDK9QLWvifUvNZLkDI+oTq5sUPnX3xOXezu6x5Djb8TtYPmQVGVGGos
mno+5OgkirBYZaIIprSkjueu//AHzULwyZHQSzOvlmtJoe7aYsRnZEFzYc6z6cCr
/jW2WIOhZ1zO1lwhb0Cjp73Fbx5YaXDPcHA7hhtiu2tt5iJlGt0XWmxUvo7UlSrw
6yMe7n0bYGZMb+bKP4pJ12fVsHoGHzpWr5Lc2+oPf1dUuR3IbDfI/W93LLWkm1uo
hYP8i6g0lmouycc22wonveWXvJXqw+DZBiIQY3t/sqEA+KWsDzfdMI7Vm9q5EC5s
daS3EPM2+wKY8pIDo3O/wN3FcYaB1oiTVZZsiD7sqv1c15PF7T9+DKgEfBt4a7mQ
7inx0Cizr4OgaFuBTJ5E6zuJQJ8QwXxeD6y4dnlx+aAc0jabGaru//k1FyYG9ip5
ZIguJ2KFiWSjWhTPHPR7qZJxTUZlFMqNmGD7J4M5DWhrDeFQeurUQozLzAIK7CCX
JPAJl5R7c84egtf8ZICCM4dQq8ben8ldl563jO831wtkOE+xZHBTdhXQyzLQObqV
Qin0B8rR7wFnxYEhRk47HbkAsvzg/dYVQBzOxjBdonSEQWaGiTPKyGF1jAo9lX9g
JatOyk/bjPKiIJHXYplDAC8wHe2vMRTmrLPkOmjgS6WDjPohcrvQcwzFJzQvUEVO
cqGXfc8H6ud3b5tDL/BdmAQQi6Q0MX8BW5U1BWfgrl0zlNQX41OJVnNM1r1MENlY
OMbdtd9CbNl4SXUG0z/A1GIbPUgOdeeE9kk7bXwUwCe1iEioz9k8NA/LYMS+SiCy
vf1Gg7CeMrCQJ/lOVpbvs64EQgr7VmJsMCsOWzI9RFaINkAqYHl7SjIkHUXCfPX2
gczIo27pA5qTMGkPkew7N/zOHVCXNhyztkBC6+XL4a4W6EZcn951E2ZnG/2w0yu/
aY0XaaWGW/dXfQWPILuBZ/lIdORIgSEnYLPZA2evWdB5XizlK4SNw2DLF2XzoxwI
BYJcophbrZOgDOVAxcxS+ExYj4WxHjUw7/C+PgW6eLtKb12Fv/JG8efLBCN479Q8
XSqVE9evIEVEq/jawYRfQKTwWcRVWNlJeE46GpUbfUCTF0JhF7m96FtiQVHxD+IM
43FDVN5O7ikEUk5PIShVpUQE0IEHLGulFPZh9yjJYZSi0zSoh09FoWEjKNHcKCtM
/GXsL1x9FR5qW99jQ0YA668vlLhTfsww4Wdq46Yruv+7GpAPcxcKbi9SrlcBiFuh
9AM1D+RrIQPyv4Dq2Jgoy6zufuiVhsqHCkRXCDiVey2DpjVYLB/790lXm2pnZNrI
z7gwpLQliWAujFmx2cc31+t0cgHFl5/Ui5VdRwCXd1Cda1FL+odmugKxbOLevjD7
W1xkYDDwOEvjcDZGHUr2eVNOW+WUf+7dozgFP4TbVFoGyVRlAkQpVT9NTqoVUaPM
hmuXuRgTlsqCIsx0pUMKSVwGbhV8ZTeP5i/Q8tZHql3f7UYMm7bRLNg+dAhDrU9w
URW0/4Wh+tLHuJhwZgmMpcAQcYBSDtqpfdkiImPNPbmXTO7GOJzI5N+gaXWdwzvX
HYg8FU6h9D0nvb2iKn3iVJE7VopBGw8klqtjVEsiku0E0XWPZzVhRomm02YSH96r
qjTdG0i/TFbufQlXaPXZEgliy02AkTyKJd8lKeQcJFfJLmCywa8jiX7NKUnxN/ly
2oIxuCn9iiYIEonz8KeMNMXRnXGgREK5OsmgkHrKSLWLs4O4fkjI0mQpCOjx/ii9
U1K+IthoqjFzzMucMFSPMAro1RmMiVNZmHJFjIrWIPq/+vldaqrjB139NFzO0g8g
BOilBgXZq4lp+e08UccCyYqDN0SOsAR3dwRCGX92hLADFGS7XSAwm3p+HNu2SGl7
zjPM4z7us6ayX+BMD7zUg8qqO4DlmURuJCanWkx/ou45UsBFr80Rioo9Q5aYiGKl
F1f9FC7mgNox8veavMUuZGtHNOgSLf0fUu0JDsPBKAwIVeqeFZOvqXW+J07RQ152
Yu1xoGK8jRKE+FnLnpJegUHSxGIB6ZiiAoklVi00r3TpVTNUaaGEbRqaQYaftmFl
fws5YdpzKyi48l6szHDeWczdsmpYg2XAWXWbEJGmcThnZ2ukuEsXjyqMEC+AMC5y
gC/UST0XC4QYSFC5tbBUuNA9kyDK79gxOTiACIiRE4/zeFQFXeNPQSSb7ImeIM0J
tCZ/PI/zpm8HOmFCESXw+jH8zdheb2iIuKLA7GXWfKoX6NfogZfhf37xjahzcHHW
EjTP6cWj/xeLE/92m7FSty1UaQMYy5/EY7AzeHDpsAhgiHDJ9H4svY/9Z+PQEvuQ
lFaNinFuBvSKidXVIrudUBv0VRIXBy0JaHD/eSqs9P9iLk9a8ZALeaezkLmVx7Fy
Hbykr0nRk++jK15SIJRbMWNXfRGDqfRYqTwA2YSt+PsazhrlYtVvonztXud5H8oV
U9t29iRDO4MET0MAbDF6sAx6GDJNO1vnRl+dq7JtzgccBpBcNc502U0yZRbyvZ6D
Eepu+VXaFAL3SvhtI1P74ZwMn0ltkuACQaFiJwGYBtma/CP7lUJTUMvcsmsbFvJT
Ty1fjLWc+JLQhg6Mb3fn3eRBw1XBFJ15MNU2ckavl7KzTL7Yofw9snnhURb+SGno
C1cksP97dYbTPNJ3Hjdx8Kwd34V2/aH4ytB8PL7eIgxRFybWxAOztGctZ2ygjRVy
oTne0Zs+zsj9f7501wNeIzM2tS8L+gYPCevj1jKM7nIZLAu7SqMFtO6IIRDEAnAW
/AIhfyH4Qyb6HzLr4t9hMC+wyz59dcXtwIxys0zZkPbyRJMIiyMNM3309ZnFtkdr
0YoCSZwfhrlNKrrGfSZZDKoABGF3zbFi1my4Qcr+QrFrr4L2NFpc84ABINwRR/RL
9oqNxwP5Y/GPpzP226w7jA5AGeA+EthWWnf+SDTWjXx0rOtDnh1qpvb2jYl6dbXw
+EzadPYVa8rdvWtNW4ji2sfgzLElbuAJqPZojAVPPRCeIQDChuScB2PaUeV2cfsi
MxLsuZhlYyYzqHkKAcWoIhjvqIaUk1fFvJMc2riRfMKaI6Uwtn1qJoOH+UkGWVjD
sZUbONLlVv8e6a8WE5hLijFXJkUCzC8MQ6r/1j/P5kN9ML273aHEI4UkbocOiZFN
xQoY3bE1CHz2KGcST51yBlIsofXeKQLY5XuIs7UnPqyQDX2CV32rI8MEIFEa0owh
rMk2Bfq6XR7sSVY4YzQfz3WPMlW8so8EBBzQHcaQEVN5LSq4+x+TioHkIF16RueH
ZAVY+1foAZQB/paRtvmsUHsj6RbdoldbAp0xJbhzIM5Al0miuK4AGomxMyzUZOcc
7WH5dez1AWBSmk9MJvC6XnV9kcmUM4q0RQ0Ndra/5d4v5gZpMAmnaUwzbSpQCh7K
OEUkKdJhmkPFk//vk100vmnCZAsSKrPMYgPUWuDJ6QOQrxODYwLoITTZGbdqNZfQ
Bqvzdq7TIJIwLAJADEMIQp3gECAGqcakbhvg+pQg1FIDVC4jLXBY3adXYPqcgQJC
C9hH03a5j4fvaAVDpJkGG79XzVBMyfCQOD9o28IP+yYPNRorVaiAAdgdKlCdXY/V
+3GSPs4wqe4bo4EquTHo7i+rfqjUOdBKx13pCCSCGrMmnCwElNSEAA+okoQhr8y5
8/SM37NMI3srPcPhBg6WnXTNE0J1aRQRZxn/DIlzmx6o8GAi2HLXTgRvpSXo3LXP
vPVKjEqJ3iBUoB1205/A0DiFUaO8nSiFOegemdMt5oO90p7PlAomPR6UAZKowos3
kNyGPqpUwfuQaoGsmIbc7fQ8Z9x0vvw02aCFH0z3W0+LjRw3d0ecGEE9LuID5Cqm
QXKvA385KQOo4UNP5vRIg36yO2EtRF5QcfOiSNpWKXSbBMa/VjrIUbCXim1OCBR4
R0mkKPyzo6Wa9uQJamLmhHT7ZvqDQDAmxrxybAQOZYfzrDqLHN/+v7/NOGjf3h9Z
Fws4waLZe5+sE0Q0mF6XXnxV5NiO/2rJC1zanFtDR5D8MVujKhY74tp9XxwieBEw
xlIDCt2cOU8gpJpdys6GLSaPncxC+ozQThZjTV35vldeCQIXt6iZWwZLE15vCat1
eNu5c48c+MTUYj8AyJRvB+4Vyr48o9b2cJyUbPgPhP7ok4L+jkwszQih48ieV3CE
1yus33QnlijqdxNieewS5hsPye7ksgFZOxfY7h68NKyOsuwvrt6L4eMn8uAVdzm+
7l7v0QWbAO1XvFW/+AdndPrbEDXLFPMtkaEPPdsQQ8TXzn2+1Be0KKFLqd3CWfK0
MXJvqXVe4UdkH+SdVFFd8zWE0qNkjMwg46gc64H3UD0HiuDmHOUb16RccbP3Cv99
mjgBbnhkNY2zY6u7gAQ+INxk/zvL0mPwPtRtIdQBm5W0I24ZElpM771HpwpGiTE0
HJv5NGCldKUrFZd/qdaw39Kis0zY2EBNswj13igLCtDw6BxVECMDn49fT77k1R1+
kjMRoiqWdkPRSQu0WgjvlSGdTb7e9WW+WKI4nEyy5DW3jh4zhMtByjDppprTQTE4
OUdfDpXRfprRqDFntTWnGiGySfu1WbuKac8Onptd1JMYymTUbIlOIHCCsjBFuEth
o7oCzN6ZS3s9tzAYVsBP5fSAAKQtjqFa12JjJj75J4lPZJ31szOnJEoeJJWbU6v0
N+PtHGp6ceOPF4R9RmXpntvKi9pZ7J+OxERkR4a/lRyw00HYCXYXSqP/Ax1ys21A
9prS2P6/PwxE/zv2YcWW3h/N7YXdlgsDAkm0JTvPwGFE3bBbIEI/ngFDcUXwazGA
vh10TGcm5SN7nvYPihQY0Im57rsOBbljZjDwxDoKq2DTN37T/KSCzFdKgz605SRk
4+zE+AcTxYPxugDBZRNnkNaB1e9VPh/KGJ7oRO7fc0/a7Jyddsd0nuocW18+inK/
UlbxesdOg8B+1fFkHhfBS/BfJuRudfB4jOSWtdyOcnf7tzO4xvkJJ6hpERgccV01
EcsG6II8mEWa93ghDN5r4BBTh1iH9w9XUVLItATw3sgxipers5d6KP+pwXJ/b2EA
8PykjOqQtlGPEv8BRRxGy3RNggoe5BZkiO0EBKpOdIiyQ37lDtcf7/en8Lf9Dolx
CZilayw4C0Dtw7+5AxrBX/lH4AYjCIoNJQ/00TSphJwRttr5CF/0PB4YJpastdyI
tmVKQ2+0Hovfo/Nt9+4Doc3sXeuPB/DaSOgMHqtW3wOt4wriUTk8hXU8m/3Ys48e
Q1p56fnsf1SSxOh+A4Wb7dRVG31W5AwTbf5BWSMAeFgRExvdNmYeHo6z5keO77oi
L9joJfIKDkL0DKLy29Pd8y0uT3xdgGvP+LVz99RvboKzPamGazKJ0URn7of+KEqi
j2W5lxtIOjO3u9Sn22TpSi/+kdH8kgN959aWjwqHTe7BdW7YDsSU6SY5lGYVyPys
vJ3i1lnb76qSP9h29YAC+W9pTnE4c2da02RCntoL5D9SNhtG9ZbckqqmQU/F8G3Q
CZf0QLGXSm/ecCE8RvUmouJsmzwYIviese6I9z7MMBbzNM2v2Q80KDGdFr/Ee5Bf
d5MnzVwmVe2jOw7TIqWrkzkB1CfLRPEQdqekl1LSvG05bLVWyylcgaeLaKlsnbKx
Qo6TeH2z87iLuubVCkKz5/PLmkKdaBSYeUliqtf1xFFWFuW+LMTxCVGe/JdpNjA+
ZqRZ1q/Slnjk8BG3uTia5okWFoW6nqMhpx+fmSB6j2kh4QHg2OvVANRYgowF+uj/
8ueamkjAEvjRvehir5x6jREQMmsSfnEsK1iW4ireFdMuJi+lLjFIz5sNYwZry3KY
OQ0ix8wpKi1ECoTVp2kdHk5mTvizD3XHSPoRvqQiK13BEI9iHJjJSgThxVvsLsfR
Em3lkVZTN3KUqsrfcMOa5V1hNxlOuqVQ03+1/VSYmwzpbHQDKvNFmRi/R/yUnIG5
0z/2b+ankbq3ijZevMWkeehGyd4lC81QdUCM/1OS0ARkoByZYUw/1sIMSScg6yWt
6h9vhkraVZ4fqm1RA+Q9t6VHM6fUaWq21UseXxc5G74n2KW3uqHQxkCLC94l5Co4
4t5hDPabaJLPcN6+zMWKukGQabB+SHBcjdcoECE+UPxrybN9DbR0tzaitp6TqI41
krWBe0qAtmgXq+nn7JxUFyUgc7QB4rqcaU+laoMx4moQ2UOXWnX19I8MpdAKRYzZ
ssI3oosqVHdKfse7WZ8PvVB7z6c/m/Af1oildV57/pHZ6SNke0d7XUeRKBufiJJ9
JYt3DLpuTLt6n0tEhEWR/wJVpET6XJZS3JJkDqFMCQ9bg7GKVLMYP2qCPzpKL8Iy
6s/VZBy/pVgFkgEpi6Bn7ny8oI1pbnjrmdebt16NewvXToK6rh5ci9CmefPeEtU7
iK2n6M6nrKOT0EMC4xAJ9PqyoV+9Xvl5m/JgGzwO75HNk8jrkVpcJezhz6dnFsaG
3Jh6j9WxbNtJf4RaJOwWKEDSI3paQgj4jaE8z6WIBUpsmOeuF88V8GBhfORMpnAp
cU+J+m1pVhyI6pqp2yEUXMMqLyR+P2SeyjGxTpESRI7aLicHjhpIAPdNVqocbSEr
YTtpqRJ47GcAay8TvvgK/bIRWOQWQ/QKg6GmKk6auR+lx+54oJ3NRxxH/Oh3DNyS
Mu1NdYgmtU2Np6mDfTvietTn7TvtPrHGab32I891H/MVXo52Hsser3PYKd6ksTWF
gexAn/AWa8wKyelpuN1nXqZ57BajT175CuH8sBvb7WOJ6kS0Ru1XRG3pC6o2FAeU
Il17fTJzBhNyPRPZJHfvpj/fgQBI+N0jLHGbBVjnIfZe6bMJ3a4SNCsexgWiFgbQ
8qKYyojhl6QOQc6sdEpYwwcq8eYnsP3uZWewvI4WK5TUQ+AJvv5a2efGGBkRSXJj
l/QNUUeyvFx41uETyImMhUj3u/ZH2mFuIDAfDFthi3Zkc5ln7l90DICGAUlNeYhj
RAODZfeYgIFL8cT4k+SLuEzbq+0RMJm/jPh51eOueuxi3wYNqyc2x14sW3P666qt
zgtNpFDzEsKmW5m/aW3f1+C+IeGq/JTvxYd5NOcVutLq+hJclEnN5zQVpjx4moRL
N8Dw6Z1F5Yf98MEixN2pPicSEDalI1CnG6PdU4+YjQVqTwAG/3k6GK0WWeQz2XnY
lAUeSuP8UX/KRjJ+BelFMQ5/mT4EFxu3q59hZ9AZmBAZAkTF83qEOjCjzSaP4DaH
AfRIkthu1SQUxRQPham5xxJ12fi2pcXUYocTASGfR7mVOyQM/Y2ps8FUWEndvP12
dbv/HGQaeIb1RBFD7mfGcFPwP0wIADVJ1COgz0L5ntQwYldGzbQoisuq9xAzr55A
9k4zRKTmt+lrW5DD60gtP9BY0Y1EZNPAeLUSjMsETKB6AlgNlV0wdv/Iu/DNCEvJ
lGmNjMMlB/VJH9V4mcxXU4CzAEwOCvJjZVM/jMqSIb9TwOLjz/HlSRu4ASd5E+jS
paf0Jo8CrnpXEltWqQiysQhfyLmdFymL+ZVHZgjargYFKSBY/MHu1HOO2IO+b8Y0
uEzIp9qiWEi1ewmd/NXpvUm5Q0iSuYotLNrDgZzs8v9VkSXtQpegEewgTbiiCkri
yVLvvuKFBIb9xnaskJmAzDqk5eIg4GcRFCzY3gZmH5vZtj4KfKRM1F+1FdwmPfqU
3XULffdxycTDhId/uj/Lkw+m318PvB9E2OZqyqKiDerwJH+pZVbKJsiSjhmIDG9T
bRDsnsPdfYpIt2Tl4pBlH5A/8vMJfw6YPB30/CkFRark8rAOI6NPVVeQkDuYl4C2
L5cFGVcFz3UszNsWi/xFn90knQwoYLUUPVyhoaS3NIXF4K6hL1/QWGg8CjZFYM/s
OpB86ZuQPF0Gu7zflETv5RLyqT/Ph6nlHGPPaar0swj+xNbYbb2DH3nz480/ZFG9
6ous7UIfPZiAImXtWtazg1rbsHPS7x68zppruxSVfkVtil/IQB7XwVmeLOeG5Kuv
x+7xx8qTDNEnnG3SX87fws1JCgiNstPlpLrJT6F+JXZ880IA4Ujt/5BUpsJgm5SS
yAIvkfiORBLmL7ma3UiczWAof/LSDiJpaeBhqaQJnPnC7zoifVHH+PNvidgLDHwH
C4oXqQbEFVuFK7zl8vnqcLjNV5Emw16HsvRdtRz4b/NrUXrWBWewGY21jiUgaJd7
Ou4Fe68Et/TYcvWTISG/FB2LBp3W1KcTg0RCmP8FQ4iRRew+j1Acb5tzGEceNtC/
I9CFyCCH444FJJGI77vICFI4IKmNHfCItQY/lqsn0oIlpQn4YtSolitcuY32omZ6
BJ5F9S9ysFVgwUItAEUphbq+3wgYLOAm9mNINnS386orastTWqyA73E2alnATsU5
3v8Sz8ZsZ+7evo3QdG72DLTxP7ZCh+Lh5zJUY/t4p93Gtmg0zUmdD3rPuFH5Nf4E
CKlXlHLCKhAcPcMcws6nr7QJCoxF/1R3FbAfOAYkhge60HLThY56LJ/FcEUeiZ+L
wfc17lDp4DyIJCS/1/Ce5dHUzlAOlKmF3BH0gH6qqn5zIG/KRWLAi7NLkwxt11te
2a7M4sTiDspYHCqD5kG0OdkJMSVBTx0LlEYVEfTvXCGpPl/9cvi4tZx8j9FYQAvW
MoN/uih6tlegrmsR1Nh1kRgm63E6d4zL5lDUW9pt/GYVO7kEPDdDtF/EVSQ5oTmP
OZiS9r3jqSLFiKpLl/ioooX0D6sCZWZN5B6DUC7+PLbNWK3ItoJeYuU76FA+ofKP
l8E5jDM8dx8omO7NFrxd59ZUBOQir26ZHP8U3iGfFVSX4epJAxVvEpxF21NpiAxo
8kBoI9Gp/cvk7zfCw18Y3iaIke+EAaTxGQGHtSu2ZZL64TBM5E0E2Tr74xVchMsB
CtwUQpUCPGgnHC0AbKsQmNNzABoA/KlAi4Hme5w+z3PH1M+aJmFrF20IlNEyvOks
2VRutiMhY4B9/f/vXp1w2c1kaEzZxlEy9SgaAKQFZHX8+zdMloiS8e6PIaED4p4p
Aah8wslyHg6huekQcjDVDG+whpO58vn/QHF5svvzg5Yrb1yqYMoxs5TycV567O2b
Ru6/fdorJaZsZ2b2D5SwC0/Vmcem0Oadi53pbYZldH4Mx4NvPDFpjr6OAIO01pAg
FNIRNykCfedV29dWJWznXlZHHzLUUCYxdZ7xBnJu7ri5JVi8E6MECHHtsnpK1AhW
8UxE0hcgU4JghrWX2pMiQhEFrl3F5K7S5NaGu9NgiprOMt0yVerKOgRYIpNlv0Yv
pQoPJpIqM7R97NwdngKP/tELSqX5Rf/u7+6d3gBCyA+aBpo5GboxK1jFGqVIJFGH
OFdubyhlm53L+LgBMlJCbrz/cACrmtvC6ReoABHdLv1dx4LagCy7uR5X0VZIddED
T+VWiCTSZH2ST0LN02li5rtTz9NCycK4dGGC2trSiJnvKYIhnU+XrIrt1uiLZ0JD
pkoo4T/SfJ+t9cEC2DgdYFCOiGRge2ruWxRG4yJLlt6sEg9Ek+UW+NQ7HqXLwd/O
9THVeCcyeJHoANcZfmJeby6hWl4MNwo4pVzXfy4YrbCzQDAXRugpQKjg6swcY223
LWlfwdxLLACFo2z3DEGcyCEOfn9BRqwhg1KNEsrbzN7n7iPzJdkJtm1sMEOoc8Wx
/v0g/9rOv1pqH36jL7mJDMb9LF7Xvb4WkAm3jZCITmqcEOC1nyK7aX3Sdfx/JzUF
jgh/gQCTH5lHGr4pVPDiaD1BL2Vmz/xJNTPedTarRvXl60AJRSl+Jw8QrfCoVsvu
FQVH/a4frwmkolWeLcnKRXbaOuREcdwNKUP0uuXvgjFGiWKhdUZR3ZZ5ksQpLBTX
eq/BeoGP1+OUFtNTPgPAoYaou10bkRCq9feRsSEUuhWryGQcJGBJw2Wbw2S2aEYV
cVOzG621ZvF8iaVKKqPC2LVa0mL7Tb/FWIWx2jHzPItZ+LYW5pJ6Rtgv0Nr8gsaP
Hur7l07YhErc7yBnY4kn6ax8IOHPW79qCTrTi5FBixWIqispKU0QgyNLNr7IG9Hy
rwNqZ4AuQUPNssL1UXkcJFSaDXpUJAurKW2cjiJ9rykccPHhNqekBO64oyOL7/yM
zgCKQy9qbwOF8bU8ZYMnLAjV1VMervE3jcFLcIrdtrQmf3N1UaDuJeD/QjPalgA4
IwohHURAchPULn2JLRbr3ZSs8RR49ZrfbeyytI3iLIIdInMXO83vtOo28UqqGsDf
DjNDY5K9xR1d4BCx9+ulYTNIO6xNUWEgRPcrzC/rpXCSOwqBjpAYrwhnzlqs4j20
V92lucVsA1q2k5nNLvpRQ2RhEf5uoPEm6AAZECH3ys0E3YDaR/ziu5uVhRTwuObY
AIuP66kGhXh27534k3abZDCe6mVsPq6FRceUNhfuxRY/2+ynvZAyuv4YaLDKWiaX
EhGTn5xf9IMzIhIFrVa4ICRfI73m1huqfZwYor77+6+SqWGMK/9kgEWyghNPOqE2
LW9XPgj5he2N7QxWzBepQLkZnSs9ICk3xGcadpeePtsHTIrp92VPi+hZuVG2OWEx
9ivtMC53NQlVWh/mtKpZQFXKiWr7es8AEGmUFamR+uqilIrS4bTw0TY1RzS0qkcg
5cT5SeqeT3G3WNsIbc860eOazALgD8081xB7Rr3nqt5UVhlRKMmZF8vJ8AInYzeY
Pja7tpcz42P/GdqYrgNlYiDbVNX2kTNrdIqEslvG8rAhYpsvSC5gwxjMoKhs1zNm
/IzZ8iQ/CqlYefBSP7f1jw8fKrXtgv/cOQVsaN4YAPGfnL/STvBihc32QKKn0ZR4
GSnfGwAlXRe0jqox3O5ok9JkNh54vPzxyxFionvnmOEXyJbxgbxvoJDNx2nWG4Ty
xGtvWXB6esHA/ZJAgaGUcWKKjEWiWTWMc7tEAo8tyOw8GK3oOSWh6GhgV4M6VM8Z
85v7BCyjWIWZPfAmvDHcRerccaDKuC+6R/lzE9iVfGG/NJ64gSysRRgiOlf2kTax
zRrofhbvPBtq13VWjh6C1Y+7od6C8wWwV+7dG7UapXR3RV7A3pyhstL514Pjq0sf
EAEyB4HvahCfkwTnqL13r4yCunePsu5lQZ2M4gAFOJBub8XxWqq6ItETkePug5eO
9VL60oqv2SYAzR/nUDpPEoHvJzhZ4rExBoEfZkRm6qQUUP1ZAdNYgDlxUvuB6FTM
+HuvhI/8q8C2jAMhof+CgxE8f1G9U/5DKx7h+B5Li6z816K+RvHxBkedymsO+XUH
rxLKb8WZZTgza56uDu+Yc+jAwI1v/wKf8UwWGPhQitLC2VQDtR4sH2uZ5h+hXqvj
t1GBPAnqoa6IT1GNLammmVzjeONne9xY/WsySO1Njc0kwl/gSVR1N4tv9pfAGBNK
hnckNcofuO8q7WwSQX1mAgVnitjUM6TjaRvdPH2VxKO5fMBFh8ZUo5VXgfycs1nW
CMbecJLXi3Ql7KTSseJVunvMNB4xx5rvDnLxcLLcVLxfoK/CGVWc8CA/+aivVHgC
zcrMJ266FzffjvrnhnPVQfqIltKsgWN3DP4GM9OC3CVoYYkayneFSrQIleUd62nj
Ktwfgl8nNQawYJ91lhshzWkOY8unW1caVbnZvwVW7AgEwQhXxoxdUg3ytvlmcVya
xQzJ1ppSK8cOBcgwRE5DC3UC8t+B1eQ7DVIHnb7qd+IL0HHVe7G2CSYuSvfKX1X7
1UzBMj7K8PG+cLsrYsIffMQzp1LvkN4+nf6ydEhzL90+1Oq0RMddSUo6YwBqpHVS
J9Mkca0LG99fyFNzJCxrGKpVS9A3BcCuu0IL4ZsJ49mLSxR0iMWdZNFBjHlJd4fk
5+MS7R2MHiJUIpti0T3LQI+cGk1rEAjNFeeSMEO3hdAs42ibOwzP8YpELYSvlQow
ZL2j5Z07qnGFLYZIawX+YhOXx5fnHYCXbO6S7YNA1/xpIJ5+6FpLXesnCyvVoYFU
vamv7qNF+H+mPKJM0E5k+iC4h3/dBWPF1/UkpM9nwOpYB1cS5gUIrkelXfnBaxxO
JW5geDcxLzUF7hfR3aGccg2j5DgHn91bkWnsQLDsXQcM5+AlyttqRXyWgpEQD7TD
LbNfRvXdKKThWI+I4/KR7VjmvJR9GMMIxgNQRzDmLZ6YQSmpXXIpb/BUc+Gt+aQy
Aqw8JRC19fUSfU7TQZh6phriFrHVabGauXUDFFnoYvVpyTdb6z0dbGIEtNeb/UUP
c+8rwOdYWcY7Ke+WdwlqdF8rgyGqEVGlYLXwubIuf70CwDy91NSUpZUv6/HDqCp6
bkL59Z0aHNuB2IS0tpwHdx6tY/tbYmKDRb7edJnPPlKQu05daLqdXreSpcmdihZE
PoKAbtj14ccVYcTCC+0oLGbzW07W4IaE0EJi7rfwpvJ9T9yjt7/pSX3OqGHwe6ao
PR92kZyywWXUANDJYJtD36wHac1UW1zuw7vq41nj8XiTir75Q+xOsMrlc1hyMdN7
rixbiA6NO5dgGRrzS7hEiUEtt7BIJtuYrQrIUwUeFabwxSvoBsoaS3amjU+zYskQ
ZfrcL8LQqCU7ErLzGLTUrSolf4SvRwGDfNvQ7IN1VNI5rCgTXhdVo5Vvn22GMnuL
avLnxOLcPLzjFPw/ZcsJiJvDN5+K6AhWmt5zoNg6+8LsNfjz3P4vZALluHnnbkl1
9yJn0DDD/6XSlwp4jk8sG2vMlz7F70CbI1uLjHgMvRuJIE/BHgp+RY5n5s4ODDcl
Uj5MO6rZKwOl14+wjeAZMy4+ygi5GyV2/NkKYGFVeTF5AxP9fhUMyAqc3yDqk2Rf
XvnA16Fltgl5H7ngz+Zo8zP0T7P5XL3nf/zG3xIRhHz3EMH2SDNq53nzKzkVEPNb
gDYgyLHKUk1DrQ1AKtFhQ8d0F3efdn3BS+azK4VPegoisrAN52ZWwjweR5mpFEYI
q3krSJcIPZp1R0gFnA7ZfKx3Zr4aKgf2MsR2tZE5sW3j8hnVs/qGImFQBWiMzgK8
P38klDDPTXy8TJqDPIbIuRCAQ5e2dbDWi9yvpxrp03aSVHsYroG1WnMzKtEvKU/f
kjqopxSpGMUuMGPiChnYkse8FfN5+aBIhi8jlKBrsRyOv/SyuqMDviUPOhRSOD0O
DyL45AkOxVe8BHrcrd9rZXCxZc80q00+UtlzAw97WdNZQN7yW6wy2F+1HlBiL18J
WUvbMlOGVWLrvQa5HITlabFExyoXq10icx0Dy3P52nYMXkYoQtzhya5qQhck8yHR
+CendnTI+9jVmC9GRmw3IfCc5rDIouRjR9Dcyw48AdoWFjoBDGUPjz9IU3tNflO0
qnPoUSoktzrXa5A5/rb8GZEb+wDAi19OivY7/rflAZpQH3rA+6L4SlW6wIDW9fCQ
EvVZQtxgWnBJ9J2dVxaDQy3zHxRumgrCSrj+9ZolKdZyiC0Bbpc/IuApja3O3dSa
WywEXiTyDZK/dts017N+2S4dZ8Ef5QO9XVTu/g4zcnrjdMPYoKYkpgrF0Me5ofBU
NO5GzntPvP7iTnjB+8NYyLzF0L6BJg7tPJJ2EPRroUsHxzUxJfXURxt+beIs+aYM
kkkCI8sEQV7Qi7RIUFUWvXFq0EPsXXa1yncXT20z19xu9Hq8l76dZJLnIrnvjTzn
uAyMpGeQPvjv31zr1u8CE1krWZpJp8v2ZXaNwAlV2n72RtTqtbEpLx/1GwVnsjru
aGP83UM+laSpSE1rX2VOjdXfEjfxnRdSb0xPUbl6FcazyE0k1nIHCwnSElFEHJlh
aJ5SpQSm6YcZTovVVBVMFCrHMOJ9InFi9jtQ07j1337Yk/N9efUA2PG+bgNp3QFn
udOgpS4jpD5phhqLVjRb/taYxSgUfV8QnCnjvdJWc7H4BiVgK+VZaKL6qyytHhVK
kYhIK6mebBORu3tP//PerB3mCd68z3LBhJNhYFnnhA/bQr9GUI0MZO/XNvm0DERH
z2sW0hRM6rnVL8v8w/vto/fOFzlUAg5I2qDkuxjn+mqcl6GMmLuEDLD4AWzl+N2a
5XTu8xO2tCBQwYGJSxGkFfwN4LuyCTbNBYIeNdyEoGkAq/rT+Od7IENOJcft0cPy
SUpfVx2LLi64Kb17UvVlOu0YOP8Vn5+QZbIy9f5ibe1NhHjEg7xCrcOft09nTVWB
5dgaJKa7OeVgMx/q9zxcbKe5ai8oxoeFv3ix9vsL3nwVLm3cejw7Nxnj3XdhUEM2
mELQB67eWCpOG/yUavAvoofW6rBeGK8evjfg4MVVodrET/Gn+ApLuy0gOw918T0J
qrXb+3YjS9msA5lDiwuneCOLsaL69K2g5RCQZ9XRGOplx5KI4Cr/271QXzKahAvP
Kyx0ugNlQY9XNWjtb3dCfZMKuMUaxZJ6o98YVrzAU3qasQEmHKGaf7r1ypOYC3Wz
GIIuutgPBa7wKwHkMfS0XR9Tg8udlqUqvsiOENAlKftIZQwGs2t+7zdHYE0Imsyv
zd4iVACFlT+ZAkZXm9jSz3EAWQLk4lBmrqLrF68klHfZk5NIOQ4zrsWqEh1zbUYy
lNJql+YfaUTlOCmZjbXY2S8izys3SJXUFvm8CZtI/lxZ1NmDw6S30VAY8eOz6XfT
HMHc5Q8TlSNDZnMAyalloL/gOcpMZuQItNSYDWOiEDGpEUwd+D4+z8sb+cYVAHNi
jk3GOwrVzdIAgpcYT4FSd9Ksq/uVrH+hcA5tDCWmp4PMi+fbJqdCkfLHfSH++TAt
k184h0g4CDQf1FUYwnMUeBMelTW8AeetbPAwSWmiJ17dc6UADXajq7eOxEOvwkto
eZ07Xg1t/yxO1rgRxlqvXWwjsIAxv+FaljwG4eeciScRapXSCTrXlcwNgqGJEoce
PucbW3gw3123JiQXsQ4Fj3nJ516J5qSxaD9L1QUtPHe6zCEJa7J+aUK3hMwerHMU
F2hpSBG6OPWCkG58OHnN78x9z6n/h957tAfOOe7kh1+7oKXZXfeTtsT7qKAEcIlh
iKTRl2e4Y96kzJU4IVEnoSsAr7+zhaPjbUj7XW/YJk95F2f8KFhdDXzy09lAx+T8
78Rjr1flCGDam7IdETl+ieGwF4pSu61EDYvIHucolZw7UJHUHLxPerSdE+J6CLqR
m05stWHMaiHzCIvQi+c4dU3Ci3XnFqNtpMucMxcjKd5cOZBj6SdMiwQ7MYC2dNhh
HuKr6VgPbuyvfy1Get8cJ8os+wCc2P9YaeK8NLVWqChWNECLI24Iq5+rQywPC0YQ
micoWHwz5UF9ZhwGr7SiRgnvCdorHm8qOixXD8wVn2fXuHRunY+aSWkNp41zWE7g
Z0e/XlVKJZLGgANRh6CU24isRE8D+jPGMIrNBTCpoUWpfB93Srr/rlJD/gQX2JB3
3AJX3n1rkT//Y8x/9PbPCly6lHC8dcymKRFNms9h/0V7xHjxFsV6Qtig4CscvTVC
C9KB61P12zX5aua13dSK0hSh5WJXyb2VBciVn4peS0UOhBSD6laC+b4poKyEe8q0
1Sv5I0+t9XImSTQQt6sJEo3a7yG50FJdzDJff82il5Yd+HXK1Dg7+21FKNGHqbLH
2qngdzwAJwko6L3CUpUDej7cXXTHPh6T1ychBzTVCm79WfSrvNprttrMlgL0uZkl
W7ZoiQCYKnkUM7c+hsTaZJd9mF8m0pIw2/TpJG3x68EEsxA1iTJPGBEYa7OEGXL+
NGolQCXILd55ssZ8QyWsM2+LhHIaPzyF9lti4H3j1/CdW9rCNejqvxbRLlCXR0Pi
JEvWfclei/ithYGZzg45f+p3upO1a1Lhu6HUufcqSUvpzdYWvO1UcwjytWfnEgDa
A2+iK08qcZYH4RQ5PqWI0kIOOWmKa606uwwyLre0yBC1oNbptCP/pt4Q7s8DbuL9
zxMySDxnUx7OdwytRMBd7fTj4ZbznANvjSXp7OR0OWcsu8fDn7o5uk9ug3HVfXVw
2UN32e/0zloQfkQQRrwjLPSMIkoO2FKoBKaDCjQoNnNM3G1hwOwtDsy1809TZ4km
X97+nZa2H7A9nbJAvYoORRh/nTJJqnQNmeYxikzcQSWQhvbl2fqF1GNlX/R+SVsl
N4HWaGYvV+5GGXajA1Kco4WP14KxfJj7oAPhtSiq6zeReGZHIKGUqL0syooVgIQ7
Zd71z0DW6Rz5IhoQt57lxGpLeEnfXVJp/FmOV8cvwWC9oZHQIxHvWlT3n4ZsqU6U
GRquTChY8SSx6/8QsJ72kwTliBpilbrI6h9ayjci7VxpCqwiQphKRgHnnDA2ZAW6
apvaQR6He4wdkXDV0TF8NYIP6SpyB7f2jQ+AXmEZ0iS6eyHYL2M+uMMgzYwQyczH
bmhPguC+xgYhm82ADy01t8eYpPYjK3WvzJAmkd6f8EJy7iAKS3dleLeiB2/jBXIw
tVAak5aUb48Q+YZID3z1Rf/L1Jd0i4e8+mhCrKJgQv14sNWAtuXbIbR2ZoumdcBW
4dH7bypWwKge/OPDY2Nlw7vhsIninNcKjdzwJy0kvoCq1+NzagHPqFa3i97Oc0xr
REqPDX6LIBO08GZHzFC4o/0yn8z3GQL5IuLIRnNZ2k85GpwKXtBSXLDap8RsfyPp
Tmn49FACZpRoxJfY6wENAeDUF+RKZsPZR3VvAloPhdY9zQtKk6B1F8Tt1u8UKQtn
uSMmplV+VcvW9Ee1MBwHDi+1Wp+93RwH2pGbB/hUnwrZBlLx/GmkD1iWMvDgjy8G
jnkyTUVCJmzvWWv206QCHsTxS4BLgDbW+1NoWZu/Nt3+M0W+0t8hsOqy+ItQ6fNd
4gr/ThLOwksJ84mOhHvT7+duBds/3ArLxKn1sFJVhX6kd0/h/G13CxnMSoIVz8Kj
ujYZkOol0aSq9/2ilIPDY5ppcnBxCtFig+RNGjKcknownXgy8Gw9qKvE/fUagSo9
0Dxa+rfKFdtzMwhrNY/gmk58M45cyjGLm9jhSJ6kq89/wy16qFwAe04hfi0UloT7
knyu+xAhEmTY7g+EoCNpZC0zrNIwpoCriLutS1MMxIWkQSKWWjFPjARO17lF9sfI
iQXrwBmF5JOFcUhwOrK1LlzO3G223bBzkw5yUI4U1yCcxCQPod3WeHb/FTdnGoJP
0H0RYAqOrvu/yQ/qqZV4UeNrV1rD4vCkiE0BKisKRi5dU5ah7A52EBd56TTALGtP
T6zE34nWb0DJUcfncLO5JRLS1hZGkGtXPHt9txiL6PXsQcEXlH1g7wUvMdlbOIfJ
CoqvMO9FnKAlX0AHAay3uYU/aKXJtgAQsL8WGEYXfZJof3k306yfnsN7108xHIpd
7ufUE3FuaMD7FDM3Ixk8iJ5rikyZBkKmDtcZFDPawrYtKn9mMi3UCbVucsoiFOHK
SDrHyDtXPl2bMjeV18EhJciRxvlLPTQRZqDiKVMMXbuC/z/gPGLkc0jslLAqpu+P
jcdn5236VbOV2Cf854JPbg==
`pragma protect end_protected
