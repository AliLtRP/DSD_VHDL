// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
RQWK6RtMOix3UNMQmsHhFa166nuAFxe7RaW6FWJZR2fygY4A0NyZmmDc/+5MDHqgMlX0XZv2iF7F
aynUg1GQjYCNUaNzaMbe36NE6/IrgYsODlZnkzRnuKk12YrRomCFmbTF4RjPFx7Kup2r3h315t3y
9DiZ3uXvOI/YbAn4IABExk6P4z9sdZNUhT+z1WjdcpzQIwlP+gqfJn0UvMz7l9IkQKL42q1W8ayl
atQpwUeu35EeQapefRhR/6jJlI+Jr3th5EWexWaX1CanyQKAGgiF0mNG3/+4DW6Q0QclfapcXLFg
TeEpVJdtopJ2CDi5Ii+XBXDe8u4174qD9YxSmA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
itgWHJjcjCJ7CW6apdP3XRjNojVhppYY4N6U+96Uun9EWLsBqpJHDDxR8e83xvMrfKrRQ3hAJZNg
M7ODgQ5dA1mZ3ESzDCfofJFA4A28LxQWCE2XG3PfmQ0yeyW5OZQheSLsQJRmVzrFzjYzLPoJYqSV
rPfX8wBjC3KCSPFTL/BAFz2x1YEQJT6AL8Kv19FFcjib+Yna+KvqC0GrXa8FcN4BcqARsqiKdeSz
pniO+gYqKscqhXGsHuSaIjE95lrYRYohLTdc/PdGV+bU+EbhnGzAT0u3c5p6pcBVRYnd5IbP7foi
JYwTHHUHeOv4nF8OXFd+SFPoYZTbF3aeL0EByjYiez/3ANUtn/qOG+NtqWrGQsum0fK4Mgi6DsUA
YCNM2ikNz+SwVZqJKAqycvCVVrnAAEMCGJWCH2r/aezZYZioTPyVKQGR6QReh81NVHOz89RmRps5
dDk2Qm3W/0DzmDCfB5YgaOx42RanzVl43Mye4K6IcRRRC9qMdpDmbSh0iEU41i+odO5HEUEIoDQ/
TyOrbB9RHafKVUz0SOMcP57o91zUYkIAy6AWExvG4QaqUzemZzRg5iWuhkm+nQrwCDLzvXL7ceUz
ObPCWDWPAGNUgBGGiO88qYmtK5994uAygfzKk3cU0SifIN84Fd8OlsxKLX3GlwdO7JqI236ddfh4
W+vQCU9HzmNi1q+snC6Fcd3AfANWKoqDiJByWKhhE0ax+FAWypD5LMFwpSA1lZw9UkDTjDSx7X0Z
QK3GHApwnJKemwbJzFCH438qKAisyveR3rmUBmbyDz4U7xq2RDrypH6Gh6I6U+otqIGVo7lJNrW+
MLeNCEDZ2X0MFc94j31FgglGBAqzZWI31BLnuf+BUtUeKIV2lrNWaxZkCCBtrgWrJmq6Dk52F6Im
7UT5fMsqx0xl330vFQG564chXRqG+lryu3yP+gLx0vcytYeRXfCBS0RGUJ36dS/klhKsHRjOTGfU
pZF8WbLl9PEPEDwWwIjmDc3Q7TlpX0W8mJZwLh/EKKDWJMFCKteMH07CsMsf2i00+YPcwdWrqTUX
UcPcSqML4LyhH4GUsm8Qgu8zPhZ7Eg4HYQiudm9SWhcWew2un/7AtF9tVxcYHksIG8zuWzhi9CHd
rJEo1jeLZKuqumOi3bXsKCEFyN+pl5p4Y5KVulQ1z1yOpCQjNpoJsXS0+nGYDBGdSOgsQYAfcj1l
XBxRJOCYoOQKk0D82wwqS6hiJHKPqeHt7VfzNb0u4QKZlDdnF7JWzpHx2Viu9xZJoMu3mDDK1cVN
xzgnuVxWohE3NbCtI0FOn7tupMIuXxe9WQRhU3auGPXUDgCDo25dbAnhaxMxtW2raU17iGZgS4sY
dXjWBPaVdc5g19nx5pnomin0FCSIEVePSj1cpzP7syCfyRh6gZvXRgx+A4uNqT5oegxL5mnVD3ua
4XMESsGIxVfR2CMLT0OMEyRMwRY6oCiUe5DMwMMWnBjQF0xQA2cs5zAcN0/XB0HlL/KQVUwj7yzd
ccn0ZPGGa4qgAQGGJgZkbRJxt9lriegZzc69fdCa3glonkAlLcGjW5bA+7tbun13SjEmS9lQcof6
DRgGQ+BlO9JT2wXKMpuuTEsWVjzcjsP2hcxY7Glsmbv6srwJxkv4J8EPBjIQiVEj6vw35GqIMEBl
XCG5Y8Gs3U6hHjo3qKPIDPM4PsYD2I1S2uJnyvhL8AEqMtslK4v61k4DaQfXUPGzCo7S7if55lHv
ZpPP99SHXlOVDLdcxBVZsb/gc7y8kI8PSID093agjUpEJy9yODBZ1xuKXrwzj3Kfk3QPd11Y+OP7
2hFbh/IKXMROsyaG5ADtcP3TN10LM11g2O6M9vFhudyRHTlgCFCVKDRglt5BXwzNBsqHbeiK1e5T
Xdk+WBy3wrqO1GL5XF9BIvp3yhsN0llrzJpIjUA8jvFVjAKfn60iaKZ7RvwlJ/vyaPMerD6W/3oY
5TfnZNlx9pzWlkqPUld7AJx26/RlcfAN1xRuNR1ov0lPQeRPm6OMzO6AEiDza+6jTDqkMoA6Xvw8
K0MqhtJTiZvECu00z2JrM6ky5L5A+0vDgLKrjjeJLK3iL+TlYOFkW3lka+YUPTTZkGhcULcJ0svJ
qwwEtmuef1R/04DpD88u24XAd3U46uNZ5RfVIkAMi855TgeQBWBR2DPG5sMuSIfT3NgdTxTpLC1Z
pjQ3wFVbtlSNDSxymweEj6po99Ab2yJMd6t/HEjR2Mg2MM8rjRSHpQhvccktqbkIMSjlI2S4BDhh
+ovteaQqwNWPfr8nNBnPR0r7JK8kccU1dJh5jc1a7nkRQFCr0SSPgh7YuWWKF7loHrrzNqmXp7y6
JK9Bz7wY2JoXRHtOAjMNC0Q9T13gj9l4ccRva5aWK44LMe+shWozysjdF/R+RbNR7QcgHZykOugE
8DaBcl2p0//7L5IliIJm2UVYQ7SeLCuHui6o6gNHu8VQvHBL2SjmVWINnOrvAM7++Wmmhl17XKP7
hR0GSdRD44Gpi/VpTbcYQOUvLP320Tu7rktoRjtrLVj4GL3YT41VFJDTU6/H8UPV6yqKhxyFAgCR
xUIu1js/nFFr4ZN8L0HAViIM7u6RzfYOMeWClITJEMGOM0eYPWkVeGp48n+t6m3UxrssU6e+DgXd
OUi5wgQMrq8JkzagPZOp7zevy72j3P+CN3ZCJzcwr9C4LniPwp5UATST6s3EG0dZGs3I7QgjCL2G
LCrrTeH68Rws/g/ZKOVxH4B7spFYMVgfEPGGdL+Jonvf0st3GzkBrSDOxOlrxEOOuxhvPqJ31UB8
4hY+3wG694tb3SWBc1Wipr2jNo5zYYK+CAbpXRc0+WIoBmDvQSEYuxK/0LxhftYX2w23DXgeuMif
Z6BeAcHYhxcZqjuY4R8bEbZQWvdzme4LDJbfH+QPj3Bm3FDD0bNduoPyKzRphi2kZVbxbawTdIZ+
FgfQAmEA0faUBVptKUW72f+3+mTXFBAETlrfI0n9UdKVLGmJEQZGDc7o46BtxZN8kTKWm6i62xql
jojInnjdkQ05rTFZfmAht3YBHYabuP3ReS/ZBynuzperkOKueTwtSS6Nsm3/1iMatZDTGl/ZJioU
8BHFs1ou3afMxZ54E5PWy2b9LBTpzuVGVlmmThacr8PKkHmPvZqN89puwZFPQ9xP53/sl4rAMcDm
WUQ82iRiPJIRh5HagrpGFIr7oUJUq6JUWgyxterjhAjhJ/QqmErKmWuJj9UXOQ40Tsgx8ycTKELc
V9ZXe+H5ftZd05bqtH74Lw7ON2eavfXsJi/zymEEv3Dc1Nych1gMl5y8fSiLppVw0fFnHiJB3Zoz
GzWbNxU5YYIqRISeod/qbnb77ukQgU/4A5CVktJaYnD6Gfykk64c4wkvY5+m+uqjd2FhJB/wSNye
9qrnOQGg9LQ2XvFoHdwHA4Ey+HtJqS5pYApZU4+W+0HIt+2KpXx+hisIdDsqWTPGvt7VLYT50wEg
SAvoNyh3uDR3gVtN6swKLbGQRQFEczofodPJdw3Lic9wzqd0Kr4hazwvgUA8E6ycbPnvI4Wl7FLY
++DOzyD9Tka0dp7cV8RMmKORCjk22pqLMq1Fqaj5OJTfQULuvXe5X9g1cPxw4t1pvEDoT5Vq4c0j
xbXe+96N05t0JpcOvKjh++vl7Am5XUXBW6cEfwfsRjKA+bVKmDGOUCQZrVP03i/P+147cSZjsFlo
gzc2WE7pdfUkGG7C2k8MBV9DrRB3EYemV8eE9A3jItRx4WsYwyrZ8co1n5m0ewjk4+e6kMCnPpzq
wM7PnlZ4FZ+vLaoxuI5XsHPs6omLRXcKxbBB7pjL0fcRgSRuBBIOG2QqfIAE1o3nzZO7YGWLPOx0
aGkI9Kf99C2IDYpy5qqG3mCc5jlPXRffwLKQm/CK4axqkk6Rn8KF3lWcLowg5Ls8ADPw+qjTKTyC
msy9ZanlMzOdVy/EImD3lEuEG1vHyNuDmT620RX/lkEhYLlcfvVrEOWhlzTmkm9rCGpU/o/Z1jhE
AeRK+wvzH+iia4EFanDMEZA4B6sLeq2scB/BHMxBPeDc6c3YaTKxnmer2aEbWLQDeoanVomspZwF
IfSVUFF+2wPPe2mIrG6HvsEZpRQfKjubksa4zLsaxlYhZOOZ8Vj4viAzoakki9bpsRgkKTVmbk5Q
OasXytBL+Y15u3oQy5Kgfh1wFw3LVvEyju+rV8rD3F7W1/ObKaTU5QAOpr+XXnePms3CcNeBOJEP
a+H2BzFLb5OPIy9P+hDWjGoYgVZi018seWz+lCj59wZGonvN5+0iwhsuwZ1ZwVoA851Q10yagkou
9vLdYtCpHy0VrWpeGV+C5DoIXXL3scShBPxIcF6NKFkL3lz6g927lhPPVoAM2EF2FBR+Lw1gCRAL
sMD0BP2EyB3wrffR/USS16uuSctxdaqr4LucRySv4raPFtNnBvB1qjMUgiSMGhpSc5RKvnsMPHZh
N9CWQFyJxmaSLVqPQhLM+Yf5CJuxy+Atz9Bf7pNymuRv5PT/UWRtA2O1VB02sWkU8uBWS7VeM4cu
Vsyn7b3AiFedfyHnckNIz12kJjNZmzGgO6xUWaBMKH0LtLszL7p+WuO+jP1cbBaccmsWqa83uemh
vXUcF0/JnxhVg1tMc8wOnJwVuVRWfJl7hzya/X66eqenDRkcMql8LF6HwlH0dKGybB2T5Y2nUtA3
Dwq+q2BBXDycf51QD8XVA5ElaxYlfYufVxcHB5fhDbMMuC0SSSkBGDQJmeuhndPWrokVOv+btT1Q
Q+LQoKh5albiOux/4qotU0EikxTWgw9+fVItqXM2mKhZ2F/u0T8TwMnqg/fiOjz9TImfVRzzxFUT
SBaCXDy5HagphXj/MYjJVobkduiIuQ9zH20GiE1TtjKCkWcjtyRiLXk7ywZ20VL1cw05Yf6Fqg14
VhDrzg2yxCg/i4T1dIxo9eLN17TriJ6kVuu5IZXZKMBFNv0aFVaKXgasNKMSLk3Y3hjZ6ybN/p/z
gGrTSbqisqjsa0bqTq/vD52Z3ijppBSBtWtXYix12o2oQO6EfyS00rIAb4HzKyAgB74Z2YC72U3A
PqMZoUTH1/btQvJyVtBwHws2wytYs+23LjwSkWnuYIb25xOuC6Y8tHj4IrMTPxiqF86N/O2TfCI1
uFKBa38BRlCgPlEu3K7Ur53oGOFWrUVGdyv3HA/S+3XAiZmYn8ZgV3jM3Gdwh3xb+Hk5yQng/ws3
XgJ1ImTwzFHebZwT5QETNVcOuX0wYF2lfEF+vdL0a2r2EWFyXIzlHBOupUD1C4Xmzpv/dW8rmHHI
qhbwN0vHqGP9vAkXqi7ma9AVzOkXrO2YF6LKajdsxZuN+DiiaHBDw8Ml+mbC2G7BwRn9+XasdmQs
QVvClK8vuLhVvuBOPt4Om6ZkFVBzGfCLKF+y3b3JxI2ZdE7OdyRfSG+strxLhOlPic8Xn6GrdqbK
tJcxGz9ObTXdHvUgRckXbOAF9UiLb8mbpby819pJmamBp/fxdfdm8wfAbSYuf3yZsDi8tL/oeEEl
P08Im/PbjJ9zUboAfs31AJ9uEIgIPY0nPt/+v04zaDrQ4gOYppbKS6pF+HTsnDSKcugz2cQAEwjQ
LNLW42HscPBojuLzqLk9518w29EvVZ5ZrHpUnSufGFDNnEoXJ1lrX8v7PWqkEQ8aNZrTXMiQSha3
sVGsWgR34WcsmHR84IOorvFhdpst9qRJtMgcWbl6qRidNk61EYAoXmaC0XWGF3OIYLShEA+K2kKf
JIEDloww3rnLCxwD1nNpwv0/XlwuKJOjMPEPtyJ+r/I0hd/EA05+zCU9MOo5eOmZfSU+OfL8VzXF
tW3Oh8yGhSLg6q7XRmmnNeHsEkmK0tNt0aThWuemEPV7KmAilqrKA9ih+g34eew7cDKXEFejvsgL
qwxqI4CVtZ0qcilFjFkM9VXfYgOTGlURACVt7mvMbJ27BGh1R3MD32pl9WIF+zBAKNQqx3Etjg6c
sVS8XbX2XuOOG3Xnd/NTyPgYNwlIfjCuXMzei4qrcJVwMqotXrXgsm7PLrDC8T6KRr+k1S5K5FYJ
htWaLAeXRai01gcZ4CV2+aQyMv3WpnACMqwguOT9waUGRmWRb83qimr70wtppn9hCqSlgmqWsaE4
xxk4QBNpqnUhFQJ61KiRFJSX1JdpkggBDXZfsmgqqIKlxcbpZlZZ2Pc4CNb4VYyKu9AtiDhvdO//
E4VBSIn1YNWs1mj3FIGo3ffMylv0dWCUum1T+mPBM/LkrK0jPS75aIctKlSDZccZG5c7iMfBCkdY
dHWXQQUrVw7Ci0XHrkFsZZChDq0OcyHRmdkTeRgeS/1TR0oqS+tbYAng32jOX9m/w7hPZ+OrhyOi
/e7zdJBRefIBXuznK9Gd1vwi3A/GjKQDobdFyUe1L01TbjpBOa8QUqSalhyMdCO521zh/NwC2gzQ
oJgqFUBmPpgGcrWAakXYpitVtpm89HxJgsJTGF2hK7DMeicjQQesa/ZLiPa2g7xctah4DnRolUX/
fpDvKMzy9CHoMGmA8efOXIP72yU6pP8JCK36DBELHOmhiXAGWRVB08TXQ/UCapAIZgu1uKQf1FBx
sOv3YlZZZwc2ztxbMSuZLr4VaUUihVxkntiEzv+jOHrT83MQ5SFRWYcXiNHcwuDdzh/TkL+xmLte
VJ6bWp0TI5ZlLiTZ6pJjoFnue1MQTU4PAunydNwdGktlXlDu0W/vwW3vch/WQAKwavTgZEXeerry
2LmM+WkcIxZ84omyc9tDM7Buk9qD5nXGjioCyNjmxLVH0ZUCvwRongk0cw2ZzKywk0V3ATyt7ASe
XoVfjRLl1lN8E5dWkKE3uqzx6gPIcAyHUSapazjdU4FiuVLhACStiqicFEIkym/wGpu7Dyx8uUva
Pm7ILE7dNEBqGbkbfJzYO6MCywL6K+Tmadd7hUi/x2jCfw75Yvbk8KYQE02CmFvEVG0ub8muJqDV
KDOHlalk3ZfZLhe9YAn7plE+qsde3mgWhwv1iTroIXJzV2DD6QtzHc6NY6cnObn4Y78X9Bsj3mlx
/MONTANimPf47k+TsV6+n2oeep2jNzc6Nclo4co3YN0fAOu1PjvMZjMwEVTqwTykRclskO0ti/ya
W93PbnfnRDXRXJFWzUiBqAHYk7NkXRS9TsKWs46l3zyXC2PBHabl4A03XZKChAzj79aKut4yN5MP
YkeDGvsRH/tHKrLLjRZ1NsvcUa3DSqoQc7PcbLPM3GWZXQjj/NDPjJ8xM2uG1PU2wXWf6g8claCl
xX5y9rXvRQz45qvmaBg4T4f8h86bpDqNlTYTYUn39d8HyynxWqC5tfk39r20dTJ2YfzScg5OpOc7
r1XNqIN/zbnlsjtqQW0KKCrRhHzEvZH3BPM/t4hcC9KKbmekhDb5xkJZaf0PH6e1KwzOMg8fZ/rc
XAnMeY5t6HKsdtCfC1zc1n6dpXoQ8diTlfpBXjtLKZW1yy6z9IWlEBnyry6Xg9rZH8lApMGEBcS7
+UJhHCsXUQm82yX2wFOksL6dZCZQcBo9hJ9QxJ0Dfx7ll+9rjeG4ohNhBYsLo1YTBKVU21f4F2mr
2j2vF+8gi1OUPhtnCTG12/+OnrXx5buE+vE2pTOC4glIaA4pKHvBLvJAcMBRq+Sp48FEeZre2yT1
4yfO+Pp1rr0WohqjMr2oUNvY40hwo/b7y9q8Pae1NogVcEEuyNJCICVakw9TKL1V8mmgqPpqCYUX
A+PmPG4sGaUChbeMmV3BhZkDzaiCfqL4h4fuDagG3kr+1A5vZJfBx0FaFsaLp0o2T4D9Pj2W3oZ9
uzstq1+yuR/w1M5lHEtwcCkvWfES/SnU8exo66X+fI0mvzcEvB34SFPdXzL4zsYESZlOJXRpwo03
VjTZQFNQIaUB8HnKeyQzeS4z15KOCiNtheIDD20Zy1UUkBMXn3y1c6dmgRjgllAYsJoCYhzETc02
qGM7+67O3iDiU3lwqiSF/7ltOdDQ35i4HmuAThSwikWhrE0HYIdf8YfPSVZ7SZI8VDSgV7eHv/64
jzI7lvhKEtTUChzLvisvqMDHYUJUsZNud5OlRdTVCN6k1+eFZRSpxZmwQ2shPQ8seNhFYw+dg9wy
2bBc/Ipk7tjRluf9mdE0tLV+Zw7YswaA+WPkdghe0nEk8A+ypNuViKdrodMkUHi2V4js3XaUnNse
7B60vbxH3+sSQ0tHlKrY4gF6m8hAIiTrv7Sjgj5p+itx9P380+Cri9cBz5PmzF8eWpSOfSBsdpCq
XcfAIAnxV/Q0o+kuMznQgUlVSYpkCbXsE/jw7bnQ6Y9/Hja1gx1VAyoyrDGxApcPFfTOGul+/IhC
2IO6Uuvg9/KiXA2CUdr0RdqEVmug1fXpuvWZF1sjxw67MucAzEtSFllKeEju9rMUY7h3xo/1j0i6
WXkOcw+xwtn3RazTJQp71JUtYZ9+5xAkfb29H30HEyR2Hz95m3IFVyuOhkNFtzWxt0olSHbVWO/f
lri1rOK4uAcZJaqGaR4IhE7eh+yGvOGTLBpDLERaMcwKmIkOZkxJWNnMChW/Wl3lkNsGnk1d/nZA
OJ1+PVldEXcUfbD1l0ur3t1Aiqr68m2aZ2XxzGha5fXlbCvowjgqOasB3kIevTYKdX20Xcl2dvh2
NFo7L/bWmVF71WAE5AacR96bwt0M6Q/Gb025dr9eJSJLkJXlUS85R+3uOBsg7dTn/Kt8M3u0k+vj
dVNCrxXKq0xAEObKJxgOhcdKzE9vqPk5IIX7li/OiTT46UJFYiB1vi5GI/fJpYNqO0lTGpZw6eQz
7ICgl/xjAH+AruqEZUQJvA5QWBHAei8A7H5nZu0vOU8/uljU1I8vY40OIYep2Bm1KUzc5iaT7Sgs
qyIdK1a64I6SQh8n+nJp/3K+d9lV73pKIQG9MVCFp9xiB72pb0nc0DAAkXkznL/IFUNPyJ5TBThU
m7FfY1HM8nhObe544MypbiJIhBehlyIsLCq3z3jMG2VKBAlww/+ABVGnVRNBiqqFLD77HsrYiInY
SXyl+8lpjvnTAE/+rgoMDo2w8T4GsgYtVzV5MJmTfqorfComuLB0av3XwXziV5EPZZrnq9ShaDkm
HB2U8IV6KjBFsk/0YDMhWf//rwk+pYQ9cuVyPwqifepFD4mt2MKe68u8SlrFULSp+irXNCRxkkEf
osTOKVPJtzZQdiMGjnU4m+YJCLG/YuxB77pb0kOzimvLs+nYXG6JnNhILPCEHMW7AqLuahNnCB9u
1rXY/tsJmveybKAafrYAnuWAKxFqykUVu73gcWOMif7u+CPa+iNBBsIAKFs1zaxAxc7LBB8SyaeV
PPbGDy662QJDzwXA1bkVc+Q9CZNkgcW7wOyd1hsnqr1D8ZyVZAXWqzoJ1o4e+QMopua3P2g7J9dJ
4fWlcz6M9kwMAGszMGBMQ22+68242wvB6kHw4ednVo730XWod2h6ogGyqWQV9bUvfjXkNkgsa1Ge
YIpPqLEsLDY9QUxGz19bmL1K/wSjGq2iua6SqAEQdkhLaq59Lhn++WDz7i/4W1myOnNyPcavX8VN
QMEaPSACjkaZgGMYyxXDx31hEwW4kVyHY98GW0l5BqymXx6a+z+tNIHzF1g76eLGIixo5A4K42tR
G7Fin7k0TUIPDcdicgR+thiKeu/R3dk7bSKBCk7OoTp1uR3k56GNiyvAbG7wp/mpP+zt88XhzuLg
pMAYACMa0D+KEv+d3HMoXaBDOlGTfEzyp0Sow8kaQI0R6aT73ej1GZ4ArjZvOobQIIVu49KKoiCm
gkrpD8Vl7890t+2w8bRt6bV/4UtiUDk++NpA6G2m6hMK0K6fq1JPXYZ4NLsKJoVV7YQHcl+KiiTy
R7zREHwa/UyLu79pwxTq0mBEmWYmuHxDee3kKcjxfL1uw1NsIO7THx5IYNJfVOKihpRXN9cf36fF
8tXpzQCTBdi6XHmDpMvRHrG7w18oCIdDC9IrskrqOkguHicxqanX0vhh9gCAqL8l+IKrS/dqmPgD
T27TCyafCb4Md/OqOgw4TycRlfFEX13a1RMKUlgSW9jLsuRdAzOItpo9Cy1X9OgT1F5uvX9ULSCn
t43beTkLUvzT+w2UkEJcfzHiS4/7DcbMnckPPevswtHg8u42zqh8AOpbhregWZtTZ1yZYDutpWie
YKWjEDWe4GY2gf7tnRiSmgAdKocAtFkEDls+iFnakZx/KZTBV5hHlpwL/t4BBZW8LvdJRKCqU4hO
B7mJve0XKeMYkUOGbNZUA864qOthJihapetKjZRKDmA41nTBQXcfAifpOQlWgidT8h+se2l7+xIm
Kqv64QLUIpo+ubi9pRsbfzE/EOZJpq1uEtFphJSrVcPHxZj0j7AgdYTDbVu7jjne2xNYVRBDXka5
awJnzqrxz++BmqTbVz1F51HR2nSjjlEvrMLZAtT38RzbvpRepWgVqJbJeU5hXdJeIpAd1bjesI1c
g3WmdDDV4udY/lFXMhz7q/e9lR4cWJr6S5xSVP2qVd0y/1ip72k6E/bMIwON3KFBk44Nv5byII+E
aqBXuNjgB5PNfOp4yxBEkoJdoi8Z/qkqG0Zp7wwyJb9hLVuZZym8doOZiQl9uMJbhvNhtmErwnv5
b5p6/voBzT3nf+DvBbS9lg3/8vdmxYndL1HhOi07GHKeqraAZKnqvguNmipDz67MOUQBF8zgHB/l
Z6DwTIqrOyF814K5e1QMXpjcKvhFNo85jRqysUivtsyNJxQfBPJnG7+3fK/whxq2dyaqm9C4sGdt
aZ/cIEso/DOMmeWpg8upbTFWMzKHZYgeB4TjxmUfZauPLsieMQ9yF8cr6hrvm7+Al8BiYDUJPQRn
Ra+Hdkr3vEtNhpDAiYudnPEJpJRqa9mYs2egC4XfrSVjE4q91TPmFMLjpUJ3sHiC86F+9g2NAGRW
JFeM8KUji2DU0bTQXxAr4GSswE1Pl5RQzAHqMu2gC5uN34ZBS3XxLDWQ7dcwRUREyRMdIumkTo8E
0ZzLbwwQuqkR4uu7zeFpV79x8KtNZ0YiFGsb5ABMH328eDDMJRVQvV8UnBOgERSdSBQ2dxq8k4en
4BhXxy/yNHH4m1vfDvu2qtZ5vx2igwGEety4409dqrtEDw+Q3qvrAc6E6MYKJx4OOnvqnQBOb8jK
qaXNKt6JoJy7r1M1WveM118SFSk9lNJF8nK5leIqN8nx7vRizVFMyne7tbTuD2Y0/2127PQPH33G
kwx6wB8nVFK/TgFu01eL+vzYv8GgyLAPVD7BW7R/M90ZW3nkYv5njYok6LLse+So/RbOhqMGWWon
DJ5bLG7jMAAkGLbEKBTlSSBmh0fL22fFVsJfPtDGDgjSA8GztJDjsUKL+k1WduleDmWTaYNhgnm6
XHnm7BJgAfuJkOZcZ5iHMONqUC6sb/H1xLJWoo1nXCLNo6WJ7Vuh/3lw+TEDtElkit1dS22TGcxj
h7a2K8+yaEsvYLrC23B5IG/W5hla+yvFWVUdCUJlTBLcg8xUOxLcY0IL+c4Y7/Cxf5qNaqEKdWxP
vv3+/ZOC/tWt+lGTmMCLAKAG83jB8LP8iPphDnGm2wsEMIJqYxr3MucKxFYeH0Q6A9bBCiMry395
q1gd4ZnsKigT6OJEX8AE2wU+Z7QZ5nNKwsw/FXWZC+sYAaVraudc9u+hIzVvamlJu5VqDOBOMsQ7
56j0PEGSc4vsqxfnI9jGJPaK6nwnmxVctXbM/WWKFLkmYg/HkwLAdnAK+2SqBYxgtagoSq1UnI8B
nzQ/ZYc/gyUntQEZWo5sbcT/maa7efPLw7tnhESvujU/qeJ4oVpRonyBImpXnlZnSt6mk6CfCsXy
9xroNO2xZOa9BYVWEf6ZlPcTYpudotNwPOa1zPR/ubynhtDdpmZV/NTvrdpjXQDHAagwZC+fb0yz
9Y6MUiRR0xn5Q0xgBZls3h76ruGEhIkousUXC4wWCvGw5Uwj5IIIsaeSGk6qkge/n+K2hobp/fLE
fhP1yzgNhvyka4YjkYQ7dvAw6EteS9JvWDYVJt4/O29kh6sLuwZ/EjWrbOIV8F0DT6vhOQ3Yx57m
mMnTt+4uZis8FB+k87s3otGz+eWOLo/BZAGW2GGTQ4bgVLY1W4FIfjf+p0qluBNjwOuLEurp35XH
4JbpwUnmVpITNocchH5Wf9cJ7Ppa4/FD+tI93msuZodIQmW/5zWUJgF5FKkYsrEqt5o5R2uZnCtH
YvR1656C5OiOSebuCgTLiuUCWA43pVPSA5osothChcYhBFjr1rDqiKmc86l6v/DkaLwhmnsrjaeo
+bQjkCFAYneeva98Eowp585PH9VYqb+vZQTUsAbGxW7I2GxOOsfC2+LcxGl9Xigg2JzN29rxRS4z
82mnZTGJ6ubbbGduhA9a7kM3Qsion1/extdoGRtTdJY5KSLXXatQuWO5AI5U5ufOSGmdWPPmUjAH
dzVnHR6EH2AEo0xHYLEiKzs6W9eC7wDtQihfPauKUmoZ9e4xmrd9hOngN5DXz3gQWtgemBbNkUcB
2VAukKyZXpdQYg6Tk7SqPaeEvzyNeRd7+jrJJz7tj7Zz1aRg15RLC9vDUu+G3J5VvZLvlEAdSZtc
jMODCLOjHCnhKcN1tpr5Pj0zhT8PNrUMN5cL6XO0GHVc8qpiBUbUqnU48dNvVVikxeHH0JCSKvjA
XMzGP9k5da1xWg6TWYvJM5rM7XAU5uTBr+YJld4YKoBk1xHe90stjmv3SwrO3fBYjqa7WmaJMJBC
uw2uenMeksJVHLMA9SaEvaAvXpx3MNNjbMKMkvkUHUvz+m4W/rd4+G3oNZ85fdK7R9z2zieQFP25
iCT+IdNKVOoFmsV6SyMd5f/P2BSJ0WLyU1XtC2DX2nFmWFFxZhh425vVFhccAvAaHD17ptGIkq3x
cRzYyC0rYpbxV+3Z5XfMQRJlZ2APX/9qOXLyGSs8ugT1xmZzPMRlXZn+mKUWbBOLklu22ol+5CvL
U1yXadRCO5/tB6m8/ICVJGfNKzgHhGIyNnIfSdVYdQkILw2zuK0gvVLQgxvOjjExbvNhsJkaCE+i
HtXwmpsJnqBM+zE9UerUjrITX76eKfRsDKekDg9XUvzMNwuvlBfuBNXUPYnXA5SO74PwnjYId2dZ
vEMYvxwBEEfPkOdp9J2ZnVYSqDs8bp1S84ygUv1iF05SOFoO+2LsWti4vC8KP2MuNMST2uVd7YUM
YvaHNaYeiTQkOA5VeWCWV7WPNM4uAKKndQCGb10nx1dOO3ea4XmKq19ZzMw3bwWncp/1M3WUEkAm
Vkvw5Nlwifp4PqWqpuVT1vSxAJQoxwcpVlDhDXOFUCl60hof+WNYnM9gdaIpy4iuKM2grUupf7u6
LSznJFeI+WSQifConrL2jdNab2tAdng4bHw/0kCkhUfe30Hgp2K22ekmdSjO6RqFbbb+QdNGE2WQ
MUk0V0rhGXDsbpMlrxbs9JJaHhbGraIHKz77EqPaV3tN/8PGMYrAizxJYSjp/Qo+Rh1bmsQWr2vy
MeMBnDsCygBGeuXpTA9h3ATLHQbJXZ1695oKvtp8ETTOZLwVrBUK7twMLyP7lOs9+zcR8Gn+hqlQ
RRs5+x19NSCC/TaxEjYPD3HWmYyiiOh9LujjgzotPmiHKzNXfSr4feow84ne8QDRrAWq55lP2OCj
F8i1o3u6svPWbYdFSx76F1IJeAq+47AR3/4bgGBI1FmtC0aRdGrWQ7Q0mWvKwc1pjL8pVZ391SY4
vEim6XX+ZB6D1VQlYcYcGbTGK/C+XQZb1JHPcXP3nHWamawuhxVMHj8WaJqf9D8LvM1kVPfSLN2+
18LeTrZNPaERCeXdZIRVijMg+OaAsl6gws9XSyyT9eLpUQ0Wd2sMuZWO7/RH9Uln6sGDyNwX8WUk
vZgAV8dFIGi5HAiLsqvSul80CUwQtE5hMHwXFMlFImIWl+nFgNp1JWpZmFM4+1+50uNKDZvJTDB0
ljhKzDureaexqhp6N225bBnl5LB7865R8113XRdnTyMgSYk0yY9YEQqpwgvm8aDXnlVB+HjYBHOW
TkdJI0grzECBA0B25EXh6UAxaTiQs5NpbmDClM4b0vXas16zR3cY+q2EEylDUzQyr5ATqmGbHLU5
/qeA4EV6C5yoGeBDMkJGSM5Zw2YAdgd11YnZ+itWZcpv3pVRPm3QW7cSdyl7j1bHfef82bQe027G
WeoNGysp+mT9Tmviynl5LY1wUSU67xTzgF86gANN4CsSIk8l8HhCo7wD6DmCCtyLdRXSUF4Y9JdY
+OiN92BevEaOMfRp/LofmDjyAIArWcwewCoktuyEb+/BEz0cCAtgu032MdN1r9N5CfmK1EFnOdXZ
liqAGcAZPZX0lS0wEiIdHJPidj6t3Oa32mQORkqgmoAzg0M092WWXaamQqwv2NuPPGyNqS4D0VUM
Hx52OAG5V2258P/nyItpyZVG9PfwCJMbEWZpwW2jiYd1z/F8iAfgqSe3NCxv3wYhhm0bLhd3AGJT
2/dxywBIJGjiqcvOE6jLPBr/9j7C16tKIBDFM7IoDd0pufV4SeERxkZsqlI873sYyZSJ+zGw1sQS
LyGI0UH5utXCzmk1/kFW/8nagnjuTDcXlWFi5mQmQ2lpK7Qmw2wZVh1CDEbuUUWHTTsK5jZdB7rz
CLjNFGMGv567ltUb3N7JBRTN3DW0wtG9tCAwkJ+NkhDjFLk7yEAAguS9Lbzs2dPodbpbYwl274rU
ShHDDXOJ3xP/H6D1DJ7k1qwytZbHpz+3ny3UI8+HGD4FIAaafsg+fwc7i8TnjfgYMtfa9ud3Wrvt
LXZ5vkKIGt3YNc2ZWxjbMV5iJZfq/rhBeG1RXX+08cVQFhLI+oLtkCP7IXbLh9MwzcDHAyfCkpdc
8+u4XuLkmctzPMDR3KEExOCZptNz7k7BLkTTK6W1HmgPYo8SxoEX3lToi7U42cswzt83MuLT0tMj
l2h2YB+hw7z4RamO92Uo+fYeGPV1RegjK/WEEsN48viK0gUn+iz1AtVTva22otcfnTOvOJcWeVMS
rVKKSR6CsmKss61rCLNAT6o9qms8rZJbalX7+JHv7U/pl+LtQ9dFWSxMUqD3nEUhA9+o/q3wAt1Z
VTIN5rLUQ+OZzCo/qIngq6XLHs8TyLd3PGMdLqaapr6WiUpj5L1EM4GimI4iS6xKy+LPEvNR6BsQ
nsKoTohyg/mb7Nu+MBYMwCWNue+E2peNJ2YB5Dj5Pv4csrrpbToIgzB/uGLcICzJVgtO5XHKt10t
OiQJoMaXDAGcwmRWnpyHhYbQmG+OJUCD8x5qfgGSehB/MBcRRycSMb0CBz/wFbDAB7HysqZQC0mk
7bONW+dHjYTG77HlBxwu4m5070PPIJfNSl/BVGJ1WrE06dK4gw82f5eXXs/FLegkCGPd32/reKEQ
feiN74p45wXJHaO+joXnR7vfpcsOtBUC+7nOAoQjplZEOxJzgF2o9Hp09bPftismlO1giYmBEb+E
iTj4qRQjYDlK6WRIQM8/7bKbvANvRf0kC1PyRh2hiaA4TiCFbeOM8B4shtxDc8Q5UckkKYfIaK+S
BTX3sTCNzkXdSor+BA1iygVGQMCdRpB9GaFTF6MPM8EJGtVYcJ5duePPQStLt4wornlPGaWt+bOM
nn92oc5Ab0U1XqtQ0XBqS8a78qbAfVq4EQFGzbUw0+2SxSQ0vEfyQhYL189LRUTGpdwe4IpYOsmL
9O8t7O89EcSZf4K5FKvKlRYIKrJKrkZtPRjXxdU8BnX+qQE3RQFFeT07uKgSf6wP3S8h+xbfAujN
sURCTX9HiQjczQEmEHm2ZamCokN/uoyhxM1gvbO9vBWeajkSOQ0dvDgCVNyzse7207RdOQg98pBS
CiURl2w2VEAa9Z//KlE2ps7tbUfCVJ1AnP0KWYN9ROl1yUd4tvIA80VAHHrktnVdB6P2anMwEd8M
/3fmvDZ6GdKBIhZ4cwmjQtrUORPOrV71s+6adt4W6KDC4Spt356wtLWtPtkdFvnp/htjDojv/pSl
Jfc6TEQyN6DB/9G9BN/LdiKmKuNg27jqh4SA+De9Wzxn7F7lhiScMfqBuhK7gLc76QCxooJP5H6+
tAIBc4Zw3XbgSYuOnOTjD5QLwM5J4Mhq/kiYQDR3pMrBkfuLxzJkmCoHtHo3+M8AEP3UIIpwJScc
S46iBbUOS5w6CpGIMUJVU9jJyMroVLLAZEBwehWl0I7pRcx+D72ETpZ4hZScnr8gx21mz4irub2x
UXPC3AKI7mcHR/ZFdgV4Ds/pSRPpwFoSK0/bIdXQ5jFe3tmZmRAcEnoweLPPsOSvDm0UQPhEJHMY
ks6/43bKDPz7dkpL4xZYCtuPlH9Puj5GC5vR1+tGYFc2leRgN+1iQ6s4EBr1ItrYxtxku/lEIwRD
/J82DcD+2+edW/nddzAa8HvnVaWDh8GpAGw3KUEJks2MPGVD+pgWUyqPsf54rsvUVG5eEA4Qw48i
IArvwo0wiutfUsjVrn/n8LvYvig2v+gc+1+g/a+N1fxy9ijkh3QixXNpF8sTtyP5Ut2kLG+q4MLl
4A8Q8q5v0Z7ghmJ6n3kceiN/yiH948mXiRdP+uy8VaHF57ExhamgI4ZPzoVO7NKf7NvIR9Xbfae9
3eek4QqZ+tDkSvLdakuxdMjrTTkZgEFAkUj0smIRZeEJc1uOk9J/ebycvPzYJv1pELHXNvs8EeTt
d+J4gfJwkUHbKi1hOR1VoA0jb7LIUtXvWIUehswRePeCxm8+Cvs21H2T+MUvPEtqt6Qt03krjVHc
hdpnO/HoD5bAwVurW0jeZ+ryQ/yw2t6u2YMkbBz2I2XWtAdDjdq5R64PjCnDpas5JcT2jvC9j4rd
KAGn2XFwLgJe3ZinJXkN2JCAduyFhEWSpPYHS3Y3uEjblMfZAK3xybgTLmrOC3MyUeX5uulWOgM0
lzz5zK91NKH8YaKjgCgv3oXqwDgSUQ+ucvJqJo9MzNxbLWWJKDEs51hN1BwbhZ4t5Kh+HCwFpp1V
L3ulT3ohAJgzVHrUYNdU7hOutoCGn6w0hn03m7nJUg1QbfS7cidIl4yumsWrgt2byT4fISZLQ6Zg
7EVkcf4wWUzfRbw8RMVpCExVU7kcbbYGPTbff+SvWZ50mbkjtkkheHBh8aIGt4lqoYRNTfXnXFW5
Y248ptFv5gwTSGTyxt3ON3hQjwNZaiPcD+RkFsCAigStHVRRuf+rYgPL8WjRqBNdFuso6zigNogZ
FfrUxABC5z/SHl8hY9VrVyOhdCKeplMQu/LQdcdFXiYeoswQRuwiPfTrvaz9klTmCx6KhHNXVgjm
EVK8eZxbbSLTsPycqwk1HyeXYpLJXOIQ8qxaQlzIAcDwob4G/UzogwXYMISeZyH5GTvJbEOVGNWO
jJA5upUPO4R+mTsWjzAM/i70Q/IBGooVXer8psGgXQBgU9UePcX/2qbWxmsazFWNIV9xX3BPzrKk
F9E103+PcatOnU5acH7fTh0m64dUkWKfCa+e1MQkQhk02hH9QT13+YSqUUOBXJfFtpxVxWBSJ7Eu
AkBjwaKliuMmdYgubwo0nuvv68ag8uCH+NwiJoIuuDEmo3CGdrBP7BEsO1VWQ2WSnn2UMIxQt/R5
1OfDjOrC+Iq1N8pwBpJ4HC5j9gbg1SOMAgB6HC8gFpIsn/rnVJ+wRhozZaDQXcIUkRpPMqJ1IjkC
B6/rhuwGv0tZ9jqdbwBpg7+yqOX2DWpsDMUOERerZxPG31sqyLLqB9gbhqw/mmsFTCHvPeGCPBkG
FRnoxeZMeeLbVlg2inMzjaYxKpjdNscFyvlCGSMK6Ti6i36BSsS2ULQSwkkxbKtJQfxedkEKJ5tf
G6N5dtKAyrkvBbAmOLPa4BfNYHfulPm2rwBUZk4RjpvokIgjBuELvqXet2sjwYQZQaPfbVUSDFM/
f8dcuY/aaLzTAXZYea0cK93tXBaRAwOiA8IakGrflUcXn0e66zLOVVwHXGgXFyhvQq0SirCTS7Kj
g4iwOtWizsEBxTT7sUxfj8iFMh+8N8W9jAysVNly124zCo4yc4G9wovQFE6Gx3e6fPYy0k7goTlO
/t81sCjq8ggJB7EWRY7rJ90Gv3Nvj0Kw0U0rH0To4fb12LAhKYu5Quu8Ng6R1YWDBSMzhjomm28v
cppjUEb3ZSbuKopi4bXc46393ceaduwf2DTQpupHZcl22hH3BO0kTtrX3W6xQ1X6lQHO3RHAqAAm
zPoKnbr0tpFxd4q19LzF8tlrAMNQkPz+P4SUOHdQbFtniUY/BBqumPyFE4lJUHiKO8x1U7e1WbSt
yigNl7JZc7fAln3rmC0U2vxmBRadgBcOm/1F6Hu4s0gmBMt0H5Wa+qtl7VvssK5rT8rx2z9j19Me
8vNDf10riab8cUCgF4hoxaBE+b07KXaLgC4c19xp0PWswqohapG3LaPuWusK32cyZoSxL1XADzwh
VFxwB8vcX2NJGpaTje3USaqvdkzEg0qFTSKDBtsG5keY9PZYBJRHv8RzALUuWs07AnvYaGB2iysc
kdSkQALoh4fjTwgLZk4edAHmIzHvrRYUF0agPwku2wNh5PPljjEzWZuCRVnnwBG5rXRMgDmRk6uI
bHqw5moS+qYHYOKjxWBWyZVgKM7P5ZsXoGLChKnEpo93MwtQz+dqYuuBez/59monDG/SdXwzdHk+
fEs4jlXoLKu9j5Yk1yxmI/t3XCCUgCeoM/l/5m5vb9S4+iaYo0EbojK8qcUeEM6j7wg81UguQ/8C
bnmUFA6No6390ptzBxczJlM2XyMdg6af7TyDspTz//x20pTTUymRL4XNOk4xHRY+Ve7T/WGf2fwW
zk2TI/lFoFLr4f3WBi5b9fhdtqABx2UDIXZWGayZd6cMMmo2pu1T1R+++akqfIPJafi4M3Y/v0wj
H3I5ytoa/stB9h2l3pvGXjo9M7s5755+h23Jw5sL7mio0/REXQyXN5QgFghAKUhskRuQvDLxSrxL
XvjOqkbAnZCK2+WmA5SHZmX5tRBJgomwSB5nxyw2hfPjpGjWGuZLP15Uj1dSuCVxwdRbj0Dz8Aiw
8znEeuNkZoP0+I5NfNd2dtwOWzA16k5mYT0aA9SEn9Sw9xhhN+uSVnGXPaI8Ms7+0/2oLxxIxgEq
XFEUcfcYalBXQftQSnUdD84VkbB41rU0JrKKJNu26w4bpXVCNkgYJtF+TMaY0PtbMa4wilAH6SJU
YX9Gir7TgP9EI/M7txtvLAxfjllaIxVr5VUsxAlTYSyzfztvGwZpr/wH+QFeF7HdByk46KLc0iS1
lZFTzXBR9RarzzsRL9+o+1eYQ+g+3SQSIYJKlV8JNL2pPy40V0HGx3k80j6IN0y6Dj9pWTVrcAr9
gMFQk/MvI3edNnhsNzfO4Xhr0E91pVkAiY6YHDZt1lD4atv8VgAhYqZeELkPzugwW4B3yrjMYRXn
M9jWkwl69XxMMFrihLypK40muD0Uo8qyMEqb/YcDuPiulFyh66KL7UhzULLioebnFEo0WeuDFPA0
XFykMGF11whkC7HViPy8XIH2hEJGRfVno2qaAf5lET5TO7znhrT8fLngQp5jMk+/AkbziyfqeUoK
jGR3wGzrfxLnIf/cGYRJ2BeR8ZFmUJbeIkw2Qp5l7Kxvtj2ksOyfJUwrS44PG3nxI+GMI/oS+ypg
ekrudD2RDiniZGpC38WO0l2Rrc/WNL8JeZ80QbneprbViRWZuIdc3BU7C3zvJq9L5x1Q6Gr8khwq
jI3nGvLtVmlxqJ0Q35pGlhWFTOA0cjWZScm99pSUIOuaboHbRnWeEcsFWNA8jW8Uf3JSefPjVp0/
moUad51lHe+8aNHRGa2U3DjFI9EeTsMnuuaRwkxtjJMhfhKHN7ye6fcZiNJNnIBf9Va4DsZ/Y2qR
0pmiHoQJZ/nvbi1puEj62UndJr2bzrUz9tV4edidc70DqjfEFYbzBvIrlSRpPcokHJaCGmLzoctE
kWmYHlKCpGJg21t0vyTXXCoXaVYf+NSGAUQN8Yt/LH+jFjpX/9mf442Qba7O3zJzi21oc0mblhCz
/RYeCcJ2kDYk8AdWspn2HHz3+QKSVoYcEV3+sYh8RAvrsj+4oUNwI/xvalph3E5nfGqojx3Ouzh4
zOsAXYhNhLYBtzmPkThv0kVUHWoXfqoMtGMnAngT/fYcs5hgghvR2EEjeUP+N+WabnuxcfSJTzWV
dRmbnqgMI8rKTwfbJiOc++k/EFRnY+eTTWMbP2NxAHAtg9yCoZ0KZYIYV3vjZGTJ8pKa5uqdqBpP
sfcFkDbKQdMM8kPMAtLHB4SVATsH1A6XUa9+JQm+hR6x1i6JH3cTSdAbGtB7ApbDc07XAb05JzF5
OVmJSKDz/7ZcD+URv4Fr8uwY1zd6l8TU5TTGgUDU2j01DC3Spc89IelikzDrjVnAkj8CGUx1Ua81
XUFbzcvZtkNq6exLmtjC0p9D+v2FfS/3raLW4n44MdSEgx56ReOFKZYLqGLqDu/2HG3qQEcKpu/S
jN7smC09a7FMhf5E8490I4iTPmrmkpVL/Zwc5r1kNMaCNT0Y9ta2gZoZZXdy9Z6UdVp3/CuIllWn
zdggBQ1i2Xfhv/dzGpbGrFf40GOWHt6XGy5L/OBH7z04d7/g532kCEn4PGE3rhAtjoq4Ft0RXHW3
IZOrYkMsH0BGzgKFMuyYhwczk2LThuk0pXM/jgTisXbAAjgKr2v9lgyCsGhNf7BlkXlZFm2MAXL7
peKQahE8NPc1kai7JKbbzNHHN6+Vs2t77aspjD4y6YngoYbY5k183yGeFCI4My587GHxOJpThfnD
PgKGrXZbJT9Y1j9v/qKuSOP2Xniw/lqyESYF4iNpQv5/wq8Av9GhbvvA25FkUxKDjHM8UddKhVXa
UHtKiRW8ifHad4Roy2ZWtfH0deLKJcdmqkjpx/KxdXrO6RBjSCYjumL1m8haer7R7NAJb/nGy/e8
jNykvfx8KZHfhT+kSY/qzgQA56Z0YZrt2I6O+5oI57dcHQtKRaYh/xFsXwZi0FvNGuv2bv8hwgqr
vqob4NFOFqwjM9tsmy43jNOxA9GYmdrpGLKS4zzl0F8FgujGCF8KbT+q0b3EFLfGQAoQS+YwoYKn
hkoyetiNyATuViorMDJvkluKD4yGka1GGNo4Xy8MFFkClCGecp3vGu9hS0B6tHYrPpZ+TevRpAT4
cdConAumC8EuSnzhiRV5hLE7L2/BHRHw5WRUAAbptLzJ/OMOWV0G+1CnIRHV64JQEvg2vJpuRWpp
Id9TVuYLOYXMxxWLMlm0gU7VmCrS36jQB10+mCKYw97fcME1QECz63dkhaNRl8QPo052vZwkmojY
lklFnZ2ZwxN8hhRTH5DzH+DEfG8v7rgfonlO35SInNlZ/6Dz9vl0510sypkA2Ml2U2LRVOqB7Ks3
SE7aAEGS0CQCysnyyogatRdXBy+mh5FLhCEJpuaRxPgpGwDq8ou5kYLEYB8qWI2cHaAHVsRHhve+
dKWc4B8ESmcnA/9oUGSY4RUk4MdyijM6ge5qiK9ipEu5zbKtSP20HMTMNhhLzSKAZ1fWFz7SWVcb
3DtqM2JSCO10tsfklZ1dHo4bn63ytXg47/CsI5r0haY1ywqZ+SxnmodEALtl9VMk29fFDhG8OgMO
WXBCE2UdwzfV4clTCeWVeBHYVhxLqTv3em0vgLRIc2vOnhBthZQcqyaUgduLqsDQiF0JDCtselpl
s4d8nEfM3lv3BU5xvDBS/onYNk28g6+pQHItkzV6QGdoGjN8mB42WYc+m3WCRPk0g/U6Nfwa1cm9
LRa20oV0f2SjcYfq/kw68S24rSRrIl1jfoD1d1oOAlsQOmV7C+55wfcxW9HyAJFcf7oVzhXPudIX
xY+6/r+jMGeMhoeU5tIA7t4rT7PrQwJpbsR5SjkoFzr4ju2GQKQtsqIA0olHEj2/EO8lbDXEdulx
cTK9KhgkZ9wu68Z1O3j1UQrTPF5Z5eJmZ1t2Tr4Bz3EGpwZ+6+V1/ByHWR6ETbXAmm3izackW4cv
LyoEMc//tO1GtJt08JkkwZO9t2zIpjS09DgMruv7N/NfsJdx2XU+2Un44EC8se1XixjR/3BVW36q
6PZHFhpDOs46Uedjp2jrcAIaCgNn3tzlJlzc28n+0dpYxL7sm0EV/bpL9dALBowFttl09Zozvc/X
iJEYsAns1XncM7n0y91qrea8LzYIheyzFHt9GhAWdHdleT5KdcsTaNrMQUcf9niGIcmErBp4MyiW
5GwM8kXOZGwGIRMfAy5ZClab5CPkIo+dUHjZJZZcqO1mfOiHhAdArguoGNIBM2PHIo2z0WlNRWHj
uku1wtaRZ0LNi9fxUoxRAqHGgvDf1H1AkSO8lXmqeQcAjBdIua/Ros1S87StQfRd/9y7bBtIGtK8
7LjJydhlPMWi8YXW52hPR9G/yXpoheoidxuwnPPlG1XXDe7lDWQ9YK8Zn2jMp/FkmX7s87ivW8f6
BA+9podEoVDdxRMSpidQhKYxnFn6OOuE4fwPIOhVKxJrGyhhRtKkfxQfryjpb9snzrDthQCKUemz
MNKQXvJSLeTWLhGkhbV2qRqAbaV4x+UfecTHUtP2GR0G1gLCW9YJ6T2PDotkUjAT4nyoNFQso8SR
n/kEDBtgZVnFPSam4+FX7fwBgZwIJwrenAqo5Td8M6dT4L9fq/w8jy8yS5DuIgw5cPKzqEpWfw1J
KckaNkiQ0w9IR1p7Z7lbcFpqSjLF0AExGSoD7QZbshdJflkqYOxUbBrCos9sCCVuLdi2rPIbQna0
VPAwqqe7vOIksXf9IKbdH4K93txZHM+aqWTaL37INxBjeWvN2uku6NJeo2DCfZ4YUpLaTjhfRq5K
e35hgGvSfpIwMbhmqW4V6Pxz1Lyz+5UuFxsr6cXMWP/fQSdWyGwbaSHVeRL6dmu+gYiMAwK+CwIv
ZgKpkz8bIEIYYhQhsA/jegSCMnQe/QWMHVMU6mSnkn/wOAplYS+rB/jHpgStwgcsE2v9tZ79y9dE
/pjmlPgyYceDQT8aRQIhQUNc7qBd8Oc7BJzpSAEI2t31sLv4uPocZ8fkVLZwVIaMnfJ4LD9D9O10
B42GfHasC6o+xWfPid7QOM9KkirGQYz1E+7pZtwU2Wa/6S6dMoeDMZ6Kx1tz4qV23X9MZ7dqC5BJ
FtAiOlFWNgLB03krzvL0MMMB3rNFQpRZ4cN5MczJpB264b4T7aTOeOWxov6q6HLLHOPMDxRnXSn5
UmrSJIx4EizYt6psVWLIBiOWfPz65eOwSt0beUd5dXTcXo3Gbh4rQ1N++VW7TleJeY4aPqltWxET
ZKTswpKM0Dw9c2X1i5vKgEIkq41u5rVxa38RSEeuFWaUhqOCJEGrxbDEkpQf2ThxAyFbD2v62gUF
rc8opX2BfyXcOcYqbA+H+gI9gvYh5+aAsEpSX3L8n4siReiY60oEWxc1T25wBaGM85m4lOLjaY8j
TJd+OZG5nTwgvxul1eLx/81u2NSkleIXXOoN1inve1a+h/2DgGXiBpjxgk8S3NaR+V93GA6I1kAa
oY1nUj3bwN7qYo3wpDYAvUam5s48MdFJ7tiC42s4Oo6mn2vi1UuYPXHolTlKOwFkhCwV9qrnRDhQ
AFARQGMD66NGvAhIr8BsATR/aXfXVIyBIBns5TMTOrCaVEwJC7yqp+S0ycE1s/hT3iaI5bMpj+VF
92TIKrWeJiFwI5UMd4HvcB7z7/s1PJBUcAqm2NOloBQFEdDOT7/rAX91ZQ+ZgHEI1dN0pB4BdKxq
PqYnC52PIMXZ1f8Bm29DDq6U4XrUmDlmgUl8MI+MCnp8Ktpay3EsCvEQsv9qnKO1x93MJJUdPO1Q
3wPdNvmTguNKW4bqpwqjiWKFBhKiBeGyc8M/4KEorp6ArrDpUpbKfEDA7+6xFs3uIQefSufHCBEd
nc0jGJoBaEyiAls/OCyxuX2e3rH5oX1unlVTPkPM2Y7AhAfIli5H/m9dbC+9ikU1Zi+iFo1HtlMK
wITPB0X9p44ssVKfqsLTtcF3X3oLq+WWbn72A/K5w9CrHXuuY7Z4/E/KrBJMAClY0/73xIatLeop
DS6WPCozqsb51Py+R/rzQYeE+fbHGl0Ml0F7//gNAGDeWfTimKvTODidAtf+FeMf4RcOVtWbKGGT
eXtA1kOhhZZTwZennMrr8X8aDWpgb9NTHQSubHkb9GaPKdMwyKBQYdFe23tenRG/L9pWLrilyADx
30Ay703VTecIqNAPLwmdFg5wmnpW4T74f3SN+eXnjYgy3afjGCEeJy082ZsNfjTSy8V+tSZ8xjKw
/nJ2m/tBmMl6tXKkOXI9Ju4b+lzDgl82pWSZ+OhnSvjMzGzfg6TB8brrglFDhR5Kf/vsQB22D84n
ZDhtBn9MSTvSSVuDLWjBQkMM7gUr0fVMTHhVEnco8ZXFaVbJtDIyze9VOzW1GCaYPuBVIoCtgA3V
WtKiByc9OlUi19tE/F3Mq7GNzeHGGisEDpIrDV2v17sHFNxiZ9B+0qr+muHCjPnWidJ/yoCcMJLF
IJ0ca4PSBCpzkRBHt/L74az/r6puORTzU3qpwl5u4+vClAUYdUhkTms3OwUeJQ1jIqeoZzg+aOo/
z82u6Ags+U44oKrza0CEBZvgNCB/SsJuNQFekLfBukOZRZUKqVaWU/h7o3Y0EZiQorYzg0NV0pt8
77HdyJuyIOYD7F0cLBWYzQB9O85tO0zo4p4OsPs2iL0AnYEbRTVrPd32hRbknmdpI4H70VtFkVmX
qqGFmhYGInB+sNMoIeLJY43hxUGMigQvdYkjt+HjYeII9iqnv6lyNlhcXvAG1hT9xvlvfvyw9Qj1
V89KQKsXmFMPlMvTViplhG+QcvcT+lb9NdQghON09FpfhiIvy1m7QSd7UCCAbdDym3jAv+GVFxK5
J4+mEC5y4eb5WObptHzUIyBIlb5j52JJjunAbq6V6ZPs3EopXU5d84H0aXwfHKa+0V6E7V1yYzcB
vaZpvWi/SjGbjIprBdYXKcSRBIODX3lyKM0MqufJP/wshI0LXihVXLJXcs9P2uMgTYKV78Yfj+QK
csUim9TQsGpBkRM46+HQUDCWoqAugV+41Rg8e6Hxry+52Ka6va2tDkNYxa+PFceGyMVqyAF+Y6Uo
8uJWSjNBedE1P9vJV7bqjepoMGMAIfY41zZIhvb7y+AfaedEj55gEcPRu4HWgjy2/3qeSUAvaT8p
a/Y0u5M4JoHc8ScS05Wf/SvZn9JDKJD8J+DFjItOnTVFGvwoFLmi0R4w+H3XnYZNZOqzEITnzm6t
53kBYooe7/38fYHKTGADWH0Zunh0K6t5cSnRNWF0KuhsMi7ZP8NnrC9rrFo53Kxd1q2felSolsIb
pjpR/3HD2Ky7ytsobtG11LQLl4tDwuDiCHBx9B+nh6OsaE8dPx39b1DZUYIvfFqgt9Cnn1OTlf6c
fEU5vkmakSK28i05IFlDQZ+EIGkV8mbw+gvZdvrMfM8fJo+plnoDZ9pR2do4Bt0KNrmp6oefJ1ju
o4fdljWz4o8QXwUyVqSo95bitZBduhu//bJVl5huJOu4XgdjNasnLpoq4Ew/GyYg8LK3OCV/VyCz
wiPAZdJ7m7C4jjQdVru8LMafyAIBiV3M81SaQDQWK5j7H8/elNoviBC4WciRbR0BH1heefA+t3Al
YfoidmSaAIVXDeRbLnmximJD+GD91FbILA/mlWy1Tkwnwqla68vZeoZdSZObtIqnu7SioMN2Rmwt
nTMlDpIWnm9/w5LiiJlt5mrVWB8MicsBLz+UmwuxS1G/dyDN3PsuCwbpqwOfL0XyzJtMKBZvyxb4
LAsht6i3Jlv602i72tDUuVjb/ICnptVokkuiGeDd1w1IIbmhfWu466bZksMVLflGdEGDpMyibycW
q9VwqSKn417a4pcaVIRFxneFO6KqzDYGP3blWbcSA3XLxp3/eGJGxN546QCkoM6p0ufa6dG2WoHt
TqwDwfTfWy7vEGvN746KLfiLRHZgpY1Rw/Sm/qXTCfSzHXWXiCSSLSDos4kwz2ji9P831ZKJX9+G
QIx5D2F1igtiL9W+Gmhjll9HAYyFPmXpF2dUpnKaoIBlybgjb/tHjygoWlJA1DXn/pb+dp7Tf5k0
Dh+BkUwrlF+mqBFmIi6Uzz7vx48z9tT7FoXZBtknVcOWh59iQcHzAd8HjPpWOBaryoug3IchiXCu
9Lrk1hzpY5otbmMNMevllXabLDUYtXmV0oyHDmA7zxlBj6kYnuTETdU2aHnKZr0nutttEHBLednL
/vhUANCzGBySRdlDgNFN7Pd4ya8pliutCxkvyeWQ+beafSum1wu3VilUKijRcAn7nNTu9BD1a1jG
4mIhR+IXVEev0IA6SktKnpfh31DWTGcyWpHNhUK7YL0p+oIouWSFqw1VJmDJOakc5aOOtBIxr+7f
VyWoBI66myaDO17X8gHB0rIOrO64EbjPiQWBwQDQhk5v53AEOPMLm80OyZZUiHr1LArSwEnMQBbn
dSuKdto6CkuZMwqbzlvitCUtntmcjJY7yXs1EMGsr4XDTXauxWMphxsipvuFPnxDvzAt+61VELZB
Q4CJggxWQXkokudXa0m+bAOfaPJUeqiwbTx7B4+luGzGIpM2DIdL4moJXgI+xfOvLIPIXgvKn727
wE0c/b79lnLhL8amlmse+wj29C/xWsaDiAmgD6nwd/vn17N2gnp2Vi0067CVpQDGLdArxf8TxzJu
/Tjjh2JeMtcRMMF5aXfVCDxyuZ5hSjxJdGJClntC3zBMK/Hjtpzl0HV2zWso5CkLyh6oqb/FgvzL
C1E6SjeDY0aUWHELBzRTwhehqPpwabH95al3ydjLiGQ6YAA4pXliaLxCn1WUNOzABE6L7cYY1Aav
sprQLJtlWogu7WiKmNYBjam+BAAgPsf9ElMHiPYCicDsBsL9L2kmIaZ3sWl91At2RYp3g+6adVQl
dTYMvl3pAB+0tLmOV5IIJig16shhnFXMkrD2EemfzDUX2ylAC2itOZtQXbz53XNhGg125iGJojv1
AKLPlDO30lB2GeNVtVys8rYt3t9CaO5ipXhpCYQt2NF10Tx2fm+0mWGkSknmHeO/UgNJtSqH0FfZ
ES/q4cBsUIV+agCa2OR0YmkqOt30YfgVTbsea+p8LoWakSrLFlKYgUWW3YogyCIrzSLsyDe5kWY6
Q8JJzK4Gzxcj8PCMrzhfs/U8aZ2+cOunpwqQiZvVUqW2qim60YIrIAMN9emY3kxztN5vosj7QffM
lB2B3h6mSIWyefrzJAxJNIKo2XARR9Lqql2O2P4q2khDgCDnBr0bABXes4ixK8krMjz9gv3EwqeQ
xCOHiQYO8SNgs9/NdfkrFtowMTB8IXdsgIa5aDtFeP4vIupi+H8++r7el4AEygWp92cfUJCC/mw4
GPA3Fo14DWbEaw0GfQCRRXFyT3JdIbzJpuz4G7lfbJJKzNb4Wet1ZlBOmBtfLUi2TokxGhgw/2Wp
OITUrAzddTAgSeJexJeofoGU34yOWn7hKgx/xOrw2LBw6kKgiOrv74xnQkcHdw2hILH3TNjM2yJf
z3EoHyCU4fEYeosJIfkqiwVa7qJ0L5U0/dSurwKcxCx79ziqdtVQhiGvfLM7il7NbpEz5AG+ho+B
kmDOc9C5rNIqVkI2+DvYLYNgFA9lvWyZDdCxIUEUjt6tDld+8RcOzKK2plWu4nNVrtzahoL68vF0
RWs9uB0EId6OO4ptmX7UzscDwxgRN2tOxrMhn4v1cIDbQSKuQhwmj41hVo/+/558T7Z0L2Arsk87
JY3YKTGScFhaMect0utGf4ddy6MEL3hV7GxpnbCVOAJue/qZACftQI0XUMpgsksIgDJvRIiAs7Mg
3blggdtvJHYneMk6rawydeQ1PBBl2BpV16zm4ptkiVA8spDX6fXbx/QdSofEPDoiijTcYCIP8syq
ttFFOiDe/2rl6zT7Dlo2vJvCPTMaErO8xuet6fLtU94+DQUwhxSDs7Z3EvMpP8t+mwi4r5UIGDkW
zE5HQLPiAES7Jv2M7UGWunI7HZ2AmRgOVtj3BVsg4E5EtMVBUhXDLy8XJrDhRs6BaGZgcutw37St
GDWrT5wWYS4FQiIeNrh3OTub2ANUrTvc19Jwmnd87bzG/pMRqLb+4vBZfFTLZlWKqtCVWqqLiZbS
+LDi4ELQaCH7yWOpYYF+Sh9vO9Izpm4ZogsEadlYtZnmrGnsd/i7rfyviFR/26DVHL2LGakyoFX2
9/JF1CvHGDd0sLlYtIsU08ukycfmhSZ7XqCmm8pAMjlTRiv8vY7y9CC9TaFpD06gts7lsyDZznZ6
qAf2aXcgnvxcM6FfSgOBlenSzGxY4Jx/qI5HJbzGhUImlYRx1YSnnlDTM9obZjED8qRMVQvrFTDB
pgeWn8QRzbVPK4B53z+p6TMyMKlyBhuTk6XFTN7AkhdOBsU07xhmIwGd01xE9yDBvBj+MG+cvH2Q
fUgT3X7VBuiVdErNGRvSLiNw8ShrSiM9RM8aJQUoLYbGzOIs1JChfU3wVPr3doE2MjBpbpzkm1ph
egkAMLWR8rvTEOvzNoCcM6I8Y2ADZ/SHVmBOZIjs2Ev1ksm+uAgFz0e/O6xa5DyY2xZXRVKXif2m
dpZYHsz6FtymEQfYjKY3jL5FL9D3slfvMW96eiC7madbCcAra2iANQw8GPQVS+tL+EF14yBCsJsf
Dw0rHU1gy8mUmfYBXq6EgmT2q66Q+/gJL0XqWm+C9J44aUGpf47d1nbMlCJp9TR8S2xrfb93+skg
8MVIFinJTSM+EVTQTZHHYNjDEfnYc5CUpDZd8RR16TDGoYzJl16Pc6N/V3Q+ldHtcGCUpKgXcPZH
8RaXB80MSC9ZBs5BLVQcn1YuRJgVxTDE83F1Zj83jFTXx0/iTvA4gKsVx68r0AcwjjcfN5+MMdn9
iym+bMqb5STrh//gdbzOcswlU9rDzwioioF3I8Blh3VCKAPVUslzE9knqm30A4qy0uP/cSNffOJ+
gAVNESKAK9HF3ZLNa+nlNiYTy/0DCCBZddXH8I8LT5ryNPA2uzEt0OvLpgPynOzoeMuPY9IFAzCq
a2gIwdDzOQdPLe4+scmvqrib39VTt4hjLsHTJIX35b0WVSkBz4nGAjioeirzexsPrUQaIvZsOAGl
K9jboXYp8QhVvbpVjDYnk0CX+l1bm416VCEN3vbN1CexwxSMCU7Ye5wyDPCUbtjCxxXw/OeXM+zD
S66yKbdt9NKRRDLDvt/UQdmc3EhBdjQH6TjmiouEwBHYO1++kPkhttmmVV3Gjpz8IvD0Is29GkkH
1qllOd8bpdfNrNLaKtU5QnyBp77TvEPkmVrA7q0DmG1sqHy6kP9J/uZLOddcMb7KZyCvxy002lmp
/8drqzj1bjE4jtqs9NBOgy46SUFWxgi9NX7Wk9ZBKSGaI/+Y1I249fVLqZb7uOVISYo6jOubr9WX
lSFa92IiVC+ZiPHpVJQJebaGUyOfpXAAWhgpCX74NOqLb5r00ysC3T/HiyA03JyUhOY170DilHt/
p04YLMpoklcQVjtrdDnEXLWQvny2JFsnqAPJM043Ha6qUhz406aSzcrU4Rc3yxr8XODZJizlKMl3
FHShgIcstnFu+yIjqSDhrQPZ9RM/sG4Cv4sJyHiSTzb5qBJyDeM0otXZRkyeQloDnJjBL0o833++
SiS2Vom33OqFj2m8Xqmbwfse9UfCOT6OgVN/tRIVDEhnCODlyWZaCLssr3m4Xgs1syEsogkSjKPa
lzb00x3vkxDlUWMfa3vyj5Xco3FSyp4JuuFvvusMtZQHhTOt0QsqSZxYll30Bjqu3kDBhrpTKqIP
3VjYm7MJLkSYelBvqQYrabaMusb1/ZnabGLs8zXzySEZthXukI+g8IgrVN+NRPS0Q6MJUOH66hQo
nSrioCBxfDV/o/ZAWBUO5Ipz2ACzqe+iMi/uN+6qadvrLrP+dRBYY8SJxpkrl2ET4Ao7mSHNE9sN
/3x2oyym5wGxaTgDufDy1pB5ZYiTMe6AoUBZd3KbwEzHOPMWSzNwzn/fef5aemkYsa+m11AZ5U10
l/VLgHJplnDrQfeEQ1D3rhtl0z33mSbsnEMqfYbBq3hvQOgru5iglIBaiqEH4WtKHv2CoqeUmKer
IbMXtGyXQ8htXoOvL56jNkskehOZ78TJ7terwvlrjU/OthiEZPqivosl0ao04Jnlf4l4n513khIR
ci98mIocLTBKA27Mwsf89b4r9z4+mxWCXJM3PWbGkI/eeJEWEizPbqU1OwndYgplrTWmdrCXcRvT
GBhH1Jn6ZqJ6/Ly15ehjzQtKcib02MSUpFwsi3CVX4HOlDIP41IWUU9g6qlHJqckM5fXKMH+vYNO
kN3HuM9lspQott9O6quqqrxzW1S7nt442YXOvzruEyGFyp0vSwvxLdMdLKkx4bngUjDbnUTL2/9N
6HEw20HiLBl9JcF3arafwSv9A59b6XRHVyWt8cca64+HHsdVNFJkgux4HgHJidS9pSH9vh17dnG0
iqI1heG0YCFi4l9k8Jy1iwsBDZPBmby7O4VzFztqteuKoSnOb78PjPm8PzlPGr6LbnL+w6i9OcE8
A6L8uLIZBaAIXBswLdd4cZlU1Axm9e1rLZyb7U5De9XjxIBHlDDKjcWNYaPOZWZOBUfmjv33KFYB
2LglKJGkM0JGnRSyDP6ETQnAKqLPYuIjWKQwmYA0X5NLQVNypegOqITkPkd/YslXiAd3YLTDC9U6
84qvdLPc3XifEMRFuztci3pPUGcYpXyx5ubd1fkBi5vSmDdFWqpCGa5HvlX69h4rKp1wHEzhY7ZE
2h58CiczQAq0/cDoTKOKRZ0vGl70pxB7nNQ0dR/yFRvgn79cHHMwG9JsSelA3RI4LEKjUZBdex4b
tInzLPYt0GCG5tvCJoJdGKmA8YWHE+ASNNQNA5F4pYr805MoRKpmkw+VFHHB9YXSqaQB803ptvG8
hq+ZDVSZFYRa9axgta+vIWQkeeO0vSTL2SmmjjkSi+dT6W0910++qsbm3M7npPfaE4Af+ATaUkRg
vHLlVxJZOyWjcQu0ak/cZfpNNc/HmAiB3X6N11NQiTrItai4niXvKkLyHCgig/drTDMWIP/Oxjqv
o0pqs7LpFg6q0q/IU5sNBui6rEb62Trk4U4YicwcNm+oaXu7pK2eb8acA6LexV23sHdszsPyIVM3
AIBZdBZYYczBNMoy0qzqC9YSE4as7x1flCCtw6bCD+gPcueetNZUTWh/TjZdEJvsMyM/pWneQ2zt
AAjSxR2bs/8cQqmwTWf0dRExc/xgTKrcDf1pLwYahjRiLggKB4ONj8m9xWmewBBuijf6HV8ErQiJ
NkJUV8s1guoOetjgq0djLNXZRQF4/kDMDdPLX3FQj546KXzzkUdsFrrnaXHYjj/lypGNLOhrbvNc
M2WsUf97Lv32YliBTUcHWnKgjsfeKIjlESp3+OdINOlib+UwrFeLQGIa1y2fnjgPwca0l3NvGgGs
AC02Y8VCP99H1pDaMWH0ScdOoF3LhyIn2W0MvzvMOuATm6elghzI1BivF9P8/UAZBzXICcFzd+7k
Ja4Hswr86ph2CkxGIdT5+W8Kth8hK6nke59HYECrCpN1Fn0IYBNE3TD4NMT7x0Vfyp8YHGBD7czF
bgf6W8smJWeJNW1B5RK5RZiXgq1frL7jBZwnRSfykn1NlqnS/Iec7rFTUuoDRBUFbWPOaNFahAAO
f+VEfiYS9sUf6q48pqxfbbxQjetyYjvPvtwK2lRfCFClUUgzkzIswAII5zPhqVSrSPYq258uLBXe
Pc9fUpkMwN5JFEVPgVHJcWe5QaZTjTSrjaz81lBkO1ie+YOLQeKfcqm0LFYHTb34T5depZw5PWfX
PNCz1/9S9P2cryLPPLsHj2bq77PCh068rwxfnBHJhTlpciFQ6WkJDffESzQ16B0PvLMbsRGf2zDZ
Sn0yhnCOBOUKybOIr08Bg1cjoKYZa+3IyIyOL3vMXycJ6lxEzzI16OHKOBcoPOJ6INfE/nAuO52v
1T3lXZuW7Jkg+TOprbrN+/PBb7RD+Hz3BQg6FA4YH5tN5E0A09xxRn5OeigmAdCZNZogCfy4ivaC
t8Le2FU6M8v7wpyF1HQWIN7ryH+L8Cu1uyyT0SYvIOl7u/CAH3eTFDJHhyu+f4xYLZBCTaUYNHhc
+fpAPCo33wAjZNj+gLHpW11NC/cIhsTXl/jUawSYZL+sF0CBeChGuDArzucBZz7xq+fwsb/Mnpc=
`pragma protect end_protected
