// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:15 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qd/W4fpoy+V+goqkbFnlPdOgYyhWSsgG3tBV/b3npbLCUCe1V8BVsrSydjzm3raC
/60H30vIInCg6wqRzcewez5uQqVvBHoDRGkJd9PeaLxewMdqdYE/PynlnR6BPKWB
f/G1Brpl8V+BAhcuWb6VIIUihCh6k3mAyMuDPaw/TQI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7472)
dToxVw+Juby9+EhUJiieBSBP2jdv4+keopAIPNu5O50kqfzuN/S7GPVuw0hGhPeM
u0+PvqUWn++d5jrOnVSZ1BchhXQiXkDBdIvqkGMF1N0PJhQRkzF64SLwEKh7AM3r
rAABhNTZ42doB0uDAXov10KsiUbsgRVeoterOfC5DrYSS7MzMqci8/7UnBDcoaKK
qc08Xm+Dz4waLCry8xKovmyY+HvcAcbYwk0asG/4Qfuj16e06hYsNmT/O9xDIMG7
q+QpoVzWvIuclbvAcfFQhF88Kwjt8+v87CsKKiDYRRe9EpgxgsgvMysjmh4ebAdp
AeufiF5qBqvmNRpXMEJryFdm1Y5ynNuCy6KkYxVNnQ/Hwd+CejhNXPHCGS62Rxxx
TpzIwFkT/HAuvZoX8WtBmK80QsBaD7ZQoaoTlsVg01vkz5nEyJqUoX+/aWvXl++t
oG2ri60hdOqL9KiPG6L0jBlZtKTpr41R6UIe4hrq0sehhX49P2sBNbeol9lxGerf
p1b2oRwXB7nnqVG4eDurHy7IIVXPOCx3lqdn8c28MEebP1xTaLT1q8aMMoaHWXqu
n3zfhx5fenCO4S7bUwpPXWpKUfvwUl/ApJ0npXWoqS/Mg29fsi7cZbUwfekLmAzF
iLwCU0QStMhxKoCsKxh3wJPyxpzCTwvqXvhNv8n6/6ANNhpxs1LpGPi7BG82D4o/
5z35VZjTycdpDwc+81WjcYkYIjafRBP5XXAIC+l4Yy6/ma57h/jcVyv2uffthX3x
x7NrE5WirXdanazgasT3zww5ox5ok3sDzD5ufIg4oPi3hpIgEIYj8aZtGvXGQU5h
EL6iUr9A62zHKBU8+HP8roYwqnQsL+sRB7dOSDSYVZtfhFYU77HdiAmiS6l//vGs
9zCwUDDYSynJNsowkPTBqROEe7vxFOj9xehbe2d9w129F9toRGQZqPWs0Fc4T7lu
/m5D6XXTwVOs6ohMlcv9pYNs9Sbx05VTvZ6lMtp6Bo+/5KKWm3EIjbQo8OivFlPh
II0LRrc/cTXUi/ujeZY0OPBXpIAk7yvDkueA+L4aRjGN4OqAg5sON/5mdLinw9ZC
QKP3kPGj1Bx1mA4dgytJ/6rWTpTj1th1hLLUEWE5Yqaqr0TPDpa2bzwrFZ00RT1b
+md5Ip+mMvxpj25mU/P2BqzlPWos+p+I3wjk2uwr9hUA+WH18cpUiuv3GAmpzlZU
/pmXyFMCmNfz6XLfH24fbpGkFAMXhOWvY3V3WoK45/bP1s47+tyumOrwqQV3PmyG
srPKJd3sVwAcCH6Sdhtm1KaFzhV0OdObCFZ5A5D/OKNVAbV43YLJRDo5l+6thz6F
xPERjlUxxyBq8CxOW4irEH1iZ4lgc/udkf6afsm2CBT327cWjxvqSOWldhOq9Mu2
6KmHOkQTwahHLKFtOyi9A7uy/6+DB6xkzNEkdQkyvX7SSpHUS93m/xUGVwTCc5+8
peZWrUsshNWz5Z/jg5ZQfb/VACL+0cSfofZI8BWH7k/xrNicbip74cWrvJlr+r9s
+pcQqzirf3tursrB02HKdYQQU62wpQCi1J7cyqPAlsemgKrbKkAu9A346TaUSxcu
j6ihU4nM+dqBoL++7gK+rAFYroaRhIWHHx8OtUCgy08kqf6iw/nZ0qtLV75r8J4d
vxjzfnKZR8L42tHEfp2O9pjBOzKpZ7fOcB7TcSUpU7YkkJbXA2XSRCKmWgy5jlJq
hgz/QcsGI5L42A0CGTp2SDzDWYH2ZWXN6C5PknYnZaWLnLt1AWz+ODdttpHrXmk7
hw6ogaEKLZNuoYffrSVjhdmVHCynXL7E3rmi4XnmqbfDgTgUIIg9A1QLEEVvCzYQ
NvGrmJOuzTapZi3PKRomLhg2MwYmTkRotiSBKNAyX4ionrOx24/ue5F13EwM1xhs
1F6QFwoD01fpYa/3Nstid/7n+bJJrIY+aq9H0Cnfxu0WQElX/9cXSSXY4t4R3wxD
kX75OiPiZTPo55/J3jjCWyotyqb9K2coeU358EsLjvx4Ma8ZrpgPsBedQz5xRErO
zMLTYrQlaYTM7AUnSZ66ZdxUpt+WMDkJOcrIE/xJ0JgQqxffzqaqbWjZyPh71oof
XVfcG/bmYJMeDDb+5KwcueSBc3gMRzRE1GsNXnnW05BbZWPQVFBjP1mDWJdMSxCH
ixsAsU+hsYg/0joGPS8zAjxMfrVINJ7Y0WW1TMTaLpzAl2lP1eR+BVlyNELTNCcG
bB1lRH5T9yg8fwiC9Ptb0mcexwpUa/Dp+WJAZVohm6XzWs+RO5MrLK2UREIAkoK5
0Cg0aaC4IGnCRtW+ebUXuRYB8octPVLur0QFBR8wdvEydzH5byHC+JnGYF7EVC98
SUdyy6sZpP5eEI67ycN2KDzU2j943eWjr1Dn1MDJaPKtvSGtuT2MaZ2T+RN0iT07
4vXXGFumj/bOFVqu/2UMl59Nowo1iMePi/5CLXvM10FywOyIDbvp2Qc8jGHkZR4P
aWdfurE1gmsiPMca1XiLMS3LnsYJpSq9abmyU+408Z0ZhX3Y3E/nbeCtp6O+j7aT
3Gd+bUnoJEvKluzXRMTSVF66v4s2+GX6EEzAyDEJIoDDTDDbsmLf/tw5O6RsaerY
hzHMZVHzu6/GauhgJPMH9HUqSiJPCXDFNnXR+olEyE6WZFBbGd6a1RBXRn8Rq3yJ
g3+RsKnMfC48GBc1SZxQaqXrJB8nDmuXfU5ylMCPN1yl7u0F0NvZo/inoqs8LqHV
2RU7VyYN3GNuuT518LDSHCcNLzsWu1xm2FB41+QXPP/nu3uQhUX+jT2W+jDVXLP/
sqAT5wvLw5o4F6rf+hHrQsqdqMz+FuxQDtd2b+mw2Y4gobzdxSz1Pl55WRQmZ+KD
9gIrD+LvWhMrNj7sJN8oUIIUiooCP4r54EXW2rie45RyMGaodZl38lfPCPdj9pQX
CVHmoIl76XHPs2vomrlwsz3KPyjhtQRV21STts+CJRGW1T2YtbXtriSsy5nYasSI
SHwFKuo4zbOgC04YZZSmGfnvgtByoRZj2mlnBk3yKKQtthdRHaQEEgCjFScQIxKm
cc1M2Cg+q/sVK8BS5c4YLe08sCLzQo1sSzvj43LEaYj3SKBCy0f1T8xOhX8P3YQX
zPAN7Q9foeSqlaqLLDn/PjxXHdsRl5fCd14q+6g+ynFNm0XlH227DQ9jqpgyfVJ4
ggWw7MiLs2mc58ffTJ1PqlIkjswMBY1FtNbChT7+Y5pMeqmK5jPV/bOQ84j/LENi
ioo0XA/AB7j4jZxKnhIDoOYmQXXozGj6lPZwfsvM9nFEORShZGOSjAUipbWLuyhR
Ks3RJchtnFRe2uxrV0vAxonX3DSSnUfvDwJtrysZ0kBfRs1tBbuQnFlKISvelTVx
JJQGP4RQdZSgRUNaV+IFc8vEq/4y1IrM2Gm6BpWsQ5jwup8RC2hz5/AfXsycOThi
wfALhT8auHnWOHJiTQfW8BV5BW3lR3JA8oILN1dWvZyEs/tyj1qG5o4ENSyQF6Rn
aDiZcQyI6DslJMCVI9XllKbUZ7WOj1OXbHMkaMqHhmh2sHqEGHBrQr+vHFXpKDfq
kkLbqqHCCry/5RTZAZMHG2SQd6n6xnodTzx3R6PS49HgyJoF4QYwsLalZg52NmGf
J0H4dJJL8vktj3ibrvsCgJ1xO/o4uyEqIaz8XPpqu5wlXpdnW4BK/wVA3xJ25zns
yTqA4tC80i3VtolTfQ4X/bWbkMLhVl/2HM8K/zeiSLJzKuRkhTuZGyZPXPfRjplU
F2eOusqzWDS3cgpiIAPtpV8L5yLs1YtK5Ms8iJYiOFUE5VaRusR3RV54qcxwJwl9
CjjKKukz/Z0hpAUagcOproo7b2fW+LVAQIzTbOXeK0JNjn3uc5AEKcMyEColiUur
pN7Wfeda8sRH+9HT76eSqQNlm5DsR2fYJx0wNASqzARBRu14DKxUhGhSg43TUKK0
wx6KrrpkEXU8jXz8lD6G8c81/iW1e1f0E304/d1WoXXrXMoaFhmaQx1Hmm9ZoTG3
jEJEviqWB5SLZ/z+vvnR4GUKXtdCY+E/Moi+ApUHKd3zCd+CDCbzojM3NzHPpHBH
mUqnFNm5eQlaXHxkMivEUuBPdG09x1cabdkPDe3/OxNZx6G7ERhbbAVBh1MhnQZ8
QE0uQ438yjRo5mD8hEcSsATysSS76eyz9GuIh6+JiqLCUsRmm4j6wVBV6uz9q3Im
dhz+27GHOGSVJVSQ9iEOQPoYGRVXECRyy16VigdE4FiI8Ag5PohfCs93TUe3urD9
kVArTKnXZlhEG8HrjEhZlz4R3IrSgYpwQ3llotMo19WhFPMBK5zEDoSbiACggEIN
5RXrVVFFYwrJf3LHKmunoDfkwbudauB0adVxIkP+wAmqGBLCR+qfDednue1u2l7O
fVP1A26B6Ipj7Gs/1yc9JcRwXMboPTKF9AsAdr8asblIYbOw1F96vo5+zwaq62K3
YXEQ9IwDL74vvd59MzE8klDwKqVZsyN8AoIPgL0HkkkobsjKylMlZh0yI53YSqFc
Ruym6azuVMrWuVg+E90LRsjSwWm6uWOtWOCSQsgOadYdf18ljMRDrzb7dfee2PsJ
7KrbmXRgMnd757NtYyJxkceJ7sOHBpiSejNwUOKCHlZcKGRRWtipftIckb43WbCD
Qqz/aPkw3l70vLQLCUaHS2WmHy6iblvDHCFjRm6CKDz3AMOzTr3L6+nhvZIV9o0+
TkrSc5zFihJT4nQXNj9TFebYkTvO1ayZr/ecCbPqZ6Kq/mbJI/S8FWcq3uOYyi9/
OizcGldLFZvR8fxky7SSiDO6hFjWzxMvO3qiEzFoOS94OIDpJZAMjknevuWA/8Dq
+oNrCeyOVdmODbgbmnszcpzISsi8eaqzQ2o/SPPbxA93Hs8ANcUrvbrYrDIaWYpA
Jy18ShemaJtcZ4RUi1VR7qQfc14HY3PGOQ+r5jibwJG0r/DL986uFfkeN/fE76We
xr6nZXQvPfEtg0/A1YH4aA1PxqH2C0UR4QsQ+9QJY9FtSBRzHralIYefvWoC7AE/
OW46MG6p+fQpgEIhtuDaB9ig7kazR4qzrKt5z3m3XZGrGFXcqSeV3V4r88FMBb+Q
tcZdCAH2rth6keCDQ0J+vFXX09KKN2x/09rMCOqgpkvUBuHEKVrB69YC25HGBYDs
asAVSfOk58Wm1eokEYdGATx6ysytiq3qisFcj1JaJpJgOWmbCAy/vr49VOhhHmaA
p/oZ8ky+TH7ImDIMVa4yD6xyYUhvvT5kKEL5mkElll0NciOCgrKwb44MFjSkkK2y
zrZxVu706z3IvZV0pCBDO1Vi/CBoIT7XayId7U+SiIktS4UDgMlJiT7efkSxsemW
pCVjAgXQzTIqI+hB5KIiU6nvLeR2z1qbbv0J6A9kT+gciCfav7YrimpnoafM9E31
3CeCnxWnYRNCjpFTnZomsnhxPjHVoG1pXRWO5UW93wVrFKlsNHnYKxInV+dqRciJ
IMX/mmG2fidgimP3aJhzIW8OZxlLwtziC2DcBpTRoUgubMkRLbfQB1MG36JPqH0V
FME4mJrMjiQGNdxuYEcQzpUo4Q86kvGmWZFu89wSFPozNgtRxhEHEKw9oFs7XTmh
p2MfBnz+B0iXbm1SpjjnSRNGvZtQDZJMbOXwqD7sciQzTJt2R/ISls8srMJolV27
59kvUL1T6VW8mu1OCibGwhhvwY0Ig6lUVELLaOVM9VAuDDPt1djF4QQVtMlyXIZ1
bVxmcQzMr3RO6hrJHIgw+1UjNip2AwJrYW2eQZvDO3Fdp2s+d9t+yNKBeglKPoI4
fE0SjGmxPX3aQbRiGlvE74d4I1mAbg7J5098GUR9YOJBrPyxeVtAH73ib/p/3Oz5
HOiPOzp9RlEewJeUdyOXNqvEe6/pP2XaVR1DResVHHVguipg5F28OhbKVfCwHCha
tBmxL48vssLmtmcJGG9i5Gx7U+mBS8CsRGbHMMA5XWJUqhEj/enLIxCsDTrAa7KL
H8vSmHQtj2pzk5TbP9guQaHv8YqgGGWusKKrPvduKngIXsavOnSMFWdJREnunzDW
pyb46RZv66K6XPOyF35A/plk4LP6Zw923g01F58bsNUOxHHKmdsS3Gv15ze7wNU9
BnMLeOChYYtQvDJwzacdHfuP8AjJxKJi9EogZSk+81/WjaI91Hfgh1U+yMtxXCcb
Jws9mRK5fAIQ4NA4E6tCAiQGLg+brwOCD53ZJ1MWz68+IpLgZQ/i8P3sQKBmv8eJ
dL5ehsctpL4/CA0+Dd41SDSAk6e8AUE4k3o1pK4LB3eCp9XFmD9JW3EVDh4lKnTY
tAik8oRQMsL4z+91VztfbViX5kdw+b755wPx96OJui+Ylf9XW5C4gRl5wXuuF3NV
KDEguP3BlvXGxSp0slcyQNLWnJFAq7wVFFEvgYpgmf/z+fvn89qw/+sAwUvxqj6d
Ic2qQYH7JPjWLAwqqPMJ6LPbzEROb9s1GX3GcCJtuE9ZSCh8sNZqliLKO4X9FO/w
IHhQtaCNNoGeeSSI/41v/mtDoas4fb/fJTyVOigPgVKUx92SPtRwxE7NI+Zq8Y3y
0PkiKi0ByI0XXerdM9q34Y9WqV69oY0lRxwLCYH0m7+RXj0xMrnsIwS/YISPqLkS
E/mxMOuj3jpBzjYQiPXBGqJKeikvcMUdI2FESnwt6kSUO+AU6sWQahzS9J50HHx2
ouIvxNPpDht83xFlPTDFKWWdaX8l3SmezZibotHpxJiX/IUNFm2oyT44xfoQj83I
wOmbgqYmpnVa5oTG/0Nxc4DBECuDGVJR/TRTNCZx4rD1eZ2m0znEDWsnQuWAIr+D
Pnecm9ktv8Ss2ym0MlsSsmDl/ixZ8VLQUjx+O2Cq4yF+26FENB7Pru1Wm5lkcgjT
tCgzcvS8qQNFpOtY4Q9Ip60j/d2qynhh6OUNBYCg6MevvZwqQe+h4n+MYGIBquzS
tZ10ZYjuNqfUsHolI8aIC1H4cueEV3oVkSrHYMKk8BN6CiAQ1nb+WnWDrIxnlZL2
7zrQzppXtTs1W62IJCAu2cFpN0ae35dlaFe5lsWksTSYw4WEWjr44GL4Rhs6gmxA
eceitQg0z0akUXI8PYoZyZgpOE/iZk4VH3IF2IbdmmpfDcw6algLfxUyEMaMia95
C9N7KhnS/iePCSSYbuEeWUIGUpPk6ED8TUPQtBh/1oSd3GbacOmTWbFwpIBgGS37
EZ70uC5tgglE/l5lHmi1TkLrlgg8xfJSBMOkFHEKHTTk+rgr3/MqONWeH/6Oe0Q7
Od7VnUlXCByUqIh6xi9yjiw+QUee3wxWpRIsC5UR2RAbRfBczQoRm2iqJjcqjt5A
Xcohiyd13OXBUd1KaXmsXUWvqucgGj01QLpW2DZHm5UqKIqX9zWDSq1FF02t5sv3
ziBBT3Ks5hlIeM29CBuRdJAp7kY0JgMFGhrxAv0HVCO9F8BLEJLhR6TOo4QC8ZWS
st85jc+XiluKxnSUCnkC/q44G1HWnEiqAHzvZdlcE6A1yxD7QtHmo2SwVdJFPahi
/liRQYp7Uck6KQaxY6/47l2nghTUv+jX+9GZhzVOoW886N1W7XbYuSnApL9rThfp
n/SDBGCO4+ZpnPymF4al8PU1wE05cZ1VFx0ln3aEr8L5K5YFYxyY3PQhIo9RlDOG
rg4Ndf5hcvB0n5K63UNKl5GaeSavT3dXMySd/SAi17slIxk2LZIaBNC5iBI0g0XQ
ZtP4Jg7W1hE0sLK1xbT3I2NppdO4SkLWcBBZ4qcqG+CA/9XuR4zGqC1uvuF0HS1P
ClT5w8oeOgVT37/S9lv/Q2RmpT8nhL06pGevkd8CYTdxKFpbxLM8/E8rAUBEx0Vx
u4umq/N/AhuKlgynXYLwYxnnhfGopT4qqL9llL5ahJmQOr+Sq6bkKgQ7oG6dOcSE
DSIHASz4tcR6seTPCoEBduJIwQQxOK2/ok/2yVWvbiFCrHmTiKbvPbWjbthXq0mz
XdggYpqg8irjOjfQ67agtLucOsOPFTt23xTSODcGl9yZ6oKYsOigXsLHvyQQhWRa
mC0IdZ0PlDhGiaL9SfW0onuCpgukA/VdCFj4SGehtiOBiPAa9CuxTKifxSqBj437
mFlALcTKgBMykr+XPqjy/MO18xdUD7AEp4fw1PfLTft0pyW1w81gy61Hy0uFnMQU
mH1qgE7U/24+HA5vDJEDVxg2vMF+vpir67WzeX2irnA6vN/Od/HL37XzXS0rjJfT
L0p2xLQZK1rc9LnoXTvD8odXst/ZbOCRmlkFiIxfwqW6cJ25gjmWOzuoklLc8eBG
I4ypZlHbJfphg9K9W/eub/dyI3o6WSrFSxfffwt10cL07yNZ79cZFe735cqQUVSt
vcwYwKedXKuQuekC2RVGYNb3c4RzqlD9acPrEN4JSfZhpRWj3j7RFoCPPfwi9FE9
DAUXyQLFXjn9NMdsQdSAKowNzqcqsMwfXy+S9Hg6aZbBlLaz/911hEovTJfWhB6A
BPXpModmMKVHX0OFni2Akz2GzkIeilET3zGUmlGPVzm94FoH2+FeymYWTOQiE/6c
3JUx7AjUSvVXbtc6H23uRyVIwzly6uFoZ8TZMp0l7TvKPKxibXSi5sJQ6JGcFs7q
TThtCZbvpmhqDGcT+UmYt77V0RPocJtOSc6kFOVPDKSW7izngAICJGSfZnnkzbV3
R2sDfX6+TrCGBwmRcOQVg3F0zBsqyJNbqxDaCHF3wBm6E+gnYdnZrZVhbsn+4V+9
k+6yorwMmkIYzCQi12IBAaQnfY4n8J2VHvtMRKmlxCaaJU91nb7PBaLOF5PCykue
ksgqlrG16s0ciCcrxWSqR/58wwcl6zYgamlsGkJ8Mg/lKq3c/fTYvglyhtD7o3Dr
k8/6dWiZXMe5GF+XSiKKgCUZwxhiFE28oal5lRXRcVkAFVsgq9V4kfRuvAbzjBYI
YyoQse3juLgWar3j6Xdh3iDQ6c0TnQ5DvVHLmMQyw611xpItkRek+DLUNqPALZGE
RCyeoyJZ8A+EN+Mq1m7BoFVCqEae+roD206aolioL+TbGe4v3r67eWx49NEBkkkl
C4gywb6NKFreCf+x+E7GBlkBdVJgW6K71Qhqtj58VmHmLp8afThaSF2nWXqMujL6
zP/tlN331+ei5kYsKhfBsIFaCUafjHgeN/UZ/UScHhLQODyHUGvMisaygg+HT77e
O+Dkz8ljRz5jdkbBu41oQclTNP2HVFY8nNMnQyGPhoulxxUB7yC+TeJlR8qok146
vp+hLa9c3oF+QzmOGqmfnY2CCKZDDgp0Xm1S+Y0aksbNgDoxYVd0uH2WvEaL/GfC
V4SJkFZcsVP3d7IrWge4MU1TsX4n3m9Y48pbKLI+xUEJ1up2YVYhdCahDHuGJwcI
Y4upOWX8aPjMH1INEg+rH4YkmOe7NKp9br25Szbr6ZJ2tm3u5h8z/DHceQIbssGK
MNsDXPebx/Dab+cSddOFBksqnH2GzTT8Vxg3EVjFyUEWui1LeRc8SkiaNvOK9+/Q
EDM9UZoXFLJ0mSNIXKDAyg32C1bmkMAmNdO5Wl/xIqyF4lrS2PQxj4d4wi8aJD5Q
0PQxBKjp222dJ0o4N9D9lb3JuuTPZxwxuW8EC0BQA1yP5gXeEYhtnJWlGwwDFS7f
ATBMI53owxoP/pKRHKpgtIftujP4kACaiwVdFoFbz88mZSIO7/BhGLnHTVSnOMd1
TL5K9OXF5b+go9P3U78BRwEqXg1rmohAq7zLRDy5XGmznipeOCWlOqDxAh28sUl5
PWyBK9GnqDrXgbK86D1dsY/LIf0w9I/1FEnkTQO0N1DYbejsyjftTQzhG8SQD1S6
WBJ2/z5u8gezXZ66Ce4txq/At4YG8NOo2sUEi8MYDqyXUNt5uUj46HpiMIP/ZS6w
AMM6F1XMxHWtyvsJUiZHsZiFXC3RnzoHrifwKs+siJ4=
`pragma protect end_protected
