// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:12 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Rx6wBC1IheHd+5wBEqA4/ibSYggFIs3P2ubb3TExw+2T7DU3zvGp0X+Sas0edykS
cep8aeyRaDYL3mPmWNsF/uEYr/ITwaEYkoXotSS1/H3OPO3k4W42+oJmmqBYfQW5
MJZ9lXvfxIkQUvOWWZ5SONCvMbNlVFXRZp1exNlnSjM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3152)
w1FTwMHMWJfzzp5j2Fbtxe+n1o5VTlS3C7D42UyFzYWwr/kRWDXtjgEifXujOed3
J48AiDT5Ea6Y3pT4CJiEcRivuHxm4YGe7fa+9ibRZPyDBnoWwFmr3tyqLu2qZ33L
jMQAF/xlkAJ6hqtTv65VzjYzZ/vdD6NcdbgCjWRFHqH4tqxBBjX8VTAXqJfy5syw
CRdpOQ1e2LPE9xEB7E27FdvtMLHzFCQXEh0LuW5+5NmC12MwfU2FY+tVGAYCuE6v
GAdSVzzFHhaGZ2I8p6BZnbipUCZZyBDtJi+yHsvqwOUfLOjOKiA1FgJMBoMtaTvF
s2BL6EmxULi+bOsV/P1ghspJ2VlMoyKk9NQYABnpMMSkM4Z2W0+ULGZBUJu7Z3Fl
x+8TYDsTxT7bvKMtQFS0VWZsztNM2bCqo0L2BqgIqCRrNyWpNWVTHTW7nX68ot3O
jpreMN+A2UUAtPYxPFV7L9aNUftJNaWjKEnreNWV7LLuNb/OE1xmFIjyz99qThqC
fjXbHxegn/iG9EOT6Eirt9ndersBPi4LtRwBIzHyR4NaTU8X+/ZTrZMTyBKUBsDn
/G1J2SjP3WfZTx97Kn+bloDq55j/3jlVITAVqDPYTOYak8vQd99VFKisM2fyKHGo
SrsbxNGDK22crva1p3+hWseWQJL3nQIWnrwknVGzsNK9b4CrshaKePwSl1VJ3WZE
voCSPZaRAEXiF3Dxqbt0iI0D1NPZE+ZOVzI9YMKD2Sch6w2F0fooBv0T60tcejGz
e5aNoisasD0FWS59bG8h6lmDQCLaYmXVYnvNFraK+QLM0FPp+h8n6cy60E5JENmD
o0yw4SgEplnj9nqyPARR4DvWyGhDijhMnb9dU8YEJ6myyHY/8X07fT+rLQEOF+kk
WWYEp0QuCvQvhVM7hFxxgJHEW86Qa050sUpX/x6DoFUBDw5Z8JgEfrPRVwmCfKcQ
vOI6cRJk65crjRuPCEHO7gWjJXNfoT7QXM9AES048bXOt0KZy126ZwcqGK93yEG/
gzqDpM2TzFSd9znu4zBImg9jxzslyPqSzScmBKZ2t5hvr8DPwF9Z3AozjFQNgVDw
864m/yD0x98A8/soRSHfOMqq/gjTt4P1fibFqRaBALosBvNzAgQ1aZP6olSfG9Jn
h2lGjbZCQ1ABCuBpzCtSt96cjBybDOPTXAMmr3eYAEFq8g0f7PaS5vn+GEP434yD
1E67AiXFGR3rJGSrLUTK7luwztuqhMJm5g6rWOMBBYUVNT0iKmrij/Mkl0JM/s4t
MVksWezhyxhmyJbGHXsG+tRUuAo/e0jIWMeU0jBmAcaWxS9GFO26HPLGFujMXt9U
VfH0Ajd+3Uw9BRal0qjX+PDW8cTpW685y8Yw+7Uc2WuXufsCIfuQUHEG+WJxTnAA
n1iEEnr/ynU//CzQC9mrgsPi8AT/Un+z2LoKKwdYw33SfBtvUWIkKfc387auHKC6
nvcPT7bJGhealfmDL0mTfnzxkVLGn2nDVVud2lGO5lAycZu3F3Jsf9C95gmDjDM8
IyYOtQGWgT0CXsPCSkq/Zjxx1bG76+SCeCESIa8/vMZwFGa0rQ+NXEasAnPJHHJy
B1jL7CFQXPlVMKXaIcRBGiJP+ibc45VEG4QHbGLD1kUdEKDAZ3grO3VYjikZ/5Xr
qa69Td/1KfDqwN8tNyTNLLMHKthriU+nsXrflJvMKY5suHksPKCpTJkfF6gofhDW
+pzrqXV1aep+pn11be6I3hScGCPnjsSvAAQUQl+GbBHdK3l+c+eKtBTWeUYEPByE
dKVYOUAzr/7CnO4uQBEo11PwXrWcu6eHRR4HbX1Ie4JcqrvprfY7VaA3d/LUco6I
5dyY3tQvZEFiUkJeoH5VsizbFEqw+49Wju4ziYzf2Di90xDEHE+py4yCevxGJ1Ba
zEQaypLTQ/Qpbbzsm3myykgLNEGrBgXWMnxaerPmqFm+A2k990Pn/yG7YcjVIS20
/GOG23TZLQE6zuoXKXfHlE4E9ONF5D1vitGW4jSjSRDCApPBIzg7jd5dl6nI74QZ
k4leyDfZkFh2OZOHvv5eKJiFigPdC2Jckb0Z7al1pdMbPeuGdCPzw9Dszn+PobNH
STOdeN3UWeCVjci5fELZGlYRbR3REOUbg4+ENwm+EHapZHfOsV1wUYetgVVye0P6
GI6NgDUxo5mXss1LWswn98785/mz0bvXZtDpkc302nxFV+mLFzo7OvLbpFZzWfmG
Kjo2bVj2RvQfuroyop20tIsc6AXNQ/xdLHx/9OAsYGZqCtJM1nPw4sLmfrTNoLDF
WdvDYjBhdMccBW+VAERxmBB4XgiBtnqM9fWh/GlfPr1VV+Aqz2SiFC/tLq1JXH+Q
Y3+92AdTrFvKcPGhiMQn37tygRYhT8REfZkSNReBBI94L44Fk6waUYF/Ig5JbAg5
apbQvamh5IS8vu57DdApOfx0wskDFmtplFdmXS8086ovUm7Xmgcu4wMHhROFo1o4
PIxo8EnmUL2s9B4UwZLrT1qBn2Xh5UIjNf8l9WlCVv2QOC9HZ2T+LXoag0MUZg59
4IZKoTFCBEqIX9yG1T6HPvvUlJUfqXSwfMQw5srKvtNWsdKtTi8OkjKDxGfM5vdj
RpWlcPk0kTnKkzLqK1wUi3NaXwGEf3psRDRjjKgORbyONODW8wFZKRyDr+kuhXUd
aO4hxx4zJp1mWTes26QlvjlqefzK2Jyex5cwX6dqkmrYejRLWaAYgxR8bVA06Iay
oUVAwuP98znW7IPNDLmLScV3/k69ZDqhNAx/nD0TWVGMUXFvemBHar9Pp629Imt0
w2em+E+2ZfS4D0SbhWu+82TdJCPh1QpXwWe6dfz6eK6DbgI+GxOI0bXI29+UUaY9
tL7Dd4YIh80YHctbbEQYLMw+Aq58F3P3PVMlCOdSwwHoukBQotzbvkkvTkiDX1/b
7VKCXQrCi1vQm2wqOD+ZBhpK0MAcDRJ3TIHLRXuUwFexT4lDnIyxnH6TFfueO+R6
X5doz+qmwizFEXeo8knlzJgy72Oz0XGs+TCbgDppuvZSu39JUl8BnwwuUNypFw6c
hb50u/35mwOxKSs3qODBU6q62euFLWQDMms1opetWfVGeAR4VYUAjxcghZ/NgShF
e7lqFlqOyJ1CyecORSo4VSPezn7e4KpwKvDpHm3SBdmn/kTify4xNcoIKP/sKD6r
dG+Xbg9Z/YZd/Ij/uXd76pVNO8xjxPa49Hy2h1//jaJW1zCxzBW4+DUpDZox3FSZ
cev4KnZprjGRDXXGeGzlRctS31KT5LthHPHYYy07hDE0laaPP+5ajSbwERcc51bJ
TpqJ4FrqVAfZl3vngmET68Dl1o02VbHUu3g7NWz/1uRF/OcKNLSfHeJPkRKGumuZ
IgmHwJULwVOB1JhMyJsmzQqA+X1N7fY1L+QTUKklfiqciBcErkozNpD25H+zW+ci
GD0u/ITuP+r7KBypAZWM9A7fEa+dXJ5wXKyyhNCKSIyNOan4H3mlmI1gjbjyiSmc
xE9fVMmZ3hz2aLTeZ4XNgFpE6hn9yVpcAvVOa2wRXUjgTwiJJFgtZGCJECTqz4RE
/I1e28uQS05KTbqabS8QZPU5NGZCGFVbIrG7ecuZ5QWN3R1kdv5roJ1nlPoHB2OX
/KetNZyQC+54gGICyLkFunSNQW7cplbHuEso9Rew/seSQpa3RT8/m4joJ5hT+c17
bTxQWoOYiWoe2RaTgH/bgQcwQEsXCS+YaKPgMJ5MBUxLGhMGTxRO1b5Ehx7NaaP9
KI3vtnsIivnKpXZEw4j3jygRQmY3loERRCW/awRp48fT/NfRqCs4svBKZTmlvE/s
E5GKPCmeIXcs8xAPudxqcU/GBFIq/rMA7y6VIB8FTx/n6sV7hzvXi+R14optA8E/
H5b7XNWanCmdRL6MP8TmlKfLPWs0Yjfw91h5rbzDm//OsAH1nmSiDPuiomw2qCPX
MpKELrsCIFfWzKUbFd+koNvNmxmGmT6LKnwbZ9deZcAKhT+8vi2pHM+FXOGnA2qe
RL+xoFNC+jebJnFchuPJqmVW7UR1zb+r3yJZnfnX3LzqknaKhN8rOKcjOdycr25c
taA5+XrweG3shcuMfoSt/OqM+/A2PC0vljvgzIuN8RdHSa9DeSoWEFTJdhF/tR9S
XAd7iex6F9RZnnsk53TEDF6bdVn4Xec1eiJ9FD7fmmk=
`pragma protect end_protected
