// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
CmeL3DVyDHKni0i/pIxsI7obumCtbVfT6wQFo8a6Wvw2sa09+gJzRRofgbJ5uRgKEWqnj6MYI6PD
3aR2wUd+6w+gsLTbYAH5gRCePXQ2abnlC58iTzkRhMYT++w+jN8TPOAzp8WoSYzuutSlZVobi3To
4fIoA9cJ5AwJn23tPMOktVMKKt1HzrlQnqnGYalv0UKY73h57hcqT3Hj4DB44/rT9larlU9C21lA
YsmWuszFdiqt7i2NAGMMi6RBoxNXOLghJTTylk0SncNyegxOiu/ezoJ48hBO9fhidn/23LUjUwp9
NyyxtwHeZWvaEc7OzqaAzIqHg8vmrzm7awVAtw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
FCYw/LY1U9QhkZEi7FePI2ZYU3kgkBmcH2uqppAp0Syvfts1EHByPR/cgW4nAFkn+HtpKUYmk2ul
pNyaQfQ+XrEs4HzUj2sjMeMbK8m8R0OvrdC7ottZWAATKH0D5n4fvaopw7o2vzDJFjILVpTLx6hl
r8IhVMEaWsRw22h1ij9gKcyR83Ubw7EDWtcpN25LIQbT4OXpxESbTW0M51lLAeF320F7q92gkPtg
EfqfVNgi877cCg028qhMwz8yhb6crccnXYd3VRdvFwc8m0tIAT3kLpUoQTN1MbwAPq1CJ77pAN9T
WSL+n7fIiahhNtqNx04GHDoBHNclJuE/uiWhAoXJLeYKZ0UfLae9Hr3xXUd6gJQAm9qaUOGM/8c4
LbPvT45diXQxqfPFyrIFjqBMGXMbMCKTeLI2ftOcPd/D8g4mEt4ZrGaF/8Sws+Kv0hk7nLY//05M
Goaw2ktR2uL+/x464vmSK7vrrwqkMwMH5WJ4CHgVWbZmRJPhrXLtQD61eYjJ1GVfF5K/ESkRsZyt
sn4+hBqInmmtFNNyT5oJgUJSCZFzvELVwtiDMoThAfpeIVe3HlLmBzuD+RZgQ5t0BIrdpKMLdwcs
lvEs2rHxERRdYUWsx8lCPtQQO9OeRXWVI92opSFr5R3UIG1UwgcPKJtg+w4V50e0oFj7lZCVkbrF
RcQR1Srf2DkiWwRRMNngPJMMUTADL5w56gH23MQtE22YMBYMzerKtXeHYtcNRDa3ASctTbCjR0m3
uMxeqnGZo0EFHBCXM1OAMsQJe2CYPBjWHcJ317Q/TANyTnYjZqax7tfxLaJPNR66tKhB10rQO5dz
YLaImVtUC8HTb97PCDWEo6eHKJeJeyq1OeSbSYo5usbpnyNgt+7FYyIBmNeFNPvgheZqXu+IxWh/
hi8+2P0yLNty8nd7NWXVEjrG7wqt6gP3rkAwBVpZZ0dqdwSluojbXQVU889XktT4C4XDE7Qp/hIK
3oKOryYgrAK0IBd0zMuxCocl31eXlrzfuKsLBSNTwOPirFBSBWq9cSGTv7HUIfo6X+8GRSyOqcD7
22+OcdbFPjeqCt/GceZeF/fZgsZdFGRaj7a0KUxjuhfF6sKGm1t71GS/d2kKbDKSFBGXguyjYFBo
IBCT24T636GuZYyqEEcXW0H+IzfGWhELZHmB+7/xjkjk5Osf0mIxfVTFcWSIx5wrOmQTk/uuru1j
zU8LPuwPiaVpIp2dUF8FEJPCnrRZbPNvODQJxbTdOGK5gPY4pecewjP37rxN2iaiZzJCiiVlzj39
biLsQJZHvgyrSx+9OZVj6WqaoFQOTMKE0CFZFnuB9yzau2jOtUsgFbDFMtwovBPyYHvAQFtUM24c
BIiQSRd11DehxmvLfTLyGz7cPcqELDr/tIszfUZYJJC4x+xCE0Idhek3ChwmF1SJL7nWlWAS9wXQ
oTTd8DAlm5kIlqb+VHvBDW/XrOVnnddx0OMLEYRb7fglNSVtZci2ZbQCwx6EwJFQIU91mw/DIsv8
0i9Rb3b9pkr9NdWwaPNRsyic9JwblnZ4d7K3qAXaH6ib569OqgkItm57elLF5Gu1MC0Ixz9gb6Mi
poNL5nZ3fLvDoIMvKhwQ5wZdxDndeNTg7PKYluSOJMOPhpYbn0qe6QsrdoLD1NIzqWkA78RzJg/m
R76ilw+bKakrzCwfWmpyoiG1r8UFoWjZSCQqde5s5Mxh9y1vFkdbdOdWzUyIPJrdh9omNpVGu/Ak
Ixj5Zyq12DWCiu4YYvNTX6xliyMGeHQpS8FSOsH9v2088Kk2ZNJs5qOZBd5te740y0qAhm9Envdi
LbQM6EMV098crZE0jkI6etNtBQ23DkusLj3clZyJ8ROWJieG53HyuY0UHO1D/9QF+CGKAGl+apw8
5uWLirnfk5msF36zAQV+QZOQJ+njras/9I6HHg/yMbkONzN4blbT/j3uFhJbibf01glFpmS4k1ja
dAXI+4v01yNOt8I2CtafI0cvGI0gGTgzgkh51xumZ1CP3n/iPscotij6Bn4hQNAXdEssq4Jgx0X5
UkNvQ7+BPoChEMbWH2VQo2xqm1Eux1WW/LaEmm5LKkB5sZb3CHKsqqGVHk77nB0uVaXmnUE+ujUi
DckoY3lblGbos5eO1XVqmsgJWwGbrN02t2oixt5gFz5vhX763welCPO5mwX0n3saj0hysi8OJJoX
ovqoDrcJRfrJGgUQ43vt9TK5WiwqeQZx2YAIjtcDqBHExsFY+EGOgpkuu4SHYDa86Nq+SnNAvVzs
k6mbVRXXUvwe4xm2SkzZ9Ln999Y8Os2n/y5YvtLDtKLORm3rgQMhhjJOpeulvVVHma7+cZzWXBD7
FgKYiFAogpExhX0uKRzdX6lNMUsUfQ0kRoRYyRg6etbZetzJgGPApsDq2Rg0d49qHYe9jeOBcXu8
DZFEqoriI+mMbm5pswMm6RdMJ7kwcRfX2RT4PD5FsAlRVOz0mPuGs765JICjpxBHC4t8izbLTZJ6
AWpXDqOB0p1QB4fPcRQm+czJFb7/k2FL24wHqp0kRqZqMm/iWIx6cPQDi11JBfrvyP5UQW3xpP6a
H7PR8QJFGrMaZlnZxaMjP2fugMQT++mhOPqaPmBhhgdln+IoF/L+MHx4fNvCWdyz2+VwjcP/eqg2
moHefcHFJcwSpLr/hB9Y+jQHJwTVvUWbf6n0tNzqJwUkcUCMYKs4CBjZeANqfG2lgnsQGl9n1xPt
15g9k6Op1JUsAZaeDzYssqFtLoveaTqChOMO8KdPnC/p7c6LgdWSrcam9qsZkipFXV/LstDKgSrX
395PhOQ2Icewp2YisY+P6/cHmztaP1rvcwTf6xMkIvZ0AEenlxUjz+cOpzQINW+0nZsWggIdpmun
8WF9Els6wgDKDKS+zmo98tv4+rWnt/ELj+fVHrW7mR3MX05OOMkbX7iDuPDXx8LrU0sc8symhI2q
aD19gQfazEzl1KFAqe9AYuNACptTPoEUZ+nGdl6sIGCMI7XCq6QfZOcbjkOHKfkHORzSoKgFNS4W
gxJZGduM7ALERj7cAvhhwQyjf0XVYltetqjda6r98gh+Q5n7CSzjvi3V/tpZqcg5RBQJxTncI5YI
6/SvcDlq0IcxtiwbjqL8DJyFCP+dU9OesgKv8TfXM2guL0Y1p4qo60Cedmd4xSQ4oC/XQOYqomY5
8KoorsNIFjD6WGkKT6YJuIUGI20I9enjP0LD0eQnK3VeTvLhqFTuo9EiA1drOBGslr9dudBynQxC
qv+GcS+n7OpJT6DljLdcF2KoFS2uO8vD8n8juoja49YxlfLeJVLWN+MWjDCSMCi3mXdX/yaa/XDp
aFULavsxVXXMGHxpavlOTeiNLPQ2szXB3kB1Mi0eaUP0iSL5mIWJptqsCl8ocpb3t2gT9kHkmStK
G0enWFt3bfohYANT2qbyYaPZF/16kau4D1ev/FX83ECO7Uhp1wWiMcnXypE919QA1PcLgAkghGG3
MuGeesRDzPv8QfRtwOTg0rArdGPyXjFaMzIl7H2RbMI62kvQKTjnKfiO4cKe4uNda8+C85mQFb2V
PnjWB5IEvaPnTTVErSymxwOD7ZbIkh3SNDJELkqGMUmRD9dMvWxSbUKUFIzibPhjdZRWCqhE74VK
pbLhOafzd1f6hBIOukA6cIt3HxVsZuWLTP9Dxv5lGR13DGpXpXcbPZcqmK7Ts56j+Q0ilXFTdyGe
TKgXK56F3DadiF177gvMqBvb/zXH/2FyqRiRWX4cG+SpGTAAs0R00IeVtzxtPeLywD7/nZC/s2pw
iWUVyoOlBWLlEIM2zc3TGH0BpXohAMp5/ZDZD3xWzqTDujqp3fCtSV+ZSJhcQS06mR8vbnLY6YQg
TV59/bp0vcJV0ZyIdZDirgmll2L3J+iNv5OZUpdcCSNE91uJ0M7FBTM/FoFbw5WYbuNq3eGui1of
NBb0dgWBiovTY2bFu95wSeqzudarGUq+21Ktt2d9h4BZouzs3hL3C4mhWHMPL62uliWaN9U6cJlA
BjrK0Oc/zBI/6u3Y66sBp7uACb7kfD/9auO/OkWJOgEqH49eecPESegW8i8yCSvPuSUwMy0ecur8
Tw/P77hGeIGernvshCZrH2ttrc4MNJmCqlaa8w20NLpSJjcPwG3LjxcK9Vzl7lI3gAvqW4TcxOb5
y0w26qeh4mdSZHDzSz+8kZeSWnLTqH1uuRdqIhU7J8Btg5P6tLv9LDZd0agBQqfMuJus7+Vx3DZ6
jvIjZcXpooJVBaDyNDKse8ADBpT0uHqe23G7sSA9RmsiKiifIVwzAwNwTilvIooPUSm76HGg2Bj4
HNeDfZHxPpRwL7/3nkG5Uzvki+qLkGRltS6RKDeG2UUUUmBRyDgwjpYqspnZd5BMenkDgmGTAFzZ
OYjDXAYWbgSrX+Xzh+RyGU07oW8LuSAVme8mZmAWuKSgl+0VVZPU85dHij1n4tq5Zch0ShpYYXd8
e36rA9xErtX0Ordp6towJM1m+b5BlI0AA1Ja+Gh3saGMSUPNSvDzPGh9bGG2vJlPD48NnR5OWJTc
oCZrhcW6dfLkQmGVuD5LVXXFhKQVLuKSmpDN/OWIEPmnHPrZBcLq+tesbhzp5T9PIeWiY2DdMnZ2
a1hrAacgv7LtnXC4LXAWZ5+/Rn3PpDfM93ddE6vQydax7kqMViz+oCMk73Q1lJaspjLXzyfd2TvH
650o3m16eGjsj6ELs7S/+O3JgfGnNNQytbmVdYI9BXks8y3HtD4x+Uyec/xSWfjhZo/T7mXcSqHJ
bw3sRQC0jQciOMKrHQNRhr4Kx0icrqip4IFV7CSeUdY1zl1Q5t+ngGCCosr0i50o5YWxjErq3m0B
stPHTuX6g81YV9wYHg9IWHXWRSiyMCkqOhQ4OmlQ7u+2Wj7da/QXi7QCIU66tdh5AVD35Yes2TYH
shvvwKaAEdAIaBSLVz7TKdlb3tvsezuY5Prv+mlr/aIkJqxbPflzdfnUg4EONVotxs/d698Ww9r2
m4tK5+UXkol+nYOKGVkzwuM0cDU/AUCX8bmVEU+3yWcXWu0n1bU6/u0Ql2Klu0DfPpzrjsRP+fMa
JWpIeougEmD08w4T0VTc+hwMZAz8CPgzrk7ktQzvMK/53al7gk8hAd0+vUJ9i/hecjnw+eJeHvXM
T/4PUYazbjuIRqrPQFOTzOs3t4c2bFpbUy9SbmWl5Sbg7pSCaNnU81vRDwrSIaISfCH7AjCrRWjC
9eevd2LH5TYsJzaMo3fPL0sXDZUKJ5emPnf2Ri5jTOvcPG5lxiGTZs+iuh5EBbj/XC3DMjDJKe6j
u5PZGRJPLSO8+M/RxxIx8kMclNcnilNVMEZDMvRVHDFXW0GYUiOyXi4DB9usMyGQQGIOzP/X4r5S
aum4KG3vAZy20bW7KvO/Jmh/3AHBCX7qDUlODQX5keQQrz9joI5a5zJ8lhBNZSyVkugjUkHdUvem
4NTEuXGlGmTeQeF1b0NcntobiaA0EmPzqbWt9P9Cq0IaXxZOWt4NyIfasHFRd3CDKpA79RyVAlIn
g4RkCwTFw08rjNjHDVT8Ozwa0y8WxFZhFsXRtG0NPSVJnBvxB/EwdPpnsTTknAxrP8ycKKUtxoap
82IEwxovR9XrUUXA2tXclWRQbvL4FMRAL2ZwRjUsu/gIlYTwmSmYwXVXvr02X0769o0wtfofqnSw
s+8GpmBp9IvyV7L6slQJ34Owm+Qyo3djSOdMO5lM93rxn4vd0tHxNYxs2REaUHjQ8MSTlnxpomny
dUP2jcp4gCidtf+xM8neRN+IUvrmuKMstfNU8wSKO4KSTtyo+VOo8+gLIQDAda7HCgQC9e+siI75
n/L8ndqE0pm57xfxU4CXamU6SmrndlmLhvohc5qMmipyWq2B/qlwsgPL3alb4Astv7WI9qR77cSX
GD+mhSGrjiF12QA8Y+GY5hEhMebpl2gYGA+wiR38Qvgla32AR+EVRVS8Y56MuOGIOY4SR8iCuK3+
EcZagXbfggxb8hoqn3gNyDbMendjHmMc5rK30M6wQTab4a/4Tnr2xTI770bnsIfvCRHpIcIuPeJV
YR9gkT/kaQzuiec+oM8txBTxiL8P+pG+aaDHWRQAZwyZxKXhy8K76v3TrsInUDhiJDF5qFzSK+7R
sSHE2mayvLgotRt0YiFgkHhEQaWHTsmlcymLrJiRWAfAQEPQ3bd2+SuTRZWtC6njh8BV1KVtvkQW
QBxALgjXH+s4jG97FVAitZrhud6Po5TqV/sKPBSjuXoOI9leKIGrzMUgkkT+fJ3WLU6q3OH/h77I
89MRXTvOS5mZbW93I0EEA1Xke+JNMKCtuCt34jmHDnzEbDFBr2AB+InmjS6SrfycaAWweBem3nO1
VBGlWuNFBcK2/5Qk8vDu2I2o70xc9ZrAIiVDS241xOf58gqmT2RxZPxLocNTrVDT2YhU51imulzj
U/EP8UyMRPtneyl2c2mHznbukHGTXuJ5uT+rl0snSz87OJbNbEdo283iLqrHNwVN3PkcRrPQOktr
qWVEdGrrnC7Zx4cOpEm0z/mOpoNvcn6d07S8NlbtPoC/cwDHx0Us/hQ/nT/jdc2EvDCNdMZb2A6Y
Wdtwrhdl8U1zDUwBCu6OAE0iogmNTstuI//7bvF+kl6Q6TpRsPl48AGEieyHNtO+ZpQvC8h9VN8u
dxCI2ImHvLQ=
`pragma protect end_protected
