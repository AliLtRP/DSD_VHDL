// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EcVTcCRAIA3ouy4IqtIwNEssGy7usITxQCkMOFng0g7Nbj1OhknJbFBDi6YBQ7ym
9pGBisINgfMT0kJWnD0r4EXBoa64iZ7jmT1rzzPs+1Apz7Ld6STpmIgcLV4oPGxK
WZC3S3WG/ehtGXx7fQT9AEEKYt1eEZ3lXx0Q74f+L6w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12176)
jd5goyfDnK7iOctbzpA0nKiXi7Yliq7Kveji2/t7UiKiZp3/miT1GZNZa9g1PGUL
uRz7PS7rAjcdmCOFe/aW9gNOTRoBvqHu2o6DERp446wZLLmTESi6WsDNbFGO5NKJ
V2V+yj4+fsnH9PeQHfIbg37l3Ph7WmUtMkWaYvUuQmcrNJTPn0+5As+8WLh+L5J7
v2V0BF6BxN2ClT0witV/KTLHkY5M0uE5HD+hhBEu5Ps0/RuWUIB3H1kJaxI3Y53Q
uVHYZos1X5XuG/XWAuQq81fC2oQfe1JnC5RvnAeRu2F+TQWt4zvo/47GNfMiccWe
ufegqjIedahMcXQWuNcl7jqtlV2kYFCI7yxCZe3VQAzuG63SImuL2DnTCmaUg051
AbFaKGS7N2H2O2cRTR2KoP15mjaD0B3zamENsU75xeiHTEWJp41piyc7iZyE1e4K
yNvIZ775kJA3jesMe4bTwtUAhdqlLFSwQnSs81ObhS8S03qccG/+Y+EcU+zW2LI4
zQ/5PF/cufXDJ1QgMs44eF9bz6hYwXegJY7JhKuA3cZZWP1q16HjKaxapWw0JPlx
xLK/WPfiFUafYj298L8GkaXFrxwNpNPWzuAartN3XuM2Fnj5lTIgrDpBECX6zT0x
9YfiAMqsxJYzZY6NbcDY8ypcsnEorKFrfVyjQxXqmuQmJQYQRykiRgTVVMJ8LhRv
Un28ONZY8UHIiyEagAntKw5akTFIE2Kq6kK8p3Oa8Co/bJtJ8ixB8gN++1nnfRFE
lBV55LRGeVnWrtIphHFFtQsCiCS0hQlpYMlsa9mtyEUNUWM0rslpV1DE76vo3war
z8BznZjmGiNvyDGNedzc6OrmuE8GxHiTTm43XSm7gi7LWp7FxSrh/YEIPYVUHjd3
Rq/GYTCgL6PeWay9y1x8LSuF2jtAlsKVeerS1DrVlfgLvswVveIFA3CHuSFfiRKE
P966rMovIr1UNSwQJHUTtVn/06GLEqbqZwRr18NDUJbM7heoj53ruqWugVIF6IkK
KGvwJf17s55R6JX7nd/kSi0qqLtZ5S0w17DxYE2X+UMiD3w27pIlZOIluI57+I0W
m7hgszZLg4NgndeW07B5Uk5d0axn37O3r5Ch8Ma+4XAFi94Zmd7xvO3LjuVmFahY
KrxtpCJ31B0I8uraCIf6W+TVazcuj+IwmfWwpEr8CV1UhKsNNEQC4++YoKewzdSu
WBCrr6dHj7aek6QBamwu+JFkyp3e1dhTbMvFE2hpYJi+IvS2CmEEvxEfu7AL8K11
Xy/C6OIykD0sd/3Xj37SRH7MHryEu4gF8xQzYznmLqwUj6fDOc1pmqDNkmqulXPJ
mSSNCThoF/+SdXXQkvFafdeHfy+v2yZkvWl/1VDw5iCFZeR5T8JQSYLPcxbA3iuB
Vg8gpv1ou1ILlOOa+yvwKxgYBy8x9d+UeFoL0i/frgaCF2DCl6iFgLDwcGRxCLm4
dytkPr1kr+ZDZ57nMOHBiTYv4e7MIwPN9M6jSMJR8O/BefJnYhFlmWquovnOeswG
TKzfHoKvT4hKBlXlslcRfBgf5VQFiPiDOBQJtyQbxfsygHbVp2Ckx1z8j9Bwtokk
RCM/WC1qqmuJAhNTdNd+alvRqVylwl1OkhyyLGY6o76AXNtWoFzneGB0eSSf6JJ1
zQO9E0ohqDYD+QoZykNnf0jknKRTbrjXURodA6AQX9OOzAsfUpLHz23qoniKPnUb
FVuRr62rW2b745t5iQHU1r8m3CSPG1coC5eljqOhHfZw/7VG5RvQkUVNGYMLppsG
MHzVO2m3buloVDPYvygEadv2xFN1iidOwRvT33Ig5U22zYpInIEzJgMuf4brGAFw
8tUm7a519InFEtdEeyeYJU6ec/xhZop6N0fNyJ1w25ASY+GDoOKqeJywxB1LwhsM
DEWWUFzekceg0XXobBy12DVJEixgHf0ENPp+lyCXbeBYbF6OcygHYw8PfQgKl8uD
5JAFxN7r9FMmbbjOVNSYY2izhKU4LM9UjxR5sYoMGZdLHpaERarhNnA3N7IBxabh
/ucS4lswrFOy2zrES9fQDf1QkAkDPIX//9BgR1DOaD7VjUiFcMLX1ebLQZTKoURg
g5rJYCiMt0yXilX9zx9PWVv9cZhO0FFgKurMTU2frPfrZFVw+9z+Y3NhpsTbjnGG
EInNfj8xHsZiHWfDNPwBqi9qR1d6gT5FJEI5B675CwzTU4PnRuEPASRy2QaTNvoo
5fq63ynO4UuisbEaak9y1hSRIQvS7lqdqtrqFhsWw+wrqR0uEkHyPzx8RhfVZuL5
4kZBowYyvptNMVBBKeklE0ob9WksPpKvOkVubC6csf/WJ24uZ7hY/qJa9Nzri2IZ
keSaz2ESwyyPEJZToUx1uZ81JTreV5Txoj4/FzS/ZNYTpba0QQkt8OC3Or9Zoq2Z
yf91Mj/+6H/iIvhwDZcPzbWgrnesI3i/ZGc76uvpLWEIVtaw5/OHdJzKnl5q0e7m
qUALM9B8It/woGvkYY01MA7qeQJxKugjwNFp/qcXFB92igeR6vEeKmC467wf4Aqg
a7//YeA53AXDI2Dj4s46IZAfU17s29cgfpRTApjMI2PXRO6zcYRQkRCl4gOMYJy/
RnsxIA6RL9mC9bYmd6yPiT7fSO6VhR0B0eoMyJueqqj4NvSqONq4UYBAbvcmBfeo
mSkg5IP/F7d0YliSlH8f6WnsYWvDo8JOZZ4onwKzk9v6bnNvApXFC0YaTgOg/dyW
dks/yx7DGJnG1aeGRP3OiIJ2gyRXIjrPbthejJQyHyE/XOibLTQetOzH2tVYNUKf
JNozZu++DTzKvME/KK6DB45D+6E0gMXfe3gXZtTW09EOQ8x5BZF2XELpY8LFzuFk
LKqxr3iIzYX9MwWfWVme4VWeoblzg3A9Gun9qCpKMl1RxlmRK+bFXr9JcZLRVnoD
rDunmgqsvu9aBZxVbrbw+rzQxCS6NyvYUh26L+yocfcd8DRLFyGzP85jE2pBef1O
QiX8ZTZhQ/tooqxIrr01WK5A+vT276dRY61CM/uxquVA3Lk1ZnBF5YLQWEmDqyNJ
WM2V/VIp3jIsSZ83ZmKWdH0RUFsgSO7paMXlxHq4tTFZeWx3tHG407hMBdyb3Cv5
mYSBGsbzOj6TvQZZNl0IRPd8bXaqMqXCUIrTFOEew9ZEaNgf7wJtYVcCZ4nU7Brp
nxHwL5jDQL2x/IC8StsgQVP8a5lrADyacS0zGkg+RBKRH1JXmLpCkO4ji5Ful5px
+4FLWQpoWgpUilBLXYWMNyH2xYQcmSWDL1zQKeqrmQUjbXPH0CyAPpbo8SDddkDv
pe4xQDgA4TsAcrF0bIBmrxs4P1IoGcZrOG7UGxxTTUf0p8j9l6EH/z4Gd4iSAFJb
k8PCmqgG+vDqk3JrHy9BBRrWyh00UOzPKgcXIePvlIFpsvpKz8mYbXZMrx2+/6jp
uYTeGyXC+0pERjwomPJAsX00rDDQ4kFUypnspNpGiI+wRcofZ9QNk//IY7t032V6
5y8msDKwXYkz2EgpZEceN5XYlvpE2k5sLpEO2pZj3UajyFwruaRL7qUmnK/3lTGJ
P6Kzd1rDKkhUmTOQkp6KO8tnX2Iasuyr3BPb4dqYMSNV+8ncRY6WSchoy9y828ux
IxpOInKEznYkURnhqNlRGN5G07kmt45AGm+rl0efWZMkXMjU30Uh1TO6Zlnc1lWe
iBz/ceOReDsDLnjv30chhg4kdWAkgYLftXRq/NmK0oBl0av0OGjNdagz88swU2/A
APlGPspMiHsuDP/rEHDYw+2mWib3U8MFroBhKZIgAwECjUGpqJdC5D2TP2Bj0/T/
kWtPqc8j7z1Rgzgpu0YivR2ZcfAJ36FQ5jfgaBK5lyy11ZRRBSaJvhv+My2dkUH+
Yw8C0UjwFUWTJda/ZQJES8f0myEksvQms6pmLlcldxSFVORQAHyr5h3mGNJ7UKXr
pu1xgxLZiIDHRVSzxneUKyDd8BTBknJAy9s7dMOKK10tIIoWtvHG6RLOV11cAKG7
Nxf4TV6GoPGSwL228N2V4z9FTLvX3J0UGLb3qEjeebnRvVEvPJ/fg0yl6sazoYYl
nfj/6jeSHXHechqNgtdqfubk9r1WuC5GiLRYgbnqxbmTOYfbONqqNvQcw3xP8GxK
Nutj6VOJx38Fw7xrTvKGcHH2DXvSwExV7bPiRGI9K+4w5bPBJBgrH717PyZYGgdi
im7MdsFk+rrswv1TWebhH2Abq+oYme/N5+mhfiNC+bysWqW9PTpH7E8ZkYQwnukC
jvZm8WM4xDnTA/oHxTNAVHCPFWrGlanxRwyGzp7Gw9NEplNVi7az10rTd3vROBAX
PEFWfB4wHURmL1BCwdygJAMHlm7sZKJ3XNI7lx3hAwmsXUff+tGcVVvnbvTTHisF
UJZNJhvPY0VKrZ4S+GRcdzEuUVtA8ZmL0CP7wwbVV5P1JHTzftzntRIqxvf1ptqe
famee3eCB1HtyMAPsK1WLjyp5/8x6Y4e+Q5q7cYxSYOpYMQ57akWNH5RbxJujxme
8Tky1HVlZLWCvyMi4jzuOjRrwGUxYW2ADe7dW7ELJocpEPkyOQGf3zmPmnuOuNmc
nMinXBFyPEgXbNAmaEaMHOO1fz4hNIxhnHPa4ipcG9KjWj67xb1fe1dt2rVDT0QE
r82Cpi41esMVsFfzg84uJuRspdkAEbCEsBZDJo8FVKeiZm/zfiCaV4ERF8A8bMMQ
1hVe4qazMt1lO6gNzQp+V6+FeKUbD1IVnxJpNDqxhaoCghwjYCXTG/eyBlgm7mxD
F3P3PTJi7NwfaLJK0DpPrzq1X9iq/SNS3VUotezhlpHBhY6toqdwc+EzLlhbypg1
5uC+XRdP2P/nXG2K0b5SMBtRwV+6/scuL286X5CFFmQ8hcqZXAY7ZvRj2eqgQH8Z
KdpnN3yh6qyuowZsq6GJwysTMDIenjHJ0pNKszM6zWcqV7+qkLoA5ExW44HSjK7F
Gwuk48kK/ogbvEVo/unaS6f/KtwJrb4OTwGG0UjIvSR2+NVVVENwKidBZilT2E0m
feLIh2AWHPllOjKXMlSJDmGGBoYBEGrVIZwaEgwV5ofOlzxFExXy8O+w2Ca3H6OT
r816E39msugsT/AIMHvHCjNREgCdXTAiHAf/FBHIEk7YhaBKfEbE5PYkrIQnUTNe
MfVTHaxBCJYHPsvYDuFxqtqsnMd4P+500LzZ7wUfk4+LXad7RXTSMBsIa4XGuAkj
rwbN1DvoUxBtSL2syT0w2KBWc+DKKKcGyfpHg+yvfJ8RTFfjTJQGmK033a/grEeQ
KXoJdqEWcz7OD8IN4QoEoKOyoiXuG+F9/cFHq80rptwXZT5d0dSNBGDYBQd1iyj3
PgJ9qzjOnQ40VxujEX1ozhqAP+kGRxfZXxxnjD+5ytMtJJVq4fJSYKY0FbJLXfRP
/aho1b4i5wUROJuC7mNpZuCoGH5xc6roNzmSUWHcQtCht/2h1kYcl/8BZ10dSUtI
Tlqrb7p4FWhFW9RhdtsHrPQ01pz7wA4Y0S3IWGomnoV51k5+zRJAScTtVb9C4WlO
Tj/oekS6td1baDNY45GEYB78DDTzkYJk13Ynyv8syVEsliE0at5eaxlfaVvq/eUC
UIYyUvYZeV4hcr3DqVG1H8WcREcIuM2M8IPRTp+DKD66u0mW2Moi6z9vFKbfIaja
QyB7SrfBMRF1TrnAXjxdsq+KvwfNFP1T657ip3c9RbGDfd1v/zrsuWfZngSMd6CX
+elKy1hVIZplVcmRL6anvHBtm/SjtM56eQxMPpGM2cczLAuW8I6jptm3e1eLoV86
gJpRY9Y9+HiDfAWLetSC1c3ZV15j2zYFsRdFiOttr47UQw07mtKoSv5HOjH/QQ/4
ujsM4E0xcbj9hAQGm7GpBRNPVq2B7I+eucH0s2yfImqW3/j67YCb8jBTeEac3itt
kdXeSoybj/ww/PUycfo/Td03eaOACCk/5ZFraF1E08nwAT3B3wZ7YuQuRY136QPo
j2Y+qt+zMf2wxqUNr0nUcK92Ingu8UljbyJdqoSKev04t05gvLTKXh83z5dZeHGb
zl7f/R+O8fpLUD9KdKplBEdC6xTuawc65i72bYsisN/wR4FsjKTjyHpOTsm+/gCj
K0NMqAPsDLkZ3zA/RNSEDc6NsgdY7XzQwhckk1cxgI8ZIpNNlZ/QuKw+3wsSMv5E
E3vinMxsDMtiQg6d0wDBRJVOoz+eRWe0KmzeqDKG5LqFBOmfEc4pv7uIRSaKPlvR
+16nZM8J+M+heq+QU4bD5zaJYMVcfIQzd1U6GZ3A8ShCqjUTtHN1kBx+FKMxYpwq
3HThpoRZP6nN0tgAv9mRxSfokDMLDjJMq0/trfgNZiacHdbZ9LkRRAOFMbStJEDB
KZSJme70Knyzd8Td4dv+rYqiwNX3H6U/jVs5f2+n+2EU/tgZ9lyijmq5DErXPApK
Ll2igcZc0xLyiIH7z+1bxs1E00A8dBPt278Z9k9g14O3EtYNA3zER4UELU+7y51U
PGx/hDtwaMqrgzlMl6eMCeqs5GvSpLZlLwsJ8oK2dwuSFlLsEuyR10wjW9txx+SI
XDDFLbgdNnypBDIYFWPhP8hDSuZhf/Xgu2VBbvocmBdJQaG6lhSrupTrFP2VCPTq
XarCnEEv/TPdAzKL/DHRu0jgqEWcCQN2mJLbgfyBVW3ZIxh5H6BVY1e/Phhj93+z
YQf2FTbz3EdgiWe+lWobsq4IShiaEnod1xtm2gWz5vyb6HqLL1TaxnEtdfKoFgi9
kh/xIRFm3aV6ke/w/iJi45WOaOsFroJFOv3XruT6XTz5LGxindiNW9xHfECkljex
sTvQNmK43jhxflHBe6gXRd3jKfV+XOoIAtr1itwqYwBHPu7J1zpRtJncEVbxS5bJ
fLnC2Ou0LtZblbCBIvL08vBdQURinWV8y43KEmkXDYqxEgjebHLavgssJahBg4eR
WM795dxGjr6mgkNp1+Y1yaiCwhP8waDyd94WghXHxdijMJy9mOFqSlyzHa6FykCJ
psSfcILOcHf6dJSRHlq8L7eZJ4/mec7i56qrKcNrmFa6GYFBO+kRcx1tTuQg0enK
Tk/A/MARilih/o/qs+0AuAjJKhx177QhU0I65SCyLDT0l61tfCYyPZ/io1asrOnB
WykkqqFwnchMmejwm/rsTV2jYo/X3E+ACgrjtWs5HTm/lppyFAC7sNU6EBOFhSIY
R5yrOtxpWQrfl3VefutFrr1RsrrxHc9KZ0447qQ9Tm9O54ZEoIIQBAJUWhmEed2d
NDwwB8msHxXndqOdiJT5b3hQ7DIA9vHqtSgCXq693XvGjF59jHVnkQI5h1/qOV5Y
ewt5ozhafe+MnR1S5g+m6nD+5mW9YqH05rkIRETGun9yjkB9cj1cpN2kdX0xa4J+
5IUMjiylM2o+DuRvru6vVOzcQkIhfe/1sGjzJgOpC3svZG9LN1Rs+xjIawYl1rw5
uXS49Q7L/Qbo3t5jtpcHzRcNewAO0Tnt0tooHo0pmXbIceVH750hbDDD8SNT8mFn
1naRGfYIYTiqE4YYkJVZnkltJiwp13QVc1xp7Tlkw1YcVuSxVri1ySZGkEjzUKUh
gAdMxJ9fxev9apYAIu641O3FCvkUQ83sx7UufWrvOBlFjbiovdnKn46umalXOP6H
+NTl5FqA5Wxa56sXT0bFJvcgXN4ELLivGWSpk+P0Iq2VqcQGI5Ee5U5RS0zp0Mwo
Dx+8NDdBqvg8OhoCTMIMx5v2Dd7G4kW2CQQIhxL11d84aMP7vSdJ0HlX3y/oOx5Q
rxLKPkYO0AAiZQbPSGcgI0ND8J1d2+KaBTC6w04RONJfIVM+/n+MmG8k11k/hdVX
8HrrqHtLlRrpWFelpHJkZLTbo8J+BFJ00xkIRQJu0d8elO838AP8nWpa465s1SQ+
/j0ZhWfGwc/v60+o5C/5RMkPLwwBv5fkS50qyJZIIuFCbVUM6CFsc2pUkbPVshpk
kkevrWADsbQMgINcoplXwRV8EG7trRHe5VdHTeVx86Lzbl0ur50yH5OcG9ynd9eq
EK7n0D6zSdwcwZzi5XaMJmNNukdErLZ4l0LAWzZDIx9RZj61JCONf+opMcoma5RF
l65Vq+6a/8DTCVLJ0vV8DYSivAADWvh6umVbqWII7o0VnovpCWUSco/e0Tb1xzoQ
qzZ7sWn6qJZ+dbgdP5JYm9vbFWAobGH/+0K8+SSOigObN/vyxt+diS18AqMX97/L
zoJyqAXUSENupDlJ9gk80/TZVWbc6YehjTpFVkIA9ahCS7rKIYn8m2pU3yxjIOVw
ao3wxXByJlcb3VOwElnwnllEGKIolwKbCr89cgymwMrmW+NOJleCok1hONOdrq6O
Zp8YhnzXSXGzrmlh+ToIqCdhSZwerHcHdrHolC96mLMlaV2DIRkXB82zNNFYzgcx
h1vKTenxhnNe41ca9IZK79CDvPJOXkQRR1v8RSbV6DRwMs/a2dWqXxYpRmlmf6aY
21zevwR7PRkP76BJHcWYG/u2evPlnrJ6z2Jd7qMHjmM/6lPGXx2B9jrokn/SN5YD
QCYqkRW3l8tIfgmWbDE39KaRdvd2z2wWwMdGMYfPaENefG6L9Z+n1hn5MDWr6Qbq
icbGFw81cc1m6t0TkQ5sEHqGqvT3wUWnfXs9321LmuFD4VNEtQT1FxMi0x9a/NHH
i4jB/p70tLBTULnDf85oEvktNOydZMnNvgOewe9/9m7t0yFUX9hZL+lXPwQ+st5e
1DNPBCLZczw+C2wOiWjmKJk4rc9BFwP4Tm8rVwayUR4rM5079/3wx0fIFQ7WleA2
ZBtbeUeoZy4qIz0XDiCkBg9LAjakkd+uZlX5RSyTAJXuoaKHpA9GDgm1GP2pVNfW
XEIDguI+0lUuHV0DptO7MxMaZiIawtqboHYxvUu4Ffc+rR9suZPiTxXPc/Ks/l5Y
pP8livlAjgZaf47H+Y8kJ+3TKxP4vA4qsb0lH0c9p/Khk4ZBLT9DhWJji/MWpPuJ
b4wJ7o3UTeF8QcVlbxLHMvcf5Zst2Xp2MjcLYLfNWSZrU17ZrCsinW3XE5KoCqwp
tRqdDgBgyjKEzMgxUL0nQMwaOvAleX6PnmPlXSnd2iIiZUFFQrsmbCnmXyQj3aAu
ClP/vhJ4TdRQXHAYrxT+cU5ckOVvv/+Y5Owjqy3YMB3sO/kTfr6Rx7TzxfDASe8z
mYTrGaz0Xe6NxkV3lap7MeLh4w3n/nwM2f0mniqSq2/Vst+dTD+hEh4D5Ke0T+QC
ka9bRfkqhWulbZK0WpIen2SnwqattehFlOdDEVDkT2SFQTBSkQ72FdalNqgTM8+F
rsE0YJP29qs2UCyjcvytB0faxftIg7cwZgjoowKAN+MdepmqSsmOZniKJvf4QiGO
XqqeDrst/lqWSOb1/AvN5J4l/XmOtu4qUN0dvlhMDBaIo5SJv8AhGi3o/jSEo2d+
Yn2lamtF1kE2oLYutlH1yoPK6Ic1ifDviYAxNEQ2dbuBnMaQph0gEZEi1HYyXcg3
/6cSPgR7d1mEhHw5KREI1neDrnP5Sp1juv/VX8q72L/Wruaq8ow6NQ3eRj7PUeDP
QMamO+/YXRGHJbG2GrrCa14YxJTzOB7Wk+Ctq264VrEBBveixOx0eQbtPzwL8vdX
vW9sGihxMA52Azb1s3GgTCY9/nyvQyfaVscnl8ViRTMayOrF4phCcOLu0oBGbXFh
uzK+H6RZslG40E7kkgLMZfBXBVQHPI/RjlwzZDv8wQbgLkkI1Bd0YYu4LzyVAQ76
7ngZXvH8/lAIiwVAR+IJRgyanHMFJ3UXQgkLOCpYSxWd3xLDYuPi+xevC5kIT9pf
SijSaxbGO6YTqwlLFoc96CrBSYuqWAPzEKGigOfYObKxFFHc1UiNkeBJWsHYTs+Q
9kaDa4/vIBljelCb1gr6NOoTTFGIh0aRF8ZyvrcmEoJTRCxGefR+af1ynVcN9jPl
2GOD93TBlMgUUxcGE961lmCj87bIks6x7EoNjzKSQzbfqmjkArMjIGWlMDJX+PGG
sY/12XKl1mVbDdK5PWdPxVmoMdDXF6H9d/LjiUqjTehv66mCamyb5JRjinq3vqwG
lDwJC1F87Ugng3tj7vGj3iqOoIAe2isM5PPqgoqJCSLJ86A/V7cWCxxlO6oF3TBp
jfLe0IJ+kYzjOq5dQzALO+Za2S55IU3WXjS9voPwEnmm1A0jT6Loa+QU4dWo5soV
95wKDnIypXV/usIJiX/jjI/+UBKoz7mahpIC5fd7JKTxFQG/jdilnTvwqO0i1ccc
0JK2CV6W8Yg6LsoxyMCH3xlf6cJJ1zdYra+6J6RZGXMHqi8GWDLB6XflcvJ9k8fo
KRP2RU9vIHbhhADtA1lqlxXDLiLj22dLZ1EMSVBw+mukO+0C61PtmFgOvlH9+YXZ
kUHiiDXMnoYh+warpTUgQ0Nkt9Vb0/rGXHCJ3Q/BUwhR+JqnOX6KnZUEZPABIBa4
Z3LCA0t8p0wfjgxLADGeovQYk42Sv03emeGzgQBZKXqpGHFjGYv4JCaugRNQJfic
CVG1OjgKpj+y80ZDN2xwvHeHY1LcScXvjzGJO2/37TbUtCeEgRqoROjg7cfk6sfg
55bUKKIelXyYI9LxQTtKT7r0DU5Y9R4MRYx1W0vY66C8+YlnPLsueatltq/iR5Yf
/VkZ0/j6IKd/cnUUjkMOVh13vvZAj6GfgPDOeueUVDVyaoLpy0raiBJVM9OQc9Bz
cBSmjJOhk9QOGPNkuOIBLiDiRKbyl/RKx/aCpK2j0U6wNeH9m2Y7VWJfTtw0YSe5
OonVgNOQRAdn1E+yTSIJL98v4hVKbhms9flpx+VXzWNTgjrVyOSP2AUXi9vGUcDd
yiJN6cJ5Qw0fuNDvP/LyR3XsUGJaXWpP09MUD1BBFUJPSkUB10OM9SNi2qJ17QtW
aZ0GV4Supsnh3jAKVrIIkJaXPZSmn7qU3DBw4kZONdfNq7D/a3LsZyic3vTj6cYW
zEKnceEEolcHaDvPiZbqxFP/wuHOECHwes5OBZiFetKKwRAiFnVMCNu8rTwHtAN2
bKAtoP4VNiKkbCo6j9xHK7D+Z+71CVD3lTjODq/j+iBTEVfcqYGUkEdRCAHHrSIG
rHP0OiayDdiHqL3VsUYp/kQ10HxTa3UBaL0XZS0BF9DcQdLaYF7aikKVj/mzJRZH
mRrMbJG8yo56LjauuDsYcmJre87aJCStu9zPv4PNzlBNCCZRujS5bD169U7KKJMK
+/obuVUcmg6BH32D0RGwn9/8+ZIxKz9ZabDUz+qgq3diihi4jnvSnGrgyNyxiAKD
fnbh4xhSHqIfYqH0J5l4QRP0DyqlrYzr6j8+RBO0pU55YkZhylCB1ZGYMCLY3XMK
JNXzrQteP8Aqf6J14q9rJnpM+9gOKDRz187mQC4RWgJNtEexGddH0vDjsEKbygxt
88mgpxk0iCgYkme7VFa3P7+ajbd8b5Z1CAAEFL57sA5+Zmd/veJA2sWvCn4LyStS
6MJ7BIZ0C4wDiZv4Ymb/TxTec3lAJLRnb/ZGX3RUpyNj6b6Kv8aa+jNWQRI9Vjo+
KAdSNhKLeV4vbku9XCCvTqsEjLkmhY26kjKjNATPAhl92JTJrm+iPssi/jzqfTwq
mlnmfwkvkJvn0MLkB59YlP8e1pVjUZRMcbH/C8WUJSwqvMUD0dUUyNo7SbrtN10r
QLdOEYJPb/sPEmrmwD27rtrxvFizgQGYypO3YkCYw/JXDbsb+y0+4cvPvKqG0dp7
SzIiLtOAY8OQmcUY5jJEQF/bQ/HCo1bdAMFsJxFfTAobOzSbADfio3rMY6X1ieui
0fdNF98m6OvlP7G1OMrjLAVY/E5mVDkHSA52CdhJih+pJI4HmD+MusoEaBFeqiQl
2pe0Ubv/Gmvd8dWBQDQ4l6LhH8EYxUQFDY7G9Hlvi55wCghfNyF1PSMaVxXqiuwM
FFVj9ZZLZnUY95ZOMZVU+AKdkRlNBwZHr7VuLs+eSHlaoWzOYtKQ1AvfOlWgAGqO
Fd/jV8t73xcRu3tpEhVQQA/kZuCbgVG99Mv9kJ+lJctHR04EkNQjb0S1ejuHDCuY
obMG5bDaxh247EMcLsGuDpPH1+ZT4lirymlFdiQTK0inha2YM7CogpGxes3lMo3a
rXOwI1YZ8tdpe8C2pCAwykINl+pZD2fymBX/sOLdwcuUnssZy6Pr98qIdZ9pr9Nt
BYWPwWGrkm6/bvQcGM4Nlu4ncWoTE44HTeiuyVSPWpqy6UqFlqhQ2V0XJ1ghBVHm
AqDjS1nxArHHoL/INY/J7p/Y674UJuI9tjobzni/OXfaWbLn3JzBADoyONVKMvmD
tRGGXBVTFT8raFtEu0VCcvpuywTunLA7IOm6F0ExNX2kPhRxh28+eN9phPS3y9Zl
DcQzon28kYbt29Uq/JWB6R/dhwIspymaWvEbzm8nCVEC0/rkBFtr9ur8szmkIfnW
GvmVpP5xwDlsoDfAYKGfvOzFMB2Qd2TrtehOJZ4u2QTCUSvxOkOjK/Eeqb/DEpWT
jpxRomDs6PVxuwsC6/w5KdXUs8Ud3noEocsHYo5RosHnLxAB6+2quvpuALIv6+ET
96xsNcfRx9Zp1T/T/Zh93E7z++7akKDBBdbHD1ybY8HruT8cthzyDhRuhXOiiMxq
dE2qiocfAcYVKp36GXkrXFHJqG+JANKUgVeyfh3wINKpdyA9liPVWJ78p0ybnECl
396FPJRpIGAZ2/pZDUcxxqUGwXNIKglvQLQUHrIuRNUYv+I4nu1gzRJ8TPfL7/X1
TKWcKL0ERDnXeklQq7KIOTbQPa0DZu1U9/3BfGYGrM5qs1py326VurLEKEwJEnWu
TD9SDb4/R1grYHRYmoYJkM2Dlsc6Ki8g4o/pHf91PjHZdDA0LfMD3M9CTNnvZYbe
JWHGJBTvZ9nxXpGh8jTz/C9woGFXwh8685611l1Tuv2ZspQmxpaCgQb/I/Cx3IcI
7t755+yIGvduEGLR6gbKlVYWxFIR6961SftIv1Hzsu/Q1WvlRwVv6vhTgNij+Vzm
5HclKcRamj7BIp6is8r8k9CukX02uwg0gKnu4BnC74NzCYqu1DECSBi9fezqOpR1
ftBQp0xRb1tpMCq/KZ8yh1GSqfsyKufR3HkXRl7upyea+aIcuSwO8XylB+Vh5G4p
OxIlvQnL0oN4IJwaX9cLjIH4n/7m0dMG5tkQJrnTuIN8fIgMKshIxKPmjx22JkhJ
lkYTUqoRXdsvEd5YJAOSiKtEjWXWM3V12TAs/C+JCbe4y/zJ7k/iLzMtcklJiwwT
3DCySXHw5H28wEScoaFe7Ny/yBjpfXm0vs+dFk0cRqpPPQp92fg96EpaS9HO9qz6
ZLD947r6ScbnhegTEKbDx3AcTSzy1nY87Jv1/WTQGBzodQxtEYMs1y09CiVf8aut
2MvOCT29N0Q/YgU168kY2Mx1CDH8ZwRHN634zqWXPjXEIDWkYgvV3dc56oNCdsYy
64/ogOwx2NkGt8gDYPfr6QLZS5wO1GMowfNHKV5waBw6ZE3Pj5q9S7QcGqAODgPq
MgNKM3cS2X7ZKi7qBNhrVJ3eea+jqEXxq5Qtqgqbl4W8g6KZqvE05VmCd7KNxmss
pema8pRvKGxUK9Kn0eeXqDnJryYDinHlIt1eJ3IOP96OT2gltPhMlqzb1/F6djj2
vyk6HXjTnDPXWUTXk3PzCwRatWFhA0UXmrq4vy59eaejHj9VI/rtmm8caAA2I1Vx
vAdPz0HogdPefHtOaUTU86VEwpfP8ZKpn/3RD/RDVXTJDG5igaXGruoNn2DgOWJc
aPa5Pb0s/lKXD/hxr3p4bI7uTkF1h787avFDHfvua8YE6c5XPek7ElPVa5o55aqS
yucTz+xLqGwDHVPOUBPFB/Sqem/hyCRnuI9TMgo5KNDmIz/4iova1h/tbqSOODfx
UBbpEAwnHP34QodSm5iC1wEcJ1NZCzQINGbsNGW3yBsRJZN0GgQEBNIo4K6RSwAb
ijaF3S59mnx326/lblS+huDyYY8EmK0gF98OPSoTqpvptMwteuokAZ5fJTnHH3vr
pBxzEM9kHophwdG+GY2XMgK0XlUusEcojI30eHv+Je4VnzDn+fu8ZMrBVb0xefq7
l0HR5m9/aGiHV85yribPR5eb8C39Yjb0BWUXZu8miU0LDqxLqrcfBFumwJoFtuUx
du0U3Td8nVaMgivmJSwhrXTffcAg94XkdazwkXAQ2FMZg5xWuP/hK7DC8gJ0RHXf
NTQ5nIOB7TyuvPy4roReJOd4KUzebsi8mU+ma9Y8DNHYrrn4CwT/b0g4vtZLboA8
+k+H2PCWBhHAYhRHMcLyJiIa8AXt92N3IoXkHTuZ2mApOGqudlsUsJqciUYwPnPq
btxkXutINUL3r+g7u5l4p7VKtM9V13uM1uQfAnthT6Hnue/fKNxnLL+ZB6MfKPSI
/gm8qW5EOYNyruCXgu89rWI0HuZYNK9BPzYPOxYUHeyfNTYj6APUZgu17M/jIe+q
VobAKsswNSZ/uqN/+hI8JGPnZU2OaR89KDvLRX849Styv4Yo8mrZ1v7MnKQyVDIH
LFtPARbjaFtFV1asIX0GErYHCYxbcYq0vkNiAY1n9ahbYkOrLU6h+tYzu7mQEAlv
XNt7RocvN9K7hMrQTF4XaxjsrZAmyG/9SncPXcXyxr/4eCbHhqL8DC6GOVpOWnHX
ydJki8qoOq2O6i5XXtIFGorHSxOKfZKy8D69zdmUxTkjGoKpwJl+nxuxJMEm+O00
uLeTxPvsUyaN48PPulifF7yMQ2LGbY1cwi9lOunc6O+iPZArhtC3FqpLh0Njsmbu
0wbrFFvTiv4EgcP5vDPYOU4LRQ6AkMsLyJqO90027fPM3BR9qIime5Gzi7lw4Ofe
63uvCoTiNQfJRSmvbDG1rQePoUCYXTLHta4P7Uj8CXa5JGiIP4Tq2Jt05NvxLNwx
sfrquGsMs8RmWQ5XMRGOTiYaQeG86HHBcxgMbae33cgaH56w/0717J2PXpa/3zTc
eQ3H+4jtvdmeI1v++Eozi5AqTy8lWmtPCTMy0YgfPVT1EuwYVkjvG++tdVsiuxkR
fCgUJCsfcUq5j5AApHt26ZkcsiS9SYV3HaPpYezr/MhO8HcMluku9HheUhpAYTgf
0F9UTO0iYre/gvoV/eWrU+lTkQnXcpKlZdKHoW9rgbBy6LrSPDarmBdDcp2JyvHQ
vm07ojwM08pnVNjV9W85D0wzC4gNl87Hos8ph/ZYnoHOTsKaAVfYF/TDSO+0p9WQ
9/1jVZ347AiNtNFHcAXd9Wu4e3Hv7aB65kMrXf21BmJKspSLmF9+PaSR7TYwmmHH
FWU89xSPpYrN6AlC9gVqYztnDYoS/S5r+8jQRZl5y7xfdN0QS6XX+bqxnO+7ONak
Lyb/1C/PSzV7xXzYD4d7on5yLMaP5Jp46VlL0ZIpTuP9McHXK88cDJzW2WfkUKQD
IjmEFS+JNYQieXg1yd94bFRzuAF19jb7l7Gv6xlo9C24cTjKa6/hWZJx0MHPeFfM
kC3wUReXjV3+bClaOIfE0ELjSPBWu6cgfokblaIUa2xgFWr4AVEjubwtSBj2cY5E
dtSpzDzNP/ucaC5itdeOsxUbpqHa7hKONlq0rJDCvDx28+p/OJk24AMDFYaCyXgz
wc7yEVInkD3d8G1gOYlM/O4I2mdv07hsnfxkZ7mD/UOESfsukinbNSpYHrQ4k+79
9Md7+EoLFldDtzq2y+zxQOf+V+zHPZGK+x8o3Y1Kr/GMlD3c53aXHTKsTAysjYhM
AcHvgjOzss+pXVaA1HQRHRUuO6AL486i0a+Wzyf6Uk6Nr97d3jvMdxqxIyVONNAB
WRMUuZcLc95wdu87BiUXf5piWMjlj4iRct4xsfcO0xkXs13Vbcso/wWpEJ11AlZn
NfHiwtDckXcmLbkk8fujTp/bomW8htmllMFeU91pZHWXQjflosf1S9l3fWq8JjoK
EheKpFDWPkxVl8TOzNWCvG3XTp0fszkarfyL0f/QI2hsiUAStv+Jmax7ZoAKH4s1
I9Bh3xyUJqdn5qFfyBI09NXQlYc72BmKUDurxC6qsh4VEozeqPDeZYnTdaltzKqh
qKlFcnUOJtQDJDi2o4efs3xkAoQxih66PNFIlokYQGLSJt7FoclPgwKzSbTnVBGZ
3GX80TI6flLpWRsrW4LMrGW8NBjarQ37vQfbJ6WczoY=
`pragma protect end_protected
