// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
JblATaLsEzPgiy2bxrIbbe2CybvH7VwzkYHc56MF9Gh/IkxQb2UN6aM6tbGCF8TNNcg7FA9wWr1W
9sAFTlhX332sUtVMTHzimMw+5F/vyWaEe4CM5ficjyuiW+zVJNGnTBwDOPEHWlqT49bAuH2YtvxJ
0i6KQ8UmQN1PT8FTCzwUL2mB6tzKxA6tfuSrg1FhZn1hBcEAjArqfKV7no7m6x6LehCrVzico5zz
Ijzo3YKzwb1as5L3dz1vDsFTJQzcmsr3o3kjv2qYCfUBsW84nGIT4qPXxeLNzz7cfCjvsKy6OKNo
c1eslTlCxlmhLJcUkSft67yvqWU2A8/lJtwExg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
HzDWc10tNWEFef5F2p7EOna8hrdyiybqGggw5vPRen9xURc+jG+fcKkFYaMDSG4sRHyfFwcV1WCy
mR/QyOTEwlKcU6ZAVZM4Y1EQSXpA7cF6uo6K7kEc1iXSGUZ+QB+hWbF4tTx1Ez8/48eOzTvuRswp
5Wccn0iNo9gwwuYD6na2mKKYNPGpEIhtedjMHb/T9G1jSVaSSD8Si4uoG9go6FK3hzOMy4ldl6tu
X/1fYbSoEmaYgLfm18My0KCv83M6Nsux7v5mfAtavvzcR9KGk6o8XFWRqQpMjsQYzp/L26XTbPhQ
+EL3vSro8DTd1NkxENEsraK9btr7FYzKlsE8mCs2zHQDKOJvYY6Pdiu7VxBp1gvU7rEs6sH/BpUb
Qj0JDfG4m/gvj8Fou4EFyahiCu9V97k/sEoWXkAdu+IQDQjxU7X54imSZVFsjJ8J8qIMgTQMZx6q
Wk3mlZeOYK2zl7ZZwfeU1GX240OyQk2QnjP+ClxOEkjHBI/eIb/uOQBzDR0G2SQ2Nyey+Vh9kf6g
EFUj5QuVlR086EBfRHOOD/H8ekBxLInW+xRyxpnAzRrdeVy4uF6Zw1ojZdhwMfEJQoZrTnhFxPup
2lp6z4NiacQxyO7nMEvmhXmEKuTpAAKvmBV/OEUrJvFsxmigsD3CQoUvWvm5KIMYnPj+5N1y6Mwm
6ay3Kz7CVo8GLHfgRofJMg8ESZTLBeaptOlR8Dm6/WYssNHlv2X6B6N6anLqlHbcLiQogblBUC4l
VnAmxl4tRsfMeUBQPMAaGEiztYf6B7006c2eA28fKAS5B6RXgqnMmwsDi3eC8/zUd84BChrvjyyE
g3u4p2WOyVcUrJ88DgA8SOovf8A0NJfl8+nDdrNjD2/WRHWaNeR/vF6T3hxXfAXb7S9KpCaSi4sk
vi5o11ok0p1LrvlfbZFfGn5zEB5DWDQxya0GzdV1YytuGECcebTalx6zDiD0foXoN0RrmPP5s+sD
PPlLc3/bhhF1lA20vG1Rmg8/Naab7lG+JTO9LfRdfRMFp1eButKfKfPz0JjzUNwgYaIzQcHftn8n
QkDsxFyDyOlxbcpoVtPjK63LK0M46j2c1XPpGmxGNfi/kxvCUfbP7P8nY78hEuGJxuNJs9zNJ4mS
1T4zdMjhRxRI8GpjqTlqJI/TUCOpI8krhwAZ2uxbYiZaCEhkp6ro42iH5o69smaR/eS6X8SWXICf
nSf/GJQXCwK2/AXYLmpSn5dsHME0GAB0AQRZOBMPHuMJPHNVfVcc7nPacoqNT49nr/VvWIsOQF47
1sEPMud64ub6UPi0KSVrZ3xTO3mSU3cj9fyRAfsUj1t1RQC/6YgHlaYn9IQr01Qpa65TeIBsD0cl
wjlVjJaUPxwtSjHfsgyfhHymBrWc3y3ADX9IgE7dGmum3HaNWEPjcqBPaBmZuYy3THpNqQ1FHpOm
sX0w/nkT5/DgGW0D2DqBh4xFVckhg5SSxupOoxKJ05b+zg8EO++qyYbqDYx4NZQejgioih0GvJTw
NsQehCzJhBBOKBgSfyqtP+Ea9uu2bBG02+hRWjj8347BpOMjlt8S3HdqlLzWiR06qjpAX3JQcQm7
38gbYSMXtcDFsJ7iUQBTo5WTHXnALgLmAcD76J3M+5IZIKHEojY0KVEcSBHwi09cUROrpq4lx46Y
Z2q0VBcCSejkhusBPUTN8mOyWjIMqzflBrZ4ZNSj2OkcuoyCNkqatxku0S4TAUPd3wE4whcNTvRo
5CvDlzsc3Ucc7/EUUKY1q7rReiOQCJmNvPyITyYWTc6Bau0rXpjZJVam+lkRpsu4E8jJqtmCu6zF
cAm/4zF44WPqpDiF8pEAA4gm66Ol1C+S2RzLQ1mABoBwWjgURAyIe9fUdXKzJFtm5xls3xL9tqs2
KFUdgmSuOTrwSqqGP7Y9GFGb6FdPTym3uAjuOBL+jT8Lgvw90MrE2akKNb4bWwPyDp3ih7Iy4H8n
2yCaW+KNbxJiMsnMeshXmWv9J2+MNvVtPeAFpBnONw/oUitxjsa9qA2Gh006l2T5JX3DPCzN9P5/
zzeDah+a4we5Ao1Eu6gbmpU89hPAthwRWOZNMCQ5WkTRkErSwg28L+X6e+b/8rGmMyX1bgjVlk3f
vCEJGN3q6xUU0yPVWS92xcfuaU5G395ySjj1fw2lHBB9hBJ0T0KnnhHvUGcmRVSRLQsyySeSMcKF
sI9lUiRL6ZrohufT1Bd3QYU+Vk5oV+9D3MhMwdSSLil8+IkO0/5EZ1Iw+gkphWAXEu2MmMAkn5jx
vGCS3KZJoQBudmB4LIrrs5QIbRmz1b6F7inVDXxUwWJC/WmUQdCO5Sh7AJ5yCWQVq1NG5huJc9Wl
Kk3sp4Lgj17ZOuKavL0C30uhdFnJkkiJBYTm7P6MZTH1fsTsq9cMJ2atKP61DwR/3Ty68h48hs8V
0QqL8EhGljoPatZrNs4hEhnx1ARWQPj8L6TOfG6yk1+v2qPNB9jcioyhx+QOheMoNU5eKr/m8dO7
GbqJ8qI/iS078nl0WiOtRXOVSNsAJtVP6Y3Dz9oIS5LLPHxz/csHhtXaleo5g5rMID5Pr/JDzsAk
YB9q4sUHx44fM43I2R9pYIs+RL/Qt76jANWk8K49wUKgfTxk+sVOK/gdx2WDt+WnF3yvBj+xcrQw
795EVzIhW4v4Vz4WY9lRae3F2tYWt39UrFQjcVd0fOi0TtosdR29UE69MNwOephe/n80glI5YHqO
Fl4jbqnQOdGzfV1QDoHihSB4qFwuAjr6lzkiSbzQDHQ6QW46Uiloo5ilcQlQk9zd/fFPtb1MmZ5X
vNKjSM574dfPPWRp+IukJ4h0hww/a9Fb6CthWXi6OyNXdBQZPYsgV1bEc47iz+TwjP6hr9CuMDih
UX+umGjXJCd1++djG9udvdReVcoghJT1lqNQR+g1dPvrhysGYZwqdvhhL6CDp3QPZ/dpnoiu+oUb
lmocNMOOftfVSj3STmRUGiOeHyNK6sZalbAAEdH42GM6HPbyiGJG1HrnU5irXIZsq4kq5nCzdqlp
W67Wpb5Qkcwj7MIyvRrjECgK0C4MN7bnJ3QDSk1kB3FX3AtHuv9w20+IwX6Sy4IDVSU7wAjdNgfb
MfDI+St2G7YDpDku7XWqSFNG0YK8xu5nQxhjeISON2G0el6XDgPPAUyp04DYi2P/em6QK94HA12t
o0ezYQNaUkIn+jlsjZr8wO6rX92/Zq1+VcFlklTdVdEGsgOX2a5s/X5KM8jqvUCYrwVigHwg+xLX
RWtsZDlSpFOo7uFMjsbTE/W3K0uWv/AbEwYWSa0oKD2glwueBTchqTruQWJjR086N54lKw+wQk4F
IjaPZ3x3XIC3uMk1uzidVM3J/LDGGuWqtIsRw1qViLb7xXP+mzC6LugZk276yAEiFo03KMzCpHkE
27F2JMq8CZZ8zAtE+fxN4zVE1Mf963OQZeDBrFK1TY6bC19NBaJtQ2EnKZ4DbvxtGhwx/RDHlRYA
nR5eDH2u+9RpgxLvXHDT42wz3EJlKRqY3LcJ52lbBSaQMLwxoqG6pkZy5sMWaSNnpdniTcqVdY57
gP1IqxLJuLelJDgnd2fttigjck93dFOAhLBN9RQRZGkIYImCO82ZK7GW/8MhTqt/0/XSYIjr53Uh
Rc34UbPrKuzg3M0Y0XFbqiCaDK+Sp69KQdMWJc4iNbscOw55FIbTaEbLi09qqOvZ42HwGTpCM/+C
cSI316GSzXKqjYWN9jutGnaRnZV/UqZbV1xtSMNXo2s4Yd3p9ykgFK85v7mOErgX/ZJIEkLhvop/
yxRGSTZuVjAj2ab8GbfUaAUcI0ih9Q4ZPp71Syz4gAFWDVIYRpA5sCNyhCWpQo9ZlO+bf5aj9xQ6
0CMyEW1kHgVh0wC/gUu4At3yvH5uikD+WWWzKqO7Ait2D0x2WAQr5mp0O1Xe7NmAZEqDObRZsLps
M21dDthsifbfb9baUir9IHWGsVsEOmZuVHaeoxeAjXDpGWCXRObt3N0soFBObHP70rDCPtJOS9/y
IB25a4upR1eAYX0ZAT3YiDWRbiUvwnFoPdij+h5bqE4gKCBDMntRFPDCPbqcQt9uHapayTztDWiI
x41W5hUQzv6Y7fPdewODmwxisUTLDb29/7odrVvesff7ku+gTF38Mr5oMwT2zU8ZqvApfE13ocll
z6LJYQtdhJiO9xBes73OTgqUz+AMD0vY6IylFGpN/6YRGTh9P2Q1wov27nP2JFmy7HF4cJUkeqeF
hXLHILjI2fNNdj4WQ/T7/2SBTARFN3gdXgY9NBzfJVPh9tX16MixJnvfzuzjgT+OnPCt+LPGqETt
Cag3pbggLcTihOXpK/t9NdM8UjRq3uouyhX0NNZFCZyIWjCdR5WtwUjKDGdMiDeuCfaOhTQXj7s5
MDGSjeYcEXYe5gtreJ1PNx6VPgQSZFcGNre5Vx5OZk+8s/Rv1n52j2Z/9XKddzBAop0sW3kIii0f
sfJ2lWkmt3FLKcQ8wzgq1cUQbVHwQQsgKf/BsE7mcRMDgIFNVygJY/R+X1hdEz+0jV0fLgOw+vvS
WohYgclZCRGEx+Tk+FM/QpwZ8jOwEC6kZrvzbRGPi/i7bv/kQqqJm4baZTj+b+Q6HuddIH5Grzhi
tJmQIU+ubnQBLLymuIiOY/aluxaLNWqmzPuv9r7dKn2F39xfYTVUVJz9+56dlCwaBRncsMBYSe6R
lM9PZADW4kat3xqbXrxtq6cvVM3tommFf/LKLfjx5Sshn7YtuAdvzaFYiJoLP9zoO8qPMLn7JhLn
dyBb946ikQqUNrYf+MVaWmJ303//H7NXpJcTYFIt3ZiD6uJSIBkxZkDGp8RRFvyPGKpeiGHUnVC2
OEf7u8gr8smCFGeeMDR7dlBJ6ca5X8VCY62WOdBhl3mokh2fV2hRaDBE6nQ57MZvbW8BGYrMSJWL
FvZq/HJr0m2J0WieSewu4xucBm71nAc+ckXzgi2a1oXg63wPO8llz6CcF/aLd23QpdgpigGqCMFg
LH0yJ39x3DT+u/05VxchZC8ywMgEuH6FIH0YTF9NOX8K0tsB3321uzIay0X8wHzkE2wkJ5v8V+Xh
D9bXrcsf77ZlyZOe6lbdjSVhXImhV0j7NwdwH1diw581ZczrnjBBjw203a5ZmfrfgE4XhoBzAz2A
QzASuDTzH659YwaO/z+GIOwt4uOXnDssrtRlkOWVURpBLSG7EQNQ0hMf4LEtiIme2rU9cSHCQx2Z
hDkUjAGUYGkRCVsWueWA884oGsfW/z/6So/arGpLr0ahUUQ7SKk1pcspDhDuJqfjkiSa9sur5I2d
jhZHQOMjwj37SEP1MB4S/tz7CTBoRT7ixHlv7UwJhdno1ptlY2yoo8v5zJNuAqI0xT3V9osqd1cI
3TaUqkgD2gEOHv32G8CtqgouhHZboM1cJTJWrgMJo6gjNSm+5LgQyI1/lKHweXX7nrH0hVJxVXbK
jncvxKntWaje1v7cED85q2VDS+XIUYZZA5bVsD0ZCEK3lgdv2nVTRy5j2zNL0xknf4TjbE1MHn7F
0FJGjRRJXxb2HOkiNDxuOPwpiDqfpEQlIWGphVPwDw683YB1237JZeIB2RC4jKH0N+Krt3GoOr0t
5bAnC6BykqxMUAnXaCnYFT0SFaRyNx1DNRQHPWyaq/y6OwTC7AJJBYjvNI9+5nedDMUtAT6Mjdjn
H1OI7w4bG3UAFFRJ5ee3poN8iqE8Ay3w9/Q2xGaIIEU55EHlmzuUWoZNwsveVQnl+plwV3Yz2+Al
GEvqD8o6OdTsR29Gm2VasAKQh+MV5Cf/InYs9749rNIuG3qFGmz/wu3yUkKan8a7N9xfZSV7swJM
VyDSpMeuZLK/TwhvVaMVKMacMiaJkIrHZvdbgWRPuhaTCYyLSr/ShwIO5y3zKsHo0hRhoNIQUSX9
4p+0UaFPKAsEJlM0scjJuoEJUc2EVX1MM+eCTOvzkGq3r9gkG+X8f+/YjIQF/2kor2/8+WmE41dd
clIr4ZRrB+FEBb3e0Af9UAvrZvHbP/XTjLydwHNlBNilxnIoZITJ6FB+582kCFQRAt+AIZmB5ptr
NaQnsr6Ml/2ab2bxJb5thGCb9U3LK4IKVeQKM05QrV3kFWWJ7IvRXRM3mg/chmg1vfF91e/D0jz4
CODcl5qtalzgrpSVlpd/ZqsteJT+U5Go4fE1hqnZwDNzIqM/kfgcd4iapmYegAAfS1RQGS1BlVjg
CaDg4f5GcHZr/sUSUFPmFrnwyIsZQBz0fOZ2gUobDm6jFZPczfxH1CWrmDAypl7CWSvrxvxodvlA
2bQpow+rBnyblKQuNFiFGMAtQF/UHU4zMtGRk1zqeK1UiwH52ZNmB3yg454TlNJ4rXVgObxYLOFL
pZlF9Osash1f4hZP8lZxab4HeIEAlEKvRlY4IovXuApABeqi4aKFtIahrJoMQ4TzYbcD0VIPF6ZL
7rQnyzOhGsnPpaGBgE+bNACJvBtwFsaC33AWVxmTkrLXJwd3ukHosAuIuyeTUbDtsdshl4kZLED0
JvdhQgy6IhzGOIMgzTe/w7u3BwQFlPPndZ108Uk8VP7FeSLQcjLroDxAf6RTDgcvDHCE9mw6ZEaN
a38xtcxr+QxNaGx8zeSbvzGRQbuafFEhqz2G/6XAGtT+uwoKciwqAsvM9uEwh5MI2kNmZBDQLC+M
HdRKhZprxdI2bpe18PfU60FOMxwOZf0Z7QdY6fYlqfU1p1aztTWz0qR1ZWQvZq31y1xuRFajhAPj
1gMVdgLeQidGESUaKNdTc0/FZAKMYXtaWqt1gsB4Zu1tGLIdjSpbLL5OF7Fhz2BrtaJ+H1cISSCd
qjNbnqF0g4YblqwTigSZJHI6QZNpMZMzaF4ZE5YhlZz33pAO1Cc1LebHhDhSMWVMXcE5Tmg4onPk
LBanMv1A4NzlFeGZh9KMBWuDKjBhOp0OF7PPlA+2xXvMAwBoeWPWgmLnMKBE9ToMksXZ/4CPpdxy
jxBc8P6clXQwpQbnqEN6iL+yHd8cM5xRyVgnfByQ1SBGiXvwmmY1OihmeyH09TtK3v2dmMc/r/M0
lwLEUNAH5jpiPN0jXoDmARUnkIRT5tNjHybAyb67vJ58Cj9W6hMwxIAFE9J9oF3okH56mTqwtlQf
qrHtISujr7chQUFJFoqZKt/7w+KHAu1bKy5SGKIAz/L5TWNau+zn58apEgaqhlVDuMwaAvuryPCv
kvX4xG+MxiJnVhZeFrmwI7S/eXvnuchL/zNHQcb2QLStb7jRlpN7ZU2Vv+XU5rYpcYJyroqB6oUv
vXUruxGcOlwrxvo/ocfgwdloyyxT7uxPWMGaTEy3wz0tgTa3LyhoCBx21Va371dzkq2Ru+Wmd7sZ
ZAwZ7vuQDz8KW4QjyNUxuekHzrg/t7cBfVrr24X7Kqi7Or78Ll9tZAHF8VxOy0v4pZYbLXFtv1i6
fb5xds9NWHsWW5P8FR9Opyt/mw2mBO3nAm0Zf6XHP3fxxJvMTQ+r+j2d4nZYyYIyCMe4z8TA2L+C
7xHFCrAue3KuTImdt/CMqKmvf/i1fvFADbmMJDqLbvT3geUdRrXvpjRYuvhEy6dRjfLxWceO74PN
jxlqVGo2oZ8qlJn0/O1mkJA/spQmAfvSh24iFZW164RMorYoAE9Fma3V8JfbnfjWFKg266OCAROj
lpMiGfiMKgGGtYviTRUS13kpS9nG8J107/nejGIrc/aCYDLVtvjW969xgbyFYjTpefNCZIkAz80H
E/lAcXkCvD1ddGUEUXPlByXjFTjdU5+GGrFLJXOHA99VERAUhDEvdqf4RlMv6+AB2xvB437hSv1V
xBjlHYXKyLI+JhBrOxBWbKOyu9ci65wXuqGgLjPrixScavnX2OY40fI53yf7G37cD6jjORLJ6hSX
DMqNlw0R+N6gnTYIasQVDAIbO+LjTp/liZpG/99dN7AMW9v0XDysSv0T0cPrXj6CNQhEGFBBNXiC
EObXooD8T7HdlROqfrjSBkUx+AwfJyvM5zsMBWIhaPewv+oIU0njSa0ibn2Iqy9jWIKVp/y95DAW
AvZg/cEfaQU9smKdABuR1x7BoeUBWtf+k63MRl5tyEOjzq47qS6mOSGggqlpoz91B1SBLWt/7eGy
IYDllMZBD/5k26qCotjIC0H3rLzNvMP6A47vdzrB3rbyOHzkWlka/FwnAqUBLBbX6HjKAs1E/rGT
QFHqXJHikINpTt+SbhuzqV+vw+7lBZgdQCyi7iEoPC2Cgmrj2tWEulN7KxHdvZD5bNkh3h+oj+ts
DqslN1kA3OdITDaWE+cgjt/KlbLjOVn5X23QA1pRAF5/dcAw4xp2tX4w60WsJfHANT8q1LF/dyu7
CDfi/D7ngHXgE1BgJUmFRstM9CV9uHsuyqEkmX2EWRtVYKItd9mr/2h7WQe1fF0MnVQqIISybNUo
NQrDcwLcRowjXqD0e6OpySbvviYDSj2wzxBfcGFQeU7M7C7lYxByFHOP9igH+sES5u7gK7mueS40
hEivBDP8r1fkr58QQdrJgRjGQ0eSTaffH2Yut1T8drzYH9BKpzd0d4ZpIdMSnoH5nZRuRuHOY/Wh
0z/tbFZBBwmPVSgTNlJVidr4eY7B3QAZfS5WQ+M2/5BwjBstdiXal9M0U+2U7R8WbIIWuZlCp6Oh
ewLfFdm5cZ7ZH+j+42/tvgrIfTe7jG6Gd3vzfpnJa5VVqWRrRY/FKsPIH9jAJkM+huKqWDU+lgY7
/4TaChE8QwtRhD7Q7zsgQ1all0NcB7d7ueMRguV+qujoPSpDwqMLDs1IcTnA30N2JcrvcrfThYhf
rYTOSEFpuupOgm9wAsC3eNOedftNRjqaxrXrbMcvEGZsLSrDa7t/j6kFZdqM8hxHZA4B3MMYl8sn
hOjTAMexuS9t8Av/yQTiOJ4d9LxetPQEzRSjnOItvM3nXv5nCMQc6GhUoK39U3kV3Bt475oJOScI
g5rFMBmy1ib/2PJWmzacjda0Z0PiRsr1dAjl0czqaNQHXS3d/6+ufjnxw1AJvibKmY2tICdsnKTj
mNXEHxLrQxtY2l4PrL4T3H+wdwS9coVaCl2c4gIh6RAOM+2+1ihdO5iqieb9vBYboHdSS1vEcbfE
KP2P/spR1h04eEQuYjVvd393EdDxMTlzqsBbtfvzMlF76c+qy0rbaC0C1jSnwXM02T8c+PVvd6YD
9jRGFlVisi3/UKWK91aapEsVHxDgGZsGrXGOpKk7ZwCLgy0GgyeRj13E/mDmNvV90LYfDn09MVSH
qdMqxsJzrnH8jPkE4o3GMfz4Z3854tbeDuQ6VducaRrl67Pl/xbgLwxRzV4b7bsILuvbjSDdS/bb
JlTVLBXvfshYWltLDMMgT/acDeEFtnrBrRYhE5jd9gOtnywDlKnH5F/bCVz4xLBWMfU1BQaLGsUP
8B9/KofQ95i0YThkpj7daSOY1mZ4iLKiZHUH+h7+DEXdE/SYs/ZdLUGh5r0ga150BQKvqrSTbJ8b
j/9xgHgXisjVTMSdI8+1448aacnV1y1UiwcpGwWIr1XuWtS8RbQ2P1A1ieDonB52zAu8LJloUjQZ
pJFbETrpBcihG6TK4GDWUJ4D1h1s4NGtZUnloWbMWl+Z1o4Qqu8XF1JoafdUzaPSfiu8Koe95Hl5
qRUf+f87KVZMD13rpZkQCSW9jaYAH9T5LmAl8S+0QzPu5KI3t3BgADilDt4fbJSm5DwwaNka3HWy
JjqO1pFQenpg5fsdihRG65vbPFXJZD5RRFTPyuJ6zlH8cP8yMN2B96l+4nqNW175w6tyVZMjyHBA
OsSLjQ8mku4DwHj5ozyu3OM9wLfHq/n8WPwsWGcTMlP4QxLG5G6SPiC3mPKYvj7WKd25O/BpNTAe
CVlzpa91y4hFwlhHt+/kYyl9n+Cde8YXzUFLw62vtLRlSPc7mkwJvZqgrmSuyDjI2E9m5iPRwfAZ
0qQQOwUTM7nj95lr7yMi5z75JPPDVsYw4bdVSKIawca/mC0Q2vVaLhxrxitEW7v4FBC71VjDHXKt
7j1pCOxKiWm4gTp2dDhTjw1q5KVf8cBk1tl+lRhAv4Ux1uSD5wzMjm8PNOhZiUDTxnrC8BMbDDDG
oCC2b/j1F1TpeEODgWwmW34/xMLQcbuxtF8ARkO3czGsE00r0tSvchnxBvm87NQh71Y1yjsbiKd2
UJ8AC/3nGUMxowO62RSZKE51FCbaOUOgs7LqYvnxAVNGZDKSrHdANcaTnRwdJd2ta4Lq5ACgH/3n
9GGNIvB/55FHXbFFvdHiZfSDRRI29tHC/unSJTggCgwYnophXkB8/63arssHNJ0LIVD5N7PRGwwl
14cHjV2Zw9PipQ85UDg7cjYyyu1c0Y/i7QTsle7uDquRrG/C/88+O4iUskTvRPj+WK4NrRMLN3C3
y/t/V4ItM8XxI9UubbFJM1JF1i+6Xequf8r9dAYt2YaNAI8xUtqeOgCdihiP6NssZMUIGhkGcZYd
IgFumcVy6qb0TZl6PCYSsDkDDC86GUANoj1NlWtiYwMRNJv/pkf4E9H2cfnZzWOQrRgiqYUFsAtr
GwSlqy86JFdYDjfmpZECLLqYEC/rsUcHTC/W/OcwFDFL1SOBnnztkxr2iCe3+VEb96E0h9+xxysb
VmdVHicuSd8APx6cNk15e9kPxKkyDlGYrlxFd/qtLjmVJqd31BTMJUVw/uQr46eustbkc/n/CYNX
ns3Qz68ipqFJf0UN9MaeyNH6gySvxsgkRs6uc1UoG5pfq9lnUTQVoPd9IeaU+z2qhv6+BvGfUHu4
4XGamY+7Q1jlkTdm5RkfS6kBMXcxVtWJBP8IHan7POuRLvGyK+rhBTT7aEHAp3U4pi7PDz+xjmeJ
Lvs0HdIrWRi+EPs+3FzAZ1abTQs8f5SkrcwvMjXLNGzGYbRXX5tTWDeNdhSjR7PTvjU3QLy6hiCR
zOIZp2taCwlnTIC7JPNr8LvM51ppi/8olEhIsHJ64DrxeHkVBRDcoRHexhXN/11KrW0v6Ob0QDb/
TByqegiomOuoQea+rQ6+KT8usjwhHvniU8BGaG4G+SvG6Yn0PUUGSdCsEZXLw+f+zzSfm+eDtsCX
FmU8WwVhmNVPCNoCcSG4iNpsUAgz+ZZjgUGOUNNVAergeEOSFwBzE8wlQsWYtBXhhJ/fOVoxbrnX
y1rfYX93NnSlR2WtrUeNdBnufAg7RtEDiRxvf9Kl/UJQs7y2+S99s3K5pw8vFqs0l31NOmaqglhI
WVDTqYpXdy8UMbg/DnltWg4Q5yxzlo2cG//e7U5iWUSyCa4niFuamKhoTZZfch5gK+FBDTYN6a+f
cWmTlQf6tG3bgzMZ1IIX9chlh3k4qbtrGGTBnTeNBbs4ZjucH998a3kb5B1gMvl29OB7pvnWTgCL
tY6dbqWx1OCiB+GeTcQXBSA4MKI8ZK9sIVGLDFMhp8M/QgNp2y5O9fbTciZdgskiKKbelbYFlzd3
ZW+LZu/1kjP+VqzF9kW88VWd+9mTX/GPgwBRf5lDYsB7CJdgbMew7+w5SolLn/taS+ORs5DBwwGk
n74jN+mhsDJuu9+eiy3NEezxgOo5UDEHzUKZdEsT46XWEsHfUkXq3nqA5HcgtZlNBzSnBy7nam5T
7rVwroNk96NgK+6S9+bJ0h94Mz+zHt4sXannMi49M2z69sHwlA9W49teJ7aJLeQ/m2j+WNTCX282
Mv3ZH0m47RPaSsshHdpRhlzSTa3mcHOxUft88jtV0YsOjP9HOkPmPmfZ7q2Hk5k/SjMTRAGlI4+Y
gD2terd0T6q7a/zLbcST7/WgsYudR4qduCm6Ngk7+onZe+LCTiLoLE6KKwyUsXDuLiCzLG8RLjue
hd15hpluHFhErVqdlgP2Vvu0uGK9zl4j8E+F5XXlH7yZGGABKpXWksmRmRWGIjW+m2hvIynEYd0P
nQgNG0aEwz3FICcp4M5ghbDbBZ2aPj+Xfkz601Ui6LFPlx90L4L5CcKl3HFJxLbNzGlh/Z9sJraA
SEbjKRYzgKXDWA3BKo67yP+IB4UEGJiqFzP6qmcoHqzwhhJVcQWnToW6qs/HisuUh0PPI6UzEBfI
duxoJYTX5efTdZ9BjLztOdD7a2/G7mKZ0IgCmmPmeNR2Sp14ltnrRTI/wkdiU9VTnnsGhgL6SbPp
p8laSPXXqsrCAOglGWKHewCjFaPl8ZzpzOhO4v/r2B5O51ey4/zSheSAYhWsoqvGLpcVjR8i1Rb1
/BhFF6sOak3tPHGaIsEqsaL+7UWhKlkuy0i9sW7HitIXrg62dSl9mwfwkwWregDAO5gsnQJDqOhg
HbJhxoukfXORAo/1BuCrJGkvLr3dYdLRNhbH7yFyNwCoA/m6gib5o5TFyISfqTIjyox6w+oOHISX
gzMlpkbPGoR6L/4YqMLvw+8YwqGfr+U2WOA5YJ2PPv3RwN7C8NpApBodl5FmoSE8v7Mo4Wr+s72u
fvdAplUthdh/M0jFoytnHwUQXUin41FtYNywbD0KCOpo40PJXU0Bm7v7/mKGmKxcIt1nPBFIo+he
1ABKm3elkIHKO8aLhcsAKEjw3Lkk7bWMFt7c8O8WCCRBTtzFI8b+ZohyhhrmFb4ScjYnRnBB8kgH
qMlGdyqNrrvE2Q9FCq4qUCp2aeg2HzzjATyB2a3+1BZ6jg+SX5XrwlddxC4vZ52PZsKbza+vlwL8
esb/7RB+sNNOZ33bBHAhBfcqGmQIDYvRaRVMKpKS0/RlHPVmhcYU4Nvljkc1jCZKHWbdpPhUWz3I
vTOudioNdcajB0pjK3AdHhtyI+o1QCSSpPundfnFQBSRfhRH50fL7kgBp4O6FUPqDU8TJn8glRmx
DoYLWmVlkMagWscLwdTDhG5qANTdiP4B5Kvj9bVV4giZVdl//T408Olj9I8MYHKj9QwnSy23EeSk
rYkFpmL6ZN8rWyerZj9To3Wqk07oUhuJEBcECis3NXn3gPl7WW5Vrhajy+vpdhTsyZvD88Omidv3
n9VQq58MVovpS1N3L3cihj756F1Wf/gjRRo9CK3Y5vdUfO8xg1Kgqj2mb5CQoMZXqgl/QdMV6HZo
VUWZvz58EndEVM+1dofDxhCMDpwqnY0Bnw6d7nfNsNj8BXgjwGLLxzWI1xXS6ZzHJgTn/oD3OXc7
HDwxhKqI41xGgZpbrfxqYCV7tLC9w7KyGfB0/iwm92Wd2J/cT+yn81b9LDOB+uq3AZDmhdlZzTen
w4/MhIKWvf+sKXj5VCmWR444X8aszoH7IFDoYqgyndb6a7+iBpDQW1GT7iy9J1xdG6M9oE9Qh2Qu
kxSS6mZTl0EABV6/iMSVQ6TGmMVusLer8AfcULwFfmyx1icKE54CYUmFf5raGHv6g12SjicxkpnC
t4kUg+crI4A1v1lLaztRUBKgoo4G3oR7jcgOEQYg7WJGgP9SWSmjJ/BQX8rTOnAa2E3jVcKdlbV+
wmd0+Y+uyn1i+zvFroyGWOqYs1/kdr8DOXKtxcEMuScCz3XDPCoapxg+vkOCqtY6tPzvtEyHCwIn
UI92dfnN1bUv7tikSgt2Llvg25ZSanrjpStaUET8KVmvnGQA3LsTGfb1OfPRHj+A8XUnIg+4Q+Dh
Hjwq91TgdAksi4w61BoyEZITNnahSkzPdzCPLzru1PJN1vE3prYR8aHBJtlONdLXcn2Glvo4k955
ZyZVhXU7b3EdrvCEf9Kfak+Fa3jO5bJUKeAtfkflkJmqVZjwy4K132oYmBk4oioGE5oDEYMBg94e
IWBWRG3ZRnwGOc/y9vQ/mESXvkI6Ehoaw4OAAg+nbXboB9CRx+9Rk6K9QfN+c8K9BX/f7ULd9a22
T7yjlHjBsjERyk7ha4GVaQ8/6EM168e63eCGLzSCuo+9dS8ZEidW/o88PUD1ya+p2ujrRLUAVk+5
fAPytX9ag2nPeEF9X6n7k09sU+bCOmFNvKL8WhHRKD/RYARS4W/a018oS1oSp5kvYEgGMtGt1Gsb
JrDKcbW2zgCb2gVDi2NmIdr3+/aOe1cZEqLFnniVCS5Ddmm9YXBcPVmSxsg0P8gnBbQm61tgymnl
tLejNcSC5WwSAIClpgyFFpjCM3gFdwYfBtX10unsnb4U6U4lzbEPcsgz42w44nq7S+xBibX2DP1G
p52LXO1rejOyRnYis6V84MFyYrtqPaTU0zXQ+KBcpL2sKR1eqzmjIUWMr+gZz9m5eNJC4LGwAF9h
QATA3lZsTwGAVMX5irDT3j6FtHiKkaOCP0qCV2gH1ODm6SW1EZKTQTz7PPZp2svQlu4A3Xy753gS
1DU5wFJ2lc+OfYzbmHP5mZfcvScZ74BfVpR0NorOcpRon1OW87WeXIJmObEM+xG89wJ/vwqXBRfA
vp1Eq8TE61Kw04kR2cbqOyAsQtKGg1PjGEGNQ+9aVFtbsQDxvzTs12mkrVJb/ULSjDawGZw+aodL
8+jpdVVJbBCMO8TNVVkVuzW2xInK+PFmQr6R05rxK5eyF0WaMnYQprUiuC6ec+NtAqHXgLemP9hq
3n1fH1vUZeFVy1J3PKW9RnH+lPMFxAf/cErOQDBcNyytqG6GJO6OtxmiUkvRZwuk9t3vTan5u76W
QvxOFz+kmmjEly3rRyUX8//d1GZXo0i8EfUi5UVpDHnqnzv6zf1s2ZabXB8DOKlB9REjlOWzftSH
DerZ1Rc3c0Zue+3nqImuQ9NKQy3/UVZ6BBQZQBcpVab5XoJzjqitokWIvvnFGBBEM2ZP1cSq79L+
PHBs8gWOeWjSj3++Mtva9OnybaEkGqrmdP4jDZxvIvjFrnRMUzVW47I8QewrMWnoizRWlkL45CBv
CVJBDTz+0YnQZugjEfnY9kTvFWByGuxpnKi2Aft/q6TlJ4RCcYNIl+6iP/Qh2/0gAcKV923OzLD4
6DTx68LDx53l5uY722sLaqFj/w1nbNzsemqOsixgMfwdItbikJ+SxUgiY1oRcS5BUkNl8QcGnqru
57WKNR8jlulGDx0BLvp1Viwn0LAw5cN+1SVPqX006wZRDWerumbLjjYkZkOUUn/Nk9we3rRb9K/M
o4yoNk6Ch9d69BC7AqqbAhfUNkSIJ48bfABNwFhNMXD/2HTu+VyX0Cu/cd7UWmJZP6OTikR7RWir
weUdnsit6pwJ6HBZWsEOT6TNeB5ugNAU8p+PhqzMEOvumnSWvSIFMfLjDWsd2Bf8RvWpMoxrg5fE
tc7uVVZ7Xv5oNs3xXpSjA8ASw7AR0Znai/81aS8XyMqOpKTfmpXNqJoUrT+U626myOxbc4hdjpUe
0swgggXr0TqBLuVroLPp9229Jr2kjpZZXQXuzlNzfXPSovpaHUwZJcfRpOSs8aSeu97eFa9cAb3J
bUuHCb4E912xdin7tscZnUcV8itKQFQMjcQTt+tBw9zVrR6ms4aN1atLT1bz8/NUuRYwnlEV1sY8
rHrEWNzYaXti7eRBL4Z36BgwBfsOUEU6g+C731KHWmZJk2WFm7qzkyNG8sjCB0sluYv7fNoiiDvB
yw0NEfmuOhL2Fj6TuXRbAkg5hdub3MH+1fTypz3WrIkXZFNdhQXfjrfYcCWRwGpLb6ij3Oi1q9Nt
yg9J4iutySvcsGW/vkznGoCNyHmfdChQJBb0jZ6ClbaXSpDUVuoGCN94HQ49gqL72SSMrv8C2lyr
HVyymxAIofd3Wga6bkjh5ZUrihmIIooCA3hxbdqVnYXDbdkibqL/I9AEmyfhzaLcWtV6/xJ2pzOS
CtP+HSFaOKZQrkktpW64SlkAJaMSnkUJBo8ZZ/BmjiqZo2GF7beIw9t8J+2AvSk+D9JpIxkx8j1b
G0cwJnpQ8KghA5xM+De5PRtjeJ+mbfS4qNwjoLsMPdQDK41X5J3fNKvQpPFhrOQEAA100EnaI0RP
LO1uO40WqWkzutt3tb3CPOZIP0HU24ph9Q82neFAhdV8MgBGDaDUp9VJ4kB7saFSvRAjDa/g7xXa
RHjU/zrdStpb/PehcoLUaZHxgk06ws6QfQIO2L91gbtoOuSQnTiUAnSGRr9qew5ATbORq7SSKf7Y
gh8H9WffS4clW+Xd2RM/OBiEKqGv/xqxb0RVa6IRXrNyLVJzGDMOMLScoM98G4cDt+BleWIlf1sD
7+8YxehFL1OfIOxeLqRUeHYa0vexzdbr87S9k+OZIx3AKnu6FEG9/lm3xv3jNyMbQms4f00ig0xa
7KXaiyONjyeUsa2i8ARt91mmqAK0KqqlGgj7BClxEL2W8bgt5p2vT1OFELwwjSRyAhOnYXu9VQlq
klDVx/a849z3H2ABjwKKbHLQK3gFchlSzdBGVIQAdmG1AmFvTwACSW1b9+aELSfiF/A8KT02rgHO
p8tiIHTRAzUEZ6+LxmlCbKb1WZ1K/0nzrtMEGnZKD1mXBhHb2hsRoorRZrbHFRPhIs0a8fNSLBJd
mozCMbtRmLOxti/u/ArebKpL/W+kRisMrsqHaRUW58Y0MNK5XWh/p4FCgUCUq0SgvoFk2B+7ticR
ufWWSBW1JyclZIBhanEbRNEgLXjGLHUzupGdpslZV7W643BMz2nXAGBuWAeA53MLakPm2QJSIZqJ
rqqz4sUry4CSCL1Q5utlC0ryKUNsnvMK6x4Q+cyRL8MBDD5h3iJLPrPHEzhgaS0asSEVtfmmPX3V
f3eduP+6WZHfkiUmbf6BfPBkegG2NzNU4J8lRdd8c6VlG9l4GElvHwe6AJb6tnNbHJe+lPvHmva7
nx8MN/bvnzoq1zEzMR6LCsoSk36Cq0qxukuSEFHYZ4W+70SrBImnwWCfX+Eutj+JpSxUltgwD9Dq
DJNVWYPWtNfT9ZhtEFhEV5BJFglnrsoYHevf9ty3xwa1iC9sR30jAZxkIGufYffFLEUjv6ouGakj
LSzS1c36ZC5WIJur/RE6bbBWMj/5USvBXiFe5WrHCbBZJtDbQUI712LmuJ4RUl7YdSE+36MFTyYh
Kgvo0Uh3zFib5KFkSS+AZnMPtUEP2ujqpH9As7clE28tzqvDE0yF0htyvX57Iu6caxa9WxH6gFm+
ArX2JiCKANMRszEFHMCwYjnJpHjC9e4R8XWbEjpOl+88d9W83qj91ZMg6BvwWGddw8YS2+6AAbvx
wFsRrxmNFe/+ct5t6q45Sq5yHx+aE/bEWQ8JIjCR8qnZ21L9cVYHEhCgfkCimJfML3meSw2Rzpri
h56ozUPFJByCJqHhh37bYy47GOSZW9/xUdzWPkHFURsesjfCVJIhYrrEtw2Ze1k2CbzbO2nc3rGV
/+sWAe/zyjMuQo0OCKC/Un1wwGDkdthduoJdI72wrG26bOvejNR0waT/civElodd+TMf/WHKscQG
AXsXPpOQzmKia5j+WHdR/Bp3iG8ltOIVY3ffCZVJpaOZWvV9JKpG/IHeZzEaZ6DVkz4RDF81KJQw
8hNOlfDswkAk+fAu81du9zLtvCvmHU6gIXtZmqxON8rE/B24/YtdNiM3A1vGL817Xoh4+BXslnyY
yVBumUyLTDHi9oVZuGHA465tapYmTgBcFxVj/vo9PTdH8a3zWFr4ofLX8Oo6jGZ49ja70MNvcHbC
Spk1RqC3s7x3R/rscVEtfUnzQ3FLMq4v82rMRi8OMDfc9xn0bju8ZEwEvqBJrumJqxxqW90x8byM
fd5oIQohOeNT4obNE84i4x6GrWZzXkruU7aHQXbC/x7NYRGgBmMXcTuOQ6Obv8kYic19UOqbBSEc
Kp92chPgSu0HIGs5MNUdK1k+ZxaFdO8X+dInabjjW3TaphWPwEF9MpWcspzbqiMZj7mhctAIjwUC
r/H1di2X5bN+n4EUGDjm9Y1mxromv+/C5e9cIndOYRjNe+HsSqVMzjpfZs8oz7ztuAnJAHEjg2j+
6ypAz2cymr6RmINK7/c5dEALFudZAPHdXIgmW3Iu22Faa60x4q8a7jJkAIu4c/j1lwobmQ1eYYnm
x5zg1dvIpf4K2vKdMi3w53Q2isMH94AhTV+UFLjrCrzzhKFT30xL+S7ardiwoZK39UBLpxMLQSp8
MfwQ/JfhRudZplqMVv4aNC8DLFwT029/g3hum+G4Xotmcoj5y8iZhycRR/Ui4yMLtXpiqD45QWWQ
b7lS/I6dqOeLtZe+FQpqavV/w16JQId42sKwGwz/V8oGUw4pcYZ/rvTywWODr7Kz4mo1w3pmCv2e
x+xPa2WD3v+vKDyX8qxV1q6HOrpTfWbLYQQ1SNGJpQsq5YtVba4Mk07mY4OCoh41OGKn+Y7NkAbO
os2smKQLCli5LAZDSZI+XkEWi+OVWr84i5I2cetF4Vw/515/PLCYrc37LuafbwPou8ez54l5YbLD
VcTwSq9Fr9Gg1hzCI0xb32VDTje30Sa1H3QOw4NfHnUSrgf22lgGcn97qSF/9egvjra+4iBGVEic
390+nEJ+I9h32BwDMTRH7yGp+sUnNgiH0hx0t+27pLU9aodOvc40iitRd0eNQiqw6Kk01/5betMh
W69zjA5RZCg5z7U9oU38vU4ieur8UFqa82SxHi1skCksIIa+2tIzvUFXHx2ha7VwsFN02070OxvU
V48B/ZerOWUhXsWjX70Y6ntEnhix4UmYeUkoJNa+nMdRarnU1LogUZsAK3mKB3dDVhr5JbbFBC/C
OT8+Hh/wjbo4WZTUVNIsUbf7m/pE9lq6BhikhfnU5SScdGtSARS3EIaZXXukhUpDatWrciNjLT0P
rrILVz22VMZ5jI8QfIHnNeW4SkqMrG0e5v2ViCIweMv2rEbh95zStv4Nc6yGujWjotMSuihVN4Yb
/kd7AkoD5DMQ2jbLrk+HoN7+1TlxOv07BX1vAzAUCSttYzcr2xLJB4ATtgCAuqWzufNz6UWUZEoN
YddRA5+kf899Z7FOO8tUHLZeYigTmVT4y5eVoLlb+IW7ACS/uh9oqXfjId4DmNg/3EOo8n2pAqgQ
I09J63Btioix2HyJjbvm5UkXJZgT6KqM/kgvZPS7GHgzTQUb1S9Z/JRpL7Jlole2XxfQcaT0ugQf
IuIAvX66EUY8Hv3rdeDNLh2IosOb8WOO8DmsPacLCsYG5Dwtt9ySiSJK5Ls2v3vLynm3v3shI++z
00XgepLuLb6Rtow6rpGU+vL7wdP2R3Y+eTnS63SVIGAOzh0v6ZVm2zUio6OlGk3A8YgGWnh9DCPK
cLot3Bd5Icsz7Sv+a8BBzEZMfdQruXNWSpxXmkxk0oeOiBVAEfTfSqwylhZyRMGLd3Hx+J7QJTgn
MFxiQWFbObZ3oJLN9Tw3a9jIhOlaHqkwBgasEU5igRq85cL+rGIHnrjkfVWx48ehRCCtfTbvPpxe
inuL4sHLMigcxWwDfPrECWpuQaZPJVe/GiOBySKeppyJeReyKA5qX88hJCGgM3v1oGMB9MDXCGWX
mr6mO0kE7i/rblTSUoQXjACfLO0qXOPyTIFxeMb1Mtz3JTGypJVmMxSRduK7IhUE8aIyAjfaw92P
k82rv744/Rkxftt31eb5k9t6CAXxY8dJuDUX1PmDBXUBGwMjblrYtyiSPbhDh0Tw6hY3kP5grB2s
qDc6EBPbNeVFgq/kyBPXoXy17Kc07XFyJqnA8yXLxC9csWJeMg1C7X7x0CI7DqFU4KOIrVdSmARn
e93AYWPjxSuk1jrEBt+x2/Wh8zNV2/fnR41+rMWXN/LwzvADLoIwlg+Qz5gMtcmJsPELc4ldPUhC
GkUFkruQ/q6B16MS/MzR0ph2tahuNi7uZiMuWMD9UOR3eeWXdoJGTOTGNv3Lev8qWQCLu0xlKUdm
VV2gI+DoAwlpaY/DWXyhN71B0C0OjHqzvr4cg2iYWzGFz8zpW6/wmssA45gosqwk5CiK1d2hm7oq
t9a+R2EvyzOXbRzO4ibsMgUPB2Gr0YH6xwlu6zyCgVGNG12P+YOsHn/Ixe07vmux6qskKPaksb3V
iw4q56wcnFaS+oIa4TdjVRN5b5oS2uHB9TKRZi3UQmIGQZcEb0H5krwAHz8bblPw+2eu8/EBz/wv
7RoALF+fs9oReLHILRvM9cVGhvDlv8+SPC8kPr6dlLWYAOtDVGLbDd68BChW8jwK4m8dK8caSJBd
lpEHUkBZcnmS/r7VHposBSAIukYzMMcpe4WKMd0L/hAd3FZqD5+DqvbSjdsjeOrgqVJHPbw75P5M
vGJa50BhbOvzAo3xi07b0xA+/jSkcUeEzr0v434MlUMcjfyGWaCvpWd89m8IK8n2cj59swbhPCzB
C2I2wg178tbo8k0vACCLieQhYU0wqkFrx3uv6gi3VQTiCxM+kSzqLohUSJZPbiCX/pba6TwjLDT4
LUerfbfDsWpjnbc+SobuVfen5Tfil7BFDkk6nF14PWRjmWzSwAmzWr3V4Py1gWr5TqGcbxibK/0C
etiGt0v3L2axzvjpfDmvbLmXlDl+fXsrq1SUIyUrZKaoCR+fzkOYPK4cCvQIhtpvcB/gs4Nfc4lj
oZsM7HHOz/iHX+tXXwI95bEGpNt1SUyzO5AEl2uBdYad6kUKREK7QVSY+w0Ke/QSD5Y0WyEl1kR5
F94p20ch8YMmquNAGSw0pB3zCcbesaLhKvxiDYUsFgs2ugO2ht8FDrY+OZTBmA8iBm7GwuLnYSoh
7yGD26Dx809H53QzMvee4gOdhr8HWgTeV5MUsJfzdeuxHEQkPBou8Z+8rfZfVkmGk5HCamX2zPPk
PRDu6pogdgLq/iLtaigb7xyAUnDfp5rW5+f5ztzhN0FQM4tT0Rgnyv44p6w2wpBJuZTkWXWiAvJ8
/3PfB/x4aQAE/lvBVnYQQgGflNl/JRkGK63DNUBsUws9bijrpTy3Lmcbn0F6Z6hyhM6Shw6clBoC
dXyFBvGlQVC+q2MMfakWs9TfQ/Oubw1gha7T2z38xgVPr/tdBZbKgMfT18Ooy9bop6C1+JzVR+kc
IwMU8HcDFn4oNMp5sTTHGDJ5iJSNMpVdQQqjOb3/9BnpVF45Y5Mx9Sfs5FbhZScLvWiRViKM5y5u
Q45UdpiUlj/T2Q8WV/6u+G/7X586NWh6Ep3CJxencYwBXT3uUYGcK1Q8qBK3r6ON4iyczCVsXTlQ
U1cET8P/FA7Mp69q31Y9DqkQElKFW0fqbjhx3IdAOAbRMV0IbCs4WydVGBiKorCiah29yRGeAUF1
xo1jrACCpLoVhwexHi1iIwSbO44++GRMsFnLcmi29tjbZYwUpTj5S49nVN19co2wQKhqBSh3QPMs
OsLMP4cJCXgccp6BEfycaCr0WlTooXNmSofCQcWZZE6QGnjFlBDd+6+/a/VAy6EpbIieasw2LQpf
APwkl/wxrs5fUG5S2CNP1nPtDhpv16GiaNI4hI+t3zV3+IP0iJPbVTbIoyzysnyglQU3tDsJT7di
qrXmKZlXhMu8UuW8y2oSdEfaL0LXSQL8ZwMnSY+cD25THkoIb+WWXm5G6nNMLwILHo94GpYrDAUG
4NKHiGjsAiXK186F6pR47WjFyhb2KfAA5ZZLWuTZp7cwHTD4UXQwA2QdHe0pxi462O+BHn+FXpOZ
umSR7keTzAcNZuGED16PeCcsFOCGZfJxWCi9Ztbwc9/mfMxEaDkNS6DOgHSHNO5CvAnaHSm92dOI
wNDo3q3g9DfoWkHS+x/KUEcD6fZzhBAkIYN3xlsheEhMQbQZxoACOMyTspp3A3SI9x8A7WykfGKE
s5WcNcf8O2UNQCpiZ2Qb49B+kq2y2r1qyMvopWVQN1sWtlNwH3YLHJSLGe+kW7pgMdWn7xAQuurx
IvUIu4b6GygGksvMB7P1MJujAmaqhzo/XcZcMIX6IlXOa9l/tgZU82cPVlFf/reibAfHrBr6/m5y
gkh1QMgHizYUuzDXHGM9yxZ9Wm7tni8996640WDJKt19axx0dRsXemwyiFvfearaHKy/u/e9/b40
8UVYUTlpoOj2SB+UQCWfbNfldcd5VWspjXChFobnPO7ZT/pi7LQXg/5qCM/3WaqAu6Hr0D0vm9M7
/nzGNARDI/tZk1icQQRub0HuNVIFiGS9TizO+9h6+858Veta4QWG47dyP/jgNYYi4rCKxTfdM0lM
Z627BXETSFkkGUeu90x0uqSEPMv7MVwUtubVDxOPDFEJkgpqaGneLMygDTJOFAsZ8gRYkmWQstVn
ZVijG8mHcniFoeGgZQMmnrmKayMpwtJQqfyHUgkMNp6u6ZDRML9dyFYpliyvTneahV+MalYs8yTL
g2g7wc9gK9BqlttYR5ztgrbPD5BDb0pOIo8n24khcWK+izPKucESgRq4Sy3MiOdpYLMmmIG3J+zB
OYyfsgsVWFuYYX9x5oZuZyLont2NLE+k/2UxzhvxFEOUEcPd2OgdAMRBE1t6JJetlb0fD58pJL3y
0km/vCJeEyRbLdQ8caLROvyhOt48Kh0Mu0PbnEfKLn5C4rKYyeBIhb/iIgtojujcBFqv7JX0hO2T
x1XEdrP0K3qu/1A5KALDtgYRs5GO3taPSWCXuN7oiQ1TB8llsKZTDdSiggDsHL1tHWAX/5ujiZpu
Ec/cDwUPOqMGs++AldG9PHNQBaGtTkb/Ox+3DzpI4XtjIzV0QDgHckE9wKwNHg2dMadHhD3Tz6Sa
WxUEHhM7oKgUf4oIIoOFbsNn6K9WdTt+DTmJglAwuQsYtZm0fH/OUfveC+JkhPEiTUCu/AdK9VYc
NFd2g7bzag+FUZ1r2h7kA2WYTysi8ZWPZ6IvUaF6SUlKlE6+TtmtqOX06DxB3YAZS6E76m1I4VpA
G60mEx7Qg5qDdF04Zppw9peWAkb/082zRCFFsh88GftdgTfS++25EX7GEexFwspufWd5YHV14ecP
zV4a9xzRhU/96UK2HmNOEVBuNuSLcIV29Ado52LxcIZJTBmhgLIwcN7v1Eet3dm7IrJV9IHVnBL3
KWdDY+V3WOZ9UsOOM0tdMQLTvlZcpkdIBts2yKVepT5d7E2dgUFOX6rgEzKTTA2tGS2iX1ejcmrn
VHgHLRx6RVLNDLzu9KLRCla7snYJ2qWpp6bzreplF2Qpa7fAphUk4clAmbeMmtw5RBUadaz5nJCx
mR2FETzp+582pTuubNcwUjG9pShLC1Q+c77ZmlXgJI6RXdoptk3SUbbgtnaCWdtVPiWGC6NbfBUO
1k9FIvEWBkC1pEvZDkqB2KzVyhqqBBx2DBxcZ/0PjmA5f4wMH9UOGzHClpHN5Ls79CgFm/ioNt/+
mlZkmkskm8Ar+XkinvX+Tqz23BoDrk3Wlq65TJm/ks76nFzsZ/sR4eolKyPxwFWENI2BYCgyoI14
L/u27a8rsXuNOedcSNcSKBr3mk57rezIpxs6dJZnyyuiiQqnGSDk585AWIN9x3I+xUGonp1tcFzA
qBeSmW89gyEFj3pzpII7vsl7AhCfjN5yWEtfjBdoPMDsHQuvgZS/nST7I3EUVUxIkdoSXU7bRlQx
YWjsQosUFG5x6mrSuDtl7VLxkBnfUU0K8NrOUvkGteh6/9KyWG+Fh1n6F7E38r2kAybC68vvz/L/
LgHrm4+6jUuYmvVjkUUfSAbfgr8jup8ZlGaWbSXkGtDsh45w7oxVBOQ2O07JWDrak12R+9bK7tTp
uGrgeY1KeZbsVkIKob+pcL8ddtz6xEVacDNVIXgM446beeXbuHsnNOl7obRpea+rZtCCsajzTM8u
TJueZ9LOwBzL7oTxr6zkkpMKDrp/0osUDafO0aeEsQx14q/TAeg1kwdgcTWvZbHt4DokSrHZcLuX
xa70+j8LSSJbu6Nt3Nnr/bXTI0Lj5TK6AXc6vZ8UVld7JA7jLPvvYBozspkVjG9A9VIpfbBgpb4S
WwPyUryVEqiw4tdRuZ6ibSEai89xBx3eN1TcYHyjN0NUMygoJYf29yo5EID7WihsYkHl/5E6xFAt
vuw7BuQHe7l8yA2XjpkHvcm9lb7yc6f5o7lB2QSSh4nmX7qvrzFZkg9a6RS0SB1VMu8r8MMsHeWf
6Ic9wSadpPlRD9ifuXXMT3t6NruYDw4HlIxaK076bDa4O4Ep6NPvB0MxO8q58qYxKDmPyPlKylC9
BUCYMsmFJyMZRrbVhKZ7rC1ps2sqF5RSopcn+ZnRojhgarDeXyKKlYzC1JDlq1cItYNtdEzyNO+b
Fbmc9fn3x/Ertqz4dnVL5lgQmdPbKwZlqqF6rbMiIlXSs6iwxJCN9GAYv0E/lI0A5PtMW+3La95B
cCGKlWRo4YuOpccuB0MgfoPwP8daLclXbTHybLW8QIQFyNV1NWXi9nhrKMJSElJ4uXW4Fla8zUn8
UsAMnSiCbvXbRqzeob3IzxC8QyfHTLuOY1O1FQ0bTl5algqLW8JYeaIkSVxF7Luj70d4K79jO7ZK
8aZmfnXW/krP46dvNyhCNBo0nhzH6+CyaVpSFS3sAoMK/BPBP257WVqcb3CwsfsL8PskAbaRFC/c
/1b56mMdcqW88uq/lnnkc3K8W6KtzoE6oSsZ5LLbBp8Qdi3iLipe2+sohPnsed4Hth5e+ynzjmfk
dxlnaUeG6UC2ElSyd/8bqD7bdJWwav02BS7nrKMSHQHRSJ5phmDYAlVsmr8vLBRnAdybqy4SaBka
jCH9bwWDLoxxTpzTdisTWe1Q78cBfp8J75BdzOg+ZEDTCmqfZZoJaZ85LE8IP0Dz/KslswmhJdRo
OwvbUP+SImSY7efxRplsCm4g2DYdkf7rrdliVck3ebXIGtTtRpR8/7EA0qvr6991IvpWMwbvn04X
snpoFfCwp/GhImrnzKlMsYCqp7a8ozXpIYMOjuMVx+kbZO4hdEIC9gd0J5esM++6iMosMyU4mvnl
D9RlGyAd9nyFoOV8wohEsBgno/GIKHia4pCdZWgWStsF3DEgSTw1MZI9om7G8+9C1BBIYaEHwfrM
MfBPH03gQIevNTfZIEk9uRFv6EKDG7y40EDJElcUNPy3ClNTU0DXQ5e8SXnE2NO7Zx+3gB34UrrZ
hmnwhhtw15SZAtEad+h1WLv73IRdx/JwzEES0TSzndUC1r8Jjzpt4zLtDwdytlJithaJMd0cs1ui
FFH03KZSZIKd0/E4P92OMRZJ0KEiqmyD1tH1znqm3SGcdjnOC3fLlK1uUazqvmSfs//t+OslmHj2
29deVZzMKxATneHre+6J80K3zu59o8SlQPT9IMlgX6d/Rm0eLjaM8YhKcM0ygrsL8+9eYkZZWvxq
R9YfEneIva6qEZ4YmW+HUpeKzONm7BvbXp9Q3/DnkDCMpQxeFlY+gVWA0LGo3PueTaQ0t3WPjRyl
Hg8tFXA9KgMH6AWdEK7xCZ7WHy+DMzNMfdhRzexOUyd+Hbyw/mfv8/NQGy3ax9jMrlg1KaE7ERXw
UMGWUQmg8DmMISQFOmDfcLOalW1HFFGVloCktIwTgIqwrFg59ClAfyK4w9Zr1SaEQRGbJfPEqkIm
jEbgOFvumP4gtead9o1udmD2aAfNYUTEYpt098Yplf9mfqyTdUit427EKM0lDkmGbnzOo4LjLIEJ
d7fV4KWCqr/XVOplJT7W5RWuv+IPgq9slEQ1Yh5Hga2CNKY10lCh680nL4rbbdUBXAuYuz+t38MX
W74fRpkoCxhVWWGY+uN8fcD2B3ELJb+rsM34DOf8Tyf0ILTsOSCcrX5AAdwEOlsKDdLGeeHgs/fF
SXd7Kxrlfx7mPqh3HaJB7YTG6ytL8St2QHS9xGC3HsVomrQX1sR3vcJgAhqzMrltK6vNJeDTnZ7W
BFLry2sqvUnWHGTsBMcA14LA8VeTZ18xLApQ7UehsMNmdrfb8/2/rFubcYA3j5hIyOG28nx77DY6
Ive6kQWN9uHLst2hVNv0S8YQNB3mdyb4WUZ0AC8q72m2091r0P1kyIGpMEbTDFWQMqDMkhD3lMxS
CTYkdolLqUjSWRKEUIT3GxJ/JudbqtbMoULRUMt2nm5yWsqSpDfngrLzHoCgAXVoTCA6+pare/fh
FBybj/65HqMrUuT6GC5yRPEE1znHkRGpckqg31She+WrdcBVqT+DKOPv2JtMSJ5FLgwdVmm5hwyr
4U1JBpja7cBSVqzV4mCUAcvh23xLU51lW0iOUcJoLTTFTVdwMRjh8GJOC7IR4ygYthUcbCG2xEMr
/VCnv1eVZptC4JJsnawge4FHp1PZA04JItJlIx94qHVmrPQzBuqt7RwY1MLDOavJR1pLC9KeIcTf
XES3s7NnUW0f76ZP4ItIplT7C5wwVU97P/Mpgp25Kd9qCKEU76ZnpHQf3E0RFNpisk6GsOBRsFRi
hg7aVwqV8XzmZiMzWEtkHc3kJRoP4htSF/9+6MSv/ysvdy4s9OYBS0leNM5F49MohZAqNETI78//
WLDOkrCuoq9BnyoctoFkwtM5hQK/xcfDPNeuSp+tS+WSGKZLFCRcYRGuV+7XIen/uxTo+6nr4wn1
p04U0TwnnmAZurlzuLspBVQ+39vuWt57B+Qo7i6ZvsipVxQCkxjixn1xIlUB/BtXeWAW3WPMVgGy
aIxjmGpuruIODE+Biq41FU0g+BJtQiLfYaCD84+Cu0uEeRZrppQ+HfZxpSUZ0b+pBPOHL7JOduuA
hJLpH3sXR2UZZ8Fwv2IcnDf9yygMe5E6cb9RKRXuvMVSOgLzdMXHUMlxQYb4m3PaQPaXjT/mZIi2
n9UFdM7Poq+N7oMI2MiDfQnF+9xyJZ+zwdk0Lnhtr5bMyEmagJuUXRkqnYRcpnUFJybEv3UQLUWx
w2FiXdGBnXyXcBtnBVnQ+AZtQLLxUX/3XevkaPcfc9oZVQZv6+I1I1kaiywoWquIWwCZ80xMA1KY
Hdyz/RjU8oOsWuUURzV+20vAKOF3UG13YQcR7GXYH0oEoDoiu080cSVSUwfQgMpeqUFxSVMvZC0p
UxvHEasz8Liu5v4csnH23WCeHlt3OEYTtzuPjxkLuueUS7qGKeAPLNIFNjwHWeZ1Pg9lS3qJw0KX
Z/FfhTnT2c/5l0Wb7m7tRP8yULjoELm8WZGihRqPi0NQ+CcqYkCzihSlo/hkDj8+XMNhCqG6s/WB
kZAcJs+LQ+czGp/j2SWL/vyHIKXm5JesHZ2sDjDtfMbqEfmKhjdPVa99kUJYo/UiZo76opjqw/zL
cVfaIMRbOKaxtQllwuUPEHx8PSQjCyZ3nFFIiukReU5zO4wuBSCdsvLPLTzZiXfmKiqddu2RbieJ
Z8yc5ocS+oVO8Qv4S/K2kgW5BVX9V5zU/lzwu1XOKVxnFgmtRDaWci44XKwh4j17SUc5wZpUJX2a
pUoSW3aEFI/f5Rzxw6DrMKR8iM53saK3lwLAP+ppDhbm1eNmfoqtM2Lxyk/kZ8b2Zi8+cYT4zjsR
xEcgzq+6fkv06qV3R9asDl+3fsEZyyvGFl8W07E40MpatQ+CMyCyIdyFMS0Lmz9dt8ZfUVykFJjB
SfsUWv+mZFttGSFDz7+YM2Kyasz99+4gN2UW6sH2yET5JgmVEO3ReFNDgxSr8W/kfxPVMZSO57UZ
Mgki3OKC/ba281DD7Cv9j+KvKMqt5Bn026zsby1XJaALXM/o59stA7stwLdhdKtzwXIGGWodpmIt
J4CVs58iKCllzOPaR6JIfYaAoMezf74ruENZTuq8kOFMKvhG/hO5d12fvgUAiSGotay9ceGoorMk
7QHuWLGHkk3PA0Kgoa0n/coVZR8cpYLSydewWwn7YOK7Fh9aqOTS4Kil2Sd1QjRwaiDOaDH/h/kY
b0zIF0pwnc6vYh9Cs/auQ4q4q/ljKEF0olxY/v0Sf2hIWbUZzDLE3JnHWVpZQM/UKtzBcY4lTsaA
RlaHcZA+cgmQQSMC1d+9K784Ky+jWblSZj9HgZhcS2I5ESD9ilpFO9T1Nt2XjXVxlPyPeuZKlwQ9
DVdZD/OfJiCPtiZZq3XpzdfwMxST/pmxLp0Aln4w9faeIL1vkZrSvOepTyDErZbwbjgpOdU9Euon
rQOqUO8mJsF3hLYHRiBJTGy8zRMrsQ67mlyvG8kXZHZhFaAkyBTR+pwpDvqsfkGU5VEWCcx0FugD
W7WhH9JqzD3Bnvxp4wXHMHLV9h3gjsd/S7cT+5t+y48lO/7BXXopZd0AWH0GJVf6yFXUEs4nsH9O
TfVzydVEQN4+PjkfAw1WksxgScIWtuX/0A9IklWxHXQEtvof9glrPhXRN6vfgf1/QuSBdwLLO0I/
3cd49bzJMIJGwwIsf0c49hLxA84gFwc35+Bor5uOZhjD0yEjMoQjs7KjXbN8sEW5XRb4Mf/NVyNo
rbspiTC90jxcd9lahyciPLN4HYQsT4K6RvBGRX5wBVux6NXnzVPhcIVouzvpVVQ39jvkZ22F6ENo
mtMNLrdhS0auXBWYdJsi9MeX0hl7HKdkSheeGDUeERGeRtvBa4BpcEaAhiZSTsR6K3LSobx1PUzx
LHdYTrFMcUpc/x2s16i6duaCkgA9buRe73BfjSYzzFrRuE/Rdt0t0viaA31+U+plzvrp2BfacaNV
IOS02vM+OG1Uch+OmJ8xvdhn07DFN8KxqCw8mmkAvJbCs4mT1aK80VnI2Hsy1ygofYAEwwHE7elZ
JqQWdV1bGnUm2ItQeqiBg/bltLWQQQpQf7a0FW7xENdhHITjcynaGWDrbpo+7w7FrmH5Zr/aINSZ
rO5SxkwKMmZ6SANFPpXSK/CG2brHtqaEggv1RH4BGQPzzVvXY4MTpSjJs7lv3BS1NYgGozU7lEgI
w2FHlS6x+P1wZYfFDcLyf4tgiWJ4ip+OHHEckfADcBFvyEBQl9xOn+tKLQiwMg2RE2e+UuwzBiEF
QHEqVkcxQQE0rC48F/M8yxkNAyWr29dAGYgpJVE5tIzLLWrifLYuTXZwd7aPhr13cjJm9wwomnbQ
YzbNGjx8hrGqLHOxHFSkLa5XsYCssKAusBK0coM5bQsuhKCbqMo5L7lEbc0QSBNmjDdKdH2QNYPh
oLSBRBtxNMHMS60AzvRR64G6sciviPDg9LlxDASZYxHqA4WLPKNVrgU3H7+582M+CPER5jxljrXN
L8wT9WxS3Ar6fASCC+q7Uytz6TQTIgdAxuGNVsB4kAJEbJa4TTObErF4RDiWtQm8JcDBywm/iCoJ
XVq0LqYnZ1/DuGu9bLr47W/xUPfT4ltuqMr7/H9jPEtiyDShipptvg4gBHC3F90Md4EO70ilGwE2
2wNjVWKMvabrd8iQJo2jY6yJnYTRc71LflB4ynUBswMmUHhqoOYH8wAjP53yhCH/ATfO3My+O43P
ZVgyiODmiottYDva6SZD2l2CShAwvhgLYpJJcCxr7vVt67aT4fIdQIIKsG3xTX/tSmAXZ803Th9z
xXprhK1KXc8ZPEsqZf01HMgTibJ8ZMa5Db+nV+NKqAZw2Tld27axGgBdyw3ppkL1CLUVa+vb1v7z
UZxpFwcUzizw54c0/Dl3MF68k1N04PxvYa7ztk1TQ5qKSAkpe3E33qRGU/vDW3SQpO3ZHqb+bxx+
BzVAbW6qrXb/HNWKTmUN+bhkO93fxKAXhRCh1dF/pcmMpX9WE9hwLfolXFOP1NU9UtIo0fVRHMWt
uXP0y7qmjRGE9JPCGtQvIJ1mFNZxiN0L3GuQaiFFpi1qEwAYA6FeXdh9XVVvaXpGMJTVf32s2PZH
+e7MPWBzzVvw0p1reSM5ep2xV2gyLuErA4RVhRf5rMxabxi1uHrE15XyCWsAwYuRelXOCoANuIxT
57eSbrAshqhHYgWtNWi66j/NzO0hajcv5/4lVBzq/WTa1EtGD1botrB3tXrjjH8/LDVtn0CLOCGr
iQ+tYg5kEvtUh0yYLarJNnXZX5lsXdgNRoEq7sfGmS3rhI7PqREMFL8hZaLk273AhAAHSygCAOii
yK/ebv3oLho7HYWK+NKs2xQ9oDwzOWgwbifcd6Lazy55fkTvtGekEYEPVbO/icU8I1VvZQ82XTFQ
bBqyAOVCk0ZTLxO7xQ9eUJolCTQ/2iM9/X8jcEShM3LrWdxkd7uI0mwOUyrSBrXYEJnIBnMnBEa+
sa4hQkgc3P215/4GGoMu7E+2MHohAwNuYkVj69XOgBBvElN1IrjwSvOJqjtYd3QN975KYumerfXA
X6Z6E4KDihAsZBy41X61GBMDB1BJELJjHx/K2KZ+cddt29Q5EWc7uTTRUSDNZLGM3mDVsuuIMsLW
VHEAW3jAcmYyiE0OpcJg2n/7yRwLnT9faQ+ajbTUldsQ27nMQ+t4W3TZG3H3g+1gRRO6SuNKlyY9
bQZ/X0PDisdaIlQPaEhUchNZCW8n0OSk42AIiE3JDDBf+sMLN3Dn5g5I3W1pkaS5byVVXpNFoX+g
MeLeEed2hbE1PCMM44EPZMxzOJwmLaDro8/EHF8M8O8hLYU9mrBfDNP3tk6rVPyMBP3US+WlxQsE
BXfsQw2BQckKGymRqeJSjtr354km/omzbWHwDqu4iUMTwBu+bGLtw9+4Fvq53ginHAQTHPdag9VC
+One1Qv3/FyHmxCbo93BjJWFn/K7W1xC5wIBw1VTsnGbkdvqwgjnNVPVhOKOVl/vbGSieGuEpIUS
fZJdUc5Be4ZATwjys6tfU1lywpTMzyDvVTwm8ZKmnl9K6npNJjDmVuK/P0qIoUr1hKIQYU7EPcBD
aHgTpjJzeMJOpCNEMRlbHbxblVWxYzg9HGHiK1AhZzHBNC/V88ALpvimmArfsaRIdgc0oDqBXmvt
YbRvQeEIRoqytW4FYMQCNOTNVcz2XZQou6PnZAnS8y6h2MsXRno9eRrm26JmW6nVkGBdf/Tx7t+J
339mO+RuGruSvwGeDBeYtaopNw4yyIoPk3E2R9DWdulkoF0nuPiKIoogLFgqZTMzNzkNhis9Ajhl
qH6zEVMv8TaRUKuhstel94d+nsOrwTgFJ06xtxe0O99qSEHUOuPdHgWGS/L9/RVjbVdshtdlsvbC
J7x8GfRA2UjRsZiyT2BEb24QN7BERTKRsV3jxGP/Gn3d8qs8ORqv7mUpmzu4q5e3ug8xkD0xteU+
HK70cxolYNSEcfTzpKR1pNQOboUtJz4BUolncKZCmI66FXVog1M3pY/E9VzYyr5QSkP4PzxGUtzQ
7YtKoNGlUvssHklBe+G5jajzlwkRSRYlhxZyrCgs+Qb+WRc5nyxEf3BlxGXYFH5qajafCE80OitM
hABLmz/5nsyN/ovNg8pUq9tVosBP6MZS6K53EYKzUiiiXAy7aByvrvJ487DEi03CYHA+yyW76gRk
r+9VPAfiKY2zwOauDCqQKUqpf6S+69EWPrt9HqodPMDpldbuHLSa9TwrjLdQy3jOf+LSphFOQl6y
U89M/MChqvMPVJE6LZ6VJqczMGGgOC/HMLGfsA3voEfOXnUH4OI3F1S0pzpUAcqjYvTQCFyMIPBJ
DGDmBbWO2uqahG01pHvzAJyuoWKxXprYw9Aq0gUM+Ila4JNnm6zq6QTA2TZ4I19SeXO0bb+QYnXz
HQDKhHxCzAZ26aHdwynhv7ce9Jlf+e9VfVmKsMAkclBk+/NU/Hq+Gp1lmay73XwpsgOXcbMZbWx/
lUaK5x1+JrG0NFONw8/QPMN/o2PEShJsUodaP36NES0mHrYH+0FekYJHlFWGWQEKsHh8hHXPGfc3
OeVwHtRpzgsdNvsvA7OHDXoEI5BaoYPnHU8RAkXp12wztMo2auR2q03+olD1Z2hgxCRnNNIVUr/9
PvjHowMMwepOXYlUkl6Je+Odqdf/mybNzw/Fe4/XYnyL/W8NRcyTn+WotoP1wUYbE25kUWDvlTql
WwC/avX1KKptZZgbdZr85/937bFeVNEzEfYuVHWQKWAzk0QnSmU3MrkEtyiwBzXX+Pxj6TesVeuf
R35JE3NSDI8JBNM/jnaxkqyw+9nwY/WxbD2cTZhBLrl1htSNG3Dy2ee8/qgpKXn5wNfPQ6Z6p47Q
in2mzhCOUXakE8HOQGK7nIHAWNiIOghmi0BADloWJ6TxUMwY03+kDL2pjbjHEl1YaqO49fyBXrvu
IMUECn1LiTJ9f0ffrkgpIfl1zYCbvfREV1j5TJs6rDCxioKt3w+np/lCCHzyLeU/db88WtKBjdYX
1Vna6/70abfyUjJwNDWm4YZAciyRro64Yn+8Fy4blAR3xGKd8ti4gIbxav3tl1rXhJO7hcf+2fXV
4qIcXKPfA7tkPo5+sBfq/pYQgDQXZQ5d14E3mcMnSCE7beFzZfHdkqtypSeZR/ihw/HSccNGElhB
9kDT4n2E3kGmD9Ahh8/tbkQGHim0KXmoYraZtLT+jKvgWD5iIJ0JFIV/dzKJtjuEq0pL0NAJc3yL
iRI+Vn9b9L2NyXr6C2IHq9rDl1aRv/lCy7nE4wstPeqbnSxEI5rJ36ucyD1ilZWn6UEzwuVfaBHs
gSiStLJiUmor13Ga+/kWybXOrbcymAhH8M/GsyC3BL45f8kOTAixzh0oIuGJIytbqD/k3rFHFys7
PvfvGWzJfQHLbcvX8VTUbDB3AhC53VMft75mEBMVx6LKy6G1QeVtjG772ewYSB93x/zgzhPTQHXe
xEN8twwYSzkZcrYIA4zaoQVh2QmJKd3tp3xiXHRIKItu2WY7EksMa0QVEYi8bfNkdQZqND1pvI0S
chQ169BL7ulu1AmvgHXXrZj/JJa2amem4iZS+HiQjp2+Ljxg48LF2UtFVlhsu2NJXUOswTxTIPoD
IxMWzL/gI1DFl+ERAFJmZPh5xC3pC/Rk5w05poen5ZbqdVMx0f+UG6IM4jVlnz/nfALW0Hxm8+Mq
Yoz1bgp+HtmjP5AGZwSplGDaSxtk661uqL6C1mvIGKezWPDw1NG/3JHve9F29J1bVEjpcU6aXAHU
bs4atcQyFTW9sqd7Him9hotU4V80z2YEDOfQbbIO9AtVjmDPibLKsLaIShIl9SrKnYI3I6NFc/XT
TypgOq0wPuzyKVHWrI6ZkCJOa+m53HPaRg6HHPr+5zg9YgRArlWo2GN+qLuX6EqDgib8CIydrjMs
e84QeNYSl1+Asj2HzS3SB3nnVsPq8T3hu+1583hTnvYCfWBhBqqUvswg71oBakx5P01/nqPUEVjA
V9LtvshSImURquk9SAMi04AM1lokJeMTb4e0X1ss7nQrfxB/ZAWKTIovaGnd6P+F12GhF9lMsbh7
yEwMIkkt06xj4p4PHXrXnlnFJHnjdeO6WXcdhD4TAaRqU4PfjqBoiYv5kHpuQ6+Yhy8TdW40/q42
/H8ngpW7ZseodtqfiyzDaGD+EknyfSdz9ZUzop9NNZGEAzk92mnUgTm2Mt+a3NnybbwM9wI2ZL2E
iRCcKNPJD4+QMrsXxpa68vytpSWMncY2i1i24sYXzSgxoyDHAYFRiRGxUsSzZkexI85YfAY938Tg
jL01NdLLmZrBvG44B56MxsCyYUb8oNJP1jkKWgiRsvDTChywd/jh5qo01pRBWNrPFEUJbGamZORY
iNYv6UxxbDD4zjC3BBNgHeDub64Y+UpifnCmt0wVj7PejDz3HT2vuBVWcORZnd60JpPpfv618376
tMHLyJRAClHk/sZDBcvav9TGdxB0Pi9Wk5tj9zrxGPn0oFaAcQgFhGSbFsfWToYfudU8WPiSJAKH
nVTljTNsiBWeXNYJoFxHanfy5yeaAsH/gPA4s2uRedhV0RrdMJZvyJ+HyoUGJCBuvO4+i6gwJut+
yh+4NiObHgkWK+gf4hgT1+IAr/tXHXXrR2DT8iS6TVioPvHHxr2nKKu5Tlw+kryIKj3e1IcSho1P
4osNO/54rxBDFXkH1xJzu77duWemc+DYBdaNVN/eAGbqY9ZQ/T0Iw8eohYV8iTya4nZSGUAsm4a0
v0YBHqn1RreWGArFLGAG/9kuv4J1DfT0wTJF4YvQiFwJHPmixOZPuV78nBexryJ4pr0auqML91mN
ukPHHc0EWTMTNw1aSupKk1zD8C9lW1eVAAt1sPy+1ERE1HF5CTArFwSWsZ/4T+iEs7AZJTacrEnz
pSC5PYRpEgA9xHscX7N7iwgh/rhGkpr8vzn5mIQi4iTfm3stw0Iycklv/tS1e+Fq3LIRtm0EcLDB
M63nz8ZnVGD2Yq7Lb7SngGLjZ83nrduk/ah/1uESxKsEC+bAJK+1PmMGgxe8m2HgjpJPUhSzhhFi
hzpqW1BCdS2IjGuqnCJGYPTfYCVOMF0CjAJCbfEpFBL0G8x58HyQ4bQtPnU580ipBNJlCGGHpRZ8
Cc4rBY0uFfQeFEs8VGxzq19rHrBSIUc9hkG1hnyN5KbqgN0EPS5pRJ1+wYjj/4EfgXkbHg0bo6qQ
+M19WJuuOFR5HZFiudhUf/PNZJROhuYGCqZNvZlQhwMKNYebjq3VhnayhQAx7hYcCaOB6cNRd6Nr
nKPXsCC8/+TOQZUEsK2XF7Harbwc0bfNoUB92IjmNSMJ97IL6WEhhJ2KDg3qf3EiIU+kuXNs4azz
kI8tc2L2nl7LDuHTgC8aqYSDNNfMKURqxU2fRFpP8dZ2G7WzeY/VeVEecAW+jjExQ522b64e/IhI
g9ereUQ42NFGjB2cque0j8AbbFcjCdLj8tlO8wyiJ9DU22T2joOHZD1Iq2Kp09WRZAsFb1ZV8ts7
cxZKCQQsmxw/wxDasejhOjHjNE+sbuA9naM=
`pragma protect end_protected
