// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:24 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
h8KPxmblHxgE+/qhiilZf0xIjulxEkaYvnR8fODEc48YrlK9FID7MlpdUMWaU0lF
XHuoOi98RbqWj+cmiecuh+4aK+j14m74GgpW7aKIYV8GoGBMm73kau/63kdvpvHz
xmnuG3tItAuIRlhyJTfAclBhb0JBdwsrIG5xG3C+IeQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6320)
2bRIRUNbkVpLfLpxnlJtrIdN7kUHcWShapaCfhzLK1gPFGaaUBRIo8WAXzhZ8ARv
wbZJtslbf0ZWBbBtUuIC30ynBIAYoIBOKQHpdQY7r48+PKR+xGrMbjUu7971LjYu
cCt5o9UUUCCpLsw49RHGHmCQc/Pru3sQgaJXKSVNwrz9tWQQl4leRFar4+lI8l/8
+DvHjC9lpgFKyNbqfQnbcI95O8vsH2IhSexMKWaEb1Hmys2x3SlBWs9Lno0+mNnx
+vCGyorMre5CEoskNs26E3uiopil09kdTY0WoOCWMJeL8ycEQi25JTOUG4cIiN28
QTEGQCSzEHz8gF1Op9DsGZayJjX2o6JkHT0BMJzDHGHNMRrQVbLoXM9R53i2imf5
pI/kqbnDBxRPqsoCo8VF8Ri2nrcEpJ2/7uq0CD32rbRndy4hqB/lKLynOW/i2K0t
Tipz9YrvVC/Kz+1kicF0iHCDW/u0BeOwmpnIvqKe6oBJOH3VFZUfT5crLkWmzvVP
vPzjWxJla+V1sj0ZduJXKBSrRoNj6V+yHehIUOeiJtNClkzllPQSXiX+ONySYWG0
1HBBRBFWHyJ/xISl6f3B2A8Iy28eQKEmr9PWMyejvwigaXZ3wT8onqXKcMk5H2r2
ix/9QomHBEhRN+KolV+sx40gOtC61h/v1LpSzFg8QMpeDgqGqbCl/1CF4ieowOuP
Hw/ng0glC5HsPoptkSS6cfejugHgztSErxTenIfPosApdfpxor9x45QAheqiE27m
bJZHCZUeV+/yATfwocUEXV8DXEWFwp6nSY8VIVWWfrrYQWumMnobHmd93L9TXex4
4COIE+BAcggN2JhSIpKMXcnCYgfcNxJINU04unxFLcEv+v7uyI0vwPPESiIM0nCs
iMYnkGDwmdYuMIQJVt3SdRZp/E9JmEv2B+7xo6ew7NhK6Bnfl9ThfPAAzuJ1XOwR
xSv7ZDTgcppOvdyWcyOwuORRPi7NO/CkOG7SFqlPlTAnvsib8m2ye2RPKbjZScc9
1KUH79QcKm5mU+NJvez7vkGepzxYZXFyfoZzxfBtUfx/WtwEspHzEVYCeLLnMP8x
A6MQ+WWLTjj++vP7q4BeHLSq44+dVAsHuUL0ED/Qpm8Ro5PMLvPIPtpYFe+Bo9Gq
zn6xFL5GCCitXqGZtJzgQRaDiKrUD7nrXjL9PsbHzJtveNBGpchDSa7c3iUGtRHo
Dhcx6TmzIim8GaaNxeQLWiY+DfhkR0Ul8+q3wMjZe6PYCIpOzv/r6/37186Rrq6U
Y5zXtQzCBA94pYTUZW+A2HIrOGgzL3dabdZLiVfp7RM4TOP8gU7xLsgL7ocvmmVl
dFB8LWKJwxTQTTlAgPy4zKoBusdwW9Gl68v3v4BDvtLEL7cL3lYWpSknHri06LeX
av7DQzzewtukVCpohZsw+CgyvA4KD84xMfQ0ZVmrWqfgep1vOgMWAfeAA+Xi+xZi
KZngYsUWoxEAX25L6j4f3DWI147UgL+9yhkIbyTSpMGrrkg0lVKRWw5t62OxBQs+
/3uQG04Z8CqaBPNLCPH+vsWx2VXR7rw2OvhXIWj8x6jarGCLgmqmqbSqUJinVbKH
+8l9GVpryV+l0VJpFAbgxiUCJgq5tSuhYltGjtLbAeFXmaG4Q2wPzjmAryQuOjrA
Q3i5nRwn20XnlhOnO2e11llRFp/cZZiiEaLqidTyAFAIyIoArHuuF/C4TSF5lulN
kuS6vahlq+fyqmKIeMH5U8phRu+n+QTO5hHX8zGQ47o4QvN1zLObuGr8t8Y4cYQa
vPiuqwzO2dcJspkI6j7OE/nCI5dGjvJdM2MYu46wGY9W0YLWupZ/hB7pmqrfmYX8
nHJ6ghNFXdTlnhMxl/FVl4wYQDQGYbIbNgpU+PBRQdlLiYvaBfEi8lBjEZ3jiG15
dTjyD4p5pIIfcTv2dcErs1MvTTkjwNgYNDHSdNOOQNEsJ5bVtnmrcmEX8DtBRVfV
8xgyXBpaPvqwKxjQHAtvFDlsHoDPWSfvWKZ71if0FGhOamyqIBa3XtJjPAsA0IiH
JxQca0xV/TsnfqKLsIwZuiu8i15nVMnsVDGgtBU/KDdc+o0E2bHlVcVnpGR/2Ln9
htRBRApKiXlJZHg5fc8MBB0j3CLdi3F7AfFTiA4XWT4S+spyCdJChUIG8R4p+/Z1
+D1iqn3Qtbm7rk4Fmm39sFPTHL+aTS9EnrCwqqV27pLUBDm/VoJD93Z7tiY2L1fl
qOLagh8IEohxq0WtFlFg3jCN53DebPP+3J2ZO2GD2F8OfoLoOlsYzcFeEz9A5SGz
lNVIhi4K+T49MWk7XIYTwyQkyWaxoe8Y8+PlNQqb7XsRtTx7meiNDMuJ7lAlaloV
Kt/acraouRd1NcLuE1AMWieSg8JlxPenpQKj2VAXpKFJ3526Y/b4RkxBmAYN75n/
TYya/VR6A0RUDygz0h005UmLyfcVFoNptXBtuKHgil8qKkR657EBa7Iq5mgXBjmS
yzoDTvHWv/oFbzqgDlwtl/qWJa2gv9/KctkkEB1hLwJV8yEYZ4AXmqZg4BpykeZ7
IV7L+I2ZRODWTXbuwyp32M1M+Gis6Lq4fEqmRMOdCeMtJ66Icq94Q+pF8JaGEhJk
/EN/mtc43px5EfTGfU+pHMhdeCcITgZvSyC4N3ca4ntgkFGbj6QZHLMHbgZSAJk8
JGE0l0BXikk33vELLtMIrbJMq8BVLj75+BQMCfmSw54a5vMAFKkdvfVtx12boZru
+qSwfYSyCzn6yTkgJ2xCRonWRlbSsbo67wcflzX1Uaz22LRY7cGbTYIlawkvZzho
gvq28oje5B9i3xEzZWzbVF2MSMa8jfkuv7nU69I4qMVRfxN5awvfrGVqYHmjR0No
3yuJ1XPdjtGot5FNeovp/QWgsLdZr49u9L5zKzaasDIECZeiQbTQ8NLsYphwqCm5
vw6gdUDs97fM4MZJdLUrF2zczhelynDgrXgjKL7bM4qUJemRxhzFA/GDfraQkE2b
A0e5Wk6XwvOHlo15vrABo/D4K9fLhUZmYG1XtzIjb7fjssDz3BI31SbcCOELxf5W
nAVbqv1TV5PBGcZoZgLV0+a9h61IUukE8tpCH4hv+6u4ypIFZcHkEnaUZJ8CwT+k
UshuJPHgEf3Xn3FdyO2u2SzUM2xFP1/KzvA8Svfot2xwZIV9vKNOZKFi1B47Enkd
2p4McuvaNvMvD0nFw9FRv/RYaVyb+NcAP5go76RLQHvxVHlmOQpo4me/SkQIUMnO
XpbiWjdAVW9xe1nfstd0EE8xJlwYhj8sE8STMduPw2xyt6s3BF+xriIOwUiS4IHE
veoQOr153/IIwrFpN3iEVPLKdjpnSMCOsw+V/HJISFsxF4P5uLpGCzXpNJP2SV0O
W6/u7l9jL6rVbKRMKnA8l4XXqzIvN3eJ0ly6WIOn14wgJLpO1Sd4tYYD36tdgYI9
c1xx68R76uzwgXhFTldGxAD13/GWDSdYGNDJvok1NS1PCHGjaq658mz0ovqqQDZh
SZ/HsaeOQXntvjkAg/7CGUD4fERUtrj1kshe0Bho9d2qZ46qcWPH3WqrxWtODDKC
vxXcY588QoJaS+jmgqYSnx//7vXIWnNaez6wi7+8DUYf147UklPUzRncPic5EFGF
rVdmp35mpQGnbJqILDyGwKva34puqmu/zt5FlPxsGBRkeayQrRn4xtf/0g5ns4Fx
NZEYkcZUZfymAaL2vOIOV4VNTHMWYKFBKnwguE172d3etYn3zb0AnZFfedRaTiwG
n88XCEnNX7C75uy9h9iIdE28f1WpF67o4WvQIQ7vcP8GcmLj/ulMIb5IYW2ObqTd
6IURo0f0qmTmPLYAGwpEfBN5hGS0H9i8H4wADiId7x5PlmgGHlLR+4zD+z60Pil2
pePjqO0XtwfMYNe6fwRM1nDepv3N4hFmK/xOq5bPHdtlnegbtRk0mCih6/EO/+Lx
qcnKKL+/YBE3GLxb0bKdYRs34HstSN3KpeBcAzOkDlY6n+4IOSlmUHuBf2Hdc9bW
DOiudE9QN03CdWHZQocC+u3GnQw2ed0AwnYjoOBYAzdvsURhvTq2bAn8ZFMtFq8M
E3LxQBuE/N898TFhLI8UzzSAW7/+9bWoCwyz3N85Y0bz6fRtJfNcmlcdWmmBJ01i
Nj9wW7CHZpsgANKAXbhuaLfOW5CZlTLZZjyZyNfIt4Q3xTADPc1lDTAxe1MNWPOv
U34Ss05yBJplPwkb74KPrMBDm4/609F04sClemPwdq3NR+QzdlkYBtUp8dnPheHY
yG5BP537d39I90oH8M1ngIXmM0bAQlOSxTHDllQJDOQCTgaTWY7NMsr2OjR/gi1K
yMPyKqR7wovF0lZx4OrANFy/JUtXh7EXuNMk2YpNWcoFVlpnas2w2jot3xlmFPaD
BIXvzkwwULhQz1DkCfSNmk/e5+eFp16aWcLA4OdpMvdncFKVxFCuIUU9avy4nNa8
JbyYRrRBVSnz33P+n1VVbG72HY3d0u3qG9kGsna1zAAemRJQi3AijrjCQwMB29+c
o+w6Rp6asaHJa62krYYUTTiD6GAtLKzXDxVe7wo5uZ2e707iDDB2pAzm+gcGYZUO
KXVATp0Lh68eUpIyJbfa+9gHhqzSGpI/p4R6HRXYtH4xVxs0pGB5UOvU3sb8aXPF
yjPpL1y3rNI+S0dakZIacUBid8t5jnaEggcWFF2oMPifokfyAMoGr9J1kbpnmGFh
dZO5Zb97Byk4O64rCtU3jrtVJGqMfMPRJ4VWIni8fB4ZYwTjlDMVpCHrRonrO2Z+
ukgLynMzOTK7264Sto+f6J9aVmoHuLFT5UoSiyHp+XzM0hHGyyhs2GyaZO/p2c7l
7c7z9FwDFeSa9Yv4sK7h7b6QmFXYKPfpm6mxGsZB1qc5SRhvOlNkZu0uY63I7Ni3
oKW3svY3seKxlrW84cG88UW1bCiVqyFfa76LsfXQDpWuZwPraRw2Na2s5/1V6exG
PbShJKFAWimVqhH/MLr/J6p/Vh8bnVi6Bi+JEREvebuZq3LAb3zZZQTtNMUfRrSU
dbcZK9gBgVys9IDFW3Cuuughmy3fX2eCqpzusWBPD5edUxEmC1StOmQ7lrkgMTzZ
6zb6NdNWo0IQRXSGnGXS+QCuRdoAVL4psJEqGy0Y++sjDqtL6R1iD04QIiySPzQt
YQC1F075YcrIRX/9i64tPweKQbBvmuckmvpLpfhIRPgdY/aw5nk92L1pvsDCUFcH
3o9U9hBgPxW73/485b5ww5hAhjNURoUDcuwiFseOtqnCT58zSlpbBIK43akmL2Da
tvYSel3Koa7kN9k9jejxUF+1S25Om0NF5fmuTY0pQcyj7lGQDIH5+ZfwbsyAcOhi
4MgY+XfqHfDNrFr9a9EOKs8/nIl6JmWbT0h31B8l2VT9/kpWOSFUD7R90TeVN2zX
bElZA1iGhH2/zdkaktX280pEDWuDr9McRJBpafaoSeaiZkUqonXLnGM28a66yeJV
lOfX5ApsLR7C7LjQt6T7voAhyfJhPFxpvPUwMqyz5c9ADYuFdQNkptIU11IGT8PD
SHtpckhyKy5WvtDlmyiRbKHk8kTmlX54g0WiowsDeGFNYqxAGAgJNBrl/N6P28QO
ahZz53iwjSqW9eM6hPZob6TAumJCJ3tdNJNThkN/jrOkP6dK10jhDJiDoc6d4/Bs
i8dPPUSVRpSk84NoqBmdNsmK84xRZBsprOUqjgQ2InB5AfqB1b8wXqyTfPhcaIem
MLLdgYiqNZWYSt7vuNEwQXgOgG91oZsaGDWZyrS6DGEb6E1TYfGSm6+qwrIccfqF
kSo4APrEohT1X4RDWRAMKZHTHMNWqeFTXaBLUGzSDCSUht2n7NPyN5xQv5d2ZfUl
xtChtJS2t5JPpEmsZ30f/76Im3znHAwTGRgrKTw928weCjpLHQxyTf+Ne3aOuHmF
l/OyDNBunrW4nNeWhoOFkPovliMHZGbLdf8SUuwXlSHd6X77mbADUpaDAU3Ale5y
8XC/7TXTY0p5ftWVfYo0zdXbAo7cFzLmQsWHeSyVmni7a1khaun3Sim+FS7u2UTj
fYWao0TmCK9QVnXTf6gWapxFx91elp03z7N+5PK0gyoRukHpW41KLpVDCtZv1xaT
E+Rt7NcHOsGrybS0PZvhkWQoaKY2u+4s/RfaoKPNK7df1HQfUEoRBPDoI4n13VGo
BPXG0qhQCUm38Rj5psZuwxeUlEhiHlvzNzeCqeomq0/hNShOhmN4fuw0DcjpuDSG
4eDxHcpwsdBQZTSy5zya2vp8h5l4IHgTbtlk9zU4qzBXts9Z2euNgZjW3LdRpsy2
cmqmNfyHrBRxw83SCldkPX76l0F+NGbD7yVA7e2wfZV/WPV++sct20Y8cnp7c3YA
O1qXOY2FgTxGFEo3PizzQPqXSMhlBWomx60tAp/riwNgt12xYECBJEcyc4Sr19md
HdiSpDU72OtQaQ1p7x8hgSe9h69J8M6RonGWL6TicyOR7/xaE7D69XnNgYa+Of3/
uMZC82W+vFeJ1CwfcpLeKBW2tOafyPX7K4pZyog2UoQnyMs25M7W/Nha5ThF5DRE
nWVdx3vG+kWnsJFjfz0i7++ZHvfeLzlZVrFt7pPoQQpPQBQ/5jaJ9KNYYyKDk+Cr
QTZOP3pExR3Df3v9hXh0bjniaOQhvTt2SRe5uxVQ4tYFUVQOyOOw62IX5+/frnvz
Vy7CSqG+DIRNC20GM0vsbeWsoTHbVgp5lysb7M2GpDhNbcNvHT4rEC9sYJoy1Bdw
T4qM9luR5DB8ISc+1Br2H3uV5ZB9HhNXJ6QVisfZj0qUdpP3CgObb/yNxf1gjdz6
XmFuP3tWZaAMrLouYdle1ItK42Xb8/4jnXNENhPFgUuuOGL0MLaevw/8Rg/GO+9+
wQv2a4MjvdYB9Tvk5NK4npT10gWV9FkrogCDkvWNUwNv7HhPfZkkQidK59pR3Efi
aPt0EWOPuIAeA6DIPvtyaB+xoQcHUowBoVgbUdqV2gmsZ9vI4oKoykEiQgcYj9TP
AoSVbC9DjUQfngU1JaziDsdAKxqBtslyV5dhUpKKdk6wCj+7PHJVaAyZ29qQL9S1
UR39qg3gn/ouNZCOQRP1cyWol2NS6T8u6IkKjecwRSGEgVAJsue4LuLqJBBhaEYD
W57WpNf01v1JMGAaRki1+oRiG8pO6Km1Pfk9cRbXHh50ouAIygWiHLaD96i9jXq5
7woYamXPiNa0vf47xd3Coy+xHiSWLYm7QUSM/UZvjWvckVuU63w/vI4SEkjFhjLP
qFASxPiG7FLAMMNjGxeWQ5mYLxG4CzBY88ucOskhQh8Fjv1momxMM3k3ld/UKEM1
qn12PRxw6jqvsxKGya5MbMFA8z/ZS92gvei547fkXKOuKAtZLjavWIwqPKCNtpSv
w1wyugIej4qIFdsof+WfnFLdaaYU+2mzE2n8oHT8i0iUj+RvVY5ncZoTaFlBUxkV
7+EXHSVKa0wuTJj8lNF4zSEWpAxFtJftg68HOcZn6VUHQ6UxOETTU+wGUn+7eGP1
pdHT4yVtJBBHoHUDf1CThDQPfryQEXhacwRzC9HQIbbGyxxbjnRaCdaAT3MJ5S5Y
+DB5sN35QGw6wZgWLaPMMi5fY3kmVBL9rUCy/1f98E5sGJ/H3dwgKfbwYNAjjhMF
qsDlQA4lHmHpoZ0i9/KkJkxXEfzlgc4vUEebkil0fl8wvq+Z8gHbxzatYF+k5/Oa
7oQdGLF6DnbMkjVsRX/O9BY+xfG1Fr3UsSWYcW4KNFnYxG/f9FPpeYRTXUOlcc2X
XDfsk2a+cGyp8+knX+L3gWLUQHSEO+MK6EWQKwIAtCTZL/9M+d2U9QAIZdc8OhTA
4Z6dA3hMzo5JgyrWUwBOJiJbLAKgzt+/aKujsy7L75Ex9pGOFxjOdGhdrfKSZyXR
G/pKs3v28QO2ESzk9BRPoLobVFrhYGmCuymCR16OVZrBcbtyaa9Ktpgwm1DunvTT
8EQalmGuZl8Gj2aV0DsZbWp+Pr+uGN8a4HfVw8/ljcxAv+bFYfWxjdce+VCkCkXl
r+bqmfsLIf8l2JdLn5/iPZa4fLbTfCl/btL5wdxRAWiC+YeBEFfozghqC/e5KjwH
ZFtqGQlC+Flhy6BthDCJrKH26Cm+zK+4BIr0S9AOrLvaIO0mcoy/3Js68ux+PZJE
6gTf3qCRrZssxyHlNEsMlQoEavkD+IXo3Kk69+yuO55ojFZEDlh7ENeY01Hvt8Gy
oBUAMuI8nNVfYlH/1yX1toOuTrxQ+V2riGU8RhGBNHNPTdvnX7VN3n7CfVvydDFe
lb01Tik1xC37FxOv5IQHg9W4P98458ry7qmjoGCVuGncqHeLIDcJu+/8EcUPCw63
cNdZ2gjvgAH05pL5Deb0TGK2enf9bUKB0lrtyXbi5ws=
`pragma protect end_protected
