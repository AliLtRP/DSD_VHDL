// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fEzgAfLdwpnkgJrV/7SoQPtSpKXdYazk0lUJJKkhQuILwW0BtLG5qR8yQLf0TkiA
qkAi2bs8Ry5Z5g5U1HUvLb0Zkmzj5URbZ7nBEJMX+AlrHPiAlOGlUahgNGRhw5C6
jfkzWlKTGFllS8ZlDDFXAsYs5dP2/gYbCwB1hHVqXns=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7424)
Cs0GZ0mS11S18jFfjTmj2B/lgxeaF4j4/vG9q0D5S4CXKEKYXJVLMpZioUik9OcU
p/qD5SLczHmSGIcAVzvdgeukMQxOkNrR3A54Dzei5E8hfhcST42rIJKj3EA7P6ae
l31/Gd4+53S/oV/seiW9Xz7pMLfQNnSyg8LuXgnuIMBBBPYd5V2jkM586qt2wVBP
i9OrfVr7iEIChIYOjLLpszAJ+E2tJ5dA9DFIRkxzvzf1SyQYubghNAIpDK7j6YxE
SpUAL615X4i4qreaAprKzh5E6Ten8VC2+ZHzGHMhi7aXiVFSN6s2njVzNsfBTKUm
zy9p/9dH7Tr86hBrkkoFuQF9avv5A2b9cQcImh4ONdIxEzGwPvG2g1yfxGsCJah0
3f7hxQ/hKNo7RHiLcnzHFB9QaRSnk57ogs/LrREtM5Zle4TrTScJQlN1KYfWph++
cfUQA8y1lC1xFehfrEFQZeAmOIEHvq/HXGglwAYFmCsHazSO9bkzKJHqs08wu/Jg
J7W7uYnv3EuFbsXc0Qh8Tu5wHAtlVO7kOWKve4OT9hc05/YQvU1sAwBzNQZNK7zD
n5iOFxEh6WDWIzf3Ytgt4x6KbggRl0Y6sISfUN4B13Usr3DL3uE2tvnI/sx7/wXe
gpssXX+OP6Vc02x1VcQpuml8jYzPk0LsMZvCTgU3YgHng0k6PW0gd2joEvmKPQxg
5QNkQFoIrJEp/dGbQzRyi2voEEQJN8vCYYNPHB1chFQ/Nf5jr0z29bMSEDyH55h6
KmPZBLRRY6heyYBIxkAod3dXpG4+QrXGyRKijfa72HZZbTzl54B6PxztnCRvzivt
Uoyrw4jm+fhfZZLbGj4UnAKjsTMTT+ywFBkzjN/TvBXaQ6zxaHZFzM9ZOMSaTs7Z
MudgOc2UpqzcXEy/QfGC/cEmRLjTAeRF8ts7tmLD7xJajTD+aDjD56mGWJ4jaqS9
B2CId/K05K+xCKybaYRTPxhQczvq2giRY7O0ie/A6z3iZldhFGsPIt51HoqQMkW3
Rh8a+1VZGRw+BRRXjrRVKJvSXCWAKHlVC6M+8NDTTaLc5rQyF3VO/vuqObsZOkn8
9xpiKe4IPtGCpWje2DsYqlE+zmWWAhtPVyKeWUMyUb0QZGUtbc4CBq/Pvq6Uqo6v
v81CXGBE25jQZ8XZ6Xf1Ma4fD5KsY5bAEIKQibKuqRH/dDDAnCbOkRi+Nc/EYkg6
AgbHy0HNEOT3NxyR0IC7uZgK3wkSzK2A1RyDRKpcdOXScBP3w8K6exhAuo0P7Im9
FiyC++cmi2J+GZXs8LXpkdB6Ccye6wnu4Ys/2ADAQ6kTFOS3ZR4Jj5FPRbAkDo3A
7fC5XlsGGEnU++66FiQBgQaC0RuaO0OG2SQYn86izIBuav8rsKeR0rHK9n6dprcu
vfMx0BaT8OSKFWQaw5+5sWjERtj/CXRKVEILNJskIf2ySctJKvNQE0N2SH+3HN+p
1uSz9WmEnNszNmmB212LgnbSO+EEQU3AVSo9yfW0tiTv8BQEUqBQ40sVVGgJrB6v
LK0qVmAsrPLEUIwSLoU8UjKZj8+Ivy1uDXT1FhIOAmm/PInb96uZ7MIDabIGtOvn
pHo6q8DjpqSLOrPvXRGQgdiRBfvlaEyJGBf3dSHy4Ce9Vyx+mfv1XZUP+i3GZHyB
AiFM+e/dEBx7CMjUZHrmNhvBtsoPORkEePQ/HZuP7m5vtIkCZrkg85uUQ6p4xGQG
lI8IHM7QwdJx+hTBw2xk3vYkU1zw1JlHPvKgOFXK9dx5ED0SSh9Ubsjjp1NoZy7d
ahgYUpP14XtFNzSc+cfYRU9VVI31/TGBZ6clLea+wsUJKOiXJCx+sPvw6TBjJPRE
xk2iUeaW6+DAYgpGmPFhWZiabgLC9NHxI74T0HhVNyxADDbphj4T3pUVDxO5CfUY
TVMAneXBtOiirkyyRMT2GLyhwNZRgsXR1shfkpZqLgb4M+m/jkVrzroaOLcsQziy
IbskSKlPZB6qOvx0JHDrPNPwbkqSj1iV5JIWqhFJcB4vcGy5iKeB+U6mO//Ii3fK
m1ZXdnXLTuYQClX6UTx3uv/fir+FGkUKEtznv3svmsDTI70mQUTCLANC05o+grYM
Pt2XO5eGm8DDt51whFHTY1YDPQOvk7yij73Qa3Nm8a3+V68v7tAceTxPUIYgRT8Y
u2XkQ+/PTuetqec1gBkITYELD1CteGcS+I0gI/iePW7BLB03LdxkLX5L2LZGCrkB
1GL2N7jGkg2qvbTKKte+MrWG9qkcPL0OKGHeghX21C07kbS7xxABdNn2Hfd9T6XQ
PG12cjv5AyUHnqbEAUy51L6KVNXnRSxFroALlbjdcalG/zfz5f3MxRJiSu+2iX7n
vwjP3SHV50tZ6K0recIJ8c5g4Cfy88ifmdLtigOBswjYosXoGgZo7Iy+Dr4v4ein
JwXPbo/gN/6ZHoT49Gam569EdcKrSKqrorzfv3+7DCqpiFaKtXKvkyXIyGSbhVZv
0rdwL3XhKlMK1RLrL6dr5jJZ1l8E/kOV1M9Lic1bv76iEMNsq1BECygK5ioatbY6
UpIDuzfNdC8P1Iql7bY/vDVck7Y4P9L+O/E2CMwye1Zard3d7vFfD9miz1MxFVC3
7bamJ0IEXaDF1uPKABUM9J3pQ8Us4prkIT/cuP4cquoAZdUsdYzcTTXDZQuOoan3
Yt+GG5BFJpa/292mEcVSHCL5T5xNCfUe/+kfpLRPgCGRFy3MCMNYMKd72mAKYlVZ
4dvNK1TFajiIn6rkgFkUWL/uNXWVvx9MJXU7PnKkCW/HmDiAfLWyqJRQC6CR2VVd
W8chfNHtMYC9pGDw8gSN03DyWTFvypxRo5VUXi3yTDSItIobxBeMha+/qj4tH2Vp
qCHH2G3gF/gaCzWSZnM0aXmS3BXSo5PjiZt0PqrjFXVoWQMxoEGvtEYucIUUXGkv
lR3vkYnYcJ2xHCBJoLyonw9X84d2gYEZkcApJaKuss0hqtZmCJsJK83FjpO0PIB7
fSnt+2LbQ+8I+ep6fP+V3zhtQuIbwCxPYHyx+qt+bRxXuxPU0//6YpqKpgHsC8Fr
BEPMkk9a7zfovXG84LIuJC+j77LgQxVInG0CYZcal1uh1rw8bgtsK7O/KLOn2sTM
Ku/NKnUUEqjzAR5DBUSI4RvKmBAg8PsEQyNKRh4OIu196kf2gNK8PaZkoHreq5np
O7C/GPt5m9VDHI4R/zCTQeCI0tDMJhSBdApZAqG1bQvmF4E1qEko/ZwDNWwOfU5g
XAVMRb3cJujxrXM9W5Qj22cSg/J2DFDCPKNAtHtD6yQ1CiBByMfnL/SKA7WTGRGN
+7cdPp2rVixlMfK9zZI77ngVezVo6ou5IMA2ANSwt0KyLC4a/fVREcCNfYlp3Z5h
HStheVLoeecb3K7gLJFngX9NAdZLsxsNP50YfuowxEI7ADwLVSJYD/PHHlNJKxLK
Zre9wYpOink5fisjVv7FUxIz4Q6RXgkg0Y8MOu4aYd85YQQlcvVHR+nqDGqMc1ye
wSUGl2jRSzm44CSQwNRN1rj/bnne2bdxu/ytd1vjiWil1JnkVa3dJXAr9UElQRk4
uzFQx0SOszd3AlGOxblZY0nA6/KP5k5nMOA2nlfwVIA8UlcvgXB89fi2S/4Luqxs
opJxgMRhd3bNpRJVieh8VYJYH39rCXVp/V+/JEULgqtogUoII88ify6K0paXEd9n
kJP/WFL2s2qitDnSDiRSBnEE/HVOrKNoltGoNQwAak6p3X6OnptTwlciUgMKZkOp
5OXUvQ+WuKLAE4ANdyhBrGNAbbtUVk5cINmehpjCqOZqFcdYqGT/bBcOEMcaR+76
nrM/d0XcBcZR4poZiezhd5GKoflCowp+044tz5OX/VkyL1HtXn/QPOoG+Es72jkW
f7ppdsxrPCyylCsau2gRQYras5yxn6Z6frZwl/VipsdmQWWJJ5iKJmMfheV8jB+g
ZuW74XfNB1EfAj/L7b5iSu8ArRCKmQ3dyARVBEWZHZ+eA4ft2q8xzv1M3chHBzuh
by6X8pcBwI/0OfEsRMxWV6EY2ozVSM7YUPWd2hAl30KYkvvaMT2HhfCNoXZcfANI
XsEltefl9H3buJiSF8EyeFW9+lA0Heg59ce3JtrwWLtkTpAT8oRUazHBBJCvVbHE
iVf3hTNRy48v9mF3fug8KrJIYu4Vn/E+MMXbs2d4/ozUKXcJ3DtdEnYKEon+AEY6
iWTc7i4s8ROqKIl8FHyyJnil0sftHJz1eNLkYLH1pxr9hKaxjCFkCTFidXpoxkK/
gvZX3OI93Mjwhwqaso+bJzTesSzzP+QChbhvaceGuRxmYKAdE6FY50oAVUJatyRp
SWoJf2s7vqKprsjRlxf9JSm7J5teMiX8uYerq0PmVtvqrfyeIT4HUP6YqPAF34fe
0Ph50TXtQvcr7Yuk2iLJRch39CuNPq+vt2t7aQq8z/xSj/FAaGbL3thSN/r0/AyL
tOgNPGuriCOQXfrNozYqRWWM1CeUAMmT/1j6rDgkWewMAqw5tIUyrL7ZarrJyqRe
IeHEtSafXlokAAyuX6bzK4CG9UUhKR/LXpqnhZMQsC+lYeEfKEMj2Bu77Ye4MVpa
uOTFyVoRI+2+82ABFO4VfmPmlsCKJDGX1logh1zIMpoEvA2h7zKxdcpJZqMX5Rmx
q1+kv9jTysfvXyDdq4i7a4nkvfBFH5Lu8ejc+H/wwu1gkPlnDh7qD9f2xXx/nvwG
TyP80Y5NH7ZyI77cStZtb7nWpWvVA5wQmUMZaoS9z8jRSioiouxLVwdvbikFDhk6
urV3UctGlcs8xRvq2jIeUriDV0JHKO/69Ukm0QOBLeo/bjbnVKIC6i8i4BHOHiwt
AoKHZbUfJLG7MGiznpR70D3QZziq6YB05tiIxlmlDSg7LV9RaLgXTceEY6NbvmNa
6zEmWZUZ6IW2tvY8vZfaPtbLtOHdnuiJQ4Cw8rvcLfPbKP2tA68L+Uw4lerCl+5y
gJlr7q8+CKEK3TtW2myMWkrhecoR7yc9TPQnK4gD+WifJmQQYQZKikoo+J/jnFlq
m+xhdwEFipPDc3KW5WTtNBlBFP9TaOLoSmu7vWiltt8i7sTVXCmisLyQhB0q0yge
sScGqlDUxdF6UZYFKIUyxNWZVOSTEX6Y7rEDVG4E/Ofwu8MMu9BZB6kldmYOUes3
216wzdcw2El/KeriInGhtme8iOHq7V+FhcGgtmgW/9qHxXokRYzkaypxSlD+Q1RV
Np7nZj0flh4kWLkCNVHd7DdxkHZpkKE+LH7U+5fMJJbZ7tT7ZX3N0UbIyFTwqfX2
aGNbhjUJaS7e73r3IzZKngkdLMqzr1OdgiEIA3vSzLykqvC4HB+/pE2gMvKXZlgO
d1ZdxIPhmNtfwGqiJvS3QvJ1hg6lekgw2SfgC+Op5dcSqXgzZrtNiTW9EthJjrQg
dUO26h90BdcXA9pquBZzdHx1YDQCHGOmgpvNuGQQ0HaRf+ZtHKenpv6Gtoys6uDI
HlzL6hSRTevzT7yZjbFiz0L1itozbknjRUT5EhUqELR/kFDIBXEpSW7mWuq2zGYD
2hcidGvrHfQDmZmVHd4cOacPAaj/UbWO2s1CElPBWd0HcwPE+GbAvoJ7Ftb0uP6H
1hd4IO25t/IR0pnOOcmqR63Fx3+CA6fOBFEefRxREyhTGTtChDSe9UcPGu7KwXI6
e7PpVrI65R7fb4HXuFZE+PydJ790tG9XwD1Y1EgF+3ReRoE4ZS3sbe/BQ/GOzuWB
kzPqkH6Qu//hfzYNO6Q3Gkr5N3aEQXa8C8dQ8E1h2Brkowil7Hk4RWYE2Mej/fP9
OsnsEEV3EK7DDC/jDALf5KoJ7oTqcuu3vJYJEy7hgD0PbYHzljYXA5U4CUrCjwzv
aUpwUxSTVnJob25pXV9zn8WkcskO9JamuUW/C2nzLjWVJcruU2B8enwJVUuAcQtB
KdfrjZrEUXPPrnKKYRlFQ+b5Y1q+ns+18ZOk7xgxWuxS2AftApCyBWXVLrY4fAYV
tzDKlDn/rheYyMOElpx+JiUu8ZJb6Q/vpcVCweXbLTL7JSURd0i26k9HxCHo5rJQ
mQ/vhm2f0WFDe7llErAZrNlrwG5ATicT06Go8PSi/xa0RRl4RfFPNN35NLgomUg4
nnQEL0zwgPcJ2sOzazKEfSaIHGplgSWLu+6NLm+SPaxioF4AYfMZH2raZ20Y07vd
Hxx26bIwW854sYTuDV7JUs+5Jhz0Ir1jLzCqAs6Pv+yP0G1gsfYiqGE+3kjDh/Tu
DMh+qfAnV1GTOaCVEba2/G1CnfCc69RCImAldBi8sXKafaZ/DsrVCi0j90Sn/LTV
As2R6ViPu31UfLGPuNaARf0B3QXWoq8cPC54qLShmQfcmKqjzqu4ov2omCETOoHi
zU4gZ4iIXfJ631dAYL73NM/eBFRJWglWrTTfZJBhO7n+AnmIH5AJggHSb6Kz7lW6
gsDgCstAD1MaVGE4kFB3a+QtQkYX5gIQNKQJDN1jpwX6hy+5fU9KL9xRR08PQPYU
QIZ2l9PMvRmbcobmdJgDjv0QHxjTI2szIyvSTi/bA6lTxvyxsp+GBL9SuoCXCk1D
0PFh2TU+5UZ8BhSeg0v6BXeVONl/5yzYmBJk2GJdU6v844/QLWgGAY2lkcavm0Ad
q7DKP1EmWQudsz1RagLCOYhByHOElzKi5bcqILcrN14tIeYMKYTwlkYcr+ET0irV
f6z/UvnhlvDyz+y2E3+dbzKjJC0cOA8FWZj62SLcuN6FmqPEv95xGkTLJtKciFAb
Ohl89RSu+8dEZbjWxclbKnyC5Aw+Jd5x3D0yvcG9xeHUIxSzAhFa/YEcYbHB2DhH
2Xh8+IM2GDzVXnboDBlPB08zoenr8TuhyivKI8ZrJBP+QwuJnc3e/g6wD/qFt4LN
YAPM5DVpaYsH5BvPGGKd9MxenM/t/olhviHiv8MAbdqZwfky6DZ2xZyLWLQ6IKNx
QIjtTrlAXb7EhReKxqZCun0Ua8xRJ/UF0/T1fF9gAc2T3JREHeQF4DSFotJL0O/P
mkSjPnSxMHErS5RW2p6GQbRhHmpLYfH/Lps2KsMf1k3OO8MePexBnRbCm5YXOCub
a7HkBgoSbvuFsK9tHZw8QFf+HKRnUo/gbnj//OCYF7v6Y1VsphJ4RM/jpeQyOU4d
QEJG+6YivMHMuUbBSSrNaghk7yOIspjYeqCQKso39lSgCK3nsWe5MpLzknRatT6z
q5K+xADUfGcV0G3NZ8AvaOl6t6rgvtt7PX45CejO5kRiwiu2IgOpRzWjCzcbvhVs
yyev82oEqGVwxd0rO+gsftzyAMxGEN9fVH2sdlY7cpI79nNsggQOs9ql6juy7nZb
a9vS2wUl7Q/SIu8fIJjIGX9ainOKBUopzQNG2BbujdNH6gkQGe9J3+8T8Wrbm434
G18dSIuxIEqj+6IBtfU9obSGmbXI603cM1zEQ/KfHUbaemsOP5PU4pWIKar6fBir
3s4wu/VKZ3vemjKjx/jpa3gFAACGjFvyIPrcllb7R1RnGC4F+1vS2ooGy7NzUI5X
2geVgJJEZZbJMQtIV/wtnXQiBLu3biDI78XiLJ7X2/CeVTu7/etvlVjhNbwY5WSv
PApJqUVCW5x91nTDmVwRW98uLDIFQ1tLh0MQfqxUHz7r1QoSHRMi8UsWjLhxdtnk
bAxPdQoxV+9bTMj+qc12gaW9+RmcEuZRMkMZgD33AizM+759KezdBxSPxVP+ka6g
A4203JKf7WUZLzylrbKwU+bhNsMqDVf21LF/kglKLpM50N8zoaK5Uw6KCEcixdAw
ldBlb5RMUjKPgDwVOQ5xQslVM7jxEkbHn4gpcZuCAHG228DdNeiQ7R3gwyXxHNFN
B3C+QjZCQNiRftAAVYUCFSWAd1tZmXzKLbvKMj/fOAe4BgSVyJ1DcNX/XnUyuGDt
nZIf3jMP93DZo9sJJm0pydYex2ud2z0ZwtGUuhaFna7v8L75dl6dgyPR7SyGCBCR
u5sCmhoemVMW8HCq0UgsgDGJYhbrxIzYEPE0Rd0M5SvDug4WJk0vKU8QFga1Sjam
e/IL8cj6B2oDLsvla654iDdEBR81MU2KiXa76U6H7QQ0uU86Tz5G1L7W3wSI+V+U
cDloeOiWYBU/hC9Tt26hgmiy8TB3KCEH2KeJiUT8M/HFjR2eCvIErrNkWqOyuWrs
WjFiF1COfYZWH4o3X8+kFkviipxkc8hwBCvfVoDwQJwYvMc72ygVOZoo2kt4NEVF
vkjPu3i+tjURgqiWnoatDJaYGEsqiKAL8vHeFDe0PyT4AWijok8qHH39+WVTV4X9
Nh6B0rTW2Vq1j5EdivO5gyycYFIXjXe5Bjby/pD3I2iGBzcmkoZ8nv/3QAYPfSvb
LYlHOlHuj/e9qwXJOhNsJNK4enJgbkIJXQL+Yu6Ezonow1jvpQfXfCmvrNb9pFDj
wHAVs2pk7qBPdmPpEclh2JP85nsr/9k6C8vMu7exS7mf1bBHleUqRu66b2DxrLVK
9pOabSwgr9d6zcVHmA9pVJ749jM02vEKtI+2n7b6dOzuQ5TeZz//M1q3eUy62Khs
MVKg5/Mc4zGg8z/d48uG/pDxVvoM8kee00ZpmuoniiSiWEUvWYtLJbnK6Q0zeWPo
TACXbS6oreEi1JoXjcXf9fIFS7xqwRH740WPjBo7HqAfmMIQ67YOsziKC4CU5sT9
j2RQYMon5AIFE5HTJLyZk6hz/J+LF9pK6y6uoGiu1+DKRe7s+geUTNVGCG1/heM0
fGAFxedqc7WXArjIFSi9x18m6QEh9B6wURj9CQ8oMEeq0/9tW+dtsSF5xstanA7j
6o9zhCZk0qtU7N/gVy+I8ggjWfd6b5+J+VRYEwKh5527cAMePzKn7A5Uj6lAs0AQ
w+XVD+3CICzW/vE4DXWr9A2+66xG/XcTkfCjpciQtYHg02vpJTF7i5yjr9IVifjx
d3BPtfLKGVVKSDe4Ma9DqPUmYYW9d863fcT+VPovAQ1WD7H/KJAuYYFBi+B7YePZ
vH4Sy1pQyjdx0o4jOv8NkGwKTh2CbSsvHbvmyC62BWCCCg+InvvjdSDkKL6Ji6Xq
vRxzT/xPlWHlpWNkSG/2I+PAyfiT/M8n8wkKtXFuQHLRQ3X+En7WP6UDZU405Ngs
zf111KKE9/7mZNMcKWatEYcPR8vYMF+aB8znHvYmXT5fV9fS3OxPdXs+DOU4KgAn
43pczxnGAN680VUYX/Zpk3jXzeiFnhOabTgYheAfV87khKwd2W8six1QZIKf0CvX
xBwx3u1QB+09SQKVHQxxWvByrBjF+HCrN6seo44Vpr8OU2HDt/J6VIwY5j/963qj
JJbblkFYoUgXGiv25aZOI84Np7vey9WShVHkjHXymDDsDlk176/XBTtgewGwnrcM
CGMwv2vrLxP9rvTluhN0h4ltdWvqPnNW9KDezmjr3lvCcZ0qhf1VF/oe0zoYkY2w
QACrqEmlhrIHBzgdFL8m+pkMf/JLt22zZO0Yxf1VO2Ky+/NndNjJFGjtr84vZ6pv
PjldZqVKn9cHEWYV0mSv9EUdYKVplitNiWCH8vAGt7khkqo4RwSl3wxNYsI4W/Um
xDWSrmYldz4F/+aWhT4umannxVEptdxGMcS2V2p1Uh1ugo7O/2Pffo2yvjyoRbn3
pvFBnN+KkgGZlR6WvJLB4fJn2sF+xnvA+Q4mkWKcCFdOnUulpv5dHmsjIbGnKqLL
kXJ+GPEtQxxB5p6VfMJr7TNjgUDD4elzDp08ka5RXHuiXZlJCJcm7VNefP2bA328
Tpfw5568KldzQYNxaSaSx6ro09H/dZzeXBfrq6pGWTM1rnB2C5J2dasQ7Bruaryx
8iM5uBiRvAKEVGgdC98qcSRmGVtK6/X+fYXaVXDc+2g=
`pragma protect end_protected
