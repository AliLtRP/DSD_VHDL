// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RdjMTCEXT9EYBY0vkqpeWHPhZp7HhhSJVseM2BGTg70s1ZcSIj14+lsJ1WaMctHS
Fkw5JHgCAJxGe8+MTgPk5QTHSLcywSwHJHnHiSW4Ue/tP2bkFfRJko0XYzB1p1XU
zFS+s2atC5Ibh8cMAAIqxMgljW6CtAZsqiZEca2u+40=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9040)
WubRjKj4XPmZ7jZ0NphhcIq3bZXJ7w2n/KvceTgzGmLt0dlLMmOrb7lyraCXiscd
QP/Jhe5sqArWLLiebJda3ji1nj1dRY+N1E93sS+OomrN0O8yhtqBYo+0ihQiIXMs
XTzJ6AV3yfHAnspf+OfmYnlYXZ9ndGlMqIkGShaflU6CDNDl6m3HKaYWKkK9rJFj
AYX6inIDsFUvT6CoXxxamkp0hkXvPAGWUhQRQtUyBcKYW/ECrnktK8YkJPi5sTeT
FbBfHSHV8ZlOPDZyBZSt349vtDSEDiQe800HNRQPilcgAH3wuSkhUKXXAnWZ3u/9
p6KJu2CT7MfzBy2QxhmoAeK71XN5tspUChUn/7I64HuRqzbQcxXv/c+OwyaA317o
T6x3Seq81+iouPLAlPHFlzzB9xVF8W2Tf79AfAfgp/kg03jsxYNPrn/0LAbKvKIx
aco+5KNNMdzlolxtOuPiJJ1TWJrAlrMMQg7Yp5pFlY+d51hW2KXe30YK9hWzK1PX
P7MovtRAnnkmWn3w6ldBWgj0KEprPrLMXdwhQmHmi1zcTGWPPWnbhaX5nSIrhg4L
Y+qbVQkCgSp0RoIn2SIBIZNTUOn4rLTPLauip7GR7WafHZqyMibvvNEeMWHVhXWf
l+wosO1Im7a/PGNa/4+OvRALUhScung9i41L3rzECmd8RRFZNZMtx88d7eFIIT3I
QCamJ+N8NZ//U+zYBmu/3oyQVhVpI7wgUX2hDJXIDMd0PgcL+DplfOKJRtqYHaIY
yhUGyXH0xxF9goYc41dEW5S7THsGEgGD/sTcb6T2vJUbxJ6S5FEQ9cEQHpqsR4m/
aymJVKN4iBlyBwuPgv/EuHlV3lnfmMprvG9fDcrqTbm3GkO4A6Z2jOwtARopnBHg
qCzKGmyPsPbjODUjUT7DSkujGxZP+dT1vnDT52fW6UgIIf7FCvqWp+oltioJQDXy
9gokKGgmtepgPMybQ6CkLo9i6dy5h4SdBq6xy1YtT1dOyY77lw88tL0e0Fg0RgqL
YUDnths8h8nvHIBZZH5Q/zL2dXMD8Z5JBl5LPXIWL84oC9P8o6vsOP7T6wmHaOx6
wiEsb9k7/77k6OTAnh/vLmIzs203ecQaYYBqRF6R5H1o2a4Ai9izbyjpcfdLc02k
6AQA+W7B71iDD8uFu4SPMt0dn4emgPGed0w7KgHIzgfRgA65OzJKI4qU0u1jdQ7z
PsaqbXscnxTTH3CW44QgU+Tj4ngYcmSxp/nBhhuIjhTbwpQYd6iqt6btK/OYsiuV
dm886TLVns62othOi4mZzncqLVRINJ8+CEZg1woCHJw0vJC0zPmyzMszTkLncaEF
qaDeQbI77xcctrQlU+8fuvRJLDXXQL4RCOqnUeOCr5iDn1QWucywLR1alvZ/TXAQ
hNaW3Hj7PEOMAmx1gGs8V0W023gPc1lL/h0SZkEMWSEdqrrs8osC/yigeSqHHw3o
jREV7z7SA83hnkCTU60/+rlreJvTcFUMEQwNa9JnE/somCu6xPFU8qCktIZeSF+x
OIJRFG6+3d+8rO5mggffWFu5b/G31k92LJYUy0JYL4STXuDmlHolzuNgU4TfnhGX
inDOQyWY+Ld2fd0TSOEeQtI6hWOCkjCqebu5/rE25H8jQcPrMTl9I4lsyzGP2Faq
cd3AiW16o35fjWNunit4U64iOfek4/Z3XYaPjV3UOSVnwyXVtiMutBE+l5lH1XRo
laxidJqAyxj0hnLLFmfPOG7KV03PdmOr+fqAeZ3Nh3JnBGRzHQkLMeNyDuR7hgwb
wKxR1NzpcX1Ih5LvChrpNFnn94snGIA4NUSihrJpHop4QFLQ+IzlZp5kQJLzSTEz
ANpmWGCuiKZSQYkJXVDRJpKTSyS+mXNYYeONWdwepvQXANir0y1z+zXm8qgA3x/T
oaBEqYhagM+ZGU8yq4fJLihXwuVzAGWwcoLRG48hy3Zi+TffF/jv+xcwvHjC7PfQ
JyCr5MNoVeTYLbgGPFRcPosaQFOcBSGm5ta2cryVKrKzi67/It/WaRHl+/zgYigs
ADhBA/c1HaVbWtFGTe2k94RGOYTxL6H1spkXgumAcE/oe137zrulQ6/0SXaHLXAS
3ZZKQ89QSFIpTDPmNk7Xu42njJRHk3e2mvQenBgkoUfqiO7YEeAozyUdm4D9E6KX
YYkzobS5gpnLoxtQ3DdldMxQv1OdZE4Sz1V6fZoGXSvgdIf/7ohfOyUBY9c1DzMq
HV+FpyVnzR0e8bCSn4Eql/5MRRQUcRH8SBCZycOmjmxeajsM6ldLbQq31R0YYAG5
jITX+2qnixJdcKPfTsN/rvQ630yqvbpi8QTQUBx3t+wmeP5SAVSzSlsn8I44/QAT
Ab2hB0I1ntiiGqbwj0lKBPNjq3kWxEM3UB2WgX9L9/+ADZLQ6dtmB+HjkqO6/jDD
e8LM9NnZoaEvVbGI2d8Lf/BUGbSUsg7xeuxoYrltiQkjQZ71DpymBEsTpC6zymDj
/hm8DjZfbZYWRpn+vuJMUjw36sscBHNbLbN64o5l6YchINFnjs3QUH5TcxdHdwjO
GQ/m7fvWzTwQjZOY9huhDuclimIN+9oJ31TNQm7BOloiJOqmIIU3UCZTVC7wSON/
PxshauPdxMR8oJg5h1Bwj2D5nmR7l7vqZwIBZPvxX6kK7AH6xbECws3Rt6cK+hm+
zqE/xXeTBdlIOvV9RM65VzE7Vz2OB9A9WOkGAOSGEQgcHtWC81rZtp1HAf+kZ+gX
KpCdSiivcjkSh/IfB+G+ejShv1HrPV2j9yPkr/jJLBZTTcqJh8NDkIQCO1GLlCsA
BC0z65VGhMCmwFpLu2DbVPc+dctMeiaTg14t8C2T08DuuhBma6Ruf+zCZhum0UaP
0Qut2YHde0PzEy74hNvSnpmAQCQfHazYjlaoEVkJmEqfnEdTEkwFu9cjkFZB8Jj2
3+QAo/76KV/bQTPRFqEZ4YiBigIGelql49dFVEyBeHLyS8I6Q3KjZjer8caYXLCI
mC3OR8ZVa9JtnE9l3gw8CnJKutrdutZMK45rOmlp45ljMoy/Baf6NDpqmo1MLJIy
RLJMD6yotyBBWgAxtSGhTpaq6vCtLSIgys9ovHgPlNQJDzZRzHkh0L48fJ5xYNIa
VmKtsjBK4GrZAYozpJfhG7HPq2jQMupnVPKzJCiCg7mhnNzF9VyOvIkMemsbgfrK
NHdwvEJXBVglL2rzWkQTnTeLWX4bDXmMTr23Fox4/H+3+mWar3UJjkoTyr5mRduZ
0Pq3b9bOMWmAWvfHkVblyUBQ0szBrynFLLzFNJRP35zwyEGEXWagk7ZioE8xhuOY
XjxxpKLBABcp+WQ5lKSZqi+UactN/gKT+n78p7KqisvISYTsVQoSueMhay1wvWEs
1iauU5zhWNBf8d0UTp0XysaWd+2scIOHXgLdQfk4uqkcu3ywafgMJqJSaWF6ekKn
wYLgaiyq3zronw41TjiF1+n6hyn/r2nQ044/B5k7Lan8OMim3akXD8Dng8wMpfy/
14KPv0xBawRpW16a4gsVQ33Jvsm1YQoncUHyCopyWxULfJJeQ41M1bQW4t3cCgkw
EJxtHWFeSZ0rnK4amZwHfKvjCz8QZKlBqOLeEtFCI7vNafIIhMI5BAVQolQ9uzkA
rCQQnq9Ri9qOpSogkn2K9A3fJUZJeOp6/hlPGS90ic8Jrtc0ACQZJChwwUA+1nNG
rlUkziZC5ZBNBeyZzVFcgl+7s6B3fNMBZmyBtI0o6b4Ksy79M1h5ibd36xz1XEGC
q1VIuj4BQZypq4UdEl6ZboD+yGwrGkkfQryRtPT9ehXIZQRznB1p+uOFkVwRkByD
o1rwwykl9ZUXNN8HIgO8s4D9S5tsH+UYvQPPxz/pXevLxqnUf201VjTdxRnbHAks
Hf8PPeh3uLp1cLaPH7ErBTRrK68GAsw5361oAD286CqlryoVRHjGUp3Sv/U2Tg6y
HI9XBoBMUfWkQxQqrINdHTCWUrAyxEv9woiXszgXQ7E3YbgHTfcb+b5QYRKdb4/C
k+NEEsJDOQa9HrRXyzoMKaGNhbNiOJJ1Aq03wb9TjxI0o8cR0riyQSf169WPbIjm
efsIykaEcxKLXJ9Oqcb24QigS3G8PaqWwKJfnU6RATWFx+FPNh+vnvEPexW1zhnM
duiZerMtACKEfbz6t2YGE5FDm/fS6wHBmrfvfJ7uSq7A7relyIW/7xsvgNkN11ul
im1tIz4Oj1yI6YJ73KcnPIYpG6iMEWAE8sBFgsH3fgSzWA0gtGDTWFgvxAtSsrtz
MP8pYLmpixBmSeuvNwx1+M/YEb/kVeHt+AzmF4O9xU0klMaKABZazdCuL0hM5yjg
1M+UnZEv4fO9VQXJ+//tJL9Lx+B9HEP6WWV/8zyJAUTi1F0fjKj6e4j3QdSxc/J4
l0/vLo18OuBlAuGuktkN2WhOLmQJhs3zMXehviz3VMZR6oBlHajqKgs+M9AUdPek
QXTTomu78ZCvXFvpM609FQXOP3R3FO9kzr2s/FAbFDE9LAF1qNAJpjIdU661Scte
pyjDsuCQBbvOvUXmjW6g2Vl8dy+lqKQ6Az1l3lV6MSMARHYrXkUEIYoHSCYqE3ZV
VXjcPzDIL/OhmbobgVUkozOxCUf4p3s5gzu+rTlhm6mJY1YzmYkfVU9sr8CVZ/6m
yZTw7N+qnNCuovkOGCE4Wf6tEw0OiMkP9zN/T+KtNsmpqL0cyGNxdjw7H4bQg6Yt
eURkJnKHlKGpjxZ9b+ZXann+WEUTPAIPNp8i6ecXsfSvgvDTomdd+N4SWyd7UKZK
5aYBdS+oNbZr733OI2T66BHLRPqmDWhyifVTgQ5snaUfjDPYoV8NVm5L8UWFsRGh
KMQt/AEClJ6plwDdxxsiYvBZxQhGANIA2RJWSVYlk+DsS1g1A1cRVVpwxTF64T72
b5hjbK31L0aS77Jjk7osWNNgMce8TeTZlaGNU5fi7jkUu/zdfaId0Y6cSqL/1EEY
JjyB6MV/jPQ3W4FIwLFI+TvD07IoZb55WMItxnEl5m+m9zAGHXoBOrY1bDr4gmek
BPVl3cw6jT4x8B1xOBAW30sZdM9sngCJeLQ84SpTeZolJJ5IBy6cAl0TjAy1hHK2
kvxkBl5V3+c5ZJCQZ19vslSZpJT6wMBuNdffwiT0TWp+W2tSf610oVri4nS1ABEq
W32O5UuxAkjoSLmNbwptrIZjYxVw5nA8fJjV3fe8d+g78YyI+jF0oEIfMw9jhu40
CWaDRvBUoyVWTuvqyGPgxps9wLYU68T+Zmw/k0HkOGlqrvyRDCB172zxeWaeIWXv
eRCBMKvitvEwPADt7YxZSRDwP+OV7tviErJfwMQ3aQLBkOVdixnFVCGuw5QO+Sxg
iFJtmsf3qzmyCVYiv9CagRuwnBw6u4c7HX2O3wSsI91OiFSXsbEuMhpqh5d7jqay
ek9kuw8SsOjlhkhQ3EjN4xubhTnvIF3vNhrRlw2OCgIbTyo1HeBZd7uLA/BJL2VL
IAoWo+B9bnmP2TD1ekreE6ehzlT+tae60ghrYBw/3dhnuMRG8krrnOAVmzant7Nj
XnXTriTuFG5/ZrmAMJLI26OQ3l+gY4eIa+pWs7H6xcJT9hiiau4s/1PMjeKVUB3m
qbMi/9Tal3JY/YfQAM7IYk43k5NoBsLctZhXzHqTOywCC4EInIdGLZdyLw6bXZXC
ktBIcjLwd8yc6FPFw9y/fsy8G08lsmt8WAIQT8o+9I07Qikos75TNIUZY00YlVJp
f7s4XXBs2OC0Onc5TM32TiDo0wVPL5U3YAyWodL+kzlFl1fuuVIW4HJ1JZ1axrP3
D42IrpdDzJJ5ypvCeXQgeUxVaobcgwDZaYLL9JuZkWXQGsaxINapzhOKiEnbk5LD
wXKUF1YvFX0cpzW0oHrEseqZ2iyAERefThri1u9XAr52nuh1lxl+Q6uqoX2/CapF
McFmVSsHuEovUumDZG01C0ID0fkna8cH9DVOG028PnR47OhdjZ5OQ4Ny8HR+Nv4Z
mOqoSJBelPnGF/atLYjNKK3hLx2XdW/78rpB/vK7lrrutfXNLVznbi6FGcTZOKBt
tY6DV3DqSWALqbplhAlWwVKJ/CWsjWrUA5bhuDDsFwcRZKYc7fME/X3AmAb7c7LJ
h5GEg9QVKJCvwfNjlpggsNwc/OPsAnfw1HpEdxnppyqSfUkH+LIOW13iq6vd1bpW
QWnmMF/OU8ej2+hS1XJdJyCaONNqBu2isxf174BzE5l0wgYXbzbbTqDi5IY25p49
JltToUzPNTF+fcvU99XrnauZmpUAylJkyOMF7lXhczLz6aFAn1w2xMzzkLo4Oud0
NfxDIf/cwBRpuTp4eE2n6Y6111k1wpRwvdttNvgN5iSr9x1WOYOy5e/14nlFKbTO
5kofwqvOk2yj940J+V4aq6+zcnvnluiFb5cWVoUxCt4+LnOmggQuqG3wr8szGyZf
Uf336bRxYxUy0fMvslorQni/B+OD2q/bwcEwxpF7uOICHNxHNzKoBxWlrql9vRg1
ihFxlYigG7lNa5IZI1l13jfJAbFy/w0o2ssoklOXQzh7FHbQ4SPXY1Cbbfd9t9IG
ttV1fchoG3xCzKMr0E6ro8BbpBkY1GlwVVn9V/pEZovBR2T24L6YgvW8appxXDWT
AMJNfrQ7YyN2Yc64ovB23E35oW9e4z4QcU2zP6YWF8LELnE/aRnt58pgaG8OqbZ1
99u4vzzSsUAjGj9KPcBee5k2+c1SU4yjUQ0gu+6qg3AAl6Y8rZJIL4etXitropkd
H6SUyx9mB2brNpn53HD4Vs33BBpbcef/A70ZHI2+NOklzn+0atiTyLhV+laRalSW
344Nkxw8aZJmy7uJWfgFxYS81YN2dyd4dPfIo17LzpKL09BJpDhIKSU9eDE/MOXe
ZNWJJ4BwEeeQ89Mjb4jl2tF0sdpwGVmMkOYBperXf0kIglanQ/2CXjCYvvdLiGag
vTgPqop9mO5HGqeuHSelcaIC1fqGOjThK64Di9NHwaR//225hpPcHmd0mB3Rr4r8
DRKyp2aeS8e02aOtSIxklE3yUxilhg50XA6hEswviZ3n/0y/q3RgyIums986K+5a
lXCyRXNu3ROtrBG757Sx9HqB3CKI3EkFS/WrljVaJltSKCGNocXOld24KLAOD8ig
NHERF1ebOmwAqa1y7XoUtUgUxreaj8IOEAhhojWdbQrHgQsOTdpEfiU8H1bl1tCk
cr8QoT4RUMKvPNR2AGYBX5g05LuJI0fh/qGjTilNQsQ9s5UxrWL2WfUeS6SKf5b5
OLbb2fQ7GmIh8FAtLvSfRt1hwmOtnrbnvrozkySyngTtYGLvr806HqvuwUkiX32z
u3W/mQjQq/k8EWQmkXNde+29mX7wTGhDT/cHX3dPipAjFAf2+IxTHwH7LB4f3Cag
ODmPBI+NHNFCLDmtOrME6m49J3oruvttDLEYdEllZ9ar0zPO1BVXcRBd/dXqYLqa
F6wv7aDEg6rpmp3KURQRSnuVCrWCLcRIhLQUQJTJv1X3H/mipHNMPKSbhP2ge7cL
+mTZAeMWAkj6QkAHTRMv9s5ZlAzYUlqe8A2ngPHU0C+mVf2xbktPuQReGphR8Uj0
7/TNHEM7zfb8WEt0BtaVUIi1f512AOHflATCC+xdjWJfNGpPPoFklwFxxNYo9poB
ZKaAtdNT0+TcOALBME8cEBWVCDFA4ouCuYOMrEphH1BgcHQokgVqov/72I62+Yul
lO0d8aisL4p7c9hGqKeZKszu2qSRqh9BEJqOTP7G/ZSwbSqMXjUp314VzWA8lAom
O0YT2Xnpe6sC7ktRExl8Mto4NySB9SklcGRunzAubmzaxX7C4K0Z8x7wkhPwD88C
Wug4IoTP9oo04VjcOkU+leBwWRrOw4auCgXIwb7d0+lJv3pG7vGrnACyD0hZVP9P
uKkf/pyNL1B1TODq4STRdQALRy7LUYUlN33nVpQ4Xto8+K/kOe1hu+HTuU/i3kge
ilA+UWc0SDWsVpji5qNI2aias/8lZ9d1eJtXFMPXR5AjPrCQ6xmYmMe3I3PE0dWk
aAOdzpiMAAkI/i0IjBfM6DumjFEdURZ7JLmRRg/wDCO+kWQXponSN++Y2R0r8OGj
qopQ4enPP2rVxsxyjsahcxTI7W/3RbZd5KJU+iwc7gYpjyxEGbCCIDMPcRPcjrvv
TK/gSEnETN7we1wF1Puf9mnCuUllYvVEuc/e/YZTlQEmVpKlgMmk0oji44alKMbb
xWgE5SIh7PWB8VbT8t0kOzMOt3DCMYKlFU9f9lt30qSWe55qRXalJUZXSJPQcQXX
KvLnnPOsN54v/WE71VvpELuHPiiu+yJ4HI4K5wm6SC2WeODBX6y1LdCLJtNBZCRV
jyDj8fO4SFxA/ehep5zDbnIcVOoLqvPfudFDW22S9/+31s68zPScsPCC0T25uGoF
0yqWF1dsv8pbj+ePiZkKNB7Rltyiwl9c3+aDWdiSczLJqwbyII0icNAD6+KHaKLZ
TORhHELBKP4CEFupnVgGrfpn5g3miE8UzbcDg91lBF8RWKVTnMz3Sri75/PbGnE1
Ev1YHB+JZJsxGrVK4FcGVTJ/nSQILujogBvceaN0iwjT8/pd7NJpZe04FeApZvDi
8686ksDaAJcGJyR/JzGwzynK1rDhVdWXJmo3Vw0wuTmVsWVi5/9inYwGe9a427Ic
2ktl/mXx8IpQ8qaSTNoPYVJvH3ykF67VXq9pgFtxSezBCDPpvAb7mkB1Pfg/zFck
Rx0kJPMyo3Pi9pgHUdR2uaMfMjmoXQirzqdcdrMeThhzyhTu8+Ibz2x57TOKhZLn
WDkbC8D/8ogl7jm9PXj8ZCKaiH7ZSh2GfaCHFv12Ppfp7JWdn/tVz7KOBIE/9gkq
O+nNWeqhLz7uo5uot74VpmH/EOCjGqPg5ASaLCR9zdd9fO3vrIjJ+3MlfqGf0zly
0P3hQFknWAHrpkNAb9JkES4cVrUyzrXpeqEWrzI7twZzTICa6jKAVjB+qPfGDFj2
Mg5ldffLjX0c/zwgeuCHay/E8FAnafYIcdKJaF6ikaAC4xAxD7HB3P6HCjRR1y7B
JBIm5SwWpQS0xtNsFjgDrzI4ez4+XcBNAl7ZR1poBgSJNqav93Vym2qKBuX1Lt3F
t4FiwR8d3xBRjB/LohZNrhBWrkAPnWbqIjitr/hQ2Mkh8ZkWaVXmcE/IAylQ4giK
BvfUMdU4tuhwuJ+ij1OVXwXVj+n8KNeyYMS7zueznw1790KB06OGujnEIpUW7kWx
oV5zko4bKrbHfzGtYtQdtxGrl3boAvr7kIS7n/MMegEXebgZDKV7ECGr4uH2kn8K
eGaCVEPHXOlM4FmqZVRJRz4GSmTiH0wRfnfcsZjgYGJqd405XtG6PhslImK1btzX
Kiibzt9CzhI4L9dHJQDsbghija/1AqXKvQTE1Ise+SVaIl88QlQ5aVHIcVJWbhpg
hjQD8IB2xJtsOODDeisaJ6ePMwtuCjdjla214HWdYOkL72nu/oemI+cGIOGmSFWY
YeGeXA9LuFGBvomKma/OTbxLXDSlrbSF9SmIGXv2s7JuANUJ9bVclaIE77SOMPRi
kUV/GLTlbIQS4oc6LeYXB4Vi8BM1EyRC3o26Aoys6590/wCvF3qgXGMZ7pTOe3xU
kpxLqE3mT1+7iXj5RN1NGByZlu8RZ6gbDmaCHMAiJFtDE+eL1rj1Iz7f0uuIcubp
3A83+ub2TOXbemlUKoTwuX3akG9hiT4HbgidcZlqGbS1lcvcb4rdw0lFqPEe7htP
oKUxjQ6aY3LKp7e1NV4V+lEPSWL8EQDDeBV9Jd7vDOcSF5h8IZLL7CLtIPI2m4wN
YZh50dz8qY1gpuOC4cMwDNTwvr0nlExk/uYLYT8zdB83r5HF1Krigj/a7+TVtQQW
gbmSMVO3K+YJhaagjl87ZiprWGxOSj7nYpwKalytn/otjwaPy3SlRjGgWe2axiu6
nyymtbjE0F0UA8BujiaXDsqs6DbvfPMT/fMs7OJkItIW9ClNQkxzR6lHqvAoYiaH
zaFFqajFAq7qSHZ7iguzDGzBTUP3Q5htwH8+qMYu9kNSfZefp+8qcEDHvpENySkQ
Ieu6qL+y7HerEobNJ4HAkz+0NP+8MyKZBeU3d/hlGQ+ZPKQ4ICojaajh36tTqKj/
qyHSfliFQE2CNHzs0M4G/ntoV4zfc57aFu7I+2qVc0ejZFP/Q7mIvgjuexSKiP3u
oSMoIuXOFD2StW8twMX/XW52zjbyQuyEr0Jc0RZsqSzaa5NvlXR3fTvRvAdIPTNJ
EYy5oVWL0LTze1uzlaR4jTD9pTFtsEUGW9e4NuqxPuHxHs+kunUhDuWdhEyUim18
IH9BmcwtEnC2WWo2ZQkXfgJm61xchTTToi6QixaPXIH3mzyzNPmMdCg+nQ8XIlXu
AmBfXP+M4dGoln9oERciuR7ZEUoBkuMTT1DRUDZq8kXghBsK+2KGFPG2/ZDtR4WV
G5k4R1ccDLq2v+pvF/c2wHQkx2LYIV0fw9Zlc/YnhkW0ymtRXdItGYLni5uy2om8
pzmulBHM6Or0wiIjq8LxgzPbmAIx0lZX/IWh83spA6Zp72sTWV5KKnnJFbe4Mokr
qZQK14uGELuLynqKwsV6DS/PQNOCuc89Y0PzKu/up8eM1r8zX/HceYEWLyuLYWsM
SLduLWIjHh9sDZsKXImUtNbP62VDzLZl1E3h2yTK3r3xQpxcy9M1kNsJBT8p6/hy
Tn+OYTfPcXl42+YxL2d/djRpu6i0tYrFZkjhRPg7kC4ZXrliUudpxourMYK21GWq
blcvlv3yusZryOIvFl8ElIoQ8AJHhnMvrwM4w647SceD1qg5lRPT5f5fEL9xfoZL
9SeVNAnWVwEy+vEcyxQPRx2DjagPBrNpJN27Axmn9/Nf2zHmugOJeShre8RD/WVz
lI9GWjJw/qr5GSZU+6nopLfdzwM+wSjij375bsDNWnf75jqv5SGOBhF5aCcj8xC1
Omr6hHZoDYTcnCfA3390JX6sKfLIJSG/xUW6njeJm/3o5iNXf8m7+rRaBtHkw+pA
9/cOY01hTUkNF8oS3fht+wUQiArMX8/ZT0wRQVFXGkklbkDEEnJurWA/239/4s0j
T836Gov0wiaFz0wifOBKnT1q5VuzowADzYLpLtp9Qj/2gRXFYS9V9NGx4UGgsjwL
xiUYyllSU+aD+9hU4Ge4mu5nkVgW8RbwvFz9d+1yXXUzL5lDt7Tlr0X1/afmqPnE
PO7gGWvpWab7fBqnC0IhJUVUuJTnXFRu+SjsAcRLN6rp+oRW8gX4YYVzThp+8cMa
XTZl0rNBD4kbyvpdbfLRx7JGoclFCspR/37ZZVPchCamCofJ6+urJQ5N2shzwAmM
/CXfA+XdfA6TxoDZLNmtWSvXPv15DOhCmNSnZK3iv2mHvMXgreiuU6ynjTMi1zIy
Kzh0aqM7jhtqKP6/s+NjDHzEesBDb8jdd3HA5VFvJXXnVt5Uuy2ereszOWMGE145
p9129IGFT/ftU0o3FK7oYYjaUeSGr/NWAQQcDL/nMwGq3zzX9HzPL/zWD9HbSmX/
JKLH5YuPhSmXn2RI6Y1/DuZ8EFLO3FaAa8I15azyMMK8d73DennWeb28Jzkdalgk
6VgHO1jsdk3X9mKnjBOxtKHU8/OI7Zizf58G/O0GnKuOzBy5ODWhrby7Saf62X17
y7tIoBnpqWlV84ROlDg23GDbQdQIB46+yoS5iwr7FwNwaBaQFr76/r7AYPpwByUT
PpREkxiThS5HkkAsMmY/6ZyXx5PmtcaOD2wDtj+48TLj07SWI5aQxxTyiH7WRQes
mJb/bTEEoN1wnjyuDhvtlpVc2I7fdxk4sOG/w+ct6LBZ4AB0tCYu/e/QG+RGPfJB
DgbEDZtQTQUznaN3rD+hGwl49s3fvCrBaUMiFoFdNsRpjKzP45ti0b1G5zQD2A5h
KEZlXTTJLDh7sR6IQBpiHDTuw6cevBRn3oPyluXB5pJu3gKnDWFGo3/kYRkj5Dpp
3dx7bImeYDVFeQcOQ8ud4A==
`pragma protect end_protected
