// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:42 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ssciRVeV0fQ4uyjihe+YFJxLaRanWFqCaPPfruXk8zWl88d4xjj8ikR8eFGc69/a
xqT+OfUpb5HwzHeMh2OVtVdFfRa0A9/yzOxvCyJOfM9/iL8iAWI8bYk9hK5j+4he
IQGhMzC6Q6WuX02zTD55S5Awb4vCdELVf3ej0cb7SvA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4512)
sZ7o9m2kM8ItmPdJc4cqeuW5Tt+RRP/DGGXRvyv8TzU6jTmTOopoee9xMWJIv0nU
ErlceXZSfN1p//26uwdUi74ougdlo4AHNoZCk4gBqRs6kGy7PUlWZvbTOW79tA0o
76uNUr/ckvDolRMkjJNkaEZTkl2ZBtEIVlsFwc+gqhDCkLlWjR8Vpyri1LkvR61X
hegnrGgDWt+jlPmH1OXxgCtEXxolk4fy1RIAMjKLCZNuBd7vdC/ggGm/R2i8yAQN
qik7GYwi0k6HyKNc8eEGL7UgMuMHFvm/O76fuTgtd+8dUYq4mcXvTNA5kqIHVO/H
vi6bPso1TXFzqjfb0KnegO+Rq2DGjJTK5eEh9pmd3y1Aj54/zu8Ry2MOd0hcSDhz
rX8iifC+os1om/1DJz/Hd+GVSjhKiJ/E1JD3YCWqPjPNOZqkQdI5VHKIBq9J02lQ
gIH8IyNhyOIB/527TD+J1ErZECqp+JCH6uxMpRyZ0h8bJmBrpZcE4jN++WhOwmlJ
p8RyF02T/ghpinRF35HwU6NlwYcRgETaCHR8k1rkJY6H1vcfvvejY4tHDEgsZtod
R/k0PJtVbKPXXA2RELswyLt4Ci5is1sJY3I21L421SczTWEEYSIAwvQxEcRv0gS9
47qIScmbkLWuld7lwuh34YiCT+hwAB4NjtNsplsXqj1ezH1KUETBZDOAKUNh5N3w
szm+vXjHy4J/81acTfRma8hSt1YUmP4Ww4lHHWXQMjlskp6NFfQ6l86XIZ3lR9x6
Bcwn3QDEIRNG3pbYtPBGQhjZCAcMvEnbfw3bZ16QlgNMUjozr/jt9gxP2251KpFD
be8qlRxhpWYCnEEhULaX+w876qQNCEoR6BcbbSBb/KCDlaqXwkmd+G8mAFQ/6u8Z
MH0K8nBTVXG/7S5z6MjwhNSyMthWr7CC/GS463+ILTOLhFS2my/+I468efR6Dbeo
NV1jUr8nNMeEEnrJNDH5S7sYikexfdA/i2o5firHB7BLKJct/uLNs2AyMD9vLYvU
1uCnePImLFji6eMsLLezcBvqr6NyLhM/OnReJnO811WYL9nQ3eIummEhcjjapyhi
PyqZtDORyQTsnQuSSs6WcI8qYN+uwuZWgO9g9WMNmWJBKt9yG07IZN1E6MO6Pevt
8TvQPtnPYuYaDQyMIYyUap+5V3rNpS7xuThFoW+zsULq1UDmQqt0bPLVggUhtGrz
oCAqnPhnYgXjTnUucPZH/bFJ2VoDzpEsocVnoR3mYVcZQkTvjD20hxvAUGW9jOUZ
PAV9Dlu3kGRe9q2w0s2/Y4VPFSz7GHomoOBsjG9+jSucpHCr4FzqRJECntvRz3cD
yJcFhBx8zDeTsccIdGNFkhJ0UT1jSr85PAo226N3DPsqOv+vp2UVhCUPzjK0co9M
Wn1LsRBeP4b5oG++zUZnhXzTbSIMOxw188axhbD1glemQ1V+hrvHIneMZou1WaWU
vNCEYIlt9YtxaJCv0F12cklJi17l+j0FmzS7GGGea9xHPt8gFyJtB7/VufL1aaMj
QXDV4WEhmGOaPTrcQngs48B5ToXJAN0imZy5AEaLGlNdiOlGMiTnoBmFv5MWSDPj
JxNi/j2WxDFLAy4WVDDemVRzVo26g3GU3hds3uEXFJ3kaOhZy47qGYt5kRjdOdd9
XOy2hmaPXqK1v1AiS9E1B01XCU+nXhosAzYfhjtLLQX45iPG4rWOb6UJAwZCLam9
/6WzdTBYsxv+4LNuR9DayRSPKuZduiQBuh65XbKAR0rJDOKfhyDtnhnFzWAHmP0D
TbbGEeEqUoxBMMFhD8nKRIHKKBJLQjr7iwwQ7Lyx9N8NZuya9Xs776tcJUprwl0R
dbRJwes9aHNP00iD9Fa6sU114yzZUxsAtYR1EOhlPO2+5UNq87J53YfxVsSQgN/x
kLnOvdIl6jmh5RUy/kzdzBP00kgwhC8GkpYLNMsoKCGpsnh1MHDLp5rx/Sd/tJ3N
lrWrq6vkc62o1GvtxKHAtXpDZrgUwa1eTtk6pU50dFKPZkt/XhYKLkf3jw9zDdyw
7hIvpg7viSRMeJbTE5LWkXuwcSUK4XLKmqEuW0moOvVNhoZphUKmJxr34nFFvl0L
DMOmrConAy3nG5QUQK862HV/ALM4E/Omac06yEJqBmtbUIFGtN2h7CeY6mLssdq4
Ri0SJsIH2xkUTkBx4/6M2eLrOTeU+c847keQJMdMF7bN44f0N1wdanIkv1JWvyhM
9PT6aIF5aaY0V77lnloiqm98KeMW9IKbL0fDdoKQ0wE6fB8bdE7Y/JAMzqZXMfrI
aTzIDb88GAvAWfTesKfhIRguDW8nkGTbY2dDUsDy3rioYuRnh67EBeYY7xJuKsF4
6T9Jss85o7Aym327TtR4EoJSD4bcIvV5trj3CDgAgY6KvVl/Ts6v/7MBAdFQQTxk
ViF9aNdqPMusqnZNXXwfy3ayuxVK3oLYx83YukwLZx3GzWSMhdCDp0t1OOqteOq1
NsVUsRy4nH/aKfwKLo8ZKoWAXVD7YHy/M1PpNM2Z6KxTPQGR5Uh80cD36nUmN2j2
i7Qmxk10rn+bebqHduGyJzYKesbBiGdLrM+F7J3R28aGLI42RUUcmHdZOv4cdsEK
3xy8MsgLNGQ2LGmeZ72P7f5MOhUHr/jaGRyQcmBg3kGOJqRzKgBBCbtGjYkvBtNZ
OWIDN/HP+N6zKzjX6N7aGXoOD4EWP7wl8Db89nJHcBXgGDUS9Frh+bxekx75aB9z
95rPfdMz0DQaOAD2ng5hjJuIh6xzhyhZWyc+wZ3j/vPZ8OLJD3OeohxM52Zu0Dnn
nATp9yBf3FBf2ODf3JVnLjZiQR62HV4UcsE+2LwZR3FQ7znN4fwVSyZfSiay9oPW
c1Z1jDIMouiqs4tgR5xjPc0H4o09KR60SAd8HuIizcvNupc+a4QLhlcTP6W+4DDH
+/BGzZF27WoMRav4q/C79vdM/pffs1hsd7Mm+VHWciHz94E8qv0em4yoCOC5TsMK
oMJHyiyVIwiOjoFhb9kHoty9x6Ub+ZwLYPGskybiUmQUkVvjowDVco5GFWr1uh2B
6zbcuOkyRo7Fm+UOmYsNH8Ry4VAZbnPrDqNHXmVKePnuhd41ZDokvG7PMsyKFyfE
CRcQ4pvbEwuzqghj0SA50L922EaWyof/3cVtQKHWKv/axoRTwZDeDLSZgJlgTdZ4
cc6cXsfIpnt4uMkEFZDp+INDYTHamh992h8W3YzfGT6eP1MTQpEU1KjMSEeJzMns
T23TWRjqHfnz289HYA7DEGJaQr2WjKP86wEpqIaMe3wP8fNF/BngnnsBLUpwVTli
x4VZ3XCaIJn6ZfVT8asNXjBvr+7O8xT0kL5Ku40VkvmspNT+KHz+DOWyE254OHp0
FTHbVRZiGFnA4ahkvKiMJP46vCHefm8T/0/D6YtkpeT5MWbay5wm3bEPMAikQalG
SfV1tiziirUNYxeXRUSVVLZXEmL8qaQpAPfktZ0Q75PbanNY3IkZCahkdAVaEj+M
wCN4mgD/1g7OrhZFwtevFNG48lJXElM/vwMNAD67jqNiDeGBsOKL7MVzX8pR1hrw
DH1F+eAfEnHRayEeCNotX5zh0TjdU9fhYQLYwRetNzVGwbO86r3eAm/xP6mz1CDW
OywSQ0/flnL1KbCsOILWFmhtX4a1YUbSf3FVpO9eh9/dOUJD0FIJF5kl3SCWlz7Q
1Gr7UXYDjd0OP2UBzjY0XQxPLzSEhBmS8uS0hWl5s6r2ydQ/LAZk/Qid9n3Weyg8
6FnuWuIjIFQUMFQJ+fyknMW5WX4gpbbPjF0omccrM7nEKGMyxp8BmHwQKBW1zyUa
Ad0VZ5bWiKJSC/d2FnoA4zzxqXa33gmpQColmCuHAqMqWGHHtbsJ/TD0LdrISjGI
gGO3jzUP+puIoNUO/IbFZNt3ju/GC0T9EBrdX9qiEUIeHYXWm9o2B9seJaEVN0zI
/pNRvLINVGpKA9+jpkGNVJxEsPFi/35Rpjnewpq4vKgucy+UdbkpINKnzPOczcbZ
HMgO2HTis7QckEpkJ39N8d4OWr/j4M6hxNn6m1nLDkbrTax/OKPg+lt0UaArR1Ak
w/xDBIVCxsVQ/QWSz3vMXViqHdMa2uL2DVN0yxVteENIrxzAiCmAms104Nf2HKYi
dlv1cVQjPSrzXONOZJTeDuxpUr36Ma2HZtTpE39ytGL+/E1yKbQhftpgEwNHg0SQ
R0JwrWBK5+HKTJVjuSJ7zPxCjzNnIFvFXO3yHUHeh3SBe86MFgn4uMrjT4/RY/70
f+XXI2nrvgqyNdX/MdD+7Px4fdCZG+7MwM468nQ3/HYINYMbMHn+6Q49AXYCXqCY
v6aiDdCPH7KanqhlSPQDb0t2cSAN83edEI6yK2GwDsL64sZ0SubSrf/9wSN3rGQE
Skm1NBzTnDyTGJnh3nk7KXWe6K5nzhYmH030qITItz8wY8b/1NXEiLEFqIXa6sx/
m3BRCxnVSRE3J/o2GPqS+BoJdsL5ydbPxPMHPi2DCYqgr7I+vCeaZ7eL90M1ZDZ2
nnBKpO3B2BQGAaYugZ6Z52LH22lT/u4ICa0Fjnjf9BR83/sw5mQ46PehE1QwhQ2W
HDIyCLoGu7/eBvSJSfxtl7SMraigu/sbhLUC3LQrxLwvoMvh9+i/zy1IWvbnx/qY
2OKsUf8BH1bQqLbolTY6KTWWgELvevWvMHBYD3LPXQsaMeICZCNrekWrze2CZfCT
M+dSLPiIxO6OOVzRAQM9ZwGjiwXR4V/TzjaPZNqE2bqSTdgZ4DxWt9R1NvROohsG
rjKJl8eh+mEbmuSHsBtgcr063lQJngzX+pKu3VBbeTRIGJdYPkmFL00pRY8lp31s
vpBxN7aUlMuY7tzxToIwFZykmT4yeg8q4uG3utBQKdpPfk0bqnjrMzpefbCmIkvO
dFYm4b08wQvZzCvhMme5ch8NymWaTYevLx84chmEs53IwhTTZHjE2YpkGJ40eGNN
jX68XfqnS1wT9J4sUhto2gBhbd5p833+rA2EXYkQW87Xh5yeagxrKXvAQ5O0WWho
oTDeBi1oJPcTDHP1mU/zRbVQ6UtlqzV9931nOAW8sYDOactZdWvfnwJkDGSMo4qw
J2Z07oZCxD4KVR3B4CB62v/fSPExvU5S2OGKlm4unRpog7NrYErTanY9KnBOTrWF
jlKatVDcuKVQjTuD1Hug3nuDYUNZ8oxlCgTRMVLqnN56sxyucymW0O7JL4lz7GAB
1Ch5nVQDoWoZTVtFUiieiu6lnetAml/THp97M7m2B+TFQviooMt/ReNZVwgdGNyE
eC08T2rW9SM8FTaEx5if5QNWX9D/ik7IYIIg7qAOZ3/MX4x/+3zW9nsvXcXuRXVq
zMhky9jo9mQK9DWTgeSFIMpAXCHT1pMmX709v1EZt65Cc9Vh5rzitqvkJoqVoRx8
3a4TmCgtApYAJb0cFi+YRXVr/bQg4tXHEPvL9SIzli8kt36dzH971FNoE18z7VIl
xCGxVhLHu/cgjqXMhhZByy8QZA3gp8F2ancTqu1XbiI/3dC5inUTDB5yfpltm+SX
zntbvmj5+UFIc03n8uVLOxLvKHtPSQEsKQsH7Wm7nboQHx22Ir62PDYxr0X84sXz
SMzlrDIy+d886InZVkJAaWuYn6dB4HLWPVz5uKf5MO4+5uVOH91SUKSBwc9xriHK
1vEE9ynfMDKkhDgrQL1lH229QWpfjWR4ftbTgKzIglbWpDfLBCZUZecbyz1FPmz3
zP49TVTvTv0jAXUQF5gzPFsaS3qYAjXVeebTDCBb9ghjK8w+sqmwjiT9g+ae739S
QQKuHYmBf2z8CZTmCK/MavFH371bFHphnhuN1ik3LJGKbi1EG/mB7DqKPY55T596
fui9xlrXulpDMzV9UwlcgjdgmvP3YBSFdKDqRS6bgxfVUNHbrJKhRXdocvQbSze8
qYs40dYK4yNkFBout8gFmRfkhr5d/7UJlsKpGp8e3FiobT3wG7D5IqLHdEBCw8X+
`pragma protect end_protected
