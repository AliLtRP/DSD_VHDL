// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:11 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Tx9oGFo6AD+pHSMLna7GMxQ8iFN/pc+S22uy/9XEqjqplt/lwznBjeU9QMomNGWm
PNBON+/5/PARPkXVWvF2/KZMiVSNUMTVuZrMhTOKRZvOgRJK3u58L3dH2jptnZxU
msrAzexK6mhggvDv8p6dg5Tv2IFJFO9A/i4tiLu5QF8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25120)
19H/MtUEqRhtNuZVFxxQTqDJwV6v2A30YYrK2VpEVwuU160WtyyLsR4giksvfx6K
4zOD6i17S6uAZX0os6wNCJozOFHv3PaA2/A0BRR+4CNsxZXgGkLMH6OgTUZLM51s
wF38fr/I18ZiH4VBP7oiYWFYVh/raGhbC9elqeiCsaFb/EcPFxuhiYqrJE4tM9D+
9xu+EB+qOsmH1xs01bNQFH7DFFDCemrQTmmyJZ7BCJvwqoN201kkjCjfIBQIsnnJ
2KCQyKicBoOJi/OrEl36SE0kItVnmwuRMymsbq9YYOJQVLClLy0uuKktphJboRrZ
LJ3PgItWCe3226BlrriEy/2zm4tWwU4d0EZahcy4BAGl4/e/gW+PQfD9mVaIjg/v
Q3e4ixqn39jbpd4lalH6+fAhglnpbXgezUivfmKrjzlZv/dxEFg8PFIA/ViU5JX3
iDhvCgg+NDcbrR+3Ufc3y9jSnjYFgDMmUh3P49RaxglgYvhleq7A4p77Vga7+LWA
LHrvvxbTd40xw3+NXIIb5xJigL0EoydghY2xw+SNfVVCjHj7tjzwugynSIfq9SCx
McfBAtqLQSVw5nN0llY5V1QEQ7wphlPkSTNpbIFTo6bIIbwQhyUIzt3LqSzTk4f7
8qP8NDGrX+F44bA9zETlZvp9Yf/vsh8kPpDhPothm1VBlRq5KPd3zSoGyThejuux
9LtVqoK6TRfed62P8DrZ3zxR5omO8XynTfBTK8dt2K0+GEdFLIQYOuNm84d8trnK
WX8m0lLlLEfPcFo5TZa/4BCobBRx+01+U2O4oDT/zWU4ngCm42pU5VsUeLoIyhQm
Msb0fKJ/ehOX3HpQkxs8W13KfDWRo+sFxjnwbJblPxuSFjTDaHaj1fikCnHOtpK4
pmSfUigcyDsTUESKDTPvePgGOWlXluan51Q12wmbP0KG3S4j36wVn72ysgJd0CRY
jeXNK3UjoGELasNt+IhVYac53x/iHkWjwPT+Q4nrHKRa54j83KmZNiuZEOgP2ofR
jetG4i0Dh4kBA+g4gepW5wyMkrTBkS1lvBuzkxtWngvxdNL4PNi5Gos1TXTma85t
KmOFedid7l9/c/TSYRx1ihv5ehb4RLTImBFZXso21RlZItpD6WsvR0XNwSNeWdVU
Bx2Xg85fo7CBamqF5mtJchCChNqv+quLldrT/RiRMOsxEUYNfgCIpRoE+jkXpqMo
0Ty7/kxbgA9Cg8fBQgW3vVZohFxOE8T2TufpAdp2IAtinHqvtoXCw4cRFJhaXcEs
BMAeRwguej7UxLX+DXIH/kqyFL0w0e953d2PMYJ1ICSHqTECmr+tF6Njf7z5mpS+
RCtfOVo1daK7cFbQb2baVUVKQk5rcstqDMRVnmRPlQ5u+zOzpJvxgMf8l53bleq/
jno8eJIUQirldeYBLkd5qIgHDENuPYks4MYuAJPhHbiTCPoHh2APT13XlK40wbFq
vw0dXM6RGugwgeyojCU8bgTnTjVQleQNOblZAY80YRWtB09uu477NIcI4Q3fNqLb
Knt9QZnOvvh8kCKtU3P4/LkchiMO3J7AdMVvCt2JHuPOJqHH416M17ouwFA6Eb9O
qgERiqIlavuF4/pNLhO9wx2rU0TGtOjxCnUjcqmDZkEcWzUieavSo7lLJNEj1C5E
gajL3X262J+MOHf/sKxza/eyVlATV+Ri4czd1JQrdCu4WP7RFVLG4nEn7gLjOaHX
3gzSyWSv+k8551iE+Ibdso8rmBfc6190nVzOX0TMBjKA18s/otp90fNmUK6BTsNC
k9pau1o/2QTtYOdbdJYIqha70cnqAWBpgDB7lJQdiLQozuzPGaVrU0GZZLxXf6Kb
zqR2LNlP+0867RYA+K2wVwbJhU69TFtYLhbR7P7mKTyOAYXF4nrmEEuI3Vdb9eay
ebIdmlcc1sUjg9xy8bfhRFFGnqnAGsnlHJBYuO3TEFf8RXVL+4VnKeM9jKTlU3wE
ZLN3nsQVmYhPlqIKIJ9yFLtqiLIBflUwVh4/fLu/47ZJ7yZjKsYCV/iG6xXhnrlg
fllsV0JNnSL28buVud7dr1xgNr51vmCmwB5cuzHSco3RVwq06/rf6MrLu7fz3igP
JU3RU+r6PFEZ9HSnt8koPy967B1Jh5IdTtnxDCYlZ3t7c0m31rxU8zNYUg6ynIVC
aKmXqSk0fgNnSgk3U5JL9/xZCHCZWGnXLT+tZJBFmWi2Na47AnIzamKJwfAMpeRD
rZS4Bh8pDiAvan7fqZ9Oq+lo6Csj1XSsK3v/MY/sZPejFHjELL+7r1btyorLh2pM
JMAjOWjN1ILscGS7gDECoD5518DFusDTxWzYOU+vpNXf8jaFyOjXI3gJ+iC4ozxZ
uUxFUPBVzA01JoXkhdVGYzpAIveKT8pN8rL6jL7X0pSuEdH0cDT56yGU0O+oBWsL
blXMWEUHUs8TKWg1YXYigphAB3iUhDFq3jMw2QNzx8alOKV2xW0ZMBHgKr/AEXBE
GDsN+JriZqi9LgISRvAoIm1PK/0TwcwFtANEqDF2sYHKM8/OKnANNg9G5xgM20Vd
cT94smIihBcXaahvFD3oiOQG8+RWXnmjyXn4dkkkPoDC9Otbj6jv+HVv5MueHUar
PZYxZLzvyxRMxldkLKwUtQyTCJ5K7Fs+sbHEZKVJC1MmFZju1Ut+WtZpcYlVHqC+
5mGDMd9BPx3z2sUVJNvLmK3cKLCIYWrP7eb9BZShboc3GM4XTnlzYbRn4RHIcjVU
YubiTXNSATOU52mMknt4jwlJuP+IRfKLOYblQUw6gMIMg7YoOhnrCawk4ItlZsu3
bW2Yiu8mKGMkFJckSD7XgyIqmDOawcKRSOqXEwc1zYLcM/ecNQV4S/u3syb6KwtK
OmSyISmb29ZSWPjWahMuWvFdpa98dqOigvucfGpcaqIuMU8PLiSDU+OU12XxaCZ1
VKFrjnmjtOqbHAIN0704+30PHn1NPekFdMkbOuLx2skdJBEANnGTB129aPcsg3n4
IOBBVNJrkGYfMUoYOjDiSy7gyGkhQ6DqRGKl7XxtSUPvXTuX8y+FicjjE3JWo8F/
y0IrA/faT+5lwPpv2u62skM0mgL+B7veBXR2jFsJHLrXeYRGZuCO+Z99j1z2kgiB
MqMXvtBsOLb+4zbwIe0E3Nz++wGYFQ3gzmhx/JhFQEE4wPKU2WG1XgM0PpaVjpYa
Da1LgKSEEl+Tpt+X9rwxGEQMRYTGiMUcIDm9iLwsRaO5Vy/Au3zmOWfjDFHHscgE
qS1+TYeyQUpsRyWDo7oFnrySrNrQM5JufwHi3xQIeo1iYH8mOnp0FOMI8UOy8FQi
5WRU4WHobqdgcQb+ePKl+GxTl/tpPZtqbQM6KZIKkFTMuPMoY+2zCnt5kZBbMpar
YB1vnGqII09gV0eURVMsKKORq5iU6TSnFEK2RTRHzoYWUqQJ2r3kaiJqYkgTUbhi
1KccRhgPxYMq4hkIcy9+MkZT/HKvLPuEglXImTixtm6M6lachceXkICsV4OiQkSY
1G+OPXjopwdWVGHdvRnGs0vmWG7jxd0Rsx0wFtKQAs95h0kctayuMj9DVqhTsenA
E70I98mHVmnKhZIja5LCTDwEC3ayhNIX9HPTumZJzF+IWA6XI0NHGVVpUwMYckje
DJxYN3SOfN+equz2Qtcn6cG3MdLkp9RW49aWsbZmT4eOKoR3GsTSXRXVC1rN9CSG
Sask3400MgpY5W+l6QW1S35KxH3UqLdhi+Ejvm9J15dabJEytgGtveCseChgmXum
N7YPQdQOXwVaL/TgP0dubc0UIGgI2SvJ3N2XtUQD/W35ZhyuxC45Guo/nPsQ5loo
UvBIkTNJMHlyS4P32k8DFgf2JoFlTU4d0q9E9RWsFMrd3MelaJ4W6v6ZqhKTtOn6
GpufQps7U1h9Eh18IHJ4+htfThwCxjmfYS6+K8mR/KRQOQLkCrboMcGfMexUiYFB
AjZ7MBd3lySt0RQhKqHfC6VFlOXN9+c4vVgXVpWpmZRuUq8Uh8yco0ussjxQMr9y
ODQ4aP5PSIwPU+2vNZDlRyZma36iBwJfzs2Gp+rUgoSJZgbwT6LJkLmpH2oATOi9
NhrD+U/pwQBlaAEfNq3eBBi/MTszLIOQw4/j6ZoTnhw5QY2Cq30M0tT2l5hafIzQ
2OFM3sV0faj8OHzh0QHAeH9dOzH7RaQEDMYwk0GSfqswGo/PK+IlEs8ACsuGwqw6
HsffjoaoULpoVfvoYxN6vCmi/yHOdyFaH1kmEK69yIOnY87SXI+TDKAS3vUv/GRl
7DuQcPPqxT+CYwiKrqd6YQqDFO1mwGCqgfgcGoq+OQyDmF8TPwkfbdlTaXfMIdO/
A2T0lOLgm/A3mtirSIo31eIYqGTFhm7lm7t0kYziRz9f9UeiEHtXVSNHOPVeOIq0
1yTzUqbeKDlr3Lz5G9lPfwyY2R8XTlby5F/grQg1RaM3o9b/u8k0WSBRUu3NM1pR
UZJeJl03tyoRnXfWRo3QJ/P1nBQ7oB1UFPf4O/pt8kQe0j8dmvRYOm9l0blc3nFG
Td1R+itdUtQHgReDDUgXb9ENVwEBcGcPy/fzr++NmIKqm7G4vI7MYS7NtFH20PaD
D8jAj1M4i9xF1zOcV3m9IYE8AvRanSvWeIq6GQOaj3JJmEd08oXGqkPAcG+Up9cq
XuGOly46rINm20Obd3U8g9tjvNLtM3roKeShZ10Un0NF+8UrHVcU6NTW8xzNHHiW
gt5gNRGqXFsY0UXf/4+vn0/QNh772sMuIOp8K400fTWVXEqwUOmwgU/M9eQ3iZIe
Qz1WOTVPqH2lqdE06gWCLTDY+xAvRJIfYB/9vfVOox+c6fG9h/nd8UiBfkIUG3Nf
VQncF3xfMedSx6kzZclYM6kJwXBZlHP+XlId48ZFoF3922xjwahPQutkigrWC1ri
25hY0B+MQ9tGzk6CnuY5XBZ3ACUNwfj31fhw2EL8XsXm9ggQqoCCmBNuMXN7rsdN
c0xz2DmvGFMV8L2QI0VsfX1QmQlsNoqrYWaOdoUbwQ26eNaZEkydzvchhb/KZnc0
mCvnHjiXKBp9XrU3rpYud/nwPrHx25RSZTcH0TC27TC0zdo9f5LrwccXdpgj5y4I
aKCyOwvLyG660a/QR8h6aPbYwq0oZtt2BDPmBj4DlhyMzn44oWv+v69OjSVYwEse
qkU3SD9fYrlzOqL0iy2pVP4cCxREcVKjCLkMeVke1iV699Irfv1G8HhEOiuZuQLE
9t5vhoEapgGMMxh35mL6gOhNmOXaIg+u+Wfbb7bn4dFGA4osBXrbl9OxNj5K33Bh
B/mTFmZNn5Vd3CFihgcXh94pK4PCNyjQg4dmrhCEkZjIvKGHyCRcucMMUaIJ4Lc+
4dD85A7m+YNsYdWlmI3e6bFMVf+86JWqgB3qjdVlJ0IsBkwBJRBqKaUs58pcChkH
yHMibOTQG0lyzRz4CtY8wK736y3UtusbDr7gmgl2RHsTdxyY2VSN2e17FIncQAHy
DTdi/5B9q2Rg6QlpRchfvFte33z+4UwF8qa7NMiaQk8AmYMW2Fzyl3dckpv499Nk
pvxcZFzgzKBnfwstOWwo0q8o8UZvquTeZD3LOcS6b04+dX/7o/QGdZPseIuSKuAo
7alng61wcGkoNGODbw0be6syO3Zr2ESQtR6Tsa+LRcPsOc+u3m/UAcJs9f7IRwk6
ca/b7EFgn+TzjHKmHbzWy1j9d7JkiDCyXUZgMSFSjH3rmMYSSczUnEEaYR62mmFl
xyOt4BdsAYBfsa2XvBuRZ4rk9e/HPzoeh3+w9+6Zfoo4nS1/uiX4GoDHAA+Ihbmi
i6rTh7a3hADpeDabMnDj+6CHPatf0gIeddeNvUSFnrwDHzRy3HP9z+g4oprYuxmg
Wl8kYmqcLn+BcZHa5lIqf0PqUJmJjQMkydh9tZ/ANhbMFmApy8AiO8QnHvAvaRNd
RbcWyPLJHISfVZ9JwwpYZdaOPd013LeC+FzPcRasCCtFavzryuaNOOAfU84wV1Pj
K3YQ6OgEXvuXkMNUFGXplQRJ+euyLBQ46E/IZs8GQC6PXsKXLQOr4uN2fRcHRY4/
XmGIHZ+3W9CRLCTiuhFlnSJK4LuJOWqAq7vN7GSKL+1Mpc1rg0tTkM3DIZ3FO05u
LyC95Fp92iI1XSYBwv0Jm0taQ0vdEw6gUEiGHHlGkN1ETgRHTepauQUWr1Hv0n/h
Iri9wThcGZWTMgQytg/KjNWQlQZwYPvxQWj/K914I93Y9wLjA6jf8Fb0Iwv1Cm6z
i8t7fchen1b1nb0yxYP78JsQoBvlhNdP9tBdVoAhW3oYr90sPxO6xrCcorQR5XiV
rfgLBPs4CdLx2gKhofaU4unM2V2HrDMVqIC1JSW+VR84SxSWyI+RmUC+5nP7gCVb
PgOK5Zqi/X79AM7upWInM+W0Ut1KShG3wMb+C+VIECaL9J4CbDnlUHWIC0K0Utzm
3FV1BwaBBrsvGX7H2hL3ZKZfErVRDLjYF1QqMaquOdyqgrg2Rf0uOBRWnpAt0rC8
Gbr6dZBNVqnbxOfVh9olMBbf/addLSR6hsqmnfrdgeeEIbd+A3oBOHco0cZs0EU4
IV/n+vojITYrlMVHb4VfO3viPkynRJis+ZipfaHwDGsKwZJxQaLcWy332ZUm/23i
5ML6mmdcW4m7K7QHNNjr0TSeGEdnMAxhnLnvhWUyxUomJEXkZslqTzGj2c/tlcal
xHudd7NkBu1lmLUwVZowjN0RUcMBX9/UX+hiV3WWIAEdWsTjritng9rUUTbmlErG
+CMjqb2DEKLZ40i9aI+1buz9mEgugAcCmWlczyF7bW8wmDMpowa3joqPgpxtapJS
q9P8WTiIbBpHMiE0rMDg+YMNZmT4JdKn0cAFt/rluixe9+enEvqBe/1woqJ7TAn6
8gUJglvLJCKk8F7tcr/mbq2j2aN8KGBFphq82XxG/ygmXW7/l6jenBf8dzzELmqK
9UNFoRqIeNTd5uCVUvOq1j3lFO0yFcdAmRbVLUq9weHDmE7IfgBr4qluJ2ZhxcAS
IQUy+hKL5RINoSnhdXfbNLphms0clvGem6H2Wp9KBIrDMew0FGiqXzE2bvRXf82X
tLsaK5q+ziZGZ2FQf80ytBuwvWXToRZL8ah7ofwuQtSG0j16UkypEHdN1dZb0+a4
+flRYUOvdijOk3PSSoA7UuQqBDHtqJ5jlWcPTvwlj0SQbMP9abJ6OF/cdn/1U5o+
I0lAaF/SgQCUfibPMHZg+4ulpVhcBInFUGI+hDjLHdi+t0qYutFLYaCVYghmvZ/b
IjpRSYmEdYLFMuDZzWb2l+ZEmDa3n16YdMyfoncdXAXWcj6KoUKq9e7vRE1oDF+C
5XKqhyvUaRnOp1gvYIUuWMRx+OKR7/509GkH+5NNIjCWmRCkXuXOlWbuYkh2tW6D
4G3Z3TsorcKc5vaniYB+gnWfFNou9oSoLnwJrUGZEp1OMJHs1qboWe0EKI7gnSAY
IDjhAiChjISWaFVHOm9DPIF7JRARZfliA6vxULUER5waqmW9j2gyt8S+XtBS18do
vp/6kgV4oOeH7rtWtFTm/3zldPObb2Uj0/oVbPhjNLo6H/2j1wPDfCDaeBze1ie5
lmQp/FNM35LlpHntofQBrn8gIt9uxAatVhX5ZDAYmXflF74OlByT/S34MgftXyTK
NqyfQmdpMVCAXVGSa4uDyiDAJmDxh9G/oLTY2xCjqQx5QKHPIzsKiF3novjUtRjv
WaDp8sedHTAL79yea2PiVW5ltk5PMdUtHwHBwgT8CbELLDYdJJHswWrLCRSk3Ph+
73CCKU+UFbIgtrXXoMpLJODa6zTxdbix9b3GLn6UzH3w+WNoOzF3ytbdalD5OMkk
/Au1mjWxXBU/7SvzcabwJdn0RblFdyBF3cE5RvCr5JoJ0uHIBlKBna95VIZ2xi+O
f06Q7yup/yVKhhAOe8p88kq80HPu/XB5BUMurnp0Ry5f/zATe7+K1HB0MKubJ5jJ
gsKw//qKt2LsB70ZbB9PrhqlejPPzbwK9YW/e/y864tddxubbnoaawpXoj9aXl/H
ARdCfmaWo2Cp7o8eUVK3428F73aOkejvKz3MNXhCYh4xCJBXlmBYGpH3FEEJsC1y
KEF/vj2s6RQowh+zoaE4fBi9zhFgv9TBA4iwaySGZ9awxcdsIzfj7m9LEuOVMzUX
6bpcY1RyEVNZwiwAMP1ZKnOA8bCEgH7GznGRzyfcoBv5ILskbraEH9DbB1jeQu+g
hOHiDQotQVypkBj8B++jnkrOTTPB13T6RFQR/lByUU5RSRhmSoAlZq2Jhs5IhWQK
DrPJme2kSEWQ1iJs/jHSraM706cxXnSIzGzbn1AL3ogjO8Yk41zIDQyGj7v8bOew
Ql/bbMkkM7pLX9kQN0v21q46IGNgub/8nwP/Ji1ToTu8HU842DK1pZ8ElAdD1D1+
+BL2w/QL+IuAjJ1bZPzhS01FddwFvUtP39SBi0xnt4xc8TLnPvc2eN1jJ/biHqZD
48Z1Rsq00j/oSJAQzO1uH9M5QnrwrSiuw5hzfZMHjWhHukIAYZX+lgvLIZY2gvye
KNhc/HjW7BnoteDGZmWLI5Q+pvP7UAfcQ3QuUxmzh/pDzUbsDgZGQuulPhD9EURK
3Ll6uI+dxV1q83ZbY4vev7hD3dfPjHYZ+UAovlLM13CBisPKxy6SXVpDDniEMaC/
KmAW6HL4EVe3h6JSj3O7dkO7EGReuTM1xydsJBraMQAXQaGVFCeppuHM+vj0JhYK
hd5LPWCI78eJCTl7Gm7wZw4S+8PsG2319c1eZJZNfMAxxRc02Tm+ASZQhcF0RlGB
c8fdbfJeU8dLQ0S6d6KbtMRNbayxWhaRYmhfPt5LFt/4LrXFDap7nZgUuUTu4MII
ElbgTtXCuDdFgEb3kpYRUY/02brQs8HUCZnVrnIbmkx5/yOJm81o/HLiR+8C7qGy
0lX90YDf6w3EEQxm0PcUo3qClVVXJdfmXZuhULWztJNYnK8Z0ZF0EZFvK6a/2qPM
DZcu+JhniZ644wdHP83jA+XAIpk+FFDD2/AF+kkS3VZLSMfZM1iLwVYyuJxSsyxP
nTF7VbMuJfdayBPonPrUvMDuAUfhTXmWojkvp6FLRMBaQri2qFqX/OjluIcux956
YSmrc5pYmzZpNVgR7C71NUsliXPSiltD3x9nYAEFEJrPla827INJMjQxRtohafdy
9yA9S5pW2td5PpafgrIynTZdekR/S8ria8PAuSolCKj2klQarrPdQW9Y3i8bnH2t
KHA35EprASEorVx5S6G8UQFOdNy+tbsnY0KOqtkIxjjH/2IkUFO1PvMlcKXPMZ9Q
VdUciM/8F9ElQnjY+z6fV3UNncWA4fy0A6IOVgk9IdqqGc9oaJ7rZVHLaKzl9phZ
cR4emInyqBBDKixAeHNWQIycKYfDR6KNl9oJp7mq8w/5VyKnq8KQESCsBl4zPl2E
h2tLdrwD/7evXSZIexBpHMIUMnDjz2Uy4SQnEi5I0iS9ev/+H14n13l9AKJmDsZh
Q7Upt41sqIoHjsFFJCeYPG2QE6wi7r+DUMEPfx+PKy94NIFuCUBa3oBl1lqcBbAj
zmG19s/csXkA/3W7uckkK4d5laI+S9PzXO65A9PfdTlBBrxQlZgQXuddczCfbnBC
dQgsgaa67d1TbWQwBagPbWE1zugacghTEddRI16xSlDFNEO7ZvFNjI0yCAaBm8xQ
sk3vl3lACApkwPvQgZzIQkmAQC58yd7rxtzc9wdeHNntHSkh69m4ibpr3C3qGOgt
xkM+M+YCSjjfU3IF71EuApdkHapMlXap4G3uSmkMePtauaOdClH0GTofKuRoO4mU
p4XmBnI8/BerNEdu2lBHmdAC3P317sFVNaN1EC6ed4ARBb8Qxl30BCtOJo8zyFev
1JWMrVr97hIMbi3D84JhSINcV12GnbXKHcrlmEm1tJ3nOjXMDZS8rLgdsGH2W7jJ
DUuKxFk/wJHr/OBnH2PZRh2rKwUsiw6R8cebZb4Y+AoJ9FD/c5CTmajGP0RuLWm4
HITpS0q0yqplYCxor/PBmVxJ82sHgaPHHqkElIzG/pkQkWCswwEk8lWDzHi0t6b7
5ZD7+DM2l26FWQzc/h3012VDTksTXvXaXXb0eFNXR+mrPszhSqA0BpEhLEmPU1Gk
kHSA6QB8FyseKTHWq/NSaZi+rFOh6gV3vz/3Yfb8sGxJL8JyZIRFfdv0YDCGA26E
OuGjOToBo0AMMLP8UL7fl+onoUy4G0nn0eM6nvG3c3+HW/yOXmXNQXmBeqsRiOrz
5jmrWN5PXGInxi4bvIODPccLRdakEkucJHAAFLBqhYMJmgjKmwa9wOb5oRJqRCNa
tNU0t9AooRX9NNn5ti7t2tfhcBFYMSOEk3hzFN4wt6SWN6p90skI/FWef9kBw7wT
PcVvdLnTv6iG880klvXEuxXPejym9uG+JJVQmypcl8GlgQC6P6dcR/q2sDTDBdnf
Qj1dxsIc4mUzsl0rQ2DdyZLg4dqbcCaLXqSJB4LOlQqKCquTRVJGDmyuubfBxuVO
dzZo2IPEEouam+rYkY2xLsiDjHpiI+VuoB91KnJTvYmgrux+KpxrqdEIj+kWOt5h
R5K6n9hKk+zOJTtZPkj6JD2pRlFJavSpJ9sAqkUUtStN/trAFHzyb6c0ai5pzx/r
sKZ4GdXit5TrLRXReBmzxDxGSjMULRCYIfEcK/KQyH83dKxhaDhnIjOcuaA7ROUz
rZq82Y/OxLAys/EvNoZ3VbPGniAwByw3RntjSQmu5+Nm35YfTv0tiZoqe7vcFQ4c
eNDeWNbhdCvR4S2jLiJjH6SjE/dGXKfd8DY3ahzuTFS2b1sgkyrG3A9xMIb4C321
hRucJnGWfvTfqKnb/6v0/8+//cV3ktbn/E45sPp3I8cUZLDzQacBwefevrJPhss+
25tfYgWQ4VmbOrS/N9f+uccGsg3arSCSDjnZcCtyVjmlyE9DV8PejrHX8PfUT2FH
wGVI5dtPMmurEr7Y+xOP3jRAQB5PaBe1y+UnnZtK9S7n5fnyP7oKJOgSVc67I1+s
72Ogt3wbbgPsnh1lYf1c4UezYiJZw7UYDgFR1cMMdky30Yto4fnQnPhRnLtvvse0
gfjxwdXrhy4aP8qY4DR0EIovdOQSNnM2+zztIYpypm2EKXwhE1/oLn82UJaIPXHi
6e5UwavXbIMPb89mVR1Dicsy3ywLWA6LFiCO13zAONy6fG3y4NwrODDDWPfqrV47
8miJoWh297s6zIFm6ZWobXZukve7vmFKpYgN2m0j6z1/FHtmkfZw5UUTEoSVDMCN
kNbnctGeL7HQtsXXVEovrZiRPl/3xX+/P6ywX/bPLb0DHppsM24fIQdDqBauWrzh
GE920d/EFLWttZANCT9Gwkbuol/8IjFCjq0bQbdYC7AE6ofoW0sNiec/ytB9GzO1
UUqfCXe7ARW6xYB1QDQE+ZS5z4Phb/X/QH+F9B0tNgLcLwdrBhv3lEiDyi1S6xxB
5Wz5Ju47Lu9yKKW0oHLByPYg85boEfjqzvTGdgVuxHV85jdfCuQKa2EatBr84ss3
gAcerx0YqRqhD8UftHd0CC58PQjDxfLOWZGi6Zovr/SGC6MmqD1gnJDXNERv/K1M
Jf3qLMmntIsW2+CFKDQRauJrHinQy3jmp/DC4Gew0cEsDu+zz0PWQPh7He+4M+9y
iQPVuzrcxAfVxjfOlu0Ic2pypqO8TjCcWG53xzjx5ND2y32pdEqFSOQat8ARQuJY
1WyKEdTfXS3zu7WLGNhMoSVVzxWnNLCaFTTZ4kHn0o1OqQB10/UX+z1NVt1fUhcf
jCA8MmUp6EQT7p56ZKA8qj6NK+I+r19GwQPvcE5N7Gzou9/msXdp0gX3P4rHFsBH
BECkNzcbVnn8FaEsEGP4blA3Bzw2Ddw/h5YLSHxjplZ/Y1NLFSrMpnvNwsapA8Gp
mVfX15DjjMk7AfWKBq6eR/oxUXY6+y83YYAioRmOXSIZA9DcdyItRSNKon/K4Ao5
ZvM28xysV/Oz9lCkn4qpUyryFh11kx4PZkViKFC21jGT32oE6LTnc0kDhdTTidCe
5QbD/dAJT8QLO5cWxRiElhki//u39GODobnBpWjkExeybrVa5PHuuZ5Hfvvhnlqv
67RIwtRPSV6/MHQS9hS/6lm/ziY0AXYW/xRVAIk56m+FFdv8bwKnxZN8os26QmtL
3X0RrQfW/5MxEXu880CAvFaiebyJdDxACI4oMVOsnZfAuKdn76RjzEvVp8uduCu8
rnmTcm/LIcZO21oGbNge1Y4K4syj9SrHmpE7iJFjWYrnAmExkiIY82PMUcjpxGKd
e3rlWLEiv5XtyCAl1Z6aiyuMjSPTfAnBbNIhRh1oFiYuABOo7joDKNtREhu3nMH9
b2cKvlLzb8TiBO7VyErRzmA6vN+gk0QrqrpTEiRDori6Z5hGAhASf/X9W0pMomRy
i/iMruC/QMCwvDG/DhMYcmnJsves3UIwpt4C+zSyacPgdHehkFKdOIQaA+csKOQo
9pBCrXWbK8tzclsRrETHMaFum01rhCcFYeqcNEBpEMHILMq/A8fcl3w3a2V3V76F
5WZq9dhPnJRw//LX1O2cHvzcnHYgsnT4Y1cUoc6QXFspbnY4dwMncjzs/cwl0w7U
FFjxR+E/JHike6TIpqm/6P7uCfcuxvnLnteoIYcPYlM2iR37nTqMbcnXpA+YnvT3
29P4l5sGSCBn3SZHH+qJ/arGPvlKkq6pWHZFnO1+GAZeT8Vd8JXRKTHfntw11MXh
Zs2zP4+32RpEI4Z4xyeANvqiVsLviS9BDKA2LZM5ybQ1caWFNs4NQw8O+M8KQcJj
BHHU0YM+O0Y8H/GUzH2UpntQV7IcvG4KX8qVaOqcKhTQWGVtv+Ip5m6FGLDg/36r
fodsWIlfqvxC7CzYKy7UQH8xC86O59D42jB9I29tsRwdNuxwpamgJujXishtbJDZ
IrtaVvAKw12/dc2kCgWpPpEkg7oS0/hhZPAvmgV1Hddl7FlMS2G5Rne+J02talMl
VuG98iegQ/qhj0zVJ8NYaIAAJtwq2gEfB8/eZXGQMmlRCt7Fd9eMH3V5zzsFfrCp
Ffg9mYKPFBOgERc2pxdptp6NA+O9I0P/Ul8ouXqeeMvTMOYm+5L+/cOKEvVlFP+u
Bp+FC9GJ2gESjJa8tFWbApU+QBpzegK1MZmzZpxX5O6J2q2FPfqzdZRndmkgRecm
GPC0TgCt1wwf6QcI7TNc/J6xFoSAfFoRB3O2avfhzydVE4ExRJihHwNDpzqXeb/E
7BAu/o/wvV1UJVIFbTHW6UvkpokH/FgGSMOOJjB2x/sKI9zKWpsEWcHxB/3T3b3s
TfCalIkXbhuJWIXvT91egx3da5guZwWyjA99BJmIVeA4x4odKEkvLjv1JrOMt2xo
KL/nEm3TRjamEoqp955+r5dFN0G23dYSwXd9Cz2+CSMu9FDafDTArrGeM1RSC6BR
V/jx9uA+yVSTkAYIESc98CGcecDZNsT6G+TWTMJUkW49kcb7sEFz2ybOnpQX7pnE
McuzCshY9E8c/vBeFK9WNB1Ym6iRncDIMYkKqt/yPrERzQXGgXf5Sw29/3mzh1Sh
89scVLU6fKVJeVt647v5A2Ggb2JzHtcerGTao7PPQuJRnU5A2TldWiEa2Mmr6WLn
K+HufqQfjkw457eFrLc+gqFXwOF/xbZCrSHP0qDFIUt2yOIaZ6SE/6JvgWa+cFvb
POL5g8suYnHPmhrP/Ovgavi/1v8WjRDdMbgv6cSdbcXfOSiQBFBiXu2pjCfHagRX
GfmVWfnO8arR0RcwD4YByaW4p6Z26vvy8NDGviNMjAKJpXiJMGskKaSRtCTN75Rn
5yawMMP/gpfbklH9+cRHGyxPljzbraFA/XqRi4HRAjhUj8y/ZsUhqfHJGnVCdC+U
bsC7bAr9npgJ0MmMOrQwpcO1WQTAnPwqMi8ZrIkdjD3w8Cq5hNkkCyG99tht9cHR
+SaYpQadusE4jpXb5noGWlhNOymfnzVPl825CKX9ZQ6MqJhGJgPYJMYupOigMcUh
jHuK3irSwszc/ryJd2tfdsbhIBsJOcUE5we6Zq7zl8lO0u7APoB6gaBNfWiIrgpr
t59rApjVxkcmk+ZpaAV9PE/nn/sc8+VPi70cu1qZFXynNJaTbp5II8wSWp2I6n1/
8MR04BU3hhbPgm873mZW15VH3yYwA1ruXl96zL6oaefJUe49T9uq3yTi98z4+5yx
b+rStpLXcrpTURg9bS+M6eyjzLhwf9vzHfggLzXn8vCRlLEEVIG0m4kiL4xosmRW
XIw2QydpPCkKG0Ur75EfnnmIX1hDI6FyDkcYAPfw/gB6CbLsq+eAT/lNp2P00K3g
zIVsonbfMKVlpnf4iKv2CjiLUvs6id4QFHS3rGKlARXCOs8GdG48Vp0KhZUoKaRI
DHM+1SZJ/m0KnfhKlnCw2MT1A2Zq+6Rrg7napv1Gye22Ovqvtil3dpvAVPKz+3tf
MbOeFnGgJWQLnZRyG3Cby/Zr+459FWvcNRlgtTH+HChAjh2zRBXXEGc/kz1DRnOE
0t9xf84ZEheq6nUA751f+iMa4gxjqcA5CxQHkY6dlyritvgHFINZiMUQJz0z3kZU
Zv48jeI1EoVqSO4fLTWCoLsILBNm+7fBUJ9uaMrHS6SiZlAXwLGdaZv1YKssXtfa
pY8kVu8lQyH6O1wu/OFXIrJTrqbZjqD0wwj/lD51dxxXQT0T35Duibrjy1cYrF7k
oVkri+nvCzLm//xB3kOBMO2CZYivDbqosDAVJM6A0ZnsD7jtlX413IPnXc1d90nG
8BRNW+dsXyrAc7cPFDw9m5hpBlUf0IGVAqns9znYCVESJmKxs2Qr8at2/P/+wH4+
iOmd14Ii97PPbbwxp2vkzBDXQZlGD9SwbYmEqYbBNMoP0MLbZK9+fgeTOoelM6Sd
qzzNKWkS7jyfqvtMnGU0J+vGR+gW+SRIYNROPu3H+icqsw/kHK/xHFtNsLAI/Vkj
JL5M6TRHQh/C+Z3FpmEDVXeWbave9s/bge2h0bVMx6H0udSyK8r87jTL6S0cF27V
FLXzu/BVMy+9LJumUru1DjI7rG4FHo46/fW9p+UIay6GBuAalfSu6YMUSJJkXqtt
VYzML7LBLVwLxv9QU4OKlpyxuL7QnKpMFJfyUhY3BTO2t9lrafvnBwt0BNV8Clpa
SvNs6w8ymqfPxu8mZhT7+QJQB2wJoATIjupJxEVegwPCMXbG+d5ErVmtFZH3ytfS
cx5qyq8Dkad/TVXvD1o0R5T29Oxp1Yx4343EBBuWedGuCz9xY/X+f8NMXYOadK8p
5A6HmTHZSRDM+y6fdQBVFG5C3EQh1GrgXwxprc9XgSCoG1tYHl11k74p6dNlGJkv
E42mRx0bsuWYS7YDnV7mce8dGdjK2c9iakMNsoYSLy6WsfEVE0SQG1wwkIUhx1b/
X359BxnfNgsuQwIwR0nvswmuf6NmI7AMi2F+sCtvFvd4Ytkq3f9++OtllKxJQsxA
6zMOkyiljTRJ1YFVt3GEHVsLMos1RUS3P7N0bSUlRA7OEsV68kbotGy4CCs/diDK
oxmfBcR9JEJ4mzdgmOLS5aY4AMUNE3IXTZC1a14qe4DwuTKCniqSUY/m/1W2klD6
l8UcYYzRZzSkTke7ProgaJuFD/ojBiX7TQWY8nkSHtAuyU5hkRQWemH0Ck0EDZtt
zusfphq5ciyS94xQLh5KYPcPQ6Xx6cqHf0Vc/4rQNAKbvu/E3VMVtMAaTubNLl/n
jf7T4F8TPPkxDGmJvYvE7dxjBYwKOqu3NGUZ+7sdCW4xotNDEBh0jfVCb3cgoWLQ
tq5RqRfz9hbgthhaCcLyEtCGxYNAqTbsJct4uevAfL9VegKxFsOPl2tOGST/eeRs
ZL8sNsXsk5+nHLO3gyqmvY7897U5EtYifLtNNJXLuoPpbWXWuEDSfwr+TV7HeyYf
RXo4LGuANYScTG6XyCblxG6MyneyfO+9UitdAW9KeUeUm68coapzsJkQwNydBplO
VenlVjqnRfr9IDCFQwPcQySfwGqXPtIAb+SQEFwxsAmZfsykKPKTiZhIAdc4WvrT
nfO5wDgmXqW3kJxvLgH6b5rrtudMwXZId19BCYe5ywsVY3MmyZ3x2jROS5dRqfkR
ind5S2y4J9c+F4lkPUosfhWxlJJxZYIoLoBh54l1Af2A3v6OkjiB7l05JW4LCVku
vr+f0xemozxkTgNaCabZ8qExezjTDuU8eZQcwMUFdH7Br0kSaxb0RlH6Ia+qFedx
lOhZ3mL+yNaMj8S0ZC7RnJsAEPKtkIHm5z8L7vizitvYJPhh0E4OA3EqdR1wOvGd
3yVnnCWhfldPcfofexftM0iiG49/9v0oxZnoMAgPzQpnqwzuT+eVhxSRttESJFUR
SNSXTBhXUJl7N3ELVvOk31obZfPAgLnWAMZrpBBPlAE8K1Qge71lh29LlEvJhR1C
xd17dVXlc5I0LeMe65gxYBDGRi5eTb8EafB/eeLQT3yq+poJA04TwutIuLl3NhkB
h85hovTzC2Vu9XDxIFPbh81WfGL6C19EZRfsmoQwcymjOLuuHANWYhsUHqTaQAyn
DKQ0uRD5SVkrHx9RLTNZnJuqAZppbs7Tll+zHtJB6tsGQadFz2jhnRaAH2HzGctN
vSiaw8jGtRodnHtUP2YW9yRTnnA1ryPjEcapJ4FPAyhwGNgba3Fo7lL4C071tEDc
hvuxSquOO4Mf6+DEI+mH5QoJYlZ5eiH8KafuNs+9cIDvu0noqt2v7HWjzREMX8YF
tOg7J2xEKqDzJCjq0n8/WPqC7QU9tZ5fX6fxuIiFxMcr45SvV4IPpHnQ2F1X9Oc+
fBiKM9YtP3asqjSDAvGT4jQk/CYGBN/7Twrcp0tbW/RjcVn/TzVEt94o2X8jMSHl
5NPnth1+1HteyDoersKCOYh+Ej32Kkl5m40mexmdYu4XB813uTbAykG7STZdxzQe
IqUMgTiAoIhWX4QT0zMM/2xOA4Ke8MXOFKI6I2VC6jSmE518D4tPbXb2x2Bx+oF2
aJJ1EapjK5miMkjKn6PjgEra7tyvWP/rHfN5HYD7n/Bmsrs3IVf9TUZyBSzEL7uA
jItymw9suQzdCsk9F7fjV5ZvDZycQxeOh99f52Q7qzfhkLP1089oV0gCcw8nsiTz
blSXqLIHfG9w2uJjT9fAE1EUKoh7pZD1PfI4BCyQGmz0cUn0PYEhpNutjWci//wD
1ayCSnzLA1Gtrcam4Hdmu9QWqNxqp3Ap7QJtX/W+siPaZ90egtxhkRMcfBPKU2QC
JPuvIn4iVRq3ic5O5WTSh787aTDccYsfQLo9WmqU4BiD0Isv68MzMdoPxDD/G81U
fF7a400DSFSX+wwaNq+3JotuqLcAi2I/0hq47xlJTB8nXnUi5SANzA8WEtHgXFBR
CMKzCbp/ENqgatZtoR2uX49G9KT+IgGWzvkQxhQdqyh7w42cweSyz1LXr5eM5cJD
VKvPG8GbHuqqjumu0WRlZPa7vF9OGtAye8EI8BH5PMc8szoCxeE2oHxBi38Uy0H6
Rou1VCq2LFkCe+lMET6dVX0hVBE2kwEd53xppSvp/qAogWpGJ8p8cyt/baBUiewd
63Fgv3WKqRQwsHC7MTRRkEkhMG/yv283Gox9k3RvNwIKnoQrnZm/ZMh5kUR7UxvQ
7BvU01SZZ1MRpt8zqKa9whJdOTHSFsDCn3a6tZQQqJAbH5MdoEOuklRdTsyqh3Dn
griUT1QOrMwAzHPNFyvrpxLTnIr898paVrStpUJ4eij4ehqVNtcH3qq85VhJewzk
2FczjD+EBA9uhqY5QbOSaen3l8od/8uOX08WsQnU2W+e5cNEk5OVeEdvTR8mRi25
swajuLTZLO94HL5YcptktlYGn8u3+v34PSYVB0p+hNIiVJzU+FsXvD8hWy7HHzOi
du9Rppc0fUJphY/RyTh//qHBxHVUEFQYnGNO4ga4dut6MBgDBFKW1mbrBxs8rk3b
sGGFV20xCNTxX16RWi8ca4FWpw1AQ2bj7ZmS+N5rITjTctLMWS7DbuGINePP5sMa
SYrVd0ZE0Ylh0PMdIyi+F9pzhn53aAjX2a/bYhS6O64QeGHqSu9onJPYCivZBlcm
qt7t6hXwQtlUqVkamhKZRm1QUds7KDL8KJCwrkh6522hHTuUiO8/wSkIlkgvfaGW
XT40ESW6qEOFvkvTci9ZbMkMsReld0msGBa9oSIWA3IfQB0b3i6MWIWG+dykXjQ0
PLCuE31y7D/SiVpnOdeZn198+MRsS7TNJqDBvgdBIumVlptRYkEKoQYz7l6rEMjy
EkDgfYIx7f0+3+vGpetEnO+QDI5yJYjHZZwfZNfefdrGcdlpxxTDugPstfpYtoUz
UpIoZjsJJjDVRXJo8K9eJT6NGOZDehCKtwKqNPtp8bhCHSioLus8UmUDNQTzHWsq
u1761VvlK65rWHm1utMBhR50VIk0j7CfmK6b6qLbvMPLPMmMrOJPnKGJkTwAzvtL
xoiAc4XXWGM3N2XGtdSudUl4jaX22lAa7Su3rcMubhP3e0EM3kwshxZSPEQkZCEK
TJpf9c5YB2r4nWKDnB8HD1R+KKJFaCDLYbu2smEIrkLTwikgQ6hBof0jO6mH37V/
0ua3bovBmQ9kZr/bIFa5Mb0rYWjX50FwRI/opanXV+C7UeJat5PQA6eQvLuJ4b65
NtLIL9odjQZGugMWBpuAi4DsQ3WkhR3016UGvrToXKlKfFctIYs0dEVbBH1xKnzR
JA7uFcvnWELiJvFEvLtiK42nknuYl4ye4dLGM6kGXV6JIEV0NfwTRzqvrorgwxwD
XLhj2pfNqOr+UrLFI2bJhe1bE8b//GBFSmnF88bRpIUOgn738oBb24TkgKNsgyP0
8faRZ5vQWTkNfsVx0TVSWat2ZH40FvP3P5//rfJxrMcTs1oCsihMFPXk83GH2030
DSi6+rAMbdHJJb1JGJOTcqEm/AeW5vY2oh0rFF7/fCQfeuk6QpvwmSQMTt7AKSoN
3TlS5QxSrtUqv9GL84ffJYFgkmeCdXjhUJpcw0Q2lQkuCvY8rUe4fr5kUb1VUruV
36VGxAYMLz2sDGm9wxngxE7mwJK478t1LBxVdztAX6NFjn6nJ1dP/NTqV+eAZlLm
lm+M9MktGxao8FvpXycVp/FkloTtyG5cnj1dds8TV+UlVZyt31f+R37j/r04I5jt
k420v6E/pP7hVYA1p0yZl+GnYfOkrg0uhVA3QnOcZQt/ASLIQsm0g8uIiJvgP7YD
2E5zWRIX2T2a2uaXQj6pkxy90sZtFXh6yPBIFYm0BBcvpu8a10o0iTWXlOwjfKHh
Sj4q39xiE3sYft2WQYQtVTImOWlfMEg3+DzIBFyg6//6lXSc10XO0/VkCu1HBBvl
6Org/Y6Q1dFbvQs/IydpCu+tL/qRZTNv+ADFavZgJ2okFrlEHiJDtvGKZciqQJ2h
viLcsb89Cr9qKzUreW/FWJrmpdRnJDCHG2BoDEpaSF+tjLAwLQZO2t7Jlp+uBN8f
Go+KAzrlnjGAxtbRwbUsKnsZ/RyORgGtqxdur3DgjyFWWII9bJteJl4zk018wH/J
p0bZTSNd+zWJRTA7rz9LEoWOgZVduNc6jgNca1JKQRk5jingtJI87tdes1qcC7xe
/zFBQsj8hW0EmRm0o2UH3LM5Hsi/jlrVw68zD5bQENoEVPdSgRSYqMIxipDQwGZW
Ny+3H+K0xaGz0fnmdH7vfaO9qH8S/MRt70fs3tPdi7VrI1yEg+rOMPVa3CKu7dTo
ikMIIVI18OGnd4WxX6xUAi0KslDlc++kXrtAj+vXJo9RT9F2xMF8nMnmeSRKQi9J
M+68DmhmAw862Sn4jaDC62nM3wtR6zkjbBao5vkgygWVZ5/E2DovUzk3dSufuXCm
oJId6R4BsamvQxupi/HRubLJOFnowExbHezDVGmRyfK8psCzQfvGYYO2bDghZ9gb
XAKvnASvOTWristy2wWYe75m0mPqZPSPYz8JPqOfYxOkrhXBBBIPm6Lquh+1pAXa
0x2eAb/JkQMEBR/QGn7GSl79QJi3h1lcUmBLRmf4dq6XREGaTbAwQ1I/AAemQv0S
c8xeQd0epkPheHH/X6d27+nH9x30ASYsxURCW4mlgoYJkY2DzvE8FrInESTOuDIF
9Jc6OnLTDYMp0KEuv8vmYzvCN+DiZb7f1ESfpUQdQwisRKczWPot2yMlegwvuMmk
iM193dkw915UH3dN8DHsTLjR05mSjD+Vmi0If8ijjR4ibJovvFJZF4dVzc0vm/5e
BqAQa0VfHsbm58YlFw8GCgsr3JsR4ffqm3RnyrEklvj9uKNuJjTYdE6oYkm1zF+L
pKfH/yzdzlZzFccZu7yoR9AJ13YibUmyWaCzJoDCQhstLNs/ue25fqdd1M2Oql7g
nPl51DZ4FkM30n6O4B/k756tDlGD5XRt90fl/oNoBkjE6/pfvNJKKodhatlW1FYl
ZwNnMIZ/t6j4q70GbRN+M0wDCM9ZQWHZMxXGkHy/b+q7BzVWHAwSBX+XkQcTn4aM
Pq6IOZIl1A8W2D8PKBuJwSvpAWm+88BF2Gz3d1x5GvN+kjfEeMcGkZUvOwTw1+rK
88/OEx8CsBXjFKyiSd/7gba9oGAtdQu/ZXWp2ybVg1maaAz7UsKCRbo0zaqmqdHq
UzxwMOa1hpQtm0FVeJxNis8KJOItxuj0NCCIqxEQzWCwRv8P/dUFGlTKbLOUD2DP
iUuMXCF1iUkqlzqG6pviC5WLtT4dHlnkvvf8lOU4DCXsEhKMft7niFqFwcog9nTW
CnerwMMZtT7rCPRhb0U3nio7pWN+Le8D2YxuCw7Y1G63uU3lagYnPqnULGQNx4IR
nGo1JJEKJH092+C6M7h6mJOkhcJcnHXdvNeU1a0N19b09dTGQF+FfKcCoF8u7w7Y
Slgu/WIlno1PADlYi6GHdnGMji+dQg2Ue5bZaCa7iytDORzNJYSzTAs+98Z4UbR0
W2u5jIBP3fGhy/WILxRskCsmy66Qo1JNvTaZ375X5nEmgjpYEFMnv76mEbBcYIS8
JTCZ1GT23xIFSGYpgFYN9uAOYifAaQXQrFYeKiRyxBeyLL7mx6IDIgsFWRNZh/Nh
p5r0jR1MSQNslzreNCn59q1l9E0wAUBZ1h22RtGYSaERqJMxc0Wd/62OiO54ITkD
RinkDfIO9OFGD+v4fJLz3Gm5e3R2idCZfvZCMwL1zj+CoabBpxxfFXDTATh2rjqf
PAime/JhAt13b4f54wYPp+Te7KNAWI0SIsEGw5x0jM1RxmQ6wxqsc0o46ELfRz0A
ILHQaRXIt8H8GT8mwhhlo7WA6AyBtfZmg8/wZddslo6yxG+JCNXHkGh/eGFeCKGg
E29ptWDSfGtJIC1do4nK6/q+3AFcHFvADj+s3KK+6wMNgPxiFToYnt1bicSr4gI9
TDYLjmeg6hGnPaBx/XcOin4RqdF6kZQ5GFnJcn2YQGE7uYu/NT1W3VCJSNIdPWR8
PPRM27+4r21YzaylaxOpBZPlo1AkdsX+u8q4U+Zl1J10WpvEjHwi5GvPSmju/kk5
6/8mEbRa0A7U20H5v9m1Fe+zkDqKmm5QpISzv2YxJp3EXFbaeCdmDWSUedD03FXz
EhHqtNmw5+qDxk2m/63oOwbTiLuNFynb9RG4JVTQKXoSYWxstrp65QCHaqDMPm5d
qqi4FQkOvintUvdflnd5+NQeIjJA5DuoBfFPS2gULoJry4mPghsSqq2olTxRSl+S
TUJqy41W/6ek//i0fqocSyvhKMh9u71UVFp2+a1kI7Q9rWq5DQf0Bq1s7IgOp/1h
3vxb6OHmU/tDgr3TWSMbwadktF0MKeYyrRmmqP3FwynEm0jr2C5FX5Kyw7vz1bME
s/yEb4XLHLvplUrf84WhmmL+tnot7ycMie4Mq0DfzH1eJ95qdB/Mp2FznZtz4+H+
FssU/gGmt/uCGUlDdV79w42wxb5G1L4OyFF9wysak+44lACR4bna/LD/JPk5A27I
I+YZmmLEDa50iYb7Hb5xZRlxQZ6la9f6fZBlbt6r8390WD2l1LtA/EQU7szxQKq7
HBkcMHy11CgBKgHWoiI0gOFMz59Rqyi7EjWz/cfNDauynsrCH01d0NYnA3KibK82
rRBwjuELm67yzrkW5lhNbUxaVg6qtkr2FvozI+mTtPzF8eQYfCA9qZw5UP/ozn9F
wq5t4L3AIRI+P6g6UJ/Nj8uMdEtke3TDcskSAy4j54HB5eJmO6Oww+gYCaNbXE1z
IXE1VU6LhOLDW8//KRzxRzU5Pkxyg7g7VfbGm8gskIv3z6REGaCoVQLYVK/wg0Bh
oo0Q0nr4OOXH3lCqv+QO5c0qDXMQv3Nnr4sdHrWrtVjGxu1I2ktLLPeg6zrY4A94
6hX7o4bKcuD+wOVabIzUiNh3XGhE2XJvDEsIwkWupGLJeQZ04uy3pmVmUeIptFz5
wIpVrQBg2FrHNPwzxxQgJIoXECLlZlBZzoNcLOT9Y9zFGj1mixCRy4f7KmCLRaZS
ANzv9dDSKNRnfIPSbSlvokpY3j/MK1fJeAE0KYB9RTdknc9k7fcgas9qY6mSfWPq
C75RzSNzrvqaecLPramIMie0I40ul+U2iBhm3SisFaoUzlGqaRmwrPCXSkY6+q7i
bSe6aW60d709xdjnQcSDJK9bzPFwEoE5k3PbxuvY0v80FYpE16iWQmA+FHOHOr+C
Wn5fSioIy3M2BEmtBIFYqzSUREFo9jc31smV8BxFwUnsdsCTt5CPXGQO9CbfxEuP
5r/8gFI2t5bENtR8AK06pLgPDAFg9n5mEq9H9zjfsaKKDSnevvpMo4R95aXv9s6n
m5OGAmcU27RBBEajrXUYHY3uvGWPu4GYNVlKqyNU29tlrlNmpx5nWSn98pRtPZeJ
cP/+VelicqTfuTNyzeGWsQpXifBZn647/zaKdwt8OFqW3ga5CiDPsIMBKvE1eATs
MOSKqAPj8Fz5evYwoG2muXcJLQ/1i5AEIdwcXA9eZBCg0pUYvmA/4Ll8jMHSFy1m
R2qFCZc3GHWyscLXw9JsqxsfNks5QQbz8ZM8NlECLo2VVhWaZYEWgr68udE2W3vt
b0nA33B1050/nZNfNLTP5Brv2hwWTHDfrqWqfuaMOYArMhTrpoEwg8ZiNELtTJS4
pvJQr+/Dl5c91tY7zGpvceNpO6t4Vs5JaRJzRXU6wzeDemzLyfyH+m4+0AACmduJ
50MW1vX8Rkae4+0KJe31D/GFJpmrThsFshMxkdafBM/TqeH3IrxIQCWng2qWZ4Ld
GHhja+NY4q3vuGUUkRkS4AIlx0bVjcnhXCA53PPToFLX1ha7zLIhaVZ3CoT7aagC
sEhDl+C27sVh1eYvsBlIQd9k56usSIBQda2/IMX6q2hCK0DIwZWy5YkQFi7a6ZdR
jFEP3cvPqncDFR5qvLWXoIgXbbl1Qrx0C1u3khyZrV87livBQir/o5VQSq7QEjh1
dhbuKmkdFtgAyknE2/xnOpR+vP3buBEbzzKFeknNF8i4G1/TCfvMICGAAHen+0xZ
oToholx0QZsYocAhnL0m41WeNowcDJ9w2xJyLD381Z7FMZCiU/9YEGwEEja1Lgii
gCb1VMV+djdRHkEugTPkk09EfmCQh+KFEehLfmcUsjCrXOsPCu166BhzjS3ZcuBi
4MgyQ1nVQbEST60LwNWcNXZAE+ECNCY1kvj/YE//aZ7jS66sdG/ALgIQSnbV60QV
chNk9siy5Eg3n3loseYHmvlD/WedrBAyDoQIMP3nz9LmsawoCCCcslC7T5B3BtId
AvLtKJucWVYXknbrznwVavt3tEM1pucnMvgzPa1SXNz6BSa/3z1553kRHiU+vfDD
4LSJaRrsZ+QmnHMPRVP0zJaIklVL14AWkqDY8rR/j5VPlQSJBwpmb6FI3houlWC/
Pkhl9g3KxMF2FUXdVaL0Qqb24nAOhWWtJYf5d5M7RC2UuKQvyj2vcv9vg7Wj2n79
YN4rUWHCofD+ZQ4sfbjZ6ut81GGnTpgVKOAYvYKAix+2NtKGZH8PRzOVKj1cWo2H
A3EmijcGcLPi9C5EcRRsl4uiJDBT910Kbj/6r040k71qbt6TVqjVw9IeHC3YGAAF
mhMRS6vr92lbB0VorJpp/BWJ3gPO9j6k17UM7TOq7IOAa3VCHTKNFiOMmNOY0ciO
FhKSFKh1VWDtHgJeDWITrU46+ft/2D9N6citEaWD93uaHI+W0a4QeN6Xgdr6sG2j
c0Ff2vNMPI/pbIVOAZgLt94atkvbkP++54oeG2ghd4Dibh8huCIfaXWRcwKOESVY
MOoYJ8D5BXtYYGXd+AkA9Q26Y4AqPOh5wPrUDa3wC1Sx53IbXeGgXRW0Cp3J883+
Gnsvac3S7uhiw+PhzMR3TYrttTL85zcZzV/ZJbv54eEmeMxU3A5ZTng8um1GkbOA
AztANCpG/p0vzal/Tw/jnPrHZKA/L6hshFfEniiQa0iazD/by5jIG9qhFQwvIm7K
7Q6L/Wzol+iFi/GUFTCIOhW5lvo6rDgwZB8iCmAxxW1a2sdrmKz6CtT5ximCzjyE
iTcQlkzLTux28DKcDXcXOFpkGnqHkaRMr44uRuo8cRC8BxRX1gvitwIFVRHSyJKf
LJ2DZ8Y0FHUrBbAfGkDcCagGgaSVwlfRGLxd/ZZkr7YF+z8Ea4V9YW07/8EgTeCA
b8A5PYG/dulV3j6OMY0+Fl1WbO49WICcro0ohB7RhMWgRIAIRs7mvLpHzSjoYqUI
7YkwQsvVAhOK33m1cDAjylDBHwvKWYVbtEbKW5ebnP2L0QR6s7vX0lmsYfVqKXiT
AFLt9eTzEZp4K4UJbnd8eAiSGdR6nroP2BwRAsodo0gYZjKV+BH39Gmf0+MgT6tL
lF/yEkQCTIuPvSzjIfIPFGAro8oG+bnkWUg87ZFvjLlUzQ1AZf/k+SwSnhZCtNzM
TIKxMZkCfS/iV7jGywMygIho39y9gDvtbzKiWV7J8O1Y2CyxarDNKM5oiGRaWPXn
mDrvg7r6kaQjK2h5o0agN6AEaP00BsWTMN64V0NMQ4Y8FpGiPT114g4YVUTJvtoU
5nZhQzMiI4Y9QEude+Ieiwm7Xo155uzeSjP09cgv2Ft3gcZdiMCspvvO3BuMsJZc
pjsONHyLK5lkDxmgwR1/q7zaRzdTVRKDxe8sJCJ/lvYGrlv/gfq5NQrwS85+5paV
recJqw63/65iJq5bKJYfKx3tKQwu2eP2GXrOMGhi362vIM6zireXV54V/4R/eS19
XnhvP5NQiDfsp3ossfXRMmst9CNQJisFQ4f7ViSUCTW5lpmiELhwJAhscjhDpBWW
bsrQF9a1JQstvPy0fKcYDcoPDrdHZ2Gw+jEt+xFUovog6t/cioIBvDsQb55J+RKt
gg9fsEoibTaNfnUaZLgS0cCBo/d+E/+Y/3xBBqwpDaBFIR+RZikHy1mJ5ZDr9HY8
Yiuo8J9nWueHASGyqiiLv1ygwO79t3Hwgmae2zUBfxiCmduuQXohTwFudN9k3a+d
qjQjVFd23wQdh7rXZJQqaWRvKabTycDTRiB+CW7GW53KqSCTN6Cm/Z+qY5DwOdOG
XntbSIws793c55o10sNX01yezpvMaIXEHTybBdjV9oKlVdPU/bXeKRWvhqglKe6j
smgE83PD00YL3lx3rrJXqa2/Me7HFIPmvvTRrBAy9Bxsx65Y/5TKEHIcdQ6XVcsF
L1aK61j+PFCrrdefjiRjWZO+MaFmv/cemkMCtKxERoUYiPZicgOJv2tgvlCxNWjK
TsRAONRThE7GdGs8leIaZG1eHB23k8EqfFaKOQgtf3sN+bkT8AbDSTtFN0hXs+gn
VguFOGfKgO87N8gx9YZWuSYC/R264YRHR+WmPfJrmuH4wtYUtjPaltbGGWJ8w3iP
Z50Mvzv47AH8x3UdGYcrnJ3MY2DHQ/PHKPeHscDyskVdbn/q64M+REDYOHfyxC7j
glHfSq1tyivtpgWJjyhWwBpJW98gz9mhoy2pHhynEDYYZc/AaKnxxKm+SAmhjlOU
6aSsX37I43xErG/+HUEYW7gaKza2iYnra+lWOhpEYty0PNBF0OA3AatO/YeleRim
PLpbwrNqShIM2iV0XzjJqC3Ap+DjRnHdr9nar8y5RgAPqyIg6jucu9eNMD2yywF2
ocPzXJM1XBGyxpOsRoZ55m+2zKALiyqRvpP/KU47LjoeQl/SXH4hHTFciSNES5qh
HjDdIpxdaR7bOC/D/RsgKQ3D/aeVmm7EzqQ+2IElCbr4Ta3uWMSvUJbJEmZiR5BU
ctl5fOusHY1kAF9FZkV4rhNmCy/0GI9N8OWhvw9WtZgypGLlGpmSOyuVRZ6QNioa
zLsMc0Abl7p/9F+UMiIOIhxpsOOFa9W4g4YBalQrmLdfhAC/5UUkpj/iDELo5vtO
2CKt/KFBsbQ2bRlTChC6vv3Ceo9CKAqdJTIo8XRJYelgq+hlhh+MFBaM7B06NzUa
uDi/0hz/YGs6TdFMlKOUS3vFAzQL1LyAOR4YxaYttWcyAmzfmKPbHsvwNUdd7Qj+
UrbfKpwiYgqMO/PExhNe/ABIL3k2RhOKy0itPs6oSPsGBsqxZzcO+FEqwQs3YQVb
Ha1g75oCHML5eDLnT84A3KO9UTT0W/AApLFQydeckKSu42yC3ojic0kkSyGJxrb/
79h6lcQF/+mQnqZgpqWUxeBlrPnpR3QjUCXq2jUYzSzNQpgvk772jSzHufN/7fAq
7dYyW4s8C8DjPoDzHI6QIFeWWUUT0/FIlpuRj7OvYzsqi+pC0t1tgu/yN81iyp36
QdaK5B846WzzFFOHqE2uhXK860/rr3lcsdMMcFX8mlnRTx6KPUObkbXtGKnvnax7
FOJoUCauZLY01KyLbuRat5xv6vfr2xX2TwKz6Wema628yEctzFD3BZmZx730vTYp
EAu3uER5TWJLrk9rYdkEdPHsiEe1Q/VCJZ/BmjNZAgm7voCyqJzTGsUhn5Y0pOMO
cLworbx2h/Vgru4Lo3xdWgd/OqZBtMrlY6oD+B4jV0XZENEoPcJb4BJLJwP17spg
M5atBnUUC+/lN7ZOEnFXdjxS3KCdiXJ9ioWIp3Q6g0BPL95Gi/JRIvlMEbS5ticQ
Mjfakbx6Iy2Tw+bDIuo/n4RO0+YLfkY5Ni12O8fwpo6dMUoGhiqz4azrtKm6ohI6
dZcLwGBNt+tnNCnluJ8xKe7P47UHlHasjM3RbBl7vOGG9IjLD5cqBkDdDYq6VKrR
bVPRExRBmq3bXPTtME6ddc8TWwGoFhXbg2QnljUX5tfoDER0ha/I069uF91MkQBA
bYGwF96pKyoUcpLfesxWO+unOWVR6/0TIsw7URmEkfk0FchNvppu3flB42BIif7q
SxZzj4szJp3xg9z46Bu8WbA1Af+3v/toCirxxdVmI4tsAGeba5gbHe+AHRj240zI
ixrg6yyHlQB3gKql2h4L06kLFaxJda8Axcwa4bVHII/OjB5tU2Q9CRM5UEX/WSLD
D4Rjab/+zVvvXmNauq5CgCwufEzMTmblTFu1D/rNeN7kJoT1G4fMoSWoX8BCyxOk
Qr/vnvSxqJeWhE4IUOjPjvKiVeEDm3hHdC0msBiUKDf/xfjwrapwh/ew1a++L6/v
yh2sIZsxZTlqkHBZr7VFkhk7bfq8/MXe1blGPwhgijl52QY5XvKo/Nb/gjRIUW07
PHDfqjMONwWRcu2Ujp1pFzqog9pSpAjbOweH7cr7iUeaH4HmHFZH8bXjkD4Pnj2T
W1sjqq3tLswJSE01QX5d5ShsilslsbU/89JbB8aVrE9fazOUDM+e4HLcE3tgWUTw
T0ru7tMAhlqj0DLNM9asS15UmIiuu/TT0seSCeCRn06EMx5hZoGr4ETHlJvl+/zB
9sy9IV+lpFMrigq6laF05OXcjhNPQenGE+vxWoncBuTeINh0V+awW9mzLwMcYYw8
R9Y4zbKkuL1xJZkoRBUBmGeZLmPMhIF+vNI6l6LMocc1/UfG5GAnvbMhgiIao3ik
lOGxi+5cj7xlYkP4QYg2hi1UrXz/jBaUvVpWhSj7x19AAwK2gpBrH1VutmLLNFrG
OMNl9weNHOwmppoK2yjGL3akaMp5JlJd9G2o912K7b/v9ecuFjEdhONKAnD7I9gk
habim7RjulcnKyal1S6qbO8aRWo+v8Kehb+J9xoTi5ei5rg6mMrYN8yIBzz+0uJv
6Wfh4Ip5yT7Hk/+5UUmAAemVfraIufM2RG3MA5Py6u8zfjgnLCeG6Ww+qBp9uXGu
mQNv7WvZqfMpYI1WpJZr3hgpqBejTdEl+fquJfosGAML0yBwjahhaAEUS6ivQ6so
5fSsluaeqviV0bn6Gg5m9PE6u7UhRs45J++rysL08pUNbPynp56S6nujJg5gADhs
Xs8BCMHWOmO7D0gX6ZAeWsyh1J3o1oPD6TMDjmwJD+NNgmBJdY/1zftoqloygLVR
OHR098rX9aVBnP4Tr2PSwNEqAOtBZv3xn+v19cLTnQdtSZjBwX4ScLonTNYPuOeF
5CX4CcwIuvIKYhagHC+t+pKKIrKiYzuDsKX6VQw9+Kb8ON6shmYHMgz7tlvjSqKm
SbCEEPjjBTsyvBdgxhAIYNoWwZLFeGTjrIOF8xVM/+bXwlRg2QUNfNv3iill1piu
Yp4+0mpPMRdCqNrTSRmEcKIoz+TFpUtJ6LULWWRdp8nzZCAFYjsvyPjDZ5k26hjC
sfiAdjbNZfT5sJWS57G13fvIuFrAwYnaguWT6Mbx/t7o6xIXtL9tQz3oHMKiJ8Xq
729bCwsJXwoSC+pAwc10Aaf17J42AoncegDqyPuEGIwZ/CTvpc39v4fC6KE31AY2
1W6jhYr/+oxgGb48xA2zbADxPfvjqFqyWWnr7oAotGbBPuxm6BUWAifG/w52VGkS
46XcQNK1QOi9AYFqezBjwu4Ckqa1VBxLbp9XWjDAC6TNzXBAHb18Kqace/8Dtfah
cIgrxJIphJzTGSBfdDCLcv695gjVioDnbmCUi+GZDjt5bgADATN7oLuHIwjPiH2i
FPkmkOJHnB+pvewRjaigSHz9vcbRisUl8ZKoGh8KGEAYOR9EsD8+WjQtu3Giiux1
FPy0+1GdtMSCIYVO3Qh9w1i0fZegEY4ff3PcNXQcQ0dhBG5QIpgdZByX75Y6wOG0
NvMDugQ+W+P3Nm1LUqwQtuoQ9SLe3+Iahf+c/q6kqCPOQNGQxHuTFOi8HT94aKkn
oiEMMepVlo/3Q70MSyv6uoQksgPNMuc0/cZVE0NZW9D5DDngz3JpMsE/tBh27MB2
oYOfDZEr2XobpWWP1yyfjZ9JqhdXpjVKENz+E3rdRd3ranCeQpT2/DBkMctGD9vS
qa9/HPD0v9FaqmRtzBOUtTaiWVDyUwipOPo6keiZuL2Ne9b4eIs0r03rSOB+jHrv
2lc7Owc4kBzIbMtuJNHvjgbqjVk+BcrZVObfhGlR9E2kEicYEJTX4wOAe+QWscpu
lNJC+FaPSyasxQHYMrHitfieKy1cAbBGqABSWoCL2XuFCj8V8rjRks6+ncSJHnyb
rtxayHJVk6z1wxpuqVWh4WKibscx6uxTEX812bYUKng8ahV280FKxjOjkdBmvcSQ
+yv4xuKSmtyv2vtNucrXFIg+MNGHUTSaeO65Vc1V1K1fIKK3NIiPo8KL5V9YREON
a9F+dBX3E+qAJZMw94BZbGAMXpMvtyZ4ePWnWKA52ezOm31MFrHpMFum5vV6TyXn
cGV0iX+qZlSn0FVKvwH37l1SuKEvIZHhhscdAQ45mK769RcwLZUcVrVcLzSedRJq
tYXTQRd45hwW9LcEMZYfX9LSlHNnoJjopNT0gWpK+XTux+IrI1JN13fURVMBvmEX
/yGV7PxqfCRZcAD0f2utGsvV9F+R55xVIy5/tAvT4fKks5F0P6/lExziZCoyHje9
fw7eIkWDJ3IO2z6KPLmcsXrHC20Mn6upEjxy7SRMF6TMOImi4E1G+STJHdRIkTIH
pj5yg5pUvsFwE8KGBJuUfLddApLPTW6uxPUBhOsr1wGavyTvVFEbynkWwvEhvrTT
fI5uQxrenzt6OWoFPPHqZodAtcMA90HcZKW2N0rPputqu73WwHO+MR0d7pcEUR3T
LRbEkG+Uhnc2GYQIJAxxqSzfpOkCmB6d94mQO4l4fCqjP5nHo5LUR45WljCVYw45
woMy8ACffRh3HmvK0iInNN1gIy9LoH+c8jweQD1Ag1Z68L8085P2ubDxaCH+N2x6
TQAwGPprzBRv8Iw/RfHRJd7Lh2qDLqqKjlUJcOOYg0Cfoz0pdOIpc6Ucmf24h154
iTo41Wodu1riQGduCTKjVcc5Jk/B1NfE+tlZHMXNmJ/p51TAjZn3yPSNiWUYJm4W
I+pEnQOzZTlm68PRwRGXY03K6VwTzw5QJaahiFPNxN1P0BxNYWyk7ytpa9nqGxK4
7lLH/Bk3LE5MNwKOhKw8vVkJQpw4fq6tmGNTcy/08G/cZ9D9NK4Nog27ug2KyJvz
/Mid/O62YTLbf9CL4TRE06Pv0huzTojBp3L03d6W2brtQu6xoDGeE4Da7aaO1iu/
cLdEnzfMLlLabHqQdAJUhiuDy8ARD+Nd11dFziPh38++4SOv3redNDZhOnEbfOzz
oCfnbCkzgBY+8jBIemq5QnqsYpSYrcyk5zX1JiJgk19L9vqK7bJc+dBTh5u6FAMB
VSXBzBVP7lJNPYjqaj0tCNLDU98BCAI2lTpA/N2xXd2hK1aa/7T4KZIulVxli0DN
5d1IBtHOk+/mkyKeDN9uFeGtbmjN5LT38ziwkcSvdz2jiL9e92sAkTnyeLDaoEw1
o4oWQSdVwhlhSikDcduiS41lAo/0wEqGBlGGfjJTG5TYUMAyS7cEzKpr7jEW9h9D
CBzFwA7Sfi5bsy4AcqqWhsZwG9dX6MTyzL4R7rdOmaUv3+PrctEYjRcXjsW7lMzG
Xi2e2C7/gc7UiMtq5Ud9txmbXSpBifgRRAKWKkc9SkyCm9hdyQ95FI1qKDR6E6SZ
6RXf1ngeP1lYHMc4eyS4SEY/amHMoQQV57NlxNImuiYyJgKuAtphBEudHgYOoeDL
nfty0WrCPAgqyqWgtTK7V/be0LRkIsXnLOholWeqLfL1HD7XBE/oI3qcPTHKU0lX
x70AflwAMo0pBwVHIVX3B1tq+n/VHbnw0S0nKDpxQ00D6XzPPNlKBLzjs94fh2IZ
NPz/+AMdjPBwhAABE4Vl1V6lViHPfCJR3+m8t2UMTgcB6E7/O2SxZ0mHyBozHn2r
FA+ZwosyOfUJa0HSb7IxPxr0nfSWo8wKE6zXGeZcEjMzog+5hT4jcuiqQfZXfCgH
V9z+jXAc6VgWq/73NurHLDXkEpRwIJH7M3grpy4Aed9gI+r4UPgGwagJXBQVJVk0
xoK9do8692sDwMpcfnR+frhTaDgj25fkRr5oqxio/WDMbP1u/FP6tzlAvASuKz7q
BN3cwKc4Hc43lZUYSmYDoeMZ6VjcFGWjGXh6amI9Z2yL2qu9w3CQxpLUwQRy5RZL
4wsG9nWNfBU67limraV3gTcdkDJqHxjeIfBIGW1Pt4AQejVv/yna2EzESE3mSVjd
8/qGiAAJGYtpsfWCW6bnmpqkQzHkUAyCMPFKQcpzAOrrJLJTpChhZJ+Vdqv3xs0a
zZAxPfmjxsIiE8oYr9oHaxU2oJlHCDW9y25oN5WbHUUT07OnQataSBBV69thzAYA
YYR9yPScqeo3kv9MK7+zb2Lr0N2XD2GXYBglSHfo5weSzxsehLrkzQFB8jlwQVF5
64nmIR27HtiYxunL2weibdLVl9oPyCxuiym4y2SgrGnxZi0E15Gry/daGn1iRSnb
cpksPLUJH8/hw7Gpz+fUegvTfK9BB+pPmGqdL4AU3sJ+MLlygjyWvkqqvhNaaR48
Dvb95P8mNF+MD/teIoWh1S/Yk9bSSlJTDPvMZAtyFAjllK60EisfMdw2WFU9S3Xj
EigMhhG9eXV3UT8k1zBCU8k0j/lLURQGdkyjtfPHmtzcbSY9iFzPD0dKUZ3CK1Or
uF5+FjAP3scG1f6gdC1azcCRoGnekQced1vMV8xRTsRHK+fHHo0Djy2BVcMDBx74
iH3932POncNqX5YGlK74LzJqHP/lpObNhuEIVcJ2T8wVQPiDLLwMuRSOR08JJdA3
goFgiCrLC2YXu4buc5YHSO1nd5ggDQ7wvZttBYL7rb5g7Vaknrh6AyAR8PXU6+Bl
YWaClsHvzapZY3NIW/j1Sr98C5BL2575gc9agOhk82uc+sF0HWF7aRw3g7Me7SSQ
fpCQqpKFKNd9ooC94yjP8E9bmoSSsA5YmqKDdJ28KYTfzqi3L4GcEYIzW4Z+IVhp
f/xRo1C2+vRwG3mbbRipDDA1A7srFH9J61NNykWAo3oNNZDre0vn+IJ9aqXOW8Kj
lPhgfwHLEOVuBb+j6xHWcSDCiXxflNlyzgGEThJKubB3RGIWxsdTvaDRHzf4PDPJ
+koM9wDYQhNICIRYzseoOzRiyc9cQma8cuCHmmdTQzMlXCCnE+RR9CP4OGm3wKmd
ZnzvnO1FYP0CCKc5+htpTOXEge3xWesZ650dt7ufj7ooM+TyZk7p7Xp7/pZUNhsT
+4lESE8SoAAzBeWdSdonW+BhtvRspmh1s0Gx2y8HsH+54rreAJV+R9YDMraJ1ilt
OFMtJwuLWHJ7E+AvPR3lvDnhsfsxhy5RrXNLVnUZLQ9yaOoia5+87wF5FEPbrnOG
hIraKVz7s6OgBA4K01cfAxaya9DdjcSs0f90dC27R5H2ZAzs8aBHaRj7zM4V1e9h
EdGg+B+29jGKdPyXK8YXsIqN9O+qjXfwJbUfpNFyckH7x46ejWDmSIvRdQe3b1z2
wmG1gzX1BN6p63xyLgAQg2s3+nkfynDm8v6RZ/wyyZ430acEu3a9izi1GwtwjF/9
4rVbhoEXzDyD0YJrs4exC+wNuYf/vnmTCZIhEPDV4Ac0rcH7x0aiNnquG/Ll5Hub
N98H1FSgSsT9Ly+gZD//Sa6WADhQtakTqIfSngcVY3X01EnpXjrrALBsf7oYQ8WQ
iyFZDT34YBjOejw/Jl7QwwEbaqz7po2mXxqyBN+I9x+c64USDli8lh7sgmXCZkmi
4jc7QW41AEpUwEMRLAb4VkKFj8BNo3HnwJzqfYFadWByr8O4UWaq+FG2fqjevBBo
EOL+kjERVVlzXl/7UyBTv5ja3DsbHVEexogMJ5Y98FQKlgqLNStNuVdT/YA8l3S2
bhh6C7EfuaBKMycPDfKzJsMBNj+/XFvsEWZr6d6wVwDPmT7Cf5jtLUDGEJmxCPud
dxYtR1J8sH6uVPCGbkhaMNh/LpuHi7JQGWWx90OfzoyftKA7pviHaXEJTmNjEYX5
MHfozivgM3xQz4LXtMmQog==
`pragma protect end_protected
