// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:45 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RvNDTH7smmg/+FFoog2mp+dP0ssxjX4clm+JGlwoW7zIOmP6NvRtZe8ND9mWrjFY
gYJv48Gym3ixU18EbKozbznapgGgxdHvMlWnIPfNbNc7bn2aC3DEEP6TlIGkNmcF
Es2kEGZ2igRgyGpRuZZ/cd43/fAVp5NmrhH9mDyKS2E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6736)
eiyR69XG2UnEKohV1aVecV1NmRgK5JSdrV9B+wiv3E56J7ldX9Q/WSiiU3sKu63c
mWNBEOXqEHC7Lal8fWNy+Yf6bFE2bKPr/d5ijB9ORsqZx3fnPRmNcdNMYtenupWZ
JvhBnWzXL5zpt0FlUfF5NA1LA4sbgOAI7mNCrrJ4tBIdfAJk1gnfLPU4iAX1CG6K
L7w7TLdbDi7mlpOwKa97vbiFMmOymCK6JIDYKIuM9DiEwaX97HxXRYoWtdQSUtpX
+g4SZPnykBDVOqzwpSfmBb47xht9jEkSQBIM0FEEPGxYoe8KJ0zg002ij0yjySFT
u8z2vRtIDEZ9Jh6ukAi03Dc4zK18/nXpK62M5INFnPifNZqCao8EX9L6RVkUhvCW
Lk7gTQyvCOoT+amw2zX02ILOKB+NZrTVRG2ZVlkOYSMvHKuHEzhYxlCM9pvzlysu
dX5QevnxYVk7f9eiWKyRe9if66vRbp7k4+ulcQ8D9/UUCweaHTBGSBXBJ0tr1kGZ
Hrccot3/gZuXBdLflM+SNhjnc6w6daBvNG8qI7sTpKDgfG+phpmD5eQVl6Peo1MT
fq/tOnw3iGRs3e0BEYsFQp3anehwyFaQj65vvvW7zzntR6fYiQ/zE+5iyvyb00yp
l2o9er9mgWxqzJff6G0ucCPWwruCWWp87BjcfvpZmvupOeOGD2veAAPc1opxARP1
LdJSTWmJC9HsVm++JQWqf6jDoMMy9bgsTVfMKM8s1Kj1atah84+FuwBB8D0C+ccQ
7Ay4pQjTKBpEeGcBmCmofKcWXxBkrtK6vHdT2FYUi7LoozAbHDXuYhJEP0HqG8x/
qwHMhHH2z9Oj6dX5n2lpvBFOazc0LWI0EHds4dCw6aasOUTudz3Cr3/QP5pGydAi
LKZphR6Ub82H8DkP5XwaeszmAxluaZu/px3WYmlTPOlbxxDfb0DMt7e3s+P1rXy2
wxlZt6Knww/NJhAgUguBhT8jL3rOFeoV5S6oP4PcSHEi0Hh5eInV+ocI246x6wwT
kZo9phOVI0vEpPcDUhmZg56ayksk8Y9tmS1n0UENn0KeA+Ro7VmKkBzXpZhiGcuc
PJWOFWvmk5GPwqTj6a2QGZ1BukMw2hflRskiypUiMz3T9K4lq4IJ4GlfDprLoes4
pRC9Q3hWoGh8ko/fj020YpY7aran/999Wye0flNGXnPB0Sht0DoXowcfv5KzN1wy
xCRCRHgUj493jMc82AvIsA9gcqP2TauvE+cKZiZPD+fyz+18+adol+4Mu3lWfK6J
zJrPbEvEf4twJutJB4AGbxYYQG6FnJGly1ue+tLU/Zv6/kR4LN7JOhycvNYrxNd6
jB0vHnqImhJo39skW7xQg8CcLT+9fSu4vdBmooUz3B74/3u0crd5Sk5HyA5hhKj+
2jN5BdCmlFfr1osbxLg965hWI5fehDCPA6tGNlJDx2YxPnQpSg0Byrot2DdipR9/
44ckm7rNRlY0mDwFK4NTTo/GZp/HnV+iZASQMfglB0DU5IUOxNEvNjyVTeoAOnZj
ESqfYoWVTIaRuppTsTrl35z/9MVT0RYcouvH8Ee1LSpzmtDvGKeGQQmwz69sW7Jr
AZ2bi/NiEdAV2w/ghU3WqW2NZkPBH6f0xrXpWJyU+gfaW0ExCQv7kn9uols8LFZ6
jZZ/qtOQJ3/ut8L9XeEjdw0lpZ2t9dXtrFd87Wv2zHw3nulYNxsjSkWbj7g0cNFF
MFyxben383I0PEvYaF4oma/ULMXth+1KjbTlLstudfmk395JgCiH4LgVkeJZ5RYl
++aDoyOLnGDV3NWlt6BqfO/X8BAslERlCmhV580fFzIa2i45dYw7y69E9YNlFldJ
R6H4odx0ESNSLPKflzlnF4sNn5neYvIvnNXR6HL6B+AqxFkMJGEY4PFbUkB0StYz
jAbRVa6tIzhfHofTYr0caMgtGBsJNRowx2dqsm+9SPaylnEF71wT22QqRT7zUpEK
OaBrnFleXPltr9Xm2mKBs2n8Mno6J6Jic9OfTSjLLpHMHeVxso6k0vhlBkcXk/Vm
n2jEidXik8HCchFH1vC7Ke6L/wACW6WCB+28S0GD0buOPxk59MAGpPqLM+lFwfaM
Bge+XZxGIvz5/acgbj4WFNa2qpPomDu94NiyWJHhGBetqSzCI+M0/RzykGxykbFm
+zyY7ePZU/kW+R4cTmTQzxBevkfM1cKjxcrZGUfetobIb2Z4omdh/SNFYz3rwjic
z08ERrzemJMts29nKch83Qf2q0EkJFllMhol7HEpusfqYE64SZcihqIJIAD2Fx1U
fBpLeLrLtPPAAV+/6jTmhZtzKDhzXOJJHo5BHfx3dUE5thG8XnW6XNcYq2Z6Aa/2
AiI50Mvggp2GKrCe3h32TmHzsjhaiGkVrXp21euL7UjPmMjrY9iIYVEm2pARa5J6
j4aJeV6T5fNNbMptFdMr7YjX60gN5ckeFNF3GqxWjAxiG5xty02ZJApxYkEajXWl
9amZyrGv9ASfYFLfRrd8QVfvRYBvKJx5tPH4BN3pkc0lGgzyDr9HCnLn2G4tx2sk
qvAinTNi0zvYlz9Iwl4y4KyRwfQAYwP1aOgFTFD5O5GNwseRbr4u0cIPq3EevV2z
xQruxztni/FZbSRPV3j03Tyr2bMTVYdHVopA1TKTiOaTudJMZQ3IXSC+LWa0kLUh
14ZfZ8pyQrbNuP28i8zyyvMwuyt0We8er0s3+G+HLKZKrsjILa/oPBALuHvFQDdq
TisyqWppyZufVSAyyV2SWqe0l7vke9U9CZA1QbD78ic3v9bw03QxMCETUFHSaDhO
N95e02jgwf/zROrjWWQFFCr+oCRp+iQIEtLmK+MpLmAZChihwtfegwEqTliTuMed
zSo4QxxP56hgOblnJziwmmCnWwp3rbGfCvNhI3we8JqZ85HqrNzgc3cCPfaXOnGQ
Iu0yATOSUAv0Ivd2W1mU5p+JvnNRGfaF90TKktyufEVm6lnwhwVntSPNmWwlQPUt
ZvGQaOkvanYpwuo949qcyyTGLYHzHJ3h9FJxq0IItuXJO7/pOgPwuFjX5rfUMSzp
yMEj47E/7SnkWXdqvKIzSmNWz1nBpms56jfbNwzq0agC9ByszVHmyuSsWSRk6VEs
e7lODol0IVRhEZffx/SNGGd7QQvEjaPDasRPoet+CIbkqSAVZ2u1g1Jg/RKl6UBu
mq1y6k354E3u83pj98gb0deN0akUraVHdK01Rx9ZY6HLUzfZpTzGP7sHlH6DVmhX
aWwHXXlXLkCMIG19gQ35Xqm+iJGUzEazqfSvVfxrKzdS6wWg8iFQRHk35ioNOnMQ
K+GIHG97y2vtVePAANs9ANeECmlX7nfQ72uqU/q3leTMUtQmlEvviUwhL1crSdGq
uXjuBgBxxED5VrFPO9acPVHAj8noTWRHj7io63iLGPAvjAnTgCfvyoa2DS7m7Xav
rSU4n0HASB6hhR83nqstDolcxwYCcPtmWQvEscNnbG6b4tUIy+zw2raPQl/gpCi/
/NcUNnn0SKkxhCfew+khMvs9OA0JRlEd3Bj1a0qsXqTx8tUXXyBzWXbI1qYwkuEy
/e/CoXtaXCANdD+hmTfK+GanmnblRBwIMy7/3e3V2l5WxxNpBI81Kev0mRDKl48i
2/4sLw9gwJ/0Lm0IZBkufowbmh7tudZhKj5ZVzmafbXCZOHPaFpfd5kdF8pt83DX
zgExDy2v8m4OaS47Z49v62FeaMaG0L2MyslrzD4N+SxHWesuENqyT/OMAt4z6jlO
2+UXQmOLkRql47kBsYRdOPEuvu+H2ZspPuEKDwqVQHyDqafT1h/x+ucytRrvyfQz
lSXHfx9u+9DVtdFpi1hMroQ1HgQmHPrpOpsAhrT48WstPQtzQ6rBCGUujas4QfTt
GESSsW5AZhmEnkjdpudQLIFeNosla4MDeYDoKSbbsqhcGDX9/O/mo1SfsjeOaD2w
APfTwM6T02+2gE6x7HiUKKZJZaf2oaybxLsPPzDNt3GfBvXpc4bZwq3I/9GnjF+J
AjbgbqjLCVIK4+EHeIuH+XtOQvOO0RygFrNDndkxA6Sq4nFxuOZ6xuiqVSpW7GCe
lnhO+deWXtYUu5pBSuOy0CdJyFyp7pstPk7v7QM9F6QoiwharSxA6VA8kHznJSHu
Nq/PajJSqnB7iLkNe3FrWeCYqDf57Q92QM9Z7mODLdgJfmKE/b8r2FSIVz9XCQxb
dOdzKPjpJTG7Bz1ai9P2wWWgVcnscTOp4fMXGZ6A0KJzzi1I86zV5RrT72gtEa+X
JaSJBfROb4TmXPY1FvX+z2N+t7ej7KGp4xZ7b7LMbvtGCdLZ0eXVqjaVglXJWLHA
508AI9z/d4oS3QFK3lE6/DeBV4oSCgoYV1aBorKuykji1eeonsi9SZAUz3UR0vPT
/ZCTJ6hNY6Jpm3P+VFo9bMROTKsq5sJfnvlthOkP1Ev2vVC+FkwB/I4PaAHas6dR
ysyT+oTsKRbtdbp70EcE3/fINKzN7nj2awxpvOdpJH/pC5GTwBPUzMNcDqnDajX9
cVTFmgvvQJ9rM+ffAQa/XISbbIGU7d4g4du5mc8Ud/6gDvK+Z4g+ScjLfm+FkZDp
TgE6DVLqpMYGspYWU4NoHHZxBOu0OBZEP9nLymUuEU1vI9A5ic9HKYJR6T88opdC
/BZ08/RkdLI6pVl6PPbZ3pYvc5WCPICa25xKjfBeayjer0GF6XLnc9WCL7AmFoQ4
wEQ+FT/6fwPF7pnbgV6Y6JQ1NCu+wTl5wL9mfz4VGkg/eMlZ4K4fw+hu5kserrio
ZSSQqD0WqKvSKT6svKWqsYFF1WE8mxG+10Em6nYn2QKXRmycEJf8e2+mbs3Whzo/
0dprrGcKyQ6woyn1JjiiaGL69jmzs2SZ95tfFZmhXfEbmH4KpcSzUUaryBDhO3R7
qMhK7rOKLhKaxWEHgVKfP4iodbtyThkz/SKsnO+M9kWbXq5kuQpOlHeZf6RMA1Pu
I5wXCyevyJxqJblOaTgqZNPe6lhsU1iXDmx+quDe81/wtYmZ+egzoSn/zpV2bzmu
Pj9xKvligmwyU+uG65XxlCAD0nf8ACVoHZr4mlnVFMLDAX85A27FfdAOpgNflNTw
itmdCQEZLRjmmj+2IQZi8VZsAeAb3YFWcXZt7W3KZypg6orR4XKw8MIlUOjpCzMt
bO51Y8DO6XlqE9Xarmju4nV9uG8E0XqI5iDWaukAHSgNmMxg24R0F5sGQvgDBvq3
jL0Z4z2nL7i9ZEOm3V6Xwq0Og74/8fEFgUsJVKmVq79VUn5pfaQNUJ0g1TEtK+F+
Z+m43Kpcmii2+bWrNhZ7ZKREkkGqvBwY4/bDdr9F2wgq8xo/XjPhXAmeUhr5g9n8
Zxwa3NuU0R1+03AH4o8nHYoIlDpAbshD/oa4JaCUlZKzytZwG+GDswqISatXVPDS
pEgNo+3iPXwTsBRcKgOXh9oD233c+2dyfVTv0Tz8kqFRRrTcT+y7V+WwZG76y4Qm
NdXGJjOmmdfCeroZjaF+RZd1diJ46PsiS4Zr3+90tcMoaU4W6vZ8oHgxsLmC/Pyo
JMYCebgyCTO0Gz1THOHfS3xa5zWhFn71E9jI4nN1msVkjWn5tct/DIi1pbkGK+Aj
1jjmGXcgson2OmQemPJVAQearLj8wBl3WvsZIbMLHYzjkYIIBJAxxe2K2N5IwFUv
2X9WFSXcCYdDdSFrJZUDgvMaVAkZbwP855t7VG6pADgGUnLBoHnASWdBHv6yfHt1
Xu/PQftXs+gH/CzLnUyU3vt3/I1K/BYCmAsfJBrU+KZCGXMVKxpx3t6LncDD+zWD
+/HwfEGrQ0+8LtOS+iPUU+AH4jZ0SdTppovLNfp+lY7cPwG8BrwtXjtHoBSjZ7av
uhS7UDjcdD7L29wirECYjLzQcTOT4yQDxeDiutmZa7aN7CiHZrcOgUNrNrI/XR/I
KaqA2lqkNsb0eXPHgYu7jZTq7O+Vv7Hpsotljx6BIIEoPPB8HdjFSxxoXFCNyF30
lmDDMftruc+1ZadcGo5iWLJ5S8ODZLWbK/jhxdTWHKlmVTw4BcUqZ81CChGrT5qf
xyQUxHCcdQ45N9g1h4+IvwJgwTi8yWz5xgE8sbKOv2UX5YIOl8lcxuJQCI4eO+Ze
LxaihUL9E+DAvYRkLbqJnDsKxSXReriKPAi3V0rh0XrCvmX3g2dmmWOLvobfFrfY
85ZuFK9hyd8FHF1aeS1a3N9e/kIf5PZnp3sllRGsiXYB5it4n57yjikOX9oqVUwW
mqgyJVP/eJdXQ1pWLk7NS2JTt5HCAJnuHAk+YkVqR4XQEOlxJH7xGNxl5kUgKOYh
/FPXK3gGHMDB+wiblYg6Qgn9GhZLx/HtliKDlPDsqJj5Tts7gW2yysbJIjuyNhqM
IPaVJimwTvn2I/RpQ6z/olB0oOUpvANWkwuoSUPPeHWeaXt9MaPLowbjrh/9/jeH
zOaGzJPtN0YzkKV0ea5S12RzK5c6RTxHPmRWViV/B5VMFP/PRZLK4aoMunhIigvG
sTTAxl1FFSqXpJtIVRy3JlEHw8c7/kz4uJLkmo0ba3zG6u10bzm5JoiWh4P8r8j7
Ts9XZblRSwfY8f7KO9YgD7o6/1YZpjdG0e0IlBYSc9ryaIMGrPLKF0EPoyzcEUOX
HL9ffh2cQCvxNZT9RmsifhXpG5tLXuwmzAWiAACt7owur47nzHRfYYX1utdh89jI
j4OYmVG89gNbWFy7nOFxDKOp0BasG0+PYT3ZgTgTVlADrbTXI2tYQ/Z09zRRT3l4
b25VfxTgctk370lW3S9BJimMW9K40IhNYnRxKhkWx31djWScnd4M+Iw/CSOH8oiS
lU2O03G2fnnxv7krBKDUrDGKcR7+DLv+1R0dxggB/t+7R2Y8xnr7ahgWdowiV8uB
Sqplvh1tdvwEkagsEqPKSan3iJuK+LYeCKLJZ69z7NnZoPVEN0bmzJciwDQlKofT
8cQYPmXRTBy/JcBuyWvgWvbiYL3VBtD32LrhjXCQFJMBm12jywVFDrJi2+gjiVK4
hjVcctRyXNntxeEYuNbDFTfdkSZD69eW9EzbyyIJtorRqyAVjNItxYGAQ800RSon
lis3d0vbH6a73oxPA3CkPJF4FVbEIkCCeklRm7c79RgOVLtjrniF+4dlArKh83RS
qPib9PnMAy2zGXzAWkcUa4Ed3m9Lw5vVrlxYQTv186+k5YL0NJgaGkK4++vS7/sC
I9TwdOjcy+zzNYV3SW/aGHE26uK3jqQ7FQXw49U771scQ2ypfl3yukg0f1mukaQe
YaAI9wgvCct15GNToQyQGDqBLhzSSjjZTrdAlDfantM58WrI954Qc2Wb3kAPYZoU
7eFHQLjjerGrYDJtbvkyuiFIV4OLVVUPEx9mZMOQJyjOr82FVWJY6Lulb8zS519w
xiapJasmBOh8ryCGH7Iz5RYs3iSNZofedxudfgUGL9Ay2pth6UXVxm/V65ic8CN3
qP8F/pY1242u07Ik9sdE4la5CWmloLxmwCZt28syAZD1H70gFCr/lqeIcOjF6tH6
cbcaP+zOldKFPKQAZyv6pGJlwnKRARu05Ace+sCQ0HVAUUvsg6YEJiuhvY7tdFw6
tzqnjke3aPOd+IJfkAfjqmL5lubr5YQTtsdscn2jvNFEpfAgLrWa/as5hOGZv8Bc
BeAli5xEb7R69cItj4dTlYeQTiTklmoytp/g+ZOF1e0E/I+s7eyqLOtn+FBAIVGM
byd5R3IA+N+34FuavpO8fPzlZtTtZSkBXgBNhS0xn1fBKt9lDl30JNMrZSi+nSzS
4bHuYzaj+iXkiamVARkiDxZrQ9Mid0M3okZS32Ju8t+OonXi4UKf0iLShKRfdN99
HOVNAKSvkWApjNnXrnKql19ixXjBjdedMqWT5YJ4KtQQzC6hj8j+OSF65GplM4dR
1LCEN4iLxm88mQQx7lsVhRAT7jB8OnDpZz8y1lOK82lUPa866I+b/A6nAAulFiEB
qYf4Hc8HKsR+ig/l9OEdKIj1pxC6RFa3bcdIUZi6C8KeZT0hWW0ZOJyofX91HgBJ
ERlcwVwblqrrEjmxd9V6TPK9jwcWYUTZS8VxpQR6K7Kx+IqSYHWBa/qhMr9t0/p2
3Cq6hRxIo6s7wcS+MkZ7NxpQZbcUUJWNTRY2rslFNIU4pjDnliSxVqkb9srGgWZG
wy3q9NNp0zHQsWlTiV6SwUDFY533tKvtfzWDNyHmolNWV77eR+CScqywAqsYp+NZ
hQvHlBlTHNM8x6/0MB2yaxVdqExrqGRlPJ0YPS9lBXjj/PUgcUfsuGh1hNUUuXWd
GJF+272queUCKYmwwDuCgrltYu3R35pSVtW9eUwE4UaDorE3okPv0QutJVg1m3C0
WchvP48iR5PCpbZqWPgFrw68NVzZQrWC2Tufrs4BQis7p/ncIMEgShqsgNqb+CiK
XLqEzc2lJfEojZ4ReJfE1jIW139K2AbDf9yTBFBYAccTMHSPkJBo1s5LD3+Z3cqA
QnixPJk6UKpNptrHcQ/UVADgcCWE2gVrJ8QxKHI/E6rP3PsehvsG2HM2ne8XWibE
cxp0ImSJjcnKIuy08VvwiEUp0BSbqayGZFxs7tkoYAL+n7ogTcLq5KAkS9m7Z9zU
vb5zkKZ7GXCwWS+zuVqcOfn+gBIp8cweGjk487amFHw0KJIpCCv/BbD2objnYqMZ
Dct/9Cgx9haB6+b7k8pKZKXfFf82+CcaYlfjNrhZwo0bNZ/JeETnfY4WLpFlyaQd
g83I9wXKJ1BxS1LMiAf5mPQSu1APa3IJBuq4OocErqZcUEK/aqJaChLixVdKwRO7
hW7fV5Ji7WdJ3hkzS6+44Eii/86N6o4XWHRRjWF5ujmhmTycrAvkVNb2KkxvLjqv
tXwoTk0nxmLmIRDizzTyARRtosRmnJ0vI5S7LxwC2u7Squ4ivfjy6rtCMWdJw26P
iGrJdfz5iskO+MFm8vMrSw==
`pragma protect end_protected
