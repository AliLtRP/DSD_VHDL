// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
VjYHW34Zb4Y4ZcvRbTxK6dkuncL2hJmDP6eO6OBlFq8H8o31BibkJUjFxBke2576GFDtMUdNtOKR
xr4/fotgb95qUw8P7fpi8xI4Rtzi0yfOV15BjqKAifQpko3UbB8pii2eHT8lAQmw8g6F68E1kJBU
/ikLxHNFiifHcYccmaYUNVaPUcWUHmbxOVLJyCDq4BLjFGmHZE2fghU9SWAx1ykhF35J3GYD5wQp
liuLh0rHyaWbPanZW+muMRaueq7ZthXJNTfna78NItKEZQESCIrt9PzsS9DlmnK1A1unWpuIpobk
ZwtBSq4o6eC4V+Z4meNfsmqwBMfvq/joroG/rQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
fNvldWhLow85ohc3JZ3fB+x1SDxuJIF6Ur52RQ7STgE3q6ilKPrpXSjh05KfEjqb6f9cinqdOfZl
PIXXb+m9La4b/hkkrs9jQ417SdlYVFnNZt41Y6LMSdya2TU76om/PCyi8wPyPAUl32c6Gq8bM6dL
BzZ2Z8TDJ7L71udXmaI6evaLX9xQ2LDjG7lvGhM1fciHwL9nIpUcHu+wKqVNmFFlVlS501rUeDhR
LPr/W43Cx36gzKLm6FfBSDov8ZrI2qm3deReNGi7MBOT+T9jJkaqj/aSoHRepsbkEm2gbuCwq7X5
kJehC16RJqtUZIKCHD6Uznu5kxgaO+4FzuuZKtI7SNqA764P0xTRmsKbKvbUiOdL2aC+UmmEsn9E
WY4o0MS/I3KnKa8+3u7xicRQflNUHLgOo3UkxRUWImpOwjnXDwfzk+ZYu/VvcPkBQeHbWFy+hlqQ
/v6WAJB7hn5ngWhsz4zO18BKpszxC44uCPfVgmdvSQlKS8jY+UVrZdX4U821aJ3MpNuUnQVmZIbb
s3KZjJBaGfe65zu6d6TGAkFCmbmno+mEt5akUEcdmTWyYuekM8stgLnMyHJwALLr377/ykM/tTMg
Y7x32lXGu3IqlHUWLhZdzAvwxH/wMdITEAY3Qtcv5LbHcamsyU54K+dJnKKW6k7mYQNYwKW5EfBm
1lqTYBq8Qu3Msfc6AXeY2bkfMo2JJnOgWIyFZmCJlDLixNQLrK2EBNxS6YOCmXQ7J/far0AzAAPr
QHPrrPqvCTM3wVGAY7NpfGxs6xDhCFAedDF9MNkpZQ2faSO/cBYpewNuE1TBSxrk5AzSKn8g9LfN
pgU86AKUturNTc9CbcT1StORucSRnNUnyUVhJQyhR0HaYL/Ys2Fz5AjJPb1x85ba6NaSOjbBTcvn
RcPFbjVHQN+XVXiZ/FWSGmjSjFDz+x7Ze8sy9v0cbdq4Dql1bOoFoUtoPVAQIzfb1zDMiVRCs3WJ
7qJQfNOJZcTgyPriotbNNCopzKNzmknu7GVXZAah+1CNNCMRo7KK8U4jiUg4efkr9wsji0OEue+t
7Wo1SHG6lzFuZiIPc5GwkNBxlQPPBPgREF1UZfi212uZENDoF7Yb0ngeDRilcU5Lm2/QqDd3Twp9
0+lEQ6cKtPLrT8KBd06bXVi7rqeO6BHG9WwMTtAnxWpEglRKJsSQve3rKFafN0RzdwPphS/veq5B
eyitikG6ytP5aOCEHJ/hHG9S8SkKpkoY0JBRGuozxyZYC2kZThIhTE4+M5laLUWqhCexjjpclEp3
wiBP3RBvpDfjhLqrDrqGzoxILqv4tFKoCyax36LAj7U28aV9U+sagcaNjy9Z9ushPryq5MTgNG5g
8TRtzslEAcN11szI1jFcpCtvkAgQ5U+8ONXxwsDnC9013RHWP1yD6r7dOsXKWjmd/GCrHQyfEFv+
mshm97NixfXZwRWW1Qee213nzbxoPi2xaSdXkdhJz5htgc7a7ma1kV0FLufS6adgS63BzzF12naP
E8rAHCUxxmdJiQrcYvEnyX3AUJh7pmwFAwiHuPIMuF5A1eXMuJjz6IpKvpQEkDhZZvsIk+V6iwaB
PurFI/aCZ/3nN+UbHqZVcTpvp/v74HPSeP+2giF05LK1XUxFz7E532NWaN3oa/FaNDk8pafacQP7
h+Dqu2puTTCyXEZZ9Z4Qx7xtK81ZLbUCrf5nyNcJd5xCDhWGv+SER+PQPZ+KBWOg4GIZ98C5AJM/
JrVI1aps8gvFKb2BARb5k+Ts2irjBuDjlRdvpcO+eUWb7lvvLVqbvP+8j7gltPuL47RAlcTqRSdO
NFmctSVD6O24wLl3NdiMBesMNZuf3Ty/MoawbKBbnjqBPNuBuFFDSssLywFg9iESZIh48QquI/ks
GXbhgHKHpb8dFACQgLfutN3fn9j6JoX0btaU6J9lps3g/03FrnhmJ6NTLsF7WT4aqaAFQ292tWvX
X4YVWWk4ipnFohz6h+WqjGCjT1DPzuknjR34tiKraOJ4k3P0Pu0Grzf8Mw2buevNzhnd5u4XIQri
3eS8VarRCJlDwOhRrvx/u3IcJQJzEfp288VBkDsCe1E63Tl6f5oaFn+hwpnJ1xDkhiDm0AXCaT2v
DYKl0pELJvzacuLQj93scEyp9e5ZqiR09p4Djw/DHZHfJEfHJiTRgrmsKSSk7TLfAiTzbTdNfT9x
tVCRQqeYNra7ziBUFtdOy51nh9yYlQDg7yJEpX9khdbEQqus1l9gtvJtYgNlCgWs2bPEm26fNnmJ
yjnt54gpyx21wMjI7wQBBwfpaEl2cAzQ/P6jTHX4PWhN5Jg7MU1C7ujsXe6sFRZ8TrE5WrqF/lTU
+MElb13aHisjCAGccGz45O07Y9ATbSGmxbB4Mu+ASnHYBiA3rz+vfh80GvttxsYgbmtrL6DZQmpP
sqsnKsq4zz2Jj1Bk0MbUA82Z+35tU0fT4LUTBhLrU4KaX/1W16TI5aqhehPt6fk53BP7wqSW883E
0am8fjQB6Ij68/bzQmkUfr2XcMp+IMxpf6LiAV0zbIF9t1pEkO53qsrGcOTmyOLRmrN2WSW9Q/T5
y19EH9V8UFpSAxQIhAJji3pMN+/U/EMdgddU045SMDqaWJomNIsIImMDYuDICE4KzGCMoSbq+J6G
o/IQ1IeR2pI01EOgnrIJwq6RhHGA3UG1Y6Zox4PJxKv2CNff5EpFqaP7m3O0eV1/5jQb+wP2HPVp
IWiKYgqjTnkOFnPF/YlwbVeb37ijMRBovS57z2XW/oghgBKmJx4rtPyZGi5V6MP6uqUvEynVEEOR
90xrEzADOt1r1GN4b/CYaTOobN1nhMAfHL5e1HsVlNVKk88DqYe36St+/1O6xh3VxF+tD6xWA1wC
tO+TbTNj/2RTEDTn/jhtjFlBe+zADKp2mPu16yUI6JRVem9HGK0CnjaDSOMGWxfKoC7R+oAI5Hqx
qR4D+1bCCrIRNQPnf18qlMMmLiVXaEqNA9XQWgnCwKn9zxVhUZ8WwafOniTs8xneNRIldoYC3W60
EK4B+UNjt0uSnb/GYVTQALtUSKGcXRfy2QGUWCgBfSWqrkVWzdp5JjTcsOeDSt7xMj6HrlSATtzy
h7thSDKOtd8XRgftanrIgkXfSVyjvv/+nXESDst83BM6FL6IFB83oYTGa3WdD2V2GAGbir/xHStz
jFunfTzlVdQOrjpHTsfhqbNx/LM1ldi1uGCud4Lpj62tXmi38IMEBNvhRUqrBmfC5p9YnvQKLz2t
caWycjw4q/0kQKv0Un6LwBjE+s6RY1zcV0OfRjQx75jyIfDtd0PN9yfIBQGgv0PQTiLFyPHCvApW
1WNiLpMlZAEsE1hu1xLgHL15zQCRt2rQHrPJSXvH3x8T2A5XgOgUsl4PMPk6lYDLo2SMOSij9K0H
fmlnziO6D81ztS4OH99fFHQ+ATCG0FFgdfiLpJjXfyt8rTowK13+EIWtxybMvhH4vV7ZMuHn5xEt
/aPEo6hV+89S/VagcfUmbJ2DVpTbqCVBrSRatTvTo3Q+vRlGmY7EOuVIYhIp+q0tVrFxxOWP3eDp
2Aox1BmDkaFCKwNvT1zcTucPgvYobnGKegbYauW/CDk/+d93A6PDY5xQ/gQgJnJfQMX21yrkFPZn
8DyqEsDO1xbz8bk8xZyeBexRZJNMiTBg9LjGHxGfgWys+QlOU3yeLAmJFQcdFCpAIhuXyp0ti1nL
9ofVvgtBmAS0FUAdQ0XkG0WK2AogwClre3rSulo5LdtrUAkD2EFthU9lEux+NAv9lmhlnRZOZ+az
lbZliaKvmj/y5sAwdmqAov/XOkC71PKeyFnwZsC2e+EwtegnX76mX7U6plUoUVh1FRCA7nDAbld8
MWAsvpnNJfVmdFHuEZGu0vpkbQ+n2nf+58ayrxmbgjxrNFEWsTGrq3GdlIVHvXPNNff7aegbxEG+
hEPIMQG2yDNiwVZqFfl77CQ5XoM2tISZncPb9ivodCk1hA9eikqpcC3hhFkrZWVm6n11mYb4/6/R
JcGzQQM6hNV5NsvtBvQAySuj+bnCqS9Mwiz2Sp4ncDAR973sZ0F+nnKiEG60iYjC0+jdo3IROJb2
gofhuARFLFpAhNJN/ARzA/AoKxJbv0dovDXTT1z4CuOzquSJQ9Gx9KFPZqvoAWUS7cK0J34TckK5
iw3qefntk7NDOhBbS0p5AyPY3012YIHic76eoqYD8rpdmFS593/gTlISSGmcwx//Mv12LjvzngDQ
Yob3SBOlhtB2rtibIdwlwzSgp2pBNTEd+C5bO8dI5O3geiw9FhfBC1ro+oO4A0Ea+FIXY7v6XWVx
prs4LR+3Omm4OiCbqsqAIbYzVp19kC4wWSWalTgJQHnGmxOAsCJv7x3zFX4Vi9FQZvm/IXm6aCEJ
t5eImRKbScNKdcwhcNz2gqmH4Or4YGuiz7fWS+cPlQxWfsBrY4w8vRbrNFWKiUGgU5isFN8q1iXq
OE8J6kc3pVW237VqXpDUfE7KLWKDYdogekZ61RPUdRR3txtM5fo/LgpN5/zLSIBZtEvgmGqqsJ9h
poakkb4IZxzpB0aTET/OsXuxwPJy8yEmvjU49MXuuAE/O3K8T8bBDkVotSsRNvDnLPZBghnmjpcW
6yVfsp0L8Hb3djyfyfNI3zfWNosaNRMaLxN56ogqYsNGk3rvSvxk8hch+slue+GrSwEUaRTKio0R
VYyaPVHEa8m1VhvzAdScTU5Ey1q+x+nnrXLIfxpl0aev42uWYT5KFZ0QZcWcq3gZ0Yvv0L53l7Gy
pVoELV0JemYZZq79oaMjf97B00vP2Wj3LT6kD7uPm3Teb0/9sEf7Hy4fhHeJeAyUhVZhyZ9uIW2P
wyZHwqOzLxa0/mN/d4ChpTFWxJ+6qssSRjGpOHorpRqI0LMidFEwkH4cShv1bA7X2lGPZWe28rI4
3Ou5DwNm3MmFuGSZ+iv3E/KP2OfUYF10cvB1M8IP7YWnVIy0V7YcDWVmbHqe6f1LDsSF0a9O44CX
XwcW7aD10O39JakTOw+/3uDjI/X3QgxXtvI9UfTgw0LvmCtJjneY6xjnXADBd/3INOQJq2kZ3uA2
HZW01/M+i6jQlBrxU4cC1+qsni4gfMsFVPMZ5AEKcVFf+cwVmJN1v8E9rtDvOzw7FEWZwWl7GOrY
v4QRlai42+PA9haMFD8DJJsoU6MoR7gqqoxubPCqyno5rQmBrW2ghSN97eGoWZPsWG2A87r8DHcj
ZShsjVm6pTyeJ47NAsPLGtrIqZbxmJu4i7F/TIxkxS06ejeQNXp9VJwotcvY1wLDN19FXXPIBocS
pZeUJFp9qP58z76FUMW2G/upIDzVloeNAIOZQWM3jVL61+dhHMbLqIneHycw41hdv9ItZZllEpTy
CsEB0vlpt5lq4vHAxIRvk7EX0yDmuubSsUn+0/NY2t3GRbRWkDqS28PhwWQIRqqCxQmuYj1AaEzD
2oJDqlfS8WuIjENZCfiayF3uLHNgCp9MqevCHHxB7K/+zU56Q9cbtjTD0dHKVJjmXevs6VJahQmg
0kbNUQ19PVjucL0DouL8hjjdgK5y2GVMIbMK0MnD/VduXUJvhFGK8kPU9JcxTFz0JstXY2qJ4tSy
VXD2uxQwBC3woj1GL47EDtB84M7sSSY0svklokVGR92jcksDzKVHVOS1aRCadZhMUSNXMseIJMJs
LCF23GbIxxTESouO5Z/MhkmBgXQ1K0mzWp3RV+HIK2XAcECudNrQIiEvvGM7y+UlRZuGmFHoxn9N
Csq+mpWPiPdIN7SyfDXUPe8aKrLA7Cp0EM4/io4l2El7Iy7mmNSxKp763ta3rrecQFVK95Nuwcq5
aLdYYgkgqliVYRByi30x2hZg6C8MUrcFgUhpQ3J9dPuTRDEil5m6lOurWbygd3ufu0sPMI8Eea4t
Xh2e+7nKQETOPYc8rJ4dG0WtQaSK+tVZNR62RbHs8hUwRqHV46oLKpXJEM1qfGrc03Zm8xcN9/M1
12GhNf16bkNFMPq8d8UZFxGc1RQXYOihOUf1eR0T5cGu817Wwa83BTt7D5cwTKRSB+pxgF+ct/am
5v3dDxsLoWGoLqAyzm4+WRoR9z07LYyNXBgGxXRmgX0QEBZW7TKAZeofhGlDo3PgT9CdMH2FML1B
QtYYgZFozBAxOoHqOrsZtAXL9LjvJPHHizp433crAtRvsX/T0GXxM6pU0JBHnNkE+j3KSW4ahc1M
TYI5Q0aCj7u57uJRnCA8Wuzge09/XS7zMPVRZ75Zh3//9A1aUq3gwlmb9gam1t+39NF1TWPWMbcW
Uti+6Tm9YZjw6TDVh40PSGUBYK0vqci1L4kIXH7W/RH9D5dIcnAJds3P5tOvdaS8BL8QA7Gi9PbG
ptzkhlORhVkDjLM7EXGipUjQVH50CvPQNv6DkUCGuc6cjCUuUKJB7rslEKDnTNMxiklvmD6HlkVD
ewxXf8ioAfGTMi1x9qP8Dna0oBEm01lEyyjVWH2M+/uL61+v0AmtJwd90RQzSu+eVlkjrLIXGHw5
fG6Gu5BOiF4RkZmxQfGEGyoWXxTGOgbzXBzOw492QkY1TNTuhqU2X8/pf8U70RroqcCnc1lXzjDl
+apf0BhrkkqzxUJur4BMDG4wyB2Qa8LSkC+xeQ4G7Zvzha5jMG76ZeyD68uimTrZN3dwED/A7Zby
U6pdxt4KAScW7d+FgQpPw0cbmx19asjsIA5nYyB8ugkqEbGhultVMPiROu0vA/KOjCirl71JxIjf
BpXrEHmbyTqqTBJGY5v6XOdZ1Ko69m+PLByyxcFrsRbRoKkuB9P4cJ+Y9gU1paCVdbJnc751d5Sx
GqMl4brWQ+XtIX3fOAo6esiNdJZCGj6Rr4wh8Ap70qvMvO2LakjiUyUAlB3J+5XboGSvdFXeKXP1
j5to81LJjvO8A/lUMh7ND1snZg+pkIP4nLGzrzh5U9RtKg1O7H+8Vdh9bCbqWMfjbnbT+p6R0bX6
8grJP1RZSNifN+Ua5SK0A74ELdcaWQxyQnR+UTWWjWWJSX5PtuXV+1c4+GTMbhiow/Awc3rcthbc
fNbC6ti59mu8WNwTwE5IeywYV3Ahu27jXrNFBVWzpxn8vwpJOjztERG+Sa/yLzRHWwMWAriHypfp
zcJUmux0dZ1VolF9JYBXjJVsPX/5OhHzppAb6YGPgKEV62zLSoP1mCmXWtwdQRoI8OoZKS+R/Ngm
heQGKNqEfNtbcGBexh9TGwwmWiTa8xc9Q5CY3IlhNAtHNQZDB8kxUL+0U/IIF+UTbV184jDfFgMM
nhk0Ud/Ysc9dKXZOMmXZ0Y180bmpnu9b7szf/S6+RKN5cZdM5vbl+MstYN88yStA+N9Y+ere+3iO
+tJzS5SiRutJcKoHD7r32qEReXDM0ypm/+V+l0y7sDWcHGFF05pXst12AMHPSfQdnqTxtZlz58rs
xtcKAVKg013jvdycPy+mQL32yFDoJiWNKT1uoVUDljhD7MR/MHFg5tqq+0Yrwvn+gxYEiTnnDMAg
nbsYu/ciUFEFNIDyoENf2nswhJyRla/aFfJmn8Ls2i71NjybkQp2v1ZYvkmdLnQ8FZiO5kBAKpVH
qzHKNGi8KqCgL98SyiraVT0Tmnf60X79rMPYXpsN4BhY2NPdWPlPlCyRSNlatvPC4v53KRyss1n3
9QuwJogdcl8+PYkr1+c7HH1YAsjV419MWX/N7dlMPGLXUGeibKWduDHq7nCNhIDmXy4h+Q+FDd9C
LXywPJRBYiuo7SVZ1bVxa2gFQL8oyfm/wVnaXH4dZy59OLcI6mjCtRcVdEQV3MgCvF9Liin2DI8Y
X4tUcPHA6Uf1eLgArF2cFHOV6mVDw2a9cNjYZ+VQL7F9iaassff0RFSEu1VG/moU5vHRaHxkKvBk
jA6dl3IbKCzQWx4ahZjkCBEq9soQRSi5AAA6Lm9HLElFkmK3aEeQrUELsbBT1y7aGE38Ewypq3Qx
ndxtEXtVvaahRCoftcldksXx5+e+Yrk5EJe4K4Glmx+mi53YqcPAB7Eq/P8yU8aUcpNnRjwP0Ncy
kgEoHSE5wOKcAVOsxDvLu9GxFyI+5qqdm+oFnSc4e1AX/1xfIQ5MIHyvmdoMPAxxiURFleEutZJL
gCmv4YxcvRHrmD14UAWwfYE+bmgfieNE79jvC542U4S8Tzdtt3kmmOEQz7B9lg0efykod+5Jl8rd
UstKtUKuzbc7Oy//CSXzkUtIOMj9jFgvzuoMJH73Aorl05An9mXgVzRtkUC1dah7+DlrvnFMsMng
SCffICXwLaGoXq+w09LX6xaGpSybUC6vGoNqjXPz1gjMPjjKHnov0kBmmK8jB96tybHZY/YyXZ5e
MXjHGYeAxPyyki9x+Linv309VpPg8gi3DRQlqEAxYC5KEdT7WHH+Q7LnjOm4eU+b7F9Y+xCDHqZr
8SBl7FBqK2EPu2jm6TtDtjX0HnZG6muF6r3/k4d07f9EBdBQEIBVph+UrwPdwdd1WV5SgxRiezaZ
xKKDKtP3FuRZ2kXX8G+fMSm7elYXPO+MyLfJc+gVtcKvW6PWDdMjShSwvanN/1aFZ5dY2SE4L2ER
NFu0a/VKxYkKatKbyDy092xECY9Zafb7MEUXeft59SEtMJ9RWRg4R3xCoEbkeOc5W5/cEEvcx+wx
qww11egWT2L9++OKRSb4oVDC36jBfI3QHWmp9py8e1lOK2EY4D5r+121L26mAaIFy7u2JR0NXPos
Aeh91HHYY1WFrOfCLvX4h5YxyvSsepX8I0yD8j6AI9hgV9lfsgNnc1peHVxQUoVv2TpEjHK0mT0w
m4qd5uyqw1DWsQqDn2XiOYCoQ7nlLtHl34WWthTBj/vPrJaWUuTWA2oNuLvuRrkc3YdReQy0n7Ct
aPJbPW72t8r5LxOGIJ3l/CKac8+zyoRkWhGrWwc9AWC7w6qdkSBczSHBgddaMLMF+JdAx24ZEcf4
OQno9Ml6wF1coP36zcaR9/Wo/N5cli67EWbab3KWXY4iCB48vVb8nHagUJvQMR8VwHqO+/fdN6XP
Kf6o9mayi6/kLVWxo77NOeNCE+XWSaKELwJIoQTWVGy6eyFYMtIgrYE1IVHt710jrR6kKFDmdK1r
O73D48mLBFpJSSkk5O2wZ6EB6AgtiP9eIu810hHH3kDvn1bavh6qIOw2UkZ6uxZ/oJkTt5bRHp3B
2pOIVxGEiE6XyOB5iuXJTBRoIcGYB4W9DdINJcuycIpVUy08QZza3fWTjgb0Tq7Q5iKx6io/KvUv
1GAsZZ58ld04EyVCQyJXa/EUqC9QYF5cjgeEzjkul6V7MZJi+M32yS1ze/jy752o/H7UDHaXCCT5
djYP39dIw0YI5sc4cGGIJI/v2VDJbt19ADO2TxIHElO4Bs2yaQ7+shDcT0DpVu6mdpcYFYy4bXJX
SQgJTXRnm5p/yJorIUb4LQC0PvYi+8C4qLI7Nz5+Zxq5wE+3o66nz2nJd+y+qrOf+DT1J4EDHT4e
tWkBBbU0JRcakRALXhcNIp8RPVhCwzOQCIqZcPvdpFhAZ0wXNN/RHnEcoAzRBd5yWeqyHGZpBl3D
kwdlvdRENtOjJsRxPDtyuUjEW9ZAhuD088hsFSW0W7VrKLDFnELvNdmu5MizwmKX8sBmbkarKJAt
Im3M66WkaFUtZwszMT+Q3eESz++IJluUVEyydu60AUas5utK+vfTE9g2wuI0/xH9ewlrk4IYlpUU
tT/eqn6cWIJwyGJCkkgB34K2Acuj/05yS+YvvvQJMyZp4WIeianERiJCCB38mloQ0zB+FLP/r6ky
wVDrzlURf80Fa4V7pmFHdB4b6UCnicLX82deAzKUNaCAqkstamXOMNUV5mOFLZTlzwkszJBtv/vC
BY92PZJ+I/0QvjnrMPN6Wy//q/A9gU3Yt5oVkzppKIPJbwTc3aJ5KFsW42xcL1/bfgZBfDVdapCm
bwadzWkJsxXJ3GYMPLA8F6wVUAVqdM9X9t3UHgeHyY3fXvyOJCUeQsnS6fqozfxwMHvvjZkHL5p3
5PPXV0LaFIPBmVEbervy0D7oJgCVskqf3fQanoY5tT6wkbeoEs10ZFYs54zQxvPbBHRgOrBf0R5Z
N78seqBow5uOudlHGxaT9+P7/Z2pl9r5K4Oy5CBbUGWd+HoemyGttSHZXbHFXsq3NoIcIoVGuXk8
jt3pCk1j2c7dZzBmVHWwCc+TCoVJ6N0AmmFq+CfInTmsrO3w2ezZf8CQxGrvWsyRTVZsRh+ZelIL
6coSyLL2Wo+AJ8aFlxgTnjv/j9BAQzUdcikyqgJrpJx0rYnEKCo5Fg8o/w/F0IbPL79uEDjY8Fu0
VSpPM6QPjcb+75gF6QxBDXUjQGCVIOeAG5shFhpnXgVwZRSVUR8RIPtFIheHC9C7inukHuJxieDb
kyrKAaSYjuopRpczjBHFjFH2EFR7ms4VfgPi9836+hgda0J5ggZxz2ZRR3hMRHZeltigWHufBuC3
UTmaboJ4g80ERLP7gYvdx614PkUBTXL4rKoWDXv20o5Yb16zuTFmyM4tB5EGCkH6dH9R/1Ghy7D/
w2ODz+TqQJ7eAzLd952DalOS46WA0Fps+1YVRok/4KOlDd5RX3CVQ8RFS6nFuvM239cN8P9pqmhE
/iKVyfyGphpe55gJ8WA8tghCzr+i/1JgIzTYHlqxw7n82EdS+FctJD9vzOvtNfnx5Nm/0BLjcqqn
3mrFOwCRkoxAOwqM8hlWCAESKQ6JhSam+Os6B8XD/S7TEMVaZbat8wVPfguSYX1LuzaXCebIZF3G
Z1RMK/XK4hpkEsJRKYJeXTQ8pDh+QxV4a24mbf574PcpEk6lR2DYgui4pnuRCuMbZzM=
`pragma protect end_protected
