// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:28 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rHeZSyIBGzphTSXFLHuMsE4Je7rEIfRQzSLKnpVaJQ7zhazf7vGjfbiVdf5EzYNP
nI45uTOVvvm9vur41bWI8ytxgjfm278vU6GNp+BAm6i0US5yZVnxEO/gVTMof6QW
crxuinuLlJ6QATEaPfdUu8nVuNjXzVJiUoj2wDbeZRc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5696)
FQkvCAHgrXcHocpUY/g1XB6ObyemB6pdBr3OHDXK90cCOsca8rg00YBN1MSfKskp
+1LZrcDDZckjzgNJHM462uI5QTLeS9auq7pOroRYGVR7rfYDFSsnjUtS/TZIBI3h
Bzgl5D5SSYsTfnS+UFCLLlbbcNp/EJ2PYs0+HYqCvO0tHkwDj7wTy0udOiL+xZ1q
jLmr2xdyDd+kd7lLvIsGPvYSBsIBaNvojr+GiskgvYd2GT2EGOeAJ/8KwTm3W8M9
RsOWmi0yfjXNxXuaZazxEz0kdZcJCjCOlbXCNTf5vdYSoed34HilJV+OWMjxefUt
gcrvuWoSt57ZJxrzFVmuHQ1hMogB+v1zMRzPNASpIb3Uifi1bxLTAwslZXUOVuTF
2a1BD4GrZjwVcFstrGS/2kL/ZOgvFe0dgrV10Iqy4nxBcRMPBv4uR8jcA+HtbvIV
fE6wIchwjVg4DCmpTZczDmN93WccCoQUYnQ6G7YSp2MtEy+x3/UiTgEhBDIi1Tgk
v5CLy1kbs++m6S67ZcgDXS/r407eo2ouPztvlm2mGAVFc+oJJlaXWKqUkG2io1ho
pOpiX//hOrMIb2tTP28Ofl6Ln277VWnI/U+qvac4TUB+OIRr6+RvNVR66SSEZ88O
mEl2XGykHdHItJs+nOcMjnE2uAnYqLRrYlp2YTWpIiPIeTtZCn+xDyTRCT4Vr1W4
/1X+s/yEqE8snkDDhrmYX01P/B1zVRjEZ12hWhgSh0dkKNHWWK6jcO3p1seRIxxn
80zVBfznYnOpiv8FQX4/xAwnNBXCEz2LO5mJgwo412E2/7oy9w9QX21b1WjI32PY
xVr/QQxHi2L4XQpSZ0T99awKR7DtsiFnGUcyBt9SqboX28W0x5k7Yp8zjmo+s986
5WkHDxZtgaZX+KRvrzlSiF6WX/J3ZlIT53X5YgmCRf/TfAY+h5jWDRyOUQOg+6jo
xQ6p1TazgkjAOiFvWf6lJnte4kc4avyHUBPSC68/752xFEb9eKiqCN2ySO3qNqAS
IHmQdtPYiLM9n5y9ZLqivdZTGj+vfxW7vjGdg3fjCtU0sEi2GY0YqVH8olajJjW7
PWU4BwXo76HUZWgbhq5FGaqqTesGZzUz1Z2wzCkAPkdIoZxz2ZkbRimCLs7f68aA
sqWC6Dv2Gi+SCbNmyiUFgm9oorC5bwkv1UOqHoeXHagLHKqsX9WzHqdSZV8eipVJ
nPk2GFwqNuk8cwV7L/spNse2gRBwbzP8U3/8J7usKGBsC4FTi8232Dup1di/+3eF
OZthL6HO+bW53L5NyNyYXyTfobL6dbMvfLpUfBDuyGLStM67GwLqEDUL8C9h+AgR
MK/jb41xbPYx2mP7U2mptk3j6BgEWkgut6ajdyXJNUCNzBC6gb1XMwITy+6UiGKU
77omjsyTa64DhGUJKMUglfafWBq2E190XhC/NVhCcZjM2dG/8p3PW38j3xIVYHMF
YaGXAOE3yJrach+9dpUGxvSSaC1XqwJbKRYcnUv1Wz1v9DqzAHVyzZRDwTXPyhnL
KDvNyefnjiK4+BqBNxE4DvvlTFkyR49eM0inK1Nrsq1cfB9YvlEA93vQDDRXElqY
d5ngMdcCLtuyQz3ySTon1PL/46NY0oIu+5H11EsgplwooARuzOzVd05PN4Rsh+l0
J31eOvclVqSiez+TycTozA1YgUzFbA4o53MxiGO3/reewSABM22j19THrvDmLS9Y
tJ0CydIx8DBizaElhCTwfs89n4YfoQd7COvD+fbi6PAl5c2CUP+HHPkZwEWsQU8E
EtMevEKnY5h5jDkNjKeBtb81zlbFLEuObjwyeO796YU8lFhJy8waq/iIQpFoCl2g
qB+0BCemT8TWDu328sp/6Iwmzf4sB+XXWIqfjAtjjMrjnZ9mYEymmvff/PiTY28Z
zCAxjuiITm0uI2cq5RqUurZhQEKBD9HBfkKDA6yjlyinq3fB97eFL91kK/8c3hkE
sCYqJPJt8MHV59cr/F46be9eu26etX+bAlJzVBxSckC16r+KgrNv3K0zIt2ksgW9
IbuPKGwK1RKSocNY8niH3FSJZhoMKDqKgEKjJRijJhNvwKWiBAt5I+uEVGXxC9Dn
GgOfM0noU5EcqB0F+T1q2AehT1uxgA7F25C2Ieh61Mas9YuHomC/pJ7S+qxJ78I4
ZrMdodzhBfJZv/mCi5N49NFMFdK9LX52tTF6IihlVUcL/seII5V0ziDahFVcnpLw
Pqy4w2WL3HTxGBaw7Vr/ooVaLezsaijpv2qZ0YYAPKSSiaM18dGjgEnjRPnCR/s1
ASscA/yI6861OsA924foQ9IKg5x4KvqON+EWGeuEQEa12oi3QjeJ4PnaWOosuVEs
fVZJLQO41MXEl/xVfXxTnqc4mlO4UyMyOD0C3Y+MuWnuTmRPxGn2i/DvHwjixq9h
o3qbnG+y/SXCoYsLjPHjVpq+O+cs1cHNeXTmN9nmcM2o/RW5kTJCF58R0A6MZlwl
X9PTI0rXvmVqZ59m/Vl94WmhUMZnHVWmfaT+sY5NZlKLpM2z4BdlZO0S+oO/aZ7U
jGsUfoyzXqoiJ3Hxney6rQlMABeORgHmeoNp/Sm0RTM4SIpBP/rDhsvSFCvE9cxx
eC4Pc+nJzClFNQr9C1Hdr0l/VhEL6wDpH0ancIguizbgtmjSZyjxgaxa8LZ39Uot
v7e8eorVgwvOFVY2cEDjItfWy/AMt2XFf1I7KvwIjNtVJaSaSwpnKy11Fqvye1Bq
X1BPoiKG6qjDJKD/pIigWwLDv/W3DO4PagpgcCHoaV6dTKh3s7g0uCvaQw9cSMoT
Su6lDBtak0iD9bwpfP5vCJ3277Q/jmk5mWGTA9EuZeVao6/Bv+GkikbgtC+gdGVp
8Mb085m9pE23XnjgJ3QXJu8l7VMRPM5c0VvlxpqYd0vMms9y2Y0/OhP+pKxS2NU2
s90t7RJGzodCVPwSLQ3YD9TvBP4oi0mknPltpT+DpZ31mls20Q+5shRUiRgX+b4R
P9M7fNGfJSNK1OFweyqkRoQVfu/WGKk4cDWgQrQvAb28EfCuDvwPPBSGb6fnQrKH
3ry9z038imVI35rdZyTU9RVlYEz9+fZCbRxIo18EIIQ4XrkcImxKtwZzSlJD0s6i
P+2dGQlBzpK93LZAUyF90wYAaX60mHAmn8qkwLaPdLrYdqO4/zFxqYwNoGiSPhPJ
9wIjlu4edcDUqmAvSxn5vW28apIeMaMPUPZjefaDTUMF00H2xaYcYwng8q5Krxtf
NlMRUuRbnga33wF97gp3jH5+TYNmuUzbUEmYIzA/4Ti9Js5RWqxqiuNyFwo+0iWs
0FBbpRtHRGnZe2uxIAGZc7Z8LTJXD1DvR8F/TVbPcyCIzoUPb1wG84lTqAUqzxGz
T9k5mp3dGdWZmR9ZJqegKT+z1i4JPEptm5lJE4l6sOkZZLPbeUNFVsJ9yL8K57Rd
QTX/Afxbu6wONrhPzgwVF1UtIQtVpeIxNcTSmijkqSbmA1dpRSf78Y17mTNP2PD6
XfNLskQ99K+TqDqNcuKS6Edq2r2aNfRKmohwwvx2J1W48k7Gj2SJmD54S3PcOEHY
2lwDLSUBHAFuoZZaX6sZvE5TupYzVgJq9ReebA1DpU3SD2mOoMgb+pr9lEBrVJVi
FvO2jj09Bi7eYUP1NokgGEjnRceinyfaWTb4qiVHgEl5xELdG4WmDcBjrxC9NA17
c2HeD0PZJiP5x0gcMDA2uQZsGJaJOlsTOBy1Ak4OY3eYLis1zF3kkrp+JA5HujOA
1mPySOls5GXPK/mWSLWOYKgAwEommCki+FpyksDNBDq8l2d+N6NXenBqmqsUQora
o8Yi75tdCfGnaoNGL72tTvimjJV02gHTt06U0zzYvtRo/hgz7P/YO9fL92VP+pyU
vz99KeILaLqsZWrISjfwajAebYsV95zK51cDT57h7X4UOBt3Zw8BZGJEYrOP/Cuc
JMjc/KDC/lBsJYljyjvV23S58JDuK+iPVJ667mVzvnlW5aFr2LAuPvPlJ5GkKSVi
4aeLOI4XAzgb/WxnmGhAK6/WuB2rbzE/bSBh3rbAYWLCaEZ+qaEkv/P5NvJemgAr
qZwyT2mhS2bZbaL1s3DYoLTLSiSHFVe8sftwfy3BGKENBmfi6AXGzL7ql5izGIOe
IcOmES4HdHhfBav7v/JRsSg0dRYIYPfgAVdN7Rlez7purW3qdV6rjeg+g3d/usKO
9aq2oljQ8VEgANRiLeWALCY5Ga2UCYGcLh1RCnrXsjv+RDpbDID86/g6Fu9cReXH
6ymmMfyCtLhafD8EIM9bmGWgWPXSzViVYIy6S5hiX7HFpKYLdEHT3oJxkW4aBCLT
FvWwYVRBZPoHh+dd+jbBKYv3T0BqpPffajjIN89m5u5DEoFf+BNPmlvLsaEEJo54
N2qZFUJmMxRInqocQi1LDPfByS8YEMXOaqFkAYwKhrA8uCVmAygXk1o4Xl+jvt5d
QUtwWxyGfoNyg4RsuzgCB5p4/R9Kyp50iYntYLD3P7FbtXc7zgAaYAtzqruWvd2d
qnR1skTrdQTfGHJ42J8R2X1qeQMMBiZVw/w3dyKgZn+N/t3gbYr8gcf4PNtD6bw/
VwoMCAQCJ/CdnGaw/8cJ9JMtUlW84qflRGnNjKWVCxqzEW+FGIpTR9WEaxUvlHsM
4ROWRp0zkO6ft6g2JR74SrOcmNcr4gTlBjOjKkOxgCHvM3ZMMLzdaVe/UWZKEEfo
OS3KsapqswvTWnDLdNQQUcD3g+dlW4AHcPQT314ZGcCMayB5tThCSop7eliMNcZp
T6k2gz0C/dq3f0xvAUORoSeimC9u77mveVwKrzOCvPc8cYFNqQ+9cgZ0od4YWnPM
IgK8P9cAwXNkFef+tfKpWH4ysLQ/oGm/GmPnx/hLsoQuTFFc/DcQqv7d4sNc3S3v
h7jnm3k39qo5EKz24wOnC1o1CDnZcCeT2bGmYyF0Kym71quUF9rHzykMa8YQRJku
J/Zk0j9SdhNsDW3thfAEfJvkxP8EAqDLXeLn1W2bdbHb1pan4vUmdi7liSmF+zbN
jvj+M8qw1Xp5BIYDg+WVoMwgemH1qesmFaUPv2HWKYSXrK+v/MP7dfMtOVGIINvt
EDRDETn/Di9jGPS2g/ExdoskvItFChc6h0hGrCDI7f1b7jpdTIKlpuKGEumPAU25
Wc/MA05Anvfk4Ux0FhAdip4c54aPR6GvF4L/W+6Pe8TcERvJx0ZbwbUDdE8Aljyj
qgt43g7a4QhWlE/NHAy4MJM8FWh4iOqySnmVJAiGJGPu8gv+yrvD+FymPnt6n+78
Y9l4ZuKdgEE9OVADIkNR7QAEPCPWZed/KysurUYIGmtJo8b7AOMeUopmH0nMBFw0
mzYztaKeK4G2I4/IE973g8o9LJBvfVmYswkuk3keCR1gIHq7M15ha6ylOZDJbmS6
TCDmUWtHreHJCMeErXcCt5de/ay9EkUINonmZ/9omDqOlhRrzbfQMj98v9jY+IOO
99yN4vsSDcn4q6riqbcWbAZOufR6imAic/aVD+AN+x+jD0a8wXlYxR+UGA6A87ib
joDQctke0h7sl5RxROnEcsdYjjNuHJ9j9sTbqAxpQtp7s5VQmh+r574N8M521VCG
PmGEBamwxS3jWwgt5QluMPsMpKKSfJNOBNA1aQg0Ht8oSA8rAGLbPBAyXYWJaqlA
f3OORmidM3xk6PrJEcBm856f3o1ByLV9/xhndMRDJjTzsSx8gEUShhV9R1cTUFHi
RyvKnn46p80ivvJkOHpctcjkKSdAARhv4I3qW4O5+VefjL2YnqQunc9ilGQPPKGB
VJREOU+5nwubrkvhC2aaXZlYYS/4yXZ90b8JOQqJ1WIVjYutQNJF904FyaW+hhor
wvPhb9oun406Q4oMh0kwc5gT1llMwSbaRazJAi1mR8eqhUhf3s6YKQfasQJFFkpT
DEYDwRUpfMKXa8BK/z9FDchD4MqQDK05USVhDWlzjrbw3NZBDHMmgyY+EYxvtjj0
DbYJUeuj/ic82cfYHScnlrKu3tF3/8aP5vnjzi6divtlXZr/G8o5J0GV7wNBGGrX
TDI3IgwC9LuKA6SEx36J5uCYW3aPyXZkHDzeWGin/9Z7Y7wiE5o8fZLfUcuIlzYT
lRLtCOJcU2f0/UXKL3HlcNF4+vyx03njVUM9OFu8ApmtW5ITj215NpR1d0NSTk3G
yCNs4lzBPXqYqJ0iFchdB+GuHaG3fF5kAUc+6plk4DtKfv/D+tiQ2cWOqGccbPLT
SUinguLCxb+3O+svYWIxFoOCENH6LrlJUbmI52OkIUR+PW2IeOOzQOwdez2FQAwG
OdA6yug5ncL+RuTklQSW4S5IMa6vtEzpYRV8ci6DHc658D+1gRegvj0Y1OBxpywj
9JDl7x3NPLWloKmwOdmVqV8te5Ta9/Ze1HrlvdJ3O9V80Tsag4AAC14gzjhQlNmk
4xpeRO+aA1XMZ/cEfv66TkhGfB8ksUTwWyp17zx0t/lgRGzCRidykn+6f2u5a28n
OAK/PKjrR9IjDn40XgdVQBwl+uNxlLOdkj3ak9FdENGIxn2pCVTASOmROIhXMKgc
OOVhU85n5vdEFoVkAMElstCBPlu9wyMrzsvmaobZQP7gc3AYB02xkKg0WDyHT40L
SkFIfJHPRztte8rtb+MVsVotNAO4LXHCNcRcEAlkF+rnNrgiCci/2yE9rUoQ+1ai
V0IhBajzGulEkEGg1R/9UuzJQvqm4yAcN0AMxC9Ebw9sQ5F68CBNs57qj0K8IzPt
c7SAO8spP3XgJPMMqwN0zxDAZFErhWXmm9/al63E6Cxuop/W5hm7Vn76n1a6IYVN
cRivr8Ks3u6oRhgTgo9FFSGYXLmdG4UvGniGt7HCTFqp1iqM3mqmX/3TiP4MxJAY
v5No0HI9RLwoagQVVVQys9pSbN3NXw6Ld30UH0dtL/UQYfljgftWCZdHs/1NxbFs
ClkBW1FjE7CElUMWzWfqQSVeAcd/M4Fv00EpQWytTMYM7DUtnCRMFi1CFstMk8R8
nA08/fQb7rKIa2dAMIXorp3KTHGt8NrwonTuNQGlOKWAod70eOPjqUCE7dtqYluD
cZbSE9SxnCdRAE6Ef/EPRAZf1JyVSbSc3BNZhJxqWs18zvd088Yjzijd5qbxaAHQ
Tmt7y/jEtenf4uiPHPnzKpzUqLwKB1wqmb/owyFBRU32Rf8J1fTFcUSQuxNrY41u
RGg7c1JhRI67suu6v6XfSDfGYiVW0SfhFs0kOi2PB6OneGSf4p6yBjtk6L1rya93
l0wobpmrDjaEnN4GJV87ynS/6F1upXDzVXovGOTxDnHTGrKmrvtGe1W6JgENo6/v
eFztt7JKIqAsM0Uxwjn5gYgLw3lp/0ioprY4PTPw/fkSUtQ8q8w41gfHJ+KMEqMB
rvcrumRAg6LN6kq7+R/+qUYhWAZknW4TDKXfe4WkljQBvhMOtrq0IVxyDyDyGnVH
VCy4OEn1UyYthQJtLeHtQnazpE7Wk/2Rwzl+8EmjOeWLGkZF7UkVRVhxdeFJ5w4r
p8ZAy73yXrX6bwQ0SedZafCdc3ubv5q5bgYjPkX79DU=
`pragma protect end_protected
