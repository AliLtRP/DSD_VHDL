// (C) 2001-2013 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License Subscription 
// Agreement, Altera MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the applicable 
// agreement for further details.



`timescale 1 ps / 1 ps

module frb_timing_lut (
  trn_clk,
  trn_reset,

  // control interface
  timing_std,
  timing_lut_addr,
  timing_lut_we,
  timing_lut_data_in,
  timing_lut_data_out,

  // video parameters out
  h_limit,
  h_sav,
  v_limit,
  v1_start,
  v1_end,
  v2_start,
  v2_end,
  f1_start,
  f2_start);

  parameter G_SIMULATION = 0;

  `include "src_common/frb_include_smpte352m.v"

  input trn_clk;
  input trn_reset;

  // control interface
  input [31:0] timing_std;
  input [9:0] timing_lut_addr;
  input timing_lut_we;
  input [31:0] timing_lut_data_in;
  output [31:0] timing_lut_data_out;
  wire [31:0] timing_lut_data_out;

  // video parameters out
  output [14:0] h_limit;
  reg [14:0] h_limit;
  output [14:0] h_sav;
  reg [14:0] h_sav;
  output [10:0] v_limit;
  reg [10:0] v_limit;
  output [10:0] v1_start;
  reg [10:0] v1_start;
  output [10:0] v1_end;
  reg [10:0] v1_end;
  output [10:0] v2_start;
  reg [10:0] v2_start;
  output [10:0] v2_end;
  reg [10:0] v2_end;
  output [10:0] f1_start;
  reg [10:0] f1_start;
  output [10:0] f2_start;
  reg [10:0] f2_start;

  wire logic0;
  wire logic1;
  wire [3:0] vector4_0;
  //wire [31:0] vector32_0;
  wire timing_interlace;
  reg [7:0] read_std;
  reg [7:0] read_std_d1;
  reg read_update;
  reg [2:0] read_count;
  wire [9:0] read_addr;
  wire [31:0] read_data_early;
  reg [31:0] read_data;

//------------------------------------------------------------------------------
//MODULE BODY
//------------------------------------------------------------------------------

  assign logic0 = 1'b0;
  assign logic1 = 1'b1;
  assign vector4_0 = {4{1'b0}};
  //assign vector32_0 = {32{1'b0}};

  //---------------------------------------------------------------------------
  // Allow CPU to overwrite RAM data
  //---------------------------------------------------------------------------
  //picture_rate(0) only selects between 74.25 and 74.17 rates for which values are the same
  //address = interface(3 DOWNTO 0) & interlace & picture_rate(3 DOWNTO 1)
  assign timing_interlace = ((timing_std[27:24] == `C_INTERFACE_1080_1G5 || 
                              timing_std[27:24] == `C_INTERFACE_1080_1G5_DL ||
                              timing_std[27:24] == `C_INTERFACE_1080_3G ||
                              timing_std[27:24] == `C_INTERFACE_DL_3G ||                                           
                              timing_std[27:24] == `C_INTERFACE_1080_3G_DS ||                                           
                              timing_std[27:24] == `C_INTERFACE_IPT)) ? timing_std[23] : timing_std[22];

  always @(posedge trn_clk)
  begin
    begin
      read_std <= {timing_std[27:24] , timing_interlace , timing_std[19:17]};
      read_std_d1 <= read_std;
    end
  end

  always @(posedge trn_clk)
  begin
    begin
      if (trn_reset == 1'b1) begin
        read_update <= 1'b0;
      end else if (read_std != read_std_d1 || timing_lut_we == 1'b1) begin
        read_update <= 1'b1;
      end else begin
        read_update <= 1'b0;
      end
    end
  end

  always @(posedge trn_clk)
  begin
    begin
      if (trn_reset == 1'b1) begin
        read_count <= {3{1'b0}};
      end else begin
        if (read_update == 1'b1) begin
          read_count <= {3{1'b0}};
        end else if (read_count != 3'b111) begin
          read_count <= read_count + 3'd1;
        end
      end
    end
  end

  assign read_addr = {read_std , read_count[1:0]};

  //---------------------------------------------------------------------------
  // Instantiate the LUT
  //---------------------------------------------------------------------------

  frb_timing_lut_ram #(
    .INIT_00                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    //486i59 & 576i50            |       |       |       |       |       |
    .INIT_09                 (256'h00000010A0080048D9080288342206B30000001390029C0A813702E9C42386BF),
    .INIT_0A                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    //720p29/30 & 720p25         |       |       |       |       |       |
    .INIT_25                 (256'h0000007FF003FFFFFAEA034BB9F819C70000007FF003FFFFFAEA034BBA9D1EEF),
    //720p59/60 & 720p50         |       |       |       |       |       |
    .INIT_26                 (256'h0000007FF003FFFFFAEA034BB85B8CE30000007FF003FFFFFAEA034BB8AE0F77),
    .INIT_27                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    //1080sf23/24
    .INIT_28                 (256'h0000002340031912423102B194CE957B00000000000000000000000000000000),
    //1080i59/60 & 1080i50       |       |       |       |       |       |
    .INIT_29                 (256'h0000002340031912423102B19445112F0000002340031912423102B194B3149F),
    .INIT_2A                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    //1080p23/24
    .INIT_2C                 (256'h0000007FF003FFFFFC62055194CE957B00000000000000000000000000000000),
    //1080p29/30 & 1080p25       |       |       |       |       |       |
    .INIT_2D                 (256'h0000007FF003FFFFFC6205519445112F0000007FF003FFFFFC62055194B3149F),
    .INIT_2E                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    //3GA 1080p59/60 & 1080p50   |       |       |       |       |       |
    .INIT_4E                 (256'h0000007FF003FFFFFC6205519445112F0000007FF003FFFFFC62055194B3149F),
    .INIT_4F                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    //3GB 1080i59/60 & 1080i50   |       |       |       |       |       |
    .INIT_51                 (256'h0000002340031912423102B19445112F0000002340031912423102B194B3149F),
    .INIT_52                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    //3GB DS 720p59/60 & 720p50  |       |       |       |       |       |
    .INIT_5E                 (256'h0000007FF003FFFFFAEA034BB85B8CE30000007FF003FFFFFAEA034BB8AE0F77),
    .INIT_5F                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E                 (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F                 (256'h0000000000000000000000000000000000000000000000000000000000000000),

    .INITP_00                (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01                (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02                (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03                (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04                (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05                (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06                (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07                (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_08                (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_09                (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0A                (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0B                (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0C                (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0D                (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0E                (256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0F                (256'h0000000000000000000000000000000000000000000000000000000000000000))
  u_ram(
    .CLK                     (trn_clk),
    .SSR                     (logic0),
    .ADDRA                   (timing_lut_addr),
    .EN                      (logic1),
    .WEA                     (timing_lut_we),
    .DIA                     (timing_lut_data_in),
    .DIPA                    (vector4_0),
    .DOA                     (timing_lut_data_out),
    .DOPA                    (),

    .ADDRB                   (read_addr),
    .DOB                     (read_data_early),
    .DOPB                    ());

  always @(posedge trn_clk)
  begin
    begin
      read_data <= read_data_early;
    end
  end

  // packed as
  // word0 = v_limit(5 DOWNTO 0) & h_sav(12 DOWNTO 0) & h_limit(12 DOWNTO 0)
  // word1 = v2_start(4 DOWNTO 0) & v1_end(10 DOWNTO 0)& v1_start(10 DOWNTO 0) & v_limit(10 DOWNTO 6)
  // word2 = f2_start(3 DOWNTO 0) & f1_start(10 DOWNTO 0) & v2_end(10 DOWNTO 0) & v2_start(10 DOWNTO 5)
  // word3 = rsvd(24 DOWNTO 0) & f2_start(10 DOWNTO 4)

  //---------------------------------------------------------------------------
  // Register the LUT output
  //---------------------------------------------------------------------------
  always @(posedge trn_clk)
  begin
    begin
      if (trn_reset == 1'b1) begin
        h_limit <= ((15'd2200 * 15'd2) - 15'd1);
        h_sav <= (15'd276 * 15'd2);
        v_limit <= 1125;
        v1_start <= 21;
        v1_end <= 561;
        v2_start <= 584;
        v2_end <= 1124;
        f1_start <= 1;
        f2_start <= 564;
      end else begin
        if (read_count == 3'b010) begin
          h_limit <= {2'b00 , read_data[12:0]};
          h_sav <= {2'b00 , read_data[25:13]};
          v_limit[5:0] <= read_data[31:26];
        end
        if (read_count == 3'b011) begin
          v_limit[10:6] <= read_data[4:0];
          v1_start <= read_data[15:5];
          v1_end <= read_data[26:16];
          v2_start[4:0] <= read_data[31:27];
        end
        if (read_count == 3'b100) begin
          v2_start[10:5] <= read_data[5:0];
          v2_end <= read_data[16:6];
          f1_start <= read_data[27:17];
          f2_start[3:0] <= read_data[31:28];
        end
        if (read_count == 3'b101) begin
          f2_start[10:4] <= read_data[6:0];
        end
      end

    end
  end

endmodule
