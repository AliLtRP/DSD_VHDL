// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:13 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JoSssmQEySzzJmMbB58yO/OlM4GiloQQt0Ehc1MWwQzlnLtLA5O3U4mOMPTrF7XZ
XsKbH4gScDydlRVgBAqztkzrz33FwMB0YMtFbU+vAf6l5J+kFT/pUWEJ8FKjta11
ChjG/tfesyH+94NnDzUX/llrP50F4bwLWH03BbtX3QM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11520)
igfXlJt2qYpUUHWxM42RYanwOaRG/VN1CP6ktxBHwv28n0aHH8X+yMo92PSPIulL
ur6Jn6oIJnLIYDOw8k1B+Odwj4xGTt+Y25QYATO4OcyaJTFjaJ6b0fpet2qyNpQ3
P5cr/w2jnS/nmShmaORk5ln251it9eZBUBe8RICOT7roZvOUhSYazpuXf1TC0fL9
oyevYo6HRu9xW9QvwyRhGUONOwsooGPZr4nh4HpFXtplh0TLOgW1pQBiCIwrkjXw
ekTUsnXDT13aMRWbqeu2zvQKtBoLjOEdJsoMLp6yYTChQnIfyufeJW+u4d5ZRNB5
ejADv4mbND0Zn4OquYG9sjA6GHtoXYvCRlsUpWywzPjCobQ+cV653xb5goMWqyxY
DT2ZWW6ySXG5y0nN1Zk4Bt1x43adFmRd93W7bIxVT9nwietz8Caks2bqu4dLuExD
OeSbVLzEEpqf0I/1fi3/5MpyRmyJ1vE3nt/iaADVKwcGHQwPINqGsgQ9Icmejj8z
Zck+LvdzlSaDO3aBTt9aeFgtf0xweUeKGrpXzftuylsRRJMR/bMkQyAwLsNCk53R
75SPvXDhNywjsTxNLDsfgX3aLdeUaCUmBPVkJYsGUVlvcD+X6QsAMhFmKn9t03a2
zmqBeaLcB9dQzAidF3ZWwcp12sidys/DkXs33ZjW7AmJdKhd84t+lj2hp3JabhQI
SrkiZ+YHrb0BCUJvMIoLCsFbL89Zdxx3VtCnDU/xhsTo6Uzgy6QDXsGT3tu/tCAO
d9Za3Av8tba0UZvccbmH0qHEPINOj4dE8D0BPVwWOn4+ORSngj5pb6U+EjMEjRBT
VPfP3U2ZiQhj/56V0239Wx+jLMSoE1cYIznyOa9+PeZ+9P4PZJn4a399+/kGwSct
s2SmiqzuURA/L6xGDSJkJ0bExyOJAPZA0DmJ1gtggBvH5RnSSntD1XHqtrmUIxRB
WOZUloEkolklaOQhGSIxCdH/gPPL/9IrtATLRgXWzkilBvGCANdFjeZeKtKt4fT+
nmEkUF9ZGchGDDH/LnCVS2e2Bnoq200/WFr6mErj1+DEA8dztY7fulyKHe42dkrk
HgTQ58Uvca0UVI8lFgDP7Niv7Y/NYQ0ThdWmoL4l95DUB8w66aQ8xMYCEKNt7Y2M
5OTaVSEKoiDk+jz4iH0HLdOunGb++x/CaafqOcXA0H+3IVR+cQwL67aAJOvJOIBd
vOTVMyBFk1fB6QizzZZS9IhLtSZagisRyT+YhntwkZEubjy/uCOBol+Lr61HWDbq
g8Mwyn/LjAacoz53pYCzII1aR+QvukA1pPC/WXY3l73yogxujQfaLFNWWQ8FYpxu
f8pWSgaxC7fTZVekCZdyuG+x0c/Z/APd21RgxLNpY5MK+K/7ahzM7tJtVdmsCZF0
lnI9i/x3YxoMkPbLO5jz5FFbzGr5oI5K3lGBLyZHXEOXM4morJ/hrzw/rUnhgCtN
HUOGotaYzJgPkpvzmusjtEe7xAeD/F7dPPM7512KTzj++pxTuiw4TzXjVOf0raww
mwck7v/8lkj9l9hdwewnItRBoEp8tJsIOpEMkjiDhQYvdphxeU64Emymi9ZM4hsu
Tpkqek6Hc9gH0NE+aBDBeUdW7F3dVlkpZAzTR61IsG9pCeI/QsKKFDj2lBGk3RHd
TR6pqms4qaQ635WRWy/zaiDkt1iwXTlhKV1a7wzb06fvymSrWzLLfUK8YV85R0+2
5i+rfz3WeFxWTRHSD02yDhJD/TpFjpfHfm558ZiKBg0l6v7x7yAPqgF/IQduzueU
PkcCQwFKbd4mcJqGWfHn0q1AFebf/e4e4xADHp4x/QkfBxLnjVVEBeqXikS1ZMo/
rg9xEA9acekgUiMoBddL0SNO2izqZgffRhUaj8PhTDDoAnx7kZCXsRbSpq9cmh/R
9RO15fDHDbCatsEGgT6kxE2RJmbAzaBQMRWBnW7B9CU2+lahqnr/RbErEt8Iv/YB
P6blhbTBVV1ftFWvW9atirDSflLQDhehkTzdV1kkVgQpVm/kT4DE4Z5GUxvUEN77
+9dW7HoTdEFtK1Q2DBuwP0ORPEHDkjXwudCeieQipMPvdLHTOGSnwohrEDl0IHRK
WWPLKz3erq5Qj6FLuqrTaqYbMHKTayD41HJ3Ux3gXQPkcWDrCCGkVvAdznes/FG9
kmwYMX1eqfHsJ5KcOaJrLyZlEIsaTPHvJVtKQenaUpbSJztOv3swGuhEkS+giJN+
x6qZJqw80Dr3EcRAqg7vP2rPG8T5SRUUtVfAJJMKjNX6BWuj/wtNk92pwS8wCjr2
6r6EaEs5H7cn0fcpwJkGGH2Ua7eMfD2FaZaymd1XNwyBx+UVTwLGJxcVNU72yGLd
phqGPUj6saAzb6+dNcpmpyLJqTMKA5XNZKu8/cUX7vjoCHNpoWb4mmzYnzr1SV10
b/nTcRLzm2StBxY7OXRTnu9FjCmKnq7w5T+PwYPGyM9bffpz+nEoMAoq9meZWlhY
nwRPaDQeS5B6NkgbfuyUk7zr4suUEYh5j1JCyjJbMawVyPfwJroHd0yHwKVNVD3j
KaMZJNZPeg5rV+6SSxLmWjUbuivPeSSVlhCgWjPaIrd8OUGVXpR7NKHzL9ET3RpI
1fXtJcOlLyPESe9hAYJQ41UJN7EsQPinng5cVq04+N2a4UwKe2LJexGN2+d71HEL
o1lmGgNVR4WzDwszBxA7HzWGGsoqM41cnohmar51HKMoafKTgvi1f8EK7smxCSQu
Dn/wgzUAilYdkzNLFpfGdtGd5tTEgeEi9B1HjaB/kvKJ3jNjmQXqb3DWA+ZTeLZB
Yj+wtSNL5XzFsiMcmKaflfuEX9iVsZP58oSGSujIVt98LYKI6BPp2s/70MKW5HkS
ebUkEthowHRi6Bc+4ulNI0iU5tvhH/tFivK9lo5wShcIHm4wX9tT9/8yEuZvSX+i
8qJ+qy2ust3OitUu+Vtjj3k2hQ4V9WrN0z9JlOwHvnVyYwm9SGkiDmepZuTu+8QM
ZPq5J+V0XwkBzCvqOc2Lz4AlYZK3NlIuOZS3Pjlexdng405QZ6JDAhXY2toHXrsZ
yS7Dm+rlc2UpRK8IZJlixrRURng2/v+MoiDvm272ol9ROr9u6O2IhImUCpL6szuY
vwIhAC7+jFwj9+Libx255jNIqdMSqw7hiiA0YrAVxZTnhg5qCXasxbne5Y2dlEhM
2XzrNW+SLPqlA30DITD54xwMscbyLUI+qXV2IAsP3Vi/d9GCv4TeKviHPqWXbIFb
YHAX/MQaT2XYEMghir5e5rSbd3hNA0Plf/v7oV47FfI2WhU3lHcY7bLY+63apcN2
Sji6R/ES2Ju1oqP3rCtZ+fmYh0Di54LOGq62U+jCqRoi9SD3RBZn+QRwAnGyU4yw
lXL3RV1Vm71ttj1JeEJkUuFXKGaoR74CJBa9IF6swO9Hz4sNV23g/TujO9/kzj7V
LMk9wZResz5SrC6li5eBE7630zYjXsWr1HEKdZg8HDZLcASgTw3N8KAi4llvvTAx
2nCCreggwEOTHUDodk2TK0mFn/SrXL+UuLsgHuUc0hs/lkKnZGMJTcDkH2fGoOuw
PKJKx5hGnTqi9ZhLaChyGfqCNzGvoTIEtvI8m9GI3fxJPrl14unm2O6DZz2fATCU
kv3bKucgjh6mjvvCyaQ1zhRY5IDuqNEWi0E0mZdYy9BdTpz8fCwk9Nw/KQacfd3j
6RPi1fYzEePrp8lPvjcVXOLWP2Fca+Suj5pskoAwIbmY/2j77GGiBpV+kAPu161+
+Hjsy0QSlSoOpmbi4B0lyFUUVznD2m4OhiUHeqekhgjPlzdm+Qj0cIuEr0U+xwlB
tEXKWG4Qo5ct8Z3JaTs9Ysj9wCEAGPp/bBqyQmqffomsmoUiNMSMlbDew7FF25oJ
1MLUMAxPpIEGfR3PmVfUW2Z8CBoDwNIcbeY5YLab3OHF1yHTLMsR4SPAM92gzn8v
8QVQ83ILPnoYGxrRZSvh6ax7m6TjYq4KMbfSPmv8h2gqzn1/EADQKG58vC+wVH2w
T9FjLg44c13IMUYBqkNz3bMprtAua7HXe654mocptROeu8/G0l0JkZpnR6pfG8C+
qw94QSlqa+ft06NqmAbFfPhexKGPImaZrZ1ZAGxAqXDPrS2qr5FkB8EG3Qk8PzHt
KHfpH73a3ZFtefQIh8ycm/VujwhFe3tiF/b/BlFFQ3geO3Sk3i+TBIYkhe5Jjka6
mDNixwuWS39xab42pRqGbRAE9bwxc7pDcAy3Q48rbGtUELgFA8kabcgzRcdQe2cN
eZtOQJ5Ab7rlelJCujJgP+YP3uYgTRbC/g0hKQuAi+F90hXjJ61VWztjZJc4vwQv
2q9YtcKG5o5jfJaWUgRxsLq6yjUkyEzrCjpvce9NdpzCTLOWHKuk3nSYs20/osrL
PwNJt1VobAKnvO8rJoou8xJ6yyOW6jrF50vOfw+UyN3OIaJyGJpxL6lrX66d4Gc8
MA2mNgDRQOsFurqLNOzO0Y/v4SN225+pPGPl/6pqmkkwNd/i5e4QToBytFy7AnM+
p53VfW7H43XYHqQwL+hJbz144H0cqCX0hoMksLC4OPKoH/Se75rcr9ED83hACRQ2
c/yBKhiA83VLzUkh5uNP9lSkP9RPdSuW2XUlvXjAbv/vVdJ4k35Od1eGYEqBcQUy
zMLma2t5t95No9TVT0M+MONBMzjqvHT44wnEVBdz5zpzIHB3moCVfGxp7cj6McrR
6s4Wg2SMIdABnstndaIjZ1CiWLZMymnf8N32mXQgGJlnGHIQxlx6hDr1O47eQkxh
yaqMrDuUq2jXsaGewLo5SgS47eUKx+oqzbtfTo2R14w1ApGiAZaw7RZXWP94rV8e
TGSUtDP/Y7mxTdfCgbo7BBBi269L2HL/KUVpEp+FiOskWAkj17aWJsaSeazwhfkJ
OlHcPrlBIBr7nTZIOPmXZShRc7EvDMgJzm1mMH8fMPfPG5hukin8kza+vPo31Fnr
IheE0xn5n1I7zkmkP2QPymoakM7PEzNwut6pejn8DkInpbgQr/VxXOTvsrCUacLW
hPHzhM6AILMiOmAe4AnieO1+qYf7Iju6P14curLychgevicD5F/8jIssCej2DvdX
oYKCoNCtd4H0AL/LP8YprtPh6dRP9E5gWGhxmkZBZJDfiZMWcW3hpfR9w1tCSBID
C2ASdIkZmQPMj+QA3KkzxcbePgLuh+hOpicmlqMnyEttDAtsNnf523D6cFlQ4a8n
1vphBST9GggHpiFl4yG5ypKeDtNCztHnCzCwFdCUpAp7moQJwM60JTmfx5yZf2KH
MekvAcXbJa+2TxF08rXN5DF5A1YrPcfgxjVtVEqZKTTVigvKptMcCxgc7RJ+ZoZl
h+Pv1QkeK500VLniWRf5k/BJfd6ZdfLq3OeybzlNFFlIu4rgyT6Kq2Hh9FAIdNpy
zJ5ykUYHDQffyHwkwwMNrZWM7DqIZRYs/ogJ5W19Z7WZJOHPU2m5OU4E/OeGUzpR
NDjvCv3JB1brWCaeY2IdJIYOd59JuaBroB63+PYwdbZoALGSGnARdAukBCrads9p
ucaH9hvHFjmfPQ9zPWRp7gcyTxWUOQJb80tHQpWaR5TrBk4DHlxuxKybuGRjv2Am
Ur+MkfUrvHVM5SBSOr89vHjmzjiG6cgOd9O7zse/nLP8MTxeBYm9TuOt0f0DGRFI
UoKoeKeY+8x3eGsQfnhc666VF/rTtHGMsYbF8aYCgyuWMvm+ftXQT3uV4Pc1CrJi
txFimc4CekKH9XlIMg5X1v9fBPIAQZNwDF4g3kMYESVItAjIS5b9w5+PVp04iKt6
I+e61nBifoTSzdFClZ7Glr3L21WDsuwSYbCmbYOBR/kupQ3/ThOeAg4NNwPwzkr7
XFvzpHj00njWFx4Tr2/cMPDpzvOA7WdZyZtKkbqfDpVuF17kN6MTouzVa+NmpCsW
kHp+xE7KBE1cN0NEuxYQLPsM/TvrIfHCcWXz0Zj3C68AFUfmN5+4RTevZY0MPge2
tTg8yvYBb6bkZelxuZECRHrf2TeO1KGWJ7Oj7Xv0IrhXZ/LGxxMAgXCF6xKte5KS
7WFxYthlZvw4qn5KV2Lla3uJltkQPl6dd0BheAyJI0jtqb9JysXnbA+mO+OWWxPo
HDfRMwSfXzGiyyD/LFBFkybvCBYL9pxaoY7nVRBjLX+CPKBJN4dlbCIhm2+AZsKv
uaZW7rOdbB+v4uTvNCvuLdwSNOUmJj9++OSJoiasF97z/ETst7mH/pX9yoBfuDSt
g4UpmoynAMvK23K1F1sDxeKky/e8qQWSGks55j+8ptrXECKUoOzClPBuO/S8KTrT
AmQ9Y7XOX3BiPn/4NGbHX4u3AH/WXRfIunKH/2fN0hDMNDjUSpgFRS+4z+cEF1zL
2XXbopeuKVak267jdxAErMUhb1ervEsdYoK5xKsKvi5fC58ria4UjBXjpWfcevYo
bWudIqlyaW3VD615PTXHIz1peq0iPrK9AzuOAJuGeuOZkZ1uKS8eWqyZIOShPH1Y
U9kYD6pyQTofQuy6xwkIeNLALwItOBR1jxZAgYDGH3C5VB/+LQP9vAMqPU4MsB4N
Mm2yLkQb/vD9PvZKzCnlGNL8gJjmYA+5IG6efGSSkb0zNtqLZmwP7AIfVa2tr9aU
TNqQgmTYu4fycbxn04E0yPCvEWi4COvncqmaxbaQCswcI8zyV5a6KsboJ9MKPst+
1gH/vP2a06hzpErGxAJUnnmpkOkRRM7NLkQ+j6qOVvEvI++NJSiwnbocp6EuIWqr
faGmrNtznq5eUdLBcawS186aPi9/wQd6mSGvcwAyU87/9kdESQUAsesOlr2q0NcA
8DGkMxxs8mA6G7vlxuj0SRdrW1VlUGU5/dNv9/A4YPqDv6diddLXQiNzGR2bm5ek
vKnu2eYF065/1iioxODIBxFoQXdnfct+N+DVlfQHlJVJtnWrwDRYKKv64xTdFBuL
64C7Ib+/tr5iZWqwoNubFQ3uXb7asaB6BX3srcgbnVYBPskGg3aLg1TaEzL7W/le
VOQUaleVOxj6J7q2ts5y1ClTox+h4ASzus5DrEpuz6yQVeB9TxDXIaz7dVcvw+Xc
7v4GAelaTf4LTCFAVIpyjdWtPuF9wcoatUvzNoabSoeK+k3qHSldwHL1GLNhiit6
CF8njNbo7FWy/t/H3s3D99LCy+AnRcLrFyZx9uufb9C38lSSNfy2z4v5W7y7HSFG
rrqAO+2PZCM9ZVuXeVNG8SxjcDR8z5jUFcwCwyEHf1V2i5RM+EpPHBeY/vW5rpeb
iPO1XpMa0L8zLrkLow4BdnwCAeqmyZQw1vJPifOvDe/mk6U7ANMd99IfKEm/Bcbi
DBiMH2Yp1YoZ04lq6PSeP9k0LyOv3e2QoLkOFVJaw4tLjakkXRq3MrUEiG8NR2ZH
8eNYFZy60a+dnnOOMbLw0KlMhg3hu8FIeZ2E18pxzBWiM4vJDqGY0EYT6D/QbQ9t
j5d4Guhr4b0XZZVwXiAwGYjT1nJisE6UU4lyDnA7GuVQ6eeblAUdP+m26M10gG98
ds7MOxXRMGsGTtlXeEH8RAySfzeQuWjswhV1r8BCixGqGAVX8mS1B+bZsH9UngsV
5aO7ZBORi+Q0FYkRKoAOfq/NFZ/Zpt+k06lglUQuQs3cB8MCeHdIy40qbrHLH3Rx
7NpF7j1uqsVd2xSiX18jUmdopwvXta90PqIjkpRp1XUo2YNuRVEJfFAeM96IwNto
02Qp+GKBmYJYDTTQIgZyFIUEw96dJ0T4RvdPmx6Y7eC55hPyodMreCYEHzJI6nbZ
6wAAlOZVRdjEXFdNi/0597xMlpjZRh2c166A6rBOOngtC9hWFJKJ6b9d+Zl4Xlg0
x8aqwPT9OeMVW4mcpDdbokEXdMOYJD2vgk3VW7l/WXB9wYkqRf5N2efe+7r4mmNZ
VE/Vvz+cVWFT1/awNRwIXEnve7knfsiA2DXQOBCSWxX/ez3z3p2nK5r1ZcQlutc6
4ksTuTYy8FZidty6zZ5NvGCaF8r2q9e0XGDrhpRe85Uq0XF7Kki7S22a6ySNalVz
WU7Ej1FnwLCDa4Ya8gu7vI+NwtL3hg/YwAXpCy3cFKMpOhgm2VURreU/yuMuMgmr
/0YJQZMDubTvzDN2X0DNsGcPiPzR84kHrs86hlNcY+cmDUuPtlyU0tP5PkyG6VRp
FW6MleQqFIDcZb99AJ7/8Bvh4HRXl9PQJghmes2KQrUgWANBj446M44nB5l//4dv
aSP0Koph1v8ItPeqJ/118rS6QGam7weoOFcqFgl5wtudLeSFGRBLYl0yZhhl14Cg
iYYPhZ+g5Ay2gGsxw1ya/C8jZqTFSFB6y8wIJCBSYhpnGAwcyQWF7txdf7W3BN/Y
IbuqAYJITQAZrBsx87oufYtKlXgtiJwfwGfHR4Q9OftSNAfhSgzxZIv6JV6Ig6of
KcnLO98l9pgcdTDunhdWAQ8CBG6UlyykaxS9iKIv8blbpckDM9rmdzqBcx3PeDvK
UXG7VMbh5XqcqwuTfolxU2jX4ST1jv3NaeTVPN9z0P2ro4uOlSOqo9Vd2x3wWEon
sK+y5E2QcNh+ysGigHRgSKVvWMcGX7Fc8nwfJfXi7a3oeGVTDYXYTJrggO/QQpA6
2kctzxZG6NKSInjMse4XM6eXTI0/qh4FNdGPpQDHkZN4/U27uNZ8pk2gWqnwLcvD
l/UHTt5xXTnuLspko/unsN5HcO3Vi5h4diQZtmL83nfERbv8uxpgpK88j3NG0x20
Hm26/ZMBIA7lYwQen9hulMN9mfjt4XIXcnBedp4i1oYGCGNACrqXEAfSd7N+NFLP
REf0jyw/fPHY5cT8Xga2qMMQkh6saQ5TGlkmtZvDy+yEFG63qCGsAazlpL78dacI
M6AD+XousmQAKJM4Vc8u/EtqszLIqHjXZPN0SFD4yo7nBz763abaGstXvbi8SS9j
FM4ePoZWuCAf40JLR+p0XlwACOtWyN/NvBMPVyTLxjT4dxjcWOc/cMhWS23lAizP
+FSS7m5dWkt0QvBbcNAQA4EICoUgMkqVOeo9TjAhJA1WYegjoLQznZiNzyKcy4XU
dnAl9MBeCAMGvxpwWOiec7RwhIv2O3LwaeemWBdFhPCrgiER6cI2SHdUryhoBUOY
29ZJ1G2vsqb8OqgbAjU2oJtnDjlaR67WEHOgfX01ocWBy9fKEYPcNiomyNQJLnP6
qfYQH6Jcf+gKsgQfwTnqrv9+YNTw2ihab0g10xy/VTzWYr1HfQ+gWWjO10R2VwUX
IWfNY4mHOfZkh6P/rvHllRUPH/UgXvLij6SRGauKFDcYIsWVPFU0R15lJNOTxcKC
I2szya0IvL9ekv6s3BtDhYhegJKvIjrALjupNnGAQCj0QInpC8PlD133xU8sqvmq
fT3heX/F/M6LFmHONASN7lAq4duOCIZ4sFMT9Acznz8+k42PxAzAVrZqXFf9KB7k
G/ma9KIfg9DZmGBWg/LyDEZ5PH3DoUDY1q56noPQiG66do6JEjkyx0Zvtvss1w7n
9+ppcR/9Gsy8azAsN6Wmb6kNwu1cZuG3g+qChE6qFojFXz9wInTOT+yC5oCrYfAV
UU/dA96aoBUBPtG6itrC5ds4eYDUfOFviT9GMa+3975fYeml3x4qiyJCtsm1f1SF
TpYVAqd3uiEZJkQWIns9YDTSEasJBw18o5S5kftpbA1gS9LeZF63fN3CVVunb148
BkxsZSeAhGNTpbFFe/piRe2O3T6YdXZXFpsoE54M9d6zXY374jki5HeY40eBaQew
ECnXUwsMrDWga+MHy+59ZafW2ulAHVY81cLY+mS6IIDqKE6wNPiAzhezxhFrMwBN
EaAe+fLt/UYC56b2YI2IG43vnW+5Ye2rBVNhMw5kRBhOOk9APoheRwo2FmYRki90
8fxpj39x0yC/yAwaKYy7eMX47KMKf61UDUtW8OeyezGdy9GPqzSv4PZ12Ib7M3Oe
VjzWLSeXWj2jK0eIveNW3kFA7K798v97yd3Mjv5wRzDXLEHKYDX44zGSB6s6b3ZG
p5i1YqUh93L+ANS/+qwk/PLvQ58rz6wXLwEyiQtq2Acw3z8zn00VeaXBr/vnLQoC
HrdTlwyOVyegBT2joYylP6EtrN5O6ytSVsyo4+KBMZ5SnhfF26nG4grgccrpCLpl
MrlAd8+Gj7JHzn9LV+SmBChfkmw1xpQjOnAvaVy89UJqxGJemss0O0naSVt5zpQ2
OzhGynGo5oZhMx1YTXJPYL6QxxutjXMkrjz7tVu2SpA9sHqmKjdNYWcHYLeAsdUy
BMhNBK8jN0FlD7sov8Zp6kZysTO3K6ma28hu8Q1zc6NsPUT+q4QVnEh0A0eooG9T
UK+vSUZ0+x+K+6h/hKWTqK9FYuNZeiUmPECgeD3Sbu5o5JlKewD3xiOPHJr6NLLE
fqKiPMX7IL+U3iWzOZcMA0bRT8Q7wDq2qxl0O0+a+UQEx+8oDqh7c10CoPbPxkVi
MxSk+oLHhnYGDyTJ6QRh7+vgJs5vlnX9m6QtNbygpM35JnApkdN5FSiNiFuhwQ4Q
eXVKjtI1yy5o91AN0hHCttiiCjoXGyHxikf/vLrlbMePVdClL/Hctn5thnAEigXx
Jw/pGMFCTrNA+LyDE80Muxok4XE3/SPPB9wy62jS+DrzVc92GdNgAX/GDPkDZ7YY
1LTpCxJ+vvV09ROMUMnuIfbJekIuCzkc0L5WHaNKiiT04OOfCsdpOIiQ2P6BGPUG
NcKx615B3H8132RVYEGlPeZUYwXY8R+mRYbknGaCCpUL9r1odYD3trJ9T2MucxTI
4E2mi6SAIpkHtDCzg7iE7uwGgawpMevhPaj7kc6kpO85Wi3jf2vda2yo393djWeE
1YeU3u0wfaUOPhjD3yHi/48TBL7SRtTLOkL0xJ5QKoLirNb6oQVjHA2MwwT+GjFE
VFqenBh1mrNzqr7HoUn7hu9n6ADFiYgSiUvEVhMSuzHF4/oQAW4C9UpsA+llMOXS
3l0gw/AF4y3FL35UPHZTMhkBp4W/+dcN8Uc7nwODlEc5h1ta0ykssQSdTdnWgdhk
bC0Fc7ry5AxY3MSVyLA7ffMbRU/nbl4C1evOWOROztN4JU0dfkGxncxtWwH7Y/Un
2ZZHrrOvECr/4zSYy2IujggR0+Cu3iPJPKAegk1NwC6DwHZWUscCOvOBKRS5Zs+d
IcJgn+an3aVv1Vx0DWphHptcDskDPK+cCUJ0y1OkbvnqVKKDRMuzo8FAIUsfbXIg
ed6706MxwDPoAUqQpsr2d4SQoI9lE0IDV31q11jaW3++c07yb8ukLQXVkVf1r+n7
cw95w50JMSe7cfI0DpGbw0TO5ddgeOC+iqoglsCTRA0RUqxJVDj73b8tqMKsT3kU
uMD7msZQTb2sD7McvJ79hytX7SvvVtO6Kz5xa+R3KAGYpKsYVDiKRa8rrk740J91
R/CYVPR8+PbBAhzBeJjy2hwgThZ66EsuN2CiDhn9aRDa3pKC3tRQbGVpvbx6WHzA
l6HuowAFtC8R2GkzNbK/ml6DpOGJebRfG32eaeI71r5NDnLl0PpCfoqFqNiBL/Vj
vOkpgEHbQWGQyCnDv0YhloprZvX2a7mfrLsiiWa/RBsxuvPUTaEqlf6YafkPiJLJ
7ntXYoG6lg6Q8Xu9eftYsIiKKvcHU+akZO0dCSUClUwDqWlxx20NgO6FP5sWsEJi
JM7ZTnD0t2nH4CzQq9gbm1+dAokT6jqF7HCe3FkC69uNzpCwdPN59N4rZrDbobcm
UbJX/2tAoBbv3axjzaFr6V7UdBw6JVxDFZn42HuP/VL+YthQloyboF4wQF7TGj13
3XCE5NW3NutT1/k63iexeWok13i3MSCzsOuIPsVPP1u1byH2MKCPEKiCMb8AWKUb
K62hYh0U8F12aAU7dt/Z1re2G27oZXVDNVUtz5KCdnnq4w1qsz4iZxneGW39m9FP
MYFS16SmGrSxN6fgJ30/XB/hGQNMs+GQJPkCok71vNGOqOSwL3MgYvyu3IekIXwh
wngdTC+eRI0JboFkpSSXDf/+FiR3LgItu/XGHciDG5bV3qhEa90dhyeVcnimLlFL
z6UhxmZnQDtWME9t4A2/GPP4QxInDuTtRXSkJ1NZp1sIJjBwJgymvs6lqbe/95gr
jAw10cSuCXvtSNbGMstDx92kU1xtCUZ3q5yp9wpYqbNEt1LaJYvqb40HlMtsnZ30
xTuhP1IhrReX9uZyYX0ctHXl0N6zdOGkfaE7M42JESpbgp+Cm+tryPuuKulOkTze
kkRfS7tfHHM+yAIxYz4W1I6Ka+xII4HUJN1SJjJfQth/twJt8IsatgiGO9dwRgP/
ZQ8/xl+VXjb+igv6aE32T67Y6XY/w4LPcafkwPuHhwm2Tz9umDDXU1C33La+y3Yd
PeP+rBcRatxFUIL1F7fO3AklYgnNdCxW9gJTYWzgXBPJ+/WGUApw+a8iqFlJHZUn
PUuD0jq23ns6F44Z3L0DTTaj0wYgmYUOEnagkH0lIUVtOPm9SYMTDE9c0O5gwABC
hZCNCn5zxw6AC+CTjDwfIn9DbRIuvUkxffgm62XrG/vPsUDJrvu5MtTvuATHyAop
Ia+Jo6lmrr1KW79pKgbf3X04/dfYoev+nU81SwIhncZL6cofv47PHk1D4rvE+yfO
82WU1WQFFTDxkYdWkM6QcwbxqfITUn71wwu3ERrvRDueEI5hRMEdg53Q/3CEh+R3
hlf0g+eGUMzvSMvP7LmwXRnJgpv9buFNXilMMjnI5f9XxqDRD+PIS2e/RIWggWYP
8QxIXPN7305Fj50wmQKEw8CyIGHIQLLq7PZcBBRgc4wdz91K/PfcPOnfNXCWU1EE
pLr6C0HrfljrjU+fqiXnsGEMjAJkbotLzy3Q9AluIXqbou5GG7KqBsMFVXDkgdWW
34oO4p4bvt9T8+zJgpL9AUaDo5cw4DTbti7CSmHYBFBFE8NsJtp142dgeLaU8MrW
ZuqYfCY6dvqQJ3A8s6aVYnu13bmgELGS2UbBU6EndLwHKuLSCKsINziU/PZlhmmN
JaY3JMMJB7mJ5rosYSWfPb9NHfddXpxJJfCujm5mSbi8iHx+kM9zo5mdh9T24pGk
rMCsG54yiwX21EnqB1PwgRDU99jj5+aTfvYICX2hZz8QAlQ/HWNcucP+NoeIyd7T
gFqOufyNgCmlu8jYgXLtCDua//E4v9Dn2TjlcPBnG97YClU7Qk8KLmP5evL9TFJm
yZ2sRCJn6z9md8osHOPqV7v3wDwIQhwkAnXZX+aMC4zRwMG0mVZAE6BACVwtUVlZ
WfvwWnJOzM9l/6t5HHKyHynJIdb9Jj+UB/z6E7HTMlhlPcixUtdblNVLv6pKqdVj
D+wQD/OkcZBjRlZNOSwSPVAqWXc8M2McCz4R1v5NlHaQdbycfcdLFUTrgrSrvvE/
qzpw8hvNBF3lH3vaBQcPlDbxhlT+m4wtkqTGgR5BwUxwh1gou8D65zthsbmazEui
TTZd7A/DmoSJMZ5hB4RgtPX0Lj6TIQ2V3qCwusD0J/A0jIQtYl0D6ppreZ2B8r9k
OOX5V+mf2ZruetriUzrvLmGVNxsJW3bjNtE91JI1V/Be4XYpcreUiIv4A5vZeuR6
vxSi9El0MzI/bCwmn2yLZFn7+imMb9Zbt2d5wPvMMrhs5oxQJF8e6xs+nDPWMRP0
D8IIB83R8ruJP/ZkOUl1Y3Yr72TPXe5uDwph1Lh/zZECh2+qHA1ZcBdZdxzlOQBr
ccx83ZETnnwyJz68dU7xzJN9Q5g2RU3gqWkJ4JaInRNLj17KOmdx4uC5L4Y+M+ji
DQ+Z9xfmECrNXRJKxulTttzXzcDkIibSTesGLhb9PrlsrQEzKM4u+j+xAJzkpA8x
0J6bt1U8eZzl2vBsiF+DSL4CyuHekVL3uUaHrGYZDu5lsrTQE1whaBqyEmdbiYUA
abrfonQfo7qGPnS1yUvIxFKGg/WV42Am+AmrdexySKVxhfIDn7LQZqB0Ec5vuHB6
Q4W91rhY78brbZkVb5tzYypX8L+2khYuNV3/pilELTblwo6AGtgY5GFtzSkcx8ge
eHQi9LyYNqApuPgjflYvocUftDOpemxIF08pcLPI8GEyGKoZK/eE8MB6/I4GufQE
4A4mnkcQaX4AW8boJxoE6e617mnty27wLAuPIQlTtuJn8exqviAk+v4tmCP570a6
kaVdgjkdYwmXJSC+paV5r/cCye4k8fzLt2aBvYDcWmK82n/kNMT4BMVJCZwcvpy+
kCFdjBzc9IPd/4Y1nS1j1EQbP55wjgC2ONkOELdDkbl4a6o/M/Xry82TK+NISC3Y
SpbhDV2xpluAZl1dyEiTVwYTpSSmkZw71b8SMEK69Ra1X1/yp1Hx1Sm+UdW5tPki
lVfT/FUIegD3/rBx6wbs/8pCNbqIvNkL3yL0WjQ9TQD79tgLkxLcpZyF+Y7HeYh+
yQyE7Cch9UHtgvuFHaYZW2GHhGWQ2ZZj6j5e4tdcqVepi0VGtkv2X6A6luW+oSQr
Aa09yUV1eVOoMm1QhQr2lSeA2Qyj//wBPOQb1Di5kfnSq+mzeCNAoJcoGQP9ct3F
tBneduo6MvGDO4wVZZznUYDcqmBPCiJP3WAP6jt1tRFdVTtyrGGjY5IZ8lC8TxuB
ge0tHqaOJiUIRvAooD16+q3DUCND1Q21F8NAIQEFttVnXwRi/4hZLwBE77O4rArK
96+Apt+ic5f6SoQBGqF9gEng5HefKlSWg8uzxPqYzYwXBKra4BiFHzla3uITiD7f
mc9D6LkahygTYpgOszkUkZKJ8OGLR9gv8Y230Bk6HiEiz4IcvlihOepJVR+quFV6
h1eaQkMQW7Q91gxEC7QgtXlPluULjVbMjRgtumnCV2clKSDMZGIaJxOAh+BFZXBG
iy+MZB0x44S9HNtukug4klkozYlamo93u1hKwwBJ3RnT9hu3NWv7O8EK/i1Duswy
n7NHcnZd4rYorQo0IeVG3260SL9d4YekfEeMwsbGwDRPrVeaJ3FLFfpm2cYqQ7+5
5Oiv5ghKTo+nBnq/xWKMoUYaWYJSqR7XojD6rAi2749Hli6HIHlOQ1BUvGmwviUY
6VogYav489DD8d9y2GTqGpXOUyuc+xF5xpNqM6TycMiLJ0AuZ0ygws5C91VUmz5N
eINDC+4i+bZiXULOVBFk2U1zTwj0YJCoUI2yeGtOdLPci2mCrwjb3/rhr1w5icKz
oB8e9jlqZPdUJIdpDhjquQdi4Ghdl6auWwVeP/SnUjXiulbAqDi6WHpNjsT/5bVE
oe+fNPo/ClXvPQEmRWzQJ72X/el8hLVfzgNqld7+rIVU0m723Ya091/FaFPzrLjP
`pragma protect end_protected
