// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:03 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oJiA6Y1qp3aLHEXtYuLT/FRg+O6ro+zOUx/ItX3KZHM1Uqad9QfN8RR4ckKf3b4u
HLPExZuUx7PIOJfbMkde4mzuNeeXSDgzdwE04pHIk+2wJX6O04agMUc4aITqd6pp
r/jn7TaTqBAOeIHYn6PKbJYDFNvoXyo9bgPRgNTATQg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19264)
MU+SGeR4I7PderrJOIs2VP2BNr6SKCU52DN42kzdVvPeDSijD2NInxPpvxtl7hug
uQGXmRq+JWAqXa6sOw8QP8IYmyldCYHKsT3kcNADsbV67I3qqfEhSGY0gna3ClF/
xjaHnau7nSTlKSmyrPtUnApFfQBFVSXZ4hlpb2N7so1DvSMTxXFRzKXqh6LgZWz/
tVkHnuXZKs753btMP788EpP1g1D5RjUs37G20y+K3wkMKNyvKUc/GLLBOQg7PsdW
EVyCejh4GI97YqQTDK24GXA/jyT5aLL2wGot3PVZzzerxpRnh799wkCgMk8B5p6A
lNzMe+e4nRDcswp8cErR1nK1UUktt/JIrZJtd6+tKw3ce1qusra3LWyfLq3znZo3
nJbCoeCvAD7krTufHnOlFoptjQUMy8OHDJAow/1pbJqPw9/SvhpdZKWUoaSdzxNb
vtB9HgXIg5ElqZ+pXJ2OYt80NhUeD169SmkKPJoJbzE2NwxyycwiSk6uEGlW1G80
UvWwPUW+sqljStnHr8rAqsHTI4Lp3sb+2eetVzLNkmakXeTlt9NVFYlP3nWK/2J7
GMtk90sdJ31nNuRhzNLrb0IhWSyapvr1qARsmG6DvHUCqnbPhFv6pNqelhosDW0f
LaMrmVRo98nuFe0JUm2qjxE4Kfe/RGPITC8Ed+iTD7OF2pr0YLU1d7XqzJIiFUNB
jqVcjBspZt1rCGegi1wfY9vb5JGY9uMrKWXlmgg+PuREMr8nxC0p32eHV2VFh6XV
D28x7vuxdNyYpRY2RNVInYm+ipRzbGAPj7LmMQO+0zrxgzHvBL8HFptOOSuhMZj3
F3wKh8piTMGLAaSmx7mDXVMb1/2f5+KLV2FS8fT4AFyAcrJsH4m//AwHf9ujvFle
quuwT4AV/YGXR1R0ljIxrwHwccsLXqIrfAIlj+Do0ciTrur9/UWGa82Hxg5p9ar3
w5YCL3M/t5loMvkF4FRp/DlzGEiBXhL7RfiyzrF9fMUiR//R4yuZsIWJLXNPE6rr
5wm3NkJFPX6+Cdt19FIvgHXjU0XU5Yqa6XOW7q0g+jKEacABf+gyv2rHqCZT4SaT
VwpMwvPbCL7rRCUb+dkO06r2ZBiYa9X8m0bR/lBjbxRGrehcuREB1RR9LgN8xEfo
grYR/67LJ6IXqa8+tEnOJkGNC2lV3K6gsGgpwuP/UwAeYzg+tzqZd8qdrkG94i6W
hoQC1u1F90aqASLMLD/86k49K1DF4ARggSKk2LNCjQqfodncGsDIH0yIb6HJxb7B
H1srslS6fVHpm+EmAdYKkF7RVBLbsIw9CW7+oP5YEiIORGdxmn2Ff6imvaXYhc5C
AZy53DGiES+6ZI2n6BbonA0Ad14ugTu9pjgwsjJk28r3ajSxOGaMnNqIQZBPZaYM
L3h8mqQrRSORWLwugON7ItbF3YjxDl1LayJl0sOGFCKsL+i/ywgOO1EkrXiQMTlS
nK3C/7NXFdpUDN9CdBYRZsOqjo9RShKDvCdm/wrzTuQQ9HWt1byMMQeuABrpH7h5
P3BKW6qe7sUwv4zdTbcXImhGM9bhc5FLXuibjslWexUoJmViSTT0b4r3A9ZBYjX5
FTB6Lku/KCVSoNjSiYGe421f6fzTLCR5Nb5wkTt9WSAARM7PSM8GlB77Si+fzPKz
yg+UeTZtpW4HnXDWKRLkJuVaNieyDxg6Soqe1TvWdQJmOvPw4qM+oVYwZadtchO0
TauMw+SWAZ/u8C3zSupYRWAWgYqj4+EXKgQwluI1y0Zw6vJ292vGOGPH+AlXyFGc
ywArrZj9OJTpoSK59+O+quJS6BmMOyr/FhPsPsWLQAbE/5L/hzuvk0olHmanF3Sk
dTwEG6jVvnUGeQGklLIbJ11d5zmMtYLpvzdiBZTHabTC/RUN6Q5D+dUpn14PUwHG
sYDYPW4YXPQiSPLfLVX8sbBZySRV6irrV8BvjVfVtay0eGht797Xq8mt8bBQSb3Z
r7RIcfUh0agqdmeumfyW+UWRumoVB6ooIEOi/kQe3HUfMXOyoV4SRW40IeJKa/OD
jbFChawdYfjn+Ov2Wo3LYGKYZEGSi08hMwXGAnIFJnJzbpRK9aWbTRvFAZULSLw0
+jQcA0I/UyvP5bLXuwDyr7K/ZiTJ6TXi5Nq6o9cdHPmO53UD99GrLXUa/S1vFcTx
ZKyHE5e1lQlz/U0nrxNVDykyIQ8SxfDIPHBjkZJj12YBT8ra/dXmAhfn9GcFtbDX
4jvCHLRVJ07hQzOnv4tPbTiQu9HMhvy/nxCAXJulGdv3oPuVfvGR5cUkapSkY3wS
xzdYaGUV2z7vbafUlb/GXgnJLa571UAHq1ZU2wk7CF7+2NB7ohlOSiGuO16rHf2s
ByjEgRNvdZBpHUkxy4lrL4NVw/XrUwLnrLD+88lNrrtcjsyVNqgVEES92EY5H+2g
lG2O+jtP1+Huby90OyhTTTjZ20ftURsYLCnHm/vnyBL5u8MGbbF6HD3xi9UZF5Bo
zEsFV2DVi5oMT2FWMz2/nl+BVO8P9lDmNvaGTfZ0PLcaozfUqPiB+sqqGvLK7UC4
1mt3o86Sp/EXDDf8foNStaQvQtzzr8uV12nO0UHDJ+2CHGWjrnxy0Zq3kJ3k6y8T
fE3kZtzk3ArkI5U28Mc5vlfmYK65+PQozHA7fFPCv7OqjdJ+00DbptGFolMuoRNr
iUX7HfBu3sAk74ylvjwcSqYo1RthdhQpX/ekeiZ85dyEiOP/c29+BYUnMT6OpZvW
biLUX/U04+hM38+iCg0eOMyoM7DUoLTuiYHOTmyd5ovo1otHRxrb87OA6p3Q1Zcz
jZv4Ug974BjpBd/4pXyvSRDT3Br7DKAxMR1nQDUNNPMANZm0VDzThqkz3pKB3vOj
jKN0iiVKryqk+cqX1YBRjSdiheMt5vbbLZWAqKRzh73W8Mdjcx86+S7DuFFriok8
RjVK70JX9QkQCaqwANINeuaV3kPKKTSdB3yrl+wEh5Og+ckv/OpgHzrNKdB2dqHL
JgWRCkZAAVpYKi+5gI2+Poiz+o2R4BG9XRlomjugO0DxpatbSdQiNv8foQVvu7yI
6MPnlTX0jfsD5xk/O212qcC5K8OuWgPQkIdnMiJB78NaJ7RYS7+jK3Ukpei0r0N4
j6QZ4SQGbH1SbInz/uahc2Mhvg5/s86LNf88Xw8lW8Rih+kDaU+PzL+sa7I9qr1C
dzxX1Vv1qn6B/ePq+6n6TM2hM30v5R3q7dU1DMPtgdyH+h7oJAmOLa0ZldJbC1qa
UtZYEykaA7gaQoX/izZoALE7o2md8ZlbEOVnucisZ1IBQ6wmYSx413h3oSgyv0Es
8ez6IapfV/Q2QEFF7DPyN1q2kPuOEdmXx0ZKdSaonQpFjA3btZ/2SXKOxaVa8KIg
vPzh4YkkSh9rKP30qipikwi3G3GLCtYGlv/MUY8miC1Sq1eb/Lbk45Fmj9QG4Yzo
Q4Bkpl/8KUqpGGDUDLqcgjKZnLCBr7EOjsodwldk3o9gShdo0NXw2rKdXZcGJqHt
/iQlIddado8h4DuoYehp9ukJe6K4dYKsouR0D2MB73Mi2I9R5QHZt/xT5rcQtsqA
/K70iaZ72AaMoTJyS/HD7i79/9iDWBsCpK8J80ukG3AnetEuL2ntIXK0mQFdoKpu
m3T1XgaFg4J5d+6h7ZD3An/77OZQTwViIvuNOYu9/EqbVnNNYLZAiZZKVOyARi25
Gv++WcrqQVysxcfSq1Ih6NE2NKVUPxmIDkU0smsTMYo4agyYwx3CaHS8YUMmrpfg
e44z9yMYYmkHGZuTACv408jO5/0mb3idOVD8X3WlUnFmbl+N1RBuSF9stMpNLSYt
9A/vEz8Z9uT95MdY8xkPDZny/TKHXJjfvMnQx88R8quPkl5cxiFXtPhFTypKl5d3
718Fu9bXc5epiw9B8Q44ktfcnu7Jp4iWNpKzmSPexq96msWfvFIv6tmqBQhNy+Pz
bNVuA46V6prs53fCZi1830TKleRmPXaDRfYCUWgmbYcOboIGuWCNOIFx78qyNmOf
I6vEDs1pCYwgAJ897zbawk5dNEEOez4pfYRV0Paf6CyyYL9Hjz9RmdMdW4RfBmB6
+ITkW+dbG2M8oCfj7Gpa80cF/asAZeCi/Y7R66asgtnTVsRNalPPnqXWZle5q1mI
uJ/o8fDXcJurJh5QBUe41J/ipB3ysfnPiaixIitYzTmKer7CoF11HkUyVj5Y0yMV
LLPHA34er1HsHU38CE7pnnLjBTMiEgXxtdsLypAzQEnsv4XewaJxkKKrHgu77N3E
fSbSctRgNmZ1o6UI5UsA8RXslQLy5FVYymzMG6TJrtOOk02DXGefwlwDIxpFxsoc
0F0n9QQSIaeQzFo6A0UNrBZlTK/Gkln16AGdz4/xQkEgQzueUinzzWHFbaGskK75
OZ2QLeF1rEeHmBzWo5tTlWN4C45HdtKmOJhmlhiFIh4i1aIlBt636w4jWBmTlZkM
bN0eifzTBI3pKC1WppP3h+5kTC+6ET7xwrEP5UA0kcBl1Fztb8OLyKdDfoywHOmq
ZVMeBi2EwI8Ih/wyAG8lg/0DlW1vIdYBcsheMj+OIKL1XkD5rN3dbedJvxcyZ/sY
48TzSn8F5MBgA3MTT8+OjvFGSahpN7mCMBj6ZOZnYznL2hn+V9st12FdJu8eKWon
lYqF4V/04PWbAYpnuKWzlHoiwIpHC7j+aaB+my11E6WQ23zPEprBcXuaqhUXwOSP
98c8FkRiI9NRWAxKALtIMIhrOh18xtzS8NQ+JJpZzpAG5c/5JZYJaz/gFFR4C9d1
9ixzGw2kjKysFMtrhWfnmTgEh3r42lRGlRixEyszDGlfXesPrqIozXZwJl5kccDD
p+xFO1cfqghmvliX5TVLIwOL5y5Mr1oRV2MBsk860upFu+XYqHsPeU4X0gI5OOmS
fZ2+bSU6vPFdMeUbQ7ccKU4CDjGAupiddYyCX40nJ+GBB3Ye8axI6H4FMJiTdUSa
bDULi/7Poi9K3T/yGu2VUTRcG8jumqZHzhgBFFrd+V6rhkKomGh5epp6GOZ/L4Hu
fhIRy7nGVZi64dYLWAWfm7K1XePQPZUmOKxSZF7lHgYNFGV6l1AexPHuOi4YNyio
r6N+3U4g9et0XdH4ttpmSML6AMHyiw7OghskGvb6tDppyJTjY7XipfY6k902tlIF
grMB0YbBhMRzGGzQvEKycPqV6EUaZyqwvCZSZmUish6joXq/QR5H4gI9vQcazQ0m
P+8dQwdJxiVRafMzPBFAVAL0DIbxa3uugdNjdZN5JnziwRVxRw3pPaNG9iI9C2Gd
O5S6GaXpdtlh8TtTPEWHteEa/MI05BNNmlh/YSryEjtB/IQCStFhwliF4NnXDnwP
QMJJBk28ldto4ufDfQZrC0d6UH/NaMfVGoX9mq0MxHgSdsOWCFk+jh3LcZZQmrIS
87MFbaqCkVsWfrGGX0mZxad+QCclx06/JwkayyVOJr7RKi6HXzXiW0rSdjAGv34g
oxy5kN9i94gfpdWHFm/CoazfW8TdeiTu3LZXru8Gxd0t3MYd0Q7BLFEieQ8an3xC
Gr1GFyNBIoPLDycsYkpYuQgAN9S4xdTXDWbbIXCrFn8FsUeHR6YBk7BGKd3NxbhI
GxgQe6/ufIv+uXOSiEQlYIy/MB/oB4U4lVJqaaRFWDtt5sAL/yVnnC5lflG/SzPA
AcXKK79TeHXKGyp2b0d17xdY1Pdz10SlJr5HG0/OjJmRT/apcZMxp8n/j59J0lUm
8T2LE32U+nHaD3wVVvAKBbcFAOqf5aS0h85jgRojjhPGlDgWjsEJ8wczEU5kYRMO
uZ46QJgfSs3hzJ9zpx49e0NC26qfRWZ8oAg64tW5z4bMbDZMAxeCFsPGTv19i5iv
q/QeNv33lqTflojmc8Ap79Idcb58yz3VsiLDQG4YySZs7IVc+3PQdyN/rUbO2xCB
OlPRZ6KvkoJlZ4Z8uVmpn5s9dX7DE88jHhHpGAvzERIQ14Nu4Y7IkVuqNi00hvuS
djSLCuNyX/PmAUCFG66GIS76Z1whiCrz8ybMBNgVkjsf/RhHLfKGtu4ojeTwNBnL
72O8F1nAAeFa7B9OKk3WpXC/2GdddRMGcjrmmoiIhzffHmKnurCqKw0UMGxZWuKJ
hC8B2l/ZxcCmWTD1ca/fdd6jCVaHdt5mHt7Gd6FG3B5f472IBlUALUrGSMuA1bpF
Y2ufUu78NsokbHg5JeEG+BF1tw7clV0iADXLED9JutCTG4Wc5IC3bXRWkNe58/2i
fF9QLxd1O3OBZTjF7IYMJU47bCWTbeJ1DnrD9MLYS62K+VXf7aSFiL4+WZVQ+uWp
rawJgM/j9kZ3oCISmjza6+ww/mNAgAAowRAGPB35G5qRY1nSYQI6d3l4pprpZYH7
emTeTtLbHf6bQGr6cdBA+5yv3QQ9+gPPQ8M5cikmcj/40ezv5as6RTLWLqnw8D7I
UIF+G2lOZ6xjpTHi/zOyjZRgrQjkul7RgcllcCtozp5JW+Mxk34rbn0KM84EJmAr
8s+6kTMGR3he2G5vPfScHy0gQ5BE4MEcu3BqzLi18d2Sdif+aYGZHZqMqNZ+hMVQ
uONMo5307s+JWUq30/rm/blzaai0qAhdU/TTdrgs3VW16pGYV51feiBYM7n8ze0r
gTl2buKl0R/8HrPqdxB4r/RkKYDPcQ7HNfeLaHV8p7Ux1RmrQlqAST3pyyGpOgDT
2JsuFiuI3KLPDevCl+XBj6wLSGBORirMB2pGUi2HG4Atft2Ln76FeeJM23vXB6t7
aqurnpqHOs0yoo+tcB7wGNr+ZRMk//R0xJ2/rfhd2cj24R+i8Tc3DVNdXJg0rPzs
6UhPXvIwpP39Oh4aAMb5VDzmbDd10QKhgHWF73SawtYZ11t9DDjttGTCSprkqQP5
XKuqKlQMxMLOODozPyYXUKW15W64WCjVccxPSc0u4bjp8qKhlncpaP0BhFR0/32f
XvIOi0cUudeC3jGELgk6Hn5+Lv978ZiCEv2K3bPCOuDEL6IPYKE22N7fXIT/rZ9r
anOCO7AUUQLMEt4LOHdBU+yckUL+fCpuyy81p1X8+SGRSofBTfhofV3tQVCKgasA
KRjVz3LksEH81KQc8egRUgIfe1UL+eSykdJrKk+saQLBlLrCYtdQbnjK4rLlO3tt
pxVv1dskrbVYHgy07WdR+mMOTaMBAIPchISAPsuSjCjL8ZrqL+Yb0zdRdLiyYfQD
V2yzqxyKvYmPGCl0Pb0OnGSq56D19u9X6Ve9i+zd4oBaUHndoBNaa1QjD3DNeGU/
yyfiFYU8e39gVXroylcc/BPE3wb28fNMVvT3RuFd1DnLCUE5cJFfJSx+1MikSii0
ZT0QG/9MIn31zU6TjGn1VK3NU0KGM8UVc6OfENLd9hqZizxHVT6kxoitC9Dy/3iQ
e8BNEU4MmCqs+PXKwItj1FwzEGOnXhkZfzHYi3qldpjiHooiT8fhyrBuIFfnXe1e
VrpqFXBj7u3VbkN6vVBrbgjVLPFZfUCAj7tbB561FpN2mX/IEbcbajKt4Zdx4I5G
+9wdlD2e2/2KZK3zcAzHIDNCVz+4nxwKOlqzn7aWLTKJpnWbl2wDAIsmRil87WXP
u13g57Q2Ml8++Oj5ZMfuD4GS/S4iWFgbm11jVbnF1ljSUJ6I6+m2Chx8dXv6ifXb
xDbr9FGNC8BOB7BfkKgcoy7efpWvcAZGCh5iCcYagsWB96BA1KHlls1JDXpstU7l
RdYwwoyOBIyQHvaS3fzVfYK4ZiqciYclaaA+O+LA1dPMpRful8kap0k1AjagPJLt
yB364a9bqqcb1zZwkDNDlm4+FfR1wrSv9EVyhEOrUjfwE/3Ui8owWZaoidbmoH0D
MEDhRxMDpNlzrD2JmgzhKVLFaAEOV8QbX+5UqiILJhfPXbKmrFi8ukqQ8t9Jqp+u
+gBkq0kK1VrgdWID+lsjH2wDyGPl+PpC86sbrQ/LjnjL4OPfsSaJ53tI4j0rvhv7
t+/GndmujoGLmGforF18I/mEi4YvRQQ5RKZLVKnOLaBiWmg+nGZLdPyKKVgpO4Yk
ky/5sDW/ei5D6tEpMQVsGXhuTRDjRh6fpJ/Moor4DpH6jl9yco/SDeW2iBGPKrtk
UTQD5QNtOW9c+oqGLIQ7/G63ECuABKVauAueXoFpNAltU3skeWx9gvQif4ZY8S6Y
0vVtYJEgPzlr8ceEoWrMq7JW4VC0xkyYCeTEOgcm57yOl5cJnc7VG+YZTZvOobHV
QcPKj0j0kwhDHmi0LhNbgIZQ8qeuQLG9fJ7BMfDI3z/5iEBQv15ETJeFRWde7EnH
8AI2akSndmb6PojC4sB/3kJX3L1uxNp/j473Tt4SFcM+P8oLfgrWNS4GGcHaX+5l
wyTRN1e+at1ygobaLB1imh3eAwB8l5bRHGyoRYgvxcqsasqCEdgk0xD25n4TJfn7
GBmUZ8/v3AlLCWAJclU0lO5XvPVJLl9eArccFGQh0M/kc6VN1hCHGU0ZahKbIv7n
uqYyEe1+/a3l+zdjjtxkovaAgHSa2Wsc3eR27i9Qpd3/xsqMplCRrecvEGpa9qoh
96aZfVEHcH7Xw4HLNZZh9Axg3deYw6o8g/5R/2ueA9Dhix4Gh/mzjucV8bUod7fP
r0sP7sbFWf/Z4h+n9wgY/c1HcDbGzuJl0zkdlc7Q1m47W79vPdNitQXbVCCw8mHJ
brKhL+wQMhJXwq4wRngJcejL6OCJ9+C/275uuBmUyo2CAZqMlpTF31IbzsUtuV7Q
dwsBRUoNDdDMU0E/YFnpYl/kDHeK3Ul2//U5KtI8nRyvb0WEIcyBSIhbxst9jq5T
CnTNe/Vo5SZo+sEstepe+OP21ABLWXD8qe0pW+r27Y70VWEh2uCfWP5GLLE74N15
UhkNEMAxpfqwpJfb76TaJHXaI05VuGlpWvBp40otGDnCWWFDmsuBj8egbaejLl5+
l9I/0EyBQiJFlV8o2XInd0AfxgRUzyJh62+H+FaaAQfXp9y4j06jz6uwtJc3v2XO
sP4qGQfwOGG81HYW8ZlYl0NCvo3C2ahm+jpT98BGyVkBwtnkeyulZAc8ru/10l/7
IXWUCabGIw8sMDl31JCaQCK8tCVyjrVuTkDWj90gFan/urDm/bvgOtap9eJxIpGj
0cjSafudOazr1+n10oWS6ctpJ+2tYFrFuUcebmDhys0flGkUj/iMT0E5lCniqLPk
upfpz2afQuui5FBibffTVSgqcp0Y/8bUIo1RByOjVhEtH2O4zJl6ITdi0x7XvBAn
WWUhP+kmkwwGTd5t5aTg2PZDKDsQUUXRXGYlNc7e6ujF71aGvazHKytzElePKiPN
B1y77U6XtaBlp8ig6x/nqwPllvgSF9vCjYlv97do+hUJ1xJH/iszBppI3OHcnSth
PAWg9rPq3E0lFEn0+1ZIp2zRlsrxPsTCopMZtmA92RrJhV26fE0yTdIZtjZWDQjI
3msxSM9+/lib3zmUykxS14c3L0kLIVv8GUgchkiL6v/F9JWoNbZBJjhZBTfD43vG
4zFB8L98Y28n8BKTieX2uTLBVTD53IqawamK0NFglNIqB44MxgW7naG9OBex6rfo
C4jnzX4uboOMyjU9XAAJxjE5/dLHiUz4Jw0NgeUagZaKEekEpYfdYlOP37TKQ93p
cUlWS2/GhniyfblJNyxzrJKhnpLYYy8BXVSqU4NIoWvg7IDT6pqiuvwGtzQ/HZp3
rz8WxRoGC9YYRbTI3MEN5rXrJVQjzL11Yb4QVQtOt53gpRO+GfK+UWgZrqtm75s2
Prn7k42LL0HvRtbQ4dZN8G35e2IFgZm+btvAGomz52j+M/nAwrFqpfNRKtCm0Pm5
8lp4bn6J0Ky0Wvck6bSqrF0Gxi1diTHjy2UH7HcD+Mt8FcDGB6d5onsFmIX7lg8K
O2RLuv65lnGJ39O+5E7Uhxlvgk7m8TY0tbuT/WENEjPpeeFoEmg621ynqLY5puNr
+2SRrzBGOb9JVbPZ+5czNrlRC+SEO54tL4fQYcoo7YIRAj51NMeJfrGLTsw74xU1
bjV6wfWhnsRQ2to/hadSL6SpWpMnfmNfrN9RneRu6GRy7X//Mc0uwTAu3pxbl0d/
ZPazvt+stjyBTw10bqb0EU+h8zZ37u3pv3zWG+Bgpa7J9Us8hxgHekTXUehVOx1g
pq5CKMFKx0rxghN1uNwXDhzojfxeDIMSJeIfwxcEY7n0LqIhC7/OoEFGSTr1+rPk
jpG23N+vKsLEyo+yqWBdlXY5gQJBRZ3G+H83xlePO4iSKsVXgac+ZQmB1dLkhVyC
+DFxzG1wB/ckdH4wNEtyT4I/340vkNbGV7cq/5/FnzjRPilHgDBG4YZf0ydYv1k4
e/09FddH1hocN6HipBKJC27Tfdt0/+p5CZUcm81qxNggiIhhtOgQNsD9+RantCvR
MlhBYpRknNyVKFc4oDMYrCxBb8g97vQcNdj9QNPBjIvUj3Q8gU8veh4SmvLEni4r
9sVoEO6KUdvF44V0M7EkjAiar0WFo8B5n3sUKhKWOUCTxkX5egjs6BOHCvET2m7n
UWJKyPnpa9p5/sh8XHSS3P2O1YxgwsZDTd3arfeqjAUZV1f86EWmoVvFlCxjCToW
asqnvbi72AcbUynkn+eIep22LRsBaBfjeetHbmNm696ZSJtjhFxGZCuYfin/QaOW
pQGBC7eHD6lmgCMgrnNPvGfpuqSFla6L6euHKRPq84c06aKHZT8iDAHXeimjYS6j
tWBgeU+JWTcUrsozcvjOPhBVaDWy100uE+D8FyLB+eQHc0i7TQYxQ7sf10rbqdo8
PUgvJ8nHZMS/y9LGj0hI4fHUAC4ZaR1F3i6/nFM1PUCnQ/V7eeedC9yQ+WNatfZr
+GVkLj+BxlQJ1SJHXMMj8PGvTK70NqG0X14dpzmxWORvoPEz8TYhK2CQ8ANRz0IH
Aoca9Zodlf2efkT+FC+Rt5aKYXghP4BBSjJNIRl6brYcd9Cut8vTBFippsI49bOl
e9MCPC71q5bb6SwqmySsld2vLY0I7tOsmSt+0smg+z0qrECMQwrwOnd6ZcgruBr8
5CNJDWLhsM75hKhWsx7WE7jsNMgugut5nswZHd76mTJY67ZljRWmHU7v7gN7hGqJ
Af91aCgqo6CEOOxFiwE4F12b0xLRJEzsd4rGp3t8ghVOcb0QEJonOlvcDnCFaJZh
s2ylefHfeqFVR94SEHIMbliNR0JUQCk+a+pXq79WPYO6gJiLds3BEQRfZkuedgRz
GheXiPVyxMXc18ul43vxT/zARRlFwYZdfyVaSK5i8Tej0cFfwHWnjfiQIpRXSAPP
Da3ioQa9C5CLME5/XxgZA+1loMHN6o6jO4NjMX5mT7AtOvDgP6cNCiMUZ38+MmJS
nLUGxH0hHMxphJEs+bcDGmTf/73XM4zXOYFYdHUyihuBFS98QMFWplk4zwkhRe2r
cdVUzi2cNtWKVCedgE6YPgFNrlgKcDfHJWpWjsYTq3xS/fTdvuS1mo3KtKX1hfnF
kv+9C7YFZ7LgS4VOTVm6k1EiZEQmPHR0YU3Yw0xHkFj5iUGYP4XjQ3lZS6NxdmoN
Q4TMtAOB1B23kh/v72PKWMHNolalcQ8sbqCXcwTT93Gcj697cJjZ2IJLkuKCJtAl
ZQlQwqG0EmWLMpBRWp8DUPVmqOwSmPSK9Bk3g832yiOCK2CnasD1fomhP7rh3wTw
PeR2TSJEqhbIkwbNH9ADjWA71z2JdYyczA3BXqy/wy/tjChOTg0tYEUvdmsX3sU9
+qyy299/iZeUwryTDDosjKgVCzZfcGd/wVWh7jQlRKy3lxhDm73R99Fo3LL9kBzh
N0TuzHV8QLfo0vlOrczjQLZLblL6KxKFQRMk9+TEvcLMA4iZ0YE/rIdZh7ScsmgI
Hh8azxT2lBnWBmpP1YhJTOxoiqdyZ5+UzNnyIr9/t5wmo4+HYm7Eu4yvELUvejUu
yn8dXn+gUucpsI1PJpfsmxiy6+BZWyg2dM6zzbiZ/+T0ZGMXLbc57UMP69kF4FUa
AlnryYeZKfOKWoPdO+pQkjjwskb2n5vharQTd4wDXYed235vgmIm4naRkJLLWTKY
BWHSNw7FIKs1tQJq7wdOZnaxD5XtaSuWpqTZt2Mc8+l2DFoGIVcmgCtw4f4jim9G
sjKckxZ+DvzJfoNirF3mNB3kHfOw9NuoG+kuP/XxVF7FR3qvsB+BpxaIow1FhVGr
A5QqbeyeVrRQ/C9jlVoL6uYwuKL4eqhq3Oq2TkU0A7sxhuF2jSvaeNcnkpgpf1DZ
R4at+Dsn/YJGktuZQk0xncSbrUI1k2TeIcFfu+oS4o078PhoK02/us8SnMldvNSB
riCcDSejN0ADVuk76VxhJU22Mbgl2cHs2Wj0pfua4teagQA02sbQ8QhMFZbL919E
knmzAIVtVNznMFKlcRFZ3DYPsKAjKbmWvhf1gTt2mS2WUq4aPzZsg4ODIsBAxXTA
fuUb9DUeMBh/n0J4RbooyARRMgWNbXBeshVsfvACZcnNCI4Ylucpr96idnXyh7rk
fVjZNtCe4OyamD2fUgsz8v9LP6Q2p0gkyLl68hvII9sR+VcvQ2HSGh/YZUFFGqQx
iMGc1MWUYDrknf/idQPjInNt9ozEzGmUie5NpM7/YEXQx8v041u7ScZHB3nRlzTH
Uu1rxY+Qnceee+9uQZEG9BBe2xwJ6G813X1yH90aYjDtKzVzo2N7sVKf7wq4CJ6t
JGgd7aNEMdCsc0wRxZwPSYfDXacOGIWEhJki8dBWGy1LFQ3wWA99BwXi3fGeZBij
niD36wsD1sULeJyWGumXjgcA+nUuE7J/egSEH5wlFZpZEmu9u6UhkP0VC+0bBlJe
80rqdMVGl4ggUo1cEyS9vvV7f+GQgfr4+m+I+OXFeSQGYsbV3FipnuPINSTFvxTR
ak5r2l0ZXfTh8d4WIehffsXrH+ejgj0KEa1SmmjpIpQSKJm8piecQkoX/IzSNT/3
+YoHRyxcMbKEhM3SUr/8pMhUxEBUQIR2C6i1nLUOv4YTIyk0f2hdcXEAHBEcM6VG
83UTU7nrjbkZlOfZFfcZkGfEoy75UeA4ZrN4pp4Ht4YYD64UXhs37WLVbtEIniZZ
WtoRXuZqw7qhirqImtN3nQycXGWKS650qWMqWKPVDheEZyDBn+WgdiY1q0GZ4fhJ
cmWA4rgJh7hsTy6VlRO4JutcMUcXRdTIXqCnbdtl+7od3q5He2J3WU1/MOZVFs+M
+DAkh6tpqjg5XrDKEzmxyL9oDGE//8FJGll4VWbVhAVqW4CDjI2R5+g6nO1Cda5O
z3q2fvnxRPNRQmiO+I68+31/RQNWXxqmlvIIPRdds9jfjMahRFBitZ/P7LRA1dOi
5+gipv3HIVk1h4Ih9+/nr8+Z2TZnyXQFmWrv9fCMoUF+4kSRQtGeTgPOtCegkimm
4QZQcpWGWlVtFngZ7mb7LRIKa1kj1hk/j42b2HPffTjkW+9havbe14Fi6Y0vy627
KcSzKYSFB3B1jvE22bMwmM6kfyww+f5JNUjSRTx1Y30Ly8pZ2s62utbbUFUfQA5c
DdTlA3lSv3GmBVeyFqDcchDdrSq+QwlEmCs0TyrY6PQ4OGxAKzdxlems5du7QFQA
t2Tfgg+LFVbRfEgWGSXVqZlmk76cAww8TzJxQnAI1Qrzo8agp0R2vs3BgCcBuFA9
Tvjzn7Z3XVOir/ByZIpg8blXr9ZWFJWBReS8z7jrLfzkyNROriiunqhQmYwMx4+P
TA/vAu0eBYAZf122541Io4DKeVonpesr6zY8zc6vfPsDd7PF01xy4D5BrjR8WOr8
K2FrQVFxWY7n7Rndz4wLMIY1Hci6jI0rMm27g5LDAler9T0YzeN5YNuZLAIrbPl1
Bn545g+PbflhCnxaG6qfd/Knn10NU2ddzMs2kcppIsMcchuS929AlMv4RrcZ4cqH
mn6kB3aoMKsbFdtr91B8JTSUA7+q3AEs+W/1Uk8FhtM58Gg4RvW8bAGbrocrrsAJ
GBotr5rNyLzsme0UgRCkKwtHSHgpdoG+wTYTzSn6hjK+3lb0aTePLTbaBY3Vs5Fs
jfhft5ju5Y3Niit82FITTyyF9Qjbafy3/Mz9Un57yAHlVY5sTdYPcNQHQ//wM/wY
uEbTpaA9yYF5yFEL9T38540A956GYwKe+A7s4hK0+uOGbJ8q2o0QPAROvYzWnoo8
v/Haz6mZFb1C6yx77wUJJl861dbzIWqRkKgmj5tKQhWJNkO5N1YqLJ/DrTPtfOg+
X04R/o/778SHQCAPY9RtACA1sANlxmUHzHlb4lVRyFHDPh+Fl8LYG9JSucz3PZ2q
9VnRY9oAFXRYMAQOqesRoSgRERfL+CeAA8nc8vt+B09Lvr521X7UnK0uzXL8C9sZ
pDZ4NWFR5bJG+5pSq7EDeIgQNMYZcHXFlcFL0JHnGmcKxXM7PQRwgJjA+BHbOp+y
SIteIMQ8n3S2g614jQvAc2mEq0Q9kqEqN+SSq6C7kPJXv/dF7caPdtEl699iJURx
qW0NasLP004AYQ07imeyz2P9aPK6J5Y1G9OYgucAdHb5f9xANAwp8G82CPgzxDlx
toosH+XgMr4/K7erTsBmKbuSuJcWzNoO2KaUPR8+MsseXGhx/uQEy6OpkWpZYPKl
x84Ad8kbSKwm9AAT+qtbH93AXbhkYusYI7cXJ15ynvcFl0nf9zEi+ryq++vwxdSo
6pe6bYgLQb2oLzSj/5pMYrTVvVi7ivLEGS23A+9Gb5xt2uV9Ptp1T9O7JLFboHLF
WkFicppmSrMaW2wxo63LuXaesqiIgmCrVDzo/njX63uToeR8XckLHcpSS+FiUs80
NSwaVZ2mSTU9o7H7vVQUoYvSKElp/A+DN2iCa0gcDa2EXPEcO5M0rErTSCexCGLG
iaPKhvzH9ROVXEDVgXGgQJzCATd1XGKZ2T3A+8Bb3Ndh1q8RPUg+A0Q1mkzgT5mZ
BCFDDGAVYm2hG/RUnIneRZu3ctl/evi3ZvpezhHNRZN9RgOwJzCOLP4gm7i+i69Z
VkGW5BJJ9fsYz3tjNyAd6SOVewMg9Sui+gpN2c6omro5+V4N28YJo6Tr1MW57efh
Jj1Ml7fah3OD21QbqPmoWVyela3rkns1wyoqE0KD5zir4VMaDcUGNYE+fehUJVCu
dqGBjcmhgT/1YdWEgZXSfkLe0XKPNJuDJLs2OKdHaSergVZwRfL4cRVIOrqDPFiK
Quvjjt6fTeZHwirgkYCh8mXTFYKAJrVbiqqocawZ9BfHmiMBUr1NQrxnQ36ETEKo
bkl8jkpUPSg4w+hVzr4dP8SNxBvTwj4Sk7I2n2H7h54wPZafjj4pUUbdTR49FHoI
j0pZYat9wF8YNmIvXmMhzyc0loVmZdsmK71G0g9RDyMWmnQvVvChRV/AgCG+QALy
0X/n+eLFQz9ysIXBHE1vLL+2qwOwPaqsylIB130OwwiAYb4TtgkSEGGhu+SjJIbA
F8fc6mJBf3I0YI5ElW8A+99+0Y/uinZPFYsV8hKKt+xI7gif55++sAUSVGaoNXZ0
oO9V7H9sj/uWlkkBOzCJyaXUG1IWTC4M4dyHhkk5zebtmPuj0wxC2kaOLWXUSE7s
/nqejrm7EaqMA4WiKJJhMwmcBhq1VIP2D1strseBRz3Uojc1+EJJGDzS2vh0G0Zc
BNJMZghtYTWvPFSc/55lsnGrQW0NbFU1GiLbf5vFEfHcCEW8zRVGXzBVf4mDr1G/
2cMaFULomjgxv9sbnt30XcfaxW9TPTO7rV0ifA8gcWq6x6agSPQIW2WR4xrQsm67
DiljguyORuaLRJsnXIVp4KQE58UUqrznumeLYG1SqxyiVzic+4qvJzp6hlhfE6Z+
4ucsjiFvRgFRijEoSdzbpdvslWg6bjHbIwrxQbwKyIyYquTD77kH3tWiNtN+JzzB
CfVA9Vz8uk2xo992Xxx0NEl9u14mY8qfEC0IA2R2Wi0S+2dkV8m386q15fWyToAL
7pwuUs3PvNq5oFJDKA8vxZ0xoqKkryDBNeF7YiTPkEu8YENZqgo6fnTnjlB1s26h
39KuzMg8RxQOzInaQyjLP6xcR2yaLx+qqvl5M0SzAQFd7TSfrI3LaX4bY1OBjfbN
lV+WQRhk8O0tXmkmqRans5lGeT4vLftCkTWCxg3T8s47Q+J057AX3+7iW2fbH/wp
TNhkDDP/yIOLE0Pdgd499EYzQ/ClM2lSfGqIUTV16kBCP7QYkeIdvB2YTHDRuu6S
9CK4H6TukzTh0mBKIlMlXy2B9vPa7aCfdThsvBGoHQVuTIPugGrAAjvHwvbMCpVX
UDrvJtvFKrMIHiniAqhHh4fdmsj/Ro8QBWppitQGnem18GXomxFL6A6haqIwAYCJ
xhMsM5fxe0ZEZbD9yazOkQQ42atTdUl/mjXXc69xjhKzuj+pYPGJha6J1hgYynNO
fcpKkDuyUdJN19tj/N8d9NQzzBsBGkz08iKMK/PPkVyw4KhuFteW5fWzAdHCJ6b3
EhkcHn3Fv3mQwYGMpRRr4sbRsHdorEXNrSvsXE3ilF/Gujf3nHPRcsneWAb+hzhN
g+rNiAIpMuAvZosoPAo8lF4m+D2nVuqdGVNfIoTqKOdu3t1lyR0ga3FjfiN0dVk9
UN4D9aITK1N2BO1RhUhWlrf2FJN6dvscVjQzx4Po0PA4/5zbW0zll9peYuBk5O5h
ODsnrkvFAU7n1pxO/syAjsOyUXNagtMhsxxryVNjKE3Evah1dhq7/FooKuct2BlY
sQDjaqYyCJon3dDxDxtdJnQ0ff5SErDl0Utnk3LoIPc8VTIkYZDwwIJKUKkgz1gc
l272IxovcWgqqTbrFvD7KonmT/oU4Z+6zBvyij4IgStLw0mMyRlK9jUc4/zcwoes
S+WYgJ4F5LNWXKQae9e7tosKWuvUadr2AdHiYNq86tGFemAbKIfPPIrU2OPG6PAA
/DQyZ2EzVQ+8Qsq6V5AfiPyfWtrDNJmmor0VQesAQ+AzL8NjfKBzHGb6eRFowI14
kPoOvlnt25GbIP7wEtIgr1gIlKF72rVUhqfJcCJhgtKiFFkoyyh/imgwTauRGjLM
7AUYo5pTE5J8OVef0AeruVtVz6MUEChKjoqgb+3cOeZnV6KBSXHm7QQEe2Ak63Pp
+5CHQsNc1evnm0XpEZ5AUgn25FzAeZhEcDbKcTCMyAtQnrvpQRxAfMKfwa8ZpzUO
+WEl7Y4kiM0wrCwXKca1/voLBNfm4ugJDr2AJ4t0k30e8Z44vwx8tyMatnIhn/SS
vZIlgfNKEKzsK9TLJj5vj5EaNFSVVVGt31YWffMvFQ0okwBHlIxHee8iZ/yg3muE
z3XtmJSFoNLqhpFqb8g+yuwS9J5WOEE6VTAFedpHHBAkc8xXiUNcqw+t2RzmGqwj
ZK08z4UosZTPM3bVTEXOarvb3+K5uVI5j61U3LVWq3KqniXfLRr1vy4khG6q6tyz
hnbKfZwwLZO8cc5Q2kN78LakjjFEEH/PbBl81Ag6WkIB41qdOYKgdaeoFkhTSdvc
x7/KVCnvst3F+DmUcU+pbFmMkwyuVNAewkiriAy9tHskuwIEYtB5nDY5rnshM9cG
ngUo2kcTk2ZiZDt74kGhgDwfUqqaYgcZUgHQfzrInWnWOVw6YhtdDmkoyjLyuviH
qDBzFH1QTNEPpWTj2oBn+/IQx5eQb8py0s33WK+3EBnGh3G5vJ5AoSy41wk4SFaT
U9NZu0MVeI+ywzEuHJmGUWWXBPH+SIr9SHfpzi0GqR5uG04lQu2ge6TvrkCPNsQz
dZ8bjtJzMzsL40Uz6gUHhgezfiwQOvRJze/plFuX5JgbJJzdySfL1hMcIQHn8CCB
PI+8ulUEPQ2vE/8bmdxyb/gPFBjN8sWpoOe0yG1Y1Uj6+OVDRCl/GIHKJg6dM7GC
PzhuvkIdjnq609fgqM+Xm9PlvCLG7t67RV4rtfn9u1482mZTFukHcoPfTa0kWTN1
bvWrG53mrowB1wcfWc5l9b4YwdO46ph57daSncFcLn2W08xcaeMkua+rikhLyXwr
ndmGjsNjXSuS16NkBsH17iyj4b4DA5Z+NeKmNOCIzGHz1QWzbOzBNmaioa9HaDLV
/L67Ahg4LcLaA56/fEDvVO7baPkenG7fAqLXahUSDodTvbTI9ln8c/JsPBM3XzyO
Y85mQmS8bO6syO0237psQVdecqMTe4SKhSojpp0+hWF09+6Ay+yOfhaK0CHOgEey
HXQNgOBII0kljGXepB8bkFvjVgHv++8s/8CzuQG+B1VWsvatbt7d+59sppv9+1aw
FG8JuAHBMEGb+IMJMUX3xrN3lmcU09tsJ566boXHixOq0wes2eIqsBvyP59yK3iP
LOsbh48/CpNPBNl5SH4ZSQ1SlqBS2s7UIvKn0B0drkzkuKNpUyVyHl7Up6iXw0i7
WuvJUlB6tmIWwF9QUvfB4iM8oea3z5B7hTBxukQdQCLl61ZXQtK+6LWPvahCX8yZ
cD5yJu2KhAcBcUyjBYZfThKt+YRb7JAhtZvrQhMiKgJY/Nyvc9NP29swfT84cjT8
nIEmCyitUcgT7XFmZaDj4acx03LtpEq1Y2Y1f7QxyyZ8z/MNEYiBQW5Yh5m4kPgb
3/SdMd2L1Z5WsoCliIq2aR8ocV+wh16Bf2XMV6o66xxHmc7QD254sSKshOcx704O
7rZDKV8PxK1SMyY1kCzPQ6wm+ymXCQICbiiu5vTi+zEvbumEVAE3UZCjwMxbbNy0
bw29DCK++FEd3kLuixSLoDJhWRJnDBwsmr0JLeq9lXo6tUnbFA7FfDX36rBnTjxd
FGJTgRmMkDUYGL1TPj7bP3vhM8SoG7c3HFYOzdspbYjJkN2xE71IQJebzOoDQnSA
dNsLDDJdFTEb91Tbeg/nJa+B8k51/8/Y0z10NHYr0CLT7wbsJ3DGBo98sSDCBLYh
ewBtBRqkPT2kQF2h/XgVEoJ7JZbMjLCCGRs1aAlBan/7Kqk+z+7vrvddLlBxMMbZ
5mqq+q5NPid/iP/HTfWS7uUd6z37RrHfkYr7lV+ydBmaZe0LrJUG6gIeMdgbkm46
WzSUfYnJ/l1zLKML9TH5z2HdN9JpcJl4iQMEb5zTxC/6LUjyLibuNVont87wiDbn
AFVoA53GzHRyIwjLjZMhpkwkyOpiPXhb/lJHy/W8CkbtSkupht3BsXrvrSm8+v+/
DLEqsOWgj2ujELU/gL8UmLc2U8xHN/HvfYjmHle+TbLM9F/PsmghmeTQFjmghjWB
kB4Yv/dfwG1Tu+QF8MA7ueH+lJhrSaTzt+hsFpXylTr9kAWwQU+3NzWq1/O0gEt4
gQsErNOQC3kD4Jyi9NIOACmENOnJM13xXdKAYSouB2Ps8ueVIe/3xER+xk+CkyNE
hWeN+0iulEz5Co4HjDHE5ZuwopJVcjyb3lsXCQ1fOKd8x8EjyJqiWGPGuq1GiCMt
prBGjZNVMEGdfZ9Fahcta6xAZxiX2fcn+NjojOXe6LRwRx1VEg7JcwqeBFrcjKf8
CPUWpsRRvKhyQti+zgV9Zm1qYYzerAQ/phFl1uUNXjfqEn3KS/J5okGZXt6yStVU
kDcLxvSmJL1SGFjuhAFvx1r3xOJqassWjkhXoTS/TPhIPpJolWch7ur7pWIxd77W
Zs/k+pH7yigdVYFWpkF2USRsjdUf8hb+qJzOwMioHM3XC5jFHq1+1h26MdCrHh23
dXWCBCmpW6aeUMfb+uGX6O3oqZhdyDIFCKCZ0utwMwEkLATzRpq8DOi20yaJxwr7
7QBQ6+q5Z40src7iUdPrjSSeKiOaDHNXtY4YEZWNssuxcffIkRKCZGVjT9YWABg4
4gZuAhXQO/eB+7wZUyRNY68cocGrQ6zSFtoNUE/RDGvIZyLamMMbODt++kcRxRyW
wUTHMZ8OSWpOi5xNXamovNo+/KVCH9x1Q/t9+be0Mr+qNiAsooeQSeXcjiD5/gRi
dfGEplJhdBh+OXQNegWF16XMPiBEFqffP1QcXmdZzfjNtZsx6ptzVe2EkaYfECzM
kU9udJjHvfBEuC1IaZ0TeGZjove7c07ZQMjbgro1QWWryBqzNX8QxtTHtkE62xHo
/waTmk2Aadno4p3Kwfb8NoubhZvscXoy5GLp7/8O7I4wTRHDorTq0v6JHQIg3eqN
cg9NblHugF5pLesAXwgYaOjggCviogE1b84AAl7KO95s2kI+nC+2Adx8FKwR4IdY
s3cdqHWgIJ7oziSC/mllB4ADq3tYHKVWix5XZYLVV8ot2xNKV/JBLf3SEvX89FVW
b8nCTGMANShpPP9PSd7og/T8P1cQm2hdp4xpSZzEf2GRQUnnrp5MkjmmrWWnI4PR
IZSN10IwGi7YXiYyL3DohW6CgLRD4RDEkut+l+vxWeVuEAddA1sX/P6Awre1lT1M
BiVFLJR0jX7Ls0K3oIiG8QUoRRPMvm/8225nI/nW2zgYshPkQ5dd7761CjD4YkiR
WvdS70ODUuuIo+Z4L1zYYBoTypLTJ65ceB/DE/dNNx0y6TMb25G3NDVGUo9beGj3
kJKNYeZzFysw2nbclPmaR/YTPNQ2CvFZXqEl3UWZkboUaQEm7OPw/qF/g67zAaUx
+AWLe0T2gPIx27mQhyHVXAPH01MgNo9KvNXS/IlnyqPMhWdbmFpxgfC83x01njFV
xS29dPy6OuXbMtsQosJzZuyYmhWnBHknvpp89MbpqZzR4wC0OQtV3FUAgbRMogU+
14Q4Gf3guOvBVFQNbeP+3MspdAR0rEZYj1ny56hkkF6jQyEgGOFzaE59gmpyOi+p
zbtL7oTGPeDvprKE4BXGam0pRHgMduEi4KB4XzyZuwKEDcsLOvw6vqTENWdBXEPp
golK66XPEbxM2n42A0Ph/pU9Yw5VeV5QGFT6iotEjavy2Rgs+0KaoWZI9Lq//Jr5
vkGnUHf2OjCbjIt8rRQjxrSaobfxdBIZowKOM8M24MLUIz/GJ2kNCyeNItK7Aelp
sIbXe1HHQ43W9NiOCcnZDPJ3CrL+BFDchzFt11BBIZYGBdHK6Fj1LDdrolpveXfF
aB2mj1zMYpNxVfv9g8Bz4FQ2I5sRHW4jf3wJwZObGrRSMPNHIoXlpJSwjTQCVwgb
zUYnkHK/N++ygcrRIx3e9Lw6dxcPofeJ/1hV2qYnWyTsWBndA8kcpvs65R/50GNl
JtB+2MaatRZNFvvP6Fzx2ubCVM6x5O8gfE4F+A4x3T3xnwnDmL8GRqPcpV5ixFVZ
NBSLiHIkpisYMfRiUXa0HLPLtLGs+HFq8Jz0VQ/Q1zFMKBeOAVPl677BCaRA2e2w
Zi5shdri5lzxiSMOi18v5HSEptc3axAK3a7z4B0Kpxt4lXyEaPwih7Xtt4xaPl7R
xDMJ7f4Ow4NtKq5slq/nHpRxGDdJmVJTk31qiO1kDsTHh6J0FXxzloyYnXx+IB/M
gBl1UgzYilkDh3+OUIR2Slu8tsHc9AAlko0BGksQ/joiEuZmn9N+mulhrxr3dYS8
kmtGsiIfMQXiWW5Ws06KWHrjH8z6ywijZKyJNxrvXk6lIqYFxc3mUcSaVWquFgNd
TeEe/RZkLIWqEUg7+P6BUuTa5s3sLphEWCDoLrb410pULQ3KFVNH3bF/AWYWiK9Y
LwK+MKvkLuj1mg7dv5J/ebY2OjnO2bHksssh8Z8Xh2fDgLEDNvVv7i3Qv4dbg9Of
u4H3OVRzdX0byLUQUbXpd8yE8M3PDIhafPobbbQeFp0fg+wgDgxy9cVpBvKmIqW7
LmSNWBOKIZTo05b88FCsgxCCKGzU674qqHXDz1hebGZpYWo9Bb9M1WguJB+btkl0
JvIgtsrLAcFxsqlyOk6A2oCJx7ebb4/wJxysvIRtNaZDLlNXJqVCVKAwTjskomzb
0zVY5pRu6/Uuw5Yn3R7G392QB0aU+0DB7P0pg+y+770ZhvRjrFQxjKYQhi/gUrkI
S4lye0mhdTEgf/rlUzb3QIIeausQE+vLQvDV88Mbfa/pm0VPhbvZt7/48mbdmA84
xDGUWHqfZz6vEX5O5ZOVxCKdKn25dtxOzRY/5y6NUB389MNweknStiRv8hmH4eIn
uhgfI6Ym6/nF4QphEWcZSLL2xOCPLovCavDFAOEKIyR3fCENBYzRshPAKmMEshpq
lQB0ScYDbv/Kuh8PAWT9LgdxQQ05Uaoa4aLNTt8GrRW4IEe2/FffXGXKfVD7rH1+
J6nCZaA4AVVE+vw0grY/sX5bae8+Arb2onYH432solo9rvruZBSeQtrKKVyeJr+o
IJwMPFn7ST9RKy6A6Q7aMlDmW40jipsJ5Tcz4knc6299p18eayUkToar5esKCVSJ
pA1jx8ZtIzQfvGhljl7GcaPCbPXXUvdoXsbz2xfFWJL6fUw0B2rkihL/KNJ0REaM
CeDJ10hYzuIHdhh499MYuPu+mAZMLgLnNHQ0VU35PPjPWYy62vmcYbdAz9FjhY0k
rqc5SWa442vmeGndmIyfxx0VmIvbe3x0EeTwKhguXefo+WKFovAW63aH9wnHsjdb
yo/kkhZc8P5A42TiYQcTQtziXFnpp5oiJ09IXsjRwkiAxffgSoZ0GkWFvTBU4GQY
TMDyrSDPj8cqtkb+TKz9R4QPk1lAWbmRyAnucKrYaCmEwspYaQlqL6NdrtmkO6K1
ofCKA/AGsTjzG82DKUp/lN4sWWa6ZELvh6pNSCx/W30zfjrSEhvSQHUhmW37AqjK
P4hCpFLZaNE8l5M/SVa5p7fyodMS7OBpyeiV8U98bjPiM1UD63x3i/3YJQRnLae2
limOJnDVArP1cZEePF4OaUdjE+FiLxOW3dLkbDlC0m3VjbPxNYUkpIMd+N8prsLp
hHQglJriMV0k9hwFKeQICcSrp7nONWi2CECFUjbkSfrobZJi8rjpMNCN2s4lvn9l
cYuTY6Dx2BNp2vrc0Z+y9j85JQFdThI3x+lAHHD+7R4k3ZaRJScxQiTB7gQzbL0G
uNzIOteLXfqajTilHiiGKryC5HgSTCcHs1lm3olGdkhOVCOsjNtUWB3lC2T6nqgl
lukuWpB8PU2WUmpG9x65M+HHTXw9VfWDzJxKLY2wubhk43lYR3KVLepkgaaoQ7Zq
62Eeiiyp7OTFkwmBKzTSNdzAXDc7yFoHvl9OYbuHKBuN7om1b+BPIVZsGg36SxXY
scwKafRzNLgF0OTEeoUKH7EJp/8i9sRMHWLlASH3smh87lckXRZwQaaSICJfFHcI
QU7T+Jl2PdMEM4y58RQcLIxSE5ttP8TkoIeC2808VZTQVyyg68H86tfxVL+LzpuF
7BkEYXAblhDNhU2v115rhlJS48rRFvjc0im2C7mMoalaPvum39jn5gJb6FfX3ixB
NpSw4uCRN6kpuovCUxFvn359C11vNL9/cgWY1wjPqGnFjUdiG5pKuuMZTyQsK/gf
YWjK4SZxU6PXL9X6SHRdienwXwEoT2bc2CM1xOVE0bCWOTwA59FZP2qTgwl4y06T
mtiO+AS2DJSTfzy2vQfid1qE0lrcNcIfGw0G5ZmZYU8McH0lui9E1K7l5ZdL1eu6
ldmM9FpxUjgkDKJd9DJxE8vf0Vdb6++5UwjQuOoQuqOJdk7iwc8zeoLbGgNHObs3
X9XGlf+I4bprYQquDhxPEFRnmeGQ6p9O/C9BAsvcYnGF95gw8+Bu6yUWs7ppG+1U
xmxJr1n5GB5XOJznKhsiyIBw3jYW+DnMvFq+8DbeKXZMhgA9+SMVclh9FOfqY0an
sy4hZZBDznKiKHagntpbdk5U0/06pUtpVHmI1zBZoLpm5eSyPk8sfDotUs34pii+
sAhOOsNkkDw0kBb+jj2OJXitkeKdIJSlpsTf3CQonbauLWgMEZUIHIO5Oz25I4+9
Sb46J8mKg8jjQBgffsQCC0RAD5wZvPLAh8RNQtTDwYGnH0QsAZth2Wmjdktt9nAh
KUNudI8iwUqrMsTuSGK9Vw/oRAfy2L6WxFaJ8BMcIsrljWh9gvCb3XN2F/+dGXGk
uHiijxrG9StGW0hTwjZ/qKTB4EeSlDaXjNMxK2EKU9Y4SHvwrvppTvaN1SDbLc0W
qQF+Vb2EA607NgFHC6ljlfvQ4XAZzHoDUut+8sGjn6Zo6F/zWQ1TM7sYm0SFTcdq
w6laEGOpVP4ZJfHhZFw0aGQKH54jvmhssoQ6b3V3ecla/9u9gmTN7DNDmWqJmqsW
ycFd/g9c491NH1grl9YuR0gXGODL97n6PqQAIlN6wu++aPztVKLqnE2M6/jnUC4S
a5dbMFE7YtOedrYVBEgJyr+Dv+XZGK1T8/UhR2hzhD+2jJQUVtpSjPUtfC6i6nnx
tGuZJ4dm4FRZMM6S/j6oTeE7lMemmuLqMBCsKVwVGksiDVJRL60RJytsSc1gb5vC
fychnN3FbKycEyv0lQfxaEeeJtvuVcWOZRbberzRSqsA/MFX8dBOIz0P4Zo4BBh0
9uWMMRiywKFOUSmxaDVXLsOJE+Uec1g9ERKQ0ieSRSTw5WNjRHYE9N0ZUCp8d4c4
ClCGMazeSwTqcwXHcZritrIl4i7V/IcZfo/NfZnehdDChXj2qvOMTQnWBDQVe0IJ
aY/2jFj7lMzpcU1qS6sbpqyG65+FaqclZNWv/ZkubOCRdqpJVaFd59/rLl3xKy87
cBl2ZMbmZfGaEFUnqOe5HuNfdpjq1zhw/B7dgzdvEgcCUPqpeA7jjDHxuw4SuT4A
jqF3KYbuAU9bZISJaYPgmtb9+p3iuFv7IpiT3XdZSycw6z8hgcruLvFnCaMfP7XL
IaVads3h4bWgUUliSelQaRr3cc7i834gIxUkIwHlPj09xRoKCbsGlpt00uMhjETK
AbsTOjvgGID0CMXbfdNy9dUGrOQeAcdwvHwPctmLX+r3AMVE1IpgZ4pc4lXia7v8
Qmn0c/pDHTAPLXmscV3wTgBDbMAYSEtBn1W7TwZ9hqetu/W2Z5xnFbwRUhvAt6SA
skkAGIDHikC4+ustZ/hNUqOLh0NU8bWGGxWQbe27Cf6cHWeLLPUmUnXqonIeZ4Mh
cq2YG1DCLpsvCNAfzGK4wxyJBa4HfbELqoP2zbeHIeLNKgMV48xfQ8bD0l6TOtcQ
VEDVVWL9XQ6KanbEHKXDZABLG7wbuIKy5Pt9p856TOUjC93brUIqWWoJBj2Eqmfl
ESehqxLnSPfNNXZdqXZi8ISwx+Tukk6Sv7ycU+X/PHjY99fgDZA/IfZBSCS52HlT
riynlN9U0K7VbdhJKe/s+I4g5mZM5mT2XOobv5ob6qRgPqgCw5dQHbZZMOOhnjvr
VvwcyFgCPwvm6hXCOqhmTtwbI8G2lJ7mOnIH3MHJ0l7hP3G/rIidMeiZeiqXfzQY
hT7yiyUftBwHK/99tpHGZvnUnW9h6CSeSlMI5vvehkWZRbV7MSYERnvJYryOrEhK
Z/YIwQaDrUKvqibyBoKl1ZTVxYDLg7+FFY7tfT9HVKKdsJDiH+Cm6lbSnvBRYwE3
9dAZI1PPxsrykJ9j55wcfjWBtWE+7hLEFXwu2T7rdEujXy4r9KpFOE5OYqbmvZ98
8GfXVocdT93zE/AVSFFSMfhll1tOJGxDV5CSZT8onkxQlnC6kvhmLLrylaYG1xWY
lxsZOz4FsK84SLAP4SLX6PvRfOtbYMTll68cVykQ+J1ByNQZ5leE+0N6ZKVW/wQA
qU0DDuz9A5HvddJ/CWH8ew==
`pragma protect end_protected
