// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Zagh+eXdtxLr+mX5t2d6MS+QgdvwmTHPxbc0zDTEs9xXxyL9M19cehXPn5mjpBkJpvnyxRm8LUJV
YmJvWEcWql1ZkamxJ3pQpLbj+BJ/b812guTyDU4Csxjmd3ifDYDiXddAduEejPaflg/VrFBLK/4O
5mGkESO7LyDQ38Ep91dRLx9x0nd0MzJjUZngPupGjlyMLk7/CeiSk1EqWN2q6TjcHdkRsobIPAgf
HQEPy9u9x87Xpgni7TzPXTXlcuBJBVkz31BgkpmvdC4aAKmqENCKWq2W4dMofNp05+TBlP9YYl62
EdrFcQJU9ofNVZ6c25RJIztMZ3+d9GbStmQ9DQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
S4TQJ2USKYWG1BuOlxM97ZUcRTI+yGDvLo1LdytWVWQS8W1wxEm4bGiae3iiCFhunVi8vIfIDQkJ
ufbG0VI2oHBdBXO6RMUXxdxdWyRPl9+tTphBzvRzPQfDvmESLwi1qDV/VXHOE1eIMe8Dom8m6c8h
+QhzObVC6D53nMClW5f4KiIRfbOPC/JN0vCD8+6pKdalJ2zbhNvvGQ9YSo6CCPpd1NtgGhiOP7pU
HSW6ZF6ef5G9aFKfWRYtOMl1WYehzo5AdaibUL4EmA4dUIt2Y33q+pCMHC2XZTmgQA/4yYz3Q8PO
uzViJe/v9kh7qBX9kafyTOWOKAKsYsvug6Ff+nEO7HLhx+D2YXnYVXxI1/J35R0BcegTzOCwTY1k
VSUj/T+M4afOgoeN/9HAWtZ2CBAKYNE3BuKInYK5ZPUo/Q3PNlg2XM18OWUw8pVpakfjnmXMawRf
lMLvPfqHnxt3rqcnAJBwd6SEg4uZl5WuzuT72S2mwuYcsdFQytcRBf5ZeGEwV7K3jc2wBk6aEEIj
pgzM/mM1+Ekfo6snwKn+9sjBN2JQX97A6gsQupx1PQfGwiUCGFsN8NCDKeT0vsZNdooIG0fR+Sta
LnuzGGijajf/YBCdCyiKHO6rbf2SfxitBAyghjylHFV9Pt1qc31ZMMHNwMpkW9t9oCzO+uYw92Ii
2XamuEkLkAcKFiY2vHCmoKtn5Q2D0W1LBspOcU7xVqsmgpRb1vyXXWBCjSR8bb+h6qUv5yaNDtfI
cn/6gmwI9qV5sxiasrE2+UBsfCYU4jKDxRclVg878vSfEZK4DAijM1QuEFnCts3Mzs9EonBR5sCr
2u3t/3rj0cvsEQM2Z2kOKmmNCcAMFZKgzOhOoS0UpPkevwyN7JPpRZw2cLFZhIvny89U4pGsUo4h
lzhQJ5ZcszurLsUjSZtHUVgFkUGkBoysexYduZreDV8pca6lhJ5gkp0GME2YehYlmDEyKHsd56+M
w+ZeAWWsIGCeMYBsM/DZ4mev0RLt+EyR3ZngV3fvzyNrZiD3BPKT5uvgyRaQ4dKU34nLQzXD9dO+
DNghbxVDNiu5TvmyaY+2yfjDWXvuZUiZLkHUPKyfN+9/u4e0ug1AR1d12zo/ygGmLABu4H11Ry2R
2r5XEyqu8hSKJhkBsmsOga/Ed+v1IxWbIZfw5P9+YhAm+xO/rCDo/DZsrD5B2oejTxeBf/NNJy01
/JZSur2vG/w7HvEASRviQlSnydr6HYgwbTjun/7SVhnMhbVHq6LDvATVNrB9em0l84+s7w0O+UTt
tOTMnfUq3UkKBOu9Zwgk2DZLs6VIwAXZzt59qz2VF8gbiOBfEbGb+C3ecj294bsqkTQhf6E1202t
nAlYt91fdCgvGkkccQF5tWPddHxO7tzw4Mq2xLaFhU0JIgDDs/gT9ANVgin9c0xdRj+KIbLEL9ng
U/VL4t4blBLAY7Pojnt1G0c/SaA6vMmisNHtDSyJWYY49u3kchFi+YXnYt+cDwG7YSO0F6dOMrT9
LNR47KE5sqVlX+TbZl0x14nPxU+hEh7pvFbxnhbBtqSCVuPqsdiXKfSbyRqUJHImXKc0FHxQv7O/
7J3QfJlRczZiy1NSM1BHUWcy0z3dFKESEG/pKBgPwu3UzR1K0G8zN8zmvZwGF1Agl0TM3/ZDdWLq
UHvpn7f1CfZVEGY+3djrhvaDxgNyNGElhBzdDv0PtEXzouSVq7SLKY52y3tirfCRvl0ZYz4mLL+p
vm6tgzldgAIgD62+i6+H42Cg1srCqSPo4ns9fG0d+KXwdVVIbEr8BUL/n+5t9qb489wzZztsxS1Y
3+yHjJgNoDLz9CHlM7Cb+UskVJ+AXmskOXthrso4P9QKoowkhoZ0SbqmFn8XOXq3leYGzHjewPYT
aZV23lN4hICRV1coYU3y4oOu5k/u6hT/FR8xPwpAqLMeFr2bK3zy5YXNCZu14+Va9keAOYF08Q5Q
fq3hdBb6Eg1lh4y7Rzk8Fj5mUs0DadjhuxfRZAJOm5niE88HPB6tMJZdwxleBKP65MgYXqdu685D
YdmWAA4r6K6aPxpJAZHt/cgFafRWRweWASAcnz0kygLrFOVgPm6bvFbZ4O9NFvEmWtfbKnpEM2zm
sKEKa4ALwZr/Xy2kogcimYYy2NVb8NGLP/4zECPSTpltfrbzdqWWfgIxjxkv07GZkkKrZkbWkFZQ
0GZAD5NrbCgoN+0iLW8lehtYL8WnWmq+R8aKbpuN2V2cIm6WPveRZ7JRImepKmK5mLXkB/HBRdgX
CUf1qmXaY8r7/Zwh5deRwSsCGoyIoOum/HciTiz2DpZQhwhm0QhApVQaWc6o8tyyU8Crg63xsw0F
l7G3Pqkug2ahfm3XEjO9h6sr0Y1NofgHxnC2nLPVxIxy3a5W6Zyyd+jRkz2viy1j1QgS3A7OeSNh
BkbwdWAkfH+AIqphBRp8cui5+XHpjaCUVxotWzrjs2CU4CvN5dOLtSmi1xjXYCg9dwDBEM6leciz
G/oYDBxi0ZKZml1vp9zg5gcFM7Z5wf8DB4bzU1fIqo1bKlZQ01Wkhkhjr2rAyYOPBNFqzCxxRjxR
i1OF7Z9yK69timbhwA9bkSIH7GVOeRLK9Rqhvoa8TMQGj+15ptSS2Ex5JeR6Wk3p9xg3w+yykAt9
Z5V2ku3txUvDwbnLvo+tV4WU52sCqZUrgQrXlI/5J7c6wW4M91rBQVHyo/A9oYcDyZAal0RZ07gZ
nKkL3kUacS225asgWaGIL0ST+9BRfUjN3v6vBI3dpd4FPBFLRUnk4evA+fokN6TiWIuZDAtD9JRt
nNzgV2CZO21lGs32eqa+qgW+vjFAP4vwqyGZ0DNMEIhI3T7baOibmOfpCGLvgkokDsN+Kr7yDwk/
ZVPf1XnJf3RSgRvHCKCIxKqilLjyikgUioAkubBXh1xKUYwmzoPtwx+eB2uVUVni/iXhHrctuNs/
mhy8++EShaCR1GzejF2ScAUPzQRaowVtllwvv2R4UoZPMib4PrUw0SiZ16t8xWAOeUHXFgjJhBw/
aEUJbb6PUtV1KXSui9eH9HpU/HQllDGE2Cm43RIzRM94VDgQrZmqbW0ldcGfNlTKZyjeJHExfvG7
fHRTo6HWjxQSC1/o1u8ZuDoIpRfixyp6WxvFgBX49HIEzDwBY8IbRUCPb7otqf/Se/TN2yX7sVjh
8cHnoQ8JXt+rWzbcqaLKWNb8Aa2ALdcemR0B9oQrd1miIOczjSZnLZqGlSIN/wG6dlnKWvd4TRq3
p0mz/21oD9rffXwlllOrSIIojhmodSgySbd3D2AU2riXNzTJi8/vroZrsezeo2yYnM6fVGaPMkRU
MHVUdZ/ggMBe6dflcpa76Tzmgb27gKFVvZCpODKyWGAJelUOxp+pupDwgM+dn0iwkI4MPK1Hvm0B
MWtyM2D/dUUgUWS0ETIqdCHTWYZB5YBiQQoTufLYCONpBbgYEJvV+ww5PP2qNJgunA5AQebdCLj7
vqml2x1esuEdUzYWte7T2lJwuxCalM8FiwTlSzFqBiGxc3vPXzrhxql4IzwLVBN9d/eQdlA7SvRI
pwStVvmCCKmF2H7X5UMm+c+cA51SLP55eEJQsSMlAPdyIA2S6Q2BuvIyVfs3jT9/PR9sT7glfxO0
x8tFmx2MuPd1UeJ0c8F+P/0xEyto+UUKs3v3zGPu7xBrh1rXH49XQGsVhi52LlcnF4/aziXIuIJ0
znR0WvijAXl44ofDPH0knkKXb/S56nDOES+l+exuuBjoR51zoy45IlTK3B9dsWbhzvo2Y5d8fjU1
7+wk9w/PZqc+N9cY6/0Bnc3HJliDfMk1/KubTbzAAxQauCcw9BT/yPxY5jrr51aGha2HwSzUmQ1k
Z9bsQ09Tb0UepgumllkMhsT1q+8f318jwU63Q6woJJCF4XFEtaBkFf8yFgNJcV04nF7NJmMwglUm
ZSx95eMebiQvJA8+nl97bxdDyVyu92zACMPC5ITDq5FHsJPCl781xuWx1Ch02Q4WKIWXzP3MiSUp
wFcJ1bHz7X2Q6+Zr6wFP2RE9fYDQf0HuG+zVBr+tsnA8NR0nZ2nQN860WbTrM0PD4SXK4uoq+/MR
6Kdcg7rSUqFtRNgGosqYCBymlCz64y+zFoSCopZ/pmDcZn4sxpKne5d3SyKx7+5bS9RDaHCTG37F
sRI0DX1UcjIsyUtoq1s3l83FTQiwLwNntdZMNHFoSUnNX8mELwGNOcEWaHCBEmx3rkcvLGwS2n9E
U1Abd2R0+krUbcpTgwdyWvK/OFtc4KDEUahmgGmOYtDGPjeF3AuLz5tOoonz19MZnguwDfvMrnqS
YlrmsTX59gUdrl793MvMdobrY3xgKGJOYmqQiTmU7cIJ/a6+i0SEHlnC+2PKJA/US4fRyfzayhUa
AzANjlLoDe01FLdhTHpboGILxUeoecXk/8VCJBs/FMY127jSVunuWqaI4nzDzSBCN7MfMfVIGR23
jhZu3Gfed0jgiX8wfbuw5081ZY2tvr9sWhw48XU1KSikpYWgnAUFI3GA7/+qWU+HpdB4I50sc2a+
wbFFjvvD30Xyotosd2KBSS29HtaUORhg+JS9FZUhbsOl4N0/vz66YhQ9xT/C7fXDjkREzMNZTvlQ
XwehRrr04TMs6PRVfrOtPgqJRbjfaWyyv/d/BFeReGe39z6FlbJv+7iHMz2PapRgD5v2J8aY/PMm
mkRUF28yCYMZKthmS9WCJfiiRMGdrHuGs5j19jUcU/TJ+hSgQHWZ1NLX/JwTHfz8JYbXo8zY6NsW
TDiDNj+2HXNmO3td7xEMS1sUwXt40C/oMs4/F5hORAlpAt3TiH/2SBLD6D/mZRuivrdMkXEib9WA
APrrC6bct/NZ8ZxPy22pkckgl1lB2fqoJzK960fK8sti/XkJHJfEQainEqiuODwHqgQlBrB+q7Ro
ovkgE7JipoElU2jfq84bk22od0UQe2zsCSNUVAs+9XB4xHcTDzClH6Y/wssb78H+PyM7Qo8bAwep
XtdiDDVXK1xZsZHDKkaJqCjNHfRBDd/VllH5kDZE+a6TGpVoAPryY0jgUXaMiwzvAp+y3p6ucKm+
AUoiqtHL+pQelOkeos8nTI7Lf0JF+7N/++B04MLulPPEuqbFEjwlirQwe4NPuEaY7HI9OBH4york
/B65KX21nrDG2srwb8CH9qVMLlv1tSZdFANKFNwADGn2SI3bsk2jhH3t9M/cz+6m7FOBAsHT2APp
8qp7X9/c6/sscpDCsKg51MBmzkbETF6afP3pZDTpgzDanRRl2D/G/uEesYqwQyxwT0Xx6EdMysXQ
MEv/a0jRZoqwAaHChAnH8Wg4ML69lYavvGjMwtcbhcJ2/TnVR/E9Nb7Py201b8gyXn5Bm0UHrswk
vIECzJpEVRX8cxSjoY+GUDBpEAKNpF2Xhd5fNrfYuwDbKrWXS97CGCZ5G8+R12BbAdi39OShb3GX
59BcCc/nflIxlHF6OnE1s/cmcoLdCbt9tfopOiHp89wUiwcnjIgAAqcE5/+1aS3M2hemtvK5EDBI
Sr5GmDMVo84ZTqY03ITJYYSFrOOZJyx9rD9m/6CwBKuf+m5B+P3TE4iRbhJob1q9akqYeyI9UIe3
aVvVO0fyA2jTd67aJEMFXO8XEnCd8tsqSV3p2syud0CHeEMfMvj5q0SHgyKSqRqNZzIO3EpdHijf
EWwcm5tjPvXSRZt2iSsn5nZ18QS7VVAt66KJD+wqd6r3icXy0Qy7j/lbMSVS1tGFjoA1oTNq70BO
o8ANs34wgWRoLFjvzDLolpuH7LWr9RBR+v/TUe4LnV7UJ4vhY8sTwHn/25Cl5fEcc8N0iJufT36J
jeL4kiU5wCnoOgDW29u2ulxy+3DowKiZv6G84YNlc+pjg152ZEib8eL2NmV4dMBxFW5o4DFi+xpK
INg+Vu4ZSG/MN9vSZ2P/grutpua75ECCqMfdMEuW7J5KfXI885OMxhsJGvsbl6t4J9AdntWybhAn
D4aev4yxNIwWBDXWaFb7PclFUzCUWY/7sWOBvksystp88j0g94Vf3REowIxtVpJbLnsQpPpLj4MG
XKszFjQ2MulFItEbbxXr/LfOP4eMkwRNJ+OEZu9T/il5NrYW40p8OVg1QXcNX1DLBxWdfcgqzYx/
U/nokTRaDNY1I5KB7CgP0oGS6m69B8qQPqsxeAAGJK8umcf2PecMi0w6vF2wFj7AYOYmYSOwVkLm
nmLMIn0Hhy8j42/Tfgrcl8UtH1hDqWDvhpRDCzPU6ikMebb5D5lIXxnQjl6EeMFlsMMrFfs6c4bg
IhY1NBstz1eZFyTd/HO0GO4cShJmHmly6SKeRB2C6Plhb5aMb7JwDdCfIj8OzCKZaALici4/pCqJ
IOke+c53Bwac9ds9qMffrD9jm86hsuMkvMA2N/5a+8gah5eK0aZsSv6vYaWMhvd4JM20kUMLpJkn
WcigZ2JCvwQ0cwgCAZXYiqlBCIf1QuVBcTI0AGx1Cp/16Kvk+ZWam4kaTnEhmObx5PVBOLnfipig
KdPwWB2D7BxlhQfGZ3HyV74NLxZe7HZ3iyYzHByTx3qaKAAjfbRx0P46Xt8dkYgliWCRXz6qiJDU
xlwyaH7TizcoEfjXSWTA82JoyMy6yqEFgN52koGjB2/gcrFCasBVzhIlWVyP6yEhWCIvOSiuN3gO
At8QrHaW1YvEC/SqwqVN7KaSe7TazxN9o3RNgIg4JV2ZUaKihyfiyNkwB0F6lJMePQY5YyX7tS3z
8GkbCF7xTTuHWw641wuIDSDqjNWiuuhh7INnolHQ0ZDZEyYnsikSVSYbDRPdvyxuc3GtJK4FfYG0
H+WLB45PVP01vQav1PuNBnvo6SeyR/DCJy918vrb+syXz2DVDGvCQFpQ/7siPPvT9kiKuHGZT77z
FnMwfAD/WfhXAd5UVCH4Hiq/jxlMgdWpEiHYQ6B5UnfHKrc0HI3E37RlIwRn4O1T0K7xOaYJIZrv
xMO9a5OuwrRoaf5Fgr6RvpmG0mp5v+3qClKTXqEDzU9v1QxvLx34/48IPmlOAtq9KfM3tT9A1qoT
QlTi+gQnAqS6cO9jsmOM8F51Vu10MdO1h4FEoq8lE1XIF79kOgO8wTZHWc+YB8slTj62rt0J6UUq
FOMyKZwum4vf/N/jkjpLcSI8Fpv4O1bA+90jEnwyOAAVIj/sPdKoVFR+9iKxjiQd87hFL8kDogCr
GxQI4+tOZT6q/sGPJGqSm1GotHw+EafPSWM71fcC1ImCd0rs3K7soAXyCtIspUJMe1sS6Nscoi4+
9wXIulabxyhn/DVI/xtSIF6Jmvo0UmwCpyouO84V9oaXquhGZAZ/3sv8Y3dJ3VdwmYSTRH78pJBr
7nN42ZihQYF9Ne6D2vh2hBNuCbQEqG0Zrl2+gh1w7fi37i0VHQoEsijruYQxPpg+TrPOZINLOQkR
+UEp2zTqiACpnDzu7YZRmHy3p6BVM9lwVP6mWOTawvrNo6LF2TsBEs2CcUaJQTzm/xDxUmEMjgNP
TAqLMuy6AipSBGx+pN/9a2KSPdAGu8u95i52Q3IJ+F8rgPOzljOX3CZXVuXQMfyq6Pej4WcAam+k
2pLfJYXRbX4QK07zhUBSn3CtrttkT/8zP9/ydTX2THwmnkBme6OlsVOYLXPoT5cNSrp/QYumduHT
s+RsjD+DQA1mTgY6rLQ6hSRxpWsxRIm34CBnwGmpBvbs9/VtBl3Ip3kVfjNv8ByVgMLRQZpa6Yro
r7qoepvUZRICI2rGBZVLYNE7dR9RDz6nXhfbj5IBSvx2/BOXx9KOtuLXs6oJsLEuvSa9A5UuLH7h
BcoD/Evf1psnvcyPEsaClhiC5RDWIQWe6IE71rbbSgmjxKkY8d2Dd57H1o5BX/C95eUQT3H0xA6l
cuQi0YN1iZilFXSMnU9HxSQAUgGN7Hb39DCuWmpPFoLnbVW6MOZ4K+9a1tEgIASYJN25xnE21K3Y
qweAkkG7bYbY78ROjF7j5oNIaHxPEXwvpxUP8/b0j4HGGOH+Qm0wVrKkqrRytqP0Iv2f/CnwTNKD
f1StBZ+eovlH8twP8AagbdcitZFFVfcQSK65VqPrZ0L536BpQc1ywEuN6Udv/c8it9hXwOZC6CUF
E+IHtsZjHI3iltCoCy/gmPvn0jDcJs+q26OSxux+lcYYmWodkLtBs5sJ8ydOWahsHoecFkJh3dg7
aCSM4+hokQGsdNbg8oEsqDNJYd9a/VBlodcMFUlgEfdNtTumwk8jWum6ScuIlaaYbKFZMk65FyZ5
jYF2chr/FicBZt6mz4BZnTrpUluJ3FHb62Hyw9t2OMTUt5nMQo6geFMfQIkFfoYvVIuXjBrAhf/w
9cYY9UhZIHbCn8Wq2JWamkcZnyeldhsTzTxErhqT8g6ITK4PRr2KFY45fmsFOXW3RxON8790yj2O
6ccuENZDHfTMHOgxgRCKXNFWHdEtBrB5bqSsTBQxQfVKGcBiXGBfE6dLsygEyon5I5xmBmLwFAj4
rQUwYlypGh2S8FqznkesknRbpWaY/9Vb7xlMMcd8loqEp5eHLPThFkjDRPwFmkt9vRsxYipE9BfX
TbJTtZNkf0vlJiJQsob1tV0YUqDIdSUvCepmEGuhNXNW4nQCsq4Azop8NenAjt77KEmBvlIINCSp
ZQlSX96aus7bVz5iJKNc7oNUXg6akggNZ8AAViynabH01NLrkoKT9/s5JNNAMQiKO7tQGchqfdwI
D+T+xlZ42W5qgMDEDpZqDDrptg/x2+QqV2lARlsi8Dkp9w0+7osRl7+uupTj+2i9gAxfMIoLiJK5
7O84Rbcf1U7UIs1zR4LuZF3gdnHSYKww3+QzQ9h8cHK9WAIo2ztt7P+uv5hvy/ifoqT4Mpws9AZH
x0koeWIdA/LutmHiHGNPMjCxV0I/ZTqxM9FZHkg0WDfHWDJvFC4LXcwAYNKjK6mUytabpu61K3R9
1N0zdo07l0LV84djPmYchZZtIshacl31kP9dOns6z4QoiOvuxsaFdzhwars/eKj4pJy8/jwU+Mw1
fHj+t5G6KSRZPultOiSnHWHpEidhutrZps28xUh2q39ifaKhgx2vEEzkJ3/gSySN52MPoWmBLqqX
Swo4Q5krIxz0KZT2+HK1IzIFa2SnziFzZai+BPVC58o8PhL5j7zJXgveEJInPOx/KV5bfkzWq9M2
xAL1vlURzOy7Pk/tIj4E2+8g0pJi7ubr92jx96GdvGAvvvrMjAlzUDCoreJBL4+hKdz0c48Kq6n9
9rCfYxcNATJmLkVmOPvzQgOl/1wvX5iungAHq4nLZc+ESoUbDViVI//DXkEjZK12wWgmfh3I8fs1
3WvOORlMyzMvkMNRamFlh3X1ZqzXEY0AQxcq8v1XJAmLy4O6zXlNVHhj7uc/ruDLvgq9NpQEygxS
eO6yfwaLbfl94pG23vbmi+mOjFUtQUuYuTmWbEsfXEnOCJ/lGrqcWiJRetNf8BNowFIsSvabcMg4
RaTYMU5c6j5NI9rAFkEfg5odd5UoRsuyblKHWRjLlJNR+VbMUIWyeF4AxgU+ourxD+1ZdhQdtPIQ
6svn7ieCf7mhol54dGBsgVFXg6BYyoR9dctFA8kCANcbox3WiKrgzidLWmrGL8WqhlOj5Xz4YIza
7Auspmuftdl8Ep+zzdeOVUYNsmnxsAsW66SOfkpvvhhzJJL8QGS7dG/yWuRwODdr0USEeFkO+zem
Ztogw29o/mwV/EAt815xC8njvqexqTy/hIyjCNDI+iPOh3llLsSgh9AEHRGVfYuBHayruzF9+Yrh
IYInmVC92yjGit2oH5XQd2u8SrU5LEFPfIFl8NurqPsKGuMyyUDOc1Bff/7sVjyJ7K4yUVUsuEq+
7i85B28FMPqqKSbtgzJyBf8THu9HEn98Hu8QGqJduzy2Kvqpp5uHIxfaKLuBN+xjnHlnK0Mcfld7
C5ZNOxcfUyoTEQY5Bef7pJgegjaLfJvWWylao8Cxc3ttKYevDPcBYz/DQvTaOdAuS4VVGJjtyvJu
jQfMDSPjgHT6EkJUujCszISo/IftuPUVyFdbeCcVbe9MN/jwb7KmbVfoTgVP30tXcMQCgOZ0NK2I
JIYl+CQGzvx/NJdVJMTUjy6WiTxQk6NIW2zqtU+IvbLXYVn/U9nRWPHl3BjZ3INkXl3HwuyWvmfb
Q1HPeG0aVVAOjVaDMMwLjIzQnch5CfXFhWuMoPKLUxwL/ivyCFRhg4Sam8esTvZLvMBlsaaIBNQe
kToPkiNQt+BMgsseKkY1LFJxAD/keCD2MMYoMd62hP87GLUJQi7MPAYueSTBGSbJLRX8Zq2FWr6F
riAUViH47aNvE2VYLrhQnDGIsLlxYPbSQ/loaIIXWFFpGHVauwmLtgZZtXrEP/d5GAgJTW4Ed1/S
jhKOId/qJNE0Fsh6RUJ9zWeN4g4sdRHuL2UN1YR4rP1VEdnVfHK2DSUIUhNd8lWUAK9tF5CZcGQZ
+f1VHfc1T67ixRK16sdMPFDjesl5iQiKSO3X6QuTb3H/dVm2V8JonQ4FBmbfvPlncHK79GTSWzAw
XpHj9f2wTItNd+FYjkDdmIjQDuioB+QZx8cH091vaRM3InwV4YH/iKAvvMPShjzPypVIunfog4C9
0XMhkVUTAGMAHqOn5gng8lHnD6vCich5rrqPHuXhDziYQsIKUbEBkNPJbfjInleIA7C5sObXcNtx
yetblvgZQS4StuZz4AIt6p+Oy1CmySTe+CH0H0BmgffS/IwlAhFoZ8tbD68z5Li2vFCDw7fWS8iH
NYupkqfNmc9zJt2T8BjcUKsZLw/hITUWl2LKNalnuZhY2QuKkf1fnQE76pzVKs3fIFnG38+EKJT3
PGePAD0HWGe+4ASGvF5S1O5DnylbNpeKibsg0VTJb8TqC1yxb3mn27ML0dq5b1msPBu/GlgPUJjL
lNOBElZYbxWMFalr/ksEiZt05bx5hAr1uIzF5XCyR3Ox1F59aRf/yujpMKevZfoLAbLwFVikalT0
ubios7uW5YbgfLucuwbwhywamvYd8ja9ya3WjVm5J+u26uZ+kPLAe4QZTC2btnORiDLzpPg2GRuJ
mmJggpcxLdNZa1HkDvspFTf9yXbzlMS/aSG1Qujwz+GerOXoV2c2uuVyBkCZ2qeIuALYwF5J89XO
sMJgaJ+kOOFcYvvwVQog0DjRzHcVfh44AH1cwoFUuGtL9+wPHRLcPOfd8E6q2Csn1rPfapcQAS6d
entiMb3bjrfVd7HtKXy4tgYma9HR51ZrUivUhl64bpBS4YI4bKMc2QGgAdGCiO5rf4/+HWMKFbNA
j/GuriMGTmhVKC5GjTMW3WEPUXdQeneKoxzkt2KSuLCEv7LpGfUsugJqNOLooSfZWeikulPvx6v0
7/TvmrNJaiKgnuA9wRhLgRvMRuSZc57m6ACwGFs/p6OyrS4DppkELKoq20NkfVEcmA4cyEKRYD5y
p7FrvR4z7WAENYF7Tc/OZ8//5XwncCY6ZxCiMWIsU4wZ93qnX2IgJz7Hi9yuJBvwVqhtlBHluyQ8
xXmjn6RocioMXJybBTzo7KkXKh6/N1iuSzAlc4PaI8C42PTT+DxeBFWhvxfUsIjTvVrYiuXXT+Vp
+ws45sfGMvoyV4ufiQcY0/Ys1I9ymPvy4k7UV5mT7VogSaEF5F2FM/+oynib7mIDXEVOHIM00oly
XQ6zvPmRooQfkElIbq2sXQTjCacoRBHQl8PwsVGFhFzy9jwgxqpn4JBwFvsQM14o+waiv5FTjQeL
T2F2X3Yol2pNz4THKyNRydlvnAfhcjYIo6/6CE2vkN2L0z8QWP5iSRyiB/I6AN5oIgt3h4keJOLC
PAEf/WMgoiFUYHwbQBIMKvpDzGjsGs+1gKnhZWPTxduH/hWG0K3FGOl/E4Z+lHtP8ADTCZlwjOJk
vOxwMuje+VZid+udAV2Pv5OxvrOLvdr4abR8EtJ2ZT/v32FhkMGeQ3nk9IoMGoHH8vvoX6zG4WBm
o4AwOyL65ukoB8msmmUACrJOvSC+MzjgPf+lsNScYrCrdHJF+3D2CQGOpT7md+cWhLkQ4w//vwNv
zUmUkA/ZqIcckGwOpNP4QQvORR4dKtiriIDG7/PLFgwQ/sCSgEZfNCV5I7KHtR3n9C+6l0AAuXps
hk8AI4bEMwYGRcYToIdWqk/IBj6hMwV8madaZCHu9fXf7W2cp9JrnP09bDPVYwtGLID31vqIS4hn
UlB4Ks+cXVjS1IERDZUmweDgazyX7ktwMNx01EZ1CHW9LlF385SKI0hRwUwS1GNcisiVfAwjLFpX
91wlG0sd/dAlF9BADNoarptkR5JZPzu/0wME8m/QjfP3xTVBvHnT2lKFIiDkjJemAE8r5DhHt0BS
rv/K5soVHc4a2ADNTqztpEAEN1NkPjbKJ2ZmLI7TZsONX6aQoaT4BHq6vaOcaYAsiZaVRiOzaals
0PevzscECIclXlAIrrz3E19MNURmdTC+pjkn1BT77r+99Dwp6adg9/PYLeOo6eeH5dk/yvQArjLN
3w589G9cC1FAmda8BkysedmkVKFjm2MGg7Ro0P9yml9IinIy2Ye4yLJwfjYrxY2pGaWjn+lfTbms
0lMm6s/ccAIiJ/bfNvRW3AKbj77ws6mWInwpeKGbBvej7JivmzbSmcSgWVx8b7wal33TOgaX5mnw
IVU3Q1kr9YQNp+tDpJuzpXiXnWewPpvMF3bXVgeK6luoZcubQyp1FnWzzLfuw5ghhC7u0Jsj0WP8
fADJaEmJzJMaAjWBMxvHwZ9dqbaM8WlVBtnTBOvnJh1aVtKFw5uEZxLVKqCXqlhvTMgg/kb/XaWx
OAAZ3POM8r64c7TIzw6CLrnyqpuuGG2AxTHc3qDetl8XVrUtA8WrlKjJtftWGvKI0E5bsMF/VnR9
qSCAVao6egthiPhFV/aReIxe+ZkYG8Qe1PaWnkG/M/dEdjA6feaQWFBg2HDHBRgcaXPF5JjEuY8Q
FSudIkgJIdcCksg/5Ehl+E3Z14wg7Fe5YKr9M2pyBH5StWCfCTIuJtU/zJGjTzgphqdYNO20fnWd
35CCafV85o+iEC88yCHMZORkexAC07dAZCKToWZiGhu7IF0rXoj54NoJ7QbyXWBFeW2No2zAbEx9
a9Qidn9heW56T23o7hP35INsxH7GbzMvsCK5iIGrz5Iud1ZEPaAGK6FklRlCAKY5FUyFBg98GhII
oLrbixZOzq4D9hK5yNnvP1LxlQTLXZCMPLBIHHE/aINq7KQ94YJUI/dytsGXPAgY7O60JauuDDRp
FNMiyiaBSKBTWZzFj8t/dGQTLP5aQUcEGe8H718DQ1gRj0WGEa8fQt6F2om9QD4F0UBhsqoyUiKJ
IlC2QCr2NuCA3F/FN5PaCCxNvP3ayNqz50X7Lt1MY/yQziMNXuCTASopuc7XM72DhHo8jRfqQz4W
6p9hTJfJBbwE7vpsEtPLtaIjHUOK6pNwQy6T26Tl08JBTLzXk1t9Cw6wv8AmNZ4rY8/NxAA1p+nb
wSiuYtAjol/D9r0TDiGQyIKYuvGERjxZLjLZz/R9lNLmxL62IzV/b6U3+7r2+52ERsBQ768qhyOA
4G5iCTynjorCO+xdEO5G4fFWPNcHBZvIJei5zKMLgaPy8w5jslSpqpMyK+Y/NJERk6yDKnc+0+tn
4oVBzuDYVgX+qgUerFgonocW+gkor9Wndk9C4PMNe3VeBHuEXvGxLhDf6y39Yloww6PJk2g+XaPM
N0zsY80HkJGcLAuusQK1NCe3dBrmwi44Hgdq2XI7aKDnJ19NF7arzFN/QRyS5+F7t3Ejh8hcdweu
Nbq+IK9DlAakE2BzJg8tA5eSCG7OHmEdlVRwZPpNKN7fO0YnEvXhH1LOjqrNqMhC0MV8BsnZ//hq
uhDyprFGNwYnJHrBB/Fwy1xOGvvwfoPar8HjohE0lM1+aiPH7/3XFfM2IaSbcqo3JwGPKxPKe6o5
IMTd4SeE/3bWED1o10c+6968zP3R/zAWjrnz+il1FG9yK7NK9joRULc1ts6zIe9SGds8SSNBiSm3
EnYel/z+5diwgni0K2Nl5clhcr7zJ0yy0MzBVx1kUFaXAiTrG0yjpNxU7E+uknWFNmF+L7rpOhIa
/5sW40qXIf4xC8m2sYhq6QArUqHkUldvDgyhYH9MQdY8zV+hcsvUQzkIoqTyXaooycdNLcI/PxGr
z4XQE56EgIDiuMI+AWgvj8eE65kB3H0taXOq9DXqNpCFgkcFgtARwVDvTluWtodm08Fp0gJ3+9PR
G+Pxi1yhoUYDnPfXMtQMcAAaHTwgB1WT4Pt4Vo49Feo/fjMxfK546mhsEQ3ZPgSQeBUi6ZNywY2D
hCdjtx8CaoyfwbXtV7Qrb7uYvZl3FmdKHQzd7Fxhavqzfvi3ZiR09N/qguZXWaeXdh/AsZOLhb3f
G9YD/19S5CKeH3zkbBCMtr9mzSxrKr1RjbjeJjaXsGk8gy/HSHPCtXXFbkOrwrni8ANMClItUkjv
XeQYvs8c0rsQr9crmJqHjxOWf29TojAFUngsWo8bkm90d5SXKxm1xabpHoemjo3rFYOv1pXdnVWG
8R2xk2O9aiUFjucq+G34MndE21MOI5baxX8rOkBFPHrDgA1KygzUQBqv92WaHJco8gRXHPsHuIpl
KuQeXKRqeNy+adke83CDnlp8XP1qUbFfAk79UYyLih1jIwLgsrfxys4ksAS6q1ysis1Fzb8NgMFL
kLRz+gttY+MpGWwPE3mmt3neWYlHmcOBAYfCxSFTLRis5gR91dUl29Bo3b3XzedwB8H8ZB0LN/Ar
/rHNJ6V+YVjKX4rTaUMggpx3H0AhbwzB/mWcMdd91MC1s95UCbvNdqVBsYilP8PzBhx4rFl0EqEJ
5KFXvQZHeC3Bh4PF1lk/S0QOZjlj/Z68S411jLVdvkfAxCdoNx0fXd2V9zIA8qThqpbp0NqD78f4
6h4WBzF3c6sVkjY/09kGz3s8/IwHjQr52qYcjNtEUkKn7ZnDVX+zkx4Uy7tdPH2v/kSYIu2Z+REu
Usy1bhoUYiYA+TtsksE12avRYnmlGDaTwdMsjcTHCvadCIxwGXOJF680j9aJyY+19CnMVv6yP5If
mx8BlSycFqH7sec77KrJ7qzf1NAnb3b6tQ19NpXmFtfRrjdWzOhvUEsU3EY/R9LBVqUIqmeuyg5s
HMKISo6HjNi3HgPt2sfN4CVc15HfVc17vQetfenS7x17VsChRnN9lvoxjYxHa3CXqYp1oJMq0SMk
X9gqjgbiQ/ciz50XDdb2MYYmsEjS2g85RaItzhqAWZi7qpbH1L75spACC/diXxB01lQTtuFoKQjh
eE0C8NM6sqrsL1VNVjdUp7AwkYRSjdiEfX/zFvc/TQUQFSkpj5nIWttjpmQiO8XwDxAAo//Fn2Ra
ZrSUQ1OJH8uqvFCVelBpGjimFNOWMQ8nMjQPLC0SkOSgP0kuDytT0lTtlp+gh2MBNPHRA1WjjnxG
82iwoJNf+pva+yUKE4cMd6EUijbDnDmxU1yaXdapdfVh6DDY4ypsPazlN1du3HCyYwPwVgkmXS+w
aq77N9Ay99/aa5KLsx8j5ZtgYTb7i7XPmIMI7CEfYZi8TbdMYPLvqUuTesQfbCtcJ+yM5M7ZjLOq
eWEQGCYeSWr2vKtG/XrRy4cLziCJ6q9d1P0PcGxLV+cooaS8bzDT8nNKF/cRZwZbE7gYSrHI7Zbm
R5fNxpGKMxUNEKwfUk8zwXtENCMw2RSB+/x2RcKX9myRiuuJpzda+uDRtev+sCij6N7iU+0pLeuA
EHXMaXb2MZzUPB2S1tnQkuE2ztSmRR6BmnB7o7ui6tS1Cx/KjlG5VaOARGPucf4BfT9+ncA0bhzW
xA/1vnFdtOp+GWOby61GNWOFCTZp4LEAKfJyaA2qao+zySvkBATnuxdh92bz7C87r2ps2ucu53KH
IFMzzHGRl2f+cmF4i2P9AV0BMI5JLi4HWQ1GvY+iO2EDhNhlEtNvrAurWDErEPObJ/lBDJZCJ/QE
OKpKLiwPRVFg/u0kFmXAfbioZye8/3YxD6AH5EEN2jYKK5ZwsRmFMXhTb7J/lBeQQrJE3h608lWw
IDrdWNA1m9KSwBpVs5UF1UH5k/OfTD+4azVUeUsCH6wzFBrQ82Yr0iz4TqrqYX8OPNJTXdgZ4jou
GSQIWe2qrfg6QbKOciJVrHxUwqQAID5UBnq9UVb5wlrtB9MNYBJiCXDGxYSvPy1+04R7/lQGJdHv
uJo6W9uILrlHBqD3zVlaHGWhgMKEKVSZJ9wrRJlrsVMZ0Gw6Ok1aSkdvWRw52qYytVk+FPRsF0YB
KhP/MF/K/oEJ+c8LKUdZAvsngNujvRpD6JlF+4kj8Al8AKv00mYN/NjXS211zAArpWBjQFH0zmNG
eox4P8XRHwWgQsXbDt3B2HW6N6Q0I5FYQv0XCQnWKmw2hqfO6lY5yz9vjWaV5x1N/hxnYrYYrEbs
phUbEKP9039Eo5v/nR6JROOGozQwDf0iYqRMMkreMJ/RNJlAECQytpysLzuZDMBgB+fvv8Q0MUX2
4W2WjJp9fylfrI/MSaUYn9jZPkI9xoOsH+t4vE5rs/bwHlmpSehAnVcl0GfScdCfpR44agQM9TEM
c9mIchWbz+UJgCElL7jrjd+tYpsm69oeHNUQAuXZy6PIvg17/v1Zkk0f4tp/itNVIMdoQVUcjVYj
FuK1FpDLvkSlRuZySrhPzlP6dy1NYtWgXOs1plp9l9c98xDgdErfKzxY+2tRjP7WpA0oPKj2dSJ4
KbLYjlg6LjYOfXFkkUuUnWRe1VcM9AYIwNkZFR1IQV/6K0a3VeaIOWAAs94HnHDiCMC7TlIyW9DH
/tksob0vPSNQdjDkBRdsBmy+ngG6vtvPQCYQHjepiGIkC9kk0u787+YWFVwHzG5/pJZTrHYCpVpI
wrAJjsHmFdEVU0w0kULy4FM7jqfohnAjdKyC0BNjgZj3a5XfAFk2AJT9JuIosMtOg2fohCYfNAc1
o1X1zeMtWdsi8QxuaOaY3Ek6+09qm0441q8/4lJK0Fm25JE+qXe0gZtQ7u5CpGJIeUDUY2bFv/Zb
S0NoIAtPR7q9PMl6DMHr2gLxrZ64JQ6mAs9i7LYJhQ+D5+fvDNOdHmEFeGcOZSbiUxX6kcKEsQv6
LgEiAgKKqYwB9RlgbTVc4/jrHOlnhkuiihPlnEf39Qof5QJ69sOcHF4cI2gE+9TwTLH2uwE7w4CM
zX7OqCj1vWbWxiRtPWgKPR1GIJrUpfMNGS5jrvTN9BspyiJz9bLdSW2hXMirJLQ68wSeQGjPjLec
Xb1ApNKZMRq3FopfkgDKTVvIqRinQYHTwPJaBx7KtEFD59h+1V4KpTe+9Gh+1eT0L/GuKcouLs1F
SFRkuRXzPL5J7plEGz+XlK6JNf6jDPYZpuY8RqUpW0EE5jTgad2iIHIPjoj/XvtEMHaBjSfY23BV
IAwvt600KVC22yVwmHcjqF2JpB491wtLO0TKns4tXSge1fGBcXZb2+Enzyvy99M4HGCGxN9ahgCK
kHGIMPtwREfp2c10V9IgL8ILm+Wmf7YYutxYEqlTMIsTm4HROiAq3N4lFCN9NwCBWucI6i3K2Wns
XRvBerrpZI8vnEsRKJvw0u3PO67r/zp8/WA2bP/wJNMSCClR0/1QEooCASJXHS69mIngYcv0eeao
buZCkicbSkm1+ZBCbk2KtsjdyI67KZcOXVvegYihqiPTswHM2p+BNKsOubUDu1k6zfdNCZEaEdYo
e0rSt9R0R+N30e2aCX24b7sH0yU/gxXSgRtuCStbSKXu0r/UpRB/foPu/+aLwEGet28iIvlpFUwO
c7zCxddSu9wb8noMUarePhxESzHSw/XpzDu9ji4BqPO8JXDm4HEnYr+bfIyUW6Gtt7c0q+XKX55H
CIRCC+PJdiERTdNZQHXOgaRytiy8B1W/lB0Ibc6O0l8oTIYBF0EGkz2+9b43i1ndqPic6ipYZK5S
kVXAfnSRNgq7pK7w3+NnovbJOKNQVhGIryEimeCfBO/Mm/wMdpc+IBciPJYA0SUaSTfuUbVBwKFZ
JbThlrEFNQLw6aKoNJkphVfARnRhbcK7vDfSEi87stJ+MNW1ZBayZannivuUUY1GYAFHj+IJy1MI
YTHQ/GYbQP3I7766bL150mllyRu4JPwCwo0E+rk4XtRRIETs5dGoRzqNy9T7sne/VvL1/0c8frkA
C6f3IQBoIVlDLduX9Zu5f8XC60YUsVvZYbjT+y7vupQLVWluhyxUwljq3A25M510ug+++2mx+OqV
y64VFBOf/KuQh2shCZccX2irIkpwx9RQEqMZtYTizPJPi8x+WKs2H/BnIq775uUpqJH7QAAzypVW
jFMhj4vo/u0t5rcXbABJJvW1NkZNYdGCQnZLidNcPtp0YynNNyUvrXzsumCxNONsi8NyFL5z4KGW
tll/q8ycx5L1xgb4LLkvqjTHLjDN1vK5wIwCNnCBWa2mYLg5w7DiPpXJpYqN5+m2mShld4Zq3k0t
Fu/sT5q2P6Td16EAKQP+LFnldTK17cqjl+sZhk4g1QfRV77CFITcSz6GlibkGPIAN5Zr4ww7Ol29
q0Oo1q6xI++ND5KJyBWsuVPVmE1BqSj+bap3yz1xha8hjF0uBGk1yamcFq5EkQ/rA0jvzwOZOgsj
7na1j0D9Yr6MX9kz46QjRZwdPakUG6QThXB8H7ENvb4zXpYuIPRvgD5eBKPTJbdBXU8ZMamcpxZc
Yeusvfkz1Rfi1RT+VF+o3KGJlQM4b8cOsaNXNReAmTPpQcH9xWMniS2IhEQWGkVbBX8S3TyYoGf1
/GUZTRgjESVnwlBxUt1jZxiY/LnFxxaNxCq9I8IHqgfH0vKpmT7Uk78ItPPNJdkfyIfBcdoOIGLo
76VnN7E1weyBzu3iC0QDRDL1asPL+HKfGqkW6IvdyV8LaPeoOytxFFqrMJ66hi8R/SeSN3cAuiAQ
WKu667fergTx8WFcfbToxJ9x8gJZlHIbubOga/IDQ1jp9L4GA7BxsYSkUe7rS68sXoLWDAYXyNgt
up4yn0+0jjIfl938oSxj9Kiz3IfaCxWAuvr5ZZ+j0szl9qXSUzTvdSantnXf2xQTnVSQscGIVxzg
cVjbZeq3kkJ8uRbe+wh6VDykVxAFNmM0wzr3aayFIe5Tk1wXA/FYIcZJ3F6PrHlX62raLWLmKnPo
nQjdsP6lTj2sDq27rlYiQizFeu0QWKBQU24U0CF+PciE5QkiwsWJp7fu0sNmYTSBdanfuJo3RgIO
LmX1SP0NvIZT26kv6ynnUYX996Lc3rKf0/OtK+SwTU9m2yu0CEhN4vANyjYW5g86I8XGLdB+aSHb
CUVkY5g1o9/N/snCNhqoFE9ZhkNO64m5AK3hQUVWc6LewPhegHLZzLjCisySMHf6e7AxUbK5AoW9
u8DgSb8D0TG6OD30658Butm3nX1nk1ZS6R2n55jvvF7bpyXMtFdPUVmq6DYokF2EHaXGQvcOEWr0
gbvGBCr2RM35Vv1GLyrevl9YEG8A1n7kQ5qLqmKFjdBbMM1pxFhvmlitQVEAxbs36BF9zFWuQ7yx
u3RzHVmnhdKcA88WtB7tGtjiYYIgO+4IxRftuzg1u/NwgGmWG2QIQLBgZPDIThs038VHBPrJaETf
xNFs8oMGfFmS++rl32d6//dH4yZ9a+mpFJUGpFi3vbFUbV6je98jYC9fnWGSdbGeUk/2gAuWyWUv
PRlIUPRPVqzZHH1G13m1e9yKWkj+SbzNeWAmqaKZ5xNEpHu++pnmOImtYX9OP4gyddsR+KtHxaVn
9yQqkNRf+5rtoAPW6pWazQAYAcHbMPvU/E5p8RHODgelRKkj6hyf1n/dNG4vaW7FTU8nC0WkuUDg
cJPWAtSIjWVBwLR+vlGEO2LrZNwXdX9V1IwhxMaAkVyyRBJyx3pO9xBLgip2wq8u4oyZhZatjkgZ
dBVEVVSjsgTIwmy1X94Bq1rCaQwx3EqfhdEGSf6VOHxVgQTk5XySnaqNPjivL8k4jKmdcdUwL56x
CWNeg3Yt1Z0GxIYNex1kGnVI43cfPS822rFw+ZOoBz8ch0Y/5rOzHlr+NmAzl5/SW5rUZMNUDzVz
synnNnsQHF2ZwlajWj7J+nncytLIolhp7MDYu6LGVRxj1yj/ot53MHimVA7u9MVBWpoEhdWrJP31
n1Xi6IN+TZXh9qu67439uFleQwwULfdguJD+Jrl9NY0q9QGc6pSjFoKVrX7aYQWN3d1bo+MK/f91
W0HgAvV3wUrB6oCNvDbTnNaDU6oEd318ri0lwbVu4Byt+WR0YaOzBJrBINeBv3hz/Jv5rsbsOOEJ
M9db1nduDBGfNUaJH98OwaVlDzFrATkFvKiuuxsSZ470dgzHBgIvSQiHBtk7HalMZ9IurpgLfZRg
HLNH8LxmWX/OY9P6WlTIstmw50UEY3dzVDsEBwQxPZXYfLeS6sKff8vHpENaW+NGKL4a4kF+IWH1
qksqaaM2kFLfbU2oe9fHBJmVdl7+X0VZ1MPO7Mx50Pog+lgV3ngNYpVtvBqkKxBSxzrFCDGIxMzE
V48O9qWqBwAGEz4REC8TvFCkeKfCPBZGO/XeDdRIYK9VNZuRDD3gqHus+5wBzRJ6f0Wsc/RBvg9Y
D/RWqnTC3t3ISZzxi++8CxfgOFMnu6+gnrhZnsvbzbEPDkXYX7+NtTZHWNx1uelPzimFeqfLCRpU
OrypQYlKaq9PeGVbCxE6xQobQ1d7s2T4h+1oQDzUq6e3gloxbklA0fiPKg27U2VLfbYzDbYS74Nu
54fGafcG5LnSR7jFuUxlNrEd9ct7lFmeXG1DL+eySU4x1GTPckU9al6XBc/e6z+2+xTzno/EtEGy
XaJx9duXCOcQYBe8yScvJ8BGxDQm2tJkQUommBuJxVQU0+XWAPUbQ9bTqmZad2yRaOfEryKHIYGc
UVBfLZyIIBvnRBmWV0upMqNh+UNoZ9drDEulF8WAiNgRPH6i+UBEOhv5cV+o5e1iswDPEC59NSir
mqaHNNAYmAgTp2d8JzA0nYdTOp0xPUjK9NwpRVb6AkbTl/ci9yAro+fh122iFm6+TM/LjF08ekrd
kt8Pd8pwjCxoFzu5JCUXtHSPZDmvaYKrzNis0/k1wQ875LEWBS588ppRlN+mu+kp9ChsCf7dYvdL
N69wYZcgfwgf6QHYIXBfm8qKdgXPaR9M2Yl9kPU95UrkPEppELv0443Q9FeiD40Otyw3MLjqETVt
J1xrb/1iVhYDiWjrcN/0NZakw0brwRAizv/WevpdHTT5+wHzAHrH7lNWKVGMCn9aEYZau9kuxL8m
i1vvvYhSTOaxh7yMDCKe5gqLkQLAqsu8EZePZEJ3YgJ5RDpGbQip9N2ur/A4UbmaXK8fT16y8sgM
S5PvpkCFw6p5dtnNhagaj0UvFdPN/nosOCu4dpS1YCZ1IUUb0rvjEJghZ3d08EIp69EIqSPYaCez
hQqboVjedSKB1bSstg5GN0Jk8/2OcX0d+gP1onV0/GvDeLKEAfvdPGlo0h8PM/ZVHLsFRziCXckF
ZV/q85oRiSHtD3Er9PZyG59REOdRReckDk/iRUHt8oOO0jNBr7r7CTIaqd/gqx32nUG04gqyx+rF
d1ivwJfTWegqdlq0ewZ6nRJp9nG+CK0Kl7IDh6C8bTnqpuBA37wAn3I3K+sZtvllNYkmQXm6Wtgl
gMjgSE+e8o0xtl9mz2wyyPEaUD7xr7reTDqBZF097tl1FBtAS66SFGGgqaSoUobGYd5QaUnD5FTL
5N186h7TaeVt2s/dfqfE7ub2f+bIU8ZcXkhexZ6HA6UMwUHf58NJbUrq0Z97yF/L1tAE8e47nkZy
rp9RS84j8/tkrG/Cs6WyrwPzfdlUe9n5f/w2Hb2OD+PVx4ClzWISmYdtlJ2yuAk/4HLIUIjL1oHZ
S8tH7vdw4xzLdBteOj0MVLGSNcStt+ByqqwvDo2Qxn3FzoNipKVmpGLDCujelDC2gVd/Sd9i5VU8
Q0HnUi0/eo5dGLxOKEw0iEGFs3espXFaQogU9hwvZVtx8UTuEiOqjOUJbuP4BPb/coTZwwsb0OxP
wqOfsiHIFotIqQEhPDZ2SUXjHuCyfOCOn3ss97T7+tlNKaPFeO5kpY1bJWB+q6cS1aQzuc0X1n79
s51pAQEgw9vKSZCRoHDJ9Fal+/D63THBuo6yOUG1GMYaExN/FZRaqXSyvus+UqA0KcdYcMG8j9fH
V7PsWKUzqpv2JPxjMrUpZAF484CVR/XdlJPR4LsYWcl6GtvKS3PK740Q7IJMfI5KhoNjezuVClOf
JqBiGOlN89AmvJ2fbYn8d7OrgeBr0GKK+sh17vQNFgKHW1F2E7GXW+sCPrUvcr6Bv1LVjWApwwnS
/IK+HqaY9ll/4TF7YpNancpKcVMaSLEp0d1YsEp9r4Ibdsb3ta4sIMivRgaE2SOw0UhJ7G4NnTka
63Et0Sh+sJa5A+rUwxh8/2BJ5J3LajICo5jJ8pw02vtikMEbihBy6aJljGqpkadUJTIzS4jix7Xm
g7WR1fgKfOLcQ3w6s7dFhirPNPkhjCa4N+X6YuyvGS9va4nJf5jlx+PFCB9TS0spxnCrtmD6uB8q
kjUqyQVBSgw4H7Amr35p9uydbVHeHwQL7OlcWI88ysJ7BCw3BSJq9/+HasqpYU2B8+G4mcgj2NsF
bVBhfI3bEeUa05EIe5PwDxuhS7SgElrDgLIZViSLhXQnOmf57IKOSPv2jB1bHGoLNWut4OBN3AyK
eMlhtQImEKd340dsaGwQYRIbLxw1kNAEs0HTre4H/9QqTT6T6DyIg01XfnPOjb7NWeIyFLn8Zlew
BrM3JLd4J2KGIqnOMrYs8rGdHz5oe+8MIyhfGIl1r3TDygl/KY1uK1/8ZdrJ0h6aS9dQe9RfDT7H
y6jN2B8+GbqMuykgZrOQv9/1uu3ZyAVSp6+Wb81bjYBt5+A6yyg8Z37FbHfNoUZ6PBc9SQImJiR9
kP+Xlh50NEf/gzLjm5le3RAGBMbXbMkkvIUlnbTImXsx1Uxd12yus4uOBIAvnU5oynAADUwQiXqY
2avgQnqa7j5URpxHlVB3rNYCkTLySq1SgaqvIhyFIvJzU/TsJJFgzPVPrxC71kyb7vEnQAOsZ/To
50+gsaEmjmUO6oE1RQyojn0n/nuJRUzbQi5BnUW5MdmuASjI+pLDIo4SW6dshQxcIuLPyFocAU2j
Segfipmcv+/VZPUZMIa0ImS8If7IVoprcVy7FENQHqUEdqTUaa9QNjB/lI6b/icgg/ckXr1G9kke
rx+fKGNWhJa870UKaaSyHtQsMfAAQBdCa98T/aTqeImAdDwnYTU/B77ull8Hz5aWsmZsFqX/rPSH
xInsxjvBFyStH2eqfAiPDaHHN+LrKcmoZVVwFCNfBa0bd4WWdqDeUKzco/4DqNm46+NseRvLYMmN
aNsk05fmSh4GpgvcHC/NXV3iUOjeraG1DX6zYq8AI7dI7nZintHc5rm5n7DMpxIf5yCwEK0+/quu
gm55zpO89+qA+sHzFnAP/iObe0/JibsRZxHfBZGprNeZuFnX8SCehddYsynyOPG50MFZm6vfduBj
EvLn5xoaBcwl8MNXd8okKGOudjIuyG7YXTE2vlOFjm3C9QG5KRRz8oFZAkRRl9iqS6ekCgcVrXAq
dx8S7OB6a7J7eV3ziazXUSORpmUgRdTubXHfYGmYkt5U5AgzOzbpQ+sD071GCUW9sIsssPjfgpxh
LN/krJ8pf1jQjBC2NqcatgLT3RpkFU1ged5fcSpMSKh2d2QW+zPoLg0GxLM96m6r+pjgURYljD7i
fhc0FoZpJwIx111nU//gF0tjeFn+22TY52m+WWzcrG4mnuWtK6jZxqCRgaFLyHXBlcB7/1NiLvJA
sMV+jMemr3f1jtG5LAKdMV74s0r7m87rFlwk1lBhCrjDm4G9NJOoR89Y+IaL3gcsZxsrS2xEQ1F0
Lcpyb1+Kew5nJkIwo1I7nOvk1Z1a8hb5JJl14hHA5XvdmelLFaht8ckMFkEV/nK+ujMnATplPI5g
r88J5ST9B/epsY+o9worWhQMH7bwlR0gLQ3UH9RaqmSSV0t6xA9zzw7YB6MHopHmY6BwM5YXBt6U
tW7k836n0ZbRdCiYVJBQojGx6e9zf5DcgQtR03xFKV2C5T2vBYbBzK7oy0HTnpVssc090DxdN/jd
v/4swA5405dxnycVkfFW0Oc4ayZs9o7u8q3ytpDSKoN78dFXW73RnTAF9GjEMK4/M64GJ2cfNxJq
sRlCRFRLetkSp3vgm+7OVw5saQQRR+IYFxLUBJNJWfnzWkak1lILk1BgT0X+zDsljLANRjhrTBn7
Fbv0PuFb5Cqkv/iDsdKtz2aQufh8xfT5R8hxiyHZ6fKj+ULSczHgDL4AM0muCOR6YZBVM5XzTIzL
M4EpBUmMYQQIMkmDlAbyaijZLm0Y3i5QkH0lqEbyuHlrp8k9ZBLrTj6i5GVbtixzt8q4o9ery477
55Jo1RTDGh3wGg8p99sjjh+SHYh2u10l3g8hicCrcx1dUZvmrR9piLGyxzokN2fMzn+gUXO/28FV
1GI9Q4G/INxR5KTb5LmtBSu1jDVcIOVd4DoTfd+fJlICaBjnvy8TIzO4fEubARXbSWyTdbhhDQcn
R/4jMuCRjH+ih9/USz+AR8L8NeQ2+EL2zT6URXQaong/UW+MYJGRmQq37bpa1+Yl3ZKTLtgNZ2V8
xJdUX18EZcjZyuPwri2qDDhab2a/9XFQL1VrSA46urjx9lAzi8U71t4EsuRLZ+6L+arfha6a0xtp
mkjuJJUO0rDEEuGI529UP+E0ArnAeUIVhI5Bs4Hid4F3JbJVx2xMojXFz+MtEdybrFrMqgokWBkh
E8xkSpoD0PlPK4kLqVHeoxkaWchZ1TaRgM5yHeTRJWFO0SOTun7BUOf8tG9mpKf2IBLsUa0yx7Z3
mn7LWpfXzCIVDvPXZoCLMEsfpYtOKXAs63CqJb0f18pWUVKtCcoNezXu65DX5O4GFp7I64hkMGpI
b6Ow0qt/TATRIl3fjHdat21Sno50xQveMjFkVuYDlzAKlBweUuez40f8IRmpgKOnLysPmYMsEUnc
i/ufjjIQJz7GJ4Uy3dgDi32aVxeco8NbbU2x+ErOaZynyUgsk4iOFXBTbu9hGUP/SMRFt2fDZJEa
sQIXkGd6IArubxZlw8n9ptz4W5LJ3PCok/Lnd0YcRL+J7f6Fgq0rlCfHfnEn6NI5khJQVueBuF8e
iY2fRKm1bGR08P4x9VUVyQvZUF2deQ2vv1TWRxuLstrlBHNUoqsiEULxScEe1sgkB6g+5fyjBy1Y
t9kfuWSKjnxbS+GIw3T+8crr5v+cvCBlvxBw5i3f5lMhRCsC27sWCPlDXecPcFkbLQrQuNuEtRV9
FDLT6LZOvWYrbOdXT66FyiTF0KLKwcdBVmdMRnMArIBBRvZCfGTTWstWq8m5W1h/Kvqp6QsVy5rK
J3FAMQ99Y9xEqmD1hP+JRwCWE0pzdm1Jm7JGnP2vF7rf3vdNt6l/J/NxTE0OH8oa88Dbb1xKi/qj
SsbtfxA+zTwQ+9HJwh+u6IzUHOnNSQbcwv/dACnCoIgdmmJWy6TRDvpd/2q3xu2dp/ZMCzB9S965
4J9zJgO3mFysIVhVGKuJ7GbjwVcWdzRTEI+C8Q97otSl6N2XiWhXemUkgZir6L2eZjTHCJF8y4MV
++7lu70DNIRv6HsBt2vRqcbSd5Ymf7/4SclzLZKPCRIG+4qcSrsoMphnajfqvwNVJUPUk7YYj+K4
FtNdj8qYIdIECSZM2rlpZaHnBUf7ig8jLYgAa7+DwqLpHw++in2DNvvFODT7a7dIDbg25jrC2sFQ
ySZozAx88AWQOlMm0UU7riliToZJiu2md1OeamQo/96KxnuuJEVlWh9qXfnnz0/X3j7v/De8885O
RwUw8kEFoVeDaNjnXfz4lYSt56hqyvIE4y2y7vQLUPD+A4k+UjTnEFeVNA3AhrpEImUbsj8YJHW7
scQRrkP13Pc9gpbsfDoVR8tC19BgDwrkuvN+cDrCwwNMfxNPq7u0n7fp92b/rG4bjiQX9bxqUeW1
djbtt8/223j0XaybCv1NP9BY5v4gdkkuQcIUPVhHjqWOdYOK8rjM2OZt8hLx17Qn+6aDCPdTFDru
D+3M7f+5+yEacUVo1Bx82Wb22Toh27+1FCd5lwwL6FewBv1wCV5OhuZa7Xpl3ZshF77XXWr4DFQS
qDjyeNeTVS5eQgBCQNQz3vgzmVEtgtbKf6hBDYzACvFqPixWp/sMdAd5oHv4uD1l9dny3GHrtTkx
TLDx6UeFC8h7Lzit8U9x1ZDcQapqdxrxUAshPfzK+d7XuS61z+dfABV3UFKoRq30ktJfqKZVplMQ
S+w9/hBcCXyKOAY7a/ASCct47vET3MCudkic4pgxOggugzeM6dPgA+8F/VXkO3TY0RXujmR6vobJ
TLvjS86ol90Bc3CSEZrOAM8w2VUP3w6/mh3MOFFt4XDhRuU5uj6jDiELClKPbJPie+J2H0gekazg
cVk4Rivz4tY7R4GViI64PlvFe/VpgeEginC3oAxWcxRU93NIgSCJQAEnerWV7dRelJsblac3DddJ
oUgB4r+ceWQ9dbFS+7xrINeEU0AyGbHUqzp88R7Bo3lGXf8O7asSes+pd8U5sGOQaFhULl+bLGW8
mqOk1G8UO2VcXvH0bjpGKDiqe8VURt7HL681w2CAE+GWQi/kLRn/2fHhoCrhpDYUKmw194St6PK8
+LQghKBkMvjocsfGdaq87DX4toKSNynsbaIUvxzHpsY3WrBH5IviZbHJvZOTPq9srCrDUI3d5Cmh
nsibOAFTn86GFhS+4cS3H1PGZJ681njgszGpfFVsUyeRtYFle97OI5CluQPOqAMkXBDb1TTWycl1
eWRdbJ32l1z9LMBAem9U1hoCq5CyJ6sGKzdXbySM/U/RRmnVhMoCtSRZb8mdpvPyTEWZsBEvfafr
/gM9bx/2HRtLfO6l6YuY+a3k5xkujxlQblc0NA6dSBvWiq4TA3Xy3xdCIC42eWjDbAWsO1jLr2m1
FeAtlwXn361/25qORXLosLh4rvT0U3lQFoGsrj7mhgDPxRCWNXmQohoZVR0ZpPkEcRflMqIkSTdT
ycuzo5i9IfCi3lMW0RPF/ObsIqPl0n1HnVwOL/u7yq3p3ebTLEZms2dgDgdlkuHXTZGpNtQemGO4
WHWId6GD+p6QfiEY+qcTQQkzLbKda6ZS1PsTHd2TvAdHsPw3uKZD3P8EYkF9YFyurLc6fimqXDIP
WKgU16/ruxhCr3mHqBsNnZzVy95Nl5QYMpsWCIGY7FTWqVYRjUlqYXxs8v4vRakVK4YBcu1T5Fta
KLdG7ufZcLx41DVcvYekXF9jjsqQsBDynFwabEaWSxlDQRIBoaL9LZ8SaiCXaFYvv7eKot5oFQVz
IxhHJ5oj1MzhsfQ6/MEVxsOjHgBgAS4MBZpJL6Kqc4VReGmqXpKPFLihO20EY2dihnxak9Vg2/bu
9ARet5oqvpOiRszHo+dhXTuJSApJ5Fz9nRjEBvXl3cuLfBV2TzO4LVInG5h+EIv86YInao8F8Nm9
EF8SIeXZn8Nal3m8C3dOOoNRxvkUHUqONDujeuSDpwcwpIlhMMHCia+7Lu25Lw2J01Gdg0sBNbbZ
+mh2meF0CQJ+cMmDFqcHVj+FMBsT62kWNDwVSX9xZl+s/6U4zw+F4iwpjEsuvEDqzVyj/MMpYh+j
HJOopKk3ZTnUfI0kqRSKqq/wZQmHtJe97/JkQFR78F6c/BxhwssWNhxnb96o7uwBPGv9c8hHojW2
8NeV9gl349fJt9wrhPtBtQ0USKK1GXxGAoP65k6VdXdi/IJrlZlILj4o8sPLw/HTD50AsYDJ2Zkh
etRsGYVBD6GBFMHXEqh+46FXlYdoH8bS//3ZBlbvceycObCcl5UdT9yim0L93ek6fML8W9MCNwlT
t12SuBoyR05BGtKrtHTano2GtuLk7VbuvyDgm9aOp/FCnV5ydzn8g+usW56F4bMzxvXcqrho/Q7F
xnVDcFvbGN7ZN0UjECXztzNYdw9Zj9gMc3BA+XX9q4jYKVdsY2996m3TxyZT/MPuA9wmmz/oP7BU
SpjOwMcbQV93x1PZA2EG3QQA5/rW3Nmc01oLnKacyvRsr90VsqbpAzSO57cSWBRf2uOi1Nl00IwU
9rNtqjAsAesgrDn17khiyme3WnIyd43xP8oXmKTaC3kdS+mDD5/X0stwKRSvd2fzSgwg2y2PN43x
+ujOHpsTZT6ZnNkRB8mdoxHNMaoLN0BOh/NhpQm/pagX6J9Nt8j0/5EBvnjgYhXpY8x9ND+2FnKG
gY5rjejVZulfGGBEMUjOK4J+Z3l8r1cMAJ/eHVPWJpQ0MuXUreD6ITFhpT4kui/DvfpgCbZf0Tyd
M1of+QtgqyiVNfpx1smTg88DxD/TdC8TgR7ET064+JvuwEr04hmfBUQS50ZvcQcXwHyiSUt2eMxL
dS5BSZI9/Rmqar5LqR6aV3Ym7tT0CvZ/UT2L8ooVwVBVrwyxnH/iGBgqRyd2+GMEbzAAQqzosS7b
Uk05D9XXTV1VJYhzz2CGuqB37qP193PLo7xEsEp8FGqNIvyxZV9QtjrBEuwzKaFHjdIQErKM/zDW
VIdiZPG1RwVuT/HZ8Wv6vpXheEa2pUzM7HAvEtTo/Nm+c2rk32IotfO7CcVed3RKLMdh1paN0Wlr
5diXGt0XtNOm1wAsWoaIULMKHDwq9SRaSkeRQypt+f6gBE2gGt174WiL/dSZ5X10WJ+UYHyf0fW1
1I7gGYLpwTVDW/6VEhchThp4ktTxm6IlDAt9B26cYSVsJI1Ym4HNHXlDz2X6ydZbnEtajaHLdXJt
XaDextvIjGINDLBMkCU8eufzn2RgD4neLIOAP7SyFeOhqVN9EDqEhq9o0MC+Z799Pz7dExrrbssx
8iO14eJS533gdvfi3p0fEtZZGEw5pyMabxFImfwlcXKbnE7zwB5YQNmQI0svtY7fR8o9MEmGwJ2B
tqZ1Yqsz056Y3AWJkdgxNBRbkWCbfToi/Vw+nv3yoRIGlB6e/CK38Z5xr5TSPWbVgJzQcl5xDdEA
hPXkvV6FcaJZfaaT/+Pl+OOl5ihhq+2ZX9NlB2xn61FVjoFxOSE6qBBd93HTO3OiaHLhMo6yapU4
iyF3l3n9v0yM/csshqYaeZMbbzaF1UzrzlKNANosWNHrcHdrsZMV9JQAJgT9KN73vhemZDv/Jlr1
BEAiHrTncym7Q86zaJSNq1BLL3QuriD0qMk/aVpeSLTUpV/JcZv8U3DvNTGntXww1qMIi9Z/FBnc
Cc/WGuo4AlTueGaZLV75TWucnvHozLDmlilupSziutVptKRDxeCF+bCcKSwbNsez6zN4hTyViZji
hL9EBrdr9iCjn9Ra4yjJQif5j06nO2MlVTa++rGxqAf1oF8B780gchulhAHAPf92o02kJK9Pzo9H
MWxKAtz0rr1sP9Db18Hu4k1rcUVv07chBJ1E8Ri/94WY+ZSQ/KHfC1sNgN+7+3UY+OB/2Po70zOw
V/qdpQ+OsBp5lRG54u8CZJs5kvl7T88lsxNUgyeUx7h35Nvs0k56bJtHpLrp8uQZ+nRbndXtb0kx
pGIL7b5JJhKXGHW4eysT2N75xAwx5TNZm13q9UbuJ2NHs09YueqB5t3wptwO1tTcZpbL73addPRY
XSN3XJPirFCjA9rJZlk1q3B1iLXVs1bDC+JF2rNevCwQyIw0mCPsG6jjzS5IKy5gQdyjjEYd8eKg
lo7S35hd9bYIy37AH3OkUYQIDV1JMSxIDpjHaCpwVHGiz7KMedqzIc4cHPsulMoUZg/MEvP2F6wT
+yN5hO0yvifDO4p68yw/EIuY6HdPdZulnlu5NRl9UeVVYncR5LrLXILAOEgwLMbyIAW+g7LqLRs/
5wtSE6Z/Pk3IvUkmwfFxVTWTs1oi/rRdxIUUqWHZNuWWeBFjPCZsuTKk+KzPrG3OC+X7GpoD92Qn
V1ljo2c3ycUdFwngxiu95MJD9FTzzTbH+0J2c5id8ZJwG9imEb+QHMqqnzGZlMlqTLbIFv5blCF7
6HULHSE8e53D6nBl5q/jJ/rcJla5zbkI0JdxZVZ25hMBKW+9g3kQgXl+D/8QR3QK4Mw1R1HMbfL6
GnB/asn0tGSRCk5S7xLISS+whe/7jSQhiAiw6BTqP+mcegslvIeisxYzQmA2LjwUTCRMzEcGqAwi
iPQylBwLfZlSGKX/F0zjC98/Xa10fXIA+WySisEXgpgXpfrRbsFql0D4o5STa+ZXKIAYx+z5QqFo
iyH1qbOoF4FUaKEdCmC8t9r67r8KwblmsKlAPzXo5s7tvA1embtfnR7txiak5aqe8ezTJuBqlR6S
7+bVRtkwmzZp5gPeDARqeGpvV1Jde4pOdrH0HKQXbRmgMZ1Eb17C93cr60hx0KxDj0q5obFbqUiz
VXNUyv95RxxGxG2WKB6QmXK0z0wK2WcEGPQOvWROAqTENoF3hdq3shZfjCOjlQoPgFyVdwNL4ueV
EjftYBG29m6z+PzgCyju+RXYBNk1PAVzmbCC7b904GtOM3ZC399dRoMfd/Mm4uw4QCrvcqDExN+f
Nt2G7/trUtbtIL2FsoAq++hXJ0VeVuxjo+YZ7fP8pMgYybqPnR0dv0ROoF2xMtByVfsrF3J9EOjh
PChxFUp8txlLY7a4FXv1r8QfQ91aOijLODC4sLDZvA4oCceQohwN+B7A57QYYW36WRaW7a9C03qr
riut5t7rT8UjhBPRFNp/wn3+sun0NfSj4EIjKjle8dxotrMu9Zq5pfRJzv7DYZ0kWHg6s6bAxtDa
nEUQcLme/RJ+JMhle0t2DuRIOMqaOwGruHk3SfnzjTHsZ2g0AEBw2koqex/qjFRK94TeYYIA+rWd
8Hy0QmYYkiTs7YyU2LY5FblP5BJ5ABa5YfeK+6FvzZgjLELeZ9xZWOBnGTWsCFYqKdPT6maJckOU
VQM5HNme9ijUcv7d0rgVToTUykhrcg0wmkpcgXaOCM8XCKp+nM9lHGoR5ZN5c/zMVUWi2JGcwSvX
peO3prdJbKw6ZcOiKYXlQGZbnQDFdxWXImqidKL8wzs5nI+umvMO7X/3Whgd8rUrZcrF37ZQLaBv
m2/2oJibzF4+/50v6Bv+usy4osaNekWBvKmLMxDAarojc9MOMzR6zPR5y82ENRup9Ap5snK3cCwa
iRbzw3BW/S5xwIAZ/RbCwgmNh2oVAO+gZ+u2WoGKn3rENx9wMD1dDsrNdy+vVtZnfnjg8wlO2yTv
YOoJwi+IPuQnA1izKUPPY9+0g2Q6V7wxBPUYvXUZqSJYHkn+p1qK7dPeF8zjzuQOgXavN8Cvxh9Y
6eQoH9nqiiRPnqWjY+ZFfRKBrqGpnBjFZAusSZ5U6QpDRvTfIhbXcv6Aw27LC5DTU8zp1mVQWEwx
FO83Bztr60kPIoyxN/iS8FuJpwaIHFsszI7DBuddFuk0s/Z2Smj5Y5vrDBiAXdAe03MSB5FZdVpG
LOtngy1u3Ico5E4w756e20S/nVVFXb3kUitUlq+tLIXtWoi5eVj2R+0ouuj2UxduS4pympL5th0a
+sI1leBgiZaT+vzms/ntViZWIYGnZcXQI2u/eUIRDp6ka720VrFjQ+idyO71bz/UysSMjndu4pN7
yejOcyIG2gW9kQlynCMhm5TyG/v45aXqBcvAyLVffu7zD1WoZ92Bv38VWqJoJ0+8fkAXRerhdd8P
0+imhQxHADzzI94XxlRM1iJjgKHgMIGtT+uJV4ofcZriFi1AGAx27ic/dFlF2GmN8HAGfKh2iI0x
p8rV5B8QKTQ4mlM0nCBryUYbuNda2Lpmlr3JZ8f5G8NNfV2Fs8BXNlMoOtn1amJfa6uGqulYUoRj
wiWQluTFkGUnWkk0AQXrHYYX21LyYmj99BqOAde2GcthbWXqMfYqx24mFfMof+0MJtrtEL9laK2o
CBcGMT/g53krde2VVs25OXgQf8AxjaYsYzFA5Gw1U1xPjyPVdnlGmXDdc1bdkDjZv6nTl/ylC0+y
21lwxbDWIEDFFANgkb8U0k/FZm1Q7rlazCS7hThUI6Ojq0LJVRRI71OCqvkTIjxU4J7Mi6AI4Rk5
mnCnlYBW5le1YqNKODpbdt0UA4cYl0Q7CwlskyTdBlrjFNfRWDquoNqdJ1xNEcfY2s1bc2At8PJZ
JGm81JIida+8fjFYDEmK8MAcs/mF3QlqqkA0Qo04Ozi1QR2521KMZDN/NhSvCr5TBziy7QsjHwUp
vZRUTGUEOj8BPvNdkV8SJluWSlsUBi6wcXYJ9qHaOe1e8zgrFyI3XoK6wbAT63RsgTDscneDzcSN
4hPmnKai0hjnQqRQI27k8RAR1FeVIDx5Lvzz/fiGxTePMM4Bq85ug3DEGftxGJQydhiS7dYfQxkX
9sC1dsoCibMbTj6mxwEerVR0jt6lTN2jXxKqBoUdsB/5Q4ixaLE5GNpGERbMXNUZO1AR97liQ5St
KPfVTdUkUGcoQWP8+abpJV9EiiIoC9JmOYB9ABPh8XrJSErWTdKBzxx5vgXhbsWBd4Y3xT8GgHmx
en4Twj8scUDpICi2FDLZ0xCvVALZ3m9g3Y9/A3IMooIDE+fleZDYJdGSJ8Vb2ewgNQSmO/xRinT7
oYf87gYCl1I9bFxgNR1AHPe/tLjWMSJ6AsyEGLActB6thVJCUCpLX55izrWqSQwDs126WxQ4rMTy
8Qakw0/ZFUEjN0IhAkzoQ6EXFttu2mSZcAKSeoz8Dkli3XoeBg5BJCJ3OVCjz0cYqTpWQlzYVCAr
kBiAcH3faWIhJFY+UcqoDHjo8/+x2l73U5MQFlXUl3Q+T3GJ6nT1SVC3I/8lFUI5kX6GrnakSPm0
PqGArptKD89lF684LPV/KRBEpjG10zwXd9M7/b8KFfWEX10pCPfHE5bV6gf6w/bKdZgG+74/fG/2
fL9QsvojTOJFVOb3yPErLAcrazATaTRLDaWrfPShz04YYCAPRfj3wiVFINjGiLRUNgUcnQ2Zfcvi
Gt/oz0AiLJpqOpxu6BuQSq4ISmxJgTekD/Z17MZ3Fi+V1Cwbl1MpeVHUnm6P2+9FB9V5TmIG3SqU
Y7qFwkgFN+QgFytg+D784ZyQ7kYAEtBymrXsTyHV+CZt8NskKVbAlVTujsAVnloFW+EQT4NQssBr
/2YiykzavKN70dc9kruJrOECOzh8KPZVWOwe5xm5ywU5UxTACBoXKluyqD2LmN0jUBmPf9djebNl
obaz0cwZq4yregCbnwNLKioOpaGzhGABYiLp8eDSnLcktdZhpphAa4M3moA54hAobapnUEraEffo
4FL2qL9DyRdC3ultp/9zcIU/mZVfyV773j5n95sLm0AMxhw0Dr04BoBrG/Vtbs0OUWkW4CFzyc+/
iKSsh/V/gX2EPvGdfnqTs0u0HNzKC0yZlH1XQzU2HZKAffBxXmnfjMUqHwomNzKdGsP9e7FM0nLI
bQoHp5dDcLsYcbX5+CDfkMjVnJdDiDuL7s3VCdn4jXnxB1CAZeNgVCwh36yIicfyK3t1D0anA+rn
iMK2Jh2+j726WZ2070OK8kl9hPf700AXUzGCAEJS4gJbLRYp38DNXjTyhoYcb9Mhd9irIA+jHAyL
TxbX3INrgc4T+rHsovMBi1BfdWDCDsNDkOYmEbcrJVWiydZimmNLyiVG+n7kr+x0+XMvc6yIhR4D
CO1QKFdDrjuo+9tWl9eiLy4fAItbId+ikGws5ShIXdQExQzhg7uEpqH4audvEfQE2OqAK16xS0+D
yXbc64Ln57mktR3BgA830ZaCQfyHryBe28/UmzgyeQ2kZK32L00xZq/XVg/rI12zqK29HbK58F+V
v7M6DxMKL1hijVAY0keoBSvP2BqV2OAW6rs66LN+RliuXA0c36O7p6DMqWGup1m6+htrY/YqfGLS
evCuNoLwW2Q7A7zMAplzyqiOwbsuhlc+PjC23Mu/qbYZ52tXfZj7pv0qOKEreyg93mPdx999eEWq
sV7EKh8yQ7Dko+FY4VJQ5UcX2x5Y9iPmMnKiRCxDbg1Ju1ZO+Z0Y4jgFB9cgh40VGbzX/NqFHhdw
YwUiWlS8jpF4mdJvc5FbkavuLLnzypWXIk+487tjPn2UVojFktOPLmcMLrCTLKnRAg6OfdWmYxmx
rwXlbAJOvMsGTrWzM+jXzDML2g1UXT+rUpdUxQlvh8+3UhGp6Z3AdVf+WvUs9cHi1jFFk9lV8yaf
9NgmoB/wVe1vc44JKUy+qXQohwHdR5POdxIcjzSTVnosL+jDCuR1wCLLpUu2z07LayV0zOMtV0ot
xDKGYFk62rtlEemzt9udN18qUV+zDfBZ2obsV0pFyZA9nSd/D8e30OGA8ls3F3X74QRForUXMnnF
+f2zPKa62z+eC0MgTGmIlrnhoTAV7nQvu5Y9zXxW34Ok166OhoHioBwd5PEmasiBtTlWILW6Onj+
VkAD9fhHqpTq9ZkFAcnVUPbN3b5Z1BeHLKPcS1m46AUeFa7M2JXD1ZCYDgKSQEeGP0crZLcfa6nr
jzZTERtn842UQGtKRuPo2P4mgxGtCSpf7oXhfWGpKIV57nU6xfn12p0Y2kqdnQ1aVUL8N4l3xeYK
5IzM8avSX0Lx+pSr266U8oGiARqPMGFcvHC/ZuzRfFtnHkmNHJGVkpbAsgk8ybLhhmQjC8Ynmikv
decxPd5MDZLB9dxo0pJZqAPMCFLNMS9TmWkSMJ3Tb/i6nTIIgUNFi4hfGiJ3emhHYDZK78gknn38
K7wAWyCd5PMRLWJnF7076G3hDWHCHKQ/RtXxd14vMftovBtKeiAbro3gMlZF/DHLQzqCYl3hXDDF
myTHe2ikr/zMep3VwDv5vUHi2BkDW9vvza815xH3meGKvKVJMa1wcR5gxMNQzyeI7PXezObt9tIn
t6GDB0+HAMuI8DZzvsPiXPSmt4kDKnqI//X+ab1IfDGQXIdHrZHoJQAump5v7ngOjR5yYIOZurdU
2bxWscSD+GFU4AxMt/xjikUOPQ+kU734aPKN8VupJU2KTQ7JD5pUaiZ8Dnx5oG9gGybp/aRbhhI0
u5odLzJOywHQlv3mc0seMEuU9doY1drKOh2qUWRY9JNuOD7wraEMAYWfV+fSXNnw6PKEkyxBTU1b
ALx9tRlTS3zrD0Kue96ylHSdY1uFBwzi+Ywd7xzRtCN07MSdj82z5vQRQ3qKvehsWLOm+S7Po0vi
t/X6TfQjFR9CsH7gNvt2xuChtZ6tdKw3so50uIB7K0J/DtYnHB73wg4P/7FB1hqMWYZp4WX/kT8h
u4fA4wkS/QIVvozU1WheVSAgmELoedwxyNz6rlIql1IwmG2pMDfhROBOEEdNlX0Tp+zk9gGcKmv/
ErI0dHRe7R2c6iMFDbpB2m0zwBo/OiUy9BabX1wpMryYItI09LKHn1CPXEYMQ5pxO4EYelwiAqG2
QCPTEtdcqCutxdh1NTDxcTAGt3qKpp1cifdK8MiqxKbCwQZDspt9B9Oe9mnFSF5XSSom1NtCChtI
EYEUimO4XlHu/zxepj+UosCZS1u9+8GnmAeE4XdGYWiRJblq0PdcpkLFyryk5Tmd4Edro2Mi1QyI
UlZ1fP8qixpbxTPfenHrZ1Cie3OpbHh7ApyL2zyAs1vwAc6KZkDoZvJ7OTAbpW+c4+T932ZMyTPw
IQw6B7KcHNJrBVNWbjypl634tsBkNSTyjKi4EP2s5puX6JEaKQUpDmMJVbcpZu9FPsqFDOq63mGb
zDCCR482I8UVBUHrKU+4toDLNsjXJ7DvhwTGni417eGC6WqnHL4ySzxB2MksQuBxgHir1goIibOn
fP8q7si5N96Tupx7B0DAd/4NS9BiJkTX3DI9GlyTJUaJbMdTQq4zMeOcf0eWqhcvciQiOJz8xPVJ
JKzVNVs7F1UvX6AKl+xZc+X7UT+QHmK0+4ibB5xqHXrRUP8ImS0wh28YOMCkYK/65e6HiUaog8xl
CPCa7tAge1MaD9xrF76WnNcPFF8SpMh0H7EHFlz6PiqF6lozyXs2SziV5pQdD1KDNAOOMNcm4Cea
pMwQBmCq4tH0tXeJFValAWEWuhWXMm8cFyPVu+Q2fQyn++43F486+gWnZ2yQqHl2TtwfXE9WmH9e
ZlaMOnUOq2NtHXfDdcwoUdCHVHiqqhM1P7pqxfECzkadLjY7kfvJGpYDyK+GAT/6eiimgweRkYb+
BGGQWRgDmxfGyQXqJY+tE+LGIDbQdIU5r+bfVSwZo9Z14Bdl5ckN20CEOkXUPggCMh14g513zwFh
I7hIR31hD7i0+6DPJ+rq049jyFvSejeNMomDK7x39DfbmuMnJx6kcToHa9QIyUh6Mnf+7tDJeR1T
crI9FuA1CvSbIjbfkcFqNl0CV786ap+xsL+0m/Uvkls7uzAyzyeoJ2jEiXcNBKQL/528qoPsV/ZO
tDAnk8qz37ztwcbi4gycdzDKM7zXlF4o5E1EKNWExfUU0mer28/rdc8oUSs46K+i4ruqvVLeGN1a
bLrnlM+tL3GogEJoB/Zke0YV8gQhY6+/tFPHnjnKQbJ9po0Hnzieopx2MRcwDvpocNK0bls0UkDe
z7JHpFUSfL/Uji52nQjA/n1yJCdPod1VNL2QspoCn4waFr+FGh3NXphObGqjxLV2Y8hbpViqm2TH
/6KdvxTCqSg6FnJUgA/FVV1xcTG28zmkLTjOyux4ifGyW56H0S1kXDgoRfomE3jNuIAix5tF/ltg
be2iB0MAgEq8ohZGAUBpSGm2+idl5MN6v3SGCnPnm8YTb0ZUxy88J/NvZ0p9vOMXAZ4au/Dv+/ud
j8AxREYzpD1wFXJf551msAeKh8hgkV58vVb739NQ0SQv2CK1xteOHTD/TrEewG6I+bZ51wtey9Lu
z0MUksqQx08d6lpUn3Ne7fF2E6kqS/dkIcRoiaDjLI/lQU98e90JN9QnzkdA/yMGEMBQeNKqzySN
iuMmUT3iNufeBs1K1Fr0t6C0UbSG1TzGLltnT824tMaC4XhhAs0HjrLBzVgSfee85nL5ey4uqLdY
OWC7BSNKFbUqRbten5vokBnQFJBJN+jkK+DTFPE0TTNVoGoYaqSgD2gxTNTRaVPs/SmK5u7lFPwY
Y5MDB/Sezbku0Gu2sPb3prZLp/OMdcdqQ5x+4DM4azT8un+9EvKWAcOhNCBsjIIzGp/bg+IDsFzC
ig0pAvHY904qCd7HCD3hjpOhsJE10A0Z50/i0vMGOHwI50F3TvW+ordxZdPNn6owvjmc1J9LG5zf
VPCSOtUYNcjzbBXKh2eotsnUVtHTdLwW5e424FG8mdpDKEjuQ4a6dcIJbgWejke+A9H6voN9J3g6
00DbRl+s2ENNG5OTkRBSYTyIQINnfjCvoBmTs/fHL6WByiABdk2iIP3IOBMwscIHGZDN1BDHjciT
i6UV68k0vgpp4TjS3EdQtKlK91Z38C6ncpW5R8NaWteCtmU715Dgo2tc4BgfyaQqisHq/4/th4EN
ezG8Rzuqt4IJE6iYvWqR7CV2cN+jBkHZDyFVWvUQ7owDnAUHsjWi5TAofuOhzHz9oTmv3Sj0i4dv
jzMcCdNp9ARdDKAo/YUT3gTdpWuP/bnsdj9QHB9q4BUNhvE+Ui4ty8tBw845pWas6SZ/6pvkGjmm
pxsDQS0vFtmkL11xaGLAMxBdWyjqKngIHZKKEdQq6lEB8GgeRhCzKrEiKOoKQMi63IaH8r5l+oH/
qcpNNJkbLTZzeHrgKBn+WwUOEH0+BALkwpMkbcUave6O02bHay2ebs2I2C6x45p1ts5U53sCBWK3
9kjR73Rlchyno6HCi/Js77cU74wEGb3V5H9JcpVEDpmQkzo1Ftpos/+zgo7Q+Z4D9SL9VJhHAwHW
VVAuO89tNKg+Hwq5q5CLucq0I4g3svk1vBdRWOwwO+lGGo7o59dpCrmyzf39iUe5sofKdMz8Gu5W
GkvS2XXw6x/ZAgK/RAOno4MWJSfer9ti8mg3skTaLwkookuudkwJnI/avxnxNhXpvaU1HY1x7iXG
wV8TSDP02ZtZwYO+eLoCdNsCnDbmu2Z2LgkNgs7K3zTtWXGyGiIvRUbk4PlMt5hLy0CGi1bpGLWT
4/W8WHkp/8LcFI9rJuORdtA8AlfQpKlTc4nhWTTMZxA6eBkc/YaF41hcMTQZ4LbEh2G6OXSiGWle
qFK8lvBLXdr4Ow2pTgM+XG0uGCiIQ+TEamCIRAqo2YhptMxE+c+q2TfrK8KOgLwWa+Y3sDRF9d64
dnWQZILIKcl8S1KcuCQzXEMjoTRWjN3dyP1pkxYooJl9wskasTbzTVZnqB/7rYDMLm5hBJRwdUSF
Q3IcdV2QOw5LKPseha8Ffsjz4hQvvATuGJKqoYGqRifZs1Eo7MZyc67U+VcTIGel6diLfCiPLMrA
o2kFXawqmaAFtqZH54YQEz8GqvjJhXfYNxieLCAkPlnOpzZxKT95aVSqVAWpQfhvmEIezAhyQKoK
jkZfRtsCDYcwBVshiEQ54NM4TkBfgqyD9iMPUp6JNPBAlikXrhZZNlafVKLbidv9o2FmpAOa2Poh
7ZFuLUb17WQTMckKx5PUNd/6U73NwhMNrDRnilaL4QrARrYjp0fW/AceXBmewzDVAFfFzV4y3+87
Weotr3oqvWxVQGzfCBZErrxhEdN+YDqGZKCzH8C0e7Wek5UNe/wAQhe/txX21HloGSqLuEUlq65Q
hj2dKTW0sgE6XnEX49beTo9KYAbZrmi2xIEW4C+TTuPgC7xQJ9uLB6iwZPfvThb6PiyRwZkqn9zd
XVDnz0pg09y9at+VRl1NfTWWPYajMjbv9XASIBw0ZtQkTnmgt+pjuYxl7PGjoe9+bu7I3jgf4m0O
/11+DH1C8BxGrMef0eD8L94M63Osg5MDo3pYKf0YE0AQ8qVtSMqsBrc2JYPzeKyki2qIAQwpEx9l
whBVnIK2TFQ3gekIVR/2FYCHOeSJCP+XY6qIQLXVnKI88vhFDpMoLCHZzwQhJ3eet0/MVQfHR+94
z3lJ4WTMRW2Iyfel+l7tbpVbsvdBL6/9iIKo31iRVz0gAui9lI14+C3DYu4wlFBnN4Hx6pS5/BGw
6V6PoTVg67IizCpBy5i3e77xekcQHdsLMy+23O+0pT9TRswmxMl2V17ubvzrYT1BpQp2atNa/y8f
tzjIfWAanrVn1Rlk4zHXf/9f6T2XnIjkRHjfzLbBuSN1S6pC6UPdr60yxSsg7IJdxWDu8AsMrtDa
15vo/niRUJT+qwbwvwJ0azcf0ZiJcFKRcRcPwF/chOE9/gVqCzbvfZmXg6bHr5mFjhh1L5lM0qcH
rhD/f3n5CbYZHant22MFQzG7blFokcBIWUa0prnr3/VOUba/uxJWdJLSOEl3a1Vmc92mH3537x1B
T6L86BU0b0pdydWEfb0TBCS6pUY24zAoSYjcfJXRPaHOXUKaYrXP1Xh1NzBRm+7q+DeHC9Fu1ID5
mChW7xqkXgraHmxZatABrlW6Od8rgtXfosoGsoGWawrhJZif3ZS2nMqSKMD7z5mikpgMPDXET+ef
yfQFrduLwhrpqfAcsVF9TPsvA3JLTsyeVrc7fpHi9fYLZHMNsdCITS6mVUf6EUtYOgUOBHxoDnH4
Y5MP2zCgKpFvM+J/k9tyMsPQ9/+1YInBa92QUp60XJr1ShEIePjchn5RyLKAMyPExUIGcKHQNMcU
LBN9/N/97babNIv0wqGD4B1V5/NHDwGGL7KLoEnnOwzXP4bi0OFgpCTJZdL2/abnQqGbE21KV6RJ
iNo2ZZyIIW21sC2JhOTRMF9hb+CAplaiNZ3EvnGuhoD4wLzhtXSQo3cqn/7kfSQc5k1HJkWWGcJ+
JIdO6EeRQQdqkyu9X5eEsRt26ZZ4Mb9DaD74N6qSYvKly3H++UqbPPwxaQz6fr2MeohZqKAzvYY/
SKd8/FNri4BhXynW7HzbhoSvW8xYnnCz5x3GMkX+Y1OQygSruVUmtZ/BRaso0w/1ypR8lKDtgCZB
ud3w9ceJCM61rqzwlUBD0wiLUWJBvgYw3a4Bh9n1uwr9mI6iJRDEgLvu/DshNwAoET2lxH8+KjBT
0IKyZseJUoPvKxH6vvYeT7feVZ/ddu0uMYRuH/1n9Mm9ECjoYHMQO2OcOYRk4ddSkajjJgNK1WsM
xdZjm2RHA+lund7uDKxce00un9r2mhHghPjiuHx2DmkwLxwgrzKSIiYyj6ZNwCGhc06/PAHv1iyP
9zHHGkAMrh55syGKkm9bmwICe6EGO5JCDEeg35odZ9QIPxn7ZqKcDm/mam0xr2CeFyVLWO/yz5Fj
h/FcuXnod27h8nKHWB4x9TQ8dsyFQhyOiNV+hfe6TqY23rXLZ23VsWhwC/i1EX6W0twUKlLGiyyu
3AAPmDcauPGiZdp3qrMGWua1gzTijlaq1QIaWQw/cLXcaxDqhggA0J7n/ts3zZyH23UHwZR/hYRw
bG1/MBpMdv36fvJzcxsSiPfHsOnnX6fnY0HZDz6exegWP4AiJYSHUtWNizDnyHeHuAc0JeAy7ANj
8f1d+frs45+umqPrDXKfNs9DYgl3lbqv7LAF455DrtdDKVxnQ+IbURoJKwGHXqPOi+g7vkqhvn9U
dQlcTlOAxkuiNx4K0avgqLDHxI+u6w5QagLMN1a+gUbaT0DPVUw3kISqO/NF0vNqmBb+HmCWDu+E
N88pY+oGL+PJulrfSmesk4+Tx9aHl8gFW3xEPtvSJsyMKWjm08jUo5h1BUTOQvkqygAhFQVb7h5b
TJMSXyUJRVpI8WtapHiVSa02UUgtUWpN3edqh6TY4KCB1tu2m/rxH7k9IEppOLMIeLaK3Ensga+9
Leh+Ce1hvdlwiJdevZg7rNEb2yNZx3FAaDahelBPnE+EBGNavVMiN/Uc5aUluWLiEQqcgioZlb25
XKmMaeu5XGFOFKKY63t2D7De4y5F3RXJKhSC69ktWD6UcFYSYZnoONO6Y6nVsMSVCM+PvjD5lZoJ
WOVwFpK9RzpH70p+OmDwOux26VTodSBkznuevUoTxkzNFCnnXECEdXem/0eEx1opzQOlCet9M3jt
lE+pALioEeD+3UPMAyDYPvu/BsTz7Zn0efRmXI5jokC1zRMGn4u8tUZCmgbgBFDeHnxJ8rdqvcBl
VBW3vhQ3vqrA29dJLTLREboxRzc2IWFaZ4KyiepbKXxB7PJwZEfGzoWn9Zz0yL9a/f563f1tc1cY
l7MI1n4xaMj35hsenqb7GEPpGJW+7a/LZMKRRgiaxufYjsCupv8he+JNIg29n6m9NfVCzahDR8UE
hF+lBog5XtPfLqbdAg1MzkHZejQy6bAeNkvvg/MrcI2Wsn4/dNj8DM4iB7NHSz8PjLOO+/b3/7pl
aokfCqh8431X1W5nm04FzbVgWfOLHqpFxZE14ByWNLzamNsP5dmFr8BE3enFKye5lDmh4pU+yh0A
3NtRe2Bm/QVlYqEmPewVwltlwY+ODCHD+4on0QYHNSfpjCByhqBJR9KtwAGAG3xztWaBmz5Bqu3B
yv6K4gVZxSUi/EoZKhZC9239AliPuShP51cw9Cpos7pu7mr6OAQDCSJGFVXt2p0u1e0cyorxj1Gb
XUv/JDayg6+ifshuGr61VgedcWyXEvMak5V7dp/nCyIP+TxUPgc5O2EX08YVRSnJ4AWvxqzeL6xy
2nHRsqhY7T4LS9AmuIFw8fzOozmPmUhRNQkATW2uQazsVat9QFSfr8ZmfNw1Kj6Q/XH9IcoWJmx1
7boWRV5NKhF19mOrP9VPvZkJ0jgx42a6My2JtEVzlVPUuYpdViUTYOI/xfuJKTwleA8uoOGADesW
a1BaMc9363MciwVhtfFgWG8NmW+5bFgZ6OMys3RXpS0SCUhoOjBHZ86er9gy6RieGMNJXf268+f9
QBDY9qvyMVdjnfkLB39pXcXtiWTNkXQEcM4ENl/IauDWGKZ/3YPGrk0Fw3Tnw4rqxisREK2kqt2e
xeKeXQBr3AO5ROyRJ5tkdn+T/0S3FE20YA8NFA2btd36j4SJl/mB3sGYfEHkI5qT7Ts5a8KHgOwu
5FYcj75sQPYsito68g1thjJMuTSRdNvzt03CsQIsvVBiREhPkG1PkiYeMYmc7eEQfcUVFi/YZkMR
Im4VLt+QFyb7vq8rwI62zF1UsweMKzeyizf52Z5ovSQ+Hr56xAqV/ZeZniC1QOzmyTB99zYVOml8
sSX5ldE0LP4RNBzocIzL0u082eYVglbmS1WX1Zj93eHfLFPvCxRGmBoHsh69bjnaD4jXz5mw6/n/
O9Cq+ecBHMKOyDwSGAzI5n/4nqRlNkLaW51/7NkWMoP1mKNtGZQU6nyPXfGTOR/UlWuVsBLaOmQT
O5ISVD+FW6QNAcVhk0qiPhXdziSH2qSTBGujbAbUBuVxuiizU3ebXq7PIaCoJ9s8s0wGFeQRFsu5
uUwsbnyYP3c/hnwoLCClFOtyoQrs2HIukpeziiXShRwRX84/+LXrA6aWA/ZtObyVPkpDo7LZn+/5
N1Q+jfgKOJnr7zXhvWecwUdBByeHWNgaGDgd/4Vxsu5GzP5ga1za9GPF4hzKGHLmYf8KVaFaR/1j
TfoPY0tulXlfda4ca9p7HwHjfvmqD2YcCUn85ER+W6BnJkf5SOeYknUlv/tVHHH0glmCtzUC7Yzj
LUkLqVcdUE7vsG0Rwmozf2qQ48d+P690STfi+w/+o3GRgYc5Urn8XGS29aUKUk6gyvPf5xbIi0Ut
VZtq3nWXjh9WoS7Y3p/k3VQio5tXODD90iAQUPvaRMMB67ZTFd8+rD1OwsaPDh7UUB/X/uUk4pVH
E4SrBt+1GmjZNGIy5Zt6VFoIdgdM0oKhidBDLQE2FlIx6OfQiDDpTEVj5fHiqfACSsF0VHup1m+h
LtaWrLT3IB7NBuKMjO/x+PUjXNVaQWU7cbD9sI+HbQnxc6Ghc6YBumSJ1q1iRDHpRYrJCq74DWGG
9YwLyKHsk4BAI+NMtg0X8v+PsqYwt/2l7lGVthQks7MlFsZoYygZfqZ9nPM53L3kESvitxiuguLl
Zywbb0/OpungzPYRVEN+NgQgkKRqu71E53g1TVlmnBIfrbxEZwBTOSr5xaEX69jPhNqdFp8vXb3G
9BiS8mW59SlK+ZYl+OyT5CXmT7yPFf4Le/baAxROencJLixk9Jizkh5ZVVu+GUew9Rc8s82Nyjol
zk5e1DFE7n9Iza1kCwbUFfqoCnTe7E6GtcRRrp5sPiR+EAprWaBjUk5g6qjHDj6UuycNNUe/Iyji
xZ4j0DOsT2CowyV90Id/zgOKLebT6LhnTuDQIzgSeZeAUi9n6MHKyBdVyv0KC7VP82wfEiyBubg8
jw6DBPLfTc7Yv+LIl9pX5e9oz6lzp49GcRB8Gqbt36nK/UC4moRVxuu6haWcpgaHaBm+pA0VXc+M
+UZGYqrqvQ9kUCOcYOnSkFZ9ILdU8ylMDp0yGashQMy7aM0LF1STr2KDNjbUMUX5i1zhCZC5blLi
gyRr0kBbEChtJPbY2myor2HzRnBoG+FrvNgtR16tjBTEsZCLfU+avNfKlGA0LmQie66be6LFwMju
u4uczBPBtxkXg+Ksd93/KxJnGHU87IeS8nC3b/myK/6eYo9D66GBpn6li3igcHXIB0ipHP9IRhP8
FVOBFeOmav/VPduUTi/iomaOyx6iVr5qkTHZ/PYsS6SsKacBmE0Q0VHSysblbLtuTFH49c8F2UQm
UXJN5ptVh2ahs3PNwtiQtDKPFXwxNo/xqrnhbEnCC0pemfjotxoNajow3xaokWVZJPqkAYPpBNk3
GFzBlD2TmD9/TBnRp6kzW47AxzcPO8RfoH6Y2SserCkJNf6zLetST5RtcErXgVtJeC1Fo43lz/Ac
1BtfgdtTf5u/q00ZF6LOh0T7kLXciTCza5Ukf4Jr4mYpZaUigk+6577rW6tcFObbYTA6Zj68h3c7
QSL43RAEASKItksuwMCTaR/MKYLCnoVU5tYDV/j5Pyzy/+mTl7/FFl+l1JrxRViQrJB/bNuKpaS3
qVkLFADroWTxU9b//GC274Z3rexWIdo7EgsDLn2+OU7fVOVAFVpZCmZGzL7oJ3/8hbV5+gi4e7ZE
jPfHS336qkO3i43IvmzA8W704ZvRZ7lbU4Uh+ucZgP/vOLLxyo73F7lIMshN7YoHGShlBnQDtDXd
1j9bp0HPI0kbFJYBGe/kscAuORtJNgO74w+NqMEVXvJVluX5ZNhZkVGSf6DsOhEfUB0Me0zBEYXa
es4DX2FzjObTDb/DUErqXonn7LzjUSAJk3ju0fxK+DcioC8U4PwDEleuxPdZyR3jOf8ON9AJ/ujz
geDjYt9/s/d2afE1fKwUdSV0bHYUOtamWyN7aTLB0HcQ3FlkaMLII/P7S3N+LPojQobKzlPARGUP
Z8mY/tpeP1jlHgHlUnGYmLe75AtOEVnly/wehX5Bj5Ws90tHl2BqtCtyPhVFSQziCaO/B6YOpQ10
xBWio0lsq3xXgqpRi6fhgdT+2bGkncimsdZTrotMSzNurwgBpCQjfh85qQHc7VIPN94PJuSJSiNy
1dHU31fhm+vIZU9yzcPo9fRFvaEr2GUs92ja9V165RWh7DjKR5jsodTV6uN0GUCptuMIIeb4kPtb
+3C/S7JRQ5eYW9iM6c/glzWbplbpstVH+EU3zRFK+geYAt3LwCAGU1UeAMAf7a5AuWdz45M8tgVP
qB2j/AOANV5snE5GyqUnHIInijgT+a7UtMcivqpN+gUHwwQ+4EuTPFGiMCYSlgu9XzPiX3u5MDJX
QQ4METdruitAsJR4HuxpzkEDH3uoXV69oaOJBl95Qr3v4b2iiU32FGTMcXtKNkKpbj55363mzUmE
4OkDo5pTK/sLvYk9gaTtuxRKBww2Usc38RQmJaC+pdMZz0zfRS6s3IakPVH4QqHp+QKIG9eJ715k
otuaPsb/fmWJAlYQSGvMY+m9xKPX2kIeJCmzDM/K3sXpGiYqm3O33Z1DGopZIIP7TFQb6x/ryvlh
NHG9WNln27W9sd0Rt5NWf/vBII/6gNPg4n2ExPhOjsOc+GPIKJqGMN6NJu/RtwGk3uhgdbvpjNLx
4v5vmT0sbABImXOa6RHfpEN67DSo1EYVikyJjNK1W2NmGxq86Y8vru9N+VyPK98Qsx47PsqrZys+
9RJ0NHxTtAgS0vmDpdt5todNf7BUwkjpmtlcCouXvkPImTQTbxS+TijEnYSMWLNFshbYYroeiOos
TYFZUtvxS37Dvl3ktKzwo0UfO5TdnHGZegpavmjV+AyVCsFfjVDOVTCZlbX6a4eh2EKSURaOSyKl
T6/gTeFpsGS+/tt4Bi7Gsnz8tBwVWzLeXFsagFX7xz2IzUJOYkwWtkZS3zmU3BKQ7lbe7lmnmDU4
37e9PCKeESCWygq7eK4iYm/JucaNSJc3Ne4UMmh1lcc1GybNMH5UmLTlRyAZy2QD5UeIKn/UMUkM
evsoKupu6Q0OkRKiE32WJBEQUifU4tr5RsLMbzA8gQAjlF6/z3phTq6KVFz4CEOxKlqAYVHjmb1m
1yqkPDZlXXJpWgrHG/fZLISV7ft2gsmskNhj7lpmxeA7dC+b8+MhI/15MwPXFbL1EPuwV4dYFOUr
3qkMm1GwQyiwIIxUfAbi07U/bGH46nM4ApYpgu2WNPW7ZfKfGqb6eSxnWcEWqE1GLdQSExYBV8T9
KGPtPuRw5XzVvmGhidNH92qjcwhDcTO8HuYtZFSBIKXKq/pdQyd+Er1ye98Z1yEB+MeIWXFHBinF
WOnXuQwfkCJINdO4vA2Mv/CbtXB6c5g2DGBdN0WHcNXtmWcLk9zEE/vnEKgjbOWU0t8zKA+l6LiP
D3wEJCIletESKs/6duei8yQKHvdERvx+Iz3gIkctjccMZcaJFfAyxzVAFUClflSrKvRzxN8bE9cn
T1Ul08QnsLgjhUSRiXWf8bWuFw9tNFyH77MBYpZsw0xDojzZmcpk8HkzhOjXvkmjqlGjaAgrkveW
m3h6scxQ0avjkeDZ01rEnQkTgqq9LfjBH8jkwZehlZXkYuXEXaaCzsRn2H3U7su1yBlF7BfxXW6N
NqNElj86a29MjlZMIJ/T7aSaz/VrtUNFsdE0KywlpVjmn4X/mJRNCfES8AeCAAiiqrxCwLjS0yET
tbkUKPlh6t9zsaFxpkrxcfRX5V99JA8UKvIwPYO/wKuOKlZgqBoLk7ZDtx6bcJkIo1N3rzhvTHBS
OVH9h56nP+RJOomgXRu4pe4YxLt4/JCuVnHnsks5jcwUnN+igQa8orW0zU3YlbKSXnzHYAwDaEKv
WdJ0KI/x39ZFAvJS74Xx4uodnNwo4ChgOFnw1f3lzIsaqR+We+rT5UGpAzqY/LlaKPr1r+CJz2d4
jXlA8a3h/zIZC1wo5zWuPDjik4lB1M3LytPXhKiS7xPIKYa8z8hYbZsKaAnUTzb/6Nb7s/tRuJDR
rJ8yoOU5HRJlTrpS81abOlXt40G5gOE765C9ThdW0D5H3XHweRwQUe0Tt5YZlR3LsU2PaOXsAtEv
Mwke5L8JVJCGJQwyzPX2ac/HLtPqartZm9Jz4Lxo9OCWoKUj5IT9XQv1+Y7UH+SD2KTKNt8jIabF
0B39Wg96b9ZMGu7EMQl7BQb6EV8Q6Y0dWMj1UAAPi7fK2oU858Evz52MbHrcbw37qNDJi2sah1ox
u3aaStaIjXMzrj4po7o0zbeNSabdtIfQJ6/r8Ka61ZCxDk6VtnHlLmuQ/foSnIOW3OkT/hf6EYkm
KyU9rgrtuUua5tRt3v3ebhMBGh2ttITIj9RCALWbXtpRUw5O/wqmefjFWQw3ZoHL+s+P95OOyiA/
GG9N8qUZyDuo9wL27avUTnz1lpvwP18FFFPmj2M4hg7xO5mc+TQCTTuZz6XYvugXtgkv3uC8EIPx
daKsUtZPBQtP9fcyf+HTYbffM/6WoINW1hs1Pq60zSQMp+o1lXh/kdJSZjZZjFFl5I5wec8iMbsZ
NKQvPVqdM1fIifbiN6/5VhLNtgk7pAzh8FNxUm8c0tQyixxdhsCRQGXiur+lMAiL3f4QhbSvD7nO
bc9+6m79zUHSve1iYz1JVMbWcXwPskIug5qGx7ZkJddpjB7IK+qR6Yuk0VnUekreK2ICxk9q0fcC
1lTwIDcCH27WnMjaY/brDOeA2GhF022RC3d/UkOzGq6gN8JJAAQgb3yw5Gt+S5A/kgjWCbMjSLio
iwokgU0NMJor7Y2EUEFAhwoqSPgxAPiBh77tqQfS9UKSn1+nYEs3XyASkYzSGLdtdm1z+nEDDELm
qaW0pDMuazuDkQSJY9B+DoDgwgVdgDHEXoMDTZM+MeDccx5rLvTus5D3iL4On6wt4vSllaZPd4cX
7ONNkel4yQn6fPT14HmqkFBLr00pzZxseu35CTX3xZbNZZeHwHH8X3cROO+ZudM3R6fKfOG+cpYr
SdejgkO5QA/etVgh6FENZybgLjVi/Sd4P4Ifh4nJ34WHuOtznvx/MxNs4wrIsQJRZ/VdMtqbPFDg
p/DykDQipsAp3hyxwOEkg/92sHKYHPPwFnJEC9zzQPR0XUlFiJDtIntXZRFaW01kYdfOrVCHKl6S
Y1uRKJSj7yMAZNXEoWNLYHI5QMUURIlPN6dPIaty5DHjd8zrvqihlVwVs47ySfw4/+q7MGrsQ0Wn
MV4zT1oQHA0TtZx1brNArRkSCz0RO8UuUNg/6PFCSfOW65cCELxzV2iIzo1oTOuJcMsmvRFtudTx
pMQLZbCY0Tq2eT25PkI1sTdPdnFf3//AA+GUk4WtpAHNoFiJE1j1U2dNby/6qpoM9U7GL/+0D0eI
aY9Jmx0Z0O9bMxpVJLqCUmCnsCHyldqfnUMkO3rXDGFe9z96Y0WpqBXZ4DVUXmMXvmXY2WvMZuMV
0uAcd4gN1lab5oCmmBvKHqqLw1UVFuAX6aOWu9KFfkHmezqa+UPHi8j0ZIlbFEmKU30gzPqTMhTO
JHh5Z6RESkMh1MhiNx170g93ogDYnMLQzQGm8I7NlPYckMXLZbDyiXlSCi/jVOl+DmJ1AvjbGQh0
9d5xhn1KpZdyGPDBtdhnoWN2qbYKagvGpguz1cErHBekxZOXGDHTGQRzm++gBzc7/UGGiUCjdbIu
7VNcaXb/y82oVWWlpLX1SXlWdYSzY+sUJ2ktfUiO9swU1WSUJgYeN4iVp2PT7cWKlO5rc0IF2Eyi
ZnNQ+T4uENI0cK2/tWwMKgPp0nXe5k9yo5qaLy/EexIyJBGHn9OPc8UgKc6kOOHU2K1E7hzWJ3AU
vplMk7Vo7zy8mUW6bNBLiCIgXz2FBkWg1tv1a7ibNqTc/+PmUUD14GtZXMDzCoSEAB3xEU0L7+jl
T5DLF0SJ6SIDbf9qoYLsbD8fgpZkEnXyOgHVDTD2pAU6LnZ7NyfBM2/Px7mI7ykrPya7GJ6cesaR
xv1OAo5fIfGc2b/dF+UvmI6OLuosoxE74JBDaId9MdpprrytDnT0O7bNJxUEw9GxzQCtJqvRQdrq
mfVyDot5FuZgtRC0v79IEIEgtynCPMm0jNE6mka4vdaO2v3rYxR7Y6pM6Pz/EONXfuC4KMgDer9N
hOsJFloeyQPMEnFOcKLJ518AXpoKMbGmMRnWFBww+h8Nff9jh9eU7t8a0NvuuKytC3MUZgC6jL8u
hIQddsUu8hSD4VS9C4TV9Y9/rNsvPp+0ojLuJ4lBgIUMADgrueiVz32oJI7cWemu98MyNKGkvMbA
dLDXbLVvKb/EdQ2J8tjw/9ixqKqRgzym90yTZ5Dlig9sMkqZhc4iGbOEbRSilaSji1TKgmJUUqqB
rVZgPpi/0/2OGY91FU7a4Am6SX1Fl4ivPu2MLnK75P7ueHUUOw8j867IMZoefodbNUuCrMiO53CP
+QsknNLbX/uN0RctYlqijWeZyeXdf6DUr/RzihfmYTlB2FJhkeOyOziQ8lGfatw7u03xjMqnFrTP
Qf55E6PvCxic1hzk141bZmLEND7FlVNhZkzyT2SniqADgA2Rqd3nSLT29jaqUeV3MSd5ufh5D5pP
EQ2u9BaIjnhvlfXZYh9bD7Q6ohxbQL+YJnZHRn8I/QP1pVHhGz+lmE4aqvLcq/6oz6I7mI13LBIB
7q8FfSTT/OG70wONkrZygDFzsAx0BB+m5rL01kLWrXtfbRkNiscy412RIMg2BLQNKf68znwtFYUh
KBq+TAxCbNJKWNm/7PetOBzILhy9NTmaaVXUIarqfwsgT0QjtD8I2QfZx9QXT04Y1+ADmhgMVnA0
jgPeDRfBndF8AA/Y0dvT8hi3mRKDhDRywjWB8hQvBpqguMZFW9Gz9IglgZWNu2vkdW6nX+NcI6zA
Sz1M0xC0mGmfnVLBcCcOnLVLI9So1KffCJzs4jWIYdSqT2l2yXDuGDYRXfR07lnwEWxqJ/SDsEMk
d7GW6HRBh3+gVRJL3LvO+Fg3rPpCyOx3O/oKe6le000M8enIaBh/FQ9pDKvYxrw4om7k3U33kxPD
gbQXslON81md7lE7r1UAtn+d3igytmGEJWCqEgbZbGB0awESUwNWQpfwiMaAetbXL7L4OXAQ0NOw
ZOyCG6TcROWl820XNMYTbdoNp7mzv12VXx7i2FZHfaxIMfuGNJJEd2ci/HYkd0iiWfA6w7X3YQqC
NRAWs4HVeG1Ju6LecYZat+Urv8HwR8wik53Ye4mfiR5ORlyp2b4ydBjQUMC/2YziDjHaYoEyISII
mxqHKDEn50c9CUA2M+M7qsCwh2lOYT+4VRa5XjXk2vtpqtuwOA2nMo2rh4apUvMt9hEgmuooZfhs
virWYjySq8CenYlywrCXiQg7+Q/uOxO89Uo62HBct6errCZnKhybs6reQzfdlZnp6ahGpavRVYlz
HmfVzR4Y/hlSf6ZHwxaPbx3WRhMMYUOifJyI1P4D7lfsEMbhYKaSI2gFeMc4yoDSJ/2HV37+qZmE
gBz4WdyzCc4OG3xO6CdRHgCcObVHWScjrOO+d7fmjUB67mOs7X/kxyO8UTRds122GBnX86l1pH8J
eQuQXpjJ5+Fgu8v9ivIKPxJ1HK+WUpoN0R5mJK5RElfPz83+KbaP/huVB85C7Efr1IK2kZDDaKJ+
vUYOIKVSTp3tCart2KI06DOy9Dc5jGi0S8w/yw2TI2KRE4fBMWoCWKmbwNb6Jm1XVefOTuI2cQNd
JptW1T9Pmqofa+viLK1rVCE9yPT2mpzRM7jK3/kTbvLXrjhUjSWEOEQJLOm/31mVUs9pbHoZKuo5
GLo9QowKUIqw/LXxQykw8CiK1Zi2T4e7G5GAipJQDYuQgtGnGjiOoWWU20TbOKFmyWf5eVwgzlvL
IR2nnqDIFpK0KeuZIflRUaQpHVQDLviwBxnkWn6pDQ7ow54yUh9W8L/3VDsAbpgZgIowgimebM6N
knf5JRIHSLWcFcUaQwGq2qSA14H48mpfGzI2u/AQLHMERzflpffIjvpF3xyZ6RThNfDrx6EaM09u
oU5TTb3H57YGXGcguv3EN7HCibiGb80hdsOgQiGq/KrVxAf/UETiiDowhmhQEzI+h5MWXcGCJOih
URx4NPe7N0J1zFRmEsxxrhQu1/v8yoz2OWB/uobRpEqXCF01PIwF4P5r3PHJlCv7qOPF6chQYF9b
RLV8vh8tygiJugZ+9Y6LzeoSaxBTJ0c+9tm1N2ku9cvwnqFjl/59uKcqASW4+cqcttsXhzF/B0MM
eDmRUSEM3m5KujJ4FbTUbB+RlEp+o+Wq4+FUFx39sK99chLggLAPSOCZG+ZWiJB1aP+8vRRyI8ZT
5f8odaTcxjJP9rtB7OpBPVNy4556rfkY5u2wYakS1xvjh3a7hENQuJW0NKuGUHQr5wguueXb/qIX
qj+ud0Lx6qN0kISZkgoH/8GJJW31ATEh7Q5c63z8sUCjQgCUcKnvPFR5mejfAS7F9SER/V3p6xsK
ybSpq043l65CH/dbMDSjBOaQ0Ss1u9qneaKe5EGDRTo95xfTDOXgcTsX3t1gNSRM2BW+SG33bN1o
kq8duLSEdlAWQzsdQPf/2fm7bobI+SYsVuCeWgrtUDpCTj0x22+FRgDOZZwtMsUaEjX682CXEERo
jgJBnvxDJgydY3cc5nAW29c5nrqTBOs7V9d/SWAFYhun9MIRBXDrHa2pZ9ys4txRlpgDvjaUOkF/
lXDFLc7M9CMYRXhej9YL3+ot9yDY8oy+Zvry0yQcqv1RsT3A6MhViBN49Sq9vzjotx2PegIM5NKH
1E3mEUuwCgW1kz3bWDk98Mw3jo8lTMW5SgQXr7az1hgaxYzyeUGNULzEwbGxjq/yD+HTQrz/J3nd
48mvSTOXUdx7IxBEXTzDtE0FFs3NyvXYJhxHH8ZZIZoH8Mp9W/zu59yhxoBwtWLO7UDwoG92U9Ra
8ZkXixuHapzS4mblxAY+r4VfJ9RGIsu9xWGIMJEUw8gwsPykB0A0YRNQE0G9XIZ1s4A90JCZwTxj
zfcEkrIFgWO0+Mp8Eepq3L/IoUcfC6pzUddqZsAr5leznarH2yn68tdwjdko3ogbLqAMl/LRK8tS
GLttRC7Jf4SDOE1vo/3R+7I+8fdTG1dRXfeUyi4W6Mttum7AT05v1qa0xyI6MyzSc0NpK7A51gpo
EhFCtYdvKUbH0mnhuQiNpDK3GlUdeZu2Yx+G3oFNMXzvY/KDqolAWjyQdQCQnjtTWtdcaum9ZAUL
wrYV0ox53LrVFlOFJkddySnyAUTUuA5XfPYURkoWrj1VKiJayfoRhQKhUeBeAsVcyE4OLxmIMTuR
DFRHyhQ0tPh9MXek3QOgQ+8macvyKq/CxwzvnxVMTpvmVV239WaQG75vmCsri+bl3XeqhCf17/7H
+VWodt09Ifo2bXu7JMz50a3UlVYmsAJOPXrjagYl22dr2dWUQR9eEaPtGxTL5HVwDc9Ni1aI0jsN
n4w5diO1tGYTBGXOnQoctLMRYWMAs+bEE17skshrVzRVl7A2kgmx13tLOFgXgvfPUHHrVa658Iwj
s+FE9mXGOdUVkmPZjr9/i12cdi5t05nHKGT5qcllWY6e6gQhPGLpsH7GreqSlpP1pwnPWmTCzzbi
QUrzkrlxRjzSw5jM68LJTsUiKf15JIbqrED6SCWBH7sdLvneN7TnVCa/TLC/0Y8KatzrsstC9Zga
pKp2bTzkqF6mIzJ6qWo4mFKLXklQ51KcW9/hVcBs5H79iw3Ygdiy8YpU+J0WYDOlWfbq5t/+4KM4
UkM4X887JFWQEVm0u2UmboibzqCDccx6ju7EUD4pPmIA04h8RTMVAmatIAbquo6ep20Jl3k4i4Xy
TMcYv1xiPVCILrqSMpA4tWIj+7mLYHNkGuRVAAdODnIC2hrdowS011bxm7s3McO76gW8RpiQ3Ez6
WDrZz3y0Xtom61BozmTUKeOzG3qHPF1uNvuIy6xZ+Cy4vVdtVhzlGQTLcAVn0/CDKKMyktQOTS13
ZK9gF8bNTb/h2AbCTCVRpZ05ywR+0yw3SVLEyXtxzEfFatmuKOuv0Iurwk9naHtIhk10+CKFkT6S
W77vkLDug60ybVX2gsWmUxvfvm/IO8+jRw40iD9VW5UpwkOyNcph2t14WF4iSyHZlx2i8u1K0UkZ
6sFMujXSNvdaYo/et63BbIE4VUktWTJn9i068JBxxVIep9jogO2ANe5mBhbvd8mvj2qAD76bcBR8
biUJU4l8ytlfsozlgzYhDBn9SkuS5/zRMqPl4OTFtKAOl7KOFhf/ZOZRH3K6/BmtT9NV8mp3LZcv
FCPnF/GYXS1JGCuJ9TKjetRg+19XrdT44qhvcivUvmqS30xa65f+kAfyKShNm/FmBqYhi61oOzdD
drWA3OnwPUl+aTzJ+z/KNtkTdCPoBeFXI879MLZNw3jxkxQQ7rlXGt+tzczmRihNXcOLMgegMFRB
nfPRsGMSbJ6hSYTRggDE7vw2V8jsvAC5qDoCTt2U/w7KUrc/C90v5LoDJvYajRxEjQPrDXKQBNg+
EuM3bLPr8I2iz2YZMJRnbw/uuVMCqNE2Cn6qr1nIhmFhMUusJQYtDXb2E5NOAVTRt4nUREZKO7GE
UIXCO06I29w/KnvRkVb5eht5ikQRbC9uK404W8OGL+oTMAKvy12QsNM1GY2QddWA4mjbNenc8F2E
BeLHxDOiVG52zeIXbXyNO2zyeyUR1DoGNzZSefK0X6oFo+5q6i3L0vOmH6pzXYRi6gSwBo6Rnz18
M9OjlRrS+CI5MC1OX8pup/VRUMPPxid1SkRaEYhUdon98NJ+qeMi21K4Q3z7cbLR2StJh69svItE
F1Q5CqvfatZNcfeDR9AHRO+jwocGU+39qv7mwKTfNz60ATKB0z+PL9LocAVcpNFBLIafll/dTPMB
tN4OT3RnoPkOpCU2eeVMyJt8c5hWcO5Mo3yBtQhQRhJ2mA421x+YnNnO3+8dRjRrAT8vmysxazdZ
bd6yFtaoWhgpZEgXY1Bs2SS3a4l7IBF3uq+iMWlkDcT+pJGKiWgozLEKYuaunf/5PRCKH/UGGF4p
tIEFpUWa9snpsqQxM+mpR3HvPIJOmWLpT1RLvCC1/iGHuD03MgFrkb6gYaNLbGvogm0EPJjOax+1
qLfz/M6ZJdhpD1dCryi5KOazjjC42SwpWmNeZ0EgfhkqiP8n2arN7qLHEWcaQk/a6AQgya137dDQ
/S+hwSrLeIJUHlnVHaV9zpgFn0HXF8GRY89dyDXjGkhksY/jQkID7RxUm5fdj5XtWyrhLe2SbBFW
JRC/IYYQv5eNJno9OYHMXlCq/81cpzYTGhqJS0hRVbsYW8F3vJ1BKJFo7fBf7cMSpirw9kaDtIQq
BOKTpGtba97sppYTeQiUoToSrmpUQVW6tq4dO61ex9kFMZWX08z+McxMLw9prooz6GpJ/LUkryP5
7yUvJYdrtLdy4qVBhjm7EJ19Pzr9lqharDDMSqfiEWyEzsHc2GObgwmf1s/6F6Zfo8Lp4GVnSZxI
fmMQhK+q7yuQ6lw4K0F1fz9KopzRZ6eW/dJer5rgSz9fp2nMFcvpD5VMMXAk+tuQvYYAo/w96Ifk
6U0HuUhRJzmYrI7wVWsfeptK4EKQkoDiZOekhzVqHNZTvycQhieO8YqGKmWbpOSIwLgikBSZbrWG
2kjWmnoLGutA954E55loHl0/tkcSYY9zR874vsEe0OC33Qskgv4oShDJroT3WATkPwWUnp2XMOt9
Aw+GSxCru3Vgy2x1fBNKhq6Nu/oJXe6ppxXLAlumnXIPzMSgVVbe7Q2xMO5zyUArpAD+buqDybIf
Q57G6Kev9GBHydi4BVNYWMFvYbGTDOP+FznsTjiVNCR+Ie7BDziqJXQWl9c8HbNPT6lyI/JTkFvj
TPJjtR6DSmwiPTNlSNVsWvdMu2X30jieCnH2izldaVBhlJCkQdhDRxjWM2x2tnTjcJ4NlE+Z0yFR
0gJBkgxl7AmU1/UArHYhRLBGd/7+16+dAav33R7OYgrwNFkMiIQav5jWdCgjgKH7F2CAh7itrEiE
xCSceucnqs31vHtpy/jKl3Aik/vyuBhAjIcGSRbO+JkjpIf1whzfh0lJMzS05V86H9VngF3wtMQv
O5aSRz6j+frA/kljcVc2/P+w6vZpjJVcWFTBBs7G6JU0/lo53fAo1ptOFGYodsFgj3JFkfyv4AA3
7QolD73WK/m05Vx/r2o0ccodeIyZ519tyvmrFDrBO9xeAcqC1ssWw8WozTGq9+spSDAgNXQPAGNz
nXhiJZFrGGqHDrFntVksQz4KK0LnyADUUtlSpIK/LpP0d/pn6k474AaMO/s3Bi1HAcd2W1+ncfgp
j5NgmFy/Uq2QAs80ZDvIYzv/Jx4CKZhbhdA1mz6mss/UgoglMSJ1mPWIAMh9DvwpLsUrAOKsU6ad
S3ENUDAjTDwrvjJDp6wiS0cUjGTSo1UGBwAmuKf/ybts17N/IfrksA+QmSBucrH6Wuu5HLb+w303
sivbs6kjkfVkuO7mR81hBFKibXxE4zjmLMAH7VTVdhD3BaXhlp7zoZpeUQQw5VhUswXnK97WdB28
3vkToCDVG6L8Zi/Lz9sEynfDbF+032VR4SOZ/3Ymn8BmOZfr+aSksT0fUXr4SRP7nwSNrXmI8aqz
+PtdEzwDNdXR/vzsee98fSYyRhi8PmY0hgSM8d8kC1unuIKlAeOcCQOSYD1lIAMsk49EV+p1lhnE
wymc+FWNK7XBZgyI4TwbjfmN2W8zT84+6ZbMfzBl8PvGy0lRq6mHG83anaiGYJgKWwP+anRid09u
H1kX3NaYJ+BejR5I7E8N2TAibdvxCejNn+SEH4tUwYHhMjN8iMgz4rVIrmqt0JGxIUWCjRVlKfet
22F/bbEHf2RV+c3P9jCLf9aqwt1FBbBhmpPJfZ7/Xp2FhycXTK3Oj0lai3llHdji7bMzPAJmH6Ik
sz9JEoZoQWO7Svt6lWYd4J2EZy0tKeeK50He6yU9KpdmmTccjlO2e5u5R4pA+SpPukqBk/KnLvPd
Ej1M2ZccuDJQG0rQ5gAclgbh0NHb19wuLLZGel1dgYKkZzb+mvnvVvtcn1CXakwSD8jys7RqGOI8
y3qo3Wzp9jzTZIgbH3XFkqxCOSIQOX+bcpfvFkPNjBCVw7BLRcYx3wgwQTA/AtzCpH6UiKITVSpc
LSqUFa+r8nZCAKhyllcF/Vnyn7kFuHX/lI8D0Nos3TMHllT/sk1dDbdbQG0lT1BUJapV5hB81Ay/
bBCd2HEGgOi3i9qN6Kzd+M7NVRCcYSPQLGz7HvWsj1OYYNQtt1nsN+n0vfBC6WJSMtNXT62Js/zv
HT8wz8d0MqQC+F2afydq19lSwi5lRiAvXjqD8+KAP6XKgC2WdNUjSRbxUZPZY1a2JdfPl1NgnoRv
xbYo58IhFouoArxdH8xuUtp1cpCb0HoVwVd4YMCK+QRKpopB2Fs1a6wvvex6jdTeSqbGmBu38s+X
ivKhXrtNTCpHwVEJijl+gwBwXJrA+anWCJjHmAI1d2cYhVZAqyWrB83W2xHqBMtmoJI1Y8u6an/Q
J98hpHADfisZwFSbkCi+oVBVmmCCTi+/1jZjZ3qtFxOOLG2DNhHAElW0/egIpnm69c6xX8+dQhZ8
sheoQrVKTNDEu6qpD/PtDLANZBvnZaATc+WE2EZXUQIPUo3HqQ+jPKy8FTw0u8Tca4ntg1tEneqS
+BM4HqbMEZP6Jvg9pz2+LMY2IjKD74jFMtrPIuC6KpRorVFKCJbq9YUXvGVOX397Rci6UOd2StMh
Q9v7O74WcgJafRUTk+tEwmd7AUobaHdzbbl2XlERTtEt03RlK/Q5PbFlTfEvqmqTZcc91wz4O96F
x1pFfMn0GgacTWURlHwaoqZ7j+2J/ASQz18wfYwgYTQUGp6VVB3SSl5FF78nWtBoH4IuOlctZH33
2me3/8tkpr+BOUWW/cuwEqeeASj4s8zj058Ai6+dYoDDeLvJV9zT0qVABByW8IQmI9OO3GXEVdRM
9mDlY5fcTfXrfdZ0x2oxk2AcDKxNZrXM54gbcyOTgMaCLIQKof06KxMbhp30KD93f9gQbO7j3Mqr
uSzNgUdWhgpAh5Iep5epI+U7ydw99tO/p7K2CXT5O1kvcxmcY1x3KeUVz/z6zDT7ZrNat7txkwjj
UsGXCVuFuGkZhj18I7TKo7mK0W7D56CGNQVj9B8tMQOQi1ArfYVjUr6pydF/qpvlLCDAVnnVE9u2
jz70Xt1lknfjDUGMGQCOyPQrNiO/wgT4VHPHBBoJ9ie7Ijod4bQyhkpRu+sCTgTT80RBCsRIM4ZH
f43FfvZ97LFfS6F0m1EQOO8VOviSJHBom3fFF29V+ym76IFmaMvalL59o+WeVAEz5Od2cobadQNK
FVLEDgIlrDtsamAXjE6zYkBCsx5RRuD6o1EI9BIBq+MkFMU8yAqfshluOwlPkeat2QGOzifImhoh
Hz50ZsUW5UKgRI7cXWvF33HCAzsCZnIftiuevigcpxuPy02IqBoawPlh52BUoCeB2lvicUZY3OIA
BzqQ0uOlG8m+XCTEbZI0NxmrlIpwxekitesJueqUA9Q55qfl30RQklfVNouhNFYl0csZK5Eanykn
nbzCoHDJkXv+s6lNzRV19/KfWSIo0e6+OXRR2dekkTnyGMp0vJXoRRUImG5V2O4xEvawkzaK//IQ
fmoetzIfB71sx+/eslY6tVU/E558zc7yJqci0H6WdfiYcXJ+HVPM5vZgxM7KmWL8I0VkI69CupqA
znaf8TffmkxG/+RMn9F2xbZ88mjDEBf/96bsTQp818Gb+vxtB2769nH/hLYZ0/FjrQoR94JhnVHZ
AUvJa7tS1fMlVhg6M/z6xsQGZacHxjeMvQLrkruvFMUL4g900WrmOUeyIMXD6qJwkycR6uuxCUFJ
3Lgp7/wOuXT+AabV1B5KOzRqPBpxt5jk4GcgjNLR5A8s2g+ra59lFF7r5YZ6j0k0uEc39OKvR7Cl
d0EYuXf1nyH0paL+YBuOJ+B36Bl9YnG5tino5T8ShjyzGoiEmTLnZQLqLvaVl9QaOAwrW2Q1J8go
2v2sHUUbr14WW9Uwf8baK9R/kGBBPYz0FymqbQ2bO5g9urrzwOG26tBImzOvgDeGN+ADWd2o0DEx
E8GivUdXawmixVqKaofrqO3bt8mIHs/kxyOmXsoZfYySVXvDLnTlTxlYBnJYRfLmLxhTRYAbVrvW
EWNtovKjGnYyqYPMz+0wGu4iDJZEmNVGrmh63VaepurIKvrCb7TLhj6zvl6h2PG6df65xTT+8jxF
5UnqNtovbuslGI4uHs+AyaqtG9mYwyvof1ZtVp91b6ew1J3pH2hKbrGo8cax7p3HPtYLGn++WJCW
eqFyAKs8n1/D+8+Ecc7CpXPLhSlHAE3IqCCPjTko6ncim0/GWpVMkbXF+vif5Swhl3MBjZ2BoRQm
jUoNHd9hm3y56/ajS50abTLFovHwCsG6oKi17yKAR+gcnfl0OEqxf7tne8mzwEzqrUje+cuXyse6
Xm5R5m+5NRLUmD51hO8V9FMlu9Fp9ZB9KnB7mpNX81sMPgksNB4PNQOP6FhFIlxuR08+16bvT9Wv
3D80bmcax7WQw8UvSAwlBBMkU6OoVufATBmQLNgECZRV2lSCb1XISIksCJ4UhvorR+scnLNpZzrD
es6kxHgFXWMeS3LQG0phNdG1S6EYS5SgqUkZEZm1a9ydgxGauHv7IrM2EMe41Bg5/MKFnBCp1Y5B
FWJ2X9J08eOir5xDvd4ePY/6Z3kkgd7zVYcxFEoyC5IbHmtTBNbpd4ddhkrdAUzhonAIct6zbcXi
pzCzGWk/MyVatycwEJHVUAM23kyI0bUf9WhgrIXQ8TbRbXIsOkXtk83QHeF3dzfOxlXCaC5O02/v
HCcCNMXNu57SuP/j+otCDJHgGRh/yR0t3Ay3D3dEbs2dgR9pbdzW5hdS2UPytjYaZtUBYxMtnUpJ
LgD9J8ToXkl65IXMvYVeHV43KD37qgZNKbB9ibmjQS0pM7uCgaa5HZa7l3Cbl2NvMA1TNQPdxcXZ
OY80d6VciYa6e8znqioQhJ7Be3CkTzE6yUivRNj9cIeN/KA9FM9c2Xhoc0rURm9ylsHJ4XShCN8F
slA0/cSWHaZ67d1YAOvJ9nQChWb/5f4OoaUDeY/h42Iz5wELeptxMYyw4vYMLsai0vZuKJNqV67B
QZouqFL5ygFHTVuNYe/kOQwbz+78HexFdTJxCojeZ2TTfVkODhGoSeS7LIncYRahuflDC6EVfSS8
pp5HuaLOFzMJxLRwSXXkgECLnQV8i4X797RPXkrX125F2czuJLtWfjmBdFg90baNUV49NzuSWrqE
F9sg9LaymjtFUKTEBNVj7K6LCpRWneRZsJcUuZPhevJeDlrhx8xR+4SW4wTdS276pb3XllU12DNb
712g3oSgfhJwwuEbdt7BmeAv8i99jg/damJazPLkcYRAyCHNNpFdq+YTzUHg1KoHmWeMsCG0MXEd
x5dnMcsNgQUw3SkoaUVXNr4/W9JUODQGkwNbXHaF3JMPCWNiW71SjfXqCHx2Jxa7ZsM8/BwP36E5
CXZcveZEZtC/b1iILsmvrHkfVeDfaP5nT3tJqR4bbwAnwl0ikR67Qsh7D9F2MbiKeg9kd9drTnUt
k1d2adfQLVHRJI/+MzoeyePWfCjMUeJlBjhqBq/thiQUasUcI46a6t3eyjceQQj5fo8/n6E3MJGl
Qf+8so1PUEOfv6aQOvpCafulkGi73usfxTfY/itWv3R8PKtfr08c4ygsTa6v8KogIHaLCZvfIJdp
LlwXeWOkQGUA4QcZNXFm1Io8XLDIGt6HCpJWpzBrZr0QDHPsTgG9VE4+Vzx/4AQ56WbMLFSU7jlA
JSEqJOYOyj5nBuQjuLcgRkHlD3wqpQAcX2WXbQI97M6lmw3ddMdX622pBCEdsuvD9NaECvMakhud
qaznHCrwPnVSfy3O3X8oFx9TvCunnlXCSkOS4o1bmjW5/KLPXjjL86cuBdKu1448UUnBZtMOmbNd
+H09dfrQkOirJOLL6bzZOf26utJ4rAaudDj845uLDi8dHI2jZcuAENjYS8C8Vi7Sgb6XzJYO4e4g
Y/5r4yZZNl7dBv8edRwxKlA6W8cGKH6zgwielgrhJRstwFpz9MHlQqiBuPRI+Da3drL+Jwg6p3DH
4KBVVoHleddKk47PUBKIkxPFTeaovo2Tni4ouWJJxfNB44TEDjOzRGlH7WLN+TCPiTm6Zqn5OHZE
SM/ajx67ziNwcNQW6vSGAmCLfzecqe8bUVOq8yTgTdOd3YyKlU2DAb3kTGtrRo9lEwmPNQiINYPG
cEKFYr8XQtUU3AfrGTCFR+NcrnQ8k7WDHl9uB9utQEcd8vkk+6huRMXq+dT9FqKIcJgW2JXVdamD
/zCcxwEQlRgoZkGa4fXBAHkCR/4XKgqj15cN3kFG7TkOQ7k1n1SKkLWs74MzILDfGEFvBo6q0V+g
hBToUDSDQQJ7qppejb6by7MdqGf/+UhekmyBbwT2UJQMx9Bnow5kHOFF8xFZh2mxiIwkrI4YVWbp
8XJtIvw3lQYnUuXUPCkLIAt9mnWVbXlr2WO83ha2wF9Q0DviPESmika7OsM84H2qXyh/JemxHugI
aejWJ6dtSzxS8rjVueRmN66i3zvkXwd/G7yjJhFrKabVMKaFH8KFIhlO1AL3D7SwnYx/ll6h3mlQ
QPw3JZ/F7rhiy3aGLJ+9QmI10GFU/S3kOxRUXvFdqUmB0zRIXLOHIriJkMn7qhJNAWBZxPtvA7v5
eRsCNwCzT5wOiIeSIr5pd0gY0riOF/QdZEczrVDmu60FvgsEhgBYFqQxB35nfGxLlakyFjMvil6g
IzUJIQPxhtJT7910ytLPxz03TlfEhmvz2N+TkaTmZuHRJKgyRcpkQXtoEELOXULMMrDHjacby05m
eUb9WOKUbpyuv/zpNtd4QOb6ymvPA1z48wrIkhuAmrIC/eDntG7iDILQTAa8ji5C5zD9e7g4fQ7G
IsfL0xTcr2/6X+6Dzi6hPsmAxeYHCI9um36WcyQPyAwq3aPYlmRIYvM7fsxyGzQOnSUJAwkoSpRg
i606cB3Eqo5pcNtXp4pH4RMFZRSqMrl8nPTqOsdC0G4ZE9ifjaQG7droIT9NZTWzrHqAg4nJk+kG
V7mWWvq6ZUW9S3oNIMBwffNBLqzlgsc/mCr7lJn/sipaUTR6EL0MNKvALiwO70u21qsFV5IVp2ao
Lel1yBhboaPM3FLAotWv0YJa37/ENEGatnVETtq3fREqS4V0uP6XGDBysqXDdBoDJBGCEuJTM23g
9cOspqvraRBQx8ISxevEqXVcvtzBs8JFodtYhM+wn19MCsyUB4R/Sy6+SU4UYjmmUJ446gk3Kjc5
JTrGYBhKO9r+k5XwOompAhENtG8tuVYeKIHxfO1vFLgq8SySvRFTqoyGDL9UDzP70jueybgHWK6C
jp+5pjkT/+ZoGq7P8PTmSHTdzYcJLCH2ptLYh7w87J2lJevwk11OF5MLIEGh/GKesMaL/JnzX1Sl
NJOVSBhi2ev7ZdqQIAI0hZrqopHSAV0fOJ4fx4lhvJ3UmA2JUVzz9qX8OgQCN6FOLrLiFmxvyKcS
q1SMNsSU5ImsD5/iZ/mEv/S68lxO/JsixLqqXt/49jP0r+BAa0CmtRAS39jp2vJPhpbmnLMscq8a
K7Z7EJnU6ksZWIcxUC8OhQuvHl1KVC68LKt8czkIHua+OdSnSufvO3Nu0f4gqnP0zv9TpXCH1cXv
QrHploW/PYClaG9nQG96936dX2yBFGTAGy3PagYOU2RHgdNnqdfD1YwMZV1d7bkr2HXONJNivMkq
hU0sjQ3ErKAs9MSBNPTX2GYbsROnk9llltw0hLfYx2gFjiLumLPQf6C443jtvR4fyhcY/uWu4sbZ
y1j/pvgBucjCIMd3Cxnncds1gSWweSGUG6/hvhv+eEDtC6NIJJqVrGos8U/4pQ5BoeSgUMnL1vL3
nkPGjwfBd8r5yAZbFU9/6uiC9JAwb2A+hAhU7qLJIF6etq4wDx1fZxLZH4Sqb3OalJJnMTFhVTtk
D4iC0IT9Iz7mQMfsxzSDBge6FpKbM4S4PmpOY3ohwT05TwybEyiqqxP6iQSLitiqQN+90X0mXWio
WeaTePhuSWN2vFjbD6QW4vR+WDyN7w0GiuQo1KF8P0vgHknBDzWeujA8K5AOjaRIW0RczHUZmtIe
BsZcux76CQROMYOt53s4nKvE6dfPFzSrCKVtW3pKptDpHo6plqVa1FuP+hC+pvyn8Z2BfvLQO5zW
AswHM2oHrQYkT5oW27gs8NpUxXZG97bdgIeqAPMUbEnyqtNJrWxC8whL7bsAEBzDjUQ/47nwCoUe
SrlSVOnI4aFqGcvxKgEsB/2BQNsuS2g5xu68RU6uWoLLPMp4XQzJFMQdBQ8Fh8MPcELWTzRnCUy4
M58L66mkMPR4vOc+PE1wOR9duBrC1oFZdhX3DiNf2xfSNH8NtPu+CdrHDIdEDkwDxzGqNjq8BE75
oyxgR3C2mxEzQL0NSz5NqYfFfrc09G/uICOv7/zc3gFdiusSZLdg6pMNZGe91S55Vf/JFulxdenc
ak6S1iVNvVwGFYk4O1e+qVjbBGN/orERf+NZlydRhXabv0UizOuJMsZBRz4SQUKC20ALECF8w8c6
aGXFwIDRB81Ao8Dp4Ym2yWN44NpFeI5TD8mZl6DRjiZWDWYPolFwv/5p0dT2spcGE7iOCHWJrXlc
nnbUVvaiaf4udp4r+NDbu6uJec2KGZkTYv26WFDvU0nrfMBkgJEDc9kXbHYCHevsbsdWbWQ4FCmd
C1LSRlVn50o1PDrKLTXIxhyG+EftPwGyoklCpD7iG49ju7iAZOBFoR44NT82jHWioQQqrLafesqc
j3w9LWhLz8/vntVtLFScQk72PJvh7cN3hab7JDGm0CpYOH4GPm4rPc2CRdP94i8qVlQqTohizfCI
2p0mJLw2BA+7XrD1LB/4rDplkRe2+UZUUek2T9Sce+G3UAGFajkPTL909uk2yqLEdnQ6Df4Vn8ej
UJGwb1afSqL4Yls5dTVFdswuJUAMEgxTy2CQMKuCQoVCLjiFyEjdhfCF9UbUVjGw4cMyaXwenn3M
ubdf/nGp2W9Qt1BHkcVPMlhxUJmTWlL/15QusUYHUvqM+tn3K2UDAG/2efLlWxLoYR/yAtKSui35
TK1uujwLgJwy+2ZMS35zvidP0nOjTvTKEiWziOCucRb792EhEN4Jcamrs+UuMbVEgevGoS+rEZCm
KKTdWfgcoJdW0bKayewkuwZL0BKoRoyNGM+FP231K2VtRBgatn4QmY9HTVs1TAR1sZrG+kagxNzL
EACJfSGFHnBDZnQ3vEQ7XzggjiR0AK43LWOj7Q40XdJ60F3m8mP8bJ09Uk4DWzezHvOz25V/jkO0
NWEsCgTT34/vURGXNyoKmPubEi7qI5WgfdNnkHen7mJ5axBdJQ/z9oMt6o7XAPC/arVxIuFmGlUr
uBNnQBb4SdMV1Tcv16NzjNeyMYLE6LA56vp1cfPXrnzR7KiYg946velppmt6VWZz6Ie/vheLdi5Q
um4xU0xKNrUHfFcEl6OWtmQayQqnG7Bwbc9HQYq2sj7XXVZgM2rpuq2kEGVSBhORTqUGfU96PN0N
50eZlmDigeHALai/MUULdiUTKk8+Pcl4+YJP4ByL6b3aIcqFOBDtCEqTMoSYB3Qpe5pGWzwhVy1V
uCQ6e2+k9gbtwdJ8y6I4Days3+yWqqv6sgH22FKC3O4e3qq/RERp2CAF1dvElcbVDCnslDZ3bUAC
ExpElZP1bbIjC5M0BgpgF8oHA8d4WFN0Ujh9Vjtoj/Cbr+DwtZfBC70Rrn9VirKYrXPKB0Kd72Gs
wOdD+MwPF6O4Jhy+KFNJE5pSNGoILvEDnbdgshlKn6LqiYHj01AVEst8GEqW39W6isrpXVG240kM
GDJGPlMAeiG9xzyY9eMd9SsUwohJFzu6VWjrLSstjwvKawU7TOnNyNR9j47Ggg3WfvyzsNLrGI8Y
/I6NuDWrWAvSF+niSOheovXY6f2eG/KQmEZmZSgn1O7ywSVb5IHWpq5x+iHh8ROCDw8igKVfxUJv
MaUW0ww2GXO8PiZOqQp4Y024Re3gq4S90rG943az+BXB+cn1Tvck6V9q0VTSQ7rQDFlJAeICyeQj
IEB0I0a1Ry2g6hoDx5BLy1VT9OcbhW4+2pH6k73a+9FabJPDD+7GJLo7P3mgJdtJEtMIyb60/lFi
/nCbE4BmT6BDncLQFX+9jMdNFdl2IQkkivCwZ+LaNvJH77mCwLeveSLPkDkb9BrfsRXpQIyeYIhu
lTW+yCWNWWGy0RqQi2At4Aym6rYnbESJWXdozbZAOfnNDNY4HDNX7RQt5U+2Akt3wwaTt8I4O1t0
9Gz05ZJSYK77ZdmD1vq+8GWKyG4SA/Hx+V5DKbqbE/VWhriUD6z+NiPvRFrSYVNIgWVlFno2c81S
cI0okZbsCaYnAnJZg4OBBUPc5lopsWPzwCRl9lvjrAHg+z3B0iOhqXQQwu3mXdWXg5HvvgeVjO0Q
a1ffxHWOm3kctjzgTsztSlJQoqcA3wwL9+clDhZFQVyjg6pEEf/Yz12SBo4M7SpSI7/XtfCQEPtL
/IEtNjs1QRp39rASM8s7x0OCUwmpMwNPsBL+DI0h7dGOx/drOtIRhOcSfhh9fXd0YTFra/uAUUkY
ECS8Nos24L6+2hZna8LIjm6rj5yZzTmMx4hmdxHSnTpGSmBghRPixMs5fX3NDg+JzEEXeEDjZVyN
pltk/MQB6t0CW0414fUOGtgvQLGVf7MUROHhQXKC6MsfnYAPle8rNW1uPnQbvkzK9+reMzutdREN
MqKuxgubpKhBVZDRy3rWK2FNeQ9W9uMLms1O9+TFAzWmQWDnumGiNEqamZOeyMLKTjAVY4GqJpyC
LPCX7uiwCD8f01ZLbVXbrZVOzuFePnn2umeKXQbXjnHMZwqw9ahyYm96LgtfYCTXagMJDyIZPZcJ
UtZlGTSCm4fyOZBZgnWKz6/Gmo4BigeuFHp5ERkTdh3Cjqm2NfoMRhhn0dIyrxrc0VQhKHRfLL75
AQR3WUV26jN/rlx6qm4ou2Uee1n2AklFRy9gw5atH6/U0qftDxnSkU/fnAzVDIIqfTgBpyNi4V50
y7GhblpphnIVggCt9av/s69cPUp8AO/s32raCV5QRTDb2vskmXGA0I9YgR1RC5lbrVK6Nf5XzNs0
22syuwni0ZJlKFwJddWyKX4oHAtQ6xiwWLrUKV/JYSvqOVIXwOLUIUuUHDsDmuoohC4oOX2kUzO1
Hz2lJ2fKDV0aEDQGE7CObqkQ0qdr2nsPwRyOYeoijIYirnc6sU+N/19vc2x+H7PKdHcL2mSsa02O
hrZesNGWMI1f6a0znZm/t8+C1YAOOvfeDfRUz7vBGVrVRApHbkv8ELoDQPdwe+M9dGiv06PrVrUT
wkQayCk51B6SGXK/lfXFqye+MZO06RQfEm0CNCUhe5IFpnpQTM4gkB+cAsqJabVBnL/lBF+P4DMB
wwpXLMdcH//8Ra1Sjm6gJyLWvt7+pHW/AOLo5bGGG+q+90e/MQANxuN3aVJ1kv4A7/CGKi4Un+OD
ex2gE1aPww8JTf3mqJJlJan01LesdKN1rvPxH2q4COo/T9gwbReGfF9nZtFKBHWvqRLbob4JomCF
j3NDEi7pPs3pY50XSsRPbYSyE+VIjbMKtYYzLpCFVxNufJF9xkVc5096Dbgj8WEaRnLKCqyVOYqX
thIKlTHh79gSqai+07TAsD71z1ieQjWvN2m5UnuYWu+41gH47EXcgVmIKLj2OM2NKSE8rF6iYz8Z
uqARco+uFkEZAZhGtAtlWVar7KXaDFjPNMF0uztRiJexO3+igc/zqDPmGpYdKfR+YHH9FXXXigq4
YHMjNZDkrxCEpZ83vULxrQWK78PMYks79Z0BvehBwBYzc09AJMnZt4Ry0jiLlFlhE/VFV0ubstnC
gLF+uBR2Ae0IBJSD6H/Ypo6UEnluRkIwSlzLV5zkAF3L70kb9+q6ct1RlQJczjLnxTQIhyXmj7hx
cPBp0ssYN9xMh6mTiU0WEXPLTAMGpeX7y6JX5j7+4ByNvwbWzqB77qYxiIgz0RWpeKhGXeMT2sfr
rTb5l4m0llyfeu7vnEvOe+ZgaHzj5nTOkDtefr7eLU+0hFbCJW3Xpbzvs2M9AjTN+huxuE01Czjq
LVxxzx0/3DWZLADyMXIFqHvo/KJ58dsWa4m/jEAOFqsm7qm5Vi4nAl4/oZVdJxPvC4kJJ125LXNt
Wl5j7NOW2a9ol5JBCuQToMIGhQ7+XBGf+gprFMNwut+05Ahk6kkpczg8DRyeupyItjXTw3KSqYMO
LZcaS+qeh/bmbT1VjmRZlQUtRIP5noOdd1lb+J1RWU31ttKKYEMpoJusMIXx8Iq1iG88HvVPTV/s
LkFmaHRlvmxZSv3oJT5UqEZHdUJWYigwxNiUoZ/mItOSCmnRoHZutHWlxzkBqw/t3Bbyg+Rk0qz1
fPrKcp5AQ047W0Zd0/Y/nrHg4GJM1+Lz55zt2QP9KS3zMrsztPnES8dxhdQEUEeOSRJxcCB0JZ+w
NI1cX4MDQ2+RpDsLFOf6ylK80zBOTFPwhlrizDwwLXZ0mBc4LHXbZ/SDHmjXj0s1IFoA+r861T50
xtwwG9dNSKe3bnLtVa8c+06UFS6ybtLhBIhtkfX7iKCmv43sOvcJiqJ7+5LRYlOporfiXjGQjS/b
fjMSTyaPLesqa+19u9HbeEsPsCvQ4BTu8GPOSpqb5HN95fvOMbPgD7sNuKCTOUZY1uRbeQVW+qfm
nucpdvjNRK5FVNP3FPQbm3X3nHHZua3uhup4FkWs7Hkd3NAXZOVl10rwYkMOs2GGw9eIZYzV9t/Q
IvXHaT1bSVvdOmd4Gg37IrkPMlcxH8NWxrFCGSxNLkVapLDQD3msc6saRKrYxXkHynDKUtUurKx6
XWYZDb/GfSdiatUSNLhl9IIgHJUohXqJBLv0gHdttl0tTzGk1iTrGHCh5tpZ0GDhmI0f8+nDETFh
a+fyQSB4GB+6FqrIQmXX+1xdKNrDeJtuLGaX1hr/omtQYXlSM/m9m4SfVncUMFL5G1dudsGIRvAC
pSCpS1I9foSfYnynBNKSsepBz9FHCSABEBEJfat618roI9gsOO3F6semhIZZd7mtuSTdeLCWQd2Q
WqwoBmf4LdipJ2BO6cfs8hD1s3e5H0q3QHxMa30gCS2cFJloaB2elnxy4ivfwGh00IvexvgAsue8
NFYnwkxFq3LN88ZCTjei7N3lY5nShv1LlGXzE3i3+7tlUXge7yZQBgSWRffu7cvIyJQPIR/dvogj
PoYV6VRdEJpRBywXtL19AieHO5O+ENdLAc1yVFvDmeBsO+VpTMchAP7hwlLIqDw6CxhsPwqn36hy
+tvvL8gKQck3Xivn7RB+nHwGFruDdynJBE7ay9Q/i15TI82VJZ58ZdAp72hRi2UhFImcunzfmYqm
yIJknyXPxSpOftjYUs9S5oSjr4p2f2MTIkI6FHfVLDnzGgiGP60hSIcQBvg/B0yQkXpgR61cjfUC
uDRYZnf1GzGXLkGD2dDIvz6QbEXyuv5+lYtHbBbzDQD1jP/yjgMuPek9VKnZeXHPk6WPwTQkdv/t
r3EM1KghQxAtv+oL9qc6B5KuRzbk53XmzPhjUxLLoWgN9biXBgz96GYFaHIZ/u/mcx56QHghc4mf
5Yn0oPsbjsjrvALp1bGE2lzoufw1phsE2EQIdSonO89SixG9as7u4E/W8ETPs84M/0Co/1qRvs4Z
2/j3+lhigGzAFN9UtfXSuQD/2OMnTjiusRQsy8IuUECAbPUcctecptfHzESHk0wHlIBJZsKWf57p
mjHjQCWkF9mYhRDohS04NSiTph4UaqBh5jzZPOifoHn0crB+pnlUaOdzrb3Fqi3HcPx/mcxm45OS
QjgRkTC+4jOxTe675KVczK3ryPLswhTKpOGfPCt2qQKiOIWIu5UHFlAd9B5vKHuCtfrrgvNS7l4N
VpGTjZJ5qD9WLpqj3as0V326GCW4cP6sZ5Z8+Rv0UYnkKfVQD6Z1ll4f/Da+p7YwSHElvbOE66kA
vbxomAwVvQ2hEDSjYW71Dx7K9uXnilcnHN7Z14mWff//1DqEsot56sJrR4an5xIyjadjs6Sljob+
/mRjmXL/P8iW/IjkQqyu8M70HMEGtI7ODyPrFbxuRGSQaDH+KIGTJ95AWEeOTJUkIrPCVZUzQpvp
xL0ce9+WLHS7Uh+Zke6XRqwdrMfl5iUYXOOYw8ta0GbiTxoVaz7ZhQoBNkVpxZXzgV2ukhFBa09c
yLf/XXaiaZK3alAmhW6sr3AmxroHN6EbTcm+tXK30IA5pOwNLPdHROoYTHqQFXlKZTQ1MykCpTQR
Luvr61+WAZdE3r8q6htSL5RF9ncqB1SU0j+4GacjC+bVA5crM2cBLdI9urYoTvDN+f9FhVXVd90R
PaJ6K/yodlyio5/wFHKWJdX+T5fWjVT6/1HZLEDurQaSAqMt7bS6oWQnKrO0cjSD6eqTSksh1gbQ
+gTfIR+P5mO77+u9fygUnhh9W6YO2dFk1YPVT0GXDU0FLX7ONp3ruV1W1DnwJeweuBizSa9UtirW
giiGPAU0nhQPW2o9kOAzffxGCzcE2RN/hMRMy9H/kJ6FXLqsxHC6TBoGqs4e/wX0p29+iHnWJjrw
+SvolcedFXVYgGrEu9cG5VXbHhwmnYLsaSi9UKd9dwr9XD09Vd/b/yzhawzjbyClsdk0y+RFpLJZ
9r9IW/wwFBKK4cPn6GKs6qjcwE66LHJyeoikCNi2jSUuMh94l6WWK0svSNvWGTDNMjNGMWZpw098
CEc6rtDp/bL+1A2dr1qswTMJD4ae5f/pmzt/qwVKt9tGExT/6sqX0bO0DPD7LTypDVrKoUZfaT6A
pG4PDjwKC8GA+MAtcpGL8AJLz8pYvNfyEoefWxxI1cs1+XH4Nv9QDtvy0C6yTDtLq58Vf3xt4jS2
8pdoErB9AqOBq7LUJSQfnbZjVrr2D0kO2rvGVo0KTLWbjJi/qn7VFUxLt5IVNGLwHP+mqxOMnt4s
M5hCjKC+Ca01qAKfRGXLKY2oy03JlobkclaaHSVZIveXatrIG4lVtnc8zPQR32ZTIgfRbriZLCft
pEhDnFFGpiApqeoYgHpTPaFkBgefGtLpcUeH5ChtJGUXCcdCu228NA7l/Mfufz9xFu6+pBykQie1
Ct1iL6R29e10WFhYMy0hTOO/nePId1xfQYrgkiiUumaYxC8Jlmv9FOKbc9cv30DH1DkRDA9vKRFt
Ef3nRAmm3gJ2G7G/ujUapT2lmfC7spsm1xz3mkBhIKipxIrfNE4pCf88Tv5ZWzgJBVY+qCKvKJPe
BmwpiuS0+h9cjM2ot/yUZ7xAHHThtkY/i1KeG4LCrnfIYw1mQnts+dSfqQfaOKJQStikmwJdQ899
xE9c7YYSkZ6BbnAgFTQ6PfSYBbn4ra2JxVmT4lkLX4Ik9ntvCaF9jPvsb6XU+ldJtRpJ6sRIvMpa
Mjf65LKgSsptw+ls4uw5d6L+8FxRhocoO+LN/64q1YTfP53hPqcQqk2UtWgf0ecMIu8JVpmshh/1
+BXO+2v7vBql641oDkkMdv/YzarE73txIBpSMCETJMQpR4v/fZuLLinwG88ajBZs36K4jN2aj+qZ
pafRrUZnVZ9mRptoIJCBRD5CbyvA6jWMJA4XapXy+qIVaAJhkuJeoa/7NYLWcJH44Z4X1PfKFMGI
zTdJlFpN8Un0XQ0nSvFOnlBgpQOWlKQxsoN6HelmrXv8tZmfZyvDL2T/Ps5EIrGcheJK7ZFUgF6B
zulzSSVBN+GYl7gq4ZZbbpUmrDEvx5/ZUaoU1WGKWXGhuIQk4MQ6gtSYDs+ruDRtuWMbAs22hnpQ
YqMXxbBZTYvY4U2I8tSiTKNmwxxSNyZU+qyM2rcmEBM8jt1joeejp68Yt2siIlbrP2aHZiehDLeT
6AuEjEjpwI8zPc/Q5CAQJucjavOhfiyA5VeiNfSAJK9bn55vmTNPAiEx6x3wnFRTk0yO104hS+fk
haM+O9f6M+iHtdrPCyB1RzHzR9phGdIN8zdMy17TdCexTb/rZwkkiENeS+F4oP19ruEAWJOkQdV9
D1oWKT7b3Td1XdVL/vB7PI5vyrYjNKf/nVK2hyW9+SFaw8GKcTRCPWmHwLDM2jplsV53bP+xTN7I
1RJqvnzaIeraUTpKpCTw13EzogLx9/70qMxsl+HZjG2tU7FMUILgeaRoOT/f7SOoA3zejYPYpE/l
NbleQWEF9NtsXlpsSefk/W0EeitGmX3TxFuc6btMGcOmCxY5BoaiBl6HKJDxAoSbWWIf5rFo5Iim
/6etwKflP+NzAPtwdZM+Qu+WPsTa/xQKzop+vHIqULY5g50jneegTiv4LiuAMmZTwUH0o8jpAkC6
Egk+o0vLjP1h9JG108jfioWMNtmg8LgBijoczcNylX82kNY4DAEwPPGLVQzj2hCJudddiUOEDvE7
88FFztTIh5zqk7O4N4C26S2AuZ7IkFulbNwX1kht5V0dhD3XS51YGsK0azcR85Z0F8nufrSb9Ot/
uDxujTRwe6axEXQqwP2kG9ATDVehJ+A4nFmuy9nfAcHuX7efW9Yaoa9OvxTxu/b+2VlX/21ib6rc
7a9zwoBtTyqVuGk4YyOJEiHtWlHp2ARHbjbU4qKf/7wrp34g2912i1GEQ07NvBlC8kg+EaLWheT/
JBZ3v/QcNeQkLRf6gP5tUoWe7yWkvX14TUa3rf+HtkYb0ORp3sL4AHpJm28ZIR5EVt57lZSSpXra
kekRzLH5gIomK9O6m2DI0fYpJXyGUzLNhLeIc/fQfYmVNbv1Zb1aEHdxCrt5iTyroOcIuWtHDIgV
8iVH88rPJhjODv9h/t1WqJjKPyk+b4oCDGOyDdJO85lZ3hwPHU5BUw8HbrToHJTOfwZ4RGfpUyho
Smih5eegqUsfCqb1GlwIkfHskUSiG4qJC99k3U0fNYPfpIB/ewovLzcIx7qv1VcT5bqykrp0h8hH
5QcBsEU4aYgVil0GiEQpYnRXEdYCdakc2WLPEmDsKw2rlNI195Dvf3Jpf7u1jYn8k6UXFUbam+NR
omeUSCtMXovnYW6KEFhOt4/FbdmYZ4MIK85Boxj2DshHUH//jLSABVOBcVaNReeMJBsyYFbRVOs2
J91cWe/zoh8DnHSIB55Ge+nZl4lszreOsjY3CnzrtotLaZI6mhgFl+PUknQYxWJO3Rg01bZff0AC
+RXQQmPcby0yWxyhSD+JshxI+8Aix5SmnaLOyFr4GvECUPn7qCVVd0kZcaRVcQDGk1mVJD0jEwNi
jvmGOhGSv121exqHCtrKlx+4+oBl1p2G6cc8G2OYMTU1Yt6syJ7DclIo7VWX94WF2NV0ffcFbc7t
vtai+gbIvgtzW1n3Gyi2E1L2YkmQyF8BCK+hm8CnOufPS0aAYGSW/ezz6k6mg0LYk/X8J+x3PktO
gKGbPv5YqgiHPeVwVJqzsjqLfJ2Zp5xRc/e83M2WtMg8qY8c8yMsHNmqZCn1MtWjeFzyh+IE3rOu
jJiV/WEBJd0tc6JRljOYPvILBFpGgXmIDGjR8NRFMdC9nm4BejF5/FoI2Qzb4pKqo9ZKvWs9W73B
9Ww8SQYxXlFNDYjiJJJtaHhKP9OxWDdLf8ijfN/sfl/vzK49v7chZXz40m9R5kpQxtjS8KI+FKgi
R/c+8o51b3x4WUbuu1BedTLEZW2AiiXGHDHcigO6M8SDQHyeg5Q0/eF2GmgN2GPxEoiyrwQLKaoV
bu8wrLuaQU1HakXq3uMWlzQsoR+fVP0a2JWErT3L59Edex6SBIH+m/EcHaTNROICFOtFg9kmA2n2
sMr74HzFgW5UGWw3dOUne8I4fcD/AP/p5PhZ8tNXrO/vHsHdFyDe4kC7soMexU+BxY+27bMYRf9x
CYmkHXyhvAukVe4ngg2rD0jQooZA9vv5WjWrm00Y8/atlSiLudGlPu9L51Rl/WD+OCfc1vP+8SDz
ga8lUYYhYQXHMxwBjFQw4M8w8s4qUlltzlsRjUz6uSjRB/PnPDJI0DuJxAThGLx4qcgb3ci+qj8d
xU0r4bcMO8E450WbkCnOBAdWFYyZs26pU9Q/xRipfDswUO2V7R31JfJf90Df5ArtIf89qxtI8Mqf
umHZoQdzCuJcNz0JCPtRchfm8qXrdZFAAvaIe4CIyfVFetOSjeq0sVS75XmqggaNOosw+tC2dKrR
2xSoAw1tvJLcO1BA0qpqw6rboUTXj1uUY/uo+P0QngR+iFWC220n5IKyoaY0+1nSDQemXNyM9uVC
oUeqjrntfFIbJKb5WYgp8cyOggEP8Wo9QWqOPETvdphp60mAzLb0zACtf2shcS4SZTOWguYfv20K
v6M1gHGNDNsmY2AcXzsqs7WHR9vkBwzSy2+p/Eiqc8nkv0wcgHhFEGjKVwct40Dil/4FGC04Y6OU
60VbEKH+8LnZt6PFtn13vfuo0qtVVb8shLYgkMTkh7MHuPzkBrvkUOGts4N5ErQGnFMp8GywWQ2o
YHF6MccOh1TUHIIyR6NY1iZ654Eo0zQ6YsUqcSCpg/SfcMKs8Djrdf0OJ/BFgg5c4wY5/ANpa86g
fr1gnEhLq8FvtaGZaOvt+70DUfpLkN+GRFOqpHNPKOFG9u2yNDC5yb/lHh8t1xCiYGWu0gObQJcc
66zEVfNcgeAt0OAtDlIUTnpI5P90TQEWqRMUFrBzDgr88SxGNdT64OfYrVQ3/tnJlmrOWETmn2XI
t3ptDz+EON6pbEdcmJ4aW9dX7t2oJmoL4rwHQdqggY4xYv/0UYvesCGUovqiE+8mB7Lw9TdQBWp2
2oD2xySggKZN2nMB/N5Jz6A4eDDPfGQ9HLCyZ1pfumHfnpVwNgCktMp1kXixgHh6iY+DM/Rd7gSk
N/ckv5NpnNB4LdIv4ZuxS/02jhtPk+BJcO2rIYGLCkoefrwGeVYYOLOElloJ/fdlkJgb/m90+sa6
5WRHaRA1CCVS5EBK+PRaBIpjI7pozY0IQrc30JZC47w30uS3X7lgB7VM7hxtitrcIfItrzaUyH5Q
Q2teOwLko7XoLxjyYMY21X+juTkr6tEboNEJl7uJ2aS0jBX7SZVHIRkJfetSiK4wKqP6ZJPD+Set
bHOpGidaWxLvRHHpH07Hshzh5WY3DLIuQmzuTbTgZM7Wjc6SOB7qvuWqGZEt/nSQHlL5VF1X4Ofj
o1bV2HNT2YPe7lVgLiDJ9BvtF8c7mAlC85UooaksaZwI8RoUNu9T9MGE6xYCkhqZluWSq4Ef7Uh2
P92PSUOd/SKL2qwJ0ZhiXgfwcPL8aMJkQUgBE3aHomlDs+UH6VEln5vuRL+hbD+wGOvuREeX003b
EHl+IsYNcK7TRF+diQLIYirO1KBqIBAuAtE3ikFjChp39L1+y7I8Kt3zAfTNcGzczXi0b79P5c4h
/yAGEcYHw6emCoWhVPDL+jT1YZ6knhsSTex7xM+A14qx011Nx3rtgE+zpz606DPwcJi3weOeZPym
cboJ0xhuHWYvHLGJqDOe1D1BV4W+ji6Pc6fEsOoelXPDFbO7XzOT0Py8GC58D96c6WPzofYy0IlD
D86/RXXYc1gIfY88roLoflgQhF2puL8F3mJgD1aTNZnxXBeuhnQWIswPFyNeBT69VyvN7RplZM9j
ZfcL+MqiE45230CzknuPTx+bt+xj1dFDnKDwqkbEkm+1dQMS93nSE+zT79ViezmVz+ZQr2m4ATNr
+Gno8i9nAgSzVrZtWrRlFbdiE6M+1cBKklqSmjlYt5ky4Sw/0cf+eGVil2HB5Mt8nGh6B7AQSjzV
Rb7SV7/Gjpl2cdpZ1OxUNGe2UU7SArYfbOE21xYN2ejgl1y4K7v10LLxFdKHBnTug0unxbYch9r3
o4mfwgj3AhDOhhtK++qAbD5BtDAT2A/0ObbMQ8fvBXsRzAwNnutXIZdwgPRUSBdOvR6UlrsR8QWe
OXeKYg9KmNzSWP7cd7axLuHbVvsoD8D+WPuXOJ1MxjZK3RYk+YQdND2Yh6Z2/L2UNm5sspmZivAm
FdCxEMds7Wvtua2ooiBP4oycw7aDF2exRRrXf1NnIQxmXfACrOc0oAjclO1ttQb+HBYQgezCbyte
fBOKTeCOiZUzN2Uet62LCW8z0htn/Mj4f2Na6hSKZBtqTZ6Z0Xdjj9WybYXaLCT2ULumHl5lkH/d
DclHlLVRpsJCiSu7mpYY0nOladP4s4JgfYpCrhwOTCO+/0HQkcxf27em4kr7WfPbvoBeBv7XTmLx
TPbCk/2sSaxo8QTFyVqNBAW6Gl+YjYZMVaj4PTdGj8ajRrFtAwN86PAom1aLAs0lb4JKIM88UDU+
X2za8fbk+R7WqwJAgrcNhj4lb+86xGi2djJCZsat3+FYO9mHc/lqz51iMbkwLMenZUawVpO1J+1P
QZIN5V3cl4g8hTcbkGNu7AWR0KV5HW6A4iLmJ3Bry1RiNKbDdK7LGVhYgYrMVAf0T67wDb6ManxA
1+P1mouSOvhhSwtmRsUSzNLFAmBbO+a6kkLwHO9m35Cuo+sHcucoqjqU7l9MhVpTeOvTY3XYGUn5
wX4CyPld/NFptSHkuPA5Fyzd18uzLLPBRs8au+0qRt7DY+RDXd44MC9xMmxxZRAn03umzn8LRcZf
+AYIwYySUFbppPG9JvKEG3OBfujcL+eI+SQgysQxdmDWZu8Fx86w+z87Eoz9XvD6y9nEVz4gz2iJ
egLB7t/2OnwihX8ji518YGjXsd5IwHFPYeqJfJi8K20fOYrmMK5dUMgs6NRPlYbywQ7rKGGlEbFs
j6cg/iKgiH8kLtnG2gBgTFScLepLkgc7dHY+P5D9HADEra8neyaaoEEbBJwhmCEzP1Bf5dgGvrNt
GcQdz3go0c5oe4wiNbbIbG0KCKTZSqteAWUMGUwH8go/IpV0MhvMHqHHtxP5drf1sUAvhgVlrM00
vs1ibVg7dEj+qANto0GOraQ8RQMard4l01ZxXkZ0J5L3BgZ3LlbiHYQ26NUq1RnzKyAcfYyFQ7p5
kd+5yqnJWLL8buudTHCR+XxXTtGwMYa9S3Hu5f3+WYkiqu2Wxz53Bx6Eui27FOih7I+yflRR0Cxq
3J6lfJUESn3/yR3XjyAazWPQvhY7aLPn4HHUmFEXG9Sh1DOgs7LlkOBynsQqTsP1/CjbXOu4lpBG
I3zkBcqTK3WiWsCczRmXWvHlPwikA6y4KmpFoDrammvnNTrBKHOkOiLYKr5XHghP7yUEAvekASBH
UWKKmg58lyn3o8XmPXgfd29F3JmcDjknXpuFK52nlaGjHhTRejj5rYnFuKRZdz7aKZ1txCEnf/Wc
W6HZpnQ4Agml8bsjndx893P08lWFrPVTIyt+Xs5MgI9HtEoTNdC9wjI5/mLC4dB5wPqHWlNLWOR2
r7eTuM57/4OXgo1s9GPcexlwLB1pmBICtGnC6/DcjiiF7EorV+myeBltkvy6nkYX39lHq8Z10wiB
XqppAWBhsrEzGQT3inJKm2u9O+AbS4iXRva3oWtqSKqZquDB0XaN56NiSBIevuKPfMaoS8VQfDSs
IAL/gM0ZcRqeXNkU8gXUj0QIoKuUDGXUe5tZE1yS+K5D/Xnuhd/Qetp79rv2erNGC1zEf0FSmtL+
7AAzhJsRh3oj/dfcNdmqdrmwLy+gjbZhGMOT3YxdajXuMhyiJXLK8y0ihsv68HJQ1mBswdJO8pOc
pT+k0YIGuBxN4nDjprnwvRQprXLN4KH3nzukeJBgaGl8XUKE7Oo22j2u6yQZ455QFLvj+DxTaPEv
cXco7ZHlpJ3Jef6USDfHFX8JQyHAI9XppcGTGASO3ZHCplmQ4oRquMY+SkbT0PTBauRzux7wk0G1
WLHBdIzDkhajNSzgrwH1HtsCHw/F6bMD+ppoybou0k67ytDWw0GAu29WzOWzEA05AfJKsXMYDuOk
tsLF7PPtwPWgT2LfELIRgMzxJCa1iP9Q42Lg1RH3LPiEuoT8X2acJxPXlUCZkout3WDw7oU8Wlo/
kSlNjAswC7a16bjXU9PMiOdKygcSBTc3iVur3Nx4Cf1A4u0fbVqQxkwUE5VJvME7h/OqnKjYfp/y
z8V2KG26hQ8jrcJ0ip0YN5G0uB/SMTfVQr1DLSrwGaO0JdusctzHDmFNSqKYbViHAtI48QTzfHXj
IaBlnDGYtsK1HXwdQB+VAG58Q8lxNLvHLu3KyeT20172CtVkB1Rsu020orYbn2Ip67bIvMobVXui
PEuw1NEZHWA4w22GIMSvU25RZQIcJnO5CNDKLeRXpxJ2aIJAB+ft7Y8oRSS4K0rnLiieNUKz4ngb
nMnMdUp/KVSS7G1m6FrSmO0Ygq4+czZ/W1GRqYi2pAnmZkQ+PW16e6CWc3gnQ3URO9XCUhp5J+sx
WQvEk6x9wJubqofThEJ3dhCU0QcPklFbl5f6/8WKY7TvfuSdtNyrMvd/0bkyyBHwi+3tFu49SKzJ
LB8V1qRwTneH4LTyibuZGnWy2rfbvCZkNNaCKMGZQXTdFZJzLzPO7enWYap+FYqfDPv9qRbBmiEr
em8Otvta/JyWX2mJi56BtRJ1r0K6e4RNTQQ90edT/RCT7kojirPVE2gGy/GOV+S99zocfQ3WsMNX
qHqKm32FEUrxAUxp4iZdU6rSALAYSzKEAAi6FIo+rhaHuL/lZC54/RYhCFzdUjDe2VeTBL+rfZLF
+iWV6+/0Y/hwGadQ1B5XyPfpkcTdtEohHAJb4D1TtcArC9+CSNoOloiFj9y1o39sfpmqpoI2r64l
Sgr4OqgShC0Xj6NVEMHNqkK4sAxhB98h0FIiEMjPkhCcxRoesf+T/DSGYq5bltZoJwHY0gsB7uWC
C9/URvLTkMH7QuKzJOQynIJd/B58WwMwZU4MSpzF6COp1XpaJt0VT5iFVuY4u8FlntVXwenBSpEU
Zzqq9fp8KSPTE9Jbw7cguB4M4Ir+ajtjoLAaRWVgxRzLbIH5HdO4DZ3qZUGjqghinnXAy8lsFuv8
LSJAcMU2p8tLJPXnomOxP/1ZlYs019Bt+M5GwkoL4N9KT5Z54t01Ug3ybVs8YUNN3uWnRnEsAfBA
89zfV9HqsoFyN4pJs3a++QKlO+3gJ8NnmPUtNmMzdB2NZrUXIumSrGIdKaSILQYI45sIlQ7OejCg
h8Y7jUL+wMwEDgrfkXXgxaxood3Q6t3aPfh07eIeTPvkqYTM7884Qnevn3V+K2BKSEDWQ0tW798I
l1YEdklF1Bh5BFqK6+wAcYMu5qHbF2+m3Dt6tPUWshpow6juA7fubMHgtml3uGvyucmClaLB8ira
p+DHs6X5A2DqGdD4VWhuS1VmvRnyMoNMNwSLle4310n3RKfgleuerrUUWvAd3DAHfTFEy4HDRvta
Sp0RpaiHgh1bVF/xUQybom06V6mwMiyva87ucMy9b0J6zO5DsvXKEMybOdskJvuCEBRJlaE7Fhj/
OCoL8TwKVPFC9rVRtq1iodS20FS7t80CWGHG2U9FtFJEw0NJqJcVwAH477fZ8N4kaDMH9AkDgwD8
kGTwBTacvtwELoomodwg659pFQsMYWgNKRN+b9JIrvcnloOV8q6LzQpTa6ux1+yRTv04pOQRMm8z
Sgl2GzJeOYOKYPjb4yCKDoAQ8CNKfIzjW/CeEAH3vGQIZZmE6R02Zvew3FvsJiAYxozxs4LWfq0P
/Y0rkupbSuzfD6TLsUZDOuQQaElngm71nv81i1FwcmTmRYQFRnqXMLvjpqr+X3ISFqbBJa6SnER8
pf4gfwpB07SZlPBgl8vfeZCaBTIB4/yTJTcVMfkQ1n8T+Mn3yLO2WbTqyKaWzJP7AKiMdFPJ3lFC
TFQHfjuCigooNyYltGAFrZzjcHcfsp49lucNMV6ltjazeM/tiMdmxs+qHVF6DNNRioZqxs9JL6Lm
zqDJlFENPeZfL/T6RKaCZeou6rH/HbLbBXnUhlX4TaCa7chSXy8YRy4loQuml0CcSNQ6WCxzfQAq
cgtmtHnkc8nPnPrBb+PjP7plkpTJqnYJmzx3JBNXyN7f0o5Ninna+QVn3079ODFhi027jbvIvNnD
rew/p07XRZy9NQy+APT50BrN/XmbBr/1KRaa/j+KSgdZiZNslnxDiiEtAkAfXViUqNOLr29/rwHh
H16hAG4O5eieTFzq0Amdi6OOfVNFP5hyHAn/Wnp53icWnuvEWWi781hO9BBLRrxXJ57y3cnrA1jT
mkXJuZs3ebTcJdt96ZNaImf96vjEXpwiVfjAo5zaMd0DoC27HUnAebYLM2A4WjuaYZbikll+CDqD
mhjrMnodRzN5s1tmDQhzgyG66CmeA41B/Abu7/lncZ/45Fq+B4pvFfjKpbtgztmAqzNEthJhI2zR
aBiayq0ezxnrp0KcD7YrN49n5nJbiPe0Gtpudgbuto4+IYNvwpwyfDAuzdJMpJXJKhP3zEs1uA9+
M9U++gbBGtg7N5m95DUplQntzrFCUTgQpn4QubGBzXbG8pJiHx8DEaT9GS/K+VDLf7C0AF0j6b95
bkfDlxubLscjZ5vHEif/F4KpFCKpwHG8IbFO2xtwO6EFYjdn8Rm3/Xwu7/fRY+DkphqABB2VTiA/
SOAVz8+M5XLTyWiTTjTx81cXPIRLSM7J+Y9WqeZKrWQF7GSxdqc6QCTbR0VZ1y66I9Hg2gUQU3sd
lk5BLXSzIwIyFKQc3nokzDhbn3aZb1kkky6yTcV1foswVq5Ap8anhFb6VagTQU5xajf3XJQ1xXDY
ZGc5VH7GBcxsMasieqUejSQSDjN3cR4Qi2/C7b4uEMLSkMSpJ9cZw15inUPDkhn4cGqNVrZeUnR5
nJtiShPZWW0Hb8KXXlRvgqACLFy1JbQH8SmQUhcSkAvCc4Idl6t9mLAGdLp970MFs+NKwNlBYy9j
bG5ZSxRMiV1Czfk+4ww0KQhOqyy6mnvveXl6kZdrxGhVl2gVft7q1tvsYm/NEXo95ROEuDTQFBX5
UsnoygD0De0XUk1QIFpn7rfFRCLg1RynqR7YfLmXwY4K5asNUGvlTN89RfxpAltyP2iBN2brZh8t
vNgCbhgl+1pk71q8T2FJTC1QnPLzPnx+TJYCtp8rsGQqAAeATvCXYGUkhGnYXhWOJAekfi2sAX1M
OLNh1qinlJ/x7LFdkgGS0ZgQHHger+onL0aeQ0yvLqaKl/Ai2IHOj8h7T4TErmwN7dRzV9j8Eb4S
mMOmcI+lcHLP5AuRFkp2wljyGCjocggNCXGj7lVIMMPWV7bQE4ceh4Zi+zzeA8lMdLXFOhdWeflK
xvFzGIxQmVT2WSJvFfRrNIvqY5pT9n7xoBB6rfPSRVpRHopRAc4M1QljPO4loiNd2C7dtR3mptQc
Mn98pXKbInFKy33D9SI7j+CVKuZHKCBhfcfHfXoC6E2st+t89gwH1lYZNkFuZVxrxYqC0LYbt2E+
TZxw8IZxmmg8aY+RSRSEawlxS8i/TvY2yxoSgRkqu/RrLZxg526+t1Og+yY4iC1gFgirvV7dyF4U
1iPppqjpc5PcenkWhqD3EcOAeXb0zuTb2/lMOywYpXcL7SIlWiQgVdSNxPzzkJ444G4XoYAIHVz0
DkCN2umuCoupPFmsXszuUaQEw3dgjDBjgrXnizHwD+kJALT09nR39A7lrpvbaruYWdYVLhRL9Cc9
k6jXRrW+CXoJbOI8sDJQQMnFfOBZWK3XN+Pi5mAhi1n9XSIghqPsiOVuJvwKGR5HCilfB2EWbt/r
QQWhlnMGtbf0IHXGMZsSTaEMH0mYBf4D75SUAXofVqdbPcyF7frSLBygqjVMHNawJjCHpaDNnTCY
pOZ+8nX/kNzAi1FmD/5PmH3a9ltsxuKztBgi5bwIHQPpTb3hyBLoepVq5hKUk6SFnCWFQQAF6RKX
97IlSWOVadbUVr6j7GWv26i6Gd0HT9/ALTF/tI5wWT5rhzFMS97CWKp7CbDI30KkuvStOkLQU71O
tpXXY1y6HOphj1Ud3Hbr5ZZOxA1WlxH2yRoAuMXSWThkqm6jsKd/1NrzjaQH4xlswrzKjpuM5QHB
G87baBm8hvpCwkvGiDUm8VbQvJ063ZFCk+Zp9N4n7AUzElHJBvzATF0i3yvfDgdZNEDEp46eqhvj
Yt7bdUlrdJr5/G1ZZYE3U8TOaLdwtOW8ixs4eZLtmznMKfyGDHrAg3DT1sjua0HKWys6q6MjFHKf
njFxvzyjwFX75UOcwQ7exBpIGE7nwCaNVQs86UNKu06ClxYpazcw2rDlhsSJPAbiT4/jR0Qpowev
HAnczpw1YtmZmL4nDwJ1yZict3xDzGbBUUAl+SIXm3uW4iTmcTynC9yK/vzuqs7okBEhfwp9nIEf
x0jk5Kt9xOf0RLHONK/WYw2bJQ5igf6rIR5z6MW22zln6aD6CiNM3sfFZTchpbCME0s9JeGPHC8I
viYfI60UKB0irWUBwtPk3tdvykXPkynH8qRIty4Mztjq1A1Yb8VKeE+Lqu8QclKO/6eCItP2g0Jw
PVum9V66pKC/PPDHGCa49nlFqhnJt3GSGORlofti566tVmaImyl2HEnEe69tcGgBmRXUrPNRPz5O
Ryte/tF5CWA8LzxSGg7hb8uuoq5qZFpl2nKtEwL0BjsplqEyIbdzwZVCQ1Jo6ku54XayzdDf7pyR
5kd60GNabrBfqKKxRO3lWlTDltIjVSt0k9lHAA4mGw6xrwd0itsc+wB1IRx78qIXcc54FBTG7vRi
WJdmJoQaThGyR4zUpPbhkBnInzokMnSzXIrzNA49DP1kaQzCknDLGixdhylLv62GCH9qovXMmsLK
GBkSIUeLqdbZ+JFTP4Wnat2kSyULvuqfm5yIvWjShcXF6Z26UvpVjaWTKAxnFFElMbL8E1MsJUHR
8dyX0Ccl+z2BpSIkQ6fEcHVcBwWKFFTJ9TEFYPt3lW300SqoDOHpQXKit5htQpgPE5hKsY/0KDQo
+WEqOdyQghC0bA2buZcOdCL0v1vCJ2XJjh7iJ6GQ0z5nbdRt1PQc1ZinRJ3NXfyhjzy3es3vbjIC
JHK1qyuCHrFYJ1VM7jFBSFXKsbGVzbu1TiH3Me1MEwXfVAAXAOydP+md6rTcKZ8h2AU6e1OSBX50
GFCsogOW+IWV/txA+NLtpQ/HN4XkmgolMiUujY5QSSS+UVuE5GQ0Cr8Ug0NriwjmyjRqkCsQ7O85
APiIB1BIaB7hp8CtdI2mf1sl0Gbh+ctl2kX4asqEsm3XlfqJBqHtgtKPr8Gzsu5o+jGparcIt2s/
unpMf3x7Sq1330t2u68GFod62f72/7Zw3LUEtP5UUTK6ujq+hLianMhOTZkOR5SNFMcxOb5FxBup
7P726m8IsPgPv3W/hu0rL0Bs4fqLgUwr/4rn9kiYR1ApGMmR47RgPNpp+VIe7RgP99o2qrdlmxWM
x0OQiy3eSByYRr7i6E7R2ky6sQZvOMSvdvIZIc3ms8lJ+xJn2Spu894Nv2ltsb0WkTv5rF7wmmu9
hshOdEogk6IRIj6l9HdbblUUOg8adchjWL+Knu3ehsk6HE0iToE+y1QC/R0pl9ouh4zN7O1MWXM8
wIrt5EtVtrsKJjV6I0TDgbP+iftMALYGRxHG+DhjtKxlvf9449M2iKEF3wDoK4pW+3wyrKpxpAgA
77AHOjn1ar9u33UQEHegkQKm4ZNyWaKU1vmWRLxnMA1yrS5vb3a5qA8kDOJXnnDg+0Sl/ur7dD9o
KXgFMhQevjcbkF1tAd3SH/B9XWULt7XBH4U/HuJkAqj5zillAaVzJcQEw9uIXaHUA1eOXFrBcPBZ
c2p2/yk5N2Ui3NZxD/F0f+KAnbe+io9xcRx9ehI5LwtokQKsv8evKrZNpUYNLCqT5kH2mAAYttie
mIFXYH6JHXMLDIR+kV54MViDEa5ubliEKGjumfFttxzZj0Jst9NXLznKf97UgMkbUvJBPl5kg2wO
z0Ca2X7d+yZhslF/npmM2TK75nT35sflRwfLfH8SrOiruRDrhoQg6kyROV25jq5+s+GnsoGA4JiQ
GPBHihC+IUPArJkmqJ47osBfdsp78UcJNChusBKkREn/dXUN0s9tfKpMIJSRXbohs7Rva4dO1Q7a
+eNfwsNAbEnixCYz10EYxXNOHylMRhEg+5pSvkF+jnIOVuUgjSC6QiZg0SfuU0bzPMxIoTROsJnY
rs6RNbwQV9jEaymGPXJaxtnWP1to5v7mKpMpTCr13hh/ugcx9Hbw7CFM1k3Kd4T5UjNC8/v6k25k
Rep/BTy9scEgkKEV4Kvgm6wUyLtEwBz5dgoYQZvOxfXmO7ipxC69feb3oegM/mXl0qKxCboHq0ud
1whLZN0NWqBJdFIHVdMRzqJJntyLvchTt4Xjfd6W1gW9NizbdV5PVdnio51hDhYZsNBmUkF7QCn5
wF9iKJuctp4LwHtZhORZtzHB18RS/nJP7n2s6Zu788z8RQaNga/ga9ALd1a7T4quxd9E2gts72fb
I/AZ3lxBkzVKvQGYUbB5x/KBqdTtk4WfsqHtayvue62cVfzdMCHlo5/nAFFkK3U9QZ+b+NYI7QMj
0v8u/IggAu3J9x4Oh9FU44c55Yx5Dg6WOE6H6MT+oVzNTURyJOMRlW+IXlzl82AGgQjQgjgZU34Z
cC8Ei8ATUAlHLlXTF2U00dt8PcFri38RmOTOQ+s5MRQ7WY+gzUhVS7t6D4JwuMi5pZHRK0tVWc+y
ofbo9ErrgVYWkeMlelCQm7UK/JpmFLN98oq/D/In5eJNJwyYndkIZPc1ZfiTeGlKzQKASiu3haoY
mq6JPUnIik2lcVYnTrz3bfOMSSiNCsPS1XJN6i/2upoJ9it2Jd7xgCo0QOgtDcf98CUiN3gAlFj6
JoqtJXL8r2H5wdhnPx7DkXosqa0CbVD1q7OFtn/wTPbkiiAL5ADeZhLUMO4joAJth6BI0j4AT9lr
7Lzdaxc4XfmiLX9HmzT1rI38wANfIRNSLzEIFSHXScjcSw+uVxIC0U7XbrJqR+PDI/hJ3igAsl1I
2oeMIfuesx8xC+DknOLyLq4YLuxlqpxkLHXzqQRYhhKCN93cpnVoQ9hTX+7N0Sb4mz2cpdlEotxk
hEZ/EQduWB6TvIQfVdlXo2RI8HAGG1tL+WZ+ZQYL3MFvCtd+YbmEIWUGLaT05jz90e39I3nC7qQq
165vfUhXTALm059FhI2YswXh3ChptCn0okIFjxoqV6LClbeEHt/XDWaQLt5jcNzd6JI54ZrsK2J8
deNBD4uPCc76gfmy2j+G8hCd650pyK9Y4f0OIvlpMrpCU5PfVPlFWf03hQST78pVfXleJd9vTLcH
V/azQbpAhykYYK/XL4jPPHTNTdyXnLeBZop/5e9RFrYCA3RaLwRN6vej1UOeeVoIlev90FuyMTt7
Tru6fB5cgQAaKp+6+7GQGzrk+nXpRyiUTElPJRP/4n2jImYYRdQxOmVJQ9+0JQlDUbyl0AWTZCJx
RLfa8RcqsUbaDVCCVWTTlRfAIW2ZZZA8vvDxD44rfitVzSswy593ck8Rg0JTDxi96lAYCebik3UE
2tSAHYdrO8jlSFW+5p2SIu26DwdmsFZjnEONeGG/13KkBYAwJ1g2/xkueOVlwK5wSeP/jpHBm5e0
uR8v74hnJ2sl/FVPX0pD2pPyNZX2Eif6u/QGFr9s2RzVYnCA8QZ9mz144qNG9ktokmlEcM0bZ9os
3DvbUQ3i9938dgCymPu4BvJ5tjPioOMSRl0l+uo4iYwAVyVmQrMQqUq7NH9c9y4mc1EITtxT1GaI
hmKrRMkYwTp1h0/iaCC86Z9nkgYLS3fhFMrv7624AhrImf+08Tf+cd5zfzu596ih2P1IPe2A1Sld
MjOicuOYZ31JjzTagRKW4imoN6dnhE714RFNjaD3rw7EiD8qje+EX/hN2iqRocTMAo/0AD5HEE6Q
VlkOB4rS6PDZ0jM9Xj6CHo8mBmSJfpEZN0spvDjSS1SDzOAOpVHZRpsSU/ybrbXTBJc34hg7YRBB
JkEx114rcziVs4JmQ1I8P17oUh3do6J/CgBGik1HoDfS0cYHSjNsvn0V8OvbSYrFBmdpjqCmegc7
+od3wzKA7SS7OIZ7j1tG50AHdxO0Bb2+ZEe0diQQbV2O7d6dXuoK1uj++uv/1eJ9jYQPBWuy89Y0
4pNAYA16e3z3Yq+jY0e2pfq80mqzHiC38ELLQuXKdaEKt5QRV3Gxu4LdNsWE3OO7GPI6wafMYIdN
C28CwZZxaNDiDlIECnhySNkWXZ+RLexBvhH30eQhUoWIa5Q+KFBhRlvGQuhCpIiMjHlndZCdYEjY
JIcdP4PSN/9xECL/PmirQfZNJMetZQS9fRxn+IBugTK40z2pjF+55swhDu+j46sNJZY9m53Sgf3C
ct9gzqJvFRMRQrIoMBMzHJux5qxSoiXsVuuwZyL2mTqHhYj4bXCaXJA9r5zyPNxm+ZTvTWPk4lQX
01HFjARHRGksEUVfvMny4LfUk0xYpW3l0vjVwADhZj4s/l/AiKGYPEwCPzIsyAq1g5CqO7RWly/p
LM+IBmKEgZru+2rJqFU0E+la/SzvMU890CrabaGpPeS5DHR6kEBt9ADG6mX3pSgoWeL4sMdzZlwN
eIB94Ky40zv6oCCRZOFwu0GxQ9poSoFSn4HVevIXNbqNkYW1SIjJMPCf7AfTq71kSFS/e/cYpzsL
mwMg2sAgjyqy2qBAVzhejvJPQdSu4M3Y2ytwWgH44RRelgonIfib3/q4XSOnlyqqf87GKAidH7Vl
ElZViy5u82Umc6xuMGKFn++1yQQuXRQCqIV6JpDdg2CRSKzIOKDBfqxMqnHvWWWm2qvxWr75GC5V
JC134KUIq6i2FUs5k5iWSRcbyPySTm1GQKkGxBWIv3yHdUBe1QFaAp7dGjSWFUkwcbiiREp8biPc
hjxO4ndE+nBaSYdmKLqj0Nt7LP6aPNQbCsZubjg8y0gCoQCBPRX5fCbeWfIeWdYYIErBz5ECXW+B
rTnhntrXFFglZzF4e73gwA3W2bpBBceVGb6UkePkMyRwYAHSbZ6IXasy2XBnvRyJm8iC/JkgSi6A
rbkpBQWy5zCHEzXOLnuTlltO5jrHCQZ9/7+VHYygb1X7Gc20/KOLIz3WaijvJqS7lqsWt/eyjg8W
SpE6/v06HTIRdpqh4RNLVCGDrtP+pegHQY6KkDo6JR568iZssCMdyx66XpyccSeqbH2qNojuNZ/k
3RHWyLZWNH+F9iDnZOfcNt12YjBfRXNXHjA6r4x0SDLxB1Iz3jREmBIoDZAjuuaMKT9vFl15EtQY
LI/1bTfzHcHrVZ0n09D4ngcZVd5SSEGiz8N/YojQyM4B6SWwDyQEmXKhyoO4KOdkhTF1+k4aJmcE
UDvip9cbTDLjLUFlKgkxHS7LK0OVnk5mnKQO9GhQs9Qx9z3KZMtdgXWk5VhvhR3DMaIRNTLAD80i
ZKzk91qicLYQBMua77irs6qi9Eis6nPQdu74UIWbuEm1iDulsluLaFuOw39/70hRM1+u8EKamcWp
UM31ebirqLgwU38vwWI1yoGgd712y5SAw38Yf/e6Lw5Omb/zf580RwsHMqqgF0v5uIuCJB/NCYt5
/7UVgRaeNc4KJkg+btQC6dmxwsuxqQYNZ5uEGKmgrDUgxo+LHBSBOe88l7pfSuwu5KviRfiRHXWO
uGmSKHd82GtgMyKvTQFaThfgYWgJnrJgcvhwHbpAtd25X8LZjcCL8cyC/p86kdmkPNt4rUUKIgTe
3u7jGOn1wto3YSTDFAKTQDGDPOn1pP37J8+gs8Qy6ID0FZy8CtBO3rrqzxXNUHni8tIMKaKYr+i2
PWHBtiS254nogF2owAnzX//AIQeXbCJfOylvtFrf33pQjvlfQfCi1LJ7Qd+WjZNdvGsl+Wt8L107
FWGibEIC+7XBY/jUZbTHRYqw9HJ7y8opmMKzWU0VJYJrJ/4aZVxEX/0Bma1KOxnFtlbdAt2X3DGU
ogL5KNsmqA/ElR32NJJz8u4TO27+/fLy8acWa6707pd8GNzAm6dA+DaY+aEAwgISzoCBJye+yIiO
V+lUG//WTeuqEO3DW/F3Xqk+zv0x0N9xbIJc/9TM59rQP9gOqsjliVUotHL2sQY7OlaE9Sl/VV0U
ArQcyx90Pupt6QvnG0Xp4xQ9lUi42DAfENd3gFljRj5PUd58urAij7hyYFcYc0amezACjymlJ22f
rxrtLHc3pzPNDF3nGMXthzTVk7DZ7+9YI6+pVMoXB64X3ExYr1NTwWDfAsT/3c38ZmnT/cIo1Dgw
YNmET0klQkWVQnzJ7vz3Kls4Qv2wqNrQH1kk8b91W6zstlb0NLomI0SVSRNUzWrKqTPtcw+OS3ze
TEQd7yZdVycaJ6yDBcnrmzZY2EaS9g5TfPzrYjObSgU1qtmVh1PP9hPI9TM/y2UzRGK9T6YhPcHb
LR0uakBbZahEDSbY+oDzfSamk9Vb8+FuD/Wx1EhHZpNWNNuj5BSBFWkbfylgFtlCq3nNURPEFZdL
rOqLvFyDRzf1G12KBmRODQt4dyi1aR9cgjA9AoUBHkooYdCvRUs5nSq3xJTleu6Pud8/IKWwax89
qtyQ1iLyLstPv7XOEeq3JA5ed64bwC6uZNiyQ+z4W8uMUJEKKN+21INjgWCbcoKJln9/fo1Ln29M
Jkdjk90eisqhkq8hDOEjvPmJOfd4GSGjQO+hYW+lDJr5wdMSyyVUM0KdO3iIEdITDfl6M+6jbs1r
Dygy5PrWLmkdLHCoDEJE2SEckvgBVpiy+3rWYgnWiRsiNdhmrmF4j7/2YaR977kyjKDaKFw2Jurj
I24Yc0hIUSbPnkep0/P3iViHTWjI2RzytHRnYpzD6IWSfXrMyg6Wms+eUyuX7Alfiu9DBaaEzdnM
n0VO/lXRWJuFV0nFtBd25uFcpRht/mYOM/eBUDSuJStdJAjLKa3BDfP1Hl1okFMfbMEzt50nTz+3
nMMuSeDmgbKR//fOtAI2KmFDKFHbuWzYezpRjJXIBR7aiOIucm6d2TRR2XNF2JLffBAw1JnspwPr
ejHbF5OEsuVXaw89eefNdZu6cERMTQZxcVj4GRqnFKhxLgpboel73sA/n3+9sw1P8NQu843dFKA7
qoWdbQHMDdHqo/UI24ft9LY7AmY+xWqTPVjg+BodsqJ/uDK/pX0WY9Qsjonx+n2woeCdSqh7vr+U
umIaXZQDx5jcFzQSZRY0SuS7bIjNumO6c0dj5vkd1fQq0iq5ZCgkJniDCxMMHeU+uad4RcQuUboE
5OpSmFhMXdoe81pYL2Uy8xZLfNy8D42yWBF+drzSbj3rEcZubMvv3rIulYEO7nqLrYakNE9cdPEN
qA2jfqZgc76ncaOlvKjGeBo/fXs10Ssz5fCRNUK+K50Q74iKDYR0qvqlX8XIg33lHleaSsFa/abI
u/ebSJivLJ49+yIC0sMLZrTEEwD1OfeqvI9ioEWXLW6QLkrdhxr10ax/MKGUyHvpFa6TRlPXdqL5
1Bkhjd/ABfA5I5obFmGCzui3Zw9bIbKzTrmnbELAk+eiz+wYYm8he43Mep/4tPuFXx/IRszl4Gml
YW4qSvvq1+g8RhuREjDWmNthN61CsXRrk62yPoVlk6TbQNjpSJynyQfRub1y0aHk4pDCxu4d1o/q
YFMv8DaqB+Pmeh39ZPR5r0QmH5rHO6IUiqgETMCxURADHU6v7YHb1X/XSsZn4dlwZKCK/1MYDAYW
mcRRr+GlVXGGnjTdksNK81YnscW86shCFJAR0S/gnFFEvX8XU7txm7yB7aqzju0Iwbt3vfqvT03d
2p7vKeKPYcOL27yO1Y4LOYDqhcmehdinKava1rkex4UaVJdwBDHKHQH2d9AqqvAdAAtkjM6RtPDY
sNTPsjlheKQre5G5Nag0hlLYxkjIVRZr3No7kfP71XdDw5Tp6ZNMaz1SraJ2PyGtQEYsn2L3v7+C
r1iyA6JG+bDyd+8hKsBoKNd+ikddxpnsBgvkt0OE7bW+W/KO5Vfq3PXXY3JBMz4Qb7iSE/K/pbAW
Vtwqf0m0Q8cOkXbdZFlh/oBVPp1F2qJLs3IX4bIEyOhbzjAJCsGel0gDZY9QwZLHF7OywxA5uWga
iqrXkqjSpoLn4nyztn2Wn2vjrltpvi2BIqAg6gcyV/azfg7va61pyEBItpTok+TCOQfhQrSo6HQi
qGEphfd4wIby2MfwKM5u+2IoCy7gGyGsqEm6rLWaI1DRPgpE0MjHvSoaV60FbJfAIej733PY/QE5
+oMLr9zltac76utAnbVjgpt7qOPyPOx6Uson1HgJmIoQuVAF2KZSdlwEtwLaXpplJfh4vXQGUjUI
mzNc5EOc7OD92N7x5AEx/kpRcSCnKip1+T8GAgDy1Lf4BhQIP4V39MWDHbZCozAxLkfo6Bbc5cVW
JnOmbrb0xPNunyRI5NbUYpVnqmvGxlVPHf0hVFzr62a0xiGCAPn/VajgUUt1TIJmrBTLs6eQE+I8
HfFCLWs9EIIb/zBD8/17mEijbH+wQboqn/qYjQVAQ9vnI+8zRkxg7/lw4J/SbSMpPXxIOBtJiThi
8DG1Jv/w4PTAlG7VeHyQfScDz4l17B+MW1zxCEnDNNcde7ISaOkDbdE3pLGTHKhB8KBr20TewI/H
IpPyiWWxvYavTS4lcoF9mnR+RpCq4ubtOg9a3Lkea6CIH+QI/A+tZi3/4NWwirjoMLfN+hT5BOw4
LzPeKLHsDKqQr2rYlAbludYkv3livMR5OAwJK62rrMDxovWq4589DSofSXEichyQoPCbzyvP/ddu
Wb2uxxxleQZf4Ahdj/BaaNhushkBDMNxsHMOpRR28k1vv6ivmY5fj7YoRlq/8TsqmvvOlyYPQCyy
tSp220xpHWiZUCu1uryoO/NbUI47JcGOjJvoLRngR84nwEwxlilJYuqV/JPzguyD2FwK8lKqNiq5
6+vqrTfiioq+qhxnAMY53CxrS7Rq9UcTPLF4cYPy2ZUuYoAHXLjye71PqOIMuiKzDUM6mF8+kPcr
RIi+ODfIFLyVcEQIRqYaJUFfJFwNzW/y7gHdLCf3CisnVKXH9yfextQEZd5BcB1yaXAqqMvh4S54
LMgglTarS++hbJ8dl+reHtI6Zgar9rnX7/ZRZbayAyhy3gYEEhX1X0JeWIcaxP9Y2G9TZJmonsVe
yuXZ/CIjw9YTzVzlET+qEqPBiBRq/7BSbAC+ZdYvA8KIlJh61pnADfmC7otjZYBHl5YAm6W0KeQW
KLjLEhMB0wj23KnKXJCV8l6piWHKXB0wc+1DguSXMMhXaKl2gijFO8fNwQX8w95SK7WmfOlXH9Ar
Q3OnUR3Wc2niJ+id+egtzi66x2YKULOTxg4vf3E/uYb5UY9oAAtg3nbrGGOArL6rISmHf2eHTbi5
CPfYOeSj+PG5sFq/6aSdlemj88jY4nRP28xS4KWufABqHX283A1y6ioV9dG5KwS/gxq+eElm4X+E
RnkNH3/0CLbRDustDcroJVW/POPLW+DhDVzgLkCq7N/6Ek7eoI/6ah4F22fSAzjr3rYQ559hMU12
DVuMsVxaIEHudXHpFCzAsjPFEvBd6B+kPq1cKOSwSOVHrMcmAl4IFN7j/IfgyCxxpcjignmC30Wh
216fEF3kaFhX0nvQEeswaDnEjO/jz23TOQQyXCCT2hI6Q2rf+mRDaUt54eXABR82SlvebGCqcngl
xQXhucZMMSm1Y8iX2hB96/wVmTJUydpycAiJ1nj05OgBeqjATV+tHTH6th+YtsQPmzP9+4ADJvJP
bI/mOe5DxBVSVlsSbbHyFspgLxR/SZuuq/HBnnnsNZK26KdNHB6e1A6sL7ju5TQxV1f0LnZIz0Y7
vqzei/hdNb53BonDU0GAUF9NM3ddkiVfjOu4wIW0N3d0tBn8p1gIBumtxv0eJTt4jarIyL2FzMQU
7UOGTZqfFGIpbzkusOKKaBjuZn10m0aayUAXUnXLqkx+t3KUWIYpxSWsjwBugE15sDKvP4wiNqnv
Z+D+claEXk2FHGbMMSVRQHh82mJfY/Ril3p5a10GV6cTf2KSBQf8Y+7gQWN1pLFJLCxtteFfZWZl
0vBtuI+ZDV3i+T9PgFACSW+lfo3GpwDkWZ8eXUA9bPd7F3BJP61ErbW90m/LbBgW9Frhz5g7QwM2
Sfshf5ESJUtTiEqe6XJxx2lcU1IGnsn6uycriNtmIhe01Fukval2LWJH5xZZ0BfvpGpZ3VM+Be2y
bL/ZZ886EnwHleZksju3sOuBeAO0H5g+X9Rp1a5iniEFrDS0indzzrVXUqTnzzfh69j16csjagHw
icSGU7tZL5GoKnt31ZwkCxkKU60x2jrzhcNiINn+UDQs4LVOnaaWzsbV0rfqZDqcoqoztWGCiAs7
OTiFB21E2INDoSurp28tXf2QYuMmJrgjRMrkbfHEK6sSXeST2MhAUupvI00t6W6VYkBvQnpXkQ5i
J68OblflhApAm88t/1JTC7zlAXodKHf+6rlvept4B08L8Y1kWcqSoDCQEfo86vsswo+yYsXFs4qX
jD4rhPO39lOwdzV0TjdAZjucIlAFYO3LqFlTeXsJu2rbgNpAXwT7bTq0JB64UBxV8bWlqd0F0eza
jtc8i9NjOG3aehWrKpnQEZrwH3QHnwcY4GfZtWeoFXObvKg9fhFjo0LPEYncFgNX4vQ9zjyzwruR
zL8/UJNeK9jY349mABxxLlbQCZrZ0jTV1xX/8fKJ1/qEb+FggvwanOfZ2bXcObYDTmjSXX4LGw85
cGNB3XL/b2QT29lAVNcgroDHWxji0K3SE0aKanRADGaS2v/5dN33CBnD2oQzQ50hcD/VO4hTSCtd
qN3sW6+ucVj/fZ9cuvtaKa67mR+iuOUvltVMl0LSpaAZf2v347IgmaoPkFlF92tTe3rh/eiCk+Qt
0vOJoxuGf3zuCljmhySnofhtPQ38om4J07J8iAzZ3Bh/mmU2Wyi8Oj2zoiXLVy1iYzKNISR4710C
6oOReiaGXHVS8S5vuPRQtdgKYb/2gDbVE/2aX/QmD3HZHQpHd9SDyBdWU7bOXH9x7mI4mhT9U3n/
ds6GOQKOi56OGpeHpDBylXCTXhEiF2cpRaPLTkVmbTKqKHIawtdLFsUD82YFeFRrxyvO5v3TSbqB
bkaPOylxGrlA2OW42KZa0Y6trbMCo4Y+tKj767+NwUfAR7J5oF+nmurnsfBkRWoPRGmKbebeYNCi
crWimEEN52pfhuXnBo2ivNSZpn1ATM2j3C9Isx7QtN3NLFprCYEn6k7Y+ABzb0NRpRsCJ7DJVLOw
IWT5dH3V1MYjEbCkLvdRR19nSIsDSn5ueUO7BIbgHMSvw2Gsyjiab+zpVRGw3OjCJ5h8bBjKuAq5
VVKSDRF4341H0dkkhpYRpbK+7Q7UxEn10VNgDSP0fuDr8yNPfm/EqsepM5UHbykxedA/Xfz5LgmY
FRuBMKeNCKeHPiUSYwBxCsCH/P7xRv1QVSMj5Jo0e6Dh0mTsslmUTlRu169ob97F6l18DxqZHzcm
OVNTknOaZVGDHABrobczGkBoMQ82WpbRcy0qy+PCJo5Tm/78pOLk9G4PLX0oSixGzKhYK4OyRait
+QSnp5mYpULYiDQnVsmhwgj5pum4wftwiukiCuT6eaJIUHG2bz8Iirazw2KLNqRl12WdXBtYzSxw
BtaCUNLTZoRbZUMyJFA31Vsg2spDVi0w48yt/azzgu4b4pFnjZ3q0W8eOv1AO+972YeA6maGXjxM
9Ggrt7MqSbG5Mgj0cHTaVONOWysWYp7B4lgIAhkVasrd6v67YEyQXMoVhwdxIBw8+AGNX+nHYQ2P
USme+JZPaWAiLtA3MBlmQhFE8PRLoNXEzyhXBXAdNNp9sMMjWHo6U9xEvPDtdVJBCKtP0A/M8LKr
2QdW4v8KFiQr90OwuTDqrOxvoZ80lMPb1qiBUTL+u+F+Os00TggT2haaK5HzK2UPZIulCtqObGG4
+Wa/ijt5t+YY38SQTCKBfqGNMm+SUf3zHv/8KJ/c6ZC7hLPtJEgs+lm1kSU5hNTN6/aK/EAKpCoR
fqVEo3X2GRa82oEwttxU+kzGuzK9b91nUqVhjsc191ZUKwD9JObOzuBx+N739y08ZC63P2FemmxX
G/Eh4pF7XcncW91RlSgXauoe8WOLUfDxN4MtpzDRTnRsrhN+BLAvvOiNI3zqXaHdi7P3lsot0y1y
k0OURGihz9WHPBT4/BzzNydu86HRLOGBS+7oFogAF1Qr9YPDa1o/boELGCTmgsRBSXAkIoV6Ndks
+/ZgFupX+gwxcye2JuK7Z1S8oOV9bnciSEz0jgRGl3D63Xb3EanO3KEvOH0qVYbRAgIRXDKwU3mE
qhQ/LhFMK+DMGX72sDhy1uwDlu7SqBjGyxpurbAEYjDSG549BVYT89nCgU6XkJkawkW9rHWGaHVZ
rONEPWtl8aHyYhYbL/+mHpjmBwSpFdKGR7u/qQ4k9R8C0tH2v7p0USHvap8IIW+ormLwVRL8cpao
fMqFzz6TgTaqmbOHMj6//W00R10H6OtJzF0tMQNwkXr/IwbrAlv9xCsmmUnI+sf13a8HOTktLe/N
YOAmwb442WMu+SThvRuJpMHyF+v1met+/oJt/YbnJLZ4jO9t5hAKjtzVijUpyHteJ/oqTUA1ZfZD
Lus/fz9i4qpS4jVRD2a/GhgrH65xGReGTXaRa7RUF2/QDaa1IDpPgtS+NqDOK3x5wd61h5r5epuC
ZRVT8fysPuvrkUuUU/w7t4e9lNuhSWjYdPPoTpfojN2oPmaiIdYXW3366Wlpo5W4a5pl4cIpg1ly
saeTAAbGtt9kTW9FwbYLyUJfEEvARvY/YdcwI7xOosPs8RBWxh5iaoRFPOKv75cjoXOddmRmZ9OP
W5TVKFWdVwiZqnS8puAkIXtdc2K8zsl5Oj8pR/kMD5cOuIdA+Qv8k/3H2R3p/9IqRJ/U4L7nNKsf
mD6vemNJEwedlrvZZKUsx/54zXpa5kjkwxaH2kuYv0GMFk+wzw8kd+f8QBUeDy+dWUOET1YVF7gJ
2p6Xo3C63g+Bhx8IEyjr6LisgFdoDT6oh4Txvm71rCW9WycKvjQofmkVjKMntrLwtwW6y/7+Ia37
grM54djqzaRGSNwj9Pctxp7eG4wqE54sEOvkE+eBRwVSFrI9wHbfPb+jtwhjhMd9vrywilRVWuBd
kO6amPwlGnyMnWtHdDcwYcK9ATFOtMJq/ULa7BUFDPaW9MYwsOPLYTGiALr48EzBt4TRzFDe08w2
uoiRESnjkSEZebRXEK7CcnZAqzCcDEPP7YjdV8k+y0SKJiv9T0jU776DRYPAxpE7pauuxadnCjll
PnF8qSxRqixsmnIcSfJP2CMpC69ASZzQIeFLJJudwWrJ15lYGWqLMMO0rLkcoqd8wQiM1CW02e/t
Ce+5Hv9/8HGupqWCfTRt6ee8+TN28LVGxer4NCqzuCgaob+mm4KGreEYnxYaymjJZgGOp3HM3/cg
zG0lzBI6zVZa9Oh8aX06EPCtBaqGATwwIkvOwKxGdxTgqbyfHb6kotJavgI787CHFVRvnFriSM32
4FzjyL3RRkEusKoeg0BqjakNG+FqA5iQiq43J6BIKxt08fMIPXyFfwTVanu2sFhCBhIrBRl/HsrD
ftBDJlhrbSqFQQKDzRc7W0BLSM5CREIKQt6ieepKJvAAFbNYclmRwQ52K7/m6p2Yk+mkkn0/ocJK
yPNdyjUblHRZfG4jywJ2BlI/FFnM2CeDVBdFyJ5Ehf1vj6xcjmtZrCcAyZvQY+jV/u+bGI2U9+KL
G9h7P16gum2iQ8j9GpjbCDvWhlWt1DovzDOohPuML05KJKJJKfeUEDqU0mDCtfSOJ9/SUpZR0vRo
wKoXxY8WTPokfIzzO21oWDzm8s/dCzDq5LKrHLiIc7yGhUFMmOvkLCvDsVAC3O0gX+pfTPB2lwwk
2wAg9LMVHMXjAjhzp9ArCc+gVVgNaDCiPeseOqPDyBTp63nOcvhrFbgSoIEBR8mDEkvNb/1XSesY
dxj406RgX+99RWI4qZTi3Wae5fEi6Mi2sVINk22AZmPBSfcvHcJ/rC8bw6jGe/sZFC8XizpYuZK6
hCUjrKuyNVGLi3vtZiQZe5Cn2lbEwekrEOnXEfU+JKuMp/rVJSHmxC4BVMVqWG5Cry7OpZXOQGdP
EOp1yHKmsuQ5jZAw+/QqkLwyDASR9o5h7jc87s7UhqMyGdTiHfkaw6fO4IIkY+KaJC3y1tYq8Gs2
UyrimBa0W6MBLEaA9nFAA7084CTUBjB4GIRJcqx3uBFNgtbhltLTLOte48RKcuGuj4lGzxeecYay
QPYBrt3vL8xGmisMXw7BM6SgIdhmkaM91ayT+tCid2/4PzB2bFNCRzt3P0HbdYlINFjkO4z+t/4s
aDkLLGOqafLePO/5kqEfkbywUc+XTgw7P+AUswKkHQvHaiOwxlhssyz5zIUed1xh5PHggWOoCd6n
L1WUdeSEq9kdC/R29RfoNGCns+/isLmuMrUxu385tXAkMSAJ+E6B3oy6mzFiyk+fSia56wFwyXcF
+82+gB8jebNiO9mlZY70wHTu4N+AT+vR0UlcuJR7HY7OASJkcXjlGIvMEnKDMtzjg2ejQaxiHnTQ
g1vlUYdDokvqJ3km2qPGp/KS5fUDVA5fN41E3Sgri1vUYjAFt/dUn0LVCgL8/djwx75dOJwgX3/d
nvFiqOSCSmCfagVDxv2DucFzz/yvgtN197eebkGy0DHUkaGpCKsg9TNzCfuLUwz2uUaV6BXzFYh2
hC0cMrUd035v1fOMBhkf81ja4s2OsIov78hycK79mhAHCaChNPfIWGSpWW8/1JSLTrHQ1xBmBpqM
qW4cGfQegAn9JvF/9LGgwsCI/fCCYYn1cU3b8iomapwIqTSM82sz8mir81eP3kY0K19qvRxY27lM
/ZBlqKqHXppza0pRWfTwHQUgfH31btNLJx/efnJCCDE7PKjiRp8wQLLZuKw/h10LcEBcEXEU0J8Y
nbz72Tn7v3Rmyv9o8sokbpJ+QMKQp5OjEZJxl49n6a3uKlk/o38/T6QANqlpxs170l4k/kw6on4U
RufrkD+S0aEPNO7/210J1MyfuUPRVVJ5bBZ/KCVclBdRC7F6lIkAeL/J4iaK/vpM/f+Gh1sUeurE
tpWUZHOXCjDKYXtjJDc2qrZ8wLmTAXuWXZWdbgR9eZPbiuOyAEo6oTU/1Y1+lV1qNQgAuQRHh57M
o7hkDpu1fx08cSh+wdMfV1rKsj0t6lJpahissQDCsEdlpM4aZexGsK2tZbr01VeC9RKMmnLrwA8C
wwxTLa2hzu76XjnHN5nGRzaEfbDM/2+Mj1Sr9VeafPF5pVxZihYVotxmA8fKt5IdyQ5v/d9Bws14
VL8srC36Y4FQKLYnX3PHp+Wa/z9Dm4XHHayz+C4dHppN2/ztOw0qfutjwrPDZ+8PoFzAYrPMjRPU
ogF1LbnVa1uwkHYGZbiS1bmV3NrzF9rShSoT78AD1xs4xJp2rlGwYITac36HXUtVt4BIYVYPQ+HD
TqfXBG62uex2Payb3jP52TUZ60iYqaC9hCTW5mzEpeJf2ueXcPAJpq9TRMhVMU2jmsiDTP3vqst2
P/575C3eSB/kOScdmPPiU/hjq31mqy4ROiWqKMZcbFCgmVVE1XVy7czfVQkhTO3gQkGz/mUHl5qw
8+ctEE77Xjc/q1dZmGjYBEw+VCCT8ttjeIZ1HF5dqxBIRvq/RrNfg/cohYVw+8boDc51Tg9KF0DC
yF/x+k5AgDiD2gbtXMhsS4lk89jemluA40isaLbepOgYoh7ZwlaTdo86zP7wyEwNF1ULtpvnvGwJ
3Qclo1S4aggiomlleV8IdLSgKZok7zeSupAQCr6xZdfc2guI2ugwmxZSgwhvZ9enXavYmPqML4ot
4OJgd2dNLMx+DhUKLk/9l8oGdW/TJ0buULLztLqwKSb/j/Q5AsA/h/vIxZSS63aqFXTbvFtiWSuk
sN+ElHCwnXt1cYyz78ptcWep8WsFtGdyugAcA87LvFvVUq526X//5OHB0cXMfMX/jkSt96N8hPr2
kA3nnAgcPPRYQmwFn0DryupsJV/MP2dKVD85yl9oT0J2rAymYh8uvCcd1uC7KiEJmJQwrAsljHID
RMQySUq7JynJpMd6ts6DOEW9GbM2ptp/t9rT+Uux994y7OjFy11lHTd9GU63RX2MRhNdg0lcL3CQ
hDvFZKVDgW7FKIHHYvZW41yvlThqjm5eXR3GefzPivHgjRFcPESK/SDN7AvEFXi+xSuwoTZ+Z5qP
zbyU5SGigK6ckUiQDTxb/eMVjctbr7IBH/+i4gIvaFmiH4ifK+ctfygZ3EmNcGs5Zg0S2lhIOBH/
3nLfB3sNraz9W+gmJm55O7oz/VkzoUPFgzTgBGWCCiOnWG3k1YwXwbCr20jbNW+g2AkN9qgWt31g
CqWv71HYjfCo8ODChSOgKBHNI+Yfc2I/GcedJnGMrpyAHSh9HtJ2eYQq2fhDhOdpf1iygW2w6A83
Fz1PICO88gcUj9b3hQdMSm5i9Q70LeePmk+JjvYmQh9hBBbd7kh7iFd3jaFw6CZK8dH0WN3ngRVH
s4HtFt/3uNcJfc9pThLT46s2DDzP7FjuwcB9ditxV3asU7rlKOFAqsK0P3s=
`pragma protect end_protected
