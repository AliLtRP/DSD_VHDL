// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JaLKYf+ScIzxV4AKz83mT+WjZ56Xu6CPCYippzqCP+khtskX3Ym41emRayBhFpIT
zv93QeZolCzbi/2nx9KOczx/SorfAHC9XKXet1z8+oaYRkWDPlLaGnntWBRx7Npg
xDI16h7NvWIhOTqrg++RKY5Mr6s3Cy3Ill3Kw/XsSmw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9728)
qMAUpdYx3zP5GQb7nEVIkIUYYKZzG2bdCZYc8kaUbKmlTDSgOsqqV5mfHUKR7FcG
+prt5KkCL4DxE23w7tA73d2sb6Ty0+ZWDT3Msqq2Yfts56648UtvE27OgII1JDUr
YlYVCehgAGlK252Jxv3maKYFCtT0AbAZ3OJh3tukksI4t6CtL9CMfH7XtzxizyqL
K6CkvVdxnsW6y5GsrNJtQSqO8cQB+lBEUUS8AJ/8ZeUGBki+EvdU/FZYQ0D/jQoh
Nnx3O54TfiA3rnKZkFJInawfKKZOnJR+u6n4Nr18922THX5am7zZ39rYAuLdnyRt
2STrhW7PbZQHuhJTcYV0F16/YgULyNpiOdm4tne6jp2dg9Yp2HEJlYzY08rok5DZ
uUO5/rZkJ08iZaBeT/LM1RNqVKEbBvAp/fEgvDaw+oRomS76GKcQcYZ/PAGcLfn5
Dtl+COHSf2T9j+i3Ecz2OrChp1VgfAKvHxjs7S9kT1saV7Gr7wq8VprbN6ykXAni
VHQ7EMFz6vo420CACZh5kCZlHSEgtuxQ79jRtJRjLip4M1pKn7iCb1uR6TDxjzae
6y8KWF5nxPp4wQGqfEiE3lP7noqpby0M+fs/1m5Cgznn4++FkK/8NtoOJmwg/wQr
bm/EtXvORjap680jsKr24kSRvXkbMDQumhIN157XPhP/DPxdyjRb9JSGPjOylD6Y
gbbURgn8naRfrdprs1eJZcpVTcIc+TF3jFfasacHe/PcaFEnrZVBe1xYuCu/hRWP
R2LzSP/Y69aEz21GzqCM6nO2LtaN9JpharEXL+WaTLQ9rJlG8o6JSVsJtgk8Q7kN
Pc2xAu+JCQvuL1OQmOBF/tFlPzQTlLr6J95rlOdC2CWOOkKQFYHN0uDIURv90UKh
j/iiMq3dbTyguPng9K866Ss5zy9Y2aywP/W7DGFROwwKy1VzQibnkc9Y6MsBNB5j
f33YUrDt8wCAE3eaFxeoV1JqegwgUO/OxbjmpSliyF397HD+SWqHmUHzYVGQKKFh
00npLhqSHyN7s6K0N5infj+hWpL50gd/33zBXDPjkpXIAyABeyCMPmHggzvm/bPV
o1cM4LSY4oVRTSj84jWr4eNYUr6ba/gWAkfpmkNUC/hCwIDqkJK8P+jEc2dmXNau
66/L6kOi4ZsPuLax4flrnGPjBvhXqZUObPfsE5J7f+Q0iLKdg5+pCDbmLMCgjnpf
dGSBnLzkbdvgmBZI3UTRf+mzKfO0oZgs82+nZg4oUmt4I/wwNmJNeastMx52Iinc
+X0uKfyzeHq4nXK50sLCaVGLdWZjYP4jY+jyql3sqhnKsNGIYYGmYK4eHkyGxDHS
qsZAyJjoyqw+3fMJLiklyIjMkZeVMrumVnUPiQiew+Ge8ZC2eFdM5AepuruwtyFW
pC+UKfjldifZmQK9YU+UxFruXgCpnyG4xk/aPfFX+kHdc4syD87XOXCHTlD4BdAr
oq1JVwaixDElp7Lhd+wxJjxvzMcKMcJJLq7x2b2v2Ga3To2FauowtSuiVL8AX+bw
0i4UTsVFKaxqvZY1+Z+y21712+OS4IOk+HZETOCgGSLe4faHy7u3gjpbFATGqkk1
rdLQYVHQb3trStHks+HKvFVYbA/WEjO4kcsldZwtcRBWc2XjzppJqYv8mlYEIqfd
5xzTt1KCiKAqw/+yeJJ0ix078uGz/s/RhICHvsFk5qgo+dl4B2IqTGL9A6+HpcdN
XS1gfv9cKx9lDPq9IwnAHeKrN0CKFrk/VSXXterk5Sq/TcpIkTYUyo61NW6snwVR
xr8HFMKtu1WokZqT43oPjB18C8VEyoBKeRqCwKfOHXNGmn3qAdhQIitl6l+yUIjb
dyDA8AX/wPKTgMdNJb7joW9vEPdPSpNSX4d/qV1Fciq3cKir8WMzsD2bL5X93v3t
lNkH8O1ENxI9heMBC5Aypi/gUwyuQ3tRhv2xhgZf2/Rtdmsm+0ZXS7mD1PGycgBm
GaGiAZ0Nb0vUp7KaIHj0xhK1cQ8UhmrQiWuPurgumvlHd6ycGavxTPqgvmjSjpi3
DSziMfBFIqNnEMfMqSs3M305GgXw0fSkHOMyYSWQ4YgX3oj1TmuUN4GG1NYhrgSh
UrK+cx/KBellzCb9sn/u9liClxjHLsvnB8J9J1NQmcCkrAUxe+CkpJf1lBe3/orL
AZol5mZsPeOqyDCiOJv2RtaBFX5M0i/tpQk8dxTW2Cu5sghxt0zbTRiuENQ18w3Q
etyKc0CAYYa8gBtlK0gJRE5tLVUK++UUXi8nT3wEex0ZYNYZlEO8n+t94WoGclHc
nVtYSDdLFR0OlEooeCYZw44PyJJ+KQ5xTLnJZlBRFf81O0F74JDzFP0XM5Gw+WYy
N9rvHhrbjwwoUP+pwr92DV0EVZIQw0ssjgTh7FuFwQXu6UuC/s/EICh0BVuPsZ9q
37dBk5h3MuKVAMN1VFgTfVBJElMisTpdOu4nA7redxUba4EirKoQit0lKnKJFHAQ
mqRTbeAaT1mKoorFzUG4F3Vdj/jdGE+H/hdflEYbLwwnBjcsIF/Gm7BMnYUGVnoh
O+4XpTlrK51+EuUAuTledUphiK+Xwy9NWHD2Cfoe2AKrJFu1JFUcSfuau+0WqWhx
Jp0YDJklNFX6m+hXkc5s/iZr2+H9Anyf4Vdy2fBE2amtQ9e52JGiYijyZtbS3iKW
q2Gb2tSshb96339LOfZI9ZudxrZCTYcmnyUMNt2WN1kO/EgSHqkUIZ2iOCJ6u3ig
4gpXD1d436gzpEhQYV4GnfB/RtA1cxGIvhOLLbS9qtZvdcooCmxb7i/XSRD/CQhj
1maHi9VO01/r62NVeZMN2GFOlpTbqXi/w4vVMSyhnBLMdH/MRSdnJwKyzF9z78P0
D52mPlrbbQJaEGwehvGlz92bEJTPMKrEonW3RbIiSTrWEQjlXOcfLXl2fcrsYLiZ
sc2jY+smqx1/gtlO+IKTomaAAco8K80shjStYfwAKyWxe/Dss+5RnCAzsWXk8Q8D
DBz7QQf7GRDcaH+0HGkxXumQF2T/yWLtMlQhxf1ATSHWajkK30j0cvZNlAsUSTWs
72nizAJgm/Xz39zpJmIpbdKW6CNRbDk/VmatOkDB8a83aNHvUGAEtsr0OogHHmzR
NcO43OxZAYuzGx23YrezmQXI7ugrCiXtvB9gRYR9jR/H13MmMX9vi202BwHDAvKo
V8YnTsGt3v8b4DuKUcA8A6bwmvBYybeGUvKLovfkH5gIFHI0ZC9dz88aFNIMfVd7
K8n/kPNgRXpRQeiBM1+SGT5XrWrBCT1/UiQRlSkGKKyzkI6Wg3VjVGO3hUl/IvbY
puROe5WTy64KsGPp72fRLoHwJ+voH16HkXHI4lM5uxvo7vyReAOXrp1Qu10NPNe2
Nm9Q76syM7cEVjjCnTCZQJC2vjp+ymhhGePJrC5picQqfGrpmqgAbh33uo4/mkvf
SuqnpCSIfWao0vUYifxVs9MYShtxu4AtcyU7ZsKlC9O+1f6xg4UFinXhnwvJrn9d
r28uXR/RtZzK+AwTx5ODwyHj0L+Zz2Sc8xf/B5Y7DO21JY47SD0pw1ekhnIHkVGR
Y3g246RGFqOVgc6RpgVbWG9vqbBN8kgApNh+j2FiRdGnKHTboEYgmfQmh20YuhAX
zE2cRtZp368S5+DCQKEDI5l7f6D4IPifv+UwyLCf8kEyFGhovfR5R9mGSbl38rp6
TY9nJ2gTzHVHa685SsSblZ2OYZwSxuDOkFFC7tN8WgG7EaffZyUMuuV9VmFIOHy9
iJXhSCBUXmHD94hwMxZkzq/BT6oH6k5yVUqot9lvCAlXHBQkkW+bVZ3uEnbvx1ek
H3GLwMrw9Iu67AotS00kGnbEE7zBVJqjnhtM71mtqtj301liTP9ONzofzzWMl9Lg
DmpVTfwK88BtZqDYtn/QkCXn5vCrEGiPnFbuTPfJvM2aFiKYcibzGGCfMd36v9u6
YB6QbEGVpa9US47Tt+93x13NBqe2oBSwVjxp9Q/bK4HB35dNsvn0uVSsUbQl965k
3FRdqhNnO5Vb+o/YQAb8T5SfEakzFdCNt/ac6fflkHp7dhaE3X7FiXfpNN77N3If
UN2vXVfefEjL3yWIC3b393+TQrFI1QTWdFjdr1XaeIx3wONBKoMMUnzlTg0FMZ4p
MI3vrDjE94od7GW4wOPYqlMGbvk3mereh3+bRYLvx/f5pmP/tShB3GKzfttwHzR5
bDIm5VcVqfc08/UCYsDWeHULe2yQY7xXTuKvtJLBg8RBpEO51nrxDIhQyKrLS+rv
WIyOTmLA/Q/PedT7a9Sq2Y4ZoOt06GhT7lYmVoYh2ZmygEi5cziY6PFvd+wA39js
0Hb1Y0ClNrHK/wR+EykHKUwB5GNlYKA9/fJuwih4YP0iDbbsStMQ1AYXf3T7GEYM
8b6QfkoF1InVzXcdy83O8BvLhbC8GlTisYYORMHOWgWGZuTW8uKlPeYg50y+opBg
TRyIK6P4s6qmcf9OM1dG9XzOugg5Ywh6WKIwOIUf2CM4Lo+v04i5vpn0qBb9pJBO
ayN2KlVPIlQv7QLI0mr8oPOE2M8yIUKBEQmToMpDusYeRuX00bExIpWBgA3ixD5D
JK8qJnQQFV3mi69GWBeY09zVyRZhntWXW8aGyR9lkQ9c5C7+W64xiCXDGX/I3PbM
YfOuf/lL+9c+lgdqO6cEVoJ+m9XLv/YdnRaw8FedM9QJuVCLt7/g+cATYLjU/aeu
+0cjjql7yCb21/XT+8CEWUs/FuKJZhc7q4ZTU0sNc7zp1uGY084oVQaRPdnvpOMR
Pil+zoDhUTrd0oRgQwAc6tFOQn/85+ubHhzhgwE2hhRunBMoJR6agRmCuBE4yEzZ
ZU1peV2ga+zIKyFFVatWtuDIjWd2BG8rmmWkGyqECEkMmPW0n9Od1vgq/vKByQyL
62Wwfd2k+R/HBdDbakJ3RdZei3+y/XgaQnmwnU/bNgSRTghIBwgMt4vqDG8S2U8Q
puo/irzCtwIow9vOGYyc8OYfwVmplhVPRxgA02R2Hb7JS+cpCnsMyM8Kn5vj38OK
cYeEj0BtBOr53tIJH2y5cD0lnNZ+Zs8TvHil7clsrcZS6ZBoaCWw4Jm1YvxihJlU
+Nbl50FPEDAzN3nHLgamtwdvg18AFKYdlHOY7KsY9La4NN5xga6cKIAOicaYCki1
qqdY19TFfoTIc4SkhvS2ndI1oavHiL7RwwPfyhwS2XnzS3zcp9kER+PvpFKlV4NU
FyYFK03NEhHrjMjsp54sSGgqBPOmcx9MQFZRa3iJ45eOh+uYujxXinl/OnqTLBiV
v6hS0FVY3ySJom7WsvgVgn+kbctAT6GfMdPYJWbRZuTsv/QAjtflOfFlRj3uOlsR
gZZcXlqe98WDY5rHoFrC9trj8Odm5yncmRFMdyjGl1Bcz52tjhROUx50/W7EtujM
i2+Xfpx8toEQaZwtK799HzIooccTBk9AMhkz9AAZTU3dBPOq2coo9G/11dtBHSZx
tYERDLGIhguEKjwBbnhL/eA/HsAPd3YVB5OVfnRi2FhlUruKZjb4SIloSUOkQ09Q
gghnWztA3wSE+tZihv7Ji8Dsb383qRoEiq6ia1/5gavumikKEjE0OZQCiKn01wjT
1BterQeBVGrciOPv50rk6vmJlQRaBKZLxZUe32kEewO/y1NrOiHV3l4m3kuEBKLc
oDQKNDvnzCOg+lFFunCt6rJIorpCmSfx3y9zJtLbR4/XHwDakrMFxJyEynTGIdDF
KlzisE25MxAWNrVKBSzoPJPmnsLaqQJKh3G5AQBk98u4N79VcgjTqmFyDSLjb/cC
WKkntYgxzAVNwsJdj8r+nrn3gMr7x3KvWDmwJRXyT64pkynbqHckDuvNxMVTjwJ9
oOMEJEtssVbgrtsIPyiBWnbkniA15kTVuBd/sm7z7XiKr1rTKCODt6a4S/xqGr+Z
K0o9eSEn4ekcRHDvk31Vt/PcyJkq7ueVERm9Ha7gEwE6HXdkyA8v0rES3SAFVGZ+
zdiOIzFTzvkmWd/yKJrgdDQLvOtAOeu1yDvKNudMue5T5KW2lCzdVKuVp2lnZhPN
Xizc0PJrwibQ54X/dsR/A73TKGgs8RPILM3Kc6sq4saHaD7haLtSb+bFjbJu2mP5
kS33yL3Sz7iTbgHMLzVCfF60oFJ3i2Qrc7MRZq7Bfyqq/ZLX+rjZYApmS3cIMLN9
OKi4jjwQSkCk00SIdtL6xWnv0oy0cL6t9rVM5mHcQFFNNSSopkGAa8wSs5eP0qG8
r8D76H/hM4iSXpLrSjsS413tkw+WfqlDyTxdRHnkwtWu6F3f3Qot1QOPV8xVblyM
3v5xqar+xRb/DVRoDXAKlyIfWKJH1RbYXzF4AoGTIJ6FIFxNWsHOdgpuAVhrsg4g
kjvLnUgOJP/hckDZaaxkjmT9E+94Y4zYkQXES5M0m0f2ZC6qXmHDEYa1SkE66KJr
538PsX3crywhHgg2xym/pxXvsCFnyl/4r7VFU4lhHOPg0uWvgXEn4PgPI1Pqv4eF
ai1l3fc05G7rub/F6gADx2008MpwePbRkLBmIg+vFRMcL+CZmk+IwUrulVV0H4rr
US8GL7Gc+0PoLlx+K+7g84jH44U9aPJRFJGvl3RKif22rjwFHdPqgcr1AYDb6Bco
L3yQqT75G0MM4pssxq7SiEA94PPsgGnfvkSXXjriuuSuLRNe0HgJ3TOC0fNMUwkY
pTwihnu70qJwqQWNSUVJkrtymnCBlm1tzdfIRyVEkOnovbR3YRqpO64kvJRj09D1
T2FwE1sI06Jl3A4GIudAqfymyMzD50Z2MllJd7ouXNuISuv/3n6eAX5SPZKuUBwJ
n/ltUHXMrZR637nSO2Vxc2zSERgNMd+rJ4V8trwSqt5mVSuU0Croo4cIM+nshiEC
kldURPRW0Bh4GnY5gyag7eSqrMavLi5t1BQUWdDeQVZKB5wia6md2nvam4evYFYt
MYKqUbCCImIhw4gFNp++Nlc9LImfkvsoM7bFkKUaGaQnfjHyNFNAVS2ihF3Mry7y
cXZj2rNHkKVMENiF6ZTCHS/djLdUCnh8otqB4rQTxGJwVAiKvU4oYS/kN3k2Sohs
CZD9yWiu+99WTgWEQeBTmSifNHUyaMcksoLz6AE4Swjf+G1uFwFuub04MGTQ9/ym
guatOy8/EW/QTX+pAqCX+7X0PAtX/M4Ej1LLPhtapDw35BgOFhBetjpRO4u8qhx3
YCnW3UsiBgCAhGF5VlPD21J/mX+hPpCyPFpLMzg8Fe5VzgPFdG7nGXjn4MR2oPnq
9wZtHM3f8hWrSIU4Pi0NjC2/W4cg2QX9pDvaiSoBd3EXL9Hb2sgJkfB+uQskMXff
6LYxAkRUfuqsi+a3rzoCS+r/+yhn3930XR1Im7HU6rnxGs4qSTO3z3IqZ25lMVug
99duRwifxEJFqSJ3rQsRFoKeDRw0WtXBMEr7PS70GnVvLCtkD6NyqnLeTtMshYnW
PUZ5fdnTFGUgNZ9h9c/NE8rCI9FwljSBy3Nb61Sj6mvIMjVnxuQXCoFWEHlP9zJZ
k2Ek2veu8jYFIEQ+iS8uInEdRoxz3wSem27wteHr28zoEgECJcikj0xepKwsX16S
Pml9j/92ztmv5OWCaxtnjvvtCTsAzuMQuiRXYn9J4fnOXdLVh5xQMK8wly38z4Uz
rYN9vEYIYLuVZlMQ47c6LZG1NaFJibDR3sScw8HRq8trcYNq4UHiKm5Jbx3vcFVL
CB9V+lAe/zvTJC+rP9btob5s3+O7kzSW0JrvbnlXhaGYQpKfihrs3u4uIeCQCFKp
t0xRI0ZU9R188BLs7vC4Fw4Uu0rukEAY/tNUicgt+Q2/eku7OMcvTV8QEsrxrmYt
yjhuwfbT8zgmrO5w2BF7wD0IdN8nGeSXz05cyw29Rm0nKYPkSu076YbhWTOfat7X
08Vb/ZpEBG31KQMZOKIF9s3ZXjap7HQ/P+68ulNOVxRLbAe0rpg2CN1IPoAg+o6e
DHR8uaMCvF60PWD+sxPgz8vaZSQmc/szUYtRb9WD21zX42Urlx/Jw+700rHVWKwb
mZxgSpd9KzzUjCJ6IAIOZm92aDNZR2OZDwthxKg+xn7XFyGe9QIh9FofR9An3FCY
KJuNJgvLvJ9KZnpJjU45Jd3XU/j53MaroaFWMeN1EC8OxQfM1zkSwuJ2NF7i27A1
CMVYmIO6N94+xnHSqi2EA1ZO1Bm0Wt/pEeaZvM6Eqa61LgvK1bwXg4ycsDu4P1Kb
bj0xyZ+quCsPD7wZ38/ZPwHMgRK6vDxCnbiavxCgPHVhMyQVQ+kqSfr+nEEhqkh6
urz7u+U5ml6EdC1IoHuvRtXwOelpERxgiLlSlqMk+l/N+uotuuR3hus4z40mhr7L
4eEeKmRnyti5GziZb0ICzMjyA+Du/uZyHFhUS09mdq/1JXcSJpIDKF2Q+lkdIEf1
qsDbUfE8+6LFzUT4O1wk9yFNXiClfbswCeu7vpwcDRwpuae62wtDFh1M5FaGaCRF
yuKJV0RZ03YQPondCYzKxaTtQfYW8W9vQBPCkpDbj4nJwL9N7JKUOhugUv7vvGtm
sbWlon09FJbijgOsVwGerXwtrIlhi3rAJwdXoR/TYAu+mgWQQP73UOZEdKMLYD/C
5yh3PD9o/BhLRLQMm3ypMrWAq5adhzfFQ+vRMqXlR1IQAb34oNuMthylolvi6ZYJ
8krLExwrionNRbQDXiuRw8jN0nGoVF9fdAb5+WlzrTZfobdrGzsQQFV57C/LJLt0
JVE1ExapRzfxmq6/7uu1tmHmYYGsZn/vBNsHvBEeRpEOVv8Irab3w3I9HSH/WoP+
JGk4O6nhLR0cid68OuS92U60rI7DyEgXRPL+YBbW6apTSzYCwYi5UZy8SKGMaucF
iwnKWIhWd33ROxSpib2jvtIKzG8g7rpe6j/fMnw3fc2q3o6lHoxOpMEqaQibKQQC
TjzbY9JxnrRrVNGazjabglsj/Mx9n1GCp+4TZvBE37mMfHQmmRVOy/JZ2uQtMnkk
pgr/rH7w/sMHFAq0+E/sM7d+z9vvUksmRxWWfen40ZkKidPvcNmtRZ4Aq38TNIvO
KJekz/YPjKWT1BOlcjJAsVW8F1/IjTYCQXjhAjajkxDdq+ZzN2GijIA9vask+nuG
w3y3DEFPURYSZGbqdxsO/HLEM3ZiGBcZ/Tcr2h+2D77W5BvM1jMigbIRvR3wEHJm
WfCXDRK+Y38/PGJqXmDWyN8AKQx0pjasupjaOOYtcHlriSwX9ML8EeL9/1crn26r
nl0Lb8LCGCoByvlVIycw0lzOoO2r5gShbpSIVyMwMn++cipidWGXyFs3cSIE3MJM
2RtWK4zVfwhBYOH1azzZawMwPq1iSWQHm+bDpfzGeUe9ebBdZAAJIgaAbwEA1oe9
T5V3TOYS6DzJGz7RUaBVXPL/QBO8pscpeiscRwvDRJeGPwfub6hOxDC7FxzbVY8u
tNjfrdHM+ihtOuW4qU/l398g6hcby575AQ5j1uU9T3PNpExA/5W1YK3eOXR33Xiq
wPGoLJ/cEu0V8WEhwjUrKUhKgBKeiZoMMZKyBW7jk98ZRzUB0mt2vZM+8vTqkroF
GDIaE2+a1EorX9h9SSMboQPU67gN6hE/pdKF6jaJHq4x8Cb5TjzOAX5cukO8+NSU
EjTF8Jgwrv5rBpYzrc2UEx0iCysWkTfRsaOfcyxmNQYXpAo2YSI4roUxZKZOaPNw
Kkt0GTTKbXqs4kFfvQk/drAd+Jb6NWJJ9Sni/V6a5dzVZj/v+FsrkDqVeE74rHa1
LdHBztZaPuKkvEbWF254ahs7pKvSvS8KgIHgwGDgggMF699bDeQzGF/6+b6OyxYg
mIDscgbBc7J83JRkCPMMaXZhizusg3a7P75KZ0pMUGNMG294m2sZiCimkG2XOmMe
QqIa+ekR6hu1LO6m42dz8OMq3lHdaHTMw6ITk1F+ylYk7uuUcF/XmBsDICJyG7Sm
Uqd1ZZxklpwAWlbcCngRL7CQ28dmg667JcIIOGYHnm9lBSdukH3T38bDaRugmaLo
dUYOMynTrbDEHx+DZCEHMs9n9sQrfWl2OcERmPn6ci8q8sVmrsJwgeVp4n7N1XBL
I+Czx0O2UbaStlnTSyxjCUEQTmF5jb3kcXNUnNBHt/PHV3hft0QFd5rr9q/na29Q
M9No/nVdhA5KK07jBOC+Pifb1jMBQ1b51zM3Mr5sdgbgST/x/PhBL9V57kYWgS4T
BNGjyGkYjOy2az9HyvDrvCcBir5G0Sg+F9zZBaEmbDIO7GHMPj9GfMAN+8QkTzN0
RfsnBrMGBfkeBAjdFd6VSTC9aECBbiWVz0IrKDV9USzI+Q3zAmu+DsxGRoOyDS3d
eNN6ZelPiukC+fwioh2f6HO/ZdLsQnHKJI19Yf7oJbTnMNBEa9WYZn4bev15tL8G
sBKbOJi4t34cMkEGeB9PTsCn9OlboCM1z5s2zUvKeqA5KPX/tn460PMwzy1Qqk3M
wWqXFOHa5uh3ZkfW5mn8ilxuaLniG2s6A2p1AZuBPPXuOLzASGKMLgMQ67/XNkff
Kmo0bg9Mfjos/lyBvk+tWT2Jc+waPibM2pO7HaAvw/7VAcmS4YbOR2izo4gNY3tq
kAbguFzUyTWReC11XFHJJ63q8IxziMLuFT3Qq2zA+MkP0XvIHFO2pi1rgTTkWjHm
CxU9tPmYj+8NPNK/SAx5zwsilf3Gi5TkVCqIexwgGcQQKheyUUyIodnWXu52Oyvi
pvquirI3ErK2rLpcLubk9ULf0K2n+mGybndx59ur2QHqSZFxzL3cdlmQA6CfD5PX
mg7ftfvhqMVtlhMdYmXKG9lKGuI2pfbckFBE0FAQ8T5vbPEw9HHMCzYgipFgtuA8
j85M1DV93fJ041EfyexXl0/P60ZMz7T0+nkJEu6srbHOn7vsTe8NupdbM7f5PT2P
RZw0CfSXt++yUKfhmoHgkc9mX2U329vGV7PCHoyn+ssiaid91V/d+DWaGKi7WQ2m
PobAITiTjT7g+4hwDVK3gPnDPFrkgEuaSTYyTXvPKj4JZnsYbunwtIJmcsEbrvv2
a9hkjUmI0lqPsZPjedhluzC1nq6Q8fYvW8AdrUkWN4QiGezS+3df+Mwi9DNEgA2i
AvVjyGwSvY0ehD3BifDtp2ReeP3AJsUA4V8RguCLX9E6sjLrDsL/4HQOS2j5lpVU
XghXawqsrS7IjRmp0DdgAGljOyOd7WAoMRe19ei8TNV23AKA/8ScFwc2C4x92Aid
InHuZqhaaAlV9xpUAWQ71S2bBLt085S3ZOHTs+iXTb6MAZJVkaCNHTogY6XP5kGH
kUeqmjw5/CtsDLvUoX/dGi5sv4/tuP5WkbkZ6raR2c7yLNRjjK8aT20CgKGVV+VF
GL+zfQa7u6QeGpEMvWeS1aQ3zNtO5+hGNr3Y3ksw8X5R9gLD3pyHm/sLU6sv6tDT
x3nh583WU///5l25peOhLbMbeKxwfP8g+JdT/KpZ95tIGF0G8igN6sk5IkdMK2P3
NBVJws0f16SkzAs202v8Sz+s6Lg14JkfNX0jJHVbfy/dQ+OnaJXU7O3qoJjuwPBW
JbKmxPjqKrOr9eg7KSDBaaAMLkL9WJan8uwoXb7ERiUXd+78sWhXLv4o0rJt2rm1
tMofJxiowCQGS2/xYYURoZpjcNzRtakqPr2VmtuAW2wtQJksVll8WuIxulTPyAm3
u5IZxyF0/lYeB+X1BbxPZQhGg0T1isXWvAb8T5PSYWzFq0WBXBpoWjUaITQIrnqE
24O+X4zYZyjI8RDrt5gBI1J/ivlK03frY4tkWX09oLQedS3Woa3PYDmgpB4FTmW+
2TyGjTpKhjiGXd7W5FihY9H3HkOYJHSrPjcNFKK7bBDmQnrZdlO5JkhsereEKJi4
ieKcmcXFexIe2TzdjPv2dZ48IkMWwNw9F2nxRFOs07wD4M5k9x/vzUHnoR9mjCJ5
tdLRP4P8IqKS5KX/AIDLWShJK63fXqLkmnR/y94mD2OT7uRr4pHZsP22ffIAWEjM
z+bBcJPtKI4eEAarZpi0IsTWg4lI7gO+NHmZHABTMGLkIuBBSXs6h0sBHmWZl1py
GW0BZRUZ8pKAJ7o71nFMEW+XUqpZoWQMqGgEoy7sk/VldaCLraiDAzVSaEa+wtrM
DFXri5m9rAR7vlEG2+drFnhK0ydQ/KJVLqsHYFCpl7MGyUQsTF0JZR9ZzQRPYd4i
zX095s++4cdDdxic50gLLPoOqj02FGfqB2w6tO4MEbfCGKjotvedm7AQsTPiyTqD
xnsZ5qMOY+Q1qVdZDXILn8hTEJMOnu/PZO3L2JuPLwNnNHs43OAaqtVHNE9mbu83
aNrUDsP4/DRaIeJepZzBsth0jZyFks2zRDljwY55nKbjcbgQe6773holDqhxlph6
7J+WYkEzTB89YI2YKc1qioHbbw9VPA8IPIN3U0uT4kzqzH6xlVYMTiYdsJ4Uxgmh
Qov85b8gyuoM+FxOr1ruk3EMjHcrZe+RTMsLGXzZJMW7sedzy5+UnTEtO/a33RYT
OCK7VE7HEQ7UHgHzL2puaP8T5TAadq7YU3FygNpZ4hrMF7KJ2iboazxGGsjj/J4n
P2eO98VE/jzQ9aoGQT+Z0ZSQ1amg4/dzb807/4no1T8EfqxUEudOKhoBnuqEfur7
1bVy1+/mxsUqWKu7fqFor0T4Gb2uSQwA6MyR7OuudAQV4/dcQfxcMPtdMb/96igt
Zfj8/VgoveYn26npnFgR85QKWx8Z7D7ALMFPvld3X7HKRTqPB2X1ngV3myrr9E9y
OM1mvNEanemVFh2LJ+MRwMUf4OZWg67NoFcziVlDf3zJVgdXTI5FUugM/ohshjZw
ABC8rkl+e42p5FmQIQO77f3ZZwsT1BX4sHJmlvQ3gH7oQ/8Y0fy51YJfvEmN6FM1
bpPK9FNSVDuxT1QhHIa3aSuHY42dRMQHpS/S05yFAWc=
`pragma protect end_protected
