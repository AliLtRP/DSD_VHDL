// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:28 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QUjaKkY9yhfwSgLLxbA49ZxRczajatvc7tHOMRz0n49T4Ev61RpXk/wozS3//kRA
TUWvTic8BfXusHK3rrSXgy4vSEFy9kgs/xkjb19ZMzeCzsDulM8Ydy5LUs6k1GpN
bE6EEqMs7bjvayTR1X78wNp4EAa1rzMO89qZcKYg2YA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19904)
IyfCsLLp6LSWMtL+M53irh+S6rSKw3Fs457/67ZA/exH6/VBLHyDbiYe/moZgiWW
lL4WVTNAtPe7SLuNwdk5n7doqueuaPnnsJPSUDy98gFxvfynu/arK1dWzM2IVCN3
CvVbnzzaj/mMwB/4nlIZYAPzElAlzezMW9ZPu/gGPHw1V22zM+KGeFTj24xHHKNH
S/A5h/aU63iotk9NB0UwksZOPiAp5i/gbm2R+yAqIk6XtEJOI3dXmKmQNDnr544V
tZgbYwEiJ4Ujre/lWwhwW45KElrnZlqNu3k8yoE7EjOF8kpQpqIwJGdIPYZHPsYt
N0B5OiGAVhisCyO2CKl3shNHKkgYausvbh2qej6jDP++bCWPUJ5EL9GyGRiVE28t
5IW73fFuHCrsEDiod0DhHCPY8ByPhSKc//v0KOwSZOQPWzHvgLaP+Y9WaLPPWynH
mUAf3IQmUZ7nMnfgRQ8N+e+Z1tOPOa38P1n9RGyhrDLWnBTId41qNVn9wmYgwlj2
YDw7/h2TEX9Q7auGAXwjz4dT+G1Aetv5w1spASqBUeuQgK55Vouz4tQAXFsmnRD1
Di7XP7vTxUgh3DCZRmEp+5/kFv+im82e/6mf+YaZxk/pqzEapXjgePwFEfiS32IL
BaUEqWM3vUqBKpAzNPJzGSSHl/i94l9x4YSC2lxlufQsOITC5KI2SJGHS0A4HRsy
m13NlmbosshnRyI2akh+IU6/pRSn2Di9ruEe0MXglHTZ2xnEvSh0sRNdZiS8Q9D1
KDpIsYyZDn9CXcgUAXgKFVon9cvzy9yEIqL6RkKOxAu4RIRuablMPWG4TLCTe8u1
Ftcy5D7GwsWEPDNsObtQpNw9QrRjaMpTSgqqGDfRURl64SSSFwweN2rmE0LfPz52
lHJ4jkfBE4hPgSW51WzpnNNCXO25GULbIuhaqiPnJBbzq42t0Kp7xNopdWmuICgu
16ImD/EAGFALTiYMzT2iD9T6mjVR3nLjwzsd7swUsEuWYgi9QIlnOwg6SwRjz4nQ
hu7Pey1hMosOyS6TMliUjB6fdfAr8X4SComcm47HTK5r9J1ylyihE4Bb1jqhh0mg
BaPlwnIl7EcUFw6HznyP6gqTvkYEkz2Fj0qOMcQTyAqiciAl2xbEs5cZdXuI0VAQ
nO86Ddd91NiUi4HFKCts2HkurcLQnReo08p+s2ruDWseeqDmQGtw2V2A65tCMul4
hEFSbfB/stRmw2zUdChNg61rJN5e/qhMQzgNNnA0mkBgXz61ixb88NvuGcJuRH4w
Vf7hMcx5yhzfA8octt4qW8HsbsOwTInOwlG8vRxxnIF1LBI9Y3jnwwI+ImHWmwgl
1x2lUsVWY6Kr6YV4FIBUi6ubNNC+/EDpVfvDYLnlnoX4/dTyA85pE6CNP0PI71Md
YRZnAsj/BQC8tcLE0HoSdX8b3jIK0n28OmzuyxzI8hlacz0bF8vd2WPOX4BP+AYR
jzWVIVmLdMBQ/unxoLeOB+NRqMO4PksbExKRQMbJrGqOPzNn1QkTKbopeOMFZMNY
vWDtcCQh02qzp39yY95ENqn4lDrMyG+pJKcULIwcBZKoSp/wR3sEQwUrlB/s+8Gx
NGnxFwc3PIxD9yRJCxfBx8qqVOJWNs+4FdbKyDbxtzFmJye6c07tV4shK6Udx+BF
bwmL6g7nCgE3qWX5WdJ08537g0IswIVyywK2227II4VaOjK9ZQ9oFX80FE8PUc7x
PKmHTq4QKnUGmD+SlH7NeCTmAT7CdgSy3kKAUlD9DYd8TxFPHsm1eCXN/URSFJk6
r5UG6RqK5QgRiuZpDqySficSgBXRqFbrxfqm+bA26z/apnRaWm9dAFlcs0OxAwEG
AWI31FxaJ9Ydq/8vlrSd9Zu0Fn73WuTRKJ3MX7C054x0XgELn9WEzJpDaswAuKa6
6VckkmpsCZj6H4tEkgtlaV6/xMhGk9KSUFEeE8FKtfQiOGI58FxdChi2xw3tELjT
eUBDIEYGGXh6Nwil4OTgF2rFBSpg3z1u6z3BqG2bLOmAY2tUaDWAh2oc2WHFziHS
SaCivxs/mARe8LR+eH+pEFvke27+pRSm7Ulzv1z4HEZdXi8i3JVicCxmy3taKVHM
02P0LuapRrXA6oO1w6LKekXGNuutt1xrNTcyuDtVy++LgbUcqcNTzUx1uy/Twkl0
sXaTffyQz/bsVjBU2TRPdhQ+SBQBBc7Jzlx1fFsKPzWFkUJtG0InR3saxJIwjdRw
yU8EfuWxdlzhbmjJXjw24Xhpztj20rkAXI9sxs8y8irX4o/DvDIAOHDIbCWnOUk9
/a5rYaOsqFxZ1GH27sAH+DE6XLOb69iiX3GaNGSsWBMx4Gi9yOCqouc7bf5/cr9a
VqHUoxGdK28oSGa7/TcqbnSHqlx0r4KKmS9G3vlbXCuHoN+pt4X+E/6C0KWgZDez
IFo7tqUSuQFzFt7ZWFsuTS9OQaa75BQOsv/LUeUyaxR+K45bLoRHY/onc99ipdo+
1eFTRybyqx7LHMabeQQ4qZ0di8r4FGff0oossBKyI7WP36fvOkq/42mDFQ8E2tTl
g6VV0ZYAiiSUIqBrXo0jTxTTYxb+fHb5lSJfdyy74fqU/F5FXIOgidzvMA2nSPCn
pUPDUajIs/PzEpDei8Nk8Q9lwk3oP/jQWBj+azAg5fFvhpJMahZ6bLP3W0YT2jCp
YW8EbukTN3jPxyjaDMxutpdMhbHR7c5c0rvv0UdzwtOODgle+YsM62gD99lcVZvf
H2SucvZphV4gnsI9SYp3JlG355KpcCbhO9iU9TPMMpC08S1YzVQJ7cE59OrXbZpS
x5/fqfuXXdYM93EbR0ExTUHrHxvIbgFCXIZVzp2ow3i1gehx9GlDznSOZ6AGdEvZ
3uGzMHD/dmU2/+l3+ti/GXArtzlMi5xiIUTpNiW4NZeiZdy67aZabNwQUHvPds8n
2qJ3LEfbfWJ2vEZzQY7DQk+mnMl4PqQheyCTBbSMQ3Xy9Xm91R3Q+sILHvRjkL3Q
HDBICI/e+nORk9B8StB/cwnWsdYJoT/vDnX3QNIcb5Yj1fWgW/diWNDEGijgRXn1
9XI6UL5BWNaWMOEm0Bn2wMZpJvetD0tHZKrMDaosD78JOoUiGy6IgdKE1CE3owyn
VSIzdrt/Mrb3wxa3AqyZDhKahKvlILFQNKXokUyezjygSsraqgJsQPUq58kuYjCy
fLJn6Hrfy4mDrBUwKs9tzKGj5CILVkTviLmIGO93owVwBTj7auelozuZUEfbv7My
Ip6lfwzAG1u+tIwQeF7pGcY9us0wVBktUYhYAChc2cmTcaxTW0+iKKYvBWhb134b
BN4Qabl99Bmmreko01Q2NjL+SwrMGpKx8DfaI4FVZ3L48eD9i/76zt0w+2/Dhq22
6XXOtQxDuIdqu00jxZCst03YMktJz6rArMa86HVNy/6hK/KdGl/js/WG4HtWo90n
uQ2iJ0Tvcbn0S3TErO2yyfWWgjWIO7Fgxsfn0ZAVEiwGGnyROMQHpCkFPARFWepH
SlYOy8flaG9b0G+M9P3PR+BlYk42MecGPv0jJ/1eQdvp/yAd0VmumxrzS+2bSpRV
UalwcWBzcin8HxZWxgLdIAm0NQlorKj80Bs6Gsq1IHzPpletH/+FhqbbgFHirK2A
KPbrxW3UtU/YhX2IdR19Yktn9zOw2MWlPI0TLETwJwWk43Mg92RT59OlOl3T8i8a
ci2jVLzqzWVvMDHb7jBDu4EucBwFGGa16vG2gQP2rG6gQoV32R5N8titGNE396Zh
p6BgsFR+3fGo7YGdOSnvuMbA3Cu6mw/0GpDDKRm3THKWv288jiUTYd6ZqKLrMwzU
ZJb4Gz5/37/DhEVciWpspPF3RLg23QYKsTXL6aKUCvtjzyJJY3z/foMBM4GM2aLm
qDPBEHa0EUm1fc606uTj+pjl43BiibdSsRpB9/wFAh29ilh2oYIqNuFwHIlsaoXI
e0WCtRnSqgYRPnKDO39w5+y6ZC45rlQMlLqqjV1XrOXvjSF07JELueJjBCOQq8FU
AeVgl/Mtg+JTl7BaohkTrTJbaLh6lUKDbpCSW6Pso4fdHKCHYIqEwPyUlSA6mQJS
NKFEmRcs6RWWXhIzC63Q4v6KDF9tNaFkP4inDp06ZerYcw4gURqn78k/3XPbI1eT
BkJo+4lazAat8GfrMJPOcxVj0c1faHx5pigw//ffYryzAUX5czJK0ijNhHgbvREW
eEyfhjfIEMOHccSHV60sBbzziVXlrv8I9gPFx/cNm9ZOk6CdcKIYnIdU3Z2uDUqA
CGSe8yjbxCap+jqKmQGywOI9/WFeYE6XcDLv+etrJYNDJ+WsDNfduRGIzG5bW/b+
hp/ul2Cl6J5+HthT13FXl2W2od8qUeKt7jiUO4qpW99tq2u4j6ZHPVcoDExL88ct
ZKzxZl4Co/GzxhedHUtYEoNESZH4vxeM9BtpU0cuawZMwQGCUnEMvDqpGVVY9vQN
CCY2276vsu+YhEoI5YyaD/vDohH+/hM2MFxJdlVklWNRiWiKIrPJjNDm+tv27wfO
Y1xiADRu/TFlleXF/B2erMNRh7AXG5bI4HJ85TJLMTY4tMoVvG3Yjfnt3/1N39qV
sZYSWAMGqb0obobV0+yBvdN+lvbMYGwTfc/fhhAD+W2t3s+iyYXHc5rlVRLRTZcD
M2XkZ6jxn1jffTv1zsT43wHnKcUjhbAOMrzqJMH9uX22BezI21ZTHwCGo0nPDCe8
CjZbsdUW+X0CGHPEYmnA/LXAHqwEEycFpoYj7PMQV5eZaIJ1sNtP66VyJPfsPPuE
008ogYYU5VixlkKvoER75eRmGnHHwo2g3IOES3StMpJpNSpNsp5g0cWTszK3l+L+
+dYEMT5+qeA4aYCSq2HZsnFQEDL90H98uSbOTKPhfKYVxxakKQ/OVJPJxJ6rLEXu
Cnvmhmh+zpN6RwVms2wQaTh5pYHR/BieILN7dj2YzwlFqwvyHcqnj6gKKS9c1Psm
BRLTnVCo0YdPhUkOxnQRnI0WP3qKEsc/bve83V1cz7hjFNhq2dBh3N4aLNBfdcpg
tt2ajWWw8f3NC+Pk2RDaA7xhQzx+nSOKhjqemsFwkhEfuuCiGlC4m1ELa+b5McSu
63sM0V5vmrV9AG0AWKX+wJuefvEWnV8dPqQzRGVgo1P1T/prLASvP1IXSMlcshh2
JenCgw2J2j+5NZJLELhmmOScNo+Y+SWHIj7ldl9zWarGXXZX6QQKezRmpTNPEyCY
0oKQfWHdVSp819DPdenALpBcwJTdHFdh4tLYdesxtzPzhSPoBMPKi7fMR9FSI/8e
153LqB0hQ8oMoWYV/VHndioviabQwk8v6er1Xs70nr8wbiQq+30aM9aYHhUX96md
N35SC/lpNmgwZFmUC1om1hSEtLjcgIS8TuA4gu4+HEIby3TZSVAbnxBQ1WKIZU5C
wasHqfSiBzihssBkZ3qSRo6/c6tIVPQHpkm5wa3Iz0B+wrduLrmuz9kjEep9Z3Tm
Y3LWCK6ZxC9peMnB7HxVXPeA3QosIT2xUgSR7cngAKhWmRGUnu+Z99/tGnoS7uid
On/V9bV0xp+nLd+skVwkiXaoSaOvBEWr/jr0l49qpcq+Burmk7zpAGs+5uADzp0k
M3mcbMRk+B1VJoMp6UWmoG28qtDa6mZ2bPG59FUqtHGzsmNFCkfmmHjatQ6r9yEm
ksvEWf750MRnmUelUKYTqQMbTsAAUh5FXmOGburXtWsrPVsRrt3uu9jG2CRPq2lV
SpcdaPBD/835pHNg1tEgYvWJFVXiVREBwQZi5HemYQDca8Gxw3BfUf+W9dG1knuY
QZBDXHQMsx/QgJlmIORi1tymi3FLNzx9mY4crvc656jC25CbBSB3FK1mcVal+U2G
5C0VMC9mkL6VxUUdWYcaNYdCSsMaylyQe7XSYPQn3trcA6pB14ZFGnT2Vqxm4VAD
SryYaXYBVof4VvJ3kYuTZpN1H0KwAXPHTd5Ar7ZDrqUnQXJPiT9thAWpazj8vmJT
PzP84ttcqx0AYTIrn8mnYxlNt1psBOlDBqIOYnxtz7FZ45q/mUhHZ82dtH8c6eI5
6SMGSX2fqynxPiLMvMT9qxyblpwq37WoXfBSaDuwGYw50TH9vLxtcDPZVqcqMonI
EXI+sNLEcEzOVmNTNtJrXCYndoPCg4J7wP7h+AC0s04MGDP1UaXkz7OLsL5HrcI3
vBodQ54vNrA+83BmfRUAkBpjcHEOLH+vpmNMkRJjKwxHi7BFy4zeIEHIyR+nBHlr
XvdUnJ7M1eAgyePZdH/8Oo83ZwWvj6Y/EjQ+TkXT9yM+GLi7TORoqV+SFfXTCD3T
ZeJZp9sl4ZLO01Stihh7M85xgCRCbp50xbfoW96N/reZ7o47C/4uw/kzhDNTTUnw
HDL8svUhEnS2Ldi46y5e3AiBwG4EJijgfFjeB8kRmMekqs3DmvVlZj1FnUhbPzA1
A6mIRE9e2ERbw2zOFN35LvdjRxyzuANSGvKMNu4JxuskZzkcGBAHJEbYuZEfhY77
hl3ofqtwhuUzpbgxyw58nQGF5OO8VTDAxiSevu9pBvqw+sFjFqowoZrVhxpm5KN5
WULw+sInetd3GWb0uH0xesaGoVMyVJVKkME+SLwWommEe0N0LOy7KR4sQ3Kdxybk
kssgFFW0iTtNBQNd3X5sSOvNjA6JgrAqqZEdrYOGh5MG4X065ZoqtBo+XN3dQPOc
muhRzpYuEZx4IcggHBcQP0sCqbsyot1O8nv4U3lpfqp5/KXinxKXQKDM9qFvvEWN
HlKluD/XyVstQa8inGrDO9icnujVepLZl8tLwCUfkHWM1lc8KnOYqBHCSGf+pwKd
83l/9V9K/cKa3EmCqQOENmiEqHhUuF3MgD5VSVoaQ0IneMZ3Q5J3rk0WZazteKPE
pst+VmWmbuaOjrnCmvRZxQQ/YWzYPUBkmJhZyNew+H63ZrXxwx0XFLEys8cMotTd
bkvn7wlbYMI1ojJ31ZM47d6gjPe+lNYJO6NantBfnjoQz1XcIpcaTY/27tp1n+mr
IAx2mUxjRBINmNZihH+oIPqe0p4+yDUoIyCcXZ6KvHe/YfMGqnXoY7tMJuYVabYm
br9MbiHZKuHqoSZkIMRe9QXdGmrS6QzMTKDyBYxfXuBzmZiVbfbmwC5dM03ABDdk
6zj9viHXddud+1trbpArZOF9i5pBlJ9BTjlZ4ynrSvi11JWqVE94g3U+LNVyyun2
hyhPpbOhTlrujxIO3SQKRdTDH/89p84LrR4YiBa4hG++e0YQmSGvWL5lTCnqdC16
5MCvmrnUrIRrbAaaVOAmOrqbbrL6mrEOmRaK96ozsFuOBzVhigl8HDU9pkb1v0xv
+xyaX9S6LWM3IkuJG2+02jltVa0yYJj70bfHQkIlbgfNtJbnomD41txTAOG5vupb
StaOmYImmak9TBHg7RvYL3+8y3BzYCDJaek9IehxlMHtkyGz6SbeSLcvDIUAVKiS
D9jnF+Y4gNTmHDAfbvd6dwPGT5CK8Yj+EVI1Zfdr60aTxN28zGC8cFVvSyA5FrLt
qdruEKQ+Fh/qhwn8nRi2yRqOqZ6ZkZOuj/P2NOEpuoXiqcuU6IkA3GP/PcK4Kqxb
tudHyJsrvIyYY/RTut+O2t2ej3YTGq5OMNzhcONAYezOnPBp81xetIA+6H3nT1Qx
7xNod3nzkb6BA9dAHp1H9F6YbWWSptM5p9Wfs7t+J++fm54ljuU37zZ74XAsHMV5
0d/bUEM2iiMo0xY2FyPotb9WnD8UmdTBHbiHr3W9cTM7bbsd65fJHLSuTYf7m1qW
QRY1NvkVFhGmCFiMLFbcyiEehqcm89qdP+D6ZaclaEm2Hh3wyXMm5JcqXxxNFe1a
3b02DgRwY8bCMsVQ1bE91rmsOKikWJX5KoMZpBQEVXUwMHk+YZkALe8Nx7HjMvdS
as5Hhpyo33EAoPekOjy1eTqDN/ITpOXZGw4vmyjj9iNL/+hCtQ3EpPSDMDU347Bd
p/lZ3wS54PMWqYi+ugecteepAeoWoB+hqA8sBSUH+Rv8lwzKP8WTVrLUoADOZ3p9
HzIOeVi+EGIOXQpbZFoPSjLQMzmn4HC3QBZ8Ki215Ze4zSkxFfKKIByIRcugP+GQ
frmKyHJ2LA/PfKVSu4vS5PT/bUmevgXzAjgeasC37MyV4LgYq2wbfB7R+hbBLOjh
acInsOT0hTtIEy/hdniJj5cN2NU4mhtOevtNkvrZQyTHRXrbziUEpDvahTkV8079
/WMxUlxSeVFIKu/6dY+ke/3R502aD0uZ625yESYarkB6SyzD8KRNGnq4L8KdPoCD
ZS+hwapIvusPR3RsOrtJBEy4qEecRqe4UNf5/hUoYUH/NkfZAweB1TAs+RQ0x+Um
a5515rSOrGvDvkiZjASF+oz/2ZA8zMm5NAe8WlAZTNlm7CVrZmlxqngzhNSqGUvo
yYWYbimFeFdTfPq5nxrYgBx0mUD73yiI71AVexxEoV6d/++zL8MqIz+zOk+bbPgr
/BgCB1C/UpkDkmPWxBfpLuEXv+vwdkJWHd3Vl0L19R6a4Ul5LsiENlB3yhcqbPJx
s3MwE33LQx5QP9rbg0gNjyirO+usSgUxH3vHl9ENGnS5D9RVk5vvejancK8f1yYa
qSYJuO1sYNNoGO4TWbFn3tymm/y4p6k/T+E/PDLHbGAGQ9OCKcVPcO288AzpeOEQ
PM9Nd+A8TtDxQbueRtGoLzf7bHwyeTMfdzBLBystyCoPawmdlWSTAphYFqrNYufv
35O8RFqhuCD/3EY5i7kRI/DmWiijIVOutYmacOs2jv2hWC8sb3OqUvjmhaBg/Avo
68wdMC/NG1532jcHupohDpMqMf7FWiTzEexld0IHq68sJCUUbCsc756hjq6mNfjp
spJNNW9AEuC2IS4RYF7rQKcOtOggmYPohh4B/qO6vu6TJPIIy9RoPVJRppRqtNTK
GaQ2Km3zM/x+MlK5MeWijK/M9ZuWln5GGsrNoirA+94RcmcejbCuU19ocCC2OWM8
pvZFbmkhs9Nc7O6eRPaLVmauJMEfvkz7ww3jSKCF4L1eyvxi5XPdRvP9GapBH4Sc
MuCsN4H0+D0FmmEPJHPqYfhuZgd7jBmhvn1Y0oeo79ht0FxlEW57pIvHZxBoXCjx
3BH8dIMhWWN15/FfiM/aZ2zRFRjdcsEt9duCAdizmSAdFi3knRl4XeU6uqC6d0x6
BLqZoMVqHJey5WONwWg8ef3F+MxYe66I2Hydz/q3qe66Zphq+5gO4uKynMJh94FL
32gjSuhw+Op9SujrHmNqTc1WdRaN+Y151iTL9ySPjFzT/LJodJn8cyBmVyCAZhST
Nsmg+o/rI1K0/MkZQlx/h1gHtk1I46r+javlBes0w1VjvECnGUkwXEc1TeaKd7bD
nZYui5k39r3XIG7pHQ40NXMCqoIUQOFp/96qn7YHhD2JD97pdBBVZxzMpjr1yDHa
mGvjgEAfPeYH1BQai3pw3Eeu9dQsX4S2PLsrU38RBxbKaaj9zA63i9oxwLWlkeqK
f0pWb+DXP89H+y8KZ5GDxThRGIlB20B+W0lJGu65vmGm66pmSskERLBXacLTvNKc
5kp5Dndl4pwZK4kSg3QpCZaQyxUQI1kSV//kfLUDFLiOc9GaRrCfbWUUNVJiJjAI
mxlq5rJ3kV2773LaBcqlU07N22sVMUDgtZ7akXOaObCyNTlgEAGGlcvkc8fud9GK
JglthZOFpc9Rf9tcdtvyKR9aKPS8nkgUzeRJZ12ieFa8RBvDLk1bP/X0JCECy5EN
AUgBF3kIGrMgkcaxlY0WgUwtuswZwusP4/3EuijysK4rsqdx+3v4Xt9QD15BFHUx
3J1Q0dG9fWkTnu/jNYCRKB2dnrWHEIiN2F5BUOZW6gc7xVAhr+uYeIxyFLtAgDgp
yUwe4nhkK7xIcjo+brIHOVS6xR1Xb5gOhIswm+y6TDk+ueu8S6VpxZUwPUkFVK1T
e9tzJDTsfKSwPjHM1OaFtbPxUShGcpaU7ffOQpMq18KHp5xykZzpDOHRntNLutbd
ylk8L7oxHWmk3iqBULVlaRoxiShPa2sVUxHpSkwzTwCg0N6p8GUz8eqvKtzrJPv5
v7sHF+Z3CgcZ+3+jjuingxqEpbWEQt9EihZT8wdYcV+n+ILW9PY9j4okJIme+f0F
FKIl8M+go0XnwcgChGKdTFyWHCoKYuWsDWYl4SFxASVwfIRuRGKkPpGD9z0yMgay
ig41iDNf0s7gqnSSIbup7gXvUzKT2KGIawcnJQ+qFNQDqT/0iuHQl1MEpN9Ip3dJ
BK0NoVeVIu2HLjZmZgWerZT8UOK6ILxRX2mE+AT6rZpy5+9DU64SDkVkRn0P6p2T
RzZ9NMhnfuEEtsqGUdtvastwu4Z96A4k2WVtoV2YxHRilSDUPs/YK3027CdOywGC
wzhhPejmE5TdsvvpCuflahvc6q+BafuvQem/JX0bdx5wqS3mOwMBkz+UOOq3STdd
0fP5jpwkkfCwpYD3QkmQeVeUSTspEVmlK6YUsdxzdOsSZT6dxq8YBx+dqEDzb0//
aajQvp6HH/cKUlOTHH+LouyFl1ruSKlDlFxTKAu2I6SRzlpNIDyZ4WFjPzGEoQ1x
/kiEg5OJhsRC/WlxU+tpX4a4bVGupHMp+MTKW0PPLiKKe+qG4pEuz4SDeNJaVFO7
eDnWY0kim/NZ4GFNaNwgbEZd813Cd+a5BHKJnLKf1Fy1WkXoNwc9d9PtQnmfuqZl
MAxPeqCDodsBgDpF5Eh+oabjozv3mmssX78aiOwJz5kFlVpuOLpMox1WNpeHvjgr
B3KzTPVZ5Wvf0wM0/xY8/bAOHMZeC2+7V4KxrJ25xH2w2lM3PfHAYqZLyQdkc3ox
wxg5z2wGPTzh84svTla+P9VrZx23BKSNFTbCqsee+DigcjSmaGrma5ELK4limtuh
CTOfsHcY37ZqmGV3dGectasL8a/73swvY+TmcA9n1IBFx/RMnM/2Lut+YQsdjkr9
52ujciDcfbVFJeHooCFt2k0iV6oGgiVfdTsS0u4Pq36Tag/P5AR1cnMsygoZBwOs
a1RqirkOSKsUzChwd5Mcw5Ob7Sp+J7C7L1ArSRpRlITh9moDZCfpsgY8ReAFkLUU
WbYy6DApYVqKwZF30JrFUokXSWxIpma4sIPfyXR2LGwnsuDqMePgq/+olbrbOaWd
vxd+ScsPNV9VqYcfm8jcTOyTlirWlIzG7fUcd5WwZ6C+LZMyoEBazA+qB9bJGoRd
8WaRx46SU6VyGFlGEiqEZyTteIcwBNnpC24Nq27m77MMfr0BnkyYO31GrNv1qEbs
TzPmuxMIiGseJRXZB/Xz5oVUhiofECyB9qdCDHSUu7eP91EpfkpTh8IdK1CtADfB
XH+HrnISiRRjxV7Zoc087I4kuLR8hxey487anEoRjY/NfuTFMU0uXP2F4FuhpbBL
xBxjWYCYkB+VL+ZAIROgxeLCwRUDBjR/XafPI03oC310bxr9Hv71jbhuj1HczZ5L
2Y1nh9pnZ1cI1tuVtMaVc/RMfg5qZTca8B5xfRWdFu2Ev994wgd4LADRaGgE/kWM
S1HPM4aBJy5cjb2AD7SM4LmIf4wUr+KNLemncoWv/jBWt8Ok/PVHVa+hr2bqdzSA
VptgRC2tMEvbNg60a22mU9cd43Z8gu6qh9ctir5LjaarwD58hXtIqfebCelUnDjy
MLjXr61Oku7tgkFBzNMwuGv8MwagcekceNJfXCI9TDdH38yQQbELKMisVPoneD4R
8MWqot4cPqL/evZAnyrQTM/kyyr6BxFCQ+M4pmfok5ILApg9u+N5NBUheRiG++U0
dFDn3ohS4AVOzs2T1YZcpx+k9paHFIoNfNNePmMNWaUg1ByaGv6lv0yGWVX7UsJL
s6Nk6c0ahs9SjBQKqa4vjB9Mx5CnqLtJjbxeVpk0iwbE2uPn9/erhRSPsWG98ngn
ty+6mAkBg6ZMW/PmSrJ2mHd8cLY7wOCGlZgglaDkzHzTrVRxL+RX7pzB7TkK3nI9
6qMgHfRwjRaFvfIAEmixJ0+iBjMAHgxceu8n6zPZ0OvCEYcptbYBJgU4shkQe5ng
s1Zi2IqqwGKJqGyu0yLlzIy4I5zOjuaqpYKlzoIe0+hLnrvJGPuvDLvsTQNt3i4t
FZl107VBM/fYj0WdNj2myFaZ167R8IyUb/xv0o2NjiBvUTtT4Fur8T1z5bmxdhK1
U6gZQNMuMh4pzUZgha8OaJHjW5lT5cQZOSf+6xFXKhuI99Hrfld4bfXAtIDDA0ws
BbdmJ14f7BkPuZIIPoe7WPchpJqyGChkHmsXRg7Qdf7NqUwlZwiiL7SmlipXfeKz
fbu6/65ChXNvs4Bdx9W7T5zQ8ElpZuTllZdQkmpPzQ0XWeWzmmMnTgQ3UQG6qO3X
AK62n+trDTTK0m76OcYacUT8seUfqhfGKhs9iSpTlhOHmshReo4m17u6HmEt7mwP
cO6W9wEAKokr1sta8lh71b7O79M4AyY+lA4UPzlvOCsdf9M5ZCAMMokgQYAWlQa1
F2PiDNPPk0JUvhdfgEGJ3yfr5CtMpR1hfh2rNS7drA/ZYIIqK/VOl2xqWFjKkRmW
qeji5HW8lYmCr43dx26iZn7SAjkzJJci8ea/nWqNnqjiHcgk/nqNmuuea0i8oX9U
JaBlFlic1MzOG96oBSKukMU5/+WT4Vi08btGAoIeNdmIkQ5VDd00PrdeOA0Pds4r
iIsn55tSkpy2OOGgkNtKTlCmb1D7VjN3anb5qoYOWHaDKfwoQ0kqzhNAqy0S/cM4
TK+ZlW5TEwitFGIG+Wi2/bkkJeeINr4ID7hEF/gFuxQ/ULpkBT6yFV0MV9ht6lyQ
96oO3Hc1gQDarX25orjy5QAt8GtfO8y7fwWZlfwcKco1DtYFlM40gSN7nhNcgU2B
Ko37rJuza2nIFQc91XhCGIZ5BLD+zMywGXacGUcxG2897Iut+YC9ozmeSU+Lh6hP
gvAQeomOjRO11/eUh3jN+hJuidkh7x1Gh6dvFgPgOKlgS3R9XMhmCIe7BZWx1XNQ
vYXPP+9aI6jS5c2L2PJ70s6YZO09Ms7HVKtAbCaVUGmZ8aTE3DaY3ewUGGSiitpz
fQmssm9e1/T6YFj6JQoarsS7ebxA2gTJolGqxxY/SIozlI2+sdJApKt6pQaTegUh
FFhPMSCuA302unoiJX1/d5TdsaIWlnJkquSJUPie9OiGTf7JVubp5AYZjrT3EXeI
0fz1jKjdwpjVqofGufSeGMTX6vU4oM3PCk+uLIMe7flk7zuGofG/zC3C51h12Yng
lWaIik/8PfOpN1SQJ7KutZ5LmpsxFnIJMhaP0UqRCjbJ6Ybjc4F231+nxScLW0yy
1IKVioncKpdU0xTCL42Zxq+GTcimCrhsEVwK9fpiW+IKi16Nrog0gPOpgoFvpOQA
1nuHQqBJnamIkZ0U+PmKS0TNvAxt9IRjWZbgoqSAiGinLBXpCSye5XTspfOkn4E0
3vH3NSa35Y7cmoFNjAQ1uK/qNfOqxduko3stkEFtw7VeM8xtn62QmRkTMWql/YJK
pxOuON3OXuqeVpBwmiWVekF0YVZAwD8K9mTdOh119pZiKWOyKpy01YqmkItSPju5
q1UfEf2x+uS2UamDr0zTREH7cQNNgvvx28cBj6FoGBWky05Lg4h8D7RL4ST1AAKE
t72UX/2/6hpFrgQbBkKUFhpgYA3wdoMUXc1fVdqoW3LG/zEUNjdU8q/kSDa/qoYz
6DYpkVdbpqdVLH0Q+mE4d0R0VUFDc/bJ4sKYr6jKsOW8V0JeMgjJvH8Kvxq0pRak
aIGYMCRPFj41l0gP/LBYb7g2oj8BKVpScGzP99ix8KADNihKiqiox+ceaSuXw/HZ
mAlRb4YxlkTqnzGfjPjJCTWjyfhlNpWASscdLye1S13uyy0rMeVdS22MwW2L19li
IM4QAgk8sXaVGPfwooBdEf57KF8sMe2GhuOh6mrsO0FJdWJvDz4z5nuC0Uy5rl3W
rR+FyCg7G/wAkVVlkdBI7OhkPMTgn3wwFlfNZvjBGzqKWUof8SU2TCJNtry0LUx0
Bgf+TyHcV/n0NwWEMjGtnOO3rMmJmyPFmxLJSNpTH/zWJT63xPnhqyBnr5YxejZh
0/rnDG8hzwVYb4NPfaMHxjc24WQFlARUUZ9X0ihK31lLGtPYB4BQjG/nPX5/ZbtW
pQh7V4nmoZ0K1dH0kZer6p+bjWChHlkvKGqNWFN0X9o9o7u07Vx2DYtLOOMmdnG/
i0Uqu2DEFIStBdEu/QdW9omNJpPm1MDqnS14yKs0KQvptawHtF+zU5RIXihZ+mVR
fquLNuYLomE67Jt4cKrhgMQ9+uWXHMBJCGjQCxZIo9cuk+QSz9fdT8lqG6jBiXNi
yiIinSrGAniKgSx5Q2bhRaDjHN2N8kRWJaSHWQ3x/wQ3nyau4b5dCnHa3zQlQyut
Lzbyk5gKLb+qfS/0rshFE/53tC/4Qta+vsUe5GRp7yFV7IhiA75UFOOjCbuLnQZf
WnWhcMtRMXnKP2e4iV3b6Cf3dZ0Lr2NDYJPb//O9cv/dcxsJl9LWwJxmScuBVdhF
7M96BXbgDZfiWS7e+I94fW41Jkz3ArK6gi/rFMJhPvUvX6oloHXMvrbp6JGlWAqj
HQjBf58pKdvMf5bpgzuetiR/z/QEeksLri4ZtsmwYDrR/gSW2oOCjmTv7KraPIna
kWzVLj43Cg4oVYFuCDa8Fl6e9zF7peZquA2+30DODkgpb0ZZaynE8mF+sJjaabFN
myhos0qRqbQZrSMM/FKNn4dlLPz/R6pYl5RLL6GDVxENvfJXU0/37nmUNcYx0H26
Nql5mZkX1/dDewp0z2/5wh5Mo3tPDfJLIQZpd5KTxNh+nsfaKjwzUIcYwtXTvO/D
V1XMJ9rOlLnH0t7X297XVnFKxcW/+L5ey821ovm2FjeFK15auCLIPx/kBPXO/wfn
CZSeI7BQ3Q2RSY2kwkuWjs0XCTMlQc0tCfPkU0KrmSfcIlxWV/sYGooOdxjOBvOc
aQOg1qY2cGV15vKfXmt6qzOBlP+vJgI5m1nxG0Y2nRnRfTdxUjIBjEFG9jkNcwI5
4fx0gLDIDZePp0CZhaSdyV/iePL3o+Anb7k8JPsWXUxh7+UXGEW7jHPtz5slEt5X
lMrdsJtu5UPizY/5An6Y49aytzqAgwW93uWz8xJQxBgZzo1BSMwMSp2bAnlmOeU1
XP8YVhaK1sRoMFC9RjC4ECt7MM4U0sKwaiqXVeWiruGe5P6zX1hB/ew0RCfHcDHo
KCaEIK8PzsHpO7wWP3twxQm/mlusBk/ftQImoW0vVZNRQwytpo/ngGbPPLWDwD72
m0rUg+aTZmfVsXk1ymXCw54/N4JExJXjp7XoavxqMILPpMmFC4tz4D60VL9RSnrk
WHsoQ7QCm3nfXiUAUtws3nGJf6VlrbB7y2ewAvYXcKmT65gWxuWkkazIhEBKRZbM
/o4zL+/4jrFbZV0/Qedt8c19WPtmkzawILPzW/8l8Hc1uI8eWVPRPjwIwN5sgM1y
c6rRZwG9xZ77tiQnSfrnG6BtK/ngasR/5OBEcfP2qFRiNq06R+WSA6jMDhXEGGTm
tQLseyhGhtQwX6wRzpPrrPY3LD9TFkxEt0VwOD3e/tqjj/E9naWtxqoUBuXzhOia
cx/FvnwRf/fGx5aPRypHDqlaNjxjQaD0UBQogbhIF2PWNSkSAgineSV76Diu2jnq
HeZTQr/yZtqbm6e1x7EjCBS5SrG39OYQuhbPYMFuOeLEIVVnq33TJ5ARwhj8bE5l
NIEX9lziBjn6i+7HUFPLjRJXBiJ+BctfUlSITn4yk2uQpE8IJzuJ46yFJdEoSALS
3la6toCYOmZgrrc4oAQNvS71SawBA+HawvhMtc+y1q4gCCe/Z+T0eTIolh0KYCK3
CwmBs2t35SPRJpsFVsXfoQBBAOJ1akgLOUVNKS0QuAutxEmfxua+qqncEisAYbQO
X8YTctgBIlrle1DDFFI+h81U4TEeF1nH1w49z1o5jkSyL+BOcP2uu8c4GJ4BQG7y
xNytfttdC1p30caVZoARgBV2Vbe/xO1wXsA+B1K2+8g1+8n3aHHyh9Vw713x+nOy
3HriJ2cU45dpW04p861ipllwC36BmLmdJd6NHNOSHtLv86zRbGM5/EtLwIIihJ/G
PFRhnQ33QngfSoDqKlOfxLJPJ4YwjhdDGYmPags0d6DFqNgWcpTD0jXSg1cx8kPP
pv6MRjZbNLWkuKS7K8DBb8CT+FivLPUlenIOLS4dpwDj6BG3MRseZ4ivUpjN8WB4
5RALvavYD3tVFS96bROeyFMYTOgflU6uhw2iQOQujmFIpxvASmbxzB9a/ifrocbD
YFx7sHRYjAmKMmoxCDB/kw/x0SMsqh5Msgbgu5xyz3pps+/z1flgDAssrC9PCU8y
ghTLJUCmhDuRyXWDLLEgey7RfRZEQ3jNW2HfwmEnCHTL+fmjs0+p3R9c5MBFBJsv
VCvwagdkW+YaFWwY/+JhvWx0YiFrCdYWo1xmfiHHQTm33H7pLBSpvEeIkLlLNxYu
eywqNWpt6SSwjbMHOXH/f3qq6Qq8fUfORyM7+DEmDNTeMTsEhwyDIpq8w2jLBfD1
OrXdlMvscxbriGJZKr34fXDFxDJOarLxXFuZpeLy3xg509/KO0E917Vi3FcIe5Lz
52sGZUqlz2Icvv/+/QZ6aHU8U5qeXWPX1lJnvqvvzaLAyKa5t8LOWywAIe1Kw1OC
GfqadxJGnbZ7TGYPGyJPC0OcfGT/wCrmOuraU0rSlnzBVSkpy/qmj8hA4fz29FNW
bCxN1OeRwAyI4gWoDhIS1lOxf9LYyuqxfmNYJL7+L1zVU5/xh2Cs5ckDhurAvBRf
AUuLilTZih9NX6aBXV8phmiV5S4ezYgW3w0pYXvd+B5NeeCPI60/zJq+/dJg+oF6
OmLflsR4knrN4kJu0Ea2OSBiEFf5on9ShZTuvD0136xz/aO+TWPq/rWs+nXGSyXN
btMhtTmtSqrW7iVVQbWPX6FmGzzhgRqGgDYkrlckL7NIqcvuhE4amikXJukiCgUX
40xgVsmjLkm4VoKNcvsPft98IxSys0TdIImsjoKjoYNi2uka7enePCs1TVKTmj3W
qsQQTBzItn+82sWK3MQOLmzHa+qVFmze4mhck6i/pcgmwGk8tmwv2BHSHFqYCwug
mfYkZhIFGWGGDVhbhxhlDNG4zWaQVxfoxt33EYli8n+Tep29yCPa4cLjOr3cGrw5
a4JLK9Ts5ECuaQhwO3lXzLDlMQJKJMWBgirjz7KBMyL8wlhqXzgNwwhRi4eAHI/a
Dx/qXQXTy0/ymu50a7WUR48YqBW5G37enEN/TZApDgyEQkCetATTOusbk4aMQSV2
iV9kd5vi8lVmIzmNz/Yyu7pqmFdDv8JbbT+srZ0Y3SVORmuD6o5BAXuNy/rVaBlP
Z5+haW67loVIsv4Tb5lTvMbv9jBs1WjPczbS1DwhnpSW0BbRc9E12Qxu44o0e0op
FSDOWYQs9Ip4M6SZrI9zpKE/Sf7I+rNC+3/oMT6SAzfOlrNXYHBZxvS3r1UTUmtB
6HibulzEWOJttiL30tKPc/sDxPO+AOmPoV8GOFgOz5WWUN95XCldvEvRl2B6a7vK
2eX8OwufjIjCvvPEtoUmwzdVNTRmN7s4bOiPlc31oqcld/ABXoYgk7KMfUPUR0FQ
h6uS9yJl+REqbvoSLudwhzMDP+Cj7J5NpzieSz1x6/A2Mi1ale5BDkFjjdzFD9dJ
qzOsC1xeTenueEX3COZby67foC282vjkpfnMq10ecC0tZumcCY/Vyp2pRFZ/TH2X
WMjLJz2b5bQQyAbZb1p2cJU2zMvLX4DWNBhG/WxdhY1sknNbe1SzNYkOU+ORXHoV
t5RIRDF6qSgtw3wIN7qyntUcjZldpeNHQazYNFAbI8IVV2QPMm3jqm7IUEoh+Oj2
NBZBXmhyNWy0AIASbePJ6sqVywiZge6GNMvnYdxRe9vDMTJXznn+2EM5Qn3yJG3T
qlPdn4fYYlK0f+w/tOILOuGk28a/Wt0oz7lP7g4HIa/gsBl9xLhaph4E1zRm/q6M
IKtyMj3hKiVMeVjoLBcO9vzT0Y35k8rT661fyfUBq/sZ4fQhSjQRMC2G1hwTw8+V
ZPc+xc50T3iV952caihcmRnxg7SN9KBNSUcayGPhFcyip/ibbLslO/SaQ68lAs00
+ZIk4oum7pi+RnVx/f7ZcNkPUuxzXWY62FJdf44pe0N3JkbviAkku31XxTR6PehK
0A54jdXFcRTrdvihYUHd3uupVPnnKgJo4HsNlqjvrsHHFYN2v/RBG2bM99Hn9Wk+
oh9w43a4QgHDMF8iUCjDnUWYpVlEF78R7Tzmdd/QwzJzWFjoUlDIbny2sG3B2vNA
jIGZXXHa3qHNGxqiFPkbhyXtwwt/sJL04J69qL0RjGQd/21egSKDNMPO9lSNMWWz
fRp+1GAAk28hPhHNfZKMqmtA4e99zDVqM0xt3uWDPS8NCwGvaAHcbjGfYazetMqc
PpcMdYloFPmNIgd/qfFJX/hcZNPZPWpvpamqCZn4AFg71jenbJyFg6G0/XlYW+7d
a0jZLb8b8lpJa44WtLx4Louf+suJpXr96KE/FhIfFGc0XHx8PzDYsPbbyYg7UucG
Ue5HPdKUzXnPB0aYkywefng45dGgg0HR3ZxR+zRMhYBLnobM+PVMQVBQ8ttsFw91
cpuDTbmzsgaoC+p4R+U1rDkwipyiHI1fjFdFzqKvCsJXXTVxKKalFyVCnc1xER0P
SbjqEN+VWWwqKIMpmVhu3E+3w9Gz+eUjhxZGgz6PplUXRS44pPRZNflRLdbBIouX
0WAQRcHTioxA1BvMLWdgb5WVR29KZtRVFnyidYdzCokqM+R5i9QIX41drSX2jn4K
u2D/h72B0rCfTApjJBJ6RFHb5F8BiEeYf/b/+IsDJCmkqESg/WZcUvqN5p6P3PxK
l9R/xCgR3ds+bfq+eSegFKFpbtPeZZ+9gLUU3nysbOEXrVSGs+wpH4GrAbMoRgi3
ezVwFfxl1AMtbb06dXw/TOGoakUT+TVTIhiGqeyarWY24vu2dIDHXjtVInYGBZmN
Yyf3Q12TkqQGupKqZcXbqvP96hQCDQg6Mo+5YCTvO+BvGC4Mp5bl24yJzKe4Njog
lNqx2ip/8sdJvaRBkB+WtNrf4TlsUBW/tHLhIdqoMWxSFPOgWjKH0JBgk8atE+it
nJdSRzX2OSY2SMkoLGQK+iLYRNik+NReBI7lh9dFzey7lnqxqfrLBGVTiKS129Th
cj6+f7eP2kuO7zo1xsCe/QRcjrL8Tq5GDjyHV/2O9XeOmnSrp2AwvWv2Ga5sLi+X
3qzZmLxinKuYQVXo5ra0NkRrpZY/9PH4PdAK2wk8xUbkzRCfTXNFH7lcIPv6ktpZ
5iDCUq5JIe1q8EWCe80quZJ9as+g6Vhx0bE+Ry+tI6OxOFUlXCHgU4+bE+O5UG1C
MqfkOCVqCdMNZ4FpvOJ8e3OtkCaV6AZEzVYA81QHXuGcmmTtpkDVDH9+Ao0dDQSo
p4TcYWGfNzYbR4u0BT9eRGnT5ylyziUpK/xptNg4A0pe6MWXjZDksIVlIt6HTWiN
W7iHQqgJHEbe9Be0p/pteyt3lxqCYpF/80jU/6+9LqhAGVAQh3ccE6HvVnf/MAQ6
Rxcd6fwtkzuCTbrymgl7JguGz4jyCRRMD4w5KqgCoVuJDIW2VH//yYlZg3542iSA
IjzS0OEcEoVKyRszCUMPdcSQ8JRC9MsLMkXYDl0hfNe1kChBYsQehmz1FPF7bdHj
9GR1xB+k8EQyuhNStifuWBaVrbcDpF4WjM/CHZ2GviJCoWJjU8o4d/owRCHo3NGZ
8I+678EfncnLT8/xbmkxGJDz/LTmyZfQXbbtLgW3WB/ikJlkyaIk0U7wL7kjJMoF
1nqFMGN4aoTnqntRX1DgibY9a+sVXEHevPmW3O6CQALxEG+dDDAnO7BDwLexAoCk
Z/2TTmGIrRxNFFU1yr/fbcR5IAckhXAaQ7J5CRYaxTYZhXWkjR8ZA11fFTqjHYP0
2j1ehXXT5K3WNZIfrZpTVQpcqG64TYKDh8ZdW2FlnX185ARQJLNg9JnCze3ipE8q
3TainkG48G0njFdRYiq1yASj4FlchB4AzINIHe35IpD3Jl1/gj4OYoyqmnlp242C
KCui12SohEas+XQdZJpJuAYzdcIlZTcNMTqdIEapq1TsRp3cr5wTW6/3m1pcI0zB
S2DohW/oIglBMK6zFC8MloRgmXEXLbnbcrhlz9LiE7tvtVnlBM16HNn4tsGXu01M
Wjwj1I/CzQGc6OL0d64b2V7mZmv/XN+x1M2aa9jrWpzsOegMN0qNJOqg+k6YTQoP
mkJcWveYV7TxymkpxEMs//d8uQZpRyjPld7v3u3FrDaJCuld4Hjt2W2W8d/dApDe
wHm+8LicLkb9LbcUei9luKt4YFPS50sVn8eojL5E8dJ3mOeGQqJIG6sFZla8g61P
T/Geeb3C3w0QmsnJALaweXOlblrpoNxIL5zjlKwM8xk16W0neyk9t73NRgF43M4/
+xrmUvtVuNcyszjFgPwuHqQZqxkJ+dKBszRnbFDESPp6crkcBxBcfZZme8LL0Y9Q
Ck1UIkC64Yyl+kRWvITCHlR82pcYPcXFgGNEHonrNpC/DV5isKY4is4834pIxXYx
2b1PopSMgfC5L4CNPZKsraFHM8iGSY5xNxRpZo6Haobpr2Bit5DsvWhYO8pjuGR/
EMu/8+x64SLwA9x86fflhWhPtvnBe5wRVpLFpOA0CnV0pRanlEuu+W1r0Vw6MO5Z
+jeZmuzPNEGwfhEnbvPDqQkJXKk4firc9z9fNNPfyAdSmiCljKkP+OLdUjpJCjax
lJPPcSkra7aZ3RspfdIM6vYedTUHnO6N28GvEZt8C5rNYYGmdcKHTCfnY+9n0iTu
y0iuq5+9uOq35QGn55duihIfEUsIAl6Nk6ynyrUZW9tbtl168PqSj3a3y6DXRgl8
8PTEvGwH2UbNyvqu6if9v6xERWr7r/A8tbbePkLmROIL2kS3p6lzfPG2aKLZPGeT
J8VVFaK1dC3R3dcc8S4YAgEyjbkMPa/VBBcS8dWg3Hpuz0IUZ/NRxI6zH4WQn2Q7
UPQXYS+7fpS2xReodytBtd1l5oJewmmeviQuwmNEQaYjxGP4I7P97gkAi6X7WO57
cXJfhVsKIcJ4yKooueVWbKnCLEG5cuqCZV9KzS736CkPHGcowqVTC5WapY8s2Pf5
goYlwj1xw9VevS1vLS2TARjtpgeJZDm1rVIF5EQysYVfwtZyRjvezygsDiUERfa4
ygITraJ9R6d28D9nQSP455YNpfTxiBOas5jES147tdsWZdiRZWyX7RJRegKWvOjK
NqnBRjVuVTSc1n0teNIuxGUNU5vxVceKUBI9OGTqDUG9ZlLn7+gp9AN39oBgaPrd
PuzKKoSBFDiNQwf8R0c/lS6GlRI1lAiq4opm5qoMn6GTJsavkEk4dmYvp4EUTaCZ
WBaJN5n+EWFjzae8frSzgnRRnplG1SyZ7svlmXREsr9cj8wSPXTu1xK/dbk5IxWo
MNbwC4H/Qud5HGKM1NzvzT3ZO5UFDTeoJfxVjPTIGKMwrM7Pn1BZYEtwzdpOkBIs
JlyPxsTFBZFc8VM/WQvlvZDXTurCjygYTR/UmrvpO4G8gE7lZMuTIs0NyPJJka79
GeG2MLkTfdBXbycXLuQ6Tvw4vvoVNPoZCn+q8PFu3cRC3cSkDJYSTg5pOmqcD2LD
t0F1r/5NzlUsntDdcyNR/k7JygML+YJ797uJtEUCMHVg/cSsRGEjt/PaubI9NxO9
WjjVd/8KLJdXUbJs86UZrtDlNrQEsjyNyAX9JrNul9j31c/aO32j+ZdjnN1Cw0Hg
M1qDhrCDxyNIHQeNBcCoL5QH61/Trko79yAmVZp54RedY7BiSQlYOiqL9kprLWev
LXGn08tvS1Mzt1KkoRXiYSdL4gVYfTdrC1UCSoVHGPG279iJKbMsFyWyWELTRvdn
oKqBKyog01walnAlE+wcCGMZXhbENvfd5aOcqHR0TbXA8lrIcctGTctRT9wwkw8I
3CgizSTGeNu9i8hnNXFYKi5CFWfBqO5EY5yIkAlPFvEo2LIBut/jnqkFY7yK+yJj
h7e5Is9QVzU6kqFYNWN0WaMT9mRX+WBvKCcXNcwrNEfgPHUzjr91seQu06U3PQsP
KlYiFhBynIi4Ul9+hrUCZK+oZYTc7ZeJ0xEMZEUShI6VQd9//wjV4rRvZdbVJPpR
RJA4YPYlRC9OGOYTj3Jd5JCy/2QIMTXlYkLSMmN9juE8+KJIKTzwljW8aLQjfBR+
AZGN0181wvA/NiuS1L9E2l3KH1PPe+MwiN3NewmYsAcOgfvw/DGOgCJeNBBxWX2x
QFZ7ttak6HGRt12zxE+Z4xNR4F1uFG/CIfQTZLqNtmLon/4waxIdiKNoXiHFKKeb
IKKXh4hYFQB9P3EQMPVfq58yDDbGsW0NVaUfNILjvP7LtY7sNx/v7jk7fRRYKWfV
QRMpXJuGK8Gw2N6umnIIpXCZdtU6KebQ3Lxh0rwHfJwhV3QiPAt0nbNzaIVmfq43
3B7m0zwhAzHNgMRXZjoaKF+6zbaUsONEW1wyDJyH2dgIMx8xPgoxAlZRYI+r6Fqj
p0ZNvmWCFDOsYp2V1cos+uzkPR+9rb4AazPd+G56ABr7U+4ynl0xb99KU/kwkA34
iJi9naBG2qauG4Pmhc1S8+9Ig+lJcoJxeGb3ce5CZo0sIZ6rJF1fyzZC13oWsNQ0
YDcQcASpf1ixgSwyn/FLfMVR5dkftU0e3wJVlFC1hY75Emrw9W/zbT8WkN//TJgH
Fki4i1EpBB5wBPj4BKw16Q82Z4LtAHXLBmS99/bdD6zqiROExKrjLt/OyqI/R3W7
sx4v3vQLFpUi2hUvz8vjU4AWpRYVtelrRr3en1+izzQbJ+WWexUl6SkDjXQ3PWIT
9hPGsXq0F2L5CUNgQhB41bH3nkEAIRVxwclpWy7t4cKVuMIQergYjm80AaYhh3rM
QkoAxZzbwI8wa5ZWggGf+zPTLxfrQ3q94zAPwGSxqghOwlyJ/dBE8ROBjbF8j68Z
qGCrlOpgJWIAFe/t0zU1e/MkyvtAIgZCKfxgBecN0rL0uBNEriBayrXSXPloCnPs
prhZK92nGmwRgzzXDsmbCz0LoCCfCedAWwfp940ahNEY3fbpHfYqqNBx/OUDUhfU
6Toog24gr7So4kOwMZh5mq5qoBnijeG9BTKdD0UkZtv6bAg7A9EeLpPeY/Y4LUBz
DC0UjZz9wFJRt14Oi5k3befkaXZOgWSM4CDTdjtLoXATQudUjJ4MCdiDz/wtJQom
yFnKQ63Db+smGQsHtNAmyfScV0xQZaJrr5Q+39NsN1weIiGqQ5QehAqB4YkZoIC+
YPzby8zntt6rWhjgLy3xAHJw5dW7qQmA8t3cJhylN+H26MOsl3kD2Had84DZvYOC
EXi5rRZN5B17n71JRgtaaHdbTPCf2US26Sju/6gRkZk5jgVO9CmFgc9LvYlMwrxC
gM0/CymS4HcT5JLPJw/9cld4LpI6YOcz5PBuGNbEH5R/bXjvc2Utbm1iF5rCBpJF
PjK+4URS/52mW1j6eRd3liomosB1j8/5A1aC7OTM1pNv6owHjCtI4pVkMbylaTNF
yqc/pSDytncZkbRyKIADIMWoKJvuAvgpRsd1jUJVMXcQ7QgtzIk3mNeGHiCuJrpt
GYIt/3V9BF7YmFhgYQE4F09eLFlasbUGGycJ+YMBlzgML8wNBirF3q1mBh9LhOi7
ZKR3kvTt4d8DSOumS9K0psNx8MIVCMlP0Zs6ci/AHppQhBFAeqXMiRTvaQnOf8HY
I0fvbaeOOaXrimAkIjtqUwIQwh97O3kJcBSDk9NsQnWtq+wxxuN7WcGIniinsQFh
lt+LuZY7zs+PYWLq6cDbPikAfKm3mk0CIPSo9gOdURBpSwXe367Et5kziD1sUA7W
jZjwRSWiWEK/qQvYZXqYFY+haL3rJoW9EodWh3lWLZavroHoO2R6oKTgZNzxbYv2
lUuvckG0XYJDZ2RqHjR2mxZelwIMPwBnNV6z6AwIT07AemDisrqxkIVbbdOupOjj
PrezJMxO8w06f4NyteI1iYV/shUBPUXXlg3oVoKGvFmGToj0ddjWsaDfpltNGK5K
50VQbvPIzQ95YlWFWEwFhTmKhK9vL5+FvlA6L9MKL/GZ6qxG2AGJOzHYuUMkqjd5
5Rxdr+6bx99XZ8dCv4Pv4pKYDW1PJGiMai8/65LM4YjUeAlNP92v1lBvxg5cVwCP
Ov8u/0vkgbpJi0x+ZTbbO8fnkscvkrho/k9kvZYWMURc2gKWOzHy3m2OGbR/IiZC
k/HjE4h7NpGUISXWJckF0YelHiMSYaw9+YzL5n9KH0aJ4WqHLUXgWki8DN4qbzIr
TV+f4hX8qm6ejShaSQdUJ1JnYgVPb7PQvnd42kRk60MuEiVj/idKM4bmAeHS97Po
t4kpJeW2wbWR4UM0+GvNqNSIkPVFiC5CDa+vLIiX/UMpLdUvaFnF7G9ft5u+spJf
AeN9cNGr5Uuc9Pn4TogvbUDi8qXRfpRxc2g7ib3UzWWY4agY/wjfx+XyZooyOc5+
FWWitoFH/21CU5iNjADjwZi65e0A9KvgEjee4d2qlzGPwka6HJYk45TzPpcexPOi
Bp748N+NmH1FQ9cY8rmAHigTH15YXRTojj17gzh9/6pBAOR3rbV/l6i91pExfMvv
b07eWzADvbRp7Q6yASbz1WkRwZ0sJRdW1BDd9QI8wMDCwGgrYhq2IfFB8OzSnxTi
Yl/43WMHVSP9IqUyw5V0iBC1Q8pb4dFoBSfoKAApkJfoQYGB03OpeZ3I8x5kt1x+
iykyv6dOxYPQrdyEFvUHaIc1o9nagmD0W2iIa8OXMCF7kPbOSIDOR07JFseqIBpY
uyh9dJQLilK1CjFO0yjsUp32M90OEQ9lPmU8s8QwL6wxcmtd8tEWWapN+2ZJwxG4
o+SzjqO9JiMILkAtYhv1gBAJ8TgHVIue4CZlXsbCivBhb4w7/oqWUmUD6yjTFT0j
8TcgcFNTRdVU5aKGcW0AfHpQgn98r4T9US8/ysqA+TQ4LX3K72XC6rVKGpSeyrpB
Y2FVZF5YrFOKasw4c/Hx6HPjbHWE05vP2lhSNL7y237WfOMWgUqt21B4FZl+a1d9
OuPoiiX/dGop6/jBfN7C97JfsUbg91g7w6kGQsod0j8LgQYfZQn6Ib5r3O01fSWz
Qr40CfKi5G42Kk1FdrVKz6jccHFJAV8lX7uduZh8j5yLxe+mQ60MD6ux2X4PXWBb
jqCRTMUtTEqMFW9WCmcIK3V67LoI7HP7E7jf2Dw+g+0QI4iWNdbiboeiCLJjjhZT
xGjU1+Q99fCsMqrV0bsxLwn+0ZZfyKUcCLyKpUyePJT7ZYZ2+m5ifoBzg5f5Tkej
9feZJAJUEcbJFVCt4DssZJmLi2tshoktOw6qqO26FvnUJC0BiCcN1aRaCLR/YUaI
G0GEBb5znn6GB0yclBsenmo/Lkr5yy04zlkz38bRhbs3k0sogVfdOphjvEeFdy5m
Pa0eDahhrelVFO9RBo5HbV60OCnyxkD/Yg7f/k34KHiDlcKp9I/DArJLIAASTWhs
pPqrfsmlLjK3IfiFw4INrKnOzsHA+0rkP4bSS9CRtRGadPP+jCE2dNh+/9UsyAuO
oiXRr5kgCl4O3OvDO29U1u+x0IxgO7E6k8I/fP4AtA+jEAFnerJjnjJalymffTbX
vucwdohdFZygmDAp/lDspXlwmfJldyp0jBBw9F+9UCwIwTNovCsG0ynh3QnLUjDs
CsobkNq+guIpIm8iyNLucj5oIuVxuSL2+9t7Ie5vBUI5z6MluuHtmpWXkDLz3FB6
jvWMr3HrRpewnqyLOOg8tu8IZP3NGb4fDwQ3ktfKu1aqUFkhRFWMjkI/yPEldtBm
UFFRLTYaIMuHwOceSky92V25TFvA5hM67op2u0c8dDKQIdHtIgI0xvmwOBpJE/xL
CsGO24Ly8T1xTHUxMtgk19DLRNNTxhM1YM0XuWVv07Tj3l86ohtyoS3uKIwhCiCF
t4Gsh1/ceV2rZ0lvzhxbhIy969jvyPBimxoQhIOKYpvMaavUF9wPpQZuXVhfF+Aw
AQbG1yv26XoU0A0RXzZzZm4IYauDg180Q0dScn0BwwLCFM5zjuytx7OWzEg9Io0n
QkKHbjlqgRnMOWLalXxn7uImm2X+IPpE2BVBM0BWRizWW5ybDg60nzNe6Xhsicnk
YTTVwe/1c1CXoeiC8wSk5IPIpeTixoRtbYa5cOiykOA3zj8+ZYUjjqYMQB5xq79Q
LdYwfmyRU4AVydpfDIiHPTkOi88JCyu7INow7a3D06dEnzpQgoUMR/9raZK7qKun
fjgyxOWo64WvoBk3WMdjj3TpzOKeBP6Ou5YRg5DN8tM=
`pragma protect end_protected
