// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:31 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IV04U7C2+cGNpqPpZevlES7EmtF1XVYVqtGj15pXd0Rvujo8EWKUADy2z45KrKY3
MTdVqsF1dbVBa0u3fJlnXkhJ44EelJfJcqBEs3ZTG0HEzW/uM7m4b2V8xSBPEa2d
kGV47mklbQIjlslMux6EDRTsEYgqUezW8PKSMYiNfBI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7104)
vdAy2os+gGv1meteD8NGo5rvJ7oMPma4Iip+ywINfCv9lN/ZrLOrqyXo/Kat+ScF
jM5Z9Ty99KhW5JpHL9M8rcvAOhKuLus4wEP0S5bncppsRMtELL4cajPd7JEvWHfX
z+8YR9yjKkavkJBGIpqfft9KiHfInSLxAYTeK7iwtGIYCw1ER5zR388DC/uWMmS5
ct5N9ajw9ocs3Dx6bngvxK3pdMWcdKSUyT35BoY2izboG7t5F0/YSYtRvyaSevJG
YM6yTHDv1rjMuNax6w4lk+XJYUwJAb0VIkvMFm0bj1JbTj86kC0H2NzDyj7lNno9
hwhMLzFX8uVCnfFulj0HAL4efHSycVAszabD5FMV9nVNi8UpAvitvWOJPd8mQ1G9
2kOve2gSM2TvPLs4qlHTRwgvbhav3gPB66NbEMGxRahuKjeRygFbGz+pku2+agKl
kYG1502TOan38o9eEBxWInEPvC+b3qWYiIs9yOzOOC6Z69dwsqZ+T+xZlDcFZMl+
I9aVKFz8xUPXjAHTINHLhXw12flTr27YIjbiAaJSe1e0n0dE4lmOkl975/vJ2qXl
AtLdb5z4j42tm8PaCuZxRex7UW70CZ0w86cAsEis/5UTe/+oxT9AuxMaDQocd/FN
JQyP0oRn4IrktkupF9h+K8Z+3crA/9WJaAL9E/109CaKPguIF/GTgCha+0C82+/W
DT/J88phzMYCXQWBqQu8TwLEPxS1hEK11/ABYuFb+RR2UiB4f9VCKo3DQLOjlMFG
jGVlURu+S+sGm/B9/s3ubb+IRRMrT2tyZ30YFLOwXIEQIQ6Wn9E2SIjzoMdImYy4
B7yO3cZApLJypRTG1QSo5mEQf7lLS871ijKkbJD5TE/Q0JJ8orZgruvX4trprXWg
14jrPrpWaa2BSJn1xzw5VCh6gFxDr2v4TcpjyZjGPSS6qsG7upWHIAbee1HQOo7w
UE5i9F3xxMLy9eCGEfM//H5yObRyyNssJQF2r3PvZpl66sZyNFHjgmW5ohtkosAL
nH2E7EJJZ+20ttGBTkvCFvfEobTTOz+oYP99i5cV2SNvv5SA5QIWrE0V/4jNyAKH
3KV8HYPD7B1tAx93Hncy7ROXWUGKM2Do7GoRlEcJK5okk9/7a23AuQGPEEVSkM44
SlgBwA1vmVTcrNY3GysSawMSeKJoLVeq7GwyAus90QenGahY6Eupc1mXei5JgSxP
i51u9Q5+afNhBc4nA+v4hZAZOv8uXVjXI0wuG8M1AF2z7520Eh18xr9dYF9fOvKQ
MoEOtKOzyV4m/wFkp/Q0UkdA/F8tDXBo8Z0w5n+3R26EMDxCA4e4kfkVk+0LlQJv
3oyQrc+vDvhVV3Cz8j6zlTGTlDVbiTGWnNVVmMTdgLyPlApcDa0qt3dPXkJQLb5g
H89c2D+XBt16a1W5LER/SRlfmll/mBa9GdbQkihdjQxB+vrG6p7weLzlu0r+rjYk
RvRJaoxvW5Ydkb3OkTdxJvjNY71QKMPvBZorHR5aB0ExFY2NRuSXxAM/Gt7G/iGa
9V5ikVTu+suw5RqlIOUwJS2mNhevYaHPiWreNWcqAnoOYOvmSlikprguLAiSGaf9
wygjPGgppF61qWUzBz75MSMPzNbipg9rr2IMD+t+7Lm3m8HwSMMHVCKdL6O5OwiX
GUI6HYRt/O553qcg0BY7UvCx2Hrasdvet6ixEv22lbp0QJoH5271nvm1OUHHj+U/
DSM7SJUdSsgERDGIH9Nnxqv3QlawYuh3hoxjuOqxg2lzkIZBEAUU029CSi/GOG4T
wEaAZn7s2ba5as5z8I20igVCuuIu7UdIc4PlVn7L3cvuxY1hhTJAsI+EzCxmZ/0D
v8svhTBGUZgYmNTZfI3PYLwXeo0BQXDQhoFcBKFij3kri48WT8E3CzIUG8CmIQCs
jTfuyjnsnfS+83TSGUYPcVz+Tr4gAjI9+XS8Q35qDuvLcaiAcZxYiB1c+MPYF5tl
Xq7XKyj8WeF2zs3tUoREeJDSl5yp4Fqtv3ROmoNMNntFNgkJWiIp9hWDSBq/4LW3
a9Ec7OVDiVawwXIxQBNze84rCUTLEGr/nYo5xP5p6vK4GPWBEzl0diCCi5iDuX6x
gq704I27PdxC4mk622RJbcNXS97n3WbJEL3KpE6zrTepqXprFco7WP2GqHaaF/pa
tyXoltCTC3Qo/CKkGlI6ACuTDdZdZh8R8GZvC1/l0ShOkzXQi4FUxn7/NQruvt7E
0NZD3yDtRMjEtt8QJjOnom5hjbeOBan12tD4AnmsFv8aDgDm6PWWNI0gl4zCWmVb
mXyrb8Rn9H5v/xY4JZuulFChxhydNel0QFH6ocICcdEmTfzexwzqdzolecXNRYub
fLG0waQOr2dDMuj9tTs169PGIgz/2rxfeYri1PZAG0druhAULETSY759CCJOXGYj
LMS5gQJoP1NAL8nleGF4Ous34ydtUrtDDf/f8ZJk9ZuUG6D4snEJXMzA3ZuWWv3N
dVrShV7MJ6kGvAk3L8FrIQoCK98ykm16iikBM/BCnaCX7srauTYOV40IbElkEajR
8/6OOyc5nnM/L0RErAX2ZTfnwnzLuVqwk5f6+JhpXOKJGRjJ2Ptruj/lpDwL+W57
VKM7JxUtjk5Q4YbCcvKyonnyOz9StB+N1U/WbemJfKi+OeULqR/yqdCD4HsGN2qp
yeqYB6iXvdTM+/GI1B5mKtY6/jExFAYONhowEV3mlVsXLJyMpAeWl9gDBh0Db10N
iMZGoH9BFLKzFxFBQtU4090cUDBdz+nx/MWrFXZ+YhGku6XF4vbwf9kCqVRb0ht4
ihVlGCGr8NsxG8o+yCkpPYpoYehWRT58qVOD91afIHUpxaFbqh99O40sjLf9y7sx
c9EtVjxPSPO1XWrZse+o9ZxSEY0yLZmo0tZ8o+sij22+CHHp9ajyT5ENV8/iJxfO
3TT5uX6fxE1qFEFJxM9XGIJjFoX9jVy8dOkzye/kVYs+XXKpOgLEuOvLKCEpThiK
CM62L5k+RXNsP5uuGAnPrpW+tWnYPclo5uWOpucaWyhWl3KAlK1d6HS+EiSGxokn
Cu5p1ennEf6MC6ZZLwpcgbBsAxom/RhtPBJrC8ie2mcBsY4wzKL/asEUhe0ne/Ke
LFUcVKVPB8DOXPJFuZHPQRJDHeawWZ1wxeeiIUql4Fghmyt/1lzAVLcRbNWEe4NT
6oFCCSNor0qsNDiXbIxHcNgvYBTFlGTmhG4s1upkamF20cdMak6V+wXsC4Nw2KC5
JhUOvIYXTXuQpm7B+zAo0O3Qg+m5iQamDv74Sz3Z4JFxHKXzM5BnkhcOKbIeytVt
dD6xIcAlfjKTtzbk1AoP9Z39+Kz95MsSIkteAdXlt5/LdjUD7jQB6IGl0eXBcaDU
EfQAJWjHG4vnwq6a6DES/ZborpZv+/RFtHzMA7a8BkRShSSXKnZq2A/DygX23SM0
TvFmBiiq7BFMj78ANuGuV03ej9E+Vwvkhp/uBT06IcC8797/2T3LFHI4fbfiu1WR
OLSq6NAC9LrM7VXLET0F9Xy704eyPnOpoCdXyaIoDdQ+PgY6QdxlzeGtW4gj1Y5R
zcbgI+KBdS67pxYubyA1U0wh23PlbIqbybXtj0Qh5FY7mI2XspYzf3kto/h4uG6A
ilrX1jWoqH6iFKLYEygP4KXEG7B5n65a752z51tRUQOexO+UaOgkiLwsmcBU0Ij5
Y+3GH1Lb4CIqQ1jg2WpybY+k9Oto2m3jGUUeqWO/hMxWtAF4v27mnZ+3wYe3Vnwh
cfa+3QCg+SLnU8XF/I9bbdODNlHA7opgN9SmPVb20eOZRVGIdKV1c6BsnDmy4ImI
eymAzvjyNk7M7T2b80fUgcO41537K/u+PK37IApe1QV9qYEq9PfHGVchvlUkQEov
K6g5sjblqLwdN8/LEEctD1y1O9Vh1HWJNPLOoArE17B7AJXd5CNwsxXpLim8nlYi
qfrBSGkvxTthkZOY22klyo0bQgPkoLaju7a/+Z5pZwlyWSYZRGd/zMjIgp5llEYn
2SJuX39mQ094o+evMoH9LtxY2qwbapmv4aDmKESAdyuyVuI5xaQCIqdYtYrLACDy
wgkb5lPW18KSA6E7zuFg9HcIb+IZI2aCD9iP/3JtvjTewoLYN3NugecQ2zCkFt6K
P6GypWzuZGQjvhJCM8nmNNkv20RnG7GsEVhu/w+IaYk3ky5JxrEtZloivz9tZyIL
CRlf8IAxt1i0q49B257YvF67XLLKLjdKaBOKAmrhpfIvEnFOAQTcYamVelIWNR+w
D0KNICY8ouJIdQfoUtOA0KlnkWVoTQwqDVv/bLolm1t8RZJmR3H2xTv7JVbPcTwP
VYmmAfyDv6f6OSGt50Gsi6zhMugbc1vsRiDWB+Tgu3bveTjUZYAMbdhglW3kn5A7
AYaaWMJwbAgn7aH/i7igdNESiW0p/1HvEX5Hz/CwYCdx8LBbTvWsi1zpyPlUCBDj
xxuOlHafCojzQiEkLZLNCUlg7MLGA8BaPeTRJVyTyltlTlXUAxgbX6yS0P8oxkXx
EzYCn4PPJizUX5f/8LDE9jW/H/kHjHWfDfn2P65aGGeFoJrMXNj9kJRu/ILVQAff
IOLldaER+qruxnu9u6393eAUS0CbhA19oZQyhb7uKwqchRg/ad48RBFIwK8T9Dg2
NuJLcny8AhanQLyQLTDdONVkO2ZrC5zm10qbdYP968vcTyX6Nf5UKV0BUrNwv7Au
RWAb9fHYDiBMpLKBsO36WBs9obKX1BFOUn/ToMdabLlvCYAPJU6tmyOuRI0YK0Db
jLoMsdxKlAvuNMYpYXTD6Micn8qt5cbdKmWrOyjYNw/bGUzi7fMFVYpFcMXS5oD1
F44XPh43Bt1sxicnVfydlcI2nJe/dw7QjnvOmcuYa5yHNHI29gphM7p6BuucZSjr
S0FnHgkjdi/kdIZUvKq9Uw8MMcu/4f87ELdrcXbYcz7csUMEZMS6GLpJwT6TUPzq
hKTqwvwrpbBeL5tPDUrmLiSd8RqNka3qLWkNv7l4hHtVvIuKDEHGgyeRT11EmU6w
UMLwjIDI4ptRu3W1tZk5K59XjRHySX27OQlI7yioP/VaMlxc98reB1yM8ERjgNCR
UFZ9YnO/AiLOPGrTJKP/2llA667f4CUorpAXSycvoAM+9ye6LceaCyGEdwUI0qka
Ioj76bdE410zLWVpx5nCtKtykhZYHPVAjsDV0K2FtWl9LGMHOdKDvFR6U+3q7LRF
wKQ6rCOhcD+qnQcOCdQfNcz8/JGlOuL1twK14obrwHJvDSkIcyiSHr+v5XOAbWgm
cDx3OqFjclLQSSqbo52aHyun4Yl5UT4wyC2FM+eSk0wuRtRyBf5wfTNuCxoPwky6
tFQnnwnJpTypGgwfwX1+2ngmOYh63GYAf1IR+WnBKnlM7XfuCxy8OKxSuwPGNLRQ
LafKWo9AozPVowxOvkGUE7zpTd/21bc81y1ieVFC5zHC5GlPeLw9m8SbGh3pac0r
875xtwG1oRZBU/BsME+57O8hofBOseUqvIohuh4D/RhgHmXC9qFNSF1RbswiPI+F
O749oAJ36OwJ8DuUqEASEH6c4IBNlHjItAez03ND+55O6+GOTGpRV4w1McHkKAOQ
ZK7VPcXH9uRo65NaKIF7fcyPOcp5osTcJfvrGU5XMr9i2R/uXz5i5ZIw+Rz75yK4
K9ZMQm/vYWimrxZeQ3+XiOTFqf6eOjA3Q4Ply1kgppbax8NZZIGisNtJ6DmCyX31
OkdwT2Rk59uZaZXMF5+pkrmveXrxJ6XFdGkUCUHamEKGbP6LM8NaxmSex9gV/RiJ
1aNr8KrsmXuho77drvQyY/xgLZkifV/R/4ppr8z18FNhjZIDPE7QAepT88QWNSN9
lWdRApGE6hZD/46dQPPJIAlkYEyO25QaoYhL/CPY4JlLlXN7qyPH9HwEazPAqOCb
enMVpwfHbQgHdZDcdZI38dhekBDUWecQAvcV5iUfxpkwMd29xw12LAThGIYQg0S4
KE5I32R2Q0uwNGBjij1mn89oeklNIy7VCxnMANogoHqEp+N8BXwti4QaXmHj/Ti7
Q8c/S1hMs2hxxUGTJnyHYLajRuJp/aDKSl6kLyzOIfKAGgvJHpqAGW9cIK6e6ZF5
adssei8cWhqlBZKM1pmJ3ZtX0NvK7qYD2vZGRbNypNfJ1/GDZbqbLAk1YLMyHQwS
4L6r6kjXdiSa6cpmkTdjIWFDSne6B+zw+DSgOWO8Ch7huqWF8RydGYYhxN+ezmkt
UDo9VLDZcubC3bdwwlQbEWHhuKzHoKb215rIFgMpyyZL+mcqOZb7YBBHnN4qCxoy
pjJjoJHa5FtkUcSRcxjp7JSwLKL+1LN6IFU0FKKXmiZs1z4b26gPkj+QJ9N3BzDU
STfqsMhWyjn0lE1ZjG2ben2JPw+O0EH64qwkicKI5S+4lk3/3ZY2S8WAOaRxkdFp
oJUvfG1I4jhM27MzGee+VzMMBPGWGWyV2DJFFitnfv8o6XTI/RxnNNBJyMz1SYYs
pOMM+D8RgsvI0sQ5zIUq74aFffJ5Iv/u//sSeRAnjryM9A9DCGimfjd6olD4hjE9
iYxqg+YFa1oUSBaWmWXTmxc4pjHmJ3OWY6V0maEJD65YFFfZbAd9h+okYZRNFmKS
bkn4Yu+k6MTwQK5Qq6Hef2PtqU42yGqtAkvceN2vQ1wFS9orh4BJYqHYDDrz3fkL
+ZMzP/uT8747I1i73hf6EmYwhd0tpoc5Pnw73Ah6W68kj9jPbalct8ewE0PkJpIi
2/spbb3jvxzjztGpTNTQDdEbgROK6NzYRGvrFAMR4hEPOYqIpVIzkl66XOi8Isgj
N5ylQHoNWd1D5Pu7Lpf/jWTbZ64Vajn8IIwl+KJBcKwykJ/bh1PLk/R5tATAkSXL
9MZHw2rXlRRB7zJm07APANLRNpPkkVCwYL3pz4KKT2jE9W7le6pHunDB7Spg4kRp
HBFxloloqxsibpQgQIwAHH+5uXmdlSel876r1XvxbiW4oafk4mj7ak277Rygdr5v
KFMqJSjtw3EzzR47gMkt6fRnnw1/QzIU/t4OlgQLN01/q8x2Hkmh1vo4um5NYBuP
fTUSMtgpUlUyQdbemquhD2Z26kyzqH1s7Qyq4beIWoqMd2KPLWdgonRYm5SbLqVz
mbmQC8HtSacH4IpMtqPpMYGQfqQg5NJrlxpbBI+s7PISjUmezUh0wPiQkCPOK3W4
ge9N4Ppw98ul/J8DLm2oRIiHK8Vb5l39VBVEHqjmMB0fEB0o2ugmCF+nKt8ZxEl3
+pgRqxTegl8RSVR23eThkeeGS2e2ldV6TpXCPyr69yxEw2FfW+KPBZfBa/n4REJi
wyX0+ZVSC/DebtyOBlZHxPpuX5CuYkaEsROoUJgYySCYgZtSvs8/+k5bUtKL/6IU
uJrqqZ8/tOQbzqIn7klsOApzeBldK+sJH6LXQBgBoUJZpJ+ioMUDWMPXAduXutbz
BTi8r4MfU4C15QKb78c5rVWYh/TjHv/1c3XkVScPOBZ49Vrv7mx51DSPfBNLslKy
b2v9Oy0YF55Ikc39TTiM2i5a9VoG5Y85IRECgGxl23Ue7ZWGvzodMUGs0kJepVM7
uCFWIcbgAnzm4dE7NewAAHUsqzXoy7HtGf3/OLXFEkjyZXHfny1ty7QZFExudozX
dRBMuCdc20ZpICbkkXx/m0UTh1wd+sGdcXMQ/SbNtGFj/03cVPXLAfIeL5glp58q
OoPdIm/NYdaTN6tKr1Y6vzOtaJm0Z8NJ50VcghOfp9MAWUzKwUlOx/b9erPnAafi
f40YcK/BQiHCfi3/MTm0uyPPE7tMjrWhEdJJI/a+/UzQfZL4f8/jwA3YSiwJtdRt
TrdgANYQUhIxisKv2cXSYTG32DQZ3RFgSyPpAT81nJ2JQrKcA2Zm7K2efWx3Ak34
hdCRU2lNvY/RhvV/k5guPoFOo5j0kidakT85PJ2/Cw4VxCP0BpPOdA+wM1E7xCLk
Z1PgU5sx8Mc0NAjJSFEmyFlzD3036g/TJcbnE3NypqnBWcsEp8ks/0cYWPC0gk31
9v6FKhLGWxta/pqVq0QxIST8yjL2LllyD+1aa05DSUQvYuU/+LSojMp2AkXw6vqb
T/AgvYICiwLqedYeFbHXeF+PA5RuTbOxfrb/z18hoEKwng0xJ1pp8Js+ZGZaVvF7
kutp9e5SJcnjGTGT0MhBgiHLFs8BAEwtwG4UUd/4pe1lpxu+ubxxYFrBKPj5kcgC
CWLjBoJN6YT1WWGP+shHCjaxOit06CU6vbavTTxq9UKJqy7s2csLhqZlxm5Nhsp+
56I4xRH7eo07HVHn7M40pVg6mFI6mV9sg8ltFJjoaF1XTF9+NJ+sHqPXuzUYg1O1
v863hQuLd+kSWEKKI5e75oZ7vgHkCef0W9Q0567vIwoQkep1sbws/78g3z8F/vAg
/t6aVLuntbW2s+1BpgaGYXMKSG67jj7uyc+/Hn8YsrA0mXsPafOwt0LyGXMnAcJg
649ZWe3wQXio2Qc08GsZz16WfDnnbfyKZ/jJfSYtVFOF3PnED63yQ0tzisX5akH/
Z9DxENi6qCYd2kmM4bG6LbfVpTE7j0r3lhElLGydORjGwJH7MVAeZ6FXCrpS5XWE
go9h7cjCa6hqOjIOuHyCsoKdR2sQZxLzzEo8IHJyOqUKEsRcUWPi2kKDmzAzoN5Q
bU1+GfV+7Tn/0L+te1ESJZk1GTrFiAjWQaHtk448YoRjFLWFQ52X6uhZuvUmMLXH
gja6h0hnaks/s9rCdYUbBrevGQJ3AIatvcMJN61VLE8XdRoV+r4rBzUcu3G7dB1G
nCZMif1WN95cAKHJjoaVEhNUthi24p083EePXAKrexIFPKQquiUmIAeoX+aNZQMw
y9ImpXThrEsxTwrqbeGCFzz8zHWqnpnjrTQQWXZL+fmPmpgB8lD30Mfw1X9s97BZ
BzXQlZsW17IM/k+JLcIVvjE6WfF/cyGM5TRdUj7llvjYaQT/eundaSFZPVv9EBGV
UmzlK8SB2IWqFnAfoSEdbG/6GkUkDoE0HVXq7SjbEJJce/FGhiV87C5Q0A+If1OZ
qWo1YHPXuACg0c2lOI74JbaJNTrudSJdAcIQ7lW+09PyammUSxBLNEh2MF5vIbAH
ztpx1zs8MOo9cKRqGNcA5R/PCuHRFYQNqejHViBk0MD0hBnPJr+YuxMEWjhuoYDl
MLyU7erwbD1NN8ptBv3YzCr2VCtSU/XU4063Zkvy04qjyiE0f45opn0n55hgAe7z
JDsp5B23Fw3OoJMUPVp5nyZ7Fx+ab7CyM5Mc8lesZ9/eulaPkmOIg0PPpNf+i/Xf
9BsEEpPa+5DNMDMFBRcU2YYCX9s78tvwIq2ivFtJBiS3YthOGPr9ME0DsWiGxTxC
Nl8g51g9lx0+QcBv3eEIg8Ilu3ZoRYmzfsg5vczFQDINBQKiRpGPT7HZscNtewlB
`pragma protect end_protected
