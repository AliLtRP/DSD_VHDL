// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:33 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lvCGBsYte+JqMB8JhI9WLvOi72Ed87izcfjFZvdSwp+hMy8OmgD6ncd8uY+FLUlp
sUgpxRdBTOXA+6Q3KSO7pVww8SSE8xPkglugOzyx5oNmk+Lb1yA4CVT9D4loO7xJ
dTDtXCr/24CfRmsX2S0LCus8IuNe4RfewM1Gxrt7ceM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28416)
AqMAVQ22PnfaZJz62vJ8ljP8LARgfA/PhInX2LZyF59EHxVaepCZ+o/CK2ppcfhJ
1q8Sws+nrZSe2ILpWufdjf5r8pDDLBW2U+Fpl4RepChsB7ZQQ1DzuNL67aO/Ywb1
hDqJ6g4NUkkQM3E466VLoGD9587JeTIBx/rN6U//3VgZRpt6UWHr5yIJX2pejNiS
s97936T/ZR19tlJNhs4MRaxd/FHUx3fmUhaa0V3nV95shohMMxaIxLtdAYftxDhg
f62XYUnnLYxkYjnJ2wxr5JlbRaWyghDbsENQ4iuHuuDHh+Rvqrw6dVrKm2o8QRJ7
cPbIQRDlgNZR3/3gTX1zTUGd9iiA8W1NwzPzc3oGmOjkN5lhIvYGalFbVWx6vSDD
as4VNEPaS3cDAWRPrdBgIL+hs9SpX+FwiBPRjJMNdK/d3SbK//DocLMdKV5jKaSk
yfVxs8++uR6ORPaoSW71nlN+B3Jn5UV7bokGz9IYMCbvSSJCYj/FepPx+uAkpxLs
FsxuopPWWQQXckWa6YCUP4dMoM+BGN4qzHcRx0sPskPWZvX/UIISSvEbHaMUTRqE
TIX8typzLBVTAHb7rhWA4igh/x/+Nr2uvzgXp4znHEFK2iQ6wvL8m36bywvQS1tm
dnQXqStVV5Sl7rAFSU5d+sESiBiR3uRumNxQ30RWOFTKPgYYrE0Xtmhg33jEN/Ow
phxJPCXz5T5d9Nyyux9e7NNanfLu5s10cdZkZ5ubtRyU+v8T7Cn+rJvCgOyeJ61z
2VqxFX8m1tiGw9d/G/StWTKtU2g2L3p+J+R4RuYbu13t1WlYMx28kWHcWsS2em6Y
ePBUbE8wxBi1YmK4c4Cq05wuT8UNY5kWApNHeDWf1ooW4soGRsZk/sP32bRprwgz
QybCOH4ZtcjISdmPN3KA8QPcqvMsXvSiffMudlrAsKe9GwHiM7MICsR+53x+kSsP
N40l3jwsFRd1J/8pdats1ym4RITu5Eskaev0g9eBpr5iLcaN5RkR+LDETqwYPzuu
GP12iuRHsnTM8D7mSE2C8I6qn6OMLBcmQ92gPlM6Yp4C3BqT7vyeWh3zs2XOCo4R
42KaYCj89SAhJPbcdUyq2n1TkZ59qhZmaXBUZGYFeJbccg+1Y7l3ExoxjQRqo9H4
gZ/686Gt7Sf9mxyyknxRWIJVdZ7cfRpXthlYXaWWY4a7McNJ81pkOk3V7rJySH91
k+XtL1CXn5dlB7dy05OEh7O7kOJzDK7+5WjGgrVk10a1QErElSTXXWPxWYwqtbj7
KOWiZeX+3vg227eS+lRNbFITSnS3vKzevHGUOK3jJJQcV8eZIX7KXwkXddTAl21o
9wI7+DgaQMDFMSKMQLE6XPUcRu7Xh95UC6VMsL6/wsT7DrXWyZEEu4vXZ9uQ42NT
LmEE98ej7pM2z2Cq2z9gKn8resHdfzubVHfNXZLbDYfUzwzX+TB0xTAtf8JwBhUA
Hqm6XdRP7qk2bA9vHlVMu6+gQuOZLlGFX36aV9e2uMXIUFjRrOPd0p8cVJNJjNUv
8D2tL3Nq4si7XVE7Q38GcSpv49M2BF19EAkwayEsBBvu7mTMP5UDYovW2fbMuDmM
iS0CVs3aukAe34jMhRbmhFZsy7kEntpCWDVWRMFEuwh4U7VRJ0pvJeH/TpyC4V6J
YvW9pGszk3qfXZe4uklVEtl965ACciLF0RcZULhqFZAXy9hP2H/YZU6q6AP8trhN
4/ZOYvdAS36xipSJGSYylDI5PeipIlC3/CUD/CS/dg/Qt+H1BPdWfNiam/Q2j9vk
moZ7QSGYmgwVtmhk60TQikW0+0DtOy7NYbHjf7kfhuvS2ngMPfpP+c8lhBYzqkAL
VKvYoRj6wS6zUYJGmtDe633383DJ0S62fqXvHYEbnTBgJbBZ1Ul/sA6PzWPchVF6
JXI5adZ9BrYYfrV0ahfcd4zh99KdRJW2UpXuRg9JsCKNGkXVqoq3l1dnDhPwKAfL
VdW6P+zpMjQg+3fIGUoJtyhYSWoFIuHoS/sR4MOWDlvjlonKKiWDqMecRUD5HDYE
rb8dt25ZkDOszYyUaDd+pKipN6MSQXaZ1+20MaOwLZpeYv1QRLOdHl6oRFr4uoIr
6QPYpyEs/Btjy7Nv+k1vwGn/iixWSS87V1Nxf3PDJCs8S7glhzFugR7KimRqKUZm
/qC/HZ84cKYJpjBBsqQ1qvyj9BqNjLT0bzo8EII+vyuOEDCa85MRTw6CmGvtSzPK
oydux4zfW8WcDKuAMkOQ6jAsvpIj93+jlDqCd1ReCWYgdeZs0QfdSiuQimAcfEYH
P3wNOL7ly+QGAf3DwFtFgtcyJR3y7RJ0wqROw0lZdaXVFxHBvzeWP1yvw7qHvALy
l4tjzcibB/164IsvNO+jKKyoZpowy5ZroWfVEccTXDe/6CnCX1icN3ef2emNvdWa
8OHQhMnIMndi1bP4Qz+YOKuXeODIIhHY7XkP6sGckxoRzOMf/i3HFrtoIg76Gjm7
yzf+2K8fuSUr+71SICEZzEYJq86GQNipKK5tRKivATWbkQJYqDeYERX1Y4+ieKQS
R3+jpyzVI8BWwm12QhR5vTOK3O5bImzuFnFjQ7w3Kf1Zbhh6+XomxqUywynMMoqE
F0wqipIxLlSlTTaMMUBf1japGK9/SguIBBfB+dpzmA4oUkAmRleP8dTETfLRDlIk
4g8r9Zyf+7CW6Wvey2eBkV4+LBnlLR4aoOKLgqYIqal56xfnyZnXVJ+Qx2pNsRSC
Ntk14xADc3l4zxSqLDdK5OPvUpojbgrBUWckVKtpx4MBf4vyiiLcvvosApDlHAwt
0146AUWn/TVBP5mYIs3bKnf7hpw9xteK/pEdqkG2wbBsmjwg+M7LkLnqg+HPtirg
qWwpTvo6miUw7XmVhe9pqOOkAZgts5KWYgXNIkpBr1Hs6tnECKzUXcsr8aqh538T
IrjwmvYyySe6Si4TZFKCjLq1VLTA3kNcP6b6XHcvxfZkH4ZX7BfPIavoZUgir7dk
Y/ly9I3Q0wcWo0RE3DVXseeI+B6r8SXRk7k9MBdifW3U/JwLlL6wZ2lEVuTzLxVR
1fFCMfihTvwnkhVU6GHzsQd8JugY4do+gxfAAbpqGWxkv9HgZDT5IG+4aerF4mDV
E+h/NUkd5pJChKZRuLLjje9B6mDx+0UCyXiMHRAbucQoAXpQGWP20gBPt6buUWlU
/bJJyREXz3BFVc2nFSadGcegse+RVkz9FXeNSSgg+yM+aKwv7bnkMvWyGQQZzads
AmRhzgNswRHrlE5LPLSRQAqI3h03OmmEXSE69O9ClYqiI2/UQ9P5yMAyrPLMoHpl
XdZqeNVoIBd03pZ7STZ5P73cCmKBPWeH7WlSDOBZ0XGxMs2z9epSAVVwUSFfoWt3
b0+fj1I3U2X94DrN7fgOrVV6x3UBw8g97e2zqw8tvEzrD4F9bbskdfdTCcTtxIoW
64kDhAfTCxntNiSeX8DpaHVUypRnfozzVRNnF3rnuAT4RzwcxDzcMlpmRb1ZMJ9i
vprPr6WnPiHjQFvivtyKb8b5tfrc+AYMCkC6ola5sw8TMmRePMLGU45dkXCbbw4v
Q53RCi7Dsd+yATfQxkFa77BJLlkj8QOj0/6p3ony0WgDxOhgVAtRBuPHDDD6HHjZ
DghcAAjYtcaM2t5dmEoboYo9UrzRJX4qKURpCqELAotFkoxxcKYBoAAsgQikZOpx
Ywkqkn9veDvaJ02e/QsvapdugkhX1tO7jKOQNVAym0p30eQf2YFEx1wHLpBls3q/
zoEkaxKvk9HzqBuXdOsS0V7aG9oaSHRhry63zAOGfjwFGLqvI1HZNSDyCT13GTmm
09yuE3SQRK5COgxji7KgQznL05hhguocHNIKvYqM21SYAp7Qa7rUynUeLVgkr8+0
tEm+Wwy67y+E0bmK3OhaLY8TTUDMIlgXepxZ2nTOW7+mIn1HePUiwwX5yXme8gPG
QXZKzvPYYhOLSWzlKb3kM04voU4DO3tiJzG5aztIc908xQiZrVP2loZExetW92Ar
3NeMxCJdauHyN0T2MYoIeRezeOuw68fWbewYZBKp71FldabIEe5hMDu1I73C1Gsn
nzHbYoU4DHm2IVbGzO2r2FnJDVayCyEAL635RGBDgYhDEQ/tOCm+HiUt0ZqJdaLV
2j4sjJ6R9UE/2avdwqssOpJZUlJqV9y0rIzKHcsH8hr33nxp4y6XKmplFfo4ETdR
avbANvIsowHmyiJcc/VgsXNC9KuS5u6pFh7+RAjcAHUngs2kdxUrGWfkTxTglj0I
Hr2zeDSPjG7VV11ascGvbN7dV4RbXRp7VctRFOLGqIWUgwg+8DiGfauh6BZXloq6
vwYvkDC60ANAUMfRGBICN4I5A4YQSqydK/Gbg4sr76iVOvsKPKoaXucxecLHbmzW
+sjCL6PjNIKRIlz8X5VbWYx0Pxch4NOGO6SMkCGkSms8haC/8+SZggfcvyW8as4B
4u1XlS4wYRlJXX/FYA55Xn40CdFFSniRGb46pNmdmRwu+sNd32I0q5nR4oyBKfND
IfZW40Zs0YpJetukEeNxIMvRF+4iiGFT2o/4tmZZVy3cX/PBPAOYv1uAIEXR96Ep
yLcMslX1ohqGR1x2nEn+ZiK+npOfXdddUuvY3TNEgd68Oroi9sTsQvKEaoVV6TCE
+domVcqbyadvWQVGjVFAjeTXhbyf1X5PNmzrYhu6Eq+oJD2UUvgJVsug97YCGYeC
ObQOEDyxmTLGnjrMX8p1P1qbCubnRlFq0uvUr3epyph7ngwZu/KhWQaO7mrMBSt6
y1oxr9t2WvyEKWwwOZYMXfa0mn+QcLB3GrP0OZlNthh3JOucckCgQ43kgZeK1KHh
YuXRDj+MQNKLwcrM2ZQXDEhRCMB3PvBdaAPCQx7tNeSgNCx8K0MDMrxij7fRid7T
N+kKXJalMri5Q6cZ+pRuhgada9kUgxsvorfsZc9RR9+S4nAoSkh7JyXMT9q+2zNS
QQFE3Fq2BYoVSSaujleMFc5g/S0l947YdcS5ja5/kVgtyg8c4MRA4QrUW2jCuC7H
HzbTuEv9YlF46rn8YskdmMf57DKI+JL3E4Riag8+QGvjACxQ80G0e42r0DhpWNh2
8fbLE98FqO2y5Kfk5ylFyaX3iMbL0nbljFmiJknJdTo2/hY0Nq+QeqQKMUKYDb3B
LnZimfSdVws5NfcylTRsmMrZnxcupAAxJR0/EWsqCFuKiEjIBE4qcUEC4mnC/CjH
viplUpJmlOihAhSaHLM7/wML0E+5apck/ME15PkiZwk7+SjBFzDKnrfTBb/s23lA
ZCgsdepT/ImEuALJ/fgHSh1ZkBFYvch11Wr9Wf93p8pp0zjZYPUW0XgROcqr4vuS
CyXZz0q/EOjtW1MmTz3pxRwmI19LK7nC0JlqA0WjlD+3jRdtkCFQqV21uhlayHL6
yvu8DmoI/sYUubi1DTjaDtBPWJKw2U1Ek+Ige8usZIdGCiiBsZJTpMCT8Nv6Mnk9
BYTvvxBRhkbQu1/M8CBUDAijyumh4tHNFbGtZAE6oh5xIzWPJTnxUqmbYdzDV/7T
R4mKhgU0HF/3AhT6cS3M+9WulWU1PzCy4zh0ffV2dc1CQHjzFHk2LqyzYONBA7os
x0N/JPZaIsVaqfZUvIqpt+kn3pn5Cxdh2bE1zqgKLMpv04YEKGATFPL1Wvw/+P2o
7w4ym1FjLipfvKdGWlwKu+z8/cq8t5cAwojYGZHGGwRUpDkAvaV2wavSaQG1EsCB
EjGQF/3HfPAHpZnDCtSIUbCsjbdrKyW7659bwvOOSZCugLxB/k3RWHfP6Ab7/eae
kk/62RXw+Oq3ocOO/eEpIChDwIXmE0nnehVvLwzGnFgahYzGzCh2+qsr0SKFs4tw
eWOmg6f0nteOgWU+YkSkKG3xNYyr6/Rs2rdNOfUd3oBDp1g/lKNveT8E8mFdJt8s
Uq/4mfalZwB++x1u3wwHV3lCTIdAf1sc7X6a+2qzpupqGuMlDggPzI7/IYVAgQVP
VZsG3e0Lh4bjrtIdaJEUd2+uEdJlnEmm0GMzJ8McFwwjm7UxbpDg/Ro+iSYnYvON
WEg0Cr6RymUtAn4NS1+3rqlg4c3IjUYf1XZyq+R5CqmsSVdu15zuk9vtkwdkDfAJ
yukCY+Hrgd/1ohDiqb+eUhsgxxLpHD9yqvicgJhyn+FWM5hL6zQZ4zvpZFU3WW4V
guo7x2defXBecgG4cG/g6CerJMd7GC8YKwUGvKjM0592mHOzD8G6o1dKOb/lIM5X
Mh3VqjrSkxlgfAkToCmFhbd0BUufnWIm1c/q+gRI4kOW1qpf55OOiSa8oU4JPlY6
RLyMweNVyNV9Dy+9Fo02xA1xwo+VV7EfoIPBIVG96kSsjNpWa18LQAdrnd/FFy9+
+exYZ5goJJE6cXV0Vxs/EVwdtXB6QMZiJ/vHyrmdki2SO5jUzOtHQQHYirp/eZ1f
sJOY8tCZkAlM4nJhfIopgqeLyTS/GVrPh5Ve06MEEBA9pi2knAeK+dN/lOhx1lGL
UYhwTzjT4qICsr671Bw6GkJTtJXY+yQx8N0grPgzFlxtVl7s60riFuqzx2hZomzy
Cu/N/3/iMHwbJKGOaejfs4xjDYwTGRpyo0RAlpZhfGIYexursj8hsJWUXUK3PcU7
R5JAxjZ/tLuzoaIHi54FCRDjZiuCgSEEkMJfp4kRwf78oUp2zO8XPNnWAih+WVDF
4gvxplbQk32AXgcy0KGTo6K+I83hevjk43HilpEDZXZSXti9ESKDHiLqrOX7ni/p
ojhFzajnuVbnCwFXMq6FJLAAnr6UYeTKO4DiUW95Zg5LzePHv/wi3HLJmslrTQba
HT8gyc8YYzqb82jyco32rHH5HILd68rSvCc+AzpV7a+u3hIkT06w8qFkaAzkoSJv
SiIU8eoUsYFC0ttrzA2Gj8uCFzE1zw89nmaAQyyirzpo/iOYjGqHbL8o9cHtKqvE
FCIsIymmX9Ur0//O17peVHIaNGefCzDkNkG0M4SQf8vEkF8zyy8IhF4PTadm23Pa
jsOqc+K92xEb787aCHl4cXchD7dKrVgq2+A7PXgqb7T8vQg9ILFEU3dyfpPOSnXm
/ulKJoLnMVghmspokPDiABqvtQQMLz+KIY/mCPSJY8kLhs2AE6JS9iPSbx6fPHDT
UOGwgc/m0F/gyt57xAjGc3nIzuwQeQsWIuKtya+UzfbXGBVRq6J5DIQGp/DtmHnc
v2i+dfy87iypTYNLF3bG+Hk5lctoFxr5QdB3Ot0+TqWwqUvBseycEG95bqDbRCMF
I5xLh86JHrIOEheOlgiUt6N0I+ag2EWNpASfwu4/iQq/n5+oqJgcS+fN7oGMAFMY
Zw9aop/k32Lv+K9S0f9KGH4Rb7CeIbIj91KT4ZJo33cvwL14b8Eycsn3m6aIUa8b
ThNcM5fiN3PlgEbG++S/Sll6rjmfjVRjLmu9dklgTtNdnDK+sEX2iZl3DxP9ZMKO
+D/YGGp8EzQRLpzvb40Ohl98MhdQ5sy1we5UfjCCDvkGWIfbdbEnXqKoemdPzuTf
/6D9MegiqhAyPqO3bP6XN3bl1Eg553vpvF2rowSngf1vKYuTJhMPIF4eseye/bIQ
e4XxGntDypRPu0xm6kRiw+ZdLplhaYiS3rHTZFG4pfsQdg9vXIpz1xvS2tu6p4Fv
Yaa1h2tgiZRv0ct+eJoc7x8T4HRWH5whaFPOsHjCHKdzvyIDFf71DGFjyvz706kk
/XKK/1XFNvze5acVH+pLOj7tQ1MBkG1USCYIunOHg+T01/9vCbj+n6YWhlWamGGP
rsJbBreeRz3Fv8zFpciedUWG3g/fLBGn1C1FUlxJwjnQj/w9DJFGBy9Ce4lPlxWh
GUOikNeWQqXZvaw/n+iBqcye9uXJrBizEHfbspJATcatpmiYNQ/MfSPHv8Pqa9C3
IggslNZcxELxPc3NCko9U7a7it8QegdUby7/D71MCmQDNQNeElZQYx3LMoYLLIX6
uyeCMflROtF/vxIGjMUotZl/1k1AcPOrQweWyCMzXCp/T7JPQThhwCHZuSEvBMlK
NAsH+mpPlUKunoQDKow8EjvaLxG1n56xKSjfA+aag5D6UQyB16qU3KW0ua3f8i6i
ovbZGXor7ywiXyTXK2e63mzNiM3eTxsKQ3cPtQl70aXalVNzVadhKQoErqxbDzaA
oTyA4jEnVyctTCwIBZiTA+duMP44syBwi7S7yfpd0UrrfX5NhqxdCbnaOXEDyOjL
4Bk0sCGpFvBzxgEpm9uzEg/pTTjb88ToWXqUq9NmdPI2YAqGlvSkApqfeh8cbz8A
TfxMQ546i1Po5//n0etcdHXyetasDM0hWHpHE7BwWG0xOGxEBg7um56v0z2Ia1n7
I46Kg1FeaWh8T9u6pfGxnbl4x61frn4dXkU1MOejrMlgAyDa74n0G2bitlZYmACN
FGWNblnWOqw7k7M69epzFetF4o3eAZemGR/UATgNKmyvjX0GWRzjJBc3QJ3TwaAf
0JchNeCpIrZQ1n5tPmB/xY61bZI7pLQOn65Z3ut6/OCOlCETX803J+n37eqUQhAT
YInk+vd9tTRq3J5eetltm1d4dWXYV8WbGlYJ0AON0Mtd6XjHtxHabIj/ey3EeRP3
YaQPUoGX9eudMXqer1Jr3UAdW5KUQcAEdsmf8sMFg/92Jwm/tYe1eKPhCcg8QdPx
CCJdlN+boIGAN20/cHTwwJiOAXB/A8v93EjZhZkBX7CVJuiNce1uzBVKhfmpjUZY
IwOc1FFmymBT3K5mgttc4Ixqbbe4xoLxGAequfaPoAtIroBAG/xAL890WI/ZuyNl
d1Laju6sc4k4ZWxwVW4yCkz5MJIMoo3jqFGYIVQ9qg0ISxxwzhKxp3hWIZmEcHmD
8wCMofeaGpLUhwS/SO8vWed6Y4xnOm6ALE9BtNNWpY1VFYen7vcXNH8Xzpxmof3M
kbfMPLO4KzTCyYq6KNFf2bL9eXIV9YKmxONW4/doqA5AjmjytStrWJREpRLZ7vPl
y+7PNeFGh/70fjlBoTMJ/0X7WHidGE/XXUI684t3GmqG6zkKROjyuMxHXbguOwDY
mmM2SWarAdzlZvzUyo/VQZ8y0FSitc0t7+O/3nZ+p9cn6KCvy5Cz6o1ZFsPRfd+L
kgZIhjQCdYOa8GmbTI7o6qUAB/5HTNhfqj8iUKLL/nVhEMNNbJayvpZhUz8Ehm4h
dKybVxTdexNfppfyAZVPkGo/Sx6r/zgtS486j6Eg9UxsUygVxpdv8DAtiQZ0eLnR
jWmnNDb29w4e9PNQ4XR6Igl9iIYmRl6FeieVUi3DoevC3tBa+gsiVdYEERvUv7Qh
osbW7wyARdJ75c93VuYjLl0+uqHiVzl4Qv+s88kI8j4HPvTtwYoVaEiGhLSRElyE
jOO9YOW0NnjYXm+eLbqYtY6nUH9jfdb5aDI1Srco2AMkDJ6gM0D4bqZRa11dJcPz
BapG3oiL0SPVuUNp72QlrPsZB9J96VqLT1tQhBU6DaD720F2q/WZYEJQfMM27QYI
o7dNmQ22ME46B5KKoPVH/hdXczjFOf83lENH0MpBSxd/Esbm5VCc1K8yU9JjfEse
PbKaTtJuu+nImMZNpH2xrTDxgngLwnOnMWgv3uMenqPJPu/vrkqLwbionNsGGZyF
JmVF/sYg9jO1LJ7jwAsPb3v1okSmOi49LXUtZWkcwrbo/di5pwDMXj5n5ZaQopj/
BzifdK5RpsO8NBdIXM+kOJv51ex116CrRcYzJ2In46fh1Jg8mNhh5lS8ySooEt+/
7BQSPOcOe6LrP/FsDPidX6p68ObtmED0XlGsVUOaFz6NlPIjdeGvxR8eyPdq3H8L
qC1xBOde7fa6pToLKfKaiWuTOwH7aNRV2tBVj2nF2HvHV7PNY4IDHBt2mWmym/aA
5YkgmIgpUzq/BQgdif4v9dQAeZTs01UDNWdP8YnZIPRqpCb/6/zkNHU7wkT/JqLs
A1ml9YjpRr+COgTFxsG5VucwSBCIHPrDT9ZHM+hdNskG9sGEDINACCfwTzeQ3WY4
lQh/q4jhWGQtUDmCgUYpdW4ETGm8nkglw8GvY+lxQTlDM57ynMRSUhfbUGBG6Mvl
GXk0tgH59TGbqNiBmRmaT+fqvC5ilXcZF8WlmIBjR/bJ90CcCn1S50iboQ6l6pmw
NBLr6jMyWNl/ARKEBql9wphpdl5uE7iNo3uMyfcK6Zkp16xnhAQhlxCHIwlOv4dG
I326FOrdeyofWfWpVnt2KjFL5LxTstl1ac+oehDdkatphSGERfo/T3Hv1n30N3sB
7l8vbNafUrHNPDgvtpHdB8XbpwVVj/TBPHeJEsCy1Fvd5/wdU7NlavENjxIlQ1Kc
2+0QgALiAd8HQ6NF1iFiAobtr4V4YFL6c33O2v5SiIXeLWNX7HVlCwf+iVhKDUkx
VuI/gsMuN4sLeRDOKukK5GpIUv1g5QGOLQX3OwFoTBSWCz/xsuIxZmC4JUSRBtS9
4O1kOFDoOcYqwI9eVDgUzoRM6R4G2+gZZuHjfZssL7xv/LQMi39r/puh/psZOUt8
34J4fQqkn4ToY7mkPQ8ymc1GQXdoY12vs97zIcbVS03vb3wWEqRkvverXjcAKLb2
rMRNfvZym6FK+f79GdiddlymRhsD3QnE6bgqnIowtqHmvUtxCk1y2TyT0ZOUWQ3R
CT5VxLgpMoJ8tSJP8G00ow2B2gzEDuz22uKoSkJK8c23A3YLx9DyX1fGxy4awA7e
jhvdJ0qJqFRgiA9KBFq4+4X3Oa1CyKS2VDOeqJQmsitZ0wv7k6f8DvMdD1rIxbd+
n5sQ9ebyIWMwAvvqpxXM7wGO1XuStRn6pa4zJZZN/aSgy5FxXimjDJJTblRLv6GR
R1orb0/O1DEaZVbh2kGALs+5xmx8/2KmTaa/rFGonT79saRAB6Tozf6p5NZEGCuN
/SNTYkH6dpezLKFJ/nxeLPTA6vf0hqQNHvW2LXp5O7xVq7Z3uQIKMLsHcQsmNcin
tnI4TBU4wawE4XfYpz31uaEootHVIwJXd+YR1qii7afeqoYfzq9jOVO68x2LVQLC
lscFiaFntcPRUt7A1vpNHo4qdi8tbDlWcUiNLAusDYv4mjXe3qNM91Z1hGqC5fV2
rxPi9a9QF7CwKSt2/hhiorhF0OR8fvcoRsUDh9OcOAUpXnz2pRg64WdXU7b5chUs
w1JcDqekgWQTz+NEzO9WjPU7Qu1ZJM0ounppbg4SYn+ti7y9ORyUU816W139IgtD
b9yrJWo2OJ33D98djvXkctcG8cxrz4eGbcsD07oXTKZOKd2EPUMET1K2APBx4REL
yw3Jfle6kn3z7BXZxdOSLg39N790So7Ee5i+3dr+Wn1Xcb0OmbyJeuBautBFk7vh
A1vUcNkUK3+cP7zWCE/lMrKwf7rqV2XJ9MyuOYr/O/b2GoQpbAb5iseNuw1IZL1v
uuq5in6YCTX3C8N0s4IcMNoCb/HLfSAIvuRSAa6Vg88ssor8RM/5dB7v5gec4B9o
H+7uo7qqun3MakBPE7oBc+jcdgFxlVgNkIVNyfqUhMn410tVS4LMA8O9dgoi/GJ4
YuawZneBmQBXryv3llmrbKVmPZDvlUlGWf8PbaNRaJEGTjbq2FHc0DpN2qItjULi
A1gCsZe8uus2Fmu7dui/snJCuzJFi0XuZHIBVPzFcJPmgJdA4pxbqdbrkE2VVU72
VdClbKHNnY4kQXX0AVriaedF4HvuUz9vzzttHzBXnmg5FhDTdm8g5IPxrso9v/wq
eSP9d6oc+Kp0H2XbBQaeNFiEfrFlOsu7yvVtfaAkc6wt3LBxReGx8u+Nb07Yi1Pv
kbsC9nvTgRb7PLR71CInjibrMlDmXYLYm+FVsUVpZlnipUqVJZbNTF+WP4CC/8Qu
Ry3A1NVCqYKkMVz8ztWA6o7bcKU+eoA3FYzYpfDRRQAxD2H9dCY9yUng7V7qdWtT
XPU/XAxLf9kmirVvh1suzbQMqpC6F1y+HHTS1KxgGi/JIe/VxKW8eqeralmvO2z3
99ZNF/hlhSQKK/t/o0XepK759xBC+H3IZCC7hwW5h2x/XC+OyFn42Zd99qZ0QVYX
pXRmdRrcY4FRmVFRtg1Zagus07fyDg9KrIb0YaWS5wKV1TGDrZW9jweRIWRAsPHh
LztKIEYJr03rZOZ+iiXKWe9oU3GRTSZUUu7t/3eZQMXnmNOynKwXHnfXGi/efNIv
LfJF32QNn2jprXEbsFBR+f3sK1CEWWPq3/rMG9mksHclM+QAhy5UtTH/TpTz6Ulw
pF773CBiJw41wv6ToFd8WjeRqPDiN8qe3W/mR9emk4v70Sw7qZyaYKmwk1LFM39c
pNIoG/m027KW9rFyV51Oy/igLW9napyfkFgsN2hYO7L5t40MwWrWUX8GUuV+ypFB
6pLXkhktQy6U47n3wWHKGuUZBMPdVUaPek8lvoDo1z4z1BDLNuaoqaQDO25pYdRM
tdBqLHieha1XnVpQjG1ziS8RTACqLDPUgS5ygavILZBVLgGW1623Frqu2hFWYXbC
2Ef8H8Fe4jO9NQtYFUoklIVl3XGe4PQZf/O6UI9YsT0dA0iSX0goBDEtN8YLJ5dQ
9MQZ5u3Du6W57wrWS6K4apnKMtMFgH37T2DlVxFNdEqfH5KBmDmLnAeaS+Yj5MpI
c7IzzJM3ZRgAiNkeLLMf7c/A/7w+e1YuaVgF5PNMf5vCUbytudfHla1EB9xt42tU
6wZr25WcX63jmtelk7pQ0Mv5015BNGMj/YrVhkO5IaRQF4okawJsqw2hEcnugcML
emBA60gonbGd3F8+8tt2hvcl6Ma7VwbU7r8NhwpIAqi7VJg/wIpyfUEk+r0JI3xB
2V+dPm3mYijr7CqVTc5BWldWwJnS7GorAadHd9tAjQVfMq95oTsfdJE8m38EWDt/
Uzv5FQceCUuiOd6Jds5h6nVjQR7opDXi0WLQkzOFVcuyGN5qBmHv8XQuLByWnHz4
F8NCiCyoNuyqNEPHWtMfqYKD5r+Lz+T41oCHbMXDHfBnPPZOfe3Ix+alSB4JJdBr
cwkXuRDyga4Hm1D05+vrsvs+9pSAbSz1mrySBGln7QccLEbMCglEhmXbKFkBj0XH
2J5giird4LKokCtDZ0XHmv8LdWbel1huuMTIaIC2vlPrOqpLL4xgcaHkKYpikoY8
BZd3no1RMdT9qzlz34vmRayB3lsK5SF9svHjsC9IiGAvLwXAe5VWulwFf7/NapOP
e3SYiZuTMyCgpnRTytzsVSt5g0yRET5voCq7dDqa/wUJB/EUKviPpmDHviZ0lnOf
0h2UWVa1XmrwoUYPyAWA7eQrYkCQfzWGWxwM79sQ/1oM/qdOh/M7Fcx/HwI4R4OI
9lf0SPM5k4QYjXMMIyZBb/HZMw38lyMKvt6joI8ocW/PTUrsFKP4ia3TE9TMnFVF
V39VdQdfnPTWl1YXXrgKoEIX5xTB3o9kYr+o2VA/3I2W4IvsxZOB7I17qQPLOnuj
YfBfIBUwyJlmLwME8I8ZPjCcTezlALvZMgPhpk87vQT8c8FDDKX/u+9gpetqhSBU
KP5YL/Xvj+Uf4tdaHAz3bP//JIZeE95d5BQDQgFvEJAhU8JvAGcpNblSsVmomQWp
u0ZeuM++qusax/K83Qv/bwgInyR/UZ3I48qAFqnmgKaJpQvcwjt0Y4UKLvc5Eqh6
muFf7SyFZnm7MorEe/XKUsx4/12J9samTpZMwL1YtAx5qxwJUzy8RVqWq45mw9Ua
8JevbxSljcf9h+eUUV4slqf1hQVNrR5qghRPKVbS5fNsSLhXbhbio3QNIUdKI/jz
TRMEJHMGDVbCkL+oZxkTd++x3x4iTftiLtu37HvmRNBXgs0QM9GSA5rFfCIcSMtZ
kL/3vObTnPVQFl5iRpgkt70qJRxCXMmZDpggzck5ExEcvvIVo8Vo4fSTsv1Y/Je+
Sps8/MdH97I9BSYIysojSMldrYyRENsUXjxrs5wzduXyNixywfydZu1rsI3EZNpp
56Wq3weOCJFkCyKOtrRIts6kwFYg7vnBuJ0EotoE10eVwYR9xmtQTWa4ZnY461jf
vureREYS6YOiCzDzEeTmAkdT64Gml9gAet/vkUhGHUaJDXXH+I437cAldlolzU7i
C1k30x+03a5NG+qrnMbGBrVPcz4AOiJibF4kgLjUCENq0vk86YLV6qqF3BxzcSJY
lblwA4CxAf3AngQhtr/XOEe7SutN/7Si7ORxCbhbMFK8pc9N//oKF81R+qYlzK/j
f+pRWWEsZrQmDi7xO4q9a3VZF0OQkn61jXtHudTwKPaTndAu6XbRO+R7G9PYdIpV
G6OBnXRw2I4WPB50mI5R2IJ0JsbZqKQDDIC4M4m8xtM0gUif+QYcCp6J5ZU6ORHO
L0hZB035cEsvUMCsYorscPaSorKhqaQJdHtFcm2lcxlSiRVd8UxfIYAzQqMc1rJb
8jflFgg8B4fX5RPn4zRja+Cr1CyYAbhHni9Kgz5Jl3s9Tx95T+nEa7kke5O47knD
DjTJIBW+l1G54g7Qq7jInhjaxy2E7E+yBI5E8SFtuGdeeVUIVisC0pVX8PTnNMrZ
XGmtNoX58I2eamIb+8K86lHErTH50i9BWwUi2XXmy0bRKuWeS368+lc8j9aIKcD+
82VmTUoxm/uT5UHre0PCYNBK9h+sg2mTE9FbIKz8DmE47ENdwjYluN3G9uYhV4wx
LKTBQXZJqNJeei34OpeLQOHN2jw3okoQHKCdvPrAgguoEM9aILneY2q54M4BE4Rg
/4Sup9L1m4dxRO1jIYY3JjwvBQzUl7k/01qgdX0xx1b3mIM93pHLtBwR7+GVOOrR
rPpwX5DtF/3vOv4BOCn844Z+4GX8aLlCMpQcawXDp3jP9g2KB3ZHjytcxnB57UXd
AD/9urDpV2Nx2kjwIut1RyOdplmaBDmr0dz8A0ZaAvXVoXTGLusUMVhkQpaofwCs
7H4Tlctn+riRlvKUmzeT1t7fUP+KDhl1m5GjwcJeAxytxh5FqikryA/2/7dFw1tb
wCOh9ehHt6bsRoA55R+GSg96/SX0qkmAM0VOjVnUDQZmst45SWQkuamUDDc72kFA
oYgGqU3OqTpIZ4l65P7GH2s3fa0dPL9kzt+61tB4O+KJ31tJp25SMHnDhWuqeSHl
buplQOMHltsIgGKpn70yBXuo2XnCPfdUTzGblH767Y4M3Fu2pPbWxLFFQt3Hlc+f
UJsmGNsbvLmUr3fI9WARAi9TPjyvv7CRWQnmrDvj2DlXpf+ci28fAf/+TItuG9xF
fwk5MLYEhu2mH/Kk2m5C8oKjIUfuAC7htS7URppXQ5apnBwLjX7MdjneVTIUEtFo
mqoyLeJTu4sReawlOB8gSFsOO8KTq43UICydYhCFvB0WXSOnF1/ITeoXmYDHiMkV
GMw+cOF0gVLUB19i+6LJQKnoeKG5yys3KbAgbZ8Vz16Ufk9tVpfd/Ai7Gps72fji
P1TXL0HUhp3QFUH9OA4fl1H4AkC9Giwt3ZpohsK5M2psByDbU9mFgobfc580zf1h
5othqjdC0fQOfciry9idOK/CAwWEZuYXG7helq9eFHZHXOIp6mMu+JfmeW4V4NX9
52keqjnnzurztvkPPiflOEAwRpiMU2ifjS6ppHaH8GOG1kJpl+AsHY04D7wwxGUG
QbrwXwrK3P6DL0zdkURjMSnYAeoWRYkZbT5S+ij2aHOs+0SFFd6vhU5QhaDkXpFG
PhD5gWj7vfVbZrESeCctoom00LCSPFylWrG6f1ntGj8HiMDswWdLIaSbDcpuYUia
nt70E9u3bXxzACArvVSwoQOQmIIuI78acvdlny0e3+savyoxwRf8i6IIaddnR8mD
M+uQBEpmiQUeaCLZ4Z7bNfhCOc8DGHYOSdE3VGgrtZ+I5mepLKoqyWOKyPPyDk5D
WAiupLCmi5jF8WWFB/z3Q45HI3OoL7BgRJtjluURLLvok1K6Yw0MFePxsR1W8uJV
79yhDMyPuhL/qG5hZgrvkBp/ippAfibygLptJKiNxeYG7InkbQ7UR+s868n7tqmA
4kEbaQGB7n+hGuIrrKugPhkJ3XngkZaNyEkAN0DjIgQh0ZLQYnFVL30BMleSzjzE
H/f/D2aZ3Y/lT1UfyMJXJn9ADtDKuVwNMd+V8PtxrFh30zx7kLrOlOWJHtN5DUA8
kaiU/psbE71kAVl9ehm8E8J72XOSpU05HHt8Wehsbg/yiwhEeMIUmT1vauOJn1C+
YgtDW8LAf2D1ZZMVQ8Dezz0KAVnavwtJkJrxp/OllHqeLmFm3dzZFjCDF7pBhPhS
IgILLD/wp6xbqSvZ6DfToj+CkJGdL7bQ7unNjbDgCQJLyB5NBTlTkw8WplSmPM+7
FE6w2gFKDyQlgAcTfGFt9vr/RqFusIF2KjlvpJPcFqiIs6NqTkh1Td6IcQ/OKSKv
xCozp4tXpsZpWntTS1OpfXWH2rwZH8eOV9mZJq8PCMN/Q6v8nwg5gHHrPgSC/4BO
DkT+pjJwH+5uNdccFDY5ZpPaQCkuXpcuBtJ5FDDInqfxcSTyy6vfRewGgG4Tp3LI
CFCNCsBfTPoAPdd+slRfVkJMxXBekEcjg8yiyDgDEJzmmnlXFN2IIMgzvHeuUz+o
LmX0kkF6DwBXQFB7avzo8IQ8KiKf4K9WPgEm9Z+wTVJZlVD6JvNy+A6rzupKHSOL
P8luJxAY0VF8Z2oCy31aDcOCsQd2jOK/7MGJWYukfsXpGWkEbyw+doNWt9GOFXlV
pR8oyW8s610ZOp/PBriiSNjM3PmDk8v0S4wnDrSOUnIrVSRhZFjVQWhCBMBlLxgh
MkJNt5NrzgvbtUwEnMX8VxIs9tFxQvl5IPiFxisrX92y1mW+vFN5G3VDCnEKqD8r
Y9wi/jrhwc8sxURjVE3qekfpuFuGrCik4D8ZTlbfuVcm85NlNhvurvEHaG+X60A5
SxKRrLiETJ1kspNi7bT8lnSp74rIdRFr+R9vX5fLLIJ+aGzhvdSeok9hpDBCPsFl
ZmE+xm6cQmOqJBE/FvPnHaw3PQgB/yJbG6v7wJtWep4S0QuMG1KBxybQyXHDcTsX
aabtiHTnalNOvNPzSklOFcXgpTrn3kgumqr9J7BRnASNMfwHtkE+A0/IeyaqqRdk
BAprjHxIf6eo87Zc7lmmXKdO/x9FEsJ4gPDQPmjeYIcXIgunzRE2LTwyQEXr+qi1
3dpRxayVm5Fv8UMlhjaOnljWn9GO1twLCa8DgRsOC8cQqCUTKxuJV+SrO+J2twCR
jU6JzJ4fuEt3rTgIBDWSLSFN5gASzTnl2JS6oH2mP5eniaSI12lomPNbxY9RlTUb
B0xYGGw669xD0HMj6OMM2j4jgUabemQRl7zaPtBZu9lkk6Lfpfp7gdLrst2o6qdA
MRWJR/lu+I/LRCutGQEAvkBJx+draIIrEnAn0hKEPOwfF9u/Um02lCn+pD9xQCWE
+e1/GdQJEwEkMLaLrCTaxjTosqK0bZ6+h46JU0T55KOlQyF+d60Fr96JBVItPMyE
gcfn6GBGzDbFPva320fvVfGDY7LccBmsWHNZdSshQLKmkagP0o/RunJTYyKsJzPR
WKtLGcn/uIvYwm746DwM7ixpiUw+uhG9jCOJ+mvbfPsX0I8RBNnHx27a7NVDfedb
L5irxpazLUbnbRccCOOO/DVkd6/YnQBHn2fuyS4OL7tLChQ2l2BNqenKCh8GJznH
2u4dv3Hl0XuqfHPYEKkHqQWCk7SuyExouZtx7DSY5g1bNI/Hjk41YU/R9P9w19ot
iQUf2TRame2vnaK/jWVxvxVnSbiwFnXe+bFXAptgf59hjL/daDMwYFTicpCoa+i9
i7Pe5y7QitJElBz52tLSVP+jpoTrpTkh3VCs4rm72jBrGbYeaTZ2Wt7RK3jwmlbL
Q9S618fCNvgBunUUKWjx6MrLuCbLJTD0LfmHvKx2DHpkJjDjKRvNosqCUj2ih6uQ
MNtSPSuyuIUSMaQHAbQjCLiRifH7ctr5T8cRd1zUPh3lxbnBQFz/xa+NOIXJkNAT
/pFqk1b6NuZEaw8KQ5emRDz3wgcBJt6yUlmUKs31YTODzVK4N9rK0FfA2FYgVLPp
vCObGaaXUm0XHxVpTwdUyUBYE6tlcNM2ZIzmmzGf4cO8tw6j6Up5M4cTImjEBRwt
OOxiCdnd3pQaTFu9mIOTiprs3Qvat1no7fNA9UW0miMIWKdl1BmXv34KHlHlA1k4
HQ3WwtokCyjrypecdbuxbak94EdwkR89h+2YDjR6OJKB0u4PuhlvjgACPOiqQzEp
MQ0/5ZsqaPA57mH+WyVunEFMOG26ib82xS5dZC2EqslJGKj/u8YAJhsidEb86Hpa
UUrwR+34tGdJEEelFmsVJNrQ5gxlbRz94NAIp91KiDtkn2Ou+FP5SVGH5npLGtCF
BP+JDI89Qee9YEJS47EMaKKwa9fkiqtuQrEQZaOq/Oig0Ha5dD0kg4Iro4YGB9EE
ODtZ/l1c1GOkujFjHrNeB9BVqtqnl2fJwRJeoL310arZlVzMz6ujUz8tVVgwOK2L
1wMvGkfPMcZhijN61/CZW6fQFcmxMCGvxpNQV3IVodtjnFHkwNxGI1M7rx1a2MXU
3g0BzAyJM4T6W1ecBQCWO59UIM6MAr9l7+9r4xU9UYDpiy1BsVMbcN84QH1CJhxO
mSZdDwE920l1aP9vPc7lkCRZfk6P/X3MeKUMZ/V9pW4wn8jiUI5qo83SEPaWCzxC
qwU/bK0AMa0gqSEybZNSj5l2/pxjWcPtnNl5sRMQ+deaD82YyVpKzyz2JaLm8rMG
e/gLKyyYAjUYVwTFu0+Vh3A9snpy2D0U/yUgb1ArDAbvOD0kPnc2Tz2GnI3o2Gq2
Po0hGa7awD99I8J8zX5cG/Fiw0NlCzc5RZjdOV41Tbkuhkoq2/uDX7oSlK16hYVg
3ypfMSqhpzClhP1dd3TOEYvQv7Jpvq7ttdAclfld2PbF+SrhC4AL/ScaMOatVhL1
oTJZrkySXlYrQVXAAXoMF5UPCFuvTlR6+0toci8RhNtKezX9th7Gp+i2laxr5wNr
gQMP6kl0WaeTu87TtAzKU52XelLAUbr1QlJIV3ksadrZvCnsBzxQwCIZrmjLQTDZ
j3wJmgpag0azWn9Ndo2wOMo6f5G1JDeMar5Q8PtWjFihXQcAfiRg1mFsn4Hx5p7Q
Sti/179Qj+vdSHt6/Bash3QzO2lqiqrostYY3EiHIyGaaO4B911EQd4KYIYvVjo3
EPxHK7t1QUsFpTItX1Blg02+XrQoRzt2gAv7GnOzvMPXWLFMTdC4vuc7ycuAfHFz
jEeOm66zmih1r5sodsLHty61QSbEII3O60ElWaCegH91ZzRdc/wHE1xPzVSdhCK7
l1F806FPfkXw5GpUMxdNYV9OjqQNaTSJOWWs/hpU6payldYezomevDnkIQL4gF3d
ctE1A9qVw+IKsXyFf7yGuGFO9XVGisFlKQuVFDfjWUGdi9ZkhCD3ocTEpCrMrcrq
VF5MT5DH6qzNOs1CSbNFFkK7bEoYLcpQdevPVQTCBiSrUaup13aSTgT2SUSEuj/L
tL27f1eweKSbM7CFXFZKa4JePo+qlGSx3RizohQS9+QsIQVYd6U3BpDopWQJTs8Y
5mRS7ByruD5Y11xYH7iST9Flevdj1ubt7NUSLHT8vstzHRnNsYc8G+eQsw4l8sN/
TkjZ+oc0G87dd2R0ZqxSgRe9JPYIBdtdBGc2C3SSVG4KP2oaaue2ue4HgarXtEqX
KgsqzkWgLqxPfFnv0YjDo59k8WeLFYqi4stj6YsqarNkdH2lGRhVKyRnPVyCAgsL
gbt1VVe3SxlnWryAFTqdgVNuKxVEzuLbMS98FpvZq9Mvtklih2vOp/dLL+58PLbl
YLJScN1QiresffeQJyiu1lNamdsYVhE6afxus6jZ2NdWNRSYTjFGdigjz3i81ZHm
miEOJz5DAa11BQg6F1FUe8XAzL1p56atsygUWIMNfcLcguO9RKI2m1/kaPcd6laA
nftjSqphLMQS9KTR5POetmxLhTDA+nryG63y3LSfKWjFLgOKPlJxohZd0AjaFY9W
H/RnOND9dprMFfFgH7M83il20rJxrgboi12gP3QobUSEWRWPVM37qNKV1rEsblsw
Z/2hIXdbS66QA7/C+vOvJoRZqxokVVIhRZ7dUBfbwhicHQ/p6UoFT+2UXucEXBFi
FFwD+4NDEc+iOo/t1lwtJjw3VmHdDkbyhKqQ2eYYRsu7++8sws0fiYTQ+Z9PyOgt
3VmQYx1WgHTOwn4BlLI0V4UySJU0oEGBS9uzyhTyeAuF1Oli/WuCRccOntVUHSto
0qotX97i2Y/dKwfJXc9/MQ0uKsXDNMhG3pUQN59KWhiKZyUGIYBkgcQi5I7Lvsp9
0BC7/r4f294Ya8NEDqX/UgryUKJwP3yc2hPWTu8wxmrPT5e2THvV5pRPFIVmVbQ2
Bs8nwJwE/pA/2IKfHT+rZbtHra2XHU066ZRfNz5Aty++K7tpgAu5/cuAaspOaxcj
jABGqP5RjEAxjfMQd05B5mXxz2811VDeWT2v76O56oVUEwNeMxu8PiruyMzZ5+GE
BlzmFykBUwfd/WqCO07NCUtmyZrx6Rt67X9gd3w+O/wxjy1SAL/0iPhZGzaHZofa
Y4OAZrxNBG19ReqYSOxeHRA4VNLykbM7e0MqBTc8NISQcXyATe7SLPkwVGBvl8VT
PdRtfS8lcYuqF5FeUFPGBpyQlUiaCZMFE/Ytwu/ixfy1tkZy6ut+UsSJzvB2yegR
djhLkIGTkLn5B4NaDgO5NLPwlrYbWHD/u7dhq/rivdgJlWW+3K8vVeIGTYyseb0h
QKzdIkNv3M511fDpVw8QoKlg9Qj+24OU7Gx8dpvvzFgogo9K0FSJtEqRF8j1hqJK
VR+loLWB25/A8z4HWV5YwOE99wk9F05w6SVx/f/vTXIGbUsol1Pd0UbuNlVQCrbo
NSe0YRTBhu3Ezb7GnTgf1VRWAG1G6S3kIsI5DgULwSu/w8zHkQVFAZf+sBHdRNFE
5TkrwKRzVbON+xks5T3WyKACvm7rtwTQEJRQT1EJuaIO4tqs/RGsRVQAaHsBLVEz
TrexnGbSGuPl2PcateXtwPwUcrzU49DvhTxSZYFXE2sMf26ABK4nzDVBl/KTObmp
8e4cj3+GgsGEM8KYbGLMv1xGD/3ZKEvZPGuo5W7b1kJCfN5X/GFLdmMk8ygvJ+2h
xYd9rQ1aZntlpAPGu1tWQbMzm1e3vJYRbx/++IUMrHOFO8VSJ8m9oBrMYQUKBjPn
1GCRopPn2mzD5gixBzNKU7wP0Ba+lQ8/bsPTpYNadawtBjaRvDa22PMAUtg1T1+0
5/8Z758NGmp0AiY1//O88wc51SMhsCNo0T1p9gyGOwpXTlyIEpLe7OMnbtV7dTpF
Tpi2WNcfJ/UXlHSskuHbQHlrAZBJORWV0V4vlaLQKDoRNeUD2LjqdW8VlLfhJkME
DBIBnNjuz5dWUNWodCh5pJQmlAEH19XqD15FOvKQiDhfNFMK3N6cEckOZ4DpxP7Z
3NY2equnbPF38ThXz/Y+XIdP6fh819lQu3LHIrWOB9UaPMRuRN9g8EPY6JDcA2OL
WBrokeNsgbwkaYtpuHUv0qhsbFylGpvF8lpY5Dp36K5R5QcW2H35PGO8cjOD/DOB
RLGfSabTlTl7Km7dayZ/d7PpEyxhJAIVGjiZheVTq1d4Bq6nrRKfBPJ/TPe4c89a
zntKxds4zHy2CwssK5DtQA3FPHbVzc3OXguyWsfb7VWzF5wSgZE2i3lxzgFEOTV7
r/BkAdAvuWFDCegNVuJOu8ZJ8TCEZT3Ws3h1GhGxDu1z1SFwjB+hsoLXPGYOHXl0
uf0xY952Fzuxe+yOkUoYpVLmWsw34t6+82ALpXnJzXOZUE4pyz69O0WLAzLal+nh
d9WeOHD4y+qUsk8L+ct1P8ileDS6/+8GOq4WObTN+TNeZlGYv4ide4xAoC2MJZbT
sshO1EvnzrTPUsak/a6qFdhWsiEqeOXeQ0KPFhuOcl2WYZuTSRRoC4HOXhpxB8/k
EhMTlEVjEyy0RMSwWSIKs/e0PVv3BmG20+9JAfYR7fKtxoTteKZUfZeDpjmJSW5J
EHR/0yJmVCkCiFmHIZpum9VxeliMO9XK79zwVWHEMxXKUIqq0fUyJNbQOiHKiKqe
nRUy0NoIDl59wNk8BgbtAEC4sXo4OcT8PbMckwkawAKmVf0Fqyf7cJHmui4/lMUF
QPnq3M8sh3lKxi/ycRjKAvMYLjLwSMYCiseIITEuOAPXpNQZFJtjFXOAKZGssCFe
h54zZX/rA/uIrr5v0mfBWm3RBuSz8GfiZEWjFIk9TPFajP+Zs/hgwWTHMOb4jwq8
G+79O90Rl18reBp2o1YmcvVxHH/pVQiG7w8AXUmFNyqj5Bf6ycPaYM5ATprPU++x
T0WLyfAg+bHR1jwavJFlj8rZ8S1dV8dOaXHiQYcExsKybIOkdkj7fWHXdRVFgbS9
ibNgNY2v91oB6EnaPPzueSwYpR6FD/j0yLSHU83aImdk/Orts5w1+1+bCIfUKZbz
CZ+V/0R1xRD+fJelOBOATgPEmNA1T03jMlRNwPnXkZvnGP5mzzmsR7L611o+jisw
/SLBqHVaIbvtfG/V5gkKFjIyM9hVXWlAFkkHchVAiM0hBaLG19w6Pt4N1zSolClm
53BnKNHnaifFylOgSUodbid/bNDEu4a+W02rKrpp3WRiml/t0qglt73VQ+g8Rbny
yogqboQhW9TeKtQzI4yH5o7fQWfIL1JXv2MtBQb6rxHTVbT/WrrBDLq4G1m0Gkql
RYi6g3xgXkYFJrq9T55Hsa9EJIqMuW83TGYSyAXW5c4uA6iAa+b5MqlO2ePuwXea
lWc9Xgnwb6ugbiC478nRyua6bG4112LQklli0VHXIimjxvxXXo9CUa81ObF7Ojs8
E1iUeXVDIFZvOaGLZaiSKFYryAx/yQUHgoDyuZ4frieZaMe/RR+A+7FULmRdjbir
ZIUGtfRf0MNkt8vSJ7uNWBSLxh5LFix8KI5S6cE04TWgzOjUn5XznEFqRgGHeR97
jqBdhj/PYv+xK6w/baXZ6Bs+3r0Z0aG0ww0Gfw9UgrIbEU8Cz+/q3yEve4NkTvs5
wSDolHiI0TkNTl233yQn312qPL8HgOWBYzac89cxfwtHTimNTb9s9rPrAq2Oavwf
ZTS5U5uQfwi8LrV0NuZu+f/EAo8M2XjyzDkMagMU0ZP3Ntikw0mp9zPpOgtfRQD1
OmjuxieabGe7Sk0TwHuEf1HI7Kudj31EBWe3CSORsivMoRafHwp5R9QmXWDWJp8A
DRqZdtRAvp01J7nYlFEoCecv2032Li9Gm4aUqqrAm7deacUyzjADr2wv5rGP5PIt
RRy7CJsmiFpeaFg5xvSS8Wj/XtiVOr5rLMbrG/VN46J85OP2zaBvOLnvVXjLAN4j
sgdS2MGTiJgu79gSrszP31X3ZrAPyQiBnaDhzhHcYFBT87V/h3dU4KR2psaU376f
GjoEMlomjBvOLRDMxLplcaT7rtv6kQigaFX/X7jrjucM1ALwk+lcWUFskYSC8yX1
T8WsP4/xqOBQ9AcY5Qjf8dGOJTtv1FpI90jKJBVn5EjpxlOouLRHl49LXIz+5sC/
9eUKwfEZ+OagMnzELY+JzGSz3X1rlwq8o+wbjfvgSakhgjGtGhkngkJMmVxyanB/
glr2Q0Yb1wgbHTracpGM+q1H7QA28VTT9jkKX/BKWq+VMgIAjKaHYu35H3Tv+evJ
zxjs8eQjpdUTWC6eW7XgqP3Wv54urdWOabXw9Uky6dHoqYqONC4ydJ2m8ookYkNZ
pjO2FgEtAo+bTmzxoEyDg+kJ+eFL6lXSR6PTav2PSz7ja7Ytnz25FRbKEKR7q8OS
x9H4K1c1e/2Km0plz8Fpa/ShP2nxSqoXilFa2WQJAE6n5eMVkOHOsthX+QfKLRaf
yD5412A1lPLyKBYlbBH7cvnWolUs2z3DE/CjDSnIR0UsoGEG6LjgK6m2VI238439
XhBeUarCgTQT6zhSM45zwYw1suUlZj7C97YuGgSUYyHzUVSKHqkI3pwmp3EmniHH
y5/Hccf8LTQw6ovZ6+jW7TVNx1cfBM+RXTIbpZ7t+zJrmz7zV9ApmHTAANJYcyda
VdECOBNwWgDOPXpq/b9RTZemc31m2ph3Wk56zmlT75NN/PvycSr6uLQJdUxnx5my
GhF2LNj7Q9+VfliXO1HDb16b6s/3DaA0zKaXGE82ReouVR2OvDNaolTHMooFblHV
LWHxQZylUrlMZENG89/HFL8pDWCi1OC/p2emWFP7bCx8mbu3qGqH/uCO1QGhmk64
IaY0iFIhemrx/6FMPOpTeQhbqG647D22g6uIXEuw+l6wzzHW2BaAhLpVcNgewWCF
DJyRtq2LZJhgmvmgolGib8b0+8Grwmm+HgN4cDz7o+nnzpTr4KU+N+rHBACrbJP8
6NJbQ7vh1l1bscFWLiA00OdG4HwqDWTHoFfiVbfrLWJmZK16WuxpYJ28zMaav9Nc
uT6CKQEuwuMZyxBwtHCmdGNGBp2i4H2xEmi1sVMN5c7N812pxmpLXRMU4USfVrSz
ZqxkxVigw4EMSLrGHJc5p4w/+XbGapoEjXaeirkGNT1KHAcSb6PM2wAyZSIyAWpz
qF93jtfRrYIQ36jcugQ4YMI+gFDsEGJW4PNkI2iqVGQtfz1roNdKVzeYkC0xPEDQ
NW9+eYXOugddvnV8qI8cp9g90IX31fI/66TBzOnmVqSR4uDgZdpGq6IvfOd4CAsX
W8m1fxvVZp07MshitaxxSJwB5S1kPnI3qQh89B+nXuvlvuj4is8pxu4211ysbs7S
rwU8DRmwFMAycgImYDAwgB4NIypxBwnB/0rfvhuGyQVQRIUaO+2dS2SRdC45FkII
7eEDHzGo+mLD5QzlHknxsxkpfzoikutY3gEKUXrhZaNh8SwYaAqXVGc4VBAg/7ef
Xu5pH5epkr77PGXf56tkbSWW442xKjhJNVURSidTAUrQQq2clI/gZnDj0SsxVfzU
2zXSj4pmQ53/OUxL/p5sh2pD+nqSbfxfiwxC4oMzRNGc4jcyBbUzbW4AaqBCEQmb
M/DqOf4BQRvTfiTTBT3j1klIkEm1lL4rzGN4RfMkdY4SUH49O1NqxVpyKcuXPHIz
x3ZE+sDg2P7WmFL7Y2TmAszV9o2ajbwXn309ZQZnUuqNnQaF/FFP9vBB4cMEBMkL
3TGYbNinLwyRGpIL+FHT509CEDFkHsvDzk5wgTMgNSWGiFPpEtiiNkUaeCmAWYVx
WaskRPPjQq876qwmZzSyAr+G5olakwa4paoY49BbIAc/etTFpSfOndI6lwo3KvkV
8u6nclZm9hZIdH83nMVZvcEaTJZq6QS5TTSuJcLT28RA2KtwVVbbVkCNk7+x3tLA
DMbJ7k0t140nXwolRb/XnzA+Afze6HyY7td5csxGXJz2vcOw11UD3n9H0ic9Qur5
kPfcCKoXKthYFis7Sp9wSEL/BHwIR7EOKfGd9Gktiqfq2Bx0FTeNO9QKP6mYsij/
K2SpW1HrEiZnzrr3jFl3Ta6NM6TkcxMf4VtTI71FT41IXKDH1F5fJzK4pL0bLLH/
aG23b8HPeJgGKbEOHvq9a/nlQPQwHPC1SKOk2rktwJBjvFIpisNUaGFFE9h6lWe7
j2y60jw5cfaj1J7lgSydDcaQukuoDki2oA7spbqDD4lzeseuu7UCkz1j8HulKJLs
wjG6G+inPpv1EcnkB01Vd/w7kjNDR0Ek20dSVFgDk/I5OC4cGLs3v62kKCxvzK9/
AqRViEcZr3uIWhOs/pZJsqHvXRbzLa+P3xp344i6A2Eb+kjPcirUy8ZNzzGGimUr
UGUqaYguIaA27nHWHbmyFDUjWw6uxBVlk1tul4iD5E5GI6s7gb5eglrN/uI5RSQw
vKgdLw9zLo2RKJQ7Q8IuaueeukNE2MDP1gbn1ehHPYnjdKWBqS22MiZn1m7d8d/0
kn5qhEmg3BeVkmXGyHdZUNnhIRppQ8D9uWq1zKl6TQDOlKBW7AYPLVh6HiuzWs2y
1oVehzj8+nIX//S1j5lT/YIUk1DzFvA7Eml1GNsP5JrMVPfF8f14cwkx8Q1IZMmP
ZucvyhWt4+CROlhSfJyWlRmsXpveeLWgp13rjNL9Ie+RG/c+UnlMzhFfn0f0vnS9
4FTU6ov8OhFfLfdyZLWeGquKdy8xHLflcTCPYHQhbl+tmmmCImTwYBP6ryfBUkKL
R8tQN9oRG5PJwk3BhGamBOdiiXChFQLE0DsBo9QIZqvyfG1Zis1KlJjA4b5aREVJ
cew9iuT120f5Sh49UAFjzYUqo/Ic28/bHd7JPDjc7EeFM61fjDhtQKZAQCWZb+Bh
PDgd/WotTrpxmGSaSZ4pXExXvctpoGFZdNkHwuy0LXJrYpf8tZxp5OClJEUK1/7N
XkEHDnw0YHx+Y8HDdBOYsLoKJnUIYIOp9J5NfyLUxAq88Tk27nYfTs0kRGWjXGMl
oRt/aQYSNjSmCQrdv/hprwFuc09dGBpWwqh4LiMa29ZD7Ustyr69HJFUnNlLdekZ
fL6CN6nEW3SV2qQv4qeVXxn3n1NgbPSQRBlsrgKcSNC27wN0PE0C+ilv7Tf8X9yA
TYBpZlY79BAgIqqzusOZveJO5i02qK1t07fzIkVv24SiFZTgEhLMr9C359Qzvpe/
SuTkjIJVTmI0Z7Tt0FFpgHkGKKekRvvcKp23jsxI03at17/32UPelO4bwW9weCV9
jorBEr/pdmQB2DTLE032SRHSCF2w2TaU+w0ADr3QBPFqsm81tTRwKU7WQE+jsJ18
mACpaTLRbfsZnOSpp0HTtmoqW8iISMsWe3MNnkpWr1lpPLN+Ks9RMuz1KiLgZDb3
/PPo41nUU34T/M4ahtVUJFGbCGvA8DYRDIcsq0kHzFsXbrKBka81NNH7btvHSRwW
I7ulNNn0JwxZ1KZpD38SMabsnwAi7vbELNup5g5SqIfmfpzn2mwUndWMWatHIa7a
ffzVOo2OQ2ivRl5qOM4I6w9G4dMKaF90Q/oLQZiYk9O9zFtiDZngC70L9REGF6jZ
glj3vrfjXWw3FT+AmBSluk2a6KaNwJ4z3e8qJwWeG1t71SiNiXEHCAImUifnddaJ
Sc6FVYgiaUAyqf9ezlCbej/Vg+sUInxTf2bTlIlK/gF7C3eCzbRvq3+2P5vnfUp/
qRT2wmBOCVAeoOJTM5I0SSB1VVaLLvOnF7YAFLZr3hxvhUYvXxMnfDKQUb4Vrl0t
NWz1n7izNq2NSA2GZiYnC679GVuHlrY+wLKh8E7FmJvnv5vxEboaeCZaU9t4QtjT
wj3ftWgjthkxPghR+627qTFpZdPMW55ElsXmzCFQ0tTChevBPiUwvE4QEvdDYsjF
RkdkLvgG65JxpyW26i2xhkvl1SNm7pJh3qdd7IuoRMxxjilJnhbGTxkV/BW4jijP
b5OHYoP8TStdMeghmhf9DJcB9+ixWcXVXDihSKp+Vn0P9Ubg0AWC7/ewLzLVI3oR
bXFN6fIjTY3IXBoeZkgfZOvmvITufPVQ+2xinomrgwh4FiMEh8B7ma5RpmqERsU6
8nMoJnvLNybfC330TIsh6wi2bob4ySXcYFk7NEqqPchGvbIwSGPHW899zaZu2mQ6
sRGZdkstfo+g2Cotxu9VzW1EbJgveItnCRb9Vj8y2I6dKsNFqAlADZZT9vBkFx2j
6VyWtKfWHzyJsvtPciFuBWzCeoyH6bPQjlOADcYUBToPcHFYe/AiBKx0D0f384OW
qMv4rFzgUQ5cNeN/cxdJfXMncL14LAlcdaG60P/Rcu1SuGZs7c5/5ECY096CkfE9
3v1oDRaqzYzXWWipoCw6K49dDDiKu/BhtHDEaMH6Dxofxdq4zN2E4o88C5K5ejTQ
m+SLkg0IQMG6wrcU/72/ECF5Z+Bp7Usl2Nw1857tUVRt64o28EU3ny+Ci/1awlCD
A135NWVopsefQw+SOJheA+GQ8crUWMZ60b7QMQI9RwbTZG35YAkfV/hC5B+UULXL
/lo/bscmVDs7wU5Ni2v3dmbGGuwZoZKvX7RptJtNw9kr5rPpUCRfUbsw1rbhCrP4
TNDO4HIdMtrS3qsM6vMyGWH1xqJg8xqPsSuCade4JO9nscfc2px2my0kEnt6Ovye
AATf5qHdNlTWYyhd9ak4uthqqX+FA9uTU7G9irlI0wEWps8kZbsnW8KK79VmYtqH
fr0J8AeRpbqwixVOHKkVBvg2btqoTZaTNO8hVuF2vp6e+LQnkJsF2ssV+ynA9i8n
I7+y/fMqA4XBV6pX804wygOYmnLLH+4A1jvm82LEbLLq1wHhRZ1h3VKgL1+Ufe/M
yyfhOpAnqDj9ULVYZZuMNxvL+KYC2cYCK0a3o3fTQl8LItbtRXASh1zVQxM8FVub
yJsL3aje+SOJ7AOWrvo8oPts1f+Fd85e+8K8Io/VvurPZDwHp19Z0366zwJGNYRF
OCSJO7BTTpb6z/u30VkvUuwz4stqZXtfSx3R6hqIf1HsHbZxfPxFcyEJY388cNhG
NqDm33x/Vvx36LazYcbVhuqFYwpVOehOZZpe/6Bc2DPdBYwJpoBwxBG4fV4tsWD+
P7LvdWJlG12Z9sE55CcGXggw022sAERDm+CWW8emrMJPYiC7IY0jYRD8KgBsqX0f
Mp2inMX/sh1/KmuZPvuEpPumKiw414QNfXqxDe6NXEBUKWLY8OoDlisbukCDtSlf
4VHEINySoCC9qZx9xn+hWd1oBJ5reWFoD1PJU2FfOw7/v1tbjrih7HM6Rg0aqSYV
oeNchx8cQuXtkW1oe5xR7yek8eaSuBr9oVXsP8GMk6vxeWi7W93Vp5t3prxZnnGV
9TP02kgPJloUdn+J3mWNRJ6Pw/OoXRo4PxrVFUF1BWGOE2BT4SM2LRrC4DZQvhqR
MXQ5WAR5JSXZcWlBo2O4M1Y/E6rAf4uY7yIpq7HHcWeIyAuHKkIhnKVyILrLawMz
CRHGxjeuYg9G7SUmWgur/CGr/LGGpEG+p2b7JypUBlsfnLIyZ3qfo0on3/lYcTzu
peEmgyd2bRZ9xKBUYBYP2vcbWJmpywR0IjGF5mtvbu1TUB1/N0S8t5XH9VPNqjwD
pTCveKcpqvgvjDnseZBu3u4OugDiBUN1Tz3F2yHRaMnH+plyHJvkc7kW/gcGjTd0
jADhsA6N/z36y0+HGOf5IGN2oIMxATRWrNYg2t+bUShLzEm9bdrrM98w97ce4U3Z
KMbIR8DdSZj9XPIVTA7fuktFHPh6yDVM1Uwo5UeU7hpXCTk0kkQUwtTacDTElU0z
RUHkIBAYbO+tF3LrffEEJFReYo971uLy3W7AomyZVl1oN3iwcFuMWJwIqGpeY7Lp
ZWw1AGojLvp2mfxKXezyH99hpOT/XvcYAy38/EjQ2t9pEHha/XC+YJBEVGFHQ1y9
ei1tj8a61GFQ4A6SilAMBfF69j2LfcU6HPa1PzXY7k2Ue30MMMbAKMMx3txqrTfM
q9oXXtROepyl2BC+fMyiWhh280SLQa6SnvEuoWEDnJDuWHDNfrfvQiKKmAoWAM9z
qA5BcrdCJ0NYkcwZcHZKr664Q4PZZ5jzl5xzsxWLwdVwwZIusEUQ7bNGejNLKgya
8HfJMgWulPhJACJrEsS4DN1HZq5IuDaiVUJH6L+xjYCHwfurBFpKjtHAtjIvEdLT
FEmQATjNQaprSKbEfFrAbzYpZTQFzM9tVrxnyj1+MlwVprASCtzaJz5WH74icMTa
ChZmN9Wc/+LnLc1U17rIUus2F47vPM7mtiwfsfGVEWXnj7Xnn5yLy8pOKVPEOigt
7x7B+Ibi+XNwwLzaLgDdUr/vh4caJ0kQ9dcIOfGazmF4AUUJjHyhrlOcPIOceiwD
3gkCu6sWlfaMCu1y2NK+AACHXwYqB5XjPDAi/cyZpl2ACQVjse+eRucD39IARE9V
QDWJ+JaohYd86C34DGeDX6GBYb3CQXoYuavqD45VOo/JhBeZz1f4A/hVzMDV8sEw
wD/sumAE0oZX8O67G/jQHkS9i3CrRmeaWqzbLbKBr8+sWDqlzTEMOHnV5YHIwQvh
RfS+EFsh8m9FU/GTr0V1XTHS+6BVHZ7jG5+U8HmotOCXv8e7WyYuxfkVRbD6RPmq
vcZj5UiK0KY33B8epaMXdm0pyuziBIeIl4Sq67gMDydkZcCHUOHxoAHnstYvPZNd
V7wvuQtUWC9oOBmn04CGWtT4p4hFLfrDtlvkmWzuaRQwbx8XhbOcSzYQ3Q7SCmut
GnAIz6VhTa/AklCNci0JWViesKHjG8qqln/pccZ60bsf9zm0D+imtYc+sXJWnjcY
h0m/8oOB1rqWDr7QJG7EsKtyDDbz+iPd5LAwoDwjINXzo1ljO+ncV9dwzfV52dz9
52UL/GMMO99+J4hygYYbO7LDwsbil1W+vMt/Do5WU1n54zYP8smUg2nYKcToulks
HnJmKnbmatauH6XG/2CRFU5mp06k3CyWsMDXUCDmPS7Uz7sDJCxEm/pYJ7aNgbUA
9dIi2drYHR53IrqRpPR1NxWdRJMMglXLneMngt+OE0qVPHFLe2GoWNUnZXQI4nNN
7OWFgP265DBoZC4RM8M91x6RTWeeVouCxWaT+nwgOMkKoD56FZmvH93oJnmEIbeM
sWElDoIZAweX3tWbC0yBcpV8VthIeiHwowaBVTG7LwYpiU3VbG3hUepN/Dw2j6l3
aDFUhOuu5QvjhnZeeCiA20L8zZ64YJ/WHkdPYeWaW99Ia4vM0WU3rL3aqcfU+fV9
FmeIrKk7fW5U82lgLVjBO3xzRaYnsLubJEfpTUfQtIgr1Jk5p3Fb5bipMXSim8As
F7S9kTfZzXSu83jv7cHqYP39d+FIyTrWEoiQ00bu7qT1UXBCT6KRkku6Tgkk8l6X
INBu7Pw/ORoZ2pjMoWXCWiclF+NmOxhLkX2x+rvvC+XVdDhJa9F2coFd8A8juhtA
rZWhNocDCS5jDeiUf+nb1MuBvM4hMk/MfDYkkv5Z7OMUveyLmEqxpY7r29SvQEOn
vz10nLEHT3M3kIyguEv5sr+QIBOIhzq64Hjxd1MXm/KWlyrk0MlrH0yizoJCHTHG
0VDYSHRXo/1VKNh0XIe5t5VdvEzllz7pU8y/pkZFve5flxLUw/o82BqYeGxPdhxi
Vp9J6MHEtfQS4igQQbjR47CIgth4rj8xIZh31iN7Pikp/VHvzGrlyoa2yxPuM8Pn
E/lR7Wi0/CBSVdzBzVEdHwSbts1jacxDrHI3Kv8SNzio21Ae95yKEc6ckZVjPwys
ZJ2eSUS0NeVpIBTniF1/vqr0Gq9hV2IGlt8O7jvUDysok+2YZiIAN0i72hcAnYnF
gvwx4OkSoCHnlHtuIsPq1JaRc0f/LPumQQFyyoAeYvqsN3xFpmAtm7HTYCzdfZ9t
/D0YkI8wcF3xuPWPqUkHDNpihKUMjLMmM5ChsJaZCqxybXSgGcO3I3MlhBUODz9g
mhbgcy/+wx9dWoNRhluYSEJvq88QDREcGHuKodSOBqOhZzbGoyvyn8Of9oWIXhdn
xotgonrelUkgkA2fsCvQQUj62/FuwwFMULnb0sHWoi/jgSAWU0NSA5jvKweVQUUF
+f5Ff1e2G4CzCfA0NE4BtvmFsSIQq8sW/imT6guYodW8uzbI3ArWLq2s+2OUF4rL
uyEaGcLPsFA51zRlHhBZNqtpjiSO051KB8p6tvSsBbIiVqldWqMurJRJ6WtWkvNk
rm/WkLJwSvJ8eJmjGzPs3vvPalrXu0JHnIcwLJM9uli7JJ8LqIlf47rbhE7TPJfj
1u9SAKxOVLkXSM+1k0724MJ4iSnkhSqXH2VfnzPmPOm12aRGZdyeCyagtTZhKs9V
ghX7rM2TpOYPxepYbu6G+DNo4PFjCashh2pybOzIsiBIrDsJyCDioleL+CrIFaru
A0tlK2NzgVw58hEQwumSpUnYsKwaim56ZWL4ppg5QCjOUIR28QwzhD/g8Lcc6Qmi
/5SaMmzw1TcVN2v8UPz58m30SAs2njdhtqVDQHdkkIeX1qtCWFrVE61/qXWNQPxp
N975mJAS/K1rIOQJPQd9fvBWQTOsHB6+8dFJMRHzkMj2brbIYCl5EwNWbbP7slVH
0RhzQti8On9wxcETFnzkLRO9k6crvZN0TtHbTC/ap96xSo9JSEaBFrSPCZJnN4EU
iRQ0kOMoY5J0nlAsv83d4n4OyALSeyHfn0o3ekmtlHiFC9/u1V1i/2M4IH5PCIrb
esT8A1DlskolwLlOtjECggz3YzJrD3wpC2aLFWM5Q9S7UwBasQFO4dj3yCNOEXgZ
nSZAqiQb1Gm+7Pb2gVI/wDcWxH3jMU5Q3lJ1In4oYK5CaXnXGCG7cqGMevD9uv7u
p82kR2FD+on0xFYixWiXOcFCoqD/1su1EIRq1i0k3pr7sVZUG1BjqYCAvK3ckMsL
Vfe1UOyYDrU7fDYNnf8uTDc1UV2DYc0DFyoRrGr3NNZGdsFp61cWyZLjFoF6L2t0
eorvdsRdSW15Kdc4NCySVvii77Tk8JqI2jRRQE7IBCF2ceXoMkjFP+t1srdcTG7i
CLbAW3duGtBsjHGZewWcOyNY06NIZG73MCzwGIub+vZwX9AjN5yJuxmkWUdYwsq9
nq/pLmrESVijuN6RdzHQzgP3EzGpDHJVYNN9XoATT5x+9icVw0p8tKJzYNAaRH60
v0PfTl6A4twbqUd4ebr7Tt6TM3BCJvQSverQEc1Khx6bkgvXbFAAvk/7NDDgzDyn
EoYA4uhDHXx9zE9DndoDKoMLDPUXhkHCi0e3gC62KPDlmM5iRi9ZYkYQnkfcuZAR
BJVAZGahMheXkgtN6AZataq67BTC0Kjs+z7wv8YRwklP72YIjgQoA1kmA0DsXiOI
7xfgnBJlG13sF+fzZOlzZURcm22a94awtF4KU6a+52Q4n76Ej0TVb5D/BczO7RQT
Ejue2wzlJXhu8AZPRlu4VCWntNBymNzuTlygluqnJOL9C8zFxG8z7y24a1tWLRZs
5awRt/vmy+bb0UMqr9eM7wBlNrsKsTDgUeEtAFpahAgpl1GIXEwpswMSBatJY8Og
BDxgOxQ1O88r9qb6NQl9LQg9QVxm0TeINiVPLUfJh9f1ssUFL1QzGKt2OTaRRYFc
YXVl8uXdraJElak7xzBtqpgeKQnkoPQ8tsJBL7wNfUpSatOn3VJUA8ZvRGmQl7DG
B3wMu3Z1efwBlSVfXxrQfX0n7e8pbL/zK/fufjTgmhQ8SiUV3Abcb4viTMTHRK4c
CEJbKwRLMWYu9I5VSOfTrckuLWnvaR2QIGTy37FiWOyzXydcQkueAeZTDlEwl5hi
UoleT9/3+o45Z27pmwoT2ZdEdHC1NDgjscCAVQI2D1Bz1B+oHGCu5ZpvS74P3qYl
G8in1uUE+WoRwl6lLQoe8D7h1WERK0KfvrgAUXUN2L+N72gsNFLa69ro2LjC/G9F
TQFGNECskGPZHHbjkjEeaICBAa24ruPOFg53/pTIYNK6gVsK6Buou9ppAOCD9YpJ
SCCoQYD7Prw/oeXPuRoorHVoVSv3ppjEm49H3NvIm8Y2UrK7dCTTYULs8j+j5q7k
Etu32b8h8uIt8k9CA/D9kKVfgFOpbLNGRzELZaIcy9+bxY0YZrpbPyLZq5mj2Z6r
j3jCD+FOZG+MQBoMRxYp+DyxM34sFW0NS8QjY3ns0NTAqli1QZU23LmI4nfiyqMU
s3UEd/LPrvmTNSXv2kGE5x/uhVLxMCN4LY9OIHzqU8MS7pVJX+yWGEXF8A1f610j
++KFSTSnQlY6/QrB6mzHsoCYcSFYd1pnRe0YCgFo+6ZKupzg67dKVlQ1kbM8wLjQ
IgnuC/1+zxan6SfNFI9QPs4oSH/IRaZhoidYTlx5e98oWXQX99QyZTjup5rCOifG
Y6CcYyTS1KhgHyCSjPHC1Dkq8fmbCstsC0y3asLUZkaskPGCctFtXtNFVXuAbAWe
2+nqlVJIh4LSnf87OmqbckpUK4SQ+/Cc0QscPSas4Y5VX3wGRGVL+vlTr1zxUPft
pBg2uPJrZ+d/XJ/XSu26EM9MQ0ajRICjEMdXWEXyNKmyvmcaQPNigdVGJfRI8JnJ
SPzHt62kBjbAShqzi+nKetvq2qPdhBWR+/sTmCWn6b6RGGevzeGI0oZ11ZiIplQk
WrmxCvNPFCm5NYPvKxw+WrIwaC28rNydprp5KdA5uTi0QzqIq/wX2mAGnQgVdLE8
kN8A1O8+Jk67pvVyvo4M3V492hkFWO5Rez2H2ME92xB79zsDd3K2Q+BRbYRP6idx
k3Q3s/4D8HspYMjmZmkJacGOL7bfPBrggJcRtq3/QJLrxf1jDh1uiL6kfcNE+fYi
+D0S4sAykoS5HUcOKMmMGpWp7aWPPDQDbva+SD9hx5WgHqg92bEiaWlg942z7JVz
FlAvvNSOBbFskdP9RpXqBjeQajp50jqPy/8doryaMATTdJBLlNe/9voYf9C23dU3
7ZcQg/4Qeh69GEtIMGI/arK57x927EWYwnsPVJs5Despr+d/3OPEp1cfOJCoXcEV
PltG8wWDr5Z89bDFAOrt3z7z1LOgwxN2kCYkbs+mYf07ofRQPJRtnXR5tYnClF5K
6T+XfM+Bvv32OdtPCEe8jhGLXu+PiOetF42ukvM5h5q+xJkp4lG7B4O4gMEbdyr+
N+qQFEAJBhG56jvcjY3IfIGylhGSnL2OZjC6vqRlMBVhG+oNcNPxMQuDKIluGmeV
fliafcsU1Ww6E2lU2opmaHGd3IEIPyvrb7gIpVWY8Z+p9ICQV4HAmr1sAcw2buys
G80V/j165q4ym0R/uxqdaL/CVGYDFjanVFHa0cadznuJWpCj6JRV6+4Xi3ZFGxWU
3Kb5C4gWalNCMbAL5a1UKOP3CvQ5orK7CqFgQlNftSAGKFSVO8uieQpsTG2wiDd4
XP8DsXdBGeejLAJ801GzqTEPjQ0R+gPelXJuIhNcgIZ3d2N/+Qo0Y6EkBTkR+ALd
li0GA4hseVcCKXv+0FQkDChbuzYaT61wIU/IstnFid7b6HmMs+g2V24yosoKpl7w
ep0ZWNBTOWWYmxfbw+1aKLfWnr/W8eDK73E0EXhidWufspxuzYsj/47tTLuTGLtQ
nbCU+JpUEjbLvyhDeBdXb+roBbDrlERFCkOi8/c75HAnyR+djcmdPE2zBH49rxQW
AsaJMVtv8JxDR482Tm8KQ4tSgdemtIx94JFqiC/XnA1bu4HDYY8OKyZXMU3lg5zo
031D8i3bhuw+b8VCexUVisDgGr5rQCzjFp/XatSgJkquQwWQLtktVwiLB4cJCu83
WVKfMjb5vsg9rNdnHjCpRA8l2yqF4LS0LKbxIK01a+FYH2WieJuDaRsf1n3uCFJc
0FREPv5R0UriYL/ioPrXV0FU8ZTcEegHEoFxyRn31NYXV93MscRLHbA1eKpJpw9p
Wc8w+y8mlm+sCVAgun7DNQ/FOVB+zDnUFvTKCgpSXNxpRNfjr4KWQ99segZ5WDzc
RJpVtYmyCe1P06OkLy8ZsMDjBvm07FdnsHHdAztg9EBPH4e+tJpIkZgCNSJ8PkQ2
F8752hHQBG1sTGeb+uQxz36b4iWZ1hSPoMtpzexlNqCP/RA6TbypKmBojfYJnOq4
LuCB+lEyECKPbLKNUHZjJ5nYcri8Cex7Dh0BtS32fdoziqqa4d9s/BOfGdU7HsC8
olTwbC+sjUn643JD+BgTB8mP39jXerAEseO4VRSp2uIAEyBdEqyzYdoX6+2xqrba
8fSTECv+mFObT0BuqD5/hDqRQ3I2UPxYmfCaFkB/dcsw3vmynQnT7exiIaOtRRm+
oXLcaAa6tMoEOGMlW2vgiqmxQ+AI8P9lLDEx/DjM7VQ/EB4DO84VRjub0cRMbdrd
uUtoWaZ7HMPvV7nWRfdMJRMNpedO9ldbh4/k1Ah+fjtAUkzTJeHgePlvpIlD7geA
+sLItqswloa3JS/+44vF424HaEA6nqCJxNsML4PTl8B/N0qRaDvCVEJ36xp7YQyi
0F/e7Qr/4OVZHtCcNIbPqfUdQwkTjqSd7Djwv1Ld+EbMNnip6nvOAQC99akIyqPi
38Ug83Y7tOX5SYrrAWfQw3llVn9ew9J9KRoZx8YTllDW/FRFeqWaa2/HMueExmOS
RIwXebWw54eM+lkFOlvydJ2S95H0I3QtMF0+A4ugKpylLhSyZhEmq+0gpSwpp/kp
W7J/qHIDU1OnkR2CMCadmXpVNAH7ZdXRJxFBS9RRJbilXowHrSV7t8WFTsh3AlfS
XfiPVs622HLj0AzObj5CyHADfPr4iXBoQxRucH/5Ps/ggyNVELwLuZdv5I6mUbsm
cjDd36Al52lZ2Kj3H2h0NQEaiYnctmSdNKOXf2G6izC9wPzD+fKRKXXLeIIPB1Xk
0mGpi7HrIWdeBp9u3fnG2KrNNWoT3jhHBd0nkezLGAcZUUUE8fAontL1xLkkrDxB
4Xl8U5jmIfANWa+MfWyd6nfd6I6lp545RefQmvx7SW7gb+//NM7ihgkwml/Pk+48
2Pi4nxNTWzRr9Ok08viGizdfIGe9d9MxWESyYDVzPv+NLYmd9VCJjSz6ZOSHPa9Y
NahM0JDfJAFbSMwJMqZfGBDo+xa0vu9vYhIdi9h/W/AV/AAD7fJs3iDwjuYMhtMq
rG7O/xSk2hgDR7rDAbf1Sm0qbfKVjELp9pFzv8HM1MWffG1RqPJ+pDANuf3N/ZKR
lBF/gztTnk628af13dgwRZa6fPqku3sQmNm8d/g/jlWMM9lZXwXDHnKo24WFjtMG
lrBy+CtzL9L3RsGcSh5+IueRb9QKOxaquxMwx0qvTDt38RmxIig88u2M+36kofkJ
GqpsQtIwHfMYN6K/AmEJc3WQAnd7a/Fm0A2SlfxYTl0J0JPKVTYT96sWR36kcQu7
CWPFENTsauJcd94ba/aOv5vAlL5Bo/Ae5pYQehceI6mi97iS2sCiCbdp/DFtzGYv
fcMmrVBNoSFW/ATHVM0jkf7+cXCtZgHIqrqxJuVlGbc0MBp/Sp4BolX8+Vh5YYGs
v1ZxnNrFZSf0AJElBox29sPvyixYRfNoubvoJ6suQwFynNTVhGo/Xr1MrhWT5tN6
oVGdUM5hj65mhiLatMytLx1iJXPswf1wJx3Hi1upXjQJq0FNcTpA2BJOmS1PwPFk
upGZ661Owq+522J+vLz4YQkD+vTGbM1YD2XaFniHtsscvs/P3AN7AFI3sloVCrjD
g31Tv3fJY+VMamJxzqaq0ljbOv2NRUTcupduGvFc6gbNXzRZE1UxMG/IS193OY5k
bg8CXVHE1CyslSslhSinsdESmepy7k+eKvk1fPOKUqBtkSQIU0S2EymNyXGrislf
XnSigY0nxTr/hwiY8HErLGKDAGGa8E+xudEJKNK/nR9nYzcjHc0Q5tu7aMDoV7Vw
o1H4Ke2aVbNMmXntK7TYzscuEMwKG//qNZtte8GVLNYHvzfQaccHtYw82mMFkMqq
r5yV/m7VRKuK4k9nLYSrDxw2lXoVQ9p4jR/MuCLgbZFrvC97uNXyfEVMZBua/DG+
0WrVJ7lislLozek3AEn91EIAAC/YmTvoYa9FweQRZSYlJI0EWODRmwtqVud6m0jt
OtAtFeQLSgPWxIwxPNxqvR6ec/eh3hligRZ4P3qPcd0D3FFyAUIeQDV+0pblfWUl
rgt6OkMB1FbmR83WF0hWEwa7WRHFAlXyxSVOPjc24yeyS5ZMGhToN7nIJqM2Q4fm
8KK+BGv9AWbNvkvY6pJhS9ZKt8yx/yhV2mjV5D45lIDlzbCAaStygKip3H4wuGc/
`pragma protect end_protected
