// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:26 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
T85KZRreUghiraLh1nWnj6cuvFwzN4woX0ODY68VvPYxhWMw9xgkOCdUtJI4/pX0
ttTF7UNK1JOVTctLzApQETmcRBCQpxv3ARrN0A+XXCoiNCqSFvE4wibICak3DBV9
2FRN2UiYlVzvcKdcGsLbccVsF3cYqA5e0BOl6XLTZgg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7344)
nYe9bJYvKUNdPVRPj3h3txaGDwDdtoqcN9vIFP5Q6agpsDrCXqeSoUQpFgrZeNh5
+H7RCvC6T/YSh9gFIh0Wja3rdZIroNbDIBhOldAkO7vK94AfqmGZDuy+tSac/lOO
8NF6Cn8RRaT7ZM7EiIjaVlN4Ga/ilOQZx50jqcbNvqliolXuRb8secXUEXvOc76r
CL2En6siwfPW91E9gz8Kf4loOCDSWRrv/kqfrpHUHLWKKoI4q0nNARwKogv4rLnX
l3li/tDv402hshL7w99vEA00JKhcsDRDL9tE88HspkggtSbGg6KLoPzxJ+bV4dnC
SXp1Y93xE9FvbVCxK4r0xfgaHBFiQDc0Ot1qPWAdvXOa+KWqaD4n8PxwJF1N+j8K
FGyUizjJNbx7lMeyT2Hn1nHFUxgU/iR3xxs4JWv59K2D38gfLetj2ns0V5k09Vpf
D4f1doESXQo1EuzdrLCVJHr9zS5jRfUGXExuUOG3MAGNs9E3sv5FWc4Z9bWqx3QQ
EO5gEmx8zbQ+tyWquoQxsOOPuFaUVZGOqBPRjLoybFiXQIGdK3qCJXpzqAkUBfpV
Vt/ZxBw3Wb60jLsF9MiH6wFKmBbYGPZZhrmrosbA20Q1iMUc5K5u2cGnqhDAuk//
Fq5c1w3TW/HkB9mljXrxTzKB6f6kN5FcouZaG9lwQ5DS9mYO0uH7QF7mZYtPDEWk
5OlqmTY6dIod/7ULeW9jm//v1b+nrmo1npvduZfNicMwZ6uzkLjrsJXEV3BmlSu2
VVIiIxyy5BnB3clzXPVhWx9Z8J+7+o+HRRY5l/hU1P2iaMgb1IZf/Rq837kRF9F+
YWlI6fKSvKaPPB3KicwHwpDbO00BjKArCZTHFGfjG2wwDc68OXl87xrP0duYkNfc
+5MyIJIiNofsEi2aU670in90k//MR0H7k1kPqcG10fh3A/q47vbYNgacAqMKhVD0
/+63n46RdN5tMyWYebaesViC5MGjoB1wNBPopk1KxkjB8KXt6c1K216XWburGG34
Sc1x1nk0aEcVcv/sromX8uuuokhLS9dWt7lPCPJcuCgs5zy3VMnTxP0HKWdBRb7o
wfXwbu6sDt0PKui5wqN2e4V4LgbfAOL8WSRJ45KjMS9vxBsuavZ73kUVnSUgBU6+
u7frEPoR2PaPB0ENRBlL9Z/8ZKNpg3qxftE+3gYB/PvVFJtxjqtDMqRtoZJQgM+t
jMXpcdnuYQFmG0jr6FUHbeIWQdUT4FlS2Eesuw04833pT44AxMCuTa5E7YVNAjeX
f4PXczUtJNW5HKVApPq0SYBwxL0qVq6TWgXNAc8u+a4yJwbhoVvt9NaE+7MD4fM/
+OwjnKk1Ug4U98DsSm9Xs18X2dSOBr1ozqa17/5c6sWaoCUGBLvIbm9PQDm7k+Ru
V85JcBG3m5pw6rGgNdDriZ3G2rofzt26kmCEplpWjONEanvcNrKslMpHh1Yn8sUF
ALk8GaRHU2/9Docquc9JYVMe12/oqSwRlOqswLJ4IZQ5205c+ofax9AtJ/mivuDI
lLY5+HwVrwQEUx//jNDUlKJvYWTG2DeGquISHTGT3P1Qn6d4xAj5M1qIDeZXr28R
u55CNT9c+sglScNVfUTlIvDW8bD0IrURO3zdM4d95xx2IqELACmxB6DjN/xzh43q
h0EvUmmdkmkZ1AtJJBftL/htlYEr7uCcCBneF22YDqo3Dxu0VZoGk/id80ADsqgL
qvJYcHRCX3bEknueCjOA1sVbe678GMXSZpJ7SxI85SxYoht1/OgSx3ByyB7A0d1V
G+V+GYl8ROawa8//mzIhxaciytWp301zcAApcFY2G7C/Gn1zYSl12dnEfg7+FppQ
e8EjUP06OHprv4eNVhtUrCBgawmcZYAvm+9p74I4UpiDGZos9IvDgyGPQc5McA3U
TlRlP/teO+d+FLxzKsSIUxjZtItuZwb+UXZ2qMlTer3qQOhjE4/aA7Z68UZfAA1/
CFYQOjwVHADqzmHGXOhe5kiVt2NAe3zp0sEjmyxsukS218u6K9vc0HmQUkf/Ffsj
s0VDB3ZPm1qEMRJB/vFlGinwDlNgfh0R1ZV7LbIIL0qNNXY4+nHQMB0OgS8vA1Ia
HkCM54OSLX1Z8uzBLZdSw9QnwnnEJmkfhEfZSS4tE6T0EsiiNe6BdudYEg3o3sDZ
PZ5+39Q4J2wNO8Q6w0garbaUx6RiLW69Pq+eV7uQ2bi//gbSRF+2fIfjvoQ+K5+o
tbzeVroNKBnmVJKZFzsy6ci7eV6Mt6z375MUTHy5pa/a/zHxEpZf2vRZRu2GbQF4
ikSFYt7LdDRy9g5LVxltfTQU1up+wXPPIqr3APIAZliqxMI60VjAYbHs4w4ocJW8
bLuQvMWR56i/FMFL3wLi/k1A2lQSA3ApQ4G7xPA0wQOopu7lXinZ62ChEhbAjI3o
UJG/VpGtqXxGdXFZR1CUOHJ8HNujedmP4SnOBcB9obWeHYY+xRBwUQuBKZFdRMj/
8toGw0LKfcuz0aVT573LUgkhjo3I3Gtsj4h5+XMkGnYUSGHlxRi8BnBsGWzZrMf4
PfhW60IIizwZmJZGxKpKc0E2IND+oxNGt1rUOTmbsIsed5ryViDZxHlZhZ29Iep4
rERvln0lNOEVow0MI+TzlbFlz8U9OMSfstiBI1e2hwJwJ2Q61TdsFOJWJrfkfoHx
p8vuvPelzU9bJvOaEKh8kmUJvd2NjWPlf/3GWXd5j+56qAjhupaL3qx4vCXxJOJt
OESgNGsO9rZC8tCa9QnWW3a/bZiGUE/ZSyi3D8SbV64x2mjuXPdhxRWIqYGf1A/E
jHwcR5Atho0jaH53yDLBVluEjeUprKe1ZB+bQXpaTtEVKUlgHr8t7LEbcw8Aw9db
b+FRPx5e2MRNzPyKoxvU9f3ZUO3w8I2kO8TWW6Zx/263HZo7QmNAifSXgF4QUi2m
/zb+XQSuV7qJkjFlyb1eWh2u69TfWZ6IKMgCbLbvhXqs2rUQPaDuELpxPNOxCzQJ
iQ9NUGwfvt5waSGpjInckn7U8wemsWxkcQr5vJ9MJsKLbj0CEypaPYy92QNh6DqH
K7CrnCHKDzCXf3vIwS71MQ/1+gWt5LbcAvepRbvX5FXzlCBjGnoa+mvE/AGKA2lp
FN/jjpSSEkA5UQL5eXbnLp+II10XkYg9zK5375DrNUudSlBGDMQhUPc/PeIgDTfL
+XAx8+IzFAdZPpGJIBqNV2n/zgEVkkb7vGlbFJRfc1tSpfBRjOsxLtAE4dzuYGkw
EDWEdfdCUGgfoBywyqLwWI2CJ23BeuOVNzaDYEQbcqf327KyyfOp7A6vNqR0iVjx
0t9shsFNnCsxn1Z64TzIboYi3Lo/hDI8zTpQP0c8yAaf8gOpDhYJoSKVw42rKTxF
dJXgfcrCemOnlNKxrEPLv77oxifefKN5jshbtpMUFDagxtS2pBrdxhgYykh/XvGx
khedSci3FF6Jw0xVBsHSWemPCNnVfIi6LXLZQMhX87v4toJjKmxoJiCwk6DOxaHf
A08kcvCIeyBB/kjIarYBms7fteN2Bsxt+4igE5WFY3Gt0P1FXAp2mqx8A+SDEePx
WJ+LnRws9AJo04XZkS4/f+e4G5JDA2305qe7plfFioZI4ExDxiIXlY14HToSHXEY
OFlIV8y61daW7QfBZ4c4lA3Sinmlg/DgpFvRS/ys/W2BXWu5K/ARtaCyeuTjQWSo
ujvhKL8+b/LtfLGEHA9+8+rTDQBJeJ10Y2lmJutq3JL37bHQ5zxh8eEqz+ctOgX2
4OAgnkmwLRXLAP0BENGUcjktp8X4DwTY8YV1TbVdJrk9+VeUrKnXpwjxYTkUSjxX
FgJTFWzF4MAiS/uAJWdHDbq5OFZyj75TmoHrGyNl5wcgS1FRLJ3oZBc4BcpeAwhm
MmiYPwMjbcTm13X12v6LQliMcFBCotuPWGkNnOVA4CZoervsyJp7Kl/SecWFnAME
5N8GH3AFvA94MJgU/XxU1xzssx832q9z/YpD81IWw0RWfwGFSfRmv6T27nF5Ahuc
uc1dZF6jmjiLpRMZeSuzkMUi5WYe4KvF67fpKSlXwc24saplZyeB/n0yoTCH8lLX
NLV2FGg6VmQ75yIALPZKWA4ERDaheGPz8NAgF7jW1v/s2ILXXS8zMjUeIBv1ZS1B
6xun995eWudYYruLN2YAyiwh1ADiUpoOQYt0KURnNG+1eUnUPpFJGPDhIt0WOHjz
2eVh4kDXwjhbVSnMLxQJM3Y2lrL4qyBsnMM5DQqavcuCnGKnpL08K6GMvMPcs2B7
eUgP9dzZDr+Uo1WWe5fWddRHZw6RD6Z9bxq/83p7ivMfPZT3YjWeAv4D2o0Na/pq
6RCCR521sGDa7nEZx+UFdZANHXhbe4J+fz8cIfsHidGQZ7/wJezKYnbqFRcDT3V8
bVnYk/eArNb+gsUwZ6ttk9nQWTfmBdLYbWQ2QHyLefEI7Ji6wMuJ7edEa4sPaym4
gXeBp3qTdgXlA4jbAaemUIJvhw25Kd+m06lK+3uIq1h4VnT8DA10iLmGrJbIMgKW
FGKW5Ea3fes5Kq0WapfFbZrOR1n0teedULbFjazNDsXgFWVweE1kQmax3uga4PU3
eYZ2Va6XueKkms7VeQPb9LEne7tffSN7n1HEUEEhV0K5iCQ4MdVoY7MW+ThRofZI
jTwVZycFxPDFevIDbOQ5CF0T6UFlX+YojFYx70cRrx2Q0nh9GMra4szKH+Y3oDGO
J8+15YtSpgOeAjfO7KC8kOM0KQuAtR0iRhKQlqS1+A63m8/kgkwt1vKy9JbWV/kn
qOPC35oZNLHxevDbHFnMNfhOomAxn/WdeAPutqTrYAL3FBl/hFxh/yqMBnSOUrao
uQAO7lmFujaRA5TxtNvnJM3OM6fuDMnaZQ79Igk4KEHxp1MKSEjj/8hRdjIn7CnZ
KebBZkpYtl4Cgzgb3aUO3opMERYq6EzhE0qEoupp9D38JyNhdvHSOC6E9JXVodQ3
cl4WUTwGkqGiOo9ohVtXCOW+H7ccXVad8ZmcICYQC/7VAvDNtF16BtS2OcbnfHH2
6djLeBRCX9KhTMIgVAsAFDJyLSbjNNW92T0D801tPINl8IGxI0btf6uwDLz6uCIE
aBeWjlBJzhKicszEg9xYPBf19kzjMlZhQz6YeKc8LEWRO+kJGHh4Srus9Fqonohn
zixLo9jmNpiNk61qyXXdxPR0VYnuowFKyoYj2lEqOC2WZMpyOrx4OhhNpwDJ6HbX
b6w1plQTUMeExVk4PGfNivPxvXOKVvK6M4gPZ8KbRKQtyCkZ6odvTa12wRfefrxI
vpYH32FFNBkXcAdXsZNDo7jhz6PhSQ7IgcXkpW9jtYEqIHOr5oCCsjh0dHjkK32q
LBgDm6TbmAVF0Rn8AmJQkznmmUbc0GXLeBXgOG9LeOFMxo5oYMoadfvmzDUh4Dda
Kuxt0/5as0zCWr3DwG3nn18LNB0RhCFba5DMwXMha2/hfT0YFLfy5+x52rn1QDDc
3ySqhR88NLHrH92FZrmgARHuJCJ7ZLsWs2esXJDsxz0ejnrVDQaTIoLx4TC6Hr+4
emn0RkM37PtgNytaXY0hNWJBPEpTE8GyxLy4WPuqHnQj5iQd4WVbollkvL542+5I
MSIip9a2vFtS+ZY10TRffwHL4/vOh20dbsiRLEqAqLza4389Dp5KZqStqCgBvft9
B1aPSjo8BnHkxfVBBPF6KoYuWCKA7cSphUL4uCA+vXLE/GFbb/QFQThamT8ncBNI
mGOvJGNshRFnxhe5T9ZmBTPnFM2+XvHY7WWIRAsQkZe6lK+qIcQu+MoBT1YjWWnm
gCFbt9lZhYedJFs8Z4XoiODqIxc+sVJkbW+QkBQMI6KJAisdaS+J+jhb3XWbnkkb
DeWDOzdfv+b7bsYrLtqCqwlNv2GOVwsh9Eke5xQB+ilCSC4nuMWTnD8AK77XrAmI
Uoa2T47wqs1/R20+rzRPIVEy8PL7cDPsnLkdLPnwxLJaV7L8i6N5WQryKSTem6mY
92IPIox0uk3rct3p2qvdHia7guykR22iQMFH05jB7xtS8Z5YPDP0kbiof6z/iMj1
tnOEgs5JN/C6l6ybbrXf2yASVOPBdOkSUSRRDWMlD9h/aW3iERDn3Gz9NWzOjjuq
LbB1zpLSAnmEKQxCDyggAhfQK5mV17NCivOD/4dlUo63tHIwk8/JhBe06MfUfv28
QAC1+yJf1Oy6YxoLUrTih2P/i0PefybHPZblECokDhn3ztvxld0EzY0Z27e188nG
KOQPCe7ln5E0KFTCT3FsTGpK/swamLvSz52ZJZzpqm5GuuUgw0Ie01jPOjUiCNPF
tKvjlaOB6HAfN82rAL0Hr5srxtV0Ihf1/M7a4ku+p9oWjoxjD2bibeTf3qSvIxBv
UxfberUf7DFvELOXN10Lr8XIhmoBMQbXEzOO8MfCv2Kk1acO54CfhnvBUJnmzKZ3
1C1LYh8iUh/jR+aYsxyw9CsCVQb9MRiTVgRJAEJzvX9dET2PFP9zvBAfeYYQ0Pi4
cr//Yc/373ZG86JVZIa0tkArdQreuEuPEh9swYNYpCMR7yQ/N40uJf0Bvu3HBBlA
CHZhUsAAvHBwQQseuA++JywRKRCRUS9f4JgQRGrOYTWLOjXmjYuDdR90Ml89xUwg
4+71DkzJh71YJ5ujhaYm7U511wXBNBPE8vXK4RJhKwysx7LPURBHayLVO/qYM5ru
8r0GEe1PuZxqr16O/HUJXoR1JBFMY4Z2yROye26P+Zjq3kJ3hJT51AHECeTTNEwn
FeahwtoCGxx8Kub1E0grpF+usJZmYeGBf9XKGJfpAy1xwcKAbbKvh0Jft+pD0ln8
eFYPaaxi9aZwR+2slinVH+/jpCGJuzW8ZPPBJ1NDIS35mnUbG3/8sBkE9jQVjBMN
VJdQLEJIzk1oyZ6HAPKAbq/oTFQK7L/4sz2mAhVzh1fHBaeRDnS54FBVmViupZJt
iAHtWT3Mg8VJqtCSdm6ViaSr8gD8Y02XZXNtAg/nKebO/OW4trssbTTh4LVLg4Hg
eMlWStc8yYl2IS1FkAUrffQ6PEVft841MkpROSBmgcKXCqUE3wRX3m3KTqe7/dJN
IKpGFhkPpxw3fL3psPURKnQiW2SEn2QGxTeBjcHcF54PdMgmCqXc5/U2g8htMpuO
fr435gA4ERAGlDjpXUh4hBLueP23OrNB5otR0AfseCIZEUXGGhM+8hABPvz+VAJG
jLmuIjTmDp9i/oEUNJPyxSqNU5bO2Q5Bt1vjnN926ww6ZfcpknD5KK++qC58zMAK
v8XaFJ69eisiOTNiGLbrBYIYuiIYRPc8s9l4IHEOHuNdbZLH5PoNbvvfKNvodO9r
YB1E1KJkQjziskqry+pk2Y102uYZV174Y3rXuwNJP08bf+7bawcimczp5Os67VCR
l0t6x3Frienflzx6mhoVS5qm06MRmBpgvuclQCWu/hdPNQM+kfTVELL7t78/9R7i
8lX/tJHRdt4UmGA5Z//+IWx7wfHBF58giz3I7GRkZpGnEwKIRyFj78kXcOVXH+2E
fwoTZgYxHe1Qtg8Xhdxj34AJltvfnRq+j5QIgYu9e+HbA88ZJAGIeynpEk4e8xSd
sqz+7Ocm9uFHpoKBClT32jzIfZyow2g5ivF5/tGnuOH6xb4moWsS/Yu3gQJ9kd6k
LRD3z9e1uSk00ZDZzXjEmn4Ptb7FcuJ4bsyJkwO9zn6wdmA2m5Eo82DJn4VgBp2O
w6MemApnNoH1hsu7kzvTpgnmagwI7x2jzZ2amnLXYDwZZ3nEoN6xKMzaYBZyWF9T
wO4MMn3Mynz8TFzlvu0k6TYkZhlNldxADrQxaYQSnT51SRYcrlYOOBu1C3+PlP1y
zcWDRsjbMGDH0t5RJ+ZAI0x1DhfMj5HBWx7tan3iGO/Q+YiIKnynX64nGye9N/BU
8p2qnr2YNfij6x+Cb9+MHh/kysbYF0RAQ38vZXF6FxjQ5tN1vixmrQP3oWKmIp0i
QSu4qkYfpna3KT4awrKVedtOowrIQFcujbLWnkd0LMANstQIsqqo1/l2EhKg8c+U
OZWLsQ/g+awVjneJ9iDWV14/OOsWgdZUH3iPqnr2hX6hr9v8VeADvrdL3g5pgexk
sxn5jBfhbuFQvEjnvl20O7FxbdyZCAbUbU7KaZXWG2v433fyxKGZpx36DvsWd8LS
MWWbrV10A98rlEl/r9q54sBwLXowHnCR6PCAIztL8DtTs1yDia9VFdWOf9ff7NfS
zlN3EJMH91ZKdM3U45w9TvtwUjG0LRgHQJSMfkDozfVsZM1qMQ+ftIv3G+WvCFQm
TOl4lsfV1cIlzJ1ydbX36RDvF+aL6fWFPlld0SCi8M8HEeUchpGJ6vYZUFiPgzne
bvkPH91otKhjtea1eXdNYqhIhhnKuXTpFI1SOvTmf65Rl/5MOiTHxEQOpfMbP++N
cXL32dbulqOO/e6GiHaQq7zxuWhHKEI6FR/euTh6ZHYZ5Zo4oPy5uKrNc1zQTZ12
lT1x+Mz8aaxeZQKQsSosvEew1/crR1RayiVxMFgoBV1VHKi1T1eks64EraL3EuJ8
tulg4ndaPas6cfcsi1NpXV7IHKz78AuJ5vf4l3mRii4xh3cFw+HOwmL7rDDo8gs7
UoWsqEJvulls1JA7gdX2eZeYzF0e9kU/KeBCVvEX2ecAlWHSo/ABYDuITVaGkyHi
IC9nGY9+QuravQkRJHJU2/KZJ5vtY7vCGH94FE3ThI8vCLDXbb5ceXxrL7LFF+5e
HOLTy/rn1O9+KmxJYam4Q4SjrbHO07jxVeK05YPSAlRaI9CwRbVFO7WluK6bnu03
KIwZHBS/MFGS+EUKw0BXrPBsw3cvIg/5mc+9OfyiY/8QJzKWwa+CnTe7fY/6uNxf
c3DzcGzIu8WcDmG2gN8ZrrCfAJjKc5/UcOeth25YrvHntgKso3xFmXeub8p+hDK7
YFUwcobyHxAYC4f3UdSDffQuUihPdMZvCcvoQUGlks6gMAktevx143Nn4MXiAjRh
6l/Vws9gzohNY2P8Mosk48cUTtczGfEyT6Ja8Y7WXfO0YKmZ71bysBaMLMDaK1SU
gtkAHwYZburxZMmCs0j0xztQLiCDO+NEHHH3MDNw8bOlMzabWb/+2VrS4VlDlcta
FdqArJFg6meeu1qNGxuZ6MaXzi4cbWtdBgA1aM6vEhCSygylteng/pbBSc15B6TM
TMjzlap4ZgaAWHjaqBFZ+wgsUi+qoe2/dIGnoexfaZFz38fE3ikuw3wC3NWUo9aR
jlrHm1wVBlV6eYUWYQcrx3aqjWTiKDkbW5MpfTBeAYUsTr5WcyfxSOZ4XxOA1Ukm
xLt4DvHU5Xp61seQMKHH6+6U1BtT1xzMFqkSLphOOu1+k2CJlfObm2lwFqVFttFj
wlaSbKXjzMU1vTjarMOf/HRmdGtmSXHmN3crcqGcgibtZCf9YN0EWb1PH5sO2ire
YU4/NwydjHTjdX4lcsK95EqlnJDaB4IfVDbp+MMCiUKjXXDAPvqAuJ36qOup9SwM
OxSBBenYpo0H4SpxFDYK6g7meN0DeM0bXBWlU+Qp+y5hpbBFGvoQP/HNGySP83tl
yzuuilvwJ9B3+chw4TGzRziRPI8CHhvnbnCOba5biLyzHj99WgOTkwRIZgu1B6iB
e5eT4ow7SYoxjEZEc18tMQL9EazyzsdjF5J+tU+wFQgY1AfqoAC0nVZAkKKVsAkU
m3MC9ae5N/b3J0HXkK6wpoAeyPZtSW8jJJPivVkOHsPwPGZlH5x+Ok8sZwwYy003
`pragma protect end_protected
