// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Tsco+cMMgsCOLmtcKYOWEX9RM2do/SZDWmt6r5XcBfmbchVrw/V11SOOr5AV7wXv7BIqozQaTo4u
3FpL5A6PdDYEbVm77OPO1Ztu9DeNK+DGM6Axpz3C6PMVu/3IDl1lQBlbxYqSEnHr+wnTd86KZJGb
lJElh0ME2cQnZ9wCoLeUlsZdUEo5QclT30zU1X3dmeo38ojAEa2nA+YcHzyHc78TIEqefeCPR/Uv
y7UJYWOPVt7v1PRMiIOW7iKT+/fGHTXNvhQxWLTLTzmEZsoyVpa4i8lhmgy2PImF62FV7A5skLzv
okwvvy/zG7w+Lv9PaxlMUw4wZLlmYI7mNJttIA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
arT8ou8jprAftLscjbx99bVL6+uCbR702ZnShVC9mh8l9mIt/jXgApRKUL5gxda7d//K40Fr/nWr
fcmlYpuyR7tFKlPa8W5nGroR/TUOBCRv/LaCcBa82JtJfGeS3MyUYfTQmE19CRNa5hXZ54yGMpv7
RL1bxfJAEXyeRe78biUtyoP6/MduDLcDMarAIoNH8GGLKkFqiBlRwQfFLMVIhgiZEU3ilgVH07X4
oP9u6UaVckpiNmjoPFwzhFD+ShM3Oewe37+1IFp8+G2tn4/XlXKihLcqYUhB31bQP5Wp+jt9D2J/
3U3L32/6/J9ZyCjcYkdN27OEb0zOtVK7tbzVppp0bLDBHcH0MZPdZL0zAqptedxdUGFzlrI8a6gN
UjNkaRhJvJTVLDe8fuZ/hnJHv7rs4WSGvgftnmUXyq/Fa+hUMbGtW9Ayb0I5gtI3/qryHlSkNwdR
7RRNZmxT5kO5JsMDwMjCw1e1i8V2ZgPbz2K2DWainoFLj+yNBz99fQN3JOMAlBlF0lZXsjyAFJ2g
nzqp84am10JvG3krYTjFA7ej/qw9uyklPYXHgZRf2CbAJjLckituhC5z8pyw5dOzELwDTnyYihtg
u4IjTfr/oS0uIR9CM5RqEdMap8fAI7uOf778HQD1zAwFs3uwtCEx3FOOLWpB2Lt5wU/rCSeqZ/O8
Oya68D994ToAVz+RpWRSjUMSDIrqXgNLi5MBwVH9STFv2gUu0fdMzyv13Vb0fTwqhHOgsBbwHR71
yHN57eOc8PFWTnOEpVQ+HVBUeWKnePgsCaKeAsjo7ckzCiCqaBcwT+4mzMfK629193GWW/jOCD/8
FUdnY7P6idKa0RJ7UbkTbxPOa6z41GPu7A33P4OrGJW4+zdAXA6Pucu43NxoMRjnSHLoEf5iaRq4
G+xMBYUgamhHYPe3a4HGI5YlOKF1haLKvLY7xjFf2POHqw5gojdqMbQKOkZ8CuaTmtOhNWELHcAn
atnvpFbKMRGGhnG7JLq1ZXQ21hIbtFEUG4FTYuKbsZDgX7P8m32sYGpUJxlh/oJOGYGmKGG1zb1q
Se1/XVCq1oSXJGo8gWiZXpOU+GAa/qOF7ftUUv5WgQuGtjuihsc9a4gZ0dSTKo8pCLrcpLqOUF9+
4gtFC9GjHNMRTsc6SqkLnw0yAWGGnYujcFU0uJjk9LfAsRGLrRZm1hYE4SNnHxENm5ytKRvtFZSM
sph8B8G9AsL1msO41Ve2/5ERLfw9WOgDbMIYMN1zQzb9EMewejIWxdjODY4sG5y3hEsXgc4Uw/EL
DGfRgHIlvK/F5yWE5FCtrKpjUK1PB5/dW8BRsZxnbBCO1XsumTyXmbdlN4lwa8ZTniUyHfk5mMIz
w1wfMx76p6m5OY5msDyW1l+API3rP5FTigfPqUg8TjiWtQ7Vg81vrJPIz/UuChabo/ma4pkNfrA/
bisPz3vi9XUWBpqBzuJQvtpOSxJgUMBRV5AL5obp2TFHtEJgrqLAu8vsuWh60sXGejcAWaHxy9fi
K/O/5Md46S1s0nkRJxXVxj8eh8QGcmLrZUrKrtFI6AWL/YVpFrB4jFk+KvGn5ahZIeAgeiWUjEEY
NCX5uXDr9qp3hvTXJfWslYHR4guPntV23BNoDDeyHlIkC5Sgzrnx1Tso+UfwZQ32ovjcUXfRsyd0
fdYpOzTwlvch0ImsxP3yQ0OmVmydhxdVhRwfvOCFqT5uXH+75Ig3Ag0TIPm1O4IfqdSQ3eY9vcV+
N97HhiK5R1rgGhOCGFAasHzwkaWj30wASFRZfROsrNoEcNaHEIJQ5AOAr1B98FTlKDSbzIQF/VZc
t0GfOrUGjG91hdxYq3jT4zBi9nnb90WK9VMN2CF2UyrFiSCgSy1vOJlk3c3g+YDZz3XocAdmGP0W
P62ETLGOUdZ//NKaDgddhNWWMLe5mmtXRMraWnP/RJQUz+zqBX+lgpK6CNaJpTmS3V3tD0I+x/LI
WDbuQUFKLpcCjO75I07mIDXMrIMPWcomXlB7zAzuFw/FWhDRAMxGFyARpF6/ByuHRQb/F4R5cHsE
hsVzpkC8NUWjZfHleqrQFAfA9LQ/4PiizNuPQSxmrzoavLjW0KcyFR1VmJHaDC2ICnrYskGZ7S7w
pWmzURmXl1ymBDWBqDy5AGu8ZA8vbge5iOcAh6y20GvQZXQHuMdX7fsnU/u4T/pTSZfdT7lUpqVl
ZYhsLaRf3ZPlXR/DGNKjypLJ8MFAfFy1oIlgL7fmKpJSRSTXToKv2tRCExlpbWZmddRDzSBEUm+c
8Y5EQvyDOMadilP32IAHNMViZp7dYKyvEseC8Vs3X2rzh6Sr1duYHg42bhkopnJ/XHYM013Dy9Gf
wEmG3HshPk8IF7TiSPDXv+cIEfB6eMKCNS2Xz26/CDxmUwA2si6mD/j6VxroNksrEAX8SZT3XS3O
+AHgyebtOtYU3JE3qxXSvarvx9k4Icvjmeo55buGOFmG2AQXinoXj6zXm8qIjQP5FQ7gLHqt/KpE
zFVI7izkQr9iOAI0jw7a+leF9I5V8j53+JV+JU+FIhQlVWETYcFczZjNSc98DqgMMjtqEwRaRoOY
i07S7QLRHZ/4Cjr03lRZLDmEPfeCqeScvrcjLtvQRjSqsStKSzDyKF/MY5oeK9h+iUZ65tsbYnPF
Llx7ytTsKArLDDK99FQWOVkHX79edqVgB+xFKYrX9gPYCQUe3A3+aMekcbSH/lHXcZHZ49UwYF2X
/dgZM+Nnl3A0DpxT2BA4npOLgFsSv2t4HcUlUZ8Wthh9JyzgB76dfCoj3IJf642Mjhur1GGtC6YX
94tbYrkNWmxTU5MIUvnPTha8bLza4RMiXjK9dq0KualMwNgstOXiqvkPhHOIivBAGPpdW3ybYQq8
3gHoq3lHsaKa9U5tP4VYQ/0LM7wCPN5kezGqQ1bhAKhBhiwG9WTsQHWpRzA81T7F/GjH5+3xS6jk
6GJoCzYvkbFwCbVaQbLaVb5k3KxRgmT9TE1LmCON75GhicHjLzpBUcBVbg8ACrtfQ8sbiW7BxiRB
bc0pjMKaM5Z47OzY3wXb1xhmoNSrvucjbpascBTYNKGHAMN5XR2Ie5rYESDnIPzuQZ5uAOWL/Zr3
l+K7V3+QiEgfeNpvMKplABAQax1IZNvLp6Lve6f8w6oYxoH2DWhqyPrNktLxCAn0K+EwoYRMFUZT
8lYwGDBX3Sdt3omW9ffaUIXr2YmX1q/pQYy6H3ELnNKZaxe12gOM8nt5MVOZ8Sr0FEiaL9wcUr+A
wkFq/Udfo1JbTigM/CVzBTCfeUKpPtHe9E1+m7SNF57/LFqKd2EzfIeKDBSa035yV2ybZLeBhOrL
VMkJwzoPSAYoJ4Nfh3/YvotrBADfkiQ/q9UZVHbaaOp0TlJyrcRUmtMuwZIMj3YbwluHS1NSvO0d
O9Yu5GamUF71klOtSnJtFUIGlFR9WIXcg2IunlhxshMZX8MFiay8V6wMqA==
`pragma protect end_protected
