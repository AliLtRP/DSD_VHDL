// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
U5aB2xYDInyceSGu/IBRS1GnrKgA+hBkNjItpz52m7uJh7T3HN/0eY6R8aO4LExgSDPSskEE4kk8
i/IafCFcrehJVU+6Sn1R9XGIwHAb3sOM2AIux+OO6uuAjWNW/EShmYIRVl9L3t86SN/YE2ah8pKX
M33dT77IFsOrBkVTNG90glOWyZRtebz6t3+jiSUi2bspfWR5lvROW7Byb2g3UQC7wepA8dIqZ86C
0CP2OZZLIdnqlDct0GJnXMzEir/K+eUz3zzjw8wqemJkq5mJxVBLJjpyMEOgwsDrm2VsC5XSPWyU
3N4ntOrR1c9A7ScWcBWdVMs8bAxfp5aBJI+8qg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
tayc9kAxxgXSCuBC0ryNu7Sz61YJ3OtYPxtVHSMqND7Q3OAnKllXcZSoeEhm6nFnwspREqGQJxL1
LXloq2gvL/f/Oq9WUcOuRtPR2xfc12aHBZo7zC3HgbAzfHIlRohG/PgJ8eEUUyssbzz76JYbNDMK
NWhcLsXDQuDxqyM7Qha7g2TVjZsheTnE9yYrPz1kwHrpkuD2zSQJxuG5JtX7tZn/t5wER5yTehQ3
Iv+HfuWVkkbYpRtFLG5A0DQErA2TSxsxaREiZLXhpKqH5Tc6U1GVLqJKfnS63Y3buh6a3BZqV7PA
5uUY9j5L6WlRdFTUlSlvEjjyqNYsa3pRMpQbApWcLAuqKInSeVJvKr04Zw1RGXIfmNrYY70hnT1U
sIrWPHdSdFVzmVvvpM9rzL2Sdc2rl7d9VHBQ9DyVic2dDNBcH5uF4XwNmKIMVjWfqx1rV/BmEYdY
u9Ixm6fMqXCdIRh8l3rQgJ1nvO4HZnUJ7FD5fUQGCuWGN0hP6ayhPUu3JccrumAQwO+VQTlVrdrX
GdUK6/uSpEJ9ZRJ45vXs6hOMxq6k1Z1gHFObGzMoTXO9+uGPEuvBdK4MJaUqPvaBwBzzPGDgj5Gc
1ciGXAI1TtZHdLxtWYYm8v93aCVHf17yIIl00NGtu8beoa8jlQHx4wKAW42dFpE9qCVtq3nzxFiX
LfEaZaQCCNJaa4T/s4n1GwweWQiJUrkPZlP4C7dRtx+Lq0tsp+c6WdOcUSLzgv+F9h/fNRlhV4x+
25BRI988rgrzK8kZGKd9Pbuij55+gwQwflYOf5sWjpJPR8cu8//SH3egDb/8KoLzwSUDfxOA6+HB
gfGMmLgLojvKtVuOfsG1FIE5G3EmJySLfmIHdqpffp2IfL4tvXBFQm4I5AU1wAwniWMMHj7OROKr
IG6yjVuh+uwDEVD14elC75NCiDbnsfz+zpiRCNScBs0zVx4631qxjwhFj6d6AQRJckUqRaOqAihP
vXTPMswNUMa5h7caPOSiUojUtigScJ/j1BLx3i0xNsSSwrSPOh+5wnuoY9Y0leWHTUz4kcksSSQi
dAVBD7rrbf9pEJj5noQBZM7O7glDkYPRuykn1veoc+NJgaxLDqRiB5LAONY1UTJEzdcbm2CpvdLE
ERr7933yUK8gSjuifl5mzM6Q8PQp8GVSTiSr9rnfur/xRl+RbuL0NjjkQ8HPV2Pt0XMBLTkxj2Yp
qj8nt7KKNuZB1a2B3RWmHuzIycCucqddqtloIEn2On+NQWYnDnpfeLNpgJtCgBADaVQrskHW0y/E
RhZ25xbmnQycz0KSGNa7YCfGQUOBrHbsswX/ezyW0uAaytr3ONOuNgohnQyqa2qr7R5yi7lK0Q4/
c0xf3GXOF5SONTJZ6InbWhT+Dgpv9qIfYfRXLwDrduvEH+WI9myKuovAJ+zLBlSDjaNXrQ5bKrI5
He310EyzLFWh7Il2oSIJ+jvJg6FrERbcXTZqfQTe0LnqgFJ6cZq119a5P8hpGNbWGib+ssqM9FC6
QPE65PZV5jnEPCedwzydLi+TZDsA+8Am8w8I1+oPasiQ6Af2eL8QzqoL9C0YDWMBkxfudNqb2koF
VgcS/StT3DPEaVU/wh/sFyiPdk6USu8bkjRuPTzDF1ttGKnMDfeY0GMhkxO/J9J0nz7yREx2Lppd
xds4pI6tgGns5ffhHwK8usXc6yjHXkYSifiEmNjDaybe9wnVL9E/cHG6MqgenIMNNx0I1urLSUHY
40L+QhzNnltIHaJmdx3ADYSmZ+SZb4n9VLt51LkL27CIdI73aO6U0if7Sj/HQrJFzqBFVDlrGUa3
rnCaFMOulXWE7BzTgxanAu0uubXxPSxe0YX8v4DwGF/rPHPSwYwxpne+3X0moA+WewB44jE3C/zC
gJUuLwU/FE8zquRgib/FvC6nNzOALVsIoHNTvYldFYJ3uGIXU5eiEsB3fyNnFN26EeIFJnLQ8WS7
h4b3UnMe0HqDf3VMX9jbpsZKMRKocuXLKTGSwtKZfuwvQhKljXktUTagLhV+G9bcsDF/aXqRHifO
2hNShG1P1q7j88Myy83rMBkAO87Yk9XwYElb9OrDdTYXIUPNNx5acR5XmutTlghDXVU0fTx8gXtL
fO9m9JA6Rir5AtOyimEHBRJ/+sfIHRPcmZGPaRvFBh0TA3rSjkMxvsxwd3srPsItZZoc7Mpa20lq
ZiPLpvHr4WdK14R8qcj0hGh0dutbLswdBad7Zn+oAs62jFVO2/WWEIkEpc2SmJuZ7y20p50nPypN
dFI604QWpGHhQ0t9OI87ixiEZNYgd3KyRiOpzmFENhsOFw68cDhvlaD34WUtY2anZtYSMQYfMdej
c4k+csHv8P4hef54x3w2NNCAQqWRpoB0BaWHHyLxLeAWYZlN3A16K5vLiup5l1lSA1Xj3dGh33/B
2X9L9epri/viLUJWzbc9ku+4LVd7t3BdgqjFiAzwIs+dnjXCK5dYouTWoZjm2f003qX+TbDAfdJP
MXqm3SusLl3RpfZcfpFvqOHylvyX4mJqRvv+HZB5La0UYB5YfaU49VH6gzCrSMn8RO2UfyE14Xaw
NfKGgOEyDO4nH4eFsEcVbz/h+bQKD46sYZkXJwoWR6hnnxyql+Zx5NQQnalkeEIwr+BQsyDUWaNu
oSF3x7xxo0LqbSGRzLyo0fcfY/SD/7Ehuuprx9gEL0AWqSZajO3i01UcKa1AKAafEpksv1zFKAAA
8n0y2OeZfARl/vEeXI+QK8q5N/QWM3h1GYTEYuv9YwnWx87m1+MroCIgO1Z8omYIjA5MMv7E9kB1
JRsYJJU3McEOEnpppSWnels1QlsYWAa1F/XTL2yTk7tbkPepgRFpdXz+2+j3dnV5DkwjIEtnGnfh
Y3/fTzePmS4PEd5b0OqugMJTv3sSFUz927DoIESjbseGlUoCppz4rLRy5O/84GqYEx9ckgORGk2D
UwK+/xaRlb/Av4LDcEpUOsQb0wlmv/hwPT9jZOB7RKbYQ9gCweZa08v5QCfZJ1VbjwFBKm3rC+JO
Bmt/swPDFwINEAYnpbIUHqjH3gu8eghZiUPu2f0b8tmsCCgJOMPiMhuW7+hcnBxRAVFuyPp5JICQ
IhkpA8CFIj1jX8utIV9c6B+iv2nTdkv/ZegFkBezbcRSZKX3d9qxSikzAbnVEq+ID+pIj7//TNFH
M6fEsW6ZyPZYrD5RhHpkFWhANITOC50RUSFB+Ae1FgON8jDKiNH8JMLJZJTv4yClXG4Oi4CUxqHN
vDlRsmI80URz+4o9532rmeAjT3q0xTkkDL6Z7rxJBNxWw3FGTfT98hxguC+GvQlUKhHB+l+YzyBE
ef8xpFSIhm9cSpR3XDE5pwELF0GgPDtFeEOY3J8adMuMG0G/lheGvcbP8xK+mp+TF3iLkGNcLsGV
ofrKYY1Ay0H2kpjGfN4sdEJ1vagg3B6Qs7V7jqbsc+gLjhK9LH+scBvWfIPG114iGBML1JoZ9CIB
hj8ftAgQrKmc1X/t594NNkd5weYwOgwNSkFN3VSkckoiNOQdqdyLedBT/v9YjEsOTNfW1PvJKt4F
hMjWEA6HOHt9uTA2PdMQw/AUhKgb2hX3FORf/Nsc67Y+cmIluTlL2otViMplHOK0aP8Xilw3tmc6
XCid1BaeSw8LfsJZz5Rpg3J967ODXdU8vqjKpBDdoSl+RnXgizJfmb/XTWCZg9D2vmwaMrSkFkGu
Zi2FlRUMhEB6TRF3LtDHqaD7YnYoU6MBemKKk6wV9HS+ph3mdda5Hg6NSZPJtkB19MSZBBzL5pnA
iq+uewA/wk4XMnNcjWGkmhSK+mc766bHkEYDmF/sLP1Z6KDPjHFjLSbi6jDvqwEF3B3EqFl7enfM
xOPj3zy5xSG/jZraRDqh9xCE45MwZT+2TKhl6IaKX29Bl4SvYSrGvVE4/ZZ/T8RBTR7A2y+Ej1C3
UNe3h3AfKzPLaEmMP6Rljei0Qx25R8Q6yz73+lwLQAR8K1slyzsolWYDrtztsnDHyxuNagAm67e9
nikS+vQq4Wi6tcL1ijT6TIqKLTiJNdM1IVjuul61crVt655SXaoyDNuiWNDw/pyTuCzfH6wSB8dF
6ZbAXPIlo8X0KuKfJsYIiDSemZ7NwhUv2UsPxEvlnLSIf1PAzlcARmWHPHH++1D9wMjgkLYI8VN0
mGUkFlLwZg0h0WlHraWfsgz42rz0T3siyi2MGpcI+IQ6utOWZYoPF//xIYyMnHeGT5WulONdfUxe
IRv5EgxxkJUxO1PVTidWwFC+2NZ7pfuk3a222jmSlCMXAzvzni3whcUPitlf+cK3wwUGardOfQ0t
mlf6tfqEl6BSQA5+f7Ur2e16qTFvMmH6OX3QyfPd6hEsTQ7ouynk6txsWsyJO6wc/tE430Z9o2f+
z2f/f6YhbETjwuju8ZjiYZd8ANiatLCCq/Wuz4aiUMb9Do4kMn7SBaPQdV3TNvLuL3FTlkfBQOwi
+aLJTRuC30AJM7Dr40JzIgSSuLv+a91FwQCJMtaYP/PvUQ+DEbaIgrkgyeKa4PG1Tc9o8ptdKyYU
9EkOC9XGC6YosA2vX4gHQhg+0bNiiDe39jNmlqspRSfzZHExkYJyK0xBdyp+FPq3uySXGw+L1Rps
zkqsfUBtTBwYLNkwpt4CE9Wli2MBE7VE32IbliPBkzx4Vzn8tUAz5fs/XFXHc1Mu/A2Q7ObN8nKv
6QehsEmzsdWjkoSTeIPLIXC76oB1RSUaHBqP+RcvHrbW1sppt8X1NWQlmqv+BHqsKdR6I2ZtL0NO
+FHEh8UmGhbpwzmIeMp4xvW407Qp25cn26n0HlJC09RnQhrQ8+fVq5gDcpwFuMyc1+k34sySoysB
IBY4ndj3btPfeFkpQG1NcKN1cJEj+vx6Fk/bC0mzB4d5lFDU9rE4aY9HqJepNjnztfdhdX1ul10K
eIjxwbs7Xqbr5G1iafubILxW7SlXSIiY8si7R4VyB4rWb7CoeGBfISteLJ3VIfmu7vQpw/l8RFuS
mqyIqv3sPVkid+Z3XdYA4DwB0KR0jhIAiIyWzXi9cthK9e1bzRxQ4dq41emrNaMm3+doZ+SoQQMr
KUJ2NltKfezZKJYtw0f2mU4eDAJbXjxD75P6p2AJOpSYqidpntdsqpxHwc+LWlgZYL5wfyrDwG46
P9ft9BmblDs0fgZcogcDFtoiCzasQrYZm/GuXciDDqsBNjm0yD5DDY6scsyZFO4+gLanNIk3ldFV
JLMZ+4oJkE+qvlhp60A6dFjQ8BBwJisvSrnacGx9/HgE4VK+8KW1xR5AFUy2g9Z8zAEeizIC2z6w
dD4/ghRV/NcSU+Yn71f5FPf1RZSaRSTKYaDu0G8jAJ1CIJz3lzDzF2qypxch889R/YyMx1IGtUMH
9Uofgo6Y2401BSBM/BJypQ3k2Rz1S+pIPgUquQ3YPWEt9mXmUS6egZ7TBmoR+RI+NmsDwshpgdZB
mLnmYKKH8+xxzd+KEMBW3WzysMLOeXTe7tyabbPJ2nPTMwXyJQ0IsQ00JU8WgTqrZT8jOB9YBqnd
d+k+rJLkDkECdpnQNqkfELfi+E+aM7duq4LJEeCETd+CqfqBntKKSjNU0c6JKeM6Q2eQdJYkvcET
2cjZLx25Dy+4+qP2sDQl0p3YA92BbtFModyYN9JtUxhvGR/nESitLeAnH4hwyauldgFe16A/ILk2
uotONTHObBGJdq5huBtlz+cBVvUy0LAkf33KTsuc7Bt0K2yNfd3nRaJqjbu++CSggDZCoIY/vilU
L9L9y+ZDiJaBMj0P0/LP89tjA09DRVHpj7pDWP8VWVGzkdNityZk60N6xiQ/uhdNHWDqbzi/oj7z
gs2rLtqIFSXQsy707OtuP4ZqUkXnrM3bPKVZOjUsY+gKcK/vHtzM1bElN4MBhHKGy7c9mA0K7PLa
PZr3YdtNjfQg6l0ar97pKNi/5dfnFQMrmSjuyQjOQSYFTYHayeFPrjHeCAwvvCu/Zw43fNQgludV
VgxZR5STF5XSGVYp+YTHMJpkDiduW/BT6xFsim7Dy95foAHmXdi8If6uM6xy3x+GS2PJiqsYxgki
2et0/ypM/TL6pjgkhvhUtVm+5G9AYr90pH7Ezcm8YIeHNudof7aUwdBCS5J5S9WNSNRWPrSY/atH
tOXqGZuu+iDPSaZ9Pnok4M3MxuZ/1aRDvdIHM+0B8+FdRmPRaCRabU/PHtXX90h3Jd03KwHnRExW
Oet+hEeJjIItlJaemnMvbLbwFUm9eRF1owoBGLt6bzJMaU7HyPQYZXXSWIuSSf6eKBKpVLwWmRbm
zwGfk+sdkuFS0uH7xthBS0Udt2PkaVLFtyCr3pyZ9gf3eQwXRy2kBjbRvfDPzo7NnkY1inMjZaD4
vRCFc3bGSEPoarZbvej3fdDfUbEU31P9U6QqZVYo0olz03B8HIQzeMuL6mHpmiQ9W761De0KBDd5
6LNpCTAX8bYyzhphlQO3tAvpN8NHpNi6W4qJRl4ZQ1rZQexULYky56Cvcj/FkI7SFXIgG4GimBlO
8y/trSi7Q32T/WohEsXaAFFEv9uU7lIFf6opD3GGs0oJWZ43wxPiksxaLMN5EzUfewvkvWjbjz6f
4tc/qY/ZPAKd+UV69DikNRfvqhDR8C5yuqL43CPnFfI4sHVwExKpDALIxO6qMhMmWT0D5L9EX258
Vb7W2miSxZmQIVvkWV9dt9eZxYR5Htyn5+KbAlaJfzdfSJ3vkn46us5aUm5Grfzt2WK2rnIjJGAX
DwAa/VqHOX7RsYatSCJ1NDVtAECn7xlsDCWGUjIyPkYrDTLWecug+9B2t4YNjwwcPzqw8Kv4IJdm
iCO6DKSBxDwY/ky+yueeZ4/nDJeHGCUD5WiG5+voU3Tu6vgKZ/Gp9pU3XGSJHf9Xn5Hk/HnYDbP+
yVxHGsjFzBBDfFJ1KKtljAdsXD8r18BG9uq0VaOyAqiiLaxiGcgt87gqL8UNrG68OVLwnaSGV05+
Itcgvo1GuaP0ChE+hGfze3TiVKfY3V9g+hqby86CmZrcYRAoQQHhQczthPGcsrqq6XOP4hRGaCS1
wMbpvMODaQ3VbCzkvkCrdBCM3IMQ3Rv5WjWhA+JOT+6Xo8Az+N5PDtwVi6fw8Dpph5VyHWSQYZft
U/m8JhF3u0/uXwhzc4RlgwmKLlxBCzG299a670fYdY+CCuYvS+cL+IfhPQb/+MJnXprqnD1Cw5ac
Uu1EtEUkmb3HOUmyy203wq2SOOjYQAbg/GuXkC4jNVCOY77KHJUZpXgm5TUNpYtFkHvdwLCWdQ92
HRSQkyo8kbcPO1hWpxNXYj9Q97PXTuF61hAUUFKwaDtJqjsf0vXYhgoAnjm0KoyMF4jMAMDuwPc5
OYo9NclUBiyRFLtOzMleQGuX4x1B+eyPHAIYtX/DAPzBCKvDN4Y7hGjV9TYHVxWN8ROcgF/fZ49x
tk0gcDtcGztnGdL41ast9Nx1CL5C0aymvtvJn37/h88q4U+Snp19hs1CvZQBdVkgfEcgF3BECuSE
1xUZihg7C7qiEp4xzLqm6RoW5qPQ2dkYRQgie2cxLqRdVbAn/BGav+pbpvcdymg8XsyNpKh0Q6Fh
AHno6/B/cw3r7Ro0JKzZ20mXzJPOH22g9XHICrA8dK4EVju/RgRkKVChj7gxILIGuuPmlwfQ/BX3
vp+kSeccM7LrHP8R1O5X7ExPHHht+3gCPMJe4Cao6jrkmiCL/SlMGCcj12ZZPzhW2JABCZtBvTpz
rIZnruoO/Kf0W89vUktSXApa7dm4mWgdsMYgP1DsXGqMpNcs/vkRE6I1gPmuN89hnVfuRbQC9fmZ
XS3QBhDOjpOgVruQ8RsJwbS62wZ1u7cfjIR1fNsZ/oycbF2tv259umTn4BHi6cFip3d1Rqj2l3ZG
Xal6+iXsHrNDX5QwJEp7ecoeCa5ejUrX4pD6EANvvKZu87vEMpUlj0t90L2s1L+/xVSAyVsjYGuz
RLKzLgaD78MwzTcbgJXQGK/OVulHOzYMxPjGKZGcJAMDTC5xc+bzUWYuiUmnu07xdt0qMB5J6bw1
/zxeBOdgTTAz5qTJLwVc7+y5dzNxMg==
`pragma protect end_protected
