// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mNv1JW4ctEYWZHwDAeZIXCOVjkBDGJTiicC7eowfXaKtKet2uIgV1iXNRsutq8yH
AJYK3bbOFCMQ9jE1gjt3A7RFxFJuL+ElKzOPhIWaAliuG4+NVdhlVkee1vXXkVEO
zJKf/22LKm9qTXPS8ULEQ2jj34qZ2Db91KKlAMqV2rE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11792)
42rnbQFFdvaT6PUqgYerZbFeavWdEoGy/CcereobUh2H0bpY6XWsNRAHyBxHQdHy
FNaAKV+GicIlEz+H0xn64Fp2Tp/bfLB0O9iHY5BC8lo/QCaVSooZj75ZaGEf7R+S
FQL2PDJoR+pTVbBBmkrYXeTWGnYxKRgMFjuY2cPyPPjPKYlJuyCOY86PSWrnOuUo
PtSEhwZ2QCZi7g8pxGIlvxRgw1FWUYLOcrahG/XD0vlQIDo9+jG2ciUrmujZAYvy
3xIthXYquZK++8r6/zs9lXZHLNr5KJ2FqTTPWzYl5uHzDI7Er1jvxYv7Y74r0MM7
FEYFc3+1WjdAQg+PiTcpnEUzg+A01A1Kx6M6J+4T2r8iCyEZ25tgdrcmXQnkBc61
h/Y1nSjK3TQtuPAUdwUkKTuLP1c5wYlOsS16BE4nKGKzdYe11e1zunkHzzEJPaKM
IbtPjE3p6bHFfpxkiqtRxLzkZH7Ol2nF+EZJCRhWSkBfBBBYf61hMfctu0mwcZZK
C430jY89+vN8Lp5cy4Zes6XwEkbE1Kq9jynPZsxyL7INFqOzvo3EEy63JvOOSp5Z
lc7hMDJbngmE4KRc4tY5fhwMMVbJ/IerlgSsGZkLer7H0k0T3rP0/uew+y1Tf5xK
fmfGWyACg96sN9BBPRMjcG4PvoC+SWt+wG2Pv08R+NrzWgTiwLQvOnsIFvlLJzma
zalTBxVu5q5Z4mrGIvUwqjQaM2BUUyuxrICqYs7gJQXqvBPvDD4+mxUpKSIP18vK
D4zAEqgZOVR+jwCtedOJp23AVp0Ef25eu0TkYiDf7Kj4EmASgfbG0cTWiWu0adRi
oHyO6AtddOtp+492KFoZ7GPPVofB2m+NjYVML+CiwAeMY75fbIi4vcDIjZ/A6pc8
vSWxN3Eqwd8NyjOcrrmtEmXL5vqK4Dd0/9oZ5w2Zb6flnzCpJBHWd5ZoX9MBV+4W
GQgaKZ5fqhcka1qRNavEkGBmrjqN4+7f8tWZWYzBWoeH9A2H2/LtIStv3QBam2Aa
8Q2BVovl0aD91NnCIQNejRScbjA3YaVcQIYzHvtktS4TB649xBiw25NoRD9D2nkZ
RV+6HxPOCeBGGrk/FNdYB5HVjcBmKu3TidFNh4AGVkRlPLgho7Uh125stFPrsj4q
cNQQrOJBX+0qwqNNSEg49X+r77VoWGKtHQyWaQSTDh9qejiWdfIthh/WfGFy151k
TcsMo8Ufv3Rl+PHMQi6c7ADb2pNPPn+bjEI+zyUm44HY7Zb0xkyOVht5+nvLEsqJ
vwom+Zl6XTg2QG47TAUKzEKLfUnrnaLd56h8BS8r9GHDMeqrUTssbkRVFVGm3EbO
nZE+d/7Ap2mzZ55V1PBw3CILkXGyWVxOldazlu1DF+FpL+tswEAhzA4JD6jJlSwo
oK61lZrUke28i2lIvISlOX+A2RE4DtROV9P2HcqvuTaYep7QZULMxsIlIZr4xvqW
m8URiTgs//gg+I82tXs8zdOF1I8P7x8L1D2xTF8Btx3llyKU+0HJ8507tBf9AYMK
+SN+Ltsd8pIPnQY3cccYJ3w+VmXJUI3CVZn1Gl9rqsdkuS414hXM+aYOYA9wzCaz
3aTW8QTKsr5yG4PZg5SuTGI0xL1rr2rlxl8RjrHBlF0UVDuWODXgrWRXUQL0MfHK
Zzk/hxbB7JjYkn7txqmARwBLT+Lls3uEmGF/mtb61JB96CgcFtJjaHv1clTuRJJS
iQXFC6GvboJMi+X849E646AMnnWo6ds0VZiSqvRuMzg3j0EUISCZ+BCe+tAVaQj+
EzLEN+xzj6VM0iUbbsyGkodjJkFRKMAz6HT5jhtmVp9tgofDMimSR9w2C5lGE4kJ
e4jr+E7+845gsomOEmakOF4fm8YIzadDKnmro5KBk/bAeJm40etcWDbLNvvneFy3
7Ddg6dLKmNpUbxFOFyJJgvPQ+pMHKcSxMVo9nKXa9m5z2CmpP54jC2/vrsEOCbWZ
vZjodEijJGysHBvNz9g7vHXoL1BSRVlXZzdCUvvKZaYW0y0DjOAbr54dYZTB9HUU
2r0NSrVZVNj8JVV/srgeQ542HItXT3vOjX7of+eeqQic/Ma51t6/+c55ckL5zWnh
mXlJidl8BTWXvK/4xlExxBfQ5cDJodQREX+cVo7vYdClw7HCIP85ru5Vp1mlcb8m
FdULtD60tDkDuJT4tAcfSIb45+tWrDTojUc+NtPJrldgTVIlPlzfwuRXMF8e524d
fhadxoug0jRcizEWpGeymoiHKGJbn1mRcDEBzFu0vK75tQDkTslAvnOhcLqF4PkQ
RBqvnaSuB2swipFjYmnLOG6kpIcCCxTDj05ASA7o137S4dDfwFfHUxi/PTD89TYU
FP23k3wX/UsIJY/E6GiA+++kMGegBT8gOWhFAW6zBe+4dT7JTGsAoooHlfb0uHwZ
68V5zd/xSSkZOmvhhrBuJR/D/HhiJZVXKGpeqorPpgeWcVBkjHbeCuS0CLFLHRAZ
5hBujijFDswy5h/N0OpSLv3vXJ3sg0FrrNfNCJztcf8PN+S+RgiMXS1HH0Rnih4x
PUjHdph3hK8QNm3DwHi5taX4uy4Y1Shs9RDZvSFHGasonH6n4vaGLLLW3BR+sXzt
9M9xSdW4Rlr/4GPgo9KeQgt71NLf4rp0FEF0/wQYkHm25NtmAv5+nOM6Z493DYVF
tpugliXaAiIEIciXH1bm3bbtbKud3015cOVwWZSSr4HbuQV+NwKQp12y/J+7iRlD
0XsBS0n3PHLWV71aRftYm/ESenSlLQe/uLTi/OMClS96IYuTigXVQNFaw4Rdg4RB
u5BtCqqS+1AAn7nZpwZ3t5bQd9VPur7WmpSWeYKfRJHb6/tVorz5/hMf4GXuGoFg
FwqRRDBAEtQ/6GYeugvTqMwgL4O6nmsXGCqkcI9/sEDjWS9SC1pM94hXpuTK2taf
eoKJqs6BVMlzLVwWWaLbcBVQBCUk2jj4nnozP1janWrUbV0LWjCkwjtyOqUWDvEb
axDYwkCGP8mIKzv1pGNIogHzjIS6i6gxNCfw4i2pMR/A8XOL8A6XU53Ro6U5bHHK
Mtx90NdHFhC8mR9zrSuV9/hmM/v1v6A1/OS1+0j9TF+/mqDrny7DCc69Eg9CO1KZ
rmmfaYbnotkJqxR6iHPT9VdLnQo9QPvNNx3aOanW046e8RSYmVlMxHLADRyzaMnZ
sDKp70vGcxeby+DThzqDiN6zq/ox3K6oWs9CU73NlKYczVH5S4XwiviCCBGnB7j8
aQVyYWY5yftMyhy4nZZkSXs03JK2mmkwbj1f56hpZ1mnCCCk4CgoAlPNI3bes7HZ
RkiXyAxIs5JcPyADjBPSnTH0se2LjLcWgrVWiziNDrUygZx0iLGl6zxg5pLjEymJ
Du1j55lc23BNcZ82vFw5EgVm7DdwJZOjhxJqQUdMbKmPv+8jgr0dLTFqa5SAkdsu
1cZZDIbF9OFE9MX4lSZXLAcYjNIlLpdpx2rGoBERNEm2hlghDQbpWS18DJ2kXtT8
Y+2rLbpjP+BcS7DEANV+vIOmoLse8y/Hr+wKQPW5HJbW4sp0b2FPGS+ma1Uf1hoW
aR2KwlXWjhIhf6oRBH9bRGEw9ub9u8kYzzfGsTLZmMTV1FijmZz7KqwHP5IKRTKx
TxwKI5lVm2lkKyq2PCJpd35aLaKTDCi5sXn3okcobOLs2Yu65AwV20PDZrDLXyN1
gHU3Eq5bHiwf0eypGXbYTbdR17B2MR/0IA4/wbebXoxL9+vuk1Jl/7tMsU92IPrb
U4U+OfhL7otEpJJdof3c6J8f5lV7MjHMGLgia6YWBtk/ScKXW4powgFrpY7GZx+o
atFIqJta3M7fVYk4qYE5MfywlFx3J2QGZbyKDukrMeBFa9DbenLfJV7GVwXajKLQ
IVB6a/mFSymEqXDZaYmyz5En3jPDOdtJY1FVK7ctwuaz6QllkNVuxnugJ8tHobBa
WAeb0Asg8uCZ6FCL2mr4Pu7hwFpd7sw0Ddgco3U8l9Q94T6KU7twDL0RZneBLo3q
uHvIhVh1nTxQ2WNEBxjqKexQ7mq1d7JWCsbsn2BqprpWqeK46yMRFLLkI4UXPJ42
OLaCkrFz2qakSuXpo0CZoUTwvLnMcJCZCGZWDX2FZMWWtPKVL2WkQbhsw5ijyNhu
cw0vhnJ84KTd/0uOI+A6sByuj/cZoIfVDe4D0kzHbxuVGfYJaa0DWNnIb7ZBd+5O
hRlkbNG6oYxjng5f0RGy5AlJcgtCe7uEDjDCsBWU8Z6Dw7Q3R/5q1lbf3aDZMIS3
DmIvU055jlJ+rft43OPHucdAAF/VSV/z3gSLr+d2enavjtk5yq8LpQju7azn8nNt
1SrrMwFP3TjkQZD6SRVbhs4IINL9YBhBxV371RZXGeEWOCCIUVEBCxFRR9OC3irc
P9vc0YRHcd+b/kUb3qJzt0ts081gKrsI9AodGaLV4iEVbSUPlqbDsVjxnQRWGNzL
sFlDWXJRcJoo7k+oB7xA4Faem1pl79q2d6EVrXpYYCRmsV8+hPnxICFVk98/MrXr
B7Jjgo7OSwCCobKC4XRg47Zfsqa/ttcmm1bNQtoHtVkbU47tjvqGdRlFOv79Ix3K
fZC21QlMkGUjpG6j8ZxDvPdASU2z0eHKgeH3IoOgd55tW3p3QX4enfb0f/9J/VaT
X1TsUoyRm2vH+hC5zKHE7OeIgLVPlocQBdU8DZZhgBv9vWf9xJ83f2vyU/1XAPg5
NoDi+eXxR0WeHzMFqByeNgE9FIC9HhReEeEi0WgoJ6MwQ/yW/ovbkR4pDiz59jXj
YNyDZRjdCEDDXP17ten4QUWcIRR+YVvqoOyiu0LT+8D8/2uvdAi64KJOFu3A2eGI
s/p5snkTSxrQwz3dS6B5OwAcXcFjPF6ONdyMeyrivRDG/WLk2TsXTftKzKSvt3dQ
WBdvjySMfxe/CWkillOy+z+/IuzsKLsjrM1yWfTj7uWor1VOlU1AP+3g4yiQlvfl
gPgRLCucRHBt5Ep3qW2lCsFrH66/+Mhb89idetM+zCmjZQEZFg/KkCtbzP7zdyFK
Q8Ybj1VDqlinQ0BHX0u0nUFSFCNwQL+pnHrCFmoiO9ibs+tLWsx1vVFs5q58hxIP
qem+wvRr4BLKoXpTLz8cSz1tMQ36wwJNIDIB1wASGMM20JRFEbOVgWxqM+onhBzd
ClzFApgOHQRwOKTN1IDCi4qIrcEVeAVqlXsh28QqlnsYGwbhplyXkbfKQD5f8pcb
+3UicIYfb97CUmegwZo+MycIsCgEGcs/DnqL6FHytQRmMCwiScbJ/ijoxAfX2w5X
5ZZLaqvvTzCpQGsy2n5BUTAWfqZJeoW73jIYtXPejxc13Yvc+pyLbMnyANW4xCtT
RQDJq/mTVaNsEJEygd3j5yemFQ/hMJ3QlLPXLmhpWDmYjcJh48Si1GoeFBdLiK88
ErbiaxhgcV6+e9UWATNfSYIJdfYk0KsGypZDtHOXsDWOf0iV5OVd22uF8D/Opoxj
v1QU3g6oBSCRL62N42wTcLX6qdros5l4+57xiHTTTOGe9E51zdbNYBQ7mVhbj6YQ
DMXNPryllMWGDjWH+SRTcOk6wTIf75P9reRtWUeQ8H8q8sNS2xHpehx3D2LC+pIa
viqJXGY5w9xqSlFswcVXnl1iREpn0+Gdu10hl6umjKcM6xyVrB43Vzoc0ctPbtPC
01MVBnl8jodK9JE0CwT10l27fwNNassm/De9hjOUWJX5PMJ00+Y0ObCqHJ3+MYoY
b9Qt0U5rR+QCqeBDbigtAzKzEdwNA4LzNPapdGqG1HvUff9DShwOR6qmVQos0Ym/
CVLa0SaOheJwlvJrtAL8nmjVEXGJKPd8tA5ww9XB+HOUJm9/LtnLE9z4FL1rgHwQ
Px3GOa8HIMxxvrGtffFYio3vcGmdUbiQlfwu3vOAuVILJEdafim3egeGv9sZrQUR
PvfS+j3CX6eWRVoolFnu07NG4MXDfioomZt4ext1Gk9LBCH8s5weSzTmd6WOVQua
KxUWRpTYdZQYzY8MUnu8covtSVrXY0S4zEvbRg7QCa4AZGzW0vBH94IZGKieM8JH
P6WnALJqzIzj34Kql0FhQFCnEUvzJtf0SFhDzYKOP1KnnLJ9QKfSTVCRet1p/6ID
7cQovLNhi1Xkudi8huI/1uAcftJU/hjOrVQU9aHphLi8vqoffx80t2NaHumADJO5
LoNtPc9o174M+uuHgmn4X13acuC8IL1UOzZJZomLsQpYc95hm6lvMY4Q1VT4eith
q5Mr4UEAUVU40jODzMta5/txRxkk2S1wVQ0/HKdAY/oKPQxnjvPByVXRQS/BpKBX
n/dmAbzj6doaXfSu2uQGKka8SG5lSjyaxS6Rc0B4YpkuLwkP2LIXNm9TG7AWZHfc
wbtI4m+wnOpYg3QmwxCJB2Yu4B09lCJ21q9ftirBEQJPRqV52p1HZsy51ekIUXyo
07J9aUMrW4V3jL4lp/JHhNgYxeIqfrWVP27NS8Aa+XMbhmmQnC/gEW3rR/TZgLcs
Wt7xGg4C3y3ScCmXsxQjU4dVBvu4+ezziuV6C1Y9RKpyVjOncpepBChpItBqAegS
1Lg82xx9N4GHrMEE0ab0Z4Gkykeik7DHP6Soo6ctnsh8008yBQgNe+ivvGpsEzXf
AlBocIsbgtyu+rmWB0XwXjAIJSrQfKh5UzTlCNx5AxQHXvLrdb8VcLM3+ZXtINKE
XDP/v5JfQkDJDneTr3vANgYUlq9ut6yk6gTTKCvwjcKNU+LdCDfWwWE31LmV6Bcw
rLBdJLp4J9RJBah5M5lZ0oV6eH3MVEFJ/F0KobXsCWOJ2J3TUFSlOjGc8VMaJjQi
rN0GcXQEueDFlb46Nl1XjkxV6YA5S6Qf6iLahyOL/L43r2AkqSWWo2rYuhBiI9Md
GMGDjYV8IDaGa4F46ngEmOSQTEIK+Yeiyhog0w3ozoltOUNBGousnIf1fn3iXYzB
FwGph07DNnNF2fBxCq55kmXgGPA9WTuIfXuVI+TeHUVPizg3avqZERapMZ0gl01j
32Li+um9SmcdaHK1twVJ0crI5lbV4wP/p0OI+aN++HIuqUBF9LPf7QCXVh9sahpS
mtflJ+npf3IXmzJLd9ErctEHEpWp7iAkkTVdvvGyelRJDaxK7pQOMpaAA68CxDEt
m98nHPJHifw+pnSIiQpRPSzh/+z5llE3tf6MijZD3cyxhUZaJZt929wUqJaSjwsH
bktUrkhHrMJyJasL3P/HcV6v7ymz30wPQt6kW52vb99XdoKPoQTTcshbCRKrXJp9
sJyz1Suxnjw3Jc3zYTZcpf+yBPH3LrdVs/DyLQL1QR2j/Uaep+rwuGJZUgMTdukV
McaOLBRAZmSGjyrsCQC3RVoPmuBIhfFl7LSnbx/YyqOtcDZFATDytYD4ZjjfhwuC
Ryn49aFKkzxTShbS3UCwJH2VJ5WO8TiCK97hzNLM4qKpzNk3LJ1VzsTgOpXzm4ZP
eu3JCX6VPrKWzpNMpC+HpMXoZjzeKpYaOIGJ6YmqhIuNIRYln3LBss+ZLKGAcbnH
dIS+CidA/PU204UdbxKEqiScc4Bd2qmAJ518tf13uEvjagu/TZUhx2NfZ653eqj2
4BAO/Gm/diwb5W+wQxaoVB0bxmWdQbVIF+rISdRGvAG1aOVYQnivnSq4roSQLnRw
ypPKDyNPxMWwN/zOXjjsfdtKT11xtfZjNpIx1i74/zF/DjS2rQrsTBtaawWD9i3o
U2rWaytmrJS3FT3vJBjeVHcEyxuzUS9g/0udMNinhwfhNoAmIDuYC9CW0RokKtfd
JYOJw5RQZAzBbqjGOq65wOxSmHbUZ1LDk5NGetwkPnfQebtMNWeIXKmbUqSADUW2
CX4P8Z5aSnwGpumEHyDFSwxOiIIipE/rtgweeQHzmsLvd61Q+rvfOULqMryECLSo
6SkyOGCYZsdE+vJxZaUNV5SNFwCKGmVg0om7esIMiVhE6TIgLS89vQUlvFGyHkE8
WPMc2SOYFLWPlQJHmSs2V20Mgt62fwGq0EQd9xZ4yO9LjB9ceqymhPuoJJ7Gx/OV
K/+9RqHvjoPCay5H/rqR/Qp018+E0uaHx5cwJIdvenIr868iVif6/xvjaKqzVpJw
cstAKRkR+f6D2L3u7bmtSj8cXI/wkSF5+6okNVHK7tiv5gBdjdVea6cJdbLH6TkK
XUQa9WgCI0lcEYleGr9cacu9jhnS8HwY5lPWCC6Xiix5hal5n5gvz9AP98uSiV+P
nXF338crygJ8LlveHXb+ntNvHs04tWtufbjisgTQjwSsneJz9XHsZRI2XhQ2mCtD
K2HNCEfhZV7MdSSpakqHxbjj9jSEFSdHC/myH2Wz3nVwZcA/dLMctBtNnKqM51iR
mOIhbLA8Gwq7cpUVK7paRC9RkRz3Lty/e9LnaS7t6cIoCVTNiqHgJ/tGSkiXubo1
fAYc2XKN51/M+ZHPRt5ayeUCs6Q11IcbGAqhRfKqLAvlCaGFtbZ8iKO3TvBk8JFc
bHgg0yMiNnJM12jCAmO59o1l3GXgxxabxT5k4dADV1HQ4c0xyToS3i7yCxmIbHUB
33AFqLmmOwvLBrmOq500yWm93N82UIeTB4KDWG6XlHQ59R8PNlli0LjD78YtFmSi
s6o3Pt4F3orjlnu5vcGpbzTYNuPpn93/7dtXsNmdBRRGswUZKx7fo92zv4ENYMpv
rnk+7bmynEDXmQgC5vm4pTJePyNFTr7tTjSjlTiz2z+pkPAb+Qr5xR1j+BaMvYRj
EuZm+hLpE4LD2p6xwc4UCqhKwq9CMC8DubTISieJTu6UoTi+26gRdfRAty46SXsu
/A2sPCBSMIzdrgUGGQUP9Gd/SoSdqivmw7V2zNyowxJ/9AEd2u2yd5VstjKIH4oN
8lEYjbtui4cJ7tiAW0biWxZXYvSVy5L+z2KJpWcfT2jdyisxXFMfx77J8TBcRFjd
YzJ52WhK4WsFlu+n16LBrYS/63LDIeP2iFxZDe6ZvgAnUC4JS7TAr/TQTwzArH7h
Cc9Q3oGwkeE5ghzKsrsKpfZlLV67Y+B6VU/TasaqOHF4ZrXLmuOCwBOBtDAUeXL9
L64UJAWgHQcUiNRrHG2VSQ1zniV0PVvUUmNABS2oE52qcloJ3vc/KH5PodHzTJUc
xkx9OXJaM0XnskDGtO7PEremhhRYHUAGMdW8eQ6v6/07W7Hl+Clpg2zFTM60q3a9
zyUvDdK/UmPuggw3Bb8o/RmCeU2rNetgeLw7dIwiJ/ngZ7M6Ps4KUmX+vJpHZaR8
8Q39xhCOlnN9R9qi+nglvmNO44B/YsK52A/WvjpqJvKt5fdMk4iTVD+CtMWQih7x
mCFNHVM7doiBSq0EO8WxEKw8LKALTXVrwjUDwWm4dV0aqBW3+niJ2qeVcA19vxL5
XxzJ9Pj+7kbVvKbu8o8/GqjkDkqAzj1TFUppYocDHYpuY4en+Ru2iPeTrvdinUsS
iPNDYFwO13wvgnrdMaeU8YjsSm5PwD6K4ce1J+TbjQPVGQ5fSfQVVkVrbA2dgY4F
cV5irpHMZqGSffLW/aYXCjKiJ8spqqA9z/S/MWW9twZD8o++r+PRMR0sUC7g0xk6
oQt3Kd5oCCB/Jm+g1eXGPyPknxl5FXGcLsb6tF4IUEXNei/iagdEl7CbsAYdpRcF
4lMwulx60VV8EoiUybm1FtW557Aa6styDIhBFxTgZgjw8SEP303xVzEFgHtUZuHs
jc/s2eTHIV7JAtoAFQS0QRogLidM0FN3LWw3byGPrlMW2Sn9eITNkHBaA7aXOvp4
h/jVjGJ5Rhv+to6mMT96xsCcaR0n+cF3Y6uat+f7WTeu7qQmgLXEAwlch/7WHznt
NHkBAHxfdrIPcFzZ6hQVHQpShOEefsZVZuW1HNgrkjDA7KC+vaFPT3OII/YBkGIZ
bT7WqRh+EIvM5E7ds59CUdlMJ8p1nww7CKLo53fpgRQqXhqnSimpY1dLlcN2OCwD
MPBI8rB8qBvAKmFjlbZYAv5xkb4WgAx7z3bkVhr+lBjbcOzYFw4qIfpw3J7Wi2PK
LQ8VAb5MqplbW8skuv4uUV7vbVs5l54FyHvoiCo/0rnxk2MO2KhRgrfbxMdwaOri
AzuzZPvbN1urZ3izxKl1tiNuoSq8962SAX+Dk6H8exuEsH97RRvXocM9Wiaw8qJL
/eqEyIPGWwzuafhSAEX3cHxg91x6mb5JUdOowYIh07KVWMIgOkE79GYoeBgE8U2u
ZqH3Yeo5LUXaghWa8tS9OhXTbO0NsinCOsw+HM3hBcTzF/VaEgRG4BQMhkccFzQ4
I2wCdvH1g8vWs9apQgGiukZxoswGkSt6g9t74G9SxSs5ZQiB/l7lT3zd6pq10Q8U
PXjpdOzPkZLqgQk1l3PYXFht6LlxRrF1sAPDVwQxsO3VvJSR0YcgNjBXathrtbur
SlYB02054tmknlmA2G7ZarfnxGG5qeTwQtxjsSzIxPyakbhq4wXH3RXvO0gz5ih/
g/0nCZKSmnpWuS8HjdRazuxJ9MswN4bONBNaQpYjwYGWgHqF7Da+E+sJzeHUEi3u
aCCD3b5Y8Rh5ZITYkGqC/s0pJGZc7A2fWiHlS1iSw6GdkSu2fzB5Zo/0ECUV/QAp
MmRSFV+MxXI4zwBMwzd94nnTnf63eodNygEOAF1aC7dewmxgMgynTPu0niO/IR0t
1erbDS9bFc5nvhESLM+j+0+lTKF0w0Su6caweBZYSaPqEjANXSEPOKi2amrSMfrX
UvDR9ngfknPYm+Y8D7ncwoQ0VDV/lRefmUm+yA7a7pgmWIaEqdqGS55/W82k0XJ8
N44pvh670QA8ubmsqNAZew/NCQ3Nw6iX73BLZD66pSMFwtcyo5w6R9j6lyRQCFDK
6sycBXXvbHCaqkhQfEoPy8v7p3ASHYMSifMhmNYzWn7MKMYEVoZqeWJtH4FwvAH8
Q9s1/TDzwbjLPsNppXCouN5ir8UeBB6CPQgzoOgSexa/6DG7xCBBEenjcvDrPqRf
+WXwKqGrE7U8qZKHRkDQg57bzj6OYOsxNqYaDc7QhsTwoIO39pFw+Kq+Cg1CSZVo
nGUcEZrLQsJpF7/ULDDOAnisqefbeGZvJEgMzjNVlooHnNS5ji2C6+Mveb7OZZ1I
L0Cjmb6zGdXIrcIkT+MFOvXjkcV5Y5i46D9hRyM5FK7Xe9qXV2tUE36Ap4zU4Rut
tT1h4NaSoHM5556+LE+x9LizvQoY3PYFc+eWeRTn5PWsbKrzdduj9rPsfUKanYoH
CGlXpDRB/wpJ9KnrHUW6U3ce1/Dbgh1bdZYEZY5nxI1PtkuIrm74YqHMLNlCX3CZ
5nvCG47k4LoTrd/YaY892fReUfW6c0IrLKPnThCg9jRpNlN/KDNS60e+ClJiygv0
5Kchegbka9amVZZdIqw7cqojF9+5XRy2PEiCmSx7yORrjKwJSRznMNlPzrrCp5uF
8fIwi//6qLfBIF9o1m6CCulXmbawZ/Wi2TFygqmhCAbBs6MIcAcDDbwhzo866FK8
VMmWbC/EPmS8UMhDg1+dd7WLm1n70F1gImNqvGPvhwZNLJNpwn9Qd7PNrPXIgcpn
+AKEkb2S07/0NiAr7Gg1bUPeac+oy/h+3NUF0ZIXd3JuAMYpUl1BqlpSzzEcNBde
mPqb3+w8Yv+Mn8lqsRmwEsK7YWongjCKcD1FXcHYrsY85LY0oXSMWtBOPmv40QWe
W8CuL0rpM+ak2cHFWdOAEb9FEyBSfbN5ekk7OtQYr/D9fcFB2u4/ut0Ex42PCQEc
FqRhTGS5oyHlxO4KRW/HvqTT7aGQQoPWeU8UH/BU4CMcKtX8MJczD9jd8wxGhZTv
xZ2WTTTvMh2ubg6KHm67uVhmXIcX0cCxaWhYI6yO21+SQe5w8IOsAe5d48PZvP0p
h0xfQ3+yi5TBW7d+tvaTvuoaUgJlYcoKeKdz5IqVBqAMMnBE8TQO9x6D6wxpsmSH
LH9dCs1QPw5QEi6Nsqvp0702kDeaCVnBhdInGEcbAEfruPq+gaFz8zJrb2YBNAWs
cgTLj7EeT94lQMoj2oCJjgCicGsbSyf3EWNGM5VtyYIv7ex9xfqw7Ch4ekFFhaAE
KCOZQhZWQFjfh97PAAX9hQro1mFh8ctOAZSLxFhQ3eKNIe04jD7PjcrpRfi0LiMx
GEuechMLmhHNWnqJUTTd4wiEpe91w5Zwu1tCgSZxsDvyrsXCrTi0kpcuuyyxTlpf
53yfZMR3GWyK7kU9bAHSd8dZfmhL8nbv/1hQiwF7cHo6mep/WXEhg0m1tlciZP4p
EyqB5LDRohXBNxToIUZWeL3xp5vtWAa3tp13t3cXmNOMM4kjLTE6o1I7YIsmfCo8
RKYZ15xiGvT9nIJxLFl74hhbnOJqt7sQRkPm6yw4DB5VpwGTz3rtCGC7/4CFtqKP
N2wAUIj4AVMYIdRnkWqtu6PuKtJeSy/mT5A0pFHWEbv/p0Zg/CB34vScRiOH+wSo
gTwZYjrEmQf/eY3EfFtJEuuXHO5odx6dM7fiH+BcsytWLGVHHRQfyiXdttYtAtTT
JtsGZeK6pPE0mdPD6xKAawjzXWkh0dj/SE7exxs4kwuSTYow0vYxh7CYCEFzyNCH
OG2Uap4p5nn1WhnZIZXQEoC4GxSV1hSwrR4zz0JeEHlPF5tPm78NBnnNWh1uTo1a
B9cBKM+tc706I0RkXOmwa85gTy9J1EVnpa7AKh7FXoGGffGOhVb/UPhHXXZBTRgQ
nFlnO4OC600IuBzaeDNvv269erpFqs0LcYrWIx7lJjTcdXXjVlJ1bu1iEmiI/aR0
azdIHv2EEhRoGmyMvS+ukQRaErqGrwnGjirH26NxlsWW8b8qZlrL0ltJkRK3i4nq
y60s/G2idcSME4EJNSvL76Jb/wxUbNWjwuabNklZsBkqYbXim6oGhJ7uxmOYAOUr
j7NlJABFUHuqzwrrQURPpjDDjwL6f91axKa1vUzR5NSN6SPQM+IE0oeL2kA6yqlX
UxAb8Lv64DUFi+GT7SwVk5Z43mA1RQT66WXgYQQlEzNeWRcdMYBMCVrM2X/yLlBK
g73Hs93EY8Vohg/w+w2s4JRdumJ2J6uV9Sz+FJqt4K2NEdNR3Fk+r4o1e2tArOwn
YYtxEYz3Vi/tMNaCp8w79I8Y+ymbrdVM4Q0lF5Bj5z7Zj6hZIXXpJ7njTtLDAbcv
PLCzj0fY6dh8b2VQwK3U8ooTqreBd0Po2T4mrmd7rNVmfXyW4xluMFa/K/CqsPAv
T8sSI5Pw+0q0A+0fKqcoqkMExPUliqDIV6ogl8ICPVJYYxX5YYOfogw92UpI1fAQ
5R2hf+Db5wSShtnL7eMVyARrFESyquo/AMXpv2uTJleyeWUhRiZPcnlXiWCPlRb0
6bbz9P1RwwT/occ625U0k6pRqGObfwSVizsAXez9CEiUUYv3YGQqjyleipRhWtJl
M+yY3qyklRAGdrkhidg/LKGMP+WV0swizxBBgl4Iv4vrl/N+/EXzJwPaaiYDRtcX
XWk0Ny5P90p8oOSPgLijDYu1JroxGx7XA2l3eIrsFGXRCdNx76VG3QCPDWY/6iSi
goz4X+TsHTM2RngwUrlF0XdLQe6jjF/9lYQ/Ltg7FUWeYy8cyJh6xVZuFfnUsflc
Txa71Wy7guExqdZXWsz4bwvYjxLUIOkqBmn5e3TOI8pLsIFy3deoOka7/sjnoFBp
7J6aDomxWpXMceYJZnJ3ReBBqaPbbA5xGF5r92sgRv/L6fFXwJcXoxORpj3xBx52
Zq7vTmF2hmbCfcJQ0uK9WRucR7Exi8+VSj7mkV8cv5Um0AHO+BY6iRCkBqqfmTq1
JnFjtBIfak3U8tmP8t/3nIAN2r3baIxjX7mug6SPA9FaXgmYrs93fxq6PybR1SSi
8PE2f2IvkKWNpu/2li3iiluMjoPQfNHpb/QfRjKDxT0ogcAIFNxu0oKGzltl1ytY
CmDGszlAw9XYAkq2gMycAiiF4zoI0IZ9TyoUP0JqcSJnqn5BB90QDwsHy3yCdVOF
SOYo9fFnMixFW4sEP0X//HuG2nB6DuNrXr3Rq7I5tW2W7Ds3m8QYbfaSIgH1dlav
IE3ekfPiq23diea6IurgpHFYBlCkIUdI74HUq+t4kb8DGyN+2VIqmSmgtka8MLS4
ry9gpZ418LpID2xyJp/K51RPjJ7ICyk4I/nLjg8zd+ypz36TfSyY1BcwhpDbWrws
PxHxNFvIkYWWReOBh8iJjJ/pNo8pVLTV8kMSCHx21IblrqqZj4wslCDnqvY7Dacm
sSemU+o8tIBXUCvZK+Oix9boo2flv3etgeBDr4rqum8eT6uL6SEDNF8CkhQ/1SDX
bldQ+JLg2KVqdklRGl9GuBQ3McQolsOX+XLYUvtmKfIfD9OBg6mngMzyoXWPvMyC
poabp6ug4X3xHzAAIZTIpbn7/OjPhSAVgL+oXDOcSCalwZVdJuvV74ZNOMogNiBg
2+7wLWR65ooPRvGwKntyW3GgalA1BevXqIAUj/e0XqPbJz0P8BtC6KZxQZbcZpWx
v0OZOZQ9yDoHZFrGnU3VrfpImZJ4PATejZaVHPkrf8r0L8YGf7T8FyF4Zb8PDd3L
cPBTV+TUHYlGrfrpUZJ9fHNfJ2zqMF2AgNWj6vifgjKKTsTHHCT5QBWythOhYN26
lOWAxjiwPcM9PHj6lxkZ3tsLrXOKR6m1i3y33WluYt609z3xTFsD5FZ+vXejxPGP
K+0f0HBdQu5o7D7Bg64jNBJldqoO6sI4i7G3yaiuSKIZdZmVDYUUaiZ0s4QbP1+D
CgJ3CRu40EkFKmnTBc+kkwzOBHD68SyQ+eH5sKJqE/diSX4CcPwTuT1pgNfnuTdt
uKlqZawgVol1fUzNqcy+EkYmWRwum7Ft8IxpfQIv/il4S8jplv71dxo9zChSxJMf
BhAxCFxi1GtV0aXleJUSCNrmkBS955AAsl7iTFiA0EFaNhaqZdi0pEcENfQzdmmR
mkBHgjaZhEpHUbpJoBKTMaA7nkF3Ur06O4P+wYbC/NFMRlAlp4xk8jE64R6rzt1F
tGXIhzVjgQhQQT4+eC6FNt/kBOJIuK43EUV8TQ0VssbYSg5YNnNAsV8EGEcpptro
cuWXKOzKa9K7VYd8JNBWZ9lJZi5WHXNeDHFk7wF91oWOqUvjYXwCg5bWMm+XX8aP
MgILqLSLecxcFN+zx2unJPwZGv8ZbBUndPci0eBIGO/btaD8Gpzjr+wHt6mvyE6i
95DGGIj7HexkVisZym5RWYuryBBrgwMPPPgr97dfXrhAmkUvyitMc2QQzKgkYo8P
FvvjZixdRYMKAMVhMM7lJSQRsiccVA8VyPN1CrHPNgE8EaKaO6gZlXRPMBe/0oxZ
RxCZae9OPztZV4YamW+P5r/C4ydo5y9znaq47P+jAbtcYOLg3aHObKR5WbXSx6IW
rP6TOzng3QoEDKS/hYUpH+b1rsBQZOUxTWny+6+8lXZmgWNxyx0DhsW1xXNl24/L
HHYy0dHoluTo8p3eONEjZLlsw8lpKYSMrd8QLp3WK6EnLdSlG0iPAOHt77SfACHq
Cjcp1cRxVe/i81H3STSbdABjGcXRmsGiLlSo4ePZnWQUASQ861HpS3ZfU83A+r0g
no+gIuEZD5tualnrB3Clt07BBlEBb4ilZw3sK0ZLlVUzxN4diaQSZItqliHrLW7Z
raDgeOvsZyIPm9uGHLd7h9ADAr3lOIz/YjaHLxLT+xI=
`pragma protect end_protected
