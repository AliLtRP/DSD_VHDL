// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:42 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VPm3+6O2g9gu3lVHkigYbM2l+1nT/3xFlek2xCk8O2JXyf/MsBRo2DpuftQMf24B
2qa2GONACbVGF9KrqjJWHUOQgVXe0aK+fal1ZFfCmL5/qTyh9jWarW7Jml/Di87E
Ihlb7nE8jP0o4HCa7+1V8vcQhkva2p4TqdNreVAkdfI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3840)
nKfTaTnerDhbc4ebT2wkvCHRqhO5bci4SARg8Kor1k2zjDCsGAdLbVRPxvi2r7Nj
qRoP5XnpLsipXZKS4oZ/qLIVAK33+fQbUy4r0rmojHrJAccCMdlEEY9dpqDbiIiQ
o0nqknoEMQ4cBPyAv5PNOibvU/aJSLCJMdWPQipMuF48/PNFAboSeoUrRHZV8I21
qlsQ4tzbFjWI1BqhlE+CngauxANNZEEGyaYcyHONeqdJKeZvPjyQawiMos26US8v
fyHdwtk2rfJc/+MBdDtf3Xk+On9jIZpV8gbBmK2WCrZVOK1jYhPUbsINmvvDNnY6
M1B06MtaIdSn87JNQuctnxlSFiUJ/dNHX/gNO5GanoBWAfAY2rzz//0dnX8KClUT
dsGTz2iqF4gGV4fsldFz4vWTEjBcRmTbKmdZCDRekUck+dtOUK2iM6hCsTYgU7tn
tdpCo39f2S+UQh7luEcOMpTr4apyUXkglIkge/dVcTbmQ1Ho3YfMf/C1GfzWfWwB
GV5y37CfiKxfy+X2MhCqk1LJaEf+Hx3TTzyD2oCh/5rwVFyX9h+uH6BqjAKAMIF0
1BDDMwwaCgnKnOdvuvqJFZhS5lYF9/pbO144UU67GiySV1MX4TUURmdv4Oo067u3
coV5g+CQGia1raI23TlcnbANVvTps8ap3XwnuKGC+iQKXWOUpUEeZ52kCdxxz0Ux
YBbzJ7sO5q++tYuyuwrYeY+0MjkDa5BL2jtOq7RcFAQnI12DceEJTJT4lEDyzUrS
SXAv+yyS12ZrXyOsi5Z4QTQuPTGT4mP/Mu5XsQPrEFjI1k1DqeKXo3dceWLNTSY7
iORwZlJQTNmzgP3ishVt1Rj7YT6uwoerM7IpeOOfqWz7ZqIMci8/075Zobb+wcd2
wSvAIbMp+N1t789zn9mnNVbLg0kxdQPOueuev95hh/z2jb7zhTTCL0E4xQrCKnDG
xpW3MMvPbJNDxk5QLOEQ9EjbVQr2QvaDkMPI54xsHoNzcp3/k6POhAMAN+niMq4I
+hXEbq8NdHT0KXHjdKIQiVJXos+pA6rbqNfFCDZW7+vN7eo7Ad38Irn1p/46Hc+f
ql+hOs4HLfnbOZ+stuURwd30xd6sLwtrLDu50mN/LBl9996y279C7Pe00/FspGl+
5X5yaOVdoxOK1mOZJNiEVLl43fJbNHbPfZRT0CHm1MN8QRnyWqrUNgOUBHjy/wCT
jtrso/AXHQW0cv5+o7iGw8fGR2rHiXTPEOzhVbAEHJTEetzwjtMN8aPbdbr2PVYD
ybMw3+SkUvMGXy665Y5cK8moDq+3dKldRjPHUPiqT962linaBuaimRrUjsjMkPuE
asaUH8NQ1V48/k3Yf7NGbD07etlLFedQoy5qjcGmT8cfrxalGiDm1SsSA9Gdao93
BEfpPuWCOLpfShvs2l0sAVspJH4SVQy6D9bq2CJ8lXhmmWZT7qlujEBp5v1HuOKE
8VL/nO2kFdPVBCmMlgfDIFrNYrK8l4GprlS8qUKs1VvHOt+xhEXRznsWfSBMxE1m
WPfNJzm+Lg4XUALJkGgbqBBmE538WfGkNSVKOBJaYQVUKUavZ5dd7VHDFGyfTy9T
MJQatcav7ceNbuiisoHhoLvVBwrgy9eGtOGHsDQDCAVFK0MUWHK9mdc8tOxm00ZB
DflPUJKR4dW2FDhrMI9Z4sAtejSuWrP+AZKCpLbS9NQzSObypFV8LiOMxCwzZbTs
Xu/q8BzByZY+ZflRciY3f/63FyXV2u7do/CsCpgR7u9BcjU627QZwb+xfmRTMpNx
7AsWsZWty8me/RChKy9E8UxiHL26Lqw+zNICM9mHV67lRtb9V3l5pCJ37Jm0DxCg
rfq3hsk88SY/plDIibmO/0ljQrKC7+9uHtcHLBSg8xFfroWsTMKAq+Vf/DgQzhtS
fpDAcdbPl+MVtw17jzHkeE534PtTtu/eycnZ1waoZYyIcrxy47jSZftYlT4l6C6N
DpbaFTxnAo8s7+gP/+ziRgySJbAeRR6LD37jT0xjubzeMAARk+eT5aRXDKAMsKIF
qjFwh4VmmIJJ9oRew0L/oQ7v7WGWdIDKdLr7Vidh53zxRz6EHa+/p0dayxGiOtG5
n62Jy7HFIluvs/OQoKzbWMGU0MTgx+RKnMS8kDcAB4jnRRnTfETgFSjmOzskPFyy
YjXN8FXRRQiNhb+KtmBj9lN8kd3jnIpPucgOQdhdW2uSFmSDOofrFQv/pLVHMIqQ
+qUooBFfx0ok3gFinS98FvH6/W//FwQqwW5+uBn1LaU84pX/YY4rcYGCIrK95TfI
rYlf2cNyNRnhfP94eQXQ3bvMzOW0JzfgNzXZi4ZjqDt/fMiZYYY15c9En3WHCGMP
rzLvvdsQ5LsRl7sNFX7srwePD80UwnHTC8Iu/nxAEDtjObwvzj176pLeDpR3oaEu
R+Cut3dOJt7mWEte9FpZUUXA/BrSneF88HR9xAnh1GQ4yiNyqj4HJumHwnLhYmX9
dGBwlEe4gFB2iqV4W30nnBKGDKmCREONaZqeYgGYd+xbfxfJBWkYrPTJYiY7qHqC
mwDkSTWCA9NgWWoLLJdmRZ9uzFlJp4EP9w8ynu7x7piIhpApyA2bLhGgOVzywk0U
9/SXHdCCqH3fgMFbR1mzmbxpDH23hBakagFAFhfRPCVXQEQxvxLC1p3wjr7NWAtB
D2pmSdY+fubJhg/mw5sbRXjZEdGAcxJRwSdkkfLMQBKYEoIKii+bz9bAgdMfvzAu
1IAD9H1TxCgtdOVc+J+DtCUAsED+Lf23YL8k4JcizyJQKkJ2iaw0IKDfxX4l585g
Fx2IrLZ2EyneUBj2EVQUDZabvfZ8DTjYCyQF9C0zh8MMTjk3GJ6PPqV83KtLiGVO
jt0qsaRxywpMn/RPbk/DtSZfhtUqNvOe/yXIDbCfcph0a90HxLDCYMUl56J/ghNv
Qgq9qQe7kKzYwRCbKL0j1lIqaUC2s5rDQ68B0jN8vaiqRomfnw7X0NeWI2EXVklh
EiUaUsM7u+aPLz3k9DGXf/hplwtDvJr9XgjcJexQCMP29+ZeYvwRyjxeQT6fgrMh
rozXRzEzSWGK9ugINiR9hhsFMT+VKodZLwAVX9BLCbe1aBDmI4vQG7svdecP48y7
LzrICZloazMA+OuQzQYv0m/k05RQx8z99XKd16OthkmNmYBj1iSxqHgfF5L+plqC
gDvYv3aMAAu/gGjTIKzaWRCLO561EAqu9hNxrRSM2r/eJjNcKp4ejZkS1NTD7oVN
tdQP8DwFi+aaRyFSSOVsKbcp1gZP1MWpQ1rXAVCEBqMnVBFRAaDTYK0+Ml7NmRfb
2jKwxkecFNTj0VfEO2EhVtlBlRmWSnaUZVXuZSDCzbNrjzf2LBksJ6XFx0j310Dc
qW51oMw4dbnSruXyRR0wN4dd+MrQ2iRwu9A1YbSzBAfOId2ou6bsIq7AIdZQSsyf
ZNte3f3pJk8SlaXqhHeA86N9A0H9j5dYRhf/qF+yluSV9AfBSwZWryV/C10BeEFO
MCkNkaq3DX9+FKwtpWSk68fXVd+ldtlsHtj0i8OI3c0eJ6JIUUXnnAFZyGNFOKXI
j33n9fbHjgYhXSOUaqGY/NyeeOUAA0m1pQQgkaZaPwvPRIxwiUlousRWmqXI8Hgn
Kuei7Z29xCeRG0TgOhGaJHfBkkQ94vjVW6sKhLRNge1bfDF1tUT9dhROqrBBhlUc
/lmMeTheW+dHYKs/CkCOV7diDJp1mKljE+R5KGKrXjlwrJycAgBPQGV1mAuuQpNC
gaBEEHB2CDQzzeKTbXiiydJFtNi/2AQZe2quR561JLgsrt7WE6UJwbHnsY3ZzcGM
5BAj9PTaFbNKPm68dWzyWhdlEXQFUKMuFcavOYWE71akd0EPhKUo51MEVC2S9KPH
l9DQdxyfDoU4ghXzB5YZjy5p9TURojdnF/pjENNmElg0W2EvbCjkXppf0mKMpcRJ
F2nrvaEqEbAT82izpmL/oAsrpD/wJrKG5TnUJ9yLU7h5rNFZ9e5huiJ7DNVGWYwF
j4bl0HlsHzZS3dUVN0HuPtxXVhgymfmnMYJghNUc8wD3xmeXS3/J9PaWt/pIfZqC
fvNgz4gg7ym3XEZo+JK0ZEyGOkv77AGYIpl0e5v6g/JlbioQwWeHzQRLcNsGc3Td
Jver8HfSMtyzGmotnV/DNENNiMcu/NJg6fBN4EXuzPzrnXfcTjn3NREg9PC/I7RS
3FB3yHKe2ROtUnY+Hd2RWgRhNM/f1fqb21+TBY/r0WDlcpelwgT3K7k3eunCy+1q
3E7aGS/3MdRb7/dVF0aWMMix35kyzaTgSjaMVPew/zjeJHhiP02+XJnpqtILvd3e
cXvOe0pDvqNbIIvPZHq8njTcisD6Oqz1OypC6SW4q7EKOlJQdK+HtumzDrx5UnxE
cvbqhvEsEMTDwZz6CHulLxu7dGPX8JfrzDkPzy51Qo7owF/MnWzY7vV9xtzFQDj7
YtLkpYidZ64UslLRYWPwdOiNBnFof5ptqoDERhKngPL63fB5PjvWr5qTnDSg2IIr
14PgeJEnSlDFYgn12Gv8uvmBxNKYYRZ6sXMO5/rm6Mdtx9x18CVfcZXKrhxNLfOD
jELwNEMTgME7WvcFteKojJ4JS6NHU/7QPGE+AdNm2yPEfbXrtWKyrhjZjDZOy9xa
AcSjA1lIYqT0Z/znlAUgd9by8+e+Cci1npNnedzRdFHzK0F+k9fx1yM6a2eG/U8T
PzFFCNHQuR7xtGljOB15a+YDN8VjFV0SUuYLqc4raIOjCgDL64acogEAwaNDZfX6
gtdEieOFW7IbKrAKnH18FDHv/frK19d6KTVBPkG++EpSovFoPzlPRPtbHu/Rv1N8
otjn4zFEOUt6oCDk7HbQsJ6VkslXDmiUs2CATrwxtCvoXhpD+lV4hjQ71I2rec3R
7lsZHIRt3SGc64XLCGIs2vqDRxNGf3FVAHDjS8FfegCuuw8RP4eVh7b4BKennCnJ
mClmjcB624J2qfG/JZ87gAibZ3lk8h4b9lC4Tx3p/u8CzYPlT18uP3etQ+uXl+XN
YbIxy+u5hWz6j9vwIlP/AN0MXD+Z0dXKqImGQY5s6H0/Qb1aYEdo1p7hIHZ9ZLdQ
`pragma protect end_protected
