// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:32 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rv1hFnGgmXGrXyMrpcYKyOHmQQA9oxl5Bnxj6U/P4YGe64EdefNaPMfc73Rxmomm
jCPRdBqOYNIRZXmvVOJ9UPs7sN8XKcQTfw/M/G7B4f04SG9IlCMzJutjKTg6hUJD
6fQkqPDRFiFDIQ3Hsv6Wbg2WVGvpZseoUy5MZ8uSf00=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8928)
7y+kChre7cTTYr0sLqB3GDPpQi0IWYbCxDhJ8rib+V2FeXtW1YjyscpMDKpQQ/5E
uM5RnSWcN6imMjTWKtLHNv7gk/RxeB7nZJS68u4lkgQs4uoGiRED2arVl6PFsk1R
c0MODWuLINA6XHTNeiU//1K24xdtE/SJz6C747yrohgJQ0mQw+aiCOS8rrge+Ydn
DSRRFd5FPQXIFUWow7jzJvFCiNYar07f8PcLoIbr7DYY+AJAfMVcOU9V6X0Pj54z
W/h1uMyq0Dw/AidLBUoDm1CB8kAJSSksGTVYS8I1O0+jhybpK0vR5AZ4bcA6Z184
jNMZDHdDgDCLDpRpUt42RZHiRM8xE8lxFGqovZ04JBCVOlgFibISDPmSHeM82dh5
tAa7IfjTmq/twNf/uHGwMPS+gyYDSMfOx8GExH7CeqlZPeGc1DrSUVJZoCkPWnUh
qBo9b3cD3cBDuBxK83jK8/UHKLsLZkgRhbGcXFTaqdC35TvvidIN1zW8uWKS0lOE
wI4nA7iotY3rxiTiU+4RHg+E35Qu/HTNVgqr4xWU2DI0kDN2YGsS1xPv8r2pKFez
1VJwFUGb23v/CNBbCInlTsDUBOxNlp+83ViIANHQpMGTI0rPQ18LfijSeY6c9R7+
01mbXYwrZybaPS5OSewFIUvi0D1B0ceSApMeQQ624Q4WrH7tD2HGZJ3usTNMWqoP
JMfhN3jI4TMWepYhDvBZJGUCRzuL7qeySaYEJF0F3o77yYga++S6g1JiK6ORsMJm
4bMFV9bBu9SsRC1sh6YPIGfLZfB5E9t0Ps+a2+btFgk8Sn0/bJfkntaIwP8fObwz
2G+/nG0uF816u8XtywWD+yudv8d7dvk0AuvR+aruYn6pbhHKULgmD1kAiX+H8Ziq
tSYSIGZGpAOHzzRSq3CZP3V8Ir1/AQBPj3FPNHrpe3VO/6C7lZWIgp/5wlYBfPdB
RaD+vcylX0lIiZ0MgXTCfFBwSM2kJ6X5awVlbXPTqclkAkgP/05LudnLAa/fzCop
Y2BvZ0cIt/EkAcQ4RZsreJjGWCa1tLHBQTSigDtYmx3EE6IV7LrovCCieWj0MoWS
sR01xJ6nsxI1fkoAsYDMW9cSjcBME1kryTqDoj706HaKANRBRBdSWdj4MjWDP3+z
2BZxR/w7ULkGj/HD6rZtniTJLJHFVIzy8agbXiczYRSE7X0ARctMzNBO/FHPkBE6
fcI0JDswUI3WUJ6hlaA+qqJEukoiW1r1l6SqjDNr+44TUnFNzB2j59ZRbFh2to6E
EOlXBurH1CRZPaOgh/Qfqj+lXiZKRMkLuzGKbRZnBquvr/2OHmQF3aXeAxyh5bQH
5QtmZ40/4uSL1vnHX5oubFGkSq5q60ZAJ4f7rZzZj1/7eqWAIdqiSyDFCtfDoVl/
d7mr/QTbqCVm/+vxntfrB0NUYvATLGzY6E0Q4Up4sgdmlnqkQCMmg82MghOn5E62
8gS2ovKCLUpvtLi+coyvHpg22vIFHCzkFjC1WfRgxHqCIaJAe2YrMVelznXrNcSA
CWuTa4mHykO+q1ONrTOAleGfegShhLkqVPEV8UfxJtOdt+8Kocco7LgPYQxIVKrj
7pYGjwzCDJOk43JGA18EiXf+rSoaQHnz/EKGiwAXSJ16fBbwzBxjn3j1acidXJXt
oKr3JXN4W9lX6OxQ3VMYASFQFbVlNfMcLqV3m/tk10MIbV/8EuGVLSBuRgyqqyxi
ja1WShYDB8St/lk/yxt3zE4shLa8dbNIynBBZNzvn4/z1cIDe9QZXdaP0uaenK+V
HofJhiNTOfpzsVracKAhSrLFvmnHgWlTlte142fVAD+ePNSd/OqENzdlcID/pBWT
HuDOz/Po0PfeMIMmiH8ub4zYc/nx0QnTFFmDO7jY3D4DKJo8msVlFoX9FDMmy1YA
g/1bvOSuxcvqSo3QB9cUSUD/sU6o/bP672VEQdaelZtEM4/SQLTELuKR+ZpXpE4/
kUVpniAf5cwXBcziya7Cgl98tiy9hVhKZampCKTDF+vgMqY1ZC4Iv7fI2tKBi2a/
0OfiALhYe0t2TyYWGAm7VVvJAkREXYFCz12aPCFUBRC7qwQ7gvP3yUUspjaUHJYB
BQrXUYnVfOGEoXgWLwe2FF7CXXvdEywbz0mLz/Oqc5QN5ItXW468s73KpEtnWgBF
FdCUa9A5hP+15M5lIHwyTcbDne1kwhBA3wdKb927+4ljOPnm4mw+l1fvVDAJIEZB
z+D86KmKYDGtk4OMLW7hCCt8WFuwO/Fsgr+mZFb7oykEQ6u2xEzWSSI83yVMLIAc
noZqmDlirc0dAhiguUJZ9lV6CyWkAjprmjFbDGmogMSzYTAbouFMzSsAGKeUgN/7
0lYnn3e2eQDnbIILNhCczhwIri5Mzhm7YKK1VmQu+/8yU6CU5/Fsmd3EphM8iYOL
543NBsdmlp1M7+S1CMf/elHqFLhH1BmS1g23nkMGqaoALVbCYDP5ifnii3pcGS4r
Qhbd3F52JacfHf7tAGOy2/sDPwCcPUULupxxvfyGfDGR0yMmz3gC4z2M9f3B/m6p
GTidH4lgbn28hHcLsKi8SRy8Whq6BGWW963V+ldlN1awkUuVT+nEFFS+fU6ACNNW
IcV6oqBUSdZEnAOmUIQikGk+1Vhtrb4hdSZSBueei6TPZ6ITH3H/PVFY3tFQvJYV
WAfEp80dSrKuCHpZbG7HFozd1QiEnnGLrJHrRaKLPCIweRh6dyQ17mWDIQ3/su9n
2x7seu4+eDs0afldR32X0eGUSdCEaZM9VkIs5H+skp5t6aDJD22AKP7jfmmEkwf4
wMQn8q8cMYXOa/ELo1D3xqtapkfjIMmIOskpcnom4ScwE2gKCgZvqCINNimUHEgr
xsZEqZVtPfgz+QFsnP7AtBHODc0tkjFjsyqedHI0u6fgX55D3xd//36ZNsDIoTsk
HmJsDtqQC/LAOsqXS4OG56KSqQZ+RFDF02aYwj2Uko/rRxBkoSGNdMlfCBRIdtg1
UheSfYaSrGAyhiiVhEBzRPR7y014XDmEiDEiHNg1yJOQVdjvMOhnzu4ZIXX430yf
d0T/TYHtLNnFYfPeuk5skaEd0V58Sz+G0RTy2WiBELDz1gFL5jCsMTJPGS5oSe+L
H+vurCVWgx90irR4ONyLgW/iQUUl+XBwI/Qq4FJK/D5hy2q4SONrUDdOj1/hc0K4
WO0clxSzCE6BfS0YMWZ09GMZF8Iw7tRUbokZKtCESDi4/KIHBJpOrXsihLN2w4w4
Aif/IGhSFPZRdqOwxnqB+h62s7wv7HT/U3yjdOakbKbfnDD2WULBh1tqwHFIMyJP
TGk8DgO8z/iCBMY1Lu3VL6xcJMw0OClh+HLC1de/GTOXWi+jBw9cjf7oysE+3CoR
qqrIyJZHANi14XSvxMQdJ6q9ND/Q0nHoj+a+1ADUVJXwuEJwGElAXI7nbuBq0HLu
m5PCSd9RtvVfENdGhFFFztX9dN8D2YkUm5qX+jSMRoY5AhB7hKJbfUylu3Uk7MFk
tSlkhhw6AgZPbpy7jFz2lvNJC3tHQSTuMtDeM1jTgUCs+PLBX9iJIZ9bi9yAlr78
gK6EZJwoALJorLfqpYOwuarZ3uj5Ex/dobdy77RHdjFmBWrI7ExR1hes2FlK9WVK
9XKZL6NXRnrP6oIXbyP3ZEw9pU+Ht6yyAH2HrEDPFIyX9bROataXWVG79W0a6rCj
l6UxjtSwhA+AHWMMxI5/342WTc4gvRtVIlk7WMomK4KXY8oEOgaFgAkaTtWWpi+/
TfVyv+FqkSDs1K0xuoJPa6MsfA20l+tm5PvSvg6njLyl0Zmb0h39Mpgo5aJ17xpM
1Au8tVE85UZ24poTcZfWH5nJNBvwGxI8t9758xHY+uKcmX9Tkfos0BThTtvH/B1C
YjxJn0SOODqARs5umgKp9L4ViJXij1JiJ0zDA9S3z9a+9SmdJXwrhDPVzSgy4pu9
vfxRf6/XBgmj1Oi6tC/7i4WiczfA2r01nxPWZj+6VcnKa1M7yHFLEy4BCs2+CB7I
PdDb4paDkYIfHket7p7VR/LOAwfgJGXOVj+leyq91ATb+3M8BXOfjGQww6Cy6Igf
3dkXh8mEinltwAECvLabF3BhcZmdP0HTbtu/2fmmtPt1XGN+ulz/SHnocVQOrHHm
2AcD7KyPjVSmbUS1VI+p02nTnK7fPsiF4Ly1q9EPOhd2ZJFsmctmzX6zagrtb5ei
hwR+AKb/CebixA31MyALc3hCjy+2fMoMGjpOTEzm+VZyTZlV+4gLzmG+GGRV37TY
fZvFLo4QbPJqGOX81/Cbrq5G9uJSLBEnQ6n1Nun6s3pQQClo0tTbjKbccWoj0Tpa
qUPj4Zjyp8QI6xpSQbw+uzUwIktvISDoCejGMXFKQOKIx1u7sBxwrqLzQhnMB4he
9egmwSfUtj+h+Ypd/Qmzy/S1o2zmUjzFdR19Bn9h45DvgBqqpX2MKSKIt3EET18n
EGS141H0lyEIcMZtmGI0pAkItbX6imzhiv8Y93Ny6TJcolywOxYELTLT2azP+Whr
YspTorv+cf2A6mtOHn90Vwm7F/kQs11/ZcShIPq7lJnOrKhMuE19XNMSOb9O490o
vjqKKrsDW90T/Gio1FCrL8yKWtMuhFT/UV1u0USHywYVZ9Dmy9Qb/8FNwL7UhkPv
kUNkaLFr1XumOKP9aHJfAeOnuS0PXclK9eyxG4/jZ9NDasbgpFjGrUYEJFUWV0ei
mZ377lzdb7VP+10aa5eAtVhWcg2lqkdhLvCDnkDCgXnqUR0+kvi7g1V7phBShJNs
EJBK5tzr9a0e5JNeEPnCEc0/NvbpdU/ftJhtzuSmNw39NfEC6/cjtV/lUiEzs3fU
1Zs6sYcZj54hb1cTGB6PxPT4jJrXPdSINvNCAm+8abUvdAZAa6qlqnLErp/bFoDm
hBT+Yxjjr4E0X3qjtfYslJh/0wbr2tHTJy+ywnkgmW/gtpBHu0LBkYJw+SzrX0uc
ZSACtaiPE5vSgRu8z9tsjYd1tnb08ME/QwPqNi3uWaYkfJT8zYZMbE1RGhSQff72
gjWREXlef947jG4zbk+PkNeyLryEKFSfoZaPWNb7dFkuQvHYoopgd+6Q97HOB445
OcMrrzExvFugeh0lleKmBKZqZp+yhwMHZigIjBDeGkoIuQPzztn4GOIeubZq0OJ6
17yFe74WGl1agz/4DdMSpzx8Ma8XKZRrDNM7iGIjFmqta15LP9TIWglbtUvB6zxt
G9x1hCror3FA0DHaKGlZtflZvW2M4LI2fKkYSjtq3tdaYxyFl1sBySaEOPpQHK2o
q51/H0Au0WxWKXdB2cXvm6WbXqhrVk9ATeh+1l7lFNjBmScCelNL6ZmIHmNtip7e
ceLtAp/7G4qG3v5ze/lpgWs3vawaNRn+D6/e5pAZHu2vOS4F/qkbMYMUsjfQIZdG
BoBt9iu+NrOyGnL1I9QA4QSpnkRo+FFGLF8vlS2H0nozELGtElV1zYE+gQ/XKAsH
Fa3etLxzp69AUe42tTjNKhlKOVjyTwWWDRY9AI7zMkqKSXCRjRNXIYIEdyHZfnsv
oyJJ511AQgwya+znlbnhSO+h8L/mzF16Yxjpi4zi78PsdTyf5oLQArO7pHoiUDxf
TZpJXxOlQITeQxzsyX1DvSR4x4lp7jy/x/VrxCC+EHt912VEhNYKYJcVodR6X1Gg
D+Ipnh4gNI80OeafN9DVNeBLP1P4AWCDjT+CI5helBNoZV9uQ9ijWkhw2KR9TAQj
+WXWTK5EKANEL53ZvP9I7NseKpKoOMtzRlpZx86gjs5SFsrILUOr7P8Hore9ZqLf
KORNc4FmlSC+9sCh6ZR6CExFAmNQIENJ7QDwuCxd2Lz/8xzD55VPczBPkl4HrXZ5
ZGQzgLRTlj+wh0sMFLvnHSd6utJ9Fram0EfLNbR88p9Xg8Kq2cwWFnLzgXiO5y6N
f93xBSdMNwPt38WuxbYKyRQrw2z/iyTNREsordcvPL9famj+64W61ABn/sgeFKWV
Iw5KY4EmepcvNCKGiDHrozQfoLRzEoQZjXd+Pqy7KFMr9H/jtaGqFqMT9jR89Nca
fQKTtGwO+WYGkRgLHK8CNHpzWb8NF2MeQfh1+QMtoKsJ95dVxS0AVjTATx8LNNJ8
k1wzEXv05to/zxQxoVkSiVZW/tFI2xxUWaKdiaMkTEAvjdE3jH+3C/BNW2SO9Zo2
ONec/IdJu86zdwl7IEaKYBjO2rMF3fUpd8FdqbrefKK4MdTC/jJ43olD8j6aJiJz
aPTxjjoQY2ehxTMIIr4U4l8sMOQGOM1jLxI2YfOqG9Ani9D3xNMec7UmD3a6Q/Nw
T8Peo05mKcbCycbs1m2couFHEYAFjnSyD4+WtOb8iE0KG11Z7FvD6HjvCk/G10P2
a71RqRvxYfYwgY6d9XbsD/le3wjlMKiRJQL2peceEFaaFAoGCvSfHwGVvLi4Zzjq
qi/HCoi0mj5/CarOfI+BaWOpOdvK8tNPe6QqdL2lUGtf/6id+ucN5VcTAHtOzsYS
9d61R1JnR3wRfvWvp78YI9Wrksj0WUYFwoX3mMidF4NOV0+1GFouBOBbn3asoVIf
X+pOZuxr6FAyEnm3rWnv+oaYNYiEbiAkfESLJ/z67URy8md4ohCZ+42pX5/uDCp/
qhkCey0eAKgM4KdoGNvaC81+l5jwPr1OqoCLE1GxJEzW+VBocpT/B5e1+y71LN9+
0ZZ28WqPyBqbohV0EormDqBH0Ptawzj+AcVNZtDglRhNbCPouZ8noKD/Dfiz/BzV
KtdujBx9Gg71EQJjNTj+B0aL5Lm91RsrSVIqQWdcIO/GectaZR60+BD9eyTwHbkF
JsS1+yPvTfS3G6ZuoQPssFTS3bOj+Lpu3hgL+V9pEHotqdHHbj08c5YbcIESapMo
0HHYbcT4dgz/MqC25qVCkB5PNAXcm48Mf6xN89TtKs3KWGDnaY0VFVuZJZ5l/ZZk
AS4PRQacFbUWN3yAY+6Ewc+3AXsJdoKVYhJnQ0XmMhXRj1+r0+iI8IvCiyLtKYet
AUFHJrCvX2mq60Mpna2ZDcH/6rsKHS0zaFI3xaFEBketIwq+Owdia4gJ6AED3dMn
1qNrdt6ojfJ/hvv/iQAG01zYQYUEKioGD1RisqfLibU0uDgO32aWZYJDjIFC4Spd
DQOXI4Av+1g3yI1RalxfCgvlv//8cYusgRq90ugC752tsfrQLzpEND1dVdMwj/zP
QOiD0rSeRpDReoA1EEGs1tEvsQnctvVyKLVMTvYfOVaS0peE6BUITh4CZ6rW5yq3
5yoyzQSN9TB8/y9pYxG3R5bev2rxGbKQrmLgVW5sIPX79PXfbQi4cosQv4PTSzmI
84eK8pS9Qkr78PttzudfsJtg0UXkP7c45iApOi05/bLDJFOQjT5/dQvfY2QkF2AU
9mFHb+Mdn8vvD07H+HjjB9w9i3gtMD83yOTUxV2KL+cNud+CHqllibOJZNFgYFd4
mGSMGt26bgVBjgMRGKJgoYobTFDrgMcWaNRrG6XFCi2fiqy8mId1sf3YB5VyX4WK
OaHjzmUstAGIMgRS0xYeLg0sFjaz0d/Gc2q0Ham0p1OBrpx4t0mf0Y6Rw/Qs7yni
XjJRcQrujQ9eVFtbGqamzc2PBvK632xKy0bKKY/GW3dEM+YZBfWF3s4cV5W11NPS
eyBZoY72buAv60mOr4g7IX5rHfAkuGJWSPJkv3hBNFt8c8spOokpz6C6J98q8vxn
zoMSy7ptjGXGJATLyquxr+/9U/rmEAimlx05F3QAv2jTJm2wkY0r7KP20msWMD6j
V4YAhQVFZjmo2d581ixiADvyNXFLyqlfTCqdykAcZhhtrYMP3Pi3QAN9U2MMOIVV
ipFXNkyTPCXu1oSBkK1/+2Njzd7SJoI65ZITSJtdYobvuhhovgfDcqsJRw1c7CY3
tG3uGqITIrlhLXSMAh6/AS5Q8bQtJM26FoK0JvUAMBtMQsbkxjRWcINu/qgxjsRh
uoN/11RzBv1wRrvEAmKzq7H82dcTvuiuE9vuISD3Rp1TLWWXo+xy89qDTzIfUSqm
2FPA0rwslffp/R4APAzSnL2i1xMKp+VbOrFpS4uKlrR0wqVQovO0vhLoySeKlmgr
Mwqrk6pOSxlUE5lH+h4wRvLNdoFVdfqxef4pGha7sqJt859LMqLA2xmTqeFQblVa
8PFfHs9q9QWPRtKlYw5N1IRP9bfLMVZ/2yKpoHNnpvXcAf5okl6dC1WNNozJp77R
g9jqcv5FBM/I91RgwSd/9QbD5JGJ48TEq6pWHKlSI4z717mNh0GnYCChjTBR1hxc
yE6Sm483Bgmb4Nyy27ga4cWMcS5UJ8Z0/0G3OLph2YXX7Q30sH+Dy4D3D92h09hi
SFHKk3ZfrH/W0LgAFxXWH7yyFJDi16Q/85swXS8pVSDGTnY9M2SzL18nmV77R4/e
yB+kZvJBNqrHsOEFIMjY9i8q4oDPL5RFPLtBgfQR5Af/o6WXyStlVmEC2GV5jK9a
2p8vSo54bnIC0lFm2fM5MFEt4YxbS8FVkljAOptO1KEDZ5ZFQfRCMRmRp6j9frrJ
ko7o1t30V/chIvx+IYV8PtQI9jg8WjB5st1Uzko2NyUo7tuSqb1Zat1tt+8srt1m
64Wl597cqXwOM7nQHm4YjrbVYC4BgXM9qyEWi6yUbFr6R6M5lo4IAbUSk0Sje2jZ
bsqeZ2PDycVCHZaZKht3/jbSRLUZyY68OswTEkUvxd0JQwhen00a+unSXrwAYjSl
GmilwCVvlInH5tTfGT/6gAMxDKF4aCeLP0RD/eZNp3zHNFjXS83ER3TGTIfIGzg+
qOvVHz83zyRaYIgOwB1PO82t6vIbZjF/yogwFL75sSzOYGySnWz9iiHZaQfD9Bu1
A9Q65sUStyMtgVF7fSHdgm7okG3zCRoSS/wRpYZs3OHc17Ccqj6+god88YS7CvJ+
mwHwyvgMBDWy2B3LFDYq/2Qpx5N0OI7Kh+W5+Y+W+sntRPkdSKN9Q4tLnuLUDBO4
cAsUt055ZVPUSsk+I3txndSZl9U8jv7J2jnfWhaLD8WosRLJvHV13WBIwnPK7q3z
shqpNXXUjXkyi1kB7a0R5x7nd4gXjmTgTYCiSnltl3AhzQVejmlidiRwa7GIVAq0
8DiR8ncnZgm2dEa1gVXrp9pol0UijjkbdkuWGBTBbnpxx28ueuTrnffIaTm4doXd
I53QyXjbsK3ZBnUXVxaXzBaowP+Hq8xedDos0UuAPwtLQue5+w2XIMtc4GghUlVS
82AuBn6c4mT0CUMhVy4OwH0E30xkZ5mEvhPDjEZT66ri2WFusKpC0FAf/19M8bye
BcXIbh/fQKUcdkJxPo0nhg5tkusflzfg/sLJN1DrEG+SJ7iCAFR6eUX/V1153wAJ
aQVonK1Mj1JZcrxkE4I33UeKOlCmPMvJr1n6BLb9IaZHDN0VDc+OGMsiYk0rEeG/
JjQYOhBFOh13SNUBsmJt8YKWuzfHBV+62qM2ZBuPRqziTFLd2YsHo2FlRSt1p2mW
WzXZLsEbAjh5Hafp5pb6IlxVNR4IeBh9AnBAGTTWK9RnQ/sofkS2JjJMspFW5AYC
mgC2IyaICDncdpAHfclvaVb24MbMC+WmjoRPmk7gha2A0MPxeJkeVsdqFEEWAeJk
TUXvQY2kuB17ZQclRIFAJqVa7fBVXsZs30UEFMIro7WSj07ioxDjZ9o+tfijUXqb
y6LVs9zfzsEqEjayzI5QPfbnEIMutgZJOLeh2jAgWVzoyeC5J5mXfnLGy4awp7Wm
DQ2tsC/5IoIZsWSvPFLrVrxhH3Mpl+y9r7eBpxpifNQF/XdwATkMX0Kr/Z1hnYSS
FJEjMQ3CSZ6HMWp/gaaIroJQT9LNgLCmNNTbrB8RzyDh5koWwy+69Xg784ysQtpR
9PJBqxySfhfju36DCQzt8VkMlf8/iegqkONlErdYBySFs+QYzCqfIpR3XGM41lvr
ybQsok0G1KzvmFdAkOBqZbU6MFieOAZSXts2IdkbbLUseOy4WiSO2yTQEys2xPii
ALgR2eDZh6OU53ChvXyYazjRfIR3Ae72zKNXs2zFW26OD0QMWGQoqLKR5kzEW+HA
3tTmuY4AQ1vBllOaHPFRu7DdEbMoEHDoUK886fraeg57kB23h7ijygei969jMBbF
pS8oaePpWI0BZfmrG8SObqy4MaaqraLImVcumw/Yw3ReiU6XXgCrFvVyf8YWJ9Zv
kdvZ1MQpU7R8XdQ5XvJO0jO/779mL3PnErDNPgYZj65TWHZ9QaTYHIEmt2TkrHLr
wPgYfIPJghKwzVMHh2Zi7PAcftNCVgBaBaZK3NIcA36DTReLujYmwmcZArBiDRPI
MFnKRX9eumeOy6XjX7eqHbqJ/Zf9bJ/AmLRxyfchHCg8m7LBiR0Ht8klEOzV77ax
5FaIniGawescFIVVlSjDYaEQ6ovDd6eluFID0eUKlKsB79O1/ToO1NFn/v8JBkOF
fn1AtZsn5PNSlGj61B90Olfgfg3z8lasOS+/odc7ZXfTNuNfC7MDLF8dSrz0WuYf
rv4BfuM/q4g80i3ixXl1Lmwnyh+YrZ5banIGqG50dMvK5IWAbEKDYhH2gyBbwlnb
Blj6Qt4/HZjFRaD6Orxa/LSUWpa4hWhcWch2dUdyt34Hdtoyv9oJXhHN83DYVyib
N4K2M/fFLl/4CuPJAm6f6O7jNiY5LYWjpDo0aG7l2rAu/nZvrMCUVGIHrdOnP9OE
CoosMzWuN/GfH9d8wf5lEntwaEj7xQaYEmqouJoWhLHUq7n7vdQ3zHqgO3NDtpBe
b5oVLBIvzrdOdDXMAZHTKrlQy8Sg8pvoyPcXw1YLnrRUbbr4Nk3W46bcIVyuzBTi
/cimhKyq1jg6Y0Rj5HNkEW64r/vvCTnjYBl0A4vR5vr4PGDYP0o9Oj9yjTUF9JPB
MW0ytV/IRKNsW482ouKItX4GdFws73iqxaPhJ50KeAIqaDJhWDG65zCI3oHWl7t0
w4ORqWlh4bMygQzA9dXvf9mDoTYLDH7hzX2pMBnkr42W+ucYYAhi0KxPdyqHzCLw
PffgL1Q38AvTlRYwrNUpaONVwuTqQaERB9BLGRj2BRA2Yr5rH0lz7DGaCspmPsHj
+37rWdwfD3OFH+sqBhUO3dmY6XeFr+ZNqAzwLHGdMtadMPx+GfGdw0P/t5d9q5a1
S/X/8n+NxnnDJY/g6mVpoOti8k1iiWKFKYNQ7ipSalziS5dN3DWNaGm8Wp5wuMQB
GIiE/E68NHYqKmXHZOr+0B53V5CO+x+XEXuZK0FaJD104XtoeXV2Ub1quZnNIBDX
EK1yTlUMoudMVrCrD6CosKyY2RdEhxgNQJ1SQR992RWDUy56f1O8A/bps+0npfa1
cdwJ6AOpbLZ/l7qBIqhevofMSOh8jCTlk1MhboWkIFywc2ccxTH0ba8f9bJn6qV6
QAKzfLyv6SSH+IXJ1YimF7d8Owe+YSMNWlGZtLo1z6Y1NA6ATFZmdtA7XMoq8drY
+BasY0/20e42ivKMtX51CtCvOhhC9iKwg9EroFadHwpj2nSiM+vRdj4lAGWrkegp
jnQVGGpS7vy74bolDqf2FUFRDaS72HGzKft9YwsQrEJZRbpOjyLjVtvMU41tQ1r7
w3BHiDC/xLCyjuJaNWjeWt4TEvbl0f0mf7ZPyV2EdiuVMDPUY4jc9bXpC2KHc0nl
h/AWvDQ6bJFJpd6cPVUGt1kz/9qiUSPIMB5PfE1+CCB02oMCHmRUs7uRMDKGNhyp
spMZYLqnKGvS3x5oJH4C4N4uqkPn+YJaBitm7/l/eMYB2BooSW+VWRcBrX9z0MbF
+nZQzCKaEfZLJwOprdkyA5S2fiPlQLxe2rX700swCbG8suTpGohXAR7uc61IPKkW
`pragma protect end_protected
