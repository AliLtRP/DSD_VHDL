// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hFAOOPoWtgfnPEFhfKoZSNre4FOlxqgxp29/tLHhCm94cEqEoPFGN+OLW1wVUvrQ
n2/o8FuUax/7NMMu5RrDgm2durfuRrAalMhb1yHi0IwCZGkY+MJIPnOzXpPEVEKC
BA5HgpnT3KJnJPeQVJFfbNrLJ6mpzz0lrQDtthWavCg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8624)
z1EWXVgvSbJmI5RLXQFL0tfZ1Xn74MYGzK+XPLnKezq2a9b4hWDWbGY/JDvxQxld
uDK3DBcvCHXdKMeM+/zpejjJhnjrpZmZaRC7edAHFmlG3eNqwAPiWQSqzB33TbrK
1Ia6FtaE3CbrGcoAa502FzuMtyDPH6xsAJZRkTM8qu33dAwJpSIZyzX5nZE6o0eH
cAzzkCyt9oDETIBHikO5k0VU2yX3mIAb6jhjWV8B7mCcjEv3KeEu5S5/3qLAT6Rm
Xs/7mI75JQbanzgCfgLo7K4K3g82WyUC55dDj3Ha+0HSPV8Ga823IuC7/GkIbqP5
xRFSdJaQiasZxpSfmM+y4loXu9e2KhF5UTWiWs1CIka0Wg/o2aAjMtEKZIuImz3Z
iAjXM4M8dEJBa55kQRT/Vy89XAnEm8L46rpqdfR1lz2um/hw0t5M6GAom4aGLF1l
NTAAGGK/qVpHH5yl7sNIVgcsFLJSw5CT7xfzst8oV+hH5FTDU5np/YNHVWPK0qRW
PaJl3lcvtBl35Ftif5Nry0nd8ECPW0sITIufFpTuI9JPoyNUCT3nluoTFAU/vtLx
umlR82szxLZLt5S/l/KkdR/IvJ4S1KSteoS0++Cx/SrGW7fqhKBolMHOPcgoefr7
Vp+Q2e5ZrZSBRKkVfjin4JjHv2U6EWcKumYtjWzlxkd/3qbuOYBJRW1D9msqwzHD
ZlQuuJnPdo1MNA44+CiFz5vBjc8VZpjocZgFvT5Yy25aMBko7vPzGcdn0rWuf+HW
O93no5v+5G0yt6ICRzt9/yzaUORVGGPssrINee/k9Vjoxx9wY/x3MLpHW3REY5M2
+LMnd3mz/QqD3lJcXoiyapv3i4dpLwI+3OF0hc4N8N9t8u3al7SemhyoNt4jlT0Y
6+qw4GAOWYO6BCxp4t2u5JObfSuz9wEwVJYeySRJ/ErVv9hQRUP7CC0Hr/Df60bN
5ry1u37M+9a8bbG8Q5oNQFykg3pcEx2beb6FuHheBlb85UfyR9WD0+36KgS3LMBE
n2y6mXJATwmnokt2wCT/naYYywRVGrX53qMvX7HH06yXCKHCXGVJXaxFbkM5jI39
9HE2oLQXEB+72zUWNupYXF30wBxemHJS/h/im/oBT2NOdfSVSwmo6Keh949tKZWl
QiBzkwcaiZo2Ctn0l7V+43U8yBW98nhgp4MfvgrjYzxpzru/ngzDwm/gKaBnOHjB
p/lqfZU50fd7QJLhUmfPnkbvjXb7VkmIC18+NMX4wYX/wysMbhCG8+SnC2/fl05m
dffl4ajra6h34a2+Evqs5OuE055Tn90DI1n7fmpopMt07pxJYv1Y8pL6CmUDKsox
SGq3+/da4+cmv75xo2ePdhV089qVVypVXWpGj8j/2aj26WisRptQcM80wpK8sY3z
GKZJS9hd0stqsagIkQPKuvVZsykqJL+MveHBXKio8uJ3tFrqpeqnbLggdoRWFlTQ
nT6ypTGmsKiD2mpjMt6qrYnWQLkswZEl9i1RuE+l4C97SZJwhtGgEeS300gE0+Fs
6Ze+j9djGiYx9ZPbPp9co+td0hFdfsVbcg6X0xToxsP2/TFoZ9VGCKfJYEak6XUY
1US9pt5dMc8kQEeAF5XREwcacemHaAO70/JJETP3kFNJ1/kqQ2DSD41DJUBVs+M3
2gqQ4f+DeO8dmuF43DdCzF1Km/lHoKsnxJQtObcR3bP7AB/c2sBiLQYmKnCTS/oa
H4WPWXumYCUS6tsbrbyykbh2POCz1hw/NWB2Hr7W8jCCVNui3UpwGWbj+V21XKjd
JlC3Ukxu39jCVHwNZN/1y/rZvLGNFMwlCYav1O4ymfu+8zTDRQQ21YN0PyFRaC2u
lMV4hpZ1cak47oLEbfVUn+4HGehZT1pyZcQuFoME/kGgI4Y4svSpv/242Zlgb6s+
Yr5ymYJUyeJ1bkv9jLEuihPtYtOxfx28826734Np3fKmnYD1wvIPuvCPGjpJy2p5
ud/RE5xMAggkplzTHhzdxAeXBcDv50Cr9WHdvfnhdpyM/L2qc0ckm32NKERm3tXB
yzEdIAMuFQ9KGebN7KaPRPwhtDLRG0z4WSJOCF8nlx2EaD4ZmX0a9yREg8no0mDS
3Y6p9NGsk3VatMMseFJmHXDqIhAsn1QDPhZfWozAniQtGNts82Rc72c65cHgahcA
rKUoXbMKV7/0ku27HakVZCvZ6T5Zk3RKfc5gCWdRgWRykjKUKSqcP5uTNQUJvOFQ
KIubVXjnhEn3yntkjs7RpgnsRCiI5ksDxiGmhesHMlMSSL/NEyVTq7mPtrC90spR
Ag6ZtyrJOOG0cepkOKBkpxxutTJWpm0prFrcp/KiryhB8GDJS295kd3ev1oHrofK
MSX2ECa2MiqyTVc8Aath/G0/9ES+4laJy2pYB0KsFTsXUfzFbDohiLe/lHRGXC4D
yJLhqMR3IwxX+V7cMNk+wohFTmMYeVT4FfV5IhzJBY4fnMLMFGHDhbVJMrQg8qBf
a0EcK6Glw04kuDA6Pyu/PVHUBX2ccsv7eeHECGJOIS4Nh/3iCuejHS5FH0KTnKZV
NgPOi9SPg5Hq59aw/v79eT6gNmMmI4wMfhiLnbKF878QoRKWRezoP4E0ZpkYeIXb
hpwimDUkB5wPJGVsZEP+J5d9VLp8OLXneWbMo2ysgsq0Bc4M62k9F0hxJysoptli
6xOmArcQzdHKgRBOlI16Y/J/sp8x1OPrZQcndwhCnby1C6cLCAYo3ST1cLzOeCcW
JXAM0r3R+EU0FxRd8hrjSPK3MN5nTLHhVGRMQvwejLoza/5LG0puF03kEDl/p10y
3vOFKuSIsE+0QnaFpLCdQUxEdjklbRKX9go/htUAlf8OiNihV9gGSEwFKMOl5TkV
rbmgXnBwZTiHjjgCuFqUZsdcpkpryVkAxDrSRifIDI27FPoHy8O7ugDcehVgrv77
PTDsoqnAT3nZcBQ27iLhOOrg38r++SbVvgta2P9xsvtbGvmG5fDFbUgei2iOirdD
p4onsVgnPZBgxgmv7MVGAWmH1tCBaKYGQP+rF1Jjcgi3B6QL9lfTBssm2hnIPjDd
FjUe+68RGJZVwp73Nlpz7rcERmkFH2j0ZJpAEhZaYI4kCLd1kCnfRq7hES3kyhw0
9alQHcvgCHMjKlUyphvJqtkK2UJTfh14GlNSYjtOP/LO7Timu5cJKooIE5u9ZHH6
9FxgRkU7sTgcbzmwtQDzCLC/4rpx0sUdgg8jPvXqPQ8/dDa3uYlARm76hyE5kCoT
woxOYABTyyxTkp8NnIWjgTdfuCSpggnQBMfz349gdKgKKlNZGYmP3ZB8cgvEs2AB
6o7jeHp+mrvVXWX7biNcoWJHkmnkIThNzlaIsEbN9Sqr65kpECUNNtLarOi0GqAk
afWzEs88D86etI4iCUk/yLGq5DOHGYTfChiGhqzc1CSBmTdXx4krcN1SVJsJyB2q
JsL0g6XpZLkX2aVtAU4t7wrtaaW9FTPqHy0njk2u9TbhhZO4AVU8k93arb2UAnKt
MhAqajn1QpaY1GDl+g9BpLY2MBuV22osbOen5/OrO6GXf8LgvmnvqzKl2xCyxS6u
vRK9AFQXtirZmw1/42kX7ew2fSpg7tIZxyt5ifp/Fy1t7tG89Y844j7tLERb+x8m
TEJcL/G9D2KwP9sAZlUSWBffkQAgGL8j+uo7FzSVWQgAyKObhHBdg9BdLd3Gg5kp
XKyLDI8VbWhSHY7J0ikshkVC18MUYzBweic8jRpnZeBR40Hl6rwtNK0sTFeNOBlM
E8ljs/sqbk3JUWnZKCk7kpjFBxyKBPvMJ5z4cwn4YP181lPz6/9r1HDOHJ6LA5O/
e8S6EjiBLAHgNCJMurQn1fj7Cgqh960WsTGKMna40aEqu+oLwjwNxMTwdzxJQX/R
Np8gynVZOgiMwY6DKEmJtLxZGnkTwubNRcHvVEpx8PxGw+yitWErYLUei1vagv55
ndLqeXzSfCOmjVWYegutslx1Z+raj9oYWCJTUw5XpEzhA7oBKS/BsQbR8yq3EO3m
OKrCWDEMD3d1MBFRdY2QgtGIIioXJhs281nCHfZFjXsoYldn38akdibaPcSDX8Xy
ZO7HFxRPsc5YGXzYAuMcFC+iSfNi3RKiiv7Jlv1X832XvY1n8DG/doXmLMvpa2+C
ndNZonGpYCkX/1xCjBaKGPSsLKnHq/UY5prmdJwHBLtY1P/DJjE25hT6Rc3RR2mW
5QGYz0Qbg630aQl5E4PJwjQQhQA566uyhYygOWK8LHJcxJK1GMbmY0Vw5qJEvvHz
ti1MUssNVsnexLw9QG6SCPG+EMx8f/HgFtoMMaFphod6y0dzZV/tPz9mq7u7EA2D
ZVTTo81OfzpmYQHxCO5+F9DZU4fXzDkHiAxQWnV50GkU+bCjtHJ1asL2DJUARuDX
vL2dd4RRq8lqP+K/wgYObSsGtlOnvJfi0x8OlfSy7koRXQ+JJl78QSEdzU52KShR
rZ8TaRhl86wEQN6Mz7m++wfn0xTK2Et4DGrYEZsm093egQq34J0de2HYJlfCRdoL
z/KzeXHVMlsoC0NrAg9mH6QkArqwtM7ZmYZA9iKwNZ0/rZiAb9WcorSvIDd3dpR+
ETK+ieTzTy8f/J/vuqDGdXk9XaX+am8d+OeaEUkBSTg6bwUOe0rvxmcnSqnv6VvU
TJgAKGV2FBmCl4nDQ3NWZqTxKOYbThg48f2nRfremgzD1L2RkhE+TS6ts2RXkGU+
qv/x6w/hRGYwB0xPT1Jea8owyPFA7OGo6oM29R4QkO+YkJOQh0McELvySyiWKYRz
uNR8TdHTPsgIDF2ZFZEXoQuHYWOi30MGWN3HoE7SJTWZVZ9rsLiK7V+uXXRePeE0
96l2UPGrVpHYCJjWkEZyF4nYTf4QNqHcckjvDfc//W/S7Q77rwpqrRUk4HmlUU58
7H35VNIc56mQfzIV9M8kuNPJ8C+sGmRLtkmEFjQx2eGUGyqzdF9huN3S4OcKgzhI
1phnD7AZ+T2U4OCMiQTW62Vhw8Y+E+/flDoTP9r1YppvYWaqRJWrOOZhGM/bHtto
oxPFi9bvpIw/5NkLC60oc0rvXlZ/hDNo16yedw42mXqMXChzqGwPyGmoeQn0UbZD
NXFFyJos5CwtWyj0znve/RDonozrFa6d1eurr31cUfD9uJcvxNOTV1w7gY1C5U6n
SYY4YmpsIb0tOWdYTbyfirTYYJUK308Vx6BRvfMvKS5FwOQDQGkCnzQoVvrlEt1v
lvYr6y2b9YwuG2gMvG0Jtl8Xdakje4/yRA/+TOG6ZP+QVuYb0QhPMz83LIvMVbyH
QoR145LYIwsk+WE1MrxCJkhbwQx0JgPPeyYG87rNsYrmfw0L7NpLclEVIcYxvDzF
9mEAaDwiZIKHe574WmhKENC/5khl9q9sWGbauO5xEhGqr8nNMVnoa7IdmtAeh1HL
8PoXioam0/XgryKJbfCqfhgj+KfaeJONNo+bbN4ZgpfVWKYM96awM4GxWWAa9l83
h2iR3LDomS+rdiMSSi9sbltnRoZHZmGebXzZdhGoXQYT4EEt7c+VvE2KsjCHVBud
IVDTTzsqviKOUPI5NiC9KhKkJl9PGFY+myVhNmhPQ7/MfEnvGQ1aleSLOaIxHy/K
B8XxgoGo4wb1+mZsf7PB8ADnZ3kVCteR+45jTJaY1ILX8XRGZ2OXdK8UyLVdK5LE
qUD/KQkOfGxKezKfGcXTvV9oMgh+1Qn5jtMjer7rRcBWpxz/hvYejKQlm4mSQbhi
glLpDbR54CckUympXmHTtJ6KJ3MZK52tPJxti64aLk8AtzTM8cOn0mrXv1Fa6AsS
v+1Nea5x6HcNUDHLrQS7nvSAwwQp5WYCevoMEZb9ecYbEF/Pu7rEb19givEsbz+N
fLNLkzH9NIBwfBtiYVaKCojnJuWpDeyZktf5INqhm+hJMBB6gNrhkzemzx0VLakk
B2ka5kCDNrvT8oNObhdQzQwpvKgJ2S+yN+BjsCpy0EcJGYiHNvNHdvJ13bBoYiGf
bNK63v5WSBgf6j21kGGE6vqmQcgDPvV07bCmdZvz6qbfaa0Il6BWqS32qzsg3l2j
kFY5rcySZkx36rI+ulAJ7ISHXhUN3Ye8qhn0b4cbAUuWOMuw9RZtEfbvMDU1E42C
1zOK3yJa/fO5ImMa88kMN8fX7KWAYwKzAfCPa1Y6Z4uZ9ytlyPla612EOL4sQWhQ
hMXsUn8cY2D8AXPTVTfKRaVZatj3ubuBplj2RwB8Wpyu+jo404zo5rCdmFVz4tYX
RfG6p7CuAVavR8k8X5pYkWmzCZ2eWVLFrKChJS9DGfPuElZUI1VM1NByXzjRaNTx
T96Zrj4rfmKjRaElEZ/J0G8uJ3yV0pRw7VtdSzYPYMiBdXqPgAzO3L7DYB78l+LR
ZmCmwlMtaqhdL/f4UHOdvaBVV+5c0NmLd/eGa0wJiJgiSMzN+e9+FskOwC2KoXpn
P8hZiOTHejy7/SW+T4k/tb8eHMfu8AtN7tN/e6ym76PlhRC9ZiLr/MA7uC0nNOTt
IKLR/RlxADZexHEwS7RCwLgO3aaSHbG+KZvsYQbD37iydVng1fVQWYekriSVyLwo
9pPGDBNowmsLjFQONPKhPowaViRl1+sIfGrs92/Gq2YQjsOUcNGYpvDCO34iaqyT
gDPmczYoKnr+vI7jrR9YIzFUGWBmCKy9bkzynWQT0KX5E4DLPANqG2wqwGBmDOxm
jXg39Rfmzq53NJit/vbAQgFZP90TuH3h+PKvemehqu/d+vgJ1TUOtk4LVOOJa+UZ
X6BPYnuBnE8znvDZEFj3FnBNp39fhZaLvKnLoowXesyoMgRgdUOjbdpM3QYEx9IM
/hZWC3TWyTGM9+z6XSbyUeyCKx7qzqNF/KYWrCQI/i7oWT4iFH4wgl5ucSMkvlRy
z32Wg6D4jv0X46PYeJMH3JhwupVApdsrZMvKqQJz/qkIN9n5gs2RqJKGVJ3SP7wa
WHmT1bPEVkEXsaQOcLYPSd2BBdYn5JVoyq2ZcZjkas9zpEmw/2vBQSvYEk1rMsSo
22z9naa+wzOo24MgsPOfcQslNMZDcwkMN3lMln36wnxFgeIm3Q0r7M5T7CtJGeJ0
gUzsyy0eRSfT49qb9azAyDQ3FSSNHn5/r+UVVim3O1pFeJLi+nk81TvJE0S+DbMg
bmL5eMssJQbwcIiYoPSKBk1xhpf+g4WWj+rxl37YN74wtA4rtlLdYEIgYm/HE/K9
BSeYmW4Wc3sdFOWpccPbiUTLFb5Fhlc7Ylv4lMc/KRUcZ23QwLYIMHSOd/fFHIUP
H28kjFDLL/JkLuxM+ohuTX/RsRpNylbUy0NFmCLc4BlDHz6vHuQlf0GF6sWVe7Lo
VRWaDmYRS+GHKIG8ALPIQwG7N4VeWXI0DY6dJG7uMqYBV/2mQJ6jQam9ZTktl+xL
RnaRbKcAN+WlrAxLw6ZSs7oX8ghmMOJR2lKT2tK6boBF38SK+qmmifNJtBQ6WEWf
U7Zw4774gIxWdErGt238UiLXDKiaAXYKuflz9K3dleIlEMu0pi/Z/ypskDLg7e3V
JB9Ft143l6UyzqhlFPZyCpG+PFPiqBN6W6JEMxkpkiasyVqflsDMzbdLq7rcwAak
q3vx0jYVCkUPpDjZgOWszCxMB4bI/7+MIZywG5fzgVoIQATYtyxFWWKGskwGK7yk
HzfmtR7REpAd5PmysetS5Ed6tWbjAYqkFNQdQTdCHD6vbzNySKMDr4pTjhCMqEJ8
BIBZjZk2sPNzxiU7zPT8mOSVVS2X932BRVzHPbJkT4Yuv+l1TQtqjaVRKvay+z1k
pfriFddLisobMse5gKeTYac8arYHCEoWAeVFau9GUa2gAKPJNShyY8LlFyWwuDUC
sCksT9ZjSdzZRTwk91Dh3ZBoKsAOQXLIezmkTE3vE5qp4qASB902slKSu2lcagEr
MvHhPAek4BroF5xSb7JQ3pfHh5ND+qscsCZ92ItEf5t2qMQAxXToCMlWvJlGOHtd
ysCmE6rpu2dvJCGGud0BG/pU5SQaP3NdAeqLCbyz5yLZJp+nbd+laVMFYbMVE72Q
Udo98XSGJmf2VdL4JwCXXD9YK7BjNaGOjiS/VvR9RHlpY/adU3pg8Y7fU6AXNN3j
NaIJ64L7OVNQmkmHuePTngM6GsTeLxUkoqbVrpOLznRbkea6kC+yr03eKh4iju5Q
BITunNRk59/5EwuBik5g7kOzTYobCY2pFbUAa/GTv5z+p4tZ+Hka0SC08XyfMhw5
PiaUoLLGbuoY2fiwe//O1iuVS/yQ0PUTkdE5B9RddLyEXLsbulp/mSUxHJt+xeib
VY88YnsBEQ+fpf5vcO4k327/3CElFt08O3Z6NWGotKf2KibaToYw7HYbfUTsn9oY
rbw55di2BZr/NVYB9vbbOhJT2vvoF+cmM6J9RgJ3yu2UIOFZ+LZH/Wa7xutAy9TC
HF54vh8vcqgLIYn1J5sKPOW3NhlS724NTVRa7gOlWUn73OiL1jQL+6fWbd+Hzp3L
qKdFIVuZpFtH0Z85YxoBeZef3Nwr+Ld5k72lRC4KGf/XckaPynNdUXJEQG8TdoJJ
Blio2ISCSsQXBhe0vEqArniF/iImLW8l/L0nSXlRjyFVvLYbXrhPf3YvJiC3Pmpp
AoY+42lQX54+Zd2xOKH6vKQ8z8mn+iTwDePX0eMRc60XSezZR3uomxHOSVWM2TFA
ThSKy71GoQD2sI5iu9SGB4Mzi61fuiLshbcXlXk/DtzOVUBBSvYTvRsIvMeYZlk4
PDWZSFCdcZvxRcJ1hfpgrN/GxoEwchrw8ws55NxPsvvFmnSGHz0AL3SxxqD/HND9
/Mccrea+Bn1EnfP3ihVydpXxIqX6pqqI6hT8/248tXx9VTscMMhWWRdDbdnK594p
7OKOhWM8rkxhn5P3Yy/ZRJfD7i5xah2QGo05GeQyAQorwTaYulJsZBzD2DjbGBMt
SXBmX4gHe8xLZk6fowEER1eGAGcW6QmuP1G3zgCGFI/abm/GpHOKHeiRB1Zd/T5L
9uAKamPUUYQqDXpVWbpbC8ldCuf1DGSq983S9w43WmVY0SUj+JXg0heLe/AcIOlG
Zp2JZ2Ut/W6zSRNoR47h6xpTQAD2I3DsiLxPfkcm+l/RG79Y7FBEwL2IOW+AM97W
cECwHgXC2XqnQJGgGbl1sLe544gPonmCF+ntvJmSZ5LJA3Him3aMPIp/nw4gB7kk
NB1L51eq/W6bFyXrpbTy4wBXdewpINK11eORzii8oaQunqltUOwTdi3uGHe9Uf8b
xUcpRhrswTZIzHnbTG2EZxcM6yoiGZ5vThZ84Snlnx59Ybz3ju9ltZuLDIT2O0Yk
boIHFklKSMAWplzcMbj1zedyoF5EO4yf+zbyycMkw7v15cXcXjEChJ+qug9i9iQb
NYMo+kzz4XVT6SiZ3lYGKvrUEcv77X7g3NBsndNcZ4yEESAw3QJBeoTVykxlsROf
jVuqSLw6wvsHQxFJYOOPPxxRNFB5rg3RcElsP1WpsSa2I8p4zcGPBZ8b1epm+E+R
rHU91zq6PjXTgK5wL3KYsGPDwX2FxU2CwD3Xx1fmQKvkFhyz8iiBjjGNJnYiUPj6
yZ4NTULpAVjsb8lHpDr65PENXop76a8EkWL9IBBJxMw+nHJdTuLsgcYQCf2dXbzC
jQRTQVyBn20B/t4lJ1QTC/3Or5/DZ1lSXYDXMQWNhTTpS+CuMnowQ/+rN9crKBnl
edVhr36NzKB+qE0aMjZfAJJWiVv6AseP9FVJN+9j64C02wC1KOAgpyzS6QnOI316
nDyRFFzrsoGmDLWaSQna8u9jDgGjcjvrxaMz5GCl+6Zkx5HsVfydfDfBIg4uzqYw
X51gEUnp+67fALo9+qy5y8qpWzQVAxR/SnSmFsU76qUaL8Kc+b+1TBVL1fswI5O2
c95Z+QSLTRescKef96DDGNaDTmYoEpEnQWvl+Nr1l/CGRgev2eqGeFIdN3qec0wV
iKyJCqCJQyl3VPOH5dbxsd0DYcSdwAz2MGcl9VmZ3xzgf4P1SpybenY+uBYBX8qQ
edarPmoLNCa0HhojA0mXp0On9RQtiuEJL0IyAlMNxg6ztg3D3m0EdyEBCXLzrdeN
s3qDHZXAPhf6cx6Mrspmy3uYMi/dul6JYswIpEzQ1nMCCe5wZyZ44mTKbxkJXZtI
P1zo8E+tv7mdKPnsDv6xfYK4GQCXTN/eu6fHM3gYLDxcSCcsHHIgXMfccv2LMspv
J9wUB0t3X0BFfKna5qtsZWxIV0fjWQA8lhvs8DQ5iQl360Q3HdvWsU3MQ1zBlctO
HGu1sT9c6rki5HcEOhp68H1LwIez5k23nq+KjUgQxlSenKl2RLxPl+dbS4TjrT+/
fn5c4z1uMJO0pP3mexvo0whQM3N/HPQRFjoEx04MkZIvJkPLi4jDeEDSyihG7qXe
wEH4E4EFZeDLJxVnQO68zAO0QCrvqDm1+lm5d/wGyBeyXH0U+ErDL/mEHSDj4YqY
LaEoLJzrPhpHWRXs9gX3bjcu2BwtC5tv+57CFv4a9lEx/KNFCildrhzD14VxJms2
cWePrlLEdMy7Tce4E5KWyxapZ3UMkUKhU22CLejJcdM3ufHq32aRlNEfrkJAxPAq
g+fAZCezLLxh6EvhmE8t9uoOxwGEMR2syLkp+3tp9XJoWmxhpLeQY5VW6y/Zfy6T
yrnRnj+J2cOczGI1lTL7YJ8b4Hfmb7/B6j6MhF+43oPriXynSgoeyPSIl+rpfKJU
rwtBtGQDPoYtrr5iT9WK4CLOhRhmz48o1Q53wxXNd3xiO1A5O9RaBY5bVmdz+Sa5
tuIG6oFJjrtstPXasMubijgmPavgJATMonaxMUdp0EKA9smQwvcmiJIqVdrN3R5S
NsTv6cTaAcNzKNQfhV/LhxJirF4o6HHm6cKKOtCSqOEFUQW8P6Z85EJBYMRFTPs4
XsLeluRquYtswTEkX6Wxob6ha0utzzxAraHoYlebDJmh8CnBF+nL0XPzppa7Q2Rz
qWe2mNMYjd3PmCsLGxCbHzcoFMBq7vZo/vSTuxHAo5vh8rjJ+ITt04GCsOOXCFh+
KubcYkMoDusQk5L0LxkEqLfIlIggHe+dw5Q6NyAzCIAZHJeUDmfyjW7/4BYU+OrB
6CW9HCcu/htuM9VE1nnWS73vLCX+6qXoywY37fbHTSoNjeY8OVxDRDPVrm/uwfeU
gG0OV7mT9H7uwkczVOCYF/kfy1ApGja8GIWPYh1g4GKseeSxQplLQsBpHQPqTWbf
nuYkzK2nStMObVicyrgkSdMHOM4n+ePq+IgjeL2WD3y7ltVUTr+FxMNQ32aA7kCi
anTZfMt1WOdM+dD9IKzWAHNmr61yps25IUhnyB8u+r0vdNbmej8w6NKQLmY5KP0Z
65bq8N6en0dhjVy66EjKkXZ+ZfntCx0t+XHFygO3AgYW/3uh8Di95mv999CNQywE
cs3QaMwKY2wycloA7GgBOnyj/24bgs8bZDPfo/ZAA7Y=
`pragma protect end_protected
