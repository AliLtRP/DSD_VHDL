// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
HaFzUrBUkqlb4/KRFO1nFmaaeFmNpcw1rX+SdX46fCqnVaVrmgcQ0ltK6VXckuESpO6nCOo1Mzqn
NoJqDQu+FOhAlh4FGKJwQAZcrrYobCN7nBd16RXPn1AD+YVuwaRGDhOlmGTKW31T/flbFL2PR48G
CkZwUJlZzayNhBpJ44KOISQ4dDomKXIASXtRSqDL8IHaI39Eu+2mwtfR0SzUqeryof1PNfRFZfZ2
ZSIpr3AD8tJKV2JTCc5ke9gwLQk9EArv4U0JaLJd8cRlJzgRKu1sSqYWRoYx+wF5S+5R8UldQcru
3bZ6ej28o6k0N3MvZ3viudqxbP2SXnC6IQ9L4w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
vkyQLg4qq29UbnonLsKa1sToQjFGYY92RaWFNhmw1bK+JyR2F34Xi7qbyFM3VfeQCxUCc99pkiEs
FjaUSrSg9OnPSPlfSrr84FtlPysDzpTRG+WWmaeAYAxARGcG5LNjy0fQ9hKpxsPSDd0RKe90u2Mz
BwLOURR175KMQ+nBX4PM+t3b7Wia/b0NXu/f6ARpsLwozMis7fKCM8jrcBW/sFtFmMVrxaQ+EhOm
h8yg0tJOe//4gBMTQnf7k+1M6uEKRpsNoR7PKfGVDq5H2TfigdmSj+x/dSaUMzSg8zsGpstZjMGW
hZ6hSoi+svhWmG2v/llnurG82CXrMwdAGoIzw/ecH8SpBvbtdME7nIe3P8ZcnkspOAQCn0JgjhkB
tRLqcSkoInurXx49SVljV81G1AC1sL/f34iNlM4cOavjmEzg8khbu/3iY3I3dHIex22aVoUNOVK0
cykb77IUEhy0s9qo3QewPJsnS5mM1zE8LNxiB6gwGdXaplLIRAu6HZPIcSyD3BLjoeGyJI1GfLTi
q572b7AAds9wFhIe7jOYQ2i8o7vfL4tBBO/tF17/chhGdpmc7QdHXoSSzqT24YzJ2UjWXYWrdjUk
mQbd/1aMWxiquA7LWjgvfoUFLO1Hqxl24MlqgehqCZcsWETF7yEXfr+YIFKjA+vyyj32IYISibkI
ZAD1Cw3NAdhZQUSHpA3NyVlv9hE1H1RGNZtrJzrI2lGxzFKMLYpJ0pPUKqhLadPCTKH2yxF21zwg
MVzklYEEEfiJu2z89Bfb2/BJClRoG2oYPUaai+7LxPb72Txy0IWymZdx8m28mPOhPez+fURQ570k
aTsBypT8ibOCTp+FETtVoIZTXQv3vLwy0Cj+66NlZwgWq7WukrKmcJYbQg/dqYsBk7Rz1p2paRgp
qEqbMwf5SE+LvHxdO/VjkiEvIei2GT+vslXAxkJJ1HcflfCpFgA0FuTVOOAVbh7fMOd7SkJWW2IX
YrJ+k0Po3Xu+xwWzS7rwKoHylGNu6sC9rDwuzmncKbbkDEhY0Eu6Z5wNC/ATip9F8K2pp4GOP5fD
/rbSdPQYLqXKj0LJ9l9iPv8jNz/bMtMDit13umR6AzJ3j6/uwJm2ndmqnUmJD6XD2trx89liRH6S
lZQ+6Womr7BOhV6Gh7xjXNCQnRZl/MDjOaQvVyJoMkOB2nOvHAIjrutIe2+lEyXl/3ky9/40UUm8
4ICgUuA6SQunVXv8t1GljLQLM1P1WkTRPShXdSPlBgZ6l0qPHiQOPFKhj8mLBCPdSPMssNsOdBUe
lW6dgv1zSZPFh8/OifK80znzYpSAEIjlJglM3Ca1vcjj8d1IMXtjDRpcdiCL1olZaVPOWoVWPLjn
xxWFa1TN/0CQAJnV3mEGL2MvTLwIzyiihVtCk4uaXjEHHT0XiWLYSIh5ahdRu1hRVQuOTY0nDxoZ
1R+WJ1WjiQf+AbiXppOQucEUzArSws1wQ6dOwkVznPQt/qh+ZKzGSeTiOxHtHRMuhNIdO0ySpeBu
AlkfOnNWDUunyEJeeKhw4h9ifc6GBAYH6hi38RemlnJ/bqYD4TRd99n0k01mayJ3YPkltoidcJjR
nABJSmixJ4AmKKhbPBJGfPsm/7UhUQVCGmwXQI7QyeGP66x/pgjJoPHGDhCatf8RNU/WpVA3RzOu
kke01GMnDUnRWewqqFWr0U13JpNr7o6+EXGYtK96pvScI5p+C2pVKeiFsvCwoEeQTHGm6AemrT24
iYSupJljxRAYUX7S9IcTQC2jLZqC4onh6RNqTezHXXfJBdimOD1qqGWcfSgdMyenIvPqt0+ULSM5
CGZp2AhgXMiTd6qCN1ncAtJL0NSbUmNcj3rdetStJCkIeJz61El/qnksTlxrDLaKpQvnie5I1Uc+
CPPGcEpIjNQV6m3T+KReFs/2w6mjzX3XpmZW0+nFyQtTB/QS8V1jsRMUCv/my5fO2M1v+igloGbb
8jLHsVn8MX5r0mfWhqTmJ7OKahXZW6LPcOUpgcphJHg14rGcOIbrALn5PeVP0FYgsM71BJiQ4xrU
byyn/sVhIUCiNh0qkqJebF+Eoql4q4yYJbhPPtwtNQNvRaWGxvNXchEl4nEkInGlC0pmiAD4KByn
qxeSjlpH2c64fniCDUDD9yKNYuvDaFBuqdemDK5s7R3tmAEkggLYu82ERo9CSqPx+cDck2WwqtVc
CZlLv/Qi9msd31s5WkTsDtwIEq0i7QAlUoAQnt3b/Hcx/WziTTqLOhKdjqRvLzYB3ldp32Q/nEnd
lv6k3IFk9D5Jj3UNFpybGvkc8RXoDyUXl0J7WWntYLNZvwea5IsgPDBGPT34oM6dxSYzjJHhmOKG
rrla5iHIkyQO0Emz+LcHXFyS4aiZwidXkOLVU3efSCu3+era3J/ZLQh2Sy+fF7kGWxmeTk7GCEK9
+mMXD4R8QvnKRiLyppjxJQY4HCKEArJsYKKxH9E5MBhQNCyAGvPKJ4CsxihbMkz4TZq8Vln+jCQ+
bxUJv7P0LOriK1ERLxo9dATf2Evk19ehw28gs5Cf5T8mXayggUGxgdMbfrxICAD7b+mcSc5WuxKx
6BhumX6S5OJTvz7CcMw5qlpERq1gBriwS1AgbHogeY4YiOG7Bc2AganPOdV1dfES6kCyrLu4vbhV
mePhx1a+mvcDeIgkqvjfEUM9BTstdQNFKxYaJiJIg/u6y1RfGm68oPxTY5prxZVE3nR0KqzbfkU8
3QwjD+rZ+P73MpooDTIqpoz4ctfx0gacAeWADf4mibJx76wARQdycxS4YhyMuB9MdcM6Sc1iC4kM
4C0ZPa4tLfvVbn6HP91Rh+rJ+hBSy6Pw4Bh+3IL3ZD2hX9fWh7mI9WuuP3C4CtPiZGYFgHfH0vFp
9NAVmWklwwJollB/k7XZz9fCt6lbbKNZA+oHlpUIk3gBcp7vQPod/TUokyOAXH7Zyx/7TZC84WeZ
X+KCHV8fwexujLTtvMjorTLQisEEH+xdBjKcW7xxo2upLqi+v/h4aJFnbLYGM5rh129hJJib0hA7
Bq/tXmuSCSBA1A7xIgQpZTtGh0FV+xuazu8S+03mgwOLaeBt3erPdTzTeiW+ApCedQ7OaX5Sxe3b
l46E6sCGwXitNe5eCGY/SmydCUKeEMrhNESWUxumSCZSfsFG08QdC0cId3WGwnK8kEFdr99uTXP9
GUIrTou6lsqSm+O/cuEawwDNIaSPRbGZZtx4rObaeucaVdbHhWqZeYMLzFcOvOE1ndod4aeCLkb/
DISu3JscoiZdMc1+FMgTZzKBeQHClhLVOwTk27B+/956YnxBLEYkdFxwVnE3l1AUSIsOYZOokKWv
hKUBZnWcgPWbNQF9qRoUsOtx2SiS5Z3m3ci1F9Qy6M/J4L4bZ1xdXcQsf1RyfaRT9C1nHZDcGvA+
ennFI3DIzKicBA66ezIG38GbzsJeYAQ+QpSKohbJPgKjBgrLI6cibcDHf+IuK5ZsiF5ytU/S+M7b
2wQPAwFRwlnkiQomplmPt4d3ecRcxKoD93ae0YeUBeJv8X1blThwo4w3GrrtdpOfkR0XQ7c5CbyM
QN5OxtYzZnfMOhjsJjw9V9moRJJENgr8o/VO/wcLik2STOz1hYpUKVMfn7UtkQYgrvKxZsuklvYf
NWTOwteQlEO1EKHGbQhfS81CipvGkM34riXyQLmPvFhofB6YMZxUs9wTRpuizvvwwY4zaDNf//GH
wkbLFC3R9L8tbQywZri/jchDS6/SV+GA+3Wm2y1asCeNe0lhYDh11FTGc2BV0mlSJRguU5MOwant
Q4qLdj90Qi+f6PPs+IWLZ8EaIne1HRHa8cxXrxuQEDoXhfUYpQBxQrkBxvxWau9qc0wlFztPgOTv
unibOmf1+WPYAm1Bzn9WsTAPyn26AxAitrFepJBkST+HMS6GkjfvDZx5xJDq0roM1gwM+nfsOphb
Tue0bBtWy4d+8m3SmOitLoyMelufmCVJGJMqmyCtfC9rQGGS3nRyNN/7jZXcEZUFAgDltRPevdmc
MLFsJWg/M9KHnr7o7iT3q1Y3Mk6xoRZJLyfwDf4LFGZXu4OKnChh5BDMp/DUMCdftKuPz5IKMcxM
lSj/JBgUKwgLUkBI+9dAMNMB33e/OxOHZTSuLpg/nX5JAs8gYsTONkXgUFvwda6oAp8ut19RaWN0
aFI0pBfW/yHhOIxhpGLX3pKP4PXxZhoa/MJqBk+q9I/lAD3lK/X4WCp7WGISJfeCXWEd2dSsgUH4
Ezvl5nWDZ5dspkdz2xWsC4dL/DG0raiJZkr8YkszM4gFIArzogTkDXAbRtPI/vLiJ6nZnK+z66qp
QAEyH2Gflnrn5ipTaxCCf4uLxEApV6cFR5wwB9prydBKu7dQF2Atcnhi2Zzh0dGTryQo3Rn76BWo
aKacAVaA4pap3avMlfEErlvJlNcOg1Cv0mdf+MELSIFan3O0wjPWZiNiDjcnJ4HfTVS8ss8Eq2fo
RTDvSCQFJjSSHzujStYhDtwHcYwXcc/jWfcx/+lUtuAKtjBjCHCDQhnVazvnhvQa2ac9SHw8BlSg
FpYAw0KZQWEnGiCCLCCSC8Rm1LBO08Zj1p1AXBpcD2um8gncQtKQn4urVyKqrjrshdZko0Qro0kf
VKJcMvfVnE5pZIqzjv3ZdB5Dq7yLrwE4b8qCw737AhSEMkygpAITXaBf770S62cc0LQisTs8KQjh
vULYhZUnsKP5Oq22oSLbyQPlyW2aIE9z2+xkQW3to5Pebk+MZ+OPKg62m1q8VzZgiFDE6vSwbaUy
unPoA3A2Ty32tdJzq8EBOmbiysA3JXEHnTlZxob6q3xJF/0qAPcUS+C08CBMc0yIPfSYsyYHSSGD
IWJUA6IiFsAom1w/3tv5j4HhmowU7exyivF8jmt7vZnmZD5yN5fINYv2Wqyc0KR62jE/Z2HyjHat
W/anvyVL7LzowoVc6P1/TtmX3a6vE4J/U28Cd3bDHSxu9tsLT6MgeoVv7zVn1NaHyY66vyWsdDok
ZZYVaN7A3ecERgvs/xWAeqTuVQJCoOd38kIo0JiTGlZSXFxeV4WqsK3q7v14tgMGdxvaz/9QCcc3
Hlg6XkEG2/jj74q25wD9/V1ft3Me5Pnd1Z6+5PirveHp/iuw9TX8QYmAai22Cn6Buq41ICHgg7ON
ZezRGj/ZcqcAI+CFkBX/1ckSc1fLEBv4D9dffUeMYkxcPmYxP+za36+up34NMxMWZxELBhTvCQ+Q
oZCNS3ZGZfa8jlJun9861GXVvWwJkrRg5S7FMC5jV6nVzY+EVQR7aavrt66l+fTqsnTs7erKKAlZ
tqrgFZs/F2ZqjBjyUeR0IBMe5VeLn/YoVRZPZOzMx5SA8XS1jsyIKL9b9APHtFP9neT/HdxlFzJy
ea25fZTwMqGKKIQQTDQDx++c0QFvaJ0lS2zoAF/9ei6Bq10Uqow7SYhALr2FEVVYwpYA93WEoXJk
ZZFTZGoege3wMhKNkMfcyLH3RAJw2gqWeNTekJ3oM3wGz+3qkwmCev/MDm5p00YwdO0s45Kizi5P
dBy3I6W/y3w/31qIGl/7v6aDwvwwpt6+cmCI4gg7xpoBcMvTXvzWd2MCskdMUmJJ505Cgldup+5Q
52bMDUcZ2QsDbHDbi9JCp5pOmgYiOSmTE2rPZ9wPXbeng53y82sD7rXOavhYPUdjENg5yMf/b/J1
cUXwpWmDy9uUo2DPq4eXess27TWCe1OmLyjk6ABEmN+l6T4t3NYR/GAEKz9qad3veRiKwR/NRH1M
+a3o4zTPUE8CeQuceZsG7cZAf1Tc0nc3XMTQWIbmlV6EefHa3hvWUBtJVxnB2v3mjn0UTZjsd/dA
egj2Y1iJIEp1KVvaS0f4EmVbUDs6xURaYJMSRuOqaTAZppqjNRCNByXL4xslyiMu6WVhc6GyYr7C
cee8uHnljigtEsTz60lYiI6Jts/gTuiCs0hcfe+ff1w2/xJ+OmT+FXfGucJcZaSzr91rgU4QBC70
aOnKX3AwaMDy9HJjnoRUH4cr5pLCS9P6+p7tBxaWQ03EWQC1TPRkit9gn3XpgHzXLQPZha/RcuRk
4xA0EZrJUU0mHVYlA3K1iolOs4xmRhquQkXC5R6LZDoFPDHzFSvIcMvYE+vFvNvkPizqutmmzImA
QUeckTle571uQt7Ryu4MrLU87IRAyTotht/U4TmoQ+dV+AZJIDBV4ilAyh0YW+f+7qGoQavJTbMN
4W440N42P8s/2i4CNEjHW6F4puXnC+nYZr81tH3UUoA8w4jO4dDD5Jprr7RE1qtJjz9G3SGVX2uC
dm5ll55ZRazNf5aD2jbT2tSSvx68RQsAD9Vlog6oqKhtp0P9v/yJHiSpO+vagRHex1OvrFpTiI1p
aCLq2xzfomTbIQcplzL7seK04Ja+l0+T+c2Aff8YCo1dbHs6a//vL8+uir65RmwpsvOUitRgdj7O
uXm6L/KFYydzFB5G8IPcfcnLi+B/TruVbBNrSP33jfTYXDC79OqgdeG54Mz6eJck/bEFbQ+ny1TM
VzYm63cOOUWa4uyFA8h3NzrUyvRQShTX8nxDJ5Cu4VaILttDPI9Pl3wsaNPYCDcM/rGDyy/71RQe
wqu+PSdCioc6GGu68+q27MgTEJdwLDdBr2fPLjGtSGzajk+9XtuimXveH1+am9pdk1oI9PlcEhbN
5LU6tURRTKmsFqKfn3Cz80rAGjuVG9Z0hRwFT5BTo1/xSpeMZFMaRTHYxtYqshXlyWIFqSuO0SEz
LxIwL7aZ1GIROPkHHSuW+iqcGOkJ0CCYa2+uW5KjK0oST8FaVKuNb+kLo9t+VDxGcKbCxfdcA6RU
FIQVxH4jqk/Q7iVKJnXKCbi6TdYp1nZT2tjmQ14mimEQo/KFEO3QQwRvhRlmjpE/5GhH2ZMpvYek
nmbR8LNreeDQbyWW9XlghsVcW2SZf6Pn7QUlrRFcW2ivWSXDiAN1yy2ZGgQcG2dg7UQrJF6xNw1d
ejdsVRj2kOHSuy9Fat/sVbkTJ9Ix4NKwdjmvicr7Ta7TnJpE4uBXS8X5B7oq/XIoJAOEN8pduejP
kaIGlLY/Xav73YShc2Jr/4OTgzikJG85fBYIF3UFh7M0MYPQCtzIvn/Lx7KAJKBDDOTktPaWJfVe
aR4CUwvJkDUIJkGaSr1/n88cuASsIFscJNG1VXcrrp6ykW6RjsZJxLMQy79HGvIIBAXDXMaW0Fjc
vFtS1+10vsO+UvKm7uJUt9OeJNimVRBAYMFpF3zVMhblMwGPCVLoBYeBwl8LxjOH1G2cJBEp8Z67
DpVFLqtigmkWTiSQ4SXI2M1VBc7F04FvEHkgOZOhM5tPkQaO0ey20/Seemrgx82MA32nTIQ4XG3G
TkLW1ZCR73sB/+2hezjtijC2RFtY6gL8htoHiEgzmbqeuRpJ4YwB4hD0+niw9VYhkoOrfUvouy8m
duBK0J8GEZ03XCX5tf+WHbl+LoHwJREkQdeH0O9p1xYJNVTFWtLAcSy+xjFPAgN1yJ3V72cROtEu
QDgyzyo3X1T8i5HWSdSeNmCNHyBUkBqRnY6AVBxVonq8lv3mwBQGsWe5Y2VFqlgsNMSgIjjjIqnu
ZSKnyF0cPizHNAumleg2HYHoiRIS/KCW6l04q0a9/4YemgQhooG906QuRtv8w+tmlUsPpg2DIAJ2
kTYtHI52afhxRi/fXOvJ/oUyFGPoziIiDaHQLgHwvUa8lbkBZiGDJX55H1oQ6sS/yjNWiXk3XPGd
mTSbmVkRBu8fgBEBIYnwyN9KBvyp7eCeh/1oqlXNk9XhcFSj2BKHQpGaip/tOOsNuteMi9S76MmJ
gOx9l2/0WN8/yLV/JS4Kj/Tdc6USJWTmUrwUvanXAuBkj0iPG4F4aL2wGziEbG+6eMTo45HAe+YB
CeBmFCwp9/w5zdZgIqnwA3k8UTkLlsm2Bkt3zL2zDSTonwz1heFXcJtAWLdzxCosLqAdXAGLq8yX
ErJj/YKqc3TTnS8MzXr8wJE6r7jpdqN3VSJ840/rTnR9JIhb0DsM8fHKaB9irDoSRIMnvY3u8NVq
z2E5SqujjPqFRjwltCvpo9wP1MbQKFvLgpaGfIvsxQWuS5VYK/fzZbqqlvG08WGDeUgEbhJennzz
9WsEaaiMBbRCwhYMGXaMVGRGKjyAq3n7OAkwv5O8Dw7RCclSuseUPdxV4enWkniqzPIc5w9IwRmB
nQyp6UDwYvUpSg8+r3AotVnmNptbx6AFoZPzFFu/d8NIC54rSxpRYA2reWdkOqCo89ORLJfMwP5P
s8WDxCssk8tmQpgocGNPDkBllX9tKDRne7JoiguZ+AUChaZ8zGUjdhKrHeR49YFfY9Wv2oIkkEdG
CkbvdZ3WySjuRnABRzlZ91Q0mn2mbadQAVAOOQsSjSq4kRlsQVW3GBjA6W9UcvTk8MSp3ZQFcYz4
hTuA0B061HFYEBhWuDVEXR4yqP//TEZtgsJBdNzJi4Xz0tXNP/9tUgYOeYml23/I/WHeboeTLmT6
`pragma protect end_protected
