// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
b/RdKJbq9Fi0S+dhoHR/wg4rpVfc4fxq5Bb1r6KrZ0xlMUXKQbM0aI3OwuhPhOvN7J2nAhgeKAMS
AmoGdb6RC6DPTHWM9xGYZfG5SeTIJlBwVvXryvTRuQLWY7zjWMmI5h4QMOiw/KRCESPiWlYRmCk9
Q7I/uB2Nmto/RM0J3gPsNBJxwk4kjVzFuLBQw7tLJwQ9Gzy3svkzFOYJDYsRb+Cds4+fAsmcx3il
WAFto6uPpx2ihoGuRetzYUUZuyvKukBmQ7bn9hqN1ZqmfjI3lB8BO+bjaPfCXYl1xlk7gd/EOeSy
H4TIgUazts5Ys5NNBZsWa4bnlLKMhR5FJ9gIqg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
TnSm5KaUqfdX/V/OkExiaZkdc1u4cCvgAneoWaUmbpFPHZFZLfqhNFrkSlj6jE2juyYgnX9peDEA
QHufZgZPlWz6Gim3Lzy6QE8buKHxNyQNKjiz9bzF7EOOqMaElJGnH66A8THsvmKzY/rYUu0kFJB8
s+RlsGgdf8IQXOqkPsmI+oPzRag/u1hKSdbDqErpc6gQBgm9heryrLUWmD20KmKl3OuFQx8indtH
7LlSOxlAfbGy6jcYAWNIFegA4d0eIUjM1Zjk8KombExFxv8/XwBrj4MopscmekNrwzh1FYYstMK/
0Gu4Za965U+7Alb11jKGeUYEmtMxT8vIh3OT2+76u9p2eYqVvCs/oQwqacxH8Dc0uzWs11AmwuDi
9U7q5jOzgLmca1KnG1RlJxlZtq4AWhEMJDPu4lvJHQ5xRl34kP8ie5eSj41U/2LR/REWij0WDDYd
kue5z5IuqPItprhrqWOyjmf86tYZF2pJQNhp3D+xqe4aCauSm11cHC6flFpck4/bngoP1EWbWTPT
7X4Rx6m3/WDvaLoVYRgXV3Jo40PpmVjxPk0pk8vrnjrEv+Lxsbshf1fXZTzUq2oCuExtIqtET9LF
8x7xX4pc10JGwestD+Ne+ZzwQVtQipkhrlZFUrK8nKza0xGc7mY79wWqyeO99AgyI3nvAJLef866
wBNzehjAFB7YzCTLe6xysvZlV8O47dQBRIoy8YMYq0z/qgAUs3oJzKZoqwJDzNwmDSVBrgsd0uYr
n57r3Li1SuN2qssQUbcPrhGlGyZuyP8YFdKr2p7UHfLwTpChurv82uXOt4tdlWvC3X4t8MWg+avl
f/7OCuaUeWPnREZFizwzd6CZdePRsOa1ZSRHpl36EzfIteAKZaDySxw56rBZYpu92bY2O9VZrM72
MdcD32iZCDitddgSpjrGghaScABE9A6k+pKs6yZJ/5dFD2I4czNfh4Bz7WcmQDsfyijlbdHJnEs0
G5F79paMLbHKmgtzOoJnU2tk0oP/ioDXgoHd2W8h1t6H02sMGnAYUAIL7I6HVxwBiPiKmK/3VIc1
+pbKKBvIfWcdu0TIgeNDX/CwlPNHbx/bH7F9Rj7hBq+77TsAilHeHGw+wzymbXxSZ9GJONN5+e+b
/hrqNoHgyhrR7SxlzyN+KwEwVnQVYRC5j9adgEQlcavKR6SCDMGfi/Odxn0uFCNUIkrZ7QWDj6EX
coYbAjzjmvnJyZjydRDO31G6/wa1Cettx1K3VLyPbTUnCLlEHhIiWs8OTSVKQ83ZT/Y9XIWUE+3J
mV7yBN5r9e6Eb5ylSqYVGF8J+0kWvu6HI7BR4wlWQ54MTkJqj1c2W9FAG0QqiwGN0pA3TilNcfkd
srpyMTOs3bFJDjifBWf7khx9aqqE0w/ZfnNZqTCcZKjMBqH3BI5EyAi1QXe7k+4hbUeo/GPKBn4l
HD1cB8lIy/2DNFcU47DElHt+CKLjobe7/iHVppAXs7ccTHT73f1gYHBSKxLSu/Lk8BWiiSZpicIZ
7HW+3+gDBazAxeyu/J07x9mvIWcw4vd4v5VytCGrdfjIQjvNBcPbmHM5ya5VM1Awd7DpEMOr8CZk
r1Ssfck3OLN8rA06pSROsPkh8qpEMlvI9UtxLmRO+NxYjhTQ0XrUr2UZDwqf7QU0odL3UryyWM1K
da4nQ00zIBY8pvoq4UYF9P2KYQRWYPXWxdHNLlriuGc9XLIop+Io/UkiiVrkOQm8vQ+VMDsNd4Lg
zqQ+F8K78vsvIgMtzLdopVjBCP71pq7IlGM96Ehl6iufeYJgICECIfsHWGjXCzde3eWOhRdGBMC8
HgZBvIpa+Vv1n9E3tg1zhOb/6uGSxTM8xz/QjVTn2vKtlobrwoIJ8PQqtB4RFZ/pZeCkjtMhY+Z3
b400M4/UcThFbY+3MMWBxQwPgIVGZs1794gCLb7jjoeOWsArnnGi1YEPTL5YaIIiEtFeZhnrTbsJ
kxEYsLyUWZz9dIIT7fK1kGBX/6fhnbqNks382fNEzrJVLehkh2kzcLJV4XL1+3RGz5Um6Ajq+WhJ
LobWPiH6KPhoH1y0Q7P7zol4nwbVymL0mPWtV91szHhtN5K2pHg6//EiDD0yeWlDjP7hJP5Sp1cU
HIHZWgOgZQlt19CBWv4iUg678rC+F1/N1VQTaZaMQbzx1TJOtoEt+oz/enImL5ts5yjUyQ89pyuv
5BTmCDopv+g6pvX1UKFqHIXtCh5gKNSRx0ARE9UhsWgOS+x9PtR54Be6D9Zm2V5IJ3frzH3992ak
IHqNMY3yZ8l2u+aZBgr30M18TqonO0jR6qHYB4c7k17+Q8CBYF3gvXcoOUBmnnWjPfmGUdlFb56q
opoa8bXUOmTG+LkqRkKzKyhzsEtk9n0n+1vdYXhUA99lqKahrWFOTYUmFYm5WwybyXHtsRvC57c0
OlEb44smwys8PGh3iOhO4OdLc9Nt3sP02VYDR2FHYGfm6hwouUGe0Mgn0KKffYPlKylleHkNHAb8
UeyN6MIrWOljoKxQyBbVGYgN7oLOcEE7F1KUBgSN4kyvQ5EJs0dGAUJcZ4V6D1RQ7zJUCD6lQXAo
6I/BeXD+vCPANP8ymzzcQxHe/BHY8UqBS2xk6gQb+VZuh63al/WLArs6GeSG5kZ57O6gWFuDc0PG
cX7voAL2sF0nZCT8vbBV0keR6JyzoyZPMQA9tkNfnrELPN4TJDxEVL9yPg2jY0tQuxzOOLpAkzUA
bf0BhRJ5ed7GqE1lnrTD0V67TPoi3t9Z06P5Qiyr7Ooir+DB98VPHoMpiM5ED0KYesUywGLE0fX3
aF0Htsi2OAoql3myCYYONwVkNAcAmr07sz3VET3y/McXcVAwx+KC82WjnOMyLZECwYWYX+mDKEev
BHmhno5kwj8XLMIskjoNu1R6LteWdHSotm3psCTZmLCyUEkJnOT+PN0KtaRjqqQuY0apck2TinHc
77dxzMT+fY4xNSxEzLk93PJDqUD/iCfpQvc1827ltFLh91YQJbJp0U+gWy04y68ZEVNH8LPVbB4i
8G91+ogw5WvJEM7rJyOxpkOh8JxvyI4WVczEWwStg3z21ZB8G+4tQc+u9T8V97kKDcTyYUHLmtjZ
HtneTKTJzUQT1c/rjesN3dERmRvChMOyMO3aHGHaRSEB5VpBOFJgBQIXlnaZLhThB0X6qxaBTXIw
O3+4TbX8RHf9TQI+DLEuoeruW7UF1txWE4RnSepv6+SACfRLmCqs3GWutFN2kobVXd6HYbRiVWeX
I9Ir4+/dPRCxdS0MBDhxL0n9YOiOcteDK+frv3cQ5NStRlrwiclaw+awUexr1V5BOe/+d0zE5h57
jpSQTRWi0sWsSzBhr3m61Xqfg/WM8Jc4EgebEUXw0xFNiiJe6Oqwddjix/76EiytQ4eE++Q+mFsk
dTcByv0Is3kkb25IvuuSlLkxupmJtUAeuHwsSGRiV3FlYK5bfTa5dAKpSRoQGLS/ZSWQSucj9xUI
hJUPj18FPivNd4Ys2lFBcQyz0UmIRte1xaVPqbsY+MxJQGt6qRNq5hHdHKtdPvR+SEj5ZKxkHtuu
4ylkRR7cOsaHmAq47wbWc3960Da6zp0rxqo7MjBkDkNcqXjVbYmGtJhpV9r3Ytggl8uGrJGn4+dr
y6ADiTLKRMUsoXfRr3riIBuohrSW49Vxg0M5EclgRoRNLN2qFYBt5+HZ6wgpv21AZgKIbVsBDVK7
Q79l8eUhpQbcEDyPCF2Lyl07QEC7TuBp4fYIxB5XvFIXSXeOgsC8j/nfPNx2kfpCFBCvpRzVJ3nY
I8QGyRvTLLkoSLmK01bvyGkIrA0dMwJl5AsvuemqyuqiZSrO6V37KVcKosVBpAUrBQKjB60TWAeO
EB6akf++bImzhLVTpd7FIDEgvDcgq6oc6Or5yy2yDRCTbpVLoGdA9pk2ziAy2U3BSSn6sQIa0pA/
IeL7lkO7chYRSR4TlIMNjkcV9hJ8PKhJjVDkjig7MUJ3OXAnj+24Ufx8BXZATpCMUcGnmiJlAO+m
3y/nP45hoR0ZMF3r2eRuZjGrfaNoln3d0S7vP9NfuTR/Xyqah18jmpvlmpZGdqyjcLEfKZAT4ki9
twlqghId8TEATgj/AcQgJNTDl3o1HD549QW54qE8yoXaTMFLpbLyPO/0DgINOJ+SV0Kr1ObMM+GO
d0t8NaLD3spYCKQLMer7bsScxgs1OwtsGiZKp2ILTujlfXL4fPBPzPAkLyL2HHXJ776tON91R3HU
dEX0giyae0bpUP9Yp0CI90GJ8xtb/smR0wNpkqnyfUBffnMU7QBKBZDG0+FssDuXMODnVh8w/2NZ
xjG+fdi+N6vHQ3qHwLlD1je9EmO6FyX0E+1CVpAl1tmgQCzzeX5OvuuZkI28C/ScaMm1lCCGNlnt
+Ph3RNTUReLuQ1B+zQnBL53yHDvKXl20zh0l6p0SGhN6LRHp9fvesJbltk0YQFwEQk+H/qPb7VNM
/4LHbSxBtLo4q+Y9XM8T8R8RGHBzK5sZujB6mS21aorQpNLux3kVEMze9xMJ/s0/ysF2YPY6UFL1
2vTRnBSN9vN3KzCV53arKav1bletxeGxlJRx87rbfGQx7rXawjmwtJcOdKA4a9b/wZuhFrUUZMfS
LFqK6ElRdhx0PnuaSby000x6tjUk3jH+roABclTcTEISqFBIsxFZj+91jZG+XCKIQtgaM9wgDUOJ
7KEgvS7sCwzMqJXmr/EFet3xx1YmQmdyit6XdWsi2N2jIjoXb2Kp87kjMDoGqWyUno7guVC67chY
+DD2b/A/OtfundJxYRdI7g6LjJPg9Wk6KK23BXpNu8mgRzcndD7d/65jM9tjKUFHGbTBX8ADf1ef
FYWa2vVvq30kZBa4g+8HB618YsH35ak5ptoGwuLKQrlT2PIP7b4BaItcEVPrlJR403iSvUl7huL0
eq2t4Q0Mhpft3xBmjKYPDkJAntF9+M0fMh5VKuoo0Gj5CiDq2wffoCnM++wm+8cfg4WyY85gklbb
3MHxHWrOiLLpGZ94wcZiwghe/sJgQ9TktaOJbZVcNwUJs5EgnZmqd98y3K8KPxH1rtaKR7gAoUki
LWXvJU6wiR4I+GI2kJSCrsU7vr/rG3ou+xB71KmobCRgsp2ZvBmM0AiNem7Zwzl6U6XMDUBWtEoj
N6pK4TKGL3ZpRlY3cxN8KshpRTbWN8u24dErxQ8uRU4JX4Y7R44IwYR3YCBrxipNqg+8LUicnHAz
ao1IeUH/UW45MaWLucpL8rEITCKUXSnqo0czTwQ1sYbaDwgqlX+XvQ2angcsRL6Ge2TLG8x6qJ+i
YECMJBddb64EdCWxvWI382USMMXSvBYAfiboEmJcm5NAnJOsBET1rtkj9gL1X0k67AYxrL3fzRY9
S50XvPbTJ/NDB0I3d/Yqr67Ael4bpeMzcozTvnlnzhwj7AAO1w3uU7eDBMMxdJ9+YVedpmeU3AGa
DJB1sFuJzVd17/x+a5fMAb6sAwnFJul+o5NkWmXlklX804Xf96qwoj70xn1DleWwDxYz6AfhCnB5
uGTZv/8zPFNc0kz9/gVOAHMSCbu8vyEpJ5DM4asb6/uWH8bqgyhIzwChKBybBB3yEUaxJdwMZ2Th
8WCcjFFZOGREcYuH5AMpiWPAumvtNNhBgLmIgoD4bmflHtTlacWlziUDvRL+ffKOjQObD4fRdnYm
eW3/KIqEj4vQSw6mqcspyyttHVvorUYf6bg4DzDpbd40/VVSbftohM3gcvUD5SZKHMpAMLJ0WEmN
OkH8OIBxZmrVgEar/AAZNwIzXokXVP5xxrw1Vl5jOreYIb97o2Do/I4DOtAvRjGCqwLjwD/UVQhe
QtsL29o4bTgrEP5Rg3tl5xZZ2oG+Z8Z+AIHvKkwOebRj4djuIYi0bYnFh1Ypedje5Kkibu839MXp
tgpSDkPFGPuWoPTHL2p90qT+RAUNPnq1OsjCXJPivvihrkW+bkh5VuQV6g406o0XpBQzjzN9L2MR
BT9lX6s7drQOACgmFccEoiMWXC5pINlfTWhNp4l48oKoKlMg7tuokNhB53nRYnv/oQ/qMSrOrl97
Rnzjq3dKDWiFL/VMWmDyhJ5Cx1vKkqfvmLBUriRoBf1+E0eQWGUoI3RZDI5I9jF+rkARCwBAIrg5
JfJICEdbVDVkaWMsK3QyzD3nMRQoIJPIkISit1MHPUi1+URFQj2tbLEKaHqlR0VzpDDmrPQwpBZL
U+ZetQe+VRYB4ZDS3ee66EF10b6tyBos0y9/fQjdVbKPEG8c7qzuqYVh2viCZuSChoojO5YZjIXn
hSYJeDAenQHJOPNNtf/SYztlcTGfc8fJfW4L/zF9hhaXEsYa7/lA2fixN0yap6uAQZutFfAKkI+Z
MDAq+o6na84ey+XWVqG9ZmbP9LBReFKnNOLGCqzEW1qTqKXwayJpmSl0QvBKP/ssw1iKrtPC/N1X
XF7xHIm2T2g8jDURUz5toi15zfou5KZsoM+0bDK+rxhBOj79EINxig+p+b2wCcq1AnbZQcaL9D5C
qIZm2mkUeoOIsXE4zoiYyzVP2531Vcny2AjdjPBgJyjKqooX05R2XvtvzyJugqBjIzqG2FqjhnEY
7cbylUMvLJgk0eSbacmGIeiUS4mMTJ3vL8nakkSqNAt9RSoCKUYokdm1kkN9YAHspQ1eLNAOgN0p
8nlUit8lQV5r/YVXOdgpSWzR+RwuntNOp1HnrzPwMQs139rFAWsYvpYYXv0eRzfLE33BUOXoXoNd
9xL9m2+i3kaP8wUUIm8wF9JWFwbL2A5iCs2W/FjEyewG9Xf5lhiWYWg+jAYxQKBZ+5WMM0I4Pu1U
zM0wpQuITUQ5jmyLS+Pgg6TZXNUShgBQaEQrJJZvkmTHsO42CEvPtdgJegEpWQJmrNu4CwxNn0HL
3uA4qzyUqBt72pqRnYlahqrxacLsVTeG3op3sttmbME44ptYY4C1N2GsvNQLpVKCztfWHqZ3NM9r
M9ddckxKCJmrVrxh8GLuZMlD1m6TxGW8d5WnqXxhMLJ5Ey/N1GDnNG+kOnhsIkTvX3cCmHSMVQ0B
dRBJGn2GnQSApP6EzctbcPRYnGhvrtGWPLWvkrvV80+og0t5qmlBmjHWWhXs8LHb47FRm4MCSDnd
ylm9A8EDVgbIxx4rB4NzVyYxYZuqfmVjxyCPajBysbFP9uogGDYJzp/lLCGbVMrtjOVnF6VJvaUb
v1Tjp9mnJvGCA1cMc3sxJgO2feztoceF/DXBcwR5sp2/gaJSM4kpwy252j+vZVfLnj8+TM0y8R65
vt59cnIOBt5kFU0MPkyUWP1m/L5QyDdz0TNsao6CK1CzROwnOZjXFyDymqdPFbKDIHLWTldl5icP
mGlbY7AXN2gQ2qlN0/X57bMUFsIgAO9oCbl/nvl4IMu2aYTA40xl+kW7q4+uAHSyszasXzDxvjhk
EogqNJ2K9ZZJc3B6uThIHq9dn1TgDEW37QqptnsnxkFE0rXsDetHL5fn5aqEVeCD7vDPz8BTVA/M
ecXt9vBDVmbOmo2KtOoZA49ZzRmK6FWPCO1aI+PjMpzYvmYDMIlfS6Ep5z9Dkz3w++ZIIAQcbR73
CFiT279iFlYha+zvo1PT/+Mze2VnyEuZjlWQY5x/2uIQYeobhOxgmgM2PxxZPJOZlVy9xr71foYj
e/UPpROxMbsm3mR3V1uZqzWtqZbQTANVukM65WBNLAEqohAh4ZhgV8u4amwTRrIFroAatce2mo4M
ZpRCoN2qR1616r7ZkKp1nX/n5BKr7+zyae3jAnO1f4jxjOOB5QA1yz4eW9NJk3NGJYvgnUnb5PD8
sByLwaC0YKt/L5zbzydr0CzyO2BXFHA3f+65jMxC0Dw6ozedbTqvmRmaKq82Mr5v4Eex56YbbWlu
WRBtOBXWTh4qmlzR8n8HlwUIEkgoPfNjgMMRXqrsMc3KNJFcS87oa1zQLcO4FThVL4Y+Bw/+KPQK
bZF7JPffi/57jrss1+pQiNr84dMCm7d/ELok/RGl9wIRkvnhQGj1uqWsyKrl95GOSTQJ1Pu3Oo3p
1413/8ojUoF/Xjlzov2Gjc7K+v2MWxDbFDcEn2q4kL4n2LDUySFTEGIP4gEG4OJIGjup3G6jsjnM
Gs41xxxlzuKmk3egrNTcczo23OvqONUBijQ0kk/lbfBPHt2PYBGJ512Mrwqwk0MDFY7nSSMvkC/L
5a2imaj/kfsQO/V/D2c6QZgc5j1FFM4xj+uAxjya0qXai6GqBLzWm4EAbrT8xNCBtri7kQh4N/yo
4SsbYX+aGmJKHOUjXwGNfiE5hzIDOsUby3GcTc73VcFcS87AVdBzBDtYPDSNiCFUOLKj4fg3sxIp
YzxecfDNOaRHIeTCLWsd2dbr8CiZi0JjTfVK3tS4UBH/spRHuOB2/4FtNkYsVcMtUFhGKJj89rei
EWqVhhehtfLarVv5rS2gjYENHgreXTsQlPqsvU8WjJpXaf0H3gy4yqZ3CMSDiUt9gByo53IfIv7A
SNWUp+nGal0RjKDIif6Q7hj9/kWTN2lOQhRh/Bry7OF8+yuHo0LGYoMEVWycGOng1eE77Qxrehtx
0OcCUe3vLhRJqxYhKlwqDAwTgAMKeKlRcU8ZN1z3qVYQRJ4THeu2JhMMVP53zknheVOYOtlTIO5L
k+8M2VazA+4G36y7yRKJ53fK1pPhFXLEoxhOvH9IvXwoSqc4hEuITP6LVwZEeVKU0oI68bLYj2eO
9wdwQlo4y+LgHeMSQomqoCAWcs+IH64bor8Wc1Rk3vZZOYMwWv8Tb7fMMTQzhUDFlM3gxbcCWm8I
GN8JamgdxDKZAiZ157XqsMRQUlF4tdV8wSJKVfzniII4s7lOfT4kJ0SedrWT7lAy/a/qCYpa5p+k
7SC/Ez5PcIzXcIS632PjOpQUo7HqQ7TveqReqItP0d6QK5NAGzys4uPHOM/PsRX3GsYem3ShPn7W
2GrxvnWhRQP4ZPbodXmSP+waki6M3CKnMwPpJlJVSLgMOGoHhV2ykMXFVoZ/0L4udYSNM2Hh/yEf
2srqceUyb5K2OVFcLgKqUYbmqUwlo4RGA5Z7GFzLxqPO14OTBouMu+Dy8xCG0yDIJTsj9dFjeSaO
YzGeHDXf+QOMVREwvsKtbPQsTpLFFHHqB4x5WfznMc77gpYZ8ueilftmYGCDjC1wV9mm2a/vyYdX
vN4ObLYOzYtVdy759/3szss4pwEmz6nncc5sMzR4hP5nNl2ZLbJesTYn9a82jsZkFTYLsZIy/WDt
0ph90UUKXNA68BJpncTuwz+HPmcG8uAu7kdA2etqNLJKNWtdHfBMDKunONwTkTq+4bW2+cAAb8rT
PfdboX+wDDQfpGjrAWtrjF+1c5bpeZNFFVw2VcJ8qS8QAgjsU0QCcJSYawqLhdWPfc5T/LUbcKuB
uuBnvyPe1vPsqLEWClkzm3PE1gtp/fHtT7pEZyL8bwicyoxKzAFBoKpxpIvdQJiq3FetBfvYjZzU
jRCMKjZW/wjdonxL9qKGGv3wRMJudNXCU5H/9zC4vYf2aTmnnJ1fiu9FDsJY+e7R0vVRpc7eMe8e
jKJxYjRYqYIbKYh5mSecI0AZhYb78GwtnxksdrySVZgNkuoXOoku+6y9iH1gIBG+tqL173HEKcwt
AfbOQzLhXd8jYXHbqFe9zgtqDVntU/xFaRINKAtuC0oeQAItcxENTZv5xQjqq/t0Odbvj+pJO1pZ
cTcDYUy/aERKID8vivQgM4PDgj/icu3tfKc7RHDc7qwhkdsTxTg9wY9sIsdHFf1RhhU1b3GZSsBb
44KfnP9zJzHZAH2tnG2UHdsUoQn9SEogmSbVh5bApNt4l90kJviOn5u3QpNx4LQrhkL1RPfEbzIC
DbtfuaQVC3sBgQuOVciDWJL28TUlYb2je+3XA/9QL0e6Nr75hbgvb1WDPMpsDtugkn99+jm+nGTY
NqNEea0gc9IWUFaW31gtmlpEiyB/XoBh1hWSHAMgqzkbvgoGJaGsv+I0OSm5QE7y9hJJM+5ZRRn1
2Xq3bm2K+UmQRHpIVQmNNJykGjRBe6IbF9AzGUrAC45ek1BshnpLDdVfNu+OMfvwpa7Xuy3ZjYOv
q/pO8qqYHHhtqYksnDQGvLvCFJelJg1xRH0EqW/yZxD5yGcWuFZuADH4da3xKLb6yKb6mBpL7Ew+
23BnAjRo8dFHjl3WjQI0FDsTBzsGys/zmdzS+UzSXc44UNNzbpJXzc3/ERog7zSkmhJZ2MwwMO5B
EOssXH6pobyM1OOHeQ1wb6y2pB1rjIWBpMxijvOwqUQi06O2JnIKQLvXH2zBYCrYHzW4SIK3EKLD
DQrbtRn1/2cuYo6a0EsW93SUlJc9JmyVQkhH4NHKMYBTKcQ620YnlB6JdVNbPbgNU9IKySBeIa3F
lpb7rtetmYlML8+AZbZjg1BiVBfRa2L2HidEX0x8ST9uC1odopEP6XWQsI4QRYtnJnLlJ03QaEpu
hRv6D2uS30uzDynDIgVTT3JStmxB60wqdgsnhVr6ohgJl9J9lFF+FkXBsYaR/pGFwxSQW13pwcuW
CYbc8ZQ1TMMpJeSstfV0kSHZnpss73SRD0UwZIHNMWF9R1WtMwnODaydqttRRZzxxZA3vNUnbO8r
tXuptLofgeUBQT3d334EGygQO65qsleow21BGccRTPqTJkAajuJj6qq/OpgrcHEbLwzBk6P31Whz
MdHCAeY2+ISAz8Hw0nGiVJmMO/Dca1uu3qmYdfwW2uq+1avYCGAEb4MY7SHLzVPzNUSD0zphv657
H7JwL4/wV270qUAaGVWoqlyqnbAa/jLLEe1++5YZ79FcSm8JYewlqOV8ZHVlGpSat1IPS3bp+W16
2/CNd+oIaXV4auKzTmA6r2IQHpOn72U/wrgbvcMxBl08rh/JRasJTez9OL8xXtlrZOoz6kdgLttk
d2EjczIx+0hIW2mxwHfoceDKYx39X30nc2Qcnn+mZXPryMnbYXAr8it3BoBFXehyISnQHoZWixd2
pwP+JO08EW0TaoYtsKyD7i2veXEGsoizcEblKx6WdeVEoT/rw2uvBxOMmmFbe5KzeFxY+uK2ojX9
rYXY1v9sW7FveMSy9TdRHexJahZIC1PpznTNAJlmHQdjRe4j0+KC6U6Cubiyh7UoYWLHDBfkJq9i
zimKXb/GLxycG+v12VG64VI8AdHy6ffw86Hn6aCmtoBHFc7DMfEMURvaia5vXYQozGTpciDfrRmn
JpHDW1Ie7NT/0Wtq+E7NtxZz22ggGE46puDOl61sEucjlbLPviWwCopTAbuCfNG+0Kj4h/wbg7Jf
zwcArmG7HX7TewAtwUIF8nQBI3MgOxSLYrj68bMoNPE9Yr/DLPnrhiweOhYhAbInRd6qe32+u79V
f9wAIJKIhPiCF8ZOdRvocyjYDWoTGvE5YZ7AM7cxazSRtVL4LUuzOnQ6ZXjSEej4ZHCjJXmKKu/m
smrzHI/87rqUHdlcnKwoa4OHMc1B01LHU2Ni4HKYzGfqfju8/sW+XklkPdA6D1M1khGzXuXA3j4A
aEUwXaMNK93Oeuw9T9TdwzYutM+ie8PXlX6bwCkj0/WXoI0LH+TlvUGeru39kgTTZtDq+2C5yTwr
3RNfCvg1FqJXtOnNpvtH2BWC0gxl6CvDbWc07E6mHrc8KwA7vjvHw7aSWonpu8KckKgu6rWk0zBV
C//Z9MFty8Z6fZ9BLx59/mtM+/3J7VpM64AfikDz6rQxSG5XIIxmn/1SsXqnDH4JiaglbB6yvvbD
CtdHxqCZQngn5hIz6o0Y8Chfjd13HAHCHY98/htDvIhiVpOsO4PUOtv6qwpPFNU29N5RgulkXfGw
g3sW1YvI6EOdWsgdkc4iLv2acIsQII+o1vGIDWG4P4FrgHWUhU8C9ihyjfV5LbLUBne0PqLuwszZ
Y0PHKBM4b+TX8h5Pq8BbDZ/p5WwfgUjAENMrrxyi1rjht6fgNTBw9REShBk+ocpdRSqWaajYuK7Z
ch5R6CIjdQf9nYdqzYtjN1cifCImcAfesjx3V36WpEhxEpRop2IEJBTdKe8sXwlpqyMbDQnjeSbw
jt9o/LqbkaDjpxgE1mhS5g1+P100cjmglrq6I9Yk4MEU8MGLcxHDRIBt1EED9OsEPVgloLQH3d7o
J1f8ImO5Y/3I59cGb3GUZT5O7WJcxYWRWp4o00mop+2+YLH7LhzBaAihHCHJrUU5Z+U8Fh3V45tJ
ONowgVfMwovGGB2j/RGwTWeYF2qSxcqKQMseqDCOG0WtuxgjNNWEmGMuph491gnejWm+hGp5q4i/
EKx/5Izqgbogc+9lMG6IUz4IGiRylrRJ6xH+Qrlm/Jr46UwyfaLVrBZ4zzxikJOpscRDHFwXyZyz
TRZh7wzgv/cimXFC1C6SD+DDwDrJDvYinPqi8tYW+QO2TiqiQTVLdFr/uXYn9eXk7ODGTTLiaMUG
ADM3v6h7h054Mts23yvCyr3SNflBbCv6Upmkx2kV3LwTjWeXik9F+PwcpqB2GAsFh8Nbo18cqNkB
49uAklKlwCcJPfRpk429gSGkLjA62DCxbw1FcDfCF3l4tJd3qdF+jcEcL4hTCvRtZt95xkHN+rgB
LEHs3ygc4DMLRevhVvdH1jARAALtt4NyxC9CFfH146KvCBgualimRa/DCI3j2KaOYqBCWLngb7IF
5eGKbSJLoo7b3xiDs8TcGdgd4K8aimFm3+/y7DjYI6ZQWUtWcrhSu7hzg6Qo/oYmxDg6p3bAJjl8
hQKOXj6Wr/6oHb2DoqD0yXgqo/MDTsCtH2pDf8htDePVrJ7qHOIj4JX0PeiTVolszCp0vpdA2oaV
uXDilZPHP4kSgjRnMfwDDZ4Ehp2hq7u8+fMNompBypaTlHC3sMdqcoRzPSyGfxnnVDKETFWRX66E
XUEWDAufGTzz194R9xFkBVOv63ozbWFiwYElgAmu+iaXNZ/NaUgKPiYIiHhk+W2cRnnu7HSlZ60p
JbPxmt3U6pNCClAzkJYM6MAfGvh82NZSb8AmZGLKFvQXgnh1yXxpPeSTpiRcxMpJwszt9ZRWJ42x
ykY6kdqTUTo+Wa1NImGZJkO52A8vximTjnGjGeiV428gXa7p0YbT0WwHMXcTgCBWrp3qQwK/Bj1E
1O6kYf2qrZe6ZWvGtbhiVdGX7byDPIZqFIKSOo38s+G4oEqb79TjtB8S/PLUWRj8F6nar2eQ0HFN
r/IlIFgfczf7CzaAqb7JmMIGc3+oLbnDx8pUzPXrtDm6tE6K1mff/o80l3xunBWzg6Jpn9ZzonLr
kukabHHPg36SLBKqeu0Szxlu4vJqmHXLQsJuZCOn8Xa5YioCF8+01JGXVnYEnCeVZO0u1dH9nPz3
CYEBH8N66mZmHD1H4b8lEsXV3KEVW+9Mg+7hAWbEvGrbJIinUm6MGByZq6OIM/h8+2DByeOP8V1Z
VlTPmYia0jip9EtKEyzx3wM+dYsi3ou79AlIWo4OXp2GOnj7Xgyc77biaLXfRWkXsuIOxFWrT+33
FCkovz3k5xlUUAbYrmfo26KLOj01ZXVFr3ndIcZECBXOSXeKLAFLo+4Hhqt38PCrstdAQP2kYhHz
OwdZZqUISw+jMMe0rM+i427U3HcWFTyqdmuneE6gvAKaQbLY9Ik3/zOb0qHoJksayuQM8NG2RBn1
nU9Ca+Kn1ffgp9wK7B9ZVCcdhypSgCZdKVfxW797CAWqljAnaPMOt2He+U7613EbGLZUiYt3M5u1
bcZ+k3GFp+cEWthOCVjn3zcwztuO9+GOnHgNB97IL+62u30tTeLJbZIAKl22kWsR6xkJyzXJPMEJ
XAy8MtgZzJ/PyTUTfkTqjA/G4X2TC+CYH/Zr1DPbrCR+L3UsFjwpFWXYDJ2/W5udzXd+o1TNpKQA
sZYNjgoBSE0cTrXLeGfWr87Oys52wEX0puzWjIvrS3ygtusQTmsQpwLfRbyQMD171tHpYR1isCM5
jlJNNkz28jMTAKDVKdM3hirsLgY/bbSHG5ZXq19kl+xMoOwG+4FaIuMPskLgsB/X/QDX+eDtgZye
zqAYEBq2Bh0NoygTNYutFZXJvkXjKYZ/k6x8Lz0LxOFGMuFsB9b62TJxZEu0BzvGsEkhWuNnD+Ea
KFvzxOXHxSRQN0LdKQw3o/MiIUaQ5ILYeDxvdtl0IyZ5jJWsI67ExHdwDA0JimA6qS2lH5F2/mXb
l3//Vgb0hl2UO+WEYQU0UKvOvG9AGA7dv0mjFJgSchIJHri5LJu49RpIy8P49UQwp64/+e4B/CCK
PR0VweLvBoB1o3cLzKNVeZ36AxXrKYaNukAxjJx0luvFT4PmtFrsa1tWJj51mGJxGOCiRtD1HaDO
kpd2ifyozkP1rUIt7TY5kyHgouW5+J5K9CgDRMdDWMQ7e1hHiLpEmZcLHiFYdMfNirj1krfX4H/p
Ya9XvmjspWShqRKGGYyeRoij/DErQtIWFFmXmASy92FHiWKZbSGSnbWb2Y0eomLzrHI3mu2oDmOM
IzC015vU3sPjKB0gK/6Inps6JcNdXMSPQzoilKO+l+SaMTP3nTR8UzjPDDCLzCggYPn0ozs6KK/N
vMtM720DHEspyKfY5ORGdRwwo55LtMW2Q7q120NSUVWZDXOk457e6CYp4DqZV1F4jzP8FHLuEnw7
OLDzKbui2UHwtiHcFN5l5YXIfCOq4QcFgqHhTP2Xt0jDjlkO5afDtgAGBklY4/FUYo/qdG6Y6XAx
oNVTES8pcwf1xpx80wml6+cUqpkMJXsmai2ENcyOfquftbMTt8KsmWcEVxk8uanDKn5r2aYAk9yj
aBweChaaUEoXHEwc4lnZ9BMF8BPO4yvpWqlZjNZKefTuQNba+kZOyXxlKw3dbeypuUD5jHUhVQBe
arM5MbeKiS6QKG9AnDDxm1/Ukpe641aX8YHppw==
`pragma protect end_protected
