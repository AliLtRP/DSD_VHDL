// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lj3R7Z0jbcEPB4YZdfVViMi3T18lzoExGF6eOFOFKDg9x5GMYL/mqMEDNJleIN9c
nABlLRaZ4NPeBDxe26H4QbcFnhi6m1EimMJzkoejzI+MTkQNCfGNLiouHKcd/hDz
D9gwDnJrqBX3/zXfQ6SIlPp4bzXSgTPtSpI7rJ9COGY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8048)
1SZQ/JgUiivdKpQuNfZBdArzTfBovfqFwcJOI+QK3wow7+ts+04PZd0jI4y4srrm
YQ3CU7E88iv2bFOiQb1BBtNyktxOooUQSKfSMFczlzgAsP74imeBgB4tsQebrXUz
R6mhxlMjCLVCbtEIXTSUjoQcdfoBAgHv3il39YBIY1laUMo/nfHqFwegxzo/SI3Z
mD+reSRIfFJUjnxbhvVf9oFJZKrgHvZ9yAPLPzdZNyUY4+PO3OtYmyMEaGKF3ox1
JK9XdKBSpJZ5sG67Vr+8x+GaANRNekXujV7XWLFd8YfQGxZ4cDO+puf0aMsIs98P
GpUBiCkDWo770oxl/tYq6v7PWbDJCxPrWV+r65L6N213vht9dgzW3a/I+ctVL7zk
1UNCwQ9UdskvXG41VIwSPaCsQ4wJh66eAGhY1L8xuoYIArONGLlYJNM9S4pvmPBS
Ix7WdJSHsJeCTKI6OfUJgwXyT2g9ugDra+WXn33EkTqPSts1ec/Ed1zu5D8PQUFq
HRdT8Tt7wOM9/N20pIDEpnoxEuawbe/tpb/ZmnyJ0rm0F0q1FWl3TJv3krFtFMnT
FJq7P+pRjAaHfHOTITOq0NpBC4tiHOEhl+0Et4JhD0PwPUN54MjBuhrmvD0/WJck
Uu5o/7vEAD/dCKYPHN++ZFTitqbLgry2WXHxk9QKfQ9T0koyfVTm1K11M1oJNWCJ
QrwTS6zLM8iSC36nNVyM6BWayVhZSxvoBpG87HciYj5elKt1OrhXR6zsjyO2n0vo
v970rHJN7O8a/5stVWno1F+byY70Wwea7UkJdLIjTT6v34sxFw+zd2hwVXEeoWQu
FcChXJ9eK+EaaJPerBjp1ndtWNUofMeJLhpj5D1tTvmf0KoUsSXo0mG1we7e/WbL
2H7lEqHnf5zeljMfpgnQhde9lC4pIIR4+bZ4jQaVE+O5d3gq9yswQKz5C5vnsz9D
9lqGrW755/gbA6TBvHmgiL7ec8zL9WC/c8G+Kj2Os2Fkel4ROPkvsu0BkRiXRDkD
mK3FBNplQNhbSqWx8WuDnrfMqYu7ZZVLMCNCnJ6qvCesAp+9AKqFhfaaoah57x9U
UPp81pcmpTdWe8h5ErYageC9gkYMR7tymAPxI+/8BcjNRQdC/5pZJ2Xd8Qtvu6dP
FVxDY+gvfmV36O7ZoaQ48UC64c10RU+oJ14DziN5Houz4qEOhLZpk/q7BlSbcjMz
lcSw78KWZN1MCop/dSiNeMtPJkz7wup2r8UqwNJd/E00ipp7KVVXglOXVYElqpTO
ZSSIm9ZlvFFCt4jCLQAbtcGZL1E1V640GKu+PkTg11dRHUMNtn4NVl9Lfr8bSWKt
gjYFzKNH1SEGw1AqvwH+PpUXApw9tiD5ssruTzgqi8fFkKxG6OVzSuT9NRn9eq9R
fxnwBeWhgl1CABvjGvlTUwO09RljTzZdXFj6d6zevreXj7ZXoOmDK0lqDJxxZLvD
RNH2+UgYMfeY/EYCkjRv3pq6oTD19eYdcdy79RvVI+l6uUdfn1LU2vUqGw+VTcHV
5yJZPVdqiwLSdumxWRF0JfmJXWIoRF32coNwH7mX5WAMmetp4YXii/+jwxXUlQx+
rnaQtRzhp7mXeRqxXZbopvLWILAZP8rLcoGYcRp3UnwgpFKokBRDFK95Wg/iaG1E
P43n4dT5/+TwlHb1rlJeYZgrhCxGh2JXm0M7tsQcO2enqp2Z5xSCrLYizGymgEBq
X3QQ6ZaLoLkBpZcZ2eOGSFaKuxIfvprMif3sb8hiADYu4qZyKQmIWqiHLytFUjUB
5IDrfw6iY7oc1u7e4tEY9itpivauKugF/e3UfXM5K2zfwm9GT13Rlkm8R1MSbyRy
fbNbGmpce9GerCQZ2e6z5g5Lrovm17BflmWNcNMQuK81a++UAJEKyVLr16NCHoWZ
W0F92H6W0iU69LMGUObpI8Tly7JjqaAQ0mZ7WsZybGmFSWTN69xzLYYjsb108cAp
XRBglzQi7d2fvwB0q1Zyb4NTJc9vZWEynjvZmLlEmpS3G9kw0BGeeYsiHIe9ypDI
7vtKc4tAQF91JDDjVfx5SQM/JAyhLUoGVYctrZKDIs/Gb+bY7Y48oPIJwvgnMK7q
hAA6ZFOeuCuZQSoFvi3tVKfC6sTSYf8I47Z8IopImmRMSm5JlKWRkZIuPW5+jqN+
xm+CS1aYK2Vd8pqvAihsHbYyB2TeFFVLU8YFDtH5riBrR1sJaZY9pmOKs2m9McFL
wyx/NdHM2JIWeSPs4Cmwu/3yE8bkvY33eGos/53xZl9rk6pj25qxeSA0iEp8cYlo
a6YCl2BBsLI8naDuP8Lo1trYIGW09KdYW5FxDnRpQAzwfwNXc5X0xlOmAy1ZbIuV
zA7OWfSuwi6jiW3Y4NWDAbHIcy/YZwucZ4Q+SqbRRYhJa+v2XSPl4U6E2/FQTUr1
FW7oGb9Hphj00vQ8tMOHv/mn5tISy8BwKbRIx/cpkgsMkGHh+AWZoa9aIYglDEwo
J40ewSodF5sVJDEp/YCjZqAiLFhBC9u6lbevQnrC14ecliWrz8hNAAAAZ4qwZ4Rw
TrGYiCoklcq/2BoGJrOBffUdS19xjHhB6Xcob8v/de9TKt6HCs/3+87PbZwbxnZH
wbX/fwf0dr34fYzuYH85Mi2zYhTfmEUol1t7z06IyGDJLFb9DJLj0yihn9BtjJZ+
5gZsgxRFbCHlECseilhxDZ0gNRnQyH87tUfxbvXMngZrwf0+W1m46k4uRiRoSb5n
qypcnjlUAXz2rQ1dfo1Dbbwo2Yy7EawxdZsUthvPF/Z37424V6VZAgLClw+353dl
M/ObGa7KSe34FuAzP7Agq+/BvUo/INPhfEbUimDJ1JNiRwG8IR/aOUxIzE1IBMyN
KVBUbBGdpF8qVYWe0GX91rOWZylBgjyQBU/MOWSDGK+DOU8zd0B+CJKA3/91j9aK
P1hceW9op7YlPD7LYlzpICqAUmvwnRFW5dIV4U1Aa8vyUX4/HyM0b1f4EXNAhQFz
ubOZoZgHwEuT7yB2iA9jFhDtfa8l+RHcXvbSEX90UekHUdmgn0du92QvKrvg6TJS
Etb4z7cXJvzZCsMkjVTUWq8S3ABN44Sq05yUAUzp2JKNcFATEaBr2vOzCEs2ndZD
zJ70DgpPezSf1B7KIILW9UFO73nvWIQlqdZwqqtcvZflsIAdzRCEzXnH0mdKWXoQ
blQ3K/mMKG6tmtzaYSlLroy0xEljz42Ryeff9HQB69+xEXaKyq4UtrdfZCffR60Y
m6tdKsnSvK5Z2lvq65PC+v0zLMQdixGT2YMx7c2rQGrig+Ge9aGNKgNcFsSkPBbe
cyrnt5ZMIXodRz7OLOF7uDHuERvdQ73XAk1DDxMLWNFEHAZLPEgxsxCY7mu5vQK4
IJW1jvsA1GyafKHFkGzQsdubql3YnUq389p+murb7XVb3mScRLNHHjFmHKA/Ljhw
Gy3qfkSt6IXXEsE9duvjChq83BxVjkW41YglRhoRsdpH8/gg4ml9zBciz54LPVJL
xMYNEUvTe8+G9Vo3lFbJJT0r89v/qH9gkjyeYokV37B1SiNyb/Kj/SdoceSmYDUU
w0oMHjNVriAgjD8kANSmb82zSe871DfXwTvh/WsJ4nL2PKaoZa05fxED0AKRTsjW
dPl8mHC0xS3vvyq0pafmP3qdHhJXgr+xnpf62VECSG4ewOKvABks+MywM4Qy4o4s
f2dUn3DNTdq6Zif+6D4pCk0o8s6nqQsJlFx3Bi25aqz1pyQ5cssG2TwqwOjomPdP
MpAtCtXWaQOFCiMpeIT4urdlPVp+RHYIw6Pdv9S5AglwtrmuMSLw3JvVt+nG++jX
JKnnH3S3qBcCQ0NQ2SJP2dYJbTieWsLmxXDMWt6GBh3q4gSCm96DG4odd/QoDihG
ifB7xFRSBT8CHp1lZhsJQg02wsFNu1q0Wm+ubRjhF0xusbsmz40FZcJRhs8ModuR
HlmVig5q7ymoLYD2WT9RTOrCC3dQTa9htCI0SBJlvwonNKk3pKKAZVy0/SHzrBA6
gS0ePBiSP5J1v7FC7h3YR6RQFCYhrQCtrlx9OOd9B8YflQiIR1qgXpPztp26+ABx
s20VqLaHbwiM9MaVosvCYA4cf2VAerMCFhsERVRqE+50nCgx1BtRYBmLVnkYls6U
RxYlbF2B7jMpBTduH2Il/vf9wuOhfOSPAA3mjRHONSU/CaBqXxm3YAkMEi86eu1E
wCCF2AQt7zFioEFs+jBs8Snqr9h7NuoOFJiXHSSvFvx1lQsw3B7+dRgw1FK0ecZV
lqIA2Ll/eZNEABT+4OIqtVZCsE6cscvpz/uquYvmvMyZw566ad4Db12pws9dze4w
3GsKWVl/+3+zBtAH+J6AZez5ju3kiTDiVNWO69gm6APKhUWF1FepojwA6CoRiZCT
NWltABX3tktOQug6cKrdVWYaxvrsvv7NzoUtsg65OYpWg6VqKYn4/AVkZGJHybyn
9Tnie0nxyUiz16wev3oWvJECSBiCQogkIuoCEWTMZQyb8XdB3b3ms/KZPGOS+guT
63x/1k09Ads9bD70BsLrEpeIYI78JSRoCO+lUzgPpFsX2VIm6kC63u4QSgM2jdYM
Rzy2S8dvhdrgF3q68t1HECEm9T+MmmzarmSVYJ7OmEhr/MNgk5aJAhvVtmwVK+j/
Nt+Qq9M15XT+HZHmgJgATuLOS51G4JlHROCshATm9/vaARUucFDtXhWPbFydHBjE
qiWtSE18r+BkW+yXbom2D6oCgdw8wrZdNPIhBRHP29hUh40HW6X1gt41wnEwgWd4
S61ixDHinRQjK6w7Oey6Rdwel+Iauu7alwRHcK1NenZxm88u+Iaf1KOX+wnjxWQr
qMgXXmrbp2bZuyThfZGPL/9i4M+u4fxkq6iq9Kn1J8/zyZD+rNvxYT/as7oKJe1s
Zc4rn09V7Em1xwj7SXuNhymGDkn+k04jdaVMqaN+B2tnqudRBmG20upabp/vl81D
csa2pFZMwTmHeZQ/WxkUQxelMcpH9e/zo7cnXpuC75jv11uQRGUFV3pa2ItXzZcM
cl4T72l5G7D4aViqYQUU2T3jr0mQGffXx/N8BJIgQROEXaDkJgzIANN/xE5hreap
X3bqGVfydmj8so6E0VBJv7dGSbAv6BTJZ5MBamA9B5VDbaGOvbTeIm5PQDkR/1Wv
p9Hr6L29XBxBgaCCwpyeAfPRrU9dpnlqB5ouPi/FvrsW/hXWxuY61nvmEZqvJ10P
r9mRkI1/PffLz6eDtf/dXnqYC4inpFnXi3b1P+l9Nt3vZNt6zv0cLbPJzBYo5mMC
clQhlnmuGUkGvUNA3ETxV7ZZhGSduDkxrrvVKiPCuwta35ZncwV+RBiZuhczpT++
woy32tpPO9VwkOI/KeUselUhEbctMfVRgm5bCFmZ1GGfro/7flhL1c2PK9CEXPCV
fk0WVfyGil4VQHOrm8MRsjgQkKpj26LeD2zwGQScV/2m6pUHTlao4kOauq2GHZRV
2H6AmSo7/tC2KkRYKZhtj4LxM1347FBIelYqeHo3dlIyr3wpb4BZ8EsBViJV1lm7
T8ArJd4Ev2laboIQJAJEcnst/0dLwmzrBb3v9orFUzZe0a/vewTq9bJSSqp/5sQR
2C7XS9kJ2Wev2xvc9aDQxd2kvgke/c20J6L3p0eR6oXAzREC8K4GDuvuM/7bgnky
0cipmHdMwMgDse9Ns9m0R/FwRdYJQhokeRSNgJ17hcM9JVsMzRx0S29hwNmSnY8J
M029dX91tCxrIECOiDEsGwffpw3BJ57UIdp7Afu5ee3preY9IG/6cIMsWEouAQE3
SbHJdaLp9x26E0NYM+wQ1SjK6SEb+NIXIiXYl7Qu0PRyWMLYEQf0DQrylt+Rz6wW
fbjNJoqBTvzwIZOC4YojbAfKuIn30dvMU1Ed8uvveAd1ix5yHh6/T3v9A1MfTlsl
Tw0MRdTtbBSXb2Q/G/x3JSYLzGrzcjNLuj10Tj9IG/CCLJb+K4q28EKdtm3015Sb
b8x07oW6AjnzFS4a1QLgpr7KIxdrj7Z0d0Z18zy00B85CShdCgjOCH+SlvcIQb1B
0T/4IjEDcHVHWA7zc6jEA/VIq+WUcWlKCFLV/jDHYmog1ic6NrOJyQa6I/rJkj1M
6xFzgw5OtBNtWejejcKu4TtHprFgMheSXF0l9Rg/VAW09lyBxTreG4SVtxNqRf0A
Z7ZMDY0DZXFDz0QP9elFW+s2k/i/6XZy9rvkNyTaluVVMEdsPrkZ10ImDs802z6R
CtI98tqLrqycvgkD3V2Hch/RaFB3/QyLcdPCW6BAoscG/ZJbasVid+2pm43RzhdS
jJaNOlx4L7Nen6HlEoJfmWx1wb57qQj0h/UGkOYl9YoqxH9TgdhwWToZsWO5ER3O
Il5mhDiuKN5kJ0Z8FC7y2B8/fEp1qiJq3+J6zAIIkgyZ2hqiv6Hs2ouFvHCAlKQB
IG9LlHiqhB0iLgraLf9K40932C7Id8C41FlxoBhIniLVZQeKuztjV7wYZvCQP26a
7EsbZE+b8cbhcYgQ9uVXdwFw7adywxT8Maj0IFGkzjrvW2RlVoWg5DLeMU9rbBkr
RwCnYzqxeiQkxBzt4jXIlNqzVWbkSUULlsYYu3RxUuVU8Yrw0lqzE3wrfA/jG1N+
aF7+exiUuJqMH2DTQbAMu/hcK+stkrAmwXjwBuDuRjV1KMG29BYit5hx/dDYA/So
URmBJ+az5TeZN5a43w1Zt6gRuvhgYoQDNerOygpt+CV5sX12Wk+g2XfjPfydjaiH
5WkvY00ouuY7mXWDeRrYJQoztXVQpTqhtFU5cECV5IgW3sGJXFbU4ZW/0MQwIA2u
bT1J7ebRNQExIeaQXh3e4azp1Qe3x3WG7emY9iNLg2CWOBlIqlD4BZUuwZO9baMx
otlNbm6+I8U/dHTBb/cb/+RHXrCFyt4nhkG57XcIhNYyAL7qMHgeMlbTuRacVStV
5uZezJkVsGzQ+gVow7vR4viR4luF+t8KW7/WPBD1gnkcJuDhJSNGjSQjhwbpASIt
x2WEIhT9vgTKfrUQmCa8pFUuk8zFKQwKsyW0Dnm8w7uCAOTbnUg6d7i+6avngQh2
9WQo99fUvlEeYiqI4fk0LYU3TbHm0WwMlg72bwFm/Gz4ZhbKNbpEvkpxJ4zAvda7
AMUb5DlCkM52fEWpQMyDjcWGjiYduyW9nYRCSbUKpSF/c/dHAaYbOBPnBFPuwlUI
Jd2G2AnEg45j0Nm92dwh5ZqLUY6dV58Vn4tjszOfoWOwKNSPZcF77Vb+kctnBah5
nEsHz1ZfY8Iew67zaNlisCtElWINv5nzhRTdNbIonfwSdAmH3vQEqhHm83mNMuP9
DtFdLkLy7Gvy5+7+KsZgj6buAvxdQgASAobZReVZYV+jw9S0q+t32hC7+/0ArRia
fG12MiF6xxkYdt9QeB+RZ1fedOfw7Krlnr4fAYWDA1fQOMzBxPinKcqkOmPKOsbe
q+xXvhnm2xLvj7GDDTlsjtswLCNKNKRoxYdnLEHAt5XxPGj0/YxFcS2+JEsL0QwT
F4H1RLLgMpO+j0E+8E1vzOnVzuGshsZWnD1zrMxNbwuVDhykz7iGwerCBWkDpM/R
fhYBCvifSThxhLx/2/2fbDcUr2eBrjZxzp4CudenCKje/0ZgWy47l8+Ydzv9v+9f
5io9IIpJIilrVJy3MBU0tPB6jUfvbAZmFX606uHBy7bbzimXW2l2I3H3iich+C92
aUILWA2EInWUr4u/EPdPG2AYhqjY3lRaIWTmB8Yr4SajsnwNmGsM/cqrHwt/hQnD
RcgPccOVN7hvOkbXdSE3pcbe5eMElin+3CipY8CJxaWCzOn/mXGFtSD6NZqYQXVX
CfTAM0OpKxZOpVfk+KYGfCeIH4ogYL9xsvT12/svC9UDkdOsXtIAW7s7kvLLX5qm
LJcPwJpOvQIDJtNU/NxHrvDWjI5j0x3o+uAEKFvuIqH6iJrLhkbdu3MClT0fZxEk
jB00NKgQ/q1rQ+/bGJQhs+9gFQlrcqNjdMAXRCqnUzFWJVShryb1HEm0c1Q+5Bgq
f3VOmZWzMVqycy5YvRURDhrLAaD0ppXO1CTMlaB5aaxgc6b3+zGvCgL5ovYSerjF
16VG7gLObJiN+Rk3H67XmRqumfYsltNp03mH376rpA4yogQx/hHXhP3cIqT73oMb
UTSnIu+2/24ByU7F9sbE3QpwWF6hMudftG7XN4J7Vm26/CXccG2Q8skyIbJVezSm
Z8jgIz0lVhgixX7QjaicfFmLn/bFd8LGbvGM80+N5dC1MH1NNxWBwu9BdCr7MrzC
qhRdeRXxEKuLBvFw67TfaRxTYe7DevYinmtPSKzhlt7wtl6DRJwPueKnACyKfjif
9/SqJfCJ2yFUs9bIalg559deQzgPSKxABXnjgjpeCtCn5Q7vCYmaVVHSq3Fyaz2H
V1HqNvM0XFj5ArwRn6sfsPfFNNM1z7i3pBf+j3rk8p0aWFBP/Fhcu+2mTrvkgMIe
PjTdMX74JaO08+mHPiu/1/LtgX/BBWnY1ER2dYK5dZ4ySmF/oLBYpJnEnV8gaGzc
UoygZ+s5A5+NXRvfatf/3f+cVgWJq7AVrSj75xat4PYlVvpJO9GpManRetCgB3z0
0IAfqm8gQkftV2YjP+89rRVbT4NyUeKB+y2heON5BLKG32WhKAMFVHgJEkouJTDN
t7U9GXTdgfHLWQHSS/NUPzVfDwL136Px22qTff1cmfXkmu880eAjD8gaJiXVrXur
zCrqQ4D2v0/LPEDtxXzXagx9sHRYi0E+jSDlacKah11U4alP/gOOqMktshYkr3vd
4gnIIV/RUwCtTFXmnaeAbWPLKG7kR/ghEw6eoO2qSWRhAgjp4YECQowYRpM0Yvxo
95Zx8VHVtTEjp3ClmD0stQIr7+JEHNDLTXqQvprhQqA9jsy4xylfNtFtH4n2i+Nc
Pcq1U3mCWQoZ9jGjxeAjNfnPApGVu1Dg7F4GvUjGG7T3HDoi+CbPhFePVCPtWD8t
+nJh5E6OP+OFXCjZ7Qty6fikm7W5gJ+ss30iLom0GHOsP1OUnNGw6lQNqTkKPtsO
1jy9eUA9vvsCh4dlrsd6mY2iY9mQSsJtVvsV4lcn4Y6coyPzPG5E4fq105Bx953C
8HwLNwK/dNnbel3c8FFVh7qZcGT1pCtA5XFFG83kQuKGVMir96w0NBpzI2E6gTXR
G3MlPOMEJzKlEpADiwDrrFm3JyJAdNynQ6pb2YCvDz2P5+1Cp9+TDCVMEqjPW+hf
4QszhZaJ71CVaRRZbubOVu4ta2TlR4wcZ4Glvt+7dQqVwZFrYwDUBGVb3yTL8nmG
gcb9vPzJ+DN+2+m24FbbZKJZbtWizNH+4NJHZl8X77Yd1hJBQkJ290HJxTxMttux
cKTkVkBaQh8jog5kB7uorqgKphmv1JWGJ+UhpCt1IpOjoJ/WjSNqVnlytET9tN9v
APlDGUEUralGXTsRhxTS/6e7WDe+UcB4WjylNH9rKFGg3bYBd0ZRW2xiAvKVqkCq
CaD3ha9PoLjr6dapCTHhHtElGX5GDpGno3p661D2/uHt4B17qrfVD04iNLA/Cn0R
l0LNAOBvmAgDotwSCbb317Ahr5bqP/yagijx1/h91mIf8NX9u2hsyJ348DAPmnZZ
fhGYZXcLIx9Q58Yaxr8HiD4mzdXHtcVGCkFrjHz4fR24IBPdiFaX2igvOz+mjeO/
jVzozrZm2T8bIEdt6gA2VhTevkleAbMdRNy+gsiq/9wfhXw1N2FFZhCjDlrM1SgO
n8906YIpUuSjOSJwN+aiqn08a27gVrQApuI1GTu1cA+guPrbNzCZZ97uYN+BFVPj
kHpNCA1iPkU6qVzcUwyI/j8X4/z4NwNrYNV4HZcIYDE947bPHbwxyUkQxsPcWDfJ
SE5lxZLuScxc+0yjaG9sGBV0c91efNOzpWPh5Q6ceKq587wLzwSjYg5ERjIZXJLV
XjLPJd9V/ZFTDnN3lFp91l1oUlxTtQkhYrJJiqC9vjTvU2WMnrCbuTkkGal8t2B0
f2jEf1vVA5ky61XKZOk+1ltUzmHgY59qzxz1a/g0Hmhni8GSg5qqgjjOH18FmrhI
HcJj27wnaXvnODVYJwk4Psv0Fo+LawYaUWRjhcNA9RWpTx/DVUg7U9YKhbNX2Lwm
gwNEFgiLGh2POLjp5zOkBXT79IqIAnui97D+MGh6cYyRqBDtqjheCfyA8V/TMz+e
T8dGzLAEvE/+rP33gkvLStsfAbVxloZTjHWSVNojASvyij2mdc0Uqb5unem5L3r6
uFX1oa7pp3jBIU6ep5VVjFvcdJ3ka0W0JhpIub6A+WcBAxb2Crf+/lxu0wzepa5y
6pIqkfAwH2plw3pzcJm9yb8isglPJfSikq8RpT1nG6T7hkBn3aQ9cutduQtzJ93O
pjsAYju/TMBMTy/NkKEYzD4H6uMzQFxcKKUX8Zm7nTM8G6ZeXFIzVpFLkre/X9zd
p6jbqRGQowEWrSVPq5OzwpdJ3gff6eHfVc6YlmQPTecNzGMwSgEaKV1r9WW2kSR0
DpdAE8obJStEEgq9Gswi6obrSlIGbUBOowyoSNGrksroK2J+ULrHv09CRQicDgVO
Qy6jVgXTvwmbRcPBZSALXxN+K+5zTRdcZEvmdLOQlHqzI87ib1pJC7976wJpx5bv
xCOayzuPsC6IXg8L/oCip45Hy6S9agP8p4oyKSzTjik=
`pragma protect end_protected
