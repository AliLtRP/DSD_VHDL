// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:20 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
b0phjOxU6fGYr7C5vQnMFlzYlC6v2dD5pfo7D0REw+o8LRQ8iAngVWCEL8Is8/mv
AApo6co2JaxU4yKN7+aSuBKHXGkkoLRGVZeJhfzPcfKAeTE0cTy4spQLzBMvXDpg
ps1Rnza2yoYkv33PowuJJt9vNB/lEJXwMcQwR13oiC4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22832)
zp3Pvq4oXYhQ2Jh/KCAMP5vtw+prAwwStfaMnHc6SR1huZBLrhlAK0zvyGH6uU1l
h2bkk1txiSG0K18SYbu6iPy7Vcvc/NJryZLk2c54VjUx5YC/4KENgS/Xpsc0zx5+
6MC9WZ3EP8Q8kTI6louwf67ptUX8RJNKsjYWKKTAXhS7uLnf1Cn0vq6tgi6voPt1
6D7HFxK15SDSqfAemT8AqMpWNnQPRX3KATWjCLwIre8uRqytk7TlHan1vtBGEBOz
JQJxCQTOMm7V/Ig3VyTnFYlWFQ17yxkZTmi44u7jgoer5feS/a0zerg02MiCQko7
YoW33KiERQ79ILXvHcsI5ksHqOzhwITtJUu7/Q6vagDfuds2270wCpqN2g4QpZ6i
Ad6LOFNwrmJpQ0cXyaarIztwc5xoekXuemgoYDUCB+Bj/g/vn4Fge7zeRqnnq+dh
Ux8SIko+TyPoBdr5SNSV5rSA1ERQf9RPsOBwAN9p70bEgH/6AGbobv1c7c/GlhJd
9kNesEPwqouU+TYPOz/szwOWTA7yITRm419diSQkFaFgU/gL5Vi76P/rvr1bTJcb
wJb33oFkMhf6QytsBZoH4BvS707DTAteIjyQWxKcFeJ4Epe1OKSrwZ0ICBGAd2V3
lDvIdHsBlDirogWWQ3Mh0YkQmYTpqAutyCP9XsgLln95P5CRneti34K1osuvTe7W
XnH2Srd3S0RjQOtHzf1mzM5JPPMUTpsyOn8Fz4ohq6oDZFil/7FGVXYT9M9lp32m
G3b1vfaBB60g8YKCqUoI3SNNK0duxja4Q5Mk0KNWDa/N0oQAMZUHqpWOailcQQM/
a7x9YuGbod3vEcxycTJ6LqQICQ5tYvgqJQVktPx6tvW8gpXayv8cFBSCCYpEgz9E
ZKEMQHZc6V1zbOrdggsb3LeY27In0wVWbFHnlZu2+7OX6PTNc1rrLo6Y0adctP6W
b9OwyO268L5DtBbjoVPskimioTMIorSMy9gt5dvJM7E8dsQr9QsgOwp8zaqLHuM1
4BMKLBGAjt7sn2RzjeEt/8dJJLgPlVtRu34ItcsaxEuqA17yjOwgkucIldq6ZLz7
nEMjKP89rLML0JDMlBjFJwgj/u4Ps2UzK955nXQHhkTg8gAnWW0T1VOq3jZeSzj0
1gHG/OeVSD/u1DgZOF6HJ66VZzLr2rGal/QJCkVVKPHK2T08+d1cvHD4n6wqDB7x
IOiTbhbManL7ojuFYst7V3VUL1ZHf4M7eoq0UQHUQc3PY2yiX0r3A9gApboOAKAE
iZLqFqLPijS4K1RXwK4srqlq04qeA+Y0ojVWaxVKhxTe9wCIzpUj5FJ2u8oZAmZq
W0blVOPy8tMsbQlYa0omhpc2oN4sg9pqNEIkpvdef/fD0oOAo2nD4Q3kg6ZJRiTK
ro9sFGGkyzQSTLihmM2UUZV82xWbxzCYCpn5Jk7TTU2ZrRYyZ7JbcmLbGdGd8jcZ
vckh0n7C6BwFpraQRgtmmyNdHBOqNNXBbolTL6Z9L5ilq0hhjM715IRbmolXieVA
1lpBGjhRjpQJGjhUI362lC2mwGMynqauXatgQV2dTbiD8F/5Flfbxt4GojezBA7a
jYIluAaidOia9oLG2ea1JgNBezKAWeWhgq/pdJnIxRkS/Ii83o3h83Sh0w4QDic/
xi3J3Wp5tPfI6+B4Kszklkd8scjZWmc6rF2+qYLL/tI6iJkJPa88T221vQEc/B68
S2J+3/Gua2c6Ne/LGN5mBeYEQHEQ/EZwNINL2hrTcPfSfN3EV6WcR00GQjgkRC3p
sZZuQHLJbS3b7V4poGcB2dLV0dhnAiQFHTj+P8eD5DzEfHw/CLJIRmzHqEx3ueeu
6zTinHQoXwzMnVgeoKIJWCWzKZyZICli59krPEmbC7Dh6UAX2wuDUwyEiCWDiGZI
4P2/89ZMWIps5EiRpKeoPpfU1uRQIuOeUpxCppQz3i7s829FfOzqC9iXuJwTLj+1
F/eRMo7QhvRSHZfCktK9sFJw2/l8MpU2yeRFtwtGA6PZQm3Jnmr2hIKs8BS2eJ3p
NN+WXL3IdQPalVsXib6I9MDRAJ13aQxNJyqaMXmAtj6clXIGs1p7hzbmHdSSn4Mz
80tq5F8jt5B/hRTl47iMmyQ9KREeOw7Dyu7+rzIaBSeWs2KIKfktTrw46pcVRryy
L0xSYdCRgvb3rA0HRpZoF+9f0gvQstFbLh3lOCcx2WGCCVBju+FBkTG/k/TDeS3e
GL5X3mUdv7s4h2xBR2j8rgdyfIjkcu1GFFwm/C8jtg1+UzDILcWQKlR/pzElxn9P
k9HMs+KR4xJC+DGMaX+Keuk1cQ7bxG8g3DV8RtQNVm2WN53g2a307AtkY5No4eOA
eFYvZkgHN50p3ZDz1hp/wv5IgKsEtfoZhZ0mt9CQGQv7cO1ws9zqLHWHFMLOdtqg
tbdITXHWZUM+tSH4kVtTRQqAE+Wp0knQzKTkUmJ3uldpHZBYnEDqpGPlFRW+P+hS
m1pmagltMHzDC19vzu94lamEqEwjbHqfVZeO7IGkzIA0KuD5vZJavOOGgcuWB0nF
OYNP/gFQqjUQZs99DhAE8rOSQTWCXuXV3l0+BOf4pSWlqzc7oxngNQRCmbGZuU9q
pHR8hVRmczOZp/8FdHMP0aTcztVZzPIl/06IveeyrwI3gNcdfGae9LFLkKGpv9Kr
Ba52nQDljIE82EOulqF9LcgtzMGTXJ7p4VaVT2eoEqoCxI5ujgj1sEz/ZipZSu/M
1gdXLeV13TW7qNabDPETPuplZgaO2ZBDnx5Hs6CziSdyebsZuC2syZf1nVizA65z
kIPDMsgGkbaC0oBCYSyjRgxlzrCAodEzP0hiaK3KO563D/eiXc1nmdeIlt2zNDAM
CPe57KM7J5AcyU99VDNDTNGZx94MnTHuqgWaaA2usNlP0plz0VstTysCDQrws9du
dfQ0y8MwGAIwFQ0yDisExELKmcieiFvJUDBltOyeOcRQH7j0U9obZDl3d94ouYDw
VleoxHA7TFzlmlRA+Cf0c6VzbhPrIxdTbPPxfY5U2HanKfjWyq+ewCr56nC886aE
UBVbpCAeyk7MyBUZC4UgwasKNAGs0qXeFmLs+woNR0/NFC7cK3fr9tHctua9bEpB
vMQFHrDPlq8cumtW+vWvWkLkQReFjYoDPt+0CVabVMeGZY2CZKs88SMfTOpYMCFH
dyFsbp/J9NDSSDm+j3hPaf6ufxGZDNqkRPvNQQ2TplNLPxtZ+4k+T3U7Uv9cm+lX
lEtHQJFIE5ujY3F2AXkuIOjwlfViINYHXQyZDrHk0+ODeHJesj7XTmgb90xarTyK
lO08X6jViC7Xe0pj4nuv8zXPZ2f7y2qyQd0qB8oZeUp6arQXIOZ8E+d2Gc1NTGjk
4LnTuKqAbnA5u5nn5IYetYNvsYzhtTDZ+zDLU3tHEXMXOsF4MqyXy1HVpIb62V4a
GGghGiymm6MqhzzVG0D+JxjMG/1/wm8QT9tp+OgHfpnXWLzEwgkZBquN3WwDY3C3
UeyBVAsQS/cipI7fR44e8QcDpYyuAx5CAaavHX45rekbpPW/kX95/MOPziw4TACt
1i0IB1WE92nTRIGsdApROZo1W55dvonN8SRYWzHmIUnhJXWKTFzrGc0qKgr0XeNK
OSfGG4zxmCgooi7EzbjaM5eIYF3VCCebdFjXHqXx0NzMPo1IM/m6OpBAif+SIQnH
r61h09DwGrKuIDykQGGppqfpF7EWAJBQNOTvqzfmWhSu/PQRmxg3KyfEESYvRNMj
+TkV3idhBOdYDjtKcBhj37EB58HoRvX81TxabB/uiGyZNuOBarHYrIawUIT2s9SQ
PyJjtfeqCla6tjLFF6MgVWEoPtK8OJg7V+3u9jzzx/78UeLsbVHhfSIbf2b+W5R8
UtBvGVnfnFlDzDVKMdmH3zKUXZD1Qb/02eN8V3YyDTN4jYypCiA29jvro98WPT0w
At+TsFcxjFLdSIX48p0VzG9qkqaX0dJ5wVoYTEm6AK+Dzu0bRkkzm+Vc7xVUluG9
VRAlA6Zwlslv2akqamORPVRQSEYzg9Q0mT6UcN6aaAHt5Mf69Pcj/yNEWKuf+fyK
L8uxQr/8RppnbupGTH8mivTrR9tonsWcJHEjtil6tnPBi7yZ/jXfGdN2KczFTjoy
wGwP17lHwk0/wK4LRiU77m0NdnVGhT01Ca6VXrgHl43dr9Y9UqPi0iOhuavACq0N
0dyISfxIWq5EhcYAmeDH+nd6bj5NzgSDuGjSy0LUXnkqx646Gw2sOSReU5sTGnZM
0J+8/8hf+FhRKqYCxdkLIB7F8SmjUO9pd4gM20XUqUo3fQrDbAni+AnVWX7YrRKk
vHpTmtXcCKosdSKHmzA8NZU9KkxEI/94gZPw0B/mXmQPjj1jPQ8/0vZysgBB9w7v
MQkHQyhDiBB7FwO78Bs2spC8H/SGl1EV2oaO/ZRM6tO3zkE/c5gcOZrP6hCV0s6r
wdLApyNYwnCpjV3/12LjhTDzwqzyoKR7+RRGgS1jDSwlebMji0CaPzbc+iHEP6fK
j7UoHpJItJ35UdwIS/kVbye9pGMVr5OXSeQQsb75DeRtbVmMQIbI8NgeP1e+wfTs
ftT3IyLmco9+RZLa3pQrCogIgS/AfTym4dEyhsSlrhwAD/QZEGt4hH648cOWmgIl
QaK0vR8eFB1xx9qwRtUcSaXvVg9tqk5J2QrR6Bf8NrmLawWjseq3kVXvEqS3/7sV
n3fgaDBnsLzJN2colybUEuS6kqDQcclC+DCE5xb13sPxIC1mcsAQmLhBM489alDZ
ZBZdNsHVahIJOAJ26fswZeCwFyKjoWt49Yk6oSZkjCet25q5wPrP/yv5AxkyQSaw
DLOjF0GuF8oJX0j/3grXOIqSaqmRf3jBOF/w7AM55g2bE63LHZYfi+rliWP2VlJJ
dDhUziA/YRKWuc44vLhkQkaQbk/ic7ym2TeyOtfrt0Oam/6kPkjW0dYeQBbXUz2A
Q3x4dzNXjHCMNyYFyammWxt6rjC4oJndw4TAiR8klPUmM88A0xjrNHjtfy1NHdJQ
nNTc+kmQRB1vAFfKgfE1yzhT3YHhKieI4D50zhYPInTxTAIFgnCYeLgqvX2zUKbA
6sFOeJo3NiqVvT6vOGEhrg87zEZOsFJRBbvZfGnEt1giMRV+49BQifbRAmzewHYy
P0YR3siCIfdnPIr8dpRlGuROgRsz4YQTOKggQm5HfjGBYifVVxInjUPqKNey79OR
ObsogaSU1FgvbNX949OWvpOSEK6wREoAsG6i0XennHNcECyoFHAlj9WRfPWZQqD1
jPKdTyhF4uUuQ3K939UnOxglNQRttPC4kdHb7QNgHf02MBo5ISPlGsWT+Vc3l+qj
csNajkVgiCYI8HxFHQuIlvMxOJJba5JYD1mS7sjjn/UQFLsKKYSHhP+Mt7LGSblz
m5IhzA5+KXH8qq4Rf8k3qH0pb9detd4OgenjSik2XryueOlQKU78lSP2wVspGDj+
B3J46tZS3D8nm5Qq0toj3QOjBxBf8Vbp8jCg45vtZ/EgwLscFMB5I03LkeUyNUTg
DmFua+W8NIfu3NoyU+0+JjTI2/OBbKKSMQZmj2Q2bV0K2saS0gymXPrqNC3+BhoX
NeXUgJUPQDWw3NZRDWFduKwlfiDQNB0tOPdl2bDatmBWyK5D2FV6+oWpLeZfA6qV
bl1UWNMy43vcbSNQpLeTGL+dYjgNqhMXIsgetrmtsmHc3ve0iKOhK5lEl2dCDBzQ
zHrig84qVT0upsAV4wQI6D2Zeb+v9nL+1fnLczw2dmLOOnI3l1WckYM5qlOVu9ZW
xabAhG8ypZSljCTnmTxGWI/DkY9DV2KCxSpV0AQ6zfziqDQc7QyKtAHiitE8fzE0
j+2ppj/XZrYFsd7LW9PfOXPeaynHdW9z3rcK5VaTh7KqKgGXbQ3cSRHuPSXTxcSd
WfSswGi50lPAFYaDhysdn0g/aOCbzl5Q8er9Ktk9CYs0BaSeR1V9O6z7mCjQnQwI
g5ZCiBv5wRgy5LF6gOvQvYdJ6a820iP86MWrjNog+/QtI/nAm6wqTx/KIqYoAxO4
QbQTimPLbsCsiq27fG7dYPP2xsOgthkF98IJYGTR8hNR0pdLnj38VKq7AFspB7sK
6YBOlJ3r+PYTFF88xqwg89DCSVgpogOu4A/AhacpmCWLRYO8UTReB0e0Fr5fBtJV
QlhHtDSauvp85eq7w2gU6jj7pUkPCxjJVAG0xvuULi26LyFs81R4H/CjobqMjL9p
AfccXenKllTSOFaGBtorYFr23kMwl0//P8VVJ8MPFQzRYoxJlhiwDZxGdgUU8yMh
bFTiHPRX2SqosKSE3oLYdTPKHDszolO6OB6muDCaALBcxryslVs7qyeuMfFm4its
DOi/PeP1Na1FHow6Rznxg/ndzrbRblFCZVCYu67uUtcz2xAPl6yTSNDcTtRh3Fta
8t0jg25OpMiD4k1Bw8xX7nGELqcf73LsNN33x9x24h1GXDXH28CW0maJCSDXMRPW
mxLPmES45F2r73L3MTvlKOFY8FT7uZ5BHY7mAiyJSAiQ29UcsZOTzO7nMT/wUZDA
P+yixlf7qf5gyCmb/XBTjXGSDoH/kvYrHtdA1e78KvB/WcKsHNhjdsuBqElx0LBb
qp3ePJZ2zNI4CM6JNrYY9JwcKO7ArrphGoI8tsQIXDWG5LI2wWfMf1WOXsvlORP1
kk9hhtIIA4OlimJLb61ZNjM164OXLE5Z8Wt01+aByLs3ynD5OwlYxOGID9feYCaY
y2IcEfaLzt6CrW0XZQJ/XdBFnJcmLiF/L4Pk9ZX5da9Gyqb/yosI+2bNuACp+T2P
No3/BLaoPiXHr2ccAHzM3EUTPXdixaTFoXfMP13CQmbiTxFgNg5XKOucPp/4M5ET
AycxAO8FTWq/mS0BtOcKQ9IY0WdJfb0TgU4K/2nsctfh0VINEuEWTn7aX/2qURzn
GUzuUXOp8Ro7PxawCb4arUFm3h1Jv6W1sE+BKhVizWvoPJZ5wTTon2Ui4DSdwx9u
LIrcSnwj6yfOVTXYUutN3cSkT50pUicBJIfY4oxD/aJpuWyzKz0poJQpdI24Xow2
U9IcQ+jftcfcgohXVlGZuVbQSuC3SAWtTIMY7EbG9s8q9tXkd9B6rLXIEzKToHSg
+lxOKqPCQeh0pmpFj4QtOCUfl4JMQ/4eEVB0d9Oifcm/ngrUjZ9Q+R+kahOL48rQ
oMHqI0q+G8COpTVD8joOE4skYhdc6EH8mWHJSqRJnWwVPkSb5UdFeRQIogGbxBrU
elFqy2dW+KRESYbvv0/8qx3vqSbsavHiEHadwEBEvKNHBE/Bzep2sj82QKcVzTZn
iJcM3nFmn9wXVseOofg7uHqoFpOoX7axiZPjdx/q8/NztUtq0KXSGsI97ldkFg+J
eOIhsQT0hUWOZZDu8qdTdWkZuna7saGtA/kE60FrJSRDhp4fSsX9DdXAxSznYT8S
EdjweycT5ntaNUdqdju8JKJu0UlHHH+wYAjFho+PELrH9Ebap78WK+0C19TP253Q
lD3t78HC9mJmWSMJ3/cw07z5WKgrBlWyFMQROOrc5eEg/C5nJDKaLIb6+Rr2Rk/f
bVOXQI93WejRfOHND8Ex2oldqon4h76HKmYrhpGZLZCG+nsp6VlqNt2YSc0POVZY
cPP98l2aVjnaiDGNngbWG8sUvlDtedzNO6Mb22KUivcGeOLDErC6JEshAZTCHpNc
wIurmx1doyoE/9/z6aewca3JiNgbydqSDVVrtaO+4HAvJN/tn3VjaE6ehUPNnj+a
SkhtsLoCofW35p6gxMYwHYRs80d+ggCs/IssrVUb2qCYNci0pk3b3Bgbf5hzHvi+
uZQR6id0NRneUupG6BzqMHSQx1y3Q23A+kcfp8bNWT7WzrjAkX1jnyTBlcAhGeoD
8cOlKy9Ji42cee46sK+FIdjZ+bAPRmOksOYytVsobRukEWwaZ8vaGfd/p91Tw39y
4i5WGGYs/WCVrR8McAtfwVpmOSO5z32r2Oz/ZIA8P8bdESm53fhjBDFPB7hQ9kZq
qw2v27/SjHkeTUB2f8gPYv1XrJLknCAcsIUb/fW7eVclU/MxQazgmvTKyJ9M1Wdu
K4nGNoBOYjMxyrXkDutk5+q0tCWD1UkAgHiCA8FQE/QtMBvg9ZVsKJWy7zEvOwLP
W4NdHIfYyTasft7/be1W5parTY/E+qrOSunQsAkoWaESTmDf32ayMw8gXQqaRS31
5E9gKXRUDm5X5cHeAHozFji0LGzRx+8YLifFs7lrrWV1Tamgm2V1C8K4q3knGShy
wTNcCmekUhg7WPhR2kHqqHlVZX1shlygtjyXpCmafDWEEeeeMfZrv8WVBdslsCsQ
GMX8tUad+zX/MF8Hev5W8qgcvspd0hgObwzNy41g/wcA1Nod/+o1qysrEAE8EZ9U
e2xLArlAmud9D2gBmOMXrDQm71duoKcXls4jc+OVjhhCbBzwFDYE99MuYZZy9vT2
c0loXm49t6vd7hFYTjnDJq9EPeTl6vGhVzyHVTgV+750Hy2Xk7/zqFBZelcboSD5
QkNhJYfoGP78B3dfd2NGtf3zTAaW8JoHHA2Bo/2+53gnIfjlhmntKrmyWMJKGAVB
/+Y/R8reXhRMcQXlZ86JocwUVqkGSV3Nynbw0r1F7JAgsNTDbDuTE0d2lP9DjJje
24J0JBIGVGy41WB7F9h+H1ZeaPLWPHBhHV+ijhASFshQO5DGQq5qd2iWCxCpQljY
AXqvI5UB5dYfxsZTt0kPxFngEZKXFj58kUJbw1QwEXuB8N4zcvU7Eg20SMyS4T3K
wTug/Sh3ls6C8DXj9F5Q7BkNnZshAlYce3KwXuKVpWm/jnElCtrM2Th2Tnt6FJi5
NEOb6l6YIWCxma7gZiiavV6SozgXknCD5/yg/TwV3orZ52B82DuyqVx+xtrv9Kkf
EupJDNH6C5jGpvbB+xVssduchoYcH6NTYyM+y4ZL6byyqxQ4Vwqd8hyZrzjGm8tu
1XrOlZ1cwT0ykZNJ9A1Ph0poiY9QQjLkSVvVJVSbHxOuPk936M8Q8GEAYcCpPj3y
8/WIL0mAoHTRwWWtZcn6Re3SyEmUhMFJUzaOtdjcb2xG5WY+sLIZu7B5aq1DcPRd
fuh4i894NEdI8/T9BYpIYXPb+GwtoLAvCme0DXd4jUlcl+pUfqTSHp1AZrxov6CX
/Yxmdv8MPxK46ng3O/dyo5pLc4x6PZsDfsQCSYoq9HRKSWbpguIY1MEunef0Kli6
YJb5Ln0GX33tqs2JpcUZnaDEvof77JBA+Im6ViVOGlLt6+HrKP7rA2BL8PQcVATQ
ERlTBt6SAeez0FGE2yse1vBcooMqlqWq7KDxTKh1JgV4u3zK3Lj9eOcI+ZplnG06
gpSI4mqLM1Gz7ZNExZyfaMCunOIWSlDTzaw7btEJ3MusvoY+57B+uGPliPWDrqH/
3vXU+hK59eNm40PYIUoAFtZqq0NcIM3N4bZT8bqtgQp7TPvELdCaMzqRNbG4PbV5
FcG69Q5ko1t3EOLne5RT5DRFckbkbg1Mcy9Zu4M676Inr1QFweDU0RrBpEGHDhKl
LA0P1tKDhnUWafDHOCu6RtzTEwpTgA8iBYOPmwLz7LqOVW1sP1W3Mof+zMLPPqwK
jef/Z+HOseYx9i7WvIpugUD9UJOwTkqRVoHdZ5Woq8m0ND4+UECwQgwlYS1KlMMj
4Ln2w/DMflKX2x9wsXb43AGFfWRIFZ3NVMO6UTHpYtdMAXabnC3U5kWsSODP2iP9
aIXym9MbHq20Ciq4Rzj+XSKO6DNVS7Yyn/9ZO4FWLzAF1FTtLKY/dYTVjyoMdJmz
fQNzqjSv8Vfp+P8yQHqwrIkFKoCWWRrYacfHjY7aRxB8BrUuTwVOrSC5D8sLqLq+
FHmhi1AB9p7qXyGkRHDS54x8P14gHe/kr3JoFJ1uVklLsrvGdwzmmYg55sjrON7e
7AFfUqwDdXtUuCvjBUTTmPMvlK3mp9CC2b1oiPyBxrrfwmweF4ra69R84BsAsTsP
JvgZ1YJOEzCvmbjbY8vRQUrBcsLVGZT1PmJI+WVjoRUh5pfZGdUKbuGK1e67sRzc
242Bqch0tGWFrardZvT14C2n9cp7LggrxvlGIwtl4NAbK9vHgD79/ip4D8ob9eoC
7neYhfRoe1TyftQGvdU58CEIDB7f8ukq+afEuUJYhoDgJXko2BlvxathChNeym94
F72u4UsLHGP+CJqUiTgdNTpG+TUwVT+gLqNvt4lXfAGWKGbd1//bWqxboKGdQTPn
g9FmQe5Ns3wrIeAJLL88WBkeRFy/tNo4wZyIkIxjB6KCOcztIga4YnQiW+F1JUHO
doAJqx3VdtWxmOaLk5ho4v/5/LfN/ZsbRJ2MeOu0iv4LBdWazhd7Ih6z6kspAN7E
WtWEJQoj/dsQTWcNxUf63xwatVOeR4qnrG2FsnNsMWWip7ugyMjPNurzPTGnmFrI
k1RRe99b5wUhSqKsgDDtdafn7K1sf6cWjiZC0MGUaTXR6i32zXp4Td6ayGNhjMy9
OKyGCTJDJjf6QzDAgM0zlBrvhd+OPNJwEMMVEL8De1m+OhncTLobgM9pLZ6uHMql
e/Ixa7uNCAYOBGp/kEwlWA0W70I9tjpE4xO9l5a6QryZn/r6yfAKRxQY9kgQB91l
yjdJp9we7ELjAeo/WzRMgVO35xV1W21P6EOI6bsdLLK56RlR9HCoA1wsulEUxbYj
g2zMEFaMN6wWG96jJgLUNlsTOcJyuRR65kapnLVsyiclDnoOZKxdNwwIfV+dybMM
BXBpDIE0KNN1yZlwnU3OGryn80OFaAM5mKwxBH8d5/dIUEP6HhoDEka9UgMwpTbQ
pBTuALDn1yX00oMsOWusCng3db5FN4t756z+Nun4xkpog9ehkokBANnKWXls/nB/
Nt/lcW4efeg9YMXoFkgPDcJNTXVCqVFNq1mBkazhUNnNM+gGmrNeai5tXo1VHv5A
VCW2BVMVw2GeJEBJoSizLLFC/YkZO8cx4oKFByXsaCTF/G4HBSp7huX9KNRxEIbd
xp4i5bW58cTKzfgo8h1Gxvj9/WjN+LKBBEsS86bVM5iBm/pUQC4MyeSrGPHWzw02
8FZiYDbhtihWU/Z5zEKkjOFmD9zCxrY+KyEMbJ39x4iOzxRzoeLnkrRD7CXEbVQr
0iQsvDbaprUJa55fkMSWuTEqhZDKQNPZxpfclIfJsat7zSFgsbhQ4cClWzDc7lTu
lJsif23tXobfbIu+9VbG42EbIc+JjZO0AZomqrLN99tfAG/c5WAtMaB/vogV2wEq
RzpMgIEc7TkafEsOg/lK2lJTu22NffKytLl6FFd6pW4tofgFUp8B0DRoNQTxXOVC
U95i/fSyfGIqOwtcSnbjpW6WCFXHcjoWcHku2yuJp/3JPHbYiUxR4dNCoFORtiet
F3Nl6cD/jKT4Ya3e7Fy991r55vUveN21etWsQBQGj1fPKmvllRtLXtB0eY6vF5zD
+iG3WURIMHrCkAHAUsNqaQ4rZFNFoPTgwLziV7r1GdnktPu3hWvWCzmBa+hOpE9D
pah0TzP1H+g35QQxNHvOZS3zA22MDYI8GmdZXBee2btK6QEvDB6SiN/4Xs94F0yz
A3ImzX7DzOurhG+ZIlHZUICJjUsts14ZKyL36FC2Q1zRdcEd4sCHi14/7Dd3Fiym
P0ikr17JAvne44B30SVepFPSuY5oZDjvv7sHNk95spO1KKtbrV9nDDMH7buVMR18
XRfTcm/3Mse1O+CB44YlYdY98yWi+T3aBY+6Yx3eenH9krCZor2K05jglX4gXEe/
6Y9FokaH/a/mRJFuz76h02v5YJKD63ZRjDwTmjVs3Q8wIaaWOmwzf6AaJhm3Pt6d
NLaKElUWl/OJaKC+PeDi7LMkKL97dy06v1q2soX822LAd8/1Gh9rDma8TylnTA90
apM03+BimLckMR33mOkt8oo1dKSMQ+TYNZIRTgLCuRRyGoi8rDe44a7d5GLKCnHM
iZRHe48N3pMF4bj1aqx0YEhIITMEAl8la2KG8qtEi+BXrbPTP4SzlD4SNQA+eVdx
+VV06dn+hijAuXCDSne1lKahaVNB+4W1LFZZmBondFhqv4i00ta/d7bl6tqmn/A1
HgfHvv9K6549Yz2BQpKWUJTmQ6yC5fhm+Thbq3Pf5djNlpiVqjCJha2L/XSgW/Vi
yKAZ7JdBEzz4OchMasIHPOlxE/BUHbirteIqZrfjhz9i8XID2EOmGLpFY/SInNJj
ip7t4xhhny1O4P3FW4ouMKpOstlqNOR+SiI4ysMmACJP1p92prxfdrKG9N161EH2
Ec/7/m9aHc7t5E24Jbnmn5dGdCc5AEFOTx37Z6MjPUOJy/GJQzZVkgd6RGFrzKEC
xV3bJhzOW+nxpeXeDeBs/o5B7ZqnjPlDzQ0MkyLgUyZCf+vKwyBbMpzaOBM03lGI
NQutFd7UGVTVbSy4aW0uZwl4zdO5LoZyH2QPLk8dpXTBPwkiGkXHHe5Kj4etC08H
UfT7xdeIXPPg0gvkoSzGAFD8FaJkNBrt0V7jdXXhn2+FCV4+7lgt0cZAfue0nSLp
oaRos6xEr/600pCLIiXXaHOXFGlQz38sNXwfT5jEtzN1swcSXeItLQP0ueAfNfn2
juYyzcR8bm5+h4KWEcNYeI826wSsnEPLCISULAme8H2ieAQuyRjWS6pU9BjX1Dup
+7N1SXVbg7h3oKJz/z5Gnuh5CKVEYEJphCMYV1qDrvJbjBCfywhV1jeAeBe0OZbA
cBES7cMhwFqg9VTodJOsQsgziv20Vvp5XoJ+Elswv43wuG4k1CAP4YVqNdlhlRUU
bJJoSPS1U8xwx2TkiJ7JMcFXH1Dc4gu2idqKoITL/o2tHayaVVUsaIHnFUgSYVJq
AcfmlIMskJljgL8WEXdeNMI1VoJRyatveLSsaTS6ul9KKRxUmi7Gq95lRKgVuG92
V2xWLWgAfUG5raukjQe2u3V4KPt8c8y96ReqI0axyl3kdtlPn1KgG5NUVJquayj0
s8NwCpAfuc64XyjdHuaz6uSbxcl7p6uEY9A6yXJDJvTWd216A53iByxyEY+WejVi
QXgHdjhPgYVUhoWY44ejGsITER2qQG0QbZLhTCpb8tJrPsd0EIc+5zSljMfWJrfn
5bHMUWH/DdeZpIcgPK1vFwvxMgx8klG74GC35vt/fZrsMi80EiTZM9bEB0N4eBoA
zrgEDUEX0W7WyB/aKjQ8zkMVB5n4Xwpv7LZY3Zn2MdnNxSShr65XXw+PCBZ5ZnqH
1AGOWLr8xuD+lVMB3SVzNMo2bKmTCN2DS8iVp3FHiDI5BrVWlVBLlaJYPuc47Yuk
6aJdMC7R9HbDaapISEIEwMhQu5KHc2TKHq4KSdNvYaCJIpUuEcgiOdmjngfsN5GM
14qh665gYUqi8KsdA1Xqo2Tckg2eDuG6IOIodB9VMd/bMp/tpe/+ZG5qFfT4Tn2z
Y1lImu6wQfd38i0jeslxaNeL0kdsJT6qlhWtyq2hO4/ryDcEYHYMbw0BERuRjYpq
Ur51mSsVs6S3WaNkkxcFcJOm+xZ1byHpJ6sZqujoT+CbVBa2+JzqYqneUxi5MnLX
wlCLdUTPS22QI/RHr6Dc6cQ7/HHlt27cvbbxVJ6PVyMxOtLazdTxy3arFGz4VP7t
OHwFjEL1P7k4aiDqMLGB6UUPO3GAWESDydfK4xK2vQUiNnSlzGGJnVglBy5O5OZ2
hDdpMiGXUWLzx+yEaE2ap1gx2DkkKtrdxDo0/a5UNVGJx/7UITvD83YYJCx/Vzh8
arUuk50e/sxV9Pa18UU/rIYGwVOf1sMlE/SWIqq43wiG8ZBAj9p2dTGdp+EvoeF0
j9muxXc3K7MgyfHH1/Dr1wcTZRuDenNYusTfjiyOrKzxV3BFlW4VVclpPBheY+cm
MiY2Wq7DL8GClSqokkE+yJ9vzA9r0uHFgkxZMF9KZyMCjtzBQdtsIxbjp+N+m+/H
zHBGefRLPKlgg8Wkfi+uwTcKixajrU670z9mAKb0oFNBBGzF1h9Cp2juv6NdNnYG
aYdEKsoFDYnYiEDRPVQdzUSRLKBRbvzNXzzqSsPj+yOn/hk4e+p1OrTqhW5bMzg2
EKEmoeMou3KmodRffB6HEB5j9OdtwoiA/CnhlmMLBQWbgQWaP0F56pfHHVtLdtn4
Ze3GFeWufRWRNgs4L8yqrRNUlpdTFOdlhS2fUO7yTZEVLY8fjk6vXNwdSiKjj3MY
iyWcOyA230jxZN3VUPag+Qz4AVBvGAZs9iuTaEYQTWB8sA3OcmdXNx/CVJIuiHEH
9MAMoUdpUVLP3vNCyJrNOD/BHksC+SItt9UVZGyZWriPf9Ppd2qTKSIGr5pzmsoe
z0ZxzkZPQOzuu3f9FJjNPyTfibnSVpNSGRsLH+14cPwro2UkMkQyynZ08ZW6Sq75
nOoUqVWuShiP1q+VxzqOvnwpKc8r9gBEfyhmg6dDlXOOLMjbldo8iSHPRIYhkg7P
us71+WGXdEbEbdZfE7O2P5KHY+pay//4RrNWWBLzPfRNNLcb5Nb2pTTAft+F8K7f
IzlZtObpQJlE/fP3xquEjsmESpp+BQuRddYK0ghX0S6QhukfVVyWdeSjVzc7weI8
1E+npReAxlB9rkH9kk2xC1jDJLIgz6jK4xH94WJ7ycNqCQf/9c1PAEpLZYg6yZ8c
dMYBMZwWlCHVVPWVrcBAWdtxJ64fl5hy+FUzBx7kncyaoqKBSn1QeC1eC9OAmu7s
liACRhm+k5P4fzAyApAO+InSEJAsmdTuWZiaqCv1gOzvWDslspnsXETonqLw8Tq+
yyfMOAEqDikI0VJk7+7qjl93hvmGFESQDQwAiVnSj4YUbHL0rFJyl04YyGCsUFMe
oYo0nrw2sMCr0f9wCrisfRSc6FU8x8K0tA0xJr/lg2bc4fWNEhHTMcv6W3GcWVkH
bviQrfhHk6x1MyxgiG7lUwprGa1zDqO3SHeNt0axAMOexdsuMcklh2Qonp2CqnyM
ujwnIgn18iRtp387FXABUoUwOYaVe+FQx/BUlHEPpix1Swh6RNX4G93mgaqB0H2l
Pge1zGRnCkd682Qid2PHoGhZ0u3BKqzZb2GurMmVd54XbPzrqb/E3ADTkRUx8wxV
udZiMKXRzMc1RRIA73buBVCMPJ7D2Wt/n7GbY79v/hhsti82dlRCkHRu/uDuhh0p
F5yYqOhJZpopjji/C8SnJM2MskaZG/7LVDfJ2G3isUqq40wAAs9GPejNvAJS9MGg
jwi0YHuaigcVfIR9x9AyPwDw/EM/+K5/S6gd5TJdtq1EOspQEE/rd6PGZJRVfvsm
vtPnkzyvuIUcFRqTcA0IjjOGscVyQvDLoyi2h5wD7Qqq2EP9RM2Z0o4e15RebpGA
RI02Amomw/T4sNHJMXt6t4S+o5tgcfke8ri5i/7W1zUIxx8/HGLgoiekY/p9VgbC
y3oWYOmwcqdVdV2k7zNoCEGJL0mjC4aApABZQUIX2YwnK7qCE+F3XkyyfwY19zOU
r/MUN/T9CPzMDmTUU4TqaGiKJr3Liv6iXeLYGVdU1K1KNC5eFAl/OR7lwIqOYHFE
jL876tnOdDeZvKqMWBArsdGr02bOwitGE6lDs7rMVxse8rLzSBoUv70zjO2bR/mz
HQ4Og+gm2vVzV89gDc6nH90u4FHo/Q8GZT/oI5S3tOZfR6Wf03roaj5+5DLvA18m
82hP7jr/CmQD0nJq0xP3YK7TNkBI7K1L4w7FSt6WmoMdquNQsCXFeyE+cN6P8YCz
4fjJyA1x+R8xw1Cx4ovmxTdQ3qtQ891mS3LCgLsMrFQb9qYeIvNNzYursiRxLNm1
axsHVnpMUlLA/zgk0grAe8oM1KQ5M+fx+wtsHf+jRyXUfo4/OmIgXPEe/X0dPYKN
mjb7k4C0yQKEs2ryRFZdzXZNHxPyevwUQbu5t5FdYMcRnQbJ1RaFCZyVzp15SY5W
0uiU5/JOVV7WkkH4H+lDZ+v0F2+yINea9WPUiFk2FmahGrIhEm8xe67aK5cM3xuV
ZLj+1eyTsr5Opwoztv/UDLlaaM1WqYcebwSBAWQsMFwbzEulvBVP3XQQFrk72i+i
8CJNTzxXD090aR79zbUEYQ+YPhegnuUAxZZDgui0xKPP2Med3H0JvRReFgswEXbw
g23czkYCWdjIUyx0jFSvNGsrB3y6ZUNzeg1diLfBnPd+/MjJJAguQBaS7vQpZanz
Gh3KgsDO4gBMoUgkmajNIP1WsomVzaAH7Fu45B5e7w8aN3y9BN0bPfN+i3hjLjcZ
9jQzUJmA2b+Yqq9isPPcsYlkr/IwIEICYPRLd3Y9BFBe63Iyj2tfUxddXNqIwWAT
GxI5gufW9svsmwq4MTntVueWhdmKsrdNr0O8uLm6IalHxxoPEmeQHJ4W+E6rJ9Mh
xDyqxBPWuB3xO7yhNi1at+Wn7zCO/lWoXjIl79Jdrmg33vCg9J1zJ7LC9jFNvOJm
/WJCjXTfypqWXZafZqW93ciHKpF1LZ+oTAOsEOZUBu3Wh4QXcWBlnLHqxJYw32Rn
JQFbTsz1rG5d9yaiA6xEjCxBCk5t11G1dK+jFsAO+Ix7AuVOEMO42mvRI5guN3Pt
wA/cg7mQtVT0fUy0B5WJZmTl0+cpqfU57Zv8wHWZWvvk5iBgGIDtJNsZsY2ff6vo
OakWAbvFwJYlOT7Agylb20txk33VtRLwDApK8lza7Rp0DkzZ8VzRluW7U7Oq8fsR
1fTJEpi0Oixu6YsdIKGafV7smuhr3nsYxqegUm8ELqOIM5tsZliIYt6JHJ9Q8i7S
7UpJkSkYqvcTF3aB5QtzhzgXUVeoGPTn3mquI452fow62PBdvtmW1ps7SsAZv91m
yoNOmyOFOUhSih824xUDhYQiOUoofiwnrb0XqoVpWDs39Hlg8trYLTfvAJQWVGDk
teziDcNTwnLWQqhcLvYZhn5hBY5e4q+2YQ8Dtuh9BLodcxQfN68SLtsP303YVXzY
R/M32N7jEIAr4LaGKzKvHlY0Ucfe+C5QyFQhI189XLzISYJytaGBGjsOIINCBz6j
r345pCExgSLnNb3jbUbLN1v8zaGPceGyBJDpVK98MqDHWB1O21S1ePNCaX36r9LT
66zFc6rDydLiQcvFD5wZ2GvRNhVeaYXSu9J6yibkhPe5zEtBs0BTWTFBjjz81pAK
txHnP/HL/dJDRKM6qUGNySZTuyy+plgEwtcpaeM2USsr0bUULsrZ9XogsarYDIHW
4S2qeGijcObcgA4eGNwzHeF5xWzhOD4YmuklVq1htxkWR1U8MrXc85e+Jy4FXsJz
bo8A9CU0hBqNaZfWgLSnibifZAwDnGf88ffoAemuuNlGkT+X/jNZpoerkU66ky1A
2Aw3uhRknkLLoA6gRo6ImAY9QWlc0TCSUsOuUZ4N+TFUGRCuiNdfJJ1PSKCUMget
6NqfUhTp93TXjZnEg1ZrLfkxaf0BlX4kdjlFB2KuwTBZ8sZM5rAzrubgOo8aeevg
WtIRXac3TDvNn7YU1DEGBlFu3TKcGVLjS0EvAj8hS4ZBM+mghm03+nnP98i7L+t5
nIR/gKWNdevhR6F7s968pD7v3Py05O9jCOwoNRfjsqKnrv1ckag8Zp9NJn6hwamS
+DeckDdRrxvUA2dKwH7K2RzH7Jp0d5vq7dfAetRnxJd1xw4vxpFHcmHHLHPCXFp7
ff0VoX1Qb2Yb426+CPRmZE16Uq6yJuX9SLdo9IXqs64GhJPdnNxTJDUFk+gp1iWX
wDE6PWcNDgn3whjARXANIWpwRNrVHym8ioDx9V6sh8aDA+Yqbu8puQ3J25lUD8Jq
Q5zA/Kosh7tEZFR8+UXqf4ADwfyA90km0T07Sm3EQlhvNo6cyabydNLIAL8c4Tuh
kMygk0ma1W0V9GqfS1MNXkqZiXeEIL1REeDqcSy/tw5oJtEf3CKrkqqX6VKSfTtK
rM/a1ruU8BbZcD2eQRcoSJ6Qi+rJZW+jWz/9MjANcEc6TnwI8UzHdNA8GKo3bw+a
7gmsJWo7MCQhyHJEIAXvCdsE2WwctmDQimjqs3DEbuEq1DN5uALYhcspIs4LIv35
+ej1elStBcpxI4n1M8bNrtUaNtOLCJKjxpvadqgomxMk+ED1+dW+marb8IFZJzbY
4eNKkGpyl2KsAlxKA4nAjXXhvNDP4hqe31nnnXyJMOLuy/gsyt6Dzjlk9Vcmn/rM
osyoPsfQEq6HR0coYLYKgUQh+dMEZxxqEyvKexJEbdxsvdbGKii6VnCDk0yFqOPI
GRzIgwjvLBBirry8tGns1PWtsySH3kLcg7LrMnZKJy8/Yg8f3xc9yYNEfLeGid5+
uxnScOfKmE/Bpz8wL6ya4EqvPEeTgdrKOHdFAumjuqWaFDEC9JFOcJ8vUyXDLKf4
zRW/O4G/KcInp/fQl4iRzF4Z015G90TWPasi/pnmwXY1ehVhvyA1TvuldIrB+Ka+
FUDSpIcRBdcXSE7kOxwg9yVlQK5sB4WZRzukV0n4i7pNOZGMMFkcl5aOFZyai77U
EJTTaqhL9M019tW14M0+lnw8btUSLKCS8huVxb1GplVv4v3PwizUSsSx4aS+nH9e
W2Zm1OpIOnLluFOYZDUlGIPf9qFeQiENlwuXzEMLOGGo9mf0nHUyjizrbTmcFL4O
NX/0HMqtZ7bnc24fk+jEPf4LeJddgN8ti41lQX+7YTOuO1+HEeF19N+hiMhwNTys
dYOjRZ9bJQCMI4LcUmxdmzI0fKIK7CjKN7buAJ4kRO0py06SE0TFX6qxm1+MT6iF
dNZphSHw7Z9vcs1JtvQC/FRlYeh4l5C1L31M2uH/X1UHznAfzo7eCc+PHTReEQxa
bYf3/7I49LulUwDUlpTrijwJAtTH/1YwkciLpMcuNJOJl8AweZHf84pN4GjzYcwn
TQh6HmDFlOIeAv4Ys8C1mtrbJuergNuuJLZQ7/UyASa+ntL5K15zwyrhOVYjA4dX
Qx35CSClcYnCtfvD4B5jkgzSVYrSH3QMOZDThuEMwNyNF7YDfZxdh7HtB03Y/S+0
5t5ze5aJFKOz926IDHpYTA2mIHzdUsFkjRnGvF3suMC217cmS0X/pXOrG8Vmsp5+
Kb7Uiv3UmU4bnZeTMWQTK06u+s4N+35sdupp6GcQOb+3etpLdyMU9dxZEuG7+cJ3
nlLCiQO25UgK+LJ2o2hXq+g7xlaXuFZfZIMRJI/nBH3VH2h30ZPL/AYJQYknsxye
ubS+Kmu7p/+cPGgNlQOuCsLmQUIm+hOR+Ef+sP90xnj/I/suMc2grvo9cTFo978t
CEtwBMUGyP9QATLWuhC1PcM2WGN/waZAms9OS16veGiPVUitRbbk1azHHLWUNOhX
WX5uvSq1vAGCK+pCkWUBjKaaZXemGunIo44T3VU0BEn2vsSVvDNhfqcgLX+bPoBs
Z/IF5vHB2/TTWGWZRZt8vqmamu9eIsSdaot4v4gmBOmRALqIwwPegbZszAT5vkSz
AGbmdghusU2uOFqCH1NgLD5rAw0vg/U8WlPV0eeUPnJkelQlMaUt2OoqNl0lpZYg
cHrvCOXwdtdsest2/KC5hBClV1dfjQR1U1tuD26XYfi1KY3bzzorEoWLVxa1D+zU
wUA7Q5qnf8lfBBQDPWEcb0cduaU3j1kZyzzUM0+pzPDSRI37w9/kXk7KLQ3VSx90
vMo5Kn6SVLFb0yTSGfjN4+EoESR/TXC0TsZbphl6QYiesFB81XuQtwO8boZTWkbC
O09PrwzT/wCHXFFC/OM1y6AqXdQM18HNn4Ig7xVY1gXvy/MLIEcD5GS2dt2/2Y8z
ZmhKLuQ6y/P1r2QLQ31RWWI/BxrtJ0/cRZ9eGbZA4ZJWQftR5rRMQ1yXcZt8kYjf
8iUg7H4XKmyYbyEw1V6YdChIB79TzOIFO/RYmUm4BW74Khoa8uQ25jIPXHNw3GAT
Px+8s9+RZonrqqWb6T0W/MPnUgcWMl4Fg/hmtnTnM2KOr5cSI7bwDSIlm+wW9BUy
ACGPjCF8nUKDP8WOvaPmulnpizw4uVYu8yEPdMm36T4J5Kp32bnlr92QdvpmeBUO
tCTtBs0Kc1sBiLJuHKC815aVBHkl+OKO4nZBcTsMvHPAwPrHmbsMxnESUrDmv/Ma
l1toH9zO6vVHj4NUcAWsNYJXPYrbeZGer3xZVjP6dG0j0nc8qbojhvN8tSS42F/p
DReacXMzO4DRbyWddAr6RNqHECGK73CBYV5Lad2c+UVe2NAkLAGqVNC7LB+F7A64
YzQZwvW1eUi80uGyecQE72YgcJmb2KGcGENmFTBvOjav3kq1z4FjI8kxKcEir0i0
UcIS3wKr42rdSycl0o54jhlFZ3SvvPYlLoDUkhRnJ8qq8+0MSJpQCwSsrU+QirOy
crXwVSpJVFbPY6tBWS8U7F367tWPY1xZ7eCDvtvdUa3zDGjLg1cchAs01KiR6rmF
nVdwjWrNQlRFtCVCvnibdTqcoHmI0MpwknF4RgHIW6+dMaFCyJQx+cdV6HaU5vn6
nrGd5aMaVcbZ4qhMr3UKEzz7vv/rw64JlroN9ZfOr2PAFhXCHVg0guta5KMa6j4l
iyaKd09bI0HRLkWd6AALES5A90Oe8rO8ApdDfL38dutWARPbxk12S5LtOWbvFZxX
OOZOHGErKDldqO2XcUdYdEMw8fPUb6cXI9nmMe7BVRPbq8/jDFNm5GhxJR8mcF2n
A0byTwB/vp8MEeLDkovcebGRSGhDOZyA2EmTUavlXeis4nCdodi1TOyJuuDQOqSv
tKhQRI9iC5Jv2FChQDdrSQt9qxPVxCHXKhZe+lyPfrLmX3d4yPOS4ABut5OTFxz5
QsGHn1EDfkT6QwEeK3Ys5u2Er6r/eFS1nWW3tQgy3fzs0RQ/8Tgk1ft85ELC4PSu
cvWQ/fVK6BANDoz3hdOR5FSwRndO9vYrfwpIU6LpplwfmSRENK5vMn1yrbMe8q0k
8Z1jkhLu6hBHGRXym9lpG2S/J1JisFfbRbiF67ITBRj+3SlhZfR2Gkstc6N1BjwM
1ytJZpXcsl2yEWuHUOzVDSzAbpqWEjCunlvtGfEGYaggpLCVOWzEWpYTHUhTL5yP
Z4hMug3cBFiqg6QWQj6/CzrMZPCCVmV/pXGEdvwxgsybYAvjR1zeuD5KFjCqBuNz
j40Ks0Rl9RcF9iK3hHcpRI1y+QhHj1PZjew5wfcH5c876mORo/t+L4M6PzvFWK49
s4wQR+66+ggp2/mktzmcZ0MrnLm0c5NCfDtdnr2nUjOGNnxiAtR0Rp+xiLNs4Wvo
GyWO2YG7/gUTkt6/b9PYDbI2z0oV1zWP25cAnXnUcHtMeuIlYC725vlCKdqp6GR1
KiTomPXMCWil8ReQqjL6vkzV6Gs93PeYTzrYQ5JgxZFE2tAOYXmTGUUhdkTD9jIH
ZN3H465ml6BtAkZ7/oQfpGuwCAzwkJqfBNeg8F//J6382vXhgthDLxLquMMscb01
SfylcOHdv0mM70GgUqTdG4DAaOm/mQ7p6QpbPzJppfots7X3fayAaNEWi1mRAd/I
1XjbIRl8yB9ytXVsuBGaaVzKeBSVNJ9FE7lU1j/8lgOnbtltHpR9+TCof14ZGPMJ
3YlT8Y/mnx81GHm/DT6M+7B5vSvTb/M+uXAMpzLHhn78g0Iw5xr7PDty/fl72IvK
bqJO4h/4GkUtGXGsAeWcH9eDS1xQPdH0POwTY8uNi5/r7udAiHa3UMATdVzi98nz
Ge63omSxMj5wtcsWIGjqmw3nl+dd1ZLJ1DMI5OwPIo15sv4DiMgOFZACpd3EjMZY
vBkEwwR4D6lxzdE84yyAFqNPKnhNLKuTWDRSiXT0drKyBlBtVG/kWdodbneHOfuq
3FCBxGhp1U1kQ2CCfmXwcs3u0gET4ZNlwLGf7m6M9P0aT/nSP+HCd8hT35g6u7FJ
l5bk8PsIdKO2qZHCy0unIRje/kRhbJfrkumyukNU3vg+akf1hPx942fPx2lIfLyp
e6ou8aANZ2b4AeCbio6Rkammmcctdy1u3StpJYJMtX4t3+vte4EAakfihaqQat/S
W7pThqsqHLXyIjniKNKYBzUB2J6YTTZcqCyeoY5FDGF0QTN3FkrbiaMqphizKSAC
szP4QqKJ4n/Vh0z8PHt7enZWur8O1QojXqFh3SAtiGI4r27mG9Z3G+DEaBskgODn
Wmad/oaBYOdnnxOSa9Gmbp08qMrWtUc2cq6AOkwyK308xdXrIbGbQls8andxh6j5
sFdphZ+DKmu27srgydlWJiiPIj1/M5tFDC6qMXiJn/2pmptiRiMOCUjFptLuZPZM
mOlXABscYOITuXsWZf1gWU4XXw5oXS1KASf5M8vDszxmnEEFBQGDrishzSqavbxl
NWfa1qnqfGX9UJCdR0DuiuJrzvt3zuGU48/AZQs0zNuvFrg5gISQ8ps4lcBoqs7J
LLYdR+yf0rj0JqTAxfmgRr/PayDjEXz2NApk+yuStVjUpRW76rbWCwbU4ck+s8RX
mjTyTeROXanQb/n3tbQ6UhZ83oCUmxR0Zc5nhRJXuMWQ5PC0W01a5UfKAy12PtwH
SmcqoicaDcxDVOEkGLcKGIDZy19scTEJ5XC4Gg3lyD7VZN/oKuMTiy6LK/pK6SuI
frxhfDiP2jbdME+tSttpZlZm2M2sPC4pnlhfDwrkFCeNUXyfXgJQTgYoF6GHiMwQ
gyt6nqD5cHqmlawS5B7A4W5qncrPqyoWtuLuBG4oedo1a1YRJ8LxAGrM5CL8V2CZ
fAXwYsZhrg5NcyJz85LUYMAb4a6hrGipXO0zX5SLWEIfrJDHvbDKc2a4RfyQAozE
WdoN8s2vxGM/R6CdGOhPkEOu/iR5PnD38oROePrL/YJa8LAceT8OwK0X3fB90KuO
j8cQ08FVD6DuzRK0YYqIPpefYl21svocHUmPSbvDBl7h8TCucvyqRcObwD36KHdC
5AU/XxJvQpBoY7joh5DQCcQAdq+0TXgyVRmKh9GDU7bSDnTOFJwoobqPsmmUsqRy
qTG+xcup9DbfggmFfoqyI2bhfZXc9t/eWmHkySYefNUfm2G04eWDV3IAdFXNx27P
9F/jg2kdbApLYHtKxjO7pW8oAUsW7tPKbhlZKk5TnQraIvSnlbvHIJU1xJ9+syhb
HkOzBRG2o0rXK49OInfG/SpGXO1q9/Jo8fVVbc8Fwg4EtNCDsob7GmdYYWvNDbFJ
kp2lMtAAaify6eA9H6rSR0sg+RbnBUtV0gAIFMqgcINLDcdAmPEsMo+gRGsuVYt3
bpeXNg3w+NN4WP2MfXmelywOHFu5zoLKlj2+r7eVvArfbqxW3Ic06F+L3MNqtvU0
sxoUdetmY/VLTa+6YWPdIe+9m2grt3nDxnvNqR6jDUrIwr0s5hk0C0vxJvLhf8Sd
K6Kc+8oBjlY6EDbSMUMBHsy9NjueRU2/eJsXF0IKwmEgAs9vfS4zmNi5+Vnvdbq5
4a8EIlxhRN2t8BS8QU6Z/yITpwFlCCMbifJyUiaX5EXpXN+9IXapXfYIkYYME8h7
cd7vfhpNS/6u5nem7keBmfdnP5QP6AdQjgSeb23GFrCf/JjhYtx4waLH1hL4NrAX
K3pgARi8t0UPhO1Mjz4Yng/M6Gu+Xw/aCX/gvgN0ZQXvUedZssybNeYrjiquECK+
WltwzD5doRQB0suMPaLmP7IY0Rs0n5pSupqydi1DSPfftMWp+P/TBa4Rt2wUYkoE
j3Nz3S0/CKZ16UWRRbwyIQgYaNzh0T7MzzGofHnj/OwLhOjzeI0zGGmtJpKVDM7x
pnYO0d7VQU1PUPSf6ZvBgOV5mqqWkLz2NEFkUnFzt3VOy2OOZ0T7Fn2SObV6AFQe
1fJv160n55kIdH/Vdno29pumc3C2FHFNEj06YdbxUEH1udYPZYGepecFp0blc/8t
pqMRTNQy3WeXAfIrKxWVXf7BClYfmQamN1XdqSdhnXTQH4eUr2bEDmadF5f4losW
p6DOetivbVajeFvKi3IseM5RZBIpE0YWfW599Je+f5JIHzqdgg5WA3qvO8aecJPv
C4KVnFudQ6NeYiE0WhD2N6h53356dLnRXiAKFyZQqaBdDFAz1ctK4ixQ9hOapcwN
Zmj16YcurxqVwE03xHQeU5xY3/ql+RVI3tdnx4xlU2cXGGRt0MR2q2B5/IBTW5b8
z5HMU7Xf9VF0LrAQS6A8le1i7PpedmRLEWdSMprA28V64MYaT/sUgqhAx9/Fb3L9
S3zzeEA/rWfpcK2rpC/AMKx4recPCxkREcSo8e3SWkxjgdJ7mf7Yjm4gS+NJGg6H
5HJ/O6NrLu54EvAIpGx97oe8iDln0crWmbw5tG3fMAi3OrtkKzt6WYHFhzB75Mmq
CUP+b6pbbcm37JJ6nIcay5m0z2PBVVHUEdW9abb/uEoDQ0K9S+1C3QpVapALFihy
XQs68Zeaa1KIP1pNsyQOwHmPmtNN/4y9/0bXj6uUFbdrxM/fyNEHhWsrL1qvWx4p
vffY7qcMZ98Hq/iHrzVzCNxP6MMQklw3aVu82hVZnVluD9NM3Jr2jX2kVE8fLaWS
AvypHFVpJ2fMFj+Mvy4smFakYFQX+YDZzEvK52hLBmRuf3OWy2354UwEzyOPPHtZ
/pWDB2xr4smzDOw/S3LaHmueu/4BUQucIfxMcSHaB3sypP9M5syDpDirnyKAvZSC
laZk2GlcupGQjRTuJkn50PRGizrcFfaas9pcObuZlhZCZ5dhHVVh5y//PzThRaQ8
5QL7Bzybc6a6TibIsSVPteupQnbmM3ZJJqcIn/NPuLnEmSxJLPtU7COjRDFMZbtG
8dLHSOxGrEgHznpe2dL6JBghzkmqIanPldBKp2hwseC52++Rvzfw2aC8HcX7t892
mvhM7Ui1oPvPyH010p7XJJXJdTVXyjthLloNpsFkQyGYRVBCLZSSwVkFnOv2O7k/
yij2v7CNfI4lIjrsL3Tv9fl6cJgiDj2vRdZWiyTSrzPNNl2/lL8VxRdYkBjBMeEA
okC0edLDv8bM+8J5ChS05g087DYFxVL6Xw+ZeVflFbZo6J+tl98gi905/1na7td0
Lss5LtEwkWt/rx3w0xzaIcH+ljavuXMa/x+bFCAaJ1KkahX/YNnlfGbalrFjF+Cc
zKScQ97bHw9w7n590GnDxdjIcPAcgK6PBxRdbI5mHuhnuftbvT+wcE3PswuZ4wqj
aJcguYCFdiNe4G5R6gU+ck0N0FJcoKxaVTwcONJo8HsCWMTtMJMK6/vHbLa7dbDs
b8KUMN2zQ/1xdSo03PqI0Li7QOee5oWlx1/4TFOazfgrBctLLgx0r+SmIUEySb7o
kCcOnKaMspghM6y4BAkO8H+MUd0cO9Je6dMPjAgeq+wDV7IxRUm4HMw/hFE9WJqD
V/pk+JB8/Xcv+PW/5J9lJgPnoonw/toG3+vu4p+mDVy5FXTVwGF0PF+2iTS077Ou
PJlEPxPjgq0gzlJBoTixETRJl7Vd/Rdk7saAc4RssMO/UUUwjdkm5uwYCJb8cUme
xxBeg6inFdW2asmmM5YxnEuMT6Bi0hmHoaU+hht8egTh6nQp5P9b7iGykdQx6E2A
DMrwd6YRCQNOlmhqtPc39WFu9keWhFGEVFDtLzdgMKOcuaykXJ8pZ+2hMuDqyaP4
zvL/ZG8QojHv4CLOBpViR+u6UG3TGS9i/NwXPyoMhwPd33q3KEZqUB/9s7bhMZik
ZlsnkXfmRObqnrjOfVYdywA+RuanqZu7eRaZJDuBhaJys4op/rs5/KPASRvHEc0j
NCgC3Jxx6o5HJkIrKB3aDTtBXPO69O2AxBBSL3o1K4ioPa0oaQTZRQBgvdr7PtEp
bbGVyf4eiWNWLiWpXfTS3IgJXD5CpO9lqcAcd8Lcu54xJsXcG4q8oCJRbcg2qWJA
zHlb2QhPXdk9hwtUUe1gloHTVS2Sv+u/zCjhXi4t8pUjVuruQnWTg8tmGGsXENLp
sHxN8u6Vuxqw4LhxYoQozk6HD9SO56LRSxvZ5Nl0qA8+Q1DMUAw9LmpAvWQaJ4x0
ZyGn7aiqLENeh+Ja/CLC75tkPI8Knf/3JsbyYssn8HnoUhGh4kKazve0kU9Z+jwZ
4h7luW+LmC4X1t1PoTh/QXCOsRVIBX0/qw6ibCqHwEqwBWuQUZdLYHE6FBSmUq/8
qzmk5FbD9nd3bbZJwIs8LXdITPjZTi+wq33Sia+IE9Zcn7V+hnkuYBWzvpeRKiPA
jW66HHAs/r2peMKlGaZgy1KYrxGoSuEtgErrkKm4ATwSwpbjgW4YT3VcKznH6nuJ
2C5lGK6Nfk/N3gqE3JZ5znq6ENZb7TSJYlQNAcTfZaQ1uXNl970CI3AWPQgAlVZ5
W0fghz49kfODP1nUKQMpabPOzkXSqLJpgoo6ueI303ddsRdki5hWcIi9/Q2ec/Jv
T4PbCRiIKYPrsha5+UhKuLK/+/l89g11n+/WT72x3OXSoiWH6g1Ui4g/1mPPyCmz
8MLOK45hfHPUC/jBEbfmdkpoBjdL0S94JSD9c7J72fQKlpTKKKPoGNgkxKWywOtD
WhKspkh+nQrWdfhcVAOxM199EUZoplGWzwTeuWEC0eTR9NN3WuudoOxFpj+f7Amx
+H/vnLBoDUez2YjB4XH3zK64IfCArg+7SNsnzs5hGpVx8lyBPC4weQcdNrjpIbVw
X9qViKd9OXPv5wkIWmWXxhivu+S8uO2QtEK0yIdy/ZsknFgxh+NZxdGtxb4kPQp7
vGj1BdZH2qsNpoGZlnBI4DXQ1klLX9JZvHSIc9EJFpNaW7e77eQkDjYNx581e0O6
8HbzkIf/qJFvorBL44icNrwwXN9oFFVGmn1xyT/g4Exlnir36DwM2PjPkvoEosJD
whEeQtLAzZAUebBCcReNuTRMtLrTpGfwJ6jnY3For4TzZVLsNzqP1yY0c45C+bDH
mlXrLebcoQAD/yAD4Ynq4X96VUX2Xl0ja1nSrgGt7sYQ5abTO/q30tyCepE0h+5V
xDYyGDIja1pwitAvRkYejiQYqEixi0eNvM/9uDSHwCu8c/8SSK4PwBtEY0P1wPWZ
6foC0LssaNLPzCsc8BfE8qZbVxVlqV7bpxjyvYCRuTu4ha+de4/f03DIL6ry5wti
VuLp8MuOB4NYvYIuWvmM0xPxqVTJ0PyTFUdtDeCCPFd2b9IMGqlDNxf05TFtzstK
aGCGAN9dNYKVbHVkpTrBQrq3ne6RLI7Dn77otQOD0Oa4QeY+Pnciqg2d3UE1j7d3
skV530GrjGuhp0xa3HGf14EM3cO3SCBE3KJzo93Q4bjVrIIv43zRoZpAD4+Weq+h
LUmeKOpJnNTkcC6YKkA335spZ9fbQLwD+a3eB5TI+LD+YoB0VhgCYQ+WPtyOur9K
43qUGydCiPcVAcyyqofgxw62AVRZFO4X0/8uMNQT3MTA7Yqy9anFa7VFyJKNXKDp
OO8uv8FvKntKOZxIruU0JRsUunHIHMe4uCqIWnSql4nIdiXyJeRqSuxlcjedktbu
CqmSjmzmz5BTwMgKR8WWXyzNs1iTN/8xckyfl/1FxGVw9whPHYUzNAW0+qhEaiNi
dvh576My7/WH7kE2tWsig8ZcqlMq5ga4zX5BN8/Q+wjJLrfAOyhGPfbUXZa28JHQ
ePnlwmk8bwAmPjONZIZLmNlwmggOiK2Bj1wtUW1c70EiO++h/xio6VpsmUSIPo1F
anU//iyGwL6GQndoCibjTPp2Po5SbcyOCQ3FzQENTY4eK1PgWGNn9i0f56V1psWh
tfPPehDD94GbE8VkUOr2G61rqvG3trNTfzO825L7W6P+rqMECdpW8RzZC0PIAwy8
RH4iHI+qShXfM7CtG7YcWL3aN5iIBa9qcIg0YQd2n87eLceSV6C1OO55OoOFGSVv
Q57pQJLClAIiiRJTv3byZTDDSy3khNUIMXYHNcSber+P4hNY1TAK+k03/LT7JxqZ
d9c2FxGkoMe6QGICAGOXCn10AT/G3UttQMXEqSGe+ICm7po4HeB2v6wDhQqUuduP
u9XWKqvn3cfo77XDZekYnipT7cZkgJBTe5rod4yNneTNaSOKe6K5LdZYKlQmY+7w
XHYUgP9n+fAmDMTu2zXMFRCxUGD/SLpuJzYIxTUziBcTYSXyGPvFkjAKfX7XIx57
KZY7JhWshpX+kzvXN/LABMbfWSjfgqGSHn8rMWTI3822fJeUUuMB9KBiOnsFpzx1
Z3IbrN+6pD7LjAWLaXZE9xnHAtZ52iJgVwZCmc+lF/2UTBvYr+DneVhIB1EeC40l
YCx9yNqQupeCgV73S60E9ahVjXCiN35XET/IYSAY+TUec1XVSRa3e1gwV0F6S1pt
4QeSVrxIJp+lye+1Rr5kqvUKU9blc5Qd7FlP7yA11KLtw9s7dWP/p273aveLoC9m
ZJLBXQ4GM7D9x5Y5szLgUD703ZxtVsSIOjmxURRB7kTa8BSzfg8xtYrLq7k66Y4q
99aOvry89W9+1Jm8fNTkJCwmpiniZEbqOHLxUYwXLVT/caZNReS3Z+Uk87Cvcw+K
bGjo9Csy/5xaKw94smHT8OnPtsYeZ443eQj5VQejtzulpciaZjZYu6IpcTfIeuRY
idHIHxJ5BePSgQ+DPAAjOUnf7sTdmVSju2LVL8UVXHYISyKaOJKbEK7zNDxf+tL9
JCQ1BVlAH2vIhczGsiONnCnh8He4f+TZ4zoOE8QhjHR709Lphj4rH0KqbRneH+Mp
5GWXOWocG9OifPrvmnSa1Gjlw6Ggk78pvx199qATIrgqCQ72EsmPfvPHHPKrIt3E
e2YCL2V9K3Bi8Bqq22xVFjM58dBxOn2FbI2olNMzkIL1coYA9+/nQn/JsM8eOcOb
fJ9N7cpAvS4IQDkBg1mwjBNukWhebl+nw9ROBb6RELw6hxmrxsN+zRgJxc3dXXXH
BcZxIvToqMwIPeQ6Yqgmgsc5ps//e03AufMm+t7KC64I1yMNX6pxweXh5WeTQEW9
PHQtam0HK2ovoVlBlpY3KS3vSiHmvSsgI51np0M1RiRzcylTBCLK+5MOqsAPqTS9
qXUWvMJoACvTZqn779rbb3xBV+jxW0WySvfz0dV8DOHpJxqhPynKlaRjWfeUkIZX
RpK8qjHNiFim8D65WyUIP8epzp1gBcChJjSVk5RMdiNlILpTj7QGCjopwYq07msz
v/beP1bvrZCPDyTuevDx+sotsGoP5is5wv8gXOm5ebdf8r1/m/BpjPH1KU1X4UKB
3mX+dETPzV2WI7NsJ0QOxcW3s9aaGLsvlIL/BCtr9tFhSXz/2u+6bQGD24H3ENyF
/GlCY6V1bVal2gj+3gfCcV3cG6JgenjgMf5qBFlSbGa7qUt9hITaijXnAWcUCWyZ
Qo4+Ej5FSngHRaPsJahbfL804UJSnwi916L6/Q14sXaAaJGc6mq5iQq74axHGMYj
mZNNUe6leXuTFbiNHVIirnGkAik9DfEcyJTAOAbTecKQ1uIinJlk7e199bMUMPOO
u0XLQG13lLVhtCGPvGuR1PC7I7dM7WCpwSJHhq2yfFgNdagNq6ODbHK/vq+9yPgM
20Rt1KWWKuAc3Bmmdvjz4agnd1zjangV/uyg0vlSsU3ghpjCDLSnDJGsd71gr1Jj
9sAxsuzI9jx711EDuAnc+hYLSTbwPHrIRuiuU/AvRKbnpYJVTSUOgExrzbmyeiEW
x7R0OUq913PWkuxAc/eYJV2V48tjsOF1UkO7vLX1Knw6hIjb0a9WWltLTWoeYuqK
UFEfDzuQIL7jCYINgeMAPEYs6d/2eD1fnV2oP87DmJTWpkBEtE9QYZbfrhHr3xE0
yVcZmHGtaje5h9pNplDtmbQWxbB3VlhSeYJ1n9gYgotktS42R4Wow3cdIk0Dwe6y
s1L46/GQmG1/8hrr50tYGLS1Wp198bv3NwWY9uyX0xTTXGehkdWC5H/vs9NwhSvZ
PyOQpy7HgqVIt9kMtSNvX87NifUi4VnLZ6e/GNVoUeWWMvSwRIOWwAsP3Vs3bSN6
CQOrsxDdW8m1v5jNUJZrkyfrC0bzdkmx+VHgWtxsHNl1BpggDVhxDtDeRNkD1d9M
6OZBsK2fJadF0TkAcR7NbfuFz/B0vucT7G7dIoUPhU7wikZF/1Iyjk07d5bZqMgR
lQbdHYLNRyEZRpnMCkTUg6gbKfcCTrPDzPf7gUXGcpRBIqukavdeFDpXM6nRJdiK
K5A5mt+zJtsCHUj57poB1HsbLuGkcPcBVBAjml7brVCtv/Pj4vv79CL3V2+Hs89E
ae9kdChOgwiVJm2NGu7abDD00pES0HWyOeqyLq2LZ4hOPf3XJ5kF8Ooe11ndKTLq
0eo7JOR+zMhxtJDBZ2dvOG/mRSR50YKHDSmiVgBiZU6x670rnuxGyBC7+eXK4Vrt
oJ3gotRQMoT2UsrYcnHzdm0h47m6a0+j3keuT7wB4SI=
`pragma protect end_protected
