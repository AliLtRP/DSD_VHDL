// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:38:23 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JF92HZ6G4F+xj9Br2j+sGbMeYoSX5jVTQZBdW4H4xLwfmQwhLBLZ01rMcuj5vdOd
YPKJSvR5gcekvehcgGyiP7pvPzhv3ETAZ20tQFsE3tuMcS06WnU2JGDetT0uGm9z
xFgQIY+miO04QBrfn8A5ORv5uy37IUWbNlPcHsKemS0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5728)
ZykE/pTIzdKRAW4SCUkiCFtwWWYdJW3ovxwS/e33w5tlpr9V7Ii1unuhwSprPH6b
C2+gaq7j3+HvraISjtI/fDuluQPr8zeJfpmxmUF7fqQhHYtAdRikn1mlvaihNt8o
E0/+VUC6gDKRsNomU5+NxUuADMOzLAHiRMvvL1/AawIuI+kgL+AN2ASJ3kh0ospg
sF/b3ylKG+/a2/Ag2Qy+73XYK1bfnDk8aZPwuEAmhqCuDQLqSaQopyscwBs1tUF3
UNV2+NJADau5jZXZmJBFG8lprN9oQRSyYN/Ftk5Wr9f8izRNt2OJby3mhCHpwAh8
mZHatHWXPmE1UlaGyTMv1RXv9TZLwnHf4Bj91PDzSIQey9/lG7Dug6qdFMK82lNL
vPvymUL+mOsKpsjvLl1i11hv9OcfW38BdFBWn8UIL0JS21T9QhOE/+TgFd70BLnN
8edHBgs2CF1tzWDT0p45Yj1gjLdE6OXDEzJrkMT7OBMC4u4vOBRkZ6ilS+VzzCBF
fPlbof1M8EgAQLE8XTnNL/ma1VdzKOZqwfDSi6n+bOg00rcm91NuoX/Eo7iuzEkq
veDQR1I35S7QVjhf3ETPy0jKopb+s/NdthxuOo7n46tsVBhz1mq/n75hM/Ihga3F
EjnuWl1k2na4tJe1SS0MPc/XCffWU5aLG6IfV+rowrrxc4nXtvUAkf7uuQb2lxbc
aPYjnF5d5JtOusXr+QE7e/MdxDy8p/PwKwALswdBg8AKiqSW/aUPAXM6GziD9ZLg
D9HKYZmm8ADPQDpSXgo3ZVmLJ6W1bVc4kGO5NXrg+fk/ps5gBwoWCYbKOAH05vP1
datFUQ8vDMUWSlNzbEQtkDZFN1ELsFmcxw3g0mzNRWpxbA9eUl91O9oPzfZavs7I
73ZmjFIZ+u6VTvTT+bW969+XqaVXId1Q/q+vdGBiMAzdrYqoKivJ56NxCMvpZkxJ
65cjqCXHyVmxFv3DuRneT7B1LxTo5bWXRMwIlAv9FO0xlGBostEXWQxdqfPEFeLd
7965KhgQ+zFQEYoB83z8wa28q4HwlBwyzUSuNrI0SrXablP2O4ER2eemtwkEe2Np
OiRFRDNmgO+GJomh0juIyaKOyqRuu1Xf5x/N4dcaNOr2jPgsvsyXGCVY31Bh7ObV
pBr/SjfQmYsv0YwJaGRh0Nr0kzqZYBbFQS9S+n2UYsxd2jP318lZPhPEt5EcgloG
gezkH1kbCntdWKSxlr+O2rfYbLiJTxcReFBM320QCKKC6LaS/SAMMlo4Ei+8Zgy1
iMVsHPgUxSMQoIg9RRW3nJIGjoGeLRsDoBXVsqlwCxkGzHr2CTDsz0W22if/PG4a
+mTkn0354JYGvcDnZ7A3ArttDvXiK3GOrg4q0jJlR77l01anS+r4mrJDEoRlAYMu
YA3t/cdWkRhefQrR5c2Jhk8pzNGGeYDO/8cDVahDkingWYTewXyz2TqSYKh09PTQ
odv+4rRO+2dkbBjH2PBeHjtWEx4eJw+Y9uQp7KXv+U5/E/Bt08ZFvqW1WqUcJyxI
A+cXfWuWyOoFIjGTYbdC7mBfuEVd86nkQpvPY1/pXKrOaEn7BHlxJsX45wv0FSdq
r3DNTpEXP90H8//Uhv59pZvRWdq36uOwl8MkJtFulR5z8zcdrEe3QIjQQ5SLSeqB
v+zMQiV87l+THYbP931/RSEm1uNAIpFw9JwmR11iHEL0en/fN0vVBYblG1mFaYQs
cLU6v4TJZQ1BVCRLUTCxkkq3LhqkkfwCcnT20ob1R9IpMRxFoBBJJgPSg9uCEzR7
AeSM92EiKxryn+9UtJEh8k2n2tgylGGBDgRFYiujrr+Y9l9D18g8m76OKJLgpIAE
lvdK7PsKrYMunwWFlO5cK6ks/G/MHMC68Dzk92hv+5CVjWXBDhj+xaVXRbdhV87I
7HZL4EHHuxRIhhVxanTb7qe/hKViU1/02QQTHnazRDfVjevra48Yp6pKryMf1JgS
TrP70WECtG7fEoc2TEcISUb4Mn73Zjwv3DceQOEJIhZ7EysinUIg/VGetWnktXkp
MLCoXZp08CMbXAkp018nVMvADgu3qFXokpMthndsAeMEefn1D3WHAn/yqSdPU70T
aCu1emMyLEMo24sxMkjoxfDjDQR5y8Lym4f9i2CwTycKDSm7P9KJDx+/9AsJ6hPz
LrarXeVZL7v/qOsBk5LWjBTQvDuNrDn87knXErAmv3gGY7sgWfOd+2Pdw5/UUQRx
g+3mT+Z+NI+sT9+Mb/iGe7FMGscVmZIPSZw4wzqCUAcFZEsa4QWspKCB8pfIhrYj
qNRSbazW0d/6/Os3JyteVO+90iOELvi6XOXBQfDl9D8DiENssdOa0pGqL53SfYnv
ICPC7YYy2fsRcfxyNfEyPWYq+JQ3CK+FayT47z4ou6wmOKZ5FDSaauTwre/Ac9VP
FqDNxSrhLN+3IEO+DNzuKzafbfO1gG9FXs0A38zRsBSLeNkG8Bsw9Bk3CR6kSj8T
1OqtwYiBum+YZEE8D8Xut9fHybkormCy9vpFxh9tSTWcqsbp3zN0q3NemsmTMOdx
PbdirTD80CUER9niDtuxdUeMj+enCrAGtkQELGSP2yrTa/UM6wRbZqFxfQmDvEAa
ndlRgB26j1217hx6zDMBvg/YTOr3IvbSTARFDzn5Qo3J1U4F0mWdpbKC/lfnlXF4
0cSDA6pLwyXH72ukgNIGO6iPwWjWlVMOATO0hFd3daLZqzUmeWLwmg3xGoI2N8P2
XmQqgXQv7CFc6ck5hSOLP5ki1U3/eL5QkqqOYvBq8Jxi8hPYwMk/iG+l1XKMjDhN
YdOlbtnXAqU0hQ3u44ct9Hus2i5qGBrXFubtR7FWTQL/eLS+nCVjX/r9fb8+Hti6
50VazHib7tPN95t/yYUXFsLg40RnbxPYUIVsFQimFKDbxP38ezjGmMdro00NxjPb
wphSawiFafk3P40o2RyI4siVkBinRwPbnvAZZH4rPY588aZ5cKTI1V/LdAUnLj2Q
DF0murBF67HsrpdPTlJTGD1kzojy1+leVvyMWVSubWuHN58eRy+npDytuAYOn7Ud
66WojLD5ZPKGYcZw44z+pl7xNMm2oEi0ebkc1zssi4U+oUcwi3W1N8SEwHhatRxe
6LwxQCjoLdc7CPXGiCtznDvy5cZfswI9RGWp9A3ER+T7gZhEyaCWj1BPq1Ydq1wi
8qZXld3+/2YnESTU5uMoEBt6MNHl4JRR98s85K/rxo8p3Z31Oh6nYT1lcF6Dy9WL
xRM38QXEokiow6ttOZXKYSrW/xARJPohx5QUonDshPyvcfMZ2cwTz/wTFAma8FYp
LFH8ChcSLPy+jcT/xdPD8Q8e+wu56YtY6b8IGk1F3ax+vwbDJOBh2JPgN04YU9wG
CQI2cmo2HnS3QunCQgvFUFZB3ZTZJDq1HDFcKPm2sZKm7GwtMpiXeWaFDtpE9iNn
zoN+BRRAS6eg/X7EvmqqIETIFn79Ui94VfN2cRuM4ATdzcRcxTXpFaLecw/NztyT
b3fp1MRN8k7x08boxAVV3rvfDzZpEx/dDO0PBIZDBflAYZhIXDlXwlzzcJUrX2mm
tNRNdJdqHhu9vS8puImgnAMTyZcYY/Ldg1SYi6nYIgfXBp+CP/t9HQJrzIRf9co5
6Xah9Z7GN2wCM+8BfCsYGTT1nlGMDzYUXylt4M372Et4I7eVlbnQZTvUe4g9pKh3
MWRoTw47hd6e1B2QZ8LCKxNHRmyjMBu/qCSHGqbA6E6KeQOm7VbhgJHhCdKLHDoR
6zRzkrh7Gdyjg7g7zoemhD01ot1ypCP3KzLB5i3fGN4nG7Grp7fYtnthuZqoejfD
Lq4Hp9cPfcynY/c0/0IFkeuEO5QAQIc+S5/JLqL10WZJsucP7N6Jl3rFaJGPw/V/
/X+2STgtQRdZiJiGgEMxpzen9BWr5//wD6MEf4ZO70TCiQl0AWSMtK7H8uQlTU7N
kbSH4+IZeiUv9pMsjxNNJ9c++3lW1dPpiLir97YFxgtiZ3GEL2vhoiVI5QMKC3lx
bsrvKA33EGaYo04FslDqg06+kUXLV2EgnOlNEBENV8GmLNOaPGDknVSdvRK6Uo0D
iUWe5m2Zl38KwZIs16uOAORvhElWV/KYLXZS/RH0JqDV4RbHAwBCTj7WgIy4WxIS
w/zWyCOjpFYcCImpe60arIeqpmBjr/0uJWaqNsHrRmmXbdskEn7IRAzW1VBgv9Ys
61TPwmUeo/plE6sRGb17/u4o9fTa6gQRbZxgCByNaurw1a5A06rgmnEcBGYMpUve
zOfLzn47on6kWUdV0y5dTV0EGipFMh2bZpUUtQ/2gfaTaUcOZc5tegf89Gtpo003
Tu3bxo9miO40C5sH4gCATSHGM9HsjQlo47EbVQiun4XNH0eJbAW3lqd5fzObAPSp
VqBYaY5hD71mGetexkYS+V4aukPjjuIPTT6BqMDokrlX+0Q82R76J1ArDhtzQswc
dV2htIlTPc7nrFMBVhaF/HZYdYktmBvoBNQfBYRgp8ldHC4gPSemslBiBa73cB/k
dqEJ9F85p47DodGpDphRJQBVb/r78RqHRuS6TD+mDfs6yja0Bb3Nt5WrOfjzX820
c3GbyJ9fz4A8INpoVs/n6cdO2OiMQzwRKuCXXQy/Eo3Ksv5tOPHF0bzzZcX/gFc0
0WJTMHPXI9TTeJxDEp9iGg9wfgyYI4HiVyMIdvvIY4oHmem6Nyt8WBg8ieQkm+wm
XKOX/fCBiZnPKON2UWXYxSvFplIYL+Y2Czcpur/Q+oD8yqHVZ0GWN7Bp71smlItx
1OLxrVDjZOAhsqya4xxB4lWFJVCDCrRmgcQA99vQmoU9caowlSa0tjIL9aRpJgAW
jKF/CtGWUtsh+B2g13K1A6vPaNuwZ5QVzB1bdSWyqExwBR/t/dQmXqriutYV58Fe
L9rTDW1iWUdF9UYeyIbSqvzxGa1skDmjPm0ZoSYajftibAnRsbqwjitNO8rgJIVJ
p/OJpzA891ueCuSe/EeDbGD8ZUokWegjxg3rikTfW9LiEtjjAGtDC/XfqC8RpcI/
6cdFlEB7ZDE+E1FDIwGFtTwIaKsDsqHfZgrimQXBXgxn/GYnMY0SEPSuzbRcns0g
TBZkfjxfdACntE5cSECFMavUDA7T+5vj/zG05Zixl/cCik0MGBHEVkDC/XYTGBw1
ubMx1/9uVSx6PQmlgwn1Ka7wSbFRcnf/+RELgu9845H8T3dZZq1tC7usX6mffKm4
u5DB18CinBxgKI0iehqJhXY8ydLyDQ+EnerXArK2IZtmFfYSIQCcKH1ntHZD6Yg/
dwZbvmsZqEAughNgaK/OBMdb0hSam/ixFr62OXLYXBzUNRcUqWojmCSI/7KG1SkT
QYTBRLGt6CscFubgbA7hbdDA0UTy+p27942EPPXCI6qgR8c0KUdCl6eyFg0Wv3X0
ZKz4GTJrC3f00gmRMRKAze4fBE7fZRx+SHLyXAejXzwYWG2POOHavkG6Xf9pUf7K
LunPw6WGub9+EL5SY3SjpADmUIjhwn34cABMC5uaOIyzDlto83K8s8KLWOcTP3Wo
ykuB9eVPKDkKStdyIkrJlvPWAwMgItD0tebHaiuqNs/aqiBbc6R3uNXgI4g3UEFR
Us4dfqYys8EIBLDBVfhwdpeXdUMIPBaHd1nQOsByfBpUQeFwM34mCp+wQPdSHKfp
vI6v3wR/JYDkyCkAvqQKYUsycfYp4kA+QbxQ4rM4U4S8VnZjqVx7Fn/nIUz+CsqH
uZVRrPEl6szRqywl6iioad2brYXx3e6rNs5uDbKq7Z5cj7/m0UtWA6Frvo3rEGGI
ApB9CkwjZxQU1p3MYWI8czrpm3zmuaxuu8KQGyPGBFBo594BaT6Lcf9CfyZ93pG/
RJmNAOvJXw3FZNf/+qZlhx9UxLUrmNm/1pVj/sIchvrae8CS31aI2OpaBMmJLou3
1D2xjXnOBZOPyaPnpoiT0dfDqd1FHRn/V01H5OC0iYAejwg8pPxsVkS5CkjN+Urn
H40Re+C42OjqW/QyM+lBQoDxxgIk8zz+OEtVE6gSP69Xfh+iUR9OBHfBZ7fxeGhp
GmaG6LZ3bc8l+oM+ouWdczOfVNeAn8O+bWO/f5PYJLERc7b7EdETTDIrzlg7RAo4
+wk4FRlLQvglsSOL+HpQWgP1x4W/ISGKZt3FCDTjckbKagVkmRe1fU1rdN2NGCR9
LSFOyYBAwdagQ5gfKtBaH2xvG3IFTWDjCnDswix9RZseSyGyqEXdoS4VY5cuhvqV
lzbAQ0d6ElLlPb9LUH2mPUdA708u12jxfJo8GCL8oQHNwC/za4ph6PCj1/y/I3hC
6UBTH7yhshW2YYwqCZXiEQBtK8W+fW0pydsM8/BCMuqPOvh65VQzu8qSabGrAU1C
vyielS1oOGnuHTze+ocVNOKBOgC4nUn8RKKKLurT+P2jmz8TeHQHo43tJ02R0Ip0
YKGlN0I03nllxVZoQer0hOPxKHmbypyIK0GKhS0vuElORkgtckfqRjvgn4RL0A2K
VWTeBhHbPEAmejmihiBPd0sPMk5PmrxXnXu5tjjlC0Y8EcuS3ctLVEBpoIEnIe44
yD7jd3NRggZmvQoZFJ4Wbbh+eJA00zgStcldDiE6QBrNknq4QO37E8UQmNwjqtlw
sKkuBCzab17YlGQm+o39E/UdcBxs9ARWs7YByVb8Wl73wS7Y5hBXwo1V7h2R4eBX
0u3BwdkkNFJD/3Vi733tJDjyGTHTM/xuFlDDRGEftktZZTgapI/CY+nvdjv1npV3
e5wOEwbw0+8HUrCSDNM+pAr6TwHIfig40VEIQuc/4b9G3Hb9J6gbrF+dbXzsYKTN
/xUw1CYS/Nyep1p5NzC8OZEdOwFZco9ZCyZOj3lUYGtkXfHPmGaU+CiDSaeXbI5x
RGdxMi/oUgFc0GDUppJbK6G+CopbpY3tvLOS5/cJDrMFBha6SYqBjo1d5bqQdYdL
twPSsdXdzHeWgurI6WkqUfCyIlAgiobKSRJ245EtjtlTbxX8dbI4X+7UKpzclkR2
60IaAdhyHBF/AWINIfSOGKqehIwYlfpHfQlpI7DCNwLRYA3sHmeqYoo6p42G0YEi
YhJBZA1nL4Z0utHaUjkJbkctz0+qTeZDrn43TGeIn+4xmilXxJjslY1X8veALn5q
xpXiHmW2W6YFTlsTYsaSgCsqE9vX1Eu5QtqKjmu44p6A15iNHl8hWfR4Ad+61G5V
3SpMBbplSUAZU18UhG0OaEG4Oncn2NxTuWBfIAYeN74kM0fDchAjdUaNJtJL0o+L
t1VvCfMSuPHS98ykR5YGF+1tIbnGZC9f5TPF1jtpT82z1WdYTWnDIan8CU6oQsyD
XNJt/5XKb1zYNN5QtmQmzOQsR5RpAPjVD2NCTU3pJYi1D+upl/RHxl7iSnzcbYp9
sVSGAfYbZheY08xKjxTs55ziQlA03OmgNkqWL21UD4QDik2s4jFJpwR+4Rc3LThb
sgXlHxYUZx7XisY2lh+3inEUMxRLer6rHcNN6QKKsGMFm0NJtBrxj0UgNqz5oz2o
V13pFfnnyC19dDNQ/oc+DShsHhrcZseb8bFn2YF84NE2+H1oYtgJcs3RXblJtYlR
3mD9A9UsWGC8VX2UBZ5BTA==
`pragma protect end_protected
