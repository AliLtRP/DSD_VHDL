// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:36 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kwpUQlYMsUc1QoQh89JMv7TW2ptNQJ5CcfBfHiiLvZm0H/kh2j3EiN2RdOOgVah0
MEcv1Dcg3iD7gPOnmQ5zQ0C1xb1/TJlOTz/xySjJzQz0gxFH+wssP59jveiX/EHd
z05wMi4gcbRDpVf/Vm8GhTr2A398WRAfj7YMBK9RP0k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6096)
5WIpLUwGdcrBaR8HKN8sz3EGGeAX8N4GWvuX1IXwG2f01mBD3PQkTspBBnd+e+Vp
dyaQFOXYQQyY+IdiTpy3uEmSKyghIKRG9bxZpRSvAzUMWXAtoBOERce+PpyHLR2O
rHsxGR8Y2uxb5O+OuiChdaixR9mq7yczfQVC+iVbQj8tQ9iuCcKxgYe/4Lf3EGc3
2OGSN4QwkImMfzwELLpifymFTaWvX6YDBDCWmtBaBIT8XG5x77G5/tqLhiaqQ67b
pFBgp++CdnOHrgs7CD1Ap0Og8OK/a5Fw2BMv9PFWx42apNWiApdW6R4jS5EVR2aw
Xj1/X1vlwovXb9TnPSoWRn7ypAhtAMNuQ5fR0OvuzpuZYjTO/aQ5DKDdzj0m77Xb
bo8R74KmQEDSYyXUpg/8An1ZnxYX/Phy8Tl7FOvNinR66mHqIY/DFbltYXwXQvoW
qJoUb3QeT89MWMQU6LbBnxOxdVIP4ePlKN1y85QFNuiO4HgbQhOqhdqkG/eAKdxR
87GF57kLoq5ST8XUDLla5n11G1RQ0kcaHfSVzIB83GrkKwtpIDdxLmnoZjWoDKUA
zI8qQMzwkQaaMiGKcpm89CC/leEjAR90AB6V7jY7tlC7kTS/VP8ZeSDzbrskmhks
xXcuezi+XHwlRRHkmi19o23OV9+ONfInBfEWORAIbnsiFdXeLSyKPtP/30nDq5Pd
tOuZecqY8SlpZrAQn0NS42KU6ntHFiKyv7h/0HP4frtS464EzvCfyElzHqa68WnU
bDyiKN/mtTpYJA5xCFjaY50+xi4k2tQ+ZeLjXnUQchpW0XIN4ehf0qxKYuUWCAq8
x+xaNK7XYLnu0jOtL9rOMwI1y1ZHE+WbPNfonIe1jSrTSQZT43jc2GwFn7boc9zR
n5qqUgycwC2Nz2y38kOLZDkW6k5DC2cpm0RllvgEheFypohuR8DgsFoPiazKes81
kpDJWDPwsZnypDlG0GCTxVZbA+bzglk9f+P13Lz7FEuSMm7BZVV7sfY+mKsAj8wN
ovUS+j0DzHO+Wf790MuT2o30s5SfqiyAKvCbDEGiwbhAN9DMMgS44sdJdatrfPWD
D8v+x63UHYRX8ra2IiHWBReg8tOMjgkFGoQdAX9WUVHHdb4TS3ne/kPhCZNuSVVG
3iReLlJjS6vCKYWBFJ0n7h+u8zqNz4e3hcREArMIx7ev5/+sZzb3WiygHPpp22c4
TCJlIz0BfWs+x4aFLQxMAzK680AwcPflDsjZfzV4O7Ky8zP1nX9ovvSriTwA29MM
u/87fPxEVZiCHhn/I0RQl0WnsZ1qpkOJZiXOdYXNE5vOK/Ttca1MDUXtjbP8ikoi
+mVRTElbuXCxcA1l5Q4OGBuL+qUOI3Vf3WlWcSrplz/jtvNANI/S2Lcr7BLI1Yvh
y3JNIr0PP8JluCDl/9U2EwDljeTC8USaga7uS2MmzDMQOUnBjSrPxt/PBXiLFwBc
6j2sO5frfvC60FZUtTW5BaHkw7QRMfjltJB2nWnNvhrB8RBqygZp7KZzWEFWuDbA
FAukK0vbDr9ccPsfWN4iB4cKnj2iduVeVOEwmHVfB1ySxQ3cR1Iquk/PJ737DqVI
gFCneF8ozKr2R8+kl42tvXQ4n+yOygqP5nMaX6Fc7G16U7NLz2+DOQmynMlSzKpM
rPGCJBQIo/DdjuUdKoJNjzqV4IFd/sxJ5hrEH37J+TDLEdfZUWbK9aFanyscwd84
OAWYL6JNhoQ6zLNy2c81EJgbc9CtBbHdMk+GEwH+10ThNL6b4JC5JAbIIINeWe/D
mXKUut4NYDEdCHPiIKaxC0u5pZG4WNWMYbg2vlRLo+p5/FqpB+a48sUJ74sTSab9
245RRtxlrvRgECFXe8eEV0EpSxSsWYFVMcHTEb6Vz++SPBL6SmqTYjONJ+XD+tCy
m886SRc13YCR83LzI9xrSpIQBi+WREBDk8aeYcpG618xuD54wintGX2yqxnw+RAL
xZ4qwbIrWe2w5keunoUteiTlcL6IHMkH4ixT65TDIPop6ahH5zgRp+kUohRR0e3U
WWeZH9xs8nDRxe8MrDY63ijISHhOX6P60G8Ajdw9BH92W9ax2iReRCnDa9WBQsJX
N7WhEWLtBGgVYPY8bFbAO2pqLHqbaC62xdWRThoXBOdyPSN73TfW8IY3VXuFZqOG
i2vuFTVILKuTyRoFgZyEXIe22mg8Rue9PR/oEiscsmRnaToHFJBIcUKtuivjaGvX
nh5fWCsgkuC7V/SRyw5eRixKrwh6hwSPkPfZQ6EZbjrjeGYK25o5bIsu2ORuYX64
yXu2KgP/QS6a1VMQj0XIjxWzIz9SEBkNyfv7NLTj7LkB6kN7jCckDaPM4bd/ouM+
NelYa3IOEYZm7zz36bUWzK7HvLuLlCDTmlu1T27cDFWK7izEUa6GXOLFPTGAf6M2
eM4WzW/5TrWKUpYatkNg4EuaxTVHDvKpd5Tyuq87hy3W+EwReUlS3bgZXWDq2Snn
WkTvOmX0cRHGj6X8KhZ2Ash+Q+70Hc2IIl4LtJUmq9OVZFNXwW+A3tZsehj6VATJ
yEf46HHJin29M+jBkSmP/PXtnO5zILlcddmufXtApC7QbR24cOfnovvQeyIOksNC
fJrC5r3lEhR494ekPjnY2GkTDDFfcxe0K8qy3blZHMqzXCPkaivifpFBb1IjtA8X
SwVrZN/jr7SaEs+705uRxIXSmzGb5SSltacbqBEARXLJQdWX+xW0HxyDe5la2Lhi
4kiaVjh6ooZjnkhSAF7ajqyxN2AQWXxmnm1Ll99IJvEpt4cDZMFi/1N0jl/t1VpK
/vcLPfVoh/0btGkQljeYTbQRcyEHcFczDQVB+4Z2maj++1lA6WBnk2Z3UZvMjmFh
i0Ya6NGIbQRSFXgtAgGQt4vcbwmZF3VYIcBKZP8js98gPEA8yhTugm9jysUkPpUt
MPvv8eOM3QhAGUHYpdji2wdx9f6ytZBn6RODifJsuA6gb/+Prh27IaYpImnvxxEs
7HNVkYEuZd3O8Fpyh0txLKVVK70uqfJT0MA9/7+TgPz+4YT1AWwCR1XoCRAWjsCC
tE2OWqutyZ10U/H5zFSS5xyoHHvFbWAz3wOvsQwR+Ox4TQga0kPLB2j/d0zlFwF3
AZ0asXKbD7ohHcV7OTcx/XPUxtGypAGdyc3kSjw6dr07rBA9ktyZoauhPl8KwK2F
5g/yG3EX3MeolvUqfb7dKkYN6lVqiWuaQ6DBECLgvhl+RCyC1LMTNoYMhhemg8RS
U5DpzEmz33ZDLoQdDUe3n4OhnJNruyK5OKppPtHn12AZFmYmUsNvY1X/gXn5R39x
29YUL4nouwf7YTuG9jzLCjoTAwe55HkPtd0RylJuh9jjzC6lMhD1oO4hSHrogVS5
Sc4tKGoTHXoSRukwcVR8tagn6N4cFZotRKYXMPS2SrdzAbcsuKmu/+I3NAoBhymq
ZkpVpydxSfLGhNHvRbWjB7T560glSXucDct8dTvlmvXOHdCLoauex8JFNAH0ZTF1
ME9XKZ4VWQR1HNmrLj4npydN4uYTXp7Z6IKctyRqZdMWkVd+JjodOPKf70FPW898
dNAcJ2SmReAu6xn2b8oAV3ygxGi2773kYu8HN+2XF6+HOfCDtgIx/iqRIHBgLIfn
8FoI6zue77NEQCHTSGsQAeW2lt9DM9eW+osuuCCdCi0/zpdfRURCTenaY8OXFbvu
uln+Bzp8+y0Byh4D/9WVqRspQneTco3c9h9F0q1NJODre0Jy4EpKKeoip9UrbJbT
wRykPe97AGGbzJXYgLxZXZtU+ZY+Vz0QIGVz+n/4evYArXR8wbyLdc2V4lDcHAIX
Nz8av3JO/FzAUN8Hoj5XXGAnLiVSZP6jkqMV9QZjugsDpqIUOTlvn8wKMnj+H/PD
9mQmkL3IiSgfWuTEWiU2EusCN7CzKLO4+FcXcR30YW4a2a2zyDvbuVsOntYQzpyf
wmJr+NSpISC7G6YalNozmqYLF/UpSeljQNUWqI/mctSEXvD7rayPey01ovFcUEJZ
y4gq5+bE4y8Aol1yGCNgD+1pUCFscue+PNgDNfWLpawQPwcQFtF79yH7xqSm6qnH
hg42bZd/nBGvKwP1myp0MTlseaEagZbpYMvdJ/fGzOXKe8O8pHrUl35rEs6g5rH0
ekcW83HkbXDPHRp0/CN5XPJeq6ZtiNuCRo7JHnKidl2b9KcOyJn20R78F3GPgHi1
0Z6bUaQ/CS6ihLv/4wJhtsEKd6oEXLKtWmG76aCSLcOk/bNSK2gY5eg86XO06Hrk
vd+Y6Gz76GW8HRO8jKaifSrz8Q3fXwIn2PqYciChqvX2ekWn5RcGSoQKAphoEkxQ
tcw+jGBnZpqVkHSH1loipYj3X1CL/bA8/p0AsfNR57dib6ClNBZrD9K40s6tRUbV
7dtNnuCmziuIfXnhIBtc9oLymGdGiZ+tduEIaEno9WyPG13f7tcyX9TISrVLItAr
eMq+60Oi97g0ROQhgRs6VyptsGwN3pimlyiqD1cH+lPz/riA5ixqlIvwZI8B9Mk5
AaL3oOa5FvVTJZQy9njIZ3pBw79HOA6c0IyqEAps1kaIodBal6QIxCDSIxlTxl4A
hLoT4OJc1fX4EDMUFgeyghURwkxgfCPfZzIkklRwWqlJ+uID205eSDQntZx0hYle
aMciyiByEHBl9FMH1Yl1zj0Lo0u0o04JUVwSrMkKdeZLEvzuLi5utw+iiION0eeg
BzBr8/PV0KXrhaqcbd28foXeGC7ENgw87wdIiGSmpl2ApOohPTq0QglTQgg4v2K4
AkTlX3veCuwqYJXqpIDkZDtN1Sbquxc4zWkiIHkd+yHYsPKK4XWqBVI4tp2f3+4w
AgYpokAJquIZzvsTh9s9Zz1B3L6LtRjpoGB/IR0X3qvJtkzuOE1mUbh75ZysroFS
4c6i5GKjlNWdvnx5PofVHXN/2fYzf4Ay5xJu910a1sO8ehM+kq5HNaVqN6ton7Fw
ogKIUdLNyv9DHLJck+YlPhRwVF5+DyAhLo/883JaPoZEh6Zx6qA/Fr6n11nxknZ8
40/NgE8/I8t5/hZNGDfYQXz5uSS6qiVAgEs/Kp7OonJN/+tk20N65SeaARwajPUR
qbNs4+pV0qkxRkTuMjmF504Lvelk7nSZmxA51AnfKqn817jh940vDpOnawgLbkoU
b+DJC0RKKIPi3kRCHSyyJB4n1e9NRiS2WrUXFD3Df9PMcMpqDoQB0M8u2EruhXC0
//i9Gpk+DBQIAlzxaSGr6D6gOur1vpAjsUU74ICFzaU2Ul/wnh4S2W40J6mrOY+F
gc7ygBxvblnqmISTlcr+3935shfQD1mKWx+tinpdczJIaVFgUd6HB7Ytqb0EA1wu
fXvU4uOOUFH/wIbXQlKYOi971sfUWCZtia3XYvqkZWpJu0jXSPXBCPJQalaY/Jjj
6woLBl26eguKnLR0ya0/kFW+bW1q63rxRhjcuZV2vpbHhN4Y+Zcznt/QCbllpUDL
ZYZPVWZmTYzMDNw9HQvo+Dx0nZTX7MfFhWeeUYZpvpxGc3KAdW/Q2ZO0/mCPqkzc
7W1+8gQ7QchpvNmsgJTYrrh7JWOQGo1WI4Qv+gamqffjvV49PAZiZEwmw9Id+Nbe
bbYdn8guupOdJkki7Gd5/jp9GSJE4066Xcc0u4uCUieeBZ+iinmLWgAs+jQgKSSC
UxsG8t/Qcyi2Nn5ZXc9/i+RP8wLnXUmBuNey26/4oeTgEXwaiI179Rgdy7+6Bu2g
PVu7NMUU1Y8Ej8Wbqi+sox4wkq5V1dyAf42P0OpywjKsnCca38OLkEUUmE8YtuO+
jFXDUmMlvbhO00loa5BvTkWArE1NE50/l2LVRJzgKZtU4BJcHRV62Ck12IyE28W+
v0uwS1MJo0X9U4rmnjiFTYgUA8GIMOxqjFvndsbl0GkF+KGJlEqAeOsaQm7THlaT
NWeYZRepTFoOevLVz5Q4AO1DAzL5U8tihrYeb7kJQnGvdCSdqBGUujGrHTWRbU/R
2k0ajSG3Y3BMmyV7GtpWAAbfIIlC/Uf+hx5WumiIq/yaVUs/ljIvSAiMbBPfLYMX
Xi6hY0A69UyucEJuzxcElfXsCYf5lSQlrxpXllKNpoj2Pbz3ni+JvOe26TjCumjb
45Kf824CT75qOiZAoWtsNqcshQ/c5RQrthQAD0CwjM87fAQxGzikIA6g6RDfHO0m
q3xI5+IEamdQ2+dy5dcM199o/iwaIE31Joy0qF+N53plOoqMq59J/wIIB2v+o5mX
iVg3oDGm1qr9g6/AyOZHiAwmQG1wj2G7wPlDmvX7csEkZJd96yiSzPVBKsMByLoO
aeiMGWA4DHFNbBtX8YsE8RwZZUDtSiW63r2s6Kq0vcIH2QcI9U0z5eiDF/aQs1kl
LZRz14CziRuU5ahI+XXZDL5NLAW+n87MhW+cpRsm0tb2RYJ+sMN5vGAuTOXBNEOJ
dq7zc99c3Y7Qcl8yv/Nb3cGc/wXlEHQCSPIkUH72fd1lKGU5D68F4YcSbrSOSwTM
lgxRT1rw3LNbZk4slMILA7D11HIhNlEU/QaDYQsGNqVksZQY7KM+M59eAl9Ww82g
09wzq7fmMT+m4y6N1zHVTUQ54PQFN9EZ8hC7pZx5liI2pkMkStKdSbyOPOAN3feP
dDXDPal+zNtwBbIy/QEGIJ5y8c9p92JrMsKqNf2dmm/NV6nUl1SJXr0TuTjo/Oks
WhUdyqtWazmHjtZlOcC1SqU3YhLP2rfxxEQEQK0NLW0yQ2LGlrhYo5uCKVBm3eHq
hFKEr3HBik4KuUYcnDaCJfgjFLweZmb0L2vufIGVtbgOU5n1Igbq4jDiwzoOti1/
fJfcumYdTA4bDshVUc8LHSW+MtVDxVO7lSo8NXWcoQ4cHnzPCP1Xewvm4XJ9aF6P
buDwOmiHbDezBu7sQfbZseHMTjpWUloGvMvjr8abcABOLvXCX6Y2AEj5gg8Cg6NR
22sab0mOWqPdPRHcvtxlswgVrapZBU6hkM7/Asd9iJK9H/oEicyk5/TLDz56vwS+
fwEwfHGZADrPpsfmp+lUFc+nAC425x71hhU7ps4QPbX2/zz/YkiJYFXGL6C7uy1C
mCridRF+LTAcSlFtjKhFu/UV/WYJAQixpKLpopSbB3IJM9XQV4lIWkg4UfwvQ95V
ECEA9+vW5iW8G0F0IxuwySOIuZrUEGrJi+d+wMAChJ1gokuS8IuuIrRZGvBzo7UV
yOBBL5qTpkx/stkRt34tzoiboTd1Tkm3Lv2AQit5XA3q7uTlyOK/xeDyB9RM8zeJ
2lDyqXtT8M9IOhNAFy0jXaa/M/QBEsOLHDgzUDeIYMaxHTUvet9e4Ge0SXJzcVCw
ju+f33yV6IAOXC+o69dzBKg0/NdPFT1dxBezTBjr7eD+b7+rpQyeuZrPpxgO/a18
rQ+REKxbTuV5oQ9Nxe4E7nUjD47GoeERBY5Ko/fDq+u4pdG59fKfh692lQZ85NtA
M86c1r8N0Fs93r/yojYYLPoWCYZmGEOMSdII+E8VMu7nqnXvmMkrRF/CaVU9wgl9
/7RM/sVPVc2ecNsX4mJ/eSDJp0UyGwPPhR0MJsm5YTInFh+nXDv8sbs0W3hgpfKz
/NY0KQi3esatl12lm4D75KR4rq1GNpw9zGlusiQwEWoiC3imVoVYYRpBAXEruHhS
H2f1k3KvEXQbFWSr/Q+mw0LjMUhkzKaYx3caHu7DQkWNUsRpC0D0DepgN7Co8bBH
YzsE/CHh9jiWywecbi0/bBeECYVr78UxNZSAa5ooQIUYVD+rKFf8eC0fEqXTvqj8
SL6CDxkI7Y6kGQWZ/ynQH57BRLxPRO2jg7yLzlf5Gi33ksmZQwJt+XY265LrIFb0
Bl9/LgojY0/ekg/l0HU9Ch1ANpERZqkP9NrG1KEW+FGnnjtXzWAZ4asjzuWaND+C
zP530o6YJHKg1KOm99SRTMpMPjsNv3oNpOFCt11PaYd58t6ZlgMJKkXOcWAoBQyM
Wv4GCHxFGWByh8UV4z478e8PZGPy9nKlR++n94pt4GHgxenT2ocsXguWXbjVtvnA
7u4fmdFigvzVXIywnnAVS2R6EEsp3u241VRk3R48d5AO0mbnGsPALhmuYLEbTAT9
`pragma protect end_protected
