// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
VUMTWF2TZ3KXVIvbWP1Aad5Dw6nvj0FkdApTuAKmIqBqiML0YqoMw/1yBfhtBmLsrulot0uEHYmP
afjc5ruJ69DvriOsshNhmDB2KiI7J7kGB9JAfx+giKYWjxPZOa2p8e8KX1VQC/qRPrKo3WPC2A8N
0iG3khgkVl7/wZBh4ed5Kuk7fIa7KtwzRppyq8YtXNGfsqVQFrZpet+kUOX57wR8T9k4VOVPl4Fp
zs8pVmMdFEg3dmkDww/i7O6y+bhCymyPL6ivLv+VB5Q7nwEoombnllnwdXmXcF0y7VVJkwA9IQFj
rI33WWxUong9fp5cJzdyAPkcZvjVqhZ5aHFusA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
ZBghhB1UuFvvwrBGH7/q/0LpIlC/v31qxVucQRorkuQjcg7nmoYuAcRDAVsIWP2ggE/pCH1dZioZ
CzKmyDHBfncK88BGC1KvCMvxk6OXrULUafxwu9xK3iHCbaYcbFD8upKSiK7JQMD4JQLAXYKiyVo0
Z8KSC7CiQy+O6kDfE/3bBaryrIEo0W58XnQrgtv5DoXfLy9muLKFc/AmrQ6tK7DhGPr/3h0hwqMI
q+YqgAQRtA6Qr/iXSHCdBTQqArKsMGHhSEd3cyyx2gqJ/XJsoACfcngLshUkIir4x+o2qt35Njhn
7jZA7CLC5UWaS0lyxD8RxPCbB8+TfSFBO6MjYV9qOYt5/LQqhDxJ2sH9TB/UexEEBPtPi0odwbBg
4sDaNPOUUixPKOm25ytvcd7q3juyNLCjHlWhW6BH/E6Abg/2hl2X92/KutQPJAuEb++V0BI+a97w
2hGSyTGIbh+fI20GGqE516lOl1GtanO6aaOshAJc0PEEmy8xm/ztTJR+bAEWQbwq4EVBwWuOHclR
d+9BB6SfNBokWYLfJPhacbzeYNoS7o9MYoB7GVh//bIKscUR81uEXZPRd2NrXbGY0fLNgpfuoSdV
2kDrXXTAfITx5kscqoQ+jS6PwvNFtT8KVC28Uhy2xKsToMVwUhg2izKsz9IMI6PWuIAGN893FTeJ
aueqnitMXY6LKtBebK+NwXZ7lC4YIfp9Fy5G7Thx7cGJbE1nXVK35j2d60VFIKryhuQJtIggj1Gm
KeKsQRpLkIMKGEQRthJ1a5/K7TAvn/3N+2ysl++hw3YwqgktonC6/qmFEfLm3F/mmSvktIqGLcgE
9Onbz2RJiD6utTe+j9z1gLnV7d8ohNB/wWhVSRg+iNwiUPXSmnLo7Oeb51x1lCDfx0Nt5GYS2ORk
hbdsyTI0dP1Z0QlmmOBeFCLMXpyOFfDqYXlJcQX7zlFALz55LMmEEIKu3zVTWtklkH+lihdff/+I
+qY41Ds+m/uvFcM9avmUhBqEsQ1qGPMrHzbodxi2SB9VQbjP2OZihaXrAzHJM8+MPSap7l9xeIJz
PmmokEvzx4jkvUNH+cSI59860dFOUVoxzS9Lfy2y+ebACS6rfu/76swfrlxYymj44nJ4OANxMOWm
BLX7YRpaeAU/xCEN61Den17EUMCyqM3wW7CR3D4gri7w9CK+C4QcvTgy0Pa59qz/vNbYYW3zvk64
iSiY0p1Et0dmmUSdjqNYL2GwDMRAm0OLRNzD96xFG75tZWFkWHIYo8jQRyGJsg5/2cnObhrxagld
MAzSeSjehkrWubWrt1cP3ipKb1Ty6J3uJnUpOIjvr8bKfVynrUG5Jio19ZRBg/xCYHNrcxv4ezQB
4BJKd9ESU2xVB7qjVNkvCx5WT84hvvOdFQqKrvddjGUgR++VxwhwxeuvPGbkDYKDEbjxPis4K6h/
dYhJR9tSr541mTfM6ALVZ9Gp9UP7O2uw/vrDa2lsqnkP225jB2wLlG/mp8EzeWuGHEYmCbwrq6po
14Je/Ujv48St2T34xTTawpZf/VbRSG5w8TtDnzgNqo5//ygw/RdNL+xt5/0/QGKK3Lv0aY7J4AGn
NjLQYpPDQzsK/lhA728AZoa8/HiZYFQfCeudsK4GEqy3M9KUCnNj2gvSqUUMMImko7ZUZkDlxWKx
CiDnoGhRdDDsKX5UFk45ldeuU0M8V1uNH5nO7GkFeKMqtLyss+8bIQRpXlau+9MjBnU5jm5167Uh
W5Cp8w1kGkFrwF4ONxzpqZQkqo7KsRISmLgEg+gdWg9ssuPpHioeJCZPvhhagRdfsdWsUZi8DIzy
tZ654Rnyx7fLXtHtSm7+Mu26cAh8CCgNSpJAhHWBRxUpOFMkFCYd4ZnC20AYOqao7PaulOjA3a7V
rDmfssth3mSVv8Zg7mNA+U36aAjgtQd01vl8rNhRBqfeXsA5YcQreE3fqfBBk3W2a2uWo7cWt+b9
6WPd4l4b3DP6jYaefnTlIRH+VQdSl3cGC7T3cMPaLZ5gaTqF0DWis/eIEPwBJgUdiKvF704jo9cB
H4xvwjya5O3M1Ma1qqNxYCi3laKLRTwr63AWbBWjUnaWC4UC5O548y/j9+OdeM5FUvzbZmc5dHZC
PbWiqQZ0mxGiDwsZTfSqzK8HXX727KrHsTMj0d0TCQ1ju5ZrOeZw10v6Ez8cqQwAKUv3YQsrKa3K
WlBtDMZ3SFbLvjMj/TDOTcyeaziy4jqCH1kfZKK7NVIPhsdUyN2+tLqiKF0N3U5YomrW+dR3U+Y+
AGt5ODIMqAJJKQVdnzRLTANfRIOFXPEmyZn8ixwVfmlpdpnznbMERgCHY3/H5pp7R1UvFx40Mytz
Jgsk8WdAU6w4pD9n9iM2VL9DLUgNpwIrMmkWlk7zS0vumIYm4NT9YwkpjFlbDptQ/BNnJjwjMC1Q
M+yf2yjzo4vzH5yISS6Dfjve95k9/REdOkHR23k7Ot6TNMYjzUIAn3q/DhcRw5wxuZn7iWXGIEA0
u06SULTo9RevtRJT7fa8duZEE75G6raZpRkE5VI7L+Nl0sKdrSI5bya+cjR65sJm7kg0AeZp2dNt
fUYmaSER0+wYwwovKZ4ftHwPpjAaHE9DVAcM1fq5Zh8VXADLwFriIdG3VHmSKKx033FQ6To6nQXe
aU4OBNQPSefNtZy2HoZiepy907oS7ZMhihzjm6mWyVWSQO2E+54oyWSJJ/XMQ8jAbCAStegTwe7n
Y/pinnlvi8On5CU3ET2Gp/Gxg0gFHoYs+YiwNZHnOJ5hkrdkVPThvXHuJKBkmmzb9+boEUr/X5Cu
7CxHbLbNlEDXbcUVKbQFGmBIpSJMHvgjmqlB/820gMEKqd5dk870QxS6M18icEm/ZBGwthGdAOhS
QQupgkPJKJA2DCqeyTKvn0VxVb+1tfuFe1M8vn2OSthMW3sggGQXoBINmoDVndHoSPeNPS9WEmPZ
rPSLw2qrhfQzFtq97uF9IID7UfpDngPnR8Rv/paL+yTJlQ6TPuoaW9nWeG/EOvK2h7lkg/RrWlhv
Udzd5DOvf3nBbgKadBFebylQLbpvTcjgRPXXwV/ip+Fs8Ysp19vIFjdObYbwIkgZXcRtU9FmsB/m
39WuDFZOH3NTLxXUwqRI3neW+FCPnwO7n6nf/KS6axCgzGCPVWlnCfT4O/A9wcA6xhZydLcca1Vc
kTbpEyRur1wDEb3vhslb/iRNNkFxqnki/poINAwY9/jxO18juARpZRNx2Lf01JmcNKAfVTysaC1n
EKfjP57khFK0osnT/aggfE8YUppeeLP3oOo6ErWvCBc/tMYAV2rc1SV97eKQHGdFPKrk4HkORrPf
V/OTOnhgyfKsMjUnH4N6xIfHGxOZyIib8TyShiVHxP42TWEyy5BSnyElu3z3TIHolu9KR/hcqeWQ
VChbq2J3QWnKjyDxPA1Uzro6B+SzHWL/NFYDRJPnCzbqIxKNrLI5vJ3UDoX70BlpRBGkyK7KUThO
wPzM/6+HXY3yQIZE6jW98EegYl2nmHXFUL9rMtlvlPkAkXl/GJBohL10XLiHtB//Gu7LOsuNi8FX
sfGPkg/cLFgTkdx5CMGxtOVmtaISOkyWI919dc1sRYs8Oh+f5h5BI1StC7HgCR2ncZIU2bCz7hWl
tBG8tTPsUcOZ6sHVsPhZrO8Oz7JyqliF4wSt89+m7TZl6pSCxPH0Y7tUwxopKo8kfSYU005zv4r2
LTDI3mnVVOHdrHGOsH/yNP4v3iUUsq0jot/HSHJfy2MNS7jTon5bFz36yZt56wGmaSwY0Uv3GaOc
oHz5Hbm2n92BAtBaubx0c1MZV1bMjIR/p7Ib+dOWXOUPQC1Dk8+3h9i2S+FZztFNXLkA7x9uLLuH
2A8F0FNfa5FNxb5Ow6G1vewMRM4wQ7Mp8JB/sxRXsnatOVVO7CHwKbp35WG6iMydmk7f0uO/Hcqt
enqrR5OyNnNdZz15H7WaMiPIriBAO5syCd5SnGP7xaPeucwGHUaskBFKn5SvDLzYsjp0vfX6GG9w
D6VUzdGpoYQCAoJOKcxXjUvGuPDqyDTP9o883mNqEF/NVnpvXP5Lls/T79AHtsjoL6OTZuBPZoG0
pWO5dbRU5ER51D6qULWH5LB1eRR2NnbJIe7PmgPjIf3/Hwcg0Fc06X1YdJmJdtkCI2kWDs1UoWsY
tjUk+7ZCmdAcRcj9RN9iQXBW1H5SjFARLePlV91oWiOCTA1MC9pRKwMsYtNv4SmLALyxQa+k14jm
GjluVXPbeZp0hI/5FyztMxT4XRlV1w9Rv+P8QfXZ2a+mX7F/UfOq46XHc0ZX/FM7O8Y3L1LY5jqy
tVN3sBFd5EqmzNFjmCgoiY0K9RG4scaKr13QTonyn2B0kVUeh8ZNG2/6FKw8TuIBeEa2LFuAXsap
C5bw9FmN2wIEq02yl9eRGsuDqS5u6eDqfJz4yeO4CLOwlR4ltywA5NIae7diO7l9pDhKpRkQR/sJ
jX9Woqv7i2yxmtZWQHVbrfV1I6TQIpogUJ89DD+325jL98wj91blBJL4lAgYWgnu4Yazj6W2Q7mC
cvaVsvKoGUkTfkgFrJ3GTn32q5u8SV3O3gCmlFg8agbax5JQEkjjfg6XTau8dPT2LQUzPuygLh01
DKRCMny4WLFspHv0ZsNKE5cBwom3NlByNQUtPKVk2zE2Fl6Afo7hnCnskvpHIbU0oKZNnxz+U0Lr
oqaSjBcKUbzNsN7kqzx/5q/8N0HsoxicewPPWZGyMoi10ly9uJjMRgBObcFHNbtqgsjLilY9VEor
LUfd8e0URUiV3TJeDJ9EFvPjh4FrPUQLCzbqGCHOJzpkaFihzL6UO7ZjTcXlRF8hGuVU27YevwBG
Ly8Rjk3LLXJ5GLB6C/zpRwH/Iyn8ggTImhzxCOWkyNbmFRPKhYDNr1sZhKqP2kUH7sZFQmVe3lBA
nn17hbPNvMKFDO44Kiy71tnguAzOQlcHEMnPlv/DvRlrqMdxo6fjY9X36+VqeRV9KaDBgBHg4zad
k6GqIO7ds7WLA2H5DVWPdGFZrU1vfB7yCuQd1uuRygGOLLURtEouKeVMXsKNZ4IfaRymnGeTLXBp
HB6nSPvq5EtlXL/1Taz04M1N6GDtJMNAII34UUJPAsFqx+9iUls7VlnKx6Gw9IkrKcDlzc3vHtNS
79GfQ1aArTeawVvYkRZvWVMU3E+afAzWCXE17hqfuvmqNfCcGrZTGa5YYalpnfUdPvS6u9gDUNKV
AVqQ6TQUx6mR6UXV3ZVkyUKTtGICLS4uEzIaP5m+DCZyX6jRomwqJoVNnr0hMZ9ydfcAfoZs45kX
j3fnXuG5OrJKzpMOhTXfS4HS8yr/c1cAdBx2DQxnkYoQlPKSakWw1eRmQSaO8H4zIajnAUb6rhRn
jx5ogZl7zE/lf+3xPHjb1WgtWo4Yi1JAvMVrYXOzxNiZVt3PxkWuW+eUu+ZeowVSLGD+3VEs5l9U
yWOSQ94hYjQ7Z/dHjl+ItTlNeYsuwtADMJUZHQwQK4SkV3YX6RUGiliSo/773/1hcRWllKFvGQMC
Kxdc6thcIGQSE0bDgrsTpz6l+3lCWpqagLpPz2IFA/r6jC1sbrHBAHJQAFjbKLF8vOMm2MG+WwSp
MhJlLXD4duGx7kzfryPd6I0G0fVkjsKmGs9att0rxZL7b3Ced4ZAqBNwW4HXVex02KAK8QO+sXzd
GEr7F+5qJqwGm96nILYiIz47FhjEKeEmf1n4VPlHIENLd18bqzsX8Pem0IZCtWghb1UYGjJubYOQ
AOPwQGpWsA86spsfXFTEMnrzv6ftE/8xPmOvQ1fFZyzdSQBJHo+hXsEBnmDXlpJSl5X7edy/0D9R
jBrNu319hvdSJHiLsbLxiUfgXfhaqt9aN7IBQkdQOaudwkDbzplcuZnqDHu5uGgfQ3t6BYxaTZfu
+LhwEGfUhHGBtP8Ovo48CcRkMWwxP1ALLCvkgT2GcTG+R+ZcUHsrgsBfh90D8bQ91GcWJ72xsYh0
DWWqy37w8MtV2Z3HMcWv0vx6xen8Cby1fcEL2U3qGIrqZMLYeeAf6rJvqzwiDqBkpGKbNK1RuPIR
QEzXKnkd+akXRxxg5ZAORp8JT2C2YnTIa/9aqN82WIWxhCed4hPmD4cwRMHoYs8ti13mHMmVLgxj
Fd+OkWUo575p/Ndehk9D/pXbnnGQrT1b7BhxPMTYT1FupWaemfP6dquhNKAh96amsGzV1KYN7prj
0CsCafbRbZsARomfrzZH+NsHtxKP6Pi1NN3IE5LBoWJKIh+JBlkTqf2gv/aQi41xSba0GcbkMyT8
hAaCj6N6fj42SPiJfjEBJeg8yVjEBEzAFyMj19Pbv8H0rgNEcS8ZNbONE29SzcSnB3aEES2i7M0m
xBg3Pz+ntzYCbeAbkMdOfnpg+uLpUtjvt85KefWDxniVlu+G1j6mez0vp601FR9ce5nLAg2kLtAr
5NdAiHBZ+UzQWHXFmClH7QQUT7BRyNmomBjeSVvHGniqIvTj6kWY/TTJHvy8YtFp1fmZ9YS9dkID
X0ZAHjfjF8nwLzdf6Eq4WXqHS9aM/fEWqo1isbFzGAAFFdgea+CSBqt1VjmYKDoTxXOxDIlK2qlS
4l7/ibvaByF0qUaL3zs6HQOS7lPf7HhtzKL4jlm4r5Td6XgaBq+mhpWPmnb2yiQxbC+aVo/Q0xNA
nUyrSjEApas4F4E9wAzE8g1I/8GfyPd1fhcWRPODGD/2cZXkelbuY5TR+LiNb4wBeJ1Q/Tdjr10N
PQ2mepiQ1hFdMX80PyD3FzkR0DxO4V0Uzt6792GTK2xdZjPH2L8WQlGp6I60vJy34+t4v6X5+n+C
P1uMEHWSbUBqQu9C/68AOSaSu43F2PAPceJwL5CbVyvL4IRItQ1cxIJxwCWH7/vUpyO8E+JQUOIh
gcDfNul+uD49ZI5wJAoECQZ+igMdWfisOAVcw/hxK5KGTw0nlCvXJnyPF9g8qD8mDc7bZt+Idf9u
l8OSchAwyiaBDyeQO3Ogncl/H6/AVI1AOmliC9AGuzdk31o+ExKg50d1Q0wfn691hRFweoUjQD3y
c8bKRUM/rOVlMklBMf3mvxwagCRf7rEikz+IQIBFGvcUW96tYZ6UbisBiJTPTghnOJlAQyb9t7MG
7cm63MjwHY+VWsZ7Pb8WvKbMA5x6GnFQIReiaQSjBfyfLIlQskKHJBjAWNMuJze+/KzIWY1smxDm
NdTwgFvJ0UJbdsCTJnKFeXlf+BkNyG7RE+R2ZZlf4WWDK5yg1kEy7x+cmSp7BwN8qcOfxZ/Ji4D6
7+LqzQVKxrIzoJIvFdWoITvUINcVl1DgU+/37hQ+2zCML9Lk84y4npyDEInlTdmT7fiZjeGB5U3a
xBi5fU19tYEPZFVUZ4a9/4WzNzIzxaGlvn2JDoM7P4X5CX/Yo7cdgpBoTNrU/7XJb7AeDIH1NtFM
SELV+1IpuAuf5/8OrfIfyJ8E44x1laaLiJEV3SsY95RCd1hL3Zti4kl/5OXpPnJL7G2qsxaS5eZR
4oclPJ3sc3FrfYeTiYF5Tfkr5JfDp0LC6TOlY9NvY3k/H3MMWfQtqlrxnMeY5QlEZyiTRPbMQUyL
CWN97F3mBsm6Nn/InD/PHXSJYfujYqEjgDPrprWMLuFR3jM0T8ezPiYZ9lv2lskL6pB5fd39VPeo
Fo6fhUFBBpuGO66pS7rJQFJ6kzSVsF5VrLbaIrTw+JhbtLHuPMSO47KgqJmLe6aOpFc3Wjyf4ggn
p3xPcoHKdjeBHUDhYR5yXSQAVl3wl7Uh8xUMkdiA8jI81kRfgpUQ1iVJn9crcJmQSmuRdx881TgK
cjN215Csw4cxrJJspL2umKJzGWMSSUKwmktJ1jZluPrsqsVcuWEHUct8iGCnVl+2CTwc3SpGjCOq
RxwMqKMGkIt6waV83TtkIlqywHdBVoGEv6jQXey3l7b+xjczbRIkXS84JKvad9lFvO0+NyGO0N0G
oxcSy1P7dR/ZgMOTHVuQPc1ZyXmpu1AWjXViv6mWG/llCfSWv8TxeQCVvS478HdnJ+MV4Icy+ziJ
T68ibZDU6/YecKpVCFtJlBo4CR5NvgzokQ+066Oz4iuxUFTl56XWVn5s9QBT4WzQQZyl2gqxB7cW
TxYZ+Zo0O+aKV1J5oKeXTn7dT8aaFZtDafkRiPQt9Si8wr7LbSxENznQMNEThzTX+GVNdsPs3uV9
hHKV9vVfuUk13P6qquy+E9rxKXcRNtOYtuhwHGl/G32NmWJuzFJCHk75cb7MQiiAchAKYAjfXOaw
u0v+XnkCCPdeHqzqw38Rhw/LVgP9lMnoSPQyehsvMiQ/0k8Dy4mTMu1ZtRzCMRVtTBkX4QIiFqVl
biYje3hQWEmxjiMvoCHY05KorxVflnx2aO0wmB7+KipMMFEURx9K2fQO1E66Wbh1QCXvn/T7WwVM
M3sG1hnauBH+OT3y/pGhM5qCFo8lCCNeda4joCMYgllDsDZTUWktAml1dz/9ltXSDUZwmWqysf+z
i7J0BK5swot09ANW7s+ikMcdilVNkAlNVEgfmiOPEP4GDNfaJ7MHfTSjsRvAzhTmdDDhmfnNrZCg
pNWP5wyQfztD6XEtFfoGfAZCChAm6kbwbRKyPXvaVtHNe8kmJU+DSN7NS5G6gtJGSTbH9dQKPm/y
mseEoCBCXOqPE3gMn8YGsXz0B/WLbvzjymOrc/1SvpdLJLQgKy0ktDd4v92BuO4NNdxP0Js04JAd
1WvRD2FFm39Sthks4Ez3f+TmYf1UKoJMTRtMDilmfrOxPaHR9bofzgIkok94heefT/i825kaJGDF
bg2BH3usDhLMIBJlnebAzJNF4gR5zZhKWj9G7d5XqN2pMNCjz5GV2DkHfv7exBw9fcMjXYczoFH7
7+UIbPIW5r90PoPEU0tr5Mhnas2b4Etyk7dSzKVYAepc3bszVuqg2+HyoUaeg/LHvrHKVmjPQRWk
MzXsjx2AJ438p0cDsegikbJM2pBeyRUDGOqrGiOHWt2kE4nhOQUG+kQN1Tnoad37ti7SKTlsUsqs
HUP/Vk3EuPPj/Z2uFNHz51QDQ4NC8YTdI/blIkclfcKX52BMsIeOTHD4vejBlWlxiVJvwfzthStb
0ZPOUJtMbYzrDl+N4c2Q7wnIXrDxyRhyrO3P/7h/RkHKUtQr6l9ZD7ycOJVUXwTIfAzzOgGnOcJ/
xoT5RWLbv2DglkKuaf68PCtrDhx30JaOPrGfeEkKiibROjNuKDVmwKuKA7gx8tJOC48jscJ4PKvU
VPLSt5Cn4Tj6XYm33NmSO5O7nyhtiZy9cxGPTROxuxRGbf51phj9kcuOum3fNyqkSffpQAJzYq1O
fPOAz/NkHPsmdxc3BLm5cUKM+Zf9hnkHNSf1AZr8PAzpDo9lhe6OZoDJ6Lk+2YlDTWstCUqcNqar
xm5hbi6SspJuiOr84i6mjjQ/eMe5fD6Mx8FXrxe6kmxmrTvU4Oq7zwPDs9EXBMnGBb3ovjK7vOv9
n8p26ewEXcXvGzAgw4N4czZxrhKYcVYO9LQaNO1qOYZcFntwZjGU45bBHJYQazoNXPfAur3aCbUi
4KD9eu5NrGdybn0y7EvMYew78yDhKl5qPEaBR5oUCgXpGon/gtQSQzSpbp2WLCkyQgpeoSojtCJr
PmHiyeExevv1tnq3C1+W+sg7B2qKX/2gFxAkfrKIf7ES1n4ZeyE9VVlSBWOuoyrb851eEdyaL0SG
KCmH35OKNg7yKXeoL/7xn7UJxe7WnUKCjYvSAK7o7+ZHtrkq/ALWWmlZpkYsNl3FH7uweqcz9aNE
aoDQHC27TfPV76SA6zrfS4LU78yk30P9yyTNR7lKyaQv94tv/zSdEU6qEFzt4f+/PPBCqeLCSNCs
K62qWQ2VzizElBnq3sCZUIZPH9itYErzqcU4CpJWEiE4jI8smCIgqMc13xgnj383lhL+MslxCG1u
aIT+xLPfyMOO4RXUqk5xp3CoIzeCid5SHftWFoKIT5Xd8GDFs7e0RcUMt/namN83PpY8ZGgw6axb
ikcKm2xrZv88v2SAAuV0Huk+YJzpTnzkswlc/yST35wxP4u2oeYpurX0aS1qLJ1wLymIrRPm7xOI
oAnL7WoYr5sSBVMsw6zZFlLNEAqveeqtIpzQGQCgaUAVT9G9L5WVDWSOpnxFN+alQ0Hm0zEg5Ly5
bfvZ27E65VvRLucUQxFgGiFwFYASe0emfEuj52ayJND1lemqNbvfYJ1WQKg9vmC7WX21WQeH7q8U
FIZgB1iu39KRt4rfGXSxKyZBTtenTGBgR2CkuLZa3jEHBHANJvr0xzRfw9F9R2aljr8pDEbZ+5hZ
bLTlH7V3yk7IScuG1sm7DHRFiuCMmn75DAWrKxjxgW8HeXpni1JsnHier+C+/DH6jKIAybuGVXJs
/8HfQ3qcHK1lCzL5MPCCr3yGwg0Ty2tUYagwjNGrXdAzoD/4PtIjQA9AQ3JOhHCMniKXavzmATP8
GVoaz3jxPT+fXbnWLWVpo3FvYNE+37n2SwquvP26wygMozvca/saEVt06nszyT2XZ221kMJvcEcx
REbTUUrH2Y13aqfHoy7U2VdsF+NHGKUp8F7DT+AQ+hKVf4jR8TeSsddFnjGJ68UzbrKPRlHf2lhU
lS+liUbFzF98zHjZllKO7xCqrTfvs/saCQf2IkUuIQdEityiwt6MNnf7zDtU5kWwcrSQwZlgl5DS
6hIQ1XIsbFZDQiCV5ZioLJnBEaXIpvvHUwSIez8ZNXRsoO9Sy4/itK7NOyM1kVSRCo3smdzMrQrm
dkJtAiGG7hUxE22IqRN6QO8R9sqRIGQTcX+CStHqCurtQiftc8PeSzZGr/tRpA63MErTBicOzME5
dcclvGT/TcI9nGrdJHuxPjUpgWi3McuD0d/qpYBPZClYte42/G0uLZks2d4B1sCnTLyPiExtnT7H
5nOjX84ELcouYhOSPlxNvJ6kHYEgsXF6of1PbG+DLh72k9mm7BoaLpoKe4At08OhLjayJBkq0wxu
SJAAshLXFTbXBNyBi3Il1dtyXBOr9gKyTxedTWct2RIMLmoRT9xtbhKOzFBxXwE6KDjG7tWL9F4v
hcSBxSvlYR+SgCgv4UM3gZzE/mPp3qZKd3x0ByQF5SAyH/ip6q4T2K8mVSdGdvluwh8MjeDvbIVq
IHXgmTnhjACuVG+2RCh6XQMt0Jfzd/W+lNPkMwyuFtDDLRsBogcXXtopC0hXLzbY3BxLO19RKMP4
qppLwoiODM4mXfsbNOjiCFe2HWT5yOd0UWb8xiP2z38DDVYmFgRQh3bLVJ4EwOHLsiTk1ujKya7H
oxUGEOlbGP79uKGcqvOPOCpXsQ8nictuu/PROIbUHYGmVpQH1aJCkHskm0uGD43OHn2RnOrPyPS4
tAoM76uUViy6xCjJw0LFigsnPiFDz1fNJ6FRhllsxOnKGujkHq+itzSgwpfi94aT1Dxhu+GXD8Ok
Xbu73Te6elT2cBkqAQ/VTQkdaGLCSb5zRamx3ri0MDjYXB0Pa9Fn9kgooGkqPLZLsFoUNtnl8pcD
1E9VJs1esjb+6xj+dKGr7o3qOzndOJXflrXaf7WpKZjScf2OUn5CF14Ic42zsvkiNshoR2fWnllr
PXLoDdKZgFLMUmuTHSQbA5PogIsbZBZsyOGZkPk3OlwFy0ZRQRZR5RwOygC3tmara6cXxkpHBMwb
HsTRpG+XafL+c0tFXk17N+Mw3i548MWNvWq/Foi8UJ931gRcpIVyrzRqZHrD5RZF0sGKrWCj6rMU
AVA22Tr0r21j+rjuAgWT+xBcn/2l7WPH96xwFvSVkfOL3v7lnZanSdLZQghIKUaSbjKjc+plUul0
F5aC1SA+ZkhEpR5U0xE7OmSEbFmO0tEbgBSjb/dwr6ZnGuZRHriSdXIWxDrbe7pnllQTa0M61FR/
T3cobS5ZfxwLaW5fQkGff943WZmH0R9cfPU5AZhslVb20f8jf0426Y1ZVNkUEOSFPVSOcc53SRQY
6uhM4GwhcHqCm60QjHOFj3R0Jaa23yNWs4QnU2K87fXwNYrAGmVCDM2D4AmZ+x9pzdgfZOpEPTSl
iPC0D3Z2+lmGzwW69X/QK4QPBy3AfCACi+yOl7QM/XkRf57BgRs2Lnwwk3s9kY09GhnvzCRj+wd6
QFalsfIBEkmWN8oy459+IPdTnDuGbVBD+frpfhC6pHyQGIZTmFc3rhX9qUsub7rUE5b4pImDh52I
djQd2uzgJYtCogc1k8FUXZGoY2l/cg6vBqt+nYr1StWbUM8t5I10pxTbxGZM86nL0uLwg/Qgvcqg
mNuxe77hKZmyDHN22q+e9MxrMfVFT6NhAy0HJ5jtfJRoT7ZrkLdkj217FSsTogbBNjJumzUynwbK
ogZY/KAMZvtJSZhLt6iRM6Ml5VAxllxViW613h5TnsRlYxMqJjtNwapU6bOV51RH9WFhtjxnHTZz
GhKFVn/o+bu/uT+sjp+rOrBFQlxtLM07qJMaW2BDzG1TzFGl4jE7mMKgokIB4ati9xEIEFg7CGPm
PjraQxC8Vjp57QYKXIH1pfLyJI3RkcD3m8MDXtSnT+WVuSPCu2HqjOQ0N3vY2if3bdOzmWAt1cK9
vQy8i9pGAPieHJqAGglTa/8pXd0PKXQWBzTMBv25YGrr2vxe0tzHXo0OPdrM/YC3WbZbZzUYyNEN
MSMAJj2aKlhRhSEahtEWzm/Xpig9TseEPB6kLWGBUfMoluoQSHOPXzIh3APXimjwnmNRZbfK81Z1
Wl9wlWcmQ5KdFZUFb/PCQHFVIzDZpik0ShClo0aCo/EBUjMXJ+N19Op1YGWvjv/uaMZ5LwwmjGj7
EAdXfkTPzqaaREadkdefykhvzV/h1C3XfTRu4vzrk382g+RbrQJ42he9joPIkhTuz0yxnuGgkNyH
qLSyLFw6Klydj1+w5mZetxc5D6i/obaB3dezQnKsv8hrtf8qmNWyTt3Yp3zfmZYJ4Z3I88ZQ61rv
o7s5LerBIuwtdkzbjyd2S8aMD3CNOia/WPrM/JzBhJWmKCh9Ld3k2lc5CpEV/K8pC+gsUorD9HG2
pw6CuvWDMVTkKSGdNQbXmHd2NNsu4JOqhPmRSUhYy66rLc624VvjxbQRy4CPn6vn8pu3xtq/uFLc
rGw3FdvOBLnkof215SVc9OQpmULSAiOlPgZF1dPmLa3gth4iv6ag0RNwwZIU2kXpsQIEnovDxL5c
PzMsyNmVPaLzT0kO1LHDVwJq3HrOecuw2WdYEMhJR147dE3qLjhnw1lKEG7AU0JZzETD4bJdT3FR
fx88hbNSYvdY1mUwSBv27amtpPBzTG/fCgrlsI0gzS8a8Ry4Gj8xzolAGQpITiVJy+9gJg+6IPbG
tqfcdZLQiibYnHlHhxuqtPQ51kUuJE/dqRERnloRAs1uMp+eDyMJSscNQYxxhb90XsDjyqJS350K
CFnuFTvtpaVC8+mpNCPrqTWbOlnMJDYJY/mOwzhA6cc3/v1tCsPfOImF3BJMeBqK0Nij7EHnPmZC
8i82cDkuXSzTIDEetkeCv/KSE8aCTkv8p+aAv1AtfOMWUYH1VvSMlFtGIEZtwoMeq8W22fPBc44x
fi/wxGuPcnJR39q8FJMNJ+kb1ACsct4BRJtx9y5fBKC8ADf65yhtQ4lpNYMuHS0d5qOPfa39X1Yb
VlEfaCOWA2deEKQeOPmsJf5D44C31tMtioEeaiRt3A6XBuCQdn8IjQ3Wy6WsB0iU0cCraglA5285
/DSPBIea22M4cWxf9CzyineWE6x/aferIdVeQ3mBvBwA3zCGQSxp/6iziqNokO0HRckj7WPaAa69
Ri+inlMLYlL31ihzoC4SDKVw3pjR6bnXcX0o5k58I52ZdNWsCEZniKd2z1kVkI7P6NNhxik50tcq
gSBMTFbmtEGhhFIpDTSkaBl9OQeRVt0scuYgbkITx3ikYjPp/GWj3a3kdcvC6RY3OMLQns5nFsiu
vhdvu3g7UskP0TSKdCLvMJRBcSS1UV3GTLWpGqV3rzQeopK2HGnwuF5+yBikfrLf9rtXb2E0XzBL
egmryX1Cj9tlPCZiw3LfUE60jZ624aN/mOaibR9Io/yZTNC8Y5ut6caLODjLUYu+ZwPCaSkiyl/M
/MvHx9GXTw/7eh4yMG2SgCIJPEZUGi12r6jLl/ugDWNoAhMKV5Yf+LrywAmm7SlPvpz7j+peoiMV
MVKz9mkVvKg5G1IrufW1wvySCKWKFsVky56L/IVXecs7t04LWCL5TSzRHeO8PCxHeODCDICblM47
Sdg4UtUVmUHOgp2twYCn7IyRb1h9j976xF2LJPbwX266KF2kVRMqwF6vvVJEaP1NmA6xrko8A0xx
Ze7UqpsqfhCtdLT8ffrW+YJagbwnudDzO+EfcUPeaX7Ko546xzZtYEPN6+eEFHauyGzdMqTZxEx2
IflflD9oEmgqJTDuTwkRh7YLMLhHXc9PbhfvJqRqVRY6UFlgASrnK5LK29FC5bfu+W9D4Zxa4Zdd
qpew5fSi+ke2TNgY6ySd52+aXAXU7aMIOpXVpUJnZULWSIwyqx4fqMAo/6FppGmFJ7UPU4oj9e/H
J9mpM6nL5wjtQ/oDdTbdcjeho43ain3xHaSN2aHaeAZmAe6T2MvCfiJjbaMaj3G2D1ddHVtRxJbZ
vuW+9vlx5XR0Qr6imtUI6VqGxjEwh5dmsnuvLuiZzspFl1voeu4HLDcSyaC1Qa1uDxUG8Y5aNkoB
tgXs/np5vRjHORO2YXS8jlGrtFKY94pl+hTEgsxdaQILXLhi2hGWql0V2VpngbT+xxB3FpVoC2HP
jcLKmFAw69M+tIk6DOKp6djbHCNXq+MEAZWBmugJMEEQlQkSrCmfq3P/e1LMKqXc2OpOeNJw6kGK
FtjXB4bNpN1ayrtysk3H90HO0cf9S94auSjlsNda7C0Xc0nFsNR6lnuc/tFYIOaIbMyKtLj0zigl
gy6M86kx1llTB8wIUjlK3Aa928cznQ4NfvwJnfI6qkdAGQI9rxtf1jz+Ch10QIOQF5iJ/78gE5gE
azIoFPl65scPbZ3WnD8aoGDj0vxIPdXl+f1lGt3tDvVHzNK2rKVTsVB0JZ6aoICn6deq0eAK3en/
haZxIVig7brRRrAMG8RfSLHWU++0uGKhObutE6IpVx1O4Lg4smbvhbJCJKmRYC3MOdOUD6686/9A
FGHbidR/P6smKGe3PHDVPaKevWR1wz9QGptzhgeAoJ6JWFiXh5fXOeyl4aQl3Aop/yj30jh1GBVw
YIzCKNuiBJ8ALLZphERsyspCG4SoFsl1KM7ItHcLcz9rmnM2jyQT/vv5sLtak/MM6JPHyZpvYfz8
YgWsb+TEKKev6ntzvw/wFPNdfUf6ldZw362pItCmIAI3SnbsF6ortxUUTku/Dnn+T3sQnL18Oh8i
pxGsFxi6jA7+f1wXvRwnqrV2oetx6kNrRXTZHKpvVlfPPe6q9bjbMtehsQGAlewEkhjy4sQ0EWjE
xpFxrExL9+zFwL0EW/P8T1YOKFWvDNQISJFP38OMM3svoi16kFVqG0AhfSP/m++cIVvy362UxKlq
uNG4mTT1HyyIntib5FH4noqInF3aKTm1ABoJinP0+mcxRBgPVFASDZbvlJh+fH2JIPaQLBBg43Q1
D5flD58hax7aHKHL0HtTfLsEDVKJxK0wxApKgayR8dJ7V98Gq4Fnx9ETIEaMvsxa3h8fDPGIpPPn
yTOQF2aGy4pwNyT+a/s4roNvdFBrb4Mqp1PJ+ZwRhxcu8I9Y+5t4A7wLagvkrS2LLMGjL0RA1uyE
mYpY8BGrmRGHujzvnNhcQXl8Xf4rrL2hfTSM73tDpaQK1nwXCOJhRqVLj3AfZlVWg1gEdOUccfoZ
CB/bUMmBNadvO3GInuwCU9YidN7rMuYHCrvZ1hoxRZywZ3Hu+oKc35PQmRrVCI7n1OvHkDKG6hCp
I4BsSBNYPEMDRQkqvpowY4nHSrxEnNZIHZa4/m/hutOdf43/GtLsJ0FHg97fYfppXBCIxcnv4Baw
mMIt8aIaedsM4AMpw/zvXYToxy/synEtETWdd2jIx6fmClzgK0FSQkDepBnUL7Quj5SE3/VQbK06
EacvLG6iMirMzEoWDzdoQmcfv5VrMXsSggX287eZS4qQsEFok0yDzxI2tKW4YT3DnU9eBzHxVe+5
SMCz3h5Xk9NgGOJ4w1CFnrPXzvKyMRdiGk9Sf4bjr7FtP21EgxTBdxs3Isgd4qb07F+FMq9Fwxa0
940vgV6eDkHoYIChnnW0Io9W5wDuqSHRzN0mKUjGzpnMCyxNx+nofqxQtx2AKhciMJAPY/7ekUqG
ggbiGLWfeGezPsXxBbARxnxUH8OAcwiTbe3rzOMK3qdAh0DzxaFbf9Ym5Ognc/suZMLFYuw+mxpD
Fjz7pv6J84VH4EN6TP3x8KtMFBFYpRnQ1/GhyZYs7hExByEY4lSnSKl7QZNEOhmUSqmMgBSRX7b9
QGTn8tf66Fogkb3eUtMVwWpXI3owLPDqRzUt0bcakydfXsvpGLpfIhHf80D7ACj5dRt1riN/BwiF
O50lUrt2Qw8OMX+slpwDC84Ll7F9ljTW5/0QueE32jtQ5B0iOkeS9tpzZkPxaCwHJ0GQoikatONQ
uuvZhgBX/gksJLbj4Mh8sY2U+9Xf4+pMHn4vsn1ru4MgZ30mtJqPZpQ+8sOFHEr8xYnjjhqYPb0U
d1gcluYEtLIOD0+Niei1+4HSW8V22o+EYInwAyH+h4D3ZrYvSdU9/YkLlykomZZOCPAHqNOWe6sZ
qZsGQHBqbG+oOFYsF2aJz0A6LURgrl8t1fzBTjC3ihVXrGgYx+BJm9HfsuZkYVJ9AHxPIxr1Y9TT
SIjRvk13z/rh0+t+9YmjwL9Ar5fSiHBnFBrXCkhHYctg2xKS1Rs9/+aXifYnMQH3yAOntTccAODe
AR1t73VaDEhWid2ptjIFiwUmPzH46vqZCE0FFDbEKhWlKVMnM97wiF/KbAT3pnf9Nt8I7g/BkFJ6
4mOttdK8fLKYHpEhGSpf2J/c9KZdYK7ZFp2fVjBg3zzCzd2rpwjjV6WzjEbQ4uhz4NcnYtLqnD2l
JF2oZU5E9O93bGkCXuSwzI2UlM1Fe6WOqRLyDp4ygwehNWULWdbfXkk//nGtLxNrM+dngWz2oEP3
hKz21pLWxd+e4bypPCLmeoEdNdlYUXnUqBP7r757H/XdV7eai3AKXEJYj86M266Ay3U7jM17vdRX
Tog5QlJs5H5/WDtLkMC5VeEViTdh75NVTMKMjhMDQSnarm5xcexABAnPvgFcHkePsahocu0lFNlW
HecwfNYO1yoU4wnPXi6JaWwr1BmyVHwnQEcs50VlTOt4LrJNmGi0+zqWLCyj5efS/1WbOhlhfgo6
RqtX4ldOBOBeZPhrK2ulj+/SFDmDFwM8tWaqprcjWH4c/eRfaNuaLCWe7UVV+pgbZ6s/scrayTT0
JMgR769uqlPDV5Mhadjai/o02iWpnK1JA6xP3C8Tei09LoJtgC+1ZYS+cFQ7sFvWSmlNqQRJbJ53
hubrOVl/JfhXc67hlWTFjXFtVsX8EWl8b+zap+puQ44yet3HOZZ2ZY+1SWBYwmY89HignYYzPYT+
opeR5nRExnoa1WErx8mSpZxUmoO+XmCyQ2K+PrPBrsCtnSrUyClin5ISvxKozCHGfxpCzUv3vYkd
bJJdBdumstd4UXPLY4HQNbp5UXFG4kQxSUz/LRYQlm9Y4bBDxvuwTixJ6mJGVLVLstZHOkIIxsVk
BIZYmZdFyE8gSnhPtquvDxgtVigGeDH3TND3rCCXuXmhThToe0GyWcehvnTRX2W4PW2Z26yj1ohL
sFWa+kY2DAA/+Nbugb56hvcGzTO6RHIyltqnxLQlwzO7j+mt/9vW9sr8rDjGmfts6KsNmshOmfk/
PTRpUc2uTvy9KeEc5vV96C6mIYBjFaLquhDcwWA1OyjiSjlbz7cuPKRiI+XS6Rskw0yCwJoODEl5
V1rRqshfOzryy0TApIcDatUjrS0SZ+vpcbmE2poTWSTEk0T+NCGnMilBstPGLiY/erw9hy+GNlY+
FvniEdLLMwrclJ+HVGTjoEuSiYbUwJciDgCvlXw/WPW4ZoEf4f5OhQ9tUZTeCiAg6QcDNvGL2vXu
PkDTVPAFhofD4aRoLihrupqiue3dJ13cHwkD/vmfHhQ4YSwMObmhDXtjyYxEcFk5mb8E1/hbUeO/
XqKe7wBmpb1SIjq8bnDlLJ3srxTHu0MwM7FQraW2A/vj1pN18vwhetUATtIau/Q+HLm92yCSjh4N
8flzAU+OI/qu2k9wPb/bCVCK4ZN8MadBXND46E2fLndwGm//YX8Kfx5wJcqlTh7t+sJeEUnXzo9T
ht3NGBCRkElpLwDbRK2cTb/3FwSgpoNY6RQjbbEd4szlWkhEXg0iuvurBkwjRZW33fo++23oa1Pw
IKQZKQZnEeKOjd7Is3xbvW9WY6XHklaHD3OVp4VJB3BWqYxGKvkoJeKJg4bd79/nVyF3A/VOPdiM
ObhmCUbuE7Im56BmyB3RQcPKXKhVWihf8hUgGmHpfPFA7G5lFkLBc3yTaL0KhXPjf8p1XniGVRnW
nf1eFz9sxU/yeOnMJ7Vsx6KukOBfD1OU17/6kxUjtkLTd+6Wusw6CTMa7C8hkmUz7kxZrYQuug3d
j3ah5yjGVO/nTTnRXsA9JK9Ppt3VyxgJzhec8z8gklHc62H2qxwD1iPRy8X1lMyoVuDnGpdEMAqm
C4hTPhFuQMjVG/MLlp5QR1LtwFtWblT5qjxbHYoa8D91TNLquflcdUNfiZaqGLm0CjPBTULp0d8w
2sgrqWqtWoPzoxmehnRNVehgQ4wp/bWJGiFcBNh7xwVAWydrGJzQ3O/IHBDIdqFvWkbdixEWPPVU
+dPseabS5xHAwy0e38qDE6GN25k5ngWezJTsaEI/60lQ5ZiuwISsv7w9VnmqN3IAoL3PYR28SgVL
WNT82hQBOvp9KxaCwv2PHYmnIyK3T4w+TDkrmHiKnNaUdb+v50aAJHP2uvUkFPe086CsGoeQ96DP
lZ6r4ybuChdkehjE8JQNqyGPHP9Q3MKmEV+BIAlcUjH/sAVYcA3WG1eVLqw76zduMyQoWcd2P2FU
MEz1q8NYcEvnJKlXPDv5btz5S1okUiRX6mfEm2up/RAk2+HvYR860Q6qZkIkNsjXch+qahc+QD6N
t1tklITxpW+kNqXquAJaXH9GIMWfa2/trlNEIb1L896HEodmzXoYSkS7LpQu9DqnyMTz3vVGUwJD
KXCvbi2ylV80GtVTt2mK0mXj5idw8xu8VOijTUKFNTYDwSv20m7PSty5EpqHeNfXUuvzjfZIDcOO
62uSOSeGGuYqzbx9TmqZmJgpzZ9FVF41WM509GY92HMwht6Oyx7DB7KvsL7iEcCkpTNAA84uvgj1
6UGEGhnzJfQaF0oSZmXKh8lxU9L+/Ga+FByTmUT82IFDiedVQLH1sLAkqvbcH8pkELP+BBhACOKr
DSvacquqL1a/h47cVmwanjXjIsL+0WL8bzst1KQTfjS12XdHFJEqIjVPe4iEIwF6piOnqAllVd58
SxdsY+8mYvHd232oyu/XlpNJSnWdSr+tUnQTue4ccj50pAMY9X2uyuFs4mXWo76w7BdvdiZ8PzQC
KBUeioug2bQeTuMGkh+xEj54/cOdskXyO+Bbb27NbbMbBk2ypciJLy722Hs26aGyVfaFgnql3jjW
ezlbukMY6z/mX08GW/wIl6hjzfexp+J2WZOG3v92IQkhU4t0F1YNeZh3t3mZz0peC5Y1SQjfNuUZ
Zo9WsAvT4rv1SNWihcCSWCfmevFzOPxpKfUOmaqf/xA9t0JSrsvCfiIfHAfMfCrWuqgqdmpVyt0F
qcwkVNgSQzaOMrj5rPewYL2nZkWD66Kf2JVEJ4qGnDOwJsbPc4gsjwJJQYfws4d3jx5jviJ26z93
W9xAx8GaSsF7ah+4hzskHTPw6F/z9MwpV/Dz/tbgKiU5HQQjUH98LnuGPpTYnt7JzEC1KhjFjWK/
LeVzdicxPMqxywiaMgpSYS+VDroKeMkzKhV8bVd4P5vzD/YB8kzk90tVmjoUcMXAhY6zT5/Pvo/B
UdjYIdU8eAZHDVUGVgapDvLG78GfDW08YjxkzFWhulCP74dBwIVShQKyk5VOQbdE5Hxpt88DZriM
BOZos57W5cdxwDk+k1Ugy4CD6oSP7PAGenhjv6W81g7/fZT2OE0GqOnTIR+1CtgQLeqxxdERr5uF
oQvYUcDfNj/hUS9jrXHiU9f0cI8f/fu6pQJVas8mNLgR4+QFBJPIJV1hG2u0ytyttDYBcZbxBYFn
IzoacXh/KdMbG+oPJPI1AA6Lj3iAqlQElZ7jpAwEVop0vbvC7qWpCotDE84X7TlWMdE1KtDvMmXR
6NDKR6Gd0KtwnShM6lIx3gBlsazurlJ0VEO7cQTdUbwUVpzCA/33XgXK2iLevFD1QTiLO1bU9/zL
NafQyM7w2JCalC8PHcADmlBYhXETNPiVLRrjyfH8x09dZV6Y3C9XnCMv36bXwtV8W/Q11Qo6HARu
e/2wEiK2nt4NRTxnS0Ca8sCB8uzMXqJAilIHUZZgaEFxzQzVD6gAQmH02V6/nGNYPzvPogrEU3dn
OhzeT5Z0ryo8gwcWr+UnPujVO9cQ9dqmkjTZdI36qenf8AKnKrHMvO8cllDoFP1/ZkgtE3rFOcs3
obrdj8uEkFjxbtx4VbxopOIsZ0FZM2PxpCOysUnCwgh+z+yRG2IMJo/+tN18hc+ND2ZA2FnJhEec
N7ASC/Now0I2uim6chHVkEFBFU2VCJRMoyLn7IxikLIyKAKn+RJhWcK6HnSMNstbSEsgrAJMKzeX
tLM+Y7Y72+QPnMIbu9uQZoLJC2OWVec5fEPRa8ED4mT330GzNvGhjqoPI3lVakFhHYL4tOyzT02Q
2YbETJdds3fFM0BKH+RDkg1E3v7ytTnJdGAeXCjPrx90qdfyp1MXFRT8G6gnxm2KOyyxCKTaY5gR
Pwshcap/tnreLcadysRc6X53ll48c8YJtBGdmdRM2zyPDipUEy1U2W4W14TfCyvOmadgYyiyET8V
dS1SXGakLoMFsbF/EmcQ2uKCbmphfpyTzeOrmM3DS3+YTkkUW0Xn6/oQuxCAguh4RBbRjHmGRmvG
gzWuf5iKXVm4IVPXKIomBUl7b1SW/iZLT7vX3Ly4l2cEd9tdcdG7hZF57r46aTpdhj7Kfsf131yC
SMr3/DaHuznqv6Suc1B6qfvd9gTcVoY0N4LeKWKUtjW9X6ObW6CVaTAF0xNGC1S2YjSRgej6CMLp
77KTzBXVIHDvJl8jqtdk2P2oIRAM1rHHN4S9IFy9k6wUpc9tygCacV9+54OJ7csCO3vU8YMNntmr
jjyXIjMjcyAIEFWsUT8mrkXPQjorjdVy0hxWZYoulMN+beC/U09yw1BLSq1+gYZViyptEk+L95NY
c/WHw8d6LQDv1fX9Nc8sWywSBPmS1h6M2NBlN60mqxIAqV+EfMzl1/X3lEyFkxXumWJzUkVFWY6e
jjuTrBd9rFYDFhe4HNVg9DeuQ/jRhU0Wfk2S4R2BHhUsO7zvsByaiDXY4+vgmx/RMEHzXuzU4eT3
kJhUd224bJk5+poBRgAJugZBz/W6ILJP7FJt/yOwYwhJTd1wMMPvFPDGjQJjGBae8Ux0ur1YpdeK
TMwM1FPPP77TiUep2XDg2uGCsJb1nfpz1OCV1j/4KfB0pevlzwB+iuY+Is0bYhxSAGcWTkojXAXd
4LEX+aHcJkiZ43P2RltfwXQjbDk8LvBRhje8RJ78GzQY3sHBhjCyMVLh6GMPFiTzbQyn662cd4c/
xfQqsOSYa7v1byfs/Gqfb+oa0CzgKmArRZHXdz94qhg5i+IkXAJh5JtHKyj0DaVOHiV70Ay2J2yB
M6b36ihQAIJNLqETdYifF8bv6mJ7QGGPWl0zq7BIb0VirGP5vbQsmd/YD0N3P74Z7/8K0uLRVo/c
G4Cq0GHQv4n7qkb4CisBmialmb7aGwHEoaUSgiIbWpIL7F/hmza/I4wkLXMKoX3gMsKG8IvUbPcG
kpIvKS02KUIX+9JXGxFHvBfK6VPyxmaM+uvJhgxs2uR8FkeGIvrMcMOHF6f+C1vQy4KwXhZIRNqN
Vqbf1IkMIQMyd9p4oT6WpWXT3ndd4+T1CtRzwHsA07toPh5mfruRbFvVFViNqw2n+RyRz1XYB6sJ
40O2Requ4dY+HScxokRGxi05ad1SLRnvYWSL+KJyZm/ti9MwWya/QOFhY/CuFC5dA0mXBXjLgzlo
A1okcUDo4FZK/PoOWhs3oz49FWgelko7Xb0GNdjCCQRXZtkOqhSVWrgUMT95QLNwn4znbZy2ZrD9
l++8/JIFdJAfiSGu9WJ4d2NbIdBZybl6l5/H27O/CY37Ag7RyjxjSvsZ8r73U+hCP2zmbjKrDuSp
xu2cch0bsbuoz6ZOrUjXIIxjirnqphWHN2hWjzm6znjCQ0wzazoeWRpBFrPtYIFTkF3QDEFX9yR8
ag2qRZEZ2RQvCPQizWd4KVlt335VmPO0ocdi2+C9SXOUhrNG8pe2uBoTMGmQ+Uix2gqbFH8CQEDf
5knM67dmvkbqNMCArbiqDUOwSDTL1rTeeKbPVi8TRPEGjGCuO9KFCY4gxB7MQI6UPcaBHApuy1p3
ccF0vSY9ZXAqCWyPy4EtmJTcTWYhbslMMZRTYVxBi7gq32UUtkG3IUGxWENdZpqaqQOy201UMe/0
7/llAf209DnyZHmd3GP1RcMRh2RI/oIWqEbegjggicX2TCU8dHjz89J201rr0UIqOMLTGxFld2Fs
YMXMmsXkKiohdS5TY33WcRHcbO6QoZ/9mhTCreq4QR9pPzRlg4ErphkAWObQB8CU3SXGTehwM3ab
sh8Y4auSA/kINaEjs3poC0Ik5C6lJhtQDRgwQYgXCn1at74eHBvtePlWOJGSC+yX9Amc3DhlD6cX
FTin56aVpse3HYtwhLv6WoXHASw7VX+waeL2Wo2WkxozliE++43eh5a0OlCjEPzoHTuLCieTshWv
VGPiNVGz1x6pxl1TZodvmHykOfXRzqUNrkuL4iHU7j/Jxou4MpgiA/LroZKt8WJG7HWQQieXJSXi
raudKOcaPs3q2TVM+5JqF84NtJkdozevMGH55DN1DhyKHQmpFPCCd3MaayVXfCOWzZqghRGlpRyF
qud/sahdq9d6dAX/trrCC7mwIvVAVoEBrdDhaFCsxcrNaUcJN1u4fjkzI3UcL4lK16avCx85rVPr
J/iswSR6iV67nKlbN4fvyzkBOZHF3IifjmhPK/YrK03k9GYYShi0EKdUU4g92WIQ5PinpZl3MQr4
+f/LFWQzqSC9ND0ffW+VFjl97/nHyvjFbmktFXdZJPIlq2d1iDAaievAy2kRlCBQkv4JNLvwzKLh
mX/AopEdIGAiU1LrtcQgelA5hq77TgnTVDc6n2sJ3kJirTgCQcHgyYYJM+RVAUud87U79FsFpKZg
Xyfh8SEulDqCtRtRrpM7KVB2PkgFhXpOeYm4ZMdWAzV+3YPVuep4pTssyCbxZ8/L7VXh7Z/c45OF
r2vQRkKgWvljTJMwcAtXP3BDfkFLfusH3vEQYR3rtMwzwyNYxttrPr8mmanh/M7TvMlOoPZJb4bP
WhiWn89T5MKBCbY3qL6nzrATBqzmC7nlW5Ovo1Otc06u9ZuD6joWj0qouagGcwwqCjBZznDCd7G6
aqCBEonsUC5O6h8PNPu/ZLmpsJRYmtPad1Q26xVQJEoaurd80j7Isb4JSDoYquUcqNUOZJAXs7K4
1lCGYUndyGBpxTzC83NMFmMst3s1GLN/BKIlIxUu1mepCGel70F4CK8xmsfiATxY7ah5frr4B6Rd
bp3pjfNMVG0wzzchq8WMplPbtvrD8eYkuVDXOiXild8oME5FvpBz7N/jLXXX7JW5JoUe6Ojd78YN
t21FjcGAkwqOe9aLskwOWY3rlqkt7Vl+ohuxOvmV7r9UFCEk9e3SZwPTTsHj9dVrW75pUVBdO1rf
aLcS6cm1uk20VtsHtUVjAi74p3LwkA7y8CaXj9Gf6GjXYFPuuuuOszTdb9jbk8Nqgoc1AFLAhuwc
VD9Okp63sRY2BwWOW9D2Do6xbmEcFrmci6cyOLeMXkJ14pAK+G/2p/1yat3rR1N4GMAQ5dqld/NL
caVdK6UMSvtG8GZ43gqMMcLPvwzmgvIS8UzQjU5ZOUws7GcEy1dhQIMoc92RjMNX+eftYd/lHtfs
iEHU/uRzo+LQ6BIdHNzyj1TgUDStjkEJUtkHyCNij+69yzsaaC70eqEBp9SCBhvY+0eOKaYmdhHT
97Kh5iH3J+Qot7Ih6EljRbalZV3pqvxm5xMqpmreVdC0Hybu0MmERPHrKfIMgnXCcdEYZ0sI9c7h
25O+hL3dRTH6Oiko9u73ZmJ58R8uwvgPinzZhHOM4lDq6lYBa+H2p7n7JXoVK00E7/7ynsmxZtRz
YlxQT/sRz0OfyJC51SvIgv5/Z9nWPNUwULzdx9+GitgYWyvUphjrrzoASInCAtnQZvFYRkX6eQdA
MtbRh9DZ/Ib3Lch6o/bazclwBPpa7t9emOE0Gk5ekXPUeQwVR+6zmlHzPHK/I6f0kWY55cUbcfcK
dJ1KJTuJYJBoklK/JdHHcdKZdzANVDLXrOdaWIn7gIbyLce59BylXSadjsU8lluhPc8+rqcnt/3q
AFBb8iZLEQCf+bcosba5Sbk+OlYbUF9OQSvbloVfg/FnnNjSxvmE6WwIYlYE3scqqetvegfPiuv5
NiPaAVwi90YeQkuitiOm7yDaFHY3yVRW4RbTtVJpSY5cEsUERY5vzGC6ECpyzu+Ih235LHUE2EoL
+NdPnXOAGq8F4m2Prq9DKdNOaYwWANM81GuDEajlS2fEZq8t5b1nP0mYgHR+1uRP2rajNNFsv72Q
K0r+yPZpbmh/ddaJS4NPCJQjYOKkcnfGMWADHJZYZIpXjsEcYvwP//vGjic9X39kLjZ/5TNYKn+U
YnXVunV8gCDP3tq2q8zt8+kkVjns0+N344qTjj4XIVX9xfFuXh8y6tHeyjdk5CohdsqAs5XZDhAf
PLXMoUVi13328vSNRUYSScG9hLtSNQTl4c/vFQhtPUFc9aDcapH0v3felDSeIxVfsqFJdknXVNTp
CGZ0UINvJ365MlfppVGzz9dVG+A+Ip0+5M7ffR29Zt8yd6av9+KuMSOua642NGhG5OWjJS+Dgh0x
faVCGySrRPcbmg5KDcgK1UDDFN4GYtofjEU17oEyiHFTdqab6QE0Mr7i8/rEdSVLaioUjc4/EG7V
w5dDz+FTIA8j2lXadKNYRQ9r8cDX+CY6ccGoNhoP/N34fbrBqxYKtpHZI88QGFieB96PX1kFa34e
qOwQaS3OLyLy/EjuKx9myQ+YDpnJSBcQslfTKCO9sarIc6bR947tj+MzYnXoiRwvjE4PT2idBKtU
4dW50TWw7p6YAMvVEqUeeZMetbk6vNuAT8ks8rocFwif5yqSq7SXSMiYE/oOacsKq6rH4lX1no/R
6AbNhgTRpZ6R5BW7ndwtED36xkc0iYtSMuqn+JoDy70FDsFCVZhSR7Xq3cr2SdRXtJCSiD5cegHz
x6h3hr8H/hiJRgc3/CgFzvNsSFSJorsW40BHDQ9ckOpThHeDnNhQvohe9HU5ZDLD5Wd0zmCppL4b
jPfxZsvBR04qM7C8x25ajPyshrNN6kLmarPvl1fpydq/tsxZ5A==
`pragma protect end_protected
