// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YsK+8iP0CodZ3duJp18gM44DfXiLNiWsLwo4MmG26IFo7wAOn49w7fw0tjlxGCIS
crnBLXjNWMoHBnvmsRCnIA3khYyGIOuoQVFGGFHTwNUyeFDyPrGB/BWD5j1kZ4J8
Ux5VvH/CfjA2ZmNtRZnzY5KxQ1ZA0Pc7hgy8kw4SDAo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10256)
6xQB3ocwtGrspqrI3GMAifmawxtzARpEFIzlFKKiT0TaW3TplRsw6p+eUPmX5IHz
kDtR110ak/5qJI3xbR8YOEgrUAxnH8BmDhfkM6q15uW2QUn8lhlfgr1a7RU5Za3l
GkZFxYB1B3jChVIeZBzdbKOsv3iUJVkhIVIbzU3oGNdpyyjZqFz0XAJluIrJ5uJv
JW8OhbfHqoOtaZBxPRLNuwdLOMUJCZ/BPs+PenjPj4x8XGXnSIivvYYA8BOJyQZo
GzgpVppJLC2BdIwC4WiMd+9PsVrYeYXo5sKCOYfq6M+GEVeLRI25xxFm7mQuqme9
PFn0Glzl8CHI0ge5CiBKM+GdRnfLinbNK7t84XbjzVZYsR0w2+o7UU7BUDAZzJcd
/7941OQ2yWwEARG6Lipq6+SHeZ8jNASMK/3tC7mPC09ntHvNwIIO/AuX8cn6/jAH
+CKS2KbDQl1kdHaHKitiJ45/AhYNAweIYr8pLGzsk2YnBM7DOjNBKg/YEpPkZqyK
arWW2ylCiGsN0BITCgYbWXHZ9Az+b2TEYnZ91mWG8M2SGt5ViVi65RUDhuUZiZSM
PTU8XQgYr8Gc1P9pf3gwSO/D9II6ifmac7HAbrUJuFlxI+rJoBaZVsyEXKw1/16t
KjRALvxw0L87C0DBm+ocU4BoeOJV5sD83A/IZSuwB84fy0mWbkc6Wdv44mNYxaqw
9ZpncmdO5K5yqTW9nyK9bvnxntRQOe+XkIzBtUvWcEYCIZxEZ6NyJpQ9eCUEPF4z
dej1A5JWDpgEsMCd0xzv7hmRFvM0srPhJWUbXg0uKH+3uIZqEro0ujiPkmgOA3EN
lcP9sQk8a970F8kBzGmm2cKH1lh4ULJPHjaRTJl1PBospRCD9H+x++Vo5SIzpwpA
FtL/0zBnzsAV/1JI/vLfTKJKi6hSIS90C4kfMUGTEo7+rir8qSQJRpHmCp01m2l2
+j9y/W9Tf6Ue9jeQyNg5GXrfsk82J2JC2NUH4jJHS4uRNodMjDYb9vnVDDjX9gGC
0v6en30S3906J2yw7uuTPyXKJDehCN/8xjr72ZSYAs3pW7Yuy0XFiKVQlWEE/BlC
c1KicdBK0ziohg36wuvvspBcBJgYVM/KG7jNl6Ar7fpVFte+T3OgOjVoer++ZRTz
AYMU5xk1NyW7FKBUucNk1Zh0yaKf0sDqVTAG+gxUmAUnts+IzpKfLVLM6diz/mCr
xO5fIz3QpZRNpz28aE7MnpudoVoSGiJMOuoMdbOs+jggFTVIIqAEZaq/XpAkOKw4
94syKu4mNfD6Fd32tt0Tb0KBGeav3xQ18L+m3Jy2C6zQ2lupZkNtrTgaBY/a8f5U
21VbEDewNaaRoBE/oO6X9JE8mp3tFnfDonXt3cbvfVqkCcuQKilZbvYpfXCQmtwx
AMqKWYUcMEqJ8/UC+h9jCCPqiAdOMnzkAwfV8Gi8Z7J9/lVu+ZUXbF7QxCAsBvS3
b1MSi/1WD4UFbVVFiFDcLXWPpIit1kWbLDIkIjUd3/hwTB0xsjMRfDkFtGBIz9Yt
O4A6sPgesbLiloiA4+nssndNj2UCzs1dfqf0uHAkuxvsjt1C4yK4UM6QAmT3iuwF
++uMqWEJyCkvF737d80Y3YT4/ubvItKowNyD4mIykK+iHCI6AO2s/bNAq5YYSL0G
H0IiLEjvr4O/WW+lM73lKHdt15T2DMLxt5kgY7vaTDMLKjoUgA+94Y04I44Q3TBh
Xw5OByxMyZnxnichQonFX/Dj3HLKDHfZGzV6SDxuqSUxjIazUHWrUXsNuB6xSofQ
kTHlXXEnJ/uj7UmWu1PrgSKYvAzQi2zY9IdmIfVyjlLDAxH2++fx62hiklBS7fL0
YEcozmOZjuT4uIBrnBn6mucICZyQpBNqQV0hDQdkp/Y9xqvrg3XmYd3fSJ4kR8bI
Mmc4KbxE8OrPTu32CbQoZUCXl73LYKDj/zfE5bOWD1b5vOLFKFn8qPaft5CDfpTd
9XpdLGv4hnJHzC//WQEyWwtNd2CB4yLArZB29smdjri4QvHJVf6MyVkbc4WxICGi
0uKbJFrvCSyXCtCrIbav9Sr8nRNgOIzrPL92bw1pmM5OpY9teRa4iRd1OBPj6wcP
fWcnWpkfKTfb/LWInXMz4r7/9IJsjFHucz2/MVNvQJOea/5yzbjl0Cm+S+GBkYUE
NJoZgoanuX0s5guWdmjmrF6r51Myl+V1EScT70RRVXY2xfC+niv6ECMI7vMI4CTG
mRcyaZ24qCHDv1zapd9Cx9OmvgY8HCvU6ylfWHra8X8rzjoouKn8QWvzSsQoTlGx
4QHsqLbbk9TxWLM/9MZoGI+xNPHixaNeLd/yhALNp18ot8ahQOCOIdUMD10Na/Lu
KAmhCKyNkpaK8NmKOV8aiBHUPHJ0eCCCDvMP4S6nF3yOz4HkmXq7GFV6+QSAhRBk
VFIaLDRoCJdofcOwZ8nV3cTQscxN3VyAdOpz5yDRyDPvSClXT7JJBvwjROwG99AU
9/1EcWy91fGSNiuXUGHZe62XA/xXTozJVyyQpPKPMd4dQPDB6wjeU9L8fbGW21hb
+HZHd4641q9rSrieSl4SSvVMQABsS/V2W5bx9blsVxzEWU+xlRotOIryb9tK9nyH
ZDzPJwYFRDQEZVF/VmvzGdj/8TqynPeRAo+cyGrfFPvyVzbxoF/xV9wpY4VbNXMi
RCUi7V1yM2izPrcH/UXfsyA9vJG3TdwF9FKFK5vgLUiJTJHnbTtP/NoY/nvr1q4V
98bnIhSo8DtnPwX/kCwo457/2XWhTsIZVmwlV3LuAdFC1RVVTS5w8C/1aORGgegE
e8mFQZDgR+/n+CsXad2HVyIaz6rzW/IQozei2lCrDSY8LHieHf06UK+20oonahHU
nEKAUKtA1VFpzYZ4T3sddM7gpRlM6PwY0UKYQk5j94ovVWugsctGe62rCjzduz4c
PGqAeloVjuldLNOys0IZrg3ilTWEiVsrItC6+qb0WuqRcerxbV/wAkXnSbqJGLoy
m7n1Ubw9PfCbZiHE6Z+zE8Eu9/nAQV2b7ZxA6bFccxcczSZg1e4R96U+UGcvwMKH
kSJ3UZP55oqApac1W1F/dlJxeBS3kc8qX+oTyyn1nMiAwD0PRyWeILvaM0Lr3Eqa
fOXWIviz4MEF54ubfDKJKusq5JLo9gyV3i/Pj84ykYr91Z4Ybro4fM6lACJ6sKqv
90tXxnTp/tKNqiBtL6tW6v+yvf8gqEdoI/A1gQzptWJ7JBeOIx9TcoDbluyl2zpp
AfZSoBpdJGCO1LE4PVljQp1Gmdu64/q7Nab2iMJmVtamWLdwOWZ/cjIYVIpdGz9t
MDR4GGfs/SP+zXX48+m9HgB7SC+B6DRbnz55TvsE57OQW8+uSZEj2yDvEetZdNA7
kn2y3dmBitY1ZhnNe9fnIiVbZQchhuR0P6x2j1Ufsz3aQFfjQhSkjz6byuK/+wdu
r+8pUiZY3OgHk3/MlJYpvfQtOhXLDDtdm0HjTL1sqlZH2ycu2OPXA+QvLyHahcJZ
uIGjF0L4qtdmuFyvUltPzD+7d4J8kzQEb07n070c2qbvodglTwgIQKVo0tx/g8UR
Yr4CSD9CTZS3KF1ORZ90jlNNY5kx3bKkPrRx1XZbyF+pSYL1mdewbDGY9tnd2F8t
qV9S7xXku/8V2LFRE/7Enil0WfGvMOv/9jghMSLpKq/8pFLzyX8Nu1fZHan/HQz0
WmgJ1biCvU+pw5XnZFpu/0XO/Q+H/ulz5J4OInBW6FhKMzRIPfoBeDoB/QyPpRah
mGIOs9Gm0KOJX8Qdljk+B7BezuPuWg3X6jWU+H6m8zLqAxkLMeJKj0XK0slSiyFf
bdC/uhn1M5J8DeYpWm5CXzZdLKfkIFJnEgqy7Ph9k5WUD3/ZtpGHzryB/tazmwlE
bpAJ9ahGmQWy7hCa74zuGJE2Pj6Gh04MFzUlg7soLYmrauBflqxDb+upvWPZbMlD
5kHnnnowVtc5fsEYlectHpEnfsbxj9AnxJzlaWqFbRE7ZfKkCCEd+0A7ezdGT7c6
HSHzpdtidBoH0tKCjy0Qn83X5vgpnAaE69wXSjs7vgauxuimJZEhKIRN94RHU8oB
PWjk4T5Nu+AOsPWBfSjI2AoSnj/dvVc5tEOAgWAtrDaOQRhZa+7ew8YaJeQih07C
TfCCUP/C3Qxb5qX7bQ1f5nDwVAdO4YSVJFOE0JqAGJCETIfTBupk8U7pXR12W8/b
WD3IEbRxvAH1k5/k4sgd5KLHipp+m2QK7xb7lD5QMYtCzcuva7X7i3r1mSxs3Esu
1IVJaQxFAX/n56ae119QtkdhCB03QsPf9npmbF2Y/hdBPYfvWuV/US93QIx8NYk0
H6ssKNTYI7PVo5okyu3UTeG3Hd3hYCE4zWTxYqFCvslxGOZSzyUHLs1ZrQcI5/S9
ro5h0kRDn0oRlGePhA+MYAe9LgxgZkoMU25v9ZHA+BwZDxlh8SS9LwE4pmGMNkE6
et3UPx2iwMPfjmF5W8SpSI+j/F8bXNc6hx9lEQbmE7eqipdDdxolzbVZ5IYWYQQn
tRx4cmB/EUrFrwVI4Xa8RiLTLhlKwhmum95bhMo16XvC64Ky3LS7OnzAGOOmcvzA
wJE0THBERY0SIOPx+ghXaiWXCKZ1jKKqJVxkDTuuLNZ8iTwVixtKSpSPTg3uox4N
qsMwo7DXcgPlaIFz5gBH/0PKpQGu3KVoi7y4nUwf5bpTHi0b80n1B4H8TApLoFm4
tCCoIa73azjvKL4/lvfj6wNw2lQxpspmuGMHlknhetqYf0v11oO3AwbvXWgecwuE
KowLzZvMO2pXmvjD6Mq1FQaBvfLCX58B/J4+3SsMOL/s4wuMSK1jMHvtE4c7Us4O
Pm91cPrRJUO3ZLcyIQNinQsubGHa8ht/KVdeKfvY5soXfpwc3lmRwA41DkNttb3X
jZmRfF4tJi9nUrnDZiaJjSyirg0Ax2MVhEGSzxtprTGeLNkX0CJZUqCzZZ5j6/3f
mw1drfNsQ1FgwbLpFT6hNk78rX8X+pQRzZ4lQh0egVQJylMmxVVgA1NHSlpx2jAN
QNt+atlzugRWxTEjc70nY1yWQsB/dDZT58EdrJHcLpyYQ9sjvyUbD0oW/hlUK9Qz
OOYOo4KqDV90A/G3McuvysWePm5gujFqlQg/SMvbDbLeWyMZFEGybI58MjCgo6NP
EoeCPTZ8pJfhUJDrLc9Q3KWoR/H6dpp9R5DveDj2EJX1tUeoiJeeqNwN3KpjKRf/
QsfIgTN8J2pi4QRJHEDYzgHodwDS3pO8teyb5ruUz5LkBSbosSWUzQDk9H5GqrLe
lF6cCt9HkJePk+NGfG7nJaBgNUWUc0PSfyEyLktLXklfk0mQLxpZrTvG3jeqAgVm
4t3QsQl31PkfZNc3cHtwhqhZ6qP/RtlUyWoOQVQuxXpEqhxBUXVl3byO5Ao1d0nZ
4jTC/KbaWyp3teNKwYlkRjQctv12sBX42PYzkpVBCCIJxtBOUCA1OVCuoHCW1+qx
0WXWvKJRs8qOkDFfLuNmUsBEYRguO4f1X2Z7+5SiRZ7bwQR+X833+h7I6KWI9RLf
NkR4ZoEQkag19speQpp/jmfTgyDMTYN/7Iqpe+4Z4UInzm6CLGBG/Lauf/6o2TCa
kHprzHa66XalcP6A59rICrVmSiiOZx1lmXEoiKtr/95SRGwncvAX2zswRwvk1OOE
pBjr58Ck1uwQZptt3UZpYHv6BrZX/2jJ+x8OjYXgXm+mJeM/Iw772GABxuSqvVr/
lJCvya5ZcyJhzEHSiNVK6nLSTaGnyk7XfEc9aAZCST0bc+wUQBVXE6KH++4seWHK
tQXgg4hQUBPwxVhfjvyIHFQEaphm5RmDPY50hxXwF6lW4KXut4cQn6KGvoeSwTBD
PRvUE+CMBQaNiC3DGdM+AFGsHTR3vl5X4rgxrFowFrd/cjRYdNpOztJUUgGFR+zN
XujTmkUr+MUBdT0OJ+syrIWFTezM21tgBehcXPjl9BG2ZvgR4ki3hNgBlK6y+JtJ
DjILibjKuTaQ6OZsOZSuhDKfYNtYKAT5vAbHdkr+ABxw0cqRpL8N8DSKGsk/W6R8
dBpgAjmbQjtyvfyhVqew/HJj/W2vLTNL3FrC1U0i2c0VE+fIN4Z9rS5Q79XRdf2B
zRVD/B7TBcoDqWw83frqwDw0GqJsJxHnpCODtlOZ7bE0X20/sw0NLfhDk6TvOt8F
hNtcNGm9gENV+My3kP8suLlbqkagT5f+XpnluVdBi7Myi98fzJePN7L91Q7XPuwX
y6vaNe7otlr+WshENvrkjpYW3NWTWx4uUuiw2VpzoTXNCd5XRi7SLHY/TvIcip1q
C8FoPYO9dlUOdOZLowTNH5h+A2EFvg8rmlsB9TxrwY/CE+NRmSQGdJncCT7e+4wy
PwdF+wG+cEjyGhj01Jvp0jTbZU6bAXZbiQsLJiHDGeKqevIn+vughN6My0mHFstI
T/pFEppj158fCs47vMfXloo0RLoJIg7gIF/faqRI4bnd5gD+1rVdOg3cpwqF6Xaw
GOVGnXAQzdz6TreMOpgARjsH4jIZoIGOSSv36SEqkLyEyct5LNkR0egfYqFLgDRd
93K4QNXb8xsVNwSYqNFGvKm0fFmWnv73ad6cYMnADPRh+thxW7pr4MdJgJkdsKYE
bGgwk+OSpfLY8dnnlARuZW8H1/jGdQeMSZBI7Rr5kRjBa68+pHg1HfXBbERAxa5Y
VROdvStUJ3UapMei3+AdSxJQ0Z8B7fim7tLei5A3Dai+u0YiIpFMxw5UHo/cB4nN
Gh2V/Y71Nz0aCtqhZ1wmDqj4mOUyxAwUcreXyb5QFFgjp1OCBumFJzbN51cyCKfr
EIhr1yiioye1cm4TCq6eNdocjnOkExfuq5lLDGr5OF1emSh6Sg9wXpkhA1G3UXRM
bEYa6y5rGcEN9FS70IO8iDBlmGKsz/Emo5zQlj7zOPOtC3ioZGQ12ClXhZ16ncp7
XLM6cJ8Xakhorad62T5eX4yg84eQ/CS38l2PJrDzKi8vGCIjcPs7YPrINDV5ns1m
/ia5MVLZLU/+qI+Lje2h/TkWajMofcz+32nkyfMjYkXkcSoBmmn2nK7ie+2xlRgn
icdSfd+Uy03twP9bvg+vujYSj5X6ct2VcJJFyN96EaD1/QBhyxCi6eqnm8i4TTJD
3R4PinhztlYGLB4L0TK9PXNkiWWs9Mm0Zyq5EOBZWrk+RB544XGNCCW7MqJKVkaH
4SHtS1OfJPDvl6Z/fbo0BEhtR5yyftmtlAa6/h0TOFE4xmvLsWRSnOZq1lY+4gjC
kaCENyD9ayhra7Ay4b+yjAc4iDFMG+vvt5kXsGH6rHj/F0BtTybeFN+q7J7lZPij
3lmKwcvW/JoxshTW0ZZAE7SJrvGYDAvFEDl9bj76Fi6bihXM0tp5ejtMjklw1Mtb
jcibLjQlw1LHt8OJNBty+jWbfuYZE6TZ6Zb4YEegToTPXaySQ7b5WYv5vQFQ3awP
ZkTagNXuUtBrfKUWQnjpZqcK2PugG0O8ASvaFYa34ISJ7v/wPgT0NlRMm4D4wSK+
ErQlg0NLqUQSEfpp/qwe2d+TA+LzvLiYd18LLh1p0emZPypdpp4CyO1qyIH8GcZw
D1IibbRMv9Xao7wLWNwpZEfFTWkdCbqoYcmiizWJ9vwpHehwE0VYPTd0EeKaItGX
UU2HFDYAHsVx7Pb5FccdezsupxmowDNyt9IsDZ6UB2weEY2hzEglGf2UwXw4IvVf
R9omjUBOGszkE2TbAUEq/1McaGUR2zGwbDpAQzm2J1NvjsPvRaRBpHIDeALFZMdA
6zGy/mI9K2VDGVnvhHF+wctCqIslwZffH1ohvb2ZFZzxpnwQRd8YQAOkUOVhYgMy
AQGQWUOIdAxLsX++eyxid8Ogvuuq9zxj4ysd6bG2cWY9P08QnqRMM3Jjoqjr7Lnv
ER3PurW6XSB8s7MdBwa73dVAIeVKeeNFUzVRUgMplkvGnN1rTKvg7MfWURIcBHor
QbMGA+UHQXMAi41/cW/2F/FG9xihy2cBsYz4C78LqyjV4kGR3CrHPE0lOM/JCU33
z/5+1jEmYjxA2Y/pc+S6Jm+7JhPOJcQQpJqzoxwoXvB0Ktdpgyb0iY+W9cQnOs2u
Ppuw8pP2us4Sk3cz2qVcaXralvKZYo329jzqTXp64KXQRFXV6LVxxr8Zwy4aYZU3
7hn3a7qPU/WGyQxMsnKTl4qd857bIvItwP2SeYZ+4KfTyj1Jg2nWhsmxTUW9MBSX
/cb0QU9NjzepwgymCjpkeuYy4Bd0WhtCnktl88Rj9qjos2WfYuJGSNfE94ObcZNt
e93NgiaWQfkYJxoFqvn+yFJHe95pta/ZA7gNZgiuBsI0OSFAkj5kX3OaUbCwmUeD
JhjAR6aFSu+lhsUjM3JZJ9Zh43oKWq9QA8LuS6KWK+udQYg3U6nkSJ5YotDEpyY3
A2ZuWHxGSl5L1tgTa8PUz10yntcl0ZSV9rcbcd72cnXz11F8XduRIcOBDeGRdL5r
tJFCgLjoyvJCN8blynKYEnarUFBR/vFQtZZ5h3ViBXcTqhtTRZjNVfWzvHIUOIoJ
A8XYUEvl+yGBeYmxREmsT8vj333sEyUiS9sMN5aTv7lxw0RZB25Rjp5aPJL2WYBq
AFCb5aserBzXWu6agVah/CNgO6IDw+czYC2mxCCUaJE7OXjHNz/Urp2kTH+p8D+j
ML785d08vpV/quCAx+KW4G3k9ZTdQx10dpKfbEEgBWH4pJPgqiga09Bu/PgFh59p
rWkUyOYZY25K1Gp+mZPHZF3InCgWa3mLgMZL8UiIqj5X/EDdQEkFLfA/dcYPP2wC
CC80c8r08TozpZAji60fCqY29an8fWKXet2Vz2B/nTZIi88d0Jj7DAi6IPFGM2in
jV2gfsHV3GzCAMV+Qx1/xlLr2SPo/AYwWYaRCtlrFBl+SqjMvkCQFFCnlm0maJ2D
836WefGW8Y9jcYImLdcrRMBRUZhHv71A7JXfWUoBMHkxzDDEKi//V5SAGAcL8yYz
b4th4ufMbTom2twCHbOkI8ZqThush7XSbIz6prXwuX19pxGy63hI99Mvs75z0rR/
eZQUs9O5dW8y1iYQB6jSHfRt8FWuHNRTBTOB5NEQqyGJp0SctF28NiwPSJxMTykC
E/W5aSYStuG7JMQSc73Zwnp7pK1Ca4SqpoLOqf8DJ33iPnrw3amrU33/L4Bd+7Vu
jDZVTe6plUcMZeiRBVCzBvm7fTVkMt8bh+YvG2c8kFBYgl/f0t/OrDXZNC0uuKSo
wQJIbKZWkHi+9LI0gnjYuSKQdHcTXOU/IR7KKf1g3wEQ0cwDreV62TrEvBMRQFo3
++haVTdmdYsmX6C+xM4XcId4VCE66lcqqD9MIRwkBxwQZKz0rvTYpuPyT8ggMvJh
suLiEpICmjpsJ01RYCS456ry/60YBrcZQ1kP5M4XPWImDqWAg3boQ1uVnPRAWihY
ZIL4YypeAjbVPXLjNoGY0ztluAx+8sUVuTLrf6GWAZA4C25Ua3KMBetyV41XW+q9
6b5cqIr8AmNNFK6WDLuMxDW9BBJPcLCz3/NIHxNZUhX4+4Mv1ytQYGuYIbLc8B73
bFW7kVq7LqMwCZL+Vwi4+Y/abHqE6jXYtvlcVDREkpXz1C9z38Gjdg/M03hVMj0/
IFiuyD2SpQ6WpI5IsReHcrzCUTiJ5mSSACY3tObTIsvAijoL+caGSLTxPuc7UgSV
Q+J1Q3MJvbxuxDK7XidiO7LktwEr4b5tzhifEcBDX3Lw3tvdgrH/kdw9KTUJ+RJz
3sY7l17gJZtHFdjUNndx+gvS69WzMJC+Lc6TgIMTrmGzmKWaEcTJht3/caVlQHpA
vQQ4hEkwwGewTy5ahwxyXo7YWOR7JdiLuaWMndUwn/3M5i4VL1uOVitzzC5GT786
Jm/fLRpz/EIiEC49oZltnC+lU9xabOSFq2ow77Kgz3IzxgRZ3txv1/GT7FE4aAU7
/wCmbv4c6N9peKQhk/pax6eila7iNHkqmSLpbDjimBtClXdFlDudMKgVvI6Wji3Z
loBKRs+LKK9WwQ2wz+4yO5TuSQkt5S4yLXBrxXOZl/5/NDAmhDUUgngojyGSQPt1
lWD2+MO4psJfvnKsrcp48RqnhR4Jndg1UYfbLvOmg7cK9FttDmsd29CTx3oKWZlg
NhkXVOt+iTZh/UokOCqL6dDd7tp3iTzDZL/Zqo8cR5m24/T6sct9bs0/kpAXwDk2
Jf80TH0nNVvCRh/aXL8RJ9leMBPanc5gWKEccPS6Iqn7mP62Th4VBn18kdqGscRR
ZETSVHO5Fm3YnTFrwha+ixDczSrMiMe5bX0TgBAZ1/jzj0BSjL29Z7aJn7ILzToW
wan88AzHWvnXqYvziEJn8kmOX52KaadzN02t8qfzh6QrkXJknEk0cxns2dnFY7Tc
gyUpvlGEFDGK++EWXt7GSIfGRek7aHaKHZDT6nxwEldtMg+vQSK+MJWVWxbZ9TLa
sApvcUUNwqkElb/QTKS0dELhU6k4qL0EMJd3UTIJ4iIBr1pJxWTvBjiniDoIUbsk
lFmVXyejZno7ohxi3nLsE85vLbMr4CSSfI/4LCzD4U6Db6j/APN9PQQlulR00c/e
usOA0L0knNSBBiaoow7ixbdXJDaWzPlCrWmcutK/eL89HRWUtUxl9oe8z39vw1CC
YTqc76AfNzgQkDR06gNp8OskgwGiqKujuDqcjaXYJw9oogMJwnJFDbR0yOh8J9Gd
vQk7ghWKL9EyuFccKgA/iAaymRxSXnCNMRtUhP8Da2U2vP+EOXAsQgAczFucYdZ4
MYwpbBvIX+nRUHnT4eoOprQ2HEYTsQBddfet6ngXGHFTLqKEE97p4QB80bGGkaD0
RcMU7vTb5yKQFEyJXCdXk+uq/3NZ/JKzHyIgtciC2wu9g3JrpWr+EVbahLrkYJiB
QMQpvl8Qb1MXSGYxLuY7vbJNKT3uVX9oz+INmaSeOUlvApNECr27btk6RZmB0x+L
j89B3KZDqaqod5xvLCyGEwDKVuiyQezxSX1PdpyBi4a97bEfU0fyY1SsaQE3o6c5
U2OzT36HvRcfX8RuJoDwp2GzWOdcDNKFjdunQmhUWzVaXZ2XBHN/guS6DcvgU0oL
fxDA5+I49pVCTt2EEzQ9DH9AwNC7ZuOkFYB0GNbjClzx8TuAMWYpMioiTz4gs9Ou
3FR/tD+rEOTuCk5Q9Scp7G9R+pfLlVsfscobIMU3X9lR2SgoNbReOgRhoLjYdOnh
tjvviE96pA5T6rO6p5LlGVFfv9/J0KgH5ve+w+cFVWnOFZ48AS7BgvBQ465FktfL
xDhDyGJvQPumN2x6MQ+S5phq+HYt9MylUHu8R46f5m5KQOKgEqghZeeMtElZ7ncP
TTobKxPN0CgXctC/QghfROEm2unxYjBlYVB75BvTWEAf29HeSCCi0Zyww4qU5ROi
RFdG/hufnG09ttRJlH/5vYATisR2Ud69LfJkiTWcpxNIeUYb0IsLVe04Igpm4XMk
lk7DoGoL87DAr0pPfQLBWH5MBMZLezOU//cmeikJvmNrF69q8x7y9zgvnDgGF2bV
GRIUUkVYoANDp/9HhyQrd/PL8BJE+nCGP/bV9Wqnf3CBNHJfSceOfddQGEKWSbGt
iHdgTpHG76fWromp77sGByoHPz9tzwDnIysfs9VNliBX52vF1E+vEiund8UJnNN+
fZYdTBz6S3eZ76ZCyLwroUpKZeHILkah/W2WtbXA8CTRV+C8yFbyGXlyvHgmNYev
9xKOEjsyoCS0zKBjbec/QNxW0Yr26wUTI0MRDm6lFqgMxzonXz7mADhK+EyLOxSo
PWrkbH5jbEpLf80gnDYqs2my8VQr6UbuVzFNIJX9w8vfM7532Py1W2hfEuC5F0jy
v7jDfxt/Ium6rIAVhQaylEjZeU5ApWoWbep36IzwDKnPCq2/7u2gmUh0T5xcI0rx
1ZTaEqatBEsstJRxoctkEHEZyGZfQkIzwMt2SUC0J/Z6qd/liW2yozD/ss6Cq3Tl
zxNYxtY5ohjGkDNqZQpREiZWk/y+QdeUpe5ibuR+iSrUU4bo1hmveBnRZYzOjkrU
04hbB89hARLMyqwHAh8yhhNmlg3jK3PQ/32Zx+0MreYcW0sFwJQwTHwCjUlrl3zJ
IEpHsZEKFL8K3PTOrzv46jXRVVxxQO6jmi6trOLrwmrFe8p5bYWUSmTyedzpAQQR
o0NeJpKCak7pdtJqVPHPf2zWOYhAQpygQ7INITieHlcjudHvN1jc7SL6nlVnE6JC
rU0x2wY276rmZevX803MzrJtkrvRn/znFl5UvHiJEAXGxjf+1omiREF3MBcGpojA
lGZB824aadgP07sanPuc4IIzbVW6wzUlKXx9FLVHpCTA9s1kyeuA0f770phQVHSF
QpFiZesKgeVT/EqTt3ngRe6gQT2Zy1fqsax9ioUVEDcusLfmH3iI42mWBG6o66ee
PPszENyg27ZqPE5yBm1EXFpthoblHV1Z1Bc998RafflB2I+XwvnQNktU5cdaSDuB
b8OByPCGfLlmOwvHzvHff+WqLdkTO3Zg2GyZNzTrdHa8ZM5act9z4iO14s9Ea9ka
ZvE926nku9kRBD6syq5hRzqL0N66nkSiAuP16Ucmmxbzt6DIfStOP4sUUwAVPVKR
9lIjzBZfZVzB7M0k+x93c2lIFy9GCWq6c4t7RWDDKFXa8oa6duxX9pgxBcKOF1TZ
413K52hqqgxVKnNZpUcHGNZoRNzlk7gP1ClCHxMms8B3+SDZBSGbiFm9TzWHV5MO
j+ONWGcxAT+JsnAHd3YDiJmEkUhmjOtgkBT0Mb/iDxBqalAxe/43H2luHDUeUpEl
AtxLvO4rFFdrKPNQZeS5KwZS0QqQ1hNmbwCMKkBTLxEEr+iJEjqHzr5n5vQvxfUB
s7/7VdGs/vZPzHnvD45fEcOiw4ay0tz9CkhHfNAPa3RZyS3xzm3hVaXDSEonTqJJ
RiFnUl4wH7yoGFSWOO7NuwBSppCxPDOjkz8cQsNvzfs4V3j2Ifn03sgYJEerGPAj
+w1hGlZ8Z2LpFmvu4+uu28hNloqU0wd/pbvv4w49lLX/x08v4e+n1Bm7Qd9j3e9N
V+8pLxtK1pFcMxusyWdT+j6NMKTGUyKy4b2EEF7LwBZuhkn/V7v6gnbKwu0Synbt
Q1NJ/5XlE0Tl5eCm36IdeacWGKpyT47H9tQMENRvZ9Cm0Y0uYIKornHQ8UcFyG6R
x1Xc6G3YBd3e+f8UdmLNSDIwJVIVWePcMT69xrPfqiS0Wv4KxmbDN+dOy6EYuQHF
p7Z6m7MGMWgySNKhlXAgNmsgzPb7CmaZZ9PCnlQEkZaKSQiwhWgjb5l+EVv/g8m3
2cmOTm22uccBgESHsXGPysYtA2dtiKCJEdo7nc3Z7SgcgpVP/8hs5GJmHci89hgg
0Cav/AtIQ+ct5JHhkh5NpR1r04Vt4Qz1YAxwqyN5r+3yQQt7YeHoZzfr+MB+QIzp
zfI1HzsE/8sXH09e5YnD1fPV08BH2Bnm6KwYc2cBPKvLOfNiprxUyzlUGxWMiS9H
+eGMlOTbPms9yPJheOY3HDSm3DsD2EqNsxObT2GSgECQIfvQZX2W8KSaMRQT7/Rv
bsBQvp78dI4K1VHVygsQWWC5q30hXL/METTrS8GxjI4=
`pragma protect end_protected
