// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
G9eKO9qfdB2l2FkVHec/pbQBYuBiCp7VeJlLY1fv6kD/Iz3Dwfz9e6FgWxsxnZs+
GuNmyCAXnhgvro6p4t9/IT8mPhHTXsZ+AIVP6y9PjhYWAkRraw1Crf5lcKzfbsck
RGpQlsXOBAiZp9/T3TT3S3HT/gEODBUubAnycAyfS/U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6128)
Jk28VwXAK8OoypodyO3pn5e9CnZgyu6OP1pOxJrd9H5vBbQf1u9yKN9WR0PNzj59
J0WJQ8utOd7BgrRtoUvuj9O3OriFNb3j7L2Llna6vFMCDuoQ0OlMLLLIPiMVspVi
qZpSGmIDBkLgVsnD7s4Bc0XQB3L4j8DvD1WAzwUN4wAJCr2IhYJ1oIkI6hau4uYM
akLdPy1FYhxQ+cL5PMD2lBj/q9bfvHo4uco0uxUKKRPO+QYEIs5prbTmSG3/RBSN
ij/c0+NGTzOHGRGL6JeuYTbgiNybrmbxROlLiSTa6r5S+EAsQsnXbqoUA939cxVi
gNspb5Hm5m8SIALJ6La6aEBtWIuMuyIJX5A8sg9eicVdB0HKUMst+oTXQec7EHRh
cOLZZEnuPKHMEWAyy5yZB70DR3HJnNf9TMUAHDXbjnt0L/PyodRwidyHtO8vlVkT
dQHF19zqxQ89vaaAgg7ypqxlMANz7maFtHQhIqV1yZXMO/1a6SfDk5fYo5RFd4IO
nxP9AQYl3Jm+Eb40EJWzhNSf4GFIeFadOyODIOw12E84WpJdEFQBblJGaPoBBCCm
dJTGndV0B/78njWbBg59JuLkIo51R16Zbwgz9HRAgtRGpREbbHDSSjOKGTFAdszC
sJB2UYj9RDApCUm50kNK0Ot8iUIpsf2ovb34He/+yNrJGqqg454z8ZSOgF91a6mj
GV8mGD2g4QFJ6B4tfMwJDQqZg3E2nhLasjCnejdv1Wi2S7x7G9Zu1p9SQkQQv27G
Ts9VTJAORekwjlNUIZpEZjnWSf/fgsDtu5BlYWNqRXtKRdWqZ7vOUPkmVK3pr/xZ
mPhwD8rYmQL+PKi6+5z7wX5Gqzljb13otwLpLH1ud2AsXf0KbqpJNINOPGcGGMAS
vqJL5x2B1evAtkWnH2hgxgCZHEkOBffjOE4r6uHXl0wGvwLUxGfAgknoOy9vm2fa
vhqyRgLQM8qXPgSUUPMyBz/6gEBMALd39e2ZS2ikuLQO6LdEEFkpPlTa+qjEQXQg
D1pzMfpxTLrgrYRTfaPp4L+NsFdMe5r69P6nvdSQ7fQnWRaftTIuL9bw2o4DyixZ
L+Dkn0EgnD3CFrQqeV+zOmibWSFZfLN/JPJM3BQjTJG03oM63xo8DdlJD0O8V4b+
q+Q2mJmMLrR7jrRlSMfR4HBTn98vN+fUkylgjrofHdHurLzYpbv6tP6BZgsMxhJo
VcMmOgpwyvDIczgmmm+vlqTEq3DrxC9dEXP7Qb8TSwN7OQGVjmXB6DIKIFuigZ0w
AZsVLCQmOshQ7sx+Jl7UeY+BT2Qv832kqzk9LrFNZOoaKQ4aiUJL7ABXfI1KWTYJ
DsyYsbp5bPjsZteQ6WxhtXRylb7kj6Iof2Wqc5exCoEqDVsuvg2Upd+iWqUojPvs
PYIpDNdjtPWizjh/R6y8CVtTvYnzA+x5rKMPP3nSkkto/VK08ib7cN2nBI3/jAmW
zGnqUdJMly/338OAYbnJVHGX+VRX+1acmqIeC7KB4Q7nsQb1r+NrlDzStivwmwOQ
B7YDU6fpOMJhRcYj/Tb2emQGI5/798ggKn0uChFhCYYbtNqDKBxKjZCzgQR8cn1D
7ZDmb/GdzijtyeYy8aTzT8LqB8KHaI7zYD6zejeST6qYMBqhMVJPjvDSet0Gc6lV
zU85N9+LzK2wKaWo0uEMtsYIs0yfR9u6vLuaxWPxASh3jVbNeMLcShhAQuqNr9Ri
DaR8ONhr+daDZjljBhGZdyzHquGPVnBUAaGRJrtbYo93Xvy/gLH1v4T9Y36FrJXl
UnaI7/km/n4MEa9F3ou+l+pKhPnnAKaVHmA7ZXfNkbPCDsrITV0e+zsaHBY2Pb/T
Oy+gdB7avIIxM9scWxvNuIaiB2Xd5ZxJl7Ig4Hx8TrNcgEO3QHxTpQZDWsqdawUL
baoUTkoNZjvSSl8oeolmIQ2/lz4E4N1XOe7RQJDHIY59Ak/1d9/BH3PxcVQwpf5M
igtmZmphK9O7xnbiIdsMxgTTo4/ak9glEh/q3hcHfxX+5HtzgHPR8yZLxskrjTQ4
L08IkRJnG6pjScEljgJ9wktcRFrni92Pg7Dui8D2luTDZlYx2pWGlvJ0lKRmuFCF
PPuW3hmnKLv4hTbHs6KaeRFffr8FT+PuJtoUb3c+joo0vYNVdBuCOo7+fcFc7ump
NPWEQopCyxz0d+xH5BhnuN/C9JiVyZebJX8iR4tabBlEPT3JzVl6pRb65UOW9plb
/2knV0QD3eYe/5ryV54kiGfEP2YakapWXbACHHnbUjDLoqRbyvGZyBEtgUMEtkxZ
7Q5eJfq91knJXG4aRitqFofbWWV3mE9bYt2pprN6GpGPzamZFRmBCWAjA/cejs4v
luVOYGMMqPFOYLljXKBOnXVhc4HWwi4XCmVWvu+mHW02m7Fe6t9CUsg578TimATq
p3pHQ78nT/uz0jZh0crJXfaT5je8Y3Fns1Dw4KMmBmEg1aZvyh+MQ+uc9u7qxu71
MLj3ebRJo6xouS0coWnqEZC+tceG9mFuVWWOhuuD2m8wOfaNjC0SHBSyVAs+e8DX
I3MdwFhkQGKLyvBlSfdNjjdpIp7Rl4E7SvkuZ0S++EbO0mE4agtftE7bEkRaH5RE
f/oXb2yBpcwLGH+VgsS7KYTRsgb+QTdhs/DNGy09pAvbMIqO5jB4UbVcTA6gk832
DVAAWC+dx3gh2rLLseUKZxv3nccHyKmVmPmGPXeQiXdx4DnaUHICCZcJDtjg1jlm
/3F9dDszkvgEntqQ7HEQavPAJ0YeJMFltAIcDJj6AF8NbqRMgNNl9XVR9BrB2hjG
VclqO/rD06vhAdjKE5fgdgVxHRB0kiTSZI0q393Bh7Kwx97qH9gno+TtvkBPUGfc
3uAIWCsb75j0cH5EnT/T+1UWr1VlwoBFA9KLnZFz9KvS6R8rqqHrdsc64upztFek
k430c+ya9o/6LwcuM2j+4yN8TOEwTskjm8S2fax1BZL5gYuaIIuctBznpgGsMciM
SVgYCMRvY9WcX0HG1Ra6CI3Ioz2M0bZrTTMllhK5r3nvKfTKYa1yFDfSTyhw7Epm
OJUpHGf5QgRCSo5KlC8otAAExJp65IVHJXtRh74Vn9FVFaWlLy/9+wgp2LJfb6YW
BJ8UZhoB/j/OWQ+y42doM0xxAdUbxazHKCw6ba6Bwr86HWslQ7pAKKOiMzEzE3+m
0Ci8tP/hesbzAFR5+SDDSA38Cnki6liPGFSx8aczH1rMaego9oqicmWTd5NXyeT9
DNp0kb3DszXMYxtTCK8so5FsYVxCWpQnUmmEzyMTQ7L8J/3Bw6DjXgcm6ujOhyby
TayZQlivlA9jZBQj/WCltnpcNUoiJmNkSzKPnyZ/GWYOKFCG3suJ4TG6cWAm0Bcd
oreUj6suvM5tNKiplPVGcGA669PtaUCO/w7HScsOG9THBRxU8B/UfOrlmQaS0o5T
YzO4vPAjJvu2AAGBRb2xiCUlSzrnNFzITJsjgSuR/MBsoKykQ3MAErIq6CJx38x1
kBJFU4DmpVj2c5ccDTCdq5nDIobPDL2BmKO6c3rZ72kwTEwb5ntaHwJ9r1RCIF39
LlxKTL+dUaZZLEbDHdZO3BSbNKwRnQPsLZuxQIujsqV632DCTlzWB6dDvenmXfBA
z9RkzYJseN/ihvNhjzgy2+e1Gjqbb9V2hBC+C344KAKnh6HJweefC9FBPnST6BUV
FRapccRn74Qhjq2Mz2hSqjZB4ukHoxK+Sf3B8/dzcOL+hyzwJ1pyJqi5qJ7anYvH
Tv87z3k+hFCBGBCVChIDC2g/bMT0EBEEZDYufcYvcJq+6FSTiQeyz9mSvK6ChEp2
xXHKTGG2FkAhPBo+5JKsx7TYcRJQ9R1I07e8qzHJV/DoNS8ZgpyWZ9Y9qiccIaWH
z3TuZDY7BYkM3/i2pcuVfm3wFf8bcyr8d43XYHNVrseMYo38tuMZTW7gGuJNF6+s
wC1PE/g1x7QxP8i1PzHtvno3jyyz/AtpovTFsyC/9sbdu8xMIQqau883lM3QBpwG
j5cP4M2RZehpma1wtBQ4woMDt/tSn1xCH4L/me/mYH2faTV5Day0HXi95ounjftP
F6KZcmxvejKCt+eVvLQeS9JnU9XLIF/lN/At/XphPr/06CJvvl57g9zeo9AzBc3Y
IQUic/6Grz6jHaD39xYPf//MBWZF/aQrEK/tRenWZLbKkFc8vmSdWrs76yYOlePc
ela44w5AVmj+H4c8mFjexxUihqYuvjfhCE5qrpgC7Q0W5VeUf+7Oilkzl2WLNN2V
EeLTljptdi7FKGFqfpROa60InkI9xSbHw4FiqrUZVPnJfuIPw9IREtjFYrQGtoy9
f3yx7pZakn4V1AWmVj3AbuPQn0nZ6XuLuXqQMz6YunSUl/NzkjB+bFEf+dfT2SZo
lSWjGIC30zjYMIJwL+H4PHgQPHEWGMBDAGbc4BWomHw8TW1b1L405/DJ4Hl5syDj
Unpt7iuBTPAtELPmx9uoZNIcpTrOVJXqH77DL8zJzw54p6uvi0GO5tbs/nabJ7Xj
xUuTiOJBeDlpS+0LMOGOJysuyeH2FY0NKhpkZlOLs+QagZktD43B4JzOHzcTIdsB
/SAI/3vtHRqHK185XmYyNA6ugGIWqwGqbiSXUXgqt2yDwJgfFw2TLMwCe2Qvlbi/
Z+GozacyjC0ObqO30TQGCjVbJmUaWS2wrhL3KVelx5OMGlWXt4d1soRkLyBnZl68
a13/QylOA6jLq/TRONrwP8bwpXMdQ47IBp7F/XrEzh2JByvnQ/Lcp1v06nVvuL2q
DfDGY6JAR80r3b9eyzfJReOyO3yAIs3nbafhh1d1ywR2bP82c+uyk+x9rWXclEhg
uZi/SbBWk6YGLOFQazGdcGy0+01EJIZlt68nUKs3niPxQYgAovhIu8bPQ6glxu+V
lJ/pyB0N/aP2NMuaUy8tsIM4AI8s2siIYqgvX2udqM9jMBARn6ulE4UHIlQhHZae
TJ15VTW1fTE4I2Sr/A3pQhCneYUWZ2mZUCh7XW4HFW9F6XZRZ4ARPep3KS6ajdnd
a/k8cBXUkwmRHR1WdsmEmu/3fDkQyFb2hKhpSYUT3FVvD55fapzdsnK1jGRK3G2y
DPiiFV3yFrDfIlK4ylnUDxTIIULfKkfpb9JJtmGI2eQYQeNdoutdiR4MUKZWvVLs
rQfFYQBJYugIsj1YZkgOnVjxNEut8vM8SZSptH30YI7bDKryOv/yzQ7mh5XyjMxX
GGjhjXUYW/aOYjM24a9LdxYez00fZUAk9BMnEeYKJA08USVXUnO9DsBLDbJF1c7r
4dDKdjfxDhGojoD1Q4DAqY9GFUmwd4AqbPVf4JttOEHg4RVCPZoiLpO4kCZyUeBX
uBqKJn2gFEqkJplM9xXOmjWDXZ2eEbKAcLEIjASZG3gqKNMg/A6FOUSCdiICbKTK
O60jrLQkLwZ1lBGL6disjB60O7X34GzR2FT8H4ANlKtW7UToS6S9Kv4VlAtQ9iym
JwI+t89IcwscMk+af5ipy4cORw5w+Ampyt1OCeqQf7OQ716HjF3yu+YwwYtHeXas
9XJtOBMfpDQtINAEVrp9mmKUC7RPqE5i6aPQt/WmDHb4MLeB4utUaaPbtBxtCRlh
TgxadZ/mLV26tEitC/9TK3drvfLFCVlwukFeyVuIOXotN+wy+3UxsS3trXQ3PVCc
klOuE14xIQLFb7TnW9knwswmo09ijlUxlBB/uPcE909eLB2wveh85lkUzNEu0/Qx
J4dl9rXWzXNUyXVYinN3ldrXbzMQ77kNaBZA4nY3I4x++Kkhj3rmVKAGrLIjvb6D
DX3VkHvrIrZWF84l6anbVqj3xgUanR5qYDDOEg8bJ0O3Pm9OHdzXQ8IgQYejLSGz
1grajnE99U18kR2FMsW9q/Tj9uGRuuroXZbyB46PLbhv5T07DB4174r7ujV41MWg
8R9lBf8kpHZ7aWdOPvoGGLT848mV2Bt7r/1Fsx9nq0TYFOcBztqN4l4p3Zndosxt
KAx+2dHijJJ1FVtm3CkSyU9Mj0eFcTCfIgKRSBhD/+sQ2vLZSYTmomqDeZb7ZefC
M8tJwjzQJa931XwTWZC/e5hiCgV7qPdmSCQnemfZ8ZR5Hkzw8i6enCmNI4WiqjcL
RtKiNHJDzxA7EvicXdZysInRp/otuPhugjNhXhmHxiJiRRA9g9JhHrZpw2SeY413
IAzvlbTYtw1CcHLkI6j2ixK/cQqmc+OUJehG1/GDJZvJK0hCjBpbXn+G1GSyilQ6
/o6dfP5ZxjXSAZ5b+x1XDN+p207mC1Cz3dWOLlxpfJ1dy80LFauTbmQ76Godiizv
qU/pM+EYx/vrrxRYat7rAScfBLsMtEr0KtWOnbPrANCbgkVMMBis5D1z6lVZT/gq
DhOtDhClPkunNFik1aC138hq0YEKT16YA/i8V2caOtvOoD1r3sBSo+c+tBrnWHMy
zaQh7Rk+hKxIqvGMdbhUthaHuMm1FUvxbhzvvqbXacxu/3PfaPRwOsE0kk7Zk/aE
dx1raqbDpUGzPVnAm7bCbpFMK/0/k2mPx4zB8OgKL5Y1KQokJ28xJFd9sI+fO88b
wqkMkdXlOAN7B6KODz+PNwQQMcBTEIfcFMlIWDM/YbAOk6TRQTb4yu9JoJbFBY6N
YkwpboPNFXZLZdXnu/voR59MKnYxA8DMzkM5zpt/AlRHE3zQaZajX5nbHwkYvNWh
3P/m4AAzl2asRhyO188jiiqdYkoLA1mnFDwNPqvNInHL2AbalhYvkl9XYDTADzb1
04usKwggR/sKlKQzAZahcnV+g7V6UlSIxILUoXtA09onSasPsiwemzUhMEHH30gy
ashoaQyxQViLQ+HJ88PRhMSV0cI7KXjZZKcsKr4DKy2qite3D46OEp4LLNSycNDg
Bg62O+xhhXA/5v5FCMLRscR7k9A4m7a///4dauCSuRJKblNOAGoSXGoZ2uZSmjEM
XcI857Oi4yih3q/5ZsRkl4Zjn1VICdeRHsr+GbCfyAUMv/ZwMVTwy0t91DSK+5YD
2plVKV1raNoQ/P5OA/jhl+GzKWyrrYC7DKyQAU3WIZBu+oZTv0jbU46DjVizyXn0
Whrj3JOmflGK7yAW7FKb5ErvobmQ1E9uPy3aH/uZ1eV6516hW+T1RXWC2h8ljBx9
JMDz3jiDitmbK9XlwMjJkmny5L7YDz82huHu90xEjnk5cn3pMMgLIEA4wiTINV4d
BpwTmiXVZtHavc+qWlgZffY3Q/n+Z2T6g1QTYRQ6AOhYs3NGkpomGwSAYaL+/kCU
6UII30PL0XmQcKPDDFRQL0GJXGH67ht+kqCH6QVZ0wdFARyet8Mw8a1vr5oaYTTg
vVdXEjpZzUvL5P7UIwzvf6Mbh8tdac83RHkwAxQAUw2zlfF0HYx5QSGz9dIKSXwv
zt5kTiWTBWafdvq9OXgf/GMF8Af1Xa4JUJwPTvcPH5pBHQlE1PGpCdGLaEtqSiqP
W/5snbMh7KEtnSKUEr2YC59bDjLif1nHM33dQl3XLp2qUdZM1Gn4Xp3Wv0mo+gJM
HigJo9bODAV+Y4Tl4D9ukcAiKg41KDdNGU4hsxpwwjGimoe39zXkVUWackhI4mc5
jw5e6oGaMkeI4j9YGKZXqlobU1294tffdFwX35uW6EL0bZU9FoqmayIr9l6o9bSs
Iiyyh4yvLs9nrez7tRvvIEEH2JofnQmp+El66pvk6Vl3cBGJquMfWipzh7kYbHsE
Ma5BKEeKNVDYA9KMHc8FJTN0dDbux3BzYrwSY/p4pKO/BLnlMBsy8kxg2PBduxk5
xZZ6nkzEGgIS5id+3IveUzSqPmmkOMH4Op3K6QfWpd31yfP1D8VdKF81j9hFg0tM
8jdx96KF6K4aSsT8Y9vk9uPazNP9y96m7IVLQtVPh8IBCy1QL2LQX0MHVgHR9BzG
zZraPHcBt97kGaPJb5AxCzQLqjhMdLBxffPZLDoluSlKfdxruzZ9Edk+Nm8FMJBk
HoGgZCqRS5Iyjm0sEXAe1hZxUPXeMpQNdQ/PkQHyWdiJAAFQ/G5GiraBXBANcg8Z
lOMPQROY/Q1l4NHlr2hljFC7jY11cUAf45c6B6hvLDCEYg40rtNYgc5OsDhrqLd0
4Gqo340YXdBsFe7rma6qUyfXQSvtfmrjbqkJ1NsT9eo=
`pragma protect end_protected
