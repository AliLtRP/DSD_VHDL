// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:39 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
j+m68e4JWboxai484eofSJKCCMnEUMpOyGz7SoLeGgrUs/NqLPpY17fmzeQH/5sD
Jk4HQs6Io4nJCCH55245tkwAEurYQr1HucXErrEyr5/GRa0RXJd5TN3qBbxY3EcM
t/6uEU/0HqmNT9Brb6a7gHfDh6ST3rSXvdBQWhT8ypM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 239552)
fKkzq7tmt6iVZXGTRZO9xmNwU40h9ypLjD3VqBYMOuyiXhCtTS75Mq+H+ur1Pitg
q+x6P1A9PLT6kr8mo/EHbfVi0/qhi495w2su92Fc2iFzT4FKywFnpU6a/H7IvinI
MtTTegi6BdeaHG6GZZoAQCCLnmhTzw1HsOPm3Ki/I4K05HNSrLP5Xorn1Bqy6WpN
G2smPryZd8fEjjkNT7ROzx5RvjhmJ5VFF60H9tGrUQKp6ztPx9jfdoaayvl+GWuR
edYlflQtKGfcxvWi9FadIyG5z3qZdWpUgTApc4ZI/HFECvPfH9T9ZneLbrRAnCna
kctNQGJd79PVGv2gfTQUv7NgYsGZyTLMx4cI7TFDtTZwZfPRuiJ5iXxLFasOxvPN
c0/mPGR73wOpZfKu/h74DHsBk1ptY+ZeG7EeXGDigGlC3HmUYIyN5+8rYb8x2FDf
MP6ApQy1mF/lHFJtWfmoCF/Raw9iz/HUchNcohjLYs/zduWm5sLTTEZSmFqNh0LG
JLz05t4lKTmoNYxnwZ5NleWzLzrno7VTrlBVNIzTwSg82rvQf+DP/6e9oQ7Q3q1g
MwdG4W6eaglIcD6992/yMgzVjufvckl+RKCAHhSoBXRKpIKksH8tJbdV2gMUnRd3
TLwNtWn0UqDoqDFP7EO0rr9TFMqLLhJQ7Pmih6OKKrxMAMt3vS7HR/YBgb9vEUpV
CxR2T3+9GTElnHAGnz4QX5GW+oPGBh1n5VDDnS5mqybno6/Vx2OCI07Lld9C1NOw
Su8QBtv/LpD4ddeSlFG5PRXHE1rEpQgoc/4sXj0DAEK6RxjWkp9o7xmgB27LA+sE
WG5lXX6FSqs3zfdYkvb3YxOut7gIkEpun5jHe6Rl3NjGLjncDSwvPKC4SQt4ug87
DqZ3zAzAyh0o9VxBdhGg6TN7gu78+GoHZGClGaHfa7EJ7oIfouuzzAQhR/4RCB2A
ft1LvM1Snbw4ho/rP7GzQZ0ScfWC//3JLp/mhS00d+TD/2t3rA/k8WMHoLNwBQNT
OgqmZgB5QMuJTPe6UFzj64nG366dIlgRAMBPLliyWdNdtKzEYhPH8R2nc1AZWigJ
JpT4tEtu3MwYDps8ZPbPAt/oWKm+8DHrNJjdfvhv0vjQI2arfqR3QEI0uPuLQgGD
OeYyEgI5Bd/J4fPfjARB+pKtL3zvux39BQAIl5pS4HuIBjMQUGNlPeSGBQuA3iUM
kNY38wi5Bg+ANb7BDi2LBh73MrKptFZ/griE1x1kiwFHhhB+EPiTVt/ulPJY0tPE
uT/qOMNWiEPIXFZCcOcdIeMyYx3lEVw2xatBmxfMNWC8lO5jDP7eBMuq/Ayexhlq
z0uNXGGr6Z/1xKwQ5lftBy5K8cbRUgXPW+Clel1LZK9pBp814bXXQY9GpVSpG9KW
wJSbHhve0GsASBREGGYrbKhUxjKm5IAZiYQK+HwYVine5HUJt78DE3U5jamQAs76
uQ3KUxXrxwMlLVDXzm4DVkbbGyWDBlWqJjetuNzlAvHD1GkL/FJI9XYp9V5tiec7
5ZaqGFzdFzmEb3bFpyij+6dwLt/6pyTR/lhHi2wBFdeMc2oBwwJCAI3kxhx+ufJW
b8arc8S7150Gof75nmyB20I6Q4zDSPTALrpQEJUCNzt9chjYU6pkc7+Ox5h2FHbD
GWGxwGRZxAuGm2S+s6XatoP0rGwwoGg9q/dsV7fElPW5lxqeCjGaqU1nyI/mKqYC
bXjYJYVoQWxeQj/v1D22ytZBW7lhq3JLgf7zyz5qpVQE6NvhEyONNWXxRIfFJ1FV
QmgcDMg8pxxzjGa8DayFtKUHXKN2klQPVhYzMqDxT55nXdPw8850VvrVpcTQV7Vc
k/iZW2Og4bjRa013StnTwXyg6shMjUy4aRI0FYqBEblUADypOLnqzmmT+pO0OVBP
VweZ78VsR65zJ47DXq7/Ja7T2h/c9iBAHQ884fZzxMGTlev3VCIsFitVkaNbPUis
wbpYXlghiQQcYEH9si2SNB8SgK6GiNrH2Zixa5cIU85qRcFVlHgaWYXzj6oSKZCN
hkdUmZejIx2J1p4YkSPjibtJM8zy8PpjB7vZ+MshMQ3aPiFtXD62c9O2TflKBs0t
l358HcqBT6GEBOsWVKkIO9KKPY4n5fG9NeuBeeYKLspaflUJWWtv6+BGneJdL45s
jqH8O5YCu9cnnsb2myx+kZ2+kS+zPNBiuNdjNPaI8fSowr9u6i/Oix/q98nwXg//
ctATIfNmFYNpbYv03MUce8b1unJJk9MBQRoH5pmHQL8dYamHc2qOGpRlHXeqnR7p
0CgRLE3/pCYT3OkBXpQ2S8XBM0YKHyM9vYEyrk01E9Kf8tGrd0OpGVcOCA+cqmoK
N8fSYT7NFnfhPC0mNKuv1Not0J0pwpWOeNMS/6e6YPRNy4HtH9TZHqPO8d+ngSO0
MkYezcPlI0r8Y46nNR1pGEnT01sh4J+J25PKZwVNuQxtwyOQ9Cno1E5bQ5nL92EE
a93zk+zx1EQ/JP80XiEBonuScQWSYgTp3WTYnD9JclzzbZX1RNepX/AJf8gZc7QL
qtA6/o9qFtq+SBqFLlAaXTjgxnMPctl2ohGYvhIOp+TBX3bSVXMbRiZwnow2TShA
7FDknkyhoU4A2vxYjwx8/EGN2y8viXqW9kt258Vu3GniNil/etXGb4bHvay8IGZP
0LzYnno0iOxmqoX4cd6gBvbHbJL85ZzxW6HpvoFzhMa8YZRgkR1nopeZHPfBq1yo
QlKovYZaiecFosoICXyTJbT9Lwclo/PQZt2SNEzWTUcZE0wmWr7AaY1roEzcYsaG
4PoL6AsA+zqfEz/jLx620wiXYQIJpdZkcZwW4DEHGy/cC4U9Hal8esmtKcP0AIhY
KAA9kj+hn3hZdAa2qRGkJTishRbycR08xKRI1bR9EGo/EnOu06AG78s3XhxJ5sdr
/5pXshGOl6UoA53dM/jED/VfJQmZnEGRej6fAQL+P9tuQ5JbE9dqPIYn8+gHREhH
GqbE3Oq5qmm5krmkNJNeWJyBouDd/PSqYHYiGsbcQfHJgNIcyCDtZCUMehy79UdB
MVsIdtoalsd3QmDF1gFEi5DUzU9vPMgsAgaCRDPDR6RF5ywR06XRE7LkzjxTZGCi
dzLVerzrTnvTatVBUBZSpeoMA69u1k0CCfXv2FTPMKWSaV5YiI2J8Pe5gQe8LjLo
CSpZnvoZRv9S2eoWZvsgyGDoow8zmjieuXcdbBGNWXOsUVqvIq/WEKbL0ONPH2jZ
Pmi65lD2ErPWaSDiJohAKAOw/6vAC7zlqIoeUdAn9W2ZB8zPyqm78bV+6sPB+NLi
PhODshDcSBY+hcfATKTSLDYptNqAyrhE3Ct1bMvjE1TV3dJagygt1thFgdxVoDk5
Eqp/176dj4WEmOus/iUiLVn5N57NnKonvDMFDMOlelB6aY98gL1kIl0EA/uDrJB4
7xjoxshGK5jNIyChVOnhVw2lUvK/j3Nn+ifg0DraSXNZ1J5tl4zR7B9OLYA6KMut
60Dvu9u4MM3AWRP82oCJuM0Ez5MkQ8sWeIvv8k6VnSAwZxawECD0tm/ayWXE2W/1
5yAB1dLIE/zvGHB2MhKMX4KK2wYJV5w2BSRo1D9S6zVTj9Ds7EO3CYHxb7MKKtk8
FYn5fGtZLvB/0EGyAr8L7rPAN3p3OWNN893rtXNuSymFsjIcszRp8ppKHqdQsxuV
64v62Q/MsXMk9AP1gjNWga+nBb3xDRAB+MEk9+6a8HeaXBbuHQN62Ssqo2o6mTpm
b/3e3YkvuLB1PTpx3BTG41lnC4nP6cjxpdvWL6rfj8xYZriWw9BNDhJrbzUMK4/U
12TPZDSON+uQ+nWZriiJElBWUvzsfHOEJr1tlxj3n7mUk8c4Bc+jz3gLhcpF5wHs
92KjCUC38tr9WIiiibXRRPRqXFVUpiPDm6QDUjfUqCvXOLEHVQcOf/dk7wf1Uc6i
6qry3farAi7kQU4AHcmvsUUqRx+UABAt8rxGcRZy5PTjniIVKlthSX/CurRwV049
Pw6ReYnX3gJMFrYWe98Uz2jENxjGXLOtiRJjV7FIk9wWN1w39Qwb1FlYxy/ChcKf
ynjweqUsYv2ArjuiaQCijFeC14B2KkTmU4td/2czQ4ERdY614lmFbW9tePFPSlxW
Ob9r2s2Pmxa3yQm7aCV+TQo1Da+wtrCNNCL4xz6sGUtOhPH9/jblMsmpG7GBf7Ux
Vu6mOjxoYYvj1v/OKYmFKMRUjNetc8kkF509V4nka7/ahG5sDIc7g1zHNXeltk+E
fGlPrww5UKj8hP7C5RZ8YMVVM7bdP9imnkO3WBLjc/umZSYwvEuSr9hWXPKH1M5T
7F5OR1ahgDXfT+CQW2QwRfvvOtHjBtbwlCw9Sk8Cti9WDmWdw/q3d/cB/vVxIuJu
OOmzyfJZL1YmRoTHX5yevxZu2uucUfWlEHcVsYbxZPcSX4tim0SXdsTE13b5oPyl
V3EAslvsCiJohsg/ZGOzixEw/l6pHCRXmF3GLkWq3CMe1QSXDPvMdYyzJ7Zmjaa4
pvZzWaWW/FCOhPGrjWaT3QjVQrMsUu5is59nMq9ukmR5BoUf3iGDyyBKN4aN59y6
tSeILsX3I7c5f55//jsSl1q5UfNzj/gO5ZV9aRhOtqwuU8PikFtnOXTU6FE1FD4r
tG9EyekW0RQT+6MpXbTi3y32qjaI7CXuyPAgw50RsV+yc5CCo4/WUaJEdu+UE820
3597EMDInQD0eEA4yKqgfThLSRg+In285KOEoz3lSx+5Av7U8T+UmG+mQCGqnTPH
toOSzlosiVWXHM+JZYJiOYJ8qRHNZdBJzOoFIge36YT45X4HjgrFGqNlgr/ql673
ADNfcyv9p02Ub9LEYJb3KLH7lztEEkgGIea3M53iLqiReUSLV+IoLenIIgiuizh6
eYH0HR9YeTk53ZVuUY78q/wdep9gkrqD5u9XTA2kFYv4QttHkNbcUz8b3qVLoG3+
R+LPGl3qsWcYtKIjaWAoEfF3HFbd6MRMY37wWmIpT9uxYYbTI+BhkMAMJCz/J5Q4
+ozeyMB6N5AkmBxxL03lH5vxSXbLlvQlzueSKipkpwuiPFuqNF6A1dmbjAT7TIOT
z093zAQ3YKeR66e31/33GMSiS0dRZQbx0LiKJf4zEUR4F94auljAlHKFPv4apB9l
FgGnIB8A2KqV/fTOmCshFS5jYZxMGGir3dC9Yw9grcl9zDwy7XEou09Y+tfD1OYQ
B1JSNE3mep5pkRT8v9bSefg9e0jLP8iYyAeAB02UxkTosPl99Y6683rl6Y8KclGJ
1Yn3noZhyErhm1zlPznX1MQISjeVLgQAj7Wrs5MO0Aub9QuYam3jGhxcsdQMKfCc
FErLPxGcGogLyRFrLiDX76bRbKC+YFvEUWfxSCzvElRB/hBLU7OWfGpOKjVXWFaK
F3/aAZSsWKt/uhr+M6DEQzqWUA+kdFZX7wMoOvSFUCe1xlo5nwo1ORuc5OflGtE0
d89/YDeidJEIyEwurfOzbu2kMjD/vVvr5ED8hRM5phk1iIOxIChHhj3uU7NUDnul
Q0TmYG6lc31fFOlKSxlpU50tBjOK3vOcFaJm2mzMhulbdSHeHXPCt3Wt0ceYnjB5
hzCiXGqtbTNdGvZa6kDib94GfbVItk/tIZ0k18k1Nu+pnGXsGb1iFdvJzgPcc9Sy
GlMXzfT/bDWI01GHcy5fPY6Eknk4iqzPvcF7Uw+GKMXXShKDUzkF/LSW/BGdtx2M
w4WwrL62UHI8oO6y3wD+tr1HO4eVQwdDEBDBmD6ReN8BcTOXJe3V3Dqc6lyJCYtL
hw500F5jRqM2AXCTCNpbenFixSgmlA9xXntYqXzPy9fVIP7nmqc/plVEdHDoYocZ
DH6rYpjMwI1tiE+cc9g/LgGxCVAhT03VR13GC1jra9ZEdeCxnlwueytCuP4XsgCa
GkLlBPMUnty/veS531g9sTV3UeCTrHnSJKWizvLYWkjU21BRZaK5Kr/riopK09Pr
yd1Ps8q/S3dSyT+SwlTJkot49fZ3zcJKYwVfG8i/IWSNfhhj1Gds7tlgoktMexQd
oa6DZ3do6JJcwg7cxTi506n+4pmZ3BLy+DeFS/h9hSm2gs8IHJI3ShMEaTnGeGyr
NtRyhK/G4XDl+NUqIbPEYI5SZhJkNj5EDnnBFEJbt/CeNk7tVKagu0+tsNxDbCRH
EIjuvgl8A7uVYzjld2vdT8+fadRP0HPWXg/jCwVBwnaYedwwpAnpyJMbaKwvcGAs
4GiAub4x1SkVC30jb0pX4gow9Sr6c0znuIKl0cWn/2c8bx2RQ1qwUEe1a8V519qk
hxr8EBEfE9UkEPxTvE3itL5LJIlPzCO7CbQz4kZ6UenPr1SyKk+skEaaDtQwyM7W
0XKg27BLa/52rNlIQr0GrrhYtCEF7xY6ukxB2Qso4hwENx0XSNya8kVdZkV1UCD/
dw9Mi/SdmqQAPbWYkzpSUABMLQ6lJjFLAfYghtqnayNRGHfhOiTq0NKNvqwCFUlW
TiSSCxpIrY9dIh150IJxnFwzuN8gM4GosNA6jZsqTCWBA8nPbLoItXg8vOeE2K1g
sqHGllOcXguci4Fssgh1/CcjOcEjCRC5Q66L8a+RqY4ZEfmEU19VpQvRHs5fH0rY
dvvxRnka1Ye+8gyH/jBXyeSAefVfAT/rmn3JodOiq88uoxKdC1Tl8LNiFxCwICBo
kAlkWnGeCeDNZpzfBYXsOT2mQ0TCbembchP6j6cFY4BzcQNBiFFbVrrckX6iqJXW
/0raa0BvGG+dG3dsqTewUF9Ouk3ckbBdZDmvig1ar5OFhOx4D6RaZZ09R1qNeHcS
SofToTkUxsZLlv0BfPnszzJEzV4YXDJbHKBizaRjwH3NASuyYb0pCGXsKzRuigXa
ciIYEwosawoF4cj+CKKYw4+pufe+oBVoYSZkCBetapr8SL5RFvL0teHRdXtx1Rnq
DdSFoAS6J1G4sIOcCIC+Aud001Gg4c8KvwjTp4Heh059fSJOVov9IZOnz72jvMNh
w+qmL8pWHLk73KsBM0cTb9SgfwiffYJR60Eu+PuJyd4z4vflEX0WoWcijm7JDP3o
Vqkan8tVEb8/WRglq6Sm9h75UfyjzTj4h36reNtAbtLNrKDLXPpEcJfZAdfVLehn
RNH1z9KKykTFh8EZTJCkaI3ZgCBErH2pYGBalnEp+96BXUdBLdCsk8ikziG8IKp5
cW2m2cyPYv7kPJecVOU37xa3gioCTUR5ta77ltxdoj42lpVqeQYzaliKE7mmYxdC
tlsayr9zNV95lLpqU+9xROz/f1E+H/gQrLW4n7WRS+vLzw8w3wwDr9Q136gIbAcD
kroVR8O+L284znjVIiLVOY310lpO/dr9k0OlIzwUQbqtBT6kG8FNZvF1PZGYCawj
EG/Pa0qu/eZzaHVYyoWXXp0IyMIDb0Dg44YAtqVPd6jy4UciQuBcvclADxDr9tlY
0LUWQu2kI2ofjLniBILVQhBe3tjg3h3vIqXeoPWAdC2XWiSQRJ4rckL8IlV4mUKQ
3zRNNPvzof7oWwEcjFJzUc74CNuil2iz5eHFjIe6y4hlWihN7JruRrbDvuntJsIx
meMduwI331n71GG+ZAUs/XC+U0jeVc26febzzI8Is8FATM9467R9B7TDrJVlPF05
iSyh+e0VMiuEdVi5Zgzs7zUO5PLup8DjLPzqso/WejdZ8BYMSAJe8itTzLtHqox5
6N327z1ST1oGN0AE/FwKamx3jah/xzaxXOIb44H36CTs1xAmwnoZDugu8gg3Br0K
aHd04RxuSgcVVIjEE1xoT3ZvxnyovjT8O/yjp78/Bfhqj2Vz8SP5OYJ/zK7yfjRo
LBlCn5cAzW6VSlAEkXsHu4V1+f0U6bFKO2a/UYZvil/yDJh7w7RdvvC89QK27Jyj
iaitTPvinP4edGLHW61mP3zAdIoPT33ck+Avv9jTGLW4ppv1hwS8BqNYi/fJGvAF
GLVP4Vp8A6rSzsX5WBLvBGGNUiNiruKvb+5zy00nuzWiUXT+rE3zQYLtiMTrPc9M
ha6gyTjcTvubKcILOt7HYP4ZFTMrvQKiwdzdnVHm9r5cBf1GIyKUh08u8J2lK+ML
WC5F0jzmuIWLpxrzG+9yW2PfIDrnEHvFGlVos375WUyP5VWyna6S9JZGtzIvyQpv
3+iiNUgihYakTWkRZvCRdRJvG0zIrGRDZRzGINQJk6MwihKcE0jkkKX03XDIG1wq
frEwlrRCi7XZhE/efHJ0kOjBtVq/K1RAuvQIgRhzi2L7uSBKb9udcqkZTg6fgZVl
CzjtvCkwhzCNGiImVtRanFhOgQuLe9Su8+XOQrMJwRSiOLLqiVMVAwDwD8eM8Xl3
sPzkSzRTG5HAvHovYGJ8+B3zV3niOG0McAZMBSvTJzKnGdjcrOp1CF7iK8fgZa+h
gHTnTqNjxVH3z4qNzWXLhx4m829EyTS+8Watv+Q94xigKXS9UoctCe/GQnFKDCYD
zrHxpRiTfnk+MXpDOhtGxPOdQliKov1oRaQJN5Tzj+G689gOrf3qHgzg/AUergJ/
l66Jy9Iyj5rpAiji+TslEkmcflLsQWW+F2qGzlbgeY78IvfD0IBUAScUPity8UiJ
CaQI57SQW4vNYHjMs/XeEa6jNo6gPYDBGpFPQsxY97b4DofaRk3DtiyqaBRkeKuF
Ppb/gh0JACxPy9PQtnkfdfzGvQQ1e7Iv0uiQpDc54tgjafxYRrqWqiFDH6b/NTxN
eJuKEcSe2MSxTnyttYf3THRl1LFPM9QdJ7EaCq6LPYr2KaZtBu9yzjSg3emTMZLC
hpl3c+kdSkXGNcI5upOGCFx27NvplPmwjP1b+rdIbPDnzE16PNkZ5EHjHt/AQSXd
jZs4Phu97V/liJdenlEN5PSxt6uSc6Xk8+1Mqjh/mvW7dq95OObe7wFhjR7KQWEZ
/zLXjU/Zkn1Q0u547H/qGnAp0N74e+/kme4Wjo3i5V9PlNtBhMccHERdzdlICftn
En519g2PakIpioRuisB/3LBl3rQa/f3o6cmbLfNpvxOo5JPQTZK0hjg1uA21iDBh
CaLLRAmuaw5ly/S0qy9VfONJqavs0Y9Td71Vq6KA52TQREYw7GXE7P0quZVyquqs
VPMv4FuV+r1EKkRBqvbrfle9GFZv1nm+21ef8dA6QiBlLwUUBTxxNDEUWu8DrvEa
bpnfJkIC+ptiCN4m93tLdG0hLQPihExFbqY05HUBdX3+VUMdlG9Lb7iHguH/SY0v
b8nWFPV9Kvg/8JT2v7TK1r689hZ/VvYWs7QTyOQxfchrapSgyvHk4CEIy5Tl42Ll
w1+muSOozGmayL63u50fYYLBof31jSB0T/1LtiLQBS7w6Uqdtx00y4Iq+lMKfrz6
Y0vqsNvs9F+dqtHyfU8IlMMyS+Iv4z5RkrjUGqIs2j250kHAz+Jt7Bu9/hMKih+9
8IFpb3oa8bx+W+w9QDgM0keyfVAZJlF6roy/+swZXHUY/A45soE25Dt25CpYnjq8
Nxp/9NsyQkPEIZij7Lbzy+q5sdTqqjAOoBAnH0f7vjIoquFCa9UsUSESoCr7oSz0
5iSEbo58XwTupSeBGYbRvaDFaH/oagxxRH4hr7FBWkcnoZhvd3TtWTVhOkIwGvIp
OUe5pFR6p/z/hV/OrMXSDk2OG4wzS53mOAUj2pNkSt5Z7XMmB6UMUezfAAc3pfTn
vDIoMhZSZiHYm3qma2cKkucmAirO39cpgdGmfnTROdR8gBp8BWH5uXpgZXofFkT3
rHd0jHdZBqvwUwcawQeDerPfeZZAcBueNQi7zTG1LxAAs8rMx47bETHlp904p4W5
rBHbRS0RiMpsZMVaWYGMQEs4msO4fbdrz9DmKGemcU7NGdBHA+9pA8krcUOIp63r
tYariR0NIApxz131UEwjhDs5QuwxqIvzOWzgx+oTodJbNGuBBCJblM2G23As0a5N
hzexgAWldTQXAfXrphTk34TIwlccGViTThEBQzkkJh6D/74xHjH50t8Eexd927iU
woq20DEXSjaC0A2UnQYzkK0GuUCKUwclNKNTazvPpAzS7EgvNxpZBNnHGFvPPP0o
fWrnioQupt6sY6YFlsBRDKusaXka2KMRfe7HCOuTJoXyOWc0iigXmXqaHGyIrOYB
sVvzcyL/Okg3OBVWTKH5kiwG1AxQipdzIOo/zvRAmfY8pzFDzUgTL10ff/SWv5i4
CTCXAL+ZD5St2HZVWkhMxhnaIIf6u13y73BsbDlXgH1X30rn41CS2KY9A4xfeali
BMzsB4Tj3Wdrsx1tAFMCRY+Pwt+hsGWvLqWHMW+0l24U2qawA5nsFcp17epqafLz
gG/o+EHM3sYYKq4vKIxDHxhKKY9yiEJTBwhPKNAF1R7Yq9EfA5SPuGiJZCYBNppL
74s5dijOJvFA+bjcSdIhsRFoLYaLyLjKS9F+37kwb2+q/pwb9+jzznZQzMqveQUg
4KAsL2DCcNwIf3WhyQ9fFgQouf7bMQIUvnMqgOn1fsL9QMesTXAEBkaPK9iW8gCK
AwljrjAfnmz0nQnrQ7qB53Kj8u20zpA1M+ZGjxmEuwPpXRZmhEerlyJ8m/M3kibp
fCWbDAb4LBpnwKzf7K+3Qn7STbnOe6n71f4DCdUPsoLMDYfbqSamvsl44BGoxR7D
hpx2aKS2R820jqhTDzi7JUVdK5TpjqoxecK8b3jKSCMk1tep6KJwLKo1NYs/ejF/
0gSG6QezeQfbVco5w+6McD2BqWZvig+C/qjMUdYiHQsQqIoqakAUd9h66O1ucKBv
G8TH3EpbMRU78Jp+u69rsBVzeVco5JSROhjI1uvYgpuxZCbjcpZx09DnIIJsY9wk
TRUWbSnkw7yXAixiLa2a+xulYFu5bdMsco2jxnkded3OR21yNynWkLXAT/D2Pcqp
F5AFWV10G6Jt7hFN5JNtajfZPIwf/lSNvO5c83qjVQTAQFtUppKibTuGDCbw06/6
hSfXUkf6N73+mApdVfamhNkJQKB/ssKxo6SkF5l89OCaIUIXSwIkiSMOpbdInVvW
qfQK55SeUbrPzyEVQBIqcYaWkxB7lheJc4KW8wttitAdcMh2pdKchoBaXIMEY9OZ
0t/PV026MuGMSH89d2NrzRJj8p/R9hXFnHYINKBGrj2iTHS1DWMSkuHn1avoxXhF
UwBB2gz1Oy67ppQ1sD0SD4gXCT62col4G3ARBLCLTXj13cTXVyeoNEU1+U9yU30v
qR2OQlQ/HfkpbVtCm0HfCbVhW+CGTvWUL6Iu5gw7snHP3fukcMvkKjnZQhMSfIEE
PwUDWAKis/nzXqK3pxGgZtI4LSIp1KR+6UqargQNbw65DOpwHFF34m85F8fgIVi0
4wVFRaQtZmjYPg2KjcgEXuHhLo7V1vvElhY1xNQAQIYt/rmou6E3Ezw52YvwiXfn
SoBclLNNBfCF4jeS4fd4jcCVWkjsDclsui+H7QCaxbzKB7p4MRw+7awVHZu+rX48
yDvJOrCwVbYENXO8T43WHn9HSecCaf6o8al1nYlaHCsq1pE1SA0PVp9vTg7RWpEZ
g+Faj2OFsfDwwLwFSaLQ+FL1plrLPH8s9v7TuZ6Lrx5mWVX3xK42id8aGCauk5Vn
50epOmGBIFd/sH159g1CLUDY1F2EctwbEN403/XD7sz3eAOOZ4szOK7Jlnkn5PH0
6uVzHg3/PMrqdvDstfgtTx2lNBf3j7+yiCmPDBj2EYlxpIkr3MJFRczq+NlR9yLL
aBWT4VtcYm9SeqImn3ch8eCfzH0z9LbgekVD/LpxjU47Qfi2E8xEPn+rFzi7NCR/
lCsp5vHx3rUmXwg7Tz+1zCRbPzetgim76Fd/vltTIvyDamxdC4guUwQHs48/kdP8
F3DuXSzNN3WLYuo9GmP/a56ayhsbSZRt14cZrSVX0UvrXJaWW+cK5jimrx76by0G
LiqHNvaW2qitGFZTlk3918B8znEhAA+lXyEXa1FjGupR1/h1uoeMT8ixLOUOMcNz
RlyZIab2NgD5NZM67AHs/md5Out/zja7RGST+LHIKAZzXwtiJEJ6ih51xPZnA/ej
+iYYCwqrhqv0u4DFJCN+mrY+sZyfnkiWrTQeP3To4UqwVx0iACtD2sviaTi+ojrR
84vhp93ZsGq0McU/+f6h3P5cKsxChWLX69SIVclXscWe1HR6jg0Ug3DmllYk7jIi
u5gWEcCxmlFuzuXdMwPbxJMBINi5QW1GkO8+b8jfrsl8eeobmbOjT5gHQctkHJZQ
oYQaP5C2ss8UWNYAkuuQEWOvqOa/V6QZM5Fli5Eq7+u/FP9n3VE/6Os4pCBNqyN/
s4ccwErTnJj8Kp+xKl7uYNkOJ7+yVTp4tsO1wWg+uXPkzqzeyVDv2RDC1gjox6K0
BCSVs7ssibBFkFXRNWFLB1Xl+RmzHxn4tJtOF38dH1jJGvxtke2dcx521r7FwhAE
1Ga4PSo3UTnNwg0SwYhtnnt5PNBjIvIrejN3HzrDKz8RM6rsdQ1yvwHelEliPoL4
V9q4o9R5Jym+zk3HMw7H+gHO/Z4RH6/zX6f8H14/5U/icKZuwu/wjcEaZMFba21O
ON0HHsTp1RSWuEYh0fCR8OAVHi2+pugof63WMAFJ3R96dbfyKMTdhP6vIoHt6cg2
kIUAho74+OtK9V6O+R0T9rAQY36fXRbJ624UyLdIy3xG/XUtjaU1MdVZqE3O2SAb
Mliy/ZN7TG0s6kgr2xTrbWN3CKiIbxU1ABd73jfyVq6TuN1rkpQ1poM1CUmcSX/K
uYu3j5EmLgbFXiLRw/p73Uk5Rco7m4TCW+ajPB3LpTb5Ko080u1EdwLJN5/c4SvU
aYoAYczP++6zLYkZGeONRnQNR9YSK1r/yRoKU8hKQvqtI5Mzpjs4EgswtqvXGnBS
nc7EzmHOGsE7Z5y9t+3iyvrpvIX7nW7jFORhhdWxTne40gEi062lxkKp038O4y/n
alzqtkcGBcjlUpcMsu+3ctl+W7w4+uYLtmtyoJvsqGyrqtrg2SauxETt+b+C85PA
p0L0urT9CiCFWLjzYDuCIoxTwaI/K0yn7rboRZtU6heCEgqdtTF8CmgkypkkUSMN
DpYmZ6whJDs82+Ta03UbwUmkFwI9FGbytkEH8QFeMrrrL84Qh5YMlrcSqC9VxzM+
0Y4ZCX9DT75ZzNpD5Mg5/3pxTohddmpEc0G42+VBGYdGyRzEq6nx+J+vTaVF0VUg
R0O64tJOAFQr9UUe97mvSByXT20iSKxcLD62jp7Lsc/xe7/7zcrHJKGB7Y6bLPFw
MNbypn27HNghQ1grGh3lSA85TIUhqtseFoPwSKu/vVGKou4U6yy5IrRarzBEQ31d
5w9SEdfbl7gn0exe0cuD0Qc0SsDGbxN6UnOIHav5b5tJ4HQqf2Ki6PNH24ppUVv3
XFx6tjL3uk2XBNDGBsmagCxnISGE8P7TapDFrqONsi8uBGznnCKiFE1LKGBeMO3S
HKLARL/ALjTa6vWv4js3dyTvszv+YOw7N690SSRxkGJZNIBtc5HI9ujBKEC9ioEd
PGAyXtAtZwWc0WAJlGLNFY0xhWB4AVs8gWeSJ6uLSSPXtQRaEht+3HAyvnAM0/pD
f1MSHX8ChfjoyuRW03WjZOrophrlLUj/t6GJb5+P6LnNqKceKKypZebqWIn/EL5j
X08iCaTMGhFxGRML22HAthAdOGXp5Jqs9fpJF4SVfaQgtCHjfc9BkGaIdb+++6rS
4px13oIK6b3dWY+nIpj+Y17hHH/nKLYWZX7n37NcGxm+SB1N13z1V5qhUSt6a+W+
nPbqSn3QslBiIIaMrDrSSszb664FtbiI4dsfc5fBfx8juxBOCWAagQm8MHXeCcl8
ADm+dwoW3DVY3a/rzxgUAYChh1grTrzTiIBzb3P1v/V+QQlnuGjuNUQSvOZIjAh6
Z/Bf2WI0YqIqOeewD8ey8R5LkoEsOf4xp/yA8meHJaBJjRob6KGBOjaaY0MaNVGi
b7C43wtEGSDWP0n7/chQB1q5lTQiK/Iy6qakVN/Uw/3ZXn8Slq67VR92WR3GTWEd
4kIPeQCmJQ7ZQ1/vwcJprw2YatirVtDB5/cG1sEJY3xc2zE9LuPtz6fJ3odjV2sY
wA7lPBi5HdQycyIinavZBiHwUTia9y2vQLgXXPv12aFasyUu8E1LcCNi3BKp5s1/
AjeFc0YaPD44N3m7qZJi/k3DLp54tFbZ9o8TCcxN7E3i2cE8U/ScwTK6sVvDqLym
dHAObJPvEWF1xBZJj8w0xAg5W1Pa1vXTZtSywH4usoPcNs1O2r+L/MzlbYu/u4yz
aq4Gno64Csp9C/wMozUzlfV6e6Y/XL5eXRmaUo8db+vBdSa8ssuPpOTs9RnYYAEP
hLTdIGJ+HfZs2vz4EPxkzXO2uafhlr9l7v1HhNV7wL40Hio/cYnwYPZPJE3A2yQm
K8nvOzAZKJ2xIdS/1DaDQlRNEr5UwBzo0Cu71CA5doD7QAvji7MiQj2U4on01US7
vtq1S5qpiCAbMng75t16MzAio9FGf1uY41QPf+U/MoUaQDHUM3/zJ2WjG/HrY/hw
jEjAuPMa0kKuCH8XPahuGul88CD/rN2hWIClA4qftsZc6eYo0vgeu4WwIrAyirWy
x7G2vQPMgz+Sm+4A5w0R/Cf41l8PswrUtQTQ6CPH8whb1mm9mYuXOUpJHYcMRhO3
p3l1fezk7wguKn10ixLo8ZGLZLK8oW4r/K7JlPot9vpmRPCe2FzJ1JgqQ+S+ULlv
P/joHe0lzb63EWdt0DAwYG0FawbGkr9vedG5G5SG02hny8FNZrTmWDLUlG9Svkdv
GrBrsZ/HIW7xZsrWtL2/mgMOxKQrHjm9/lBR+Rk2iV+8oEPaEw81bvVuBCSEFBrr
kkznZSxLUIqDSV4+fvbkjnvUnWNB6VC1UBsbt2VTHvYzrHjllkY/WC6uomIUJwf4
DM5bl+hUxS7QzsaBzbl6Rk9FtlR3jOgywDQsNMWrW5jXvJb3eluOolx/xMzB/CwP
evZjoWoCtmM+Ibe/qGwu4vXBC+Ud+cKBgPgL7jlrlCS7LELqGUm2V8IYoVEPk5BU
ZudcDEgvEOkGNwK/+5ykOfy6acjYYasfDEvm7H/dxxT9ph01tiF5S2xPwlLNKVZo
g+6e/8y+xvP/wkluxyaUzyyev7v7nf2Hhy3MBymsi5YiNDqN2/gH+b+kUQ0AMTcI
1jA/B0wQyxDvfbHTBPniCqosW4fFmWXbhp/UGQ/MHLNPujANCXq6c1biDg0poQPZ
8+38dMaXVF6OtmS2h9XXInuWjWd/GQqKxkc34NI0kZyW50VpbtAhwk/AURrNPPvj
QlhexRiCGLrGHi5CZ56nxBN822reuol8Vg3tlmIPH3i7nra1i48qlQac7ZFs/8g5
9N8GArJsboXsAc5bcsAmQcVKIEwZ4ozWWGj6rXMk5db9a+XQGaH4lcXp88V0Lgsv
lavZra1mbDAWMVCL58yn2TcBphgi/MvWTsle61qTnXhd1JbwVOhcK6NwHzhVO4xh
AteMtxa69HUawR5OBRCKgAerI4FlQIyvpeVGWd1hMiY84X7MRvzhKeuIyp6Ztri+
G/h2wl/I8eKhJI/pvuvJONTZg/JrOBelPytx/zUQuvdTeMUKdVHd33+3wN9scOn/
8Jyd0X+zJnSexa3nBpz6NmA9JNc60lDmld9ImKOPG+4B5YPB1SbCl4HqjZnG/epc
UuiW8pgMRTT4MdUryaZ1Wqb7SXk3B0DwYRIBWmTlZNH89NV+w/0w8kpaYeArWnaV
0Fa/Ws8J+B/T/gg68ONHQRq96Gb7ZbHMQ6vuxV4NhwTXFe3xzeOfpH/MN6us+xa/
tUrcLopSLq/fa+dyhnGyEBeyNTxhrrmuRCAdTs5B2cg0TUGT4FSsdav/Qlg1MLUI
I3eNeAfFUVzFIbshN3V4nNe2N9VvRb1Kp94Ymr8KgFU4KOQHvpnWF+kTP2J1e84a
MNEAZuD977IrO0n7wqOT7LUXuLcoLLhMC+dkR3IY51belrIB78SnP9lYs8Bw0WII
Ak+RaZ/Ts+e4Ch70X7fd2PnMvMDEckeaZLsMIzOM5YveCIx6xqKVnUelUJgKO94G
bAzcmbDX0Elnh/BBNVOw+SAbks5ucffgZFyP3I/GMpu33DU1MuctKFBNa9+U1/zE
t2G2WGNntnr7WeOG27kv2IiinfEcprnYf3YXaCvUaemVvxiZOCciajbiovMBwFbP
nXMG2KntfH2tTT9kpRFSjGXxW2gvHCs5C+NG5QzvQJbY1fletcPUCgGJfgyRx01m
5wJIUvcDBt3YDLxsmYr6WqCUdhIfgTdTKlJC81HhBGKxxplNl+Ri0DS1klHnBvHd
xfTTQOCxjfO2mH983BY5DYM+kIoeVTTz5nE59Fzj3AFlsMTobeVA4pyLRNZaSTSQ
xpFAb9hZu1slL0pVNF7lCoVdnpJm5Pxszz8YERjTIz0Bc06PP23M4XhSAkpR+we/
U7ryTK4OsecWWSPLhq7JhIwHcLj5/z8YBj1LSKsOX3BYZl+fINcClXRQYKR38DyQ
6XyTb6YcntYxECxpLIl8GUer9hOwE/rGEEvFbYGwvZ2Bt6LSxzrIZe5rBXJC4xOS
0Rw95P9/N+5ffsbaRNk3MVt7YQKULKh1lVagjdyz/eWikLgAHl14rguydfqFKpus
6knktkt1+N42ISTune71O2nOMoZ13R712BCgWm9QWaMYm1tUe+chBDZKjrjzoN/I
3GQPjdX3aeHivkhoSWNyiGmZbdnEeNa2HRN8HYFUo2DuLK9sdym6pYbJzRxTeLSj
fUyRQzJimT8KkWU1dYMkPgJwowPiB+x5BaZPKRMLBbQJXZV5bNGfQsUsnkftHY6W
2+yGKVTKD48VLWOGgRYXX3+HLvPRHElCoOE/Y1ov/IY7M5THyL8QKC1TgJpjKMDz
eGwzJJH9htrKGrJBu2WLUe7LmyTurG5EutY+n+92YQxou9+TPzhvElGIkRpSr863
y0A59d04iN6M8wuDqWly+vgTH8NGs8J6OthGkfd+aV0Ug1P6+qi3JesVFfSuyuXb
iuJAIBB+iff4P7KJUwJ9T36mZX/LG/YfuGqS4dH5kqcNtrpmUErnBBpZHHcZhifo
NA2V8ukoqaT7O/JetypLLqHWsO2Ck8HwqZYFWMOoUmEwovO0o3GNmN8tzVKAMPSK
IYyy4R/11CCYDU1QcTPwFsoZL5FUbUcV54qiQyUIxUgrm9gCIIG9WYCqKjF/MiFw
zYtVOzTMN8xZ7TS7VAhrWF7R8rVAbXyo9qAxtBkW949pia3Gvmw1jnkr+alVS3AL
+nxRKhkRwCpxeyjwVw+oFT9erJ68Gm3VEW9FB8l+DvkiiSNgd7dSZsMHfr4++6Ut
N75dcQ41snOFuf2+FHHhhOorgg/w/HugtRY6oVnuSwMUJdndngyB7g3DBs72KDb0
ZDh9MvEBSMLL8cOCqsfy0reTX1rvagNfescw221pnDTTsCW6Y1YktDb6uDlGGI5D
r7/1qDFB8JW3PE/+lM7uu+/09OTUNDqh4Fvow+kRuawIujQd83qFnApX7mbKpUEx
vUAIZ1aGON+Z1OcnPDIHL3crzK1TdOVfJLujLvqB9so//ouli/46NsdqVQloKUcB
mJzvqYoG0Rn0wM0HdoSt9IV2AF7GKjEYxZz7gwaxK7or1YiSTWaRJ4zQ71ZST79Y
n4SbHkvra+5CJMQ0sbw1tlvKzm9UR4equab149eDf8wZUK5dg6BURukXbBpmWsRH
NUuhAMXoaMJw8FlmThSx70tOlkAF8EAc4mwvzHYbLPDoxQ2HpTvoHGYkF2DxDvat
WE++WW9qmfAKeUHgSM72tBIg4BYuUp6vugP+X9yand+o5QUtfp7OCBrJFnUvXnGL
aEcShOVfFtOexBPoUXMCsfVJ5zHrSxjn0S65pZc6x78M5Nm2Garv2H1SDu8/Vr1k
SVItUszRhm8O53ydh6zn7weQJeUKKjG7C8PFlUOzhnzDeQFabEITvgAt1n7WtSP2
bRTkc+Sk45CcY4Hjml0eybscO9Ypg5WjVgHsUC4+myJQvC5MOPtGPzyBuAvBnN6o
X534RVrOb8DjSoTm8kaiVixwt6xmjAwhCa2wzKlmVrewLnannJ6b9W6RQkmxW5AM
EUqRHGtBtSoTXCdilt6hZ1SLGrL8fHA2VR0mHDJMXJ0MKWl8BTW4JwLJrSP+9wlL
Biom4XzFQJfxDSzL/Z8Ur9XvW/C190Xfj5NJSeV+uI/qWg9WESG3yrJyrjPzgJzh
7efo1W9HOIWTTMqI/jZIZWRUhKZovfJpNk7FPlCvkhKZKrV9lGOQKcb9kWl0AgWw
OQPJGh19jASYGW2E3dvTPTPTzegsRZKRRAmmDG87qbRsW4bg1RiDYfj0+BZ+nEh4
LYTy6jT+vnV3EU2H8qNXSDe+YXgHOSc3mCUKZoZIC+469oxGf2sDfUtOzDFSEv89
FYHxVjs9eRxtw06DMXHCy/DxETZmsJg8hkjogTv3f+vdzBqSC3tmimYhgh4xKA6+
x66IiJXnCYP7i/rZUKNA8IdRWHwknuczZMz3y7d5TBRgEJzowjcyimXOIrUDNGNx
Rg9hdJUpJBMUoE9tCg2+i4/csvcwEZDnoGXDmcHS1MTNYqoT144JgiI0fuOrROxz
iUFgDQRVJvPQ/1wiBtauiZb42xstvZqSBcohQLEtomfgSrD6u2jKYAd8zEzEcCuC
MT5++4zJXdUCW84tnA/x+oW7sTYx67OTT6oEEr7NGUhM8M7yzVYdzh0ZpqrSc0yu
mJcW9XyVH9ztqjuH3YgSXges3BRsa4UJeVHvObmbndegcA7DaWKdswWFVkt4UGhI
KecCMs62kvhPjbgR2rn4tQng8NjE+3uMy6qaLhqLuJ49308iu95mDL8r8UfrXPhV
ap2NDiRGwx/M6q0TLpF4rgMzd3iNWZvKcwTZEZClXAq5AKXaHKGnihXzkyaHMxYF
gHxaHYBj+8i7F0e6euH4QsbrSD8MHhr75yzC1iYI1ICj4Xpnsug0QH8cN+waZf8Q
/4ZToXKydh4cuFvDgK3ng8m0By30JF4oPbsI+GHgTzg8cnSeydyNzioSxkxwAKYy
JjJn6TOkGvYSFRQbDrHdTuOi6EjKm4bMTVUmrdJTk4IvSXSOrk8LYov62EWuVCZu
FA1ZqxmQ7LbOViNSR8EEGu4ublsGHOQypNshsTTz5z6bmpps/SYGYVUKZM0cbRyS
akhhGUdF9n2JU7svX0og+RJGQC+aJanb0iw83m8A8tPHzc61glnqtPITFFcHCv6M
e06rbLkjWcnIt+J5cREd9pZ2TPkfcBwvVaKdsmLATJNw7htvr3dGPm6+XYTAjffB
icr5wr/CRXpEazN2DMB0Af6yPEqaLCAaJIhYKfUZxh3GGK4iRho1eMuDie3i6oz4
UC1CxJ7ldmazlM1HtRxC14aazYCKvVFQc8CbZSKNPjNK65Hq79ULxGzQg64BJdgY
LUOyqeKpENxLxECfaM/rZSIACipk2YNDPrIY+YHG0gsTL0zaPt6BL3Xfvhj0+ADr
/M3Th+Sh57yJVyYWHePScpJT/w8mTe0Qb+cIfPq5yGT9aPRSTQlYUhEBJxYx5NV4
aJyJu9xP4n+Ru3mi+R22oPLyNdEPwSUlC+x3Xg4vqzycBkL5+2dxS543Rqrlb13G
wvbR+36izd4Y6TJAZbny4++Jye3eh/wkxW0OzO/57ZUYm7ihtIoxig9j1/Ar75br
/Me9g7fUzXiagmN8V3mbA6HPcFLpt/PTUYZqqfVY2WPu+J2zknxxazR1tGFTOgAv
9/F8EBPdrZA3TBEBwKqWFFKmjlVfhUJiSXqHVRnqAup2zEK72CbJRhYl2pmzUpTq
MKVMjY/Bh94ZLIfCBIG56SXzHJKF9TqalP8D74eM6iiav6rmgyHSmf78YQT5MH+k
SWlaH9KvjOTm97LN4OxZd/eN6ei/0x11G+kpUG3uTlUbdi5cJPWXfkhp3+lQu8l2
wFzET2Qqc4d/rP+MGPnu8wVdVensCn9kFZhJFt9uyzCSw30opKAMKgrJzy+0Sxy7
z64Y7IrsBLgiQlHoRg7tP683YaKyQhqA6Fk0OxrCuT53FzXsbercqCaRp6sefLrU
d8htoriEtxkVHWr1lDhT6zOPTY5pxHDt5QhdcTgKv6323RtQ/+KhTu+BhfmbmiT7
EtCQfsmenTr/MsYWX29W8Ss9KI6CiEiMI+ALKNqcVdp5RJGJN1HT24UgOo/OKjXI
fRcCoGSX7sOzMSP8HBf3he1a/lX38/2Jl/mfl/IsXPHP9ERXDcdT6u232a9ijwIw
g4JaDWgZ6aJjbF+XCk586djDOtQS7ZgSw8GgjroXMJrZTAJXcd4WerQqbQ3C9kxe
/A+6krcF/tjjSqMU7aSC7Zpr/HgHJcUk7G8Q98Dt4D7PeS3+IgDeTpVGAPlpW+iV
UCjStCaCqIrvx6dPVs/L3kBeI+zKU3Olb5le2yrrid1YulY7D0Bg3KtYAH32dUGY
gPq1cosaNXm1DIAJZnLHC+tkX/Bqqi3tmGv1xc7cTfEKGioV7J/EG/8ElgsMKQ+T
KnzoufzuHYsTgeMLXrpY2Xv34CxNfSkTxwXj/kwmd8haTJiA7gnfYihFyuUHprt6
+rhCt76WhbWEUc3yrv2E+e12xLjgZvdiKMhOFoPxGx3P7Ur/7pMBJCyi4RCmIfV5
xzgF+nmgnOVM04C51YLcpmtZP0EGFKdjW0PLGUmd6NBqMaBMJYYYiMg2AhKzEw72
sZw3383SoP8fROlM+0WlZSlA2ddBzRufyTy5+DHxzykQ0OUpSyAGwNN1zOcIak+M
eYGOSt20kxFLGbZP0K2lFVSACrUwdE2kc9U/D4ql+SWKfISBk3rQUESfJKJl/2KR
kIw7AJJrWda6urifUnfEFru2w5ERywa4Bvzn9EyIy7z+gJnuYDOqm0UNJNm10PUa
sYtxCFCuGHyVL5C8KKKq1LEzDFTI9sK96XctLolmyNrFrXq36UM3oO4BULaJcO+W
KH65pbtKKkKQ0hx2ZlH7684vlKIodW5R0VOxIRV01ueDZdTxnjCWKzEDQOPcVw7J
K0cv3BnYQKh+1cyr+5VQasPS3JdkZjqruqc17qNgrq/mFM91lN49Ahlt0pX5AL5z
Zqy3S8WYC7sVKPi999XIF0yNhys3nHokLVg5ciz1ts8xaDcxEk4VEsDW9IcuzxEO
C3qOFII2mMWzCe4Edkog1dEbcPz1Y8I4cPO5dFyCMyMbFru6VoPcTJ/6F/EHJydG
2OjB+Le7ypv+LlmPTRPw1cldBg7mmSKjcbh9OfjxrgPL3IuCpJ+hrYd9IO9GgML1
KxlLaJbaSRhPPq+R00Pp735pIWEFYq0k7S9Px0scoo2xwWchHuGQ7/GFyjCUoMX0
O+4YFNYTtAHq5XAsk7TjHNfYb2kq62DbH/QikcTV9X7SKeKQtz+a6EnP0f9vbvER
wf3gjx6Cbdc6kcArOOOSzfzwbhkWeLj6hpCg/HN6J+J+4plQw5ucLADtMbO6PHri
NR3AVQMpPCse8swcTCj65T56mTbnEb6jeaiPG2WvAE3H5n5O/kSWDQ58jKekxm4J
18WFsHl/f4FJrZDoB5+zeaHbADMkuUMVJkcwtOZ5z6BRY+gaoFYHSWjQ2vUF3QW5
PEEw64qIxoFjnQXp8+zluvCr09jMM2GR8WyRHpKkFyVe5XvqoC+4uAICIYhthdHP
iGnimjAzVSTeBcKfH3thvTBj5tou9yoFDIEE3+LfRXEpcdtk0GrWi5SL92QYE9B/
eWyX30kv/X3fH/E4on0h9GQYWpkVbqocieJOiGfuSOAn0PrZfrWdBfK6/O/eaNs+
CWfKfPi2R2d22Ag5YtAm5HGbwfSlYMa6DFSuB62tGY/SyKMnk/CDvoBEIkWUskmQ
8mEAbzCBRm8Qlf2EI3kAnQEklM+RE3za/aHt8D2OXToPWIIJUiYpVEGBDSc9w69O
8KqvOjYdreBWggwK2rHLG00FZKjZmrs8Dx8n8a5OfMcY/6PcNSYhQA7xiyAR8liW
12dxP1NmecqhvHTRzAX4Wsx5hvcG8qbRrUJJPBZOotJFiBuP2d4r12JnXmT1lEfq
U5+sD9cZrdRFtxUInMSpGhHGJ/dJW3yciG2mETkUR9MSw9hzRRStAg9utED4AOHC
lpP0aRoAQcju3/zrdGQrwvoHSRFjvwMaOaP8vAJCQzj8bIbmRMPxieV3zHatMoN1
8p08Zvn3i1Xed1BVfzTQfRDvSkOhJgocp6v998DLFlp3SVIuY/O/O+ENLUfAthx6
qWDxJw50us201s55oo7b1KVlXHUWR3T+v7VeyXcVBsw0ZfMHn8up2UNZj1YhpjBk
+ZnIBOdnCH/udBuvkNvMBTuidKOfOWu+2xt1T+hqQP/D5MlL/k6Qdfd863Yi4u/4
rV8EhmaaeZ/bBo8vlcIjFdPBXvNHIQXEJFbeYms4XViydeHLL9o1ritEbJEw24+2
pjWefR6rvDcynjumu+Dp9PPuIKeRewVHzAOKM6hL46XyH0X+e/x24aNXEHckroMZ
H9m2raow+w/QSG4seATk/v2ADh7vdAIJtyK7878DKdFKkC2D2a7BhvZ5JihbXY9E
OpGbFsulnK8R+u0akLRl/TPmirQJmn3pJzp8NIYQ3dbk4J0EqeWwTPyID/ZDFj5V
KAeNKF22h9vEkm/aBG2Eksn++mzfMHaL/20/DS7pFj/YBv8Mln/awTGrbxRPe5dI
9y3+ZrEqausoPk5tth4+KGLY06UpOeLgUcf7hnhBvhiJI6F3+60DWyF/F8Mar7ji
6Clcbes563889SFewcNBmhEiJtQm39mzqbfF8sWbEur2Cpr8yc2ggF5dN/JyCGgi
V3hLmzL14pzP0PQYQ+2fJQK3mw47Kqtsq3qhsKfTDstDvtztvw9AvNiL8cBiRZIh
+QuJmGapZeQIyNsusQQn++5TbHRJh57XoUg+LnXRMnQ0+oeJDMIrt8NSXMIq+YEI
7NdZNVlbtuNCuaGU8IaBYwL0yyP/2CRq/eHZBBdp0wK3i7XBK0fHzt+PYuhv4PrX
PipV9WCxqpyIZU7T2z4UHIGbnAEoU/XR/erRMQz7rG5imwP/DCaIFSxcRi5MXgQp
A8GNZcDlN79Ge9FMROzHCrf0DeYPb2dsZD9aHC2jWqQXabd5jGlAh2Ztw1+88a4O
rk/2+4hLHpPYbtkcH5KjjR17kdO/Diq7arg0qGec3D6LMGhkdN97lmbpx5fKrZTX
3x3NIvkR9WVEsXZANetmXkdXLiwejV0xJ17RvluKfSN9XE9g937sGbqwGltJhFo6
oVCLfMGvvP/pO9DxRykW8CdCdjkqH6Zw05hjAGaDvGKNtaeBYSHm/PGDDs3eeLB8
Z9E/5SeLu9EafJtRMAETshmFnCLmDHOyyHZKS/ZimrtCBix70Q4QWVo+nsJtMJEK
UxLhf7CsIKAtLuzYxXrzHxsxu9rpKHAS0Dwu1oXy+SuQSIelCpJWkE5MrVRVXUM/
SCjQkrldwtqSZavn6yvKU7oHQWr4rmQtdstdd3gFIi4F8VSlQgYeLXIE1qid0gko
3GRFtX7JUw30nk6NBZiPMQu4lisqtbfHCNXrE+fNRtBo4Jdwxsiuyx+wxIIl96IB
fa4TTOm7cMRQccRHtyeJjQX9FsL60LigKr/96zq3R49VFoRLKJdacowD/CxsxZap
2qexDxo/+seJtgMqrOprrST4dlXmIyosR1UrLtHmfrrDU9KV8wmQSHxEi2C548M8
2piFetmfHSkXLKLrL7ThEvNTkkxMSEQxOLuja9YSH9aSdoAm8ZoxoQBBIRBnqZCG
s6d57q25sy5mDBrTwthNaKjLCoylT4vo7KBH0p4UOHIJ1Hx1C7cqyxGHagCf4SW4
Hlv+faoZisiMzouqJBLFRveg81NH0bXixLcN9LyEYYNP8tKRVEaEuQgFLmzqBJIq
vb25+cXXzMvNPAhcfizsMP+LXicvh1MxvPQj0W0068SpqC4bcmpx+iS2ZkjwQZyi
kXxCLE2BPyjtjec4oAu8kIQiduSD2qgypInBTxDpkpHzsvbvaXAmA4N6VIn4ajOp
nkuPaclv0OWl4uMeUrOG0c161uNVZxPKwS7TJPdUDDigBktzZPJAhlMOQ/Vh9Uty
BdAOLenQsjBUbT5VuK0qPgemcq0BkIGsDv0lQDPnEdbBXnYbgR38dTP47jOi7d0N
+LORWmeFQeFoAjVundO+NdwGtH4nWPOak9we8jH89C+15PHkM100KcW46VCPyLX5
qXVKvi0/YZGOWVnQ4HD+SAjNb3r+Kf3dA2zXvJQ23TP4kTVL2HKAKbuHpJazZJez
+mWmx/snPCrQLjiO6uI06wzeeqvveDiPEN5l0AwJB7agk+9y6/aNNkzH84fPEK80
N+Vs+etds8xxzEy+dvKUMmJoXhT7rjEAiXNz5UTVkBqIQMwERa0gf7xyQ9ppWLfn
X1+GjpAx3WDVusSdMOw/1y570k5U8DQJJsFUXN4IOvXh7mHaIggmn8TJoU1gk781
4RR3ygp6RIpGaCezvTDkBQtBpc8MYuGJ7xq+6a/SkZUBrYaho/mjjLq8933q2FUP
Vylr+3nvThEKcr1MQZSaJK+knmrVI500mJ1M5YjA6RgRxMxMrP3npzrFr5AZ2KxY
mtn0x6LwD6tjIyCgdMZvoXWpCrNe57e1dHLvquSm7wxhtXgH8Dmz1d0AM8GgRJmI
gkQmoTED9EHZpdrq5DiXUCPNvojqrnzCEv+Fay6o0A24rormiX9Nd8Sb6tfzvpSq
1Fjogr8iMsXXiBWtjxKTLzOsY6Er4TB9DWuu3meystPlRlR/vSRDvi7hYH1cctdU
aOh/6i8Ban0GeUL9Jz1PqCzQkA/2so5f/q7uPaCFlvscfv84NH1hUv/WUUscRi6X
3/TV/4W+W5E/5q+roaz5MAKfW538zRorSjNXA+g91GQ6mbIpx2n7AUJNBW12dAsd
QyNxBOnrxbmYZ38z5eRpjze0UbcGx72Enf+6IpE1xhToINdk+4wGOhO2bIFLiVmz
ifwsO/GXLMCsGh2Vi+hMYi/XjN8FnZOoelnqDQBdz9TmRcqV4kZcjAwN/5e9EdB4
9cWPgLrH5Os0uROcALp8AdA5ocAaP5UGh6j+89DddzwA2Dftwtuiq1onvvqkA+Aa
MB0TOrYWcuzXkJBpXZbxw2tMULXIqYr6dCqp6P9CxvpIBmTOUXGNZ3vZOGyAgU7u
cOLFATc0Yib0lwF5v9hJ1CCZa6yLllwSvZGr/lamS8vv1/kydRg1uxPlfGtxx0sd
/kmhYYaeObH/KetdIVaDWnM2+ZrDTrMV5N9vVWaxMfbLQ4FevAMdKCASP2e0jx92
iIIe5ZPF2pL3fPMx8BTKkhWtjSo2P168hE8iQqFZq4Nzxi9aLbdFaZOlDu6kWqQX
TvsEQduUwqrjUi2Nb/lybuHNtprL3O5tifIEpxCKPf92eHNBS+KIh5bhtudKFWpa
vYHyjh13ESSjo8oglZC6837NL+E6/Ws69Gmp2kk6iPNlLO/oAteifINvyHH7Tnk2
CzjgWE1Ot1wT1T5ktRMgA8qXUQta6W3JxtS/9VSjYepiojCDl0QZeAODvgkxQfrO
p4RKrvLUStUqDcV7Gy4EicaHR2UWzQ18JHZAzJH5L7AH6eqcvc6Tf9egKO1WZezq
KwMimVkYx4OmPUZyCE9zRUfuUW/+dzX7dlVmbyaa1aJRI3iQaVhpC0gDYg+SY8E9
v7rMdE8WZ4WpYaHLbqhdcLHYDb0yBG7ZoWzlz+yTMBkFRbH+hpk/CLtCY5oZ6kss
j9pGTfsXEbZBJAvrbncEJdSAZOZTpqNJvELCY1qcDxy7LFOQ13vlYMHjp6qIz/UR
nfFc6Y0GN5DQ8bEBcKLOuIkCLvMbWLAN8MeWeSMcjPcIZGnG3mhfP/XaWkyQ3H6I
gdTYYP07Qk60qtBHiZishtSQzb79TaWvRnwiTSXeJilG6Vc4huS9iDAXDPOWTZ0P
ByrJjymCdauvZKkwIKiPKwHGL2PMkamKWfSoA6dAobvOUZHl0qQHlYy1MyNPPiA1
AmNHb6hglwo1FeixkBUd2UfVCtR5LwDzH9CpaqhLFcWC+C65kRKEwMbyUtGVDgYt
B1O2DhtPNvWgC61eg483CZc9JzhS48om9tiHTTl7AeKmvNL3ebp8eCODin4CpGNP
xT0TCL0+OQ1X+OHpX9YPgN4MJ4nE/O7+B3fIGMdNvxT7p0Icx/nqyL70Obru13Ux
PjsiOLWuQ5ExM7beZJILYZvaGxAg0d9aklPQMzO+UV0KaVJEhhZlOeFWFl+Xlytc
rA5sojqUjXZt4s80EBszgzkJnAVI3vdtq2ShqdjCeZUHm3jlTRqpef82bNjorNp2
Cck2IjveUDqzhxqV0fAujGkpRQ51stlTTd6QGgd5FIjPqCTCcjCwrX2w2qg+Nbbu
Ap1gPnvLteyOs3Wt2uCE/kCaisiubDatWxG20JJw3PsLUtWTR8p6rm3nTsYmmNQD
pVYBuQwoC+Gk4T3JYri+td2GvuHV+W/TCCCfrHKwk563UOCjPjGzaStmrWekaENm
R8EWWmvwLpYayC6JyV+gQ3vxrHsw3pgWSIZKjbK5oKcKsNSo5RpyAlMwyAblOdPR
e9a6vMw+gXqWHY7UwxCg1sh1klxf2nVDMxCk907pTsal9f6Iebwl4F05CFTcCv+3
/344z6dI/8c5/efsv2vy546E0ZDjJLhtY9gKmh6YX2/KtqcpeyvocDGNjp0xflC8
5XifqiiBe+rrbhoa8pd+Mr/osTYhIWJ2KtzQtaDc4FcXdFrG5oLlZZbpuSPUS4AT
bAyOfGNGAV7daR9rTXtPBnD1kWayDmtB2BToPQXjFDCyvcnQC7A3zkVt+FCNsf9t
Z0UOPzCyYFeIp2XGTQHSw9hk2nuXgoNN21xttIy+OGp+4dEBYMbbSDdNg6lMmIcD
XRXOfnDYqezjPUGB9ZvlvTA7vKyTYqRNZexjPNugn8YJ6zlaNEKKNoCs6cHJ3zX1
9e2t5Mp8bDLlkn9XqnTuMbskei3H3QGoyLNYaePT5N3igv+wy3V8H4lzjWvl9LPs
EirmIFdWmUIFhvGaiP+DXioJ+rHsieY+hyy2D3cy4PzEcFZJVRhi/nTFZeI+V/Cd
DJud+Kl+n2A2fdOiIMQHgvhvu6GAdM3NYJLpm1cVJdrPntdoIQzL4u79ThOdhFHY
u7FsBVYMJ23fRCHppwBWSBW6+RtHAsyaKFAUDQ4/Qjy6hdWtixF+H6mU2uJuSzaY
IlxlGYqJeVf+Dgf/HM8W1UM3pohWW2uMGRhBe8Xs5VBg25VOBkp3b3eoJ7g2CWsW
8wZKGcJqhdnNNONcZbYiZRzGahANwLHonHzYhir69UJ54aFn+d8WhEq0knQcDiAx
I3LjqGffb799fZd9KeNPEeABlZZbqfTdxuk4yUg7I6zXmdLbaWHCwCRv2VRBaxT/
vCn587N3iDwECxgllaAfiowO9H8Q92hiMn7VImzhNbg5nPOiyUlIdtZwXy8xGhHq
rMtSL7ZBAW46gAQh9mhpd4pjhUeq9zV99nCPvuHYOhRk9t/oVdqgDDvr0ORaMbAa
7b8A2zEvP95HCgqyiMLbbwya3NCaBPMTJZhsjNPqakv1S2L6C0zJ8IEOgK0WkxfU
Z9RB0B5xstr5uRzSlTTWNkU1Kab8j96UgQ1MLpyUuscWQAS/6JjAEQprVcaB6nRs
/q5sBlZLMFcW4LuAUwV9cXG3gaK/kr8FHrSnf878WRkz3UYC0Ot8VqOjvlfHmlUc
v4e4gBTrXi7Gj7No2srrGJpX6Dp5q+fqFwRpqPxdw+mobQ+d2rbxNN4jqnQtr/p8
7zh5Py6YepB1/CbqMh7xpgpTZF8g9HVpluDKydoYeOM3W/mCeKkOMCQYjzwV+hVk
6Iwv2dMRF8UUDnBlILemjIG42fNeytITu2/fwzJ6KqckKJed2bdLTFYwJF5MmvAH
9C1X9fCINJAGuC2AUHHECinzcMBMFgFOtRcAWnmD3Vp/Un4dVAUmrGGQEeCWGfLO
eN4JBoG9q/8sxEsMErklSaUbNHLqKe+GEX9N+qX1NDOh4hsUgTY0GgfD3p6rrGjk
9twHfQVq6m2pAxdjlt+F4vAmlpSxAFyoh3n1BqmpUYxLruz3HxtLmddNK0toyNDk
z1ty1Jcr+vSOQMKRjREMDChVBNq/7J094HL7KtmOf3y6cM3Xt+JsqoBM2e095JmX
sIJhlRTcDTMM+RWHiKqH+2LVFpuqQgVzuFh1NdvUqh2Uh8OsUNGgYk0jsuvVPJO2
CaITPNAy3k+6wu1J6jLO8v2KRXg1Jh+aUQC2TRBT333FdWhm4shheB9VJfBPFlrK
zXLMOYF4CBnLYVfJKMoQkM0qNCezijNv2RH2uQsSuoSVzWB9cH9UHAO5BFv7+gKd
n1Bo8lRxVX8Y2HK5BPGA7GxVauQ800XBDMgArp0UpmtmikckZeCbU/hgM0dn9KRi
j8HOWgvg+n9nQJMm8LUx3ANkXZn2rXff8QmYP4xoUiS4RJCBKPyKqwjhNIif4PHG
NlcEb7mVH/AuuvjV6vZFmzqPGSvG+SjS0AmugsXXr/U4abRCF6jSXKT4lhtzxVAi
08KDujVaK+NDdcjUH7DnenW+KF+mIoGUboMyyXQVJ/w4YNzeyO7BKUaKurAo6jrp
teDL9bLHY0gPXtdrA4arEXGdzUX964Zrjg9VS/0bpen9AZ8Zz8OwHQNOZ7e7kKsR
k1F9pMQD49eS0OHKFr3NirijDOWQ6eDsaJd+Y7WbY4z+zUkVnxU/AF74ibnC51HS
XrHwm+LIWWIdmryg9g5tlv+5zCSjBqu/L6LSrivZf3h8bzHcH2zzMioUNLKNvVMU
9iQ4JjYPxMakR3AzzNYnIh64p4XzaU71Da9/jsr8uC7wxGWMtUbHIp2ZhvoS5Qru
DqB8EH8PzS7tM5B94+PkcEUg6MqNAoKsCcu3rZXjb2tewHdAZBHo+73/n22tPRE4
7AKzboDkDQZqL6YOUGCtvTmTf6iGozuhwTtBbymFpuRw7ZD4kmScxeVlNfEAcoSg
Y+oCSRHzTOtvusMNzYOSymy6pmYrYSrlLWlnAMoS1YBTdxluImwy8Bs/kwVIuIsR
F6mh7D7GjeSPPJWaHG5yJgm/srx8ca5L03JDy9RBsakwDBdGgxA/U5bZSGo0GC3e
hX/9j43uah/zbtYr4xP6HR5q11JLEqmmIhfUZAezZty3KFh3KP+lF78Cjhq/ibKo
g2L2BHYGl51Tgw0/+pokqaKj76WbDamU3AxWoNC/Hs33RNqKkUQa2q+isRufogas
BgF86CsM9bLSBShLkkIzuChvbmjehbeKzZpL6/rwITExABEwFlLcSmJtCXoIEAkp
SYWrTXMZ7F7Xe3LWlTnh0EKRTd+kebxETw4MmMe4Yfz2qHLf0wlkc9cFy2F2V7DR
V+KY/jsN+411/RdwvtRx+C2R5Ynpd9UzNjmWPTzmDrshNTmSzgTypb7BVyJDlChX
Me2IWG/mNFqI9tN2GcNlPtpFs7uvS+9uqf35vJPOS+mecyzf45VeNwlSR67z87Q0
56tFb6qfnPdqqAj9ds2/6wnIndipPNNBpuJj1pqBbQKz6z/rn9tJt7COrl8VTxt7
7Dcjz9P+r0dGgQXtIzXp6gXo0169FjYZBiFOrBi9BIpPR1A1Qw0zixgtzS5G0E1b
J7qbToccrYI7uuAEF27Y3nH3PYwYcLWjTDjdfTB9XGim0TNduyCKLdRYSvQHy9Bu
ckeRvm5dyud181sl+dycO3FlbbO3XP8kBODLj4SimpSZa5hnxlzq31fiIwU6+Z2z
jprDlhdN1XUYsOFdjPPE7wa2TQQKEMI9lLCGLa1WRYQApF77euwVoaorxHWgH6bG
p6sskqV07NJnq7HL0lEmsfBT1uBFbQfpV7nhC9e7stitS7q4Z9Xw08iTuBVt2jwP
+1BsAsp1pcw2jW+hVe61emQmq3YarqEc1i641JnGSFVxUtdVHSDgm24BIpSKYBaR
ZPeeiSQQKsP0Yl5N3KHCvyPi8Si9M1WWFeLKjKWf/fbERxzYiTHktmp0BNRIQnVj
KYVQO08COQ3Saurqq3+lss2aQ58zuSkSy1WGKy/WPB97+fRnqJj8nHfsdutmV+/l
4764cgIEZKvQNDSt5B/o8A7nocYHMs9v5np16LXlQu1dmykDv54ND9a3q+VrqR1s
vK7MERZkSfGAb/HBUubDvXyAHwL0lCvT1rDyS58LhS3Ox2UCZGOW87OzArCKKPsc
lDSmBRoskGiy2ratOpSQ3qXtFkrSEF5UvsOH18ffW6HOY0Pw5uUT9B1HGND7k/ki
Z0xAB0L/Iyy4Xhx3UxTh5KJ04t0qAx+YiiQol5ixgSMhOeUf73XrchWP/C3AM7Md
LCI2q0NnFCpUyoRw5nfnZHaI78GY5RpMdDGWwymnKPw2Spqx96Pjn5ZvLN78x6LG
bN/v7w/0c8I1gtKKmd+fN5NulJK9vqSXnTTYeT9+yn8DJVy8H7/1QSQGwuABk+T8
AwdO78Omsbfaj0/Kb0Qvvhjj+LNUcuF2abnfUwoY6+GejvHh8meJsEyRi1SI0iJC
uxXLiW1IFCPDjtLm/tnZv6yCcmoRGDo2rFI8qPXTtNPISN5hRMdcddeDSa29/ouq
9tZ3teQa7qnpJu/1N2BQJjXiYFHg+RENqh+JeFSL1q6RA92UBsLzmC/xDe2JkCGi
nfVUW1k0zY2is9S6MKLOoOG0m6qOaNolsk+qDt7VB6zT79/CIe01lhWWf9WiWBz1
538DxoniakKneeLvBUxt+aTueIZPvgsF2DSQFbVCKbn+5G+DLrShqA61AO2nI7mV
rNytHtBN77EqvW8v8s05py38dZu4oKFS/8MQak2kodVaERhTaGDqth2/64/Ufuny
jArazyR83+pw1Eibui3qAKgzDkGTM44torZzU0nIQbmVa0SUgGZAvUfNthWdSKnA
xNgnswRvQD18s9f6aRrM5QMReWUY/OxcE0Ibdio45xr+kQgATnI4HLulGDPhc/8G
D0pA/ddoKbjPJpeNdFMStxToalX+z1XHbRyHmLd4eE4oahJqyhFS02O9TuVGNShB
hhYk2E3nMbUR3oTIwaLA1wGU7pPTVnfuGl7r7Y4v6huG+J80rLKmhQpOFgiTFxfC
0P8Y0X8kESvlWeVIvJCync9agU8eICgTVLG3aHLVBGCmStBMWTI1hve2n+Ftos2z
R41/9y/i5WyeV3OhUXo6S4Yr4WM9ciCpVR3eqgLTe9t34H72MJKpI4vYik38LOiZ
WLH4AXwUqmEdSyCSfa6b94ITysTNGzlZdLeYljNz0rQTi8NoNJYHXbiGGGIoDbIT
WtGgx7jVaEpU06ebvbnhHxRLN/WJ2gDdAu9fIC+gXyXJPUNHdPsi8eSF4khYUl0k
uNYiMHsK9if9bxD/4CUfQON50J71kxvqDtFOPFdhieRr8aO40m31bgHWJWAGtnrG
3mv0nn/eNCG7Zk/4vUbuwqLZHCvQLFsCm7W0XY4aNbGm5coAD8dR4ybuoWB5J34K
FPCVC905fuiylgfzQyUMG8whHTytautsAj5p+odwjCczYOh7tQuCIeB8RphXC8fi
D8oc1aUtawBoxRP6AU0BaChx/N/bfhBVhXPezWSBKQ1M3fK6yjKXbdkoJUsve9o7
dPZcwEyV/FA1diB1L+idJFN0XDdIibsNKiWYmtsjXVuqZFqptYjmKG29NCucm7Kj
iZYl4bPuB68pn63dONDsDl6QLiJ+SCPpXgNgNcI6wmnw/rn1O+NQJj1VwKFiIYcH
tUoPEbfHj38BY40wZJC4MrWGGBNZ5MtsVaISAptD5svKVrWBOj1Zs69MupPhBpZf
EPLnyMx6XKbbE3cDdXXkq23ZOEsGjafzwLyOpbeq47kiGSYCtKuKeaT+QdJf/pk0
uN042cAT9CtWFA/toSRtTm/hMUzKvzg6GJQN0BvByeXeHiM+qA/TEHXfSJRBRsIu
pvdqg97DNemHl9lcQxiE3kraTA8VyRvT3XhDdmJJLSahOBoUP+INh0a/R022gAjw
Ckc2UGmPyfjQv9YRJT+8iP72Jk9huCuXddlWcQXFWM1M4LwoLgCeZWjuSXqmwuEU
nu8BcT47Lb67bLJUmyApWsJCwT7spe5ZXcSMhWF3xK3FVpoxqKWSlNWztYzHNZEK
V1CkDvC/i8i+gSHiQmsHXaQ5+WktYxw+Az6xFqadN9nXU4pvAv2/W01rBWjtSFh+
pkVnTQTBHLH22Iw7xWpcj5dnJVBlWRIxd4Ve3YeQaEp4ReZkj4qRDmGGd267r8Cp
SxxW8xghm7RoobKzJ78ofeKY4yqT4ADViAR7UmTZSV7docIEm5pHAw2GPTUSI4Pa
+O0h1zt+MWWnhxI8RgQObChGm7k2qO/GbyOpklew8+PfKRR3NxyYfxC4x4zkGzRz
Smm1C5evj51ZszhdtprGSisV3gZSt2oNyatDWVJEIRUw8OcZmddfj9dcwlYEtlVq
KnMyaxSYxqMKGp+GH55vAzBYqzs7UmBR4p9iKiwSE8iAnkDamyiakdeykRogxgAP
/LhTCBapVvuQW6mWhFfT+OITLREjy8Q5MFmR5KAqGNG+yLZN/uPAY9VOcu16ab78
SCTUzY9C3qv/XOkg/tGez7uYli5BS+vmVBJL2YByiUw4sqXK1libGIjPUv06mbm9
Ta54AaBbpC6+l+Ih0Bw4lRT3L+r6hzpz86o34o6Jvm6GxNnYBkuicQdykoUR31N3
a2hyFGKviTEdQjju3RHgshNPNPF4ZWCTFgFubGVEFPQrVzdTXOSzat1riEsvW2Gx
FpMuv8RMlIw7cbryFM+eMercXfZp35IFfayfuHE4m49KzaUE7ywM7eF2X8p6jsIO
EQjJoiVKaMsVNNS8OOrXjP/jLq8K/lyoTU/9iuhmGKzJAV9+vVe8mY2IW5TQyVhK
C8XRzGriUpTKOzzJSXGHcLxzkVNlnLA2y/63ldiB/FcQAWBicVxkP5HxFbENxjVs
oB4eu5hmO/aSgIw71pUwqXKqV+rLudGDKMtU1RSxnhT54MFQNncTZVoN37NyUr9h
U+emb3obxk/Y8tmdTz99g762r6cEbm6cJGqhxEPH8HZBOHog8G9ZoUT1+uECO9YA
CLy8VCZ04g+gGHOm20mgm3tnOm/bkPKxmraSxHVD+lpZSFWxcSloo4QnA5BzEa8u
Pp48xC5oc5A0YdK6jrVhYHjo1jDYXyNIXZTES8ECMTcnbt6/n9t15cz0EULoDxo2
3g1K/B/kJC8oCT2A0HGSu9V6bKrRu5PdHf8cnaqvi5Dw73BobSqb2vLZSY+t3MOK
bdT5s8v/CPY0b7MhtbOr1z8P72f433GzXL3eZ/IWI/kwYOiMjx9KKAkXO7aXnfKf
DJrvBy/CW+d4TO8TBKsm+Zj53zedz4fbVy066wUXIOZQMPPX560MVge1bD7rzUtC
XL/sOfeLwmhSlyR+bxvFUMQYPcQMOrDw6sNkm4Jc0qJuqBIeBQKgwoqFL2UePRNz
ilIii8qZRQ8n74hi5EUCkdG48T7AExi4mQo0jkRfvQAPJKLyU0a0IxXzvcRQUE5o
cr6cV5NP8M62n+53WQa7P5N/rXuOZ72Ply+XCKncG1S7xxEYYPOMVOYITqqePdQ/
jpClsZnnEuLN1aasoD77d8eOo4uPOqRSdZyoaM+4detnaf1KQZPuGRtaFMYIw8GM
GguTm3sX0KoEyVQdy9KIYgfOeJVCNMxhWRk6YUMTRELF5bdRIPYkcrGb+dRz/JTj
6dPIEQeha/SuSMysReqC8GQwy+9fuja9lu3jO7Fz+AP82XTxeD+n8d0gLS2Idki7
18xNKPlypr1EvC3ikTxjC9cWASVL3Y0iENjKFlXl3qAjwtVp7eYVI5498Ai4ubJE
jPFP9jzMvGaVNzi04Oq2CwD/X9dZPIQmZzWPFueZhYFb7eGc9NanI0lya3xC/sp5
3IMOOb9R+K/TOk0JyyVbOR0uh+C/ckbkpT35ztGQ0GCvr/k3YhSg3l2br3b9HP+z
hKytg1GGHxQETjkAzjEZVcbNiXCJN8vZFezTMRHpQkzdjY9D1E71D7nspMs4uzhR
1N6WhxF4wmvc3NNUN7f5LxGAQ6qBoKEoOgHESSb7+j8uEOs7Q4y7wz39ReFlJZ9o
BmlABQd2FE0a+GWcWYv9XwDwORsgVF3Y2fBm6KjKzu1znML8xPmlf7H8a2bNzwuZ
VzYNaK6GHs2G2HniZfjx3iDpMQsrtJHmW86f15D7ac79onitxSVtWV0Ib9+TBB1m
Mtnkpp/hrRLR5kLNQI8x8T9mSOq8EONoAqEoe8+SUqygadDKCrqN1TfTQRr05B/N
jJO/FRkr436agfQ4KT+k/JPtrXY+2xMxzjdzRa3oE8oMIlBiX/200h/IOckPeQCk
aa7fjzyogR6xYuZdc28DnhlokV16t0BqjcU3sSpA18sBc8F6R7wtrA6G/cGc4cHb
JXKeMfkcNxhhRkCaFn1wzzpQ4n1zxr0qdK+gDXss7Iyz6MIr+xAith7qYqytBZ4v
pegm5LqW8jbNuYjRfio0WsCq/lEeVy21aIwjk3OIpmw+Rgxfcl40zf/hKdh5+jeb
1Wj6nY7wRaAJAigNRCUc7irWyI0Dj/hKMp1GZF+1Mv1LE2W+OQHpykW7OP2t4Dd2
ZEKnzvWoCxnH0y24M+RJP0Et3vPpODwnojxnLlVxC4kUjMN+aa3NTiLyn+jGAwlO
ZBoU+ShLbyS2cPPcZBBkZ12tWbqbycoN8Lne0rLuv0fv9ali60zJfuW63NpgpgW+
U7q+vvdXbnPrtP1LmZechYzeMl6+zX+kCyLB/RhZCsjFZr5gYbx1a/O9s8vIhG69
wo7WFKL18EBGq6Bv+FXpXmAhPy6dZYvaqj39YIAuh/a8I7ktQqtVLiLQLL7T3TJi
oi3p7Jtz6P1jJmjbMQA0Qu0cJvShryBLLyUBmOr7IbTvJHOj9TWmyDLU5//I7OA8
SAX1s14IAALIasTMy0Md1aTjKDSa9CCXWWVl1rXIcRI/njTyiaShAl5ePA3j1hnD
yKiLN0TzQ6bcEHgET4PP+CRfMCXUi/2MQ3+41nQ7psYGNTF3uKKyf1uQNFW7dPN/
vhcnovwVzOEFkcx3v5tuF3UFo66SRIGkOtbnM+nB8LQrEsYrm3gvYG30sL7oP6vc
euyFgdkB9evGarycAlimXymEDkdb0Qltl0YSuv54cq2z8Qo/0Bf6JjSrhNnOsuM+
CcCBPvXeb5vllf3SWAhF5GY6SzvlBnmNYhHZh0eXe61VUDDnMz+iekLNSRX6jh4y
kCdQJILjHNY7qrLjVPoFIRNmx5KCkqYXBWousv0c2Seiy4VgdLZMJekD13dQN+8s
ktNFu7wjAYeloWK8cEADBEjmPYtDCc/u+cZD19BR50sBMb4ajpuCShD6eD2vHf7X
XWhNNBkuRmPZfMzJqcgwY/AQd8wJQ5NSsL/J97rgPVvVRtCgI+K3nfhdkphohhYc
XVzYDhPqCTylrRk8MHNWgDbkofoM+ae46jycT+pev2ZS/UN9blhMAVyBpMApjCaz
ARaTbLCrqW0TjO8rv9pBQbAPJDMaUn09aEqj00wKMbFML4DCIziRUaR9IAGiLFOu
WnxZt9pG/zvtGBPgUpVJs3rzdFS1eWo1EL+BQKUcxXrTWVMmPZ8sV7I56UJg/pqn
kfdESBzyJBpUm510RFF0ZNi4djQFh72N3ru6VuFK/r3FBxDC52tibQMgpLcyG9gI
jJDx5+jaHeAMYxD6+WUZbRST1YvlwKEqowGf9HRuQ2Lk5HTKTkMcQ6YeLr5aYSw9
xakViI8RD/tUlkWowXvsKiXvfOM80e/CaEBtfMFEQv7jMVDdTY9jZthZkD30RA84
iKM9//x/mr4l9BlH7ETmtRe/6bkfWqncwrcUibRSYzTbpg8VxRIYG6unb2YlN3G9
GO2yf+yMeDKpCYNx39OydF0QEkB5+a+rOmGzePRpV5ki5Kr/SsF4k6I3wfyIwJM+
xrOVMGTuRweYvdjM/2eaeMR+3L2+jbOo56nLelwul+Y0siarkm7mkFBjP/xMqyYZ
JuWs09dRZLcMQ5DXjpeUXaAy/jgvB+HrpvP5E/kaq1b+kFEyS6zY/3GtbC8NMMp6
uh59HDyHmf7pxa3i77ZR3gFTKamPidoOkwtHSljFMl6ORhSQH/59BQBzeZsJ7Rg9
oQun0UXnID2ODaudSo0iaTYDfql7hjTDxlJvLAtbxOTFggEEZ8JFG4eN0DKyfScX
psk+2j53OyIrk1NDcAddQnjTzmov3WI63VKwAQP8Z6zpI4zMVgiJj0A89ZeKhUzN
BtvIZcZMXx9R0DsfNxvYdaUm8OxvbdM6YQFFDrKSV2BQb56DlX3UsT4HBnR3jJ+o
Q/4itZpccT0H7pfqrRcHIHHCXdos0CRqV68qtcTOcvxEPkaXDjUI/rIy1Vb1LElK
qKF+44ffrxV5aUBOg/9PcZ0l5CB2e8RC7LcwMYY1oPc26hei2mt86YwSj5I4svOx
jCOJC+GNvK9jnG/XK9JiInwHSdNOr7Mp+Iipx3iYv8wbYmO35pFE6H4RQDaCoCzX
/USrjfUFoCqdNa38E0dss0V134xjWjsUxVscZgV/oQFW2ciPiFzTLuJdzUK3ZQkt
vznOMd0hWB1WMkqVvK+O254czP/KrvMGKHMF4oHeJRfEsdO/c2vmt7V8UzdWfpJJ
F6U8LYZZqJlPGy1j4Ui4vsAHtQZrBmCW3WdVfg7ADHV0s9beD50+nwr2glMqu1o7
4oVAQna66aleWYvZ8PA8a1SWHlvnk8h8B5EvM4hklGs0k26/oOE6bzT9+B+wc1XC
Qpm86hc6PBvUO6qAt1KE/4soNrDUwGm4kuVV9Apf1THTfrmWazYQtWtes9Gd0YDg
he0/WAD999XdQ93x9kNMjRjnROqFq+C7L5R+8cEyiKkg9ybTz8ymbvP1HP5sxCUZ
eLX7+YpERNtdksbOTWgaSXyKI4TOHMBjA4PbwRrKjnx9g0z2Ub0R5Lj7hCSKOBqe
Bi43fhFUuHYzw1wpLRhjnEtEarQ3MdSsT1I56OxOP0xlTtWAwx5BVleobwFK/8mX
c0a65l8shXwVJPHzyG1D5QZeNA/BPRrxYTA+/iS0qbfThoMj0RciOV199v/uZPQb
/0eWJLFU1XMGLM0ZeGaRoASUhn0CtgslsTBelQXNTFxcpiiKewi3KFhBWkx8/7MH
NXmYZQQI1PWSWKzLdd15K3IHgxZJ/qW/qV5M+HrvhV575pE0ivO+ilEXQ4TV5LUu
G+zBLseAVAeKK/JV9OXcK7M3c9sQ4s3Fy/fusjhqYYcFJ0/25N0hZ/5tcz7ZldEd
dIwMGidaw+dR7SmrrJYZGbctjTIc5oSYbsNZAQ0mK/WKMOeM6IpNUutMLw2c/FN8
IH0+FGUjr6DSVtk0IUtAp6m87MOyXpsU0FviVbriPYOadl4uiNioZON8Ng/FJnP/
CLWze3NvajdvoCderVzN0GYOhAfruxoSVq6zQvScJIRHSwktDatHUg3L7vZSCS23
QOH48KJF6kgZNMSuFxwpvJEcQvel/QfZqocIgntg2DRCboR/tPEjO+41Oxohs9z4
ZvTCMrazYjbmQqLqFQZyN94+qhz8nwn64Eiz6gqITRFALD9H2sUSzOO+f2ZzU6dU
UjzGkO2aqjfyMR/CMgO4Ma1Y1nqzJuXuj44CUqvyLQ2yFwq9xKTSZXYDtRUKM/Oa
90CGGUp9RoQ0M0Z/K2vmL6ucTJ91myo5NU7S+lE4nTK3qyE64gu0j20MkIzcNXPl
dpbvn/6rUzFuByCUaPhbPHf2OCt/12LdcXItQvlSCeXzuscy3S+LTdrHJ8pCFKkU
LNn/Tf3RAZxVIzfZ4LA96Gw+pbW9hOBkyr0XgbAZjpXuQcKslV1kjEPvVgwg/uXI
IMXXP1LZjO6yGwol5kxv9rVUjZ0fwgWewf3fvOdHJBrm7kyua7F425+3Vq3k7jGp
Y9m/six4+ze6ODgzaFGEJ5dclIK+dhbmw6qV8j+Pz0jXr5S2O4fOGTjH5GoEHKNt
dnI4LGQ/b4IPoEnIYKGbIh7ly3HoDsviZt9+3/WGEk6HQ3JdbCOMFpOB6agiZoA8
N6zSciLb2Vny/m++4kGai6NtM755LCF5fuOrfDrXWKVULZK4DDTo2vBABly+RTXr
Vf9lxpKprKVdqJSGEiOyqIGXE29VXqbNVO4taH9JRwJNIwu8+iIx2PgXnyxd6v/u
ZmIzhQgtIeh4YjWGhd53sMvQwpEazJqKsrUbieGwM5qneyGKcwCoaFzkA86gPGln
dtI1xgq4BeZP0WjHkFr4+pqyWzsXRRjJC0JM1f0P3DWoYblOGinABvJ8kE6XpG2h
B39I3t/ZqDT/6f+qs+Q+cailCb6uTM7F/dB9yoGaXAndHv2YP/VWMuSD3BupvT3W
Da0du2bvfovKjyuqFSn02H5BWSpxLx8vi3vcCWCsd5ltIL7gCM4hf4ExNHoJVkK4
3qLPQf+t2gWrEv5Kch0lsMMAfDk/kmmGjei0e1ufI3MgERdXwB87TWr2YIhd8QM9
hd+k+d1IAm/yEYp6CAbZJIm0MQM30GgA37YOJMr7xazxbWKE+Po2SMZorVxBA/jF
41yd2zDuQOubXeYlIoRMol6FHmM2CogS1jgohCgNxg6xfKkOJnAwKSDFW3Xiblr1
axjkCOobP74XeaJqeQG1a8cN115MpD4PCVlIWK9iIPHy2g/3GcfeKmkZfajusrBA
KzB6AS2gJjfnvMoBbqVsvK5ld1I8/o1Vlj7noTNEdBm2XkeyWYtyjD8mE2u1jgoU
lP4u36ECEEwz5oYNgczM0GaV560bwlsZSWRv/QtuoYs5yC4VUk7U3hQfxL18/4C3
FMpT+fdr7y5e4dEJNinaDfkNhgfWAmWyQTQhTRE617lNNag48Zvf+wDnyq7j9POo
jbHQQ4u+6Bd/MiYzakFr6ijJp0Y8GhtYbqi9e97ttHdhCTyuVTbewifDU1EUTAGh
76OrfuuHK6rggN0XP7T4bSVFcUjXDW0mIrIrP6Y+n//4+4DWyaI+5/lNuzGy+exN
c1i8JAamNOKk7ZvuG4Beme9OjIb97QkZ+rPBfNFSvpMLZjeuyDoZNZ+pq8oM37O1
gvv0bpgT37RKTsvrsZa9194EQFIAWEohjCpyk00KfAYE9ZIEqg1MRPeJRy82ZmhN
SXAe7qSWbpMwvXaWIttAZSguq0zDBg1GbczGzUrUpRiDzC0s4hXTLb2mG8wwB4Pe
BaJPMWoZDkgkd+ajLv1Um8JAJa1PoViDkrSibrO3+dU5Eoq3o7SsWX+cjTDzSqG5
XgRb3Y3/M9GbkI7DYk9eiklsgMvEgQj6s8M060Z5yKCpWBJW80kT2v9FDIRaBs/2
yDcZL2evQoztBF3mHMEpSF0GQmcu8CFkL8HLAmS/gQ+9vmRIdQSSkpPNbsu6fh8/
eXTPoM9qPbsnEcbEB1eN1OHSWCSF7agpAdtPhRXYMCi+U2dTBltDYUhi17S2JRMj
mkVLeZlDedcNO5sUkCJc8OSCIddip51sXZUkyzA8adwqtSkLQcGFUc9/5ID7wVGb
cd+fXaea1LhJ7GqUop3tlX1rqdUO3rMyduMkPlbWS4JnIWMgZ+afwg8ZdyeT/Afe
XZB2FU7PNaEM5bLkF36snhQSth4lKaXUJsvHvAJszvTssFdsGoY3aC0EqVwbiPk3
hU8mzPZOP/+Ts/t5ZEJHDX1rvFDyIRGULCJ0dFTOomjqeylzGMJLJ0dlIS3BKaFL
3CoSyjO0Q3NDohV1160MHvTsE5mbzVRD3NjolF3xcidSc6h7SVctRI4ndNSQoLut
8vLOsE57IrguXlk9Yv65i/O2N+x9epLrkdeLQnYkM4edTenGNsBZL6UV9GOeQJfe
rBWPUjJ+oNhk81nnXkVHFRok8KUVzWsSZKW+OKjUZaqxzbsaw7SlX4Y+dgaStUBG
UXCIRBurydoJ2glv8ZnGVN+vUIaozf4z7ATo6iwdUrI4rVajCQMocHxC+zYckmG/
8DthaMMmqnchtross2a2HqBZTv8yiVoxwpbhvq7RrTSBROY+eKTk4uiFS75agLfn
qSo2FsymMHePbNd7DHibpZ0jH5pNpN/u69osJxabpSfe3my66JLEt8K6NeAWGrx+
5zgMhNC5rmnkbHkrJI3ixS38BvpQ0K87tCAa8SzgygN6SJn87JxMreSw1r4g8W1V
nUkBz4OCjFmPwWnaxsubjrMw5itKOn9PDi5/6/ZrkdICcbA1LRcvQbeQVJj8pYr+
NgsKW0kbJscsqgZncrSBKTZc6j4BlEXSX8yY3RAHPeUj3bF0H+9jHYLbUwCNpAY4
e9PgyParbNvyEUKb8BAmWjKJ/3aaksV/VnQJKGhuL5LSHIrx0/bGOaqPkQpR+Xqw
ROpLXgP+zJTT+6DZTNwLuCZzLkIpTLHk8YsJi5gvsw+FBWYO5ZD6kxWJh/Dn9oOf
sTq8oX1BHQEzYT2hB+9rad0dlYDo5N/ogQmXLKS20p8ULHK4q575IBALhYoJfV8c
uyNkoXGjChCYrsamJTow26q8hpEsJ1nMzKm2LaiMjGy/LfVD6aqvI3d7/GWgMv06
jPiHijt/WU6q7OK5D+/uN22CqnWfEAeSv/7pTJ2meNTiV5bV9pxYe7d9r0nzKPdW
PqtoQ9fOQnQip26FACTAH3afhryoKZxVv1s98fKYl4sI207ACdFeJX7iNav1fZEx
6/dYu1+bc6JA/tT8w6uJjyRnLY0iZl0lWerAgQXAJA94ODI7g7kWKAletohoSDjO
5APf6UzQwG2GjH3OhpCcyhw4gUhrzpWnlEa2HZp1qI3e1bnZh9lTJC+tpJ9Eu/vI
xoDjOSNOhXZ5tjUfJBb9jJs+Y9NzLYdUh/vJFXTaeGwUOpjtvM09oPtFZlhz41OW
RLUGvBm7gFfOcsjIC3izHzW0cfnobjbbXJPKZE/IiS6a6e4Mz6LqvA6MubqCmyTe
Q6ePulQ03tmfRO3iOhtjPtClHTVxP9dyKt3pBQ0FW48E2JEbZlevUnsR8bI9n5GI
pjd+l9KS6cdG7JZYlY2UYgLYZKKp6fW8FXv6EWkwXtddJ2h07ZjqkVMjw9fq/hqs
MbhhvD6nzCKtFTT6feHZH68Yy+zfzycajY+AwWN9ZVHYB6R8v7a+VOavJdqCRiv4
KqAP5t2D8zm9iPpLAQtGDgtrNU2dmjgX9ud2LK0NabrtS5qVNCuZeieLiTbjAA6V
PHbntOPOICthEdzkPpjqvvE5fXJeV7qRNocjEjWGy+cksQ48wTRax5ZGwRqJVIV4
Vn7K/d+Uq72OtQHbge74bI8R/7pM5Gm9JpcdFy6CR7yGgRpJgvbhzjNhjcj+E+VB
WIDKmfBplPGsYleoLf3S3a2pGlq7S3YcVnmYTDgApNwBV94f4UR7rE1caZLJ/h4N
/xJjEQJ4GUyhWXmPLgzgwaR5GKV6jMDCfLp5qRjGN9FapCbs1m+4U0EKWWlsebTp
/uEhFEyxVa6+jr/a4zPyFE4ueIRASPRnAEIbyAgjmqk+e6IYScriPkiIAZRPo+KI
ZrEv9OB5jdB2kLhnGmo7eLTouAUNLMCkyoEctaYZT0mHmzGF9KRu91oTZHYB291j
yED27/Mj+5SvwMgwUxT5hmmu40rEUSOzToSvvcxbDALpIg1p/EJ0T5wKmFHFBnc0
Nm9qP1Rk58yBFq4uaHnJXq0tvLdaQ8mAYF1lBgmkMNz7BRC21ItIoyXJMmxKQFmL
FSzNsRdkT9fDP/PTBm8uWIYYjpAXFH2VnXvjn+sQBChLv/X67fHSARWcoufpbu/b
zY1Pd1i/3gkP5HMB+UlAN+dmq59SfrItsL+Ys0v4a4/JpMYNELJD/wMy9PFsh9Bq
H/ymjGDlkDIUvrB2zGdjK8391pNzJAfz2UkP+RcpIXIk2JgdLFfjYsCG8SsY4TN5
eQbebXV0oU0y9pUouvh/9tO8hJgAqsuPQ6MZ1mBbjy+WhnTpGdg9T4HHkHyP79es
lDdW5UudYhfVgM8RmnHi416dPpYIJrP9gz98zp+LTq+sRP348JY5tj5V2HFmsYTu
7Jc/uhzA/sun8vZApj4w7oARF/+zAeEWLRs2pPOlW3sO4LiO0h3i22QRmeoceQgS
h5k9f/k+pogqptEtm7MOuClQuuYpuSQl+8rcCljKEfZYpFQ6fLjTOUqwEsNIa03J
ExVWHwNDQu7yhrhyUL6QTr+hvrV8d0Gn5h3Bb299eddg7W9/ZK5TZ4I/AhCVMrpe
APLskgw30fcIuV9g948QBx6PpDZEYso46jrG+c7Xt0LpV/byU5/wEpoBFTkop3zT
r4xUXQZ7zRMy/cJmmZ4xJNoDoUCrW7e4/fetGXGRM2be+P0y6md0A66uDVm7dqat
t5zYmbqCUVc0GsbgZOuFbemgrrKA1qI45+66OLGVw9283SxQlmaAP4PpyNFQ1Y5x
b+FSM98VFjbmSez+r187APkIxJOtU1wqC9c9MI1F9R/ylOevaBSvLcW2JupAoC4n
4/6mQWvnUW5IYHdpXVwrc7pnYjz9pi9IedsslYlZDNrl2m0AEm0ZoW+4ueWP/6VO
SWXWgrk2pRIpUbL+14lI+CuepkYPsLzJnY7tBkAW4/U06lpO73RCngBGFe1wLqiv
o7B4LPlPRgY3aFTSeofsn2ayDkVr6gIkbpFLyEZNsglH54z+bLThCMuZ4abC/Zat
rq49y1WPTIb+sHBVsf+EcfV7/cBJ6i9uj6d2KYi5gMayU5s2NWsjGnHgSqi94uNG
XcBNCF2m0/lGimIv3XKdoKHt2xpkRt+ZuJ866AqSzm0BJ84heGHhFXE45k0+B6ZX
dw52L3KLkBMIEnCnxjYa8UHbmKat6/xu1JNR3CBdboEq/aTsHfazHARD1B/hrHqu
e81CcCAOCtfYlnzSRMx4AMMsE2gmcmkG2R15lLLPjNOcQDk8VydbGfPM5cCERtD6
/IRoU125JTVf1H4NNfYPBA3cE0vI5ZU/askB5Ng9RYbREU9aWdIvyR/ZIBLA96RA
BZgAq/ESmO4Ct5FuSdov4BDMLmhbYhwkwGd21lF/mcmzd1XzdNDpc0bdQETOf6l0
26tyG9/n1Iff7+wgwuy125eoljuhTP7/ZNLCduU0DfV22iODftfSWvvg/Y1PmRH6
14L715zpbAjz/MK1VeGNbY1VCkw7p8PWd0GLaGAO4lhRDEOD6jjV4LlhD5n0+Vaj
Tv4dc2R/vytcsYeeoU8XgY2vNuQU0HmyQ44Dgz0woNP1xxjZTiV9fG0jHixwLnZ2
P2IO7SL4tutESYggqbmIllxoaHih95nSSNqzWTtt2GgVaDK0KZ0LyOFTwpwTLliz
k2vGn8sMa96k6ayhpzi/YB4WqUJxSCV+WOvOPge3gbBQolTcA7an4JR8zJOWsBZN
lO8xylBIZYr1sDbY/KySwkQsCihdfYZ6DBKy76CTOJLRCA2h1/5E46Qs7WAgx4cI
wRUuWM1TFYA80A+X1zcd6XzrA0iCNWGbmf7ke1xNaCW3fGhuhXUD6wjJ1Ky46w33
JlKvksP/thCThqNKpKoP0OlUFC3I0zw80PzAlyppJELOcofdG/H+1UbpMMceguSl
WbBUqxtKLdN5Df0OMf8ViUZ5STLZCZCpmB+kBrZH/vkv5+KfYhW9sN0K2xCzgh0N
mvQmqmbB/LHswFLvTWRNFtAEmB29ufBOe9xMWWqSdqhNfllBCiaJ1ZNkJ7M9nHHT
GKWqdpqE3a3bSwX3DhOy8iTSFciChEzDyIo2yVw3uAGJqSIdRkQkzwET90y7qj1K
P4TIoHx2zLIR45WCFqWf4suNpYPaDIWjUtB/Wu9guIS9eg3Y8h9pnGQp9K0ZaYq+
3pDRQyTEcB596J2NQsIOatuQAw4QDZwffsCePDByKRJtUDsAb2xPIy9eZlFBeoKC
ZLlq0ixpGyW/P9OPZB8IZ8+p7YvLWToylCQIKd+LR2UvmNRpAumjLpA1WAu7hEP5
FpYDm0Di9GRyjB56+U4lerzeTb9Gzg9tzIy71n1nhsysB6kFj3hNdx1X/+ua5UyC
ZHiQkW4ElsykNqfJSHP7urRmRWnn7A65awosXpG8uwhQ9wUh4Og1kkRR1iM3ySt4
BezsvcTO4CHQuWTlBxnl62xcez1iGeKcpkM4DF6/H8wAGQNl6zC/kr3BX6LmS/86
cSbrs34jTmgff6TnmAqCDSuA4e9ywFWIyFkd6vLkH/8GnMCFDi8WUHER3oOpQow+
bbAczOPVfs5tODP2S2pzdD+T2vkKIZ8ldeVt9yKCwIamUUrExjbehsHX2MRn6v93
n5zibgfyFNjRkxE9RmrFT6jWrSmdBKhs+U1zTPY1iuxMe5KNI/4UgHecUB83bGfb
cTK49u8Oibe5rDN44Zk4Zws58WWbs+8cWaRdiRZfy9T52CMKSXvU1ceilYcz6c+w
EVPaL34VxZF6MJkMo8LIriwvDbg1rFS4yFdabpAP5wj+TDl+LVSckRtnAPXXs1ap
TY/KXICnRSvKvVq3R2qf3TeZxQqjgVvHm+fKOW9dZ/qPtpqzNErQqh4ETX31o3r9
962EDe4yKV7uZbLX/TJAPkKJOpOfhqZVqi8g5dGkgCX+PjC50k6tJMlcMnxKe+/N
8+5fOcThPVnhePpoXwYGAWJ+20kiKxgYRGlueEM7Iwbvu22f2I/3Y/yBfaa51LzN
V03zSS9K8HK7g7Ik6nAL4So6SveZESow/xXd4/9+olKhpu91bSnLshtx674+66JJ
UuZ36e+vwsyyvWr2kDGhGZDoErjyrj1prxINeExMwchV9nS2JepVRe0XwDtv0nxW
6xa41CnU5I4cCPbgD91P3Ty6GqZ0P9oDLMLqIu4wJ0pVOCHWZC6FeFu4X7aiX+Zq
zrb23ARXgXknjyqIgfWSrTGvGWV3BmPo725SUXOnBAOJRYXIqwHchJHwYMBSUew+
KTewXbx5j7if9c5d7FWSu7yx/lVUxAVV87zudtrcF4B4fDQLcY+qj6LHKkDqpzHB
XbcpLZYEJns5hQkN/f1alM4e8mIMUlCnDyYqiznf+vui3xzHecjvHVSz627G4gSY
TGdMLKEMvglJz5y1fVq/x8PVB6XdOlzP11PW/4DpcusIm/lI4ysKTbvbzhcHXzPw
vxXTMiN+bWcrkv7DZcRvwgb8ZGewjAQ0ce32BzMFzMOQqiYn/t5APrYaxDDEbsQn
F9R61+7cX56a4ZTeZsnn5sIfjuPeKU8YM2YAtt6pn1jH71kgsPBHxTnX2ejLtTVj
+WZ6Rtni5FI3chp4IwSyLng2+cxnz6IFybzOGCgP6U8ZRVGDG7EAkCPNcSV+DXy7
9e9rQEMN8ZhyStbnWyGj7PhLZvnew7S4uTi6umXioeKRzeMB4OiaVqLdoedPpCr0
TbltcIlgK4uO4prAiYdGlPUi7uxZ89ubmLTORQNRzErqrQ3xesIGmAVIo7SezSnt
j50nw4+fwMOk5ubMhre9FvcfsTT2dw/YkpR+MwmrDpE3+PU4+1ROZIiQUg70wWKR
bOZRVphnReLJ/6ssxR6auoEax7UViOuCWlA7+xVz7NFBKJx1RzypnjL0iewBGEjx
qwuNMokDxcsx3Jn9Lu0LtVLYj3Ilp9+pQPDiPOTF0HvFxD4Va8NsFB64GEiJqUdL
vyGFMdr+F/iKNW98nZfsWi2OpMFp/Iroi7Y1h8h9uQYLp6m4SlTWuw30Of4drglV
zUp5nK9/RyavRaNdxCMqCXU/mwHZOP/AYnIf8AIDP32ZN0wadPNZHLaoAhMvfNKm
ckImC9zGU0Qz9nFrWmrFJxbBul2m0aYTLO+8KAcb03D7XnDPg8YR7WVrfnT+Iq40
a6MxPD4QPOmXoM32K23uz9wTuAIlKxCUWf5yNH7aJPxAAfJ/e/GSExGQekWVYGgZ
7y/51Puj1bhKwj/xVdODByQBvg7Wl8lGSrV3GcGbT1oGAEeEFb4hdD9nL4Myz6Jo
lmkdiA7gwi/R14RdMqh6PuJ/HCxY5LgfMI1oTasQAKMfxZlK0183/7SHnCwAzrTX
Tf5BjnMcT3nm4QcJMtQaPubSqUanjHukWytSRzeNr4XNzr6HiJdvfs4KY49c31rV
c5UUDn2+DFLnkgrhU1WXO663lBDe581YbRtoKS3KyRR9Qa9PMMqIubygJoAhDane
zxNnhY320p6yrRXcrITtD+ZWckhfucQWXNKGAl4rxsu6Y2ZVFuhAXjPI6+D+UBsI
rEfM8IeUOxEoxJH9hgK0pte6RjuWsX23timPA3Kga+//X7tYlPr9hgmB9RScr4lP
T3LDIeXTSyw6O/EEM6X5FA3Etqg85LY6MWVtqaYF8s3LdDWueNorzx9zMbsRMwp9
mRuYtAkM6TwmScLQhO6JBsxMFDMYE6oizj/Tudzbn3FUhKMQU12+O51DX9zh7Hqm
/wVuUbm+zTKTbHRIwSnmrHuUlT8goCh7PVx/vLDvPJfQ3/ojuP5u/5G8/+D/XySB
8ge8MRJRIzKmQxcxOqgsSdiolMK4ATA7Uwz+gBkE6yhJal7w+xBEBJ1UaXiT1WLE
6ZWNGXJqSBOa/Hhn6FsfWPwLA471U73x0ePqjwNr2YqD0tvuw3qO7jf4B0vlpIv6
yVv3aM88jp8IpJXJCPjFtFFiS1IBFbJ9fQA5LPQZCTMvX3372xLYlpiH8ZzAtxIl
tjoTV2mISkp93TZrYxpot8T94JhmuQIphuykZMNhZmEMa1dyyGSM0gv2O1YGUVkP
lfuTrwGR4eJqWKwx0LH6MPFh0g5Z0NArYKb4UvkpFIIR1vzueFNzcUstV3sR+x/U
rBZOz8CppGFM2H4hxqw5rtdozaFuHypMlA+GJ/zMXXw/3U62l9z+nLmutvvKQGqs
U/KrV+ggfaDvvSfzHDASP/Etael72Wxkb6ezvy9KFNDC4biR0dh/YcZRr0fL79V4
JQZbObYxR+Yp95VTJOcctOhlREcy/e4uNntslZcQzfDiRJfzQx6u3qZTYwunSP1d
xsVl1CehxCwV6bF2S08lfEZrXhE5BkjkUqwWC1PL96QPG9JSFxnquohJB1r6i92g
jUuLjffaGj1lEObAPUWg7qZRjp1F67SLrOB/wVkTF3mvoMzjHIkQjsSn+bKK1Nfl
vaOIpd+U4lRpZXut3ThbSAHAcI7SIKBliv7+A5oKJB847I7Jns4hh91IOkf4ZhpD
s0UQqAIFKk+GOamV3kJc3P2NqH369R/LoYkYkev/UAl7spOMOnOtk/aHip7S3VoQ
Dsyi1UseCks95kDB9s8bFH30XdnbwKWgWQk8HiwdludnCPdwCvjZKFTW+8i4hwTr
JRDTCIPNNkPQL88xkjzLwSZH42YZjPJMBpjuORXwDKVwaX1FPRlmzdhP9XYqHb4k
Dw26iEspBtcVUn+1egfpvp1yKGBQ8E1uf7qreQhJdwLZb4KKlQGNfV1uZe4dEOwF
exqi68L36mOIagdJiWXR2y6kqi97Q5Nhkr+WMb4DTzp5Q0SjyU07FPwMfJ6EC55C
LeOsct8Fln3NzMnJstD0eE4wPJDjq3gHzLrBOuIJbZVcBjpJuNyeLL8yRRAi5cj7
NTcTNb7o+gHT4r2K8xoYyhy2Nk2waeHpUHbnyv3VT1pNaYPEEwmfWqvQlQRa3uqt
fNZ/CdLLER87m6OraZq6rQLtPQsNU+ifdq2JQcD2g7E5/I9DVsfrUqVHeqHzfY0e
3Q9MPJ0ESrk1gtkSrjpuoOZl4X05suAG0Gd7I81H5xI0zrDDVf7+/6/eqfgWl2uL
yuyFCo3A/Cbjlehmma9RGhym122rasvzjwU2joxxJ/IW/SnIZMpDr2yi8NcC9j7D
Va5xVdmnjdyr0sJ29X32wDyx8sc6UmQHGwJ6cuz/dKRW9yFXAnilyy6LYA2lUO0L
5pmtu6U9jt6EqDEQ4+PGAyGSQJmYSF0LGU2BPoRkZjHFICKF3ad37GXI5735oRrl
I2E9n6slxPMilss2/adoQMN4n4nOf+M3nFNON4CFbRsqeun4N+tl+hnyjXZnQYCk
4VlU+SjIYidkx2NmIAA51FG6UpydXLG41R9v0wiNjxKK7FUE3WVoMnYC/2JdkltZ
NwgOjypFSZhSJKD4jLpm+7QCrLe4SM4JtjXR2XcI7si6Soni8xyZuY8aACIzAy5U
SPNhPr1litasKcG4VWblp1icW8Rxyzr9MBeGaHuRL+7JWwFuoMQkZAJ8A5SLOeuz
nQW7nVMsINjwGzaJLH66Y81ELliqfO2nMFGHzuAYZG67NxPhfm93LpjzZtw73oak
RQ3YTuATiT2CLAkCDqLfERLPmmP9cXHcX1emIEtBpc+wv2c2qzFbVkglm+lhyWWm
/HG1+sHCRJg6uwg89NFCOaOBU9zJ/dmBxWUTnxB2LGVevab4zJS6LBqeIhTbEB1J
mJz2hLeJ/2kzo1n8zSbLKfyzVc2oj+pqKlCHZC/qUx+AIDmvoE8oUaiaStPye0VP
FR3GLhgqP5pkM1ip8iOW4JNhTM0+5ZAOViAwkHTTj0wrdWnLTDsCNVYyyKyMVE8n
cDPtqTUikYWDPx5j2LNNlGDRVfHmQD7WQe//zqCDrEU21c8b/5ClQSFClqZGNQtv
zvdE/TtA7zA5CnXNKp1pZgbWhSlcvSRzZOuPAsjemKeEwFRb2An/geqk56RFhWbw
onR73FD3j1g80sDMvS82EQW6dDHujapVIe8SX++Z4M8R3ODh8/fAzk7BUq5ClgsD
FsSwFhCXFq88QG3lRtXdFAuL9neDQOAFcj8cnpz7tlKZD3Z+aUbI9f5bopvLDfQt
DGDZgCfUI1CL+Vtyulpa72nrtw6i4SpYxvzfPhLMqM0IJd8ciCmph3DAtUYwXhkD
5gr63xcwwsJcRQqg8nMR3och+TVQ+JNc2W8eg1WeHljX0DsicEc9ojA17RrjlOFx
3cEJDSZUI6O1TRFg5L5+eKqAltOlEBt3dAHZpMs7xXMWG3vIpvzpnW7/rX3+9pZu
WjFlLVNKU+7D2hCrsemyHBMM+LBEgoCRFddqQ3HcdtzSfJpkeH0fl09+VzKZsp8f
yuw/9filPmAVyP0OcwKFeWwleJOC753fKV/4yEK5RoW5waA1Vt5XCrYGa+cYrkEX
0nYM/zpD5fKov066NE5lsxR/Hzuic9kdKV7vtAievGaXm7jWu4D3OigokZb6QSPe
Zq8dlbCL6533sGIB7kZ6ikAQBgm0vZINmQ5vTzOUZ7VhXrtDId9PTeuF0nzdqh/X
ZsFhjHaJRB4pjtPazJVBfYGRIRlW+p6Bad/3NHOBbcBo2YqIwaSczG+w7OhF8QK5
9jcobYDU0LD/3KL8oY+N12tJNAP+iP0aVpP+0FCo9aeIOUnhqIoYrrRvnYjv1mt4
QQjQpceXb3+4jaif8uhlBW8INVnSWUNcXyHueJqbi0QBzjg6Z0ld8KpOqXa+CD6k
Q0CfQkFKrTdhOH6fx8vs2I77sVN3GuwMWWGjeLjVJ5746Fx9Vg5mY1LEzVMkpwl2
acs2gN+TBzFmEfyrzkZlCd3Bk2x5ePzOJF9VUNpjhnxQC1FiK91RxRZlhj/8h3n3
MXYEYMGahPY5V2CQkmNcTSqKQm80UKkx0lF32qWRB3q6Ko0l5ueoTKex1CdUUIT5
G5d+KUXmZrsp+H1mbvPXJiyFLXvAKbX86cz+59rlgWS5y0JMai6EhkPVuLG8uhO1
cNrvW9c7Kx4eLznOFg5iKhpVRC2Xx4fdc2fl3QwMAFmSssKc3QB+aQkL/ig3rboD
npiCiH2gsdtXXRcPSJzlQZg92mMmwPiQmw0B3T4MkQqxaDC0yjn3gkuyEtypCKaE
lb2z/RVom/kn7PdXfi5+iRFSjoLqrVju7P4ndJD8QnMhBGRurVCTOU50O0aYM2ta
U/YsVsLBpGgrozKVfQllZQtc82zcOm5kNWFt0qpPwNMQjsKlChbqfW4eoR/7l+Jf
v9tbbjr99I9Sh28DpGaxtNH14zwRNgF5xthxvrOKM8UyHURghAsX/BZ3vFgWn/jF
SPFuJlgHzK8Kdfu9SK1tAPPuI49Cl0mX9GKJ6VXA6NoPBXiEcqLDcnG6BoQRMUCp
+ORhk8l50g2XsCIBGbGry4tvsYBd8DPZSePOupo00OopuZ7cs134Uv0LILoCMTsp
T6KGzeSjI4LNz30yUMkpP8Yxgd2xwYpCC00eePPGhxhpOWWTNf/JQxm2MaD+EBi8
Mrc9+68F7/B0ucA+DRmOAWqHY1ktY1PRFnm4kjpzskfK9Ks6hcZAFCdRWoS+cwMd
PIM8KWPotlG2Uc20Pn0pMSXVgVsuXb5oece4/zLJJqCRpROiDfOa/i/r1i32HjEO
tptXTda8w60zjYxK8Ri4h906mW13x427mqy6AdLJ/9qLop9b9vxo7xl0V/In/Muq
Rs63wu7kjWTJS/uM640qMt6jEok4GSXEnCxam69mM52BcD6ln8iBBQNimevyO9Uh
xv75tqTwVgcnhBdUx4+53l88NKY70QzIdKEvht/uDGbwcTMUZsb0LXpGpppALbWG
M6ejcosdFLI8z3vloSkgdybS8PpdZ88aXH6r7Azs0gASsUWj7S2K4LPQgytREUrv
chJ88rrK0IN2v6zVuFU+uzWN0PRQhlVYLi+osABBHLAiYblrFrinyLjyqYUQHZJ4
rszN81mzyM3hFUSwDfQVeZzc4lpBd/Fqu71tbm+fY9g4xI2Lu+ibb4ox6NNbqHwY
aas7hCJiuRZ8/tl5T63vyZ7bIHNS1cEs9Iy4KylhFnCCYoZymy2btpSGqpdwBpjh
hnXpouMg34ui4sW61Bn6UR4snoqauQHck4ptt1V7WZD/EeDvcGaVYpXhtpab+eCJ
16AO5KluL+ByehM2w9k1pAlML3jJxcNWXqu9qrQImhIUN5F1JD1ikc+DwRIspm1K
0yBHzUxmBkrnTgXYjoxUZ8DDmFXDOfE2pUAL7Ex+UgSUm4jaUcjmHl0CTHFsxUgW
BsHt7O46KxqaPKUo3hM91U2LsXffnOiLG2Z1tylS4aYwRsPcceOhpLIeQe1uIT8Q
t/qEVG+Kf4KaFLOIU8QKHjmuca1QEae4jZB+bR/JeqWKfmSOMygkulJUcKn2xNDI
2j0E1NlECEYq6of6SsHx2nS5vDkC8gTSH9F361aO/ypZpkR24K5uYKzR812hrvQs
zkIv30UF25O02u/c2H+tmhtBgd5zJbF9UlrxSQ8jf0dSbpimGgj2VAmvvu5Qu53T
+3QM4+Kl67bp9u4vCdKhbVzAzHN63Cy+tpsyW5vJtmC1Wo1+uZE85eBSqMrTwdTB
rvNwiNdGGQswnBr1RkMjy9ikKrrBX30C+k/p/tgLnn/OnBBYRwH5ajElvnRq7g/7
a16zxyCh8nFWz5g+RaZ3p82Lj0g0aZ8BmW1x2ItWvO8e7MqyasBoSvZC1QvLVIYk
wJLrDbqTwQsLCfelimR4CKAcQlGx/pbe4EmEID2CYg8t+nxgdgBjetcr256qjEYj
Q2b1ViD3nPoR3oIQGM8HEr6ZtkQQOHlNu07E26ePMeKzXGKqrrf4KtNGYskWi3do
rKSuppvkUFFQ3R9DvnRQGrMhaqjvDuu/CSoyXqRvfH7JZTocWb7J5/a5qs4bWEYl
pcQpkxty/9ZGz9rRjVU8h2FnrkTpJl3faX4/8ApIJbh293Xfho0YNxpaPyWLKOYP
RvG2IKKQqTTjKkAUz5qOTRehYzryx4txH0OMKoRxzxKdKpuFSMM+Nfi170zwQSI8
bGLJo82cFf/Eck1davTSzh84G5gDr09a3O2FUKazxzXE2bgI8JY7tTXt8lH5euqs
cr0hbrZg+2raPy07IPaO5QwYnDfgOl2qSjfUyYPLA58aprGNr1yZhUXUhvySbJTD
W7YyO4Drv/w0HSlBjG5fXUoXNwo2tNKlvZXDXE9M+BpFpnVL8F/L/nGDBZRJ/+qZ
NCAcg85OMNU519YMraTWa+W2TrzdLBECvy/xqoGbbjwIpjat/DHD6DfsW/cfVk5l
VRBIqtvuzr+9tsg7nYyUU04bS6/emHViteLOCZ6UrXIBo0e5uhT80sJAT3Xa/jbq
BLd+a3ucY2HGbPQDnW8Dxu2pRmONAGngZ+rHW02fI+fNcA34gbACJWi487Db830i
ECKc5/Db6B8LT6/CjcZhWtJXmYhCUIjdlTKZZmku6HqWsqJYztag/Y1k/8YLuJRD
9sWXuioVO+JuZ46GnSkjt2fga6XGM2a2gefoQpvAZruT0vL+74NlCXT+bDhpG7My
cqUyiY8lCHekL9u2tvfpDqlZ0g+LPZTBBMWzby0t3HbLkRUY1+joWUFnPcdsGsPG
nU0eEhjUaRjJY8IYLXoq27oUJbjlMjO5AO+h4CO+2c177bhi5K+eiLuQVN2C2kvC
2doebrezktnHMCx0pexmkut+NBQCeqG0A3mq3H4qkeak26j6jQfdGH1m7M6hNUwf
PiZjE0wcBUnEU8uHvhCi05wIcHjZSOTdXmwyFjinYVIQ/6zTsA44+hdz/T1K9Nmy
Ka27rxOMPCOgZ0E2DTUKT8E2yl/ftUIWEbKX2yNnnVq2ICThVqu3i3rMUisjJOha
ut+Zo+TYjlg5P0M6PFfdhGMAfCwpc4dAOrNyMH2BpqLV8Y5XKe1stVkL2cGeNBlp
QdF6diB7e+3RHUcxhPlUWuK5PlQnuq5ckhy7q9jVRp8aiNqIVgDimHhBfT6SaTB5
FyVpN+L36hMi7bWyLXRj7dPZ2xWqQM+WKKxnguiHa4KEvAsJ5VRe+ToKNtt1o8Ga
05a1AFJ6YCCGaACiW0RPHkLD7+X2j36FVi3L1QlDkUD+dX0Lm4WxbxbdrT7q0enb
Z/O9ClKXRRnk7y10mfHXMupWuA1NZbFZG2IV5DsIVlVFHWrd8CekjkASLR22rasl
I3IMxuTVki3MzSSALm3eAiMOZZhvz8v6teMzf0SEcPp+ugeFaKOmnFaInT4mES5k
T9YGxcpxK7bIQ7wHb8UInsJc4jxkH1uHoUO1Q4Gb9csy64CddCZ1+NA/Fl7/cfy5
4zlpL50aL5v20Oix3yyQRrh0LDzsB792FimGu459kh0T/QIzmkTFi5wi23IlWXt4
nODaTK7ganNqiSgzJQd/fkoVvWjmR5nAGSd5GRRwAZQyAEjvq89gTNZ9RK2CwmTX
4PuFXv4/S5w+Hmltb2QBcEx7R1Ft/LVDXsfhNeprdWC812pADtgNk7BHdlH8JxcT
wVepPd2wEiJs33zVMF3oWiNYGvLNxIZo01TiY6smZ33lWMyjWl6kJIl5SOecFksF
HFRUamBOAzE59h4QyCoqrT5M4i3EX3v4nC+NS14H+VQ/Hktzx6PeINzK2UHqgKnz
acUIStMsSN9wISiPMyHBS+r8rXD3bfX4CexWEVnffCyi0OL135MwND8+AshU2EZi
WE5ZQHUgm/F7wU24yd8oojFv7DKBcwR6bPgsvGONK32DsMFtKcJqZCqWd1iq/QYe
v/F/R7z4Puy/mU3Upw//vN8pOBkosKDa3EiQXWrUa6pJSSeRIYR934hKoHLf6IYH
wky7MJVFx9W53hZyJsbcBGzt8w5ps6KY57zIoe9I3j/mwFU4jKsNUAFdPWbgrkAX
mNmV9n/qXUhuvOEh7JG7ef6zV85/QSd7r+6gUFtD8sDX0NCM23chvHQzAsZ5fMiu
InZk3qmgg8kQmGVB5f2O+7EcTwJKRpHQwEn1H8zxnBmJFDWJ0GnSPlJAu4LI+4cT
OTh8u9br0w5zOoQ8LhKkTeMvvGzsYq1LOFvq+S4yLzH6ddeeL+il9/Ywtbb9IX5S
0AprxkCzbBCMAvA5YHZlRwwyKKZPUt0UW7iUB5PSbbzP09H99AnAV1X7aN7St8bc
KiDra6i9akm2kJ6eAE4yskAJ05goZc+kwU4H2vBkHI2J94Gq1YLnBR6JEaHmS4Jd
RmniC9dvd44QFsr2viD6TOv6AgpYITHfUrKlwCzlEscdLUUJapPXqFUl5q2eCvfZ
MdFgwCao/WsUE5DxCMu/oz0Y9sGJLi3JVv9WPN0gj2ZrEpt6EDT0Vvg6vNzvWqD8
eNxoOLOffzWvrAXodBxLFRtctKOaGO6AFCy2GoaCjWEQRppX/VEuP9rAcTsBTpxb
GlKmOoSHGz8b1d+TVOvnBBSoL8Lu+WRTGO4ElvDO93hoF/WIk2J90OHrPqO3+BnK
J5+iLJVlMKyXDqWTJ+oxvHLuPtoFs5LMFZoFSZSXHvyYxpCwZ4Rr9UBOmHvYvrXM
+eKIwabiW4+9BOiOpHt8j5I+m4GlHRrUzU6nqkkxu0rf7XUniQoGYZb+HwktKiRK
SOuTQgRmsT1KYpd5acJ6oJJCIaAyBoFCWpa3fmIgXKjNGOUd0XZf0NVtTQviCnJx
myEVmSW84dRLHDfb/zFv/QME32P380R3ejKsOW19RNk5eG82WqSCLUBCbnK9aKJx
tWqHHNaxyyjcvi/GOOKFFz7rwSdC08SQPnmmCTYYDqA/SStyG1Z4mnJB+F7EsBF+
WCsZYub1ojFEkq4YNmLuDcMXnrFOdbvUlxBgNrCmvBuL2S3lS7F61Obxzs1FkSAD
9FpnTKRinIjYau5lPfHck18Tn26aYxFq/3XUB5p5zWsS5jy/2t1YvPOS7zdOCDOY
ltIGzYLYRsxW2IDaS4RErFlYzlaujriSjzoLLSxynIEPNEjoSuXB1w9kg0TqCXR5
uSHGI5ceuiTgAxJy9Cpuo2CeqB9gj5dh4D5uT8aAr3x02WcQRviMUU+3+ngWzDlS
GhL00uyPXTS3g0a1Mv1nFUcDrPZtFAztU1xdI6U5207rJ7D3g3k1yRHHj+WWnqIA
mqjIlBkR+EwVuJN0LwZhr1H8ncXr6bl3Lf2MNMo0S9Kw3quh+cwT9gVPiWB+d5Od
2fzY2PWpua0aBVl3e2AEcvHm5VNqjUh3YKnJ6kdrPrSA4bfiWDHdydeIGMIJ/SSH
pSq9R49lVWZo9tA5ZBJJfvklzrA/aTQ5o3oJDb6f18Um7+u1f8g/l6pZHALAyz4O
kCrQ2XtdnUFs1eo/qcaiQFZjTCd7dDnjUcZ4Z5Ma6Y0FJyy+Ij+OlXrB6slnVEzW
GHVERz7qYkmck023R1ZsDXcgttVA920CG3GrFLaAF6nrFrXB0zVTYG3dXQdIE62F
vtr/DQltOX/5C+oXg2U1zl0UDF9asRkV8tUnoLU2Ky+pUBZ16KMOuQxogCA2ge3U
PVIE7wAvrYTpjv8fOaKQhGb/rOuNH+BJY5DICpsH1JNHPsNIcjP10Fj3UmE9Hx/7
Kcqilh3rHYTjQN+Aff5V96Mx+LXQ/KVnHkqLhhT/AsT/9AHp10KlMritA8GX7+qt
hO7d8vshk162dtvolZ8dZ7ghCZzmtXx2fUQhGl56FEIYDOked3uU3UNHo54sEnKf
z87pYZMw6m6RqS1KmFyHnVLlHHHxxyx3cfUDLm/01Uf4AiCKTUrdwCEBTMl1QHzA
yludsGsleiNIHnwvA3QcRASVdbAS/lrKHM8T2r0QsPkx16zXtWWNKUzqxo22mmCM
y6Sz1zAdDSL5j02k6zBp00Nx8mchxy/nI1ti9yNztVV0oxaSo99772TXnhFae2fg
Z6Sk2hSFKYyQI4VdNtnAwOiIUw20dNzZS+LWeDspADkpXPQflchuTXNdu/setOET
9vY2km1CpthMdGReZlOJlUyjX72mW0iHOgUdk6LUU4Ih1is0xypU1dLas4/gMcoN
UQu9QmRPe0PkP58D//GM+A/5YQZEMa9gb/Gf7hp6BdnYVh3YZkwg0RW/tj6nvepx
3HUfwFS56lU+R0I3Wxmyq6+loO+NAUwH8VxIoCpT87gSnakdNKnLU5PXxRrfJc/r
cCpMb5AvKX3VL/XDJzIZah6ZUDpNdyx8pfB6cGUkYtM540PR6JJKzRk2mS38FHE7
DAMYfJ9IkVsUD59fKw6F+B3ts2moGv1OhVUb0b8tKMSAK2Bxx+gl2YuMBxX0LGZj
QXDG3hV2KtAzklYBStJXDH6z5QLv0ZnjRAX6eqKziBbU5pu/MhCvqbMjnZHNZJn0
MUnTQU6jeJEtJcbtvPSKr7qITvtG9LG1Bjon7X1qo06b7s3ZHsCs5Eo23+VrQVld
+c4zINPsuLD6daMy+udWmwixma5auHw1aS1ZLb+ypcHZW4ifG5cCAb6/gm2fvFBX
SHH8akaEkDhxhjefzug8nm/bb/jYBKc3ruhlvJCCnG6V2DOfvgQch4zeben3XeJU
JNsy159MwAjH+sg++Z9VLoGnCZzVYFsmIycjCmG2KUyslPhXDwoteZMf6+YIOIBY
PPjdrN9/bdrVeMiIrnkzqTTycU4mSLPglpy64qCySvXGjOkZvPW4GwLo75n/Ekx3
qiKN9GqoPyHFDajnEvwLRT21A3InvlBMWLAhJya4LGmAId8UkGqgOa3pep5Ct8qn
DP7eDps80xr6NPBTKS3ua5Iua0cvPDUH0UV+iACmzgoKpDl4CwWUhlhaUw7tHbfZ
N0HEhk05u/NVJ0xIW9Lzl+Y3Wyeo9s7WbObnpcJFmC9FohFtBtBUtebSvR6Gtrbz
QSqdY5OuRjBMt/Szn9fB0GFRaYonbIWK/9ioPyjmchOIEyav8WcqnRnK5cM1o7XM
ibnnmsT3tId1XHCe39gB74KuaFvczP59p0p/1pG4TdVQQXM4buvkh8UA2YH86rXK
BLT+J/5S+JQwNUSLk911T04h3oJb4iHM5ZSth+V6t3L/gk9ibwX65NN9eegd6QwH
9+u4jV101a/bMkZ3YLErESYs7fDa09Yh4vOE9Ji0FDR/0LBZ7tJTbp/S4aw1x4V+
E96OIor195QexLZcH3qR1ZkcKv/rQhXyU13Y1IGRGEss2w1xbFF8N5z+jll5fPAy
Dlp/Ikel9yEzkCMO0oQ7hjxTG5dtEaRBS9RO7UxZiUJUgjSdJjoO0xXNEg5WT/Ox
7dn9r/bkE7Ro9hOTrO0UXg9dm/uawfuW7kUoYemW+5wXWPYGtdyAvsgxAmDVvwpw
8+dFNUGs7qZHeariGEV2jL27+nveI/YPL3Dc97BxRqcarqNBG40ebPPSSg8oRbh2
rST0WDufWLxfgRq+iHgSdSYjGYJYaAOUe5Xl9pDYoVWMsVkhJlKxe0u9DBpaT5PH
nse/IfwCXkfVigoJX2b/N3febKd68NEO69S1a/SLoh6p991+71ZSv510GMocpmm2
oq+ZCXKGPtmUHym/OUDfiVzp9/FuyQS00TVkp+IeSF1g8ElpgM09uMzDt5wLP4ah
vv9Cznru/Lzpp/TlPg42QAO/JnqEUtCBfUqM0Qs8NYEvbpYibYoBZJIrwoDKDNpB
ulL7xlM7fWZCNkCvK1+zIqpnLfdL0hLcEzGv1G+PAZQ/5vDPMNUCw6ISW9vafTLL
cx35Oxic5/CUQRlhAZdMvxc0JS3SDwCF8nZ1IAbJJl0BrgAdQKF9ZffOXYcr3mHU
jiLVUj73kDWJ/xYEssdEL+Qz8mMCfg9Tfi5oHd/ykbX7fA1KUWsIZmoVVst9RCsl
pLK3sDZ0ePPfL/VRi6BJSVYRhcabGFr3GLBJAy12rmp1pbaIaiGHEIYSFhl7kkWz
aXYy1VOPjpq9kEawFpu3afkMokoNZRgKgyca145ER8aoLDsbjhjUUSLm3L4QVsXH
tUwTVNDG0r3fsac9SOOg0UQl6Tv712EMsLJ/Lnblp9sOGxF1Yygo5OkE0iyAesjl
mN+M7kfWNGLrVnnJHz5hfHrPKzMtM7h9kB4+PiphK+Zsh1+JaC4kJx8+HItGBEvE
LLVmhvsn/3WTulrhwe29toLstje7hNPIMSU5lt4t9R1T5Bi1bYemRx6TWIl+avIn
gC3khbejtZBWiIyyVCBqIj78AaLaBpyKDdCZpqQHJCDMhIqUkhDdGyfI6kaZrF1B
hgkdC8t8/jm2mCM62/TAPObA0qHVW8jXX+O27xc1UDkrL34caXBDftUXyWo3KnRc
zWLQ/FwpDidzsO/341CvS/0qDs/mAHMW6+eLY2IPkbXbivi1Pbvntz8WS8zZPxrh
GLm9a8R0ZUfJ1Ce132/qjmlf0A3EmXqcWL2/oAgyKkqV/K6yfPGb0vMs6TRFfMiw
X+alYXfw2hsZjXjWPkERqTdjS2onY4nVhiTQdhwfwSg1F9C4qxMMtp7tLXwTOdoM
XeW7+CySPTsh6k7LBMkaG0zeokfzlQjcX3IwfWpCi6wNlMkjBUbWf5IH0e2m4+E/
doc36kXlTlE4cM9fowSjTSzIGPkeS2L3RzmlAvm/9uKGYxM+suYjJnJc2nRQTdR3
sS29mkcHH8cve14A1Fe/xRApbMolL8HoJ+GnolpO0EK1iMKloOpYeWwvwvfPHsZV
Vhd206hspT3gJ0Z43C5WiiSu/xtz03/FslykmptB4WKKfyNMTjMG0NMIWtBAeRnP
QKHoc7T28WSvg9Q+LJMnY0obJv2vqga063jerYfQXdaYVVsb4T0Dfyj+V05KMJbW
s5XhAl1NiKAgJGHd46/Gr4sCUSH2uDlY4VI+3WoZjeXGPGT3MNGQ7tfAMu2b+D/Q
I44tbnoqiWDEKpLvy8gp6jXS496zeupRPxh0acoMfeSHh0/vPRHCxJHti4M2cgus
Wbbf6ZW73VuNNiyHULyXo2Mw8+Q8jFGKBYbEpdaBpveVcUluhoumc7JpR7+/EZmy
wmgM0flyJdSj6H/w4gsJu6qSpU5rHGWsyb8YnM6vDCMIO3gBhsRet37VhFFcBj4R
GMvXOaj8Ctcj2SxQuBeRDsIhxkVVLtDszIv4At+B+ngfd7/t5IwpfrwnTv1R592+
HKFXecARzT/Oa2GmumrqnDGCxGAVUfDlXSCZqNgHPozpI4LYFKKkeLaS+CEwAeR8
bz2wjwfnd9Tw3YXyV5PsaERvWaCb3t5+4qtY5s5h5CbfNJueJDH/RLDPL7BsF0id
eAmENcCviJlfais5OZt9phcMszkWayVzMIZ4u+jFg/nzhLspMky0GqBT9DZrm0eN
INjwHtehUJ8sXlxTTBGwrgXDn2NvemrZ3JK163R8EW4qb0OaU/y2mRgvqbXgamCi
xY5pv82CLRXy/lZ2bHcrGGiAAtImC/Te0Le7G4fCX2ZN6TP5EdskMLIzhllIyeUX
bpM218v3BuI/It+Dunss9kfmkMgUk4nC1N3vnUTmTKt8BKbMxXsRJYqITjRrLO6V
JQhQ3/fnBnXRON/bs6hvgVQGfBGKvPlC2WnegZYCYG+1QCq2M5EY9oub/uKvXzPn
jBx9LLLHT76Af3MjMuKFUlpWNcH0hbZo3CKsf2RopqFfpQCPh878XJajprtyVoNK
AB+C82PYfoQ0Jx99pLDkwmgQJq9jJGlAztvnyofytzS9/UCNiChGVwsrjEuJpz8c
WoVEdiTTNSuDKilKAI6c0Ngp3EjSpVjS0qye3Hi0FuHvQXVMslNqbiIliwFgl6gn
+sLAhsXS3uT/jF1U8qo+waD0gxD/hIKSXa2J6pJpXAFElqPXvzxttvoHKznQ51Ae
LmtwVAdMM1g5xtMcipBmSlUwPDC3J0Wo722vbqJP8lv62gyEkYuLwgIycedWpaZg
di+lSS65eLTkdeTxSusxbAGrl6DpaDuKlC8zCAeCCPkoYdKVM5LfIMTY5qcxSAMM
TV5qA8NgtkXmyVe4vtnOkc1MXQy17qwGktxci/0chdPV7tOC0c/PSYNOlRKVHAUZ
uToawEE+6nemyobSd3w4N+x2Cz564daqrk+2TS8mLO8sqT3IfFsrcEHQ84MzvWVb
T3PPhpoqYsxjBfo91kfi6t+bKl6L13v5JdKWf1gsK9i5gAVpJeBXdrEhTqrk1NJY
/FIzgQyt+gS7c0othjnYVQ34Zkvqg/4gVak8x4pnFyxYdZnihtuDoklQLPnLji0a
RgU7yQyz4ibDME91qLRViZmN9g2TyZlj7OYRZyUOHq2doFJ2gMrLvds6W0MoA8sU
sidI6jJwZGfMmZdPQm5GJ/JIDySDAqgbmNcUHp673wFwRp4MQZOr4wfly+dtzQbV
RAyAN/w9jw+zZv1UcCTBJi/Tp6/STh6H5JYLBlgqYaSe/OhgeHlvyfq9pNjbEpVL
MBOitg5tli0eQdxnjn0eLeX0XFNaxNIb6sHpPgKgNHZO/dg3HWnoJyGK+Y79EggR
+bxXaE3xbyNbTPQwvwkwxvpVovx9HeOJbLuJLES7fpwV0Qd6ZhhSQF9wCSvZw5ju
TuvY6NrMDlcUrcU2M857Z/FMR1XoTT12G1EGKNT7y4gKLTboIs7Vnd8vmEF1g0qj
h9U/SQEIGTxPrT2tLyqnmobeY/nOERml8oH6DDXELL5fNl5Sn903hETURSHfuxG8
zJc3l8L7zetOkJDKIO5q0D5GLf+enLwpLuLK3IQiniJ+48zxnp4gtk/Q5fPL/PFL
PFfnWc4pJiqPTO205ijO92Vzf1iXx5j0tZ8nGE6vYi7L/SRGzEMNhphzpgqYaYVn
BuHkTw9IbuL4wxtC+dhW6+Z65yDUumtIHLl6by2apldWFmFXXGWnDNRnweNuw09L
abtLpn3AK0nFQ0FlCYY65UCf0kHOn4+gQV69CfS70k/fQ9qKgjlbq6umzVBwl9qi
uYCQI4WPDJpUwEtJFB+m4KDX9cHhseUSh0fqVI5ZZEy4iAYLzdd7sRM/LZrIYfgh
b8Aiep3KgIG/DxeOLfui0pUXT3x78BdcQIKrSHRfvbvG7JsuPm+q/AA+LUZmCoXo
LHV0Xe8AJF52S7lV29YCUQLT53lOiawsNkefPC03XoXvNp7DMMt6qj7j3EHGmx+j
NTrSR2a4BV19YlV2MqsEbJ1JvwLiKZ1n2ekSI+7UQl37gXUTGHLJSoilpnVK5DkF
Nu5pHTfa1O+/U59GWtt79hy5brtHqnf/nTbfwnaElC3jDK7VpoUMiVvRbXSfQ6eU
mLPVz1nQiV3Lmt3uT/iBGRMzyYhLfTyVnhoMhvtea/mz9JOXXJDzuZ1EBVf5AXJX
4XfQMhVKoj31NdnsOMYv8i8BlSLSPDJCiajdf2BX1vjnYUXLnfcofTf2/a0IKYQg
LZrF9DY2r32fcyWOfiRMXbXBK2RuUlCOhUmu45egsb7oVkLVMEn1Lj6Ikp1f2ojy
13+WWMs7MBOqSSOu9/5rsZ9cuqAk2qW7nArItEvzgXyVvOUI2rnnitGWwXfmQNxk
6W9Fs4Gq4o6jSb4MiK+hKw9vJgVlY0piX5QA9KsSQn/1ehgNhL7KT8NCvqDFiaPY
fs7NanoBxTjYXtpeZwq+trA7a6ZKJaoNBobdJdXyqEra970ZfnIDmkIxf2H0RoyC
a91vnMYChYOsTjcbJKEITsO1bhPJ/mDuSkEqDcaZA/QGoUUrL9vusE79v3PPjwD1
xtwmtLbkayhdQZoA2K6t8jFTk1B6ta8d9fZCc+wm2CF6nAacUFC8mQLWoCHmSmq7
Jp/wsoV68ljEE82PqJmXY/E1DIak0ro0BgbodmO0IXbshEgNjx91kLOfjJ/DKRI2
c3knH0QdN5WsAZrfP3LF0qfJRynBd2V6iKSQ+rTbBWFQAMG/p/4r/QtqpnVsk0yf
f7zwW6W9MRi/24e6MsSRNT5kUeSn/pSj/jqNAgWTHVUzuMASW1sBN6mRkOEEfGGm
w6Uw19zamC7tYdfEZv3/z28etDvpWVwOCWdCfswkJ3BbDrwKBPijz06cy3vuq3FH
XoF26tEKVishDcucYa6sQ3QALWwEn4X+EqaP0jHIXDJEYWwadVVykA7eMeEy5w6E
5VyCwfqpBlzRgifGfX/1BhgDjG7IEzjMirh8ocKJEPdAp526Ki/9A3JtVu/lJJrC
rtQOTk9oYVCcy6d3mfL9no4Bj3rzRciDNocaG2daJX+CCBWFPGw3ddmgxdlg09OE
fX9CKTXU89ysMHAcZ7xY6adD8qilk3ln6/GVwY7A6i+K4BPusqu0e0nr89zdBJB+
37bueNZMe97A3i7kEKJiqdZTTmcy5So9YvnfT3NPqz3jaH+lcAjjS4rYqCwDKuyB
wVH1OdX17PexrgXYgmXrIu0IxKppnJuNGBuBZ0m11rEls0HjtxXJSp4htdbRUWaD
VDpTL8R85ERDauw2DHmRNYIpgJsgFJ0kU+5M6+Fc4h6LWGHtH0AoGVpIoWHaiNeu
ZE1cpFxUQJnawR7Tiv7RnteNe0Brdyd/+qEOp7fY3fq+kAv4Bt4hdN179wohCmJp
Q61dNWaH2z3gOc7u9qYLegdfTMCnbps4OC9TCGpHM7EjyBXd4HXbo5OG15dyrU+y
CS18JFrkUh33/AS+YkXAC8w0KYJ4iBFUtbJHp07gkLzUhxDHXN0drHhIAQI5a9QZ
pQKi1Q5G2fi8FqkAyPUd1yO2LbxnaKThBySUasop3aqonwDylurkkdtG5KcjV20H
NoRTcxvl3mkUZjo/1PW3tj4ETDSdp/XVSmecVqmm1Xtw4mJGjyMnmW82twdakwv5
D8g+t0WBmFKpNcIjnNrBGwkKOfi01957hq1t0G8VNlDuSvbD0fXgsmjdZeKwPr16
zrOYZdvC20GeLpNvnjxbamMGqSLbWuWeC4VQKHiTnLXkeHRCR4jMVp+WSq9yF1hw
53po4P38GakD6M9GuZzJEk9eA0hFAJlQd62UOBJBgO1Jfx7g3gEXoF0c+xfTLAtf
ON38CI+q5DF81DqAyPPnQ94dnBqkTakgKqqcep6TuOvUCsXeNGtOWLfRdVRh0NAe
AVa4QRaW0GIDxORpML1c6e4NpVoiVnl0Yjxdlh0EC533NdbXoPJMHQliePGmYXE2
t/jayhYOpFPK9CGDcyJL8LLNE8LeKDKKTm2FYFNpbzhBRDcVWhADNWvb9AhTVGHW
HHPwD7QlNK/X9fEb6gpU67zZqpzQ2M9zITQI7FUk5AA98bzK3tVR55f21cx2y6mx
Lfx3Y0jlLRp57v0FUIWj65A9CKeOJmP67GtStsnyCivW3n8DWfhpmaVC1R/216O4
8/4N4aFSIPFfPgzhm5Yt02u5iFYSTld0zBZEU97t8ZYtzTJbVbCbxS1dWhg/zyqp
J2yyXlu3qTpanp7FBaVoxyO9+LxfL47+IKh30S8fEkA7iR3uSOaVyF0RR2CN6GE1
nnA/Xh0lAKvOD72qYaP9eC9d9++iO2D6bjbTierCdrKjeT9X8uS7x3BT6HZJsdxu
ejZc6LqCPvPab97OQGFW4KtP3Xp9rGkpEbcdqeIONQcx50na8Qh5rTIORvlGaed/
1lECXhtPAc2qQ9j1evxLOQbP2kCSIvtb0FhMukbD669+wkhKd1LsQuKB2CXJfSIT
J5L1wV/MfFTM/1tnkkvr2j4ojqH5k2IZTtPxoLAge/n0WgWgPRabLkfDjrHQZ9Aj
VGdmT3QkO6DAbXpOp2a4W88XeKBKUZRpgCk0MxyFjHr/1GtXDyqASYpPYI+NcWxQ
dMauOWvvxaCz8+rdbDyUVJ46iyak70ijUr5Ji14P+jrA9BHyCeAaeGcTRdPAGU7C
2cad/SykUAOM+NKl7vyUt3lPGYePRkGf2cRmHZmSSOTxT7xPWG+F+OXMsOfsQhoK
SxwdVoZZJrc6qLNV1a2hN4nk1BVZVKV3qqrCAbQWjM7YT/jz8wDjqAgciCqAxsut
UuRK5cWTbeNhDPuyiEGLuWK5OvDgVvjKM4ki8Yo/7k/j/I84sjRyeCBFiRc6KKVI
m3Sbz2+TORDYELWLF/isDuES23oiy8n6VqIZzZzG8c8ylgWKqRFsOWyf10mXQsy5
YboxJ13VxCoJwlUYkdRBIky3YaLTxJJ+fsMNS43UAdtuid2f41mfSGrEYmc9iClf
czKtryhpJyLe1WE37e34wulBb7ovvfX9XjFusObcYtOMoeMXSzVfcd+rG8bhNiQw
QBr1HLDlPwNl7vskrUQaaOv7Hr4Eax4ozE0TdN6f1kQ/MmQskEBJs4V2r7TzKSOM
FzFgvR6hTPgoQLpfyYjQVg3Wo5QmApotFqNLAYvXf5EJhOH0rFW4Me2Z4Cyw406A
i0QXq3vXMymSGmXH5JgKCfs1ML6cl10JckCfyOYQu6VCUV9uj5ETLTkmM8le04kn
68vJtuf0sS15YtZlVcqnk8uHAOKvxas7tbxXmRiutEgdMU8aEwAMjxzuFNHAHUTi
FhaB8xnYscaBPVXshNwjrGe0+5nLoh1BG7uyK8DqNFaf7UkQvKnEeTzGBf1WQbRk
eZj1BMF6ibTCdhcXGpFek/MsGO74Tv7VKf6SYuQE+kNI2Vqhdot9ZQBbtkqU5y0U
Ha71rHEpwKF4NYc191mtJdvZbzYsKwdOuyF1Jds3mr67OSZAM2e8RzLoMRRU5Czx
mtSr5Cjo7sqHyNEpzRnNA7cE1WabV4iBbHReKt/e2xd5h0yUkaSooRW66Iz4twz0
krPJn4kVYB+4j339tQIV3jqvLHTHfTWzsTXMyk6F/Wxc7QN6JCxik/0TLohbL20U
ygDVEtGpKHLShe4YTwxbuDSLgEPTsiSRTGZ2yoD4Zq2B1i1GNs/3F5xE/x6DjpI1
TlZVPtpa8Lg35FykInZ9ZVc7RaKMg+/Mii1BEqUk8QN9aHfXB7LDvYSLvgpHdVwv
rK40vsXf8GXzoANtNiTGd665ztiT0fzzZJkp2XIEwOZtPnYrGt9yu0hfSi+7jpI/
sYT5l8zxOrE0AnBwImIBDI3Xq+CkcIMMjKZ2JyU8GFRt3S859wtaXFDKPOS+aGeM
kdOEI5a/y2Gk5+JkUToKg6ZA2OM727tdVo7WVYoyqNnmCbkCU0LAr48IvaQ3YMqf
x4Yjfdurhl10xmN/0eHHl41gQ00dxjf4JBFp0hftSjdNwvBjiah6RHczimWS5jh9
QWDmTARccWFMsWvfH7uNsmNylPm2io3DSaQ+79h74CHgxtzVa/XZ3ktKHLO2GPrL
hVKpdF7E/65035uqTo1kjru7ZrIcq6D+3Jv1Cvd6FJQu86NqCAytvWMhYrFHPGos
+gf37l/MoQ+5Mx5YHn1cJ3IOJU+NgsH8jH3rTHV+po8tv8m7m6vTr6QWjBzzqwWr
PxdR02RVhT3khjYz+S4AxIZI1eJkAiS0MYuIFjAzPUhjyu+FyLdBjxp/w9d6+TMa
mcXb9x3AWt9o8Na5dTRsTZFK3X9zGhLBSSpymBfVZHlEAw5y+yv2F2eP2I2caj6k
u/exdmjAi+LK1U4z9xX+BEQRVo/PHAVrZjA2fSNoN6pIfao4gHwTooG4wMwnGcXv
Fqh99a4pyZkaPRNGkFI0SQGvuPXLTzD1G/IWv7uiH0qtC/lO2BOAqNO8PLjosiVd
86/U1b0JKqkRlj7jrOzEcIzUvQX4r12OzHP7CNRor8WhcWbqWxCcYqxB2XR2hB/n
QoX/WiZwBXSqv/YAjwpP7DrB189deEtJINLSf5stgCCcuZ11VXm28pby2xUlQiN/
vBIOdNCXv+eQHibTXLsxySp1Fk1mpZcegt53GHGq5u4LBrEP3cQtgsjqbHytYcJG
EJ/FRCyhaoVDMHt0U9AngGkGMQmIFRc8E4ULpxsudz+CG/cxqVyLrjsUlmzPjN03
VScakbcdW72KH0/TrDM2zub78wQbni7UNcBLWuLlIc1OYwRG3zhJ5L8ixyiV6D5c
zbbnc9rIs+8uxUg8O+LskX1P06fH7T+xXn1qjGn5FSR+E27Ez3pYygNILjWdStPj
8eXEShfAtCcouxC1613MqBOsy5d021AdQCLLPzK0p4uis/Isf6+nrVXrSdxfhofY
gta6dAq3GAbc0Zjiig762McP9B4SLFuloo3+ls5+ZK8NwfxEasX4zVkzwKMB7mbO
H7YyPS+yds0JXNojMbKTuHryAzzw1d2vHi+A5HR6ALaPypY++IsZILnBYGhPJHTf
ZW3/K0bkXzQe110ELgCJWcuMzGk4J6ppzKZuVJSoL/TF5S8TO/oCorrllw7VK2bh
tZsR+HI8S0gGuC4ieRBkdgGcZPhU0iifXhTV7JLJk1k02OqRhurOTCg2ZB7l6eVE
FklP4xpHSpj3aCBGEp5NcoJDLcyAP8uvqHNznqcOnH3VFfoYVoSSq8BiWQwAab0N
DZt0n2hlZ9kS7aVbUCgGBhHog4wBILsCfy0xBombZiwhDJ6A99z/m3P9b5kNQ5pn
VGYeJP2PneGy/8kCKi3gI1Ry+Q1VhmorwEfYGn97VxAZA7JNOJUU+WzwOQzhEml3
haTs3ltuOlwYl4hogS0zTw06Ywo+gmYBn6NZRo0NZLdCZush3MfJPXjz5EqTNdXX
6/xGPpH+gblzU/uwaOlkjn0LT9H/1xGnQLKEg0UPrwWBVJ8qy6k9b7jCbyTO0a6Y
oVgKvO44yJBUS4MslmDtEQQjEOJ1UtmQ8x3+/Hs7UJUCJ1dwJrx49k7qZOlctngW
v8bNNlvovTCAssSvOQzE4iLpSXwHjwiRUtM5D1qxR+OULOXFwL6e+NCwAG0FfsUf
oG2EpFC3cHstEyrRBQhZCYsUE+J3nBrzYtzqBU1hBNFhowt/2NMGUSrZVawevq0P
mGH9YOhTXdq6rebwPimsGznb/8nf2s4ksV9KbCBtoNdPWnVbfE8/C03IdbW81X9B
D4Vz/EkGe4zcqC4z6vz+SbyNVov8QnA5tnr9XPWQbNShqmNadGli9g8dUz0Hyel2
MFRbjwLEEEPYmozOmTwdF//uIQcrTI3NenLGl8PxkwE25i1EdeghMWL4BJWwpKqC
cogwfPS4GfkrFmy8jkSMaiacGOgc3RC9/CLOe9AWjR1uL9u/N8zxzkgHFDN6vz2m
BDtiLTlPbK+N1lBtcZCdZmNSQ+NJFwIynyS8qZLwviJuPftkT1StjN24MQGAr2BR
3nQqQwO2z3Bcs3BzEdoWeS7jFVwgv1TNRR7cORVPI8qeNy/XqqtgyBk9SzLC2Rbp
8uevsg596JFJfqSObr6yNchIBaNVn1ZwECk7W2ZruUb7crkz5kuR5jfGZEeRxueR
W6/jC1tor9lUPjCXb28xHWINn7h/77H2zl1JIKiO9KQHPSyxRixZAf1FbmlzoYps
23/9OJub3DcEu++BRSiDeXJiTrrQlApouCDDnf1ber0hDa1fxsr0gnYU0enGoT/d
NsK/2N7ANlYV1kchTylXPzY/fVKmt/QH30jiLf+FnfM5TT5fyjLkE3lEBhQOlTMi
fXqt9TBnHgpf24pGJkbHuFiQ+E1eT1nJxrsQ1U5K6Vkifk+tps/oDXt1bTbJUV1w
GWlcxCSrYHeKhyiXEVGn6xRY7Q32IHDMtciTh2w8GT3bXx98VSh++77Z7uaieNnI
w1kjJxPToX/+s91yGfblrqZc642ToNPJDEiKgJVmIgfoVQzH/VKmmdCbCjYTjsoI
XrdDzJx5XAronvD6JXZwXjl2Vsb00IQp8FMQhgc0+L9LI6PQZFWNyDZghjn2WpY/
TnqnmG74C/4ZvT6HKl/16h7FGXfHQY1RToXYmlsHKLUIAI5PL8UUMaoz5dKqytd9
TL9fmkO7iBYPXxqmqiSqa2FoT9lx95kSlglmwVOpKNmpLOm1vIplv+GuvXCl0laf
QtDFK7S6WK3XOqXvwsPRtdnt8sEU+PZaN2LKUHAuoPFCCT6PCXwFyi95QVuOlp7r
0/t7O4NSbWCzdv8n0uRogGBEMXRna9cJ+LiM6TzMNZpjpXQoRiowLhZ3uGwzWBoZ
9GbaG6Nabqi5gJhPOpADQ2Z0I+0VAa3qkTCYvZgDs+IregrsClonLqflBtnAUlGG
z1xSWIf+BxCMY8BCYayxIDo+fg0e1iA18higyxpCsqZIQvcPFNiXT193pVobF9Fj
ODxC0rA+xOMPhzyzLQ1V31spki0/+unuuHyswwFnl6ufxcNUdXA3xJwaTRB/w6Z1
Z2vHg8AymfNl8Pms7e4tjUwq6viLQaj3kWZ92KPV33kikl1p8Jnzdp5Dlthk08Dp
P/UTwaKYpeQkopv85g0pjCIpfPtI+oBWW4SAeyAbvITOa6J+HGfFiLksieKTSiIs
ONoQTEHP0arv3I9lqiGkASMN0ODgQmDUjBOMp1v2CMiUyUsBWPmvYK1H+Fzw2C7E
OGh8EwfD2NXXcJCFRFgGxjdSVSv7yWKfBa+LfCkVO8pH5M+LZCxan9QCInnWkKsR
lAmbonxLNv4sYIM2RQcju/hvz9Sk3khyXwOsIbhU7DhMjELLGBArBpsdJRZDvxIZ
wWpCJRekXx3Z4Xjnh9NHphXzk3XsB7SSPy6GGxs3fNDuhW+cM7XzowDZae1zNPk3
+vN/j8xVybumIj6oQZNaNqpg75vwr6Ge63+MEkYnyGJlpMwJN3Iv/yUSA9Khf4Lg
p13jqBOC5CqRX9VhHoV22654MA+oLkr5tKpuFQErs6JA15lJS1gKb+erMyu5EfDj
RBx2R2DN6Fh9qMqb1ZpgPbvTmX18UROOvWdC4njaMaTRIkjs/RuMS/dhOIXTRrMo
6cKYZcO+iv+RJLDn6uiMpSH7cVwz6PhbmLDImu/2l4TPDRy2U0/OgmAc6zG/+u3X
8zgysUdCJL/pNeCLL+qV7koW4MA7ZDrSMM/6cSnRTRJahSLtPFVORbCkF5liotCE
1SG1qtNjtvlUCmUda3hCQy4Y4xtl43w2IXE2mJtasSKYGMTa+S+ndLfIWUXx89OL
w4wetpSyFrBbZw+DeamSCLNjAgXX0gk0YTA1nVg2tlqioiUDDfUHMO9hveshA1E0
MTaHhWgfDuvboAzBlljA7twP+oNKxy7MRF6kaQms6FrawVA9WLQbyJxgxcMmj80E
kxAngnONWSH7xvTy2Aczw3m2H9ph+hkv+qbXHUuIv42d1wFfa/mJlAKoFqz8Ore/
khiPKa3Kfjlr2VaymFN7AOTN5PSVf6xG4HMghdS3jwUfGqtIeuUNMIhP4oO/RclU
QWoiUo5cEWNOx579Esb9TrRoknNnBmB8Z73kFffNobiv/dsyEZmUNfKBDyGzehLE
K+zPusmXgDl7tfkqsT01tBs1r0nd3WbfS3GMHV1vt1VpCq5SnamakjPyUx2jOMo9
wME6e/bL6exk3zqW6HLyp8Dn5TL/0kZJNiwYGKRMouZDGHezhMraL53Xv2mT9ucg
Q6mC/tW9IjW1gG7zEccPQb4032811wsreFkA4ZF6aCHeN0YDkjkDSSNfvpBbtEEw
JdXDZDIe0faBRhg2eMUBaSPcygPdGIondpWwAwhc4ycJjSegCIFwY5JbXoZ2YvVR
l27nZFS2uZLQquPpzIuwMyZsIcRqSFMKOs/zmFZBR1OWcVqysC/49aNakwp2L4tJ
BkLqPXLVRN4mWGntwoNW5oyiWit/MIfw+hsJFVpF+81tBWTIwp3KO8SNbfMSC5EG
r9rucTFxDmBdEq/56Bp0phZLWGNYbrHTeS+1MlXx/cNgtqnwvSqC1Ud7uNaz/Iyq
7bu0wESQ+7Ij/EcK9oGFUKk0t7KNPIq8s2msJdeAsTbHzVnBYjhfIOYdtmlWPaQO
BDuOq04+6yFgKnzTmmFLIlLZLF/stQGKAOrpf/6CFonTVKz13OJdNwHfryTZkRK0
X93FunQRI/7i/Ne6nG1fVgN5qdiI0PCpeLaQHerPjPMguSBWyjk8pPXH311B/yNX
nlg2X4HDQWN+hXvNjdAxJMWTlMClt+7Jx7mB6I5n11w7RXWrS1xeORWtKIcVJsjW
TmcemH9Gmmew7aAp2/BvBWsAWgRF9nB580e4xKl2deT8ycuNP1E2vJXFy6EPxbIp
wTjiIW3AOrq2b+y8+yOs+0kw+vw39CN8K82mYBcxvAejXDdA3UWNpt3yM+Xwb0iP
AFx0XsLonj/KXMd+UZHIbzHVxIOFQbIHnyGhVZi+HhcP8R/sbqVNuMkWVFANXOLo
IKmS5Kpmj5sI9pFgfNXxLyoANfdlPh3uLgo9bM4TuIv/DxZPQQnfuwx4IQ0mN0bb
anX5qGe5PsLyhbOnrbrkuMc1cTVHBIvD8ZJnBd9wmTJA9iAsihWgMLlTZBWRiYOS
YKAZBvqJq93NasixYqrd4TQ509zcsI8wGds07J7sH1QFWkPgJWxmM4NfMQFijcno
Y0rK45iXLDthmBcMtC5GcqDuxbPu7jzjY5Hj47l/25qZh30XrzGQztKopS6YjkSy
ziNaWxmJuIA2+c9xCOFO1JBr/xJcphSCmHkaFZ12LUXU976Zt5WeePBmogXdDTRC
qsJlLj96TzQOYfWdbyDkOJWxXfCWWIt59tI4JizSGi7WrB8FgjcsQfXWsDQFt6pX
0jmX5ExZMjoJMuuVB3/u1VqERIyYSGApRe4EHYNmzt/pjynYGp7QfSH6DTmnOAFg
5YpL9ppjVmeKfsnipj/dWicWfSt1zIcOhpkVgJIU/yDhZraJSLlQ5x3+Qw0QpBjZ
aXE2VmON++Vk/1Lxe9VC92YZcUIsO7JFl709lSj/2mxavL/7zAzsKoIOX74PK5X/
9SrIoUBUgA1+8KUTd0Vl+kZO1EWvd5iY5xsO+zOdJT4YFEcKAbQdhtXFkXQd9HOu
JRvk4CsK4PpFU+Fz9qvywfNQ4RE2UxSqYEiWoozNLYmKX6OAyGhK0p9AjF/rUiU7
jqewHsCn3sBOXyeQzSMkykijfrhFBYgNd4Bzjw9kEiI7+uEvkbO/oVwrZplp5iwS
wLRhltq82lUE++en+tAMB9Bsi5Y+F+tzFWUo0RMopdhn+h06Gg2iavnaYioulAeb
DtawjwqBSFCHIBB39Y1jkiqQlBSWVgRv0K6kAsgw47q0xEmoq//Q8aZ+mWGJaX8f
lne845wFIscZhZvJCuNRdKlQPbwYixDGd9p3Ijz8YgeBOzVL+VvJdW0DoLydDLgD
L7cSq3RHewXLAkB6vGj6E0uwVb94um/1XIVzuEDQUnFiQrXmo33SicvzneaCsroL
3ijN04Rjc+gQ1b3TiyBkv8zA/yqks3Ej4CkKO2tL/uAXbXBI8MjqoVgnw9S42xlO
shKRpnnCi7mudnadWvue3PatGDKQARl/gwbLw1D7FVoM+Yrq4edf3ZSyI2taLRqb
OBoR5+Ogpy27/Ivxwao8ZP97R/V9Du/VSqxK5GD35rm/ifsgS30CE1rYHP8HQ2Yb
EwHn3G5QIWPA3P9JfgpGMpAFQydNh52eYc77uFCW/EDfsFQ9yo8TFMLfTLqPNIxC
Ep1V8Kgcq8UMF74TzbGZyqFXo4Rranz4czh1UlVFiPFas3CW+oCndeQ2BSmhmHnm
oHhgVUzyoMUjC0cY6kx7xNwJo/HMuT4m+WY8+8bzAoyK5PQ3x11bsdskaG6o4kyd
aCsmjEciQFtzUVr3/RrFaL9nWXfxbgsmOQxG1AiMHTSvsaIKE6BlTkFCfZpZZfT2
cNaGfBGL7heuDxEw8jj1YvMwXYTUNOyfy0pQFMaiAC+zYtR5tSsqMZYcSiAnaVI4
P986T3VQ92t90p20A9W+a8jXTcW8niQtqus3HJNqFHFfLixBdkTHwDLXcz0BrgKi
b18HJxtyOFjns7h8wBliU6Sz3IBqQ4q8bQgBqfStpUloEsJ+YUwqJmdbo8Xfi1IB
8h5yD1a3FwCUIYn18oie2jbVsV+EgKxdklQ2tzS0FILUXNED/GQx3o/CiNdCqe69
NYg7LKaHPaNGjJ60Vs8uYMY5POkOVcEMt+E+ooiqomxkwc83K8bI+qTFokJVSy12
0PsQZJRaQxtepjhu9YvgqFsj/SPCUCjAVD8mOaRz1Qi23RDSKVN8W9DRD/4Yy20H
3dX/ITmr+EfEu96cKgMIYZcsmQshnKYo18hSZCr1nJLXnq/U99SCmHRnwF4EayLI
HTLwchKyVvO8gTbac5c7Z3bBGRMgLPKgbasvyJuPHVeX1NHmD3y0pK+yZT5KSAwU
MVzmAyKwCgTO76corOsSoJcLVchMinJNsOXI+CxHkHPAL+ZR0LCWsAyvjlRAyLB2
jUaH2241u785Td4XXlV5vpYhVNVW1LaV46wnax1eYhaObkhEAT6ZBiyXrcIfBbba
UfrJa5qBuKFS4GhxqKCknbHoORF+b1PB4UcEfGW5rhy+ZWkxy9dXwMq15/NHX/lY
jCdktMVlaGLemeW98+FY/n2Xx59Ez2qlUjyB1Tv+0RbFurqnY+bgM7EAbb1ykzip
lYDqW2mXoPGPhNgbG/Rck5psvxegmWPnYsHxhVpiVEpyJT5vMVMFQ5d0yUavE8mE
wnXZ0pwP7Ud1wxBJZFpHalr7thfcbq9y9tpWCYjJlLmRhqE4BrbzQR3s8j2K3UNr
gFSaCbAqP0vQfSJPeNJmtEEpFXNmQepk0JDiSryInly6nwSqnnyCCpZS+Oq7DLVN
Muv44LjIXH72gUNxvUOl0a/UnGwUcAiCLj7r77Dt0Qe4gk/LGmnUGZutLC0B7PRI
p/zSI+n3EdCVJU2c+JQ06/cFOJuRRKiiovieTEjtLQstVD5luybKhtzhgNJYoZ4Y
4hxjpljVeBVWMWrcEn/FLp0mz8af7kmnC5BbwfUrNs2w6ocn1+Rb7metgK/yf73z
J1VvYWSUulM9OUaKjV76bG6wDPxgihPf2xozPY9+eWj5eXl/JELVV/ZffPtTwrm5
c/USMH9LjtYh5qNFnesAxdK48/1NXpd/h9BR3z6Y3VSQvsLfWIjIEEVyy5VOS3W3
6OJ3lK/Z0TgtVCOjUlrVR07GzXcJvK6VKGVrK0y2RPoep5Advt7pwc6gmeAPAhSq
iB8SRMpvhH0hIAX9h6lgk4AcsKWp1K4H3r6ssZWHOH3/pgqN6PuDNPgTQIS2T6ya
v2YBE9r1sUs5b6es9zJpc59xLhew1sqYWYqU4CUwHLP7vssdk2WCHinfqphd3Qli
likhpn3I4NzAz4Br2WQc8/r/hZY+9fAOrJABz5T6rNSDMjIsU/AMgX80UyLGunF5
GDCB0+cDLGNsTT7V5JXDhUtoD/zFNE+c1EMM/T639x1XGsFdU/Oy3iCpv5BC0ZA3
wJ2MVTnDIeHCOFPL2gKGh8WBa55Fjita0NOETmvREypBRU6htiQxE2LiIgadaOh/
AhhQOxsM4xbD19DkwexZzrOtY1hYlwPK2HNU5CLDiPSYmDEQBL/Lc8iCj5wHk55t
gSKaJUFpFcayQp9Y8VgxOg4/AXAFEPp0D+usCNRcJZIxUaSuJz3vb2++ecBt1zn0
bMiu8nuMX4/JOQ2BQEpojgj4HJrlaQCyVCYtjBjFVN6nr1bdzODq90WmDMXVwr1R
iHslGq9y9ovW66G3OXkBGeokvMVWlLOqzUqUwqWxv9Frb1bVAG146QgRnk624UjU
TfxjPRSkI2cqrRz/yGXSkAs6a46dk4SfGALA7U3tl1yBKm9NDKP7PAGTxMq/K6vT
PeHzYsUpzTkRX66qhwO9um3pjlZZc+CYBcVaAwjTZUVnyafDR7eMfqzIdqWdheMv
lLzw5R7CVdUg+soAwAjLXHNHC1BaA3jIqEU6JqKj5SSnya5ccTFjfaTn4cHkAVKv
XYmMEQtg2trINKsn6gkhuPjKFcS7lxxxbyvN4Ga/oU9juHxw1YjbkKzFdsHz5NvH
fl36RVasI8CQsKXuxqtfFNN9jYoq+U9ouhSWyE7229JToRh1jivMIJXWjUKBG3cG
Ec0GX9zlwn4rI6RN5IG8OrZ4jlqW3XsGh2Fd44b1iRo8VJB59FIBM8nHrUHR3bWm
Rw46HBc3R+NbsrC8rhsdGhJ/G6vEcuMC4wVFxekldNTA3kU+NYXacyLYbWd/VRH/
/c13VEV7fq9P9mGRhiMV9vrIUPQveqSv+OJIQo7oJQlakjF3Ih2PNTaZnsCqd5+T
s4g83PLfu4dQIKhIIyGZo2Ta8R36dm0zHU171Ya22N1jOALwkvFjrEW+L/cwyd/M
MXOuT3tVWbHcjgptcKz859T5/I8Q5un0mNp2Zetfc5NShPtgfey/JypU9zvfHqJ2
XdLo/XPfSMiM/WlVjU+eohx5zyG8TbHebpdN18VEhqKG/E38VAzEaFP9SGpXLFAo
MKa5uVq7QqMOc8S4B8uUvgfGlutXtV2ZkkqJkzpJQA95Gt0FTy4h2URn6vexDhLV
Oh0FDVDpLcPzWvGY+358+1rGDWisLO62uz17ffddbzY8ErIB74Go5Wy7sITQDrB7
iMOHAI1OxxwJS75mcla5SACB822iIhdH3rnN6nKP/DNHafmuVYZpeLS+cQM1rhwU
4Uyavl3FVrr8+Y3ghU6NgLqwkaffTS50hueYAKIdQxnkv3XtP0YiMDU1G2Yjhauy
XU2rae2cgnoWG/xOsc7rJ9/eBjgz/Gi/V7IqAGve1gplX9JZDKhGLSZZHvzefrvx
ampQPPVY3ckheBUH5BkQY8CVuCzdCbrzxMA9SuNv7ZLUreaM0xy/uSis/4B62pl/
iVDl218aIN9epyeLeBCUZC4mvx1a2zPMyg8VrilkpIMff8NpDn/yI7+/dXyzW3xh
oIYd/1/sVxqTrjqz5P5oZnsLzHAtFHA/MeZGvjEt3zYJWqG0D0RMqFWAP4ygit8F
6+2Zo2LQqRQQgVhZCPutoXGSeZsJQCA7VUZ+Ndyo8fTH8VBn4wLz6D96Y9VmKcfW
qWnBOBTFRHVWr9T/ShFGhSWhd7eR8zPjGCf4+JSDI1Ox8ck8roC82ecBZDO52kBw
c3fs6jQgyYMbJVtGbMI6aG38x4GavzP35tpJSnFvrk4T1qIPzSGXww3zbRYT6qel
Wx6WW7VcCGzokNh526emj3CC7+Lm1pTR4+2YGBGGTl2b4Pzp3bXAp3Oxym+p6fmn
9xb7l3v7SddqJ2fO+SryQnPbG9woUFt8/r96CEq/aNesQOFP+YKjLK6JQ8+FRA5I
T0VnX42sgkQi/jy+uz3JOUNs2ORnzNMUWa6k03hGQPRmuWq0XuRLLw50qiC89eUc
RNZG2bQ+M+gfJHpgE4Usb2dHVweS4JLGdB706NF262Y0UCsmBSfG9Vr+H3cEovcb
+yuLogtjOWomkrCq+b0TuIQeu6mJtvm0mADNhmXkm5Y3RYDvhKV5b5Kt0PWAPTWW
c69n+fChvF+c0Mi7nYTKA2E7Eh746Emi5xWtoy28FMRd8pwsC2LPdEcOvTC0Gjil
YYiqIa6iQzC+/UX2VQoFUREZ8kdM/REQizxVnsHoBD0i9RbXSDYvrLtdG2/zBZxA
u+dbsM+1qeqGzHbAbRIFVwTakuLsSwb4PwHfryM68GfFdmTtvSYZ1dzQcBULVbA4
rCnbPbilFNt7bJbh89A+8RLCIS2oR/8Y6o6LyB5FipNB7I1SHegZyvHyDFwP7u5V
ywiFtm36ogzioSDbbbV5sVv7DbkeND817aHnVu/yzZFHgA6p1/jKWR/iKieM+f9E
BrVzXzhSsazXEzR1O2mUGx+nh03pgb6OJ7Tl6l0ZXfB9LnoqFXYGXzyEmI4ib68o
6vJUBUM0BjBGKF01HPOPQ4igVwq982V3XhMWMjuVTXsS9ExwubMYTTV6CJbRLgnG
86vmvgOFTOln9BUZMm6XOl+4pnHJOxUM0PZpeitiWzrdl9tXaR0ja+clNdoohZqE
Ihf+1RZ5qGPG05zkMKQS0y7cAHdmsofbu+BWPhAG76j+WU895BVSxlCvjT+NjMWH
ylZq/RMGmleA1Beo1slem6uq2UDh1WCWUsSJ8DYtDVUwLB7JG2hsB1KkYuWgW390
XcXgy1D6n7pEfsa7nalg/KOvH19hARp82Z4sE9WclkpEMPiEm+hUxNvjDRLP0JN9
USwUIjiaqFsjX3BaF4O+L5FfU2ZQ73viu41X9JlRvbBU4X+3H3w2SEH/zQgVo2hO
Eye2XvKDNT1/lyYflPO8NCTwVOJC7Qkc2MBrXAQj+HJqU3FWWhVS1Zq6BBtQwNOM
hhIfKVCYljgxpDV2QeCkN5R4iIsvqEXA9iNwIrdKu6ZxuX6d6pN0aKmgb8xIX4XQ
oxX7bz6C7MHJJAxghCGmbWNX8/EGZuJCY65GAaqjVeko5hAuRE4JhxkOus7BqKj/
Y1EQ0k3yji0zLmknQxrWk9iOgejjSEjNiSWTpOJVwAgSX6qogzvUMUvJUmiwtlWW
5GZtHDwe4rbvuD8rm8kIQ68KvxsochYqZpBvNJ7Fa5/XGPbCBUSwJBG9KZwPlgB7
PK7r/4NUqULgW7g7RzZVQo8HDXSJVGkk7tfmw2jtiOXm54mspuFAvkorIn/DOMwJ
btBSOgn1vRaFSUV1Za+ThUPRoYkJFef2bFMW+aQLjDVk+3Dx73XhGGXJTyjO2hiX
8rKQKtu6BBT9v4ZjP+bg+gRZePKaHJ0yYIew5/OdFpWxw93f6nlrwPT00SXqV18j
2s3gPEzenanZbYXStB1X2C0gOd9neDcLcPCTKkaPaMlbvJqvp63CwxHK0OuMzmdF
MQrFtNjvAVU20KdmD2pPKH6Cpc+wJYC1r/dUq4YgfhlAwipuELViyI1XkWDeuXFy
5qGsDIL0lbA8UmJgisVX+RObT5BFOLX5LB6P4WliktUhVqUSl6RQyaRCxgBgyjEp
SWrtZnwh6G0aIicZ+E6Vt03es3WkA+cR0HKks/wXkCa4A3CGmKRP+MuuHFKcV4vd
3BGigLTSZwT4UEwL2UZpRO2sbCpRR3nvVZe8Mwz8Lk+bzNCt6s8XQPsGDVQvJIt3
sAk1IfypMGNoeOmY4eW3G4Du+93AtbO0f1cW8jUY8wKuK7Ye8SMtFs9GzCf/baJ/
atdCvyexOo3ZRTO1XFJ/m9+jrti/kBCaUkLOLvVQHfQOr0znIxYLGg2SeWaa9JfO
Q/5ELQa2SnygfsJ6bOMEBULCCw8TaK0TwgHnUqeFEIBoFnOB2q8STgTc65UgmgUe
Zh40RkfzrbgkGEskPt37dcMkrMS9ua9s1hb6kjo5VeFpjRW9SkiAhjm+uq3cINyh
iL/hXLSCqEmsmtptFw9puxIgyDivweFsy5oY1uUvy9gwo+5u66Bc+pBvAxGVK3Wt
KLuHB9ng/zYNx8BG8/u5MylAnIVBsr4+WqQ0VvLe7DNsVHnHWVV5/7Idn4WSCBTf
pnShBGd+JWPHDxZZiUt17PfXfULdi192IOUFfTyeBCQ4mzKbOeEMAfFBafItwBnO
93PB3nW32Tkmml80aKHysCNpHDhZ9wipVHPebnuwMyHWH6I/dh5FIomJBZjO0mvq
OIs6cnCcssh3oZ6ocUktpZ1HE6SBQ8ZODycf/+nV+yhiVkqF6X6Eotx77pw4VUrh
tjMmYOyT/d5CVLyX4w2k109O8EA3If6qZdsIAWdkhQRCbc33sS3I0YPgCM7eE8Zy
f6QJ8ivuZ0MvvN+kW+isvjmv3BUXIH/B3KUwY0RVvI1AVN1ch100zmOouAT3RlID
LVYKpxngiRXtnNODdlODOYKkcfet1bhTQzNU5VkJgfftNiSeft+hypti2z0TDuIT
s9JXLVA6/LhRBgeXlZg3BHwLECbJznILtVz7Axz4ENEcv/fezzX0+axMofVmul02
bytX+VYpJxO6wElm+rTeU2Qs5wsCtYfCPdEtdB3rZxkeOPNdiH8fXPiwCERjw2Ey
OjVm2cyzLMk1LyDqRjsNTWEqOV5n37OwGcjSXcZGELQnSp9lx7s9GUMhTa6Yg+eA
OIhPHep5i8Pndvn+j3iNzAkp243TXh4RuTQompg47SKmM5OOQPTRZCEQ+6mkB7P0
JjfAoSPiwLHCjIBAAXEmXZE9Aji4eYIJxncDT6krx7iRFb8BlgHQk1ZkpFx+ZWmp
0FOt/1L+LefjsKgSDHgLcUtniUL3wDKf6NMDUFtA0wF2zwvbc7xKV93PTgkE2flR
k10MPlGV8uINweJLlbBH0TyFNqXXYmVSlKYBtWsabWpDZ9QJkOU6UjWKYKH5lv/P
gwZiv763TSOVkL5l7zMgLZOUS6WfP6uXMH52gCgw1Mj4xUrChV2lHd695+jtCCR6
Be10eCV8FVjzzG6+8tTkNiWmjET5AK4LSqZDFBWwg6zKnTKDTelxa8tqD18hHSlX
SVYlfLSzk1fE2Ue0oaZquKfxb5w7JEf1pUpvr02DhrPOC/rqQIT4s09AJdSujEiC
VrX3Y+mKfDpC+tCWt38npjcInIVukUIsRyQZgYAg25O1sv9cEZ8PICtM2bqBfiyT
x9MGHP1gTKp+bu414tnX02j3zWF3DN2ZuYa0XEW4WxEXUJTvSjtIIfqGBd7kWlAk
OP6vnAZEm2PU8Srh6tvPnCR7eu6pnSYQf/LtftwoxsglNy7AIEpvwLOovO/cBdPW
sbECX1tF7XPMlr9JTYSD/43gUvLZbcuGOaj3AbdmUrDCOWHxpaqpAOe7P1NWdzfR
DHFdeoesgPtF9T7Aiy66HInmEH0YNSchmHsVKd88mLUoppXV/DmH/vIU+xiQyLqB
YrshMtRL0Jw/CNrql8dbz2SOHlLjJ1c+RX3xVETwAT3aXPBnAMbg1yC1U8+HP6GM
uaGpiDAY8ReTOeTI/KkC5vPO4lLv9ximG9/Jv06A20XPL8NJUdRnwz9kJhUHeNuj
U1R6FN0I++3v03Gx0kFh49s7A9PiHKOMJmQcpQGe3LzH8fgHIFtOWLBRoguWzupe
Y2qBks/0DidurEjNmh3eF2SACBQ+/h9JTFyqCx2svNbj8nGRf0MrjiD0YO6MQbx4
GHQ42gzwr/uzF2dYh0ZcjLDzpzy7fJp+76ruhHGOWtabdIojx1duWwn1qvdVLp2E
H+hibvOBIw/l6lJHXVy+D0DsLuYTzCMTVJ7pSq23RCRk++ee+FEkm0btFzSMuJm4
67faMyPX4lA03AdV6LM9z8+J7cFg+RMxaQA+oGiI8VlKMSnVQ4fgFGttOGljg3dL
jfOJr3XFQnc7wDSlVQ6vPnPV1IEC0l3ZhPJQjH6myv3b/BVR8lr86qe7VmZGFMoz
DBfzp6B7uz9evCw85G+z6E6BVpKTJB9y6kaF8GHJYz3II8GRAy56dInTgFAS7BFe
uLe5jlIF5XlwnGKIcaNjTlz6ZMYlHv1kEA/y69Rt6gE+rsesEBM0YgElm0/YgVQx
jk8rnBhmxVVKsHgH545tawmK0Lua3DxUyntRUXjfg6qxZZGfi3Yxp9oc2bmpENVw
L/jG6jWYY+aKJ/yY13mcUdeSHh8QK1OEFEWJZmu/Fj4yx2gvVfiikI0Tuak5aQT6
ODraQhuac0IjIlrctK9EgaKtsIsZW9fz6xxURpfbPV3/LlwGBxszr4yI1J35dTtm
6bgBNoO5A7MDrI95lE05aCFAExXybYz51aCQs4V0Q5wwbh0vLI2mAwyC5YcNutLb
q5a5QpIXd+Yz+K8KMACe3Lu7ptha0RdVPO5vNO2poAjk3yXbqMi/XDKZ/loqB8Nz
r4EmzJIBNcXI2y12HEwOhUpBDkMEwcP8J2RTHx1pBre9bgS4sSRF2b+5NIfKbzoT
l+yolAkOqm/ALFl0p4JQbg8IXB3GV2Lm326iKCxcLimPR4nK91aBKELsXRjlrcwp
cq6Bp7RKJxe51tmS+KyjKBvl2cLcwXi+YCitIJTi5zDAzWdrEtAMax0QI2mabfAg
+bY5scwynmH4HBqe6pttq3OV0cWSd46fQ9SvzvpYKDuPsxsQcZsB51i5MVESgQBk
ajm3QpGoBzypdsdl86nesIwwtVH0sE/zQXArAhpt3CX5tPIo5Ab2i7HhAMIGItgN
mjeYI8vpPW8Zs9tOcR7smoLElsZjzj8q/dBT4DVsO4QX6kwjwPcI6b5V2jrl+Htx
vw8ZzCJi9s9qlRf6A+H/r+Fh7JU0cv9ec4LeyLxUhuYlLY8VUpHbixgnaqryhy49
GfLS7BcEZg/vWq2VfFZMXx3S8DFC+nxAH8uDrWcjbBTHS2/CMfhXAWRRgM7Qh6g+
PdaqqCrmyv3VBKios3o9/SfPGjJVFcevffmb6GIuh8/qET3ZRB4OUbAUcr5yTOZM
Ho8Ktk0w1Ly73+2L7LaHEsQvkp/kVinefLC9jKmyjJK2jmB968zoXN3mDOPZr4Ys
tBRBPuYIFaE2MhtcxqaIxTAgDw9AkDmcqOps36iQSgjFcESkAkhBpgKH1Xqh2k5o
F79jIV2OtYniuCFoGJufTBEU55wuvj4YPbyxbXuCg0AmeJkR+8tCh/0f0bBA92Ac
XuoPvnByZKsXN7RLFXXqoXnt64NphDUbBMlrmVDzNg62WbDXjexEHAXJKDlXVfg8
4mYnliL6efKCM6YCVwsRg5RIQxtxyRFF68bIulKda0F6FO7PjpZkw6jGw76N++l9
ePTbNjS2LT0Bbu1+O4n1bg3qHHK+6en8L+9THZrx68kNofp1vQkmVo9+NBp65Yxp
E9WVjTBNv/o+ahRMnnSoWSycxJDM4HGED8KmpXDUZ5PBOwwwcF1CtKQwn76p3omk
+RiLuDkBp6kLWsr6HBjqBKiJ5wIqOKabq4Y76TfPpZtxzF7qmBkR69nNZ7iK8h7J
qentXREXrKl9uujtVwVVpWAsSjQWgqTLjL2U2cNVMqVSnuXoi+Yc2bDtFk1+kOBj
8ikUayrVe0OqondY67SG+A+l2mLHxvXGAnzEgLy/eud1kDiBeLH6aml7jGa5ChWW
eVmvOsfDhLRNJ49tbBUqL6WEtq7Q3xXFZkqaUd/d49iljWce6bSioWaavCwFYbKi
VK4PSNqCY0vlh6ZoqoCieAYribqF0/kq+EFCzSdGvFoM7eolwEbi7jczd7ikzXOo
6Sc1TRkssJ4shZwln1wjecFKMq2LJzvNKp2e9E/rV2KJnS6kvaeKyq1N6xrREny8
wYhhofcKQW2Tog3bygNdvwNQRaY1hSf7JUPJUZJJwdHAo80gi7x2ziNo6ZZZhsQe
z/ltOnqM1N+gQfOmgR62pVMUruKEz95+MaL5ubo9NeYrW+Alk3MDPyu8VR0NnnsV
24SuLkCyGNMz500JhedJcITNfmKF/xrZuOABNEsvjbZzOkjg7ULuL/Q3ViNlityb
wCzOfqnbEigR2tPsZ3iBTNs0fEPFOQAJ6/wQnNrfrajywl4Y3C+ceqw7NOpRGvY/
RA6M5pVSVaasCLsSXX965aTcia0Zn/hH9ALoHHc2UVeV4JK4XiTRqxr4lMJVJ3r6
AyBsOiE+UCZr8wEgTVRRFTtI3kcnNXuSMlI7epVqR51B0OEhLhJyc71emjUKSqNS
oL1/NQnpmyRQdVKnXS9bvYK52t+CwlOi+1wAyalusGszO95qOmU/xJxuA3Ryx1u7
SGJwv/CWD+cYbR7pH2+36By01RJOhictW5v1j3h6vglWF/h9K//lOQLIvTCCX/QJ
N8M9v8FjGZfwtn+3k2vAhlQTlmB9UB+4/bxQwGD/jb9jxkG3BWmtFT85nEG/VJaw
dxkegnX3hcC44U5OMv7GbHr5Mj+zcllnEeA0H2C2kFE8S+O+W6Jfb+250KxEz2bh
AAZRYwxNwTZrQUaw/ehP/HSL6Fs84W7pTmUML2WGUNYfF1/MN7PLj7BBA+qkTeXs
1FWCCLL+viC89B+MNnK5ZauL7Bm/9RsIOVPJNFUx5R4GKkyP2mTiH6FiYetjFFCp
WT1nbDjgvxagoHVSOB8QTrz+WXAKWlMEumNKOG5Kq/6f7Fj1QTsYDj3tsk/e4hUK
HJU2CtjiJyeV4q2G81LRO4205oR1rp5DUU+R8UTS6xaHwFicBLCDxi+m13+EWEsI
Qn9mN1PksEdhHtahmCEE4HbS4J0RduLWxRmDQ0tMjw8qYwQcpWDqEClxNi07cbyL
KUOiE484NwnElfiwfOjyEjAyTCtqgO1SgNOWcFiQNqGpbaomhYSWPpQU0WGBjuNL
8+xB1xe28Kz7MoCcAwiKCu7l9dUkTX2d9XKYri74shyRkE7XbWurM4JaOEyhscof
BA6VxlvXWlZqSixWD1iF0xIO9f5kVYddn+zjE4aiAYGskkkoMiGXi//Xb9TqrO1e
IjnDfr0sdwZoEjC8U+fuSw/EdACQdJYJYLVvHUICBC82mIkUhxDAylCjm2L7SM//
0+kZjaOoxeQszpdxqSfbXqyz2eIT86QfM68FDK232uSs4jhyhdFdnxgiZIyi3dti
ASFF7IwO+cZFZxQVjwNiSbdL4TgvihjjUFk4C3lq1S+IXOxQt+pYuAs9fg+G0RNG
rnrCx25+HoMwTv4bFIsbl4cutS+zFiSQzjFIWKdylhe0fClUPAC/3RIM/21ljTX4
7oV7UxQms9loS58uUTJ2Ov8UwLGvcPkv+Kfm/fyV5gdIjet4Vr82ArCIEJAycn2M
BI+b1ejfhcrVuMYZjaRqsduFjGpmCM8zt+rAVUjDJBqCTqiO/yjqTNJAOV1fdxuV
Zecd2NTJuwv0rHQJzxBNx66usl3S1aWmr0PqYIYasdoaEJ0SksTZ7Q/Fy2YqnAyP
QB6J3xMpnLeKLtzx0VVKNtazDKgtGjfQRQFwsKY3jOJw8OzyB6afb9DxrWJj2OBH
mk/urtHZTG2YYzoApGKp8IjCZFRF1PSuxonBR6ShEDvxFviPMLpObIcSS1NcKjPK
UNelFY6jtiMji6LUq4etJl7cIP6jsCLicocOre258tFw5xvewpQ3wdDM5JmpU9xL
9zw8vfY6hpfApMlPQ+K6VPTDfy+U58Gv2JmRS4h2Dyh2wFWI1goq7vm+SqY9ZQzY
Z6NVFfZZWCP1RyDICs/B4E21AtNlV7U0JBKfJMjGMHgQgjzGOXOy0tPxcle2o5yj
3UoU6PNV8gSTwyZ55OvIYH3BhoHbQZ/bveOdo/lM5tp1L35v+XEpJF7LESlH/lGK
fRd8T2FYXqkI/gke6AFuWP+0KTpBFPk+5ncc3TI8kiGHGR1uJEvkde4Od8IOcfQb
qIrekGwqumRBLfkLeoiBA06qkb8vixRB1Pfu4ZN4YbCtTVCwg/ZUPR2WIaH+24Es
aGfiv06JzgH7O0Nd2IyX1z4xYn6fbcKMY8TqGgi4A5o2XzL6FCwypxPAWbc8SMQp
KxRg38IOmj9NtuuXbSwG6TxOM2SQQpl3JhCR/XsYbS2h18FaY3zaRPSTkiouNqFd
bZNhg7a4bcoQNwcescBRDC+3X8fRXaL3CKVDbYuQmryYnIQiHOTv6W/pcNwCM3rC
9+KF6N9g/Lo95zyKETMaoDFJsrB+ey2Xyz68tuzaczTbsj2zmbsq7ovOiBo9Oh4T
zec+c5aSbVIZMKQClXVL8KBh5u+E2q9637d12Icopk0LPfUkzziLfypO+s7QravY
pwP87P4jQaXlivgTszq9UbTzn4v53wwUv9na496R+ibsCNLFnJkRPbTSJ22F3wre
AEdUL7ctTHDhg9TWA6ncm20XONXFHqol8SpOO4p+oYVLawhQf14AlCpARJXNJ++2
ImGU04psym0OcV+yuyGs/l2YpW8mMPtHCFXetFxfEiMplBjJPljxM6UP9MN0R8yd
E+DQh87WjyN4jVyhcbwwLrJ9tHzJ9ZsxmMic5/7tERIzt7NsePk45UaJViPI2Jax
CpwOSwqjMPrM4SGwfyHOoerEB5kmPObtau0FQbRfAN6sjItVhYxuw9mSW/8VYK7/
PdakmSca4At2tycO0ZT/y45wO7svwLPeekIOLbi3cm15TLnu7lOt/fozWqBQrLfs
NnH3k+chCqqnatdGyeF1DzMpaEOBtzjoZBWjKRsy3osYO/1VoAFW3L/LldNnt+BB
ss/lFu0F6su49UngUbhELqOPOD116MygTnQvkLuAdWouc5JKQ18D4koNMzxxOUEK
INOtoN2bdW93+VmA6o5dgaO25Ao2lL54EcEqGLvfDluWRRVZ6+4dV+6qebRb6Zb5
0SCKJBmBQbDo8sEPHMISazrIE6zUax9/nGotPv0erED+d82CEsq31pg9RD5JJj1k
d3jzKO5D9Ijf8iWi/aBOtQitxLTOF/eCEQAFHERRl15w3KZxKTzRqEVIC/Adm/rD
wC7TcR98oEeKwVGVBxNQ+GYX7dC2vZaBRXqa4Kqqq4Idg7oxo2zJR6zGEIjbT7Ei
1WbvV53xtFOoo10RlN5vxCDlsUU0Md7X9S7dpIO/dFsXHD+IQ2OKCgp9Eyoiu5Ux
RikUg0EezUA7JAQU31nkxErN0c0mmQ27Td0V6jrr3oFK7CdWh1Cf3hmJIyZJdwDl
iaGwCKxi6CezTTeBwq8i2m06iKVcxFxwFovH+h4pPUY9I9qIFYzl1c+NudHl5WT2
w4OlTRJrT04hl3cHJUm+KbzzcYzTh5zaazcw0qhr52gAyZUz7mZDqnm8NCROmzMx
Jgf3oGt+fv0rW3QeDhUndL17OUCJKqHzrwdgEoJRnODelXNyIOaSGLrzr7kB3eEL
0X9Lwd5iN2f/V1S9/LrOt6exVKeCUDDlY4rOD36QUOh6qrpyNBKpf6Jnu8Dckuao
jOLL6z1WmQGKp4JqgQVR50PRHi7eWLGK0Koo8UhZLZr4HEtA+5GEEBa8zppWRytP
KottDU4Dh/ZDGOCT8kRNYDu2RZ7Jl3p8hdLQtr232DpEoeD8lOQegYTGsg+m/P8G
o52aPQ1b01N9FSPm1jfSgd3XGAlZbRigrnJdVVNDLlFX/CIhOe2fYfxAIrn3pBYr
5v6WvcDiJArzWh51x/tvJ/O6t78nQR0JmiQOyHAPNNnIJOUsb+6qKBRp6MZEm0P5
4zfiTPhNpsC6kkcL7xSZHXhWsExYiMvjbUrKPw1uCZKXVseGExxeS+lVimtA3o1s
3JznsB1AiVNpBwDUO8n5dcK/q1VuBiRxdO6kNxkCw4GK8TB2RJ6FcTLxi4SXBtEG
SJD83lSGuJAFfHQJu+OY/kN8kS0n2Y8+KPQwLYR/Y4c/fN2gh+hM6DDGmNJ7MYku
zbND1Wy8VNt8oMuf5YZVjgyTkz7RUMkBi8YmMFEsPj1csnYa668XgsqRHtCxhIYF
MZLORIn0i/Eo06h8CKysg0DE9SURY+2mACxT4LBt7keHFG/0h8OGyPf+0JzwyWKG
pY7jVB2WoivIKEhFovthlRuxf96M5qqpAC9dxqqyj61abe66bAx6uLCq/zz/3o/v
IbOp7NzNKJpmPdsUBBfl+oou87X3mgV8HIBmqTFkXWNNosnc1iex9ud1QTiZ0wVO
wJJHh+eHFby1W/fnKhk86E3LJjooqyGp3U6Sqo7w9kEI7f2bLB5QzBSsdeq9JAn5
16TpC1/hLu4k8sEh40q7/Yp3ci9v3L1cFK9iVAa9PhX6BueUn0l4eJkqjhdK++ZR
ZDGVzgFElghSVh0MGLLoRGAexqXNsyzgDusYM5YcCYuVxTGdM+y/MJrQuxl+0gxF
eWsBy7DSCtfpZXKuVBMv170ucZcw7vrtRblYgB79FVv9280dtpq9uO7KDguivEpp
m9cQVHqtFhIJXTXeZFGZvgtP70g7K8aNIeRKqqFAd5ZciKaHPj//K56GyCC1Ics3
V70ZJ0mOFOlHl1x0KIv3ws7GgZ5Zvf6DV4g5GoCZwmCztjYBnGRfSlpyjmf1/w7o
r3ZP/lPZg5balWLRbsc7E8F6soOl7Lzt1KAoiNP3bwjTIkCXC4c+UUvrhgO3UVY2
p2w7/qM7blesXqHga1wyfDFO5/XX2+ePzOLQCcUpGlGzv6V4QBYi3mzwMRP8qY/m
nN9t38Jx9D1GvptRKbpozqtxghyxLz5DUwmdXSoi5vbJbTuQIdJ/1y5DWg/QMz4j
qj3T2JWKkFSFE7aDUlVM8Q4UVHbQM5FKLODvd7PkQB2UkNC/4WioMBz7ytxfNR/K
4Q6uKC/BiCkLsf+bfogvYkQGHQv/t/hAkVpfAqfXkD5AZw+lKu1pM750UK0vfDRj
ucVKAPGCqkbxu2+T3K+r6ceLFPeij6YGFdQ74HmyB0dWdMvs4fNR5jQjiTBsvnw1
adaKMh9m8KXJYzTHGFbt+wBrTGgzZQEmy3z4ssdjyoHZSCvzF/7OvKb+ZpiRZxBM
RKiXpQQmh6XfiOjoLcOTq5C212mERjrneg+7T0YTaghCauDV4jJM6ZO7aKgODWAw
i5D48UvOKezlbQHQX/k++bIXyi0+9E8GTXGCvtH2AXwLnefaDY7QixfjsJiwKRQT
KcWlwQTA4jjqWjQZKc7CwUMaA89XpMkYYAGQ9I6ChqQImZO8RRjpPKUTtgQfB3nY
LxlTqnHN98A6R4HHfrUd2/A5M3qk9XiKwmXxUhQ3fo4aRP4nDp03camhJpCA/fJB
YVVwcGF+Fu7lUdXK9J8ZNAgFqUxpW4og1tDf4+q1U+nOujs/wKcKsM+VF+RZtV1U
iwxuYp55GkRGymEiLuXh7XmAoTJH1PfgTtRXEwEE1mXesnT0AiASdZ0aexeFuEKz
yZ4VIIP/k0WupxQrHj9Srhh0isLZQXL4koD9a60zEIhFHYJKqNADuqWl/dtWhWbI
T0F3PYgNigmIsel1m1ohNMErzVDCcZ1D7MJpnlg1poaBoCC2t1+csDAzOWAyEgik
c+J5G5pGT8g3iBKGLCFcTmIk9GurFv5dDGt7xoOrX0xcUvA4XZs4tVCz0Px9sZqE
sJJ4wEM7YexWVrBCQU/kEOQNk9JEV/sLe3JuDt5pki18HvYV6LIqeu6Qt3/Uo9rA
kXyy7yR4Dlz6Babi+A7xzAgNoqaKdng2uKrih/R8XL7mIFXkAFh9dxOF/E0nbmKO
UHZVV87jdA8ipK8zY6P/EL09x1FULlxpa3Xd6uQEYRtrf/CQYxJrxeMRo7jaD69P
TUgiNIrPNCnWwQBR5Cc8IMIIPT458kdQDe7I7Fp4Dh4Ilq1vwGGcP9f+VS93EDPw
QuAFE7APg5hgJUepI6QNk4codGP5Ymt8UXLGvHD2I2NS+NJHey9QzRg6M/tGvCgq
1mB39QZPfjKuk+a2xVxCNgnAXNd7R15cxGXRzuSpUVd+RpsT+ayur25VKKaCVyQy
wJ1EUUzJx0z0UDl+qUB7WBPSQqqNxHW9GbU8X+cw0V7SGlnxzvkRELVtjx1ltwr8
DX9Cc5gDITELp1nm94Cw5ImHu3cSF5jJHqaALCgLWOEmAl4ZqKZN1bGPxQ4Rioj+
BbYqEkcSTTQGyLdeB2XaYW4QOJn12pBUznx9Ms59A4EE+ZIL2kNIABpH9bWlkdrx
bFRfGoPxqCNrCGcilbH9lJPPPxqN4JjxfSK6dysHB+uz/C+kW1LH8ekJWSPJSR5h
pPF0Fei1zR5xavo5d1lTuO1zfCbo1h0huFSIeyZlj7fMyeuO3fGrXZ35OfuvmzPB
Vf+s/wCkuaeJ2ZVwJuNdjVEH7Re8BS2Z3ZZKh4WA6x6Z3V4MDgj75zg/yTKfbK9L
YZ0OJQ1Iihww+4bA8Xc99XXh+0UweZGWMMuTT0JmF3SZmJFHqe3bjs60WTa05xiW
w8rbxTsamwC3mYPACe7uiuKQIyTqVB142LmojuyDphkuS6UoMA+TnN0ReggDi71t
1mER3uwvCiZmmdgmO7hZs79gu96ww8jW038YHlzLsUCTKL2U/KlgBGrFj80I+kgF
HVDE3OP9OucrSKuwx4fU2uQOyTY09oP3K9m9lHU1M65EHBuzQvhuay3UaU4Q5nC0
oXW5CMnQjNcto2gII0fj2fbaVrRvwQ+3QK4KirSElJyOBLdA6hgMTlxqFhkuBSqY
kvXlrBC88+sShpD0ypI8Fi2VgAH3Cd9SBqmJPXz9ixiwXUu9mi1RtrCIhri02CXp
mRbncJL5N7JQ8xmQtrcVGyV0b3uSmY6giEyaWBw80H8Z5QlG8tgk7thkWfXvfXAn
tJ4Afwl8iLGD3+vFdWkzPL2XpIA561UZzbVuk0MSBhd4ReyKBDztGuXfpuIRrLcM
IJrXXaxhrm5c3wcHVMXlfD0FDEK5L6FThRja50s57QQFjzQGxh8zM2DouxWm6INW
b8VQ0wha7CDyfHTeLMYGobemz55e4G1xGw7/AcZfJXTT1MTfvozDiI4wD2z5o3H2
royrq5NtBv9CMPVqsU87Jg/aArjf6yRDpfdC9ytd3faj8205UVNal11ULw1EQiP+
OFRLbkeXuW8D23GvFQoug9LpHsyjOH23fMqpkO1HrjIpc9DxRPVK6RYuIt3uxoTF
eF+30WVdq3F9ylfIDvBVShAQm7KABo8tjWBh+UPNUUvmiWhxGL3Rql+b0Bsoo3C/
e0UnGLKnXrzyXuVobSdoEt7bcg+YOlHyqvWW0pJyYtzrM5f74WVzfJ866xhmu5Fy
N9A/NOqeEv7U5oTX93lxSJxyz05hvdUD3YWusnkgpEfFAiYq/jUPCtR+K1LEHTUd
mKazUnl73io8hqSBPXpOsLawLqosnBgBRxpIk4oXKqE9NcptwI90oZFE4TGOzhz7
v9cOc3enOKirCZxyEyPRFA9ddNV4HQTfZYiZeoUjBXrQIHkialVxnqMMat7HrnS7
SIoobjR+Gvrp8Wm/Cxp/gdK8N1K0QxPmOHDeESYTZSTS/mtBx6rKfOtHjje9f+/D
j7St7vPweetId8fSefxGhn+qeXTA0O61PKRPPcCm51vyf94gsf6M16fiHW/ojeS2
h3KrC2TCUGfAPK8GPk07Wqh2WLAmSYRsppf/l9RugDhn55WiFfQogXrCr9D9EnDq
5qJf+apH0zzGSsPYCNKd6FlA6MW2RWXW+9Swofhba23GdstlboLjSWYaAnPy8IL0
X3GNLp4Gm36zTFiQjlH+tE+5L+EGcCV526tRGdfhIC8gN+v/SWGp2bb8gAoHM2R8
shLOh7paUWKXbST8aC0RxCzoX/LSmTbBWm77foVcbCj1FdGkkDJ6o9d7nMDkOsRc
Xl8y3fc/8Iwqhub5c+HcESKOyQFFbtHzhrECqjqv4kE3dr89Wx10sRbj/FL6fzOF
KkButvWE2XsEIvuqavWwbwdoP9on8JlJMszfa+AIaanCKec6mzJkVe4foSxTfE49
RIHgaA5V66YabZ5IfguBjKSj1PaF3vt6PptE8NCG5K+xcTv8nWCXrZi1gQet9zaC
rkYCfLQ1Ng96vbQ7TKrqAlA7O/NX6/T07YoV+3X84fUjS+3Zh88/Hpc4aw9q37KG
+sEGHlPyqO/Dr2OU3aINUXjeSMceBLnXUz6FH/ZfILQLRmgNc/JGrZMtbv29zli9
9UQx2Zt0hIbNhktMczVNxqqbxjHuh5WUlNf5nRaFOyqQ49yK5v6m6jFe432hABUT
cTfvM/Yl5AoND5F/tOSmuFkTdoEIOBs3BsMHKkzUC9I4fO5qxZPiKhX1XnGt7bGg
JdBr0BaY18baP7RBMHKn9JenKMk7KRnRoMl8WiPtE4gjBj7rnRGhVguPz/HAJQ5J
B1VByWevz75EKi2MLK/AWsnjXkFecHcelK8OrPVFdkQz34ZQ61Eyk8owko063GI0
1pBygueKXno0FJGRkp+JrRvJDQtYlfNiTuMXEn/wzEIFcuBDrI7vMTjIYwTGFvUm
bwd6OtDSfrDMoyEgGFuZ46fqoH/ql4rMuJGv11mzkPSjSHZs0EMQNPODHmDosfgF
K3+e7QbFdvz7URfRf9MoYwXJke5u37tQo+C2eWKmjXL4A5SXBoU2TeP05OU/CERa
odMksvU0CjbqZZgk922tHH8x3NFGUMIlqxysBkPOybRpIIjWxH7vsqe5s12/7bUb
6LrExiw1A0C4lsD4X68dZPu/IsVGwCXTqYW2MtzvD0AJXPmPrbT3wHfGUsTA3yiN
P2nByjhG5Nk4nfEyd+pd6fmO2i/S+HPhhvaHnbYzIeAE6x18bWkE2tHnFKN9r62s
dAqSVILghLpRsXVEPw3MrX4tirhf+duTV880HLEBdn91+IWQCUBcShe2+KkhxQ3o
A64Y49LDYsFcqEWe8D6sWuy7XroHAA/pMvUx4birz3QqpqaKBhL0E34+4n+WWU53
RbZmf2Ue0KOV2devixcDwJgNAmKNW83rU13Mw6n3k39/nZtyh3Ix0kREDE2FxwCp
xE7T7Fx63Eby9HKe0OGDNvda38F9Q5zU5TjwZmbRNKUlg+/qBB6/QLiy0jpF199e
ui7uMIAXXOKkus0F2Nr+BRAL8DJ/sKuizZAIehrB5uRtdDNRkRv5XOhqhC2R26yL
a+Trjylf7yecloGthcYctq4El0syyCihuCphZSLel4hDAOX2dmT6pgG7rDct28mu
e4lj4aOe5OjHceYlVcfC8xCUjUVYvAO7TGzrfu9YsPxsRYNAyJq/+R3XIUB68z4S
ED4+kxOzkA1kGrJvljshKqde3CbrHMBlvMbLd7GvclYxms/8lAxrTCtlFMfJYLaw
S+3VYIKpAaJPMlef+oU2XBP4LHAS8dd5hyJGuvId0Sk15rEuy/VmxqN0UeKrWqhi
m8mccfgPum6xmFW7J7t6YuneSsFPek+WtIeI9Wuafm4ebRDx9jMTX5O0UFfCKNWJ
cLB2mSfvMGy7XOUOvpLbnWX0RPG/l3OscIA0Gah11hKGDOv02dNB9gVTqtPPI1x5
t2dxgP9tivrq3Tp0vUSGOcmbT2YHsrUdhUWsZsBI7bCMpTEUQ1SfU1x7qA7yuFki
r9Cnu6efe/QCy8m9sYh8pV75J2nFV/t1E8kiIxu7N6nbZrwuInVDTnK80iXKQ+vO
6j7lZrjYAqgeSdgtAXitf303Bt/X91H6+MHmkvYK2+tJvvULJSV5XO0V5bcKNy4l
C0lmCW7UrLEaUR70hNrXcVDUXGVOoz4e8b4dzZsyZ/igtbi75nLzgMLrXyJotMmZ
bjoe50jUjhKoia66pXL2E/ZzyPz/krkpMwOfKtd9reMGJ0lA21s1AQYYLIRXQv77
APlTkADHDk8iXWLnk1OSvpwWgwgfP9+HY3Q3K8uOp3mSbIhEin0Cx/y5f8Mu3qmW
V2iGR6UkezmER2w4eJzdfMm1WDguJcPBzt7bzneArGl/tE1eYFdF8sF/mgQIGgJ6
vtIIw7jyZxqOLb6zTkYsjd6z1ABTma1XK5Fm9XxaJYCdV6JdIpvbOnWIMD73YXVG
kFy7algVsb2gLacGgxQ8ffR1DXFLypR6p1LSIF6kTg4hUhM4i7OVDmnFCIGVty/Y
bR6rmkiQuljRpr9MUUEgo90HZaiH1ouJ8o+5G9bcF7HSTuUAEHcUoVODUFt21mzg
vUpM/4lUOf8vU9rlgr2kfOT6Z9/p4pE7sc7ntXrT+j3ZUXLIGT1RIFd0SlZctvbM
lCJ5+7ubwuzBGKYzUV9R4EyAa3brCAJ3O785Z/QpzhvCMBVkzp0blyfH7UNCukox
pFybNJLi3ZgwAkSfaWhr3/LOZpAz8FgnRa0t2BqdsgE8bZvVi+JdiNF35cvE5mPY
bpVD3NrOff5CSSCaNfjw2ZDRo/ArVRQTR9X51Gj4m7LEe+FtgCCqqco2WC7uKDPi
eoRHNe7Zo5Kyn9IC/JYdX2kci/zNa8B5qOUpP0OQZ4BPLeBvU/3gU2Ovv4VYlR1o
YaheBdcBB1o6uDaJSLrw6xcDmeNR7crfjuVawGLUChKpC+NUsel2qrEQeQ9dl7st
LscpuGeg0FZdZPyfmSe2N7uBujPGRDp6qMSC50Lsq2yyO/r6KjIotHkcFLAV0ZCX
zABmH3zsiryI47yeXTK6PM++h1P8RTSJ1Ii/7mDR8nqLpthUkpjqz2kDV7Tihthk
6bg+yl9IAeibDPK4ZvfSQPoRH3OAP2CyEpcVkqO/zc7wInv1S5dPL3IA6HV9gGTF
yLBh5m0tzGBDakva2QqTxByXf1Y1m2G6atcDtyvieidgxrnm1YZDxOhwxv7TZPWK
FBJsLP/lty9X+CyMmp2jv/il4N/m48HyWJtLJsiKIinAWSN4C47QEc2Um7eMqJR7
r2FQHboh4rcmhxR7oqjlqMo1X6xugfIlOIK8oDorb0x/9QzZmwg5FDWdO6DppFb1
A+xNtkwAu0VhIIZKvReJU+1b1tNLHuATxgNj/+dI8XkS0L6IzJhlnZvhN9Hh0SB2
AuHaWtZAfmWFr9o5vdiOxAKgJ5ooXSlTY3uSksEWMnWt3/J1/4zDuky27hdBqU5g
62WQ/B0lG1VlxQmAhpOH9Y7PiTENpV5/G/iITzO/ZW5dIZac7OrGuP8vYrTHHXuu
HKvXLrdx3vjfHIy42fwnrBLaTNJTnpvi70ZEsMUxwElUNWdOYQhW3HsG6SNpDvfX
EsgNYQsWLKFT+aouKHN3k9/YZgx1k2HsRZJ6qKgRbxW63y6q+se/U06FnNyzK55/
EjWuMAPDn6OCfjHErWSLlADvtwBoOJC6VA3/sPTA29Eo/SDpSDJNKlQTpDRs7C4w
QVrYo6kVf6XUpYj5adhTWNlNilg/qgMfgBlBgr4NpFCLIKAFDZFAm96pbgoNmpZW
dbEjzymXWBuwJ9qxTy3i6k5y/BpTAIT7j/P1ie4VfV5MLgZ2gAjFvQVBDHjMwKD6
4e2n3BW8gVMeCOvuhbbW4BVN/mdgJcajUrvAPxELxtXszrsuV1yg8YdFVEgwPu17
LxCQSG9y8oyLAICXSUwWgtUMcPkmDxNl4Fxya5Lh8bTmPdSMGC1wNjNcM8tMCxPx
59Mh0Ta7rdx4d9X11LHb+AHrcTwVfZnN4XfGxGaj1PGWGNlzDvwMhatMGU//Yqwc
f9n1LiRUowpKDbEsTgiAAsR81uMEvE0m7QCcwmcAKQzEALD6Z6T6rfcDJBnhKaM8
zLEpTBCcTZxRmL+MNpcc8fSsRYWIpBSRV7gUUUEmz6xxe3SGiK66uiiHjw7DHPNa
tM8rmPo6qHl96CGxLOI7nKlzbT2chlrNO0EQm8OCtsDu+ObsafzPBugu1U9yMVaG
/Gs/lAspYIpCv0Eq0dmXObWu+pXqM4jnNZ+y8lT1DbUosokfqCf/ntVeMp6txT9x
T9euS9rlpn7Ikx+bY/o5SctQE3fkKPaKtt/t3HlnzNSMZSX29TjoEx/75WWVOB8b
ZS63tfd92uIp+4PCBYuK7ZGO2AQVcHcAXVbBhecQneEK3pJaihSxLBD7Q6VzBuEW
iTNq3uZJj44JYYWQX3Z66xl5eIGtfGfpqgAruLqTQ7t+0XFXoYtZCz2oTJ0loLVi
IlN2XUdwCgEQkfDeZL5GKFCd/KYozUzZlQK/QlPfpZ8u4dHZOCh0ko0aaXAQ+48w
HD0MjuiOYV5gACrnBcXGF+grWrehM8WinnGspKOXZB3xHrWg9PdYJn4w4i2RiOK3
6DweR9YgrM3Iis2TdNcbCBCfGK6Da3SQV2hQ+4yoOT6cDA56yj/z23fWSB8HlyEr
8q/pr7RH+KtRBrrSTRD7rAnYIEej0Gdyy3AXX2Xw9bG/rbvjg+LCNhrAp70KC5Br
Ps9eWsT3behhQOt8Qu5pFRdqZSNOaJNRQmQzfN8iDvdZYh+FwCGDA0Ifatm5g9z4
uX9u+pcglata3sXDja/L7+rIL4ky7YE2/ZGfdCuoDXLKAcsaeuXuZdEf0aCGqEh1
wllcJ/4dWHDokUEjR8TRytRWBngNdNbw8mzks0CpT0HHXfQ2QGUyI1PW8nmH5ZZC
NBkiXCBWgBTwdAQtVDUOBMhSrhDaK1lK/ccLc9zDIOsewDCP4Lbs97pxy0KRwcU6
hIafXBUO8z72Gevy4ZPrAu8bWzW5dMySPJepnonQ5pszhJM79Gmd75w6SdPN5YgR
/N9ls4fZphOItek1cbOAcFpa812FxFUZi2B8qOwMVxxFPBNZlQF0xoevFmTd3eih
GyxwuSHAil7u11XUICsiMSMBS/kol6xNBOYAf7cwJIFvRe3C4RKI6RjE+eL2S+ez
RKpD3ohTr5U5WprHU+CtgjUBJiIqYFVJoVGDBYVd5HSPjv8tZuX0pFWjhWESlWWu
e+mWU1g+vc2gcXVCMQ5f/NRYqLT1tF1JfiIgwC7OTQSMiErIoT5MUayqYSloMiqR
MvD9FNUdq7OKfUlk9XI2buP3PjTcDixHwAUt/GLiwXjS1nlKdcU2zR3Cw6qMsHSN
f0BBv79SiFE0sQoYGHb/DxiJN3ajtRLJruolr8i2weTITkDJl1HkMHhpRadA6kgR
K03A1Fw+e45u+skmtGQ96yuS9cFBNT8WCwtpoJyBaxhIUfhe/OqsF4ApnD3IPfpk
yDxbO2TiXxgVxULNdgmy2L/l1faA467yJmFyRcmsxRifBnDea79EErlN9tfAKCEO
dQiilbP79+Y5FNeiyXjI9fwO9oQJ/DM9qJq03ydBmsQ8/uUs+7eAwOQ+KJRCKHFW
plPGlY43fU55jgS8tl9STOdplrxXFqtIRzWwlezH1nwqwqafg76Yr9l50VtBzFXg
aOulhlfGOlSGPRykSHqMfO9V4B9lGg5iluy8b9g92eR5LE+MGP6r4gSTS0Bs953p
t++bov5NH/CxLh9arD8afNdmswMewijoahPi3xH+x8K33ZZe9sxqTz+tb+5rS0QN
l8MJYrutrgA2uEZ2AJIINKDEoXb6KKxURQ7k2S0FTik8nCYB/MWR52Q3p6fV4ys2
32IhItuTcqBhdSWPoXrye/d/OUZACFfMLqvVkF837aEWfav8Jt6gPVTeaxAph4Fh
aEEjLlbGl/4RsZ7ElYpb91lvF6kG6hvNVZRvk1ATirShUM+A4qrQpIY9d+Wk375a
Zm/QE8dwWyea9oGhMaNC70i+2+F21M5nlJTI8qs2w2n7THKKnZH7AQjOJ9/Nm9q5
40APoEip7l42UCdr06p3lUZMPEKVKt9IYiUtO1eikyAochNXrH0aGbMn16paJg6y
9lR1jb+IL6ppoDkqgAqBVb7sS255d1CBVOl1mA1XHAtzlF8+I0+MS13KV35IQ0MN
dYAmb4B4qnMwN59R4dpLWM2TTuR7pjBguOE4agt+RjweJ0DNZ32RKFt74yyhTNTM
XVn2Evmu4t/c5VOf+n8n4qNFiY+Hgh1unN7UDYjDdKKJDSGj/uNt+ox5+AOZK7b3
p9NztDBmf9ivVwyxrMg4FLc6ye5tGRyTUBJ1HEzTFDp6yLKyqAwtLxLwSFNhJpWY
T37AblpaHcduaYXlJIFn/aHC4NRiWhXeB9jwWC7q9qPh9LQZUTNV8JiD7anhMkdd
vNRgzHOEJfCvgejvuFLiELVsCWz/6xvkW47iXSFEhoL2Smjth5yVf32O1oydp10m
d0h07/1OqZth12R3kClzvoBsKDQ1c8sz9lzgDYHpeZGs9yKyd2YAWBmv17MSl2aL
8BfCqXJ4a2kqlBsWsePfloGlW5au1h+Tp0RDFm7uxqo/V9zQ8mWkCCwFFilbyIHg
LZbaesit7bIxLKVtCJNNqepKGIjm4jvmAmx1G372bqmNZj2nhvwXGQOlbmbd3Bor
/DTC9kmF7w7O24DZs6Qy/0FXGmYRjTLA91pSR18/dU887wJf+qP10Zj4b7hYd75f
W0GWtCLdiQNhDuMP8xWWiCU6lCYx/SzAGkCBhNUtAVNKfkR/nl+QBgMM1eMMFBuw
jlrZLVDlbE3OIlvWiJQINWAXv7Cqiy4y+0TOXwoIYT4Q9QxwiQX60bniSmpFQRJy
FtgiRQG39lqGWVcS/jryzbbjjnrduPJitVjlv5/Q1DtN3Qqm0cjUD+zfjZYY8BwV
2uwwMMCwti2MyKXLMqS3ErKv+9JjKFIoLy5WKQfIDfE67hrqMfAHSUv/HJyHLrf5
zBIkLCDbldd6whXbFdOFom99Cw/C3RoKfqAjduUgZg3ZNPx5Ur0PalqL6zyW2Lv8
Rpgmcs4M1/VItWqurCTLLxYpb91s+BbwWrrwoHAoaGvTBS9DW/6VeFgaG4gdbQsW
ebzfIUzzIsvUSXDPDkuH5xAc7hVcpHNseit4CrDSv4Z7Rjt0q4lFMee6/ahSiMuN
1xyVTp1DGlJI+eA8fkj/1C3A7yibJFc9ONBU69mtUNJmPSMsZ1r/vhjZUE7vM/36
FWWI2ff+tVAvhQpeWA3bPvkkaiMH4o8OzXDeOkjC/d3UK/gbVynZ0lc8oyHdk2/l
RG6VMO3ozJsFDEIBZDmISHnfZ1r7ZorxT7ofu5NBxAw5/dj+fgmS29NFvi2JyIKX
6J0KQTNZSdlttNRR6uq6woGKIeJKnGCTkEP90tMusXR6Gv9X6rHlKcwjCzZ7jb/t
kf3S3rflksDBtYBw8YoN9tutHfa5ugF20cI2JlcKYZI8IkPbJyGFLgb1FU0vsmIH
52z/XNYel7lKCf4aKaKBHvmUs8Wd4UvIfXOMeFu93l/zYGEMNRFFOazmBPYZ0C8t
QuF98OFzrIaLIdIbWjjRPRSkEraAhki8AVBP8zt1aItxXvzgayNyCRFfzPv1CSGQ
/9kgmuAXC4V7RKJgpL8j+putPl5eiZuwY9FwO6xzuG2cNL/4SHR91MFXtm+cD8N2
3XX3HVt45Fr22iXfIybokntleDJmRjsEk8pS4Hesj+ZCUoGpXQ1OYpKVxp61/OBz
oxewP3z341WqsOhwsygnX+9roVK0xvYD3qqifk48xfCzZFtzYw7TzvAGHDAZYWEk
w7B5sgM7nXBEJRzcn7tvyL4LJybe58YTffoYntbdSsD64Qahu6SVUPaeXAWS4IbL
RO8gzSRw+AySWWVODkXZUyAAyiA/Iymew7YB7p7QVpPSr0VSpu+ww60dups7enMX
BM+yJznqk/qOgx5Dhk5LUv9TSrett6RfaNj1l8mOvbXwjz2+9labtEcKolAqE30k
pkTN27lng3F115PfztjpEQuEKjy3knbWaiUAT7LgpemMS2Y9AeBXNOzn9WALQmj/
wq7nCwk4Q65rTceylnxtku9qcee3nw2Y7Vz0KMUjK5CqB4szY3nHxP5AHjQUtgsa
vBNtHAbrNHZo4h9TJtZ+168F5xIYPJXfPah70vY4Zjqjy9ln8aPYIKgdTESHCA97
R9coErIhauIISyOd0bLKTrGMSJydHdQ1Vi8IvVyErRv2WH4te78897FvpWK2CBnd
XH/6tidtZIVQlxNw06LvAJi3e+0kscqyDt46+NQYOnFq30Qx77LBe8fFupCuc40O
FJFJeGYxVWcRlrDhCKbp8/gSgeEprEOEdKzlfg3iZ+s/WlGpuSN7x3xSIISXcECU
4Uvnb/8x93b4KoNfFTA6J1F5HoRfr+5oJ0EWlJsKE7b7z0qYnQHn1pAwFGXv0JcK
1N75lqwIsM1I9m53Io7TPIcdXFSqw9Bd4p5IvrqqTe1a85C1nQudF4Ax/wZLSSDN
LMfHoKbeug5dgT+klbSoZkgQEMheYwWJcOW29v5dURwtUZ9CAFP8rzzqzDyDRMMl
w15Y0btnIByrfxKB8oxuYRgxMIB+UJzJ+wuKw5S7Jx4AyvK02uDlI9rH2/VT+HcI
eURg5LpopqDfXvFOckQaXp76kJ4hlX7fdeIKHCntouvE9M4oc1Hb/HsRimViwgJv
cYvkeM1F0sEJbqb6NwhVm0U+xR2i+105w4AixvT2XAvzH3eqK9gm4DL+Sm2tceRZ
Ycln8K7SoIZSkhV82WouZEwY1pn74Im9Qy1GaMrmi6LmBPbf+/vGsxDRWJcITmh7
FzzeiZ22VuqWNtrr6X50zuEA3q6gzWFXrqxhLYT6wtIlSJNauRh+gXImcNGSYiW/
9ynCNtPF1XMD9LCZ44A6IxqxBiRLcMMF+0kFZZ0TuTib+1vGFyJOrknrovFZxX2A
Da6aclvGq8ID7GfK/C7p2+i4Dqc2IocuTYpRxiYgkV1SgkdasB0wtTEecJCSqhcc
ruGBzUBLpZIvGZlwDq7IkgzDLCJGC1RODfj2dzhrAWlxNa0b4EH6XXMGJ/yXRtI5
n7A9lpLKpcoATaW52f8I7ykZLekw1IjP0h1Re6NZE0RnYGnjLG92jziPdhUXhFds
AGtkdL4R5Qpu9xsYBnVv/X1Aq1Fv52e4FoQnVwK7vHlTLTRRjLzCxwGRC4cLrMyZ
I/5HECpn3NOn9fmjRDWYFUQQSZS8aKddNxfDxgapo35Ed8kCDVWFRjrCHI4yTy1S
6/e40AyJeiir3r8j+4YYhZNP7RCPMBnIU5BxrziABn4gL3DuotvlOqQthKAid2P/
SglNC0x0PgIlgz0G3f10X4bhz/KjRiTaQLlFDXbLB3QBkUjOLSJIJsfgCMqJCdzR
a5+NfFXjBpAsL/LQQdZWj7JGVMmKOt/IfzSkaQbi7pbzxpzilw7I0y6xzKfvWuaJ
rOsQm5z8sGkjhskmZITp5JBK67APSfxUTwo3mx+DJ0blahW6agch9ZcbuqSvyQRY
mofLS273SZPdu8lsklUAxjZKHERzrljN6OGab+9m8nzh8UcP8c4qU3IQxud30eJd
9DtNUDqe0LIirlIAKnl+J6S5xEshncemYofTvsFyBlhsEzimrPlj5fUblvy7PMWL
FpzZfOMVxsAlHrXnH/UwyaCcsx2Xy6ATZnPmVHnOA5FDYFNO7Xscb8GP91yKz/5W
5LUybmthgODX7xzwS5GFvyPUdkc7Kfg92p+KjmzKQwUHapUeOhfCtio+FC8pmSjS
JaBvXD5wyfvNSwg5IGKqoBNsDDBOBA/8QAfNL0HE4vzFhiBL4QUtraNXNozPsRDW
5ULyZLdwDcDDKwjR5nxGUbwyf/5EAgNJQ1Ibn4dzP3DYUnBCzUJnLW4cXUBQEEzb
ODhd9Rv6LuxGBNftR65LVBvAPN81a5Qw95GbO1ahSOwQfghIb9+GJiuh9/EJg7Pt
7XYz7Fzw+D/Nhi4OuQu1PJnyrl6Y7cinW3zPaJARw5CRAgEYuny3dtxEdqCV7zJM
RltD0N3W5i/mejauA5V5Kj+5J3IVWDYz8kaoWQ+y4vc5iA+uH1miuRtyZs8zhozC
Gj2Hf92weU7LQ2do+xME1dFYffPT6nM+lH/Fn9ZiIQp9RSpeGpanyHSmRf4MWsDC
303lRB9frmM9N1Lxq5ZyT0DH1UB5OskPSia26iwwuhBebgkzyX9Cjmx9S7q+fn4O
mSaN0SSLEc8BP+8NILx7Klr0L8HL1zbsx92XMqUAWJNbZ+Pvwwgpq4Lpud2BCq7H
CiOStZS04T3FQtp9LaGOjOe1Dkxqkv1InhFrfrX4F26S9C2GrKRh1TW38xyI+8zZ
uJVlNqxrVIuPowQEB4342yjf9RqZN8ZAODFYD+tUzV0VzJ7VYlL4wQoT3tUGV05X
/2nZrNUm/sH+kDPMpd6ttRMIelDNg/NSTFGrX+XLlSdPv+jwsqksFftp4unixCiB
cTblTUjMtOBnx2/1O1lnlJ4YoKjsHxQhHlhazF1QxRvBPd5y/QQnPuYap8z5ekXy
HjWXTjhUS4hZM1pY38BLUfatYYl5/Ui4TEchex4VG/d6bGLyF4r7xu7ruqcvNKYC
UhCqTj4RLLSfYl3kdIClFxfj3rVjf8S7b+RSfBzMsOWnlhXKtnYL8XBVTP8yRQgX
xkzObc9K/cM2YEKUknF9wVQniokMdws8vZn2179OKG4MYy9JhJZFiX3Ypp22/g3a
n2rLlUog7J9Zv1XpnsVc1HhesSRRKm5IsMi0zlytTMdvy1Pk7EUlzgKGVLeOfHfg
UxJlHRmlquS8w6XogGuhzqu3ITIjhPcPWH7Q0WljWneTs8FMf2Z+906B+tiZaJoX
MLCztel4Nqv9lvamrKS3BhwNlrXC5UYnUCuL5cj0GXuAjZgbRaQVrkZooMu4IQF3
vvoJeQoDEavwcy3Om2Sjr7mrQeTrCGoWAYsnvD0GgqgEN3hvwjRYBRuXDuNiFYWD
3Q1JzzpLzhtnrv+EPD/wfWAtIE7XDNVtqDcxsI7jZhtvkEFBYnjNn+AFdoId4vm7
uDtlEAdtabKhI4VBbpQj37fw7PNWzVotInfzzy132/UHHVnfiVhwACD2uv18QVMx
k4ONY2RZ6QIoQkNGerrwJy9ASeVb4EncfDOfzbihH1boBgfdEqTCV7WVBbvOoH7Z
l+aSlJabYMksACB0MKKDeFZi9tnty5JCt9/tfpw0FMzY3OI9Um0Cz8Qo/Hic7mJK
n1R0jRO9oSwlPlpH3miXK/BOwyzk5tArsoW0acfEB36N+bRGvkfRVrf1VtqUEHjI
4YzP51VDHvd7dE5zwaIm0Z5G7XtEvQveZrxU+E00QR+VvOA8SvIAU0sZ4K+N11GG
Z8oWvH8KOpeG6PcaOQcXCGAu8+bU6Hi8Y6lXf1yDGTHf1GOw0XhtkjISJ+LlEkv8
kZrgzp0ckiYmJVLK7cw4b/dnVCGbcJtDKoZJPpAqgJ5Awf5oFSMvpyy5jkAxPzsB
n/G+0MaToB/sYOa1vF27SALD1yvNrqph8uVD0TJzxUQIb9Gvo12I1/e6XhNwiWVB
7xnugpz3z1GHI8jdy8Z9/uZGBQjKP32clO0cFNMnmEnk5Ob2voyZLe1M+MV9QYjH
XG1yKUKwC/z7+kpEdGYDwW2OEMiPIcEmM3/ovBuFBJQl/f1lAQ1FZzwKbSkUEX5A
DH5EDIxcOALYQnyK9b5tOv5e9mqniFvIFEgVj91g/h2XVbYfRWeEpCotKgB7cxUe
KxCZoUEG7aI+P1870dgKK0K1Gbvw0IzMJJCcBPMZ5kY3xzmmqtVocZOp4YHY1FRK
ONy8+9Ykf/ilDV2oi41ER6Qb2/XReyjMPSkdbNBx9rq8IJmmKnFnzajsYhvEVFo7
N5xpTI8qLYaWomVsi0NFqTt4ld5jBA02XtGZRKj7embk3GxfjTOzvmagF7TTnuOU
eYn3kj92ed3fof60aEBRoBZinCIyzICVDPtLXk1j3joYnuqHir1LLQs8tXF6CZui
ZWQZ3yIPcmyqwv/ylbnLEaPIzeGXa0VJg2uVSnidNDb1vvK/rQF6/l+n+f2jSlr+
9W+6nluLXTVyhMFSCcM+bKnYX8sblQGlYpf1y8yqJnbaPcfOG8u6bVKobRpWPLQo
SLY0MwEw3oR7OlbgxNci88nfE6GxqHmwrVi/p6ici4FQUauhhKiBuxz4r3AWbzyB
k7MaUjFzXl/U8mYmSxYAl/moq/mSlJpuOVI1rS1bSvd1A7ntV7hQLFLSif43B3Nc
Q9L+uLxWMMM6Z6SzuOfNPsrPZo7ZX2btn53D7WIsEGSCiBGyC4FBK2UduCgsreSK
4SOWPwRTnHEe5PSxr2tvA4Roe78JHV9EOJXQDt16F1VG7ze8ExcEJ5A0Z8ZEIVtT
R5ZU1ljrg3d1PBOgia/wL2zRBHT1zqbwInU99DLu/g67YIGBSukCZNmCCSOSAxZo
IwtqEHtuPtbJIfUmEs3iyWLkGktOvUXNpLSFRyi2F7Zq3GgOfYTEWdX7dcuLHnOK
mzQ7w7+GVfXRpsGkfkEm/wBlQ49A1hQwtqFf+gspjEhgpoucsDEjJ8uSjb7B8Wea
x1YPXmS7mCyHjhFK6NtGx2NMp4NJyqYoZzuoOignxrAs+sHJf4aZjTZCoqxAAmCz
4Igmn3+6GqaAI5qDBzH9zaPpOW0bN1/CWumaQICLdZiZyu9IdCWnPjST+KhdIfZv
OmR9OEiJmfBrO2+2iVKuivEY04baoekg2PusRpEP5sl8iQhbdiIIj5cB2QMbvonH
2epZf1S6nccaT3svpAjCrTBR+53uu4co6HcHGxYTo5R/wQ/db8e5aWiucg7dV+1P
qIhJ64jJqVMSwaF3ma0QYgL23S2Glgo5iOoIqeJ70nifLOduQ3mfmby9TsLxvIO5
78aniUPd4Le2Z2e6L84GsvR4K+fDuxw/uGDYA2pAlUBY4rcSQAI0nGSiE8/Ng/YW
xiqr6ylXRpDzRgSh7irZTnsRg545X2/LdG1b1rZNyN2CxOBLoRDsnTBZfXfdsx9c
1AHv+FHFiMhyk1NnVwY+cts0jWyDUgO16bpdKEA/Nj8MjMMwF8yMPNwNLRr6kCvC
waipSt5u3l35m+16MlJUg8MBflim3ZxWCRIxWqfPe44C5795h/GVBOiaPMKTDiT/
2wDKLJkwjMC0dnrZ3cSutubRjeoejRxbe1gkIyKd5Ybw55hdv6eiFaAYbtpZkupe
qI0glMyD+oqCzPY4wEnhAIqnxbeynpJjGfFNG3r+y/xdvgGWNSn+OmFrTaGG6Mpq
CViPnAD8xtOwGrlMEXJv2VKJQ5vSoaLjUydIGOJm1KP76C2g1WZ8nTZ9hSFIpHX/
6qGKdFGZ/wOQc4Z6tYWqw3WnC54SPzxeuFaFPxsBYgS2TY5WZ0ezHcWhTiesUPJL
vReTE/hqcIxPeLnDJcGduMnxVdSI0NZXr2d9U8ZWj18GKpwIgKFZgSiF48gXzOdv
GPOBqK3/Qf8nE7fBUjiaVVjLFcHirFJQRmhjQKEL1Aups9xK/oRmr4q+fZgoUxiE
AwQ1gFlSDXIsQ5oNYoYNMSxkDKRVldt2d5bkQk06ETwCRf85ICfGNPCvE3a4Rei9
aVapisylrHNSw1N4lMBvIE5bnDnxnDXbIkPXz9HkygWBP6SmgSyT8cKhUQs04/eK
tDJybKRe2SKIEfH9gvkscUeI/uPhHIapXQoiozBSkyxytjJNi/aCoZ4Txf1eaD9E
58YHfj8qJnkRn8RX7mULPP/hsRsDOUQlQ2nKMo5DQ/yX4cRZYXO8oYeAo0mVjxhH
isKWqx0uxtb93jfxKnK1sTzNfRdtqqczAG/N3kbwlrKUXrAtJsqnKVMbTPT+0M3f
TATcLulDQGzJAPHK6eMlTGUUWf+ELOG0valf3KmgoD8B6Efxlxn8VTB6cLNDBwSN
zjTpR7++X0HsIjmthMk8WMIMugxqtuS22WT5rFUkXhA/VTHKhBX3YY3oIU22c1G5
TVG3/vCYLlLcMrqr2Poa+WLWsTaUxhkEsFb9agNYg+9kzZz2z7mf5MVUUvjVhcC5
8TWYuNASuqubVnJEcogqXSz3MZ2OvECim03ku64P09i0nxXBYIXBrp4vw0ThJUPO
gZ8W1irIp4iKYdR8ddXtvnQIiWYJCUQTZ2lUAZacQNrcmkfVVDDCWWUAS/Bn6mFH
Gz0ghauQqkLb9cO5WoxCvbRttbmhB0frnNM7O2dsEMjZmNIFrMV+JvFozPn0FZjh
3b8Rgx1YWY3izqq20uhmFKAAgT2j/TOhQMKn5qDcPBJZn8c64UC/01hpEMRmVWzp
dufqUwpvCA7ir9vBBZpeKwOE9z74yAjxyqo1Is/uhBL47BaGshaJVFsQd7uQpwpL
O/BGdukB/fvWmnewRe2GEF+NDQa2DcDRWky25anXrK6tUNrrf60ZBRjY+/An6E91
lKcyMRuGBVKUQQbDFTCC6goiJhp1oOp43TMzOlT0ap7rKYhJs7WS9q8VsFh4cj/l
S0yVXwXUi3RdOMbFDlIE49KJpKaSgrggUZflUst6T6VRsxk4fe/yR4RWe9UJWUAV
YobgL/GpSOWGQbKazpdjssKLqscD1868jEekJNXQSZEUgDJsyKdR2BgjUvDBQhfa
XNRT06bnmHR6EFY49GhapfPKEdSxu43GOF9lAgPRi9copqx9gCkf5Du5JG8NQhe4
wOwAsgQZ6sfDqZ7HgR38pq4Ozm2ryklOclAQ/7xp597WGZ3NvHdCECqD51IVe1sI
Qyuo/ydXK3AumbPdOzLm2ryYEmVEVwUEqyeUqUkpwPrpYBcF76EykaZdqDVxTeGM
PQERqB6ul01CnYLOaZMPXrnFzS7h9/s+mB3GWXoO8zRu8x7mVmQdHQd7SmEZU1oQ
SbrmxQy+M3s2KhXOfCMd0s05Tu4D6Cm52ljUN2RcJoa6GfM9rIZtjDmKC2HU2IC0
biNJRkezvTU3l47+TtyNvfnTJsSnj/vwYz06W3yXGySJhMRg5LbuD2Bj5gYXp8RB
PHHcrnauBV+HYNPVaFWP4ceocez6IFH6xy1sCKNzTBFAASgpnnTIUB+8Md+QmxpB
DVzXyZHSLXb0mo/R45OwOXkHUjHtVNyFArk+Ercrt4PietTf7OC+wivnHK5+6XeG
GSOsL7CSfDW3GjJWjv9EgcBW8mNX9j6r0bCQKdIsnhiu4iU0DJkNs3VuZSEifnBm
uJrtLLJEbog2/WZS92JOnR6TN1Txy3E8Y8iyMDiLWwUflm3DPmqdfKJSpeOzQBOe
t43P+jNGJkbLNkrMIc+vOMKB0dvmXolFryFo/oi2KSXUFJVXvRO6x28Y9s/p1BOr
pcVmMv46O9OS2r5QhIcLDPb7Xw2FVxPGQEJ0IbZGYSihEUpfjGEu0qUWvl91Lwkh
Jb2UjXeCkhZhZbSnmVD55mLJ25Pc010Rk7CucwAW1xNFxHQWExOQ9erEbi8q5MQq
lSVALRNHnxgIfDXyFQR0spGi0DT9kI42kpBK1BhL5x30L8l2Vsg6u55C/9lJSe3v
Nb146hk7+eZy9bz4g7QelGc/cOYjnJmQc4+c19WDPcivszPIEQjJnrRlNgfmOsk/
bSDmadxKCy2QVjEGwauoX1mW0o8PxsMQslcEgTGHQU+opwu5Zujnu0dsND9KqMD5
m+xvzaKWrxjSBOKEqyegsyX4C4JDoDTyEnggZlCx6bTju/e4C9T9OSsJt6bc9ZeV
A6oAxkz8iT09tHCs3+S1sMSt26nEy/u83Cxs6HDvHGzU4Ngx9njD23gNjd0MvHi6
eLHOQubNJtdKvceSEL/iGuirb7vHI/f7mqpZZPJi9z5iAPMrND9VAjShi+ElFp62
pcLTds/4wOCFwdIuoUGpMM5HXNFJw2/MHED0NgqRtUtlT46h2KurBrxIOV0hZbBy
F4xOaPLimlvXMOB0KF0jP3m0UIAA9XRsh7CZegERc0qt+mWyOFYXAhehXEsR8rD4
qYrvNAVkzPIoZYlNKeyNWMgXGUEwzGw5PnbGLaPm/uU2689wqIfI2hbOpLpJ7z1N
NoGqmefB5BDpqW698VCxR07b1XtzdO3jd5fUcf1DdwM0Y2nAAu+pfvtGmWZorGMN
RdmzsLPELbZAcvfefVJaCQgHroNu0pI5qtERK+AOvknQ3966UITF/tWyMwHgLL2J
8WXRp2vmkG/S+KKRwAbfdfd0KF/tSBHLJzitHP5LZrYIiPC+cxql1ujTXoVqKqvE
FIw/m+Ur5c2kTMQMF0QFlKvE1ssNM9ijdACFC/aFoJ2nuECAOnGPDDb9Yo6eCqjq
U0zG6W2DO1z/4UkimcTaB8oDsPiIuTK0YBo1BfB2JxJ8ZUyBgfZmUXiI2kXLONQ1
c8cSeMaOqV/oQFnE78pFzcs6yInxqiXGYx4bbmtJM235F+KGdSPhJqb6BkcJO8cs
cOmQt9KQ4WSO6j+H18z/NGtGZxcfsQaN6RhDhCABlD34gy0l2yh4l0tSmV/fw0l4
GHiz3POXXTcq9Yd8Zjj9tgYPqhtZjezqgZdm0KZ4Z+EW3N/c+Clf/P6gMiW5GXxs
wrt0bV5wYEIDcEcB4tIhqVWZ+Eo8zo1l7OBmm/zNVjI2jhIF/WgpgYvstaJMpAS/
v36LXnvMH+sBQaxHXIEM8f+wvBcuzn4umlkBV7XiDycEmPXzd+98z12H/7UQT8fN
++6/KiTnEgMuLWjjviI5lL+mGh7sHLf1sQmgsKB7rD3HBDPhSwx2xNbWDAB7Qd4l
eXf5YvZcIAg6zxNPi4uMtqTHLsNtRsdZXdIz6/5+7M7r/fY7xHHtDI17ZRMzjf6q
VQhbakTQ7rDD5uZkqHBrXvIt/oQpOOwNAUeKoRZ8G4dk49LZYyd37pCfY5JlxaQj
83Z9TDEjBHVnf3wBTz/+1yayhACDmjxE4M+eI+qVbxPf3ZqOTWh6VkDqrUfTq3b5
xk+Uo8cw4u4QRKX5sz9zDSZb304XDwikb8uHfWhtG3wUxtLT0jtPsrvJ6ZJIboUl
yK3PGKZY1uuwXMu2oyJv19rOjs+yHMIY6/wgDEG2XtJbS9RgKPWg9ENgh2p4/Zmd
xeYqYQYfWB3oMAgLb19duJcK9Ne1qfwsxcU85DfZe5ydKYqpB3dSe9i/rEF4olQ3
+7jP98uuapqeLw125dnao+pvSBBDVEU6mPvbDqG92oe+TmzIadLevpMvmFWzZ2fl
H3Cl3NlabSMFdTK81X3Lu3f3x6JvGUzig0sPYWOO9YQJJ5cezj+allFhIK4ZqxE7
Omq7icWpRN1kPUtXLSFW6oKpg2hafuMmTKkKDcMGHUXjMVi4lnhTu5TWLsqmpRK9
otLan+iPoTbsTG6m2kRzSF2BB0BI/DqTYaRra6Y2Wy5F7NTpr4clV7YjrqMlCxh0
DYb5+9LxlKy35O3+ffweW2g+qfl20RtOKGuFxSVwMGTPwAzNqFnNjl9pBGQ+1pH7
YYzkPxjni2nwdA5kW5ohzL9D8DQvyA4es3J9WzJOrSbD0rRlAueAgjZj5jHflVFo
XPKViB2Yfh9luXBDMEwGtXNxIVeFW6AI/TXMXpU+GGSsRr/HFl20lmHB4og/NlOu
DKlwo+FJ7HfTICFF0Qk4ELS/dxuzO21qwMwwpga5sXsj0vT0fswEaA1NbugM/+Nt
yTZqTIRzRMAK1TWeWkOW7ZY0ETDC3YN0gtwzxf2UlcSddnIWLLgvBiTWJGRpHzEq
aOWEYdB4eEPDjqIIWNObNeT3wCO6N1EulKjPVHfVpE4j7Rx6f3EWmXpV29sPS7hE
djSl8LTd5ZOWbKGMw5JiA3oFn6/SPld7mUJPlqCsjrkYbhOZhBryTbYLvyZ/t25G
S49AOZ9pfJ00xt99xnESdsujRof4jkstr+fQO1cY8FldrmFLiuIC160wogNLig9R
6ikwo6mt4NS8VkyVM6fzPPG/OMYgBGVoUqVVGkcFZvoRlUezMy08QPkXtZ9o+gKJ
cNffglS+nSjkYfN2VUJjFzgePTGC9jdvySK4WCKtieC0JPOG8EmxsY73jFt4z5N0
Qg+PpEga2RUc41v9A5f+ug3diR6+WqA5UKrLzLpv49RTTvnCTx3Szae07aYVgdvI
wCCAPTf2aiTGuy+6v84RQHL3GtsFiAONW95C/0+Qyf8ShhkcYT9CIi6BSHC4EceC
J+ajJWjG8E3w1M03XcYG06x8nxt20KNwT4by1jS7hjdchNywjQcK7wJm0p6LE/r6
OiyJT8QrVAE4Fae2M9c637ljaVM9TUlaBEvxgt2rh3GRS/A0Hmz1WFDU29Q+gCvf
3l4WQTgy3JDqcA0C0qMjDu0UurjCfd9uCzLdsMdHcYemYRIQ41y+h+yhy8IRgm8J
D0ylHklQPgbSh3RiHcaGo9aZQ3CFrdSC3lbvM5AdfEw/T3OzDX2uBaZjF4F6nebE
PFEUcBKqJHpPY3PnPbnU16kis8RxoMlPMw81MolqRSdQmXUWVWb/WH2QY2i2w2a1
CNV7K6GUc8Kehrmptq9wJI5nJjwnixRYCWAe8hdFzEDBIXf9N4rVWEgpr+7jqm1M
GidGCjUV7ZUbaQm+PrbyGRuT1PJnzntxlbBPy9e19st1lid1iPtUwb6zufmcLC91
5/s1bgSUsiAz2Jkf0dxK5uHaHyPSzW8JSL32iFBs2o6kcQ9Z1ta5OodFvL1Wp0EY
ceY0L3q4U96HCbReyhe6drpsI3Q087hYgSQZywk4fDlJStKAjBRa8hAk3vUxcF5W
V+ZUGq7Y4xxXASvNhAx3hEGnpZm99F25ICkuKleYR1+l1I8+ciyT3shDlp8uTeOo
GjaYaMBU1D76mzTwdVy8nM53LgdWftMQfMU3J4+cJ3ZjoGDlb2+Tt3aXNrVF1B0X
3BLjbGSTiuUFZ7HZ6osGAjFHaJbQETadJhYWV2gRInJI/yJfASerEcnL1ttaQ7jC
ZcJmsB4XgH1Rxf3Bb+2I4lJUd5Gb/vox900+eeH4F4Vw6bIClgMxeyY/ZRa0F5pm
zsDNVC0cBQqI9/p+C/uIaZxik8uF4Uzv28zmi8SFVzcBdxwhi6J2XRCFkIa/h/B1
c6UkvAulzXdssyWaYe6YGiXA/B0gYogz9Q3HWv1DlYaRRZfI4ig174rx3i2f9HmV
E4ezGHBcSYVprXZ+5T3J5eLtJ1R3QhNGWrDvJVfpO6GE08c/8XgBFaCRrSdYC94I
6LasdgSI76s0klrJvOds8rHLDL1CiIb8XBppVJydLos/k1fW5uK0fiXQL1U7cRbE
3ajK0H0v+n89dsjaRVXfOY6jbryQKb9PiqsuI4rUci7INddDJscYdYMC724glq2C
soj2ZoicrC2pdmf2Il8IZ8DiOm8nZmqYfqSYOgjm43uoIpkPFvcKlpsnpCdVog9A
r9i2dtf227R8cZh98V60Knwn4PcPSgHi0KOnXi25f2mUu+1Enfs+FyrnD6FepJ1f
61aEX1Vf5MdDjP1Oj6PN32Vdwf17OmbMVv4GNGOHoJc++H5hIHLEp48S2LJUOR/j
0FkyWmk1fEIhxJqwCWBhKbB2L+Q5Qc0zCjtwShGa460UCiGuwknrhvgswRGYf5co
96KJe7XWDIgybs9/zQ/QHRB4jFRWYayZFLs6ckWQtr7IqIl6UwSfZXcjSJDh6f3d
4N/IWcq4SZ9R5GAg8XFCpW/noYmwhqWqzhYplU9R4RTKGNlQld8WSu5hZI5M6m7U
zPROzBCNgS8ig0fVh7iDlB67p1KuCICHKp/mBqOHnxt0qkw0YwDFBK6ZnH8Of0js
2UWFvpl2FmcJnyU9oLhw1umMPSbWbs2FmzYVSJwM+zUtZyYnpEzNkNFSnibpOzxq
+f6oM6hFyMf7QZZM0/o9X3Tj3ir8hToG4L05xlqxOpT2gLuRn3mmEuGWU/4AfwYS
5wvSUxQ8nfcdKfgxCOtjH3qupLDsweU9yto3xT79IdHP0FI2UZSJTiEzpN3wQsti
fsziPUpvN4iLou70c07ItE1p2WUYv4IhGSN3yu1PveQMSLKbHg1FhmFfJsr8eEG1
vCv1w8R7PuZnQiODZ+GfgKqslplQvVbhUsSyjrGaMCSeuVXqV5+iErlEFXU9+lVg
WKwZPFaoV9LfBrcwrMlBwWcOIybNyzZKoNbWCHCDvB4U68A6H9jSciTMCurjNYJS
EhwZjvOM09cGYX3yXNiWhDHbO9GSJRFjAc6lMkPKJeIyFTT4GSarnOVRaHbTI7IZ
NGgXCdUsWrLVfrrIaZZY+gdggf3zMIOU6GX9WinET6RPwPfBEVT0dSlyzZpXOkzx
mT+0rFNIarNky43QgMBYtCytME1kr0hcux3l3H6rAGpnAKuo5L7eG556xKUQyA3P
T46sd7WT+brWgNMs1ah72QWJlEwYfbSv1TnUxl/ILllqQ1Une2tlhdJ0QtxkChTU
LuSSxiEkTiJz6JYe7fZy9JLCeZhPUdAgCygAW8DDlqxo4OFw/E5dl4L9h61drQur
9xYUwWeFHyZnVTSJ31Eiqfi5Cry1trXnV/Z90WZgTtzW/49/Z/lOc3gtRS77rj7u
4srLVmkMUZrg9Hjath7ClAMYuhVPtesvaWuyuNw01R+I8pHsspyB9i60Y+l4daMz
0FHUPu2FVUykxenQv/RglIjxt3r92qfvgAkb3IVloOee/6dXZYnvkb9lNflRqpV6
2taaa+bwB1exApBFVYC3r7t8wGbI+KKbo5W4ASoRQ2qC0Sp9k5ZKUlVV+fFh22NR
yjVd68wujHA7yPBKI5z/NSBDOeZ+0RMjJTCZ+WpPi5CrXlozhAj2zIbTuCtfD+JQ
ovWxGMGY8lsU7ADBwIQAeVyH05DubIT5U9Z156+6HtUw/TygG/Muauo+NNJTrykG
RK0YYcnsr6Mp86RzsMaCbTd+zIQkYbLHxTRQ8vAX9VdspZdkoP2uW58+ljHjuREz
bxlu6n64ek9ge4fsUFIz0T0obpaLr2dI4NsEmgAzaDIC7PxWXhMV6EFw525qkWYH
YJ/enLudQW+TVEboqVlUcdk7Uw3acgpX930ToGcyXbFV28dN4yXW1b2LFOXvFaep
twpFtzvSNW2nUqf/hi5isstrf0AQjHAFQQY8fGgAOjsah8w32JCHBQOX21PKzELN
zxPpxSNEyrpTckmBm4URCmiJZTf3DOU6/WZmWv1MBgm6ygqd568EPFTz4cBpTE03
SqxyQ0Ul1o4l3KvXcK2IlsbpwQDGKe2ltpP+hZ+VTYwcCWzLfNBJTRv4z3ql3x3e
6puqIolwI5g7wQGGh/29iaDSFKlf9aYkVVzMCbmj5t/41RPa3DRPxUfHT9pHgEZ8
3Z8AISYHneL1Tdas8U6I/xmlcfWxf8Qi/j0Y2nbPc0IQs4DQz5YCWxqpO0ABcrjU
wX0wchPv0mKkH7ioxUDtqpjrKoxMR0EFST+/hhHOoANWNpDo+CbAxOX3p18mlw8R
ypabEjjCeyd0NsRh1+jlrnzNWXyYB3FYWW5NT9RHHB0w6dUU3ByfEUj4yYZIFAxP
t/O1VczfJDuPmTB22smwVLyFjNEOzJ910/OCDGiPxajnC9+7X08LohLrEjSnY95l
Lb6Eu/HVxsq1eHhi7SSmkSlh7xEXbET9n5XciEua/kD3ziGF+KUOantKrjCMZxcL
005yx96AGEPhcz367fGPqMgKtEGB6sHjeeemEJeXB2Hm3LzXjUEqd4IUNG4irUkJ
I3lynBZBGso3qY9VJunMvY4ie0GweMeb6QgNByPAXlASeEiRVmjeEnN+EpujpGzy
c346lL5zgddyuxnZdku9SOr8E1o32YrQYS5F0nBDxXNTUpPZTmgb8tbFU+HiVJBb
tMLU+3dLpA80V1X0nRV8SWThIEv/Yt90kBAs/KcK/Dh8dviCVUxvkh2iwkb0//y+
gtqf8ZCf5/cdLrIqXty8pJFQ7+L+uLsYSl77gMvMQeNgqNYCdfnOZzMXV20Zh1fd
wo6Mvmr1Ag04ryrgBn4L7DilLLo4GVl/4+hj6ZIuIPxuDbyo1e/7/mshhAvb3yqv
RwWSa7d7MHwOGlv3F0qJqjndeXNR8Az/u7VaXBvcJsLOhmKHQCZEobqQ/kMfHKHN
jBe7LqMb26G+oBG3uxdZA4CDr10/5Uga2p9ycN4A60G5GsWnJzZOJwa9v4PelUq0
jzM1davZ5NH6OlVHjW2XI3tZStJH/X2dqDJ3SMu4BgzPd20v/6q4tdbbVXuwUwNM
85tnS1wnUX94v9u51m+QQeejWO/Ju/OHOC9uKV9Ze08dB383mF9TMAewabSsK/LD
sPENWP6b+uJC7pkfInPbu8OnhVI2JZVHIUCd2rpKMSmOsQfzsABKV9tqyjBxXtyS
L1Bhb2Z4cQSPuFBvF9ZVRld02kjvfHq2HUN/SCpO6JhL5LC4OZq8e5W1kD0DOf1U
poMSa4P8S0B/swW5fvkL8o06FnY9FE5NoCZt0CUGM0mHZGdGVok3NvzAPZFj3I+u
TIjm/iH+6YMkEOlGH3KpzBArL0DmZ1km6Tess/0k41ucThXy72qK4pnET7GdcxaR
KOfNJ1D1e50ZhlFmDbf+3dUpHAVASqGd7Xn1z5C3sDPfj2QJIJnYlUIho+gwzq6k
XwsXH6NMxUXZfBR0XTrwmVYUW/Tug8DGbjGd5ioOGsdCzPk718v/QGWt9bW1dBJn
uRmkyyc1KiMSdIC4uQ2ZAALGCXIC2W1vuOQOfze0zoJU8G18UiKylNfzKZh0tlTW
ic7wflceoY0CXk33PM4JVfu7rT76z6dmKugF+3zlbcx8Yomd5x5/2I+qWVWhrLYx
LtQV5Ocsq3d3klIesgHcW6a6D/Lln2Bqb1QxghjlO52V8TdRhYuzELbDfHrLpMaq
08K4V9+W+1/bcbucRDIb/rZzx6pH7GGFKPQiCIx3VfBlCd7p51PpDxSq0hCwnvRE
zR18AM5fsjGA8hwDVDpBul93j6yY3bKOlFSzLqPQxC5RHH0XovQ5UsJCIte5tOMh
FZfVsLbNGepjaDI9iXfTedRU3A6XMGx6cF4kVZ6fN4+1exKxh7xcT1c62fhSGwLI
FD3/uy+1uizWaJdUso25HHXP6y9/EsxxgMjasftWbpDOcY+0OwGyDNZz/pI6RcQ7
B0Jh3Nq/1pp0PmoTgGTCQzQC5a4sgBfpLt7sScgqfln1uPn/yIHpef+EfreWqHzI
rL2E5UcBqscPOHaUr6wLA4Q4eQAu/rVLoW9FJM+dgM7F0qFhiCdD/jvVrwEuvHoT
XW8l7OkacBIS6BwDTsRNr9EZuSUVNajGZHFGLvZCqiCz0shjK54Gdm3CJb9jEGsx
WoVk6EEA5TnkgO1Ee5QcczyCsb1cnsNMssRTZ/UcrzOzzr4Yweua/rLnfKxgGD06
UZy3eSTIkHyDcJ35eAHH9GSDPOHBMTuJZ4QtcJhAIADTUVrdlnreBxpt6j9lUCmd
gH2l4IOfsX/U4OoOozc6BkFVfLrWeGRb6zppA25X74VyhcoyGLrhcDAaDBMNdS0C
KrYMWKZ+FYr+VKw273z00tUr1AOgDyNpRIUalSNGAoNYoj1bYozbCvdX5/Lz26e0
qcANKaRdhfA0Qp9V3TcWMeYWP3Abh2vbNduaDy6TZ+M/ncVItuJuRXTYJjnoYV8u
8RxR5e1viBbIV8X3QS2WJV7V2xqNDJqTiPzhEfPPxU8E0DRZFkQtC75STivSzLSx
4Wl32Y84oek47ET1ejEvdzeLszgfDe5BMn0hHS/GU/VXne9L8nY+iw2qz0TZ0UY0
4mR1INPdQE9RaFuntgt24SLFbvyuPi+da5X3sB1UNROfI3kEqv7aDJILvJaDzys+
j1qz4EDNcHWziCRDdk3tSsWs98plpxciHwtKl1lcmhWDh21hZW8/wZPTn9G99VAU
LBE0ynZxxOVcQ6XB0crEewsf2jBTd62CdYr648IgxFfL1vtLWOZYIoFWnj2gRUOr
TLfHlGgO+I4wPSf0w5DlCqmWAxhWcX0HxAJx0vRE6F2iVNIlPwZq3n/R6aTbbDJm
fesCywGiq5SIRzPnGvvYHri1oj+cG6wGMhe/6VS8kZ62vv322Wt/HJcD92x5whR6
QXi2KLTb2dnuReHuyLsIq0yxPuXO2hWATn5ec4k95s8VomazfGDOUPHr6D2z5BNG
NYg6YqldQSqyflc6VuX17T6Pu/juL1oh9c7voTI1R9RHHqHJwbfNvTnupNlYHbbd
ZjOgHiio0/efU6XN9/c7uXnM3JE5eFlexluGjaUT3+C3vVtotzy9uwNsJbeq/MFz
vXaMvHyXCzkxXb7MO4m94HiOS7CFqVchowtXlLF3iePXy3AzVBJAWbl9jHa6/q6B
qhA4amGEslDldxfeisICGnnOwN9b20S908oCAB8a4Wlu2VpS4bpgvwnuuRdbQmC+
zXvRpcTuG88THcvb3il4XeqUAKVqNvFRm8lYdYNb07kbx/r4n9ZrEvHjUpSl6L12
IUEnC13/q8AsHiz3Ohfzl4muXJSAcO+c1hs4KUlf3jmyzewBO96K0RMjeq/pPKuh
AWTU6WVsBvshJjez9T0yySKw499PNkcULeDzmzaIRwGIbs1VZDKABmbgLmhLgRBZ
6aP6sb40YqYmNrbPS+3ZNlHXh1WWNq3Ymioosh+MPszNXt6jzOLaqdNcayQh7TVG
d504VSnRuAfswXm8ykWRX6mR21lrvOf/Oa1fkxQ8H9OL9v6HbBMGPCgNwn4u9ODc
rOS0PQzvaYbFVcew3UyJh7YmetOjnzmb6zWl06dpQ/kv+ls9shbT8Mh83Z2y/Bx8
d+HaxdgX0ll1lvH0dB2/O43szOlCi/uyd12Kz1RQj0IyDDQSlkGL4NkqcOtEtbrs
8TzCj8p6QVbUsGsumjaUhTrLXd8oidMeYE8TJFD6u1SkcJ357475LQAeMYnu4O3G
p8dOU2posxCK3ui7L1wU7kP1luoM4dDC3rwRwYukbW+RGVlEJ0EsJxu6Pou1k+6z
KXEeU4xfMQVgYQb8mYDPWzUQJBGweRZfLrjzTm1FkXZz163NxNUffJQw89uPmiM0
R9hjedtac6hghvUpVHIFOJ1evcSJ7+Hb3+aWUSTcXoVtHuzit1/PecuppSIVAMmA
U/h7m9ODXa7h/IGQ2rbyk1JrgFn5ekG5DvMbs7cfrxaOjGzUMQMUbKKBpdNR9GXN
jm0Ic89zusSJYvZim/X2rTFlzgtCc9ejp0tLAS4E8C4rYRr7wTMypTVpa7tzKqMe
G1IESGQb0fj9m+ANE1WqpBqGGsILKafQ1ggJKsuIaMOs/0SBokW09a+Kn9Wp3O9s
kiG6agJXqVQWVl3rVfA2PVOUpr3/JYmUxjsGvPu6rdOhPc2/gfOOZC1dwCGcp2p4
B0m7WhuP2hu+kx16QtDUYR6LlIawlN0Cu5cb5hv8GBoH6oB7tjdCk9v2MUmXXy4N
PYx+LgpaAlIpESYCp83oTn8MPu8ROozTG0jaXf3WexrxEQ157o03RKULyZpBCEBR
zo99KZ7aYLb9e7nbRxF5aHLBxz6FwN27KzlHJIM+Z9vhgRMAm+qybjMYg4a7wywj
kgG48tihdqml6wrv1EBHLDEeOrU8yopz5UJVV/eXyPLoBg/ddORi68JBYP3daV4V
4InHNNCzGLGg8ODYrn3gLCusMF4rrhqgPXan9kHG4eMEeNPNVUfNSrRxbP2mPe89
MYgGlbEWhJMwJHfwwTHeK7iZNsN9ZfVnfq27EuNskovydHHbyjwMs0J/JJ8BwzB4
U5WGKQ8F174GexZJNKMGIZLQ3SNh/xHVlebnBwT0Feo+EMLxf4NYYWH3HHzGRg0e
4wMd/XRNNX0a1S9Ucw8PXUcvKSgbgX5Rk6rbu/aSL5lh1LrW4y13eoHyU+6QLaNV
wWAvUhtnNUZxIMX0pWmUqLew5Cth3tJh1pDBwTyLErLM2I0X4UMhEYXFtpKrs7uu
35CQiTr75/kp4pmQ3bpY0AO8Srsq2kPJ+fKgikHcYehs4JVuOQosNN7sxZ73mRh1
u0GM8o+3UVpQOlO0uJWTzA3mlgIJjsXSKr7RRUUIBDk2dgpfqFfY/7jeuRTPwsuz
4mUv7cv/x3oEef82ulkh4OipPmH3OoAjLvGA/OL3dBmFCrgXLzcQY5+Ns0MCsyc3
UQuLuGFUbbEfAAwFv4aoh4Uc4Zlj1CHsMN7b0JcMDJQ5DfgSegrLlMNiLBdqYtAs
mKAUv9T7OkYh3lTKfNeTYwYSZZ9qPZn0/9/2RDHU42h8vFf5nTFAb8YtWt7WQvxK
F5hyZNklx3Q3E/7dlfpmVTI+zWUAm+bKmqgKBPRQO/JK7DryYr8/GRZA5lKvO3Ub
jyi8pcqqaW/LrXnyR6Rx+gu6ZFHhPXzsryxPM0+ZaR/LeuZRDfipm8YhOPNR11R0
7LDEpkEI4SKJBs+tGsNZde71B6Eso30NJr4Wl8ZlVNuxv7nWD35S1nYpfW32EhAP
mNYiUC/dR78FnR8NBCiUgw18ryscKO51rDprz6BB+9GQ3F09N40Dj1EtSLlC+zOQ
7ePXE6MzJzIi8itSO+4oo5CxCbg6VuMheAG5kmOihRwDoKNqMQTtfhV+N65KxJrZ
K07F5j0cAR5nx/A/3Ut6+gJy0c7hfG4ZtFL+I0IPzmzR+iwYc9RtibH1E5pq+EBE
8JmWbkv6395oxhU60K2pOi1F4GGbrmuJo5Ni1taUGB6arpLEq6l7V5LUmboAWedx
S1IWffipnU+WnOLz1wlgG3/ZS6zOtZJTI9C1LrlDk9By5Tl0+MHwNj1OSG27nEX3
MYkJOA7UJPUbIzykWUY+olYUCZKEo4wGq4G40q15yzLPCDBLKwiA21X4oVlMR5Wy
9Zyr34BMZorvWFs5iiUxh/xHobV5A4eO6vwuBW15VIeb+1MSSb+c3scRC62A5o5S
9QAnHW0Xior+zdJ4DCcvrLg+foCKV5tusShIrWLrYW/74bt9yvZo6MrzwAe8fcp/
Gyx7C9h69wvWqAKLLOQpzBle0nfh34UxSyYzzJNBlZ9yE7guKYxT3r4ZKUU6zeAp
ognOo+EJRDxJXmzZY6PDOUVXkZWI9MF9fLEkY/g0nTLsbRLuDP5qVPBUCKK0sA/r
qOZesbfZ00CRf3Spluc4P3dPMC/zsyHBAyYiUHGpFh/+eGfqZAdQRLYXlJjtSstI
MuevD/eJsYgaHLU1z8ziLqstkL9zyPuQycIfjwEZSGZf87zqj1tw3q9ofqXVuwlV
9RT4R9kWIYqsgfC9w0GyyrVsyNFMExW7wPc0ali0BDGt9GP8LjSOQQQrckpqxKYa
y1E3d213bhYeHEsh5fkIMbERXCRltky7Wr3dpEz5T9mp1qR6gpvI8J3RltMLLk9X
keF3B6BA+OthcxnzcIbpyfLuAwFdFCrgv11Ou9bgGacUl+VDzJP2Ee5ltedLeaJt
WLn0baizuGIIPG+OpGgVB6OMIFZc53l64FDCyRf4Cm2tY0y+bGgZZTm3WAho3VJy
a6obHINW8G57ATPWoL209VguKrg1VvXGfTQOLAdeg2brpkNzqZ5XBXROvCF/wcG7
ONTvd8LVZKX1oUmn7h0z1ANOz/zG0f5R2xys+OGhLR40eGGESnU3qNHp0+LaSruq
lxCs7tF+LHuK37hLI0IYOfNolI+9wFWxlyprUH9Tuer0OPX0ryZBtmzS6qYx1Lgu
hKBK5T36HOZysnvI0Cym+8OonVo4q9WApd5jCKZy0Xsj4vYffuNxOqXhoFvFi/KS
Ch5omBz1Z26l8CYWQNTP3qcvgtqDFLAIVVUJ7lVV+3B0SOBNvIWSy1IcJguyRjXU
5KrRzpnp0ODyMNsMtXEjBbakBEiWPKkHAsBCcD4dlkM0ykapvd0DQDrfYJELk8fA
TvHcq3spvvflGVaK/3bNL5cSZUu8hiNz6eucf9GG9UIMJXxys8vg7B4MJvaZUyWa
LEB4O2qmn3K2vnc4rEN39ZQaUSxC6rSF7a0GjS313uW/b9arTZ6wFxKF5w5OD6ap
fx6PlJIwREcLqIBxtJhlanW+wO4GnFboR7Z1rBZ71IvEDIJM1JvrQhwiTLnZOuH+
818m8jdV4GzjJCLWcgky+HohmdN8FSbWs3L4PhnbsZazqbVXWHDJiKrKyXf/n4Dc
FyhBsQJRSEc83LfOtENSN+TPe4qpgoBiy3/rxXITnjYd3VGHJzN83et4bzb53Dnb
zd4k5yq5OOyU79WL2d85KGjnmnZE9Fa6l/79en9hAK5lkCf0eHvVU1q1ZqiquPJY
O0up5xSmOOw6ypjFlLVSTB1aTapV0e6k/qGGfVrUPG0hbSKBogCGdnlyMNM/VTOx
5f+0Viw7mlart7tSp3gbEqSKEtCYeFUXAu14AnWz0KtJIMWKVz3px8EjGfPW50Ej
ZDSysn0KEe8NR87ogYYxKjGlnD8RBGWGzGfJH/WmULHzjkGVNjGdP5rxl26zZBIV
dfj2FNaQuhUWZZGyeD2rAkiXUULhUM00nxNfbtaT+XgBGrTcn3CUdr+0ItS8MpOK
1IyTtUjHKC8cAry37WLfTSDGQ3CFDrZYBwHitAqsEg1G72iOIfTeo6LSCZ2P64SV
H1YM4c5xIUA9OilnJ4fmeE8jsnp6E4c/PA7BHX+39BfhkxLSAuzRv4tI+WK5BVIU
uEKBedg/Bswvjast+Ke6a8o7ImXBUYyu2G2VxtGdreH/mkSXhFBdb7Vk4kDbZB0/
EswUlFE5Rw/Q5zQVQ6H970sVmS2JLmuEUnz+NP64xuRF1aUzkWkkt6TnRAcWIzdm
NiHoutcBbbfOJUFI+lu1bt+N556vxzqSFwINWpzx762E44ER64utewZVQtp6UlQ8
e43QMgaQJ0PT8ZRVDs/UaP97e36LeNPMoN8SzhBDFaa9fRBz1I2OUOF0FmGum0Lc
ddm1urnfVDJMbgt9VIp+kMzdl8ybchTSWei4x9//9imrhcvqAI60pCDMRUoofgUC
uU4BYsBzgKriJXdnTd2/RTh8pnyqXcQRMyFOMi3pNNO60RbFFpejcnsmuNHVyBnM
QEphgIYxQzTVXpx2HWX8wN45aifC5L0KW1vFSQrcjIdSfbmPe9Nu5u+RpJEwvpXp
vi7H+WcYpi6prr8u1f+9SxveSNABDX0uvY191H12TNU7SL2FfXkpOtUtM2eSBa0G
0GFvUBUIoyVP41sQ+rBLkDYMe113n8t3nZ8c5kHP85JcqfG7E+CBsKjJGxznaXpb
vKoEOPwkXrGHSrCTPE8uVU2+W6cB6qEhlE8pWmUKfBLX9qRdgxsLvI5i7fsugFrn
iCwzoiBsIZhZHNds+rwCUxpSEJgGTqGDJ3ot+rar/3KwRT3sZpTHdR9K7b4z7n1b
V6IWOtKfQGbdy7wBMQ5RbY1TPDhIzCSi08APXy8xe9pF9DE8vzt4/dDJJh9uP8oN
ivwtR6SvI3j3/WKGD31D2h68+HSxp4Q4VjDVculRjtk0QvZQ44gMTVcj3WqR0MoM
jpv201PYAcMmrq5GG36DoE4JFivzT2dTExX2362FWUitZJuvwFzn7mSfQXmd58XG
pz/VnxhoV55cDGtiAhIbg1feF5/Q6Y/cdCyM2rQtUVaCCRojAOodFBE2wEkbf4lh
T02/S/TNDQlvL0b/uI6Jqz/zB6QrkKve2LQUupUtoOoVTvYLO7QW8Z3Oxr70LJ1b
2+DicORY/UASyLuUBsuaNqfwM3Rfc5NXjT7wsWKaPIRHN7dybQ0UD2X9HbaO6/1m
YBkrSZgEwQiTNofqdEuapln0wkrJ5Nf/k5FBDxTXy6Xv7ble64N4C12vj7gTH9Qd
Of1Z+QiKFKhqXbxqapAhkmswlh7NQx1P33KVIEugSgImTDV6LDk3fvGaf1eI/mw6
CjNkEbq/DX/czdkkSg/Zo2EVD3RraNq0vXSfUEzQpyzNXYHoMIBWUoNMfCRBhiq9
Z3qtchtPiVMrjJjeI8Z1uAPxEjNTe1Q/YeOm8BKy1gcmYg8zLz+rO45NTOgPIxO/
H7oEvybYVy621gms0a/Zx7YDawDyQT9BWRKTC0Uv3VEdRYqHSl7VjZYHG0QjEv67
iLeXemQTJ5X5C5Rt8apO5qUalw6xZ408nLB768wnVOxO3+jS0gHBHfDb4CYN5fac
EWifqb7nSVqdBLqtCA8D9ldk9tSF1OP9tZ8Y4U11ZDh2hsOZk4Los4OEc3u0Ntqu
mOB531MOBdOGiKJWCMR/rey5CkENyyI2ThXHl8OzAG5mmHgrzJIaPGI0knsCxnsI
S0M5FVPaK7vBkWtRP08bz4LzW8BwRDCWukJMCq/QPZiY52N6g4OCdhQULrIl3RDP
FQDpEUssGmx04jLbXve3kqxHFQXwsl1yYgW628bTo80G9Z7290Bv4hOjd8GTOUrF
cfjt2FrsHPyr7wRb0MhP7Qog35A1SchobbdYLmUZfOO0mT1cyx2GF1p+97/DKD7X
FL5ph84zG8EuwAwuYh6Hkgyqu8X4lzYLgHnyTYcL2PQ/d9uYLfxZFYi6EHPogTYR
SNmcfaBvlXHiFt7FvfDymRRy7Kp9+NIi3hahBOEVFuNvbj5xrFOy8kVTOSPUnOu8
oDqEi7AFXdy4FZDhjkxxT6+rQNih87e4G23HYID8AGHwjqHFuwXlQqw7OsX1y/Nc
7s18vVrV5zzvTt1ZD9BcuhNKCDsA2Pv5MjAstw4bpzD1iNoAF6c16VrxKkpdRb/i
y4EhtRMLMQcIhlYo2HPEtrcSNNRp9gzSeTYIt8465U0MH8npXOSHzoGgo/kQ1jcb
WOKrswV8Zexqbdz+P+9jhnE6tcxYIu0BQc3/ADt/zQ0MfAa+qyAqTTXjw5PeB3/W
y1UC9sy9pjAHzTUBwuAjh2HdnorbR1yIOtgWnNMpdASl9hrwhZhMCnxRC+RYfoQl
REvZCM7bI63nt3xKtwfiPPsq7c1ZvpGk6Je+D1b99U7bbNisuEtqJfbvaTHTGHiU
6CU6WdgfqiXklHCsINTR+16N17TbBbkB0oUveKTJMddjB0SiV6eAO/mqPJW8gZzT
WRk/7tsloBmfD/O6UbUjBdGNHKoTt8kgoZln+IGOQQIdbgnOmaj5+fJWX0ZgshQH
tikZ5Q/T+6ajhWFwV/P2DZYhjRxjnd/MncoicDRMEmKT13SyTc4vwc1rxfQZw3My
CVm74phnGyUtJvZ2jkSyyXv0KsbWTkHAFUtWw1i8RXhJ/UyyVJplHKnUOHff9a+E
adP3D9nuPPx4/KRP3Q44DMpqeEbPUnlYPevRveEAwtrrEirh1HnayHVUmK1bUCLd
wz3bXdF5sxKFVPnKpVlWaCFCjW5Or+aGWn1yIPKDa8tF/H5+l5yjlNBTYfeOfGMK
43ohK5tOAoYg+GXZsDhZ7X1kHWUl9MUcq9hMd0XDysJU1/GU+KpK4PcOkxKVRiQj
xa5Mm4bZzclMtwdgjOLSphcAOrj+COufQcraBRZtAAxrRt8ZrYz5P8BFfuVt1W5L
Of3lPFYFMxQlCUjOgsBDgBVKK/kUTo8BXrb2tskp7Q1Nz8zCyW8pENpFlnLtLgVb
BqCDdzb5jgK0y393luXJ5dVWCtE1hcpljx6vyxrGtfGGYF0CahurNbpOsEeqXZl0
6EEam4UjlILf7I5TTSJQo2gPw/2SzqFsSdli902+1nRj5HVyRB8cINDc8VsTP0Gc
/PyaRyTVi5VDTfsrX3x9QrlWG0YA+RwIvU6jwbgJjsMiLMhSi7OkPjtYCkoBIeBV
LGos0Y8nWiLf7NQxKCaAniT/Sl4dOTV3qfJMhG2aV8Dn9wOGOt0Th0wmYK8ElZTR
hOk4gf+JNQMvB73MGlZ163BgSLEIQWvIHs56PHn7hkBQVODsHPxB72OCZHfFhQmq
jt1A1KxafGb+fQ9SMItrtDPZsYU1UjBTF9vFbANj91d0kgJAhIkPxU25J66pXEH8
IdGUO4ejmTC+L15G0H5xVgoucKFxI60A3R2Jz+w67/tM3qe0jwjSLetDbxuzKj/v
9ddPBdJ6CHLCw0xKWFqptpevBzQYmGpWNVzAzrIwlupHWdNnH97og1Vv+ZM0PeWM
PfG7/EulE2G5Zk7XUhQAcymJZxjm7iBl1yRacmOq6502Hq/4cnT9wgDJP435Nqy+
ID260tpV3k8gVDg8Hjls1kb6BIBYkCCs6JlX48ahW1i7Hq1XeM/IhQbfjr8NdrdD
/np4ZOWpR/Eyq2b68OTHalk0C+XyK+ConxNpvMpij7plvMtTPx0gHx0//iSDJuve
lFfmJUWFcZ7+JxACByipega1pz377/sViDs7nJKSoxKXABXbFTgikFbw1bKx7vJM
5m9hSmfmODrmEAav8aI8Jk2vXi5PbSVEONpq+ZNZvToKiwC4V/eNjLcADyzzhZQ3
RrLL33dpIZT8V8gAu9MYkv4HgCmsTqDcE+H3WSD+7GcQSSSfAAW/UH/ayhQX54Wb
kVvVeZHVY0cejKgeLMZwr7D8UDNc+VBr7g3nweh6u1sy6KzgKjN3LIFPHNJvkxaR
1dzljhpx5pmfymen37Km9f7ozZaYJN4wfM/Tmf6p/dieDlmYJyBcPIILygZt0Uzu
DC4tV5vBjAQ+5BTxPp2JyD00gLT5E/aE6NuHRPi1kFqEltJLxK/Ngd+DY9NZRdWK
Ig3DrJ0u9zystcc6Fmb5jimmjGsxuRU7K+jC5o06xu+oVUdFCpxvM2/6JgW+vkG0
+wr333+cVB1OlwVt7ikdWJJyIfx3o2PiH5rT6tPP/qwa5daV0B/Ifi5anCDH+rzm
RNibHZzduzMevE2eBLpIzuoUGIroUOA4hzW74oM9aDwjLixZo2lF3mJOsYpK94+R
vwM6W76EuhnbybXZ7XEPu1Kwq5fFNxD5LJgPHF0fYTTYClLxaduehiXtg/7KAsup
Kd322RTvS4sHjaNS/xsoTWBTP33ysPFbcrtjo0dntLA0pRQT5j62m12SkSqycqDR
rLaYVU67vcMoQX1WR3fIWj9w8Niv2pgQorIUiVeV5+nuZDu6LycdXbk5rtSw+4y/
C9CSDxTk5MZTo+1ISd4C9k3h8/xIYXMd4CrioeAAr/oV9nhfsKwy1hVXLrbMYvuc
WJxMcrmGm7ETQG7+Pfkt2lmX7Y/6qenencZTcOjV3VClJRMkftBEEuFUsbN6x2KC
rHNzrQeU6wafaMQvuQpWpdU8Q6qjiW6D/qCPhZAnxDrkMsrZz/JUpxnD67JaDK1E
pNSU4VFUT3zxVpkrt0CWpi/wmWyhS4KsmsROY5Mde4HZhMRpeoVv9EnKleMPfU0G
A+qJIETlk44NRsHUO60/MKhEt40Yslb1zWooWqPlt4ZOpVJZX8pGxp+1hRcYtfw+
GwrgkfoDwfh4tO+zI+exIDtL7cw/ub17qSOpaCcoYGq7iPEX30+1HF7GZZ99BY44
tGPKIJcSXEDxonY1uJR0yNYiQa/7uFiJ1s354VAHd5XLon6+AZctxRAxO3vNImUp
WM96TdtUOYn/+sUAoalv++9KkkNvtZ8Y8kcNfjKI9FYo90nKLkVX5WIKWrPQveXM
nkD6lxrknd8YceNVsKPW8bP62MMqSTtafdzSSwAJx3qfyTmzMeZHvrdV3tpocySP
GGVI79+QfbAEFyGq8kYstlOWOECYXx8HbJM6at1eF/bpPnP1C3lVJI2iMA00i8nW
/F2FxS7GIZEdOgmmH4vN+kqb/btF7oKdUEIu8VBlQTCdNaR/WPQ5rbbNGjXmlVK4
fPxWIQ7N3gKjrj4N6jtt/EbFuNav8GJswpcRONiT+7nw9YbbumQSUWe/SZX/hygZ
eWKLD0HAw6+PpzwBdiLnMyUyEhdNw0MQna/qohyjwKr3rPhw+RKx68DJu7BC2kwO
0T8PH5X/5opT5qdE2KrfjESHgpVZOIaR/I9szsm6zARFE34tLcMctWPHCTcighxC
hFv4rsElTQDAnqgFFWWm9yBuZdOugnSAtbdbzyh6/fHf/OK8fb5W4YOGKd0lSg59
9K9iXlgcS09gqq/ndcnTUQuPfpH8wFwaQlXmWzv/d4vGuh3fyiNcALmPAt/8lAWX
9EdkvkyiPh85c6Ftw0a8hUVUDytVZTk5TQxROCOlXRHSuaoA+eu4b96gSYutDqhn
gqXa8ulQ/VpuF1Wq15qxCi0F0vaHxrr7b+gj1NZXDcfYJ2YSq4qGBnODyPGI831U
E12a1e0Q1TW6V1dVdo/d9z0SgDRCUa1U71vGgxO91xgn2iY1cufZAYRJZQ041bNK
XJqgdgopMYA0HYyAcK8sFZIpb1SN2byK7N9N/3nWXpoIyqmcGn83uhc1oeW0vZCu
bpasa2ppX2QW757+wQYOC5SkAjCDhSZlopbD6dJwajilaOmMpPrsnMk3qGD76z5Q
lQVDpzppeClWpvAp4M5DVhngVDN6KoDoFN/qWQ3XsvXectk0brfHiZesu2RPPwO5
zxRxtO85pLjA12rkuGfQfid1Wx7xtzFaTfPB++tQwDvrhQebdNfVCSwZt1boMSKD
Wh+NMG9mfoHRDVUE6M+qyk5o0rZGYUVM3BjLhO2/w546YEPy8RMFx6KWtaJc/BZU
LkwgaRC/wOODOb8Pspf8u9ga9XqzKHe51YCibDN3bNbBcRoKYXuCO+i+BmI4VaQo
GbnkmSOC1UQltPYGon5a8EXafNjTfX8bsA7jilrhskWK7AL04kNSWYDPyU/e9+Cn
yA+QY5bakMvh89okf/NkBGD2npgLvp5COT57JVGDm1x8+E1rosAP2SkGiAZseh58
ZRjkYKftJ6ieWpXzp5fV5UY7178kA81W84AUaNONAkNn6eEE8JYg6j2FPMGR6Wlm
0QzYJqJDoVV5aGAN63QgQ+VaJMouThZTgHb9gZQTbbaDmK68wvJaDkCVn4wqXA5C
8vC0Pt47pfjrrWckVhcmYpC0PYzL+AkSCf0Az4n2MO5N1lU6CKjVuM60L4hn+AyA
HAMipGOBHkBB2ZT765jtZD5pjC+SFH4t830egw99vLyd+6aKS0nJ+uUFDGiujl2k
DiB76COSxciG6Zpsel6LYTwyq5qkn40wJaG7N/KQ+njlXKvIZivNRIi5H+9sq7na
wA3eDlJMlWnmUAiItmSAMiInRS6Hn8/0w4Hkq9Hq++7ogyKZ4KTuljsa1SkuuDZw
/IkyYkSsYz5UhloZJMsvoUD5H/HKqVV1Ywsx4ouQgdCSV/TRUvFTqVjuJ+uWmDlr
uDuHGTbbUYGOIr+IyInXMsYn09QaOqdAndtK5+dps9aGleXWthM3Of1eWPnwnKSK
VB84tNXzR/nfU0d2onMmIGcxfFvjy1siBCc4LKk5GUBwIfq43sfOLnJOCZ5ykuCV
f96izvLjlwRZRVWEHTcpREyLSJxR6TbrrzJQcgWYOSQsEBL7iEORwnCOcxOvHqNy
J4kdu5Jl5xpNpn7v6lv2DrqAQkrjBExq1aEAaRLcjs44Q0IcXcupriobl9wDMAbT
0jSey33WDrA+/UTkez3JSyEmPwVnudcX7xxHS1JjlezOqzaLBeb4XSl6JPhXoBkJ
9C3uvj62p0X4cfExN11nUsYwu+r1G4CkGNBJCt6bXsxuqTYkk3gzeWy8ofxSkzUe
Lz2Lm4ClBQBAt4pU+uL+rAJhkuGi35bqhZ/RegejKksk9HQa20wK5Zz06poGNIer
OskQbSa897aYAm67lvZ6pmQ741FtXtm8lgWKUgJyvAfGApwJGZgzKeg5HqbWU6Dp
RuC7aYo+hoPDcPf5ZuG0lBJuTE5p23i3SMqsWkPGwoDIe1B5ZOaiUWFLeYRW58qw
/Sx5lJBJ1fAiBp97eL4jTq2jiVBzjmxY26Jt+ageOxxc1HWQVVKYg5h5JqDFQAfU
UKYVhHI7A6tLoK13FfmuELQxl9KkYz3L9AAehYAUYMT7ApanJ+ru7YARJX0c1NDu
hGGLl1NpfnsuuUVqVe5d2BUEMyg2R5nvTwEQZjaip5EZKatHqJ7ix2JRUdkJFltC
+gUBo02XYtIaaze/NWzP3AU64Xpu070QsxFLGHetUdB7UQUHgBMMqGFBQcdJ1qO/
Zf42Sa4ZdCvRsJkfUycGSImi9/M9UrmaQ06x77CXalcUBlDk4Jhxk0Vzmh7o1T+o
Iq3O5yYBjS5U2nTqQOtc4bAn94Awo7icZ31fAo68wvbWCM/gKIkbAz+9YXZrK5P5
VQUr7uB09Zuv/THsJ4gY7JiMzzsLbN7X6zdD1hNcGblndqaUJdHoqNB5AjAtA3k2
Sh1H22Fw60Qf+wKf94pGjYFkXyxWMuVtcl8paD3lYW0XGQ4B5y1b8C91QNjgrBwT
POcZVG7QHMm1J7XZ5YGOOFRH3dlgVcueYoFWbfsE/YrDTkBl9AVF2NEbZZp0749S
uRAYFdNjjAfYJCApafzy3zTk+ZZ26YTfqgal4Mr8o3H6kEBHp4qbVRyMWB7jL1Oa
UnvWhGjuZjy/Fv55A5C9wA3S2AE5lSfMXbkCvwgthgmE1MYHcxSPWF9t7b7+Rhdg
XlzTBgAFC11itLyaN+9htgGqD5SRP0uVg/yWs7fkxeD7g+Or8Lz4D2CUfz3WX0ZU
J+Km3hGC3RGYSxOa+dP1nMZcXESjTGuskIXdXrwAhE7/aK5/ZK5KmoUxKxau//2y
hJmVqInqph5aIXcv1ICcUXVzQknDAUcZ+5rIpwJN6Hz7vhw8aOmgj3DYZLMelWw+
5gADLjuFUQkFpumLhKoaZkaXYI2UZjseB75k+nbJ4uT6bc1Xvn8V0hrvT49rz7lR
CLvJA4/hKSCqUUjU+scAv9fW3caybKZ3WJiiGxt61OwcWv+MZgIe+W7r6GNEgV5l
pGMK2reGVUwPy46cwVOuGhsG+3bU14hzjFpMOXvnlwdVaiyrCSdrsUiCudT677v+
9RoRs+q0FjPXyeyqP1ZwOmlbApDjeMuXSmhnLwmJlNWsAvJneUVGfRyX6ipSVFdh
7EAiUdKnglLtgTauoSndhMjvpRa7iYsbmwcpFPKXbZlAmjoGdSHB5ckKgX8qa7ZQ
mtn6AQPxc37e2EtGdXZxElot49MP1mzpgbx3m52WezFJVpYi+IsSbNYCUc/IZUvI
n+MHbtpt+ThRhpUISNogeMiRshZ1tXLxNAKJRkyyXYOnu8gK4d78zNOFQwdyKv76
7kn/SYpKL24pU4GPD3TwL660nzl+R5mQRicZ9pnilQseZE7fw8JkI6Unq4/ikd17
6YoytYadcuRhm0obzJv2TiJh0XVKx3Y3XhzY2An42pW1B0HEN9J9JTX1gt9GfG1q
Az34iquofpOkcxSFV7a30Dz2Yl8Sw5M8rvZuYiFQ+UzFMh4HBuZ47Z/O9uIWDqYd
cigUlzCh2R3EB35meN/GhSWTFlHRKQ5l2BY1RXFUPUQLLqcLf5G54cB78i5iI7YF
svm5bCx8Bg2nwOb8hisrR1ykjeV6J6I0EG4sR7hnmPVq8Z/K2Oqv+iWmZEmDOf2/
aCXTkSrLekpy4HrroBJ3LnrvFLTAOn6JQ6tigMfwEjkz8q5zj9QH4RgRj3ifOFZj
dh2AI4OciGyUgZq0pZjcKNknmhCZKYLlRowwD9p60o5wEz5QRadRnJrpWNRRKBIK
Dj5DZW40OHnkd3xmjV+4yXqVcxniuYVliEfwUY0JKLP5hjBs7xsKjsbm9v94Yxjt
duxsZtILPjo+5sqNoaqILmwRqVFcxCoBSQOncjHv9dk2xPfpSWIq7EBYY6PAlv7h
ReE3ODz5ZmYQOOPDy7nI0RvAB0fA3C4q0NlnLEVzjWzubAtouye3uunTrql8Qjm9
CIzFygc7Dku7hUeWbqGe2Jf+5osvnG2DUw3sz4WkiUbPOSM6GxdldNGy1CXYp+mf
i1vB/nmoD2XNni2zzwPu3Uz5ZrNjlyJhB+IGKTa6qNrG/gsUIqIYwfx5Y7Mb9RPR
EwugQ8Y+2pxiZcsnTQES5kxzwvxNePB/C2RSLi3U6EqMs9dMpnndAcwL3MOBwuF3
Y0cUMoOJErA1yQ/Fh37OnRxsxdJxJnSrkKIU5tRQi/bNrgwzH9dz0BouPklSXT4C
Pl2XG3ZUbizf25CjYVpijMC7TzXhPROwhi67KnR/DdwUydAQAGlaPaFHB5Q/FCGE
No2bQo2Y7grqQ+THj84U7EYheamAOeoifZOQW+2avUmixKZ6Yb9UE6R1PLPa2rvp
Z6wqGIULQ/PnB3rjecItPVeotcmQUrTMEPk0KSqu3iSHT0WA+RmoPn3hj+b59g5L
M0IVqKq/0sgiGnBuC2tFCdCsBtLwfumQoVxePBvrKIqkd8xqSafYTTENKPdbxQmW
tfVzyX+f/7pjkeBXOsFwUVucC/6VMI9sDlikijP0Y2FWvtN8OgdFllQpswF0FYVW
aZsU2nfKsC8zSQhZ2vaNmPifXtA/QZgt+tl+LGHdgdMHRhGiOVOr6i0o/6nauS2G
UOi6jYH4GpwR/uhx7uxeoLd1l9nXHAMoeBBs57JpeZWVd8FZR6ZDqUW0cWIFvBuj
hdYhoEi8VXjlsrwGYI2DBt+/JLEbO7Kl6q8kDIJat4iqdh5MGv/3i6yaHyzr/LWg
AckTnDrN17XdTOpDa7IdVIW4gwbVdCidF3nKGnXSyZ1UmmAFFBZmKdigMNCitWc5
3yVq7VIeU0hsod84aBAmYoAcnxcezsoCJjci9a8pmSdLOTFetP1hJFs6bBqFYTTP
t/L8OyRI3ogJ9hES+UT7OBh+UyUmUbEehDqJKhukUArp7KIzcvJabNXKpY9lKDBl
aTkbZozY3wSUQ6nJ+/Wc4jyxA1GMX56MEUJqRpdDLNSZ7qZye2eYzth56KhorPM8
DDklZqQ+NQ55CY5bjFWLo64s1LSpao8ZcdEtHkJuTP6keRUa0qs6IwSs9PgeSziM
jlnRfN/6do8AIPTmIy44WNFRLhjJcgyUYKeMjfrKkhk6h+egBIGuqqHLg2UNpscg
Cte1bV55frlMSJegRhqZXTmZOpbw/at4YoBBomt5hkK9EQndlnOmNL+3qpW2+QUJ
RbWGgtm2SZ1b826HCDE8YpgdDSXNbO/x3LJBvjRPUB98xA5QoJA4JN48/5gjgdX4
T5DA01xAoOoQ3/LXbZ5ENeqAxVhHE1vflJ6Mxxai5smVj+j2hRsz1uPWLufdUjB2
ZplJuZsEh05Cr6SUEmdYm1DMHtm0PtH3Us79mgoqd528FF/lWrCiKO7Yv8B4aHm4
/UEh0CiqSbhA+Zcu8HAeLlbDczkMqaxk0Rnm3PuwA95pLY3emXkmimJR8YQw4dkb
WW1Ag7plYtKPNS7ItcMFow1SSQiSO00e1vxknYYLY+bMCf4jZ35Au1OjJ8oWH53O
SlLZrkL1hsIVSomEGmtDbK4Au8K3f+eP5Ty4O6FAtX0XzDQnJ4IOVzp/9GblUUeL
Zwjv0/TofQvF1Xz9JJuAUtv8ZZnJjKw7uU7h+rOqRfsRs5cmrpQ279Bm/ZEwwZYn
2AafujX0KHRl4Of6SE3I9IymGH1y4BXw6pOkJJyJeIsM1cSQrVaIZTTX57hmPolp
isI6a9ZndJc4DbGYqUWZG3PY1cZ9HV0dLoqjZhqf9xs9P5jj1kFIE2ggjm3hoo6v
7Og5+1a2GYFNHgUG/f1hoxnG2P7236G+kXqQrJlnglQDkWLp/kah5qtOgAqxw1kj
Ef1YHxHE4xW9txkKpLs3nVarOtZqT3SkhaiLbGCrGG+PUUemFYOsl0n3tY+zrhHC
nhAtYhyx+kuHzRC539nN4jn4VcASakyPGAIaZPLqE5UmpVA/bmixUrIg9upPZFDH
aFSe6ep2V6uGVf0SfWH1Wo59Sfmh2qj2NC1jz700UDQJTuIqR7KEbVPXyBbstIUo
MSiydu/+UjJBQhvGY9zBdFwBPFPBFNoPQJcUbGXpnhoj1nB7Zz/ABmGJ9drIexZt
RLkHi2v7JwbFdcpNH0A+8rdCpMbmA5Or5U0lsFx7XJmvJ96MAesKC++BsXEuuHzT
auLOeJ++AaOee1Ax2609YwexVF1yIzbx1vXpNimvDqbBsNHPKeQH8/JTE5KR/W4S
G24Kji9NjSg+form/hGWWOdTFuGrUMCufuwQEA9pdXLEwNZjBWms6sHQ5iKRqL72
v7dPswmfJdI8TQidI+ZPmPC4HjCKALLPHUqvegV8VD+J8PsQpdv/RAtob9cwQMng
zFxSdUEzd3h9tAoDX9bWYu2b1jnkk1ast09rPg5mZFqqGwxD92v6Pzi0fTf6jBuJ
fcjw88/Zx4V7Mn75hgkygi0OuoUAuCH+NScWHxeHkJE5Gscx6B4BqsnJOi7VNRCJ
5bRxt44hsw13YD/0CUutihGKFn68bB+TCOnmZRjXWUwMadTvuFv5xi86QjLZpqDM
vORrmozsnsS9TCMsAMas5bVlVGUDy7sL7RdVDXBGriSm4USfs09Fw+FcCw1dqT7d
h0MCM9d1MyEFYJCQLjxzU6w89vAYldNebu8TfbPaiMrlSUFXkJZklcNoJSUVGZdH
QgAmn6htj5gVhF6YfUAzNgeLTwNzbsoPs/EBmD6Kz4G+XGSustQgFkHIDX8PQplx
6FZmmHV9TAL6YwtIqy+o7exWwQjnnFyfJZZXcI9exLt3VyYoFVQXX/YGJMa6UuAW
NwMa+uGHQWclqE3Zb+SVHkia2C+A/6W4Md8Fl6379UkkjXN7qHRSHj0kj51+Du4U
beZdEvp5cTj1EwPAc4o5fn2heT91c0hCE9A5IpIM681LT+xCyC0q9XHmqyidS0Hg
mhRKv+6FHnrfQuZxQnhcSWHPjDCqwcXAJepHFGfXmtgAL3GCe5H5PylG4v3Diba0
3SdCrvi/wALsc7cVWXd5ZTI+jGh46qp9eDbb44z5QdI2z30tPKv5FHsxMlAiXFIj
O/zsqzspf+NCxyzbmKQ5DIDZAxqWVs1U6Y1zVCCMUOoJvjaiVFXYtz1wqbH6Wx39
R8XFF5enJmX9IHUKoNT3aHVhICbs+hxNXWIMhanLFFS8Wpx3Dzg3bo+4EtsKRGln
wq15WuOnJ74VqQ97HdwnvrhCjI1NenQMpwzD+N6q0ltvhKOxqXowX2l8+XqJX7eC
pWgUXJ8eOkW4ch1fN1+N+OpdBFcCcHjDvCf70pXZVFFPmQRi/r5gOhf3Zo9HDfI+
qogkOUUpcYbzVVXAHPJDDDWdz7+h8you4VFC3ctfoV1nuJVu2Kzyw/TSA1CQ0HcO
9Y7EICkV54EZtVA8NkmO1ukxdwlk8NhJqqLzK5Hto8S3Va0+HdF4w+ezzLtM6VoG
pt5Rd8zMY2vVb12VeseqGPGpNTnbJvM5T8ueAk7ZzyfxrtfAbJYZSXlAyVVBpBcF
viaHtnBihVztC9zQY64SQE6q/WZ81Hb0jSzh7aZ7RJsIogaHsMVd0YsVcWAByiNp
oO+JJd2TnkVk6cU3e9V4aVX9K/+SKJnrDdLM8QzMOybzdSRhRiSWzf8/LCDJ1O5/
g1qWuIlB4GXexjyhhZw9KzwXJOjUBNk30/z4YPSWIgySn5KdSsYWCiQoC/Xi53uw
BkCYi+bdWYy8sWnna52f+u94ZMhLcFA9x42JhaBXHmSqgOG8a82+8TfybBXrhko+
tbXN5OX24JUGDZUYUnIQKvXKy2hTr/ZjBFWw83PCgLWEcXGyY/PuY97VMNQFcQT1
7s6PSEwgDm8pj5eaMAJ7VPbt7efDTuutjY+qZ4UKRgrxoRkVM0T9CMVFkEFBAYGm
SASe/qgni/LS1p9Eq+gdPEVcP6gaHwtFJoRm5vDoJUN/JO3DNdZWB7EY4zNUhYRi
NSmf5mp8T9pk4GSHZ0OvaQZebqLlToPetcBYIIi1FCWqte61AFT4jxt+TStH/bpF
XvCqgtWh+2X9XKeCY0+PvGR23YLmuCfRP473967w7QybN+0UeTa+x+Ub5i+sH3dr
lFvyLSx69Subf1pUgh2zRIl7ndASHJsMkselCFWDeLiu+f14NDTYPSt3lIfRV8VQ
rjzoNya7OdNvA3fWm/ftwrY8MPhYBJzWzdK5y2VWmG8R+8LlxzE6apiWGD61kgJa
85HAZbq7yPcEZBXGIBtmSLoBFB0VTXkKzX/U5F8oS9CeV06PMKcrvMU+2pWAVFAw
5TQY5kGSqHw5OWIbMeGH9K0fhoGPlgcs2I3IhK/Rzzzfxm6SQk+7P06PlJokStlx
QXK0rmDOPBfkp+7WZ5ty8yzqyUn+8OiSpyCyJ8pvgf2cDlRWv1ft/Yjx3yCAusF1
HZN7MMzuKEw+WkcPmgeX3YmXw2oiL7mfeqZ3qyj+LTrzS9UzFKv1LIQLRwpsp3zr
yP/4X6Z6DDHLSa+CWXwRPGfxzK53sX328wis7pAm0mSWzUpBbyyv5e5++82l3gi3
DBY6StISuG+8LYXB1woaaA84K0ngVxzaYRg8mMg3PYpHtQKdg9hF7kLjAf+ZjiTi
uzNUpbbOCqmTKK75z2Elk7ZoweHpdCLPtomT0DDhmPYN4AbkC9NuZ+eKq9+u0AkE
LooNUtIKQ5Tu2JwZqxrvhyVyEGbZ/a6DXmkvv3laACo1WZambtwV1xP6rLCMu+Y1
HerhWOznzAW24zj+hLBB/hvkYOZPnhdQlEsk9iKbX0ujcgrCWkzpGKFeCrukgiYf
QE0zpFO2KZc4+5ai9Df9kpb/yAdEH7m3rFPUeeF1otEMEgypZ10dph1j+UjBBzZk
HdoBkVbfXCfBp29J/o0p1L/osXGoAVYr2+WsdT04OBZ8iP7+mJWWeughz1jimV29
AqzlrXjptKkKQbfsgR/2fr3NszTzg7+w4EVHD9xrgZkEy/aB/AUlDnMX5VkqOnXl
DROWG03MVFIuvCZZO72mrNgxB824mla/GBLc92EzZtmTD0E6MKgsBMbtg5BgMlbL
xkYWomx9CYxzzPIwSNIcdlqbLX9dprvyOBgw+6GZFXnWkdRcnHBgslcNm/YuCu/6
+KV/SItspWsX6Djg7p1IMwELw6HPXChgbd2VnVdjm/oVe4IFSJ6ve73vwBRQfgy3
V4cL7+ic0dOL3G5j4SJY+wDj9iEEJdHDInyC/jT5ZCzmU5S9MIfACuals9EuOrkb
YXCZU99+2/4JPFW05OR/5dgMHWd8/w3O7pcO4HwY032P3oZpaS2TTNowxLCddTdL
M7arsBoFJ/LlntHIFVsT6s2DFL0MIXX4G69LiX27ZH3+nwvEOJqJatW/Q5WtD09z
/br1my9sVfNeqC48+x+RWbUmvJkYU4jfXRCJsFhEGL5iNEUhWABKvYF0ls2Lq7dj
4za9DSDVECnAC7B2nMkAXA4ZvYb14ECCUVZnUpdYCMMpEbMAlJ3PJDnceZnVBpRH
zGE3+bKCtwrVB49BwX5jplZ7awDjNFrf9fELpcoWjZKZCLzMdmmg9Y2a39B4tjdq
FX76lvMDAA+BkeLV0MRfmV3SCvlWLQqma+qLqAlpSh9JIlEK+nmQ5UXilsbs+FJZ
MbkNzPhDkl6IBRf5Yq1Gl5ir+rC0sL5ASDIkXcmcJqmAHjc7GeIj1601UpId/C8o
Dsg1xFKV/TClXHfLCMjk51/tCDg8eGjjfVMJcQQ9mnoeVwaLlVgDexapP8QsC2Ns
TPlCT/QLolJtE27DHjHzvv18e02Qc0guVXlIean4Dta89blkpVdxTsw2gTjCPgBk
5gy7n7MZD4UiKoE9ahx30aUPn8jgKlnvCOxxb0fr7tzN03RYg4a5igq9O/LaUlWx
WXRlKk3cEZpmw0eyPbGhuF6t3s/HMVf+c9XOnkMJvOeIiVwFBGerZZDeYZBhp62F
D6cVolR3U5n6cWdY2PC9e6FPY+wQXGxLiykhSqUE3HMNRT+/0bzU/zjVr/dfc2aG
znpXTZcuMA2ebZwwp0XiD8/w9uWCJ4HX9twwjyUyYxGjIsCGVTDWK6ht2uZWTEMl
w6hGEfrmu3MBrSbvhcZx/UXYT7qTpLNW10K7F2ZBXz4fOjrFTlF8Ll8PcFXVqDtu
XunF5mu88Lwr//Txt0BO1jeZu9gUgxBvjn4VJrFeR2RoUkHmE28BatvPExJuVKn3
3ygL0+60HWn8HbgElfsRTze0h7B3PziKmVr6K+dJEoGsjS3sM0Be9qwHk/zU8DFx
flmXNs/dXfC17N5WgmptlX69xmaAUcgbXWZfj7OLuH12sUtYOznBrkknJmto4rkI
HuPdth4F8KHPGl1gVqtHnyR47RKyqq/xvO/6WTVzMG0LuSdSHNPfqWdIKmqJ/0hF
yNuoEd+C4da0Qqs7NJKkOqvsDwIgUtvwj+AYrYa4Tegod6SLjUcHtWxiBwzpZFpd
Co6UsmjMXiXtRxzLwJCTxd+j6Jcvtq1M5aSXm+qQtnVJEEwaNQY1bkgPdewvSD3m
//Z3sd9eiuhltyJ9uWBWpJ0OW+tu8yPi5k46V60XEpbOBBSItb0gImoY+0VK5PW/
bQKgBq8ODvdf5xNgPVsjriMkCF5elk1Q7gWM08yBkSghQLkEcHSrXKFqWKk6+Z0F
uT3x9OUflexuInVbJ7v0GRo00ipTA5FWEmtPc7aKokWiBEO2IoBl/d3RDapInyBL
JOJO+baKZBgsy/vlTcyQ6zgTUvrQU0YBYZk5LniZnkVSzXtCyGiJ2m8Ypt3albJA
2jujqPGadlbn5Wmzo4qqX5xU2ZFYuGFgDkKBv8FQ15Sr6vlDlrecC+hzkKiyA/bk
UT4oPakHr3MZFulFrKCXO7FX44xXDjSp64pFdsma8NcFYBBm/2KYYzC8EXD8mx7I
bVrBdef4XAZvklPJc/EoDOlGJaED0lw+YBTA1UEcWi8lw0WMhKvaEk2eJXjswT98
QueTifi2gIEfbk+Z+CdtBqXE1bVfqgwUCeUfzW+79K5KRwBOmOmwqnWL/rEwz/g1
u+5XMCtGbEMEcBlFemaC/xW4cAve/8FfzWVtZL9e4ztpTPr61O5wzC49DvAFNKgN
z33mN1Ow47E8SWQWZOEMRwSi4flhVQ0/qaeBPSzsroJX8pvc9hFSIq+xf0E7j0RV
qaFl0Pj2mjmYjePb0SEFhET37ubP6syLnhRghs8l9FMZxts5azTRyuVv77lljd0/
Sf2l4hbzdrgRddmntwP8maHI5R83DUSLc72m4l/z/RjdkcxoGHgNfPgfnD35HRq4
PLxhaPgb4mQApraSezeAIHxnuH6DiiTAqZ0LC1hxDqljkl96WnswfNZoBXZiVVaK
rzuC6BKc9Et5IpT0RmDDEe19ZZzicWWwMkmZ7+XX4DwByhSUkmvI0hA91Q7Xf8hH
ziVU3CLldMRpJgvg9Xc4Fy26qydySQkd+TXJoYEfNWHr48NcYRCGa7s8a6jPpjV9
WJ2I9SAQImDVPlISliGtwH0lqgSPlQC5YOHz9QAbPe7l/2k1T9ede1XujIP4ivfg
lQLk6x5QvZYcN711iIZq9yUmXtoHXUAw5CbQfPZUnDJOeTe8v0vo+kGnI/v+Jeiy
9B9bcyzWlrFyTkMtJG+/iJ1Nb8AAiRkha23LITXxNAuQrp5z2du/EZrUYjQVgV3s
6n+XVGoDYsHcpOxuHOrlpn+NBuG1UZE4axN2qAVyjgbbV7apKqOh/tH64lQ8K9MZ
4xC5kh0slbVBssief5gNl8cCZKxhJ9q0y3tnxRCwbdqm56kGzpTNvaLTy5f0xQbh
ljBqb+a43x+QmWW1brOHOiMF2bnUaHRQHtaEmRYlZSMEamuo0TaGTpKAp9UlgPCt
zGzDggzoDk2rdnsBQ1i3KUoqCqikiUnKb0uX74LNt4W5fsrj4X6Hn8D2nlnUm4Qo
iuny2o6dRo+vSmuVVZ0e4z6tFFLUwW6Rrt7IVg/4urGVzbMji1F3dXoh4LtMQqZZ
Sfi8zszXPubglXO+0evbP5C8YL+iG25LuRFs6Yz86nqRmfApu4UqIP1vb7gspTuX
522G/OAfA4v/qww8yTrwavNhapY4oHvVL6HmeXPTxkYKG8/hSff0u2Kgx8l/lrvT
HwsMqK4G6V7DpU/n3smpcqfgFyY/+4Uuagvfb3CQNFR9EEB15iuQxzHff2gxV+AQ
E+3AGgnRrESKD3BAQr1KVC/Hts+MDv7qOv1M5p54hD3vXp3BteEBd5zj4m+gAVDi
EgXzjTSd04N1eG3d278v8ZzPAhFRN3IZT3vcGNAAdvGyNF1LN6ZczhKT2cKNc1WN
sADgw5ITYqWsVkcMdTdO9urXsAuMidQUqeT3JHsSkDeMorR6Owa7Zybm8+4FFE5X
vfZTEUvsaVOcbhSiEh8MRhSwk4d7SQV5JWonVjhorBrB9QgopB6rkOg3+0wEUnJN
JNvgkpUP7obiaA/Yp+FfAHmPGDeWZs3uICwm1Bu5XeVcU9EHp4D4i3zNX5+TWH0v
9hJ6Q7qWB61dT385RzcmEOCBXKXO6GSxqf8rjR8lt10NcjfxNS9+CLx+EyuTwNKx
VgPGFrTzqLJKt6KKn+ytHHtgvmiHdPPZNk/kxQm4g3LYfqdu/bferzPoRi7/Z5k5
kWekR2241qXfCk12V1/SFB4ETnoEUGBBUwyYHBDddn1VO2KmDZoUcUGLr3xhsJGW
YDeFrz7kH/BhHzrMb55rONKh+YSuxM4mEpYBD7MYAf3P9Iqf5+nAD+QMnFYq9o2i
DVEy/SFnYLCXcSOMUPY5tdNGYjI/49L1X2SYa6YRnaNYyUrQHdO7FWpL33EMfSdp
Ls049hBy+icZLQ54rIXomBG+ohnTvtTs/80Uo8wmHd3Y/TBVn13qaOgk7QJBVMxl
OSB+wUhjm4CSRD6TgDe0oAWApa0mUtJ5mzUU+XlvcSw/zX7rp2tfCUfe2/x2Kg8d
fTAP/592EBG65KCD18cZUNkevynr9D7cWnBnFblhaJ8GYPMRxKXqiyikfDH3tnyD
wDOB/U+DL6oDk2DlDHsGQXNKjf5GEzAgoL8osxMvmg3WGtWlrkTfv+VhLCc2+KXn
8LL9HQdN6r7ucPcxEPTd3OPWnl8D3M1Vmki5H9gJ/g+mjeKF7+aPhkZEQi5CAKkC
HGQeXlUf/a9JWWK2aGlWhTEzoxR64HInITQkXa/J01qq2hnadiEQBOm2d87uKvW/
dSyuFq3E7/7sksBu4l9fr+RT95yLolX2QUQ3X1cUVmEkXaKnJylN9d/J8TWfp2PZ
lhad6hUwZneP51+DkxZuUk9T7/09Bu7b2bmuzP+7c2vF8/FFdNguq5X4Rt4KGk29
nkuDeiunR6JnxjjfL/GEWdE/wesmQh63FeVjmYWS19FkIuEAEix0WXFBOs5pV1S0
BTk+siKOE48E4gaSpN2mHNrncSuwwgEQC70Mua5kBnjHx/XySbnjG+97MkTcVfVI
Hgf3lc59/aHo8d4HJBIF6igdPWQtgzmJcJNaikHUzwvjnJ0u478PNn/Gah4XIxz/
1vXhs/1qjLnunHQKvP6ewFylUE6hSE49rabGhAk3pcD+WqyLk7VY0bvxZsuWIEPD
A+GvntZ5k4AhjKmHP84JD3FdpjIhvCxGxtAGAnXY362sK8OmXgNuSkMh50zDolGf
6zDr7oXRnNCyU4x50P9IlpZ1VqS5hkCTUguuA1vL66Zd+NnJvs/pyi/DLTxv6nmi
yEV7pbPoql5GKumZbmsCYHXI0fRX+E7ej3czaUBrVtW4I2riJrqebKJji+jE6sG4
4yEOJPEqz1NPrwntKR94UAQTB1kB+EVJ50aEJ9qI2jweAuhfw5T6VSluPBxJ+YLG
Sd4vPug3mDp6gI0LX70oEgXaz0MEg9xbzZ/7tMkSrmaAit2/iG7SbsCasyeGxOk5
aMlzBMVe76bQUyQNPzUpBS50uD5a+4+gSG9M74YeC49xCFxL7iFHpbhAR1UfMNv+
P00VqHZNkColi7xdTj54fldoRIXQHaTxqN4WiyI9My75PSlhrkj4Ezzmj7MV+afL
4ce332RVUxRMn2Bb+Q63LQt6LRwpPiwJZSN9cGhIOM8/sl3NkO0OEoC4eLBavwLd
ntLcRkRDEP+yXThMLsUB4I9hm4rw309FnaUuhqlTaNR8KAc7CAiv+rENvA7YX96o
4dsNpnYNPKOcS5p40IynYXTvKpQPUoCp2bz2gEKcZMXaTU9vvmGitmJ/+DGaN1Ds
lrsziBkurUSQeuCxGBMET4XQKB0MZGTBTmEhjbbm4L8Nij330p2oOr9LNY0mJwu9
4gBU/q9XpZAR7gPOn4LUShNVEVFJg/Q2iT0s7tbaEMNnISv7mNAVI34y8iakMrTy
7i2fTZ8Abjqz0eFYynMYUUwe2GuSQU6evekOGyKtmDwoTECRK700gXu6oCy0g+H8
O7UnRBR3OzukHJMX12PfWDIP88XhYrAbqxMYouKC+LzPEZAaK/eM+SxkxUTRqdV8
E4bteuQ/v+DH3AXu87vApSmoaChkVeaXW//+83DzUUyDLi9UCeJKvdUpNBXsM2Xz
Llp3WTIL78xR2ihlvQNb64at/nRJf9nF3vAvZuq3exjvZqH1uoFoecy4Yp0M7xHX
advmRCYvWJ2e8/xMiAhiLpBMnK1lWjg8hJjDVkYHJN20FJmSo7goXzzwtqpWcNA+
EWIkqt0GZNeALXOvUkBNIVo5vfUX0zkW4l7oyJrVPmiIfv9jNQZ5h1oEPaL+2/Me
qyqJGckbvSVlNu3FU4vRspSBr30zNwSntMBz45O9vVwvRuHkmfwe0bASOZHlcZm9
xu2uAIYF7lZsAvBYIBU1dgs79gjHWR10chFNqBEfBaZfzTP3oRo9zrvec/aodQsO
Tg65EelWSsHlpU7egLCilDmhgRkyN4A2q1q5sG8uslV2AdNer8JYsFFRmJvVainm
7/6EEVibDxamapqo5dYG9y6QAv/OELLQHkee/YbKTkqEaQIMCyQ5E/1Bc+oocM+f
FwfNc3ksenm+PkqFbZbHIir7bZwgpidTMemRV06vnEx0QZ5KBhmkN77l0yjpJ37/
7zd2HGIZ/L0bOe4stffKWhltpLvIw9ut85gBjGrRm+Wl8qTs7ltj9i2pATdqGzZl
DteH82mYJDx0jPGbGJdJckZ5C5WnQqdLbwNQjyWCOqqnJZb8UKPFw6jcXFSJuBQa
E5RGNcYdhrEHhRfMT2vYKFGrpIpMhezwpgjr3VN2kPbHWBQYQHD8D9A20wNkcyyZ
jPjQQOHNgNe1XLvNnslOTNIDbmhOuHS//z42Ap7jwxHUziefL4BzNKaFLOgekt2o
EY6P0lZtM5f2Wx6TZXIAWxHqfB20Dq8NsbJGmgW3TqoWMK1AAwN5R0e9ROsyUzmG
xETiQZh9HnoaSEp2zQm8fUrzjwrbZin3GJ84UcBm2CuxoKqq/1ibpnc3w7ENHch4
cVFJ2klmFi8XOmxxa24jbpkxCxav25DyF8eC7+UibkiAPzbP9CB67yyM5rvYH9UG
9nN14J0lPhxtel18yMluIQiIJlMN6njzxSlDnZ9qDkGozfjZrAMfCbY5F1aZ/Li3
xag4nu1MPUsPMr917OK2kLyREt7oyOK+R/+Sekd/19yqcba+dN70A0x7WBbmH2Lu
f24DlH78UsNQnkk7EotQuaUCBOKoRAyIWHCOCsl1+tj1DSGjmL+up1DMXLX/iotI
Ev8C0nxEqOvq8j6LRmtMx6f+qZ+8q/24fX/zh5ESSlhz2dgZmvVQWoFOm9ycBO2k
9fqftfFtEo11rb7UQl5vF8jC3wx2Sd9NGVLTAQxfnVc9QDX/I9ZNkRlr21OGvY2v
AzfF29fXCCgqVGClIH6BifHvESOfnVWwRV6LBq697VWO5fXGjVbZYtZtpdsShDIa
39ECDo4g4Wxtt2XGb8rMNzxLsY4gqpM45KpoIlMsO8vIrE0a44U/FzZWTUj+/vsJ
6bPaCc76/j+qPHHXenXgDedie2kamBqmysUn1OzycBiIUH5wOUbWjq8ENbV9Ju9E
pZC5VMmvOqqJ4337eLygR7AXDrs10IKob901g+vyYxPGtPONTpBqFUHi7bZzw/pf
GeNF+Z0xb1olZLaY4PksqBPEBFeVU7QaKuuZ4m3EXKPzatIwbW3PQFd3IQ9ooUTW
s79uCsjR/AanMhTtty4U8+GipX/EH5phdE4DKzUCoqqfZz8o3hgZsMs/zkslYOqc
VEuP/NWtDY6ABoXonJE8fM7k9WWIKgrlaUJnSoo4Xjfo+bldgAUO2iN+bqDs8Slf
oZnIHj3tb+9R/EM6y45xLT32MsUwQieYCXl8LhsKKPX8VIXLQ/TVmkHpCZkmF/ov
d6T5fbOMY7mbzUrGaReyR4Mv5dnEUmaHCZiGuLSnGAiv+ML4C8uUXwhLjTXz8IYD
eTFg1pcwleeY8uNu7Wb48v6H1KlA/QDDf5Y2NGa7fM1PuzU8qgOE3mKNOQT+QTyF
gzqpbX11jk9eqmwR6tFX8Dk4RZKmeoStfCS/t6yGQsGr2d0jQ3GUugwe7i1gWZ3W
GxbEgGwc2nmfC8Iw1T+8MFedj/5hi+VcA2vAbr/+yiRrvnMJIPV7Sjsg2h07mjYn
ZsEZo5JLUTD3/rE8m8/FftI1TzBfFnTdKoDbcEwGMhQB4wQGqfrpCm+mgMQQ+k+8
2mC5/3/eRDFshkAd6VJ7T1eF0KdlfIYWbdUATLVt/DQMQznfMe4xDEq08a2ooyPv
aOZWLIJ5WTJdM8Xas9jR5IgKbYRIBZSOvycbdTz1uRzrnYiguOsLJ2o1aDsDZPYF
ERN4tnvngdxQO1h3CD9hgap/0tL3x5V/SgJ3f1GKNcgTq6Mi6sqDfL0jCZRXOkb3
NgGKuEj8G+YrGLJ+td/Zu19Wx9Dq3cHBiQ+CfiYEJmnA5PtpCHqQZUghqBpU0mNN
Y+zYZ2qlvfPGNDQ0KhnqqAGG84pfQyLjgzYdSPwdCvshTEugzpPqC1yUEN34TM51
EcBZUdQW0Og/nob0Tl2EOFvJJz5yj/PKwJ/LIqOoGH1H7FuMuIgLRS8+vLBi1paw
MN3iTPLCOqEDftvsXLBA2nbkb/a/HYN3uJwsdBSPhCUWG1iMDO/E0XtsEPUbTqJq
KG/eY3iD4fHiNgc52gkruEua+z1SKkurHeY45wzPh6Uj018utAE+ps9zHWo8Im8t
OE9RqAp8hA4MzFhFib4C6xOX7yQkPkC8TpPjO+8rfEaTt4tcRPTV955q2pjgmqzk
j08jvbIQTvl5Ag/DCCyzh089tZJnUr22wQIS2Hut4sG/E/tAGHy+E6Z4epXBBoHq
b3NSlIn49yHERMXdYpB/lT6En8/lrHRwx1jAwiHaDiP6t7IDYReu2DS+rHw7Ct/p
Ymv8Ie2zrE65hxegJ7oSJlwfaDQetICVFTgeiJyLcqMRqJQu3ELLwZT8A22Fib/D
y1c56QPKHkpEqQqkO1hrCtgeNXaKkAGLVSyXKS6MjLN/vDq32FFclyb2zJxPCu4V
SFax1lHHr2SG3lZdQ08X3suWSuy2/N0uzRUe8RM4nbcjwBCiS47MUGn6mfCgrN9l
wQ1gkDRwHY/X6SxlMB4bbZ030J24NKj661QYUmYl5kFRO92d3zJwm9ABGLu9YUW9
XNTFmvN853ZC70tsoJCMwuvfLBpR0l+ZyeWeDjISsM7tVFwv6U2zdq3mnguLCcdP
imTATsfWRZXFTHtBnGvoOWV9OsFpCVZbTJ+NDwZcfUcdnstbd3VfJV/buM5gA5tw
n2KDVuX5JDTcgznUI1I2PVq0rjNQUcIqr3bZVOmHtcea0ipORiKZfHPCMSfiQnG/
ijQKFUzZ0GREc6+gXR7tSum2130OwmdlhcXPfjerodoziil1ibrnxxkmMqz6BlGl
s3uCgpovacTpyZk215KHaI9WE7AUhxOvy7IA58olYRxyqs2TkQt6lCTzJr9v8yYH
H2f2LAfIZgvY/tTJJNuL7lQ5BU5xZgcoClrm/jb/1OZfL+sxusWIlulmuKsWRsyp
1Gd+ZOvuyi1miTRY6oaVLZ3C7OXW3OwkXo3DTYZM04+R5kfd51AnxHr+cHCNi+Yf
Zr5ZmrCCgxITJt5pZ5DVHJ8fVdI0t6Zzw02LoVatDCi10dggtsXAArVtVyLd/XgD
vnOjWAHHPb/8R5AWtdqmOabBq924l7xcJVhyFkiMU0CG6KHtfxSkbX57FXwv6jRj
LW9XP9P048aaZN3z6oHfpWu45DzyrcdQBo/V/N6MfTwB1bQP35QoHyj0hvVq8K5b
/88R8cgWtyKCLmCLwIuTSvlsHueq6+Bu7j6i0uMGa0WVPWaUgDJSBLw2mVz4xUXw
w/rmaB2sPD39P1U9NYhfYeEamNdf50SqKyQtYs555amZOeuTAoT9rsZLdAdQ6/LO
VCL9kQxcE7teQfHUimyYLfTT1P4EcoK5pvaOxIj29/CHi7jwYBH+5VEdGAZcDXg2
F51MvMwPVR67zvzw2E8znAmzPN5k36T+ta98E9IRjHIflASMnpu06k/57XOqhief
XEe93UVNYhLq9u5xgX3BcoorHuH4d+MORhClvD431HL9GW49C1R3I4LIue3727vR
twrgHmgSojgPIJ9P16IubJYbzZRK+sHFi8oDY+L4ByDD0eSa3QSUXfCj9SA5qoTl
k693aTCpfLFe0MxiH5kjHkZbo+ZACP9jGhNTRX7K7d967TFd4o/3QukKE1p7kk7Y
dzn/TtNstSDyIupXVfdYk/nWY2Zm9mxDmzq0tYK6iGYlE+rLjvcQro0p41OAZOE4
eORONxWIC5Xjt4eZ1f3Syu0ArDdSwQBqDqC5YXiQ3HzHz1OQzqDoZLut0x2KjO80
fQ0gMp3wNuwNNWEnlvcPaKug5G0SKeo8HskX06XBUn0CPUInhc/quN0iUO8ogunf
wCDnkj37sHqpGY7SQYZ0gZnBaFQhRa08AYwujmyqeZLySH6aQfLCTm+3iqAcg3yC
R4tqEHbFrzskCwe5EPvHC0WXDqmO5a0jnk/P4w51IkklVwXatZDs/95nY/y/R38G
cORe1Rl4pxSBH79ApYaz+TVi1HqP0jvxHyTvWJmySpicwavA4/kAtXBqZq+Abb+3
CzDLJgp8cSlB8PkjxW+jLZFAe3SYDa8MMZRM6Mf2oMliT0z9IxJ4zLo1K63OYW+h
wccX5pTkctKYxI7uR32as/eJLo5vvnMc38bsxYPfNnJGSrdh4AThugwcf8WQiZMA
vlAbFK8OXG6RG8UVS3vWNBmQ/NOTH/WOJDLEnDU/VqfsxFXrdrHfBknewKfNAXJs
vvf64c/EMtmMSkpB9py8q43uaiJUk6B+T7FjexDXtzusIGc4TvUIvJ6lSe5HiZ7Y
JjCqAXsR4dOrlEyOPpDJggxPudxHM4M6LxMC3zUmnnVO0KFnx5OKaukAEGCWmGzg
YUImiyHrSf43wWTXSfkIdLttexSRWuTNQAagVHjiOFBIi0AqO8I4nnykNQC3qjuz
Z5kG+62aAWmnRjGgKup1ZCjsSuTtEOvoYVvHrh5v8DEXXnfYdmeDzSr42t+bbG1k
IT3J9ddmMMNvgXuZFhapG7lw6kxzpPpJbBMJsA/3JjwsyYOemqpyBNzsXg7MqtEq
b5NQqEZ4/r6ReE8R7wE5RkwBOaf5h94g3+DgnBVWfRCwKG2FU5NSlRDLf7ic6TBY
Od8fG1Xc/rHYC2LzADQhHg4+s22S2XfuQUcrdv7HOR/L3ABcK0SR8+UbQmyjIAC0
Ya5NRjD2ZmvjWn9oTR29llIHl3l9KKM/I0NfQt2LKHWJEUs9kQoJmVYtP9ThmLVk
rVRS8X35r7xqtbCLuhZJp/GR1MUpcQocPrVVECtGhfCT40eA+sGG2KBjhsFCSYyS
azuvvG77wYhk7yU3C+qUCgwX7r2AqUgvwNvVO0ZUMOVAwBuZwxwe5UNK5GcUP3Ej
ZiAnwwJ5WTxNOPwZarqRL7n30oUFMEvlbd2FXQxZnuVExIzKxpjt3lghqvxeLzBV
HyuDCIvYyBtnV+33XxJ8uqNk0xcgoN55CmmsrEFgsCCR9+J4NJBQpO41pNe5iZum
6vtnfAlEoCHgLKbWEMDGUxMDe4Mj6FqcoOOiumXCDBJLKY3xBFOXiX9qYnWmuFq+
aeaxaeDO9dRF0rimuj1DXtprNqYbNbjgooivw250Wv1cQyxXATh0eR/snM7FOJbD
C2BsGSnn/n8+YOezbCPWKawH+JfizpkHLgS0Om+MOFsB+LDoLdOVkwwiThhU+axs
oYZGvE/IUHcJ/JirJovqJPl8ra09sFPI/xRK2uOLrgZYT6fehOORAnl1Zlp4U/4k
B510kdPeWZDBbBaYg3+7UTdofGDsT6radz3uxPyQA5SQ19lX1QfFxoCwrgrqNzwJ
BvohNC97Ex0Q+kWTp8writjfS3KQ6iQTxDGOvZtmgQ3YdfKobheirs5AnBTtSY8T
Y1ij6/IZxDJrJfesgfN4b2zM5cmJkBkLa+j/FKzQO+kKIEncobW8MhihtEYBpngf
LoxjBRHuGkH/RRqVJ3juKEWXnDRmLIuDD9wRp/jUFyz0Qaey+q2CyfDM5CHM7tlU
h5iKzyyAoMhBjk3a9xP2EdmjiNyF8ryRw4m6kBl4eITVzko/qk+u9N/Pz5ryVnX5
53byn9KZvgeX2LoUpQAf4WLkb4KnmM3sBavQcUL6ZH8wOySSm1gc3c0diAKUMZwS
L2XE0IFGQI2TcJKLL6OUidh7yL0MG8/x85MKGfXGUMHM2iQc8HrdEgteArHWQRGq
3n8mNxP33LRr+TKJt2KiVr76ES4b9eHuqVEp+1KVCrc2QhGqupO8c4iLZwsqSyf4
G1Z+0BTXvsaqMguq8KY+cvbDRLIHAB8Qok2f2K+8nWpkczLkPGOpIM3yy47QTFJF
SPo4JvXfjv4PEnbJ4U82qx9XF3GcLxuc7EHJbtJ/6OhZ7x2YybhTasUBXTaPzfS2
pFu+unx+XfVFcCOTpzyi2+5/cSXBcUjKAI4rUVzDWGslKTzlAfeCmno2/ERrEPCY
jWzhTtyApOqAe46zOmUfpByUidQBfD1FoXx8QOlFkMWKQ37QfEfQwEsgI5hxfeQw
/vSmt5MWxWRMBLcldovAv90d8g+wGmmo4ut34vt1pSciJy6AeYHw9XU6Sn6enGZ1
lWCAQ9MoaeDAuwIfv178WWCtxF8QBAYoJ2C09cbrBWTrJ34YFCbWD7NzF1jk2hb0
+ar9j0u4SiMhc48hWieyp9UAw69x+m+rgojCwc/PGEZ+yMF3GJgBlNA3Q/W5GN/t
bAGZ7RVHfu8fO1CrbD4bCvI47nZjDjzqfkgXiw9RZr/G7AYP5WTxFDv+Mq0vZNDC
jRUaPkH8uFjxcLA17q9B7OtwJycbADkVQMy/kbpsqHBqB7VEf3hdYaXZEH/ULNV0
9YbvCL6U6p5sfw37zJ3D5sCROQY8ZHN6WqwcX9hqwRFAHBp8w7FJFMUfXDVx89+B
2wnlLU4sQ/LiO47Uy/oCJiHgfz5tVEa4Ip63u6MLbA99mIDfmAiwO+WyIkyxCmFn
IpTZuiLCwlbHkU1cHSMB8YoT3VMvVZGCP/J1VybHG14uKSNWTMFROvuHfRqjX9TA
zpY+8w5PI5Ep1ECIvNQOX3/gsVMMdMTJmCfGHbP1iTrNjqOSrUgPrduwsczeTZ2Y
ShxZQmMTV//LZio3Jb+BJpGE/uIEOCorV45qHDlnyfZOKsYV9flVOdv8d+/Czhep
AjuTFfhj4uhlIUpDk8qDV6d/63Mu8a0s244D61STL7utmAgLq8UDLQvZPrsje28Z
LAksx6gsUZgabGfNTeABh5oqRkrKlyeUzlvxKQkGksbQqzruH01rAnPJjvoHj3kV
3+BhFQIPWZhfQjg/yXS4zGLP5EJUkMgbhHbE3vs/raozYBW9St/2FGXTT2NmWwQ5
V8cZwDDJ5sq1Bf7vlXPZSfZ0qhqqz9S1QeTlTbU7iLMOqZaFPz77zCpBvw+EUg++
T3Kp1RoVeStaNbUCmi2qQasG4ZpgLKGe9cqo483FOHHzdbL3HWd3zticlWL1ovEb
ttmV1aJPQD+elQcr3/BBDNO9XB29ivt/13qmzy6AhjRmpTC5pbaYszHBJOuMuUzI
298yUUyUYW9j7VnhWL1gYUtwboES9qDlOgYAvjx7IWeiHcwqk67alfmCP/WMxBux
gmxkR6EM+K8jTkl57QsWf4lbmmW0iYfD04+ubSt4+QVQEagkwg0qQ2v6AcUzAbdD
Fe/IXfOePUZPf+vwuiaU+78mBbDiBFgWkaS/WqbvAv2/BoIlfMqwLbhyyJQ0LBAn
npxvDQ92pbpK4nouR+AsraYMpyhsvQrZmIUpJzPvKTA6cb9VggVndZSvYNNh0Ibc
9H9Fz4IqjaC9bXPR3n0n4FwcMhfdjBKERJzY/6MIymUoxYaHDhwuiaGDWaVVtzxK
SBq+yOgNRGVs0UqkGlUqPfnns8nJHmQw8AwboFd79AjpbdETUI4+PQK6kD8lscUk
xmtxDWXUO+fnoL4KtR/hNwryy3bLVAVzjZRrClOuZl/8b22mbCtbPZM6thqWnbbt
oeP8Fs8yMlRtFoE5s12EGzSE/1lKFWfACNvf3Kf7QeraPbKvf8ZA/+avmjVk0LZW
oqVUjrFE9dpU3c+xgIxegH/ChkbOfIj9ZvIexYP+4c0OUUYu3pkavQruUo/Pdkge
pVvdvAJJ8SzqPfeBMJx0PEmDp+NHlbIVhpD0L//v1JbXmgm0a5FLpwHSKrVNVYyQ
jBpX0q/qow7hjSQd+NsWnn0sHU+Jz+YoIOjoG4RkpLgoVW7l0LJdvxiJ7Lj2d5+V
HFjro1/E4onm7U1DDn0Evw7lCkZNccHVPRKjAbNo04L0WFg7Eygn8vQ64vy26dmR
GcjDrwa78HdB9kWWA5evKNUAogHfbU8rl38KSyCuDLUrfpUFgyT+uxAm1Gc3npkh
IgbTCaTld9+5QYuOrETNDpoPg1hrbnIKqGcTbJKL8a325pe0A7cr7NwZBNewCAs4
QpV2s9uZzxZ2wmOmDAvxBCj/tBs7GJaBmOh7AE2+2xwKUh9DNFmf5txMDKOj6mkF
jsXeyjTPjgsj1p9LwDhEJIXxkVuDhxEAyoRJQPsn4okSkbOkEksbSMMKiPeQxsUu
87Z37cJ6o4V/4wb/2Z58AUi4VXHaSCk2qb9nWI4iuRGXkOq0uGopZQORmaQQNnOq
KdBs+L+SsQSEwWimjKCSVAHRWP3sJXBe7KEHOSEQjYeolHW4/mLJcn0kTX6j6qtH
ltAZbo/NtIQhwkpfzO+IkCrlaYd3oqSiDwJqR75hbviOXzywoGQWSDM7/NzteewY
aF0oR9Wg3SaMPEmujgEknJ2M/+kvQrsKm+zrHx97qUP/GMIrlMRgQ98kRGbksHCS
yo67QC4AN10fsO5MQekq9pdSAHsSpD47B4GI1UY+86vEvWykteWqZ1/WmQIsqRyJ
DsBSJ1Z9rANXhe98h887IwwlZ6clm8a+8zYReQKONnb2BieRD3e366voqU2ya/KI
FwkkiJEY/Q4FlUiWNRsc+4X21l8mBabrHiVfyHiZYIkA+W6HeVemDRUD93i5iMKp
WnLexGJ50TiWb+/eahu8NX3KvwFcvDleKnx9546v+uYEzbtspi6OmzVnGyVcPfDo
sfaR3NADMRWWPxkNbaDe8etlOUalcsdct3BOZqbrw6TrLKGzfYIQY9RiKwygnXJU
fyj9YwsC5mbGEyZ9CiKZzL5tqkUGxYORfsX7EWh2xfXTXUqfa6NTiAaz5aUMsbsl
kfihLh9IVeeX1TLtQKZ2jwdvZZm9UgfIOnyrrZOBM3kY90DoN8hOxH4Gpiwl5uRb
1TaLSj0NXvz7iS5FaBBvWtO3FhFHBmORsV33Pz63JAl1PDfJRpwqHkd9A1YrdLkz
VMra2My3+XbTVrQz7aYIqD3M7MT+BAEOmXyGjoo7bqUeZhZM5sMg7B9e35sabrHl
cJ7Jct9IMDEJ/U4riez/DVC6yRsBj+Xp24QqUB+qdjY9cYqoWDyh5tCUxcybs8BF
DfTEYCfZ6A4MUMPTx3KBHOjGH0uN33CAM1N5Z5StBx8ctjQq+11YKRcfqyDP9kzK
DG/0PMQQNrXJAbBpCSIP7Yf4nqpnMYaD9++fCjYMIp9Z/4UfWj7rTeiWma+svG+9
bylx86KWQzcfqfCsllQGUNtUFD5+cmh97sBvNIMrUBJJbL85EzOEuPvY6DNgu7Rp
u828v46rRrCjsSF9KC/Fq+FXpc4kJe9M7PjKS5r/gZqXfKxUnSCf+BA90i0Eaxu/
2YSpXRmdF1uMT9UW7Db8//UyGJ436MZMWBcOdUpJ+nd2M3PzVB7xAhRcpsM476So
avwaxD54km40s0r0XmYJNUwYh6ISrZAuMx56A+ysXP07Mshaoa0Xa5G5HIzUGCJu
Ms+A7E3LUVUuKLIEdg+1o12cHoi9NUnURF9Rz2FpL7E+Id9p054KKW39AP39H0pR
4wcifEiD7JuHIIeeBI+oF315DjgUkDrlkuDQGeAUoVKNBq8BS68ebTMZyNmBI8Au
7KpcAyNc+iF90zhrgdRcjdMJdKvpY9BN0wgkb68asa3ETjD2CW/FgpihQtKKZolc
RgkJhUMFq9mmhf4z4YJO42tnbv6ZQwGrfKV4HvoqInE8HVsMAgYnoWfUKsuqvZP4
2ikzlrzw0ILJ2A7ygreejFVEs4nWhJMGDYYvbWn0LTG1WBF3T16wfsIuLY4guEcd
gAWQNj1DZsQ1kLYVzTpj9LNdZwAuSSNU0vw385MfKHVd/2sjxEMB/RZfrH5qLN77
1rxlV+1Ovlj7thzWYog3MkXvC6NqdXjhEdcIxemSWaJFWlTGhXQoZeI7WBhd0y/+
ETGgrRXy3+A0/XyAoRC8MeSbxpdu/vSqx0Q9bT7zrfBSaVwc93Jr+NvJaR8juUzm
PGCiYkKJL9AKHdhTiWqTJ9IvJ5GVKZVYLEsS4W2ZIk6jGHpQ/iITe54mRd3oPavy
seCMi82Bf7z08+s/zd5RY/+DnRVQqTY//hjVj+RRE4FYU+1KJg6bEQQRgAyYxo4C
d5TPXSfGNvmhSnMJzQHx24arszsgjsvAv+3fWiMwWDLUuehf6xbSbsghMlpEMsQB
ie+hB49WJXnU2/0Br6idCz3Oo5gIk6pt5KJtINy9MDYI1N6DFv7p6iFp0IvaMo8C
Uf3JBdu2MCfHW64qCy8iRpHitd/AGGBagF4Yb5PnRjkf1sKkWNLae6M87h3bXDbq
Tco8Wx8EL6ezt87i4Dd8cEh3eKaXh0loGuJ5psRST0M+e+jtUbddLes2OvN4tltz
5d53xKzfQImTDeh09esBK/7ggJhKBZaYiOLTy2uRoPhHgDeD68Rt9O2yU7RwZoPM
0SIbTWydxIL4vMDmhGgQ5BIDFKm0RVneIWLi7f0JELGJz90/t6Sr6D0MxQmOfziv
fyxEa//axbtXiKv8fSHpaCiQT4yTQfGzOkizFeWUBDHtlXH7wpbQJeDi5ddPgjMn
E5TlN0mvMvDVS7V9FVOl7/zOGikIc42FAd3fC4Piw60EqMZHa/J4YI2wHd4wy+YC
RUz6vN2DigifOMNMC7SJsgTPPrTJiUJGuRucTJbB9udwG1+oW6a9Zdr+yN3TmqUa
jvo3OsJP++oNMf7+lcMLN0Me9j35mId0ePtK7LjITQlYGZ2TLTwvCiQnblXMoepl
uBPDKwDteMh7dVQvjyQxHVpdh9ZgbGNEoZG3D8ktJOzlVZKzyhqDOshJc0e24Ujc
5ooS+QbJ8k1Pg22N18hJEwYO/v30UvcHO2L1AgjaaD1EG01nSZhgishn5grhuoKO
xjlb2FrC9aJPID6AWsLrkbW5LFHCcDDmmheKhfYh6xEQuQK1cbvuNMFE+WDiIesk
MSmwtot2e/nBjPv7CSKdHWBDhEpvX/t7rXVWynpGRC0GyypVBAVwaT1QnP++Tnda
JwLWwBkDoBUyf1b0pGwiCwDu5RPbKElGhX+wjDsWeGlsUlhSngsvfFN4SNOdMf8A
FrESodio7DQ8qVKpTqeTrkPlqnN2yh8v2TwMZEiKXlDacljkFtrt236I+z9p38ct
vw5wPkXJDeBxD/IQyvdjqHFWqAkzUyFavpM1Ct8A4Z3NeS593U2s90p/WmjJJ/Nf
Gl0eOMt3hJVTDiQLHqlX1q2uwSygyprRfdWvtlykPAAdPOal1W/duSdzdWZTD5qf
fB6tTQHTA/d85JPCz2ex+erE+gTqPWnndr65RUS9askXA2fc2sDJ0xxJ7BAdUTP7
bdIj3hriRhNRUmZB7apKP4LiqHZosBx2vta+lslh5E0QazxOd0LwsfugHdpraQPX
wtWVFJYM41lDpQo1Jomu9V5p37AAACzJ3rSlenUZt2pMZRbRmDPgiaKnMPbIBxmw
CTtiBYNa26wiaq7VZspBxHdZMMbppSQfOj5oi4ltBnjfFDy6pPiiDc2+Crq00BHU
2CBCyy9GtC3akJV0LNQMjSm/Ne/H0coIZc2mstAL/XGxys64QuB+fHlYwiweV9b9
RhmMyaXilzM4dFA8/auMVstBefI9+F8A4T3xoBWWeG1nWYki7EkKlty9D8e3JUA0
bEnwypX71br0un1icdML7++S5VawZYydYwL4zhxM+ercu2uhfmYHSmxaawyU21TB
AfOeD4bXd4XjR/z43Fi7s2oH7kOrYsXOCLI58a7M6oplTVT+9teKN/nyYQMzywvW
kt0UK5GZc9gwOaRkhRU4VRkmorj8JPPpfgX9P2kQau9hR3X9cRSmtnV+vgJqmCuJ
nPf9CgGLFp7R+26FzUeM2muU/lMZJEdiZhcWvrLelkeKq8CJGN3B+5ycAP0cce88
SY69hRNNz9MENlcT2Q48tzjUhHEepW2zZvYMmPoVqdMeD+CFWCxUMH4DvU8dMkC7
5fPtgmgv1Mp9IAtIOqcQV/5+q4i4iBSFdvKDd6a1ws2IFOcXG2jUfhWsSyg7oOT/
1SSL00gCXD9R6PzfFqjaBraPEhw2HDyj4qNGXsRO4jVqNP5p7eW9msYdYdDo1URn
ycgrlJ5S2ejPrVMORL/Ejr1pHcNsk0lDYAZWUVk/EFSbzH6nyNxCr+8T0/FQrANB
mDFawjr/Zmqpgw7PG/N7E+RJnexMoeJU4/YjHlRhOHTebIMSxJ7zX7oKBN9XnWTx
hPlft3ZnjULtkpFyuR7kF/r6qUNi0YIX3XWvF6k5HlEmzsS/Y3EJa2XetyYrSKpp
/ahDFLLVTF/QEVBVcowDd90C0x6Rb91HTPr648KThmp/FhipvRymduSGTIXJaGMj
ak+9bghio0lLqcjQmy3kSkvG+1ciGVAFplawPODouxL6gU11ESswXAzYnt1eK98y
XF5oq9QMfx8tAfQxnCgmLvh7SBhuOp9g/vNq0+iSy4oF7RsrPIDnhl5wy7yZdon6
ygWCZWwSLkVX3ZTb02S/MS5oYo4SG6c3CDSi4zLld8ZuAHDTQGQSnaYEWqw96kng
Rf2f0In16v5se5Vy8wkjSRNgHlcaVL2T76Yp22JhpWaqbaB4xrN7b9pugSh2QTaR
uffPpeLMbKBGrf4ljFasayX68BOLn7ZD7Y6Ga5YfAn0/O91/l5y3tM8Jfg3puOYC
WVkMuX61FaZf2kycbrjSdiNaHw1U3fs/kZ3yJJ8PX8lOZICA/90fqLjYV60NNBXi
wpX//Bb9AXo2RQNoS8jSmmMOYsFqL4U9XZLVnzEdX595u7LzclpVtzhtbxlAGWUL
vdFjC6q5vZEubu8X/29RsMFIxYijJCh/klnUy2jecLObZ3/O+3J6sLx90tSXSELq
pjx/2+18o4vh00rcVhU+kNFstZXVpzNzaoBFLCc89qWmA0nMhdupD/wwN7SrKz/3
IGbNStXv+pBjdpphkAGpcUxvMrCyeq22yg4NUf2c3bQxsoGRFWY1zsl+FfEg9Pf7
J83OwcYbcH3t5IkvAR2ioUTADQrjPLIXncJOUaY5G6Hd9/3CiPX6J9Q5+VXFUye4
uN3vS47LeMuB1szqwCTc/3yqR7zTCMC9BEidu/EnZlz6A7VbawelF/Qf2iK48rNN
WAtaAGAQanc1DQy2vqtyvbqmeC5+aNy0jRM154eZgSln5xsY5RJpBpuPNRwjT+0q
QEfuI8cxr+bKmnMjk/TkScX8B+6MxKAJVKCBtVPLR9eowh0Vx00ObZwu/b4a1N/K
8kto0+UvVT3ITY7TZ8i+eS9u1s8EIMH8z8R+kJyt9/JlBx9hBW/vYK4L4lNp0e/l
VAN9yvq3lTxrfBf/RSA3Ct1aKEZ6V5/BmoW7YmyWt+hk/m9VMJZrsPn53Zni8tVW
BQumaSjE8Zuj0a7cSLNAXcBAdv8vEpX/x5HjJXQ5pnYaM4Lu1HNON44rNTx7KiIt
9rJhwqDIsKBBR98k6YjzS0qNmItlq683lKtHVgZ7WHOliC6y7rQoi+oinW5LwEt3
tef3SfDfrImFBDQDMKR0nWbEWeFLfq7w8WdLEM1sXl0+x7GDeGSfdA4zQ/Lima4A
qShCIpd/ta/1YZKPaACM99ISq8p0R3tVBeI1zfN1ygAysivLptbcpFpvTvBqiPCD
GX2Cvko1c653eh3Mh2B00mh6OrLqvLQAf5c5b2fpOIEq2kWu7gxFTR3xHhjdMno0
wFY2Q/EX01DNxXED7Za+FhlvQDripk3bq7YngF/g72aOiDzGJaqaf3qJoGd3K8Ph
BaLXCezjPmaSQCUlWUPSUdTsb+FbNxcGfRLTEvSV8UZV+qZosWOfuHgBMectnCDi
G9efgJ2nvilSr+utQogQZhfGzx4vCE9tcQ2tHmD//QnAEE0880SBT2l5pFz2Qqnd
QPuQlOAAlPxwQ0wUb4Sh+JqE7usehnUQpc+LGbqdGld5LiZldY3B51yI8CweeKLd
lV+yXX+W7oXFk7Id0CeyCI5vyfbs7CehcpIOPI4qxEuGy+Bprn8BMk1tJy77m9ZA
mBrLDOW5YzTqh9v0WISSwlq4+JiodOZCv9AZ2i9gJsROYWMPVRonQ7SB5XcOCNyE
xbzwSe5vJIZu3fpCaXw5QW3KFFBeNN+Nns0c2sjQnkA7Hwricv5UR5ZRmGsKYYaZ
lKgpeRquOET/mp3Y9zulnkmvkKata9XLFZsCGS5Xj4eU5HBCXrdYgwbZvWHc8Sha
M9imUSIUSqDT+iDYDhOr/YtpY0MXtANWX5x6iweB/2Emc5D7EAA7/YLeDvl2I9po
kUhm6y+ZARhsyqOsycap4KO9VaEW3G8dfRiFlUb5xYQcXQF2lXbALlfltW9BC6Db
5nRu8VqaboSl5im3dgc3QDLcfJhDX2mcVKBg7hIDtEYehzHIbXIYHFO6v8z8EchS
+fzICjnf2NDCYRQveW+0hp3FTDTtHcJmn2KlGipPy2Bo885URlI6hYkQvzoyDxiE
ILsoVJ5uQC7XAH4ouzXyNdsCh8Hxwkpbtad14soUUTMRuJNY+Y9pm8tS2GjKnSBf
015TOi91HrY2PFm+qOFG6w3fR2sa6HHPPvgSH/oEiu4nYIcM0RhZhpryceGszQb8
NDh580bwMri7Ws+myzT3jU4wJIoLTHV2aLhq0EwYrDG5V9gOURf/qCMGP5Sz2V8V
jcCeTRY9s014poS4d0Gd8sbsef41Nmyh72gPcDQ1YenLlrbbM5+Q95w+gxeJZ5sH
SHs+VQa9NLgSk9uevlXrsAP2W/GYh5rTx0EAhNkg02QWY1rDyoi+IhoRLKCPsimw
fHHvX0X5duXE0uglfVdwTlEn8n6tSTFtkWwW5wDtYtMiygDfReQDtGZ4RdGjgklq
h2MDxnpmJqsiR0pCemTDCGHh3BwfSyB7lTfY/rBRK7ajdgMwpPZdVYpgQ+pg5oTs
1I968SNfrQ7r2QUi94VOue0UDeFAgwmaXoeZpyTm/xQ5mIsJBJXCoGeohHQEsY3p
HNJvfXocIceLP4WzdNKKPeY5Mx+2NNLKe8mJOP90mAOjfwwCGX+wODphwP6C1tVK
uaaUee7oGBXMBGfmQrrymIH7JKQTHUwQ6ECCQcVU+1oFP0CSZV06eaB5Mmb/dwY9
sUugz1oOqRLArUI7oZEqv2+5S1UMYXBJ7FnXVTj+T6tdC5lzTYF0zKTRLt/dilDv
Pmy7McX95+vBepuSNOKfu7QwDddc8vElCV01pUMHBvgtQTg8dVFuX1Sxq4Z6994i
8aLKICkbzhfRVS76sZ/n/MJQ/+ZifJoJLDSSIBBjyw10i6uMTEqNrqW1zhIs0o7C
peUBC/7MQA6Q7WvjMmxN6LFIAq3oVAyePxg1jsZLCun8qdzwfipORM5Rz+ZDKboA
dMksuFzgSvIBTNxtW2YOxaa6PgOVFT4omaRewjitUvCRoMk7tCTUZlqNlx/fhvx3
mJeiGHYeEt6q4Iyy8XCb7rEwQ9xcKUR9ILXKj5T8vzCvNRGtButvkQ6h0rwWcrWO
SkDuMQ4kl9IdkoFbusxZ8ULNvcQ8PYcEq6WXooU/r9p6pSXwtmvDj7bbY7O+nBgo
r8E4vB3AAJXdMuJF0Xe/X0LEnB5SBMVY88LIMAFU2sRVyVuxGmENJmMNOB7Bo4HH
BzMqBvvYZwsUPFaEqQYNCiNrGNyudgvhkT4mb10GNQps/5AfOSLO38gMaaFvwaxG
iTPCzhcSc9GDfUID6ByeYVzaDoKUfYfl9Ig44ZxFa7ncngYwgklWI20hHiosg+8r
hxPfHx2j/kYTwUCjZDnt1O+AtIpnux6CW5y/JeXxzwT1b6hiIUwAz12wywFj7HVf
4AjR5YiegMkYLPri46UXBWy/B3rIR3yNWcwDcYZijAH5oLPwiJFFI+Fib50R/Glf
CtV7cxTUc/zPvk3Kj5mT0xN9j5BCFnupga1PwO5RE5OxtINIfmWYlJqqDOoUFiZi
zXznJYWrK9Dj0zu7CHTQO8PK2wW4QPOEBsn0x0R+BkXCJETVgSkYRXmbtkOxkcfB
qmC7IbInuelh7f90geuoMTSHD5g+Vftw0dnqde6gmjKt2/e1d+5j4YKpro7vHh0O
neGkEh8GEpncrei9cOTbtjDM4enZof7bIjVqFNBFCLqCkcbDpNXoIjjyY0/929de
yDw6NtovrP5Azd7u2oC3xLDIis8JzggWJ2SUbmKCd+kAjnmMB6SuzFZ8NWCtJP8J
bJ4/VpJAbuggH39P40W/x1n/dCiWyIA7G6YeWicSoIfgr3jgsOym4SOu2v1VSzCX
AI2GbeGiLZoDECF3jWjhambK8RfJwOzg/vHTf0yVDKinx/gpGPTFd2lNK3iE5hGO
WpR3Cnbtj4ukdlLjEt8lgIvFSMZrL15/qkdek/t+WGHAkh5OjCysv6KIvnntPMsT
R+p7qnalSTOHF2/MuLgLacUkiq1up7qUoiSxdFnhXCHGKS4ZeySWGWfk+oFyIhLB
TpGR8P9p8ONhyZxOZi5a7Zs1razjb9qXgUaUmfP/cRnylc4Aj2NGzU6Jrf1a9ppd
DYWFEDlZI7bGHafRA9mbtEdHoTPF5YISawyjwKygiyacW+9mw+fz687cLIWOViN8
KiH9yPKOUo6IaFKwXgZ4OImFR7CRPfAXRYREb66wDVbRdqjca8orX+/7UPuuT+T0
Y6qXGe83CQktPzuU6A2spZhoiZa8cuY9PnWWd0LlGlP8Uv/TPK1nam7WFCkBPJL2
/UGPbfTTAqblYpiDFlZyNLlqJDGYSLB1BXYPxkxU8vMJ9xCxz3MwvP1YVRLjF6qg
iD3MDLCWChJfMnChq8iX32G7qTb5qajYreRV1qs8Nv0JhLjM0ITEa3RDBTp0t3U5
lxLOXSR8D/5MGaY2JRRd6b2/Uue5NVGU67RP/NxVE3UCyKE4fCcE0c3fhk3QLry0
SPtZbg7HFFzOsyrc+Q1VxJDz67108Qj74lhqZAmKatYOuhREoPVWVjpe9gO+ILIv
uJpAPQMA3U6UEN9DQolph0PhKCZ3Ljcsn7x3POeR5xjS3n92RWyJpgqGiG8ZOMqG
U/6jk2iCTTW/5q5bWCzv1Iu+jvBoMo39sE3OJ+mlGSFK78FdI/Mebv95n6AoQhDQ
OdWozXffXRo+FnTef+HA4TveMXuBA8KXTo3fkgrukUvc+D44YwhVAlNNVbrMe1q3
WiAabgvuJC1hmGaxyfdCBO05Bhs42fkLWr+ESSjA84KCCqc6gFJO1uJpeiPQj+Bq
YWnv53I4AWHsnA8Kg+ScRmMjzDY6SYDubToNylnM3fVCqCgAi2lvIu6Hzy4zdMuT
X4smiT5qJfIAfD15KArYTNkeJIPlZ8+d1P1bmmKbZ+bRCKvrlFbV3gumzfSMrmwW
Qskuo3WfcODo7cWMuJUznqz06RNje27Dyuj/l3MECWPClnuEAI1aAf+wXur5pRPa
FWJco30B80qgsML+KOupgM5lWncYum+b/+WJvTef4dsV0EapSk/YhtgANMvKfeG6
9ZLpBqvLs+jrwcJhne7+muKkC7Q0Hjy1sl6SKQxxGFcW3lNi2PCY13HuGNwnNJBz
rd44uNehpQUG4LqVlw2Ldjggdm/NUfvt3Cl8+fJAphaYueow7Q88idzadMu+DCLV
LlmeA0nim+uA5jvkDKAN5Qo1pRdzfgg/vujLIVzH9gQCs3ujiB+PChShTN+OArOd
07a0Q7TNzYmL7ZHIA6CevlGI61tAFOwvccM2Rgos/Jwzl0B1VIYaPmUdbdpRA/W+
7hySIGuvjEIWnbTaxkvu2QGArKtHZbm1HY3g/LIH+y6QbCgydUFxaeLIV8rTdK6q
D2zq2wcJqSd7MFbHISxV4my8X3pG10GdOARX+G3mfYCGW2/dpG8rsmT0WKXuEr0u
BPdGVnCgphcaU00wacV77SgXIt21aDpn8PqBK/tD/Lhv8VO+YpO5vQ3NEqeHC/I5
apQ10LmP/I/XsX9YLYvSaP0CqEngHQMU9czb5ToS3mfe6Chsk3sFNwFsDY0hpI7b
l8bp6J0Fke4dvZnT0q7837h5QNhG2gHZOARYY4QeMLtRt3jk09w4EUuBcu0vsbEi
9zwuJ6rVbA0WKdIU+mkZfoeta14rfO6cLgcTuMFjyyf9UQ9MPhazpN4PiTwJkfoR
6EHuMFlzSv9YxJ4v+UYRvmnfEWXkCjQIltwnKLRapPHud3k3D6kWtnXpFiVSFXRQ
s+TEzClWht+8NiSXd/5OcVCEC2R1iMsKWdeUVLSItiJN/hPQefVx7+l1nRfRkZpN
lo5B+rm4CU+Bbg6s7F1QoVFG3YIkpwpSlTr+1T1Rb8hg2BBLAaYbWKTxSniK4s9G
oQ8biLIYCxhRAUUndYcsbBQz5/0P1lf7nGfEXjihW37JfXDdEFdEp0q6hy8VA17O
mA7rhs5yQF6arBnlEML23z9g+mSUPlLsNsxvvZSIzCBiZthM1vyKjlNHya2tBNmx
n16qQiqWlbhj521lpncKjnkOxWPGVBuxc6hQXRupQa/fcm3k3EQLTtpzcorsTcDe
a5m259LeYGLJpFkDxy6B487tpEc14mhGKlUBQtD5gFS9QE8orzKit3eReT9vnlWG
imZ9Chv2b31Y2XrXSRKBK8DMe8g3rRBZTH5g19ByD+/qRpBKdbkhQnU3hVAztf83
tNCQnjjOpqhzK3NPEwXQ1eHM9ZwhVzt0x2QuCpBonZjPfwyqQMJ4klUzHXvprLNf
3oNeRU/Di+cZKuTi7BAJRk2LUYVKlXP6aAZqKDY8Cz2HKPmiEIC8PyVoiQ5sr708
H/opucboGwzqYECSWxJlcJk8zRGV6bnKxQNRkBdiK5i96S71G/zLw7UULxMysbpD
7Qa27DSa8AXfRrVDWoQzKtCC7W6LcLnPefJxhU0IwaaWom4DqXid0OtkaOq35ERH
CcNsQ6tTg6KqZm9bY9HUR8bxiEy/hiwhE4wijRgLX7PSSyHM5HiWEs8VM8Vbhh9D
H38yWq8uxpK/4gy/GTl3fRZuYW5r39Oxl5cE0kzbz7tdxL++3W2N1ogDTkm1JXmO
tPL3lgCkb22XE83HhSm5I5WLeGsTFk/wBNCUZib5zGPKS/u86zI73hgl7lKh19k6
jZyiM9ykCUJRuBX0dQDI7uCH62ttS19JLRtarOOWkrShSDX9+vTs+4KJYkx7gKFQ
7Fl1P9ms8DQU1IL0bjMtC4CljK9xOJ+c7KMQnGR37zFPXvpjCWQ8qC3Cay8uqgU/
d4T4hpdz6Dxs4PF40ljTW0Dtd/zygYjWOKpcw/P9E/aubghNi2M8pnVDuJ7BOFVH
nyFY9ifc11S1ktDmSdgY7LOID23y2TqBgAuek6VBp5XHYxpwvu69711fU8GTjWri
r2049UvrEqAlSTWVKi9Q62wNss31yMUSmYV1YVKjgTyX6eREUIjEndlabavd1jqr
0hoSy4bs4pv7BY3ozbk27kNxp3apHUCwhQbq/2crczDMqf8ypNaDJm1cKGR4Ay+r
h8xfYmuUyhN0VI3v/KtRuehI1BLeXIZZPUnBKoUroSoPdEsQXaFlSA9GVS4w/p8Q
lPNgtKfOP3DZcU2e+bTE9A5YOTPxYkU21TL5vY5XAI5ylMIWXA1G9Y+tGR1kQ7ib
ePQ5bTvl/rRDh7wWfyUJJXgOGl5aZIgrFYj351Gi/vmcYPzIBE/Z1FBGrtzoUF+U
1+TJT+wD7lVbPD4U+UmhgdaiPIibqH8WxHiN0py8cr+VQSiIBbWI4Rkri2P0aB3P
4K3pFUN4gDTC9OIur4lEvRyvNP2Uct+loaAz/XV3+j1faRsZ4aGefJ+jR1/vUzgB
qxdr8VuR+qGsFjK9IWeWgwi8RYzsHKyrAfo+Y6SXz76chQw1D3fXXQHOIXChQrX6
xdDitMZoO+Aq1brtI00HZO77D5az6gve6og/JT2TG9r8n0LA+xycs8HdM55DQUdy
JZhZTZmkfl1/oDuRZ1Cu2naUOft21yLkNRpgXhE4kOVmWa0y9JIZSr2aLgXELkTS
s2j76siL3E7nbz/vXgOdCUkXmRoqMjtjOtCSo4KH4nZU6pJM1vW0ZOO785WXV5mi
l7MbwS5iziKK1xv6VMABh7vPhymYlaI1G/sb18jAMcIYh4YHHGOJoQ4QtYL509ny
yPg0zLBmwx5atHQaNZMu5bkrE4qZSxgC71Jp9ooupA6iRJIyFbCR4jvfdj1N/hdb
16wgLXSWfsTHit4pvV26e0YHxa7Fl93ClR0lBs75Xb1SiFyQltdNpeewdfeo95AS
lDJfCAmc6dtZg18UKLPWMV83KSLp8rohN9MLp+QkjORTc+ECv7Xm6WqdXpexvUhJ
KTRGeqlq1zNCw1Hug0entWQLY2ocEmKw8cKbl8pQ9leKOrinZFWp8ouFxGrP53us
bscDeOTO7T+V3HEe+2TJrPPn7/M3AUUUAkp6cto2G3YSHg5000xaS2Db7bi1mg62
I5sTS8pxso5ZXdLLgMm4N9zGDsznT+3lsLhaSIrDdavAuqFzw8x2jg4trhxotmBQ
UM5rVivOvRzTuzRxju3j87/vgwogB/8P6HQK5Y2Z79h8U18Rvf2zr7jBQrA1fd9/
resDZ9YNjrAoTImYAfHivF0uaRZadflBLEw0xtce/ho2bbwkE3mgy+gAalwzCa16
x1kL1zUMm7lRPZdweHCztgFZeyY1sFZhQhAYURbh0eYKueTr6cW74bB9L1EWTGLa
V45FZ4NcO1xM6JvVhWnCb+YLSaAYvhjnnn6OmYpu0LkUS1zl7Ari/oRkrg7lJIS+
7IQHq2wmbjnHAoeduDFX2Dgy7yOODNNMTDBgmuKAYkKWzCg2pwgMsX71j3BmVqib
vicBDVp38s+PLrzCNvclfyuxcg2U1C5pqYWjGxChHesDZTglmxaxtk5AKfAIivBw
BgF/WWZAP2kI2jjMjS9arjIwSIMvIKZqPWpFhvsBpNihMrT99zSQ5asSEwYxIWwF
v1t8EfD9YqOhAaRPwQglftH/C2kEzT6xizte2z8ZWpV3z9rjnSejCo0fu0lcW+Rg
GmbHmK89gUDTvxYgbM07cWJ3baN+PWtr7yAeDR2nNsRnkcsGxufDBK1SydRJbyld
KVFKHgcRjxCU6Ml29wk/uwut8H+Iicqe5S/uZdPoL7CAQDcpSNXz8ow1Ruc7o6ak
wtsixm5jHkt0gy1sl5PaSB7TV4ccciL/xzt/0swrXIX5Vb/M0S98afhAMDhNqIWf
+bGcX2rRMBFfmqo3tmV9Jk3FBtlvD1tZqWYKYh+MysrOGj4iMx7otzG9Q0XMz/3D
3nafb/131G+jySvDbP8J40+vjDYzPoB3nHQnw3irhB0iOx61w7OAhfCBPtIMtlNS
jpGIpsXR0u6hiPwz/dYTPahI2xazfBybhmwIQ0TFyTenPmvKbgb4hNl2h6cYGV7/
u1jSjwMe1tZ1ZQbo86s6/diUb68f5GIpcS++rffbuQ4oHd/Ho2DOE+shndpi4h8a
MByGOFVYtUvmAa1FRmSqelFHpFtnkFDpeykHkQUvw+PnOfLCtbKtibHru/PMI7vs
qyq/AhoKyvIfMONAJ/B3b6GLbNmnZOQ23/er5ekLyzvqZdsTZjsEXzv2e3xcqcEm
MgfbRJ3S7feHY03NqCttElQbnNKQdz9VGxYy63SD4Lw1QEf3ZT32S6gJnrZ7WKug
iyhAF65/zXYVv1d+pIjR+Z4pOtmWs+gW7Dh7vnEKkPP+AyynUHhw4dnTjrKVanC0
vHFn4EVyV6w6zaC7ZbirvM83SbsxgtiJ+LQ/rDGmVjiFiViIhN22ewXD37tUPiUU
th9WidrE/wQgRF+EBm8A6uCZ9ziTkKrOvWFiH4hLw/TnPpIzAkLMihYqREtA2yiu
t7NjMZm6K1UZIT7nDPxW7rO02/FGsnWlD7BlrfrBIqN3/s8L2z0EbR4YmLitv8yv
d1oQleROEiSyTLaVTuBsB0wsz7J9p/M0siKxYaT2owgCm0hmwwqwG5P4uDJrScVu
4QtwyxKvo3yPbh47vVKHOgW4Afs1m4IDXhiGCBEyIw8MsultJClZFcRMRHZQT/mt
S6eyvnS5lm3f0yEgUoOh3QfLGKfyJFQM7qZjEPy/deyq2wVePaUJITtMCC/KMccS
gh8aebRHMp6REEOgl8+AL/fpU/fAs9hYNb6p67E/DAq3sFlaDULPv5gsrdm3cJPz
ATQ+ZUolIrAfDf3N8Yo7M0ZPOLoA0uz+SF/kMtSbRZAQ7od5De6nxqR5TRX+V1J7
pJI7TQQanCMCCI/sWfa5zqYUGfCAbQLUb+kDbCzYKtUae+dLhrsIosoW1quyspuB
8m3jOkLz2Xpg8ff3MEASku9LQ+mNW5pKqRKSfExjv2bo1vb0B86/6uCHtM4ayYX0
HaTXPHyz9OZsFk/UaGdid1ViFs7CWrgZR9tDaaCS5WBF8kT3iATzoDI2EMLWmzd/
CqJqFakDNNQ5uNi0ytrxomPft12WWwaCCj7RQ6CwKn8PtC1B7A3la6t/jZ+EWsQK
iPDXMjamwWPa+2QfdCiC1mcP7RIDBnjyrpTGh6p+IghKcR5EHyqQM30kDKnCyvAk
O4VZ2PjbJTydqjsIfQ4rzJ4dNRPlfREAJBOO8Brl2n5m92oH7Vn2rV2x/iKXHPle
54olThFl0us4dA9VgszDOVlL0E+r/RzfglA5NtX9XP8sJJMkpUsm+Be3GHSYranx
WkDAvdALSsq59Q5hDUfLYgY9ipc4/afKSaMJZ/RbuqpZ9Y5R+4QPl8ZCamNJV0/K
LMlIpHhbkEBCUNIkLRlueKJFU6aUruAGkM4bvoQ2fRLUq379T/Z4i5Y3OE26pWRz
+jnCzr+nqkug+04fxvnXfI43VXP1ecdWfYOmWsChbM2Rj6nBwEzbVChnFfQNVYOo
J+h6YR6D0RKDE+OCezVMwjTBUqWC7sCSjUDiVaqOWkKO4tmgxohk2m668ULLkzNt
1m4xtq4XTSi8JOsLo4M03Gw0xTDMIfrGmAhu8sSRNDtnLekmDzMF+7jzdgYpjcqM
5reg28bCtQnfkfYJJCBmTuuTXZUpQXGskd9mkM9S1EGT4WabVJsmnGGND9sTZfLs
DwQFTRk4fNKq0tjD4vRMB0lGbyRTYUOTz0g6izopejOg/UJSxfajmxr5LwFp0S/V
xd75mnasUrU4QMo5nYn53DakH7ZMyqU+zWEloU1DgnNYvOpGkr2jK4bAeSTszUYp
04dOZVB3HRBclqCFBegLzEpjBNTG8uloCLvFg5i9dcl5/TQH1v0X+ix7grq4GY6k
h4twoPo7RWvrJxT0iwzGG3qmfvPi8sW09ezRVbvfd9PQoFtxzAcjXTJE8/aUYRPf
24hI4LVPXj08+5D+tcqiVE5WK44KO6Ji6qQaY/gJh3VWShOAhdCSW8GkHYKxf+UY
oYgIRJqDD9r26/NeO3AUFFOuxm7ouS4ZGtBoGg1yBKRvYXiqJCKAZeKgAlEcILOQ
LGii9e98pOSxBrNqDkbFkbV+UG+4ocJ+p2HNnpchX7KhSGfgcDkgZ0GmukP4X1Sy
SKx2ulBtlDo1dUBbM0AULehW1RGT/xkqPS4D4BwbSMdykZvPCJRwPjW351hdCayk
s8hCntkXGB94m6MCt4BvUIl5LX6DR05fymIsRxzqMR6fnRcl53sMi1iud6WYu5hY
rkDtOZwNVWrNJPovAltDOXgPiQwoRZ2jGEogaFa/FMBpxBTL2HBcX0+4arFgG2Db
V1txbGSeL8/FG+upULLB5MLLpwM5NHjiFvJF5wc9C6Fn45ahOfdqyxYaMZ8HIwBE
xRWhSRXQrgs8cFIEUVu0Y25VdI0c0uXr0MZWgWZsvbMJSYf0aui+gz5ORKZcsCPw
6m06q9sza2UE2u9eUqeI2NGAwol6i+IXfhvzvit+LKlaGrwhqOzj2iGP4ZkXsEPW
bJK/u0qlzypn+5ZZtcaE+1MyxI71rLgj/Qz0xjZHjIeCu02yeGM4Aa3Lr7iWomlL
+nNImPpCigVvLEB4R6iTLLyPrPjmgkZcYGcXgM+zVBP4puHZpf/D5Zxvmyhl5zAS
F/46KIlKG+9Ka+8zgVdQeAB9nDRUaaENGV0gZ2EsWrojYeULidL/KPwA6nd27UbE
EFBrPYwHanvuWP3QwR8a0Qtv13Gn5HgEE/ElzKYnxAkWZPUuHnmyi+2zNAVr5iEd
di/mgILuzXWu5TB816y/7t3bm6fXe5tk4aMH34jg/e2ILaaCvGP3HdjyYuKI9ZHt
YIHmddeY/hZeSEywFKZc9RxaSkos1gxcCKwg6CdPs3nxCtuni0hGAGP6yuq7gIc0
KcgOX58xfbvk2OOFrU5z8pqP/UEwB+3BWvubBsFxOoYm2HKbQtcU4TVf+WtfQujs
5g2tOg9WzWRFshgIfNp8VSsm6FjTFOfOYn98i7vQ1NDILtGmHoRUs4x093z3kk/h
YibQbh3HswwB61tidxolyrNOPmbXULZ5LE0MAQHboZL0SPCIBUAMIgOw13YXf1r5
DyaoCj3NNmQSSGb629ASnLq0eZbfZ352jLPGoBuG1NCYy9h/i5G+3fzuC+hwFH07
MyC9DlJoP8LOC76KYzOOylpCUNf98uKNmWcEawnJLzrG9ZFfcbAAHBH1SYZvMHPe
QeNXeEF6XiW4gpi2XjQlTDk1i8wHiddpoco2X70IAw8LfbGbl/7nFMKBUvVae+Co
p/HWuX83E2GriVcIhCTxib6wtCZRDRv966V5ebVbv+mWJ1O3l1I39LrPKgUo/6dW
cuOgdqUp+iWxHjw60GEAt1ywZIUAtA56nv9sgMgGiOW7wW1H/joAbPetXsvR0GY6
312bDwknH1uTk5GUWsRpG1I/iwnqxgAm8vgDBzeovLE7/R0H0iP/3NMxWnSHCWlD
zbvRtdtK2H/MNK76AXEoouvY0x7DgNhKpEfjEktTu/KGwmH5y64W7Mvemc9P9QmF
sLB72zsOEgff/197qNrM2XijYA0NmPomv2Of8mXTqdyBxBzAMPxkFvsfVPhxvExf
qvDr+DU/ChSUubGcLJ9Fkh9QKSzIk2wc6GAU4Tu8zbJpAz3BI3Tq61LrHqNFN0eS
D3TzVerCYK/jORn8Orz7vO7/Z+0j+t7ft1M0qhoeKz9S96swv7/QJkqGVETOPomS
vbFq4RIn2QOrcRd3m71OdqopRaXXlZAME8izA3DuIaUXmlf2EqA14Ac6zhUKpJEX
BBLgVVSfjSzRgOuhHfiYCa7egiWisMvD2H8DvSQFRZfAFss7nPxypREboIXA03AM
yuoEMkKYYV02BW+bdcILrSxmC97fr2TfqidrHfjP7Afq5BnrBpsGb4SKW/vsJq2b
PVhlTc4pHGJQjSfKik7N2RbSRORDA5equMj+Uut15xszs+SxlGqk1URYuDCSGTWM
I9vrPYyIPY/CR6HFQrYHKN5IU1SA6K7Ll0HhCEcEakJg360CHM8S7DjyD4AYeOyp
LOJr3kELGQOJfQwXM5cMfB1vi7q1erTOHU8g9QIFtWDECKUYu2DHI22VdvHd3cEa
MYBsbx+hdO65WTdgYyD/LU6SI4FoVEH47XXodUUP6NBAz8OEwBjTMIzhbjoVdEoJ
93FqdrjLqBlXpdQk+VAWnzrrQalTXcySG5BUMUX7eLWEfTh+zQ28so5WIDa8WBJn
9LUHLbWjXjVrs9B1zA21+VSLSFuAm4WTP+JYcK2DtBquLFfiIEgi8jEnr/zNTqTC
nTtbThMdN0nCHEJgJS2kSsN8YQBMRYrwwqS1wwCV6OKTqGcL/6Ws3IZn4CewuHdz
EjMcSy+5lPySZH+dE9NaDPwjl/X5PcIat7GKNyJYMAsWpQO0t9jAECjXKNpulFcI
0XJT7YT8vNI/1Khq9XoEPQcPBbuPH17o2tIYqQbL9wDyrp3ppCi9dIPR4wgcCGZb
e7e3NUkMtLB4M79wESXA32oe9UWd2Au43NIWAJLucxnyCL/nsUM7famH03NiKk9U
CgIbQW+5/p577b5Bftz6tKG/GWUrpUzt3RGXRHHzBHcSu3ltvqSzwZ1obHoDQnFF
IyIVNwbNbO34zK8HIy1Rh3K89N4UrguVhgUo9NXJ9rENDUk0P+coGIBSntwUxYcj
G0g6F4YGPhkEH1Ch/DZGK25YPkI4VeAD5H5mXOD2n3J/Q6OgBPZ0AHjnZU1bb7HX
XqAJvL16l/S6eurUhrIBSstb+PCVs9m0bKB+uJpvxiaJUQYYCXy4bU3+u0lpzYli
KSx6E57tiAkZyNPPzCLI5RlXFrJSyjewbhdDtxsJs7dZx66O4PXY/LnUpYg5GxfV
/GMPkhQwr/y2RVdgAm4BrwnFF4DlpkISxdXaFLsB/9TbkdG27b6CClASeYUiR9NV
y5K1zxSjJX+gGq0pdhxOhgq+P0TIOkgm+R4WZNzQLOgvT+KJRJVeulhLaTJW5Bwv
UUXPtYFKa6hL4anPGEMaVHYxiKZDWxYq8r4sBpBAd7GShB7956v4J4EhNaTdWLIi
WeLc5CI1FzJ8BYHcp1EG7SfkNr1e4OJPToScnmh4fyL+pRwUO5ga1ZzEJqT6RE5m
E16L2fHJAgckBYfi0DwGcPf/hxK7faN7MELdaIHZaFfkwKjbz63Jq8ZcuARhP6tQ
Tj7NBMB2rY0fLFf/AkpirqdAu/YrJj1Yb9kryFHOpGcgkXmskfE2lZbkZ386OyP4
+Q0CvxZ8U3vx5ranDslGJWXgTp3B4/Egl8IbUm94FtXhG1RdQuYxRWBMKKXNinWa
/pTMf/27t6wMl9kwXHPAmSlgs1AcZpUnlTcQ6VIrajd/0X8x6JcSyiSCHn3e9E7J
EpHObT8061A6J6auMuuaprQbUzueQF5WazTmDV/jR4tXW0iIC1nVwsPqflWkkm09
Rj0/4VGdlnn6up0tdWGd9EoyNbbPKor9b1Eox8VVBQHN8jefaJGmOuBx/qPuPD1E
8hYW16Fo5FXKUa6vBN8KbGPgI5DAr1034viiPCbXP/Se0P+YP1yNc9ToE1nLmdKC
KnrqcSgoge8on6FV95+Rzis/yqqbJiUjC7SVNTJ+u411fcouV3oC8sIonNNxIlSW
QJBIBy7HJlbgXXsCdV2V4GwuCAo7y2/AUul1x2ohRNFCKD6Nz2N5w3CBtWTD/EfR
ffhtSUPLzZvE3s7jt1o0cKF4KRaZV8XDVsmST2vAqVI2z/ImJYpuFppEocBx+WZ6
MJ4SyEWFyP9kaPjXnvSnbBE35CAskbPeMoLwmN2UWwS609J9565XxV/u71aTXqHl
iAxxGU/QAEuk60nkmRVtwdhSBhGhEoYtv4XPHrAiNCsuK0A0O1lVb78IwekMUmMo
KW3o36CCEKBhXPL+FwVY2xLJGC2ewAXgHmvC2+uxn5tifULdPZadzcOYL2PSh3ro
mvXHqMsqQhHHxJSXsSOmAngfbrMgUKNkC1WiurHQCEz0qtw8ETHrOZTj0MdOx6UD
kO1i5Ip7YkpAbBUmWwg+mngaKTnJSuEOvZchgej+YXW7V9zovV9wmmAIZPKcKFM1
UDGHx0dnb2fXVMnyMlEl3ViLeG87OenFGrtqrXchHLKymDeVFnqgnJ78m4oUAlv7
v+TgZybgM25Kv+zOdtz6Qa7as0I8Cg0VLjWdPp/gjcPE4kbM6F7n79gJP94eMXnD
8AqFhtgHTeAO2/sqgar8spZVNSVZ403uSKkhDe72AO17OWcwaeDqTuuK+u3OHIEw
EkcJTbCzLd+4n+91asvz1ZVQykZ/DwOhzR2VARV2ggtuFemPqHgMM+Jpj64yaxRS
ZDmnlIVlfVNPzn+r5AuhuS2ipwxDl23y+oO+U3a+k2xfAS9dYZLMBNJoVyw08eNQ
rnjUkBKZeDfDJ4IaMe9cy4S5phGA8eYmr+MOsCIX8mV/l5WO/bCJm83qbcFMHd6m
DBaKMWmwrpO6ZxhFe1K9RB8FjzdA2bPh+WmMKNdFFHfTKBG0u82dFXGj32lNIsgN
GiKyil6Z88UvKfF3RPu+6L9ubUImi7WHnE6tFuF2K1enAuSp1UHELovojCTuttNq
v68HyPItpRkmIehFGTOpepnIICA51uQe7lmd9Gq/gKF8pwqKYhfFwPPy8UZ3QAEj
dupNu0aUHOKQ0SRoxXuRJol8oQMsO4YsohVMHv8B0fdjmistJ/j7AToaar+pwVU+
cpMsStkYutleIc8oT36W0DztWUU80/N3prKTm/9tGji2hmWYdQcoQTAAqb0q1Llj
5qA1vENphgfUXIT6t6Go2busVn4qlLSraO/nhDLdOi+wYtY/fwvXhbc7hXwFfxN1
xh037DW4hwu5n9zL+J7i2sTqXlcHRS4v/ttU4XI/KB/gysx/PCJ4cx8KuQhapsUZ
W97Dm0mFNVtH03aK1Bpp2My7D1AXiqitEji6LMQUZXA5sbkjD1cCzmje2iZtc3V5
SdTXzDDXjJrVLT1FWvErVjT41u11gbq8j7Ga25Hza0VKNRPsa8XLpzkfx73eNKXt
o6eKtUPV7I/TbVTsD/KD9tZO049dr6XoDhsUp/VWsp1IOfqNrkca5MLvz4l7TPqW
2A40qkR8/JL/M0BbtYZtx4p+NBqHEbMUTlJ+pz1SjKp5Hl0unzqgmU6N7BV0cdSM
I+pBhvh8OB8TNgYzOHMrgI08tlsXFozGLI12E0o0I3gx4qP6uwPU7yTCF17oIB1q
ARKIt2s1g61YawTyiZU36YAKK8vnS3/EO65ivOSE0aDPjSuwTUg8SSH15NY2eYwq
Xbe5vbeM9w+CEjNCLvBshS2G690B5Di67Oe81p/9jPniSIUPsJ2jODEpT66EaM9Q
vI21zpnESaPQ9EBdSGVUfcoWMVJ/hc6MWDGC9KrcIEZDeCift9/RkZl90c0ZBLp6
CtVAOv2Iv5Rbsm5ynayQI0likaC5EtBqetp6vpRys/NiN8GXOfpfx1D5vh6ex7uk
fendYmaScRmxjTSV7v+9wGiEkqw91u56qTVhBXWWitRpqQtDNcyVdwH+9pBTj4Wf
3QnBnDn1WIvINyrg8+fYV0HLd8U1R+GKCLDSmaiqxFA69TMOAt+sLy0E4g25QfAG
Fo+xGiJcp5bGz7GLraYiO1A9Nd4Uv8LlwHWf0DtkUwlB7jL0uyANMGnBKTkh3uOi
osabNUtx2IPh8JqHvB0oQcLhzWciF7wFIf1Y+hTrbmN9Oy+6PB1XA94Yc2zYJ2Cz
K/ZtdCkZdPsxuagkAdlzgWZC+QtaTKvey4dmKIIj42ZbzWgTFchDi85jq5Kvt3D3
39sgm3kN/3bLuIlB44r2hOFkjuIGUfnWs24m5P+QP3jEAeJDWXx5S1xQnjdLX3/X
K1nQwPnmwfBm7/S6lH0bviLo0RaIJbCDwJszGofHNwiIM01UO46cVgiEHQTBHfzT
q71SLci3h5EqNquDt78RqXADZBOQ6U1NNK0s4T1LQaRAz8eXtbI4+/y+tPUJ1z7j
O4rrtbQQQL02X7ycjoxzc5/ufPcjvbFZnh8opNs9bcQJLZatT88Gq7reKWDsFuet
0DgUmQWLmdys3MCIKGJCHtKJ2A04DX/QCxOBe9Uy5uZsMN1zLCvhg0kqG5yxSQj0
t8jDzGIItKVkwVwPKsQo9vA1JFkoavXsxwAXGw9ES3Kv1BcTBPZi9/bSiiPMe7K2
wbWIg7wBkr7o0o6YyeMigGR00B8QQEvAyK65INmKXo2rQ/3Y2kJm0QDh6cblTC1v
QhNftpZfXk9kxFtMe26n7+jQWTOU46JFAm7tnyYXuz5EMTzuWH+FsCWyzBzlOKhN
6QVVxkWZqPbLkekZO2Z/0JhzG0C/4zA6HNP/+rXlNiA7ZJF4w7FA8dzIukNEardl
i/kJtUSCl+CrieZfNG5+ZF3ryM6esi4M2YVk/N5ac0JkH5kpnnT4aVMf0cQtwWGB
eeLy59fw224Pm7lzX/wB00Ga4bu2KR3gyPZjpsj6lw0grxmiPk2X8R7zSIPXJs7k
LPg+cW1skh7+c9jj+faGUVGcdZPgDfK/M9SbDceof3ImTPK8JqZI7+Y+iK5ptJgF
HFtBbcSHT8fVBcq6f+r4+h250SAePPcYtGn3nRwhQZHzuzK5VIs8lQhkD3EkyNs5
9LaLXuBvyQjOF2rGRqm2R5lmO6EUPcVYfaPQIZDcXPeH6wN4BEGeDv1/goejfgsK
2AEZwA/QmHXgxFT0W9hq8GnYK6Dq5zNK+Abz4A2ahl0SXMWItIsdZ1gpgNT0xP2M
+4MuwL4bZx0SwsiTufRCweaWWrAWSGdSq7Aw/C4qLV5YQCzDHB5SKsoieAxkEHRb
4chDKa+NEk0gWS7rtTncJratw/3Z+66QxDRL5R1qeYz45OQLLWb1c34klye/GL3p
Dp6REGT69C91ilt+4RgouQ3jZwAuF00AmMo6mt0e87JPm0AJ5OPLTz1Mq3gcNDi1
GTQ5iBuVqEp/r6Dg7LpJnbyY+KMSKFQFzjPtfelgd1o7lA9XK1VaYv02OjX05Ucw
MHd1RF+oWXn6G2/3ROfx04B379lEUJeUP/Kas1ulsPnoOs9hJTbyeCBfCG3qrvSh
ICCABnW9HIyuLGxQUiVbkIZ5Eyq4Xx+3CNN8OvxY4naqBtaq6OseeNCg9p6GKL0W
BZAztB8SxhWyqvj7mwMy3C8Mp3KxBbmQnt3s6NwSfPfkEAp6XZ5+sedn5UC+zLws
vCdTqcqZlOkD8ArnL/Z/7I196AcjVw/Gzv5wPWKroBSkkevj6SM+n4EuX3Da2RrJ
f2WeGFYaaiWDorHxqZXzheB0nXbcoaxTta6YSHOVHN9TjjVYpnqxMRQVXSFktinC
MSH2MJUXfbtIMbIR2DuWrXjjq9sqbcVb4j2cZVYZd06JEErNPz9qD7aPo4rVgh0P
7YXVm10nmRdDirdlHiYpdzxbKpVVSQTzNGTzpNZIVhyxhDoVuN4UpEhrmhISYFVG
80byM9rxytpVfpHXWmiySLbIMuRtc4ynrgILH80SKPujZzD0PhC3JQpTSdHNM+wv
rGNiJtG+t7M5En+RdQzvdHSZhw7Rd+cYWrzvU3Zm8SDv+YddZSmnqSewJWnxE8qT
/o/CIYAALElyKMw1eo8+wb561ZOGaRVxtYHxoImoZW0uL5GHcQvwObl0hhh8Ach+
FN1ApdNJeVY1WzReE+BpazXgyZSCuPpq6Gvj1CQ1GylX+/jvU6+VoosK4f5XpTsQ
uALsdp8xxN1QZ55MBzRHE4JKUaPW8DlxNF6ReE6deHYvYmagCPS9OR4SLHioDBvF
DMaB1C05fpLOSTC/R/oz5hSjaHuMRFCYkK5Bu0Tg0gYk8MmpzubfMtD/btahoybs
+0H6Ls/Lo5os4MlGb+wKgOWVjptcjL77sSrQkRTDJT4h56PcKiq6ypoxCG7nd5QY
u5LO2hjyNe3EGCo5wM1wIJV0/O/7OPU1nDEVPbeeKf3JPCXgxfWnROWBA/igD8Ph
vYQwg5mZpQF8Y2MDkrlS2QCF6DrxqLeXvFD3KfvRrmKAxiNavY0/7K2BaPal4WBm
Etelt6iRro/jAn5fjDJ9bbXEyAwOwG2Ta/w3E/7jpuykFIUjbxSHH6x30/ExJK+D
gSSVShJ79ATIOmqmL7++bCo6IQ8anxCCSm3rovdCaDSPzzLZ24+jekt5DotAU1qA
JNCNWHdudEi3qR2Ja5hQ2wrapSuUqNs71mnRQKVYHvR1Hb5twPh95F3U/mWqhqLe
bKqobM9m+q1gqLZrQCXI7HuJQtNLRCZTqE/rt6a8hNbz1aiRlxc+UJq+X9AEgULG
XgSDXstqNG+sG7nKYvlF6lbxHXY8EzTXt3jbZmAezEnszOUFHjWLKgg8UKjfSmM1
/GKft4PtZCwgki/kua3MEJqRW9bOoRoCRlY8jf5nZLAZ9Es/akLGJ6cVKL+kYr8k
Sdh7oGzWoADPLTKvNqXLKvfdBMdzaEfNU7sDZC7n7xHlcOqNAgsleFpgPxi5kdWJ
Eaz5iFYK2n8qK7MVQ9vqpBujddsYC/l4fhOwP3KVwr97LcJ78evD2j8Dp3soRybR
EyrnDxNhePN780e8Ir6aKAfMXF+6tq1BvKhrL2vAWJ8yl2LXEb5GjBWHOLpcBgis
mSDTFcTbznsPfohFMj4kVpzMtiKFKsF8jt83++D9MLzRM09iQ+ifOe3y6qWMa5u6
0aTqaye4gp1MBWkz5yIpS1JezyUMCgJksBG8JHtZBpxbc2vXbP/ThabBlFFRSVw3
Gj5zFjQbgNeeUUnbmNTw91jvw2/gdlRyz5/INDw7cgtiDdcdScBo8GbRu506giSE
T7Mw5hlRT19WqVFNpHQ1xFiX+dDUDbG4rWiRwtaWJzJUx5162HdWudTrWl72DTD7
y5aAyJKcc2qqUshWeDBd/waFfZfS6GH/zFYhLAl7Yqnj0pwrsBqIFPPTMPe3QSs8
Ci1UoquLDMOAhoE1yoelWOELPL6qTizBZ9/UuPGq5ONP5DRoShvc7iOEbalpElW/
Q89GYpw9HuchJ/124PZ06yBdbL7daub4JtMzURVA3B+Q/6p4M+SF54pM9GcIBB4d
bbP23U8/yYDokvtvcqIRicTU+PYS0jITMzlTHvqeTuPw+yZC2bUwfiOUzg4HfF8O
N+8yiaUtyfrbJ4cfWhemMZbMNCTOzKl1s0P77OZkLAIu6TEgSqTOkEEsXmvwBPBL
d6ueiCnda1Zj4rwEIIpHjtmferBZp7KKoDp3FVmd+A3p6j80COp9nY39MPPWjj5b
N2nYRVsnU7XSVQ48xujvnrJt1nl3GhXF4UFMHr8yEe/DZSaXOxfRMMl/FHwLqEDU
4+BRLbVNSIjpMRcSAJE0zPQ94kOD4a2JAYOS89GOY8zrtoYPQ8iNfmJ97IYPxRCP
x3CxnMjrSSs3Truvnl193gTdcmatoifwyQ4aVPQNE6cf1g3dlHviMN0iPNlY97b/
qqg9JhpIeafvRuromxlXfeyQ0jucKyDguhk2EMatVjrWURMBPWLNzgOBkfZ2Y9VO
uY0VyPkexmrJQlfTQfpqE8tX4Y29MMd+2nYyfE+syVVOoQRQwGxpxzrqyWOEENXQ
7GiBAADnn+QBzzvCQP6VhzG4EpGEcEgtmH7fg5UvmHl7KHS6YsAk4YhgnUT8ZdAT
el03S58W8Ss6W7G5jB9yuBO5TfKuTbO9MzFIOXlFDZ+4H3BRnbyNqoNYSkJV778w
Y1EhiPUr2gdk8P9N38dZOOSzAi88wRexiobGFpKiggk0G6ISB68mERaMs27dJksK
q5xsqLUP8bvZjHP3EtnXeMscgt9PN8MrkwUAJdHCpnKjDxXbTgTNcJ/hYhCbqcS6
7ID90mPIoSGMl40W0dst0adDri9HPAaQ0KXNtKUZrOHhlBQ0cCiELuavCGZC5r7F
QYh6hJEGM0Wo3Rzbnkjh6y0db6s21Z+y4a5ZaVtYtZhMBPFW1fv/NztBqDVCYMg1
LVaZHJsHVsuBgmDBtEs8LcxR+vpAhYxB4MUc0M9SRSQbWLoSs49Py9g6SYvXTH8v
oWrSEf6nZJq9NS8blxrmJx9mON2rhW1Tu8SZhlvMRx+hgQdsHwVozVAPRIcQbeWB
oqADftepUPnHL/XXzj7Sh/Fxra+aq1Xf7eMDLC1r4MYASLXjEbY6wnF4nSpHn9Zc
pAhTRDJytgRa5P9tLtiGh5VNI9VpVVYk9mVq/TMfliO/Scw2fo5GrQiIxxPf0RDJ
xHClhgoZrQhXYq/1e+zFTzEkB1GzBJotpTBoDkaU4eMnL96f/PRLQsYMfZjiSS+N
UgrZB9Ds63vUl1n638KDeCqmnMwmj7nHQtpr0ZIlyIplXEp6sup3LQLqH72ePMrP
sbBW8LBzVudFy7EK/TqvgjPmTwj/vk/x7KsN0INxgqEqT02VJkJdU0pjq46Y/beQ
3lms6MB2gKEx4hYroQsXPztBRLrwUgm96KCXEPmDRod+DhaDnqhKxATWuBr2WBDX
bUN2LnSEqOVr7FdMAvNPhcfqwRSR/0o8rs3TitfjDql/TgtZIxK8s4uHsdzeTOGi
ChqMzeyfBr6ki6sKdeVGJjJIExAn8Stq7obGDQy33Z7ceFFgPrYGfZ+Rt5Ph2std
yOpjg3ynkaVuLzj4AYI4ObNTOr1wDbVnFS1JhI8stCoTKQk9F7Jp25VhzF7mciOH
qMKqTAcoXkLV9u1snCO+fJGAOeduAGFI29XMMtWQ7O1YawQGInnQPZuhKX7R9IIC
VcAbYCAr8F/kefUxaX3hfblokhPNY+6ek0bWyiWsTi/kR3E9COrZoLxOsnlcj/AG
SqTWe3fBUS0euCC0mtj474pRN0YqRCVk7KUlYcWbmWTSgwN8OIPnNwuh2BwCaMEo
FWmcQ3N6CICXEnlnTS9v9C7eKeyP413FTLoRj6nuILmKf+2V6RyznXcdFB6PabtF
nOJuUqn3cUvoMwNgY0lnvIh0t47YQTt83EH8xIbjHxQvYh71ENrizH8RZRNxb8B7
o80IS3Iq06Bil0yHuTQUNW84EV3cbVS+FhAPQiRGjlCbp8wXOaSu/KunA9l/sVJJ
X97uX97EEJb3G3MScZxhqbt2fKGBTAVLM3Nc9lwfdcY+Wv2HcRPR8JBAy5NNpZCo
84F1t49K2TJ3oZUDO5V0ZphBeeAPTjdRfBFNZqB9n89Ark1hHSra03KuNVKlGCNB
2s+eyIWQxl6pblT0k7x0PAUs+0ZqHV3VehZgP31uLqLKACDRI7tFM/2551Nacrdu
uXGLUe8cBxFz+5HHCrbjJfYy89RV7iVmzsZbJ8BJhi614PJ2elUpZMlW/kmPCyyr
0I2hTTqcylUNfDVhQ2zVkHyozonNnOJyumzRC0R1tadiCB8yv+W1tIyKWtFJa0oA
lwaAtL3Rgjuj00osHUztIPaTLGGi5Oes3J7WLRc1jvY3VzPKE6ZGrFmEkdDQEXuY
MMXTmNiYvHIon3VP7DoZaUvGB8qnJeX2/dOnMHqOoqxXC5QQasYiuvFpdvqugvr6
DNY3x5edMNwAAh2gCv5AW0V/kCs9gb9mglQh2NTrCkRmXwnMNBn6qQ3ADhaWp9zv
jSiUZ6Dew5/gy6T1XuS9zfSd+cZtPyFLSR5R6cQ0vGQ4cI2YyhKXNT4FsBH/T9Ay
gjZVGjRWySHnW2BeaK220gWIA5l4p3ydQKtt1C21xhVnhTDAACvC56YNEYXfQE6A
2NSTCLlrxn4wnxXRnYcG8bKes13N90MH6W+ZodKirDT62GRlj4H8GlBOM1tZco1P
bJSPljcq1wkcp2rY/F2waFJTV9n3Jbik90Vgx9y0NfIxEhdUsW/Z59OTgHADLuiI
iad1noiqrmQovFV5kDJ6HN37/v+OWfM3EHQZoY+x22x0z/4xnqeh2/aHOQwkifD6
cd6pb1La4rja0jopVwpjLoheOPWSNcGGmz5vzvevoUwn7GWfmMafbxqBFdZhJD2V
GS4g2b0bgFt9AO1tIm+LvVMM2fSjMoMX3mDojkq6XLuM1D2or6J8V5qa6CpzsDsQ
LiBK8wmgaqHGadLygOHwRsGZztmgAbtvNTDbThgOCi3X3Lv+HxAPTinZ0D2QLXfw
oGV831BH6j0MLFieh/lhlcABh53pjQJnAo9zjmEWV1jMgVizROVUulEm+NHvWs6y
Sf2CsBBAdncHQWR+WPsBbK6r3NTjJrlOpRdEPNRidvzI13Vrm65BHX+Re8zcti4A
v48oI7bipqpA7EsGKYWqu9A3YttWq8xjyC7wACYSXzX6+1XVGj649z32ranlYmEU
m7EquUp2hy696geMOsyz4KeGTN5cOxeBE00mGm6Wf7E42a8HB3LTAIonXHOdmyC4
NbWyb+q/PrnIzgloQzPz5xnTGNMEpW3mmfZwEVewz4XsDDj8VxJobKWd+woaMYP3
PcCbBaRKYVe+prdw/aQ2G1ZsezxrZ0jZTci8RUN6zfBPfUuyGL4gvfp3Itw9N92n
23XFm+ICVICQe8mXNUoUTGzHijt2UgTCCQ1a5uNvx86gDakEY8JoeQHlMVOxY2BY
TdiCxPayVh6HnKwixFhM5DudAmr9jyO7RXuV6au8/xyX+JE+YAPA6T8YjRFV5q3B
2oQLHKPDUGAGusRXBU/RuV6DFrRpCSfEZf94JHmYHXdCYMAp7h2TbK+iXT1qieQK
fHR/OIVat8ydobiMrodwmyGdI1HoIGcb6XkyfhXjxyLom8l7iIky1jQwqTNfB24b
Xs7htyWrSAEcgnB/EUVMuuTRTtPHVEdExE/jJ7GZUoKOuWzFMWIm6Xpn1BTQM6IT
89ld+Nrt/LbDre8Z5ehpR12fg2P4p5nRB0QO3EKyWGP5OSNkMmZFxWYviywridbF
UdLMgJq7tNIQZU0q9t+PmTxKn7OmTm2VvEb9IIXbmsLqtB3TvjbKzRSk8bC1SBzP
Iwj1nUwEUZ/4PU1HXiOJdiytcDHJAyziVfly6pgIcKGvacqLhKS1pI4X8i/WlYRD
WqZVBT8mrcWcpJvvAoBKG3GphEDKU+SbLBKtU+tiErgMgmgctlMYgrj1Wh9y0D7P
fwl3C7ospaW9+T2rF61g9Vx9XYVQ1XApQjhU7HMXirTOHmLjNMQEdoGuj1qGZnPw
SvOxbIUk1zTGPadtwS1LtwuNj9ZLPOe/kigw9k5SL74B206stHtVztARggUm2+vg
8NpgqM8iXyj7jlWhTKB1KtADX6XhH1vIEQ0EGGUMSaC6yuhirCn8Y8H1ILE2ke8W
cM8z2Y2EqXvjh9KsCk55yYyLca1Hk6QdKfYjOdTsUqJnHOnDsUU7zLKB6Zj3xIQJ
+0HlSMjRJgxSezxQbUEOYDPSGdaJxLoownZlZe9CCtD+yHgCwD+d/PA+gobDILi6
IlAe0asMzRQda4OEeLN0MYKAxXYYLVqanITD4Opc7J1Qx48WkDUbtbD08DKMw+CE
7OdVWQN+R6QcM+OWTnfQoKNXS7SfbfH+12iN9nWOPGmIbolWpM8wAFUR/WBObUdF
IUEy9zVK8GsAyE+9Ct1ZPg/QA78TzkCZOjNBOOkWc1BSx20LnwDr0VLiSjc2dPr9
TV6MStzDKMD60X5s3254fAzErrNr8VI7EZE/rkpURMldo4IZ5asq5JBPDuUvXO8L
c506MSPGB7tRcssLsGfztvvPQfA7Ge9p7z3d9d7f/m29UoJijrwGN6GdnsTwbF9D
zlXihxeus3vWNvhoAvIV6RRSJzYGr9C5Phtb3E/25vl9atnSU5fpECmLfpvSLGMM
3lMjIT/V1gcDC6I6LyRFBFKVTqsyPqjl7mZ9e+p1MHZBm8jA4QqSx1r7EMDTnxYS
1nisUEiqCqMUlzCJB+Z50Vbif8Rm6d0NO89dUIMy+MW5foKyPwENjHNrWvCfmATL
zdcJdz6qajn4VD623N3GZfNer9ExDQg9BsbGIsjAHFv28v5okbYAl7GsCQsr/GD+
HX19/RSB3ZZQKHpDcc+926Xh4zFZ1czLBWlAtdsaD4Z80l+gCZgRAY/4O+3XwOxm
bzm3V/bD8wbMiAhoNPwxT++01hqIVlYRbDUq3LN8IfiRUej1CymPdUEwLFMTWZvq
TNmoj74uM19waZ66LktcY7j2q6g4W0u/UBA0IVRkuigJ1wui/Bfqt4Xr8JPb7tTv
2GExY14oYTKU6z4EhSPjkZYGTzj6f6u7xWypQrvW7xr1+TsF7R9mwwMcc1WvZKpB
Vj0dqQu44AEyQa/USYrjZ4nS4vkIO6Mv1cKLNFEsoyQRJnbFcGGvqMjX21y5leCe
24PEp5bhsHMzrotNmKQWWME95MkRGmOe3egRtZg10jDJD141n5HFmRh29UXx63pn
sc0m8OKTN7RlEnUV7ARVcAoSi5hBo6OrcymTtDq1cJfYG0w9SPuosBWmD6bdPvkG
MxjjrBJDDOcjtCogCjjOlgI0PtzNdpWSVmKIELz3NPbhFLZjJB/R9j21pkq3o8PV
ut0vZ6z2diWlUv2Xin4ReistjOgQVEWgb+C1Ug46SW7UXkP2lBjYdzYLYW14oIjC
99Aets8crS3VUnEzmfLNT1BmhXrkmSzpeieZAklR/g2xzsJyJD+55HgpZaD32DgK
zVM8rEGaGak4b/q7mENtbYeIacvG6GgYMg+XvPriVFbTDjLHhkNLBj1Y5tqSNgYy
WFTem6/NXieKO5OGaX4QQyv3KHgr/WZkvpMr6tMdbBrJTtj/4WvX7wwYP5tAg2Vh
PgGEpKteTOr5IdVD+w2Vk5Mws3LiBvKvEBHl617wu6BiNQaKBPZcewU5fzoHCT81
pL+DShX2bhqmXYVtvMLugrLtW1+IaUf1Sh1Mgn83+X0P0tN7fs97cQOBy+J4PKUA
8Lkc2FRfNjfkcdxg/yp8BgUpYHZa/BjwM68DN9GqwB202tq55lUe/ZJHU9XeG9GJ
GF/yHJFwYOgFNcJ59X164iIwmP6ujKO+TCIB0f/PF3RxRDZwjSPYGwApQfLv+vKF
3KY8sUonWHM0psPCRmp6Nij2A/nYJwcD4H4T0ku+muue3h5Oowi9/tY+Y5207jG3
GVfBP2JCV9A/K06vL7dL2YOvOYOrOq/lmiEp/BrESCcuhjWi8EkqMuIyLUsBwh6b
rHFSNYoANyP3f7C81Z5XayPN3CYWGdo731DBvx5i960tP4KzUbb9eXmVCGxsBTxY
EXld+SorgeF9ebgUZxrxXYO1FameA+ThYGnlLjwAvGeTq+Ody5KzhlCn8YezKcj/
KZk2C/EHFn0up/lCk4oghwvZcNHaDuh0ou0ISIbmefch/ZFdBBXlyjl8k2sLP6TV
3fuvRcEdXpRYYtQkRT8rw2pCNcDSuM8ApIBCaNh1iA+oOcaWKsig0w93KLgPuxQP
QEtV7NRtZHc3z4RDnv8YdVwmmgYXuNQI8Ah4glxD/T2yDuuJrf0fp1GoeJqD2XN0
vZbgiG4Ql4JqO1vqSl/bbdiqkEYEaWbCn8thwFcZuNMzwNyTlBlC3Ck6dTK8QvOr
yQzCsW2nlRfDU0xc7RYd+6eu30WugUw2IAgBFNvC4ZQ7/CqKY16gBhZXVtUpTSux
otpVZD6FyuUaLorAksxQOIEJop3JtVBxKZs3UOigAb2yRg/GQ7u7R1oR72mSpZR+
rOwbqFsLVAWvzk4FrRoqjEvGkiqP4rYaXVW1z+49pMngpcgkGXbZI4hLeNpzZ8SP
6m2dTkGkz4gwiXM/MRSh5ed3/Bhwhe6/2NRDVIg0BfBsOfp4+XMi0yxcFr32N033
iv0JukvOsOSL51u6QZZodgvb1iJ0CDHx74mfWPNl6fvi+rgRVRiSufP94pcJdEYL
jLUjVVYdLydSdQsUT/lp4eHMOX6bYhXe0Pbw6/EIQ2dIb8mwl2jTLpbbDYEC9Z3F
h5fXYT7aiWhqWtLykNjxpPVL1ZMEDRQIv0NtchFalHr/9A2XnSpD7dt3HK7iPtOt
LyeQv/OHvuQ7encLpeTnm9Vss6h14w/+Wl3tboLwXxY1Oyc6+rHP8xGuEphfE3FZ
kMp7nSXRnB5FIjxCy8QCZhGrUHqK0896Y1i7+ObdcOrDsf6Clbg9ACw+u9c338g/
cgFFaZV+UzMM1550xJzrCBEV45Nh7/pU2LX62xQuiYnWdFBHqnFV2IbcJw/VhOHk
av8p0XmIn76Qh3k/CHuSFrd1NuoiBJ60Dy7ZTFP3lmEfPtEMJeR/D20Fm9dLc1/q
oM2QyCVuNxM+24fxpuKdjkQTqvjov2Ofis9q50dDaKwX+9dKwecBMP0ZMAHlWYyd
xSbp9OMGI8VFBSVDUJf7dvfe9GehthLsXQMORY+E6YoMPRflb34QAMp8KkEq8JCm
JIGyesv8+Ix4Myai/E3adyISFPW9yq7Q3SiF2pFWsq2W1TUhLNt7P9GBESB9dEO4
JqLhmlcDiPyESHaZubZbY5jbHlIiWWKTCGa9Y83nB/Eam0YjBpC0HL/PPRh+Bvqu
LIf3gIgqhHlEw+B2LJaWevM3Bz1YDLRnxgYw6y4OoVxo1ZaK6fB0mx7YQdRz4nB6
29VyoPF0gDxbO/Yc+/13w4K11Gr04pfXzCqu9V+87TIgdwll6UINGyXVEJpOLEvf
w6V+TGG00TTjxEIc6vq4KuwL1LDgY2790dBMq4LVSlF0KJTj2ALmdpZA7dX9Tw1l
/ASMHKS8icdMiBlLVszodIf9GPobBK2WfxuxaoC81pd4/6lW1UVrWre2Z71G3WBs
7am9Q1DRnR48mQr+DHtWpQ2JU4bAWmjnQCsh4Taw2icEpIUhCvX4kjaCRiZiA0Xj
Y2Hl8ujLS94o7fIFcNYDz0fq9bvSxxALmAV7prGqGAdW3KYu2PjlB1FC+jRCuxU0
W7wcyK2iuFPKMRDd67Qoosk2qwaRFUCixj8IBWv0uhiD/WV0zVEzlwO+BNgDUXqi
ueijBWoehMh5cz5j7Q4KbmN1IZhNxqfc0n2SRwu4GNzCroFPdbaR5MgsAG0ssL1K
MD49Z5PYM2NcxFrqL8q+5O6WduKQPyvvoWeQ0fMDbVl7l3JLVf9wtaX1yZwgSi5C
OKxZhI5HvGq1tL35iAcHIBR1ePH+A4r3Xk4UYVFNYFrNMCTmRFQVNWUVwQD/u6+q
7CNixMthKW8IAktPSRL6XjP72XZUCoBWoMLzywrCQe1DjrVbcUrCZXuwmYhMyh0H
KAWWm48zAwtpWvkrnDJ2hC2y0oylbWYdRUumdCB5dn7YSguKc+Jr00rcyECfEMIZ
Uf5eswjDuasd2Xm4aS/GOeEMjv1tns9nOPjazxPpzKxVI/6Y9qdRCb70jdSqRjqM
tGqO/W9al3l0Yonvbx/bNfx3/KTVITb7Q+MGpNb/YV1RPD35K3ZEfjp0dZ/2O988
KJ07BFZjL/sWP3apVepuST8pA04QOK7lHJbc6G0w3+qKpa+CYMnrHsZUKaQffIgf
ylHdKbb7djByrWF29EPh6yiaoZ88O7quDOeo8Dp0KsB2MU3ydUE2WOfL2PWlQu1w
Fe/cYAvAQG5jsmArKK4lJJH0J9d5Sy+iW9SXcmcm6nUNyazd/aLytakUyctA0zpm
kD8U9W6ZVX8DPi93i1/N5bRkpuo68zbdrjVDpy659GnRu4NxkkrHk8gqTIWnhm7y
EWymKUYMH7r5iEgwgL8m60RnubZC7HAjKnfG57tHc8C4XBKz45bRlBGGAC4lSnoP
uS/fNt/QeU4SonsDkXdpjlq+EhjKzA8axQ2ISB5SLAATmRGN1mK0KxiDVOEkSt8H
klYoTtyqY6Om94tVn2zRNLt/POBYrNR/WRSp6EKI2Wr/+66pSWdDOOQA4o6cJrR2
PodRU4Rro6FrRZ+b3Q+95NHiqaFmNGOwt698ZbSCWQ1e5ttt410rMBSSLgk0I4Xm
qPTuJQYc87oMBFQDvIlJQCDw/8Ggwz6cACOEHPoLxxAcKkzDeL6BfwYAkUkHLnD7
K0yQdPaM9Kna146OGEm494pa+yUh5bn8uTFfHoLM5LrRbqGMRYeoPkT84WhbT1xm
4S0wpotyWodDrpPV/ugV5XIIw3PqWNeQGmM4JHyOsyFlwIpuvfJD9maS4IVVphV0
9tFeWLlYgzWgOaV8fYqD25nB10VlniUpwZvZH16Z9URlEEc29LERd4q5GaA4auky
NqZfManBtFIt8KsSir3feNqeYF/QOAXyA2ZOCNYzmXnb2lDff/Gk5a+K8oDHNaZt
FkjTyj3LyUqUd1XyHee0r9jaG4E+DHBgYF1L5/zNzgtozFDRtRoa/tDHqJ0NHf8r
mBW8DUrLUEa52GfCMpp0IliNYALCKKerM+eKw/15Bu1i8QH+uoSQQRN6YwY/0fkq
ztXDuS73FfOn1ZAPw8ILOp9PzudxBRUV11GC3qkd+jMfV4upwgK3ondU8UPiCtMH
zjxfCQTvXDmMJ/oHys47hwCiumWMMI8Ph8gfF3hndhWx7uynUDH7gb55zF89itf1
cctNQzfYPnecPtGzFBtmZbfrzKSISiKm0VVj2H7wNCUhKumRfv07NKjBtQg+smIH
YYHgsg+nmygZ/UzaeXYIisLfHtfhDQvBVJz7MHO7Fz5hM1ZdQaSwq3ODbFmuVJ/E
WJg/f0K4nuacyLs0TfskiXKUaLCWIlNpnFHbqociiMZP2T7ZeosAVAAgXF8H5j2t
sXylBrfmDJB9zcNYPcTKMFC7KBbbHjJrGXK0p+G7AbSpXkwk/ChZNYJVfzpVWMAm
vDmqESl4gttKIpQ7qwjtTZxgXMGnFQqU/0TEoML2IxcKiunXThdNSq3SQ5voEJlv
35z1XnTTr8zsvOa6sem79yhel264vIoxPY5d18IoqO1aTs5K85Es6RhrVo/zvakV
tIhvq6Mmyo3GBzC6fEykD4KPLU9w47pOB4OiHJcwMQiM3b8R72grAHStel5qDOcR
lw0FH3XFdZjXd4GCxOiSlzeI5heQkcpllyCFFkcHgpwYytlyEu32DAuHfZNddGlJ
5FFcvX/JQBcW/XWvKvWnD8cVth0SFAip/DjEq/+HU777Qj4r4+nNV2uSzukTwUS+
8yHQ28jV77CQamet672WaCGdpfYpXDVcVlbmj25BkDLTmDoV92HJqkfXBy0qPmtU
WHpj6rHkVsG6taaPuXFRAzuj+vUbpTBuyI+nhJaMnhgkpBESq+TCMuPgS2Fh73/9
1ov4F0gGOcvPGeV7yWsGy6wOKfV9dNW2j7AQNdqyHHKYVAFqnYzE/Uk+XV+agbNb
rtQvTEgVDL7LEf/gf5J7vzmCoeIQ0rPpd0wOJUj5jQuxjqKrdRsCIAKOsLKBrzOI
IDUEYb7ADIAJV8R5HKz/9kkkYM59xYTXtJQ6KEGbkjzQL0mKTBru+3brHZu6N3hp
mqwSKKXeJrFrV9XWIkJyU2ZE8ahXP/SvY+ZjUJRMZklj2iI+27VoXtjQR86daba+
bRKxt5z9Q7pZQ4Fp+VxF+Y5wh/ePw2khstNcmJG26gOSRPe4HDI0TEgjzc6lJlgZ
lbFSq/oGEYtvUbFFR+twT62n6XLZKQXhYR/J2++RZ434GYcnczdhnOw1ae2tIAAo
+muOjJzs0hk4g3CvFLaR3FhXlhsRwCXWZ7C7Kb96aP76lL+g1sHS8sExpJPNhNae
OVwrgClDhu7itOS1EcIUHcvQKTjmn5/NblVgF6zZ7XBQQj5ZsLCOSFsTjsus5+Lb
viBx5F8P3pe7M/17/pccd3yLgvsOONZ9jujqCaA1EqySgi0wW1TICf4dMh9Mq+J3
Fq2RrdYhXQUETI0VlWf/UmLXQQ+xzoZHIWaKOLGPZxkP1yY7+Yd6yT2qIj16riMn
G9qp1LvnB4SWAhqP9EIQc3IVtReqfkcm73tuD17vfCL72duKNoEH9vSk+bw2Fdrr
OvR81vNRxtppUei71iH1uIkwKqSUNwVN1DGlfbWzW5TCp6/bS0/WA6SnoSJUvxDV
6tQlOh32kdK32DaoLJNy5M/iSucuNkhXqHKRcSdbz4+YLA6EBZ6kbxKo8+ggqUW0
iEDt9q0D29U1dyjVkwZaOygKWw6FBTaXeP0OpBUt9UYDlG9K1WRQifQKc6uGkrAx
5MMNDTJuYBB84cmSO4AM2AIo7ctBq3M8Yne6gpOE7OV2h9w8bTFv7hyOGtcGMMIg
axBTPRl86A+zDeoL5uKTlf+1kYKx2Y9U3b3U9gt2rlhSI1PDMgrNeMXRiNu1sXoe
vKdPuw/VPieaQKqQJtQ6eVJmTF2QyL7YUoMVq+dEY5ocCuuDenP5os04AqQOSxhL
wNr/VTetGRz05EM2Bk+Oxbxr3K/Bsq3Gb1nXhkfk81jphTPh6U8ue7HjMRum5sVc
EVJLb1tY0DYzMRahykTmypQ1zw8NHfRp3akN8vr7cs+R/pWMoNLxgfJCF3Ritiku
91HT0GXr1GZt8g0TzilMcXtc010oqSn6LZIaALCN+R0jlGpeRS5he/O5ktwKHWuk
g9tiQ6d3CkkvIM8BgwzZSqAhci/n1OPK7l37/EK12XgASmz6sBsbzA29/526xxYe
uzDFe1wbaglyPEApKp+f1pzEKj7+WVyBkXtKzSgNZBvY7/5Tn/FdN8DG/1820lwq
H/FU4jwcAu2Yn5+Y0lOnkLmG4Z/x4Jlp6hRVKKfGrcO33V0qDh5wf8aMt3mxHUF9
h+/PUX8Pd/MisF5mH9KKhHXnCxegS0wAXPjILpGPCirSN6t1Zcc6WF6GCFetJ2xM
hSq+6M3o4/VIV5kAP2saPjnmI+61Yww0HmeV3lSXScQEUfQdE4QmyaMI2XWJbBop
CLxWVDjSDmWoy3ljbc5bwIKCjGAuDqhXki8eEITBWytjH9ma0Wzu21t7ZrUSJu0E
gc/7eXwN1gWYHWz8LJvaPfdb/hf+fqoSw3AeIEo6yJVSXUUcFvRo5tfwoJnetAH8
gOpzxJ6FNbTeYlezuxvD78TXEM1oguwxmJ7+mFDtGQjXS6+gLpn3nZ096od8NUtX
vMb/uBe0PP2MQds5PMFP3hErHFvYZIHfk4+2OIPuxtLAOtSBB3KFp6zPdMRZxBOo
tkNpBR+RVjmvxPn3ZDFrpbbPhhJWgiO4wfA+kPjm6O1smPS/rN004RHQdYTWEfYR
pkqtVodHd/eQpzYKlD1kW/uxix/6HhNHLuQaUpHDNp2cd3C1YfrgMyWRJoDVks3f
5Q0tNGobQuBfuCdmsK254WeIXPeVialKGl52tRmIXi1gMbjGyVKNRWE4zRCg0292
1nmaAOOfsSihXYKfHZLSjz3I/7Y9fA3VOb8JF1DenIEOYHcK5hjy3n3YtW/ruiXX
Aj78w8ZUzfT7/U2/V57YB9PnCw90k+EL+zh6BmcJWvGvNaj7Lwgg6Pj+mbdK1SGU
WKDRW2cgLbkmmlTq9yzwAw5Z7+6SywLCc5VLdUuFiY4upOMzr5P6giuqeo1Vky8W
ZtFoTWmMPdvdDgwunEvvV3ATrXOvpBoYfb2MY7oh3vQnRG218L7JcQlyTAUnabXw
3JxCStUOhZkEcX722yt04aEB/R+ICxkUjLK6wXbAyXY/AjexpOw9oa+pxZteWAlx
iAW8S/L36NlLpuUnq5IEa8yWJ67f7YmL93ZErVjkdJFLBa+ErFEH5DsPg8d/BC5F
/pY3aLe69UnCnKQiKCJhoyrL95z66jctWPunbr32RZ4zoLd9JhtX2yZhmol4ANev
xTjPYhKgj2/D57twnapOYQhKh9KYGlRPPar92Lv+73AVQVCYNVc08PVELCaqub67
n9+M1wZAz8N2kIeqdLCkgJYj10TTq9F7zeQy7Kvdavb/vQop3NMxcvcv8JbrbfHI
mRSS+Y1OJAINI/AMSWV4gcN0HSlkgGT/JhuQX9ub7u1rr5LKcBKb+yEb6Mjb4CBa
8n5ZELlBdVu/Zcs7ExSalenqq2N4I5m/VKY7lNiI6iryU2Bzxn9bLP/Ngy9Q4z5x
vj39yHk/qCqBbCmc3NVTNThAjP1BDc3btbhNUnqQSfGLPF0kA1imrC+yYREGRB86
go2mtLP6EvHc7JdGADQOp5zHHf3rS0YFjSnaieQeDtjcUF/Nsm4gmRLm8uIaWPxm
9usKgBAbxI7wYzd0N5QmZvOKpovxJn7zlIgDEopPlIQj6OyNRNY4/v9dnJE0zjKB
hecv9SBWHbDUB048eA2UBvCFY6M7t/WGUvuDlQwmAknsDrXf64zHXFrbKwzuv13b
kteseustLRy5bL2UQv5Urz6QOVhamHwXPk+maBPaMUT5hOGTqbamV7a66LGlXvf5
UBCLFVLCuFqSTlpXlf56ZzknQTWZDLnbV8W7SLUCbFnxoldnnfXGZ6mFxgROAZZx
6A4B6aSTyqCs0DrJRWP5CsLKv/sGqtNlwnbzBbxrlPB500trsAEzJp/QM3Fw8H9n
o/qgOUrFA0ppEOctIY4sNpY5Wnr+I8tOvcZevbPY0uVewkxXZ7+XXaKtGO6rzsFW
7VFY8EdLeYjcSSc/RUvBXDOTpHsREl+yTG3VVxEyAopI/z6gACfnq7ffqpZnP4Qv
dxA06rPHKIU5Vd91C7poxpNRjrp3oNQz8Z2rEzUr1BVYpdskBjnZqtcd9ZunFHNP
EDCLf33xKs1EWo0SCRkXwLayFLlqZU51iUN0BsHmyuaXInBQrJx6jH9vVM1Jprl9
EjxrLZ0yfsjEeE4OUGyIXwX/FqVzNMPVNsxwOQFmkev62Otn9NnoXI0tAntHvNah
hMmVMUHag58pcd4gKS6GEPGUDAXdaHKFS9ZQoekace+ZMHFhm7wobB3OrQZxqsdN
rT9zc5Ee2Tuecnd+9griHikT6yo/PCVEFbztDnkIOWZ6VMFVoK4I0Rn3JJJNvt+t
jfGKd/c+iPKY8dZNKCOnF+nArJPDAinfzpOwVB9K+THeyyUWL5aYD7OUrsS4kg1b
SvODeznXc/BjRg1NyhRz7QdNKnqXvEkmhZ6VqFiSbgbi4FWY0pLD9W3tjHpUonnw
6KMsX1Ocw8BYuU+RvnQ8uLAduDBgMorUGIj+NBwF63bHh6M2VjyD3daxDtk8Tn5M
hqIsfYe1LaJyy6MWX73yYq9apf01Qin9yLkkX1yH8orhuwN5Mj3KiNvX5fyX5MId
w9m8Eb3jhzNqigkPsGs7H9rnrb2b34e32mCAkNPeV7kucG35i16TWJs1oxduC7x8
yVLGO4NF/OAAJtNvlmr2imDaXSRzp/IJxogGwkKQZtvTx14ETHHZTA1LA2dAd5Ak
zVlohHwRnrjl6MYoGZFMWiNg19PygAJ4Db0wJQ6UOoIXk6M7sbzpovwFvfxkBKGj
T3TuZQComPMAcGxzsteTe6t5Uk/RaFaPho5t5CWmGw7zfHcc5jYMjbAxbZ952OWh
7XVaGEdL3sukBYW4e1XY80q3owbq6L5B0z7rfXnRE2A7ZS1sXOawJtZuvirNjOuy
L5hxRUBeH3Idh3CMla8w3cm65BsY42r17Do9sWR/7JVbrN4rkPExpn1wHauCpzZr
IRM3NQnwjT1lEihk+1MKg6nudYvwyCXheZM8NJHofGvuqimPSegxH8UNdnHOMEZb
Vd+NAvBbA380gyaAr0qBojVqYM+WWOdej4YWt79EtSibPHm2+4j10/Eexo5u6BCy
pOYnl21sw3R/X1HsSNmNXaJ+Fy4jmBDXxc1ZFl+fIdnQipI+UIPdIfzfR+7cLewA
Da5jhH1iMtqtZR1OfRVpeePVOC1Zy9mLZBaC9MJTQYK8a3WLh8p8JsHUq+9+OAlC
ah7RzLObGTevY5Q0D1KvZAPPIcMXeauCylUX2NqFI/RG2XZs0QhZAY1i1EUo0Dyc
ItCUZy5vE0sM/pSuK3gSRKXmMLWYU+anJsO0dtf+XrGokrBUhSoK6LR0EX3/Lt81
Sr5aclmO0mPUnr1G9+u7BBWHJhhr0di+lY6AadrFrI/PA4eraj+KbeSYicPeKWfp
jhU1O84FpJMesWdxtPjLpjfz8nU6X/vUfR/Jzq8aWlJgkMy1dpw2pFK7NC5l7d3h
HisUSLpIwdGlbTqpcGn+7a5lwm//zjg1say3pV0YgEgXaTXdSsTQlPVK7U5oe1mf
YrOtsNaFuMlM2nsVGRn3YXmm6xBCAeAepc7RW2vtnZwWFFX+z+5+gVTlQiaNzoZW
Qzz8m5EdrpVTl57WWXJAEwvXgFE3wu4CI6xiXKfXUTPGNsjBy4yUkV2inP3GxXar
ZjWxbalg+zSZ/JsPLxL6TyImtC8H/lmuV0G+eNSrIef/UYPWODV7LPGhefeEw/sM
csuPvluQ0t4aV7+NEZMNhL7pMzLS+HT4kuVJmfWrn/PY3YI+eM2qYYDBbRUSnBhe
jncT15sv+fWmkB4RvLZjUcNWdFLZRp4eddUnqHOSdaCvxm+aAK1Fads6h7TU1J9L
NojeURefUPazGo59wPh5/JUX/YmQfp6Fa0bXI0fXbkjGkf2TTmuhJt9kWUaLQIRv
eyj2p3Yxojt84govIpKyJl3UDdIu1U1gSDo5zTXqikwfrqXj8t9zUuqXHLGxcBcf
CSETfnQn1uEpUaTW7aot/pauau2qyhctH+dNKc8cGjWruRvB9VMU6ua+WT7p7itf
8uGvHMH4y6/WMTWObwI1ND1syybN15osLR/xJQWhiPLT3VBp8bATYdCvevZdvMKw
EmF3RRZgpdZW5rcILc3Qb/icB5pFdKc+yxVCqy2o6wS7uoXhHmDYHF1C0Km8x94R
duHuTGA1Re5Zkh3PzUAyC4I2DtGQR5V+57Pb1E9PfNnSzsfGObR686+v6f+eXEir
Sd+hqtOq6GLwJFkdTlxjRSE0UnLdsJPogZiukLs5+1XL22w4yQuCizOq+TQJsGQn
qJeLs4VFwD7LtOTWZxsx8QNtaQ6e2pFnJp+wQENTOjqV/FyygTneAGiEZgG/2wMs
Y8e7zslfKdAw9difbi5bOZuuletNkYhEFfIFUBlzRDoJIqUQgmbAF5GMJu9r6s6j
gWaPYM90EH26arwxiOyosRKdvag4FaJvIryU1Q3saBTBY8hEJgg5uzWpfwYTnhun
HCxuTzBl6xa4ufqNHNfuC7+WsWLC7Jnwowyizi2GDBEzA85Vr3wCP8GeCpxiAIUr
F5Skg2Gy7Ea+cUqIpHZ94LX/AoM90UK3AvTlANJmxTin8Jsx6Myio8ryfwEdEjhM
FsgkLh53/Ix4S2mCqAU0FmeBv4Cf0wK2QmVo6WWJQ/FQE0AXae5xY+RuSmalbyW1
gM+IP9N/+sJHq3ZcGFTOVKq1OfeoCzGO6rA1tV6NrOVkOBfRca3r9rPnib21XTEx
o6EFk3SWyxgPAKQ+fbT2blt0lk2zFXjzant2Bz9FQsgPheGgSq6huX0O92wbsIBH
W5jlfr0zGr0ws5m23vEs5L1GmiDGkzZHFMPgCU7SJE4IxyLKF1qsISwy8gSYLH+e
AxhTXMhR1O+KXbljjnTa6p3jmgYdub+nhUXNlZ942hZk4QybN932JdPTxOOjl1op
4cWV/IsZW5m5GS2MuKtLy80FRcgmveXHBRUbv7H6DrcuPD+iQZqtVsZ/i1qlRJ+k
IBHS9NNhGKNr8N6kkdGsd41RVVykEfo7r8ry6YaGN4KOA06Jvfc0CV/M6C9DWkO8
U2mg76qdW849jZQkqeT5jFqYyu2J61YGQa21ESXHJRJLOVVLyOGZvVUw5LJK3h8c
a8iKX6Jq68X4zq4Jp9ia1dKS6ywbjZDGsFmpLn40yaysdFNkIA49iXE7NuCJcXyq
nWLIYqa0m3vk1MRDekM0Cw3YKKMFCGQUnqAYt9zQGDCXk3THO8xGbcup/aQQdJd5
HaTHrHUvnwX1L2eVrziPj/qikqTlHjoUbRN5H3wgml45LyQX+muEF0TWl1oz6RAq
KS7h5cG7jy8gRXWVJmdWz9qq/t1RjxZqu8KqjpUhvN3ufy0XRUiY4lHrfjCvw/rS
gfNyL4aLp3VU4aw0IRzA/7r+ODUXpvkdx3CUGVBx3yYfy/BFsUYDrT3BR4uU9qRx
sSIIED7006xXYoh3pw02Mub3150CZ8VUJm3BMOt+Sud+/bsm6x1Drp56Y4nNi6Jg
eeAfkiDwNVhtyTjyjyDxg6vnvnuKqUCT5pQFBKKukZDhw7+JpFCBV6X4NSYqXgrk
UtV98o/smpghmXdnxf/IJLjdW/2BugM3ZQ7Lk9OGuuG8iQyFb2UoqX0JWsmAkweR
2PXdQby8vIYYaOs6tnsQ1QlA0NtuhKZifZmVIg1nzuBVBwADL65g29YCYRVYxX+t
3BWpa8GcBz5scNdKuUIAj3DlQaavVQqZWo4jmNvaaMwrlfF+LXj8SliQpMtd5Bg8
db76MiUUDPaJIPbpMEo6A+eKT7zRh2AdYATvX082b96yu3UQcB0KplMDtjnb/OSE
jr0NOZFDXdu564aWUDmvMem3CDEUWnr9ccpvTRwspPls5w1/x6GhB9AsWG+AaveP
Qvz8bU6aPkPb4Ss/UPJncN9EjgZsE+EJauxBFKNSgJdYgltiSX/eekJorjRCLAF4
MQBHJY6HuitlzGfA/CZTwmM1uwCWXxZhlNdJHyFuKuOvppbAvmsYCVJ7Pk2uwyvZ
aNcMAOBX+AQ/AE+WcNDysY/6X2b4KXxwOCjoK17hMDMooXPD16zcYl5vUyeFWx7l
MY54cVFIca/kcEZkxJHChtrbz5DtO/KSLwULA8V2ssYe4mvVV8AlNsU6OzQy6xs8
AEkdBdWFGL74mj5YT0ZnEbSBtA3SvnJ9+7lYc5Utk4QQaW7pCPvZl3iEZPftT/lx
HIVBSRAVt1TTUZlXPidnxWklPAm86LA+DK8UnyMFBjm4FM8qxodWYcd18R4MnMQ/
l9FXxoriNLfiJWl7NjKGSd33g+1hLl7OF0mAt4Vf2FRMJsuD+RVCFU5P6WWoeJla
Ax4gj4Q7RdPM2G9zbWOfRlPCZcDKqzIxV02OnkgtduFXa2Y/T1sefwFjHT78AxuD
rFU32fpd/1HgxkaV1lVnIE01kV2Vh2J2rpXf4Xy5BVxFA2HOjpGHZcUcKERrnyFf
zcL7Ieej1l0YceYcBNtQyuyfyslRaXTIBt0SADWhnUNewFRhu2yEG2xiQ8rPrTR2
ZST1oqZ9ouOnR0spkntT7OMkDR29zbmS9+bsi8JVpL025rh4lKA/20R0g07HmXPc
6Zbw6+73pJbE2vkyDFvLiCIUp4Zue9CI+LR80dyv0dOVsRpk993mfgiIBp5pTLMe
643VEk4qYvsYGIA6cD0/bNqmxvLIYDhGIvsR/NSUvnQsW5oz/TAWux2m3GpPApY8
o7QdnR0pflmjukY1UmMbELXCHfvOGoJ2Qv2GHq/5rP5dFB1UfoHszkSKWFocOtme
B/KqqYTNIiAp5HuYT+oBKo8PoiQA2Pb6VDhaa5VBCghSucv47J0ZZ+Bxv5Eih0ww
x91Trl3IPPepdsLtZrHYb2cfsSXEnrSRyVeDWGnMYwjZU7Vy3FRlwZycmGVxaWjo
c63atdIdfEQjJ2F22RYkbkyeReO3LmqolklTNSY1B5fPzEV5wh3RX2BKU4a14aHa
CJhSUBnoOLoJVO78lx57dC0R2G5tQCujbiTR0xCohdzQzGw9M7j3kYWlkeMGTeTh
sQUHyieMnnOm6aIbHvCLb6gtcbQMLQER37Ypi0YPGqBOaHI5cnd4cJQTQmODzFzI
BERELXqSrRPLANIORYekK3i6SW+K66sw2Ef/z6Z9lCDkJIE8R4/uhC9T+mLvufxI
YqKStKTKPGlUPqdng/32QByPAc9FYCKd0od6u5OGwIO1XMU9htrDGbGJNAE/H0tr
swEXhoOuVRmSpSvRQzrIW8OwMagSN1UwYWcAwAB5+82AoQ/Z6XSrcotRyB/IvCaV
A93Yv3gjpSx4uq0ggrVjX7DeCtgpjTdBHTaG2ippaZxSHexT1fGHeUzlXZ8WnD7s
C6koARrPaQS1X+eEPOH0oCds0l95pqieOJ9jzmW+ToHEbqUs+uO+DQMRKckZZfaD
djwgfjsEPwnU/mYa2U5362jP0DSqwszQauStsblEg2ngoOgvHqWbDsGBRVOX0A/H
+r9vcqE0WeqsZ4U1zyRRNvOEH3F0JM7xhqbD9S/L9Q1rN2CRiWnNnTfzldBmSBos
qSrN9Z8xQaAPGSbXS5cn7RsclZ+ZfE9eyfPIqxYZqimRjaGf0vHKuK2z3NZs87EE
RdyyxUcfNxuTPjAMgH7CeZVYovWXE81wR6zkwvT1PSbjdS9vQkO8jABBYXFUwb4R
crd1oHeccc13oZ9l96/vgnhgrF2bHyq+plOhqdBoV0WTPOTTyOj5g1mUdnnmYrz0
DIZQRhEtMafO2GMWPw7NRYD1MRRfckZ1vvD8eG6JpMAdNM8luISyJvTCMB9FFmy4
+3q6yPW6ciW8mOfcdiI1pNNgT6xIRt/88Rsy/oJ0tUt3TG4HX6CHhTK7GuPFdDfp
nIrS7Mx5ImRh+CYY3x/PMtKFv+GHlGVK7rZMbb/uDX35bf7KUNXfLi6ZZPjAntHr
D6IH2enl+FV+RqDR5XV28U3onMlFDlP7AMwU8XhciQJ6DQCsbrGNUbUbMD4fD72f
08K668r9GHX1q9EpcLaVhpuBF3Tm/blxY1ubSk4+WmVQrr4gjRSiT7LZQJs21ttT
AFgGVGcXUT2psIrRsBIlFWvaxXVIbxIH5Zp14qftY0QnJY6/6lB1MlPYHsnMbaP5
iTwX+6A0Q66/O9BIronbEessibCkM1Q2T4aoSp/3NHWzagNXOY+sOHHoh95JPzDq
/1K53iHvEuzr6QG8aiToBZHJIZopHU/O27zMaygD+Ef0xyMgDogMbU15r9yQvtld
XAO0SLHfcny7aJka2aFsbb6wKD7AZP9LfpeXaZFD4uGFpIWky7L1JmN4c2FzKzk2
xEaNIJ8NE5TgqJ08s0tAdtcDeuD6P1WlHqVA4OXsw7R68JlYRkAsDCmncTdhYPme
QCeZjeAXbDpg6Dex0Oc2Yk0j8gKnWYmQT6QEoXLv+/ccPFPNc5m/7bqrlkwuz4qI
9ykGsV2IWpYnCK1kW8/q+VQQpdAkp5AIWhKoAzYBnIpS/7Gh0/KVyPgA/47OHSQO
0oq1izRpd5Oc9JJqqEUgStEL1c06MoQnhqX4kg5Rp90cZwa0/14NE/tbxXNRJRdT
UxsEyz21SnHAoaKNkeo0/vIh98Rz7039GW6eIpSyv1ewz4dFZ1OdiyCbrzcUGyPU
Tmd2L9JZaHyXOMpwzswIkcfo/KLfv0DPSsU8tIyX1V+J1ecfhoPyKrnGy18sbK9g
TNhwIMw1BpZophQJpufSZeca/W4qrUlKuuM+t2dulbp/91mbSWGAdBYKSak20LYK
aqtwMvpxQp98o5RR6TsTck/VvCnBn/yxWtKgxLha3TUKxVlqp6uqf4xsH+G1cH9M
qOihI5Tfx3jOXecyZtaz+8Z6loE2F6dUNUYTXZBOH/iNu4ZZKPc1ZUn9ilV30Em/
6w2JUd3967vCBFZgFBq/2xy/+CAlGcK/7E1m4Ohik7C36+YNwR1ChO4l3Qf6y0NC
22vUs1HpAZJGBn0ku04+DAbB2vCokAiRG/6JQCQCPLTOYVld/0JLXuIbhkvyKc/+
55fy2fPEp17BB8LouOHzoyQh/KA+f1o57MkZt9hA6F7xU2mGqsVeSk01vT+pd0/n
W+DE9JBThb34qOHwzo5OqxWIE1BgWEEIDpV2q2vgauoKmwBmE3ceHkfW7dlCj9o2
MlyoANZDxyas1uhMeGAUeikEgvdlEWHjeHigSrfaFJtVG0DNNsDW9JxcY8ZZx7Jn
gWhPronO0I7FG2lP2x5VHgDFoNdRwlnm69V78AZ+SeFPm+JPiNDp5nzuewA7woPv
SYDqS3GLwPKJkQCT0x2h1GL6Ho/MsYFshmX4G5hnseDM9KpRDaMU24q0TPTPpgzA
LQc7yWZwsriRDPAzcsoTG4ODKW0E+W3lNLhB2ueiezaGQRbJZVBMGueFvDy/H+ln
nrsczp4aFcz7KHwnXViGx2sgSSJv6evLxzFz0+2bzZHxwAV3IlHDuita+scYVN19
JHLSkybiscN2uZ7I7N/j3/9XsR0tAF/g7pdMpZwOrnYe6f1zQlDNUP5QOUFvXoIb
NVIAM3VuPBRrF6nSaWM7cnvd9xA/wIPljlJhkbHIngxTX2AzuA3j2MBPlRyLnWWX
m1zJHMr1ivkaCPdMFtlGPkvq56b1qxPF6fQsqfUFmIoUbMQImJ3DEyzhGJl48DWB
Hwh5K39DoHjBw8r9lknETzB6emILrS9WXeUR+oxOA6tg0xVUdynooD3seX7OkRa4
u22ksKGpGfGRc5MlnOulevZkiZD1tbl0dXGVQSbLB+Mlzv9vt4YmPtU6V4TMdxVn
IgWnyvRuXD0jAqfPzeKkUr+JahjqcglOFiCHiKJia26SKo12tZG0DPNUpD+ACOd/
p/RxJkKvN9gF4eYJMn9dVbs9hEPcIn2Rj4712paqchdXLBKvi1Smct60VtKeGS6j
rIw2wFDevDFc3y4SbYxrevaakGSNFlBDaOvINiNwYVVKcm2nRYY5XCmwarXSHE+B
9mD567S4lnO1pYxXTCFrQ1eYgqDdPR+WU+OkfcNwF7gil0Zfi3kLqx/Asmo+nJzS
Q/MN4Kwt59R1qNtYuCCBoATz7kWlKe4DFexFGlPiRUTo7sMxAVTsG208tfrY2ag7
WvHiD4a/Epf5SO5A+4RQlsH47gcoJ2VbbnnaKl+SbwHFMU2vKqWnmfBatZOFSYl5
I9RW2JCxpIN2ohda5vtDy+1uEQ7d1eALsR76yOzdcBoODZ0ClxU4kBc1LjGHi6Eb
XAfQyCxa9YwrVjMrP62OtRuWB6ISCZOV9hKk0w3k3PZPhn2NNHgzylECFiGUTOg1
DP/zBMCU7Au7XQEpwqFY+RUMcLE11KaE5aCVeOhElRkpx3ZyoqJeL4/+XPi1e7J5
Zregd3mGzCH8BKtGtCI+YKHf36PVqGoQuXHP9oZI2ZeJn5I+58K8QBJXo7lx1Y0v
lttiCvi+slkhpu3XM+dwzJbiXVBM8DU8Zs2zrcaBVXnIsboxigc9ZcWFE3uyJsY3
4+jwKqUoAHFCmbegb2COKROI9ASwHiS3xS/o8QmWXi6cL60PkyqdUmBgAI2MCvu8
6uFOrgBJwqx3nzmKLIfhdNARiKucHN8HLtrFMSrGg2aOM/UKrWdKObVR+V7SaLOa
6tGrgh4/bnTdTU9WtzJp6NKT1KUaXO9r6eCPicwog3r0wqu7LQfdRuviP+SaCFW/
C8RRerjgCjwE8DIG1AVfcDz89SZOibFRgbI80XFnA4bUdghZlWsn38OkgrUIOcbb
LcOIuvVmB0ZXaSMZAu1hRaBK9948TesKn/W7vxXQdz7ZUqmkqvEZwah6tNpE23Cm
VgCCOB1Tn84e06Iw046rolAQ0E5TFx0VmlhrgbZrCcOnEq35EX9xhOxGc2nNYY3q
zNcipqY+rDvgaRx/hADR4YUCQG8h90h4VIUAHpCelMpySpW6987A3tNcH2/8gV4b
uLDAVJXaNwWJ7w4DmhSXNswJxJ35HC7LxBh6CPMDeGWu4sYEjpK8RZnJKhP57/KU
wRDPxLMhDYdr/NYsBRQ6vUPk7UMIbVXb+1KejGIoOINGtGdVaDFdBXt5grpWOt8/
cZ1xERXdfduFTZe4v9vjD9Z5Not/i6x5xmLTx3HcnVYfck9O7ohFIrKgHloj8z6x
xc4ot9k4o7CcDB1JBtD9b0QPgDBl93Fs3QoHgVN8gO4Ux01sFmUka81I3epbbCDt
aZGBQnp34iIK1qLACDFAEOewrcib+fkGuhSd+1BpJWjzROzOOQvIXtbkQaCJlg8l
jTf9uZeZoE/E3x4jNEqEBm/1rgYZzalfiROAH1wQyFk0x7haE7WbNQRD7QSRxOfl
S6PFxvnfGX8q35m6j4HWWooJqiwqrCgJYJESSR4ufSk/vJpktBDZ89LEDdROjLfp
wuctMf25oafaALKQOcjIy7bG4+yQq2ebkWkmHVN4VC0MJKHX1Qj+n8XsLFGNRJDe
pW3sxvktA4o0XJQL5CBHPwO5O8PlefJOOP57AZeEM35ow4cCwMMVVHYzgYROrBtJ
d6uJV3yaa4IQJkYSF9+vfrmTp5Fatmr4mjoZyBJrEJfvuSGfguZf1H0wFKcGrmyG
y3pa9eiINaHwqvk6LvMMdi4cv3emRvAkow5igdlXvvxhD66wjd0yO0nyO+Fa9FUY
zQoT+mCZL4cb18dVW0rX8ZtU8wCCu51ZgVGd5+E/bFhRMoiMTgh2tmb0+Iko1SAS
x8q69kzTVrYwjidn+8LTrH1CkSU/l/ot3ad/IBQcciX8ro/mCY6RKBNvw+F/j8DN
qdlVLyMI3rdEP6p2CZ3jCykCNC7zZ05SW1B9i0D6dEE2mHOdC/YLesIbE7dAxbPu
xUVrdcaVsOYpO+w7sRXJ307d+8beV/d3E/JJWtpIap4rjorW2riSwZ1aNk7KkHMT
vB36JCaq6A94OfhTjq/EcC2YTJ+Ath0MWt7AHl6Dwz8XU3AESUT1urq+4nx8QERC
BYbzKiKbNsrIbT5gsWAfqt6NhMHemoleVNlB9jU32NtJuO1m00uopjLy8oxaNF/4
NKHbhClUIZ9FcbzGJvJLYtruyuyQlfd8R6ZpjWmjdhV9y/s702kvUNd+/tQorwr3
pIf0gGit6EeDewoIRE58wCYCcS89dkvgMxEIeW8LD7bZDMoXkpGSQkGOr0ZugB5x
3zV5geDTIWc/Gr+oiy9RMT6++/5f+nKfWF3N4KyOdTrM0PaKObr1Ht03Ua4HPZO+
Fj6tbU8mFJaCYtGiHu4qUtGvpbgHf7neUzw/AhIiM12wyGstJgU3DMwojR1162Qk
AUyS+4fU65PCaQ7+Kz2taBytyuIGmw8zxcyQKIlG9dAC2wS+F9FlvIPFL/mBFkV2
CQT7HdZWkrSGINTAYhMeUSKQpunZ55bqcxn4XdM4525NOLpTamf8wuC+d9FjH5Ms
MLBUiwfKnOCcBeUNbHcY8FMjGUrxrLkPMxcQvvEyYv2P4LvVJNEIM7MlgPGQNk3j
IeddOtFiY4oNBNqzgMJBa1JsifwcqSqCBANmQ7iiaItoQQJA8zWV8E+z+EDitMZ3
x2MvWNMTuOnOH4rsfWH1dBMR55OOD7lQa0g3hwUjvNXVJxfPZHTNJh0AB/QtQgVL
63d9ncGMCAwVJrcxwbf6i10qXJeO7Vw4DBYWNsem3x0wFWNSKmaX8JoJzndLQObs
YfqennWqKJ5KuAx1VuvcwwJW+R+rhu2ZUqo3zhRuIPZpQOTvXbvXYLqXS3711lFX
YfqwCyPCe8nTsUBYARYLQAGS1S3kMdwaNa8nuJ1DDTydVNlvPSzIeBlnOyHmqctm
cFbxIJA83+d+igCVDDHkCd8cEKVLbXePbvPMtPv/oEsyJZuHGdBTL2qxb1NwAZoz
7dgv+gSnZEPq6HvZc5JCWcngyJ2sUX4vKfztbT9M5Obl/ZcFpK/7PQooEZ6e/OdY
Zw3ldtAS8+CSZKp9OrAMSRANY2+u/b9fkbwZAcHAKqxyTmDKAB4IPgHgzWBuzljT
F8yeTwSEmYlxWEvPfa6BVNDsh6iWHJqqo3cXTMAgeWw2+QHaVYfQFf0zi0SZNaSr
EkE63yYxx1C1sBuOVu/mLZczhK1u70G3rVarOzeq+morNeVsSJozDTRsFRZDvUeK
GDlH5lnKbjwsUvnfrc7GQrfggvae5oDaMFJ1nbCGiHifT0IQBs410oGAffT5ndMC
bPdsKRpv2vn/iBdBxpeutH87Boyy4h1eICw+6+ChAyS691f4X8sf1WPMUEC5EDPV
v5OFVK7xGFeluRfKxczZiYtAJ6Bkk4VQaIoLwVfw/WniesY6E4SKA256Y5xMi3jW
Kv/hRjc8loDexGofUs0ofC3tP9WFKlu87qLuDrL+QjvPJkKSYzFKtCBjRngMn8bJ
7iNm1ejN+likh5xak2Jv8Kw8zV2vHJpVRSpaqB+IzmHbPEru6iAO5pHpCeTAz/aL
Y2YGdXk+isuSwsq/NOlXki2y7Kz3LfOQrJcUVZfMymHo6ZR/QK5ks+qk6ruszCMq
Irv3vVF89l9BYobqAkMPZk6ZcGYhSB8fS6j4oTvL/SD/yEaWkGFfb08gb1ZGTKR3
Ug5JrGtvW1M5ieYe/ZzOKA4vO6GLQA+DwFnmUP5oJPiNGaAK9hPpSslHRYvI+Tw3
ZcDRu1Ya91UWY0dXE1w0/kM4cw57UHXh0T1uMtlMxbxto4OFDnGt0YJ22BhOQf7t
W/sOm+vJHPwcFjArjcKsx8NFd22wdqsytnihuBhmfiJIK8tnsCWIXJII5pz2oyCR
DfwCqB22x9SmfjFe8YxvB/+lBdyA190blNWQkfjOgc0wCy1QNhov2PR14YkLdNEC
boTXuqhaPHT/uY5auUpJT0wfIIlufJn2rSvEmh1QIIVnBq1CpBsp/VlfQwKBXEZ8
UAuZjg3uWxdtCPLRHFfsBaB9CsoYK6D+kBZ9UYakYc7dXdMwq97gTBPpITiv3Nl2
7JCl/ffLIn9dD0PvT811s/DDSn48N7iyZdJ6rclT11PSJd9l4aBlSN6KCT5hpaOU
hkhWfo196T7puuI8x8fWzKk99qc2iBLKCEejob6P2Izj+ONJXyMgUJ3t3JuUnXrn
WQHarno73L0KbJ2WobPjAwsuQ3FlBCP/bKRLcJxD6jO1Wpb+Kg7NdOPVZOzb4n0Q
pHBCz+Hlg+jCtPD+h6jbH2ndnwTGKnd4Lq/iq5NboyqRHN0FwUai2NlRHiulYpoE
xsGnGfBLxfH8eqmkHVlTi8SDzVTmuvSKZg3cZNfh7z0r3QfS11O9UR4M3fKxgNji
pPbwP9jgTaZC0p9CKcGROmaj8w4A7SJve+3qZbHO0SaGb6924xTQQX0g7RGZPvqZ
LnRy6ixXk+oNwxBEzFWStT75IBby+2/JvtdMp1GWM8bttQJQ4fGA+MIFNvaTvb0d
UMauMh7E/02EdVCexIMQvRCyHrVmAYuzMuu/Nl6DW1Mj6IDi0AJhFO4EuNemMccj
WldeeMVqUo9i4pYo1wvCyY2zB968hlCoaNG/ABBSWKTzAf/iiSMqRCYKXwV7JPk2
qEboaa/KDQy6/5o75oReNIYNEiZi4jftS88ARCDOfe3y+0fVxIKdwXKMW8CsQbPc
kYVEDu1wySZCcDufxk+HkC332EPVP1TNt1TtePFivGriAwqEmVpvDuT97g27s291
FLoM4jPzQ3gnFGpxfEnsrpPYH/R6nJbTKUgxWjRBgG+UYbd8h1gU6ufMqU3I64qZ
9xvtSpZnn9aflE+iqifM7dOHu7C5NSXWCrB9bTsJ2qw0aOWoGT68y/Hy7RLe4tku
boqkN1EmF0rJHK3aPEZOO8R6hDEgkhxQ65hCa5CtXT8T9mNB2TSQ4RbFPOwAsgYO
EBvHRkiKf1kB2jwIBAe/F5DgZQlTms3Y4uFh0AnBdkJXBDjJdPh+wlP4Qwswpp8G
bL2vrSuCWgCiqGfyxRjhk7ZnJtZAGHvRZ/37fHyni1mqzCywVyycvu3IyphR/oZa
7J6uyWWjhQvgQU8k/nEwRZ2sqFGKfzEgx0f9G/gXy0FyRb49306qofNRd37cu7BE
wyqTqReFensRnlKlKWBKgqhqaOJ9b1V7Na+cCRHkdX3sAZtiYS9QmL9Fmh2MGGtw
PCFQDLc7GwH7p1nbP1NtLyx+MslFUiJcYh8fr/XzrfPPg4sVjbTiYKgVaoVD4UOv
/u0jmjx2vE6atLdo4/FHjhLWWUv28rq5UsF4eu/vftEjV4O8/MCDPjhShXIFIdmP
TYfkkXSet08YdmoNkBdv81khZXHVuZBg6FU+wm07NjjHEVeioWYguYE19cobR09B
ntgOJOwMhi39gbqDXtg9QsigZ1CL6YPC09ZGPIIC+kEwGmjbVYubZBkTIB496WTQ
BC6nrdULNQDCWY3wpp2h9BOv91cgetCkgPKr1Lx63Mu1QxSCr8j8PXoU1NttfvhF
sHBNZrxIkrD9UsDmMVQk3Z5JtEoW13laPn6C5SKC2wje6q/cdxHl56e8jRPGDf0/
vYM03MaU3j43zfmqcbr+iD2QBJC4UfGIvpyuEGoIX04oys1mlF54GidrLYZdT9vR
nU2iTS9e0jJdeAkye5U5vADbPVvZsAMcpnReo6E9Nfvl5YfQxReLXjrjjWrIQ4F4
XNr5cR3LJ57EuHFJhWcC8h/usgEkNCYmvHdfn/WfjcPaM5qssvYvG47LpNlUeNBP
hqj6nKdvcs/eRUuPDFIGSIBXsOpSlrl/L4/XSiPj2lpNkjUQM/DUQyP9ArtoBOls
ENnUBhnwtosatqIrwc8F9eFgMi8+LLe2BcaIfdrbE6dyV/1UuMGmeWxyOlPjFP9r
EFpKCu/7nD8IYaVBeFjMkzBfChGWvIZ3pYIc6jY3CQz9wYTxA67f2bbypusDv08i
r/H7CAE3/ZYmMjVgOf6rLpZHH/mmu7eurLu7voDluELj8GewUWYn8EQj/0YZXMDI
PjpuqZiJB8DntRJSiAZTk/QwdXDBXf0On5vFdaQmjt0L4NliavioD84A2GPSeT4C
LNuCau6DvO31J9Cm/YquCov1bJClysxOguXKikygIBZdHA/ANtUK3nhXSF01TEqj
tSTlqngmeavqhWkMM95QYvJby2i4agLTqKhbcF3ZUsMKZ0mtw1KW7qClFQBzzHDb
uq6Zvz8yV72auGqf5q0l/oDHnMaxXJPFxk70IfjW/j9k08xCWpFG7KxzsoxmDzMQ
DiZ6OoBDvRq/ZQh251eVxBdheDjhZXq5sruvb9gH3bN8XZttx/Lgrbhuv6w4Kz6F
CrF38aywLmbyg+6/UGEMHJ1BWDt3RjK6d/PMJK0EeA+EW/lKP7j9G1Fe5TDAfTVh
r/ifzOBPtkboVbToQ1y/0nELRllHGGdeo+0Tja9t1ed7V6Vf6nzZmJM7wdLtt3lg
HR5eCWuyLA3oNQjppEt7WXZMKELfYXxGFapPsI4WVX1306nbuaZzjg+4rgg2cYbJ
SykiAf+SIg4c179k5Ntf2E7/H5S89lv+KzrXX+LuykhcSt9Du8HkekdDZ289XY7B
Q3K2DnKTaolaVK4yrRlnv/+Uz40LJMZkLw1YTQOSBT4CwXIglZRKIS8TtR93z2En
0xtv2bNLFcf2BkxdPaBbquaIqMgq8yVUUWXUY04gdjHGHs3fd1PLWkeXUEQx5hLW
hX6Vnk2aeltxHI6hjDEMnHQx+1hunUecMCOyUFKhMazCBBkAf8NwFByTP+p66V0y
bIPT5/5XxvcKp0gk15IGmeNhvf9b6LnHRAImYPHWiEkMWeRvBTvcKvgbxfcr/DKv
yU7J+lqVdPs7qINXu7rAh8QkAV/S70ttxiODYWZDzeJDa6uioR2qQRI4TIaucQOW
xBDH3BDABq4W0OX4PodkBWcmXRQ9tVpjlL5u5UFFVhk+8SI4WOjd+UMWsfD0xr8M
JvmcDxcacpyRMX1umljGybgTIDiZT6fSAg2eBpLmsKgKd0Aw7RisS1QpXmqufUiC
yVSBP296RdIsxxys4bBSvVfYJNVmZo+2gca5ov8uXhmTVBnwgV0ogAGNnpmn8KUV
entP+brOatmB6DJml6AjmKo1QYQBNmbQ8CShF1t0pFl+Q+fPRpf9gZ1X4/Bprbql
3Wjn7FJ3PHAkAg8mfuhdkKd/IUTx7oA36LPJrkgJ68A/3UbZnw3Gd6CqrZpdKx3r
jnW9qztvOO6fvzIrBjaJoVSNoZl2qgMOWU35MtI2Gtq+cbdb1xtk6UrVL/oCosWE
j7yhVFUUY47loGPjgOBtmoSDEEqDiwJJv6QL7feL6LojwSj4n1+qvcYLC4cSdW34
sSLG4ugqPOwHqsIAb/ECrRGl0Sos1tsmrX7ui7OrCuBLJwnOaNg6ZyixTw+DBqPZ
nHOuX4KwJ60PUpacVhK5qyA2CalxJ3VVgCZ0LuK/I5sV4pe07w6LCW38oDR6OQro
B3ZhpjJ2Y+3Bq5TOWxt3fIW9U6PCOnMe6tfnlGlrCmZLWYcab1slGOSUd2t8KjKj
Cp7sp8G4koecmGyDaNiMl5kfGLztSqUqHNpoW1oEplCGjaKel+O3sTvvYov9MEK+
oVWxXwqnzbPRBzk60tgZn9b8aZc7GQttncNgOVCsp4TkscVTg6sZ0RbJ6Dr45IMA
o7kqrSxdGv0itiVQhh+FPe3QdDNcXKQ0BFE4WL5w88UzOwxkfSbhS/5U5t3aa91D
Ck/5CE79Qmoh3RLmBlsz4ZcGUvukTtRM7zWWEBkeO1eos3mxeh1VLY8qKqz2+26l
AwZc5UwL5HcBdHId0CQgmxFRKHGYNzAeaCVl4QZEAhM8afw0pxH9nu5exzcQJWJp
UMgeVBuZSZ30SkWzYY1Os9ZSQ+vxnlBVpw3DEt4JPoL1l+W3X9jcIXJ/OqQPdNDl
ai05CuYo6ZoT0k5SIvAWVzTUtIN4L3o5+odz57dsjeXFezkkS/BQyRhKyuaP6enV
qVqN8mhpA84fVY4D675XB1BMyWW3jdfYqxNGCb3FbyX071MkmombECGzEN0g0mnz
/jqKrjF7a5w1/a3MfwZqrellCQLQypC7KzgvV5JW/AYmSEDr9waWy0DeLCUemBol
emF1UlhRPLfWrzezOA4RyomrXS6aRqilckAMV2UhUv/0AeMI+zUA6gpIKBfQXhnZ
LqsMUvz/dTksfRM0Yatdw+WoGpswfNks9oRgReqf8fCuL1YKhm/99JiqcDQGkQd/
aloHDUioZ3F5I4Aq6FJ9waPWkw042UnuEDFxq3b7ZHsfTzw+6mTfLaG5VnSe/b7B
0zUF/CbRThG8om+4V4dEgmKlVuiKbrEAgwf2dbjp00omOTD83m9BgJ4w4eEZfT9C
2ROBrLnbVM/aBXN9tUkygd+eAd2yZPKLr9Tr2l6qZAbKi54Mt9e29NJ1BSZlky/S
sC2qJlvaaM9H8u28e4bBOdHG7I+GSGd/R1CqF+d/d+Mj/Y5o4vhkBi3QoR/s1hGa
Kp52A7pnZ4YBqCUhF2OWEDPU7PEnwtuNShKM/MXX3lnQi+09gsupmI5cBfWFScdi
5+hDJajuovY8KL7aq7kjXX7fqqsuaNbki86nDb5ShhyQmn9A79IqJSgZ7TuHE54F
qIP4vZaBNpUSLtEOZ8I2ezVISbQR9GxaZvUXQddyt1UKO1B8Q6e6f+mBlWIsVemj
A1NT2EMYzEiLsfT2/jmT7lWIKIKg5ks0XkBWnkWcx6LjySPIePFowLOkQRnR9qdm
9BLDxPibMN14VoyKFP7f2TIy476FxlvwrKCLs2ZbfbEQNpC8ddAIUvBWdY4EgaeF
oQA5kcRnhuXwH+97uR5S8eiXtxRTIhuY39gSAR+baV98CiPHEIevrd0qPnNbIEzu
fCrlsb3K8Rxd1PDOpiOV919gXR3flkzQKhdXnVS0finOrL+Xi6lvzomxJJHQlcR7
VuB2NmyToZxsm8TLsikCDMqz7Itt2LYJFWWlDIAzJysgoVNFr6ocV47132mGGvfX
lpqMe6JnqvAlcmjygoZIs6b05+rYLpqJx4e1Virw1wbvQ88k7+QPWAiIzrjFikyQ
N6vT4sTz5oFLAR8ouN9bMvt/wCqTk2Fb6sMdsxPGoqxKsKYpuv7YfB1Q00K2y+rA
B2yIsVli8pBWQGmjjtPA0TskcTaJ3OjCAPOgGJyq/zgZ4nygeE3ekRTMWLoD5oCI
icT98KuhMlyxgecQczworIrB8zmeX8bsolP4razqSNKtSZbNgImF+DjFatbOV/d8
yIuZZjq8HR1zTe38RLzHjU4FE86Q/ViJ9RKwbLQWcCQ+mNHEFvV02P+NPrArC0kW
E9qbp7C58/nUJlEbKayET9NTes/h7gY6OoY6g2otjNpuZDFyoYQrMeJ5g87LWHGk
5l7xYlGbjSV8jqmNUjbBsaUMkPGgHOn4x9r5iXu7dojYpUip/NIrOrsduNt5jBqs
cCxd+96YAXujpSJzahxI0u/t3WLk2R8unxq/Vl7viYqbKGzWzfwXVApk+nK0kAFd
pnC+7TVN3NPWlaFIrzprqMx6gFIr4KznZ5WZZza4hkPBKIJYuAsKWRl/1UQLnrtS
QyAI9pFB7W24tOrRrXP5DKMIx6ee4b3kMLZEp3Dvr4uzL3TC8jqplShdACJII2tH
MENGDtaD/N7JaM/XNLq3n2RJlzVCOGbNq0a01yFVTqhxo2LXUSZZ4fuOQtpo+AJp
CiryBaEgV9gR9mPffKN7RHFEpK96Nipj3UAnTpz4FMpPVP7/ruPaiGrbOPDbAuku
+lWyUPaB6qS+xAE07GnDvhdte/vXlHiPBsPlh1Qfg+PbMa6vmtsqKF0/1Imc9SU6
Bxfx3ii3W88iJCD5ld8rymbzKWwDV23fT9rPmmQjBvqOKeK/cmtDQXidEq3lHYp5
K6sASHaFBZz1UmObX0kf5IcBGgLnCENvWR+IPl0Rir/qswtSh3kJo/gG3jmoF7x9
I9dbA8TEfH2f7LiP2FCMMvah7maG5LoF4XgGe3E1etk1UR4DmjM6dQ5+29TIuTFX
uCle0i91ZGhTbi8cmPCB+HGmAODW3GoOIcIxrCR3jSjOwjYz9jfr/L0ZzJzm1eik
mJwCPYXpQlRDRQAR231c+p5xj1oDJPZBwIDwmmBUuJ8xlGJghgTGWEeHNqIniEtP
siOmDTyVASwxgkBgP4qEtRyc3iZLzTwERQkQL7ucc8SdpSj8snyNEiy+QI6x8spP
vzZnHmipuh7k16cw1ysECtae8NFneSTLJMbzCov6qfdfJQV75S6vKbSNxvVnjHFe
kx8AcYb04nZPT7lv3Aljl/yaNpEe3zNRlJShOyBf+X0WlChRnhRbhyVLhGX384mP
SVM8h6TWq7B7lion95fUMC0W2iEajgy/0XUyw/D+C51rB3QX4CpWZ+P/E//OKMVM
aUyiKv53vXmQ4L1gEISO2UuGT2HpmjQ91aJYR09bRArREv/ELvRtpShyA3rxAoii
KR8494CRMjckokusBuHBgITXJzhTFZIpeEU6xWcwrXsDBCsjzYwQd9QzLQJXmyYV
5AU72GAjojwRp9rqgFgRQf2ezCySanL3wVGQpSw1KQvESoh0wteHpZp0QklY+Zw0
m5dxXEIe7P7ZlnlaiitcdSN9GIG3Lg7XqxWnCu9bA9B1qfZUZKxbYZ06pBoOf6kE
upXSZYEe8CDI2e19+CHyEIHxgNUKOJUz5o27vSTd7ARiKR8av1arqjy02iMw20C3
SrSWd3/9HGyrJEcaNqNFcsS7p/W2q6G2SRbMxlgae9tR8LJQ2AT2uOPoyXczE6zj
l8b0cTHzxmrI679Ye6V320910y8fC4PRBh0JoA6cJ7GoARo+wvYXm+9QIsb9mkHU
WJBq9JAZ7n0SjKGnPvVxhC0Y1VRA55HTPGOsG9Exiekr+HibRlsSDkdSwsNECHus
TA9BZyHkXBfKCLyi1X/rgKR5J/nCD+5Wg8nGeEFwMcTaXh9EkmcGraYiSEU58Eg+
9O5TDYAed/u3cV/AJp0dEVyp4L0O39Y686pU4Advlr+vMKrzHG+DNj9RPG97WSX8
ZSWpL0cWpwRArnYLERQ87oA++WJN9zcdMD3it5hhSsp2aoVCjOgdl0Rny/Cb9CAh
DkbdHsoJAWQHr0Itjh/hli7rejqeNR09AzYVKHJjYLi+CUI48HQUev5p6r3f/KfA
xhDghLWb3CsYcMYuHYbOf4CdT/+vV+mtAj2VlYlBk1puj31ZAbCW7XMdU28foWQd
vD7y+h6W3Lj7lLtl6UlLCRqYAT5utrs0wN4rlbNVO/N8MYO3A+kUrDBQ3Ju5V6n/
Y0WPO3F5fEp8HpdGph/XZHbyNUJe29FKCRAA68EYMn7zOEuBaBI25/2dEo/r2058
SJpqxW7BW9+A+5nR6G8n5/TrdDjvXwSWndgEA1a91hV8UNptRj4FfYoD5zNs/aRM
EP3s9iXApV91lVgEbh6xHmeCqOYDhtRCk9s53G0BbNh0B79ETgYb5Qi7H7Q9cAZu
fMQHufHGHU/ZPRiIa+PkgY4Ag0rq+pQL57gQvMQbCCeJV5wgEgua4egBdEaobClY
1Lir6kVPemOzQJ5bLLqtZQKyptxZvKtm5n/bClvzJbNXS22QvqaucPN1C+CRHjpA
TmdnLHQxGj+Z60kkg60LJJFelaiUWLKdYwPaXa8wufmo28rcqcJgu9EuCRZ28/nR
qvv3dGyvU+lH5UNE6PrDUW3eMtIO4+0kHOo/mRsB44S+wdFd4k3voziJN7p+7LK1
LhfJBveOfQMeCaDJnSFZTiJsPawkbwc69haYtBGYmZcWUNI+0WDJV1RJgtyAxVBo
AgEzvgVUaMVPzcAYmzT5Gz9F9Tl6tAVf8/B3Kj9cEm/WTOvRyInQQAl+I8QdNO+z
uBJdX1uCWkHn4Y0Eakyya6EpZ+KqGAmXWE0RUQAZvgFoBksteCHLGUtHvbzbD2UK
9sqZrncYlM/Ek2I0hjW1ulChROP6qQVecAgtSoJUtjnMl9dDJSsWtDhTz4SujC6t
sC/yJDdvYaqTLiI15g1dkaauaEvg7UAeGkrFRblcxfDbWQ851/f67Oatyggrq9hO
W3/8Sxi/36vG+v+1b1csNEyYj+7sWIzgvljQk5z//39D7E9VNvA09L7ng5CZn7dw
hqX+GlYzVbwEypmxz/+vAr6aPCTDL0aSVxS2c61IABa8DKO6JoH7VBkceVLBL/F/
PcihH613L8pIHnAjkGJdYyxKHt3phvMKrSI1r8rXzMQHkjaJagX9mEQs3tDgZja8
nENTqNTBVrWd+iDUBeB0wG/vZfqNd739ALAuccc150wyFvU1Aat6+K7mfZUaQXnD
oHPykRCUSJRm2ZU4hEVIqlphoANZ3uhnMfO/05OBoSHLHJr7AuBN59bEhJxJmThM
UnvvTVgwqapyMLrqVTk1t5ffk87x2EJZKK+qqFP+6sVG+nOISeEXkU3DmBswrqRY
nqJOnWAQ/TSR28FluU1Km1n2CR7WjdvFRYGG4rYaw3dSqFs05XQhwxpWWpl0IHpc
UbYR4HCDXwXGa2FYaITEQONurQixhhhvDUIQVpomMhndWDe20JP3tl97c9E/Ei04
SnhkLUVIJuAkWM+zf5/w8D3zDmgixNTCxEvchFqXEmhOkLK5x4Rq8YIQD9s4hqvM
FuiW6xW7REkssyTdcGEc0QMI59Cqmq+GX2bJKBGvthb/HY+dCjLEWjcoZ2Q2ILS1
vNN+W2j/DXaMgrzZ58BWw0tpM3TDmrZOCDwO5ODaAT9v788T0hRFYqnP8eLJlB1n
g/RMUbm6yTfUe5PG3wUCGKWG5eFADlBtIwXh1/i4wxbwhs8qQ3u5Hagaq0o+oBeT
uBgzSkw8hz/8aQbFSvZ3c0aiFpSkqjn2+p56zGcasjY+TXaZRgOq9y0vNaHObz/7
QbgRHFikNZ2VTt8qI0cOx10FKQCNRelk3rKcBY8+SnMdx4SRZHKX/MYxmNtA1R3A
RG+MALq63gX5Bat0+jl01WDacB8QaKV4jMzGl+oa5gKSzwDEezTvrY4sZdrgV/HD
BXUAw77SKR1LpeKJg/d9RCTlwzGrgLNevgSCv3e0aFayw2TuAYydBz8fpYJ8UBiQ
71HHAr43/2BuC8Tvp5l7BmbCN/2J6CcQoTD9mFuxi1Boa2q8nGQJE4EMJuORS70j
tgnxCoDOYfQsWWTRDZ5qCSig3blap9xBUHd9RUSpmv0jNiCPy9JP2aHaqhVjt/oP
WHLLM5CTaULQpIf3gu52jU5vtxwVeI7BBvK7FOELFSfpI00/8OWUul/H0qjMioXt
AtntB6kPTiml/V7pMM9faP/K7Hd4kZKON3n1Kn6YxL2/8UUba9OACrWh8CzgJu1p
QoBWwxzfferXV5V1z+sw+Ny425jD2u/a/tPtARDhvTdLJ9sUkIXFZrOHMuAS92zR
lE07bwuj87xTk7sWrGyOe84shvr/0ShxDJ4aQ8G9I58EpjlkcpKQ+dbZlu1pz4qF
SuwRj+MF+Ql4fBZCRAC6+cvRraePFHOdLEbgCHPQo5zDePTci+uc0olGkeif9Vt1
bFIjMjNy2DMfzedbYmOH4W5zIPE3JJa9+ajMT1tcVhDHSTR8ZYVZYCh+biGFL0ex
seXvKmIC/3/QxgcvTiJe/FFun6Qzwpb31d8ME99ZyP/6PEPrPTw55M23YObxgVJP
ug5wMDIWX+ocDcmDdWFuNa0CN70IrcVySTGbondwIe6QExNFcQNpJbSZjLOq+CQD
+05VPWe0b/xWG5rFve7BpvSh71kQvqJuWaI+n4n51ym6gomZZ+q7mhbvbn0WrGPO
rtI26wDZoYL+20kp6K3kO6eR+ky9+FMleJ12vE/a+f6ZKvjtatH2llbBgzf1ApTi
QygrEMLFbwW93nkD/L3mEzJLySqkIgJUDXRpHHhSnIz2xgECDMbSszGyEf4O/XxB
TnznO/KGGOiS+WHm1u1cjUI9VcHheopDsMkY15y85ahCSo4A9EXD5AdgB1NIebZq
4cLo0pZpN8FMoxo0h32G0cm+OGlvpk+EYM+WYAVme0g4XRUYIU5Clho9sLpOqjM0
L7repsENFCa1UXxzk6Q8ittCfMHr+oqrD8lpTyKkpIs16AsvEnzcqIe+AZc5W13N
3u8fTVTBNGzOq0etc4i4HR6s6PFAWRjeciU+soAUm9B08diqJw2LYeJ15nZVuqyT
D0SYrbg3homkP//+sKrIsdj3tdIk0WCiR22WYdaZ4b92OTtluq0koh0izWYZW1ZE
kY/HNtP5o5AVolDIYCcSOPMkpY9g9YMI24+g2ebcWXYGUGDrx6CmXLdcmNfZqjPN
CHtYWd/3dLjbgTPt1cWS0Npeti8qtRyMSnpGi5W5v4uuyPSE+A2jlwK9NomgbEkk
DrjyggDiu3thHJcHy8etd8yyhhl+L9fDfaRsFr0d4oJxCGijoer7a/qA7d+PEame
LePDIDT2KZpNuI5lOCWInOfQYluXokfGU+vh4/5xVGlEeH4m0758mkIN3vUrQPXH
QVOls6NcrJRUjP3tUGplPPLS+lMbcazcQvXXdCYr77ivIjll4rEDUSclByaQla3X
ORfRX/lRv8sZqqidSiQoPr/LRyISlz0fu4gUbwi6qDRAYHQFh/cEt5c1iOEGrJku
h221Qjl7/sVcW7DW/iuzqhkuQVmHOHvW2+rcydpzAyeo9GHXtFEygIhdDFn+SMY3
Cme2YYFtheHO4Uj/evCTAAJdPQ7Vq4m0ZcxN/w4uo/miE3expM4gj5PoAyftsoG2
90t2bAC9I+CJ9heMEYfp1L9RczX8yM1fxEz4K0OzZp+uU0wHodx1O5LAzczApfPO
eLh1o+0X3ZPPkWcvBbykcYLZJ9CV+3EH7yXVLsZdDysgIJnldKjHGBdCBkzm/VoC
pPqRfMFYshs5dpgEvpPyzBAeenZgwKmEaWwEgz04295grp9bExlbtnDF0HRkiMJN
jZ+bDfCQjxSHpQlEDckHC8bMw7B6uTeo2kkBEqadE/DUDFRJbn3wREHI/cFp9QXj
3I4nTekli+BOKsYODY6LEiAtVzhDSZSNvKIVO+pV5+4Xx43L33ycllJBPbpUVSG9
YOF7yGKj7CnOoRoX99ZNVLnLHCcARxIjcopkijGqOcqIQ8rMPN/KSiQMD59U+/Gj
uJNgyBI0Vrl+ISuZCbJxvUnhiVXXCg2UxZssN8fr82yGgKslVjvJzjsKODQ0bMJm
iLhqQkm9QZl9E0rwWsMCK/3Ea9MIG3Rtrc2Hx5vDcnRWb5kVq3SoCTJSx2TcPv6h
bc4PpjteaC12oifzszJbeszLVMaOIyODQwd7KlRj0pDDS7Tn7wQ4iodyADqyJtct
5E7a6mp4KvySVkFmiXYNYg5o2zh5JSf3jOjMGlMG606zkMaac1pOe2sSzgeKQFuQ
d6myf+kVXK67YBYTuX5satNhu0+PYIf3TIysqEJdWk7Uxic0rbLgNZf2+RbalOI9
qkvp3DFXF+11kMHERgEJXK6kXgOE+tfDIr6bb0qKz1MKZCSLKsR1KjbhfRvGgCQO
afB+6HCN4dPxhHDSy8SGRa4EPJ7vtK8zPfjtSRKRFGUjhH4qqydF8BPs8mC5tEc5
saq8RzgYPdQpKhpIRnnyGIFXiCfcnwMuspgNnDbhuOmp382CBixcLQ7N1L/CSIKb
GztdSqxrJ7sXeHBZxpwaFKNvFnOeGxkfFI9IcdBbWOiyHTOGFEIk/A5fh7JRqRxm
utMyBpzwy986eWKKIkAk6Ut7YudD7MUsw25MKr9aUzVAL8yy8jZAWKEmih+YMdmV
pBAP5bkkpCS4Zxr6SClyPmAsZoz/bvJ9bGTWjYxAnD7b4EMt36tOjTTsMP4VCZWL
Pk8pg2q4olAXYmyysDbxSPxyhPVfobRB8WmlvmHyjaWjhY2dDiXA1OVI7opcUe8F
MsJzV2aDV/Vy4uDw322WAJ+NiRiBJ5UvgKSTBKQPEjXPzjw1YVhze3Ui4/2v1ssj
FsFFePJIigwj80LVtBErK+AaMsGP++1hpqMELsybvR4zT1PWtjqY2sEEwGKy0ORD
h4lABTT/0dW8y9J+pZBBh84dyhg1vHeaY5kAIpuYSeKadvoY3E824ERH1kWNTqyO
llHLR4QkHcygpWrXdZswQtCjmLbRT7/nwnf1rxJf1dVFhinPnu3cT7Z2UOfrvytK
fOeSRP053kBLgGkD94xHYbYT4Oqbt59NslgH9qS3CzYjmDyjlys+50Uc7S35EFj0
U4iSxaw9W+4m5AeARViHG0QosLq03+WCxXy8mjdVXd0tZHiw5aHIuwqyf0yNL3/r
ZDT5GIQQZBpXfbp0+qfVykV+njTuS2hnNZxod30z5pUWJjQBcS+jDeu2LN0dSoKl
sIg4d3GxPZqNLALxlqeXb0jPdW+uvyFF7R7HVjYW7gA5OdxHnJPY8VGJSICjikk0
Nwk4BibGutpa/iN0zXokcLqmO+LlfcZVN2fKorASiUlLbeGMYhalfFji0LAEopbE
OusguYlwi/59z9tIBvVuFpK3B6JfGhQO4XwooiQMw4IonSBdIwXuvpDu6CrerwbQ
oH8d7gNe4kW1RZ/qxLk0qz3bwiSDRstJZjmMHTtkwEu+7UixZ4L+8MV7X7hmLVg5
G6fD6lkBHQtmzPBLG3W01usteTPgkZjwCeCSBFburSYNfowGYWiFQOVX0zszFvJQ
fXxPNsh8VoHn1ioU9BYz/mYwU/VMS8arHBqlbnjvf8qoW+tw/ru2AZe7A0dymYd/
JzrTuTAZsnr2U73KIeKs/JCgHG2Dqb8RcdyXg4d1iR8cvf/TfzqJtHaqBYOBs6/G
M2421uKO9YcB1NEhUdDyNcfD5e/PtO81n+e4QgdYbz21gT0l/se9yHa0afI6TrJZ
HFuFrMOQTqxSW+V8VblKeJ1TR+rByRVEKy78ObVgV9afjf0JIc/RSRQdWV+3IKl4
mTspmSUgDOwu4rwYg2yS1hFhS8Oi5VzDTqb01ODgi4Sjcksor1TaplXNHu3h6/zK
M9kCv56RKsYU6nlIJJpdPqfhioa1Nud3h/4XXxWGzsPIYwLyNt2SRnijCqIN7Npo
GQbKEK7KOFt1/NsRDG4hPjR2RJ9vjpcwrdHdN+rPDQUsEVEFWuRn7FgowHp4MyXA
1FGlFHljYaH9lOOhmc/js3WKrMVsjL19mqyykl3gSnic5tUhIZ8p8Gq89SWjhZDs
pd4Rl99oSDYyz9g8KI0Z0GTn86fFdUEOQeI2MvmFckhBHxc5Iw/c1+ro6y9wAaC5
KxhLjMS2UR1ioFFRgF0Xvc7znJCtjWwUOyBrfLuZxPOEWWUwKu6D7d00GsKnZAmv
ew6NC1aNrv88+UD0qQmL15O4ohcp1raR695QR4V/alA1cAFCJvBtmbtYUUiJ+kVA
d4JkHcWMuAhTHgaBRQdOhIdXfyIFhQ8NHUZ+HTY0XovfJ5LVJyWbvrxoHxiDExGo
MNyfFq8YRTg4C1ETXaQcojhJ4d9eDIZ8cSDpDYkgEiKZfI0zFy/oXB9oA2/Djo4l
90behDIss94biwUGGfF2rXLOqir+6+DXsOMtPczQiyBPnI9uIpnF9xG7If7/a/NU
rMlJKsOMKim5TlS3oXwfV/cmTeejGJQ+WuReue8FjZZ5b3w7fso0pMbWN53JDfDT
UnUld3EKRTtk+/wDd9w2RSs29VwKegyusoI/j+BLGuo9qJcUWr9Q9ii7rL/Yx1FY
ocSx1pHYVIR9hticCvjZnHGcTHpTka8Uy/0tXBxBG2tE65bsCiiVYI2u+hJbbJcC
AW8fXpwRdKBNwGnHQQi2aaRu/amNNDLvPBoYKuNILF05UOsk6J6vtZYo4Ujeshbq
kPP5Q7IBiTPON5BZg8C2NmBx5XaDP3LmzzaEHb2khcB0B/6JPWrngsfHuFyEREux
ZZaugMilT/MkVPCEfto6IZjBOiesmSm8Rol4uWaoy4fuVW5Ph39APgLza8arkNJu
KYv9mHp+bkL4gMxXLE1XMEd8GRzS3aTCPQ71Z0CL6Hvlzh5vxi6E7AOBCxf4kwwO
6cD0/AETZKZjUUbRuY8YvmACOALhVsRVtLsm6nrvuBJ4RW1M5y+hAx2jRmisly/L
xCm0DX+2w6SvuUXstUc4US5feknh63vnE4wtGL9Bb+E6vzXsBugAyXEGh37Xv3hu
ItmSCqYkbSflY6dbYWqm94gdZY9sRP+Ld/ZWbYzcOY80Z91ER71Sxcferb3BSzlA
628e7KpZoRuU8yBuUHm/w5LlXHOs9IslW3rJm08/Ruz2q2sPuT5rzXS5mJOEq1T4
TtJl23PghuSkFtac7gngqFX54UNNU97LattXJBYZwJxSA6zXubKqVEgGOyyuc6IP
UUbvE1D5j+NXgVI/q6m0RZK1IYm5hZzEyLN7/erEu2W9GHUG1tAvLymh1JtjMAZ5
C0phFRfh0e0/kL+uYfOGJG+z9rwtr9rwxfxn6TijHcGwut0vKgPFqL7U/dD0F+pL
CSOZGYZi8yqVWvmIcbewdmxIF5Pbcdurg7580WUR+gEj5c7QlfPhSHPfNa8x+PSr
oOSrQfJBT4fqN+MDA03fRv35idSILw34FayRiC1i12yuxHcK4Ci1F+J8afnKSSES
SJ0anM+EBsBee1CR6MYMNNiNj7tSTav0F7UGiiO0ezYgF8uWu3Cnge1nj/gxCIIp
0FJDDou+/XGRTbkHT5pxpudHbNGIFcP9C8yZlgwnjbNpTdqj+4OKNNH/mNTiyjyp
d8CSoDZZca07tKYrui6UOTYRZqciD2waoJb8drka136lK8EX53omlPzBxRks1a7f
Bw0uYLTLjWi+vo7hAL44Ov3tblRQlRyrjrcHHG6BrkL7DKoDZPhA+OMZjylPaW5G
OWBSE+yoHGNmXtf+yBNBxEHx0vMOqKKJ3mH4Z+tNGfCclC5TmAGhjauY2/j7Rr7z
JwZiUKjQ3ZMXov7R1539beMu8YnLSuDuNG2olFf+j/rsmk6yvDU1pCJZiVld3lTi
kP5sWZ4UiKu2sJshJRWiWdksk42tJxjY5sEDVbzuYGXNfXGZ7vGQJ7PgwYjRhF0Z
aRUxNoqhvewZBmEKNNqrWBEf7kztwYOAmsuGkolDRE0dgMmavlYuWGlhZNQN5R0t
7yOhPBUAKZIq4OOJtn4zxlFLBhZMDAL9H4X3NLFtumjhv/x7mtN2yIh7aeY8HUam
xF+GW9ODYl0qJP3rMjmaPnd0a1cXM5dxUGn6v816HlEcJxO/UglYTXzazYd24+SK
SnBOBPQHmb60ui9MPd2ZKx1VpZ4HlCGqQej23iYz/WuQT+hGQygXi2h+aRW4c7SS
KCJncfZH34CgjBDxaR6rzBfR7KH9G4Kj+Y0e5FO8vWL044yegWrO0yEIhn4JPYZD
q3bQ7vX0zUVFuihw9QiVu03OJ4/2LH10TdRm61u4uBWacjHEf5Gyx3qnzXGXpRMy
BTqHfjnQS/j4PnDz+tWmdi+UMx5xPLhPgAyeCc0Gq8HqBVunhegwENLnkk4cPiSf
LIG/w9KPjhLyuhVkYLUC7v+Npv4/h+QwB9S6PTM+Janpc50d7nesIDomo2GCQXTS
djTjLKc6FmToVw4/FbANO8/FYRrZyJxiXgUq4LojIPXE8xAKK+S/iFhmItVJ6xOe
54Tzdq7+zfpX9XuJ6fFfmcm7LN1xGfWhGi0rsJPL86FNxkNd3873NLBChfeYuROo
Izg7fML5BzI+JcET6Rkj+gYOY4pXNFdPofqPVs9a7PZyzk0AosFwwvVYgq2FAmTv
yvyohbPDuBikBUsYS69ZgQtYmS1sSOxbdWB2n6FycX/wbYSK8uC9m6v3rcbTCZmD
5YiIGPNiFhNRaST2X0KVlRNPy1ilPEeWJYMJ0+rtwyWasORprUfvK0aD0XsdVUe/
4hJ1oL0zw2pverLgeFxJ5/pUZKz0ZXdmZIuMewta1/iKU3rOgeHJWUKkexrUjfsh
Hz5Nr/8yDg4DVfoDmHrr2qUwSwVi+YROanuDNkUX41NScbuLjOEIuezlhFvQMtz0
nK1Jx6CHBpzzotN/Qq/XMrm0wQOtX3Wli2mtyItzglZ+NvahQBpmM7mtAcJOP+92
8zrNCve5dSNohgMTNbczeCuE56C/pWW2PPnrdTmWoPMY4RFrik5Iz9iXE62VZ4HS
ozcgmHYMepOX7/1hToFYIIGeHJRjh79aJlrC1y20mmpgQgeZ24fuMAFiv6EtWlI/
pllf/lPbmxLetlSSDKMlv37Qq4Lo8dILPCv1zQXVsLTOHbPKsuIJdC6/lH5nXEev
MRg0ZChPz5uni+6dZTMmpN++F0JjTaYPTdH5oSzN5D3VsE6F1dAUp0spjXSs8hTr
BUeF35JP7QnVjvot6uw4Hs8YbUG2DSn9o5Zmy1KF8KnR2eeFy8n82Mqa8FOtEl1W
YwDmvBI4INVubqrpBsLtmzsUguCiRJHpABJq3HUOaO3Vte09W9yGT4x6WiUR48tt
BHve9BoAr0AKUDKD+HS2JaNkrmuKErzJ6C4JObyozTthWsc1jKXsxGplK4K5Amll
9JPOZF5OS3vi5Vf7UEjSbNZaUXTFPT8ZAqV5ePUAtEX2m6rdCYAdCwFuIoQhWoR6
JUvklLhp4N+MNPEQ/7WhTi68qnxeEtiSG19iPtcAIQyOu+nXz5CbloGsP2KBvv7m
ZH3iv1LT8FkegbdhDfAyFQvxKkWlGqdjIZeU0WZzSGeTSq2+28XgFL6aKDn4qbbd
8WWVV3h1+Q5RG5+is3xUtu8OydiILx1Pptrt+0k53WnD25hqg6CR9SBPifiTN14a
bVhkjRWVMizJUvS+t1ab6fI+zhtblPJv9cNVahv3nA6nUrhTmRCFacZHdOdhyzQ3
uIJJGOhqAdDB+vdKtI9IvhPvy16TLghTb7tH4PfaBLcIvi3L249WtpYT45MLCUUi
CBKOSigWf+Oit3jw5zuSATmTO04nQxBkYiBOFCSBkd1fqPRyqXJK8EYgNdq/xPhg
Wc3lP8Xj70+3qdfM0uc3c0DJwKOvqx+CdqGMFEgopnMv608Qv/FAsLjoFcnvZ1zA
3jpgAmLvXB/sn1DKc4WPWEhuZpen/9t632nbFIXL7FNvXr+28pyJ74YqbFBafpG6
BKKthd2Ql8fHqi5wWnD6kkLRegbUFatGjnU3eAH+MuZOHf5DF5JrZzOyObCGgDUK
yB3tnJoVDTKnOL3nVAtCEcupq7zClrQVUC1liBSO6Uqq/bAru/HMG+0yJ9qyO5XC
KBdM0Ua1CVc00GgwRZqoXD8IifkDP+aqS28IPLuKS352IW8nKoNElw0eTMJHE4iC
rmp02FW8hkbP+Urc+OZ0HM3/2cI9Db61ebIX+dpODWchK3x+bR8wtg8/pDl71UJA
YiaXLgvg7mwTeizYivC3vmXzD+2V4VrqR2Exvj5zBWX7ZjpxovJK/JHOf870Fwt5
D39hm5JnPAsfmcYGYVYPjF1a5yozLSfVievLG7C3VlJ2zxE/DXfvO1e0pkRo9ZCq
Yh7D5L78ksyVNRVULqX6pUwyLXNS77Mtn9jSXH0dKIzDYl6WTKIlgTmesRcNoSBt
0aMluKB+cbh9uKC67uEtQoS+tXiNpOKot3vLMLWP8ss67ACKEopBOmANQ0QzlKuN
5U/yf4+cBKRI+oKqFX95I5aeblla2gPn3zN3VFnATgEXOfY9lJ+ZGn8TNSa17NdQ
BU2t4k2pboTIQhz8EAQZ5CTuVAbTcb3hOM+SsF4v9GjJmNm7yP69aUtaMlF2eaaJ
9o7zYs6zc7I91vkt2n3EUfnkmb2KjwPOGD9yN9QMENFAVgGhdwoVyVqbQ41tg2vc
wmHRAIxbIjlznylg/TNsGmMAplGAmAG+fDrBuObehyzWILkBiEeASe81r+6UP40g
99dyPNulSbhqHWAuyq9UCCTA1E5CwaOCyqU4ckVFkoAUx2D2A46+LWXG4/+kwN/s
Lm01xQFPEO3L2cCU15ETXScNboa3PxxMcifFGR7javQpW/BoqVY6R1rmKzfyWYMW
MbNwonwL5GGoGpI5i41BBYeeLB5Tp7EKJALD6rDw4miWpnnVymy8St3VKKlH14i1
j208gvyxhRBT0XJBG3uMHFgfnNeNTXVZ3fDmUhv+gm9z/R/gXAdVTNmCKXD/FDAQ
GvXfT6qHocAFY98Xa+rDY7oBTC1WTvMvAmXTAjFICBmIFhx2VMbMkB7tuMvl/QOk
wdAWxE4VDfjpRl0IsttOVDBuYXWpInVDTI0+ifnkzh53nF9/pKKYvDRTjdEfS9D1
YhLHi2wdvRoPTNPsktCVjX3ZxnPqPQMOfDvhdQwF7imtzmapI2BFxV1E65RLghmL
zMkQSsOwpwdDbP/S2Wp8IvP7CFEFt0MIfRX5OpyjC25aDwG3LEs6Apk3mKHdLu+X
7nZiNTt+QDm/TPwbVMMBjUNVnUwAjQzG61ohKWnXtFpxSAxHq/z2i8ZHw7VDHgmI
vh/JUCzOUYLDfke9sH/1+8iMo3xgr0A7EO5bvsV6OZV0anYCl8TBv01M8YhFmhBI
/uZ/AAWnMQopG38ghSEQJfe3hP2sTgjsDotVV8ex0NyYklFhGhtRtDSsq8I7nxik
3htU7eE3wgPWL1VXeqUUScFgP6wzmQlSwbxwqk2S8S4K+xCNL1wWTbo1MisB8VEB
6cU0vaELIWpP6IxppCSPGl+Y351c/PoZVxkiIg5dqL8TPt8hWP3JR+tGNlFI5N/+
V4v0sqMKe3UJ4J5a7csGFTElIwXwTmQ/ARsTe3NeBlZayiIw4115cRn5n1kknSZu
Q1VFc8f8u/4MQF3EEwx5TOOYtdNQoXB0I9TNxlwv2OrtYtYz2ukj6U/6omFE4XQ0
fc3TpKwMWU1wwgSIa71BCulRSezKHTnbF6ncpCD/1+3eDYYZaqiNYFfDLr0ELD4h
9Xaa73rH/JexD37rRMRvGhhxOuGDklNZ/I1xK9cV2iimzzxq26IeBfoCCUw1y3uc
UcVFVFc+SWE6KYN55dJZ3KkAVrrDN3aFx7PBI+qMUSZtFDveSN+mNUlUqTzuUP3Q
+m+V433fSlepLzreJpDAxzK53Qdvjc9RdtIh7q0/i4bL8vvhsQnQ2K3OJVlz7G3s
RFrH0dLJYAOnsOl1LwW+8Q1Sx3HfGz73D7I+kfybDq+ymMrirXsz5c7oez1GcOLv
hsZdEW9Vs1qJy2wQomtAeEhWNeV3h7UwNYlYQDNwMRlO880bjb6inWh3zHIQXfMd
/zPm5zo3H+YLycrvgIOvst5oT9zXI62tXXuFxWrQYgoYPDskMxC/j3BDfUlYvovE
/uRviGPpGbaX4NsKijarXBPVtc1NmMuBQHP6imQX8KU/MFMysxHpZ9HKMYJozhsv
fUzDuzxOW+h/wzeiudsZ28wnVz2VunX1FnAHY2gkhg5J84sNdL6WMxCS99wn4poB
A+HtMguU1fAl6gCarCRrOI2Wj0Ge3pElwRUXN0TEnPf09KewoT0ErNVAo0OjXTrR
G4r1AdUQpSynkows/RLnO7/nn4by+qQhK/UNl4QnVRNcyebwF23WA/J2LdFVp2ws
89Svo9sgP67Z3YKbTMKg9vBlKka6nCmX78CqU+TCpr0COBeRrMT9naxmgnGtFn5U
R0H5OI2zkKQnphx8Phrnle31uuaknTgYCUKKuvhZr0AtELo4g5tBKFoPcJDqj2v4
4u2br8Co5beHpRVIOvhCakz+8wY24YZsdHiN7C9vUf7L+n5a3IpPyWRbQYinuNAa
UevDs3ylZsf/LbOj3sAqGbbEBFhFRp6S13ymCiu2rTa64mZJK5Tvs6wUlC4C3Idy
9tb7JoUiRMVCCrISLR+ZJQNc9gcH1r+1SsS5WbPplx1FVA3PTlk12x926e31tErI
gB8wMeIWSoL6r7GlbAvrTvjMYyvYeq8D2iccn7WxWO/WxOBoGkUJUrsWO4S7p8m0
5wp2EXaIJkaiNawcqNuwzJvzGc+YsU39GYI9L2n6vlr6j0HLV5JVaivhsRU4z+YV
GkVTrE1Gpqn30DvtIuIk2GNgG3F87fz3QVDhimA5zcgSaKY/drzYK3GGtHCgyZ94
T8NEifKIPfOA8LevWdRmjn96YlXPOWBxAecHkFGK3uDBu6AdWDsyVYsVWxI8Btdw
yWEuFvOfyPqr2v2UC0+ZZLRm8EDkpzjD+gN/QbB3/34Jwxp70ZdRZAnhTXbh1nvG
1Hdr3pr8HqyhP3rCilbY4u46yHrcHt4mEOseIPn+c56Wf/uFlf12XNfB35QAgFuX
wqXHBiY/8CLcokXOGr7n2ey6rqTXmB72n07bfBqvs3oF9xUuJuYgCWJpbspt00Qd
MdYPRinYwRv72MMGj8WdynOSO/MHk/EamyxABP6iDPRu0agXk/MgyVWNuWpNfXVM
eJmYcW7nbE3Ui8PjOcSs/IbaOcYdY1R+irlVEOU0wpICS51eeyLrKaohzVvBNMXn
UuRkv3rX3ue0Tu2Ann46DInR/QsJ/ykGKkvtcnbN3rVl2QguGtLUJ88bA5S0C37T
j12GPDR4JdCadEPyBkX1z9gfHvm/BbpJ0td/a58L8tA0xtlMWkhWePQRhgx3SAsT
eHIWT/TV+zZ+tGaQeo0QNpgl6svHZldgW8YWNzOxsE5VKte8nQ73wSRlVcxF2gqI
bMJH3i3pfZfKp0Ar4C8INRCW96lXPxBUD9uv+oqVpLyYWh3AQ8VCsU40s3tkWtLl
kKwOwUWDAjoAcIi1WYZ/6PMdO7Tw190lSYNARiIzdvw4qHFLWUWKxLLE8jQCSHc+
PbcnK+5uSuSI6s2UgouoqthSA4fHannexDgaDzfxu8/NKB7XbKHNxasOak+iSmnZ
euiUfOu7MJ23Ow3pDNlNG/t3n5lkQJCXnjxMPdv4nnyJqZCkqRZpJf38tRDjjXwB
1iHdccP+XWmqb2KDaAlvVYpx3e0XoDQh3K+l7GtBVqf3rYPBnAPqC9NArHSOolm5
RvXNmcvbiTpuqye6Hn94AZR+mnUjVQ2p8hPMcQWSNvM3t7w3rd9LnKX6HxhWufIK
G0fx8Ltzr30TKjPwPyTjv+hU4jbcLyHpJLT+h0a4E96uptUW8w8tanb69cnGrfnS
HtW3qVAVnRx7xikpm3VTNDpVVNV5wCxtkELHltvgG4Nt9UAOWlroVyCts8o9FpUV
CdPdF2rHXiq2GFLucbcUh35BVCUUIc3SDZh9G4WNZ9eImtzArWoRDBhCRKR5rRBr
YEB2zm+1gbqLTU+06skps5R1q0CnkGCLT45mx5sg2Z4DntsoywEvQKCKvtxGStSR
am6ipHDZ5qYtbSYmVrLpzYZeeA1csDocr9JXPju51TR69rLJr1Js7Iuqgq8p0PCL
J1rsZ0y+/Lvs+E6Q6KvM3E1tIaN4b2NCQ8aV24j6oh0laYip9sCLyCL8Ne+k57yc
pPkDZaAMse3t3T+O3hlIm+sF4eBh4PlRYRkTFluC8ujn3PDs5bfkItZ9Ve54TEJx
/80dHROa9nIQFDG+N2o67o6JabaGPEhKbuI9DIZkD/JMm5v4Dl0+rmAZdYpYquAN
IB+h0C9N9wjqGcEyz6o30WiT4OU2PwyKiBMTnMRJXuBbeVsE4Nv7v+1orv34rHyz
AWqm/Z+xo2khnbrfqjuPv2UBp6slt0+F1uXVMnFOsPO5D52jYbqUpogO9pp9HrS2
ld9amty3zx7XIoakH7E9VyUkx5v6+niTK3TsxbiLSh+JKTSvxs6yFv64C86uWglR
yGvSl5ev9GdAkJAQnv5wBij/wbMc4HDXnNxzhYIHNvMBbagP4jw5yaMPL/wpQ6Fd
wBxhIkDR1QLlpW+rZ/UtljFzTpGGwrw3sxQ0L4Q/BELSPoNxqt7WNFtJG3YGNXHc
gbFfXN2OnhLznY5NaYcKQs0w3stjPgpQcK1B8pnyksvmg6VNad7Hi6nAuHDLOxFm
BzuDPZ42nx+w/DZS+qqYvZq5b4win5Swwrle0tLDAq0qSIigqQkNCa7YNNHskN/j
YXrQOb639lNSl2kCoD7b/NuOqErOn22n4Ki+zfnCp1x1c7csnXj9rgywOwwBbdQh
XAxcodO3swnI8uTfL1K4jQMgW/c/jCFanYkHNoriMu7fV8DDl7mJTvFdJ8JShcu2
DoVEg0gkXBRFAtfCQmefc4VNYHtkOQL2KZFdJAYwYOYsr+gjsbaZHPtgO7YVRlsN
GHWhZR95mBRR0PdOK9/wVrLHFpMPonytwrDSuWNqwCLrHEkIjqgzhWyeL6ygZxDm
G6jmbGaL1tYRoHoH6KUko6sBJQ81TK4orFpdSusnd0O7HmOoRURywlrOERXWmBzA
imEAO7/ZtVDGqeG5NvlYs4sHnCRTY4DixtAC5HdsFe2njBpGqlGgSamZ0X4iWW8y
nLRlu0nNVnExpZyRCf9vM2/ij2qLx6e7mZV+NFPm9kp8eEM69Lt97R78LTalrn4t
9kFrkQgKrn+NjAa+E4+WUEA0yhxR6VD0FU4tCnCVkOVqMxm6qrSb6exqLMc+0w4a
4DO9AjcQ1WXbRTWjFGn04auaRR7AFNJE//T6I+3Q4C3iqc/tUE+8aRwH8yGAc6SW
sFM8hljiHp5S0h+WhEC9YFGJa36uQ7kMYJwy9knar3gfdVMr7xLR3CgvbbAnm0mn
T0cMG4u61Q92ZP+qZ+NrPvbI3irOo02NQXxLHRljRUG45RbBH9et9jYfq2VJMCFw
CVy318LgbJmTsn35HzD+b3zMczCwoNlFaIFsTLjUgDoHwHxnTHcOwefWR0QTzjyq
dSVNg8BzBNSsHLvrrEZrBHpk74JCTidzg5hNyC370HePHKyFG2KaKCAAzu6HLYcJ
8UWf9mtIaGunbPjo14IE2TYcTvqMm3MX3aTbZ2uF/xq/EETX+QMsiskLrNrrpXE1
bzxJpAgl2kdGy7z83ufUazF7pzSnUUo86LBdCjjb6l3Y9MeoPndCoON0dF33BQyL
0fLpQzKoGGEuYaK6d60PhGIog4HpNMSsXFrMMiR1Oi4FFz3BJGV6cThbtgaVU75Y
X3hmHzxRy5xG+jzwJy6zSz1ZUKPeiuGGuqSSpB5KsCVjsxnpXnY20pVf5V7fHkEE
eDuSl9dZ+k7Fqn1wIWgz7l/EGhlsim8oExWgawUGvcCPVXL1oU8tn+FYTwgl4z59
hWcxC8YtBJlw2L31vFrCr+5Akz2QO+UTi91o9cKgsBvyJcJf56X0tkFXGwTMml43
PsEa9U9+tDTUUmtrWQr+gasx6unxOyBeeygD2/cLgX7Spwk/hxlZ02DYSz55ikKr
mMGJBv9vW/PMbRlsUwLyzcZ+2zcCIYwf/SOIUgNaY4coTNlJ7HsX1WJQMhGu6BHt
5y8JEyd1e+3J/UBanHn+gfb3RVGBKH0ma19dgPOfeRUT3xpr2oPJsHsWwftzYObr
Dlmc6hhbRrKQAHRAlDvG3PSVhazVP9KzCb1n+oAdFuTklSJeHoGptIfmdl0GsLIj
tJOqinSvl0ambVPQ62KC9cn5LbqgHAsBqJgydSKPn1LSTRlFxTAeRcFOnG4QqC96
kd4qGQsL2DneCvBaoZhDjOXx5LxDckLTHSJr6Eg1aLQ4aeYqR+PZT6UOJjumv9ci
7RAePv+Ns/hQh8dbE8NIdQAU7HODybTzeVU1/mYq/SlCgNknwA9b1PlrHuq5ePRA
lbjcXK+QNythmHCoKKDWjohKp0v1wLV5GZKIPtQpIk23ZAlgpF6cq/n0y7eWJR4u
3ajG1n4+aPZGQylsDU8KSrh+sf0SBmMQqGqM6PLsfeeCbdlXar+VHSQcbYTiGQ4E
3laj0V5LlIxNGvtU3cVZNIujmkogjWH0JxTf0lhjDHP/CN7ERG8tWxa5BzYsib0A
4ZU8RAV5cJ7+R5wRUjmkjkiMxCvRM835CdFF81u1JqgIrhf9Cl5DnCYM+FzioBGu
VHxqdyHC7jgwMdtHVanOdaIXuRDrovG5rb9n/0Ugrx4bkLRRzCFJvaji56W1tj9R
yt7+IC9hhKAygK+jSFICFBlfdKUfA/fskXAz03+u3y6doDGqOF87r37p3cP+7C/D
gu730oX80ACNJGvL+DV9ZgSeR9/2DdBq7LQh2ToEkwXWaVhq+2PYcJw/2924gt0x
nc5UYq8KehIQZTqJWZa2AA8TROJu+j/nt20vctAQKTDBP9Uzs+ruyxLb0jVRXgbp
KUzgoDeJZkmKakjfjLxhVAXm7BP4NTK4gQ91SwCACX7d2bjdQh+ffimiEOZFPGBP
n2KPhT4dO7bkgQNtBvi7mVxvm1ZDszX8OP3T0U5zk2EQUIzrY3epfLH8ZaW50VOU
W/gM2ks/PE/OanigesBSeZeKIWj1yj5nPC0f5ysUpTtPp72XL90nqEiAsIb7T30c
O8Bm7m/7TMEJ9JSov2J5UzA8ejXX0fUZ5TfibVQCaUGrAQD1kFs6A/IoL2FLo5i9
4IedBN42QrekcmohjhQIB4gfyIjNHl+X4W/aq5F9+MJpRpzJFK6I3vbAC0vIgOzL
6KolPEiVEOFXNUVqFB9FS7UgDbT2PR5//hdYmnpIXC1scXv3riS9ElgG3xSH1PQa
nMr22bYNHQETs1Bqze3B924XSZhXTMOmlk3IrLM9CKsV3oltWiXJf6G8BBSWSdtF
fWr4Kg9CcM7R1u+DPHZT0x5BxxMYrhCFiiJ33iM7xzwdXBI0m3XGSUsx7K0SVTtq
SdHUlzRQPgsurTH2b8MnIQk56Q2y4ZtqI5V5iw5gqqEU5wMbL+BRvcAKXAW0Bml+
CztloicaLpftahsE6pEyUzo28Z17OkTkKoFBgbd6IdUCTQKwgfnQOv8mxLuiWEU/
y7tkvMnlhhhv3C/Lj7i5ZWNhxkoHdMwgo/ig6+N9BXmcX2Igy2zlypJB86e3owY8
rqyOJz/xol0t5JqJ4Ge0hDpDxO8Ex1xIzj3y9UeK8uSlXul5nu9x816DTpLdT+TJ
FNUhpBCireKJ3yk3EXdkZ0PWGeo7J3yuoirciXAVxTa2Xh/B1cyLy39lMcjY5u1t
IZHJmd9Q/Ex35XGf3a5vhrHZOIW0NlyL82NdOUMHkbv2Ij0wVshAfg2u7vH8gaUd
M46o/msgJgYWzY8NE7CFeK3hmaYQ1S39pQq2wJ2/nWKyoAa9bmfYanSiM6dzDfBp
YlKv22CcSUUH2i/d9HivsHAP/MVc9rc8hNJNgkdFZVLiby5qN5zqxcIdMo8jAah1
Afn+Yrchf6pI/8qXV1E2yVdgvtcwGYt9rebpqeZFEOVyMIzb3xzqkZtr03CjQTWO
+MsI4L96qQh4r6fduk3F++ELyiVkB4nRmU9zqFiHPwnlORSFkuci89Al6vUCss+r
MBp3JAOeWaE466X0SRnhrlvX/0kH4O1T/hk5h98HKkUCeGZiwVdy+5FOuO4vWBlv
d/YqDUIZFX6bLj1lRMixp1TKsZod8t/m16gkEUo7h/58tooiQl97Mw9EInv9ZuWt
n5Y51wQXPlRvh2C7GQsg3L6vCojn6OoKuLJvmy5sbe6HF/ePa5V3wr45G3+X2dty
eqDUmuLdfmvDtbIym7CP6WMkDvwIMq0LCPIRlAi2s2Wrqv97vsKfP7RMZZu5OODU
wKAU79iitmJ7L+5qp4Rg3ZDCUwtqv3SGg/TB378XacXvj8/tf+Tw3bHirwoGQ+jT
lw6HQ4WY+oZLSu54jTXX0sy1DY8WS/26/fuWt0LlodEXYJ/I6YtabqqNeEnkaE+b
JWoRCZhef8WJsKiExRxyNOihAjwivv7FFTTrEYAdHifd+35HEYIbjmWm+SUdn8bo
/VkWbmNPM+AS/qqTuejhGkN4jdpQqF0due2hfE+fUPPnCaEDZyUBL9bxsz+jZPr7
UcUwy9zv3Et0ogVsER3lgTbQ5dAo7V5H8BDYpnmGrQUi9q+Gge49rBkYRCDTg58Y
DI01kRMzF/f4Z76/8388JsuPODWdRAWkH+GDKkVeC9UKk8sCMY0MUwfkzyKoPSIx
ZLPnScjjeIpDkjZsxkzZaleJFTuv6TylTmfeejuxm2it4NZ9jS86luTXM4mQax9C
rCDW8gUnFLMANwgxRDB3bnReU4UiERq4l/sd4FdqmKL9QNyKmp82OG2Bo3aGobGe
PCE3bHv4IomEPG0AWgQo6Wo4dg9sx6NsG5F9FVXsY8IYru2E1ViJUUR5RJg8dmTh
uSKAulEHun0ZW9f2ykpw2mKPdVFLrPXwhDIKhJtgpU9Lw2yBnrfDPW2BJW7a8Ak4
NPQyd339N6j3B+yKoCOsxoKaX4jZTH55kuzWRd4fuAMD0sdsJqecNZAtVps2V9Hi
ziOb5wlnxuJJIjczgsQJu/oEAAwE2fUR+vAKIO/5I6p0C4ym65FGr1upGy+IHsjo
R3u4tHlAMPe9wt0kycbl8DFYf0KAsKGn4QnfW7yT5MITURVuautmrHpqnHAojErP
kyb32y03K2GOvDIk92APib9d/iJcEObCIbuuff/w2gR1wzJxqfdmtYHvvoHN0266
Y6V6qVxl8J3fkGM4tN3WLpeWBNr/wLc+IqiJEwF8PNSDjOdw0bvnJEP31PAZBJem
5AxwpNqsy0igIt1S0VeLgDELaYFyUnSOVASiiWJtSuwv3TBML81rA5D1qG1v3cd0
b17WR39pB4bjnJCGthyrL/f4baWI2FtSW9RAKx6lgF4Z3i5XZZuUaLveMhdpOdvr
+aiw9hjrmrFLs0UNPq/TQUEIu+ds7Uk5G8PrQPost15tN+dhNzrdUwLvLAhlq1qh
u2BwXoXfw4RY3yuKo5YfNasmFyWa7uIHpJD+VyBK8PDGXu90xwc0LQ4ckxqu+qbM
DJJrm9xYAUmNKLo2fbFPzoe5jLiBsMC6E9f9AeD3bsrGxZjO8A3V3xcl/GuADKUz
gM8IZdPQ1TlK7Yyv5UmXzTF/rumIjpsp6w0kTlRgmSpCNhVO07WwsH0Mga3a/jN8
0a04o73K2yZODBQPn2b2ePy9aLELwOIyAUftDpMwwJxRprWseKdeCw3HAEJ/OtCu
ij6/pb2hR1iwKi+jpKlD/6YP6s8lQvAQDTnzK1bZHIVk8QWNPqAYaNPPkj0ue7HX
aTxRzuB3XpmC5qTi12ltv4qQpKk7DPPYqJt4+L0xnzTD7mMSvAWOlIiis6MHLaOM
ih7iIBpfy2aZpYA4HbTfFwLGAiunqaMQ5lYJrkV+UeiueAy+vBwfGQ1fq+4EnG1e
heXHXx3Dsc4cG39tlz1uHnVY335K42RoWva6xW39US6WxsRradRYExz1KXGtf/1l
NQC6JNdZWbD2I1HZOzB38XGeWFPYlbCp/BHS5m3vwBXU2+Fjqf2EGQogw2gzA5cP
YFJxOW+WuY3qcOY3Dh4pI0dKIZodUJpdgSLsvCzx/EGUEZRE4zulw/Q7/86D0qFM
karxHhd0niAV7uA/DFj9U8pkqs166Ko7Al7gnBkvRIdvGMa2GsroMjHqTXVUxQuL
VxRIkEjC3EjyWcNag52kLEGj9rJ4t0DY6fHvBL+iminipeXD5e1NVtzEyu8NA0RS
UzYtgb05baPHZDRj0zAsF7WUbZ0Iiokn1TSvFFhj+g0NHs8gWN8jZhptGUOI1CnB
J1EY5abS0N/AiZFaSH3uVOOtzUQDfC+2aUF2rvyuphaaJRceqF3SNuHG+h6BNzwi
6edEHvxB6Lw1OCoF0ZV86saF3s+qkyI7nj0/jgK3j0iEJD3wgWPDzQ4vgDhseyYU
aiPAI0VGFc+iNIso9xRPfi0QY7dY8qJDnLeBySzLaAnyM1+hNgUBxoX3whpAFYWS
2Iaqun5H0Dp6bug27hl15em3ShXczHKC7VfxL5jxOwSrOqSyVgVxwIHNK9rCuAS5
fiQ7hI3bi1ARFSnsSkga1s6rz6Ll0lI6CnaRg/IPUewQy+kIkKKriPonGzamwt9v
pTESL3oc7lhVt2RKoNBnQkXjG7AXf1/wI1M/VY+vaMABgblHDgbl0EVRxXmB0o/I
w8n6pIvnXJc7DjZnt4RE3QCm+BT5LNJgHEAxE4BqBZaO8cpSVCWT15SctKsnfWSX
AbuvAuIVJwA9LEDJxKtM/4IjIjQQIk+tICbElW4DnsQbtawKnAD9Ss1XAT9NPBoA
gVPwSgTHkDiAotIc1iYsNDPu2C0eMZke+ftL+JYo8FN8qKKP1pDqepgefX/o36PU
UwkXb3/TG8+330v66UOt4rtYPTOB2jp2jJufZWIpJBsZiNnIba7GlZibrfVwUx1U
X+XIzeQ8Iff3qV18fY0HslNI0FP4AQi5H41VBQTFAoMZmWt4NG8nkG2Lw8xqWQ83
F8+gjjD8eaQJTVBT/LjzfUpJ5n1d6Ei9iinrYmLI68aWT3ImmjLd7vskwed8Mvy1
fAEzXAV5hpRQNriIT1YPqgwM781AVerHv22wY+UjB9baRdVIxpNxBtmhkPNwTlQ1
dnIWOPythwh3o/iGbOOQO9fCECI9+22AnKgW1Qu34gvtU7wh64k/tB5YNqh0RBKD
KORwuLeqr7Or7D4BKNdla8a7WaSnD2tbQn9x8nSKkTt8qnv0kYQZqFwSWHRuGfdk
4JXgXCG5Z7bxlDQ58dA2vtLKTzRXM7jOIVfP6KqxsmdSFm4bQx2wvxQQfFBNVmXy
hOmXWKJ0gY5xqlo5ZaX4vqwFO2GD0Qoq7WFdvUXxQLwmXahPGdbq4pLIqyho+KDE
c4c+GMNXZb3TDWj3ppYjPlp8kh1sVObyc6d8Gux5MdkztukVLMTCEgdgplRbMqZE
6YwLDN6+XZjCszxTSOvO+LRjB3OqKwDzlWUpSYc/AwHLmwTRdPnBCtaOCk8/QVrT
akqOnPpG+z0woyM3wBA7P+6irutQX9HXgB4obX5AKALqpWMEP0AxAbCgB5qteL/8
Wh/Y//XvQ6TfQPWt8JN9qLUoqinzLwWS3fh/s/xfaLq1e+PcoX1NDoFBoMR6k8EY
idCBxhkpceyYyzd/msGi0kQ76Zc3+VNoymiTDxbJH2Cok7coYD6X6NOGLcoJKxCe
KBhU6+R79wEea2TlUeFGVHFWVfreokO5B6YYFvUD2PYX9n9OkVo8gRlk3yxLKWNf
XRCCI/6EEpMggDo2Cyuj/N/IjNhBHzx15XHzHZKELIzCGcIzT3pCvs7SHx9Bd1Yx
/N0ZlautloKQGigIbs7INImMs89IKDEONs1CLW0TpEh5uphqwSKkS39ZduCpIf6W
6/fMbpKrEkJhwk6sHfO8bNhp2gIZ6osuXBTetehgM8OLoLqnSie2oXge548+PNfw
/B/LAumjF5mzWKR8aQPE4wBdOiiJ1zjmTuYHgXyrF9fUSxi/wgqsq4H9vIOfWfZY
CKP1H0TuobQi89NnAy7GpiaBO26+Okd2K2P1ZBPSL88CKh8ATSf1Ob9atFzzKqrM
bhwG8ac9LAPvOOs/CSWz8YExfWC8SsoVzkBNidrQTgH/ySN+O4kYLmF2iKlsMmPv
Qj7DOhb2Cgg7jjTHQVpHtDSANuPn/xW2Vl7UQReIet7RXV1rc80FtseUBtGGcnJ9
LtppuoND+x3KkOB2qTHvaXeT+ijwl7lasqQrRkDIzAw7bVJ3oczh2jJbM7FB+wfx
m0mJUo4h/kb3jw4pLaM9ryd5Za9V4t+Gfg00TJ3Gd8rYsyOJhwxNG+U/F/7aNvjm
ZQXD+UZ6UAS+Y0+agN8kJZT8wfGbVklfelP/JYZniviMcUyKdKp6qsbGpLz5GiUh
Wd+YNva5tCU33Xuf9zsh6bQPs++65gFeQiXWI7hhOrfDo8Bp1JEBWAlWPxxtjZa6
/xHLb5LAXIBgajbFNBzQJ9i+h3lQFaHX0NgFeT829CvgXrv71lC4zLQVm4IEgzrU
mTV+GKprGoWDb8iMTe32FV8Hyxc2rc3WOheh/eVqpP5JPKYJCCl6rPbSKATKWDFd
d//qrpMXqw3hmmIJd1o+w/Z2i3J1xq3ncKk2qLRjCT3+c+/B8DkotvkZ81HC9xKi
+7V8PBdoFnEzqpFKMAZ6wIvj7XzbtkYu0P+PhEJs1aZeOdSv9pEMpmH/R7V79DNg
JyP/IooRANchN7cvPWjTkQHIZP2UYZy9FWzysuM82RrrHUjAvaVY3Yv6ZGVLGl/A
XVbu9sxFIhtJUVUVxic7bI3CNAVv+TVIxImGwDBhO4cepe+jq1BWy1gPt7aFW0a1
Z7WiQ3YEQ9XXOKpu4ixtnDiyvI7873TIVhtdP41bW9g9IlfNdFlfXP0tNea+Fj9o
vLRVYxJAU6lYl1nmb1En/0r86++MTIo7YFC6K5v04vuyJUa+ZbGOltS+mhFfsgaA
MFTC+dIVfsy0IpoXx9kdiorF/SX8+2+jbDWubBKRR7F6PmSiltKg20Pbicymarvn
FkZz9nUNdG1IvNihG26Sl25BDQ06DRXziz7tzu0/hLVcOQH8R68909BjI6VNaqsa
G2icTKyUrtSKmuzysmGstHq6wl7WGhVX8MBOdRWcijDzJ6hoRfWI4wF/ZWroAIf6
OwWUjYP8YdPRfN4g6L6BvW63F1VJfR2U1r2UGsjCZlKItOygedIKCrdBrn2H1OPk
6hdW1tkb2DvbKj/tW6sYfVF47iX00MkUDqSPx9PnI2BgfqqSoYdaJ0eZINx0GQ/I
lK6r7Kiq1SyPhNUU2YfgIueMLkCSAWYJVaCptrcUuEWyxhln8QlIxPJR0LxByk+Y
BZ0vstnY+CnrKbbohmcz1iwECqZOgQ0x/0yblIlr/3EuMBqZh2xWd1YFY2+MmtX4
Tn5WqnYUcqprn9Yz9is9HbksF5oVrYcAvmFQ3BxHwTgGRNPiaPPZdM3ejXAMNN6A
9kDYZ27oSHPmydWsFZdVi+NZLk7l73NuJif+TD9tgTUY+2kH/ZE1x3tgLnTeFK82
AvseJoA79iJpYO5KRedP1YyLO5AZCveyxoxhIYk00NpVORuIkSaBfCU3sebEVGIp
0PhoL6wdLqyM6wCrSwpnVxtBsTqdX8uHQUrfrLt+awr3E4MxDmZWyyXRcRRThCUQ
u0/uBQ9T3dF/lTaIBVWAz36YSAoTMuLj8wC6Oe3tZVhG3C5HDvT9XUK1uYxoIETR
sJegLLbCaJrXQ5SjzSPxqyvYVR9CE4x7RUy6hqEMIT2QGiK6fBTFX4/G4o7FweCB
HRMgCKF4RYgT2XeUhiV04+CjCr60Mhq5WCrSKFfmK3H5znE7fxFb/Aizb7PJhAaG
B/exPyYZ9+EVgdoOxfTZj2VRxU7nKkS5p1AsPXHTRCpP+bqoLXjXOTRyuQuPwGE5
VBsq+kxQ9hAepxBEqN5ipPDYzT2wM5gTFnRnKCe87NxhxpW9ZW/QjAczClqnVTyw
BhRdAPe+U06frN4vvRiVLnYb+5ui6Qs1RQPnx54Dmyr8SG65KlOELUCzkHELqawn
tH64RcQwcP49AzbA490D2fpQYyG4dXO4+Y6MbNwR0GY6Gz1kGtbJryKPbQb8dMBR
MP/Qj5zLATWUrl+DCRnVlRDqXHcrkjvNb40D5nPfRBKvOpAnMyApF1kzsgglxt1m
iqmHhiSgL9f8Dkt5B+pq2UcRcO+iAUEsLZE39VowivAzxRz2CGEelop6i9Y1f0Zo
5In6P5Zki/o1BEXs2YEba4IvP/EA8eWZdQkYOeyETaQJhWlxfiIS2AjiT70bJlzy
XEapy1f8p3rr3oVaqLS1noac628zZyZL5eXIlGIhq4SFoc3odcqqfshBJXX+hRjR
CVrcdx9aQhUzOycAxsGYOgsd5F77CctO0pnabk1anJZGDU5BIsp0JxWBk/gso6l0
nIor6BE7dsnDGYEndjt5WvnhXgxR69Er+UTomegS6p8Jm5lWoxMwCnxo0jrjv99z
cc2Jo2iUk2Qmfu13vsdYSefSsy1MJXPpTNJHSIXUZWdpYeouGXcLQU3HvC8GPFCh
FCX5UCFhoFP49pD4w/QVxUSOyua/di7GeeLoMfS9rrKCrAq6IyNx+X2ygbycDsqH
TXrmGoEqiaxF7xMCmjJyFp1ngx899zkjT/PCwwxGvkP19wL03OHyIUgva6wqxWjx
gw1nEwyxQePUzq5I3gpIPeoyii4xrjUtcVBAaon4TX8dGiGIPpcZyxEitcOfInem
J2D2Sor10Ryo7Jh6U2MY6vk9+Yiz8Th/5DAFiCZ3E4cANZSy1voldWGc+u1pUE0d
GrPVXYyG/rsTWLGDGCZGCTgdhVYlMGTZkorxrV3T1bACnXpTW55hdMXBpNLnu5LM
lFSY6hy3BUYZiXuxV0DI5NGs+TuJ2cy8c7tPvRoKJ1TCnJ+yI7kUOx9sTsX7NV8X
DoaIb/Do+0QgqHEe7dKQj7GvUSAwJ+6wGB/+KNjIo6i0BwZMhPFYRh552pIkKDrJ
OvI0dpxzb2X3tEWR7iR1NKZ5esR+zWkMsfAReksIY9+draByeGuLNmGPuFqboc95
UC3O9hbUG8ss8jMJExyABmyxKJWNUL18hvTvhNOtoQ1tqjH7II2CZ5XVjYrsa2Ex
worMyGZQtiMg6YIA+DkVWhzP1tIHxDU9asV0L/LTbtgpotVVg4sk0cABeAXovcvM
HUjJBqQGtm3YHG5ejFpgTGJa5RIgVVmQfSmEMQoXgOmFeMwWI2T8PEw8X06qhWI2
qkalNaNO5VjnS2/PvxHn/SrrS1hmGkVZaeX0QGJBt5iZUil7d9BzbobSX/CrKxxt
Eep/9+pSRGGLJ6ERhHUzcJP8LceAeWcOfHSlwUQiUflByoZcRHsJSAoSEEismmPx
diSi4yUodZH6p5r4iHHDkF3AdSlUfXY/qGPfjb4uQX+zKLwwJNUh1+iSkQKZbwcP
+r918makUBFrAcSUPeu3oiECk6W+k0AEZEYeRVtTbss7uVL0onex/zqTeMsvIwRj
0M4Ol4But/ayZGfXeoY9oIDndfyL9H84j8z8wiooq5KV+jttWtC7dtoDQxFyg4Iy
JuJsr570WRklj2fc1h6u8kd8nATDAZbCVE6AsLfHjwCF0nmk5egGuY6vtZ8LoefW
YfSIckLs2YEnvmqVZ9zE2DLOAJh/zGyz2pCrEZvT2I14guBvsABpUFd0e56xsnIn
uNOo6OdvXNQQJdr/q4KleM2sclhaG3++e0k9lWWbrvOA7kopXf4v0u90gpJxjw+j
nuRzUsxPlp6P/EyBQVGXJ4CPu81ZizSUpe60D5FXhZpIzpKh3T3uIkIh/XzUqno0
fCc2XWTFpAaZ2AGsVaIPf7hHNMq/NeHod59MYz88PJiSSEzDLZTCLPPdh1tbVEGx
hUAVNl++QceVMQs0UIlGwoK6NokhY33eVe7GFMLDPJV2uAvqC5OowFtA9lQLS8PB
xeZLve1G87dVUfs1Ia98Mn6tL0sC0CQkYCDUXubrTrmqHQwPPMgMmRvvG+tI7Ixm
lyXLX80Z2Oy/P/xzefOtmYai6mNG2eGZfV1Sn6VrekXwtbsKdCjRwmEYLA1UDKfd
54WXiSgBkJMoAJYH6UjcBuwNutCbfnZTQIcA9w9yrDjDBH/ZAiV5NQfIizla9ci5
jVgb7+6yXoCuGB684JlRVbVq1L2t3AUaVrlDaaJtUTgbPBhXPeivFlsTxOjZD0N8
s2ppEaQtV1E9iEgfwZBSumEj9NR95papiNstT0q1iim7yfmkZBoB9ZvPUkftbLp6
3p0LzrES4v4Nesu852nUEAkDhYzhJSQV6KIcE4t1MyLahOYe8JzSkUHAUAMSjdzC
1DC+7fdj1oSKVo0oHH+oKM+ysKkHj326n61AXjaTnntL/y6ktxgKISiR4VI1XD6x
HIHrdtSOdcTjtOvcxEnwcEJmY8/80O2rpmU1GM5KH1Rfs8/QLsakSQh3byhfpK6Z
8zFgXBT0B5z6TUOJhhYK0bsPDIBqM42eaC9Cr07UoxdENRE1zfoWpnb11BEys2eG
QMma5Mu3YzbJI9dpCpshGcrTrQRctjiZjZ2ey4PjcS3bDMavZ2sUmR6WMBNLhrAu
lGT04I5LfYfuGX3aeixJe6VyCZ+lBQHilFWEOeekDBIldqgQfkUY5MHKT1tufxZS
5xSm0GEter8R45ERn6tiu4/lQSE4+rxVtES1czm6DSDE6Q2p9f5yQqPN2IayAPnb
VTEgHaXwuFK8gj4o0wDEVUtDsjPu2u9biapM77tJH/C2KAo/HYsOMA1xk/RhruAT
Radv7OOJ5olhH33uoCHxHi5unVYqUDEFdYTAvSenU9YdRggGTUlAPb6lBo2fxSSk
GOB4C8MdABkvmYTaT99XFFdsPZbi1EI2LWwmGO0FPI7gbiEz+6nKoXzgd/Lkeows
8nhqdgmGYkhQFDDK8w0D8/b87bZkpnVOJntILbwsGH36Nj/reweGevs0ConEpyO8
9h0xLmtfy5Yh9365QB0GOpyWiHI9DG+nLRCbuQpvUHCSuTypUNhU3LJq/qO3VSm5
2neg42ggacExg4BCXED/GM6FB09w0bnNm19w28KZvaJ/CpmCsOjgOGQZpMlLbnPH
/hRWDPNwFEINGptCCMBn/rgBqLI/L9tABgyJ26XuET1QPw05NRCo/3bQar8wcIFR
NjtQbMTkH+pUu3HlwQaLp/IIqZcTD6PlafpUhweOYK4uIjYLC0D5r5BtUb/omC+M
ZwLCcT0OVse+n5X2pgqtT2tG/GcBlpWMb7XjCWi2MyVb0X0ImGKm4hcWev3HCmqn
az8X9saNYNed6HQ0S6NsqZE/p8mF7wJj4H/hQLkMqEqWB0LxPHlNhYyCR4iwagcd
l7rwZY4/0708RNolerIHp22vUfuTAz85wpKU4rT3gHX7grhh2H6pXVvmhvucGbEF
yTZJaYmEraIzdSYtUJUEXLvM0l1Llvj2zH8g2qPX5/0xiuPAIbTGKBb7/gz3rOlf
Z91JhnUUtKNUzBVb8mV9tGBNnGa9LhbpUbpqM8GSWjbCFT0bYxN1zkLkZFHXoZXv
kA0DnRLhiTOovnrKTnojUwNZCLc6AiEgDAou/Nqu/JqA4m+Wt1OPTykvJdBGJUAG
8NJBxCIOzpZWm+c14sHm5cuCdKg5FrOwnBa+oTyCh88UdOdl8b062T3mARnqzdX0
7ndbjZDSD7671DPFm5BFFN+AwO05TiS4GDYHw18W9kSCcQr2+WgZH0EqKBOB1Cng
eiRbrNHsimVyKjlqYkQ5orDWLlLUXd+cR0T/O+EKbqnSHS2qjSI5mxKWdNWnBcj4
jOMcFuqntIW6H2NlB+4XKQBcjua7kLaL5rw0lZXKA2rGejJI0nY5GG78ZHojgerv
mUGuejLcQ2cqDq1KlAOQ7K2eb5jjujNW/nXki4y83UOJyBv371i9gaRKo8FNk8cR
ir5mfSo+N7ne2o8Gw5aF909xDjCw86e24x078xLcFLUHF5oysJ+yozPkq3iVjDzd
q8jkmmeEf+u8OLr9h5mLucVc+S9u93le1whugX9E3M/NaU2a+4lkUfoMS/U0MFGz
AoRDk7etlILjdlLssIcTTgS4QO/PgAp0WLREK7bFTbgY5LrllufTg/sn6JAq2xWK
f86v5O14dMKEnrbDME3/E5XyXVW4ZJmAPfZBxRB/sMECDj1ZofY5eUo8pTdrZrrb
Y3XSN0xGd1koBnAVrQNGBaI8n/cNFsK9nr2xdSZgQBkJ6xHqBUTPOAz8ayuDmpR/
DBCRJN7t4p2OuDDN3YrMGO3yBU+3NXMNG1xXsip8IhOIn3h0nWMoy2Ce7RNQ+act
kCqPs6x8PTcTGYRdHOe7E5u74J5lFf7rzn2+AvHe6aP3VmcCPl12aq31eA4g+Gy1
0t/Ngyf0M/o03Ov07DBEZ1c9/RX6HNiONBkx3vyHV0+fcGJJMW3Xqy7mc4Dmbj14
1UY/AjfkjuP34XQoDjVQ+J7cLb1BukPcvJmjJI1JrsTWXorSOoUTsaAh6mCf/18X
37W30Y7yOn6MUUKTBg0YxlB4I1QjA7myceWrnGkZje9RpNMIMhvyG/B2WUrCD0UA
W8BlszZMr7aNM41hU3Enc8Bcw18k/AuPecwm31KhyzQf11wodYSut/gPdAcaFgv1
DFsS8jHlJkdd9mPEp7RX8N6+XhiA+tYpVT/LXM8R8/ONgdMb3LFA+JwU50167C3b
J7SXqbkCmi/Wzgbud+VN+9zPDrQv4QB+BRvB4aMIvqQ16VBR467CrzPkqXOIXSXK
TbEdcdJvPDchfFiEgZ4yoNktCMFyOLRHyUyyv3mGOU616V/KhCdYWtONjxkq6rUp
pM4Wj/pyDALVd5eMntrD1zMHbas0KpZ8NRk/EaM6u5S38gGTn4+Y4sITcpHGcQw6
fHYwfPwrZG1jxc7vbrvY6hpPhLAVDCm5l2uGWUto6w7sMBHpkQi6Muo91gU4P8hp
XDCZO2Q0XtgbgDdwZC0yFCCddCNt/UyP4EEv52DbB36YJlAcFSJup60rLXxoaz/8
0lIDAdR4kusCGoyxhXhF46xp6xCzRp01JvB1EwA1ZFm8AGQy4grHQQulClqU1CWg
TKvQFloS23lQ/dS7V9didf5prhE6D4N6i/tDLn+5iV6Z3wd2JlePI3KxgAbRZWBz
eGayFUqqxm/TYGWxWjnN/zYF9pAxZL9uG2eIU7+dNcLLG+9qhIMmKMLVZ0chw+C/
bfYCpc83jmM+cje5YKItg77nB/7OxMKKYkJo0UcTYZ7sWrl5rINJG9vYFja2KYyf
+U2xoPJA+dfpD+wOPlPc3ZRvMKqvIgnVBdjmrAZ5IIgHJU8pHxqczhp2nVSMVwQQ
ngq6+XSQG/WeBbuNYPOPZ2E4qPWcGDkQFTMugbuT8EZxAr249DPeG3mvuYgP2JBt
Gb8wBsBqccUsawDPzb6YZbEzyjkXpOqh2JhFbRAWfhG+aUfrMfhw4kxMucEDo4L/
NX8d3ugcJ6ezKTz9g4D21T/MbTX6jUsTY1BTBC/XOIXwR++bwuH4JA7COD7xQBbB
o/4vFlo6x6S8CNA2IRH833Bc+UPeP/JtR8T+7lktwy3w6kkegxd2PUFB6Xh5EElZ
N6W1e6eaVC/gsGyYiZF6IpN+L3vLWH+a/UdXXnA/t6iUWDkz3ILblJpCPE5UJd1t
Icj4IjZ2Q0pqb8aEiTHoa+mWHhfcD5aZc8eiyKg3OalTR2Uzj4OMNEtjpTuks/eu
Bb2nORlSLSVJumYZWepqFXfSaVHcEZir+Wn5/cnsAGQdtiSCnh4Le3zdwqCVx7I+
HIEw4AX1rfQ5js3cuVJ2w5cycs662qlCfh0KphAzRHxey01WwnahzinluZuVtBIb
dQTZ/ORlj80XQVieHqPiEO7zw+vsqhAp/R5XXEEIwSii0WSLqEmaRZgDnAaVr1en
vlYBL4ur5QdCz0LdVNmxvr0cGw5tmBzfk53ztXpGGOVfANyQEPQwa+zXLpD4wMfr
NgQiKFPFOdbyFWFfFSZOVDtivTI7jdHB2ksRkGJ3a2OHfT40573UVV9s0MfyLYP8
CSqjnU2VbM12dVD9fF+U8oxfu92tu079flAhPLEFDe04CK1+q9MZJx8f/SF8iRQt
rqnvqr2B2mSInlnH9Ue32yfPaEUAwVSqHvPevI9ikLYtxnXPg/5hMnkr4i/A+41n
b8SNWWx3RJG/OzT5tXAx5SMmnoVEklqV8gaOLzEY0JGE/n7+LfaaAwfGIC0Mtat/
3SJvlEKMLNU6NCFYwpy6iu0wJWfKt9A6Brtyy+2tTpDvETnkEDJKjFEUPARYVIS/
QJ1tpU51N0f1rCrAu0SjBveLFYdcMRlJz/3g3fQjFfwZBlUVYnb3k1Krfc2TQPQ9
SplgrUiCOTrEx9CNGMV4U5Tv+kHhhMogPOtbZ+sJhe8ZT9nFYd+aesUKe5/VFua5
T/4AVfIQyaFct/iVdxavr4E8IRghavBio0l6vGC8ZjSn6eFsT+xLPWMl/rXtk1ps
TvlKFHferYsvXhsTY9ZMYPvzjf3qfY72pXh6wuqLMJ0HjEOCD4BmqiUxMii7l4/z
yQVhKIqYAwJXwTuCwzH5lFx12Bo3SJS7tWriP1Zo+Q515ypfQDAR6hafC6CRIOIQ
XykGKthQkVUxTQOMd2oaWi7GlMGP2dhQUSrkr0zYLvVHy4s5AxwPUrTRebPwfQAu
YmkACUkiw/SpLJRO/XQJrIuq/z24cPVLqAQiABcj9xyOsTjEiopSdjwiY9bZXmUB
id5uI732qAIxgriPINXYurGYN28IYBCFIVYQqySzVxuEFoTIdgb6TsGZW9McjVhT
cAOlU6nhv9DXFfVpauiVJFfYmV1RzFVkUg46WkF5Wes6gQRHtP/kctGZAP86OI7n
F30LJQlYL2Spxx4zUTVFHoTpODIZhfvK2ZSkvpCGBS+1ibp7x7ixZhYiuSvcij49
IQpGgNoCNB9tOqMNnG+UabpTrehEXay/zpZLyKrDR7NNOmcsTbP7YfE45yIGSuCT
K4/H2oot3EFm979Dgu/e6C7TnIeMqG/ZAd0HyS4SjVWlswTAWsZ5qZkNKtiWf8+D
pdbiwfjNlwREa+ZvV/gCoQ4HAo8pX+8pK+VyhLZMKkxQq2lVTr3oUg27lZarwI0h
Rinzn2deNtovA2uCEWACSM9o3R8E5Mgzqi+jxLiSBG6LOZTh4Xnpxg5hmKIlO9MH
vzs4645lScfYm0CvRii9dHA8AKP03Ns5JLXPoE+mBAEzGqPf2jJ/RAO/hCNMjYHX
lVPUNJDrVA/TkF19LP6UOivgXg9rUn/Ns8mJdW089+T+o69kceDzPC45B9FWtaoQ
US0NC4PzQqo/uOrT61/FG/C2FoOB03TcOwrlpDv5DTznyuoulbyF3j9qRoTUYtc/
Gii7cToKCNOqg9zxUTQe/z2aOb7wYcjQCzQvGA3gFCMSHe8oZlHMDKrYBbI6cBgv
7f5XdGKXPMCVaTgrbRX88sGFCGCTyI7KRhlPp+KzoQy6a51Q3AtXKAIrIqQltSyZ
J7HXNKNI1oKup2mDkluk9QY4LSvSzSiFVtPJrJVKmHRJkt9vF2jcct4ChITNsATE
pCJng+nQiIKcKjAXicsqUnVmZqmz/znhqTI6UU/FxZN5guttcDr+aBLaN5EQq+Yj
Cgq+gsmZi2J4mQqAAZLMwLAz/FZ4CCGZ6E9P43Ehzviumh+KRtzdTCTwEyzU1Psm
gfJf9uhOURe25Q5zUcCctm3gR7dNztgY0nvD4sipmwWmh8+uEvDMy3gbDxuD+FkV
4MESxjGqZappmLz92/YTUbQ21RRqXa4xdMGgTiFHTZjo8viuYaubRRoJ+NlHso0A
07auH2Hn1xP8pCTQ/oCGXIRYJazvBFGyrYvhaZkpvQlygy/uWDZCATPdJtsX3r82
4UCb6wWxcypXqEf0FNJYXLGaRwJ6Y76u8GloVhM8hjcdjynoPMCVy461eGzR47mc
KeRITJHY6ejt4gaPAROonoolgt0TVM37tRpzHqIpWwKZYAQdQWquc0KrKzAxA6Wx
YIPHnwA0vERwBdIIA/YtX7bF41em+72F37OW1Z+zwwszuERnQEZS6AnIgEQXOKCA
/ceS6iL6h9U3t2n3TkC4MCB5n6Td3OQFsavK5cPpUg56RZAZBAALLTVSFML5LelL
yJflSlERMo/J95Tv4L42qKoHO9/J+AtyAza2HnPpQAoFrbnIM7SYSjheocVFIyuX
6cRNv8wP1lLam2uZdlx0pGU4WLakupR2QNf6nqERmHXvktVWIKt0mMiWm4Wfjvsh
HU7//TUojFYbo82ruP1478lOKckTWisOZ1WWsJ9VV2UGQ6isFHs17pNI3MgAlDX4
fH/BOwO4UB4pnMZjiyIpX9s1gtlujLlS2nXWo0iX8ghjOByFjvrqBsW3wfvLMHKz
JElJDXG6DALcRNVWA7aKhW/nncsMx1GrOUwWifEzpx2lstGR2HtKeO+5tS+98F3W
SSMx9Qeb9GLWJkD495XXdjUjM6Jilnxx+nosokeIQKgY+S3K57GH5vUtwUH7myJ3
tYi/eyoz7BC7i+shQmYhzgqQfFu3woaNfeQzV3G+ZjkLPFlvj9LZW3CkiaI57gZ7
LTfcnvLdUbhuHe/fPgHLxAV5uyxtXvto5pcTtIFMEzqk6bpjQ82Y0a090XN3KPJ6
RuUe1vyh0h5eQgdhbzjp+hl22jmYe19TGpKIbFsy9I2vRkIooc8WVP3zP1qEDGkD
MmCPCbR2KepdW6CgPeFHesx1jeW19Ch+NLfcZ7xNpzDGJJmbyWQu7ER4KupED/L9
s1tceyBHoR5BIjBi6Naac5a8pl9qxNRw62yR1pPN/znvRa4jVy/DGhActCohyTHo
/L/U8vdxK7XogzusVGgDYaOwsLKzVoH9Xt+t50D/TDCRxH78PiWjtpH2rQ0D15tC
+OubNwsLtZmaD1FOzmswFgdc1szIqhuzo4Nf66H9Sc2lEV/ZayRCitVmmP7LduBc
coe5gmJuNHQEXss/aEk4aynHsMpLWegYwfONxklwhf8+fUD5wh2g4ipr1J4LPxdz
gv4+jJoF6JXSSjn6o79e0CSK26o0O1pYkzSBWkismP9JDzBWr9M1TbK76fjEiCkf
p4dR20LvJ05gyjESW8kgpkctti94JyKuhqe5n0NWgweWNXVO/AHchGh29lRS7GAf
CFzIhynTosjIKpXCHAHSr+Z1Svky9t1ohFlv7AZIQBatrpULItN+x0X6BpopQPHL
jL/y7uur+JMdIo+yBg2NWNdIpKiBBIkJ6QKavjujs0X0HT0gy8Q97B3u1aAAirKZ
Qw6N4OVjI/4ilECDXfUW2io3wi+QkWeiIV6GcmwywFXIVdqyNYzfQjMeJTQSSoKT
WS5qHETYZOO0HolYSrRGbOZ/vdCBMXXuJeeMmm8VN0TPE0HM+CW7Ort0UAeDns45
Coh0+JQTBNkoQ77mLBVdXMpx9Z+vs02snPEL/7LwTN2/cgjUh7IS2rgbvgFFHZIZ
bi3q2SVPTjI5hSfxlKWx2bNrBh2BXWA/W5ASmaqlrL0aRkHcdjM4wwniUkpr1UdX
L4V05mJxTXNaI6+efVLPb6ME2NCb+FDuc4KUDt4yglnhhL6uBDNVDGtFyZ+I+dMs
E0YV2v5BThJNXUkgWK/gC6GoFoaJ0/wH7K4mysLADmBsnSMovO+dAaXmqt/3F4iK
UXoB2cKjTbOiUk4kW3mcIBIuarCSALYsy8Gme0w3AHuHEtPclC5kRAySWFheWBbE
NHfoIUESUmNkKXdNXbg0neCJ1fKCgpOV6eQLaUcHJSln4MGab/IbBdQwYpvmwRoO
wms40EEHeyYmBRbFIAPtxaG5lOOekGGH6FQqf7wWkGiQFDTSaXatb5jJKmSwzdci
HRLaiqNJ1zfrsIRnsmr9EJkA96YXY7DAi6M5APChvgvtVPoAo5WUiKEjN7Yrn901
w248Ir0mj1T2erS4nCybtSgEF+q7eMgWfxau1HLjux92iOcdzYii961My/svY98W
q7d23JWdVKSYkbFdxckIvOEY0wwsDLSLBeAjnfVBs4vw/hABEh6zh6fYJoNqfOC3
P3SrzdAM6TrTm3x5bCLjjUb8VVIz290hjKjo+oXQtMsJRX1ME6rFiLB98Mn8telC
svz5ISGzWW1Vz870AOfu38aswc62fMElZ44oFnRm7Kbz2jvldzNg0523xlvjsdfc
H8EWhIYrjYQPR+3j/gjfpge1igvtnb7zxYbfnvQbLeiZpbrEWRxl1OaXrdyDfMYW
pqNQUJxpFkacRQ2846bk/L8w5gVR4zqA2YnSurYF0f7aujpN2PMt6Ipy/MnfX+15
1qY2ZjB9wT8N3SuhGbSqxQ38ovvamUPkXfx1i7sODFlwMO9AXYcKd/Hg+WaCUSK2
gSob9coMgtIPBE5ZRK/gy4z48k33++pQ1AxHlmy8AqL4IRnS0gCqFKcSOgzR/+2E
y8VENCtL0N/DdjHYmkre8YYsxQoG7H+UXb6rNk8/2qw6coWAHCm91m49zARAumzU
TaWd2a8scbzfgInAQlY6p9DgX4rLJtHeW9Qw5izd+0Bma3FAwoSJWdKULffesGZn
lh7gspz/oIKUv0Ii9iFPJ+dxlmRcpWL6+DbgeM2HPyGWK1nQMLMQ4usJHkrsE9l1
8nrah6jQHMI5c5oF0v+hULQdAzy+ByOJuZAUgKn22kq2LzFZBlE2PRv5hhnsR4uk
9L9Zuo+Tj4U2clHIR+8HRktc2REMpWLTT4DjhppzDjF+8XFRXonWhcRTpvE50MxJ
B2L+kQknw420F0QWPaJriWLI3pl0GnKJpgA5CjjMLQ7vEX7O7KihX5QjlpPmvODl
K0vmRU2w9GrpXNFK8H1hrr7vanJ+hJImCPk4unGOUSjZ/FkifEJxf9aab0qWUl76
ihfHZkB+Ba8YqO75NPDqybLbQh97SBhm0telX4rHRoxs5jYyNQhJanY/ZnMvytRo
Kky5FFoJPN2sXJ+RtCkVm4lxlwyoBFzs0QA7KkmNdaFpisGPZBL8a77hwrdd4XQ0
1YhnWv67zKj7u6277dPqtPrt4JA5yf/8pxwqE294OP8KqodR0OghpH8uvaEAbk/7
TOQwiMLQ77tjwdkH6MY7OroD8FPbiSDy9rOiEW76+8OdQCgjYm5Wuh3Sx9v1wAUG
dnMotLP71xtAR3G7Uwk2v09E6HPJiPcDNCtK7eDhYkrToU3XNhOvatBDJtfZJt/K
D4HW1PKjA9hQRm/6DrwX12k9LPyHlkUZAOZ3cocQxq8X9vrtbqzykYo9+XAGV7zu
B3ueu8zoOflvIUvPHsKDGatC+J21WiFyhbgfIqvh0Gpi2cEJioaEfnOBSry/Vf8m
fmIn7rQHu2uhztjz85LPtXcu1vBR6+sjbvJmjF+Zq0dfj1KCA03jmr2TySpHyr0z
NZm0Gt3RzHxueZheJefYAjU6kpLeHRXQQXtTtJ9cua9yzyWIKd8cgM1s8LCEzQtE
oE1m7gAc4JSrSormWlPDZ0/taZ0g75yhXOSU/gWaQuj0fGOPwtFIVYx1PjqEPott
ZVhMkXi/LNPl1ZYSBduBKzYJBdq6UtlAi6U4eXqHdXD+G7EPOxQoGulvRmD5zN0+
K2rgJ/F6s9ZsTn8rvOG4xoKJp12jg2u9+j7SupQI2T/c5OQ4+zP91ke+Q8zZLS1K
UaQk6xB2IRTg2lFXepWjRqMd5q0omTs1DOGUPJ5LqZIzX7dYdF7Cj6HCNPq960PE
D3c2ty1fEMtmweTtImNr7OeFgpw/CnNyd0AARHwgRbKsd+MF/8hYZTF2tzrEeOT0
Am74Fm6/vAPJApkGQhzxqLHGEpgqdPopjlXuCB+lTu9Uef5tbDbHZpN0wnFzCwBx
TNKtM3ZBEIlUBSbDRQx0vJEYFQLxa8maf53YhL2s4yJgPeqGR//G7nP1L73Ax2G/
vrmSJYJa8xA+SxP9yM0PSfypil7lEHMpHgCRYsq8cibBxqDCb1BoV6iBeIJYRFdr
mRE8V4M1hzjHkKbWCPa56AOyFeoQZrQcLU0FqgpMWdvWxiWdsj56NxD27zLl4qNt
AWN4dIENCTbhJRiyVzBTu14LcolhP07w6zDGSXqFV1xYJ6HdGZeG9YU28zWNZlM8
R2/k3hgiQys090VvoNNkELzGF1yU2eaU2hQ5h1Jyzfy6J0tTUIVkG1LL1N8iJ0yg
HELk2G/M93/mNXCyMyyKtPnb8QO0F3mBXsN1p+5kPShMaj2orCRqZRw7WdzPua7S
BQ+oexY+LuaTQFNyXkZYQG1uCVIJ2Q/xZ6lm/KGXskpyLV5goR8elg4HHmJdwzOx
U+9u4omqdAJzy6YHq5q5zX+P6rv9SxzqKQ1rqVCg3G3BQSmmLi4O/BUqjC+inp/L
IC+jXSPmxiKhKHu0vzoZ1TiggrOeURsaU4ypc3jca9ZqtyvEsYke03tmfDqB5Pbh
QMjmjolz8xzE48nWCmb5ahiOyQfPeG+L8PtsOwyHcm3SNz1AHWYsaHqlSrdvO3hi
QtD36DjgTiw7rwVgHA6ce1J2/xnAn8lMldmefFB9/0hD/wb+qOZxMpkZOvlSV8WH
mFEI0gxE1vY9/Ij9ijDkp12MFd52ke15p8tCoc0XtrpOXa5T9C+8w7GT4wWYnWuh
dXHGM7aoCHCdC08eM2UQaArvhOE2rZpiKt//QrpowiHe7ODvXJbuWOemoMFT+GNd
Rlihy/zMrM7+Ukaj/EiGskyl56bIjCdTIli9rmsSZ2X3jC+mIj4RXiZCyXBtiE0d
L0rL3de/nNDbtaNycEpkYy8MQ0e75TDbVolqflpBIaAV1MfHYILbeVNncfGpE2ec
PT1LwVXr+uvtgZvM+Hw3HrYbif5J9h0jWDgU1/cFSCuVRLYQn/hEKRdKY7g+G942
ER349vivzCSmjaRj9rvytQVoAy4Kp63YHFx1zgZ04A7lq/flprJXGES4td6bQn9p
V/Ay7ZzVs4YlF34J9oNk+oyEabsY7nuzxlPjmhvjEYK7PGNGDIdY/cCdpyYeTRcQ
GEME6v3vnfq0rNhSfXsom69xRAJcN87gzFmI9RQaHJyXFQNUqSIf1wtooWgucnme
2kx2U2TjftZ87NGITVkG9SyYmD3g3Tho1rjWJ7n1f6Hp2OFB1fh0nfxgszltw3YR
MQ3CvurOf3qnjhKnyHq5Dnlnlok7FK6q6xDkN8L/npQSq66Jrtml7NdCFv8vBH0W
+j9EiRhz0BcRF5OWT3GIwXzaIt+XGOMsM2LdyEQ/MSYx9/gKqklms4xUvPPWBQWR
WMEsImzsxmrB+ePIgwCeOBxwZZUJxbPWLRruEpWtj9ythGTOnHhk1KyF8S/M3sOc
4xbDdpJwV1P/tin1Tby2wBpHrbTSBnSneYoh3X/kaBSsCavKvw05mE2fykIR+w5i
kc/PLrFh2jOIFTay6GTAGwr2MNcNYP105EJ8u/IRBIbzzP0g1grK1lA7Vhqspmt2
haU8b8avXTTCMpIZ8Wi7eKoY7ZqUH3844x9Hg3mocSRsXmVEyjrK8Kl7vi/Fimrr
DdbXXwxVGacxcJ7EYq9m408SAj9pZ16MwlMqzqspQN6nZPfQewkinO0jO/ouT2Tj
q/p2fJiI416gVdqQ1h0VppnqPtzYDrS59Ld7OLktcBffkkgAYbx4L3rHvpBl+2XY
dojSAvv6LMHCTKIEkBmvFaVXsGp1MMSz0nNEhi/rnDRqDs7wejc3nLUfM5CcofHM
8Q4s7ZabCF5vI0dcarlyXfdhmPHLZuaNkEebtEYQdZSYfv9Bd1MyBpbXWMZ4hO+6
BybFw3fzsEwrc9g4Sz1yUkhRXGgaB5L5C/JGxwFTjb6yUzShTsbleF3VnhWQ67bT
3lmGb4Ypq6+jnkxzQHk59Xq2eVyW5N7Frr0GTvEw9d2ZXBEHIZf1t3o1A8CWivZx
nMf24yXWwSNZxDLazzu4v0FEXxvItc0z3uYrVa121+b9GqMUhF168fwQZaSC8PG4
ToIQZk9fLx+Fn7nVMMDN0TCBiARtNdatY1lTHJiVP7iBGZjY72fXPQrA7o0WjxMB
w+XRDxV6SimeTMuxKoufx3tpwqEeY7lx2wlnJeOjpSoYqg0b0yuEeKXkbBYI9GtO
oOYCNiTUkGEkjcXHK1nJYqt4k30HqAaHXHoig2zDEeFE5yGUoKKFT4b3kTO4/r4A
3M51ksdWiSubikUe6JfsYLBz1IeW9903mWNrEMkVZXU0yQJQZ5YGGCHLy02RPiN7
8k3f6Vi803M3Q8I68ErjADeH0WpYy1aSFL9s3py8lg+KmkIXzmCttyB6r5WjVLn/
Y5dYRXr+FgTbk6XlGAg8S11DM9TPy/kC1LVQGIFpy7IvTVE2LDfLx95sNREcPBma
3BvBJ7pw9hI1i6LebWHfdHzJLGuvAnV3W02kk8HV05M2WHF2Hi05rkcD6sjNOzjF
4Nz+7NjmXc7uNhRS2D7sAocXz5e5V+F/WNZ4xl62glMY8jx4aBHkAuTz9wq9LuHj
Rzrc91Yxq8P9ycqKkutcR3+JtxYdxBCnZgntaPS7HwbsR0RuMBDkWsLXbtjeZ0TH
0EdRNfywXpmhRZYUCqMgq0FLGbyBHJ3ykUgKjFdw96RNUb3ot/lwLmzXHz2lDz4d
oah7T3dGhpNY2NpE6gZnAsry5ZfP/hmATEokHLHCYHScWTX3RV+p0VtmT/O2slQt
sudRm5qCNZSAjXDpX9aiqXGDcUWu00zbOITg+95xoIQGcCbT/OrpuxVuLDp+GchW
vtO7CYBaahdm67XWkaSIkejN5BZqVIOe8r0CvokpVVtfI8FxhHJe+lJVbquCEFvi
vk9ZfpWQNzgScBkEKGboVpaDJUfNUuHPr1Tse5DFRPn725zDYzp3i1w3Ian20Nk5
m/Ap23hf0Kk3jB8cLZEPLKHtxPdJsZw2FRrwpSgtD4WqGoxJsOMGYR2vku1obAfk
M0INRmTqONEbK2PYf7Yv9P8o1n0cXqnVc3fpZ0NrKnL9eFYCEh9uxRr2uxTD70la
v2aEXxfP72dD4vpe2RVcxgwnAEdBaLnw7V9P6/M+qu3tzk4dKjrLWYQRYgT1Zvu+
U+E9SWXxf/HXhGPP9arZ4/uAJ550aM/Yrb4ApmNYZVA0PwDSP8+yjHgrTn60m3bl
NBEBWWgu2OjXUCeWv+tBFLhjPYTAAlm6YVEXScKLsiL8xlySeLKqkNq+jWaFn/2q
TXhSYrPXo9SpB+z2sPR29HoLvIbpEc1+RBTOYVGQKY/1ukLdNr8ylQQqghFfrvYA
FangBUox+M8ZctcVmeRJjvye6CCHJ9BAQ3mlX22xV8QVeeLZtcO1BU1E6DfJ1emF
6OD+ZJoOsbvQw9/SEzeM1N5NAJxuJeLRrJTjyZxHCL2U1MLrrTRuv3zyqDnEi8Z1
tassp99/pEVcetTYdIk0VnQuodh8lsclcKn/oClUqCMMP5do6K0xKadjPolTn5wv
x3vlY10IMUESJZdqNJ59+bJYDXzr2i1pURAaXJzAYQUP+A9Hmz64bEvUDZt1rxZa
LGjWCgi0vp1KB9QnjRW+g+rFVIQ20DzmiIVt8uetrZhgKQm50r8FHctf8YhjIz+W
qJCZUyg+R8x4xEeNpDA91DR2vCr35eSzrbn5G48ggt+f0wWx/2K57FSWKxCB5LYK
ON8gBsCGl64OJ6oozMmH6/Q8z+pXux0NTtQ5fVnD4zBp4d/Dejq1RRnKbS8DHUrW
n5SRZRlNntTkIBQbc/bk7f6vAWGNmCVn/tWOok4QBp3SR8wPSmb48FJGqM3EU61j
TyAtKeLFPA+7TfUezMi8IbedZLsgDhpoQBG2Zf92hCjI5+WqBLKNpGVJhdXYrwo/
YylsnxUdSljPkEVnH9/Eg7q+gNNL2++RGqzn6/y+dnwU2+VtcTiLvZqODIdIGXQP
AnQko7yutTX27VUN28LwdL0d2s9+O9m6CEYOsBhi1/VxxCwpAOAqnJ5DA1VfQzsD
Olhz9YwGPcOxFyy+O4MstbeiWJsJ1wsJAfGsBTY6aEV8xEuGQRLKJ/wzUF9K8XLA
B7JrKFdSAgyOOGovHM7k6RupaCxW3xn8CMmBzasWz/sLb8qU+OpE8H1Q+QeAn5an
WS7x0Z/dP4Vp75rxrMJMFgYGVYbNLBNYcCc2s+nZLP9MP76sDazux4ZB3iX3ZjFv
ItXIy8AJQLn/tJPWnfApcOxA6b6VizKGHxj/OOoeM16FPZKCYm3pE3W2d7PQoxkL
33vEjVspNn+7rB99Xs7epLbxnPtQ1HNAP421/bqAJNhwR3r6QB2Jh54W/+A+Man+
TKoIxsI/y6EsUKKpPbsjcL63xTiqSspbQw/MZRMfXPbqotVCgJ3ku+2sw1hOGnn5
4Au7iYp6q5VyIJITXqE9W3tb91shWnx0rIwC2Ixf86zhUOLkuE4Lxwftvz9+GVuw
YE+X97MfGs6J3ScI6utIGTs43YiH/CTjaedTZwvj2eGE0PQ0sRIM6rEW+mwWODPJ
qlt5zBKqe7UphEy/YI0AaawUvQzaynkM/qg4Y2q9s5DbwUcu1DcBgZmrYgaJU2OT
Tx8q9udvSRo69KmftQU6hGUv6x1Gg7C8HRfRWMziXVfpfXy2GbWfX34j5nMuDwcH
YlmMNRAhA9UrI5Vz5ukuBNnKND7UKgMQIbFXWxcce9bHs597Tbanmuw2iadUPacv
eUvPhqsv+HEjawp9zZi3wmNo9EdfLd/NqNF3gNappGuIdQLD0slijjOugYhu/Uk5
wBOOpUJ96NNrp9QcHMzxPDqCOw3o7K+b10gnVHBfa6y0BZuORPr8Zdcdmw8pXPAA
l3lDvw/haJM/sXqN1hcbK1cfkhEVx490Tr1aMfJ+RxMWbp8wE109950lYxZGVXFt
RmWDX4YKPcle96W+j4vExU2752YS57l/n1z+vdmp9Xt50lz7ItewBd9Bs91X5BCs
cgLZGfUHO0WdaT+uKRE5XcC3rwDtKGBJuMmqlGfVQyMjxc5I7H/5+7Pra50xiMrf
/xxO1Qx7JSnEW8Xhm3SSoOCiMUm0E9a90B47UDlACJXUs05tSdM4AMpUSLD1Paob
mhqWBCCWT3LcIFTLV0nlXZOItnghIJ+oMj+KgJcGb5IYsx/qKYMJ1Z0k271JH41+
4986StidaAf6UXnYdcOonE+uJJ9DD+oMoWn58KRTQ2F10PocufZLWtNHKqWpuCtg
36hezh4DC+OdfVjJq/TusFLB05XRz+ttPB1WIywoeGO29O/N1nyU7l4id48eoMu3
al8FrwClH1Hhlf4qTCgPFuQEV8374ht8FZAMTPorjb6Jcr8hERjoC5GTcpOSuPvE
XaeUSHD7QL8Pg4THOmi2XimCMOlG0tdEE0IOz9V0Zh50TfJ8dA6+3VM9kwNNVMUo
7NBmFfLoDEQtZGTx9zb5q62Y48GsUcHOGw1dqNvCl92LrCxbT77UfCqP/6DI6CcZ
GJY6po+Q8HGXXywi411QxKG0A+uydRdBjuAbUkrnD/B8GHAr3JQC/6kbojywjz9T
kYgsv7b3DkqGMQqArLRREjqj9jNFoK0M5VRN3wghLpXcMeWbp0ueMRYM2vQko1ON
Pn2G1bU/MairZGi+pEW5VkwunOSkNFblSEsHyx9Mwv2qTtSLVvk2laWZww/XsoD9
tIZQtf1QzJ2Tn/hEdr55MUroJZKik+MInce4nOozgrzaIuPpNYtv5oquUkTREE1F
zTq+y6ovuSI47gRoW8iY7zrznjuSmNLPKWpIHqsA0RZjc61o6FQ8LdMqpdvZM88M
c2AWK/3Vxvew6iEBEs0c2bG7HLIxYj63D1egI+vUndoM6y1p1aTsq3E8vB6xeapI
lHhOt76CieaQKnQEvF0ANOpUgJQoI5Ndr3tEirvfZUWtgaRI3ZGlhv8XOKKntGuB
dy0r/saP4TaUPpVNcDjO6nOET8ZZurvgT4MxaQvmrM0x1Dr8y/Z67ZaDXVWxz76l
/auvM7n3rTae9VTCHQMzKXUmTTXd94K9SzyT/Ve8iMEiOP7AruynFh5JgdAyOdLU
PUvoBDQR3WyPm/p2ONpu4O18RRIlWpevL2oPgau2MfWF0BGDAEgN5n8HHVttI46L
40ZVvLKKpxVmwueI6+PypD//6UvlqfqbNegNXUr6w1yWZc22LnckDD7DlSwnxghc
9eG3tdLwRjvOC3edSOc3Z2XZpS5tz1nk3kkkg2yCV7CbmK5X8PDF+vpwQeBhjcr6
hs7oJSWaLYcKtHbXpui5dMiQjB4kpeL6eOYVyzwgbXK5th6deQcNPlG3NZRaTEqb
BsTdEd2eV+IkKvvYk7Y4ZOVCHeBWcaGeRMwVSmU82IorUZ/usAFOZPZ4ACbKQiZ3
j4Xx/f54ghebhYMoaNvLyIuNM48kBz7OnVBcr17yaxEpGoBCF/Rz6K5EOFZJQR21
LqF/ymppBfNOwiL//4tqyxRTBKm5mB9G5Hj7t6Rg2OT3WNsLXCLiWpyfoZ0Jmtvu
ZTTgnp5HEYmmLdb3jvr+lUCpv551WgYwMjulGY2SPOZDJ4+YCYYzUnHEp8n+qXvg
OWv0/2r2p2LlG0sSdxP7zwSPlXP7DVijVnocU0fqqhvgOyI5EGR9Num8+ykErk2I
yKiAra5NMr7pHFHogMupd+xwYnr/flkvbUaXVzgbvpQQiIF/eBqoDT9zukvAdjLi
ETXU4vwogAJbxAG1trpRihrgqRXY5pV4wxQgvV9PukOzIHPVgT9LB8VlupIL7po4
vmybHrF+/KOYxkj1Dp0eMmKLnrNMPY6EsKFSI0kBry5fCVmVPBNYhUqtuEwMlprQ
NSdt9qzY1zK2h36W4zIy6kHibjwNX8e3d+dW+J/28V8Hz1N9aLBEUNupjNoH/5vU
gaQ/4UAz2Vcv4cab+unddtJHr3c+CVucoUyzqNJVK4lUOgF8CPayUNXEVh+uBCpd
neog+rLeMRs5knxuGX/zZKdJoWXHDBAAXawowxL2X7yxY0Uta/JGUhikJhvniDhM
Mu1/aDd2pF+SxvRZbhD4OySDbFwSc7gVxRjdoEMOt+VhjTGjjVd+1x77hfvVxmGB
gJjMzMY16bWuX2Jb/ODft2utNicYrv2yLRGxsE9mVxctChbIWQ1vU1ArZCeQ/ojd
D5BaTsc2eE7bumC0PnhsDmvdky+pmIaqyrDCGwTh8D6dwCHO3iQnFXtLLA5izAtR
x6cV4XX5NMRj9eSutuoUHyRBCT3z6mM4b56E1NagbfI3N8f7ganKXLtsTqu+2/Gt
6p9zjoLQ7Vt+BB8dyAd9GrbBn9M9cd6g8BzooGD6FChtviQ9DHl2YzhRF6xoNpZC
AKt2laSdgnbdQpBV9KquikSR4zJ2+DWMr/efIeZdf9WMLer9ddqm5POiVnBF+2Ra
FGKNODedLvA4ve9Ne5PymqQtonXRWl+U3n3ggJGeUee7UE+LhZLMfnvU2W8juuTO
Q/ZFXOxDUx/zh5xLS5Dcr8tScVJTRetwFXu6ZyCZPqlv+bMRA0gZCvkdE1neGVrl
EUhwFzlxK5qHd5zmk2j4z6Y6K9RySoSYIz4soPhFjRpgoUPdGulocRDmPWhIt/Sy
zTSJI8nSGAineddxSvdIVrLSjVX5W0SFitCAeMhCY7mggMcxoVMxmwEr4ZOzQ3nQ
oa7GFTcp8J44Uty1GqTPbRqH15rh3861XR8TLUhWjdBzRZMa71r/EtxayM7OFiU4
viOVNTHsB0UslEgRxKZoZokb4jP2VMwY9hmXLu3FbmnO2Wo5jT62kyfrVQUEuN9t
g5O30K1O+WdouaA9ziNVbDh+3pkcuTDNlpLm1rMT1zHWqGjkNSf6MlyoOGvGSwHN
ekgt26P5UiNxCwMlbcIjl6U8g+hmDS8SNsuWu1iZsFWzZS5Py4HIizgCR/vqDVQb
Md63b0X6dVG8BsS3/WrZPfFQBCe2lW2t6szwxcMTkCqPxjupDqCwA9cX2G0LymrE
bO3n/grj6Fjf8Yy3XiwkR9yXoa3AzaDULuyTv+/cdTYVmIUhL7THFCDKNlesoudA
U8S0qcN6nJ50dNOK6JXzUjnuvM+9WvmkFp5WA9vdlvRx6HjgG4OSehecaYApa+hb
IyWSAwIxdNGKc44KwnWyazo1LFx28b9iAnmUOyAlF7f1k6cmPuzDcnUfgCHbwtpr
YWA++BtagHZOCfuj5LnjPO5PgR4XZKqHXvxqzD5hN05juGbzifFZ6BiqtL1EXTz/
Y704TUwBu/E1SOYX9/NKbhkmAIWQrq7c1wW6pWGr5gM1lze+YlfhGhcv6gzhlVXO
D3Xl6We/5sLYPfWg6llYw84ZrbujySg0HQnsuLei0NhUhluyFRuM5ilH4tSY/4A/
2PO6C749GsezHSf9EM8DImllCLTDds8anH+EL9AVMMep2zSLLuReMKlU4yh8MUyT
VsahBZcDoOWuUOWOTPT6vcyRdAvvmGsFJo0VLgSm9U8lXoDySJUPBeZbWDppYAtq
32BBO4fIdzLkd7F2/W63lk2Kqruy7VhSMIn1Z4bqcuXQxe9y1/vjPKr6sjtijenZ
16YqdadbuWYR9G56YyOtGbClTrLZeJb6xPZNYbxYHNz5exfcoKrOjxtYFgcrHeQU
TbcyWSHSub0KPL6OzZBt4v2ac3lOtVGMTgDsfaWhsknMa1NKqbJkBOczLyCF0sNw
CvsEgIz6UblmRxYZ72c5m7Mgc2L3JL1vnlBzBvL3rGtsxg0sSuZWXxH9D4P/79se
Waim0MZkSfj6xyS99brR3ARfueUw3Z+0YScMcoYWilkgWK7MVDTAbjEvsz5IHUro
yM8+Ep6ovkIuHqsYPfxQ9fKNuPYFFZ9ebnGl8qFUiRkOUPbmv/vebDAOKGoT8vGi
1txkbba/nRBorLDiGY7r2lmlnRgmJYGlDrhyBv0SHvL0K9eLdp1VHlFo/t4dF/DC
QRaWaYpBBUQ8KHJWgyoN9T+fz3uLP9A3eiPriLgOwtz45JpUex6OF0G8+d/9lii/
j1MHYCSiia0oN0gK2n+mZOFZgEGfhcJbePzirkKIoPkU7al1oT2mNUjsDDiVn9Lj
xRqcrZHne215YEHQvvexBbHe/4LbTUjRulC7vwqSvdEMWdpuZ52bP5YRqx7q0r1I
dckRtoxt1M4EYPC9eONI3kuTT9Esw4ir5ZH1swYpDRmCektDso0SNIPOXO8rZ+1N
JtRK0k72reQGZQS7Ylsncr02CpR9qsdWFDzUwRFo+IR+5WvrdbVzBFOW0dCHtftJ
mYEMlcUW8q4zOeKgRHGm+QaeE9/163QbutNLxgMBEclnfPJRPAh1jbSA3F7epGw2
X2PcW0bg9XidDvPAybE8dxGFKDcuSEgl2eVQcO6K0Us85Wbhh4S/W8oV9F6pVeb9
u1effNPvRIs386ZSDi33xG3hLt6ezNgLIXgYBIp1vQoVv0Vh+dVva6gN6ioaO2NR
b2YCE0r3tH1JfKnMXTsf2TTGKkeEH1iynziklKrVLLhQjhEb8I/DMSsB88Lj7WT+
vv0PjxRystBy+UZYYauRXJRzzZZpN+HLIFq1aXy1vF5dSBQLygavvWUoZenH5Ssn
PuszqV7FKi8tNAhw8r+DUicWfLLC1/PAUvSGwa3twhrZTxz9pbxMY5WuhUmsV36K
OUk7F1KCmCQe25WazH/kfvuRDl85TZhjfsITIeWj9vTgCqmvF5weZcwLRxbksm1h
cGM7OHrsdQjrGC50vr5cfCNbFjst7wLYxcwZkIGFvGOrbzQDBg6Oo4p/wR2gSMB9
YGnmzUhuS2PgxNc3u9NP8vQvU27LQXKp1MjVt79mNYa7pNAtNwLwlggI2LMIudjM
9/FTCri73y4T8QNy+/zfWbyoQ+cEw/zHc5hRU1EoCzQwjLWMzQWlUk6cgHJJN1hd
pOSy2cF8I0mthGXpMIukKcruhLAO+V32RFHFbPuGwaa0BBhmZ8RhyyGRt5/yv37k
RG0Gp6Ryl5PQV2LlXN1vhsU7FR/5O60sL6ApIG/wMppjS2zOagDJxYB7URMLGZyD
7VTFZ4q8ANlZzyxYcVFTt/XzWx3TwJYQlcU1jk6A7fXC2DxbU9Ja9jFsaCO8q3a3
cmZJh/BFw2heO/yh4zQcd4fmeHOsSSjdbHOqj+z77QZIKPG+PmSzQ30OhfCvsuyO
Q4ffZmGAA/iAkpJB7W9NzyA9lI923LASXTlV4IhgJL43IwIm0TsTJ898NAReeZ+r
mthVa/QF3+TTCMNHCnKcE9/EvMcMg/+nbNqJ74sSGa9xhXmXN0garhWv9HPN/YqM
bn57gLw4WLD3L8oQ14aszUHTeM/nQlmuwbDlwTMIdgAnnCTyz1h/69gkfWGx7mK+
ewngNNKrH9Ddo1t6ttLH9ikmE9ibXiqO6dJAD8EWIJ1g3o4ReQyQJTIqoQZTeYqq
w+n8U+SxjdV0EN59d3m51muMBWSo55Wii9CfEGJcZ1fim/dQebOwhoUzg7ihqKQ1
jTs1Dv6q87o1Pxgg8elUoLWRwEZmuzFFC7OgsAM90ElFGvSDYaK+3NeOLnpe4Dx6
6z6YX8xocpzLfXByu/agwcp3bhSqZUEASDGNCMu00AO3V7YtMR+qSLURAWDFSHml
mmz8gjcfbOeh6vI3fUJDZQpNnn/3aPldzI0QeJfKnxwiYYX6zRO+ITNTHErvemkg
vS1ELL0U/BVoSKuhNFA4znR1fmNReOQv2l7HgQfgVKQ2n7vTBv9F8EJwJNnA+wIn
xAYaA5sZiW2+3yNitQG3XQqIhy3V2l71RUOtIuP/fuCeC1E+ZQsmClBLfaSQHNS1
58X//TPDzhpikfVbLwSpYWwSCkMVw2N4FRokq2n8UMRCsT/ttyzxlzY1xEQ5ImS/
E5/hA4AOdOjcq6QjMg8WZPCpYWmwNu1u1TAd5vxgAtapCZ/rTUdHns2f+ukg2BLE
ipXmWS7VZNqqO13CBnjyRaUdRRdx+dAO2nhnA/uY4g38W13T5SQZS2idBIuKiHtF
7dW0r53J5KOOM0tuFI+uVFF2Fpa1GKePlYl0RFczoT/7BvwX7lexrmEkrii7zTyr
2Jsjv6hP9kCTIIpFfUNAAwEkTJcoLvYbyP4SqdDuaWqO3o9M6cqp0TFuO1zPax0z
4GOFOYPEsXH3OVFlkk3m5dTYUPHQcZNhOMcdJr1ZbR2t0Ut8w/1ayishEMYXvRxo
QX3Z7uAu6B2rXxJm6wbpXaFPopDexsJZkdUGuIdwZNGfbrf85KiCFi42AUdH/YWa
8dFO7upKSec2qk4YuomfpKEgkowu2Pmww2pQBiU2mv1gScZ374piTwfrl4pnUuhJ
WxEFSvwQZ3f+edTkCGckmgH2zkThPLtk2XlB7aQ9MGgze/86qig26XP1dG2Ebq+9
CQ7QTP2iNuhQpGl+TDuSlEm5vrrXdwnHOX8kCzSu9U4Sdi+1DByjUlzisqgk1R7o
zwtn6y6XKAJloCI7+Z0D5lkVfbEB3WM00nrExqSGqmUItOPk5H0shfxGU+yBz2iC
7U7erECsW1x0EDXDFvldXCbY2yhDWH8a2YHGrKKOJ+PS+nC3vRKXnoK7yuQnfqxN
VlpoSzg8o2zsNg90TKNjdN+k9WRyBhSo1trW04KMF0878+qGl7VvZYF/E8C1o/rL
ToiCCuXujf3tiC/EsJioBQSwWoKqBnEisVdCxyp4Y//ZDzExZhly7P+e1xqtWRRr
9WbQ08NrvqNxi8SY6IwV6MphnvuEGZ6+402d1YAfstrnWloUAV9dGC8cInqXZkn/
BQnpwVxuhba0wjqOrXBvZG8Aj8Sl0vLwbXjdAA1JTKoCrApTKScSkys1Fk1sALCE
PTddemr/pZv3XSAPc1n82FkW+upidf+nWQMmWWuZBeYBDMyAtWaKoYBzKOm01btr
NgbbOH5dfAixKRU+wvv93SR8U6K0fCAcu+jbjZ5nu7UnARVqbwQqxn/njeIYRBXG
2f5I3ZmCrR2BzrH+fR2lbJxdn/cwpY7AlpLlcCiwcxL/xmJRhhNdVAXHrrA1Fah4
pqhTX9yEDGVBL3+/2H/gn/2EC5EdcSo2cHtppI9p8fS3lcqXI4ZK/xgaJCWtw/uq
zu6egTqZA5AWIeeBk56qmvICjHagYPguhwvPdC0cKF0J+fehRNTHkIwY2waOGO4p
M/N7YWqfET3cXQ2pDkW/ypi49uaGVh06eR+gGVbd7a8AzbCgz93eI0rNCy2uDDz/
AZ+Cy+IViB1kd/5+RgxhZgwgx4/5yTfbgUgW3suZYcPB+1v+Tr0D0lrAZyR9i2fH
LeZcAWKkCEYbrFQyWX+e9d/jXU3hAtsVPEvNBPRCZNpoqLhrACgXkESR1gLjlRQg
eSa1CZA+IS2m9u4lyvs+HTUAi9uft1A7gjt14fEG2gY21STjBBkhHrEfBpFY57sT
wFgeqOtHk/fyN9MRQrg5WbsNAZc36gw8LU0AS/kfY+3fEp8nnaId/JUqF6vADpoF
JVJhi3hI6D3otz7InItjBEInQyVi8n83dxsvv6+xgNaNCz50iN8xuKnCYWVEubjM
Mu8v10nffljpvjEWyAmG9i8sJd4hEIFUoE+w9EQgk61+uLXdvWNHsX5cnq6qQmon
fSWKE0QkuIXsYQksmzLY8LZAUN0oAk0pqRvWg7vXGYBxOVztKbiGu8ja5VGyuzeN
ub4eSKYS6DFE0lEhICbS9WiFNdA41ekgKgX5lPtwxFSQ9IHO18HY3+rQcHFTpAue
gn2TNEYXQTGhos/3ZeifaFCvqEdZ8zK8q4CPT0Xo9t1p6BhNZWBF9B8oTMb7tRDj
pfMdYE4xiO//vKDr3QLmiBYPVsWKoLp9EA7x+a2OjleGBLuR8+FwHQRkU7i89q5E
bO2GOGQcJLdn5GOXkYyUoA3EZa3y3fvbB8RGCSgnd3AQXv4xgrHO62vbcKM3/3Je
cVevTrkNuiE6lHnzzoQTewGNXXe8Nfk/7kpurxGEwicfnkln26nYD7WX3p6mFze8
A2aImweYHiIVUqOovdiG7Qok6UqIRycjzcNOaE22FQZl8Wa+W1kzlIlrUgS+5h2I
tAcVZKupzxkZGx7IOzeJ6RW028HukLi86bmiBUgdXPKSuXYGSACldRPqb7igUfQX
Kmq60eIO/YWwdPAHxQdHzglp6k3MXmUur0wTnL3efXfUm+9IhFsmFikgsgGZ8mZb
lrae2g0trunlWIxVdW+tObjxHLuX9mG6YdkGVJvoguXAIhvzXRvWG9FYc7sofB9n
porRWGMtdNkC8NyjS/gTSC3OQf+zQuakOCKZoFdySPJ5afy3Zst6iDZTaIveSi3u
C1Ij6CjSqm6DcW6i0ubvaLByhGe5EH4zcgh9JvLtQT/wB+t8ZZA9/W8PnF4ZTvvJ
GzRk5ZCYeq0fACm6JLwXO/Z66wGFLRCyUx7i04LISclbLcJzfotC5cj5grMjOdYz
948l2cYanjSlcRt9TUbb5mIK8A7c5uDf41+T/2Si7cL2FH3VkPJTUb5c3gTrxWjU
csj1gOCgALzcqkM48eg7/JoO3BjczRf9kH5hX8sSQgyA7DuWaDQxjohEeAGnt53X
FTtYbmV0uLJ7XYKEib7JyqB1YuVrcIJaUhTXru7EjgWeYTIWmMcrz8iPxhwedPak
fBvL2EHo/PPhwBJrqer//MaJpQLN2p07bZO4CbK7PkFZOOB9QfFihx+GXzFR8qoh
iUfNelZomeLAZkpb+0Hp9hkNazqSrbOEi8XiWFIU0HEL7lcW6PBV2M90N9kf+4/c
y5f/cQdQmSz8z0mtyFHXT9kMgCfm5SjgALFHEqOL3VwNjBhX6JWKcApBVF+fPmRH
YJQMwqI7KUIbfVluo9lJZcOQPQdWZbNItAR6vqh16y05FlYt03ucCPg/GggWiHdu
fcNIoXDgoNxWOjGKsn4wMWEFUPQd04YIiNLrzdMOlYa2E+xXZFn0wLSlWIDxrRh4
XUNzhA+yu7807nbdxdjsIWv9ogA/mCQhe5zMb1lk0cHyquB+9WMpEs6opy+DRFCS
EyKTADOhXC38GOivSKENlNWKvOiJURinUjhEgx5T0XeQCm257o0mz/bnxLY82S6C
LLZMrMc7265V6O+LTKauo7Oq+XRr1NyKCefczCeDmaxa0PCZn2cI7JBz4vVm5sv5
e/fpRPoGmv83ed8wCgwZc9gB4XFqxtT9A7716cSDvUswEMnMgTQQev1Az8IggH4b
yre3kWf1TgZHNO2Ppd9V+4xm6w/oSGgQzOvLXsB/i0NShUfKVDrZybRs/bW1DfQk
SbuPyGmTziNjPZS2nV82GVWsyrInVusUjqXYctVDlETbNn2PZZi9SrTUlhJWSDtP
qJFfDonTtw6qdFLH4KimTZMr04fZhUPdnWqEXUuDhktrNx0njNOo6Q0BNARgDEeS
XXGwa0Cx11xjz4ES/a9rdhGwW6Z9bBc4AsQUlac0KwffOgB0ABnkXWisjczXnrAT
r5bSuGn38LR4JQTAl1d7TE6thkI6Pp++BT3nZT0ZPUZXx6SITY6xdpKaaInhgiOy
TU7f/AA+JjKO6HRxaugC3o3SLR2PmcvAMtztRDUtclZRauDu+AU0nSJSbmQ1EJoK
OAwUeAwjW/n2yzyl7qUA8CzAxR9UUcXwQKH1uySTgRFwfNF+3NrP/ItdFhbRkc83
UtkIyJwsmiWXHHZu56gCL3OT/f5bBX0emZ8JAO1C1h6v5gMVlG9bN8NixEWom+9I
otAl880XdID4W1XfUN8eCVwWwskBm8ToP41llq4CmHD30RSN5e0rTVzDjz/iGEAy
Oz62WFcqH3koUvSVKcMoGcAJ9cQAnvSyHwVz41wrKolUsN5zb/QTNT4iNC+iyNj0
jjMYBDJve8e9f/5Gtyq4gzdr4raFduo7sGJA2qO9+3yJF6GeLvNpddDC0B2w1ukJ
9Y3OTkmYvRWtIqp19uhsBzTX3n76l9JH6UCKf38tGeO5x32cGaez/loZDDibUHHk
iv5q1xjYkYB9uQHuSEwBhgFWTm1w5YWkW9c0d7LAb2M0rZk0x/zMmuj9gPuISzmy
C2D6vreBm15knwe9HLlYh2DEEtoh57cG7HYLWhr3aSCTT3pUgtobFCd+b+gvtsw9
MMDcDGgRY7j6ph3/qqL1h8kKJFmVsTRfloGFvWQ691KwMbss1fRQ3zWIBulwQB/l
B0PCjFFHNuDzZT3aA6VUINdHC/2ILPQBRciDOJ4Rfafn0qzmnXDFq3C6wJWrrzXn
QO2+1dFtzzHJmMDB5zozhmvWYj2UgEAmOLAip0ULUlIHX9cT/fZUuwB9lKUBpCLq
gUR2uN+iVzNNyT1mTbpVfdnDgRDWbW2svv0kmK4DlMVeiikqtq9A9OBbRrUfDAB7
hJmc0W/KwqhMie4N3l1Hvk9hJojPbLH2G6FxLYJej1Q8li2sME+ss45OiL1zk+3r
gXT1TULOwSRcPRBHbphZE2fsA4hehUj+aWQt7JRZeU42AMOz8OhArEe/JS5OD9I+
X4kvoN1BcjJfNNRNazP7xpTIhyDOn+OpRXfJrrGzdtZeuFUgHij0IPRaBrVcCVNh
iHDW9U8VZxRailSVBGBJVKTLAyMgtC241jl8106SBsUozhhDCzOHbeXk+1OFdFMg
rEB8ix703Il0uWwg67NYJ0igHEiL7aRPBSkLAfAnl9sYn+IvEQ6Mp90v8MBZN8Rs
9eOcUH8v/uKmBKAx7MbZwXib2aD82IG/yTl52KzsC2XQyhAZrUOJgsJ09WihiZVM
qZtjt8rYZh0WrtEXEvy0t1dlbRWEHtzvUolIqOAlXXQSz4r59pa3FmvT8DuOm85g
E/qvRdEBAtQkUJur9Jo4rTHRljkr8AQLEAjn6cPNRaTWTDPfDZivpq1oPyN4oxkw
EzgbA26u7S25doYG6ZoV7qtOhBfzSExaVqvlxksJYXcf+SLXqIAQWuWFM/Z+X0G8
VLxIx4I3bEpgnkdxSUrucw6tGdRvQOZ93x8EmP4hDHHqatbvQAvZ8RoY0UxBhfDl
dWoNnQC/F1pZGLJXu2P+VofUf8VwfC64Ih0tPW/0GIX6p/IIQ3G1ctF+YZQqgiju
ieuRdZfwWWpWGrTH4fw82OUBDRPi/3h5Lm5gtQYpBoVQzPFXHlo2o3x6lEa3u9XX
YxE4ngxZHa09XUmzPlYqEv9vmFPmqEJ+njt+PFs+hzm+ZMiWLg8gc/2jq2uMWjYE
6d0hGcV37YIfpSZg5sJlU+VRflobFBar5/KKaaWrtA9kBnMs8SaoxOQ2LCsPGJ+m
jMNw9Wdk5DKp9IhprxAeZ7SCC1MNVhEsnuHdLfgyl67PRVpN4ICb44WWwFsgRIxp
BvdM01b1W6lsI3i0IMStDCUjX5GA0Vj2gdNZ1nsnfG+DyJC/7pZirPTwuUM78VRB
+/kerUqXq2Ggaye1kIffLOG/qMCgv+v/NJmkWdQekE4w0H6wbvRrue6z86KYREt7
SYgDG1yhxfe/3fjW3DAszB2FsX/yK90Uu2Lmm1ZFi4oxZ61QhOZ58uz2aent31/i
MVrK54rlttn0oCjyXKWR2GYsQIHNG9MRqBCE/1sTGRQAhn2F3VDK5raC5FhIZrM+
q0NXq9Xw9RdwSnIcAxI2K7Jz0PUoi+DRTQWSnOI4BOYG4s5LL/BXODfg8H5PDB1/
pS5eUxF9i+FzUvj1F7ir3DT91CEaGVUM8ku4SCPdj9IM/PAPYCkmBhmMly3xMaTA
F7aTKyHTzMTv3eSoEIf9wpAp6+GXQvsL850J5PPddThziZU9gDfUhl/HLAijtIzW
IQLlBz4NUGtMEiJuvHfLvuI/qSz33K49rX34rkg5WAdiPOw7YaJsuTemYyonPw5j
jVBRILEKOprrPENsGgBbStprJl3CIXf0v05VRMoDHh6DNahdt8udxKiYsjLr82Q7
hmzFAtc8mvbRZDUBeHOq13o7wYWDoKbgt99glchgDopbleXOg7DdnnL0diDqJsg9
6is+zHLk3u13Ou7Kn3aK0zVgJlRxsQHuR0SYa8O8WSEUc5kQxXu8rc+v1PIvGL6O
30QEgHuHhZYgXs2knbMz3ghirDyvGKriXkvSyUerghqCDXWuraaJVl0mKDZLZoc4
UHkFl3O3Bj20a6CaG6SR+04lGMsceEJGo8bCI2xVoTPxmTqDYhEXpQAOfEDQ/YRH
LPHkjQ2ADKKILnKXG7l2pEfrhml8Ak68AiiM2Z+QwSv5VA04ZoF7fVtFAOjJd1p3
cquj4Z1aCF4gj1W3AfG9bN35yAde/iZoZEEbEh2uZQ7/HEhuRNgftUU1402YSrT4
swGFv5RTh5m85GHsKFESkd0nzi7Mm5PWyxphhQLSXLgUwmHYiVp6n3POdBn51vxw
bCO/YTWjOGvQPUPJTzCbFqJmftoT/kgWhtYdYY4+gPJYXUFp0EwhcjU2/xw8uXQZ
0+DXdW9EDWsyNnee08x+ogdarkeGM38brYh89cfl3MVonehPIN1ncU2vfItjZcGB
6vxyXcKst6HKuxmWP5F/uKc+fo89RAppw4f2JroCVYltbWoJTbzAgIVPYTo84k4n
2u6lOrNbq8P8jDqXA9x8Mk/ZGD5JPdtlCPT8byofwAGGMhHSFkYkDLOyoLlBQlQq
wQ0hqw7OPMpP3BDHM/2K9c+wBMm3z2J2IkRllefXvN8vZMNif5Ym8Rx6H2XBHfZB
90ZKjN9Blp5Tkxw7mvAtXSLdZEIblkZ3NfHD7Y5Fg3wsT7hw1k7NvX1SylrwWkoO
lEktBGCxcm1JqhmLBSzJurZGLxos0eeXU6J+uh1D/IvJpf3Mw2N9b9GAsjPcM2B4
/r0evbD1qo3/FUrzpg7jU9IiSsOiyqvokfcLpUMw1GwIXXAu6/t78y+L+MrZZ+Cp
MzwVuVMTzrLbHqkvAGxvRus9VKiHj2ud+VWClk0ts8IBETDHdOYi4UFZffccIVaU
jH65PPhYXvXna5CCugnGWfvOG/eS5rVQgZs40K4HI2b32m73Lg0dH75wE9seobv7
g/T06nhP3cz71KVXvFvNj7/j1EwJRS8nqmhDKAKwfQwUjdbwRL7qXQOTfb6iNEdb
6NPgnz1+nmwQcpYrB8GqljlMD5rR5CrxmOJ68oXugxpTWba5XcMwm3HoH8iJuw84
wXThFxMhPasNIfmvvlFFG0cD22eWADSmJHd+hTw+tvKWHk09i6oUmHa7WrI2LXNY
fQCPwQP8a6lXOMUJHl4zww9p7iqsa9Sd+xfNXCEkn0szs9vRD5tGZ2jL5VXzrbPX
AR4ljpU5ypQVCToj9/Y9foEzSd2pzG7pTm1PZIpNmkQpYZypftokwX9iAKUpL/kd
/EdwYrfVUou7SFzp3fb3Qzk+ycXcfdtak4CbJfUpHf1Vfxo6E9Il9ttjUvaKqf4m
9PMiME8fneUukcMK72F6V15U+nF25me/3ucfJhE1cOCisJ97lA8eebSapPW/WL0k
RlPM/R/hzQPh6gz0apckULMBUSqgCZBCtQR5gtbZskgZlKSa91LqmcPcem121fAu
KYkGEEN/7nMcpLjXWcRvAx8d5spBvxiE1agPZA0/WOKvUGz5tUerdBJ33+yOPr0v
haR6p7OVNySziYc9tpfYr7byFS4sSG2d1pHrVtUF+4DWBenS/rm728PLrO1PbdNs
M35JDhMRFXs8WfcKZOZK7+YqDZ8fym3nqVHs5x6brMZxnWU2An3e1yOBTk+igwVs
Yiuw5H7Rb+sF6ORhMqP/bEQJNlD1ajZI+Z9bA+7NIOKHqV1nztEWmdsg75MSLw6K
TP7ci0g4z3ny7CbKSft/et2pulpbwiORxgudHIFetYW9q0OYl5eX2Jgs0UOP4x+T
C/SMKk/lDs/QSOHPA91OYsCUQlCvWPsUFf3P1Td1zhsVhj1qE3mXV7SGQ1j+ijKp
6y/JKiyndyCxjCBrxzT4JgwzSPFUNfIbkP0iyTa2ovlQGW3DeJ25fnkLiVDaXfDT
pZmlrQA8S2ZStsJEb+y0VMfU9KGFpri6gO0Dh6T1egdQZpGmjvG2g5syhEcusC3s
IbJvL79cXljXhBZP2o3NDTmZbHrAAAb0wjBpDCKY2leQQS/IkIjy9yt09j9LTIUZ
nwwfJXboMcowhZ4CTUIiovvdaE7g/sEcT9KqdmjvokIhhwSO2Vnc81ZEX1q2oTLL
GO6ux+SKAfhYvaASaIr7J3DQToKiCIGJX64LGG/gNHYWaU07IR/aZh7bmAJ3vRL1
Mb9ff+gwspPRGt6bIbeXlphRbI08GWR4B2P2vHSaqM6MAUyL1nwTlprB4EVqtwX2
08/MYPTl1HjQisQP7YyfkP2+p9fVQ1koIDHLlGZ6MQSUgLterejMg17QbU0uGs5y
pIwgAyUUrDrQtfmyzd2w/5uFqy/VALymd1x3cmDIbFOiyJGDAjYGrrckCs5KmCcp
cDlJ74lavkWCNwLR42bKYJbXN8fjPMWLsJllvxo00Mv92gtuVSTxuhIGYSmIpo3f
6HI/ueMxORvMPtuEG3pE6jwaxTs0XYmQTbKPqmJM+3yRF0Hl8PXoy+oGjzRQW/tF
S1lM5DNv13rn2Kl/3AB1RVyIzTFWRKk2NXn1iz+12hsSWRx/g7bSCiDvH/3NZi8n
rTj16OQoRum7eBG7oRiuOdac8r7DPQZJ7USS5B28DySFGnwCKjqTcHb2kMEvDq0/
uwZQPQnoR3e38oOBaaGUhL0J+Afb8ERp/mt2KCHeQNW2tOAxbkbLECavXZZLEC9g
XC1BCaYxC/xMgW7kAQIWW+eKW0ugCLP5rwkeU3fXe7MeE83/rCrw0rQwLpWh1ZfY
JbU1Lt2nOuRdNp8MXq/wQc7ppGwjnF87cZScwhOhVz2POuZcRCc7h92yjlE7Qaeb
nZPFoV3K50+M+IEyTZfdDfdkZrnJtbt7nJN59WCSDyqPSiWHxmmmfF35s6sBYFiJ
AFvs2TEgWLpmOF1AB5qPygwSSTgAygO9D6no5M1X0iewljLnivNMrMa6ByRayBvi
4UTsvtYw4KAyj5Dkh1bdzRFuQBAG1cd2DsCuufcQQVJw4nzy8JD3pI1WgwA1BXiK
HvRsWaGwJAmzxUf9TKmReChR8/M9LV6+LIWyqCWN3Hk5czZvLp5uTcTCC8L25Z5g
b0mubNqs/B3rPE30wnRPd1BaLwee6Clol1UKZJ5nEf2SWZEUlT/Qq3bMBCxR0aNj
rMpGCwUN3ujdKmnYD7PrZgIkDr0BCn4yw/zRBRBLa2R4URxkIvyIt5v1kewEBQTJ
kwAgD7B/MIMfSp++d85YOxsdr35qrMmFAlw8ouRdZEXkfBAGH2SmiZTDV5a4MPF6
ri92IivZyVrHkh0BoXD+weR9UxzO2A2lucsrC+oZ9oCcQWR12TYcQYhomB6xDkUp
sE4BMguO5rgKjjWzxv2qP3kpPR92s75lIr8rz5iZYY6I6cj0HCDp3Py2V0iCWYbr
cBP5xszfq4U2LXwzZ53ue+BK2wXTmVeeCjJMyuzsWNdEPnM17itxPnmlcLdEhZHl
shstBPlsRD1xLkEMNZUogsSp2rbMbO/SayLIFW7hQ/dM+Fbayyygv9E/8QAprQ7T
EUtWaC9DVpg973D3HlvUWaKeEZ43bjA6x045P9EAXvmct4mWT7aiYWzpkemECpDf
KDgNib62ciMw7OVc8u0p3a+p8BjbkOyNdyQo8nWotz67gl+3RqRWEhqJodD/7SIG
HERVlGm96jesldHoJ8I6/h/AwCsnFf5be3TSlYCnk2qAOksOJLk+Rtk0knkn/LAF
QzBu5Cpxu08nWHmud5UUP3Z2FAa4pkABaXZpcbf5n4sgiQ+o7iFsEjygD/vwy4Zs
jnlRrXPFLikEEDoOQpvbONv3fmqFhE98nnO6WWdv7V9Xf6OFyqdwCsj0OcfB26jH
V8bDqAij0WPdAMVT24KJrFhVzb34B1wnhu5170PpAN1eBk2t3s6dxmcpX9PFBs+J
QMObFHAYA955FuUcyThlP9bYYiQ79fOIgRdLG/gsK2k26YSSl/tdnaEq3y+9NM7Y
faLwHhteCpiYog1nEb2YXkufqHt0pGMZJSZqEgwi6lzarPX5em0dz+6kjRzj78Iv
QkAEI3inbucE9PD5VzVS53gWrjxpps9XxQJXuI1hGmtbQUdpDkx579XSF3ps9680
hQhI011zgMmF17oUp5wLEOReorNOTkbFnqdh77364DUShxmw08oZUvTGUzY58rxb
Y0V9CmgSJOZmgeGVUgNz8LZIBxlla4iYvOIafWyL+FObqtllCyCmWaClh8PHQzD5
HZ9RjOnkdVy1KCfF20GvqtccjEBkWs/B9TsJmRK2fG80GMVRzoJJjCE0Y3H3iFVC
r5P+w762gdg/TA8Qa7wssp0D94PDYKma2kwbuZ/jOQ6/s/dLYf/vdaMjhdopWss1
lnKVAMd1iJe6kM8E8VpHlgT7J74NazKjIszEutMSnEiaVvqac77FOnkwakxIKfZN
T7m2W2rUmsJq4dimciz+KG4MKXCw0eaf+6vhjIzwC5TAVOaOPvj93/BJSILg+Cu6
I9PYv0YR+/QnLhuUf646WsO8TrekTVQqMX/j7mpfKGStGDrXfOGtjBapYci6+suO
6E3qA7Tw7ZhT0682f/x9q1/HI6DFqTQCDxYysULX/7vVIiyTkHyWWzKBCcqPd3RI
jPdc7gY3J1eb9soz5p+QRAJ06Bcq1gXXq2H94QP+/JYjQ9o2rvDAO6HNpBlhSc0v
AUwkGAfIiGQWYWjBunwIGtTf+Tv2/vXV8TOJFuqdCvmMZMql/Gh/PEfLEzaWNrs0
LJ5MGEHB5mxWr8FBULiCdB+uNHnnpSyaXzO+/3MUGQVMhuhWEjktAXT8UeRai3/7
2QBdmMlvWMnYt8KDaDFVD5pgb7qY1UVJhuV/ZnP2rDhfV8yyxcuUYLdrxKIaRzHV
+ZrbiuwfhOUlmgVhq1xDWVH/8TagBH7FfLSNE3Xf9F2Mk1h8DhpqHcOuvBkB8gDe
S3bDQSV+VyyAVlFDkaLoDC0aSrUn5OCnFECZ1wboTODare8KSKLyVAbh6c3DGDjs
tTN36LPLjg+dNPHU7HxZselXFPaOgxJzZjT6VSAdh3qWKTEIblfmknavvJyixT/R
ZuQ/wNUO2WHZw+tvQVVmIZe0NmRWXiBfXmxBO6IWU+gRl1ujZkWysuXdsPvp8Pcw
jfXuhlSPFTJx/zr6vflZiuAEEJM57OcWJx2mXl/r1U6FfsE2D6CcQLo9i7do+gtZ
JBnn501XqyHLVJwJDq9CMGQTRlMFXEGBSS7zhcd0cSH6jc6OfvZXQhMf2vTKvit5
tGMX1ffn+92XhZ2LKjsbBQOvds3Y5gibIGA5xDF+rb0c9Jz7D9HsKHhudxtOpkH9
ghsSUeajSX3bxJ1RtUJ0gjnOVzLN05nol3WcFatdE1QSmQ/nPmr2ewswejvSoV1t
uDQNAPq98bxH+P3YPfsuj6m4Pkx08LPvFwYvMK0ejvDMPxkK7a/zWzfn5E33LGPf
6BBzXUR/H5GULkghiMN3sobRkaSvJ1X9RNhX/6ZsZGw98vi9aZWDzJ9Qak2chLZT
To0hDKXq+Re11Qw3oa02TnF5vgzQqYR9RVai0qbDuK2VbFgGF81WIYVR3Xs9l+HS
SUoBtkEPaE+kd6GEUt0HsHZnLJ2r6FBQ6ZMBH+cIkRu04gRB086nMrxwifXJoyxp
n91MJRr7ygTp5qsuXddmVmPqBhdniVuo1jv7/Q7rQqE2xJ3RTa1GZAr7md2lVBD0
XDA2UmY95xWwUIrK4+2c4vuMK0lpeNHWUlYwv5QCQq5+rf1BI1+GZPK7cZZvDHN9
uQv/qjbS5Ic/wNaHWjEDrF3pqHbV7mRbgMumzrDp/hztTlCBtE83IqWUTtxZqAj7
9BJwuYY9CpFnrG5t1vRwiiwG/9ISSs7RLeOT24WKgSbubVsfnpnGkdolwom94z6e
bh/d3drfVLLIfxW+3hCpKFoWdYSxwbDSX7N4yYTF0Nl5ICxvK60QNWXpGJzHMEjY
xsPmDbZmi5vzHNEEilzKfkQDRpsx/CPBUUPF9e/kYXobAU04JnCT47TEe6B3wKKd
Y1HqyozxiHV5ETmQ7u5fVPuCI+sXY71MBQn73WUMF5EEuqWvB+AExLyH40iZCiEw
U2zN3WY+uC60yQhu3K0iHM5TBgLM9711dVlbiwhmMtwbLsqQhxhSg2va8PyGYLj1
M5fyhaXm7J9sHRXg9fx1ZDjEDdQh/1IkJhAf2eiuIZ5t8a1me5oFd+7NstN17B9x
N4eOpCm3DvIRlUXhm8NokfcqOATvDlItmenPSGTJy0l4BbwqebM2yAjumKFw6CS6
nYSwQKtpXAdf4WSCDpAVBhFn+YaOUt1Nd9Cm1hXp2SXbFvbc7nCkehFvYlvE0iae
KEqZlptw90s2Vza2nztxsQnktY5gdCqgBg0FLAM/VzvnuJp/uVozQMtPhh9Vnhoh
lHyXPA6CVxuvp5nqLa5edn5Kj+no/4Bk3DOUn6xddSE0cs6+PSpmKJKMHVqLV6Ki
B6S0CKLVGmcab6Qrf7XD98BAJLTE6IWL/QXMDO3sihi+zyjog+C89m4y6LZ9kbbv
y38l7q/j9o4SfxOOnLFczaLxw0wKTxmbq+ruBmm4N6fqjo+FxW2cH9YqDrXRxwdj
hWfBJF4H7EmKibokfUVS9ZENpuYttwvo5xZMWq2vQQGwCKDnt/vxd+Sw/mrwK0oi
sO8BYVxNRcKnT4aJSi7XfMMxOKPcfzOijfEhSrhURCKeNM/B6ypEQjy5HIIMYSKI
oxoVnMdMWsGT/O3eXjwz6WEDPA72fs4X624ZtocPY9Wk7vUzTvlNzsYC5RlmHpKe
ng1/3i9UxSmlZPvrFjpziolP5JG2owmNCXLbO1N3TOHZM0PVdpRp/sctatE6xfBa
m383IeWjiHiMcKBvKz3AIjgAYbXfSdAsnU4VXCtvZkcrIuVgCa3lNWr0gaAq91bN
79gcAau3GaM1iR5MVlxXcBGdeEtwyUS19Ra1nTRm3XWRrwcUzes2pbWYbfySGByu
yqczRhhAet8gVhxYO139nzd0/MD8rXLgbgXBSaF58rOahLBtkvr0TLmJLKFxZzm9
QN9sNBtQERsX113Ndz8DUvOAE58466mVKxzay8uPhkYTwSNjxfyaxst5/hS1VpS0
3zknvYb2+C7Hi8W3lWofKRZVDpZndEnDN8CEd5j0ue80LWRUNrDoWI8k35sIC1Y8
W0IHQCdoghJIFMF4a628K2Fdg5LXt1XjFgPVL9kxAlQTMx5kqs8Pu++NxKA4tGfg
njOqQ1MU1C77dj/uZgpUk8O810o66Mg7mc8kPcxFCnEKKRkADx7LenDrG4aE0FDP
ij55x7Z3r3+jFPt11VfKtxf6JON8NZk9UCvr9PW1csti9lvyc83OuCzNV3tZ45lx
/m1BAwqGFfrLciBY36PYTTsUAHAhCKeKNc9c/OplrdD8SV3RjwLxT8JYvqzlYF3g
k0s9BpwN1E2Lo4d4TQv8sSkhntbFQs45mEp2esigp7CC8kUXoD2mGCdN9dp3k2zJ
ZqahLx+F45tC+e+bPDDS1kptXn9obQX1KKXg/AzDhJ3FRRMpBd4ya8hTXcRviV5z
y60mZyZKvnsnDq1manXJrxfoX327pIG6XZy/Y+aMYe4RNT19wwEAUhoQC9GV7gJk
nyPCX8ESBNzWLsUXZBZ8FJitgJBzntf+d0+6Z5I2S+bJHZq+kGGJ9wF5vUJ5qUfZ
mF7SMrDRah6aE0I5badB9CmQG15oxlyaDtgwiFh4lDtoHa58/I2BIuJGFsK+1kvV
eJJOCZ0KqkmsZxxkX6NBOGnedgVQfMfrgxSpoFhTWpLg9C0zLETGS3xAJ8K09M4s
eNjxmCHoRTAPbz8QkfbXq3UXhUbK3dY47a9qzSUps8aPQhkJFFBL7YRWtx+o4h9P
+J5fRYpVQlYMI0p79OQYQTrx+fkEq5+eJ0NRwEKJUuJgzRRkOt6npQkOpua9GH2a
LkfQ2zxunoU7jzSvNTHROHi9uq1uzz7aVEwJWYZFBfBPBxNAiI6M8OgyMTECe+s9
NAgE2eA1YYjE78kkF9p4inGC2hthgkXJmBJFkyVJ5GaxhRa9+te48D/ittspT/fZ
HYxuXNGIsJCCScFH8Q9oTAs44kw+jKhTLr99Oa6ZUQp/qWD6icrOozuC7Wd5jSEp
BXmIRJTNqLs5WAmfVKBgLzrfvxqks154pAx5Wuo2NqMpw630tqOhvHq4BiFLLszy
appZGAJcodd9qLixV6gRG0rKzxzLOiCQZ4oNavZA589H26ttGMvL9jwf898ZRnwp
/icv78vxWgb5vB2qtVA2hj2O0PR36p3wLBJhctIsnhQL2txKEWngdRGAnngviDxR
Msbn6fxAfuaUDZWf00hbQTC5KBAcM8aPKKJCCNvYnEBKlwbjnpoQtRZ4Mj3HJ7VK
OPfXjIb+67Utgu2hTbQwkH6RHNMmz30EkNy0s97NiwdrkNGwulcOAQfqdlwZBVFl
PVJp884hhrOjRmW+PGPe6Tz0nqKj92+p2SHQ61Dc9WsmJARjLy00gBVnrTsU02dV
rgxqheQI+qjletLNe9AgrLA4F5vG/BQx3rqZXqxwyelyWtyoTqS9dT9MFmS4Tg9r
3Rzz+RD5wgiHzyVAzcs6qnp/K2d6Uu3XHtcIbiH/iWUR2r01kvHMtjfcl/wOPqk5
QV1T1gsiPVsCHfnHUyQKIZnxVbcaXhHLj+NO1lWqJe2g774RyHqW55KO9EBsjHQY
m+o46LLLSVOBqB+mNnq5sRDJDNEk3uUxDYX4cRYWcG7PzJkHEhBR823GhAUyHa/e
Zdp18mEPcKC7NXG/tvxelavkKaixyN0kr/6kD7dC015xOf6QVJdEvSFuAjD8gExz
m4+miNvYR5+OvDJbrwxpmr+UdVQqKzcIZYIWQWHeu8yCXuleal9EIU65oIDIM9Tp
0FBMkeN/soeb3rLXuQCb97eVxEnpyW6QKsL4gzg1iQG3SQt3eQKVU14sUQiRWwQ+
W/d4Ch5MD1OVrM8bWLS1hR2YLyjDvnMKOoo0cdh1ft//OKLsB28A0n2mc42mJ3T8
HPrlpDIZ5wPzb5dPfY2mfohs3ZhBVm/zv4O60du5zIipJf2BlAFHKLeCkO4S3XuI
Z7xCYlX5sD9MYGRkqzxJW83+1SEI1hNnP6rIWJpFP5lrfd+1kCWcBgkAQk2lYRGo
3Qphjo34dor/jJvhHGGqsvg0zLws9eXa1XwzF50WKcPVcqrplJAZW88XwDjoF9Rc
DuuPXEgOLcAjXpAbOWsTH8Vvau7Y259zfgmMGVN6Qq+YytIc38ruCcO2IGrlqdb3
8LPdcB/rtYhDpWOnLqOfEaBsyTcya1+phISOkiJkfiwcVjC1/oznt1HZHv5qEpGj
KZHSuHkA59a8T6zMm8k0dwfFGn24dIbVA6F55S1XeMhIFwt/6/n1V20m2KZhmRr9
AeSydlVDjR0eynUP+zuo0Z3MiIO9Lw0Ig/M5YAT6jPUkuh0hBOp/587se2C8/GUl
0BAVD3r065epwsiKXEkWgxlVa6Rfa/w3TeW+FNktAbVRXDZ7hVBIO47lFWsuYexp
gfJN82j5EP1AytZFafdFK9Af7zRpA35QxoWQPU0zUW6q152ePwPHc0LRA7TXg8LS
Gwl1nw015Wia6mj8Mg6Wia0G+C2u4oITQRcK1pq/CYSQX+OLejlrobOZ2pYsHRTu
PlPGNXBn301x9FpN3JtP6VICXMXX1QjdI0cCVozfMIjrJzLqQcj0zNwJg23qOxMZ
G8RR/mhWpOdY8Cg4hHcyL4SJEHqeARBxLY6s5p1mp8eyFL0YPe0pc3BQa60UE1Hs
Xt+vCh3zv7bpHXysKXKbVGLQIeOqBXMIwWWQ/lweHzkrSqmGqrngLZV5cqP04tQ/
3U1le7FpwLw+ten6p7HiQVf4pdQracKPW1AYTjelQZsFW06GjR84Uq6oA5jsgOSF
ooeZVPSmM+BO6Tc4CzHN7iWacddNRHL0+z3oVJa25+f+inYVk/qQ6cYzrBqyAjBB
Ozto3Ki/BXZWE0V2rW8kCD+Qx85XPLuFOgFXK7sKmo9jEEmoyNXeaGt+uxWWch8h
moRlzn4pUOCBzeEc5fBuFGvxgNKcltWCfvyP4OD+NG1gTaWi0jRxepJzitfRxfM5
L95Qk3hAL/CVXa49vNYVq3JhXyK8OLldYylnP/iAXzjJMYFjsNPcQvu3YirKKVz2
bt4RM7oSsM2kor1feISfUKz1ct7rxaruCDnbSBFqi3P06cAq+CKmi4am1Gmd5OUm
XG6ip2BY30C7hEIQa56LhU/NbzNT/rtkLUT4XhwM22Ud82+2AlVkUkhFiytbSdHC
WkAaop25mh+qV7AagKng/nkaXi4SKVQNRdxQFsyhQrt4mGLuQGnZ7GRRMcbH6NpD
mTW0FbtnU2COsoSJCJEHBXlxxPdFrFWTa3U8y4Orl+8LRm7no2yKzNnh39UgMzjx
Ad0rsH+DLz7Mt/7OnWvCm8s+MGesDT6sp3BYyalvJlZs5rItlmp8xaqoNJRReT22
OgdG/iSuKOTqNSTMvRckme/jc06IMM/c00yCawH/fc60q6eg/OyB4qwXVM7w3RCY
asiuyQcJFoWR0zcqo4VI3DtZpRWq4+5QDbdeBwR6nLOtXbBiXnY0iLCIjKWxLPGm
UUh2UbfOEcma37WsmjtYwADmuxQuRri++6q1OxAAex2/rZ6JZn4VWoKRhTQSQe8K
MQswrbkUrVNvu4oVzhMR3fDXpEZXjbJl4U8oNCK+4F3o8HcLnBzaxBAJmgVmTnKQ
+cZTiYkRvPJYZHykLkNDhcLKD4jiJoYf8zEXWehLjvYTkxqrkKyXrOgMyA9SyLsq
CVmF2p8hSov4vAOZe+E27E04LrwJrEvNlCBwFaYwhA69UIiidp0iIo05cPdV+C6M
WOd+VXckbI0pWYFxF2hg1RSsMI01zQZDbqxneeSgC08Lt7ZigQnUSyhfT4G8ue1T
CjOOCxdmPSwd6YoMCTymnvVcPA7ExMA9FTRvrtiFIHs8nsudfNuaRJGCxzWmgbki
42hWh6RB9TgBe6snEb0viTmB4K0Ow33ELIqUdg1Mmh/lvSbYBENFV4gCXox4PxjF
mquMSqPOQ4OyLs59KuGO+F6jmjlzw4e4WZ9PFOxXSC7+IsBU56ixHqcWOrK/ELpa
ZT6AybaGyKtcOt8tcuQXzy0LrWJKZcHqwcSpNeka31VEjOHYaIkbb+J45gHOej2E
l+G/yrJ1FI/PHRLapr1+fWvkvVjGkdirw65lVrs8xj0fYYN0dhoNodU0Xa1Po4Bi
LkJUXSm4l7o5J3Dc9DXr2RtlVBEkXiDwuvaw/KajZfZ9O/+SQu4qA4I1AmTVFKbR
Gih3gjtfLMxD8np4yo5SUyebqr/QPju9Y00QOSJ5HQhj0DlRWrgtLXRGL7ApyMY5
Z+/vgLVpqjjkSEV2b4LMfgIo9+ZOm8MiTkJIl0HlbKCmIZrMD11SFNg9BHIUgwOG
49NlqI93ixiGITQphM5EjV/MeAYDFnPzJAPcyoMIt1Q9eG/bRq6iAX435n+Ok5gq
XSi0ovl2kj/z8lWEBxYAzCjpkptuGyau/nvCPlwVc5fSExRblVLXqXurRhnn3DfH
Rb+fQzlOFHo3eql+apL6TzaME9npzlTEZIu054eO980t+ZbHIjMMRVTVMLLCm87l
WXK1AtJZeBkGx8p1qK3kVY/wWvhk3BtXBe0F946kZehnPYrmqkoueMk1Bu0oPIAA
vF18MXZCVGX88y+HUfPS21WdFQuiXj3K2HnDxYE38gdB0dyBY8zSeCgtR+SkGXZ7
5aQltDYLM0eHJhgN7d674K5ANKNaDOOim7bw6GHyMpvqhrgUrYB8vEZTasOG+0I9
vMA7ImL5KxuJEGz2oml6KK2IdueLb4yIYkU/HOj00mxwn4NgGRPZ0VYgdnm82ZzK
qfvkzlQwStzSxbpPy8TnaWyOG712VfV6k5upfWJqcfWKZ26Vd4uqNpBDY/i+Y2z7
QPtoQUTZtL11/r9nIBp6cyhEIJkn1eMw723YpMhpEoHQ/VvADE9y3r8vNDMj/DIZ
D9SbyqJCaF/Ew0xvc2LgA3RqTPDfpuBJtYo4wagUDoJTBtwEBgxWNy8chyUlWhnL
9ZKsL7ZPO1MGV5T3D0UuXc+G1eh1R9Hz8mktFRcstjltC5bdpqYDVKbT3hvMLdnq
N1qPmIHMMCJMRpqP0L/g4/SkbDQ2J5w/2YcKWzYJbgdsgbvcTd44DBATd+uWfoiH
vuelf1/lYq3bIarcUIy2BHOvj4L0tMYSalaGChSF/C93R8/yvZYLvExVFIf9OmFI
XHT62SRq3tmECFV2LVfx/zYLZ0njIGpd2zsYWKTe0eFvs50ZkkX3696bVVlJC99c
7lJJVCuE++6kK5rTjiaG5xHrySbfd/oMzBKRyeQU3B9wlikSukUkmOa9zQZpyEPf
5p7XHV+5p0QsMB4nxgATxfpoeyf759EtO99lWc+k99yxahihX2xXJ2Q3lvlhtyzc
7FKnFrNR/ILPm9K09dc81GirJqjBMvwHacVtfWe8DWC8ENKYKlzK4JQljgOGlR8v
khw/+VHzkZxgL75gF1hA28Y68PswnYW5sM5lNH2HNt9y0oAi4+MkRo2dih6LOmjh
+0lGYe9pUXuaQYuBz1ikEvPuHK+XYS4zQ1RhCmZjxdP1rY3PJ+ajCodTL9Yd7TqP
g/T2PlsrI6UylMTmkV66+dKNgkvUmgAz/2ofngsz1ul9KKbTjnsuawD9Mck1nLPG
cOcFinj5pMiuTFXUqKh6whIsdKN9Zu5nYnpHN/uYRrtL1gDMt23lcLhJFEM1urTH
VsEHuOfMZjFqaHJz1GbM5UPSaKAoCqdBIM17nqhEvqlJ3nG4OnJ5tWx/ZVq8sIlO
LZcV+lTg041+0kDypOUl3+B7F6WxTJvvynnKb8ATQTSsAJfs2h9gRdMBcIgo8PFz
nco30KNzGIzaYt5DSj2Lz7nog4nCz3vIY0+/TxjNjI74mjeNo09jSIGMbjs7zksm
VdbukuDw3FJODb9RslZMFqAkd8hyHdYLUbaWVTeprNIsFqtdF+1G9iIVefBv5YMj
5IrOGlkyAZquF8PmQ6Sg1xGl5tk5SWYnyNPWKL25rE5NXzP+ekSEu92mq4wrEsRN
Uz0IoIWfNpG0R52sI//YCJ6br1UV5knmHZTa0uo+RbJD0Xz0US3n0vr0F3FQ70Cs
yzxhdSLNRCNlror/ZPJS1RhlDgk/egHqx6A5SryuJGNY2pRI0C+NCpsTwgxOIVja
9/Fr0mF21AJh/m+rlLUKALWTCT+zdeqo08LG5rxGat0QCnty8LsCtLSsLoPMiL1N
dMTZhUQ5+KQFi1nbCrif3AuoXaL2bfLI+O7+2P98cvhgvB/oigqWusjgf22X2W1b
TzcDpWGOethviuwsP31bhj1M0FU9sBdbotBsKatMwChgsh/GcibkDsQI+jjJ2Tt7
1oXd84GWYMPvi27xd8TVPdpjnjFMgeONI9ClMfNlc2VP3qZduPZHr6qnH6aMFl4v
msquNy4z4RM5ESZHbpdStgZvcd95r/6in9uzEoypL/+0AG29dhIL4oVzb0lyLvg0
6Rp+/T/qiy33nXRCdMNMSh5xaiAZER5mbPMhoD/HNLDlmKXPSzfEEkoy62u//N9r
r4+5ys0rNlUAcUixTqbo1hntrKfj0gSSMxkbqnM64g0nanT4/gbVInOYkWDp7gU1
YnDTnLIVYUe69+tGubo7YrAL8ZelkbgddsPwvfKxwtsOg/BCZM/rE2FmbQqhesED
rQ4I1IizPPuheET0sLpedcVxKWvyvGh52wnhWbS2+7N0qpOJFwqQvmGcYwDvcit2
2mV0sotgfJw7n3BoJWV5NysHqPaj+xomJ6g5dWftOR54vNVejq9GptPYM8b4QF+U
B9xAWemE9QYZW1rczxA2JEmYaWRRx8AseZYauGd/za3XBSc7j8JIZ/+A+iJKVL3/
Ua+CsAI1U9MxJCf6fCBGXhQHB1WWLaSRXrvAsuvinpv71qkV6Jg6HZKjvO/SZHgc
Qo3s+MfXa+sqbqVIAbek0Sy+HJ3Ze2oHAvogE0KzBBzOM6hPL9ALuI7UlxQUZ8Hu
d62IFQ3EPLpGXL2HiyK9hzUyTmxjss2uX4LRzLLuhX0YY6OWsE2VxP7y2aQ+IEeL
jAuHXOxpwxf6oGsDgSfkQWU9ZsuLiYn9/fMVZIIor8wTiLA241tdVakro8JlDur4
WFCjJDozMg0tvmnfgyXrMlYwJm5dfaFgAmi+0azBcPmiAf7oE8Dg7BPcSchJIuYZ
4SaqxcQyKx13IQdQuiykWW4AAyUnYAslf3TmWM5Rg/Y+5F315rjFJAYPnhj7nVDH
yDAA0JwISt3r1K8lGV5rsOZFrY8Z2/ivGonjK4EuRcW+vvmDWQ2xrSmNzaAJZUmg
8D0pEzXkc8L6k1BuFOoJbeCVcUVGj/Kaj36io9XaN6XK2V+RdymmZ6sQDt32X5yH
6PSPENNk5aTqec7uswbkoqGJdeHi9oRumg7aNHdb7bX2lGwgoPWuHpQMIvDO3cin
+zufCyUyib6CJr9HARmwxAxRSabTtxDtjOTwCLJu7wV63TwUZpDce56GpC+vwsYR
Q7eUwQnCF453HUYa+8c6f4dKCGD8sZvkg+CNYSN10fOxxwrTsjREeCPfHdzdvM4U
rBFZPiWvEuExmBTsCkQhZFL02Tn5gNsaiJTrYEHEQSuPRqT1aPJaw5AMQnItc3Mf
nL4QsqayHQxPDcP0Tv0KlJCGbIbiBs35NLbkORpgqpKOGv1p3eDD7zKSuydy1PPV
wncYSqFvEH//ndJ2Tttw7tj5ZLV6dEul/vFpa4wKAwIl3SaA7YwtG+bKbOZX/+zi
k5o1lcWVypyAhrrOszMQsVRmuwLMtzYseTyHGQOZazetucUqP0Es5Tu6+bJipHAd
TOh4crYLedkgHC3zGIn6q9IOdi1T9StZvlaIr42472z338ojcHerjNsyk2YRUGS+
h2/HQktdPOIBp7XOGIFe8cENIU+SSqyKHF6qCXZZ7Tx1FISmOaMjTJHNYs0KYFVe
OAALc1HHxg7144ntY+au1nt9KDu0WfDHKN/hpOPrL4E/KwwQlUj18MGpQ1DUsFn5
G1VFXO0edI7o+4+fojVDfZiwFW6D5QC9Fd/ldIy73Gz1MCKPjGNTHtH2nwUPfkF7
PvIfEqKcLIbbBL3rM4MLM36a4YS9XK2mFg7IQmPX5tym+m+5YXFql/BwmEdQkU3z
3kd4IA60hWg+rqJGn7ktwCxi5x5pJzMohM5MYAyEslgYn0uuy7qnwEIkDYhapFBq
SzmbUQpy3kt/M7N/MQqJrnAfEHl6I7P+P5zNyfd7q6SSihdcygXz3IjGbhM2jrCt
/nPfCibSpXQQAo0Iqx58RnLrMWvFUQsuMtPI3sO47JBKkFKoHdkV+CPUyRfeSDbw
vXkbJyyHiAyr5YBJ3OuGnrmdcwSjykHmVXGUFqpAhbYt++kj0V4RcVzlXnYMJf04
/aFiBc5ot34sFbfCVbvTbB/PdG1m3CiwQTnUKfjmp1fPdxrfQSfZ5qJ7Dyo/lVHi
uFM/0FVzTMPs7b9Jm309sOQqMoAlAWLMDDDDH6qZpXNCESAHQpN9hVXffldLg0a/
rLZAe4VWcBKYQY7gKYP5VGKELTUH6xQ9sC3ckgC4zqRIC39wofRUYEZuMToTsjX4
fo96nOY2hXXp6FMYQxDT2gMgNcS8SQr2+Eu9oZk+kpuVhp5GQecFdI3JkhrB2iUP
UL6Wwt2+0riu7zM166cCp2HEL+2yLrlHnovq2/Pt1h2ldRFHk3Q/BGhDLszS1N65
chCeOJgiUf7/47qhdRgYi5vf0m18kKrXNr3L0k6y+Tws93zUoIxNcPHfylXuQNJy
znCvUeLZuOSPQiX/MVtm3LX6HPvpNGX/Uq0S9Tw1LlQE8dWaVFgNz0AI1GXfzEim
OlIEufZJoT3cUW3Mh2ujSiFNHWRA8r1KH1m6uN/49VnxDD36PhP4JNdm8SBTumxA
E0nk8biXMa7QKI+Sx3B9YJYBnx6A0IKL3uNNcCM2kNlfsVAHqMSxXTOBvNHNO6jV
hzMSs1/oEh0btaygVfRZYac7PlWvzC1azATkdD7gb5QktZXJk+oeNRNK9eyUz+oC
FAUFdzgNN9Cdd3czFii+qAV2c1K2x+XfCHjIMaIPgzkYNjmPC4FL0f1RJp+SiTYF
SGb8yGZjFjBOnm3dUJIcVirV/mFssgrP/ozTQsLZdURgIiIcHgjkHNDkitvwzQON
lvjtztGh0mQlySmKgIqCLy7U5TzBAbhOVZd6MnGugApbC6KKUUHwEn1RpeOBr4DR
5txK/9GEZP0AYPoPeR6B33E74mQzlpNTxRtARycBVu+eBXzcky2lgGpyLSm6ghXu
PR7/Wwj4ORxMLmv1n8XGslir619X/8A06KqSc2EIh5qQ7BNBdt7rW20yI3OkFw46
ZQCxkCFtUpD1tEQS0j50FhmhmEscVhsc7dTlQsx3SfIhrx9gZofI+1PPJZWHVbhJ
TxHbRmna+ZCESTEQBAcUplFL0pHFwSvWcgTML1HCCQKJRvGnKEe6PAw8E0XRg4PX
I75gIrvfm9zoJPdQdPDdUW+oMA+nUkw7m99RzOEbhuzopPhVJ3ZPRogUqkV4jU5b
hE5HlFAutd1wNYqd7E5P1nwyBZrK+Q3yB2DbBji1b14lCdks7SLLd3d8rWIbxV2X
yb9bSm4uh5lLXVfILqyVwItgrD5ZV+jSqf6PFX7dpknB6ucmQ2t6rHn1OYUE2a3a
Hw9rzMagNXEIYjsyCKIzCM9r4FfjhtZKmMVYfLT7syCd5w4QogV/yHVFaOITKqW9
F1OVEolXQTxVuUKZftaseDHR9Mz+6OoJP+ybhT2BY1V1LyZSk1m/9FPNWoNxtyO9
34fnGRV2Jb4ZQJcX74aaT3XCuaRTpEzbFOP5aQxkEqX9COjpdH6IZBgib34LlbJn
nSJmS5Nh9C1xSocFLrZg/ER3oPCDU9HKC2DjCDR50i6DeM4goTUlR89557T8VAb+
Kp4HDL8LSgz3CjC/2v7rsvMXNnyPuOv0IbIV3U5k3e1mbgQnfSKcsn0+/3qKbY35
VpaBbsqYky8nuVBO2bpEqfJMq+3LlI11tthlVXLBoKoYm7UlUFdRCbg85WwYz7Y9
XAS0MKlyUcm2czso9F0so7n0gtIGyQ8QtbaKTu/9OdMPKqAr8kQYOmh/bxdhxBJn
SJrXyvrcB19DrcN3yZ80kzPEk1T4LBC+Y5Rv5gNs6P7fJ1XZMDwDzsnw57RAMxNK
4s6fF7seFcbKNbgssNJz8Qz6xmdIs9fHVLSgK3lB0lDCg3UoOlvbcZmXLra7tfQl
SjdizDUce9KT5f77xUAScdA32qKNZXt5pPWGMA8oO2smTZEcYws4N+uGZlQP0mqV
kO3BpQZ58HJtzsQBxt7LgQjdgomVLbKxEnk1/nwWPrXN+PlJ3vRrcE/s5mZBFatm
DIvzVsxpTAKZPufPVEVFlM8HEKLrPVfePsGu5eXmQ0/QY/DeiUOSOxy41KXy9Yj/
fnbOG3tETnTFIQt4EnKVkXyY2bpXUx5fEa4H5gmveoE2CwCJaMHVSiuqtjiTY+1H
l0weC0HWgS40E8tNy/lAsDiF1SFr4Er5l+ZG5BX5VgSnFu/pj6jDzxqD0BLLG1NI
nRUMvqkmFUVI0dCIB8HXAQrDyxwqC5Pi56MNw6mzHpev4t4SmO+4vLHziNnqi9Rs
+nDaHtlTZAOfpw8g0VbgEUHeATSxmYazc71QI6VHRgfbjYZrW/cHsKr3fYEMEv7U
YdVxOakGavVo6aKhqxRitV2fvJomrqas0P+qjp/INHGYU9YU+rTLArJfQ8fEKS1H
dr1/yxxPBLU4ytEEwS6oyXthbELgWzbtbG/ZQ/MB3SK6E/eW78aGXtGnQjof7pPs
qbvbHwc17HK0Fxdri0N30zSdJKA59B1mlNrCOLTMh3Sk8xKkf6adWv4cZ1Iv+5yg
VqeLBlvE6VzZ0a59CQoWBWO03LD/UmX8tDrt0v6qcnXXX3zpnIVeGZzWnBCUi7OF
3A5Hboij7TSoUDsFTDNBTj7EH+/N8jgfpfaWR6f8uePLSh4Zq0LSWlFphWLRZz6F
vT3fqeMz+skElEGlqWqPfB1Vg1JSvqAEMsFbQN69ghDcm6sqOKg+Va8jrsNZOAOB
Sm3drAvwgO0skUq5WoP4pDtB+uO5p4mjxr4QkyAY5BB5mNTwzlLMMCQ9Faf+CUh1
9+dmaNH5Osj45ttYJT4DwH+UfGjiKo9yF8DMMbkMH+qI2OCKI+uvHwICeuNmWu+f
EI5DJiWauc/jC5KRwIiQM/a8r4WwXxyDJgJzPRsUXbxLjpjNHpXa4vTa9eIKOIey
7aDBLdp3xyYzTdg1bmFWtlf09vCUGCJlIvGmy4zUvtZ3OUQEreSHn4URcbXvbfNO
7tSXFQg2aGqBR68wATc35kmPATl7t3UTpDkOlQk7m6hDujTg+RNJnYdyM6KLnXQu
7O6I29AgNqZH6fOpeRE+2S19lfCZW1+rIlrG+0+Ni4Twi6bRtNmRCzGK4MI5k7d2
ZsO2jYgnh0bGBcQgOQ82hhYBIwAyg98xRv+zFEL3JXrN08J2G02Xastisq34EQ3U
ZgN43/l0iXwUihJRc5o+uYfhEoz6/4ichw3Wr6hnnchp9yhOiNLGJBQryH83Wl8O
lUP1Rnd8HG6sjW8APueRHFQ6Q+Vz1Yd/6jYXONrvJjBJTWaiu0muoT2kWqydWolh
iBOwplbX0lPRJWslPcD5r+NRJI6MDrsuxMBHSjytB5+c8Sw+FWF9aBLR2uhyo8/U
NMVxvsNztLzDjHnvhnOQv08ftTNfHvk3trVQrQ5XpYn4VLYdeWvlkVJWv91TS6b+
KWGV4G+dAhqfn5JKPE3VJ8677FWiDF8e8BTY52TOOOjqZrLpvC4TKzz/cnkCZhuC
PDMk8BmVv/5yhdn+g+IkFwTSn33TQD6entdAItwPrcwSCvka2be+7I3O9r95HuNe
ELAZl9MQ1ElsPjCJQZMGDFREFrO/oTyYdHGi56kfXjKGjrgBE4nSO08K7fmuLxdy
L9hr4zYqCPXLb1VaUuB/j1YcUWKYdVlYP4ZXpjHyeE4dJ+6TCn1dk1vd+9wtNY1B
fwHp6fJdXznQ+ImjxdVoZHelOupHJfn0SQnFuP3vx4xBXPRD9spIfN1Sj2EWkeio
ZONuXg4UA8jfC3DFH6Ex+l1Fq1KNk1nZz6x93xORG/EA1vowsX6xYTYYD5Qffcpw
qUmMKipmH2cAQGIwSlRFU1l6Gl42V61kAUMGwtkwk2uwcMSAYImaDW38kx6uwPxt
iZOUTcQdz6RaWwiZFJ40mAQrZqHf5OgwBjJ9i2ZLH2bHWotFzrB6SGgUekPszvGs
QZa4r0UpDoC3qZlLJK9V2pLn6VyU42yYcotA4GEdb3MdTe4MP5VDZkGkk7FZaQYL
VofFl5DgZeo116oae6KrUBuzij1+0uftqUVLsu9neWLsnhsDwO2faQhwErRlxjWi
ES2YNjk1OhxLDE3ulbZjRDE3NFkx0qOAtOnpeu7xYCuhazXzuPyp/OxBMokv127Q
8tyCtsP664lG67/91L6h6TLNpcjC2/DHBBEQM6zWIxEKeW87IGgPbFomjSF9Sj7K
GnIl/mM7/1DOkfU/u97qTp9IKLOYLbkTpGa3k8ZBOPqn0vRJmDn2Ci9NvkPt2mi0
HnAd4u1ZhGskbhzxC/OvJuYm4sel8fIqnfxusST0cSbwbMiqFbZRbhMcrY5mXK42
FDF6spqSBnjz8MxpvDGNA/nBRUX48d3clhE6oeY6EHT4YfqIfGu0iNhD7uHV45f4
saQWUBMyC+ntfD84YTc8SZHDrrnxdHLb3IcIhaTt6woNFlMEOxgZUXA53o6g5j3B
59IrNZjpNmcKupoYogVFXB7CiYsimjTBsAXPjJ2035I4WOUJ3pxe0gZ3KzhlzhV+
yUu2Y2gKvkV82sEhP0PZbBT/hLxxK6e/dl0dayvB26NJzVrU1dyArMd2Kuv7QF5K
ZdP7jGqY/f4M+PIpnwQXqxWLTNnOiNsJv55+aeJ0AuFV246nT8YyoADtOOKdizqA
j8v5a/nAG+iEtB3IKcTRLxYX3l/ND/vDXtAZztlwMKCZbl6isGZ1G6j1YtAO3p5/
uKyIPDRiFVcF2KGgxjIOoDJVKhuGYFCR9j4LkaDihl5u5b1VPWMN63UJpm4iONNN
ktQkDhRZoUsvZHHTjtc5stZmKgJ8EHSHGD2ffTg7PfUUQk/yAYW0zGEK5algk5QH
SpYH2rnyiKYvOyO1H+RNNpRwMtg0Y5eRDuCQUgmHqa5JuRfLukMR5vq/6XJgCDNP
v65f2X0AG2GTW0cxqPckkIamHuSZypG04VVRIVLsP73aR3i1C9bDlSVKqLbGe4dv
aThp+0ObRk/+QNgbIlUBsyq31h1eWW+ubazITQoVceqHWgNpXGlmtbnbl7crY9kq
hcOXBKQ2oNQkd4EIuXQ8Ao/gUVMH7/ExenrANNh2YikREWbZDJmKLPO+1EFTQsGT
wvg7kmPaOFo7l88evR3Ki34nC6o2XcqFXerP3+RE0eYGmtUtqpalsJIBAK5Y1VsE
kP6QRvmbaCnawc4er54XAffpxk+o2g1aThJEaeYxnIKqKGFW31OduEMkjtSfU9ST
RGK4p2RfttGhxVNIg+lcgLEVJXM/ocDzoQC4D/3aRmnST8VtRQvAGapG1ygA1vsR
92cK3c4jkqpIztpcYVMDZozU4IXGrropzwg59PEtGraLHXBO/xWiq2JvM9D1whfQ
9yiBXmImCpdDNeylxh5/uw4N95KL2QeTKdw0+6yIq0bVSW6uOcXFEmedh4f2vPWi
zhVnF7wfZYLW5bJWGP6wwFA0M04fpULvCuXAxHG4tTsQjjnkPZGqBAEzrntZNPDH
9nCqzEkfYjb2tPKcQNPk95rCGoYMM63G81I8fEK8SJL1dYT2CdXhUspZZxflKV7H
7HnQQeO8X8fEyWjO4bAbxyNxoAAvim4KAjdZhN5KVT601BthvtiaXxUDtVliUrTq
V0EJl/CR7ytAB0vJBJGfTYxNYiehA1KbQC+FLMHTSlbEOGzT9+9XFnzJLXBZ1OsX
bWEtJyCT9rwwqH6sPstYtZdnfp9Hwtq/1ec2SR9NmsTLzdgYQm+v2dd8iDvRdT1S
9eLjvqldCKx3Vfuh4iWBD0RlKC6AGcN1EBjTlacSmjdpb9Y7N4KvugQFoE1xjk8f
k6vPA2ETNPEU3oEDVJfv+/EFJrD5UFBPtcsds5h9j7mPyh5SmLlAFAis4rvVDS28
pZQKstp7RrflRVcuz8ovV7o26KpbURhm4tZTTWUd4a8mEu5+N6WxvMbI/uDi1yrL
oM/XjMiYDtucQkky4O0LcIjzih6/fmVfLkpbMnS9M+z+UihfNTM3JgKhQmd9BXF6
RLPBUMs179GaLmdNDUQXHGMq2kC0Rk5TSzelbTGVlMse4+67mRqavSykry2gMoL7
HQT/HBsnVbafGvFiRXILpp0d1KtzQZBugZdaF6PrCF+4pJ3+4qk+YZrMJgQsNCiJ
bweyt+frMTl0vsPxQEypwZOgGoZANx/75VEWVz1QLuzqsDGqz7Q4LBMXXNX+2ubA
qyaazHFtgD/vnCvaH4kRwKIeeQtyP0/NPq/scJtrH6+Cr9wq+GXCS2j3w1byfdOZ
FZTFdd6qKDZJZH/7NOzt+gCWyxAm6Sez5qomi9jxoA/BwBfB5X6bQfyXbHw2RieK
yTtXfqRNWaWEi7BUqe/1X8kevjWan6F2XUMqshU30z9AqPA8k6lAA2MZAQVqomEq
E2DZcin3nSDlk+5EvKqlm3eIEkP5O+vH1KBkwaaFWRq9dHDuXMXKStvHjVFOGFm2
OUORv5TJmfdGSaXlTQ87IwwlzW4sMUSj+l9KcXKUcD8u8Dbu0kVcC/P2uM0Fmc43
XXv18zCRPp/9I7AadwltQtfQdqZWCPSqvNDeCjiCDnkxhX9gJuJ6zc2rF9+c/cgK
eWWnrsqnr1kuaEUREvKOWLt04XCfPU/uDke/Ic9Y9Kq6vHL8hNOYWTU9EwFyBHMJ
X7BDihEOHqpbClqROCdDFjdI6ENXaKIR5vR8vqNxMDpQZ0IDUYlS4befE9ymWviw
ZPRc5VHaNJXlnKx5HTTpQQfMSCdbS6AjvSUXRchY15ale5whCdzC93j38QBlQ0wx
CxrHunNLtuGFRmsj2ixbE9KUCkX1fYDRP4VETeFMKnhMqEvTDSpXCYFbTadfQddo
uiFJlshZy9pDVXTOdmNclim8gD+mPLmhaX++6O53MtLUwM/K3hUekMZau9j21uGn
1QgqHMlxkH3awmyVI/9vAAi6aqbcy9bMq5x4oAWB3dTJC2pTcxnALG4aG/5X3/cv
cVKKS8AePzsxPZjDx8+/x9MxyzeD7Kbb7bcrHVms75jYQ7aOe0CpOU+ntTtWZfEm
4d7MzO9+JKspEHb4bxHXYP59EdhSoBl4Akeqpckb6l5ACBFS9p4GeQoJUFZ4Ho7U
iAOYojIBSE3myGkhYruD5v0Q6pw9rAGs87aztDPVUlQP0ZfbQne8mPxjbOjjbyBL
9SYX7DdNumvXP/DTfJPnWXvYkjp6w/0PZXVbdAiR9c1IIc/SSMkb84NyKaROViZz
nlg5HveSzaip3dumnf+WDD8tqwQ6eSoK4bJoVkeVUQxVNhzcHRTF0gzQkITI0ezF
U9IdKIunfBwQEPEBHm/vGdZQ+shGStz8f3TyYZB9Li4hFd3h8I/PPDFQQ0ZYHsdT
KETYRTa0sXT843kqyuKt+BpnPdRX/2dHbUf1WWSazAp5qZ1hCe4vr9D7HiDC0xKZ
SHE165coL669dYQpBoDJX//FV9+PZBunSpNdSffSqBbhw6hU7NV+U54WyA7zrGQr
gEBjyXBCiw4oriEcAPMZbCptrmtfnRsrETe+IloUeOdVuNBaHw6m51llzInyjpFS
8C+Y8zDnYKVXB1/Fm60/x28Q3364fp194M4m4jGKiFz3Yk7Nu8vFQ6cEnZGZ8Qzq
LTaw0J/A2ENbXrAuK7BB/3TO50EDf4OIGStho+wRx6LqQAp72UK7fvsTjxK3nk2l
LmeANImgkN366i4NYpJKGq1HNiwcHm4IqVEFJQtIvCrHbHsJQ4dOVMgKPu4H9svU
4hO0leeUaxeNVo9BPGU5/JmVoxny3vnN9Oze1Sh52kKgWiYZfldEe+BaQ9iRYNbT
TBysF1PxatBRxfescRMCJQ6B5RmhZTcS/y2zlK+MOAAmjdHTyL2xGT/VBlQB5I7l
n3ME9BM2dOIPFtTwtzZ6JOjnWV4LFVcZIoOEIBjvG/gLx52rD4dMZAMyEMLu0Q/p
N93aWg6oicbY2jMX8vBQvp2tI00pK20qHI1QQ3CbzfMC7Ftaayt2HpX/6heo8EqN
Hjfv5vlMMlto1/ewz1v6///2o7bf4AsBytdGS7UzCMEo/vsTGqzJ1rdguwLzPqxZ
gaS6X1ZaByoPgJga7YuRFOossUuWJo89zp+OOVocTrhe7kwjTFU1kLJOhp3N5Y/U
5jrqYkckx+RmQpeeMsP5zgnYkmwf/VTiow4Rg7P8r4xnOs/gN0zvhhPmez+Cw3dL
1mfkmJc5+ty3tWLQ2GBMsljQxj2hOdNU+o9pqpzAU4HGRKPj2I6pp7bNYfAdYrgI
aZg9k+VoGzX/LLBKa4KJlmpQt1VGT4xlsm4FgGtQyvUGRzi5XZJpHhl224cqhnzI
EKByjIAnI0XF2SveAojyb6UCwQHVBmc6Ag+5WE/qXKtby6j6wVdO/6tRmCzcm5Gz
YJ2qiDC47a1P1zCi3X3uPUwTbkmvcit90QbRHrEfe/CFbpU8rQH2LSNnylBTIpPW
FP4ikzZV/qXUSEtC2ymNYBLObKWv8YP6mbxIbZsgEotFkGr7bPLVt0Rn77Bj/HNC
Hileuxa/XisY5R5zZ10lNDY0VoBkVXVoy+8mYoVlmSYeXi0lFc+ldMn8TkDiHFZw
ueTMkUniGdrXjZfbLu5gVl/HeE86NG6S/aqRMal7AqPQs6aRZhTcvqG1DIKeHUnL
/4/OP8OKPA73+c+NfDuoA4d7loDujQ/QeBnVBEzj/hcFzS3r4AWNplq4Q76f5F/z
Wzau4TX/Q2MPAeAfZfTaIGvJqqiameJVpgfDvFrPxjkztVeegLNjcbQuNVTUgTQb
6Fa4m0cIEp5+Sjf53vw9WZ3x1dkGYVOYgM9/8eP5dZw7fdXDqmaAt6c7EhjtxYRS
0VEnOjOwjp+ngozRHckpKe+a5zWXmr6zs/KWvC8Hj7lcKJWxt82+DKCq+Ev/y7pn
cEhCnJPiljEgVX6I0TPKiMF8IesVD0W+cjTl/6Vmkr/dN1oZlQ8jmlLQlX2CTu36
zQzKQCowVHP3pxFlfWa7SiIJJS0Snc3mBA8V3yrPQLfI8FCVcoXQW4y68ZNL5Xsf
DTPplyipquT8jbV9LOzyim+LNr/7aPrqSHv7r7JAcbB3Q598IWS6lAlIKKVDCKKV
mhAtyou902lewtRQGKBgT1MGsj5vreMPFwlCa+imMmOcwflfvDH8ktcvWfvDk1KE
zQ1MObuqpnmUQ830RyRM4X/McxV7tn5EW5rUC0mLDNrBBjrZg/p4wF3ywoH7VS/7
Iuv+d4KIiIQnPPDEAeTJYgHke349BJ5TCmtS3vZb3ZM/V0N27OfppTavJct1vlI3
jpIKUeUtA3mc1zIa79fuVUZEtnhyld1p16FSScTs20CpsPvc0gSoCgVwsLY5cane
verIAgLTNqu5R9zWm6i/yhWFBTW5PMNxj8VG2PJTf8C7ZOiNrS5XUv1BtjuXILdO
4jraJmz0ErKIEr8HJP9is7S1DyTBkR4nqW3fUwOtb6IFPknRG6ovSgsuf5Cgzmao
gOlyLoXbwY7xaR2hgtPDyknvuoyC2bLQwmQq+NkjXNQcPYB7k+nMH9ESk8cZwCHW
Lv3lnsAFDxFtJitI9kQDoNaGjPlFfwTKDsZ5RKRfWyrueGZdXaSYPBuZzSlf9Z2A
GXxFN+Ww1ZXg+7xzhfiurBPIKhzTLrjM0sREMDXjqMmO5p5KVYnJ1xYb7iuxLHEb
EXERylU8J47leuAGxUGViGAp8e1BAv0+61B/K5t0Y8M4gK8T4HRHagKs9bXkEhE3
PS2nTrAToW4QbexXiVZQ7ZZWSY0Fnyicm7SAMWRabm9lzj+bIRkj8VtFSfnX7+ik
2Zkr6n22VTqBfvjxujYQvJK+v3W7mWsyORwI9GA3MJJXxEAsDXXUIxgR7fHk3bAa
QXdTUJwOt0VAKlyes2s8/Nfn0VfMkqToKJPT6yIyx9nznXoGNUvFDMfxz/iEwaF8
dP9IEiFXfonmUBIWBRxqyzqvs4Bv0KknzQJK0uBWGaEjyvqnypp9W1wtEa/WO6SK
0t1LYYa/+QrN3P6z3kcoL+i383hklw+n0m2bRYzMXwdfPq7A7yRArGJeKOksnT5v
k59C5ud9gHt5p0EjQm4X5Ag7IL8+cbAjndUDdJrloKlf46xDl+xf0p4PV74acRIF
NR5851wshgAssrfOSkaoHQtVSl/lG9iB9t0bzCKYon0atJZ4JKjqwLLdynLxA3jD
z1JUYJmNWqr6SZrsGZ8t2F0Ga37LZPZJ2OVBZP0iStx48y0HCYgoHgsYqDX/t/Zf
aVX0zaFvsqYkb6HwCR4My3fqN6zrI9CDXGBDziE0W/d7W1mHbRgq5+6ZI5CvPkBQ
CHN1+zKVIdx0K23ewOAY9PCvrw6/hcrF1qeWapQzQiv9mdvUQ9fnP2XDQMpDtifi
dHayMrn4gTtNqpbNR1FIlXjRn9d5pkgK8pwBNnGFSgY7EobXe+uduFIGW6RTBM6c
vHIbdJtsHmuVXmweSzMK69FOszQqy9xf3T/S/J840nEpKu2jHAtU7wj6PIRiCh/g
eRU3T03fWuU0LsNkiXHsLF+eHrEhIcNnO9B55/RhKVbNqF3BWMqSvzYFm1KH+zJ+
7x1cOy/Aka4UVGBD4sR2Ibv86KxpzplZ9QUBRMnjFjAWVfmp2A3zI4G86wRWiXRH
WUUSopw80UyyIa+8mx9YqdyR8HSjiFSAwk8TLcAIyAhzKT8gaaUg1tcdmsMT4fXE
+okIYJ4ncHYhN+0xhyes7NQP3XDxJugbqb5GtViglYzVIVlaAZr/V4cVsoOUCpVO
sSYgtC0KhO+SsYP1uXOAb+m/J0itVhPdWXAcZSKyUsW6ZX9XqeHdQ3p93Vi6rrRz
qzhRq7BdxBqNmjB6UZAT83YZimXxw/aCmj7aKUlY67Xd3i3EWIMOpClWNKWltVhm
zggxttA2jrgip931ehVMULzgBEL/7pRdj1ZNPWxC4EYMjXGaoqirfUhqSr3qPX6/
uTIYtUL+v89dpF/wHOLBxyKhnkQJvcM7uyubNOCd5jBVdCXYLXOqBKZqWf0nK87W
ORUXnq+de4GfZS6ojRoIQblCsi6Te7kQqLYgrx7HDKmI9zvC2cDzwMYlVJvvZ/R2
sr732Qktf7pv/JmyQpxmj1BK025qogD6glQ7fps2KZb1PeNGATiVqpNu6UIcBHHS
k2h/6Dk6GzyCOObHo/cG9ubgf0B880G8EwJPVEJRv3yBcHyuO7A7ApUS1ziR0hQK
pY/lR0Pn4ihYo4eth5Sx7cNCXLJg7JtUBLVlxtF4U9F1cqpVX1EzYvcPnAwtMJjd
y9d2MAHg0AWMDqP7qhkdZAobB+TMzcxJkI9qVEUEaX5d2HIbPF1S64AfcvoiLB3m
4jeYYowDFMVVeBbqoWqX/6T0xYZpYTMGBH3r4ueTm1p6BUHJecd3TR+C+Ve0WiLD
0snW52xQMmfM52ZedEWqQoGKK5YJS2nEe7Dg058iDyVOxEYI1wmC7oFF9QD3mqCd
KPEGE8C7EWZvFKz5/dE13Y/tgNLrDmZBIl17YFpw2agD+8T2Z4IV55oDCgsJuI6P
LBzblNyhj7YiQImFRyPp0meK61aV5sjHNNx2HtOcIz1PuAU0QdzAJoX5ZW657p6r
w0iF2KtPiFVC/Iot3vCMHf9J7v+dCpx0DpaschhkZhOCIFKnMIvKy0d7ErNAcrJ1
wEt/pY5gy3IotELMG8Q9A3NKZSsaYfrVbf/BYUfOpl6wJOnTYZkYXqpS76pZAGCW
mWCyxmnTkHMYy3MFYDvWfeNVvcv4VDyAY5L89Cfb1DAfV7jeei/zxq9fFABth+eT
SvcrgiiT3zkes4EO5SLSAYSqLzWc/QY2Nw+/Ja1L/X2SgDuiVgSmMQJrcx0XVKnE
9ccwcj5wdG8I+nYMrQBOs3FibpE0cwtdR3ixSxKpOUgcghJMM8eqbXiW1fPTJTOG
4CHGk8yZbtPdLeuuHjHWL/VaeQwpeJBALGymr2thvosojK+AtJ02pJbEyn4hBc6E
9ue7EpWOgvUu/g0T1xHBwSkcWpvJYwSsoRtU+VSIfpAKtgUEkS2JxS1ZStG72kxZ
jFc4CH/qRhLWY4s1dXr48W3L/2BcgrWIIgzdx+a25X5AE7utQqOdFJoOGPEdiniR
sF6HJfA3R3+IWAz6EvcTSfUtxpsqK9vke+OHMR3cyvFNDl/PXk+mQUWayVf/R5Z2
gJUKRSEqCtHOjCLEVjl9Er+tVqMzefI5VX54JxK9Hmax5BgIr7jnfXxAHelgEqEJ
d91WOwJGz7c/hVdvZQ3WVt3kKF7FDIVxSUc4g9tL7oHvH2yhquP0DBFdp4CiTLMP
hIbEX9IsdJvMQcdjejhEq05z4+h0BXKqWYTCQNo0i8f8J/eQbBtel3UCitz33tx6
KGIFVwrClZacavbKL1gZPERDxJsRD7I4N04kATEjdnVLxW8nwD+BtH3jrDT8UTQC
KOxTY6KMjukB56BaWn+Q85uj8Qi6dVu9DFw3gD0lAOyBgwE4u4fzCBJTyzQ1o6Mc
VsOTILQtXgKG0ixr4RMdYyf+FwiANBBPTXzPu8Is0Uw2JldtPfI4vFtD35yc0tgy
+dnpoTxO7OMgRoY5lwj9t6+vJM/LnV1T1ExyYhP8zl2ZNRNBWLLmLf2lISrrDzLS
m19+fDdtYEbw8sW/angPvyhjilsJJOxHN+a9cau8ZaYKrpLkF3U+8VlQc4ousZX1
xpziaRHfd/uvUChUFao8OLDM+bn41Hu1iRnqLz+XOXS+BZ8iWa3JZQjqWgKmrKPb
rgR3JarB4RY18enNAOmKu4Afqbz3H2H7cbmXQDjrT4gsy0QNHvWP9at2Uy9/xpP3
OTH2Xg1lbAgHD0twvlgv8kAibleruhxOzd0KVjuDYXBIEpF9qAM+9OUqsqim0E9F
Hr/oAVUHUsZjuig5HwNKjArVFXq+v+F3FUEwaXjXXJDuR03Z2nclbxA6oC0PtsoC
zEWxAI69vCVpXE/f55xuy/14yjtN82RhDI6wJHy42l/9JCj85LEmVGIKJIw104BS
nw/M03cYVdi0AqUHqQAsv4UrL+OhyOcpx2XQxd4vCepVdWN9rSIgRYCddUW7Sas1
NjUMFNLOaBPIzsJhplr/pDKcqMzOW07PMP2AxXr+IFgYV2xFPTR70EmuP7LmsZIa
uMUiNgk+sehDb+hKXDv36qOp3SZOo4b6CViwcM/BGjG0PQyeVYzvhLpNjkrv5nsc
q4o3iTCxPzGJYKnS7DoZ359r3dwi6ZJqH7FCo5PBiNSVzjJtX67uHZMWbzb/wUJY
HBQ7bAoE1aYXXf6J+aYSjIxf08xEc2soiZFw1TKmuFX3L6wz4Q/VmRcx9HWK7bW4
5iU7NUBMDljaT2FkLvwXbudllRf92Ka96QYBTbRM5HbVwJe2XR41Ew334WcUHd/i
LWI/T0ZmSL+hvLe2l8/8nKv+EG+5XNTw0ljsjkcE86xNNVB+BRfRltGeHNHnKykf
O5jmnpVZknsHhDWvI0Y+5LuapBCjPvkVgxbav2GWOqCmpSbmpHOs8lWrwYcocv5H
YrWprtSfvacfusapq6wxdbNMx/R2Ake4F5ObUGv+tkWyLUJuUp+zlgdDTgkrh7Kh
83pJJTlAzo/0YqBG8wlB2Q5LO+GgkfeecEqKY3vZFsyPwSLYj5MgGP84chsoNuzm
ykwRdOMTaptqdUE171eHF1+PzSmPjiLUfUMGlzmUpQNK5kgQFU02qMc8Boy4ahcj
y0WtryXQxnipVUpPGlWBpUaS1lbW2rJTT/UWCzlnyGlsGztaoIXSOUmVGJGE5u6/
wMUONWfXiQvpE/tT+vBVUrBl9idTpEqRfwyHrNRbIEYHEMDtCBtH+BEk/I5gvjnK
l4IaTIlYGdRNwHBeUQGpW/efYZGIyS6SH/HNyiS7Obf2p0a8/+X+LLsMhXgxbCKD
26ENOZwHsf4++nqAHAgsy4WAQUpSkNQffyYVFvamIsR+eBG3iBDEh0HgEZu/mEqR
xrKtCNAx9Qai08OYCQmQ5LBv+eYACMIIiPjoWqt6EV2amkcJ4loqACd/xeMgxeJ5
hBjLA8enyOH6GB91vI2itR9uGQSmQgf0NgsR/Z5wxMZwSQDHOZykmIkbBBb9pEHS
Ap18n02/nCq3dk2TqVAMvW29EH5o68SLAIZj0RQuu8qMNGI+mP3wzclds1t9Xe4F
EGrFgbhZrXuLdEPFdEKqqqACmDMjwZXmmsROVOHLfIaPT9UPlj6d6PwKAxhemNac
l2laqBhDt1Bcxpku6muvIOW0rxxnvtWYQrVTtHRu1JQgnj/p0jfj8s8T9qTURx5O
E9t4CYa4qYFvPCklrUmZXjtaSF1yRK45ZQ7JT72b59wtT5J9ymFL+PMMxc3rNl7e
Qlst/XjZYcMeDyOKm+xn4NFksdBXF0bDCRIJSCJuPohbL4SMAGC5hvdEnCbN7lBd
GZ2cGtryCTR14eS+cHR5rDDvOaKSyWq8mioWdv8FwpK4PiqJhs/RQbgGsTrTJqLU
1EwFawqQDZu8fudFSD8C2lEu5NG8VDmve7qurU8PyvduzMkbr248zOYNcW6u45bI
zzPCdIiNiBYgMPe3Q/E+s1GQLKOollwz5vxKybcFVoYMBR8OGaH1SoOAGUIm/mel
twFzkqft5XHTTTCynOnY+y8+ubRJd8zf9+5bT67ylIKDfto0+HZh6+mCIJVhoU6L
sMzUYVoW3P/W4ezkJIEFv8imb/8y/rJk2nY9ibGHkJtKv6PXqsPa2yd50FM2mdhd
niowq3BnzXCnwiGu2ogF31gEjXnp2G1OohHXA+Mwxw4dKPdAbL+vNCTbRIJo0AZ/
suFV68mJApJcx64Syz/iTRmD/wMy1aC8rX+k83RltO+pwKDz8tWoONbzxGm1Uf08
zpOezq0SK+A17BvhX6lBImpbVRdT9Mitt2pQnEPQRQCcwk6bRGhbHPnqtTys49zC
9kiT1YS/2hsSsB3dmTe72qxF8RWPZv8C6I/uElhe8EmDuKFzDE5Eckhot8dZeTR/
vvIJe6vgFDnJrjeVTQn0XFVChRSpMTSm3Cle6v8kZPQB4ULXhPgb/oMQgcRmYxNY
ONhROaplAgXpaPu72QLunAaesgbvx8WRYXbAXtTNUgQWenIpc/5DwUy7zQX21Xj9
Q5OBfsJzd0uRAs47IMNEyvdqxNWFVaXECBXUIYj8d6q2yWu1uAC6pf/3zRv+C/HH
26BftR5W0sORm86q5fDpn+3N9y/ZcLsaj+iqj1gu5XpSJojhNhPBmwQoTkeVf5c0
n15FhEgYf1UQy2GYt7QLzwxnC7lhav8wylquGsZI1Ht+6rHrnIYOawC0HMLcWPFF
j1uw3JqP+9TgsALxRp58Ztvtj1cY7PMidQQr0qrJEAKB+xPZRPoUjpjvUHOqgErt
rY9F7BTY4HGqxrXVbA3K0f9HhS20EXDqVEw4YzInpcxgTLFJiNZ3JkNnrdhDU2nC
gB0SKQXQXgh76FHtuJFV2a3FQAjbq7bh6Z79YPQpTS+7/NHsEDTc4Xo6XfFgzOSe
ncafaZG1xwMxdmewL5Taa8TqHn95fkvakfZsnAHy5XduWY+2VMO2j1jg1IG0q0T0
TwLcIcm5+F8HVkOzwkSW0L7pBc86lK4/gFrSM1Qj1+RYkYuPciH9fyyvozqBA/tP
WrXlCcATXyk+SDwOdr6V733PPMCenU0Z0dRp1iLGSzB2gcqM1KTrHIJB7bYh0zVp
w9PoDGNYy7pd1x5dsJJEGSpkUOFO4H0YTTLCoUmQw6OiNEztjdRnE5fHm/vfOm3I
PwcInMdsvX00LHpW/5KWPqBj9+5eboNtHGV7tIKXiYswrkjszP+lWjas1eBbyRxt
kKBWCBPSBeg04hnf65hdCMPybwzbKX1n3/xF+JPUC33T89iM2isoDLGXxLLXkmUe
32dEMsU3NQjDMMLPqLHuUuI+brybqd3l23b8gZ2WmMvBM2lpp2Jci/Dl1/7203I0
gYBTMQXbCLD8Mkj09tVXZ3uHZgf/qYOInx48+nhIigboSDQNfmnerHxfxffKrkfO
s4CXCy6o0p9mcUX3/qvX9VZUXRLoGjL8VmuK4/yDpxj8yVi7eUhDzxd9g3acaQhH
clVlzxo6k1LZZGZD2bKoTaa9QRKPShm7e/sAvf1Db/8JZXtXHJRdyIKvRieG4owG
5SR4PUQrFZai+tWVjP6avuhudUO3nE5ZtBFaWDCt/dPiALD7je1aNGLFOgOWHlx9
jl+N+F5ejUCuXl14qMC5cVCQGH8fPVF4KnqIrJ518hceUtlU6sIaQBpV3s+GbKQj
pM4kN0LT4ww5O3agrgBAkWwgGREgMJ+uc7nw3BMKZ2NAJx7BW8tUBfDZ4RHHbUtM
XFowVdFdlcgFKGhbkky05qHXvwTEn0MJbnxMNWYKSYmTBSN7lIP5TraljJO1R4YG
8953mADAHsB7jWy7Rgj8R1x23KGuG3FVJGhkSWQd1GrWICkQ71ZuzjNVm+V5mMeI
5N9dvE++pylUDvN9D3uY8Q0qobJx4siVqDArzy1s+OwJnCuO7mVQcwQ2uDopz5MY
xaqiNmGzDRHf/u3fMPx81czCrS2gaOHFyoBfaPLif0xatbSVswI8Qw+qwtn5MeHI
NOcm9Lb/r0Tp7igrHsncELFRmBTTSWRwstMl7Jy9iBYbZgZISYWL4Hp50piKr4Kd
I+OibTgwI4m9TeX0cWALMgwzme3L6S0maLaQcy5tBpRq9TAp/D/QZ0mcryPPOk8j
amNfXFmxlYZ8fMmbCygUAPbO/5xXCL6lCk39MmoFhAMFgVtqsDyS25HdkX5uE+dA
Ud4nmDQwAz1D4ZH7+DRoW9GJFNeUfcapyln71/uCBhPKkLpORYjSdUaFIIh++umb
C62km4+B6dIFjZohm/bzKAr9ofcPeu/cflYwdSA0mMFsHW/Fu0aRVAQSgEViyyTW
4iw09siYa0kpqdWpChkMrFOuxD02fdd/uZ8B8FhrU/52Snk0ketANR5znWwYhhT8
hOIIKv8t3qCdXTrh4YptLInFjVcDfm3P5bWChquR6a6M0YL0L5dQD9F11twm0O66
N3qgbP0hoYuZXwazpOJvG/KZCZNkidXN4dQ39oqdtb+ivOeeXp9+EKAlgjC68X/e
FVsL0F8rhGZ03rLFwddGdcyP67dsddmG9LTCisq4NRF19JrqO+kRxN+WZUWva300
9T4MI6/nmQZOcoFPqYvsgLcjXnQkhv4GDmU1/h9mX7zw5xUuUxXMnd1JICc6ThaZ
nffjtaeapX5YmEqwLPIl4PBa/4TJWpWugSValSBTqfxCvLvD15l9d/qQGRglL9a0
qJw9dRqShxqYO8NHzRlq/16wJ//1pgN8fs6NSuH6fcv2xnBfkhfqlynGgsa8xdqZ
Zh9Tct9mK9+ubb3GcKe+yxJ0GmRvb/XK4DU45gCazk7f+CZ67vRICHs6t/4Z7pcZ
xNeHUM3WsDWaErzfyMNXs1ZkFFeOiNNI7/ahKCYXEVLrDGM/JgLvdUW+UcSbZ/51
0fQwKnhD8KrdJ2OtBdkH7E0d+0YZFwu8fpOLheUoGpDXNQx/bqox04scxJu+aujC
68w7hlgodGlyMLE0u0JIi4I5rcQYTD5DRFd8FmIFpd6hOWXpbCpX6wX6fxA0+kLy
aTKdUjItrgBu/tkeFMnRz1BYrClQC989yW0bmTlU7FTYmmo2ynDb3aBHUjgK/HlA
XQ/UFNpL5vOkMPVLxoNby0G8BraO1FW7lae0uy3DoDO8Y1PTwRk1nKE7V+yXPzAf
y77CU14k9TtywWbg03mFUn9gmhVWFKzdEiYJAB8/4kz0/qiwcvecpZ5LdxveVAzr
mpyuoVsKpNQU2V3ZMGQ6IM41SKW+arr4+o3blEkE+of5hNwWcxrLdbTvI1MhIKnz
Zw617Af2bYGnJkSvbNQUrakqAhlBiKZpioXYJXXoRjYMXwSDNXEU6Ei2c+uXhXnL
D9OzScymyhHIX5mz0ftwJscTHxTEIH7NV0xP1+WyJpr/klbHeHQ27nzQ5klKYx6w
ZT82/iHVD614pfK8ULV0XoDi4lnR3OyIrr0R9KBfP+3CeucIBiErDsE91pP0iwXc
0mXfhTp7kIX3BiLJ1NkZlMUMIx6l68rIRc0C7gQxq0AsibhfzUJTTpBAG4pWi176
cqSQzsL6Ic8LH+ThSxPImi1SSol+fBPA09+9kWTm/gmLxV7TQ+CljXhOFskuP5E+
zoycSzIv61yXI2UdRvzryhQzLoiU33F/a7iF20S37w846PHFzq0dd5zUGRh+eQrj
vRduq7AbecECDXD5l5e0ATOXl6QW13CWv34UFkNl/KzWSwl8JD13fIm+4Y3P2tu4
2nXrEeVMzzH/h6uEkh2mN1EbTkFqEfApqquArPV8HKVawghrIdANIvrZELP/Jius
8MfKYjBzxs/pNRCNMYCll3IiHhmAbRr9fpFhcjm+xhF3TYhRpvusDEWEibqEr79D
vi0MkukUptvVhLMl3qGzAEfdTTtFL39blDEG7ACetYqPbfCWtTq1v/P1yF2otqGW
4rTsCSY4SftJ5ksdIkyXCtMUtAp3ZNJVC2RWxjCrj00TARn14P74qt5uZvyi9cuz
72uC7gpviJd/TYZ9ieCsZvbfo/nQY5hwWYUBlrnJXm4pU/CsqRxigH0KNVO8h5i6
RuSWr8E/Sx6EYASuRwlE7EW/WmJAebNrGeG4BMdVpRhGCjHH7ctDhbpxa8eAhfCx
+o9ZFKZYf11Py9yW+4AJ1T4e3rOeNqEwh5oYuywLxQDDeOs5doLPDleGFjve74aa
Icl1nSZRYB6GasaW3Tj5vDawFmmuRqcNelBJl8iR9L6Tlv0mkpAHfMRPskS3zPG+
u9fINeU6kRiOR1juI5npqR8S5lUbGY888me/nXcVn2cjCeVM/Vl/c6kPfm8V25ZQ
O4sGCFNSIgvSpSzGBKCcxhrVacUqjoKpj+Dyvjei8Wdq+vL27/pPR4ZL1XH70QBi
hKvvmajja2Zp2Oc9xFr+xybbXfgaZr/BFElTyngNehfFiWuEA0Ox96JTEiyB9mdS
5DHGfIJbcqTSpy1umrPDszHzpHY1XLodRc+ZE1lqRLQyOkuJh2qWx8PigBI1fZ6V
v03q+5b90R4fb/pQjd9vMcfrJgnO1+tl+95nYW2+lyXkyJTiBhL6Sr+2uhH8ubYI
reUakCKBcsZ1iSW5hc9w9kh7Vm300D9KZ6on6c5MkPQmHvKlKlWJbzBks7n8jWhM
sNfAzLslEXVMHllRQxeVnuxtmbMBxpNQ4wJT6EcOK+FCRzLpadH5DX5MffRV5WI3
Lu0M9DISJRcoQ1iWR8sizJYIzhAajSpLqfpRDyoqWyqTcJDUyMi513v/IH2MUIh7
K6osiWycIvY69OYhSZQ2v3qdmISr0gQipeta6DVd2uYa13s0U96qhGA0dGWZW2SM
WTkrLVaW60jZCNah/OAm+5vpL0VBQxWlSfSxWuHs9UXekX1s5+cP4e59cKEfBMPG
RXvJebbfpzm1E2T747sY71CSfMb5+dY+fBXosZFdavqSQ0TAOyRJ+wN+0y3uaBji
498yy8G6E+ykWpB2jK9gQNblFgzwDV1+Zh+8x9ji656016KAWDEw8trUSClQDFX0
f8EhdBW68WO9m0zBHI3S+hRnl1ZNHRw2zZFNbczIGhakGKgBCjt7VOJ/PyPpmxcG
bLXhDXe7HTBNyjZWaSupbLf8bQ0jb0F/ef1TqPhffXo6BQNkqIy+nh9rk+mXnM+s
8rbZvl2MDeLXgvyZxSN/f6uTXyvvaDCudOZcCcHklB92Y3Hv+LUjTK/U7NPNpaXa
1hQJu4VBV4s/FfrNc1ZDWi737BPMCaYroD/oCpThY69Cn94tp/Dh1BHhbOZwyvIX
1PkJAdW25qfvcOdMVgW/93FL8EJULO5VmbgZBpmoemU1D40Os3OfimCl8k8mLbwr
QgW4i8f3iAtpm9MeVaTOR1Wc3zKG0svhZEQJxFVsptgrVpGsM4csvvx7eMgxR8U3
oJqItE+14sZARn5rxiBnJIT7nSYwkPbb8ZrqfGu3uMke1p3cA+v5P6jxAnPj1oRJ
PcxZH4WW0uXItgQFSmdi+KgoTrIGgxyPbobm0mDuJeb0urDDOZ/b4bRieALNtZdx
ZsclGOOk8uAkTfx4ZH8AqGyiZcvU8olPJf3SgoUw/WgwMs5X290VkuOAHG8RCfN1
bjVIYjZn4O2JkybnT6RAbAOk7rw9AVokxOH8zrLgxOYaIvtiIjz+CJRLlBUqMkzN
Hrsz4WrGjihbSj+qkMzX2h1DKVsNbul4m+nPDQ0WJ7ornOpI2ED8oIAXNQfd+0Ct
3S2V02uY4iilgrReNP+PQNvjp8Y3wn5CTJppcCJkIHfXyiqr3BCEqYlFbXPcfJUQ
StJw7h2Cqmm+7uhTWpvQ23dddU088qciT2I4SjRfQfq2qQI4IIzTeZA7YpeLR2GU
4zPnAbW7ITYz0vOChJFKQSXbmLUoN5QXri1G6hR/xYX2hfaFWZiClv97vhsvzwWk
/JciEtuZvUwo+EBAJBGTw+Jm9C1TqtYc/4HylnUnvZFTyhMTXrFLibwqJP+LN2Wi
OTtu/l5SiWDdtkpX6gzG3kbrZ8GwCxq3XMoKzG7zZKtAM0pS1p+y7ksNuruZHgxN
wooZuSOV6Og9kSkLDCXQ27cZMt8A4Q/wjJMk3JtW9OTW5qdDxl/g3jtjxdF4407t
bUadMsT5ySLuQYQynll+GHc7MEGP+Jrhad3SKA2zNFDjNYiRnbImukbFyfQUbUuS
tuCgD/KWmg3ZLHg//Jud6csr09ik9qmus3KI4zR1N5EKYaNgZynIwe1EwR6X6jsW
jaz+xaDfJJ8IzmdYjyQ7KL96WLGqsTh/fMXshhNzJmeAudHRzm7hJ0KvXkzbVsnX
Menvvy0FYlmS6SkCFBtZTaaR6CJQGWkCpqT6dE7SziOLzwcVWK3zI1zMladvW9Q7
moXm+N2FJ+Z9IixOEjFcN32WEpSC3/i9j5qpW/1kQU/HpUT+XDNVo9EPcvkENWqw
A92egAX5BqRqAMhbfyENJ5wVW4UMc/H9t7O0oc9EqNJwWVGwzv2TxLz0KxbQgWaS
ofmBfBcvfxJJLsFRmASbCeEo68iK599jRTg3kRtug+Gzv2aQR4SDKzmQZJwdB/0x
wASYq30L5KmXET5hAs5VEJ4gnhaYmYZOel4TL/6ip/yzruzUTan7na24xxje7bJW
LWhj3E9+/Igh34IcJHspOs0hsCLdg51BC84BkJVMM/H+eMN+Rgx1G0i5a5sjM3mf
m2P0nM+UcvvY4kRnz+AEJWATecxtp/1F/bhXIC/4OEVt0XxRCrc3zbqXsOVSd0WA
E0ywpisrShooEFIsnnBXKy1gcFn5as/yffAg+n8Mhz0MBNwON7aDF7KYAQi1DAen
fve7Qnb/8podEuU5HTuYUZ+zvhNaYgSM9NsidDci7/87IBsGxeDAn15mTlqi+u6H
sYzFmUiAWRlRSo2TVJLYshm7E6S8gATGjwEMPeea/hVvbET7wijPA+5IJsKp1Tyl
HqRE/u1xgzBZ0s9zQYi0pRAJj/iP4Wp6owXDPdsmD2e9EwL1z7wly91CVbIdycNH
+Yyk2IAu+/7NcXnFcECfT6GZX6NXrkdedVZs3624Xhna+dsLzqeuGZDg67oHJyaV
H087BSy1UHx4AHJmn6m57xAmGzh+nfxKJS0CP/18r7tYXnkJzWsu7NSKSeEce6XI
mAetZ/dQD6L3EdIkVDGT8H1/1ZIUbneyoC6axTtSts7jf7gMzhVQri3BbNeRsNLY
p6eHAZQWQCfyybdptO9FfQ7/bvkvropc+LOE8NHtMysq8jU7LAQcMa6Z22/3vh1x
7FsY9KuMqpBWi/7+VT5p3ACXIerrxsy9cuDc5YmGJFMJ+7/ghbaIeU1pASdQuQgM
bSmkqOyVlyWe9QwYcu1TMtY9iSMIEkxqQYsMVUV7HOML8nVR+AZbtvK+qU9X2neS
sjkA1bfXRfQjXCUK4X8wdzcWOcEolcIq1OXZX+xBruLR0e4fffzkSlBpGW1kJN+5
lZ3g+8iWyoX1cKKKTdMta0H8biVSn7Td2o09rAh2hSbgMNqOF7qO7cFp0qGIdYFl
PfCXIepk2EL42iZt+D/8kjHsTFA4z8Yj3Q6xqmU/3Yggq/QOeiNUdoutc72c7/ff
ICheIDhZtYRNtFZGwnVkIQi9NdSipQ4aX/L9OnMWWv4xR9/DC2lJVTVYyMCPLZXT
jn3dZwyg2OnRPAECqdraIciWRSWCKt6l5MsJpur66Jaizsf5ctout21byJePAM1J
S4zJRcOGmsRVloHATfwU7a1s+myQM7a6p3wj1JPjkD4ucTsJfwOhHSJjk309jAYT
Lxjg3h1JMRVE33ryRk7aRj4VKj45fzJfPcJ6fwEsCMJRQom986PbxH+N3v8KdhMd
rt01zcWxV5H1Rnaha6qXi92Dz8kAakrTHdUqv12f/7S9PiHE1pqPND0LDMhwqBva
hQgzEEwfCTUs6n57SYIKjhihN3mRnuftZu+L5Il1sfxaXmBBRKZmyhx+JFeYUO5w
NVy+REBD9U9qefYNsXYpFeJfHA4w93YNVW1s8pf8WFvSqHilFSUvH116w0Vk4Amw
Bkn+PzSIe+MAdw/GfXzasrV8fl0s2vUKIaRBWTjaDI1bt6VzycjlSEez/MIVLg2J
vGlGrlulKH6phTBhA0W8PuFpKK4Bl+Z2WM2K6nPTyX/K4PRXSq855aM208PM2ULo
SSdyCeENls2GLj+NL1LsztZH4VlJzDewrsviy6cqgigiQgJKFqMgiG0dfHTf58Hr
qCRWIfMAeFA1AydZMjI38kKc24tz9EtBqL7rcRe1NX/6eUo8+UOO3AsBn0C5H3TJ
ducLXaMXYqse6wwwlOWGvEPPw0OsITHgeKoDdfOar5Lbxv73w7vf3EFtB1zboxiW
ZwdWOCq74EIOnn7uwxTG3wiv7zs5XZAxYh5+pPzDllQcwT/pSsdJ0mYeeHl/vZW1
ofuuE9Zi6pz9tnQbjPQTFW62pDgu7kuvlUObqVeuaqchBgC0kG8GR+lHtwmeArBX
8NfQgInosYyJLCIPbJp1EyGibTTPOOQ2PXUUM+2ePmoQs3i8Cog1GcTU3tmFaRAx
Ge1g35Nd0xj+/T9odml5hxiLZ8gIWU3llrqD/sw7rKWMl5Wushmb9b9nPu31Cfp2
2cjK+omhJDx7Vq5I+tGaMmee2ie2fQHdPeE1KpJjYNKEW8bXbVlse1UnotxtbJfM
O98mV+HkpvrPbXvCAqYFklCeJY1lgT2IIO91uCvnUJRIr6VO2YSACv+2IO7Em7bl
UCvFqOd0ueT+KsBOZOS3q3A4v2b9HrW3y6YG8g2qiS3ju97ily2vc4iezvbs/8ZR
CAt0zm50XgsVoUG81ABDibIxvHUwvkmhRv4Z1k1Usy2WEAn/NLVjAGIFkI8pqgQb
ik9QuG9u2nmDHcmZ+KihGVwcp6AQhA1iOrWBaVer68LAwcnRiibM8PlRMBkzDYgd
5Eg3g0dClqKJziHGRwxQmQadP8+R91aqCjpSHIv1wiO7Yp00RxB3fVu26eRXVVZL
ILj6aR/LqkD5WyvrrFbCi1i6mqJz7uxKb38HEhGQhMJN3gG8STKGddfcGZgCjfp8
O5+zW/gbwHa2L0oUwfBeCWGFgxLH6TDp7JbYte5WsggMad5+JbfEz02JWGA0jbkm
TRZIhsTM7xPkWP1A3IppSQXCR93yVJDOZ5VXZ0Y/PJIEiic6WqI3sciNRHAs0tSA
YCvaqWivIq7mVus6snJZnZrEoQCMVZNRlxULdqOXIqODVIZHRXfqypzVhTAUqLID
2deeaBoI9zjG8i5v7OcOpDd1ZA76PwG4tT4hyVOBoVI89l4l3kDfhxakuqEWcIFH
g8koxAIT+uwXBWwcA1/jS6IBZ5Lh7NXBJoeo1XK9EoLHiMAwr2a/dt2yBj0CSrwg
Mm4kVsTHQbtYLYiixAWVMJxNkf5mHUpf90Podpdc8BraMqlTFcZJsqgA8AFz5mSG
dlLwOfOXQQmQVuJf1Mk4rohKFT5lHW5fIpmtqVR30frfOB2P5HwH41YxNGuPc/Pp
MEMNyXMBY2VuwsR+zD9LvTnUGxTqEWNopP77kv+E0kKbC+a/2uXYD1LhBKlGDxia
+7KbvDqqS2v4sq9JG1mzVN574qzD2s4PwwZK2KOr8ig90dqwklGq0X0Wae+WZxzo
pBX6+s8KEuEk+nIT7K+zm9Tkx+1NrRAtMvQaf5rlNmoF726srOF8QCcSaUxdei9C
NHNkAcxC0xFVBDqBUNyBQWVc0/rftXUMIBnEoWk1xVqcgxEJ1L6ZM/Q5cIPSPoML
qhIxAuBZ3JPMjIEgd3OSN2/X3kPXkV+6wAq/RSrB8Pe9DQY9dMuHTaJeMwvCIfhZ
w88KdLj/BKdfcvP4vOkcbnaAQtT+tg+MESQA1TdUpS3L+Q4jvdtCfs3nnYjSeXsv
CTBv5RfSs64BhbpCtTlLHUbjcYfM9rVkMcZLww7uIXn2mUDOGPL2chCsuo0jhgJC
G6r6sr+MABb7GNMjQD07vjaixyCndJLVuHQz/04bW71b9AIJ2ApIJLAn9nN/PgwZ
isY5zfjEbhAvsydEnl/N20QYGmhMUFVekfFzjxnUM0MDPf91Uo5JqCoo24HB+Bpw
UfmJQHrHDEvy5hGnFfEyD3NOgsSbv/PInyLRjM4pADJr5G59quNMS+BsI0sXd2IQ
tgSxovBJQh9c3hewJw8huBmIwj4naKh16LFPLU2a53Wfr+bV0fTgSR+vYy25tg9+
aXJofFvgvvKCzoYkEIcgNd9KiS3IloiL8zpke8zfy0ohugcA4Q6O/libMoAA8mXH
Ajalpxo/EQXNmq6cnafq3A8QzxHDuczq76P7Lznt1scbK0FcAGNZAmqDKCm1TF2I
ojhIWEIwtsb4Ff2Ci14V7XPJXE/qe/aLDcRhTYrovvXFUzKOCrtdOsGyBkB2fzjY
OvnH6qrlwYOEe3o6DHUpla0SfsjwEjO0QVZ/DguRrDvnXKhsFc8I8QUPC0UsFfbe
7n+ld8pRAbQ6WDPAYP1z7yO7xwPCn/Am3sfVwTNbqnIeGZR8OD1PpFC11m6CRqWo
G9mpfny04GLwpw9h4mz6xoSdXpKx8EV+xIEEQItIwS0fgdJxfxbEv3C9xo348qqH
MV3pN2JPSeNIuAu88FhBbqG6F5W9mLL+H4bvAAvZIWgjyk0he2SnEW1MVnd36rRP
eHtUExSBqF6s8xkFg96acL4AS9mxBiyIA1RrZXln0uS1aKbR7hmLE/1pInmvjdnV
JMu5T7FMeTG92H5QwlFW+9921IaNiwlXM7rP6bIRPmNYOUiMslNolozCSpBaXjZn
10yytY80VB6p5VaAi2Bm5I2xVOYfvpwD3Q8IUN954Vnz0pn4MduvU/3Iq0AaFadO
T8kWhxV4sCCVv0GzQ6BOtV5iBqhSI89aZKgrnYotjp6FZ7teBGX/pjYFbtTG5FM8
wlxZR9br099Xn4LHh7JkasLIKOwdTuNk23GAIhFxAZ6A0y7ZGpAjsYDrkDSk6uLM
RQhaaaWTDKp+DmIaVKhtHE7fngydsTUdFPYEhl9vOt3LgtZoTP8ZOU3Z5GJ5fyYg
hwa+EtpBaLYf3je8Xy7oRMXRPVn1pDfG5oIaBMAmlPqaxuWfpgW+ZMthCPTdHphp
PDthevx5iaxNRdhbpcS9tmm9UVARaLJUqbaITJZVt3XXWQbC+VO0sor27AKmbohM
vkHhMqsuNKIF7sUACUMlQ6Ocank8AdTn2R/GrdiE/XOkVQ2rV6oGoaBaiWI4tnQJ
AMVXtCnuaSPjLPG9FKcsLcjoi5S+rhqeccDcyVQzdNLNARZjfXESh2NasTELQQrW
uzLGWxPffgLFYNBqDOm+FBa4DnSyspujC7ZrFHO9JO5ruAkvgIubfo6YusWP8848
2R0w7KN91CBpMmCNOlRsLKaJevGj1ZXMx62pklbcpXfg2LKcAA2muy9YbT7ascm0
fQCjRg586EnWq3USxcjacJ/ChgyTwtnhP7k1plogvrIQ8RGQdxbUzxVZB6X33XwR
H/P2btwkDYs49na1cdWxZ8pwERqgomrN3PAGqHZtWb1Aj6FUK0IkxolXPyM10b8S
ogjXTJXkNAoBLIgTEhGqm7mPLxKqCgetGStWZlSS4lB+SznEitVaT/eDhsDOPLmE
sicikvWVRixvBxU3obvdupETX5GsvWZR9lONCgXjB0eK0/+LFglImMsdvsQUFs3w
WIt+ZewkBTwRN/30A8o4ToFD7BK861zju+pSQic1k/YJfBm/Kleh1kRasHMQOYAM
z9AbCPQ2nOsY/HEzU9A02vxXldK8lnmJ05mr6nF6tsAb7K94Im3puFsqcAFw0TCL
8uvb2F4S758CzHytA+HBTIeRmT0MjJrwLusPkG2TLgI0ZQUSPp/UoCdEwtf4Qn4H
h+KLAubAw8VfG2kbzfOJq89QrnHmIlnD/PgFShJND8T3XvWyTwR0ZURjSla8QacM
EOuHh7hW9SqRN8wuu9fMdy8sIui2Yi+h/WMjKW2B8STeg1qW1DoTcPQNDGGLyjHE
5Kuwjyx/ZAiNcIVcx66N7XZmLJwcqrXsoHZN3t9yWJs0DQ6OEp5pPIHsdyJLIq67
sYGFTBfCVWY6FWngbjorjBTIIerU9UCLT6VEAgBwyw44uCgutNQpThEjK3sz/rFU
jGOthVy5MkWN0oNZ+/K8ZlhBFe512Uzsn0I5FnfjWDk+rDtol2Zjgu402GtRKcQy
cUflKWConeWfKf39t5WsVNs4/MqT6gkO6awPC/pmLFDTXmLqKtdjqrHYbA6QupHY
0VGGxB7R8Me1FEHn/b95V1lTnrPqfWPGCxJss/HJf3x3kvR/NVxKUTD84LhFO4bL
aLAPib7iivhvHUbueKXqzY7EOjR1fDWTfaAAt4idYc7wpl+vhH7C7o+IU3D1iemL
tvCOhHFqja3XEKrvxIa4diuXkG6X9w4fICkAW2BOxNTFRb7H69l86cSmxdMIUh2Y
H3I3aWrHgNx1txnT/CbSNxEF6hxhngpl88jQDWYRVZTnIIsuA47PKNtGdKQppe4X
YP5kh5I1DnToog8twM4JzMPLbYlIxQc4oRf+2itVhOpjCRB24QXnInRnSEN3Ujrf
Td/j/oGjsRQG/rq8Ys6nYXf8PgJn8NqJ7D9QOjZtHhL4HSAI2VAKR1uYrVFlFtIv
6T564hluZ2AFEm/GmEitlL3veg84ojZ3PIPJiRwdQryUwM2BkEr+BF7Y4F8NmGuY
XGPrTS6vvJ6e6Ks5qB37SoY0h2XlPOY7knRRypxZ+lCX4BLqTPa9vfXg9rwz4eqz
CtmH6DHxcQqShuDSqizr6KwDLmGdiy1DgBL2cwpcp+OnhMcNJWGqZjO2iiGXFOMv
oatexdZfPbcBxEaJl26UXHynzztVPdB5WXtmEjY6//2IGbqixXLHUT25WRc0ONqX
vr/y466Zt3R48YrEmtNXkRrJLnA6KiYxWLLfYGWTUebjgytF3dLYPg71v/+Q7moI
BmQ82eZbepnnJBGlu4AoZ4VA7EqF3GhdiwJ7k7K8b7Q6cKRw+pGxG3oPzc2XZXNE
UAXNwoQI7STIdPysKFzMNLXqDxhgTJX0m7FedIvrJw21Pn6isE4Fo5ImO5C31Xr2
Kj6LgeduqVs8M0Bq6O6ihVXBLGB8oTR2eHwG0TqFHQiveAYAe3DbnR1el9mJxlaT
nwyfC3hED3Q0cN0mJXSV8ZX4z96fsAovGojZ031XXRBS2mj7uz4EiZcZVnDeKiSL
X2dSOHwqnDNt9Dm22y9c2554fTdaOOzBgcJ9fbP2/K8qGVMUFAkMEVRuSJvxcb90
WjxRkDMjtkLogoMHRLcGYhRiCkGeomkVG7OCXZXugRB6KhDFHTk8RQe4XO2Ky2/8
SwLV3ja/aD1h9LzxJi0a2D81lKg9WpIKhacd2bcGKR0qcCJargmyNs5jfNQhkzZq
q8GH0aiwFqpgzurZDxs1hGGlvDAtizL2x6gJ/itLqPRN/I3PfTXEh+Z+DFE9dsS0
tRhPpFkPs1KBhdZ+hYV55lJL4PwOM3z6yU0xupjTG+UPtlkhW9nNMeFOgRB0/aOP
l9yYxNJoKiW3b+ns1T/x97CJrTcCUKR1fEHiJ06RETxlMEwL6FK6i65WkOsljl0c
DiN8mJON5JZ8y4CmPVFfmPlUN0N/E3+U5UMBfIOCSK9d0UnSK9gLU13z8mcuLywX
LSDuNn1FFFpoV7rsGKXlHNPDpUcmQLfm9NSG+/zj2/hyJiaOPTlCSWf2a1PN0JWi
FX4fJWjBLxH2EDh1WtrBrqMgmmhDxSXYLmU0mhELxz2VbmwYnF+KWQjrQJQ1cFew
Y0E9sc0A7vl6zr6pmRaHRRN/7LPGFpm5z0pQQMPxHG0+QfaI5dvQttrZ0KZFV5Sq
6SVzQUltxjkrVSSpJyhraxjLTV0eeVgSFoOa9k5NLfdanYy/DwTFv+N7pF58/OjO
XTISf0of+zcnkwxvvjagk4jLLRZ/YsXrlDQcTJZDGtjBYzokDBRiWzgA0bavgz7M
Urwl7/apOCF/O8sD3OOH/PGp2sxWnSfzmK1IVy+SgMpnR7kxjbYl0le91W12dzV7
mZI7f/ed8l1DZD0Q7Lha+feU28j7tWinyqzICF07n4NwqJcy1MiLddjLjPgtmVIt
hFRhl+kMthACZNnh9vIAvsVzK4FvvCRm9cs2VAzOTl3NrPyA8PEPNn+H1BHV5z3e
ly8RwasWvUP7626w1XiEoXK0c9uzHgO8DHGfMSE5BRh4lPrI+eKn9CKvikUSCTB+
QbdyXWWL6e+iD5LuiCMfXTQb8jMIFceqY0ALJrEv3Fa/NzqSmkZzZBf+Y+E0mCgu
Quns0Sk7d1db+sKSolBnaqiKwFL01IcpEftDiJhV7qJfGWfv7b6tSfp0fCT4SF0/
e/qL9QX0maFRphsoAGCMPzD3pDiGw23zJB3S/xpPHBRcWvcvdy79siNcAO234wCl
YEuOfIQVAZHBqL26rQchHfiY+YTVe5Bj0UQF5RU7zwwYUSZjSIsplq67wQSFSIiV
1D4JIFJpY8KZFYsfQ5V7YI+GaIiJsU2TzC0851wS3ofoxOColyDqQEj3PwfVRNcj
FL3fhFv1Ufyvb7/Ywl+r2AujBNTheGNZ9W9H7Mr271AREd+5qDlzPQiIJa57hlmz
zn127E/jKGCoGkl5LyKBaGkaZVGSxUrX0Ar3XjCDXbk0kEdaORdU87GlXGF19edH
Idb/J9gF08IZIHgX7XKgOV1UBJQNH6WOiBlHRKWth+EflHdb4X28hejdXjJLM62g
Ty96fdhHErTP22I8SwLx1Om1xHMMaScGJLWUkuMTNuQ9ZjJaTwKkTJ+l6JGfw3lp
Qxq24HpzkD7gR+Md5lW4AYKPmSmHukkXacaRhxqfBZYp2YZwtXjfsT9lA8YGV8SO
L2onr7lnuDt6TqlaG5Nbo1EbTvciEYMS3p2bHzZG8FZTMpsQ6KZWKTPy2NkjG2ev
voNE1+M9/CG80IGHiZctJEtRvBAwWScIEcVqP2+PhGJW0Wwa7kQXMVljYoIzq8jl
7j0Xvn1J1a8QiaarBX39a/SxYNA/tVI8GWQuJ2YUnuYaNH4YPdfRQ4J9hwghtGgv
nZbqS3MK8CGWe53Xcw4vOAkgzhCp3fhPFAqYlZ8y/22aJ0Y+IJHFzPLx+5sEdlXu
87Irnh6AF7A0K1WtVKjklj4Uh6it7itBEulJb7Jbp2y51o6jqKJZ2DF6qJvvQ+UC
1NrS4ioVvHqPzymYK62WzkOHzQ2EqBJS7DREJ9l1tK0rGJxMxpss5mCSpjdfMBWn
s+wHgPhumQcg7dRO4QfRfdCHCEJZvjzjNRL1JDgaZaKrvZuTtjuhfMUzePyoN73y
K74Qfllaip2GbQjvuaQaOdHzOd9i/0AzxpAMjc3gB+MeX1NtnNAS3VHQJODYRJv+
uMEHZTxe12LAchALN74eLp2tVL3uZKB9i786k36jHG+uauEQs8gDa47A9LC9RU6D
N8uM4amRyJ/7V7jCV2Eh71r/fRDScaEqCNXNWc9EsOgGpU/B2CGQYw7NPmHdDSd3
Xv0+zq9zSCPOLaQPP9cB8oVlBeJJUKflZrJZLG6NOzPpZKeUZU1qxpd7AIVuICjz
0zrFsjXY5AvPr3kNM7b9n/0ZrYrMFlGuJ7HD9BbrVPYLUZiTSGSXF8DwlbMXtoFU
IjuOigNnuWRJCAeBSaEQ/1G4b6NwlxfmUWio3AEbPATQQPAAnwJ8CMNvrUEYwWfj
eYylWVm5wRxfo+ZlMZBOlT0FkTj8yuRAZ+ef7uhSvP4dnVFsWhpe6wnZyzHwRIgc
GXHjrhQupN1pNIUTXZ4vlgVoU4CeuvFR3BMEv5URYdnB0YLFTqGgKTAX5y8ZNPO/
lILQ8oGYfvmIegQXMt9jtU6jjBCdYW1/xMjxmmJCwcjt1pD/idAdvvnz3stljZ6w
4kM9A4qQePO1gSfhprbVqa4nN3v7sPBTuSGD4Tu7NVeQ/jm6051ld7x+VGQguQO9
mN2REb0rC/P39lJOf+7BzAam8TNYMhgFromfMUprdoU3DdPR3Wt0eJl6RIv8B6y9
8w/8Pq2dnrYWwGGrZUMa2TneUyJy2Q8u/UYAHaCOPQCnRmhHt9zdZ6mkvZach13c
28TQb7H5ZnR3QbWoT4fHCWOeOZtSc1O5nMBXMzc6e6Pzwh1MJAb7EM1Ug5nirqrP
laUIoKNAoRNoOcnSjMuGKAskSfVxRFdW4a+jluBAkR7MWZmabcQLC1zK4jZuLFDk
bkGHFk0HDsnF4++nq1kTQS9HOgxOxYQq8fJwuDY9ysOdvmJrYL02gQ4PabFjHFVO
/1kUWNYTHnixXKW+K0KVRSlFK8r2hdhz6JHagV867Q0F8qS0Cbx/vZdbSqLi+hhU
ADOwmRmU796PmgYXT97zNSoj0HJQxBmfAUeGRWb8yce6hcAE4+VxTKUGjNszDlxL
4TXEcGaU0UbdrPA1nRq3Rcu6YUK4lu6rj9EAEdXl7xFqsQO6JCdwhqSD71IoYL7Y
94idyCDXjqcGI49H9xB1r9oGotP6Aj0M0yjrWjjbH1E6TGdjKjK7J7gvArNo8a0b
jgNhNlBRGOD8PpGJlWMm84mMYBTzzppeQLAjuaKHq+zB7ppuTv/ZETIty31tO+aQ
jod0noEZGSOpT5wx2itkqS8j577KmbO7fREaes+MA+kWjgMgUQQzaW4ZUcxG4yP9
7HdlSW+pmzRcDLtA7FFG/40khDFAQJ87vB821IpyxAP1X6eyi0UFuNHJ6HiqldK1
ZQ9/Sa3g+BHEGxv8V42QltNyftmJKHgqWl94CPHntw+addAv0ax2/hGyJyAdaXHu
7ifA5IAOt8gAgvzLnBh+/6j3/0SNqpuA25CA56FUXSLP9NaBCik05P+IxCv2B5LB
oh48kxLVxGZsX06FWOWlQS2PuKIMpkOR4yXNYJzsXQJb9MTl7/Ipau5XpXZunVUw
e1VKC2lPHBOZgBgnCCvqjBJcTIVrVljoCPevSUJ8hxH/NtKuNf2lfj/X2JHz+Wla
Ng9+k5YOFXl8rz3fmECPtqo2cLpMcB1DUL5T5DD70Ah5ceCDsA+seVJYXgntx+Aa
cSEnPriXE2oZqoCVs5c2jbLfZFyUQnHjRLHHRfa/MLdEs6IN3qz5y1TedZF399KO
OfiXV6gzG+N/bxavxD8LGeY+kzhmus1LVTrPgl4D3CV5iL1wCcA0T4QoWzIL2s2d
LYUF13HE+wIMoJJtshK783bJPo765S2YvTyp9hr85ENCyylGpIEmuwRorsDvg7Md
/LzprjWz2NvNwz7xZuPk6co1mpZMqcRh/m9YLJUTe+X+1YY3YjXvCEExCdOQT3N3
dk6swEgHH2fagXsMcf3vNg/yBagFwZYaHDbc0UeMor8/g9ny6pIcggAxKnGG4AT0
JSCFwcCMyiXoCCzf+ZWFARnAav4fzOye2KXOGfvEgfrNYBqtx18TOJlMHheY5E+f
n2aYXbLy9A3/CDxUw6oDU8tAf1wgJf4SJOiXrdiRTeam+ljGS94o6slB64iZ1Xp8
11ItwY5450VxEYc8s5bz3NoFKZdOK5Oyu1Lzfj5xUFxturQhLPnJmhTt73fwVzyn
JkyljaXeWMV50fiJW+Xw4Owrm06+7bDdlrCbxzkspO5Sh2CCunef0saDJ6m9h4hk
5cYr/nhKUFrb+krzfXU+suxieJ1HZ/oXJ4z/o9fitsN5BLJtMG7Xhh65KJbDe7fG
dPJ3wCq93GtTvvG8NE3cJzb0WmwW3rmfSdq5ZvuYSgAGZCHUMwNXvazOZOjdS8Ui
a1zGf0B9m1V8c5e8wET1tTNoNTmtsjRnK6llcRSfBgpIT80oQwoe7oD3uSrP69bn
Uz/Rz7nhsg7RTEr4pDRrqGth37pJ0ey9GJ3maEYwwja/6Ksu9G1nmdbSDHTOBcFT
QSGbhDYWUeGp2GjVID9neqOQlKTCY6FkGZPKAAU8TNIUBX/iOId7QnMeKaBd9Tsy
i5GR/gRViJX65ogmDjXEo25GIGLwi6mZdam1CHJbU0f0QOPKE9xxg6kX08C5at09
erpus9I11YfBi2BTez4x1bynNWzUk/z5hycROTiwc5TEuKmBoYruLtnp9oS5y/4Y
aqNLS8H/xfv/b7bVtEb2eLKnbnzbaMD2vTJ3gZ5qK9e5bth62llzjf5BXGzjmZcx
frWpUdfjikbg3bbdJnxhyhj3OLXIjsGeEUPuHdYVrt52wYrLjGt+uhiWvNtNWWh8
KSyNvaCDvgV7p8r66w8IQtguW2vwwRH+jQCMG4VZNMiS+6PDliP+f3JjwRvMyfRV
jzDvyj19Mdm4xbf9AmHLUr0mnRfA9vocN1TSwLeAIn/cuV/5IQGqm03zIX+lLlEf
FZoJ9xhS0VCbP+zeTn1+6odTPNqTAZUXyMhp4m0RcgVNtxet4Qe3HOJJcqAEVA9/
W72PbhZBM7fbys6WWlVu/RTI9c/j0m3y8d1pr+VPTjKjLolp8kh2ZQPbEQZi8eXc
kL1HeTuTbPWnNkJN3+wUx6WFL7eZeRYHyFxtPemFUnrwL44WAHY/Kh45ba6GhEnm
oe/dq6CgOEDxSgZJRwzsigjTVI8LmVVCM4SdcoPSi0+Bz6PyJSJCJdSqyx0zoCCp
6om5ZZyZkcoc9IhVEFLdZe+qQnU9Wsh9QteLipBqUIMKsHF4eJ6Y72C2cVggV36s
dus+LLWXyfXQFF+OxCZeKX3PIiZilzu5Mb5cxe2Q17JWxNZLScw8no68myBc1uWg
5RhDoSo17O+6vfIu1hxKopai/bUHnHNdTNUqGydBM/EqJ0m1PIw1yZ6A8Sk/ULK+
AZV2u9VmKRH0RBDz9Otw6ml6jlgl+SqXceHcXSgUqhtbEvEFUW5g0RmWygvL6Oyy
SLe8DnBLVR9Yd2E+t21a/zjZUda0w8XC62wHD+am9OFbQwB5vJQ8Q/O5bOQg52JJ
xcq082Rbnk5m30zfdxlnS91HPAwqCG89qrdHeBqF+hl7lViEcsou3QTRuyK1KUTs
IJgWOkYNzVM8TlE2MUYi0XhDeUd8P6SLY6bGRDl/8vdQPtOh8ofsSr9PN3prJALG
CDS+eL8RLG/kZQnnQe2g/eHgt6qGn7zd60otkuNnHoqhKbSVDqKyFJwV/1dgqUih
dEUjmyei4Ycj9xVlzksg+E7QPoJlrdQr/GbBUUGEtGg6X5KiqXO16TbNV9jyik4V
CSr/ou90rd+LaP3GG8AJM1aFfEl6dauo1NRoyjH+1P7eJq9MVffEFCsJZSDu/6vA
KMq1JZEIBpdI/1R2cdZncNBlCiCnJrdSpbbPj8wnQHlV5ayFZ4d868lrd2fE1Tt1
15Mtv5ea5lCFc7aVEty+xzpFNYtMGi3fsKAbbxePPDcnb35OrD/BWY4ZposEcuSn
Abcrm+hcrMazlTCPDsQd4XAWFjwupXonovCmNmZwDsSk1tF36CFNf12vC+K3G3ND
OHX25fEG7r/9b9c6hROyRDjKckkuflpjrRDNCbjs9dMstq7sU2mfLsHiVSp9P8By
ROjUUd6MykvrRZPS+ycYGKnIalFfjLfceJNNs/wxFXwSkw+bI0OZyDj0dFDQZ+/6
NDMDN28y+slOuGTk2qNRH+UgytbcxuZGJG/wW0UtymC7MwC4TzJwMb3Zf/xrF9fD
NVbzHO+uDD3ZpVrNBLLyM/82iVVr3m8pUy94vpJ5NL3Nw6zS4TRRW5jbOLrRQ7xh
T8iSgCqkRSwE6/3QjTyK9p1JcDf+G8Z76uRDHTUM1Oyg/oFaLXzPzKterk85Hrv6
NCvcBSj7MZr00EVtN6XLZooIJ3HsQGugTHo7tc3vA+78ts1TjfXwa3u9DTX0qP3y
Iy7U7biAvc8IndW2XZxotre8U+l9ZLW4um+bcWSaNg0ODxmBKCnfv8l2GanZ03CB
TcF8nAKF3ZYz9LyXo7eRyEuAxW9BH/wMmWmvFF6o/jV2xHp9tJfRxeoM78Wxgh7q
D83yIWVBZSaNyPi19ojz6duBY56gC+2xJEHS9sCoIGZDdxIUWeVBfPmYRhEaJAWv
aB3RE659boCs3Y+7ipFhspkc2RYGantOD9bhNV9pL3W5Km9ZFRRPhy12+xQ1PvlZ
QnhEZMEpy3v43dYtw7AMusKtO57rr1w5fcVmtPDTfpb2EngKizXPDd8NJcoyboCp
F5m/wa3qCROBMbJ2SLyG2v1jRs4CIZKA52EeP87uCcNsiKSAEUwCSVxAM9SKdm9+
lIHCaxKHULahkZCJqKBHQiPIPLGgAW6O2mtIv6vDr0A5zrl1rZUb6ZMQ9CvVLgVa
3g/MTkBoSYxsnkEyaPXDQcejPJ6DyPOLVvprEqbClZDN9vBH7A4uDlG2hIrKIqwj
8qKBTSrGGwr6Zt70Ei6Q/7fAfk9WvKq/1iPv19MmcpwKcfiJs7c0ystKoKupxs79
nQd7Sn1DVb4S4yUfXLrNs7WoQfzuHR3wvdFphkIEw1icd3U3FCVN/D7Lg0sQ1spy
TmFTxbwWwQ5hl54iKz6yUn1TPLFu3Jp4wB04RV3pOiu3zLxTqGJAVovhFD4q8xi9
wLvCtyZgFkzA2I3xW0e+FyZDLjgOmvF/2Kp3CK1a5F+hqeNIsUJmUlwblDsLCIcx
dag8lKCanEkkAHUk9Sf7wWut2Vts9NcaytVbG55oBL87DSwbkDyLpQBF4h+aIoIw
2a51rlImBTbdpJ7Q3nQcWT1TxxD/zOeTC9BqbkzRxs3aFqOxzM0gYTWDJpnhu4KE
MjkXM5W5AGHUGX4uC7+7vdH0FxKb/qrfLYTgBB9jpFQtsa1/D11I+DTAw9mgufYr
NIzxef+vQd4+ezlnD2xacSf+r3sV96COH5hnpilD7A+Ckw7gZOEq0j4/9ujGcLph
cmklY/V8CVYFl/apI67yFCPppqbieTL1cBiSlBkGEuQraJYmGq0p/wTJ3micQoZC
1bXZnedZPqoP8ZYLgdM1E2P2SpJi9yVdPzeaGYJ6Wkraa4QkF9YoldhZMvd2NiF0
ezKhk44eBamIWIshF4Atziw06MGPS1ebRCh8t+e5t18CVZic3FUuSnp838le8HbX
o5DKlOMA9ZRQp5+rVDdhNraygASUsBIwjVsePQn2xRCDEkcB+xJF25Gyso1EOSa/
WpMqobH4A4e5MVNWjoQNUJtrksxJgxZqimD2SlpLdXKc6ie9TcgWBGcfxKCVK5A3
00mZ0t8XvZnZRG77QqLMleAFCxED0ca51fVXenV8KkgsxLkggDexaqhG3L1EQ9XU
ZLY+NRYtiEd4Lo8gybffKnX8zXSVjBedjakZ98wXXxfmeyau96KPO9qWZk7KHxNy
Mt8/+C0iY/9RBLiKp7O1fhyqB3M+oPbF+uL3Hl2FB9V+PSohW+vSOlw7AdWIQTHz
eoojDirmc3GGKFNbJv5if6uD3jKuYr9HqKB7BFbTE2cRQR5/gOEmZK66JtSLuq7e
lCptG6w9t5oild9E5OT22i3VrKU+Of9sPJQ0oO3Cz96w1EV7d3L15+5d6ihu77S9
d6a21eybC9accTK8D1R3vws4F+ZV8996DB9e1Za5s6uGrQXzOU22iWuFXixD2VdA
hks7CLJsxTBJlJkdKHr4GqbRzaKI3ANd2a34sqDx1I31RJ9FH/SODYX5cZOHIJ+d
mXf2xU8nDvJ87IFpxnRvioXeY53gI/6jSAZALJ9jBvv3IuymmgHeYoAROODSY1dL
2YPKeVWFssxw9ohvfMlUOQGJw/AJyLY8JN5Nn4RiY37cfMU47AHsLotdKZCadb2D
TkK6wtKOyV/upZhoPmN1G4CswHWGCDZ+jI6nzD6R06xbm6aV+gNdgRMaQIZhl4G5
aII7CLdiBa1ohGM75Xtz3CGGLtKl/M41dBOifve+9nFUh1OqnPE8u8u4xHuaa+ZX
gbi6atqYH86cD/wKm3JxF2te/w8FVTM7v3qKgto9T+h+jsaTRxGj5vWcpaNDUTY7
ICzss6fQJ44//0J89f+CB6LaHRKpNTHRc259k3CEhuv0do6K6STrDigI9cO/8iRW
bWzQZ/z08XFcKhgySa9bMBHMPCGaF8z6z60A7vZkJwiiz+Ev+xoQbL2BjCc+sefV
Nl49ruKUjfslm8St6IhCOAtYrM6HF8PNHbt5Piet1dbexX0WXPZdxB+pyB2SscPt
sJdBCczrjIV1Jb8WMzW5q0BP/PT78D7Mh0sTCEPL08z9vOAkCxYn3fpoP97GDNKV
Q8IK3IqRkaLOVLOfUMAmVwkffL+Lx2XfqycLLRzMMLHVMOfGbO0+3GUA6ZrnWNhk
fvXNgqxdpegFknuM8tkO4o+FStVMQcCqhpO3j0oIJeZwBCpVM++aDK/vwjqPw63C
Zz1pRLDk1F//E5V0zZJCy0vgownYSTpk/SdhbSeODNK355f7sAFNBgb4eqR/JoKw
WAf+2DWQAIgp4GjhU9MpQGSEcxxuiOgCsr3SWNYnzW2Q0XO5tenYON3s4q2LXPbD
xWVjJit6eVRPaQPQ3oXwDVQasY2agPBPZfP9UBuv86t666ecd2ppehG1Z1BGd4we
ovuaSWWHqBOIyrfeNVPFSTe9dQDw1zMQgBCSWpDthC/OeHlo2lKgkH/r+AT2/XoN
FICdWBKZUoG33TCnz4k+xykLqHnbyaIUhxmK7OTKBpTMEo6LYHYsYjhW3prOt3zi
vfnPnGrNGncmYBNwwLOr4Mv/9GKlnsgI1UroqbXh+J2Fid9qG0g3beAKsEJhaAF9
44YirODJiYGZvpSTiErxLQrPxUGJ7et0ZXj6NtmgJiJkqCXFaBpPijlReYbK9F9v
ACSffnrzIfNAm/ECThDu9sSATd9oHkdu1OPcfBFnWuxBsKQa5R4sAQI+XzeTqtMz
Klf6wwX3vE8mih1lw3VDCMOUSBj0/ia4U402J0Ec4YJIa7aUA9KUYgNTnILZJMK2
8Cm1eeLHgNljKN5DK9Z6wB3Wag0XwWUdXtJTfCCKl9w9cPnI4LwL65ca9/+jVMEO
5ON29DKUCV++m/BdKyXwNWq4afkSXsCjeuKNRN+bsc4tIMbL/M9clAaMvr4cOv83
bEQelSy+DcFfkCWJyYZjCktjsr+hIl2phcG0eJnK6px8ejECuoHilwI65QT4QKZ5
1eBX1hmGsk1mUqqw6FKdUYPafq2txh9EQTqqPpBrB7x7a+XNzlWnOsVX1djsg1e5
puwsHCUZA+By7dKYXtUiqJLATDTumG+AEyy4EF8/B/DH/hkPamPXclrOCNZsE3sI
Z72T8Eqj+HlvX3SDEIUQAomceyyGj2DElIr572WkQn5tNawCRuOAmJiU6bITp9Ng
RGV6lIGh4ZJICo5lNxWwoNW8Pb34WtWWEEHVoHhlxqg01NMFgy8cB7+QPrYQ/p1j
hwTqk+J0H5vqn7FpCGfl6W/8iHgtLKZWy8qdmCH2uUE5rg1aUEHWJJ9IM858xzng
keb0bZTbhpHzqg1KJXF0LR15z4Rio/122F0O3ogMkMTUuYr4p+dM5jF+WqQHB1wR
2YkdT6PUFism9+F3CcZ9O+yf5Qrc02N71NBoBZYny/YCS0mRDU3lHULGXnBwfUGz
2NSUeoDyozpnx0th/l4CYogXoOFfZaei806xhYLBSjrWfqky1cpBhhihckbuBOnd
UgEbAqm0pe4Q0cX9aWfVnDr9XC8TAT4pSXj3twDVLkeWrycE3H7/UR5nn3xTL39X
veLZeTQwqfGGXGQujU0nlYYPvLmgaAWx1qALGkPGNMH7LZubLJ0A9JGxuEZhrrWl
BeXwrIn45tuZOHf5DDpnC0/X850TIdLmNpKs+OjfKXqY0SfjnrXvC7yNv6aw6c/T
QQ9UEwoX0TBKrUAzN3vs51DUOoSnntT2ioxAve6olvz37otb+0hGzvH8+QiVnh8r
jQcnhqpRfvRvDzTDHv1hjn1SlMjdSQl+bYaPpuLOWe8IP1WlPz8a06Sy4RNa01Sg
6iwueDF7o+rJmynl+IUUkn8Apk7bpbOIW8X+S3QOdWmsuEhvIkLOx1GcelYQ8eds
tRjcy+SNHJH7elAoworn383qR5I+xs2FFeypSJgE28GRkRVneLnztX30t+WvrvWf
3lJLma6JNEp1V4VFYP/y8NR9gavk+M8Pxa9rKeDFEotHNIrkkKsa/dcgc+NhQVUx
bCJLnuerjDSXEmbjuoSbauLdv4gCploAGQOb68w0I+C8dL5hF2ZzzsIPSrZG384R
aUrpngNUu2xutJVDqRo4FG8uuZe9liCi5/IrzdhEEsKER3O6WkN1mQ1/A2PBcFKS
LKIhGedmEpQ1e1cbOaU0qP8YkgH0CVq4NUKCp9DlAk3MtwgKCFVFEbrGAqlX1PrP
FSVGOrWlrPfQW++uWZ5l8bT0ZiqPilhYK+yALZzjbRzgDfLt2auDTB05mqo0RlUf
fDmoo0H/XSy3usq4XFvlpbALZlCkzLAdgRMil6Ds98GBmx6KmiAe6UZ29M2dosI/
ggK/kfpQJEpO4A001tzja9tUUGVdAKQbmvO7OeVQm8jhwtb6mXTiAMvxMMWkn7cb
62RTpMywgt44N+7/YuMlpA8mM/OPikUwAeYLcn2+lwrcrhU/xxZ6S1oJpzYPZzhs
nONE/wGMyX9xJPUqg1MbsQrUxJ4Ky/KtbGNPcS5L92qf3VDvp3sTZ0ROycv15HJX
H/AuZhoYVNsIepUERmI40Y8sI0bUMFzeIxtxY0eYClbhY2ZH0TE/0HLpJ7V9yTw4
bvpveGz16mQVk83okedFwYdWeTjAIegyVD6bhPzRqkAPgr0aQlC4XBMQ2YPJzlHy
TWhyPckOifqPPJH1M1l0UkO0dV2vr/gRdKPUu+E8mHHnOZXHmBFOT9+tNVK/42zW
tKxOglvRP34bgDHx/aDaApt7Ny81MBk51W+m5+dX4CLsqi33WGNS/KYeIMc7OH+i
9z7dWUDBusH0G5biuivhRjG2S11B7PpSfwu+Omuy952O3ffICxM8ga3P+JoA60gN
63hErwZ3pu2oCSqDykBQU5xjqFltUdjfBJZ6XEErDK4grRwIfQn9yXAwMk69TNxn
Q+9lDKyiGTCDr6/mRfT3mOC90QQJIhyxyhoKfGb/P/CjFIc+cRN4+k7V4D7LAtjA
vexest3FM0NkHjGiDyW/tQpwLsqzwBpny7A0m71ZZkL+hP5cwbTbHg+ajWOJ7rPA
O0SvO0OF1ShFKgdwcGDJpK44sgQ7gldsjhNj65oXqX56IGqfIbit0oSm8IdZkh5A
H4+YUWmsK1Z9B5l3i6r462n2m/moHj7SUWb7muDWCdH2uNLEK1hGdPWFelKgo8wV
QNLfn9+5U4+gfDpEd8NkCD0UWHipdN2evn7x47ayfRENAr4ls4dmFPJej0JEGqOw
YNuBvhUqqdS0XorYnxGtdDkPf5+3EafHPXw2VAplfwjzgLVgypPda+Q0ou7XPlfP
8czIu97e3/jO4bNWNstd7bxFfqujmW0Zl0Q05wLyl42XU7/MAeaUvqH4jtBzClK9
SYIq3buSgXteCz32pBjCNgQRjeq4a8eEHkH8EikAqZRJ0M0fqxZMiV6DHTmgU76F
k2gzN9vTjwI5W5jCidL16kyeBUAZw8KOf/+fOHNT0QDVRihaRyTtjQMNpEv9gjW8
Bfsaj57IfjMy7EZfwn8Jzs9NPxmJEPMPfu3RCTmWA4fMA4j3mEHBjUb8Yo6yEZBF
e+LuLai/rukmBrvfvBzLlWFszykNnrEzQLXNE2Iu2ptatrV7frt7r6d2ncA9W2s8
sQryog8vSCd5Ht1tVaxNI7ZYHESO80QCd4OZp23QsktIccO7Z/svwBBNQC0/NFoS
6OZr+M7b3SA4isIDIGkpCdU9EvRwxqaenbI8EHb++nqAdAXw6AGhSo+/whDmloZr
DnUE3T9949skM/nOa7gM15Ev2o7f8+LIruk4yLCcBXMDW40JV1Ng539GPxMYWyKM
Wii7FOhhspMHNRm5p7Uo8h1HpkQbFzYAa+Q58VOzog3WW4AVErJwDsDzNUvAqAcF
ZqD1chVYNmVDQ8b7lLF/nh7MkS/WjnsL7z07LwmoztMUDsBdgYsauO/UWKmRUVhL
jh1BRxmwuyB2DUIOHKu0nJ+hgNCQ+bsjKHbWNqLr/8geohzibU7fGdKfjjQ1+MXD
C5dzCmJTV2VUpuavco1gnFDvpqwRfvN00k5YViC9lmogx4JobYmI9+9k+Mk/cVtE
n3aK1sQhGmaAVb9h7Sov2BnUczK+6vLJwz7qjmidGnNK/ZJJMCW8eZZ7nc3R0b2/
2NzvC6uaUtuc301J/MH9E1VdYGyO+2o92OlBRipJKxleVNY4OxJj5PgEq2S8EB3D
lTHw4iKjUW2ZzlztBPwIxpL0b8zeSaiXePFvWQD8pq8gRj7e2a3Gze//+h7tIG4I
rBSDLcX4WwNbo46VfsfNiZvknRfYbsu1sdmyhjt/+JMm5+I1aSgtSgrK0NWU4lrY
rhlJHbQ6kJWhItMy/AtUXmtLL3MMDrxFKRMg/3hKwrZTeLodt3NY6dGh8fy8xpkE
ElcpfSz5masb2quB3D6ODAOszIxnyCOTlVcndWKYspYHJ/gL7fBPEQshypEpgRoK
Ja7wEQkPpZMDz20/J1VI+KDwY6ChtCBN3K1G0WK5EK1EaWuL2vdlm3L0/7hwECxM
NIDEcygltTXaCW8kuqRfioUsAUNwMDN8VN6zfyCt9KP0s/SHuNBkXnuxkOeB0hVm
fCEZyObGgIHaCPx+Kxj6iuThVZrXxsbzt8upbPI0Cwm8A2aJPuBhj3KSyoRuu1CR
eg/dr/mYfe9gS4Z9hRb5JHbU8YqfgaeK3CnqWpqhZG35tDKtH4YIR1LfugtzDf4M
eTPsqVBc2G2trbDWuzvCtritQOJP+4li7eV4G6Tu8B9nv+jWGA5zw5u8kKuYitOK
FWh8jGWOA0Z61vqMKvggyFTes3/BljvjF1pcv3dnvlxg5wdKZOvUb6yCHnBt6Xqz
1CBfy7pUdi9HW2WHe3k+DIbTLMWr4QSlyxJ6IlSwMZlYegeb+kFFwUgLipBgn9Bh
Qj/JX27yOPzLsECmESM82Rd/ztyhG8rpawcwHmaSxuodkWYrwel692Z9K97bAjNd
hjTRHpdCM+XJswNs3V9tfQ6dXM71lrR5eNMOG8jqIFM6bI9sXeuR64VqLOJCWMDB
GAP5W+7uletHi2paklpdieIqoMFtiA7LNW1Nj2YC5kXk1itjHDPIxc1uoGWHNPTn
IQbppwXY1NlOmiCl2Rx8+gJRmZK9V2LIvX1evP40pqyARYZ00UWR2RfRkO46KvPa
bc9nmfCHTTYdx+0W1ag3FU+SdtH8vVAoDSL+NZMQdrCZBq1NhE+ztdy3jhKqh11p
c24Ub4r8Nqz5L7u4lZC5Qed6tzYjMRPZXl3rMVQdSgQsatzX280CPHK0BrA9s+Zg
f1SASAU6annXfkZQxtizhJjEv1DYEInevNKaFG5N8xQO4d5eJ+bEujr2Q12IUctS
EPtzBXVGdNicCyafav4p8fxuLiovHZ5G5bdW5MAPDC6KW5eRIyMOoopoOFTlO9oj
7WdzaQZHYatR/+9KKTqETuzPxqiI/NW3yPVzPaKkIqy9XEGkrESo/NMtlyojOQeh
t7+bv0A7bal74JtgX6qrKryhr4b7O5fYQGAN/2b+XmcYGgtdB8ZH7Kd8iKHozpLP
pPrAqK74fspS7OwNaZ1czDDfjs6JN+Jj2ec8DXSsX8ZvsD82dFxTCw44BxYAMTLE
H5NFA3BUemkzL1ZxEm6zkPkVjLvV9/bugVgqh75eun1VsgHNMvLtq71NNDK2OLkI
tMHltDzBLE2o6Ljt5QbgYsvYYjBhacrMVQ81dSkc54QFwyCaasENUEUs0eud+3ys
V+HSgS2TjmNL4SGdBLi+n0LqiS5GcsTr0mVu7YL2MeaRKmBRvWf57VJYbpcJwnxe
phLJAzxqau3HEm8/TN0wYHr+CuzoacZ90sEGBKeEP47Zd3QomOCiXSBBvVfwfFRC
THJR36QIJayrtwAgQ+vMfulb56R4vVHnUAgLzcOwubFPatwUT+XX32gRB2Ciy77f
/hfZugmko6UGwM7PCpH0T8Gv1uxcyweDJYwNvsoK05vV9bNXn4YdKII7GD2oeOM0
01xd++ygeSh/qEI43kr0W3z4vztjd28eX9axicQzh1KkrOMidX5eYaOXwxpovjDN
YJjZMZ5UOjhAIrS3qG6MGU6ol+pjkFMNdrKP4wJFk/DDRD6vHV54Kx4SQb/milwh
qQtHO4hLU67sdF7jaOin+YDsjxzQIs+oip3yk58SLoQNchosVq4Knrg/f5Rg6ltT
/t2/mLkYEasT4AWhWbgsaXVIu0JWjPMdaOm5Lx8SlCWmvDQaKWSf0sq8nNjVbf2V
wKVrSwPX/XWMr9xglwZX0LXRUQH0NtLPgnGs/jldkXc5mvtDWZzTgh+HMGHDEf6a
+KClfVN1a6/pBSO6vGPznh+bZDecPb89LzSJMSSZ/GhrjqT79gbDZFrjjuyui3ru
oa3+csMoyK0c9hV4IU9XX3bArKnQbXWeKp4ZS2sL/4okA8gFs8ldQeGO0da677DA
+FK/h6ijEW8cbTiN4LiXYgiLB1V8Q3p0c8rapm43Q9689HQGbKVkmCq8Dx2NFlvO
fDQ1oEnjfJNb7cZTqHYcRG6PwN4/MNstgehQzOt15UmAYU8SMYYE/ERdmO/CYjng
QbJFy+QGddYO76Nl00EvXvkc76w/7i7ivQJETA3TIlDFlFLByBbp/pjkO3sZB8RB
XuIl1oI4Wmjv73KVm4SUiu6eYMgQGtjB9YoQgL+/LhtvNGjiXx7okJ7M7WVWkizw
PZCbJRBj1Th5sTcHQHE6R9bu5Ii93nn6PUABILsFujOIldZyg16DmH2I01fy2o/S
i35xS8SK3fSXd/Z4Xt0trmi+azbej2gU1NsqQE4rcxQo7nBG4Zhws1uraBIdNkpX
sCinpnJiOpa1bQLWo7tfTIR0VQiVAzEOYj0L7XH65LrFBwZujo0vKByU5xo+NVZh
S4mzL18IgHqtdHNHBdpHZw8gyIuN9LPt9FI2HhhgyV7YjZXMEOKY6zBfzDnnRPE4
yzdgdEAi5lS8GJcRKkEAIKTsyMqmZqXX9KhLcpxquambgQCCNz9ndNkjgFQGNeKI
a3x2IaDF70//cQwh4S/8xFwClfJhk7CP8HgV8DpKnreIQp3TvGQnrzzv1Mnm/r5l
gWyeYXP4jC8Fle8gO2enm7qdLfk8Q7EuvYFd7OlUH38elQ+B37mOifEvLKlMzj0B
a76yDTNQF6oOlq1/94rOm8Q0J6Pu+6Ce/X1NBMo8NfIRQF5mqGkk6BHQQatmwJIg
57umhaU9G5IsTbYuMJguz3yg4Br376e9I73y1QAMhs//3SPafQuz87sPrVZETivS
FpNX6ZersBsyHGw7xpDpxB/gEv+4M94bL1RZQjjF31CC1ssZC+SdY4wPlDUYisY0
wezH6i/TsPwec8c3xX3wzbFdMF8qg+dZI4U3qvw9RPFvmPCQarZbeRU0lSfJQOFq
oGW8Sc1JAgY3pWsm2vga1IkBfuHb/BTdlBIg1vINIDh4UpywfJGF0tjzbQTQLzTH
Q+mK4ab9zDfo4ev1DVo+VmbHfaVeGDV5qwqYW4zE8FeF7CxlUkz2g8SLAct/rvog
DaWTwsb2q2mcXnV2ZcJe33+eBGa2gWWtbyCSrFstapw8/2kQtkr144XBaK+/OL4O
lbYthyispuhUJRIJmT2WLxAdVPWPmhPvJIe/FNB4zFmPs6pth/L4F1NJDRwaZG7u
1oiagN25RQ+WFrJwEEi64+kIi1EGDl/wh6BnusPRyOBjc8+d6HIez/Po/m4FWccr
iLOPBLvXzEz7ZqtE9da1FgeHuyvJNi7sAdT8vMib7U+Y5hkEY1Jt/MVbnTNTah1a
NqVsNv9dlvt9CNmG06vpU1l/Zg0OK+OIuMvL6JTO+FSxlFngQSCO0AwxWlip6v5c
APgvbOoenlA7d1yxbLwN5jE3KjN1Hv8HavRD+SyfJ2IhAapWfUNjPT+wrd1+RRAp
ViUy8uA4+uohH6LYqzhLjd0+YYOR6DHswi+nAsn3lKw2Le4TW6ykhWG9ZFrSFLpJ
De4rFR18Atc61T+KP+Bw+NTIyPDz9iWXJaHBBlFS+mX6YqWBnOZniYd1hKtGKL0L
v2SaiJsafAVn9Z9kOZhY+FuatgLMpcCgRsxCThKUF9elG6RsCfIBu38ETjcZ/gZi
FL3ErfBGrR1WrHy27Cc7y5G4+Dl2Q/REO7JhPBns5tZe2Q96CLYEsFty3qyTJObf
CBL0KLFOAtCH/g3Z6mClHnObroqWeA/t+QO2xuz1g0odmjd1dOv7kyxlhRaFNamD
pxe4Mz+T2a4Llt8x1yFsosw1uZbvX6d7v6WIxa8vJVYQ/tr1Z8j+wepb/tcaWaKH
unsCQ9+O3Z7VfYrjzcV+/Xf2wyR3859/mjlf2YLZanHHI/Mkff3OeaSf2x2Q/Eyb
tNewZp9CwSI6G+2MWrn7S8gfFz/7ipwYMrEiiM1ovTv5k8OtDFdooqVXKZu5+9m5
khjIvjJ63ivZj4thaJ3CHTo2nih3X31NpGBYxUSbUaPwnmq8j+ilKACsZ3A367KK
jliOl0/inmabsj7jFjtKsIgvjc3zzudiRRfKr3j8sO82GX0oleEkpbCVi7/yb7kG
otx1mQFr3aNZs4dR6GlBZjbHuSrwhzu2zi8M+jtHc3BNwinQB2ARnIKcFtIBYOok
TZI0bJjdCvaCfErCVCuIci/AOU5EhtDYkaOIs+vpV6E1eo2AMJdpVtsaGY0qmAdg
2TdSvjNbJCJqLYK/w3hrBhkEWoT4GThZU8WrFmf8F0N7K9p5sYfjlWph2DRZ/k3M
QXXmcAQprXQ0HZJrKgIrujg+bdAA8GznX0xfCT3j878WKLJKpxAPhKwzhOgaRNM5
b4+pYW0mPl9J2uPwrRL7xqtVf0lpMfBFbcrEbfapSFNrBowyc+xoMj4JKv8aqcOJ
Rnwzs41K5szmNyiEkoXsYMk+/mmTTnWwRhCQtyW3xadiy9csSWmeVa8Dp1cSHZNC
YzinOoPlzHqvyRkW9JHzrSEhb4nAOQXamgwQd+uk3ktvwztvOIXl6VbqUPuHbIJ7
yuzwR/7RxiX1SyJ77P0Yf2y1cR/NMHUg74XI0UJnMvvx1mG0mSQfiHSWiEURZlCZ
qr8+eyzMfkvlatSyyMpXlK6aryiaS99N7GUo7plER15bwge5ab+cXP4HnXfjppJj
B/oBq7m+TI2xclSLKlbsjXwaGdAOuoCTByneIJI8sox5xqMkAlPbTgb99Xm8trgE
RwC/W1FV6LjapDUTvPKA2la1OkkMgAT1PdvUSXs3RZAad2yTjvLTvkBaDNatpqzL
P+IF6Mk4xK0t95ZA38UdhNTG8ivvCiL/8/t25hIvwmFuMHqOePNNPsUYexncrNxa
3AMcKOZCPSQ+l5Sq9rFFprdNiwH67kM9q9VOK9dzogZPKQDs3uFJ43lt02fZS+p1
hptgyTvjYv0qezT++B3G80GLHnfjncxc+aua9jEdh6izOGsrs/Nf07Gqg6sxBRX7
gBii45jC3A6aG3fwWo6sP2s7toD5bT2LYGXlIPCrfYfXVsOvCcAWHlX1SpSLKgiN
LpvstdtXA8+p1KnvhTKH+uHfyaLuLyh7NW8ITOIUb7tBbtl8LcboZTXWJqr2AQtO
CK+ZNBcbX2HWptfPV+lQ54yh9olLoCVJCOSNsvTZikYbyURsuMB23U/gZ5xmzGf9
HqRQaJZPc77nNRVAfJbdd1AS/zTjd65klGAr/ty0lX0tl1GzW+poKQMP8bWOixtN
RiFIm5A/Q56iU+aMHoiJwkD4q3edO2Q6+Yvr1r4QM2fuJxmULcYIUu0VaaW0wLK9
fV/7H/brG4Ghet1ieW3EjTSSzGtICtRnQsfrjWhMs3Y0kvF715aPkPON+RoFPLEU
xvj5qrD8Te4CJw21ddEWqZ8nU6gJUtXzBDRfdAAbZfrhuzqlPiXk1wV7bTDiHtrO
LCH/uP6aRWzblPrUEXeccVwEk1HPSDJaExBNELll/aV8KHCFBNPiEjqhPcVnqokT
2UhU6jeSUShGYyKWIVj/Vrk+9cDU6FL9Plnv99dS1+nhlETazzLt91UcuBDk0ddZ
/g8EPhVHe4hFKvaeI/eRi+LOXPga/3F3Q44rTnnPiukbJofu0yYlQbMZBZGq4BeN
bALQraHTxttWXXQ+aiGx7L3X/+aGun6RpXGQNMzuW2BgWZ6taMqi4Cwjy6RnySEl
nek6Ld7r1GZeHSQ60sR+IBI76X5D+4smojdkc2GbcNC8OHaTGiSmf2qp1CQi2zMS
899shNui7Tsi8a3HUfeZkWOLJLA9ljcSMOVSlDYfvLfqDSsNwz5WrkMO402XjjgO
ADK2Z6PO/uOuDpstE7B7NCESdCV7949RZ/mtP7i8ggEyex7EtCfVCZnj25WO4lpw
DPJ+WfYeBnlzB6s52tDOONv3QLFh7Khmj0J3grYQUFiNwzKXSxpE0ZX5NXvXanDU
bXxS/N6oUNA52ISl4/2LkInEmee/dYVq631dyBjZ3O7+fYgA9Em5WxWhvF0Qp1vi
6srA+ON10SM3BbFIuk6i6bm06r/2fLEDGC1jIhdgBleJcH8cnBkLLep4KOW0E+++
/Brs/inx1Bgl32b1tjVKF+f8Mrv96jizc7eCRAhDfNGyA7HfjQTJTsikIFOauL06
3MoOSaLLZvNobuvF7AopJdfBlBfY+0DSX+3uGfjB7rF/3IouGsOKHXwapEa8gKd5
yiNI0htoBc2Xa6mey4KtFdZ/ha4EanOWyul5mMV3iVVLPwk0IUP04GUEaZo5emy1
dGh0+CJDyLjs2Kdx7fCCxUQnADcdBqPTAxenTLeoqzpyXGz89UQTwBHJ0umIUrh1
t7rLTQDMhnv98SIuk5sD4AkeENP33LkiPNQ9rWGBCEikZvxYe94U9CWKszdEryMe
D+3zvq16En/+YZQH+rxXn5Vo2LbHEjXQvyZkRfRpGCiX03IZ5clS0XJcdOC3bApY
LmCqxjSMLgZn3BzCQ+ph65kOnJ8OuVPTEKJsX1nSt6VNdgR/q5uEQE6qFGEOcR+Y
soePKFo0c6gK0FjYAtm2t9heSb5519pZpUcl6vVvxawPMCK5IZDANOYV2pn+KGvP
55EkFMM5hGFrMhSv6YPHlBHfguex10/Woi7R88qQw9S5xmI3qVxrqWSkN4dUizn5
iG1/3WNbrbZBIiShABXAaW/06ojEJtynfTisVNik+0QPzuCscLlTWrNJ/A+K7NPv
2EQ8MlIGGeEOc52ynVMQPRoK8u4CmU4kpNvU+X9b4zYwkgkO3YOmIwR0NsPqwb4i
uAjJkrVPpjOHleHbAd1vRkmXYineI2oMoSdgHhIKQAs+zXZ73kVXqQlKN56QyZOK
OC+MFg0qK7J20nq6foJFGVbSeT/3xyIX8HfsX5XQYDEuAMrOt8wX2AGYz0Cd2Vt2
ewd+BeuHwrVE1rLcmdhAltV+UVnfTL93WSGZwZN9vEMCbYOVTAnNT6c4vC2lpjAC
YGMMyAyhXhktWg5PXXdLBHdqciuCChrfRmUezpTD86XmlgXAHK57eEuvppGf2RyQ
K1S1Ak6TCSsXE/3uwyhWRH2Z412COrOj0wRhsrfqy3ZG9j6cqgAWSsIL9KVp+uzz
9GaTvBWNg94H5f0NjrH9crLiYP4i4pERS54rS4OjIhXgNEJ+2h8YjwUoXCJKv53a
WkdzlNaRhwa9b7kYQG/Hb9vpGZpVUfGI+F8hAoDJ7ff30+JXdLIWdDs3x4u2XQL5
sJblWac2lzCmRa2I4XmumO/Z03mGEv4Vc7DN15pEIy4iageO7HPIJ65zAmIn+qCU
5rjQe36CQPyiSj2l1TKLu/rkSc78RI2K66QsaIi2Iy+FbKuRoDp1EacpKCV7aRkM
MsEYxXtyvE9PIqkH714vrwCUVjKohx37py3mgd5O+qhkEs2b/9jEt+wmvaSf2CAk
eYoy1Ct6yx+bj3ly2gHdUnS7Vwq0tn/LF8pXdWUsEz6YO8srCWAyYsHqLmHjr3Rv
wzHi6uRISw4l/t1A62CRZ9FO4SLw5Zj/7SRICXlKJqCspAr4Hprh4lFzWuAXsnY8
/Y5OzGYKz+FufWlygB+tMmFv31QQIwr4B094tx7dI3xzbNP+ou6Q2v5GQfKXvdck
me6dBlPG+fYNzZogZ+IXsf0+9cLkaqwphvrub8leC/3oylCUXQSAKs1teb9qvlUY
v+up2OTngtapalTbhgJFMEBNEJQ41LDmx/lod16aA9TDXbOzraFY9mq8I9c95dFt
x7jkVVD6D1dfCh7wXtLRbTXD1c4tv+TJol5O7Ikzq0g=
`pragma protect end_protected
