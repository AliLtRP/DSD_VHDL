// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:30 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZxjEYv+bO8ztwivDwbU29vv7QkdzLgWqj6LhGiS9zuB3LZawsk2K7d4p2kbm6TN2
Wu9P8twg5+9EO90MO0qZOju2af6B7fSiW5gY6HRk07xdFCcQZRGAAvA9WMh1SHsO
I/51Cp3bRNFnWUNTTaIyqSzRpDwGuYJJ9b17du1NSKQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5600)
U4t43tHuG6pKsJmis+k1x4uGu7wbxDlhPlyaViCGIidszjn4QwYZYUV8fKk2q2SF
ReKRz7OYRoD5dGwSy0TjrN6kkfmMnZ+GbRU3AJEA3BOK/uweht0RljAqocOUXPiH
0IQUtF/dts06nosLYCZy0u0dVGVbV2KzZ1gjwKbtx7xBXi2t+XhcdE8VWVMaiOlB
5W+UTebvukXpeBKupMWsvz5xq0DUII/2SyVOdQKd6fsNGcXywfZM835cpe2n+WYr
Wdu2XbenkscV5sJndkhhlhFQV4eNaTkx5d9cu1zshzlZj9ERqdEB2xnTxOrJEM9a
uFpEoXG9E+GMON/NfXM1R0sH26fGpT46nDOYRbvV7LOF01bwxFrP+xh/8xAssQ5a
RBrkEu/a7eWRq1+Q8FWNwYi62DkOcULeY06ax+nGLn+2RLar8GueWkOBX0Iia3vl
f9KcHliMuj8FEoV05P/nNmBYuDazrdYhANvGWYHvY4bIBODa+p1FNlByo6trYB5l
pwYxKZ/LqnKi9h1c3AK2ToMkmvY15kxxUiQW1Dx2Q0SOuS4otkuWI8E6Vdk9Cxgs
G7HCFerDCFwypQ6aHD95+DEr+EkaJ8NB0oA/J4iHYYR9GpDIX8T2lgU7FtdWkqnw
oghhb0PhAtbUUSV+ZwN5vrpBcnr7tfqtQNsoEzidbKOQnxbwDNnO1Tj2QP/iGUcY
hqy86ti2yzi9IWOZ43yGtxzUZhUwr0ufHC6+OyoDqxIdwEMKhrtKWMfRhwYM33oJ
kC8zOhrTaX5gjHXFDd0xUNhwVdW1Dl5zp+2J1bvhyb4TznIop0fSWrfpFh67dfX7
AXQ1xvIMArxgSV5OrXkMxQYzA9BH/dJ+Iq7nTO0vJnZdAf7v4yeddZpjUNMc+5YX
i1d7XGXsrKsRKdceGLg22arlicbejEzpNPFBCTTBIN2fjbcUWUm//r7H+aO7ymkA
dEShtpl17BPtS/LzeYGrq2UdLk8iv485MaYkW5/R30Cf0mQvDQMMS4p+GMl4LvLu
wbBhUlL/wCzC1jPSq3VgfKnVJGvSFuDuRm7DzWbRDVqeBXzgsyUQQaTPpcmqaFA3
QHUm3mHhIjw2X1pBdwvO/ioXoClVMnTkeUjuhCHMjLiQQVD/nEsE06OXJeHM3HhY
RAF8KsqUG+T7rtTW04mEcHUOZILfD17IzFQPZP6DTxDTo4wrURIuExJ9Qmzux8Nw
ROz63VAWKxSISyXUTCWEjk5vINhBmKKp2y+bF7qT9R3jv9wSnWjxNBOkOALKO899
JoqR2FavEkDeE/JPW7D0ydAVf15Vowg05sVof6DahtbaQYOsGvwE7VlO4x4ZdUYT
HqBsax+tqSfIcs2JdahsjyJxIm+bn1W0QbZMmv7TFPsyXP49Zj/kDG4vwxoz0Xb9
yc0zMZdtgx3kw7JNoPHswAE19W0e3getZiSPT4/q8poGMIRbFi9uaV0nwhSr6O1y
enTTfB04I41umOEa3j2dFT0WMzVeTnQNrINMbOl60FbMc/IXe84iFrtUgXfPqAeC
8Dl+bXiby+IKhDq9wkd+4ehu7ljkcZgqCxKsolKgGHF9Qo7GUj7qKFl0gsfmyzhc
YvLv6CBQcoQz/0nO7AZukc7CNrDWoi62D8HP7RNhCSdQ0zMY/uyZ1L5xmdWdLJ4i
IiY+iaryO8UIiyDVQobhHfRXaGenHwtGslAPOy3PiO9doYTpMIh/w+j4yN/A8UIz
VlcitTkyTpBzM4DtBO2eKVlIY4PJLmgvo84mDZC7ZkrTpZyk6hf1F1TSWgXetovQ
47tbmPyDP7nzvicpbmzAfMae0AQC4d2Azej4Xx8f8LNBGWBwtiWJ6rgtA4j7v8Xg
3B7bvCS7XP53GRYGmQKW41toRCFuq54hu07q/i63SFGNEKfUdioG/QZDSsiNAIbJ
dVbRBffBl9HN9I3WUENOElRmmUTD7H45JLq1MSs3VAyfKzxKHF2B8s2i3hblvLoa
aj2RsV6igx+IsoWSEnQ89+P7UG4QniN/csY5M8duQ5BDZ7xrxVT29d+g1wCCBEQa
FyFVzbSbXvmibYQX3FLy3BNpW2E8RSMXr949NvMlcK1Vq39NIEcNYRIArtARhjuU
mNlHJAprskuzqFTEkur70tYAWGz3SHXQj6GdFqitgUYdhBdBhcKNCqDfs5qghqOR
RL0cxsZ+Knv/KgJ+d+B/9TSZLfA8+xTceeQamJQSqi5XQ0FrPxC/76FyYn6gbnbL
JInKirt0X/tCwnnFbNLh9XZ4+aSzxDtzMUtmK5ngjq7Uo6nkvWu86GBoGtH/dt4/
4S83kViZEp9bJ+jxxhu8s9BcN5PASHXN8wRMJV11mm9aL+oeAgcqjrL0LY/FwQ7n
/9NjUinPZFCr2LU5rckSYZELC66TbbY0mqEh89pFMoHn2kOb21Jq0qo4UI5ZnUWa
5+LrXsOQBPCwi3TJtihE/Di99yxFPAKpcXUZ453dSCv4KE8RUJWfnf2AHOzsQfhg
Gp/edhsdA9Ckp2NJ5UulM14OCXO9epD04ufgpUB+vD8qNoD1fZdhkBlMaqyzOdkj
IFsvYgxUZqrYrh9p8ac/RcibE5ax3Fg0BdUhFlpssx2EURRJV3rKXp8QtgF7tjgM
duq5+fk7IRNEUQ5/i7rrWl5GIJuHz8frJCCbbvAPg/FzMj6/9aCgu9ocT6C73Mt5
24wPmKVAeJPXrstg91ByM0FEX/ZzqdGHI+8sjuhPw4Anf5sl2UwBjOLW6LbqlfYN
fimQkd8e79eNs6JKpAZnE71Z/j6+pTB7NgSDONK0C3cFlNrbJ9OfH648VNODtSed
IeTwHuZl2ORu8rTeMidVOJR5OgVOJNrv2lesA8Jjl6G6Gu8zE8gKskFBoVv8xoBl
tMGV3txUq4c/2IlruMfQpptC22iEiZdtdsYfgWq2aHH+BLOLc11yKn0ztIuTyLT6
/yCtgHwbQP3kxakeafHmUO0fsD4He7G/dhADVuEYvFNShZXQ4bQorHXUufbqbsQE
q4XbjYj9wp4/YcDW3PeWLteN20p+5bugTKSe4hm/SrEBQm3EvFzNHPYHhOqIcsW4
1Nn3WHQqHVeh5zWjAXD8K0lq8QJ3N8Np4jMY9ri5HCiSotXGCmXvvuSbNKRkuQyu
BOWjjYXAUqHMgZnL2F4bi3rSmuj0IpOERPxXWp7lSHLxkXCHlq34B17L0WSxT2Jp
GVRX/8IJtrhA/aw7G9swoArm1nRTDg4k1y/4l7hpSZsN4fVAsUFqh5ZpQNd0Y15O
QQ44Xk4b7c5U/qFbpKcM/pi/mwZsaWShcuEvjNUshOBk21/BoGQSYJnEi+9Np+Gd
kItA5sUAeu09V2ccBOlAu5GTbgCvOxIkZRFzFxoJtGdv7EsCg/wD+2idA7s98XhQ
cjXlOBoRVSWmfkwUhzswDxp5SzaViaEScwAfWC6F+RniRHwXqUkxLIkGoRXoQ3ky
jEv45SNMfQzkLDNwnAvJU8IKaVXxsShIJCXuLYkvnLOWjO8z36FdKkvvNFYudTI9
D1JFk2hi1LRqZcNBagtAKeWsI/AL9JEYjz9Y2ZHECTGQgadF+SHHnGTERu1UAEgh
aCdZq8KXbWefvaemKtcHNB+T9xhKGl7bwUql+9dFMyfdqyAhztnjzIi/vw6jyjYU
9pe7JMvJlAAyuIlwi6gNmSKSoTbcgXxz1HotDLmx92vo2zdinGEApXMZVkp3/ah/
2NPk5JbwTsxwuguIlmL2phJab9He7k+A5W1RTAhLrxSLHB2gj1gO1wkBSp87lXH9
RgvIISb993ey2InQVv4vhjMUFDJF74xa79mlFjihxEjpf62p7gq1cRO3hEbNK0CI
htKAZTdtjQ3XCX6ZomY8NCzpUEg4FxuGJGQXxFxdElGwlJZmTYPSnWC2/bOLkb5S
hFK7YMbsQHH0qeCLpUV84r3BM/0LbFXP7ghhbuuc1ojp7UCka5lao7+uHxCW39fR
1l5305RI4kqyc/zV8GqZ1Ap0Gs1QC4khjp0uOrNLjKtVMQTFgwiWefLXGEQeuxLm
9qIhAr233bONjSNlHJRqibBmKmTa7SuXSQXT7G4IW8uj9wvnTRn7WHJ22WEEpsm/
GUUxIHJc2gzG6WjGByH3U5vlCYUKxQ3fRyhATNKdBVNP3bFPWHyy2Nuim+eH9ahK
xJjPPfSlEQqCxuvn2zDZ0mo6EUBudcgrscgMzjTHSngTwemYpi7POyIlJqC1KDoX
JFKEz2ZWXlDx/ySX4aF2Ofto9WyxR9gcw+/8UGvzaPwt6kMCQVdpsRb+viw6a33c
lxDkkZADuwSF7Hje87v/UQ4I9WqH1t9VrLwA8MfbvJ3+Qsfmzuqb87TI6ogLCYrH
u+aIwdfLoooj67IxyXOeCRd1cez1RPRadlkozwX+gh/G1VRYYPt69fpHC1jayGIA
htgdNcbP+G+urX/55myp428Ed80yJHNCzragoP6qFTVM27HlKODIHU+S+6ZXJbtc
g1/Vs2B3ML36zLdlqNt0Ntv6zLoMo5nEv7as5uOg3Ii9FQJCxUXwkPWoc2CV69Gt
n5qlEwQX+xnyRhNdfuzZ8QnOWB+VPzLxGb5yjK8+68KLD/WiHer3nVNSX7o6spMK
b3B41O8kuj7wKS5sSBvV3G4eozDBe9jI/7s8Ct2zff9HpUInfNj0r+WhnO+tWzzu
yP0wwstbVHfZRAOomMItTVWvjkX95YDFQEeykQnDokNVG2AfBmtrppTNotH8SGm6
wj56Mdq5wE92SFVPFXByonmqkR0bSg7vUsbMqYLDh+L2/dGleJuPLtCwJq5SRPMA
SSvlu+WDt663rF6APesN7peX0k6cR3AjUXTkt821qg89iTyIoiv+c8rLaZJRi5aZ
MI+9I4Z1nd2NR6AIS0+zwqSEwDLSRCnLHR83F0NGAxRCIafWq6+KpNbrMyBIUtyw
CM973SWniU4RihkSqI3nNxAuAL8fHPgyh4bXSrmbEIe84ShzAmd5HSZxXAH5C3z/
YNxw/oUQJtqZG+CLGQ1WATkCWrNV4KkzpriT7G7r9ToPvYYhIE029V73luSeYAwx
oNwSitSO4LlMIbGbK/0UY7B7CZfXS58Jm7VWB9pdBnv6Qt8oIYjJ6vVkogcLEoBo
6IWphq3Z8LdTWKEJWhxDS4MywmcR4qJeUAntEKsFKkAPblVAVH4qkCq2ya+R6LaZ
lZL+j8WMQDZBqjPhwSUVWo25jyk7cip5ETuVec+htvKvoDxj7r+EmzyXeeLEChtK
lBGRdrokPuKyzQPCweA3Ndy3aSha9YfrdvcBrIJjPEUKN9fP8JBNf4Wl5ET6BPb3
hjJmJnHeu/IXrJShEIPvZ0D0q6kItqlX0qXIuQMM8DLVTmyyOwKEp1mLkWx4dyi3
nuw0f0iVPJqShMLELYgsExoN2W763un1NXHX0m4dtYkJpLk67MA/TPsMlccalAzL
DeNhVeH33BJYPz7Bywt+ZwzfGM4Q+q17PtPRwJTIiInxmKAqI8L8Dh527J52WOEx
qEusicwdWVW6XuslSiyuFE4vE1MAAom8IZgLEN4UzJQaX08/8BdxUFcYZkOdnMH/
W4pHTZJ29m1UmkxsuNuUxEi01SIsS7wsJJgX6jrP9clxSxrWBw4VvrA5kL11g8te
nU1oOHxW/co9Rwn/rPElPjul2KW2ejAjl5/UGsbVHhS7e/mTEodDVoksQKQ9NYy2
aYsG7maxZiXSOfSGhHVfuZth/LoqoZyugZRU7s5uvgEpPYl+Rn/yTJtd3Wtc7W5/
XeMlgnzfd7hNxsijCLyY3A20y1DP0o2nxay1tSWIVnYvKahBRVXh4UjRxZPoBxO6
DXpWGsF6bksjROxQ87Fq9Iv9h1K91v4CtslO6LJ9EJWPN3xDWqe+++KNtYAUXbNC
G8gdf9Kn8UxrY7Zzzj/REqSRxgtrCA93OaH38X/pdirioJSlEnKFBhM80/tNK0No
Lc1qemkOjCk/RpiegK3zfZpdnkgGur2t3XazbQLvGPCn1CDzuIUJn/g7XDpoxmAR
i4cc45atNDKv4D30vEPWdfaJqBr/jXJBlK6tm3TyudPeR6g42pBauS2UFtGjzIBk
rMUM7vO9Vb7OTsTcCgzsdLlLvQKCnisQ4B5X59CTNmTxYfQupVxq+ARXCh2p+gHe
Go8Bq0R+Xa98RYT7lGOldTpc9QGGii81GXuumYWlk6q4jvz27NaldNcgUJRFzvg7
N+tUDLcjexROOFl0NZCGAMgdc5s5LL1Qn7puIfiGOaz8DapnAPaG8Z23Qi0112Aa
ZQmQ7BU7sgEA3o7K1XbVF6KXun/bXoA6I+li8vqAE9pL5IYc9anCdWwixFlfuZ3b
AQH1VY5x8FmPl+X+Uh0XVkQKkgx/Wr8nMWh6zs+DisbeOrM0sfV5N07A89XB0wDV
XA7PmEOIWIPlKqJ9zLeMGuBbWxK4i5782WSXBgfys/wH4cHlTJm0mY3HvRcbBgrM
0m3TDocZ5wP/SpBtusCiC5q51U42PnJZ8dyR0/AwR4AhR1s5zWgPyQJyNuS+TFl8
SgeRWYY0fycu4650JUyfcsw6rxaGvTQQtaSWEfQRlZOCtq9+eiHQoznmykNvxJpa
mL8RkSeUKwaJd8BTp2xjsE4RZHfyRTiu0EaUsfoCeOqoog3jgBN6tWGsM4eY26IU
xCmGu61pkZdyRfMBWMPP2+mydTQ8xEJJiajuccnincLYa86mAnxmBcG17zVSZ6+2
XWvK9Il8TFKbLvKpwoHQrOled4gRN+MslYtrc2cir5+O+Yklqx5eXMUf6pI/zQP9
i4Li4imTklH9HkVdYPYdjiKbBhy2WkbwY5YCVqHYTkDJP0hMc/TsxcB8rsnzE9Pn
hKq1eWb+Rp9CTOb3t/54+q0tdnFESKAkicIKS31Y+oxXf+8B4ExcVximbT5Wicig
cMv8xbku57eWm4fHSoBhGhMqrTDwMZ+u02DMNejgH/TBn7mo2LpMBZVyyhX3Pudn
1SHsDNCthstGGgP5ud9IGKNa/Ac8iV928CBRTZGDA7u2B6sE+Ve0noW90kUQM6f+
jTrIMGQC92lhtFGhHk5LU46NVVsNZqYQRF+ccUT/bxmSpPIuSvJ3xTUpF5yGlWNr
2HYBd7+Qe8W4H/A5Qp/RLWujo1W073Aw7nd3dZBWIvw8lfNx2GVq3BVZWKt5yI9Q
4spPY3eOu9O5Tz6a2KAjVKNjcFcRofXax+VyPqjCpS8v8je1DDUhkEmjVQ/9UDh7
MX0yngAfGcEpYDrH0Xdx3HHY+TX5KKwRGTK5s0LmNxHBBE2bNQWJkjPUjLMK2/Ni
HvHZXK+pmkba7TM4CS2PYX3xxaKgVAkyN7K4Byz1NDfyVZ3h2IrV3aiDHSdFJC+H
fEt8qPBtEIvpYAffktD5Yi3ZmatoFUCKoDvpX84tkNgbv8YjV/FU1oj1xelohr5U
dxRyruem1lA5TCIhnzNrT/h8fjge+WrG7BuennK7gqE=
`pragma protect end_protected
