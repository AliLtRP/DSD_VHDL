// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:17 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fls0PLz4ZBsayz4YuXYvD5CqBA8q+jWHwDWV1zKT8upMHznVAQ605X1RjWsykt3o
om0wi+794RJbFdgRRGyv9VamCjlVxek7cyljPpU/l7O2K9fE3owx31fflCnxnF1S
GXRpxdiMLyMBIWL+a6KU5sWtf3BSZb9LlMLW2xm8L7Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13184)
4MOv1qZsEOKD86enHrVJjAEay8ReGmeokucLCcAfNdpgdTHvfb8Ct+GbUkq6zjpQ
oTmsC+QpPb4jxynW/yqv+bN9veGNjtMltgDbbTz6QAxgmhU8uO4a5h8J85i7zYSI
BBgXqHUiPPti8Knf8K+lrmlX5IQihAP2VYxB+P6/wUbnCRqH4ROJwQkJK58Imaws
f5ptr5kI6Pkv5/Jm30gNRiuYIxge1CWiWRTkWuJz3V6aqcRW/Ds2oU/RCYRxF2M0
2GfZM0dsJEtBw/i0tpy9TrUtyYL8vacrnrrTp5Tz20l9QdTiVrBqJUattkPBIPAE
T9jIX/hDTkCMwVwYDtuxLVNtqNCmQCC6I2LZJD8wis3hOVBdFczIJlQgNXrEm2TR
QOK505k+5JEGewva8oKGMR2Zq/tgXi5mBkk/9+xa57sL1JwlwDo0jqtwvyDZlLu1
dCx4cCSZ0ba7E1KvkweNEAi9w4HDDjXmAhngpm1j6XtyDrPVNFdznxxqiQ8aMkcb
SVgrbZKk29eBfPJ99famqV9Xhj9ZULInhLwMvj+wcG/DnmzjiMlP14sOJhcc0ICs
A+QpBFU34s3PeASKZZUMGCow8uibX0iVH3MgXcbjw8YpaXyvNNvNq7xnyhTrAtSF
zLzTsMe9NCcowHrWgFHSTZEkM1olxLaOucJROwv+ux1EGLQORxm+vLnfLNSBwtIJ
729Nc/SXTKJPW7PUskrJJ9CqVJRux85vd681jLRaMh53SQlKdqiGwy5DKvCP2gD3
7aNawGwgMSuyxYJBD8waU3jK9yN7RhkOowiH6PjdfqlIV1DP+9tYpga7F0J5SVhb
kOyCww0+qAoqDDD4SNUg1JuvWfZTR3ll596/mz+jjEhtVnJUk+atDlmq7bTwhEdu
VlwCyLQMABW4aMJlZM3cQlEiI/owEKeqVfvBPgCMYANQ9OsnBqw1pi7wDYYPEnJ+
n0AdIatU/ME+6oLeTJlsK3e1FNBhnZ7MRtPoaYRVpoz+W4p5SLNV7jJHSrmILKdI
tZ/YdCw0xT48Y1Abw5msvQPKklGDAMMkOqxhl1JLXJyAMKYXC9soQytXgovXaLbo
40EENdS/MkuuLufql2Hf6L6vNXHzumAS6SC2PD3l43en3/yb6RDgOXQiDZTIkFUx
0uhQeXx/WvxPyridFRwUa2UZzKwsUlpIM4c7B2MFwnYkDgnEPHxfqMPlfn3btqIf
hNzZc6R2H5gJ7p1JAH5JAQlDRCFpTlA4/vLXVSBQhBc0qID+yOEGd8fU9Ir/w89M
0ivTWKHucLNmXzb1V+Ht17iNPMXzxD0pT9t92TgZy6AVZRxueW2aDQ6vC4U/ACu7
YjfYT7R9doCIYRp1VyruqxcxmimXz0/CLsKts6vKwqRhDyCZEshD9rx4SbqaaXWU
4G5m/InN5Wfo0q1QGFarJn4Sqx5AWc2jQfrIG1HLPgcDRhZinCRlgyc+/V5HzxAt
T14mvj2flECI7O74OOgw1Sy35/iLZ86bpVdXoVyYunump0nOXPiC7n9wJ+De0vLr
Ibzy82afJhe58hu8SBYUzInBa+19YDh2VolUnnltOrMuvfysNtQwH3aAVptI4Az0
SkY8VHQkmz0Qy8zk8pGIRkAOPcttcoAyi+CnloecCvBU4RTWMYsKN032EQMZ9Nhn
hVpPHy1V5Ie3yHl8QSIid9qKM0ka/iT9oqml5kZ4yUwgg7JVdDmMEUHOxZJfnH0N
Ywzt5vSMY49VuBDKMqkiOwkxhTILExwv0kxGT2QgxqWOGX0W9fyEmsinMwFWpA8T
X9+KgvysBA8bhurK8XGWKDFxQkVtvt9LL7S2zY4TZGOvZtwINUOLc0J99+SZlLgY
FA89rE9GsnnePPTwi6t1jAbl4ulQSxnvD9VICRaSIua5Ri0ngBlK4bnTAUnbs/iL
8ClTcPFRUa0Qrx2jVCqfa3vhkj+NUHWE2BEm51+T+GzCbeU7mLlGSUxAP7+CfjF4
5Dk9Z0NVeIzrHKVVE23Ar/Q/JnCW4xL8NzNSjPFza8zSmVlUWipiR52M/P9sDxR6
77WzXBVsd+5dVKLJqHnyLQ4yOGpT/ZDUiQHTYHxW7ez6NlQdN2XyAyozXWhwJ5kf
TM9jYu8UzRSMNFOG4RhaVRoQ6rzubwMtJcsmhUrMrOCgYUTQzZORSM8mdUmmaY7w
NtyWUw2VGDyOas6taeSW4jfzY3TDyJ8jsgnIMm+7PIWdWcUiHobKh0u0VaVtKemc
y6I0NuQ5nuDslpCXPOmryinVVMm1bRYBbJGA4zlUDiDkcybjayYNSndToxDg1seo
vjZkmA2GLGSv0aaGKDuPZPj9BV6373FTCNvsKJnOyO3KbKB0ZwcDyUQbHZwnY6Q3
rCfw8izOFQ6k+q4rsqD6fTJPFrJqmSfpiN/ln+PFGBp5m7cvK2RImlCZKwlRnvvk
zWxFkQ/w9BJAmkaiIrTwT5XDUFaqISop4egbSC5V0hYTdDYPnB8b+6I71iUSg+KW
Kxqb1QmEB4//Y3/xRYGJ1MmTwKY7TlgIX17Lzp+4/KuwNr+PLAlcE6Pj7CXek4go
iOLEr+ECF465gCiXIhjLWfDIOiJ050hmpZIohSjJsM5VJp1xy23yNUN9ubBB6eiF
6seqHhL3Ki/CXssgnVfBVuYz195j508rGN2O9ou6kUKAjAF85/0NmDr4qZOowH2I
l/cmgQZD+FafH602KH1EVZAdGZvBfuger/GnPpecO7IKOkBc8/WZreyipCAyYP4m
/PgEh6XZb/mfXgNKWJx1zNstLtVt3QOVoN1R/YlVQFm1HceHUy37dWjnyKA82ten
je2zN8hjG3rVhbz1IuuG7WYMG0tqwUpPLOZhCE+BuAImV0npxH1UTacHn3AGA2yc
wsq1mif7ar7c0Ebs3RplCCAOlquxhk84mPgtEibgMT2oKc/uzIvA8whLXyLtYDHt
8bODwkg1P5UVxPrpmQNypeA0OSyJqXGxTIObdGSkB7SEiLT5oq2FJ0EEIC3KPmyN
08mA6TaRWb0o48XGHDd5sxzYB8st3h4y+yb69HAE7PoHyF6LOXGdXyA8ZN6MD+kZ
PEOrpUfPEnv92Rw2injkrMLidtIPITlHdxnnKywmJJ+KbY8ujF2e057QYArgxXQC
W9doCUPTrttPHcfZCF9erBaxDdXllK4Zbts7T15nR9eSkbaoNoc+xf01dpUb9GaR
yxWG8NjUmJ16mtlz0j38EW8aLHka2STDgms2jAxIy5Hq9DTfSGFEd/iPhQu2zHgg
7wEaLO3aKKWBpgdM7ddNbzbe8rR5GYlj0h3wdRyk/AMD5xLdIAYHma1RVGcp9ntC
42sd5CNH4bxv9SqdGilvIkKm34g6uLoHwSHmgcvx3IvVB4POnp/MqfHIm5IkLIS+
rznLz7wfDSV4KwpJW/xTWOhJkSNovD2IbdB/lr2B5Y23QyTBj+LK/IZ/sHrZM91N
ysGrXVpQakSjq+jWBBDz1HS6OQ9lb/fW9M51kUkMrR/MtvmLc3lVltgwQ47HL58l
ffk3yhaaACnGVvezYlCf65d2Sr37vCBsdhBvLGNLFen5pai07zyrjc47F7PVpoc5
F6172QiqrXUHQaxNLSaghtbFDehqr0i+zrmH6E0Mp6NYpLaMdpGuvPtj8V2SncXr
hyBGdbj6VmzkLeTS2gweF1FplpoBp34c4VZP9izKqwOBVNDWg+MxF0eE1rH+7z1J
LSJfjmcmfDbwq1RCUpEivBknJIo+ASqzVip6iqCl/k1fa1qzYqpMuN+CjcjYOJMi
jZe0XC5TN++QIfR4ZQZfdGtxbcN1vzGewxSWDHMwEmfkVQGLWMk1BrOSn2touXib
sFBXXOHALHELChELhzjmtvp0jQsck8blmQAzvZxGMm/vis9CteXfqnjgpGGQ69L6
V8ZbcdZYQVmjiLA4AiPcGr7EY3//YXqHWdnWO/IwlVpZwiCS7EGBAyeOLNPfV+Oc
X+9cCgaFyga8YpnTautTMUqttnACSVUODjxfEaX/JlIYJME+P2GhSW99kjA9UwN+
Zf5AhUNUdUpEcp5am0EA5JggTZxzbmF2b/QB4lb76HEfcn7TSHOhkFU7ULZxskSJ
FU4xn4Vi2+njJGPBS6IK3TTiM7dvGmE3S059cJA5lf+voVEwsemaQekCjM8lCn5e
Q+DQwd3DyextPSsCcdg6QHRoY2gSVTCP6kvyZvLG2294+YWu09Ha//ZBm2NcRsLh
MIJEgQNHxkJhotrk7WG2pJOFbCSaY8YoSpG23FbdNTJK2L0dRF8iXbc5UmEgR+mi
VFT9WqE82j254ZVn+iNCl5ybAfaUBXvkWdfmSgKdnNE7eUVWRmiDqOhTF04I4hNJ
a62K+OAKUdokxH3ZzKmQzWlz9btTkm1Muwkv5RoP+bbDB5M2+/EnOxk6pma5sLjy
DLNfvPMuQP3fH2ad2oXcAHZZcdbhkxqo/DfOiQPfJRWIXtDU5cmhpro1+/Jm3k0h
3av5ufw1gTVJHOEr7HD3mqDFtRfMwRvVhV+ysrTI1XPuoFIO8BLoCaV9uJXyQj24
FjDiZ561YqeTAn37r3VdlOIv6wQ55uV5alCbC3uD4zrqRI4NEIIluYajD7++EtmY
ITG6ctmZngkVHPk9HJqZrpysRANVXBBZ1frS44irc+svJ+QnBsFHQhmwm6DbbRua
DAcsZqLfQManuCCwEkNrkPo55kwSZQeDphcBs3IjKm6+3c/bwVVzMemFQh0gLjQ8
5SPRbr2YtIcLs6iNmIxCw+/bFwyEXHp9o7/QjDzJSAv3rvfFYBuzysdXuHq9ERuH
vv8dbFxj1YYx+rloSqPHoYnrJ5y94+NoGaQTSZfhnuNgcSl5/dkYZWa5+G/841si
VtD7P++ysidlqLaZ4TMwoG7CcARgcIUKbWk2jxgS7N/9MyzAb4BmFTbultPK+FGC
k2b/DGPyWhfTgo4j3tsUEn4jhM04FayEEs5rHjYAfMYEL9JOlKnulCVxhg2TI6uU
8hCCZpAyUhMKwiJZIQm3fRxQQK3nh1V5UHVxhCKGZ0w9zn6xDJwROU9idMAWklk6
QgkW+UpODo9VHdSf8VcgEjz20K9dpqDpJzTVgjam6fmqFWXXKf3+fBJWCgI2xtrk
1x5zMfWMsrHao1NhcmCVY8KnUGiSJs4jMtfV13slI++ovs4yWZFW98FuPXyrob71
wBojY+D2MZc036Ah6TUrtptuCuW9eLWLRu6toqMs419h3aIP0CRDXjFCjPgcEbKV
7vlDBY9sWWPFfIsjkBoo4anbmw2r01Ye2KNJOGsnRU9SFJB1YKfRo67ZWC5IYTpd
sevqB+IiUmV+FKLNuh0A7+QaWDDw5G1D+TDtdL9PsgFjzHwdVA8vRY3sS2VVW8c2
4XJgW1QfkLoTUxSccr5pIpyf4ULRHB6PkOn+eMQ3MmxrXN9qZTjfwf8OEAi+bShp
pamDWhrDWN0GeViVllYJP62Mx5HDLDHfV4FGFQRUiRSectJljEWXJLLWYK30X+62
l4f/epH4Z0JybCD+idz3tgG3f2bm3ZiXBUEKf21Cub2fgY9Lt0om+DGhnx9aqeNk
lfy5toiSj/imEAcudsklcdDrJT0jpqZRqenahqIXbw+ZHCjYgzq/jmTb9HZ3veId
1vTJDQnG4WKLZBD5r+UmTUnPd7ERpXqXERY+q5cMGMZSrK0Zwa4Ug5TMt4SBWCi8
SwpwvlAU6Kjwj5jfMLA2qoQefarDGvXSBW/226V34cfHDVJBTKJAbmXjs+dsM7Ek
P4MdEPtwcpeSAhClil/d+X5x/X+biKuHcv8H5J8STiLgAt2jsRSjhpUyxiXS3+2i
jLaUQL+nybW8NoYFoG1Rt+xo8+/H4KnPfkEpcpRwAbiLAI24jT+R6EaWyNjPGDA2
TxJHHEed+WKXfrFBkofOf1CuLV1h34ao3+vPsE9Xkzo+hYXlA44OJnmFhcJ7LrTw
5xqjOu6dMXheuZ+UeSU47VsudN7b9im9J4JLtCxvhxLOhVr2CGk84X4VfcRVifUN
mvg4k8u5xyMB9Ko5zqIVu01VmYXQS5IQmSwnVNz8OoBsnP1Z9RvzBcAGkFaH5iuJ
3QzLYb5VqMfBTjkoKumPh9e7ar/xGf9AUgzX1fHeHP0YWGQ28gmecB70llAk+hSh
ckOIjj1Yz2/t0qT1IW3iJFaynUBzN/f6TKWCNS8blcOlSrEQ+4Y676759D4vGPKu
+g/UW6PIL5RjV4cUBVsvKKxgcBgHbe/vvqoHw6yB4qKDfiFUVS0Exyfuf/EQdQ4W
NGoooz7QcgHUb9USL0Z8aWnkwwzyfePz+iC+8w+/STvjfUcAMtepyrMtdN1VVnnp
u46p+RSOMIDKTjUEtmpNfs3JubE/K7jTLXgZtl0oDPIrqiVmmj/IONK2wvsw0LrT
rUVbkuqkLprY3A4QDc7y71/0NSrnkBfi/JFYoJ+XPEKq5mxSoGJhBMPNytNagHcy
1Kh4gS6FI3lBOmpVQTyv/gv023KzuhP4jlDFJfbQT8u9OUVJI5q73/KLElkT0iR8
c3cYm6ktgEPmCshM/yxUwAgJj+dYYl/Gs62w7tILDyaYXwHIQ+5uB1EupELkhTRx
gRmTpc8/vui0cHKnTH8Ey2gKds8Y5qp41LcMP1A2dqYoedwfcBymyO8daPS2im3V
U6o+vDqk6xYg1w1Nnqz6+9Mcfm7oAMGN12OML2/cyluxGG4I2q9VywWPlsDSNN2I
Om4eGRyIpnRre8CAvNmYAeGXiu1L/wPr3qPTHy0BdzXGsy0/kJ8RR+KlfblsI0Cx
ZjiVMjSpzMqC5/d3fczYTA/nb+B0EUhknpmQInA+EBAUMo2b/opL0cp/rZ4MPLeN
M5KavRFgzly6d9XfQzWJe8yLKpD0sYXYrEKl0kNCsKq3y+ajIuxj23Z0XW330lnS
HxdcLryL4um0+QBNWVPATRdMqOoGj1girAi3F5d0ghbQL1zgWzhP64HEPpwlwSSu
YCFrKxWgoBlUrW6sr81mV/TZMxPolCbz19PrdpPiSLIioNFgwvgEIf1vSmYBN/NW
+3vILte3y04+qTxnYoczc8uYjkXAY/GWDsozOlFpixT+jBdO9qje10CdlymwVEyO
8tZnImTFvMIi4O0T5VBIS6wF0ktHHQkh9IwxT4AqFrJpS3UrKL4H1ZYHLQedIDb9
uBnhmjgFqQcQRgAEfFsL5zKKPgeZOShVu2cmqIG9tWZ9tmHGzSJO0Bi8H7LA1Vm4
OAjWVyimmJUoLIicA4HC5Ci5xRMX3oec4Knu+1Wl9RUoOeqPoChLKbkw6PoyFJVl
ZK8TD5GC6ckHkwocO4xArL+g3xFvJ/NJwty82gaHzCEfv0XDdd70tB7Mgw125Kxq
D+68se4LipHqq/2JXEsySofN36SX4mQYkBfOqGnSqaj4KcU0ua/ccM3U9mGSIwtH
hrlJgKtNJf3j2/oq2pm5Oxy8vi//2sWVmvbOHuwbMd1ScvGPRVP2BmQc+bcV//6J
1Cmow62xw6yrRO3YJljA0VAdGSCEp4XsG3CndVrGGvpxYRryw8J9H6C40uepafQt
/lQslbUCN80aU5eFEqd8SOevJC/94vxKy5JpvvHn7fGWivZQQDC6gbDBK1PAgU6Z
ZRgJ+6EqhmsD03het7ccqp97EEXQbhp2EqMC1v7/sBUmo3AGQ3CePjyf0f9v6FIx
TTZYCdG4VW4bOCsvBmKX8pFDoCakOmivsdKGBqMgdCLnaKDZ4XtdfH4X9RM/HM9a
mqI/1KuptfBrfAhwHA+E8IbAE4vvwbaOHr5wvk5GDUFCm19G3OrpEOx9udvFaFHS
FrNqhcH8dgDZDHlPjqnLaC4H66nY/W7SrISedXv0oX9UBFkmC3l7Hgs/8ObOBcLF
TMYl4COuYe2xxqUurwGQlTj8/3m6XkQGXTMUkUwCVKQWHKUhkI6tZLaxh+sFSnO+
EaYE1DcHSaRcUNVB+qEl1+ITL7cA3JX2v0Nl8OxGV91+ahVAzEu3QP0EuqhFzKsZ
9K40mp37/u8n/GNFWt47I6Ku5tb/oaueXr6s9THso9mmgb5OkZdKT6mvln/OHYmj
in+cG8rdVEaciv6qn+EkbSSL3+DhHeVanj85RQbStC8VY5W0VQKp8xo/9b5c/tFF
9CL4Yy5slkFFDTM/nwY3nk96Qd++r6PiwzNV2DvvOUAPtO7+nw27Fx4oNnPlZN7k
adCUZeDQJNSQYuH/Xcopd2xRc1z/hbGgaCI7qT8TzLLi7Ra2y6mwbR68c6A99dSl
8WpO7YBgcTjkqP193bBO82O4vLw4O2fg+ZqZ7w8ZTR59nEd1Xq/tPV8LVz/IhRe6
NO9S0lALxuggUGsllUudyIMboTPRUbMjlg58FiQ3tW7X94lJxlqt8f0eWdrBdBpR
+woUkcm7FvE3I+lPitHP/p9b5lmKeDf5eDzzSIDj4+lGRk/L1gJpbi4j1YQuKa46
1YYELQfJnvUQffSyx7Nt6ic/DHtkYk9Fzq+EJET7hqQ2jo/PxcvgkW4RZy0gII3h
Df98EDAuDsgAEkRdDP2j4YoxSXEbRw0eMIVp/23NNa4CWJYtvIv2wykg8HlpMH4Z
ArCD65cxL005/nef+wxR0xf0ZoBLnyVO8zkaejd4S7APLGWaIbdS+zULboTEZ1Om
CsPHSyeGVwp6XXtPmMCOB2LjAMG8dd9GbGhaIlUYlSO43nh5A2U6X+w8GwLD+qEs
mc9hIhPmbtyFfZryInumcYeYJHQhJAKeR25B9LI71PQbLpxer4/8rAE2mp8krary
SrVGJK0GgXNA41gc82lG5+WbpfgZKOIOD/zSPwjLCG/bXEU+tn5qIB37djalxxs6
aNgE88+UEywc77+OiRtrBgcxSmLxcZCc/ebNEBoatrLUKvJtAlB+UdkFmXNyjqRe
WgF1xy7k31UVmmdpGY5O8n/EkuzdG4tCpWvECPHeG9Cci+0glKp4RXAtaLN0n8hc
vIgkzUmak6GtX4pXImS0cqg/NldoN6yYCM3bLpiugfcw481SNbkhdDFGVOiHQn1m
12H4MssRkORmZL3HzILnrHmp523MVHvng8SuxBY0XNDECc/KHrFubmp1ct7XCnC3
2NLSEbT/pDbTFPMrFDjjwgZoKltNnzHqcphclR01t8Y/KGb+yNtgDHyoiPyKcOxf
doH0TwFPBvSp29GsdnDc837xfPCO6jhBPjhICrER5GbkSTjkN6VOr92yU9VVxSlv
Q8uGsdtGkn/FfL62OxTF/y70tv0ZcO7RIlukwgTI/ZE1W84L4D13jYznCn581Vac
y6UK/oZiNUlzwKZs7riWvIlfE3Gl+BlTzeAoggYPX86gyFvWRmM2Fs2V1I6pe1Y9
ItRdMvFYrivKkg3R2vIKdhth7eDBB+5MeSfZnayHkyr4TnvCyFMHAKR2tEiXXBbU
v89Jk2wW8hzjFPKZG6t+h+Z0KGSIAVTeFyOOsd2UL3aiLYQQw2zqJyDBxFJYTTQX
kYSEBrqT+WQhzSXgUEfR2c+nnabCMVupfSplxdz4xwAAPui7KvAiyJxtT3HYhvi1
Djdg4kVKb8aIoB2n2kbwbrKozpQtxGyz8luqQ2e0nPkPZB0VhS7AT+hjv+mjmGdt
oOrh8iEP+gtKR53VgtLlwbEkafeJ47sKUV//qzMccXeSQsuotptTMcoq1FNL4XTk
a5hnLCpWJAIdDV8ZC7zpH8T7T5XxohSvByXlmdWalWn4dZkGttFASn8hcbobaugM
GsZmz7VSfKEsE5gtl83GJ5/RrjzOieqktESQXjCJop6epiVfisxp/C1SxfdJRHFb
cq4mJuNXgvaGsiukGLv/al139oCDVDxU7YwJQg4GeoXcsaThjD3wfLaD2bjkvgoM
u/9WDprq8akcxgL3GsZRcTGYkyyZGPqOHn/j2nbMNUq6PrmFxHOTtbHl+nGcbQpc
l+mlrPyWRssuH4TSL4uzNkG1mF/hG/5n0pJGb0BgXpilcKChN2ZJ9YFU7zZOxm79
sakreSeTog233SBcnW8V/ZHCrOGjweQVtkBnZDzIr/qQs4L5U07jB6MUi/E8+Tsq
bxyiVxAV1RXbhesLwW2FH/cwAnGeKG+FzOIH1wULqid58Ya8GZP+f4YKDxDoxk0W
60smC+z9cSvJmcL0sctnLrOpkI8x7qjtnc2TLyXpvLfrrxGfGQPQ9eCMTYAz0KOL
ludEk89OPWr/+mfynFe17cgY5810lP0w5KHFFJvq/7i1xQODN9twA8cUy9NEb5NV
pV019y67QSA8a91QtfK5qE8ybDx+NnbVxm0svxrz1ID7Obq1lM+jcGLZKTm4Puwp
KL/++KcnMXR9u5YU3WhXBNONM+Pe+of6h774jPCXHN+8UYqQ0b3r/xSx/KHTMpKR
lxj1V9SOdhguRcg9yM9iEoIj+J+VlWUc3jiQsLOypfNPeZ+p1wPIgiAkFgLyW3Z8
MQht3AuRNlIDE4FrBSn17Nao0HQaGGFc2NWCA2vbDi9Y9lE3R5p8zFH5OnM5CFZb
ohEo43kdTEu0zwFzWTlb4F/D62iwd9b1JTMNTa3lfiqxSxuQjJKqxnqHxvcFUMrl
MpiPQBAfJg51X38/ntNqhih8+n0R7PWum+BO7penMeFwGbnUuqAagbZz3Hya/J6J
mIEQ6qYs3iubU9HHznEhjntsXG1rO9l3tywE5ssr7efwEE+mu73HyvqpXqlC7XeP
RB0zuvotsUtah8JyVi+EigzNTO2cdg0uJXxioGmLUbZODZyo4/REieYpbp8ZxAkq
mXG3eP4yadmCPEDhb9+cEUgKGDAyDuu+Mqd6sZ7pw74ciRiHC3+3sR7ffqJQyE/v
wiAEoc5MH9fNYRQpA95UwcxUHuBKZ4omBPEPOcTj9IkfITEcW4kf2X0CrluRTWJC
r+7+iJnfWgJ1VG8/4u9rPr5qW5VsRDPCl/LU8/Nkxa/0Ed8zyRcqiqv5LD7KpoX9
jzhcxytRRau1hacy/aBjEoP0pYSTZB/44aI5OHi/xhU4jK50cnuSm6gbPkqQ0mEb
MLAMQaa0trS5GctGvK9M5x4Is8M/4jbwsJFAnf52VzC0mnEAZxXGxnjE06wdCBd4
oHn0gWU8seAaBRN1BA3fbCDEiJ/j89S4/Wtli5Dk5YXgFrBZ7Gd3D5l2erqZH9o0
lXV7v1R7kTFNTf3cuhH/3MC1yhL6gG2dOIZGtTJHvxEdGIR2BAFHfgka71eoBeVc
3znUHJnhmIsuHjh+f1nf+rR6MmWDIpgUtbjVNm5yn74aB+S0loKj0ts0DEKA2AiH
b9wTQ5enQBOctyxp2Rg67A0gta+AmzTuZKrP8K44yVmgnGzqeTaUNEfRtCa8K7W0
s0bqK3L23quqbfM7vEi5AJuAvrg1ZZUvTu/ITlkgv6nfiw658ljkfZv7yaGZTr/n
aOtGKwxaCbXpu4EEMOjOX2N9eJtXTycnKKn9R8a3Mic/TlBQ5L158H8CwUbZMssz
FmspJy88kf33Fpj+nNHSmbYrMzaE5DkwggqZEEs/SzroyXBaHdDOs3l6e5GtRidF
b7aIoVAJpJVea1uELelwqB+o6OlAxaaso8nJlHq7QLtOrBMeGRAWsG5/Pq4SOoB9
loWOfGKtlm6DuzWhW2had/6cld6IKv8kbcaP/NhMSU2eu8dzwG6afFFVKuXGFmoE
eQ7yCfZWtEmSUD2UmjBOtVSHbN2OVPlm1zcaHNbdPjE4gecLHsX3LTI5rD+MbXDY
uHQxHftgZUssS6C3UUvVzld3gekvPeVotGUSJBcmo5SlakuEtGIhsPsHac7GahCn
c9ol/bNRRAcnlWOWx3sW3ZnR08WCraN4UwLs2U5PuXeu4XEcVnBhj7hp7Ir3Ldwx
Fhop4PvdKMHr1cHEDiwMgWgUxC+K//hJddB5FW817ePFfhZaHlAs5ZTqYdXRbCeA
Vpqe/SpwtJm0Oz1gpCx3eFcDp0LrTU43pSQIxBwEP+nVml7F0TTuohTq0KEgUZ7/
rJMFRQSc7g0el+aXIwXs0pKIutFfx+oyT5qnRUB43v0JQs9kv+7UgS1IlkcLTzlB
LVjwtsRtmrVRIf7e4V2o0xY7xiHET+qa//6ods7JK55gjMyMJj6N9WY2kjSyiFNw
NqnVmqYNQD/TkinrnbNqLn7lJXIicmhGNiuqRJ5pfz0DWHgibRQoaSY+JvA+ymo+
g8N/Q0tHIeDhxLj2YdRzf1MNcyfuSCOWrUBZmFv8XmatoFsZfkSCFonUDGvyGaE/
z+JpMrsDXcyBuuDYUHowY/qiEnaHHWg7HxRYXdPJa7cU5StkjZnzfGa54qQpHoDP
VAbvvDjd/sh8+v+b00gV2yMM5XYOGl13RRtwbJPrynXvjUFdCBEuoME/Dr/7Q6lu
Ip1HUoSgdMnAZIVbQatc3jeMZZHG3ONy2cA7aJOjnHlaPFzdEjAOvKnatc8kTofB
tewbuixdDLIGZfncICrqfNQ5D81zLy7L9bR0E3GKzWBRQnaenRXaFNxMMUoePQ6W
rUOUJt7J0+c3iEXEFMXeH82CTpaWpsO6Q9HMwmwhCNatxD8s2HGe76/DXR/5uc38
EeDDfx5ptpH0CHNxtQcO/OF1XFpQdNEoTarFUI/C96xur1UMKwb3usxV5R+yrVa4
LtoPYChasx/MbkX9RPKC6Uj/T5z747NGL7jnmU15fL23D/JZXhajqxNXnv85/tox
7C3wgKo8h3ewslXM0wuaNu8uIErvQzdmb8tASdudKuVy04wQdqYiJIfF5UwIQUp2
0iNStS+bJQoWYgwHrvQP9yhdAxNT25CQtSPITXeoda39Z+TvA3KIq2wwQTtb2dNv
1SOOJQvKh5f5Mo9ir3KbHn7DdGjJjRowVGYyn5Ex5SHW9PPAO4oSGz4Kp6Esre+Q
zTHEOlO0utVsHoYF8CfFlPhR1gqkqC7aUIyekS3Dk2lav5en6o8Sa03rvMVw+rMo
yY4Dq0PI0XnssA4zlclcNQY4JbackU8kTFlZGDiYPQP6+U+AdZTfLJRb2ZhAWtiU
xJ1+6ETtL6zcDFIzHqlIE3HOkdcTuUKc6IQA/l9aOco7zgP0nyMj1y/U6gLDEhym
nZ7YWYM5f8tGdKteaL1bt1Q/UQf0AAPrIybmvIuHh+QcX9wMYRXd8nj9VGbcL3LO
yHeoS8pRObhOZM83UYPo81Sh51TQjmXp3ArRqxXOLZ3AHZtPxZI3XcmLxY111lWr
pJrv3+TuOS4QGPF637rR/aXXyh7744FBs7U9K3oSj9f0CQFu+01LDmoHirZuFXCk
rIz4hV87oCdPvV+Fvpne9bYN5QQT+ZwOL7WtgBSEsfD5eDRmjfdTb4RDnokpGeAa
BDvy0MciASpIWm5BLfVBklBCUb29lbRNV4hod6C9Zxhe92b0ReeFPM2UUXXgQUoI
8Gu5PRSySwhpL6P6P0H0viVkjUIcBnZ0NhdJc0fW7HE9kImjljH54XQfA7VH+wI/
3q25xaKxx3QLjlfNvQHz/ENlj7JJdRK04RdK1HxWi+oKXS60H4doqD0icpxDcvE0
IRK81ZfBIxevP91N3Qs1JbhLzHU2okwAZBpXXhOw+u1EmVoa+JAiNWJa+DvZf/h1
Nf0MKdEc4gmAovzeuIcGAoZ9BIlvqV1/L+aINohPD5b0HGPvUpBl0t8o3srCzNfq
OWchuhWMVemo07ofc8Ez5nTTBt5RDVitsoIh865r7bd1izlgfgQ/+v0PVg2f2ezZ
DJygLUCYh78ehp56lbcxVarjR1++EX7eTyONjjJMf34RGLfqcDbbLuF0hyDHkH7q
4T6yx40fKpnsv5qNhBiBeTzgwI2o//vMGm4mQ6iOEQaJeM2okOppX3XNKytrilTC
sTN/ytAHPOfwDl+M9B6U1+hdqHWiPoRx/3xVUUlR6YhPgNbUd7R8tUA16XbHSFBn
dfXahCzBDsO89bQuIl+pg70nfsgBgdZvFiJEQ43WyheuhNKiTaEIpgocSf+yd58Y
3kISOnzPbzq1Bh63vg8LMxehpV0h6eA5diS2VfSlndu7w2QgxhLtZrCxGxYsFS4H
E/GgE7K9Kfz6pSIEqtSsM3usFzv/+whLgjyYxowH7gaXDnSFtOmETdEAB1DibdBE
OmQc2x+/TOdB6LYBRmroKJeBnSF4ltUy7r4fIZez+pqDGeFuWeJhDjjJxgNrFBOO
NPY3GAsmpbA+YpVTQBgqxkB6R47Ea11fqiwc+lowp6bmT9DQP9EvGa2iXkIDubsj
aMdXiwsrWiF4pSbI4XZ25BzTgNDO6yXt+fs1ADxRZ7etsgJ3ck5RGsAGpzXr9rUV
hICPmoZZRxYgqERgzK6SrSyX5gb7rl7ctKtoM3CZ1yqiZi32ZZErH0zys3dEK61C
uUdl7F9KJYQf/zTaT0d76jTou/s+kWNtqFtHr7HPj64aE0wxH7Xi8xmzq+wK2mON
5m7Dw99sy/X5C2yg5JUxNd8V+grsJJcVhAbab8t00yXxvZ+U5/yfM0cLqo8tUYqL
avoXatkkwdzrP1SZJkPVkAil+DitOJyBE1XEAe2TqgR6LM8LTrVuCLSqt11whFNQ
MOVk2hLw3XvyWZwPMZib0gjOhdkn6vQFUKJIC4PjuGi08xVuePFzNBeSdhOvfgfz
GS5afMUQsInUD4xNbA/ngm2Oh6vxf0lzSBd1caRTtRBIrvjcefarEFyMdViTFREX
/ePoUy6AW4Os4facGjv0dtuxCpWbcrqvSGai/Hfr0sE6QlregnCtyuuTOtJyjl67
BoR2lqcyiAfb0m9V0oVo00ls8qG5oBf1FPGbEMS3wGxmxUbCufBd0cR62O0yyIw9
eAtcBx8oDqX8fDPv3qjz7bAWMOXaZ8hw1Q1MObof6B6wXTtrl9Wmeq+qG4EF1FRh
zFv01Jueu51Qc/3td+LzYzV64Nh3YGlvGhMqBCoQ06PO9s1xGtZYnfjEU37fMZWp
MJfKEKi3Wvfyak2vtW/r94bFyX8CuH5IDP7Hn5EEWXo5fwgK5L5Gsb7cybhgYuCq
hgGVlldGrt9mFUwh+X7enDOZfM7pgZoE+53r9vHIT0qbfncY1HMJdwXSDsRsEoGL
aYbHQls4f8RHH7vT9M5E+36HMFbvCFpL6v9kBjb+yR+za/UBnU8FpaePD6gnDaOQ
iETEMA5iAI2WrQU9MfCnmUII5lYDE5vUMq44Cqymn96w+hlVlJjodNeAcMrjHBow
IkeBtMftpKtme6cfciv/1mg4i89oPFI8KXXfhOKcmdOOboxukKM78mV8ykwlXf23
0QVsFX4YoafFiJr8K88tRI71lJwrpOtXjYMfJ3rDev8bNx6ScmPvGhkUBr0vBUT7
mxYXU+n/VDxx1HwJ0ZoJqy6hOCjrNqdRGJHRDKgLGrOUUcK+4Pw5GAI4KZoyR0Oa
RdbgxuV+vj2mkLbRh6YEw1WS/EGl7b7i7SPyYLlDpmnBNxyqnt4MrT+zrQkalgQL
/QKQmLsV4H3GEU6XgOdkPunFNrPDosXTobVPja0qL6O1lvnHohjQdgsFeTlAQdbe
CRJnbHy9p53/1avC9zB+9QLJSJc2vBbHTFVM66kZRGtN3d1P/BAEdmcMBBQfhLEZ
AOZ8LEELxTMPMul2ekH2w2xX/83dLWzAksF+sSSwm6sL+urYosiZsbL1Vz0cgq8A
azfWqh0ogdKgioXmCuKsh596BuZy92MWr9C30hFYhta8fZHT50jcKdDbERU35Dgy
xzHp8aaIh27gxw3psuUrCjx9Uthi7DS5oD3je6yKaht7C+d4XvX/CVEl3XqQr2Jo
q7q+qwiI/GAE3TzLqzpltzNlmGyrnnKZWfIRicZU0Ug8aYg94iiy2y1aI5OWamFF
pFJug6oK7de/yCV/sr/uGv9j7nuHOAMJwvkjayNkK8lYTCtjv7ymEJ+0rpR12FWG
t3RaD/5N2hAUiv4o64APF/VFcxsy5wBol+YE0lCBRka45QrWkWtnpL6qm0qEeUAi
8T8QSe1SGNSt0OIV7S+rUDEpIDrhFN+0OKOvZuE4uLrfPq4M5UyvLpEmqa2pxjEl
nKNTScQL7NuMqCLCk0Px28JmPHmbkpF1FTJZjwctYVj4+Yeke7TReDPzU92ncMDp
B5M08c8LZi+kPhd7S0hpA8sm9izUldFJEEJfiKzzn5gc7V7W4oFTi3FZgPkNkMrO
iJqQJpEAySuPbSIG53ZBqLugse03HyxVHEy0Onz/0FOWioShZAtEg+VKzfiOqcn+
yzn55TvbjbwJfeAUS97vRoGNTIRGNu1hFib9E/SZLQ3cTy+EDJOfT84adulAtsLV
4RauPpBZ/zT5C/I+RGTRRMXrssooe6jgsXJwN0QKoKfkqYdvmbSH5SFonp8bW6dH
1542wGyWBgVG3YFVx87r5ZhbAo/OFDXKfZ2e5rWMs424jGsw4jHKQ+1NxsIVxXrF
jtk1szLJnXhwynSrkpYAqF/sMOPmElD66qqQw3YOzTK3vdbGP22JrtaGj7kQC0Dn
O2Ovf2QHHfib7YV7m/h2mouLzTZFl/fFQwbYQvikDfFWI7Pa0XYUPGfir5Zv/Rfo
qJl4Vhp4BgPDgJ//Bc380QwGlUaOkX9Zl8vM+N3eO2EPKd37gyLdskEz1oVxC1Pj
528+f8CLEYDZsGwGW654aTBwjSwegps9iaXCfmMfba1ui+mKJuX6A3Ov6E5YU/Iy
5wN4pv6rvz2zL/cxSukazUQ8JWODMIhIBL7Fun92yLm3ZDrVlTP+KwxcpoDVcWCz
ziIqMY9V7VqZu2PYseVPddcWbdwpqzxp7VgVq+8P+ox681hmelA4aQunow1eobvw
h3bukKPO7eBlo55cnveqR8NAmZlJmSP7e9J1H6ceArbxu3Xc7jTQINXJUWumHKTZ
TiEsnCSBEdCuPjz/9IZ1ju7h5CipwO7MkyNUfGRCgLNj0fCIp5iA0hTMqlhhPIZE
H391zuwB6wyfItQsPJZP4s+1C4GzK88AbpU/3RZSIHR70pk+B1o7DdJc2DBZ1QRb
OffuPPrkrSBRKp5qVo3FmBrLGYxXRMEAjfuymeW3c+qnUR5FMk++iXnPkpRFbNTC
e7o5ZtOk0FN+tGxRZQpOLV5kChA3VMc3I6Nu/GOgZmVX27ynG5bhX0hoblCQv4Ct
9OM0ATU5uJWI8MhHBj4SrA9XtCKIqqVYygzov/18BMBq+ykYobmcFxAEoXzWtH1D
MOReAVdek9h0qEQjMjZDpBhQOJ+OJKjdMTAZ5t7P2tlhqr4811cQenKhW8fOXsw+
BnInYSGpgxRzxN+yUXrUX/WSVI6Pj7meVwI9/vH+SVQ9UdM+/bpfwmFQ/t5Aqrsi
9bCGfxYaVsSUjvfyXf+lzT71dcTs/lH3SsNgq1NS3nBOtJJslxh9Ybg3uhAtwGjS
BIgn2M+dEoidhs/VHpX0oefKXq6jK/qLwlUAs5Yxw4Fh6W+mRXShjethLQODf+eG
0IDYeO2ZchjAunLmkODeUoh7ovWkjJ+A6cKHac7y2U6xWtRBCYwreUct/f/tiQy2
firfPnIPwlHpC7kWkY0LNfBwORDSyEOiwfJ7NstMwcxo95zMaubWMqRYZoUFzwY3
XbXjF32U0amqt863/Q7GdlY1mF+bIwdnGdUUwKJhmoo=
`pragma protect end_protected
