// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:23 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IRRaBvPyoTKo+HyHpUm5d3Iu75lc3I8iaDyLWSIZb4CAgeqlt5liQqSVOORKUp+G
QlCRJrRy6LirE5zaa1AtsiikMu7EC9Mwd+7FR4juj9GzXP0mESfBuh0eAo7TNqnj
oFnocVg0Mqya+FcsLBl+9YpQRD61Xq4f48MdykzRCd8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30640)
Lebc2I4KzFKuv0kg7OIQ4CPruzwAvbKsIfkgbqceriRX7dWDQZaZ71MVVXEQjTtT
RwtULnsh+N4/yZqAeeK9hM/WAvXZze2r1xkx0WBeAfB6kHGGIv1ASPD5G2ziHRax
AGdamj5QU5qWtDNxIKKVCmQCL9misd0Bdb79E2WHPfFRGo8X6LGbwx2hfXEuEVP9
y5MoqLLqHS+8mEipH6EhLn7T8OS9+TyKjm8+7EfaOTRtscuYNQB5pmF0YXAoYfwE
TXQSEMByfy+8oHbIMy7CArEIfNZQDC7EHji1AI8LM+yYpFgRFtoVpKNOB9ZiBLJH
Bksnf/N++2CNzW3B8MacDVsqVPzjGdEtWkG2nrPnhTxNmD2gJnaf96G4zTh/qbum
j0WC2j0G0GX8jgBqCyY7KjeygjHUIsJFD33JhB08hE8JUgmSteSM0ZObrmjYG5tz
Xo1NWb8uEFQxZnyrr1i4SV22NOJ5DlV61byLMrSyNJo0AbHkioQRLnMQiO341xvt
q7QjKKQdwqTthPNcClUXhEzu2P6F7icMc/o1xtDqm2Rc4mya5H5ToHoMns/vIf5Y
IASLKwo/lSxuWuyNzbpO1XjaaBDGkp8UQxOp6SXUYiW/Mv3d6BrkW5nDcNS+I0Th
8nP1r3V2YqqLe7LnHtYn/VYOlVX3BXZe5yPppObV/c0liUO/4gq9+S7cwPwFowC1
K31sgTTHvTK7CDt97tuD59S7URy83ie5vI3YkVG+LwwGmOw0ogq/vMHDsav5L+6j
3o+PWFfHU7E08AXZTx5SKE3Ic2ovc0uj/9UF7JQLs8+2DVeWjUsyrgAZ43l7+gbY
K5EUAowsCL4W2UR9tCfSUG1e6Ya9UfQuoNcdtLFqao6tWuYtiqdJpOs5i65QpSNm
Z8PN99gC/0wNNt4c/hREp+5ZNXU8Kw57j6gnv8EyYStEA4QuWaYFuYWKR2h8fiiP
EnT/WoELu8pxdd3CaN0pf6VRDuWDvUBcpK1Tzbo/hVoNYU6fUyyxD+9hn34Dpikr
1ZcTEiXOXogO+G6WWr6xyuhw5hv1v93ekNEO/xvzYZdR8HMlCHbqlNTGUTxfa+cQ
6GPfkQOZbTThNgrvlL19ly+2o/lqezGGXmy4CNUno0Dgu2ysc+AaZdCgyiUzWjma
7Z+iiNzYKzTVMkNWbQHCdtraw5NVKjZuY070zyNQhIexz6xlj3u/Z7IPZ7CdAZH2
yLRAfS57lLTlio0102CsZy8t44KJQ1H1TRJ6HrqDP/j76Mtxq3t8LjrpljfpF3gt
ut9BvnFrut7g12xHkNWKjhFKr0bEz4iay8K74dY2IepQ9JbblXKAq9OQLTZhceaY
L3yOO1novWpr7nKzlmoD3u31Qos0G1oAKpOSw3NAUtlw0h9rIlY7m4xaQhshS1hl
7NHoUCY2BzhpPypPjQ9+ICqfQCamLZhEKEQl0N+r6AV7+Zy4rCRAYXcnc2YaPPbz
8YeIj3yfsHS8JryeeuNrxpnnOfR/pHHCjwsUGP8fy2SU6BOIfKfA93FBDPlcwqfg
MViwgLkY/CSB+tzYR+LzS1yMhmUwiXBTfOJyKHwyG3NX5r3kYFyZlD1DV/pW7tZs
E2dksx1W7qqxGx/qZ9KbEQTxBEnvH/1PwobdQR2f72XgK8MFg6cr3qLwtQ3/2pbQ
Zlr5UFt9UDeyI4RYn3mxLSP5vnjBWoEJLgbWl5VDE1g7qlZwctYJ5YF0xCrEW4uO
L3BrOSFCt+UkWEOQjPI6Yr9pI6/G+YxTifhh/VjQaVYsnS80v/5DAYsEO7O0z0m6
XFkyeXeN2hqUTOWYNjzInOQ1tJ/duZ8vHk3ANUDDtMpuWFgN1H/c1tLgZnV2ZHwe
UhOk8nBubywv/EUqPxd0LCTpOa7AUTqQRYEu3OC3b6tYmwOFT9aH6Urtl+DIle/A
UuCdrlc5joqf+hetYiFPNuBfa2TuMr8W8diGaQbQDyjJGues+CnahUeb4Kbmcwp1
F627iY9DzfDKlHewbmgigTeS74yx+1KQhCZ3NDUiyuUbq9ED1v1QKiS89z3mxYOF
k16QEz9upcMV8f5cR+uVjcF2yhvfzYqLZfZqeu9sGwHOtHVWwXJIfjFUw8/0LL34
Ylb8a1a59U2VJYU/eBOGuehbXiOC70qEcuf36g21taJhoA/gSEBIQ1/AwxsBB+Pr
niVhdlZclKiHsruBd/xVJ56byKB9v9iWVPiwwHhFCyb6D3BrffAQNJErLDbmpsFv
YBlj+4QEF2IlQPBCICZAMUqPnKReIvoUHGuCYU1r5Bee47gG8cgp7yo+u/KLVL/B
WtMkrsuQfEulgEJoABgZzyc63Bm5qZCcjb4nz0yiJHXRp4+4C0dNBOgT3kpKKxC7
Ru5J15n/te8dszVVmlXtwc1wCfEitsvPzb6b3ClB6fs85mj8fpXvqSkY910QGDT3
KGzEYlsJFIz87gReTAOskdX8VUvFXrt9YnJys+YiCmwCr8+cIsY515KBwFz266eL
7ZG7SC9JPFJLBwxvA1H5N/uBibJ60cFQVn3nHcAO6wKmTuAoL17XtPZ2c0F+RgZu
2VmOZSN/E0Td520dxMro+91F/kmuGcVDKCUUan3l2HGK8DAFzchj6bD1OuIMpLHk
jKtvvWeYDQqVgYhL7P6+27Lgw62UWmfnYPtt2MgoiaWgYQf35m+nc/vN6xibh24S
MwayVb96DPVjLIv6UHdUmoQI3ZfmXhGxMdP9cX6io+qv9GpGcvrE1bU8p9tYJpPX
IbR5yWnd8TveE03SiUAoArq26AfHItFqVyPw7muxcoDtR0045oI6yj0dKWTgZ9q4
zDUwCOlGOt4q8VDjAKUeI3nvvY4SiYuPu+xGpXYq9o8ODVDYMccvLjuomNuX2Qb9
HkiLT9OUXUsCBpIdrYHPr/rS5mvgJCKp75uIUMAEhueQStbAiYQNROjYez3Ftnf9
/q/1irq6pF0jpMiiIrQVPF7w/ldHjz4dVuO9/lRujKZnrUxg52JG4RanVqewFGno
Z0+RKSETVikrCFhBswAaObglnCL96vBa8RcPgglxcgc7DXYi4FxDxLI21DE7LgbG
HG8IZtu4bfavCW1R0CBG9fdPM4JLkGZWBl3EshsQfiQSUaa3840l6DKdHclnFQ5B
Yx566DwLcUJrtTH2v0/wihHwVX5n1Y9vsJ2qV3xAxoj7C27/3gL7EHuYygjPCy1r
VEgMndT8pzDwH5kuLsVYk3CcQbYv+ogcPbHTUqdvOJvaAUnoJTw7R4DGGW8isnk1
tJXgwAY73sTH9H0lRUiA5AZHUPcetM5dwRg8+u8bMhQRV4798KygS11NAlZfPj5h
5toUsAQTlySnyHFcx1y20AWBiDDuTgaH2Eh9cyN42tb7mk+XdMAYyW+nVcCIh5On
u5ItN+l0atUcNHW6d1Z5ib/BUq0kZwP5RftTAtr58VsbuwBF7Zcyxt+i1YpOhxC9
61vVpET8C8oAZxdDFLICOETPyVS4O0omXbCF4P9DA+Uo0PCKL2Vy6A2H6F365aui
LsWWNplrFaAxguO9+97cgp9fahE8tAw0472nbbEu4KYEeeLJSlAzi9b8skI03EUd
1qz2haBL+OuYzxffT7mF+u4z4xABNlXpyE+8HftAvnQ+IxJslqmM1Mp3zABDGHtr
+W4bGkX0l2+fp6Ljzkq1C1Pw1tK8OobLN8h/dSD1OYdcspNpwAp9S45eB8kloBpY
Y/9mSIoE2HMrHo76Sa2Rkw+voV3ORO839DFlVFsvlL4HoF9+71IwdE5UlSX3A22b
PcDnRHMyqCCZiDtndVzKU8cLj8cr/SOz5c4xuJITt+9D2Dsyt5ZiRxwqKSalPK2X
KBULQZUV0A04Fu3HaBp1admXdzzDJVcU8FUajzGLIJvSQOY+CqGho/YDCsgq/lXe
HJ44HKot1Fxq5DI4z+idCLPKKF1mGx2MqF6fS93DA9t2w89Hxf5WasVSyKyWkBZ7
OpcWp9MDEmRyXO1ywhxTPXSzPNuaGZMEMWkwK5fqLYmvBjopkcPe3KoY9qPnCpUx
GZG1k42uROHKZqjEvNkvEncuM8H3EHHFDE+fu/L6z//ERUQnTeas6lYpbd0v7gEV
afTDfq1Ez+lUCipxXM+ST9t7ctzOgvEQEye50YzYzOAhvkigcBZuoJ6MFmoSeIXt
pJAVF8Tb2Ac0ktR6rnyLHkvyPTPePQhKvSmBTm0lpmdcDXEDdq3qrSPZfYL9/Zty
dwFJAJr7gev312u/i08nxOEKV/S2Jsszw/YktYbWTJoniKuza9CUJm6aMEqTtfUQ
gh+t0Mm7AafzRmUrxctjyLlajcErqoFwUn8MIX+F0R/+oTuGk5wu1YDOBjhQnasg
YAISqok5EeCZ3IK9T59eY3vxi7RLYn7AEb/29Q9Nv0vupb/QexwwTOBJDLMD5pIS
HsuUFqGDAk1/W3uLuzVAIM82nRaIbvSQzQVPMx1eVI7owtiWyEDAmJdObwHMcpbA
ubXLE+RyOUfDKZkgqnu/RPcbHjOO2GWct6eywpvrRTov8GMzBy1j6o2XwhAB7qEe
wRHd4cKCGkMzKBPDS/qiXl2f/Da4KY+wYmWJzEyafO8OiiRF473aMJRNp2qPPvPP
/PGyqCd+c42jh+FccvLAqqs/BvE5oU/MW5jDkSnVjGuwdu5RZ9Irvx0CYPzpndwk
sZMEf/QnV6UDgauWSsIqcrGgzRIWWP02o3PqV9r89bBUiv+5L8DuqCzeMF8/k80x
O3pP7ou0cZ7qUdRYLC2K3rLZ7z+cYHWTHgi5rbuyicfYjZp7PSwbZrucVsUwYLVQ
AuVExYstjajK3dBz7I4ducXIarkVmsxW52/u/8TRGY/IXlzKgqVpRVP5+qd4WIp2
yKv8Q+Mf/PDtrgzznOX+FjeiERo8EenY2FmLzlgucK4hyGkVVi24IQbODW23pamb
PY567/yaSlroUV52SSertsvQ/7gY+wq8ZeaMHhUdFOa8sGjzwJNR0OmgQODCvCsR
h/xk+farG4mLTLuxuF+ugQW54xZcxQNodjw8J+P8dMSgfhNMex/FfIFVF+W/osvT
Uo/0nMIsYNGuLPs6WaRIXIKrONWbaAJmxiV0b/fI2Xo1b26uMKedlBX6ilaYz3Gp
X3BWqfw6RITOlZP9QclGeEJUQsP3Znoc03Iwhf6gDqqJh+/i7oqh27yVppK8nFpW
+NYtlQ+4kyyxH1q9nZcaZc2g6yUOFZEIZ0enUAORpI0NTJaB+35AAAOikCoNkJVD
OuSK5y87AFkXFGukH6OGP9QTXKRRM75qCzoykMwTHCe+mtzpLKn9ULvxRZvkwiMC
GgzSosfoF4Qq6LZplzBR9nFTiEZPKHPi+CZExlDXUb/HChto6oYzTwORzYXxAHxu
/nmEqKR6+ltmQdVb9q7DuvRSqTsksQ0HL33sPDNaoUWUtHQ9392W1Aahr31dMUjs
GCxczPWzaZH4qDUmK7EPJLN5EQlcPNOAuw8Cb5SfGGOdnC0VAmwmloMO/NafBywO
Q/GHOcPZtLy7efgno26nS0f60LAlsA+TodH1l9QIfypfDJQ7ECnzOMlTigDKZDAH
uLXrtRq5S5Q2ALLvqpM9ACWtJSuTt004cAwJLwENe8iuZjbA8W3adabNGxN10qAX
KO9G+S/8C+Ol08eIBsy4vlXjXWpm3eOhindbkvl9kdgpDy+nYmZCZqeVg5k+AE+s
mgaX9sFoqYYldeiSbSRu74aeTFXF8YZplfwvuovcUgeyCy1eAP9Gqr48xs9+Ov8z
umWj4l5fuaDMLil0TasKyn1vpnq9mFU+DyBRBvu1y634E+YvUPxEwhPDndVPYEu+
+EuYjX25eJ+sjFWRA31I6GpWDRMu3pMUh2NcKYwxiYN6cuSB0WEwGFquEe31752y
7u6VQnspJHRVWQZ1PLvLGD/bUQEmmsed6ShBPAhdw3MlYgKcfoKm0zRW4PLNAbgW
RdmI479UoMXBKrHKj673YzzSNglFtfqRYROVTYFAqfs++kk/v9gaOuOTXD5FDdDZ
82Rnjmxclc049K40kWqHddgxE2su6mV7HrJeUvDjRCHXa0mWVsqO+DeeSH9MYBJz
IX7HOXphG4QUoAs3Le9pNLbAAJ0KmEQYwntG4rRM656/adgIbg22lMEXqqS/Ytr5
KcA2znl3TdnP/6ygCPkBxODzqxBXEiM6JWVmP9Ferx1xkhFSgzcLnO3wVyN6oInU
Cnn81buS26ubX0L79uCTR9R+xm1aqYCcDI3If3a6u67RbCYc9vABoPBUvd4giUQr
rOK9iDdBJFjVQlIZPAlE/ROyqBQqdQ2o99NJDQPqfaezEFENJ3oNPqArXZdiGxX/
CH2Ravs5hSyclh3jZKI+FwuIutmvMFr1N+hFHGUYboSDoKnggv6kxqJv9JMWgsuQ
fEabgRj/BqJCvuE19IWkHb7LSjJKHM73InFtxTgfyS4QK/gcqPfbUeoKo76Mhq1b
Tfglp+pmQtYCaZb7uDAYE+JvODQ09QPjSfUVsI3uFVKh+ymU5mfQ1ea5aDYTAHX8
RQfpSdbXgttQ7T5zdElZa22HGDoVzRm2d9GHfy/349R0m3aW407TehRYF7yED9S4
2cgmGKX5KOigAvgMYRp0TIPZAMqGggEopVCJvqTN78L8or/ARNQSN+RET+G4AQ75
2QYxh4Y+r9Xkxj0uoU77ERJtVglk/T52f0ue66Ic4wI/1XI09lcbURoDP+erWPp7
h9j1TY90NIIkEa952SgjRX7iiI/POgj5Rr/bPCSBxhF1GP0pxiLA301vodTemzVc
Xs4oN/pHBFqFZ3HGZKc9bbvDrVJx55uZ6eQGPgSxQZsMJnRt4lBFXnTc+vLnEzGi
z09DfvkQkJKhaJX0v99p2N516WMSuP5COCraqufUXOkHh0fgbpjOgg4Ejr0+qnlm
vbUbnCenMo+SGPNVnRv6kmAnZ+gsGNqfZQexlyHRb6C7bXVDatk/1k6Owg1PPBng
baOYKcxZrTLXN6T72l3AeKMDd/noYL8bzMF15Xm5Nz9LCsURD/YAleQGD3CXcv7B
fIfoexsWXm2fg+ZbT6KPBq3okjg1Mp+Vbagpj7fMAMzBqeoVa8MCIQR7ZDQDFR80
2FeICXhrx+L7eGGB/KUhxouQG5Z+Ll9noV3V3G+NQaYuy5Xe5USz1Qj/sJ5FQFse
fc3D3QxoUCB7ytrINNTqFpftxnLlnr1WUUUyl2YB0+4/mTu2+0V4Hr0ZaLOhoq5h
ckNLIMHIYJK6W7/rc1BwDOoXUlvROoByFGcumwJ8s2MKSPtj5qLkqbbqUCo1tJyl
LnDR3JnhHGV+KJpN/GXEYgusWoC0eGQm6mEjDAvzDCMG6vbwAkF5G7VVWeafdJo9
jijkTdm2S7Zlv383aQeKEPzTPZhmEd3NdJQTXb7StBn5P/g5NrVq4pLbRkFha3H/
/apr8O+dw3M1EnqQyjHGcrXGFpeh/05B66VSBdAu1wPNuZ4pJ8lv6YhpYDN7yKz0
4tvFWb6jko7UAjfhHbkpc9ejsIqrU2iwywHZB8IEDtMKmPEvOamSEHgzD5a/FeK+
sQpgtcDv9cjhFGiqhxx96zjeonTn1R4xyBpb3hAiGvZFKVrqOPVPjMF7wQqg+YLr
+4ukJIRAACEir2KIU3WRGe+dr91paxtyFaldbiDEgLZ38rVMx1DHyqO/ZoxWHhlP
jtwdzEphHw4n6BLGBT6CqtCmdP6jB0Vx6clGXlWDUMhCpCkDaVe1t7G6/WWFm8eN
6HVAWfDc1uu+BigIglvAEwGr5iUIQ0xo0rA5gKZhNFEDrstX9XxK3l4UZVqarmTc
fU3eoo29eVbLJVjach5AEMOfsCB+UOCIlHlYD53JuD7L7mJqoKUmv3idkOjGKiTz
TtmMkfcS7KERvmDmCd4URkD7ZyYRI6y0bLOFn2uBOSDFpRkuugrWnbSBQBlZTeXf
wY8BEoRDUqT8dzoRY7eEfV1E/OfzXdx6lv0FF0TmvRQeEVG7I2NGLro5iHmQxSNa
XC65SXK25BIXgsIWUyg6LpSE3JTfDI3v7eI0P18WO4bkOwZBzW2rgWy6B1NsfZSP
PxyofDC+fN1rPcqOS8N7skHPJey/L+WVaxSafYcvJo+mi4TkER+cK7gi3/1T4ZZS
wmZyKVENXcxJsKaXfwR9w3y2fX9I7rjEtR1PHNxorpkammDsc356u7SQR/eIs7Tv
pAmEntu3YHe2/COweQ27EPH+VT2Zk+OkxuhoHZ6VbhI9aoPLSr5kiYa6jVku+SBk
S1Y52FGC5RXqb6fcrNkY0iGWMFE0kUeMT8WVBETlSVlGyhCzow5P6hAEVFOfHvP/
CqNVuFsfnKPo4NLm2DzWUdFslzhQe1M5bK3aQQSp3b1YQQZa2ufgZYqKcwY36eP/
w7oCHSpJhhh2vd4jUy5GLFz0tiUg3cimVW2EkP6SyVlbiyHQ0nMcgkkc/s5H/E1C
1CCzqpKqrvErP+tH/vXFz8utZA587kMqxsgGpqdhQuKZpEG0nw7ZF2n29GLbLnnf
oegx9faplYdtQKjUAcEHxlq/CMnPLU7xDSCBaHmXCpJNGoNUlmTrHYctz8ObFo+O
5fGuYqmBT6M0M8d+UsGHDTYCvLbEhL4L2wgioi9tGZ7xJMef3K6NjTwWbP9SO06s
qazBHKpkvMtJs02LYqtM8id1cV9cyj6+XccChdNVdiJ9RdL/Qrx8dQnW1kt2lGLH
4eVn4naikPUTwyFyQtVWQMddHYWzlyJOgrsWuwOrtW42njrOTfWz/WX2AiSaq/I4
0j8cTVFZqIgtqTA0ajgN837dl9v5OmzWcZKcDYtYK7Fra1ZLCu/KR+yZfE8c26sp
BFGbf+36wOh8oUl48F4eTqVviI0dZg/63XZmhYoEI0U2D+whCSVv8W4GUHAwhzHn
lU3o6yIaJyOYmHAX4+RI+ptAdV18BCHVLyskAKgRBt0TV3q9bKw0y/4jqRKwJZYy
iOBvkPsWFJfkrldcIMTPd37H2+i8ElJIZzuSrG3+5i4pB+RHVWH1PoXx3IN2QLry
RJ3ErxaNsjwsO0B+jNgcYgqYAVLEgVcI3mnQLvFrh/FDs02MVQQVjbkSl3e7LTkP
uqJsRYK8SPnws6WI4BSP+QaEDxCzO7iWYxEn+N80hjczIJCa9KOsZ1FXTLJP2AWC
rqg6x/LyiceZWt9z1TZdj06HQiUo0hvjdvbeK7VcPIHn5r+vXazF0KxSDo4K1tnF
yJvxxbxgVANETvyG815/EodenJHmHqCt657J33/6hHGWQFTujvnjVi8BYnDYz4ml
GP0YDJnoPict/BaF5VF7G1hiIOMg2AtdEWPpm94dhAx1eOqygouOtA/oV4+bLuOO
kIDqKuTUVk8NDYiVH91fnDpY7zjpIMvvKk2yT1kGVOg13PncqoiJQ8IauqQtT0vK
RBNKNGR+kbnXUX6sGHJZZ5M0sbwNgJlwNS0teZCEJRPJ/Gnd+/DzzYhCG76y64kB
8A/2gP9dPtGHwVr5ZSbFM16/qS5aFE/hEjDepJ0fhBlcfPpfpoFWXI1hHsm1RkK4
Pdem1K7Ksg6FLL0Qy3EvZ/sRqedx1lEyY33wyqa7MdaSHRg8IL2qznr/ImCJ0oFQ
T0DdAcEymGlUXwyGSWyagLrMdj0wPnzALYM4jSbtNHi941ldfyKZJ46nZll566aJ
MGGNUPM9xrPPwArXWUlcBPvA1LVcp8LSBR5p41ADEQYK4AsoP47B7/COyMkhkp31
xStmWQs/InDYxrC2vk4M/h0cqRGK3/NX/HaRhMzeE2vXnJDVMwvcFghtITX78Lm2
4rf+XKYFqavCpAU2zJ8hN+6w9mR+wg5tBWIN14lAGMz5DEGSdTtr6I5oNE8Oq45G
lpHp5VMMfPJ5BGby4d9xp7sotI5peEcsI9nPNDSmWP9mpXY6g1fHuLyKLrosv45D
fznSoZAa7SkMVz7iWekmDFMBFZTnWxG+R8TDw0mYpDyB7NYGC1DkPWqTxzMqiP+z
aswlCOgxwLufqRl6p57So3cK46mX0Oyn+qs/PZCD+4Sr71zcELcIzWa/L1Oe/ZWn
kbOINXgWtZZi0kVwC3/Lj+rrBFOu6r9qboUo/s2eW2uXnCM52kDXejxLOP3opGsN
18iyWeGc+LE/3tos8vT0hTuFYwp1/OYU7PHCdsVstJUULlQYuwKUeiaN/CThTk9V
7dHzGOpQ4fEa9TEE7I0ed/zGrfZwOIGpdM4fvxebGMWjiEdtQsrrlrPnroMGJ6NB
L7im0gR9M7RhbHC5Mx2yOG573mjohA53h6F+O8mV1fHuYH7OQM2/osMvKfzyCc5X
F8gDulrSe118AK57BIr8TcYWbLVeqvDFqJzgTkkxY0Tfqotn37ohOdDg5+ICnKh4
RltBt+PfmIJ921rUx6VS+2HNrMgXmc88Qd2kjis6YhfpLgHcwZ49kxhbN+OeBMAd
QLaK/Qgq2PN5JGVnVi96RdgRlEDNDXxdy4ZT3BCHWG6iXCpO60Q9ATiSqQ6+sobu
UgIjiZtZxsEBlnq02MtJ3g+X8IKAtpzVPeiybPyve9gYBKU99gEveEUo7/TOC4+8
B4inBWakcqSPNGw+oKMbyEkXvQxO2sIUUpJFgx/xYOAP/sC1oDbSLadUj7px0y0F
/DlSLdgLfoQ8eBwK3pSdlsZuqRxaI0YWv7pzFiIwXXUqgLl4M+7cIsUhEosuLW4F
xyR6TDCdKdInqxKIwFxG27Nx6kNJjkizKbeHmOgBFz2e77SIimfnZ6YauY5jAtje
rudXE+ZjyflrClJ4ikSS71kynVRcg2FZfWAXKIFkKvxdueU+u9TOAcRb/4RUdk0B
+88/Fujw3qaPYRcrYXkzwLiGxkjjKJfDNLC+k3JkNEtaVjOODVfjM5I4G175GgZ3
zcufr+zae2lUdZT9feN/iC99xuBiI1fQsK7DwsuYaJSBlHw3PWcjuayFCC0Qj6wI
6xXixe9f4ZraXWaxBMfEJ7L6kRcRz/ovFIcgp6b0Xtq2T5VwwOfg9om8Mv2Aqxal
SwKHw0aNVQKBQpxy5WBcY1pgzSDPf/T1Rc5KFFsLIczfV4zMbkzujN0xk1n6PuXl
C9p05Mh40iBU6qoUi91+NhKGznu3GozAoTZGEr9NF8gnaytNpaFn7Gg6bOrNczCW
9zm/YsnPLSZvSfCAptiNluHFrous376WiWvIxhsJge/hfcl6zM72vMlEECs7ybnO
KpHsgcRrFVULObgNX2ge+MqI28zzNWXrn0Lnq7n/ja0Ox59EtyGpAo9US8VWdBNq
3CyuGuZzU+fLfAKxBjhQQSD+ctWXC+BG8ftDxtORNJtQ3BQkdThh0JN8zhBJwxFj
ZXBIuTZVaK2Z/qklBCRZfd+CZESSnjmhINM4cT36237b/LLL85H5Mw8Q/twAM7S2
ABfOL8VzcJ1Hy0HHFpU8Bn9eDUwJV8XJZhjo3xyt/sOvsCA5gXR9sGLvjvUd0qUu
DR85Qig+xnbMoor001VQQOp5KX0TZn1yv9ens8fBGbmb3arrxHh2qrIe+84flfNt
+hTrLiEKnz11UOKZaPfJfB25TWGZi4mN4S3p1HUGpyipDPF+slKtg+Xb/aUtRb6J
yvKWuZi5k1FtWEOCFhHxdJ0bLMXFC7Rpzhy1567Y/JK4R+0Utz6pLPuPtWqpcDOK
MNiokOJPbmdlIc6aN8iCaIag3Q8ExTEP/WKOTuXcV1M1AOwEtxRqTKhL0FAbtD08
aCcoV27654iDlcr8emEMkcW1D4m/ql86gzOTRNCbJa9Dw1kZChO4HLx7sYqMvLuh
tM6ZvmiRqRnMGYkykf6iMzswN5+z9Orm0hYbLoXlhy+ItG9PQTkxU8eUFrkH3fp6
PEfKZ0bA01z2AX+/nMMhxd+3X+1umLFlvtozW1vzDBaf3rI361OqUhhVRR2RPSA7
IGWddvpIS/7GIEtf8aB5QS+eKxlsRYBeQwUB8BySVYkq0tLzzEj3A3XnTx4rqdCs
dfd/LlvHt5tAPLgBBmsF0yP3QzL8f5OfDNOSfaszYOSafpUTtewXSkC4bWOqTCon
PwdTJKE6e3066l4yV7RZ+IABpp56QvSUb6YeR56NJ3bPYRKbW8zxNCjwRsAVLOqk
T+DpyE1kyZgHH8Z711G4Xj8pT/9aHo/tnnBJNRPunRv++U7/jZdDMtwnJUQF/wdt
xgRzsoCCsHlvhJrdAn4lrOimC/Q2UuiFiCjCOgIlJpwy/OlT66cBz2IkOOZYnYQm
AVgPmvYdostiBLadOrp5opsUycIYsxtcpvSm400juCPm381oEHGwjQU0jSFEGtC+
JCfms3EYRHYbTQxrgL+WZJdcD7IeKjFtrOjiMC1e2jSLj8uQZcMwVl5xH7wGOHsE
XQmUWit3N79dXOZfWrTvqF+8rV1insB97mOxpI1Ky1Um07gAiwpTpVNHdqgDq/9Q
0jjl2HP+kK2jlf70cgFnW7nvjW0DmhiHYIgUCrxFENDan3bNGJfHys4SRylg1rCO
TNj6mORzF+tQIlNUp/xRJckAJ4+ghP12pKZIhLDVdUiIkGtL3g5oaTqQjEaPZYAX
VfGcQRp/7zzfAZB/iMMbfHa1EPdPGWcfSRTw/Gd4E0XPo7lgufsdBysHzIIBCHV/
Lq0bkuXeAX1pneLdSQbhi8GEqstu7QfLcVPIo7zV0TVpcVdryrYo/sev1jdFq6Ny
WhkPSpfytw3gFzZoYcQP2OdJvRY/ijGMtEPReIZJ6YddCAiC8jfmSsvubo1j4KzK
ZDl5vRnLt2Ysv76V3BarmQp1FoKnlj7OCs0ufFDl0JWQa/IpAhHdC3VtHlnGTzHw
M4VmoabIaCViHZnfducYR9qNT0FF/OVDFiCFT+Sk1vdMJIAPOB+H4f1ixk4+xOh0
pwCWPdiUgn3MU03bCaOjnQ/RpCLY5FZN0VvpQAGBIFq4KjRhT/ZzWmHDMaIIjHE8
R2GMnOx5PjYKknlt/9JJFQlpXu7Qd4WdpIp4IAI333WY+Dnwk57r8CnnQ6FLW8N2
/zq4N/34LO49H+zFB+PKER91g+V7ovhsITG/L9uoxVzO2+xZ0mQUDry+QMlazDqS
DVlX6PsLbW0B7rltpMcr0uEDUC+bVnpMQxr87uJiiUCtkfaLfLLV8RclOIU59ln9
hOxwOfPbg79m3jzFW6ETX2ET55J1Z4FiJ3HrustKRL0vPjFWD/9bjB3WHCPXQDw9
LusjwLGcJI0milker3QMj67rTscNtjG4Zkj6O+zx5ecZjl/iJXKJd7IOAUQlNT31
tBoVE/AL/385LFq8lFrfV2xZd36Aw9Rf0LXqYGbqiEd7hvX4zEGV9BTm3lkOIGxG
ye4K43kXMMztIIjr6I2uHAK1PfCwGclCA25/XKrx7115NmbH5UTA12rIiC0jackv
j0FZKYGhrSaqqWf6QPWlWIkyQUZ8wEJRDTRKK58o4W0bkQJlxHJg4rF1AXai8asQ
hG0iuTk4iD2OsmKh+ebisSvVezAu5GnBkhAtTbxbCaqeGiDyyqNGd2UCT+dj8R5G
ot/dmQARjrGr7TmEx7TMdOmU0Tm+ppAZ1JVqpsy1FzYi+p3n2yNkJ7wtea0PN4cy
2iS/ePfz3pGQmHi9woK0Fq1KMShIiuz12ULejwjaCrEiP6EAFQcZoR201F3zhzrK
z4rjIWLC3KD01k5tsh5zWKZ1LIsoDqqmitbimsA6GbX0cSwaVM4Fdd03FX6ADXFW
JBoKlxZzr4a7iMp4+zulyCGaQ61rg7cmC2DbOWU5gXjJHELPH6DmC4WEUNxn2xYK
ZfEp2A0DY10qbk5bUWxOykd7/s4Q7DUwKD78L/WGBDLqlLF9RkMaLsZBcsoAxOjl
I1HlPlAtskFjA22mzHzgUsJkQeBSTPq8ZdhM/59lHdlhkJisRbOcs2SVj/m55Kwk
0d7pqTWQvUZ+tJ4kWB5MlJU9avzdjD9j3yeHxOD3PQoCQZtiQClYeniRexpL42OV
PB3REa7Dk9RLO0wLcMclQmkz9yaFVADPL/TE323s6wiLpo86CQcSX7tDizdaJLbG
d9YpLd79IWYWkzYMrvflNdtDxwGA2X6eyCpiWYEmxotCofrDy3fdDXnKurKf8wS7
WKEU0ORWYsshWU629wX47o1eOI3gkprILTcqVnxQGNzt+sSCaI51LyIvcMGd9gHI
6DoafYIkXXLLPcd46KarurFYuR7Ilhh7Ffor/CQ/6mwei5yld7IgzMm1v3hrNM9L
NESg+YSflOD1uNfK7yht+tGP9Bi11L6HVEBSV0cF2Vs1jU1rMWxDaFAGoVJ2V7Xq
0R/oUyQOkHunaH41iIVoVDMtOoMhVIA+iEdqlv/NxD+/x4SLgy5G50zrxKTqDZtm
oxxTw10BRZJckghgzkkYRqXftfMNxfy7BB72v/9fgxBwWjoNpbF7lc7F2OZDnfC7
DBNqGpc9TiJxgJNWuRlh10j7MEN+hFEcPOrEHtAJ6LKMGxILhX98ad4w0OVBmXYK
IWLUlNwHM8Xt80BeLF23ksLRpC/KqU30PlAy4QObfTqJq1kauignNuLWBBzeUh67
iSKdDGyO2WlgoHHxn9VtOPYTr8QCpxK7+0yhnvHVfVvW5lDU57mVK8T3KirO/RSR
RTrHZJdq/ELTwmg0indR8kKCn15cBUdqXHvPLjAP6n1+25JJ3LPscRNKMUtnxZPT
gWPSRUfobAxb346ZOxs7PTweBfQHgecqiahQMtngpQfcNLGbTSZ5XkqxUKLXVPMy
yxiez9r9FLD+XODXndVOh2xwg5YuPndx2xAWY34SovIgPEQhpw250N8sY5DcfUlx
O1R+UzYFhyoWHiBQlFkxV8HKS9328AVY3biHMyUdL64KY5iJiRTAFbwt3Nt7R7oW
1AOgbVR/hJ8wnS67iV/fAitvQ5RwWHTl8YSO8+CirxTA8rOAoxhmd41v6GfLP/fr
GckgXPyxelyuXVDU0shVakTCcSC2pZ5y6bEr6Lb2kbGy43V31pP1x4OzyqxjOT54
yrV4zZfbAtjx9+oZj5mMGSMUNrA0+CtRDGZ+J++MhyuVEQ8KkiW/ZZOHQIVSWiEn
l1986gWo7JeBzOV9Q0dsOxeXq0PCd9i3sYWj+ejiDd+Cch9b+/1byxJsMd4dqpy1
aRSZBW2nVXUHCh58yfGn27Q4hTD5YUVf4fLWa7okuP3xNETMY2L7Poy5rl+HMQOL
Wa304Fw8DXqnVskneO4B1MzsXVeAMrTIqR7kGVp/GkwzkhdKUgDh9k8rpa5pUzUv
FSUDvqIfzfrexiNIZoheTFY1pd0gEUfP9+hrT5qPtGy3lZjCeRXbx7ESzJbNjJBQ
EcyriGENFVKv3jrVkxoSQChQrwZ1WXebFi29Rb1fGQQopOG9ieIegEYHnp6MC2Ic
A6Sv4wi/B7tqXYuf3hp4EorcXX/M0lEdRK6jO3EguvHWtVTsx8DKZtJs48AnceB7
S36iFG6eGjIlx/vir/8fpkBgs1HmQyJYI0xC9pO9s+G0TOCnoSMKol+cuHk+Yue+
oQM9b5AWr7ds8t8g3iCeYvgLfZJAmVzomGPQhKPZMbPwPAmrVPIef5PX62RaAqMP
k76nyODMZT8D6OSFHs+9KcevdcwtaVildZY10NJwG/Xv6wnVw0yWW/BpdRK5vBme
vF8hFHZyxI88gXaFIVZ28bPY7f4zli6t6lr9JOAO/ak8/BuCIta5ix6VO8sPQR0D
f1GkhPfTggev8No5c1SVykCgDL2KdcQQmN/BerZeVLza/oq2agossP0ZRtlx5sRx
nrzQmzodVS+S1RmZQpTrUPDIJx65HUZrcVvaEG+4GrfR8uSmNpJKYXCHRtZz+uNg
RiYisEzXI/m6/ts33/yhg0oxFpgCZ+G0FiizNBdma7PUztbBQMmLtaVgw0pSI06c
YjbMCxF1s8NE4+qWmdociTT83AWpJIaUS8jB1/wzk5sesYMPyHuWaegftPvNCg7r
vdzh0o0260yNEs5nbzku0Y4UIS8XXSN442BAxzHzvC54c7Yiw4IWF+eB12Gd7hrt
pe7P6FMglrx+4vBVCb8sne5Or3Oxxce6eTXdP+r4hcY0ndFKYWUv8CNrBLFmbuZX
KAp11zqXrXmTz/mbwf1MIbOJp4248AUWFgehdO+kdYAuzWGZWCJwQgJdF5iusfnH
Qy6jh9Shylnpe7018cOr2QL4i4+fCYTgyT/vSpKn0S20ay7Fijqq27T7CbEOsTP7
kQsakLFDAwEIjcDmJJ7fcgX2sr9zBtAikU8P/4+GFbxtgxNmOPQFvlSNxt/b5j/t
GliUcFSwV/Sd2koYshrUPcuKPAcEAopKqsNpOh7OgiBoaS38G/3U59a60jpEv8G5
sJfpVBgRHeuhY1n3xed+qWWyntlDj8kcBLuVsstOYa49NcJzaIt8A7L4zVMzGeAL
0/Y8GMYv3Gttb3rCwdF7kFJoHdNmyGYodjf6MPbfgiF7zoKk0Ecq+cLAiFWpCJrB
mGoDcZXdheq+nHHQ4vP9kGfMD2fmRahS8VE6gfLfsN426x2yi6i8aps6P59bfb/U
oxwSRjHdYmk4JCppKxtxB+M5VbAxl8GqR8McELVncBdVaQgmCQqi5DJQT6yiRmSJ
P2RGP17FPN1YjtpEeTTB7CYBrVVNqWr7MF1GCjoJmztCh5JmqkH4C6me39b4uX3I
3ls2IERtNTGmWreJu/ui631/RAP+LL3J2V/ckqdczAgCUQdKdLo1P7fSKcqD63YR
JWY2DE9oDHyQvfzO55V5/Xwfo4dRLwuCkpHAh/kmB+zo3nMvbQRNOghWhaSnz83d
Sjtc5zTf9+emoSEPbsRU+c1Y5Mfko8lZznIA2MhZGLWZQCBRimIrqncSz951qEiq
m3OifL2YminFP/8zilW/t544xvBcw3IqrRCELAE+TECvCb5xfR1zKBDoJrCZTk6z
661ZmVv3IV4zKxlcEHprmH7f6Pg1svIBLH336CwE5dKj2PiPn5Iz7wTmxnA6ETvo
T5y+JEIdJ0nyd9KkmIO8C2Up3olGcnwSHKSbXa5p42tQTsjRjrMkpjazHbSjubuO
Oi0L8gCV1Sc9v9ryYVI7fnJJyqIYrPDykeg4VIvhtEEnl6M5Jc+zV8Xa8GFbp/uv
5JP9OlJL0HUqGxTua2LFibXkPKHEX3/TmP7qoKaS6hUk7fHuC+Xy0K5ss4NXjASf
NU9X9MzK0mV9wy4T5E8RylgVZM7yRpcxe+7Ms5HwyNtqYy6qWbxKYBNPZFGigeSF
vOaLXJVf7Z4ts60yO8OHtzQALddQUatX4AnKa3AqsJsya4iHeGYtVc08/EcTW7El
O0Zg/BFg7cLp/FCYFqFKfqqcEUcOCbChaX8e5AN57plv8Oi5CPtp4SnaZdDzpf0/
8y062osJr+rGtV0lSx8IkggB3NPVJBhhIogMaiR/ovJsd79KuvP098ETZ7J8KRRY
nM5mdWY6KBsTsEfUY9yyXC+rTIP1oGcZAk3ikcoBZJssWvXtOjsznI36RLK5eI4Z
4dKY2TO75e2mL3+Tsxn9chZn1O7kHq9w2z7fdfFp78qdgueAgDQOmi81bg/zAL0L
UV9wkfEkoQuDFHkoqgyhQa0faLPYEEVYF4b64A0Hv7Z9hjLn+ti44gHzaAMr+HHe
+7+Qi5AHtEMQE5WT195JcSZ0aRrg2OzyCTmD9S96a5436oi4Zs9UUoRchoUwEYAo
v2T5/ct8rxsPR28roI04b39jMGefn0HwJYXXn1kNaN+SE6y6418iYq0cyICEt0an
n5jDZbuHaH0mxuQ+cAMJ5D311n+5J0IynF48SuOiMYkjsOPK+sAAAeCc4/eiITbX
Dy/CH3jtwj/u8uCo9iyjX1vR3xPjZu2KoWqUozpWXklhtz657wVFdl08K0AEaye5
YBSY7zuwC47o2/sdDgZqHsmOizB68z1HxRwVRCsDJQOx7KtxTC3DP4qIKB2ZL7Z1
94PNHg1ZtHUOYa7EixgPo7jvnA/77oo286xeKaqymY5A1a3kXZgNgnT8MnoV/D5e
MM58MkIKG+1HoMV0dcRSi3I8cj0BhOwPit1CUue8Z7cB7ou45OKX5dk4vCP/1BjE
zX3Mszh6yfo1gWTtUjwiliF6EHO2ozSHWht+xEhrMq+9KrkKLhdc+NbUb7sXL1G8
jSaKKClnOB1HDT6G/udhbDpSqO5G/sZXxhZtZDAQvSbyga0S8Y6rlideaPpYLu38
p5jS5/z0IwS3IgOwJu1ywQWc8l3se17GADgd2XC1FR05bN2QpJ6MZX43mwCaxKpD
tf1GF10KwPGZ9i8cvWafv2Ub+qGK16HRfb2L6/FzT57tFKnxuGSuYKhLi3QzEA5T
2zaI4jtDMgsSsGSepEgbj1hJcXyHeNfpC04iimy5U6TXJly9nWIhhGXFWp9o3TWr
bTXu6F/flyx94yvnV1ybi6IWfHO17OyevNxiay/ZlWdPM19lOW47OKjkujJpUUd3
KFsv7vurdq1/Ku0k+dG3y/dflGEulhSr82kVg8Blo0pJvjIcjwl6dC3gTtBi0Q7L
cNBMhm+nl2oVH6bIy5Z5/3k4Ck1CCEOVJJQyDIh+X/3OH8q9i9ySfWIfbdoRrSML
ERnl+FTXAxVU3VsmYKzq+Kv9NWCZCKJlK+iTMwJZR83mq+re3zXmHwTqRW5RdV5L
rnPI8CZ0nTfw8dZTd2boO6r+X2sj41siHinY3Kw/jDCP+oaQx2GhF3L9cIhhj1+p
PWpH4xxYyKT72kjPVvrHTQbo2CVajWRZHQtwWklOFMOFKxNFT27X6lLv4OR4o9vP
+0+A1z7o6fO5bSk8AJa/HWxCqf1sGVIBD2vmJMs19BS/OongeHUMcaKrVSwg2xWq
1630fhisPgP5nWX77ahGmluObUQN95aNzriyP3mMo9hDoZ0BKWjR9uyalNEEdmBJ
k5nxRfBMmrog0HolyPyMCq6b7Cbjom8huJgbnadnEREtMeKX8dYiQLZZj3QNQwBf
qcrJFXeEHbm3mwRclrDNanI5HBfWD6qVTz2trKarAQeRK1gWbn/oT/5vYLnYO5HJ
nSBKw8Q/0R99phzdPry0OpMx/kNDRVxmy9EWpguE/lORzfvJd3dD3ItgGnaf0y2r
Pw/Wwseb5kQUsWxtth/iympQpoB0A5D8jQPdPkrv68Mjp2KknQa6WXWXVIbKJ26+
aF2tpuMjAu0cZPzPYEWsQFUg43ID4B73iOErllsQBItNpX94NOvZEdQXAIUWlc84
5Syuj0Bwus7CXoRkurTFleqBjyD5ucrFsdxhDIqRSuasYjauI5I4vKZhwo74ccmv
lQMiSn0EfpFf4weAB/XW9F/jonmPDMDX+d0BpsN6J/mYHWcTLA78VqaqbvJhh3dN
YjcddIKiuBBb1H8bxLbVe+d2AyN7vNJYgThHNm2wZlQNd2Z+NU4O60DO0PhXGI/9
EjQWVfCjtkHhzn1No9WflCXiqYFXGa3QAlU+Jvpkt6ypy10WGIiQrJIqlB96PpyS
2J5nmAvJwdV0d1peVm/1q5AWhWLnmXJm2kANMYyfnxTG2j7SWgULlME6EbKPdtx/
xOtSWsqYYtH9Qx7AqKz0oekKer738Ojavv/00DElirf8C7owtdOwExp6n9A1hJL6
sk5eEpSTOmBSmcNEYshePCiwy46Bm/UtrW5X3dtpKerUWlvJRu+1vR9O+esB/3z1
KL9IOUbo6Xd/9/8VJLt6tp26NibCtd6vz14Xr0JhiJ3D99CKeoLzK8+KgTylOvNG
TmKkF+KojZy59yNePmFNwaC+LVF+i9S79FO89P+d3GYP8goq5uSboQBC4/tsl81d
fcpYMt10x1rht8wXHpgxNbZKYkWlmCWfqtiIJZ97AFNjlhzvCEYAhd6u3l6xcX+/
smLMqBndZZYlqmTmirmyQGi8azL6cvxCLhITjUz/5BWwF3lc1sTz3FCeEv8kNjQI
WPnJUNvw9RIAX1MDRXxfBMRV+g/WZuiHDLYYHBrOze8SSavIOxzhth5j6li8jqLN
3keaN8e90dadWvb635wxMtL7v5Ihfhq7BMykRb2EJup1qVWzpS+lA3YIs7auJDsK
IFzc5OG9sNTLTZmr6D4AC9GVwSKRSX7kmd3ryuQoGalrnuc0+vuCtuo75CY6FTaC
RJPlA5lTvKOiNV6Kb4eY4ZAStcn8OBsXl+V5e+OrBxilijt3afSA6IOk8ItYLLPu
fdpkCDNrDIfyLPtVogRkUHPGMvcnveXB0ZsoaheClj6es8r+nzkLdlu3yqaKyLHf
RlKZFjuuA1QMV91d3NdYFQxQCUIo7GFh6VRPzKhZDVtQgD4KizfMZVSGuHzzMmCb
oB7iMMSMqO1+h7rONy6YcZJvVd/Kq/asu8xWjGZc/xA+AXLwzo35ASvTIArVuNPX
VMkx3kGvExpWNvPVloJ1rRfITKEJmiUUa0UDto21f3E7mYFbGExWRzRwoRgPstG1
a/X4IGwxspCFns83ZR27ka95EFbuy+2gqGPc4Xxa6+/Gh+iGzTMXThOAasBdlUXw
Iplt7HllBu3740fj+zz/8MzsXAWSswuMNnVonw5uUlvN/8r8rGfGVElZkDdYFyjR
S4qKSMqLZY6PYKWzO0wSxPpL7xCuj7Qw+r1nR+CSKdo5OFojgs92V8kbLhnbCwuP
TF82ERmT6JOLy/PMkok6ikmG94Y7ZTJ24SGAeNHROzh3UF1NFJ9YNxPdtOhGOcsE
JuE5haElYIviF4vot739yWcx3143axGHAleObm1e9dWVZUIJu469xOf5sEPqhOGD
o8cXyEwnY8FWzhF3F9rvYWwp3gt1nN2SBVZqFEozsHP8Xs5oUb4jcDIIT7tkNMYC
uzCjL4T1Iuwt2hvHX2BrBVJGiBEMn7FCyXkpuOF1OYq5D1lxpQmFG4y+0/OGvO1a
nUhWPhSIhSJutifUCyg6pZpuO8SHKFqtEWT7QEghUKbL0ATZxKW7vdAKSDFnlrJA
SgctBkpduOL96KPOy1dOWa73f203bz2O7j67BsMqvHHF2oktYdEZLtZ1xn1xSsd5
0SXqwyaN1A/m1jsaCyN3GAGHd8HxExjvxkcvwZBK8VbrSLSItls8XT2QlGOFXL9T
Lfsgtzg5/drmlZH7C1hMjihmNlXwjF2Pqk5WFhIQkJm1GiJa0ygLv7JmBsoGSn8i
mke2dTXilgK2lJz+kBdR9+VG8EBDNkso+pAorGRX/fJx2P3D/ak+lbDQUfDBJaR/
wmL9hx2Jwcr6Buq4FQgYKXUqOmXoDFl4x2qwzPFgZ0ZMbDI9JznZFfDy9GA0V8VW
7O8tlvrtCorLC6LzQniLIOBjmrQMMuEN0yZLH+jCqxLsQDefhqaCzBu1qidJ9qcu
A6UWTf/Q24MEdc0NRGcgVdMeD72FemsCvGbfscdW8QsRGuAgX2k9E2zYMtdG6Agv
bqfP92v9WtXAbUOMZCKGNWTr35iWWpEtSFQyMrBnJKj6NcypD74B1lbW20EA6bvL
E2qa9Emx1lBnJJJxgcsYB8rFUNgeTrMroo03tLrinELAdCzy5k9KPliRAIOh72F3
D+8RBjhUMy0GE+w9ncJoqe0ulw36z4ES2oaHyKijhK6zBj//mN8QHwORc+iU5Rs2
K7I82v0d5LAw0I9dpAj6BZZQQleirU3pmKAtvejRc1hpwypCWKRBB6diCvKju5vf
Bz5SRN8Hw+6zNh9AvaILgZvlyWuGfgtXIdVPGiTiiSXF7BlQmOQ4v1Wom9cBIe77
7NxQICrMZ+MGB79iNs49HYGumtP/h8YQsjQe9M2AGSJwbwt7LAwJHJIFKe23H0C5
pVHGy6830H/S8JtgzhO3rhNd3gOJmlcG/VYzXtE/PugwRx0tc8wKz/h/oeK9IqXY
IrciGzLPWmr0b184fqMZ42ueBoabMXE2RrACym+8xJ5/mzu3rFTY26RLLrkWQxle
vZdil+6+HiIgJmssKUw+5wNF+bMWUoUuM3eGQOuzcAYmr4aUJ0trzv6eVv6wzitz
TKb2v1sV+htBTuZYBC+XybBXC1hBfrP9MuMGqjZSivSN4gcQnQmcoJ7sXrtwUVl6
FHjzRBIH7h9hbUHwE6nPrsVtDyrLHdLuFgrS5J2iaDFCj5LP8cVrbIO/ga4KMKOd
dGC//belbI6WhRpcwVKeV/n3L2Uza2FX0US6K7y06qP8XxHOgdGXxnbedgDXHQs7
8MUP2Z84m9TvAtCFckQZcz8mzev57+CvwDIO70Zr7oOWmIzrdfZ788lXEqeqBGiN
c7yfzQh4odQtP+tClJ3u3/TapJCRri4/awAwhn4CvUTphCL6fEzqBdwmC65Eaaes
nF3R2HV62rj9ssKTJF6JSUsotafCBBG6/l67/kDmgAClGTrlRpEL25dHuToKjC+Y
ggeJsEa8aIQihjxkvnHcQT5+4G0oVMelwaZtg3Ker9Bc7Ayxx2/F/nbFMHPBNLdZ
D4ir3dg8jezqc7m7lMSyMkegGugoBODcedYH04lJ0LXkBrQczIHWNU38iJOdEJdv
lirnT36+7VqztNx8gLZgNXfrEsbD1Dfsvjk1ua8hGAuQW3s262urmcTjVaQAXPV5
PZgah1C9rhdgGQ6shGHNGzuA9xh0uUrEa0T7+cAHKuQSLCWmvbZDGMEWF1JPCK2u
QxVNJymyq+padhmAOp319Gr08f4UZhNvZscb1NJOfm4fJB0t/4UesaJPU+3s/zBn
e4G2T+OL01zuASFM9yEFb65coEQsuo099m/ADa2Dqn7M3jUDDEg+l1ZTlFvaveyQ
JpP4QGaWAwTtJ0QigA4EG9zg+UuyCq0Et2vZb9FUiz8sCrc1llSuZ7OTBcWZk16o
IM6zaNLByOUnzhVEQiyfJev4f5/MQEKrqpr8yliVoCV+39hlxwd/o+08wCMdQ7++
tDEI6mKPqcJq1rK0kDNOrf6K/UEb9JbnmC8A4wKlQ8oB0iQT/ijnIqTfMxLkvrhL
NR9fiPOr3I7DhUaXjOEoZocdz8NIwD6JFv91/ZJvxoAKOZGtIJWCcdD6D+m7/LBZ
vRYwTgJ845i6BtK+581M8F9DTrCYZl2W1dSRWdHs/f6mKSop/DABnF9Di643Gvwd
/FOqABcRGmW+BWsfIIdTatyDH0+Kc+KWBTOp4MW5X9c/hW+NYc7K+ECmvjWNx+A3
BNS5rR5xUhYT/z7M0SY5pk2PKSi5sELPePXJgry5xiWK5gVff9nYzhV9eQMa9LJQ
KL9m+SG0o86aH8DTyoYB2MrduMrBHyod2VT7Uw0Y6n6n7xW/3fMDoZm4kswe3uwm
s/lwDg8PqSHJbq0mwkcsNaOcfqgQ0j115pjVfumPB5EDgNhUTUt4bAO1BzGZfJGR
dJxuCweQroS1uWC1ZpfLja84GgFT2GxzsJxxjmOSfTUfwhppWhxui3Vkx3LWY+04
iuoXFzbQLjAnE94tuFykJMT/mb4ckys/yw+mwgk92TVqp7viL7EisrRcRX/31cUy
BTnMfFm5u/kDwNxu9mIx1f1L26MnZmySpe1lkgUP2eoNmO1DWQNbQVFdnknHWSfI
n3TCGsnyK1vL0eMkIq7ARb+V4pYng5LBeVfih16vPcku3tE5GEZFXdx+GxG9P83u
cZi+y8rIysEkPwjLTLDc0ae9Y9uZwbMN36MXzShbX8Ld74D5Wod2XTh4+M5VM8rP
g45r3XOHc6xuqcAgwsD8hFI3Wt2rGTLq3J+feQ9X5jFBP3brn9EYpYAHcJO9b7sy
xzeoHEa1aRz1ycMTt3CAoe7SoV2mzJPdv9j1uHFX2l8TPLOZVPyE3L/qIongr3dd
BhKDpw+gTbQyBzUcEYgc8sbEnjoE61/ZdqFhJyVuNKpmkzozq68qEUfiSK5wpc+J
ASvgKANw/ZXWRUAZ87eHD+pVA7XhKlqRnsl9riQuKeUm0W2rfITKNFYY57m87x2B
naEBsd6qVyRbpryLFDgyOX/GxrFgqGwnVRVbcQ7rINKLa7/IqZAoDHD3KHG3ZR2d
SddptH362bPHmKqNGKC7PCwfSyyLYaz1hRH+4/KqoZmyeCcRuWLjb8P0gYBw+aVk
RQq4pXNiPsDiNBim6pGpnOqdjbGL7/TzSoIiueIXEWMPuI3xO2TZDc8Dh1O0QuJZ
461rkyqvAAwQenlqqIirLAOjkl3xJEQPrXb5RG7qdKb4uHr5oxL8SNNrEtF0Jb6n
Hlmwl4Ug9RDN9zmo0wHpsV7BflRWY3koFGeI16eDptmqCb9m6Q3jA1kSub8WhPEX
c+LdeA6RugpfADdhK+CALXtDnL0XRFxqLgbbfoeE8RpLsKWFh5bkRcvOgchAcEaA
9g8yXqnMOaqAZfCecSaorg3TO6W1OnI6PQTuFUQpgyMfOcXWzxOqbX3HMyAXTnLx
PyGDhIoGWUf2TrNd24fBfFg8w6N59jLrCA/fcajdNSrSgUmGIj1sZ4xY5XGXuKbi
eiDkt8cVhIj6PxaLBI2EvG7TVjaDlqQG9oNurVIBb7ecQRH6cJIv9clxAxGS4/50
IKx4648o5h8fF9WGFNU4CkSG2FtpJJDzXiquMe0NFQg9aJJQaCORGh26hiE83I1u
/BApADhOwcwLN4IbE5UzoNsjZv6E1DYFOeGh4Y9n0TDvwyTYwv7nNzF+Ud0pfGBU
/yv6E067zZ8d9El2D2ZROj1AB+iBVvV3sK9wcIkFYYZ30h8K+9oj/poL6c9zT6YN
B945Pi54ABolIU7mDMHfblVK2hFgbtwEkhaVneJ4vBLvmD1f+OrNmtjGVuU2g+wa
Gae6JffO7fXrap1CmzyTFIb2Z8lTbF24jiBbWSNtTLhD9uKk1yDfzBun3PuF55t1
CXmHLeN4lhRMClEVRw4op8aHncMv586lXJBP8O4Q7PQR1QUwrdFGVl5fn4pOfHgb
Sb+6+9/GcjH6mrc/Fg9dMslMRqwblxYbxr3TxiP2M30fgratbazEDNCp+CJdwoP+
Vuxs8GPujrzRBusq6FB+rP6elfJ7VxiWp+5ozc4ChhVhmadVWradm8x+5xnWtuMT
bzmNi8eshu6ThfI13/ZXhjn8MP8LUO9hy1JaDHO5/DtP30H//Q+EfIGP2yhEapb7
UDUfKP0xh6+oz8Xqx6f9re8qbNvnIKDSz6zgwagiN0KnvkFmcjCeVtMz1kzf+8VN
YQ7JTPyhU3USFtqdNbZyekmmsPrtboB8BlZ309thD+H4u4/J0SQmJ6SlpwJG1mXM
CZ7x63dTNrUkNWL0ETAbTdpZodVX1N+pKFVgt3/+gX9+thPWcwX4H/abd4XIgAbK
nSu3B2VC+xe0/9f4+y8Qjp81N1ZCQB/3NQtQP577Rt7mvVBPVPpxdVA0IXrdJSo5
FE0F91J41LJXaXP2tYyPL8cwFFunlFbgK8Em4n3UqD76ORacOIjhrUp1Nx20nmrq
ndTYKAqiYu9gTRQy3USL2FLNEvO97rkZp0AbjpjzNeNyafwAncelVYFOfBJdy/lQ
TTbighg+2rPouusnRXVFWYM2sZ+zyDSZF2Rqejhn3ZFH9G5IMmJBnZuAQmZa+I4U
3s1E9uHsPBtzAAcOOv5znwM9kWuUz0QXjxzBfab8yLtMZWf9XhkVJOWseU5Va5yF
j1Eom1RSDjloWksPFVf76LCQ9TWG7tLM8/Zm69E4YivRQXgy2ixhI44ohiBnFy+i
tPLr5FpdTBZ6+NaI67PQ3bYtEvLOb9Yp0HGPdaA9WzH9jJTrqbf1RmMnO8TeBV84
pETJHocPDL/gmDWgIf188AfPhTKfJHUMCri0RsJFXIuw9DoPckP0ex0LCJqO7IvZ
W8BpGjG4WKdbSmLzam7mz6JYM+LVIasTsBGMry62wmWAWhHDH7GdFgzqAJ9jtxmV
GoG3+GmuUMh9O8QbbnZNuQ4113gojiK6MNGvCOJT1l1O30a6h1fxYZ20QslqtKej
tPNm2nvBOg5zXu754V4m0NGlCP5c6b0PnxM5beI1SWB+Uj44ptZF1KSLCYLeTufZ
Zk6a5bLeK1qiCR1PAuaMhrCtpEIEPMsFnXJT4v3Uxe5MC7Y/iQ2ueTvwaEr9Kv0y
hWdxDbu7o4l/UylS1eWKHANWIWB/OTlVyw59fk+XnqNPO29GfyMZ279M+B3Dnz8O
w8XhnOIoHqjgS9RjlJf+FDUyEM8SSeeGhdr8N3N64rszUcA5FgFRu6WN+pgLSfB4
zwzU6sOa0dFUkqurXMqqOzc4XnjSB+SMy/6uPUSoXbpt3JfLuxi/teUsfIPhK9x6
oav7rLTkvUd3dhzJaPteo+42huzE2iwtMYuEY/7k45Pj4RRjs2pUpkmSYOaBmUX9
DiWZjNSd2eF+6CnoekG9RtszQ/SjbOKm4hedb1G9lRn5le5YnoKOLZs28R+6rH/L
uR+AfYsaR9Xc3bUpRWBTQdcve1xC3yU2qcv2DqCI9srCWnbeKmQP/d4axrbFCB3P
bVbkc4rwgCOZU57RpBxVRYlO+9GfzFR9x+wJFCs4xJhV67BbZmJQw8JLPIvNG+20
hKCB337sXvM2f5N8bkvl1ef6Qh7N7+aKsqa/sdGpvs6NQc9oKbT7ORGExtWnrzO+
WvfACps4UAA4glwYgcWCptgjEXtvoYALnyAdtePblllWyWumJ3KT+QhRfjCb0+zo
F5FgdpPlJT8uZg6UIgX/4m9Dot2o8rnxpL+TP7s7vcoc1VjmgxqXcktv6vVCq9BT
OSFeloADCw50eTPASJz9/hRl50NN+0nFlzuCfJrOPqXWQD9G2Iwatk7ZTt3UJUT0
cbByzSTVoY23DWZ8K6QfuGOkfBbPVatm/JMJvuUVveTT2Y9sh9A3qNnXHVT0TLmG
mVIcU0fA3voYJ49pEOQTmGX6hqdk2/db73xqe2E175YCCDWlD6t4GRaJ10ufKELp
KRsAkFohsWKxJQ77apb1cu3lca8Bvo5wF0F2weVx30pMBztE50PP2Bv+V24h/H3Y
NFzFf2m/8DMYRjiFjAH1Srvs+0GZoq9PGumjl830Bk5g/WDUe1gosBWZSXyBeEZ9
PrLVOgqX1VK/llHV//NFMNSxsNkgKjY0iHFVeZkUhh4uOqhi0NKHNhMQ44xBRhQM
+Wzun7HPvNhMV3z4jARVnHyLe3tAwuJj8uGtxDzC8FB/v9IzgfYEqd+wu7/KAEVh
25qjrL+uor6heCnP2lgv4ZRhPbHvoXXf1c+eWiawSiLDQX2IZ6aLfUoB+/mb263U
/pXpN2j5id2/DOu7kf+tC0oAqTrUfJ9eeE2hdQ4dZwY8GWdnxT+5w+2fpiAcIbf2
4JLx8V8Hol59DzodbkHwZ/8dstr1xPPO8jR66AXTGj4y8NMXCAlk6Y7X2kfyU2l/
0+x3Z6HaJZKSnHEs3b7BxWYfeW20WHEy/JUXffiqoSxYUTwhsWX5ktTipMXeAiOf
NookJanv8demtzshwm9qI0MQxnfBtgkCvT/Vkd59DFSNqfW9f1num8GL6A/7dx1A
7koM54FBzXI7so+JeeKWYego3f/nsQvTpUYoUAAoWrHB4ZOu7jpKGFmqN/iLp8Pl
xwEL3Nu8cpgDJvGqiiCoG98bY//B5ud0gyJqzQIgnIwAC3lH5xkMO5yrxw5qCnUJ
ZgIQvgx6B4imqVplBFXZMv3OGmY8wAm8dHbH8CtlAq3oTxWudTdbOQvEnHT+FuEX
zW26RmsMm7+JDGoh6fUQ1qvb0J3nuEHwxErCsDlUHdhBPgCm6e9sdFQP3obLLdpM
TFa6DO5osWPet0qPFa6/lW+uAFx4Cffld+tnCGl4YvYoHJpkQyG4CH55SLkvpYLK
0JEdFNNdWNINORWU09+JOconBV6OSL1ozOy/SJxYdCbYq1F90tT0z6jWOHGXTzOf
Ecb5PPCvwXuKMAO87RtB/wRYo+3umuDeshR2/OviUirTj23nENuvllN0WyH5gO+n
aoww2oJuGk6AMV2qLuZSqut476Fc8c6IfsnYRG/0/y5vT4ZIduHgdHy9rnkpDMHN
mSPxyouuhT1thjeLnFZ4Sqt5i3cjs63/f75nf0Es9uc/VmM+tCiVoUTonZzqR5Aa
5j3Wm0lGRFTG00XqcMRyeQvncpMQ8maBKcOXbBnEQlQhZ0alxP1oCimt31iTCCv4
Vh9BuiW6JJ7vPrYVmn0/bx8BzC3BHeAHrDWYk37ajb5E/nGv/iBd/MhXuy9q8iZP
LJqdOGxjFOw/T2HIhu3LPUHdgSmvh7O6Jtd6J9lhO4Lldq9ncz6E7GxyJTlNDqgI
moKQExPTDBmfifkP9S13r+PjyEwZdJs3Em+kZCiAp1ZdxTnVWZpoEBeQ9h5z6PIo
mq6ySumgacl+s6TsR6pvUw274ScMul6xzMaeGBaI7YwP7VZ5W1t7NQPkIMat0+bG
o31xJZjrv4o49Agv0T2KkZ/xuuYW6WXAKPoaIQf+3xMFZSuAeD73se44FINAAltk
cB08EaK58jfC+pr0KLi9y+zYVEIb+enQhecPue6fcuZZvkSQtXtBpkHEfv5yPVPF
cBuIEHswaVnXsp8MKF9waYTGQT8th8gaTsdFVJwt7tN5KE1VM5A5oIup+frF5eTk
LB+kVJLZFfkDrcB0zJihxrxTz0pKb4fAiVE+VpxjNovTLJaUspMjf2Jdcwo5Gn/x
k7laTw6H2ABiwGsIq8aWCEwGCe9zXjxVpqpcVWWgQe6g5s7Wo2bBqqRowA3W2H21
I2Mk6JHLSCrzD9nuTekRHYEVu6sFGCqWmuEzQffxOujOK+dQKxnmS4iOPN9AZAvk
59QkM4GOaeldkSGmf2Z9ykTmpWU8Yofni0JmCljH0fJHe2Bif1kTZwDLTF9/7MCC
m7RGG8UZ2lsMFpn/IZrgckocWUWYx/D46ktDPSpDAQ29QLCLijIN9SWEsgPjy68v
iDM53PU5mgLSbBRy3Un6WRklzVOIJc+pxvtmf04nXXrkHSy/2+x5yu5UEZw+a/vW
7ZU8u6Ydiq2lZHNTT8TPVrtqhOxS8DRuH17aRjk3H+AgLp5qB09Ikg6pCpU9fXtm
Y+W+PDke5aR8XPu7eI01x124vPMKFV52jKwL2/yh2BzHhG9c9n98Py5TWQ9Mus9b
SCjGWRC32Lx5CwD8zR+w7SXo88Hprff6tnKYD1nmSlEFEq5hyQBL/f13GjbbcMk4
gKxgMj/2eaI/tz1FSaU3dnxX+rYItI7R6ymPLXgFOdfMWl7++7fRKxig3f7qXsZ0
ehNkfiFsBVdksFFX54gn5Peus+4GTygir96Z2vm/EjPMt8wh/IH8ND99JyhnZOht
gcRwadCFXxPo9iNHZ5bi9OzSOp/TxCd8rxBai73yyQvm3eK7O1fS1snN0QfaqpB6
vZvjMQxiV/UtVT7pzwh/A8URxhopPAGZztulwAn3Fha6w6I2SLHYzy367OTdtQvc
uksXdCJvsXG/jMB2VpoiRsdpBu4VUedrxVK938Om61m+mBayU93bLUCOTj0nsneL
eHH6MffJ577OZfV5Nf2LbFkfHJIMVz5txPIdqnBzjsQF4qMgyeItwx602Dua2Sr5
6E1kt3CUv2BmVhVkhBHUngtaI90SfsjF9Rr+GP2pAYeY93UNAzZMmn7a6z+1QSio
MXdclrLrNMUSCjqAwXxXaY3ODJIKrgdopIrMjpHlLQA536N9uRElEQnxZNwJLdG7
DRNEXannmtIIWmMeHbI7lpGGArGEORvcpTusTzcvy/jJJ3AgSxGnKlYS/5Bo8WTa
mQfp5KV//cKfqcicUcP/9sWozdVO3u5/XYMpJUitIFN4Fe8gQ9WcXs2C4GMQbeWK
oYNYNVZgJFQ/5Y/5eTfOwfEfoVbA/5RIOS7WQcsG0/HnxfxT2bRQsw1msjv7nXMl
KQOGBqeDX3YzBMVuY724BFw9FkPA+2QgJuHar89Z9PvpIgey7tymvvpBKU9SlvIY
3FdrqyjebqFb7os4qBGc7HVJEceP4UKxkbd42U3tX43ILFym4xlMy/P4wKtS8O+V
S49JBetk9CCD0DGet/0aHRbscPy8Itu3oqAXrA6SS3kpMPeKGYBKtjroTnmURObr
qAiK6f9YCZ+RvHFWRAEFvYQA6AynkShXRf1wS+YVjWnYg9vfHPPHENpAm0QWtade
2Mq+Srp0YStSj4qjxYVjP07Fi2j4X/4OYp7lRzG77cxNm5crnpFJv5NZ2fGTgC0j
hFeWpYAvLLzGzSHbaWc50KnB7TTip5meRjLQrSO9MoABuW9Ax5rm88hWqAmP0OqF
Wew165f7avZkNpL1AfIVzGLSWEKCEye3gU2/0xCsmTy59MM8EjNY95PSk3KId/P2
mZrAdxTMME8oRDQhnYS+Nl8o5ANvojm96R8zXN6E8MjlYLHixpN3Pl97zFKisQe1
glZjN0LfE5Tjbwv4gHn3NMUxLhW0NHda9UXnO/ahSR0xI/0cKNO/g54tPc7qL9sY
vvAON+9gohTBURaahThPayKENp//orvKBjFbykPxApvzaiKO0C/orXMZ5qkClG5Z
V9eN0P+Vjc7wZU6czI67aJqDfEyV4ei+13H3hVVq7qGc6qGDw3NEcayLQbOFK91N
kdb3Qp1uhL6WZY1HvTlb6Ta8upW0O5aW5cbrtff9mirLJ6A87UDMSKX+L3v62sBc
R5TSHeUAqfkUo80uo4qPlYg1GiTS2YEC7GGw5zRtvgcvzv4NHRR/bPk7M/b4ldCl
HBNIojELCNBM5sfA44eF6zYMeMSNWGNE+5u95LvzCXd3lFPz20CxUSyCW38hvpG7
v2WiHdekRHkpWcORQrRZGNImDPhPQwJahJ4I8d4bX+wScD/BZb3gURKAjaU4GsZo
ADPX7Xeb1gEuu/pXq/d2qrf5bKoiuoX19R78amHzUW4ssLpYp+1tcp/RPqa/OfII
1i6OaVyc38S71kskpLPNGUjEb9EXX6mERDlOveQBEJ81TVfYs9pJf0gqUPpz46f5
PCWgho7Hqs2cVlAq7vmgEUMZa8KOccfYQhh8UAluo5adYORYMMpdyQ6CJtyTLqRP
kQw1UohbwuIzCj1WbZ7ZA7DsNHjQ75IrhKnUy5cemz3tJ7v0oAJN3pUOVzPs1eha
1VLq+eXSBSSwAf0zILD7gxyJiUPSLPtyDRJ/3gFm0ksSNHHxnqNn4PP4u8aPnnNO
SVbbLFjw1srwPWwByBGn1gTGrCVP/BWwdIpj+RHEDRU3hBqTNeSUvfnDYXK1nr32
8qkjHRHwXiK0P1ug2RrelBiSDqq2Aqwc7KExJBtDOslTB1JHElO0A2Indq9MBR+n
j8wBx71hhkIknEKE1Tjc7rF3gXr85RHI+lnyQl2ckxhO8BATSdaGpKPJc0S41h0P
lo1r+4gOejGdstEkqYN6K0KFREy1cWYkyZuumNwTVygc7Lswuud69NRHXgg9gF1X
4vhSbwcgcKqOVx1UXjaVcTflNZSrhEOO4fiq/LTpN7MfzOoSuQKrP+mB4k6cK0YA
T8eyNDEES02FBlkJ264mZSsXMZIWOqkaGwT8/ivPgOw/R36cJ+DjYveO9QkYy6gv
/6UGUCNVDqvW0gzAponTzWHzi9NpXuyhPOR499SG6DKjkK8Ga7l+2p5u69uMIZqx
z2Q/bCw9RbBfjHhqwrNnCQPzDuJWCtB9rQOzSzk+L2vtfWLjYJ7xn3ylssGxPxER
ptVcdB0vHR1kyTyaxlNhZJUWin+RyuBn0YfOP2YGI0NTd0kiv7aItCj9yL/GBFfK
4QUS2IsHOss7dRg+Fe1oIaT+NsoFsHKnGh6L8xVgp/lwXhsw5H/t5j2V9M7ixq3D
cvrcfjoFRk9M2caFFbg1EdZryFRwtTTg2qJoJ6NI7o74ttD9qsqN57lUeNzkO718
gTFsTLSAgbCWpdwMlQNrqnPwrFxgO58wDO+rftUe6pPTVGppdxQ6WwOgClEZyAvo
QZRYHOAbQgDIgYAsrAO6EARzqXXfmyEpdMQy7/wg73WSUeWH2J7qehFf7u2E8/RY
+MX6X3WGLluho2HfiFEbjmqyQhwcQYaPpl7dKw0tYCvs2oqSvSHbFKaiCPmVEszI
OdxtV7sv8RHB2Om4l35YyNNH/c/C2fU8a50+BcnZ2LBe7ZE/+Sg8LQ8dyKZGDQAU
99GehFv6Y3UQ6PAOjgGaciw8xaOjqJXQcb9cd1Tq5lV/j5DWZsyT8zr3mReIa9ZJ
oP+0ZfxPBAnmDIzFA5fEy9A2+q9TOWcVg8Dko5ux0LX+yVu/8KVHXz5MBwvk4UNk
Kr1NLgQ/zuaTleBZE+gFLRnnHT6GfnveqiHcyrO5zGzor1DPEr+HDUgLEC1P8YKg
jqZLStrP3aEIKeen8Sgouso36UNn9+RIe19IEH2azOc06rBnO5Epp1/Kk/TCkC41
VWOR2q9c0swQwR5sCOGL8nLZHAgNg6J4H0YnP3Vi1n3EkaabkUJUakTwWKdSRjSS
MECe1baGZtbsyTUoyb3KziPElNHM8wfjuRw+p+rtH49bJSONyjks0VhETF4vb6rM
O6PfmZruccW+HAkOh/F+GwRXys35uPtNde6b/eOj3U1fkoZ0Dc+OgWqDVXbnq3EL
cBsatTSqL+pnvw+91xxcJw6dOfoHFRwIy07Q0fqnydcyMTvuywZ8Vc/f9EVGOdm+
w08Yp3MKo/B8GgeZ+5fspMORS9YMfpnuJ4WErZ+JwEjq71qG4B+TXyEthLrla6Wk
mfD003hHv/x8b9Hz96Y6HtF5EST0pGvisx9PmQhSFPuXyGcFkzsFhJuRCkBgwaU+
EYl+9fPZBlk4SpvyDXuDHnJvJEowpYM7lE8KqPKaLZ8qu7j5YVvD5iFy1pUaMMt+
NA+8lUSUg5gp1n4aI49f/hSJ0W9YN/AVRWRCMV89F5d5lOt6Vi4vzEhyuFbzb9Me
oR0VYCZ7DOJeicQD3WQaiVA49b0tAMO22sCw8fC+MTR7d/JN3iSY0xKohlg9wlvk
JxTzKClVmCXEmT1gaW8S12syQHkP0XWGOMEbFh/YUkyFN9Yrd9Xnon1IpKydBWWX
o62gN1JmfFmAyfj29zFQ2iDMe1yxLc3PT/ug914I+JWNj5qoqBnCugRID+6428Qz
RwV2dUJeIwGoojnyncDZNwzCNlrWhf0RwUvdCbyKrlzwN5Uf9h22QJVMSwRn5rQD
STHW+7DNjnzWIQTqTHRJzZ16KPtPRzTv9zpSbfgR+7Sqq21OPfGjQ4TxQoYqYRG8
NU/jtqAT2Xw4vTZA91WSggLzcuygacM+hOIXQN9v/jRktfCnEc4+TuIvPzGmTrw0
grRKNr1mbOUVv/NGoKxOqAh7ojMqV2hCToXUv2B9SU96a796uBdHm0mXql9Z4uQ6
jqhgz0l4Zr7tLQRdP1vNOuYKUgjzwrEbe4cW+6lFERhpEMgonST/PSDymy//N1YI
PA0rk6BbVO5H8QVMOZBqS7AcQ6n+BBd/Z0VWsJCLseatJDi+SY3sW+pOTvsKjn/o
QCJHISqhv0St8NO0VPHtjbCVLbzmgfIMpZglKN56cmvQ9GnS0LdbIajlp82u0/yD
DrgoM5eBPVYwR7w+ZvrmH1mGJBfoYHjdg8m470FIAoeoeuh/txRgDSkx0qEh1gFf
XxS/snHe9Vk74k4KWrcIkyOHD2H8OyIdYHINutpZTUvHNlDeZgc3aiIGfV7cLv7o
+En4ysCkeovMjq5h/sYFhnURg1zXjQXkwV/9JyGPeRjGBeYMPu8s0fA/UNaImjID
5rGJrEHklyribfeRu9mkmE+IVtA02gXgAvs7P+RW5uJr2RKi69ui9B6qh0GfgdN0
kd+ZZcKI6UvZwzsaevKwV3iuNqgqvpZseeyurK1IkdYydKDQJByaaYBmJRdQHAC6
GxV/xvpaMA0vVggyZeMx6cuzNYRzfjkgORIlwgUjENIqLYbV6EfLwkBTc3zJluNC
f5KnT7/C1CLK585TTl3rA4v5pV25CQhi4NFzIfQvzickExMKOPyEjYGIgQgIAF7o
4oCcy1KFeMCM1+LZ9ROQfFMfkCS/AY/PvQHVj2Y3bW5dHJEEbRwZk524YUJ6P5ev
4zrthrCXbzbS6oi4lqrhpqZfVHS19VRezNUTYgRBMrO923+6HsqWGd5b8Foq4RIw
UWgyqqaRq8nwtjDE4F2HCsIa/TxtKGZa4X7wUtohbYnUvPviViaAtzCZxXlmc9Ln
0p2K04LTDsiPxYU4fDIQ5zXAixE+5dbP2JWGv6rcullYkQB3kBiZ10pKiO7OUGu7
IRif1UAHUd5aaWhhPCy3t2+HDcWfSis6KSvUewSX8D61YezPRFqAG5gf0emuszZl
LzSczhJMDxelK6hKbE480PAvnBmiwRqw2XSusLIjKgH62OsFlJgKtQ8GherYUW2Z
gywpokOOyK8ZEWWsKRw7Fszot4hZHsZyDoT26poYcmVehXsh8lxs30/4RHn9UAOZ
GWquQ0q8mVy1rnDZmx8LOj1mJeQm8Xmp58Ygr5XxNCAtqoXbLXv9atDiKdBfDVIZ
5bJHNBV64J1V/Ck+K+ao2JRinU2C6wM35yDX9HFoKiRspLD9Kwzl2tfMhgLpbfPo
p8HxKe0rdAxOdik4LyekTmvOw6sNrmD5skwqWW315WRb70HsIrX/R/aK2oyBizPF
fHbyt3BcPhyMW1n3geYTKXwbgjHRFcQrXROdTHvLSpA/G+SYgHL/s2VheD/dg7hP
q+DYJ/AetflZD+DwO2KEwXK8nR6IiOLsYft8F/18ilvKACULKtSPPqYW7UDVMH+t
gwdDsWd95pKsrfcLgGhUBi3k/2k+uuF0F3q5xdTZBebUzXjjCYG8NXnXoJLxSwiY
l/bsBqF9Ol+SAM8Pjp4+4l8A9JHR7SRPpnan8zSCGrYEFJKKe9OfsTLLQAWWT+96
v5hAmDWcY8bVKjxnAWDBCcg0kE9GqIEHjn0gJhZUrJaUdo9Wr4fMKEHkm0n24qWB
+3IkVTIyFePCVAkNE8YwihkciBQQykpno6/pJrqHVo6b2A/0pwgAVP/o0GDbLxqL
9w1FSgqcz9BHSnW3seUhRMJLW6hnJtlmHYHPLLzkrrewoIiQKx6i0wc+4MziDe00
U6n3PPJYauZvXK5YQJbIgQWAYvMFuu9J+7IkCZ/C+N3mj5ijCd8tAbJiWMHetnp8
6NmNpQya7+7efaJtTCJ2yYZdTo0Aid816EeGXqn+5UH5M4QFsLmaczb1J4gjq9BT
EP+1ifBgufwwrec4FnCzXKYeKZUBQoI92HKhDaCPE5pjanacawG3CppB/fJFFSz3
6ET9pXmkPn1Wtf9p0TVdTOf9XMv4JtNOqG6fzZxZibWMHLRP7AAeWVx6DwVXsjnO
cSoEOiY8blgqe3QSLEcEzwQ5pSgOSh/oKODD5JEtnUaY9G0+UTrvoeQgkFFLoUO7
OyhTx+qV8/hUmkVtmhefzskOcWkhXhvYNYuppQH699RC7jesk6l2LYSCqskfOarN
zKvT//DVYbuwp0n3SGm7lng7EKhnBQ9JprkulwAKNG4xZjlqBGeaTU2sEVH2hak9
jof+Wpio4N3zX+an070H1UOsDsgqC6f2UvhXP/81zyzshgUAxqjMgN1EDcFUuOiX
N6anGgWw+AmXO7kxb0mqoNrIic7uTXGBE3X0OXRS3dT6koFRY5wPyCHnRT1acsjU
dUUvZ+YjuJ+SQNe3+A/dQaEDZnhFfJsq6j5dn7nSF5bDJKE4DWC0sUJQtSfzQ8CK
E9Kin2Mgb62oR2B/MVUX1VwG4A43eiGz/Em+wRskIsGyd6/lPvhMTZTFAcCDTjeG
uwQnhIi0R0coO8a2Wd+uU1qN8UF3VI5QANl3iNWOOQAxRyMui1sbGRBnEJMRhteU
iflAifZa/nw81b5Ov5eORcOJTJA88tw+6WoMoaPtS+Rr+aOpVZnVVwjZSABrH6qJ
uQAZ/+wRBr7RYA1YV/HzWGsE0wCEjkvM5Z55eI4swIzjwJuxkAxuap6iiSDKrcWT
6QMXFVuMNNCFuTDo1Gia+yEm5cBNjIRHKCuUfWuMxkKTPFFd2M1w9wpgqfTvbI+D
sH/5Y7GN679Jy9ToxuSDf1R1Mgy+ZIF6moSlgu+T4PfXXjfRXpE/NfFLtT+VG6Of
kzp7WKdreh7mFsaMR9rLqMn9pjoVFgK70IATYj1kgh0v1qR79mYzhcWH/CV9dHVD
sQYtXZ8ovL4Bdm9zJJWoUECNBpFXGZ7sY5xxoU4wMP3FYTjq9XahBUPyCgSZZgrc
46ClYijpNMaxDRxv9oUWU+ysuIl9c73erdsaPwpbHh9luk6wFNYlhswbat2kcXkQ
31vXuWbTTOH6q9ut0S8eMu2uPXSutN3kyuj/xmNd2ilTRSuXxz91Z8SZvRni7PWO
qu12HKqsdj9mLYJLW5x03Sr+p8VxdazJDeZz4G8Ijxl0cNC0wsRQwD4W4MSkQByO
VuTr2FnVMdieinF256b3SuswS8b1bkUtu2DJa+lO50fkh2kEGwPhXxAbO+t228/2
mEfUMpty4LL57QRSHDbmgyO+6CeYV1lJGA9SeSZUyYD8zJnEXH3JTrq4/hB2Cbfr
QHdv8nJmJjjdXlMGo6PS5RFU/Z18nNtAAu7Cu/JLySPvNdSrv4xmP4K6U0QoVmMd
WO466OnIAC3ZGeDNlCQlQIGYqgqscUzPhTYYCY+bzPB4G01EPep6KBFcrxmsdbKS
JnS40kqhZJDFapBSXXq+I5ZTgh+Pc128UPnPTLuF2q0slGoMCXD7OHuZK5rpVGYf
nMY8bX4fn4nzDgdQ8GQePCBXsfpB4EiFKV6xaQ7XZ1hNvwt+o35RArynhgtgfhz3
Q12oAa5sx/rs7q8WvAp37ei5jPVGUTgrbhbovcLHTha2q8EeRiUhFzGPqf0duWdN
UB6EYk192U00WUOMQvNUIaLI0bKvmr3+/y3MnmQPH2plfjxp9VTf/IfBBrK/E3ZG
q9m8D+t14Dyw0lD9Mpbjf2bJzeNHjAP6bLS+rN6wibb7JzC0fux5720uEC3YkdK6
+mM6MyhdqQwkMDe22e/nbcldZrwjgGjKmy6wNJFhclrfiS+Qxv3kKqj8O7aPSWwW
xS3Tk4tFFdaUp0BieAG7F53C6N1Ow0ndgL2vmuGmaMbc62Q6KIKLpodSLgteuGD4
5vopSbzJ1zeZn83QKhSWn/kT3g17zF7O8ihTvoEBbtAdiVftJQtk1Mjmoejid5Q/
hoFIOGqG+nS51odaiaFCXwj4dJgIRaADF8voXFcGCIDgMm3ZRLcTQzCSQEfruNns
xMWPHsyARt04EPioiwPVNSat+kVNXXfaBhIN1PqpNYCPT6CqIyncHwptIfT4MN7n
WRY1xDmzUSmQsjC+DLxlEeGygc4mqsnLItNCp3wk7lA2LVeRu/FJw+oQF48keC6j
YTJuIoEq7xy01YQAOZwhsAq81pFmM4duA8OcE4wPZjlgIEphYtFDtK/jP55pLqy4
99+/rVIayV0AwVpB/ovvXIZ37Rmuoo7AqpkD3c9XfEEodmvESUlkTDogyziy9Ngi
4Do/AKOT9lwOu1Lkpji659lGjV1Aw03HeVOfL8AOrLMXfCVAZYaWGPiM0L6i9h63
f8sPV9T/3ZaEAJz/i5A2ClY0d2LAjiHs4nUAcWp9Uia2G2MvFhfZCPk1/fAtMsVV
W0quaSB0JnhDXOuvISvYq6KOG6Bg3FwrzDN6hm6EV+fjd+ptIz/6GMp3bgPMvE5m
HcqduzNdmNkJKS4F6JeRMjppuR/FY6LGPXID13CwBxu7dcFgcKzJ4CIUu2ZFpqgt
uYN7iWJqwXI4+c9iXnvDJKEd/5fIBcvvrJpDT27MNiRskJHbk5qXiF4trcmW82c6
+jYYdJfQOMsd94duXpg5cSENDnmtH2/PcLe9qlJQux2KB3VSVu2APtDSqCGrd3t0
Kk/8rSSQgKelmuYTJp4LgIqGaRPX24RkY+VXAXXPs52zB7prCSpYecp39GIuNVvr
2zudIVOBl49ln/1T4+iogUU1Cg0bpKe6ijaSUx4cqVccl4GoBEBBhwAG4wQEbQ11
mBR4PfA5nVBa1ORqSfBKUl/N+fADqSEYiZoBHlOiVhPa2xM2Y314yTkVKX/S/d1r
oSUvKAwealp1sJulfNCwEpGrpTD/HggT6vTuXGvX7x2Brd6sUBqqZxkgvH06Ocd3
XEEQ8bthvMf4kRPGZhq1XZPWwELbLiU3lEqspfsmeTCS0o4JFInFoLpSTq9u9PFG
HB4GGQfXujpWey71wDcIlFQhubJKGWIHXiRYr6q1kUjuRsykao7u6FRQOaBPCWE1
h6qiISnncD4mOvJqSv2zveUMVzFqn94sD5qgS+XQlJIyUDf9tR9XbIyCWebgOEQr
mI3/bGvYHxvYbe3NP5RJivS4t6reGJbQK4iOTRJKO7Kq9rYwM6cILAIjHHeqKcW4
evs7lgONIausRF4tX/lW2CAlEheqRowRJkodf7o5c2DWoASCjjIUMFv1mdzJf5UO
oox0HrPUGCDHzo+NczxW0fZ1VCWjDEJ99qzNUyrZSfD6dZIM3iEHlV5HyVtTh4+p
nFPCmAkS4416a8971mkrBrMx7iycVFSLfeL/hf9toqHMbNUVmhor5yVefCT5XhSk
qjkjKUNFcLmh1i/UmXue7srmozztEvLgAdCctYQJElo9uYUf5IXs8DdwwtUiitLG
Xh63taLL9aJMSZhwfZTI9JhZ2cThZcR/rmvvlkJaXTYF41qJEAdYMn23x1TWdOO3
JjUyoVldlV4TDmC+CFuzPV/IXa6YD8k+4j7GHmcF52QHcoCuyYsXQwK0O0BwMvl0
UmHqYAOnJDratHEtuWN4bGsQU06OC7wYAxYEPjUIm8jE+P9p8KTifDv6H+DS+1Ob
elOOxbNbZjkupoylezs4HwO6IKCIFTxh5HPo7gsi03rFpa53vCwMUZsUCPnxnCIR
Jnuey1Ur+tbhJRkXbIr5lIf6J/nRO8kMVmWYCzKl5o9WhHB/Qzw8qciRmfI+BJst
EuKomUpxOeZuvsvHamycTlPSldVYUqZMV4p6L3a/ShJXjL6HgZygGHj/fo9IfwAT
HaaHu4ykU5IZyhaq2XBlJSk3FFXeEAwROAj+zAxJ16VAORJ3KeOQVxwf2TMciT+A
ShpB5iSNRF1XABMdfACilD+VqvRt51UEW6iaYiyoIzajrLLpJMVj3skizLqkae94
qYEKDATRzJnURrQS1uH3c9919KVH8j4rQp86pkgI1XbmDeuJUsuCzoJ2EfHdNsTD
Vn0TXrSZjwLaq2ApOtqOiLEMgAZwPWDQ33Xbth8yvTo1DO8DF+EhShX0OwYwScTe
3BHOhtC9nYkXc8jsELMfuBR22/09mLZ++LCwZVu7PqXueLpSGyYl85B/rwgPICgh
5tnpbSkoZV++ne1Ah3RL5+r8RlAeYDLRwVEznX/uTpWV7TF8/IdSrKoeuDj4o5so
bhZjg2ZkaOjqDqRmqtz3E3JmxZprc2hdYxOw0R7Fl9e8V+GQ+PuRkBxF49vUbrQ9
hL6a6P7seoPrMH3K7uZTamlfwmDUljxiSVNNGURVEtasFJay+pI5ZcCDx7W31kTR
Uwuq0pfXV36JNsDhhdVosmMvk5tdy8vvqCjHY5ShHL2R42azn80kLijcj5a9f2WO
24W64DHwIpusZX4PleOIfRHQiN6YVm8UiEW5nZMEWIa25ig1u2wy8SnqaiuHxFas
z8e0Iq4FjWvKJg/4/foNmbEaAa4xsUVoxU1rx2D4VgOKxHbSFEP/Uz2+eLcChAUP
X1Zz9F5j6r9UFVn8ERJbYdmaggGwzefrSNyZmIlX41tgHKen9RjxNQU1/PzSqEtj
FKveXKyy5LjkLGQIFE3JRN9TFmtn/HhKglknf90Xbqrmcc2x41GuciGj5ahz08VS
IwFUU//qXlX7JdoKVBf+bfNQBibEys2SNvPYsy+mdgLizC62XV0q3tfei6sSs9dY
PZ0rv88dYgtrjILQaGBMSOj9k6wYjtXfac1TcoONOc0RTno3I37lh/bSGK9QAq15
JR+OzEWxTr/JfJiX1hl0WAjOXlAr6H/js4SA/qu3NBT7E+zatgyvuFPzIt31n9EX
e3MbxhS42Y0dEBfNhceuuwmhNDlcek4VaFQeRxtXg1HYEqLupLaG5u1g3zv3KZIZ
wJTK4io2FbxdEXP21ndJSA9INRAG4JqOy1OAj09KNdWu8fEeGcSMYmWaXrgzmr1k
fubvUbCTzUJ3TZG0Uhm1MHz0GaIeQ7s9oaVZGtdvYNIwgxZEAVlZf6YuYUnG+7M2
QuG7AEp9O8vzKFpC3g7GMxrsNmk6GP36FJjVwG7xVseYEkUSzXSxrk5X7qrGhBub
7ARfXf1eh3L+5ZwPxmvxpSh11UEWxHE2r7T9T6TZDdMlI7cwqVGa0qw1kSsMdiFW
9Ha/bRP5mZ2GNc6G97S4AMPo/DjgzKu3mmRk2JKHoEL/gCuzd6tzbxBy1YZy7puL
cWvZFLHaTtG/+yYVrv4gjBtoEYu44SrQhdzlngun/RRy/5zDDdMykUF3029jbVUc
pad1Q2GUdQXMSE1dTDaww1oH8EOG3xneWRCul6t4miU1ZFtFZ/CmrQPA7aamh4/4
xxFqRjDGcWuvPsJVPIyBVSRk/DHBSJ6FkOP/oTw2z1nTwqxrpuTbT6pQDpCC1pZL
B/pwB8Z/ZC5zTOkd8rQLH4RLSMKYQa28gg9s+x6rYNu31QK0t5ME02AjAuORqE5u
giAix0YxuTpKFa2gLZF+YepXMy7W5oBnVhvEPlOkAK3GdPRrRrvF5SIOTIic6id6
ISQlusJcnB8NX0kFxw26xwxds/SRHFtVya2hK6A5Veiyr8jbfBxYuEeqhqGR9ycy
aAFpEmS9KKFtKW7DfDUlJ0D6p4Hx7skRlC+Xa53mtfpYiRU0dwV3W61RzMGC9Hr/
0Rlt4JsiAPGXN3bNn5ON2hsl73QOCETFgU6ekkbL2cyB06JYVCo+3rTlpU71m71e
KFLSBfiUWQWN3R7tGaA5kg==
`pragma protect end_protected
