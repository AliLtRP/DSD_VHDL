// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:24 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FiwN0eR0edfamZ9z96m97y7RICJIgNamzCX+qC3bHMi/S40Vdxg0vYBKPkNk607Q
dKMNZIRUZ/xx0THDa04RCdOKkSSZarOwrQP/4On/DkAbtSmao0smdIZTjwiytjH4
MXFWhG/fTcYTB+IpK5SqH7RC0qNOjBePIGYrlNuHw64=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15200)
T7Ui20uay67NZUrh3u0e9HaisAFe0Er8R2pA/CbDig/feNCZ/AM0U4lEzzof6DjO
5cI5MqSUE4n9bYn+FzB4kFc7XacRMyr6VBpzHl10kk3tLV6cpYxZsIYnFz7D2Pb5
cjftPAVXEuQtlmYbEU8+Qm47TKtZ8cYFRZti60fyhb5Ygjf543/NQTvUppYUDYj1
cdMQkOdeLfh4lVEkBcwEBMgu1euYT4H+CztxtQP4L6bYtW1+wU/vw4YwlMeBTSrx
wEQUsSdcyHPnYS1+m7KjpJlMYLNMJY6atxC+jhW3DO/iWtefRQDzOGxajq+o303o
vXoDHTx2cTvVzKjMaCV6NLdl6qvH1dQz/MhC42Y4Tneo7IHexKO0zswxlJ3VUjHj
q1rXno6itdC16QAKbbviSLdBELWmEVFRT4F+JmCAokpUtz5TQVYQChnMJlp/Jmwe
kM2HvoL2t6BK1gMNkiJfXPdVlnMBgifWuUUqJJw3iXxtZgIgp9DqQtgVA8GjgUmO
t2xU8961uT72nUezCKWmtnm2nhH4SYxlp9fPqWUHG1pJT/mBERHOg0HDihPucYbp
jP/SBe/UdNAFIFFWzG+ucgJsv91Blwpowy5rj1NeNHjubAXJQt0cepfKV7zPFR0q
zsXbJDK3qlRqDbKxyE555xf9nZe6mr4uLMalihAjiZOyqnJfpHrohShKnHuQbdx4
ecq4QJJchoBLX+mdaBl1O2IY9EHzU2QPG0rGVsC4l1RUIqO4Ny1OUkrfwALfYnq8
w1g6DuENnnTYwwOKFKzBy0pzFpkwCYR0dtCwgUj78fbhPT+UV6ZMwtPMOa60LeAN
iL7XYFdzQXPZFesi5ZsBgH5W/YrJgsUQTOJdNU/4UoBoaSvsfDQbiZmO6Yz0Nwu6
79iYnv7KDPmpjVgYmQxGfUAsvaK+xqUBNfafBEeMR8KVY13zv3uiswibi/JDKGwi
+L1L861r8++zWWQ/fIY9ilLeLSwGOTErB5iZzczX5CeEQSiiZgRAQqmKFkBV70WG
fk78uY3kFf03/mktPZFGCIrm/wkRx++sFp9VIF5MTUaMtdEjgZSZpHM9iAViAlpY
m8J2ggSIDBCpCuMN1d7uyGpYoFFMOeNFVmmP2F69nPSzAa4huzWcGodOViAfCeje
FqN/mPY351fgvac5u9PCLeryQddlbJp8H0IVXkKItUOsupxuhE7bF4KGg8RSVGQQ
ZQFHpuGdwycLM+TIxN1yjgbXMOop+J/w/ldFfQdgWLbA3FYLs7Tt+e67ed0t1G+J
brLa9wN2R/yES5RxwLIIxPiLBzvPYlItIpiYNPgWz2hhUxEKC4sw/i6wCNXkPqbB
+PmfdHIH78vjQNGVKOZZsxzEs3jysZZsEF/q2k7A9JPD7NuJDeHA+DgW5Z7EJ1wo
7+naNLT8Aat8Lk+ysBNbia81GYnaivFX6U0cBq7GOjfsh9aE4xPdH1vOSLTfFgcE
G3+5d1avCNNhp98ms27BoMxAy3jl95yPFYrWNCCRNOAwaCPB/dOebZnJ+3BoDJqz
fC3/RvozgrDttFFwBqCajPYeIS9wfVZPs2IV9OwE7x0PuLgo8bbJd4+mqHcJkENC
279A2k36MSHsbLNapUamy0oq6dwrrUyMY3t4lg/y/AgW6bG+F+COPOy9lqQDNOPL
UkiKGp5SbL7DpauUQKwfWh4khYAgXkxzjNX1aen2cr7lndLOh5GOmzvjHM55Gc6I
kGCxkK2UL+6IBglpZZ1exYAjq96GqwC9jHP0mizqME3HleCOKjrGx6JspTkRD0fF
jRMjcSvKdZXAGg58ULtUzzZb6VTBLGehGiXLvngX/VN0zc35ErHl1ZkaQjSvvXOO
VSrb/iBtyAgt1yvOAieEV6gMAn7WxoGUmp1rWOsGBxiSVS9/b04F4NGoXr3hmcaW
Mm5oJM7oAOFyg7Mf+4p/x34SOE3fcmDPZM0PpKbzau+/y6PFNCDwvfZiMju0X/1B
UvZPijODsjRY79lN6YGEzCOHg4hFBh2LcGxONTqCd2esK0Y4EIlc5VSir24PkzXV
heIv9+/q+GF4pBVQPagdgwyq8QrQGOJirJ9AfnGhg3eP8e2h/knNaAf3Oq7Urf75
+wT14/RxFNjhLXWUFTX6mAKI4f4dIoNrtIhmU6OAxdOQd4KAZ22gdOULRd1Twyvk
6BC2I07yfzh7iwN/EnM2nSfFcjtLreNYA4JzwkK16RuvGcC3iDSxVQji6k6JRVLy
jgayF5QHT9w2ug+tKW8O42GKKvXSEDNC0A9EdcYuzjZ1zbJNyYj4qTxC49sWm6SD
HNiygHBQi87+NewDA3dHr4faUOYYyqsP5ZnpxwsuOvLMsBsakYSSROH8x87uNg44
ZBg1/eaFLK7SjrRpfrMkKnp6HiaNMqSB/E/w3K5rmlIvV9hL2O9dZTN50p8vtK8i
o39HynwNNJn4z0qlMXAYDqfXNOPY64JJr+rZtXHOO39/vr3kk8JCYP5sPYNRCBCR
+WpAb9SEf8vuNub/eNsSVRFARrvjGJnD9JFVU5UVmXYLH0kK1uiYxr4IjnsEWl4O
SrCx48uopIBDm2IoY+COvvv65JGXdiZW/h2lkCFIh+pEn1K0rOjBZCaX/L/jgDzL
aiYXfCajkpco0wVluqsf7GpOFyjE+x3jklMiSggcu5paBhZP9rD20c9bGZO9ytsL
0kNdkJCJNUhREIBccyC7JvMmJbWQLPI4YdHNbBRWWLwG461sUU+9Bkw5Tkm7OZRQ
SQNDL+9L+BEdIDhB1Uxazpv3taiejlZbS4Lp+06ktpPml8jvZcQJXSqsmgzohl4P
ecZIvgsCilROn7tVMjUT9PGpZg0WpBxGAUuG8Ng63yIuomJKWPru/YI2J+ZUIOMz
IeThwVCPo2iHdT8GcValgt8/7Bnt5ZaxhQctW1A3f8ET/9BGX61/kFT8KTph/pxn
NS1bSQSLqogTUAVUjvnHkeqfmzdXVZXfFAJCDCBdMvL04xjp5J3XM7sLRECN3RQ0
WSgLgeJx+EEjpo47r/unrAroUFtH2RLWY1vWMqkMahgN59B2NPWVCQ1K0U0RCSHj
32roW33XZzlI+1HETiKFE3PKsXK+tlbvyGmVOFxXo/h8l2a+oNzJt6CyHcnB9v3i
HRgh1doBtRt9bLx158PkcoPugCGG6hra2o1ghBEpYYq2f1y7PADzPOxrNP/AWaDU
UCuN73WImg7KbFMW1PnxdWeE6DtkSCWpgxovOQPBCwhSoPJYKA+GHlczwyf9yVIn
/1VdXy14p613pgbxDROY2kKbi185ZlwEY/2jW3OYnDqp8B520Lp1fToFoIWsbaez
IIWevV/NJT3P0UyUIxZlf2xcSVAVqL3r7PvNCVo6T3C78Q+NxjvDe2HSMkb6grjU
zVKOje0D/r9SdUELZjEmy9LLri4aLM5wtuXOO95QftH7Ptagc0Znw+cL+1BlfHa3
UHazz62XODiJht1WO3k6woiC14cze2rMWOVD3gV+Pkr055YyAfjtExmiyjF2UGtH
mbbZNeXauUClrynJ7vSFj9MaSOsKtmV0mMnMQxAWXr0IqqD/S1MytAGGnkxVIlgj
cuZSZttkGX7OuBRkVPDr4RjUWOKcD1a1N5SmevYCbMKU6InspxEt1rkWB1dQAv8U
uU/XH197DFkwF009oyHwT7LLCb/eLEwceRF5zvJOu5fdYB64Hb/PO/5cMMBy1okS
7QFGNaCJlhV/5Y325K76q9k9nDVY5r0tPCJC6edpqfLMyU5B0UPyE+EzTlYCGCuA
vWWtxpOq9gKBxZ70mHlRsZMfjmR1BufFCz+5OAAhPau3s2zXlY0r+NxoL/ayU4Rn
qVM+VNS0JaFQsEHmtAzW3Ah867PzeDirZPJmtHXOGuHtw1iPFtzBb2hcPp/VFWnO
t8B5jEIzNoF0dBEmC1SdVQ2scFrBjaYcuOv/n7ijuDz8bAfOXS/vaoWnMR4jrWZd
JHMhxiJ06p4mXfrYanSGqBbDIlNuQ3qGdzkGJg4Ou4ILvFb8LOaTU/34FgHmPaRB
WgzaCzQjrkFExn2TyOuWLvaosB+/pO184HxcSHmomXooiTzDtv4sAfF7zOx++2xe
rN/qq+mJOWkPNGGz3vcTy0rlKvANmX0pkUIYlRgb0+XWsQqfysBU4lsee6lxrqqq
mKKW9Ll4KWaGUanWPU9Rr88pd6qWcq9sN1FBB++BPjPxVjO4splphVyja6Rp7E1W
zR2dBmojq16XDrOkSPr/Q6kadcASOtogwRmzJSwtQTtt65oo9R+WZnCied8j1Xud
jFWXFP8KKEEZBSSUR/LTTG+8NI5j07CromidE5g5PZZiegmZT7+08zIKG9LRAS3X
uO5fuBmLIPkfCJlWkZExRykvfe+2IYQrsuD+wv385+b3JmQoQTX38hmrmgtHRY5A
fJMIFNQh2tg7aeBISn8JE4rCHljVIEJ+aro+LIuVkNJ9ki+BFcXIzxMBf+fVTfGc
pyE0VH/roMEGqz8Zw4pqSlnZ4BPADkm/yFmaTry7NKKcPnmnyu+guuyCeF6iOz38
FXYEK0ooET7db8KUEpzC1Fcg+CDqeIotdk3mgRgYZpQ9EzvJOfj47OqOuQFDKYOk
NrV1ZqW/CkzmvCmF5yH5OLfR0ojo8UPxD3HWXjVuwU26uOKYVYgVyr27ylmARUlQ
OrlOgRh+4XrKpA2A/yudmyUUXQ1XhwkXgwksRfurovvNSgO3sZxLnF6IgecVqtTP
3SKf5QaaYsX8a3FKH2Q/iDkrcDyGdWITaJtHREsHzjLO5Bk9LqF0V2zj7BdIUsZ+
I0VPw4rSssOBdQLqiJ/KKUEAPXnwlr+gpXgJnm/vaABxHHO/dX5ZFllTAFke6R97
V4bGevE0GwsftqG4nmexYc3+/8a4jQH/j/LFMpNDQga32s7KCf6VTjTDOA/BiaT4
tq1+zyfOdOVsFMyQzr1TWRBrfaGGlcHm72gNbGQwRnrrGc4J7fjxuk37DrRMAVSl
jS0nW/Shn1s8xZ2JqMRqrtCKB2zT72sdTyo/XStiep/ZK7ux+OG8620kFIgMR4yz
afItvj7xy5iKWD1iWtT1jaWPPLOOG3LYcc5UyxUf+M1QCyhcPV/pId2udasWqyOd
zxR4nEHyPQlcgUYkTcPHY20/OYdgZGcfdVsM5Z1VcPud3m+9ov1Autoy952nIbSV
Rt4Vgdl5OKAW3T58y6dmMQKqZASOz/YwtHOQtv1uE86OF2reyXgruhOZ0Xi4E+MH
RFL3/iE1b7yiVm1YQ9BEwzUze/UrdmCdrgH5bozkR4rr0oYyNpWXwYh+U7xUK1pl
YdFdkTHCiL2w4fsCSp9jOOSYUDoJPJ1W07192bcq8wpD1uxqG827wlvBHQ9E5CQ2
746rrQZNGIj/PoPw6pEOKUupLIkINzjgsa6vnKEKsfe4IaMODMRXPpElCCLAnlB2
jeXl+8TFI9eek11U2tyZAdV8eRqd542malbOpRXO20ob7eAuDdyNuCI5ccas1exR
gsRJuCCh14Gy6dJ8ohzIIIRdejwIE7uBcshql7+wM3oNDxataFtQnbcNKcfvViqm
vkuizAJzQuENqSnTEg+/QUcq/2WV/RibNuLI2N7bgVv/O1pM6SG8pgYANmbmGaIc
e7aGZE6P6TzSI2k3wJPWsObtj+h1599b3pu+TyWbQSZSlOQlz1CKSsGTwoJ2RqgW
10nogbbZz0d7TCyR2WdFnw2BJjjZNTDcug9HaMp9/YP/+uvsE54hkK7KTd0sa91v
2fwfv7osLZwjgRyCPvaEgwmQoEEXIPUHv7Ua/RecbLMZnfu5Nfy7jUgQ3l8w6csx
1fi0xXK1RNwvv6lXJKR9UtiCgBI/8J8uoxghe5wOxp9VtqqfGs+U4EZeHwEvFLJn
rFUFeZJm2zwnMF7k9L4nRIHp760pQmfhYzmEBKiWmOYb9AKpdfERMHjkyK1joBch
TKUnD4rXpozugdQqx+xlqvVIjj7mgOws5rpBus3QGpo7foKSRtjvh/b5FC3494kp
yraG1HtDANeO6g6mqfmnUllDEOwJI18X+IF5y7XP1Cpu9+Za4PIwRbBBg2dMNRlv
CTLmBiu8CQKQvCIVyTN6MxR9h20aXv5pM0u383R5vx2lUFn+iamycRm1rLO2CcDe
AejYDqMOKPi63tvZQTWcwwbnuZ//HMIT9Dcexg+NZPH8hCILGtzkz5yO4jq/AinJ
Dz35YySiw8qt8e02dGae2fJpnvVEdApcoqVmnRkKiHD0fsg6jeqAd+NciwgU+2a+
G+rRByBzPJR49X1kIqBXOgXsAYV4f8j2MvVjLePmwucgE0N7qQPjx3G0RxA7iDLS
eMwaYv8ey4YSBVlFZ5Jg00OHfd+8zplyZ+1xllX0Zzurr5+KnNbc7WEzW0QzV+OW
tSvamD1UnFZrbkfMGGF6jr188eE9k7cMzwylCtVM8k3u7NInj4FymX2DFrLSCUEe
y24iLgsaJiI62+pF5MNfN1PirGGb7K9gYcNX8X68e949UeAL+IsEQoidfOvL++8k
zR04ezyg+sgNfVFEZDdqsoARDMWvr6koD3w2yxdBFY6O0dJrhB3+bSZvXkyx02vj
DTviJA/KEelfmfI1PRkYUuaYo56S5IskG6N4Pc6oiuiI1MT5NiLnRyNdDR1leDYS
QdWOzHDTeMvF1PGfO1VUIFIudS3zRNw3PJ4VOnBfMui4+eJL1llIi7/+xM7EyY3F
BZ+wYbu+HuOtaW09Zg2UsuJoMT/ponLP8GdSo5mHN5qz2GP51NlNpL7z1gbGdWWO
PHp6nfH4ykrYjLuxiasiyoIXe/NqmYctsh5s6luFUt+TdKGHKh8b/Rf0jrjWEUI0
G5bJ31hI++VCadk2KdmER+s4grI4aojO7cu05CP5bDkaZbujn/Qq0hBNs0e40E6C
4QUswtr9/Tt0DfB7tQFvqUNaE1LvHoywLVnLa632ga0Kp8/xGYu6SW82sIOxo972
mNYecx7mKjyz9YSSRELO8uH2k/AtIn8wF1sp+ADMhlntKCuNQk0f3L65fm5yARUH
Mz/A6o9VfzhonqQqXkyLbPPwH3HQnjWH+63CtscdsrNNKD6xy1jl4P/OnZg8LXgF
h1e+mwJzqlLTW8jBD79mg5IPVgsPIdSDTS08slFeYKsd4xdMFXURWvvQ8tjSflql
U8dAXsIYjUHIkZtkZI5xHagfOeOY6lBYQroLUL6xywG8rKvr9ulsa3hdJdguRaAh
BXHlTbX/evorep+cQd/yqJmXG9Gtly9h4WbnS7FCtZr9+5KeVSDf5LIcg+/44h3C
+9VUkv2D1RmWp8XcwvJgMLVXFz/KhGeh+uXLwg6bYpezYCgZqlxWIsQDe49tNfqy
+caP/2GQ2sfeZgk3JhsjrFEce9jyyksklwh/xBVQ1xxU7q6Ybg2Vj00d/kWZ8KUw
hMcXMi0hAh5GLcT/ZaPcigjUbCodDsEieZdsIV0CUfJky1Xu7MzZNs3osGPm/Ufd
1EBGZvT3L+qwm3FUuN/fMTq74TUE8odBOkHPaNMLbSrilXStzA5LSv1uWjXsKKa+
TRqgQHFVM7qpkwXAKdEG6jmVqwj1OBSTDFIJx86vG7X0BY/V5LDrSfVYIP3ZzG9d
4XdeiqIJvjTsqXuwg4+24rP0Vl9H82jAfPMCi2cLwhGKM4LFjV7hyQTwOFoLCvO7
i/CLAMGO98kCyVa1L7YhKBNhITQ+hMzaG9DQT2GylLLorLEBkn4YNRdch2Ld/bne
uAMy1dVnOR6Q3JMBUFgHg8SCDvT7gwsWyPuS1MSar3Iq6bx1LojKxUKuvtyNcAOK
YKMFKW/ZX+yBGfEEFoN91W45aHuujbUuiwY2bS66iO2eGIzq3AI6fsxH60x3sPVY
mK8cVr7wJquhldWHtgfE06JMg0GKdjKiT11IHl71Xg9fjqO4dUGqsS8oMqsLpj1n
/sdzwnFD/tmvfnS7HQXL4aYjFEQ8dy1mhRbOCJmG7flRiMfRgi+AZxkMY8rsW5gw
974WfTN+c9xg1KOmzoWJMRUGxA+nyav+CuKzORc/RV9mb44FDEaChGmp0mN4cX4J
WESA7+DM3z/sV7PCnJFO6podi7eCUZBkNaMMFCo0GIUxhHkTQA4QRlTJZClYMO72
ciPN0COf6WHrbofY00lzNTStWMxlP0+injpjOrjcj1vN/hSNkE17wrPirqejEkZN
gdsRd232PGhLi8fpzdiUTwJfwfzmMxdcexryilM8yx0SgwdnR6Emde5CIxerMn4c
qNfbrnHLEdX81hPYunpSDEoQVzaHsxoiOOCpzkQrGXaV3/IiXT7pavSv3WUBIcs1
v05yWqvwbC1uA1JxhXng9P43PVY5wahzNRlqEs4r0wJdxWvrrBkBIbfp2cMoCLWc
UuftuCN8kwF+UBUprEc3Z2VsqGtsWZcHrLiomjQ/EaMS3torvMOUfdfzVRcp4b0X
NB3BQG6YVDPH3AUhpAgHtDZbL9PSdau7SIQaZDzy/S2D3qNvKAv1MfV/XZIN7xQ7
fmFJ2YoKMAiw9HCdC/9pqEUVf6LhB+pHdQC1usohZ2nTKNO/fVGnZ0AM8ssFJo//
Vg3pVFeWtYKlzVb1z7+whoHRWqRzJAjUXBhvahdQIePqDflZpmCofdjrwOROTSw/
qB71KMqQjWNid7bkjEIDzw8nGgMoWkWO/xgqgZKwWICBfq/h/cs8kvyUXbxI+37j
8bbfjbtjuRqUWaPftGIaLEOBYUlssEC7uKY1pQ0WsxBQHHXscLNo4jD9WXnR4MKl
x9RsAXalT/mw+D3OaykISNhHenrwzq3FS837ly0syooxCRR6GfPCQ/sbkjT+1KJp
Skx0oI8+unIFg1BtkS1mnKYde8bSVy3D5OCdFTVrFRR4+z0flceTGRF4LIRaN89W
gH5RrYgGtIsl+Bjfc6Lw1CcsOfRez+ltHPNg6mbVQmyiNSI1P4C8EtXgG1HpHDzY
MgEz9PObQ2VQKd9KxDDPUPGf7hMlzf9CXEJ1JHmf0pcZxBXu9YHgWmn17prBEc11
Ykt7Wx3aOUA7aIjjxxQYhCEmfmuMBfHLozzhz0BzgNN6QVJe8pM0A0NEpbjAregw
dYWwrQR2N8bRqCY4IFTW37g5ZefRogOQYso6gmLlOfjW0Z9m4t0WseCbMxrQKfM6
DAaitYPcYBPY8cJ8rJsRk0DLr/pNYNEix2UyXYCAJROqRumKN0BWvPp+OT/eXWie
tkmZ7YE8y9kvJv8lqGrpfpXw6H2PsB2oY2XzEw0mkx1tsa/M4aGha6RmvFoZHtcz
tlDp9MGg1CLc2pfeocMy7CbZv+auPwhv82gkfWGU+LQn/g/R2aOwwOazaU75tkNo
dMKcZh0/BtjkuDp9BIz8NMcEMuE8ZVBbcWJMVo6RD5/iG4uhHG4vP00kl1Og/t7Q
CYCTW0YA+6xhzBNLlJYs1bOwFAS9XpasT3MyUqhqTRI4y5Mw8x0cig+ReRxHffGW
KoR+kOybb9hpTFbXrSVXL9MTWLKRJolxw5Zn6SbwlC8ttqTqXrQbSKi3grhDVEMr
yP7y0rg+lo0CYIGlWOnJRlSxClbUiIdr2x6vuM/kLxDHNeCZrkEMTDScMppqx1Bw
+TFS9FUaxuifDcXwPMkeQDucQkqpMSi2J0hA1OFvs5Pa8MbLtaQvtSS7T46Qk3gJ
9TpsUghL9C5KRmmQPV0pkBCCmo6uA2yrn9RqsADwKiX0IkK+ndR6WszT+pbT8iRY
NnCpFE86BFDbIZy1RTIhNHxer3iIA1bUwtHPb/+cSOaZkZ/l1GZ9Yue7JFThA1P3
N5/z3hSRDjnt75XsfsjW87Lxhh+9d7bRaY96DXbeG3woSdt6Z8KFMTpH6V50sA0Y
6PCOHsaCQwKKHD2CM3NsC1x8xwBm2HefHOlaZUiFzumE86AXflKksPiIU9meZ1y8
XSerI50y2DFUGnm9AAMJyPo9RvG1GgEyY0HXlqswaoHjM+USywBmdRmdwLzqc7zv
nKWpJmNkxdy8+Wj9YrtG1GlXxPUNuyTxIFt6q9b9FEoqLZaG9LRKXiyfdGAo8OKD
mxnTHTP/tITXZRExQtYXwBb1JbBlTEgdK8rVS3fQqU/yFMHEg0LwtIHofejbGHez
+AVMNTaqncZ96LJXMzx9XB9cSCLLvvGTwSbk7nvBbxLV8tzSvp/ZDYfWPCNrWITa
/iwwL4+fl7gUUQJEQZlgsrmLOGrGD1kDY/oMj1tNyYBfta1vQaXXe01JlGCZ1GlG
FPRNwhjiiFt/j10DOavYZ+bcpCFgwxQ61k1x3JO698PpxpHDuFEPOkjqyadTG0wb
7/q0Ic2aWy/wlsPUu+3FvL0HjNSCZk3gXWyiEYZSavySZSrrdbP6T09mZoTomGEL
Y3QAnBQT/BhY1kqkGJRelJxNNt6l5zFrR8mMF/IWDDvCm8I6jyuzs+tcqDsrtBtE
4ZAZqWGmFjt90fULp8f7i7kjpo5kixxccI2P8mxpkQKDTbjt3FCw9DkmouyCq2z0
FyXsJdjWTs9FMpreABu1w4YReTfNE5pSGtlQGHl3s3Dsfn73KSufUwtMQ6DCSW1N
A1BOuaOeh4wt5NR41LejmiM7NuKOFJR6s5gtCMutGBFZ2SYYiqroioXwsCDrQ3ME
YPcD2swLIuOf1+W6BOD8LE5ZTTpkUclKg6M+CrvPUJK/FEa6eWyb96kBY/LCM+i9
dNotLZG8H0bUrJOUInjAOaoiUYa9QwEX2R6reQhf0THVYk2kTQeNlYqTEpKHDZPl
kPGUZtRG2v3mOGuEX6XI++pFKXMwxCmwkRR3VvVz6XxBOJsutfuv7lAVv015E0ri
jAAkEmihqkC1CwJYaNAaAvc8KWGEdBS02wrpb6BzFVRywBWH5muKECpfp6s2UmL+
JIxD2Pub1tNgnj6dINaBYxAKpBWhR7phms7cM4/AVI0LgvwEYiQDpIWIaol5fKJ9
xqob5N1L/OOaZKlcoIqK3Db/+bBXE7dt5Qm69TNwn/UaJ2kEwkcNze0anAr/GJ/i
nP84C93CiedLnLYv2HHy7DijHxaSJNxf4AugKgeizvt64263ZfmdWn3Lel83QLKb
aZv7y9ULxm4JZh80AhsNaTtfdxaryeFXJs9LuVHh1QbD8wIsnwTSH+L9LH95+I0J
cT6xGFvDMstYDVYPVlrO0wUkd69op4o4Sh2eFJtd0rYOpu3vLsRS+PAy68KP0nZP
zIvKSUODHs5IVzrF0vvxarmRWlVbPyCCoZqzMHzWoeEfmEO91DTn1/5GldEqotRj
8P0Z1g/Lw++u2WihCcomqP1UhE+ropTEa4BdZmL8T6y4qT5w6sE3B9UXrzjYWYIL
jIoFug0gIAIVbq/JoK6R9NdauxEpA+UlmDoFa1jXlregfp0X759sEbhiLfRY7ecp
DqKYp8usqPSWiwGi8SyRubjTv9SA/cTTtxNdWwocAE/7rKB/VmWJkq7M5csNhWJ1
5LWTnbpGm4+YOwwVlNN7qHjeMUxHNntjXrWJSn9laKh9+DbsyqgGF0mcTeP70RsP
+SdEbESIolbprWXTXruMR01M4KSyyfe7f0F+WufKWQeacrb/oPkOOMLq0aUJrpNX
xZsD9pwi49ivS2z4MNJ2FgTACpJbt8Mk/97hkmn7QhCm2BJnt8aKafyBkEqt1X3h
S2i+M1woy6zDOpxPfoNdNZfJRB7ME9O7EA2c+v1ZSQDkLIVa67sl1RV76B6Kbdga
b6KQQk69gi3HCcSj/+OXKssObAt5yn9bHbezC4EmpFHp/34EB7tgliFsxiTWU80c
xUDawodMSNhaDYJL77opMvagaSkbt5ceMIzzLsiCe1Z6W8y/f8pCzE8Iu/urJKLd
Yfbv1iw0887Vm2COgc2QBdyV5B+CNPQqF7PfyJ/DAV2fU5GRrx+icesOi9xUbV5x
ODI2EwmfISdmvsBN3q6j5uJr3/6OmKpfm9tl4UhouPEOw46cUg6K0N61rwo6wBxk
Qv8tvHXTtHEay/uTJzd46QJWN9cLDkYr5CztJLdmJKO+XvmhcYLzT6Cmf1m1N3PW
prD37e7PjtH6+hpVJM6dAiqnMJxCGSAhVaJBVW8gw+ax44+G2EGs/vNMv4SsuaRU
bRoVqNl4wXTkbED49j6+ki5igqhmU3ypufNuhhJDxmFpgMCBueWcBTkMsUxyN7zt
nrm1A9O2lGL2jho5xPstnJ0FAGvLCzHwv5vcjEuzmQKnkZYkgZrrf6zW9rP36nrm
zPSG8pG3YyPJ8GhBD1bxBrO6FR7i5ShfX8IM4DO40pEklllYIrMZ7GrOMd4lwtG1
eSvlHYL0CqpqtT11MxBifBC2i/Kkep2FTxxxvIZAOIFJ1PMSSMblXhpvQPpSqvma
GokCkWBCm3Pa2q7S9h53H8o5Jeonq/+GV/94rwZcHpzHGKhB/4C6Tc42q1nDbim1
t4GzQb0/5PcpGJLyDnoQdG/vmqV0rDiFZoE8v4R0SdbLrZynjlkOxTEUO1Cj1mtk
02pBLLjvFZQil/97LricIlFqZNdyED2AyNEoJ1CZBxylOUiX/Uy+kg04NGJFEWOn
cuJmHh3NP+rfLaPU2SoZhegWIP/UBidfPKLkOXDNvyXJYZ/g1c6A742Z9IqNkGCR
Jfm4DHA3F4IJiWmJkSRuz1GXnFu65AoyeoEMqgE13q1v7OJW6vPvRAQGmlqgL6aQ
l+eEBiXpvSsyTST2jUCFbSu29Spfx27ecIlB6yh07vgord8cyWnpT/XwMgiZCgQZ
cipC1q+3RoPd3gih2VcvY2DLOx3V/lqNF+SIGJRXzQX3AM1Kh8pzyNeOSHfaxPtM
ieC3GmgmcCF+Pxu7cxxk9dnXYHDL16OKvReXwt0SBtW5yclPvIBu2d0bY1rmdSAa
1zCMtrVMfj5nDuIjJXC30ZQvvqm9IO368ZR+MRDAn+1l2yUH3s8+hCyWhYwC7Es3
660pYWkf7HJ8m8aajKeC+fAwY+VSloUqXrIiVMYZ5fOxlHMoesU+rcs7fos2MLUI
HC+4VJdUpF9PPI1JIRqCh/H0syYXSxs7CJ8v5/K9BtGnyz8e2rIJuBq+tRiLaRDq
DMdL4GNB6Z2mIBy6VVTQgXjk6gftB5rw0JqqBOvh/vPtIsg6wEVK9BE0TKrHKIWT
a+On8EsB1CBCBQQLUt2oQuF0huOnOZ7NsfzGOk7ijHLI8uQ3OCtQAlcIBbptZCe0
BugV8VvS1nlL/l678k/LxR5+B7mkcbIEZNdhye6w4TqO5MKfJeLo+q81Q1Fm2VSg
j0rehmpoQxbjH2/LtzgyhxhFhcCp5WpfGaHTvCh6wY56xmzszPunTE5Fsnk5U1Xi
oJUKqsgkefs8w7QnOZhMN4NUn1G073mhydl7rdItiHrnfvuzf4E5Pbv4KoxCJE42
X+beI6acfuRhVSnfHQxRdY/un3ECOljwIXlRor1CWitlmA0cdkDm/JAC5ZSEptVU
owPyYjdFAs+J8cwjUkyWs9y7Tg0tuY1qujLxEpial6Pl24P0oA4+VgtQtQyccnN4
g6kW+PprYf39xt8O5XpJj3ie80mqyVCSRZq/v0NmKLBnkvI0MIt7v2CaSc8tXzex
wwhWRP5kWVvGXpRrILnMixBA4ShkMMMbJKgaAjgJ2+P8qgrLppFYSIkoBUlj/QAn
sNSf+j9ZPrH4/7MXJnrS9YrQaNIA4oJQ6cHLZtMQbVj29heez7WkNjn1GhR3LFQ3
j5LEk2J03w42KlK08ZBvzaRSL+EJajsrF0uvi8d8mc0H/2trz6m13cWl8eiOSQtr
MmvX7EEN2eUo09KzPctFJs8/3RJN4XcUoSJf2Ku1PQBZOJgJ6lJvJHwT5zdrkcwb
zBaPcPClihf/a/IQWT3w4K4icqV0YcUXSxDLjDLdb518tPg07bl5vxdJ/bjOotsp
Cv0eaPLwnZpUYn4EUOVJr1/5LFszIT1VLWckpZUsHGGu7J2PDXeKHigXuYcrQxCj
4z6l7rCWJ4m/ZAwVYuUu00Y8X3mnJjulpbPKJT7gW5ya4S2IYFIJRSmilUuTnL78
t4/gHKhOPrOo/ZSjQkZFBW6aYmrVDaZx1FMqSmAY/S3639hr/VQVAQ+TbcZZlDGX
qF9ANxhH/q+UwWrObe5nVVN8EtHt0d9GKsThMu+oNGb4juKCAbj3OWWTuCrnoW9T
/oLgNe04ODO+SXHE0dig36rD0bntt+iNVZKVjz3e7tD3VLbaMDfJEl6pA2Ed1mDN
prRwiPMzEIHISH39fq2orXXYoMVlCTCfvZzWBEXzLwMIOjCmJHfE9fkAYYjeQmb3
TxcYNp8JOnHKbzKMHA0KeLpL1sKCzBaQce51OiWX1xL1CWKJOcliMRuuhAd/mbO6
GW9R+DNLGPi+appCJraz6H8Jxk7/gAubP3RzO1yfSWta+XGAWjGfM+QATPAoyOuX
s4WujOTOtxii8JNMg+VO8je7qM6i4woulZ+Kdozcf0J29U0u+lRLkYzWDabLyAEz
pmbLzZSjsy9TYZvhdf2fj2kWICJ1RcPCPTpCtkKIhR0RaRQUZPeOvrIu3r3M/4av
qkru0/orgs5NOgXpqUa3RJ2Vz5xua169oa/qLZ7/+RORrmonxyk+PmiMKuRSwruP
X7Dkiz/yr2qZF1y4gQ9tSdWNHhddRUq/N6PwRUu0DTA+6nJ3oLxZp1p3qajMhJ49
zHW8PHsvvD11JN+1KFQCXX9lxh5L3TwIgRLGhoLz7Rz2kfKzX+d7E9d4ju18uywh
um0uuDaOr6rcrcMtvBzdC/fSGj0EUIq4YoBcZU0kLjz4rmsWfyCwlKbgnU9M9X/O
50Emn7puxDBq8vrC42SLOCRLaRECkfby746rv5mpRElmVHpEonWzIc2iRfx8SnOr
hGnazLdKhTLIYsT7v1X2TzFPIIxlwU0hDK9rNTvKK2XxMJ+qpIEJQoIf9kUBTa5r
1CwP+rFjK8eiExfLprAciuUbQfFYsQEp20urcICvHqPCQxS+Dxr+xl4dq900Lq1E
LE71SG/YquOgJhKM7egBHki3Aif4N182L6UkGyzd/7eB5lFl73S4b4+TkB4a0WH5
dEnlzjg0iqbuFgxSugdrkl3ngRrqlu/dFYL7SVXb1w8hoYaV9ixibdqfbAS4Q1pb
zo62C3fL4Z+KlOeORiZejRAa59FMLpXjKDpCIn7VUOHeXedYMgtI7DFBYGD4SXku
AkC2TzF/bTX51DnAquSLa1rSw/bOXpGtX5rRS8OvE9vEge8rrrGoZlWuCDKjV7g4
EVyJ1DBNCvKhdQu4SI3YYuHnwv0e/djVdxjBHllyqZOsYOWlb5mxDURZrtw2d9Wd
ctfkHZ2t9AcUU4aBfmqiNbqbZOmhvDeBZ1KiE4fYxLROUWV0GeXGJp58m4grpNP/
r2Ckw2dAeYv4pcsYDDAKI/7VEmN91phjgRpmRs+Cian9Rdp5NZIew2ttVbE3c81Z
g7Lh3Sl7VTe5mvB/Gsrir6r9+C67OopiI24xXsQB5g2z+JIoMOqNnXTFSLiKbkEL
/I37ME4Tut2qpRgLZWfVT1qfcFwMryRPG1n3JcUEHSy4hMpwAG8mvVDHZh83Xg46
InCqt7kQOl3xmXh8VMHF67nXaxMji7sLuMrbE5FY2Q0UpYb+PQOGXf/I/EUiLwTJ
u5wnPzAiQfPrE7F86M78OCaaEbLCqiUGuu57OUeIis+Tl6Zz2ukFurWUQ30GYN2Y
gPZFp8BrBfsQwtnFA+LpgJqFlIBywprQ7O2a8dKfkw/UwQ16GGgfVqfxWuaXpTBY
h8lUZZr1D8IfKyD6eJRxGtCuE97snFIJTSnOLrE3dJFw8IaeXQdDXwcDb7OGUbdj
QUTsTKrPvlKU7HBOJf6vARYXu3/NbEEZXsXs36VtB29ffaPTeq95JfMTYBACwhP6
+PgEIjwjKUWX6Z2lNZJgj0S3bDv2BkrHUczm+J56mU0JSTrYs28ivfplcDbNR5dk
Tvt9b9h4p9vhuwG+gaCZRO3YrvWfCyQTD89iTqaelXgdZU84fk1VR4R9PbCBLFfD
cbW630Pbb6z2HjhEQ+WJGCAw5nptBafFCyo4GNBjhz8O+CM/edU2xaqn10dP9pj+
PW33jqyj1KlzpZRSnmbHIjXH2t1gKyFh0XuPviG1E0SDXX/zH4vAPj471bFXjbRB
SUVd0ix/0q9VYbQF1Mo/zFiO5HYG+qWn2DSvkqbCAYb6Z0FwfdW5BmdJBW6mpsDt
PUw3Yl6Qqo611xrdik+rilgqC4/m/VKv0z9gMHy+EfejzsedopFE79J5fCTW1p3F
gxj490psHwtKeAjjsqvc0bY93WP70PsSX89Kt/FDwG4HXCHiGkszhm34iKAt6tqK
qeBUHh9C+tiL5b3ZSqrCSKqEipURRGJM5wVAlTILeq93/mLWW93qQe/brPz2HhJX
J9EOiqKAeM2ftVsEJ4ZwcgaaCvoQlSZa0zn9wA2p/G05hWkLsGIyAIOuxcvWa5r6
0xll58i3Uy6+hLBIKTz1Na2qQvBQmpruaWpnE4fvGs4x28pyNmeimM3iZBYDoU0z
mx07A7kSn+8YRBqGoeYnfZk+1tS0rJKBfbl0U8SUkXswKDizh3TRA+FC20HbCx/X
Aawt4YTe1x2OeVD636lqkJ3jlChsL/PzneFLshFI7vCHqRsMgMjgSLLgkTe7n7Ur
XD8F4kCl9xuX4iUvP5TPWihYS7Fc8T7pE9yt1EdyAKxcHD5G8LS7wbuDOLVdufeE
aRVNG6s0OFWtUf/rF2GVbc8brcRwjJFv+bDGfHlq98WvFcqtkaG9PnyEsTcWdias
IpmguQCMk1Trq7JILgQsW9bGNrCNR06fmWFWza/z8ZA8VtGwFPhzC8n+FiGhyuQ9
CNDMUjQz569F8ApmctqxRuDByUOBs7hbRKDK8vzk85ifQcrg0FhPzfA23tR8y/wR
6pZBuBkD8E8UGY76ocB2jvKQJYIdCuiisUrMpUCbNSRAeqXFk4Po1K8gqxFT1Spv
0T0g0hFHWx0VMtSKxIkzsGC2D3AQoFx9lLaXBrK2PuYtRYm7HbCT+3bx1JniifcS
CIETNkeqSA9WHpo7tgSDdfSyAWlRqGBaVr06Dy/O0dFK4JniXIzc63bbPFygCKvm
gKx/U/CzaBxQH2x335tMY9y9EmwEg01vRx5j7rVypv5KceqXCOgfimOvjor1Lb04
k07vHxoYNqYWlNedaiQUmSBEXUTg5yVgHVcmYSaR/JSUDf9OQRCPTMgtkyf0/Apk
IpVxmBgmAm39+rGslIxgXqwwf0vAZv0fBAsC5bbhLCB50C/D2R7WN6U+s+SEQCK5
ZfumhiHVZe2E4G7d8iMIrA4KPxBZgrdNm4P+BZg9X5DhZXJiCHMWz1GhGeNf9/Az
e7BuobtRkaA1ux3X3usXV7yfFTs3EvB48JHtMIqXLgBMED8YoPH5CYo3cediEngy
3XPRHUjhy+oMxi44q9Hg+FzSUuV1CilaaTHxyXJGRneE+3Wi0SpfR6FP9eC4Cag4
3O4DuJFLBNzLN9FzUMAcD5L/4fZCIlNCykgiPLuN8v3FWUhMGzrfxfn2ACOvKfeg
oWOLpxcZs5HWvM2+yx1FFkI7D4ycERoAzCTQPS7u8ssOAkcHEewqkaltAfg3Uw2n
fYSyCeH6l6ZXK+s+4ZmoJrVcdjbWcxrRnAZ/V/+7LF5O3GvXVbrVojZOirBAZYg+
ZU8y62+Kv5KBzs7II63lsEiM1zJ3J1ZMtPRC5116+95QwCIYC8XgH4PAGAikfe2u
eR3Kj12/tddzml+I08WbbbQ9VoJ6Bg9RwGexVSs/AIyheuLtSJeGydo0e+1vaTKa
ZmriSyUTpM+Y1PDgZfkoxe5GDsNfsLvn+jIq5idZm+sYNGkHttF8XT/gIPkRWra0
oIC8LoOruBOW7d507mjXFKolbHJm20mpEMhzxDwzLcyePnkpNttQarqTVrvcIip7
lA4KiP8MVySAmTUEzXU4R44J96WjjCee7/Y4m4eJpmk9PDelnXxKBLA/70d7i0ib
YicxEtM3cPPH5cG2Qm3fFV2BNArMLCPsFDoNlungwAT6HoFJuxVDGFiGgh7fleUE
KRX389ywRLcsH0rlHbGOso43nTfOHhDMU4BukGJQpyV+bz3vX4HJiDHYHi0/NYg+
JCvDN2Re4+bgsI71Sm8uM42AsTHP1Tcf+NkUWm3VQUbnO1fcL9qVAGJbtzDcEWz/
gIP0VUlOcy75SW/HPpdUomI3NrEOrM+agogvG5+tPyjd40Wye/YXsg+POvk9Lz0M
C6bmH27t2kOfInmmnFC+rmpz3siIsyO3Zkas17tdIaL31BIPZJM67w0iLgJTVLA3
JkbYKxFyrNieYG5hWA4vHYXDaT1np1jxenG/Alyocpnx4dfZ5KoNkD19CrIULtSq
8sZ1qJvm3ftk+H8Qup+FRM//hrAtDx/o/xzSdaU3Bvj9QQhuptlX6D0V+DezGygl
l/byUOIgrUCaQr5n4iX/l6HEDiks0zb8k5ijO/sVNnpdNY0ho7UGbMWkhJqJVeg7
uyXPqZwpwIGSbB7bEaswqOMWUaKRubos9CwAW7TbtbA+kbe3+3bqyFlLwukX7TF8
XWVoN8NZMOaadz7vS0WX0obGhHCYZvb2DOtsIwWYutVwmERmQ+ZBdqNMVMfGlZM9
eilB/Ap1M5Ne2wGt8uaNFi+D5MNG8OsmVjYpEh7CvmFUFZMdtQAlD1kb4LpCvn5X
Sp7zjop3OHYLRe8eYvf3o7/2sxEpNVNxWUEJ44dq4ssjDdq5WLAa7n1iObqsRROH
8hWsIUSg8AX5A7x6Wjt+0Kkw2F4yzSM+wdcVssJghOCn/xsjiO9N5vEyNls3jQrB
/eu4QNtV/2PY4K2U/KlvdO8T58ojhy449zGSJOH9luDHOizaGB4PbyLZa+0nGcSu
B7lp61AK0IC8X6tVE5O6AsZLkxU2h8XMKMViv+/4qeX+FkzbyktwKV+8EylMUL+F
dG64Me0gBISXH/JZaRWxlPkP5Kkgv0mGhH71btUVvzhcBatgQKBo2SA6cpQG1r14
nG4pC2FseSnkr1aTzZjqxHFKmi339BRjcWPf0osrX4SQjU4ke4ne9ir3r7A5TV8b
8LPA2QIkzUDb0YG2X97T5PaZApteNDaC4jC6hHXEeVsIz6b4kGAcOjLSzN2UEwN/
bzKIgp8Pk3qc7EWsUs24LrRBqfuVXY6nA6+P3sSAij25IR2MPmQEZSZamLNaH1K3
JFECpjfbvGfw07RCEC0L5o3RjMZCxm4N/0UoKk1qPg0J+8/px9kDCm3yYOAvYt/2
NVsp/8DIqnVCkBjC69IeoA51YM3ZXSizO7IetAEv3vcntdh9KX1OWDAGzhNmrD3z
Q4a1E2vTwbNlGS9ezBhX+PIzFnjD6qInWE3YNblvbR+Ag8eIcQG7OTVDklLRnXHH
3fjqIWZcyObfGL90Qv61CNK0GYcGcfmDD5OeTDreiS5VKyz3aPGnQVYhb7jfUu05
WiPKP35YnpI1S6fKFIYRJLl4NjUfLyp7MOYn9ibhS6cfUFSDJlxDHFM45RHiITkZ
9dJR9TyEWB9MhY2jwaRAq4D/YPplVvtkdvzT3nJUeITRAnkIlAe6T33biKpirIK0
HyvPC16q5nMFCEUjA8crB4WsmivJtqUd/4iE0tIxgMd0gEja+tyHA0/G0GV2uDpS
Tg74qPubqDgwpGmR1xNOf1QzzWbog1UBflfp/2mUe2ZnXEsN2O0BdKO70KnSiGGr
rxYJ3AxzIOo+GEw7wZqDuSqpfO5pf8Knw/OZ4fyBXzwfdGwk1/c9sPDeFoo7RYnU
c0Wxh3D9bL7kONvrg0L3ocnn5BS4e46aHwUcm6wy+q0k3Bcv+oaEyJYcfj1hBRVC
R3GokyPimNF50/Qm3j2nW+W3AKeGnqS4QNcc+ClYtpEHhwpmkw+c4fZHUhmEA3CW
5hZKSm/Pj665XwUZ1s9Ge1ARpDe4QGWjT9YPbq38aQaaeWm9EYFuMfLAiNkLkI8v
BnXkOQqu3FZSGeHHBvpchb1D/6nmIrlybhkFCFh8GejyOPjpuwWtI6TXtVlZRFdk
h9xS5HO4IDTLEkoxFGcS9dDTF5DYhJREC98pZ/usDUotAvlJb4NePPBl/qsQSm6N
+jB1L80pkjiWlA3PXBlUjrFx8a0/sRaITsjllt2jXIPgXR04spClz4A0eNxpfXCZ
A19a+yKaFc1I3N/tyyUSJK9D3RCl54AMZKYJK0I95kvN1W02Qv/kOXVc/qvvTC7H
cYDUNZ/4xi3AXln9E0tdrl/q/HO/fza/f3Zlle1/MvA=
`pragma protect end_protected
