// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:31 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sEVAWbHmNI8YF2QiAeQLzMaQqkeaRAD6QbonqTMmB6ly6v018Lnf9feViaLb2O5N
xsGHNaPncHh5Bpnsy5MywlfnCnuAM4zrUby+11H1Mq9FqYPz1xsXVSc99RQMr4f9
7JMHjFJyQi4VQCLo0y2K8v6NMJv5LQ9iaHscMQXjkU4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7280)
2NpFPHkz57/48jc//zy9Q+aMbdx+AM/15hl45dxRgXsKUWp1xANDxnWlbP++A/o1
4zS2ADa/I79Muz7YQz2pgqDnd7I3je5ZmdpyuidsgYelMicqiGseJBiIyuEEk33u
untaFPeh+4vBN3nO2k03haqdL17zf6bCs3ikrDTEuLMqBfcsYOy7CSbMiQKiPVa6
cqkrNYwNhViUfSMY++qEexMUTywP6BD76igcbRmplDCpDjsKckquXXtewVCj1kk/
QfN6R12tVQX7+Lor1iOpzkc26AILLOUTm2a1LU+zX31we9tsuOMxnQiVyB/yakwL
pREarFvfpYXRPcVrAghz924iG+u4e3HtybFi/6HGaUI7Hxcd/5cFWzvVexDHcnjx
6+CR/AwNy2Hdr4AFf2GNqWmf2Xdvd1b3yeInw1WC0IlmYiKr6cOX/sJdGAWhE4wj
Ye8waEcAtZN8x9Xv96mz31wo9r6rMyUEZ7RK0W8+cZplFqvy3QMrASBmxDMKvAQ0
ZrnNrwiMCwsn0JNLRKp0wGRacUmTlZbcNUhE2KSESQGDGMxvgpsOE2HApngfKaQ3
mqBTs2VV0NzrNd+il8lC5ccTG8ThbVe4Lg71ORc9y8a0QfCJi9D4pIhXYtgZcONt
djYrmD6fkB74NtYbIaZKxOOwR1VqcUr0SJQtEJ0Rnx5aH/slX86MMtshqMruApt9
SXEMECM7/KHIBdDZqHo/OKV2at5Z8JlIGwOnyupd57omyIsSowJ7YHmcZpT0IwYW
v6ZqcuPgPcgLOtTJjMVL3TNp/+kL/dRbgSGuh9kWTJoISU06pJLDQLfZ2i4rasRz
O3l4QpCiVrFxWxpufKPl04qn8gvVaDBdCYrbRlhTwpWej55q2wubEU+khDoJ1InO
pbrJZMzNpk6HkvaI85xsZpgi4Hj4RhxmwdatutYXe762wCH9OD1mNMTN12DfRXMe
IFUHboW5TvFbOENWvqzs4eUtIvlNWUxuibWAZD39w9yerGKggvorGpeUxGk6gX48
pj0l2CYQAWwhgAxRL+D15vdviVrcAGtkkxVeMG5abT6v+OyJTG39Kf4vcT6bDqaz
p5/9i5z7ZRLCp1i6dHtHYXuw9x1yoSIlFuhEgCKlCu+MJwyyRXWPLuAG7JyEOtkU
4dCLZB4Jt3vjDPbY73LrsjgUGCEKUeDTHpa6Rvz32YJm6QITq0K+RBVAT+cTUcms
J2f3zNQCBa2hR2vFX8N7xcSum37fff7naSnymCY1KFa+ACMrJM4UZixKiva1k/3L
aJPIYltPpLnE/IR0eisJx3CQ1BV0GE0h8L4jj93rkKxzOQey2/8JOAi7yv07j4wk
iBbteHNqN4y/B0aKrmZpE+eP1yg+WUtmK7+QW11A9y1nBxu55O8E6NTSZMmAEZrW
qomB+G1RCb4dCC3umrVoX3+lcWX3ayLuTpy9Mx4VncGYYFHgg7Of1zHsT24uLGaq
8AoflnYtOHlwj6SUFBvr5yked9H6WtPYiVcdxrHCD9l7RY1mT0R9sfKVpmW5A46c
ueKeQIHJze+OpRj9o9UTag3CE6RjEozgjLcv+HiMZQDrJSgZOlhtEoy7n5eUW7jY
i3h/nIfocYOhdAqnu+ixQ+G+rbdVZBsNeDMx/oP99tqla/SsJ3dSteajFhhBMj6C
V6sL1ptGlFEcyTZ//NoJMO/kUrdUvOoSkrADq+ga/BforWUmEbKVp664A7yXM/cA
aSqtFG15UEwlj+DjTayyhzgJQD18yqRtM+ueyo2ekVx1lpRL5xfmg1FAutQd1rG0
U5gsB4F/dOqkx68gNbPmCa0BzngohJzD+sbs/yFS8Q3y0K4ffInxftD5cxIudX8s
NmqX321Jr6/kb4LIxJUaDUXVJjUVPvsTPVuvHAgF+VZZ7W476GSV0VeF3WwicvyB
zMG0Gclc9xCo1OQUdCfh/DrKl81fgt/gZdx1/guosXkl/kMJuqG1M35kumBTP+w0
SiKm1aLoURYSO98IRfcmFpy/cl29vcLdifitLwSLH46vxdtyGI36D8MTqMDjaELt
bFP3QwUb4Tktj0aa6KxfdqM5yWwRb5iPfKMgDuPgImc61WtfjcECNnetHa3JIlAG
pPrDBawnxyrflos35BOydOst4qoWtRC5LdepOg3Smzj8fCbFiuJBOlDp7ohZUrzN
TrppRSKNpzY5bqe0M+Llpp+t1vpf49h2plzT5v1+Sz7ff+7kQpSRwYHlyofffCVn
OpfbU6ZPVi7pVz8WzPsjenh84FhIdnAJ7HUG+766Dbbw+C1vpofB0WM1quM9L6gx
fuUoFZSoSsOZAt68F+GnDK0llRZaQmf7tvE0xg+CEPYlK8o60JRG7WiFoyGFqcGT
drIAJqH4T7f+V2u7M1tKYnpqbhKJ3SPW+ARA/fZB2lADA5PKCSoLX1OODCy0FG6w
BD+eGKk3xdX5WGw5AThET1Tg7JcSBi9/bu4jc87/XTuUrpyoE8Q5VclHfP6qpfwi
ArLFPVAsOwB/MsDGRcXc94KbyqxNMMLK4N5+t0geC7EMes6BJwc5TvAITN6uDC8h
77BYV14G2Q1K0AEYXw21AQL8oBgD3Zh3lxvAQwSk9nIHJZNUtI42jeS57qTtahda
ZuNIGusAHviOYbHqHkPkYaYq7arKqjO6OT6fhXFYlqTLoKb47V4INEyhVmzGvdXn
6YC662TWkTpdiFOGNhhMR9r6UmWZ4i4p4RJ19faT4renaGafJBb4cW8OREnEHRrt
qTYgucsVfDfSO6pgKAJcM28RYVOF3joPVCq8szlLQ+xCz3xmi23ekESjgsZGXRni
Ae4AbE+6WQF0Y0pbSGJED5qA6wSE8LIfL+HUdVd9IVg+YLg5escn6YKmNzlNjKBg
KyF6Pr96D7SgfBrXuvRU2PI2m6BAbP7Fv+9+i6IpTG7bAlTJcSI23MRFns1bXvGI
b7kUuo7w/yec08MobgmucZ6gS4jKyfT/dMA1pJ477jSp5JVWCLHidzFjcZIQniIy
ln0/fgtOBWaceIG4VCeLKWipQ40onxE37otEjlkhYnfvmWi3GIdR2jVrLBSPA7br
LRfSLv//PZdXFLevm/fapy2Q+F5FfedllB5IfVZhQsU0yxodcB66eVIy9usz3AXq
WO4hHdR2w2AFBiDADigU2J51fvpNEeoT1XTpq0ZztZSQiQ/rHWpe7ScNI+W/NbqM
KcyqVcrNNELB1GYQmQiQPF7zhqpSZrYouXtpKKE7qQmsjmGGipiYzeAFgWx1if+5
5l5ujNUaEM/x09oGIK1lAYPjwHiq66MUtH8uNx+VbvQcuFjhzX0BL7d5mOCHg1y1
PKHUuJL6aVwB4JtBdI46B1M+t9DkHSJ5WIsn2mw9uD2kB5iEAGODe/4k+R+/vODq
7BZof39rQ6NKn8in8NJlsjsF+Szrh+mJtIIJSXlPZ+LIFtQbPwgJdtr78zEmvzlM
2vwKy5tl4GEVhT5PWLEzmsWlfU7SzIl4yPoiyeFiK7EljQMTEbIst9jlvKJv1hlU
a26Um59NM1DxNubXjkyiqrj6V0YoC2NCF3WGVOgPE8aOJTlB6/FoDKc5PtQFrkfw
5Bp+SJ3DbptcKv4vhYkLgZDlH1v9DgNoDce5eaBBMVdoG95Mqzr+k1DqxU9aQ0A0
TD/NeI2jqcTqO0O97l38K1M6mQh2jmzHvy4epFycr1p4WpAjTC6DRc3o3MdYHNo0
razbc5gtjzHAFH5tiQSC4xRmEswMCk7PB2mRFgUj67W53GaQL7eUNygnkhx6Iyvt
/QFq77ngSnA/UyjNQ0GPaj0GnvGF/fypztCsiyedlWERqEbe+kkgpqCXcZl3aFQL
9LN4eTG+F/sGG2tJ78+LpXvzWjBK69TwrQ3BZOFzEDhANHpeL+PiDwaWZne4v8MV
ji4sRwYW5RhCCxn5slJ45gpt7ZhjZDiUnNnb4riDwtwkg7KUs82HcFGCjX2O5LDk
zrkOR1+lVs+hk/a/aXGwNvm+r3PXKsEvePTz6eaGz9rGSWWrKkkFpBNVKO0Dv90+
MnDRxir/tPraSTo4i3lgLM4qoQ42UuPb4/mUAYbbruI6Fyo0v+7BhZ0DIvFUhEQE
JnFdzsVR+Ak4o5WtNbqUGWDWpZ9QgTxrpYKJ8TkzE6gNnAzMNgvuvxlzikfPd9CQ
1ybjPnrxyhlO1n+cXJGez3ACaZOBLGYAamwn1BYqFwRCrv+5AkJkBOG0LlCRtXpC
ry0QT52c3ODLzBmCBeHyE7RdRayZFdhNjzqB57pXLAdz4BhMuLYeFAS49PHY2jQw
hecrOpbtyMpraw1SCW++iaExL2H6CPayeisT2w3tL/LFyE4IMfncH+l2WJX81E8v
3Vk5SulCZMSKO9NRRXKlrpbcTtsVnx4iWyp7G9WqpxX+aax6XjlsXu5W7ckuEjrK
PwqKg7ZkqY+e4tMaVhqPRsC/ypMEenc8mgL/aF0zusmVGbX9xyFcuWHt6kxynYdH
xL3tZchF9Bfw3OUhj0ccxatwGBQqRY6KENQfSfWMcUPpPGOqYA3Kuaac4/C/fYna
65XWLcMHm6VmCmT4QW4IbpZbG46ndEDBWMDxk4CUsUsleTj1CAYgKpJUKeGx9kth
Vwg/yOviP59M45vZAvx6sCLv4tfHercvR6WktuuO2gZoYNVfphJXq/jveNBHg+Xl
zmPP5SVhV7lIsg9o3/whZ1QAsYwElESQ999kuAuyAR90ddOywlnTjuert5U8k78V
BcyXia/l70CGdD5tZwOT/Ya9kUDIdX/5JxTVU/os4Z7+kWuaik+o8lK81p3GHxXU
K65a9s1xF5FoszwzY7dxVefBH/1sQVEwBtQxlQwwKe5pVO9/oafTFTXQ+Edi9FOB
h17ph8ThtIpxN8uVLbyLOOhT2RqmI8kIKOcL9w4v0sKqVMv2Ide2Mf+4RsW93ysg
GZfuDygNeHNReS5GV/TW6M0lp8SX61QRC716315u3vDwNj1SPnHw5h6cHGEWa0v8
lfFcd5vDb3rBEpL5FUDpU3owTo2yj6tiMZ/1vHvEGm4F2brUP7Gv8UdoPzHEMTfJ
ckt/7yPHR9IEOiNHLgCFHND5NyA1nc8WRW8FJxdIXRg8l74tmVLdXVJt7APyUJHC
3I/gKgyp1TuMHOMEiBLGI3nsnvt1kShqxPj4O235lk9+jVONf6oG/Zu8dsToyG+V
8fd7e0htrf+srUXHFmSRUCdbDBnoLVbSjI6eh7tkdm4uIl19Rf/kxHjC57aA87TV
qcTL7yp6MusJLodosvt8kYb81+u+10sYI5Eoit/OjUPxppQWFcpnpOhczhnJ3bCK
BWkpOxvRHnt7r1q0zsbZEahCdao+14l6AWe0wCG1/M2OV3+nhv6URZ6ze71z1+Tw
EU2eYZ3WHRxx8TpaIfs9O23OoQGA1OsV/WiykAzYTKRU4HX1DuvgZ09Y0C8PmL3V
UDhTvSpCFxQJed/cGL4JT4Q9+933e9dFjUgdevmQ3Gt9WS3S9oCVvW9h6kgad/0i
KIH79MwLRxMl40rI+Nr2HXWfy9uczjsCircx4Qqn/HDtDl4zeJM6jb+OXG1lkXYF
C++OcgAtZA9oVoIjJ4Emk2IHn5T5W4C0n63PP2AZiQZVillQqvwFM/zTWbWWzuZ5
swMXFFmrUyrk88dMueQTz/CRly0XfhJ6PdGoQwEO3mgaM8M208UPVnYYJ4xIhybu
qQaTLWBn9OqXuhBhbcVOUxPZq5Fyp7ZXy4b93BlFye6rLIVj31qpG49rSpxvNUTA
txHEUD6kWv4zpBAePSGXHF0LcXYFVRRWUKUGe6VHZwt/yZZdvjUmBbgYwlAAmyzE
scR6Rv/GxKZ0E1+a/ajN1oqsGL7x9SvtogrcwdC7Rlsnm+CY2pmcr/KJPWDlRNeH
04Q61rs201RL3rGYlgZ+EaCb7epAOn++Yd+bxigdxDYJ0mbKqGN3QtODKNeD2qMl
Oy+zLYXsbvwJK0Y7fw6oUMFQcXz3P6RDGDcXYPahHmufzgkd0Wdtb1Kx5EEk0SBm
QYn7C4hvshqXDws0YijkH6LbVECqfD8wPZKu7wO8beGSVKA1x+QwPXdfmEV4SFA7
ZILY1fzcr1qHNpwa5aDTHen+HyMk6kTlsDL+KA/m+LFEEqiUcUtSoW+YEs4OsMqV
I8W+MM211DEAkb1dtdmkuEPIWL7SO3dtA76D+AvtXXV2IEfOwqENYC6MjdM41Ouh
eWGlo/Bt1y49r37cPgq5RtwbEnB3m9Wmz4IH+6fyA97ibRkVeUR5Hzb30NLejl+q
d7aZB0hMExD+th3aiXPAT+Y/php/YXiGdiQYJd+B4ck3E/NqbhqhKd5amjdxvfYz
dGuaUl8RxTI/RiUnsfnPSJzyC+pJHTw0NMkgjiFwTJbZ6Nw5Rlnve4Mdt1QqmjU6
uuwPQN9Kg6JalrxbBImdY8yIQh2Cf3Ek5Sa1Y/TZMr3hiLGDavNCEZUpjyE9SnwN
4pYwrIoH7YEMjkPG1xuqpznlnFECp2VsO/xQ6CIshQMuBwFIhukltOMsjJbSIJGg
s2MUyhkdG95UXSc6tDoRTU6QsyuxmisQHy6kE0z6xzlxqM1wnUF103VAxBqMoLl/
czdGAJUbyFmMAPbQiFsWolwX1t7cEPro4yRvUaENryh9v79qSJ7RHT9Q0mxr3KbW
xE62rHwhmQBHxl0KgYh15CFpmEJY1kJnDwLwBctAwPh5q4vyubdzTCOUhcwExwtg
Me8kGHctMfqtu57Q0uqElZqdjO8K6flhs+0OqiiZ/Gz5J2oGuNs4O31cLurHpCn/
HsmQtKPjqnHifvOVbsYMqytFNFePDkJQ/n8oCKPuULjdeeg1R8n0MvzcTQ0YO4tV
jdIyDST3LJ4i0biPxByUgQg2YKXSIYGEPLZK8hRfnDdhwPDFk99UteN+ca43e7ZP
5bPsxzLo5VvgZID638KVp0XQq2K7xYA+TY8t+qnP5bei/KEULZsmF1jirgiDCD7y
UeUZzyJae86hkzPW08qIkLiTXKum/YOD67shTyVjqmPBtdg46+k3lFl/F9sFdK3N
tJ84G3CN1CAeZd6PjySzqUoZTOnpr7MbuH2rqKTQgJOHjRPIacAG4B++Tdo4ksMS
GoewBz4Ph8AIARtOCP2zUFdjap92S18aka/T3hKphqEZ1Gag5Ec4yb5+wEiR8H8b
v3Mep/8Y6hfIjiBJj6llFli5UHQYSyu30hkvr+KLO8RXJZCx6FoGWLxZU0omZMw1
/h/EaBn1DZkPuT0KaAJ6GcuHSTnmCpfvEa6lHOgXk7eGRfoizn7v5wpN+DOjoz2l
YaLVctMmbautTFd99pDFBZkMJT98mnjY8BiWeB869RJkrGJXD2UoA6XqjbrXb5Md
sJsX2v2Kzog0jkHeI9VuQ5e31VcsAQl1s8uxK/Pudjh0/CMQWbm3BfA1VuB6mzhm
n3dkfMWoRwIyHbXCxfcrVbJooky8aGF8hfzHaJWKcudEfb+1Ba9S9yFgyTKBVslj
G/wAp/ZxlrnKF+U3XBToVhmssHW6IcUgIf3mlTQCkcJge3q84hp1CKSOJ10TymkT
oP4gKHjhVxxO05u7eSQuPkzkOoDLRFh5WQ8FT4P04rjMC97CYAbr13sHM4lu/8MF
w+0jbAlU+hkqwYvQlBPLgR4xdG3YFFvLacdL2JVEZPhYZttV4Bgxspq5LZKA/LXu
hlFIc0v79g/TvsihtOzFpj53FFTgxweag5Bn4JR7X/d1d0CqhPHq3ZNID6syrekc
65YQ06fbeNQuxHQeuk0D+Q8aMW/hT1Kq7sbOY/o3YWBbw0YFap5TGbij4rYCrpxI
4HRPmCj4H86Ks2DZ4QaKkCFjOpGE02HiDy7M8H5NH99vQwqHB9C1wiiNifZPzM3a
CTa6iKjOlLsUoFmDta90FknpaKAt0E2Ku8ScRbFQBDOr9EJAIWR6b04dk+oQxrq1
RcNPBhUaQb7fyh1ytm7uGnCLRLnXpfPAOGJE+l1jAgZdcdghRqQI8UDDsTLs3BaO
uP1RyiidqtvJcGLR7yBAUDcoURzY9pYAjs8IiWu9VdgQj5jTM1YeltbK2Y+N5Pnb
zW+zHHmEcxWJzIWhKd5Wov/fgL4hEncu5mHX+HKFQ6XqqH37N7y9qzX/frHzhN52
jmMpFH/cp1aDpgWCODYXgnEkFb+lEtGfzU8UJzizDkm1f5f6WY9CBh9HXcXDJTbn
ZtBeAudpKcYhRycT+kIp2/dr/0rLJrjxvP69tYQucjqq/LiJErrmzsiKDgg09KG7
xDOBKpzdwwMerMF+gAkMzNzpqE2qeWwAITzfS2qe5TXXRRrSU1lFaYRE07k5n4W+
bCOSGF9u3PR7oTV44R7VtSXYqMMpculletIoRSMfVrslj41j2dMODb8VEQ410Epb
bc0dVGSkD09wczZuZAW7LGwdEIjFdEQRjdHsfcVDgrwEQspiizoSKIUdSCQeAJwQ
yEfNYKXQZhqsXTdqOULUV6eIgJvJ1yPVx1wZEi+C4aU9rNw03H3WqbT1Qvf46TRS
Fk8Q3DlCUnrhL0nA1wpw5Oq0p/1/OnFPuoEX5cP9QIe3cg9tjxpGLv4hQ9UpvGj/
p49CPgo/Fbyim0SIuCxzG/GSyjoDg4Cz88SkQUfWGQjxv68AFNqGidElqmvng+rd
VXBRiyBewIbocnFQ3qmq05nWvzu6oX3fmb8z1kR7mSXa2j5pOPgsw+KbXhukqYgm
ssp1jIyjEJ4WFsFVnSAfy8ORshng8/z855H7AGzNjfAm7ELEfI91dFbk5vlQbdgD
fELiwaV0NhuV/66tLiMdr3kywhPW9yVqLA1c6F2wBXjogeR+oPi9QbPSyxipBGpg
Diq+DHiBsZ5pPBZ7cG5naUXRluzvVUZx3Ey6IOyLObH1lsGXW8SwozfAMXDQjJks
MvK6NzjuX0h9BHE8mHFcm8mP6fT8pyStVc/ndq9/bEKCTsfiXKE7ivvjJujTkqm3
Rplp00h4QVQr71VlxgScT013AoOr2YYLpj2cy30aTe9AL+uicbIsPj28zr/ylae4
j4bxNeHXS6CpZ0JTLBm9+t7gOiG9kI1v4VkIPbrBE0PRoBiPUzkan8LxFUHcifIu
v6ejWOY2dSlHgiF5QcK35wMVLbf50+GaN0jaf+Cq5cR8Wk76yzj8KsQ7rWvUoQvt
wr7Hb/jmL8fSXjfe1Be/Uf5K9L7BFMfw87dTpsnrlIrqxsW4r3Vrg5aZlPi48NZe
uasRquG9ZB+h5LZfhoFED8jcZdLMN+Auqq7vf2Mtjnc2uaTqZJPW76wzz1hZzSVj
t2VwLdrXy40JzgzLdg/8L3W+Xx5gnpEj2JNNg7J0RvbFJ3vECCj3oxUdcW49y2Cd
u0LaP0BKjAvJQfmyMIeL5LNC+ThIVC98heJGCC8Kqk2VUiiZ6BUHXnzo/cIoLgnP
C1zUBvvAqMvICdIika9vTbUn/H0OA7TyiF8Gq2a/Z4Xh+8JqyGaApQ7dIL8RwfhY
iKh1jM0Ue7+VFH1AoPgYPWC2+bo6XCHRlL7SEo0Wz7RrwSRnrZ4fiAOdhTRj/AsQ
uOsScKd3cx3CkBAY+zD4rhq2eqyisevxNwtjL7fhnEJ8fnOgKUA4nrCg6A9RP4Rb
cpONVjV9/WaR8KswBV6UfaoUzqlFGHFNyENKaY7RqnvJf+FFUkdVt9zDuUDr3eDt
CAzSZi4Ekpkz6VDbbO2hwsOkO0uC5aQ+wxJ/0Tt8YMg=
`pragma protect end_protected
