// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tXr0LzOoUUGBPasILquE4FsKR/hH2dfnPu7rDGImlX08FIbTp4ChSDu1s1JrV1lx
KQr6TF/yFCu6EjkfuKxxRjI+5GXOU1bRBZbCayAa30COEcXttOOLlFP5CQm222gz
pvg+jlv4ZiI+E5uKb0d9NuNhkoNLfkBc7q27w89F6UQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2720)
Sc9u5Dxxz053O6ryWIrUAn0MTRsijR8xnnj7UFPEqPS57tANNfFob2rdf2OmK5mz
oLA3xSGkksCLg7mXuwto5HdAIQ/zCQpl67dn307I5uNEjJTvuK/V6au7roHa/uN8
gR26LX1gkBUDS3O79/tzrmnLSnhbpa5Mma7rB6ZPGHiKG0zD6UZfvzOgZG+ij232
kZNStxbksDFhGrJEaygIPrY6CeMRYU0MifA+DnClrNo3mIdpKSvIeOwcYpqOX1e4
zgGL569+RyH312j5GuMRKpIlBeOJNAQMAqAX408Lw48aN5QOsp+8HfTBXRiT5PwR
Nl16fwcRF6abck5/V1zZILYS7BzK4XxCS4vELW31Afi4tdZo+wqBYOVzNiUcyzkk
LYEt6ZPSw3QHMhrJPbVAAMfbTFWjzLxO/RS3pGqvcSMNMx9Rz2ZDeopycuBCNuc/
68NzJVLSe6OHxQ+lx6kgOK6j6V+/hyOxiW0oHYxOVeEhuU1DfGECS4B7s5GB6sF6
cpH2+XqImnq3sDGsFo6GMW2dc9mZmI+NcQiJ+sEl+0XbOE3VtGuX+KhCVQEhWQKC
WFTlWBRfV9+7CYOFO0bPDJcV0BUiwFq607Rc1jFxIWODsK7y08uemMkjSWHk+8o1
imVE9+wevF4NooGPFEeD5SBwR9R/IncHs60Q8nuD8FAHczwgiVXwARODEohJxyvS
EOlVY39gWo3ZdUNso5Tw7obR4MzMk4lJUQp7i1/ndGrX3y2Ba9Yu4Gzxz6qEL0JV
+ryc5HUCEnl1FfpskG0au5cl3ZEBbgG2aa920tCFAtxD5V/3aDPkY3TLu8tOIQl7
EBfD+mNlQ8IMTcSX/tuxvGdruuy/969KFGKJmIwLzEixWPJHxBACWpVWWpY/NZ1Y
dnRCXtSIQiFZURbejWgb1uzLoptiFBelnSv7nrzsLgG/CeeveW1WxFRz9dfp0X0r
QcqaQCwuzbh5nxxVeRF6qTI4gN3MSaPiIVTjKzAXW33Q/CajDYEKE4+vnTLIuFLR
hzqH+jgg2GNYnuAW4QnO9Y1pqdLCGESGhehLZLoKzPLgQ053hQ67TKSImUsttq4H
cq4CVx6/W1hXjg/2nmb/RRdPpqpF9ZjjjdUrcE6DAo8eW/wspsYvSCp/dXH1vBNF
wx8JxKkH25zbc44dxs/7Zx4F6idWEoS1wrF92j86NCxC0fQodKwPiFrjOc2mNDhR
T7DN6epDrftgExCcn2n5hA9mEtWRNk01Aq9XSFPFZmpbXIGFl7iULZbnOvql8sAF
6fMYo+RBAdbD6XPC37Woq2Obcjkqayta9HA1WnBCvQYDtKy40PM36s9s++/EAEl5
mtK6/dbL3YX/n80VM3mtp7Ps/9czbJOateusaVf7YmIkujeK8aErOV32Le1Jfzvg
zF978VkuRejjH1MAOfIyS+u+LsaMXGJuGovjbI11YEiu6fr8n3MN4aOHwDD6xBJk
9e4PwcShOxi9egeQxe47YMln6Nv+QAneCvln+S+S6uFPuTQSZrJccpUtP6ELyf7L
lwn/mcUUKYCpSEEo//QVFuavi254Q/sqp/aoLbsXbhm030j3P0rQjm4lloez8jya
qr1YRRieG4QD2Ugmd+Sf4l61J0lcmgikLAOlsSfbFPs2DnArr7adfpYRrGhnwI7s
XAFRVfoV1GPO/du3uq7LA6ptHN+lsHbZzc3PnVnerrEgKYp6eiuj86vvH1WWPO0w
o38gDz+iSC759CEN5vJpTvHE//1IyK4mYP8sxOZarbQ/PDNpNDQGmUtYqPcCTFBa
+e+y7GjUvl/7WUd+IRTnZHXtgVzZvXmIj8fnODrkVlNt/at3glxGU1KvZtha/lyn
UjxqTb5/iJPG6bfOanlvvfbULy2Yg5sVZAcS6FsyvIkAF3n/V2Qp7TJd+rRMFwQq
tPny3d1YwBeAU35QjCZ6LLz9iVUOpiJw+68RR65f69XxjxyYodp3SXoPEsZHWAuT
783FdGdOcpmvXfMlNdwg+Ji+U2zbTAEJQS7CeoQ7pGDrTAIFm9AyzQxYABkwUfdu
/m3hrhgCPWgFMvtMMCB4d/WuQ8TOyp9+jp6Za0jraiwwJGsrw2MQqP7G6eJdlMEW
mIhwYHKUuZJanxxr2QbCmbOCqRLfqm+CiCSOCOrySVBrHzbXTeLWo1KUOxacEf2Z
btNdQiMk1Uuz6+SWGfI1Nn1hIFP5+scm5QvYWpzulxKvk2EjDArW/Xw38Bwaj5mw
mWyLhS7xfJjPQ47fRVQ1U8R0c1/pYy7BrmVHMcV45RjWmNA4U6cfdlPy+KZxvAj8
th2pcO6hs1b2/GoBysZKg1fhsW/8UfJGm1HQWgwlYkPHejaduYzZpalG8mgYlDMX
aHfKNVzky5DrvTnw4nKylmaAUTH+CeLEenPedsPlbjBY0/krbCHIFtpb10AQU0vc
g8aKnls/r1c+yqfbq5l5PLQnxHzSi39mJzXhMcidKpoDu3gvZTsvgyH71HzN889o
egxGrCFkAcSLBklai3ngTCgpv9Hji7Qy3ojRzTF4djdgBBRNmXTwqhi7FmoxcAjh
uFVy10O91Z0vzvxJnsGZ5v6kM2k08FFgb1tWlm44fltwpHlDAvkno7b/eEFO1ukt
x1AdHv92c+TOeKgyaAEeihF6mi0BQC3DHSAsipqR7usrim8o1kqiNMRERGzGpKuJ
Tf/0tCD0ccOTJ3ijMyQXmKugoLTPpnWuNUImite3a5tp3zuddYdeMo9iq3PHSYu3
nJQ1iodJ1nMiRPh6wailcten4bFI3RX6UHhOXbEKdg1GmbjkZO6APe1vIZfVRgbt
r4woorIF6MCHAIpHxWRfZYTBJfqw1nOjwLYqqJh+DyGDIhbO0r0EfAXZo0cYaLON
I2KX+qns9SJYufGDnrDzsV+QRC8myRja+l3BykCnJ8KmaEDy2dTCXbZxkXEpJFHh
+dW0eP0dm/DXhMbpibxK+SBeIySeSrNexNaSJUWcQaQSuSwyBI4wJLCLGnXybFmE
GADCYIEAaZpswv3ChyImcsH+9fkoBT6o1Xayg2wMRfkBvm7l33o7gGk8KZ8utFyr
u74pkW1k2Ryn0ANbG791QMB0SKVb0OCJFF4SKhpr7TITTNLb0brGZliouJXt8B6j
KyVyBWpAO9aHa8SsNpr1jQw66krzkH4KB3ZKRaN0wU6dpiuVw30WEqIPirJBCmHm
0+zlGRWmNnZiPqUI1NP3uAjOUUy7iM8fN688HX6FTX87GoEr90LLQIqetEnQAHsz
XoEnMtEW+rIan9SrbE3JOoGJ7hC9tv0Lh5NDfQlnI3lctDWdVIAdHhcXIRjSkBbM
eOT4m8ccy0cTNBAc4E4fMLvKciprGRQvCTTV3lVXTvFPQliZy75BBIYYrABoQq30
ynysqZ0zuXKvecFAwxplOkavcoDe1J9TkY4C6usDW90go2vaNBgxmjI1DYjWD8Ee
h9k8DYvn3s1M92/27kdPoNI/ekyD5XCgjGkOKqjXcNff01824SwExGACI0noXOCX
ygi3uBGzeFK1e2DxUpnLUfGJnr8aSFmFWxYMJLq5e5N5tD8TiCK0XnIT0ArNusD0
wPuaWaGnnpGuvM6V5wOED1YlzqnvFEwmt4mGXpi1TH4=
`pragma protect end_protected
