// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:24 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
b8nuLtj9v4PhzYTQIVVYSX8/0Poe0P9Gv+j+Nxz+JgGyaxWzRJJSMgB281/tgZw8
vfkqrbLb+ztkrFg+AcWuAmMAcRltvtTREALKMnKzeOCs5hXV4pthA1P+KAYOXPvK
aW7uhiFNfP8DLkhJnZVZNFgpDl5n2j60QYlA42bOTUQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6880)
4Vk1NcD6tEQ5BSOFOahbatryMJfIjKhwSsrRQTHwbLN8bKb9RxcpYp/+EVsUyFUg
ReUP0FXxeLWODZ0PCKLBoXYhsO9585z+21FR9Wq7fqcgNXrUhcfJTLg7CR9JXWwS
TVec9cnttVAIOfvLr2OPH620ALgMRUl6ONCFVnmZAgvRngVQ2DLiGHMD4N23QZxI
fI85HWKX9pSuHnIt1mRMreJ74oEnyBrUsZz9BDOm8oAv0HEItapeIymSsTvfkwzN
RufXr+a+B2RxGprX2BIykcSw3uTmGzAQO1t7dlFy6Dfi35harBxVcSzuKEhzosIx
nTUwsbKhMD4kLmzSP/sngfXeEOPcBu8hlbn63QCnQvC99SKukUlayd5JYauBtHF2
hbwxL+R5oFzfcpXj9R67Tpv43VC7m12USDPq/UoCPEvye3s8Mm8tJPdLGoWazI4I
BT6F8mf+o6ZjZhp1U+cqgoHsg+kU1WLIXTSbsKcRr2tQlPZRR2gRUxUN4xOQRR2v
ahlFCxkABbpQpL7QlnIrR8+0Nd6utz9FO7i0Fo8gT+2rpj4esvPF4r5gyfv+xDPZ
sh7JSDACfQ8xfOVQdj5ofnE9JzCF3b9euRFH7aM6d7KX4pRiN+dxKGQudGg2rWx1
PPvTadSqA5J7TRaW21YgLpgIrd7cbiZRWS86IwbL7Qr1P71H4vE8FKYzCTYyIuBZ
1cfY/thGHhb1GKdFiuPlfmBtoRhN0Jcd5Mp7+3aMcZ7pi4vACDX3n1F2ROazwtwv
VKyK/ne0HNf2oHGxDM/egHbkH1UdqC2EXQ2cAZZRAfFL3ucq+nm15QnsYfDOAtmP
Nch19Fa2sOhV1aT+fkcBGB63n8hNWDduAD2abtobvZzCy3OCLULAn1d/9BVC8N3E
helU/zlcFYMMf5qIkQa2ehfi6TCTmQCk/fYfC1lCco1V/b4rCIQyaGxRomGhy/HD
xWdf0GvYJYPxmfzxZ+UOs27I1uADGbziTulPLRBTVPK5bYmYtNaHLo/98L2pGWML
lUFTXXMsasB94SBBLgcoGRZNpJBmJ/IH38icViqq88rjG/qKal1CKUgRUuEjwApN
Fhr8p5j/DGfSG8NyDL7j9/iY2B7Zqx7EEMiOb3AXAMvzcD5k4E3JQofPItZ9KCWg
Q03aq+xFNajQxzU+VmX5st8PsSlDFoF4hw93NxU6CCJjrGjYUXq8iP/L2w5CwwtF
8BWJD5Wf9o3vbPlRsIpF1mw7dix66yUMkdUw/xAwDvw/6pdjBfBtKQPaXs4NhhxU
ek4p6uIWZP70URyZEjBTLzQmRB8/EUzERzFFLHHkiDBE3T/P/PB/0NORtCYTSeNq
vD9oOmR1M2dBs2SFi2g3P56OtU9QgAFKcP5uvffRz2ZdRq9JkmkVMZjmCDBo+xGq
h0wSFPrycLCoZpvCmwHgQTJ68rauvWJmT3Yk4ZBxS5cBkF3e3ljQd3znxGGnkNNI
Ow9tluwdRnV70oIpWjAqcUGOVCpq9eRG6Y3lREM9D4ylLPmj75sXfzxX0KG48rFH
LEKdHHs54Q8cdlVFkL8sGrwPIOLuz1OqEdofWEXx5IwLAxBZN1OgLE2WpCBCGf4Q
ATHKgOw+V2BIGe97P96tIa6pfWJfx2+IyVZUxmk5cba82iM1yrJmKYZqjG7MI+b2
+SwPkU+SukHLKr+XNU0tFWYDhqJvVoYwzd3fst4hymiuP/JVY67jtbCNb6F2MdsZ
6AKI/HRHGTX1rjoLRD8MCVHE6ZO40812io702AwwdjOX8SfdqeuiycIRDrnHJLee
qm3+2Xfr2ihHUS/8Nx2IR6wCv17XRkibYFCOnqye7whAiVDADFy32uy5c3cp+F3k
oIusHx2w6XI0arMWDGaYkHBDnPCCBGS6nnIZthJK7Vw7ONAfgrlsQUR1WRJRRJNa
EHKUAxsd2isJwikfJF9/Fs5ZXA2NbFyz+9MY2e16/IUxwOCYXEnCsQomFCaM3e40
98l4p5z/ARvP9a9ySUTHOEcnPUETeEmoiTJHVPno6Kr3X6rRINZab5jcM5QHHeLw
H4q8U63YR1h7fIyqoMEzTE1ucmGJhQ7MhJKfa/jDLzkpZVvfRRUK99BsjmAtfj4j
f1o/b/g5RqYZDvkXICl1jAWuVkWoSlgh1jeZqN5bi0gvU+aAwdeK40kBR9CgAoW5
0x/HhC83CK6N4dKWhbW2ebzZEEsSa67dzB3SNmrESBWOSaCE01Z9YeCtwx0uI0Sv
jifcPpaP++dR4LA216YhYYWJvtn5dp9CjsYZtLqlAorPRoLaCNQithkXVxJAL/1D
Qf/p6kuWgT2CWdZAb/B2qsw0cSCIDzIhxNQ9a3C1CAmHvCWi3JhbvIIsfvTDJ9vP
p0p8zhJmY6+lyWFJ5VVMfih2RNTmb7jcub6PMnTpuW5Dm+cKUWRFwoLUyvHv+dZy
dOZO1llREt8akJevpL/Moe7dkfZBgJn8fU5ufh95a5t5EerWmfSF9K7O23SYIZBZ
h03NULnh8TBez2xJSKk4SDfyP9NgH1ra8/Hb4F1wqQeLd2nONOkJn8gOcJ3OGcew
V+AzYeH18ufWVJLCJXZo2IeFblQB4KdIK7xNx0sIsmAgam08PHhd4C3NYBMDyZ+j
J6/k+ssYKiD07N/1qjCx8i7XjCMQVkXU6r6mgCws2UFcSC+t1y7oCmhuiBhKO7/h
Vy6l3W0z7qHHZnjZwRe/p89WxnjPIeUQdIwII5x+HLQQJomIUgeEsm/J2j6tGSsd
CELE9tZOsog20Z+T3sKN/zez9RSt3bdVxa6yqwOla3YGpGy8GHUdC9QTDCGAlL4c
aSmy/DlAYAzXrxoOMbRIF4Hj1GRFE4ZgjpZtQtlt2lIVVwRx0EgVpASH1tiunH9J
lVNdrPF3Tq+2qC8s1UkfQl/qGYg1IGClXOmgGVtpYNTvQakmSv6XXR5eNaF9vbUZ
jomdPpOwrTJME3p5ZU+ttwkae+wQRNXJ6BZvaQK3iGWWNA4D4DJx+vvzqLGKoLIM
VMPiuSidUPDloAz/iDHNDopAK42P1UU+cilMj0Ug1rn30gUnf13o6JlaOWqpq/9y
TY+SWfJTrWPZbmPqdmPkofAgnK9uAaSQAdJ/OUhTJzwyXMoW64cGIoAG5ilDTAKq
eEfto3NypYH1u47U+Q6I1YADuFi3GpoPQU9zwLegqttTf6grRo1TV5Rlszi0kgmu
MCLN1gxsCsLYMirEhKhLYUbDifSUPbRyv4I83vItpsBnRyqLA5AuXWRTwYLaOoAK
Zrx6mlmTguXZkOOU6MlrTVB6m5wK4xJL/xKrj+BNDhSBqYp165k8/Sf2Ae+iOp/G
BzvC0Nk5ui5sDgUorhCl2xRnQxjL1pfIc8gOe8SBCu0kSp/NkwbKuaiIdq5V6B1k
DnFrFUxNPVfk/oBIbkRM+Aq67HT2ORprk+iS1BIM4tX4etBY4jilpONwb/vOR3H9
wl3iH4SehUko/fQ085fA1Uig88Vgi/CzHQR5kkC2uPPFS5Awtj8XfZZnTsKUoBq6
yNnZmFX2o+/epicZ6CwJj0oza79fC0acF4lhM8Qnn+SE0/B8L8J79x30ArT/3g6J
HUJKC1LcomWUKPV09LYOyif0X23Dop6AHEznG+Z8hBWWx19bhoFm9NxV/OTMZy9j
ugo3UwKRGgOkEciXx5OGTFiSqMjoFzqqwKUM4X6kcQBXDmtZFaxXMr/Z9RpKsO6s
hqIsHAnuT93tOtoWxM/GHtzaxGrFUmhqz/7t99o5mdgC69Hq6Oq7SREbH1X5TBR9
Xr0Pkquow0jtJcjaeoG9y1THVXmZchY1IoZHXGvMJr6Qrf7x5jJbQC+evb9b5nUA
FWnxprCoVWjlVO8xwC7R/jcOS9I77xvatt5DSCglu4XBDWP0GRb79kWdM8RZ/3Q1
6LteKatIa27VwM0hmpCxlteoTsVjs3rGF55SmknkTYyGNdNhPZHzgaOgzSXWRSyu
O+gpf5Glei6awlKL/wrd8LKtL+1HFjUSMSxRk7sHrPI+XuVBu/QBcEKMGPWH/S88
k0FSXmi3dGUaWrNxWfj1ERemPqJny04cA/Ite7TUhjJG9Fc5vEg0hGEfCf3MuZrx
kh+sQB/CAzksTQBWos964cFvus3dXHKeaqkXPqjj+vLVazzuf1rQGH1OX2+sQPHJ
h1qeqsgrFTy5PAb26WgTpINxNx61rfgV1cMo9zdhkKAt8GEROc+aRKjr781kH09M
pjQ2cBfQNeCkPvcSw1PxGhtD6CsEVKd2h97cA3VuPtUipc7/iqB/m8RyWSxAbtKy
Cjf6E/SL6z3RUDPDeVtakJN8MbKLIv0B2SyN4dtbtABzGXfZoW2e+8Tfv4VaMZsk
T1PBwMjFkCrIeIle483ukAqdI0dkdUCXP2C0ZHsEldbc8bZM0Ws+4rTOcmc3Fbbo
3xQV3WaPezON30nK9pk1XzM+vDb4ktYrJq93ufBDF34FOB03lXwSCyVTlqTgO3e3
asNNtDmxhEi6adTKhU5dyq4GazCgiureLGn8KoaOKI82GT0MC5ysARzlvYMDukdd
jMO1zuO2xETIz99tQQI063dBKrs2fF7m4IHKvml3nSjhZi9hQTIjG01INhhBsVlU
HX5xadEMrDuUXjd61jZ/8BcLWfy5amCEBGRS0g3+cprXxfqkpT95K2Zx6H0czj7g
gT/+FJj94qnpEzck4QqigHx1KmzGaEbYpl4h3TF/UPi63oAOkZBkiihW/tEqEz7P
doHnQVHr2qzypDVEFn4B06AjysNPQpF1xFfxg2jzN9svnqRZBN1gn01sotBi5pPJ
6W0Yo86CTsrvhb7ZXZZod+pz2gENRl/CRfH1p3RtnqDyH6QLbwIfk3J0a65lZk8K
t0ojoj27/lw00aWJWCYKPlnZhlwGe940K/g+JyfXw9Pi66PklV5NGcASyInJ21Y1
KS//KWZm9dVc4XO/m+k9HfuynhGsBCpbWc5hrQKIXNsxf+XWg1HJ1jaVX6aLCDOq
fskx86dJaki+2Tq7dSszUnL1jTdlOoZnzh5pHlx2zlEfK274iX27ILplmhlCzEsk
JjKjlaakcWfVO0Tu9KFrgIC4GfMOTzrTMAFSh8JdV3gjWdo9/TcwERh5BpaO4deS
vieIA2vMCiihiiCsxb0kpdWDYQkQnzlSGqZqHMqHEgTaFiizrGD9s50acKfmXLaG
jI9QQ2A3lVrl5ffy0SNqIMQjr2LDWNc7kr66t1qrGdrPvAqD6SiW9HSptAYkTTLG
/v0xV+hXkqaSolEj5o+jDYEyz42KkB6SydmhkVPJu7D5PiJejCoDQq9IHVQHu51t
p+598QB6Sc9hzSdYVgvXgIjaqTqHAe2pfFmt8S72gShBxG3ubiFislHtx3c1+Iuf
Zkdl2VzavEhhCSahtd8i8xYyJbeKWKfIp6jL+btViV7wRqohW6huDxP9vUpO2MmD
KSOo5W+OwxPMjGjqnlYmPyzYXV/Ewn83baK/1SxjAbJHFyZZnMyix2asVbMkqdn9
AyAcTit8DXth5KhtFFyK8Cq4ghQxciymgZc6giuXI5TGlySRNDyujQIDxqj31cm9
rzjCLFcfZJCifwoPP7HH1KxG9+Fdr3uol3UAveB4gMPwiDzDY9D0fQuZbG+QTFn9
Hmr60uqyQ/WWIY4cI1U4Kc1fBzINUkujLwpMvtxB5De/JnNfm2EopzU0bvc7EGTG
8jtJfyroyPHI3UyNK12hgVgR7yuKUY29KVJ6DZxhGmTbLYqHNef0HT6TajCKg2yn
STfrIz5k2HcqGzZ9IAwWgI02mQ6TU+CiAgDq1gSn0+OpHh5WnhPLPYvOvmrWSrj9
bO2ZOje1RBJP5EEZ+p+eWzMgMXvLGxOnlY2pwwGB0navzCqNfsYxXp/oFp7QrNqn
/x6Vz8mDJLupTQvPAbBF8iI3LSMQ3FlETGoMpOJnWUvcAUf/GSev9AkTQAEVoQZ2
zHcII+lSxPfSXE+W9JJuDM9Bgby7Jp+Pp91xtwKZ9YQrEWW0I5ciMwN7ScIY4rWs
IwkRrBgrP0+BebWuIQJFdiJROdtGdmTh05ugsR7/KGnZVvoUTPC6lnUcEJFQCA4k
pDilMBKSprpbkNQ/Bwok8qInBNUudteM5/mzr1e1Nps8BjhBBX72nF/7jI1ADWNI
eHcvb0iM8iqMXVY6xAPefdP/m9q5iiFPb/uTGwn+Q3QoCkNXkGR6YmyAu8shg6k9
J1eP32SOX0TcINCZdpr6J9+wkhu3T4X7NhCXtk4ZH01PlhGBobsjpYewPbjA6UED
q52skI4i6UyPvRiKX2+b6oXN29FEoNHA2TGxs2d/9nD3dGaEUE8lSoRlistrfr1+
Vg7qm9P4HoBAVloRlCA+DK8HQ1QQuWlrvwwR/JMp+UVdWNsPEvhKg5qonQ38ubkj
2wq1B5R9X9i657mmgeT3Gbwdn/LbznJqcOm/KpRM2sxnmmzDTZz+lOXwXdh2R7FR
PevUf8lF92WyjqJCGhvdAkIX3gitAxuOkSB7OKlqdGmwy9lUAwZoNXIhc3j8sd05
9vbM0LlgDqp3+HyGbFhix3VfeK/m+SUwL3I5bLJHo17wTV5/fq/t2qRsBhUDRPGm
5zbqKtjdOQDUmOq+fp38KOlD2nyAMG+UThmynzzjNmNVqYIp21g19TaL55Uc8ORc
feM9kqJfCYRImyaRDultdSepNXVGEP2VJhAXjGVtSXIo9RS6Dhfaxx2KqTtutzSR
drQqUs2miyqbT5BfT6C66xlpSpesYBdztdwr2J6roVj338qO9y9IR78JpXs0C5vu
xMtjGJGrnOF25d/9srBiZ9EjcqOj8tv8Etx1a5LKalmYuv6qtJebp91lA3sqIyL/
V9dxoDIQgHmbXvsVd7MX6Q0GpAdKda2C37flFrIt6swHPEv9IoZegEDyKswK6gBN
pyyCig815eJMK20+AZoe7SzKskGEmu7l8po3W9kT7vceMjiVDLsuqnmuVTvBHh5S
7XIfI3MlZqKjZGqUT0F6FprvN5fAo8Aom6a9wGUAeiowQXSZHaHlrVLLwYH3GKFo
DimWMxg8Vd+EWtFQlvtjlLTbS//XaVUQbzRVxhNtAsrB+zO0V/tJ7llVHntEyRKY
/h0eN9GjWRQDMLJQ9WpFjaYzu27vo/kY1EUXVvmE1WOJ3ziP8Je9To2/vrUHjicp
9/1NcYRBfx2ZCJxnbrkaP9d1faylaUpiwxFJu/akLJbxWxPozohlVMsm+FiffDI5
2ftpfITChRHukd65GjZYHwKL+dNDF8q/SpmhnRcEfylCIwOHJFa4mdep1NxTt7AX
atxQcXlasXku9RiC+j1dg9srPvWUydGm+J7RUfKaoiA23+Ms5Ym03fTEJ5HqnQbC
CRXyeHnLTg6W9ViO3KCdcNo+eF1JYMj/IKGK/6UrJgr6liB4aXtisZbPVnBhjt42
8JZsrH6PkQ6c9XVoKR9H3KPD2R2tr4qTAUKvHuZ+Mg7r6KhNfVXg1K32eRmh35GQ
9+zNxamPExPIhbnDmLfhQgagiS+xAgK30SlpQRUpvwQJuFnUGcn8v9qx3Ui1MJD1
kalj4v9dU2ces9qrHhlP6d5zZeAaEuNRPRl/Y2lqwmiViz12Iu47S1krYLa48VfU
zt5f22ySvQj0jr2DQViOPB2oJGug2bdAnqbe8gT+wohhJ+d3CnpG2+S6VkRI+0TY
o5BUftA0cEd07wzXrZ9Dc5RNMz8Y0v2vcjHlA+SSqg/1Ab8UBHBaVDr5Vh0duFfU
C10h8re+54sHO/WpYcf6zmlFrJxbfjeEYKQ83sgT+Rl7rYwY+FriSbc7QJt08TsT
Dpeq3j7pKHtVxx2jDXuLoYULAYrBSQ6iCTB/k4hxWjQElpa7j7XYaaML7pL/q1wR
F+pK00M5yD1Kkz7DzRRrEHpMI+dcqsWXg9Y9b6bHzt47DYXLrIh2B6dOOnznzE8P
RPzuq+krKikwGvoznOWlxUk20UliEZwRR2MQ1t3dfZ3TwaDr8wkBSvueKPQlpDYX
yPLAya6okVtIgzck89iZX7vk3dOEne9f/SrD+32eAAml9U4fJtGXe/DRh65H7+iZ
geANeKC5rn7U4PMjdetoI49ciLZl0BuY7JULy568zeoP51XzKR6QAVtACp56UiGm
9uAcMAtc1/JlrG/D6OS8w9wMeQ4c0o0pm4A1awGv6EjPymRFXIQJFGoL63Qqd1a3
G34Kl+LAi+MtU6F3+g53cVfhPhjTx+Zy276pvzzukHea73+BnD0pAundXepZ/skN
CfkTarimJbf6/M03wAt6ULK8wBmmYh5I19q/ANb2R34fJnYOoQp9l4n1JibCOpE3
A15S+stoy8kEivdm4TfTUqLMiwnksbjiVTUw4BhxcmjCzvBaYt6l/852BEtJLtQT
Wb2w1YeIVE50NMYZARi924F+ice6zwsHIh4jmYRK14zhLLxEjNHnfesTmo82Gv3w
q4q9fuoy/OS3DaiGkXtVWAHDmUjsjCwfEcCwoBHzAysj0EkGisUElUuXNzAATWKs
pGzudLiXiCEAJ8qRI11W9ccoobfE4PDTgJMV9ME46DOzbRGvnHvI+DAu6jd3er4N
kO1kmKqwScuG14i7zvHnN7FyKIGyqHJYn6X/K3Cy4K+glBzn53RlpwXeGQI+58gh
fySUI79MpLR09xxGvtGznPPqUTbTE/MXPwPRpIomrGqL+V75QA2OuFbebFKjuFqm
xooRdlHq9eVwDIPiZtCuPsDoSsKDrNNc89iTP3Wv6iqh5fsP0sFcwhrEOqNbOCtT
6LlQDXfrfOhChwZS8iJFsYgMhGa8ScG+9jTKBoWK1O+3qwYSyAbiJSVzMvxg3Xr/
XAS0DpQWWAqyp2glchrULh2Dp4j3Gx+EkbZSqlz+sp17gI9x2sF4mYHnicOnqHle
FZK7CJAjLSog1eITkT4EV9Q2kSCuLKREBaEKqSJQazGp7njl9/OTc5B9T6+5MwQp
fz7w6AXefIf9K/2+pzgB+noJsWKdCPhHtr4kS4Rl0b3GXi+SpvWYTDLjH4fr18hP
YW4ZLQcxKjQqRiJ2vEgJnHWM54TaON6z8KFpJWcmULGlbe8AqSxS7y2n7UGkaAOk
SuFeyLGsO0H2Hwsm2KleI4oZDBKgE8RDzfWyuXly2jTSTPGcJVkgnV2E8OrowJfH
Ggxr2q4UynY3hh+89CaDgw==
`pragma protect end_protected
