// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:37 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GqPwP+CbqfSO7yG4vUp9eZvxm9nsD1+UrqAS3/hOtPWWzcCOTJUO6Y6CYAkV3XuB
v4Vq9zkNzkGPV+2VRFDPaZQC159bLgUXd09EeOgvbn41Y9hUTwyuMdDamhiIwpfH
d3XT3QSmxdSz5RlVCRsh1vOKXABwziYxuiSsVsSGzrI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7392)
V1SIxDD9mwjBV6HmeQd03ZEEdu5FJqZfYJ/u7UwpnyRlSisMbalYVU68o+iCKXqe
ZsT58VF2bgw/skEO+V1aFPNL+nxRdcMr+zu/gWX54IkSmrFKqg1rRabFw4mRM8nm
MB86D29NtAz0T74QYgND0bj0LIkxzz0uJu8V6IBfUkbnF6NXrISxU/JCmr1l5Bft
emTzeA7NXLRvQI04GXsNV+UAZC7GnrLJTrZhck1pgep4BBXnQp0c6PrjMXkNOUv1
6QFZNWBxDV7qVsOvfYFeVm64h+N1fvo7M2/OE9BGduhCYgIzRwqZz2VLMsMn/gD9
10YhbUwO8vOILi4t7EKahDrdkqY+1qtO65N2gfeo6dpkddx2A2tmFWceo8Q0P/Kd
YYzGO48+0pwKlpCVxrdEvIZaORGtdoxrzD1pxGtbeo7bi05loM7hzW68jOkmcvL0
l3bckOtN5A3y4ec5Fma7r6JL5NssRgO/jDD43hq6Y62gYoKRtn+ACjAXVHVPjZ2E
kjQV1ozue/cHiNT02pbZMZgWORF1Rt6G/mCL8YVThsblXOzmsVm7HLpLFEl1tjik
+n+1CvOtPdcogX6Qy7P0koLhMFvSEFgVjSp5zTirV2g4NQQOAAiu7lyXy8H9D+r3
5gKykUH6VkfOK7n8xhUHqFLZw45CELJ0BeYJUPNG6Mpp123iz6Ns7MhnDMevlSUu
l7vF2VJzhgv/Qw3zVFocrDuf0RKWZK68edQfOiBQbvNHLe2drqqpqyq53j6hDlmw
U92M60h7UenRuvyVDu2vVGK49poEVAE/If/n9ZV0xXqwb5IMJA1ViH/sOMEPuccA
tNfYOpISUEyR4yUExmPEzYMRsZJcfAhGFwtMj0eUapRGGVsRW/5E93V1l7FCyQ6G
rCpcjUO/zep+YQEylqwMuLK3iKJKo1wmhtV1mdWLQWPnmlfBLg/mEfwEl07mTbkW
qhgNXGVriNHunHEKiYyXIAmskjI8bREwwwnkrumw0FQ9SoyZJCvt5PtynKMDiEPQ
mo1cURcWMhXwpWT0hN6+RHv5HrlUn7Iui4wj/ivrI4mwzKyalkAcKYdTHRvSB6C0
GITdZF3XtTCveKraVnAZhkYSHgUI2G+Uvrv4cgLDfdRgC1yC6LzqqlUgdQzV3ANt
z38RyYPtQl7i08QTDoVO8YNSXds1w57Y4ypHNT71KbMc18G9XRIdx+7ad8Skf58C
ZvudrL7T8GPUa3GscdCIwvBGx1OROIT8Rxp3Gud8M7eoFffPbQFZW5+AtdLKdPFM
tT8/IUqEBVKX1muZPif8qAOUrRJq4C75PbvXw1D2IyCzlkY4xaEQpkzbec4pidig
gT74PaGJEb6n46GO6dqsr1eImchLXTywFf0pi7ecqo7wiLlmCWyEBFLIsCpkEZ8q
PS5/gLbEuxpa57yP3HvNhyR3aWDt8m8nAkVvH7VHRlPWAefvnD16eInWCWFozbHv
RYdMN8aBIDybjTOJsv6LBGozDFbZYUcQInGHDZZTjZtWedlmenxRb1MiccSUZQyB
YkYAIwePPu1hSJ91Y1R4QqfhIgfrl9aV0RdSDAtULivxQGhj4UX+jTJHTtY/Jkkr
Ptw8vmAFZeYUi8Qv2A5rZ9pSzyoSaN7LYhXySOStWdFg6FX5pwtz7BL0EzgPaWQu
wCG2hCBkz7Y1PP+5o3jq/WaGGXYFPqWIWylIraK433d+EB8DvRgORg2YxhiOFFbk
gGRab0fzcrzaNwQxY7MSLqd2KjwGUM4PaGDWBhpFMF4GQOnyB3x/Z3yTEYZvGYs/
fp3iuyOF6sivxbzDaZIi8he+51KW8Z/PZwJ50nGzNGkoOO1UpMFxbl7B3cne5YJh
23G0gs2ms/QgKtkBkEbR0xMFEmnlRM2EYXNrsTZ5Y30VBn3S+1BIenSVS2DATZUY
uOgwmHuyZtaFo2CmrLNltOxrLQ2qj+Q1+VeWWSoeF2uC3gLjfAxqRl+uYj55d4gM
nrp/fYj/nFWZSwjXAt0MOD4X1HRiwqasukPmakB5Oi8LTz3IkVpHtQWgP5eOWQVK
Ee0lFhnjWQZb6c37h8k7LTLeibyu/izPhEhKnec1gfG1eipcFBhzPztaOjFUIOTr
Y5C6FLr4kEKLh+g7z0iiCj7Y0oHaAgfg1Sg5WXFF4zu+yQGKXOz5JovBkWNtZ9zi
NgWpzHzM4s5aCRpnJduhhrqLXS096HbIdctUokCAoI1nqYgZh1d9HSiC+KWHjaRH
A/wY1CLQY71yXrBKJIEDIMB0D4XmRkL5wmoKeel3Fka/0Sss3w+fzYV8HKq59mB0
+cYqJHumwiSAMy7bo1VIkcnx0oXJeDDAmOJ6A9xNA5NGR2bMY5Yyokh4Eoj5PmUg
l2ViCaOC8uWyQmlxjG6ZG25Iz2yYE33G2aqey+JeMUdXWLjjTjy7G/rC3O9w3+X+
8oTPc/gq+ydSgN1JfwnEub+R+X5sXTmRanBY8ncuThyKvOR3+0dbckThacUz7qYG
6hyT5WgoQ/j8EnEBlf0JzlzX6vRBEWDE4fqDsFn5mNeDzVIRabwdM2M0BxY1uPFC
7Q51/rHAf3S4YFPLc2Xq2nFvoTHg6cZ6e8KPeTJey1X427oCNTdrayF5XzwB5haw
JPi3m2P06Go8l26cYlk9Wf8Z8KZ+gm7xV96z08cVgyT2gyzvZMLiXV87UIPa4d8r
pvHRGjjtedcQFZAfcYCbm4R/aPEG/F/+4VMV0oS5qwf/66KB8BXU6F9yx3Wu1/SS
0HwNcZXDN4dUtJAX8ru9aDI91/iG1l2nCrtvBnJ1PiYMr3oDJZ7Ulc9n64DhEy6X
POMaVmssibakvkpnWFBnzv2w2mGg/2OpfMijPFNrdt4Po+w9cN+TubnUndNrG4PE
Xxx0vci26PEaD0dNMdLe1sAsRFA3Wl394CfcCe4Z7PibvQ1eWKnJc/GE8IbmoUJL
jLXPqOwDUgEcDuBfSXdu652+h/tX2xRj4rRmHvXbB4ZruMb8sQmGlbIMfYf6jhMm
yOXLvweuSdam9596mQXc8nZcmMkTN5s/cSDnN7UbaOlPhO1L3+uL+CLW8N87llp/
TbYDREzmGw4p2bdR8ULSsBCf3qnSz432EBu8fiGhsXo5uQGAhpbiTH5CZTPGwbTm
ytrqNR498drYYye3tm7m9MpdaJxZiwjRwF/9xDnnCU6GSj/ySKGqIV9+7D3cgX2B
WmQsDuMZJ4a5Ro5ZjZNl5WQP8OSexi9hdcpq0YNCdp6som+TTi7CFNwlmqsZNCyE
ZCqJZMsrIEr22gJZjcceBfPgzdIOJpCp+IF1KAW0KZ+asQQhOdUWpjPHoAU/QYaq
FcvwNeUnMaVJxuULZYgDVE/YHNaKadqKHMJZA9fOrCiaDnNBfoVawjYCAWofYMWq
nFWfpJ/F+gZkWl1IkhIFY6/Jd7tZ/su1iPAwej2W1RMR9vUTYvPfzDGCnrJyOvCD
3Lw0E3+jEYfYUEOl7Lfd+99WWmMhz2GhbHMMZlj4BvhCkhgmbh7QDyzOS8swce34
Qst5qhh/uNyGyF3ZApVV5uxJjyg3hvics3N4hDMNZ+ADLAzZDBg17PwFDi4VpTU4
uPgaO3yyWaRSbOzxfgdWqFmf5sYBR5QzOg1MPmEt1XNonx0BeP3iHK1q2kyikzaC
kGBfyIoMS0eFh/ugMcJHwt84qMzYcVgGXZroLlMSSu/f7qfn/sa0ojeGQyV2tUyz
Sj01rp3fOUYA4mkFQJzq4PFwZZooApTLDf3BRTLVQNj0L3bgogetDfN3bAw5fQpj
agiPLaM103eNMFNcFmJaMnDjhki4ZZVb+8mOEDKOhvdmLh9fkpeRFmBt7I7430ww
p19SEW/hCBEGyzlTuOADiDy6n43hFt/43DQ/THouRtpXhhHOnU4gtV5c9AuZoUlY
wTEyIGSmTBzPHjnOflAMdNCZkkP+9dgsCnmeswW8W7FulHkgSQagXdh11LUa30JK
rA9tQuz/0caFY8nTrWXly53dO2IDFpXXdNtgwBcHp9OeGyEYIkhr+Kg9tKykeEow
hR264M0n6EiN7RfkJjy+XjRryxCnOrai7FQ95EyTro/OkFWZJD/LI0qI81vzXbD/
VdjyhmPudTXRvxZan0A/JWogZC4T0uzAd5Wq6X8UqWxbDVlr6SXvS3BHXmBl++i7
s3TQUnhAZt9hHoR0FkAETD7F2xOx67YAx6wn1clNGt4nAoeys/Osr6LcbDPEiVFM
7tpBZmWzz9e9xfr79GEcr6LXF8dhTI1yFmwCIuNFGHfYCJ6hkZXxRgwsbsmU3iUN
jXYDo6yAk1UElxY+yqFNsewOn51rz3ZqC4Se2fpEXP1KNR/Gn+vd37Bau+6SRUqL
LfyOCjDhAznOGNQlKB7DE//PWereqTlWk/KxcOSntKuRhKKrBCkoB1RnafMY6uV3
WyHxIvzKeR0tAQDB2NSrPMzUtnihHBBU/THaQD6MaRRFsO9gk5xsOphG5tLjqzTV
EZ9LcLGUw1GSmOlSdqQ/EDWt+xKC7eCJdDd84a3LscokjkPOSanChAfOyEtgGUEK
zA7LmUHvoVVA1bbv5VXhE/G7Mnq5G448XAlo1iO1s59mBe+Ziltwfw3qhcUa0Mpr
8OzMBoVFd/2G8OldXH1OggaCrPJPPdbm7KgrC+8/3npyg0Uwu2QKWOuF9Urq+o1Y
BBSuNHoqRPUs8qlSN9o+G6mWppWdqxzifRCuTsr6/1oXofZ+O2Jd6MrIQ+fHNHjL
z+I2T6YjZZTxGmUykF/W4ruwRJJ6dZtmiL1pflyOMd533v95cQTLNgtZzH09Ol+u
ZQTqSNF6apQT4uXlsQAPzSgRdB57fk4opldIK9vH70/CS1wIu2Ar6WY+7glocZTC
YCvuL5V2ykEvh30xAJp4UjVSbqKz25mU5KeMPOr2RHqedCv78e+ex6/n3sK2HnLq
olwH7xTTypnrbHIitbELYEaQlL0wLT/SUNW5nbN4MbrFT8lJ0x6ra+1DgdzqTKtM
PhkMHJzRT7VnZI4RRAv4L5oon8dtrmrlc4YOpdoh+pUk1yrArus05G6w7dCfX6QE
sWLrL/+rt02XtctEShleU6RqRhO7AWw4T5g8N4yd9shCkxTvHHupIgfAEL0HjW2m
tzC4KqZOb3xdQ/leOz8INeScxJtusd3n8Hq2mqz8pD3Nzy8v3SPdpJkiphPVNs0F
jSZEjadXNr5iXmWDv6WXDo4lqAsmAo1qqQ/yJGSjDr3nu+ldQa7SOZcGYvCLZ9kF
Qv5LTJQTKDF1EmQcua+ygih+RYKYCemyTRHNWaACX6bhGUSVPBXxqHpg3ltekzLZ
6aNImO6GtfFd2UrhJ/uAqTL7+3nSnTc4DcE6GPChtaE4PCzecF5n1kBlwMRvqvdw
ya+c9xY76jlnprzV9xD3n9V8rGUSu1HlbyqL1crI5lRa8lkUv0RZ1/WHC3oI9mpF
rSm0g3c0UD8WDe3GKXSa3zk1efxTwp8Or3AK8i9/XvkboN4oOnP2Poz1nCaUrUxH
DiiMcl/F1QfdyQKWXtoo/LSY+KKlwLgg4gtasEBbF4cwyifVBJovC004PsyFjBaS
DPABMnO7ScOzmwK45BbfjqYbqQlDTgZCfRC+KdmY74pvlEuPYNySRmO8IGCywUgf
+AvgdU8sR8bNvC3mJ3ArBeVIsQ+tWiubVAkwuWetrKsFriGT50XqVAMoa+buJ4RY
TNWyjTwPXxtowQqplvEDmmK4OiIRD8wcivI1LwiyD3ZgOPn4riDEDWYG1w+BEf95
k84xUyx24fKLCGBkxDWjklsWIkKQnpRbeqFOkcayMuWTG7+Xml8z77eKQy4le655
xuz3d3/dafIbJrTGN7Eha+wVSRQID6JlX0EtsASs94P4ClWhveu0FErulVhke0Jj
dNPF54eoGiHg/bw6XW3AnT6Gk9brkZEbaFWAHJ4UFK4Wweeyc4wKj2iYPylWdsSd
ttwP2t+522hnUFnpxlM5Nw3rxilCjk0q7ibu408x93cZMTcE6ACbjcS5Rj2xQ50y
1DBhKJpkKvUgrYecmnRLIsnAfypgeNv+gJBUemZ+q4EInOA1t1ygdwj0YtmbdscU
LAl6uxmKOHZvtwhLd60MVaedws2sO8VQNa40G+iU/ylzUzHTuiOIVl2nZnshzBlT
KfUlWpkdx2oKh7jum0KJ6aU392ldRttupJxkvYuAYvf+iglbIlr/BbfJL8x0nU+R
FZ2TKtlkhqF1mV91bzvL6HTGzyMK5bAV26A3AxiCNPNeUAFIaTvSwp3Vu8NQ+6Qr
kGLn8Asg+yuyq6lr7T70tWIxW7z0IgAqls1KocxYZtW4p6aKWSQG6ik2mH/IwYG9
mySEeeXCDjmFDqY5KhCqa/HWeQ8EfyI9TKMnzGUMnL6D9rcn4M3ymYOMjNBCDibk
8hzxhJiHQup6fB5SHsnP6JiQjMJfi0t3CZ/ajVtwEatDX0IayXpEmvhgLD3qxxdc
i1FihnT5BaXC92mtiOocSqt3715sCdmEeMTY/X7bPxrndNGVS7TVV+scPd7XjwTI
Y7CovEAoN4LxAzeUJ4g9NNavIgHaetWzMoonJRg1AiXJd+Mz+oEN+azLoBYWkZjx
kNTHLz0aptnw5Erx8QJIYVYXnZa0dOG4UJUCtQfq2IxDdPKaYeCPk4sx9qcZp2ii
xSKofqfVGMwayPvedjkWmLt/ajrBfMg0tzmUOqJSGrmXiIlXmrRwqiaWTXgxXxzI
2E56qzG/fGaq3DXIyWeSK3ulkN/hFxED4l9TBiftXhTmsW5Hx/4Whl/5Kcs0xeiJ
Uxiiy+Fgj1YzdaWFAnt3PQ1+uGC7FEMsnzusF6s+HWHOaoKPzPUa0JX/CerhgLHN
RQelRAb5jafoSSx3/lIAXvdXSU9CTRjHRrvnu7SRbiD0fyPMoyhgUtCzA0LVOQNZ
ptDKQn5LTAGLc/H6k150yWamo3sy7BRGbcsxA2Zuc6yszGC6F09NEhVrhXQTLdmJ
Er0fdwveuIDNQQF3YQDFV+a5YDioQzQ11HbwZV1ZnAe+xMIC3vgDlOnmJVWE1TLL
c4NI/8hPfJePKzbSOYBGuORsTsPa6oGMRbJq1Q3oDVS7UFVS4pJVh+l2ISy1+wSM
5+vbhvecZUnCZcmjhNbbbmE6Gk0l7HriQcK+XYM2g5ICjfzUkVqVPrfAr2npyPJY
atrEVltlbYuCfi150xEB2omef4CrW1FLSRHQKR2OgpwpviOkbuWSp4IqEH+oxukv
95eqKLTK4Pgu9Cx1TFR20XR+IMXUjE/zoAn+oefdyzCQ5Rvb8IQZHFHoX47t5fxm
vwIWgIGtGXx0DUUaP167D7XztiHEeCXiChfJ/RY7yot9u2A9FUeRhAAnnIAqaSiL
djboR9CC9knz26nBUXbvgXxsu3Zuw/DjYD1sKCJYeZpTrtU58J3cU+RuLu+k3OjI
hvCfI69PIIIKT6woVpaT31o1dZ6BlAaGQwFhKUP9zPVAKuZjZVHb3UID/LGVJK8b
yzVmo5CjJx36Pd/xXR0ZwHNJhAIV03cfEc4YopMmtDNn5EEyggTZA9++kwr2bgco
T8+4Gf+f3xgN+7fjJMVgsU4r25OkIBJwNMLoiwKSoIOOEN2rMpVTEKjQxBUaIGt7
molvnUeGna61qRd+4pRePRnQsAiERTKivUkyutj4ryN+xRzsgLXkUAMlK7X+I206
DtSQhgwoUonzMoBz1X4uhFvrVQNBUKln9bDI8YrTj7yJ91aDq0p8Qm5XwMmcjyCA
2cHYNz3EcXZ1DivRPv8WytXY2vHTgl39IqN+G5aX77JB2QcEnjOJf3cSXhUmxYCg
5JdnKHkR1DtJHDcffJmXayvalb1DFj06BhJLuNwrWjWGIf+E3Q5gHcCOS3qwmhlF
EXKl7NNPgXrcpA8cEx3fWWBRQ6rO5w+dHA1Z3NsDD5LN+zDuZ7KxczjC5JNGlq05
2Mxfrk0Pi5psLSdW9e2pdHk32C7azSqF/y0wFCo424fSqrZjH+jQpRcPEMX/51k+
Q7SBIrSomoDbbVwgk82tbZPwkaIUi4EhKv0lLAqNlM59YU+q6Ln8wK+Jrizd84BC
K9N5edQ7janRtSMnQf2Lj8ifhK12sHXRTAZyuYaauNQ10eZM0MflbiU0E14PIwhN
P/FzF3yT2CUSl119Qd3Y3dQZuzdTWIbr7H9gOCOP12iSmFGR8rT9kLVh7KHzGnNb
+9YD8caFuM/kjrq6duFYTkE/4s3yjqtcUKMAA/Lvqpaxwyc1FBeFz8M/EniSTPRF
V2LjYgnu1C4mHk/rY8IvOPkqay3MiIHH+2yBRz9dMtKVqWR/EPtMd1f5kbOLPM4h
wcuC0BAkrd2fm38jqaZgJ/nM9ftnxPmyzGmTVU9NddGi9fL/e1C1UapwfsXDPQZc
zoOid5/vfFvHEGjBfwkcEb+gOAThr0wDhpSC87Z+CyiyNsr46XQzU7Cnlf2BWgzX
DArAhlRwXQawVrnhfhubPthR8qDBUNfMHGGYjGw7qYAYaXMi0rNVe8ARtKwbRlu9
zzmmyjj6H+KJQzKFwszZ3342uKdAmWCjBegR1Z6ysC2Q3vQ+AaZmtEh7NFjPzZ7t
pMTK3jc++nUqeh112xdvD/bxSC6cX74SC835MUbHaPWBga22xKwIzu4i7hAREauw
KhVldWrJBYpMJh9V2qdkOidjsaa7BmWtQBBFLFs3Op5T+HhDIOrnXgHp3ju9OVnn
zqnjMM1cq9DxLxUME3UmC6AN6S5zqx86WpfLFNe+vymJBE4PN7kFUEXOplxAumjM
dCVOMWLZyHUqC3m4ssdHId6Tbgb+oRcavDeakapUrSCwp/n2yhTotDJ3L2b3ASsF
nJkrso4hay7/CSbTEZLqfpfBlWR7yKPAUsv81YcLPpjsxUIgV8MdbX/t2LW22jEP
Q1jrlHuEuup6EpN5FkWxU57eNzkK5Sw0SJgcj39lxT9hZ9S3e2AEtn8mKPkiQ0da
jsQJbRmBgWqGUcRHWPouvgTvC3g+qwMOmCp+47VAwJJLUmeDwaeziCl91ssf8yM5
zdjOW/dKjuhRVrCnQqCXvx2V1Iesa+RgGTeUQaiZS+0pCrK5HbF8lRL1UInNoNJa
8ZDiYQLb/rk58vuQxw1lDB6GGL1NtpzdD3X6WDlj6P0OHr1Z8rQlOnGJcHCX892z
4ntewW2aBvqkxO3mdIgIiWvbjmxxgJ0FhejhoOMNaNKP0LMt+on7XkMmLsFi00wg
DYiEvxg2ohoiR1OkwY9CAL8CYjcnaLmnKfoJR4kfamYYpe/hakQ6Cnme3Vn+7pcx
jpRwyOHhXRRonVRZJLUnL3LX/qwcz/tW/oOwib+7VuJyN6WXwmqYb3LuLoAHGtSD
/HeWeRREtoGl2vepLnV0pizAft1hV9UTdIOO4RFt81ydF7peA1zS5awgrSIgDqJV
JEILr813F3hiijA2htOvw4mXhikGaaQWPOguXu0Sar2Oay7Jyh0bZ09ON+L0ZSYc
dY69IdT5IgvaGt04vYMR2NtM0QyP8Zd3brS9BH57j1IlQcg1zt4FQWfPLmKwJ0i8
MGnmbwYbjll42XZrEFndWY9lFCiJCOvfbGTKtff8jIaLvArWrjCXbWeoVddnIXEc
/EQPNoYFH8IHiWObFth41JvgNsAbJuOudKTHFlBE85qor/XE5ukWL4wtT2Pps0Kh
k5lEZQMj71esCVj5/TAkBGBVilioXvju07PQG2eurd4Q4OKH0aE5Zcx7dBRdXvGS
UEpDU3SHr+iD2p2zPfWH35IJWdIL9eU2hh57WjYoKh6c9e6H7Zt0x1egCR3/PiSf
wl0kljABljFFFQ4v1jgd/dyT2eY60tLsF3kekuzUZOr0RIUbhptWX5nTiFT1nBit
`pragma protect end_protected
