// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:05 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Q/fA11Q+ROCqoGhGEdIz2sxI9MDyYITDYZSYRfwkMY4SRcAtNuV5LBckMZcffw8A
MDSQYrMuuSZ+sGxwCdWty6Z8Hvn6hEfpv/qdwLKh3Y3cHarkT0KF2MRfmnT3I4Yq
kf3kynYQZ0QIkxGrezK4u6/FslWDQcxUp6PYFSdVLTY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25680)
PwfaBMnf3np66zZy0dsi55cBe8T9gvfRWBgdUPZdzqcexYqZfX1eCx2dBEi5Xk5E
YR+lmAB1XFQdfmgLdKrss/QoPQ5pJO7mZDrbApfgJyOOGgQT1y1C8GvoC6eo8EQi
JExB9PYlqhJR8oADVIojT5xaaquLuOPjoYSJDDMNHQO+S+M7N0NalbXrnPrcrXhZ
fDVfwMZoRAf8zxqxhOcc/LOYOjSKycuWYdEdxllStKpbWU8OUagkrccC6RYtSBze
H2Hh3Wb/iIbop7LOdY/1FE/dwDpeiwQIQidfynv+JA+VDK7AjbZmPqoUMMsG0R7n
6ks2MjLr1IgCrvHUIs6fzY7GYL33Z9XuXfDGDdDTghJ3wGPqDUdz9uC50KSqn9zQ
BnaVLEsJWIYFqcXbZqTbThc1Ew2adQTYonyK44rlR6z+zCL/VSRoqv3vDolznBVg
csWE/TmlU68lY7bzzK5iRzRbJ0TES7IUwMHAvpO8p23E/NP8rXozoOSx0qita9nJ
znVW0YQDK0pxzTSc3wey+2NlsMHK29B8UFm7/lyiAUyQiW1C/frkEQO3a29zlQKc
EQQlnv6grmnI/sF02BZIpXSE9r7xZS5JcwMZdNp1WGxJ8gEMp1WblDRFpdM/TGD6
Cv+rrJpyY3q5dKLmpDZZQq48ZOy/qkJaikMZGRaNNYqB6IxhdY+KmOn312ZSncXo
rN0VGcZ1EioIj6CP1L64Bh66/S33wZQktrKpPzqqmwZ7UY8kS3ngdijB1jPfo5IZ
46XA7Uhs5zD/EJVIXlKkUiiJ3k7RNPe7aRN6I0/L7TOVUhnL81aKG4HFQGTHUtQO
K4weAtqdaVULQmiDzP/F7bJlKtRBLAOHsn3YvzmRG3gP1EYv+qy+xQaAaEpLGoRa
DRzVfLfpGpNJqkvhhscEalmZ3hmnWXvEOgiDBJEH5jGGDik+ygxH/A1Py+qeUJbd
j71ChxtrBIm/+iVH8askJl+4/7XKLOMJuAuk3UmuT4aJvyy5zE42lE9RyBAT9OcQ
IzY5kVJVVq63IhhlNgH5FLlxHyDZd4+Gqd6y+SStuJlX4HTnuVc8uo5HOOzFI/GN
XkA57P32o2Nb5G5tslfWYpXt4H9jk6YNXPrvC0GFqXukPNGENhtrpS+M8w5Q2eOE
AX0KdKlmD351PDsu9upwJsnvULFI9raakPYTxWTVDvJRr/sElvkjCHQucSDFXSWk
4PPDWUNIt2ioJcsHmSXOavjPcrl47TS+0hpuapQeZglgmlWV2WYzTDs49Tqt4zwV
sIgB8kaPwYtJMk26WkUOuKeJi/uECkecs62o/ftWvrmTkntpVEfvuV8hztZAo43G
Sk6L/hDFjMx50elauRmmg0A3kLDEPT+WLDBLch4LMb0CvMiUvd3IZerDMkk6Jz25
8tnkOMexHTbcKf6A9KGkJ8FenwwOx6rWg4/L8vrkaDS81JdK+DZpHA3NkzcyKHFZ
QhSQg+JBAx4c759e6BpWmMUbHL9KVQBqX6DZCGlbSqJzcZ7x7DyYIiROztBLScXP
xlrpVyz82mKRwknHr/8QXdagxLfFB7kF0yBk4UREFuNCT1wENxm1B8R3qREJDiGQ
p8cdPanDS9Bz2ibxm4H6aDK/yiXLOpvVSh1Z14Q7ILoFPJlokLtUOUH5MoMDbsoM
G3RF7nWOLeNG/EppPACKz1bVS6+WO+hwO/2zLkJft0DaxKfcD1i73g02TJQr1yvi
l6O+APxMtzEZASlIlDw/GtCR9Ce3OrZcMH3IrRywhf/ZcGupKOWD6Poam6U0zyMR
4j19pVTH/887KWphxfMGBNuiRS9hPm49x29ZvaIDZFFtReW1EJuOSZ+weK/Rl5h8
x/qVdrOqElWuKWzykvWewgT4S1tFLuDtoIzHLdJWRHvZoaDplOsI70bTf7MOl6cw
vBxobzwdqjs+orCnHUvNIfTVqmednGCxyQnm8/W+0NU4dNHZsJV1+s4qNA/5i9z4
mVBFn3cCftR2ssZIlaBjRJtZTCnEJ4HquRP5BfgszwJgbHw1HA0Kd8PWztOv/sQU
8W1OpdlF4UyqycqXLR/Hl3Onk3uX4hmq4FEwIfTujMysjy47ZWFJxtHI4KIYkzCl
YF7TcZHYan4uLyTdXpDdNd5NOYdCHyYUcZ06EmJi3WphfZoCV1E7Pe2Zg8cExPoz
Hzc6CuRyAos+Q8gKBfDuw8JaxsWej/HMBo74EzqepMj4T8Fnbcgx0tv8BBArS07r
yzNBudD4sUn2YOt3boRicpF31PIDJoKx+U2LHkw32cn6A9XSyb4moNZbrQ0NaWpF
FXeJM0Jv8QKhwDN0wsSJcPKJ3taiD3ExPYrX2PGFWZE2EsxepSl6DQ7hejNdn/2w
sNXmC+Yfh0ycRYawuoR/+H44F5arAv9a4zUMjgS/yyzhrue9c5bAoBEJDFMT4S1G
Mh97L8VDjt140+uC4Y/U5NdENq5SwH3O4zC71bOPP7CwuY+YqF7teHiRfyoV5+Dd
WtZGFTQr2UmD721gNU4wPnk4OoDbnuNthEN4/xe2t40D6wiRUAgMW4UZB++Vu7e6
ye7oBRK/NeYKOj8Wo5uN9J26TYSl3MurkmpypA1Kd8iYmel3FR2MWiX+3xf1cFaN
JzXTL1KJwl+1/gpLYpRvtCNLXItWr6xMPYan4D99ch/n/wQJRUMyitZ2vXWXKg/Q
7ATSoRUZj/pZQbQ1wAIDt1e9DsAygaIa4FlHlmAK+o9diONPwi3r1vKsg2M7D5NJ
qtJbrxv+fc+2ZlarObXMLYxlEhIpfrYp6EGLPkeZaniNZ7kDVDG2XNAqi/+iXGJs
3RvR9/ay6fJLfiX53j6JoCVQkLMwk//lj28WHR8jiKPtZLCL9ArA5U+WiRz60luY
SJepFcdrUL7JSTocpb73W6D97QuzM8lakDWxeiTqR4s/mkwMOF2RWkuhpt9YBBEA
weKczpnlxnMC1yZ535pxbAfkq10IltWLx/flPDTacoRsD2uLHfPyY9gPBw3stGVd
IYAOBuNKcONgQAT+lGheQdllbcFnkWAzMoHkn23yXYN3BCSQa/SyVVfGU6QT5L06
aOduUMWj4TczaLZcCTkITatZfQN8tmhOdtoIOFufLdmRFGyeS0CKRiKF2P7Y0k79
W6/UTIdeMxwulzqhZ4d4X1dEj9GXtMJeKG9FV+xYs/371dDb1VXq1mc0RWTHrXy4
vRVgNhtSeq6J03emgh2aOzcKNsASjS/T7jh9bomy4n9PRAcZ0oTTS22X+1l9ef3P
leLVAPVdqvKEA1Zf+VijeLHaK4NMusHMMpN5zSWNvpahsImM0qyxRev/tXmG6KWm
COg3HUnvHOnQL6/n8GnmofCnh3vw6Qdxu6lTwE9V0cmajzwn5uc81gTbRkPhQzD7
5Xow4g2lvFOivqN2oUPlHfjsZGpYzk1qXMZJFoofD4db2HPPWJtLNL9xOe/gDux+
5X1sz/P5c/LZy2ZbXqurojB/fP+BGpZWppDcxixB1vE0/Er21UIzQf8c10iFnS0y
EtXmmtE+ZnBu+VdyxPls1HFjHaLf6oph7wChVaNizwyTIkvrHB62Im6KbStuBhGv
C47PgeIof+d7KadYTA2hSNjXVEmY3ErrS5fJ9ZQos2L3jZp7+KdzHes4sILg7uTG
gZ5NS9MhuHPTDaqv0H56qaLkRMDqjgrinPaPiob50RTCTpPICOioCnPUT9ESYjr0
TumEM8r2wjZMM+XaZ08Zek0dyU/jYZEDTjSwVoYlmhlTTw85jQu7Qg63UlfjySF6
w50uCslAicNyBQCXMAURprculNkXn8ukx8JRZ8+VcStGn6UjsLtZKf/0UzqReJd9
hRMHYG9QyRJ6ZSPcywLZMh10tzutvrYW/y4pCdfmKOP/G7MZmB5PzK9eaKTjqoWP
pTrvICv6ujDLoiGGCoqwSxNRyqt2QtRR3pF/tcc4qTrsfDh12XAJbYcnwp+4kQ+5
QA6omnBqwcxY5yXLI/ZOoAxy5tksvX6EMuy+UbKpNwSKP7M5v1FmgmPK0+DBcGGu
WxzUr8GhCRcsM5hP8OC1VlXu+7+fhjwiZd+04p0ll/mO0zJFzqUPyGZcAqmKQ/nZ
Dz4WqMdLoT5Gfmuw+cK/VK4Y6ivSojXfoJsMHhmkrj82i1+ZN1Kl9RX4ByMJr+Vu
PwvRo1k+l8o+x95KnahBeagV5qahZORfT1mk1OXmJgEenodGSN95WagATyC72OGh
/jW6qJjnF3t/g9QySwPCpEVavCJqattYcakv0xauQK8kiEnYDjCmzmB06ji9o+sg
Ni6qNa4QK8cF+3nh9GtrTBeGG8TMbZpNAcSyec5qTLUmPLxM8FVjUpNVqWX6PTLb
1mmYIudgmf20X4tmhAAHD+d9gvwH8+aF4hMdjeRBmeth+SWb5ZELzZOm8J+lwp7W
FufNJqTWJX65yByYPVFWPkhhW0gsM1PklbNd267k9+0sUN6bopHGuxjeQpfM0TzR
GK6DKPttPuT37I7Awm7oabYKmsksyksju9bgNRYpLbk4mTMdt2GDmpwRlEa1MuIc
o+BdgpnpYmh7vgeirwptoXL85uexPV77s7Vg3IQRj0P/6GJHYhuV9mDJTLH7k8QE
DKz5ZJJ/aVl6JmR6apmOfZQ1dV4pB8JYej98X9DN94PB8/exzG5f8lYluz4ZGcSS
3OQoh8MjCpHRvO+hJIMlMy84+GAquVPcHI15BhTb3YdGu0hhMRAJApg3X/aACLR9
aq44H7yaZbdrS2vu9QYLTs5uxDXieo1e6Kz9k/Mp1JgHOwE/nwXiIZI8ZCgNZA2m
C9PBxKVuKG+zO64z0bOVadMtdnj7lTSHnkz+LHOTy3/TVS0vMlxdpVfijt4eGXmi
IwUnutIGLAwrZjI1Ce6Wu8hcqQ4lVxW7oATpQgonJESAT+Z230O8VP1lg0Z4sc/4
9AvfZErIJ3B8nupFyTZN9Y4+q1/zppTvfreiJ22XlQMLDj/h5OKd+TXeMxCY4XeE
uwg0geMUPdRPb95leKepJllU6zftZbb0+7dQknm0YbUxp98DQMSvfQcBfXiFrXQA
KZbhwIY4cX0wnFMX7ekPSIp9OcOmY4UVADoVQ8TrLiQ0CewpqdgrerQ1laXsmQ1N
pQaMBhwORF+pygddoqdjQgjHmVhew1ig3XtMyKfImMOHimZIbyW/F3VF80LJY6e8
JEgpqgATK90uXTw8KZlIF6WOVLwydSVPTxo+X/waBxQiq8dFsJ78IUJ0rYTGSACt
TIkEojtg9/+Yu83pP9CChWra1nlqv2PB2AuGMKPgUCuicW+tdv7T5Ov3SXo7Uhup
P1wKWIHGvQofdJaj6c/m+T7QFhgc5OvVX3aJA9+TjMjUrg63oQFYdARj8F2Hg6YG
P2pRyRstaPdWrku/tTS1iMQZFULGqFk30HYLlrVKwecw9rSAhhKpghukUdZHgLs/
7TmOPVjyFtIyvWb9K1jh6H0RNiqaFO261C1fCjqfaieB1majFC4HSmc+cuNVJHIL
yB7C/1oFCB5ICle350yb+5xwjGzlEUB+ROQIYvSXoSPAu/SJd6xkhMg2oOTwgyYC
KoPowvMbXYG8+qsBpYx3mapvsFkwGjGrsXPLg0PDhrvhAfMziBhhDs8Vd7L1UPOj
QhE4fZmxSo/yFlqd2NzWqXM1fLsZs9qsEwNZk2GigD2E4JJY+CxuU2G7Xzkfderh
WhuoFw5sY42XprbfoiUuoHhpcafElfS8lkl/hxU90da8N5zysFtgwZg+CErSj3rr
HjfeQ7fiIlxG1f24/tq6UXbdmQr2XoxRxR/0xxyxsSS55KDCBTw0Ofgajrw2WEk7
T+wGbpRZTkH6byU5vh7rk9WRIZGjDOX7KJc9rdYKJSmXaz2c5medg/zeR8SF/6/g
DKyL4fQB8OW8nh/jFUoOky8v9cEzsYts2X+dmEyAfPaXpab+BgvgCS51l7t1hsvR
1BFmN3FQIXBn4jNHZbKG3rnbvmcU8699PZJ4CXu0YLa2gw44ftiEUatN+hFQoPtb
A/XY5mC+fZGuBLcy2DV6J37QX7DI2YAms28nK4j9mDvAvQUoctK7dRd0z0yULpVs
/vtFHGagdNgfGTgHnW9CwUZfReRxMDWFV9qpJgBeVtnGb2wxpyoPeTGAZZd5RfDw
AZubiBYCbTiTKshuuB4nqW3J6i8GHL85yDWTpRpD+qeeKB0oBtUY6PPcIU1BWv02
XK2hnSYhc5esotOtSYKZDUYEc88k7zDzQCqPdjm4vr1OibjpLUMHXRLu5XaXW2ms
ya95b7AjY50AggUuvGLO6U60AYDcOb/0T1URvsudiZlIzQkkbpMTFqVOLMb0vp5A
+dlB0uzrCayNrTBMWOXwTu6Ky3QGS/gALoK2YsTafA5YlHU8A1/f+oIf1u5ZnoLE
uL54qzaRAgMI/edDq+2GZ+v7QQjwloVPM3/bjY0p6UE7L3fQcmi8pu7KTIqe1381
gt9KA6If8n0R35RC4Ie/qx63tkKiANIf57nS74DNMttyIkELMmi+vV0iTqZAEW08
igoJ779yUTyHLrHTeUcT2ZDXeCLm33kFE282bhqInjZAQLm/iGZ3LmtiBArAwvgl
V7WTaxsCJXaVrmZhE/kwGI52bwfi0leh1SHXYgA3VVLAXz+/nMUHyzRzd8qegqAM
ZjXVPBtuoxK9H06sGPSFVX5lxZLZS4vsRFoK1/b6DelVZG2lf+quDusy7pQUlKer
XgA4jPLwv6h9O/OPv8kMNdp2iprGW3mcoB5Z9BiEJ2yiWv19C2uXxyvIAEn3h8c9
0H0NoBWshRfXFZ6WwLod6L41GYQYeQXmQw6ILMaoEpfo7IhP2DpJsjZgh6EZMdM3
qTWp4V9uraFtKwQtT6wwac11ylCDYWOJy7595yOy9V3yVky9cF2QnwzlfZnQCFt1
INyJWm30WTRsggdmK+7Nj4rDjf34nVDSXl2QKeUDB6HIHVOO4TQx32bemS12xkH+
q3ting9aNWyC/IHtOhlwt2bAUS3LphTUK/vBJReIboQu8YKkinU6WVsva3wLOW9y
sHpS7cBlh8BkHfwa0CaGx4Y+9TQP75fikYabB6p2uHSyaP1QY+eVDGTRnSw/tZKf
L4oEV0w0YdcEed5iCRRRrhkNQxkb2Y9FEmiJAfpsPC5FtB7FhYCt9f8eVIYMm1d6
WxIslL0hmmNvXzRiKPBDgdcPTJ/bB3e8KZp/qqUqABPEIYoe4fwWROn4fG1PSBVs
p2uaScvItAaUQ05nsJLN7XxSQx1Tds6EhmHRHwnFhy6u8PIUiT7LK9WTD5pURIYh
zWK5AN1+1tNZPHkhXvY7MKDUDK6vXw6uN8TG6ojtvVQc+VAd0f2F/VqtKBzK4HiW
NoHgRaIUvGt8jp4WYJSSILeIpOBHKUFRq3Vsejzg12WQwVGuyQtF6Ty3y4TCJ7I+
2vZpMWSTEmCGQwtmUvapzf4Rk8vshJ1FbUvZ11Fg+nYYixJ8sm3Cy9/714AjDD/I
HbYGtEdg11S5j2MSrJo1z+MXnIjkQ3B1o4PGLiu0+50b02j/7mJVKy5aiuPffEHG
fk6cN84E8jsbIRR/q1FdTT2J6y28m15F9nkYUewxJPZFEhvvBX/L2fOe2BPGnHX0
cBFnvlnjVEJ1UTPzTUsbEU7qtRQVMLs6CGeQMJNE+5BQ1LWxiTgthzZWaYQHg8rt
5Apniz/VipN69fTtXAR2g1cJrfpXvl0F465oVyesVnpEc7PgPhiqBZ+ljsgvjMer
dHU3ex+tc3zaTydKLm9fg61gjtReAGaSrVwIO1YXBV0uedgOwKUUlJHV6UX/neGm
L1LYWqDOpLP/WoqKyL2A6TTcAmDeHjBXSe9pnzis8QlqUk4QnoO/iYVrU+t6U1vi
6WaxZvrJxCp5LY9F1MU1IC8FMCG6fzN5L8stbk4jPD/nE5F+6nwgsvHNO9hO/u2m
paO/3+Nw5f2GEV45PyNwCM4cgBoysz4+lxHPZmsnxcST0m18hDC/Lgxlly+SaHL/
GQv630Zi1xsW9qinuoNkIOrtr2NVDHWS/7srqNvgpaXCfcfsXpN8YXNWaNLu3rOQ
oyCBKKkDC6tjKDtyyQBWI5XBlfU4h2kykH3n3PoolVZQ+c5onK4Ld5dFHau+pMUH
1q3Z0r4td8jR3HoybafeX9Lp17S8RfEdrwCNkP6QUZg97QlqVmiCZnOUeb8d5RiZ
Q661rzrsf9sxoCrPqEyRRo9Kg/l4hYhezeqcmY7wMhUPKpvNr7fiIXjAi5KOdsly
BSegY0XYAijazU7LonSI7LGK+2ZPteamg9UqgVZokWpiySnygwGOyhtJiFcmlsG5
AGURef2Z4/fziVqSP/hqXLAYX0iti6suhW0dc6DAUDNrehRUPRcqtMtlr3tiGVw2
G6DD+06zEFpjvUhbkIEt9e+O4mcDydX6/SkxMtt96uzA78Xes0Va86XqoHLnrlLZ
Lz3Pg6lBxLMFyQIYoEFtTzybhk8Tcfmcv5UklSjyRUuaWYbqF5FvNuH+BGBMy/24
N+1tBQmN7fzYUMV7FDin6HrbNWI7391tvglENvyBYuKVarVYq2wvVdfvxfgUdwmt
eqCOry/NDQ/Ck1RizIWCmAscZPAZuoA1gc46+zLhrZdP2T88y40ozxKPXrmDBqnN
ZNUNnjty6DdJcEYgg7ttTAgpPOgmpzCXovJLWgtGl57xLQND2kAB2Lqo0zin/1lo
aMrw5cIIzpuepxp32Loy9y325irrm5u5kA7AV+6RbOXxzZ5mGobYCe3rN+t87D5D
dHCOXBXJ6ieyUv7PakQVin6vUG/w+YYIu+Nwj+cz8/tyB99Is9orofYGpjAjJ1uJ
niWEIQCFKw2Tdcz/i/1aCAmvPaseuk+srfuaPm2CeS+yuKFyyHfHHod8yBqK/0Bx
eLfv13WcUYCTZuM6j77SVEFig9FzyvST3Zs2ujEp7lrR1E4HK4t8jd1YdPasrlrc
vPU5iBuD1hJHKh0KpCJJOFgWZLdhcakkXPZR9llk6q34jt9F/fGePxOoyZi9iz9R
0l9dQw3c4c26u64A1vmR8BQukFo/74j9T0OrDHfYWnf1TE5dZu/hVB9oFrmNTMYQ
PrS9QbOdYLm2vP9Gq/9+xg4vwy8winCPfJzMeTOxqEnWugsADEbBSvCifYxhZB0K
kmapNlwBZ/iMzMs55MQ/5M+NNJmH0uflBpLiIjHJWTJp11/Jk+b/VCtMOaV2zRAB
PAJS94fkAXOyPwJbbEj31Cz7zmC+xWlDiJbph0aajbWYu8tNLlVAF1rDhcEnNSsn
T1h/Uo9PW7wjTjtw6+dsdOvPcah3QRDelGmTZhNA2u7cRtiR/tdhRXZHFuHdvp19
ApNAs9GWf5jE1oJQELFwOHiuyZkJRgyhSP5kZI6a/S0kVcBbNwWUBqZBEFGhB2nQ
FwVqjGPL9h/BcsUuXRPTrrZlJ4KbTWshBY7pX+5OPJfGgRY7J2gX9myHbnu/XTwN
YogXuQScO4F7lkyQZgQWyil28F67xwMiMQDLMRIXesJh3RgzLtzgBii3iyv+6GcU
k06tD8v9K2Dj2C3JYvOH1uJb19UMhUaLZxZDzCpE+FoZ1ck4e3GFfp/1utWTVdXH
yvxjAg33hMohSa9u+RdRi4IDQKhF47kHBC92IFLQU3tbFR2KJNpk63k0ehlilPc0
YRmcXllCZUDwZ46QGiFRKLwHeSBj301iFc1v+R9le3W1NZ7SNlLpiTpB73yfZSyf
S2DntHcq+ugOnZlHt1HNTlZjoXDZPvRuGwP4TBypys8mFGkLasIR4eyA1Gmmc8dx
AfOp955qQWFpfiMsISPl0SbN5WadQEUiiLG4Ikp4+tv8lJ5/DeMG2XtKwhKexYoo
4rAlqqOUz/vXaO3kRG7UC4mlARMqzeVwu6QPUOV53ny5T2snt767r5fQ27stfw8X
1TF3+jS3yeM/E3ZZyWSD5h9b6KflylmUO4izKhZJx0rh6i439AOU64lqmzx9PyBX
AfSaRdr5ivkdTc4WdhzQE5FXuQxPdQYfLWWmwWckMtbqDXpCggvv0Ah1p0a3Z60C
KN+S2bWNCszwsWJBXw9fDfw6iBKFv9JKYg0UQIrgNOZO5BbEDyCywJN+zDMlOiqG
JUfs6nWU0UWvl1e5cvHYRhefAs8OzioxZ13C6Vo17DlQ4ad4YR/Op6Uvu4FcxkYl
zSc2oZLs/5lvV6z15bipUcPvRdExdiXBSM0y3PBZtn4sB4dCVcFmL1goLt+Rek84
2yohDhxHIhzNNCzGU9KkZVkyrubHN+5WhGyMfqTS5BjZ7GX0+vkSb1wSulBPyCQr
GVLhF0b8ZnAybU/FFForhQNJ1J6RiZ122egsLfDXTT6on0v4vXqe0JzeUhutJQ3B
zKsXsmZQtaWgTbtSGUgGxmAk99X5xlWI8BgroH7dGnC4f3R7J0Dpf/J6mpNeEgwM
RG643KohSpuNpmdLB+u445qh9RZ8wcBHs6vKHztT5A5N8WqBcJmlmSPhIZ0JmFO/
6Xmcpj6WfkMwiOm6CZVNdYvwUXwxcoS7d2jhl9bIGsQI+UecAiRprJbYfTyT0siq
rlamXibtgSbYsNp6kuc+gow7yVegRZRBeK2Cyk3klvPTuQWNB5L2nVKdzJkrySBt
JUaC0F/M3UvtUWBzw2rwwEhyJriPdWaglRrsucoZ5OGxh8S1KIrBJV1ohxAUzDd2
f1tVIZ9Xi2Ty53ueJqPiIxMa46d4JIcZPCqrLX6I5mpCbWesgQLWiOP55T8I/iD2
qNDMSAYdxEa9/CymvSmwsbFCQd6yPSj7wwhLEahHuVQr0BlP/vrYKb09+8eST+Ys
j5R3veyay9+uy0773rW7CttAZV77DRkYtoOzaJ5alZ/FDihFgHr/bDJfPRgj9OmI
McLQdn0vjGeWsjkFyZUAfglLhCGByACcwYDwr9YO8KhstUNXrldeEli158HmoV3p
Nyx+pNvsWavSpidkFqXCaqnuYb+liy5l7GpMdofo/DXianAlHrRnscQoUdK/QFbg
Bgm69JqLctF71bYQihINMkuzYT8Fu9B0eORTldPNk7WDHOd6wB6mhFRysnOjFHsK
xnALZsKOhoWZBchi6Wn1ILflFDXRxPcuIzzBFZDYUXXeoXeZJAcUMHLMGjEPZBIF
vJJkGl+MqHwMFwdBdpFwqXIxjE7W6vlKbrHeZSJI6VGS3DD+aFTJ0VyrpX7wJWha
drfEDCtJISA4wpWs+fJUhF7PYRZVwtKC2Jh71WX5VyGrJGCpGKVntLc2DkFbw3MH
O3e4Ux8rTu6C4kNismRmJb8t0fgMkWCaDxBsRQ53hGhR27rbn4PyBWERxRLs1wgo
n60UmuZIfVKs3AwV0IQoVgjiNTXsZZVGO3Pw4k7YJk/f3ryGMKRU+mMBKnEM9Imf
MAkA2MfWpI+89ywpA1waSXRKd0Dl9R++W8ANy8sID8fGxERZ3+QRbYe9hUQdlEev
JSLVkT7bUfhprrfnrlZIUzayd0wgcbsSRPt9DrddIcM6cXI1k/ZsVfDWVDAV4L7C
4fXp7MKzSQ9W4AnoP9of9LeZBYI+/uc9xsEqR+t6dSGH9GzPdBeQtLzD71BAtRfH
PEao/7ZUCYfj/dIMTI68VKTl1HwAS7TNWK+YORQsIyfu5lmFgkhazdlPVMLrSCge
5vQANfLIHL3C7EmisnwimzLds/zKQzj/LvLMcbsrmLbOvw4sehqE0pF1U57SNErA
slXXjN9SmIg6gs13TPIedRt1VE0nySgSqOs03bua2fSaEDASkUGfM/NCE/BWbkcQ
BcXU5mWjQ7LwpVNW/PG33SUorWahYYLNQAsvCfrsJ9DlmxtPEAx1G6ZTrwJoKG6h
OrZFWxaenHyhEuRz/XCC69AgSiaQ/mURWbweX2z3BsK0ng5TrRMkcC0IQuvmQVR9
iDV4b3632LdcfjXq8Q8YpYH0K+CvWqVVAGHZMB6UCiYkgED3fufBea2KzZw4ZFT3
waBrkA1GzM/Z50VMXXJThZ1oLfIDlTGklo5CbHcg+hUrfZnGxWvZ0YHitiTcWbCz
ub1b40RSGvo6mWunFevph4V12MimKrf0PF/a16oq+mrZrGGdcz4G1vpjnUeH5Uzk
0o9xfnMvNSNZ8ASDn9B0SDeGpUfPH5g7gj6GbQ6vpkEIfbQh3Qd28DmvQH4HWtjr
Cs9aGvmSWKmKCFZO9F9vVNTlmXsrAG77H1AveZF1dWrVcjKP6DpdAyWnLcH2gt33
9fxdP4GxVQ9Ky9kg0+jnut4qX5Qp6xJlQNkR1LMi+NUaEvxzWP4XIIwrsTgDSBzS
GOoVsJ6H+wvUzATwu1BviAvAZrvb2NWE3FCA8gJAOOCOSsFfNUixqbDRHZacnFs+
RmdoUnYn/UrkSgR3pQuAGCuZB0prwkxov+VZCc/ZtfHkEf7JJtla+6VvNCx2EPpr
wBJ1XmzYlexmjDGTFr2B5zly/jXk2WU/Li7aDZ6VbqUtkWDh3AY7w98kZJE8SEGr
gykLCS5LVG/1sudisddo9aJ15dz1xRh5K03oVuj6vHrtuLUlcI3WtBNO3EemkDby
wtzSAfRnBKq25iBgqXqjWzEAJECPl+8ZZuURNwmQt8D+jm0e9k315ygA3eVfVlXZ
dEgZxuuZI8YAafcAYGgsMiWqXG5wcbiKnpItBajude5kGP2X/wxLRNHlTdCtBy8Y
OCFoCxEYSSr60F3wlgLspr8+3DxvRQGI5W/IBAGoFwhNtLs1Uty/0C5im5QVi1eZ
mebM6MnSs6B7Um76TptYCfi5qXSo+zYsh5BH1dngmNQXvzWMOaWVjh/WguaKcWj5
9FGF+DFqNntXZBdYDnIo8XWIa9ggnv7t5dkBsoaxCMJF/acmyh3piVMv0LQAm1ll
sn9XZle8WuW7nhz2qpgoTS2+8eKSx59IeIf/xaRgfhaWVZX8DaLFfCt9Z5ew8CAv
w2bA29Dx36qzPIncvGUPYbXu5r2K8nZtoAbZmwssa4cTkBUh6K6DuViYwNvyAoBE
J0iXR98LxVrf15dj16gVjqOyBL0ClLaUFFDst0DrxR4/7M+TvUQXChYqyDvt+03b
E0UMgQt237nXKJoUCX/4yPyRBJnQ43z16hVgIDeEsFUkDFLRTBdzirh+//obXHvD
fnTi4+3sgi9OoVf5AoRJMEe9pxb0qluZIWyP9E5CXFWF468A9jARWkdBpUfR1lYz
GM9Qj5T4kYiqij3sZaXwtvzodu0RQnRIY4C4JcFS8tW2v50loLgIPXrCqu5LZm2/
P5nCilgN1tQpTOAB7LQXKwPti9i0lCZRey3upOtRehCYlt3xkCd6tv5KaMoX4PUT
9zaGhpfKmKOyKW2yPVoHyMYvHI3Y96NYM7QjMgZRySwXDbjmXi/V9Ik4HVTAjnFF
6YwlCMl1vxt+lUE3TkTX7IPMa7bddWa7yLN+L/TtdP4aM0R2GohmPG9vPlKddqxN
0zGPo+mFBubMpfESnJtaI9PNOxD8glBPA91SoQicQVbrFNJNNG04EuQJ2XBkJwTC
rGDdw71zuWU37nPCy/UjgNDh521UyNrSlOHKoaEXAJpLEMxFE1Opn9PHvIoLGT79
OBp4wBRoO140QELqtagkmDHDN6dRI2ECyzmqjKttIMmUXjfRfcvgdbaE3uvURaA8
Nn9d8DyZnO5u84cBTwm13o6yXp0kulz3x9FFYJzEkNNvykWhD6DIn5/t3VRQ6E+4
NDl2+cPvQIVkQcOPOfN8wUvHK9BzUhDWuWxSSYfnmDV36QBJb7sc/yaF6LZ1KdAJ
GZhOTfyDd6/pGuNo9c2vJhI4pAXbxqK2JxAyYBykquwvaxOxfg/IAAw4LO4HwSRE
7L0DJ1tHTsxD82TEyw5JzMmpI7hdw3MgMTdLHpF0uh7HX+yFi9EcD3HhdVyAU/qv
22gZjWtTijOX5fd0GDeomnFNIGR7aS9g0eMs3MIsgIZIsOe8ubnCN/S4vani0UbW
O8MUdlWoRm0lUEg8cpyGgBsnIDEuWn5jmuls2XoVgRIT4w7mhcvMCqfpkscIvR8d
TDk9PjLkXoPiATvrC3R4T5ll44bW9siTuN8gwZZ8aSRziJnNZlO8BfHldI2YztP8
4j2tYW6diW1VYUZ3LtfqNs3kkmv3obgji5HmYekyet9d1/B5mIKaOHKsqDJ90wxC
00fMCF+R0fYBcqjUG76jgtnUF40Htb+c5cuW175tyokMXM6TDG+OQYz88ycmc+DP
RF/379bytEbXVxUHZgDMXCMAmFPZPAIPrPJzx7Y4Q2bcwPc1bqSyrOcwZhLIsDbR
hCOkier6MJO+t1JKb7ECuzUGCkdU6btn1GZNvPMTFAHf1OxJfcTa/Cv7v9LGwGjJ
vXF5vXdrJlVmG3eknjJiFVCmpOQGRUwW2+eTctQRq2zmLag+dEZGMzOjvZZExgWE
4o3LEjiLAKkNkzisEYZwdAHZO11Fir/FjmDcBAR9LY/KKCJY1bbysfEGKKMTEMwG
fSoG6XinUP+LhNn99ZG5SnQDv8lNwAzm1HYvsJZ+fgm/SXCmgno16/DbuLN3poi8
41zTEGEMfsCTfUl1Guzn3+Gh1G+HjJn35FdXWqX1NCczqWevdroceExwfqKxybDB
HXtt7+q+3oUrF9sa6rIF11jKxneBJeFlwXKrOVEmnfaG9EXMECVh3vMGXOx07XSW
4JxLx8a2QnQxY/vjXwRamEiPDDHPBZeNsErEtcInzVuF8v5WzomOdjwkH2rxa/lh
ufVDS2oMBzvM773Qu4Yrmbt793Y8k5xzbKTHr1fadSiXFjYe0ZvmgpVjAILGQARz
YHZLIlfgDUGGZ15iY4GVEurCeNSTDstKE7TXprCoult8/daZVaGssplVTkeZoPvA
EbdOUGoYBin0IoCiXD/g3C3SH5bscGQn9CvDVuPz0Blja6OAfqcfb2ohi8s0kEYH
PytsgXz24oZV9VeszFPrmXB2zwEKVsY4H33qVMk2sArMboInPeieOx7PNOoLdE/v
KkU0Nnw0RRZOF78YdHN3hD5gnZ/C2vrr2pq8PJb4r4Ybn5dgs4df2SsiZycsgB5+
6m1YQOcZ9wlSMV2XRRLEypFfYB3J5v8hmeWKWbV5Fb+bLgeisfX6aFY0aCKLAIxa
OGGWOLIRrqmaQLUoi97dACVzHl5ALSLp45mBP20cy9tt2b3Tme1UQvFbFdmhgAuj
Wp5jWTQ2ouha+utuy0FaVCbbbkT85e4h0fuXI8823ai9foZwUU5YPYQ6VnN9ssT0
Iv/u1JVEs0XcDIi1+DAm1d6NJFqPqmAd1BSOmEXlJKd7g/VMa+6x+WiZWl0E2o0f
2Q2sr5RGnEBdlifJgDHd/ocCyQhMG/tEwFOn8KBvBOORlhfyTGiNthZTzhtkmxEI
n7LDmMvZuDTebRSmpQPF8Arg4hvgBKrzpLqSZK8RfUG0CMPTdoEk0KR/p+RmRCRa
Sg4bh+cLfjJsLaATwqsM3GPLCvjVlx1nlVr8Yu3q8wx6F1lsh43arjuSZCj9HrLy
67DCnSYU4EG0D/FvGvbjrZovcayDCdQn+tmm0DZWkBoYlA/nfz1XfasRc4/kM13Q
68Gcs5gMO0EGhwmfSPfGpEd2gCA58aVAqKg4nwVYbXLSLUrgOmO54Ft6D7nUurSo
x+iHbEM1v67iRJilF3dljlUDCsy8UnQoiamkU/kthgVjE4Zc8fArGR+QPNlCUgeU
fcO7kajxHwW9UQN4t+MRk2TMryMAG1apWZIYbRFCx5Yui7vNwkbFW9WANHjhI60+
G1lQ/rK9UCuLV3U3VywchZYL8etVsgEKqEL59WkgcEznS2ms74TjdDdwy1MA/+z3
3LJq8RrKm8HmCsEVGoq+A4YmYeJhqLEfwsntCGMLdmnHKv66f71GSM7CUiuJN+xT
cjlqBxh5cs/W7IZMQuve1bolkNo3f2YPWO+4IxPQEtcJIVFrqqQ/UJQv9GTHF5i2
UfsvcMkW11ZTekHGir2J4rW53h5ptNGZ9AZYShP5IO6B4XfM6OUCl8DrB5kjnXkE
eEQ/HtVAVycIHYUZvULeQyk9PsRRRMqhTMfvo+MwvnIToKEXs4dDjw2gOqQwh1E4
qgOQArepSJrWSFy9ChxPtI9KEO7EVw34IXZ6OsYkf2a/tfx93+TltoU6AThGhSzc
eT2GArwbUftWx4TOfx/R/rhrb552Z7huP96gI2JAu2lnKD/UEZf43J/1Hwn0CH2N
BdLlqA/ixVQvyWAXe8k+t2XI6UjG4UywQCzS/b3xLA0oEt6kqGK/aA6DZITBI0Ih
9ziPy1JBYa0b6/jcWyQgzCvXbzc/ihHglCxjKxspBPMfjjGGblz+1A3uGRSaN8UE
QMzA3tkwkOCG1iT+qXux0S24aI5QpG2EC8R0FPWGxKOzVZ6sfJl4jVMzBvWiv1nK
eQ7SLsxKkFukYYw3mEef8SqtB1iwdds72r4LPGtHDTFzeMi0klnVpnNlvlTfudnC
ww4C6cJ5yFQ6fCeo+sS1DQq6stzpzHZ5JNux8YKa9sloXD7duqs5VrWygiyJKWnc
ZaXwnYJr9dxidp+YE5meApDLPzuT9Qkq8Cl+VG1CHSHr9XTrWPZwef95lVBBpqzT
wQRi8am/7iJ93Eu94xPkvZh6lR6SxTz1MnwE+KV2qwtF0lQS5U3VoDds97SiEuRg
W8HpjQRNitP+O5QnlQAKMQHKg0aXfCsic+yjcahXnopqGG1NmvDeGJ3+Q8tQrEjh
NWkzeCaEdo1BR7AO4/B3sg+vH2ZkHQ0b2fIygtYqgHDjnSGKokn1rouNVO+ZcJqg
Ah9t0/jjTotXNXj8Z0f8ZKE0y3/raE3tDLqUi0nb7y3+0FiViQzi+4xp7mp32mcy
OEhZUGS0TREAsPrUMUASfIa5HUkGFCZG4bpel7jzC5HNSGv6XYwHlE68ewzZpgc6
G0MyyJ/D4MQcsnhz/+o7dLoJkWsmlHR0zAS4VUFtSHLh6RNRIsqoRkh/wysPtLMA
CTsQxXMg7W1ilHjC2XEvSsMNf9u+ReEiUSmxckUgisvFdJeKBpCjVl8JKGJsP3w0
Q6BpJ0B0IClK7SfdTzJRKACsu3s7lbn7wrlRPRkihYxJabE78GPcjGp2INyfi2gY
QY/4QoCxSzkEzrHT09bM7V2VeaxUu3stjruOG8iP07Br2xKsXo57UKaWNKa4GsSk
73x0IOo0VtZzAzgnQnOdem3BREiavErq8Qqty4QAcBoHxJV/I7Ch3Tk/pq/hFsQE
4crnvwfjPqBXHna1w7YZNYADSgSAEJsE53/UhD9OeBV77P0MSIyCrbj+yHajxvKM
0hkEBhCC2Dl7vuJu8i2r3fgCyM6eeD7scYP+LX4Fyg2ivPE5KFrC/bHowrVJ4geE
ETqL14iaEZxzKyjELqATjJB700Qx/hoaomsM08eE8Y8NoRBszr+f1AXoRt2qaKGM
TBJ17Kl22zKEQ9izoZ7slqqp8rCd8lk6819AHsfTuzMkyEhHuszjdqBzGAfiBSb5
mUvJz61ccvR0TppWiT6gq91D4ZxW1AWSg5XaDFu4A0/olNd06uZ9MUw2wr5H1Uqq
dJBB6+CeWDX381CgK1U85vZ3ro1PlAwUhmXX43dceutwstCFerPSNUwz8z0nW4Oz
2S+Ssxu7M65zejZoRH2YRpoWt1EXFhdSTHv4cYacmLCglyeeNxG/iw/9drSba5xQ
bexNiyCjwXektHUIC0v1Uf/z8In4RDzsg5tqLkC0gNAZmQaoX7Xe2zfbQ3vUm0Ju
rAMMKkyUKc6ssWFbpNHzqraiu6+496XZqknhpKFIq9oh7XpKDzd6RqlFxa8st30z
PqdxIw5UNcfqvudqpidiJNP1OPfCdhCUm3HAnMWgNUd0sbTNNHQ0E5VxZlojKysD
B2Wmjg5m8AHzWO5lk41BjVEBn2jcO8jDninmMuOt1e1WO9kh5HCJRHk3ca001qWx
eJDYyIzIkwkq//30gjLrpUfb3RPcbn1v6UoemMMvxMne1o7BtZtOAuUDOsaOj43v
Pc7RbquuV1vrDMGnUpsOAGd5e13j2S/d5Oeqo9AuNqp9qBkqUeJAtGS+fQDVSA8t
eVcuVGUp1wv2qEx4LVXFLqdV5kirpxO41XTWsi4p5xDM0K8UgdNEGlBaZMX6ONxW
x9D/RQH1/bpvkEebZLMwDs7ccc8BuJM0Cr+EwN7H8Rt7zCzk/VZw0ppWPeWOyTo8
/Pz/TNB2jTXh8DE+xV1RzZ8henvh7dBJshKyjO78N5lmwyqct8M7onaYbdIsS4qg
6WynXlmvHvE1p9xoRQT4H/g4alv5kfmJsN89lM3iDp1iZEFYzcsx3zeRV5AnHtfa
NpobgbNNPEeQi6iv51/LMwevGdEgYAYe8lLeXBnFkMt5aC4mVLyw7VrPO4fPIVFn
1r+0uoKBRBDdDMpogB1cHlLEYS2uclfq/u6w7TYl8A2hxnIsLSn6pXGxuMu9sl+P
aU5Rz+++NrZoI98vCjhY+vSJ3BQYtsmW/8s9pNZv0rY79iVQ3dBVL0UYArlVQVb1
u+GW2Yn+tUSLRjGwINpEaeTDPWIBHJLimjUeoNhZmEOKaleRE9xheihdACvYX6j0
UVwYLivFlm+f5wsefBVfdMayU4zAyzSTVlplet52Ud0zo5U8OdRoBae+1wym/ZlT
O0R0IEVecaFl5K1d9JZjMIGukW3jmeXP9aLuUKfn7Udyq/uVGdo8g3AwSr6dDsYu
Cv6TPXXP1znmAJmIJts9DzRBqrhwrOeD3lvETDH73qg23hzgU5E1KX91A9OqdmUI
hdcvgakblnr6PQZDM794+LT/ZJ5uBZ88h//BjzPGyObF74ZvqCvEMnr9TfFVwILO
OfaJ+u1voZ+jhEfrx2b0qPU/nZ36bD37fkyIdR4O6jjZFHjReZEXbIgzByWvQyWs
8oh9gWvVcEVxEnD+Fsq66Uh5hfbyHG4DG7z4xkKl45IPkc7FgKNr9zDdGVuir+m1
ibaDBO9WB27Y3/K+BXhBBQ7kyW0NSS3cRwfRhSZeH0QpZqZzR2HprsKguH6SsCcZ
fup1w34Dp7HMNeIKFutUoSVYIhlm3Zhid+/K6a0nXSuQlkdmk5eg2eiK86kRoBy/
OrYdGqEI9TEh5gRCgxg+P4+vFJ78qDWi7rgf3SVeOB5rncFSrQp6L0v38ZRXgCsK
lJxWvBr/44Hq6iKeUf22pQLQEmWKpraK+xRuSua3DBnLCEU4gK8SqPMgpTlSWjjU
z2cyZP/RPZJvG+vLyid0Vf2/RRa8GsWfznNXYojjcmuf82eOd6QNXZaK4XyVmoQX
st5wRLTraW1mGAepYy2qCdtl06pWsHKogHj2S62tB9sWKBAEb2pZ6bQhFEECPvIZ
28FIE3vZif8u6cEYWJp1RChf6RkALTg/0h4bqylFyAXbK5CEginE8qXtC8qKRUmL
KQ4hls5utTkmxsoE1aAxHxjw1H0OtBD0jwgqsCgcCbIOOycsA3FID8zdg5Y+YIp+
/2r4S7L/HuXIMiboBnlWi1CU1m4Q4GB5kpssJrwrON2JzKPZ7Ctpu8e/H/AiH+Lz
7v7VXK4fCKaBQKy6WKcS7Sgcni6jzH6NuY6MY0jD6BICrtmzlYkQgju+WBjR5zEW
oD/ZG5SnrvIi1Qg3DTVP/7nGpz3dx3DTslRkHseCQMf2NtpXfgmIgoHlV4KgVril
wbN0p5o/L0mIMn0vzl4aOGlaGUdDhmp5ltl2Q3zhEK9wRXIAS1BOk+mN3ixHA1I6
ZgP1FHGPvFHqKgPx9bGEFDzwK91QuCKJ8qwexuBje4lkAkg3SQX40M6DJ7TliEpa
ZhKsUr7Xt8LFt20vHfkEvyKChaYEs3/EnXr0sqaEBwvSkaZR+Bq8dF7WS6MvVlNV
cDxE55ZImQ/9nZYBwmra+uSLZyzqVOPriPiqk33XNGD7ti7WP63y0eBnlsNtmVrO
so1sbBtO33bJI60ImK03+Yz82S991Z+J5cbJ/ysSP5HmqCMEXp6f/zdOMVq1iwaT
EWW1QpZU5rIhrFIDWFgGTyc+yNfW3gTQa3kZlARV4l4oZjZpAFqQdus42K3wc3CB
LRbmk3lsI2e+qf4uH4N/UL52Dp8KudT4xbTkMyOjJjDXw13633pvo29eVbpBlqd2
Kv/PG4sDL3n16bgqktkYXfS7gtTHw9nYwlExyGsgSwliPNhorR66TzXAMKPeCFJH
l6CP4E7mbrzPP+nXpDtFYS8lx4mnNUXPYg16qJ0SaNj2DB2mmkdF92MoitLVVtSt
Cz1NjSCjoj5WOJAbVS13JjREVcF0+pz2/MHBnl99GV3vW11xyzLvWa9gRx0QHda7
/OqnZ8iwiQp3pYmClQbRZRyzdZ8bYXk866ZOd/serbIdbiwaKthXIvEqOtY215FV
lCuRSErUUZEPp4KV9aUhHQvOHmUyoQhbwGTjEZBdlR4pzuc/fEkiVFgjhWiRY+W6
KjU5Oppm+8mKwW9xl36CNpMzkoaPwdRAB6pLe2XnVEwRu7X8rJW7obvWRIRZU4SK
0FGoJf5/G9tjtXk46RR3qHYAZAQOLjoqB8yVagofERxqSP2n1f58kkKKVSakCZ7G
E4e8/V+8XKBD6WDVR5G+a7fWprjP3mLFBwEFYreEFPJ/0lyEElBs0jKD1TwK2UcS
vaW7c4nQf13EcR7F82/xI2d8AGfR/yDMs2X6zm4mtaQtQJDhcI/eZ1iNScIceG8K
BdZXQOdrXrlvZabNllD1AphHFWuHPHwwMNjdd9jPXwJxhRHv0/PDP4//JtThK2GZ
YkXzwnDaxZaFlE65KVNq8xlaq/NCWV4O5EUboQC/Flrmd1etGGYZ5ZQW8bpWZJ+H
+QYO66j8cm/tE5ajP5flC0kuFxHqeFhGJ/pcKNsslVyN6CwOrCYng9rYeTbOj/0n
4+AnRtM8tZl3V2gIExGjOMpGyiHfaZHyMceYLrSXQCkQZ45wPe3F/0Vm2+1f1Enl
gzlOKfNQ1t/AsIsAuoqHL3Xr4KmzZ8Z6X8AXNw3QYY431/fK6NOJhYspgxQy9eXX
bqRVigd/D9RGw22Grfm8oOQpwhZc5D2oDVOOwEiPuTifYHTrl1otDWhit5uhmV4V
1S2+Ej8g3Ow0JNoYBMO5dxbUWVTHqJmWq+1ZzZK4H3Ch1FdYKaWs+/OQAecDQxFc
OBXjDpuD002HmFGrot5O/lqobpkiaY6dfUlK01Rd8az7V2QV9wD8IXK5UBHCrkSS
CUIOjrqAwUZCoksIwBh/zErfIMijiSC2FT26vr1duK61Gm2abzvaAuqDr6CUTD0T
pdvkF8gw+uidyVJtb7kf97ofaOaxPEFZqdHhkZooKsFTW7TPM82p29xVZfOZgsDF
qVL2eR3+x4FiXckWnsPXXwQXJqLkAtpNSfJNm+2SYyiiXandMlFRNnlzmTdklIOY
HIiD+BLu3IP3F+wX6/me8p7c5wTxs8iwnZwgJEFKMnBaWzRgwCA+P0suDNDhb8zy
7hm3dQ7g9sTnEJu9sSmg7Ib29R6jO/e0RSzrRNUu28cAR3XGwTAiOhqU/OcBZNkw
cBRzOAvQvYAqcOZpeCJRMhf4fUoLniqWvAzRXlz2G+9vzq0twjyeFFNrTvCK+/9s
3jkqVTkx9flJLouSJiIdr1QX89QpbR9h6s7gjG/Ppt9bbGB671nvHYSikdyJTvFT
wIUIvAxoIHf9Mj0/L7HTId9beenDxk8g8rg7bdshojYxJ1outhb5ktlaMtB0X9v3
i0+OMsUdTQ9v7ifP0OX/LmR53TxVephBH6WdDeusM/b3tmjmR96HF1eYl+2+1CN8
17DW+HU7xXF8CJ6/WH5n6i+XZ8Zcs/mzHscfu8JAYsSCL5buQRoQto7/cldnMf+t
/+KbeMsKTQZ/m5JkZcsBg35+WJHC/TKcmGQTAEDREcdUd9SKsa5GL9Oo6w+XAjIw
YMoq6dwPBkgZgGPp/LWBi0VuSpzKWTYyVuVZs4xs5a4t+WrAiUjhnzovBcRRqQPP
kJGWXlqKGQc39E/KBHIVHKmVcdkXBA2uXBITXXG9hvvuOkv8euQPCB1GCcctB6Ao
DYCAL/xSX0mTvXsfXgWiCLQDU712pojpw7bvwIolXFwBrotf70ApcMxEJisyoXjP
BpG0ze+k9rHzNFOlq7PSz2vAN87ccxryJxJTqHs1A9C9qo3ZyJRqfFgWrotTumSD
WqB0dlhwVyfPvEmZK75Ryxpe8EZOLvli3TKuf/vfcTBIAwWvvfKNrynsWHKWu9BG
z3iY9Bu/2PCzokkMQExzm6sm0wRjkuaTJ/iNweKGZ9X3GfxKcwxRSw9IYLgXX/sD
RKGGv8tjFS7vOsOYzOET9Ny2F4LRl3Bl42Hmu3FVfdQW9nMMgUeVDUbDpdZcSnOb
xS235fcoFwzli56NLhv4MtlaFN/B8JsKqlLcSMMhSlOn28aSCQ81vpXseVA74sl6
c0vwhfbbv69rTIkTIIm41tufq3Aimz8BW1wIf/uwsOAi6LyAHaRII8DXHj1a7zJa
Q2m3mh3X/KDw7jUOCqjO+/vp+D9IlAAujwmOCRlgjDqgBvNPJ5134W56uUcUkXh4
7tx6U6mF/I54JmqqQn9zF9QULEqNo/NnXx6nguPqakXzf5OzBzCCEaEQA3jXZOPy
ddn49GqKKFw+3EuXClKA1hgJ0qwVF0tRCPT8SJchEt4nEEHQqz9Zn6GKQInNuwz7
pW4J0ObkrC8xG6u+dajIDIeJyOB2iwytZrd8TbE88BCKHXG3y3LJ7lcHe3ie3MXS
wrOXnMuaLvB+Indh7Vif5wYCX0tsK2+DNc/NgL6XJL1Koe508ApV/u8o8zO05xjq
VsCnaHX/Y6d2cuAiKuqNV+gM6r5nTUPU8xo/WUuE/DT/Tcke8oBBThOS/58EpT2C
8LEyXjVgVTuY8Tsq2BAidrlDveN+DDBOw2EnHZNVDpeGOe9pqRRa3byIIWLF9ejT
DHAcZ6b6AIcmk6lTOrwdOqINUN3SxkW5FYwse5abwH6VCm+bHh/FpD8UT3bZayQY
RUc8L+aZ40zAnvyqd7HXq31EttcuZya/7kWrz4+LDpvzRXdKc2me0J0Mj8czw++G
vMHjJB6rC1wDIBWHcD7LlKgGx4ARTAwwuujAzbuQ1WN3gFCeT4QpkBmLvQs+XLnV
PL4+glOFZ4onNDfzziJdr/WsnlvT4V0cSieI+Jgxi7CkRBJxWqocosXCGcGdIhyp
YGcXHR/8wRjRe6OAEwCSkqSDtvkre5UxbP5FdRxEO1LasxgIO85LGrhpIilInrNS
/VoEcOU3YIqfqtO1shqAkSXY2boznfrhtK6OMhmpaOHtnTY0rpZuFHn5SRaaMr6S
SqqValqjY6zFrzLurYWw6CwlIi4N6EjEb5ypFeMaGTiqwyIGexkIbIar+7va4SWn
P1UN6ukWpY2aj9ilzvNfMphaWVD+WmJy8hz8FzrHBTtqdINbCvf55sAO9PAUHms2
xIWFyqqtM91SNrMFsQsexryrnux4l8iiGGNTsXMuk1EPXmOPlNfOhHeG0X7K/Fti
GenvM/xUE5wXTTXLj+FuCVcDDXYkAjO3/2fV+gvleVrj5kL680WD/Qspyma4jHqd
5yBy1+Yu7TgWO7xyXex5WCp8wI+Ji0mAwImiqZCL0eG2bx8xfO/NH38orHK0LSGK
P2siI+ARQAizy6rS1P+xP3YQSaquXNk8K3erXbFSeWHwUtsS4SxxkMev8WkexH23
TzAXjaPtr8sb7xWufJsWe7MHV4rWnWNzia8+d95E680ACQ1XrwJOgFnGHYRD5kUZ
oFLqVzPMACOMwSwMT/7RMfkZQpHOyXhWVC1rHvkVXYb7Jnv19QKpkPqXQpkuZeeE
0QCLnLv0HmDvHSxzrOTe3WZnM5qJsMtbnMXOsRcRkFjAXoiUtzUov3tFP/+AaQa9
KyvdSHhx+yJ1Gm+5SqCRXWjZENm4Cp/7yEJtPPIRYJpHSzv5Svw/TgTNlDODgMAj
xg8mSHevI1Qe+BF5FjWnQSFpGPOJ0fKkIdVJWNUbbBC1R8a7hTetb6JxmxPl+FYP
m/qHyMn3uv3E3bAhmN4uuEB4lWpAxtRaPgv82tTVnFtUzy1OmQ9a9bwtCX9ZsKo9
IfqLGc/fDLMvEOeIzXvSpibIER9e+EyOVsLJ3sWFmcTNZYghysXu5rq0XFQUH3jb
v7Tj5je/JB+iUY1ZpCmqHITtPKjUufIU2JtQVNNqQEQsNHUoK50S4xCVeQGFWPf6
Ip7WMvIUbd8f7xUMS89L2JBnu3Y3ZAB4L6O5JBuKdbqZNbla+N4XDD7KBq8a4qBn
Fb7/P4W47FAH9dgfjy1VCSzyA35vJyzTsRbt2XlYUiNO2kdrkDo2cA8Mp3h25vd5
6rbRlk1GUN16k+kIonb2Y/+7yzMaWLvvFhwXJcEtZHGrvxL2CA/HTOdF4yer4iML
zbhNm5Jd3mAK36W7g1sodrG0jLFVc1WCO+OnpCqtZrFGNRI1dZcosKhEIya/bB4A
U/v0OInuuNfTW9X4Sl5y7nIROCdQq8jHulaulS8rRl/cDERQxGRsjWajzCtrEnw5
BEQVUxVwu9DH1BcHn1NBKG9Vby3MSqw+QZRMY+ZNWN3pS8J5dPcw8Gw43iUID856
G4tvxfePg0r8cppW37j08LijBqA91Y9vWqbSiynQW+5MAPaCt95o9P9ygVlJu1OA
wFhmg0OkNOYKRPIxM+/42Cz8Cu+GtFhVZWhWZOvO6U1gQn/OFt1IY3U8FtG0znK8
k4jCkkEODa/Io66THv47a3/84pgM+E+vwHCryL5/9s/Zjrb/q8pm0XxkrsyTzEUx
viKgz9dIvggt7mhq2xMhXJWuuc0yQAmJVzfaICV8o7sjiwso//+olxAJ08u8nIQj
nzI2gAkuhcgAct4/rIbm8JPDRIujBYedUuI9RFwN70YHnap02AX9TTKsRS7teyaz
CbZGWHeBCRmwrljG99REiwJHcCZonFgJVHLDY48Eqxa31bUjmz9kRZOgxqv5aqzf
XDBWhB/AgWgN7aHIbIbPgZ85doMWOnyDDrfGSHQbdbJNnKvTPRZ//trrqNf2e5ZD
rBKYF0y3ttMoG/Mv5TuftyyHotDotSssfqCmv/aM/OeSrwbEaCKcSjBaIPNwV0ke
8nYgqSZHlbRlfPquW2efkf9H2TkHfnuTv1xrEmU14jGa5STAQHPn79Hc/mBAbrx+
W59tUCAOMx9Eo9XLvqGu7TskS2TWLzyyB/H6qU5/amKEgH4J2q2Vtby46aZGD+kx
umcM/yHrrkMecyWAaTt/qDGWmRUUVdSTlogd959QvDYBdxwKshQYFJP/KNfBgTgk
CVZLTQ/s9U1ik1ukmqb9iIK1KUV85vMIiHfS74MZIzmCYpmmZyctNjIQwGf840Yq
lc1uiWns0kOQZA0RB3SNFS08+lqUYYCM0ZsnwGOvvi4uubh3wa8ogiHjR913X3rS
T0LHbsKHtnw5bcduGxzrDcix8gH3vLanBNwUwBR0JgBkAnnGJPKgUYwWsXuQKpLb
bM8X/bZTgJvmNyyJgC/yqpvg65+oeVNUFbu43IFFe8iHZEBGEfT1Z4PINO5/Nkd4
AieyCG8LqGmeXKQSwFHQyZfixakE0MfofEmiEU+Af0jp7f7cSAd7MM9y76shYrN5
0aL9QxNd8OsLzNMNq0nEB2U6sRg7/wya9hetFOD8Jq75LU+FWXTCBjlwjb+0xRXn
WFvbL3r5yzq4py6oqU0G/CwbZNGzfsjyRnF2BmNQ7cXh1Lhx0iOTfwz3brX948rn
oG7+tYUcUGmzEE1CoLQA6F8KrwJnqa0AN539K9/HsC5cBWscxb9AO9JHKAglE1lR
K/2iKf9V9KwK39YGiwFFfWMJOPGbKYw0kLRgL48Dp7VgYipfgkFUhTWUSvviKi+l
fWa8HikKVio6infZwYmCOc0TR4RT2YgFCZQwgY856Zk3TjpgRsd7L2kPiEkOiCct
XtzjepQQx/YS7eOUglQ5bP+91CahfJUKXvOApNVKeeTu0s/lNi8dQWMWiW5/fEfr
y3YuKYXjTM71SEkr3Zdp9/RhsXNHzk4nyH8LtpEEvHAvOIlbetRuMq77VEX8l3rV
TxtumOJMWXei2xrHSDcqo26vo4dMSRypGC3OFtQbjkD20WSMO3wsvpavy3xQCkPc
S2S6ddKueTfHXL6OgrMBXwA1dsL/If12ucVIfHGCMQfJHVgzX+cZnB+CVoJTMHR5
B2aVpdDi0JwTeW/5WYPdOk8ahp/+sfDl559mwFlJoLwv2G17nyH20BKSaUMpW7NP
dfyXd4htfV4/kNejug2dxPnnc+H3NT6En4dkGMDHNsqO8eCbyoi6rkzJt9geMiVB
uWeZGY1EfwJ191rQrDoiSlGcjtETzXcrsjI10Ye8yetmKxy1DG8wLVEJpA0yX9rw
37/0Wo7zd9jGM6BxzUWD4SxGDvMkW5OkRVf1r1XaveeLIwoU4yHQ0rjXG6sa7DQA
MkdWsNIZRvMoXAY3VrrotpepTcgsqwfX/PLmjdWHNkeKzPK3sKTluPpnPeKt6xdk
gluSs8olLv/CTB5N3wzW15dTOdSkEoaGU9BG0hrnZ4zjttbnbUVSG1GIUOlSY1hD
TkcrplpXTj5V5zQj3a/ojOTQojJVLptOzrRVXAPnbsfVPK6aN0rJoOC78bDnNAcc
3dO3aPuuFPrH+7wcsyX6a82mDuB0u/KTrvEuqegBi8W5DRzUrOKcaMyHrcar0Sdy
v50v/oIxt6f8jDlC+13qwdgsXAmaIYle6KtmUf8qj2IIX7m8rHhIXdY3yHSy3t9k
yLBTxG1ODH3ze69honzZfiNHD0RNfSYxEQ6X/DwnS8s7cg7GdpmvtaaRkBXEm1LR
VQx6psOTVgpOzCDxYuJJt4mF0LTBuPTGfJnoXU12k5sxjvzAt0ogmkUTeKJbPlqU
H71e9BH/KrK7u3xlfs+26pbUBeWYi9FWHVXSQ+Q5i2cOezuxUFn45cAqqpDMLl4G
MMXbkainiaiJr0OOAuyfmAYnabNkzmlGhPAOisPVNkiqxyjoUi+o3LE8Dag2tzak
1dhkGKSj9HkYs2uOInBEUAh/cQs0byDzDY3ZrgXB6ktCNzUZeWwh1qD1fBsjDJZN
95Z6JUEQaXAuqKw2yu3Suk6xHDcpJp+Cb3kXDvzCTSl6lr15fiCd+iAaZFNg/+bQ
oCVKJt7mBsGqYvadtOXF7Vb2eJGrVZ/21nsBu4gXoxJT+xEYkp0pEjVZP8gq/7wM
F+v+hPyOy+NeIREJXbXz1cDCKZuzByQjbE4t1K6WZyFLlQOfoSJMoOYOJxHxtlNE
ifT7nGN4irU9kJ+J4Nje1/h12ciq5UJipcG/Sfonr9IBeRqveWq+Wmd68VXn4cZM
FLQbzZGmtV16izZAfCMzCiLsxp7mcjDgbD2gAweLau/Nxe3CywEwKhNCNSwImPl8
DeB1TCk2xQWRT/GA8d8z/fO3A6xt3fjYkZKbzhgCdwV/y/Ru0bbLC1s0Ct4gV2EF
aYbo0x9i7dFTEuQ7b70Y/HGoZxa5EuQQ4WXd1a3VfPTdAM2ZcwgamN96fVmpk6sT
fHmAB8cyop/+XI7cZXt3E4V6nbrXM0/U6VXvL8EsFo8U63g9NKZVexjmYtf8AidM
WKXzpZvuGq50ZbLvFX+I295o1XwVTjgpBEkt0dGGFcTGaUHIE0s0bwGbdzqeSHcA
3DRuCyuZHuZPJ58DvswaSG309Ch0uwd6SL8lK3GkPvmDeuK1yrcvmuoDXnTCWcHT
apM0hww9+zHa0N3t0bP1deraqbUFAuFWTH/ecumltvm3B5cUsPabTlWZFG1rPyQb
4S/mWVtPFuN/+eOj4bpKfamTXkWPmbdUF6MrHWZckYMLfXaiba21pHEk+Cjfgj45
68T7ZGzro82xiysSHJXEn4eCVjku/QP2CZkr9lIyWKXexnFi8u2JujlTMFGbITTS
hBHlPWnOOBgxxZA+Rk0M2wLqKGM1aLlYUkk+FyUIKOmYRS9cOpYld4BY7dN/9BNX
3ezSTaMs9H4GJtCmaEw9CDJ3WnhQNz1HmbGL+3jrbLbF9RTzEmmIsB5gmCnvnmPD
oF41Jgr5/M0hB6f+1ExyPKcj3fg0gpAWGl+sVuE2is0YyDS7vALDSibxBP6iwGmA
/6I6bPgQPW3ZVfs4xf5LCibvjlHIvgH4sZjU4rKRayV5LXfnGMsOdg2zjg3PQJ2T
fdhfDHlmVtn4DfiDu1QHld2Ub51l1ZvwpRL1zGA6Xjz/zPO/Oyj++mbouiNHAOrX
yjEsnp9H/vTxEw5YM639x9S2kw4xqe70CIDBeSZ9bm5rCQXPSrs9F0pwl+dePt5w
p7Y43xdz/V5GZoCIKhG6Opo69hsFvyiNgn90yV6nRSioMSJo5lw+CjOrdEJfl/qK
+gjP0WVlMRnpqQ7Wqmc7cXK3GVb4cRHFxjc10p8nABdjMIoNGw9ITGp1PByWyidk
lBznxacoYXrvywTAAowbK8GmjwTdC5PYOku87ToDteud1/Eay+jrOFDLvsZAl94R
ClQ6tSgdtfATlcd5f36Z71ESouO6HkXdrZZwvmZxOKX0U+XRNxzp7BjaL5IZYnKW
KKNbLFcWDPEQTDLaxryJ2R/qiTNVhX8wG+mryUlQWb1J7aB6RngEBW8b2N3LJqMI
D/3w2C6HRRlCnZbJXWS0RgzjhctOBvQoYxNwzsD3lPittNrkRfxlNpaGJ274DFkq
9M7mF2hyb7fR2kzWkzp24OEMQGLVFj9K8udy+pEE29CHrPIqX345Oi4GkSrX6Jtf
3ohjx0a2xZyPxuQxPlQLIymZiEe1D5UM/FbXLLnPiTsLAfo8eHIldBJNtTV+NXqu
uEpka+xPKVHQEegY0EpBPKpWobEUBOcfiG/ZoqKnF7Jp8QFFCwrcghC1hH3iOB9/
5NptdOttXbM9RV0gONNkKkMkNR+/bgrHYnbGUizyzf9Yih4yFE6Vren1GMl2CyLE
7yag0Ez+xU8/zWncBfH75ZNDBp5NEM2RNeteI/SbNzlKGUNhKgrajq+9JQ76L5w7
JNXC6QwIiK+v+4AGHeJdroNO36Eq0uFAP/2h7/eLpLPFklQYo3HltaA221xAo7x8
HS0f7QgVo68/nEMyokxbf1/ZsvSiJ9y3ScTvZHoa47UVx3aC6XNSEiXngjG1BC6q
2Xf/k1ZPrQUc9ehjKV9aLeJEp+oYDAWbUwB0T4TGXIRjaTEI9AodUhrsEzYzuBA7
L6Eu+Is5Z2F6p7H3BEQRUbEiMccVqH2J2wodIlJ64DlolP9SFW1Ljjh2SSI1K7nV
dIvhkonMIvbqyy91by1+k020SnX2BU2+rJzE5Wn/C8M+eoC68krPTPQmOLZMhPwd
OQ2wa+vujfavL9g/HYYfH0U8q7BkVCwyGG17uH3M7SDNd3mXjnAKqyRSft8OC/3z
0jxO0Jkt7ayk5Uy7EaGPjUztYAr0oh8J5YObXBB4Nfa+baCDBzjoaiKKBas0hnvY
qYfTJdBkr3wzXvZiEdctGeRYCWpKLQEz/eHV2YVyrGsOG4UiaNEL09bX5XfGPL8U
UKCAvgs3tTZIn85GRrQoSRORHakFAtYh59XMCD+3k9u85RTSZKuXvVV24Pdny4h3
EJyFJFlFa4yYQ+Qw7r0XFDBLKuk8bUI7wLJGyvd34Aq/ecPiR+wZM86AebDZkfAj
pCsqF/I+U5Kwbesjl9nk+ZNupjLIsltIuHBgJCa63KHt8CKwRxAyGh3h1zt6ETAr
EC1psZ6gk31Sar454S+CNHwcXP3aybtqQF9j2QEd+nx1dh90sWQwu31YOW87moXD
PWMDBiJzuf2MycF7e8HSJ0ktk932YYPFuiPn813UiSwPRm92Xi3wlFP8Vt3yxgsS
SRjeAbwRvAAzxV1Ypdwsj/lfR4Q3QNsmNvqbtx/R+lp5Ksm0SzTiUcegk0OpuXcS
EGnLTp/EKR7T/l/SIxroVoYkOpmsLLQ2ozdH/Agi7tk+7CJGdofcKUZPcGDbdrnO
c5knq/3iqP71A01omzzNJ37WGjthEuc4x7HpBh8FNAZEq0MrpjmFzl3f7Aeecgtk
G5ZMYuQX4S8+niG1MgwXTKsbLsb+pUHtCbObR2dXn/uP4RWj0xLgMpImpSOWNRLW
FqSQZ5kSN7GqEDVb9xEQIzVbMCj1Aj1qEw1qBQR8Vl4q4jHYyGBW64AMmW8xikYm
zhw5RPTciAsB8mhptJAucqt5mUJ5p5VcFNlPFUkTt3NNsK4PJxcRTv8eTjoZBwl3
ksMgcf0kUjPLvnS7lTEhG4v+K6gNW0acZeSDJU7TOeFuct+4ZX3WFwOtw3LOqCv7
3Rwoe1C8PcX2zatxDI4MEb+gZ6u0zfZqvBpGizVrisDMH0+Fs9QPZr2lHgvRsZN2
lny1g8+J4l4mgbxiz35qt9c/q573/KIDXakruV99kn0tU9K9X7HQLrs7YaDsZBgW
f3sUH2ZCpiO0bBO0HJ80j8l9iA7kvTgUMqMTLJm3JADvfzxljcPuLAmr9lD2Q9fQ
s+v3rD5QlAGWwNU+Fxz6LXaYpHRrCV/h560jD3VMiBGq1Z7p2cXl158azKUDJu+F
2q+rW0Wyew1rZJ4wl2J5kzq7CEFZDrwvG6Ertaeshq70i9Qdvme1DSPybpAOjrG7
8jWrVNGTqkTvyxgmegUYpb0onzKSgfGwxlCb6SwBw93WcACvVs5bK85g+kC8+GX1
KxnH2EkORX2gKgC102i915vj/BY2H74Zd6LOIOqmhEBPHTPJjRKDXH8c3gAU/PoJ
Szm0Aejfq0fUGV/GDASSx0IcI9MyPhHUprmpAW38siBBEyBOzDHZSxb9Y2jJLJzW
WjVhg4og4T5xoZaYBHN3CDF6agx0NiBTlDOWcSggCjKHujhOOkl5m6FppwB6F+yb
IaJS/iNeAmQwUrYqcWanTMhtpAeecse8V2u621GoLUFlt/7r5eDmO1JrqdD/uP4L
NxSOTOAj4DPTAt501ul3cgVNkyvIiYuLUBSxtOoSvsQyK6+veVnw6O/0Mu3CH+tC
Ql+/Uioyg1OxjXjf4mAIuw+ja9iBwjA/dnPe8Xf6Uiyx9e/t+39CPBSDrAkSzgaY
uill/g7gvSOkGEUEH7DfeJS2QRR/P84YN8yQ6xB1bl902VeoPRs55+jM2ShipmdY
qd1EJVEfqlhYcg7g3gl8OF17AzRlXDoW/Y4mv0lAKvpNbFBuiFcvobYodZ4GdE95
5BDtPIVnOpljKkH8W+a/JymBursr1hBBaHosrkaDQFDAgY3nFtZfj866lslnRzzq
P0Li6+LIIbn5ECDTOX7m+0FxCLQSQGMVQ5Ma6KDM9GXuhoWS2cUlp3ukNLOBsrGS
PYh0RWL0TDzo97WPZIBJ84ucVqLGCxQupm7473pfmu9hQmvBl6BmL4sNNdrFLt1i
DhMucq34tOH7Mu/5PzG20lu76wmQPhzpUPcb1YXRlyofEpFUjbJXRP9nHvzUg+iZ
YqoYlDU7BhXMAK4YPvs5TK/Bw6Kel+53kcuPqIXTpBcJ3GE210ryXzarzHSVJ6Tl
ye9gWaSAbOl+rRxix6VY3h4HwnkwBYwnFujLd/uYQRQxOy/mnHg5SRYXW8WDo1+O
LBzGu6aN2O7a5KIWt/9c4+3lwaJFrYFAKWUXJyYBjkBJqCT0niEnSf/PngcB2yke
nHu9PpcX8lcwI8xJrNrfIif+ASOeLproKhI2haOeeUkANbNUciunnCJh7xCgeRFs
NLZRNJdA6gLaC+rHNeOTj1ghhnvL3xhk3aTcVjkayn6bS4L/INz7G+b2iHn087mf
VoP9JncC5MUWOt4igzdXwuvh4oMffe1Ot6sA8xlmQUnwjmAUqBKLBrlcIgyXR6xA
8txI9jTwZ9Pr+3DqcndgBFZu2e+DipgHo4/X3SmEFbHmHrrJsd7HwIHyj2PtcKKY
b7Go5HHaO1rTh8iWfMmbI6epoSjcWQ3UYxZZxw/XmLTMQwlU6v9wp8UkFf+f4fAV
rYGPrBYnmzYjlbSx6r6/eg7CqSSgQIeaY91+uP+cSZqS0KkOTE6f8bRWfQM+w8JJ
HgzU/J/S285Ql9sIx40qKbLpVlpirW39ue1munaUgXsXyPx6uXLtAuvI/LUzjpab
8fd5raHXixp0m60jjhTRLUgoF9k+sI6Dd7Svvf08awT6N8UelBsGVxjnXtUFKW9W
w3arvEarUhxtachYNhJ8W7qpEcN3QZMHecpaSB+PGyATv/F7n/d0PtRhFaOWtN+9
lOlN39ALCYfJkmlpupKQiy7JAEENuU364STrGfRqRQtaiG/b/XaureZ69NYWaLPy
f0DMGuGZBrvlTH/4z50D05V3Qy2ENk8vwfc1oZoE1yQi7949+g7fEgbyhLHJFq6u
29AjpAfSBA8WMFLFs3cbCMVKI305WwFTI1QrTH7zBpjWgZahzfIakqXU3LoHD97v
Er875vrlx2Mhq8OCXIMGf+zTscFOY5Y2OGdDxyEHL/XsZNCoj5fTZEq4zny+O+OO
FR91DNwuU98ziPujRndp3jtOl0CTlwzxmGE/0y7Tr52FxWwTvxA93hTnjnelcMhg
vTEImsynXEa+S5BfaogZgUKLoXeOH6A2L7clpaYbAR7MdyObqlYfCWBbpf2acuAP
CdL+6YPX6/xZV8ugxctT/fyw60BSlpc+PYHHUruA80mqC4dMhPN8E3bGlTqZvFb7
PUeqRNw7ZaTKWrR0kDR4ISLYqpuCPW8oAuBZhFkL2H715yrzgDm/RaHxfc9CzCC9
xd/whgUo2BUQha05eF69CnFEMwdLAJ0ebV7VmYniKhE4nfY5LD3PKVCVmBxebBR2
sGjDSGItIGuktDYDIQz34KAmoG1Rr/0aFS//23g/AhvBVRyQM4M3aDDAGewUjAN3
3sSTVbYeIB7IqbX4Thlc4bn3x7X51CSuBZpaFrISmr+nxop27/66ZfUqD59nuZ3v
5fC+Hr4GPQyI6mFsyHmV4JYWmO72L+lGKZnz7toLOHr5CP5yRC7FmAupfFiBhj6M
3LsXkaGN643B47nlLXvb8tiBw8DoCZdvjX5IWLwnyOEDIey2Bjudat/83b6oZhH1
3RZ8nKF2/B1Uv9nifwuoEC+5gf/3q2U9g4R1y5+Hor1cO/RHLAnuPOUfr+N+dr0k
ASWJsf91qiwZXGX9/SPEsQTJ8VZJv98sh35kBhmAk/EfEEzM8OnjQJMY0SG00/Q1
5zywoarK/W8W5iUANyMEu+afZp31Lfgch6BffV+VsR072GjiRs9/QR2oC55rJEbe
ksWuPGsBMML6f+0gmBT/03YY0KVwpSwBptRpRT147M0IgiB+1L1LKnL6KAUsU+ui
LhwNlEeQCxT1230r6IwZJeScej6xin0x6P5oysqDGELT959j9uDjT+STukRMhGUm
n+RyMNjojNedm0YKccpoCAz1LchNWf/gI0bQe6FfcaP9RqgYLKcCEnSWEksZErFh
0s08GNfopoXe0bzRJ9TkEStt93PAy277MzpPBeQGvPPP6D5V+ikSmi1LceKxMf9F
dN/gdzojvowBkoXXS7TAR0Nc0YrYMM2Qj/YkBApE29hX23ngVXLTEYVixidtQ6xY
gwl7Kemnl7t2grOt4qTmB29ctK2YVOoo8IeD8pTNk0UrYLG3IXcvcwv6uItMS7F2
E/tP7T7dgjNEdv97oLmkULZGzRQuH1B6iNSiX9aBlYK1PYGZ9/L63Vyv3+r6OG7c
XJH9tXVGnB8HVtOlxjXQOoo8cHowbIxyUnxGllPrOc55NN36MrqxtydJeV1vx6pR
XRgYHjw2r6Sov8BB6CE/C/vFh0XK8dWleLmX1dqp35tcI4AlVQPesQCSYW50R0cJ
XJ1wRZWt3/0tw4nF41K59h8kVLqMwODpOfOBrWW0LUmygs5ggoebhuUbzqQsEMv6
qcyUeuLxX3eZ/it7MMsqjRzYZ/P/gU9tDDZpCoUw79Kjh5P9sjLG0iPnXN6F6iWt
55hDFq/lHXkhY3gj9oxcoXVPtcLeUcNLhTIw1ijbuFfIcx23IQrFKfOM/Kt3Jv21
qrZTNXn2PF6K1wHjLr/viE4H/z+2FqXr5dfsDxneuIWl1aD3dg++Tiq+XK5lSASz
lv3KPcTEYHf+nckFoorzAcL1Nh/9jJvVJxxqzxOUdxLzrytH8D2cdLc9U6kvOA7S
kTmZyILzAjcxdYz3PbaT4Y0mg/2S3E1neJtb0uWM6ssCvjmJoLZAdouED+Qn2DTl
8Trkfp94zWlTLFCgsLKFSHBAUgrglfewT3cEHzPT4dYISwfE1c8mIo9qVzSd4LZr
`pragma protect end_protected
