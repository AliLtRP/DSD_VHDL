// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
iARCqUjonHoSzp4Mg/Lk7gtIlghoYwCTZ09YDFjzf/0jAbp6zuE+OiEWFZV3teJwRcdFkiKmKonv
b2oFCqDaTfg4T7dhbTbEqfYoNWwDHET2cf246e/q+C5Z74WEhYow3KomxA493f0avNThBUOsmC6O
dVcOMEQCXg9pkuXc0TqgAB+GNywTei2nAZL+GhXa16+qiIahmWMoV2bM2YTIIkfna5t2EDagQbQs
7CwcFXeAi/Qt8m055FbJX6UJlAWekZ0cRP43gcKy0RFxUr0FLzDpzq3xFQqK8ouMW8hs2tA93fA7
DqfvqY6AW/0vkKBA93aRirv4YdjNeuc5acLEdw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
oXLixGkjMjKBCnmGFrjhJRxEfkygG5eRbW5YW2XIcU8SSjVyi7b35bWr+qwtGhSgUN9XIreflq+H
iydNchfXbHxsoQ/md5cRgutf+9xagys3rGiTUjl4xJDue+PSl4GYluTp2fYZ6/6PWAVk1ZGZrY2c
YtPjj2qQ6NF1wlRCZsbMtJ/0fHYfc7+BtCEo/xT7wiBKHtGZCdXhk8dv6fysOLpLfVvNTyKrFaHm
ZTndKBe3Sv/7w+JCGeXXXPKcV3Jdwj/pR+MoIOySIdJLwXdPAQKXk8wO3ZeFwIAT27/I/eMJPURf
a+RkIEtrjplvbonJDa2aBaZVcJ/4l2nm46GGEY6QLTXJGhUWpEfdz2pSpWZ3tBOJE+rMvYwRVlAq
Z0dUv8oTAOMqq9kzzCybJb8g8hfyhcJc9Qou+y58Ir/EaRGG9wNmNeoEj8cWE9l3XsY8Q0C1V3tp
leRRBCbn0QdGwjrmYsTRGRZTqwVzvrJ2zNtmKj8doCCVPYW7xOAujiG1MDb+iD5nkRf2p8pmcBzq
Wnj7GXemytzLi5O6tVnkOTiVWBTaLWMJPaeXKrzoBsjL5VAz0fZj4p4xOle6NcgoD3eI1+OtW2qU
JdF8xZqsviXS9rnH/kjiO/IZJQgETfBOmfII23D3n7EWKa5oQkpctX5vEOf+viuE8YbJd6b9KpRh
11d3y2gqzbSK2Cut43BnEqSR0zdP8FdUMQDI2G/VDFie+hMnJ5kbme6X2WtMZu/uID4k09tMkFDM
kA4cEBIXueTrFvqmbRWBlIZq1G6Ud40k30hwPrtr7q5C3Q/1jao4kJoHOpBaj6vtm2vAP5deaNvt
4zshFgATXTAA7mEd5AAmDapXGku7xJOvw52GIy/AZenILUMKob88EdLdlgbtmdNohC7WbFBDuEdL
/NnViNDAatkTAUWAzV+fIdbk79/nndVsj5YevdGOgrzxovb1asx4/1XIZ0QjyWcJCdKGh1T1vsou
lrV75xMiFvCJwFU5Yf+nwFRwoxkv0MRdgG+0rJCD1QoAS+Upovyvpt2jPNC2Tt4JImw5FDeb6Q7j
xAkjC5LV3CjGMoJjuwlT8sZrcQhiJ8IGsn9i3zpDbwlpSFL0e0BUIh4p6rnY4709Ua+83E3Y6EJk
yhevbZ43gQmCjwfUSw/1lZkXrfzcLFjZ5Asl7yqKXn2vJjSRu6QnY870aqhnXvYwiGsnEYfBigMV
DmYDO9kfW8C/SV4iL+cfy3KRw/XPNMNbegUQgIxSxnIXhvNw4TK+3+sFhNU0Zeh2fKkC/ptnccgH
p3s7EhKzkMPOyXpDb81g/W8GRQvdaJTFQfUq0MMTQfusdrsRJMS47LKQUPlXMeLM8cqny3hYwXok
vOEUQQk+XgQHMB/pQODZfvWAMtAiyVkQEzZtP31zXGfyi3o3qt3h/1mTk6+iTxGys+u3WwuLXhyn
Wtfi1hbSnY/r4mf4oraqs/L5CrzMInUp4xBQGaF0tWzq5zPtEzmAoX2/tistuZPClu16OnONC5db
4VN1GUckMgAQokCExw4r0VEd5PYCEKQ9zRN8gQ3hPzbkNg+ZYQS2FYdfns5tuRJA9Tz8NpXjVvra
fgT42yTZPRJBsTqgd0PCws0RFA0ALGqVmVwuUsbPGjRdQGY4uNIXLugornTYPAWLQWuyHrEdI9XT
aTLkPDdf3uAcKc+/IJRYPMqjZ3HrEcUwolrXxtuD6xUJlhvUtrMdC97EZe6uRwgHuqJXzMGrzg+h
AfuqKgSzrZ1eztpwsj0xVVGbaKTCIx+FcDQqW4EAkEKAsfvuVuQkbjeFWDcXyx6gmk1QcO0RYX/X
Ac+UO+/0Z2WrDYoG0BartUJ5QPXIQRBAQNk7gR3G/fVjgIzU/POGLF9Nunav4XX37Y4pK7uNMZqQ
BLrPkPOK7x0YnTaxvRhyil036kmvtg92nugjJE82FZjGeYPoEuIrmnZfm4KGuSstmy8w3nbh1eEk
wlOCnHuE7kiQNh+7MFf6SXANs1LN10+uhwNbdnojxyVPF7QcRidujs2FToIdQjQPFvhFGqOJfjNs
Bui4+l2GnzSZU816YcERwlcSyEqVRCkTihLs87E0P3iyPfXWbPiWMs9LS/4wJkAkuKij3HhYUdAC
RsDhelL/+aIGbpDKgAKKBHaQq7H0N/bmXTjfse+29RHcgHJMdVtOBWNn1bT/iAnMccVaxiKCpnsR
kK/DnOQg8IxjvSBO3PBWpWx7DdJH1lkMtpLQQLHCChgapNU1IC/b1ToFE65Wc/a9ksT1MSvEr5tW
qrVfGun3tL/i/4U3Xiww898vbPKGzprwUoh1pPksSiCOwqV49tEL7QdXytJWiu6K2ZhrHuWpI949
hAevzkSPNmaGPNtMxgb0V3GiPMYWGenxAGp9F90CR6DEMjTZWKKtxENIH9qPcU3tHA4TJC8F2uA1
5ONZFKq0xAv8BaWNFg//apcoe+Hi9J8iszRxvMV43OKz1U86XUuNeVlCqvti8s51eOVVmOu/LH5E
EVdLaCjmtrrK4e5ZvZS5V0klTjpx24FvTXdm4LNEKRQKypZGWEOHsqtZCP0SwfVHROJTf5UoW5jE
ts1/TrA0JwIbiupz/0cXIZQl9eVLmCahwOS4fHohYLgKWiPcXdhJSFysq3jgB6DX+Xj4GuHSHCw9
0ZYpWW5IguLWw6FovbNEwURdcTz0Fr4R+orTh1kpmGrO0MFC6uQ/xZErTbATmjaY18/Vnk67C0tO
gpL2AinD+CsuTGuM0Rqa/s+p22KEHxiJqo0IRb0Dg9iEUDkEg/ra3JFigQslvmzK/Fm7zzLK6SZh
Upgb3YWMYdSY22kG3MUjv/0+b370E8B/4ZA7fuaqbrkxbuyMfp26WyB4CpZBE7qShG7ZY4w6dlwk
4f49k0ElmS6tRb3svdZvxwxlYGNdMTVGkCh8wYISJ4Vevh1POAonk6YNfoqQiouQK4JFwfjWYJnH
dHx0fCcbSQCzpmoC+Mhx2E5eOA32T9U23/0EM2YCOeNufe+LzcgeAMNmMrC3xpoEAgrwjTOotIfO
6EJumCQ9xQ6GoQuIEb5yNd5MdVSz1w8B3FrUARnnwvAk25SBRzUQ+rcTWxXD4mB5UbFUWHb13WMT
W9ve7mljFdATXj6iUMlVItyB6hyE9/uRcjX2Kk2ssl7QTv9Bd8xtpLf2BwqOhwmXHqC2iPqlp47n
WEwErFiFCOlaDYJO8HxaC3BWi7gczEaDilsKULPVGkdpSNuF6n9U3oayAa1H4lwa+HDe5sFGG0pF
cvbMgKo3jNYRZ/9eDOpubzCLPN8CfeBz/jQ9Zr2TZih+TdHp8hbj7EKpfaqZYkr1X/FA1Ka+VSjT
9QA8SCOOj0tBGJ2MHBC1Sa4gbud2NJ+xrG4U4yeB3VkRAB8buop8+/Ayhsvu1Vp/sWgUzt1ON4d1
EIpBwRvFo5aybvOvKItiddHhp4n3/7JlWy26DQiYhZYCn401IqpTuW727FrOPJW5L5Qvy1hqhHq8
uQtpLrxZpZx/uMhdG1fpDrIlGjXbZTR7qyBhGJ/Ft7gQOVK0IRzu4nMR8EHG59K8zEcyehkZL19/
LR8gGzvaiPEJj5t6pO/Wdtyy/FsYdBPHBE+O4AUu2IQVubmFab05oDqmhVNZm3jVTTRWnhCuPcoX
dgBfDimpDYdrWeYmv/4VxdyNaPXWjkNNWoI72OSpQ2wYFgGYJdZHQE9joiU8aVk6c8hB4UBerB64
0dFBQ35ZAcKk6hBGM/3q1WHsEVJ/aKIDG358qsrueAaW4BjcphKXw+FWay/IKvqjaFTc1mOe5OFY
xf+vzgxQRUCyEHkNy1OR3D3A9D48X+SZ7CgB2UB6sTzCAXMRsEV7o+Gac2y4NWwqg3KpiHRlwytG
p8ZYY+tN5KEVCZJM75RW8OsdoN38h/hksaVDyxZq9XILw9t0Ri6MxHBRmHqQM7QLNnjlkxbDCSHm
XfLty4C/iQFWr2rVCNOZZAY36gjuw/il8BOsa7R0h2SYAf2T71soTnrJUTyCpsY8DF8r38wodu6n
5sUBTteU79WhZn3fSz4mU7RiAF+3dLvo7TL0H6h6D+lBXuQQ312AnImnO0IEgnpm/alEcBYMNqZI
oEElWYzmpcLGH6+NlkqE1vdD9F+D5laZrvulBzg3ETJsSp0uAJkT70cKsOZZDP93zzj9x2yb80Nd
EmjeSNOKKj6uGiy36QAfcFWZokyozhSsvF1HrYwKBpVW84VJjEwHp7zmUyvw7p1tNqwmZZCMwa91
4N7rpPQ03srJnY+W3zgpeBg4cf+hjgUEaDdMtc9ng03SVw7W/zA5Ms1wiI84kudVuFJe+YzknpHI
8eBD49TUjBcRsr4VbyjLznVVJERXduzJbjz0cxw/re+w+//zpzNhX8dPhHUuX9JCopf7UEkDq+PB
SP5lQrqddDq3Wx+rq/xaePLVpyhguYHnNcuCyQ2v3CtylRjR/vDkEGqmM5zA5DZOr6ECIBSq6VGO
dM/JSBGG0ZkMrRvUMhsLUm+g1ucmB+dADEHwgoja5ZCtxU9euxqADqlOEd/ymGZb6gA+58mZwsrL
2e2ghEDx2MCOx7I0WvBE04qVznKadLN90sJ4onZlF5afDy1FhMgf37tVaX7H6VmL6RxZUgjjEjNp
7S6GlVJ0aBWIaTCN3qqa+ku3KPmgr77jwyh1g3pWr+vI+hZR4v8qFEGOc3U0Ex+B7HVX9aPhLoM3
AOxn0URUuZ98jctTVulJnT3d4TOwXH9vHtQ+jtLfFZm8VJMfWGK+9qA1ksYp9z7HZozX0vyv0l33
nk//D71IZ2c6laSPODgJWf+36Yp1id9iRFNBKKZWJtC2VKP+0PC4DKM8XiobO7UParDcrDJ5EoY9
NFlynC0X++/1TisbV6ESFQgPuaERlbtTtR37IuhvCD18ZFx4b6v9IeTzbyiRuuSqQOkn/LURijqc
8LHjlNsbhXZunzIqG5pPnCZUKQx98Ip/nPaT1nhY/3EBvEZ5A353T4trAehgAfH9iv49M0X1bYJI
ZkvMIujS2RKczJJjCPzMkkkApPc9UWupb1Sm4G7P5IXwxg32zNADsxBlihaOvRgZm9eiqlEMio7L
DzpRjswdFslVHjuWaK42ZZKRJghheocDDgqSwfiLM1jHxVB/ivNtEyudr2Rzcxj9Dc829sXBxB/3
5+5nGDdAhdc9PI9B8bDv8mHGIQxLJH3jauR+nUi8F8zIgXUAzdnVSbbLwoLjqrDyl1wE+zZv+A/+
xQiM6xbJE3O4oCM36MC3z+rdtiGPnsqqSzqAiHVYO2UPqhE7DcHZOEYfhc0CLmRoTWUa6x7sp9Zp
eRmr6F1XT/ZG7Mw6ikcno3cMLp7SCSo6iblxd53VMsaXVLKVbvbWQw5dqaxNbAdKbfOB8kK42u06
ITuSE3CahzTAqp0iakKxkXHlFgp24u4sD+C/EU6mVvegmhL+mbsCJj8F+MJmBJq7v3hx2wxmqf1n
HZ1qJadZxNoNCEv/MT9/NRwls1S6cRe8LKR88Dn5wsqcgrx6YvvoKzq81fuGQc7iQPnIep7OijFv
2TJep+X7ZXSeqAkPzknlC9Rl3G0ULKQ2HSECrJxT5zU7pU/eLSEhayAXqdLF2e+28DBeGQdNclTa
B1WX2YzK0eTvXYZnvK3ZePqolgEwEFRadXSGJ9wYI813r3C1MF3FbwsoE3UOr1ILCOph3OdURwNe
NSpDguNJZ7G55wQzA9pbJW1t2xDVMGFb7T+yYbSlRqVLdOsq43nGMWR5LDzdy91IKhvdbs2Fv2Xk
cpdvV7S/YjgJ1MWksNUkAC/2/MtyisQEOcloDrd1MAnkQVb1+cIwTHRcJ2jiE0GIUg8YZSfLUg67
2U1gm0GnQ5742P3UNGZJ2upfrUjVPVaZxwIPmH+T8GCysvP/KHoieQhTLDQ5NBtnUz+2t856Sz7O
2Wlqn9BPXJqF1vC3YlcAhazHey4uV9+tqaNga67Aiz8YLnxtH3jfZVy0R6YeLZtSFzzd50OWChgx
MztBMM99XsXdg2mdY/P5k/VUOr0W7RpY861cEJy8ioDWutM2+XNcRY0SSdoJtWeaexaor3+3YvJd
OsYnetey5WMo50YK4Y1fZeK/BaFIzDlsqhqGrpIBvujjrujLwPdSJ6I1l2TB1S/RGK8bs+dG30k7
9CsrCd/xYQX5Kw4MP3j4NVsYCwUFTryEuCC2ChlbFxG0YvRKbITScnk/FvNETZ7gj+vwsPML+Tx8
Cf565m590zWa4prn0caey7avIdC5Kc5JJC+qgD92lI0e6sEV+qdWrarYjlBvmXnNk9Zzt65Dwxf9
fuRPGnqONcBVNzPn8BSDsZSs7/Gozi1VGCfx5/db4+DS343H14eGoG0hdQSpEUPZ6T4M4ysqGcvU
O7H7huNXiFZzI6h6gMC6L6TC7LHVxIqJgBhGYZU3Koy4thgMq0cQzO9oOXlfcV8bIazMJNr0Hj/n
9AmRPqgRx/dYSTNP4XjTBiZLZvezgiFBXNcWM6trWVpSOU1khGW8wDwtbYa30vDAaakw1n4FQHg8
+GA31mxmm2DacQHlO1CjavZkPbJroUcyLQ8hi5zFE+B69IwA9AoNh5Erbz4PhGLw117m0AoJvNJD
MZVWgOkSwP0fTxBhDrK1rtS19u1LMYf5vOO528GVEzAStLxrQ69koxnLWI9Ir70EiX1qqX9abA8b
N9nw7XenEFqkO69BYP7861iiAicVz/93lyRx6i7ZQA4S3UScZsvnUFG2DmYTDzCfjjuVLtDfmU4a
rRlCR3VH5sIPMABN8gQ4Enguzaw0fY72jG7SOdi6x2xtdQmLKFFxyygFcPrR8H+DWnI6fOSEs74E
5JqpvyApYz6OPvDqmHr4dSpiYm+8FdDUhszrQoYy4Vu2+vB4j/9jcQxIDa6vmY1mrj9PGUYY7s7n
XPwh9AAuPqoPy/1LawYdxPySB+vQr07scvpqRbivJRfRVOJtVkANQo52VZW0fgg9Wj2pNKkwzpjd
KurIZ+jXZ6Zb2JLTQvAvq5GtyOCJpMtGMlMkC8iUcAngCkjpfSNoahypzQOE1fPEY91cgCpvIWrO
CIx8+eWUNcV482EQZlS4oQGxyQqJfxx8D4GhqbBnqp8Q4ynhNf5cvFJvB60TRA7czh7QR9gnfSn9
LV0y6VPotWwmsua4wPt2WIqmG3uV1XdlPHBrBM47fK/MYp7tRk5toQhOV6f0ZbDm5wo/dfinhyks
Gji6FlPOfsP6yQaCnMMqu7Bsm7IBX07wzNYEuP9YPowbcB2OWKVGArWh4BkY0pgQhAX/+x6mP9k0
TZiuHgwMXZ8pkVKi2Xm5qGaZXAJQVPMkEKy6bjfEGNVgHS9q+2C/4rCHOwYYYGcAkk37Lrnhx/Lp
dBsAZjPUiDxIYWa7FpVfwS8nfG3u3QWf9lA/a1IDsEjBHVxlI2XxkoX9zrXqL5Mph5ooo7opEa2f
AZfPwR77Pai4XzRYceh8+OwUJVf/eZ1UosSDCcfgONANfghwPH/Dfu/wiaSBCUQ949hu60sU4Z2d
57UJlOS8ZQh82M++w2BQgTZZhxfSCskiSpJB54gXaubT2dEoP97h64EgIiG7n8877GpaGObHBhX1
6DzzbwoNKU+UOOX64oxKl4RtxS0qKQuMMJP/ju+GczzXzi7ewC2wywkeUUmHThqij6MszPFVFP/C
XxJdm/5qn30b2xP/TZUklFBSRAMrqwhob0q6uLiTzpVcpNY957lA10MswuaUFEI4WjLmoWnV88eu
aG9+Nn4FRUemcGFjHF2iyJe9eaQhVV/GP0lrgTvatAGkjpcYkR3QrGxGyXCKjBPp2tQ0c5/HBNvG
J2hgDOy7HhMeKVrS0aaw8HiBOM7yx0rhtaHZWzcPOvGapOOgWQSmpDp6uMhvv0Be0G6RTH8tnvDQ
RfFqiSITkCQUcqZwxvE9gVvJ+HPN+wt8pbeXjrrGAzgMWRGx/kM2aUxR+PmTMe5XRfnU3YwpEkyc
Cd5vY1Fmz/HHvzVR8YB7M+SGJnJn4UFmV8HNVdxdsEpMhUU7kF2QwcLoDjBorFMSbiDxnSPA0kTx
BxPVADiOrRh44aSoSp3GZX5Hnhaopvt35g2Nf3co8wPiJ6oeRFJdmLaFhZ4pl9YhJlQ4GIoyOV9w
nKFNUcPM81QPaeSc2TX/zulib7LtoMJt2udvdngx6XlO5bFCuvRVliiKlVYtzHna3G08I/cvPUxb
62dJ3BltGWX15dM0YUnU2yAUja/g3JF2JraDBLgSMVKAZWWBX8yrikRx+sGwEa9ZR4OngGXY2Ayy
kh6q6VFmR/XbypOzVNQIC37lguFCl/1Rir3liehVbP8AixWZA0vCPaWt6KaS248nGRM7xg26y5SF
yrW6PujH/eHV5QyWk0Mqd7+kg/RQmp9tbDDXDOs4KNFxBcYXeqJfFVejiAtwK/1vaRR0C/ppIF/e
vcZpL4SEsi5JnvDT8uW3jNxqJRfV2F4E6s6Xa/o6F82TAv6IdILsAhVYo8jIXQFZLdl1zeT8ZNWn
f0kFGqyNxlJNA0LsZpUSTJFyrLd1tzpOc7oUP4Ofco1y0D7EQj56lq85pGGHEBiSUuk9i4K8eIM8
dGtSi0aDOqbaAKf39ffKVbSFly5cB89gZm08Q0t4DbnUMJHO+Fhdmb3egON8k5X9Hj38ucFwEgmA
mHqjYQ9cVDo23RHBQt9Mw/ELAEeMFbGavgb8MGgG+MN8Ae0LPJM/cOcwrCoSe/XnJtu5pDb4BFtA
ZhD8oHg6SPcivK8D2fIAi7rN6D+5yFeWrKz8KpxGElAqpCj7s9YcAjBxp0pS+P0r6GjeTPASD4dQ
qrwVuuQTxPxChqy0xYjkMySZknfuFvd5aTJPIcv5koqsFDwmxfb5QMKGm40udiaVqcOGIIttnrv4
9ClzHSeCVPu03d3PjVjTWtqPCVnywFBTWuhW9FMYD2h62J7kTrhKLMcDF3m0+4l5DlONI/BvJu+T
NxGJL1Sb42Tbd/DFn+c+ZYS+cWbM7/mOB++gVT16H6dhW80nNDfXcSc0PC6d6ssK/9clfKOjVoOl
YuWlwxK9/QiJumdvE/sbmOwcq6XCG9GNKdQzPK1MeSfBazMueCwGmh1y8msHMpGEcaNmFpId6mOd
nC9nQmAux65HUPcOUjgOHsa9wrNTjpxQNhSfaty/nx4FS0yhLMwfMdH3+SyRmgLDhZ1jM4ZtwPyA
Yg5+EEL7rTHIxHdXd/G7OrzXQwpQY7lus8+O5qUcd0vd87Ir4s5GhYDSMP9mAEzDtP21wP+h/D4d
X4GDYtjMgWDANeN1IXtE8loFQekAh9PpwC0FdjDiQbDvYeN27B1YcKiheaVfUZ+IpHjLbQHrRo6i
J8VeIU/AdeeAGLfS+Q8/Zco8nbF0NRG5halY4hy6fUizAnCmV9iMDHGVSQmdl60n2+5L1ZoJ2GBb
4LcQ6s1qnQbUris8T3dj2BlTElYyTB3wB7aCWz/1jLpta4kndRFVbxHErLTMx0eztUR3otsafCOg
bYC5H11mOkw/mSPdIZZz5kEbQ92AtjG9q/bib55DRz0SSlIzwUuAtriLMudfw8lvnrexYoE+BemO
3o3CP6VXmjOtUVoZcS1UkTcVkTkdrDoLHmmZPq8x6SvHL+El1vpzPTPJ0vA9LPkI4XmtkP+JVHdH
I7i7dZvBJCcmcnoThcQZzE4TnRtcjuaqX+EhMBaYhWo06NImzEfWjqgVd3bFXjIm8Ni/5MEkl+vh
wB+QzQoVSnDfPWTc1hl20qczPz1TEvcd3jp4RdOTYGcytXoxt86mvUCYKLQhw0N+kbJaThAMz7fl
wh9aPtKKe/nZK9FcNMXV4nx8fyJqDBY7wEv3QeIQCm+Qqp5wLVKYaBDiRYA3sFv5zMVM6Yd0GtrO
ASSp2Wj/29oXVg5/Y+A9foupmyGwegFUjKJZEVnOzbxORfp01GcUzwOmuFxmXUYjTIvjS0EqsonZ
uqgNsAjZ3FRstA/mFH2H84rBEsxD9P8yBtWZFyU9MV74QRthubcaGvKsgzOQ7qGuCGOPt/CE/TJo
e+1h3L1a4eFXTmMQbSWsaisP9sy9+M8Rbq9W/VX51RCoPA8lhpDq7My8Ve0mR7Cel41y5lkbLV0Y
E7NFTkXDqBjLxhDPd4h4Env21K7lQ/yVQDtva0g7z7luKvFoEWxSagB/3QxyUUtMWYWknGPBJBwR
Bql7a63WADAUTlDosfSSkWwHgBW2r+IM7n0PPdwria3ThCdLuAjBoa5IoetAPsTkDMmTrv+TMIqC
NeWHn8cUJhZblvOW5Aj7rUfU2CSxYwBnhS0TttyEOz0Z1VCUtjid/cZI9rgZlk3qihPpRo3YWu6Z
iiDWWI9TE4cGvey52DBMaBzpHHcaEQDJ3JFvtgpC8Owlt2SucmSoF7gEYe5RTHeY5nXjTl1nvnpl
K2s0sCB5/rN9++LjlLw7XRu5TWUdSUWdelEYjFuUXdfn9SVJAa6mqMVdha4I1PpR+6O8LehtBw3O
MgvKDOYdJGXBffGm4nPZQcWXYlkp5S/0ZHd4kZuTolWfFz3kip7QP8I+K7erzjZdy8jSci7gi4Ei
cpQmgwE3sbRbDUZBSZF92IsZXqtxxu6HhBx3k8lk1eAO9eHRV6nrCfNDTl8teFl3AFCeixt9Z/Ua
5kDbu6rLU4rRq2hkxXUqvjW3WhyOJeBd1n1GcsHKFDY1+dMI7UbpVllk6XUbC/z+Jb3tZ6//Nhp7
Zy2s9q/uUeuYmbS5bQZkrAq1c/6xiJPm4CWuReM8fRZdsNmhxwDSQCqJnaE5Afa5CmbY3k+LUIXY
BHsCBDv3BgiNZscQUasP81n3ZsBQ0eWbvWXihKym+PJYEXjRIUX/qPy5lzpSJKqnU0eWtQfNGK0H
4xhc4jhP67bk/WabCi9DLdbEdrsR7kXgNspdYwglNm6lFHHfzGttdIRUBlzGWp7thZHfYWhJiZLV
PXIlGto4kJkxj685GDg0C3hmQuT900CJ1hEr6SrsR2YQzyzfLyT3YSvsN2Yi79mKrjIlNaPU+l4n
qwNZ8vZhK/W9ubDZWDLRNfTSqz7IhEcyqBUIxQGzBzsuctw1nxX88o6Y52/JEMCAWRd64O0/fgKt
lbmbMh9vl75dmgp7NhLadwZCKLF2bJ8TqGP0H2WZ2H+do18SYKa6oSuOTHLy/cNEJC97pW5rEKUY
8MYfwbRgUGGwrXeogNJ5mcFjFeb2u66fAuiFiMHseVPdVmouJFTZkgGAcESdU1IDH6Dp+Q2VFhfB
ibULHXt7D2i0RfIpw8RRYJQm9510VBCCbz4a7Pw3nAFeJM813y52C0IRzgvkdhVqdVB1aayNSf5F
pAO4EovKOiK2NLwMqX0ssSBjXsNErK0EyQJYUkDHmU8vNmnGzT9QDNg9BVXAGhevrIwOkDpJ9DRq
c4cDzpqAYQyZfScoBQKHXyO+z4Lc57yVObX0zUCu66zG6uYd7T3SF3PkYTwL3Vw8AjiUKp4ZOU/Y
KpjmgQKV+cMFyWPcnttdkS1r7hN0Ue8Vg3XyOiXidbze+5gyGjmVTkIpkz0394ljBtmc2eOLX4XQ
Ds7DIUlG63K+RY8VWZzkQiCKbD0f88faatLnq0p+7sXaGXYrSPJigCCd90ONSS8iC6XDL5eQIQqI
GyoRxT+30OvCa1Ry3YLS+/RNG9kro6DtxRd8JAp6I/nwSDzZvpe4WS6IvMIyIZBiazLz8llBZ9ym
UAOeicNVuqoOWtwMblCAXSDT1OtT+qXnzu0RCRged5O+NA7UVksEzz3ldNJ62BZNzN66HMKNEjGe
UqSSEUaCeqrvrCUVCm+XjRremJqlELEhr/O/TdIIfKRyhIsXMmYMYRfGPudXHYzryv2NT3XRosMl
GV9R26cIKwfu0hVd87VDh85ovBHRbwbObUsNkojdab6HGwZqwqbmLnIH8e7mnrTgApbjLH/KJ1Fz
NVOIkrofN/GQXYT2zS1pggE/RNKg7KHYRZZ3wNW1CT5qiPpt3L7jUzBDdk3n2EWzo4LSrDv6O8Lm
b/MamIJtkAbMz9v6K1ctsQQ41jQ02NGAhLG6fE2P0VlcpK8b1WI/nzgNoxAx7/dUka296000rxTy
kzBPeHcNWWsVdTev1uOcWjWmOcONmhrlQ8Evtf3/8ZCo5PcmahPo6pCsoH0l3UVl+EHpJ04QQLpG
rlXaFbJacYqGgiKOz9OrDHLEditZLS14n1hwdyYnzsZxhf0S6H2daebSHFe9xrQo/KlUVcwHgkb4
1k2BIrsUS5LDAEptIAeUcsSa6wbsoumyxLMvQ2UdZw8V6zww03twmc09U7paWZijduNZZU+C3leC
B2/lmQ0LnfbnEhVlR8OmRd/Z2tZTYXjj1ir12/yz6FrBAXHOdskORAm3l6wZvFyYsUH2o4uT4iJy
7W4inagWr/kmTU85rrqw0roLC70JD3NXPbZv/jagmBDiy8z/DH66EO4R/uufDYW/M6Zm2U+cVXon
rODMS+vsB89DeLW1FKgsqlxuBbb1iiRJ3ipfzDIN5lV4MIdV0YJv8HFUQZOcO+Mc91FbWSOLyQHD
OwOF2AiTy2+folYfLBB4bEMmLdR5W78BTGlzsVlS/99ZxhgfcTNVSx3O4yJkeb1rocK3d65K2WJa
p2bkLy45mPvv48cKNMRhO1RrZdvg+YjLAK6EppjizT0iMj9XiP3aj6tsvHzScStnuMRk8Om7CZZ7
Rp/yZleqGMSetW/yDxuC2zZIGXKjvik9L546hJfLi3kHgO2SbKMHou7vfS8IL6Ai6LhU99YvQTN7
GOtaZMT8JgG4zNd3QsV7/W04lk26xgPCHXNxcMjjrSLpm82OHU3Z9/5ucSoaaFfuaLIYs9zv0wD/
QQaR88+oHfXPXTaPu3mFFyCJFe6sHbVryzDQyVM7/e0vEzl5qEQDHzS0uj6zEUxMrduSeT2FKCLO
Khw5lryMyOhHFq1gtLIZ4ZgldhlSCTuCT3nTUN2702pQj8FJiwtBbWFbgf9DmgpxkGvLEZFg8M3l
ZHaoYZ+sIrBv17mNsMEjRj7yYjjtEMg+nse/FG7lXuElgvgwL2DicUQes8twLiCeUjfnd1R1Xcib
x5KEYH+sSU2jh2TF8qXYpO+NDOkTmFS9jv64ASJlXWAHnX34aHqD7NQf/UJsY4C4nKLe7jWlswaT
f3I23SXc2WyRR8WJfEljL/MagrJuLKI8r6QjauBxF5d+bVo4JSFoAXIOezFY+MGOY0Dy4hR0Wp3r
D5mBZQ9gKtOc7EHUlbOYEJDHMaGee93ukYB0rwfLCLUweM28mXEfCi7GrK/RWTvqv1OCQRT75B5I
ZpPw1iAa7R77Zi/qRucwT9ZFGenB6ppye3A9fjGyCxEGK0YpU3vQEl7ZikuLrf1M8+U4bE5MuiGm
nWSgx79Ho9G33ZDTCTHJqQORI5c/mOx+2SoJMtxoaBgqpFOLlM9kobdwzquTLTMtfFOioAFSpVIw
Jlf1YINfbTaUnT3cS1s0igiYoRUa527m/CRCH7/Uc+3wOcelaQoUqbz4DSMcqkGWvFIcUhuHgKRw
xN4ESX+WHCA2IAKb+yA/vkig7mHFeYKSQ7mOBnm4klFqa8Kld64quK7hDwtfzl2UFmI5ieVTiqja
0xHUQVFVrqGJUi9KxKTNCkffzSx7Bm04Iokfn8V07gl+1Hdd8H63mMm7Prvqvx389384/XxwIHyu
ueniix4x0BbFk851cVFWkyOj8LyqxhsGdNFeFhQY8FOmapi+oX8OocA+R9LG5fZGXgSQfmTo2k+J
sJxkfvmhE+zAOSdYBHsZLvlIQL1AVHI+LyZo0fKXmTDoid6IMhwCFJHEAM0NyVdwmC9kaUzod7XQ
uh6Z9z6XJ3AL5fiSePDLiI+Bcemdk7D1ykhmrIVfZBjoouXR4Aa4cY9UQnepfY6xIWwBg2rXmKF7
RPkzH8I4KugNCc6PE3GM6MPmE8mzhX/HNgXc7bCi7uddnVx1zed1xdOtGvNiy+PW3I8lCqNkq05c
0p6xUrlcjbJ9GAxDUlTmE1jE96kOHHgEp2mWruaBXn6Le+LgoCkjODJAqrnIlgLGMeJrR2PypDtO
LIIjSfSJn7OWm4Th5xOsvLf6Bjg8avi8Xj8+jhKv1WSCgADg65tLo500iXDygCNrqjeuz3bVZwQ+
jyf7ag72jRZ3oEV91Blz0yHys0eDUa49qh8O1qucjE+jB91Nar6ybIThe+ACKp+NGiVYgRN+aB3D
jrydQi4D40+T+ifRv3hK2Nj2FjNcnUv9jBbn6NnuF65btyPtxTNC+1sZMSv19sj/Sa+bAbGZkjcY
GS5Djlx0xfkdgqyBHMrAHQLL9a8WzzIpUCTBduRjbKWcR9nY1C+e0i+okAMlpiABiMGzSLBFdhi0
cCFO94edtDQ3aUibVNRdV/kDXNZAdhIf//d8btl2Bgn2CTHQvGoD1LkySRw+j/oBo/znerGuCsIi
Xz7gupRJmhX3/JLqc5yej51mVkFyyApb4MpVt+wW6g4JM2n0lMeZdMrx/dvYV4rmPfOLq+48lY8n
SEg/NHdfeSGYpsw3CjJcTZD/FLlrWd093AJZg9oqRu2Fkok83HEVyl9gcy1EAsuiwiWten6APDbK
2Zf9Dn4ZiabfKT/pRfvMMMSw/Gwr86NNowxHjX0aJnhiU95xG9xI6i3bKlC1XZuUpMTzQvya8Q6n
ucugmU0FYFzwhZUusb4yf4P68WRK8LZkkWggPBBVKs/e0iXwHq+fW2yCLO5Jr42xPVggSaZWthuF
A/r9UV0xnzlY7BDCipYPSzlaeNnzgiFC1qadCBUtta9FTRzrdLJmGtgCR844S/o9i/6HYlW/GEGV
t6S+VKZqqyL7fC1x3befCT7N+H2p7t/zFy74pVZjXHts/JIc7rErO/EM1hB97Q4IG5mZazRPTb2t
mOP/cJ+oKGqLZJAcqsk2rnlQ7oaOM2YU47kENvI1fWIARhpL8hD+ZYFO9T1qKI0Cgzg1FsRVCR0z
7W3j22lMEDIk/Wscopsk5uydbVpzyOo8PJAjRX3cF2XaQ2k/dTBZx32lJ5FNqXDB9cmjuaNK0z6R
CEflo/5iayqUk6GH7l5SAkAiy55FDz9jDyiAr0PXBPqe3QikeJqCYBD/bPh42VDN21LDAFHTAD70
qyKL45GxHaOPw/bSfNMOgt78dlgZToSDxmVJGNkKXrllUXZPla1CpfFQFK0ZEw29393EIU9OtRC4
9+n2SZ13fjsPlITwXpX0lGoKnDf0fsE05BgDPr2R6JDu6Ohs1vnKFkNgf2vpVwAaJnHN1Dyv2uQ/
AfjFUCYJABQbSmQmIRgmyJ1nEv72SHYruVOR/tdW1m4GHkxfej1yT6NuQlEuO9G5F+ze4vNjTLPS
lxF0uxSOZ6cq9K4T2VyRhVqh46t321j5X4FRaanorEviI3IT+3LjsrCDVYMaf95YJarvjnL16Ef2
HSgWJ39q8n8OaHF3uGh0p6Ux//fcU9eHBktYdWhM/xNWW8IdLoqkl7uQ61eD6rXOW20MSwtTiMVq
0SoMlQuAciWiJCibwAM1cOfBEVjbdNmzU/3JQZfNoPfW8+2cuTA4aMYJzQQpeq3PBcGvaOvumeAb
xUSZCzhtdxLt/EXd3Nu55OvYrcJe3YVhsh1zMbC/Xcg9gyhGZ6YOaFeQXrFUunY2Fb5dqjLk5gVn
2WQZJHomJ+xkLiQpqGlf6HMj4p9P/ODNaVBwOZlLhQfldduo6au828ZjXqMO3A3UuiA306bocszw
+Hk9a4mQL59ChP/QpjKPqO5P41fAvmc0ZfIjIyo9dXyCnndRCm+jIfPX2tLW7WvIZ8c3HVntRwR9
PE2RVL2HM1T3k0qE/KpKPpG1/zKYLSPD94+kHErMIWb0EONvb7JPyUK7nhcCbpdU9Iak3P7MIKCD
sg8WTAqtEEMXZrIv+YNxXVtRfFpaK4pcdweRVeGf5I8Ho3VuvAwxM9VwOXYkWghiRx9uPRXC5gVj
1egWz5j/USv9E99nsWEky0Kfb8/gFg7eBKxW03IRdJK25yjJDLbwRYsdNZlRTskyokhviDobrmNp
iq2NmVnWzM6vvP6wG7o/FLFmEVzwEy6ov5ue4NsswTSwc07R3X1cTXMPRjwFShGTk+DjkQ2W3DNV
O+uXGupWGDhBYjRxrcQL7RxtdlMb9HzD6+GjswZYYeVTocDhIVWBEASkErlQP/AcILLI1HHDLwkf
FU1TowGUaBxXcY9YYHYg5VJrqwhvwVqNMDTfViCfRp22N36T0cnuMNGC7j9tvsIhxYtSHwjAA+To
K7feTsWsIv3uhB4IHtSIulAe0KEWXZqDDgfPNbeZLxEYy2dTooCtKrZxzdlOnqsyEIXEH2r5otYD
SGe8s40Inmr0I70lWX7BAFnVvyAueDSojFlXmdLJFbmfGD+Zk0fqA8lzeri6ImH/1kMTa8+MGMTY
i1xlQ9YBP0Egg4egm9pGJ2FbaWBmnF9pX1BkiYP62/L4qeT9IDfsWqvQWlORnDlxM/b1pg+/bFHW
Bv864SXMbBot6kUzjGsdilzcSEGXJNieGj2bE5uEKbyZqBqEfjNu1sFXSOxQ4dt6X8S/W4zEUAJF
bSgx4tWc9mHSaAgmnuOPRZwoV+fgpN6Zrmd8JQUED6Oc8Sfp0L4iT9DSqN7b/9u6ohoXRg2pXZ62
imzLeHYIyfkPZpRuWKJ591mSnEjBbTf9TY8Jd0gCP9qPiB9H6dpH8uAWhBeFSNmILAMlD+dl90yA
GURZBHjRL6nyqOVeMANDxIGWFVprWaaT/McY39Y8tnsKyEAW/8YSrrYvc749tB2fIAp163BQPRGh
DZIP6kYl5RZALw+tG/Y7so0G2nB2E03ZNWre/rrtbXZZVQNlmxC42oPgpKd6TovqNTLhS6RJfaXr
OxlLGya6pTUo0eqqdfQseCIJO0Pyko4p9Y/u39iwonmKQB+j2qZwRJAdjCQvC6FjmP6bswuxVUWr
PpzbJ5j3TmOqvTcEqW8c+qqcwAaWsmK3OGPaw/ieY9faujPZyC6S7PCDX+KKWG/qT+4FssDMdDdX
jScYiNwV8vnsLVtQTgflaTimC6o0tLfqxUn77DHbfkXM/LjpFzPQntyWDHieIiTPRl/arQwKbSWH
P30wh8pk2C6YkOhLWLT35HO1YDLV7AXVGCE8kkIrgiQZGPSZDWxRNjMG3Q+/ORrX/t4ECq61CW88
LL7XGYuY6SLmUG1C5flPznyYlhC/WGuiM0buJ50Mz85Ob3EbCKMzF6rsXWrMZsSJYE+KlVKzHw0a
crdveE05Vwg0sLt1pnpgjx1qbPsRSa1CQpNLc1p9UDOdKzQoUPO6pibglq1OEfYTyY4ArvXJueW9
ZrfJ2N6ASnUyz1KOaclt22cHEdiHiY7MRv8R6EKuEFGM8dxTb1nUjH5Bq95G3qQeTlB4G+VrUunp
DXs7yLXHQk1KnYu5Q5H+axotelMNjjz8ZTXECtmjyJK836F0slr6xQWfuPBc0Jmjhwy8Wk1r+I1X
zAQySNgCFd089Jiadw3DLDz32bS3gLm7p3c0WELygZYVcpyvBIczuOazi8eLpR2J1TALcdcI5u/K
hCxSBJINgK1T/7OuYSRGjcFWnSRV8/bo5/R9e0fL7EGqgHRPmtDHSyPXDYDCiapWH+lteJtDbjR1
mojnFqkEs70obqS5ng1wGtuM0xAXTseeOlUUbE2DmG/5SsWgZr4ObrBlTaXQ1brGKSW1Rg4TMJrk
PBsPXY5GkyiokVY89+vOq6iR3zOnMyZstPnBdBqL3r01J4DkyWdUkTZcBv3pwhWf/Q+yXkqnDe9+
b+bVF60eE86VqqE8WGhPuyKJ7sNssxjtUo8x1nfGuG12MIXZvAuklH3h6Udhs8B4cRlo5MYvDPrp
br9tvONKByYkxNzTqcAZRPZSYpPN/XySMCK1zhYsBme8nRI4su7eSeKkGSQGVXEhlxgC9U9WaVES
P+jP+SvlQL6kjr94iebtKKhHfOMMhzrNj77NGOXxx96g01EmYJZoUGsxVCEsl4hNhhkijC9CDK6o
OUr76D+X61unGZerLp7/SRkZRffZ6KeqAU8dW9DintSRIPO3T0Q1a0miyg8F5KscDX66jcRg2g7U
pV8N21YMVOQ/G9hgLqvUw61kL0Bp152ZMg/vc2Hxcz1NTw3dz8uleSzThNvauYYnXHHmyaU1K52V
eLmWnTIItkCaSn0MM1S55LGt1XD2gJtzfyjuCboXNWvnfZ7raYZFa9BCeuGjd+TH9FAChduXhGNo
7oDKXJtSJmUJAlOM9G+1YQ0BpGbczm9YumEcwxUYg2o2hXh8TB+5Bwb01s/ECr4UQNuFSMIQJbUg
f70ar4UwadtLdNl9xW4lUs0G2JWQbrFS5iduuPWYiteYlDtRz9KhppSogphY44sZlW9u4LdS+SKo
M+q2/j9DrCwbygZmFpk6HUWOSNeHvyBSAQ/vNYysJcnr9gzGqo3lndrU0nwZYyZGVKazH8U7kAbZ
34ARGzm+G3jneIgedn1D0UhqHHunuVGWoDYwoNcTsXQe1e5tjSEggJXEgGYrEUCu5cmFMJqvHUo2
6nKC3DzeJVcXwEkJbLxQzGsYxU6O2b05MmTBwl0rdqJRYpK8tcJOJW0s5ySSpSH/H3DZ9itfawy5
vVLOMDND28xXUdeBa9J0+ohajlRajLDKD+5X5KIWkiF0t/m6fLSGUOfw3iZ3YlEhIXi1ilD2FFO1
5Q6Sd52LAc9RAL8pQOZnBbeG52re0pljaBk5bzC5UXv27qpRf2sJT+M43jSs4PqGjMS3bwQl7Ew5
KbuU/fMd2/l5Fe9QI36MzEXOvUYcX81ok0NkAm7yzxJX0QCKY+gX2DrBJAEL08IZWPGbDWeKFCbB
VTlrSiJt651G8j9hCI8jOR7526ePqozUxz/gm4hqbwCcKKPuMtgeuP26tG3ojPtn0M9VeO8ju+kP
NOS9BHu+/zpYRXsAY73Vaj0uS9Bh2b2Z1vbmZQpo/wQfo8+oeQCnrSBdwNmNY8k+sN31+Gnb1yyB
22Fc/euZkVpFgb5+jO/Rp/Nw+f8LOcIrCOP8BnIGSxuf4mcxANVRUJS3LMjUjoG81Eq8HHh/Fsb+
bDN2YcxhuMWGBFwwklGoatvQgmUjGE+hJ39emkbVyxJ1fn/+ClYVfZ+EHHGnu/c2y/+kbRk9gKUr
dj2s07CZ9X3CUWrtGwRDxCunJ2OnoaMyWcauJt3SIJpruRmWWxvll3NzMo74FN/4tMfr4ydWZkXV
oKz8E/0xeFBDUUcqln3FtDrF7+1vjCC/fTJszTTLt7CG0+DBeQvIUIABh0fjKEtLq0Yv+FDsOS9A
WSKxJSGvV6aM4glRVJHuATO3v9ycCqN857OBTq7/QnfMC7BlakxUTiyzshn+rgzliL8uh8H031SO
8kP4Vbl9YN9GPpDBHhUkUZTEaGDd7Bujm4kRcY+UDwPWFNeru7bJ1Ypc1u0dVZXE1jhCMlOIN0Xe
H8bgLn0KOedwM2KDDYQyzMWiejun19WC3i6hiQjvIlU1/oDmMcMqMaprldX21dAnNEwYwW5CVl8M
181DQV12TIgu5mBalKCbBWdu+ZR6+GvUY3MLpKs2ojgYqJ2d8rScQ1x74zDzPbnfOGerBWh01+cf
fFDUN4oGDovqConvIoWGKrvkUA8QDzmLWt4aSBTvPvg73wLb2Gv/eKCUeM3MlVK0uNGFwEJHSmYI
KUkrgwalKQUWl2OCrmz8GCG0Xk9Pm1ymzRHt8ZjwOclkaMMEQ3K3DCKckHUSMeSG0rRAgIG76RiS
NAGqlKwS56hJ6q4tf7WbNtZHpsNOu0u6MUaSR6nFbhHBYV3C87cOu3hLTb7ScMmxWS2XtjgHgNPX
qq3F0hH887Hw1oVU7sjHJ4txuhWsCj4Zp2RzCsKu+qHebRIhWlunWLUFGUJbOPfKL6pdUSt6RlL3
u14hEdgtwKwW6vjWwMjCyMLCqnDL/2fS6zBq+lJf1IrJdn7kkC6mDqvxaFXMfAJNkCG/OnuuL7tp
AXH7GeyWs1M2x7TlSi01a1U3nL7eQPxitpi1bQLXKQasf3kfMrJynwY/jF+k/VdwWQHQGT4Ep13U
9RqrDiX/JFV2pNT3psW8O8mAg8qEkt73Z+xcfUEMWU86kzVyNYl5BBP5C0I3YRUcupW9APA0PiSU
5Pre6N7t1083+ar1AfS2sWBazgVWugQope+ZHV4XC0Ratf3r+1snLoWFhh0/S/5C5Nb3EZNr/0cI
HQmAjJnzjfn7t8FtC2Ydd/JYel+yO8iPheZC5B/AG7g/XRiOHlk9cPZku02vhOfTDyOCQRTSSu/X
B9KEwSuCJB+GVYGvpcEC1HDcJIFm1oU7zAluZED9PcluqQmdsBqILUuqtemttZph7vcauWeP2Mt+
AbU88WdR2wyK+RmsGJI+DMsbYOgVafJ2wtVxhyCcreawnge3Ci3YFUnUa+pcjOs72GDcmGx34M6G
3H1xLD2nhDAA4YJrqvMkJu4ruSl1949FuBoqc7+1/JEBN4ZT3lpylxsKA7WHYiXk960TPnDSHG5R
0cNmgRqY60mGVgtdM9JXsVz7pdd3sZVq7KDZVRGLB8YRpxw+qfzc+RNFMRSxoFopvGBinTHIYCS/
22opB6AbSxfIW9tBv+8mkRUZvnHyjg0u9Lfve5VJTgT+rmKW2FD/WljhcsYrVXXnbN5Fc1gVSNSP
KZHjanaIXlnwGzmiRyECvUAZ1YTDd5GmI1SKT3ra85FrfPxmENbJX0DzJn6F8OaTQBCxAX6ocOfT
z7celNa0y8FKUFyuw2tOJogJaqnZxXyypReGk63G9eLrAC94FvgTkw1lauvmHdjmQkBHXMdgaK1P
Y+yiu+8buPGOcEYCGebiFtet+vZNIOs7QtlHsfl231lAO7guqTC/xptUeZimFf4w/4oFNmoB7D7T
HVCnIwNOTgg2cT1X9/iNVF+ZfIIAfcC3JCApMur2prNCrL17a2u2iWN87Gq+y0KWJRrU8JfVbujb
/6MKGa0ZsYoUQmg7Vo/btAZqdp4uHzxDmKKNokc4SGuIVPqY2mqmVXY80vD8U8/oVX5PIjsRhEjo
+abJ78+VwlfTA9rS9QvUDv/37yHbhlaRkH5rdObJ19AFK7J/AkHNKlfUkKszGvIgRkCEzGmMAtR0
tKekeNfdwraB/hKg/6S+FtQVsio1zPOt+Hn6CDK7Yg4wsly44LkIT3f4pVgynJk8T04KUNTIXjh2
vD5HxqxpWuqaUqAgKaNUrxYp/8KWEZ3M2iPXEUUQjvik13DNmG5VnEkjVimS79imcLVc+Ne33Q2H
tSDMlDXLZ0HeT05oLTgInYo380JB4n+yH/FBsHO/HcvSLgI/EWJaR4idxDni9a269iV4nJ2IAFbR
PF/LKQl4c22C5aWCQDUsttAeZWSidb7vcPPyZeOgfETucH3Jf4e4oM2IyOyFDvpBkYBN5lJjt06o
nOCj/6PD4YYrSw9fobduStiXmYwe/CBHJqWBUfRWARbgavp+4KuDC5ZMUSbF29JiurhpuWwIalt5
TylHP7VDgHizH2XP9ciNXnqnOCVaDXGlmLmP8jLMZ7r+7wx6Cz9464m0GqrLTEfuNma6R4UWzIfW
TV1CaN4ImfW0ovfJaYHcnAOX9u0SNWcSNdq+LPj791jh44atpdPjMOjO3IijY0rCk8DNbJmKou6U
vpbKMc6HF+38Dka6kV6MPe0yETuX+OKmWpHe4DtTj45XVS5sjFEBxF48fQYTwTgSCLwzn87Xqj2l
3+HX/LxNuH7G3c/m8dzIsFs8WeUvPizRuehmPrDU1x9D3rU9WqSKaNwQjwpyKKTcWSyZ5e2NVwUi
UTz5+Lj1wkqPv1AY6H0jtCzHiCvNFJFdnOK0E8T4J/RjS1Sy7TuQUNI8jwOmqVaI3lXwnzAkCg8L
B9LuadwB0XmK+B+Z7rQXBgYgVOgIyUKsZeNi1o7ko+YhkJdYbKCDrFGCTom9aa9WYSqYDIxx37PT
oyKnwaEzLJpau7PHflv6l7UP9FxIF9kXd8qwMVy6BiIL4Lt9TBZMrfuNS2ax+23ULoOxDMKEfeyx
Z1QOZsSCAUK9H5u7KYnXSz7vkKyAossvwzho1fUBWUxfsShKKSblJTr40CXw+uJqbT97nsGrDiBK
qOYek6BUMp41vfxe6bK5vPd5awpeJ7KLjpP81hif/WGXoOgXtrmdIS6n+FCIfxNd8rqHMglav9in
jUTUtXXX1Pv9zBIBdeLQ5+/+NRnYtAV1mOdzApufiK38Hk68RZzEJ4Y+sE1xpIcvNjkPt2oT2+MP
y+Xdk8PDY0xVAM3rz83Bto0FB79NoH8f+LbngBfeTf/MN0J0+NLIUxEEofn5cT7zZKIfmUAhRx3G
QzkdFQL7uxkO3Qeb6SA6SZMWFzQ17QNxVs9DvLF6Jc8aUQgJP+oGwukW2YV0FC+DYbNbdfUV+MbZ
fc62pQjC5t5E7T9c6tqpkjpiieZQf3CoE+YFHKnzIvfpIARX7jjyK62n3EgHkbr5hKb9qS12ZKno
SDt6+Sbj/Cq1ANsbSIhDavXxAMd4pkL9gO+jnmcWqxKWEJzvfu5OqArhf1oiLm77gUrXvmCnhoiK
nWOTq+HxtXfDoenMCdsu9zfIsWqABtzF+Axw19WRFBF+jA8KSDT0JLGJJtcqyr61ZPZdEsodWCMu
uiO/+d79Fg/ydPaG7kqOIh8HqqOs1EmARGpEIjJgz76/JPmgC/vZN1RZcKDrB4USADUdwGHQJIli
CDtIn9hlE25rxYuslm3ck59ofwTtDISsgGnn0QnCASxDm75nTwlCn2fF8s43wkjgL8DCFrFwkomd
bjbe0ZtsWVZ+CycQN5G9xpOQ3JInOnCWOwLO85KQKFer+lIlUg68K7Dqu1UUfj9SKuqax0z3BWhC
UUthkGM6Uyk5Ef5yDsiyUJ4+hGB8afJwXhj0411DG1/jS3ogATRwN/9MdoUMtFKLLAT6IR6lkVzB
KgE3uj0Bz+b5XemGX55p8QpGxxpGyKdzMb1Ng6SpYz2zuVJuaF9xhiM0FZt59IXQaqshb7wOQ5DA
JUvEjVPqdQ4RcrJI9eR/0AzO+9Kiq/rGgLXhBeejG/I60KBmq7a0J3AdaaKo1a5/rOpqMh/XO24n
RL9q1tWijFi0G/jTIDs3tBdOwdPtx9z0XRFPnX47sHzL1Kf0OGMIYEeMdKT5rWzilC6I4+SsUzkU
WdHoF45YFg4ae49V7XDXHLgUWdmW4ft49gBPgMVbGQGgXy93ZfwNaNsS4VVbd2pXCfcTPOUjcfI0
H51Ge12WAG+ZFLGn4D7W8IxxzBLU6l4iNbMKrMSq/Z0th9PKmOL3s9MrE1uRileDOaei0GZH7OS2
Xqe0gnj34OSViJcmG5IoSpuMkMbamXfNsjjsWg8r6KkGhcOBUcr8BLOV8yPts3IGqRo72daoulT7
1GSSUZlXN4P/fvpMKuUhzdFgclavivrZp69Ji0cCPh5bCFV5YbwXsSfgIBL+MzqPB+rfjFKXKqNd
r5BubZc1hdukc1+tlXzdNWps0sKRfV2lHUYixw3xWGLnWwo49H4tdWYp7hIgxeDPENFRcZgRAGV1
yzBy+eS6BHzn+ceiNn/EojqnDWkZs9c1HGAHqnC5g3NgchAas+ZfUU75WUh8MqarflUk/m/qs5ty
Mnsm6KyqCWTrHFlLpYcHGPXZHgBPUckicawSvUpVfN4bYBMJkYxYafjxBV9kK8pIXtKMgAMrpWg7
U6naGbZSlZv3eISuA/G+MK82BA9osGf1LqYqU2AxEbz4OqC7Qopc30tERxBgX8Qux2fKVaXo3/81
Lj/a2mxRGqLUuG2TbKeUGV74QARQc43MAbc0WoEb8FD91w+QaX7DAfFUTrEmhtcIEsV9jrh2Fu5w
HjDxlY0epmSJ3rKJG0SdIYKbk8pd86+HV49fj49pFu7Sv+C+QOuEgfvg62dukST7zsSt8zKtYqkN
BV9EG0cs+SmVKSCAk0A2cx95bcvhUPs/lFZsE6gx8RC7OkQ9a8EnFqBCEhUCXlLyP7ru3671GE1M
l1dZXPBblEmaQhhK2TeEsWiy0YrnApu+TWYAvSYzNY7lDpO1H3TcqYmzGGuU1FLcjUmK2W57knVc
mHSO6wgfT3sqbSMxDQKLCqE/vxDsHR40J60JReyEO0DHmqtc6gfwyMM6sySwaMzZmFfPfy/FVx1a
ckfaUiswNHl5QvWzI1i7QoqQB4dcqcHhl5KbEuqn8qXBKDpWIR67hTN3T29DBwg1cquIoo9Ttgza
+g3RzAb3Q6oLMLwLt490XDD9+obA438kgJbGSK8TAg5AD7mspN+GnyKhIOmiF6wtbtTSdJ5EpC6n
shv0UB/CH1sCpi2GlTBIczo0JwCRt+2b2ezvgXMyEWszqg5i9QaVZqIk1lLoo3PcEvmRqcztyQXq
3/R091DCJwnPkg5oribvJgqeEoBdS7ENdEukbb4xuK97jvPe+Q0nf4dXqSWjaZIa6EYPO/yyUotv
chTCJXT6pJQ3Qgxil0tkxBcf9GmcWbbqNkaqv/Do4tc4TN+85UBCPqwa6iD0shkbSc3B3JF1o9bo
aKcHxZGPoGuNVHsu+LlB4Jkw5ey9FAEC9waOJqsUQIfNRUHF0raT2wrerFJPJ0tMYH4h4Hf/HMI1
HZCDGRmWdeTx6dGTzVX5nY7CDygorWy/mZFs5VrIFm6MtjDYLe2vZVNsqkrsDknaS9E9PN7cH+j3
+tHO370Uu5IWv5unOlT/sIDQcOU+k+tL9S+gQWxQ13RqRdNy0Y4HBsExJI+ORTzzmqzHAuWKaLMF
bLHgpzuz2uufJNugzvAimvzlrTN6HdhoCT113wH+7S7qkthLo5WJzucdk9CvN+2+sQNS6vYJ2PEA
M4peHR4R5eWbby3nxd4vi+pzUnqC2wrVT+tqS2sFFXlaITAQeIVgA8NCU5BHaZBTnfvnCJYhtn8S
o7fVyNjpBbr25+trwlryHQP6gIF1idRhgZEO4qDQDcEmMzWY5qK4Ofvhgs/wj+VDNcSR1yQ4FxG6
/OvsZWur6lZoCSzk2G//2ZHsy7Ras1E6B5vgDZ0QV0+cRFwKx3FAOwTzguK0rfzqkfTjC15j/vK0
XVlFiyEiUWftvOpuIPwC5WU677RYrXZkP77uhw2FHVr4PARuOvm+AusV9OKd3xegxhRR3rM3w6MG
b58SxHIvnV9+6al4B0OsLVqf1dZrUQS+eLVhA+tZgQUHqdQuaDdeaq7kwEEURLos76Xb0nEW9+Ei
nZRpnu1Z2Uzv2dM0XVddeLhYLZny2d/vDHksmBgQP/LmN/7hwKY5faqltYq83PRzU43SVsbp+S6/
f2BY/ItaebZzjoyIfP/RQRKLpgatAz/HP6+hh6cf8g0THvIUOIhVS7BW2CyCO5zyKlmdCpLxu/i7
GwOCO7jywWx3aofbs2W4wzbhn2/2gp7EnUBegU4GujNmNH6GE21g9kdpueUGigajCCJVc3Bf1NAc
fDgcTe8r4J3udGmP32VKi0nyAICc8rZ7Uy1iTmEtsm0F1xCoZRBUML8mdegXauq2qAyLU1LxoHYj
h1g77S7xANj+heMJEykLKHcDZql23SZh0HSVeGth2y76mbJeOe7hVOuDl7CwLdjXndZthzzcuWjr
NLBNKShOnj9zyopXLDI+jgATqeUA92xCm/pBbfWX64rtfpCr7NDCHCgUMP7EOOrbFQs0H8H6Pd9f
yrd+Xk0/jIETbBjQea7A2HFGEQq5HcLpGYVCNKdcAd31hYdudFgVnPPlLewww56TxBSo2AmUrDdc
f0lb7wL4hhd4hR9EBlkcoDnmTOopAXZw0yCZXjHr9uDKcMKXZVMhaS765a395eEDJPssxsnyLFGt
U8SViZFayw8v6rKXbeU4BgOk+qUmelNrIVzSyPSkJeVRxjnecXeAgIzTpGX6UxMKmrawIWaqtgMk
OzBbRtSifrmPZktz50RTKj7w4OcgV0fUTpq65J5hRUokZRseDuKtivjvdwsAEll3+nsVPVMmIn7W
sBU6PMP31l0psvcRnY6Ep5neOgb12oGvKJ9qd9Sq4i3jTyfWFxY/Ymo8H/dhnlVH+obBxf3USKd5
zk+pYmLRpxeK0TqfNppY0D+8/ol68bhpC67X7ntjgMMPvYaSmwyDRhzTEBjWkjUQERG7ZKupDK4Z
5Q7j12rlnmSLSQlkP9lbBkZpWCACy3iJxhNzDZIAiCXCIXYa3v6Acle6MvzvsinrlFeSQR71KFSu
KX6cgwBGEJhN+3GQcksrZdveWS+wG/tKoCNnTEfT+dRafSWyuB4Kc1KTw+CKz+X6qjJOO3fpWPK9
Rq0oYRm4gJtY7xKbtISWn5ZIP3hV9+jIk9npl2S/D/6PLK5JnLQDc+o9kt/P2DdrCJY9+XkKON4N
4DLnMXarNzAQPW1l2wNTN9wBMgPYXaEURs/A71PSTTf8IUVVONla2OPrTk8bMUG0EGCa0hUuW4R8
Ed5ljndqk/jSRpX0OU3taGkqobKxvYE818ltO3EoVFddreuvTSigPEQAIFKjdIvcxxWb++1cEDiv
z8pAmAT2e0fubQ0jucbLfmpsxxf0eWAHQdR7A+0XHIbYAm2k5ctBEqQswb/eZY/bT9YLhqp4MSw0
hCvLZgW9fg2cGow1ZogZUmnIqGhkhphbqGniqLB6yW+jU5vqaO6pcRZbU8Y0lPpsFgijumCg/99w
+aJHh9kZsfEiKFGOjJEnRFufixyM7RRkOnjxbsTSCjZMj6QKYKz9jg7m4SQAMt2c49uk7A9sMNJm
RoBFPB6ZgmsJZ5ts0xtoaacS9cNJPBphLjmjM+2+42NBwoATjXSpBuDlT9u4eCLK67ETw+KouGMB
k7P5il18PTj5mbACfpphYqEzFkDXwd1rnUwsgSHh4po2VQ6s6EzTsQPloKwSaDIM+QUrH6woihi2
MPSidiJZ4UlLjmdZTK6NkxPrFdzn91Y4ZGHq2nyj9VWiCYyIp103SZEEduYrfruBdLpAJZ41k7WY
6k4ISW7VC7NmEdoOWJwuYpMPcBe0FDUKvSSCQhkBz7YJ2VI0/wAYocav/kfqQcxKwXFRP2RkqFei
P70ntm3RYzm8U+GKoJKgP4jrsBV+y4OMUz/yYhxbS3+/aqYS/4J4KH7+Mgl7nKlhr6hlrHv027cE
th1X1HQgRGOQUQsd3n+6h65B3XNg1lq/xfmoUcjEUGjc6D1Ml66I4/8m3/ShwmIXAmO/wH1GmqxR
mXMWYK1m5/XnMbr6vKQfCAnMabpjKkVbD+YU8ajxHGhnFfBQ/F6mHUVmj0aiUn7YMz8glW2lsEDw
Pu5s5JBa+UT+j2+v+ifHa4CwXh9bHhpkEA3A6WOVbHLRmEDrOys247dEDy6ZOn2UjQW+/RUZIybA
vT+ACljNNsZY/tm7GXULpANnG72c6cI2IBNsnrx6BpuCbVP4NbUOXUxnoRnZWgH+RjOtgj1BduW0
QV6VS0n7TKw0flTXP7cOjtLJsCKS4jeowuI93jacqs48uC/usQjVG8MVgaDFL7lkJEK2SpeXtHuG
zKpow8qaT5gufwUcPLRjOa6WNofWOhSxcTFfn/icka5/fEsn6onDMxbCGyJaGUDmTYfTt1rZaCEL
4dw+gsDesCho/Y8cs3ky4/IYodHfsTFE4kBfbLkQ1OLcgT+Y29+rkwrdA91f4o1pTk5+xxrB/mMi
GRmux2kkwdshwcAvx0UV71CqugdexyMPxKi5F2tGzUnY6ZAj7q7XfMDe6wx6kshW2vRuilSJB2Gj
X6jc1nF9B+5qS5zQgmT4eJ0dTDpCPF5AXFyaDf7jIFdILSZoMqRkCvs6LOuCUTZJFFYQBGa8Mpgf
WvUZShlir0OtE/PBxdn/sRzLXKEYS70y4+wiqEUC4NHBiUbrEfJiSD4Dsky948WONBCVdH2FjMxL
Hji+hZA/pg09QsiV0tHy0mIpjywCR4RdowGepMlQzA6elx9+VmOgEggZpa4H3MI1RIES6kkI/+yf
dAQe9pA6eDYUYrP+OmhV9s2MImt/D/GHsoQYV3SryhOOrViv14RmKR5U3tVSqEFlcJwsNjx7ZfZf
kDX1EHjY4EDsSfuyruHVPz7Q9FCiikNOclcCHcLeC9vMnLUGMK5+qKyiVaLoVDuKfCl1GPL8IhEa
8xoVQKMEjuoN7mV6KC9b4emg1y3dYag0l+tnTQidjuIEUdV9RJaga6wFnZFJPE6J/vvpKc9uKEtT
zOSN30LucAKcdkkcAX4rqV6oy23YzR4gphX5YlyFfPiU7HCLtFeW7VBtFI7WbP3hrOYdxE16IFIX
ul9DKawzkm4j6WD6RCitGWPueyOG2sj68mUu5FtUMhq1Rye/1rGc01O3MA9S6RgLSOwPBL7DFadL
epVLkBFwWzNuQezMMXyB7E0grZ7cC3tnGYttFV6FWPn4DSOcFIt7KwxVfGbAjFda69HN9yLyi6df
veqW36JcXuVkza9rMb2KUdYXHrrFEAGu8m1eSqxzJrvXAbBcuip3CcgRWyc3KvWHQapcyd4S5loz
vfWmgxIjs9uvRnxWuf6HprfyJhvYeu8n+RIdChe10DzJ7hV61TnpIjfaYJIw1PotiLlsj4ZkcMCi
VWb232IcT/8oW+MqlK5r6rjCcGWap8KUb7LheYbGA37zaxGu3MSdpaT4qRG7DhPgxvO0ulErFhDo
XChdG98sfowkYQEt0LbUZyV848aJ4plcEh5iJs6zFOswYLqAkcq1MOAJpzjJDeGuz7sB8XAP2gbm
RP4txN+J066LvurDvlqlsZBwb0PqIlmnjoxihi1prWHPsTiwSZwyjvF/qPnVHrwB87RMJiw6nJn6
HsbVnze1i2VJTXr1nZgbduHWNdPQ48kpGSi540PCFUvQYOg3SR3ejA6Gu6jhI65tkv3O0YvGVBa7
fnd2Ok+zU//GPg0vj9jMcpsoN3OOttvuKf1GQSXR/rgAtjTTMv9vm2ShnuPAALSrts/ZavTL5TnH
+dGTY2aZx3fYqujxxZJasvvmvEtj8v7tVs2G/m6hbLE78AQLIlFOLyWxI9JzHwMbm+bBYBpO9/Dd
kG5JYF/Jk3DsEDE983keFqqDiXWZDLhfHz4P4gMAWLyt/rOmuBdx8jSWRCnf33Cqd2RwJovLG9kB
/vOrzfTj4BCpVFQV6IGiw8bTdvrgMKNo2qseizIOeTkzu4GIQJtFWbl4PWa17qThbKHZiXkCpely
WRGNUYQsi4gj4YMijbIUCHc528OJH8NjN05SudGN3KP1nu+dFXf+iCpfLzi0pqCA3IccZfSCoWnt
Iz/PCV69YFspjWC31O8T8mVNpUZAs4s/hWVOLR3avbtYQq3PdxtL08Rxuu8JN2cLL5R9tuDjZIed
O11P3cZQCrw3QbuM3A9fdS7N7VTt7+jfrmF0foWRToDwIWTglP1itg0hskTVAVlR9Qf0jRjrnCdi
dxb4qNzpsQtLyF5akWnukUWkW0rFxfPSf46XvidMgzf2d3NqVh6MNupFPgzE041/GSWO1GkaoE4j
8Tgl+6jXaQnc3vz1YYrNQZwYiycb9cHUEAvfw7btqzvF6M/ToKUe340DYLQeY4TpOujVsFZp42tn
vHVjMEz/n6ULBmpjN9eNgNeCrjm2gTCdXMA1pyDsQutafeK20ItldUuHM1hG0hdE4UKd1kbLkc1L
KFJzu2qsTZk2eLYItPo+N8c7OPMcajlBzfl60Dw6cxVKPWdggb90osK55+2VKxDg1KY36PD0BWnV
97D6Ent6OsahVq+X83BoyDxxtzQ9z3I7a8hX0TuU11xITFVxjJnj0v2UDTH8SsGij6x/nR1eBwAM
79x38wcY+np+suU70mBZXRLWN1uS54ty/Nm7vs4JwUmBM2C4pemTOgmvS8UwGX2lwdWZbaVyfJuD
c1X4GBkKNAtZDvAmaEjp3fgnteKSTOS4dBH/g9RRSuXSgv+v96kCN3OjKxZ8dNNShAA5GYSVnbw6
nh54jHDPP/gkdtfKIKCO5fAX04VRg50bjPxYEiv2ix5m0Nc51k0VgQFfmP/3hHn+yCgL7uVegoQp
Q+vpRjeJLSQ59mq2KUIL0mEg0axDz6eCRnTQo7zfwM92lqvyJ8VpLucOv8GkdjOldqaBtDCDqbjM
Rlxt2DNg1W+JKhzb9vVsiW9jIF9tct0UjbOGVHWv9iCHKnrmMo/2agvGX+HjaTt2kQ/6lm3MBP8u
7somr/liHUpywtPCgOEDhjovWlOO71KATZuKeRDnc0nx1dipK0LS5GSv6kvq1QWE1cZMY/XqlNQO
5KGjumyWHgwEWjEQ729DVVw/EjbJ2p2f+4nbxjuW3kiwMge9WS68KhZN6Max1r16U2aBPIK4mFkX
dn9VKjl8bCwLd+YaRV5ldH9vHRY5lxWYcoFnxZ+my/jPrjTf5En2wNtVAM7OD9DI6pTPw4WNwint
Qv8b2Z92lBw9wtCu+WVHM8fzajQHunu0LSXQ6osCs5m1BDeFdrRAfhvPicj/QbeZzpSNmtUClwg5
NsOU/HwtO0cZJMj+FjJRr0NdgJzp1SDyXgGbIRBGuf/swtlkWEgyhWjZDqjy4gv3nFyBF9XsXh8l
V6TbHEWHI+BaNQWwBNMTTO4ih70tqusn7HFVDNFxdDpuDtFJRpkOq0aCRy5FTf3zbqopkYZoQvHL
XIBxHucXTUAF+SNShKJ/Ki65bDwLOoFwUMTQX6FutMfS4HZWW7d6UHxi1hCNnPa6zBniQFWm2F7V
+u9GbSsMbZ2+QUFrWUiPbWnVcKSKMZIsFzg7xD4fNVPmMQ2BxpVdloAmlIIWQzo6lqCV84AAKOuf
Ngzavhqk1jFgJelLTssiMMezMYuGD4WMLisshqEbbqytHyYjDmEymQaJ1ZaN0HTgvJ+vwf2D3r7J
JeHxpogoa8/ebNYMIZrJjaMN1Ev61QR2jMcKrmDs1uU9ygShXR2TTrSzKG5PApw52lNAn7H78NZx
XZxKZjJie4ceuysrG+2twGc9/6e5+hvLywF7KufOYthrwntYWzfWJttgUix+vacKErma8ZyhQ5lL
giIYPUke1LYBIAFYX8a0yZnka3lGKSt9297jxqwAwjlOb/2mXiuJyerb6eG2cE3a7yIl2XY3d/Qm
R8JOMulurjJlkEr4kTufMHpowU76CojAoIBZcpl6I5xok74XDB/QeljgJ09iYwxd3Fvj6/B88+Q/
oHKhI+Jw0msK2cQO2rUw6j8h1SWcqyf6B518Hysntj0ezVIaOmJq/EmtYRYguk+w0Ri2yaeK+CN7
AQ6PRC9eJ9hAIgGkafxQ+ixMebRK9UN6mzmp1i1hbeDXsmsg7dBTsrrhay/O+efmX9Pm603D4CKS
qaw7HMul143g8UdnR+qWbcybuGZe6hYiBIWix+Ob3dqtiG7gX/M2TWnmp18FxTAetfN5npt0NYb5
HKOwrVomxGNPeoT8bhqONSqEbp+BJLNStfbtil2O09bXJO4j5wszVOc0SDexXUaK+j5Zxg3fWISq
WTUKowvmylXbcE+moHkXy7Zny32CNzUxHZKGrGKoYdXzTl57UhjN99oXqPT8/R9NW+BIQLLmlkYZ
muwv8EEKq+OLg5M+Xf1U2K0Rhu34Dg1jH4ae+r2xKmir79QLW6DaJNQ+J5kzChx1qfjsSO92+5YB
Px2mFqj9dmc92C4F8esits4RiIDEmHHczJ5fUVdB9P6REt5RIu58CEETCAry6EW034RGpWm3nijN
weRTl3zn5DjcbI7DCVbY3psZoaPcoetlseaEwRw97gu5PBK2yY8Axx2paprEMuJ17C6y9z9TNS4F
/0PIohpiteIVfFM8sV1tbfdsmHRJSPeRToLeqvzQV6ge105ZQFpNB7ldXmzUMwhC3craL5Ov7OOZ
s0acH8uzb+L9nS42g44XNTVt0WxwZDhNN8rCk1ESRmZUvyXeYKulUcbYUYcRZbXQOEMD0zWeqlrH
OFssleHd9DJvEMvStktrx4w+vUGb05e/aASNWJiCIMct/vi1sgRr01MROcjOjNiKTlqLF05wyLoH
URWRjjqoRRXY5xv8wzhnEbjd+merZsZx8bY5PzTWtChnyCBathJViPHDzHjREmgFfw0aFopved2a
RsDGVP3Y9atRRzhbAwYwy1TTsaMUY7W2a/hvZlA2snSunw9O5ZGgyDCb/Tb04lK9mTi40Yxtdrqn
ZOcpEoV2DufRnasCH5a9xfAO7I9IROkSaLSh+lupziJR7Gj7TLyVJHnHFsnNjicuJHqpRTN6hBbB
YAeXJQPyTp73V1dmGnV0Vs/lmKoTwE/0xdImYfZviJzhhOncdS3p0RlpFXWwTL7xRUZAchcw0cvt
R7Z2Zx3YTDuXvwFrIi8Gg86wo799jnju5cKiOzHXC4qZh6wQQjYvuIdBylWu3ftoFusATse/nY3u
FgjlUMjlFRWtO0Pu8Xx9GWZUyxUv3lW/7VxFZNbhuSv6UQT4sEJLdePhXuE8VCcrxrxYfDEORW3x
T9tQnazb6dupXfbmDTnn13zAoZcAkmkLpfZlqcaJpNzllplA5KSQGH8xQx+pGicUW1mjWBt5fRSk
uOVBRwkEUcUWXvGFF4/DVA0Mx7bjkFpfGkoG1pA/la8uDopjsNBvv+AIxRqvp3GHCUy9YsbULKc5
FcjcrK/V0uBNntXwOr6oNSGteLbOF4lO2eOMg9KCKgFK2HpJdYw/OMw9ReFN5CxTZcDWSpP61DbT
7RI7tQDj25l2EXfLm6jMnFIWICsRGI/rZh1nnVMyN64QpFVqjL6rjpBVks255iOpX2JGEA+zHmGm
mmaMVklPtftx2rGQyzfsWY0FimkkCMJAmssRlHgy2fp8/j7aBiOikBfDoCWFpMK0QT0IQSQGsUrh
q0yXNFzvZFC9WBQ/AXfUvQVqyj/+h6xSrDjJ6eoF68/KBm5UMFT9jLA/7Hd7gpeoeSk0LP8IBqad
Y4/Grw4uzjPhB34zJOM3jpBZuUl0AdjosCXJwkIox5DhFBjqBd3gcXKItoyXEZe5odxZQE9iA9Bu
kuKXd3XnFsBwvcDjvJAlDJO/aq3N+K11261sBqVNrggYoDrifjSQ7A5bIelDp5oJ3KwgwhIU7F0K
1J/lrHBy+LzXviIUaVgK7ZOWgeeInOh//w5D5aXDYCTVEM6ZeMlQ0UqgK1xJvHRG1mehpZ53eMpa
ZzUtMc0rkOH4n09IYkLgv/pT/cf1vK4euXbPskKTA6xeg9YwhwGvxtDAkgt8LoB0VMg8VHLeL1WU
Q5pYp2V2VbjOqjl+mtcac+5iu9hZdlNS0dM7Cn1G6Y1qj3i4BCqIOyjiGJX36AFSJ8Bl1bBlDYEC
jo7VWzDNcXQR9k2/tQ2c29zwg6d5aaQkY2HsJFUCBXnpTtH8D2KJ5TfOFqYdWm83nTFg20hrI1Qu
VrUiLhLQL9SEqjAcxNRBhYxP+flgIhCYH/eBSMkck4m8kB1L057kb//ETG1YrqnrlInkxVCnwy+1
O/r8huaV1gwx9FR5QTiGyVPiKDVNQHGgRsoaN4Y145Hg6+p1JmtT0E8TFkP4iAs2eTGRUlc8IGN6
jkv0iJwSJtsFdiei7BOsucN7b7wiX0CyehOBmaHD2HmWZ24gyQGsVtpFmG11in6NC3TcvzL0OAah
6RbtA2GFBwUc7vco7BOwqLRCWmcTfQ5owSLshOUD3OGKiQTnHbNiCCljqvCfSGHOpQwF6i+B1+/6
QvUa96vAbvsoa13psFE47oyUQbTQ6VVC+SKwYlN2wKQwzxJeK3QgjlKrHhVAE6SieoAZ7suYLsoH
Wo49GaVwI9cbrJZlTaGA5TQDUzed4YGlqns/1oXwcC88UDTFBMjopsZdL6P6cwoQPEDnH9WBTJnO
yYaODG6CudFG4S4Lg5NCNv4rZuwUw/HXnUcXiwREH+cLy6HsIgVi+EVfQ1dO8uNvNRd0LNA3hASw
ly0BADxh6QGMo29dZ4y5nh1D5dbRaFHYPUY1ltpuwguMRsss+gIvxPgS0RYN7ad239az+2yWqM+E
RkmL7BVX9ewpdbeUvW8i4kPXI7rvORC2i1I+FamoaowUi/xjg7+0FGe5FfRtLdJqpkWgwJK79k3p
mYSeLkHfxouIOw01amyHg6uWNUa1AYMNfUVqf/CUu+BVstViXPEQaEPuxQSxR0o2SwNmvKxo1uq7
UMCJJ9UUXs4lQalDNhUmGikKXFFzxUyHpTgLdI92zwN3vIpWPsRMhhr424xsMbj11ayHgYdtb++W
UAj3S6quoObagcASCEZepOoB4XcXwokOi393KVSbJDd7GhSzjEgtPkUu8aXhjGnYurTLpvwnlT2q
1ycxb4jN/lKf1a+iUD5OiWQLBNgfkn2bKYt53yUin1LWNh0nJNjHfw0d9tic7dO4Scw7bszfNGk+
p+tMwIHkztaAHHK/enQUwYDcvCPIuZ4Pnz/inR6svQbhJEK1K/0mNRXmPZvoXVWN3suNo0cpe8Fq
jGlZZqfFkWyJRgeCk7X9YGcl95XWFclcYW8ak4fTug/1bVzWR54n/oNUcsC0GG0Q/bHiTnhIPinJ
GJYqDKO5GUTrT8UVGdJaNVjYghHQey+94FX8GByYI7pjRSmVA387NAeETNT2ScX2tOw9FlFbZdKg
yjn97lJ1ijKLRklcHiS/eSq67JNqHIvnY3b12qwOFgZsZCuJqzAf5L6hn5zXeZot3AEaEn9TuKv7
J8OqIqZvSjfQXJC6VT/adYeEKEC7+h7y3bGZ7NhwUqjNNEp2HHMDnHvD73J64Ap4vzfO1oTgMUNm
L1Jp0hytB4dxfbn5+pnez7RFuKeLFS/N6DSLwF7PAKVsNoiHzfd1gSHFqR5oJaWD8ErAx76XtSXT
wDICGR3feOxUPsnCSgt1ZqTXlkn0v2tbondwul4keuTJkkc9aIHjoFs2sG7CQWWxK/2WLU3Ry5cH
lHMa+O5etr3rZpHbbC64mP5YPiZAnvhVDTkxNwLGOb6FZd5Ix+HOUAuoiMUgTOUh6WzvK7B7uvGW
mNHqZ6m3dgSgR7lnIw3xe5XBmCDb7uIjkddkyO1znO0VLx+JX0SJFyILQfb3d3SeeTgE/AQ2IyII
vrv6zuqV/uYfH+c4+hzr0ahksHLdymGjzDV3rz/ost172r6wAhxepBM3YpKRaZ9+ygG/r2joGNF6
Cd5zHXqpwOw2Sc7YJRZ12bHazNx2kd1TzbTLPGPnvGlawhhrRtLE8FWl5YZVlLdrV6UHqh9dBNkw
ToaVsps4ZnkBHZDYD0by06QSKd0OI+51mkDNpt+FF/+L/nEH/0KIDfN1W2GuKNDDi6fvxykCvinT
WyYuT5NrMOoRCp584atzMsNsDMJCJGg7hGcKymyD9X4GX7AOXljaLkh6ysozW2VrPN3sB3U3aQMs
FyURXnmbbXsNaU268LHj8Woc4SGoPGNvhjMZZeajAw+RrCCuVGRusl/SgH8pMD7IVE/eVe0dp8vZ
No6D66lWwyO5gDt/FjayJHYaN7u6HkS98Zg3ucWWJQ0gGElzdPPwVa6YRzoirAzTrLQpxfoHZsyo
08kXrQOQG0Re7lYosgQrWQs2fWoFwcCXVb6WxKuex4VDRQ9moVHPiDFhgOybVrdduI0JC+Q7e8e7
07CnaRVCVyqg5WQbms40q/ShCvMKU8ymjnX8lYYooknJwtCBKFgg9q59c8shlWM/zVgGibgRJ9pO
xzSWYoeWaDVowv87aVtGZYHCgtAWcahSqEbMl+NTy3vogK2mSZwdLqY7pPZ+6Ktovrn9iPXi49oT
SDtHLXm4bMjHZmuVdmGnXBG4oa0hnO7CQkzUjLOXryuJ9omPIyaP1GlAQjRPSJVyAbEmcox66DWx
QMKMuwNjE5JQy38+KFh4jHQwgvHv/K+dmvpL8uJeO1WdEM0Vc7QlybyHlgg1cH9AuwGYnw/LrLTQ
5cQuUE+imsJFSoLDu3iJyT3Ff4/gXZ3Tulx/DefDybQxPMo9HU4o1YokhgA01KvwEoPqbzZ7gEq2
w4H4Z4cXt0xlDwZQEUHxuITF3H5q04g/Kl/IASyqiiJXOIDphzDHxA7L8UgLnhgg4vLXaYXh3PTZ
iSsWvfnXKFYnw5XqMjWC27NjnqGmTO0WcCg64mpKsfRQ4C9z5k8mHcDC3En3CDScaD2GYIFViCGo
xmlUH2gxJ2B5lFzRfqCtl/iua93CM3s77Q4kRUQ7JlF8BdYAeuB0mb7k+aKM1lhN7NHlNvBdbQPS
rtUZdcCvJUVoYe/z+ikFfX7AiEQyv/1t/F9QSmcK/Mxqcr9/O9RWPGs+NdRWhj8O8SCnVeOk7Vcu
oJl0ZWXFREogccSHWSe4ioWx0yqp7ugbDkzNXxvuBGP1uYdOn3dWhKIaxI4Pojj8Fm05D03b3cBJ
zWrokikqg6iO/UV3Qti89v78wB22ptGVx7TRHfd2l9ysJtoTvaeLm8YM928sUMxRUaplImXbAs3B
+jjc3tSDi+SDg8ptHlXFY5/DJfZ3RRV71eSe0S7gc/uvCogpfDLoZuZl8N1p+OqSdanOCPhZU+ev
pUc7IoinTW7Yiar/veoIYo+W+zKLl4hDnflV12nuJsDHUv371l5vbdDcG0xj5slh5c2N7K7hjADC
t/o2OPpUxrzwtSbo55KLYt5dfNz4jYqX+dLUkYL5H7VqJoj2BmWnuWx15Nu+7aEbgiwrq+PRguC4
FV0newOJZEcRusnNH7hchK0W881kmn9XGWkqEhcIsAG7ywvh8gfYYa43x9H/M9Vk/evSOTaxNMVX
fgLWaeFWkRpMJPyyL20I/wI0EF7cHhkwCIodyGTY0tKa5aIz3XEVRnTJmgHMAH+ByrlXFag2yD5B
s7O+CfdNQazHtd8/m0dbYbN6l96CVEPRaxHHsn28szkb34YDbuzoM79frlXqG6QGoQEXsZOD3KaT
YD8bEDsXpDw0md45NSaG3sKle8u5PBlRc7j7YzIASVmaBNzp47SFD9Y2N3B/vIlTbnFQfi/H1HCn
5jY6Bd6zcEfCch1ZXqsITg+gA6B+OlzwRSRnQhTcIKM1WOcHe8MY/cVIOJNMrULhxylaAQWm/jjV
zbExMDXbf24NcyX+xC9abBVRE+WuCdtxS8drb7rZMM+cTrYz5UPYWw9krXL41aH9/iLQLzVjHS/N
sM45gQtpWyjrUJKxHuXxbneyuuV9QVzBwPTdBlao/xn0VgPPYMWl+kS6utCg9jm5vUCk1y8wDTem
iEFJaQYvaS8dCvBqXTltyyQrhrRgHadsdrswHLthfi51E8HQizlwLtFD4vKldzcF07O06TNF1vg2
jSRg6SzEI2kSMHI9SsIjvjqC4rX37SPa22g+cGQJX8/tmi+I78flCw0edGjJ9xqKjiJ2pNWHPC2T
CXqG+VX7tVDWEB0/8+QJMc2/rmsPVpEA+b0DHaECPe6MojaCrvwr1ZwaPvJxF5ldb206XRxvNmRb
6hiKya5yA2tnlZIyUmdCcDMMVNHUgziUXg/pFTAHhtr8FnmQGVOb3k4NADIlc5ynSj6rV6y/qZjq
kFe1rEjMaDWZB84tyyDLtekYLXXv3aI3DTbI1UR0K5AJ1LDijsIhQWB8d0ZnDzyWQ9qkimZb4/UY
4ztN18BtSflF4Qk3qffU0JdIWniMAf8wLQ/Q5g/HZpN1BqzEyASryiunQWaXbRRtAw4DkiMDN7cg
Wu+clIg3YWQpaSU1tEnJt8a4obc/NHsPAB6CP1y0zvmkkaPcLlKimpxrGdOg+WJ7IxXb/uzwifqQ
5j7amcjKxSweSeAYloinb0mNOh2d1LxdKw7ikphoX4t6ncYjdKS2TaBMe6XgzsqXCQKub9BQ5X96
s+CP/XBPleOEGQ2EjLbfznvSvA/LuJ/XUBYiz5ktZNx+kuQT3Miqncbii1rQG42uFZ8kMxAkRhie
4dlLPvpDa1VvVntq4lRLLfgXHhDJ7J3N+JuPBSxC9QSCBmzmjEYwWziFB+uNUPjB0TeLvru/et94
3r74vn9/6IOqO2e9zFTifsyZPT+6RwCpc96p4UAvul6rEL1bEwZr3pUfB2lHMsN6bQ6PM19GkLXa
7Ec1sRlI5NtubEaPajV+6N9wSbHgEIYrP97PIcTX8a9yML8Oz4HuKGKQXgP8kltnyyDZ2m+JN13s
PgS/ASn5DgLUYrx9EH9XBhBJQrhVFhIzIK9IIYbCjJfwxcY6H7NCvKqUELloAojeu0h78JKvthog
IVbqqNv10aN7Z6oOtEuH1kLNSYUYt95gRwdlbgFuoAeIbTJLuHRHOji5V5NNwQV0b15xdH+/PoY4
CVfUgECqo55RIXs43qsm3cqXnIN/SsGVQHc94mZUZs87dRUKOoUe859UOMIPJM2y1fo8n5Xem9io
xmMp3y+Amoi/70W+EjeUATTv3GaUNJaE6HYIkHwF8TwckdeXji93WvVugHrh2p2XocAwTUdpAqjY
GYyenP7MEZtkHQ6gTmy65XIRA680x95+jyqTGVoLvoTcWWTio1b7Uj8HyJHc7YdmvJ7/wffI1XzB
mnhOykbqLAssZutZtGOMl0S0+/W7ZYYtpyc51zs1yKZigIRtR3dpjXWHS0/FpiSdBvx7QU2WUl53
yAYL+UPLZKIauWnyxAUtiX59Ckr9Gbl7UAuNjCvxkGi5CA42k7py9RnMY5O6ft1dw220dIA/LGqn
6nk3CqVRL0ouxdZgRlqJrp6bGDBpFET1su7vopKDxTBeAf/pMmUXYFtYLMxm6rtx5Y8bbd2hkVL4
WY2Y4lV+cUwAMZaklNVUVNGMVAr1wt6NbdxQfJBXgGcpCkZT0xl/d8+Moa9llN58NSS1S8KK1cJF
nhqoTx6U3HdUqqstfG35Bhb99mm34kCTm+QlsmZymDwnmWTNtY0vu62Ptt7QZ/Si8L3LYQq5QYsH
++GmRZ6tFRc38kP3Nlztqjz61mP6ER04eJlcXHyndBdeKUYTLDGukiqzeasuJn8O4+I1Va4g2+Q2
W4MZSty0Q08lzaMP00kIDgqNKy9Tv6QxfMTwTCm8kXoXdflGFxsBLrYwAtxnQISs+LsrHoz9Ybik
TgvEG39LaJaBMbo9+tgxP2AGmowgJ86RdGWcS3jvN2azMQr6CirHmNqaWWVBZIkbBMCzPi/cBTi5
gHWddOylf0R7rqpCSdQLSkxlrw2bC87C72m8w7zN8SUyYK/4TF2yIxNuHmb5Fg153FNyZQQkzGLe
RsbdVXU34fY1zPGsWIy7EztcoVxFnOhG36fTCkt4OL8W4aaQfEpnxdlgo9TTOV5Lm9G+WZsnpZ8Q
abL3VHGgwfiQ8To+G+VuPlAH15H0MIyXY2NRTEUaxu/UUU2ZNl3ZNqFtxlDKqrt8Y0clQk+YNUPU
3Tb9OeRmq5mL0NBtF5aGn7J1iK+6OWdPJMRdVeTYjzctUbolWDgcaCm0rg9NUW4fRO+tOxiqs2ww
+fOXXd2P+i2qH8zLnnspc6hZloAqkBW2RUvhZ0mJ9DVUAz7yEuAeYQELWMR7SkTXaGXSQVFCJE0o
P/G/XkdJuuEuxD/6cq2NX0XR15AMOKHsEWZH7zU6GA1eb0QY9fYJD4hf3W1WIc8+zaVLBgfkefGy
BDjyV5EJLtYgqGpx6mqgAjYgwlSdx9OCmA1hCsepX2I+IlpMNMD8b2d0IdX6Eci5FwNkkGWrh5W4
6RUopd9t9Wmefv/T02Qbel2tWbKxo+F9xuUetOMhClra4aiyuI6AcRmjqSCcjkWvucx2EXbR7CXr
C6cPIL2Zx9/b/4aRShlCeXF/aI2HjzROsMmgv+nNNOzaNWwu76qTVMtJhNbGkZBEZYjegDiRb+5l
CKuHs+4W2h8lSawZOm6VCu4OT75Oi6MCh9MyogYcZudymBYwNwlCMANjuynfOa5TlYoTKEdixn+7
uGQ9MKoPkUHEThOEMP3HyDgPEnAN9i/KtxLohJSzFVhBm07gsXViM3la7VZSlqSzeoMvhdSFxfCo
jjtqSh7wT6q95ZBZupY/kMwo/81mmN7TaFpof35h8kM0ZQY0tP9LcP3bNKc8Sl4DDvUuDQmf4qv4
a1dzyL0sc8CGXx0G8y9uxQdltkbp09MA9Ur+mQ3MTp0OwRC6MTMEpcmG2BXNknHI3RzZAyozvWEP
5IflouTqnJ2Wp7NXV3SNgRqGSYvDjhiRW5K8CMANaOHQA+pLirOGPTAwg+hkdPK5ql9TJ5pmkgm5
DwSDAE4tW178IsJePuAXTgpnl1bxxHvysdfsBtJoZTKJDwM2UDeLzVg9kkg9butWjc8qjY5SbDRO
W7yGqc+I2B9KdUnH77d6zOi+67hCk+hUHnP1DOiDPhxqzzavvfD48mMB0OyrzfIWjHUwCWf2yf7l
/cThK1hFzCDBNLD3kmO3VsnEJtbUbi+sPVab8+YOtfM+5XDk8CioQv5BGBrOYKDX+fE1fEjz69F3
gCfSnjCDQS2SXf3cfws8G60TqM/33JkPa4ZoexJAOzbCMLTxZ3QTHejsjxhjo0Cw+4prUStdzrGL
zyws5QMPlauxQ61NktCz3Omy2gjTuf+hObdhnmOvkq+NaR6dBPJOjqfgKRbNSqpKMM13iSfURPYl
Jbn2Rp16WIVs+a4zHj+8aV5q5OiPfjsq3stq+NtdhujUNH1wOrnUz7rsNX0coBZK1vO43lkM4Kek
4Sw7QXOAlGWltP6pFp4H7h9OvGpNyrz2wCzEc4hYNlvJAUjahyVpdA4EcJXzOorcjCQgEoLeZCib
0pn/CucwCwGQrGIsbLaEpw9tmzVLjNeHKo5OlcTR+VYn1HM/QefbAOuIInwFka4j22mlQEd2MTCc
08WEaL71G2uEylN0P4U5qt+Eixc35rw8Ek8AEAwphZ9jvLrZTOyFfc9HD4xtYVkOFJ4I0kJkZOxT
i2A0IE1iISo0UQKDwltPcoEYemb3PInVNc2ShWL83MgQOgsoTpGGRjqciF++tZgmzTi7vKNRwX/n
qdiNiSyNyYA3ZXIk7/sPj1cRW8Ga+zQJoDPkLkVnQWZwD6cd/foPYEclMoK2WBlW7aQxLPXAg5Hi
XG34kp5uxr6gBFPF0pIC1XoC4kSGAJKGYXko3Q3isKZIO6Lm6Vl9HfSIBEk7hiY8igPkZ4pO56aQ
+Fmkg/dXj2HMgJNVujicN6c3iNPLnF6pGiHoDQEFV/NHmMxZEXTNyufglIoZrFJsvaYcoeq24yyC
wj3uv/++0jn3KeJF+wVRvgyeJtLwqRwCnOTRLXgLt2y/M+31tDRzDcNCBOP9QrTGMa3oAzGoqSn7
CMrdEOmEzdIaksJniQMDBpzgsPjnh52D6CtwIFFwX1Gl5LyLcfDVNL9E9xCI25veUWrrO6bqupwQ
j6Kn8RulE/a5JvZrrXrKEOYCd5MECQWljKTDepP8+GoWA+L4mT3ITpPBccnkaUdVpgchYeJpIeW+
a0GkGl7oU1g2ECb46EyGx+OeE1cLPpuvWBogJDWiTxlmVOfoOTcFHdjRMqk9vL8gVav2AcJY63mr
q8jDdhuJCot+O8+IiguFSDXRQL5MuDR6itG3bxxjcCFrYj2WauaaSs6NafivT7sqGEWGiQmKbGx6
r7u93A7C4CY+kVH/6SqMORJ0JZpEe03S6EW3HWUFVx59a/VoSMVYO7ewrU92pGjWa97ZXdOgc7rk
erftqtevLmBDnFcLHbfr8r7PdybTtP+QDr3XDEcVjoSthbU+uB8zpUIoY7VxNFJrrhvVmP5KL9oT
BRwupafCnXrsUpNhRCZzQfep61zUIv+UMLUm5HDumQr4lf4XgBfNnOqQkeYO3ZHkYVngzEeEeRSn
0SPRyaMSg7sbvA5/MTp2t2Lje+K6+xyT7PRPZUHENiQ6Ib13Hfsv3BClCDB+QXr9ceZnE1O/EsaH
/r54ccgP9k7zUgeSjrhqLhzxQgxEtqofSbXnHBUEJuDfFlPUXghJ0vyJ+8aG+XQb/LrX79O0gymH
bSL/pNGxjEdk/GG2VQLX3ILof0UvTZIkK7LqJaM9bUhW57w8ZbDWSNrVzYeOmiOKgs8fmfjLFJ5E
VwzDsuc++YPZdaJVSOKAh5DAgp+psa9MW5SjBz/wC9BxMMpkQOH6SHRlMfKrJAnsKgvtWOGTUQoE
dWUjCBnG5EemAcSV//P1oQlHqDkd74aMD61H3zQPULodVxzuv86a3rotkxQgnFY0d0IommwoMkMg
gvQjOoRBRhcaeFShRj+8hrl18Lh/uzkxXzGk58r3ZLLjg6c8efh0e4GjK7Eql3jZ76/RvB+eb+6J
uaPJ010QDWp7b1cjJH4PLm7euSGNskl2XR6nj1UQJ8684M6luMlu3JHQauSIvCf3CxXnCe2JRj7Q
f1ihNM38W+5uiT51OimH3vH8Xdlu9eugPYT+VQ9zT9vlaigduZYH8yg4tsBGUuji7i2G5Tk7pQR4
UYr+UESTw09CbErRC4V7IyW8mMCFObGZsTiW81Q08FcgD/tJ47fHZZayYg7CHu5CQLZF+VbuSAGd
syUxDBCWjonUKm2+8YnVJmMqnmidIQzAtn//aHVtUpwVMcGQZ3nhpj+kJHkyPKBCkDjFn83fH9Wj
UR2jCtzBbJZRJvGptn77LO1lpd1uXmiazTp6wu79k0PCzEAs62yAZCsz1yzIUB9OuLbpFW7AVE2l
gvhfP5FFxBuXQ+XLmS6M34nUWlXD2/5JPzCBMMIVUXXprA46WGG38pNyYnojaghn4HPm1jzu86FA
GdA64rIYQdWCl91XIKqFtnXS79jRtgLp8eDcPs4ufV2BFiLwLrdvF67CccZj3A1SwIu+vgO3+cfE
du99cos37gIj8HE48SL9x1e9Mdjqgz+dIY6fwOnzLwBj3MFS9JPnhCu2E+vP4jO0TxrRjkwKALl1
oq2JhT45B+VgcH0ECp2zG+/i8n3l+d1Sh9p850j60Thtedlj993ED6ws7ryoYgP54stma5ISN755
NvOg7EU/uG9JcmaCG/+iT8V15AZhIvL3f0rk5gRJ2vkX4izZ4FeAT4RmVCzFrhaqlstKg2ro8lc9
lSImuxnorR6E/x/gP42Les3g55Sb1P1QGk4ASj98c2/7nSG4Gas2l/h8ngZ9fZT6aPP3g0TJhJex
zMn9B+ZIvuiyrFIlK1YCxVyJluDoGypskj8cvJIMDjAzqoHnLvgbgIahoWAsM4nPpkRdBFvIYReS
zrsC1RYe1v0FbtMFnNTVcD2XMLFY7pzQsgh2PwXgTcB5K+0IHbbOxnlv+dwosD9Ykf9li9dDx5hE
KTJ1om9Joe2yro52JszHizvs9tVnJsjvjDZAsDxTSkUmr8HxdrsD6/bA2wOQwCvd6ODA0qT9c9W3
Kmi9eIhzfJ8MAjoyI+W3Om9EXz7NtDpyqxokD+7KJCMxd30I97gUqy08JVwEHEYDM5COZwtg1Wfh
tIoq8LVnOKA70/o57Jal3S8DoWbKXKWYMHMANZcvuJkSHobjJtZGSrYE7bYPOepyvmEFa4dm1Etl
Q+7xi0ObM7Ksd+75WlICtuF5xK8zKbNmdBbISVczhtO85w9vN0JZxHWOl4X8aRuRnG9enJT+nVRm
xyvnhpDbiWdbwfBOGCCfL2ZME+CIlpTiy55MC8FXEjA5cUnIHNWFslyGzsryRrARmbZXzg/RZKE7
2vKrvsckztwGPHORAZLUhcI2voKexwm579lqTma+0uLTdJi+T45yr9ZbmZcJ7irqbvWb9i9oVxQn
jF+hGdhg/yzk/9ZgNp3v/aTAwGSckNJbdX4mimYVCk5bdFse7Iij37V2sBribYua2QDFz5VjJBR1
JuQGY0gFn7ZmPWtVfqaDVzDRwCkjQWDX+dIWnSdY5GhyBvFLkife9HXijoxZKSgk7tFS9ZXRE2v7
FJrUnLwxVJP/Gbhd5bbKGla4D4krAvDfMNOdmeudLVdht8GP7wgdb0i3TZLClVc95Nr8Tk69iHVK
iia5y2ZrK7fyb6F4uoEgbPvhyOO7bCDsPvyl9cKAbIDMxxd1Yto7Sf5dxBMqB834fpYPMYsqoxnV
4dSJiNoGg2KGHX3GMuFEFwugnQFNQRLVxYYBeQ/P0iio3VGdvgL5uQVBBgX7HPffRlNW3vwp4msO
mQm5D0IHJDrxUZMooWxaZNyXQ5zfbVjoYh+nL60NLWcLZQkS+63seueAEP7juiLRyHKmGki2ZBov
BItTEgq3Myx4+awcpmL6Og4dPKAE48GumDSctMz9bUvQyAL1PvSHsLR/gboMm2ir4ep5q/rcbvtw
qR9a/GhOw9k7U/pZ9pFf4Z8PsM/PCHZFyNF1zEHpUZ7kKZFnX6zjpR0nSmBc+JYoOTRcbem/V4/6
dIac0IVyo7tlKzRuUTpoo6bmQvImAWzBGASF3K/pb2xiAOO8RLyT6gLoOXaBpsJoIpFhXisGEzJm
7B6/z5AKNcJ4YUYVxR3rhd+OzOgzWGoYSshtnG+F31vJgAJLVCUNWiU/sTH5eFGMAt5B3YMRx5G3
EqUHf/pJw65vakrkOJwyRxNj9d7zoE3Ga/8O1hUHK5jyhL5BoC5RzTHS8z6PSbuI7biZX7bSIHNl
GI/nAKq3cf63fEqdPDNgsd+u64EWOtAK3AAsc4etQFoK/SbbgpBuC1HLyk5qQ1T/bCEp4zBCRg0e
B7XnOn2J1IP+SwTDvEZjC03EYqo6tEhJivGGwx5vkOk/v9OxZ8UDtPdAg1lraEaKn5KYxHI2QNc0
IglY7npm32yRCqYwo8ggFe4fS/pgcs3HXmE5ojvXFsNb5dFE3eiBorrDLUzg7C0JplOTh/u4mVbH
cK/JSm0mDf37cdapTUA4u08YMKD9IiejKKicrBiltQ9aJhMIxsvD5Dp0ALPMMxK9UImqcg==
`pragma protect end_protected
