// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AewMfMlxfLOhw1QtUmmXzCd3EBsnnBslInFriQendu7pMZMxyMHLw1DVDscI2PTS
QvZi+VGK8Z7mAFiI/c+qY7G6Zt5PToi1amm8HOG+aUfOPl0wbDnj8FEBX+j/GPnH
/SGURUFOFt+1po/PGDjpCE8KZ/SQu45Sz/IlZ3x5t/Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4080)
E6zThR8fUzDe7O2n9nGVMcdx3KWAyaDIgA3LCndH/dUmlvcflxhxjKbIx6/ygptQ
jMNWxAjY9fnI07sd3QGT11FxGHj/XOE5QG9uC3EjUhYCJH6oV8kBp/Hp/d5v5peg
rk2p3VBAJake8CeurpaoHllfliHYU8FlFtGECFw1wxnBWWTC7IZR0+4fon/nx4jI
aMrgYl6nsFDJPLCK0cwk6WxXrQoUdu/opVmIPnjYnDkhBsHH98Sd9W+pwoG6Cqss
Wn9OmfEtcEijIkoLmrmkDR7Mu9f7/pnL3P7sZJT3tzB+4muIt5gwz8Mv1fqSCJfK
FO9VS6zc0nw5od0fmibK8HUqp1J+nDBklVFH6OFaXBAOuOsSPb9DnKO5sNOWrNNx
pg934OZv5Z5y4tGQg3XElp1j41p9Q8iawACC5RHJxk99RiO88rA5a5F+I9rTKRIu
qinRrY+nRrS5HpVjEcH5yMF0QXOFbsKTnrXXo/6jO3mJk6m/R2VBqJ0LzNIAHxcF
VAMES9+ufEsJktPDsvFEUSqfBIRsK5ewZ1d0zL6sRK+jKMOpe6E5PRjXUEJE5UEa
oRI14v3IjdU1mCXH756CJA7LkMmDl9jeD6zFuWiQ4jPtzL+tNqYQDasgeQegcFlt
5C5iV4JRECXwb0xaouCQTzoKE1FK5CHS4LYw133Ej+wLO+Ezlnj2WVbcpR1Ne7ve
rL2C8E9w8vTj2ISO10kUSp5rtECCXsoblUOtjpCRx1zGplK1ZAni04vIyyMn25pg
hicku1J5vxgHUEjDyj4dacM66eGYWP+OjmQHFas87TMawbBpwCqV1BVj1gYlnHVW
TAe4S7nFfHDPUD4P9ChFGio1frU9SKbNc4d7n1vcntbcaA8AKgdqnoVA6QU1vePD
Xr2pWylR9QDNTzTd4yHDJEyc+rkzT4NjGil/jwpcptWWmvIn/3F6ydIwLDX/hgyE
qpepHEAW0CXcaTYRzFV45y2lFjskoSN9xE4G72P+8p9Jefux/JZDIhr1+JZXOM46
fTm1PX57Iham+cPIjzMMmFlXnjnx0N6u2BHn7ZsMnnUpPU/PzocqgIMZZlAjQfmY
YxRKR4/0ty7GKrCxRjy33tmb4F7DQD68ws6u9n5YZSBIbKnDU6uIxI9QHhVoSFZO
hUjyQVvjlnE9AsWjhPB4Bwf4yZHrinrx0LbicWcwVa96scZ+e9FlFrf1THbpSGAV
hvCW0+mrO/c7eIBuu//spU2vR7HRxzIJY74qt1KBH+vGU56xujJ/rSNzg4GWWmJA
4R2ZuhfUqHl+j3idSXVlTGzlNiXdHtWK8OlTv0mk7vj1bvizeBYkYuIr1HiAzol4
6QklAMshAdo/9Lugp40wo4I5uhA3nOXZJXVdSMq7BiVbqP4k5tOa2SqYynbxk8lC
kNetlSBwFP8CH4t6bZgbiof7UoOvxsMvcuPoYMfRpfRtevhae3+LxDcYzobLoWGr
gjxHguQU/ibIQFhwEJiq0MBslmlQ+ATRxeLtMU0zUeFuDsdP+AAqOOzfGWCY4H7i
FeCFkZVdnTb75PQ/8FhdFQe7Yzleswhgwqi1RKunFBNB8OYdl6NiiMlyIav8Bs+o
9nm8jxYznamYWSNtffJ/qElO7Y5qJZPOKiAiqRncsUc2Wi2LIspAjqmRQBaTrZAX
jLRf+rZm114MlMRsYhy5/5Cqj2ER9fFMRSC7VUfu2NuYz4CDexRdYzZic7yzr8wY
eldC4yR8sy+td0TmT88++JOEvgIh80tuOyccioXll8/vRmpvfRc4VygwX4JcobTd
i9ROar95vrOZ7ecwAV9KGl8daAXBtPqmF+v69gWIWOwE2QqJ5y63FelLa+BVcoey
J+smlvWyhL9OkWOyBYo0/YCW3Ap2ESKJhAHUo2OfeSCmeZ304qSHQGdG9LVRSWRl
OLV/CTSq5qsFTUcnNvrwtLhmhahNEQCpe4V5IATlfgXckrGRiRzSu895/V35D442
CVZbkcSM4QGd9koZbvdhfBT7GkHVSMIXN/GvZibKewdpblqc2hmlTYXHfrQRG2So
chb9Kx87XeOXmsSmH6eK2PCqF8jTBn8LJP7U7mLuYD2862iz9Pvph3oPUCHxq+kA
qOSO4GG8uMpWIC59OqHm59lw8w7SK77kaEqD2aQI97V7vdftgptQrNiAyxmktTzi
OR+ChqNudy6ivCijOt3aIBVm7ETb2p23pHcpOxhG1MZzNUn5o8r9V9t7fdomdowK
hQ+vCP1j/fXrCONnes+y0Vyflmkv1p2o3QTMOVC4zhTgS1ncpDmSTcPikyaFO1Q4
LWopw0Mqag02hBBtL8YeAyZj1OBCHsDmc9mvxx90Ruo9C55XTlXaz7jop1I4x1eK
z+hIbjTiQmkRpoGpAa99wQ+obzGg8iFakJsW4wD8OYdZVEx41wOuOwbYzYXh+Te0
Zi+PZ/C+i5wwOqxUUhj79nmchhjXG9LlApI5NcjFbAH2sMSkYhPN79PgNYNLNRd7
9tDiCN4PGLxdPfXQHgvfynEIs7qtmkp9z75XHGmdHtvxme8fJFXHhCpsu75RR7TA
tlUt9hkPn81okeQuxGK39lSAAbagAE/ya9X3w597tiDcgiocCNA+RNHwdE5wCCHc
/HNbeU99ipfCbZfOZtUqz6GOU5mbY32nxVt4piRLxn34fFqDVnbfxLzRAuIJaPB2
iOCbFQg1MNZU8FnjLKvjCp0NGELpgH8FDf8xflEsL6A77CV+S2m0+T33+6OvLB1w
KEfyyRETLOlWB+6I667whaLOI27Ik59FGbcgY8rKGzxkHQkj8175lWR+iYy9DoS2
J18ZldQNqgyh5bAxJ2ZViIlY4vjd5B1ha+LfrBhjQWiqg92RPj/cQDjEBOdHX3Gt
KJDMDX6HBCzR9jO6YeKDSXegifTmA73+FdDcfDKVW0gkwHGY9C2AEim1w5GfVjds
m/uL84N6qtOvH8yk5CUhU2rfYwGKQXcEKf1IcDcbx8DKzkoiYDBTSfhpB7BFMat2
J6TVy2BlqhQ4zWn4sqNEKt++HDJIXd/7B8/L9zOSwHRD6w+BokhD3mNpQG/S+B3P
mgrgdAlrUHYe/kY0HhN+GBENyR/bJbUiks7H+X3DE3essHDUyv9rG+dhcGJ9KgzR
ZPwGNeDzKx72CeujoY4HQll63B1dArPGN3ig0ICmxCdVGPTuPM4qt0QYKBPYdUwS
W2+Sv8c2n5B7s3wFIxa9+lKjqLn5sWTupl0K2Bcp4rV2eLRcgN/RNIHOccNrn05H
BqyOsNE7h0u8pfv3B6cWCEc3tvH+60bQbUmKmQk7iCRsJmPGR2x78r1bI07+XEXY
y6j/UGKM5VefAa/2hPnzcAII+awAOrqerPmklGu+Y1XyC0pABi4/EaqdrYzYNDeh
kxKViIReJHUJURQ3zPesjiAgf9bhozFZWM4bPRTC5kDkEpiw3s4f4GCdmJUsdX2x
/vv/UvU7bHpIcm0Jnbd3H+FZE/LWfaODycAkpgC2OgP4XGvOBf7fN7A+AK3B95nm
cINv3sMvfELwe9ZwcKnu1J3XDBC79BiPwywupbMQo04Kgqajh6geh9XKog2z4h+m
YhElBz/9GMv1fp7EZi0GDggitWX7T44O1dOaOPEbKXJnUcqP7xf6crsEsW8DzKKA
7LwEPmGlcBVijE4GhSSVtrvf9g1zS57U3QnNS8gISaTIMoN0Yvv10Tkr+jLArXiF
rPFA40E2JJnmVxVPOEGcDaKJaQPOVSs7MQmuZK3d3dNLGUUKpp5jFODtdUAhV8rq
/VX9mGSXb/CCPAX1U7XzRJ8ngFPXT0RKu6Ck0IZ6+ETdjOrWRiTl6Gqx96TQ3mV9
8hY2P/yjAB4NB0yyEf5qUIzCpGE5B85i9vKcPyVNsqHf+hCAUjtiRA8v05VxHsyr
6V9ZthsJOd3lFZtqwB8f5sfSTumxCEtyJyCxhGYcihrV6CcKvK78pHBwcKHMAkrE
fzX34VfZJ64wlC0ENFAWt9F/l6TyqltzdPUUFc/h7M4eIhTDHKeB3elvrWCzolGL
lieqnZ6XuGP0X1lci0TIB1xLomOcu8jTitMAwD1J6YqSpj+i9Mqw1NLlHJ2fbucP
zNCXnVaz/vHX/f2yxnrckycAOZxqjUt4Y/uwYbFLm5hV62Xy6RDSYsNYWj/pBeKb
EqejR3ijAkeRPjrdACgV4po97sdaLfs/U80R5BbZtwx4opr8IGGIjwdl89wNPe28
I//SR1m8F9EzVlUSQLFGeTGVTDFW5t+Dqa2ckNv9e2f419di8FSE70BwGzwniKwP
1eHaDarM5NkAdbzoQK+S8G9Xjy6MNst4k3BfuHpeB6TriiOmTIKPowQvJiJrLXLz
EM3sHVHF+J5sFXbCdU36sZflFDTGB0eOpBkne1MotPSWC1QlRNoM587IhITwo5T5
iS0oWIOOx/6yYTMNr9RYmJT57JJtvqGU7wfpG+WOHgcyvzKoJk5qJTKQBQOBNjyU
1llu4Y7JwisGDum14yma6dhDv5w978MG9rdaVCQSBVlEC+eI8AcQ9L+8c4yTg14i
HAK7wiLB56f+b/feayUq7KkRQ3UaP/s4aJBwYZOW5dhO4pRujF3hlqr1d8KothLh
wmQ7jZuHYqJilCWcUq/m6UoK5IpGZ+RmwOnsACqMupi0o1w1WEvdbHuvrMd8z+UY
cliyy5MZrZBractjNQAZa2kPIgTUWEJnVSKJMnf8JZCVuvbTZrLFr+wBzL3DYju3
HBLbEutnCGf1+H27KaC6MJjqNpumn8qoJJU49WegPonj4IZMUD9qrL1Y4SdRAEYY
TMGW4N484B1CHKYIh62suietlcSgBrzO1x6m/kdPdmFI/aH+NnWK11ruwOaxzTnA
ObOProF3KmfqkZetTfW6722BHHAw4Jo7clm0c32bXB2AsFFnaRnmnyh8rFiL6Jj+
DuNDQHkboG4hwX+ieiuDbQNLr5pk7RIkF4R2e9HqvXjwVMtL5rr/UpluOpHCKFs+
o2SDKtQ2VvWLQriEttZhMEW27tP8jsCjmVnbe5CB361K4kXLxpclxp/vaurhgWCe
L8v7p1YvImY6gUPB7HFr9spJbosEYF/ye4kMERL9iBcl4p7FNvmRW95lS6lbWrdG
iCrcI7VH0RE1zb5zy0Nw/W1ENoM/tQQ+Da7YpKlfEe6bDKBk7Z+l3yBcp6Te2IZL
qrVexBbhY/7lsFJI5sUfHKy+XNJj0y4GkpmK5iZle/Ocw0kWkVx70Rm1bTBkJ6M5
bKZdc0ubPBcv2lRGLLvipKY7JtyLG5BC6T3x0d8O5OtTVRGb5/WXs692Mjjmch8t
Z9DlT4DV7ToyY8cWVRKsm9rSUZ+X4N5OomrzQAQOOfCBpSow7Msqhp33LfKs+8NQ
IpPmP4W37P1cO9aGG7Fi1bwBEs+9xYEd0f0LaPbJbkUVabCagON1CQbe5tpAdJzD
`pragma protect end_protected
