// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
ImIDj9S3PqsZmdRPCJjqvYv7WedEmC+BzT0RTtSXITK2bySM3lxToOWA4oWk3i8T4Rpj6iCCgbto
X2hi6nuVqZYyJShXdrBKnPOeJ8wEQ/MHXQC9Ut5liu1O13Gw8Vr0RkIma3+zNR5rg2SUQdfkXvRp
z1/JxXMy3UMF4aeNM/CQC6go8EWwk3H1u48MnQSBX3hgxNEkLrEv8eXAEpr0ge57OqedV71SuSPm
AocqNYJKXDkEmwV18h7nbfXNLLChS/VQdSZnIYcTJugwh4i+9K4KQM5hqhBK6UZtY330WqpzGudx
WvMktIlG9/xZ4Pjdmqotr18B+qMFR68OK/SNiA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
8mKnQTSGGhOvji/H51T3tLhHn++7gkGxhWD7bpRjdfiefxItww17fjo2DjXTCBSsJBIowu3b9292
yyerEj98JNCcjK/NCxNVXdTZGcBippCUZa6a26BSVA8VbEn959aOTpsFKr/SoCaiudOt0Q3YKIXu
LrBwaoDxqdH/nZeASC1nq1O0NzA/1NqmzEnXne+eFRCLjKW6wA3Hp0/nAHD5iqE24XXeIXZstBd/
SO+pF0fJCdDv9zcbU771bTeF/AJ/GK4I9Pwo/j0TMoJjv/19rXPYnPQtnMiZmxNMBeQvCoMwv1i6
UmPvuaWg9B05Ag2eClFy/UfpH62kmuW5TvlbqBU9cmfj/+YnDgMi8JBKNFPoNaA/XBEkoiB8Tyjl
gnTlW7UrgNJSgWBDf78H/l6+nBp/KhZCZbM8Ws0TKK3ageX9KsQ5qt5oEuJDYFm00grWpnFOZ9G+
1rVEK9EJbrPiEgNwTJYEm1qvuNv6C2h6Qj1wLN4FNMcdXt6pA0VHR9/JLHWRMKQB95DWIvDcxN3x
W+ECFd/XGBXEY+RSynN/o7R9ag/hodzW+gKJ5sU0Aa3TtCmwfXjfGGv5C22DJagYMIxmep+aeeXl
KvhivglhedCh2tRbx8Bv5J4+NvdIkdeNhpdqQ7mYxm6mnOAnCC58p3T3GUHzgKIbbRvZ08t2rY5V
F4nG/K+who4mUnpUQcoL+kUoSlWo8+eKnjgK4hb606Sd7qdLPlNu+HxfeDV93esFCxp3ZSZ/BbaB
J4Ywhp6u7t9axmcVsFWTxrdVyG/38NJf7hpGpyK+xoqvDn5EtxdTBdcfZh8PgbNJEiAi0DTOFgvj
2AdJe5lUsg8lL3XV3fub1R4GwY5kYToEkmQ3Kq5FXOl8CIVQEMXBZNVcrmIeQ92YwyjqE4tDE8UG
hom1UIFuBaqz09GpV3CQFofImnKEYNl9v0gsW0dWMeFHGtOg+IJ06yqOGXCo5OvpjqqrMq5oJFDT
qH+DSSCLJ1bLPl2q5pqA32isALKdWtR82TaUSa1Uv50sKlsL/yeTRLL7oKgjvuwjMAE4eiQLKkDr
5VbeY4+XxbwKvzMwTkrLxCdU/Y7a2LexYiJ4JkL2ic7avyFBf7DjfSWjoHUxNXXhk0Rdi6o3JAtU
R3DcjG+vjtCz4t0KA+BJPufDNDurKk6ZVtphNO3Rgkmxbq4EnlSkt9zw2WejHRwXe5bD1cicH5u1
ji9+kDJuzyvzeatLFaFcxmHYqZ953Ha9OPsvKQJ71yq9DHrIH+QuyAjHOIFV1SAFEKFaSY0xg+u7
olWPDnjB40y7i02OJEKLCpp4J9QK0H12JERADWZwV7udQcdfmmYduRtVX7hfAxWqtgZyEaoMRf/M
xgsXIO/3/qJfsvOe6qP6RiFoBBuuVsf3ob9L/82KK8cvApMTCVTjyQqGyVajx/9oukOID9Cm1e5E
KHPmv00uuq9M+ae958w7q45ua0l7ZAcwXAQ/Qfg111eOx2E90dt9+PURa4UAc5ldFo6JZH7XYWPm
rfMYFT+2uENo7PZcv7E3hUaOovp3qyPeW+tfAnRf2gY+4yMINBEyDaQke7G09ZGgOuWc6/RB4LdR
fT+9nTy1Eql8FQ+TzASkNigXDyJUWl1S2yWGM/dYELo4ubpMSwEdkJZAIQm06nolQwSMI+P1gFjV
rTr3h+ypmyq/IEI1SbWr9n/hKFZAbreJUJQc3/84xdjFHSWBs+tuwilTd+4KBM5QWqeRes1UOoG+
zE/qrH/CrXO0c3ibAl+t5A4sGGjmaMJ2aHvjdVtbll53DVhO3iDTR+SwtHrTm4TGXwVFo0+Rda1L
4eS+2FaauQB5WzpjrJFzKz9lkZ1URBqlHIJzuBgu1J/nFlUfeLvOnVA/PNN4eW9MJCVTA2cyYRZX
wNAQDmnLsWF4SAlX/lX7Sv6LwEhwLsLNskk5ParykoYc4sbwFgZLrl0N81uBULJTC09Bd+z6Dm5L
GM3aB+N4m/x+z5JbWxAsH20mk+r+2I9DildeRNomOv5Dv4BSgUlHUm6WtPePTwDR4UMfq8nw41hu
mxzlt1e6ZhX7sc0Zp+Iy0hzR6YOdLubHPiJT2S9IUW+yI6lwmTSCgcGrEwD+TiPxmhOJspvWulCf
N/5CCWPp3ZbjPM3DVfuGyfkFWGA99Qf9+KjjKChdegJOuOzjA2opsP217hNPUX1C6sQHhOXRNYzm
10Ki5to9e8VHAO23A/vLz06wk4gM1Mi9MFjAxXZOOTz0c7C3yLSIda+vjEbHuYhRFWYrNVKMV5KA
3+ZREScRopYVJCTnJaj0XuiQFsV4rXuQAiOJMZUxSzHePZrVmgaGxCHi+0e3870PwTGB+1+hkojf
g0u2mz5vJHyglGiePoeg0XpPfb8cLK2ZSnluORaeW6MicASCwIGtr1cyI7U65eSFmoHAYiOlxChF
CAKBNDJhOlIdvYWCiNo69Z9MzJceProDd8ayHpFv4qwXcXjXwmzQOdQwv0KWixj7XCwqfRdz5kKh
g3z0t6ZdOHPDUdUnb87C0VrJSpE8gLW8+vOMOtJP37Bd97R9A8HHlvI1MMTztNCE091PMj7D10jq
X1ob4T9q1MWbheHekJlZVr+M61szG3/uUSUBa05yLfGZ86g3jJUkqn4adsosNMgwuYiBaRxzbXmr
mLiK03+gECPIum+sUwTAylqFlyVJPF/VOHHkIjju9WjrYGvwdXGa+LYa4DT4WKaz8agmXe4TEFWy
N0pVeCzHY86xsMa/Dx17+Z2SSWRUZkZeqn0HnpRghHTToRJtfQP7elpasvCDc/6bCTwIsJ9rGOLC
uqB8i3ASqnPxwPm3l6Y8nX7VJXZ0GUAUUEhJKZpEFr1Oa+75vJMWkF5eBGCB3bA7LFQ+PT+6bpfd
4AGATh8q5X74D7PKRpbotR2IfwnloMf94bzeDedSKUbe1VaY/IxczCg/aKztyAdgANZ2pWO4OWmR
p+9DwtwSba3zzVRla9OKCfDAExwpf6MW+AyBz9zfmOpOKTGtS1P4LaM2f5F2BHFTQsUlg0DeBnMu
YDSN/IXlJrvbu1yyIJPIsZq/E3H0mj9vQZsD0c1HIR+h9ubaZ8v2aA2h2k+5mp6k0AqlfMfiLrl1
K+dVaeERWK6j33Jc/tQCJKau/DN1bl48RwyRsmZCn6ykZmQPEdAC4vKBCxg2G/aq/pCY1KVR2kio
+H2VTE7J+Kuq+YNODabbgXn9W2YUNPjSmJG1CmeLpns3w9qAJ2bVAjBIwdib924dJjcPreQZCGg0
GgcKTPBwRId36hWe3XdeiW5FMUIuYbbWh9xEvish52m9y9kbuz54e9EsxM2XZTZI04JECYSpSKxn
qGkc0j4Bp9OS1xIMGuR7daFyMVev1PrXze4hz9RMP2iXCrqPp8LXFi/D/yMqSnJIaOiFiwYs5+bz
YYwu9tqX0Vk9t/5E6TSgXLervMzJX4gaCOe7q6rlNnHM7POX1cvoZO91syDueeeNqEB8MUoRvqZr
osY/Tu0fuEzmFF4mHDwaonUjKBGhfViZ9iPbJuXWL7CIrDnLH5TCL6xxBGWC2NzOGwy6dTEUlAOO
llg06YL1MJuR/Y+D4Y3gEW38Mbuh0JzT+fwO2jonrmZQj8j48Qo2NjR9CzKJypW2YaLMPguiL2gj
zGSTedOY3dnZd68HTRprugac4rtVI0hit3+mw2hiWrr/JSm2AArClJ8XBDaWrkH3D7I6ydIRTbPA
dVkjzFbvue/pwAVz+MADB/JKe0wIe7MTeeJi6IIgfdgKuZ4MW7w3z64trHU29DYWcW34VlbA9Szb
POqI0LUVDrm+F4l4rZ5zgULHtfSilciFMx6C0joFHiwI9NFsu70g8zQcNNXxMPXtGylFLGWBwHAN
IDE/qb3c5e8m7w7QWlBXNSCUbxQJulGxhQsFvi/LvD+SGZk+v2knNdCKaB9Jud/Smbq5EPUv5RYG
AAQnP4t4qI/YeMduAxdcwC3kzLvRj6onJxMJVAFSuxa6rsAxAT1Kd4po6EtvSL3ZKn/gxvAH40Yq
Oj47nUV7tlateeHgKD7Mx99GPZ4SI+bdeCznaTV/cVoAR6/to6fuVNeTL0soWHJTfwbPlH1/1bvV
t7iXJzhMFZWjn+tv4UV9SgggAT4+i5wdTBBn+2/fL0FaI9qwXhvLXHyouM/ZPacRPtLladzi7u8I
0GyPWbDhuHA70MErxd+KuuuPCyIh73x2tDDU+gKYRHDq6f+m7FfRq2cYGdMRiq8WFVfD/554rbdM
lMN2ldh4kKx9H0N0+fdf507a3BRn4GZCF1BQ8lcIo6vm/BNxTfiAvqJci3doiI/bJ8cqIGxm46jF
ao13SY+OxTxogxqd+k8B1EGtuOxidod377jycEj+rCvDPxatAP5a39+FqLgiWzSvDqDIAogTTcpW
4MkhBCo/vpbF0BAsXVlT4RkNKVHxQvxOo7DgsfG4Dq1S9er9Glvemwfn88CnbNrWivbYaEF8WdTm
m6wIMuHlMjj6e4UdSZClCV2vkNgiZuj1eT1isTift85oCa4UumCbYzJ5XdtwR+EqF9Yw9nCcKL9Y
OxoqpWEd+jRAs6up4aZ0I/g7qdQQDaLE6QuMSukM5WPVmWtiqfcMJW4InL7YdadkFzLoeszMVz0X
Q9BwbDZtCW6UNdM5x9v/SebhVFmmS6G0bQ18F6B0al1zPeJSxLH0fIHh6s1KHjLCqFjy4dqrtSnJ
y6Xp0AFfyoXXdXEZrn22NUL7dECpHOJfJ5N+s91eOSFhnfHq9CZewFBEtvewhgNbIOscEJpVOhty
2aPVSAF0hQ3V8b4JeshnuRv5i64X4soaPlW7XGEXeUFgtXf0SXXE7QFAh/fCi02QezuyjaywsidO
VBCcOnEbzMhwKzC5VCytndOdKmq5NlbDkOYHp0bkREJ3iN1Jlug9t1aDC0jOaf6ARSgShCpFVPd7
WKeMVWA6M84NMx5r4uHAhwdcxWBdApYZ05wiGrOOhcDcwTxODfLmx8lRFtvf/LvyRM+iXAk8Dl3C
yPnoxZynctwTsZfZwN02v4KQpAE3h/6EWjyJj7LjBjPIyvfhBmPfTbWenueJxMjtXyP6avpYysqQ
LcdfLyOVs7n0NpOuca16g1h+GeNv3R7DaTvPb214YI0WM+KG/+04Yjew+3y5Fm6/kxFcQcBfz3RN
KOMOaWzCTvtukAaWbT8HOksA6GlTtS5ONIW0nDr/U0y908m6AK8ODqZ/jvmkyPpgvVo72GvkSJeA
Ye5crmV9h/XJ93ymD2p8/ApoPuCFp1WDrwWeUrB+er6IQ1n6QoNZQJCCCgCrGFitKzTfTkeiIPBQ
zUslUaEl0AK9fVntqBum8uvDHFobnFZ/A2217vhKsKqcNbgov//mClVRfyooVUZGiYWiJjT+mBFU
kU9ApJZ1qkt/HFge6CF5N1Kk0wXBqov0a4oUDA5esizxJqQy14PskkWi4r7rN+4Ts14xAHn21sds
XslW6qA8aTiKfK56dOdgqsHdl91vRBgd4yLYgj8KsQAirU2CwYDwTcIPhWRe4rYxJFb0Fyrmws3l
p6FuqO1C+zkbwlkboFz5JuFIkg9jQLKZFl5CTQDo4V0k62Xg/iUY6r/cBv4KKeLIuwyNkrN9BhSd
l6lprSpyD298/l4PIjZvmAK2hqd9T4BUyWVKUtc5nz3JIeXnuJqIZkYjuc8qrMAhzNvhZX/kfMpG
3TZfKHXUbU4kvBZSoE/8azxWsLByhoK36sLKGF7P9VvCdqZi3AI0FddF5Xab5fM8WYwMOHGUK8bW
pFSHoMf9p8LRbhWbOJAkWrMIB+JiP97pBCCZF8MHWvEnj6lxiL9RjpORzv2VpkiQ86Y6k6qtqi82
JoXbnZAH6QlJz8CjpI77U0riDFG0r2SQbJ2FsBAjivonNXYnbneSow38FXsaAB9cO0qYSMfUgaG3
UuEiFL2uAI4Mq4rlKDamd7HEEYMZDVGfrTxNe+mYDUa2aN9Mnx+C3Evq7WwKmXpfUcE0GymqHq9O
60+DRrCBwSZoTDffGnjM6L/UNOYyuxMVWMmK+EwyXMlaW/egD+qwwXCZhjXqRdP9FaGorRRRMuFv
zx1WjFY9BSlbA/jbrNVWI56IePKLRQi6FdRyfAV9hTsL4rO3GHS0G9KogMuRY3oUWYjVrs1z+pk6
W21HTrIdcCPUu3FrHoXyBhocnw8hblHCgYLCsFZx20WMqf3fQen7hl7dQq8wN20BTvCFsmd0rBHU
OaFcI6c1h+NxB8RdcMWTJr9Ntv4w5SatyGhlASCGXqO98P3nmwU5r5b09J23tbPXFQbtoRY4270l
qBN+TNzmtzdxZnWTjSR9fnB/uOuhnF4v8hRdq+exRsOpkDYmBfBOubBFZQrHGcj3Y+6RPePsH5Zb
iz7SLHMhmGEJgYQ7cX8v8uQp0PUWZe5XTRB7tGBPxLfe/PPWKAvxaBWNf3wJvhi32X10X/sa+0jK
m/nriQIWH4qhw6v0Vb+/WRBzzqaQmifrDR3yExs9s3o8k/BaJh0hYuLBMTlRG6BCSpE1upuotmpR
ib5GXK7hj7N5gY0nKqrq8F3ANGg9oxp4aPfErrEloxlM2lCMNiSbCUkOm+ALBCdT201NcHDoJGc5
CuSWYAEd2bR+wzE9VNeLq5z7BrUKYduwij+qtX69PU4pI4/0jKAfRGZXD1jiHngGhjnPJ5NCGSEN
CnM0hrxavOinSR7v/VIYEjUtQ0gW6rhSYKaL0jqF5sH6jrn5W/WJjljFcDRgiAaGBgbv25TJupf9
I1Qi2w4m3a5nO20aPhFi/sdYJu/qP7jEoVnrI1ohXXJDQJnhoCPYacmbxrw3aCnJWFETIpv9lkKn
/CPPA4WgdWSmfSHsm83v4+zflWUWAb0VkSBe5jWOKEH1n5rbgC8JoT9zXFVDqG0HEZvBpb++7aRT
iwi8FvwScW0ZCZm4ZxpeYybJ7xpTrRna2Yvoxm6hjAH8MZLdagMtv3Ym79VKdG8veLBXcoK+pLbN
x6s1AMEZbfjVExOHXo32SzBlvWXajCtpVSfu05YjByH4To4/T1L0n6kj8dZq+OgrS80ji0gbK5an
sv3nEyMJ0ieRdnkltOjiXgtK/qOKD7qJ4dkkjLiqtLiylViS68Rt/rmavLtjHQIkDGtQfXrhPQA/
9G0yzhygKRaZITwkA51wLiCNRtyZrG9LmANBk6kQGgu718qLSh3Q0NbDsaeHZf6JixosulkBm6UY
39FrHQkq7bMePJ0BPGe25uTdba9b7wQHi48uvL6k2lEl0tG6+cKR7eZQcUzlheyubwNRLEWfRavt
QX2zs4AveO/4A/18q5EYN5X24vvtvV4/JkkN6TEAzrr3DrC25ZwK4lHTIUEI/8Rvvlg2Oh9Mi19X
qmo+PN+w7zEMtvrIJkfvuHNWH2S0y+HYjluZyF6c5UNQPdy4LyCS2q9ZraUVNLEYHFergHl4eBpu
ZS1+UNWy+nqz6Pwwr9sHCTtPmPsrWld1u97bqwGiIJ/P9Uw6tZFCZFiViHYgCN7/jq9Vs4H/DENt
kApOgNKTFzDRXKdqlh8t8vT5XG07gCgo0aNu1pRo3LQlO7o6NNcAYUcpuzbmJGV6/3s1KchAKiSV
PsgQYvZJRfFJl7MMk3qu2dMCuKoGY47iihZwX+2KpEsDhadLYBIVKC/ZWCgwrIuwxaqasGIzh+uA
AoTHYSscmQOtGliOPOV7r04ODTb2LK8aJh9hc6TVjFxoHYklMZ3MgcuLRB6TrOPzxdI29j20Hgfd
1niFyO3xWoyoVWywsdtc2Ar0JUdgn1j87S6a5/cMEkjrcVtrC9xxoHEU64MDFLwekblLdD6Bgi6u
ShpnIxL59eLVJnXuTniFDQ3YIEdeiOQsKLCtMyTE6GlALeha6FFvnnlvpddjRt94lz/2yk7LQSQo
QCIS5A/i+9H7g1chfb09p3llmKI5q+dh8LJ/LbKUuX9KIrOkHI2Ce5jwUsFyqbIx1ddo6mQdWuF7
LnZHKUR/5t2TNSAzP4YpUWlUKP5BNLWrUXmKHXtcn4rzObeza9B/u0cCRP2jsmIPNDvl7lQnfZCu
PR0A7Yj+lxQ/7C0c3uMjXcejTDciwO8eeZ4Q4uVsRDFcOrAMr5ktK1eAmXVTLLnkfU7lVtC9Y/jK
l58M9OetCAfmqvCkbXOE1dmvZZbCxjtaMAEsJyrYjAzpU2RMk+2DP6tscnaRyc/EQj1nHSoPiwLw
0jN5GRaS6UsHsQWjnic8wWCX3dLzVcOtQziXuWRjSOA3IDxSbltdsmQO3z+0iUvFpvm8Wm1vTZIx
s/kSpBk02u2aSaGe+wX2YmRQVGSpcLstPAx/zK21PGDN/F8ggS5Ub7RbjlcOwNbpSTQJwlkC6DQb
JXj2NZHhfv0ip17qCB8jqwlL4TEjvVh8HjGBuG6Ilr6kIFaGFia3wMlEC5k9s/DBp7GX5rNkfPLr
CRGLsGD4N/juaAi1H/TO+jQ2H1WhG3yvekRxHB/A47MlEWBDhCWXY49rB+zrBBKLR47iiv1qweke
tfujlqEh837tpgcj5aMevYJCb8mf1pRG3OlbFVxQBWNrXFGXG6STmjmLuT3vfEuR3aDxkO7Lbwfu
2yKM5wB+uaLejj0TtQgH4D+9c7RwxAP5/9lG46Z6+XF4VBoMyzdvbprxoPkpQQWXmqD1kzokScmf
xiitIWlGQ0Scb6BJnoR9zR9MDgvtJPkfjvNs1BHLPEI7ApF6SstMgm/W4VApvaEveasp4Ex+JIL2
wvK7itxvmPsDtGBagZFqWG2u1xzMqtIYqJ1QU8ZFKLL0+7wofxVUfqo/f6zS9OFJbk0VSQq8SIfs
J6NuaCha7WWOHfZOSRG9gP7EoA+Stx3Ye6ejV800+rA9ADvKrIppwuL4K/n3c6swlDCLDIxtXvMz
uhk8H2j5AhXRQZ0ld+XqLzadH2Mnv/qTT8f0liDK7Cll4bb9w6iFlcOM/4gI0vGGvMmlFHNH600L
LfVg5NDT7Mxi85ll76936Kw7DfY2dQ4c+fgXgDqIQwfdB/HmY+eLLrWYcO67XYiUJVLihwGZg6Nj
u/F6XxmnSTR309Dzl3L5JQpEYAO5e0+ELVHupNOz9GvF2AcCAvGwVXCrX7a0AL2A4WpXD4LUkxcX
5v3n1jZ4MOtniV8SXCJxZ9DcHQwl8vj+iHbTul+vS0t9Rc9hL9K4DajIYKWaPAP6a8nXmg61RMET
E28fsOxWLGGzMBY/CvPM9J6Pyl8xKm2TKDgYhj80u/QTWyRTnkt8KoUPw6+QUMEL0nNC4Y8hmLdI
kMQqjKSJL8VQvfhJAG3mqF9nBsq+ZcFOlEELrqk5wKzU4pK9r86nxJashuP3ygKx6YD0tzWvv2RR
froY8ZLqvaX4H51/f21Td8i7NQBVky+aCSI5puBveaiBeei0+5jLjg4NQpLwqkP6hBDmYbGs3nz/
1IeEH2LJmxx9+p6bVCjVa3+I3O91pquG5i2J+u8jUsSbcpFG8L7dlppZmxD9/T4VqJkbjAjYiDLw
TNRVFk9ROjoWT6zwHq7mhfWzBK8a1jLY92MZbqiaHXdM+6zySC2p92ALKrTHpfg09eotAMfu9unv
JeGzsumEZkEWs1aLxEvBI0BJ88joU/1LEocTb21xtigGHdD6mj5DPyID9qgG5FIM/FxqmBerx8fF
/0LoAXJTOA8du8J8BlYrcr7kLuJz6ex32jaOXxZPw8bAGiW9oD+4Bw9sh/3mwu23hItlNMfo9AE1
Ti7jliBuqg+rlksAyCEytqneWxdMu+z7vuKrfCsL0NkCSfLw2n3KVOWZgn9Sj4HjfLgiv5pD4hhg
PQpovF+qfAZTc23m5vqYJLZnTRPpkzx/+ibiAS2rsa1Yagmf2+FzvLObcapWk8mk0yvYGCSEFAYu
V9ZtudqjKeDC2vGkJKB7+sH4CwvJwRkzVB6BpN6i/NzHrZWVvJ7IEj1ZbkoKhqVE6k35Ozel/gbK
rHBZU0EfmPTBZm45HUQXGa9jjRpwmpElueUeY45/LA15tqbrBLPqabuH92ZozUXwH583+Yb2bsTB
vxdhQg2z1RCX9wOJ1eM53PYBaCgldv3mQSD22X1uSbEvoYSe6hefPca0/nkIeoWYMziuesi0iS7r
u9V0wA8JmszkhUTOvGXlVWPyNH9LgFNOkG3RiDH4QHZwaBfml7rLkF33Wbw/gzVvi9ZDsf+leEkA
YQfcu3JFOFC6//26nm6n9n9J9+lLwjhYSl4EXULETn4XR6KW0snbciIXBo10SitPMW+7pu98cOiM
ObKyccrb0tKWv1TaNg6XZvGZLG2JJGvnbq/SzeTKHpcZOnkE1Q4hqhUhALDGT7bsgpA12lBDlls0
x6oxpRef0aEKwkFUmGwQQ6dzaGEyHym8WnV0fouRNuxSdp3t7yRlPCl7739TwffI5ZMkCHE/dsCA
MMRHjlF5jmn6ZG60s2Skkb82Xo50QUwvEjXkpw4qrprsi//pFF7aTmMl3hDIVzAorna2vhculd4Z
bJOdqOZJXONS87fxniZO4EtXLy5k32Gy6r8azb8cDtbYB7iyiBapPTeuPkeTiJoiQ+6JvoPvvegd
ujX2pXZyNwXczjuDd8yiFLCxTvnEYjulC47RHrzaQsIoUqSXtzNZ3RTTcJz3ckBbTkfxtH0WWNMK
BHo0mNJHH0+WQTVyWEEPkP21SXRJcPOgfE2gJAtms85e7ukW3bdQp++PhddFGc8I+TIFF5z8XhGt
qN/QCeLoreGZC8Gc1C6gAPSrY5sYEUee44Majd3R8GlRCWPwG1EDWipuT1tDozJJ7c4x9dG5PX44
oOfLKZG5fA2Xyij5lbmlfwi2sAVm6yTK6/yRty8yLf2xH7WvMoYENHObmLfK73N/aIhplS29SonR
5OCe956YeHIhE+dZ7d5i3bR7S2/0orbNWpFnp6o+guwtU7Fc8lFGz+KgyMOsC1o/grNDU2/q3lJM
x3s5EddhVApoiEIYBu8jMx/JTZubpLtmz+/C7eRNXXOKrdPTdSn6rMqZb+k13z5h0WYjdYz/RZFJ
3mbSfgUL6DdsgYWzXcXzX1NEnyzur4TSd+3Jmz9p++58zgHorr47xs0NZah5RQAIBWtXk6LHsGYz
snL3HVv9bqASMqVqB8P6lQe7rRoIaPVvVRGhcQ41/Vg9oWoJcA5RvmMnRmvx2wwaijNgl9C4rQEJ
/bSWQPOh4Iu7+4KgXRMmbqj1fwA3N5trmokJWLaqBdRrjMZ9Enzzxbu/Y94K9aR6/gOb/+xAQ11v
GBtasvggmA7+yNbypwjNA4SF7547+BKJILYFAjvJn688VSI3yKFuv0l3rI2M/NVyPjc45zE3ZpQN
uolLfZ87GenY33SODg5U950yEJ692K4jCw0eF5Vjb3OUyjhlSVMTJUjleNnxU3gdUyhf84PhxUTR
7GH/pGnsGu+cvz0YDXMU5W3GVCn99NThg/twz67hDiOYbdnYhVLAMADOhx3ne+0KoRuisS9h7UZL
dmSiIUabvckDysbMyNMKjl9g5UygRhAJF9dq6bbJj1XgRxUa95lY0OJAE5dSvStpGXjoRwLxj4iW
my79F/TbKtRSdQ8G77g273aomqy4lwkYp8PcDxbnFZJXUiX2N2Ljhp+eqAlNm2f9NuAzQF/LmbrP
78fbCoGRLeNopzzvHTnU5z7IIpa+xpCyTSucbXKvwrRcBGVPb9sLgPIdkLyQCvdvyM4AStRk5pAK
yCo6C329DabPRw1EPoZAdkcqxWCaVvveAH4dxKG5Rs4LmSQJpfiL4BCrgqzPzyJI2kqZVxMFvfex
/tpUFpIByNLmqTU8cKANSjpHoWej5jnO/Du51OdS72jTahQidYWM1+evfLcSfAC3pNYzTUcWvS4W
JBILl+jMLtnYvtcXjf6fkX+ajEmiD9UaN0SMLt/PfGUfrAllX/8zlxye1EETCrpOdKlglszixzqm
uqzUcs1oA9zV325Qn754kgL8efUxhlnxIKVp2ZXbOYljNHtxIkU/QYTwQQQ6dF26AjdHnIj5p07c
D6cUvbIKVqWIBSD0cxwXQj2j4jmJ+JcD+eQItsyab843ki5PjN/6poOOBUlgCPB5EzG4N46JVl2q
S9Px+YN6W94vqFnIBl3foawfWFzRi7YUxlySOqRPmKUi2YborB/gNTFf0RJcOja2i9/4T+g5+tN7
jeFUAr7yEsYuL9T8ZdMH/qQ3xN7fxqxdr8rZRB0G8iuQMUnTiDOd8A9ggkzKnW2LGyKyUGjRYNi7
hdI2K1Qa/j5M1XvliWyp0u8WhzJj2NtRs5q72dhfKC9EnAgKFg5g4WKxjnk0rH8dFIr+9LapeJTO
gPY+gmB9w7GUp0bJtGVwfRsUzlsdiygbdTnlQdZwvPfnv1KApGb/c7yT+bPgdMfnWExI96nYEWif
xmg68/+x1COPPqPspr6ukMQE78QsEKpbFinPpx/JCOj3y9jE9QQQnwAFUEQ2WwZ0Ak5AZ2O/psjO
qzuiJvivwJvdx7xy39V31+KtCtzoiRMKPKEt/IsNkjnot2VampP/PR62IvkwrPXaWarWqEiLMBOk
8hkUM17e3Cfmqgv4/TF6rqyGWvviOkO+ZypychaSoTG35tDLRQQ29vmoHQYy740D/x1gE3kHUCYc
iac0Nq16qvVsw68fjEme5/IcU2zT+RRKr9fQGM0EMu3zRz7cHJ8x3gcmmJXHMwkdmsOoCfYYsuA0
fB+Mab51vbaTFVwyenvuSJf+I6ksZvv6P/9MnLmieawYt4f9zM4LmZub4ElBoCySc06NV+DqOV/f
E3K+kcKJtrPp2OYlbIprZU1l7/x6Nuqm66eJ/kKPZkIBEuVVDFm8s1dXKZG3ayncY/FgNGfoSxEc
1gVKX3ktc8tCRYKoVVAUNLHG5PyEqVAWg4mYsoiJCOZfyHoah2JVnHcp93bz/N0zhOFnNnY9ZlEH
Ie5CO1sHF1cR7a+Jaw6uG7SqjnBFyMeZPwErH/rQyMg2ZywTn5COZoU4Fe84YkHsncEAUNxjn+mA
l5p+AH2xlNOR3/2vWJCIa6bOBGrpkfN4GPwgFNMi1oYicgisrEYiT5RBFJwjxTIU8Wog6SLnZ3Ta
sVrFzMAk8W7KbbmFiCcAUziWBxE6ITZdpTZQ40jLWYi2H4I9zszi/vmjDLFwQk2t6DkPPMnHmWiz
g9zlYVjApyjEHhfh9IXvIPjBZONGSaMg2Z9BiTfE9LMGkWs78QIX64S8e8ELU1yyLZg/t6nJi4nM
yUrqXPofdYTYohuaggvAsQxrWub7Co7vj5cGkdbIrbkbZ/Ze4Ho34pv6rEe4Kva6xp6g/iq6O49E
iEZlrJHUq4Pv0Ei+VSZ/Y9lxCJADgww1kwnVpsKA/Z55Bl8U12IU9ZjeUgj1Jp6VMTZGuBY4Ct6b
9PwqD3b8p7fn5Gs2Yz0n2oy57HfpFVNn5FcHsBRgpgxLXdK2yYaxPt4fC1tw20t0sc19fsHoVDfu
g8/VI2VDpvU/Cx2qkHRobL1fXh4EvW4C+xXr2Fd/aFQxYbSMVoHIs8p8726Vp0Qi/LiLsELZ3HL6
osLJcy7ZwP5DX8h9ZH6IRYwuA5MUqp57XchtWwxJKk+Zn+qgduS3oWYpywbvS5EmjC7x/lIK9xco
2CrynroBZ615IQScGvTc9K4TVh5w3S2If/gPC4/dA/fxrORlxuYDQE0d16gPFACPjYccDALjtX6A
eMvKVbNgK4uU2myq6+uyvNbZ5Zi3fcqKCyiemUL1WmOXAZ0qyCx4cDnM7S8apSAo0/Cpd/KvlEIQ
VpSReSMXdvPr+vLL5KzJg20AzLYbPaIl4pGsmxshKqQas8WmulIqZZ04kRREfqeN4XiXOJovXZ+O
Vsz/ma8UV4MhmUhajcW1Iq0Puc6uEJ+tEtcy4BBPr4LrfbSZdG4d5b3JX/KZRMtpP8pO4XqnN6h5
AOxcq+LFl5D8xGKv3jIILkqJdvn9DppkR964MexDRg3r8U8FECh4859ftTb5/w1Hc2eDm9CX1yJl
OaBK3vsP8XFpbaEPuiW1n9Fsh6yQoZjqbJMVP2HhnbAS56csibXZxZ32KiqcjkB9EHU4bFPXUirG
QvBnb+sOHHI+jrgz5QOkE2LzcZGQOFEVEqMOSZGMuSpmIwrcVRUCpfHKVXfSHdSWq4nDWHA1jiwi
dgky6OILw2lWbwyNsro0YunY1Zr+fzGfhnGEYfFFT302UTzOXuYo8pX6JrGWs0Z3UC8Tu/silqYN
oD8eybDFEIplJjWiUEVaA3AyvYXWuSXMFxgl7w1Sm8tfLrWpcNG8iazOrheq6T1OF1JJrbKgLY0E
jBJwlxuqDMX+2h+pkWFll/fT+tw5N5E+MheQQXu6l3gJ1Rfyi3yKlzmuI+OJzQrC/b0xLOlCpXaU
ykwJCFDdGfjdfzfjBeWT2yxQIgccwPKAEsjkxsHCZLWaEoM2h0NqTGsMJF1kcl2uRCvp3OrG6OSb
oSAYDMAFkZRPeKIg//pSk0R2ROYTmhiNLiruvEYCJiNzJh6UTVAb7MTLTaZd31zpjEBxf/2cbSpm
tacEFkYHTwtRfgacxpIwx8emlT4WR5GceDYSrZKs6WUImlm55MJw/eNKIvOI99Hx8oWP6cyDu4sN
DSS/4FJcXnYs08/itHg3e4ZKkzghQYupmZ9MhpDv//XA6bOLuWdjhcSXFSClb1ODizd8NN/mwHi6
o7bgTncR1OMeRDuH9gDjIkCgQp3DAplxlao/prFq8vDcNgNfvtLEYH4hdaG6WgrhMl2zsRUgFSOe
sglp2l+UTGZhE2nuF0+kzbOCFyVNGcPFesoc7wJvvHYL6mghv1aOkQMBzd18VETIMF0FSczFj5PL
Zg68iTNsMlP674VF9CZOn3mprlzX20N1/CEUPXsQIfVgZ3wYcM8fJJTCq88AERcClTuKhtrQjiHY
Z335/sRS+We1+kUzzr/k5dkm82bKF4fLIXOdyalpEJdHh3TLqZNPmTwm7Ai+LcAlSajh2713IbsW
pegPLTdLMQMDmpWsnEffYJtNN13JrBcvXypI60M2LJNMToNWGWqoP0dzbYYKMAyAIgsZzLgmoo/0
tiTwF9MYAmSJQYs255cFeBWOq6nT1FwnbhZg6r74tXF679BlXkUC5jpwkUfS7hWUBNvgU7TQyaO2
aPBUXpHrfVeF7lHMqjoaq0OYzWDKdh3qgfO9yMbKOHDPjnRXD9Ir+t6ve1mwwJD3Uil6fP8eTcWX
uA0rZXck7RVjHw78ozDOT09KiZOMrw/tIlT47p+zlZfUedNrPX20NRkTuxkaNPb/JgvUNNxT/vOi
03oMUGMrbI0h1/0rhYMt0d+YWucjpXE0iqqdGbjovg77R4JjwEjCGdjxQI95ADK4x+6Nb58Kzi7C
icrCHRGRvEu5yPwllfsjUUgVpLGmoH+kujdmKH5UtV42atUws1FGh+72j0bVsw6dvZxqZTkt1SS5
9HmWGZOF7E8bIB/+fVbZ04+dey5Fpje+8AUkRX+SzBDk/EWkerHwqDxSwBreD3/XUuBmsY8t7LeM
xb+3czCr+0+pKNyioLAv5ysivGWyDlT0vyrxtjCbY+VPyuOkFqWx4jgoqGwddent1BgMh+dbqg6u
ydsJ5Olc8hVuNSsJCc3ttlkLEYI0CxjAW6t15PVAHUnmg5gB2STGMIdpuxe5WfXSaI5X1R+EHXDP
T+cNLWu2ye67xO9axajxlDHwxq2hHXKGKkpKkqTvvV/h0LgoeSGrZmtGpyUkvy/qY0QJB/AV2A7Z
KndNonPmgYYT+5ScymPjXuTfLwfkDiWRS2T+NmuNaq9gdAyGRMsMJLU6XghNtdAH8VJbZrrHjEeE
A68STs5ZvphrbR4VpPBlBsAL3OwRMCwdxpnQldF/CE3DVSE7W48t6m54I8bLgBXOGNb3vaVyB5bM
FOEmMrOuyxpkrtr2+nbuL5iCTiRWfvSr3q5aAlnptQjsPYkhUPhnT3Q8GvqQQAi7lL3e8Pxovi+y
q7qMu80KMGaUp7Gcv4HI0shpN/Z3PrN361I0sH0AEQrIj2Cmebu0wdmhWRFQ+C3aCwso0GxqAqHF
lXKQTpnMCoG9ZE7qCPp08AlgaYsOOksqhnmugb9/qogOmlIzs8/0qsCHmZLhXX/NsIHWVAKb3oFu
l0ObF9Gv1Dvj3AqZCxP0fyYvJoFWes/FiuiolRsY6UprIvvY8PIwihohSlwykrbDt8FkhoLrOkU2
fZgUn6DV09se5cMJKrr939RXTjmLPA8ze2n8AUTB7hnDBz9A9YLNHHqgSjdsbZ8thaWykpBzbrkY
7puN/Pz9saUtC1lj9TnRrj2CpSNyfUas9EphO9vf2t1AyE0ED7xGUQXafsVY80Lj9GNkk6Sg/g4N
C7zWj7xP4yBJb1l7ZIHFDYLzx3ywhc1ABJb4vrZdtek5j9vh79JtqgdlXf/IYzIlZUZo+xIs53T+
oBQAwwP6Qp7iTmwlvA4iy0AD/OvXNgQ5Sy0bDaHzmh6CGYa16HkgTBxhCzryP42D0ZUjm0dyP5+W
2IrFdwgvlH75M5a0wN+2H8GvBqfzY3dJEUUt6eoIhsLwN3KqebF5JIGG+swSiqSEWuxkKbsDNFXb
dvaRsH2jtL0tWVgGSCP6va19mrH12JK1p3l5igHkr1Ex/rBOViIwmzUn7LF7UUJdUmL9tPn1aX/K
V6qb8f0MWdkdSrdhPf3eDOOo/uVw7B4zGixRbX5fkoh1bgT0RnKfihhpiA6dEvlH6aQE7VpWpk7Y
BCT1V3FB0tLCCt3/jJmKapwdsEsedRhVd0oALnLSqz7ryE9aocdn/SwUWIwhy2ZoQEw9VZmGE1ss
KpaKzKlSL7VprrPOrGLGEvLCdcKkusjveNhWnQb/CFcVCYt+n7plfjs1kjGhb+G1VPhw8/dPt6df
tBgEUrPK1eKk4eEqlv0oZ9QW6QJeUfw/LLec4+Vqf26a87ZE40aHxIu3uzlgBdeJYuNj2lzxkKHj
LTJ34QD5qFv5VtntX4/s5bLuX+4PMX4ViQEF6O9orEaf8Tta5mU0ljeYGP9nb9StpI3D7+YH+jt4
e2mvll77otwPCkGWJWoViExSmKGUe1R+U+1B+MzzILbiY8rjSOqsA5CV0o97P29PZu33LZblRnkp
JfGnF5aQmC3cxTu/h7CAjhOeEmRDcS0gi35VvPPZnOEavaDWPHUMHyO+wI1JjSM4umqp06wCkTzH
tp/ywso9HIKUhl2oTcsN1R3lbl2N3DDbFEpDfGAVbPRvoOtmNZZoosuPKwM3OiHuoSso0sdtsS3t
CP9ZL9+IXiQ8qjbxwCI24OZgnE9+qDId4VxMBFbiR4UpVuxZEyqF+BDXs7OkPiNHJS7gwAcTlW1V
uQEQf8qXZcazaU6qE1L7ifqs8JS/bZVISigQuFDJGm/l9Ah7r/AcXtdrKK9xX6guZDgQJ9C2Gqa5
XDBFTCjURWk8a1Uh9+l/uKoKQVQlPbl4LTMLj7dbTgM8eOjrufeI+V5GeRtQYRwitl8/8/l8d5vi
ymx5cJm8ouyyV1XYG3y234gN3WbpHxRJO2w0T1ydqVYAKzUHgNgXn50NonRg0+3JQTbXqH0swuG7
1RSYcf/t1XOOaT5CBGORhzhGZV7AfwvZtvMePTK3y1+/Rpb8U3paQZio29pG6uy9W7XcTmI1CCw2
dE68j7jaGbrL7qtAE1fD7uK7jy3dctmuxAfjItHgSKX4rYhuI7l8FYEHifzH+GDOe5pagYIB+5eZ
Cz4ZXd7r78OVcicrBEX+7WOrP+p0jwoXasyJFgJLIg2EMsE2fAiOn08NyR4CUPPvBBx0Ykh4SPer
PljT4UoCxnpgWjXm6oAVsCG/Zvnm9xkfBx8v5QOZqw8FkI8MpdKlPMJzWk72bMEprG6I9HPcb1WW
n6gB6VHTS2XPrt0vWiq074hWX/jOrDS0d1Tu3667Ah4kk4XH7LXDtt/HEjZ0HgCIocY6hULrVBLH
XHS/Xk+5/cpp8wauOHa+QE1xGuckWeQ4WxrAIExwGKbJcwwHlyCeoRlfNYs2HLw3CvIpJgsFl+f7
wgNey/yMrRQ7jdcqUfYzkiu3sakl+X2v53iVUmiX0dJzyhcZ6f7/WNobBIxmKICcV+9yyh2LZVvp
lrTvlBP2S4ns02/343a4f6mDJbKojTJSUz1ujhdZO++JAx9YSetRbSRh/Z0hFtMcLYZoy3LmPjLn
SQYIzqcZCgWrqZjcc/vKDr+5VKwrPRy/WOKeinFwhscLFUjuqAk+LLTKCqur/Oz6JUAvpLy7NfaJ
dEHWG2adjmyrEBs8MtiJHn6zeU+DkCArfUBGH1v9uRPZk3gNafdH5KuA7nFDs0bvBEtu1AnXiM+m
FzZRgM81PAPWs2tPjkx6C+cMd094IGhyo4I8Hm1cq33/0uiY9t+03s0mUkRfTgny2EqjKmb/TPXq
O/HNeH8sd6+76hxXJrinc6S9RdnjQ+aYPylxnVuRipFrF+fA0G0V+whMRtx6Fv1OmBq60HBZtbWO
SLVJ2wZ4SuKoXIxKIykRuoWADY9EVPPwiNkEFia8VCqDmqJQHsQr+1uTRbRog3CG6OEuGgoy+tXx
bXU4eGx9GbSO8Psbuvr8A9EF047WUIlUkDKDp3FBgtY4mZqSizDJqWdWSCLpkKw9Su7mB9BbzMz2
gNDOMDayzKv9/MpgJWwafuwtRFw0ATsfg3/XVsjSqKuQYtojwU1qwLbYsrrgaNrJgEsiZI7dUZoR
TEPxBBMZB44TqzGGO81llQ16Xw40NqvWH0NcdlmYmRcsj8YUrskmh7Kl5RXC1TQYh3kYf5jQywBx
x7cQIZVKvukRiNVw+9sWKsCoaasEUj03JqQyYFT+VtvrgXDgVd1VRUGA84K0C7Ds2VtC1diu+6eu
FdTVoDDKHlUlt72/4rqzhZ8jxl38P5tG9tsqTPLikncZYWKpv3MwoIHjN66/iORUjMTgTnd6aNDF
p9w9xQIRJ4Mtz8TsE6jGN5v4FlC2hANwj1FIhWBBsXE7YUur4FO5BIbu9bU5yDDDfoJRCEf3ni8e
XlWNIU+1qW5sqw+xUhAiAslZt2o5ezaHv6AA75sWxTndqdFH8P5w0BYWU/QeFNGTvB1nkwi1uEk1
P6vAG1Fof9V9q9u6ojthsdJ9qHjTjTlir0Y8j1Did9BHIQ3vC+SDt6ZtBe3c6arQ8kIKIhlPFsfa
1snQ0bD3OZptpQSbSl10VZR6oMUXcmUOldu1CIbwiyCpv4v6/rLT7tijW3qwMjJ/4nGXDThf8lYk
Yrx35Prazs7lsbvDUgqTCoz42MBJ/mO3ltiGQ+mypYkWw+OT36l72VrsvvPPcebv4nQA4SsBAgx1
yJPvHiwx0qYXmcPYQH8qmYed2Raht8Baa651p6JRDfO7XM/aDqhosoX4wYIf785uMEJ057Uj2juO
nrWNkimOCTpWhTVqPtwIDFEilTC6sODdpnOAopBHcKquYbSjKS5To+VkeWegm+KhHcSKHLlV/6XO
7O424b5uL82VavEmGal5jGl3X9pQ+r/K9SBtDiS15UarEz/zRS2XAw+TxnXR8vWk0qQMr7/DX3/7
kS3oMNmbtyv5WJ/Sg1/NHh+MnicY3VXy+4JKDOGjExemYBa96MdJms2znVyRXpQLmPTdw+m8nwGy
rGBJyngqhjJgMXhNhmupFuqlUkkMQ1+H1UH2VfGHj2qn3fVmvKvaXeL8nBXHLXvjOjhZVIFacQat
nIu8EkPVkzW6LZfe2IRgOZ64UrYn5WPZjWXg3a99acAYO5QtpYo/YYYXQ4+Kk80UDd0xbibWFn9I
hzbQQX2ADvkCKGm+7hEIMCbBvptBRNrtawuky7G0CbL9uA+xMg3+FqNByR/RI54Y2s/VAF/6fcFB
9BeQSrsuRJQYAo05f1rvWyZ/XWiF34p7Q4rGQuH+AJHuY8sDYCHVXZwmsriDo3QmSd+Pb5nChXpV
AieYJTR6xv5p890qq0x4jf2JFJBs2BTPN7dIdfUyQfT1f6lU5icVhQ/yzFBNXBHGaDhTc8ejyqNk
lWwZ33lh5eRqZJ+lH/2Id0SLlrnNVikxb5bmzmc2cU6BCdN9lK7rsS6yRP2+1AeP2Jjsyo7Ts4Go
7nqT3SxI6Jrk8G0xdj4T2hbtnNGbM75Y/tvxL5eZ76+Dw36+QnhEJne1or/mATiEOWdTw21rgBnz
7mwXkTY3HncQrLkENWNblOrRw/FW3LOwnsA56g6YwRdR9x3xnxiVoavyhpJcKUuPcklN0AeuL8Wa
3yLdphX0WAtBf3ORPy2yBexn2qb0qp1/75EmTXx7whPs4oum/xOkAunq1bpQjjxxHdoVfZDSn2ky
YHpvXuORoTfYWdcR9ZJGIHoL1VWS/0HqUvQGl7YrQvExp8ss7Xef8kidMy9t60nnMSXg+jmPM02Q
f8MbPs8mUBl5NqzjiIXd7qVwCKw0Un4JpD1wfUbVovLH7EgVR3sP1Yl/kBEUYAzZdk1xtlK8bl5n
/1BDzzSRZoY5vfYnl3DSyV2+/caT7Id0VkqDIFWkYdPSEs8rB9NGo1wNslCofx/MSSWKuEFM1gzb
qllRWOj4CnKuw6CFUYzn7WsNWoX8DZ1OWaOvVKOqerNl/eDTwiQHruiWk/KQQK9aXODosyUqqXWG
9aJ5k/w1PFU2tpED6VsOz9xRC+/c2E7oDTwwMi7QDn1tOH3dcG1L2qzneC0XVdvMb/u53knhGp90
bG2Eky7j3cWpJYFeWK2brS2J8KwAVJirJz7cziwFVFsRoa6dcJEhCXHS/NM7jsNc+k7/Lm2Y/PD1
j7ukVPgZjEPYcJxKQ0IwbEPwxMz3EbiQU5xHqyVtfTg0/8zDopvRrF9k7MRWyeBfjkMYNL/dwvK8
OmuGhvfRt4UuYnDuTON5YQvXPNIFgSHO44KD5NSB66jawz8VHzk5l7VytBsT0+jUx82r+DSpmQC/
8q0Z/Nbz2ULvFfdIpDgGZ2q5bRD1QMBYzx8c+I/GNZ1Fg0DQFGeLA3CxaDDtMUmOLVrpGjyBmcLt
mM7GqZ5r7WXJwv/eGWw8dGbOGaHwii7C5HfQVvtaklzaMFjs7jT9H5CDyYbl230YnzhiLEpLi1Xw
IkWPBTQvQ+qQIZfc4WkYaZgH4KVnYs+6HMHIYVQot21645ciEhnl3DASrq8d8eTJAVfgmE8XNokA
5bDDXC7Vz6iVFVQDbiQU6cqPu4ZXANzSkgjaeTz+dBZEpFXyFJhZRZ832wN6IVnhCAEoYKqMkKwq
DHLjcCmOVfTjBPyAevwgTJhLkVuyXtqn6uHqU0fUa37dYgrCDDwiNWD9VKAv1+wNS0YWja9vjlWG
syQgohkZmiWAoEXlHKrLkXP8PZizVFd4ttBLP2Zi1cLuq3M/Ndp2Xf0Dzlwu7nokZDs47QxxTj5M
FlnH5glD5pt+IoWadtgoWrK9KoMz/sBwA29M/KLDL7oPgZFw+Oc7ITAkSZmwUtxxNChPFIyxf61R
Ho90QC+rpN+NE2xNKTCSVg3UUkEFoAmHdetpkxbe7SZM+DS4A7cjtS5n1SiTndl5tl0UIif9zjEJ
INMr0JxgCfxpCjfVtn9gajq9OZ+9yUzDPtVOIn2EMNK21lpDGyLvTG17zIrcgTDoEuLqmVY3becZ
H5nlGyxaeF891/BWgNUJEU7N+jmELnDLCAbXKcZrK1VQA4+2sG31sah1oFEFFgHKmJiTCC2dzfwu
6E+9oAH7M4aIU9XEb+wVGLrnxW47+otJFvcQeojxez3I+zGP8LZDpjhreey+LDVtg/O5RRzsvpVO
c/hL+shG9JGCECdboLCNstEFfa1T/ScjDd2KjPzWyExXtTNPaDs/22tlHv8kBNJMH7/Ly0SE96B4
OCVR870Y/g5ZmBYzFOCOPmJSsZQ9SCYC7KMbLMZmjvPsUGJu/ihUjAaZUqdg52MVcRQntbK1nMfA
gH5XT7tnspFXeIcIYFwtmAf9b2rAu+EOi8r1yNh6dex7l2lKiDeDCCpXJePxZKTQBjIBpv/64KDf
MZKGxgLYQlo/kq3K+tx1YRjtBxigXXjlR7Yty45/kXThEAsdyoaOQT4Ag9+8ioyEDqOSAuloJFeT
ecjRypvuxtB+ei3lGIYmPd8MBSMPWPCmOLtWbGJPPmSkD0nBQ3QAZXK6vlC7e9g47vm6cECkg2Zf
Y4i0o+Eu6wYggs8CnSmL7zvMBKC7fEt0UnUGHlb3+jQ5TWhy/N2ApX6z1UAygzJjKWi4aijPTwae
qrQ3I9RHWtc5xjI4///PFzKabWDe1DAQsmpJ+R6Vs3qfHbMngRcbF+drJPohbXUvDyp3pMPnKbJj
pFmQEK5MFl1i9MujdTRLJBepcKEDaiyTs/nshVrYN/ARI5NiyOp5gMdBUtVAxTCbyUxks4ZTzMdu
Dgtafq/u8YhME8neJE6OBhESp350H+nukdGPEUuFC3mxRDhAE13PM7EIHH6EEbPKjDRsIWBxpBX2
yhSS1nT5AgW5s3vETYfY8lXujXGuTojRGtf1tT/oRWpeapJaaj7G5vPfQBtk1BD0jo2mdp2ID46l
ZbwafW7mFMBkqQNntgwKuUmj2hdhe3YTj/gty6kkMNXHNA+oqVP3vw8yMzeah5etYx9jS1coefmv
Pf7JOxBv/jgRp3ceO6w4GLzIlO/zDc7JyDywLxXIuxfkqae+QPgbD1xuEB+gynwgaD+acbULSGQe
UnNnBJqwgeSIMwSEz9G6UPDXb7rSOdrWusHyNe/99VbxDRoZFnFnP5KrFdpx6lK6zAAIM8VYizNN
+iW0ayJ5f3CxlluZxlmJszi4q9cDqdegsqOABIXnaTCBpygTKg8YLZ1sWOk4EgbGpsgF8YzWh7CY
2/Dh0DKkN0edNd6lXqc9ypLssuSl0yBqxp2aBEHNCknui2otUyz3nwhd67M4qNqe7Hk40ZCsL+FR
q+q0RU9W/t5Xdu8qSGEXKaK8kqFoig7P1WXIIabq6p1o5OGEYO2m6lopyKKxRWpIUotoNUhDF3/0
9mHLFalcQLlsYZznoxCPWYQvlVDAdBAKMKfiJOPJtIg9gDLjG/Cyr0AcLhKzSqv3EhujD9cZAqpl
zXUcO8BHO6si7Zttu9JF9B00qXBEMjmy24/Zl6WyMOlu/nlBGpL7EAH48d+qNy9/IlW3A60s4r+c
PIWplY4AaFTt+v9rMMu5smKrF8qPL9aQAUsZpFa/ajvTeksD1EOUT3LchQeyC+oDmulOvs97tpm/
W72Af/hfxnl/xIF/2lkTrOguHr9wQRysKlWovMDlUAeWDyWSVUTyS38rDyZCe2PsTpG/gVOZ7tBH
nWivDQWLDV2hDBX/yYBbzmuY1VaQcimMryU2hf90tL7xC0T5kNL7zqlDdN8PIaK2COXa6Am4jZcY
v/ROHt4Vq/OoiNfYkFFIfJiY5HzWwu4/S9BnEl90GO7EN1UArw5tBMepcR5KUgg90/Mn8W9pXeYU
EYKifcz8SVMw1t/eley42OkZUmWUuFEswq0bs73RFhxn4MJynteJUljkNPxtE18juR+oSBA36tzD
H7jmr52AXm2B0xozncPqJRTqMaCag0hR+xd6nBAM8x3NZ8QgtXSez3OgDT4eXJFP/cEbitPGVEic
ahgiSGk4oTLq9o8oFdqYmlF86D0Q7swb0Vte1zOUSA5aQKSCYBgeDqz6TCSD6NIkhWJn5YMN2cXV
DpqB0VCiEgGF8ukIYPq4WA+TTTpGAfbYep1WOA1NfbCqbLgmxy9g9+mF585k2vAscu3sktZ7VFa+
XFbHq7+Bp7WxQKjUSP3F4zYVHDV2TqL2jOgCd+lkfWQHJGwjE4v7uEuJbsu5js6smitUrVJ241U/
+8AXZ3QESJUD/SGpPy2iSBKmdSqi1M8ohsqqGZLqQBCZh+IpxQ6xCvc4zXuw9HjyO/dBMKa0uyn7
K/mlRLA1q59WdrHt5B6BTHaw/wD3hztv2pR8pFmESR8RBUEipOSMufhn5BR1XDTQMYmUyvtY7+zv
dq0GFciIDjHNPoNQUafA/5rO+YAA/aitAkwcgpSjJN9vKPI/VmK5fjP8DKrgjXQ5aW2MtolmjLdN
FFxuZfJiaTHRsYpWHjYoQTZAptXZFbpptjRbvbEW/pat7wCANBV/cB+d0h5UFsbPW51N4p0v3Vd9
QtIH564C4cGZIC/0ur+qgPkCH8Hv8G+qCi1gD7fXWE2r3jLKZJR5U6d1iWYOCYyLkgbK5JyE7mcb
OQBG9wZt+DRqy5+aCPa2POREc43CXdz0S4O8iknSyL/0/iTvGQhomQa306f1mKXLLj2SLjO0MVjw
EVcPchTILEvFUKkO6v6X487+Iy/4Kzwg/Uu9+Zum+e8mAZv3k1ts6ZPWEXN/I0tu8H6hPCy3UOAM
Wcv3LbkG6fUZT4LwYEEzK7bYKYI+rZQMKgjt8+9r+Nk3HbO+l2j6g5j7SZaOPHKA/LwjqKR894Ee
E0FCIipl4V1FeBO8sbc0W5/fMqyuR/shE8OknTYGPJH4ZPHkCReWP9cBQfWfqGxAQdhDmb6L9NxS
NtZq4O20VULap4cydM5X27ynPcxNo1AGjNSpRbBgZFauAbIKC1OEjrqMSglTuBiYvQahe1yX9sz/
2s3FQ1Fz+YytE2DzUg5xBqfwy7d1fT5Qvbb3v7RNAcqAFe3OqhfQj5XvBPV8W4s18bkzw9CoyWnK
sCyHqR6vuxwmijOZ2zbi+sK0mjEQIaOtc3sAV0wrv31RTnK0GGtZU//4qDMkPoZy5nhlyPWpn3vT
Eat0IWhgbz2pKuboSHhWiv3IcIvesFVzeBJ3XifC+zF5Kn93ig4y48MKYGoOSHHr+4Ai7gNx5Sm2
UzA646rr4jVzeZMXLjTjtSs/ZdVj2ECTXVC87ZOU5WKhOOZ1zXMqQRheN3A+1ND23Czjaa0ryQjC
JLUF+Eb41qHjoGebApVSKFd8gz30keuzUEoLcogkZ1IM4PhcwxKb3qQRbHPk3wcVd0aE6xsm/f0b
tZqHflw9PUInKZ+nWCv0XWCeuA0bY/5jyhwvG5BwHRkyN2GkeEinRdPABuqESDKqw3YQ+nx6+Pzd
bc93thbDrQzOz4gkf0rvBnbWce4oLIcnRciojFIzm0QjElP212pfsvbp6ttiXyEslgrI5ZXHAWHk
CMzOvNsB2C9EPlch6Uc0ogxr+mdmQTUGvI0S8EK6vEi0JmDTPmV5XeovgOrzcU+bjXuhQKCW/6Hw
aKw0aQGqsEl7G6uJ421+G5J9wDL23rgx9j9Pg8ab43pre48+gzvDKnPh0MjDxNl1aA7tLkDVoV9N
NupTARYhv7nsy1HIZKwEIsvrKE8U3NQ6unSpLhjSqJ82uaD+6D1jU3Yfx8GtvE2Dpfu8TgoWirab
FoLMNw+LD4wJGJmd5ecaF9fID2KYzSqoiAD7LoH90HLcuMtzF5FDJsQ//KuJ7RbQxgrp6p7l6LLg
BDBruw4NHCa/NGnN3ok2D2PiI/G4k8Q/x0ubxweda0DboGi8eJcTd7opFLNUxM+NzfiaWiozmDlC
AVqKf6BJXEheQE0VxPsIUtpaxbA4aNyE9WTSk5fXf+l25kXAUzmK+/Qw6nsb9akCqERlC8dIw/6L
2/ZOCJvUpvTgeDpL0kc2bBirga8od943O2hm43Ef2dcA2cChGSnGPZ0nPiu/1do6Nq13kh5aJSbP
xQbawnHOrDYjzyleS6bbONvRHx5jG3mddebmP15SBWKx/4LJBzE3+CDQO8suM08BnO+ub5HidHlf
0QfWyv0Jes4zeqqrxS0qW7pqzdu0JdBcvAqXH4gb9jgky6nTypM+MWFi1Mfl25BA/mw4DoYnWlb2
w0eCW4oplHOEhjzmIakOk4krgoSt8JgebsXYwQaMtp4VfOVbvUVAi1VkFMxb1iLcvtRlatOReB+P
4gqosvL+EeCjLTfOQ9YtZ7f9nxOrrgd9P7/2bfqkAu4c1Rx35sjAZL+xc+EKFSY8vZOs0dHICFBt
xpwWRN5ZzPcIS/qfftRqZVABqCrRhv2M2+hZkVwqzP3l9Dxd6t+gMcIahWkrV24zRLqNGm8Hj8Ah
SNkQ3IPGInH3czcx2ny6hTmb44pIa7ELzDANjSJTaGzGTdVd64+Bgmxy1ybgx8jVDkW5f9Kx64lA
IHqDvcT14joBaotk2ToG4iNp24P0psgSfLTTQgTqLnWjCNcbIPfH/kJObsevGXPK3PdfU3KYDTGk
pNcQJkuzTgi6Y+UET4LY5B1meWdFb1HDPtp5rOL1UlRbTyXXHM968x2opSHv7mE02aiI/MEGjrN5
z2KxFK3N5TgsUgP0ZMtfXddEjf+tGA4kKhu0eCmr1tfj/J2/qyekAumRu2AlqOe5nNnfkJIRx8NB
RXHEkeZ/g1kpQ0FvyE38OYeYLqIlio+UsL16zV+3Eez9HwPuvR6Vv/WNVDL61ngAMXnG6oJ6pPEV
JKi5xDXO7pDeGMiJSnSWGhiTMOHtBy4oDDWKa57HGTnpjfy/pOjhUfCDTkQhJKdFsI5C8BAWoLoX
Cz+a6XI39bW+hNggz/uT/88f0onDBOwLSUFIPBdO+kXIXbnoZB2Fv0yM/fVaWPTtuToh3I2Ui91r
1+LsVnov8OprHLEvvKheUcHWgMs6WnUPdyaiggRWyvIb+8jk79ZfUoobSPbEVEHSMmutnZ2bc0i6
JwfA2Z4lZ1NmW83ApYWReCnmelErtnwTit2ADOp3LwWYTq9kwebfMF4z+eSozJx7gv8ueiuLtmLM
oEQbeN2q7pRWmYKaeJ1wOE651o+FML0u4zrMGiCrScN3cTSj6DOvf8ryLb0E7vQRD3+Hqm161cBj
w3M3vSh9SFOAqFUpJfN0uh1O43x34pf1fuXov8E5aCbds08jn19VUhg7Lhqk1sHuPFdZW56ui1Jq
ha7ByRtydExJAIamG/o9EZyZQtE/x6kuo1Yn61W5I2mfGDYebQnBFX7fmJp3zuXDWlfT6BENeHLw
ajn6YZBtXI9eWLMUi1OqgtlDVMiEM7d/tSxCskMhRrNmR1R6Wj7kEuSbbFAO4nSlTcQBiSQBptx1
5SYT3TvZli0FHl8p4DFBKSdFVAz8tR8UdbD5rZPdV5S41lC1IxDTLLy66D3tq2HZN5qwwDmRhBXn
1ciA+k2j59D9feuggKm3D5erqtZJlvJhqRzE8cyFkvd9jpdE2hLDZureOUjUiz48hJ8212V10f9X
je6bwlcSWThTkZPMEhWEYGTsxFgpkgxYeei3e+fXwLlK/fNkxcEjItVYSIIgboBflg6AQQZullxK
LInfHRBfjVrKJy0qEN3M8G4FWeuUAzauoW/zqqFWjJyH4ImxUS2ijJfH5t7Qn8GA8ai5vsnfKDz2
FwgB91ezp6xiJk+k2QrvXDFMALXlQGh1x+LMdgcYsdRrYbMF80wZHLHaiqXPiEw9oXgJPTC5uFkO
vz8SOYktk+s3uiEmIMf8n6KNRvdvubNQ9WtJ3cnchTXSFAktpaC7AGzl8vGSwSroQ9yQ41llx7Ej
4EHNs1oHeIF3qV2PYyIjzMVwIV8rAI6e0okU9+qdARcmj3WhdFofnrnwYNrOKZuu2lCe2XLA8Kcy
MoRmbsSqPFnWrpmlY8VRaFh0DxxxL59bZHG5l2pKPnZtQPhJK0m+HL8p1a1nPdeQEqYtaYcFSkw5
n2ssgw2QftYA6qOk6xiJodaer9Z+dCSlkNYxc/qYlIcb/kGw+KY6BcCa1Ga8jTlumSYNk+LNJMQ0
4a4GC5L5u63B1LTaqnAyJCQamqU4HZl9IEepWetQtIJzFLDw6jlfMG0r4gpVQuBHO/vXlr3V6XZ+
UUXzoSIbaYV5DOQsh482jx7XuNMVDDOM8Cma7Vz+PYyOzOhL468vwSFcY7lObup+nBFK8Bm442b1
K6Nr/syZpgEDeZqUlqhw2beC3JKutvr4ho1ZA1PhoNkwMcSRGEgVH6m1tLRy3sYg4qpE6yqnwZOd
KHrGq+1gP6ZmHKCD5nrFlqECKa0I8MYyNzbfnlY1YbYc2YeI2P1S02+Deoy1E4/b+wP5cpH84uEL
R8gAb+burTuUBXQeGYAcTx5eInnBwBj0H0whrTij0hxpXM3I1FGczsCzPz6nR3/kgfJwVcnBt8Wd
bSWtsgYXfIxOseRj49fyAiBECBRSgL9YBSBbd19IyZxbEtvaMJleUJGcKQwyTXuUiWIcZtHr+yJJ
48QUl/WNQiitrjkQvW5A0Hg3Q41g4JoNqIreI/6SP8aD7720+sZd2oaVFzIYXBMva3pw3B0EvISy
OHWNNmEoPiuDdo8A5uyqE5lSRszToSKGnUrFlsfbuWRUqbOSMwXo+Y/ASixAHM4bVCkz1FG+0kKl
hFA4CI7YvNpUpYV4nD3FFo1fEXO00dymq0kCd4uVleuekt1hiJXqkmIEOCAsNMlRcVQwsQ+xHzLG
o44Rkt1gpgGRvl7W1EO34qHGxdi7vlJ7vthHUjHmETBoZ7U6n49qNJos2YIYal1qmdHsM9VqKVH3
lYg7hk714hHqq5qiQm+2zgEPXMpajjZX3cc5ofqHJwh3QnNigPxj3Fr3W4E4chZtEVu7Ww5CPwIe
NHUv77o99W4DEuaQs4bkwwj4yT1kARFEBW/Y48Dei/NDyIwB3cJw8BMQqBnOydO5O+HCUMTCihFB
tURJG7WGdGZelXjt3/HWPuf8EWgBCx0y1WXcMoTt0H1Ftog0NVheD5gCL0nVxPeJbf8UaIzcIoda
1LVRRHFUj4m/0l0Uog05ND8j6HT8ThSNjdEUZRTD5bOZMLXqIv0PoMe1ktFqAH+sfNp9/BkDOaxm
u6suu8Di3G/x/e2oqp5EEFMsI380YTPyr+P2m2ELTgWJF/qeC6wjf4a4Grc1tRciHsijst0bn6WV
e7QrXay28PjGrpB/pETGHCLf+bfQ+zSAbM3rYOwXSbA4OHJl6XvOGYPUtR9bNYYNM8qwYyP3dQ3Y
bX8Yc5SdjcETj7n1eWsi74jN1feRvSKeKuO9re+jRqu4VMRMpgvmjiHgLvGuNUTxCp40FezRwD+M
u0uqLSjDSU7XfkwmIpw7riLQyQAKaJyC4hWJwBLtuYLrD63kSwsFdgMrrMHD5eS5bY0t0VKLNSx2
P1eA6SXttMCXF0S+3BS/LjnaJBomi7ZNaq1WsdLo/Kj3zK1xdW3mOAE9NGOAi9cwn99TEGacwRHe
gn6jvbQEB6Wuybf/lnQDEM68KLn0sYIk2qzUBndLIX5fAp7IiTEeIPWhOTVEjGFiWT62HwRvj5rm
Hs7LvWQiCH/eYi1oqjzCrjR1yxXOld2FvNq4C/wnUH9uQ3nk3Bv6nc10Km5ecDhYjqB2wfg9k/ix
ns97YVx2OvjgErA9OySNAA7ehxNhG4ehKGjnfiHbLDsLnmL1/RmvuE3a/jXz/QCnnDZLYDxLESHG
Tq9IYCbAFjrOQe7KCCqEYiGf/61ZPMwtR9ZmKTQXmKqZx8VoaOm/a4P4W2EwjdMa100WG6ZtIQrV
jquD7sapZ8gUw7l4AvBTG9FJ0f31/lsJ06FmxW0jqG+Ll/RlrAXIenDZQyBMs2krDk631NnxcBbm
TXnBmJ5yQbpX0D7yHiHUfTjum1lBsjgsvJjEDyIFCuASgLq8zTy1RnlumPQt25u8vu3m24LkuFwl
enlwv+I9z3ePAOMlPIVLEHCpBffBNMOrgb/ppDAgjWBi/uhtmTqfFFk9nq7sndIa4b3MgbELTOFj
kq76zVbeZorMK7aJdgCpKLHyE7EXDMk/58r2Csrz3upr6Kbqg0m4t0vp/qg0b7nCFVy3HY91un68
4OibGi05ac3llackQkmrrdWKP+2J6LhFdLLTkn1FvazjhfqoXxRytqb/Q7iTs2PlFTUXkafoHx6y
wEm88UM6fiEvRA7yAIg2Ay+0gyky1Er+0Ohh/MPcdPU0ULkPRQhxGItjgRz+nWt3YbAa+NC6hhMi
f55YRThJDTejFzl4vpTmucBGqMJ1rb1d/yex0uJ7PJ24o2Bi7lqnUlLph8dKox9MSrmD3rfEUG/C
1v8h75sC8iV63MY2z6PsaopYWOE9qRZx3JBVJrM1IgOWuQjka183ylAKfm7KPs0FtnSx+JXToyqp
/OwOd2FyLRQv1yEOLe5+MIrG/vgGPn1yH4CtHaHBi7aze9PpnQerf0gMPc15f/YimneodUluRbdV
yRmwCuf+G76Pk8Zgt1qQv20f+ttK/ioxnUVFz8QFstdKO1fgKaDFeGR6YaFcua9BF2uYGa7qxLeY
vrls61kjDtwR+1cI98YhPJXzkjdaqFwYt9yGt9Rz9CwXnVcySTUnG45Y9bA84ovota3swxOdvnyd
nd6hneCPoD73OSuk+mkyVM6SBjCGFcM85p9Uv81HVKHDlpl++59Il338oxJf6Heatw8SW0DEI0Ah
m81xa6yMQukADuXGH0QIliibQ4qRbWyfI5z2byE1arJeHTdR98QfZ/HQ3jCvunce079b6DJYaCRY
R4pyaD4S4uVZKJIl9sg3pikniLbFspDpZXF+osvR0q0ISyFACw50Ve+U1MTOOUEZQPnvz6279Rre
FJC5OW2vjxAu0YG/2HwgkqO1Btiwru71A6pRF9MxUrqdGap5l/Qi4Mq0L1WyO7OXsgBwOfUHcHiN
XGlhM7tGignBFo/uC9FqnO0wvdWABWFNsQaN7yZrs1iJUFE+1gh3H+nUWLZwNPTRpp+btzmlfHBI
8F+bGNrqIlsj1YfbsNX+VqnrOeODGd0P3AiXfcgv9D5P26SOugl8QY+iX8hTEM4qgyQJtvUczCAX
BTtJSkG8gOTLSHcIQVjaoXNZwXT+QZ3J1l4j/FdNddDvDZlC4gnebESs2o/dt2YntpqICWNPrsAO
bYeMRfPB1kduEYvg39bv3vCBe80po5oTGDTTbmhgcnkZdnZ2tTW77dwSMLV55tpGrzSY0VvNs1GH
kou6wIxDCUkhw2A6CeA1IKvYmsZicJ+BX3yrC2TAVPBK2lP5IUqI2j01LUhN+Gx8ToI2lrNkSQmA
Ao3XCnM+olug8qV+XqsRYeBQaxPkUexIg4kgRE7rp0wRpVahQKL81sygKVHxLNqgUX6d3gwKlYW9
GSYlsIMKCxqemY/zeDEseh6HS41dtwe9Ak/+Qpxtd/afqYYyZmoCY8XR2VSzOEoVbbaa8FFphBWf
Y+0m20sPwGFZ7/VbPr7Nm6crnQmlNUHTR/66u3ojk902pFRGGNwJ0eqD+OhaqjQT4LdYgX+9Nnyo
t3AT/KRucrqSyM/G/PGvQrqhv6ma2lERCWou/WbBCecgTZdEsDlev+p180qIgdDCPtAawzPFB/TM
RWZ/2dXI7g+pWZczW0g+mGtXbDxSoT7Mm3MSHcGPSu/40O4Hiqu38+BxhI00UygsjrNkEB6RANCL
+N4d8FmO9MOIuxhjlyRcqJ8pVH+6eFuXGn+V4/huks7JpHT4D5KSxpjZGmDcvy5dHIBAjVm8LGz6
Mw1ogAWjpv3y6wZdHnYhJIGrc5SYQtzMV1EVI4SboynAiFL0w2gyxKDIgFfWA+tAGoWKuJIs26g/
qGvz8fHK4aSc0x3413DiNHgp+1qSE/PHqON2A9w19qwjS/UlsWt3BTbyqW6EI9cvTmEq2YOaiKYa
PO6roGDkqxywWXJaa1G79Q5NzeKy9KfanS+nbY5l8V9EvLKqMh1CkIwfE1q4PCXn//f+1o+NGUe8
g7ILnDlT8Yh1VJ+2akWZumvvR4S7u73WwatKB+RxkRL4+wyzuSZnBZNfTYGLh2vzJeF+10/jmfil
8AoEBPH+1sW9zxCa8X5nnZYlPgbFjv2avGYlYUYetSvSrkBLxyglaL+xwrtKdai8jiRSxlTDDYg9
rFeqyzdUgVreVE+JuyuzFJ6qUvjXxblv2nTIzoVzZhwg8Y7Ain51OCTJGt60v9OWdMXXpBdCOaYH
/6RpbtH+Eh8vvcy98V02y9+op6FGvjxCjAcSQRDtnSlC8jZ70oAzOCjc+qKk7NWEoFbyP4pa8mVZ
0rTO1iPtOqiWrx5Gg/Li0PBMGgZT/CUMh94z+cIfdm06wqbmMM1IGDKjmJ1dnF0Zm9mVt8stXCt9
5bmEjYVeNXU/yV7qY7lgNm2j0MPAjdKxcnoCkMBFsckD6/z9Naa5fSxTc2ds4id5kSBWWQOeFRW9
2cl1ph0++wXqDbYYvq5gCuckBCMWz1NIxml9it+sxk1b/WqkvnwM+uMxjgUR1PZR/9hdACextsas
g5wot7NCED7N+EuieAUTs3fWj7xVbWYu+c3CuVFqJr3ay0Cu8Li2KsFIJdGzS2TuRJg95zmFt9RF
Vj64QhMJkpRrInIgKVyXDAxSoSyfVXi/mO7nADs2YdgW0TG3FZXNTy772SLz+fQxzdMIS/HwObup
Q559Se401toRwoafrmAhEVNnkpEgdI16r53K7E1lKQLwEFZCmh5zHv7BA5zRT/zZBBWhdhSlUKGR
0BtJshNRYV6B7IhtdptcbiFK4GkQM9jizI4vr8YBgGYsbhZl14YXQsm159uRT6BoIR+Z41uCaQke
fnwZR4drczr4S5e0jX5n5E4T45XTCnMUm14eRaYrfioKcfYpsd96/yCKGCjW2K2HWN4khSsW/cPv
FciPOvkxN6YiVm8eMctt6UDakNyL1x5qxdnS9G8tsQei/e56SXs7GJ0UyoksZR0KJzWFWj+A1Q0s
9JybJWu8P0JYRZkqC7NSGv/BlJC8qQx8MaK7/9RA6KoZ2joQsaVYxDM+ar8+6wCDxS1R31msdiOQ
OJaIgitK1LxsLnc3gnwLGGCRNb9UwXJWJ9Bzhgm4BdA2K4F5Ta1PFDEhgBLpzFlytRtuUbQsKqlE
P8mpnvLZg7y0Ux32UYhzgHNnaiWCf7LPDR0BK6daq2Cs+3jB5aCumZ/+EVk9B9b0r+1Rm3AfwZqH
zbIAwUbwIdsHh6Ec3golYtYwPjaoZLRk+EFf3Ov9h1DDfUZL9z0boikjVbhcl3ivnvVyxRuTwCqW
Rf7CzTj55pxYQutdTCtxNmppCIASuTOvMsD+IDLd7CFHnhiVyujpDjGuq5QYkKWxCSUGtg4AzgiH
A6i6O0LRzsPn+R6YUc9or06jFVyZVOms/VlRtMnCDoPyADgi7Tuf8/oRlR54yZwPfObocSiHpo0A
1FJaWia1kBrvSXDKqdoxH8sHG6fpjOcgly7pKUAvj8VP0rxcWJ9xcPVLy3WINNZDTFWxqZ6XY7dI
3xZJuKRABa7TSETQLJSbpizYQ0H9knPfR6LEpSOj5+Mm1Vg5uFCIZ9uPelhcSD0aRdqyBW6klOTr
0vm/lPNQKKI6BNrTTKT5U4O7fSZO1Gp5+NEZINsCnRpb7+Mf1ydbuP7BZZDtR70j7xKjq7YXfX5k
1Is4BWBW4MFlJ3LqVzEo6UR0gvOYVDoXF/muWBeuMzB0wjFnM5y+iOZjZU0FEIdlm+M4lM4qmHxm
D0Bcv003tN4pf1MGOnqJtCJkPKnduBxlV06NNKg8pLx24VUCQLF38vuajyHnbFJuL9ciqVljgfH6
dVvnlrGHmSq/0TDjgXtrlC1Tjug3Ykd24RSSfNcOa/HP7Gs14Ja4wFPhXXRwf4+nWGrlkHACeEnD
zX2Eaiu3+s9FJ5x0TZlLlrO0+C4g5egU++pPsBOBNKOfpbjL9WnheumbrshlQkKZGcxCLTDf8hzs
w8mhJcNfUsk5HKKbj7caiCWVJp/shndikDZ/wS2FH5CORmBz9EWGFtxu4il72pizChta6KY8sexf
eRR7t4A0dWi/RLL/OsPApkLlWNhzK0khrstB4vC/vZKaYFA26KwiY1X9lHJ1j8ZqS07qn1VYEJ8+
mXYFxB0xXCHwmBWNCw03fI+jClrboBQV3ok/yVjg2IxDGHgj15dkoggLNbXETZ6/xRzmLsgMkVG/
X/dOD5LWYfL9IRQOGvoaRWRshApo7ywDC0gokKuj4JP5fUGBsraaXNg3gLh+SivpPOFV9Kojbwk+
ie8+1pqiBSAJAKuiH6KkZ5lkWaZGE8ebnRe4xU08Y6OOTnxBHpH4mMPcGYu5hF6RvY+0r6YqEkDk
oCAXuTf54hVViRelIQxUkLUizktzm/lxs+ORRrzeUGbV3xkY3Z0JJBTk+XZ74GlcYlHeRCssddVD
uQU82y6nAi4qhvx0umzyIgk/hU5GUCV7ksQ98mlFQibR+pWWwCeXfX2QpPnFvLk0WAW9+SAfvCgw
TXJ1Y6oIZmUYS0/ROB4fVYaPpSe3LjMN0G4CsDxxb4VcCGkFI4jQuLOcRXj5+h0bb3Vhg+MMSnae
N+U7+RXEyLAF4r46809t4W1b2VDkuZjXGvGYAmBOvN6F9ubS0Blv3NhNCTgcrQWAcd4aTYUhYlii
HJ7SbEa9CeD0KsORsH9IMKmayuQM6iqgIMklf67lBxn30mPhNDKJaYU63ziRpqwN/wChX7nwTRHc
zOb5pg13V9gPa/7tugrWP3EpSHTmn+zRA7uVueS7PmHbShfz0PmDGkvbXAlOXBdmB11yXgHm4R2q
Aqz47wCWy1ETY6BLGXk/MWsSaaAnKKhV26IniwG4PRjkrwO5GK4dkSvmI4y8T4T/kGBSdayg3ZMr
0VtekEO2qdUxcMKJAVWJJdejnJau3qG/GRVttj1D3oE4EhfBl5Myrb3BP0ncjNyGn12OKfkPD/ho
gO506inkHV2Ix2lUfPW4/NDu7Y2AjxGM2qLaPqLQpgAq+tw/vC4XGvI2YzR16HqASFuV8cDm81GU
3IrzNmBTePTpQV00yP7tlEtUTalHXsdys/9yWvUAkcigmEyGLCuhDRqIdaI8kOg+IW4M0M5r5vOY
XBUkQilZGjuAGuxRFUywJLKh8HJGUSiSq5FeqRe6NzwoFA2XRYMFYrtaqtxw/z6cXrw5vk15RfOI
umwMR7XTnwij8sq8R99Vx6kyCuXe5o7wRyyj6aQGKruId35tk7cZ0rzehNuGo9Wq4F86kdMMQCbM
TojwZXjRa4yFRwfyKdceA+Vfd73tTmrIuHC7mgGHdbx/pvZ7LxpUPuyIFrTNPi2RqhzAjhdiS62U
bwuVzJexJsz7CbCFlEYF8zHneRclrrJ8AtKq3ZR2m5a6AEnopMPLlMokdYNkfCxY6eQydP3iSJ8J
xczLbWTijW2EKzgozLQg42hlx4KMInPJnspS0SfZI8Y4SDy71fLuQkAVAROClyEC5oghCjxsCpZG
pKKtrv+iTDyAIuPfbE7926Qcu+JA/7s35uFZkwX9zrVTgIgJ0gQeP6FuQdafjRS+8EkORA+/Msb5
y0To86ZsJ8dGJ4MvpxunGXknv2yFTvb+C/Gcz5TEM2kfaaS42vcNjp31CDZ7zCeuln47h9I7rgKb
4m0Bc+oCrVZc8w7GGcuoStR5rBoU/WssG5dF+zTS9Nj4USBhlp8HAdSHqIG231dRx418umNHoLcE
XGR9fTShIHytO7WOkhZa5u80D3dOiuOO++7q79rqeMWfuWM3B+D/M8Zk1j+ZhQVI1R+mxmn75f1h
ahMyWXAqKbwbX9TP7zbisEnzs7BY0DnpNOgQGXPAd2AWvZSl+jioND2QxB4uUf8gvCs9iWJXkt+g
P3Rl7o+lkYKLRbHwXtc+QaUAbDxdybCjcU3xxz2Foy4TqaaRWnXgX/d175lSmZnvx+VGxWVCJd4R
8Y+9ugqCp4LtSP73m1ciHcx99WZhpE9etseo9bSVFMYQH59ltn7qzl1IImC55vgHDBeB/Gz+f6E5
SRdLqrruY5Bltsg0+ZtdCakafR1OodDPnw2XthVCneyViIq8l6sGrrexunnqeLxOxIKrWZCkV0da
FQbGqmkyO/0o3UKUqmehU9QtgsKR/q6NMBxk9hj4hodBf51Pi/tg4CpV82NMkXLhRA0wmS374r0s
9eyciLBcmTRnof8HH3vul74o8ozN9a02oDpQnXNHiG6NBFTjtzFRmVwOtIJZmTFRW8/uL03wjJtZ
EUft1n+DRMygFE9p1FzgGNTs3RBdtUMbtd4H6grt4LYMV3C6JQjf6AjnqSnQJ1s1/pvEZH6OYtxn
PnX5xiI5qQu3IN7aE5RqKZX85k1enbAA+c0eWaoVgjT6hwI+7qb0OXA/Ja/zHRVMRYTCp5/tAyrg
jrLpfk5SUJFeOLlissPtgy9BUB+zeXVIiYFA37VCLZo690zuJXikomBkONdDGIOs1cPwFnK9gNTR
wB0LlgGbhjsKSxNtKi2Dx74bl7+SgyaNWJ+n28zGlUCusIT9Dui88plWA+Qc4zcNoKRy7P5HdS7a
Bn2YukdxZvpScNkCVOv2DlZ6RXGvVaNrWW5KQGs/YsmFXHvnv9pG7Z9vvvDG2XIsZMURkHq3+f+A
7rRyPwsH/p3POBhc5ZmEfq1q3MApdRveNB0FmEQwoc6TYwMSCSysBH66KYXsBnwtVF1mVgImCrTh
udn+o1A7p2hGxQ+gdVrjNvyjDoX/gxu+x462JbHyIcT1Xj2Fgn8IAeVjnQGf1vRB1AiDSZcSyHwT
XXg18jNN2QkO+fuo2tl8XAPkVhgeZeByZ8CNr2ypkPjIRyX+0dX3nNsm6olIPa4CrDwWBMenvzrr
rrEOrZmory78bVTiNT4bkn/+d/wlFSCdgzbV720m3jtBI9mTDR2OULYIv3PCScNjo4+1mwtCwMcq
5IHeTVkz8NouOSzAv35hjDfJaqTluUhqSfFdKat90VG1ANGELWMmrIRTV6g/cIUVSoXtG3Vi/WQ6
9QzC9YmQ5OLjyJIb5LKXAIh8b0I4CyhVaLyA/h8k960N2Avu+0j4rAkqQHBxa9DxWodlJoXBbqpt
6wXFNepDhql58IWSP49hpMmhgSyXlrzknHnLdTNkWTnfvJGlcnBtVzjfLVh4JyGv13iQiYvlwezs
zrxpsehMt7J72ddU7+28whjnr81bla+gTTbWTPFsHdZjS/pLG6k/medr6DBorAB2nwvpYftMhHZt
OEb6lr9OzqnU6F9itpUDeHzHaGtF57Pfv9gwgZny1nIyH79249POziLsrlSI+qLg/HZ566A7ei1j
ZAr0VuwmYS4eQ4vOuR8qEe5p9HKlW4PrCJbEZBheS1wR1Hx4O8KK2bl1mc21augGrzcQRmpBTXgE
b5msXDdvYRlre76DaADucrldJqedrSMh4sWm+5xTw4pmz4PfPKI7BM04XrjixLO+u29eEt59WidK
gNLuPHHLT6lAFisNyXo1AThPIDfeIhLPcsQA3eOgJQ+8m66aHyTEfsQ2QX5z8IfJiZnabnncze1w
Ru0cVIkBUlwGwAxKLcsjKxTRFOrpjj+PhDxcGuprUqI+b30SZUohKFRizM+vqs6FYGdqg4L6IMB1
ZZLhGXB6ZHJU5WJqa2bRc8hXASge1XV7KExt//7zJ/W88AYuHhWQmxSrquihjlHWDUpH+jZCJnaB
ZtTzWt1ZxCi8sl1KG+bNB7spwoV6/MovRC9U+2DIh8J6WLmZxBIHX7aAmsl1FDjap2aPvaKUhQUg
z9oz5Ank3BJ0WZVfqR43kOQHwByhqVX+4ab3981try2RREPq8fz+QsTgFhdUlSvvwpuVDDZxjVXo
uahQU+B+iyn2d1o9IJ/l1phfRlp8vq8EV9P6Iq1w0FPVTyiClru89G6k7fNnBJDUjrg3qd6Tyjb6
rsd61ZqenKbCagr+ruaIVJsVxYPofrpvEwq86GEe7kPoPVaphwHIdszEdiejk1g/dZNWP2jxruqj
18HppxIFUJupbRhXx82xqPGxtawMi7zskLovRjTf6PWxwUsxnuhuAUymPfiMdxU7RedkI1I8hLEV
VZpJvpvaCoSo3GSNe/+WDeBGRIyMLm0h4/E9PpGcFj9N/VzbiXJyDg1nPoc1ImvKrxKjTfqcK14l
0ehuEVgZYkVZmr1vTCvVpB95NJgYE/GFaHGKpWj/gc5BH5Ft8kELVzVkW/l8Y/yjh8bxrfAMue+c
8uUIC1abWxNDMkXWs7rYaiMk8l11eCQvu6vyVMuZm6UvkD+zgY0k1zg/Dqnni92c4fLuRXfEEr+Z
SQNZgazWDWDGmcDKlafcdM5JP9kHpQ/fQfmAjmhauXAzNZdDfKiqY/2gExv+EbpAHuFqperory8p
kTrsj0lxMDsGTYf+t2jYwoCj3wVcH+w/jX/AG5hE8rgCsxPH5JNaeva+n0Pn22ToiUW+aD0V/Bxu
tn7TPvu8bmAwkYMqMZQMaNy5YoFV1b4YoypSwCVg3FwNQwuyMOvp2V5kPvTmZUcp4cU9LENiAyVe
YWm8uulHzsMGFNUtjvknFR4ULcZhqY8nZrFIec/vBD1YrFOsMkBDlmr6XPGQycm5Df7TvOaColiU
skSnfBIQhjKZWYGyZ2iMn1SE7+Zz4X8r/VDFKxWIMgIfJRUmOWeJ4cXk8xlVHiAcUlIxhIt9N3YN
v3TAeCZRCnA914M2xClWmpBwi9Bp5fL4mWvp7VAuR4i7hLPk7RhsLIOMnMmXm7tneLSkfVWe3VLt
B94g0zsAQ8dMAXeZifDuk79mlT9KGnZ4qG6z1QUlTBbt6TBNIZiB1cS/bvL9GTaUPYiJPzuMGYwM
Sm3KSCcnBqZjuuNwnzXGa+eCybh0tMIYR0nI1Y3tZvnXtBFoe2gRaGxXq2AoiTFTUjhC2VO6bve5
+fD3w00rU0oCauj253ZS7/5latBCXJVEzRz+M1U2/lVaeBsenkwPQDUDx1lrD33UJeOyJEpEuA2U
ASfgMH89fYx6XDbk29y/TC3es02KkTsqSCUOsHVk+DIxxldTU2Cq2fWfrPEDXiSV2Yb+ZfsUyCRa
X99zU40FsIwpjqC27sSEIzX2XXSn+6U5hGRESOlMKw/wfM2tG5tCnLvM4IGpeNFZrzU8G6vRTYx7
C/6pWKdvrzMsiPPNNSiSZaQ5ng6chCWMaI+3yOp7WnsmAsxvH97NqEZCjdtHB/ZjjWa5brZG8Dlu
d/Rz/rAMvq2A+GMb9Lwuc/8q9bvrNJb2Rxyz+A0VHQOFk9+gcmMwq2MY8I4qyYwbNRlx1/L6adb4
nF3yHkqCzM7Cyum8cmizCHWRzZci8pSyj0kpmd0Zw/AyLeE86LTkJp3DIjUMY7a7gSQm4RZhKA1p
4nY1YdtHI1fHCLc1O2xtGxaYmkA+AeC4F1WfcOpVd8OlSGedh8/QllCPA2U62ALhA/+WYRM7cMV1
6fSing05EnWub9a16Q/mWN2rhybidN5Hl6YF93Xop5f1McI9740wNcZGES/akcStbysFfINHow0A
k/WSqGHuY7V6xn2SAcXnuMiM7kVvX/yHVYLczNzDfHr/t6VtbYQiMODxZEqy87Iy9D8FOLeCcs4Z
927D1Gq5JxEnja1jOGxH4V4FFEovJubn8GxGtcEKS8h1QUemLTwiyWjBATSDjFSNyQOcLy07H8Jl
8UHrmS8FN9odIJxlRw/V/9cNUOL78CHPeJQQY+Nv831cy47XugnoYgighNkz2mAzb+gJwDtH/lJU
050CaIs/IDcW3dW/MJvd4D039HcaGjDQB7I8rtRMuhmogXso8k3sfm/ANUBoCkt5WmHcDCzPKD6W
Q3LkEH5cioEOpdqtkNQ6dwLIJTuKS6w54Ozh/Lhinn7mdATXh6KT6q64vYapHwvjcAqaRE5F7LFX
arP9opUlLKoLXquYlzJQA0LtaxLNaXxnPzqW4BbQ6hShVLBWrsDNJkDv5UzY6DYqivmRe5rrwcRM
/22ZbKa1UAfaJltxKUKoP7Qiu4IjXsao0F4A8wG1ZtNdZg+3FDBGoCzSigbhiMEEW3sgJNUXj/sq
XGLC6WPaTfbrrDTIL5ktV9YjmkZmsqXoVsgypW0YoCE6lvIJSw/Vaj6TtFYCDOAECw1iDZoZDngP
hgCByB2cInzYHYA678RwfytHK4aFBhsCsUFBkhj0nGptDWOkpOgdkqc5zXzsVBOQBkzp9eGTDDKG
jrccbeZmpNWi9aSgrhKA31rrvujE4ctYGtUdXmgivImz4N0cnlFwkQXlSqHrB0GyaxoQmKOodoaK
zOkoV2d21DT2LhvUlvq37D7Eq/NCX/x26TWgFdmDlhUVms487YQqoZ9fXBU72S0LD5LNQpfo9dcc
sc3Wm+C+UyIp2Ml13GOmFSQn6P99DTSL/VLaEL2rXyO9jyJGkNNb+KUBn1b8frOs/MAN5GLU7B43
GMlerZh/0UUDNKhYyr+UqG/3cvqvwdhuw85pQeCZyNrEWjtLqOo1Fy2wjMIUGY5sI/p+UCS2CDHi
z3EpgBQTCDYx1QfcXXJX17J/8H3jre3hR1eDBO86FVzrJtJXxkNz31My9KlL2eFeZ0bWuO8ZCyRq
BspijQuU3k8ICDXzrJOh4KJX7Z9b3nX7z4b3b+g4i5RQFg+nnMKy9Pg0VYi9gKlj8gDXiaj8K0mS
d+j+6NuBD9aaoHzWiZZEw9kwiDSZmkdr5W/VnrzEMW3ib3nhlYpKrh9YdeXZ1qQonCP/knMl6nsN
JXsMoNsQC72ywTRkVORdosakY/hoxJir6A4/6NjUvrbU6uI2JRnOq7qZL0vB4gR6aZL84LgFgrU4
FAMC6RFFRC8Hp5m3goHwLydayo6r/XDbk8aGgw4JCa3V+HxKZIkpuDyXFuwM+tLO9Qibvpoh8Jp4
GmH52FZOh3kPAidmkHon6Yedc8eHvqQiyguqMUSsaKw3sUwbKudVzREVvIdLJW4G7ukAyeEJnqY7
53HR9O2Zx244zCpVUdTP1U2zXKZyui0QQvwzejaJJ0TEO2REKW4QrbKbGLCdLLJSVdAIzo27wQ4I
ih6b60BoeOqVkvDwS+c+1jZhF8V7OAR7aroT4n/0cpnjbugP0UO9BDwJDTLCXGI9TJwnbmAqlCec
oY4qLOgfX1Uooo47ByyngDkVsZx2Ig3ESVxASqAmAHGzuaev6iZjYQJiPj3NAmmm0ASWEyOYeF81
fwWWSJG3MAKqdDS90dH03U60YQIhEjwSp32s3ppCtcM69GJr+bfJGfi2gqmhahiQOTbkNNgvIXmS
EXME50kjBCVto2kXv0jjVlSx8kzqQ2XF9uQ1jhbqJdrYMgE/T5TOfSkN8W3u8gMg7HiqerSAEl1k
QNUHMiOM5pDDCDB6XD+rsew1EhGXC5QHdgMltFbGskCx45vMqW9Y6QP0IrqOtm77sjCYcLx3dhTk
D+HVfuzYGshw3I1GgM4aT1GdNOL9FmJ6vajROno2bFSU7N+smd7pUqQ1ipYFch6fuYDAUQWfNF6x
ibRc6JmLKQGNWn+JdIWhmReXsmAXBgCw/wIdNrJHdTpUTu7gP/VrzK6exSLeoG0W3TmVg2dNBNuT
gtSeRCiD9fjEWHAiRKhm0O2DszMYIbEdTeRF6bpPVnqEGvPxAqnENvU25njt7ThVxT1c+PKIUY+0
rq4RUSQnx22F3M2WYMnEQfB6a/1yegLkFNcmd3vfMwoWEGgNIC5ZeHI4m6soXVXtf+R0ZMBLPH0Z
Inu5ZlUi8MIpejFk/ISq3paLytmOkekEtKV06eCJkSZTha2v7CLVpGOWGfjFMn0mOGkLrL0vov8F
Pg/5IK7lea/EWmo+hr0mAjWBQ0yte1MaLhGwFQjl6sgPCc1090wQfoiU+q0nAUaonyG9co7Ru+vE
VEqXlIk7vW3phFUNbXsgCE9slc7ocgj4phIz4TEViJyXpdPCQIqgzTBqr8E5BR99AxisM+wl1Z+0
cWHFgkDlXPjFz3VDb07i97yYAqf4q9eQkwOm1ZTsza2hB+/5QnCKjoJWqdMXVMSANogclSQ9N6ZQ
Amlq9tvVtSlVPhgQHqN7jdvgGcu+U81CnUNmuOHel2kFRWBhi6bJP1vNJtntW5CevrP8GfBuPRr+
E6AOz1EHJbQeTJCn8F63Ybpj35QQWmulN8ssLs7++KQ4LEArXbYZuuUJwXmFKVSCjwjtMm9gVp6H
bf/nH3S3pGrAgwHNBHIw2n86inagT0+1esj33h+3LqE/9bZ1VcCOfprud0Rm+FElN44HaZy2V9y4
xbm5+GOIzYL/M8BA4f7JXXj3cEeMgFWVARWz4lSP4FYUkENEDeyCoZHJy3KTSYZCz1esW7/hls6R
bBiIieLIVou9hv5TGH+KYfRo9KKXXVUepLirsMlOgOyTi/IEZI4AClruHV830YXoif7z2jvy3FiZ
bs6MyRqySnAWFA8z1sSZvzOpMGiYhMnECAlz3fAiIUaOfiLMjZV7AmkCpUSL1VKABe/DQo2e6CMS
+Y440F4G9yZ6+7lUAddA53Xbbidxwy6VpYaRxPxvkmJ1CQ+y+w8T9CsoxyvdwHnUqnXySG5xU+db
Pyg8pb1Z9OmS003Rk6Yk8rv8M3gLsXRYEFhk6RJuKUpqBeezF04fOeJrbB44BvF/h0CmGpL206m1
0WInIpQUIwAwKIvUJqSVB6zaCF1lp12pPN/yeS9SsgXSIp0vqWmTvAcLvPaqyDJO2f0dfr6soQJn
p7Xj8IG6atB7D8ezaSlHrCHmrvCDGs8cncLGnTwifxhO14VZxZIuSIaVMLzjiWQbbGqxBL4sxedy
br4fgvJ19+d3gtQmWumXVMeOrW0IaPgMgNflw/ABYt+xCrskWxoYxmfyFtjlOuW4t+ItqbfSsfNy
58WtJTx+vSb9uqeiZWwkAZss484nAPqkYwtf1KT/2iENw8/W45oXutzdRb1B0TRkR8+9rNi+u2AP
M9cTGIIHPv5E6RdghbwYZMZvOmKeG2BlDSU1xINuJ8kP4mxlP0PC8ha+isGC3zrBSRLl2n/tIhQc
hnt8kIt2JT45X9odhgfnGLX09XaypYc2KZL9Al6CFSCJE4oaHhELhlxrAfqqwubzwi0enZWe7VZ5
KWF4wqHv14aPdO+Wva617w+NssGuDNqH1lEValanQ9ul35glx3kQ+IXQMYcSvcDUf8mj2fBkGiCl
Q/dWfjbUTi+OZ67x5BDyhuT1UaMjVtEZFtSXJTYT3A3azFjbPeWAbvbXLXMZLjUbIPuAeUGLUSUs
nwDYOhJD3BeF91j6cQqxaylDtttIY5EBzNc84+lp7oc0EL4unMdYUUnNdMLp0AYF+bIq8umd0Vc5
kBpyPrbQywQE9R6L8t+9Y2GkRrl1gZUgfkn3/3p9is068PC4LQFKNByI4auRjeJksYaWpHh3rQbf
2Qk37yTAYdoKu69p7EBt1ncmJ4wGtNK+w27+FMY/7OX1vJysmn6xZCprqMhY4p/+B6YWTVG7IAco
qh7ND6sDUCiCgoPRKw0//VlbfMaAP8Dw/Jh/9SmaZ6wImLgkiXfqDhbU7do3ZKf8Et/kC9VoEoE2
P5R9QAz3clX23skR1Hra3LVYcoNDjGytu5FmKK1EOGfXGprDwWwBXNnheiJP1MgaOSkmwVmaHM/2
pg+Xju/w4XL9hJe4IzU+/kPDgK5ML5i1ykQiuxhP3+hijTdeBK7m/Fq720ErUu0wejX24nx5aDWi
VZ1QqksJ8ZmmS426Z+0Nr5kzuNiIgPUisXnDcKHHvMjLKa4NgtFM4kKOQNoDYUpqNbG0rGRBiadP
XyEJbNt53WZzcrXOpgtQPaCH+J2Dm5JV6shXnj8o+IyvEfn3oUaCJxtnz9kjPau/0exhMtaa9p8s
tS5XAx0ak9IWui8YJRAW1+l1KXiQNSpA7+su/glvesgQpDdvmyjNI6TOZOH52w5WU7qVdN3y1gyA
vvASAc/U+ar3JdHNDNkacswxLsTmSFQ4GCPOTze/9odLndW9MsoVRFF4cxbuQbBYmedIKGY3i7h0
qL/q6hjqYUllAgx3GV7u0XOhZvDYCLYiYl01Z2VdqMbcUvKZBcLCFckEpPG9YrU6GMGQJURN0cq7
13kLO+Pix08pk3tb5UfShaQys2YxU61/4Au8XIptPHp1btoY14unQUyO16Sd0DLIZ05Fq2b9Uask
su3RExliWtGgV0r091pF3OYrVVx4cyaT0KH79kRgme7lkYnWI0uCRCObNpaxOThTg+YyjtXq3klT
8YLQfpeDoG0jINXFR7QDhK00fQIM13Aga4cW0Cb0glOYsHufCTTrweRcxE58H6T4AlmsE4w8Gzvf
pHZQ7QnZLWPGW0syd5j3P1gDNBVHOkwMOTeFl/ZaxLy6CsAONF1jlcsch+72hyqXRKEeWTBBCgFo
Q7+8JIra2zumLyj4VC12b0Wftzprq6cZan9fNrNiClHF4Aj6NCg40qumPl0/O6A2MqwMp44y8m3u
H0Gy4Kt4wIw28nodyMc4zNcTd+lHOispHaa94oan+AAFSudBE/stQBrZny33E3jwvX00QUhHZU/U
vGkU4ekRB8L0EmdA0Nr9tmof1B0tWgBbq7DtUADh2ToZaNI37FmT71xuA/9dZKlRKjjY8Hm9z4UR
SmN7scXMMn7lBfBSdgWX3yKyWN6hHNjcbIS4g7LDVGIUnIPKyXlgf8gUwQan5igRUkDQwRT8Gd01
iYtCLBgv+Ur8adSSvfht0T/TSAHjstaNw0CEVLoizmGw+TfHqDE2CVqi1Yd7j72ZAoYg8+00BECX
poB0Je70dxqrHPpNFgNqdL10PX7+Sx59oFjayYkXpX/K/LUXlnwHyVwtgyvDEC/7TO4D4531zztE
bRya1h6YbEFYTFvMIYEUup9jGJJV5z0vBOmXDFJWmfGpZFH4HgeOsHz9ZvOeO8nP7jC8RipX+jd9
64cGv5wkaESJfLSZ000L4EEcQ3ifya5Vvhs6i7aSW70i+Xkfs6cWmKb8DPOIELllXZzipSWZz/Vc
J4j1Kllwnw6OMLEfEETbuuY9Bkhpw4iVFtmnk9jLSXNbRFDpPiJ1Gy2x/TvDUxpP3XSEt5a/x0Bn
ghtOdB0DLiRAoS7DWOsh14BoHt8NOY5tBFJIRBqlWxtbdlCZDTW+NCtr0CcabTH7ESQRtHgY8O7e
c0ET8KEfFFh7+FlKK08hUOpJXkV/J2LW0u7BBsLfW/2BlkwqLqP35qRKQwzKC5tmZgpAUJV4lPdV
es31hOzHXnWm63vgbzS9/9Ph7j/Jw2NB2IDpVmE6Sm1l9ttJEDPXzDnjfkLF0TE13uMoGT0CQG95
YeAk35LuzDkHfMeV9JCLf0oWn3pFZgfLK94/toajV1vpMarDyUoXY/1E/fWiYd1Jido7G0UVWpQx
Q3GfHmzlG1Oyppb39UOJ/upIMcQsk8+dp7m659Vfyub/6m52FXFz3M7PSdBXPoD9ATTU+dd45185
IzFHtAnewL91a2LAq6P2hMh/TcylPbxBn05DxMDgX1ZJfhZl7ZFhjUCs5hp4SUS8gWhUDMv/IpB7
yIZ7m54jOfiCQiAFpQVQGQ64b78wvRtJbGPr4sk3dN8Lwg2wuV2ffNfwzBY4vrzU1FZJmP5zQUwD
St/69ljx3x4hunupdUWUZyH8JRHfQM1XcuUD+8t1Mn4ZfhoiTHEp1LYS6shgDMRvyhHgHziVm8HN
1X+gxDgE5TQXsCKhKzht71wdeYui3hXzefOjKrEinlyUtpeec9mFaOqc8PMGqnHhsotiWBMirAV8
Lva9p/6zTOC9t2HPyIo+iZ7aLRJYQmHdzGcVZQH1s8cSoejuRZ0aIZgUchSBGwvnJjcSc4UtF9j1
84HonLYlIkBVYKVWHIp5qluXO7F1bnoHmmFdrZ2VaOLJcZMqN5Qt/8SkUanV9hMjAIz9dV7DsQzN
9S95Ac4KeIrgJtAhnTdO/oESfP60T9r8JmjKtOlWlK2gocHmFqtRWSfV3/I6GkG1mOi5UcV71nqA
e+UuRuDaQMJwlfatuNvcYwGLYx1XEqlluCkOHkZ76Kl+VPE3xiqPgUHQtLNo9gLn+/T2h/zUVkHq
sHeIMuqQZI+XthGLfdAbbMgE4YPRpBII1AfuEfTBoz7Oh3+ZENEsCA3k7KABCsZdkYOUYWM9778D
Opg9a9hm51ouKt9iMZlsIpluc0KZMqPj5ukeX+oPrqRcUa+HaYC9i9uGdqTMVwQBjxzb9S1rwT53
XAyumem1myz/FOsa5fjUYppExGU/usLWLpCnrceAYDyBkO9OyDeE/3ITYyf6Qt6Hq7GI7qFxnmMz
Kp/rbhAUZMir5RVGnCPHVcC2i9CS0nSoijckBaeRoEPceOUxib2r9vqInWCEtituXHGnEIBt35wJ
wkVBOofO42LUXblmJ9BQ6fSiEkaTJpLCgIAPuAcZk1ujTCm06v1IAE+IQ9UF1Aioeknv0wSgylox
dimQv/b85wQKK/zHEAHI4lAg+IqFu28wgsP3yyglOWas1/sJDRAb55jQLpKWAvQgYPqGCvaOIi/m
E0gQkAmFckfy+QD17TOYaBkfexv7uvW5FodwZKJnAbFOQ2weHdamJRUdeuUBL4JC741oWE3wihDf
Vf3Fv1cNIDOFyDm5yPrSrmmWTFvyt3Zy66j2trdQUC21h2bHyiYXhNKVx58w9IkNmSkd9uErx72C
6PemP2I/xbOp69+olqhUirRAdHGxH1MV0dLzUUMbQ9QMiWbDJtQKwjhzMXXluPMtPL4HNPEAMcH9
PjnWmUaBk/voaqqn15WDvlmBlvtgEaXyrlheCYRv5M2s8B6hOojPgpDdlrQnuGBVWrRBDNbWoBsK
T32zCbzUysJvbLgre9XwG64fcJ67fM55vdxtHwESsacOCcZya28lL8b0vxr9L5UO1/XNin+v8Fyc
o3wlfGbZGLHSTNUvMP+grdMfTkNX85l/kUhYGXsO/TtdlkggnKmXdIV4LxHz2UNMF7tUguPamlOG
AuJruK6Ol3NkyA6bn4oYmPxASkE4XNb1nWPwr2ZcFxfthIJw0RiMU2ualdcSYMtsq5YTAFpt8vTo
ci6RdqXngY0TX2pf7/5hewhGxxg1wFsPIZlErcwoq4bdgmtZXNz8ldeF6ljJQT6TszyuK6q/hKU/
HXeYdOx7xbAJNplNF94sCyueiW6gPEukZXF/Zr9SJO6S7fbFzYcV+6Tf3XfXBkL1/WSDh2yllX63
CnMtCwYv/EvfWugczr65byqN1WFdgzg0rtPRWWkoY+Orbymw+a93/OuheNCj1XjyqENu6WzPkfke
qfEa058GQrbsxRKMncgpv7w3qs2VuhPKYzKHrnfqs8y7rki1Sgw5wYgzCJ5eS8EFo7TPimY/QKTI
2/uz3csw6osiW28ZBVvH1sry9TqooA+AaOqXtKY9zqlX2cxT1ozTmP8lbEvz/n1Y/LqGyS9ei2wt
RWTTVqKJkt/jbkOsG+L2lvDKEABTS/RCZiWUdOR19rK+/DgWlu0ncPr+CqVyCMtb/gdApXK6fLol
HqtoD47IdOHK8ioLfpBH+uGIcm3yAD+4bUWkNwd9DVY0/Q6EnB5rVTSXOzQ47s42DKHGpSozzROH
Cyswo+1pG2YD5XBUV2Zx9E5Z9oQDpYu0r1vAUBt85YLyAJjQbhBhsfrtNcY5ZkjowivVKiK2yUQC
NKz5IgVx6AVyN3f9S0wdKQJ6UykD3savyUUHu4/anfLN6TT8vqRSe0R14PqVXF6zWxOgOqITI6dD
PY9O9SUPyd6hGK1bk4OQUlio39Pq2gG21Cdo5KjyBolok9UrM6u5noSh1mX1cgrVL2wZg+ybSJQB
S8a2tVBOD6YTCONEx8HDfM/7o2mRjO0fO7x/6XCkSATIAF8966GFlR4iUB6BZNIxXynLO9RN7x4R
dOHiiE8Aop96/6uuvVup3dLo5p8kjcMEFNSaRe3BhDoKDkplZFhECCZNHBYYtP0T+XUG0z1C3Nie
POc+wr23uUHgisRkSrViK9K1Hd5yYqbLPkVkjC0v/MQTXe+ZWk0ICHgY6Jr97aWdw53Y2gkPcjoO
dRVhOpbgEcNdIZcU2cOHUyuggyd+brUz71zpscCKg7fl3u5HiTNd2JrBQkxc6Ehfh74jRRYXuAv8
yJZwmx56RAI4+iWq3cR0ygzPCWx7py8Gn3zai4lLr392zUuQtFCr/F9rWYMwXtKY/CELcCxw2dRB
+a5iDjmuh9wf7bVRMXQ6QImEcg/a9DxpuZpwKcUdtp7+3SO61QcuSYE5qrxR8lVBz7pjVjDpn9mJ
f1tMIpp8tXojg3TnkRN3DuB8iciDeDsa1SYYJxQHLlJ/iSUqbIaVCa/pKbLilaB0vn3ljdfR4FXj
wbuERdRG5BTn5/9Yo8P4EttcrtS/OlvIbumMQ2TvAXVAjlssxhpbnmsTLXHT71EbgzMtBYXgW+b3
/y/xKL3pLod9QsZIFX1x7DP0rbuLdRRdsVSnSq4tWJ2upeQ+J+nSH/XWS1wmS7WCK/RD/7fQzzyW
E52WSkmpUBoZvc9m7xscM1kT6s/MPUxlLTDculQ4n8Sn8uVsLPmafFjatb9Lv6pBNwaz3dastL1X
mYC1g9bcaAgEPOBoO3cIcxQn0+Wi2BSxYtGocijmOY3onBJCX3DVGv2y7um5AE5p5SvGiv6i5UGM
qR1Yy/k8CTaOd0pDGdqvq0mB1VQYurqsf30mn8KuLMuA6zZsXpELPikoLi6BVS02MMrDQPQotP4H
Ehx7P1mN0fwR0NACb1PQLtFF0fGuWQanhSgO23pEjvWvgU1+AVFH2orZ8bqdb4zOszHmBqYiQiFt
dGAoxnceCebKMTlQ/yngabbp6oP+lCh+oUJ1sqlO6v4HbM1cCQYiQo/oB6BsvY3RABs7yGUwZodf
1Pp0WU/kIudME1Q7pnNQRYhsoAVLxhr4l3BLPfqEuDEWdiTgG5cpXoO6D9R3KI50cffGOjHOU4pk
WKpv9D+0kPhCnNn/aDY5cF8u3JhwWIG6pvxVVF4QrdlrGNb9RiK3vAI9Hki7Q0v54kmnBBxHwJvg
q7YXT0kE6DnP63ylTGNCsjnr2NgANVgp/579H6MpgrbfRJrLri0XCfxPAmQQhZ9RVYUYKlkNPT5p
gdb4ejA30/XsahANqgfNGt+XlYgmIupoIwWq0316lYhDoi+hydrjYlAsx6g9kQyCJTcCgdn5Sbiq
ZgCvpk3OOCbBdN4d6KtWLPI2BF1jXr5Dn7z098TqBwNF7pIbw9amG3Z8VTtvR1maLh30OT0Yhtrf
lBgZGpVZNhTHir1ove318PYu1KvVb3YLcQpCUqsn0lCqxJWaThyLCzvbKE8s2oxyU5PCdZiqhwAc
eAIQTqPCqK5wXfdyn/n7QdwROdhbfsPZRToh3OyArTB0qXcJ1ltPylRfIO1M6rHUQ2Z9JLMj9ziB
uatwNiNETWsHv6LyXHm2uJLCD3A1WsrSMZEvKqC2bjrDypo4Y+kwzaXdocuqYkepIKmNzlxKC0xF
NxH2uMjBrSjxNlXJIEzFby8mO48v9mSdTceJJ4bZVJY3P+LQx5gAOI5wtsYigGEvibMy2/jV3hOR
eDLmlYjQLTGhnxNRHRxrkEsXywYqR00QORwUHVXJ3acawuOgwOKBfYKvjoeoakHD/Dw+d4P9tZ7O
/wPdTwpk2v4asohBQUA67Ae16YFnH3rUDNcLLgc/7Cdah4j8wAmWerSeYhkHES0e0jBMSIYIB2FO
flQTtcO5XJb7X4QRlGSHP7XmQywr47j9UbTl5bCsFDhCIVh1pprhlz/vy942/GnC3a+0aLJRYtS3
7dn/On83KpHthSdfumKGJcsQCnRav7+tin6bqC02xl1hMKIHaWoZZjjqRWrL2uPv442t9YcgOU0k
KJDKWRcQn+eFVsmQkO8aIbm0fO2an/dLu36mFrd6JrcwhCwfDznT5XPBWR1o20gJf99ochGkUFqr
+0jlw3MMeJgRIY447sW/3OeQDoaNkRcc4kRXaej9+Tts7fe538NpORckIXswI/M4OzuhMWLVbdr9
Qtub5OlpjCnXXkzNtrS23XH/n1Fr6rP1esV/i6cpHQUEaQvpbd9r2EyDEtBG+ytAs0x78CLhe20X
YwWSRpUcOCSgLVbTNQkRm+42OA532svq/AfoQve4wyswQXwSwl5mJ7ilK+QL0nze5FazPtHMAIk+
mqx0cLECG3sQbs+zTq89NoswgPJbLupca4TNGpCuANppHO1D1ShEjaT6EBgUufwrOuxcPY6uDYTj
cG2docPPnmO3vXKmyasTSqYVhgMeE3fvWbR/5HVEtL6aHQOfJp9MXRMUku/n3vs4+toAF22WjjpY
M58Cf2bXQjnYDRMwrIiwA8FzHERRJXGZlhidbs+YSgxgq3GJmnkanwOIdGkA8+c6uiwXgSVP8FUy
2BcOnFT9AaYI2TPN8BSP8yJPb2CdjBrB9yQBnkkTF6tecLbeOAmtOLqFG9sb9sAbEU4L16G/46sv
CW9Wbv8SiHAjBcENIp2Q46w+Bwhl2WirvY57gb/+EuxH59xYjHmxH2RaQZxx64a0lcz7OK455A0l
tNiiR5G+7sEDenaIky88ozRJLHkfWZAnQkEewIN1rxYnD6pieBTXbtUSpDXhm/no61suRYKAQ65f
7F23pA11QnLp6tfh/Pr0drKHcOiBjKy8NbNaVd102TFJgU+XWosJO2pRw085NRVetNyyI7yJC/S3
RmXDif+74rOdLaZR+iyxA0Gv2QsSQl5ekez6lhgv3AIqYQEk0DcxUwvUHIMwjk6HgL1rmgNiHDzq
Q0o6Y6v8Xp5Zn3jFXlOHbQ5mQ6eLiOk7eKPDaPLrnT3x3ePfuivrMCvlCx5VMpFjV8bYXFs4r35s
ewSWc4LSaJNQFfB39TrL1wexM9VmpalDOW0kxpYbvOz5v0KodY3zd/h8+48BCsNN1MLj1AWyNqa9
U9QezJLeaFiaqmtuTtEaxzYXodEUxT4evVJwIWBi8tcVZJoowUGoWhJYDwyit4Wh6iibQIJJoNfU
pVH/EXRtV0dNfmBPJMZFwtKJ0c+2CvqoangQjIaHVTAhyR+29G+XJha529W3gi+p5URBI7p9LxHM
2gzknO9T/sYhyfl02autBHtYMiqSvKwhGPvv1ze7N73jcqNQ/kYOKzqtCubl1bycZ/xpJLoGhhmd
fYHntAsKvHgdwU1awioDm/ymRkY80HhQ67I8y9VB96xMAXTgyrh0lWDw/6p7S1g/uwFo7+9Vd+og
hMHKC2eOtCq/PQkaTErT3A9vjYu8GnfE2QmDQoHh852uaNOpRunty0OQPNR+6lCnR0qhehvQk82M
vFBHe8yNs9aL6ZwlWF09BP32mkmVyEmgtcsVa6M5W+2anKR6WTjwwdb4roYNKoEAneQmBjTy3g63
r6oGi0j5tCh8e+eCNWH7G6JM3g35Np/JCsD5XCgSwnCyheP1pLgN7jK6wXj1dc4z7L33lL0aeQiX
KLDowJ33tZQHAYYF2RyglH/JmrRNzBaN53TU9EN3htXymKJ1uRXrSkuW6Gf+MCFTHwDivhBY+Uuy
kqbVMKGwKBM0PFmyv6GkUJvWbnUXUmIw87hQSVdaahugEl4sNdcmOekn1GmXuLKgklvrj2ZciMLj
Sy4mAtyf2qTGasA6X/bkazRduZI+N+MPpiQhQBUtnu7fkev3GfL/jqaq1aCphWgbnSjG+qoo0RRk
AkGWIYU1pzCMIf34FbSc9PWyV9PjyAGeILrgWu5HthVD+rIQK7K47gYwaRFcJnahwnJM9oe8rUrY
5A0OHOCYxPpGe9Q2DTYYoUg64ar5vHvz2UxDz07XmTkwK4ccf1MWSzcXcq3mpkBjSWHtdhrxkePq
MHL94znC58ZEb5JER1lTH6PNfXpVv39YqDEKz2QLM73I5owOIH5Y5isnGxWH+WwFcggOM9Yh66yF
/n4TwoLCBgaeZZkWpbv662nyx69nr1K+Fty65KW35XQr2PP+DnQqam9CJLCKiwb5E2yBWvi6TlY+
Sp1S6BDGUC0e1C4Vyg7c42L7Yy8d29f1PJ1sEqoHXUtFwkGOQBWKYePr2lEtXylm6CSSnX4HC8g0
RtK3YGKjoaSDoViXG5CHjh3ZoOM8SzGWH2PQSGRRaOJWIcY/mqKzFqnDizAn1xQY7g/ebH+G1Fg3
FlxgL5F/xI7cR9xWBA7jLl8b6mPBfCXPm55xDjP6s9fUPPLQDnm+2yf7XuRq0wO/0R1lS7/WBrnA
1cS68wJHdRmsbJthDg990RY/FAvtgFOn2BlFrS9Ter0lOl9giTjfRYyE4+b0E5eaEjaVy8tz5p6i
m5qi9aCdmPpqal4lUa3Qw5r8buDdJISAeNPIvFIwjDR9hOFYV/CxK3WSMX/Ywx/9R7KFbGAjpHDZ
BtEcYAPsMUaJBMAHUUFvPvNCN2Ybh8JbIAY0/+3YaOqd1OzZuY2SqSwrGqCsw33ccOIcIiR5w/o2
SLgfqzbwLfb4WDmNopMPV6pYp2SlfapKe0f+QeSf3jmTplL/w+TK2+G+S0NSA19MqXMW8uRCPPu5
t2mBSeZw0nQUwgkkVI3BeRlwinLtbASlrovZUfS9n2yBKumj1L/iylYgXpyWlEYAHGEYERvnARBu
9K6S8x9u2wpqucxM5OqarlPxyVmZxq0bCGbcbpm8V+OiB0b+7vOnGTMjBTkhPrG6hYOM43yA3Qs0
wLar0coz9I3AYEv8h7M1YTa285GQXUgCFaFWH/AkT7Bk8t0LZyu3EWYzjdztAeVqz2dXs50z65e0
zpoQnEiyurTdiuDaaDZrmNrOSHRuQQV3h5ucdKhE34DpnFAZxnth5ihxEVgmdxrrU3NCHkZlUUUo
ByqOPr0robFscDQMH0EoN6Nin6nGKTyqc9WpA8fhM6g6BrG1947KjUkZHVh93RAfIdSgjjLn53lm
AwBozV3JGGg1Xd0dbuz9MwuPixpf7McMa7GN+yK8d76jsE9e1UVd16MoY0MCSpaV4cZhFJOy2bKe
cOaX5//UhP6YKOzndRH6wXoTwrDCQy6wk33glRf1JBevx9qUlMMAly6dEnhVrT7X6LGZaaQ4mrLL
egXps1eYYvyiSVi3xa1f3/agYIJZzg88qRk3Uk7NSSuQtyp9SWtcHXMYQAO3EqHKiLbgrwtttA0G
t7pT5taBXFEDajby0IueoaMmCinpYzaNE/62r6H9yCYiL9ZHdw2z/Z2FS5vbMxTH7Hq7dMYxwiMl
x6iest7qbGNXi7CPZ/qOD1dU/s906vpzRbq/dQ+A0jHOdIURqarZoFwjv/xgYQXV8Afyq8unB78T
W397dU6NZBMG/kXnnFjSk3tWbzICt7qUvfW7+2tYDz+S/45g/gdWclO6xE/YCkZ3SN70WLFbd5+0
cNMibHzO7AJsX3kI9lou1R55HZY5gv9jvg9QdoDDl94W6n7X5ize0UUFvVO1IX1lS4gqD7T1Xxdo
B3UYQ5kkAWw3I1ehxolkWYK4YzVmJJKligBWX3eBGHcPWMqW7vXAz3P1Xs/k2CA0n93Ic4i7g9PX
xq3gXNkupJNOOWZX0fao6Oyh54ClT07Xln7e1OjxeGBvqkUah8YS7HT7WUNNHZSznU/mUYKCI6Ug
KVkdA7J+wS2dZiffbz6RTUZex7RfFiF+/+OWaQIUDc/4D55pDl7coCVz00Aj4zwWV/NRL2vlo+nw
Mupu98cqMIMrmkOAgZMAKpZMfejL+GOHYZKonVENRQSWQ+aledlSm2GCFlteBMVLt4uueqz4YdWH
NujsjejCQC0q3bnRJgJldUYruosKoUk2eLrm7UJZ5KFa3dbRsZxFeLRuBjmjBDPL5JtJzwPcJVPd
899XrOsXI7JjhUi7LFOZ2jkcZEB1vUHitQhkj+sjZFzTKl4EMWOiF0r9jh6gBg4GirLC+n6BDHzL
14RzT/1oFa4Xg/BgsFqn1+iJtH+297tz+j0F6fN0JQcAcRzwicsKDpbFyAe1g9RrgUkev1eHnZjP
9i3G7yh8rDtBDc86zu8TXCUuVPeDeTBnL6yBcec/zp9bxaJ0N4DMkVapCTJ0hGF+e9LfHL31xk/F
r3X4Qc9Oepu0Joz/DFHaCOiDf0CBZeakW4DolT2gdYPhMtNS1dIYSViwcPxubLyqgM8OYhDKWOUP
vmVDm4rjYMUfQMysoPhZqai9x8o27sjgjkkYYEK9khwN7eyPlgPYCiNzFbCLJjZiIGDgonw/w/qJ
qBx/SzNkS/T5wryZVD2tNgAve6Du/HG9CxBjVb0NmKjiu7p2X5XQn0QXXqXMtfA50W8Y2ymOP2vF
8PKkJZHlj62cP4cro7xbIgg7Qo1HYIpWCznT/alVhABeW7aarDMyu7GP0ONL499HhXqX/INKC9Nd
TOf///Y8PCj3aqJuA74xT7vjHMbPEhln17bO2+YC9v2HoRNArQOVO542t0UwPjESLM3UMJJURbq1
UVla6j2z0p2Ok0Huij4j95bkQEcDEK+y7am0DxHm7diAN8u7oCO6XLKPin9GOqTV41kswGRBdUl6
FN/FGKqa0e5ftfrMb1wo+2zrai4PFcXtDTvnILaqHcb8sX8zNTYkusu2TGeGT/CElTK7CZZnjqWo
9uzcQhO6BfJfOw+fJ11ATY6+Mx1AA32uXWmwQZJoK6ipoMgThfZBHlw0EsmftlZxm1j1O9J+fJWe
Tkw87C6gn4JgCzWnFZUSbZTpl3OMqgyn5Z8VhrlaFOnZ42tdflNSOdKTH9I2LEbfw1jgKgC8SAId
F0nkvDVndLEYdUJGcHoKxv1TMVFQ4xwxHY4meYuYkqaKs+/mMyuVVUASLSmtaC4T1YKEeZBsSwzM
MwGyQMuLJ4iLihQ8Dp5o5qBulCxkR/hoM0xPdVJWetsnbeLoH+o38kfCizOFord845Fs9DwxIVwH
yiHPDYoDUxMci1x7wi2af9NAtJsFTDic6hmAlSsMUMTBNOaQKZHa/2cnzSaapc+G8L+St9GzBoeU
Y5KdrZw4ONdwwcqG1wmEiBm+ZvbkAdDNb6fddig2IT9OVCzz1bn9JNPiQjtKE0YOHRYa9z9zLMHR
v0NN7rvwS+QWcK1lcpbXJ7L8E7EjLdsScFWTSbgBh09z9G4TEusMFn1t9JyGDpgG5pSkjZc0U2L5
Dk8mi8PiUweWAHhORIjSrh9zW72r2FrbJkpTTLvvxkPdYUEpqwG9gtqaq3IMlR88dNBn45FHzUS6
sURMCDFOvB9EwqrNedhbf/a5npLK6zN+zAmBcn6cNdd9MeUez5yX4WhnMq3lXMBU01txBurhg9CJ
s8lt9m1/HirMLq/KPncYKP0ThhAbVqQiQrlQ6UzHx0WBaKfBzIK0F4swCPaS1MXoVPcPQy8qyJx+
jjM9MKWNyMY1jt8vSP9Hd2iDrIsBg5btOCSI6UPV5XsU20TGK8gYEoXnms+wxLljV1BxZgNUW5t/
SMw1rGrXRY7XU2ROegCnmAmpekcEjr6WRKyjhXxkWmTrbfSZk7ocWREz9SGbHGcKY1YFzb8xk+K0
xMXyMpe9UZt3A3SdniXETuPGgVfh5aGZRL3+En5nkb9pJm+DM8T0QCYueP5HnP9o9cfr6zgsTFnd
7WmD/C3oxe4xEozo5/MlY6DTEzuiFqAS6enuEymAwrAZLpK+LGH501f+AvEh07m84cUug1PHDmIM
BArDHmIEe8l/Xv7NNV5BSEt/6yly4aIsrs0XK3xTy8NeVl0QEHr0blqu1qi7mEMlOta1mHi9lRFv
YY0HH6hR3I0xNXmQfwuCfCCMXmYo5cTFOQhkyggSoj0dOYGEM4E+og1GsPlK4HCZ1U50l3tdGkxS
okYqLnSb9vlrC4WpkTfcO3whdUZQCop7nbDqpGJFfnHNA9kn0eaTLPvZ2TMdzG/To6fES0VvHVR2
9qeG8hv47Y7l3vqLgBJTqkIg7+LKyPlZ2YCWbQ80o6njSDV4Xq1K6+bDi86a9RMkQhfPU3gJgdqY
pSH1eqw1srf9TDhRctVrMlFU3p2Xapfhv2FCNdKKbLYbvSLHOgKAF6DVi+iCXfDjrDq8OQ+mz3as
6KQ4M24XVe+8tPpvPn2urNjL7sYveEc8s4ncDk4+lkRKklMSE4XwREu3NC63NC34lfLQTEI6iLZt
eFC1tM+u+OugpfCEpcImHauG15vlZPkX99AazFPDJZP0bSL+niMafF9FgT2XbepY3jCUvqCe+NIj
PPdyFwB63E7rEEzqBlr/RJrM0KObgTuDz1hkzyg7vks3g4kwH7zPhNTlti+MEeOtZLl/HCSUNEUE
2iy2w2rFLC+pDvUHOZBNHpl8xIBgEBGCD50gtFxHzejYkPDcM+Bzqg0OHhlOu/UgjF7H3K+Gh+7T
6oJWcyBAIXp4hTWFSqioBqzCHIrCWFaeuLrdfQ03kWSYYqkoukImug536xzRo5fR/A6db/6OGTGs
T/EA0b7VqZzJALxc5RpLjiAftduIaLLyBIlui/iu6kZf7YHNjFmzNHpu0pvgRM96i67G03XLo9iA
tY00c1XsIpbdW6qSxhzSYh9XxAX4CB/kQ+3y+wtFrWh57bOAK3HYYCQ+Sv0/8eq1gF3iKAuAd1ld
Wfkswf9JOk7Vb2JGleaBrbOYOqldct5VvGSxaoDVBPlfyLY6de7i+Yo66OK8T/AH0oai9ObfbzmU
8LO1OV7kgjYnT//Ks0USwfB/05C8wB6RhMrMC8vLtQ84Zsx+i6MiCf4Bd4WZ6x3I0IJKF0ozlQn+
VjmZHE98BGlXgkOwYftIHzsbZ4Zys1v+7tbrgzvqa/1i2mToXTwR/U8IJN1BOjA98EeMJxNBXMfC
kNyxp61jH+3Vt1kNEQesuDcOaiUEGdK+VcgwP7dsTYFbE5X2aeY0tpvDyyi5teWzI3fpv8YBqkKI
lo2ud2qnIu/v/jPEtPrMRolITez/uAtt+u2ikXGIy1Zwtgi3U7sSNK8S+12sopRD7iacEFdjDtbq
sC4aOB7AcCjwzn4gmcrst+Eh20TujIskV3MNVDOX+QECFrvgyNBt8dys29Wing+Jb9jILHCAzbq6
9D6H/32812Gzt8KT7BPzocFbhC7l9IWIQlKNByiB8vsBAFCA7FczFwM3TjgAa1uDg7FugYBbaGHx
mpEH7OsDj42tGO1nn4BA4e4tJafolI8KB3YjyEN55rxUnzkKYnLV4e2IMi/h992L3+Fe00GegmVy
hw6KzAjERHJmBJr+3s96PJalz7Ytq7rudD+Vuyg4scq0ncWezNaXoKCYso3uWenIYpslMgYuMhdl
eA4eyx3Mq8tA8sUY9QD/z1DU9u1VqiJWMUwP8qviii3k/YYW+S7NXg1oQIxB+uZDRJK7CvcY8lBD
eXVs2wWhIECUgZ/0wW7Kdt80DtGXyn2RfjdfkU0tQPx4koLJp8+Zw2qMwIGeseH1qjgo06UwYHh3
IjqwZ9aP+LD1iEpeV82+zEAdAS/je2k/esPVHKSY+k1YxgJpFBiIBqn4DzBD+AHaNU6R2Ba6gH8o
T5Ovv99ajVMgfJD3I0IFspIWrawsIIMOEuc/v28Mv3h8VxXqfKZoF8DNUHpG1XwqhYXltIu3Beiu
aTnVuVtWJfpiFS/5qtKm8yfoHDL6d2O2ZzyGa8c7rW3oalal0RBpy1Kc8OXhDlhIJ0U26UKljiKq
DcfZaldksTEIlr+x7PwahoOwU+VlNGAsueIRkj4bFeCKt1fz4oxzl/jag0FsklKf+LZIx0cX5RjC
Vu2bgOQKamTzExJ3aDS4GTybZrZL77F/JVXk6ynBCHAnnNPEMrRV1Ho6eZAUyZFu0DtulMH3YazK
CQAQwnqbs/VsfsJaugFVOC9mRc/Zg7VXN/sUhY/SX667Ua23ZzASpjqRwv5zWpAjaT4x0aB3gBrz
Q0Vc8VgQKKPJKrKHByQGqMMNGytjUrFgq2yf6idOrZ1xTR4G0+7CQZwwIfxA3IrB3VbS9D+HTuMr
PjaHVoKHGbiYJff1Fw01cYlHbbJOM+/mD20v6XLwLFpnWvrmkQWQ3zAlCWsupVfbOk8K/kkpApty
5DBtVd8DeBr6RY66D0wj/0+urvCaHS8eJ+bksAFI7SfjL8XBaQ5MEaHrveS3GfbfT7dLhzQ7l1j3
rbFMGXV+FZe9JM2iJDIzZfmYavvglDWQlQxBTg6rnOoV3JWDOIyO0IdcC9zaNkB0tJF+5E4QSSPI
Cy6BUbqieydtII9t7e+j9I6EUaSqrUTe3wxzj0ZGaE5kxEY3Lys1tJyhbTsIVpCbhXgU9rF2MOtV
2L8bn1tDf5xkuAPnmWpwW6HslTLF+mAnpk1YM79D4wwJ2yVH4QNRdDrMnIQpdMWZxWjQby+Htme8
DvypZps2JLCco5Kd5N6KkhDa5/fDSTH9R+6mbaiL4/bJwYoWsEJslMo02ElGM8X7dyQu55x0PUTp
pmcH3cpzcu50qfYkyLqNk9eIMbyLSvORW+0zspxpRM7mq8BCGZVgFKeK5KXUdwdOoJE5gq71iO8K
Ss4Ijr7VNhnV6LbMRYXl9oQ5g1LY0HZj5+FnGK1LQfivDydJxllxrse6mo++Ncu+RExbM4RxKjIB
Y0nrfnPh2x4kiFkilPRELWwdSrgCPPCyBcA0QUKD/2jvzLuS9JJqredSqWf/kARxW63C74xm/bNF
eL9k37jIBRzWZuFGW+sXi0GhaNMcnU4CX6pFJreDC56YtcHMsTWoBR3BqxEabLPEWJOc+GJoTGT3
iVAxb1KMeHIKR7G2wEtjk2MBBrlhnaeIx5m4O9P8XYvcYsO4dVbp4NwdTakXRf0q4G/RveRDZ42a
ImXetq/sXh0E/Qg4Q1+37crCaZFIY26oav8E7XKOWXimVdAwL8/a4Km353TRqOYNt2YElm1Kdgvq
v7nAQfOPLRwshYTSb38Z9Pt6+fIjmZP+esK1gecWNFRU1qbWCbrJH0ebvTxr3SNfTDQrMGOTWNMV
qvY6LkyL8GBsdKTJ+gxTQr36IeDvS3m6R/B+IK+ljNpvXiYQhxGWKBFXgt7vMtCw0Twj0vbmvr3e
5NQpqgXeu+dKdw3CylGFgB7mr5iDdpqVzcwf0vXCgXlspb5UgD0grKBiLoe4V3mihpIlzdHZU3dm
rNod4xKTDCQZpEvEmJdX1z30J7QqPdsxvjhXZTiKXOekI3gaF5Yofh6ZifMiY73qPchXQM8Ste36
7AU0MmRjsqEdK9f013YIGbwBfFHPiSgn8dgrlXWshlnFf8v39OHyM3sFSQG/9WUuMcczL/C2yYGm
J1scWVUB24SABAKuzj8NhlNz3Um7DZ4yiM4FLoAhkJXvYkOmo3qXAXlgefYPHubeueJCm+i/uzji
ZNmQFbuelrkTgmJaXZ1DsuNlNLUkQVn9yFcZQ1i2b7cZRn/M3nrcxq5pov23U8ak3hRDDFGosxHe
uZ0AHv1rs1TAJQ9a3k/p40PtAmdreE7qnLoH3MUR1rYJ+Vc1SkUWcivvYbWwLGappvCF1TDcFV+H
taT8QRD5Eew25X9xIuJEBDJvUxnpESj/OO2WxpRqApl3FrSx2hiLWhmgqVmE4dV6hV6pk6Ky01i2
l7I7PlmbwymmdPQ38puhDq8Uu/Micf+j+6txBNxqV/LRmqBCyAYfXGq6BkXjtJ8sFFQBO8ZYEcoQ
phhC74FDjceMh23USIn9fQVFSoAe168nSLc9Fk2ZbLgKpDV4bEeBMxjIryzKLBr/YA3z5vInkio9
CSb+YEZ6Z4i3kZIZHHtZEuh+iAkJ2X2LjGG7d8P//gf5Nywkwnmbj13chsaAFiZRGPii0iSz4Mxz
phMsLnun4oSaInja/nGCw3vMbbC/XZa1UospMiecZqGyXCbd6UTYBWi7dyxQqjx8x4hluwrZ5kJE
AdWv/1BQSrjZmVbgXpUvK41nwCqZThVn/jSzNMtIOqY7rB9HJxWZQSlStI2UpAx3rFdeadCmePMa
+XudpyiBOmbH2fKnlPogsox5KWyf6m7oPk0T+ULvcf0lAaUZTuEgAwDC8ZWgkRRPvx8Hotexow1q
n69K+DFmFFaMtu9G9b/NYMgZ7JvNklnDO0SOdHStD939QyGq0+tvDLUwb7bY0O+382mSWWC9mT8O
Wj8ZawvLObs4MC/EgAAvJM2RhU8GKPJCTXPgAuk7ZQZ4tvEWNaa1KlZ+RW5vbWCU2rHz4dJDVRYA
/3Tf9Y2sKKvBwkoLL9HNGtMgbtAbVOflKrXSHAfDmzM29Up4IO2W06ZrIrQc+bQwa8xPpxlXPM/8
wLaaEDxnrfeou+VCNRpQ/4sGcqGx3RXQu/WrQPESREpZUW0Edk3PYtLWBDnmJcbukbfa5FkAHa6F
dIq3PA2MRtTScK+Dg4iPjfmro29L6xKtkT+uu9fC/pJHtEpFMVKwzxlNoMomeNH47I86m2KGMley
bToMOr657tOrvR/AUW8zb1hcixIG+0BoEGe26p+H+mFaWspJ9aLz8MGz1yuCOkYSe8UlyDmGMDhc
tqR6l9OiMlajiAdeUHCH/4zj9Xs0Ls+TNQmIdAwo5dx+aJ8xxuaVluc7jIArpBD1efcRHHtGatRY
BT6nC5KVdLW/hAknVoNGh+39syTMix5tIooGWOPpi4TEzJ/lAQOeN8Ttn6/DOtYpgQx2HJuoKq9T
O6JD1nuLkxuTTavemiUTuA628e7K9kdL7AI/kPkd9r4S+lKHxEv60peyZ5rBEx6nr5HGkV0J2/AP
tfXRaiznFz/YoTSFKZm7NUgF/G1cGqus8UIkUO9LOnozjH4BbRHiNwsmJrTkLyMIMLI87+GlGOTv
SteYYvuxnPjtTCEmaZ0GFEab40jt6fq4RdkYrTK+L0UGwdeycAGvRbuh2QGadySczH9OpmJUNSAy
y15J7atGYxnlquB3hOS/tm2uV+hshYNKkhz3HP3dL0uPRxs8glbwkB8MpVHNQYtCo0vmL6KD0QjF
vp99n0CTfB6Fr1bHP7kZO6UyLoM9GRZ/Arh9O1TAmjKoyQLl0086wLC8cOyGXY6QzCfRLqpY6cHe
gjzYWXSaF4yEaHW+x5CLnL1kzQSEWav1T1iE2fpP7ALfubL0FhzV8NVvcPR1hskFAMEkmDtS81Y2
bkQXYAUxk9/tPW0VU0MRq9COf4xbor7kwxwqIExB25feopEn82w2kk4kxrqA+u10+GnUri5yTo1u
ZVR9xDbx3sp4baGSgKEiJVngv6pxeCorK83CP4v7axV9REqoxq1ztH6hQFTeNllunxgKNr/LTX09
9au0psof7NNyLboE77s387ShhwGP071h4/Ltffp2R4jKOwUXdXl+EsXCG619weM+ian04V4lU5kl
ucBG20P70+7MSR77bZb7A2H57FHsdDsUlg70JXwv9KxqQ16vW6sRVUnMRQXdp5A6uFL6O+FQ1Rgo
4sCVvtHKXJKW6cUf3o00IdUDFO/lzjDB6ihyb16xvgmb69SMEFupJJA1yPZyVABONTTJY2s6c0Wi
Wdq3JIgPtL9eQJaYyFLBHtzgsn+VJIBxf4vE6wtEHrzZsEq8bxXu4q68EDPeeTEg10cRdplz/9ug
AZgkITafbvcVAmBHc1sRr9RLmPkUm/7XlH+/pdRdxSrmhWV81pH3MTVtnz7jfsMe2sIqsznyGnRf
qbthcKNRP4m1ZfpPWeUVbzfOa8Al5niEhJYdDzIjBDG+zLAe8MCsR11UCti9C48vqTnN6FnBRqYx
qcGkkqxj91L2F2Gxvl+rSI0NQVhRH1HeB59HBGMfALPDaOwjCqfatrHhLSz5ce7uXzx7HYJ5ik8+
dFVD/WHsJk90QXkcdeb+CeSrS6nWQ9Zi9aAGEur447xm/6SytX3UJw8zntHEZoOIih+6d/T/iPsR
7TwY3IK1ostWenzcSh86Kelcas5fc3hcaNXXCJFEDK3UbWfxRYQuNx+o8t25slIx72EcEsJMQ0fQ
ywRRHGKH6Ed+Ix/lMMbCG7W5eFdhwD8WnNIOJcY+f+KKzWzpT3I8OtcC6IXYpNOn9jFOYltStnVk
pY1N5HVHZm5tD11WW6vpI21u+C/mHWdpw9KO1INGGIANYl5GfO1hnizBSbJyA2abxEw2LW5Yb5N/
P5atl733oggsgCA524JWRfgJzlL/w86wDtMZS8FaqGdyD+dx5J0H//aavViNVVW3vfkp5BIOekXI
GC3C0ZwjsAbMXZQN3CugDc0CmXGpBSv9BuyYjlQIx8LORA9/O+AxhRu7P3cF0SvQkLS786GQsaL7
cBQmpXLXJwajxArc21GktJmxsFZS0jZT2cmqOTQtO1AdwXBEY7s5bW51qWtr2ENcxLvTjQLsWrCV
9mx+ExWTYaZylHkt7yvQvyfuAHgNHiSxc6Vq5eplmFKFdAmICOxjW/k0ZvB5dbsw5i88r+RKfVVo
W2penacfkYeRbf84VOPzXpMQlfC7st1cG9fsTs1hRQ9+AbvsJVAaY2ZXfJ9veAA4bTiNKowKDgSM
0N9SGL5cIvo2SLVN8NDNxyR47PxFHrA2rIiACv5J9huO2GM2pb/P5ZGTEVKKknqovSJ+hfp9cn5t
M9VxrQx8wftu97y74vTafJfJeNDfjf8DTMkS20xAj95nXmeMggv46zh32rw+FPVT35oDPeuzLzeJ
FrOTdrddU1gIud8J9ueBFPcs/B8dUVzTYHqU1sODfzy/nfcqU+JKLD2ei8Blgx+srbutFKSWO9T0
dYPp/+5UxTa44hhuEUJTH8Y+afl4ZtllHZvnP4QXV6RA9hrKTQ0ctmBbP6Bxxdt501p6+pFzBL/x
rDE88jC4SVg2aPZxl9lcVcmAHCRMFXNXNhwyGg/4FWRLCbeXv/Lznxw4uygojIV5fVqO3sMdx0gQ
Iy5CXx8XDipEy5Bv8JABiP8OTV8jMc1cWmYQlbg5KMjgmb0+4tDiTMcU2f7l+AylJVN0de30Dl6+
dbLoan0aqi0GtnonQW1qwgKI292YD4/08luoS27qRYunDK088pZ8OK1QrznyFiNAgSpPObIiJBQ3
9wL3hz5gV5+66X1XzQzd8M92Hy0DQXMBl9OJ5jV4g96tdZ5Bx0tknnhJLqrD//ejeJmvRz0mYDeA
6UkUgejtmdz/heoKEaeU/PO/m9iF6gCyj28GcCQacPP/Kz7WH0XDVQ+F3b3pjzyXGvRbzr04TTZ0
OfrlPzlVowH8zgOU91vptjPIVWQtL7GYz3SduQpx4UXVTgeuUd9zdE6fK0WPpYhXqWM9WS+zKr0P
HHzAMbT81Wmqg57A5ijNUFqxcsDGYU0XyLuOCNaPHyHfLSOCkV+P5MhpHjepPBswZ2yQG7usk2RI
T7obTl+FbEm7nguJGKvTz3eCa9bprh0e1aptZ1Q2ocYbrojFAYLC934nSFar4g+AZR/nKL1XjeQk
G7GvGeeFzl5ny7eXpf1kIn+ykwELAF0+MKJyb50ztTUIhddBF3e1tZ9yqm4VoP3pa5KQOrX6/H7f
zEej3FdAet5r8xTV5FakNcxWKAt3ypfX7fqGmiSSm2BU3LzgSu99fr5XsvzWjVLAK/+eRHB9lnqm
TtuhDw9+3LYngGT3f/DACMDlkRlAbszE3JvpaG/psnVNWmIs5xR7Wu8w2QEyttzl45P8tl7IZN1X
DI1VYN7tfGMmc6SdqOg9X1NcFfzRzumdOzdJPujqOkx7ry5n65myv3aB52QMOe/yOH8jSDRps/qa
5DZAAFn2k/q/cSNVjpzGmLm2xVy4C/T0GgcVTqxXyxSJB6PSZ0x3QFd7XqdRdlcu3zPmi7ck6G3a
Fp0alN1YA6s/cJ73qeXup0Rl+PN8lnNQDotz5IUOMpj+akIztGhwSEH/5hdpfaH5r0EMgiNce3mG
/ptsk9VYCvxf+Aaz4Avm33bGkbScPBn8NAKJtoQpWbg617vUqgiYGlDDxKNfZBWUtPj0xwBEn4hd
GahvEIm9L/tHWY2NGTv3hrAPxvPwWH/bTwO0JKuFiVsKNg33mI8MCMHQCpI9w7yyfwZ+3/U+HSDC
RXBcRvQuSk7owUjIHDHV00pIJkWUBTkC+Z79HzfxSjWzD0kx7ryuL5WoRun5ZYgCgStbIIYitb1s
VNn8RqzrtqWufkT8GyYkrM/UZ/bSfMFb5FBo21EYkZzihdmiR624KTj0eMMjxLYtTXCAK6Tqescd
R5eojDmZtjCmm6H4AkMuK3dLr4Pp/MYt5xQOWP/futWu+72P/an2yLbM+efNPkWyvnsuMMrLuELE
BHkcYecNi7U3HS701ua9/kbLhs0oVEuMLsBrgGeA5gSiCg/RDIQUxpP6JEr/piaTWQhrsgma6RJs
/aoQ+Pa9JLjCi++DxZQHItjEtHImakmdQJe6oNYPTJmigvHfKE5ggdeQ4O4w4yw7pJv+ap4jW9DL
tqfrcAJUkXmLvUZQL9VxN0H3lwF4ViQkJQutbIVGFfoT1n0UtmdzKD65OD9rDKJoOCaklBqrU0gB
ZiO+Brk4bwqZAEi7RXQ5lPKNOCrxVn2eyfsx2HfUygGsW1tATu4mf+jG2J5dYE68+keHdWj6pQzL
FrxAQ2rwyeMGHSCOoTetFJMw0Rudx20LQOiQGZC7VUdMU8qla+Q0aCMNeHFDl8NEVXGr420b1kWn
0WzFpZmehnvr53GhNrdBIPrK12nmtvGHLo/zwvX5sAi5FVAJxnS9+XbYRDqPdqKpsBeylV8xjcrm
TaqSxS1qa+ZnPyfQ2ZhWaz1OdhKpHUe98pfi50TzTW3X04OetoCWpiWtScvB/lUZspG4/D5NGJDH
1UGndgAam5ejROPxMQ7xdVmht9Dm03PZBM8LdYOXCs2Elmj5j3HsmKCyXU2xOMx3/28Olsg5ulOQ
LtX6QeKuabalceYzK4DpHXMlYehZS9c4oYlU5yH7+EZ9XHr1U1UdjVt1SqjK6UtIn+XUREr7O+1v
jSFL7mO7EyuRhyDozvk45d+D63wPFGVpzsi+UQWhKNz45sobCa5VBjCgiz+B5zJA2xXqR5z5QWl/
mqiU9tjetCA34Fl62zgpndbaHnYB52Nn6tgF8YZsA/2xHwi5MptnW9Qm4kBOzqxEQXPylVQ2+AWm
//MRZli0CZPomHDWONq9bKUk8FnMK7Cojn3vTtRglx8zEu1fl+c/243P+NaH9XsexjXsAXKc6H4L
07JWn8nEwbrgaKvKlBxmEI9MJWNY0ECbZgstgz6HRLXnZ+WtGJnqyro8/AqHUx8HkgRjf+fNIgMj
26PA7rwjLfDHRoJwqH360YI7yrtiz1wBoOC+RSj4aj8PR0HLoQE1hiWMQaVOLrwzXcbrIdj3nJBQ
7maGlm0vKZFO7eboO3lfliX3jEalIKWjTx1ItU3erbh5E+tUoQISwAZy2y/33GnXeTh+Xe9WugK3
zdAwDITSYsTIyRE+MtQgJdvCwGpOqBOOHi3254YT+7XWMO1sMoFfBG3cvwGWzk2RjXxyBO/0kWf/
nK1SVwKbrE2fc7iBlNR37o5Ph6P4Fgu6HIn2qc1tk4rNjngwxXx2QgQiap1OS+tXNeLoVGiZWlQg
u9BpWyZkNgLVXFDmE89o0JQhujmpbHwQL7ueRpNlxPb1+aF5ijxdTMdflep5CrAyD/SAtdtDVAEp
IdoWDUtP3/R+i2ooJod1ItgcnPon72ud+MiuZj7jonGHM5kjDA5tAYYZ6XcfHZialwfYCmbUfm45
VGj7KoHXV4Vyry77qHOiVcIv4GWqRr52UxmuEn5v3el+K6U12IDFW6WcMwVXBZPE0eFwYZ9Udp5R
3yXO8pge+AvJ4mEuOLcWLKa76SKpx2scat8U42olQIgj0XJ9Wn77+sfXLPlmHQ4s9+owDYl4v5r/
JbcGsPj1KWOnGrctQasQGDxEXxbITGvfmQ1OU5baCHLlMNZBYinD1vPrGUFfNLhkCaUnQUddEQxC
e6fIar8Ks3o9Tei/n+4BrfwyLjrMdNzTdTkl6y/hKeEXcmhroVPYqdgKlDW87xsNWuNcMOF3oICJ
ieS7aiFC/S767Oy2xMHk7YmPSYHPayLzd7yNM5jCwSeHt/ALUs/uwD707M2aqFxBI47s15QRFbvS
z8glG0k3vBLVEchcnNUFyKcojqVlHOpIRI7VrZYhNbmtXtinYNnGdXTSy9DiaU+LBlvhnxWlzuFg
IkJIKPqwaGngbVfJr4jLT1rPTa36n+mAIXv6a4rhm6HPVG34Hyl/YNfPc8I523lQ2lVUTin4ZELi
e9ze8Y11dpk+xydgNFJTt3zDQdonibd6D2Z9/3C1ygaShhiFAyBWDzNOZyZIEFjPMj/HGnC39RME
A0b6Avr5EKqbcXO4pGsvP5R0DKAQonU6hFWOgAuw9s7ch5zV6CpFLX2LDkqlDrcYLLFiQf6hLgM5
zO7Y+UEbQ+wdxfrRVI9GS6S3xZdqpGCcb5YISjBVGgBUegHO4Tmj4J4Wf29s/IAcqbti2+1yoDIT
mbmln4Lc0E6eQzjeJvVm/6rgrXQ86u3l7MkPjbvt6tW9ucv1484klwScDLNclBZnMQ+IYqu/1HB4
EgwHqC89YX8Qp6zWHSfJbe8q+joz6laJPwidohgUKipU/rRl2j2OFeBYIKWISWVJRV9TUQyR+jNJ
s1jYGY8XUVwL8W+OcOB/GKcjJ1joKaLBhemKVQ1ATi+MFL+hTEgoxBDy+JbhgBML6c8fF/yDrvG3
ffp8Zh87dX1BVCx9E4bEdS/5T8EBS/Vj88QiHvyTHXb3xydLV94Fjt79wrpnG7RWJ2NAR8uxYd78
AE0+fRPM8vCHSaD8SFmGm+iCaLd8Dh9Gn5NUZ7DQFfpNWjXOeMYmXcp8VaENZ6tOOgdml38pwo3/
UmRv59q6OAbpe0T7xMMFU3Cx7yAIIBRwdGgmmbfMBw8SOUJTUMGzKvmpZrCD2FD/hyLgrwDuodVn
3SSDGTLJAEVBUtjlfLeODO829zjWFRvoCPs1QEZi+cV8MhFypFTjTRH5kXdnIDSF/IDhA3zrgki5
NLgupgBhnPdKfBFF4AhFDyX1awUWV8zyyVkpUmR0+62iAjLdekCrKWvXCf59JEqe//jH+fXlJJau
PST0/AnDWBPJeKkhSdVgpavlLrcy3AVo+l5n/ktc29kBgqnL31jCeNa197IJ0otUKO2T1aih/Kyu
5gmAWjUHVLSTKf3VVfEBHeyUasaHNXeabljufakXK8ertf5mWhXAEIN8I6KCU+weBR7BDa594I6L
L8v/3bZ1Vo/lypeZ9yGWyzhgp6pcPPSUfhIxOCx8rDInhzbwJ8qmiohmsncJWWHDrAamcQsHINPp
aCU+SL4o2v5ExPRmnGSZmFAvG98uLvJ8mp77Py6p81s0GJKMYTYGmxPgSuPHmmMoYQhI+Kg+pYBO
/JTQAEB8HKVT9YL/vhbRsRYI6/q5OJpW5l+fA5Vp7jG1qt5cjeHOiOP59kHxn0IVFyRJTZFTQTWx
pq2pmNvNH4nFa5F/oKT0Ol8k/9ZGYciM/rXFYr8awanrm+X1tpQ+hagdwicROlVQoTmpus7ZkOOP
5gF2m5GP5M+nIPvF3ewg3enIHD7JtIvAaLxr4m9wN2aFr9RPYsnZlrk5w0AlNJXo1m/t+fDS8h4q
XHw3j8euM1BOTWtLCZAsDngjFWKQU8//potxStTvaSIeKUxF3rmRsj13hdfsPVXVmCjH+JGJ8RHa
8GSoLuXu2dCF9zEwp+xtqJuM9NhR9W/mMLeUmLMEvxP38WFViaFndwc6fhfrgx64tXY3FwqHtQ6f
SI48CacriSQBtTatJQE0SVHrl1/JTtRlomcUQ9TZ3BjRCheeQ9HI7AZR+FUhxgsPHKbgc/EaV00O
bMCfg24weJJ0nHoTH9PtI3l/5GAKW8BLy48wHhIUD923vjpuX8JXO4xcR7LWB3FuZTrExXVVdugL
1pfBWW0ZXUTj6KYUyhgXkpPjKs1H3zfsbHToHYtW2mU/w754+NSn4CS+6YyVd7jgc4SHiYrMu2Ss
o2V02Fd2w3sXG87FTdYnRYoWffO835BvKMRZj0Ksphb3WLZuUbtmDKFI5F1ZhPW145xEIRoQOcfE
Bk1AwbL1v519wUT+hKC0Xd8z/p8Tnsy7eDo8YG2le2p5Cz0RJ1jNaZ2s7u6/NxW5MCPs4IBc+dob
TebdOb6XwPnJVNSnJSNj2/qgelXrmOUHu7YQx1ZnWSYOszrWoQJ8gDdlhQLRpcpj0LjqvM9/Jns3
akhxECdjSS549BS/0OlZGodv05P5DsTWzFVqBQJDrdc+kFiG1PcBopaqcW+JE5sJhnsa84jP6MPt
0DdjxykFGnZWcp3riP5jdx4THMnkSig8mRHZh78I+8JYlOADwm3nDkPpVBKBIyu11bsLJQrogXDp
ohf41b5ArCufdgr4nhR3QB2MMUdRZL3B6vrHgBV0MKCw+kxhFcKNO4Vc8DGLKrfAyVlML0ry9W3c
IUqFGnR33hG5PZnJF/8N1POXX6Ga74X+dX8x6ndggZ1MDNBkL2OKdklZOf16LLUG6X8KiEYcialR
axogSPQpH9Mx/SRPJZQyO+xrrLGN0wDc5HOJxB03exs/n2XybVuc4dLTyKqp+9DAkggQa1d2vUR+
u/2B11SmRxzMtSEjhI51CPWKKVqkIvhx3EIRzDOoLhLeR5m0tsNTePJ73rzrQPf+5g1rDki/68Ng
5rQoC8pffzCEhObLcbcA3OQUc5R1R8UiSSOUXaLvoSVuNj3Pfh/eFGDTJK9hUvuVaMuacBlIuW8i
NMr20EwDHz+ykB2Pk7MyiHpk9YKvrDxe3uRCIoPI+66Yq7UGqze1bkJyxfXTqHLftkL0qrqRUPy2
9CTSL2ikWlB/8aBRXoA7c6D9Q0PfKmtjbPQHUr0tkuI1B8j/ujjvcYfa9Bw8CHIl0dJ6Q/5hCRBe
R4ZjgcvvTi3wc79/fFAk6WSfZ0PdWa8M/VFhCSICf2etG4LBxHdx9clyFi7rFmv+VVmXC8yaHvC4
1I81e7jpaPWE1BIKBzratoJJMj3Qq7Rd81z/Y2MjplDCzk87JLuGd4k0M+rOypW7tuNxBcc+QoHT
iYQ5niCYw5FW+8WC1BQMDXDBZ/TGhVV4xIGx8V2+mvVvtzj1pOPhKS/LjEU7KDBQvQKGPRUc2nOs
ey+MA4p5hvCfY2LzI8yfJYrlngTKMFCwCY/4Ow7mEvvaPicYmGgaZnnRi9G5m8IRRTohnbkVSrmY
vmyISnA1JQKd8Oy7xEWqoJng5FDcpnQFqPkp8xYckiJOCeqMv3Cl6gLGdDGlzWU6+sTUmG58ae0P
2I+JXw5u+gMKF6wuPE1e7uQ/JhvqH0LH/sbtAxBwbhvNlHVilVOO4RAkWhVUGLJsXR5AIFUr69fr
vw1FwsbmJaFfjyDMaPITIgkae9WNg0C7hZLAC/WeunX0xC0m1+A3Q81GNKHjMqCvTK3c1CLwXmOL
yD4pp5/jJumFP4QZdjN2px4g9gJVYYFTVdw4aFvF30bz8+bwdVwJeoVbCQQbNY6QC4r1/WPyKRNa
jfQ2Gbx12Ae1TrgaJXhZYP9ZVrSKl5VxnZ0vVsSh8jB1MjQQ9auEU0afutmkwzHEBdUWcHpYp8Cf
i+xg193qC2YPxO4YwOgT6uemGbGge3FvieBaDmxz3cfUkppIGjlYbr7qQyfA/8DVnOXUZ0fV22qA
SyT472hi/X3vyZf46PYt8pFkhB1xUqi8b6sxCf3OLnuMwqUCtqDXtnFuhVwJxxtJdRu7tBzTUkEP
PZfQf9S6CSiUcIvb8xxx0o32ZxUCbQpfYQ4q+LE9CKwFXTFJmIBadGyEDdfMhxHJIy2FgfSj4owe
8JUN0a+HJdh4YZegZXgVHfAKQxECkWDsHCbfeDBzeTuVf5kgymzuQ5IqQH4MERFjBf87YUywNb5R
jyhCsCgbPIHrBSKdJp2vSFSJU/NSotaNCI7HCdqO85gPPlLfFIB9y9r2//vOmYc/DKtUFB0FqcIO
tAMH71tLNKt9ezUAKqewXndwOvF481el5VG6JdXqcQqxyFYSfaymeIP2f1icohf3oh/0LSwkH5Zg
q64uYCqXsPA7KgsNzzAV1lrlOQMXHZLC3Uc2h/eT8uu1AhI8oMf2xhB+tNBKGQS1Yq/vZHdQPkpQ
A180SlqYOhIfkpWDB5Xs92BGfcTVEkrVCuc3bL7wuBFKL3kbo1HStr972lCvKD+h1nccCONZlnWY
FNZL0Mm4fZmTpTs34Uu/JBK7phffHm+mWwIncXEmX5h5DrI2YsRUhW2SsdS/s3/uUrn1M/laqlc6
z5313VogPa2KRa3HAytnmmMMyEdaXcGt3obdiZHKbB+iPb9vElypVp9qutYaT3AGbbPO+wJSZZ6B
50Va28msW0f2jCurS16yz3OSDINFUHpO29kROLFyWKNo7V6drdPJ0kOrf2QC/HaIIXsrpJ03nut7
ODYzcrZRRkHMMOB3vQtwGYaCNmpf8QAmZDTtXfuZzDTPC7B5sHXkXjrcEgAkbFb712OxWYZkezzT
YmAUCepqPorkQ7V9W3YH0DUXwQuYynVQntLRkQ3yWcgLLvs4a0nALGZfyjk6NoDKS8NpeO6WjMd3
ESqE1NHEufJjXvmBF7vmVNHEddyJyq8SKQXIpxsQSoN0dXBJp3LHJOR6zZDiSlBk+vpQWKqlIpFc
wgHKn8nqm3/gfnKUWGXg+xc5MRKbKe7WqBP6HLdtVcKsS72z3HYMgr0jmDuw8fu3xVi9XBitPvMp
4UpvJTp/tects7UppBPx5abCRVwDmFOVi5K0tLAYq5SlggcJo4YC6IoQKWgOuxTNso2XxktJHZ5F
kWSG2+Ty59A7YmO0fZyKCzVXXEd3/lALJ8Y8m+jceU68AhIeTdQMYTjY93QLB2DDZ1n1Z2aDFaRD
FdEpLgfqdMJwca1vHdKXcsJHd3QW3l97FKIsotQ6Ph8CU/A0J6J2I5Wm9PUhUiBMfKCZCOYV3Uk1
CYYG9knDPjSCBHAyLcHY8HnLQVlBKJ+lEXpSqYhUAHwUcQ+8+VSf6esN9cqm3GeYZxB55zqBVEQC
bCm2h1IjtjqlTC7Aqp1u4lvg6ELZ7oHR0bPwaO2C1ANOEYsPT9hfEVEQayWjvbqqI2X9rf62KCVo
EqwEfzhDLoVnzmFf1jUQSCf/ZdqX9Mg28hASdkkENVy8KGKBkt2BFXEIpQd8gcto8bWthBty/SFv
Ff/UCwTKPVaS+PqrGO0uD7V1MtAWCny376XUrVDEUTO8scn0fKD830Se9bBjkkDkwV0QAbYJvAAJ
3bgF3aCNeYIKXXXlSZVEgCQO3JT9ImYHOzo6RSWGlilDgeg2xtIwCC6JMJ469mTQM+w2yNiOMzja
jMztMptvtfPq4a25oCYS2AuiFTz9cDFg3x1+VY8lVRI5jrIaX/S+GfoWD69OdUOw6tly5NHXF5m0
Fnd6FYl7cvpOqdLKvtOeRCADH1r9p80E5ZbVJSCz9u0n7mTd5iARMi0VFKSJTFf5ij5tNOhsIG9o
jx/YvNAb35agAoCXhi2RhHsTRvK6K6wuNkuf6WZVGlNB053xns5eLW76tVJjXo5LSs/QDe/X8x93
eTUMEw5IL1Q4/3KtsplOm5f9oCkpE0hlHqZtYI/MRc51hdKUYAnYwf5vDOg9/DOHifvbU/xLYKCQ
TFr/xLHEfxYKkWBb8JE4mIU4PGRHsD3KJEdN+gndcaE0wH7+JoNciSAc81QuPVn3RAC9HItc76ax
YoC43tlQf11f5b7hOnG5ij2Fw0UGPZ5yAbstx67QEjs0Cf1LLvdxjna9s2IPBCFofX6qZM+McgBg
OKBnds4tvehT0pX8KEwQozc1KYsu55KKg8AvauhCuLKQUFn4GxHEznfo5TUFQX9QMl9iz+Nh0hg9
uWaQ8ERmUxIaO1q3Zl9c0gbtmSvHzRjl4kROpjE973F8orpYerH32/YvlGHVqJ/m9NHCYIKaO/Z7
CHO0Tory1/u7MghOBfEoACTh/fZvdZDFsylFWjhKaUw1ZWBraSqTwjE3rIX9FCylT9FbKtM3A7n5
wUr/x1lDf2SYnLyhBI4oYQZED8+dvI3j18qaLfSQQH7k5BxdkDKUfAxarkQtkDKP6Gn5mV+4eBBm
Kg4pin6VyB300iuzU2sGOoa2zcPH92MLjFsJX+UWg6JIgspNR7Vo5YVoph4FsOMSOzNEFZ4TMFSE
1NxkpxsgZ4KRETru/dYaz+7CmIrFs0s6mpuEqvayTq+g+EspqKZTkLRk61r68TOr6LKmIOq7VT5S
dq3bhFBkjchgAl5v8e6wefR8M2SO7pRZIFCHkLrkBrTuskrnAhOU5i9fm/DLiI/MeBLY8jSKWeW5
tbvt55sU0WdJoDwnbfbP2NxJg3GRhjrtaey2aMThLzLd9BPdsen7TMJfrNqFmN123Ul7IYgcoRA6
l2bMFjm0gc/WC3zei9g+Fr9Kb1qqukYT9LPxdXuiz977QcuTCT5lXETQJd49FDEiLEK0cWM2Z+Vc
AoTIJO+tL2HzkrufQzvnbmkPfEDk4hE4zJHi2MzajCUegpdDaMliNbmDCjZi+loCw/08lIdUEFf7
9xmjeKYy+8Qfxq9yB47ZAjbcPuXM0wzS+Y8po7NG1iw/4rzLpE1ps6NTblsE60xm5Fz3x/IeD/9L
S65zH+STUqhFiTSbvJWkMK8unJgs8X+/9FSvnyxQO5bnZour9mi0Jy14fenM6h/3+w8/I6xXrjMO
l15rXOwL+BeN2cR2w4G9+D3zkR0sJSH2oYfsh2CYyBI32EkK3B0rA2z5OBtnnQLFXD1YJqF4gSSO
JPGKM5IsqDVwe56rtGw0Qo6aVZ3X21RbhxQQC8vQelwWjPogthsxoTHZs4u1nFFLPPbQEYU228eQ
vCala5JuwapMPAzXWEAVmUzmGza2KBLwiG7Ns52R6o6aS0eWDyB1U8K0MShwiuTKhRmc9WDl7bXd
rdNGSnUq7uIwbsZCWBB03/IjyuO1bhYhsbFgLoyivFWeZF7SQYg+BCPxHTpBGNozsglhl9cUWgQn
w+rxb6TWq/RNOf889HvY+dnvjW1YT32MZj5bTtpD54KHdxJoOr9/zhRsHmKVFzxBfzkIJ+WdKWaQ
c+1CgCtgt5u/8Gd+xE43rU89B6hnT9LDgSHjpaRl+KR+dgGw9mlcBkl+z4umTvZ7nK7KyBR4I+YU
3xCO7B6kMN5f6vtTLpnacYGwvsA+cHDAS8XlCsyGggJk7IT607a/Q3Suy+KhyYwfvgT5nH3MHaKO
4kGW3LOGkxVqHAocokECvP4RX5Ce1tCo0kdslru8XRfsAxLFM9ARMGhtSsg79mRwN477UGYLf7ix
m/2qHiALOaVgw+KT3OzQ+0gFCzlaCczLEsDy1bO70iSZpkgeHd2HojhvjHjfhazgE+1PGqCMLdb8
Y49XzZtdoofICPZrm8WV9oKeAJjKfJ2s9iMmWZziZQkA+5mjggS/CQMaJL1jWQ3THiCtmA8eduuU
bY67UdrocWtK+fiKf/QBX8QEnZE2Shn2jchP9ZzpNVihl+i0eh+EdKkQ0wCKnL+MV0ruRSTeoMyH
uAhKR/Qus3jR6HJsxQjwlPBcPj12pLqtrnuinDqpkTRrJIknUcEJtL33aTAkXFMfCF9PYBP3nCH9
5P++u7Fxls/jw/QceItwbEXdcGY3Qww4opT0dB8x3+z4iH++a2gM7yA8XTNDadE6gwS2jAsUu43e
SY/4n5lb+G/b98glpoajomnwE0T8OG2f4BNBCHio5NCNxaTvSNU/aZvYKAq5ISwJ7cHMa3tK9pkD
RMm/zgM+AWKfPyAVwL9JatZCeAJ00rLx1DJT1xPCtDc2a8CG6y+/sJTtwQUJbEBBgX6fpMebk6ZB
NFxP0OGSVjo0vnrgtZEzbBS5ku/CLPvCdpalsPUqNYDeMtBOsV4JVAOhD0hMeMq3ogtb16Qa5YhY
b8TYfPu7A1oxCXwKGFk7haC8lTITbDwXfOxj9E5GeDArQsonfz3Wf6IJFKRGWwFpzyE0E7HNGqaS
9d5LBIC65s7MhucVGm0TnmwafpWFIohL371bh4Ci8GfpXO5Q/3nCod7CyGfJmeZmFB73KkWPP7jT
0ytDIMtJTXArYdpnk9dcFm2xbkReX3+1yNrNtA97ROATOJSzUYy+fmJdVCWEfQ0s5S4rl+c9UWL6
qnU58dn07gYdCNWyYQoa9bunsrik3mP77D8snlYVQLV00XSG1t9ZWGKpga8SeNkkrpuFdOkY0GEf
SqXlUdP7wUEp/TaGKWylik9s4ipwbIv7/crB9UBjXrFlp5fo0KpvuChxirFbSUA1IqaH5VE9aVI9
Uftq/qh3UhwAahXewXoOLI7KSqD/WIvwBMQEbEETa5zir7kVddXbK1iwfLrX2qmpykgHgmZpuFum
oBZ+RUdKQftyl7iMwWeR8/dZ1bn8GwwK25Cz+FsyTtDBQi8B6j/Oli658nXHhUpT3x5TRaNu7hod
/6rB7f7+rXCrAxh4+SZjcG2knsr9Fv/V7sh4Bk+63yZOxb+5dzS8GN4Zr3TirjdkqwwIgUgGMJtW
qm2gU0RHdbx7bg8Qx7/masa0tvOUE3rRjBfmjgESoJi/FfrwA5D2NDoyTQY5PPbbnZHtFuQSmdl6
or1nrMNkWY+8JU3/wnHq18czaJaiXqdQjpm9ou59WQasEhQjc0a0Ol5Xhi+jTZRJs1JmIORFWMZL
PKrE/8yTQatwLiiLgODt8bxkAczLlg76IapSLTe2d/G3jn8KdkfqKZaDZ8RX7tYU9oVWkZye1zQP
NRME0OMjXM55IazB35mB0P9NcrfsY0sQJohbx6eGQODQ51yPSRvUFbgBn5U9aq8y0yzdbJjjoyvR
k23PCbxI8kE16XJu5c9ttxyRCn6by5ryIdFxIX+uJa17Wqx2iFdfilG5fvKJ7dwGkmL1z2l9I4kn
M9pamQDlwgo8u1G6xMVDvM3ehXV/QaUEJt37PQhYAmmylZXRimm1YrYsIEMWMyxAgTNGdrxDWrNc
Ynu0ppxZg673W3uHA7yReaGBG1xdpMlViIMrhPpd4tqJREtuHnwGb2fAQtxd5Hh0sVoMpsRwCCBa
7V4FGmOqieIYCsDVdkqL7761oxyUHTvV44Bu8nB480tfxcCkWV4kU26dZ42pPfPWjQH7YlOR5Y/7
kzgMcbMN3MoRtMqJa5fSWMrsWo8Zv0rmM+PNivQzWiempiqHdOx3zsPJnDsvRSgs3dg9RNzhcU0t
TszAvQxzAJef5oH4Nvci0KFx2/28d6fQitBA3wjbnrIBdzScrR0sPRZkDStKx+CnCMMDJy9EcmN0
F4qqtOx1/K9d9pYCB2VzGjusBpYzWOv3xNUrrUuncPHlKAAwRs4K6Wr1A8so0LjgD2m4Z4neSsdl
kBuKl9nSBphuOoR9ZEoUeGFsbGayiKlcyJZq/mPqoaux+3deFPo8ChVFmHJMo0+CIrzhR57tpkr/
X439BMw4ArrbIlcZaMqsR3iRpn4RKro8g0wwhXqE7hPxODjK9Ysi5nPpdvU4c/KDs2O90lEb8Xm+
e5LD1hTz1IPv6wBBNKujxZGZpeUPCDwlfASos4j9l3JzPsMBnA4TfST0/ZIoDy9seR386LJ5AW5F
lUQLDBWNHqvDH55WvOdtmhGMxHSVwCvjmGZ4BhdOGiEZFpXgZsj1R6l3fZU5rDSphfVDPJOukE2T
bYsCCuF71x5XSnR4VDpL5crivHgWXFWZv9eApDRPO2z7FLgfRpZgfp/fDhXQb/12nI6U+rgXBhxd
nO5L7h8k5oUYbBUVDZXDYtoURGzP1a1jS1CTHU6fN9NwgCP79/edPGUfAOH2qw6pLVDWAz/BCKiZ
Me8ETiF6T2kejzlg5hXQKssTMIEwUDbzNAgmsW/Egmiw47ktAhxeatup3B6AfzHpr8qV4U74zIPs
fjBkAKTcomx0pPG4ZXCEzKafOsOf7yBfcFB8htStBrHHREhp0shtRYtWchRHhGvx79lx+gGuhrYX
sMaGr23GthtM/hDNGLyt5ERDnLjNR0a+KWvVXnPIT4R2jr3VXXVmiEu7WAcEfqa+AeNw/zBD5hE+
zxWSm5cCe5E/36xAgAc2Gp/Qes/4UbFiOSXKfhakv19dDGTQisDvX8Qm1hlm8D4zwUrqkzwjpnq/
+luecLnMmQa5prmfDGuyCjt0s6L3XW1bfak5TAk919Oj5m72HyshZAaMrD406Pu8urpvT5QwhEJW
DvW0qawcUeFCY9m7eCAW7dswoKkQcu997VbMdRvgJ2gh9oVyFSzuXluQee3gM0vR1UDESIaDpF2G
Ed7k2nkCzG6FbgcrlnzxJZLgO32uzjAkgebinRDxlxtK7Hd0buJycQybKwtcCCwcMcdemoTbaD/b
r6KbPnWriVV2XL2aBS6fW3pdZmqzdoLVAxdluMZ+6ostZZWp1BF9ZuP9aUu1mnWsHM/EMSIxRwfi
zhW5FlqCgVZykhSQf3olw4kJmPgoENyInD+H923inhTcPTjq3UAAoyN3+VTVMdDL51jR2KSfSL6n
SLJss18yP4Y8cXZbHZ7J5noFc4ra/nk9J6MPXeZZrmv1ejSKKAABzCg8WrZaONyS5Oa6w/5gntsK
AyeqMQx9HekkuElxOjFSQsN7AS+3SH2a5u3am15KycfZOJJOs6I1uogsPyzTNUWO9buuHEUDcFhe
p5ChKdekA/5uRwc2CLtgc+5m8i9zmJYOhM5pRgW4AJHJ41VcUbQyn0Y9bWs5uYYDh9KOf/IgIYhp
DSdVomy3c0KFqbFev0Qgg8hPUk1t2V6g0OLY3hymizyGDeGldCLOIi/3NT+MuNDvAd83Qb/e58dr
q8A2rqf4434vUJUJSXElkYhMgssovFJNdKzcZRps+aGRp7O4UaXl11Y53koyU0pDghoIF7QkK6wa
eg0pstGEJJOGSuwBewOfB3OBf2nFdwevLJ5o14+77xzRhLjYUrD0yJfe3+pMsfmxHx7+f/nhQyxR
3Kb8+n50BAp477zFT79Y2BvvGZnuTTGbKAbgOqmCbvDY+DOUHf/k+G8e4PSOJ3uDeyWNJax+1Tc8
0lJagYgKCyvT9ft1TOZ5hwf30vG+wTY5MQDyTU7W2oJM1fj5bC+pWspU1+mGCdi/VfMrIqo8GxV7
EAS81VQODFAVsP/0Ydt0Wkl7PRXPaFSdDWT6rmEzCmPzCPrvmi7qUZXxCSmFo/xBpgNfhmVPfrX9
7/3Nm0LgTfWssVWhf12MnGVr95MMAwTL/OXbNXnNV5ZUtjXDfZ5MOpt1jru6GvfMBBUuEO/6cnjp
s7hByQW35OrlN6Q/4Y/Rp+jmqpoW2Z2Nw9WXgdQWt4RT4rp2XEXNfeyJpZqb/nLLUJXf6un2fAvP
MCDN3IwULZqjfndRCrgjVlBiTxbGILg2aAWm0DOCZg5iHezLbKXT7mISIg0oW67+OluzKI+/Sqra
NcrVWxXTgta9GIkuOcnP6lDxF9ezJzJemz7pF7ufkNfoC/O0owbx6H8NK/Kai5LmC9L7MysUOS1s
c5iEmVcsXSUWp5VdgvOUTZ+wIEQ9+ZYYfiZTB4tWzwD6ru0/ykmmuh5zZtUMxQgJ65F1O2X67a3Z
s+37gnvdg8V6F4Z9lFhQNp7BUDGofqzcZOReXiUyyWOGbxccdBvpYIwUxKOIi5RYNbVdKxZdKbMl
iI8UKK3QgF8G1ChxgEyGjusk0Tl0E0h0JypxkOdqHRZH2xircwhURAjZfQesL1WrhmJyu0UgkHb+
sBeVHnELtz49WujO+e2cysTqhJGyfGeUQhiKx6XI+coSJFijFkmfqvUjFnMeQ6ksnRJpn1Zn2eC4
0+x4avQ8/atxr28ptjESqtWKcMWtyB0KsjFCapAy754kUkmMXbMgA2pyAXdEQzRcyD/IiFcz7u/f
GocY9V6d6xvxJOlci1GKsvympjrB8grVgxkuCMM0Q8Q+0q58PoR5Cd9SfOev7IpYEwsnqIA9r7SJ
cvrKEcAfweOxK69nE8a8c6zwcCYX/3NFUVrDenFniW9Ky2Q+NGKx2n2rmRM8xZ66r76buaJFvaTS
1J7r2YXsx0BFNAVAzUN6qwEsrUwOxwkxrsxNn+RLB6wE6pgt2nJbCpFG8HlEqmPBoc0LJ0lXprlF
tyXUqBft0Hm1Nn+gbR6G6fjQhFabEcAkbDmNDlINm9qinUXjO2a3ima/emdu8AXnZn9TJwNH4ITl
glr8teYlujKBwf8l2i94YpF2F1VhbQBAfYWlA1a0IzixqUlVZR3OJSWKELi5NNM6w+tJ9q61TVQ2
F8mClfzp76BPIl6i7r1GYCAdTmq8IWqg8mIhLzLW3BgFKlmVRQhRVziGX8XWOEE/0PrfzRH1Ooex
Rs/Ak6ZoknuTFiBo8Yk0eJWbTx7jiHubjtcJJMrtu04spZt+sx+ZuHyT6kqQWhM7NKiNvk0Jic1T
CYl4Lu9rlEtNAbjCbyf7lGqeHBx+I5l9qSr5JJqwt1nvxc7eXo+Z+hZZi5MIT5kX70VIg5agJOgi
RJqwOt4SR4wMs5lJo56yMdqG9yP65A0FixclATihbhP6PxJ60+bJvRWmVv1r7uHk86M2ySIMGGAT
rsUS47C/LFt0vqFGrh4CTY6/K8ykHeHTBtNdkpzA3KN1lGNFNg6vsC0s9tXoJ8MKr4kvCyhNewZf
JigGqa2AEtRW7eansg6PREtAmsDYhzZnloBhigBuQzBwg4COj3KMR2C6dzIX/1f8b2dBOH/5oidq
a+yKlgIgghDwizPkolljivxvHqjZpAULCElMsh1W1+TSEewfsbMoTIkHSCApxJXazIJMA9GzEXx3
SmCtPdAsoQ5j4AvbxKn15XEi5Pa8mleOz75Oz+t0xP6Q5SF+ltQXdHYP+62xy688Fx2dKNGINywm
bRf/CeN3m0VODiN62pWQhW7gmMvQMu19mIVRVTSMGwQk1r/I2WVFm3tms6y2H9gF+RqmSKF68C1c
FpoSuyM2tqauLYSTM05YbrA2x4xX3gKYlBL9A38d3pOqM0PWoAxbWo2ZaL5GhPtNwOY2hlOoXuc4
xnyyBd7yLKKx2GEmp/vmi/hu6sLDFNWU/HGIB+OdoB61LXzsV1xiSmfxyRjjb7EKmGHXp66v/Xre
GKsor70lt/vqpDYN80e6yF7DAjAO6NdP+42+MU3bArPJJaOiRHydugKKKAYbz5zUE0oo+yjWslCh
Vig7Hn1lZpwFrHDCY5T+WAnO/uajDjxcuJqpbvxRQuteDDfuJ3caYgyq1xMx3W9OcHPOQnj1S1xw
APDOS9bm4vFceGIk6mijfZghLn58xu2LlINYOraUPNx4D4lZDFxzF/TvkO+PsKgJ55WGgryef8Vy
HZe9BCTC2P/PB/7w9K/77UI1v3B/RzlCkkGJYXlE8DbIex5mAnwdQ7eVehkkpGVwuk1mKXSXibnU
H4Ea5ZuHDW0VeexkcJRPQ/0Ks4lMIO6ynsHTxUOPed9sgU/1OM7GCH86HNK3F1FkY7+cT/Wg8l5O
o7JhTYz6qK5QOHpiG03GKWN/AgjvJuki7YC6Yc6i24RRmI0Dh1gHeiiaXFkc9dmOh58Zh4d2xwZH
/nFezQ+HDovms4PMJVn9XGg9phBC4pX+L3tEYtHQPU2Vr+TFCt+Dn0cTQNlfAdOkCH0UdNqRXQ0J
Vr4FLn+IHXCX2z8XRTfPS6cq5cUfowm++Ivp4OfFm6PvbG7fZ3qHbDqu/RfTuCzyUswrDJpow3X3
z3xiGElxbdShsUVu2VTEhXahBzXrYyQKvYt7EOQD6tWqMHreQo4E0cFQUeY6PoTGezujNInglb3I
w/WnjPcTZeFR5IImHJajM5Y1qNw89pXOQs0Ly8Ber9iLW0Ii1iPwfTNkQ4+m2iv28MvCEwi6C8Cz
JcL4K/4XsGfZtZysqf3+UcAhJWQY3C9PEWEyFvVggh93bHj6/dWi+EgFP2TYxQ0iWBLzEhWFGTWG
qM+ah+W0i37OdNx20q7dWgeFpgri+a6rPUZOf5dvOYG/z+xQklgmgttXms6qiO1RmGEBKKtdP/iI
W9UXA6IlvnTRV5TgOJrAtKzB7zLyOPYIXsjyNc1mcxapKCqvWnLZBGLyXMs6K5GELi5/iH9mNhVN
XXxeXpo0HcjVQ69txC8D3TxHZkpAuZrqPIGz2EbtJWS17IppAOIjetzCBgwXRkBuSZBtGfqKX5lA
jl5w37uFQfYnK807QwXdjiK0XEOqOhxe7k6v+FpLMnemho5g9a0XtSOWErBWlTA7Z/7eVGYS7PB+
3OYp7bvHcGm/ufnEgW0HvJhFmP2y1/dinIXdRv6HlGysya4pdX1bLuM5NV5JTSvqEepeRtUs/LTm
mDzB3OedGOVqTtXV5JzpIXgtP0GRXER8M8tWZmXXMxQ7ODQ/bUuoPYntFfUepq6QbuC5rzyInbBj
nr2xNzOPNJQ3TWBFLB4D/V44ULGsy/reU8+/WihdX81BvyHWMbBwldYfq3Z/9ceP+QnE9WGTVmHw
vwov31ha4s3sK92P3bSZ10QYPCNc7YNqTIiQUFcYXHM+wkCtlfIZQotqFnr87X+f8aVZC4T3FoXw
ai3No7jjN4Y+0JPNjvyyu1r3OJzvexOFnQ9tCuzZ+2lTHwlGkzm07sg473ErQ8q07MieEMSH4KOc
okGRjR9rpwpQGcP6iemqUIDE2UMStpvDTwBxMbYOPITRJ1qho7KSsbsP1vVPeeGtym8TORDvkR0y
iTFyZNzXlwUbTO8D8Cj+PDc2CwHFyEaXz1VjqtuZ4SMuRykrSTSv8NGlinAapd54yStLaHg3Vu/h
bAR7GGRc6IYExUNHCiD/AEn6sTNdDP9xHQzklUBII2hzcbnf4PUm3VqKl2521fD9QQ7iOS+1STGF
ZQeQXZJoDvnLZ/R4DLlAlgqC/8sbMudxI64Dz34RRNhN8BycWCXVdpJTuh+cclicumSAAePjvGLG
fh4qdwxXq3PdzdhTxMdH2+gfGprMs8nrzfXq7juhSs4eQ4pUWgsNTfBXrlPhqhVfEinTgzGeeLGv
FCD/PDfl93zF2338p0mD3b61RYqWxJV+ACdzVfvgFtzjK40hnpDp8pOMvhjyiSqpzew8z6mkVLC1
XcRbc9FGcgweN2BAJyuCL3Ce+smiygNWJ4eZslDWm1LjBmvIMnviBIMGSTccw0MVq90S2tdVBHJ8
2Napjrep4IFJWgdPHWL1H/8TxQU/9Al/gYh0IChwFjw/czuYU4hp3dJ3ZNoY8GaLj3Cp/DkzXNd5
7o3rCMJZHT452fscIM1Y4P/Z66DJGaM7jOIzrvNj+heCw1CM3wsJj/ThgmOPlGGD1yUJyjMJAkoj
KFQoGGKdzMm7Ykg7CBHZguf7j6RFA4t4Ney7O3ToCSQ+uI7cT6EASxKsB+pNa3h7U2pIIxJm5Bxi
7L0IgyhWKaWSQQLVex1ADzAqRBbqa2w0DeQPj4WmTQxsMfWSZaEMa11BsDuIeJasD+eGjO9a22Rs
q7Kfu1wJkaHC0rP0leE+
`pragma protect end_protected
