// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
i+v4ZhYjCPqb8Xwj+V40Yfip4MCYiJSE278AEphqrEJNZSSBLVEDdfIqhz9phuZq
6UuPBridxO8jhYI/tPI6DMBJIU15HB/wsC8wUovzkh1YmeUYqEFkqm1lcATq8hyC
yvlXM3FXHmLSjYab7G80/qVRnFCJoyjUurvpbYY14m4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15328)
fCn5W71i6dVkpIsQFBhGnA+PrDl4/3JFua/ecC/BTGBf9s2dQjjv6d4NAHPmsMEf
4vAgB1IeM6Gup+p7BJ6pJqqC4CaQEeNc7+piQI4BRGg+YV6JRblixS7h9R+lfw3t
SOz7tQbSOjUkoGks6t/w0WNaM1JGOiMbVMl8pixF/1+R5ip29VXCZjytYp2dyIjL
AB7THO6+5sacz98z/A9estTjmE4pz29y8ttII2K35aFW2wJEQraceRxw3GBDXM9j
jcwyf20V+WxBVmrLFkwBVn8KE9poGK1SWavu1DLMBr89v/HVo+VujmMvEu+Z5vS+
ZxJJX92V8kiIzYam3074kUcgnTN1E8D8QuQYNJUX1VQRoM/VQ0UvIbWz67WzdwDk
T9sf4mqkRIVydBHdhxcj3tE2wfUTpWl1Slrc2FWphZUUcm7O0HDDbTnDHPlqx91r
DhUBWFG+j1EXVKOr8neszcLUMluGHRy40xwUkB+JZC3nQebvjs1fZxNEm60zwohy
a80hKDxUY2YBODbHhe2tUfvwHdku0eEF4C1Wyum4KUcaLIM9PloWsyr2RIiUYtIJ
mcf9xwCcZHcZ/nenqfA8WfYYJycOjJWAuBGkHYvm3uSWHssD5mHqwdJnom8CxN2i
mU9MZIpOasNLKPn541zGddSgIntZ7v7nocB8rqZVnig/chTR37kg8h0ks8uQzOyA
xOn8PU1ql2dv0K2OXxV/0U1vbc0ildS8FU6sGHjFiZYW263OETypjxGVDqgXOo0C
uCf8kweMALyTo9aVmkvsyiPmUdbD2NPGoN4BzOMTSLvlFMYMPE8oVrFfamTd6BQr
TyoOkIiR72s4TpSGrXJdZQEDXUFcyf5ctuwbvRXQGeWFktEoAHk6H3x9vKVO4o2c
WW2qFLC1kgeFXiUfmkYWjWr3q6Lg2drcbBOAh6tP/sdvEtwmJV1RP26yEvNCmr6U
IN9s+yJJuff1A4/WZbnKz3aFQS2A2TKE4y02loe38hS5Ca4t3AdrdjUlwsn92C2f
ROLxPm/K4tA9+nJ0NcrqbDT/1ucWwMZGGjSEEZYgV6JVsLEMmYlGUO1RFlubbYBV
3RWUtEl9hjp7lXhV8vxeDe8tP2NzIqLoaWYucgEkR1zZ3dwqTSZ7vXhVwAXTGcTm
1ONyDwtAZF8BhwiqmBjFlh9AKZoBeOMHc1A/Kmdrf+gWteJpgEgtByHL8ST0knXI
4xBCAQU7DM4tQKAEC7LLdPAYttHTLF8oIii9Ic2wWYfubv+JvEdji0lgNR8UeHic
vwN/l1YUxsXWqNxbO8yBrG/3NfkLpU+AQ23qtu4lhICnvsjJ+mH3bDtdMvftiO1V
XGzS/qG7Mti8QCQtVEGWO/C3DuQ3SGtn4T3OdLYa1dWKfi9crp4CHL9CG1Sw0B9R
fk2nWyHkq3R1wtec7rDZRuDWIV4beqNOGr1vHo24KA0jFPKOPwI1wEq/Z4f+qhSw
7WpLPHAXnYQP9It8HvNj3wSONWs1iATkbRvcaw+SLOwOkHXIBBe4Tc9PAToBoYD0
8doYN7vMmYluuigKQoZRkJIjfPqh5J1PD1g5k//mI3M43+bzRYWiuaJrLBTkt63F
m0fiBLR+RD5CRcsifvNwMMLF62TouFj+Pb6F121jpySVWU66vPdKiO1Pf7HdjsJx
vkBqv8Lxq7JOboEdv7RnDqUEf45mte/gT0GQAojQ1EOcL5J8jMnRQKQiD2l7TeC0
/91FfykQI7hFt6KExb+ThmaDH/rdmGjmA2RX59GA3sa8MEkDRvbRm6aSp3JOrDMh
IQ95atjtaywoyV5URQb8f2v9s2M4pcIlnlPxopwjnwLkpPvaVpxY5vTg8AaqYbbq
gOwJYFWdvAbdeZq+va52/vBD2pVTSBflCzAjdzpFUAfGkKFb3I9zGI9aMwJ23CY3
KSx7uRHcI6BVWysANLYHEXaBl+Md2yBYpfqZ5iqAfRM6nL71GYHPiDkXHlR3ZBn9
SXtcrEYYrJJUh4OilwjIH5mJz8bfxWQQTLS7wpIkqkKKdsd0I7y13OJjdfgwzQYt
ftZuZkwTa0SUyoqMq4x0E7I7JC+L2p74UQA0e4Wxb/+MDQWHQJk5VOfOglA+lhU9
SFJ8ZpQ6SQ/KOZkgQfGpSaGCr3W3XM3fq7L3yKDkdzKOxOSAd98aXzLTrygwMbCB
1TvAB2oQIkY1yO4NfKxeA11fk7M/wicknMA0uWGyo3d1oYoOfe9L+CUCUv2OznJS
/kh2n3lIruN2i9/U9WrxNg7ptZuWMkrAlPLo4tbx8HB5wMoHgV8vsvGffqrGQC6S
KeOXYqfCjMLXqBtFIrhJ00lM8RDFRi9AkzK1kMpnxOiyhDtFAXfxGsTaviP80vOb
IvXzlRW1e3ubM2jdr0t08g//jTkCRqPQh0AU39NpSgbZiBM2eecEG0myi560pHOs
gMNehCCZGTBeCXkfGu09NLO0gZeN5JdPqfAzMZxlimvF5Z8ng4Q/oHieKTCkb2p3
saM698r3pYZm98TtkHOZgoiiiJTlsPbcir+mJOerDR3ZDHhIZUgNGQr7mlJrv7Qn
Ajxuqd7xyjj5kpNm2CcJJkYnMgHzM3MKfOzhxQgiNv+zkyY6I9oy6jxqYU5x+gtD
XDVQ9Egf9K+ZwHpdwxQdtVtWAUmPje3vfzSODc5rOnLuJ9zdXdID2joE8NbXVDsF
VU77JbXLCco7pdp4Sk6D9cohkfsYkyS6kQjeWzZfCVqB3LMpbSJT4xEX9HbK/iOp
zgqjMKVCHzusinqtt0gqUQ+ykl+tG/eEXNLNAivjh4fKRJOBFKsjAPPwmMITKYvm
p/czV8TkaV1h2o2/J55aHeO4LieK7dML5OeYlgHkvKjymVwwX6jgZNXsJDf7NEml
K5YEHcn3hisck3DHE22E5tcq+8G0xn6bOwo+RSw+kg3b0Z3mE2t2PSGQqP4WAuSB
+FMovaGa/u+NLpG/fpKYqkMff0g1RPHGCJFteJpwjxoIFlIbs/8XIwo1cjjxXEdF
Ss2JXtRl5CuF4A0SVkjFTvQFHQ+VC6pO0VzEoGdEWvjlttidO5Wb2TWEFmqyBt/p
03Hp4hfmtHLbPS9RyGYs8KKa5osZbh+Z/Sb/LsgUlvzdG9uY0xirCPfv2KU6E6uf
aacUCyCky3nZzFfImxRF4YFP6z01J2eUwHPqBTI6ewoNnP3mZIGrmGQG8JIIz8AV
qM/zomRoSmO4WnF2fPGI8aTlU7XRjwEeM8/cD0nXHZPNqTnEB0+ci3M0IRwaiEF3
EeX3mKZ9wE932EI5SroB9t7spT7lHe1jO9ZbwSHzRknU5bOXtls8Qz6RMrjh3sev
FsxjNJbvTQgFZ0W+ucIdvq9QtCX4TxRsB28YbGkrxZPt9KfdRWAn77aPPjvFSPgO
JKEKZwYy72AeO9o1WzGuIDVhtN+yl0U32/5wyW0Vrow3dzc1m/n3NR0x3enAPcu5
bSaU5L9CCpUGrEoYqpLgxwviCw2eCJoxTOR6brwuvHAnNoBzglDhI4Q7v5HoUQ2u
zjnydhS1nwWhiH8Z+f+8GPY4Zve9WzJQN/6e6xal6Qs5OM7B0strPGl+aLN0prPZ
bKSqe0iiZfkusB289Ge36E0kAs62VSJ9xMc213gZ4Ym5RcIdSJqQTyU/d+mdsFMe
LmdIBdyvf+6+F1jauGy66XaRaC43eu7UkcDe7sTIh3GX78ivqilKLYFmPCtSt+Kp
P9IKmCzpThbyqw9bY2Ojaof7EN6saZYdt2iLTcEejqTMY+2U6v3ftSecHMVTP43w
ghvnxuNtJvzR4hLe7S9kyU2+H3P+ehDqPJSmw99lRKw81G2H26K376I+0UnADIjm
aBNbegiKxhOz8K9K+md1bylsMtPaO3JI1yxs9rBvp+Hej89r0S53xkRy9FgSZ060
7Pp63eNJR3s6KfAtQbnvfIjIFfaxhr/RX1zCYgeKzrskodZVfaweDmuysFM8kfyK
iQGk50LE7a5wVQ67tQ6gupi+tDreg/NYyk6DPwhMh5556lzH7h56ZxdhBNyAE11N
/XvZAan6DALcOAq/Bz9CXsmifYilKdaU/LjbKv7u4fbDREYjqlk7nAHEeodpaV7P
vBktMiQoveEsF35KQ06HnuMaSSV7JP4pymHukyKoe0+EluPiGMrOlwn2gt12FxBS
K6PuitXWV+XxGmC7pjj+FQe0IPHOPeqLiKYEhiDDghtqea4KElph8QF9ftYvqZkQ
ONAlNykmQ+DH11XRXIiHTRe4pQfP+fdGDc8W/uaOLvl5ALzkOIQkqq2IikiWsRCY
iH9nurVSUT3db9m4R1j4AKL4jKPwrNLAMdOA7D5O6jzJT9r8MWaW2c9QTih8Esdo
E3nqMk1cti+dUCC1moFKo14hZ9fQ9tE/C9ezBxgoXuH3htqNTx4voLjshzalz0Ld
Yza7o0Hvu83gsn1/6ZqZ9pA6Ft08onMg4SYVAnJFES8LskJ/L5SzSEZmiL0vsPq9
QftQESkdM+P8O1cDiB7FOobvus8U5QxtEjxX1g4tUER43+SeC6f/l+3IBhUtJEt2
jH718Hb7605aXFFmtmWfpcRS+42WAOXZ/zR6Y+YEL0GyTCi9MyO07GqRWsqmh1EU
wWXvGOiG2MEuk+faTnICqz7xRIbf7NfINsmzJjBQOwHXRCTU14uiga3IZSilLMHd
PVkodMOvYcigpvWyZPwsYxu9qGCbKhOtPu01K9U/T9xd+y4wu7PlaqbqilvicqWo
0/Om+cS2LbMpswxlBh1ElLQHPOwoFjSOcxeN+TFucpHMrehTl6WvgwygVR6n3szd
zB5YLQF7ELnunDqYfbIw86VvA7R/LpFardqkWSmqmDaJvSOQiJuTYFADw25AiyRw
j/Bs3qUoh1FkEeZj+Bkm8bTSNMrHBnH8Vswk19qQoAY7I769+8/fuvNXR4+vCkSN
rc8gz+baLaSs29qegSupABbHFDcq2mplRmOCizk+9H9SsWQ9AvU2R7JNpXwqvjaT
8w+YSn4xPFVaeq1aLTAAFKYrSGmzDKiliFWp4+S14x/bL11EKMlYviITNsJbZzbS
JinMlTirEhHsiw1leCsnvOLnHnGQrS+4hXfLlzlLSYuefz5fbttJk6mWUOZbr/f3
gF9jRTPOJvV8UvPahkneUEZJC4b2gmwBlHDU6Y0kAGUM8t05MnYODPqryhtxtTix
5WHu8Im9YJnDiDslfWMugMCUs/2bOxq10HLpLhorZinOm6sREDGniZvsEgHCiGJM
Gb/5HMMIhk3EL7jfW4oUv6j98d8vsYfNxokMzvS0Q3jwT+yEMRu4XiiqQAPRCJsd
ROGtPlxbZmKYcU3hRGJJ0ntjH8Bb2SaRSsRypmISQc/18IJy+k7UKOztB6sy9uRG
MQ+8gx2h4tZWXDV1qgGPIu0mu3HkB3Cwc++SAbBASCfMowJLNv3vwubVkvNo0Twg
RCZebgm7DAQQxCNunQrs0U18aGUK0szKxInuKIWGzuIg6CqUq2fui1SgdR8Trknf
VV/yfVDTfkgMictmZi/WErhjTxzxhnjf+9VnLujNEW54wfoT2D03D57PZTLsm/Ro
0JjOGrvJ7Nu060Z563Vg8D34RW/Rl1NwjgPQhQtkrj8IP5VPWyH+xttj40lBZkFU
NzKtgj2NXDGrPzngv3naXufTP84ETFFof09Q6zFowN67zNtT53Dr82w8ZxcaphdS
3Sejxo7WQioNG2DY0s3uXN6Vq6ntYwOScb+saAdtBIuR9PtwaemLi2sCdeSrpcSy
JbH7CBSQGdV1W3m++fy+IAmghK3mx3ANzGyLAi74Bau1bfVmpGs36sGmwzxwARGQ
yep3MbvxKYjxgwN8NRIKqB8H2uwm3e6M5MFAzqtYCwQ31wJc0Z6U3vZqynZS1453
8MAo71jS6SS3Thtsn1HaMvLdMDpsw0bTBQs/4t97dJJOv6y5FeEPVwuhEIrj6FAA
FeEHIVOTVzq+mXfgszCWys/Ad5gRJwx2n9OzA5aYFsG7agbj3JI4HIajUzL1r4rm
aYE7WdNVo6Nxhs7GKRCizjQWZkLN1zqBPZMuC93TELFpRVoM9wyYnIWMBc9t6QwA
e/tzrLRHV+WVxmCNJJCXlxb298qwIg+g/a1u7l0g0ZgFjCXohmsNeq8YQ8oKiToq
NbgAzkz30QuA+xDYrfULIq7zJhdLmDCMv5sfS49C1buQ0Mf3+ET0RCeS6C+ES3zJ
thBabxilWdZdVoPgAB4OBxfuDemhrlBaOaL2TGrThQBST0jl9UsdM5KZLNS5zE4j
v+r+EwqPpqpe1YoG+K1StI4N7F8cAdcmD1amSx/twLybc/gltL+NTVaW7KQoz0cn
i3HHCM2O4Lne2R+AjnWOrz00CHjr006Sp6FfEz/l4uuwRV7NVrk3Db39ZkCokW/G
ilW5tRU3SCU+aez2lGBhZmbXEsMnTvWuuqVy6c2TScMVdIXe8/A32GCm43Zjk/Hl
3NHqc3khWCKXSnYsG/Ywscm2FjuQOXtFKgmtQi/Ydnj3qr20nTP8hNEG6vffZpqT
xdkHMsLrkal03OTAvpNgi7EWeQApNWBK+nv6PlywIppD6tRQ0E0owIRyjITOC58x
oqg/F5Q5EhNhaGqOqxCagk99DaNUycN9XOvO5hcppoRjmIHux3n3VvXDCN2jSwqe
EjNVsd33K590wtr8DojcCOCTCK38DqxB6lieKQi4nwIHmwEzQPWdZhymJ8PS2kNt
nlyPdC4/f7ZKCUwYeofiEUqxAgtkgyqXfx6h8AZlSA6/WYlRTzjV29OflD+E2fjN
Kys+sw14Jxic53MSC8MQ8ROMEB9zMyVG8bX/mQXShKDr/w8FxeM31skohwhoG4zs
y3JonmnXVzPJa5piCWhuKnDb6rmpvzqzINcnWpzKPYEgoAe5CDlE8Ng2LlyV/d+2
scSQ3JkbBVgVh53KinD05fjdXm49bqXGbG4RoLdClUG0tOwlovzMLfmGw8z9doyY
TqQ/3KBFqr9HKqaKhOsxxKNE1piyIU2tQZKCSDv/bWVbXDX7QrwqCBaNLYd2PncK
VDqUt28RZo5WP2Q5YkDg/jOPQN3xhM1mbdK1sG0bbNNZ9IWldAUzqRfXGaF1uB78
Mp8WsbPANsP2OXYAJKMEYnWLetqPbk4fgksaAshcpENmKFDLh+IgULe+lPbkZgJ8
pOJJ1C85eXcjjhKkrMRzExtdaP/OBMVt0Zyl05GCArP7txThGkrxnwol997/GgGb
T0fe+7f4Q44bMvZ0wZ6DqI7HjWmGfXvXf37L+PlkbsJY5vOvDmh+dB4kZ8SLD2jM
Q2ZEqpaiR68vawKvbYxA/Lc8ZWjeZSwB54q8OhhwBd2V7I6jCTectKlbQGFsyDc4
WIC9uUetlFcIHhtHkFktiGlaV15IVvo5PTn87h2oLI1LJEjT2Rk7cZ1TRRVFP0nI
ICKe1SPEpPmwCFe5idcjVP/XYtbKwDMzDm+Bu4O19+kBiRrT0DinjHjEVzvph7JC
78Z/Nb5FtEmCfkJ9fg0bwBZLaq9VALJbOQE13TcmaT7VyrB0c/fSRWhab+XYLbR7
V9G3HleB2FJkDhiEuzvuti7e5jILXx31qe5QfahayxtcAVCKugpI4Hq8Gw0Mxpfh
xryp5SH4ZQCuqoq57u2UvV4AYZpln/BIRuYVOJBZRfXZZSdJCQIe0kjkP/CoLkMJ
sgo9GnQGanHbS36ngbqcEloBCIWAbeiAffdTFAmQjw+vfI8csE9I7o0V/5rnmlkW
QxSSe6W48X8OSXBU5JEv+KJivXeuNyuVg91aMDWtGvlG4kI12Fle+WUGci3gepGO
QfLCKsIIJPrxj93JExv3AKHf17lzatrD/cb12Lo7PsL0sDG9i18cDxzcTH8GQMeR
se5Og0IAfpaiMoJE4JP6RuOnJlD3O5SRF89H3jvNJFzL6LaEq3pdTpFuJ324sSan
pe3x2snjnzNJxKTaMOGX1652jzH5m+VgfzFcHhcTqEwI0xPSznQny5e70tuAt5V9
T2GZWTqly+HNv9r2Z+7W2TqVs8/16I9y2TYeSRDZ79eUGfYveCRo/0gAXptmez76
EeukWTednajsJRvB6sDUV24CcsDZvrt65xkH2/vOZQfktHbcDNKMmAIFTc/RYxQl
LzVnxOPbep5TidCAhBQheaG5Ebo2rVMtzwxY+qiVb4vZm8hHR5H089ht17nBnCv5
sEcj/JRSCf18+t390GgpD6weBahyfGucyKQ5qLRX6Jhf4neNXdtjtZgVi9Cm1cPo
mJsw+NPz6AofcJdP2ogLD8y4Wou2gUnskC7EtRRzxL8ZRCBi4M6hWb1++DvkABhE
uBac9DDHnvyz7iPah9aE3bH2/SJh5VHzyNGXV1x0+8KihnsO2/lPTPwu/7E0MYX8
SPcbOJvwNfwZ6fFhbx8KNXVVab0IdqGyfrvSRi2fkbd+IFLMb2/+hrrHjF5tdJa5
DrYz/pchaaX92iRxkg7QtDjJlnX/ZTFRgkXa4YTHzaJEhtXeMLRIMpSAMn+GUQx3
vTa4vXgMBsZVVhN+cn+TBpNRXmbPCThbR5e8xUid2rzbSMoDJybXeCyOpfHr/oCX
R0EnbR4o6qP+nEkmX7bfgjeNhqmpbXsPHzFzoRaYCBMdScF5OwJrmnuuEKjWiG8F
eSP7GMRJva3gqoR9Yu/HncW3UnwmwOWsJOtpdhBJd6vGRQHTZvjh12A0N8th9zUI
NW0FabLjol3j0i4oC6aNzfCGZknpE8+Qq68xUWKuQ0e4Yut283C6WR6QQjnSwsE0
ofuzTzBw87iKarABqx+fgaxrQ9IkgQvsnnwsnk8HFvzs4MqAHbwOnKw+JtGj03mK
4NHLABfxdQlN1irPR1xFMyv9ghcCrT42xH+1Pyuwy8o1FCPjJvRufSJDUNsu3XiZ
XkuG0vUET7sNzVg3nGWe7p830edo5kC63qOO68iwbRmtB82Ky6PT8WM/f7BE2kEj
83fG3kHfReclbGx9XTjg+FFe2NLejNma+oAq4va+3RnI3FboHAfAHtehZtFgaDFt
+6jsh+ABYTNe52oVz+SixGJg325dGetBzy+6RJzkk4ukkS64/kXgHLpVe98Na/D6
NE8qRfJEvkkjZ+OL6+hef9nPfe1zcaBfwAUgRDpKziPEPEetAZ3PqPWAWXrpNi7A
mZCOIqKxRK6fGs/XTiDUlRrMg73r5Ekg2mw/WKzDOeGuJ6/6f0gaYwr1fSrUOTCm
VgdZeR8my6QS4/8qlk/iOlLzL73b98MuJ2BzM6nHKRs22NNCfeetthYxkiBOB/DE
Wyd2QWEBq3vvYUbx+bnQSGYrxkZpXDa3i3xlx6YXoF/89yoj+aZjc1HUVJdAPkFY
UTzIqjRNHyNXfdBhMzl//P/tIh/AL6oYMyPbvo3dGdaVeKPA2L+js3tac7PrMXBL
0HcMlyrwDk6yAva4xkNrMp9umOQ5V7YWkz5s3RaoO968ycyf0LX+AFkuuESHIxhp
elrlkyzi6qDnGFuf58V1OFLdAkFEyCGVaBQBnovllcAh54PHY4nMXbRq0Eck5G/t
cLwGDsFs4TkKkUtBJAxC1SZ1PV23mCFKJWzo2I6AWlS+YKq1NpqGu7CNc6v6k4Sy
/kdT3L+HA8w+bTWNf5AaspM/Gf0tht7WWiF+omFH+E3ngUrWVr9IdQlQO/y+ckDO
At1NQuafQ2Gb+x5n1gWyZE/Cc8z9WlhhvwUrMuO0M9wNdTzu6LQ6VSG/PyJRZMJz
Ri/I30d9X5E7OlUsdt8GQ25bVuM/zBUpnGyIRKegE5w9Qh75wTo0FeeuhJsnQx9C
cs5pA/1Ah40JR5oGdZn0X3CFQir8zahgBuA7VdYx3ijDGWgq9wFp1hSx2wnGF/Yz
Kfi2YhgtOXht3SeZ6/8LubColdYlzpXLu9ArqDofxw2iO15sX1yb8kG+TgxWuc5R
mTXp3qzFY1kcwMh/QfUEZPPxgm0El13HnRBSuEkc68hMOmKgN/mH31ctoQr2umCu
YuJNS+lsV0GZ9hITi8Lxb22TRkA6ZG3ZGiE7HvOU7I40QQyOw9zIAsuN2adbFgmN
8CDK9PL0cGIEjd5VxMbIR5zuJIs4YvvaQv+ZEI19Y+z3xSpkA3MYRWe6/ZsOapPQ
DOaijREcYZz7rU9wVefI6Ux/tJT36YbOM9cGHjazAjUOrTCzieTC3M4lGOnE0w/2
b+bIt90YRvMdpo9SDZ1ZiZaCSn7EMj2ZP5PmM9amkB/BN3juluh67yPied7/740m
8JUcUpMz0mpfBuMX7zsGXazCEpb6RrsR9G/UZs5XF2f8HVzSNDSTw8TMCQhf/ptx
1yavZ4i+xT1HFSml6LhzlixKdA4Xr6YmszJ1YvogSBRYsOBpyNxtraICZutni9Y9
q59p3BbTIjynRUuFa8r8Vt68j63GzTu9jsSAxuDexwXenuXFPtM0IeGODqsj+etP
3klyRp81T+9/29Dn4kYW8PelU9FxTBcr609ZV07P9W0aC9U2sm4OX0WL+cXHPfbM
aryY/DVYd6plsYL9oYOCj65Ni1soFYu85BMOD7RbSuaa4ACryB+Ip03jTS1UEA47
GjPZf83Ea9Avs/Ee+vWw8qLm4eA21k1GafslSI59a/zQ+nsSDAJhMPhtIfA1XhTn
ZgTwmC1WN3LhuJa4AfTaL56eNs3SD2ErHAeQcm5CSrxuMXKMIOv893d1sQx8VNKz
xTQH2rLOh84mC+lAXFlC/tpkdGl3i52+Qwik1nAzibSnABPSh/tvHOgvGc4PiuWo
p3npLOrdUhVQbKahVdnlYNnJnu6mA5mFpNcoAenONOQeS6irVkd8YeN35TiQw+sP
SAPe9qsfQ+4k9gatrLefDj59FfTNSy9ooFxW2GlRSqxV2E3fACL6kvowTqyf4TLU
yznl7rTwdQC50WHSNlpm2OsZOlIzYcc/zvhAi2DsQrWdBIog19dI3T5VZX2yt4LJ
YT8PEHnt3bvKsnIbP/Mcjs146mawkgCuNsjRFFQP5NkVzpVqjRhx4xwBuvDUS4QZ
BCgWo4cAiWiYQNoEcnEXf+JCLCyYM7ftCuczdHyLwoTJEWt9Sc7DZGfqWgoCql+7
upb32r5BkoV6zAbDwCRe+h6npsO06eXRU64Jc677b3qE3UEnKpZPCEzmMelVDVam
AlhQBdPkhRH3tKMGgT67tW+b+hQGwNRWyOc1rER8n7oMXzHJ40xXCPDGFLqsrQeH
R/SmKBzHo3LNUkCL3dIOclovBs1PXDpLcsrR/5t5XtckcvKzSP+0E/X1ao16pkAO
GcDKz1r+hGzfv6q589NHaaF3towmYMH7XEd8CGzJQM85R4QygGhwpmkDAFikysVk
Bgm/ru1OiYg2RWMd5vvK2lww9JRBTbTY0jq6VyByqNcrC67gtuFKYJFr25SKxx3T
Imb+P8n/VrpfEALlqbOrx9BGh+QLt8r4wxjzNcd+nl4vd2PpFFDvIQ8u/gIPjU8d
2T3sWKIEUHYgR7qBCkNflYQFGkCTi+63H06vm9FqrOLk5AJVKKxTQ4F5kxLUADLX
Bss1adE3W/NfxhOc/eiNtzZSLpKbCGE0mvz9G6jKRitkPisj+0NKP67DezIaSDiV
wSMtKB4bIPtQ9UWonnE6jf5s41nYhg4ctQqM+UIolEErT4RWd67UQDcMr6aR5LU9
JgZJHohBV7BJ2x/jOQkUfPjnxHJY3ESH8I3d/tBOC0u8iSK+0K+emm6pip2naf/R
MAq2vycs9fv0vBQRSt79jfacXrBem7w9d91bYUCZTqOjdnAI92vD6APisOAkxG2P
UCNaa9EFFcUlVtE1+eSdAUX9No3o4rssPqZYQC5e0j6lQYMq+IbxkvkxHTsNiKRi
vaVxV+ZcIDnNoOuyYN8Ls/v+HvJJliPVS6CRpAnaTo57bLWckCpimFrdFbxXot2s
5+f6c3pTkKWa47Y45nI79fMMF/n2AdU88uY2QKahrJ2SUOlip8ZJJM/m6BteTuAy
PhY3v4tO8AuRNpHHc6cMi12eziDamjahc0xgz+9IKcFu8djfS73Y/IxpJPV9eAxG
oKnYA4704a0fRXcunlIjFMzpAEq37WUtD8PGzRrxS2/T8wDHhQOZrWEsLuXGgjeN
2Y4BclzUpH92uiFmPB4TwBlRD4F8a91/rJBwA+Nu1cJAJCF7T1U+MB6G/NtkX7ds
/F7I/tWWFcCaKemSe9/W1f4LMA3P/xXIOQO9Kd4aJK/vs+3uvU3dWD7DKiq5cnE9
wOhBivTWUe4EwzMyVHohWTu8wF/pOuaIlPxdMNLX/1heU/1FdfTazd2vH0oclBr5
AMqI+e82nsTbxkKA3IbPJqTbvcVRX7GBX/dpJjKWwpay7Ld8X39Pz2MQKfF2//26
nd0MHR2NiORtMXDzjZcBWbsZsabe3PJYKIYgrY7P92P3/RyF9goJ+vkrC1ugOMsj
RVclt36IQ4z+jw8vnlHItpRxun5XY0bZveMkUBJDBep6GfI1y39twc8oz3/n6rMn
3UMqnsdKG2kvdoo2XJxdxB5LbK8Rnvr9XM9sGQKr4MvfN5tchp13t0SQyb6Izzgn
f81ohMVsWC14jnahO8iUQVIgpKRXrh/UD6Rc/6Jeh0BTSozh0HXMTn5qGH+ZcUfv
8FPLXio6sHBBtoMxYG+vHZR/QIQlX++tU0qdNAmJ70md9FinD70DdyhAbgZu/wm+
azCw1Y7785yoDah1g1wkzSSWq2vdMiQYKuuYt4UEod486f6ZSLUNIGjPR0ubpNlF
jQl27SBqGMQSlHazZz9WzY3Nnma94VcZ2wwMjZjZ5w82Ds9MmLczQJc4GsaNyBdC
HHDHA/1md7crluxMD8RstZidYVLYRu9QqPNn6SvCmZEJu3sRWXByKX9bwUOAoG/Q
1Q0WkVBhLdh3gipM4HVxkTcG6DUDAMEur/5TzVqFsVQ6TMcUkVsaUPAd3aNROCEO
SP41lU/SefzrO3tJ5cQjbYE7WE/KAk+tx4hxJpvMtseWcJhhOq3sSF15dYWbEWZl
dAVpp81LAYXGDt3W07DuVcct4V7cmNnB61Me53l+Q38Zh0sU8SGPtMks+6s5I+Le
m+D8bkV393VmHE5NTpIwuAFNzYQUKRxYZBv+529lU5tPRgKJnKCYg2F9C5n2OidJ
IeiJH6xMkothdf6WpQk1HtNPDvYs3mw39cHsQeEsZcG/cKcnVfWJbjNlvkNLoqUM
ul+tSoBVwUx+wh2bcVuM7v3oWbO3XxnZ5M8dcHZWCn8DV0Cv6oKv8f83kkyNKgST
bZM1lZl3xhpYKNMiN8nRhjJPCsSOPyRtW6g5tEA6r7XDbk/KvYuqd96vw3GesMSH
OwkxQOELPxFjc2viH9ihhkAdaCIHt0PotGBJMmPTxVTZ2c1iQz1BpIVGaU+kCQbW
PCQvsvxy2Wy2+WisqxIR0p9rS5I5qQhA8DuJt5k+jfXuge4evpESVmF1odX514Z/
/qbEZYEDcbc8wWxU5AEf0H5CUYdf79YNALfwZIj6FTleE27vbsoyak/TenPgU2nq
rY05iPAJ/RyN8x/RkOnHDYq2mAQ1mzflpmp2l47IYPYJokF9o0AuQQRtSWErNgt7
fzn4jSTmW93AjQuRSiXEPVW39Ay7D/b8FxI6IaqVYpqv4HWYJupHkPadxECcJiro
LVkFasu1IZsUR2wzdK1KL5TtBJvw4IHsHyNOh9Mhtacc21FKknqwZ53E/FyN4y+L
t3aIwJp44kwgGD5WLiRDMUsIczyfxHdWcAWX5e68x4+aLo5pyKqb2uC5lUZuEa20
bYhUbPU+9Ev3CscsX3pgbQnupEYD4HccAgJyKMaFCB//PKDD6WE0xEoyIMhH4k/Z
MWN9/eIPlP6HB96cR2zd2U3sqZt9V+8lnanX3ifdkcM33uaDfhaz2OfwIQkqSfKO
E7f4Rf4EMRDaZipht5bIMen01PvR0vC0NA/VKRu3GqibrSmiV79U3515zpzUl+QG
0TuID12rELjM+mdUL+/QBXH0UsGL4CycJwh27JKUaozUzQToq1SW2DS9eS3o2LIF
kQ8NuS9y/sBekuhJSdBM8sJEKByg9bL7nUzIBOLBGdCMTnDY9N1XzvATLESdB34V
EjZ9ilzsdHfSLdVppNO+VdBet2Ef4apm7EsbClUJ/lvt0hLch2hEjVxAjI9SvwHG
D1M+UUQT2OGuiuZyDMpnT5EXLWsnnCz+2HKL5uvi99olW+MfnkHzLksT10NcXlqs
x1VnHG4AipHAyLHksYWk1E+SvpI4U9RZbXzaCFW5uPlwlV5vOYx1IEWs8tHexJX3
7m/9Feq0Iov/jh/tiINDy9vebYVjU4TLBv5SNg4O4JIbWokAxLrraVnvhZBob6KB
6/q1qgvu98TKBVzgCpofwguzo42RGgPa+4XavxSEsASg05rmxUWx2+87jSMvHzxv
AQxstacfhQOni47KQRxaKZXIAak73F1J/29sbPNtwlMDi3jHV1Vr1F575yFCKwur
/09r2rEtCy4TVBTmqEcQWBzdnDRtLOFT50BAayghNKgFBsDgmZjov6av9w5GKdEa
BS8PmPYpuw0vOgHTT+sfJJ65Vpv2oMDPM05iT+JLAm6HBrA2DN9EmQy6wVj46Oks
Y9YEhtXZB89zkdKh9ik7nS3IS551X9f2SZOFA8If1Kzx98nZYfPHC9cjyNsvakTB
RW7nIeJf9Z5mGoN6eHNDvo2bEyYcFrK2iPklLDZTUCvr27KrhyUZzygj+vMRrU8+
VWRe4mY5guxWP2DTTeKHIv0QqeVfjO2jCsgJnPUTlTsJ0h+zP4SiPecwE7b2a7x7
5RGkGf27XD5BkiWVz4NC/6/2/7wN1CIQPVLb/g2gpE9vrWa4PZqHjk20EYgkbDju
Dr0Wcf453yWmVrHt0VeFV1fYEvplxSZol0uwcywqsJXVj3VufNVovOO8iyu1cIbp
lN7rFlM27aenRWJQBX7JkyFZg56NOm1/mCeSfXFsSEZCen1qstxBko3Y53GoWAeX
Y/aG/keWdCI8msTCw1xYkQHI2zY+mOhxI90V3Zim4Pj4LacurPDWgHS8gL5AhbRk
aYhrzGnadSMXZe3yHuHGMOkl3jYO+1L6oh+so6XBuQQO4JOeElBaxopnsQHUFay8
0h4rL4ouuuc6M82uVzi/aLQ+aCM5oOlOhY+bkCR760zg+2FnaDEBA9ypwIHmDBXz
29bk0jDImt+vzNhoSLEXsXumeibOb6Ou9rBWracKC4qfSn9tq4LrD/cxVQQ9z5EM
08tnloRVsmqucF65XlT3hWOK7OFkTzdX3yCs6iZ2JI9o949ocFBCyy5ZKJR1F68C
SIcnTRFZd1QS5s04IP4D/UKHfdXdqZMcn97fye7mHpXXQOASe3hgQN8e1oTmzwU/
yRT6HRZc17oodPTKsj9aF0J8UeA+H234K2C0XxgURns+z2nLDdDAJUIXegCkrogN
MW+2pZbZnQawM1+wHAI0vYhHWVFIB09Uu+cgdukZWgRmxY87AaLCJNKDwPFvvE/F
HTzgWPRpjxhdxyKxJ0CrmacxhJso2jgibHBW1FKxM1qf9rpYvhWyKuDhKQhZUeFn
ba6sEIvVsOy5IaynDL2kW4zdZqZxkzGFSEAOBg7LdI46Np2q/qvPsgtAruEfCHzO
VN5uI4ixFRe1wDgmLUOjC7Z/34V2naNp/NLSkDeuYI83K92VgkTrE06PQYlebt3h
SEqyY3SZfQQdlq93E6n3fjuFcTZs9Ql5YST4m60+gag5XHXFpU+GLmYPRTzE+Za0
t1cJmb/ECQCfA/2mmadQIuTiDBG2X9XP/gSa66yR7PmqIURwnW63/mENaA+KUt2g
r4QItMvVvvHDlE35bquih2Ocopt1R4qR5bC+ezHtnYU6w0UjoRz0V6kKLJ+6AK1z
tFV4wmH6fW+LtNrLOHKnbJ0O0uaT0MFlfhMoRhkURVKE9CoL04Abb2SoHFc95Z0L
NYissCwO8KndQlOoX191ZC1GIkhdv4wvqw7wTlOC5hpPlSdsjBUy+BY3LQJtu3Ao
FrB4jUVo2vDURTq2DpBDTl/zZGpyYznUD9t8SxZ7dg80frXaNXgHqRujd8VUE6LL
ZhbdCQUXzmt+JEWNg5tjdIdeK4BU9XPnQN1bdIwymEC7NrpFI+Bq+ZdkagqCvhJs
WZmjUGwF0KJWmCC/yo8K/KhjvFU1nmmWev0Pc2aIrsI4BkJ4B/4rqZHA61XBKx+y
2EOd6do9mPpTwfNcwv5rCoHPO1AvAj1xmPamEyPvFFnPfq8MUyQEMcFEfDDP0hpX
PrAl/hl3V5M9U649TfdblVJ9IzoJUa2eC+2O7eb9BwU9RVzdukF9dOGg4WSgt9nZ
WZWsfpqXCDyvvF2hq6BK1JElX7n0IcCS1NHSwGER+Rk3oPNL1pbfZkiNBqmMAsOu
M2PAlS9PMmbIhpKuydts+F0ru8CufgMbP4ebiQ/6OSAubTjwEQNimd2ZrnqAEFhj
EpYZO6oRze+Ui5651Iy3MStBEom/y3adQidC32DdYJ+upHSHF3286gZ2xjOw2qg+
d0cXn/cdAAzhCI4CdoTh2LJv2YwJHBdT1FH+Z1gFOk7g6BFRrMTIhwWslpuGGPAq
6R9ldN5GAZKK84HIyo5KkkT6eoCaj2+cL1ZqJ/acoYxhWXsZ+SkJkYeELUXR485W
oQAWtVEhYGcWfScXyaG8FdtkrfclM1ij2UeBqLtMliw1yveVGdQZ6+Z3PYTTJAAi
iUz+xksiKCLUJTdBMNjTSXtWlGroRhmRX8gsYgOnSP3aAjAP2IIrN3ir8KdwncUy
lveN3BgWa8VUkbQwfAFsb2ZQI7/FnTMSgjqu1BLS4pGqn4UfKHwmSP9BAESbH56G
yKLyYeYe5h0AGIrJbSAxQ/wyrmTxuHZKQMwXWROQhugRtxI0ocgzScHZWGhJKnkT
suT6flXfHfW75ZFsNlo7DPzYm0pOuD8rSHI/7cB/gwDidyGq3OLIdPz4Upt1eKhE
zPOrRTgTzpjj88hCr+m+elc0iR1VvjKtIJsaO4RkSs/+Zp24vZjUYD9JMv2lVg3R
/uy1Zg2rl51tZaF/I/cb2wiV+KVj1WLuC0OvIdcTHlC4v4JtcezBuQhJnd2+WDvQ
YyhgqqjwLm7aO+qqbQ37Bn8/Y6UW5uYwEh5Gmtx5rsJu/T7wUewrdXOSbT3PBpaL
eCRm9eZCD9MghEMq7xc0xtEymRyZ/B2QR4Ido3n7jz/yke7/2AxiZqYMx3WJTDqY
7czNTDLJUWFZfpO6dhKRd7AvQ3ff4mS/R2IKC9gLQ4oISHzi/tixHIOvk/glmVeM
vzLTr6kKT084syTs14/WXHNvtwCIE+zv08wn2rBxwh9VRNLUPMBhfty70t/o9QJ+
H/2kJDCMZ5H0IOVlt+DnGWIoOo+7Tjnqs2EPhB5QQjeMJ4q+VFLAKeLYW4R9C/8f
BsNKmdNAJAww+tlKVgNv+aBhZY3jJT7zu1hzmYye13bbPjVeHKPZDfEfOzwV05VK
iyI6vdRcfFHWl2ABpx7019wx0DWVXcVUfppL5iaiXREewCHgnTqx/Alt6nzXpikV
DrOBKUuC7CksRfO9fFr5md7HOigltzt6orcGqhIhjSw4GI7C9eg5pj6fudzDAhc/
o5hs+cpaAReqvoh/xeuyzJGSNZetkIXigQB7it9rnona2SNCwl7vSPMucAt7sA1n
SQqOCH7GRncZZPYWAaKwT4X2L0Bz8ZreGs9r39IpH/dExyszRn7g92hNn4me8K+I
AeXuvhYUCp47IiKWc7mtfgVWbkZQzGGI7p7sJLZUHcVwYmx9uU+eONXtzO7cw0nD
aes910dEclC0S4ZlWCgVdfQb0IRkRLy0eulYyKJ6/C4GtSpGclwjRHUF2R/5eXd3
t9sgcDHY8Q0goB22gnhaotkUSS/pjDr64WoV0SE91ls96h+BAOYCLw2vqZ9a1iAZ
NENj1KVPGhmaDIi64Zq89l62GWYzjTsd6r2D8IQONzTc9Xm5lb+Rs3Ktv4lk9FFV
F1hLsdhC/BW8Fm2cuNL5w5fcFKQyfs16xhDUMeHu33Wspjlc+zEBru07QlktQIrq
eAZPx3tlz9m3qgByJ9a5bLRBlJybgwae1czIQIxSeLzN1wGRY77GRsTm6PbUIrP1
NsG3QueKo3pfcvZEgGdbxi4ihN1+kL91yb/KrBOfyugD9pAUYXApflG9ijx0PCM0
7SlQGg4uhHYauRTQ3rJGtegdTh4zzTDvAvs12ujAl9rljmm3LPhbr9TVSRlyKb5y
4pY5yKV9Y5N6b2fFd3puWih501zNftoce07gzCvIxXpML4AZvkj0oHzdEaMKTAR3
7lTcQVgxtSYGY8ngkFGpFjHBPMWy93/UyPYTqpSWx9lKsNHjtGYa1ykCrMm5whQ1
2PVr1eAc3HKdsj0HGhVC0fT/LkX+m9OaW3paXS3HzA8taa2QDMFfXN6bW4ADv/Ai
lbTcZTnokuRG+QEPPTtGsgU5PI+NAK5XZfj9wmPTirlRyiEzQ5fj01Bbrd3t8VHD
bnIWl9q5iMmjsCPKmHq/2azlkyVwQ34fjkN1+sfwljaYFZRJxw5bGSe3dO3Xzjja
s55asn2BNxlpEpqEIjNJVBb7uzaXIxDtkBTMVtKkp1cxVIewpyY4MpgHKMSUOuWO
BHRjGHnReVzCu0AqAuAWxnNIRNuTzaCkGrC7LbFPkk/FSGsCAcRtdxqVlIYJYJ7B
37iYSjngM/xdQEu2wm3gypCU/eT+hUepHnBZtxB2LciKCrbnty3XZ9uu+g2Bh1hI
TnErsqjUt8137TmF3FZS9anx75qiwa65c9cqicF0cG402OQM2dIcqE7iDXXTl48Z
jHWuYE5ok7FAyycgsaGvVgQg//0jScwyD8jIbUez/D+eZXgezNvAp8wslmMJ2WMe
pV+Ilvhyzl6RpBm0VQv3uuyoXZZHZpHAXbjMqZgSy2oskX2cYHmi1zbMycVtoZL8
bUIOt0QFo1ElEoPthg3vawneeHM1ew0wfTaBSONWsM/4Dm98v9ZiDvb8YsXSLXxu
eWG4f2xeWCmkEtVdoJEOpX1GdmZhJ33CrSTNv06DYcia+zGpGrdBnhtMxa7r8s9T
8j8gdp3trrJJRU61Bs1j3Qn2UVY9S2h2yAdx1y7V2dHXLDAknu4LV8WTpiyVuvC5
wT8NLd43OWTevYNjoy56twIVYsp29VrHPEDI5sPMwjyQ9nnWG+f1pIMHeOW+63X+
ZWjV+gm/Oa3JxKof8HT+7xbOWRoN+xkjKd0Cg79rd5S1foymg1thmiKuthFuRIZW
yUaG9GzEctoCcFbXQY5Goe9h1cICi0oyMiKY3IlRYo90e6SwtGq1fgR4KY3fHIa5
aWjF/0bMVKRYnv4LAVd4G0CyavrtnbbYWgFmxMLxkUfjZaf4Mxec4zp2bxfh74H8
J3T56ZGm1SEMO/2oBNwQh45aUpxo/FXwPVGuiLZZAVlALnZfDGr8FpCUpAJjArFH
RodYrOH2gf6RMvpDqsY4KAuC/qZOLZyFZy0i8Gjim2O5KX34zPYHrkjiELgC3Xbj
mCxR1Ns7xNA/FtDJynS/cU64qZbbuR6JPso5JQOWEwp13c1SKHaHbVTiZGvDgGDF
5obqESeXdJcMbbSTETVKRlkObQuzsNNcQVZKJOlfYaHZCHycm1JB222tBfY5e6Yd
qeKeTmQ/70Cuf4tucA1uCCHLmxjRevzKXXcHdkreatQ2qUA4FMjOzjqQZ//0Tm6z
VohZqPXhHqDiSUdJke7wSPUWg+RUIerc88U6n+qaOrGUo7q7D0RPDVHM4/AgFQga
pHVgqBVTtK0kTtU615Xp6O+DkjFcdzdiafSqpv/hIt5uy/TSKVQEudkCLpOgeNRw
mgxInMmra0CQl0PrHRni7jzZ3jaqigcpVALDk2YVlMz5otVEhGpVM2iQOuo9v0bl
fwjw0GDY7JURFVECfeGQXw9XCfQ9sP1eUyBH1xMgyY9GVSmdjPMAxVrT3ouCV6oj
J3r5dCPqNDfqljfoDJK58qAeUyFhuUszkktxhMO6TGNy++DY8He0Uww1/8zDYXkw
MBTgDU1Bc6Vs8v6fcZtqDNpQc8LolJQTNwrUv1vvE3EJ1CW/G0CXD2sWn36Dorlf
mpIq/Htg1n2SJpURDeRh7qEJerIpHqpiYlBhhTvMKL01lh7m5CoCPMY2ZmBbADNb
70y5u9kqqbwBLTstNEwYemx+Eyy9tCdFKF0lRHsu+om4tuUomqJ4F+5bXfH6MJZ6
djefV4tdss0+Q0PyG0bJtwgbEQb4ZTK7Mnfgux59f8KvB3LQIk/4UiD/PxEU1Xa5
e3c0f+6alhGKy7FcPagK8bbf+iZGov7b3J+7zrPZonVlT0AZbCKz5voP0nheom/7
KUjhsYc8EItTfQL8n0gMGjCsE0Bhgb3sV3XfLtwDHePLZ4s1lFzQbm6MuqNlLP9G
aX+whU36/j99blIqHk0WvQ==
`pragma protect end_protected
