// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:30 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UpRwmQ1SAkK8rZfOMAK26D/z2bWQruGMlBHW9waQmD+Prhh+Hgbq6P0XKia/r6uc
S1rJSmPaakWxMiXqFNss1qX5HNBwSK7nhTu8u2dIhAADoYbYNjKE3DijJJ1Gp7cE
19xhbXHN1xXxB6BxO8j2iQ7l5Ud1HovRHojksuaSb1I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 61648)
04+FIQM2Jq4j+0+oLOzhU5tdrbouS8D1MYwLkgLpZU3zrrraJ0EN/6zIuF0xNDrz
el5GaMlHwRRIRU29MFSxYotoVCeIqGWU0j0DEGXG9wKo0+m0Ru4VTl8bDQtfm8yk
VQUvlXRYbOlB192I4r8CYYZTHVCUbRHqPhCkeSgalcIbgNyn7BqnTLtRMkpY374f
RFJqiOSwp1JuK5mFDLmQi5MDD+PiFdcgqMYBS6liLSxS0m7oiHjdrFUr1zCZcUDm
vwuz0m+3ywEcT1Z1xuakRS3rgPst3JE7eRO9xJQNcLUSKIlPDB2iSIGREvWleLxF
rKAcVB8h42W8PWg78aIfjOyZFUiiLM65yotnwdZer5uzKxfFc2HkI/iAQsTvs5Tf
wvCGBkr05wy4x++qNulcvHcSeMYyNMq5N386rRZ6J7cpXSyPXritaPox+47bg9D3
00j2ATFLkCPyAjZKm3vWVLxfpyZ6+jjcRweHf664irysQ39ZoDt4XgyjjJTfmDM9
87XJhwCrcuKs2zAIP7XjWq+4GzR1YaT7aIgypCCyd0FPl6dWDeiaNo4W5YmETWDE
Kof3WhaxXmTuaMnaMSxmccx3k8wwLL1MfrBi+ljFuecJAGn9uDj3wy+S7uYGrZU9
mgwo+71TWBRipcNuwcVkSQF9NltUvaHquPGeOnq0yTGFDzb+gbJKhsjoQVvZ0vLb
YOWUBvpEStIOVkCEXyfXsn0oE7/LUn9UmU5gmDV9Iu9nKB20w8IhDbpP7X0/DY+o
QuKKIJZVYw04ooo/OCOk1qjJ9sCeqNYa2s3wIRTCtv7B1kAuK+pMZ1k71Djzz5j1
mGMRpDKPYFa16fnFPu6NQzuteDkyzWlveqwaww5Vac5PRIDzjHksXobbU3Qlkwkk
3yMrN3OZztpxiNcwCuaKDiz+zBTAnTe5Yqvy/TO6K0hCR6Z641pLAQj0Gob9Lgxq
L9NOt5Kdtob7OiTsWLBnZzeWwx7kvppr+fd8ZCcN6aKxBgy66SyaYSKUYr+CcOzG
diTc2k6V/e3hoSSGMXaTJx9chtfZQzfwvLDfauDd6t9aXvLeJRCzDbu1UI8PtOT/
R5T1oYOozkoLivtHTCyI2FXwUK+Nzo+NzA80VYqnHKjDFUDZt789PRVEaOTGLmCc
CQHg3IXy/RvwhP6yJDQ2VieZy8Vipq7t+f3o2L18/Qk32wGYgjJbqOQu2ZhIMk+B
WilvVJoaN38lgmM18oKZ6AR0968+4aFExn4dQguO/RRli24CQTUIEQABVMLnJBuY
JE3QQbrecrJmRw/+GumfkgzsDpJMy5cKAyf0o2bIy5YyoN+e9IeSNT7zAcNoxL70
69MbV81Vt+p0YVVfunnPy6eN0FqyUxNRKcA3c/nw+u9moBBvKUnVpLje0grNaZnD
EsjFSmhrJAfNCRh09QZMedTZ2Zg7XLdf8wHE9qL2RxllJNqb9XRMzDwWaS/8M+8C
o92/ydIfh+QQv8xI7gbslMdK/EHS2BWdRaRjCu7h9ZkN2DCLWqP3JNeHh9PMKLXy
2fT8EZcUiVGBHiiPusmnWi1vZ4YFxWS97CvOtLCE1Bctek2vpUxLAUSGlF5qFF8y
kjjDM7M+Th1oJ7BzwtkN8uEX+wr58mt/xq4sp7xwEBEx2CywVmWtfM+nF+NZ2bTs
d0jakRgeoYX51JD+CBhxKjui7b2Lp1DFfB1V7wC2R5FNavf6VNfRwH6DVy3URoMr
XBDaoI8CJM0wJiA6cnWN3/4Kczjb9DwBWq1+/3fhVzoYCQhEaHlm/psYMBZUe7p7
w1TZuSZ6Airlj1FaldEMCeOgZvAhAhYx3C5WEmuZPjNsHfZ8VXQzLWivjGxjtdUH
nJfK02i4+NHDi5NdmUeSXLn9ah+AUvzNvoxLCbR7OhATXW/InzE+Iqx44fximqYg
5cT7KEzoEZkwd9hTnghs0t4GFdagwbt6D7k+Jz2g+w67buHSap9lANh3dO1SsyV4
dSxGvvJL8aePPLkcauDv/eIxld9bgC/D92uFXq3f8M925OohPJahXfSnLhAmjxXH
c5YGZTPngrAOoocfe8ugifOFkqR+xkwTFBQffP7iXauyDQ6mAlnksGV4xMd7SIvm
1CjRbyBZ8TkgnBqjSzi9CJJep2PECmV/04m01JL5ouWMDqujSehDUQwZKNi2nSVV
yWOOs+vgP8+6XyrxSL1MPm241DFCVD3tbRF38dTCBO1SacRVFOPc62dEGZVG1KGz
iMN20D0EEi7bP3WQowmSM2P4/v6Dn1Q7UEXiBMLZTQKnUphhNLYrxNPnHi5OZ2lr
vF4m8U6IXAULLbkPbCqUPClKj3OUpVoWc4v9ao44bC0yjfoAAfxN1lC7KrTESQ8v
vwv33U70vCmi3xZKWXL0hIxfUgkhD20yr6IMdC6UXnBpxY6SLO0abzwNlUDtN97H
VFGYbxPuUtgXjSlChmEptCmpJjvNgpOA/k4+sGLNf/G/fs/eGQrxgM392Z31h2lf
GwHJgEcrXczrOIlNi6Qz3r7KK05I2KeoAVZAKxHYvKAKTc8+K0xFei2W1DRAssU3
Ark3TTziUBpfLiXv+B5nwG3wPdhDbPhpRKUGQBL9+BHwHtP1SLGsl7LzaY5HKinI
kgULaOwUXvvdsPz7SPJBU7EzSj30BPHHu9dlS3BFV6kYUwDY94GXGwOt3edjGhXN
6+j99dZekDVRE9XQ2mCyKcNJg1UBOHbgPXCzJ9NlwGwL9m9hm87eymMjQtdsn79J
gDAr6Hpee/2lZJerhUTTIkl+gOcP2q7iETrV2+VchLD3/dg6a0+ZzT5fASzzmcNb
1sRk7Yx2ruMTqo0KxLFR3xgH7GTUgYqDmxIHX1gGFJmjFMLPPMjVskiiN2ddEWUz
XnolzPTzMXxkXkUoyMPoIJ8l/CBhfkoRjDn7RbBEDooRebwV5xjAbSHNFHLKf9Cm
pyX809TlbdL+BJqMEkS8HTS+gk5BbesHkQfaDyGe3nv4GSc2llaKWJjVRtOJRNk5
GkOfh2WrrGYq27WXYafhjyl5MyhPlaZONs8pSPmJnc7CGNSiuQ0UY1OEYYm4UcEf
xwdAaqIQxIuCBE1kA40ohHb0oYqKe8sfTG5va7rK9IM2DfiU0gLESkBTOEd/Bto2
YxcMWFajG8q5RuVrypECXUi55XvD/EKEdubDiMOh6YaYXqApb8hn/tb6r6bQHcR2
EyzlidYfsTouh72A+Vsg7RP4JDAyENfzqDZJ07BADx/njXszINnR26TuI6O8jZSa
EiRtjn53UrIEdhY6uTmBg2g+kN/QyE2qFR0ZpzGPQwJxIBd06g48zo+cpYaOri+C
dNvKzuqtdwX0cGs6fyGgf49WurN4HjtOroO1/KBvlwUyoJlXND9NsrkdfL2ej1iO
m1q5lhDOOlv4cAQy0kOyhaKhaxVmE3T61q0LfsGPiS7B6RMLJXbbUQybyCwxgiM+
fIO8AscLXQQ/gjx3KrfYJ9kk7dcqDAMFp1wpMfnc5QvXDIz9MUsbpypzt2YOTggw
Tj0yQEMp1npPEqBvWYs0e90H1EGVxwXFjiMSekW0u1tXHvthPsmfYvkameRzngkx
ohtxNgliKcpcsKxUBLGJrR7LzqjaQtTloH5yNo8bo8CbXQSpcTTUpYnXiGEM/Beq
+WeazKCHXPa3Jke5SZC35JGsxSy4VQUgiMn0AQDf77JxBON3h/MwCPkksTuxOJTH
dC6IRuMKTU2G390xLruK7d2Jp3Lr7w0Sylq+vsXCDoYmfHPhssbLIaQO6k6gbZTA
mZF9G2oIa6kdReIGam28Psoi9FG12VVUH0AmdBUNnt39yPe3QkItYwWld47dPX17
WwPQXE4RL9l1H0zwtSjuwkOF+GQW0/J2o8n7MBv4qJ/JIeZ4Q9HigKuAEyMuQCx8
hI16IRVPJ3d6PeDU6MSeKqUY/NUXXjKS98ZDCTtLOyegTLOdAUvOvNwcI8O/kbkr
f1gaadlRxWw+5uW2Ik8L+mjBnbfz4S/ZP+1tvt+YqX/AK+Pih8mi/yheq7z3qjGp
ZNChf3EVHuYLpUE2eKXEUXCUzgzvqXbGyz1s3bBNIVu26Q3kv4dlPNxJMLC7m4lG
7sPqiNXcWurnOgluo4HEBT6ALlG1OEWCFHBXm5XoH3H32V5iPxolSSXFWaIVMdYn
ervSMiNgRP/nhU2UK3ptysjYrQsYsc5Hd1GiIqOICEB6zhH86j/aDdMkTvc1LQ6O
RjH25gvslhys/BlPrEObAgKZWc3XWnOZFUWyJa8OLcBPSH4fxHqHakbBPY7ISYhf
DQVwCn/Glx5GMeJioPJpwpDbGP2KjFFLedpf6YneNzKR9RA/l1unQLPhiXVTyZCa
EzedWnEDKtNTzxmy7HUF9gdhA+rsCzVsShHw44OI3v0iA2OhKt23nt7Iua8QbPOg
p6/As2Y/NB9jJoHhVMWVM/5Uc2y/U+cTGnTnYcUYGc7q1UX3caijRtsShxOd1Ryn
BXLdAGG7pIwwNwwrxTvMfR3qQg2n9gCkrlo7VuxasBac4fEUAPDvFrupoQbhDyBD
/lxF45AtU7B5g9QyzW5xwjhYm18AUkKca79qtg21yq0R8QLqoj8WmoZBwK83TwDm
Eu2sO32EopkOfTqrsImSdGiKo2+vACyTGkovskPlmCRx0c9baA9v7NBpu4b9Vk1Q
0gsUYKg7TJoplhMQblgZ6z3/6y3GJ5f5leL84OqDtKa3PyFdm4xxW7Rt+0oWwKpr
1CNjnBEz11n8f1ILTtgmITfDfb3+3jalVmWHWSF6euRwSYYg4YxcUiv/JYPenNOY
fC0HK897Lr4Ec5iD999nMTm4Ij1qR5gKdsKWho3G3zVQY8+EGVZpjQZAh2cFGG6m
Q7wG5LzBnQSdhIVJ7CZ2dEmx7YjPiabY7hyUSgnYiqaziTZakHwqQ6wfI+3qLya3
fmzup/jJELlR1kjkca6DQUqGJ6T9kqGNzLbaIQWOVsyyrWhgB7Rc77DRmBjxsILF
kkZ8xplgsmGZ/ltIiQq9/Os8aOLLxjlsfRmFwlnjt5CTsRpuDGgj+QPKOJ2R9kQ2
yr6cL4Q7uiw7k9wTqGIP8hfpWH50pzdt8VRns8I86IPfic175+zp0z8XB85ehTz7
ix2h89e2gpppbRq6I3tp6ySk15yv3P0Tnwjk60vmhAjoqZA4XdibywR0fv8Ga8zS
7WdRH9KDeOm4ByyzT0JWhhI4O4INecI+2kspTTreZOPmmTIjBXGHFFhLetvhB12I
whi4M+IFUhEoI7V9K/Hf3vkbEoBFUHP2L5TU4vqQGle8J0yVuUeqg8BEjy2PJ14z
QjD2rysXYSHm601ZaqXyGeh8jLl1G19f9qh3KNysPPmDYKFMVIXaX/JVXA+PUO/e
tCEDdVlxfQafijplAjHANddDfuNIazcggJIlujqixhD2zQm7VNJ7XcDSEDw+vvOH
YAvPyoBtzXIHiHuYXAIJtkP55zB9V3YwMxI2H5Vdr8tybinGBk5kC7ZmlAUVucQf
8CzNMsjbxObwxaoTngm48pUMBbAWaIhE9OrG70wqgG67tiac3F7FXYnB2JfFb80C
loEHOe3s0mh3xEjiAD8t+d6WozoFhgTcrAq8sbEl4I3AsnI/nrbIJ3Fgh1pAeDex
mN+BP2IOOZQFiZ6LT0n1nH/DVaXmFYNquBzPK35AFDJx9mw6oRMfdDn5jrB4rTHd
0ia4xwQD2U2jLj2DP3XGMeO7ZXRYKm0LqF6Me4dNArrK8ycq5XjJC0r13CLp/SKM
2y6moShR6JBQ/Xg0400lvWUjsnuRxsT/VAZDp9DTB9bVjDRbXw6nKb+EkLODEHih
V9g1WgNyZ/apOtHYkRivd/5qHlHHFGsDfPEHlNbVYB3gh7Esm+GDHpuyY+I1X1Ri
2uSpzQXyFjZQo18wcva15Sr52nRhypjFKFLnNqEai5PlovFDTZjNkM/B4QowWi9M
QVVg4QCG5LPJc0iQNjV+2k7huLPLlErKmi7VT/jvwg2tb6cwAJbb42hdsG1Y1ENI
Nd3Oveh8Uix4oGtQODjhha7EjLXjwBQ72+RRJ3hsaD01YPTQCI/akvfVhstiROqA
vuv7ESWVuwvA7/VikO0LiBo0URZBe1W2kk9LSVuxnJczxR5K1Yow4hxJq+1Hw5WD
zYiuy8qWogh9vtj3lphHw9v39fsRcMIBLdaS1Am5mYK0nELOkWrciC9UwZLUUSFJ
XzbIIsnQzcNUZj9xUxduroIv2aeThBH9qYBCglN2q5AKSL/E4Hqppbn7Jz4TTv8U
2UlQqr+pTV7F5J2BTFSTdEok209EtW1VQvlNRhBY1yAcwEmNTKXOQpCfK3POChNj
OgP6IaznZ9/2RxULEPSSzJlnuphRA7DTlXxFyi0tF10PUGO6WQQ7VHKWahfTliQD
SI3FB+whJHUZHcBlWO/ocXO3mx0bBGXahlZqfCCcq3Pqq1T9IAyC/rEM14mBSaYz
B/gXPZ1xNVaRJXShhAIUbhm4DEjv34aPDp9HQKs4mQ9++h6TH4O3DorJKe+7WhL2
KZk2Bei4q1XFSmPTJJqgCz6X+kJ+FqBwC7APyDwrR9ZFJYDRilvwOGpG3DIQRdFa
gVmp38bjuYs/YXJy3blaek9zJ2JDET2XUgX6Dk+IyXo4fpK9ei9bUI713UhnTT1P
DYC8e9CnePyvXSckTOUeUf97H4LoNLg9q7wZq+ze57/Iy3XFeHXsZQfXDSgtBLqu
1rtm9t1MlQpVph9rxn8znR/j7tJ0ewDh2FoDj+OuUCxucDMpAw+ssMch96jXAwZe
4XEjNR7arLBsjeTPPkU2/zjkZV18gr8qK25eBUbInu/HMySBvBgnxrIKQ/TdX46i
QuAdqNxV9H9j99cGJUcdMPG4FxsAdDgWXEviy0/6tCpkhXaAztttUJDwsE09jdiZ
oBseT2ZMml8JJGE64jMFalJ8ry8p4W3SVDLaHj6pGqLHFG4OjxxMP6894WlDtKiS
w/aq9N6yyY7DoGNNUBQLGC7wgyVFCMWj0sI/WRnh6xvyRY17DyOFIzia2yLSJwxK
9L98sXMJLIiokB3b1YcS1JTE8ghcs1jT5cd6tZUJcwUUMsEBTawteNHNQWD1a8Pg
Zz0BjeEyYm7GhxEMj5tIqOmXcZ5IbchJ4xpolhTkuhlfyZOB+zDLIS0V/wmrN+vb
PbJEZov1hldvdjJfPPdK+SmbWS0YvMWkQ3yIuUe1fyLJFWIfWSs+N80T4/zRpgUr
uwabfVeY9qCAGWEgPPYm3XJ1RkSJwm2WgRwzQ3C8kPxHrEZIqU19DUvVvJk/b9OY
9UA2GjC87rRM6wp2gL8cWZ2lcwdezSVXPYIo0ycNOC+Us3PCAti0uH33ao78PWuZ
ICKW4HaWQ2VHp5Lgmp/wt/LrIzDwG7+LsJYooTM72Wpn7eteW/QYL2AjD1+svikB
zNRF23irhseGX0xM/8NbzXbTuGcVJ8FbrI05LCrJEcT9DLsC/3KzJMfFQYIPQBfV
zsRL+DrqnslTrzLGMNisBUBLL5viKGqJfJcmuCmHFZvt9oVJT/RJl9Agyq1l64y8
Xqh9AtjbX+oNyYV8DlcndXpoUDJOlK9H4CmupHDNiXAoA0PDjLKuXMQdNYXYe1X+
Y6t9lww7NqSAqGBZBRx1ITtVHZPIFF7hBi623eyx5+FUF74cfxowv6108qzlydei
2YlpwCr8yLgs6H+Vhac7N3sCY1LwPcJSqmnb4qdSWr+3eFwl3H+lw4LrLjRpY4cR
DgK+nnlDn2DgLwvc4NDEPYS1CCIOTXE1F6lBhLVpUP58+bkvbEfH7FlVbp7siqWm
o7Qkvd73eBfPixoGCzjUu+UQ2CFxbNSxpgQA5+9LbNLHckUKuOVlyjmMxs9hdjnj
e4POCmP+tCzCLS9qN1mFSlvQHCsHtOexon985BBDPMSzQ7uHExlI3mv8BzMonsyO
KhR4nBoDYq2jn682d/uXgvC4bpEcZad+UeRMhXFy5qKhjKp8QwnzbQevbYpReIUI
+dQ+OF4izw6St/6/MvaBs/eBcdU6bqlwq71yT9Q7F2kmZOWLT10iWb60thu6thDO
osz6K0mpNL/dK6Tp93NMXC2g/4qlpwdsRsm6r45Ut74dYGPQX00gCaX8U9wwZurH
SCgjpt1OZT71P1J8WZgvEc+OCs0Iz2S5smmvPgotRumA9GWsRn2zi2VTZaWNk+FB
noLPje11t9wP/n1CbmGIwEprcSq9kcV1zNILzavH9OolCAwHoK//Cx2pjUX8REvw
fkARzroy1HEc/ytTuiROtZJ0sl/1XuNPX30CM9ScLka7JOUENPMToE/7bRKukXsT
jIgj23Oq3HV3Q+S8+ZtOD6nBsBLVfjDgZ1Opq7jQQH+gSGGi+f+g1hQgpsUYGbDF
3lpAdfGxY8OesNoTUBJUAUNdWR6e8MxXWZTVNOHW+u3A9G3ppsNtqPWdG2sCLj6U
ibG7qhOVZIvJNivYIpOp+jMiPo1nEQOsq73Fit7mRftF14s6fndwD8xATmjC6vJH
L0RPf/G+pIct7AJNyoYQaIjn1nqpJ8BiXaaGtQsI1Pk8wmOiOSOgSNCUBYTFRD6d
A7BohVVTx9mG6uQMj8WrAWZxM8rqbZiVRnJICJ6rRPwYcCVvpLgIqllyRzNViwXg
9/DYPn9TgpmKqiDUVGH/Wa3fp7nN1Att3h4u5cLWQAkdQyg/X+RZe8obdFsWNBFz
0qs3da8GWv6J6eONY1mi18nYjwjYdivQfwapkhNov8TsbtTjdU7aVIvWPpiIjwhn
zFk6xxgN6HEolCNHUmPRfbj4JVFixXtd7zbqxUNeU45tMnsewFy/b2D36WtJFZDn
ERHemvT+zyC2tstIGOhgZ9VlRNYslxS5l7N4oLBLnF6cevMUtDUCrsUDvqrOyY3N
2JtVOK2upW0/54XJKws10LhOQ555Wnc9GuRhr6qTmsXnztldBdwJetY1UD8y+hos
mpVbShv6NqgquC8moA0lp+6kQG59KuPnjuFn0/OAMHHhdlJlNg6DALfefCFN/lYa
i4ssx0lEsMqYUvgMphyP69leYW9+ywA2Wa8XmvyPg/X8657yysedPHnw/bAx0B2B
+WD3efoDQrq+s1UliOb0x93Fwca1dT6xFI1cT5TGWaCAavVtcJY5aEoPjy1SgaGM
Mnz9KswyIcNl25/clia+NHOrT89UgmDBwJk9duEKbtwTY5N2GHUEiD2ZyqF3NaSd
1Ki1tdFJSJV7OvXiEtD4ekdkw8SEE0ssCZ1K1n1sjdRkBrDOTu+AeHMoQVMUq/Lg
iJw1Siz/Dod+fxI4ynFtRGX8tGgeoen0ppWz236WdvGWIi4Y1cQpyZMckfUPdLEr
a5Vr4pDacY6IWDqFHhXqtCEGTOeAzoHOp3EX0Z/cEz1a2ynRk18DrqHPBc8poWQ9
qAlS8cE8Z3Famxy2LPLnOEvXbbqOU8VW/XzWd1xVwq0LlqDopr4dEtrKryQNsELQ
k7wGX7oCFBvpSi40yoIMwr6/9yhBgN/UQ2N0hwZhZeEoQ+1GKHxaSYNilSQAfC1M
fHnm6zD2upYBDeNoIUN74mvlSNOgrlHGn6bBJSVleXVaZ2qgKoSRA7pbyxV+lt3h
SobVoL47O9boOtkpROZ9TD8I52UwRduwSg06+EABLSLFq0T1EdHvktK8pnZZy/Xa
zigiJtvME2XuSTbDT2NGIgeVxaQAKUR+miPzNcC00XyvNrexUQf352Ce24B56075
ya42sfjyECOTVIHCrgs9lFp6q6PMeQCxbDKSWDNFsPjosbtMwcf5bg5d/JbyCHQ2
nPQkcDKbkflYjFhLfhuksNjgDRgpkH0WU9X2afSO/MFnyvnK5EMTtpMuw9r4+5Th
Ao0wdai2ZmfV7OYHGn6nYu4dPcfvy2LXl664Xt4AMLi9Npvr4ntNbNnoRFs32GI2
X8wfVUQBdjVtvt34Gmap6Ml+rDPF08hJq2VqSPcJVdvGIkVpJlCntsSs04bGx9QV
zrHCGbnFZJYHb9WolKo7AoqEN2VTk/DERVWtdZzYHy/9A1aNw/nxwTsqYeVDHbja
TSP0XOuB69tWmIkWBRDTY52NyaZdeX7X0dhba/dEINRXi7h1o6xF4Lj0KewnWvjz
xFe1N5wwknQTn6gsw7bf/saq+ZfOM5aAySD6C3nYCfR4bEsZ464xQP7k18m/vbuu
1fgEfMBiEq9gBm53GR/ZrQ7Appoc9ReFGN8t4y0ScRCzeeKlQ7Wc4NW1vzQgXRbm
gUKoOX9kJ0NT8cP6aJ9JXh/Y6kqwnQllkfR7GbN6l8J+srgBr8ZRqvbYpekLeS27
GejHp3cZBUTP8oZEi+IT1mCbUxBzFIM3AzCayQ8llspLE7w7D7ysI9bd6XjPc4w2
cvNGHFiVybIcux2nmKdzosZxHW23dTnnanFSAJoFfoY2pblnvwvzZXAwy6hqSAQK
aYmUw4jwKMpzORHdMFcaEWB/0KflVbZH6dd4w3eYg2uCusb2dPpLv1Q10Rby6xVU
eoND2A7rUH8c+0wWhXkjR82iB956tBkFJOpxdpWWPGzQDE/3u9KfJVugQylS9BHW
OM3SioxnjseULjhQo53t4eeWC7w9LGWIs+zaPIsGshb+PQ2IP7mWQj0uuuY/ZmUY
bJZAnBJlg1gNaDMJpiDT29HZVTugP4ZvcaMhqethuRoYaB+IcEmhstnyXGLv4jQk
cR33WuGuxy/95JGaLUn53IpnBYjqbe3xbjyepD7paRZ0e5v5rmdvet8ddbp5y068
z7e4mVFfjP8SG3fwz0qV8drF7tGtWIWedJe2xRr5lnhxlAsMGib4xNkz1TaWl9mr
eJOcm5n+2kduflUHsx5cCGnWFUkGsYWw6gd3c4usnjQK3Mfz7sDQ/7dbN9aJibcr
H5A3QjsMxNjSS3E6rO6i9s3wNEITMX6vfPV2rDqWEadBo+/FBD1NRMRQmw1ZtcAh
PZblpSuvrbn0kzXeDAEquRa9dzXYk4mOfQ5zKDoCwbHHnOI9gNdQeF/x/05sV1X8
3PsIytE6XV2gFRwbB8dtLMhfoZr6s8D9U+0ocXITyBdhXEVq5LO+eQTvkXHACOPG
jBYHAr3ykJtUk+2nRDGz1HbNJ7yyBqMJQ5YQXv2+Os+pTYy3bh+Qs9eRr8ACGAeL
AvMl7k+CypB6wMeFQdjM2pQ3p0Pht1o59j6hE5q78yPIal9vxoQt/wIF//vwSGKb
Ol1CZVH5qulRJlb6/FwRBtCQYMHuDLE7k81QZptTBNCRhlYQeMhaHyest5fGUHtv
D9LhM2BNyBJi+6LlytBA+p/VI6oq2emcsYB3zyTczHTUF4CjZ3MKU1eR2ak/o0qG
NAJj2ZEcodKRGs0y3EaDTnGyt6Q0k/HxecDrBvYdp6l4BpJKrmxm3QpufpGBwAbI
TymB1UWB4rk/d+sP1MAjLO78TtzrDbJrZQOk3oVYbO37/f0lgjI5yQJydnrnLBjt
DDSW2ojSGNasOF8+mbVoJkymNrVGT236an31UV+dBYqu8qNSObkodXH+jd9o591x
IRo2qNmC05kKrS97C0NwnKbaPOj1LsipjZGkWeV1DJ/tjlNVJJDXmsZ64d8hPrI6
ZQ7bpw3qL1CTpn5F19IYyoDx4L3YWVGhyyrZwNYl34CboMH/TX3aW0Y3ZppApdAQ
d24rVJZx6wl84poO0q2EfDS+jgfjUG4KFmr18eOfoH4zPAfBOEB+jc65U06Yly+2
EQfsXhEGAkeHO2WFuTGaJwgpmWzl4mpyA9Hir7FTeXF0DCIAdsbF7RKxEQs3O6X4
QzWthviEAPbMnSnLJhe1OpP5YYDbsXSfSVcUrdnZlRjBpbQRSdEAZOm9W9Z7zc8+
oB6PUJ7MqwHVEFFx/aJdDSViUbg4pKHahjf4xfJGx1u3n3LE9WAEFvXYDK/5aetf
3fWdbZP3bYTqZLc+rzyF1sse6fCQ1BG1lA+JSiIHRZwRy6YmSlOKJ1OF4/foXwIz
NPzJ6irt1xAr84I6uRnN5+aj79YQ1iOBA0tDFCyPbXB0s8By479/5MHE0supc8ST
kxzjvEKpoponxvEjBKyrD1iD2HOCCkzLjjg5E3NRwJ9pHixfF7uz17z0sI111Icv
rnW35xH3Eu1aVroUiwGhKT4V4H9jjIzIn9pIVittwerTgTxSKqrRK8hJ0vFXUJNa
pXxdak0CB2ItjgQB7MRAwQtflkAsLLoNuJutvSQAzMPioiSzhzlgetem+wV7HPI+
FfqTwk4QF+0uc7YD3fyVu6jCi8leo1FTLcoAFVUmQlcIpSS6ObLbPMVSPSF2cxss
KS1LFXUErdd+SMFG4B0LTP1DlXuP5ogTbisWMCFMoKKNHg6Fbac3N4vL4cXPwiEx
8pd48tjI19ZzHIxZRYZhfb/mzLSLBpgc8I3u/a3CvtL3l2kFVzl2OnJMC9jpqVv/
vzTAikNjZy6+kHtXbkEpthGPhadX7KXD3nBV3Vn1NOZaXdRuzuFQYrfhyYLD3kTE
4087D+9gkiuaYB3+RVhFKO/Vstm2fFD94QwVa8We5bTklhI+LGcaYd0W9p9g8J3/
Bz4YQ5njK4djGlc/IhWQHQFX+lVJk06yoLMAWgv/PH6tZwloyiTvbbSeYOXZmcNW
T3ViHPx4VDC1inF2YHjoXpx8/+wS3P6FEyTNiFVlG6zFgon9+KPvjSyGTkt9ijHP
amDobRyTzpjHr+cQhGZNGxqn+eBkPiiZxco0sLlVU/eb5Fcg0czMvtINEEz5crtg
M6D49uHXjC7xCuNIaHPer7QtAqA0TPHvbvjoNFfmbs2WUEhXcySszXYEyMLp8sns
l3DSn4huOMzGaaVW9kCPL5VXX3pkzBK5qLbkiYNvgOvg1ybvjiIO0gjHAHLT5mf3
m5lr2WTyDyQGS4bf1Aho8I1CMYRjbfxRauRKF4VK8ydIpAo+z4P+7ZXCu0rj4OEX
C1KnEAEmlx88inMeNKcAGuGjSjkAzt2bgWf9kKnya9eIitSOPyEvV+FUqWy3ZL+o
GT0OhYeR1a1xwKYjsNaXxjqGDPatCD7IjqX5M8ZKvBmW5UhfemEW6DD8wva+dQ0d
HVkVH2b6jRA/NB/eJACfqDdpcv45S+I1f6iVkWyJ5hPRHkbkabk942rXgImCOvKK
N5zy4KfYRIUrVJkL/sntujOZru29Xo47apUq/vY0qeaFnofwlwOFSKA+KBEgZVjM
srTx4gpicIXyZ3QhK2zHJUr1ZCqOdHQxeZ3AY9s/kQP7Tos4+3GvwHSyl9NudgWK
0nvWR9rw4AKWd5qcYKSFNyNnkT6B58rBcynEAZQ31M2S2bJGEZisFzVPt55mz0V6
GYNoHkqQwud07nR3wB68gUVVXeFnPVEp+Fr972PkAGwdMnL1q4vikx+3w9OrPqz8
+CqTqjFJ6d9Yc3txO6NoXwb/bPdqPNQRuavuosmpCqnuLB6vViWzHb+v421Et1WF
zkkAvCVVGgjBFKyS2jhY2hshAdsJpYlzuCN0TXYiWzBu+8HLS1QTg/Om9snJ3p+7
uXRZR2kTgBQbiov0nTeCRJqhND8+x7BxUkELdIBHAd/BAcCbzpK3YxcvNiHmCNST
3BsEK3cnt/zZiK84rm+3BzmsIICaGsuRPUgr+jFtOKi1Jva5UFKB7/ZeusqY723/
6r0JjXJ88LBgAl48NrQA8N8xvHXf4AEtPzyeIhLV0QC49NcRUnCLFlxvsyDZnxxe
ip8NEOyj68HJ7rQFDJwC7UvaEGG/xiHRLnXnsFWWo/dpYVwMS7Bpxy1wrp5y2M7y
MubKcq7gJcwUJ3yfwoXWiqOniPiyBTh8ynELm0r3MJwNda77mWYzidFPj/Qr91M8
itZyq+HQz+Qyt9jITUyS8FM1toYLkKNzM993M47RjKRln4MtgCDcW6ZZgh8lZskI
TY5p8w+1LCIFwYzJBEucAMAZxTXkxqpYHEzFFtqWsXTsf99w+52/vd6QnYWiD1r3
y6J+WzIG2AgMG6My+2oHGTEhSITs6Ya3pTLJuNm8Aei7CdRhpzuPgga6e2pqCjpE
znAQp3qX37ra3/Qt8eP4J5Myf8YNeFdFa/Ymtf89gel1RBOhV5HJX1mITZAjSS/i
Crf/etMzAeKrM1agKEg4Lr1jaSCBOggGQ/bt4UsWUxixW/5/+htSvcx8UEoVR6NP
6VxZRY14CkIl7xihcpKVtTh/on1rhDM5/ojiGY3q/3CYSduOGxDIZbkq7NwXNwWM
GjNLOSsyE/Srsimnr0q2l4IZoUPkxV2mG8+yl/e0u9Tq9p9LCPi8LCl9XFjC/4M1
cUtdTvpEHOoJXuk8K99yDXrItXk0sKg/oHfiwgoE3UJ1AHnZMaOlBzS8icE/uUgQ
Nw+mBLIK5mCYHYd/MoqifjTl+TC+CFrPhwdXB1j0/bQBRG8JG31PSsSCGr/tkOLK
WaoivD2UY7269zWqbYxVh3CLqH1849qrRwL+OLMZWzVJbTO7Q+d7r9QdNB79+Cd0
LqWZid2rLUSQrBF3X1NcDind4ZeCdLwhVCXTVyFoySVYTPEHi3D+z4b+XtFbeX2D
0tPcJ1zAGERZV23r7ds4bWNkloFQCzWjn3rUtiwX8Qe7NRArDLt/t52GYaAnCMDR
3mDVcv5kosNyLWqS+KmqW7V621NNxX3+wXT5Lmvhyd3m4o2OOgCFfXpqZLIcJwPx
NbYf1EQfduQXF4f+vh4lqcqGpystyq51qQJAhuNH8IbnTs3+c4H4YlhvTE4aJDzZ
1+8205qn8hKgdG0mGN4Ds1tc0l8BGtsi6gJX1hwr4kvyU+/8SXaNRqNDv24ORpc0
MZV068kqV6qeKCk0A7qmEsrittaM0T2vBkWcdSR6/aYl5t1mTkZi3jyKGsV+tK11
nbGWxm03DGcudwsVpoaWkpMTivn33pV/4d0j94/z9L9d+NZPTiVYy8TqRRT3jBWC
k2nc1ytKtdF17Vu8y5FNyUEOy1Pm3JceFco8lAfrWSsuEbGb/VblIqFiKTXhKWuq
j8TQ27LhIS6/+pedQpYcuqo8xwLgfT+s/jbx61TX1v5zDtAYHKgJ/UwPzaaey8lQ
c1BilRSJf993lzrnrZoPBK8QuMiSyGj6dOa29rjkyrDxdJwHHKEl0Anjsv1qIDDU
uYI/C6FhEv3W6srU8JAkQJPyE+R+F5E82GWKEJq5vlOr6LNJZa/e5hvlpbRLDCUY
nVcFfVesKKgegeUOGcFDC2CFKZZnMnsFqdj5uFducUm1nJSeaK0zoyy5fA9yqj+G
7DRliJ0PW8Ybx8nayecn8QQL3QsCZQAs+clmsN7MGHmCil9LGgGhj+bUK2BTjxHV
cFj0Re7uLfqw6yd7bkt0CjcywoZ61SKviY1klUHznHchwYNGPCMPZArR+U3Cnnzw
sKiiEVSQAf1u0Rkjq2cQmfeG/iTo/hRqjwDhtGfWgNRG2QvMd8Xu65u7Wnsk3S6y
uetS7kgmbRaMya1WEkJuxg/FCBVYhCTYksXo+w/rxtftUG8E04ss1XpYkMjLehpB
8AWIDkvxHoNF5tIYMsXdGDXIpS2ORRJ5jUaLUbTttwhDiq+EGjjL/ct6WfYvzCSu
5LXt/oHHE+A46CXR2xocZ4l51EUolLCeVsGVVwx5RY6b/emf5kZgHBoWO9sJzYj9
OkGjP4688aBIC+seFB8xwaR3jD5uLkKXlvygI0g1wEF7LKTv3OMNxleHJNl+6/8P
6u0ZyQfWMisY9LlNItnXvmf1GyZBzdCl5ZYcgAuJsQulDmQuaK3zaUO9DhgUEXLp
vW0SNfYWoJboLkguQ9NAFBoZhAA9XS9b4Z6FGKwdyJv08Esn7se822iQtDhNTsD3
IWmQ8NmMEXN4cWMTJYtNV3eh/1HYGVi3/uFG91NxA31IKfMDHXU+tmNEZkGLGtZZ
twtfACD8XWrHMHZM1k3CsQA0ICqWZ/Cv4Xts0yLwptqbRREM/VYis0NnMsuckU4I
xltPCMtExL+2Ndnr/Vp2MRanxR/Dmxqftip07O3VH4JBfR9nHT5qJdCh8gQ0V8LI
VGGRWxdip+V0D0okSuFNL8lqs+GMFDZIJvTEcZ/PknldZ1yp55RItJX3GMoGFFw6
12XEAgHunwNRqv2qVGlMe0Nn0xG3zpCoy72T4H8j7xg1mKQPGZ9U1j8//ijWMmm5
WQtZ87LHtGrB2kJ3TR1VR1X1gFCtFhCnKN/dk2SpmFkU1dBoivBhEz2Kkr6Baxrv
lmXrauzITOl9PhjlbgLk3PljE49dMXe13oXUzhO1g888ujaevz1uQG7TXfsYh5iA
kXoTz7R3jEEYqPVhX+fPeM5F4PcMcNCRw6icoypHrU8Yd9pgnBGklmSM0a35Ul4Q
f/fI2kR+3/36PHD6fVEAEBikfhnnwCBoyYtmShc+xSLaeSi3NO0J7xn5dzi+ESkb
0bn2pvxdiT4plpoSuyasE/NcIoXv6aD43aT4BUhF/DRCA4dc0zHim62RBfuob4Q1
2kKfL4o/ij/WSVYeB4iiJT86MK7YpIf08tfIjtRoecXGKHZrY+UhHzkamSmVnMjA
T4X2l+g6MfSA+WdEHMfuZLQzd1g38mxFvHczWhNkb8HGLfW5FUbVwoXyOCtb6J7e
kx7zCOZlfRQY107qV3e2ycIheeIuEFw2sPA2t6SQ0yC1r/JqZxECYtH6I8u0+wN1
pgXdp1wVz30lNJEwFrZ/YHegKr8F02aZa8JZvJfdXz8ccZbloaVDcon5h7a529Im
CRoMaqm5VRZSzBIlK92/+bnsdlfgq+2e/1SkV9EdBw7gopL3hqTU3xvk+/SbIN1v
9HZffoeSt81PnzPxtGhGi9XvYmjOYvmA7xdyrM9eGotA6vLK/L49Lr9b0vgVaigG
2AMPURHk3MK5mFNJ6hBHn7fRY2XNkjgd7EvZlv8njnHoMhYUAu8HSIz8R1AHNP0U
GbRLOgRPRCSv37m9s3mfnkdfUVJ/4/ItUb2uCHuRfodGGPRSf2EYKYTD+h46Egqq
O5I0toGnpBDUCl5eBiL9nx/gSkrzOiV0oMs4avjsCCr6aCyO6TnLNEwzG0Zvf2co
/tx42sGlh9qvO3aJ9J2EubiWszfWY0t183Ltt2RNVRcboyb/TCmg5AtDDJJANlAt
wadEl0UYbWwdvghOtL/CyYPrJsCKrVaWXnENWtFt9ZmmOBq23UQKsgLamdKyclUX
xivmlsFKPwl0ynvUQIOnVxXaR6AY1D+4BOGm3WcpiCb93iVLWKk5NTY4xi+tQIQO
YkGVMKBmYptMOQQJTynaJ5IpEXgJRRPtGYHjZtkfb1BhBM2LizuBsGXls9p5iN1S
Ia5avBFq7CCKs5S1J/eQ2YSfMkRFT7UhhyFRSTkdyPQX7seykdzbgnI3oe3X86u7
eqw6lyAZoi/gKxLlbeMZc3lkcQ2LIsIvYNTWnnXt+do/TFnR0dbg0N9V2H7VLev8
wXhHDwvHAa/22o9WfaO3ESqiRZ0MCWdAR/ccyT1NGfqtHMTtMFuF3jWpz0DShC9T
XzS9hHE7jI0aTUPZFe6AOze8eekRZTgso5AZHpcdDgWtbBVWxHRg4KZ8kcd5O8St
nv3bOuOUsrfzIxA0wb98nT+MpUvi8/T916RwTjc7relduiFRU+Ga010oURGYQQE7
0aWl0lZthFA8N6a6XlXoZXv8mruub4oCzWkVBY8qUerrteCNkmaJ7lWSI8zRH9DS
N7DSdxTu+08FbsuC3KZZQKji7cTFqixAp2WDzoGcZZcUH9WNOwFWXOrL5ifaBHh7
F8ePyOBkbFpNSrY/WzOi9dc9I395a93Y66dLFLKGYahfsgpv4+bemN3yJWwF007h
yzfyN5HfYKmCCfEgKsC1turzB5NqeXOL2L5rRGMjcha8RM87oCKKOtDDmTP4kgZd
xRRTwe+tLFAYmi/aIdMR5y31DSgy9Z62xL7LYwX+qCnE/6zvjk8aBxhBCjPIuLy8
TPcvgsrfbqNtP8km/N8UXI69zirMBx8MM50cGbO/BJxNsSfdtkH3xxUv/lYjddcV
vdRIRz/E+LnhaKskCpIiheWzbkoz//be/r3BEpE0IdM86jss53jkPOO9gEkT4gyV
704Dkgiu8o4sUqmWyE4dIfiaFIoiqGQkN/bdhdgNe9PVafso20pvNiz9pSvFttRF
7OBwnu7kcrbRQLs7tTka7svXCmFGgytw9LkEsOpdr/fd6LJYIqtDnhQi2Jy0tlrs
IyMgZrcPNBdwPCf6ZRHsSJ/AF/jYz6DA0Jqr07CquKdrCY9ihM8MmpICLOvHuLeB
1PTbNJIMMqKwOK600YjZsKVPRNjwBfWFphmooZpO9f3hezz2GzgJ6FD1hOuo/prV
GebwVn3exnd3YuiU+Q+npOY75TSn6HIznieFCGRkme10lEJWUm2BqyC/5QZLrBD9
4UJxClOhaCF//rp7nxlg9Z0LmH+sLRDkIa7a4fKNlqCEMVSQo4xbo2/Wo+W3it6Z
9p1OnPjosy4NxiX6koEfzvFCgICBm/kH4jC8vnRD9xDT6OGnjmpHwFClQfGHyQsp
bn288BEhbAw6Wk1/DlOGOg/2qkK5H3L/ZuwSZg3+r5qm2rTJ6l80ubcoo2RC6AMq
M/huV9S57+QzbPl0IwXmoprpX6ozJICN18qvpfrMPWCFZPafjueSHaBEUF8OQhxO
i1KLUMeTiKUo57MELgQRvNZNhSLVK+Z1q+4svCXiKz0aH580YB6gK6Bo3w1HIbAd
i51BjzUDmtWqNFYhBvi2CqprSweMFC1TNCjhknhngrcqkpzL60MlXAEdjoUoYfG3
hySqos8DbB1s5cM4FxM8OE0p4/zh8v4v89NM3JydcEgC0u3obYv0ZhUDb/6+2LgG
AG3rHZORYqh5EGTpfH8wF588jEzm17YvoT63ZZlr5MryyrWcRf3x8FEkjUZmEJ63
qw73unJlZRyFvcrZI4kmJpxV4uOYD1XYDU1N3e/ayg9kTuLP3EqmRZiSYGVXOiP2
3IaCKXhzKmbkjVBgOiA2m1xK7XgJ4xz4ZWGobAWq6S3EBSkEgyBDHjRGncpuVRTj
TcjXF8MEcake740vDc4p8rGGB2d9eYtcPHMLNHo94dkjwvF7erQH32YLAy0Tplf2
kspOfkEtkZkFx5X7Jw2grE8UHpPTh58h1dXhAyKnJy93AvcZb9HI8pM97omCuFdb
1NJGF+IvWgpdiQipygPZgWsdefPnqnghVWHO7fQ5GvV5MAiCIQufbcbfd3wdM0Ei
6fjfNDJWW6SC7oegwKlJHWBK/h/MRfpiivXZZXItomnnm9eoos7Tic8HJHEQLrpZ
OEd0eJC/i8b97U+WlIQ9hhLn1pY8HuclwTw6DHtO0zAUMaSvt1mL7DfHQ/g/nFMc
vB9o8yLcqWE3UuqKD7rB0Y3jZnAKPFCzgjTsqt7F00TopHP2UhvvPaiAYG8W2IWk
Qh0QQLV1mZjysC67OO9Dqg6tjjnAay7u63e8i3LO49AX4irB6LHKgZj6VIKEm3bq
dkym1pMb6j9s7e1bFoUdQnMvrDOEwM5yPoRTx8GqevQpZgD/2KpsmsHreFXwlS0x
Y2nsSVBQDcGCSMOlvx6z6Q5dRk+nbFhNciW+jSV+6mE1Y3ABBd1h3zZpjiLJ272W
E71ir0Z6v6gDVRRKs6w16BZ5NAGXd0D4DydD/BRPvd4OCuXUzG/3m1fdsHxwoALO
wh8+ZT3fKvVdVi2yDrJpY5rnIUhWepzdY+6LfBGY8A5AjqQ/bJE9JIkHiHFfotN4
iiCrUMqK33uFg39za6jeEg8Uxsbm03iM63hCV5tj8BxQzM5/NpiXLHid2Ra7bBIk
qtQndE7ZFPJNaq+yCWUu/hInOo/1sFN4MM5jEHYBybOxV7bTmF/zbdYTgXAERW/4
CfCCAFwyt5jSHBOaJNyTNY55DScZswFoYKP+7Cjp2hAEGo4MaBzSkscUBKXbXyUx
0FPsTzZvKI9YJZiax3VbJXFmmLNMJQ9xE5mNOLJBSKDrKs31RnwCBnYRtOrUiq0t
iIt+0Y9QqhRgxf2by+wpUyW1MSASxzzfb6Z0bCWMdbmiwqEr2UDztlAWj/ogujdB
ylhYwvw9GNaQPg1GW7hIBb7hKO/41Xe7sBHUGfGx2G9wnFECWbrzP8vr40UwJnJ/
fQDZ+VTc8HOZL+RHaJ6gOTt4czmUFJqa9LMT7I7bxMNu/95n4nvhruyvi0f+S/nD
OVc0l02vS7BGEKe7VwdQXLkyuKwcNyKMPNFwHsxr7IprMHeknHTWsr5K+71m8uyw
5rdY0CKWGzMlk9y2Nq4i3xhoFiwVLYurzryscZg8vjNBe/tZAu5p8v4IQeXSR/Xy
4dbTRYBHAT5DagQzI1Z+grelgm8p5Cxwo78/RqJdvuGajFvSjPzD+cGUVztEYhqx
RE+O3fbsmuAoIMTObHuS/LwH06RIirt21PqOyx+tOlNudhkYXciG1F39JVTYbYJc
iTJh5LENibi3CqREC0OJfL9NPqLQTJ/rOB2QKnSaVv9WSrgOymswKTUlsjC4Ze2b
jWR9DmrM7a5TI40hsirO98JrmXhuG3js5ILWbzVKz0b7gAOvcSvG6jAmC9Rciwtq
agzefM4TzQm5AsnliaC+voiEK4WZqBWdrTHW8as2SVA80LohJ1nSu5jtcT0p1GKi
5IExJlvDtCu4pFH+LLyPO7/tz8eMTbz81si1QObXkZFXfAUQqI0qYvwIISnqQa0W
1A5CySICBMdmf4s+aEGGMWWG/SBbJs5aSkg+5bR49/7NFTqjcw/0cmqXgjslOF7k
Zeby8SKcq05oqfMsAyWZ/pAW0JJ04nM1f615AMF7CwNTLYBNL8tVxGx7hSluuoSO
Lrhc3M3j6VSV0yT9VWFDAuPR10/6xSmQWEX7lzivjDSJEw4AFxADd8P44PEDDhX3
afbcpR+ID3ThjntVXOhyzlyKrwkLEV+rYtVLqbo6FYIQnRMlJgNJlhs08BkBuaMP
on0DrcYwuDtxKgu065791y4ghcps6kkyc97b3qskafkpFhR3tbYRp5Vq++td64TY
V5ze2WkSfUlfaOeDpErw3l7novkgXzcQ/6pGaHd4cFt1oqiDBNx3u6A0CUkvyOjA
yrjI+qgSOuGc9v6f1PuZptobeKPN52Jay8hWbE8UDZUAQ8FXp8xVZnhfsz1W6wyc
CKl5BOtTy0/L5JOdCXDlS9ZIKCyvpysQOdlx9pS+VytL3xbGeCAxXzwnBlptSe6B
6yzWu3unkkdV399+7WSImgzAJbl/DY6GmIzt/VSfQRBuQU06XJQbP63V9HoMy+mn
jdzcSvx6NtYwRIDl7nxwo5/rTWHk9reGSGpYdwpKGuicaYHqnjYJidddss51VAZk
cUzuGIUHCEJnOLgqV0y0iAXwfLG2UU9+FZGbZvEY6lMkCCJGUdMuVYAeqz0XkICk
E/LD0QLJh8wqp8K4m1lCsqjaKITcmyZ16CtJ8AfG5YpSDKyimpskIr1OltROKap6
Lu5uPlPjTWZeDeZdS92Dfj/46949YmYr6tDim5wNDW3dvTSOovoOyNoQeF9yc7eA
QQT6HKCrMf+5QXNgpQtXjDImaT1f7uSGTRbx8SXJdUJPBxCpp4UAooNa784QaJ0N
wBFFxYmHvq48eXfp01n6zk+YHIKj4Qiav6zJ/+cbd29qSJWkBxXrfXoPSd+X5BLw
XFZafoV6qzIyOFYcQyi0BofPrFq1qnIpl2dnhyJ2J1+JPtPuPicFR+lgwukB4hTx
1ttw40A2fZb/m0J7hkNQWHDof+SnU8EJ29PUYDPj5cm/+e4XgptbVNDU6tKTYmbh
YZoQ0w1gLTKhoIoXg1ebLmO03ncvmaMLxZ2uMVta+HKKGSJzlO5e5mI20aA5PUuA
nr4ygqdmTIJeJqaZWgcXSzcIawHK0VMcFsFhXHdIPOrk8MRztpHYW017nzzF8CKT
BjSCYIvoLJ/CleZ7CTUoO3xBvUsi3FpV11AsDDCq1/junXYZfwLlvGqk2WFt5cvm
K1qWfxihVqcq7x4SNzyqs6Shoygobiw1C0HDf4BIEAqRzAb75ZmfGH9xrN6HDjc6
R3DIC19wpk822fdbdH26DfbXjj6GfxBjdKNZSsxqV/pZ1Q+iWofjw/SoJqA6I2Mn
ObS0Ab6LxSGCBxjHMnl9QckMqebPNgHRyLyEmsbnbYF8/xj0NSIJ63PqaccyEqAA
uZgZnLatMIeJ0a0fzBDewfpQtk1IRTUhBhXyPi9o5BmX2Pdij1HXM0xSiDkro9Zl
RFWH0SCAqYC1l6xH2EFxJWxw7VMQm/bvq8Coogb2m1bysHrwqFwSr7SMWPUhIwnA
d0OjWDucyaWDZPYwqbFyPh7A1zPuXKUw5uLQm9ARIyAxBlbTKp3CUWe3v0wLsQMk
C6Ic8S1Fm2lHF0ajGIaZqMTh3AMBZiZ3wLin0EGFohV6fsvZMCFTb5MuDRUcWmfL
DlkyjARTBxm/QFxzhDXml5ObjXKEYH53yi86S5iEDyju18bJ7H2n49AOE8yKaWay
cQO6ZASpMLbvWb2swFTBb4k6whFFdlaiQNLOvNw+hMzWnHuCqlUUECPEkxIlwIHv
cfz9cqQDo3/L4lynnwv98ZMBm65pf01PbpmJEvtQuJZF7tm3o/7CjI2NcWO+PUNU
7DmZo5IqwqJsn/fGq8Bt1hTo2qXfBNbZ2tjyU5RYBq28WKMEMCUlbklo5YirKkv5
Ovc2k+DJ/LfYhtkkQA2r6BEZ0FUuw4ps3zJ/2tQ3oeD3EmN3X1lplBmev7wB6Yaj
9sp0LgFfHLGWXzFT81rE7L6+oeRWNpV8O6U2ltZfuA82R9DMCNXAtnn+/ZdMx+Yz
wON0UYYAG90u2fcJwTdQXx1AMOCScOXaQRv8icgFUv922YBIL0TOf7iO7mexPUvL
MYwG8X9NtObDlrNCRi4B+2ywgTSwY+XbQ7admI4EOwp8xYj7rEKSpMQ8apvEHwsc
Jj6hK/jutff6gp3ZLKxN7BraG3+H3cIKq9ZuXS1wN24bWxqTern0Z+dyZcC5Sa+q
IKkMvJJXq69Btk5nPiiXtnfvbLXy28cQg11z50YopN9oQFWLfJ3PkDtHkF7G/k8N
yukQ3bqshcIE02PRCrFfZwJS/ANvTeBUYsmj4sIZ0+b5tmPSqRCIg8G8nDpYPbTz
ErleoFqliCRtfduET8uDdBPKbdEwPmXevZyom826wkPtei4Vo1treDE0xqEzV4+F
KXC3NSSksIohs1OyZ5/xMTZpDpmp19p3C71RvFVMfIjye8OehKQEaykXVpSrFL0x
AfoHiQDJWxsU0VNcgM7KVIZx1RHyyCbArCTJ3V2kbdp3BktV9/lveZ6u0GbsUKJ2
tQJUPGWUoXAeo4368t1BxNkMFS9TyMpmjq3kCg+Ye9v27IZKH9mP14xDVUs+OLfg
0ICFHfR/vs8+kagPLE/YD8Qb3G1rfVHVeg84qnvpfsWucKf2daSVFRrH5WXlpm86
KI+JwCZPeif2RxLKyunune300f8kgREMoH9EqvBopS5LNXhUq3qPvUiCcJ28vCWc
kSAGoiyQAOKAoWRXi0SyLaXvFdNuU3P4GfpLwW1nTaxvuBN5dM3Xbrv42Zb14PtU
TxaFd/2LC9GLxOEiMF4T4D4/OBrsJ7N4UWyM3dtndvW9MmJvfZQ5mYfIJOlMzcor
uXAbuOVc5n2fNuyRKc5gCzQReGvZ6yf2VmmfsvAgDXYR+ImTeXGMHklN6v3vatto
0Pe3aPLm6h8g90y6DJUmgnljA3H8Qx7BsP/pdy1SU+YypQtb2JqtfQ3F7XCNJrum
GaPnTrJoVSHP3HHZ8J5nz6WT/nsN0sYMghmws66RueeT9gApWd3IaqMWWut6bUB4
Q1do9FihYKLv1Rx+m4/a/TsQdF6Q/nVTFZdkRAvrA7kmNjAVe9rEG00VUWNZz3ev
UqddHYTXmVG+yc2djW/Ws+OHAnxKYoxS6RluvzkN4d0fVawjIJlUjjMjsJwSaO7O
S6BLU1GV6sZAt80s20YvI1cvEimbTcyfML1tANrz+sBIuo1LOg+jTmRigFNzbDSE
3Oe8wv+DSvOz9vnkHLz4ltxCBAeks3g2a2zm+T6p5/fLbp2fNbjWKOL1/c8+KHLh
ltEahaL3pOImxTATPiSrhuvzCrTyxlWt0L3D0NnHokLM8MvhfmYa2jmwoV0kzyJl
XynZQlMv7dgvjkXmGd36ssVG8DMBSV8Yc5c07JRG8Vlk1uGO8J6FOKZsW/WHQwuH
9/+frG3kyPfUy332nBBYZmVeRvKVAvPE4FRhvuF0j1WGuiio6P8PsIUdlIyoiCdg
xjpmg8RXiVx+JXX7TzO4cEDoQglk4Ct5qK3sR70zxPnO5Y2nqDV/IQH9zsNK3WT2
bPZ0ht2rVcKcswogGUtO9NJ5gtRs8rCpm3E82S0qwhfpKyFF51qFhmby3X9y/lx2
mqAPadG1IvieGYKjr35irB7CTPaFaMtQE5yqpVuOF4R/8p3FVCznWyeFN1iM69Hh
wyOY5GH9eIFAE5BpjwQJvBwoPSjSREyb8bNHUihtYYvtRJVtX0OLKxSZudWgEgeM
OL6ObJ+6UtT4YGZrPvgQKXCoP6+ZUBKaYnxHlNm1xs0MSkLWZauNrG6AVkPdXLW6
JOwfLnJ2/iNopAP/oOSrQHzUKD+aWNazpDabMZlxYaGmkDmdcp3ooVmndIVTig+C
C88nwuBMb7s+Z9AyipINcYqhJYJWNlmUL9y3BMlTUGz1KIEC774fcpSpu01Lo/2S
kysOjqbwsnBIBmx0pVSFOCtx/NRFQglR3sT8DCQkXIVWhkglTTsKiWbT3xVJkvM/
kxGNOa98HQsrvUfyuxZDJsPbeGlQTafLywxQwK6Lm8UkzxFPl6RqgzSoKUzD/muj
/4MzQXoa3/zfahUdOSjWAsPwKeJIdhjYzU88BG/lmD46uls3M4yCVOhI/gZXIEZA
Gdz/SYH9W54XnX96yuqk36dYp05dTjzOQ//8GMGGN99paJVraJ2eYfEt2JajDd2N
WeDuDsnNCLculxmnXj9m/vtrZTwTflr/04vRGF6UMHW+QxNouWZ22TkhZEIHQZ2N
81egU2sxw+oGsM3bMdnzGqgH8tJGSn3V06aLAdX/Ma7rMs3Q6hqq+P1CC8EoBUim
cXccv9JxOffCTgZ8kg4QnleE1yFjHg31DsU3B5vC0htzPvh7o5V+E4megN96s2e5
j/DaQXN9BZQtKAOrRaeF5UDB0q1XAyNmV1hCl4NgdHu99k1CdiuFaERbr7GWKf+b
Wj33bElP6ojf/9hcYAABAVKVg5cAwDozubTYBjHLNCOGNO9V/6y2K4kWU2D1Jxt9
7aUq85kgkHox2r5/YHFXC//yo0xS9J9KZiYmRtInYQDFr6+BvqEYVAvHdVXduiWV
tj5QaOUDAhPlb4bhtF4Q1u+BGvDK8hsyNl+YRVusBWh0dfsXNT+YMzfvsJCpDQkC
rzkRwD1iPNC0zUcnxdYS3FcKR8icm6Zbiw8/5hriDsGYY4bZPFGDJkeKCfrZzIxE
SWrPutzBPwPhijxHMHNcJnqdF+twnaoWUTMIGYjFmKZOBi/dMWnO3tACo4mdVKlI
ZgOFYJ8If0n/mikUdsmpG5Ob8ErvtLNRCXwljhvjtYKuiLbUfNALnKHilpzwAaLW
Qtzg2hz8Scrrblro1QMbrOjCZtLNv23YS4ha4gzvnXaYsGFOhJeFO881aQpXqXtM
cXRSy4CrUn0Ky7DElPDJv107xY0LWxv9DC//MqQQhzgGT5K7eMPf+JakT800IQN2
MPLXmSJdvltydecRbAtAnuZOID4NoZ6XuH6TjXLP1Lqob1m4Khn/9qErieI9oHnB
HyQuFKaeipkhaA5v3KwzC9nh2qwVqoJoTK7cnKPZDObq6RUPpVGC2mcyA/bGn/ZX
3kIhzFF66mDG1RPZX6aHE6GXf7cmjJ5n5Zx+KDKxcqgDky0N/2p3+id7Osx8/xXa
CrSxX6mhTDmOmZli9Iv75Xd0Yuns8c/LTSZmVYf+EW9H1HBE4+83hsa3HZIHlEkh
Ytcu8t8A/l/FlFoDP4zwPZcC8OsTFa62PyOkW3wQ+HfPVpRvPsaF2mrHJjmrdK0P
RmqtLqMsF5Zx8xeWMdE9ZCEQR1lNOVcMULciNHfGLMBqcGTrOdyVBOo2SsfcdvZh
6kEPS16Ij2sClMtFVOTELNZpwwopWA+XFVguUdngdgj4nz7H0rFNboI66pbYW6W+
bulna4G1jTwze4Iicva/hzPRzVsDtUH7wiBz3eMHBDH4YPvQjy+c6nOzxBwXDCZr
47FmLuxoEpw4LpK+5ipUqBJIDPP8eMPn+b2bq2c+m22CJwTafnROsCcZiCZgRNrf
tRbinB5vmKxUv3lsTeYadVdIk1SairAdPQq6VCcBllO0CGZ+e76Omf90x5ZjUvHr
1tgHsf/mShGeKdtcNtz7chxSzkCLR6hriMrZSHLT256agBguAJF4nS20A/SK14c+
9LkvXz9vcid3aXYa1NsXeDE2KKEUabvqU3Iaf4YRtuQ+7lpSYiCb0ShlmFbtTTMA
CeTqxFY+B8Z9F9iTAgBUOmxF1GpCzfpzCds2Nkt4oLZwmOd64HraPbRoewmHKhQV
+7b0VY0lG2g8+4uRUAQ//6elGYzXgM0uVW5BND3wF3NTzpCcvqSrfRanOnxPy0WV
iJ5kPaONuwakXiWzU/QZDQzLrpi0owx8YtPur4uPTR2dcu1RHcgOIYNKm51uNTkO
HZ9VmUXALyC0Tx8OOrxLpc2KDydnVP9ittrgzhgnM22Z2fLeXsWaAhD1gom7IHaa
Owxi8PP2Du4MNLauERuS7i4BJFpED+BrfydblH8pExqWDkL3ywBw7VU6uXbHeAha
xpRiDbvyfH34+TCnqjCGgumCzTTEkMZVFUhHUCd6GqMwpwau8DFhNL/HnJ2PC5Yh
WTXT12lbDcWZ/f+JxxJO+oixgcU3BymqA4wDsqF4GWHqivXLNFOFXoCGmX7qspZJ
CdGywJQzsjw/15LYNPvAlYNF6zJnrJLXKF3KsU0UJ31xKoZkz7fdlZl4OcEkUVzi
6W6POF1JiW8OixHO8z7mD1MmfzVo1ZcbLuBFjU9si36jHpCT1Oja3rgqA1GKG9cH
TELPjaVddy/lVVx0SQz0FlFQI3/3b8LYIlAgsYSf3syesv/etHZcN5CgIu4yeDrV
UABXEVuG1Xf09WGqhIfNREc5Hnh9C8hKdKhLgGyURwqBdtffr+2VSsPbp1SORGjk
quSKNH9KrMqukb0MhK6xv3YD9G1Ep/v/1bciF5qmGFDofribamK5yqI6pW6HvD6Y
R9rzmzX9STUaFZ6ONDaGk0E1WZ7JJZgsubLRLzsPnoe2h3wCuXlKM001/7DqZQ82
qW7Hz/BF/aMEBOLLyr+d8vlQ5BFGEF0M5OUIffkNVkrwBhsY5C8XCtSMk1bMEW2Y
cMEj0R+HxsGcm8BsGEy9qCTqknAQfdCSZ7tVgCBkkaS639whyQ7zxAA83Xa0yHgg
O2rScl2j9o80Za2JRDeMAj9uiaTa1meDU2wVzjlsoFCpZfGn7sL0yu3UP81gxTCp
/rpy5fB9b/ZiZ8SdoqoQVC0gatyB3bB0PTieF/uVGyJD3Vbaz7S/pIoivGNNCnOK
OjUfD9parZlwQ9+VJ8PNbBYx1BcIwvyyKQNRhiJL7p1EngKhUd2UxxyGZH8a3rtz
ttGPt5QeyFpt2My54uC2Bf0KervvZHOiGkS26Iw2QDLPOuymccfBF/uRtRmcMHPK
fYicGwK+f2qpwzA3jxmoi5gKqM4jToIFGzC43lPXCxLveSFrZ11GN3HKG1uNBTA8
O4daqHNTbc9GoYMHNqIVznEVRl054UuGYxJ6g5DkoVOCOL/ONhsPUB/VhWvESDU2
UgDqykNyoi9juus0CVFiy6KyzaBvW8IQOZRnPlbt2ybSqZfpn57w86svtKdIsc70
QGZsiUCvdeKChi9X0mvb5Zj3Ux25xN3EnbedgyBDQXUt9n2uZENTz7SJpwD8G3dY
ITMPxFZX1yzX7f3JYqmw4pF6RcUDJ5NtJZnNo1iNwyvikVvdP+K0jJkSe13UztFE
4Q+Hsg9R4uR6klmMfzY1I+WKmXn2HMKd1izN6ylc1foP11xlJtXhK433H1vAIHqq
xvhd3Iv6yzAEWJeWob/kQOFmsjlRkgz1YtG32VrGt4fEe6E8K88bBeLFqNS55Up7
z1y0a7FPic5IesAhRVcZZfY4DNs2mds75zbFKAfBZyGbI+n2sntZiSrafTbTqgy2
bRPvNeew28NNHssCiUh+l3E9FKmgTuL6kYHRJ0gET+GeE2CxcEUils0SfTgjDTq4
EfVQiwalC8WrBqv4gDbnJ7u9chK+RcPPTKSPuzb6EGMxwnXafcu0oqN7Fo25m1UL
vMLE0lJWMfwgiUPBs7YP4Qq7pg5vEdlwEJPKUWUrrR/RJRtOU5ztr7UxGUi1oZ7B
DfqRWNdcr55+Zv1t2LYWlitvdrmqfRoyxu15UazVYatbiE24dWtE1EJDZObQjeop
Sr2zSaEK7CeG4otPW6hwFx3SiD5a0jLw32XMkRQO8osn+/xhfcUSfUmOlAgvVe1j
hCM4+351q1uZiiVqxHROcb3wq3cm+HKyPAerSNeVEoKINteFLlWcyEzJ2LLxcDuY
WVaLwrPHosDFcnSOmjf2eHK6ihydiOOYeHPV65oLEKQsGDjwQVRviJGXs+mkbzrq
lfVs2GY8M7FNjEdSJDe2LyHHjfn/RpdwacuU7aENrU7sFyI4sNyIIFuWF0Klxz5l
eE3CuCRyfUx06fe11DHPkQzd0U7cFN+uHbhF5++fzvM9zMcYpAvlnBEax2UUAu+Z
TGT3JOg3KwRPxhPYUmkoBHV+fIuWTySHnAGhoXUyQKda1dYjLXi5I9EqEKVbPC+u
T3FQ7tQt72aVS1znXe52fpJMIvEW8Sn33S1I4XGLdYtA8MJ4IUnyhG3D4lBQrom4
0OTt+/ylSsZ/pjPtnfDEgj6dJu+YyaX6USMDWFeg/ovhnONBr3IptO/sufKEUaAM
sxYzW5nro1SB4cu4fWQuzV1loC0wf6RhtU2uIU29k4Bg+W9VceqOqajkAW7LgFYm
rEL23Hc53fhGVzIVHBlk7rLWXxlY7NPOgIzONUz5MGxIgKSF6iSlUe5fI0N5GcAr
4Ho5XQlCg/RRAgc2MoS7OMM+ylzD1f3EJwnTN5Sx9nEztlGC8h+gLLIwl8OsQLAt
aaJxLuO1m/GEvuiz3QzLpVQJFDxR+NRjjxRIELnBXlyQP4PRkK/lwNhWxiaELuYW
h1N9WVNPjyjnSvrucHpi1vGMY4ANk3lVZRmYGg/6avfwctMi2XfXvMimo58HS4a/
ooym/wo62TYH/29FHOX5BX8BSU0zjEO88hTEPliThrjHVPeXqTAmyT2o4BmVtV1G
nrSSybmn2PRg/1PpJChhXOkdwSgrWHjevbNzQrB6zRmQkEQ+rBSQv7xjzvJ6kOc6
rXACczjJW8YGAUXabFhg7kLOFxxMfIiGA8yFT679R3TIWWAgl5BBXJTw+QxfHvUq
/vfB06P8em9YR7Aok5er7t+lVoCqMLckEZNsvl1/vE3bJevHC1rAzp7Gz+KDl2KN
IQPY115YUvDW7H2OSI2UNfpaPVKiHs7DFEnog265NshX89Se8q6oLY01WEJ4zTai
bRDaWxSDK7+HGbYhvQfN9WZz74glBGMGMGLTvfAgEMTldmF/8kCH/JYQywDAQORF
JZYHpOY4bPmI6Gk7CpF4rQuXy69bCUhvTENzRWyUSKVJ1WfEpQEs38DpW3ooLPQZ
kvg+LilCTkjKDnZPic41tuaTDk4y3+knGPAORmOZgYNnEFPslhqgR+dxv/c/huZS
ISYQnXXYOTpYR6FZKyq9VqA0u2Cek8P1GcBTYcm8agsL82hOGV3r4Y/mr0Py/mQa
INzcxjgTbaHI72V1rQSN2sK409IiF8L0SYAIrll1yujptoWK9fRwwGo/6513JHfB
d8jmG1i63PW3hQdXDfepQDOnXBTOCYAjBbCvLL4/iE+yTrGQLXs1AyJVs/leF+o5
tdCRnWVYkIo6CCGzGDdtu5aZItN5nTpOWxgIilePfqhqFLy0a7+yriWNUfypyitv
+8BmlCK/brddKgEM79dY3K2ub3pZKZ0i7Cb3S6gDbppOeo+uFhDk8utZ1MfaU4lc
pmtl+L0dKiFqvfR8HVhDVDJpCxQnIYZnhGyvt4nUBH+6owaXZLkP5AE016Cq2kHL
O6nw7fIrPgZU86HLXzyoPBU418BX9o31ENI6JVjq+qGqs1bENpTnNACtGSzcCna7
QN21d2kMciOr6QuPCmaq2HnstBtFyIruAw6XzZebDSiwVW9tIihde87n9V/dmEsI
wZ0KV13oIn5dbNMeqRjBdKSP3funXxf8AZM5EQSFqHr4WNtN3Lbrt4mtupEhALFo
aVtYxaBiQ9C9Il43z0OsQe0d7bHlCYiGgaazmMf/qM/24ZDWJp+ll81hmBqzRWH1
ERPCvpf2K4WlZ/EEPdHZ8IzhAGQtqUk72RCMofPOGbe/tzSDpvnOhFaNH9ESmTXH
yrKEQwlMc73LmX09ufhlAgSpcBV5uqMwiUhhN+h+9cF3NQlS/V1zB9LCTRkRXK3S
6iw2SSu3FzikxbTo65ia328SMCVxPutofOsMaDdfNhMTpO4rpeO5SlhMJJEYTGgg
GK5+IKxztUICRXsQYzbBhneaJTomDtvzaVkCHvWqJFc4FhanlXHQe00gPPzVQRV1
tZsfT+Q73NwpvWhmCGMJnKxBfCkLrzVfMXKUQj7Fmo8CRD7ANe6x2C3LrlvMNIkK
wuKgbL/Er0+q3QjAHX1gk2DKHyFNMz8McCy1G5ZcDpo9h4wZcoHvigQZNzVWpRdP
YTWGhELLspi0B+kcRtmNtVnia7n3YuThSSjjqKpREPExg8BzBlR3wx7PqZIWo8Zb
+X4n+ZezBLTbh2YjbDPgUujbFI7PGEs9rKl8FymAUAEIC26PpG2Mzb5cXQYfQSrO
btLBjkGEU2iNPDbqAtgjvUI3pNLWT9atxE1hX1j8kUKg2Fiexdq3LfqhEiNI8yU9
Fb1bITxZi4hiozz4CMrG3OkRZHh3TpyctE9xPw3qRw3pRztJ3YkDaF2ZuoGTdvUe
kNjdYMcwNacZWHgi6+u0BDxgnbDNtmLi6X54/6jbfdEGV59x0w2lFifim5nlxcqN
PzKbGcVhu0fNebkCAeZ9RrUf5BnpH9y9nmfPeUqDnUcEhKHraXiMyAUzE4r3wRpS
2/XiJDhrIWdVtwGjQs+25u5acacgkhzzikF5alzvnII3juPje9TnEwWz/SjaFX5f
girjq0wig+pXJ/owA/WqeSRpthlt8Fur5Ya8tD8oesk+0NSJT4T56Gl8pSX8wwbg
QqryjorxBHOpsc9SjiP3cB7h15H5BwkfR7HtnYbKWzPIKTuIygWosggXkCDiT3jq
MkihvrbZegvoQGktP3rT3cxWDPt4obQ0EVGARIFi35pBp4byqKqqyfLN3qcmd4iZ
ZiUh2eutuzSbTHQl/GHFOjdNNKdtZEbr01OuJIrw4Bjtk+yEmfsCWcnZsSS56aUD
s27aXa6mU5spggp9jQ2CZ0DquXx0WONJnfTlNVEMcWhRaNTmABOLJOttmthNghkG
Mv9uHuuWIQQ7VJ5RdtOesflhddc7w3e1zxjSwvZ8WN07LAQpSrC57XbEjVM5DFEY
9VoQbbVziOysZXAHERNEnR0taD8VyHSMHRIny1rLYL4ydoorpPRENz+M1iDBOJto
UPKyoQ5cQX/0vjNhmcTQpERN7Z3bR8hnfqOv+D/d9ziNJEzhh4p6qxD9PovG43Ni
jURQr9ika9Rxb0fIfQILWAbYtL1TOQgcuk1cXECkgKc2n3nHM4KqbKWfd//6JIo8
xkcfMH8gKc5XqnbS58U5BR/RqUcWDaiodI5Tj3cDIc3ngVFI0ODhIojSyKbelKs3
DQBUfe1QrJe55gwH3CrKcu17PiH0IIfwEtbpzGfrA8ZcLkh6OyVSEWzuvkZ7jzfl
5NtfTHv9t/FOeegc+iwgpF9O6z3Y5i11J3LqY+zB3h2mFqnwortq6/0Nk2T6QE3I
AMbVEqG+RXVSMWxKzsFLonvV4N0Wr3CYIP+VYu/sFNsBK5OPS5aOr6EjMOA9mpDM
sA1ltCDkFDHDy8vu6TLnREhpTJnIF4UJ3My66tghF6GryZ6KEN0qB3C7I5FmKHtE
5QYlQpoPuEGIu/FzAelGbWXIXCtXDPLDac6deE6HUiVpRBnU700EasByichfM8XP
egqmOnywrMP0WG6zrCCqpryPQ65LDYaE4o/7tXPoRI/f+01KWGh0/OM1VDZjaiv8
536CH7z7kDjBHQ9vRZhcmUpMPR5aVOmyu1NjIaGQa1y+V9BHOX7TsHA0+LR4vQo5
gNKFrP+s7jhmHv6BbGt5h5KmUc0l521CZ2EAhB0Fh586JfmGIzRIv631qWNZKz9o
N935KXdUD4fdV3fehuAZw27wOuEAXd0+X15cOeQZ4rYzJaFiAjOOVrfGIkoudc67
VMJ/tsDGwJsJmCSulkyAXvTnILctiwndbubmQ/TwUDCgZvbXk2lV8/+IV/sPTjJN
gMe81w+ZkznGKisnCyc1QlfklynD5sZxNLvAI/btHXgpfFEkB1Z0zOc1OqLASTJl
318jZMq/Dyb7tebivledKq00lncU6hoQ3PiYIrDf9LB+RG6LGdlKft5j+GriPaJ2
kXB3fbj16EzJ3uWn59K9p5ALnf3E7N8L7K4ggAQoa+yFdUcGyG0JL/3HZUFZZjGD
1RQAxZhaeXRDEpLu4PZ5+XMQdsKnOUKdBJu/w0RXgpfEmT67ZigTwAolvdrZbWjR
Hi1RhsWGMRE8Gm6HDAlG770N0Z2Tp3LQdOZIAt7F8pQR4F8NlqeY2uyNzdLLO3Pd
2Gg/jNjPNzq3VKjkhfUDX7jOig/jigvpsPi2UgPy6WxwWvXrclsKb7btZl+LIqYp
ZUuM9DRdZSWu5fA0jvhuPtcxSCyS8wNvElk9dyBFovh0A0gru9rqJvS7GKE/dEaX
Fxbji/JhtS64zHHq3C/bv3iRVPSwKQDVm4LtGXiV3IYvO4npNfSyfotBoXTuuu9o
9F38Y7MayYxeCMnEbPaPyQUFgVssKu8bnKrUiEBppptCzJkcWhqEauUDWG0+jVCo
zashRRVSxuIq8XBPFdpgRwPJu7pu2YX5LubHccqpoqFgCWHe2aenz0OAZgHpKRHE
t2VXZqg5wIjaGDkZ6JUATHEU3D9Oi2tV6X2s4vPKlgbi7UxaJx4rOQcWuOvMbCvk
SRSMTcUM83IyDkhT2pX7Q0Vf8TcNbFWn9VXSEOITn5CMStWHkhkaDG4Zege5yk9l
ZC6+B0h+Yq3rzIKIvRN0zjWlB2f6bKcO/khCWoV/dF9E8I2PheIsHQbhwsqUsPCO
3U/eyRmg2ZIcp7PEgAZlC/jDaGjqGn7e23WwjZzzXWBoubVsmCfZDOpwUeVbWQsx
Zrsj+x1HRF6wPV/U2wD1N3ByDAdidYWe6/jP+0jsNc5jowDjNM3gtZ3YHzLA1rjt
KbxKwptNot+VunoBhK6S96XdEjyDGtO9YGyKiG9feGd9nBv1QsUM/8NDIo8ifwOo
ZOiplYN7yvrxtVKcwD6vAnFI66uW8wyuQDBooeleM0/4emk3qUJmd5IoS9Nd9h0X
sVNBg6YjfdvHlXpBQ/oHNGGj+Xpaw2Uqk1QP+dTDH+vZ83QMV9ON/S/fHOQiPwRe
9VgxZ+mjU6/FQW/lDp4PqFFfb5+qj444HddKj5D9zCEkPMkkCYzFlCoZEK70jTYp
EhrLTjW2Vv9CCtdQLJ7EfgE5gv8nVj9o5wrzFoZAb006H6Na09l3lEaCjUUm6c8a
bd/UKnXqvFcIJalmqiHruDQ7QFCNSQU+o2ZZRqg3Es6wnUcYW/rD3aBO2ziwCqwb
tSme83Z893M+ZQu47OQuopZNGpyN298Sd4ze7VvDJ1NpgkSrE1xWA0u+dMNQ5QA1
/ZgIoMtc16cHq/7BvyM9MRkWC3Vo4LixJWwXnImp5p+p+uMUrrvSxaAq8bp8uSbo
6MHT3ExIBDQrwm2kSNF7tb6zae1MUjW7AJEMUQPWdcr788ZvRzd3Fag+f0hD0Ekt
lHBUKR6WXrd02w5paGCByA42YDicdTaeWd8mqTCtP2OPRCBWwEC4OvdVyPkudENy
fcDS/inqg5UjarCbNYD7RCcjw2OgWRQURx65eNAlHuqoYJ42ziTBHISoAYCsYTYA
HcQNvkDhV/qOL4qOKDLCD7vpopeehvWGvimVwyvtwgnAHf/duXq/aBURqB1KmpTJ
7w5CtQfuOdQcjgXIdv0k/DsUL2aVV0g9wbaWF3bZFZkc1d7HyeaW1CPjcX3EesfM
7HKk/qK0JnHGn99OwzMovz74sBJzBJMWUQqrDprtlLxDIaWa8BOM1Hxn7ov5XJ7i
krCQm/dKUajxq3TSDER4BEcLn04boCOhEEwJgy5dw7qn93WkeH4PNCcVUVgJqk8X
RitoIN2a9btgU1lt3GPGFxzr83uq+LaLWXF8qmJZa9HAsuZDVcWO+sHROCqSuthC
uZCBuu435BRJci4VRB740o/NSNT1VJkrADula0ccSjqJFUwSWxyyjMiG3Vc3wGAp
YmpmV2Mi+Rl+llKEx4A/9abcuXv3jaLbct1ly+XfOulT/NkKPcVhgwuxhVrMtPgW
vC4a58zRzwc+MLfmJz8sZAzEIZ8qARjRXS3pSazT7gb45wmINs+4Kz56cfgAhCv1
Y9VVjOok21DAGl+qNyiyBAyutRqV8eUu4JbJkftz84XthRKPwSaggJRDqPDWoFTu
0qIM0AK+8IHh2ZYek0oM5BT5wc/Z0RIdbaY55K/7JJRvzkY/T6twwBkf+3HNFA5/
WMsIkhaCb/tnN2cCeixFXzNVkn86Mx0w51IfUlyTck5545W/BALalLrM8pDhivvy
4Su1MeagLriuRaZL1P6kLMDGGsEuAwbNg1BdRuFLVYd/gaArzAzMoRhavD1iBqqS
iu2Wnk84oPww5DLxBjc28gxw0zr/Op81NP1fDNc7bllyytjFBS1PM4z3dfxUMNXT
fXyGBbpXgMpd/wJTMq3wg4sKD3OJWHV9kSBM5KctgyZtXM9sIFYpF7mlyUYBOZ/A
Ss9dyAsrXoqbsJFLwOsi3thxDEF8YbHUbeWov0IX4Lhb0/gItIINRsh8CppXIlIP
rFmEcwm93aNx1WlVwWB1qTI9a5e1EOWH0i32hshpmxRyxxsb3cBLEKm2SYTf3KLd
H0S89FaZjdYSq3h1/Rjt3kBspixnjfx8OzDL/RJlfHBlTiFyMfLBrkaCrwL7ubfb
qi1XYzODdQmoHVZaEBDzwXmJhX1Hbmwx3OPCqbCRUj/aM5goYCzVsjUbEle1l88R
5//Kw4KMjH14hly0pUNes20bWVMnVWJH88vSN+3Dt35PAtAw+OSEe+r0vlj9VJxt
Dax/ggK2D5k7gHueUFcX0enOjWFoggXKJ24NgJp00GI3oGFic2PspUwRW/PBAiVq
Z/EvTZssmKzRPqYPBQJjO76dsZyXyddaAZ/6/vmQUI1UdxhXB/yiFUaCz0uwQ6Kq
hpKR7PMg5tyBwyoqtpzQuh1WOtC/DKSC7wrH7BhdwXypyJbNRVUxiWJKkU9yuzfW
XNvIjdC/WcgJPm77ymZEC0FXNmgOvduAp8vfeNVegCuLw9i2fTzHfWTP9mF/Oy5G
x658D1Pj3uDOnd0v5TEHRnyKcN/E97CWEMiE7qOxE7T2RTBipC3D8nEz19emGbmR
nLOYmDmWuIv1DUXgvodHrUA+RyMl6jGWP42B0cjkNQRt8fJrguKG1BOi3B3S35Np
rMnH4KHrPDZxayofghwDm+y+RMNQ1ZLb2JNmiwp8Zrhtn4Qr0/zu4coKEj0UN1iC
3YVCGJ+29n6XoVUKKpA9lakNVccuukoWbHA+DEYZI4VBbO/zAJ/hKxzmXCoTcftt
DqC11JtWj7QSYxA1gmLx7hxSjGVHsvO6F+vbHrDZcdIHyhboikV3NvkjWM1KKR7K
6hKbNA9o30UdZIg7TmVsqdaY7Jfq1Vnu5WfUHw1W3Le3S0a6t+vDSGxSPhxEFmT5
QW3YhpINYkp2fUFKskSRrORezT+1F+1sOZuvnHplMOwAxw/cpAhwmdTjMN0gmPM8
YA5KFl3sU/6LzLOqLY3czXCVyqoroppPBBpiU/WeSCwTzsyAl+iHYyDiJ3J7l6OP
ZZFnNGIHws9zBFyyfgOSIbmWQZwHK02NsmwO1K+n8EFxXz2Mla1PTMqD8Ot5s9Ba
RtAh+p/Tx3BnJZy4lFBB1l7ehwcz1xO8A9H2umcZ/6EXnMOscXe9Ev4f+eP+3EyH
WNEMkpRoOI5i0/lNwuOAQ6lu5Jj4WrHLtboFq2VMCeMox5GjNOer6vPNFkJOFezr
xMAPZYTztrmzAnwTo4e/JNDWdJos1ued2i0s6CVPJN1sEUCvq+XLivia4arm6xlR
nGuTDGaANGGIhC2awltzWwUy8pJG/nxY/MauWDE1cEKvoWZay/sTI1Z3Pr8Gdbh0
M9feHWlNbIkTnvxKBwHrSTZaSi+zvzcGgCm5Ss84EfmgFiqdP6VujuaFnlNUu47w
0a+s4omTB9/6lmmH5VPkdDeuhFQL53pKAp29edY559dNiKVWltw1Zs5EqiJDKOUS
GG8corZMxRQaBCfqOpJz7Id0XgdO5q+Nbh4/6nabmRuNaOty1DaqA0RhdYS+Y6d6
GP9IbcMTdWDNWN/t3FHw/3bMC6kAT9+QCObb20nBya6JB1BISIrJO2yTuVgk+Gzq
YNHFrp1UXZS+ngZHKgYzM/hW8HP1wtKasswUI9I9nZkDCDu7y5pk7Ue2TOIrMmgM
OqDQA9jFamLEk6brUvCMZaMqv5LU4OpwNf/42Vhj+JPl+VSL0+cWay7Y9WXu7f4i
R8a+jE1VjKNXrBysPtZn6Ds3+2FtH2giX6LJX0aUSgmhcRI+KArWke0zr7zUCM11
0TnZnWeT8PpTPeJwaFrlcmecj4GBeFFq9Sx8Unu6VdG9CED4lS7/hilIrxJAI2ef
qykQbRDLsEmNynalSyoGv1orZJmzTRHuQHD/UGTsCel3ExC0eNeVQ7RqjEPY4OOB
vhQdf8qtO6E4szzDANlIRC/x+5h8EQ2Ikj+fEt7W2uT28E92UsHg8HVbDqWxgWVb
nndgDmvbRtmecUEKb4vyzjKLT3G9kolYidV3HJM4hpeQTQwu0DFLz9/kbMHqkr2J
V9ZnvfwjC+9VDPQ2T2RhbQUX8AjR9gTnBtetmfhYFl9nxYjaGBJHb8qKppUI+Yya
EtPdCCHcbDEknXbmvqfCgMRqdvtNrXmIaq7LLNFN44mcx/ByVjAQN9Z8JBa2F0TY
8NPfImD7eH7dy7nmTxWzmXzYp3MhITV1BhdzSU4lbc9PZY7g+4NqbEmLAQKISzdh
NSdppDGbB6wEhrRBv/2+yN21R7jn9YoU71DOip4fu7YVQ11AK6ZE43i08tzTIYTQ
dyPTt/CTVsuzhcDGMulZs2f1p2NXHiSGCVzJB8rMhAbocL/DAq+pDt8y01VPajJJ
Fhiq7RxnzIeC7c8uzdnZXjgL8+XNQaFGSEix5G2Om38uh7BAWsgScuMyFn8UuX1n
rnWy/CZZ43HuY/KFmTRb2y8EMR6UHbIAwpqbHwCHClnmDSncgoh7Yd+/HL0BAM7+
lzED5LDBO1H4+SF201QQ3OUyINZwTpwhvO4VSodnq+AjCA2lXAAwaRdQwhOSDPr2
qMPIXZO0Y8xluLHZwck9Ir0T3LKJB2OPDE58dTkdALnLfrJ29VMDCrnaBNfCdFNx
0Y5Xq7WlkDrCdR1h45eRYI4iELBbEhoC3jva3D5GVOka+8x1t2WaxUmTLbE6+7Bj
slIBALzLqO2kZ5XED3PVn3gKvOqj1LwMt6dQHNAKB8al/oVRyD04Heem6an7tFZ2
rsDNQjVxTGLFzAIQvBuIrleaFk8mplKJKGRrc3ypGSM8SoXrDntHwLoCgsDH8cb4
w+Sy4mGSgPsiRP02VkWvb8zS5mT7L5gQlU6vHvZ6V5qSPswOphOsOvquNldJqYtZ
fzbZkieWg6eDx4U/N3gCoCj5OH+64Eky/MqDsg5emq0mLEdOQFsh2u+kaPYWPQ/G
DQIEl5+76W1qe7nYipt+Ft5B9fb9t2Xk/aFvTubr5G57dwDJQ/tbn4m+eC6m7yjW
r598Cdg58SKSzUvEEVVveIUuHuM1x2UTjwNF12mTF5THuUWoKayeY+tWSbMVVYo0
I3R7Yzs58s9t4MgDeN763+/BYIx+mG8HouUL961H/fFKicydcwH726f2W25OJ6v6
cCUzhgD4rYSNPRZhdqaKebEasbFFlM6FHNkIUBHxGRcrfMzoNDDbT8HaptybUhWa
HaUUmtuFB+bzrN+sp4tGHHJGW/Os/f/65BPAcTUiLcf0A+yN9xDSOb4v9QydyQY8
NWgyDRtV/ik5UALvX2wlas5D87a6Sbzr8IyGatX+qnUICvTfazfEojxw8pLH3Rtq
FmkCEisLxwB+ijUhqzfB9S5X9Xd5ybd5ypcwE9zBMPVBwafGnAz+LFZAGedU+SDN
btyZGsl43fennR8Ih87qyqzGmgFBnMrbGlJIfYTtPNv0wKGVxGIC8Z9lrd0pmzJJ
LzTwPHPZY8LfswBB4q8BpWHfqD2fYjyR05+Mh8AGvyrWlwvyGoTk0W8EmJ5XmtOn
3cMkJkLIj3Tirh9ppTRqKRu9oM6Fc1q20Iiwvb8YT9xbeDHKJPTF+T2RpROkrQNZ
7h7l8KER94nprjI/AvfNS13EjSn2titWBhn4mi06G5AvUZteOmYxkBbs5+vgAhIR
6FTJMWN40PCaiKlzkFipyFGWWkWt+CF6A1bWFk72w2OVB2WkmV9XkyULC6s5ZzE2
7ACxzXtamOZY239ejTGXDgbqNMldghYiRqQqXkQlJoRUPqk3bcBG0EOB4XS9sZeE
MjaIuLFrXfY3BHAHw4vKNNWguS4SCTUedcMNVWAAzsDzOXd7Y6PvzHH4Jdl/fKSX
DaDU11wJTHqin9t4ooTXV9pPlbeYtUly58rsXJHDJqS8SzUpxzwwu+d2Dc6C5asJ
+rvqSPU6WDz2PAzqh4pWLKhPmYw7Ie+JRSHNmlrmcFZi+lA1pLPHYiOKCx70Or9B
XA9ABAQtyoiML9WwOFNdii5pceiyzvE0lFqfbKDa5G3cjHUKvV1jQENqg35C0TyS
xxI752EhdrlvgdEOZo5QxSJe/XdqYcrllRGZd7fDvScGkLhW7Gze4EHxZrrxuczV
NCa2YO5FxhhKyCYwyDlDYf+DGOJbtfQFgg7iQcIVed0gUIv/z2qL+inATbKbYKu9
muTzAXlnqkYFRGXJow6IciNN0/qKctzGyvODB18I2TVmTLwTxX9r3vys8xIDDtuz
dysnMVntZRwYDdx8LwuMoSagaoOPjB1IdhOXRv45MlAgshMuNn7DIBp++eXUW2rP
fTam/wJrZ9hbr2Rf5lo3oaszNsjZgWV9D+Sl7dwpga3Xr0Cg9v27mOQJAdWM6k6A
/Pieljwta4q9gQlNPxr0YhagswnB+10TDv+v+zgt41VHWRIcpH+thJXDp4haD5/j
GT3HUFVgLvy/meA3lsbX0BcisV03yIZWB9tM5nMgdKGvdJZkrHJJlHdcPgD+A4st
T9E6pIAykhL0YCCbXbWPmLjiyVsjPMPNAtTaxPDLKhioCLEVuVcz0cLDHM9xMXk+
mjowe/47vzZyLZBR6FU/zJaFtQxW59dqYhGqWgLRRK9XFvUZE6eGYkb2OVRw0idL
FOVL6WoTbHhdMEbKDN8IN5PN+Fva4Mtb1sPsR19sZcMIC3W6reMTWweylRdgxlb/
IPYihujNq4BBEf+pZJsKTsNlGWf28c5r3F396xDOPeFnhRcLcxaKsLUrfH/DRZ5c
QGsZtZSch/pz2szcFhw7cvisGfKFXJw5KniMBd2+P/OuJLgkFqtBfiQy5PEyhtQV
+62jFzV8BQxsWAgP6m4Rk0DtWj2MaF+lPVx4VUQS5Pyy8rx0PZfw0FN5d3qB9uUg
n+H9svJE0aMxcGwDCcAfEIFQK/rAoWt4o/znsevY9WvpeRVrj4dqJFXyOtZguv/t
wLOjXvg9BIh1/Y32rO7rTZ2w4vjEIy2rmvnPCR7UNfoofEB5Nfmx50FLzJWuG6xM
yX8PiKTidJrh3oQuz+UWgWdCnc/pGwVa04l2hgLdzVJRzdadDe57FBHcwR8lf+5H
vv5H0zVnIIhH5Vesxogz/p27zBrkCcGBt8FXlvpzrb3W9/FfAWIAWyGxSAkpvRDr
G+/G+ecvlR5SSlRHO7vaWbIyD9HMGcm4OxFNBDCMdBKQw/rWU6cskoVhAKldvDjy
QG0arsREEL0AB4AEOAAi0TFJRqHfVJqICq23VjnC96g2AoPjoABYKVg5QwsuIe1L
YBAAg+nnURN/0YW5p5jK1OvNTKvegaxSkOi+9Vt/4wkdfpkUuayFA/W61CM4zPpZ
Wu0ldpg65N/VSiPGW4y9/WjFFHmBWnc7lPXa7Vr23xaVNazy2I5gjYVJNbF0LikF
X1aKGe9+Jd5UJZgrchBRJU64NvUHAvsyQa2CMDwdB1E16U1ri6eHMaVZzBXaYEUR
qkMyN4pO0LjAODFvUTuLoC4hHFPeYi+kpXJHpujPP1TlwjAP1YvwHfpqlyHP5ieX
1seUKAatW0qLfjFvCsoUUSHGWNz0eQIjMG0UdJ7EfBb5Hu4BDcsHHeqUoEX61k6X
082+1OVT8W6QP+zbybinnDGHD2XCAqdhOn/U7VVcFKzDPBMwmMC/I7rnuIcCm579
rRUVLC3pLscNr6hriVkbdi1wl/NLqQBoKj7WzcYfXConcDu+OTG/hVhebDT4R/ZP
9OTvmY9K6fSw9C4Qb1o78ZzBdjLf6RZ15iwrQlVYlW3z+KQh1suhZ8bisycVK9Cf
OBogVx29Bz/wo2uyib1O5ZVHVlvW6AvPyiggcNWxYEwu4qakroN9yRqEIcxcRvff
ui7njyjK+bjAA+lxoOLkpYunMlPKn8w9P2u/BwCPRfPp41wjKRHy/VyhHUJgOWBj
EN2IZTvhzCbH1OqENWqDNhWeB9IFoO9EpsBd5LXKF2IqrcbDhNuOLcpGI3OO6Qx2
mWm+siU3FRqT17JGT7dPUPBhNpTuTyBWVhCNhubRywTVqZrXRByOFY3GlkZTEp4w
ZXJ6BDmmw9LNY8e7Q5NFzR7bVe0tAjoqPPAEQ4PkYFZoCYc2t7qawyM5XuVKwUby
Kyxl7tavcQENApjql+tvJ5llFG5xVBMjPAh06uYlDpaz1pixl6pFoPUHhlBYO4K5
nXvSFJ/v//icxqcl+I/In/LZJRCl+jewnyeVgNnmh1295qj0N/ARkpIeDOpbiXz8
X+n9nr+hZO+qVtIdI67j/8DcsPLpX39NDpdT7ekhfLwc3sood0YjewsjiLdz+gaI
OlgQ6qsGiP43GsElTv4V0cx2sk5+qs7XzB7gJbfITjE65KWw7fI8R7BOzVo8BWGk
wjxjnnjgPpzZdasOd27rEOWHtsOvyPw3HubFdghCuOZAyoHmu6mCnGgiPh3bIfz7
Ho1hqBfdytH19T2Gm1LGSNYzyubPo7tiMLkSerd8jiSdYkdNV2tPkwVW6K/RY4vI
nU1fX27iP9etDD36LNxBlrYUCEDEd/SHgCMjJP9l0jLkYquXxYE+yIiV0qa/EjSo
XBvwPS0jm6k0blZkiM3o2YmBnJT7Q74UiFbjD71xI1y5QzaREWPmnl5MBvMGxJRf
PyR+smvnM2ExhXDDhKGYACcnsFUNPU+/vmIwQKD3Ddf9MJ2/GRZr+na+myrWZZGY
uODdmLsIIjJFBF5TOegaYJHamvHhdgbdvH05/ltxSCPOFL741MGq4t0Qc154owA4
qZwnjwqA5Y8pqCwlG1FNap1boKFXgpQZOyG6mORucH09f3LTm5KlegmE+jxGdtxt
KQJY7Bol8EB2+lZgpH+0C0QdZ3xIYVjlB0eMwtjojUoXyQSCalX7a/mqfGXNujB9
s4bvnjYWKhvC20RPVldHECy6uUwSkM4Hys+rl2BAeTMWCP8W0o5/uwni27f413lo
obeZk5FHIQJ2fdQUmNQMgBfUPrs7IcYdUtMoNunc8xu1prYUHCHs4dabF0enWbfs
Bdg4BhqvnW4+xI1W6v2ggzau0qkw+x9i/g9v8hGAYQaHK8kY096F1Silj3DqD/dm
+GPeV0tcr13p0fc5jr0hJmss4pYwv+r57Eaeia8gwITj3gKIiWJL4YB4HMoCI/mb
Ma3Ukv0n0E9O01h6Yrj/Rh0KE5M3nRl9cG4sRY82ElmWA8TN3kJ6PnQdHojkUr4Q
JFop7hD+hPNXmcCTm+sogwA1FjnTvkFw6UC2pdigMeTdzxLFe4FJjxSUHSQxGznO
7dAvujn1iTwYURg0ldlorHqeGF5hr7z1qeFU2Pziwnh3brqf9Cwgv9iXbyAYe/sF
q4CaRhQ5JgQgaw8FTNVhYhKBFjNOXXvnHc/p1vGxVHTZ++zfcXJbY9obWX0+xUb7
pWMm2oihxLxeNK8Ee0DHnr66pUESuHxAA20c+OXwK+dGd/B+3oO0S7ztV7Pgjchk
cd4iWN9vlLtCLGuWRdhMuYIcfMSZPSUEc9mUkIsdNxR3qHMh+sW2aDQjIJhdYUiq
AN+cqv6qoQMbW8Xh7kBs0hGIY1jSEGIpnqHHjftVXhcmVo+OpA0DiwXNnV0X9SGd
1OIFzh08uj+BqMUxzNf3SqImgxzOXS6OPwJv1xCucnalXWCkp7QsFvOTanasovYM
X1C92dJ5GpKUxj9NzaWuAyKCq3qC1lbqVLTM/wkB8NBSoTMMHzpR7PAh6hAtEDda
llbjnjUiErtVvixPmse2KLpG6kZi4ANoxBAGju34c/zN568XCiJYIb4w3I7mLJMp
YcXQ9DSEeXTPmriaX/U5sFHEhiSYcgZ/Se2BdK42K7HCMz7xqgAPDyDx5EI0qqHq
Wc5CpaMtVIsw/nitKsow5X+s1CQxSMEGkrq6RkPp3UYar/8GqR0LVSxHjf/hwDpz
IFWfSnQ9eEtyC++YIFmfA32dv9JfaJhRgh/DUh1mk1IABNsD6sVH6ze24Q+71911
5tyA01Th3Tv8Z3tkwsuNJ0FPqm/4MKrNq6D3ln6P2aAX60oZO6RHs0vXBcSE6r7R
4c6MyV5UqrpoNakMZxN2Xlupe4Jx88SwfhjWZowHpOtFVDNQ0hvRBDC7dzIbdhbk
RmdKXOh50gtuWZiH+G21GlLy5mlg5deT3RWY9B6/paVJc7A1PyS82BfSulntAYnt
U+jtslGpVzBCqwW0yrvC9S4sSXFJAPJ3GrtwQWAxLQaZAcG80Y1bx+llXG92d806
I6D3AWZKlkZFd9uZXf5PU9VhZBcZfsslDNdihIUevItnqNXTnU9rsQNXzB+vFjwz
SuN9cZCILLzN9CA1IDl/KqNv6DE7EzFSp2rHGvVXpEjiGatDGQSC84wxOboQkHQ6
bqsAM2hGWQwGhJ+lLD+b5LMLmgfPDDVXfBqbTkvh9gO92Tsk5L99VPGklA+y0LoI
OaUyXNldcjGjZIhskaku7FO7U6fhk4YXESIJwr33vW2Kt+ybyd3Wjj8a6csH7KYW
mh/rOam/jL1nbDIOyQ69I1NnEGt5L2IKVE4RG8TI4EZ1qgjA7EQ6RA/C95VNld2/
B/9S4SV6Yqe6EHFFd8oVFRkoFYlTBmdPlh4lUEY4YVcgJNrDXSkYOezIto3pyg8G
CJPeypEuZIFlQdX1zZ9lbHrQ5mYT6TvODWpvOqbc+YWFxOXR0p/qaMaY/mgqMFQB
k6NcdF3rKFa4IOUe7nx3Ydh8ZkpkSi8kg4W3IDJcKER0Nc3oCyothiW/JHMN7WjY
x+nd75UWODCON7sTiCW79rGUYBV4fkhJIVTmNhLGjyxBWX0FyMJX8cawNMnCiR+L
Lkmxqi70IyrGgzFHVwGEqKT7rVnI3uylHFbz02nyS51BeVthvu6ZbXX7PPN9yQAy
gSNiHbNtBxZse+146/S53ObvjYdnailu/r9zMQ6JsVcAFC1XTg5Nh4TXISkm13ik
JFi9rUnuO7kTAfBKqnZOgNfS0q4pGD93FxisktPgZwEUr+fAswVQhyq72CkWFohv
LwkqI+m+Tp+nBSwdCidt1EeS4yzJGhSCp+2hj/fEl2c7BDx3hR0bNDWuXrkH92yu
CjvODIlaYtQQYv9LPEiMMKvNQJrC0E18TKuOevdtTS6LzQKja3lTkD/cK5xTSgiN
yySKeY0LVaclcO9QFDO5A8dtffIN88se2Qg9BJ16hHjlskUz7zzlr9RHYHFA1QeW
AHf8Jg/Cxi8IRjNDPUluO2gcknrqXbrUmNJ345kcCvIHIG2vErZkqQDlEuGRevnP
HpJyTH6Na3EiAhqgsyMf8g2yYHXzHn6j96O/6VODRrXsMQWL3VjT8bTFGnCv6mCn
AMGL0db3Yi6ePPgcJyuSaXBrP86rTXR9kFOdKnCS9eLK+Kr7EO/5YPP+rWuo+Jec
38FEckI8XxANZ9RxZph//tz1raeU9YTwe/7wmfX//lvW4Ey5XdBdrBtec1pyKC1j
E9vzMevAtVg7IaZhERv1S1TeCaQimxMRmmAZAKSUp1UqyOkS/9XbnJbq5Car1nmV
+v3PARxDppUtktCWqnjRxdn2+vmiIhRH6LbW5ZNCf20X376SZqN5JnFKB6cG8c/C
R7J9cuoUZQNVGi5EegbtVGwwClMUNDwDMq7LHxEqnD2GiNjP+uTrxUpLA0PyZJMA
pl5Vu5C1kD2+EmHP/bqNP+RfAtHcXvMofOY1P78rrjyAVv5Sr3UAipoaIVzJ51aC
D7bRtzT8AkZ+9/SHpDzVcVoBrst8+LyjLCYwworAXzaN7hxaf/6dgfe06bu6wAtm
MWoVw0rADpRyIiRwE0rNRbZ8aaX2I8O25iaDyjSTZEZ8oKBX1/50703YV1JZr7NV
c4LEXqrtwwo8X1zN0Zkv+L08/65xHWg5QW5cvg7MFyJTtAxVEI8n1hInOFWVN4D6
h7Y6bZ9Cw0i0fFNPWcfrZgjC9We9/c84bjvWqy4wK0sCyHhWB87p+UYSOnPv0HQK
YnCvur5BNfQVK7re+93PxrLhU35qZhCHlEwQ7cDLEw8AQWRKbk+cezRKC8b5m3pp
g43+sacDwh66W2QZvKgwLfn30X9HXYd07Ki8lzbcBQbbKdBq591tLvZCFcMluFi9
3YXWDdvXb5JVFUKsApBNHLErtMZ/sahV4DCKzXwAqqusVDiTX7RRcg185GT4M1dk
frCMonYqDk9cOo4argd9W7vC71PpHWvw/8Sg0wnX93doCqKiQNld7x3THitBnE08
ejMES3RTTi9aaVuWWJkS+KJIKFhaikHe4Kq+lzZzrs/Qp/SVWBa8U7R4eyzTk3Zk
Xwk/KYW+tfP+g7ME6caukKga45QYXoqmqryyUDYRly1CNMpuzQ3Z/8dxGyMrTC/8
GkTs7Ev3PPhgIJh1Vp6f3fqm3gK/Y4Sa2PcSuolS2N7qzHPB/R5pcm4eM9GLRTFt
PPJmTWUYLCOzKpf1E1ljTHKRMUECzOFGvGv8LTWVlJeYPy1muG7Xwj0BvifKIE3v
pNN3Zc2GoppMSYyMmJws+TdrhaM14/N6OlOcOw7yReYOrzZe+yu/O0nZ41Zgynfn
TNCFekGc4lbTc4gLY8FY6Ty2Gtn7vPV38OyDzl+/X/qQjN3tuau6f7bcMxy1bJuK
JINoC3TuIkDPspUdOOr+Xt2JvBy8haqcRj9Dkcau7PNis7b5M5ENqPVg7tXtapX6
oJOPO/uLrJ51niQGAqUresWjnL8aCeYqYAy+yDdbh2VgBm2GUEGr9zhCF3YYoWOo
rBM4GwRNMcskgvlPoWKvLqjAMDhGoh/gn7+FlZFThU2VMuXGVPjUVJz/QlDqE7Xi
7jW+asYQDh9QcCM3mMUTWreMrtiTc6V7G04S3A9EiHWkdadiDbYt2XyjtvepdcIh
Ql7d8uZMpHT1GCR0+mUS158KYWgac4TXeiGBB4VfS6YoQH9VM34huzvQz/6crwNL
ST+Xf6rwVKvwJ882S1ErLQbaqfsHfiILCb4n/sBHpqrH/9oFN4pIB7tfnYH3msdl
Z28fEdcrplMJ+Si+x9C+5sSBqMAslSvRUA7FjP1S0NozDfxZZwDEimItx1vRvXa+
ycQdpG6LLF0bjPXAvwbRCLSAGJ3kkxFVWtzsMsyvVnn7e+MZiTmhZVMtx0ltqNTt
z2dNBFdDACuXHgOppfHUhozi70kNei7Y6c9DSxI+sNC8Y2aBpM2yJ5sekuXutmG+
5tHjIuvGEBhZVqaBUSvwXCUZU/UrNYCou/V+InE8iXWJU+PnMijmtTC/DRV6cYtz
Iy7lAbMAyJzTYZAyWDfiCLsUSwY+lSxgVNHt+zRHHzqQCBQypPi3wozM9JzBeaii
GlFPD5UK+JP/j53Pqm1RkBaMWGDcQTTysB8NGG9H8WmHEkwH7Ar9x09/AeLn3xlL
35h/R85PWe+Jo2yvxss++30gXOc1ThYXuhTXtNO1t+dcjO5pIId82eOXLN2HYPy0
LKLATNKKc0QvdIg2jbSaaQuVGMEBFu8tAvWgftD37YYeF9OaAs24vt5Qosp7nUqo
rjCBv71ofiFguFuxRxb3Lp8j6BrVqBlIrWLn0BfslLhnen9sSM/Z+QeibIstYmW1
K2f5eediT3tkG3uiKXbSCO9zYwoF72sPpntMiRBjUSIt3Yr0KJl3WRUxEnbbIGe/
TcZELXBUuT2X1F/Do4OFYcFcrv27q2oILrh4HZhjwSjLlrma7Wwn5BhKKhFTXfTP
XyKdnC2vianjvf8FW98/DkIW7Zqp/XM7lFylXqmbjfpor1BeV4BKOSvEbZr5dxR3
dVjAxNLIaKqxGJW/6KA8Z3fWbaA3WztEexGAslac70C+pf3h3R2kcLgmcvR+azi7
8N86hOQHRfVbN23ALU1oIaZeB33GYx4Z1ZIRDGPgzcvZ5p85durOTQbeebSLXKOB
AvDz6iK0Hyb9YW0nkK+3vSx+ho7T+A6n1r2DcEchUTyja0krt9MbXuGzgNOg3wQl
0SA0x37aTuRXfn3Cr3KZad3LgYPlrb4WOW6jDkmhDsCeeLzFPMnvaaJlmbmbYuyO
HQUOO7Afq7POd2CcQ1cWeR44iMw/ykynD1hhdmDszJR9+NFXj20C6dU/RRiUrRt2
6k7+aePRWGHBge9x+Wbs2gy4QztQzzm9FRx+IOKgZDAe4ki+eIxA8fAyTa5VhLAk
JA4Xcpa11YdGJf/wL/QUXgNm4EnAxdtzNJC1MN33kZuuwEIKGc/KvmVRuCGYSDNF
z71+q709TLO/iaEBaSiYNqIak08PqziIe8tQRXuOVRNLYVLEjEcvRFcEsYE4vDpj
VrbnOLxKOvVtM58dxFw2dPoVQsPb4AUbd81ZGqqYoAjXIEoaL/wSKMHIPQ/g7VHS
9LW1Ye8V+GwmqQbKqW+QKiUZTUAlz+oXMuO52/1Yc7EPzeIPfTL0fP0hrNnnFdoT
XY0naiyqTt0/10vQ9usAHmUfzQLgJSY66VZJMZyH7F9C7j6hpNkpemsq0cFz6z0Y
1pHS2uqxtcwJt7BBLWd2YO/VTDxSIXb18L2/kYFmH+CL4AYU87ZAbDllnYwGQBMR
xAdgm96EjS68Pu6WHS0tOPJ7yQX4pyyInHHtXD6EpaS2sj8SEJWBVSMPlSmt9I19
iHWv9tNjRlK/+doK0zFGGq42nRLJDoWxfDJK4NyPapcUOeqYjNuP/mQ5OsdQpKiz
v0KgKrfLvt9+rzMnSS0n6gu+0GcCczUlHjbFQhyish+y296TdhpvdM4Oj8B2saTp
CFO9W+XsuOkxgTZ7wy49bQuenkqmKmE08+5BqrPm1lIZhsuBRBHezj3vzX4FnZKN
ToJ257KSuXnzrifnFO9v5KhRDERWGzkDniIbjxkCmHKEl0P+N+LQup7GxdVo/j5U
AgSt8cXci5VlYa4odX/xa9LJ3ug8VZB3yxbgvuFvt3L4TWTsHsxWyN1G/r74rL+k
OOwK4xfayVHmYI4Ldf/KnjO4BWsqPuHBaYOtYiS0n7cudAbxSRsEYE0ashNPYZyq
L68UfMQZ3tPnl+yp1iwMM7x3Upxhbfl/5X14+IEryXpQSWMMhIfUuuW+6Ndz8lwT
+XJni3DeY4MR9cEEg2X1r9w/JeYV5jKfELPoLuQ56J5ajDBgcSFHOSMRJzllbdh/
n9/gXs0loji5kdFebA67ztk4qsi40nrslGMUoqxGfVdM7LiKvdxZgLzMMz9Ic0L9
kW97MQHkR2mrkNXvjWcS4Na20NT2v0qHRGKlLSUPKkMRr9VOp9G8SZ4ekfNQoKhb
puPPOXWk2elvjTaX9C3tIqY9N7r4mweNXj/Ys8VuvQkYI0qHb8dP8xYiyWJptMTD
n3lmiWFY0rY3UprRV5xrHpzMizvA9IyiGavUaKcjQF4UWPxLzzF+kwxwwC3ZWlIO
mGdWpPMRMg1At3eEzJMqX0z1JrQG2ZNfCizHJEkTXA0YdWGmoRfV495NJUWIfNmi
bcnRmLDspZ3/JCF44IcNHmNxPOGxKR6lPibZgSiN6SGFSay/2kBVwlqjtFyYyRSO
pC1HoLPfhX14SEJz0CKw6nMO9pwwycM8aRSTyWf7CgkNSZu7VweIITgBm0g9urhF
FjIKrDlp7YAgKG7zbd4CtOsvoB8tODFB2c9ZTDGDqGVggqu9JuyL2BG5hkiQ9Aq4
WgrELuUwKAzep8Oj2om4ddxsChajdZjfkchGt6+hcKZRYWH+2NXOP9y7cBg7VN1/
KzXRwXTsAbER5zs7shDbOhSmo5tG3wbrwRlLp4JQBS3TFrZ0vyWjMHmqEKZ83OZA
d8tQtsNsMkkNpuqUw/FkAeChBDmntazNJ72zWgTXqWRAVfdPcrpWVkcDllcrK7Tg
OQdxGhenSOWCDyfN+iqNUxo6uiKorrkh0aES3poY9XoN69RFrQZoHr5Dje8YJ4Eo
EVM/a9BY9nGBUoHq7EX8C6D0+YJklA3P8YLxBYqigTv8KY7hSNQeCIJtomZ1msG4
u4vm9FtvPUFTwK+PlR+K+wz05qyLcVrLY/UZSRKMh/rkFiKZgUtUiEReZRrVFmw7
T7H9QrwwXgy1KolEH1+PdmS0Xx1SohUkcgAfPK9yYEPGTJw4ve6rXWR6J6iaEgBI
u5R2Y44x1BdswBDJ6ESCyV1LLO04GcGhUnB6t+KGzNTSXKWOXIBtvRAZwsMXo96K
D+JifwqdWoKHrIGUbqJxgh2DpJ3cGrbbqz+QFcwPjdCiLCD8kNnZcBPSMlLEEhwR
eGUaWu6gp7iVsuPIGgvPnnCPiAmDMfOr6qku9fB+6ju0laHZSeD/7QJuAzyDPl3C
y+6O3zcSbeq4ff4S6yuhn1mOIErx+sYo4rRfH6uAJ6KVjEsY5IV3o4/PDatSaVJY
pIGgbK/oHBgtd7P4gtvtLum9x+LP2lOlyd77Sd/K779CNvFItpETbUySDIZF+2tR
BreKLDd75ySBJz6+WZN0hzs86zwhBfNsIAZWA79klcV56zCInEulsegiKj4wp0DR
5lTCrJwt5HOJ8DSjRaSArBOKxUsCUD9zEUX2xgQcw7R5QACQ0cZrTEgC7lGP7DjL
hboB70wX2ftsEE0SDjfWQSh1/32lCDyy6PeMI0CZvzA3x+sv3xj66IVBfJ1Ght1/
m2pGNdM3TVLq4aO6Lm9GdpEoE479PDpIWIDnhKHL70ceJT0A+RcxBrtOiggHfMao
kjqCe2iwfhmOFm7EV/rIHtYjFqk/mGQsXG+8ZepqFV5s0x/VH7fadvC/4EQDjzGR
AkiL2GyRBABur2SXf5bvjlDXBhJwweeJ7bwMf5Z6T8tTYX3DrwGAL3WlUHQ7VLgU
pKyffjgt60dKxXqzrmoXtVE4whhXzuCvHeUYj3eWh6dPx6UZEsGgTujlv2gARvBn
kEy9yUH3ZXagDKZov9zCCUsb0Fzg09S7XFBB73O7ai2GudhSJGEHlyXq48ydLFMQ
qIhzl+sicwRBtEpqIrbBAUjwxr8Z2njPDB/WDhyxnhU/WeLAuWQ19unqPqYr22CI
RX0G5fwRuNaI269l27e3OiGh5otBywIGTe0Fy7tuFpZupLgn/8bMow/tgzMHD+fx
FDs0gzMAtqYRkzemBWPXsYnNobB3cGbObjNe7SlOYuR2iiSbRmhAM6V37PahGCXN
ixqecjE7VkUMHBYn4zZ3fsRuAXH/grvy46ApB6QIVE76WNJacj4uHNB9/WDqaL/M
oyYHGi5j1sgcPTpIV7UbjtlHUPi7Ahq9LMpq7mAK8NnAUZz9IfPd5SfsNd66ALdm
d4QJDI7BSTYRTnZgOIPaCw6J8Ru6t1Lw8qtsPYAY3nWg6CFwuhZ6cpkJZeyFDokD
2mF1JtjJsZ+e9wOFk0jC+aAFzDPXjvL3bJOgupqG3LAmimkcJJOGi8KConIesyhx
M1HL/899+X1QDXb98rD0QveCot0dw2pVWI45H2PEcw3wb/E0RuC70MX+k+Unmy2E
a0E0cWX1HGIeDSqLAfWMaGx1AvnprLEFNIV8g6x93WdFeS7O9rVXgfNoIr9EUkI7
n8QQv7ycYhrX9xpeBt2qCY21oaFsbZQGrbQuqhMEhSAibxhpz6mpnXEWp7M61nMY
H0CO+i44ZzvT0di3h+35V7WZLlDrOMp+ymIUKxvfFafgh7lgiXmAb5J0e3T6nGqF
4DKfjzjjRqRcmUi0lnP6JpV9hwnkVlmMiStRjq6ar+l14mLkbA70UAdJLBEZ/ZyA
AmA30WvQKpGEgfnAawudzq3/GNdTkP5rdZ9/eQPFy3W0Y3hBID/GRbz0CHbtuN8E
YIQwNUkC3QGbUwhYUmNVhOQHCDmRCMYveNRJaUf5ngEQXXMjUFS1S3Z1df+Gi6ov
rQiwyU5bcGElwzlfWhT0tT3Urtn0yIzfnctG+rjaOdL1TbO57ZqQ8potf3lFbwCp
OGkyX+MzxTduEAV3zZ8zs6GjHQPWmgFfbIX6+EmOTnPawVET0mY2vAXAiePmP3zO
d5nxAIkxMTS/cGjGnL5qSU+Eyk4BwfR4HMQ8r1PIXty1KCYazRTfyq3ZpmWtu4h4
4HziCSLs7QdiCrSROr3tBp1KUI+yoxf5gw/ibHjmmtdI9gYMpyLWyj5TOpeZ1Dr/
eDmzKBlix1Gjnwf9IZaTYesoueR3zuiF4l+KCBdMu1SaVlOiknqvRSYYhMWDJMWC
+NI8zSLjRPAjfFEMONy1YkLYobP5N3wKVa+UlCbhui4//5b+pBpqVGs9qeFsVbOd
jxpHDSA4nns1rf0kOcUx5tELdrTVGBup5aSMzcA6/s940vGO9axYn0gOAGDZlOsJ
7frWFKqulEFSMvAhXWR9ipPu/YpoAptHF6kdQ+AJq9jBX0QWfx0XyUALOFcVCYLk
LIVhwISvt5pMi2rj45iY8xCRLiCdls4P1UGCQk/2u+i42vPD6+YU5XSb/McgVtqO
TC13VsW8miaUZFbO0cgRpOoiZI1Gai1l7EDlNP99SroQ4sOoX4X4JMbnZGhiS8M8
PMHD2MSJzxuX/GHRjybMx8ELk3zicF6NZaC8KI1iYpGLBGYwJmUOsmJbmQ7M+HsY
MQ7iNwNV6Fjo5YuvEozm0Px0SHLVIBbzaZwSCoacdoyEXJmXQesIYXExcLS4StJr
v5LFfWnIUMYJDz+x/aXnL/ASsneXBEqrJiLe9r/LX3L/XdzirYOVJMHFLbfklUAr
4Z87GR6DTEu9fhiyBI3D2FeLPJsbvRpOltKTTRSAWLzVdXbbHUAxc9NeRKF/kYLo
lvQ2TadDivS1Ph8HY9vKWdjvIjbd6SntQ3AXPtfnFCn+Qhw+Kvt2+l3NGFxoH0fA
a62LCLCx7ZKOqTYOT913uSH16XzJSVppzw8HgUVyY5m7g4e5NOuMhBIjSB7AniKx
CT2ndhNkZf756PcwqxgCfsEV2ERy5XQMwjdVb86xBS1t8mHL7hveR/XZkKr2xe5E
Ujuiiq3Pkj+liSv5ABebk9aSIosHNfUtlRJRu5pjZJ4vbTdHy3xuvC/JbI55Wxdc
K5Q7eEA2j6MJcf2jhW/7EbGNUVYN+NCGKdAEPRIWQw+BNCJT6Xhrt5ez3CPxdcNi
tseFkKaCEDGC62D7W7Di+9VYe5dW8Y0+/Wtue00yXVHW1xLiherdxTUmG+bwWcKL
1+svEjB0kM2T0t3i7kkuINXt6YKi8+hZzl2/NHSNa3kpOaJIgxfPgCsp6MaDaJB8
Miwn9rFNl5n5ZrHtDFsh1IqPCHiCZzYuTscdKB9G+GMtLYqR1AO+Ai4z/fizlBFE
qoa5gbeVDiQPwiHGuJAhDEkDFoV66fmGUvO3LGJKFeyrNRAlGEfuvKk3Vacs9cqT
jWnUSa8z1VVSbVzfCepCZqORgPRcLBia48GmMfP9MHF1HBmDGFD+g092BrUTr5eP
ZmuVekixTt2Y5L9oS9NvPddpfDtDlbOU/BA+ufumco+KDrzjRWUEIPhzvt0S0B3m
ha5Cb+lgd4FRZaxZ4LRQ6LtETud9gdK5V4LYlGsO9Va0hMMHl6hZ6NeIr4cPo+U0
1wnUf7xu0reZr6Gik035BhCP7wIsY5z/b3e8g0K2TEOdQwD0fAtA0t3MRlCCxgkh
cM6PqfExITQAKlJVDt98DDsbnGtjl9X9Cn38IbCbAt2IgtVksEkxRa/s6p7NrhaE
TOwIZDqPJJvWHIph58ZZ0C5KzmN7Xbuieqh02Y3P/bbNcshQbbwdWeTqk58LhZda
Oq7c4+MUb6L6XgdvDfLBHqnsxYuidYKU6xI001/LMap0g2+N028xPggH/J3byxBa
jZLBM5XcePHceV9slZe6xmLoko4HDRMCvn+urbvpS5bc7NoX0s84iz5vnIKfWlWr
heC+DUG9YoLOSF27Yb30ku9nkPQ3/eNLD51P/1ePXWEjBu01b8NsXVLcijUbGlQV
j9zAE1uDdg29nH73yg3j/qQniDBPGVxGsPqAkTMiLedqd4tYUqyVljzk2kCam+F4
xfGdaNKJpf6n5sD0GSwNBhCQJ1QjCcUHj7mmaesRx5fiFxnp2QlgWVbEVsoTJknC
jBbixKEeM2G36Npj0CrWLEl0a2y977XRSsHyK/jSEX2sf5vo0gr6RHQx5IFEOlM/
ZUEZrY4nq+M2OR+ZLOR3t6vJ+N/ofgeuTzLJfvplIjR0lckTQNL6zuALIOVxaqlo
Rgdtfhd56h9D0DdAu1yrGl8gg2PXH5mF/qO+FD0UmrZzqQ2sQg7qhylcFDoWnzNI
WgHrgT7XlgWxPgj7VE+sueTiQbD7uteYc5/TeK4attxoEphA2Jqaxfi/kcZrK+75
L/xMxa2gRUMAvxdtrOgTMYzK6aTUS5tjAUlyUfEUudzW57qm7ftDMaTlXvBqqInj
B43ttMc42+QyNFz+T7b0/aWIJQQl+fjtMflJmd3sNVJEbqyhZXDcmeHmzluAMnsb
ZVC14Zy/yFvsO1kM4j+WUplFCQUTGFUqERxjjaXMH8pu8f86CJGxxtVTswdkiCel
vcowNsfMcr82MyW038KfKDw1pXeDXJpZy4thjB5gBgOQSo9NuTvsAqr2fS77ruaZ
DNeDOVmHnIP3X8adAs2OJt/f5D7CBuzgSwPeMt0K1SqZyiVPqqf/Qpi5PT31sjtC
Go/yD0y1vYdOE+Ub4PhUZ26eaqPAf54H+5M/GWcZs7bMoXi1Nxar0sCtaf6+lmG3
ZxEvtt94ANpaUVIKd1GZ0Dp096QXwtYn6QNr8tu9TuO72hjk7Yom7F2JUlj/0ST4
BQYZVMpcrtGv0MEQ6H09fk8Yzx20o+t2vOEM6zD7xCZkgiEby/45AsrukHw1CUTw
G6ObXpayctDgstEjP51aSKh9cB3Yx5x0OVL7DIiDmK5/6eh2rLQ/bUEkyxrEfP2w
Cn/0jHooxuUrDUnk6jO+eJHWyST5biZuXruCzgWzf+pdNCUYyJxaC9Ppeb51R5zt
/u2OIBLz6crMa6XvHuafj6SdPabDsjNYyqUdvAz3SfvF26Z5cCzzOrJwTK9pJBf2
5pLeizV0B7ZGO/FYTnQhQ2U9y7Mgfh+De3+RmoMCC8Xx3GgXR3pdzuloZd2lLeMQ
x9R2J51UsnuPEeQTnT2tT8NgrHelifQYLQRPB7zCl9Z1446lKY2pBV6D2dlJmiVy
glB+C1uQIcBhePkmPjnYTqjvQiQF02Txyax5lOzdwzLgLuwl9G6tpzOwY94WkbEq
IjTOVLkn9y7RSSXHdwvBKoVVu3R0tAuHpg9Ie0oZOeDZkbk3VXuoTJ0bjOXe82V0
e8GNlhwDJLCnXnp3iPvL8d74rgd7C7OxAwJBRiovi8CVvx/U0gzwnZUVQZuvfnEN
Apu4hmNTdq47fDcZioN9FGsYoj3Wb7s4uFnWSBguj0pdYCgIJ3npCBEvcRxTqYQT
trVZG4q/zAkyfOssukh6E922VUKXXLibcB23wycE+pfa5HDFj6T/lBhBp7oktcTB
asQX1uZVkG/EzrpJHvVGzfqTnX4yaG5G5pEHarabn2jpw3kYwhpLwwLXjk5DYEtg
wSZCqrr3OzJg0u7bat90QJGI7MHNC6oqLe4XHNf+oYvzwQcTHOF6UV7lU7eDx3w2
sQUVbxgxKfgo2x11yipEEQkzs9eOCMwi2aHFrwYAHx3iJsnkD2Cqi0O4TOXyLqKM
IDBfnz4joQslLsPgKoO9ifxJnpGhbcrZSquyGgMuF65tOw7PyRVT8aS+YHeorSMK
11YC5Qi7BD6zYp6KGH2d12LJ7nAROQ47m8uueRi10AYUcLQqdfyI9j3Y+8aH2XTm
49EzTJk24k0Ej/6Gru9IUAhUO1GEYCv4eJkBUQRT+Li8WRreA8l/SdkHTN1YNz78
h6XzhiMTX+0WiLA2O9fqNxoUK65GnipOcd9DX+yUyXlfdMoBVZxTADaPn1ylw+1N
Wjye2/+ZyimvOxi3Bbjhqe2T69AFk0aOgaEaLhLB/G1/xEYmmCXijRrg1zFRGOiR
I4+EmSxww4OLhJDwJbMgvu2Vto1cJ3OAkBBzi+ZDY6OTQn0sYL5pwmmYe3QuYPGV
M69FRato66Q+yAMieijSA4CUQjENmGVxlGgfG8tx7SKguDdfRpjZwia/GoqckAWi
UTRess4JDEtZuXeZjkvL5RNU0T/K/ql1ni66HmGIVrdP/PeyqLplZlQtNoFXuCw4
pFQezMsoOUK7j9SS7sLQgagtWO2AI7ZFNhLDsaOLs64aoT1LJy+hMMwuyVJ8PnDY
/21zPVpXubtqqUpWl5D62dZX9jgVsB6K3WlY/2pHKWxJm4YcJbRIJZQjbYBawHTF
AEeS7KDzC3dTJuGjLazB3zKDk/AJ1cuGk7QCtdX01aC4CW8Lg48SLby2FR4uFs8w
GoTIQCkI+TXDNK7H7eNaPhxUtBgjAO+IPTwsEJroLu5K61mCFr4DHHhPQVL1MDYQ
wkceDu8961DqIwgb8dscFxLSbqcigAcf68VOLyEctEjJ8ndKZ9ldvVy3VuLT/hEa
tIP33M2ybkTvc7rnFDLTcWQ6xD9q3dPs0XlvDCm/U9xGtgkx0jz6LDI6ItLOWlTA
k//BNcrzTuUeALe6s2znHJBN/gjYz0B/jpJWsUIyd2z0oDwhhbi472PchNYvMRQP
C82Ii0F95em36S5w+/gZb2AFJ8RlkwZ8CqU8q2nVS5vovyJ9ro0iWAw64N79IaSu
Qef7N1dB8172sJWBE5kJnaxvzkDDpNPRJXvWLw0fN71Yvo/ZepJ1q5TQiRdBHIaG
LQYqH7x4yWMffcby6/doWhX6GlxIEHMYsACmRWtu+SJiKO3+hqAgvVRIgCNGcUkk
rJrVqsMZosXWRSvEj58zHg8XHN1ZaC2yz766rlcGbyP0TurKqapg0s3qmydbfItx
8oK6QRXCEDD31GWaBkbG0seQX6hYfUJF9qZ7dqdea9SIAbyX4WTxv/FvARafsFjb
dM7G6koFvj6JUIuPBZouxxHdUzVY9BuNqVfNi0mPMSy7N0nZphZpU/Kq7WeJ9Egj
XBDaHPaKI8dJ88Mr0OVu7/FRFsLro9BRuXKtFDfxYbhai5lfFDTyfvk1I/CW0wOs
RCvO1Jyh6lFMIkAz5AJRTZORPBBRTa14f3bYNvdGQfY3KJpBTKI3zFwsKCcP2Fyb
2/jl1ytuhRkWMQj4D0b+Bfu/r+hBoNInDjQ0V3hWlU2nZA8rq1KLj+0nXejSkavH
J/VKpA7Tt7pHWrBoAjIQFsJFNmY99dnnm9v04Y1rCdglcLMUFllt9/xAnKz7tYwS
U08BobzMq/MEIc01EtzFwBBnazstynsovOi4FZ/wRkYgbA/zmNbMYce96CF0WVF/
+W+QpOTLxcjukvZ9QTtlD2MZpjnGFSOgW1Q/S+s252qHH5U1ivIri/LzRylLuVoT
7MbkTveMlG06Nq/8cudRwOyab0bivbcWUn1TDUmBTZnvYczRuuvdll9zx5veIjiC
+etAN4aMXRBaVEBfLgiNIX9HzNgIlg6LGdv21DL8ZTO4PtosTI1982CZTU77oSdE
4ymzNQpAC4JFo56Y+B5eRRBuXB4D/FN3Y7eNjyl4KNIb+HwWjlnSvrYlHn4QxuGT
54z6bw60EHhuyaK9k7dp5PkD9P2+7hrtbZiDp/y67vsQlpqwcAVU/rfrbbIRZ8Wj
HbZFDuSrngNps1CdAqfDjF204IvaeI6dXYcnyavF5q/N/id4L9lCKexmHx7TurzA
5OeETJiV87ZOlGIJBONZbyRecJzp+KRw04Be0xJEEBJkW+quSF33Olh4MGijHRp0
RGQdh8PXRRvnqQxkw6IHRflG8YUHja8WJPgmyDQryBdgk/XonhgzlcGrVRN+Sp38
CeWPOvNYocRYKASn6J/AfagfcSp8dgeiIv/1olNp3eOIJLuyPFeSkjSxtpLNEcmS
r9SnhzQ289/BGLX6g5P12ig92rmEzYAVphia9EwrmkIhLJFHC9LdMV2sx4yUn97U
2BDnDu6JealO4dRMe+7I5cym0DEIW+vB1rKa4vvHx2YbfNSPRUfCP/tcw3g4whbF
SVvXE8HG/2nK1Vvm2UShi7mgk0zMTwt0eIvNLyyCmNQuu3+VnVXlRypPV98C4Xql
O3Jxb5Z3jfR1tiHMaiQER5Dp2bsA6zwB1A4p9DbzFvxPLRlTgoRFLrK5KERCgWJ8
wgwsRq4gQ+JMIWi6TxRVFiMGS3CHN2TK0c5nTWLt0TjeYzT7K3i8128xmlkMiDY1
xsVeIy1SdM8LGjq/1dNXiCZjlsgiugQiGN+wSLQuQsSh28/M3z2/qkG4/NDd1WxU
iOANF4EWMG+BQGnB7ViDyhLU+03K++yVE/L3HnNnWxKbr0sHf2t4+OwxITVq1YfU
u2cY1LyOayMNAbb5gznd4pnf8vUuxSYyE3rwYBSunUkncQpkE6EGuBhq1J6WubiW
PzBVw3ULuFIIPP44Cc4Br2Z6nmiuhif7nn3GyJMhp6Q8jxT/JHkSRQOKaDBmVC17
KDLNE5Ojpzhi77GnGcmsFxxUITDi3A2EQN0OyGGq5ihSTq7DM7TyHO23qj1UbxZ9
K/eSkMt6rtOY3wSI9LjqYmbagyyECla0J4V+F5ZYJMd1h8mhNUHT5E8ql8hzNwAB
rRGHzEyY63iE7qcZmBYjFwA3la+L8I4FyS27Z+FLuTpM5cW7g0ZoFcGUE2M7bbtA
OeZv7ZXaDsJysiPYqG9BwwDDlHBNbBtg7W11psYcqKQJxjUmncB5AzOiaJYDvHJd
3V8E2yyTJm29sXCFkLYVyoXgXfejGhhZBp6N1zz8ZeZNCgss79P/QZNIHFK7r6Oh
au9FJNOMReLWpXH5ddLTWMu/+39uPs7ZbPZ2l5UWHnHKaVPI4URSJahusuKbbnbP
hvbe5D3paVjHx4Bbw8KhsZH7OzBJFdnYIHX5eAblGsDWYBf1oc6w7Mo18+ng6skm
4AqZo5eJhxvqjNb/JLcR1iXa/HZjk8v2e1GHZyOnFb6OfSUOdj+qiuj/mmS2NUDx
hZ+BHo/IR9IZTbCIpn5+hTCglYCKk23mpZTIP4Rf7lP6W0YNfsJfBsoOfBAxziQp
zDM0/0gKAC49O3uLeG1GxZ1BUz+NYw3JCtKhEmcOgaG9PCcP/4jeVLNxXWx5R80I
qTdPYL5X2faorEj9WwR2+qsW8SOHeqzC8p9pPjNt9zcjr3mcQ5viUFQtJmI3Kdp1
nkFsfpAg0KmmvsBWDDDp4oizIzObtCpKA01Wfgj0ZVtTsi1yjTZm7jxNU51Ufj0C
24997VTQb9LVKlJ7H09A/nagYwC7o9B4giN6bhPakIdL258p1+iY1Lo0yuV/8r5C
G1dmNT3AMMpw7HPsQFpqQT/9T5QnmbZoUdHzLLBB0CUQv4u52RKPawQRDgLSdDVq
GtuuVqKAZqB8EmrR9t4D9d8yXjNbwQHTZI8I+Ym9wPkbagu23YEATKXgotzza7z5
qRC+zTGTt44JLvgquqkcot6042G+D7EIAgpFlPWXUhVMLBRuNpdQbYJP5SUuHeNc
yoUabFtDAo8WuzlyEX/2YFBuOhZCweml4Ha4WrIA55ZJ7Euar7ZT0B7YAaMB0K3a
00Xf8R7YNEsPZZF3kY1UB5qRdJhgoIBpef1wlmafDtN0nMQ2LvzJS2nyLLQUcenV
1uKLUN0LWxxfZIWwVODI6VhaRQXGpaqRXtPnZoL8WDNNWwcDDBRDMBQJ0Lolz0bk
A5Ws445BByYTmbL6M9WDSEkeBJnuaPeEtwpS+z1SyvzICDUr2W+87psxTSCr9tcF
uXTt9qizOsVZAznoKG2ldD1emMFfMOBI26Dte+dth7lX3ic5jKt8sYxSu0cke4iB
QBlfUa0e150e2EC1oJ5x8VKp2d/NQVQCGhaqNMcDR0s4HhVxxBTD4FeAWaWM9Byf
hAiJYV/Bw8uBusruqJe0xHFdzqaxCGsJkcwr3S10GlCT0tI38sDjLSJl6vUFBWSF
mekghwgsP9dF2Zas7aUxpo05t2qT3gUcAabAQLP3Px5hxS+vEsQPZT6T3sjWURW4
8GfMS29UA0ymaDGpUFFAqCikCj1FECNv5m7iT2r595fvcZN6BNIyEoBeM+DLL8ez
AoVl2VrogiK8e/o90WO5oLsp6q7G+I2lQjySSNCOb8J+g8S6yk58qKz1D/gIuc+W
+WwKl3ldCJ1jOZIkw8g9XVe5WTubS9OrMdFfH/rAEWnv0OOob21j8ao6X8Nyc5NM
0yWyyUzfhnCcoYI1B8JnWbtT0MUHwig/vbb8sTj6YEoDTiNV/qEjmDmU76iVCQEw
9NvgJrruBf3WLnyqUKy++NU0Rj4j8MsYlxVa7RKOP0Qo6G3yPwoTc6TPjfzoV0eA
VTNzBz7V3e9ZUOCPgKItUXB/XZg1Tv0AsnTEndRWoJbH2W17XgGuNN58+FSWZjiX
V5iTFgplWJIfme2AV2S+pXQGZRTm+/Qd0WX265rjPaGAk2EShWXWcuAzA2nVl1gD
aACUnZM1D8GNmrVcNpbv/ZRj8H7gvjIX9Iaj3h5BfKpBBO9g8wWQWirUBf7iuHfo
CMkyKHKgjynWWzttNQqomU19dRujpd2mbteGn7edIrp6PHjbeSm/ObYKp0LSpBNM
jkKkWzW6COKL1/A1XzXG42twhYy+X2yJGUJE8+Hnlf/Qj7qtiaQpB/LC6Q9wWW+K
2+/ShlH+yGMcFk9oni97JSRHheAcyFGD4ObqWvOeHUOMiKGP02M3YH7/5HvUTViR
NA0jlq460dHTSH4mzj+2mt+JdpCYxBSjqaZHO4eOB++6DbOwRhaJ4A6tJctqvqkL
+bJpniZXP6LRV8TtdS1q7MfDVwRMF3ryLLNnkjkydTit+Ir4uMoeyoGxFJc9XQz7
cW+pCigSCmpR/lDwFYszOtbBBv5G4CAvTGOXon2L7W7EbJOBA1y2i8HLh4oA3doi
gDQtyG2l1tZ1lgUtKWZYechO9ktL5OGJC7Xpj8u7so+mNmpY9THhyiuksXgJly2J
wRDqG8vy81gi8Nt4uNTArCBlbOEUKEcKERqiKs62uveutY9rzIyJjE/3ouGU+BXV
VlVM0GCRPcRvsvz6a5uRV2Nol6RvHGfQgybsLP4xf/yAKZv4w/QTO9i1r+O7pg4J
Zncz7WKMPd4I9yC4Af1dFBy0Id+9bzeY0jZDiYrddbcx+19UDTVYam+kATSAMnx/
1rbtEkC8OyeGLVa2hBjW9ufTEhMvp2oBPuWHxETsi8Qrj7SsjDEokDGJJu/g+dJI
JsFKIQZbyBdyz5tqlFSeyOxKRm2B03DK+2aA51+fx/q7IOKRK9CDQR1mus5u0SPW
Bmvn+YPxZGZtBFMd6E0spTNfiuWT5w5odJtIuCJdsHncxOZbKg6gIurR2Hd4UA1a
YT7qR83tWmnWzukDLhEkDC8Mz3bU6a+BZqHWKuznyu/NDM5TfSMf1kcbCg1uu9cb
HkVmd0btRdfifl9ztSsZPhsaWPwLxowE+fIrIAmbVNbyPyS/zQ+UWO7EQC79n93V
sdZOAzjtjJlkq/TocL20Orh7EBcT2yb19uUJIsdOdM1JAk+tjtBNQHInkgR+5303
3JEssbFk0vbI6P2p1g6TJ46u7HypQKtlSJ83Ufk1RFfM9Rg2wMcpOzasnInNqXuY
nCL5LpTDTwYCwHOryoA9L45bZvmbcZeMCAfJYt00NdWRffv6EkXJQ96D2hgo6r82
ccX8JdZ4iAga1GaALREZ5Xc9ZQtlLRgBR55Xn1NpesrQR8uqOefafFdTsLI75szf
Mo8/3DMZue/oCoe/35p8TFqdWtGjt8Qz/G223i/6yWkvOB3xj2+bqE44LzkDu6xc
zmkvTsgmG4Ei6A3PdJFhdcVnNbtlYbGp1Xpzkh56XUZG/0r4yv9V93rBBlBgcB5m
PWKWQ32wucMrl7qyKvZJ2s8BMjnSdMKjxCIuLHk1UpjyqQEj8MSpLn2R2/59kZ47
q+kkKtwT/4xTLEMkvRF/DNo9PsEs8Fq8GGe4KJXmpSjgTG8opoJYH30tipasWyHp
NnKOCsX3VemEcnt57wFALAKBuXbsznXhh6mQPEyrljGmX4xajcwphKut9YzEOYqn
syMGNnXW4BPqIMNR8wbb5+l+btpOWN7ISXoLB9kkW2J8Iicjc/AjMadvIFrrC9Ar
ArDBJMQKFqU9QCVsQTnfCqjG3AuBSjxmXP1ChRWWTiUBfRfh7knTqjmmJxyXR6jI
cmZEzZenhNkdm8gJrdIhigfLaz2slcpVOm5koNZRXdincxYK57aIR7e0pqSH0qhU
YtQouS0fKAO4B50JvrAhGhmAtOXoLHTg65cNBM7OxjbLV75ByBms5nohsMckKRj7
0SYeI8gtsW61cSCoNaKfG4kHZPDNNeo/LOOatpXs9fZzvyAH5ALwY+Atu3QTcBlV
MWUHKn7cN0+5zZz2wueeD/QL5d7Il3liuAL2HAIp17oc56KRD6ENCYXZTQRYh2BB
dD7zlCiDzN5xJZDeSHeosAkVUeocMRwbOzN89sMSiZmMZP4LD5R6y80qd+5OnSpq
APDZu+Nbb3Lpd5tywkq4McULSG478ovG2GICLa+0d8Evf1z5c6Y3W97pSaMG0U7+
vqzOCCL3G9ow+LHEIAlsZ1INJKkE1ecHCn9ssKpJ9XGbXKryDbbhUkXN8mFaV2C/
7e2fGqhARc7keeezTRjTvGeUpxP20mmWQB7BmUHznmXt9xW2w7AdSTrP/sEWSA9t
XO9Q4GnWGp+JlfGLtHFYQ2FL6qVJTDXdU5glC/W19fXk3ZmM2HwyI2ft/Sl/Dmsj
keNNy+ldQJeeL++B020/iUHVQsO7KnkSxfTAwarkBsVNyE+p61iyA4pKV1UDhnqz
/DvuQiy91AT7+fZ2hMXAEw3JGZ77RNX1jKx1KtYmhqqUIME4NFU3zBJ+tom2X/dS
uD4gibisbBl7vCL9BSdPXQcbBqvE2gp6tqVbaHI7RNXtCkc5q967oOi0c4hJSXJX
hJiS49WI32o1L/hwPmMssfwZ5lLOJZ6jyWESdtDiOoPj4s0xkM8nBV6AumgJwJ9d
rGD8WU6KT3R86b3L0jd2zvtuitl2WPo3XvxvF8N7VRkK/0Wyafeont/1cpKMPCmx
kSiGUDza9FVLP8HnHzQiD4PglLMwxb0byqNaa5KgPqxf2iB2WJ8Rkfsuo1T/n2sj
YAjHZkMvt8GBvd1MyTgbg5puCbWdtIpqym9Trvrf40LWXZiYDs1TCoPknvpK1FiH
vTb03hd3DAir69H0NU4VcFgSgfL28DIXK7l56qSCCzwQH/1mzuAJR+kbsxSSxOlO
tb1JoGoBJBmuQNf5cecd6+8HGoU9h+vAacruvTQdcRLRR9Zn1vCxhSmtzPmgATVN
urO8VGcTAFWmyQ2P2a+x18ngxMLyxIyMqYc1h4goR/Sc9h75VVqzZZaOJa1/ojwB
JRZjTa93sX6BTaf4V5sIZPQiTlAs4Jty0yP6dAw66NwDmB6Md4N28sIsp2cYEYAq
XKr7MAA5z3C3FOWA8aHgFpGPHR3sNvO9HgvEGIkN+KKfX3/WiYY9I8fn40bgQTik
0p+WAPx4TsdVaczOz35wcg8rO/mobzKrQC1C6NeOW6cvam4bk0xYS2PI0mM/7D6+
9fJjyInwu23jmeIeVPEX9KjQmh04ODKxzUyjBFVYc1B0fEw/2EuQOIs2JbVlku3a
GcSE/qDlIbf3O9nQVg7FV1ilVjARS9nL7afpWnfkOhyhLiGHYv9C9ZVyN8EVL1sQ
HDi3K7aFux+gR+oVLt9M0n+p4+a0NylCZSqLW77AIDbf3pmw/rilttyRo6iTFNSx
wj/Y6CJhTIKFxZjaMmo4HNxxR6mLg9KYv7agEv8huXrYZP9rjfi0X95OPzXV7hw8
Uqn3pSAmcMi1QxIW5oIDTTwm1JZqW9O5anuJ5H4ClYTXmEJndpjYgSPmJJ98yybr
efzlJz1OISwFhY7IgKuTSNpl/iLk55w+cO5o90aPTVY/nC1xNa5HVBuH/gkXFHyC
BwTOhTRYZUMY+cEgrySeEfXPSiX4n3bxGHJYySYXmgAXXjwQSLRrFSTcGUoNnRJW
Wi6S4OiftO1FWSx9G9aInprygns0jkO/udTJpkJLVJIFyrrpT24mBApCcxLOzbtF
TwaV+rAJ/Fx8d+ygC9IRy0IIYAwgk5Vi8Ae6OpHZH04W0eRmNMaVXOFOr8dTM8YV
5YVukvdfNuKRcOgaZDkY1xM9tej++9O5kvb3KagJbx3/3ac0HJgt8V3IAKr7QAG4
F7VX0wu37JsrJgBFvQs2GcIF5TmvKxf0fEtd3vzumkDumHEuOKIXvOCu0/6+oHmP
SaAaApSJTrcXaNv3wzVxAZyBU9jX4vJ5dvVmuMKJPZJPjQtN3maM6czduQG8Rn9h
t3Xvhv+OXLOkhUiRVzQlETvfEVa5XDlfKCOhiK8yOposRHqWUdrAUl1QOYtirxOp
5JnTIkXUj9lgpNlJ8a543ly1nt9W+UJQZNzkclg8tKMr+iQr/xCOUzoHGrqdpzLs
3j+kjfunILHKcxt2k2Z+VN/C+WMO9rbl6euf6l/ItpLRrrgNZaleuAHYssLt1oWw
b8W7BuqaWDpqO2SSypIJOh5iYh0KHGHiNYK4Xd9uMJ/1Cpj8dESjCdo0EBRo5zj8
Enpc6LinCNTzt+bNu69/8k4HgV5U8Rc9LnSGJbMVRHkIxSRFTvUdU/r9VBdWjXNo
6PzZAyqSA/TKOvjtGI+3h1Sf1ENu43NnFQNu3gsblwsFnXXKBndAOhiU6v50J9y3
KUUWkB7Ze8WCT01eQBN+1gHv4Flcv/uOgrZzVqbGL9LydrM5S4hD43vA/KetYhij
QAoOxga7kcPiXvoHunP3JAhNXP0YOGdiWDoUX/uBPk/gpWcIW828aIffWy+E+3hi
bFkiMX/c0Zwlmx66l1KtOI5+lSOiObOdekUh7oZvi3VO+UvZ3JdoaWNHSFZGAkJB
x3692vHbm10kIwQStg+4J74Mnd9T9fylBFZL5ddjU4pcX/3oaf9Td61K3foFbePO
oRi1c19Si7NnwN84QsAARvJioPMwPKn8q8y043uDLxyRCCh6SqNRGWVJaOKxxGFA
DHvgQ/ggOQUECD6GZDglW4Ryis2YnOQsJJkBX12b9pduu43AGofEHiNKNqW0s7Sj
YBDY8HxNwt5wwNQlbxSjs9pqcnEwnKKHnPMazUXzGkGOFgvGiF0uCx0vE9O74qLa
CBdFSj7FrjxJoaXjJRvC/arL8nD82HRuKHh1yiYYppfIcFx41N2L1Uu/stZC6S8w
bH5S5UxXQ/jiTdzlPOtMqR9YOWfDY+D1YcDrI5d++jpr2b0wQp6fN+vDmbtzJclp
g8aACgRSNzVu3uNtqrpRvYeWQ1CZ/Gc3KRDcO0c5o7Vl0CCFlJuySEDy/qjacdgg
Ni7yUiQWflWdX/T1h7+HmKg0WCv3IVal1jFs7zbsixU8hdkPU7gZSeBeL4HcqtY0
XT7IsanhPsRO7hnllXFfZduuyywtYNw9S9mZJYZRKBge/TKR14iokMtPmtFjIPLO
T7ss9jmJkA3WkXoGlMKTCnu1wMgk+Hce2V3Rz4QNYCPj3r1lWKJ1Ol9RWVr06IRD
lH9d3m9Oa7tYCwXSa4b77tvGCiYyK7qtbCM0qnDOg8mrbaumbPvUcX1bTRdykWYC
Im7C4TQ+MpWrVXbAhXgYtiy6DSCPE/G69VKByN6jIGkjWZAp+twT+sOZakHKkstg
ue/F1Dh3Sx7OPw1narz/8zHYs9IdJHWS8IXy0F26L2A6p3NAJvRHRaJbPAp7jZR3
UOezfCxqROe1h3EVr72IB7v/d2bgMCfRDFhSGxh3tSigzmpSKRAfhmH3xQE3iAY6
rtTmDBtujVWuA8eovJoFyUocoYEM7A3O3EHc1ieQZgJ0NcSBsdv7ak6vDNCw/0ux
3DmLGRP3aTFhTuUCu0yuoqg1gYsjkMPNJM3Wg3ZdteISTSpvlkO7mOG7RJMDsscu
dIGnuT4JWjkknii/QGytNrqkaKvdthi88dysXMvq8++P5XoVElzNTUywoH0VaAl6
DSkHO+DMoMoCklsQXjE4UJSHUjUs4kbJ6PcB5u5V+aSpbM7Afi251Y8xko1eifZt
TuyGyq8OqluTHkCncmV2MmkYvAcODpUZRsQGUoiIxz+mauz3qwZ03ULO5WTMWNOa
1Hn5bj1SIcMcJHAvodejdtk1UhyW4NA+89zEqrIeVGYcNmcmZy6X5deQSHlUajTa
OFq8WJ5qtucfFdnVDkoH0goqZK9VkuXWY+Fj5sGhN7oK0mCrZ/BdkWDii6xABFac
HhKlsY9WYGC9+mF4pe4oAKa6waUQnd5yYHML4mkHbnM7fFASeqvUscSh6G39cwii
YF5i9DJ92woaeetbTSqOaQdrKmkXCLRDeDv3IDkNsw89AdZObFQXb9i31T8isaV8
2p/KuHq3CiY5IjHm4OPeOIrmdTGHvGJKo2CMoK+hSZri5fhuP5oSNGFEZSGw1hEi
8pjyDPxkvG8BvmHxrxjY4AoGpTkfWMhIJkTHP7HmvoHLrCG0TGXaJTuS5xZQ9g3F
zi5WHb2dqp1lv434kf0C6omVo/NcXU6ekPShKh5MP10qrxLVR1kTNKPI/6ht1Qeg
nacdkqpS0qJZe8JSbsCPWR9PU60zQKP8hQVSZYSSTj82aH40/q+jvpUfABhP7Zvq
1U2xiyM1OYgvR606O+GjwzwGo7wmAaOC4ow/9rTt6oloeZNcnjXXkXKmj0yfE24Z
hFVuEBoll+yMARY4bOmUFh9RtCq+E0F/38QDtMgNCETYQr2Z/bkZOt/jEU2HBago
6ttt5ncb29L/4rzaGZ/WggQpyodnYJqEQ3pE74uOdfb/xmkQFw8UJQ59wdIbE8aI
jOq0ci5uZhBLD2HX+mFemKF38KAx1EY4t+ueasYy0HswHHGZ/Q5b/vgm7RITKRh/
puP/lIKPxf/QCE09gn/eShZ0B63dPVMbFtWXQo8TdqI0sJASnDT86QMA95y62Z91
vXZsyeXXdOTuVF3h8knOzUfVrk6XBlaCQMvQwGZyw1VRffH1JUSMJKimzrCHWyuJ
Sn6mtpYutsWsaI0ARWuYbow+CpxAhKFRPVr82ccWXEnsseYm/Z++e+1wRSahr7gV
xiuSoIUnyX9bxA1C2gW4DgI5FPW6SnnQqKP4CuoNs9CMuZdmn5sj3yHntdMO/xG7
fkd53WwGeigRXK95j6tDHSgXhiPMGOfNE9z4QCf2a71u1Jng50vglptoNJ4vQwWE
Zp3Bbb0KMI1eL9MClSK2mEdMWgJlZT5HpQkWqV3XYbf7lakkhaXkJh5TTYkyhRwi
nWcenYbOHzLdHQkj+cxvMgbMhxZgdMzEsC+dPsJ+XlLBAiKGYJMk8j5A40TsPv71
/30PNyJ+F6bMrw/+ZXUXAOOJ1q5F/0Tno2atbIBdD6zQ3rQr91ZQ3yn0QzCjYW0T
JgdPPdIQBMU4HCWyXom1Aprpi1LuVjdUDmJcnG9xXMzjgG8bXNxnec1OHoU8sla0
tqpOT5udWGt1QKq4UbB1XmxAeWII5eukXsWjo7Uqwiv/9yg8rXiKKxFIGY7jLhJt
eEBWh9r4MkGSSHKu+5Ezf8QpEPhJrfBFvp0NYxlETCaZs10SHxXWTvHa+3uevjMi
77MuSNfwcgR4UmQGKYcjLJVcdGZ2096w6uJr+Gsi5GVViPtKj//ANVKNbglNCvq+
q0b4AAPqfqCoSMNlJ+oJhF6Gsb/9Tig0AT7dhPRabnGKk3jFHnjf4PCp82OIbYNu
iERdYZRYscBAApC8daAtpNPcleTvNOzxDbAvFMdXxkZ2eXSlcocHhLQCpCmnECAB
dutMsLv0D3BdC3zkV6bT3Y2B6c9+ke/od55IHvWLPKMXr4QUv5GoZGb0V3v+UIoR
yBltH1ikZi8ShXNmMfZ5e5qcA0GQwl6WJBtdvF//HROyFk38NRUknx0jc2mjiCfH
qK67aNlxhOi3+/3w4aCmegfYEnHbjoNEiFTAmPk6mQILvpnnneCjakuWv+CHORze
JUOl/9/kajOZHYW5y8BT0gBMleL3sbJTiJyGXSMWGGKn5FEgIfge8AXfPIn9sVBo
KGKzK+jvB5uNIs6uYb1qeYfYKzLaXUDNGU6zz/wRYkeI+5odevc1LUn5rpEWMYGx
PW9tb1g46iCwdpfpS5XYCA4KKBDiKZTWEMvwqBPtYzQzmBfwXJcONnyaXZj8lOi6
KiWP5CQ+rGrUPcrR8owEzoox1C9w8pneHs22mjTiiRxujkycekstyvqsaB+ua58Z
K3nBVlgV8K+jy/MCw86S5SlxEbnlIc9bQw905TyHUkgg//yfvmZk3rKabwx4yMYT
TXnla0bbkCiDi4iTEKrWL+kavgSowNsA6Urnrjd21P7cfOIaTkeNYi7to0RUP3N4
5YGhYUDB5NX2f9ysG9k/BhcGIFBbutRTeMDwB1Ejk8w0evZ9GRQ+b7C5/o2Zvtw+
6yA3VxiD99+foGAh+xZIBq0BkJzy3znoRrigtbFgoeXPS46YR1YMJEZZllrx5rLG
j9IPe26hPCqGM6oSCaOEJEO5jmJPuo6QFMheRL11aH/Cg2yR4O8c0xGj1TnODLnm
G72VOJ69r4UfbuCBWmU5JfIXll+4v3ck2bQdvsi+1mbpPjum9hIO6Uqfp0YdVxUy
XmgXbs/YLW1bBpBIQx6yhh0uo5rdWihwgSBIXHweaSBaZd1o3WNVsdd2RWeE7/7p
huPNqZVNvVSk4zJO8OKuSZ3SWZvID4KH5tHB9dZclPOPFdTShClKP7Y9VCild++K
qun4QlC4gnhkKrqHZTqZ2JFVhg3FZAdnnr34l5aKStBfo8AkDdp5BSWBk0lWBlsn
DhBsE3aRbuD77sgWEbLY+tStuJmfhQMRb60xCI1tOBsWOoQ5IsTAcTJPO1bSdcAV
wN4yEzs38HOrDQX6k5RrWu56FjFStn4xbdN/T6soE8yMNQiO7MEgGSUBUZXPFJ52
Ozpj1wAr90hhJ3gsvaTH3qHuJNORHpWSTFujmgbMlY8B3F/Lw6CMtgLhLVJEYQs0
Em9ZICuE7wDhpw2nnYpVWp7JyK8sFdOSBS2KwEtEIBj2YTL7fVPvRjbuu8jC0cFu
1aZJc07Txx5U4zZ6yJ6jyhMOz9acANnX5nGVNFg+yFN4XFBxvqJEuLG6zSXpCYlU
wyp9oXeNShqCUdd+mmxPzsU3M8fI3qY6t0bJFjsj3PllbL6xfZWggEQwoDINe8i7
6KrMaENvdzchhJvTH0p0gKpiE1ihuUvewjZP1Z+suWWpa4+syoEN9OuEkc7gBTmr
WuatuwFNDrpmKPVJ7n6Sqe98poogp59O89CgCgMui5gFINxaeupZ7dPBJndZLsiy
TITGfLJtvKhRrR1UBJl7sNHPokA0dUf1CRjvw5CGSIAgZOrdvqRD+qbF5jIDn4rN
PMMJkAwWSz/PMa1kAB2JQ5kX2KIUy21+KLDj9faQDpQ1tPMO+nhsCSM2UuzGCbeW
H0AuzLtRZJ0MlJhhIR5fv3ZwSZlaqCX0mbFK0brM6MpItXAlaBIpVxQOByRAr3ES
PwAJ/3Az2OS6VJ5KSPsbT3fxeSPgi1Io8karH/GsJIM85SsdUbF2Y/hYbjFD8Rg2
36/kEHCNUDMSDXA/H6x75IbaKT0m0hz50q3DHEp3tdXey6UwsberNUAxNTgeMiLn
2qw5Ysh9PUrngLOp74L1QfQNt+Rx+J9lGzIZVvWbBRuIG69XJhq6sM1KmHGYkg57
F0xhNs8A4/ogXAdSfJl5iP8FpWSqibXZnkBCl2f2wuRPYYpPddFFfyqWvU0Ws9Qt
QTewwf0kHjnsr+ksQnC0CTvWa/M9TLkpOlTWQmTp/ZZVdzl6X1XlbkvT1jV754Ie
d1bbEapyoZqH32Le5GIDysL1vcvY3EUp/B0YrgqW9joS4WANWuBgKZ3jS2j3pANg
pXSj5ONtNwPGeEF2H2PZX1w4mAvBEJchp7MMJdVqqqj43EOkwhBmyM21qp91O7OX
6+2ufMxz8lewxTd2TNvJpqnbnjy2pwzncxunf6+8y5++yuTTRoIWkTATM9KbMmbl
BjlDIMR/tlynTbQukdSPf+XjDJFP8V0ztwzgacJ/vfAJ+K5vJdDFfW4GuF0LYZg8
rwyphL/3l66vX5hxxiiCG54LolbI3pZevcMv+/VkVG5eVH4u9znNyh5z/AF1tiG2
vhcBEkumZZOu1ZrZK29KuLn83iKKMQAzfaeJfbkSbVZv4eZMXMzfnOUuWtKAr8sz
eOBXmw/0ZAKabj2zxcXyiquQmYRhBUJtSWi80mBRqNrMO36g8BygfvEAIzc0r1CF
OhiLq1YIuSCjrqOZATlDXKe1SdRkTsdhjxG6TvDE/vA4a8wEW14B+qaT5vq/QTJx
9bmsz9n7RbpjZM5YmrBjpp7ouNQ5GbWr50IeQgPo2KzGFRf/oc9AensoomYc9pLx
kJUorMk1G/TCAXJr1aN8em8k+kt1vcF7hNrRC8QhMI2svukg2lc26KhZEubRG9JE
JyWI26r26Xn09fqBt+aQlCC9zGedUoXiywd4C2TwlY1/yHQfuvTOkmhAnVD/4CSF
EBnvH21RS/2MDp+q6h1QUO4UeURsFpcCe+VKcit7FlTZFpOdiYFDu20RNAUTPMh5
Y4A7yfk3T56b8/mY8bXitvmOMUMkLbetDOxb76KPN5NCPw0VAsniAV7nkyJ1EZ38
K/ETKY8EEtimHJd/v15+9BK+IJImkA3TWpsWVQ6fBe10f9KRXWw6MEbwY9/77fIN
H5i7COXQz3zdbQHtB7Oxtsxtv9Yx+9qtUOlMqy4t69SoftgQnxhJtYC23uZPcgR9
bRQD0xQ+WicFwYLStDmLITcE7oxxLjFojz7McwIsHLcsvzrF1txzLxkDYJRb19a0
cDa/kxdyAQFjLA9yYpdiWE2+gIFWyC3Ab46rF9uNoq6IN8nOEwBH25VNVIwVyfpM
rRwFQT39dVxjLcEQXTLiPgXEcTAPisP6Q+1Fv2mnXwk0ohpQ4KwdoYOAAsi8Wip+
5/3DaL8xICc7xhdWFlwguREuDP7ZxhekzaG0HbooE8/P5hegHXkMH3Ke0j/H5E2s
HDBDeuW7pO4nTDj59w7RWc8fY58E+xnzKblddiWXT46wwmYxYIplz9YymgHoo4dD
Tncns/WinSeuEgqTA1XG7vvpooCxVXPAJU65M9cFIrbAE3aAxv2Z5VXyiHuCbmbM
vN1FeDs5A+u2Ne3qSElkv6QDwtUt7+ytgkORXoVvjFdBq2MH2R2MKvNNhjh+zXg+
F3ArddTJjAzjog9NXaNUMviV12VGK3fV9JLvXcNO3DVWFeVAw1dufDnCwaOqMzLN
T8DbSttWdPRSMGYU3h7iEqnCEAMNuXGT1Cvr67YnD6K+R4a1Hy9BjL7m5d2sG9Jr
eUanDKQxLvvmrBzliqUUrq11HskPw1fY8iwYonAgp3u1ZlOH6L/cPG2En3ZQ1Zvc
7JDcTdC3RYk4gD9SxqrjyoxmsKZDJQleCTjdSjuCe3Y/GFjoFYN8KCksHVIjSJmS
VeUkWEWAoPpfULobkg42o+EYEy1JZlK3aQW5tU4CieAVuvRwbjMcYXBySmxWnlLL
40Egui64/wYvHcd4/qz6Sv/1EAVa8kr2bjiS0VG3soroHGK+MSLWRVkGEW1dBm2R
W4F9jOTRUNncEQS7QtZAF66cKMngI+sPAMzF/6+7qFtrZuBT56FIGTR11w9Rcwkx
pRxJ5l7CcikPtyk2WamDcwYYJEyeq5SujI5HMd6IfM+eiboluy9BgkQ7vK6bnrCf
pxA3Wiuf2CzeallRrEC3soDU6daqglWWnoOmrCxG51nGlSagvH9AKUkG3sv/SMQ5
T/YTS1PIm+vTZSd7gMOapMamFHI5Oo/HNVCR086Ikca+g53VQN613aZ4wU6a2bHH
zVm8QG4ZsEpAKsN1oTPx6Vs1gS6f+vcsWIMDGp3mHRk0lGuKevSVZf1ZWY52B26W
yJ2Bijwd9L5D3ngzIrNBkQKmq1VVAxeEMoP4dIrMVxzYaP9ac8e/Z7h/oCm7nkQk
SBZbgq4Hk3ZcIGP4UePeLrhSWD2OluLAsqi76rXrZ7+z1gS4e6FX1TRuVEc5NGKB
ApWhh5ft8A2cDU7xIj/t3qISpN0Y8GApcaEuiggGRHCHhxjeqctrs8RpGKPOyAnA
EkdXbZ0rhcCPVOxrqFWbr4r0V/b7eq14fBbjJcdqEGUZ7itfT53UeiLLOOUFq9EY
OGWfFLdjfuA/0aORNUElewtfvGxgtDIFEAM1V/990QHLNlmXmmYZuouoj4G0sPnL
p0g2hTFPV+L90YHqnTfpJi+xX7ZpnqqUHT5pYgSzGLMMcahL9W3BhN3grFuI4MCS
l7F2AeZvaeLT84kZHs8zYxU9dPudNTDrlOYHhgPfTWegRMWXex7yZVwaL3nsAfci
miGjTBo/Ms7r9lfkk2ETEzTqhdzDevvCj/HdzfTw/mmg7zQbWLMSlMOttB7BoHJp
VO6PHz7ZmdEg7wAOimF5yhdvlzfKgNXSP9WAdTiY99LTaeMI1uM8RM9GGPbX4KVd
jWqdAdiYB4/3kk7X9ikFS1uESaWdFXMOHFeQjfbOJlVS+jSKTdqZ03XobZMQKPk7
/dT/r1Vpr2YFyu6eJvezHsq6BSFL/R+/9MJjYHJq1JZfFB5bxoNjMbri0+Bd9B0Q
SPMbDdivpuVMxRnhGNBTAp0RVywHOihySyJRjwuC+NCLhXj8imaaJchM13mjCUt6
fNRkWB3qIAHTUreys79Co/+Q52psfgxMcFiUeuCEHcCyQLCWlE8UkVVHlqrTToR0
vz1fXp9ZAJSeaGWYewX9mkxnt3ZeOtXIj/nPptdw20M1KmxrJ7YBOr7WPYZ91LA7
eCPWIGe6bii53XaO7IXfc3Im0CggWbipz38N/x3o6/38YNR/Zah6+yenpSvfsu9Q
JI2khlP2rtS7Qh1Yjyh7H2MqUAf8FVpvYjdYVSbs35ei5Nd+rqLS20LeMrueHf5A
81xV9/X/8SRbNrwACprUv732U3UK91o9MZs8RA0DYRibWu25+Ue07xQpfGQPbXJu
ZxfEWWX3Skpl7Q4MD3nMYPhTfddPlkn2VRbsKjDPHGZrasVnGd/lYdfQG871BUir
DPCIZ447ZiiEWon47iQ8VCBckI/GP+7JG40FmdLv9o1COLaTLGJgERZSc/LQxGLE
pYt6FBA5FQXXC53iWPZ9eBIiw3PwX+xJzASOXbPWXjCh/ggNVutleVUfabuoPFd0
qjV+xqLwGTY2xiCaJzkppEz2iD6ifW04p7z6P9iNcKRjG1a+T+e+NatifOMKNhxg
xIY6Rg/6ve7jmWrkMnCN4Ks2YmIqIczJpA4Mk/82a0Gtn6kTB0uEjTTYu8558P4G
eF85pwVhf/aU9ASyDUCkpeiIdEScJqmXjxOTART3BL2QTE8NBxw7sIWgMEGkKIXJ
QWy6B7H/gpfv+kIEJApdooQ2mIsXU2Dgchi++zzaYfu18B/DRMwTblQL/PP8moRP
FtPhKJQtkV3wLli/VI2EtGdjVGRtWsIrQGl2Dk6StsP8dgfPiRZPUGxdeD1CS1kh
AyBy0RcmZycJIBQLf/eWHN/7cwhKyedcQ0v6Cb+affncFdP6ZlKUDYEHJnxA/Y5t
HhwFF1tZTgs/BuhDRbskkiB1hnuA7PRMBpOJLOq5QPfvr+0oq9MSH4HgtAM+8H9G
bpgXhiGlS0cbxB8ZHvM0r4Hk/5f8aL9U6CrDS2lOd/ObA+Z7IvAtgSMAXoSAq+c6
hlWtYDclsCqVfIYESElb/CIrS5x0XJAfxwcO0nTXtBE/axSHFGMo3WtOmtTXV42e
h71OBeWqu82aM9dVlK1wKzJxol0Ph9gAQMyTL6QGDRT+UmDVsB343ppD61kb1w2P
XTwzqcMIkZwaPetZjTyobIbRT0wlH5EfwIq9M0NrW5tdP3XokwPa64x8dVaMUt21
fvbgmWHGQINiYoygSWHUp4+23EXKPPI/RE0VSAzAPGrqD/frNLti8xnXLPkUPqQS
rYkHy312V0BmqrL0DhcJ+ip3s/0tgPgprEOCkyaAS/A3WGaGJ9OG3kFps+RtsxV8
5fLd90Nmym0tYwGVk5iopFmYnSed7ixp9898yErtUYgi1+B4vQh+DW6pyfxC+Hx0
3mqHKDnIeO+my9fvWR+AEX1Qr1OCGJ5fF1kvSehufS2BuKBYLuVc2D2v+MMoYlRh
pwStVOx+OMsw/iZAW74B59mLuE7Ylefj0ZWseEWyhLR3HQ8eVfyJUI0V8KgqhSTL
Yf7Io1sOEBSpuGDIMg8gJbG6n4iyXhLlRevhL5hypxs4JWWqTIXoubcYECXqXifT
T3LyC6gpiH1Pt4pqYYSEs4hEQtCH9y6vRNvwCo0Wh+GWEjTwP9J+sgkQ4OsWVc0l
J63jWKns7ANzliiz8t4uHUHKsBAwkdZwLU/US/QRnhVTcgNlMbl1RAszgRMq2ujt
DFrhrxlBghegqCYzhz82mUSe8SuS5oN8+gXV0ec9JX+dIfhEQFfnzlqqZE3kSUOA
v2LWNTHG6DzInNIRsfNxLF2B6urmclELsAqgvhLM/wWbCghPkMZ2ZAKkdndzomai
ZfRKCbHe/b36m9uXfznAWHaFVSbc9ZwkPzhGeE3Kdf7vapxi2slA8CJOEaZfnuHz
fvAvRzkKYwOln6YECMcZw/06GO35Mo8VBmKn0I8Gua9V27An+Mb7E2qaTw6ZTjlS
2UIT8WqM77ru4Fj/Un7G5Zr1qjZRa5WHderJHpU7LEmHBiYi8Dp92JbJSKjzI7I9
/bWNJY0uyU45c04d6vS61saezKTHnIbBmE663VKnnjebEMVqg+PMmc3tkOabsKvl
VENHd2c7mHVsFDEZc6BMWYxwxAYqupcjAJbn/bmWkn2M51pbm+BmLx4KlsxAcFOC
XUv6RCcWdVHD6jE9+cIM1f7p2Um/uQbLxJpu1nqj4m51ewj8JR6cARnGUXyyHzNS
seDOCvAuV3td+BOEqhI5tgC6Mst35/xQvmdQMSueDfY7QcH+wGNYxs2bdVkC9wqU
fb7HdVNOkGGYrq7lx/9AVYjw4dMBC/fkBErXXj5gzgO1o9n6B/qELLcPiXQIGTM7
LhmVxHzvPu9NcDNCEDQFlBtAiKcCu+gKobjiQCZkqIxTss0llFoYb+2BxpZUFaIy
IRUg5dtUQF5GYmL+4tKFSSEoC6zUj0xIV9mp/zr6p+JW722bztCLKhC7rUx2JWwE
0X3jYs7AdmGhhdQgyxUMOzNbZLfwTHzTCdtY38pGDwJEd4NqDABNJrubybJgtYSW
yvBRdG9HPAJ6Ak5JiavtR7pj+c3KjG9kVtPLt8iw7bCjoObhnbc5cQ8p7rvwvXRG
yacYwLeR+3guQrMrH09ixrImmnP+gaoS48FDGZL0TSRYXEYiifZtba8D6J8H7s2x
yXypswNmr/axTEbFTKCcweq7U6fc+llT4wUUh0D7797RYCUhAHxEQ0PQ8KtRxrnX
qDpqk2LFNTerNpUPmspYZph0gLeN/mJfZysCgG54zEdrFyR8G1f+5vt0PQMwKZw5
zNyh6oejf1G8TRwR8q5rvWb2n12rGDnnbsJpW8+ZgLIoACueTb+ZhyEHoBKMl8F9
Z9GeVNMkv03yLjbWKCu1qJRyvULQPO9jx2MCEZkMqt00s6vHKgy038B971AnbONZ
FIdq3IhzWjT41U/y0TmxcGBtmgVU9FbGbLtfKPeHZ0tVt9ggm4VKMisxiSRzchPB
knD+YLDe8kA3J7AsPmT0EiCiWdeT+MJP9/uVRPiK7U6BKw0gitWM0ONVv3tgZEai
xicScdQ5lNHdSH8bRBBELTQ0z8swlLF/ovoSaiyNCfLE8aDLBG/q19UqNY2qL8N9
8ll8wqBIOfjP8L/7Lh92Elhykc2HkfyundHo1dtxCMT39gGFOE8m+huoorcazvXm
+nTSD4oLYuA9uRJBEzKI56AUJd9dSHsj8vlHEbKKW4Fjkp3LMyGjeteZcicTiShA
7PE0YJccZni6OG2u/EWgrSCAT2XJWRsXe++xudtFnUOVgAeICUVTSu/CCr5HUqPl
pkUAq/l3B7W0dLUiuJMEb3B/eFq2dVi/1xg4yozVNLufMJaRV3JAZD5b5QJ2uEk+
Geo6bFVXT2kHef9TMhwDG0qZI0cMKxtmAWAED47S3IfVBtm/0CgZi2te6kqn9jZS
ZKwDWf2IFHfNbBaZaZa+12P/LkUns09oexeNKmVF/gMp7N+QhIrYoK+zHGGRAa+o
oZiqV1eDGRQTOyZfVaPEoyoD5jC7W5fmm9ADHzMkUPW7M68ImT4iCPVHy86Bun1u
PoBNi17hB8c0gnfk5J4t1LxBF2Y4VEorfM7rdiIEgMQHNfO2O0XrONTRwlxyjDKN
Rx5Bv1oHzJXQQhN1qdKJgb4BgTs/UsJb3NZb0zUuCMwNs5sXPVlq7/Cm47X/jSLE
JHo37cfRpDMLVPF7p4dW+ulG17lHafi3a2Di7OKlXkDmFXRLcLzhGujulJYD9ZJP
nelo0sJnomhJMU6JDGUz+vgNKtqQRk9ohHX/sNQRhxyLJ7FWH03gp90VDDKkNv13
8eMLDj9REV1bFwfSak0G9TbBDRmRH39zYFRjsXvJoam3vjUT6vyhsZqqyShTODxG
Y1YGJqkocXm7zPH+nbmTt9f+UcmXl/Da58kkET6N8lAxOoQYEpy4aZMSKNKMvPON
tSWvFHMi6+gw68kQ+AnOKnW+OqQM98Z3iR5W/HFHKsknULOP03PfDtPbIBFYL4NE
CPdtZM5cUgHYxLpdqBE8YLnchhjTPeTcgTY+4MyJmaL46mYlTiZvFUtIapZ4bspF
GxDc+b5Vo3nsCYGoiJHTDbIbPbhBxvjl0fJnKFqg76kAkVdQ807dMWVBDRzpFo9F
KuzZ+P/guI6gQXrDgkCajXMz2xc11BiwiyfW7qJB5d31ipOXXwxP+JVExaoAspUv
A4wVwECa9VAlESbR0ZIILsCaCdn6TjLn6/6Sv6g0iwkL2iwrqTJOgHpZMazQnZOp
EaQZqWn4yl1O7NmMKAXvabbJc8QvxqWtF3LSJwlgi810rhuTBzsS0P2/meB9VG1H
4HHD6hYhL5XvQdtkNRR/a2pNWhjbUvRxSATMYHW1wvsxxnfKDe85D0MjA/qZUAKT
nAIWPmOlZVUUs0NGT7zGsEL6GN9SiN6m8NEf/c3YABBAjRi8Kr+W7jyvUo3ki/6a
AmklvBi6CXBWqWMXA9vjhO+5fYrfaHEp0pLr/TIco+ergjyyQ8wGmW+OqN91EMyy
yL4gA2gDuBYgiMVwQiuZzA7DEJ8VtJwC54ntQf+6ORu4gz0Uu/T1BwtFC2z9Dwwi
4fBo8oTVFpR4l0sk8BhKjftqHFEibmzBg8Afd9fb9hFaqWaQR7E5Ai04yuVZcay6
8vUqfucF+3pzxNhtM5yvPOpFp6zYVwTnxVjQh1DTW7hSOEuD3zVeF+2mF0B09BWY
PQ5D2GL6GRNXZ4wuUOfgA5PeRCyZZI8QjtNG/g2XPq7ggndc62OEOtxpmRWw2mOx
ImDG3Fugm+4V9KOhsOxfvzRC+U0zfTrqBTpgpjZwKjUkjvgD+bKuEu/dUyEcaCIO
QCCM3O5IBNNrp893iEnC4i34OhMt9SIlTnxYPFk5wf4BdbnGW0TTxF6WVn8892x6
U7/F48xm0HgV7nZxEkoay1dRvXpqAmAnK/W6u6rK2ffZRJm3FzSBNHhFaZExOerW
i//7WIW2zTFre/OU3GCXiitcaB1L2EUZBGzPxGJv2dykheLEeWlc9uXBpS3ctExt
6OuzCXPoh61tb8cHQ1gjNImH6aVeKkGA+dm4XFGwS/lgB7HaHSUglQYuAQ/g/gU2
wccVzek788mVX4T4VcfkUGigo35/7N9qB/jhGAN7wzv3/0V/y+mQNZhtHYBFFpAU
/EaD4gRAzKdURYpNEJaw1jBCqG20mYeUiJt+hP6zIvaBfoJqLlVmTBXf4ppB1Brm
+vqf7aJxOW75EDZv/5EaAshN5RYu8vKfrAZ1R8C3NJSZubhk5rI+wA8EQfkwKUJj
pt+RiBAO7ATbjyXe/5EY7qA0aIMe69t5DZAsQ3WMHwM6r3v467JemVpm1dtGM4Bf
N7wj7EQHPlc7tt+2B6qAD56TjhnkirqPYBkb0peE8cIlcbGbbjJ9pebSxfi4L016
SHd5suJbRom1vPf+AdCJFe/Jl/tto54NLtIMR42jrYHzpF5UywswXBBOaQpVAcV4
iXcr014aPF2qnngxDCspx4n/hFnsft1CEyEFLSvy4imVal+NJ4qRq3HADFcZvvTh
kp0FvaO9PDWRrdYve2kTkbuN3o4HcjSD/Yrgg7P60ok/PHSJm6ewumRRMyftwLqN
miTOXXddnCeX3eaHed+59rYxGGdq86RYctRoALiRS/DMZ/PDB2MC5UGM496QZ950
DvGEyDtII4tMaD/rCLlwSCIWyR2nHJiAft8a+NO0j6YdMAJWnvbzKwbOPZgrLZ7k
H3F647qYWbcVeX49VpPmhxRtBonpTn/LJ7kvd7qbSRn00L9IV/B/GFDaxctyhJTL
0WGSckll852+JJXhP5wx548bwclrZoQV/24jsPI1LrzfVKdl9x9aV6l3pVuJlbPa
AZFI4FE8VOyQDa8RFcNG984/FthkCAc7x6c5daa4c6uktafUcHBsB2MsGS4ZAvXv
R2o/4d48+iNlusB6OUU69zxkZiaNxi8WbRcWXcUww9gEoQX2rNJFONiKZkztyMKp
xaHtXnhdSTZBtTLHtxKPg8LQjeDEwxGpWKIQDdMQ2qqUzfNbqKk9G0TlfOYeO2B5
nUaCZ6Z65mTtVxmHYnmidtEg0zymiQjogx3SJZLIr0oMaw3aTb8dByNqUJthrUgs
gkSntVYzsr128R5uxfm0hcoynTtIwIEDiW+xL3PaQmHxOwemfOjIrg8wJoBqjDoT
08htaqhIifHl3ZNT7IZrOzQcJCbjIOYtuW560E8Tx2BhXf6hh0g4q2nJovxyJGz3
COrU3gzDpjgswpPgiiRzfytRHiJiYO3sYiAuA+kAJpQVvgAN7P/T2pLZO+GxOhCl
PIEq9Gy2dzDf1OK1WmQlXydmdL0YBoUQNBoXfX8CJ6TnMan3pvwpQ4h/+y2C6VMP
Hman8o6gaoErcBcXHIIpxgpjSGvTUbyLFxzHSht6Q4Csgcpo/3P7xdQxPFE8OFyi
U6jRY31J6zOqVKk9gbwIu/B2HVz3lxx3r6e9FSptyxCPG6r3AwwPTe+8WZVnMO6z
kwWTZfCSkUf/8j6TsFMoiVHxiZM23A14BEkOziiQFdUmRvZ7+OBn4CMrGeC2aDcJ
ta0W5v00LnJNYeG8poZuzl9EJ8Ef1+cFrJay0N3tND5lAXGa1DyhEWhBmvxrJOQK
G90MQfhgBwSoaZ8Z/hBBU/Xljuj/gyRf+sjwre6xLvJfKnTeVyQE/zPZVtgU8fwX
i8MuWFH8wGxlXfykR1Ptb88h/sVEWklTTkXYfaY+btUyoOJOvnEvKy6DuLZjliLL
aovM5hjqTc2aav9X4HTPX5T2tOsNO4Roj6O6NZa3Z5ZHAge8d16khyMshv55ojF5
Wo1nxnFTbnKu87Diu4hVHsqzLr31fVZgKYuUMKWJDG27/ww0+X+ca/SNFYIfAEBA
sd8zguumF+MnjcC/feVzjeYWVzRLjNHOWpGroPHALoF+BVST2ZcHrs8j9AUBv6L+
nXCVQE72JG4CuoqUw8WhgsBYbp96ut0pDgbeAlLBFIHZQrXpZT1x0KzoTrrEt1cM
x0e9EvLKvbzSLwcwZ0lKE+QnlVNqm1Popj077vwyjdQDMPibnF+OX2WvpLAWNGzK
NguY7TW33EBXWhnY9TlPOAtuvMUpJ6/czjLP2VS+TMwMAvOw2jrUaYUNokIAWqUU
BsaUWNv3/zOfS89P60y1p18QaSv96NnXU5XPX2u8BxMKWHuUtMV8vVDKC05lsWS/
V7cGtJ3y12g4AFRBAsAyDpWOpexRGQut1PwJLhck3k2HfH6KvjW1GjAZmuo7tPgd
jU7FP/khVnZwgIDxdjxfufJtY+FW2SZScWXA6M9RfGhhPTDTZnTX5+/ZYLad6AM1
GhczcVMJBovS7PDitYxcDlm8GcZdKzlahUXGu6umAyxR5HZHuy/PMTov8W7761Qa
skoXhJwtuNV2HhBKuC4HMsF/kHCAooHEWjrbep9G/+CFe3SP2gY3SX8kIQyujeHJ
MvtTyy+uE4Samr7/FW24GyD58Ky019dKquF4rGz2ZEtgJGFFn2I4wK5bi6u7ddgU
fwC/cHqtRGaSpWk96pEQyMGST19ebD1sMseYsnrM6wOtiA7eTG0WZ4vCi6+EnDT9
10DfXJSBfSbdFjt5nOJutmUNdikoLvv+O7fr33x0MT9BSZgl5D6zkMBpXLiviYEi
hB2b0H1sN8iLG6y5WsV4o84G0enqg8gX8um89+48JB8joI8JtbGtVlLFVA2eJRz6
aPvFl5oJuA/JOl+74J/YAtvlF14Z7Vs9qLQTrDgNoRapnHsCz3jxtRgX3eM8bS0C
M3IL9qiaJgs8dmIBn50dmKX0LGBs82OE8WqpiCs2kS1ZsqzlxyTmVKacWCR1ulXu
cZzmiFIudkV/R5G7wfDKxTObQTnLZ4RFbMPc/SPuDhCmk/GvqFALu07ILTsnWq2+
m01bW7YTq1kz+GwpGcU90BWTe5TjsLs01eSo3Xn3h/zDcqPPri03dJ6hEQHMrg7N
u0y5m+uzKyj49LPaO29nksMpIodWpQE8+beJ5sKe220Nlpsow31Rywxl5P2uuOLl
ufIZ0bR7o4j1/rP97kBPdUhNNZQS1EYQnu7ia9k0aNBmAe09oTo+w1OviwERS24M
59Qyl0r/IppkxCGnQqR7GyPoJKWv8BRp4713gRAO6TcawCM1j4QvMcdkKFwFevIS
KyzrrGYMYSXhVQyjRgbVN0tDmsSGfok3HncZxuq5DMVCS23nVAJ5f3Y3Fc+KnBLJ
kiDNjKroN0tgh4HD78pF0e7UfrA+OVR45AdoN+0QuTll+aELfQ1JGOr9gVrKDqrR
YP6VP9DCGoFUAwNr5C6lLFHhsotc7hFf8CgqBMzbqnRwi6yThKVY8gkKQmbRxaXb
KWpoAW7tprhJ2W2428/Ke1fVh36By5uUBL3jw7wj2JsOVoFLq2Oxlc63d5hAlfPO
aK9cp+FCx5rikzj/lWPdZIdEj+ndtJmJeWeliT52qVoR377mIoXg5JoI+X68WysB
j+2+IlO6Zf6wL6C6nG/oJCqioOOP1XfgWfoej8HUIIl2pOXBtQazd08/Edj6pUkA
I62PPEs/HP/ycX1aaM3CWG1lDggKZOgVF71pCjhVAGEXvvvQul1j2/lUG8+TgYUb
or7ztSdQqz+IfTNEFVCXy4QN0w9lFQCuOU5/oVlt/VzCW/zNEiPK6TDO4GHuTbar
a5Ri1BMEOkdK/X7XHUvtFMt1rrctWMzXof8Bhzs4+FbvJ+omLaSKfeYT5XH0hl1U
l6sNutltQwhyIcefFknAeFgKCJdS0s8hbZCPHXO/8gd6Xqd9BUGtT+IAgONVKncm
xYCXsDGta7xr8WjsVofFP+QKtpEJnVBHW0Dc+w0hUT+t9+wO9yUzLmFtZ16ryRpE
723Za4ytlH3aRNN+7ztE7UwKkx6DbFM0ADIwhU1LcNvsaN0K8ofAxSxZACUkFKrH
6V2LaTIWxJH6ewkPFsGPnoz5AM3EyrTv0VIcwh2PmdTHHt7aa4X9PYn+yFli1t5L
FXXddyQVRp+16GTnBIJbxtCQpyNi46HGyS/jU8feaOtBAVtbZRS4DfmWwWsQ4dYR
6vnAqju/YxK/8N++1/V62xLhk7kDYrEyzlztiHKvwt5aGctrKkaL+ramjNR+G1hn
2ngdYzp0/c/8xbSaBwsaKX6S2411KMbW+Zel9olOU2pVmCi0cMReRNngHUXewNgp
Gd9zIlsKuboRt0jK9zmmtd7XHrNiNRUsx2t9P559BP4MbseO0JTDZ9OC3IMVN8pJ
GCZMeCMTjeOhzmC74TOUB+JeJ5geOLjLNujrQEkfIh6SBIQBQ61NxAAWpCKomGOU
lE6DAsNmIQEnfuFBCOoiyszXDBOiOcb/8BIZsbmDX3mj2/Fe5PHeuz+JQ7Bhrilw
mmij7i3Fyq6HvA4CI4kqyL55Kx/AdwzARVlxTQaH7xJlVX2jUcFoKU2lo0FVbPCM
DtmmNrV87vQ4WTnIS4mGp1o7U9j7UApuDOxQ5Yez1prVydqr8omPehCawkKobqZQ
WtNp39utiYvOvoKOr04KtnlZy+F2n3JHmiZQasUlK887tuc+YPp2eXLXhldh1C3g
H7csMFjsIqkR/fRZior9rR5AA016dO7otjRpObJNygxMKvuaNkqluscE3zjzJnoC
yGW5Do1hRxT+IQTCf1Jl4tpgug84SNC+3YxT36Ixbbs5iZJ0Xe8HWsNoeB2oQQpg
j8xpxcZiDoKM+rTl9xfnWE8GgvpkIipX6Aqnna7FXqDndXMXn7jzvxEYpd5BDrng
Fi+7LpYDPt2OZY/snJ/LFquUDeTUECWXVHxCP560hbVZES0kglTNblrRhEDQVzDR
+yK2ISQYCgP9vcRuLbx/jRSSwGPjKx2kjZ9CTlezSx1MLTWRzY9z9CxhjNlXLswY
CnLF6avUkayqNORvNG0XgLdhJn/hKPSF6f+d1DndPKEuRcXpnaTrr3EAo1wHgCZH
JImWce6vbKta6gD69ngZaeRAfiOAX4aIxsC8CtiiEyrmGIbVEEHXvlpHwFbwamMe
QWwx9muaB0+i0hy4xd4FgsGpW5tvZR5jR/fct6sFFtFcDIaHH/pkwBSjPpaxGMt+
Au0dZzmA7say6VLEC4tJffBd8TXU672EseIzO+ovD2U98QuhZNnHPL5K0b35NSTg
BC6Bf4z2sHEUDtGDPmeWzogevch1Q90fn94Wvkml7zaXgvqC9PjaJuGzPrquZvNo
K3mhM0kUmvaud5RgaRjF/No8aZgNroZBLvEAURFvcIW2e8/FWwfr29dCjA3pI6Q9
hweOXmN9KxYAFoa6ZNqsaaQ6qQgAyHBh98z+XhRx4jhffF53icpXN3MgdRwJobV/
90ajS52WdRy3phtwVtKe8g==
`pragma protect end_protected
