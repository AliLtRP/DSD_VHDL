// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Fe3kURCTWxHPQsHAG7jdXexp2cM61HyJ2pkXyHf5hWKmvZPQMpDbu4lwmbomZTnaksGdcSEHnAa1
yfStXtc4DQo/rcy+rFMT8jwQhadpfhnd+MaqnJ0KjH+x2I3l0guTrERyXZd+zOXBwg4mA5BpJGwv
dQvIkpOzn7nVbzPn6J1hWC7L0hBEdmn+/Mkfp12dUJEvIPVZFyKiP69E+zJeFBBWrWbu1xqfMn9A
xVa4Z0So5ZhiVAQ61t24LXr5mZLGd8e0OyXt5pJpk+oZnWaZoRS9jKkxzDg9tHgDR35/QGB/C/AY
kDly7kH4t81uScjTvE/+Sv4ycLN2HvQ1SBA0Yg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
5mrKeAdzPTcj29r7uA+lwBzKeW8GeDVtTBIrmXp2h7Ap693VgGzJRBaMDeZO42XzJOMPC1O2pTsw
s3/OkB4f/Q/mVG7ZyXb6n55772mh6aRoZqoQkkLh/URFh1WQOSS37iiYWVS1PzKlQ9axBK5UItfw
MOaemn3XhP70PCMO7p5IkDk3jbLKR31drO396RyDFDSic9OaYkZQnVOTTU5Gkei3wURvnvgoykOw
dVgE+Qu8Yy67HPjrPw5GTBb5R0qsEM2wnEC39C2J5i+kveoCwK33v4OGBM84lwUIpKAwBB0U3/bp
E86poBMVTW89qDTGYTqMvTNVFwRUizfVVJYqziNpQHQgfokU2m8s2IgjC+fBj07Imf6jB8EjWkmf
j1rTCrSV9Y0zkO9n0Mbug0r/g7GpXY2yS0ADkEJKkXIEeM4bVNquMVEr/rZ9APSzqSlbKR3UMe64
4kV1QZeAWZE3W9zgoqnaDviiQRFJqs4kzwNUyATaZY2NC2ZbXrOFxEvJnWltIQCkTku9CzklJzqB
jxra8e/4KHZe855LhIrmpIDul1dks0qjvmjz9fNjaroVf/M0KtYaaVbJAG6k6z3syOmznVSwIYr8
NNH6okzB/cnOrEPVN6N9CFG8U6xGqjESXLn/TymdNXr+/qXaSvijPquWGg22LAmvczMC6Wxj/Lkm
NISsYvqVZDnazNKLfsqEJAz8GPH8aN3/R1+bKnEqnODj2oNghRYZKg+fb66jT2y6OS8lcxwlJ6Ef
YnPwNJ9O8U1KLlBwsLtjnyNOMGmrryhlKl763h/B24lzudmx96DPaJ1/9XIhUDFG5XhiBnPZuIBj
HIvCrvQeytjiBTVh1bY+gsOhttL0eVBEwTRut19JYm3rpWQKiGH6TIfyu53aH0x1ub646zkupQaL
68+gkcICWFYncUpkGVgxa4lfAFXM2DWgR3wLlVXMTR0Oldfut+oY7DVueydYCOwG6q9gXArn1j5g
AKOq9XjudDcVtsDvXHCmoDFCSu68g+/MAd6NsfgXIRykzkPwZt8PKBBHhzu5vMlXT6SeR9c/e/U7
jOoff5a92o3xzdctg/OkoXhfmitOuoHZkHb5OnDhxGyRrQLLDuBbY5EHpWyJzI6PhmKNcsWhaIzJ
Gv0rD4Pkezn2S9oXsERSAW/TZtLf8jAJ+ZjYTl64yncuLAjG+f8HMJpEdRSiqwdMzjenBS8k0dsJ
bDa9CtnKXQ8aERrDo7MtnpHA588EvmSgYA5AuZCQ//y6E9kT+TTdUzfS9LHXx1uwC4h9UVqEf/n4
jdGQ6sJtVMMaYynyX0nkeMKOgoHvCEx1n7nexfx98EiotNJKam6i6zzO2fxw5+P6oLZfBUJKPcFv
urAN4ydCd19JQrjRaxHwGnDXqcbU7fXqZ/IbSA/GphECXVyWcUJuwiJe1EJMiJbi8LNyK4rDrmnM
dQCwPZOM+phoXmD2PZOTq8ythbJpdGAhiRGGqbzNGZBqpkIenzKijdvI5XQkUCq8Ux9SGaJbcwyd
DO3xV8QFFHX4NGJuzCAsDQZKD7V7Xo+LAeVDimDC1byziqqjFfTm0dFRYJkNAYevTelu1Qfq0g5E
F/zLhL2ytdh1NKr266ibAz4SqLwzbewbunDYTwSi9CUtulfR8W/pWxXKdHTsMGXXa9g9O8a0gBTr
eEPMt/+t7sXep8LzydrrDV8VZNaAiOxs23CeIdNiJQciq+VyzWnyPqBljt8sxuiqH2THFnzrQzYv
P34/X0R8GgktESa2GRJ7k8AN3efeTzrLs2exWiDrQVSBR6Tbc59aFH6bVKv8dyqjulyEbKf0iodz
/WQ4qhCaBQTalaBEfe4T+QSCAs/C8IQoPql0nPf8H32ijF94XjXP3WwLacvNfl5q5M0AiCKKuVQD
MMlpcvvXv9jtfDq343IvEhZ1B9+QDi7f9knpSboYxU/bBJTDtNu37EYv0NJPnzn7qd4O5HcNv6eu
j9nZ9+B7f7hLpjCp+6IJtiRXw+s6P4AmClINEllcK+mfJX4cwFVYLiEsXG+0QLZ5E6ZaahGBsW+S
lV+ncuQ8CtJbts0liYQmoCn4P/lnd3ndNmBYDiXBggr5hxw/vfWorgBXEczEhbxat5At79VfzCu+
RWPGgTwOK3RdXLH6ESNBTxsgkDw3FDXP9E7hUYNBKLkY54gslhy4IDi6VAHlxnswrfXjC2saYR/9
fJfHhmgD2o6/JFEJy3mPvTQsXABqdxX/mI2rgoynRtr5aDswtjAc9oX5fsKk1LwrM6M898ojXKY7
9wHMqARctkuSXUPVFWwW51lk+Nosdw6ze3SDe4GFKwdnMBQKBPYUQb+pM6p8l7cr3hjO8o44BuUH
VRzLUaZGH4S8cHKSi6iMnpkT2rkLcs5CJ0ko1Rx8Hk5Zc/zdYyBRvBdSlt7M84cmB+VLSG2fCVex
J1cDimZFFImk+j9gd5lzPpo4uJsGW+GfHjzDyNxJAgc9SpaJm1L5inxp9KYipcZAyIeKWZ4bmD8J
R3zC3qHUWXyT8xU5UoGY9N9yvdi58zF3Oz558QqijAAPpzWCWXaGuFEZveiQ77XMEqI/ZHOx0utB
BCtPnfqHSVFB44AeiKcAsGKb9S7Cjo5zedTXJkOK6ZbrQYtUU7vhO47loEGPcdmyrHA28gDGEuju
X5xGRerUr9+JJPPOKo+eg1rAw/Npjddd0rgXTUfHP+BPjsMkhofa0VJzRH5i03rJaYLpARMj2krr
l0JTmQMh3AO7VAKcv1w9eIK5DBm7NTWtuhYIBzFL+a3mS8bFLVCGPl+/I3wdYvHGG66yeTRalY4/
W8E9Vz0xu0OSWBWXKvE2rgxhcaRYlWssWso0USg/ah4fLzN99dJLni5e/6LZKj42pfucq5dZzKcc
ZYWze/sNhVrI8TTQ5S4pw6xsM5njzIrJ1NCndfU8aLtqfh2i9Msrj3nl0MgTDAndpuYz6YHlbRwZ
ZgirwCMo2Fn14FIuPIZKnuk+gupSJe1rLkI3oTEfXZgmP0ZxdxeX8bMHHSr3aH72sqLaXwWvLbYY
o4l4zBxvaBAOg26WK7+ztAhvP10VYBJEG47EasS41NKkfOBkyznBmRPEctqXyO9KRt3zG3TwzbOt
OfBKgfYLJBJU6Ae1lqibe1Bj8Mpht4pMc6jzhwmqQqnO6i4bdayaqpthHJDZ2KzxAJtRE8x9BBHm
cCDmJgJCM7L0ohxkhhL3AmV+VJHKd/LM9DqOj+YEar42JajVY3c9RuuSkGa7S68p1o59IxHABHzk
inrHcMeY2oPD3zGf+OIwLcDp5x67WpwG6k854Nu7EtWTJwEl3S01V9lE2bD81G12o/Qj8zBw7eG4
cdaKcZtKQrkyVO2JIqsz7sVit65+6/HuD5pKKabWEi7kwH7lPn8SulN05JWUB+hCjZXss4nz7gZJ
J7U5ezXufeRbIMmsqq0G2W4AfMO55Gx1IuaZ/K7z96uVDniwpUNuw81L9m7nPOEO3/MXZLUBaPjG
cIUe6cR7gPk8pFpsq2KWNBAynbPyigUIx9aiOKjnym793Tzj1xIk7Pf8ZESM1qwOv3/s1OCD9xXD
mCsdWQJLtZRW5EvFvzCPDSVSSFlVZ1fKudQqxxhMymweQHaceph/7W8jSivDW0XP0aB/oECIT+1n
+rzgv34h6ahhtgbQyVm7dDpif3c6WtuO3/zEklladrYf8H2aYIZtTev1N82CbWwr7qNjshI49UJT
TPxHdwbpDjNEWLzquu5VAqrsBCUb6KB+86QY6RE1DDEdJpgD39EL+EwgDqxui57bsImb8qdsttDM
B4oDknHGCR/Few5jm04ZJrfBnNBDWsLJlpGk6W0T3ufIpNHcVXoRZpe41OoK7kP9PGJEGhL1E09r
SVu9rDl78IGjsaSjUO0qUvfOKtiKtfR9evVn11EO/CamnZaVTG7HzITvYTLNYFfWD65uDi93Frg1
8HnjBPK6L6RA67ucqVEb9iY9ugkKc6f613qFuHZA6dyG/7Giyrg8QJjWI0aDAjvep4KFW0seyGkH
R9gYn8PHLbvY7+n1M9zODddL/Qprw400rCy8ZiDqPvBoARP8H80pr7oCTfNiPk6Hez14dGsvzHCj
LilqlN5anUpMw1cHVgDS98qA8XSLnffRTBW9dLQywDffYZi7XlYMhANoFx3aX8U/T6NnEEQPYeRW
HTZtVlAyrdXF14CjXhrzm5Jv0+6d/lgJSujTo86/HC2Q1Fn2BIBiTNIkEPnFfKaa8MaiTzinQkov
/FBs+Hted2L5mX8nlXST9eJCmSfGgvVNpLuWm2EXWbVvKGJBl/ki6b/SfJgK8hYR4cxiRclLdhWe
C3w4I33ocYqwUyQ/PRYfMIWMJ/QF6q6yCPK98MmAEeamYDFHUS4yG9NQbbgHgchtZvVVkgN6UgLe
mZowRUD5eHfFjzEGOXJusBkZmIRcFo39uF1zsb4WRWEW2QdkFdviV5wU5fs6KsCQ6ghVujhM+h+i
xYiAjycSGGDmWy3yCfUrPTgNMX9k5Qvw3PDbexPxeGt9XZVEx9G52EkHY2+yTjOBEJD59h1r4Dy0
2WQHPUQReJesk+f2N7x57rHPu9YcP4z27o4E7TjMe9JAZSLzHZBDWAFcz2gSr4P/9dIcNNLoHRzO
llAPedBc8mhrmxCOMHRWZg8IjyFq/UNzAtPyd/FQsNReNMLx9ohOtwj0gH2Qcs1jcRAN1euSaYFp
jLnymuTAmANu7a71kkH9+KkCAE9bGzDA66GhHY+4l3VfrubvASklrJCeTC26ELpCO7aFGlA6z4lq
AbrEEyZ2t0iAA3YaCqzJTxoaPQSY836y/D6EcahqZ7zp20S19YiUvcAvJqmkeKr7I4ra9CC/wpvH
PdS2AKnSjOMn2Ms/N0rjQJ3AX9N/z4h9aqrQIFlEGTyBwmdqo+tAc0zxTCLbq/qqcjLuFBgJYOCo
YsiQ3T69+GYo6gyM+qSsoROSWRhVbQS954iuUdAJtWAOaQkRN60zFd73vJpj3/6Om0tvWruJTHxf
l1gWC8FzoATnB7soW/Lts9jb262HEVeoMQYcx5gesdOpXMpk4E2GnJj6t4ut209vr2f6lOn/JInA
PWy3Kx3TwFIEwaXFbimlVSOdDekAY5wXKexztxquolfRLEPxvEl04TeztgLZ4KRWcppo62y5xU5C
y2P1zOGTvUPMuhjAXL57X1zAP+P5jnaaQpdTtJA9P/Dxgx5O8qRCCQgshCOkuKnOfDlmoclpNIiJ
MCiPj0BcUT//rW21Xt5klncfK87HN8KpduZSfqWWQ8Krq8S61uyXvY21Iqq8nUrPK7t9b0kzYTUN
/msoZ4lPYBZMAC3/kWLNzt7qycn+be2bv2sj5wLqrOvXdZ2CqEo0QDdISUY7IOU4qVXUK/RMobZS
YbtMNS6SO/K+i/pHs5H7cRQ0cMp62GmPS2fKZiDu5vWKkvFd/FSwzn7w+g9cf32CZb2kyASsTNtk
4BW/f6kzMIgYRISzTzymSpAWo6nnVi4wjp4OZ16rnZIYWlFQYQ0vxS33I3vZllMu+IB2v+bxqVK1
VVBXSAbO1a51R2aDUeJLm+ygYqwHXyp6jn61ozvsrGanzi+MDaSF6VCOD8ipIwJQLLoII8rfb/A2
3wO6UvakerxogtQPjd5CRggXDflDxuFObiqKQtlqH3mQK3TmIt6EALAcnvQLNz+0f0tlRE21ij3K
VV+E49cFPG93IMk/SNFTD9jr6rS5EZYdjgn2soU9Ft/if4H0F55Lp/G6Ya4owqEDI0GMiVv1w82/
k9vr4w1tKSp09KHa7r2Ji6f4qKX98JISMyQ9zLlAvkQvCz/l/RhwcP6WP4MlUVemdh/9SlqOQyrN
I432/puHdCzJvz93A4Ot0+Gk7B/JbL40WsbycyDArtHPZC3a/py4M1iHAUFmG/954wAe61gTmEKU
mL0ZGyYQutqqpRsetLJUyMdCl0EeaK6I7Wjs8p24ifBaw6OMlBsWlu4iHbKMBXfDlTLnhfYdI3az
FYuItExhVwvRlWfCO7Pwl0aq0R7f/yz6ToXjx3NRJE3kAW7DKA63ncikmgQe4JvXot7rOr+5gU83
j71z9rGI7L0ySD0GmLVwKLFL4eVsddk/GeDsbAyjDTTQPsCV7n8990c343/mUuOt6u+5C5Z6SEn3
gpjBsOppTZ7A2V6qae8wDMAqoj1HmYjRTNJqXVIuo7lw0+09kNDEWfdydO5wRCksclX2kaAJiT2x
S8i0ZyAXtrx+RO3UVleBs1VhTlDMdJqYao1cVIUG5gGVcYnTAoewUuJT9yMq7XQ5SWX40xOGQwNZ
79l2dcjcSnREgptAO6XzUDi7pG54W232ElMI5HlJUu2EAoLNJhl01pR+HQhrT6eoWoiV4RJlLN2n
CWulPoPfzIUTI07hbjUg+Uo0K3gvDA0FcMikTzl++ERCp2Ad9cWClYWD3qUsowYngB/87C3JCoVq
sRUlE9RgNNfkDNokogFLShG3W7TleUTkN7ib8rXYfSFHU+DFM6fieqKRA5Bp23kgLFv4LRTBGUE6
lsCZWBzu7+jC5lEDsYAnN8L6W/RThIET6NuImA20go55/3/1aeYX9h1dUVP2k9x1DfYMrFT2xAy5
yMbnNCsGkZ/c6XEP5DHMIwseGksnxXfSZRQZY0jtibyCfYwlDjv0KlLdMDpKBDvvbHpjIThQDkJ0
Q8ajhgmueNMxNrU9r9nLk3KP+gQzDKFul0XWlL2HkABM6isMTfT9QgVZPQ4oAD+EKHOGrZPmF3qv
zYyuCpPUOWq2HgPj7Hj1a7oH7SPjRNm6lD/SFer6EQo3I3EK8QsMG7yEDKcvC+LGgai3PcLGT2pN
6YGUr9Pi0YxLH74o3FAnhv9VCzLUd2a/AQ/mfLAUXWpBavrKS1waNrvdrPBzNKLrwZTH/bPLPODB
3j3eE1oBtqP2P1WkdP8MpHFllyW4VqQCK9v1XYtNm49as6eOFVVG/PMTtlCAQ6LLXzCpkaG+wGmn
rJU1xIwnDL1ZQwZ6qMO+BOFE74dOlWf32J3Xu99B693I1aQ6+QFO4VvV3bHdK7syOygUr/RVnoG4
cG6sqfBnQ2B1WSOJbfGJUltiU+AAFC8kyvOIpN9uDsihrPSYicOPeEdvdI0wuTD6q66m1jxNpdda
tqsZ5AqZzZwDLE4XDmagwICjwwG8RjxzCi8nEjoZTRlau+Mu63Qq8XI4MPHKZbC32//jFU4RamJi
igZGOpJxNvsdhOUDXu+km58A3p8f9brJjKco7BSWMRMb0Ph3/RSPsa7YSi7bXwqcZNc7XW2VVyBN
NSfQyUHZiaxrBIP9Y6xvIO00oZ6m2MA0BAd4zTLEx1lI4Ieg9TlEqOc3VDjRUI+YOQNGWCuioUnS
bWVsvMESpvAkccSn5FiZRvCkf7sqKtHI0MVXWWFhUBPQ2cAmI9i8LTtTzUpuWgNu+rmaGKTjVdov
KUs+nr0U//EqP+FWLyRrTMniLi/9abHICdObRy/l6qSMeg5e2rPGE37zuTBCrMZbrI4I0wf5SiGS
wvxMHbvLOOBJugpITsvN3M3i03jhEWL4zmZh9IjwwYjduJxjvdaAwrezy/hSG2Swlux4OzC2nrAU
9Aj/mRkA33kF1Xn4Dj+5t0Xrl0aSYNRxaMwy4xj/0CjSG8hlw0CsB8PgzQh+ZIXZfcNSqrBdcas3
Ev7FBo+8MniqWyjugKiaYar2hvTNg0UFOp5PX1pzqNDeV2DxfXQlZzjgLU4wHiFGAB8f3zD9ApLT
DRo5s4kptLQvpQ2vbfduoualz+fmDw7O2VKt7GcZF7PvddMVx8FY206nyk614NlYoJgBllUvJVsy
StR3hHF7k+yyZxUG+lpQEtsEpkLP2agrmT0emfrVrKsySZhuR7Uh33TQPSbbkJN0zX3+lw4jzR9r
HX9JZqD8N9O/mHAgg5hsZM8r+60E1F3Z94JNPys1yqSF+XLZZfUlbFvDJvQG1cS49tDfGjc7oZO+
2fCqicf4jsUnktayqbtTqKdC3uz5WyEi8PxVwbcR2spEh+WAVsx3pZ9Cf8ifExbDxUdIwtx9LhGa
l0IwaI1PFOdjOdYlJRYIOyKZnV45RWoVFp3b5U/QxZSLUzTis7+lZGskLYXRDTuj2QuiB14klOtl
HoK0LXLWq/D0dIIUSDyFDq01yo2VLHJhA8qJHgc6Qk/GFJA/4ASYy0uE+aiB+PPfdBgxE+4qg3s1
6x3fDD79/pir/AujWC9E5jazzxogI1gv5RBavGZnrxcMf/4/rEXCFBhn/lRozWJ8NpMMAo/WxPdh
ykDo0pQdyvNc6V8f0SArV5mhiJkRhkaYeHZahbPHrLtCYATtXoPkdkxJ6hlEbxj8Hf9KrrSZlsFI
tPxHqKLw4BpLgrThupjIl2dNcXua92kYTsaUrRrjPhu1WERqOp9zfZbfcXbH3cht7anH4NUcPm8v
QyAo1vmjt7bRC2zSkMOwkGRnGRdzCdF7MtghNqOyHKZs0K7MkXsLy8DLloKP5dF/N6VXfN9/OjEB
YVJzn3LGVPbqrTz845y6VHT8a8QDnwLjlXaC/jwZBJenETNTyMGrOkLRCYsCIptv6cd+e32GUurE
2QyuEScPI77I1W4eogJIGmGts34IWFjEbAAPJnVg1kRqXoOr62kLLopu4UVEgxFXa4e8WJuVXWt/
XrSh7Fn6vBVtf9Pw7TKUzjXRM+UHxVUOoSo82UJyV1DEjGiW6esauxj1y8wzqsKE9JXtaNrCV/t5
HfwThr/pvT68bxUOuz02qMrs5rM3X2nYrJXH81JBd8l1iKRxJss28Uc1uxNZDLpJ8Cqv1+XYXVtp
Khu9ND/OpBvtCyc0ltqgcNRBe5OWLRjK3j2xMCCdnzobGnpKfkiE+iMURZ1Qzmd8CknzYnJm1+aX
SFl7Idg6B4DdjAMMgo6hewaJkqr+tY4XxP5GAPmUwDNpz5AzabCgFiFjcqo90KWotXKN9/L8U/R/
2gDo5MeCIje0Hn2G1mj00i0AGARJ3xMTkJgMZckP2Yj72RKmka49Yx5/JdNAotzQUVb1y1Tt3oSt
Hvni/gRGPfgFf0bTKwf4IpHWQCrsFRcBQPmn/1GIoR+CHzM3hpduBKKziL6wIGkZxZQBphGKD0WT
1+GkJGkzjW4NsP3A4U124DHg12UToXEEeNqhfIDXbEBR+ZRcLOeoWby6B8iEd56ZVpZ83zc7bgNb
TTPAaO0Wiog5ExvYw+NtIe2iyRZUvDRdSFhS9bb/bfJSvKZ/o6zdXKDCrJKtdqWZR5yDtQ2PTJBG
6wmkizLY1ipjz8EGgufp97Zx4Ir+V75wIpD3/l/lfPTa3zljcBqV2veaV3/9RAqtQPg33W2s3qkb
IWRwjofrJNq8JJGYE69ECFv+yoK8rNdRMFuGoaf1jqkLAtt73mFBFWXfwPWiZkzC7ZS3oqsIDloU
qaWFJfmSxIbQEku16q92VXQtLPjvRVSGwx/R/QLbJhK/+/iOAfzNUs93FUBKZIK97+F822kf/13b
S421xoIknbj2jkBJmRxEGkqilvBMHm6LnHHG/hxpftwaOR6GC7QCHjye+981afxahFDCGRUQYBzZ
myiYJBDEkuBUG6Vvq8yMK3E2v+gJOxiJrwGqqiBcpj/Iv6aYMZP4hBeSa9lPM52qYoZmSqWAWrEx
vhu5O0OdMKNZ3porVi3TxVKvuLcUhfd8g60+AY/QpphHyJ1JOTaph2rxVbOPBt076q4yps6sszQk
bys93X86oXg7u/DAV8sVv9MeSLmy7wtxm791vprF76sDMdtxiTFr4bBlaIY/2vKgNqHUTezD5dB7
GZ4udFi+D4xaywWHoXuf53mfcdt2o6DyQNdsWtLy2dCQ5kg+DJSSZYl0dcuPSAix2aoYqdyc6AiJ
jVrRsJqarBNAfDi0r1jsoPOasYijZ3uUEDQ3Z+91XdXUl08LvBTThbHGwS3z5kNfufRiBl7H8C6Q
0pD3r9xuFXU9hE9FF5Au6Dx8aEiIokS816bZu5hgAxjKNUfiovPK2LshlCmq1EdjetzD2ObxvWR/
/hz76+E9Dm6KOMcLRISHNq6HRWhDYrw8Jm8ppkIV6vgHV5d8YfpS0TIC/C1jwvPvcfwqFUjMQ/Nk
Eu98qAUu4zu4/ipCwdVEOBGrbZEGlFxLYotvaBN4ozD4SvSPMwNmNRODp0Kdsu6TSICzWwu0ACKu
XLFcPfuscsJRy+XXrs06+vWmWSB1qTBWg/2DY4JMuW/OYToj3bZ3yuMJ1/UI6Vmwq0Jq1Nq4stWg
Tiqw5T9p2yQcKt6BBnEdmluDMwpmXN7WPBTLKG0dMK8B3Bac00vEvnLKQTNfunpegYR4umDOPKnB
UCKyrwzVRgiWWckO1E0jDuldo8/ZvqvVgT9gvrQT76192qdZXbF42OIcutvjVtPblJ94srBrBbcJ
HtANgMwxQwLZ3rnkFkqWcMqVhVsZL+j5DhLPFyXliuWcb09JubEdUjiPDLegRhvhalzwDB63+cdg
sEdqM9DXizxIDbP+P0GrsjRBgOPUG6Yj+73tvOE/qMMA7jRGvf8JUh6b45h/D5sMuZrLjlP8Ifwm
/1ZjDjnNuSLGAb/4wMHJ8VlTNMItolq67sw6++InyglySV2gBWsD5ldecn5B4dPFFf4Mft17NRcY
PiCujlwvEonISRvpGjZxj9HCojl7dWGPClY22kFSelbQesQK6aNub0CsqPaQ+GI1dPiMGYIPsJqC
EvaSRnH3oWmfAz6pox0mjeF09OCDzY++ndkt4ztRVeFofhSjXbkc0xHbWmZS0vBEZNUWgso4Ppq4
7dKuxj7CzThGK1ftgqF9/7M/6cosFINy8jn2+g2zGXZkkI445XkHeYTtG0e0nA8wCZwp99BhZ5sa
RHR6Y8YWoghcQPiXeDL4E7GicoYqwIvehJk5pNkEMxgy/u3XonwhvrPc8eiCMQ2GW/KcdhkYaEtP
58h9u+O9yqEAfvqlNweOToSugyb7YanLEQyHw8kjnL07f4GKG729IHR0XYFxqGcwrlOjM9ffHqgi
f7MVdEoVC9e/vH+s+18TFezwrfbK5AzV+QH0u2Tz16KxKPBXaMPCHHbGGiiOip3EbUf1hXrnjGOn
JX8eolFaCPwJgkYR1oUpcI14ntvoH6abefG5RKuLHp2uh7x6jXMnEfHy1Tx6GH5inEnsVDiaIm4F
F2l+TCBxXzsUnNrA3oDm1ai88+MvN4rwUx1v+YwgsrRVmOjHxD87ZRPdOnu3Ac4le0E2kR0ofaSF
5qtXOqZrSG0Zi1f35shkzts6DSUHz0R4bTR9dPLGXHpIvThGf8rsVCu3sgMngV8/HWaip/MSmZsZ
XRZUI32oqIPewJNbKhvbfpdjOiOIIujuv7YtaNFxWZxMwL7dEBeSB2qkRL4QgsgNKd2CBGbe5PPo
9kspywrjdL+4pbluYAecKrjlxD+ortxlxskwtlD4ZQKaJ8bb5HS7kxFD9u+m3Bmps6Ht5Uh+Vfgj
FLszeMsOYFfhVaitXuPSXwNK4XqC5XF5oJYuEGgsUVyZQykxF4TQN5JheeCUgg20TezaAdFMkfpR
kQeR/Ap1kfyy+5X7wSId8Ka7hCD+DjtHLJ0S5BsKmNg5Y7bHXfhfsJy67Lx1TZ7AE1/L1+4vv+++
fekJrE/HH+Jdmag1Vm2VP4Lg0OdyfBgnGljW7bWNICF+5hTzDmcgH5i/jULLXEF7EffPvYtBzeb2
L8AbdEjxqaGCyM1xoRV4XXagC6G69wbLCBeCnSsyuAK1lox4yx5KqE/QJpTJ6ltFmQNA+eIip7E+
08qDCawyU8t6BvGX3pMs3fz42sOnSxO6LZqJN9AjMmhb3L+3xGSB0aI4OxtHjenQK6AtbqRFSFm5
j9+z4uV0/jUSsqyOg8P6KZck/eFmNw/fzGjdJsUq2/D+8HVdeBoLIgI181y7Pg6IPxWEpc17N9my
nuHiaCf8ccd/KG7Uu0kpZiD1GaibRERjuhrnmgkP6WRmFtkRo1VgXIBxInEJDcfQCfqp9NUcre+I
mrl4GKwl8BW/Ah8cIHF547boqnz1HW+x/qOlknI9oKLxHQ8zaKLt5I2A4+iFurIqYdq4I7G4+8sF
8wulrFkkFf+BoPfHpmX095L4K/Ea46Bgnyb+dWWtNEv/V/if9ePXq67t+WSGj/YIv3c5iafYCA7D
LOYlK10Giq9pfibfscNu50MmS0e5crXvfgSbnsTeDdJQfV92SwzeXrk2hCIob2SHaY1fwYsoiOkj
Sf7w6fbcW5wUFgzCdGYLf+x3bj0P5znuJ5jpeML/YOdB7sp4EiKibSPstng3lqQvWyoJjlb2Td/7
ypKuj0xl8nXfW7cKXJJSuJhGoOWo97OFhplwZ47DuwDP75kgeB0v8O8l7BoBCazamiPkATKbwhfw
CMurNS32P4xwBPoR/Rw5vKdf+RBtIADr2Nm89piKQFiDRVIov1rqQpCWrPNRvIBlv25U8MhOOF3a
N2Li9z7DsAVtO/mt6BFEl8wwYDWmMFCKJ1mLvyP1wPQZ5ziPUSTbZivpyrZGYYmG0ppkshbW50aR
Z7DCIzLU7+Aq6QUseBaqpyeVlRo3QZW1yQorLWZds17DNqFl4ggGDup7DUPT4WEZWWskQlLz4zsv
A04ZQlCtxx5sK5YL+2Ff7skR/zsOwHbEd2bwtCZxzqozvjZQIy2gx5OrxvEemVOb1zv8HNUoPSMF
dkolBPuRP1Vgayb+5Br7B24quWIhvqHvSMjubVXA5m+nDxeWVJqAHH8Qyev+RvNDulgq3tMGMRI6
ehBCk4o5+qAlWdTKh2Xl7xFqTH1GPYCCeR/CnvnuC+2+bYd83dTbGPB7I/THgipp+Ixwdk3bHgkq
JdJSiq53l0y9gb+dmFSr7CQofyuN9LyY8XTnH3+ypWZgnYY+U3U0fVPnZl3RRAZjsjuvI7eJOt9M
5YXeGe79K+RWR3P2N1/H98VjeBZGDHefH2Ne9PTHFzceN3SoKl5dBfuhaGvYYBRDR4ynMQd46NKv
90DdxfAt5I4szD8QPvD3sIxp0f0JAIj5K+3lT7es5iFz1wJmeyd35l6QbHdaxBL9jcGqkgTC3Zta
WRv27x63uNCS9WobE+tiNUHerLiM619Ng8jC1pHi7SaHiaRS5Fq5xmBnlzVKxvMY3N9qftM5hm+n
JP1mYC6DO+N0ffnpj8dgRzYouner3QMKiU4w3ezSLV5BxRSi1oyKcO3j1yM/MVUt1mM6yWVdcGte
afM6UWpd2qtpd8/6Es0E37Wxg1K+YELnTM6hTHL4i338hrRpcZLHJEtU0zhF75ijZGh50x59onKC
J3ze0jK9nQRuD55v++Zh8MPIrx5aDA4RAbD0fRETIeTUToe0xWK2AyZcS1M5fOYCjKhTZmKCWAhp
bwiqhzUxDMtOyDaOVPrhAJprY4EOrgw2/l/k7CEAldWMc7gloEGuv+sjk13Ws4mdIs7bCzLejt1B
uBXrHplHKNgXE0evrbmfHFVxp1i+GX+480BLJZiziRumeUCup3tt5Es/6Y5QpBXlG3wIs6V0OyAE
iEBEjVQrI/2NuwKTgLJH9VFIpVK2pemKr/o1zEB82pPiETZ4Z7L0uRAivjcfLu8rA97nNCn8Hd1q
Ec0/uBX5pYOY7hO0R45g+9DNaN1EQ4KjtHAtYG3/OfioZ8JpznsDTy9PobkXaIDOFjDebj7wnr5G
p03zcemGzxHsVLZXmV8Rmmwc7MRgK6ZD5BfPRohBLbrTBelDWKb4cUqGxpqoHknahJaTKgvHR/hP
Qr9myQDhPvycJE7wG/LBt+e/JxQRmmRm+iVoTVacnWu7INp204LWbVpWfcYgCg+l0EMsQaDd7zdQ
VG5Jm1iECmRgGK+NOZ1Rn2QvcZkIGC7GhD7RAre16N6rwWsOpMLjK87yBSI1hftUnag+zI5peTP6
xVITmDqzGoJB5MZBF27s/isO81Nq6Go4TJKOswzXaAmELINEmWCEU32uAf7b0tiZ6r8xGT1Xdg6b
cSCK/LcgUjMV5eEs4a2PDw2wIZH6LkFSC3FfJPrHsc8bPfUBL1Qh6bs/1K02m7geY2xWc3DgMqdA
t+BuuRcpQrcJYC/jJVXGsloOHzYY40ZGD35vxfDIam7CGH5LSeqNePKqZxXQ41g5ZCgCQx0MVeb4
KSTqQOlZ0PvftjVZ9KzDHOnfkxaZP30Fcx9kmcsMyqmxGoPaxlIIsDRxg7Pss/iVfkFjKYyTt5+q
IZ37n6tGG3qL6nPOtmMc1RyIa7jSSd3eNGKmJb2/t8+Xm+UlDNMN5DmTmp60BOv3UZrIKtadgHrW
syeHoYxnVkt+1SciGdkIGTfDhRBbMIJlt20rAKy/v4TgJd84Fv31bw8xm7vU3ULbA8VC/N6uhj7x
t/aGJ1JwZhWYWPWVpoYeYUpZILPy7VwjK4Ant2gKLm8J0lHNhNv+FEX/lG1oOFoycoQ74vXz0cY3
Lzs+9azgdM8BIge2grRmsBjdB+m5PJrpv+kFMPAWH1KYlzLlZKNneg5NYRyZpfqLzpdKQUFwG/R8
aNiIEyYwkY3yqo9fWJ/+YfGNuK1Nu+T4G9HQxlXQtFnX0CixDdh0nX0hVR/PIDmSdeQrwbvRYUWA
7dyJJrmJ8P/StldoaOEsK03zLyl/so4HzJ8cuHHIBI5gDYPl83GHjRVb1+NwGyQH6JqutNizEL5k
egZjsQlsrGxQAnaYYm0I/WS1zlquxVqi0ZLIxS7kyXr33XFvQQ55uZ/8uiqGPjXfng++9Ur4eKfD
E5AMhxA9Clyry446T4Q0zsCThBrM9S0y/TZaqfx7gOgBZDtfjKl9PYiRxMCLuaYXzBpT2p6dudpg
YmxF0ZadaLBzzwxDsydsnI98mfHKBp743vytlaiEegsI8e+pGeszXOCLlKjLRObE96ONjp3VQ7Jp
7rldUG0WjorqHb3ckDsSJ0qs4ot3GDsOIBUJZ5C/IzYtBVj8UiSBRBnXluhv44/afy67fgWdlFb7
wjL4rWcDebwA+3O5KpKuQo7stFUhyyTPw0rVSieNiVNh1fcxyfMDfoz+tJIAQZkLjYoWDHQRZBFR
s2e0z8SyWRc73s3JxXHTAhakE78OPA7F5I7VKTEdMtlpWGdL7xwS+0r4bB35ZeaU3USjze37mEXW
liSiBFgXxB4G1QmrtGbD1I24Cgt/Gz0oAi8j3yn8RpyTKgDwAAbibWLl6JhMZiP2xRrFgLnN6Mbn
nBe8YIOlHXJ+E3hNlnn2UjoHlkN0GNHCIohXR5L+q7ckt8WoCUnUy419yv0Bm5Ox+/huNqJ4vaMM
F85r8x+fQ0wNzyVeUG6Xqn6JBGlb9szCRBibtqrAQENg9RrcHnDtcCEW4PnPfwF2O78K5p9xhkyS
ll9mQY5LZG0axiTRMVnMz+WxLpjN3NLrmyMhcbGGoCX8aPQGB0MQz5csJ9FPDtcL7oNt7XCDF/aH
DiujT6fXWm780WjsBR8UWxPlkJ3N1rwhDY3nGri/bZqdctkcPPHfm0vZ2uP+S3BV5iPKSn2RHAHf
oINGr9aKpszkeJc6arLnYeT8d2SIGfdHB8gRvMjXpaRd1jh8lJlVo2bE1AiPVhotZ3IYihAIRtG3
6BTlKgccpo7cBc0xPUYNDqSvLhUvKiPHmrMii/IBOLu5cu5X50fDqyLIbZ42WpzYCzvBFFZ4/CN0
3yFKg3tOp2zeNPw1HfWin3J5tGn0fLqr12rsCvBN3TQ7GE+cvH1XhFMrGT4izNwT8VOzpDCtkvb+
dsk9dUHUlRGof+0r7bbZ++u3q/oKc1rZP9B5fjpvjky7Eda5G8bmsjnFhrXDhrzl3JEHi1Y3JIXp
/iqrpoXThaTsK8sb76EcVknPOstviZbo6GrIPyid5Lge7d6x4/WD070MJPwHZEsENvzITTwtZTB/
6hA4BFduIvOzgOBgeg9ywuXfjp21iMd26eiaaFxNPqekvPLKTBkNY/gZiB7M6q1uOvjsTyJWXNh6
4knngBn7uu/yVFQ21d9kVdk0F3BWroDVPI3BYT39VpvnrxYH6UB7goQXx4/IFvoAJvHAMxARVD8a
Se4y+wjDYSeaf5LVL7yRDQlbjDT6AdM4eSq4sBXy4CyTOvT91ufcHQ4VlTJLc4r3Olp8teIJjsyr
5LOcjqM1U0Qv7pWw/wJCYnMlxvRZtEGvlFYQY+gM8k/qn2yMmxQlkhmjzvlQyqgJj+qxM3sgTLd0
h+IsdehbbSDW5jxPWouVtQaf/F/zK7ViYPwZpFIgCAgylc7wTJ4UfofIo0ujBAkMxu+LF53yGk4W
TkA5aU3VQRxB/OIN8rCo+psIeEqCKClcBi8oeYj42VO6pDk+yvwcEpGMG/CykPf7YEPj6rbdpghe
BhOUs2pM4d10a4bjhn6mxDCxvirHu7924tTNDfRTY6EiR0lvwJBmUYW7wdXJPo031F7zGmGhUTfk
SdR5dQ+om8gw42OuXBzzesPi1Hn0xByLToabRKLpSYkBpYIG691Qzq+KgLo3HvUS8eJvD7xbcLcF
xec/OlOcwZ/0ZgqEuYISIpZM7Un0cJ0HZNqvOU5zADCEy7mZeGBSb3kDijX8vVvZ0Xe+VA5GKV4P
i1T/vQJjYpgaCWYsp9qiewKwDDu8ScbNcYfp0VfkD9Ae6yC9WKXzcquKWHSomJ4b+GYbEgAzXC8N
SqwaBAKAJice93Ht4/5vj8Su/nv+aODWMk3RVWGvaeSlqsC+ACrOi4JngovFqDYFuuJ5jQEY9ZeY
Eqz5fKhg4fGNixHhHjrjgbYIUtlgWRS+faAtnOYhoUa9UOzfaqXpon9XSE35N0TwvNN7pgZ34t/3
PAYNWKjJd2HUb6c2GHgax3UwUKKqWgfg1gy3dwrNAGBc5LzrVjZhTT6ObJJr3oMpdK8BqRrqrr+M
9wirbYRGNd6hdsJ067drCsaG3Kj5kmk4Nj1bIucshrZC998CN24NK6ZeySfvXjTNeOyN4B5M/5QO
ymoQIpi2c1PMh3R8wuF4pY+2cF0wmVRyHLT+/JQDVmNePWAjnKz4b+9wYDkhmMFKYD9WofJBI2n+
2FdF4rG4VMqTKJ8uKoCQtZ2tFC2KYaOeK23BZtXlwnqILS4B6dmCW5HrLMtkOCSD76nLvz1QLmNO
AeWQ+ljwhvAPOE/YRwjNPIufIwaxWwpNGKa3lOrjVgpLOtUgC3FE1O0754PhCEW4ZVT+HJFywxjN
WzIwbBZi6S8uXwd8z47tdChPR4nzfpV+PqvPb/GgCYVONu8JMwTQGirAQAbqL1+flXrbzJ927F/A
zkQd1AjY0qho2IFqLuTMiYFHVjUv8lyEOvLn/aIjg7tuuCyvepmDaUyM7HSckg/e6wlVD74+VWJY
vGWAsMShFQraFD55/UECi5fhL7dWXmR5U4Mje0ufI1/wfs1w28g+S9jbrjPfajPpLCfOU7EPDUhI
O+eAyjqV9wF09s9ncDy618CjvWel2DvbKmpUMyWEuSGKi/Ka5+M/gCzObFV8DECQKCUNbcamnIBB
JHIOHWakkuOvxRsjCuZQSXvjMWO/JlJnFYwyeCQlUhp9GC00bOXi9jLS48HpWjx9+KxjC4g56CIW
/O0gzZgpdr3S6gwh1xYmbwqM+Zo1Nik9MdOHgGClut+f8GFOhzMoCcWVdhWB0UuGIxTqEjrVcuKz
xxCNvz7Dx2O7hJPLNKtyVSzK7gnejr0bid7znfS+dUCPny5bbCZoGBLYbRQnZ6aiAl+ew1/+clwp
96ZPbkkKPYviTAlvXSi2hSQK8o/KPpxFetEsW+lceCvTcUSh7V1Lqbx0nvTN6EmEp8r9ATgp3IKl
6G6IJ9h1aoarPbK6092JMLqnQzJ4gjeAalPwUpbm7BfokAN9K3JQFSR321LD+g/DEWoKJSrv7bvO
camlBoenD5urE16TyjslMDRIBTZezQjtycGy/uyfGTXq3FhQaCcA3S3J8HcTKZjzLrVERGOZlohY
dsp2xx0gZuTeB4U0BYR3KcLOHidKGHxh6dbYTybDmzKx4Hs4qWJluhX2CmL8VeWuiMpqrVYbTp3a
R/HKb0bdms+6LT3NzDfrvvaT3kb5AXIjvapWrYnU775onJntqPdPZC4pgA702O3HVeVVDgSMomFx
64Ek3mCyJyH99FV5QDHJYHYuswfoUe5wSODrO578thZh8zgI1NiwdMrrKlLM6FCHZENjFVwe20SV
AV5Gi/s78yFNYu0RaVGfsKSxgA5RDxr+Ge1dJLP583S5LC6XqVMZvJtMcBi9fEemwcuUQdtmZeRF
nG4uld+KMV68+bc5XdfgzFxrpQbcX2kggs5hAJk6vzhZyTaMiKmj1MCs82iNHAULjTUv0LXndeNK
tS+QvtTv4bSIs1I9gVircKbKcF0RlUGbNVu9UhqBQJyPqSKUoV0g3UrtsT8SeDHDGvCQ+LbBaaxi
pqwX4KQ0LEfcSgn3dSZmiiGaLVFwD87sOIaUn/SOooXApqNTo1SSgOp/3VNMn7ZFL+j6YFfHj98u
nAev8HE3lcWsALQPyn4hr1JW3K/Ki4B4mMqucYckmIR/ac5kEYQ1mlc27crGGXC8EcelatHT8aPo
hh8NOpfxHFUrDm0qy/TKTKnMpqBWUVre6BAozAudV7+Kpw6NZhkcj7BviUBbj4/BwT759j5Z2sZT
OzoXVaEgmqoSaK2rp+gJKLZRRNYW9fZJUs8fDjauCdyipm4wzto+GsNI/b1K8QFtwjMgNGKOt0qv
6lGOER2IMvHj8Gr5/G7v3nFAAt8XxGnT97b07KHpEIX5sIgPYIvTQa6vqf78AUS3sdZMubU166fM
yKNFN0M1oWTPO73O6o1UrtvcMk414DY6butwTRz76pznPESGThGWx8Ya0BxEiwfmS0Pgf/DHYoLA
6qXPUjP6G6yEjiD8Tv6r4Rq4TYNAfHG2uJeCtWdK5re7Dxj3RFDd7qmzhDOH1Hswz3ShQtb7lFUs
zWHNBhfCtO6bLFfONY+9l60saVf8+I3HRnY9PKtpjnf80Xd0XOMJQJqzMMGcqgG2ycYB6kfJp5n1
7ppDfjfmxgF8fwrQ6WIiCSr4XnOd1UBt/5/Jba3ax50g6bpGdDRC+sSxMw5ATx1RLnY18GrB3PM2
aZ02PNXb1f3nHdBTY4V28dfRvSIEzfb/sXNOkIhIFyis54Yx3kJh8nhErp1iu7Y3lOqBYgeHajge
9E71z5L9VzGlbzLzYyIDALpKA4Y8W6HlwvXZ6GAFtsuOhIDvzJFbceyRoRIEw0IaTqWgYmlevI5/
OqTwypzMGX3S5OVhF2lug/Imgbu2wI4HNBnL6nPFCyfypwEiWk8xsX0G7DZb3QxqT0xbhOKj79K+
MnLecl6pC1avjjGyww3zA34fK6JL7aBwbUKOzlyjg2Eap8sorv5c4wF6Wfmh2r5vHRL8dm8FwBOK
zfQ/T9eHG6Z4h7+9ePWQ8SsiLFwpgdJ+7hltCkqQXXhE/f7IZ02oOtGazUGdRRVQQQnNFjD/5m//
gNBUWT7b44kS9owZeJ5AiFMPb72xfYM2wvJo1T9YhqoTJdw9aB1xxWDFDBcjFxfQ+HKtr6asGK8H
qgOUb+1x6l17RclUDstVTkJvw6YqBls/uuJP5AAJALsXau8VILDkU8XZb5nwQNQNnHmk8bMvuMYt
f5Lw31ydPk3bYk59THP5l/qLUA5oxC8ItZ0uEV39ixP0cP627mtDttKhkq/BQL1Z4G9Lgrb+kl/x
+ESxRpYw/jUJhFksRkeCpZ9spszntMZLPsK+5C2XFBYSsYHaX8jlj5Pf4SN66Csk/mEaxrpZR3yo
j4m20oueWKfweM9/5AMdv/mHILwLVfh3wgm5k/4xswCPn5UNk1aevsUf/QtI23ktAUPzYAKM+6Xi
3TS9opWHnIimtXENZUeAYCN1RXoWzNIl/eoFmBqhVcO6AtYprxiz+TMWWOuImWEX9bWzOpQzkluh
xPdjFwfzB2a+VmRHXJrr5HeoRDqaUm23+sZKeFfWENLDijCDeitOfjpF21Kc6hl0C3sDdCcacAeB
EUK5+k90NYPrGcKIdzzdVpn5r10xdXK/+NjrpXfPgHkTfT2suI84qVGBYZCSBzpe5RtpPenitg/F
hHKQmfEcQFhilI7V8xFU5mG92OH7hkvMN9ScY5ZLA1KnRqwPwcIeh4v7ioa5IqGMXxHBdb250HRs
HoHFB5h/xYh2gdjGri+dj5WLG2rfcN/SSmdq+pZg4lHVXdAmJCMyn6edwac1PYttuy+n8vvyIuvp
pTNT3GkAetfxvnOPgYC6zRRCkJWcZD3DdkIuEbI5/FJ+y7tq00Vj8gte1vi8O9qoJBHKMZCAXNpu
2mqK4/zKCEN1nPopsaN/NoPPPEaWKVgVZO7viyqwTS+2lLFtEJ4zVX7lkpW2OKn98i4JVtOpfy/G
iUUCv056D7ivvvMKlSti1ZyK441/p8UnuwHn6SwHCOhWcTRpRVnUvUQCGZNl//wIEp3qDykr2Bqs
F1Qr2b3wiAxryw+VMzbyI3vp2z1U9E7c9JFW38a3/gX91rURxJRXiYixsEfO5UrMCR0j2EIOVtJf
ZsmIh0+sniq+zUQBd85Rt0HWSF8wgafBVKSDFcMfa1tGhiGTqu4Y8KtcK9SajTZFJElrNMNSnzjN
rQBNn61BbP70Ire0IowuaxWEuVjGKhQQAOcOJLiI8fqMT6wf9xHvaTBVeCw/FSU3v7O7nGVuQ5lu
JPiyBwk3lk9qcVuWr0kwsQrvsp3Flr1hejRAdAKVIV3VtOdfY73FJv9GMl+jGM5alpE50tJzDffC
0dtzra3yU7YQXN/tYpUB4n4U5BtIciSaoR8c/Y29+Sow+nFBYKIp/y8WGhd9sWzfdme+1+hD7Y7a
dmhNxMSz8NtAnVTwtUoyLrTOqDDtPlpeYpl4JKzAENoQu4XRfJ6U2hWOI+//h28+f6A96nnT7PJm
IJhNAnfMIRs++UU1MuFNKi94era9kfSqwfOrCmf4lJTOqjPRL6d3gg70n4LamRMaqsqhUy+g74mH
OSGBmXqYmLW/nTk1vUkvqE+91DsLxVFjl2JS+AqDY1+XkOYTEHi6ENF4WKS/W3AcPtzXBRmD0sYI
N7Nu9ZXuVuziwXpIZuSMT05acnPSX6rzZ7WxvFCYei/AHMZwEFAMrC0ReqCGpl+cQk7joS0t4p5g
bdgy50c7u09C3sqW+yfZge9hZKHzJccVf5ssifILAEOTQDVgJ/jipqhe8xEuB0sB9971Bv7XMmf/
B4QCHTsub4+ZJMqYscy5KzYW+tvumj6nfQY0OwVhq5LHJlNxxjMVNrmndrz8fVR/yJVzNf3pXXLz
EsZpIRpGsIN8o88dYm1DGBdnWh3IblRJe/gGuy2tYI1hwuqsbP8FNfyWLaz1WxxFp7ShJtw/uQ8X
sizp+vc++JqQi622g8wlETxMjb0q+2nSInbO11bUQeNVbbydjKZ0+t1HcZvG+0w9gQdmKtKpFd6u
J5vqCJptfIaNSpQW3yZQVfDQ5TTOw+ws/GQE7PDQ7dIusFWmvUR5tobmaD1tO/5V2M/fE/YvQ0vM
0e614M07YbaJR+rcUA9DtGVC/TYiuHjO6jJTnwTb+nJQgjwjIBQQwWo1Ewmk+Oyo/FItQ8yUpXjW
tYMLO3HT41kLwhKn55bBTxIr6QbDMqkePm2d80ydzV19440op8quj9zANAU5036yw0Zdmv0ObKct
wFodGYMwrj71/yMm4C53VNb9gjTzdlcKCWcBDIdqo7Cm2GERYuaSURxOBKYcqWa5FeWMjf+G8grb
SZKHhcMyAnVWrtirDYfll/4GB4ggk78rriLnyK/iI8tdXZSCq51aimz5svqJFErARy6hBJP4IVWN
McPxQ/GHrn2h3/WVPPtH3CGGDPikDM8O8SnihS/EAS3ApC1kEaNyTUUo7lxGoGF5S4ivhwRh0DMR
D+nBNYk0Uruj2TOnhb/qSPdMY6s3TZzv2I5t1RiBoIWLenmxQirBOHY+y6wx0jCSHkd02RxsfBrl
bQVHfN+/WLMgkukpQSSr2Hx5tGvqa/tqNDh/48YfJtL+/u8AaYy9dt7wfLy91pK9bQpZomuuJbWH
CgSo269q2TTU8iL02uqgsi3NzH0LMBINHKVux9U8Haw1xyXA3zW2HZpP13d21k/+6awX8CJzuaDH
vxI0LgsnpMYTnOQ2xu/cQdRLwikI0yAjihHJBkrnX/VX2OYHEiY+pHTzlNFJ9DIiDO21ee6exagF
SiXh0OIpvlZCxlSxzqyFCtlkkZLnA7FIkoVelN5U+5IaYRErpVBIk7o5CcioWhFWOnjhZVHLh+h/
RGUt8VrkmH2SSS6UFGwgTPSmDKd05upIYJEq1394ETkoPHpqvGV2dCf6fMgGXhmJ6GgzdNeM4FQE
njzI/Ypj+3KRhrhvKio8riVWEtL/VWYEqkop/SqVWmxwoaUUcQ8kl5VV2g4NDlKmyanid/xheP2G
ZKVh7UrEtDSdm8549PNiT28wWzSnsMw54Ws462FXlPDI2NXaJRjAHjyI6JVZKy+tJmEubfPSb7v/
EJrfPY0xhlPKKMddnexJiGIXqMYmaVjkD0X6fEkNrb8a0BFzsxJgvpKKHIZ9oZGo22+03eqeDkni
hO6afHRPfQul7phEpkkvu+eVTv0dJVCMQ80JhqOSyYTalPIDA5x4icbnrvSF5bKZbcUHb0k7TTst
Aekti76BmlFyZwKssBfF/PcRk9TKC1E3ggNxo6H/l6PawtnfKZsGkpRvNwNfZElrythfqg8EVi9o
CuuznJ1fQLEe5QexOLt1t0J1/SJv6dGXm3R++hQg2t+6Njrmj+IHZyNI+ZDOit+Vw7HekFH2jrEF
JgcipRulC1084G92HqNb8CcdMvUIlejgY7wW8tgAOSEH1nnIbjp4sxJfQJftAxVyfArxUb12qmyN
8XI+2fT5IFMqcUd61kKJSL6rlMJAZJS2aJ0Zyah8H9strXwHcucEDTcsdzYS5GfMN9i1HVZamhw/
8FdC+ELrjaBwSLHdjFKj/GMrr0ydL5mxJbvN7nUWuDKXgB6xXWNc7u6UCvTzrRMAbfhkbS4kQU1C
L3a0frzVsf6B6A/eLB6eYzxFT9YgCGGazjO9OiZGkyS+9R7lh1XjFyM/t8495NwVE9Z6pwsPa9gg
5MuMKW9q9ZXbJ27jkqh2Sk4hyEUhVhafXFCSuixZeVr7b7hhjQImMozpVnuahP+SpxnIwjEGWKP2
Epr2FV4Bwfbi7OmR6lcREyO+y8Eday3XYdl1FVLaItCgnMXgVJSUK9cDgS4+6ZXTE4YJtKjyBEle
3TiZWEkf1Ukjm7qnVIcdjPDVvI74h9Uc3HA2Tw2rBEslwbK3ILCmHiyWU8TJol+BozJ80CDvg7ll
X4UZv59KoCQSGQf2jbFVwdnLk7Z372WVBr+uUFdy6TmxH6rtZspaA6ivMuOAt6J+jZ4nf3JxtEGF
ke5altFnsVPyjnGp2FSqaq0xeLMDn5kUUs4+q4MoE0sufv9H4HP6W7wfeJsxf0An4C8zhnEFr5iQ
gE1CF8Uyz4X/3HFoE11L+OQ9yJewjIrY7CpfUqbIsHMeglgja2SzEO9WdSyDhS7ilI8uPHlxSSy9
2IDslJvo1Vh55Mp6L9rWix04+moAr8KYW/TlHZwcni/LR1PNmmGUVy9FyHr5NF1iYullIv3B1Mgf
vqoV8ADzx1DgjENN9jxTyYmTu4N7f6T8+L635ZQSZNpsYg3KMzBP0hyJBejQ5ZbV0pV96ekDpHdt
oyUYo1wOQ0dUevtUPEA+f9c9VtOr2mMh09QObNZ10L8GiKSdPfyygGPFGgudilaJlXs5ocmxAI+v
pcq/IQtkcWhm8qDD1Wh6tqcSQOVf/UkBTCqBq0fhQ3da9CaGKjx9mxoawvKDHgguFlwAYr5kgcYH
TQ/yP9QG+Yrqy6ke/9v5g7vswHO3NnWgef8u8GN0mZbC2bGjr91r95VJ1rR1SBjbL5ShYafe5G0U
qQpmxK6gB4RIZ3CVoDDhT3ck4eRXPYJOyOj0KdjFJznDGllgCLIi6XRuEqYunHsMORCg0KFCzBmJ
HDAvgkQ7zkMnPUIuWEUkuPriXmSICwIdciIw4klq5uG4/dEK+xKQdfmbDkUtHMvsXzUh/tUcHM15
+EhHmR/DvajLrvuK/pt7qxsScsT59mXay5fvkrs/bwgfubgMIB82/pNLNmqRQhkomO2Fx+Wmjjov
SBjFz9KLrMXEA+rDgYNNo5pEgsrVwF2s9eicu9sTHATvxQFJDW7rZC+CbcdGjZhrWTWZx5X6qCbp
mvDQFc5//GC4YBwGr5jW9or/5P/d8rUzxrMioeRT5QYaQF2t0o00UMEb8t4OSbVBdCW5i5KJ7/x8
b1TOmsPdhymlEQgrp5Rz14NufNqa0qw3KsZovjJvl5iTXOV1S3KP5pp/42p9smJmHLGRxVNgfd/s
VQJGNK3XIqn7WcjOishOXo4Jo4daf2uFRuR+xwVoakc6YHymivgHa8KIbLxIhxJOkg/an8gsnbrb
bgAdb1Th5rxbffH5COJrOYZz3jz2D3NBPsXGhLaofiabXrbBXl43uGsYz1hYVELKiXVXNtauazE6
PpLjaPZQCrXkobpFf9+M8o0Fj8IOHCTplsiHfLWhdMcjLZxCpwLamjXxmAgQ/6Z5MRJU+AlyU2B2
78z0DUKdm2j89i19iHyhsS82Tmn70S41DrBnaGDfThIhcWfWAlPcCUi5Jn54NsjnIxLq8eKOQ3HB
YamTSSHSV8iufllqTK975dbcPbht9uoDLvUjM09Sme91LLjVCHzjGQ17JUbYx8GIi2VSjg/0Em/w
dUgIl8AjzFZSrcrTnp3gYCSTQ/gR3hhAeQzW/+SPzisdJPen5dOPJ9SB6HqH1uUqrJZfC/WN2Sq7
MoG1YvDE9CakUpxYaaFm3rI8Qvq6QnzWATeuIUzzs48Q2hHHNeT9u+dQ8uiQgvJf4Mwiy5AlSuGT
V7l4e7X0u0swSjcKZ+xHdQeFNrw5lBAPDJfUv7n8ZSPSvNMeQV6EzPEgJP6qtSKfiD1L/ziIwydQ
f4fMmZKvAtiglLtNcht3tahn4rTaV6b3cgjhaaL3U8NJHlu8Pv1zAShuwd2l4uKhSqKVb+lO2Idy
5e1JCgONsw0HF6BXCtWgPAgtBNI741ghIbbGze/XrUG7Ce13RALw14ynu85nR57aQSWc5yvU8DY0
UBWEonMSiUh6SwvPBs+2KDtecQ8niGx6xqHqdaPkh9wvMk81W1uj64i6VIr00XbHfMCMbmHsejXU
TzStuD51H25R5lp+axgeG16AOB1ZOUs6bPqc8zuNqvnZWxD4zXHMy4Gp/6X1Fz/OgfDZWExMasg7
rmSa0iXih52vq/82l6uU4lGLcSjUxbpz4S5T4mb/XdtItnUvNoBHJHsFQrkZgDeHszjNr62wABv+
Ex18VCY8VyqodAjP2VBSdPJ6yEolDSVGe/o552EnYi+fiMu7WRYqLQMgaaV8Ph+FsIkGDYsNbyvh
b3mrmioTehXbemoXNLSmZncWCVwGw5kGEN2u0UcvjMN6apRcluwEkOv8+RMVhYifz6A85VchAOuB
NgOv9uuJoKNQxh02i8aMbjRrEO5qg0azQiA2hIn50V+RtPhGiBfgzyxjf4zDW6WnaI7ghefAzBo8
Mbhx9dWSZY8CWcBfH1AQttRY7gaCaZpEN92AC28/c6ncLFN4t1rpSJ+9KFqWWTSwSt+vrQ+7Dh1Y
t/mdBhFep4b6X8D3yMEg0R/dymmF0vhbg9fh7K5zsK5O4S50gJksSGnEynMtsDzTi9o0gzCxtv8A
xGubJXsyFG9/qgY+LUh4mI1OBnU37Jqu0qGknwJrgeCCufoyq89MYiuZkyqgBi6sCnqQZouTJVNm
+btBpdq1IuJeJ9Qr+ISBmxZdkpNWUTVJUnB8ooGekNPvcXtcpQ9tvLGv0459OtaXCanHs0N2Q0ts
aLNtii6G8U8wqQOgoSZhqI5qCC/6dZreuJzZnlp2tMthu56L+ayhXNadMbCFsvsnzzg6YbkR3tFo
YQNGGby4u7Mwo9vLVs1VoAv/Wp3vrLJXjFAIYqbdHk3kVRckAHD+d/gDegaiBolLdtZLKE+i6yb2
23kOTOZGUoKzbbS8PKDb0HxVRFPz25viNFrAJ+TPAx5k6kHucMCu0jyWp9OxcrImOr5BJFE6T/EG
/rxmuR4mp4wGCiizeolV6ngSkQN2Z95JWlvM4YcWicBgswXLZHSVrg4QMSWy3vfSvhUkx8NScTiR
tXcBvvz7YAvVSn5cSXvB+WNQXKVYVKQJpAjzqgNuls84UzWTRX8lxtS0C/1VNfqoYH910+CB+p7W
ZI0Yp2czb2uBSZisBHLMqXKjbzGFPWN/OZ09d9eO036Kj1tcsfspZl+xrOXG/cuE9xglQ/+Cd52t
fQht6sksL/a41xihQl85f+PN2Sl/nWKT4iefQY3eYzQ8Zz0AX8Lx0zKdWLGLHHZC0fYhlM08hD7d
YowzIGneyIZkYnKYFOYdAgjanj4WyscAae4PCFXQuzhjLxF1kvIGg89n6hbRQNsued3rrZBF4q5t
lrOhZ4Nf3Je3qIgs/EXPAP4Ph6Y0bc1PSsPsuhwCdMxkQcCTqIBmYluqimjhsS0469hntanHme1V
iSHTiebImTB2iHGDzNDAMPiWK7iVz07hzqcjxL/K/fEAu+TmBioxx4grEiP4qsSsuEKVMPKlmxcD
myE6e296u7+DhFy3x47rFd/EMvigWSvxz11KYsPWy7SzJCoK55LiQEddqWSfUv/NGFYGqpkiarwp
brfrgsGJLRsO8t0BNwXzWZEfWbwJCEVPhlQBlqUtMNvPNkUkz5UddKotK2z0KXetu/iWHBhG4MPi
WXPiIPEAwirwKT+uNDMKFjIHXRZQPXFOVdCLUfDZuugzloTrHjF3LCNpI+f8Vqu6PW+K1jEqTJjo
ws86vk0saKGUfhRgV57JQqn0A8/XjBucXFOEzEADyMgLTbFVM4NY0lOlLBrLZ5tb/fJP+BjVO3g9
CGebbP9rJe2g4RgOutfPvwLPl8LK41Csd+oTRCeHkWRHrY62vPFBjXxxII2+RLOKJX2zLn0r5b8q
5DMeYTlWqT+ivew5u7rY3ZdlON6VUq6vGwo/BNahHRbTa28b/EeHN4L0NcspoITHW2gjW6FSUFAF
d/yn3g5cYlw7pcrqzFrYLIhKPYegKnAEycfHoAY+t8VTgI5ss6g9eHNLkuoPR5RYqqa+MngJejgK
+MFT/fWmQyNJOqj3Z5URXIqcAp1BlKHcnlKEfOHOC0uI4K9Khz5zBWO4ma2m7hkj/WrrYfW4zW+7
QmKHew9ay9/GMl9TIU7AtaqyyIVrSbqI4Zk3aitWQH2zTneTq5lc0k81t42BwPKj86eNaKWeNgYA
bjT7QftJIZajwgYxILBFUaeX5UZJejXGLjHSiXu5gbjpL6jmNh9FPuTr6FODb7/Fyd7qNrbIIw4f
ViI9TMHWvIgXtas7gfI2K5Hv3/3C6tgAd8r7Ngq10CJ44VpvMK9mLgTT6OHkKQ+P43znBrV6do1q
0JkWshJJmHGCkiR6GECIFmtIH+Ufka9cbdVjwwDdZvAN9GNsUU+FGsl5YP6x4LhjaoqZy/bGPd9H
i+L/fkoD9fNpZqttJhBpDxbqQ6DgCc/ESBrtOowcEImI5jVAsvgg4iKMsiVs8Z/RgA7FerhvFBkY
cefp4Q/Pu0QLmUJ0nU3gvuSUWKSLrpBsP+4FN1XqDlx1AiECW36sIOsfqCvrwFGqf+ooWnor6ah0
Fa/0U/FThtZLz3BSZw/0bla1ty0Nb7mcwZS7FAyD1tGq4CtMZrGAkj2KQBMI8IbxVF4QYZtsKqMh
diObfxxZpCVB8yOB1dqifIPnzTO3eF4IwK0fwtdMEpRu3pNy0vyXnT+wwTOW3UtwpH1xIy0kqWte
9pfPVPoQBRpgPITNQvfQ1exML/6Pxq0D+3NIRZ6tQ2Tos5jMXiO76HGacu+prB27Q8aYfiYeoP34
c/B2pH6ZUDTOCEmQbnSsKdBDt0YYxug5ecyLHAmiHvK+1jEnKZxyQYszTD9qA+uBqoM0ElkXXUOv
OrHsf+nGFJahFbGeFixJoSt8nVPzfIMhlz3BRn7nkNe2kxC+YDSMkRis3F5rK3Vwg2LDRM2oAtwa
789jEGNO0qhQeunCt+OytNlR+DfjE9feBHudscr/wXZlTfVYi1shAGIgIedc3YieetGYn8Zo7DxN
4Giscpr98m+PXp3msdqlmSstvMaP+5J68X1k9Y3pI7V1tiUCKycYZPEcA0mjV0AVkkJYh3QFKGOg
296giJUUsP6Lw8Edo7v+H2KyiF1mL+Bpwl5BHSFOYBwv6lJaqN/2kOpd9Bnb2K55nj/C4HCMRnvh
r0bUgciCYSB7XUGVGdr+20SofKp4JoFbsUaTQNBgBs2lZdgUxlni05p9wwjYS5rmAfqsDnt5AFN6
HP91OJ6cVcvV8Zb18NLMW/DURo17hxwq7lI8Rocxo4ycGrhzUH3AVYai3gijXiVL//kzl7UEAgBX
qNxZtu3SGdh57FSpFt1o4f6p7WZmjGjlw8CR1ePi0H6CzdbTe1JgO5vgIqiqdldwfOPYgcFPFlNR
jlv/1TKAIVKDDRoGsBf+NtRwNsbosrv3HbADLpAXD73PZjpgWgteE04cVACngrg09vDDsofc5AwU
HIiaC62o4ugV5tnxBloaO9yDRmwDr6eaxqqN62PidpVm5r9CcrddTtcCMmA2gLVCHzDIB0BIqDny
1uFuer7Cr9dRzxOoFT5fZ5k8RFofQehZpUNmsTkxvbdBQtW1+INUNyq2qUX/j2L8mvFbylUET73f
Mhj2hUc63i7q0FntBRDMxG1nyF7P3PckGcgyfFUaThHXipYicIu+x/WjEzLtONwDrjkI+/ClbjjI
y6Mfjh2qKRhjDQbc1BjncUg0B24rG4ZVKJPp8Fg45DfuNk3F3stUtPP3G5LQ1Ycqs7DQYWyzN1qv
N1FSgOaoLq4tz7X5X7P7LSQJ4fdk7ar1boCfGtHELLBbF7bFxczwBWgv3582sinoELij8tsUgrZc
fuSd+tnzq1pVm/vLEF2DCsDY+zlQ+kCCpZvL6OLSTzqzdvcF1DXDnQcgbJgwnTOO0sEUjdV0cuQz
BMjuZHEwMue05IYG3gCUsvCQdPkaM866jUpWP8NoBVFixGofT4XfrY9KA9kgye7T5mfHdVT0uw4b
rM+cXyCgOvbpMFaYEHb65rEiFvW8k7o4WCldLxRSXqcTgw2EguwJre8Y22b4MgrvGscCM47PdU0o
OMDLYftcp6w+5L1MMKWzpD57XNXNrFoLw7e6Gl0vK9ZlDA6FSshWeBj3XUYNJgj6ESqxWTpEhzhj
haVTqTHUZ/4px3bOf5o19q+AWZ4aQjy2jVo9z7Q2hzn1k/r2DszNlmyLPZ6LrdqoE/QLzTcaBvJG
M26hBU6R7Sy7czuD3EddIbsnwCWlJH/iy+25U1uOCj+22ao9/Pwfd8T/dQdWIDCkwvzBUloZC09V
3Rrl+JD7/jRMRHfv9LvgX5pAmLfFcTbUdv3HF50oNBwyMjsw1F20y92K04xO9uiB9TQQhP1669qQ
A+g1+q32x/fCTpS3AulwfRqbCo1nVbs4SC/SAlQ78o5gfHaI0oizC7+W4g4wEosJ0/MWPl4B4CtJ
GSVfFwYZ5W/hyPKjHBTHbW7APXsOPBmkQtNOSD9u3QlDrA/wacj9UgkBRsNXmawYXpm2PK16yTGA
SV0RwuUCGC4/moXstADfoI3D8F9PzivoY1z9mHqekhl6iLAilmFvO16HDmqh1Y7d9nuvfxToNH6b
kuU3HSiGG2+Rcx1K0FYopdqGQ2+jtk4yy3oID379uGB16MoWs0+4NjGPY0qpuW5FmE4TPHf9e/sf
FK8yZ3Yc6opJioQzQYPlARDDjcQ1FsipkbSsAgy+gTXS9kGGv9j9vPyojcZcla8rsbj4PypiuOj0
Zm6v5Dmf/n5zas/wPP5kIQmomI4RSC16EZUXl2J2eVNP+E+3leWARi9cooDKD94I/4XGD1+YVe4z
3WryufNm3nIn+kKqN0xrEjHYNeA+YRbDyTyPao3m9HD74wAoPClO0onWtWcxaqq5jvvxQ9quMXTn
lGhefElebQc/G1NEEZyfd74kr8Ogh+/xWwHa1mLrAQKbBlYjNlIwrjZsfzlgeybvOsLeh4pWDWjl
1gR2y3OiL1HRcgGZotrRe+fbS4Y9a/03K02oavmiuAODThXX0pPDyKZes0r5l6LkWVujKPXg4DTI
A0XekW0s6i6wMoR2+kB9rWM8TOnexG2tK8+UH/GiObAuRPZqUJZC0WLFv3CR6ATUvVW8OOq7MoWn
3AzDIgqI5f0UTMj61XIF5QTEQxypqOhf7gBA0yWhhxwqXp0a0mkLqQABqtCskmvewmNhdWKF9BuW
hw/fHQAvBvbr4cGp2zr5W+4L6oAJLFYsd2zg2T2iJqanCXGAopcexMXD9PbSPgNtQNrCSwd8oTxu
lgyj41wXxouTsk874i5TQQBG8UyfB7kP9CD87mqihlvGq0SDDW5GVqj/qec0nvxmRtfZHMArSFxQ
ELHW+dPWw9RvDIXl8p6g6RwLTulEUqHY+Ksg41FPixOtvB4lhGbvxRcLtfZHwSwCDcJ5g7/QqCzm
lC4GxDK7eYJJbEy6anMGtxiLFal48Urem8+k1k+QDzUHiIYc/jiS+HW8BKxPO4SMHagHyAJPeMQb
EZtoIdehLqGNd+FbOXzn85HhEHavCLWZKH67f1hwyqjFE3QDXlJBla+/g496lyAOg4G5v4ebY1SC
3E0v1IXbA8Ioh98rbO32eNbseNsOQVgFlQCYStEUc42MOcP+2XlSF/Kn2tYF3jWYu7UZBf6wJ+Gj
8aWPqpyXKQaFhu1Rswh7X38LlsNY1nLEIY+X0gJN/QdaC/qev4AOtmDSbl29xjqjO9CdaYrjDSlt
tSFk/imK/7NBLLGV9w51GXAQsjHRQGgdWY6XBOG4eGSAdAecZLKEgpn14KURhnQR17tqYt8vNPL4
7IFWfZQ+pRRFS+E520F4ILxjIoXVm+kFdjbZPi2iWoNnY9aCqb/eyQpzColnJfOiRtRej3SEmS27
OXmZQwqtMMDUEWnV4UKD9lAhlUZlVOvLnzmsuie9j9insaInUKhhLRgtK+NIYkyT/O1EGOF9Bf+A
WKe53pJwfra8kWx/TfguQwvqCRvfbIfEz/wI2pgO5R4OTwx5ExFKB2Zl/nazOriwKwH1UNSbBXQq
EgRzJ5k92Krpc8D87jmNpLgbscB9iQLLy8ROHsTdnnLofB2N9KhkzWL2orEIQdrsHBlWHw2Gv9hZ
yeEgx+CSd1+fB5qGZB2+NXpIyii1FysG65svfzHGYfp8acEKJn1UQxTyBX0V9tsSjWawtMQcfRqs
DF+UbCZLYZixtxZVKzuTAB9w7AGvhTg+VVOUmkh0o1w8NMEakMYejVpjklZ3Te/5fWDVy/el3na1
l9el+UhS8u8vVt2/XHn7jWtggKewKopOzwIcnYpUVExNBCRVaoZdkTt+s0XaRK/e6Bg=
`pragma protect end_protected
