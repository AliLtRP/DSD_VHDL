// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
bg2V/KprEr2jgmyzS8MNA88nSTHARlzA3Z9ouJc37VJHTK6ssfzhFIKv8gLxysVL8lsBrkFKVCNl
iNPHHD1JEMnnLNUJ0tdIeT7rcpuA7KKbgfet5NFtvEmtlTnb8LMhP+jA2SWtQAJjq7xgVSv08QyC
4BSAC2zNV+YFLB+oxuAJdA+CAJgOJdoXMZgeTvh/VJP/KORUOFUDtguFZ0rvjncDUyM9U/63p/81
ra4houHiqHtvFsu2GIR+HoUcdplTB5/ZBvOnfIifysgZcDrUiUaegD3cgQg4et4HeCdfHKoVy8HO
uthl3AhcjImJCAWU6ngwzDCQFfIiH+ITgeooRA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
FGMz5Jqz5fugrMk4zcHD7w2F0F3PUUFLjR5O/gdKr+j3ZvRQmbx4+RdvWE3Lhw1MtmXxY9YdV0xA
gYgKOlgpua2FsnzUvFY+FPM0ZeFHrQdApGyZJIdKVHI9j6OsO37OZW8MMVWCB1+xpFYCZp2XBL2g
WKBTMoyaStbeWhbpPWAh53t7huMfGIyKvjTr+9CogpTNaXgUkMwETCKJY3z2TWjA4eW/OLS9WBGV
9GANRaqXOYahkqlye6ALMurmXODfv3WYVRdX+j+v+RsBC4G2ePUb52pRe0PdE7W2v1UGLs4mdIw0
NTqrpbN8Sw4d/GsoyvDijkp2kqa4QEiK4DTt583ji9YpWwfIB8PHvmaVZCJRH+sBK8OmITisEBpi
MrvlwrXlIsYsinlz7VUUkS++op5o0wVMJylp3w/w2AJ3Ko8DpVKFkzwRzXku9dSmCAm5alZHjF14
Z97o2GO2QUNoZMlcLmK/2htCzKBPaRnOYdrzsSBRLyg4fT3vMTJceu0sY/0Gw2faFkiCIXAPf57R
j1piUIPhCmBUrk4i29M4ZI3GNHh/b9Td5dgu8ZPKauzBgj5NItKJtjR6rXnZo//AGjjyrolvWW2a
um5J/1G9vdZXVyCwu+WTS4soQ9TGsB88RorrJiItVTyIzH69YVfP/j1XQOZDjSQOl8qed9xnaMNI
iIwhQytvs1cI9X/rRMF8Neu+i8ElEoE7+ufbOHPzYjDIIeejoFY936kpo9n3JqRsVlzr6noNytQ+
DtPhp+OOAtNH9FQnC1x9PQTIQFVpn8UzaMXyEChY19HOnYdaF+KfXvb7yOlA0mOEZl7n+KR0Gr1L
F6nVQx5wZnPTrvQzA/EpcZ4iGUASdCRcok1fZnpBqfASSBm3MUxDGsZZxbtYPUY3ab8YN+VtVNG0
23Q2WjjMAvhlTcnjx64+6WQpTOoubGxCd/0qBc8HWnK1k96BbwHBBz9GQ4O7qAd0GGcBtriGnv3E
9D3AgnZrXpY83bSxb82j59/oALnJ3U8xG/gsYgOuAFzPcaUsQJFPSLkpckEcaCC2RBE+3iOaTkhF
FLZ0ucnP3Pdui/8iWLyXqWYnJ11krQxOoGEOlcaDEzPTrkZ1eRD+AUm+XlHFTDGWwns1B+vrsDOZ
kNM8MTugMboddUdZNAoaImeLnU5869DFjJhbSXTUGPHs1+eCgscYJUsWod6HdOVz4R6x8cipany3
Cg61ld0IAWFZn9HUkjQd2xY6Ci+3Sd310X7/ozlFK0drs2BQws8dpMSXCl+emJctZVVxvpA8gs1A
K99SAxbp+pDRduaGA+dKwnaTYwSfxT603BdXmlJFX+/5f/UzKcw7YLo9ASnPrRuV2mD/QT3nGkfY
xEsQbnf1Dmn101qvG5zgI3HXMSJ49VQqfseXSGjjKtozF3wBHwHv9W028VTr2ncCLrlGwWyMd1Ns
4atu9HBS7nbW8eUHEnyttZokuM4qSsGJNsoGb00DpxsxFxOl0XQ6os9xBN4B1pyX3PoZF2a3lzQk
0pW46XrIS7MM0X23R36B9l4FBuPkScwSHPXmjEhnxy+0WI4QkjS+79ME9EbmpW+XzEI7EudJtaO3
yEyVuT6AvdJmin00CSGbWGSjozQL3Pd6Oapn2bm94e1ZgTeqXAaPECAflDYzxStWeYE5TFIHIrNS
Ezp+VixL2Sm1HxoJk0ofRMPmtwqx+ZQ9vUwXQKD9jteHzeHsjvJBafjLBdhE4vPZhmqWJu6wfocy
T/VZnLRdjPsUl+rxnDogb4OxEpRjzMyDm4qWrh0kfpFIBdeiVivWjgt3rIk+yV9LGdg1KTBb852d
Exxe1lYZZez1SJclh4AV25kRVbAdQf6VJUUwQcl1j4SdBTbyUgjEi9MhURKhlgYcqnxvjpdk6Rxb
b6zhVRk7Gdw9Pp8xhux95K6UmlEZewO1FH/Jt+CIP58V0b0/np69hdmiHYcoylCFO+QMYhG8kuNI
hLvb7lif7kMP+CgMIWdLRtTny1TJYpQsgr02ow2rLFxgfJIh18XZeQ1IR6JcGJNeV27UqsIVEHJL
rXkW/Qr8x4U1nBtrbM07JCh22s4G6jswCVRRskXBR68pjCdPBBW1tRChjZC6XTIcb9bCuUziVseA
0HQd0TF69vj+j6Vi9fPq4s136PkEQAE4aKiABlntWvru2vTBzhWSNTyvh1DrEWrFp9QSRCEhiz11
zDno03MNjLAjbPiyfPAgfNoY2jGV9/mQoTLIxXZOcAZN9kFHkCYZOQGsLNlgEuiwd/VHYcMVkn1L
St3m1ytoRB0ao4QqqqZy1S16m0Bm9rpzw+KhKMahQnJVRjZkogd3DZTA2aIjRwQwZsJoElSl7hE2
JRuIigzBbkkJ6dcgC2GwsMd6VpGCf+xHYg/qHHIvfEfEKudjmhHr6rLIOuSw+tXlpfeeeOd+re9O
oiLpJdKXjUR8w4R0qbX514pDFDJylAG6qLHp60PBEfJaQdiRPv24j8r5zIvLuc9ORkcuzJ7ectHq
6+XeKbPr4CbyNYi+oTyID/oqPzIKGwVrP7X8nABtJH5UW3FvexT6d2Agpcpa90GngyGP5eowntS1
hZPwYgHN7cHvRDEJmCEpSjlHFfMeHQvQBFrwIsEyHOHx2Cf3RFTMgKk03H/a6GitVEdoe8aHmOCu
FmpBiQGSPNSogPABKRneYMNDTzK26FCg/NuQt7e+Sx/mbLSsdqejFXiDHp14mVTFkXlMuKuqpadC
1mUBojwI6crSlHyxJbxWuuAfQUeDKhMaL3qyTOXhY9ZUSiGC7KFExfZPxrDAW8XJ+ZOUeOx/KB7C
UwBFtwIVEAesSNV9/5FrGx89ag4J9moGlF6DuE7plPHMQLBxu0yG/2qADpl6vS7jX7bVdzNlffQ5
TpwvVR4bEZPtPuc/CLUrN0MCEPzIlkgY9gD8BYLABkgksV+moQgtU/vXa1nKzCmvzE1ZyZrfL+L9
eEuQYdcUTjwOJUwnP/p09DRq+6+anHvyz9Mpr7e4/RksZFEWDOnZXo2OWQ0z7DEzgAtvZ5kFgNl1
i6gbAc0F67h7qvjZo8UZSm9q30db282sS+tEEIFz0D8Ry5pww35e0MPveSfitzuDS8Dw9EycAXBh
HnzCVOQl+WKovJ0gtXC/FQ2VeiWPhzv0IMpz4AyFMb1e62ZvEu1cGZJt+j6a+Pqz43lnqfqOLHM1
oe/+sjANyACqGzKizDU2OuFftyMcghpytvsqEo+8RgDfjsCJQMyWW9/pRedKE9wX7rEv7JbFWF+c
J11U8VR2FztGEsSIyVXaLOcrDXP/7u4QJV+InPd9rtS5ZMQ8HEaaUbmelnx6TDtAS9j6wU5br55x
j3vwN4F9QPckKNWtJQGTAjCjRBmr/l4Ez0/Fz66IHw9L3PrhVbph0Sq0lya0zFZbPeQxVhFf5chR
GEZoGlMK3OzlnKrbD/6IPAY+kuDfK6oZw0ZxxZL/PRiMAs9Z12Vx1gW57/gcnPrLuljtq4iGFeaO
/ZZ9z7I0joMoR43Ck9X84Lka5tAr8TOr4ViFICSIvCQMnDG4y3x/kc9v1GLJFG7eMejNATIs3zMQ
v1AvQ+k1kwENTPD4rEUXKIq4CIBo58/E7neBtG/QkqLIsY0RlgrR0fOmWNMqnbI7kGz6PCigTXCn
RJyfzZINdrgPbwbTs6lHK7+UFwhPSoFw+7tQ56YejgK5DCA4N4R2Rya8HTuniFoQpBl56dTojBoH
FOHvUm9RY2Bh9zyUevXGB6Q0GpJXoDaMKxT3G4QqTj42yy2rs19fkUsu0s1tpNh+xfqvnGWeMq2C
AHAnJcltOxgE5zyKyexsGUjhTMySoreCTAi8DJiGhwx9VBuHymsdhNUzY9+a3a9scWnu1NQelKPG
KKL0KOEV+J+/fadVhwT6N0+B1KWXhOQ9SFb46keLjLAKiX6uT8U/mPS+H2mGGAtvbXoPxSimETnx
NeZwyIqcOneQQSTfmaNdOJ418ihv68HVdtAcMhfCb3j8DwGMMUQoyEW49RUcinmi7XsW3w4Ky0oc
6BjNMdy31+D7mN2+gLbQttQjkg9O+cIpOJnmSWFKaFRG+3QGfPV+q9tE85vykHu2k6haMJZ3fbsv
3UaYysNyOMVjFQXqTkI+Tj8NmAfioILlPHSmdQ6B/6DP5tdKlU727LbFFnVT1OjzNh7w49ba1aVc
MsfZ84VmLV5tcvUUgPpbeLCctjv8EbE4vf5zomCsvW6lEj+DfnK5rHUoTJONP9/At56LWn5ZesV9
6a5IJs1cQV1aww82jllTgCxI9cQfcz1q8BJlf9omvM6Vz8ex4r6Qg0hvUcxuHS7wv0dmtl/TEGgE
7toc+Qw+f3WrOViCnDDxmt4twezMsUk2OhiQEegJiSO2frB2b2Qj0MooK3gOMUxyger11rCQ3sh9
9iLyUpkfpm/ttvn8GBOzOeY1z4Tqo9Z5sKu+4WvXhW3hYUKRqf5O9kcaw7G0UQBamaPpEdtKak63
NGNAslT+jHgodUtIbg7Lb87RSoQhFPVJqqONHy+t6tWOgX8WVkiFYq0gAXo5RqxlZTNDF9tUmUQd
UyeDSarhj4jtsfEyf/M/taJ7B8QpsMZOBvcElARh82kqAGMPfxxPcj5oB2jAiuKdBURSxnOi040p
2HPJQC30IxSfuj8AENRSV78ZhK4Sn2UCDKveVoa+jbmn1vS1ipt9DAO3k1UG+lNoOyhpA+E4Te3s
8lWs0hRB8f9fkZzFzVgRm/M/GboywaDZV7Tezo3DU755X5oFpyYlxpRntAIookstRg0tpgL/bmfE
WlXIxIvOYtdfNzhhElIRlQDzX+aLWTnse+KPrdlDwsGLe5vHMss3PbTWlOQS1BWJnyyZ0KwDyAg3
vMq11ABPX9VcBTBPC3Uzpr2maSuGv+CUctDl5MVPQPkwGKVFqtB8G5cMf72M1zzx8K5HPovTXthV
jLjhrMdsQ71OCiVBlVrczpe9KpOwJiPaj55+zMQLs82KCh/76QGya9Uv+fU28Ln1h7W37L5EUPge
yP0qxnutC5FKKF5pFadwGlBH8vvjjJyJJCdNf1qPV9jew5RSDgo4bmshlIFb+5EcGrTSgEv/P9IZ
ylhdGq2GoQpggRKZhu8vhJjhSgPIhn/yv5vawcxB0LxS/k4Fxc1OTiywhXAZnD1qglzL/3uUpJ1M
dZLrVzYTQmELUcyFp/2wp9z0PweQLh/HU3d336Qe0mP71ZKbdZImCqC7tBfIMx37Uc5qZ9AffyAZ
Hrhmj+hQSjH2hT/W9SjmeRI6JjFsPrkv8AtgZMICAbLByJJDmdUFuLoe7+KYnETsNRxOYYCFO7Bm
6VLi/ayNGqYfyxwXIBQQGGXnEJ/QiGKZSTnspQcBzqiAlejAh2tRJPsXL8Mk15jk1xa5A381WwYa
RtWX+/N8PPIxws6IHi6LfMspOBxSZXdq+lA4gavaZsdX3LJq8j+3ty3+zVmmXfnY/2PFgXnLJVc+
AI/RUdq89Dv6N+zn9LRQre3uERakvyVsyneiefL5Yixq4LebfD41VfuSIao4Poaj6wjjIHq0X06N
+tTQQZuzALC1F40mhWZP7Lq233JuPBQPrZEsbvW0y3PI7+S2/c7cPH0/vcrXIqgxT7kmDbPrXjFr
DxLRS58K8J+ctvbo/SOQDdVhdKxmhNDo9RS3KfYWLaFBYZWAy6b+Zc6Dc/pW5KixKJYQQhyPLh/g
sJzFTGUDNGcBEV5eEHLnf+9Gmta6XxMBSWBh1pyFRqiFUi5LXfTfTHcEnl9wVk1mmt1MnQrhrt2v
zxczLphBf4y1MsfoJ3WG2HYdBZn/E+1gXkL/Wl1m8pWUnhnnpTrood+dplSQbpDag/toqMFifvZ/
qOqOIWYfwZiY8jBGMKS9XeXealx157roSmK6mA2eepCNHT6Z4y9JXrNg7Ntam+NIXqkEoKiFj7Mp
kUPmHco19MW0Qd5auGJfZkykH+x9i2UlR94mIQTJsaurl1KamXegwOccwB5BeRbLrB47SaQkTPat
TQJATaHoiRQa0SWTNn+WXA2T9C5EsPGOOzhR7HKAMpSDEYrlRnvW41dl+e+fJYu4uJSFH8PIg4/m
23nAg2h8C+25NHXIHbLfekSeHt6y94O1V3E/tvL4nsTt50XyM7u1hyhJu8DWW6rBcJ3i1Xt8O0Zz
HkTjS1xpi+g2WT2YeMMi5oLyhz1qwuJn2aT4YvakcYk8Csl5I4GwWwsGZouCwUbRDJNDE64nQ5T5
bEOIVbmk6r0t1L6iJj8imMQHakMO+smHpbw++Ufe+bVzWcHOAVGwAjj87ciqiTp8vVd1TivIWswT
CgALOKmnlPlYMwEJKwBTssXwgMQOIxWyygmwyu1H5iHWVb1lpci1I91wn/4oYeYCD99yOvEaaW2L
wbqeHYCytxgted2G5VCah1pkQiGZiVnvZOTEU3e65VfrBz/tGvjA/OOcWYtojNWayTLOHHn6NlS+
F1a2zQI7gu0MH7gh2TPHeJpgVGKsdUzBzp/AMN75w46fBZiW6EUHfnxdU5EHhRVvI+uBctW0yOMx
rMDNVrGB3eG7dpJpjQnBSv3rvCQ8RZDQpeNWv5YXcIdiBuedOZZLu5xJv4eVlfs2fzd7j8A/SDEL
nqZ8hA0dZRRGNK3V10o4Ii96VoYTtotZwARXmne0krIIURlCOF7ycOz0Nq+LfINAwRoyFWQ1inL1
H5rmmM3bJHtCDsFbLTCCeYZosa9vtwYjVUMRt/W2Dey0qDE5xpnkd2s6lwnVY3pMOBlKwWZWlbiX
B11OiooL8rtTsLi+y7XNw13NPJ1QfzMGstGzoRdXAtzW6EOXo4rgv94tklvNvRHAzQMDL5imYH9T
NVQiN5WuF5ACTB+8YzXvodwxGg4xTVkry4Tkr8KMp7JXnwX3v/2ExnXrUGpmD9/28u2IUTBkXUoO
qZ2TTteqnzvbP7HcpA4fUkPmlnyb7onQmt1xT9L8o4vWfXDW4JCQBbAjfnKgJbWghE+xDKIpMUuG
X0ueV4QgClu3k80EvfD3CteFNMhxn94GnjoY56iby2UHLUXC2pjo9VfNfLmwt6JDTf7IlBOpZA9y
YxWHguawXgtDDAQZf4ydmLkPFjKrfkE7hX+6W2Fizo7iSDbNgLqNifyctGJZVPX7mv++PS6e7aJj
Lzr1A25SCOK9Yl2Fwc8vvCntmZxE3SYVBTxLRm1xmIknjmAFPvuKGF3w0hA+5VpzVoFVlGo7LesG
jisVpjz3yr7GS5QPZoHzWT9BV3Dr67kcrbviPauFSaqBgzFeYVbNW8ZhMZPkHFCz7OEAREqMKPz3
rOTh+vTI/qjUPVpEh3M1rLvfoqdhXPIdLEPMAWtUzCi5NZ8D4fkT+tAXAVjEsmSWx1MPRb2J1In1
/4eOP1hONcim/vh06ch4EIUyrs3cF7/sdPxtajrZ42UL12t5GQ9yzr7fQfe1g0zArakJqP3w929C
e9K1AUbcnQuWzq2mZB1bUCdYDpRRX/+QvfzITGgZ8bSvAraKnV/iKR/kbKGo+pLnbtuhNq9hCY27
DVBPQ0p5P9NuZ45EAo5dEsFT0y4H5L9+mrhA1X6nSZ4JJOWIENSZBuAwNpLV42EhW1KPa4M7CJd+
yIWt9+5Tar9uB+OrfXA/731J/fNCbt7Gr7AopTcqf+l9U2FpBF7UYCSFSpNAEIGR1Dp0vwqo2bDG
PbrUdE+8BL7weqmLM2eJ9sxvGQU+MsXlDt0/n6QgPwfJ3psIDnFVd1nlCd0xcrUKPRLvbxb+ruPB
mNe/rICyU+UZgQgZMpAFd6mVk1TSX4NYjot3oYudTXOeIUIiy3w14/osug9k7iK9NmBh2STlAY+i
uRKblDqVUSy55/pZjbInFAxca4YsKWcXIC1bXTSFpj1MiZnnn8t5agnGvg/wSEQYhRTCM/2GxqOW
PAm/jiCgChPXTVE8F66JQxdVs4+mA3UwkDg3DExK8c5sdhzucEA9l9XxnCgsTWzflHUWGIux2noi
eF0hYTYrDgJg96xUZNARBkf5TKThIDhilV1dup7Beo/PBKbynBjT4stoPQJPTmfJ8z02WYo6uFmY
aaiFHpHd+cjIh7d86hbhqKjXLdpD1GkMuE7+kMEsk/5qhRGj4kZnZvChujuxntgU+uBCHyCymbKA
WNtLLvpKDmMFisxrJfwmr5w2h4B8tLxwG+4HMtxmgymygCGjOGXznR3woX2q8sHUuhpCAaZ0pVPq
BbdMY8Z0rN1xeEHOrvqUHQP1XZA6WeWQeHZMeDg8KVRfoIXIXH9V3SBRFn1/cJeDGq8QEWrgPnok
50tIO/XIjnuiAZijjUCd/HRWmKO5ZMwEQP38ixkD6X7vplRriraXZZZJ8UoRrbzjuiQttUMwLlSJ
O+alY6HtVjmvWp7kmxqecLS5KOKQL3R+uy3I4I61+myr6Pa4gIjsSeiH7rBV6vg+oEqk2ovRFnF0
po/nBc3JF6/d/glHvFeSXGrb61027qNhLNVhdv/N2Q5fRajOO2if0sSteuBS16ByWi9Cixg52zUZ
fFc1y3/g7d/JHCe8WThJrZOdElzkwv/dqivaYY42cAt/LNOrUpLaAcgQN0Qps4ZIK/45/zt65x3F
Y2MD0uIUxM23x4zTI0T5WYppmXI4Aq0TRZM1Jgs9lmGUjUIGxBi7dTEtSMfsOz4JgF8PXOAiBEqP
RnevS/Y9q3FAveEjeWpE2D9CClVIdpTE6Dlin0+YyA3ejNHF7ET84hPvG+/gbNyy1Xz7cJagWa4n
vAKu5sjM231k3Jcq7Kr9lc/QVuNPFb2kGOtwVnpJJGg34aOkSzY/ObRviml/h2Ah1MB52l0yKvvV
aPcX4fAGDFce0KKsuSZeW+bXF2CThuo1yJGZTkety/nfL9OQRQC9NtXRArOMJIsmMNwT5mU43NYN
tfAbDr6/iCDg9B5YhyKnqXaSlzNwhXWEwCINxdtdbofdrcXJQwMomULmXmQZNvTSruslQ5otyJMR
eIdcKILScJrZyoTgMD7QgkEN88r9OZDt3vrVVreq+7/lHx/ijqsq1PdkRvuxRmPHeoR2oBD0KzE5
tKeRO512s0rQJOhTSDn6fa1jtiZ+yS8K1b7Ph5xd2wXs2/oqziRjsJgZVmQa/rVlXz3Q/95HI8HO
KgroSYyQ5/8ljF1tP8Tx3MJuoMxUbv2IlsqrLSSQ9Y8AZL3XzdgmMHutpD5VI7iMrllDPSxcVWai
FR1cvtZfN27pxPJ18krbKt+floCIqVT/fBVZBSR/ysihvxh0PkAOgihXNp/h+EoN0M4W4K84YQgx
eZrhWVK8x8R69VyE7UYYoEyzK1xZP69qISurlU7UqUr4XOs8Tmw5CWiBE13OPPrWQvnr8Plp7Ezp
t2NLykZQqWFh+/KV2/6MMrTUtDhpmb+rvL80QdJe3ityN1IP8DL5kDFJhRG5Fw8nGucK+ID3/3wa
yN3iHZ9YjxrpYjHVuCrdkVdVRn/a+af/CaY7I9M9NUCG2QuMZfxBAoWvT5mis974Ap9W7w6mhwAE
3Atr2vO75ngOjeKyIPDqTtULkQvqyQ4bluNwrWWo91c4u6WPYIxXQgsc5FgXSzQwpUZsLDoxDbTV
RFLaSKEMLTSAUWekacECLae38c5JEg3lM3ecJoeLQaIIOyxoGSjiaMb2GeIfye5gPKVXWZ/QseoY
Ez/Gdre2iegblc/iVsoTXT/djjZ/40mKzhR5fVZE+Z0IHiTE2LQpodhK1eWAO2TsAUkTnRP9FFOH
a4yKDjahQQsn7xKVFRU+L/DKYZfOvizJ9ThiA/LAujJ5dpfC9ookLzneJMZ2Y6/7XR0dlyhAUJ8U
J2kZ5ehB8NR4WsRdqo/O7m+NEl1XhhuVza8j7vnrHzx2B2DLMa+tp1kmxD+nOtBaFsu64t6wVtYm
z4Bp/LuT1/Dvb9isYkq+iCghiQU9Ws3Mn0aDMckSZTe+008z9rlhArJgqKK8aAxceRNXIZHZqRpY
AG0onJgRwgDKC0o6Q31Upfh3yPd97Vr+X23vfu+zhsZoQLqNO9i70afqCJtka7PBZ2T49S/D2x/I
jSuCVmBbn+Fx4EOtrkS3m0UkWYx2zrs70SU2kegxykfvx2bWMb79yyahumRcCM75xlqQoy0IQkz1
XFbrhx/ZzMzzm5HPh6xski8Q5qh802qLkGTM7lWdx1oIxFCd1rp3WsfhpwHm8OnjMbfUEU5YkgKE
dTADCgVSq7MLK6t9i1LdnPTMnijdaHnV9KRbtL6ZWYwRu1ACmRnibelA6dHGBVG4swDdKvcEi9az
1+pE4uQ8zvY+gzgga+WV6uW4ywF0Pbjvo9S89PosjRjeTPp4tLntQjl1VG+e9sJtVW32lxWz2tHc
NgoA8+NOiOvkxGhjwiXjRwSd6IWlGPfgfNsI8M/Dgl0wbBJpjPUWsIsSUw/bbk9AUfpQuv4kMrea
Jr/n2TJBZv+1i4r5r9eEqLVkxkRMbqtSThM52x9zmNIfdzUaojiLgP0+MbrprExyZocFY+OO8KYR
IyduGXm7KE485f0qQlkGTUAX6aPXkSvrsK5fBBCuGS92KBVrrvHIMbnoHSzsJWnmR4N1C/O79Pry
SgU+RfF5AogRhQos6o5VuDnjv/iVv1EKwsroeWYMLP1D/Aky5gNHNxkV+OZtFHHYreCkj7nGf3Tu
odWKJ6EwCF9m+/L/jS7GPSfzjWgWd/rQ0qRaH8QFtPltr8fNmFan4hxVHIbW9LX01Kc4ah7NixMl
GdxI5ad/1lw2KErucR0eVMB2KvoV57YCwMDBVTw1BFXXT6HBNRwQF4oMhphxpyfiUVLNyX6SPrkc
+rinkjY9vRq1ZHqRpj3cq9lOclU8hIVdbYRBi2F29prTf1gFW8nFUnzCtp45GxUQ0pQLuO6+BuNV
5vdZbouEeO8AOu/e1BpFDDjXGQhHuzJ6P7LT0Q9fNL4u6XTKeUl4n+lQIwvEFvfluq3fv8wxxJxO
cYKjCa+BB7fW1RhDucsPEXnkjZ142T2B2jXaNKwvR6eUqucmxoikZTGeb9s1aBIcpOVI3/hAl4RL
DeMqiPNDiZDMdHBg69icGxAgllA/BCIid/ww6TANwuxwNuMCCbB0Zu/rMKlfgmCT/NXoQ4isyBNS
UymYFsLL43uKdLHge9Ujku2seLGAbclGf8/riqsnvomUtc2U4rDDFwKQDtbukFVv3sm31iIbrCoG
viSvOB+07gLlLWvbB9mTS85979hHKOYVQzNp6y2phpWvxaUYArwF0jO+nkcG41sQVUBpVY4N0dI+
a+CjyVW6S+vyNosxAxPWNEvCK/lVj8YD/tC6C5sg8ShAy0dOpwlbgjJRK0hrsJPn9wJUq2u57FGx
issD4VNoxuRyO/lDDQuB0rd4ENvqA0TS+bxHCUn7vclPOZXwmocvQuprfxAn/H2Gly6V0FehcbE2
HsvFwYMINWxobUGUMeOP3PwnLaVqLTZgfLKyfdilGp5U7cfajZ/TJDDciZpJwBTr48GRoMNDNN+j
HZD1zUq8JLVOP2Y4jMFlM8EEKYILEZcY9lH8JQQwIlUxFcuHe1Sgquwr6+afnY9SjQd6tNtf7cJC
RrXn3CWeZzkdtlMuBZ+lKmZf2GMHmRlWcUSK94akA1T8rlUE2P/5f4HQxz277N7AKDQp/YBYnSKk
FgNB9Nifce7CD4BibIquqSJ7HXdaVTS0oIRtZWvbu9gTgd6f4yWilLLzQnemleXqUnEhDYpYkHqt
LTYIhZ5HN8nci+0nFpdn8pLGBOB+QD/cbqZGJwqGjCaSAeXC8dDmdU9LBzS7cwYFutaGjlFEXPGW
PvBE/aneSAcbezbvpq5UuYQs4Ksux5qiSb06amDeVkyGKfqsUyillFY5/p06pklmMhc7/5r5pq8L
nYM7xYldQwQ+DGAYrR6CiiN8l4RXqtFxLjzGHolPaEaROIrhg2B9+p1RtmbLApSFdAxsfVYZ8C/g
1WhGlPv7uIw5asdIy+WE1xBPPNcNb3fCuYH9Sq2hkFx9b1V7UKv68KB4Cp4x9lBESC2mQPNbSZ2W
dlofUNKESQHr/cNVCOzUA1Zhhi0H9AF8wZ6WppfON1XkFABz1wg7TBZuyNfwxydJ3N1mXaD+aJmq
lzEURr1XEoQnieBE/s7IiNPzU0sUO7NYmfNIQ9m1+V4e8heB0cRvAUuOibgiAFfgVTxRTrf6QxQ2
nY62dkv4ros8E8yN/4c10X1cyJEruCzP4Yc9ZPToF+P8i95xLVcdw0hKKzLW92r4dKYQOgyPfw8q
9M4+OzNl3YIND50WeOXbSQkrnqFbX9KRmDyWe+4rwf/oJEfu7EXqYXj5PW0BNQb956fmNNcpjAja
Sqg63r65jiYByLCxU4KOYSsUHiAJmAJngPdM+RG42ULYlcLQzjQ5mge1sOTerVIHneWUxKKMflHO
ssZylGGfENICJEEfGuAFWvGXHFTGiCQOsKBQBFGwBzL99QMWRbCPugdWACBFjbT8ehJmior8twcD
Xe+bg+tcwtwhA75VpIxNmjdWQmPNPSrFRWlD2mEa3aOzg60V187KBjDfCw7Md/u0cEyHL1xSvE+2
x3B78GYpbLMgMEaTiq/0SKiNrTtYJJtrY2c1K8PQp9huL/jHI+Mr+Za3S+l6X6liiVSe3fNYBu3Q
kVLtCU6YrWhlXHwUaZtyvbM9hk51jgBH+B5xUPYUxQ2bXmlFpKIQh1vSpXQGtgmOQsgSXRfJIS1A
cWSv5OOo8umgaC61PKF65KmriEPP8pu1zeXUmyyjVTeNj//hOJnrKsz2h/rTQAtfzBcK81+w5zbD
fm5wF2qW2ZSOi2VR5RKPPUy/hbPB0yae/9frMw7jPMKuI8hnBQh0mtZ3KoUV+GeTJRYn8wHy2gDJ
6GZARWbzN+g0cUWFdkaDJ33mN1X2oBsxneiAPHhAmH2qc/+T+Z0FpwoaKp4Y/4oF0dat6ABGKdH8
1MZcU3bepY+2erTQZK+6DWSsAUowudbhFRMn9qXV6uPvL1dpVDp90cFkKSO5/ZExrU86lnk/bpFf
qXIx07QnlmBPuuc9xE4gy2VYIl9BbX0/Buq3g0rG5776n7xeJ5Dh/PBGjIVE/0FZSKjEFtMMc+t2
xGvmvoyw3YLH9Fb2tB+NmISjrSIFspfonxqVLB1GY/A7iKZgAIH6EW6aO1O/7M8rClrqq0XxtzEP
yxp8iX4OIJ6m3eywHNu6sSTFeRl0f2aWy+cnXC14PrTBlMQcRDch6fEajY+tIDGIwOHzVsrPIm4H
fHVLbbk4Xy7zgKFhfpKoSmhYYNvLzrLAHqpynK2hHA4tMuCe7GGXiJ6OA24MJwqR/HXwH3+SrJym
1C0u7S4s6kZFVcSgh8XHF3g5UyD4oiPKzbpIJkH8SIiH/6BcShF45TA4xKagKKeU5mTT30OkZCAx
PFJUYD0nYvVeTLEl6Akd3T/AhGMRIRnYM63jrTkFNp7W5arwqWZoWqfF/x7k1t0IQuuw+vrUu9Yk
zNxpm1rPQl4HEhhXp+UfX84EA8cuIKzq4SnqW16xn1BepHTgCkdslnFrdJFy9uhJd/fdHtYjkfy6
w1frUQu0JxsyaQXt6ybvZPxqCyefuvEzxLEB5kXaSICR5mPWGem7KQ8v/JI6N9Snrhd8oDMwMJ/N
tY9MeJ+8EPaVlGG/IfENaPlJRHsRjUlF3b1dwf9j//BV8yh2HRvDtjZqmjJ2zJwi77Xsywbq8OUI
FX5us7jBEX9R87BC4f49omMS3q42j1OiukYzM9W5mYiLWe2QIPdsH8+SKmuLqhOpE09xIXFNSbGC
6fN+52Z1pPW8yMdUcV9bHAaiX25sW96v/c6firyX25yQiIG8oEAmRiJRPhPGF/+tHmX1RtJDhWQ2
yYRG+OjaMQ/bbJYeW0H6URKkmFNOiGimWbg/AdN5LgdY3VktCouhy8CRsyJ14x/2bPqHkPr6c4mL
CDBrmwEfsJezpJFoIEquQqi+afhLs0RXlHx6Ym50XMbEQ4geEDyqU7zsS0KBBTbxlOUD+bSDLcwc
lWU5gTIiac4lgY0L27KNWDg8fjxM/YNyKhBORDIXK2pv35q4iCKFtDWJ85QzNjdwQ2A0PrJRfoiB
Mn3mvnWbYFUtLMpsnLk6vnwLpAer1k5HpCvw1QQ25Tbuoc/s6cyDZe/hvA4rGX59pJDawNppfCLv
2fZ8eAW7+yQ8a9PkGfeopvLkR+vOhaflXuoFQRcIBBtqhWvnHf6lUzseMX7qyDkZqkF+PUhLFCAD
FDcWz5k8Tq4rQgFU11dly9R3sc949OzzJb2sPike+kU1RQoGWjbPaMCFFSwBRlsNCgmbYz+KFQ1Z
zr6Iw+r+EMmahNG3QGQtnLIPl3kzsjQuJBelkQj5OCffDIRTxtPXBF/WljMRj6oN09AQ1MRq1M3Q
27IaybPDlXewBpx1vODaQltO9LfDMf6182OHQdjUnAWvsO3N0kQUyOSUkGj07G0heK/oS1ALO5mB
eMn50yVd0Ovc/V2/dTg4+Em436Yij3KAbzedNvrHAS0RCQsjVQRKaVLYEfPlc3bTbsTX16WfVML8
KkA9qQXRQEEScodETU35JyP0fIv2DKp9fwDCc+MW39q5EhfRGi73xlad6QP1tlK2TOwZCTpHCKCi
7A/OBDUNX011j9frZEJi5tcxAp3R9cuRtPOomNSKTg6ZBl/DtOTJUAsJkefa7C2fk9hRk87frXnY
K91Si2DDUarNNRH/nGr0r97zcCmQkHXmsDZxTZQgbzroGpOF2VPm0jpvumyr9bYtGKQkbAyUnAow
/GzeBlpB/axchv59g8MVPuy7QYcXAy4FtZ+vf468i+PcAA4whPHMBP8Upc7/sc0APak7PTto03g+
utodoiP8On+8/IJJcPqZ7qVpMfwf/Wtk3Y099w1TP0l94p2uH3F1xU3965qqMHlhZCGYELNA/bjx
y5AxTmic839fzyV+T2rL6juxfcAG1XXEnZqd78ueypoKOKG20AnjExIBM6Uf6e02KrFGRQzOkvQl
NxaTnbuu6eVdKOnbkLZ7O0g82apwd4QDJftO1Avk4Gm9JmlWt6uWpjx38zKwi5iqssW+S1zNRfCQ
yH/+wEMCjKgolLsrs/59ISNePhznWgC+tp0t9U5cgKTtfj5a1nHAUHDbjts2HngCnigCU3SUWzss
dJvTtmb1v5mqW+kN3up4MS3d/nrTVb91ISQrs9tkWCsqtixIbdKLj5iuw1qShLgTdDp2GpZUtVtY
7kLAE5UZsP6qD+G9qDcywkb/V4Ycv0kmE1SAuaD40R1d4xM/ybuIqRoyqF6hK2QNH+cZMX9w9kBI
AUbjJ065swxQgbDQ+fOGY6Ds2NMYQbR0+oLMO1tAFbMuzVwrIhjxG82Cb4bMzSbVyPr3WdZJhMO/
oTJZCpf/2CLE2xqjHOMF6K5UDnJ1UHqsHyPufAbymOSfyxsbFL4YoyIYM0YZV3KEkI/LwHmrc1SR
/X2EFGUVYi8lnb4oFST5uYDXPmdrw4V88UQ9cqXWZ0rCGkQx9S1QrVSle0y8JDz4VJ+wGs/gWDYw
8vl3B9+APkeKu9rCr/yuKQi3lm3afv09NrtAv2TnpoAP1969tJss6VJgX5UiVMPE7iyQgGD4h9Oi
+Acp1FBHDdBKUq5EneA5eGO9smWHbxFiHCLXda+mxRSPTiotMY+GnrnmSMjoMoZNAOKZc2dwk6+B
oKRvMlPWXzqWyk95dMz3Pl8ybnGAZCNo1zh7aCPQwqEzK9Uuf21bg9xZBYWP+BwiWRDj9LBXdATx
vY+AJeTpYcJvqhqfYkslWQVr6TaCRYYRAsc6heBOjP53heyY08scGaRxUfqE51SNEaWyxFUaeCNu
tvUeNrU/KCyK7K1NR1EtWXe7zdUhH49Ucd1MQyRK17qqZjOV45l53RruCj4qbxHl0yBMgdeY9auV
FqY989oWIFufZ+TV2jxJ5Dq9qMw/8czmmaXI7vOn1Md27SvsALVp3ZHWFPw063PkE97gMNjIqwST
mxtlGIeKbd+WqeaqknySw9Ejrh8698q/k4J2HV5FJrj/Q9Enl3MsAIeFcfnmZRWn6Ml/Vu/vcDOg
KJ58Z86PrqQTe071ltqiY0XG6UfOmLo1hWzg4Er/8YVb6otwMATOMlc5SYstJSH31W57fRMVDWOW
oDdeLYDQyb/C/om9gLc2GjGd6PklzRHBre8C/xrX08VHsDm8W5A6+S7OWoJTljg3faDou1Ae12Ck
gKuj3hC1P1mV2biezAO/5rl7+ujTmYHiVOeR2KrvMTlgxUxhwJsdkQCc8+uuS6hLKkfoXiNX9dUJ
zAREASC+Ki06rkXqYyrmcrXYLR+njGOVYxv6KATFk6ym6PnAqgPEE4bpAuRkozx739C8kEUYzHYs
3684QcAygG/wSxQ+w2OtYpzgD7dECyB1F07SLIdxJBDy5mgDCsVJfi7xJ3FWAg8xPra12D4YCgm+
0Vzw9DWQL5GdRMXiIDwpvmke5gJB1d3wuoavEU0SZ6FWKT3utzR+bdz6iNnYaggyThIWKa3dtGHp
J4/o5+UDaKSsj7kYuGZx9xPitRWeSQiMGOpim/OIpj9vjvvdUcANsYxlHsermB/ZWVRYKbzdCNsl
S948WppeW2XwD7MJfP4pm3P1lGYFkq8YSQhZ0OCw92HgTvQex/sq1IgFfiOc9Iz573D4HCwfuWpF
Y+m8hxSbtlvJcLSkfEeUK8emmFoRSg0sGdLpROF900PUoGEZLQe4OCaBQDNPnMfVvccJ+xHewIlU
eq/izkykQDT3uGRPptyeKBqAyHkLUEcZzxo/rIwOd9KGwlcb9W27XSNa/hKTrxPkAgftiAHPjExW
UHRtPpRPzwdvBRzmcH0FtIz3mbH2SutyCSIyv+yMZ/Tr4bMxiWnOmYvLFWyniKEAXOjT21Y9luy6
ednqebxU7sYA5lKLIN+m55wygbydbOzDArQiZ5WRsOcsMLdXRpKIIUbN7YEfrrEJuWfzrLevqVAe
fKrVGEEbK4VEaw7EljqfT35uPfIVFgxjzpmYaSDlnJtOKQkdpwBPCKi/lMOk9H6DgBwkLZyEc4SW
HspTbfg1yQP+uQStb/qRqm0HHmMn2/zIuko57alnvjwbTKnRUzoPUhJBtqXUgSSCaYMZID/unSBr
BVFGNITu2pTf41vvgZePBr+1x6xbldRgX0M54t3NwhTLT+VSTIz9GLM/PTI9wriCvOxqcWhpyeOM
vv6f1ohVsmqMMu/hSTuK2i3fOKBbavEkbKeArtivezXls1HGa4xVdruwtV2GQjAyDIVV6i9SJoc0
Wd1HFKwOIQIw12U+g2BUujC8BPZYTbfvNwCyibYl3gc5cutNvqXo2Ng5BrKkb8JWZndGw/L+q4IV
0mGs3vaGCoWnWve3z1l4a26u+CG5LQGbSNNO63aANyAkX1dolWvgqjs7TXCZi4CLyhkaf421SJzC
HhiA3wTa4a0LajMOfExoSUi+oW3ptGFWaVtlo0XbKxremDmXRXpwtyp6JmZjTmfToKHn+p7sREzP
JBXtWPIi9cmWD2AjAPdyahrxR+hgn2IV492fw6uNvkaHoqsrghxVoskP11pw2gpRFb/zB6QFqLDT
Z9ykVz6pdFKQNHaAZIhMHljVmQnDZ3sKUSmw14cvb1SSRHcblgiVkNwSKXK2tELuA3ibGOhsZXeo
3lhMA+eIdIVbZ/FqErW/ZSvv2IaV5t3ciQXBpvx40uwWxrpadxHIapnHilgmEAuuoDaiuOHY4T62
gVLhPhEXMDIidF1PoNpYWIHvTgEIR35l6sTps7tdgghJBzS/f1lZDUxQPZ0FALiFQTpFDPvbWmLR
ZQ9xF7qSyGjUM12igowPlDfA5pH1KnFNf2KNtRywSFpNDecPcQAqB4RZyK4P+UmNvdApKUsOYabu
cQ8e4d0d5DX3tt0QgUHPFvxYfCReGQgG6sd7e1H8klxjdOVsB2zLBLn1O6fq7kL8BgtFiaVeURab
67cbi8L2YVRK9y1mWOAO+9FjP/sxDKhC+OnoBKwDc5/3vpmTYt5TH2iN+AHenWAIEIQer1zMBhwV
ZITawwRPCE6ZocbU/o6DqPO+XAwJLa/R3KCJiOMEjHtZKZqI7PRolYgDVajws7/iwVBKqB46JO1Y
bnvxy4ePISq+L3A44AxMAAzofUtCe3yldsvqT4CR2uxCvSETMDVAzSoGCc9vmtp5+9x/63IcFq1U
52vNZFsgvDTsS5UcZ58Z51UoDbUp08svTlMv5P9VTuIao1cjdGCt1X7wssjOH6oZOsmACzh6PtuN
4IFPIp4/vIoLaRWr7eGJ416gQzbizln1v7akG7V8/b/bHk+y+V6iGWxqNNGu5ln75bT0OmUoSAcc
csEWTPGyUNtorUuUSGqizEAQ1mOM3BHgK49/uEg+syxxlyn70HCYyllt4RX/KyQx3FrkzuGUukIc
trU+k1Y+dvcPzMSu31axgeLyHHOT5Zc0GhC27y5aCy4xIXPqMYJgLXb2GvayhbNi6CJAfPgh1m7D
Qe97MCrgehYWGzikl3K97UYKDkfIiHBW+chFBZS97oL/BSC+AslbfLVYS9DmORpvhhqJeWHYSwZ1
OOvKB1J1xrsAJ4K7UlaWzZMAksfPk+Yet+Avk/4cEadWTWI9ABOFLIXlnlzlT0+SJH91vVYeDNl4
b3mjjMTIcHcrBa6NYMeNnzrhlNlKU01i32Q/+ERN7QHVkh7xzm5sEkhK9OT5o37SfqYr1JEomVi7
ORcvBZ/Y1IWaq8WHhKnggDA/ovAy9FBAE8r/HgpB+TCmnaqXBxxAkcjjD5QPC2mUm++TUf1fdUS+
5EQiT7ahvDgogTMibSEf66AAyaLTYsOjqfGfJFg6vYRqCiaVhIjPrHht5s9qB/HnfGh4KA7TbFmb
o/XGgks/IJmxg9hYSQBufbpHGvRxVRFiEC3W1O4uW6v/0wpP38BpWR2tsYF8KgVt9tbBchNVTqSK
ICfar/B63JNbU0XzzB9waxA9a1ggGWgdq8yXEaPfFUpYFYTDhsvx2C6tHyX5Mr3XQk1SkXAxau9O
nZUpOck0PJc1pi5ttdAxg6hvPvG34OJ0smGQ5t3as/hl4FRj3OL3luD/DcxwLjbevhCvL5YhyDha
iDKGVhpqdcdLy8cAfNDRo/lP4B8OhTcsJoeLlylA36vmq6hrC6iq4N52RPzaLRfuF3vn7tF0Q5NO
cKvLQ6i4JfZrrhDSU3IOuO+A5xHc2RH2xm4JECIa2jCe7c/2xlT4p5qNMBux3G8wMmXza+pkttLK
ipx/e+mqSqAFUt8KOlJyHM2k4VFN5i+lD2zg2GK6cZ2t0XxE7w3Tn+5SYCY2hVN+isEXLM+3shrQ
7JAhtYBVLC7mhYqA/EcXD+/zF21uwJufZy4om1ucg8IeaG4OmtbeIqFrejL4Nvrjb0MmZt0F5hgi
DpeKv8Mu442PxHfajXvpFJ3rAJVvFeuqjJMZE3rfn90XPA2fRnSzGVoZb5IxBuIlUHjhYVKk0BDo
ZaWhUGSUapkCfXOGsEeQuiJhO8q8YAGXwZlwew3ZUdD96OdfhNMJNBwsxLpQCU0fKwhjZnZpAAdK
GgR1r0A51zVOiwYHoMg33rk3yHALXQLlNh46QPyftZbEi24iabM3ns3b8VtZkSa8YTJnKF+3GvWM
Nq7bZ3vlL0yD0axBFgw3CL8IRXPJJIZ+YcWtNuFY+bbROrxDcnTdCBZF+nBJ5Mqzq4qDGDKqCcCx
knd5i7g85VPfMHj91HsUDOBwFjh0YNQC1Gkmffhd2qOaDfvCe/fLuftwfKCtViRaFc2vW5fhgjWq
9dY50B165TYozGYl/0fGeY+TQZuFo6JSvdwNFYCd7urpIPdRYo7qt7SBtoZMb44vxv2Jl9kxs9RD
7IzQLOyPOgYFRgON6j09kyEl0vN6X7fzOgWqMzUds6tYOjesrqNOSrXoknPZrDEq0J+YRo+GCZRj
tVIgC6n7RzWCFgqzYJed5oJczdwWrd6HY9mNo/buitJ50zePHv/6n+DdLsAHKC/QPLNQkAjoZpQk
++vc1eTR1l+vEqXK0x0qW4pbCkxWQ54MHh+ufn2BFlF3y2u0G/gwfB1H4pUlJyvpNTnfKTgVOaXk
LdaiOJdVvSDWTSPLhlywLFDcfsOG3SzgOlWfbdOoWZTZ8x/9dZ9EVaF5bP5XEVJY7rrYyPzq+yrI
8G7oCxFcqPxL0qvEGwSjCn9C2IIrXvnRW1EId1QUbPEOHNbktpV8HVfMhsUzb+wGL6OGd+W5UpMH
FBli2yfUzAWhVX1z3sVlE9wweuTU3/TRlMHAXSPX8fIEEsTLTXEfyhHTUZYb/5rcNP0CVp5k/kmw
41ps7PqUGZE6Ggo0Cvxn9vC5YH4TkeAX/HVTz16RRVaB9yy2UcJQYoy8PqX5tLEY+pWtiMTxy4LF
MVnmt9LCpwASH08As6oAuMdbP8R2phPj4+0I9XjH7T6hYh7v3D1G645xwZL2PkXKbVF80MLSIOjV
JTU9va7Fa2/WX6HKcMns+vX6SIj6eL7cw2jIa2AFrcpOLQVlAjby+pZCCvX1/hJHzDNslHtAuI/8
wX5NeWzWB4S+WVanITN7ay8WPx3YI9RoN4u35ubGjLC77fzSwr/i7b4enLC53MJAUIl4+9GOMHgk
tXaZIacy0FQtKUYtsnyFSryqDVI2SzjtnnAX+PUDovKRoa3M11ddsy5nq8Skri16bW2Q02tVBQ/s
nqIBOMVJ9ZXMYebwkv0y7LPk6k63N8e1uohVYism4t+6GaKp7GRYWhHsSpmgVn0XQ5b+oBGg/p63
c+jHNSZcpnrpzKoWVTf55Qt+p0irmxLxJYAbkoiFACgoc03sta37cM99/IUKxPojnYnBmD9/6VRS
LMzXouGaIVgq/XQwsqPLN7Uf/jovvR19FMg4fMhl0QN3/GRCyAaAz6XZEm6LST7ObiHhL88oLO0P
Dcj0gA/kvlludtUVVsLfqBFeqVtOittEEcoeTFFoFlNY/X6j2WLyBm81RvmmLj4E6ZYs8MSoIjGw
mVrJHkgYRzbUOM+hUn21o/qtCs6Mj7Hm5tBhUG/w56OtBfDEt/qjNl1y8rgX17ccRmvyqgpKblRj
ZgmdFpzfoflQTxLxfwTasFKgRsF2gcdOcnsFdXhWQT66U5G8Jxy49HtT/5+GokpWSWmix4AiNcdE
fbDqZNSGj/AX2/bOnf2KQ1uSIVFUFRoPiJz/HWeypVi+1ncNSG7z/mcZtL+rPtc6Nh2R9RlA59VB
mxYsSblB4B63I4M1uLkiynkIU0j2HitC9JIcC4DHX/lsZukIqfilUua9tyWXnd31uxmU1NkZ4bsi
UByCgJ+mDZEVVz7n0cCGXwTmA53NohGZu6Zin4cXiki3E7Y6+9wuAzAl/Tv/PMm1HLSeQtzFtmEB
/k5sox0TYNXN/Sv//6abE4faVwQJ2/MzBx6fEWJ1yYXSQAigp+6MXIm8aMBAKRwvLbYo6se5hNFF
2Jj67xDO3brxQ8JXC5ltV+okYE2OyCs49g4uairjxx6aKdqmKfxh0dYiWsr5NeXdRkXIS3/425Xj
CeDEFRYvZQrErykUajGE6Sk/QND79DDqaFW4GSGQ7xjPduELj5BiK0oJJpoWq4gIMkdfPU/C9GqX
XdH6v7T2WtprsnSWYwLlrR18yEsWweBXRs04xkEoR0yQhjx/8bl3/rXcazwE12RFqmO58pktQQP4
eg4YbESaR+jm8ZAAWKVTyFOPICWYkK3A8J1NbShOqIAByIaaN/FR0jJ6GI81e1pPg59manJxD+OD
/jYbk0dHKlWWKyxZgrngfrHeiECy3X1LkTCtI9uHeZBIAkR6Kx7ZMPSRHVYc/bHVbP1kmG6mNoLL
i8fnf2YrrWgXaw9kpOSbT3vS2zLkrMYl7da8AOWkuM8U2XVUbOFZGGGXlPUepQ5RJh2yTBFT2uTO
Ldib56H9QV6A8M7+1h/BdfeI2fk1/3isR2m/PP6pALiXFr6xpnAVYCCsHDbBvAblH6SomIFZdIZw
UjV3kFzWZD/gFiRICyQ3apo84vqhhSMhxQsTg4fZbRryzpibaAAz8VBweCNcVN+oLPgS8ruUvnFW
xtK/heb8KURFMkUlfEW7qLe5OG4gROBAW4ZZZiYVB9mg+1jbv2HeR4I46EeihECW1720Axh1pNPB
uQ+Og9njjlgwAvpdIjKGMjHWCMrato+l2HqhwZimjeqb2gE293qWfSxc16Q814+orKRK1i1ymTX2
9CxRJ4zqgn9VYFrKSKjdKgW9agOZwQF9R+/OF6tpKuS9ULvKpQJ81f5N76HPlMKvSEN8nXeEC9BP
RrWIJqOJvEzlNwp+l8EagmUDx3U89Qo5K7b5VyTfKbW6IsYA0bmL+My+qViot9IXb5NLeV/oEnMu
GosipZHA+XJqLTEHQtMQOrwIHlV9Q5u4GtfLDR/jvaddrzssqoPVRIW06xorQOkCq5/CLLvxfvFI
oGALMavSbBVxqsq15HE1S5qQquVtUnosKCWHdjvz6u6eiBWdyEStaG5r7Dusj6CDaU+ewBMBdKHz
QFXboMxiG1sxoNNzOUftz4rokImgyZxPtl85svQ/FShjX8DGyClLfqOw9Y/BI3OzJHLsgL+0h1zw
/gHPXrLDZrHdrdEt/hqmCI+/CekNyBxRMUVwuhVw37Kg6uvPjHfhRVgLUavIHt4WFyl9hIW3XlNF
1Pv6UacZAjyP5TbkWlq+KcE69Ros/0LyU/s0AL/WBMVvnBY6j7sgXMdh/yIZrBk7efd+nvAWZALl
qa3NXuVCb3AwCJcDD9+Qnv9t/jeZGap8hkwXxVYPiFBBDJlaT+lUN2nPrKdf9Xbnfdln9GDHCXvV
F126XEQgPDvBkOVzq6Wutkvna+7UX88l3lgliuZand+O2vMBPJujupbz4yIWhaKts3d4yCz6k5T5
TmzJR6jFb/E+IC1XUk4jW1Csnxz0FnwfbVA1fOtPi7JMRQVk53jPHK+kIAhxCWVW8m2KtYKJ90lO
kG4/c7YDza/ys9gr5vBLaAdUKPh7SgdZMYh2JN47c7W1HffCyQ9G1oD+doGNpgza7dz0xtG2+UyP
Yw8oTVME9Ml9ZqMpZ85klN4tFpIQOsvq9OHUglzgPmXzF0Gw957OBFYjj1FJMsFRk452IDwMAddu
mZ7LFHPqlzzyMwFxEIBMQQao3S83hC3x3xiH8ZKaFdTYPdZCnEtPQLmpTqs+vIhGm8o72RA7mufG
/CHMXq4q5rWWwmabQUHTl0FQJjaPJpJU+gamLtm/lEAow1B0wMJO/WzZTAfYLY7MkepZ0fJFFfdJ
a4y24jLr1R0Na1sf5nzIhUkWTs0ue59sPLrWRl0oBmlUYWEANgM4MYjCKjS9je607lMsYvMEEZ++
0k6SQfgf78DLguGsRcIdp69LDTCpnTOy+OMDpyAEgavw/SP6mTH7HhfNhArZolwubx9yWOLU+Xel
uHx0+2OOAliY6kAvSUO5eWdGLLYXblHFoi+4B3h7Il+GYNLoxS1c1xSSNXgqMdJgMZF88Z5gv8IC
yXUafqEKnfqn9LmlXS0MgQEw74a68OSqIZ6jUY7DQ6DiU2QgL2P09hAlVWKQmJFAkQOztIncwKFm
FFaDfEAsz2jd5vh7jUg0KI0CW2WElo2hxlCSgbi8h1HustZOSUeknFhtIDJdLy0SWiiKD3cKlqz2
TI0AqvJBxRnSZxVa1SQ93uQuE56TEVrK8GGzk8Gg5LA00TOlJ1Ag4b9qr81PzTzpbzDrprAJzXuh
00JToND1HCvJJ1rjb7ZtDObSzEzBmejcq3Q8hdgBiDr1S0O/UWAHLT+qUM1YdAeRHHoziz87jEck
kd+B68a/Dpj9AtPBpDtwpM7YHdZjOzflVnHxu2O9JMnBud5PejyQVZ9ShjOf6TBZr6Hu8W487JSz
DPCMOFX5iNJCP5MsjCFrJiaR4l9vnYlMEEMMe1A3zlbgDs1gcZN5BaYklrTL4BtTh5nbXoludGSl
uvOhUj1XTEU3om5rjaA+kZbJ2D/JzTY7KRbKyDX5+5ltAOfQ7+9sYsYtGczUJVwAKaV6nNMB+24O
LCKFDnFbcY9H4xLDs4SixNqBgXHYwwe3D9OHImJCXe1jKOT1ShT4UAR9lyUW3+dpS8HTDaxfqw70
MxFsb4/XfXbJpUCuGfAIMeS+YViQZTczvz6iH/P4dzDTZ3uJKBaTRHRm/601UbXocVdEGFUfi+md
cRHH9HMP8C8mkcK63sYfgSfRK3LhH2b3yqGNv3lnCG612Q3516chan4UIdycW+mbc5jzdjM55qHH
EDBD/YVL7cVoY7iQHHgMjp9E6lb84BLst8+/kzjIqhet7c8w8iSjwdLx9Jmci8W5S0iAN1AOWid9
f8oACm6xInR6+L9nULIj+YZN+hxCBLVh2+V8+3fR0kPGWoY92XzG1x6q8HkTDOelqTHt/Hxo60rg
4JF2iQbJnoaXih8mWT27KDlpMh9NC+H4uunHp2oCyZhNXBiwpjqtldlzg7ksApfUS9f6moQ/Hs+5
WcZ09OJDxJB0hw0EhtYHESN08a802WGj97rY3OIo1cKxWkBSg7zB1rh78YyPZmj4KlAvPdzEosC/
8WXsYixkIYiu5QP1c6TnRgWXkI7taNMKt73N7mzJ4rMCVVjukETgNSJXNnuK7Y6MLOwb9ZzeVG6X
swzKzEf+FmWVM8rRn6isXuZlTpEXrMKMAeXM5D6/LYPracPGFPfGH8oqfCVPE22BsUJt//f9xjch
QzhDQIj6PMj7aQQELCQl918cElZIWwKEephJSt2xILKDYyFXCu0AaFO/TseNFrr9ASl6LETWDKk+
nE/HqAN5GFVI1Dp6Ujuc/JL5lUHgxec/Rp1deVM+NogM8hsNzMc8rWhYvS+a2njPFFsAZXClaoyj
hlQ4y/bMyTiU+tk85SFo4N/ieUiwY9ghMaralGwY8vrIFvYOM2LyI27c4nfxQcp+znaYr3yw3Bhd
wEYIGEcDL99WxZg0/cjw0+OsarlbgHe2Y6V9w5Opl84gmcDEv1c3RJCkRiac+VToi6zWl1oIt4k8
Olb0O6gXrD8HcfC4PydAzztXzeHBqXMUoyiG3Xq1LHWKMxSkYxCdM2NNMSUL2X6jwX9cWy6KTJkm
OkK1JqgeR1kbck5gPMG1zDjCG4ZFXZhjW9YAVCRm41v0/7AjmSmkGm2TrxOk0wYHW4pd6kw5m20n
cXCRI15wwvAQ2zWP3Mr222BcWUjFbmATXI0KqHnO+E76fJJXnppKhb5VBv97OOzyfOjj6mNF7ytW
U2n7txsO1DnvljzQFCcs1Pgu/fd9eQmjnST1SF2pD7VTi1R/yNem6jBbutHHYN1fXf1HZVyQDk9S
Rp+IKXIhmFBG7KWN4CH1MftjCzNfiyVlPuKPlj8pDGJhAYd51BzijHUQ9e0Ntn2CwFGwZ1EqDfsp
XNS6bi/8ydhhWCFUFTck8dbXw7xvH6uBBGJoz5A+eFUa+LpwBOFA4US9QBwUxrnfidFSWgpaF8qd
8IHr9MAe8vU5yUJdbpRjb6wmrztHdp+C6iYzaakKoGTxuoW5jwZtpxoHm0FDMZ87TppMHbuHnE8J
h0qbSdne/0n7hyZ6K7+DB3sB/7OPQYx+iFuFNmO42jj17zsrUFsfvi+PfY/U9dhBDerAnJlRKpuJ
t1Cj3d6fLfV8D2OUnQCIViUQbbdd1bcG74Z9WEd5HQ9SSPhGuckvdbzOYA0qG+KsMj6cMTXG9i6m
wDjfa6n2FxoznKbXeidupQ+M1UkBhSgRpu8SLmdUfQFCHZoWCVgEMY7NTxJQ2i0Xu1K+om7CmAcj
r54btgpHpROhaHAiYbLvbkjv4gFF0g3/KlS4aJutcq7GUYTqFUPwwxW/c8ghoDSzuFY9ZFJEtw97
W2V5yZuYvaa4xvlNA7M+IkVjXOcI6Qnp4YAFfdD4guiphiGXz9NSzjMpiQeLuO5alcr6HqPGZ58Y
Z0udP3CBwJtro4BcAavzpj+f+Y5PlNtZ497Ui/hmCbHGLIqUJ7eM6+fAuN3wwnmYM3w7GS9ruHIy
uii0+lG+e74hvWWkMuiDYDui58m9cE26J1xGQ4lVjQfwYl+j/FPCn6kByXHLO0k7Z0J4BON9FnTv
IxPWi69TfX7xMJu92VuUO7eFR5lhy4LCtn0YQ10S7X2Khp0w18WCPU+1oFBy0JpuFG09BAexQOsJ
cg3PZMc7JuPFm+yMj0rxqKAuReDi+SW/4f2aDCVIyDyv0gdgWVw3T+/4UhMRgfqxLGLMU5crzHyG
KmBPvcZjkgdsigmilXGX2NiQC+K1B4sRoV4LK1EIJiTXz4HTIzGrZl22ZHflEpcsuSLH9WH1XO44
Eq+QvI4VFFUPwd2R7AdAv+4hhcgM9WRpC/CEd2nmIAQvrIGFZzwnShLwGGXBHjSO8FEP87GiDIvH
xCLGMOqqcORufHtlVmQmBi2NgIaG7648whJJpSkyY7f1atx0BdCB4e3CoVTx5uDbzHhX9TnVtBSF
YUU23mQt8lPlaGwlfap+/fe4BlSnBVT0ritB5Zxsn2zQdFg3keozB/gxBsxoW15qwu9phLqNcjBx
sG1O0VwlPJlQvx5B59Q1mEgThI/l4ITnI9CH8daSO/+39o7pDgXfY+c6wwyBLlRL4Cdo37PP/f8K
RtiZ6S1mD1HbANpzLFSQp9aH18C17o4aTdNpDSX0FxPkgbAV5s1p/B16sh9SEJgcyDfqauIEOJML
myyGRu/KatUcLXVKDfmR5vOUA246or811StZ7QrRYNVZwiPizNn0HhwoDkhag/uL//ISo3Mam9lb
4D4OvR8ueRHbF5yIDPU6J58/yfjR+h87hKjDIiNMoSVfXqGK70htw8VAMhOoFqSg8HlrGJtlznBP
subBzFKj8YpRw3dKiu6F6jS8wuV7+lN2lD5OvF/ajLha2HoxhndB5qQl+qE4bF4+ov1R25unFYnR
STruX8HDsFYSRD5gzSuMUuwdLnl6rrhTS06UsjnUbVlse1jeNZpRrozwescJDkwmOx0Pxzn1vcqy
2sN8chacNjXT/G+2CFU8lEnngphlfHRms9arsIs+1ACJwXFvocZBPpoRYU7sNWK2HcB2csbxUxvk
BXpkpg0IxRRRgmoCoOPG5YdwABSsGOGqVXS3KmdMvuLSFKgoM5zZyvm3u+tSW0nxxixNlaT84AoU
GLNlt7ImEhWv1iXZk/Dau3mAdQJexLQF/pNFRDXqUqjVcfPPZGbY8i8Hpn1fGteDAO6hh8ycGtt/
cMqtmf+dgvZh73D4cnFRztc6U7pCP4uXM4o8uSk6jiU6rnluT/jk2jtXX+UPI5kFoW5058qntpUX
pKf/7yrJWfGyj9DwxkBaprFJz9NQrVuzCWOLCGrcisudGza7z5IA2cbEGH+VrgjUNPaSejYcIvPL
83Jtwcvy+xoINZNcbhQwNImWz+qiAQ44wedco3scpThWdq3zb78emvFK0U5vdaDiFU3HIbqdhuXg
nbWsqolbWNnEDcnU3HPWHniUAEzSo8oUp+HQD8DmXRX9Ys509wYDKRE9X0qG3faTZuzW7f6eXvnn
T7sT9Yy+IZzTVzNzJ/nBP9mpjkubDsfgifC42cUbjgl6gaKVV4718weFHNAg9tfByuwKy5OBdozw
WBeWIQkSAAQcP21sGy42nALKlMVsIFuJQ9tiHXDLkvzm5L4tw9hwqKa/PNZ8ANj9riCftWzyUQcg
Pcd4zHJTBIdyZu5hbpF9ZbcCPZf8W1aplvxgmxsaSE2o+ZkUVeh3vsHuiautczAW7dmBq8xyUT+k
Sx8QulB1n5ET/NJPrUYQpmFwcBNcywFqWdclQoXtihN7NHmvnAaMrzx/2hLcV0UDQn0D0r+ZISMJ
2ji+kxIqUILLl+a2yby9eXAhdPffhxj9QDdRJ8mIauAxip7hg0iN3D0yLmcn6RsWB+iy41hMSBvV
BE1ptm+AIBJItyPgFNAVdE874cjqpmTyQAOnsyuXmf36ksiB0O2x/ETY8iMxOyHPHGgumB2kyZ8o
BnQzJVirwotbJJMTCTM6mafTOxfQYHfKtz8+O07/co5X67ARuB28ivNKLnMQb24zd9SnXHXn8mwf
ao5+FLC9mAx9DJAwxod9SL+lcFBR1hrTdNM13oYFBbKWbo5jtya4QW1iuG7jfpdMaQeqowPdUjSc
ad8d26SjxXn3digfReokn+ehfv4uJC/YsOR2sfUyKtfRAlQLWX7/ESzXwN1uvMpcJKGA7YGgvsb7
JFz8hzjQoJi/ZESakofalFQ0RfaVPskXZb55aXt81smhGhUkJ3WYHkyOc2nKuOqMDcNJQu3i5Dor
fV7RD//mTxllNlegNzkPWr+eHSJK0jxgQqDPThe9FodxD24owpaw7AL+Crg7BLire6uNYTNshJU5
Tp5SRHzzz4mhSi6dldnkTfnBStY9nzQKQ6LQNFTVQm7LAtZXAcjLXDL9ulm2Bz3m/THhhXZ56now
fWfvMon/qhf836azcc7J2SpThZ94goSYOiC01jlD1P2A9kaCoCcCg4ZfPOTWZC9r6mUHdAqfRAwp
sBqSlaKM9fuMPvF8J2V51uZIh518woTDhsiIS2Xytivav1vKOcMxvZ9PVqhpGjN9JGDhgooSjitk
pHI5AwRnoziXG8VgdpD/Xsh8Luv+rbo80wwGJ2Y2Xm4ugr+Jic8WjyS8wvCEKUjEyn5u/t3HfRc+
i7u9fd5B5MuHM4LJqhzAgqX4j6FLPe6FEQoHqs+hJDbLt0VuNMfsGkbJg6qSaB6UC3IJc1F6e6dZ
yfiQwxINnbSbQsl2mx259aUuFtyyHLyb7cTpsZp80cJoU0GNlIOiiT3unDw4BYPjiRLy9TLOEz1+
rbZ7r6917hzhc7qkBteitKtMMt1HI+18DRSWXrje4TmtaJEbqBHs5O7MjUCB8gGPGGfybpp7Fgo9
NNO1eH/FsaCZf9kgRmkjIbNOnqGJoRV+WIeW7Klcj7rJ8NjMCSvIWGiU/qeS2GhBgGhBa/JoXvDP
diDXPOQzoaVC8dLKzCPAbND1lQrsXBI42dgcDdydDylzhuMMMbqozUsqKUfLPk+bmZM/ZysIZtuS
GwG7Awqa94ItyDFp2f6FvFv97BghIryGB04G1eqv34OJbCuKPP2HO8TBSG7/PBIgeCLVIC8/1Ys+
dkxSGDM7o+ka+E6eb3pYj8qehJGyupuZmRu4X9jlaGA7JSUnTPZGNZhZHFZ9obLD593eazJVw+/r
wqtRcrUZW1rIW6JzRN5hB3LsKhEMahIqUcGcy0yDaWppPCgfN43wYHm99LP+L5a3Saa8n1fcnw1r
PB4eqWa/ugwXH17qh+JyfOyp33g5/YzqSzkZOU5AzaNRSLGDNRt5wrcWn0IVWnXA+TjOZHMHPy3X
xWcF1/Ogf0D4xYRXZ0GtqyV3Hc91D0Ma4Bp1+uZZU8RaCFB1cDLnQmsd6MINt88ce12GG1Cb7iid
3fxLnEOQ3Y3JxH1CH7gWj2adO1PIWP/FikYM/vdSSLCcwY2pu+U0agCwDo7MiYx2+MtQTSfkeD+t
0LrXY7cGD9+qxtDGwMZfEooglYHM+zUPfF1o+2xk+EC6qJ1atMNhkkdbO2YitLF+JyrMpoTgemP5
TwSJP6WUCPpPciaLyKeBSj80KxdbSfkLfZQM9EoZtEt24CYMPjVqTrBpftookmsxzUH+Qnt9ODQS
hOGVTurKGVZQKPdXW+75KAeSuPrWnenju7ovlsw8eyizttC0bWUN9keIMDpPL/uQiss1Wdm7M0LM
oT7verEFOflIPFBSppZUtXVyLcmrkiPzvBgCXcnR8qFnDsSZEr0fO3C+BdCfLen8SB0dymzunpnG
0ADSN033qySjajcQs/56bmeqnKM96D1V1uQB6rsOijLIE09MD2F+cIcy4FvdVS5i9l5NC929UAIp
3qxYJPKgsQdiY1hAzRs8B92BwEGgMunsf6Shox7eu6PoLdUhbZmvN0QPgLNTffJboRhWroImknsh
a8ivp3XG+cG4TiQebiS4yElbueW+DDU6IMvRCd2HaAAM3Jnp7Ov/D2R/ahQibwSnEbx2cQ7TRSJH
t437OcpJCBFO/02JAMf3URprUuCCXp2Spr01X/qVlSAf/gteCKNwL8TTxzpkP0uYrcpwjgS301tj
AMkyD7lGVaAeKvOmL0n7XFH5aK4BclaYQTQHH5oz1jpyWRQlg+0qaHbvalDieMScMtAj/fJbluSp
pjWHzXmJf/3jjPT5PF8VybGh0pmOcbBuRQXnbXQs4t0wb0AAmeOYbFf1U9VEVPC3TGgb6fZhcS7u
XgvIsY2GVj+TKWx/IuHsYCWn4yICsqwn682WstskFLjN3gGjJZOvbimtvVNnPqVQHg1XQiWjXBdp
mQYS3ztO2wLXpT4czEIBDVn7ZrKzI+MRv0owcP8+ac3moDCiH8ZGy+8kG/rJASwjKx2csZbPvsAl
qgjlUA50uINoEfTWjywOf39eJo1z6bfbwT71LcSTudIt8NfOUvXd1fAXFJMVGrVF1Sf7dSGKaJQW
RIAa6BNFFdEWapc+rOC5VXAWvikyvRNCmSbl1voE+fIW+kWSf+X8/WqZrZ6P+RFxNMj6nEUVISk7
NMGBMyHUzALblnXHGQoPH4PBDGlS0tgOB72QmfzpcV2IdX2D8CIPelC5W++x0fdcilLYLPrnTrl3
CR7SMl6eiFG2WBlIyfCoDjTCuZ4XfJghuk1KZT4uScBQPexczcsRn8+6yLOYyqSjPi3XUqIQhCAJ
J+4y+ii3CQE06cuC9VHlJROzLkAWWW52eJl4wS7AeCwC/dhDsuDNTamb6fYIu2lz2hrtP9KcOu+4
rW9ltjOS0X4GjPBKbrEQpia7ejgLgBBXx7Lle05i45XjDcoUqfwgIIJdFWFAClEN0dP2EnsWKC0+
/hd50l+nOyqoWeg9b3ekjkeu/dqn56ys4sV+krWvePeLM9CAUeh7LUZqoS6oddyIZCumSJ71KG+w
2DSS78Gd00NehTnbudw24GsDYNeKPVBHyxTsUl+K7ye2QC4Owi5u9Z1Gr4/LjjnTMPsC6xO3fQNV
62O65it8k7ByUpXbMca44QHmFnwbqf+c8jUQ9CsDFKTRfPosdSF088xTtYNZrilAMXC9pnAf+CBc
CZ84B+2PCUIMc6NK4jjwB/an2qqIM67yCMdvV2yEVSfdRqkEt5+yUTxACFTa7CwE22/UvAegJ2DX
mNFWvgL1bWx8I2jLwe00FVjAkD0hW7ojReaCNs/t06lp80cli48QxxHTmya3iM44jp5Kn/D7JR/U
ujiLL1JEJFWH7NOkNLGPyxyaK5esuoHm8rx5fllG/bIS8SSC0KkjsHzeKC2XrkYwSkVzQONjmL2I
5TbAy675xzL49CXG3NOO7oQkCYt+IixTbrcMMdhX1rGDQV4U0f4udTZkkp4kJXTBTe7BX8KfUlAu
VGcGCsfNm5+KedQyyfWHXY3tw0crMjBLtjX89yuaW2SSWtZIPAWrTB7NqgLP0ZxZzDoORrPveoQV
5rgpj1sXsqwu052vWXDqGkkJmECyXI5VyvczTDyz+nEXu4tyzlv8QdUXCaapIMtX6HwDcSn26jrn
0mpgae6vJxqT6PjyoKlD1/bMx0HyNuwgzvhyc3G0bao9SRE9nuXCJoPm7uPne++7n+S4SMp94PdU
Le101IYL7WnxvoRPhuVZOLBoL8vU4dZaxwp8hPY3zuI+1oFBBEhMLrnSpiFEh8CDJCvzEPiFSmYM
hBZI89aiOmebGqD6ki2iRoyGzkdphKSzGqlEqLDNZebivZcEQOoXoI7P3VEKyNDr+gqJ6AywP0wU
NziItpIcScMC8Zfuhh6/gi6JJhZBtXi8WRzWOvl9vZY91QT7TzaizzS/P2UVkTRFVGfpZ72GpcYY
pB0YXdlt2dzO2iezDUwsTNJNjRu1jXB8ohvx+Efmzk/mGf7dkCgYONofTPNmO7Hj+YHW5FMHs9oN
j1Qi5eDwlVf/gejh/BprEtDniRgkCV/W9CAC+iTOJayweXDFzmlBv3WFdtS5N6+dCOz2Izj4oVq8
Uip7uV3QowlDRWVivB2aiTGcI6LvDVv7P/RwFjjcrQEdU3ndpCAx3q8bnDM2ss6f4qPqu0KX5agE
dRx4bGT5F87zxVJk5hMSnY86QdENwMLgSIxMlah2LUynjq6Gm5MDwesnc8Mh+5ZoIV39xxNhazAW
LgMq2lQJEmiSDM46HItr4GMORMh3QqQDkdjvh9YAwzWLWRVkcmo+EedjzVtKZez/cL7Kp/5EgXJE
bVlapurRCX83VG+NHSztOaX3NXVZC5ZpvOUkzmXAHw2MRE7wSV6DOahKKIF54hsgWBwDfMN1W4Zb
1ybMy03xb26UCk2FdRHCHPULsq/Ee4lOOwhQL5fnqsELmiLd9+JaeafMAYjYPATESKtFGeTvT0F8
FRbBomAAEpft+WPymkxl5Zv8hI9BBJl+Up7TaBld7PEG9yLekCQIye91us4Lwu0KDJ2S/yb7eOYU
PhrnJR401QpKu4oV23X8QHAso7kizXM6cOX0Yx1ic5DMe06TNeIEwa3yofwXw80PexuFNyedpEMV
Wn1qw9/T9X2Q1FCRr/tjH2dp4+jBRdXm62A1/MDktYXtqPVk7JCkq4nhFsb9hrgEIOEgur1B5CT7
/vX64fW8vS5h6gsebGCQFMpv7NKLkaU0nSe058Kstj7OIC64yzIzjY6TcdiYsOcxOTVrJ7Bs/vIL
rYiIizK02Jv2gPvtlKQw3TACr9qswaF5xzeK30jqyXb1mLIS8Cs8DI0ybgrVTDMceTLV2PN2oa7f
dmNcHAx/LDUPijkf9PiNkcP8ajVvWZZDeI8YO3M6t5cN8PmUqUm8oo/nXj/0fM/PSkl6RWIWcMeW
U7YSgmV8UTNDPsQBxbnR4mxrw4KwEZ+2eY3JDSlj1t/gfAbVdC7AzucJsqwcBZoB4//uPQjTP7zy
Sbng1RF6aMlzBZQH85l1/DAQrEJ06LAycQKKBz8MyOcTnfdO4Lemk8VzxQM6KZHbTXpRUFA678Kg
fEHGZvdOfWzNwDzkGRyxaZZ/3Mo5x5AvQ6QqKF+dAQOgCyv2jiPI6XsB6/hqOy+uPlpefm9DZNjc
0uJVxYiyGs9KFXcajg7j44/e6yq5bLX1CwSWIBRJS6KBrqOAZOhvBQt+MgAbD3WKZyfqcHpWOP4A
4MfsitbAiaOGAm76C5RnxrbgHhgjm1qbtfcRhpXXPpvfVeRw0eWtEpCGzsyISF3bCnnHwnbh5UAu
d8h4T/VRAIh9xHGTIqw2tiNg4Jp8eneFEGrMdYXe363Q+R6mKF4zbRx3rUrEiudXiAs1hetOJQUv
IrvKBvb+aPwG8N4+bvfpNOtN5OnSNFPYkub1mTSg003KmHcttX3t1HJMBRar3ziObvdjMkBVkwPV
yg9xjiBx8CxmXb3E6XoG7VMq2/oQfNgICWm00gDvMhm07PVYP84nTxY04oDeAk15vhJRcYHZErYR
kUW9X7vMa91wADaOl5dEtZmhGK0QczEZL6A7XT5Qq3lTxEo0ixvfRgvVmON+vb9LaEUN1ul4keHr
aiRsQ0LY/adf0CRpoBUvF6dSLVPikY2JuL7h8UMV8gjSd8P5Br1sAYhbBxizwEIYxQRpn4Xcl35H
4Alks0nM7GlgDTbKEETyWii2IHySeyHTyD7RhW28e0gEXqcmX9q2obaU7T0xCbbye7pPinG+IW9b
vAfrSgBcSG7/s0JWqUNlNagp4mnI9wjWfhi+IsLT/q7SWK/Ku56hJU61gNGl9k4eW7DNLthFhvTH
UnH/UvGOH8qFgobbRHRU0/nCAi/FWIs7BfvSUaPpx3V6TmJvbVqBDW3Yqs42ZdMGB4bL/e8P9mLn
SH/ubIoCh3RwsFs1K/fGe8xnkUQe8hjbWqbNE626wWVgho3D52/GZK19SX0l4xqVVwYS/Q40ePfw
/ZTKZGMZNS85pitdTb+wekCsF8vf4XL5tdir8OPLWDF1twZZWX+KoBMZiLwlocefh+GLqPAij+ll
BaWToHi7xfZs9gB1lO42HmMjdZhjI9d0RXJfvviR5xoRcGc9T9aVGJQVXYpPpEfYlhjp8stpsbu+
gn+/5/saGRABKPOgEpUbEFUJkDzri69x/H0N18Kc1rir+zVXHdD0m/LIp2fa31cFki1W1IaTSMeF
gNGk8YH2+tvFzOtx29psIsdG74QMkQNYMHp4Mg87a18XkglNnnuZWOXfWrKXJe0xQ+ubzl9aZs2X
6jPmr+avfuhprQkLrIjVK4nhRrgx/VG+1GN8lP3cllKn7nHEGM5Uso9KoA6xOi4yTk6equMfV6Gj
CqYQg73YOKgHCeihzjenHAmOzG+9cyrGt+v0WNFxBdMsseoYkfWT3JBzFUuYuNpbWvxYyItkfcKb
9bBmzssL50LI03oug4zowAtY6ntAvSxnxggMNWAK0zvlCLpzfO8NFS72TBlgx5RRrlCfDRYBFqMp
YSfNkwbVSCJamDXUTiv51F9A2g4FPU6tmkzZtNVcjq4wQg7/sErcsjx+sPwWtahkrA2nr5aeZ+sE
Gb7QaCykE5l0wPYkWmgPKdHt1yzzj4QrRPjMVyIoq02Y5NhgDrVzyxuA0Rv7XbFg22x9BMGAsfq0
lF2l3ScPQyHQxqa5L9qzrySGuXXc6TTmBprpeviTcR+iIm79SLFwjRPtlrxpMOD5uYMfq7FKO5QN
1UAYiYUCrrH8HwwpOvWGsue8wuaO8r/dDXEnWhDklInXcUD7TOvytqj8BA2MW65PpMX6qrw6DKv+
7EHu2D46aZSaqhzm8QmL9G3ow+n6P9EakRoZb95KJYg/f7iOpYlOV5C6I7Mzkc99EqEZK2WBTCIx
+9F+38KEaC2oWRID85cP+IuAENXwrW2d769J7xa4isrDb4ZDvPdNc69uKcrYNd4sPZMdVhUZ1HCd
XJfsrzw6TSMUj0MCkzjBWkVuD3HL8cPmEL2J9Yum51szYxgYzn4AFJf1opafrmHCyKTaI2wOxYVy
5ww16+PxXFT0rVKZlRQOoHnIsC1JgH7ETIJngzGqrpvNrJG3xIje7CpjeOWPdXextSmRQWg8mMoU
B0FjaJoRtiQOv5bPdz/rqvmgyBAaOOdA4iH1EBjoYe+fG04kiLsgBFKfcHZgAfpcxEQMunscp8IE
NbNNzGmbmXYW+0S9cm4Djs874KY0oBuQTByvHJwefHzn/JjIdcPJBp8UzZh59ZRT8DoTSHbyUW19
oAQHrcLA/vWVY/SCpREC9gxpnTrzTrCtSRNjDfnr5YO7IctcwDqq9NBDgt6GWvXv/ei2xxn7MKDg
DSBpizYwGFL90ZtOeYUIPvWgXiFbum2EDyj6c6Fs/qcS0EAlOkZ34lqSZmKRJtwD64GslkymuHZO
BLJ6zUuNiok2lU07pamsCgjmgyHHpN0JX6LYfrt1B5s5mqb/FqXtwifulCRq0d94C/sPJjLJlCrv
rCszz6TbxvPJ/4bLhiGBcfS1RISULPBILn3re74RJgzEAPFBw5pyYD2bO6g5EEebiEJX/dtZH2qQ
8w13sQO16+mQuYYygHPVeubuaxAw+9aKh9sx1n8yG8q1rmV3UhEVcEy0oHefUtj447qhao8che7d
tjxP8S5a33C03WdMP20++WGo33GHdW43R+7nC9s+Tzvp+ztRGDgpDg+TY5PNn2GgE2k6oIkRS3qz
Zb3pmV4gU8dZ0/xTvE0gKuNmR5QOZZAVALNMmyrJG5Fc9H1Cp/jHW61O1V+XrSUpYxG4S1cpTDDO
0iTzaPZSWX9GHSstCNzscEUx6XzhN7Vw7DVe00rFdav3eiN6yGBHs79cRmCTKUUnFUaPr8KgGNvb
RIhcfdJ9Oyd/4BpUjFuRSfYbYcMxHxoT1adtmUDiWnK0YinGE1V9DuGzyVFMOR3G3d1jSz6uAgNW
lo7WCIVcBJqpk9tzh2qO3OKnOG+hL9uxxlY+fNN6VMQjP0POihPhAxneT6ioC4mPJtG8Bujn41UY
AGEY/QdWti8XxO2a/hDJfSvpB/WFBuZ/8XQws3/3Xvb+1l13IVyIoFd8fVsCJCQo9HhACepgeqEM
f0QLfsTw2nNBFPcXCuMWYXf+LYLPr9n5G/322QxkrS5zkEm6fruuUNDVj0hH+sbsTec4NPuOgmPe
r5utyl3nwWivKqm1u2Xo+gNOFVLtxiQMqym2j4eGFcesFogthiRCFAp1ez4jNNtC9l2kIrVhgTdO
budRvJ7Yuk7eaR2DekoXH0uBvmvaPz+t3XESAzJ+GZ1AaFdAmdvMrhoeew51LI1EgTxEyfu99RUS
ztqz3198BRVN5GuAcLII+ONaaLwjZ3/U9Oe24FiwVW0NlHTZo3fBhszdzKM/RyBhn8FnztLXuHIv
HOfiYuGxbiauT83CG3QBcbQIptaqPYk5jn7wv8LT0E3QdWa50k/U2lZRLRG9LON1WO9RZIV787N5
uqdSCQ+OwV2gXn7CXjPdM/VFydOzm+Gw4gZP3k9FvAu5v6eobPOZi+4/U3rV2jyHeAIqdJK5/w4V
2XV6cspU2uScIe/B+wR+MGMt/jLktjYmuTnvFUNFOnwCERNKn1PkXLZs7EKas5tGRLwDudiIVtFL
r+ga7ZM2/x+MPTW2OuAI+E+k1sHl33oSlXWYtarhQNJe9ZXpIsNzOKIUpX9wSyGPQmlAOFS/GotE
2fN7HnFNSsMSrAiy++fbKlLasLm021XUAlB26ZDWVkYQ85CZ5H3lhqa6kv1vOQjJ8rXc6JFhgMO2
O8kGOyomzV4Sbyu5rIbCNCkB0+UBD6IQaAFX9l9q+jWlIPSVm6ljiYLXDdhat2feD6I3UdfoosoP
Ztuqr0lrbtdVimQjHGoBTP4YqjRFJ7mtwpRFuMx/njJjCKXeLnLFUtMh21TIYLffYI5aTX5JbujI
ilGddw9W1DO6qDKsxNPbYw2dgsrtYUcZUbHqmGzpcnSNgaJD/GC3VWGUoE7S20JsG45z2B5/rSkr
3z5gDm7ykLe4DbhXUKY0Z/++inKbHXv6krOFsK7oy3UEH9IOc1D/8TRyxqx0dLfNZpvzHL1xC76K
6HhVn3b45jKnXFk0NUxENy21wUK5J8M9WUGsb+QQWviCNoJ4J2XOgTSEwIshnB5TO0WYqMCLAmMm
aD/rvai9+53Mi0RpydVxor3gHN6WQh2arwSIOJFy9Bnf7fI+K7mOgENcviHFWdBGVmSZixZVn3u/
ItFXkxVQW/yQ52kvplUiwVluG9kuR1xzg6DNxNRAyydvhrnzoeCDnnXMb/4J9cWJkYjgSPs/FT1P
cVDxCwffRMURUeTyN35nN45Ptsaa/H+PgxVm9i3HhwWZe3AFYqgc/bwc9d+5ACHvj9AIEII7XPiD
y8l0SnFQBjBw+UL5tkTOgDEjI5TV16A6UsvSV0RX8MCgkG8yrZd6Oi4LdkuD2Z2AX+entOexTJUK
j9csUnFAsg5WTgXLFhY91Rm8FQ8VuibLBQmdPHzfA7lim0Zl4C3CNlIK1J045u2H/iUwrQR+adRM
I3EeLPVbF0h5uSd7VPYwH6fJwx56RfJzTtTzC+ckUExNATHbCqHYfztfMwJmm8sn5HdlyT/bdkaC
GLpowbWc1TfNXEfbqUmAtlpvUxOOS+uYMA2HxialyFLI+i53GBTztS2P98CESc0R2ijWkp5s2DXP
mahEnY5HN1S9dtY6E5dxscIU5GD305Hr/H1uOMC3lP+jM8nIIyt1cmwWCROXxioxuEIWcTtdcUka
XFOK2Ws4InDYcKnNcf0y/tN1z6ohHU0Vc2LQee93l0SaYQZjwwy6UAY15weu8qCdR6K9hMy/AlZj
M3TXwemaAnuebgUBtS0S+CzXnrD6oaEaOGgT0YD6aZac+qutSjQnkEUUkZ+Zlx5LOw+pFJBTj6y4
qZdQ/X/2kQSEfmAcNtaXxtfbPVSveJS6mjPrKlElCsrvmCDHfk4oLwR9+evjBvUnXI/Iu5wQMfdY
fSiQgNReRZSoa0522czSGnI6rycllXJ5b7Swx2H/F/tu+FFEs+/MtVgyJcm84ajxg2xO1hlNniiD
Bwnxs+xLckd19vui/+HucFtPH6mxgzP0jPdA125R29z5iyVIt7Qcuj0UZyedyPU+A75iAR7tCgzx
9F1+71MGGWScbKSRMNFSLs66gR8S/k/PHGtvX9tnyxYPhZabJZFcrapxdBXhuMtcXOFitfPVwhCO
rPxxetNxi1rIzZ3Z+5NnWk73UFaJkJLBKYxyL6tzEtvWh6MS5Be9mRgH0k/ra9S0ircIrCsKAwDn
KKXpsafElgYKhxKqtcwk2oa29MP6BuMlZxEoAuoNxIH6ZGjkaIH0XQdf8V7HxBORjbUDrKCyqgJh
xz7JjnGUS5Eo8pRtHJNdlaa0lYd7yRt7ozfjGWLnm+aAMxF3GsUQCE4A7yZW9X2BQwOuJHfMR77u
AXZS4zhXmXBmhMAXLf5ocl2X2i8Xc+YdHY1zouRea/ckyQF3PLm7kpOLxBDUN2yyzclW8AofX+Hi
pPLgdVrEydzEe1gcyzeAYPOl3xHf6e4+29J3THezTWWKmJNyllvRrhZhI3u2e06oEF9JQng7dJzr
TkHvwjE7OXLIn0LS23Nv8ycFZ+HBPpzCMNX9+wwI+ldAWWtacP6Tf15Z22kuo97nIYw6eNq2+cyL
RbHOgUbgTXNTQIp6JETqDx31znuCgAEergeLzGQmYE1gy/ayMhy+nEZ8nm4aB9/HeN241r2QLc0K
TyBbzvuwPJW7vC/+eDD8xM9JcBqsAkq8tf/TK+5icIMJQ8Z00XbDLo9zwu+KDfi+m81KOossdNbv
RwC7+xD2aYwKPuzTPJ+Nhq7HqdrlhXPwzOFbED8NU8IPMbWsQo72XOtBLekkZxpssDa1c94N7CRY
PgXXSnz7ESLH01/mgZXc9aBAtyu90Q917ToM8cFXvIRLdCDkjowgDs06pOmUFQetbz5e450yvb9h
0EqFTspQ4Ya86UE3Od9HpAs3QD13qP100Wsv+gE29dVfeSVFrTIOwoxFAqEt8yH4kNBNjAZ9W/J9
DmUh8C/xw0cAqF4ozbXF5EhphBOINU+oEwm0Hbla74+SIpbLfYsPM6XMesGDuyO9/xexsp7iUDL/
k9jn6pywMVhe7cJBXbgFm20H+Y0Y6Cvd8npdl/qxZNZf55FWDwtYatHuRO4HBggsdyFiEgACXvU/
v0G0WDTJmif1Cmj9znowFxj/3QhMFfWq5wzfi8SY84v6UCiMlQakyuuXoCaZDe0mjkP0gV8+JPG1
jQv96hZSYGN6z6xAt6IcdLuDbsFVfsKXVIIDkifpwuBoBg1znRK2qOhVRFCLtSblfIXalv+vcedE
TTm/m3QiMlCykza0B2LMBEBxRgONjb3VbBiLkjRxpOgFSXjo2cE7Ra2SdCF5VVJRAMg/ttrjX3Ty
uTBcYX2Ls+evnn5Onb5x+ZDheN+MjGHDSVKFBIrdJXkt+BYLA4yA/En1MieX04bw+iPZkNHMWqf4
pjdzjHvsb+GlACNJ2opUFQS8/oOr33JfjHWrB1LI7SQfFhl5lBXB126CU8Y/X+JU9CMOKH9JpQPj
oqn3Up/BiBxBF2rn+o1vvFwvXdoKlHiaRFUE6jYAvggYIXIJwGD3mKr+/KNXAjVMYKe2H6Uw7ENG
CuXbv79GHipFAG3HcsgHgWDQ4adEIYYi17phQkaaxFIiwLA7bOxXfhrmwNS+4BNEERbsZKzsU2nX
vhjcCED9whvS8AIKw5PiGez4KC+3MRCdYN7pElx3iF1pXb/d6csPmSF02IEcJFYya2clJBxyYPRF
3YFvdQ6/oojQgwv5BYXUUaRDr3fsOXNtsmS1AHOSHgl0jnaYWoNBOyJwR/1FSv9uX9bDH+Nrp6Fe
cl1Q5nTdi1cEXeoOU2jXJKUkNWpDJLT6ZM67H7glJ6FHnbWx5Kzwd3g9j5KZkP1lQCXpBO8Pr5gt
rpGyYJ3OGU4dSwSesgNpxS8IqPpfxsvP7oDFI1Ldr+EdF0xirYcNwQ0JSuvy+JUeXdxFu7L5IFXx
bWeFiI2NE7EhIgBRu7gUrua6jcy20LoRAQUURJgIJOduGjkLuAoJdpiE4CxfYACcoFt5kndwdXul
4JZ/8zwQJqSzS4h8OPcu8kndYTl/KX5TW1D6SFeEA8uRWE50GFvFLTb7LmmSwFWj3SHvzC99v3Is
rFCsLZL0YE0tKa8uP+1zteMAOoDpa46EWBSZfq0uVJXFKtDZRlzhe6F4S6Oum7uPGrjiNwaE7v8a
lGTs/yzngA4UMcQwDyeBcLh07YnZzIU3BmXZ+8m+iUbO1SXHb7S387Ieviy+TgaYHIwwKPcI4klV
7KueEkqwX1bSCJAv4ts+R+jnEhLjBCcRz0bU92NlW+lnJdYysXg6YS8Bn49xJnOrUT/fFVFmUgFG
lbc4Lr2+0QMHnmhMSkZ7hM28PrEj1LloxKxPxT7dPrUbiFe7aX2BuKhwHOwJebuosrOLJ+CPuKNc
2A8BL55Y4T93dLDQRKZA9bFZeeSPG1B93Ob4p/DVrcM5VC+GAGSpoXGLRjLw/VZ/eWRwDyWc07eC
qFRKtgAbT3glBCQCzTSqKBGF7BHN0AOcgfWx0ynIfBxpr4pJDXbwn+K7gkfmpcazXjL3T2icd/kS
zLaYPZtqhBkF2UtY8/m1BxXrwTYm2yADJSSHYZ9rfM+QVEEUgVZqGGNqZdDpU2FmJYAGAAR/aeDC
DA3clIC78w/xQGese77xx9dhuJDOCJaqhGeXmoP7ZBPKi1EFKSMW4um8/nrgBcV+yeuf/DTFfFK6
9hFerlzuXmmEY0I3A7Xn9jKwQapxWT/bwZCq1wxG6qkdGBIvpjzSBYyRGXq6guClUEA0jPfphHkK
fx6KqC+Te/fkB4TMKYGN9xAa5NqmlEkahhARLYKecP4+qumSBIkBdj0j7gMe9ArMspNsAgQFN+J+
NnO0J0fktPGsDVly7+WtTIUs850ohU074MMXO9fX0pi8Fdvb9mACzDE2Ze0foaVzHA61+v5x
`pragma protect end_protected
