// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:59 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kffTi7jfGO/hVm8ud/99huiiCohw7ocQYz45/WPFQdi/K5AMUzyBOGFoAVb45mkd
0YikSctlueEc5szdOvQUvnQ+341NI8SZgClHnBMbmCuHP5QxGwB6rJwuDp4koGlT
6uJhKTLV3QPWSuEjMyWcOEA8RXvm69eGvZKJdBLx5MQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1856)
kwoO/65KI5dydsRG+WZlWW5deu4C5rmdr6PXG2Yxjm5hXWu4xhI5P8K/NS77w8DW
d8FMs7cWujHPQcTvTzfy3FB4H0akt28F9SCNfHcxjTGYcTlGSMzBlSfNs9AVYU+c
Uh3MWC14NPYL+7nZ4SNX2Jix1N20GpGbYYtU0KFuIvAUyXp2bxUMPDQFBsRYBrEX
9qwYRboNCLVnXeOhzkCbKA4zzdNS94Ffnnm4p0lmYGJZKB7ggw+PQPpDfJXY5k5y
ebv2zcjTwS2iZN14zW7n9wZBED3rGa8ZwlxezwUVlfe/KsRoCSlTl2NaFYs1nFDP
x5lic9spSlCSWzvydQfME2MeH5647zom9pllQKezcIa9BKqMlFKYziP3iJgAGrUk
OSxUI1sWt91iHh4Bg13t7n1FhxPIiLWyCjkCOW/pZ5NW1XUosk9VdVR7a/LNxGmt
HH0eGY7pTby42zpBodoU+RWI214ux0CG5hc8Q4zh43B5i0oosajxAMMmdyqgwaGS
ud0DJH4NRymZeY0eT6j/YY+UFgQpTp6NHJVqjZXuJ3xgS4xPXiPmH6zk7Zddx9eJ
AWVjMU5ngN1AsCut4a38eFi8HQI2VO+r1a/jUnATgXuNm5LZgYDustIq0Wa4yrrR
rK8tH1n0Ekjq1RxBbtdAPnh1NBgBIYIWmwLB1Tl5/COTOHbca7z7Ju1HFj5JhBj0
268ra1NKB9kPL+hT32KknyiUQRbXlZ3vF3IoLWlfsB7Xo+meHUXNzvgtZBUDqIL6
Ov9LjhRLf2qxczP694yvkkzSl1n6/Aiat5eNaAk5AiCcV4PQliA1C/stohwyzAlK
EgTANeWs6ex71VTpztbRNhqgtPt3UFgm0ti/DqEiU+M60REgReVjVgApGsA/sdam
3NrU/rxPyAeZ6dEkGbLIrcMPI23EhVC0tB5HmyHYwFGGxbk+dAAUaMOKULiz6uzP
kRZN6u8HfSME6NXogxJp4c2KDFn7VnCF0xRSy/4l7WmA6gbfkqGy1hoIl9QXeLE0
9PNVG0rhbCvy1FpVtIkMwTqaX+HwqQC5jwi3JVZ7vmh62NDE7osEgiK1tkdWzorM
R9IYqi+luy6FttXYcO3qYk7Ongh2t+sByO0CEB3/fIPdNM51iJ/QRczC2dBKuhpS
aeD1vfQCxUdIa5g2khl11L+jPp+hi+NITcPr8WSp48RLwvKjCQacp5uo9I75lIq6
vY5CpIUBF89Z7qXNBpLXgvdxgVC0NG9iUCBqQzZfyJixtnrfcF6619TJekInXFXg
jJPAumD6c+OlbOopRvzSQd8Kap5b8JOWIZ4u6DqSZzjcT+X8PMxiEOYqG+Wx3n2s
2CFrdlueXmCoSsVwPYYOg79OWZp1t91zBpmNWCUTIVohc8C9qCPXW8fX3Qx/ofc0
EbGGD3ORAb0061MBCsqr5qUkcsdNnuaU2/7zUWyKHFbatyAglgb2BzVfDlWAzqpp
zeegYeutMdb22wUw3L4pezOZH1aWykluryd8plq58QlRNqIwRjsQQ71jC/RTvit2
6OH+74eqXltV2xP2opkJydqy7OHcndF3mvGVt8Dw4bfs4eZoCZ7ChpEHtuAJKKjc
Gb1M20YWU+9MK/PWWPiFM1BU0ykeG7UXUvYjn+no90FP3cRKGJTzwzLqcoErLzQC
PTUsX12UIg6ZXMJNRM4SCLYLFuCS2qemWRg7707y0A8QZ3vyjy4f8xGCOu5fpJ5W
z39U2Eg5Xe62rW5SNsJmz0xiKCuZ/Kor7lcbSWDwDmWAVVM4DmOPmuHmDXN2Ed7W
KgwwqZT1k5pEQ3Mlp7xb7mxXmQxRWa/sRmlYoJykpdoD9VNvwVEhTAXS3cJDBb75
BThtv9UJfEiFC726gdOE7pzyUsiSo1SXKLw/oMgLN3sbz8Z5qGR6zGT/1I5OpPUz
U9URIxQ9XkY157kJ7tkF7frPWca6H5l87cQ9AvE/ZP0C8O854HphGLMwoFHaTPC2
FUfF/4iN7VgbmQM0q/454zggtjaeDEqzltCUurgdbszEjZ2L2RpwaSep1Vz7sWVh
uoUfXfFTpTMo9W/CLUfQiHS+RaoRqxa+kjRp4L6LDvHI83warsheYoJ/TX7m253x
9mSOHdaADHIUvRqlLHf7ejxx1v6wg3pozKR9b9mIZBLoupXxqr4ejz5E0CwrJLSr
ao22W7HgTnHhmRNVbh1RKkl7CxazZKwyp8iZQICsl2Em0bJUwKy4vBQC7vBPl5cD
YlY0skvf6IrOhkbh68Zc/k5Ap62+iRR4EEVb9cDMRtyBULBoeoCmI5Lg07RSav7P
rxlkJpNusGi+cHz4PyBZG81qG9Hs5z02dCRzdpGg7cONEyikp2WzHi5NTAFkn8gb
TDQKzN13aQvsn0FGkRVWkTq3TaeW1AtSx8O0exatELlPgIuo2zXR9oQh1K+O0Xai
BjCbfEzllTJ3CU1aykLGwg+LgW6Pc3/xmcmPf0hK7ug=
`pragma protect end_protected
