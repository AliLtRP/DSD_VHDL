// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
aYO/uuh1UKhbp3hEuUCrSj7Wy4DUECvO9oxpeagizC1kioWzWFexQALYnSUfvgRpwYZsNB87UUCq
EZeYp0x6XZu1wnLWbjNYMBl3MpkIAidyfktaqTCZJhuQrEElKggjCxZzkW2UsFq5rafZKtgnPm29
t7vx1dLvw8eoB6VhbG1ZTw7rF5yUYafMZOoT/dWrg4MDPn0Mazg+339aR5gaSB3QK2HkIw93r4n8
z3QbaLowd69ZUwYpYn7hDPirm/sRMQVtpXM5LoiqyrAjpHi64JGrxcGrDbXlRELyRwHJAmLEEbhJ
374J7ofD++FsZWX5Ee0FxWx6xwMNycAAoCdBLw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
cLIEnSaWb7n3ZR90WwAnUo5gKa5pIEW0eDGTN2hoO06K704gCATgatmEODIiaIDEGaNJQ9vhKwU9
z++c5Z00vRiKuggc9JyPYwMUIRlKM5xDtIiiymp/us7SpYBf7OKOIOC4JYmiY8KTtuUDUtT3y9V6
yUviB1ibkKr5DRvsfJQgpp2gQ25FPsQdsEE5XEoHauqieH7A7R6lPdNwCEjYU1GavaMfvBI+dJlZ
Bdjvs+ukTNP1/3X8fSWWAsLscGbBdYeQLE+5RJ2kUed2Cqpr1Bw4/cEQTHJhYOacF+znIVa9yE2x
YzHbNalIOr2KCIQ8TSMlo6a5B+vZo0Vx2nCnEPCflwlKK7OYeHF2BxLOiLU2NPfO3dtTPxNauoEI
xgsQqpKgCbWzmdJvpDgan2EjLtZFrcWhIakVNHv8w3N6tV43HnF5S2GhK7D30bQHie9ej/NHKHd8
aPrPxu1Aiac4lsXnzrHQZMbTG+J67R8/dJkbfCxlaTlcRHsFRWf2bCJSDaZLWodqdXuj073qb3vm
HMpCpnVBobBmufqRvoivq8hyLt/sljnJh/1fprWNO9ojMIE95jcij4vwFgyfaL5bftTv9SfjjZDw
h+eBayshlJ2dTJmWWCfiBGtcXn69AFa9MwTjjAuJKaLe4L9wPx7ELFh+u2z4VnH/DwqxX53sHH9S
91XlGOk6kwAH5UcFmWQ6K3e7j31q9UN7FQlK9zDWldV4h//6RuiZs4vMc4ZiWJKkJkPVwXf6pdCM
fK6FUzqHeRNxacPV89p+i1wj/cI3hlBp9OQU55MbH+gjP11KhlaDr+UHKssl5525LYDWPu1n0OHC
oOXLZNbCXVE//mxha6NnsH1sk17afT9HVGHXlR+P/pb/LAo5rU1xw2uWl5VMWruzeaOz6YN+PKUw
ZXmdlt3mtXUoHgJ5j8ieW3jFoYni4iDu2Yn+qCJsYGgTDmrvTwtzbrxLXFM41EU3WCr3mHkyDuAS
/h58gy6oOONogJR7rVa/bTc9HpfkLMOEgpbaK+GNpAnv1CsBG3Y2OllEQmeixzfy11V9lmZoVEcp
3utAIaVEPDjY6XF7OGYdYQZX/xQy7NIZPezE92/N1uaIUrMAajrBepVeuNPDfmnTohIb8h/CZimn
zJJdGHgUi+0e2hcwq6FW24VmGRD3NApdwj1MFGVFq1Qx+FPUsPQLffC7IjdXWO0IQVuzjlWJ/kRX
euQDtQpLliHxIq0+PfmY9WRmmwFzmZXJveethpKJYViJk7bDvHQ3h47u3osdc3d+WFy14ip0PTKd
KyTyirQuSOI/8Pt+dQWuMkT0t2g/NyrLrrtdzHGyMZwg5Eoup1g5w0NpbsPvvDaLI2F7bsaEW000
UAtQJO1VZq1Tq9Helod38V7g/2Wx468nBig9xPIjAMKJVu4iZQ7MZjRnnzHd/fQDxATLVNtoiWJ8
fH9MaV6C01nTiJtWIdGxeqP5ez0yEundPI+aFAV7bHKdtDikYlTlA2zcY4aq7uyc24scK/FCvqJo
u89NcF4scPqbvwLq3Dvvb+DAH6cGai+bEjQP026IP0oBH50RSMvjIAmIZZv+xQvDUhYBugmyiJy5
0H7+uWhuT42xm4F0hp88yLEkt04fs5A/79vLvTaMtY2NqSo6RVrdBawrmuPA82S8YQc2wOLNNZIy
Zm6Ls0B8Ge+JS4jiP4Fg+22OR8PmfckgxP6MMLPXdrSYHbt6BieJi8GWm+3Gki+6ifw3pywfRy2o
U0QHNSSLVWXKNBSKGvfYwb4+cMCLNcPFGnhhlbToCpYAfIIaL7ZO9sVB4DSKwE0AbTiIUv6e4PBI
VOgM6VWknwcVlC/FtHwVr9OHJsnZmimQRtFsn5hy4yG31UQeKNBw7+axsnRbe3F3rjXiOPmMeyCj
dkRLLMfbiy4pCeP0sZkm+Hv0aTNXGPm9mO+gMooVCKDcBc2io/bRqlyiUnubKjEG4f/RBsMDKBUx
yBgWRsAL07BVsr1SMLgQsYCByh+yp7byHvMcFFHY0lCjFnDQauXqJpyr8euLrpWCcpQ61eU3ImVr
9hwA8Mz8aDSKmLndV6wZOiSj4uakfSaaXx/FGIHzYnvAwNxzPVAK7gNq8jX6+fVlst7xIVeTijM+
o5ldg2ofyDOo540Mv5lwq/I4Xodu/jI/V9C4qSPJTxNVY4EW3yXVFZ7i0fF47zqxLsB1nY2j+or5
WAeEYfJWNBtQz0xj+5NkJySlNEACRpZ0YBhHsIB2jFjm1i0xb+JGdSC3wnLY5Hz7jyLrCsgJG5YS
ZutmeI6KXymGpvU+vpnv22DypGLM1DWXR4K1xHagHTeC327YTWLEo2LFEUFsVlLZZaCuj7b1rdSj
y2CA4CkKEivog4MY5jBXRqybObK1uvT1BjexmJJ0KWZPdvRZbMlCNOucqjLJic27ZFpdEFDgr36B
oI5t0CabgLT5wsWKJmIDPUnHcIA4DRruKM+AbQT2zzWnxL4HUqAVcjShjq0tFxpdY+HHEzoM3H/w
6FdFD6MtUMuDGD7iVTuQZcteVCwyTZOHu0vNhFial9QQwurPdnv8ayYS2IMqbS5iolclR1u8NqVa
QQQywLwIqB3hQ86QqM1NPxjIW8i2i8cyM0ZKkFNjRmpoB5pOuoT2Bj39QA3Hk8BI7kKZBsqdK8Zk
DYnzqFPO2pio0hZ83P3vOkd+tVFk0cRSYmIhtG5Tnb/I87lv6mND93hiF7sZFt5zxJM8PUazQiUi
8D6o1ppGWlgG8YNhroY0Ue51eVaoHfBOTxJtAZM19i3ittN5+sSh5Xu7exPIRq+GliZheMW4yCsu
nVflJDMzjs10kaO9J6CU8LcH2aVS0Rb604Jbk05Gf6SaP91mBeXKNtw+WzJJu5Z7dv3J+ij64mWp
tJ+k2T2gEynt6vIKMWTxZKmII0OGXv5aLZtRhekVfOwABQofGd7ZEIeaARkwpgaSG8R+YWZMf1vG
8DUTYKnxAog2CivuF+q8y/F4qOh1IhBYByxogwfkyB7N+plPxwWzhVZcEma6wpCYFqmJCqfvOVoJ
/7CZpLMsJ34utc6UPBzQ9BdW2blz8Lm3ws5AFiPQfubJuPjK04zy9vVctRHSEGsEb88d3amY4qIL
Tys/+dUloMso76rlFrt3lwN0QDyQnFPGVT63+OTJ+hy4iCcZYOWlTmrTjjh4KkgvS4OMiLbSkPhS
20+gdeN6j6gECStNZpoZhFp2jn/XYEFfEeDoH+9agU/p01GpXyQv3soXnmZQTGce7GWuXhRaeKpF
ZAhTu7puOt/C3MAFkYuyLVoCCnaAwnLh3+awoqUg/UuWhL4GtVbR1VFkZMzdOHfRvjAS1ACaPg0n
wcXZKxrsUwnTxx3R0Naka2nStSoP6dUZAMm3374KToL/qx1DmKUFC0h7nRtMGehot3ZO0nKOQI10
zrq5YAjYTXSitFh5jEIlq9YF8iKY0J3t7AwdtXm9mVtNRcQYVSRgpBovhQfyLgSnno2gdWaA1bpz
fKs7DiQU2npJ9dEEg8UIFETApMseRyd1lv7ItAWxLTDfWbOTEzSibdsuaV+jJQfZlHa3S3BV64mO
i21WdgAV8pD4RVN/Ay+gptxn3X8ZZtawph//Wt4rvIVotexVTQF5xiSVr0Ui+bNdcg2TOSgI05ML
yH3PQWJBfaHUvLkeUHDtm6Hwx5HhK/wB9owl4zxfu2v9F6+9MWlMtz02OKxJ1NPRPfdeEiXQPwsM
QaQ8h4eAIV3IhD4gOrgrF8r/fVjdLjw8B30PwY9i5/GGgSQv8M7bM/92BJcwdaZ8ZBXt38rf06BM
Sub7Zeah2gZjXRK8T6Lanh8bNBSyvI7SGkgZBelYuo6cjA3tIhxoF11r7C3UXs4R1FOCzil/9ed9
WhguKwcZv0NKomRBmH43ABYmLgetDrgD3ylXTF9lM2Lscck0rUwj5C6Ocmh94YDYej9f5aItNlDr
4OH/k2qzBm6PhaClUm8H6LDIm6DSbBBuCBj6xx7wwuI7HPBuywxqXD6EaICxDTOs2mfXeugFMBoM
suOA1BZMdl+xR57N6Odv9387m9FB7tKbNyvFpHEvLUY+avz7217Yyb7/aCM1x3hWvJhza0Tq6laK
DkybpeIcRJ+e6U0Tsd2CCc8riM3BbgZ4+m/rWpv0vkqW8lUDZU2sAya1FXFraDL7vl/RHx4L8b4Q
OHG/O9DsbfPQk1EE0fi5+mL5LwDqqf7meVBuYzyN0vMkZnfxRuAnVJet8UcI6YecQwm839pRASfz
V65ejUCyvtVC4F8+aW7iN3+sMzeeYqZgiyDOeNo2ppoq338fwIBx1NEqhVMoI+3RppJPnZI10t01
9/YkTIrA0XJDkCGLZeracppOiHneFw+mAfi/VlXUaD4bqnxWnMR+TfpXkQCpDlR1c0szsdgKeyeK
fkkjf1zCWq31jNgNuKHG4zjUpo9Rc80a01UAAsvILeSo5+Q8pwtFNTMJ0T04EgataIrK6SgI3K+h
nihOaTdSjLuBxO/rNs5D4P1Mq8/ZFbpaxRnXec35HAt2ZmsNgeCwLmtYulSSSCmyprWfgb680v6K
LtYZ8tybavKT7tuPyvgGh7yMAq6yEowXOPtkU0pNs7Crkrn4eaoaulN04YaZCzd+4kW1E++MC4hD
l3UrSHPtc4rKJhgzDvtW9iiMixR13pL6grcX43gA8lVDMwqOX+wNGGmK0ebNHMxWqJjzGC3eVlMT
+NtZEvSYMeNnKjfJlFqOvmfUhNoDrtiEozIKGs6KpSgiHUMjyTV9tNzBSxWSu7HtUrNOd80Mdqxo
/HcTeiPi4EIyVBOYvOSgLohQvagioi71scynHKnqo3uM204y/aqeb+LEmgVSidFupyq8BwufctCj
J/+hPDzhK24rlnnwmSyx3AKU4jzZYzxFxN52gaGH4MaZjN3fnIE2oiHgekt2/tj7CvGIvJOBmPo/
IwnCqBmRr8JdvLx53PmgccVj7JTfH4qPhA+uWmV+Rs2kRfkHEWuF6mQYfbujEl5rY2499a2bEMqv
fWJXcTaEeE9KexSSRd9wLdHfJKnsMQZBv2FLAe6dAjcKiQ/RZ4bV/2SAjAnbFO06XnkiurF9uiW5
1HN0DVl7VRClBWhzXr5v4TguVR2vUh+3ZugHTFC5jytZAqbEyXdj6bYBa71Jyig4Uw1l4lY9sENi
uO7s7WVCGgn+HSX650BK5cpoVvDkgyk1E9Ue9jpWDqhvt/JUxoHpUR8MQP7RreGRJ9Lu8jtkHzIf
Yy9uKBrvWOyMwQ0Dp5uh/ZRc5/Jsu7fHyuu24woGDHoIKW3u6ExZ42IdCoEPKKExJ/KXWTKwzzgF
7zcEf04UESUQ9YlAEf+1Z3WP5sQTz9aWc7XlNVL+tVNFbjV1PDPuqPHY02PMh0ZAIAyjGSZMjqoF
5P42LGPOc/I9vpKSdcybVHVQrtSHwdaUXRzP4q4wEPqTjHfCuaKcJ8zG8HwwJ1qxRVPSCXyjprOt
Ah49IqqNbn8+6ClRAtGdwOBmDgixw2x992SE8rdIbhJsec+e8waW5UL1Fm6zmcemL2v8T769F1L8
2BX1iMtQp2B7DtD0XXzC6/vB8CWPvyDSYkdOWowj21nbtGYfl9B+vs0QifWqgr07/uX7LbDALM+B
fP4TowNTaq4L2sc6dzYeoaPVuifMXRfxq7fsZ8D0msjiEBXyhLYuh7qRlSehiMbEWm+XqRp/9bXa
8sTAPK5s8/oH6g995TKjCb/55cG/t88MjgqJVGqv9PVrBWBLEt4eoaEY4FfMdHn4iLez7YF4qfoA
rfYxEnyTl/Mtp7Ns0iBSo1jVllaXz0e4xZazFUwHSKJa713oYX5cHKndg2Emh15F+5pwDqLXOeL4
2DEpYYzqokt9UQcJhWIBaFN1BcGcp7R8Hz6F5fObmatqnihM77+Ks8F5ICprXA9DPqiKDJ4yRxQE
rEW0qLCF/Xcfe+yFgf0oPmiigUyrsrR76U6cpJipAWFhZO+4lUR2YB/Kk9cH6yJ7t2FSh8Dxv4ZP
PASn9xQ4PBsDH67uJdFMyh9KrhHIzBfLVMbtU/P//lb4/lCV8LmLqYG26r9rMEcTvz4DlBDuRV/T
lXWwWR38K//1tKyZ2g026e7L4gN5phkT16PvIpQbm8LIyLVyDC2Chv3yri773HqFlCxsaLsuk+tT
TkvaWKZvbv3sUCJe0hbR8ihyon6iQcze2fDFGSBwnPkpe6HlmwqpkUi+MPT6IuTB9NR7I94Q9s0w
bOxwEcihgik6tz0mmME9opd60Y5MH54TthekkiBvj4M9vg1lTCDgovs6jrkrzuZxk/LB4XCEQVS+
nRDpi2cK56aj6Ewn3t84To7OPgmpUCFtMWWDXSAXLcITR2Zxes0wfglZqqSmbKf+RiK3piwAooQS
7FprrWxs9OhYgn6gdTCziZ6D+1aseTKovk3G/upHONnPvkMMMVnir7kpIoqY5Q4/tMkCryRFqcum
L9skcut0LqOVHUC2IHpseQ1w+yV6DgTTnMpIN6/uHOKqhJWbp/CQA9RhaTGJ1mgPKvqd34y7tQms
dreeldp9N3MU8Qsk8sSE52mU3kpgT2AivM2Sbb09M0fTn6fWg3Ys5hHkw5kyo77nRfqgXO2d7PJD
b7awjLZvum0AwHOzrT96ZBsdakKnbZ3gw6qpkH7k0YhFvlmql2e6dj6n8bG6KuzmwOSK0WUBwQ9C
OGG+gIDaLm/Ju+3ZQqjSl0vWOCwFDXHF2VaLe1YpTIe0sxiw1qHf1RqFxCdwFGcfnKbXcRSf8sly
9mTxWopQbhYdxAchOuGz216pX/MO5gPMMnTsvhDhgmfzrLvlDjBjfF2Z48kJkZMh05b+yUbVNORw
l8rR5uGkPSwDCpUbryQm2rDagaMr3yxRa7bBR1+wQ3+uZ/bfRl7HQNONhBsygQLrbXLdo4+338eQ
7Z4ZW0z+5iIST+H3U5mFF+8vxpRR5u69CdlY8bnsXlyYFQeRzRoAOVI6s9z/hGUFJVih1pA5PsN1
MGEQaXegsdiQ96SE8KtIGkUV/m7n459kA5//aeTOE82sj4VWn7ZqcC5lIO/WfhcyYv4U3Mep2uEg
VxuwGWZjppjv9Bi3nOItk5DsOyS9Z8O1Uvf/N4LV6FkQzYnIHJCUGSdfITztBBBsca4zhGT473xb
2aS95AU80sau/R+Me8Og2YGrF6t8ySvSPqtdras0JRHdMIcqEIcH2sbOZ4sjZWXTR22Je7wXUWmY
8xvzBde+L2LrhyfUdTIj9jdRg8FnCBsw4muSTOAs4E2vtWZABMhbpSStCbae6R28N18CRScR8/JN
vUNE37RofWO+fbSewpj6deTD/3vGRU5+5cgWjdSJIrmOO7PtupmnJLck2KAvPW5Y5DowrHbnE5yC
ZVtdRnSClj/jFvU5eySWgLizsjacw0L5KH35j61Lvly26fsG3ILn3JGPAPSkBfFSXgzs1x5i/hsn
w5kTFkRtjOuwD66tosBHepOL03Sg1iajMBsoZaaDelq+aq4wubKQB5VCejGroEdJS3P0eeDWDI84
UrnPExjZEAHCYEdnUErwHmscriqGRRGrz1xC3OKYFGxx4mXZKwzwwbUbHXWcvxcHepFSA3gdNfdJ
bbTpaS329J6s8D6f8VM0cLznehGtpFIhYiv8nnn5znhJVF+1OAGEfey/2Q1ppoxj4hJO3FNVlNDh
IN1VkHOzvCyoE7oV84R22+lETvWeCEa9EkT3v9s2jSPiHBy4ST5XYUxdeOu1XNJSebcV/CWC11vs
2shLMIwokwVpr1lSP1qmQsIr7UITDtMxSdYHvsqzVX+MfhQ6vGDkW3RyIvMjcLKT+nHfx7wGv1M8
Ids3Uu8XBWBs1T24hzwZF7z78glhq3rQAlIfy8Dt6ju5gFLWOgf/b5WZb7YXfLGOQfGTGKpMVNMk
HRQgbhiPHzG6lYcc2O7VT++dfDPvyMCqEBSPHzUzqZTU3RNIsMAaYE4c8pIh1elACYFNAog+wdSz
56pTqZt/RpVuKwQ495qfyzFSQIRJR4/RHd21glprCTTDB5jbnBIDmiRzzH5EHhLXcUshI9c5AAhN
KqJO1UwRz4KRdeH/DSmxkfLff7X4zYyu5aBzN0nO2V50xAwm4nRdUcqqmxCKkDD5loEuYF0/nxFF
fdJWZYj79uhZFH+TGOLm/B83L88VOiypKAjcjesXAo45TjRVrwjRAFkzJfLfTlGlk5LmHbCJc4o/
ha2ZR8XdmYnI/JCriEJTU2I5WUCu9XQzHTE3tsVlxx5n6Q+5EIE2Xa6fKeIzeFEvfSRRNRXuCly/
Oxt9gDpCOjZ6K4Cs4wBTrRaj+NNEZvfLSYh316s0r/y6m/yjyv6ThX4Nw6FbSwn2iz7f6QTMJNxZ
xvVfvSyT0COZcX9H62Yn91AlBgBoGP8mK6A+4fVSgZViv+9lgvqZpIi3g2w6oDon7pRbiM3dh7I8
/aoRM8T0a4rvFcSX+nm3qVrxMgnPjAVxpWozVRL3heCeTGP7aYy41Lc+G4NEQQ25KTHWYcoYxzR/
sIUG2Wz7X6dCJ8rTDNSos3OKrdW/WjgzDkn/rowJEzmMl/6hDTEMrli4X86/tT+wn4iO10M6deuR
Pvsc4xJlKIKralyfAqJ8X2Zt0oUPPMBWBcHgPA67pEEBTqXH0SvNasS/9PcoWiv+okCVOqjA367m
EdoMCTUpEOU6QFcUKvKVlNwAigLOPp5Rfua88PMcS+wYSqCEmtnDQaUoU+CqdW2/nlza+wZ5+pUP
RfWsG9YKMQU1XUKkKGCnLn276FoOPWtL+0CgWE4QE1m9ozC/4g/3JSJTWs5kUM03kjBD5YPdgRro
SomEY1IMMPDwIUvngq1WMLcVa3VGtfsGnD/z+onXsh3yUuh5wvhVvkZyjJnc4Xg1olSRIfownWFu
x4tc2uu9F1jgkGKBqUYJwmBlY+AIMLZgJ5wlM2l/kyAZ0aeDsjhlrCkjrvYunUi1T81RBu8A/V0x
Tgm0kQB8xQcMV8aFfdiA9XgvjPgED4G9sa7MXuEfYTr0QyyeP7Imeu2prbBcwad8/ha0lfhivEob
dPdS4G5wUuLW432Pgn1Xi6vSmsz9xIa84bnJEWJ2hNpNJP751iuFfjxCPaulFcxhLpkeTeLc9nO4
Hr5Cm1k4d3IWR5MSbV9Q/oaNanuXrj/vnIkjmMwQpG0MjaZFb901dPbiRlZgLAdqIkoBV2vKxuYW
llFY2KApV1SJPb2h62GroEom8/i+SK3XRnvQQnh75Rj7quBUrl7p0Kifv87ivp0kw10OxocRlc9L
V7MgOtm9RL1BNJSxrNeCfgUQskL0EF34tb5wzQjOwr5hMfOQXcjlWkdG/JOpi8nyJXKX4qiA2lyu
UwwJaNVbRtW1bR/4sVN5e0ciuaik7rPDzY3hDZm6lCnGg5NTQYdq15V/YM5Kd4gJ8GeLHNwSTcQf
jH2DcsKrP0EO94HDS4LWa5sfQSBuDOZmFJYWA0iov5wc3zE27PoHD8uAAF9LCV9Uo/ZVlzoQNmRH
dPgjUFNUqdsnBXOjZwXaJMGNqGpl9T9dpeF16i0R2FVGYUaiCeNyZb5NZubZhaSlMWfDKOjHeXcO
SbInSfpQFpNfma2e2s6zpeLStklXPFDQ2c0cCQ3dbCEdzUDSc9Igf3xPvSRm5MPQn2nlOibRlCjX
n6BHek6LceM0b+qdWK6mqn8+KojgfhKf9u/ZGdR6w7ie9oHccnwKiNmNZiVlGk133jdqclJRmuiG
18TNkkyfdQReB3R/o5L4koNvHwS4H2csm6Yn30GfGlFoKhZEVWwyoi+hfblPtmyk6AAcIMjpuLSA
ZYVQ0VyvqZM7ndyggjyX3dbo/BhtmUp06ejlhXdgWh6kuh0+1l8pTKpKnadnZHL8Cw6QfbRTy2uO
cVmBmMtadwEuxqYfX1g03VXU7OuI/N9UHJIOD4yz2gvp9b1r5VI52EARKxwkjeZho/Yy0hxuTANf
t1Z5O7kd+QrLAKoCfsj3ajv3/JH468xfHy7Sb3q7MCrrNOYJ1voLpf9y0EwIzI+D6SBi8ApYA2zr
VIlE7nyqijubzN/U1Pwi9Lp8c4xTUfckJ6nSfy/eMkY6nMuZHW9J+2/TAjvPauAqKiUYPGZc6hjW
1Bor2O6XEjqb0Z/q27ia7mLGQXZg71O7MlRhqCwoXBC4KVCvqF93wVElRMLIpZSTiOEiFVh74B5F
NH7ilkxF1IzBKsn+eSiobofhhj90sqUii/gGFsNem98BtNscvvtTXEbEmMbDWXg8pUQjzkVl6Tq9
ZZoQiJI42/bJM1a1cqn8IZ6q4h0oMR38BYytC6owUNjXIAmTQtZgja0g/J9Mg7NP1lVnklvt2avp
Dx5H1BEot/YdyKl9nmz6HhAMoJWkTvjI0KCyM/E7j9xOSfukXtuQLUe0SsD5m9g1sKlauxwEe50h
Xq9Qikb9Le0YWG9R2KAQ37v5WA6iB4WYKhoj8EvMMtT48ykTwFkRmrNBp6J1SdS2I/Q8PPmTj3Ek
yWpfSiGa66vqOt/neSkFNNCVvB/eA4Zk5y4RVDb+K0bKzXNPiT1An/3irPMFBfvkz/vT2UyYeNaQ
HfY4qpA5TYZKq/2Z83AY0uSlacqZac4dQtXa6ePmm0fA0IPWrjuqclPvchHr+Sn0DlzclsPA5AuH
c+WpGBsdnUfw+8zKqbN1fxGEJEZ4CRwd9m4bnj1DwY993C6ojYUBJY6BRuVrcQBsQvbWnD3wwhgT
MbtetigzDKY51F2H78Ee6rJWBelQ/jKzxbepn9b5chO7ykc5IcJlEekKSvMPx0gygoCKL91Zt7t1
1pfoOj/yi+SpWgm+BUtXMYLvkn/mOF+anSQS4/4dVNrL+FnSsoU3BCJpOgEbgOFyCviNFDyCR3mb
56mPzjqATC23AkndHGhm/WGjBYpIHKPzMpj0h98MGLqEy0PVllyU9pPFyk0RWO29Tt5kA8QZWBif
eYQk7XVi7E0yihCsNleXQtNs6f+cLjtcUrCEMxLAz9rKgmqADF0rQ0BmIb6K+G4yx5R6+eQPDL11
uV2bb6P8DZq7I3gcEaFuyR2wIDyYsosm8ftg1de9WNN9JQq8Z+jP7GqIzALnM9qQPxWE0bDg+9Kx
uuPKIj6zsAhtDsDrQwOsrpuewYqfx1Gn151IlScmLRaxf5mifdSG2pLDv2A7koNfxDh2mFV21miK
7fvMvi9vLgZFwe4G8m5fb6YKBSuezk/RsWgYedzsb27wGO5QYL/rjSH66jcB+0a1JYQJJIpm9Lgf
dWpmEBWW9sQGImf7ToBLWRKUNGtpmuGvjxt0WfIzUvPl16vyRy+QrXcI95gZPaZMXBa7CW96EWRG
XOZGlBKAMg2IsdzwjazOZ5M5V+zX6V3kkBzDQu76JBBNyzwP1j1sCt94LKZezewKlMKVUFrSWaCR
+YsE60K/ysDnuIBThCCwREgaAoGd7xgfJNjuBk+EkLNlb3Sy9syafGy+qzlzdV6kLePKjSzh1Y20
sSf95aEOXg471BAsyGxgwsGjZ+hKB2K10WWTNl8QOSkcS1wJh6snwxD3zYQ4bbHThXq4l1mKf2ph
VAt7Vurq6c0zi5mnIx8EQ++sdU67VXIfA8dREtmCHYcKADiBrO4XSXHc5DMioooYwYvKm45uqjb+
XQ+orjvnfUru2nJY0aoHb9kHMbT3xl8rgEiC1xaxK72mukl0Slr0vB7LlLTh5r4GfU1rWS7hkd7W
JDTF9mjlqD513ScYlcHjiH0C7drFE5N46lYUJxyjgJN3VNwnpuqeTyP8ku/Wzs1Zg+zUdKkwGell
JboIUy5lmAPNOLfL6Hxe8DMSBFxfz33lCE1tcvOF25R081EhSw7L1CVj+I82eP+hnolTguwQTaXx
2N//DriMg3m90bxqsQTbTWb0m5JDDr8EGkPjLsaUTbJysqH1crbMEr6cj9I5UTig26C3VzrzVwOZ
QlLL4ccLEyEleNETyBHnrJ9WAIkOCnEyhUXV889C3QjZNJtXn7kfI19ffRFf6sstqRZD6krV4tXm
YAkbD9YueHPzH9cS/kuOmlq9MSxjXi6ESpTrtZPO1LDyPkzdn9aHZkuQSfh8PiaNdQDz+7lT+0jm
nhRyUoLGtCCpiLtenFqay6pawGhrT3eWWLVl2ELnke27E2ruIyt7F0Ur2ddHIcDcXV2vI12XQ2+t
eTUOTtyjSxoyXsCWCrSS4Oa3YeYT4oeZZDGEQaVdIUexBzVC2MXhk9UqhokWM4daRvsQUQTu8P6V
+w5x2senpAJ7onSQ2BA+qabEfLaHwTSXAZgAEftSFv+jGCD7wrVljf8Pe40qBIEWnm6Mbamvjt9B
gYik207Dg/70KZcHwNWtzNVNNu7StDbuI7zwLzQL34XQaKPff6mqPZRstbhTV0iBTZDYixTyvYBP
KZ3sBmtb5CHL3o32rRCZ4FcWTUsxGSTmzUYEpTc9rkgr/mpFnEpK2rYnFJCzkVwvEHW6tVvCRBlO
fkwLwQTY1birqGPj779QqIBGpyeAfG7zBkXlDIeV4MZ1v6z5jO4HB7I1v230+zuBpol7ks2F/USw
8e4KwLPSsHDYgxatX5d/qIpf8tDTWKDmIP0+XU6at0Tzt8gegj/FI4c7n3QrHlCKKYeF0HTJ7sin
FBKFVniF+bdGgu1j+Clecn7KKxPqxvn6BVv4fWKkizCUBhQ3x+7W5B3lOpm8f1Kuthb2bAi6Jnq5
1JEs99hmF7JqtPjfz+cw7WeyClARSPO71bYVNwowrz7CYezIlm9105iIE+quyhytbyw/yVUCgCyl
45CGP7hUfPpnPcETFl1SabDQvkzQ2Z3zfLtkCq27VwzFd4q+L2GFSMycneY+KhAhx8/FBoHFgm6O
xuNwBRpz4lsgrsJgi6JLsi6FDywYPhGCcpbWjZpJHAn/3ZAaAKrIMlXrR/vV/4E93sOO0JSskm5z
Az5gfoLdllKjxGIvaguSXhy2OSag/808OJjT8xjQJFRN9hOyQc3hGiJSgZaMKvQEP6i2Uoo/ckEN
eCcqnO3ylNV1q8TwH5/df5WCwLQUJEZ+3iMSbRjq3VqOhRhZ8yTWKehHlq9M5wlgHPWHML96cVjU
gubXHFX8b/Z4NQdALEaaCeEfUDBH4ydbfhIZMIOA6Gywd8BF+aVuYAsBeGWCcxR0f3z/iO7yj0fY
beVwckbjrrIKs5NZbSll5MvYCmZMyG9+4rp9HZ5az8wZwPDdx6YVLJU+i/FBUsLVKRAzuKIDilKD
eC99iIYQ3oNVG32gsxsK6QNWJp4C2jNk532r8ny67/6lvEn4aVckmFfKzq1CAnjKZhM/lpJpK16p
MxNGKlpZoX9fTxZqJTYk/tQBmfmADBbCvcc6tfeF/6VoPJfPwr6CLAeoVN9f6rpZcwqX7AiPExk9
A5yPFSpbPetMA9aDyCOZ1HJipmClvpwyZe0UR0+zz1NT2pP41oSt0WHRCMrcJlKwSIvFEuromvQc
Qqx4HRkmF6GtaaLB7AH7HuZzuyImdNn5my3Hyh+L0f5rB7pLiYcRcFBh6fS8At0wM9jyPToDVSVt
/WyYw6qwrr95922iIzbm1Zjz3aBL/VzxIVAoNiJwXCYwLcfNj5Ug2KG2A2Iyi9J9Sxj5DGlD8OdI
vZYGMeuwEBJhvlWcla8ZpYHNtOkMZpiNwPbdbEeDzUo8e0y5JTlcohmApkDroIN8aBnfPEdwIDCc
qsBD3Qx9uqBTRDQxAcbnBs5FWUYHrKfpUEC2GG62rssOHelMlAkWT617D1SzmD+VsN7CJbOlzTfh
y1jjOPB/2uCwYF9fgX0ebFFkMtzJ5LPwU6jfeVcZL03SFMjVAVMYF1QnMBUWpA89vXdqcloeifJw
Vpxzd1y6/Y0zHD7aMo+h4Jp7Q1/JJF0HOX43i1TGDt3YeTNxvl1b2mVHzGwb0BHFZFoho0Gwtt1z
L2aJ6KLR9zKqjO7HdCDyJ4WosmilLpW/203V4qies4ss6n//P2z0t6bfuLOHC0GREntwfI4hFmax
rNAUc6SVGVCzq2C7kFiUyEWVQ2FmoIK768OXQnyiEl3W5sNn97RBiTsDl0iIWt78cinuuaxiiY3D
xKyxquUBxTOcRHjKFiggsMHDN12kTqpwph47LcqRbm9opACRm2cyZbHoRqzfHYv7OTmjqXuh0NWE
8d+bLPcQTqOko+t0GXaayi75DcBeihAYcSSqCAkYnrTXA2zdat7TZToVfgfVQlOVrJeYEN+Ue/hs
gi0ul16Ur0iubLIA4SYuHkdZT4w/cgXqFXH12wRZ7KLLs1tsT79r+MlLfK9a6sd8+by8kB9uM57T
pDkBgaICV57YYcwZBwLucvDHraab/KpnfLATqUylqA19O7I9gkSnG2vEtPfYAE2t6PbqNT61VISl
AEjRhYXLM1gsLEa0plsyI2/1PREMreVnUbnqn0Hqi7kFzOwnoMryk7ZXlTtaIT+aNXJSUKB9ytQ5
/iG/o1rD80UUFYs3XJx9CmGnLwLbpiWnC4q7eWdYT9RYjOM3Z6/Yp46F/8zvHviofzP9643C+Nmn
12eWpMWVszucMksIu3WxWhsLnYy5JI5P+TjpU3bIaghWiMxAW9ZkrZOp8rpGEc7SYRNg8YnWWBrL
1mpU18o9kSUuAqftluPokF94VA7/PkEfT5QBHSzTWTsqANqSyairqQJixLO0GFKwdoKHNOB0wSyz
f21uKyH9eYs2+qz+NJlAL4THTG5X0hGBBlyGhtLCUmvzDtv+k1eHfkOk6lfyJvBoQhc9XqDv5P3w
cs/esIWNVR08NIx0avmC9WzSJwhL7gYMcmEc2yhrMijHFHwCbRjpWkxiGofeQlf0AI81pVZ9lSDL
GINapxP/YUYVRUn4ys9USxpWPb8rZ0Mqo2z8pI1W2M0uZwgELtI9KTC6DI0kVrYHD9mEasDJG5Je
Sv27B4spaz3afyMRgkC5b/m4u8JkaP8vKXDzbNtSQxfZsdaGpnWjR1JXqSnbBHH0WTkrU4gSuQB6
NjcaBI7Ec60X0iUYu6fIUOrpgQZseMHUdGUTTJEsv5PA+iEPtjrjuQhFKWrOOQgVCPCKKkehvp+L
Vu4tRQz9oY71wPjDHs5FsDdd64N87sFa1Uilqc5R83A5TW1pSLZFo9Jmf3BxbKzSajFoHDw5SWpy
wxH/N3ng08Xo719icYexIPVeZSAY3txcUyRNckatgF9wOiEHGCXy9v2vH8xPYrQcs+gCo0rFgkgP
t9YwSK15nR8/TqkmDPFkDPyPfUcCrgcNo19W0M1nU463TGmZfEC3kAmuAToLtACZIeo2W/7rFmrN
Lz4HFYaKPZkmbdZUQQxMb1bFs6TcWjbuuA8DMWutSaChAVGy0ByUIB4l/9ShaJoGTUWNaAf8JR2I
Nq1kKkYMnLUPVzBMV9InWk6qLDzv0UGYvwLc5jUBrwdl55kClYhcKiJFD3cNH7Q3rPzohtE/tLL0
0s+0BRikSJGjNquNej7KyHLBNzyM6akqM1YaGh2/Zg+cepJ40gz2jeNZ9+hJ5AfWVgsUsu/W2PJJ
P4+YofiKoKs3WlpiMTDlm1Idw2eqxcWUcWG6f9h2exuCa4iMx6UqYGphs7CyF02Or3Obi5Nd1Xw5
33DrWnLlhxbibdOkXvCm4qfhNyTOW7E3jcCCWYZ5hp5wnrgEfgkUiBwSpSppF9ofeTKQd1PIJjVe
x6PLX4JkwmheZ8PhMPfpSuVGTNXqidvHsZY+wZYJf4V5VXooDHC3ki+A+CYY/rYGsd5CUYyJNAAa
AdKun367F9iryKF10NhL9bc/zjFlbPLwz6kmAefZfLxfSrbeHd2XTlxadu7zTA1AybKqWhwhPIIZ
DVl5gSBwjdM8SNE0pQ9H5kTItPJibsktYAcbAJnmrQlseHCC+BIu7Rr2O95xssB6LBP5DOtrmcSQ
gnHNQ1rUCQ/MYwN/pynjp4ofcTUUztYRnns56QnEXWau1d3zwTWMyQDyx7tKtOg1G353in8rXjyZ
SZrR+0Q1caV0I/Hh/TfN4MNpLfHe0c+0nVOcOExwULzd7+s1PF+zVabi/svN8Hq0MmL8S53t4Fwz
LigDxf+PC23OooBh7rhFY5/ZiRvnJXqUbTqQwnWrMKCI0cmcH/E4q8VNBeo/V5ZZgBsmgEJcmnYr
3dwVZdqcWJ558wxG5h+QGSS2qai3gbKDqG/Os2ATj3Gw90FpXyRuaGlXVji+4BhI3qE2OpjjPWXy
jojSBJjiWA8P9JA6vuCW9dXIf0CSHUiyYNkcSQ86O7myxg7pPPHKUKBLvbYl1v1LeYE9Qk2J7zee
cH5toOMNffEOMFk/Vf4ZuqQi/SieYXC3CBC6A/UHN8M6kSS986nRaOSZ6dUVONzchxOiVT8AfZB/
Kh52LoVQJ+s34bIwQo8WUsimXSZ4MDJm6rGPRY9lTDFqrlIR8yBVYnsoskBUNxgyxjGnSRNsBGJ2
4Hu0Yq/zEFE0YjHzJQp+Jd1GdxTeR9amjmUMNnU9hqL1XrnS1HYgepieP7oS06MJqhAfR8tYpopw
87WhIA1y1H4xXI92S6lkx5yXhSRCOfnJYHTjW/qI8Sm39sXVUovLGjE8Fjg60/ghkozTn/cYsNG3
xrmi1cc8MCix7uybMeBp/2qoAXv6kymb1gTHrl3tFUAEIDkuFILsE2iCT6G0E5GowBdQAPjBy8ji
NwAoF9/0h6kHEPMBDGE+87UHOv02hBztHwwRcwfqyoA2CAjbM1Ft7Stm9QdiLRm+Y0/MrArNGLO8
H1l6ADw+0GmdtR3iQ4leasrXDJUPRz452TA9modKDfGoAQoRNibYWWNxqYfYYe7otEiWGvWFcGSI
sN9Aly7+qjcll+qp7huvcYEcjiXzpb1fTQOVjmUBrA+730hQxJHiofqcXcijkJ0NCEyRo+zAGKSr
Iz0PRl83QDVQsR/WJJCCeWQEocbNkaB6xCVZSrCFqfblKibNXccDLf0QO45AUBAEwvc7W9+X4z/L
a9lfIkyL7DYpOlPTwQdzS7PhERZbi0E/odrCgVa3hJkJJ2eddT0z+fy7WnlhK0ikS7yjRkvCyIRV
+gK+8yXM/r3P9OiOt/5nBEMUrOMX/eDGlpzn68MVqtqJwt61nVTpNo0pP8enOYAfZRwMlzZ3GFsi
Ka31oN7BqOiw4bE2Z6GVdg8NMPBpxkSH6DqcOkU1aF+QBQPNb8Rf6k0RYD/Asrc94M6i31IJwGlG
p66kAbYBfafv+vqojm1hX9O32I0QAO+80aKgM1T0BFR6f5OsBDW+GZdkN0R9GA==
`pragma protect end_protected
