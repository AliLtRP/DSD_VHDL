// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:46 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RdQvk8pubDtk1PF04TnMrBfSUMEDT/YIh/9rMCEM584yp6dM8fWu94HlJpw9S1kS
RH3oKfQagSJ8ny8NKZ/GtuiVD2WsF8R2yT0zUHhXwj4VtT/acwsJ+1Q2oCtPwc/g
iRS+fFFQCOLGOT8pCxEhf59g+jBqWDCv5Z98zSQgzRE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28592)
/m+fI1tXoWHKHtwir2lh91L4wNoB7RJZS4Ed5ev5YkkEm5d2r5+gI/CqRlYtni8E
l1lLS9oSEKlBddE/9RRWAXsJRrEA3PUDZKSvOaFjAAyuwXiG/Xv+IAXyUdby4QUX
oOLRdjPNStpK1hvt2puBVrrNSSOF11YlyOxrR8oKmzNZlhgptt8m/JQOHQtcC1Oy
mhopdrJXuctWCa4+/YySK+EXAWBIOe4/Iyun0mFjXuhtst0AAxyhVx4+oizgSU1f
Wx7XKUH1Jw3thmOclzavNY/tUox9dYKCuZav+hoziIGxmsVXnc2CYPThi+vBGGO0
4KymUnVumZ5XAYWgGLrnjNoLopJZ4Vl1kZAwNcAsoOS//lp1UxtV5+IV+2BnwtRK
C9q2K+jAr4a6wPmnnlt7ozFh5SgdAIW+g8FharXIpVno1vSVnbf47EmuQCQOE9A+
Q2ae783gtWYoEFWaki1o5HsynfRzLqsbw+J+xFVAo8jQ8K70WFB9WX8Evc0LrH6z
nMv1injYX6X8ay+RDGMYU/g0WHZ87dUDoryXegdYXj6v9NXy3xQ1V71DLpA7+iYd
CaDFBAcZSHOdrytjQok4NoHBOshh1hMb/zThqWtb0Q4XF5MeORgr9qkG8/1S6fWf
UEw+qKfwbTVe8MT+JBaq53URa+bZjYMgQrY+YZJ4G70BEYLoZP5IBR9TDB95gi6o
IWBjJD9mYraEtHrtGhGcD0m9ctmQpj5lJcpd+CnRzhz/NpULQPTH4kiFIBcQhE8f
88mrop6hfokbz8d8pxOZ/fyg1EPF5P6Aof0uoDdsDap0DVcEaVO9jNdDknsNDWM7
x8LDW1MVnrvhAIu9yu8blO3mMLcD0kEG5sDcj9sMFjbV23E1V650PE9y9NU+E9Fy
oH2eMwR9evUnRr9cq7ub3Af540cBGpX197l5oPvVQ6yMKMWdbfK+/mnJJNLmccVo
weYi3F3k8w22UE1em7UuE61euGv/iDyD2woetVGWU5oKENvxJ3QJB4hZUuUG3QlZ
2MN9dXSWPYfYXcyK6+5SiV9/c+uKiSm2bCNgGYaPemmBc8Jaj4Lyt0fPO6+lWbb3
J7Bd91RHvBs8SGpg0lIMWdbHcpXQZw3uoEhFHcrPj+5xM5L/q6H1xtGwWaIKBAqJ
BdEUXvyYOLWBy9W/Tiodrx84i42ON9VgkXsFhLUrY1eJivK8gxAoA130dsu+/HPs
XhJaoUGhQKhJxXGEcXFkWuqWk2GV8ZAPS1TU8BvUiXwyxoxM7rFCCDj7Bktg35Fu
ajB17q0kCKqS5tnMCwnlY7Z0HDnLj7LEd0B0UiJilFo/fju2zYEfPbESKQHHOnHu
n6oKsLH+ujRbE4wxTWXyNjjKZP2EM0KNDAJHDxlXXxO9ka5ocwyHJ1wu2TXPsedw
mmcNoCufAHl7+o0BAzFpt/uszVJgZWzelbiIc3ynLIYo9PXZyW0CPTmNB1swetlY
tKIWuh+lUbqqrwvVTPI83fcTRCj5hbuhNiV6bX+40es1et3F6PZmddWretT6Nkoj
Kt95Am/EWYIZR51kQiDipnv6jseID67qKeT3nBImIKAQlXK5XlOdAvk7gBLPEYte
M/6CCnMrbiOVMHkG60Ts3qKO1Pes3MjOjkJ/3954TJrYfUV7/ir2jxYOLI7rmA8t
67snI5c6QbtIx15g1jt4aEvkIEfpAu4rmf/QPgl6qyD5IIizGDGNhaoo8jM+sdmG
XxlHSczCMbWFHpn5CL0edzoD2qwDulFS3HJM+SAlqQgdzkWZ2YBzPrJNuyWTun8U
WdeOKMCdmNvFfgzNcgKwjVCV6kxRoLB46GSuy3RiYtvYtU98jeK2+Bvqs/PCb4Bj
W0+o395GfjFKIdjgYpUdPA3aaNWaQIVKBbfwF2/WbmTV+txSP3HnubSnBUJsQItb
z66hNChBU5xV/H2IlD+VCfSWIbwfOniHUKDo/9FZPpLr3tAApjNBl+nhhMqDND+k
0yyv3QIYxqF/SXptkwLJP+PnG66XnOPlU6RASrYv3ggFNn/n9aEOtTI4wmoq/yKC
DtWTUxToFmVGrxFRv5JxUEpLCzFNKnxOagDLkMjIfDi6fsoQuSz3o+exJADWhftm
DlL8b2Htfu8kb65egxBAj+jCNJM7pA62GUmsmNQCRwNL5TP+IH9dzFNU3mDd6E8J
Rw6x4NJ7MA6ZNS7QOFzvj919YQyf3O2b8hIV/JMSNj3yDmHmJCXGX2PG0KYZLHog
ZVd7bkktk3WJvi2lAj8Klgh3Zsrd0bskydkSKl/HwKuh/LCW+ITj3OTs6zvIe1ya
SilaIkMWR7KHg8wRiQCHOOerCczOTWmwpCPg8KlDTI/TuO5W+1DhxGPSWP8MkXLY
lkp2FiRm2RlmJGkabMdZFyUWXfK5I8J9yz7V1+cL0ghnScKzutxFX4ncgOVbjxO2
/SG04IRoeExiaR5VDXV1EFEmUJMz9ngRqsuywna+zRA8SklaryEErgrNeeyvl+sa
2xRCGQppaW4PxQFhIvDW5uKMMKSx9pPSmUcRPz/m8sXFDRMz6686aCV3mE1nz3m5
GJwJsjNVIdEZZDYdqIzI78hNxyGf42icBx/rCkvY3BaX+QoHy+gvbZ56a1tzisoi
z4j8yT2M7C+r5++OfkzzFj/jgJ/aeyR+rSTGjdWzAeEpE8fKXgb6SE6ZjfEFHTAL
oAjI/iE3zTgD8WwgqT7BcIKxUfUCcjxYzx7Bx5dsJL7XmffD+fGvRu3cDMMzSXV1
dLkiT7/b+qv5l//yLW2T9V7Xzl3nIb+94Gh1vHjc28GGYwYqB+IW/RYV79rxAiOG
P5GiSkTHLWv/wHRtdNZ2HQD3ffj4Es64wR1+E4BwXnPZmIjqLODpB0JsM19ttrIR
OMfHUOvtLwhrpUFfNi+8Hh3540p+NLbZpj1Mbkhf1Ap9SKnhTQpSxf8O8WIrACNG
v8kHRXfWBsgCnLDzQ1NW3LzV5Qi7H+dwBk6SJcX1uMF6NucSGslWwj7r9KbTA8VM
f+HQvwc700mC/um3fAwJnX5Scu+YRi3lrfQaNeFUd0p9DIG76tX2U75YrzfycaPo
W0XmQrExTFqOf1ob6pXTLVquvY08sRtPXsy/tDzScu85zjwUZ3BZiwdtKQVZE8Qy
gi1/s3tb7vKQKfxn7Bh9f+7n/lo9tgTC2cbDv0JV/3SerzIckPqKhsVVi92zirB4
3X81dpCmqd7W0wWaT2hhyGAGsFJycBlFkYQBr/xsNrUHdXpTpeBCOnBnr+EzmP0w
Xl/BuAsBaTHcdyu1JplBSVdFRhaOPlmtiEjRpet8B0U2CNlUUBrwdNH/125EeRUe
iKi8EPR11XgtmYgFSFZ2ezguo29A4vYgsHfTFOVBd/Z+dqmGNjeINL4RCJDQvV1K
eIDrDsA+u7/z6lYZyNj2pEutSYzbPpup/uvq/RG6V7gjkgoSRqrOYSqkgoumW3CK
n4PoZWzBu5GbMkg0bOUxQDgeji7QqnqCkGM3Ezs8cM4waVPR6cbp1nbc2eLmyE4p
swmkZ1oQI3vyS+MT4mufOs/GI0ghU51mZOX6KegKCzyFjZR9Sehyk6fVMH+TsaJO
9RHrO42gqznAC4cHNMxUJNvI2ZxSIXUjF1Hv1Slhz1f89Kjx6w+OsrQRWTsU6pfi
Z0rVEr2eUrJyzg4TSuo9Bnw09MlLilu33AsOo6miiYSba+DVtpFSFd2cKmKruCoi
cqaNOh7KGTXjDOw139BW2prXtdLjFzCQp07/BZyPn3oYTfRrHSRP0bTaNtndi3OS
3r7HPTj1Q1HXk9gsVz8Crf5724Pt5uz0p5ltC0VIuAkrxJ06jIT/gxcufFbFcNI8
6IwXEg9347QEwiXzhZqc8xXmyKfz3V/GAHHXwezyn2Xx1UqMCNtmHHH25u9g6spf
6DzplAmx5HRvLCjVZmSfIPbU0BEydTJnQGFDjZFGq+mtKGUVhq50OLm3R4okUjQ7
F+sZ+9DOXiRGQLqwToZmX+3iQcZI/JDQexnFY/WeCxSHgC55W+HXR+rRWaTNPQA6
dTxKlE0syoTI48ip93x/GRWbgwc1CpO6AhKnVJ0KghWVG+mnJKl4G31L7dqUyTPi
XpOJ3zhglaH4AkBkp6rxwjJiH4CO7e5y7n3sNuMm78o7EVBInXqGmE/VPMCmyfm4
IM63uWMLcKFbtBM8RLtDNgkbNMni1HjiOhqH7tg7gOEZFsQQFEvaTamYT8vJmrft
PrabNIWko512fJeXil5zpv0bIPtS3y6YNjK+6xiIi/+DDW694csbHR9z+oZIv0jQ
LIFAEQIRufS6RWbIOaQSS+PSBdhxdAXPSt7b2zlifHDl1knjb+kg4i92Vcw6ZBA4
TtrwSQgAS0eFjquhpnGsN10pmeUcS7tgJBN1Beh13xEN0yNEZTibQ7VoHItqhWlK
5nmD87syNdOAp4BxPLXQVJOTRqOGnbSYvr3lx2/940S2ojQTvnSp5RhdukDEpbM8
/H5DCGdxyYkZgK3M04By/F2/bTr8AtaDu0fLcrfUyYwUcVHCLJ/7/a3hgmAjOMML
cJ6DzOD9ABKD+sS9xJXeAUXmfC+M2YHBuWdGsd8bp0+M1VmKFYgJildU/4bjrD+5
IwF3o3DNiagBjPDtiRsdGjzPdQlyn7mtUFLBB8jqk5Aob4cp3fAjoBDNIju2FXtS
y6X4XZiJzz4Xf9X10yx4mJN4qgiPqWoHKrvOR4J9DcKQZFbpTPnFFcneecYJX8eY
NBiFfAFGlutjFDgQQQ+h1Zw73AI763LiS7WIGSQp3jSMPYpHmjjcx7Vhfvj/rjCI
PgplEYvClh+toFNz+V3j68w1R8a/t/feFY8Dzhv8WjS9W8rd904WQH1oBNFXV2hE
CJ8H/70bVg7Frrzec6SDTOInTLOE8McP7Jr+N+ATiNQpFg+MCGMIY8b5leyhUEus
m8jP1XOMq76/c63qTL5Gs6qYFquN5z/2Uv1fM/99MQm80Ry6cEumuPdogxVdv0Ha
18WoqsHrsNsaKqFGBxcxceOyyyxNHguU0KbDvZlPqjoTiPSmLhJdCJZJm+3eisdA
APD0ExdhKLj5Z80tey1pdbw0K52Plr9YXet16TwelKJPD7fiQ6gF8+eJJyaDtxLd
urnDpf5l77NUNlgw2nYyt0T/Lncm2BobEZDhRzF9EDQpHAQOkvT/lGJhCAAXq1Bk
rBWbD+Axo4tiir+yQETfp+sDHqPtLQ3PjU9m70sf9Gy8Xi5JMrKrHI53fzXUCeu5
apTyIR8PTHgtjCcTQcGxj+LQ96RWkBfz87kIvbxcreIoHweABCjEftorLNoQw2ww
IJ3/Ja4jI5vvkzcK2wud0VpLsH2smKWkE0DcCGlImQoEGZYumMvWJkjeL6BLZiyL
6w4hN+dS2TLtC2GYp5+i9Wb+N5HqHRji0IyXLR4HFw013Jisv4t6y6AjbjElG/a6
j4EbyjL4QNqxHK4+Xm8tL9yzlKx888DvD5nJE5h8H+YF44Dk78dmGA6xgFoZNUmV
VRkokjtk//5EADB0YVKylBfvPTChVH+N7rjdculJ/vRTi/YyQ6MkuofdtuuZ9fsa
yc/8DuCJfEFhqtjB1B3ZgIj14RQY3HtJ2mptxnM9igk1VjbDeTiVh02IVt41cInk
UoUKoorctO0HXScJvLLGVeyy7+GW3h/VrRwTZlxDYuuWeqr1fxMQW3Ck676P0dcC
dgz1BFnhLD/JMHDMT4cHy0CsAtSe70WYdblwn8+AMXR+FyIcxIew+qc6pCLnjgcQ
aWEL3mRV5idoELRwKcKYYcLeaYgBBKX7YlaEBJ38EMs9h+14RzRV32a1ek9RmMlc
tNMjXjd23YMR6fKc137MAsHT4tugQ+g7iFJkS4O4G7phNgUw0KiXGVTyx7RowUla
dYc4/3KP7zl8GoNWBNDnhbpnpjp1evMyxlCyyimFGlhqFjJw+Qq7dgxF7qfRr8io
6/ygHZ2La1C+OA9OgyMM56jAMXtTc/QoABEdHNmWnxBko1hcT+tyieQBCOayMvnF
x5wYcIU7SlNUT3v51bZftBsiMgoagtgTMhSvQ0FuaMYSowQn1XwahrAmp7Gjzgu0
lOQ9wrmSE15sN2rnjztKeLo9j5vkIMUkJMofnDwWoIvICn0sfxTFcxJp6FtZrOEg
FDz2qIKlwzryZUItdLWcZPfKNVF4RjN/Ga08lGNRIVL+XrwlwC+6ckJl25M3hWTL
23+YKAxUypxpP8mD6n3hx7U56nm8qU1Sg/Zw1hZQdYa0ubcFYpvgy/dMa0dlQdzg
KQdgMIVol3s5NUw5fozJtKUh5tc6t9v7DmV1VuOK5Wf3Vd+r73xuYnMoDsxNjrnO
oEgIttumDHuN9oXKK7gjwHD/FE8FdWmR2O9HpLZPIW28gFLnIWJ95Kqvlzjhz7+C
z5AgRPvxQpo0ymcVWhbQv/mQIaPBmsmkQ1x1Puyuw0kkwvjG/kL6sWECFqBiQIRr
ODvoiCOa3OxY0dOUZiTfgiq0jmgMzC5OyGlhMYZguOR9UFl7t2MzLMXhPrv6+SUe
1VcDiE/e+1XB/gNADwsXFlil56BFJFWKHrn8jHQ8OHVon/TR5whtL2u9u0+2+bOi
cGaCeHz9s7FRheCoGvljMuyd3Kzmdilx15PtvZSqAgmijDHEGt2kgwlzqu+HjBoC
vmuvE4C4i1Wvic+YDGwRGzP27NQW08dzRm5WXC0cg7vUMQcsCLOqSKHOMG5/Wmc8
LikPi4EppM4dc20ZuY/3aUX7voZpgYJEj74r2OP4SEGZz8ALL/j2tO/x1sNTAD6+
tef8kNbmXVF2xetbqPdyjudtROPSxUQxE2Jp0Y+b1df56JuzmsoX6TtuI535ctlq
FwslQ3YT+JtvJWiYmKHLov2xiHwjmcslCEmTLz+R19a5e2rYpJJ0ViXCHfr9a4cG
eyWZUfhkHb2jYHCFzRjXxP2lSDsy3gttl6HrX7aRKBx8k3PxsapvRNYr5Tbhf2y2
f+11BjGAY1SZdlMxriqeELi2va8DQHWLZY/kP7M2xjJbUMCSSzwSyovhcT9wd3pI
CQOhG44VChpZbZR2MMxVeaYrJJzuX5ST5W7NhVuy1rCGgWnDIVLYMmVygXDVLXM9
v/GW4l3vNk7e3updf/+wvumsOvWnsVEhZh7V+tjB2EMp5BVXZXO9A4FCqUAfFcb8
NEYhQZYf+Iz0GEX20lwgMA9y85IyZLIYVhwyM32SbQiEHqsrAZ5mBtJVN6JS69dy
/o/5xE03st3EdSTJCGuG/v210qRbIamYsBPhkYoqfOhLG+IwmJtzDIqCDXoEcTBC
bCjudX/vRlzBToRb814nIpioCkyeGdlcG4kFuEOOHc8vdBc3BRFmjoU+cD/CrmZT
F07IBhM3yNy9LjJxBGa/8ueXG7YpfXwWvlCEpq5YlgYeOGWDcV13/VgPDVB78KgI
NvTx5bszbrKuswIgF+WH1EvBakCpyv3s6a8k5HzpdKro4drroX0jAdLryr7iD9AJ
yBf43Lb4740TcNRw2T9Y1wM0cNJHqYK0t1cr6MtG1LVIMiSk3cxhKhAfiPj280+X
7lS73tE9nVPyp7KE6py1pjzGNfiVrwBHOS5UT6sIH9PyFXplsM2AAxPnubOAVDhc
lciVv7y6w5J6EeZxlsl/SqT4UWWKC365+0y1q92+FPDrJVtEwIwxYarXOfUIfg8M
uzOKwpe7uf8EWKJ6dic3IrD8mrvcaTBoYMOfETNAmAacrMEy4ALYdOE1OWX//yfH
oyPesky4i/N99f1+7zc7WF1UpcAnz+fyiLvV0ZR/v34HQp1kE64c0VwCUQoboAqw
wzCwZoPYE33LIWyb3GtxbwBASylhScJvGhDxKnWpobsqBBxzruJj2Btez4l04B1L
9V260btjPv8ZwHQRIbhFi7tOyc46mRPSD7o8JSUyJI8NZPiHlmSQbdAOUWeIGF8S
ZGgRmiWr4c2WdCpxNedt9epmkNUfCV0lhPh/fAqFhfcuhBhT+ArYeXFedFIlMHf5
SHR3qGHnDFU7kOwIBU6ET8arZTXnGmpViuY4Ak1er7gjX1WCVM4c2CIn1qeWvXhK
etkvF4pb9ge1mftc5KC6lznluj5q/VXePIvnbhWHGSzcm/dtIZ4eLgh7/4Uh3acs
5kgfrmZJUrEcoHhsvtstEVtJZ52P872JJxiTUPu/KYdw7YFpQ2mZIg0RkuSZdvt+
XfFUhK9mPX0O9oywcoCt8hhAOSDAfihqXtq/+AngFA6NJl/XcrBQiTaM5olikgt5
rkEqbp7AnKLy9gw3IKQq579BEHet8B7wwY1L1aWeaCp7O18sE9W1zSy8nlQm43qy
t2UnKFoIyZ+Eg6BVEdaE9FOVYBOLZYYM3YsXDoySCbFvAwk6O3la+5/+NePe4s9z
9pv666MEkUdv+e/13tlGxVpJckO6AEglM+J2/SAXOnG6EU08BNZSZy5v6CGh2Jbw
dH87Z/N3oVw6UxnS2j2xKtjkOBS0nIbJ9ovnQvcLE/BX95p+8YbONzwoQOWsESwB
hnRbQo7/dyNQXZkKoVIFvySBIZ7iWMqrzximqt6sjIpJ7dgCwvtvw4RWFRphfv+H
Wv/VTfcn+RjsF2/o6Gu0SMVKehEU7E63O9W67qhuB6fYyrGfk8DwD2nTn7CSZ/JC
DUPksE51rAbp8uP9p+3oR/hSFEJhFOL2vYKC2vKZJfa9TeMfMV4mSfFzSkqey0MJ
89f+6wzJd1AkNu6RdJG7i2bdgs2Vzrj3MI1hQpnbk970/ln4oTDC78GLOmSj85/4
izlGNdjuvdmeRP5Ur/7Pj8mKhxnm27tk+lrGPWolsFbcuy/IjdttN0rFVrOGC0oD
dSy6K+7b387gpWFDVr7KNqxGp2SPQeIoWttAA3BnVbCYWL6/w8uD3tAhLxfzzEIS
MH+FwJRzF/uE87BDF0PkpRBC6s3kVEvB+bFBPL+5CFNdhnhxoUplvKvdnKUZO16L
swYOkR8cwC2Vai+1oFr1oZFIlYIUMyu38FNgbqNKSJhcbOQ21LkV391hDHDrUqlF
VS559N+dyNiTL8NnRcwqOyy6IkCxy5Xal5cqoLhEq/Y35s1Yl9MaN5vjbT4wm6jW
O8uAXMVWnaDKVp5ErJ7dpsxM/egGpZxXKn0sSxGgW6dyR6TLmlechPPi/h9XwyA3
blwZH0juElG9c4gHJjzzf2xAYDQCmnV4848LNgwsPAzoTQ+m+jWSLL9Gs+NdI0C/
+OuYoDHWUj43tNTvxoyLM1gwgWllpF/FeM43AvFvKFIfxAPOYoR2TvgyecXPVJB+
knC+yOrNLZs8CC/RSrsZbGeI7rOjlY14rCKp/mjW+W/omJC4MdQJm4QWO/zjqNGf
DAesShLJ+oX7JPXmB0HecmABQlR8vbEq6cQbklzZFw0jfIiwk1M2Csqb0P7owsB2
PI2kp0uG/TKsgD3Fa3Y7P9GR8ILg1yyaOh/5r7mYPzgy9M8GQ07dX9FDS7OxFO4m
NIWyoVBINkCKFQN+5blklJhsNLEvbQAG1fer4L/rBNPTAVS/CxSyEwrSDKAfW4He
uTtY67HzgYcogXygrzvZ/cp9UvDgUqdkC1iYI6FN0tX3Xpx0LEgw27MPR4mwKubX
e2uCfBxPR4a8bA1dtchLoa6xPvZjAN+9oww03KTUMOe6b2D2wdv79kn4ezGKaaD/
g9hAlzhpx5miPmHTxdE7gv6hDsBihy2M9emCG6OY8UVHOeO4VIKSHcZE03Xb4E1s
R6W/Xxw9sT4yqTSOKyoex0b4xdTQ7eUB866vZ7vIz8MaxJo8katt/6FyoC1DJSSs
018AFfePaSgdUbMkgEsVTTflRDXM2a/AY09vA84BvXBN3JCSJ7/zv0f288HJKnTx
VPomOf4q7QEQCIEecS4pb9h1vjmIE+AC0tGp22CPDp1cxr4RPYjGFCXp1wHsccIX
hBC2xMVbHkkUpbTGyAgrb5jWuMJFmrk5XTDp678MfApStaodf6RyxOR/xxlvLjn0
ZAZPYwjL4PUUW9XeRoAcTe7Y19dvGlCXTdC7NcYjmnbvcTVVixyymV5vUBH+CHbB
U0rUM3UOA2d8GPiks5Vevkt3fODQQ+pOFZ/A2u4LkA0vbbCGlv/qg5yXN/KuYrzd
A2T4lywBtLqSOTc9aVkU+TIBkyadaEUXWu+Ils4tzMKK/bSJSe03FNpCfAPQ2OJM
PaEgit0KKodNNdDi2WlaElHQbSdc9pVodS5S4B9Wk77fATc6VK4J3qD3YQVORju0
LukWuC0OFysRV5vIKGTCFaRM0/Yd/KXeZufUxEh3cHoxA2o8Nj9PcRcDFFSRNlgj
iO3KPD1bd1uyrvt/7dGxvf4Tg2v7Uq18sOBG3Th9DOxub9ZaQDMrdMb47/t4OWhZ
EcbLlYxdHtcEQ03LE0210qjr2pdSnvB5vlxtfUv810Gu0Oj+sm6txUhYDH5jXHtX
+2J2fOuSLIm8arW9LtNKfTmth12M2HLz8ZOhmn8/1yOSxqBFc5/MKw3VqrgpDVZQ
PTpYwDWOt5k55OcaQQp9Fy8qxkm5bF6Iw2WzyJw5X0iKmkPjJY9LN2KZJCRwMC5S
Yy8mQkyzr5kIygk9MY8UBcPzLUZ2nG58G3/1wMDHFBd5tg3FhP7OV/LGh9h4Gzxx
IWjsVY61HaxCErsnxiHfNd/Ll+oGxeIEZmUUFev7PIItLpsWIz+a8FiSbW6GcQdh
Cee74i2FCXF4qAPKXiqJen4zGspdA5YxOQTI6D4rbSRMxFtM6KfUCTZUZK8TtRgQ
/U2XcSnFQGGeyrFgyivKhVBfAI7fJ2KhlmE1JtSGPGP4LPSZEBnHx4Lkvh62CIKZ
oBpxmgyjl9Rcnv/xtLJ6YOkmd2glwpqNg5VJ4UInh4bh7NuVY4zCigW/Q5r8gND3
EUX4VDNP6lr2Xm0j65B0krW1eutqApE//hx9XDCiEz0UoGIkLckxDMdJqYUm0JHS
G2GUejrCxo0lVRnu20k6xRM5QuOOyK/1vFaZx/efcQK4INtLUU/g/TB1xaNKMmHh
1Z+rmex0XUJ/adg4Hd2ZZ+vk9hU5apfKxVZBj0/ByhMBe9KpFSxWwbgDBNdSl3z4
H2X3gkwo8kfWxCXO1nlAZNBqYq2v2NLKzaPD/TtZU7ihUQFN1gzdP3nCAq79HCrQ
aIZ1gEAIgxG605HOxEDKz3RfNp79XCf0KflZK/qqTWI4SdrQv6aeaVyH64DGoD89
Em+eBM2FpsWOAq1PmK6YS2HXDfLRSOAUfVefqqdDTk9IpwXdJO/BgKA1ILZQEV1p
ryUsP6FnjJngLmPlrUDWX7NaxEARxByc9QRX7UoyE3l8/eBc3c494O6D2CBYdS2d
kHKrRIUveWyk0S1m7N/vZSW9oLfVS3t/sr769gw+he3dZsxAFHt9uUykbVAq75Wg
ZjTZ4jFOb0tyLXo59wJvttJ8Ivlbpko3Ob+yO1wXU1KbZwdfMX7aVBwiWmng/seR
3VxfQWHfXrBls1ImLeuDfZvZw9z/qIHlLTbyeGGAu00RdZYXIlDYtnCuHo8WYdAg
K+rIOOhST+vg2jyCGe2ddFtr69se4F3Z0+zKlAnRGBuqOuAp8Znb7aQEsYMJBEZL
bdXC/sMTvXWGZndbO7MKgGvTLo5MmCkhNnf8wMwt+iCNepsB6Bn2Sje77lofHwbQ
9Yg6KWURJg/FouLx6tdtZ5MgyODla8bElWx9w2Y0+JuJIpWsW3fPTXNMBY7RDgkj
wFYvOWk0H4drGsxZxYL6ejK7x0+VtxTUNrMitB8Op4AfqHuzxHvqchNuFxpYhSwQ
F3P+U3cpIeENKN9QilDZqn4NMrkSCyW6FR/oE++26/DUH19/dA6FJ1cIJTqbjhkG
DYpzT6gcZLCmgA735RddpfbCGu/CTBGO6GF95/mWRgBsWfdkNRGGqCWSV1n7nTE6
RbBR1Mg965B6oZ3xD00t3G6VWUUzAHoTy/Y1t8xVeVtyib+VqlT6t0oMv5tNGpC6
NUaBGOvW/o3PlOiLUv8F7iTmeqXkZdhMQ/EzhNwjQ0fIDfy6dS+ozE9+4ItzWjj/
zerDdfY2DVwceIczrOdnxVcBQsSk0yk0B6tfcnaqoFvcIfEgeQyN5ngii5nAh28W
tXcN6ByfUSnEeP0kce50c9F+Dv0OJTSW985nZHL2x66glxl5aAjrDH6IHlwmLKA5
hUNtdxFWcnmo/TaSO1cHfgKY3Edh2Ap5EvqMoWgJwa7wcEDjWHPiC0Tdi37G8oxN
YhNOPqMQsGxtTJZkzxQMy2+UCPFcNrN518LnBoYA9fCwtfIM1jQ6zZL4hhvL9/NC
WTnWaejsx5I87nkPlX94wpPUJuPsK1yWhqHNCjB3aBxkOxHrukxsbYYh9KEdDNpU
Z4XB/Lh8qU67xUkPZB5q5I035M19YD7iGi2t1Eq3mYSVIdyyeA6pVmLLsUKQuo0N
jgyk1MEVc+gJTk/pEuIiq9nVdSxmKvDOoKS8TcZ4kFiUwYqBsKzor9ne+Ujr9v1d
KWqQ/ksmQWTotG5Ku3bguh+0wPpfU9UMULkWKLjbg7qUmghyO7SFOC+biBEobMVf
bHm3nsOjYHWFFyKav7C9iwpQAllRR5vhKm2iX7Yu8zLcg/nsUW8AhiFNPUEB4f1w
a3yOWt7+NqyASnx6SuvVUB+8AX8zWBYMAg/8AjAljYgtyj7RzN70otWdSvhO0Kgl
ISIlhcFEMLMO3xqOX5m+EqRqH22Es3CBmXAZEizFU+JChK3jWvau4lrRFq3XTEMl
T2unyDv//Y3cFY2aWplNULRHwPe+v1VA4jOSdrHC3FjQ/FJgX2QAUEEcN2GCN6CU
xbo8gi3z5RO9bclsfu2qnPedoqEGklcIdnVKI7SrI0lqdVzO/kSrdoIpzPuV3p3T
H91vYAmXnXwRHT/OLsWwx0IAVQfy3Q4ARAIG0YXeAnixPbvkuO1GW+NCJ0quqLMp
m3EA6pYo5/iNkfrKD2LiuZgZH0KCjf/3CGxqftgA/AzvvV3jxVZC5pSgTKfh0MUJ
4LbX2lAWdh5ry2SRVzSWjy3shetnTJyiWVYTuyo7f5c7yOd8b4bu0sV3TyS/Zu0x
mQlU6e6OTvDGKWTihUjSoJ55dJOSmXKmvVuFdaRgOPrmwnW+2+lnyonVboYM+ehZ
ki+qEfS8CTDoUiUEb24uwYv36pHVokk2pRHRGoCJzTB1VgcU4RyS2/lTHE4cstic
hCd312r4Fu/sZfjMwsCHl7X5dAcct+fr0qz8Fu+44yw8fwNqNL0SIjgwSfg7tc39
vmf/WN0FgYcyXASPPLbhbnbwZoxzgSQVIQpRZQm0V27P6P+xLOJgYTWau8lD9xoF
brdMUy02C4R1I53JFTfYyXVGF4YZl/Tk3f87F71q+fr4PpJFlVLfcKpQXkMfMWCs
SMAg2eiHngHG2IPi5ZLhJj/xj84Ic93vz9JDJST3Rcqm2x+HolUpVlG14109PImb
bJculwZlut0GwWkciYYRkDg5JsGh+fWk6azl6K7MBmAtt4IXgAytJaaFshhJizCm
nwhX416EB4CkNOMY/jVUcv9e3B1RGkRLJ3QUV0KD6WW5/CKccDrkT6iHwh/rUCiW
ImWSwEHKGY7PXR/fI8PIfMzmOg8ldpxG5gsQAGWidA9anEAE+Y0fVnGQxA0LEKF+
jdura2uQb37OgP+8SbqkJnMvGAGXgvkQMUG4zBXWAARh3nf7v3Ea2rhajJoUiFmg
wxdrwZQEEeVBIptbzDsWnlZBooo+fX2I/qccBgHdezFm01kyUYX9bCLnggaJG0bV
CSVCSENiKl5ru2pQ1rRkAzrNd+vBZa5R9VMKDOuIAlgDcm+1dyH1LGzumJfohl5U
PhtTRpLACVOZz0Ae+MGfYQ/lfpgZLTUduN4W/o/KXjrImlM4YcDZFO3sSZdtEIqh
qjXfkwwrqJNfFMhS+rIs7jlPnkPSzdodfV9HBHS8GQeu52w8nwcOU+8nOX6pj6EX
9oBDXVqWwyJpcEJoLvtQnjU9aAveADoC/YchCdDbqgIZ83cjafeQSxI3wtleE6Mo
J+zTPKOQAedjU0EOq0/chUUAJ2Upi8yo4y4SBLMWpxTWQd1474+ROindtk2OcUCS
oy/+GDqgFrWYfDMNBG1txFXJx5i/ik5q4fJ/vlCCJDfXJzZryoRk28DxtbFtOw7g
btfKbDKqFtQvsjiSQCNUvh8pxNMqinnRWEmK1NkgzqeAMwa3YnsQOkJBwyRJFjj+
0013Xyqc5fXPZ/KaXuvOXy3S2BXE5hFnlqGhLEU4LEoZ+D5WFa0W0TPNeq2IKj8F
tNHkyhsEM4sUcO7nBacSsI+HvSS+U2R7TIRgJ3NdAEq0P4cExG0MFJGrm7SsGsjg
lkExOV+76hCi5HSYq1PnLQrWoc8P7zi9iAhTt+PG49gXpDybOSROceF5GGOYf+cc
9A+ICpmC7PF2vu2AN4kuK8gyjA66bIgpGrN1Ix0EINIxWFT5CFAjq4cYi6Sp+Cbv
F83w6EX+tlME+dFc4RxwPkb5i6eCcgRkoONL19b9NLFjNs/erRmAr8mcNaXMSgxC
UW9+RGokGab+FS+ImdsfSqKOZqJTlqYxygEnTEa0GxPs7yDz8na1titOBhqTX8cy
jSCtXWT8Gqswy/VN/fyaH9kiGqiMfCZLqkGLOYzkfYw8DjiJwX8q7ylx5S/IgdwU
6s8j5XdX/ZGQkiIY45Y8b6Tt20qE30SIVkcAVhI/A4+5tp+DFk8TZevpkRq1lwR8
p8L4i230jHJ1yuf7bpubPLOnQgxkMRW+uUDv2pC5IcTjBnyZ24UdA4yZdFz21gbX
aYjcknhWeIdO+vGYZpfCDFS4oucLCx0FF0T/w4dDUb2BsFU7Zz5y6+G1jJnAx2Hv
z6IYil9cNUbfGc7l4NXufT34FzAl8xtWEH3RvHgt+aJohiRMiTyhyLruz6fLwHlD
lINwLTqzbzUdVWGtTg0QZxDvO4WGbFh7NA9LBLRNPrOBkxy4pzNJ6yToIOVpHfWU
OtUNnjVWuVOBCx02ZHrvxeqayFWcUVk7CflvTDh2dXbO67nQFS+XwcNK+l/jiReM
ICCQ8C2AWFTvE5B1rGuEl9ck8XeuCfGARCSHaRKp8NcZ4TafBnoWlJb1e/M1g8AH
xLANnHyKcJgfFjHUxaT/0pVRrmHRNdkw/uX1eJsCEF0HC97LDWC+vdjoPNPDxIFq
uG82uV4gfRYgFSw7CHy7SvM4Lcd+LKI171zAd9jbc3bxsLSmUg7PFRIq6B+Ybqid
p9XT8/pf7VtEFj20p2QMY+h8KXod8uNz/AwyfsX/LXB835ny7IGwrcovzpseqDDZ
9ZH+wmfgwLNctLQm9LRz4RH8VpRfsw9pg2f8d2aHZgAxLWOIq3LFT3lY4+Yp8ARf
RO4rl1MNtK+py6eBHqVFLDgAs1MHgam239MM/gkTs+c2Sifq+fQa0BlgZlCu/8Y9
RbMcGECueWz7X/mSEblgYIMxntq+FFdVtA7P0h8AWpS5bVa0rck21KQXwBwOOXLe
YcCnASMAqOnVuIQ9a03FbNVd3pF5SfBlaANZEv9/kgoE10Dsdv8R/5C0Vgti+nmT
h54aJH6L0We93SoZ54GlJNQ7MtnQn/w++qLA/6INQHYxS7f3R8iPwc8ZHH22MyQ9
m15/qMTGIxUYHQia8I8jcxSIFhi8ip1I6NhaJE3pxDKrQtgLPcNFJd5y+ZgKtLAe
wYJp4qEjeZvFnugHc6KpWaLbON77W3y6kpTdHEl2/UFcNjSllzW51lNUr19h0ZLg
ZlpvJ6Gb8ilMoEyG3PgFIc1f58I9Rt99zpo0jWC0Ol9PV+KR2/AQBw2mU/5KNL0z
2Kq0XvPrumcuoI5UoWESWHRfs2hyqhtNgMqVETVlnq2vp5AdQHjPC1kePJqtUmH8
cvm+cWj/HoLtrt2oRq8dEBOcME0yymHHe7MJmq3OBFVGwCxx70iNcnWo6Zz6fyMc
SjUs1lCm1qXajUiUQrnDNDt8tEjl+qKjM9lSgLva4OUR26XuTy7DBDWIAqaC86Il
IOjFgxg9sVWWss2gv8b8Z84T+yuZ3DlkmCl2x1r3jE/0ugerf3ULR8ZWzQvrcTAX
NbGFRen4nOcY6mbmzZHFCnMZe4/XZV5k8PnkGXEhDwKTFu0x79ISnuIHMLdJS2VX
D4f/cbMRddZyS8ohS5yTDHuXzewqRBN+Vn6KITR5KgYxUnAQgMHxVLCmE1dko20d
Of6N8YJcL1B4pfqVeBlapx3FbRZPKVcq8OoPBtLPkHVBjzczv3a4zJA7xkwOVY4o
zRxMNrZ8t0s4RfxpEbmheDadn4T03WiaPHEG77lX3j5LGUOC6lNIVM2CST7Y22lK
9ygZS+RwbtWxA29VXIyVpYArI5ifMs/uQdqronot2oKQKcHb9BbHOWidPPi9Qjt5
GAffxhgsJ8DsMpPZddSopfV2Aj4iCCA9VKpUH9OxepvwiZip1bRqbwQkPUBwWmBP
y9fb8jh6T+xG/eGuWeje9EnntFunFimdFjcg16I3IoCgnUQO1q1+Ey66NJ4U4SiW
JaJwpwzufNRZRKgxKhEcuzo2fgsnmTH4cqXASHg/6zYziXcvVSMJUDBS0GEUZpgq
16PmJRjPSQEUtOswvK+2UoXwYAGQ209TZEjSu+9Gr3ai8L0dqdrcrtuwKHyBPUCM
bKjegzahtn+Y7IbH9Barxh6O/m+LbWI9UuUJ51cnTteXo2Ck9U5akNukCcQO9PHn
yZtzmw/w3a4vh+jr4krav63ibj1xojs5kZIC647c10fqahIDFJtH1r3VQWHkvkP7
z7cjn3iUASZv143rvFSQZmr6XbON++LX+MpO930PgIshxGg3wwPGjE+6t65W7j+o
S5wGCAHZzo6Yc+0LSUq+ndvRyDmgfOEo5na1h9KOsyVtusmYKVcUG7gagax0cj/7
ucifyyzlcBT0Dud6K1oiMrXlyXmzor0WIOXPgxyRzn789URhr0DaU5EKCjyJzdPK
2pZP58O3IuAes41x5BLhBAJFZL2DmOpYjpu+vqDLm3+5Hny68dkRHnREp6k08HDN
9X3Edau8lL4RzOv/ulqJpwrizE2XtkJI7MOS/FCYBHAi0FOwWpU0U01vj3gt5vwx
KmHSsmw1sJjE1+QWxidm2v2DQ6rNWcXisfH4IlnlTJ8alyIN5n+FoyzFlqtlaH4s
FxsdcX7jY8RBv9orzMGFwyq9S0SKIigmw0xhuATTFIeDIylmC7kE4CCP+DIzouWb
iz4MrTXDRfrsGxkP24shpq2yYvy5mWOLFd0949+wnjPhKY7BjsqUNeb59UKu3Hf9
c3+V4+by8AqF9RqcjHVuBI2v4MSIZIPx5NuW8jbHXO5j4vL4STfrfBQMMeH5LOH9
R3FFpJAcdYP2N2rr1SxnITBoxOzkCzcF0H0iDo7lfrTUGL7phqr5TdY7qcEMfVB1
V0EK9YP0VK66PKGfhSWQHoaFNtUAUMZTqDb4lrt2LUvUyF6lZ9/KUqdRQ/xiiA9J
xiKJfAuJGIZN5c3uJ4zFXAaz5IlScyQzWMOMgwxDqMOsEu6mmxgeadjPyM5VcezC
p9moSYBnojC9IL+tMob5J/agOG4EatopgGjffaIzAMxho7NPJwAsPaKY2PrPHpBv
JtRCTxgM4B9ieHYORpx3ZUK+qiLmYAXxhkOtpG6KRbtf5Yk5UkW6iEnzGjh3rmfT
yKEmvGoq65IW7BuerDEPZNukHvTNmuYz+6Cc/gvFewrwSdYXO0uakIZP9iEIfdr9
Ej+BGGqPNefvCeBXITqMxPp3JGGr1DuSXmTKZgEQHbPvErgDjDsb2e5po0Bt4/1M
QK2+oRsb+HHPfrar52yBqj4fkQLGyLsAj9RFxcsbpcM8+w1HpnxL+QlRGsk4ym8g
x1DgfN8eXaWZpb49vhNtBinK4QWw2g2g1BUsabqOsfeRQwjEkBJ0lt47+DelYxCf
Tc0LO0kmseKxuUT6/ZRtE4M5vRowx+y0uGSEctrARH+pClDnAhWPqDXJNs1wPLnx
bXnuow7LQpMVGlJ0w/ELU9YVLip+ypWV6tCoIUkXVaEZknFT30u05mqTZGWBtXoN
kIyZi/t61eLKWktm1kVDxbkaojt3HiE6/5vsW9qDW+c1ecyleob6fYq+gjCHGBFn
fGZpewsrCi5JLccJ+pZRikk4VJK9AMLNaXKzq2lZssUYag/XF4mt6ztuuMTLqHRP
CueAe4bB3rIT5WvoPXSo6kKXKwHknk8imJOkhppWSFrVkheKXhVFHWZjmJ7EqKy6
NXak8fK/Pxf23bpqq2S2w9pq+nMVz8LMJgXGZLe0uJ/yrl/2OFEbrKeAHVwtvZ4A
bqHeBPYlTfMXVURg2OeDpjpvmC/4lVz+BPVnV3utVFOhFLbYSqw0j+rPpmbp9sD9
rQCvlBSjx6gQdLN7jG4Cy6wv5bQivSXWbaKMBrdqsAzHIWztV+uztGyvbZOfjwx8
xI7jTG/0YA1yHmGfK8QqDLrhT9Xne3UNZioV6HI8pSrP+nuhFB7g3thviF+VfIq+
1QWpSgvHtwYraKF+7UOzdXaurC3xyb5zqX6F2P9RGiWQTI+o8agbHny/XZw+MY3Z
H0zu70fsJcwNc40zMYLJYRnsx5mMYHDuNmHpgGc+aVCJdop7VJU5ox74R6jndQEK
8G9UUqiK6ieeGnsOEQuJtY1zV9ZohDEcXQPrLFQObQY0+4/6lzgAoAxWVcas2v7g
logRg76O+OHoPzD8pIxKsgUBZC/UEW/U35niqD/YkxMa/CaYDTi0lStMVEDSy1d4
lbwUeZoYekuR2bZWxLgnaDDJmtnCBkwDHlKDptncBz5rJiqdr9FFCQCzAEGTFZhr
lsEjIdCcvj1yYPAY4P//V1gGfJJ/c54CzPcG35heXejTsW0z74259gAOTXCzQSVq
8FnJhNuVAdYe8GOHsE6JsL9aSv716UaLZ0xt4iinAbk4hyNV/nwoQ+1huz/75+Xf
hbPs1KlhVLaGSuPpfg7ylWRV5k+uenH6/nUcp+jhmX2V4pwtpaQ4yfc/9/WcWo+K
aCw70jGgYoMOWAEED9b+qM9kjR1YF1bIqYRwZO+BglG3QHNI3SnhjwDgfQHMrOHb
08pGWIcej7CROP28htCTpH11AV4y6mzJ511kZ35AMzTReIOixbVyZvzNg6sbG8Pa
FCuS2HdKzA54TuChwKtS9sNm0v1ltuItyBrNgK++NcCF/r8sQGepy4jgVo1sRBUH
fULlYxcak2kxRkUvBo89QZJxIbYDTr9Rej+oPmKmaZeB6XvOAAMZWT47t6YjX1UF
riKT4k7bPYjB4JYchPlt14m1ovxwYrJrFE5bsOnLAN1Qmj1dQnzNjUvfnk6Tokf/
qnrpy64IydIOtigYEzA4RxGWlkPTlT5S1tup/nBzU/goUHDXqCDdqMMs4eRQFoYq
u8X1HYGWDyTwI+mHbwTqEoD6gWVUZdyP67YZz1dI0Y72IB5YJTAGkt1ue8ura/Dg
qX7BLJEvT4beFlrwVi5R8OJGdOsVLlUisPgijgG2Tqu+SHLxV9033DqSBiasV89A
csqQ/eP234UdsnuzDlOv0AI5KVJqr8ngANA3H1pWjAQfuXIeWMjica2E9BmTpuvq
f6jf6xIzMwcda26SsO0s5NIjGCuJH7RBH74wmxk8akbhzbcMksER27OiTMdwJMwE
k+eopTRlMaXHVstfi8fv98yubbIKLgucWwyFaRrEBXxcZy6Kab5Tg4kV+FB5k22w
tH5Ks4lWhDwjwhP/0R84fJQlJ6+6za68O2JJMJPyiEmXsOUdFRfJvnUmh1C57QX4
UUplXX571MfACirQ7WijyKa+/2NaOjOpkKlq2xXSBMd1eeReGmcpEmorOP1SZWUJ
bCmBEuUhnNJZ83WhI5d3KTbx48SgWs2gPcia5Yz3l4Hd2xGHgUHKjZ1ibCLvQ2Xa
2lL3YiTlamCHwjYl/GOlYZIsGBxQu/+0qJVeShcnQeGv9vxD0yP8wVMtRpRyaggD
36qWUQtakrbF6kOQAB1T0s6Arst3wxSvu1d8Az4HKGVwS4ufrreEe+52QTvOBPx7
0HS3CY0h5X7hKF9scjutMssp6fmeyBWcvDmWO0nHf/lCEcqwBi0mv59y+oUE9xW6
q9JompKNZ9paJ4/kDE9B57/TE1S1Cl4YnlbUp6enu1VvFD6bv3sw8SXFpb9JXDtq
0vwgb0Q5PKfyVd9gsMAX8oOtZGbsmzu78mlgOwsb7E7hJX8tYEozepek386CZoTd
gjMeT6tiqW4iThFFtxuJ5W7fKvn1Q6jdwEP/3/tw+DYLd/594EFmkmjGKKHdSnEh
fEoVBG5OQe3F/4iTEYaRR7IfS2BtQqP6uo1MvIru0fpt9zH5/dPkyih9TmRLhOLg
cmn86T/BtG2oqOQ8ag0CsPFmBF66qgr4qFLLkxWDT0dGP//tLxKBlric0ro6iHQz
7hof36IjLa0QxR+9bD1oKXXzWhY2rzynlX72yz8yncoqSx3plxgibRZ4D9sMHZOI
vXVleWjEQ8ncR5fmf9+6rzW/bp2B1zw+YHHyWehaVgRIEvlv6O+xon7gSa6Mj7jf
D92jamMa9Q7EJSUrIIaCLqzWf8qyGzQ3DilapEZLUfcDJ/hXHf7ix6KbISnmZZ7R
9ogLvOIjbgPcGC9kjOjvk8EBeTj4ZA0pGq2Xi3wP6UlIcHTIrGA2E+y2iFZB4SBF
7IOxE8s7AT7ffl9JA3EkjejcuWg0+ZfBbIDJg67Qmp8nBcGYVIXv4SVVwo7a1Bgw
O8TKMIzWix9srAr0o0/JpJHeTGVpJCyi0LIu029hjcWnPA8YeBuBwGVTLR7dm5u8
hoH8d3CjrKSCXcvm2R/p3oMLne6MhtSJiUCCS0DHzzFgdqaqpxlQNFTgHD3fKgs8
+EGF3S+xR8yFWUcknp/NKBrjf7LXW9JERQgbvjozmm2MhHVDjs7dC+qwS2JMQQfj
pCc79CP+8MKxWpyRiU7vX1J+ycO/3xvcpG1RaF8TF0A9cWQqv7nF1w8N9il3lKY2
SrMJQNNAh3Pz9oSBp4aX4L9uP6ANCzEE5Yvlh9oTDqDoQdI3G8vE1xniNQw3CtXv
FPKQRyXGOc23XMYUQ+yiVAieGBBpCJ+E+dNGXKmYEAa6ISje5Xwz+CJHXrzeYNsO
fEtMO76SzwJuWffjoX/Ddfjzoj6wO+i0UNDYWkS+JvjLgi7JEcv6Pb2MG6muiYkG
s2SrGDpP0Zwabk4V97EzL6oL2bJM16zC5rGtVPMw/MGdjos5XFPDrMliIvrmqq0C
nTiPmRK3BaWAhV0ZgFG1p4KdFTLcyr//SxgElimblpXuoRTI+VYjjxhGGfUta3oy
C7tfSaqduPjTSHCCSsAi1k63vtEx0NevqYgVPW4uMqcMDUTdBo6VTZnJXb8KMq65
0CaZ3yu9YppPmSB6V6tD6PpoaLOrY0HXx0TGKWd4QgfNj+FnnOFc0uxRNORt0RIN
uGuD9Iga6KivN+oK49IwhTJ7Br1LbHi+LPAbO9VSipgrcBlEsA1LGKg0ZiN9+kdm
Ouid1iY+aReRwWzzTRWP/S7oj9FNSV4E/D8b7dfY/ymiuOLBYG21KNDaWJ76v3wW
lr4xjIhUUaB/ZcazQxhGxcd50SGoos+3PiuaWR6zFZX60uiQ9prkcCsqCFM5Xsn2
t5Iwow2MzzqUt8MoxsqDFuET5ASqmHfvFhLvyvzFHPFnqEISDVaQVfVq8m/Wpj9w
8f5Dy6YbEHIqRKZNGLYdkJUGfRwuDkYvJVv4oYUYuzTsur/X4KSYlv8PKqclTh1i
PvONgt3aktvfhZwbWYzNQozVd7htCjgnbUxDVajxblWo5qe+ApvXGD+npUrCCDmk
F+na2awnLC683FjOTuN4KqgQXTOc1Io9LN0b33AJAH5ZtjuM+K7BLbKpDx4zbXtt
i8DswTgQ9tUI2dYizuOC/eQy4mCrq+Yq3gY0fLv1u6H4zfzIZ2lJ0XS2d9ETTQ4V
dyrUnlqE35YkSVlY+AVKPDgk6QemQzumuflM3ndnhEen0TooclR4VkINxyhH8UGT
hVcjQWSfZu3nYWjkAt/kJzcGaB6lbrBo2hRxslrhQLY9iodECMuZ46Xyn7N4u/Tz
WgV8srBmVaosemSoNl5T+eoS+Jb/AYEdtX44CGDji+VWtg2mJ1siSt2arJyNtzzx
IZuSHBZ8PV777ecmWGE2YMHibTHRbmOxbmKvZ28y8EcZO4wkjMlPrOYnu0cn4A58
jyxsxZMgz0Cdum3xAiNmTH08KP7oioHyWz+XX02S5S1r8/c+FUrnWlFG4k6SmfAE
bfiJJK2XU0EGgjoc2p5c6VpdxTEbF6D8aJ4ka3JxAFOBWor8vVH1bEmaIadlKB25
QcN+Xnip4G2lOJGZmy+ze51Avex8liTJj+zGxZNxH21DdCg7UXgRDFT4FfRLB3l3
LBZn1SgPwjRTtl+tkpKNhPXZuLJow1BfSSEdWPfxePMvcoDFck3VoSal+X0JWzK6
LtVsi3UW4DApS9Cpyb1+4IqZ2b4Vn83dx+C+Eu4lh5kIKMShkw/daSZNkfNkXV+d
Hmcx57wUemxbDD/0yLhIp+ACR+te5AYyzuigrewpy40LTOfX7qSGhy1jHsFUl7nv
PIx2qlK+vtAJczB1v4Ov5lTWD0jYBvwayO8ApNwNEEINe56tVfp6o/eGSoid0agj
nfmO+6WMh2xWOiC21rTsXAwrZtDYt5MheacPYJefUzvVuBvhJyfoUzDs3gLf6Jfl
hgVkjHysgxd1pF77Cz/lXV9ZxQbgO55jVw3Qkhi9zdH4QVRdvrHZbRrHARsz/cDX
daUmhl37VMdTOYyfARFZzZTHZmFGOAVsUtiyEQHmZmwTzMBgFKKM9ZNpAvs+sZC8
kG7LQwhrwm3BFHOUXaO6mDK8nZ+Ms2Nu/3mb0gc7NnNqDLjHaaiaY0KusWRZ+YXn
cnXvfqxP0yH4+Hy6jfi1xhNjFzFulb26+0bDgUvwx7/wkqfch3ya1dGaS9fUMDZW
IueFlmR5QFn+8KX+3m0o0DyxWg2HN+QBcvgFFDAjWy0P0nUcUSvdzU+Sntid5+e0
c4AuQy0llvZUyCyVJJ7MI6eoKAjVcWaR6jHR1ONN7gnK3m7yhNFNJRyYAUJXyZGp
PO2hI7hMiLJazOAjH4r+CSS354kCt5PyRvYrHIHVTpyQHgjP0zMrVGaR28BKLv+w
PtARXFfC2DsnNgvcZRH24hzBEprTKkfpRt4xXKjZqYaX9eDF2s5cdLugggkiD8D0
2tu95ovGsodnsQfTcyswYzpVEZHv2Z16zwTHxvR+O789uh1JawyzWw7cWk7FLW+k
Sn+ssIjGh4WUnARr8pRoOD0xUz7kROTydt1BWDD4LdjFZhGWNqULk6ljJ1/GKZRL
lT5NQgdYcNcIliPuaMgzvP8ECbEq28rilflfE6lYx5poWfmM+bTgEkZVwgiHhkf/
7H5WNE3l94e2h8XybKISAni/0SzLgItsy61dUmWmQDMhP+axmwuPCRgLvniVoxJO
NLjccUPtIf1i+DlnpNK4/36eQTlG8LcxxT/RDgxnL38WsLDViDb+UrzCOtqvkvAp
Q66+uSClUaJIv/jH99vup710t0ztnabqGFUwD+w6GB+5CdT8LNKY+EcQ3twgelAS
AoHaEiq4QKbw7M3LcPIIJ5haGu1CkrqQ8b/vwXIHZGMyPHqu88NPgoU1OY+0OyCT
K38aLpCWNVWyqAoSwywIiOW/Bi8GrMuLDZnJKNs/oS1WYdTcFc+osofGO52NdxBX
rsuYYpsuRoFRp6+8Pg17Otg17oxtTl0oIBb6kx/1hxs5Ok6TJZkKYR5Kdbzx0sUb
q2aRI9D6N76iX+3LVX60TWfn/14/9YE1XmNYEBB0735ce+Xr65fkZlTGJbYylNgS
Q6qkviG3KFQQ1Ay/1sIMS9KB2+dZo4pyN2r2Xy8RfvPuW+HEPorlp1oKQk5eWUv+
RtnJLTsjO/1wOSUMhlBfoVgjDtQHHNmA4Kiv7YpDYiC3iCVCoaUOeq/j8rjqgsyC
Z8xFzLBttL3hybVKNAHfkj0hllDHfUq/GVE9O83y+ZqfHeeBeRdwFzG0MHruIcfK
85lF8SrCstYJ7FPbvTzQDaVZ8F4ZZPhIp/blVvGdGkkX4ScDJG23tqrEUCSgGNfZ
Lrsb5t8HkKgMiHUitWg0V9VNIfvXB9UhvEILABAsArt54sL2Rxka1Txq5alE2/5c
dJ9oEr3uF9CzPUdmVEayuhKWzNOI/rYyo3mjgugedjClRdezSa2IOyoO8Zg2QjJO
iwc6rb3Da2MtZnQu6/u6Fpigj7C7yLB6/aKZwyP7ML3Qd9L+9WPJDIXtz96G8UO8
2khIB0dDN37gegFKglVSVbssNvclGuZ/gKNN7HvdCttcvV3jF5eRP836sOO3mzMz
4rgewufnbtUoEOTN7hpXij/v6gsQWEQGrUyuQJqBflmSb29TCBZXJM24om0Ct1qG
EDnV/mVgpBmmr7hPRWdf2Nt/4gP7Y1K/ukKXlIxW1iOWJrxrwEAWD4fEi8XqttSo
pUlDJtD3f9TQgVLcACwy+M7FdsEwAxqduELYACE5HWZrs4qICXD6d9JmHplLeB1c
DUfYmfiFoj7/uxv5sTi7xX2H9zGtl8UoI6E336N7Ip14/W2EwLVisr3s5ojw7ZUc
ZCKGq5cPcTAK4xS8AGS0QsLD8Sr8UKSV7qcHGDi93zdjuKxUb315h2JVXJIvfKb0
NyxIdfZsIqlMjiW2mVbvKXJXM+MO52CXg9uxyvN1kGYylwZj+hylVqiwjqzGxety
oC3FQDKRFE6H390D3y4pz8gAZ5oCbtzy9+7TSTXur6ulrZxYtwXthq3OKxICQZDL
4alGd5RTLhJUEkbU68KlZm18DIFTEDuz4B459rkWkxdV3duZJXYgDLI03NiM5fOG
KJc4WZMj3+m6EIRHgTbTEOLGLdpZrjLudhuGg/2mwNwvb0JyhXUmlmDbWJdovQkh
H+Wj+SzhNU1D8qGuKxnW/1/9Qgqx4h4PGglBaj7R2kUKx8vZmZQ8ZTgjaR5x5+3F
uqNoFxbEWWK+k0XA5jU4mnm133tCYE7t6BXLqlLbl3FEK5yj2TP5p2/Wx8JSaX2c
WeBV5vkcNYSqjbJjrrLiReNogHotH281NX8bi07/9Z2yjps8vU+42AI49egSak67
Bhpf8UodNbRjKu78hhKhdh1MKjkw4Pj8mrdJXKl6IGW6jqZQsdvFGAW/I6hh6U1T
WDkJXSgaMV5t2PCwO82HdKApAK/gScQAceqf5pXxeC3pZ0ezUNVbJbYdxtK9NfP2
l9srjijyfw1jdCZOUYNHJtwoFRXzVYErV2M+jm/6SROacsDHGstLXGnjpTQLJwyA
uzcgw3fDFmkKBsIQa9et+/8xvQckx5/eFPXSM3oUERNiX5kReiMU9WR6O6q3SzZQ
9meyZgnBCpJFRCi95v37ipMrGr9pYlc/4y1oZq3rAFuRwCu7+L+blLPGPkv1CwD0
cICWP+hrVnZBcOC95JCcJJLukSLyMS6DwaP2XGps6mtDufBPr9IR3WjMSrYlRaA5
ZtGoSaXZfZLAe6eVQ+IxR00LsIJw3XgotzQ3ko1oP0QidOgj4X0q9RAvNDCSWvCC
3E8ziDWQvJamR7B5vux12bDX87DkewjxSIZgXKaexIH7oYmGxuX3M/7FSMaTTG8M
rcAtXP2+AIxBQstWlbKAVKO0hmcqIwr6YfUEwCPjaBPEzT/0a/7qaocvsBHYaAFy
yw5geo/kTKMuams3c2AY3zVrhZcCHHbZwTL0TKZ/amekcF8VBs0w60LN1v3NZfKs
KmCfJnP489t90o0MXktABpAszRj0vmFmQzo90a5URtYGa/Z3zESIIKQCzS0AMS1q
p2epNFJNNm62djtDJ/woFjDxqsSHq8HRkduUgq9f7bcVjYG6aFB10qI2TTwxXb9f
i9UqFq02bRFzWwbPFfBDfcjELiLTZSj/eHlbjdMp9/4Ntmu3pa42dwD56UT1n7+P
OC/osVcZAd/RyGCKH5ErXlkOO4RBQQmdW7IOFNH1ea8qX2Y9H3717R94+SKemXfe
6Mcwig6dCciYibj0syxcYarNiJktlMmZlxeXtq1fTu67yfG6KUknJVR8HDNNwNfp
6iM3was3oQpYU0P3UqVPQBf8ojcZESBbP4iUO4VCfYZCQ2t91CDlI4RswmzI+zFr
SgQy5MxjKVVzXE3s0xbJx9X2yGBF6qD5sBKF8+x+6C1uGPWuKS33WOCFmRnnzLeu
k4qhqLXbV1g8MKe9DiJ9fQ+TZEm8HZfgXW98isJZzN83l7kxY3jbEb7N4RfU/Snb
csYxOQdViB+TcuwgzRT99f/Msco1CYcWfTlLu6fimXFL/7QePU4Y4++G1jsUagG/
Ih+RKr97WCHyFpiRkIBvjtG/pxKfzvDsyg4CStM0bjJkOuVWCHynsTmXCnnLYJB/
l/F3F7I/L7sHQkYHLRWZC6R/CmduoFlheclBI0vWfIia4DsaiOqHryMJcrXqcP+e
mdF8NDB7p6VwVLfwpHDWFqpqEBwhZzxJ1xo+eR2nKAa6dz09BWXJr5f308cWr66A
u6Wv+GoQXu8XI5CRldYBPuQKQqIm9F1FRyAYwXJcWLx79AGUofgoszTI2OPpYhBf
/fic/3GDIgOYBGH26wdtk9xCnGwvY5V0dLuzoX9OMrRqaV+JgoBQMnynFcurh/M2
cjCdPQNq3jWa25kQkBhLhZ+DxOp70AWFjbJKYiuRPM4W/AL0H6omgCGCNMT/qqBG
QwB4CE90Zly273KuaSlO14FypBfuZ6MU3EWSGsi6CjuIyOXvF8g9vgmLbqN/yHkr
dX/nniMKjzyJKdfIQX17mSeKzdIb5ZapigOAEca3WKgb+fPmnM3UiGIe5INFSvWa
XA8nJojGCfXef+zBDhay5I473LFs8zSdJP5Iqb72wutZtXyzzFkPPXFWj5YnPTZO
neWBzm+JRG7reAGzzofRzvJXeiFR26yLjTnd167U7z2k15QIs/R399WfN/0uFwJK
lLSYacCF5m6gWlgsiYFE7t/CYBtdWVQ8/TE7gP1jSL1x30b9BL32n6JWNUfx+j05
W/I43iQxpLUsIhxPpjKI8lY5D/wfC3mO+Tlzy1TMWbpW2ZoJgYNKWCQv0ac36t9p
qYvvjOpse2p8e4QVqOp0pwhijcbRyR11XbxIhHo4knvBdZwOCnOsp3PPWhoR78Y2
qnhSxuE0nrSV+Mm2mqO3f3ZjBKJ0jYF5Xh9eIWF98mTPx8RtxTnMpPgn3tS0Z7z+
e0Mg3qR+JefJmXE18lCuTwpCe2qTyq7JGYxsdqrzQZIlIxyhuTOa6j0FpHzbCTIf
XGpVnJWzgMzPrentoaJ8wAKZzEsc7toCT4tDrhucb3TsQisBLjK0+dw649Vh8sYj
nF/UBESwq5dmzBzFiXKpe2kaVY1nTzOSxRWN43lbdbf/fwJypMiY4LM4jzb6Lfz1
4jk7EPhVNRROv8TVVCcMCJAruMG6jLO24dB06UoVNzUXPF/dSOmB6dtVunTQTBcf
I5DsfZwQ62vbRFlc/CZRV88zFodjPQ5rPBchexyBcJnSNtbGGNYg9FL1hs5JceIT
9yMnx2LTEuS612HbC3ftERUYnMulOSxbjYFrfCGEjwOF+byqhtDRzXDOh77S7/C1
mSmoUmSnTia5Pg0lqRBxgTADRAoh/w9prW9Nk0mnI1VWE9+z893Lbnlg1Rg+lkWB
n5ISpOMKNk3kcImpv5FqGijWwXTUOdOuecOf8tHTG7gU6eX0MpjI+N+lFohcso2Q
NJCBJiFVPbFsFI9akv8IOXFgZyiNHr5SqIHUeJncYfM4n35Oh2U3sTQmuQXOGnJR
+hNd9HIhC8IMa531hcw14+sn8sMqn7FIae9R9DkGG7fDv/AJx20sFEE2ftg5FvBL
fDqoo2kw2xWxQf15AYf+74sju6QfLm1awW3pqqii7i4FgQvBc+qVXP344Pvvi0Zx
uWFbDL3GK1R01SX6MrSZ+Ga0FjLbrlErzzKnEhDknNDz5mVVGof48t1D1bjISu53
FDMJqJ6A+tD5VA9OHccOK36jEx3CZaLgIsMRiOJIzHOjp+1hLc3/lMcHZZV3k1ES
O9FY1NICzfK8ythhIUxtZT3zZXKk1c/kiyLEIryuDw6JU88m4nU/ZSpPhD7R99fe
cOpIXopoiUlVPjwGmArhOg7Qv6Q9+EF3kEvfGNj5kYuw8a777a5HDylTLAOD97hi
WINqa8PQmdfom93PP1msI5lSsyaE46auRAr8KXjRbUZBN9B0OKOdQey+lup7hzqd
s25wZweLgEnXOITR+byaWlzACjzvlJV+UyWalMj7eafwLUiPi2/1kkSTt8+jXoaO
v1gKWIVwJzrc+qP9l7RJlVBZGdrgQTDMAYIFtvnVPKcMpuqoaCF+OGldRg1C+aPl
Cu6HklMW/4Wep6TXN63L8LLCfSkM/9gNVJDaFGIaITu287F77x0L2Epz07RLvnfS
QwyDCqXT8+3hXz4XDIRKUxpXh9dpGZEISLo6M0Jka2HLl12uoMeeV54gmc46IhpS
hudDWoXedrpMZqQbCeXZwE93Z16k4/sntXoBEFGbqL6HhkXep9lViUnK2HO0pOma
4I0aiMgCyclbnVV12eYpKXnWashReSObvH8Y+DMVW+4RKIxWl0W/WvFCFzC9+f5t
JIkG0qwX7zg2bOiBKRc13aibySp18WvyNfLMsiCvyfLw4NWGLEfrG3haqF4sAyrQ
vc1OtwPTC2nEQ/ajnSJCpfoP+lOxZsDfalLvoXMOavfK/t134pWobPa3x69YGEQ5
K7dXBL7bK/WYf3gvxQ2ZJacHsaXrQfRGX0ik0vXlTjzngKXulrV8FIrdVSOd+uDm
ET0FLeMs5y9VomL43OwH1lIKoLbjFMKDK4DoIvoaBDDPKvIOpaSLUK2Z2a7XGzLq
C8io001mK6ovbcUD7d7/NXkVlU8/YpgZBWeNBszMtCqxtnT8sBCRgiq68tmzIy8j
zpFUhDOlK6Pa5WU6qKr6RpkKWHPYfiuKN7LPVajYOIW1pLpcrRtWADDw9VcUd0xx
kMDbw7FX7r9Pnlx/yktBhYta2GiwHhdPx64oNjXJW/dcCin4gRDqexGaL8gKl7xH
zC2GDdy+idTTVKXE68koJIg6+0m05eVUybHA3MIx0d2UMkrlS/wyloaLaiJentWh
TcQWGuFX6sCfUEgYe8DAu8APeGp5/c74uTUJJ2SjueyY7/E3ix+XJzrZQQ2dME+J
LLnp0/si5nNdBvig1M8Aang6gnc/cLN3IIUtnfG5fn/tFWpW9Z2PCgpQk1/dZO/e
0OzXO8YqvT8YTS7sufIStEwF25SBp74tcOUEEv/GWA6XWlg3oQSHvpwr+n2hKRd0
54fUwx2pRRouRHmljNtzUw+yg1PUIgMXYVCNS76pLpjEISv3H/9TYi3Px8tDws01
WZ1HwoQTcZIuUXwbeMa1WmUk4482vPWS/LVk8e8urFktS879Q0J4F8whBrfTF0Te
0Iv7+j0HGOECmv7Lh2lXTl6bHjKghJR/R8u4Bad2XMlA+VG1h72C1gJ0bhHZ1ACH
zUNNMb9rw2+jQl8mm8UeO41FyjRibnxLwIvKSJHVnj28f8c7nUADkWAuIRoRsgTP
2VOQwvBb7nlzTwiifHzsANxcJy+NJ8fHp16qqUD/j2mFYkO9ThFfFMwFD1mqqbeT
AwQCpO9kGVe1yrl+hjJ4prLuJv2GNpJwmRWoyYSCTWz8y4Tp+vmFGxbJdDBibCA7
PMo0u4QS2r9SsuDjt6AwPbAMyH8cIFky9zloJtExZYOScsQO5xShk7mlCNyFhZvJ
at9dHgizSGsWSgubrDjXUtmUd39j7NAS9kp/9If36/oP6xTUM8h7/jNvfv7Vusze
aHUAPYQDcvTvr9aIGYaK/T0QC0TP7FshOSjt6A/SCY++HjLtcpsr49EE65hOz4In
cYyHGmuNi59CCWjt1VHKNnFD1gVwMV1jRxWf27aUklbBwFhW0ftS9DLYu30kMTbh
nVMpzLtOf7ib4CWcSJm+ZeCd2TZ/hl7X4HIrybn25lqGB5zohuz3AmrSqRg8w9z2
ZwfkF1z+bsXiPFgVnjM6yzGlT/ECIQhBA8TOlKACfyO2lIxjdbxLspsEHCbzjFQm
XSe9Vj+8RRDwnh2tFIkL+BgxrIv1iNYUVVJnOTmmjTz2F38E5AhaqlHU63uF4xB6
rrTYdTd/BtYm8u4pegRJvcfDwXZ3KfD5JmT4Ub1Ztt6FNHEaIKQMRDDn4sKXwMsy
lYESsABO1YS2Qk0WA61XX3p79Btp24IhEeo9NR/c4oszU6C5koNhOn29h4C++VRJ
GPOgC6s3+kR1p82jvQKjCJ7ghTXObgwNkIjaVx9yCUcnMcuFqb53lIkW1wRKco6u
QCegwcveGlVZPrgieHDrPulwfmEPo1E6CVg0XEva37ZuKtzYcAnD676g6iWIUPTl
yHjxCd/W1jhfxg9rg6RQvcL2cxPf30gcYTvF/DSkk8gQV3ZvAjMW0rPvBxBc4uSu
qXurHyRN9vkA8eqP2vlvAOeSCgRAMsKwbUeNRh4fzFwtmhqO53cubR42Y8nqDiYH
HegZIEkcv+TrJq3JwMoI00WcEyoEtpVQgtlrnAq7C+ra917ugUYLjvZWDvu7Ygwk
A6GYLGAhOrC0rhq+f/TauoQlxCQnDRsYiUN4990TW+9h+Qn7rB/EB2AdhFBVitzE
4Zb2P+XBESAecYMBhqVwIB+8DG5ZhgjPjjHLZfObEjBJYfFefbZE5XlEDqyKaenC
/d567ikX1yV35/x251KUSxesIz+V1aASgrXRwW2Oi8xh3W1V/HvgJLnAIx/tl5Z7
Kh/4UuaFILHir9bQ00dSgikftSya9Jp4dbR+lSS4/mXbRiJ2RZ6Z2TDCFTXG1iwL
TAwi8qkVBCDFY/+NAJFKWklcMtDB0quuBr84ybIr7HwU+VttcK3Dz9Q3nXk17zPk
dbwdfq95RPSn+5Ze+BUL7IFtv3MVAdkypN6Oo8BVqRitJybbR4jtbpRSTlBM3Dq4
04LmlG1f/bKSmJrxfWQ0n6IYznHDlUtqoRpSmXYCbd93DUu2Ng8cj3c+FuIl1i+/
z6jxAXK3UVRfThpig2VJOPPH/dSXE6gfbfMkN/X0p+uWWc5M0UFjWDBthF9DXAq6
zSrPBKbeBkwgNZpwl31q9n/fj7wfx838Rlr4AFUe/TeZio0ehBUc1ep8V2Al6tc6
DkLAJU3Zvs8uSnoa5HOH6OD+z6dDBL65Wr0E+lPXceMPfYLpw+dL6P24ZYYFdTem
5F/ulLEaiqdxYja5HOw1GDjx1hyNxtNBLpHG5hPFmUhDSSA/wLUmSaGiKs36K8Po
6B9FbBYzF6h1Mg2CWVl8ma+fwIfZipUR4zzIqFUARBaCv6vsx5NDtABzp2eTlT3Q
/1tSH51fqclvMg6tfDtNHNCRR4jVxPnM3CmYrj0V/oVuUBQjQGVPyotHaeltbpYO
zclmyep5ncuF7fzwGA5rD719Y96SgIbZmFSkPZydfFXGarkqq0AiWgN6BbBmBe/T
p7zvdRSl8yraOfu7b9I7mb8aHe8CMX3Bq+JM2yOr0Y5Uxcfq+AtDMVc/Ee7KWuHL
YRGI0vH8g2rj5bnz2gY1XCgV6lMokXhN1vtujm1UO1livQDPxmJ4qvor2hC17lS3
f7t7xxCWF62zXrax+Kif8Q4RfEZsId0IUQ+iVmWU05vRVCuF3hu6q4+qiBcIAWEB
EAkpOxfU6w1z59FBObKvhZ7DU9b+npO9RiasnyHFqpDi9AapIioH4NFIWIOdzy5I
yVtzNTdWyPR9xjiWfoj5e13Ptmw9GbBb6sfWNQphBm6HNCLvdTPNcOmDxYSKATV9
5On4DjOudB2TEV4PhINoeWHPw/SSoEgLgeWM9KHQJlfUPNLJqTwHgQbd9q2CL1Z/
HoGCm63vUZ2OAp6JrLqJuu6kAnEIkbPG57qPSjvmLsuZf+dyfBObDSbOam4HFNlI
xV4rc4DdKgAbqUaP5OAQxRWxAcN4gGVvwqHEX9waPaAvfA8UoG2ect4ltwxiDbdm
VuwDgcgRrlKSrJiuujzVHFWAKM+d5sxAjsDow2krZEhRZ/xyW3L8Cq0quZ1q6i6F
i7Aqdwp167DqqmmATN2Wy9WIRa+ayeKlsUj3hAm11J1nQXCY591bWR40Y/2ntdcC
bQQb+r1AABaqM1nAAXLfKzCRDawmTHPR/X9uUnKjt7IncEAG5xDqpSczMt7kysI2
FeaV0W0hFlwjuLpfcmrjItd9/FRWa00prfmmGEGJnPYA+plwTmgX6ehO7rPwqvXt
phdgxDD+1bECqB0YQXYlwDs4l3XJVwdWeY+6eCmzJAUWct0QOraStb7b5iQo9arC
VFAgO3QINxl5hWFgIxmm3XuRQHv8+jtPdpNzC6aJ/eq486ew7tJ4b8FYci9QK/ug
/nuFnF8dsSQgpfgj4Vxd10MZct3iLDMeTEQyCW/QwAkK2yID8MQR68zu97Db53EV
Xl3Xqkx07/4akXVQgt/SmrTc6Eu4t121bfbUdOHO2OXFN/CM4mD9u+72FQhyctxT
Kbo2S11gGtQLU7qn66G2dy29ocdWxzCH37Di68f7iqmWCxk7z4y9Z501+/KETwtb
8EiWNBCWxg5tGsNXlRPADFKeKvLoX5aIwxWaQnFCXFrj45ZAXQbIcgevciVUPtVm
lZrVCdZ83Mke/jx3v7n+INzs5nBDsHjcYdMDf3DXwC2xSBYuOS3GR/Gliz45Htt6
Q0xIMLmYWmRL5J3Vq4yBJxSDCFSeLbFeoxMW7CIS3oj2bti6OAP7DotVUhYLpXBS
3BzNxbUBnbXErqIqotOxhjHe7upirPm7/7VPEr6RkY1iiW83XyjDOrZUSLzlC+iH
5sWgY2SrA7qAYdz8urbOx0vzHnbdXBhIi9ndJSEH56SwdTNMcirOe+DredOK39xu
Sv7+p2/G35u6MTvwoiPOxfpEFFLdLZfIABs+JWlYjpdR9AanWvIfg2+kxMoJIHvX
0uhmZxoeMgtsO/iXgvIt2tt1JhvFS+vgr98vkRfDo1qTfiVQMzW2bMuFC6ZTilEm
1ROXablQzDgFxRQ455fNi+sb/8nAtcyHsFitfbU+Fb5khOuUA7fyYLEYm0FbXulJ
dujcxluEt8C/tLT9OHUWzWdfB1SnoN2PTKgSxOkWLzCtfFVDXbaaOZPCtEpTgCAP
pgburCabaE/ztA+aSDLnKFAX08OTyPZn5OekPBIKNUFMD81yQSJJwghmndrm9Fic
hF4/dlrB1td+sUH6fRhEVeku19H0KsAu1vnCIbJF5EQoQx8ToQD8xx9T9tXUQKx/
+ZMNzDAm+MVDPv3C7m0edV47ve08v/QsCF3ssgCk+76KYMKvLxPjtWFSe5sOe+Pz
3vKpPfK4KtRuHYxj6RAeiaiwdg3iNzc9AEjGoJwAYGWXg22Ap0qlh91s80eVzFrw
PGjVWmwqjF8w1WGVohlH0pEk9e2sGjNEMafVz2/NQsORslPIk1CzFZhyn3Y5hw24
Gqwu91aK5SxCgDH+O5Sfgx4AYCjZ2jJwO35zz9uWTEzD7FaQB1o8oUjioN1MKI2/
Z02HjO6hpnbhbibpAXNUzzxOZ2qwWD5aXEkcyybgk/gsNKkSx8hCEDDWb649GNJR
uqDY/kIc8Nz7xfEFae2j4GWFLl5PeYlt1VwBpTZm2HNEhjC+/1rO/PBmKimQX5RM
0tab8qRM+Qk2ytoLzqZmG7WVUMaEYVgf1PVp4nmnJiT+q8mBfNY0cKGVh7G0/Go9
BlTz7ARs60lCjo6hB4Ghjtc5HjiUKb6Rxb3nF7LAFZT3halFCSaBYLurNG7pZTc/
sreCKSo0BE5t39hjbLC9/zMEaaVQ9UWULztyuiSSdKf13yxJN2kxettKnqD/zbhB
kfULPJxX/m29BtADXI8RNqcW+YtjiDuWSomL7At6s12HJIw8Y3KqL65hQIu70Gs5
GQFaEb9aCAxdiVAbAMF0eDPhIceU5rjgxbeH69v/8Lisicrs/GfHpHBnqtcYBGmy
HAXJNF+KGBQIqh8uYGghgSE19bdW689CojoH6hK7f3oIcJaTU7CFfA1z6uMtNPb+
nKKi5snO+CNq6qrrbr5IZ/m26rCajvKkyKrGy+PSJxQGrcW5WSPku+k3Ks6tsXc4
K+Kh7UJ2m9TjfIn6weKSafre36C9UgbmGYFJcXPF8gPM+DISr8Bv2WE09aCc/7It
vGQkTCkWeIslHdcTQahDQrmQXz+fknP53ndpupitqRX/EnatvWsEcNEO1reUV9dt
o8xz68vxU3XzdQcfS2JYXFa95ITIolvBiLSDsI5iYzM16mO3++qzMDn66HYipKRL
l8D+lGGzZh4wKxIKdLPvZAp6VkHf/CUqQQwJuPpPeP0lRMdClCIBzKVjciBfKF7R
N9QylPmeQNhVJtgyKFzrRPaPR3Y79RYVhzrqKAgfg/RMolJJ7qm5syUXVIpzhCdi
SWnAkp+ks5juNogY26vGQeMjZwPTVafXM2Sr5g3MRFjSPdjpYROFqc71632NIZUj
ZMdDj4szKvK034uxKOedDfCMQpVVVlwZRCi/ZDhO5qFeVNTYklZqQmVvKhgR8zVg
TfBRGi4G9RHjxeogdfkE2QeUMqf0pvSYyHcs3uhX9RPDj0J1Xn6tRUM5tzGmlDLZ
CSXjsXKIa7CuFcUIX/ldO7+IUPSVkyoxvF+OexpStHmD4bzFoavarRRYDoFlRY+u
3HJrInz5NC33DbvvmfNmCRILZZY3w54jDA4c7j0HwJ2J098ErjtQyb6VvrhkEGlt
wC/5LjrOHtYdcEzHFB8KRgNtMobT22LsCwKZhqLG5Rm3zeL5KXFilx0vXpkO7eqr
4KIIvCTRXZr0rFfz2V3GCBHlSPK2mHZmB4iWhKiphvatjXutJSZMXne7IyxpTKJi
e5+oSa47SY0hKf3Rt5gEuWCUfv4IiFdOeTn32fH9AAow1Flku677In6GxMTWeiEl
IpyzMGY5RQhCiwqaEbQrB8+i42zx9n5euohhnZm+U7zy9I9kJvrit4fHjMlSmfFR
Poon9/ks6DRCc9kbMw48Y6LIuAXqGQc2BH1lq4ZtHAWeVnToZv0gzjK5qVGxdqtY
2C7J7duQdKHRlVR/UpJNCnYcQWfiikhisLZ7SiyvND12AEmLisXv1fMq7eDNgwLG
q1MYb9ZtQpBmC3PzRe9wDc2ROFrIvvFvvXEjQ0Y7fbIH6CR4B3FdO/fONDVdyOtb
0AoB/pQh+TuTt3AxMr1P8mGokQFBqgQWF0dTpaGswt9AmF6ID/3LmLsHsWe++3nP
4Ss++ResdfglmAPZgcKKtW9NusRfxe+Fibq+iVw3DYyCbkxL32q3fbfjMPnW6vT8
V+jzYwJnW1yTSXVqf58f3Wn8aQntDCbplvwdkD8t9nV/u0dAMLycE4cgMUPMIFj6
BEmhYTWW5MzLvvGJW9gBFYK99iJwiCpaXiYELMry4/uj7znrajKM54IMmOkdYI/E
bCLjROhborjNiwguKfqXAC5ShZaOoohZVpdMBMIsyn8WeRJ4Cc5gCHns+Ybp+KpD
EIMQQ4Imz5tBicKZinQqLtlA3yQnzOnB4epslIre8SCG6cnTNf/xpU0JjR9H8VUn
O9in1An6FglI5P2UceK1yuTaUYoyYiobuBokJaC2867zjQ8dAOAQ12iLFv0bAvra
dgCwAK651nvY/ucsZMHoQkl2Et/kHV1QRyWEs7D9ZNhegxRffePmiCqr8Lpl2vKB
H0RGSN6PMAnAWklqIplWrr5XW6AsPJQ8Pg4tPBRVupUGd6kKTnft62EUAl0rC56L
0Xs5l8yU7wagCNGfVxIceNV4/ykrWarLaYe530RBKrXYZhtdWyoXkrTL8M++YtTg
PA4fpBtIvJqfvwzD4XnE+NX6Xk34HVPx8SDB+Pw5hDtCPPFCdqBW1vFzlcbjxPYW
16wWoeQs/XXJEK/nVl7v32LoczYcXB8VI+0RzsNO5f76LufQfOdOkjNs8OcnjBwe
b8yXpjjM+5JqiaVFYhgk51vfGrg1CeqIXg1zpip4xpIM6vJq4ucYzSYjkomAFf11
KQDl2otvv0L1LkqLfNG2rfsBy7uHFItex1qCrvZPlpaZQfPWDIla5XUALvuD56GI
s3wGX3biWULemJ5wGpmc2HgKIcnDzxY01e+zVXGKImkX4gWf9IhXobwcMNdSaqI+
bRWqTazfsjS+FrmsGZmFzKQDxQaFouYpd2dipbEZ+h79+sT8X67DTpl+XBHcje9r
94fdKT/owd4x9URIwF+BwUhd+jUX8to2qQTwxVxzl8Tq/7NTr9YkHBlmcO943IUl
NWetipNfFHH7nS7XiUENkDIs2nxR0uNSCInYF/QALxCGcw/dGQCgOBTsNO0lLjtS
WCS2Ok0cSAHLWAsiWOo3HLrjdMZ24x6+G+mmCvbMxUFo2eUEimViwqF/gSC2xDHh
dXrG8rQG8Dj/xR2hDgsAWvn6k8+QLIrNVPCtOnHh+Nz6yDI9vMZHwQyJHerpbL5J
HkqbJCKjqnvPkKKEqfSGj0U6tZQCcZslcWzplr6nF9nPt/AdD6S5B/VBUNbLkH2+
xKhwfzbkfFmd6xTovejlHm/JL6h1+2hE9d7lWYHdV5ZLEWyHVINGjyXcP6gx+qZD
cEXv0EsHz3/wjcYnZtd0xlD0FQ/Sw4ZLUczLMAqGBqbCExxLqI9Xa1NDVgNEv1lN
b8m2lepVaEurIm0cYrF1e4800Gfnho5XSAgnUthjwXCvpE8mwDF/SLK4m2dl381k
eT3TX7eZDO3w1Jn/DwtqpE4DCKnthUPedH6kRn6UTFWIMOw488euyGhI6IbSecId
3poX2qxVrYebQokoZ+u6KTjoh0fA1aBhYjrouN7INLtbMOcE3LNFxFddG6aHlk1X
nMyRwn6TItxI4FPfkPJQcI2U+LMD53nCtyxCU4e1R729jpBeIdUyEyPHu8sJZGfr
AJ9oP6DdAjMcbHXK8Y8bJV2WpA3vfgqYVia1dWar6BzbjvplmyuaGnikeMu7xO4y
/i/d/SMP0sIA0oC3LSly7Mw2KK0EwoKNrTVyEbi4Omv6pmFsLYJQjujcQUtE4Ole
RpAtB1WPhWzL8qX5J7idVV7PYklhJJx7xaghAUn4TVeqnfUc2W7f8+kJZqTnhYaR
YEWrFFCI8zks1D5sTC4Iwbd965HM08lJVa8buO2edn6ZKx8M9B7+rjwLl9JlMRw7
SxIzqRvK3AZFohKtDRNLqQuXIphRmm/8wkdOU9jwshZi+9Yxuo51aJJyiVhnS2fX
xpJWkOCr7qRPjn4DUcv6GYn+6KrZyfYLdeAin7DRNveoU/Hnptd2DWtmP7keIx5Y
F7KD6RPYuq2eYabTW/XUCogN46IOWm4b56oIc6TUwCw27Z1JVUIGlCkvDAJzzxDy
zktFRNQqter6aB6xRtDfgornUYz1Phir+HhxsaMhtzooBvW17YNoEvyy8HtEJduN
rhJdhPaTmIxX641VTCH8Vw1wbAK0Sj3L6HqvUiEltZKYve9IIwdGA/WTtIJ1sH1Y
bwR80TihBkiOLtjGxXuhQfI4Py40YRGtuGrgAmkEQKkb9OkDEUyTJryEp+vvu4Of
4H8VhCjeFOwsduIKblmrQJIdo1nHFwnjQtvYar7DLqGI3eLW7/aiZxjvneZA0TYu
xXRsO4Vz6q7D+ltF65IG1fpdyzKm2rJKDT1ITAMkB2n7N/NsG4F3kINiRPgws7+t
UWSt1T9jN4jT4dApL/ya6g/i1W+280T1jwPaOmcl4prz7vjQzWKdEkCQ1JcXM8jA
D3T6bTrbxKcF/w6JaM82yBwnLBM8Qjqc/krD5n1omilpXLvsVC4lxH1u9tBfukRC
dt+tq0/jlzeDbJTiZMjOmENT5FAiMdUCxYjdOoa+Lw8v66z5n7mmgVpKxslaqOcx
E6mUkayfuC7RVFHcosNOJi+wMsIm8ups6g+vEOmfP1Tee0ePI9OjJKQRV5LFkQSm
ni5V68BWh99FmxGsCgr9mbm4uDqz8Zm5JRfO8yCt5aqj7BDkx81FzxXKIuKR4D0L
P2be7G8/XTQJ5SX3m+WRWtI75c2RMTnKKOTAE7ETYaE=
`pragma protect end_protected
