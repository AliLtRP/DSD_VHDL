// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:43 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lqIdXmHgokYMqRh/LyqvfwCc4VjwfBl8O0BPVOa4SmsdEtMGTHiDju9/0zxLyhPH
RPceYGPlRLDHvOOLchAMZPVNxqerLM8v4HzvYggZ7xus6++sCp+PaK3YPx2aJrD5
9HMdevM2yebT5qN0S3LHENyuW0zgRWH4Yd7lMAC/qqM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5744)
JAZUvvlAZuy1djyyQUH4wrvXq1X8/8JoaOiW772evYqauHSiw5CJJgTp4kFYnSVp
zBKfpQ00XGfhrTtqNwURuDSQTIy2i9LU1sJ0EI2JrCFHSjvkS3E9TDJeJY/L9gnd
ExbehZPW5nhMR/Y6v+mha1OwJO7SZxyqexhrvll74MREDK24XEYVqakKJCRnF0X2
sPNvlgvYA+v3ApO1AerhRrl4Y3dVhgzdTikde7k7n0AP4qWG/Bz7cmm96gSlRMQP
RavTMAiC0XXivfo/HO8t7+fCQnC6SYVhqgKGWDczVAQBRn4fNCl129UDVEcEBcYO
TCSqcTDd0ptwyrH/YWmmzWlDfBlGPJMCVSbKzZFjx1Mz0h3ShPwLNVGkdG377Pio
0D+GGEhJoaMRF27OHJNWIQb2jvdYZWlZeCj1otnV3m4B32nEtnwFpjk9S4AuPoT7
hCWdMFgd+UHj7nwFpvBcZJG1KuwG7HrC3IKUyQ7cg0cATMd9496tRZ9DgOC5slaN
crIvoE5j+lu0WbmQFNAL8+HR2RvRQJpBsjxOZm9vav4fODEeGsXjhgFimhSKgFal
HjDTJ8nx8Rnla+CFflY/exT1DdJVQGKumWJbcOcLTZU0dHS1+J4WHSY9lsoRNvcO
tmU7wAmRqeTpO/djcfzfbQPh2V/z56GhB9exZc/o8ipY8+0+YDKcHR/sJ86FRmuQ
4Fwh0+LC4kOI17YsMo8OIlWj6xJmcLTIweRI7xsEVvtJpgD+YHhV5+QYJ9FgSjEV
e1oZ2K1aJN2fXj5DQpnEHEHbF/HpQe4ZaxwbqfO5M8Glea+wpsHcYEQqiSCDduP5
Yu/O8tYzjHW+QkrXPhQmWzzCT5Md8Tx7vyzbT2lzuQ4gBY21FcinpO7PNxzaoveF
c5UNGiKNVgVwB49oVxpSlD9zJEXcueemuNtmwk9FbScPj6sSBUHHdBueEZSVLGWV
/6fBSOF9SySpo/PtZHauKmOo5W9dtNJYlLIMk5pcMBbG10l8gnEmEi+Nfuil/kxk
1I71fZkX06VCmRgJ9LjS0KYwHk4/+zw75r7WT7XleqylGekuml1CQ7khbJeCpLqY
+5tEoRvik9QE49AVIK7DnfJNwceQjexQfKZH+Azq1kBNayyS4uLUyMzO578ca2zp
Zt083rbHdJb9w+Qz2/AQggD0fAcktVc2wyOQmSuaj8zV0ppWd8lnAMff8fTj1t73
vDyEh5TfUXwaKYMw54INyC8pKUnlWi669jdSlu0NU11VE5RvFuxq5HVbK5ntRrKI
GE+dSUiJ+3ct4cbTjF2xJdEUPwqnAc8J3Fw79CXEXaKt8osMzix7W/MHzQ5eJy7d
RkFCoGTqF7v63stBTsFjdNE7wRqUMCtiL1Ybcbja2YZkhWRtvYXEFZE99tXQdFx5
Rf/sW8sx+2wIuoxZx9MCvjFQOAZNhOr7mggzpXXOh+BPwWprH8NyKeI65K2ESVyG
G5aM2Qsx/Y9jT/lxMNrEkK2hFf1ZsnKklNHezPi6wb0xBikomvNcBzFYsx3B5/Hf
roQwG54S6Ab10ayqoX5LaLNVs9JIN/t90FbiBuOd1Mdl3lOiCNaLA3uhn5kYytKd
L6EI9YMQEv6bpQ4TfsON2rwKmQZyAwSW9gQOotM+FCwarg089Kfm9SQznxnArXlm
9b1thFAPzSens3/otvdiRgiEKfQ1sFkxFB2S4hzJ/6dyaMkVMjyf4uXQCaTqdSSD
8EC2B+e/0eSiX2+Bdr0PrVKf4kfcwrIqekK8f04wo44hRGo79q82IWSL5I5Nc2JU
nTFtsGWyUsKQAfQ5THGjJDPHUHI1JlnC3VAfp9kUNsL3u7wZFCzA9nW5zE9sr6MN
F0QmoKU+Hy73DwffN2JQop47Xj9bqAo+HICYPMZrBZgDfQtK0n8mGuvzgtU14Pza
jrcjPElazL0sZL9koVmbeNgJUzh3JhK4KYdHCnCBqNoKWL0+vnEb/MOGwbmdp8LN
CQpTTbpvIloDVK/Y4dK307aVKa5Cz+ae9VNG/O6S7mYLykZLAHwdCT9zSaeJdT/3
0uNrXWJtBCoxObIheuKetIKEtCJ3f8PkhHmRkqgFYJMlglvjFwUAkOctHedlDvVv
vRgh3/2p0aSOxDJIXRhsKbciKdTjd8OVnLnuNmxATEHGOL9UmcTRjH/ADe9gHPZs
StC8xceIQD+2HWsInMsFmwEWtBkC0f5SmcX1sLW5B+hNF78KtKLLIKob2UrzL63b
k96Gz4iJ6kJJl8DecCTZz237tuqiT8h4c1Nm64LWTJhvmeG5TwQr4OvJqfNvkt4S
AScApnJlK5tsBfWHDb4Gok6PBu6jRF9aT9y5/z+IqQlo1lWFd+C1yPFR+rlmcUc2
I3oEt65J5GUBZO339aOmVqUqJtHLulYfR3gJY7hTv4A9W2Ovwg68Ud3V3ynM4SxP
T5rfT2JM73giXT9MFSK5t6hDwHg+KsDt9Y/GA1RSYYfs3frcJroOKSvbos5MpodQ
kbVNBtb9tQMRIKz/PzT9VuZUNkvorD0CNzezN1XWU+2at6xqjw9FKgy1iT7oVNHx
7sDI++NHuNxHbfs8TmdjOe1gklBh7w71umZjrPgd+ZQBIN3e6RZe2sGlpeEYlQYM
ctpFei9fIs7VvokLBEeXZjL+9QlWhN8nI1GUgj9izUizAuIZHPYqbWeD5bNI4xyS
MO8/FGhS3kxtm67Ifhm5KVBPmIo9a54SEBfW0WfVy6a4mGvYkEegmpFHb6UCyKH8
xsShY5lyO/4wg+tN7b5Hk2t9W84Gvvd/KXyYTYmXdd66eNZU7ynZSwQ+CBYMCXeY
Mo/uNXzF5KRLmysd4TSSeg7NFDAOHXl27liYs263LPgkMWHmXoBUEGmLQ/VGXrfm
VElYm+wdTbeTIbh9v0kc0qaDP2bWNQmkB7yCWxYHnWOX4kQ+LfPgD0hnVDjdg9fV
Tt6PNbHng4jhVZSPFHCeibMHpR0h9hkaQA9thQSGBftubAvTWbhTey+BGaWMh62f
5ZImldirBwi9HbyuR1hoQDIcLlWF39c+vz7Jg1Ie7GYvTLCUlVDCpQG+RqzrJPKk
LqcVo76826LEKXTz+vSpf+pHaoJgKUt5i5Lr+I0NwrBwbzNERwVKOH93d6V94CWg
Qt6lbT+tDKjxxMBMnDyKQgkDOjjsJaZB7FdxXmpk+OjSrTUY+ZybLPx7Y9XBFEFg
Y2rdB1fU0+q+29pDvP1j4IljZrOChhhieTVE6LtnMauAWID8AdunrU855XOdF8v+
3fvvD2GPP3e2NQ+QmObaBTQNE8tOmODzvBkU9MtbsuAOJrq5e4+d82PfPun4ooaE
IVy22KcmttSziRMoEX4TGVjPmDKlpf7W9o4aq4m3IUOtuKXLtUx7wTyvFca/daWy
1pB2gWSx+KfAdGBwYufkRR/WT4lpoeNsJoRR2Ztt8fUpnQWS1846eO2XNnr01Abm
7MMUX8z7KxuJn68wlupSFp9OzOtn2ixdVAkc2PZ8o8kLkpemGO2CTCYfu2RGfHFg
GOXLe6HZvcpVKorO6YWGnclbf7YMSB6mL4OdNGnVi7tqD8MAAhBnUDgm4HwMGB7m
Iw+1LTKi3ludzWEDMQGtMEqFgqnHFyiKd1RgueJzRZCrfrDint1fNzz4+EA1kyVB
c19li6lqawATQittHC0RtEtPYaZ96/MnOKknHYzDMkNMnP4Ug5qqoxtDlq7+2TEV
bAalnh1DL5b2c6UjF11NtZZvsQWkNTHITCx0UC0CGhI21dNC8US3KjrJm94aU0rv
KIZq4vW3HqtaU0EaDz97WnuVOm5KEcK32IxHCe8ARZVdAs8Cs38IvnoYMjvP/xY5
4luzqFGTLpwXmMj+iPDNvIrEquaZjjZNzkk5yhIQ+CSmosVa3zBYlLSA/A+HIW82
Q6lOQS3+nG4jvAZLsy9b9PdFnTVlodoAmbsFjWnUpnkBGYOhcLSuq4oiIj7pEOAa
xUowgzS0rOHn0FzdxvelviJ18atHZvvgUSPgQg/uM5TP1KrhLjo+v6SLCs1z0kR0
RqbC0P18qKyJNYDWugvQ4gXZwS+NN+8GhtdyswkGeuEZ0O1Nv4Qp5eYioqWa7eoh
BpY+kE6G3Qgrx5XIrC+zmnAIiobBQLzCT7FgD8eOo7ceDp70lPX+qhK6+rcWTzhm
UxIhIvDP5+nxLsX2FVbonlUdzeGTYUqvrNmk4a7/uuSW/voz9G7aYbCNARx4zkAJ
rr+fy8lSazpEggMiZvZ4fJuor6TvAYQJMz8h7u8zk6Aeueu0/4KgHu/uJQpxshQ9
viMX8+VnrZQHZMuC4kDxxGUQ0+CbzJYyp1D9/6L49E0Wh5vje5g1U4iOtjCR6OiS
XRejbhcNr/Z35n6noKOvIG/QU+/fYLFQ1HvHBh+Q0zfoE5uXp8uA3lp6UaWWYBRO
egB7Jmi247IkzmFjBLpmTfyiCJ9/LVS8gN88T6601k8LpLXuhlx3Db89dohFfcWm
CztmBIfDejafpIioq1aKVj1Pqu7cIAyaehPw9OQUGcm/vJvh1u8njeZTcc8ZVVO/
okHzXkSkgmMVDz8PGxx0hY0zDpN28UwemMy27EVmy3est8oZHLdsip/XBvAmWMfv
OJSHeZflHmNmtwgbXNOorowxBXBcBD7XmX104ZOPWySH/vQwgTFCpxvRetmxPEdx
4enxOHvy99LbCLZ0XPiTx6+abvciiO1aV9X4vSZqe0cIUtgXVFY/9ZCp31qJ2R4W
Xwo694loRVQwCN/OBUoUZ24pTHG9hlwVDV1BpIlkF3XWMg+pqltZgQhVEHUcT3dY
o/UAi/RpfpjGayAGf/DnIMCEX0SHcJ7KrPVujWv8XnJO+MODbvnqhTi/auX+cAkZ
F7yL8hs4FI4VWD/FM4x3uvzS9nTUFGFhg66EYqgHhmoFHUbhEkt+TTIQzku5wJ7d
Olc9X1R6nKbhbG2vW2/au0WdE5OR7U8OJfGEsGuu3vnR027ueVlaZm4ihxHxrpwG
rhrNI7000iAuXqRKnsOHLJojkahCpGYjiaZAEYU9nodmg9voEGoi0CdldH6JjGAj
MxKm72eujFPoM/3HhzYsM/8zkNtFxoqRMZ68Zlba0nb6rAN0ROS3oqhJf2TiYbag
bmZpd7cCB1IJK+lPKX4sDCJh5CybzHWBjRLNQ4Ck0oHcd6akYF2/H5qUd3Ulg7Iu
aZoM7ViC45AspQkZxBbGARWyWY5Zc7HyFbSMU4tCW8Y7RYKb4q2xLqbIuqoynps9
ES5AAwOM95LtY++aE5P28ZY59pKB6MlxsA9AOHYbH/nmN4AXxacltM53IK+d03vG
WtHkfW16yWX8LxEyuh+Ev+uellhltNFvWaEi2d3FRKarXxuwAHSmLcFMDpKbTii0
TRnNXIZHOdO82wJa8eR9v67RBXnEbtNxWyD3NFjZiRbq9F30ZhUhlgPXk2O4qrbu
tVGPkHplI135hDRmH8y4eAAK62W2VGIVxs4h7XmTKxigeHm1ZE6vXVhZU+DQwT9G
lrl4WqofcYeBtYM3MqwFoXf3jWvIAx5WxT00/FeGupMcSqbVZsyYvFNXbbYRKNaE
v9CBKdsW+3daqMU0J3903qHq7D9k7gJD1g6QKwYHAu7Moh3ZX9tAj9/K+wobVmyM
9HJ2n427D7oysZx24oOgE1K4+GIj0J46ad9AYeeD2enWhv2lJjtoHnEBYzb/Me2n
/hzY3oArQXY1R/YYv2RG99SJ3riBUsXBNTCpQVhtpKBUvAhm/D7/KwviB7VgaYo6
N3UA6lEUu2C8gmdA5Z07zCsV9fe+NkKrKzErX6b0T5IIJDpUVwjtjHJ6trjCPyQ5
NKlh+GaQJNS2J6B0dbLiIRHmwtrKxDNcN9k8KbMOucoY0ufuv5dGtrUD1WGz+Q0g
wFrHJX51+3ijuggKjIxn5I9hvRF09FnU3zNE/7TupkWFpYHSIqQFYqSuDk1kJHnp
NeBQtAVHd+QL/P+4GuPCy5gdctSQXkO/lBThNBsw3h18s9QLc6Eb4Qic6MZOuN+H
nRSxdeRxGODu3KRdU2f4L0DDwzIlm0yGkgj/XCHcywBs1ADmcqOYhwB5RxsGmX+4
OpF9M1d+Mvd8S1a/d27A5rtv3eHerXSLU5Wx3DKn+5f7wOUTQZ/UNDQdILuGZPXv
osQRCxe1hjzCNQu9MsHFC2tpJPbHt6CnwOCtTvFHCZVgDDlaRGaiu3Aq6A89L2iI
FjILaTkt4NX0WddckxwqKXy4E3a/iVrodMR6TdSZ/rDZ2ndhbhWf9S0nkBT2r7Rm
AbHpR7gy8+9wpPERQ79cxY8y0+7GA9+yghGmU3kwKRCivemK9s7zZs2bv76speRH
lHU7LBKxM8j4N9a5GxWwTLboY0gYCmb6BVX2f2AQdtDGF+AnsCVkQaSXZxry8wkI
KTMbC0QDxZBpKJ1q8e7WsjZGIUilI8cRDd3EkvTPlHsif2+Eo1+9ztTq+Hmxumtw
di3EBuQ5x6FlI1+LAaqfmOS+xjlaiVYuZpjcOG1Cj0DY7Y+gBZ9Wgy8M27xU6HPX
iWKyvo2ESEn+x6MkgL6KVMXYcQ61qhrKjvzxTJzxAJtpMH26HKaH0T2gS7+X9CeI
Ut0dKqzQopQ7FDNNOqU7UbdX4BewqfRRWuZZq5wV9eo8uSJI7SQAF2h2p8cLJIXt
DZSLIkJozv9h63vwwG4M0M6cXEKXVeP9Ne8eQ7d1p8u/+QdRPaSH1QiGQXmnMHsG
aWVylaVolGbJyrwtI43XsWm5Ia9D5zNdqfaiMQRMZ5f/XdwNH75ribvhrz+r7UQk
q/jEZf4ll244MMMhXyFoejtyHK0d47CNS2BX2zKKeAADzbqr3UuEJhx0OVc7CLR9
jBq8iXd6U0XtZ/bPiz1LNRvNYnvg5RUxb3035Ao2enmlgkWSXtQhE7QA+vpoN4hw
FRoay1r5qkB9S5JB2xuz3kBg7B45Idy+jDO9/IQNzMbtcRtU6PP0FHgJq2up/CE2
pBR0fzAN1QGspcxdjmUASPZeSGj2Nr9U6sGjDi6a46irUyWFC+LDAzrA68P5nXva
2cDu6aLia3LRZK4IOKvn7myibljCZCEAq8kOjqkgLi0xbH3ycmrkphv35DVSYK60
3irbptiokFoVBHYVu6jktDDdy8Qx5ytnQa+mvPCD556zjWfK1/0ApJ0PlwdzvIXJ
shVPApaXYD138k9ZFq8KXvxdH4p8ashHiCRxX1SDy9Pb9lXMpmrqU3WWgdsC21sr
/v3kNarGrI33EoyUGXqcupCF0PwEGdb2Ko1hM1drCSJFxPIdk6g7UXd4bmxcUuxu
AfSfZA7+2a36kM4dD1W0uZ2sbsm1rxH8I9wSBGm2+nHpb38PxRb9wBzC4UHVebhI
vWzJrfmXLu8C/Vs5g0orhZqnjzBGXdoTe2zPXzNRsViRpNL4hs49x3nIwBL2p3i+
C2fOgmSIcGGzdq7SDTuOFbhG8IjZSpSMhthOAhaxO0VBwsEf7CEqxtcxcoxB1T/U
RUXmpXqbOVX7K4oj/s7HeqmpY5Xg+SHOqWfyPlXEq7dyWVX7skoU/+tXY1bFUwP6
wi4u3uCt9ZH+Hlcgk7xv21PJGBkNFJvJXIObCTpV2GYVa47DS1HzhuKX+j5lqMr/
+Ilb4YdZMhJn5cmhCuE5tuLMZByr0jsbtZKx3eoqEJg=
`pragma protect end_protected
