// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:32:49 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NDJTmASHbr6W3J4PyJKVXIt9KGWZ7YWJrFG07hhBB4OquULkAObGNnZvq5ytc7Ss
L1L5ZkaJueMETQI0P/duOagdT7/P3C7AdtXIO0V6pBFoVBkmqh1sIhYAD4dFsyDK
KgYcoP4B1xbtC9xItn0f398aD//O071YhxRDa1jBiAw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4048)
lR6yeV1kPpdVFeGCSlEj47KhCk1qMm6g06j7r2rNTT0FZj1NAuKXV5aSPRC/cY2i
EC6JK9+x/yQdUBLdU25pBYsDJuxsUgF5+iKsVvZKF9ExlIUXcyfWjD3ekbXAvWs5
gfpw3cascESo2ETzz944d5pSUrTDvsog7ayEnf81Jpg4JRobi/cPED2hPDBoy935
kuQzkCG6ImtiM4J1I+ydmqOau/sSV/tKJXwZR+yMLWfOm7z8cBp4EFDaXMH2UnXp
XaunQ79Yax9a1i7HxGUWiR7CqzEyIkrJ3mqLtdJ/0oCvTjnoF97pi8e4lyKFinEA
kFlyvOB3Ywvp0bdFon/fqqwbLtQEjwUp05ResRoxVp3s0jezbGlYSoLQFx+j9glt
qtCCnfoVXzeQdIoJehAcB7eOzs9RHvvZB0EwKVDOliTdx9a+C/Kf4+e8RcLvqzzv
A4zZVCNM+KybEsG5DXf2JACZSFB3ZVDxIN+z97/UEgaEAaGlD87JsYcQt1qK+Q/v
se1Bwp5f3FsjrCHZlj10WljJb0LR/AsRbp9iv8tQ+KAuAdtg7qBH8XO4pHAO+yTe
hePa7TPByIcYDCzobB3sRJ6GAo9rqBm9fQosqJWGpomSwaYIbSTgAMi3m5pPx70Z
pIjqkjuqd924gf6BmNHZZkKZTws2OAELnJL+UeRZNBPIZuFVw2xQTWFDHudOgayF
j0cOQoYBu0cvzADz2/Ufu6XWqGuwXfz9lenzZYrjyLRn6fkfUeno5vWwzDD4Bh79
mgvVwGHa93vBverHBvgwbpdvY9C3spbsBub7JrfMxdcA3oREwzmLZ7HGVZgsFbja
Dv5dJiDcbsMJz1tHk6725ZTTZXIwBCbCicrUt2h5Cz0TT8jsD/arqgu2bf9d4HVr
Pgk11HI23Pcmrsda8aXiv/heB+Rd6cWy6I4fn1U31K5FCPG9Jd8fLXIRqD1sBKQM
horrKgQXJ/yctSwv6wnUMWLCZ8lMVGIEEJgNqJpgNGqKl4Wp641DIRO/yp2qwYtG
J3RFtPwU7axQu19za2T0QooYB8RdvWxT0sHZAOhcU7ad6NRwK8/TVikxDbc08Jhx
TqtnqQIDNNDX+lZWewR3ZUF78kESkHALEvoVN3xnEEHs62WvlQdSjjFdeqeGDhdu
IbUqhK51lRVtetMCVCVNJt4wsGc3sYZGgTbcvCCzlW7mmFMQIZuL1+o9uN1Sqs/K
VL2i5PCkLLd0YOi3ipjhGMxkXkKGmEkfW0/CNwjb7WQWXKzyCYIFK0NYA7GKJRIR
YJFSOjiqwybYdn2AKavGheMJMYDzrYP9mWEInsPR2nsRuIXfRB3ROd2KuKALRSpn
NwvoOvywyBtEuczueicCMpO/iE7zy5pS4Ae36oUHUbXlZIWckkpof8x107MoMgMY
uDG32+dLVcMcME6zZg/Mi32um70/GD3Kv4q3QYslkL/S4gIj7xzfXv78eo+Eech3
m1Ca5bBoI4hDFl0UzUqjNhjxh4RPHj9RyxrCPH/PfqQl5vSQU11w7SK5LY/wErM+
McOHw6GgGT+IvDBJzUffP6w0ctht0Z1NgwfXpfgsF8we7ugCdHrTIWvnP0DFlcBm
splfEszz2L5IdbAW0OMIxJDWQPgmhVnWDjuQ3JRKv7CEfbv+xBVNfBHPQQ+b+r5A
HqQT9OKdgCLTd8WrndwGRnqSgjX+4Bb1rWs7OLyqlh8BJ+j8b0MjBRXkZVI04YtK
PzXo9YQDdzc3GxU2mA3e9D2zCf/eu036GEirX04cJh7mPFAhKqO1b3j3+keKIX7o
9i+YvcBsH15drY+mUMT8X7qw1DGdJeUlG1Vq8emZ7j3pV/Y2nuzMG/Ehsx5/tqBP
w01+Z1JGfHJigcOwCcgVegkAdQRLfpWYVvqNIEhR2uaS/AUjIdqcWtZPOxswSBMz
iAurM8+fg/s06peG8v5UQC7BLLl/shPQCxZAe1i1rRdmLy2SzII0Z4FBxJwL3avP
FTmf4JRhHyMRJXNcfVQIoLDZtqbieVOaiZsUIoojDI9nRO5x8GU6aPUFNSWh1yDb
jaabf9UGRAb7I/f5+csT5NZOKnsA/wmU88634zDIE91SqjmFPZe7I7vli1AwTkD5
R5nlUjRLR+/fnoaiUSMR/9a+04RT4VmI3JbvydoFAUgJr67JxeC1ynCyLSsN9tqR
FhexG6nts0CMm3pgWP7wnFmsZgxLi20Pu6D8bkJzgkK8VkqzXx1MKZ2oCWBeEEV7
fhoXYz0ZBw8DqLn/woRUNcKom2zQiVyfeuEEzMHHh/yYXysq+kWHQRAykl8JtrcS
cl0Gjt5Mh8FsajJqU2C94rDg6oVZW569F98bqi+Hg+YeUqSeM1X5HWob/m8nbwOG
m5PPIExUbleB4RcKIf75SFjtGyk2EbDyR/VvG7RA+ci3LjomHZPhKvSDCVJNT8Ic
OmPMdtO+fUfJpWfZgtmMiyU0bp4UpvKTyqeKaqaThsvf3qL/ItPVRGab7HiWCXPW
MFyO5kCY9PkKJBRsngSn7c61inD2Rg5aqvNCBchbOsQ5N2OVvebE02pxKdolB+xh
j+uWlQU5Cx7i1rvIxV1MPmstaFJOTvWguR+ZPSgySM6GzQTiNCG8idTP+71X+Et4
Wx3r6IGMxL8i1VOmqRAxinIlN7ljUSNS1v8oRkVnup+tpTpWipMxOY8l2pEHK8tb
3I5NoOzL6ZmqL3ig/5l1tGt0QaZNu0kCtnwFqoNO3BwgfS4TxDzyWVPOZ/jqtYCL
ToCGD4R9j5syuIH8gttpbzqNC9Jfh5i6/PTWutP9zoio4iIYu6xglWAbbZl2YYfU
b17TmhKIIg5TGrk6O90hkwYTqOjR+aUbQiVl4sX+nzYpfsdAZk8zKMgv6iGajeBV
Rop0/8GhRFVwbc/aaYLb90ui5lDWpxMXmDTJ3ros7/xPkc6tGwdnbvCDmUkg9Yap
G7+eTl5KD4RaQeZo7DbXncUZwyB/I04uPojWHRZpQUI4D0EXn3UFblKGIZ+QPx0c
kpN8gXgZqyfOg/5YOZkuw6FOmKj1yrD4Ipf73eF6vvnh4Ia0uP4+kuzIrOnkloIs
F4Ym80dwqOV2P9u372RWvzMyHsv3AEWDDp00jTNxYlej6IqFOrU6bfA5sZHfOGWx
DnWNQ4Ms1venWncudy9jI8nT7XYgxCIqy7KNbOipjjGmuqFXwz7WXlfnwVmqIdLW
ZyqGT3APwfA6J6AhchuUP24sieuhTGSr2TJkd4C05v9ZJ7LuZtST6ZFKwKxFADe4
GSB4G3VA71wN9pcD4AHLHOvc8ws7cRXrqGwkCtFmdx1uYCaD3athKXMCfKkUMK6O
5pdjBTyyJyY3/V/qFAHeNx/BsRp6B1crYW1mwjfrG7aiWwp9sa/hJ0FSr665qLgw
5nm6gXyEQAxw1jXybLn3tBjddivXbWoAOsvLflxw68uHb65n6vwUpCIH1aa3EGKS
62owdYFXSQLhLySy5mFXaEuK2FtUcEY2YwpUtZOkqdKEumG4fMUqUb22ooeCdTPK
fYjXr5y0bQynB+n4mp+6Uhihz/N3LGSCZYZrj8Pa81GS0p8zafkG1i6ccX+HZaon
yyIYLI14u+L0H+/a8HvgMbmCp8jmkAOVfXqWTQEMq/f/dEdAx5sDvCUJvGJaeVEA
rKwOWFbo7ViMoemXsSva0mUBpI544FnSaquy2U2KH2k7nE18YkP8OH0TatNLzn0n
dLsBJM+bQLXQn3PpAwo0T9ex6DgKrq98m8ECfJhfaK3LTgIIIEuZ40mu70nzSdz3
JhQme3uIKlH0cDQu0e9PNdG7V2ZauZ/TMceJ0l3n8U/sFjRqH9s6iTvXuLNAB/Kq
LeeWKkMlTD3IhaNF2jrhlWQHMzhgPOXmmD1O4ApVV4BvWGYvc8kv4+9ZAQKezy8X
F8GjTFp+Hl5Be7qvzZ2QE7nD6tZQQGX9RnmhG9/RmhfBfvCxYoEMdJgSBdTAoqvL
lzREm0YFRkMOiUSCPReANpw2Vk7FbCWvBQgmggY7SxcYQ1Oro07YdR7U3czrogf0
TXLQMZcjQPa7QF6aDNovvrhZSv1b+isVV6WRJ0ighQjakqQrzB4Bqh2bevCsQMZs
O2SygrzaCyA9IZTk78eXNaD6Q7kPsgMTFW/hobyTPMUrLXJJy+WohR8JFSm2dN+d
yXmroP3r4cZkchARKMeMs2yMwGBBo9VEksQeuj95oauvovDfUvz3a1eAsiQvRFrp
kbxM97MwJpwzQgTLEU7hzjdbI6EezUp7NieaC+IqdWMEmf15MbzY+1SHCnSizNz/
yvpD1wW3FrmyHoDMPLEVvDYd0Dc774Bh0Z6dljjSG5nFHzK8P/BTapfwGBuqfVWU
/7QLeEPKpjjLIJPGzq6gLmZV7vZU2z+wPXQj8zzM0sRyH8ZAUMSyBqaIOAyLatc/
HSA6fLE0HHzqFg8e1ZCCCHsJWjIGOCWlTCPzM62KXAjd2ESRQZvd9VlyJ2+5XXBK
yl4PtzDOmgG+gxtX6bRMll7NatOCdO0g/s6nAlyBwN4vr3E/I/yxt44dCaMtAVNP
wgEuRdL4SwTlrrWV12Oe3hDdHCrpM2HAzJk5BARVWgyej0ZLuur+NWaZfAMs2leh
5+fzj+L5+NOgxfQvG4/STxwL6UDNgyr6TQy2en6kiMlWySQpKre3xLNTA06SNdr1
HofGy47kZ3m0IAIr6Mn+BFG80Y3DRQuWNUKg0znlCl/+TWy/g9peCGS68blxjEQw
6xRqTg2lKD18aIHuvniIsmug7FRK2gU1lO9Igeff7Ny7b+vXh28zFnb/a/ju6ssN
9+DzO2Kdk0XTslgP4g34j8rv7xRFENt5LAF/RbcCPCsbv1RGLj3ZslgSNWlR8CEf
iCYmpOSdrF0QBfmTuoqgiNQkvtSTMoFuvVx74+Bd//XiDBdjdQCRS6NBy4PD/4mF
V5b4qAR/AIda2MfDKykztFq00P0dohpJ88v667stQGmUGvmfTOwPjnEfrRgMk0q1
JNkkzrhV+lN+htkGR1euzIejKSFw+hIoY6EfSN6QEE+kpPNKnFFhv7y8Jrh3tojF
dC5HZfsdw6KYcBUSchXHwE8wck6rtQy9W5uYZUxVGKVDjF9SukFfwXSIH3lr+XtK
iBDMuWXgBs6Hda2JZtEo/rijzPFa1iJL2TFvJFyerUYVI/JwCgJ5RhkypTiN/mWy
lLNtq2IZvikhcKdUXM+rf8+IpmbWaQgosBRQAnzL+2MG7awEStd9J/sG6I9oJ5iN
UgEP4TmFgLg/QB0xxANegsJgQMncm+DowLR3dzz9AiBFTDN9NUrUvtt0uLaf+2jv
TWw97RX1Gdweqf3xEX1kBat59vPb0iSLETUsBKBs2XsdZ/2IwaC8VQzKZyeHG9o6
hcbLezVUnex01Tmb0E9W7Q==
`pragma protect end_protected
