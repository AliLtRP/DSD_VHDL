// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:35:45 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nTqQ3EAcuOPmblVDKzw42MhdAhXg0ekRt1J6SmetKk4MYR8rpxYeqzk/ysFWKBYX
Ve5tD3UEnZmaEDGC2NAt9b/2edGwLmqOcJ9kKZZdCw+c6cGXZR9/nzbKOwsyiNt+
WVMWRTcsmilekL8hDum7mGLqcNzEuOBsF942ZTxRO/Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6736)
ZBllmBb0DJjmooAgyM80QgPxCopVUEjxDCb6rTDELchzzHKw/hH7/UJsf+8Uhd4h
G9glh2wM5znVmmjJnrrpZj6wkWsj7e5fgeeaeOd1qPj99pBDEzFoJrq/N2ui9X2v
6iDxRm4FPpbcuojfeg+Am2/K+jGNZQywIQ5Y+2Sw+Qbm4/cE9jdpeteMoVXUzg+g
spTXHNmFnj1gvuP5c1WQ2OYcUhV/KQW8z/4Z8ykw5MDstQWJSd0X0VH2bXVEJmni
rio+bU+tQBBVN5qjzLMxn5LrMNsN/UWOrJ/B3RKwOPehY8OUgogMA4vWReQI5TuJ
eUoZoBTDAYRJY0Fd+OfhCz68OTysfVTBh+pKFdus3EkZe6RkbgBctgvSWuRILd7I
30RIpSLHBsfzMYTx9E4Iaf0946WCRm9bDAy9oYAOEfIBje5yA07uq0bZuLQIOT9R
5+iV/Jm9rO5KzXvLKvq+ExaQW6o2FsMRRdvqvUnqFEc48IEAkvAOu5DHrmWXwOov
NZ+vX7Yf4lMriTpvXUevIqPWBApoaFEJX9mJHj7fXpejPjB65wCOt8Tag9pt7Ypg
w1uuXokhnloEHFw/T3LuDQZn67R0ArxlOR/XQfX0UlaU2sv/aEM+Miz33vg37otx
L13X3P8KqoCSJTLqygSO9UOyxzehx9vD7xetQYVSf/9VnkRuxLfvA2j52we5+itz
finK+uv1nZ58C/SFlJ54L+kLm911skn7xi0oS8kilGgV4eN/DrAgtmleVhoKNVT5
OWMzyb15vajXxNXP6OaBUgXwgOV2vyTORrD2A3La0FltI2GDyC63mviIBwOy7RL/
lR5d2ryi1gg2Qs15ctgwLg7fZ0gYcPaVkZjWJJj5UOFzvd9+TJsFbiyFlLmkV/0S
Bzv4ZWzKH0nL6vHs68IoVkWNqFrRwseUtpfKmf6wkEtr1XkYo1vA7agzO5rUuCbO
igOkW7t0QbwURP6uJ6BW6iQ+QcmzphQBS8tQU9FATIcV4TXuxuN9bnuhBIQpMqal
FK8YSb6nUgEcWdE6CxS2C0jWZkdzylOEBWbC05uYBH95MjpeA6zk/hnuh1eTUw4f
9VYL7xav66sVEzsunli9wcRGhsNm7Anw6FH1KPMFfkw5Z3ROrpheGettDqCfG7oI
QRlr5Kw36AAeTyqQM6h6xvBIGC0fAGJFWOnPZxhuANmZujZPGyIgiskuV8O7iE9V
XdkhzUt2897E85nrndb3bUq2to6Z/R4h7OfOI+lg3YgH5kIhft31hsFQGI39EHqB
eYze3Bp89fGG6kNlYpsBOB6JvP4gWF3UuqGdbe+c753tM2Bm+QDymliPAzRvlC7r
CSwZeNWdfxYriei3nm01T6wBqUQTHbh0+6InqdShuGKz8RMN4E+4nZaH23npmoUQ
WREFsaDbcPGuR6z6+S/6MLRuRM2qghbvQ2obLeEoGf1XzDrYrbf3/z/N9fQcZYcG
ESNVJOXZIoh3S9SruFZf+AbV3nfxt0PGib27N80Do27HQjUm5NhC3W/41b5Mdaby
OFRA/qoXR76FkeorCzHUja8OXiwUVuc1GL02BzfBuK5wDNMeOo4eLSuAp6xyneko
RIdn+6AcvgHDwQQxerbLUQkReEJJPpQ6/wiCo6WkoiGXtttVYyn28ihbz51xTWId
b/5abbkyhH1Acf3hWS/02jeDAu9axontYBVo9WCOl0VHtRjHXXyj9Eg6zUt0paqn
4YtGWYI34qGiRucIFMRmXvsFYoZWLiL4QNMNXJf9k0bNjGtT0vOZlPtorU5Z1Dt8
OrrznlxuAQAaknHT4+1mW4JA0bHe5rFYbzSMJR0+lRDMWMr8tT4BPJYV3xDFsiR7
glyQ2C5yIgpjeHHyKd7psbpVV+S4t+ROAb2MgppzPeIT5uLNBf3fFXshF1qju4F4
JoR+hSuOrSzNjNE7WTVutdr/dsbThOMM1A0XMpCl5JzNJmdAqosoFW+MyILTPFCK
AxIQaoL8n8NXSoS6cE/bLM9EZaJlBfcrR8tdFeZNAd7zHAfG6NF25wKFV24exyQn
TN1xkWsht6+bKzq1FE1fymtfX0Eazolpfn4ClZG/oLbFs2D9m8Ey0qd2X+BS2OS0
c0KPbFprc1iXDtg8G7+XIIfsc6Mgbv6YLhP0PfHndltRVJUXvpz1PLISn0qLm9g2
hvdOe0j/OEtcBAijfFU/aQjr69QyMaNi8rnHzA0SYhOQnClyCapF5IsJ4/5ouW72
flLygD6vDY/wdPFLAv7FAEHag27VniSbHUfLCRfAqq19FE7JBSIwWf/agFHQVwz6
8QCuQJKFdo9y+K57uzeMFt6YNNkdl6I4FPWGhxBVddtn6cSuT8/QOKaRsSbRloPw
HjQetApd6k+S0Va6b7MXEY4DFHCSrDgRFYT6Zvwfa68hQbpiNzk6tSxAvzqBOe7s
Ngi7oop99/01/rpwkzCtcpmMgXJjegB9PodtsOVLg7jHshcTYY4oVlP3pPP6oI0e
WAnDxfpSeNBfrKOS5E5g4tS4sJYkF6RkUHdg9ap14K4WBLhhUKKxfjRbCKAosl8Z
Q19V8P0OBfYXVKMZaEuk/v08bouFb4mJT9KpXWj3yfkUSZalgrfWfNJrmDI+eX8p
7AIx5oT+LYFQPEh0Ia6pR5FsKqxhsn7+XmmjHqtlJ/htifXLiu9e7GYIWj/pIrTu
22xRl+1R9uEt1yrFloW3SOIhyL7B1aW5u4L5PaZ7UD2ZmkZn1HAqFKDIbFot5B8b
nfs6PI3jLVaKMuBUB+Y8czOpZQqigLcETWqegB9jPNlpywH28sUO4PWvKZowYdBN
6cUbh5lwUeuYUZj8uj9YNjQd2FcOF7cFKZG4XvCT83khLkU46Nmk+DYcqSjAV7wy
XBZI2cvR5UmO5Jxj20McWaKAFwpP11VrF31+KuHq0l2HOe0Kuu7zybCoA7NYzcvC
IqPgiffN4N8yvZagGE8xwfY3btlmWFCSrgbx/H5Sq5U2vn6rd6aGF18rkrb8zNG4
A223NgCSEV9sqqkIhuScSxVFbj38HZiOi758Un0qDJuwPiB8N3KMA9jx9S1cBu3b
1t3VZ8yCK3oh55JlUN3rzRDgHAVi5FphnNXFbQ7N7OdtiZ1DnoTA23/blr23cf1l
6EyS0LBl+/jPgVFTZbNq+fbfz5iWjfwnnhs4kKrch1vItUlHM31OctC/5MAtOZtJ
3zk0vaB3F0nIOn6x+edI6d2P4mu6wybiNs0p77QjH/2MaXw3V3nA0t2tRdEZw7VI
kaS+cxQYP1lkRiUghPdUYn3ACM3Vz32Omnwh02CE6M6vx3G3Q8dCP6yPy2pTkTl+
M+BvoXn/MwKP4YGoG6S1ErlrbIC6wlwOVgjPKmjAQ/JNpaCm6o8zYr1pYQpIUo54
Lfj9JHCq0q9uzXx/WQrKFQapt6HhtatLO01aBckyv8shBq8wL4iUplUM5SzLppA2
exN+FTTLdEyexiBqgNq/Tlgf6UHTFr4fb9Us+yTkKkduCJz4XN1q66twsjoIvUz5
iCHED4cWf7kkjqpW+woQqnbli8+oDucUIZhnTMTk1R8dTM49G3OonR0PP2kNTqQ8
qQcTDIsVo8eANvzO3o/p/rShZE7/cxTBFSy73ShRC733pMsSuR6V1ui1wzZjBida
K35Z6r69LkY6rHcnc2N+EEW5YVrjWJcaK0tN411OgSvZYGcMdsiOF7JGcLaqhaHZ
Zwc0GiO/ncTEAunAIf67FeW/8Rzgzf8pusedBj32IivP+sc/kYUGVuhxb7GbTyXm
w0wfSMargVR3ixO9xQXLq+eiwV1XE0gfeYBRIgLPCKN7fY4jTubvox68bxEmdsP+
jo3GiN8xMgetUxuqHb1GPdILOqYdtCMb2lthlPfihYpg/saCLgMJeljfMAyWAeGL
a/LM3ZeKrTJYvmDfWbgbiwL0/RUbdPt/YIAiiX3FVlsFlMsm4gvYOvImUG1zEHlC
ZOlyjmtDsUZqMp4Zy+zzfpF6ebHamhrVQWl8t+bYnqccevzPEmtq12X+reTt8J6Y
YHKg/HXn1xIIci9QCkrbDA8U2Sr7QY4M5JrLUpY7DIvZwVLLD/inm9rFuFcqRJ6j
pEhO2Gaf4gt5r2mitxMYsXujrFiGGRDHXCRBElP1MnDzb4WvLp4MzD+RbEpb4hUK
7PWJPih3zV5UCqNFuBa0phBNpgeNz6KXYLADbOAXIC+XBn7O511nKopOfjiX+Yqk
p142//CPBEoGhz+N7TC1sV8X4BwFLkc13NQG+wtE1AlcXIMybNptMbvR2tqSA629
PTNvBK+/sM+JItisCLeyQzFE2HfXwzdOXMzEJD3r6sZdspHyWvvRyGNcv2mrET10
LgofTJs5QM4xrFFEAL0UrD0ZDQFSJfZD5SzM8mhXx1taopwl32StjDKMxkCw6XtD
7770P20aDAeyglUqRlnqv1pctLQtc73TsQDyfnJjveInFSEr6Q2LoTLzwIY/pOrP
pr/YajL4aMgnaGpgOFAUFQXFc4BQwwKXt5HhBRbfk6G4TK88ilmytvP287TVSqDD
U8MGVcK0xw399G+gflPxhzPTDrMIDenYxXKjFsU8QjPfbDUvGmz/uYNh6DnQW06L
UpG57m206eQ2GAOeBcjOQ/E4dUGeNCdAl/E7IVgr/d88ljLeTpqFT/PxsoyvHX8X
fhJwqADqekYQYZhFJ48X9Shek0ff2jxKv+aaCUj4aL3nUnRrFiqVYHeOnhj4TXA2
B1NzJFZNSDTt8H58HgBwYzoWiDzaB/c7giJgdN2atAoyvE7+ruVRzjLfB/GX9PZP
3JtHOzJov90Lyz3TSOaG7xgC3ieTSYFOkN0QxverGHu/dd+/GZSXst1P4nAl2LQq
OP4M74znemNrRo3fRanHOA6QXQ04ll9Scir4QEchioSdj0QW8qWDCRAP8SEnfpag
e21BlY7dau86DTkWdh1/IG9rEeN6/AxgWR+heqOvpL5fxhO0VhCg/aUDJxgIA7Uo
26AYZ8+/wGt0662w8Uz9OcHY1GhWSOYAnYzdJ7VNIUn4rPUu7nsD14OQ5EcBlBSH
QrRtZqOfACUMz6PM9dHhthh3t1eePwjKtW3Sd8DCeprEcxBfi5pWMg8HnuSp9OP9
heTOoMgg+yVjezvg8W8ven31YSJVkLr92U8tMGMvgWUkP87/5J46LpnSyyjUJ2H7
VLAfZlWNTrII6VTRSozUTm/TRsmOgHeTaYWDoiTeD7gJbSruziXrrlZxsOws5WKN
p2TNa039wM0Xfv3tC3bKRzHMk8q3ARaey+zIEAv/1NLrzjtwvf4GloI56/e8398j
1PFAgHWVps0dvqMcRAWSQwck61CSdXvIcINaiR0MtNa3UtXmp4Z1sLjvJjIQgLzq
Kard237noLnCimHlK6CDOSLPmg1zX2UWJx3l6Qx8Cnlz8+FYswPJ7CY5YXbTeCWg
osRmykcK+2ZzgbtwFgE+vGNmE1kv6WtliXFjRhaJ6Z0+EJCZ2A/Eo3aNWcmPEfo+
oRysi6XhBwzuSVVTkbDjAVjPoQSQORVa7wBv92VQm8xBysJ/9ZcAUXc6Dk2d+trl
fMBOM8B990OAREJamSczphtM414+dLru0RrZAkjevVqLXEckv8hvGalvD+vq99X1
VtWai0XHHDxuee99cNjITVj3jTRkfpB2T0nCckdFixhi3/dtZO/3hmi1t//rbrzh
cyGKGeWgi9tDM9ccZ9sQmjrrc0LtaSLZK6EYLxZAyWYclWAt2AlfYbHlrenxtS9J
QFS6RuY/tAZ7FuQNLqK+5RCJzjnn/YgxLXQUJi5SHe7hXmy741HPpuxOXuh2xQfU
gxMcHB1NNvQARnZu3uZxl+Ij5dVooaj3xNReYsDH5d9beJhcHp4Q5DB56VVdBoQq
SIzkOF1hee2NjiduBlOxzRH1sMrjdaiFGPtDArwaQUhhQyHjg1PA+x4HNdsBZ5bM
j6NEupNyGWXK2dVCvetAR+iFg4FvQFf3lYgDfVBXi4CmtN8/cuudJliG8mbmrOHt
35iWGjQiXB3qPb17+AgiMsPMQXicGl4rE7Md6Gj3wZoNczpJYxJq/lLcmQiGHDGd
LNQ5dPDuKhgsQSJ8CnEo7eUIF2vwR5G1Sw5dpADBkKXPBEDZeTnp4ZYqLOAonNlp
2U0QO+qr+8p6jrM3eh9tiu8E/CDuMQhh8a+fz0Gt45j9KRM9pVl6xF1xjN5uigZ5
re1sTKGDLKSPT5f4qm3xLmc7PKzzUNaHzg1dPUpuaU+FjsrdTF2etBVkOGekmmxt
HNyCNvc8xYN437sRCOYit/JJJ3j+PpEPozbUytgHVIEKVVciSqys2C7E4EylEliy
+JlK+62+H115Kbe8XVVGh3CxHVtcTqJhlow+nJvayzrZeezzRABz54T20J5LOcrk
JetBS8i/Yz4g/TUorLYXNrmByjPpw9/g69h2PzcY6AlsTmpAitdPB9hV7jK7FefW
nsRUPOLB8GfLDlCiOHX0i51DvLyPMw+PRwlGRD2hSyEGMM7vfmLBRbTdlbrEGZNR
psHjpcqvxLE/rsf2j1x6BpMpAs3x3VIfr0D+tOqX/SQz78vIlQHNBBczjwHAepSc
hQb2wHUDF8gHCgfdYdtfMADn1AFn1s4uds+foGh2UiOnOj3RcgVoaW+/FOL76n8K
/ySOR6MM3lboZvfePNA3hQLgzYiA1PY7uYiId59X9xEM3roCGXCH0nzHUPKS2VgA
XqVaIpW9gsnKjf6EdpHr0meVMkE9kaFyBZ33wMzhyauuz30jrIgSjS5mw43L1xFC
P6FxHuW9oyz4cHGYCrVSHdcVtlaYl5knBUvzmXH5FFAGaKeD/crgoXvhnvGxUshi
VozrpC3GjIk2OvYCyreHrIIgZFm6NKdd7SoGFJGbXz6/5zOFlUXI9P54evy1j19Y
GC6eIEYZXtUPkD90ErbRUM0bB6bHyu7f3e+Y2IC9kCbor8+BaM8Lh4/DohvtmGn7
PdvuoTjrKHDIvMU0+BvB9z6fptf+z2NJMQfCjv65zsyJFOg37S9J1rAXNZSgisI+
RCzVAjRjqCBIBY2OvdohVmakMwejjqecww/GjK0Jsepa31l/AWAW7O/p/b464Few
HtZHJzxLqShpXIGtA7lL7yaku80d2fd3TGx+tBd9iIXBtL1sIzB7TxjzMte7t1VZ
m1zahQA8xfHXVhsocKMMuEMySanT9/D9SmIcXloaY2e19/BBzBU8Bgz5j7nm0hmv
3yWEwohWOR6f8m/I/j8UzsOEOi8+H5Tctbh7YQ/5CzzG4BnxlkD9wSEC6PgScV8C
z/fKslYgn0k9ZRIWT5zFlduVcWKdVEIbIQ5IXmhvsH1R3pBqxx+a7yKoC0/HHJjI
Dj0Bd2sun6R/dSe++NcGOKXpjgITcVv2D0WjaS3ViMbrZoItFjwogSGc/+gqiHEz
0iNsugrAbCrbYfn4MqyLJoYsooqDeH3TRaXq3lsYM8hTibl6D3E7LHQswE/qzYpR
awFfSzuZlujmSiMYy+xUirr+cQVUcrI8MwzNLh6eayVPu7D3HFHT7su7b1YeZ0fx
/a+KHK8nFbzrf+yE+Fm1oU/yTftywO71NQNwQ+n43VnfbggzAAv4Po1IQMxT1u+V
1ob1xZ+iGbfk0wFH/HVVIJENDVCQM/MtulF89D7oXK0/vkpH17fnzSg+qLAmgX20
Ojl/kJEHsYhVDbCD6agPiZjHxFPQOjWfC3eEpJu22eEEgS51VtO5wi8i5AAvd17k
faxJtTWG2k+S1m6WJ2QLWFSwUUZ/h8Layydjq/aKqTCxBW+aODXRvlqGKqXw6Ren
C7cLoTClVLCkz+AfZojSoC6VKvpow9J/hSR4lTwIWwlsDddYHgvndgI49GdO1vq0
Oh+T+X0g+zyY7rKGk4pIasW9Ms5bVFBGlTeCr5omqBVUq4YQ69toDKnub7TiFs2z
CyUseqKM1C5mUhvhVBYAR5hlmOiOYbx0JGbfUdnlFdInLNZLNYjRfaKsVO7agu/6
4bAFb1RNF3bFSrvCChR3Pdu6UtHG3Z9MP7Z4fQLMJyDx84iXkjRj9NQfdLCSNYHU
JHdI4ntP3A1Rtz2klu3QeJF6kvf/F9ECwKfzGzTMF2B9eZL3KeW950FABbGltghR
45W6wLrrFRxMrZDd6h9LVWBkUrlx7GJSSHRbaDs9fZbgFAB6lWuDogKRjT+bV4Ov
nNve4KXHPz9tzhvbmN+jvMrzu6vNnzYaXFHXIqutpsPiNQE1KFYfwjWb2MnIQQZ9
sGXMSut4gbaKV0Qa0wL11I0nmtej+1DZ4md6la/SmvkkTQMa/bBO6PMO2Ryi5ysI
DVV2I5ehzMh96ucGk5M2TsWdpdeS11t//uLMhOZqLNYEYdc3tWDMQRAP482RW/lk
UAmLoNoJigHQeZ/vRIT+3G30odWIK87uRyygfx2yMWM99morIF0FV4m5IusVItDm
cAuISXWNMbeEkKI2BWsEQs+Bq5CLGPyVVIIHxFIPdRe6eJAqwCdG4o6S273VH2VN
9jWqNk2U9SypEdIXrg/u8H3SM0F1iMDPO5r7coDXP4j7+qygTbi92rOHqy0/aF8m
0fKyrv01adop52t0jxVOdNVQpzNQfnIYR5Z7FE/BQHgTLdr5FS4B17j5rmlMgSny
4pRoxgvdZadeg4xXPl3gy5RBvakqiG8OeUjus4VjsOuhoI9m5MeUtTDyleWXgZJ8
6O7XmklQEqIynGAqhI80fgY1D06SGYpjeELAPtN+u4gcoIUhD5j+bzc/4Y4J9aBd
+qPPeNirY33cJ0F2MGEPfH38rjwaMfynWhOgAEd1mXfgRuXhYf2O4M47izamr1T6
Grwuz1sUIj+3emYpnCUKXxOecKstKayuYCjsN+GFaeLdUW88ozztX7MPJBH+txnz
Q5nJf1mpEdFhYIqaTNQMr3o8lnPe1PBMGz4JFvRKDdyM1RVZ6oUqRjSw2D72EH9W
xVVbMIgr/9hAvlfDeGtpgQ==
`pragma protect end_protected
