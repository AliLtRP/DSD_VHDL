// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:14 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Z1GLtAAirOOPfT5DQOSN/xCydTel9RzgnT2Q6xoLq4WWRL3L8F3oO1iM4XvUK3gB
/MyjFbr/A2JqOG+3rk5f0MbktGo3trnZGDttC2cmb9fZ6EEueVwG3kfkMB7DMPcH
X63JDD04Pm80fdYTpX2ecziHPfNwnP+cQuWTJKxEAdY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 88224)
f7R2pAlkLtDE7FTGLNpJCEn8Qv4ppvfdcKbSD5+mJ98r8bXA2AmPpGlseT5QA8Mj
VJwtAsCqL+mZeXsJ3l+cLKNz6q9+4xUA6x+B1WCK1AzX8KKApWEKNeCTzjnGfDBd
4KXBCIjYYDFrc4573OAZ+1OxjwEVzCXp5xZH3sDDPwYlB1MPvVTuMxWGSSXAT8ei
QJVm2qboFVVbey3LqBpAxpYr3bbIMwwrUq5bWA0Y8A1g5DKSzpY8wGEhsTXA0li0
c5Y2WkziiByFRDyv6Lw0l4EzGh/HSn+VZMhRf0z6/dKgCoAHiEdk9mw4QUvGtO2g
8MIELURU+dOiegNjPEWVIOPHmrldhi6rHwpcQlk+KLNfC2h02rHQ4oHsoK5jERdV
zs4izvbCSwr0DlnMmzS3QbssOJMuPRFlV8PkaoQcRWSlNj8waK0Sq3u9+B4xuv+s
MpBlR4FgIND0NW8Ua8U7I1YOKw0pwYlbPCEAFWmnJnbJVeBemad/pOnP6XHjvTrJ
O09O/yP/2GLmfCHDkI/IYhflX8beCBgUwuhBSHNslvtFEHzAbeN2PGwNmaZacwF4
EuThHPMkNnDK/ma/LvvZ+3jVwKipZmEOSQnk0XwzIHFta+NOKxyreHTYgT+ji+gU
5jiiY//3Li0ZjC7GaD0OhO3ZOhjdv9ly+67U+TWjY7ZLBkUP+LtXvwlCQ6IxZNwI
Qbb88TC5A+OhDi949FHwu6UwoJ+SlGqeuQHqi4kUD0SwmtYeg1rwuMyJt3mjYzlm
lVEaoz5dEMfWALQm4Ce75YBVDH9FsVo7LcSb0tMTDZL0NcS6q9xIpx79YZtzhUcK
VmgylTCFmmSmvOJvGSJPgzNk/1fYaL+AXAEdTFVgRiR1xZaflmINizuzADSRgGcw
Hn1ob+mFmgswPhoOtvgQFiZxeulXqDcCiP7b6ETHCAlS/7e2vsS01UHBkmZlzIeP
WR66Lu8boyU9lKvZkviPtM3RRunFO07MJhBraurrB3x4rutgxvpmjo4+HkKbCyrR
TjFALwFDwiKAWlkK7jfC/9qLMjrfiVie9Mt1P5HVwmHZ52NLHrGlJJUKoKd4R5Vi
5VEvCRKqQUlGmYYY/Y6hUVV8AQ3GegZCTdYTDqmUuPlxEMv5k4/W/qvIkVk2tOe4
XuHucvcJr+yr4cvBhIQRYTGgoOTnKQUehs8N3nxTRSl6zVliHYbXXEh0U5c2R6e7
AiaXH3YUFsQkBmIZ8FIWoWBChe5qTEDLxtoBB0EiI/Gdzukx1nCXY55c0IS5utjV
ZlPuxjxVsJlAedTEgGv3hcx7FjdSDeNWNCvfV1HUuOxr8yefx8go7jvFfkZmVjDs
NPfl0RiaFurUrUConXu3DJJBNWSS+g/9modR30Q9n6ULUhLecX2kpFB4ws6aXcbZ
Hl564cO04BC1cna7PF/4CHKNULbHYNJ/7+dQvKQpC7q4sSeuTqbPC9J1s/kmO1p1
kB9Z2Abo1PgnhYWY8ub5xaiA9FQ08FRtZ2dxcXgZDe7Qr0O2fQpBJg1FD0ExRdZx
923BKq8TmqUoR7h9HnvamuaWCvF9qs8OUvAGABzcPhuyueoNLHLzimfrjYaYL2j5
ObH6p0H/2IdjyMsB15mJ6mODxHsdx1FYOpBKSHex/KIuICjq6xBH/X99QlepgGj2
4R0/0W7zhPv8R1JUBBLhcYybbKJEtTm1Bo45YBrNiBoLC35XlT2G3uSfhk+Tybt0
Ta3w50w/XRovjs6WnjnBN6hxAd6BulGnpCDk0XuKMe5tNrZsRZF4I/ELK9ea7VMl
L4gt1uhWAuNmX8Xn53GVkUcelh+QUcLZJKNprZL/dZN5afZEPlpD1mbyL1FXTItx
4x6tUmTvqO3Qe8+W/AvkQJSYTCFzXNF148UAqslOPGwUXdG/ZwlzmEsCSFqSX4zv
0z4NmHy8VygU6bG0CGZbQcMI1waTbuHq4oHLs5IF4yKe332Wu80jOayHWK2LgHbL
ep4SweZ/eYkEA6yfMfk/rbVxJRHW76YF7tIs1Ox/1PeAZhxc3tfADml8arPCASoa
o5JnidapsRvwOCHNulvsGvbpotmr2T/BvAbi9X8VEQQf+I5Ih9+cs30rlVPUkX1z
iTxvtuF72yJ/9bu1DuaScOV0eoYdJtiGZalnAyi4mN+QI7uPb1uIl2vW8pY3hn/X
LA9KOm4C/JexePjpOq1G0UPQ5rP9F79JIwT/RRfBhBU5rR91gwhkGMergkKNcidY
EHqJ5oTBvBpbtmv+gjCK6C9TsbLsmr6LeHw2vCyaLptQbOZXE2enZ7gVeRfBwW6u
9/6okEOEIWsjoQNj/XI/qO+5yaTUHtBp0V3slAjIBYooKlGxAg4ZxWCvHpBcJcqL
fVIIpotCGJUGnK5Iv4xqhRKNMc3KSTVBvTC9rBvrbn5IOlSIJXMSzq6Tt6Cxn3Vb
bI9T3LgsWJijItT18E9iK4B2FYVo9h+Jumo168uLaSWC6Tqft4LcAgmZ2IdvV1B8
KJo7HqFli3Ld/DAVcLcJfwdaMoq6N/wyKtt45Z+KGptOiLDdhtvVDsfkuBrel5nR
88I02QvbpNXeWJM0hrMiQzxNeFok5gXfmXujwmNrfE2IjEWSdp7zyXyG6LWZAwcv
jzjnBTmcFEaO7AUah+g7/kPhVK5Hrf9PNZLw9FYn/wvSyQQDGYglkG2OBdOkQHON
Tl79FehSvYtOenWoS2JbHsqlDbrLxWKNgITzHzImNBoaoGsRGW4f3refY2681t7u
n9pVxtYQ3yinCpGNnH6r/VJdZ7c0iAhk7SmbJbwhlTZyh9FjHGkB4YvJViTjAW4P
MMneYKDj4Q6zMr40GJwun6zSOLTKRaHQrbhXyda4HzaWBspxynSkkWsNFWxYNduz
hXcHiVxqJy6ZH7OdMRayu3saQv/AZi74ciezt0w3QUZXxRMalrzPSlYJVzh77fTn
rinjRYR2reKX8vPjmJY42x9WI6v0iFH2SFKyhv82he/UXX16WxdIlh6kslP7tNFN
wi9WHSpWV+3YOmFlavUmo5r9owOTEjRnvCdr89D39K64N8xEXg+saZ0jKP/+x4gw
7syqSLNh9DS649iSMF3yuBlXQwWWRUUVjX2T/nQBmaYVSk9aFMQE5pCy8tEI5k3J
KnGUtE/kHWVeZYlwh56g/mONeYn7CoFzMcU5rdAbdODQh4Smz+ohX72OJN2L05Jq
uheftClJClur7Pz8V3TUFsnAkCAAkP9Hvgm3ZzOGWXpZJhK4kHpv8kRlP9dk2kT9
aJs7yH2/Zz9uPUIDKaOgsuggwLHLVlhO6VJDKz2c7y8R1ECtC0jS3A/rC7yr1bO6
56OjTq2e6UoL4K/p3unnJRAnvtNoprzb4qp7JQguvR0q9sgas2rR94YkXhbgiz1E
uw0kpkU1Valv0xjqztCsJUFKKABirhYfTHXx6G7EdObuml80QyieZAXtXyzUIhj8
s5H4QRY5DNRydGHLr6IBLakO6qYTmB/Fq7aDNKOsTWb4hwV03SNAlDVB3eyGl9VI
F6zAoyrKTIhX5BTqy+oY0uuGEWMdkvM9b34tSB0yeuUwpJ4DhfMwBvB8uvhh+2gr
lEisnZ7jsSLEHIvk2kT8hBNWYKwOWSXEGoSDFna/rIrzYhCQq4vqK+aXIyLxQwIN
PYjTr7K99o5+orGWYctxsPrYnelvYKtzHiKAChm0H74gB+uLXcp5+AaJuybrzG91
KLk5GkDCRSa33w524a9Lt2alGvhFt6Nt/jm6G2Uw4RAKpRPTzUbLKqcNYyO0riXN
GdccE8/Wc8Drf6zk4seWOK0i9CLktRVLN7gNpAb6eLienA5g/zem5XlqBVvT91I+
ksGbxot8inLG/VvFOaepjS5OgdyStbDTm8hozgohiE3P1JgopM2vOqJZt7tXjhba
K0CjSHhtXSN/x/BrW7NrleHgp2+f2rLE1nyykSCfdojMNZM48nKk5Y6Zxc4m8+It
PuwQkP7P6AjA4i+s9Xreku0Mwm3jhR5PP6vu5Idow0aw/lxg51QGCBe9demirpSi
y9Lxbh6GE65N0s6worp5nctr4E0yjA2bkXMn7HmF+ZNSo9tW/AQ/RkVoyXfFUIC7
JPu0LtofaRwre+owDi43ddC8L59LIZ08HIrxz74qyZjRUPKVAdMGZAYQJIwF/h/u
te6Ut5U1WA+yxK1yrhGBHQZ4dfgbxYr+9MvS6vt/0ztRUAMFW/fQ8Cpnmqt+pP4q
AoWRxQLlNyMDXauOT2jVgE6J4K2MCS5mhZb7xjVwccn1Rp7fE4zca8f+3D9p3SbP
wPsJVz92GQpB3rUOIfw2jThGuhgeD+RULob/FGvq6ehSGtw16ZX0KgzghkfPjdeN
yllgSCbQ4CbovRFZR2cejvnb8IIgYaKivNmrZpgc4IfwgO/5R5f/3XjHHJ1jEHR3
fh6ac1X8K/woOSxzI02diA3DH52IvDM/6JB1/4K1O1PMEynAWy3IicVq//uOo+in
NgcPZ8isWQVunuW6MgiqNpyryd77wnW9JXO/V9swoWzgIhNHhhFRMUEOtHx2jede
GgHK9obCRfXPsWzjMBrs4ATZsYQ5vNu39c7RhncvRZZKTQ4zMEK320v0Cos1oCfs
QztNUx4EMlYMeOT7V1X4ZL98+bAu76zNZwIJ9eVnaTz93LQBySvZpKRf3pmLJC6M
NH1yHpKLIPy7syx1FRxtimR73IlOQW8NP1AIdixbuRDxMLM3wYJd+gVTlpRq/Y4A
mzpzVVOeAnWkcL8fqMuHCkCMvqnkMkwpyXDpE7+wLGFsKB7QL2X1mDQyEDLThc3z
d6VzF+1eysxwQz3XQSTZbu0c6Lz/qcLT/mo75k2+wBtQBTmkJxqVaGTASTtFjhIO
DdJj/bNS0HMAqQtrO5WzJUenv43/zleflJ9809zL9YPDDHhP+/DTKqod95OkmIeM
Gj9ixAXIIoBEb52inPco2XJORoaYsBjEQJ0UpLjU5OaAi+zuDK31XSm9TBD1MgnQ
FSgw1XXrc0Sa9l4S09TX4xAw/7QhcmyJBTSgxaQS+rhFG/6PgUbd+cVAgjZbPqEj
JDFDPU1wMK2gJZR4W0DEraliD1zonofyUzwrPRm0r3fdd6VTZrkrLqK32bPyoM6Z
u6yugVQdjb6fcQTlTN88mwnGPloYSOJunI/7SbNFLI3pAwhsUNqV0/Z3Wzl2sXRI
aoWCUTAsd3g52h2ykp9NMQNHA3RXFg+aU4qZq3WFA13fROJpEmGTVejqNJi+7Fhi
lLUPybgTcKlM4rlBHpENQ1d/gdcxYQHhGZ+n+4KKwa/+4OigGLroRogYlZe34nUa
iN3gWE2nSZQ+Wo9w1GjPrZtM7xEGUHOObjpT4pJlNZFXHOk+/i6m9hHedmVMc39h
qN71GP6MQVhbeIUthOY7Di0Qv25gNcLYmuxXRtRXqXbmistuVfdF8WLLt0BiUkRK
NXTCyd3MHWEtQmJlRJ57m92iB8dQCFQPdh7zc7LogLSdWegUxB8hqVnCX9GhKWx5
9FEwBYma8ua19VhYLiYF/sU0CTHQE6JFPnHTRwdBgwIdbe+kchWqUIQZzO6hLyXc
W/qW81zmIKkTzzeZgB7bEpjw/cFjXegb2ggFRCeEDxq5L8qPP6rj566EpnePe5r0
vi9huutqEQu4ZVs0g/a8l/fHUqofQa4xm1pgZyNA/2vRH8nVXcI5KUAlvj7RCnip
iz1DzdrhraoSMrJ45O9viML7BnM2vZfewbT3xjtr48tMOHyGZ7aATfSDcncKklRq
0GxvpwKuHwwP40itKuBMPcLiWgC4Mmu5PQEDzXSsj2875oEf/U7ftPZRZJvhWmqJ
S6sMGanDNrCIG3y9MwIHeyl+KKWd304ThvnAkuVO6FWLAomTev9YJDi23mJmdTr4
4yZ96wOkXT83ONsLTXcWKJiDOrIaKavR4rlHsD+Hen3UhTcEMe6FrwQS0KxOR53S
049P9Dplg96M7J0/Awaswd9rZPw5LNw4Ko16cRFulHEzbtTTCh3mImQyNNqVfUXf
CFxO6sL6N6qYoDhQEYtTZk4zDefIYlQbwZ6I0162Yf7YBkGZfS7P5YPXEeUbJWRO
v2gwV8zckkrqjGzarhX8Ts2rN3Qkf0xDWB+b0kGnOS9QdcGUpL2A49f4tR4l3TTU
9S7J3HW8REAi81UWQQEIw2U5BV1u/V0z3D8HN9lOUXb5c7f8tGienvngSjF3PcDK
Rf6iKeGaQqjHV+thoxJxgfxfgCvfJR+bWkQ1sSkhCvItPDqt1mP++30VbwXwuAPt
KWEige+MlHXbnFY1ATFgFYKfvdu/zRBNmt0p5kmTblYAJJ9BRqtIMRVmLj4rQ6B7
MKighae7QQFsesE4jBxHvD6Ku8TdvUJ+1JkPVBrJmyiUD2Mvl5/PCXJEuRuGI0U0
nfnPMcd+bluTdUUhfQ3fKzQh4u8wYr3XoXDe7mUYwipFntf3JfW+0uHowakCvuUZ
p1MFBtgl6mA6mFL7lbdOyrWQv1Pa3SPB4LJ9tLAzOlazyc+IoKtmGbAaMDAJuzH9
Qe+hNyHk47wi349A6tT2T6tkvOM1sRJDtB6r9LB5nLbV2dQKTnSYqOXU7MWXJpED
jRUkDkUaLaI18KetJ9tU0pN4cO1VrrH0Ee51chRQG4McSGsgdp1bDFrkaWImIKqQ
MTKk9sfRQXNfCJdfe/+TTXgeZJFyhuSfedye0j6UnmDyfLL3dga1HElMqxhS7OQi
yaPHtjeCBrCtwK8S7WwylN+JoSfsKSbl15yj2qSU1yoe9OOytfaaOCv/9exHvlaG
Rq8UjzGPX1jypzK5uVyRQ9BrtpniOKn0Zpj9jrQbPPz5YrlsJBjGOhFvUW5dcOoi
kFL2kP3WcHKp/Zu52QS6yE+/bX+bov9ly4OYkTw+u3T0Wg9WM7PIJyvxuUxLFWRO
fIc9JOg+DscvEYkCqVMlz3kl9UVElQCWouvauBQ+Gdvzk+FHa8tsBIaGjtHA73P0
oFPcC9bOhGSaGXXb/eCl6LU0WqHHWQ5qQtQHyfVe2reX9kvSB7rvr6NfS5rhS4L2
Cz+K7iKFj3lw6eMh4ojxrJcgNMaZxyNgUJwTvPw37hMngIgYQRyhPAhvQHh+kOQm
/mK2BqP7B4EksBowuNe+GKVXBJDE/1DFKDbzkpmhXYKMvLmqSYvj5AMLVIdyTa6W
kRkSvROU+rjdslMmG5qpMSSOvxH0TGo/0imjXtgIcFhd86zBXJ4DPi96OgLvVa5I
4TFK5F1LN9pzHSD7ZhlgPjoV37kKcRMl+BRO9VFEqhbooTe+y0390THdBKjc9PIG
e3P/FzbXyHBUvi36JdlvQ2gvd/OmdlMkub3hMWY4nh5P/M9sxV4gzTF2rnruX2VA
3dKoHu5xjYeF0yweD0x7OZnvIxjujcyL4Edbubgnyunvbgni5bV04xc/pEm8QyyL
QvjTg8XG+1BtbMGbZEhSoJwPtahAQij3mtETJhZ2LTbcf7Aj14elJPjK52iSpVRV
kkfDE8XiP0wUAPuRaSW3UVRxHYAVMbW2lA1zDSUIvB2mhfrhIo8UQScelS6qwgAw
kCJ59QtJ/bnzBB3SMHLY7Ner5RCNuvZq/Jd/oammJZNKWAGfjPCKVsHIdw883Kmx
LolblWMzBXcKHN4a7wdmX32mDUs8viV0XORCL4cpi6rh79b+5v9FwfQlx8mwDTXF
VcT3oh5oMIjvIN6levrTPrV6qYX/7eOBRdsHR+E0A8te/+kNr8HZITvZzE3YoVxJ
dY1Oo3r3cF+Yr2LrvmXgYpAm0bF+iYYg44MtkV023IG6p/hnj6MFBJIhR4o9NzQo
pnfiNvDxm8FYQZVob6gBXOzaZmsY2UARpcBJXzYrthKqvEgguIoL7Zz1jjz2z1Do
XB03pqibv33BCjqInW9cpb/uJ0mjrNcwioClSFOVS/HrGszHiBf000Wkru4ftUKg
mkvqZvUmC6UKhWtIjmJIMcV376pJ8Y7kWZdMpoOcy9O7cybulrWAQHIKktFGGcaS
WGboTP4dJjgZGDr0Mj43G5mBklVMbPBLNLLI97CYropvjpZkIBVShis6mtOO6h4l
Q73aQZ4SZS/Qi5NAUugdKZIXJFXfBLpnbdeD5IoOWKGQUTXxhFb4fUqzMEnIta/P
2FnPI8aCM7OzHKwFKSmDYaZlapGBgBlKKX2COhxZy9oGwIzXHpx9q2G/O3Zmffyb
F9iBrLNXYpCwtF8svm5wSn/8gZ3tSfssPFHSBSpK2v2IuY5UoE4WzkVmrnnVqqpq
TDckCT76awMTb9dRi8VIPqoNPiwFSVNxlauJfBB5z8Ea1NzzrMm+aCK60mJ0yDgG
Jrl/X70ov8wWnZkLIsqlLhjtELUACoKZn3loIahXvLS+Fuk/NDJcurrRYrgWcXJH
WiEnMB/KR8AdWwdhIwjeih+9fnnA7ARtlhwhbv0sWmS9B/36hjpFxo7n0qTT1Rxz
27edylwNhbi1VRvifyVz3Zb8Cc/RUW+90Kj73xigShagSszckZA9KvH5v3pa7/K7
WCarj2+XsAzOJDEfZUNluWqMzsV/N3pEz8flViPke5CktpyoU3K/hfnZdtj4I62S
EPWtX7xYiDTxhnW6Yr/cyVQ/7csVZvHKu5Z946hPPFtVeQ9LfZx9/aGi+I2zk9Qw
0Gwd0LpjfuXb0n/5Rh3OZg40qrP7T03rkng/uEQocGeaz3KiXzo3Y/VxVrURMacW
LDt8RNtp3TRlcUZ6iscC7pis6men/ry+7WWjiM83+8j/lk/nGKPVFR6UNn15er74
8q3ry5T9FQNJNbrRDoK1SK2J5UjYNXk0OD7C75OBHSf9JOK1DYZq9tZd1U+PBI2L
tXlPnfHnkegWDsiwurluBj4GPacsClmiEa9PnCDiVjaqcLkgza05lkKJwnVaA/Li
AAqiJGkXxQSMseokLOf0qE2f/Yql1fZidGI15PehUoshyVZYIw+cQ6xGVn5OpC82
xzi8lStidIKq438twJv9yEKKMeZIO7m8So3qShPUkidrkLwApgBWfohRR2By5T8f
GyH5A01U4GN4Ru1IaIMhF6jZ2Xle08+mAQ6AOBNqE6XZB0g+1nrSDKx8cLzfgEh7
clH8zyNalz8wHriCROqsomiky8wA+P3z4ZwoJ38Ffskfssy9KN+gHG8gTja0YvNj
3uMFSrUXYSoH8m8POxXjVR75KQbaFVgSyWKCP7unmh4BB+f3+b6uz81hqGvqaC6q
YDIiiJNr1J/lXxxZQl5v1abLXyyQ27ZFI6/gimWX0WbtnusLU2qYBH+J8Ax5N3xY
C04tJwbV5cn3/u1H+wVwotS2t5gUoGzm09xFF6iV1mjnvD5+Cr/3GTr4GxJu+3dH
54MmZ2Pq/XJSfx6Sq5aoiuz2tk1ht96FxDX0jJ1WyvIIHxZ1CfTuW/jnfJXkC60T
eszMfkw4JRii0PiYTPOo9YsL9QRf+Dzad11ejxhWMs2aJffGe2ZMLaBD69HUxzYq
quIX5yShqvWH27BQ8ehFRAUC+qXLZt55qSrjZBVFrjDZzSe845WgWQHMnJR5lvpU
D+kmrKpqk/kWI7/Yra5quSNu8JvtqQmSh3N+R6a3yLZZh4+7I3+fJ1E6LyNosXBV
sEbKNzmUDPh1s6abC2Le+SqSMnGGMfEjhouEhLj8FREwRDteBwRDJykoGodzqeNI
sj6PlUycVbVvp7w0prCqQPBTHRTZsenkNtOSe6sSlt9C1HjizJmCOuKmpGk8yeeF
vFyYpmwnYbB2olx9diJZNKUj6m9YgduXqIYpRN7SrZkCC+AS4PHOZtka2qt0eOfO
Bacq4A28b9ZQ2fl3/chqpck/jJdOOENKVxOmxxZG+uxtn9wegCt3oXyPA8LnCa8q
zqpehH5U1Y5aYMDLBBem8A9YG8tyUDMNtwei52jXtyCIFdbYwBBxdkvYBnZFLbOk
SQrFw/8OFovG9MFjsKVuvamPCORVex4uRAJ3wQrvc6XdJazsfG/Z1dkfMALTozeP
QJwBCeNzFfmmvOZXwyV+Cpug2BEdcD9eEgtdulRoyEKC659xENTwOvWzBU8hN2Pb
hhQSYd0IPi++MWWCaEJP6OFy0/EcStaQ+OW7efSWVBeA9oXM2r8aXziImDZrCHMj
cQ0/qFWGJrUcmDkUUP2bqs67smLoswXQ9dcXIuivLyfNHbq4W7z8KOQRg24Jgqwl
TT0c4NCsnDztQiDVqVse7jk5PncciSyey4WhyVBVlg7XvniaGJ9uOpzHDuVgS/xm
up59BPes+ZltpzToLBZtrN5jsKqG1QgoPv8RfqJjWlLAsgwnoRmpeNqH98whEYNn
dkBoPK6dRedt2QBoVdVWxJ+vmKYDiaqkwapQ0WycAIPjRVkUYRHbjA71iwZHBcab
GYu4miSgMtsGhitQ5lN5zdrnTWStpAJmjenAdX0cSds/0dtcccCP+jRRk+t0gZbq
paHYA0P9oh9l8UCsmC2KfE3WPahFfltWi015GjQnXUz87WCLN9VGBq6y1+60yBsB
Oiz9zSTpwQlZWbX3IdjPHLBZMYIM4Mu7I61g4iWtBuHTNgORRf4jy4xh9ToOuzZK
UGMluTXSdu532PPa5YlyU6lMgn0tCPFyxTK1jUuKNbl7qwVZ4LWaW60C8kuDmwA5
sjvCVvqrVoyxg6ysgjSlKk5bCHxtytM4If6Mp5EsrATjXEg+kwCfNT+NVHeApgJG
ypCIZZ/vagzvgmfrIpBi7KxwmTa3FYxaoImt713b2vQxd/GH5WhPa9Zr7Spol4bh
7eF8ZYlUQaMmE50PkUyLMcLtsH+KmKwXwVQAxoG0wny8mfJOyxJHzqDgs/yX9yeq
fmFA/ATJ/r1jSPqJV5Z66qjUul/tXgHIjJwHW8Wbe+4X4hNws83xJI0Czv3VaH6N
1N9hPWdSbFS5xEnqYLhcNLWtEiP6vPzE2C8sOivJOcvvngeMWZp27nG4dXIIHgFY
S5apyX+kxRPwN+sLtu+zRse5ZkOFzyvGj8ld8ELKlkXwcPYnYT2Fcu31SS7SQ/7p
cRpderNXPcUen/e2fu7UNFWmLtH+jeXXRTMaEchhyVV4Gu+BDD25qYMuIGZ0CORo
VeixjJjSxDkRPrrmSHwUXpaY0DfFKjZmc6Arc/K3Ap93AQByE3FBQgmlxQkA4Q98
86t2bM6QDg0TEF86WG+3vWgQPRtQ2mBhc0ofYSm+UnvhZJ0pHVwSzMLPKQHVi1b8
SADLtsM0zn84LWa1GCqcTwvrdUfE60xkul1Dho3jCf8uXzpHXEiL2ed2wrBnZCrF
Rc0vrdgL3SPaI5yRiOlKfP+OeIulmRt7a5xNe8DRmqMkl81cekagHzaoiNEsXKNW
M5ce1B+sgB3nwIHHPkoeQlu4Rh4ZM/EmlYzNOE8AcdfDkyIb+GX63Q+ooEiQiJlW
Z+cx9k+KVUX2qR/+7+5kXHRot8oQdELbJfnInjm1Qdh87soqdhOvyT8jazGlec58
l/RYcP7caWZyy5mqjXsgVfYXSYlID7x6mLkBg87ijlY6hpqpH+S7WO69QS+h9ImB
9SQ5dgiRLii//3ssS6wnrO9VdLiv9+kPPJxAwqNzpuTHB/2SRqs3DJW9NDS5MXuL
38yIe7iTKvmnhPRQei397f7J6CjQ4ZZR1717WaxySKBvvbMAfjdoinMcOfIj00pd
xmQq5WRmOYo2IvUsQJ8DPzdIE27qcLKRelvHPa6L5UlJqyeUvBHJi3KyfxCyDwnu
dVPKBvV76j3zkwPKe9WG5iLnFJViOnus4dYPPHEIjOLHM6fMeBnbxm1GgvoBoN51
Ss436N738qewGNii5N3X6CQw0uVZA7KruiSWYZscwsDTCD2UtAyZmkJrtaE5fz/X
CpFGDvXwzoUAb38hvk8jfFy5ZdZccOmOABt+Xbq76g9iwmfGJur6TU3NLWcMk2Ln
dGH+D8XBB15LNV3t+/lcLxIJzvk9vHfTBCBgscMliFRU88O8BfEdSc2NYWsR8mUW
6hywwPii3D5+5Eu2DLPKSQPLPkjtnOsyrYxGRltVn6cCTHD6uD+z4uLf1DF5eJSe
0BfH6ZsswX40NawH4/1wi74m4qbQVIP/NNHns+xhFWwktobD7VTCurLxJWoBnvWn
YPbB3wId0NuC18joYRVXOPjXxEnwLGwsnOTOtgPbsn2XGLFj/p6OemLMeZqIQKaS
nLbdF/zMR8yyA7WGsxu1q+0mSb3PJlw0xZJX93qTxr5lEYYLSnwzO7qLwfQHbl+7
t4+n0En3z488aN5ZN7XgAWHAt0ubQZt+BgEPAWiV+LMeFpjId3SrOC/qFQrGof9H
CHnN2VHEMGUV+fxWrGLC4ShXLl5U04qcW+RnNmFed5xb2SbhaTB51BsEm6JmoCdc
KkfNW/vk1tBDHORVLnhFPjvX4Gdj4FnmqK4pW7VEF98Dciyx+eZr8aNCd2eZjfaF
u9ejmRvXZspluCYR499g2YUBcPczu+O8dBOXR0wSceVdpSXVRzt61yll+MFRMNyT
jZuMcLpbpeQLMCT8Vj7yMvIAUC7xdtQPPueI6iFVxtOUwqpLv5+WexogFDGSDevp
NPSYwWA8MKOmR25loszQSEA/A4PoRSZQDO3fvGPCHALv0BRvFURqSkIE89hvVU3v
cfOTO9GKqzUbVgA7g5K7E/E5bNznN5HLP6dKpNTetVTGlvmSDhoIZLXARAt6uYA+
IiSBaqZjEtWhWMpXVvIiE0ekcEHJPDkrIDw0WBzt1elrq/ppjL62MKLWrPhrB6YR
iINS6QSHPwZN3CvajFXyrL0QeU5oQ1J2MZAauDdhYlZloPbYWpeqQuccgGWOcG+e
V4hZuvS2PrlOnPL2D+03PCCA+qZN5XKa28LL4q6ahJzS5zF8KPflZWR6/JtLb0Tq
HkGbfDk7Rp5+/BiEzXxImTPIzQD6FiOsczrpciK/HnrrR9siRr0clcFuo788CF9c
mwE00iccW9Mz6HxGLkHrjZI0gJ+vql07kTQbI0rs6zmEQA/T1M4fQuuhB1IuEqUB
fd99bXb2u89rHYmc2V02v0xsXXLw8nb4NALHKwwikk1/MmrNrJUIr8yeNAKu5t17
LpxHNgPfOpG5dDmoqj3R6TIobfKuo1S5HTyUUpexRqa1vM9vswJyrYQZhTqn4RHa
X3EKIpj7MJ4p+gW/n8dYebbSyXZJcVSW70FMXQziRqj3sINDu7S5CpdlHjGGHUC3
nQsw9zF3UgvsKgKSlznd0xvqyUdSbi1+PsAhBi7f8xBmQ3abDDDujudVza1d/RHK
mM0Tskq9lHX6615s3tQKDY717Tgd0Jd7qSbF5waeHszea8g20swZDtpMKW71IEyh
FT2/ORN2Tt3lZLfXVgQrZi9EtIOc4mGtRa7u0cOyRuzvG7W5G2KCRkglAQ4cK2Vh
fla5zxOEp5e6WE8bHMekFciDAcmDDfNc/vam7cYcpSQ2U7rY3iohtXGNuyRVMhxu
SS6y87fYXfR4a2QVJkJ2pOywe8h0m+QN4gya096jiDc8BguAuSIv6Q0WrijftPKa
idkPT6wAFpE+z5aKE8tiw4MuhVj6Hr1uNs1k+KqTdzdntkINzbqGtFx8YqrRApzz
oEzCIg/AF/Fv2F21/uakLLgiiT1HbCkB76jU2L6ehsps+OBLEDUKiHqOMBstLGiX
+imldmsuVB7cUqbu6UVLaTmPBfyGVanc1v7j5E8UxPkGQLEJdY5OiEy6JUDiGEWb
uDOKUhwMCEeEPhSHup7AdaiQGQvecOO47zOkA4Nyd3q1ytn08xhLpM1+KWRy+E5M
RB1Hx3e8U8xadFwZ/cjHLxf7k6Oatv27jFqprUkASIfv4cwQwBbwdPMfeiVzf/ME
bBv44LZz8RZtYzdn3upG89UcdSchGdX1YTOf6wG6cDihKUoxiIh5FII7tNt1wbWS
GReiQ6FQVoeoFQyxo65Rfa2wco79kA81Cy/x/oJaQ7/RFx3Jjacf7GfqqbE+sNjx
qDdzx3awaHsZbFdXocKhoEP7+rJ9FeY9w1Scead+xL6LjIyCfoawwErCrIrnAyvG
OG3itY2pBVoBNELstH2c68GLyPLi42hjtIsO9QvfQNBknuYcxvPLvZoOlHWonMox
ETvwFk8Y+h+Kp14dgqouKT/JY6OqRJn8xYKZsS0DF4+1LukZhD8IiJFJr+2uAptD
J6afM2z8stpshq89W5kD7iU7nRHWbW26iXxYWNQR8cNmS09VmN6B+yu+A/gs13ib
r0aaf+wttVDWoHjfd290Phvf4kvldvdJPUhHYbjpRy8JqjyAJC1Ancq6AqTTqm3g
HuekmRPs8lF8RUAmNcCzPmKSNxB4cyfJ9HgNtQn1HQ3q97BtcrKD/rDh799SkGTr
fPZRJZEJl34jwtTLPhEyTubPdH8Ut51suWqeNsO9poVLEnE1U/J/S1GOFQLz1H9n
Id5gtYlmWSaTXmW40X4op/sB7lcRAz95WWBc4qBjNaQmTn/WVoZyC/vQeeobAT2A
Mvm8il1FW3v2QNqKu7YZfEEIuiis7Dm1qmlQ5kT3IyNWBtH5UZLiTCt0SWbGqAx4
YsUL75ThT00sKv2w8LzycBaNfckWBhAu3tSNaItizVd6nLdu1GM1s0hcONYRNLjj
bzUs07P3VkxLcl298narMZ7U15jCSCHnkbjPXDoEAd2nrT4qwUyd9ZGtyuW4lsbE
f16Uh/N766uPk7Zs5SmsPfrrPGJWSaJOxc3STpEF1j0+YqOIaDaXihkr8Q2Oyd1A
LuHlSnu38PovfeA2HVVByzJpnMqG8iqUuPEx3H7nAXzXbL6VmRROsDiKs6jnYAh4
cTMfbcgAwZrT/WDQHbMhAEOEtfzucvFFpVI+bw+39JEljiTv99TXRZ7XHQ3hmQHP
ucoaKhGu1C1R2KMpoRAQVKf+fIkBnHtVuSMu/rMbSy0IsQjs2rbZVJZmeaH/2r0S
y0cYxduup2K7RXN8l6hM1ghKIQfPwLDcTcz0LbQVzKBtVK9dvZjMO637YrQP7Gh9
DSxazq7AVz8ypeADtpFNqQChAXvpTgL1UKshMqZpX8JyHf4Eh6TaIPEAfXRqREgC
OdV6KEFjmxE+V2ptIJnfH8VIPn8cQQwc3X6mOVtRBD6e9o2cDdetI6P6VOOYMn3Y
I1n7wIadcUy4wFnvfxOpcfaW21dQitKdBXklPP+WMGCWD8Mo7A6Oy4JNmEZcIKPE
C0xh4oNI+genHjJFWsnm9GRHC19fjM783dh98doeA/Yermryp9psMcRP/eK4DO1J
iql1ylO3L8j88KFHs4k4qMO3573VTnyDsjtGAunTto79j75ACsyCZlbl6m8rZ6UD
uwH2Oca0WMbUOritV2cvCHDG03uIJ75yt0HsO/n3BUplBtBeu101oLESCsJ//p3M
c4lAs53PqI7v/Rvt6omcEu/9Ak2PV00Zg+Jf2nHwAOF1Ehg/+EvGX4Sw/9AiAoGL
O0o3i7BekPGoY+Jx/ac/gw3LUA+AbRWBXbz8ROx6Th3VX8RFiub4a7BXWIYzIyht
Fe0h3sn770qL8GN4tTEq/XIbMR2u3cwihxCs6hd6bqRmcMj7Oobj0XLWwM0QmgB2
5LX3fNV1OWjlpLo2V6nCgcZTGuNRUP5ZWzAW9R1YMwOYuzFwsIU8RLUcoD7Ovgc2
QWUAQ6QEiwcR5U/FDJOyMSeMH7Dt/XjMbPQJfxpRL9s7S90RegZv6k5FoONEk0nz
HLQpmQTzoxIbQZf5xjjYno1iG4rYEt6sI3nU2Lc8vPpVUurKBFgcKFRKmFF7fL9O
9LqkmHRMfLJQMP5Gnc+470mQwT6LJG1rseWwC7QGYtt5gDGwq6+cVXAs+/Nn8WHS
tUpPrs6fOOfe1vKTT14+XiZR39iRKxJWdgndA1uWhLjDmqHyHlfI9cP5+1SRa3/M
YPO/PSbEAFFotMI8pIUGKRsRPdVbeqK8u264hZl1t0ZghojDFXiNhYOUpqNZBAOW
ZbTNB/u1bhi5pXRhVpZ7dZUyU8Og7HnMHxHekZD8HtLllZSla2qoBbkz8HE584wq
+k/vqOdMlSZCnYgr0/ZGYonc+v9mG0+ml2Y2+/jUArTGr653rWiSrVc/850QAYUP
kyzzwb25Qm4FqsCW6j2l9z1CGP/GGYkYqMOayXLBIEhazRiTf6KKDsEV5H+8zqWS
J0BQxZPSUr/6xsV0z5vOB7NoXRqJLJMq+PoS1SoZOieHhX0lAXobO/Jy8ibp6Wgb
IWav9DYRH4t6NeJQUtQFIHerrRhHvWT7oWrfIV6V6mlBihqOPHq8KB7VO94Sdjqn
puMP9PVQDdnpiNi4/0XJyYAB/2g93fbCPDYkYE14zTECCeITyHL7AOciqvnIwely
vrbnO8xqt5XAVVxJEc373zHzQTgd63i7moByhUjxDqK9UT8CroDlPr2msTzG27TI
V4hidsDC1UZh6DBXyszuKsTeabwpE/BVnuU8hxwxi4ZD4NjwkK4Th4jbt7Mh8HT/
kszFz39D5WjhpvbgbYEEW4BGj0g7SGlvMwPnJB/T2XjEfqREHmtt921QsQZYMzOx
wEhT6IJFjj7Q5L1E7xFCzk7xNzyoI5dlskWt/GB8osLpAcUbFUoff5x0vw5nOM5X
JjAjes4QRheoYXO3WX/U86Gv2758ze8MS+vgEzLjKgrSuPo2egMSExuMmiPR1ax1
hCBu+ScQSvtbVFa6i95GIjeT1YLeuhA1DwkosMqHmJggvl1k+7XOwQSXIvkilWBY
rcy/++EOnAzXuaQKLJUbhD/efCkQrX55htOF7JaCGNg8/wUd7RXmgZBxmW+rL0hs
PQu23YQnxcoFALqzomFKxwankCcGAIVvcwJAClsbaqkhuyki51I7zJSSOCoxoXpv
Zwphn3BJyUOiTLuopymBVs9N9qh1ashtutAgH2frMMi2KUV0oLklGHhKqPK7VeF2
RNzV3qi7BT4GoLbnee93drNEnM8TgpgmyRCRl+dX1KAQ2laoKWabZ+keCl8lBO1e
AqWbONTIhj3QNr+8DAEA1LTIzQkn+eMTX/8ncA5DaDDQYfFHLd6q6ndl07r9rpkP
wlfea6GltL0rHcfv702tflSon56m1wsvigKMpsZNkA+5oDEjjzgdAw5O/ZLsXAfY
ePB6VPTpm+jHrwVRGZs8+yDom6moWYWNSP5b3G4kq4XiWCExUvG+yN4BEH5u+zcD
wk2y6WCczTGQE9fwdoLY4WO3dAxEhycAh4jaDgSklkmunhx12P892SWlCxZUNaDk
hw9X9OfNFcVv5ekhj94TteliXEcJMUoXnF1/BGODMgUXxMlcxq/jvWi5Yk/85Kwm
69moyL05WKo6/RcCNnA2yk9/B74nzPTrbNa9Yb/rZWJrx9rkhF6c/pphFxOp9Cjv
DUNAGnmlbnGOPEnia9OG6BRoW2jPFNvHpi90mZAymKWSrHdWv2vP7ZJORtLmLB1D
RL2Lk2bQ34pJZo+P00PHYmAB2vpsvSVos6BB00HDwaRmllHWZ3E6T3yHS2BnJLRu
mIcjjiKktqA/7hJP79U2sSJRr3+3SYPvrMS1ZV24uAsw6UxqgxeLyFKyckuebMGQ
d942uPVo+ru4bW8opyEdRQD2mfd6Q/EIzk3HxUcjBFUHbjr7LvRfLdh1/H0MjfNg
JjKiHle6P/HKOmXGLLBkzOhWlJBhITU4NZdCUtn9MVkyCHOneQ9SGGpCD5vt/NXx
COHKiulmwmMyNjBOYnJsX0YK6cOFFOuKdkR0dc04Yc7bkMgOPmBoYWJ4nufuPCRL
vKeZuXytvc2QKU4QwHVFQjwxb/ZZ+Fc31BFfHXOKMkAPdKdM10EOL1on9MQl5mJV
jbOcGAjuNJNSVIBl06WUjPtJz+6puH6fSnsciO6DHjJTsxT5qBh4laWtNqu6nfqc
188fQpiVulcxbyBKFx0/H8Y8yXk43FevUPbv5ZV8nKVhJg/CHenOtkEKBiO9U/a0
WL6If1s+aUVmsFUmsbYsQkJJeUfygb7kJs9JFaZORCCwXFh/4QOTPC930TrOOU9w
XdU9/our7wYiPbkGFH+hEodWFOi/FjimEP4bFyxXzUnGZR8d7KETIdpSDyOsFnqi
9rvIL0O4EwhRhUc5zX+5FP30/ICbpdxyHIACDZwbRp+namC7k6h9xmjpVV9K1UA0
w0V/gxvlU1hcos2cq7YqkThriVS3G9V+UUDkT8GBvWdPIHCX0XurJu569JDa1BUz
dV2daSiDp6OCcLYUk78YQp2j3JPnFSTLyReL7mShvxI/sdyrcfMHKwtUpZouHKuJ
0lxQmpgjcCiTriLxt3y9Sf85i06PaXUAJLd5WyUowOROdk98HOZY8jShUeIyhM/9
jhILptjV7NSAyVVQU3PrboQ93Z4HN8bY0teASbHDStIAwQvoS2YgFiU4PvyFQmEy
DsRtIUpvAw2Q0f3EnTN915Cw3MXLgqOcFyog20K7KNguYD2lt4FH+APdj4eFBTj7
u+JzsxUIeWxQBG0dDrjoEJyHiVSl6fhLLK51Ee3PIuxzzNmyUmas3bqHM6elZ/n1
iS7Lx47Jkq3S/UlcHeBLY1DCXmO/OsGaIShRj32b5J0acX8yyiOJta55mQzGmDa9
Y/kIaKI1pG918uK0znExIR3c2GF1yrYbDqOHc9XuWIiF8zj/lnKus/0sDxch/SyU
C3JkMKkHx+PxPEPykz7JxTd91ehRS6QTGfCV9hWodW810it7Iy9PmuiaU6PEw6Df
lsbXDY79DbdFJjOzWZzJPwEa20JQ3HF5xDSWWhPQEpB86qpmaL6mLNaGisgomW9U
otJouQY/lmwqTNc0QWirlsn+kU29Nl+P6KLJ9+jy5EddRE/Rd+21OrvE8QrbVuq/
eN5yd3dBdypV2pQHs7OFjpZ0+kp49a+LZFbpIgyc0+234IHTWK3mBA/gPPr++X1z
KoJtE084eqKR3Vc0Z2fFd2t25/o2OUpCb7H2aovigO+GVEv4MbOIwkh2wMu2Jss/
G7KJxP+x4zLFAFbszD6G2sCO1HgnG10MyOUwQAQJ3Mw/xk+vdDL8jXoecgsZm4M4
nwbowoKhdn99TBKXQTYEbUBXrzpPzteuOFnTmaqUU3a2IpCVGCyZU7YED0in9Ky4
5qfL84dRbiBEuTm6mhFRvTOY+Ocx2fNcCr1EqcGda+lqVp4aN9+cK0po1Bce/Y16
SCzhEtjB+U8yDrF5aHC506dlRwh7PyDyGdWpiNJwX3Enh8v8jkyLWuZEtGE1KrV4
fA8bbuPyL+RSmYITWxERrB6n9eJM2bBBHka8Sheoh4V7MEtCst71OqvZ6er8/Wde
gyNHiIiHL+vkM5fUgeGYsjjy6u2Zn5Vz5NKhyD+Xcqwa0BF4BYX/OMqaCJK1AmOb
gszELGslCOU9gSXspKH3fdcUzLIWK1KJiJH+45g0bX07ML5pJxv6G2YOZojjgE0h
AxaDn0hTzEp6BepL5M0qvC9o1wgOhOWUGg+9C63aqlANAHWQ1w42/gTpRXqJuAsB
SWfEYnYZ9EYETmslTKmCYk2dl8mPsjzcGBEudoGTFnv2OTuaCJBoKsN2Vahy0o49
eLBl7AzGxdK14fMJGzyFGcWTQF/SYzUqwL8Cf3QB6KdKwzc4KcTVmebr1oaZtGo9
n1NNGl4Ru/67Pb9qMncwFzsLDkXwwWKn6uSt8+oGF3qP0m4DEH5GCw2PUvm3qanW
XGvc4yrkmXhwbFB1ct/rjRVzNcCh4orbVZ+3MwUEg/Llzy99Tfp8e7LhFHLqGrEW
Fu8E/XFw6u5oGp+PrXP9hnOfD2kVmsSMLRz0bST07Eh8LqUqpByAi9wCjzw08Bmb
W7sdQKaYdyJcdSjgrixxy7wX/fatzvuPszHA0DmDy4G4FAWSSejce+AuMLGB6j1c
vzICGrC9joIl9lvoqGiA1az+tWB6MxX5fCw1R+albZJJR7wCHIrT5sCmxD1XDvxl
re17+s6EBE0cmn19Ezt5TK5WsdRZF2jXBT7YN5uk8EyV2cRdenXIPuE7afRFcxzz
A7DyByUfeP7JTQnDv+JC7EnnrwQwTmbP+w/FMxiNVhSGMLCaPpTljQ0cNMWJ/++i
30L98ISpDN0U3nkzl56UsFAerJXz0rJeRA9ZogMihA3TUvH+OY7+eZqXdNlxnvdm
mfDA9L2HrWIICqAKZVRqnrJC5OAp7DnqoIZGlYVEM0OnMepLiIesT6E08AR7d/oA
/IxgwouWKntMHe74TlQ5znAjUgz30AXHUmxe2ut5BnPWzAUq/8LGldiC4I/XRc/c
LF5OGuGrma7sjA0JWDKfToYaogHEDwYAX5sSpoWRpLwyA6HG8b/biAsDFblU2eUg
i7z6mGNdSB7OrbffWb3rCGiPPfaO+C+sYNDltb/a4bdi9wNZZkVYl+XQnSvuz/IS
C5fDQoRFAkOPrWvUHTcXp4g9ghcFv3q6gPmjdGKOPbKfeyRAIvh5PGMhbTz29fAM
uTQ4coEt87vmGT2xbfHdjHgrXhoIkiRZwfWb98FVVQYxQjwahOfL/xY4H1s9RTqf
Z+QsKgIPY4rGoGW4ubK3isILL55t5RMOvNEqmzcTm9F7ioxV7qFtr5AoHMmasj9M
SwH/wRyVGmwOmVyebR2cCy3XtMC3zWdNXSRRpfeAbRME+Nd/szqfybjDI4VOMFuu
il8OOhp1yPvkvD6zb1qGThYJGwW9Lyc+nMWAPcyif5QYcMscns9LhF4JJD4pkU5D
tvYIAuZrtE55Gn/ZMCiUWDczMVB+9RMvk2mQE3guEBsNWoAIggEzBeBQd/qmoygA
WmzrfDVKmFfRnT+EgXlkOHu4WoyDaj6YH9Mi+OhHtsan5oqDNgDBak5IX4AtPjW0
xboZv5Z6gZYn7FKhYAIphJ+xFd5TPrZ9A8dcfD07x7wM26zke8sQja6Z8yY+krEt
59DteTdeGwP8cp5bWUbSwjTfCvhItvtrOzPEyS92ymc3UXS03bSayQDNIZL/xjn1
KWynz+JxYHRcndet1FScJHZBQ6aF3qfiO2NWsd6/8RdhhetBU/kEWNiW9wgGW1kJ
njjyBMMIWPu6U62KezykxfqTrrBkipJDjtU8bKCwg4HzAabywlIfGSmTWTST3cga
BjMRyVBhxaK++3BDXDOYLY4OduAGfGmykeZBfiREu7gQxpx2NbBcfq44ZiB6uW/r
Y8+3MtTGrjjiuF/MwvIfzW6VVBdZjMzaou7+BQAT8mmBbqxlgGrBlksZ09UZiefr
MlhW2Pt3AhWDfViWNCGCHl70v+wE8yjQkJKoYtMkJEfvox2RKMXr2VsOhm0H0fld
CFl+LZSZ6Y/tGdV7faKG0RR3UW7f+WUhaLQuns9oR4gN19IYLGH91hE1XRj+TDmy
YEh/6ZnxWlkupI4ycloOcczh52+aIVHv5ZVhSYhJGmWwJbXAsTB6y6fbxZ3Y+vT5
Uco5du82772wWkNaJciQQ0RZhaQsxCJl5IlewIXDDMc99h+5bleudQju0l/iGfht
bGGCSK0iszgo24b71v/j1rKN5dVf9kCYqssEBd4UxzyraCIsBMMXKXID0HpeCRdt
dNyj1j//Iih6gLg9/dDf2leBoODytGlvXmVc58Y5u9K5NpZJiuOKbTmdKwy7P+7b
sP1l3XlCoVXYBHIL+8qEatjNNjhH2zhP3fQ3otRHPQASlWKv3eprfGb1AYnVQoER
uvd3nH4B91VOPpVqbVpZSPvSjlMlYxYoOoAYm0zHDrQhrB2GV+uG1I2btEQ1sfYO
p4I6DQfoJLeZ3MjAw3NqYljp9I0Mv5U7ae6/VeiAKUODzgKF4nkhg1stl9XsFI3G
Dx23d9RJuCsISXRFEKqM86oflOqsxaj5bbR39hxVaJ+pTL3ALw5UJUkDoKkAqUud
up1fsg1OwID5HtVeyBQHPBKTviwu12TTnCFSH+uz20xRjM/2FTb77rpa2Y90tFh3
rosaEmILH4rDvQswD7TkfskX5BOuk7K5k1GAHsLRIIv4DmF4gkPdxwsyKitipBpw
t+R2m1OG78t4OUzqCi2C1l5AggKEaqz/nJFWzzLLUMB+KFG1Cllnlw1kTU5hpxCe
a50Eb2BEbQv871NnErOuinFCeet1mOtwpcR8+AZYu80JjPWUun6ofJVa7crocr9M
zE/7ofSi5130BUfBwO43LtRpaWB/LwQ0CdOtHwFIu49PpkDdFtWOv5+yCAJWCimp
WeV+ZrZaTApqlWcW5DBeWmoyM37UiX75fK/57s5ryrfjmb49byqbz25TsFbZkh10
2BQnKYd6LyRoa9Ul0H4Ti0XBjZb3CqT/D04FuUiNHPqQMxaumkn1DW1sEl4NVX/R
MQuyHPkPZqUJd1C1Xt2f22akf0WmRBV6pllwzi1mRdg5HMSh57Dd75X0k6C+nJnB
z5vCWzjN+y4ZSTDO9ODbi+NbVnzdAJ5wrU93smkoRXDD3PQPEwsGnyUrzJTuppnc
8YU5NUwu4p5yt6z8p8F5Jpm6piNnwR6o08vs6VKIkukY1EXr6oqax0yVXfTIHqgE
VqtdwWx8NlK7L/Fv0XCR/l7LP7b5QEym7LGYRz2DWRyJRWWcyZJipVd7Aa8HHncl
YgtzYReWVwSUiR+EIZkW5Qsie5gVM2hfz3KIOfETjm/WIGiivpinK8wsQoI9bCAv
Xaaad2KXI/0y84cFwZ/kmwUEKCunGOsYd3f/tC7KDlYen/yqdoUWMSGBSiYS5qRA
1Gmrcc+ugUpocaUPHtTdvxQ8gHDMp5WLPOG1Eu8V5JrRnZjxQaRiyxEC85S0wpBm
rDV3xbmieNUvkTlmH2xZJRjNEetpt/B/n3rXRkyFT63mP3uzUbrHZesNlE6j1EiL
hoKP7SAv36ozXyNfxmGqBZWMTIZQs2dbx4tDdhzZhHH5WAyTs1kCIRlc2OKbwmzh
RDzA5ih56D3dV+APlC8ESU/GOrWnu6rp+vDSrnP59WTOJf/T9T0Jht4HZlHS/ZSw
phvl0jUrTQKAUgrgK9XJA4xZOix1vYXBB3JfQSZEObDE2eI80vLqt8dkFcRIcLeo
GTXIeF+AqAw5NsI3yBK8u5clPTzXqdc3KvwMhQ2xZR0z0oSuvN6ybalhGVNXEmF9
Sl/0LBnsFiV5dTcFuDmp/l0oK6nr3zBSzhcScFoXF5h0o3TE4+OpnUodtlc9DTWs
Y4/tMWiN2xQdH4N3QSQFjwYAyxaydkJvFAmWB6jAhXC/FraPm/pr/cCb5gu1iDVv
QFOoWgZktQH0mou7106Tt7uU+2BWkLvBIX4UMgLw25ri9esu9kGRcmxHqnD9EKth
du0HtHVuscNvYiOjver/51+QMVjh9/fDwjFccldFIO2/gb46BN68M9nT7y/4JESt
fdVtE0qhkUU9BZ2pcguGOoTW7XQAv0sezlrwxbEUIjJV3poj22j04hb/OD8G91Ge
mSkvSPR3ybCijuFC2DEhWDVVSU4f9FfhyM7iSWWRyS29tJSePOYhp6rzGbSoTG9w
PZMVBCwmZbQZybuX8e1mA2zwd7MHhe+QEjmyILeaTLtedzUamapgKpMCzq+fnCpT
7cyyIRV4kQdi5ngACwJZK26aV1AoHCiAkckUgJMH4yEZTCOZaBvufrLsIWTydvmZ
rzcPUBhGUxdBIbb8wiFsGMbOBQvcA+bio9yfeppm+J5+URZONxzADk6cQTzRP2ho
lCTTgd6AvY/HL+6yz/2O3j+VPFRHXPfmskl0FOyw1nXMY//0yhH8INmiy5IBacqr
/mgx4aiiQnfYqaK0JU/wZ9RpdbY9rKoAPjpqMzePL48QMfT1FL2FtjSFrvGbeV15
KyDFoN8SL8siPb72gws/c6ATzNPDP4Kp89+6GwMgVsnr581srNHWiOXpkQcCEdFf
aOLk6pd4MxtUoubYpBmYb/5HyoYnx7cW81ZZcxBUvtXR67iF56PjbjKpIdPXNv4n
OC2pn5McP/43LVE7HtGq6nPGhLXoVA9gcqh3F3zaLuqAmr0M+zq7GEgqpAFHiNhi
QPCSajO8NrBV4S9L/yiGvD5Bl0/kF21STepmV8CPoEtzKHXkkQ1B1vevqGnJQQcD
2xdNHJpw3fcGQsNMGwywCNjgSBbTqWS5nBfAzf/LoqgTAL/QoCXfsfC8a4vR2KSV
ST08lIPwLpmjv7QmOaL3b47rvpmUdAteVKlQhAm4wdsiMpfIyOm12D9uDeBZLaCc
2tqnVNbKYIlzZZ036/KgRxQisEwqRFETjkhNUH+YJdvciLjEFa5ClBo/GuGn5HSa
AaD8uUMe/PuAS9eFP1Lte16HBIfghXyoRjRFzl5EhYksTH9gQuInSoUzE6eFoB8/
1ThxViwa+ylsMK+CmMCxYfl7kVDO2oC3rA6ANC7q65w/lyG4OYS62HapO2wHReAP
hPYTR4A3faABMpHJzBn/tyJ8rCbp0y6HOE/addmg0tuFwwwIoD3iLvWtFbsKeY9n
1phDhxAI8ValjoUd6pMfTDtC+YMOjEPKmZq7xW0/s+G7tbFT4o1fELkIarU55lEu
ENKJ6zNrWZ4gCiNe02htSO2BWJwMc3B8NQe9GX6Ej/aUuzYwr5lsxgt/EPIkXEas
mS0UL/ZcgyZ2Kxuv6S1Bdh6jPZCeeSC7nZ7GIoWl7Udar6B0s8U1r9lgLbgD+5fU
qIfBDdw9pqjBC4+reTIaYr4uxp4eWnK9b4XuSON688oHyxL6pqybVgl/5A3DfsdZ
1BHXticF54z190HEOnY7E+0LUZ99eKyZ5rpPjE0WrDVD004M5ygPdLyu/oKH2BuO
UQ6M+Rmts9a1qX9yReUJXjZAx82vP9VcTLReOX0ivL3RK6qhL+Qk4OJcU/CHpt2A
FXcMa348xLNzWEbf1hAizg0Ly4TcAZ50IzXdFFCW6G77fok4CVjtiH+/0wSOhRP8
k46hg2ojc8cdZP2A37sjMJ7S6kgt16VEmV0oQtegGsUmhmhCniV236JOacoux9hg
KBSMBke9OBXbw6q8+LCojqhn4Ukwc/K4dpW+/5eA+4X0Ivb/R7gPUe+XJ4nDZwxO
OmKOw+rLcemySRqYnp0bnLlyAvdqLajr1Zg2C8Jy8XZweqURwfs87NXzBgofFfZC
jn26mdVTK84J4y2Br1pd4jX1CdGbKoBldAQCEmif+HJ4UU+dqhre1j9JwlkM7ak/
9U9KL7z4HIpMexCwSTzA7mqCdniYRHRUq1M3AXpjKM3rqlpZByIarJls/HjRwEsl
FIc6jcL/cvXqMt+kt0lehMqq2yCoEEkNzfVFWDorRV/S4FxNyU3hW9s5ZfkSPRpw
83ijd6cxmt1FDsLlRZDVrPypnqS3lcxRZg3kC+Eowpxm1d3W8MY2qnPFIdv+RpQK
tAiHcE/Z52hyLGu/BIREuwFWO3mGg40fIdq7VxTCvWMFah1HmhuAeG18d3cRgij4
yKslr/lrxzG4yP3ZABO1MHqJrSv4FeAlgIOqATCmqDpWtaBlJLmGzmZowVzirfMR
gUwcrpTG8nZJxhBHlrOUPx6Mt60k9qa59exnssSifXLbZuWPYwQ0JahZoTGyh1Sc
rUnDIEq3HIlZup1SnziHiNXcmdIrj3tsElNHD0hCnQnyc6K5dyPM2vqPb/VE/UDx
KYrxoJx7trMyoIPcr55I/S+vvyHcxGUCgnodgCQmL/6XSJS46P2ObaBYhjFQzPnj
7M9+oDxFFQqH4Yk3UdLp4ozmcYW4Xz/U2d2Ds5VlbLJBe/aiMytuGXT/myX823wC
17dYMLO27xLafxX5hHlSCoRWRfNc//hRuX4ID54IQPl2EiP1FZZAVAvCohJWFJCq
2Xf3FnjXFEnfERxvD3vo4JGVsGJyiI9E2ubYow4Llg/4tLHXJO4Pz84dqZ9dO0HJ
XwukvpTs1U+SdcYnXtX3HzpZhX5RjiB6nA4+OdjqleqnQurPdXDdoGJTV5ojRKl4
AFluTUeoCCItJLWeov5wnVONBobbd54OKENqqk1Fjg87kVBbxIoUUcIVfxOYH7h6
V0o/WAGsTI88967/uiOPAxhGCW+gZMumi+DIMnz2DlKTRJAQvz12sdFZFfwfzE13
t2o4llYMt+iJnFIgn+kXyZxUQy7mxKHwaSWCtI0KdOKLObEDBwucFPymlF6VWuY3
cBZxc4DpD62HY0/t+VR3aPdbzrSpxcharTXZy077nQGoEZelADY7pHb44vsds8gw
8pC+VTkdRmRKsu3/TuOlrIfGVMxnaRI6qx+499bSPoVN61yuU2hUpOkW6ma/+1Ne
bU34sBqS1h7d23IyQcqS9P7R2kFJarIRSFwBhJPOIH06ZYVNjMXkZojI9Uklsol0
0E8dS6efZLxj4913Ro4yINRePXIQ3mRrjV1HFFwolxiczUB41bLoaJMm+4ScbseA
qux/Ua1UJhVl7L79iuGlNtQPePEdhgwDvBJ2Cei3/gRzQmBaLHx2KdaPq3Rx0jOn
QlRvdY2UVWjs5FMjX5LszImyhyaUpX8G1cL4RHskPrpgwfa0/RaDp014TvgkYQ4B
QoFvITuWWRSA5t06l5VDkmcUJhM5sWyHsMSGbCSQl5lUlcCo+4WttajUkVuGIpMq
0ca3EraxrIYH02VWKSFKVTwLE7447Wcm6oJldmnu03Mk983/zioN/MG42D5eVT12
kEaNUMIS3U8+RPKZg7U57bmRLRVCDR2EuKsDVlcoIeT2yDuG0a4iL6N9NHN75Aqw
qC8Z1ttjaqiKuFtQhgSqwR/2FQyb8XrL+mGnE25LhhuyhGRivFSsLKKU/RHLbnSe
sYz6OO2UUl5Dis17ZDHIl1H8CMWEckjkwXSdsNZFiY6HG6iAPZT1wsT+VgleIBlJ
qquhFF0AJTvR7sv9SVSXhbQRhJI5gqe7FyLecDGK5tWEv5b3KwHkJRxQOo4cmRrf
LP4XuHMrJVvmepd+TiwVxE5BaCwN7d4ys9V1dWiBkriElh4fP8kAzLv+p2FZrPUU
sLOS/wAEsb7ORbIegOGge6Y6zND0BKodf07QshhNvzqFTrAt2AoYIjS4gfGbFXw0
1gOk/LJBWIGtbPI1UQMwYvm3yWGK0FJuNvxOpHCOtTZTca+sPvtrSixjPk7v656B
ml7QY36R+JRurGZ+SJGf4Xbnwz9CEm55U+oKTVpG8WvNVJxs2hnnDtyDFwfGmpu1
GSaW+tMwYE3MDDrEVJJKsR7UTxCUG1CKwB3B1KsWxH0uIBYmQaRD43aSdJGMOwyu
LDNq7CspSGlMNsjiHQvEieFYb+UBT0rUhrihyP/Fj9juvAgfeGax/s2ijCwSLQVX
Lp+xZdruETs4bAGqM0+rpE1GCPIXMof4OomtGworfUKBWbp07oL3HiBKAPE+nwLy
uOGjoliPNOlBpl8O24Emj986vq/03Y2Diu7L66TxrF6wocOkH39ovB9kKooYgn45
r9yrtBeEoYSj0YR9+XlHKc5RSdhSOle77A1ckp7UGOCQKrliGcJ6E2XalH4aw0uH
lepwimVCFdawlcCuF6g8BOc/4Z0PYhXRgyvsHkRRll3KgPwjOpdZzApHQbi+KqG9
A5BVveVWaRzYuzuzp3tv2E7au59Q+aASjS2N+VMx7GU3++rB7FLHs89OX3jjoLPJ
PRI8loC0VZWhseKT+DymxQaT456iggI3gcofDrmks3DmsyEBh8nNW/aixQEqHi3Q
YeBvRxW9RdPLXHMaU/JZgKFCAemUMuc4Md0/EJYrUcs/wp5J5+gBLij0cdrd7ziQ
sdXsNLZZ9t0PyVAVqFFFGPftb8eT4cCxHQozLGKESdVuRuGfI+J4W9+sbdRiHBDJ
JqyfAoQNIqijZaunKUYH9HeuVmFPORW3n/OJ3AEhX0P6D9JbR2n/KRj/9vM+NPWw
dYyKxznd+0TJgKd5mo6/zxWGQ+STU2JRRdTGeNvEobFccCV3nuFLqJrlhsgv+5hT
8Ww+cOQ+h0HzXF35v/Q7g31YSaOU9jO44ESe2elLWVfAYILKAjoEccpRVxy+s5a5
iDpf0eNy5KP/wf1C1PyY7j/l1SZa/3NxawJ1LOBkdNdH963rVYGE3+h7SvGNGC3L
6mlN4ZAFPleg3WUo/lEvSdwoKIR23OdKPt20+Zlqw17qcMbZDXKIBJrIVzpseMBI
9gt14TeZXyS/QznF0MHfXL0gDUlVWw3dCa9p42nrfxIYNl2A3yLprdkDcaX3qkGh
5MX6tuEt4+WTuzB2R4BJHTcqsZsCuK9nbLvnIvuLeCugVkBgTkMHs44Iq3ayMYSo
Kg3kBrgt+0AfzJWAL3Rcko1bvaDM08XO4bIwOn8ZjXWpK1jFj9M6GprwwViAN4hq
MGFuPg++k4+yjeYNI/ZZmTP3JUGrEfRDYnXeMTUmT8U9ms1+S2/PqqUuejw6wDGG
CYKBMHmAHFqAf5i+RPzaGrq64V6v6koda6F7pJJfOeTxorXhiKwaqCWxht//DOrf
QquzGEXcaEjfadFRv0rdavvvS3ZCV0DzH1miLP+cZ5gKAbewg73qI40X+o1+LYAD
pKWcRb7pwZCFn8EqSO8QDg6FjEgdzPPPgx3WRO/usk/RHo8C9R2z7Kkt6Lrk4Kvo
iV6RMt0NDMbsGs3sHQnEHmLLUJVwz3CCmDjWXT0eF077O7h7kZFoYENax0Xy8OvV
K79QPU4ijew7ieF2Km2mafRayvC5w04Jk6U5N8wTjEO8ORFuJYaxEjU0BIioWNbZ
TyKxtgL5UUd5gFfBTxc+TS0Q8zTy/35Xj/GU0R9lO/et40xi/4UG/mblrQai59ZP
HjlqzKMHFtzJr+kCQ449k/9FOChlE5vVcSiahWhHoBTbxEvxoJ7TJenU8ygZvcWV
QMLu6nIjXKnE1ZrJmmqnpnwEj8xSfRMd8ItdU2XA+7DvrJunqFQP6W6usLZrX2XT
PxL2DBV6iC9Ebhdt1lT4s1NHRZjYtTy951/g/6/7E3v2NWlTqmNkt55Ds48RWQZ8
apslgUjGXIVZCjvCWnOnzMgdh62KWWcGmSen+3foxWn5WMigHSuYbTeAQxrdmKMJ
Sxso88jLXOu1K6uGLYJA+81Ry17dfo/exxpRS7/Si4OQ8qCSgRtfQKXFwBzKAjG7
AmGf/c2Ux2bpXPwP+OU2x+S61RB79l6knfPJZvdqTE8Ul5Vi3LHseh16xLniewvJ
A3faunnadrdm8k8/qtEQE9DpoprdEJyQDtwEkMcrN/cvXiEGMcKDfVtf0XMVD1kn
l3uwsUrMA0O8Is7OMmK4qAUjizF/vr2vLfH4xU1HfSoWvuxH+z3ddIpw9vYpyXTt
nFp72yO6iV4MlruzfesYwjN9MwNrKElsDD3pdw3a7K6Xjn9YaStzz6yUxWcoNGuT
fHQKmnyIA5gKpB1SZ/jBqmcUIldzzMhhbffgs5ohFjXcwWxXA6CvOqJibxdrdJl/
PvSvi4nY5HEZBoizprS8SH2NjFZjUqlPjAhNWbgH5M9PFwmapSDH93m5n2jajHXn
QYHHHhqNeChpp7lzkg1R3Yw3VjSKYTkU0KKsqyNCgJBblRmHDtMGT914kh4sRMqj
WbeSEhpOG6KhRSkl9Ka3OA2JbY/rXwSVqdkYJ3TlRplBmWzW7JNKut1B8OOiY/E7
ncmhJJSszIuJRjYaUyF3GXonO+MjFOxJam1bEU9N2ZIq1pNm6raNmxnDnI7f/z7p
pLsPeZjAiu2jMCxAQuutGRLilEV1jrt/xW8usWdKJioHFUASZgeXegWDtzwIEsTr
vUJqDny/4myMhG8kGCPSDRZ1hciJBzWD87WGkJarubLMDHe9+gbzLVzikajqIuAV
mwpOsH85yB1iWomHVsPceLRp3iW5fM1igQR3Kp6Adr13JU+qkotx2I6c6FWfir8d
+JX28A6BM7p1QpH4XjHcIVyE2TLs8PUfyR6uC0AkQQsvRHKWcdevrmTiduGIw/iQ
pFjZhndnqkBiBL0VbhTRnVYeWVyK2ImvgIG/CtYX/0PuQOb9z4ItRy02yCTXaNSE
R2By7DnbKqLZeqTHQRL4pkNdga1kXkLr3hF9B2tmO1cPwZCrsovqSVMd9rkfP2qL
oOhiSbqS+9ukitZs1uKWKegV/tkFe/o4jSAuzcnPKtlk1ozD13ABD5sXCtYjcL+y
n0Yq3cfwJ7uTTNtRdlaZ9oiFwRSUi/NkqJTv7q8MZpsits9MZEjlOrng6zndPSEp
9y6ms4UNZgaSyoh7jIZjdHQcbUgq57Z52acEoloQsG1Il1BH6QjAOKyDiKJVIlEc
mmJ/wr1EcIBBJgvMTyKJP0vYR7G5NBppExD9bKRYTnLEXGcsgjImwMHCkGVIv5fr
p+vgmgaY9xfBGHkAjiOT+7gmD5sVaEF2Mh1So/oo9dmdHl+lsGta0L3UnzcNW1jA
yABN32B+728G04hO8IYWYTtTZQ4BJjP4u+ckQ+NF5SbBN/UAU+p9DIe+AoV277Mg
x2cSjvuwozIfukRyL4qTtEx6Hbq2K1E+h9Zaoz6rI9SAVstR+ROIcSmEwPJgQifv
QeteHRBFJP1cCVRIzfwFS+U2idTtiuvdA0BouehCFgWaQAStJ9x9XHzyVyB1q8Qm
pKmqK74tjmsUzjllWJhI48eYB4n0w4rbYiemRPC0RKXQsC0zwU/Fa8o9GZUGy9AZ
NTWfF3nf8i9kg7g3BiTErx1bTxzSlzM7PfvmluXp+ByNhihbugr89TbRiHyCkVxV
UFqxoYW01sjo1X0qsC4oArEM4NgEz3j09m2gpymcFQxk7lsKe4Dt3AKQm5WBLMEG
txeVT+3/204eoQqgOJJ2ZLvEMXdjxInt4TDBjoxFQW74gk8KwLxbaEIqM/M+Pd5U
ocFnNFhbnMJhAvZb0waG5vGA80i56Gjr0yOdOQ32B5h2NpqWoLAoHftHVosuRJfr
dLwKuU2kTjK2dczLM/Qn2NDRt6yL+2U7Hd+h+6ovUK/ssrZ7zTvFcm/9t+T1NlLM
VPsGLO8rd2Dw55qxJIf7sXmJLDNcLliUfxgixnGOuKsSqmNHJCEbJli1+zod+ckb
fP7bES6k/RJPj1/dKxnQgqUSVg1/lVs9LTwPxi5eYYNNJ3stTBQsGzhhK5omQzoV
GIJUipSdcDVZrfx1o22k4gqhEk1C1ArzOizDaDXel//IWotR3IPJjHNA9BIkPT7S
p0iJ5BSZfF4CTNJ0xwhCMXQ+GifNsP/T3p+GA/S4JQviv42ikjnQ6+RRRqJs/Y0a
RWOMgoDEk4GZzyf7wD8jBTy4qhDx05AHpbOsP37V574XnSiuiNCKEZsn8F9KHiiz
mDgs68Ym6ttlcRBIhGF1OhdXjkTlHRU0GXJRzblTXHr/qEj+j/SJUVINEdnHYotf
U9AYsqeiyn2/tGieUew4vyrwgTeP9lDujMYi0jCI6JlUpHHVvYP+83T+Z7LA8TRg
/Gg2CCFOdphzxpaXt/yydOj8E1gUnxv7q9lA0BlphZgAZ275dfW6Pozu8ddE+Sm0
2MEGAO8mU2ktiQvOYs96EGOX3A+/b3xixdoRfqyn/QngmYFr+7WNrvKLxw91K1PI
NveFfXQKXkXNvdg3zbxk1sRtCfAq8Rn92bgcxnEff6qg4yFBEN6lwoBL9pSfnUdf
d4yjvrOsqZuTWQTUG41KzKCt/9Colt7Hl6KHWei7kHsCUDcJrbdgRQ4YlJh+Rcb4
QtZ48HT9ktE+9O/yzTUVkMhnWRVNVgOtXhxAC0CnOQjPQoZsY+yhqaGUbOJhTG2z
tQcOt7CkQa1tbtxSU9gRV6OTnXCYcPjdJnIvgRkiey1NSdbFOpOodR2DukYP/yXW
YWY65Fqzrppkwu71CfeSUuOtZqHCANYv3XvH23fq9po2AEAtWayUwrFMb9uhkRiA
1XRk1E2NkIQ8GD6Nxe1a+OAL7z5cuWMKm7fdPX1ep9srOx9IA7XWn3hxHf/4pgHR
aOs//PnqzS4aXSxdQacpe0IXfj6dcOI4X8TpMgIfJ9xpKuPNf92qKdfPAc+LH3Ot
X8mjN777nYM7wfTu9Dk9YlRa0nO6W5ye05vaOhy9uuxcFdV8479aT9JU7Iszvyw0
CE3C1E3FA3pGTuFyZG/pZUB1SwWIpbjYHUOKq5jfIoCvFBC4jEYyDdPm4GKfNlB1
oycIEzoRB1t1zFLEh+6sfmfOTAidst9qfqX6+I1tnb1kOPu22cdtwk9wFNEqRfMN
WIQ77LvfpLXlbdxkOhGeC8RA61/gUxNwHk1vl+6SBZCWgzC6Ihp+EVqSDu/AMwiP
Lxop/f1gSlrm9KR8t80AGplPzliXqXoFWpqlLVedI5srfnM3dfCBGItoP0jwmYVP
fF5DnHihNj+peIWubn73aAMJN+myG51QB1RIm8RBQPX9m1Z0AFyTmBnBdhXeLJ4C
xhYlgABGOYNHbYIDPHY8gZaYsio9FQ4rKhDNJwkN22zEQFW/iqOuDXmcS4xPUsys
+zcHANO8Q5DARQjleCbvr5P1h7iK4eeLauqBiNkG4YmOJtYzSMdqD5hituVIqh+j
GddC1ST8T8wTwxqIJgICsc1mmNaEVDxXXGvJFZcxRunCi+495/JF66yVdapTxRln
o+y+AStyR46kXZj5YCzE3yM7zXK9JeE2/rztryeBM5OCQNJNjDU34FQ397pHBR0F
AbOxFYtAhvFTRcCm44s7xC42VUxLoiRExybEdQnb5S/PnMUarHNMlt3XtrdX83VP
Xh2f32CkcadIOxVU8qJ1fbdst1roGSULbZiCRg2vuEYn3V2MPdGLS7HIPC+fQKh2
9n4sEFnghUW4G8wb1UOYCfKeg/x4HVkP1vi4Zl6a6J5LphrdWpcDOAsqd541wmMf
K19pZeXP3wGvDVa9Maa4Cag8BkWt06GH9iBsfd+lFngeEchVZwbwlcnsaPeOeTwS
yPO3XKUhuHeDWDigz/0F0H8NgX2AaAr5ojwoQMXhUcBFD3sBAfB8imYQea7S1jSZ
HaLaL87Hgl8nvFwAaTDLKFSC9x2Gf/GAC1YzBIgKvgHfG81yMNTUdAK15OheZ+QM
Zpt+UNORh3JyDTQdbWUtCEoy9RhEiADHAwKF8FFEpU1VgmMJVhSEB3g/zgEQvAOf
rB4F8mSAuUKN50rOUjYQwtPjDBN0jNZv4lPwdMxhNmwG3La7ffhVYPus+qp9HceH
PEjenrXBPwDv6nNhszM4UWurF90xqLcgSO8UZ3KRluRQxUCnWLrWnj5HKV/OGBaP
GtScYWHo2wJg7nEPe5JPzEhdlBEcpsafhygB4ysge3OVV1MCuNI4kalYQ1d85Zqu
wYL7UkbK2QWfU8Gn6/EVFz6+BOeCk0Hox1lsScU2QsslgigjJs73jL8dB3Xgw8mp
LdNkt4tlIrlTVJzxSJDqawQA5ji+dHauD1zOA00hVOBjZTEpwyKo8+ZQxQ6v85Y0
QgVMK4Ehh/Y6bvpvLkREwnHpoattLm+ivsgDZQPHKJlyVeJsJZrZYLScrMEY3NhL
FL3dZSnD570SXwPL33OI1A0hS62muZwC1mhdWh3HQvIGhETwzwuQfEVu2mWZCJ30
P6HwTavKYfU/Ozp2JYjNWENLefZoKMilelJQ2bpq8QingEWudDyjiso/yKF0kfx0
nm3A1rhQVKMkS680c89L04HfwVnl7lQg3bjsc5YPP1DOqIEtGJuSOMaGXOOn0TcK
LsCTIfo8fuszfnUqE7DqpdPiiBJKECcTo0CXijQ5v1EjGh46GKkGru3An/Dkfhtx
NmQxOG9mSMT0vq2skrQaP06T0IaQRrH/IpBWuCPbpwNOuYx6egj/+VbIzZQqtJcg
Yq7o8bhhjaXVlS5wPWU64XsIMFcgu3iyHetN6PW54ybxc2rOJlvm5ajMtGwz2O8i
xvaftBioL9SEXcgpcitQ4p/5pMKtSNj9+pP85hQBdSrC2yU9g1AkDEYp17Gb2+Np
7SaWER+DVNNxBaVOE6qKAW7W+3XC6DR5sxVQABu6kpaEi2diZgDK/cI7sr1t6kPJ
/DM0ml+3fj2jR12ww7w3mku643X/LevplEzaXuiBLXJonv72epZkeSYEXMJA8eIG
BUaTVo0mt/Xk3G8AiB22d2bsp2Zi5cmtQAAyK0TZ1pHSGFKxX30ER+CULjwyGGND
Rv07YTQqL9BHVP1wRLrnvtE9/OfEluP/bMF35e/18A+Jfl7O9Tq9W7wAu3ILbd+G
5UoTfxxrlS6StTtFRVo0kMm8olfG5Q6Csk1siEGKNY4kx0Eru1kLL3m9boFlQkXh
I95JTkzFiaWo87mPuAy+n6twA+kNT3fJ9kHXvxaNPYfXr4SXm1I2JlKsxOK04lJS
Z1KgTs9054Ug57938gLVayNcYf89VdEKbipPWYdtOfZgrjG75tFvHeYdsRcfXPcq
3I/HxnigjTxsDiCC6XNc7IacYX5BgwwtI9/M0yEYgQTVKUdmNfedwvUUAXNMcbxJ
9SeazB/bQwSEPHgKqyXKnJIHk/cVzyUOLEgxygqyJxrs3BJsMP+8jukuy1c5b0I2
I9NkIGTFUfrS+wAHJRUOBhqcktQbmwiHlRoapZLZTLsCqgxD3nb6/YmiU6Lj1Inl
JNUEGtNJXIdm4l4GS+aqiv5aaiWo/Z2WBH6CMluX0EdKMYmznXvgZRA3Gx2Jw+jG
eQ8JFpIRi5y8M9ke+pWSiM+ptwkTPKEDMlcvQVBhjRY9oinIdj/zu1ruPcd4UCkI
Ya3/tSUfkCKZtr3/4ccHjbYKKq4hpOy7yfayWnuqsxbv8KJAynLuWKxmdbNMIhG7
PlxqfEEXS7b2tf6bfADmlYyVRUTG5Eku2/4dOfPizaTxgkLSIVXhR25fyNV/LI/N
WTmZHRbhMG2GBzfeMTbfpe3o08uaR++EwWnpyCQ9NOv6Vpe2b9wgFi9Yygvs73YC
VUxLGJdBiRh+UEROJ9Tqe3Kr159aEHipWdiwE9dJaZWTXhhUrbbHz5/AAITxk143
+tORWzURF98ARAmjuh9qEx7ac5x+esJCAlW1TroJ5hhaG4WIIMLf2cu6AlrsLfOW
IytfaAOyykRC8SbkhYAcHZUpSQ5j0L0wCjiTkUIYsmzjgsKMyWd73IoS8YC9TeNe
38+dc85iU/o0T8Ct+9tk+i4+1DZDFinLW6NRY/PRJ0b1AmPg8QU66M7mwj19ZuJW
crBDEhq56XH5uHdrgdrNnwZUF2g1C8WuOYdzXHPMwZWQFAYqYJXsHqMzPIVGiPUS
zRu55AluIEsPDtQbAj6jHNKKbPtT1hkoLvAke9g4Jt+3q4TSKJMWfEZGL+M5d3b7
jBhtYkL7VX3GZOyrQb3oY/I8IX9qA0RF9a/ahQR17VFka2SeftHveLjHfBGq6Kjk
vARH0KyTsz32Jl0RGrUqLM68eCQlCiIHnsMW6ZxCHUMvNjI0R8C16/LWYPVdDQf6
KJuufRC0u9vTfuG0MXN3nBlXcoNljWbxt16wjIHFvxIpgXnmRXUsQ5QmuTjuGbp6
0xcfze9DbQCE62vX8jrc7+mxWOujHVpohkVYxSd3PrdsElsuz5RwTyPEarBeH/ZR
DuZnWfdolreW5t+f6dg3m8Wg7DyfFFoYNo0PuCktd1B/n1BF6bOopD/pc3k8Z/Nm
u5Tm+hKz0YhhVzu3xYhX/NNgxaflmGseYsQROl9X1OLx4F/NxG0Lk2NP7lwG3ccK
a1T/o1WlkTlj+ATSVOrSl7zQvgIqEvZ8gHUiCFLm3rLwZXQga9sFXbqdfMztwi+4
FG5cTeOBLvW8fjqbgNd/cGkhY45C0hIc9oMcEgx3ntcDjkAKKh6ZDkKXhqKt7Dwj
M8izoYBDj5jur8n2//Nm4fPPhX/AxGCGTOOg4eWnqF6k5aun7apHppT2ERJ0HFv+
dKqWBV7/DRWOp7jXxOD1xPZf/Ys/ykndGfNoY29Hg6UzS48qbZg6DKgfT8JANI1i
TXsYSfqChiuAtES9C/r8AnbkMadlsTvrvkS3Z292W/udQMxDwfobggUs3pXnJOyo
uvp9I8xFJN5dmJtFy4ns8sqb7BFY1ZCJmPUf2OsrAIBk5US7qd3KdMCXtWLTH9Aa
GzmNMaMD9E2MWqhXiRwhz2NSIGhJC/+J9XZBvNuV1NYk+OfgFTFKFUel3VjBm2az
vQDWz/g/jhpFsAPUNRZLjEdQ4GZIxluSRHiatzRS+oDaOIc90ktgmJO0Uj/l8Ji2
8n6y/D3YxNwjqFGGaM654sFvR/dEcmenJdXR5ptg/eolRZ0Aq+AJ9PjAChX+9Itn
SqZIdDHncI/vRrjm6FXPgExTftDE7JoinYtuPgkxytYdHQ+u52pVX8pQ5AzHkKJh
wU7ROnfKyfNqdnsaJIuWblQEwnK5tPJf5LolRzB4jygX8o8vvQBEopqybNy8MgKA
PqU9Lw3QzC4g/q1V2lJTcEd3k4H9h+rrPhRsCpQ1qH4fKBWlOiy/evBBBIK288HX
0VLE5ccJStXdNqElWdF5qDsJMeUUP8vpOyGdEBdIQ6W+MrEjuAPxMBFoxwghTpS1
/Go2xnsMUmu62UW0ncuF/04sL9jFMUu6A86wXtJzxVjqMFM7OGJj8otxbrv28T68
v6KzNkXGl1ZUezXF/zAFWIF6gHqdCJURt91QsDU608a/BRBPV+YwWwHtTr0E1Hzy
qiaD1sktQiP9vNRRUtV5qmB8YU9yW1qFF8RTYqC6m0UEScvCTfgKit30eAU78+41
UIRTjmXazV2V/SW/LwoZ1nTRxBghqn8gIURy2JjaiL0OiV51SbINdIxfEYJCvShR
L4Dd1efdxUIgl+RxqY87JEOmAxHICGlE6T1CwB6E+VRGdp5I1GN1T/HvLAJ83qhN
gRE+3gPxXo2btd0s1P0tQEaK6mtSa1sNp/WKnYbAMjmRBLW2ethWOzS+T/ssq2br
TVr0ME29uWK0yohWQGR6MQRHOR4qZh4zdKkx84CR5+5uPSQyH6b8xj26R7wDw+Ru
qatA2H8lQ5s+2BIbty7XFli14DnL8LIBeqtxGgWZ1/0R0RCgUgx4X0GS+iHcKz0M
9XsTqgtsrupb3dCiUzc3bTDaoEN+snSKjCfvMqHgRDsellgpz5fmKUUX8ijTmUze
Aaymgk4k8jmc4XE7lTvH//Dxeq1nbpZTbK31V+xRJFulRa15gYUEW7YM7LOcfnj0
A45yq55ve/4tlSxDp/M/qPQPaLhCh03xBTGX+H3sYgyXKWTAITkVR4RCSJK5Ktz8
+3tVAHM7M0oDnLboMcsaS1du8n0Xm64i1HIWBtvi80V9xKu315fmjpGHfPIZc16d
W1CIxRDNhDmdnfeU+GdgDZLPdhv7BpFZuUrACgjxqtTXXZ0arR69ZMLGtYBbzebA
PV65lG/cril9x7/LAcT7yws1IQRyBp1thY0KKqdzXt6d/RQzLT51GipybBLCj+rr
JUN4A/+7L7bR3+r8+uoiGZFgs6RkZLBZeaRsQgnqe7hiWo7sdtbKWY+gs+SWlEkv
+G7otlrXuAZ39yZ96L1PnIkjWh3yhYVtM29nHPpGc0ZOdRmKkPo8FAUZywm6WZ0N
ADvkRffNF2EZP/IB8YjmObGWW32SaifAUZUkS16SP8KXAbU47uEPBZPp48dCv+ng
iUTQ3iQqnWT7cT95AV+ANP/rq6O9/nS11cvXbglWPhTxEq/cBAXZecO0w4vFzy/+
cd0S75IlQuV38n53aqTstL/gLdZvriUfZvN0AW6qUwF1ghGkYQIP5bVGHVsps8An
xRKoYjqjIpl10zubCJgfAusjbSgsIFwe1jg7TxWLlQc9gDUoIIfCVT9iX59+Chkc
SHLGuZm2rSVmncla1DwXmArkQV3nUF5y33IfoAX00xK0KG+lA52eMqX4KH42ovqM
E6gexet0fFa65H4fP2dCqvSa08o/hnLzcgix2KZUQPTt9EMEl4Ucd3bojZfJkdNM
GAP2iywX/ycZEIQlXyKEhYoZJa4h0rWtD/2igXsVg32qNIIeNpRvh+/x4C8WtrNq
4PZy0H1xqkYpvZVlUmuXGm42XqWCc+8HcPd8aOZ5jW1+cEDyuG7/qH2xQq17xnba
5M8joZ6yLrdJo2KXeoT7xEv1xSG/eK5KBwcHZnO+K2eE0mMwpf8LKGT7lAdmFvB9
UIDFJe/bPoJikxheJd65PeKCcjUhrROwElbEotuUdS1/P8lTz9pxm5xcmo3TOQTQ
hw/E2z2On8XNTeAhnxwvHkTq8iwBJT7ehl6/1Lk8qDP1O3eF7tZyaOHFkK6SLX2M
tHvDeggbalMf6/iSycfyaTBf0TJom4AixwuAHPcZkFm9dJyrM6+Jdb/jLe07LFVg
8CwylG7OQxsLbBm/GD66joPHNh0GOlP2N6D9dndBKhGysZaaekxCbv/MPOGCKCOG
ObwYN1XtsAlSGYuN/K5+5cA/zj1lzqgM9XG/RWu9fa/rUb+THoAC6r+hnCIZLiZp
66UkvLaapMGiQJ/2n7oNc3mfJFg2p7X0FE6TcOP6IZ76STR/itAKcDRpy3jr8NMV
RbdH2Oxk+qAj17hD9yNXIWCMLUGaSUt6SVrlysHkCvX5voiLi3NfgXoL/m3LcNNV
xSTiTK5Z0o9MOL2acPIrFMN/MhEXEAlca67DKxPs7DBlFSbDd1pUHMVW8VZ0IIce
m2WF3k3S0UR2JYdK3vNd0eRjV8k2hAeO+PdVoLIp54WwzomQHFlKnu0pVI2x4pCr
j5VSLXhajnxmU/v4jRoBbkVsTe/NwkMkIG6ECKjw+bw5rkn7D/ZVPI1QGLNL1mRZ
4uwvoSTMq0T4dc3feWcbYX40yv/wERjgyU49Kxl5+pHpwVG3PZ8TMMOl17lAFTB9
L6/cEQtYC9HV8JpqWZIrKqnP/jFz4rvAOjhUkfWRnDSBTIc2mUrb6tH1AznyZ8bB
9GtK70N6pnoFY+WpWaDKGTqsaBQBeOTXoabEVkGtZxdWrqUSGwxETuB3Wr+ou6vw
H5J43yLH4ox8xeZdM/fl74Z7gU57AhTNTFYlNIIbxBQvkeZ15fbSrRQe1H67Wzro
/Y+/6daA+DZSa80iD2XrpETHJtptp+EI/P/ZWPI8XXStYIOfyWV7T6Mxlsg5oINH
14A20CcDeOBcrNu2Rh/lRFvBz4R7mIz+pghP/0gx85QsO/8WllbrP1ZwIEzXovHe
jtsNJakavhNswsjYEanAS2X6B5QkhCF3Oysf4mw0mlTQwALTl3uegKK+tZ/pH39/
Kbpv8XXy+x48CaIZDUWu34KewB6sUKHJyW29fL0RdNe/b4Gg9p6zqNLyASI/ZD3S
caA4QHZX2Sw4NndWIdkoRBi7aANb8i/Ez2fNRZJXtUIwgcEQ83S9th5iGEvOrkxA
80uzFVmfBsilZjda6twy97i/6l3ku+5JbZiGQ4UKDhWXldAKxnGIA4R+/F067+g1
m2afJ1CPyObCThXiXQUxS5880HMtVVHEHNCKMJN7cpa8g1KWjYqbbUDO0t0Q+jz8
19M7IXb0eJaKMkMtq7fNHHDEJWdiNTB0I9Vzg7MTYNeMJqNZBtYdWTJ8maRXDMiU
BG/NrrPXXgAMPcx3jKCqcnUKtkiIVk+HjaGije4uM27g5MKaRXyclGA0SzwgR+73
5fezDp2w375HISjd6lV8BPMr9KXuK/3ylXicbTmcgxONqlSbHC0Ok3WxZGhnV/Ev
IODj0ZkaNzL2yQRyLyJXVoBWRc36F1KUoI3+mJ1EUkv2lhlTihMCjwqTVDkEWzcH
paBrnPTzrkn71M1uG4Cb33ZR8cZ1Pc+ZqipGQzIBVKJR51UqgIEbcVlL5Sqtwgw2
8ueP3HBTgm9arEPx25dLv2RliSX7xI1EMgYZU39HiGidR97i67K2O0Y1N2MOrgeO
3jfDHt+6rW9a+TwAxiXlS2Hqo5l3E8v71FjRqt4Rwo1UqBadTKnbBD1RodfC3CTM
Eld3FdkNtEc0GlsiItXhHiB0M47UpCroUHYNUFHzEohA68cZHZbZaiIQQrdkb4JL
cZWpvGTNR+j/AAdutA/NuNJQjtvmo1tKPt1EDQSxydSYNwSifpB/+6MuV4S1TRrv
ppxZSrrP1u+pfsZiWZPItHxzUKY8cgVLWAigvcLkE/nqd5qPn/lk3LGGVCPKPwoh
b8cQXWU5J/ulE8KEPQT57l0ZJoJ6KMdopq6+Bb3k8UuLeNZ9bWvQ7D94et3DGwSA
iWnQdqNjt7epo+pBE/F+8l6Xjx5wBlfMo5xlmF2KOmrAHpAjY28m96jWyQJtY+nA
rcfXGfeiBr1Y9oE4cFc99QOlqLO4Nfh5kwzFIoO+68fAzaKnkvGQA6lDxWKf/1Hw
BSPwNT2ZtV92iQQlI+qfWjLWmUVmuzSGDiCy7E+ILDJwj2HNIqq3Nlj5+ZntvmKu
1F/rSXXB3gsqEC2WFdyPWQj9hRY5eGqatvpADEWGGCV5gvKe5caMiaiftefze0So
+uxlbJYfQ5rjO054R/bs13S25Z0b7J+7voEPNYwTm5GHSBtchD94q/CPOReMKrsQ
92ZJhycj261aydlRPtHgCEwaOwh2SS1NUNLnZSRAESk1yVDYwy/RNuYYjlGrIj2N
qM/TxXkL4Mckr+WMObmXy20rr43YO5XmsMFBIixKTVnhCN+BXYMIpKi2CaJB0C41
Z74OWfgeicKlSaIR5Ovn5nqLV1Ry+vdu/vnczb2YkJZ6bI7KbHJQpDhtM+o1HcSa
RnA3k3nrW2EbyFcYlX0udAxG+Obx8C8fPyUZ4q3pbFTxHLfX83Fnat4fZNJg4jJD
7Fj3smWFBvZbI910DyEhGV9F20b6247tnW2z0hvKwfAmZQLvVehI1IdjhW+60hPc
UrJ1/b6yAgHapEPfTURnBu7bEMQSL03BOgKaOb4yYsBcrdFsa9bXvXvDtmGSfb9F
xm9Cv7SM1DlOkqe1PtZpzNAJIWX6GatxiAJ/qxMq7MPKGEdx389tF3ts8aJj+pVC
c09/qCTvZRyhB26xkRNEGabtYxfoqWxjUKWZgjYKGiE3PeMYEms+nFE2pDr/FqD4
b4oSQPipS5xkWQgYTZC570BA9TQTteTMue5LFAVwZOEnBIy9WDkA266ylBJBX/Wj
cYq7n2+G92uMtFMXqAeQ1/Z8nwbqEyInn5HXMQkz8d73Iz9W4n0kjtJsPXHiMb7E
y5VDGmpGp2TX17cGomCjCyKOAyg/xPTRqzJvWm1mWLcW1htp7GX3S/OwpcD3pPCu
o6oWb0puVcSM0XQ835uBY0NBvUaD7ZLiYUAjDXVUw2HhivHh7IohTMtDCDlgg4BP
lYuRh0b1tb1uxu0hjDXWueJoRbKzXkMsszPY6sMl+dq8IUUuFuGU4yRKl0/MZTaP
AZ4yus5geMiVU7IVaYIm/bFvYg1W6D+G/DoLplniS4+l6n8/xDVJSMrBQ0IvMYF/
2szgB5wYKSk/jmqgrZ4WvFOq5Gj3nzyV/T22u/JhHyjRLJ/ui7nREvWQ8LHhOBhI
mivNjj9uLQKAfceO6aYdY9ZXu/KsoBxf49t4lO80McNuVcCEnOcqjg4gUWu6m8Qq
CW5JrrYPWdFXN1wTpJ+EMSL+PsNsbvu2/w3aOqIk1e/slUMcSpbodpkWhyegyzfP
44VZZsEGQu8ZT8WNn0ITFi2g7eDStkR3ECo1ZwCjkB8XNecbbxEZFohvhA7xUVOK
jtLrFEKxpdqLYjRDSRTG2UX1yHjow45sfDpqgp/M2ps9Sy0To6zSho2AiBbiyQ00
3RglXLmGn7SioGLeC7T0lICJD3YpKby/+nBOc0Q8D1nc6O/Q19N+bsltySJIKugJ
dfb8wt0aKrBF8JXkskhi1tSdMW06ndhgOndp228ldTRToDyUJJDuf+JRue0DfR0a
RUqsHGMZvuejVXwejzlcd+ciD6s/UGyzBQxnMtELH1R0KzSiVVba1yV520l2UWQS
66RJcg9hDmFr1xezx9whSigIaSs3fvBSeI+cfJtl6tD1Z+FzStL+AmAjCwGtHVsk
xyveKBWOZ/bT2O53AZmr6LSHugOAB+l5r3e7gvtEUMiXW9hfPNe7/kxdS2cPRUWy
NQyjHpZNDw1SJRvumvk4PzkcQOCh8gPHpK8KVYJ80ItTF7ezoYpM5Q6YvMwca7wj
UoHggFz679WhUHPedsi/kJhHPKwDerefPzbQL7QZlxkZB1SSGoGqKgDDCztbAKMX
HpgDNNmNRpmNo04rEdHO+hnl+lVNa0tWInohGnI4ah2FsVnaPQVa7T2maNsxkSzb
NK0CaZcvyBSpO7YPB1EP+pvy67MPKobE56g4unZYIWV5SDva7Os70ti2+EWywGzc
u7ngqGBK6tl94HpX4BD8dSHwafPoO/mK5mFVSR8RYks5OT9sZ2Ca0XSTQcbKLEdA
71FRnJvIlDdgCr+Y1v4PsxxLxGZWAJfwhfhWIMHdJ1vwcQS4tvwncwcdQzk9VZuq
V/OqT//d4gDD/PT9dC/cN8Ewrs9RjFMEOl4SrbPoxJ1isDmobG5ZmxSioIMRhUgC
0wpo43sJopPgbpVCFGm4OJpwlHnSh9T8HCrJDk0KM9RiqoEUYamhSGPCg/dQRbZp
mHQvP+sHMiOOLfJSlbT6CEhY9k/ddG7+AaizjRQ2OW/aSe2Bc/mjPfsfc7jwEBBu
igqTMNjB9INo9GXo98eaPhEzFAVquBvXwa5nQxAD/tVJ+W08Yg5lsP2PpJsiuwyI
ws3zijIU1jCau0sVHwOgwCEflvup+TvN6zkwlyo82+zSwz70eIai+XSvSUAlq2AQ
iNEppoWRSBgEIdMz5F+RnMBpmycwp9pKkBEcKWE4WDE3Mn7M9g0Kv+ehy9V9AcJ6
72oJdwSwjcFvcOIR9OhkD38GW0SNLanO768Wp6UPUjDt5NRkSPLbIT6TG0LBERtY
qQo+a87Lf1Fso2qrFobnBjzflNrclsuwbXkLC3aAWHDbcpzblaZdmN0a9SvQ3bXA
IJoXAdZzQsHc8o1+2AOALT8nwuWjB1VLBWuPLrNjnh61vwhhcw4jhbzSP8CJxdOT
fSy/uzOjA0Z92yebKrxxAeJh0Pv9zTCkErOZNoK2kzr0Lks9yQJGUuVpiEhe/2Uo
Px55omEvgBS9r6efKaAe5VNZznMmXKCh2j4NFSXQzxFVHK98F7x3nu2VdWL6a2Sw
mVsKz8aEq2vX4qZ0dhzUb8u5l8Bns7spDIG/ZmSHw7F7JCzF1C87VmnXLLGW+zBI
ifx/HICQGjkFEDJj6NNmf0ZkJJJvoJl4GVLOvFcjI8QKVTDwU8MgES4O7HBrImFp
hH8eLq5BFbFTBOgVD+gikc3cwBEcuP27UVyC5tlEeLq8zzVi3TD8O7NBv7wUh2q8
T/yqqqelHMAVqA2/ax6heOKuia6m7kr6z5HspB0AaEVys+8fNSzkY5qfiKacXHAX
2x25mVYxMm2c+AD4CLNMdAvvgpa5JgIV7BKNbawGfeqUfOJc4iNA8WrgBXRgV37t
L5b1HybVxKB/4mppcT6WNd9BW2Q5WJUEbWvMh87cFObn5js/bgZb5FQpIiE+LV1Z
cGt0HdFRcB8aLkU1c/GwlvA4+2iL77778VDNHL6cOlX/ZtLV6dPHfJMgQg9zGNxv
/p68HIFOz0dgC4D5bgVu7IoqJ19pMx50cJGLJLVWR4lEtoGmY+d5VcQpUCwj+JWQ
84U2WRqXwzPYGiMNYrZBqS1NDFpsn0uTv2vUysr/BKpAPS0VHNqKRFe7tY1aFW2H
MaHqZCdT9RyZDmOV/jdM8AUv7po/PqwBvRRRAG0CpVM06GEEzYp04JVUjNdlsAw4
tpZCW35zugGjLPxaw9t8i03TGclj4YTuBdsHZExWajgldmUvby2xjrw5QXbnbSD6
Ca2eWJpSnLxqJ4k6DCNPpoGbhKAj5qBDnZcIF48yuS3uVulPSIbUeqw21G5eIN2c
IyqlUypjKFuHGk0cz5MxCh6n84wtgqPXgZINKI70syGjwcmduv7OUrtnLMmvtB3X
gt7Dn1B9BzxtPMqbMI+QBtDBeoLjVSN/ESb5byQX0Hka5pCUJ0KRVQUYvihS9AxF
mp/S8S7Nj3++RI5Ory+505wId0Hg63NVI+BI/DN4aiYBTv8GyCEa0V8s4u2na7q7
s3YeUntvF9XaNHTERr0UAzAvDl2bFhJE6P/tEhE9v34pUYRaUGGmJ5BCsPUeZsDP
cxszuknZXTIbWUVeDSbnKNSaM1TOTV0bIAozdS0wbJxmtrhvriRN6CxkhE8kD1wK
YFCLdjzAmCLRY3BWa3rv0SrnxcRaRINgt/UkKHM+shr9F2k25aIUBbDl1wjELiZR
QaH/bLn/KMDZYXUZ7b3g3tmxS18D3TffGACkitID6QIXAsEu13/MuE9otHT678YL
tV2f0CfFvdFumaBelJtXu7Aicd60Ue07oJwEfNqsDAM88KWv2Dr0L/8rOT3RMLbp
RbFZRrjOHq7gRKI8VAPo47wxhiQbaXS3anSwxhL+Cmgmu/jqqV9wpPvspxfOBZNZ
rS6o4hEJxT6t1AG6DlutiP67R6YQ4kD21sL/nDkoLvD9C3NFwGO/yezHnD2kG82J
ofFlwAHgsXCaFy7auxDKpgP+/4a4PGBDKJVbmraA1dWXXtWh6T45oy271t3p30ft
QBkZfDPyfpHAROi25QrwIOnW7do3YE1UhP7mRNax3sx+Ptarr5lLhYrUHiIAI/Rt
2qnP8sIda2K+YieWID9QZpNMkZg1uckxpU9PaTUoFWmAkG6TQM1qqMUJdWxu52eI
Q+odjzwR38YWOt0/PMd6uw/VPY6jngWiNUpNKcwsvhc4DRSGYAQG286z8fZuO6+d
dfzK0hZYadgjknOMuTz1/gBpSXV3+9PH8HglOdX5sArVqtzjKkLxnFu38YpNAFYc
S1MByvEou4no8UsOUZ4kXBjG2sTvMGwHu0R1caPbHJeUcgteVCXydirq6NfQT7f3
n7Y3eV5t2iioru6cl3+2cZfYTmENBimXbIc5mtH9TcIXbQe2qf7BqnClpqYigD5m
KOEq6cNe0w7MMXMOQ/QpuAAeoPOEknoEjDWOaDtwfBx1ryTNbewoYECWzHTX2Pd3
l4muknW1de6VHaB49K8O7V3qi+q6bDnPAqUXW77P7jRqkPx/ENI7+QXV7ToXU9st
x6xnF5BQTvL3AvCD+QOtF+NtN20QYAYlRHqEI0OoSJMv6FJ+/JHUYX5E9VC1YFDe
15xLTN82vMOSZ4sxI62aiJBgzl33bXdCDaHJrNnrL9xe3IBXol2oW8Yns3bFGqcN
wRX2CtM3avfHcyAsr7oIZHJzp+rrWrWqrLiU1kVqVH5Y4yeljC5uz8Eq/E0SKt8d
/0aOM5B2JMmFqAi3HGo3Bidp5ABvSO77jxQSu19C0CnRzJvdaRfOVZMTcug1vNfI
RkfRe3QsnRBwfhbcQZSop6nchQTCs5YGi0A7dlGmPrxyw1LQpEtYlq672qYomnz7
g+Oi1CXMMOdoWHt5NgKGUr6J3qEyaN1CR3HrDrVTKwFg2yjiqtdUBF1GP5EdWLV2
NVar7zPETklAbFL4ZXNWmncSoF0jRtVUfMk7itjXepnNpi5isHEQL1AqRdFJrPRf
RQXWVjFQkZER0OYCdQvnI4cthDfkM/+hODDuJPvRmjn5G37ORpWBoONmh5R7V9Li
YZFClzQl/FuLsJNf7gxg8viiXMRUOJ1IyAqUG6w8vmz4+zxba8MkVtWQSCDJbNHJ
Njw6/2Fdn/W2DhrLCjsfzD8PVAH30SqEccwy3NWseAAV7wYvQS60BJbdOSEbNPHw
6iKXVHFKc+hh6XKR5sBLWlEbHAaN8x8Zq3LvzKdv4pVDyPXj0NaH6aDJqW4YXRGc
aSSoQOcobXYBomHsyUR7/E38gbDKQ8RicQ8anAZamT562pG0cq3MwGGQY3pYuxqM
1wLxJCTDlg7/VhM3y+eujLLBC4utdAhc0R9avdG7l0e5ezqY+C4BsLTv1NFbJtBo
tQIZj3/HnMItfiq3aGTi9iShjBj8FGw0RAIMif8eGIpGeoZs2le/yu++NJAiqa/w
lIg1v/obgRvG2lzivNCjVvBy3BKzn5/IXxQiJYML9YfmksFerdcTybWzfCw0zmeE
t22Ko+Y0ZHy5mxhgqDwOiO9+RLIGNRTvoEqQioKiU+SyxmeimMXtpEQUwa1GnGG2
USgfxaCro+KC57L2uajwJ1zRDlAe3rAla377FrDsivejBb0qooUU8jgoS7djq2JT
62UE9mz7PWS1D+kNL6+S0PvV3B1qQv2s+oYH3vmtPUcPKSFRaWELgX2vUEcNFZ0r
f5fLMAct78CHIC0tFS0j//TR1Jmoxnjv3MN3vjC1Fs4N0hTcnXnbSeTkmaYim21Y
cLhyfYUte/AXvDzQgiolTtwc00mBY9oA+VdGU0vfGxkhMDtyff+epjsc1rNJhMyP
thd8/gxBvSd/KYdtFIPrqOzUt7BAxqXBgyOq/cKsuFU2ORCS9X2L4AUHWZSFgEwl
gdk56xuTCwK8EBv37Sh3cnwVCcAWUUSDQkNuraiQ/N/UDEYPnt+1O2Ng9ORPU/oK
xEBUDIO+h3pgLBntgekS3Rl2Y7PLqEPTzkwWDMjanS0RMKdYHF4nf5dBboj5dsOu
rp5CsaEbdmVaAriIHpl2vpC7LHCZItmGopyrFCkM4hvsxtvMhYc496cpx2rYmnKG
z01lwQlE+V8VZvyjnVHocxJjvhpNHLdCZBLC/7Ags23Qr9pTYwqrhKlsyIHV8eOh
XUlkWI+d+qearNwWqSP7RwbJHZPZD+sKftBrAMifxo/CNnhMYGDwTQFsbeADi9Ro
BiIYKUL8xQmrNgGKq5cDnE3aUTKKBXTRHiCzwZ7E1s/5Knlx9n5Zbu+vSPQgMc/q
JRBEBmyUJZJZdUSdIZ+ry3PvnxG61Jw2MEeO/voO5VvC3h2zjOf0uyfYbcdrryE4
NgZ0BDvLVL70gDkY08YjnOvnyznAm+gXq4W+/i9NR/QLf7Cog30OwTkjvK/R7lXZ
CDPE4XDNnrldQO6Z58nMfburKb+r9HmCPw5D8d2/0vnMBDEL6IMXXT++PGJVY2DK
fIqs60079yMJzQKLqxokDYE1yDXlbg1PMYUPzeEl4R3NzDYKDNDjh1antoG9M8Vw
XeU2uInE8l+LDKwygH34aTLeKF41n1UXTiUfP344guA97xDW+fb71HTRb40qov/e
feKnQXCxZv0L7dfG3aQZ100T3IIw0LpaQu9rwT3/JrQUEJ/5VmjQbRcRY5uahCTx
3HQpNIToLomty51+6Srp79VZk14Bit0xXEaUb0tQfHqDfsRHMD4RiG2r43PasmI8
Uw/yGnNDlVFEpkU6+XRm+oFRo9LU+nNRNyEXPx3XCZI48uRB4x+syHLx3BZ0oMzG
2qzeHhMAIr/850z1IabETlsmEf8RexjGJ62aOQhPkNIcxGWz4JTi8c8JDJBX6w01
iPYBqtnXmCdktdSlvxvc5gIC6BCq/ArkfWIYkOdDBriPqlLknguN18KDEY/5HLCv
RXBXwyFCq+Mj9wvGfIYIDxuTFpoMpDyztpEa3Ei36urxqe+wPbyJCsmHWrkrmHj1
mvczQB0y8sdvQbY33AjzhNgDRxS4fQcE28SQ6VEtLTPcP7TTq1z//nw/BYDJlEmv
dDOKce4oQ0NnlSw31xeaCD/9zwV2zC//R9ZNclKVuybL5V5Qg+gSsgQS6ClK96xC
+7stzftc0A+Q3Arkwgwol6qza3tJ57+DsC1RpAZFh5wb7eITr+WSwaDTNL9PuP0t
wFx4CUWtQaPRgzkMJj3MOkTvOnLD8+SHyqRtOaRUYVM4cQRjfklsJKFeJZrj1Kun
9j6LS8JbrRsHWH000LWtlkOLbEGuwhPMlT0NEOEAAUMrht7qk921BqkL6+47zEGg
4pMmzhxjP0krFGZ5H6R5xSNST/KWNJOC8S6Wuc289EDnhjm0PjcqO02A55Mdidgb
b+vQtqQCW8f4v9VdTWbAASXN3g7YmeA0X7U7afTK8FTXeeXyOG1hDUFaGsRDMM81
GeLlB966NA8ZvRpLH0tMRqdazT0gkn666qWke2/zyod8SZEGdQcrHXJmuX5ocu8T
45tF3O0lx8BY19Ka1hnHGINLPM7pOS1uBh4Eod3/QiMgcUFvGt/79jLHeumF0pVl
DHenTQFURn5dweIi3SVw5IoZifPZZh9sg5zGuSFTNtXdE43Vk3u1eBBvXZAHAqev
I6Bri95VIrxfdKUdrcy5MscUk/kC9NwBqP9x9E52dEctpnKa89FGw1JBah61GUVN
JouX7K5OfD9bw7Z3Tbev9D0zcVtOgpf/5Gxx4OEMlkpG1ReqINI/84NPAXAKzv0G
VKRk0V43UYE7aKTgPiyP31vcNz2M/mGkpiFvEpmvAv1V8MINwdkkYx2uIw50Cs4u
+ktvPwS3jW2ta3hse95JfwNHXA5CoA48drTSC8TfeZ/A+Fsbm+ISRyNHkykxw0Lz
C1HrUbxhowiFrqbt1xHLPVgm+AcJMOv2mGyu4QiPTYweCckEea+6Udl7TYmBNFV2
7r0J6qtPQgP5aDWOtVXSvLyaJ65fXlJ7NYCiH8UIf0gUYScddWaozhGW9/LavQ0u
lyfsNVLY4cZgdHyLyKGlJwZZ5cavqlwO/VtVqAIG/tvL0P2L5uBimtjlEy8L02I/
tykRhCSyUCDbCx4tcsmrBg05xe+a1+F78HFxb75aZhbAWgALxFuINhdmN0SiiHcV
HJtbnvZyOHzUYK5mqV4NKcxmO6iSNcYemkwNj0XJTzjU+TM0OTwgupwyr3MF/8jD
/rNQMf9k7/6tNPuK3kKEEFX0SbM9HaLCsCdHxQ/qpALI7/M7k2MSSo2yJmiLMsra
dk7kAfe7Cb+dw+b6toqUu9lug+RmbC7eFd2+TtzGxrL5l+dGxwNcL4DRiE7TxF5P
kDkjUVKZ2uG6CR5yiFytHhlMTxXLCVr8Isu/wWt7zi2upNJ1w2lib0rz7J+QOXY2
wmt+qLbsIlsLzjb2pyap1etvwSPs2u2FVvl7t2FJzjou8U29PaRI3oAfoZRSHnXe
YxRC9tXMzQd3z3pI+KQrq7cP1/QsGByieCjWgYHh4Cj6/Q5EgIsRVKmGMYl3Dori
Yd1M+wyoHZ4roiL6N8YL+WOZtH4ounepMNGoqHWbEKJRp8+lVE7aJFORHaJMMukM
LOLs3yw9FIvzKPyhvS6TpipMDwgqRrUDAE1Cs/ryZDUOwhOetftbrIfZVjru4zXj
JZR8nx8g2IXvWU0vDuKupkvxHvPezyYhdTrYNIEAiXNzMyoQCcObCFmtU+M40/Uv
8xnevPfaHD7muK0pZudnZeDPWn0lrwMd6dcY53ixRM+ACV7H7HqYFlqLjLeuCwwt
MQmmEETuNq6Etv+Av6Tyl6+QpEhSQZS4Bglwnjp/ZWkNCjcE+8d+KFdYYK522ZKo
LOvWfDySzOiAlEGd23sVAUZ4U9Ig+wfClkpLkmifwtHdbZO5X8vMEjo643QuBn19
iMlyQbuoUWv37cDiSVOtKBxqvh/EaDlqMaZcNLKZhqh7CW4eH4qeAmWvir/yRW4c
aYJ8gmX5YmS4bqmceogDZZtIEJmgCHzvOq4k9Lk/2OUis4e90JoebEUbSOEWRc4A
EalyYUcImwzepG/Ra6cVhNRKXzf7vqznIkURMCll2nUp6I5ch/6v3sa7QYn9RHWL
wEs6+WvzcOMXXZAdnKprCc178OLPmwu/FcG/vWa/nn6sPxxLPccJ2oo7/IQxjKxD
SOt7aEp+vrpABs2vv37Ip7ZHDLQLevC5Uh66zsUeyoYc0piqHRd7ui5q29/7fjCT
uYM6WcFYdUvSEZ2w0HMPd7uFUgAnAVJa1aU74Q9AnojcmsQs9DLAsdZmYCf3jb/S
zhg7YAxFptPuO35Fnfm5NOw79x9q7tvWchyQzBKXNQxkTYwTSCDIiv9QxMrf8nqo
s3359f9Z/pKNjT1DFQnCPZAmy9HOmdeg54y01l8z4dQ262m8Yv2/xkv6ArhtH/Xx
21gXoCQrsC0XAspOzAd08TFAwAUhgALjeOiUXmf2M211TZ+xrCXGSpx1X6YhHxDJ
m/QWxzba5WMSjdJRqfXxhnPjLEVtwSjWpOxBUrCTX90krbN+BAI6eYutk7zZcTql
PghQ7XvjjKrW4gIP3XT4vXBHTusP4/A/L3RhKsAy2iwEO3h6gge4MvLKRMyqjS8o
4HZ7J8digLFBbGa67/HX+ZOHLJJ7G9Y0QmYqaKs4CinRQyjMxhmW4v8gALiXhpm0
y03P/t3HsBc/pv39FCFkyDRcUYITUvz2C5iPKguuoHHJo7W9nZOu+PQMYm07yaK+
hjLuTZlGF2pbhFfBrpdgSKNpxMn5OBz+qwDIU7V4da++I2ngKGrQcCcC0fe+Sryf
iSgcK6rFeHJdRyWoWqdL5VAj8F79k1a0H9cjGMVZGXsHAS8NgSCr04TRjB0PGuB0
RWmc+nW4vDH7ialbXcobUQfWlhxa+HCDAgdjI3CWeKyYZ+3t4NJVPTqsezG1Ucy/
Q0rTrsmJyvfDFkHKp1yGOQQYWtRZr60m5sGpqtUrb/kKkyj4Fb3QbUdNjiBc6zXr
TRNJSaNRFEAzBi/KFF6u0kahzewsneR1be2B7SGlkDbAYcoUTxbDh7wD+ftaIp+A
+mtm/mvBi5T2eRBDtlxd3yPhJiMDoQy1Q3E97/F3TP8rqp/K2DF21wX3D69ck/gR
zdBN7EfxWvtJOARA39wMU8rmdcMGMNlrm5YNeVF3Rj7hXwZgd+mi8Hs/QisE6fYp
UFjcNc/cJMu0+UxxFB7hXAaGyg+aMImLszv6uERbpvE98oAPLNirIbiPKPj4hI1N
kXNpj8ZNb8pGmgUTlmGQCl06w8kPwKLabR4et6Ee75A3cMdcENdCH+SRujQPvPBi
EWRiGExqXgei6ukzMyrBG4mOnZQQFcBwJzDbbNMJqIXOm+IIqZ0hOKcHT6HzXgO8
SlCRqCs/4JTOCk7qVA2pBBqpRYHYwq87x99KHqPJZRdvTjNDOw/03DYMWLpCroc/
cnUVkAKJRSRKXa96BYsr3+CznF0JAIVlgyseD+DW4SgqpfjVkE8gZsorNqHEyTkY
+yZ61J7BV3hW7lnNs5J7ObUGHnCukRX5E9b+M1HN31ppSSQXx4IX6NqUP4jKvCst
nmQ5eGXsrbDs3kUg7QqU9HR0D5lgRXosxWGHNWExH/xgd2p17m19qrCtOwLABFDN
kWLUATi6wzXDToZMaJGVNMEfLTZ8Uc6sNbAOVs7G60k9ifwT/4LYLJxj/gAnf/T9
IkmG+M/QuaossNNoY/KUq8/YdFhgpfqoGQovtOYCQBpMwJJEwSVRZm5dsvXqE3XA
wtTFmbPVUwOWTfqu3BcHXbOf9FVWtgofowOMylgUkWf4ei9DinDjmcFD4LBRzM0i
9nXb8TnEU32mM5x5i0xtQfuaXWmvwrKM0PMRiCRZvH7rJDodNQ0BmtkZQCdmPIUw
QjN4sqAaG1/eyBb9CvIYn0SBlV2aHBBaLewYTgvxMFkh6v03WHTJCMUjbfWXLLbZ
hLgrCqo7bDkx9ZgE0SX/jzuV8D/eg7XYqMI+fERZNoywf9DIfTlaR/d9qxOSGUzY
Yos5UznqX2f9rrNWC1aqThg1XGOepwDoxousWpP8hGUdXQQS2mz5yC+5PGUZbAYf
Ps6s1m78JqZvFFIqflcOUdDNAGVkueixAZq6nUUBZFheANBxD6mCYTjG8oINe1G7
o2YZXNYmGgyTU2+xdREnnb0RIbf6PLkFEC+0iDfezJq4AtEZ6G8VobZWXoXqLPps
glTNrSHvc025pNomyj0CklQ8uW8ecnOIIyzYLFOF5i5w7LlwH7/HaOhhnfKNNF1D
O1JHRyXzgohSqXeQa19LrY7quWZaKTbVS6m2QPztillpYhze0TWAh3gzqD4P3VG5
E5ZITQ3gKadag1ZGwxiDhP5mooprGJQLAcvXLGkXO9WV8HbVsYxRssfwKY1cy0XU
H2JkNJFR6cX9fH6d4ZR64JCX/NaXNBszkOc+NfTDTiN31RWnapZww6QmO9bTXjDK
NX1Ib5ZtKgZ3JOj/Gf6fZyKnBjHMMxILqOOJjOqVpSHzNEs2yuwXwHZj/tuQ2dkP
AZOM0gZe2DY1u+F31JZyixFBL6OpYMM33ohQzuUi5jug4bmrDBY7MdDjkrpRJPSN
MjqtwqRMGqFz+cGadjQCcfvGL0A3EPtkc+Y88vuGSPH+Qb3kjVejMvizQZ+GWAnp
qoYr1rC2/k5niBT4YqWx4m0MuVjsS8H5bGd8eJ3sB6kHnnux0pZE4Fvad+DGHbv4
4T17rhAYd2v1+wNnGdr6HbSW6Sd2DEiw8qbZv6dME4uxXa/iUhNX8hb52qkVVX0P
fD8/pK0sMiz9Rdg6ahKxUZmtINcF451jryJNEzAMF76RE5tE6ZiB8/VVhAC28wyy
2kS95raXqAiZCpakFg4i9yfBc/HR9ZXThHxxCXDVS4L9HCaZ3Uz4zBlbm5IEPdC0
UcqGQJg6/taKWgBv/uunfC63iWSj+T9IUztXEykcKOhXzHzd8zsb7IQPBMxuKDTK
0D3qdGDC+4cZfkd/BcBUmJY5c50xEEliEImM1uolj2nqRmfN3TDfTuWa72UhX7tS
q82yD90SzOgV9LsU4U5KfaL7elSbK6pWP5+pM9X7Yf2GEfBswFVoWipQ1p91vGOn
5l4TVdT+ZzVYNEQH57kmATE/rBpfQYWDFCDig75DLf6ukHsXNZoeYFx47MCdItPn
TtwaANbYxgJICBQmQRFVDwIN3pE8iARVTmG627+rEeQT5fOL+2M6heH6KiYbCUF4
pIykF598uxclRLvDXYvpuFQ76H4LGh/O1lO8B8TU9SwxPgLTy711Wpl1/dHfEw6E
j7zkskSAunx6i9pUbgpgvRj+inH3T253nwB2dNcW6jj7YG/relOuxBFLmFfOYfTC
UN89jT/SuvMaXHCzq+zw0flT07B83psMkLQxR00Ea3LYfG7APgOSdXLcRIyk7gEN
BuCihUsS3H142gm8dBkQPDpSaX5tFcRDWgXr5WVd7BKwcfHW5T7T7QoSxZvu7aG2
k0Ua1mqWho8QojZC0tBN0nOrPq6Kh3aztemSS97oa5PewgvZ8W52ADEwHxLK05J3
FOYEA7GVsKR2DE+rSoXGjY8fPgW+xBrj7m8gGIPLKHFMj3s+7Ub9nhF3XTL5p3ib
T+p6YXekLFZokAMUbnp/UPmhug2OtTFt7ey86AO5/7gmkCREQXHIvCDM6C0zJJBp
5SZy3eHe9STA3He9eCedlYM7x6/KZrXZCd1Asi7+ATJWh5BPFGM6mr7T3pPBSFkX
ct+m2b8H09vHReTFAWrNw1U6T7u6PkIpJn4Z/pH/CsBhlS3oH7k7CerZDYaDojg8
38U/ifvDPDMOh6ifbTlt+cROjgK5ApN3fsYkf8xP3EbviIditgq2cewoRHiFY8bZ
D3UzM6onqKTZZo5/XCcB6hibvHEEFbxXi82qR7xseGZyH8bkTsL8Ps8VBkiZDyQl
RoqgiT4X3aG8tnzbnoVaNh9aMZeQvpxnCruScHKbmEluQ9YzmqgGQa/pBk9rBFt5
MEUwSszm7kepz70iw/ZMr5Z3ylYqCHKhvdisKfJWJ5xvUi/b+N+FSE0hekO/ea05
gXotp7eHsOJ42Dz/cDWJj2wDQLSR3je9IekqhLujeScSrCSZglEhCCZLtx/HY9WI
U5b0CkjFfG1Dg57gOvaAQtj81HBtJUkt3NwFPrLynj7VTv+MKSKZN1jV1yaMxPR9
CZQE38c6RT2xfWlrJOCJGDa8a6Htr0scmh/DMUAwt6/3SFlO7tAcSYSN+AeDMF9e
wAhgVuvHo94gFYOnhHwqpwy0GtF/00bxkoNicYr4sIvqcGLCo7gA8qGfnPYUnXe8
8cs9xwVlmDXQkhuHRY4pcbWCMhdkg6simzhIsxB8pIbHa+wwRFe9zWffpBQdB0Lx
9mGrG6IRn3hymB0Kjqt3CwfHvCX/u5YIrkP/dznTlcUSh1hDC2WyDQH6lXd8suZy
JisBQWWnRK1zQWOUfJOmDFJzp1W5fpkByCnMVxWR2YNlil1gd5c2v85zlDRFx7rV
P3b/VHDdsdr45uBQhWfCa2j8RDeUo7OgV5cc8vab9LuM9jrelsnFpsnutpdTvY2n
U/9LzR3tSVQz/at69pkdskVskzhRtEHjLHskJ9WpHBwWQKT3oHT5WithGR0v2D3B
v4VKrW5Ml5mWyIU6qyTr2QYmjrLP7jUXp775UnAuPjLC3Zy2f9gR+ez5wkc6WGdD
v7GGWGShUd4pLIxyRdQhQrI81ySUla0+KNvy/FQIcIUdrrGNA5wMUW4tC4yk5tfD
j7YWax5gHXUpDTldDiuoUWHRHKQHnMgsK5Cb8ndFQXCu65Egp0od24YLWXJha6Ns
ylXGh6gI4aIwjNXLkR+q3TmKKoAoYXHh0x3cm6GMzJUU7kbYZqf5MEbMrBRgI1JI
pksFdgCzYsQZbas3x5Q7PAiCXAJqUabXpJAz8lzOwBT7id0SOS+CEDpMDFwx4uiN
S5NxywLYr+bYRIIpm3TRFKdrQyi4F6XJI+Dqng08yHPO0Gg/I7e3VqAIz48zbLBu
c97vQhzLWMgb2IXknZhxwzH9fhx0QZKeNyiL/i6YcjoloZboHplqnaGcecqF69gA
NEIZLiMymDNmoLQkT/I9EGdZIpUqrItbQXTQ7USXUuFLhQaN2fEJ55pY9/4aDA9F
QYVMwrK0fLAOfAF9bU+E6pEOd0CJEEeoSqa7e5fNI+++O9jg+VZlfFY1Zwis/VBI
3ueAfxLHwCqW3odJBn4M5kKpZ6qarvF2OnJGmdEmBTSL/Hprj6VyQ1Fpe31K39ho
OaIp4CiWEDThKroppAW7+hx6Y69RdA+BwQ/oHxDWmaD4vgAjgtwU0WfBWo/GYShg
zWP+AioaxkAjaDdm7XcDL9EZ/1BQmcNa8xhATeeGynH8RA+Z3iUXmaHUNKT6WagH
LMa6DOGJzwi16zpHZg8sNkXEh7drL6lQz4wYB3oWLU2g2l/29EfiVMUYhC+pbJ3U
PuMDJBe/d92P1LT6crZhHUah6BZ7L6Kv12iKIhQSkajmyOpZFn5ccDyfUbMyIOwi
FAJ5AKsqzqu9+WBSz5SolfAoyL2NoqVSduBIZj8z3RgoL7AiI+dw+Wiiml2ReTMr
Y3UOStwEwASImXCHOZG0rzof9HLfX7qK+/8YGrghex+RhaTE2LxHx4LaTDCwHSZW
GSS4Z1DQ7O4rGwnDipBy7sZBrYpFYoJr6IY+OVCWWYXAQLSNIynIDWNjdVo/o1M4
q+dMZRoO9dLP2grlTKTZeeeVj7pl6SW0oDe/5IdfWyYGhFpZMSJa98czR3659dxm
49aFP++sV+ZR2Zehfqzoa7yoerzP+XiXGySCVlQ4iQA+TnqgiFsreMszca0OwsD/
NKNA1/ymyDySgF7uCyZMgTI2z/5Wlq1inhMb6td2AxTDZ1moQvA0WbN1vajTDCl4
dqbwQm4VUBEwSEBafgCLU/FzRsKmo9MrBUBznMDm0Rg5RvUuXkL/HKKtb/D4wvxf
nl7NoSrkPp8zVsp5+VxYmIufmi22U4Ug8oO2RBtF1PbdeQEJGfSQ4MYUZWbDAl38
VIjFHh1f0qn0Bt2GawohKcy7gAUlS+veQkhKy/dQFOJC3KQL0f4i8y1Yy600/Lwr
xzfR8KcQIiDQ5J3BDUuOUgqaB3p6hZk2HloLFpCAOnIKioTwSoTPIcqgFCGfoBtQ
R9FHOULCUe2i1Oo7zKfSqk/KJB5iamV+95CYucWyvBwUWVrfK974ZesU2n3lTIw/
0t0rUI7nelaJJ/x96YgFAkFEGZoTIErysS+vo2w5d03gIniGLT97YpBwZOqS+Qx0
erkbdNXa/xKtVo+fJVQ2vdRbc6eeV9SfkRcURfPLtViYr1pZ82tdt46On004wb0Q
LZgIg2ymcsfjKyRbwd+1qvaZyRH0pUplkUBGx+wb6RTQ8HyFA9UsaJPghEPvm5tE
rkti+rCk7aQBICBJ4kl/xf9ZZvRg0hYp9bW+uilJn9mNcNg7iifJqU95k4MetAyf
+86UiPvJAnoY6tKSNdv4G+s1BWAzaGaPQNxPzaBGfViSKIPzVI80q4yku4ODN05T
WJr0xZBnCuugcrj5OZHdug5ktLNT6RXI2i1zQOpbJj4Ld1nQDi7uLlDMOC9veB+H
Iaem1XPMNJNlUhECWakZVeZmJ1VuhoLcQ0+XKJBC2fFN6JJ2WRwX22kjUqxogugt
aKNZ3jFl7F5sWe1t0+YnnjI7ZEDevBk/edqSQP7mjY9whIcOG2a1ipvzbGAjSsph
39gdUZkdjgCLj79MCO4O0udm7yeD3cLKA9y89OwalWqWVsUWGGeko5bSVMsVwo2j
YYVOmVN3cY04H78tVFdz3xftqsYLPPscorWl593P09yfkMhEQ2kalYjFW2twaKWv
vQU6K/TApwbqe1WkHtwLcPeYTv3qE2+skZ9t7069DGAmBJBzOP88MLmJVg5RIbBW
keKCiNlqcMhW68Md0DrhvpdPj1SZ2s461gPyVOQP7jrio35qMrTRkP0Qo3LH9TZh
lD4lVAXwBQbNVMxB2GeeX8pRXVAtIAed0skJAvZWStLOa5cmBFpDsd8Y+w/QIQ64
kxwaitAJL9r9JFKgGL5JbqpgdGKvovpG6UX2BSAK0X1urMJ5P9S6nmr2XR7DKe2v
3f1O/EflyezbaOdA0lG+wpFI2eZrBylCFt/7EJYy7dSiBABRwMKcZd4pUjILifgE
Z29wVwCQ6e4Jz5RUk4lm5nSnjaabtyKyrUVrz10leolNbqQm3H23fqXyf7kNXvvz
5NoUf4I+ZdTmExxKJ/YpCB8zHwEkjibJ8ub2za2ykYc6Vs/m7hLk7XkR0lVcYaji
s9Ck+4NZnw/XlTW4M6kIvcgDfgLgoRuQj4VmHEf+bBNPJHwDoiba2FRsFBkMwQRv
ts6usJzqHgtP5vL1ni9i7PEuyJB7NAjl2ptYxqqDTdBJDMR0n3u0EI611jQBtW0F
IkE9YFoPXjJhxLf92YEMxyliaZD2jexrBHPm7mAJIIP8bYtsRxTGYnz/7cPT+Txi
M7taZi7nTjsql+xF5hAQD/yEQ56JYHzuX6whEohJW/TiPLqJf2JrazaYVNXuRtdX
AwyMn/5nkRnotul8KJurlvZrKSMB5PQgx3IRtRbsgZ/CVITot9fN4DPV4xkOh0wv
mVZGl/aYWbno9trAoMry18Bn+usbMIyaraZRCsabfAxjBNle0O6NnToEIFPxQIdm
7CNKRfHaFvl0TPQ6rI+zLf4M1o4ct3+khmaxQ94TT6vRbks+LywUW+K+Rbz9y1K+
XOKkVldnWoIn1P5bQBOFG+w0pPhpIwcJ6sM9+GCio7eKPdz/314t32MpABVSKUUM
pk8zKNEzoQKSq5LUF8LBfI1xxxvVHwTGoAVp0qTx7UpQr4FkhP1TEEiELDWFhhBH
7EcTwH1FUFGHwQwZiSd1Tt6aLHF79H64mg80kacPd9O3wWP2YJvboYd2lIAltIiX
92mBOp09qDEyeMD6JtnL3cC92aJ39qofXZ4UVBSu9ZIlIF1RmCdunz2I/UUoZ0US
9aRDGso81FOE5hghICzCYfvD720hBMkAJoYKmHD9ehD9JQ3wkKZOzmIBMixRvfbx
WcQK0P800Fc7lyYl7+13mG7C2/PZNT2RJ4c1fdxPS7LoeWxo/ToNDrzFedp0/R4I
/CPg/XeyGe1SfDKY+ibpEJdCq6ASQbXiCuxrjX8osTxfCTAXEbM5wxb0fHcJcINx
ZLxxmpMplaS9DwQDLkgwsRUNcdY6l9hljXne1bnwTg3bT2NfV8RZNWC4bbhKyXGG
a1n3Ty7rPlN8SVFoC8gzhJZc8qYO6rm9KQtggW8guhv7e/BDbhCVIXLnZb8HGzVY
ykp4FUmo//rsGULucjCLed14zICBvaJ3eVMLCiGB7dwUL5NpcLmh2gogcvGNvZ60
kvqNBIwpeOjt5WjUWMyLmqWBrmOzHUs8f00/e6fqNDWq7PTIiK3fUD+URVziV7yK
3ryYlSL5HR2ZNcZU/yKEpEtIieIy9Cp0dzY5tdjJJLAnrAVcbKB4q0R3x0CMc8+3
74HUjcxk542/Nwpja/0FiqsA0EL8kcLE472fJuDfx1w8c+azCCRK/a0OYF1V9xo2
aqnmuBujMy1+VSPqCepeOe5rCjzKB3nL6ia5dJ54QFLNonEdCpVgN10BS/vrjQbX
xhkuGeyWiKS1blIU8IKaxH57KgBn52id8jfnk3PVNrrWWz4gggBjakKhPW5Enbji
DbfbHtzCpulL4AVROOhJDTjxew1tAobp0D076ec26J2m5Pm8WYzdENJwUZnR9zw6
YDhWKTDJl2CO1Qlx0dYbMBqOjBjTOccdtJojnGHJEwI3DIr85Puph9b87GGEOLqe
+lU7Bwh3zugD36yCqSocRdU69gJY8DnR9QoLyNv17x+x49ArkhQNbcmAXv9soq9y
pDPILERxIh8A4XXWBfWsc8L1GH9R6AetRyMkY56S6I6mrrdXwQgUrn1szyHqLMtx
Gsun4sMyky5QW9cMdLIwZhRvZNRovMR0wIuSgBk66vKr0HIROefJEhqxtyXzEGm2
3GLlmu1EkDUMPzJd8Y7bnXUJijt4wh5Me2o3cINwKZzdLFQo7Wu+x+vW/DJBJWjx
lhjIyncPIT+1HvwJWBbD6JugW1P8Z2HMXLRxUchnzX2D7YQ0SvrvFNYstDPSGU4w
5+aSJflXK0I3X2VXpYJemQQs5lrejPWxwOtFFk1f165TLXoHg6WPAuV4ZyYKboOl
sTtKbydQqcnFAnnTQlbnwsRUqv+OZGzXWL9kM5JA1zJI14m8awcbjRVmIZrKChSo
OGjy+EMJQMhjypKvWrkxZKeTa7+KUptTd3OMmCUca2qYlY+AEwzZN/Yp9rAwLb8L
XYO9FUuuZAN0WtzlhMMqNxai0M5BKOz1g5E5JrHRUv6XC4EKfy76Z2z/MGW4zpxq
NxYx2SkBg6z5qmusW0oIlUh7D2usXUX8oIwXNKDl3LJ7EVtheweuw0DacC0qzQqt
FLPeLqQdGQ5mmeMI4+ub0LPSS4i6Xr1X1ou2jC3+lbpW5M8LyUJclwwgP/BOAQj4
DVRGAZOHx6NWvmkPxiaSf6S7ftIrZFuC2G+RkwnuDtp3vH8njxjS+VfPBmNeIdet
0p4fN1aFvEEjarNYW5fHhfFWY9t1vPqS1Wdrtxkdy/r7p6DHcg0DPjGz4FmKKIK6
6PuvGKcLoFAkQOaJEb+ykemvFYAoaB24hCK899jW029jMhzf9pOXkjrmd/25I0a8
5myTYjugxXaVTHk2hjgTuMGXIf3c3rhqkOpMPmGzgDYE0imoU0dB4QOPtv10vPCp
Hzxts3zs1khz0XlKfojDoS8dSaic/sOQCuiRhLrW0JCxgvk+J7tofH8p4nyfWnmx
o/dTKr9OiTdP+8aG6s5w0W6sVacQErIp1udWHBio3HFPmVVOn3wOKwhJsOLjqfc2
zVNCA7tZAIgnvrFFOC90TjCJTVP71r8xqDJQ1tzZ7AfzMwjMTwSnIqaRfg3H5WWk
Ie9ybuHKKGhU7ppzmXbccjS/IC3ZIrB3OcTW9Jm2MYfaCxsx92HZ+HShTmg8IoA5
htOQX+9rqmwrALz4hnHY01DXFt+v/g9K5jq1j9uJSNUThQk4F2CsXfHpVsOYO7JN
mwQ4VZyFVQ4xRc6MiOBqnxLMTsCUyeo3vH6FCYT0S+t1Es0U4OBaAz61bVZNGtiH
t7vgqwtoUbqAQDBrjSZjE6g8ED/7I7nPWJxBykEqemtmU2c4BfMZxQJR1blUJP81
Hb0jyee4+3YPJzyzeYKau2BytwK/PvrqmIQ7psXtrklcdUSVKqwd4V43QOntuBce
iPgiYnxvZg8akd+b4GDQ7UmmVszUukGnfhIEsLwoHKPRn1u5VNFDPcLhUMShgOP6
hcHlSmgHnPnO87lVxVrmuDQNAwMzozzwtXgTS66ahfFGwkQPK2Clf/Vb+y1YIqpB
HlMOaFpy2/LbWABv+VsLOHEKJ7tiJXCJhg5co7f+lll+eNFQ0k+xF4ZAagkCrSak
54NZ4Y/JHAjwdL2OsLuC5iMLBuUCE5/pwo881Ga8pnQpOKIZoAY53JuQnJVc5IGe
15uxHzKYPFTzOtE3Z50x91dBUfD0MaPyf6dgmfSAR2b6HxP6J6dA0NAxB4KAcJA0
xx9ha9IbTgYU8WYPTwz3JNjx3zoWbd8rOJXWkAibVeNJOoa4Ib24ydVE7csTlTFh
ijUiQ0ZHXKc4B6YWKAn09NU30QrAEool2VJDc1GUdCbk51O/En+7z4m9JXM/AcPp
J47wKf5bT3TRsQWqhNap2ZOjpE5AcSd0x+LK3c8q68hzcHBixWGUmuk/TgVWUZjt
MwqB8B2ZGsxI/7DlX0WVIZZqccrmHNKACLVkede8dFJo2H41aIc+gFLHdZHpo6+U
Ru0ZhRpy/SQB26tNteWIGlCDJ4voRHf2G4NfRtp41Ze3MtZh0jihy047QyJuHAP6
/uojv7la6qZwIIfp7e688mhH5iL9ZOuuRgiPGg39T1anXi6KgHsByrRLf8q2MpOd
BY3wHrcsf7mu9V48jhh+VKdfCJHbVzhFp2kD4n2t2s8HhFp5f6+gaBYeqftU7kfF
9wePugsWQqMAZ27BvFBTPdCKcVQiMh5+jwk/vUWCfbyJmKTgMvMVv985+/0HF0Lv
l1pcNQMxLDuLFgoxgg0BvsrYbVh3eBroCpDjkR7/o0nfwvWs/Ez+vrFSw/K7ni/k
k/1bZu4ZGQiHB7K0hLNrgN7NwiR/562AZvJrBtp/emNXwUrAaAQZszlL9IfQi7It
i0r1DflZhPQpU2SMd/Dgz2ffdr82pVG0dvESeIixSDWOuTqOLmwEJxBwJufWgGaj
eu4RdPuRogisxKtcAqtE8CUNWA7T/DUOufNFmO6d8tVILN8+qqzwT2DXII6FZV+I
7bGtcH0QKVPh44lUdppvvAsdghq4dQb71DuboLIWGKe5XzYoOBPCO4+p4XMVk6yY
wLJPk9wk3Fr5BW94jrryghuRilyvzdsL0KtVgtCOD2Ms3YiG2YOIXVyy6qBRM6Nr
XQi1y8OH65s/NAqI11b03hE4BjLyR2O0WbQkZ0QJPtSJr5kgnrG2mc0aRD5afsj1
mrrKD5NAyA4JJ16CGOLKFZDMdUP4xb/C7zM0xSAtJagO9ZcleuRf2ML6TYx2rtjR
qRdAViZKROmvRpR8KRRbN2RPaVt/X4Ysnat01N2U1212/QEgAYl0PGr/KSxPGpc6
TZM+Km5f9O/zlZge9SrThG1xyX0o+S3oBclmMQYyXZirWoI8GMPJIKSg+nFVnUlC
eu86cTfvULHUPhfhw3VFsFn+/rSORFloL2t6BEa615se9lKYFIlOSCf8DSmyKIFM
BxnNgkevYi3/ov/w/u3TXtDVBgN4jOaPMOU1PyZjY8rDWGqwXuCJ6rUWY/xS2e7l
BXNUNwRxxo3xWpkYQLHUM0TKuJe5kGxdRU+qu7wkmTb0ujWG8l3KdKghemJgDFxu
QATHGFYtf9u+BKFdhA23uGFim0kxG9k9GB8ZVVQOG+L8EtoyIaPH/WIAtR8oQ6yV
ivv+pbndnM2GMiEgSk5daRYJyldum1/pgcxxjypDGvKIevqr6Yap+KKkJxddX+wI
PFOkaE7F5w4SoQ7X+rbtG5cN5bCdkBafzCvaUJC+gHIHpYC99QIyqLlhG8/FjeMz
ItEkJa+Pi6GBnXQwCj/Frk5iXaghrCOQsGvo1PdiWGRPXz694R+jU+RAh+/v+fcE
OVmJphGx/CDC//7YmQUtlVBdX+CDZFNqkXd5IYlxsxL3+qEsr2QECgvLZLWc0lDJ
ddfCbzKajCtd1qFdUaiC80zx4da9+siNQeGr2eIa8ppR8L33iWlXytYDn5u72X6t
MW4I56nNJTtdmP2EoDPgUBT+TqWJOqX03Sx2W9Bd3CFNzWc7kyuBmlZxMP46aIfG
O+B8dmSq0sJccJW43K6L59oK8A568FdO16lEV/BcW4nwWUG1C2nu2BfH/Gt/ndmQ
9IqI2cWx8CZgAMSXTBMbLstFRgx9Ex+C8SIqhz4hKlxn2VAM2+pbbMDkhlKsmkuf
EzmMDPktFQ6oj6Kr4ggPeQNnsbesAqBkoBIusRh+dz9VLo/kF6/6zmjgPhnugsml
fyrEErpMomXJW2+u99Y5sK6ZQie25lTAlQBwBn+pZuTZ+/VTnURQG0xUrubpXIet
4WcgMViDIlQTQuETuvZdYJYcuZVh9Rk69cxJLfxwaAURG2gwVSr66Ms4rkEBoPJE
pmld3lg2ZiTSucBSRrrNNPOWH7m2O/VnBnSJb/gKYa2vnOj7BkcF6/PyJFrd8f7E
7ZOvezLhpQxpm3bfARjuWhgvyBOIedIvFw0SNDcUI3644/7GOcmR9fMoU0HN4Hed
FQt1wxPdfcHAQTBXg0T+QOBj5gC2w6PdNAkcRIgsWeTbjVsEPFWbZKSXrAIocL7c
0VHjxpzGE07ux6Migfcuy5l9HbEYE0u4yM88zfoyZf2UH2TPb3xW6IAn/WruzFxM
ndIcCEb4wmyvCGR3fOitAcQynQGbC2Gkk6FjyFaOHwDa1okp8lKkbtyf95P46FFG
k/rTX6qcIuIZ7i6XP6gzzgq28VmM1wTYwy7SOLiuUy3Q1P0pBB/vs3U4YeS20++S
G/VF3t51LW/4YS2lo1ok8gJe+BOH5iT4uSrqix0xs4SuCi65MlodPlAxwhxAxi99
FiHjMvEGQSekP3pZweSGqsR7TSw9pDn1ZQ0GdSSvK27MVDWq1PgVM9A88GuOdzqc
QdzNvxdirA8IHUIYSmcEo6+lGCgZ4NqYKTY5r8DpIFkTcFEwdinpw5x+jdgvCDu1
RxCf4NEMLdWq5EJ7R7/sVFEcmlX23NqwDV3fGU6A3eIoBMFuXoI705z+sXlejI5w
9V9YWt7XlYsPr0eI0w6duDNmhosU6Zh+sVuJcjFwLbslXq20nOfX2Gs3gyotflwk
AZ06fxTO3hg5v6730P590ftbnDPgpxPKFyE8/Ue5m+uswRCwmAhAViuUc6byl7xK
N4uC/y3gsMEvPnWP2UEgZoMy4cbRDW6z7b7mMshCrLd6QpisJ2Fh1zE5anS3hTSY
eltLJ/HuujTyoGkHUXU2sVn76VW0stLftETSkGzvWqQYYPiGKZfOadDndPqtO9CC
Sy5N3XE+WSs8hyjxNc+sioN4G/E2v+A3uUwh1gaJtoqx4AD5ICoce6Sy7lSI71wi
/mMroV8bimJeu3815UqK+/tTrKMH76FnJQ6wDEPohgytMKOOtwJKhNzSuxn7JzeC
Dmrg98EZW7HiwGufs3xk2PjXo8w0/GYothNFrUQTShzfIBu9SUtNAgQ39gWstnzP
WtY3rz/WMdFsSVUr2QWiEua0J4/3RsVhATvcZPI77G+ddILvZTcV08pIqrCuyUzn
WvBuupowWcpkenqWsmNINuvykCORwFd7vSuOcnsl4+L5JwTToD0wu1l2c4R0hNSz
n//Wx3fHkeGDYXwve1YUQVvbU3TVdvH6oObGI+1m8JXT9Mpp1j4Dit8/oHGTb+u3
KqylEty51m66jE7R67YxK0HpnOHJUXw1lA06D2xekCEwRMrwKAyg5K5bW8rlLWGQ
hY6+cDfnyoxfic9fWVIlt3QYB+/WCP7htVSQLHIbzj4+ulJJMWvoCDHfaz5o46pY
UtDdTwyKxzAcL3LGidLMD5glRGRRC69nVSjXeVWI9YE7MULtGGLH3JBH6fOKFGeq
jLMCyCU52Tt9pIy7fjY68wHDFCNMCtnn3B42jHRObrZLelD2+jroRBl5R86NGeZ+
CCmEFbnYdjpnfMo6k1JCKYR0AT08FfIjgXfGod1o1A9jLNcapVF/F3hPxlex6M1u
eJPo1S3FjlKVEYIKc6dg4+fV2eWcVw3ClZl+TfismQw9bRJK/5HANqc3VNt/zdEq
jb3ByvcdKpgdLJvEF+D3IYCGSRjhCJWzueIK+411FZXPt4Zta22mdQqyaD7Vj5wY
Sgq546iviVDr+RK32I++1O89sZIGu0lsCjVWrEpRZzwMifATVoABPNL9CdsbFnuD
+THTVOEkSrvCASGyT69X/oWoydtKX5OfpqHfNliNVZ/rBgKbekPJOTBKSNrkZmEB
rDiIC+Ujhr4K/Rc510nnHLUHfzbUnOs7k//YIwABEdhwhP8jxqOrm73NdaRouBOz
h3npLuTfd4agQDe5Bw+VJUA0skqTt36w8YmR5KXihguBKU79PU779TkPs5omwxkE
GixLgzBIrEUiSBcrxjRK+6qg8EZm2R/qa/c29Q4iVpCXbnWwHeqX905gJPtNOJA1
2CppZdvPasiuFZAHbKuRyITCNnADLH8pnQXOQ2XLa6p19xrHcI9VTiv+I/4jsQr0
cTWg6M80NA1KgTxDW1/MV/LOjOf57gmMMqFFdp+FxvY5Qh35mTjwMFIk2Hz7nOSU
oZ2XTutFcpz14KLWCSVgW5p8MBegvBqe2ctDI3cl36JXbM4MQWBaNHdoTMybHUZD
sUYD00vkKKG+6miZuPvFgxjHcUYSi//Yp+OoxJnmadCtu3BHzKJV7YL9TKEd5Co1
OXDLqJnuBuioDnbXyhLmtk8sv17KpzWYLEjzwGqIyt6NfZim3Y4EddgZyDNeczJA
iz2RNT45jc5xVSD0oW3tZjS2IGHrm00Qpu3SMk4HplwR1nm74y02tYBixeDnN/j0
TntI64X0tgY0eBeJT7bAq7IiIbRlw6lSd8l+g4jBfpUqx7jGis47C6VtyTMnq5yw
4fBf5vcoZoBDIA/xjl9gijqBAsAeQgU1bHhy/SY+2O9bnTsCoKPNXonr5OWi2Vc5
mwWpSiFcfgMpkie69KPwXVGoCoMjx9yNGEpkP80pWH6ltgKDlZofRXe2NMO6HA21
Gt+owfskpw26NfzfyndN3PEk4u+ACLis/5BdzFNEmRyHcfVcW9520toXjN037lWV
Hx5+1K0s3PXYfl8r6woCcdYENNgg0Bao+/muPtiNoVUAe3xHI4swGwd6E2tf1xns
LIffyg6thMr15RRUDUPuhFVoRGx0pttTrlb2K7i77bPLINUhdGwuv3bpoch9RfrA
+mdPI3Y34tZZDQJj3q6Z/FqTs1TLT8OHhhpEQ3LMyXzMMIbVEd/kPdO+ctx0IA4D
DfnJaxp70OCKR1pogqnHjGX0y3Jgq6OLVU4jU4SnLJyDsFZFEqpUPpdgtkj/weJp
7slLnOxyNS6Z4txSZL/MISnEgCWYaiM15g+g98htvNWUoOsFzxZ9KTwQSc4dq+bL
ZF2puFLWDo/3yayDvnNRE8WT+bJ+lhOTaRofikGzu/d0R6HbMLVXofOjChF7qqhU
i8Gt6wH/v3pOe2QSme9TErSI5gffR4l8MFeEJ3MDvBLoLIV+M4yzZjGZBmEccLyJ
6BC8Q7RDVnp8MwmK2jRy3DINeFh32lFxC0A5s7vdAmZISOKLEraCuICB0GhVX1PX
zhxXRUq5dp6mmBTcVjJ0npfKXcM279KxKu4GBom3b5MCwXjMv8IWZduYXw0iosSz
Yjkgtidymkx+Ob2cSh/dNcvu+JP04U5LQAZ6JlcOWPzL+Xtt+2YZmfYSz0E4PfC0
eJecEx439Ry9oDO/psZOpZTXH/zYA56mvPMWiZxgAKymjLndcJHM9I2eoRI4Hcsn
k+CnKEa0mLnsEfreNDlo6QKTTFUPOebRUl7/khGvxpcJg0Yf4GeKCuBXqC3nZjQL
ejABSRhHrXu+MSasc+tjGv0TSUYGS0GBT7ybtCbWjZuti+VMHwF7C2LX4aFFT5Gq
ISqOuujws5lgWAbhE5H48XOgaxaAUQSt/26kxBBhgU+lBksClge4+nACROIr5IKW
u7wZD0C566z0gNTRa46INRgHBnMDuHNdQyZ3PM1uLpnCSWf9TK9iXZN1oH9rJ2S+
H/Mbm8wv5A0GH82rmeXdTUxMQq2w5G7oe44NdYYwiCYqVfAX8suKscw8cenM34CL
gltqe1AR6zYkOTOAhjlJaYHlzbQg6fzA2MJvWYD6tfnXeCCFjZ7p/OUr/BZlF5DO
zBvU4i0hG+YGGMiC29bpAV/GhgpzYMV++RHzVH+ElsQXYV6ThYtSuQ7T7Z2T/F1N
E6CsOW/EJ2RAIzXmTt8nRj1WAC4fzUkXi6D923wkipkgFQBelWOSNi9JepKjhRxg
zdj2zCfZEYlGcpHdTpGB5RzvHMCRRDnqRumTNM52jjskuiCJqtPVL+I6L9ppfT6i
elX/pk2EXLZFoAj4tjh1YT/64rK0aeCSJoDI/QoZGe4O8j5Imh3XiNV3bNnUnV1M
KBMaHIAmC+3EMUjtrdwER4U8nKeAaDcmmZHUSwBSUPFwCa+hukuV93khOuOaAuCa
7RaYJwxU5iBLF/YSIoySEeey7KPKNlZkBemyfEA0z0ibwfIh32Wj8M4nihM14zc8
0Zc3k4QKxifI07x2PY/WXbGA/56xxV6330qYCNum4wJrJXRXzWZpH/ZqrrvQPvSF
ufRfYuoFn8dQXCbK/4fAudYfujIMCZ1IrIfb5vIYemM5j1bxYG5SDeyM0ZaBQvOT
5PNhhPwCsKCtmH4VIbLZSdIvvnqsAqHkK05kK2ntZW4uFvpDuAGrfIuP5GbPxL/O
ATD/iko271pSXvf/acfG/U8Rifj4SoK1NCPTwQaWbDiDvHOUflFW10is9GxYlDF3
CnO1YceQWmSjCpOH1zbchIMbJVJgbIBlmC22xoNMl6Bxk6EtDLEzD4GXTSi/CC20
ZgezFrrWd5o5J2ZJ9BoPGh8PFJnEqrX8o7aN5O7Nj1pY7F/LDH8py8OsVUrsGd8q
RBhe5tfw6XKqHp1/r3Fla1gYNgqAN2j6yq5WBcw4wgWWksxuORy5tauIZV721KBO
gmskVF6wdNxDUPFuPMXbS+9HT+mQeI9JBGO3BXthwagAlULfx93HUJ+dfbqPLnIQ
dDtp9R9+oeVrZXl4BeK42UMEqqU+0Fzs34XwiE9Y9nPtXoVKhRPK3RM72AL+g2gA
Ll5CrCaGChisz0BxV8bwnIFfhmr5X/cpl4v+319iD16/SH1Wy4hLXVp56MO0iikn
YqGqAgTUZLf4HNjpmThluMrFq+yk21OcBKZ20B8V5hrf2O+kNJLCkoD+LyiM8FHh
KnStGqZyKywiSV2sX49qJp4cN9rCvCkTEwuvdpLyRRF7SaHM/kHUdFLZrZK7yQJY
RfMAJd24fgkB4QZ8/JlS/xVnpfWifxGA404vfmjDvL4gkGweyGcM6eQPOFD7I8Xm
TfHAK9EusjOGMmUr+VLM/0JLrbKhJ8EDaUIxZ/IWQePQsNVj8yH438//983NEk9W
Ju9qCW1+QkJZn1m8dY6FG1kL7UdpNT+q21reQ3lE1hku6+AWESAjAc40nAJuUdN1
+aVelwOlXtl2hTPNbRtJcw8HA5xPVOCyFM5t8lNmhyFr+A1fA6wD0vFor5Jya1LR
D6M0C000Mpnj7chyknFGhjPGTRXInf+kD8+cH0BfW0pbpwyltLWfJNEFea53TnE7
KQ8brUdkfFdSIFpq/c41lj5BO2rOMSSAzwETcZMGxKTBS/b5/fwT/pa5XKf9FNH1
YfhoZwSkp18EXEFiJw2p/LuIjI6MG6pUf6CVZo1AmQkAq22lPg29U0cLvGYWgFgt
19bTvVYGnaxPgnKY8fu0MdQAle6aXiwxjhfU3DWswxH1t6egnd2P/NoJcj23X0ro
0nFurcBp5tnd/H48Wq96pQzmZArmfppGsKhANTxusohCpBcQVlbrk6wWwPcWKGsO
LAvKNrrEKmVbcRyNAKqJYk3z3SdQvR46+RLSbrCTdAFjU/CP40JrRVpNgQS1k/5C
D6zeM37EfUh+wFLD2GWKPuBw8s4WJjcVG+O6vs8p5T/RuKfs76mBHwicsV3ZtfGK
jzYTxJMG//Eyw+1qDLUA0yKuv43cDX9sLetBPs+oVa/FgFEBPewPaCfoqdLjooqO
WbjkkuaZu/ar9Z+RcA/lY9T3/beaa0uT6NkNcPqaixTPzXY8WhRdQknTRpbSLJbc
JurhXwx99LTEdf0q/oLUTSov8+qk+74iYpNim8A3zjEIXHWomfTblLyYBibSY9JR
LMghAgNe5IBW0byQXQ4ZBDmYueSdxcQRqY2gyRwhtGgeGhdylu6tUnuZl9oDY6u0
n3Z28cglfucIRmvCxH3eJa2gk42qL1pmM0HprCGaqg5u/qX4JxmSp1JGVtCI1NZw
dxJj44sONXlf0dcQcPqCIYrq06M0nZRqSMR+x5cuW8qKQqtlBGVbCc89Yu+Xp8KB
w8c3o8TXCqFdk5P2dWddArcScbOj6YXd8vxRjv8PpyM7vuOutk8YV/CWzaL0JlbP
ZJPLfyZvyR7y9D03b4TA4E21gZkXcQawhtsIwuFEy0PX1ANyLj1p0CRa3H4aESAX
jbQo6wT4BbmXsr80WOCSQTG9NtqCf0Jqg+FBGT/l9Przrj2bP+NJ72mHs0IwtmjF
CJZJ1W3TYqcwMfjxUHQxLdbKJToaj3cSR2JyCRxlZOJUs925QqWMAHuyWX9UjewS
bW3D+R+pp4/hQF2CwTLUj80k8guO3qU82wXKf8x887a6ep3t9CCdHevMxWKqm+Yd
aSexgTkB0Y1z6yePNfBI5bwggh1uylyAI7ZiOnD5cNg4rykT+OF03aJpBxuVWk+3
NCTHmYdOow4MamnI4kupG/iZq3JrEfKAisNbIgxuHwBvqNEvr/hvBGDwqQ2amZv5
EeeWXn46AWtm1JhIrdt66iGFE2KvV4HuBpPvg8YUJOezSsUBxOYqQAymxgJjol/T
x2PpPMA62geS4ka/pRjVq9wFju8uGD8QAvcH8SZbTGBB/qSVILtQyUTqhFB46WnS
01X2ElJQUhWZFgUZ9yM0YZxPB6h5Ito4x7FeWcyKZu7Tp2dZ5mnu0mtcWhzz67F0
bFhGjgAcR1GXYLJ+UivVgr+zcE8SNe5cZY2+raJQQJKv/CrFsEQcsQagfPUjpQ/O
NLp3O25kEsNVo8Timh9n2Y/e2H1wRJWCPZeyUNEfLxZ2FVkK0CF3rJlg4m4BiFEH
o9eyAorerU0qrxNFaoQ9yHGFx9cKdxVCAMxn97JWhwAlZcmV4mbngDo1NSx26VP9
T49XcNFKND8+ONfcy552RanQFaPbKh+yCSdJcpZupUVGXueytPNJafON/wUemhZ3
APXhUOulToaMZ5JONexr4y9XlVgbNiZdxzPIUKFkEtY5MuOOSr+Gz9zCHNDKvwqo
M9QItqn4EKqtuHiXtarR2ViJZ0QRzrPwStWI3ig2whSnQCBlAKAGa043LkyDQGXh
J7bJHqJJ6JW/bT3zSU9hdKIRD1fXzWkk+lSF8PcqOwkr7vrlYm2i7caBbpUaF4ML
Eq++0vcXKflFLGjutnocbpRnnDlxJzv5J7BbD6iEvc5uY0IfAu+Jlvl7ccWr3cfR
khn6g8CY4gZMqoUJnjBHQtyzFeqXvs47Op0bqkMRSwduMfBEiCzeHfbIfTq3ZlQy
vmDXVsTNxbB87lS6/h65szaenI+8/4Hnf1EviVBduk40cNXayV45o6vusKg1Zenw
e44tUI6XtUlIUAD7p5shkB89GOnF5TCrGScYpPdTvqXsS6+uJeZ48D41SXwpcAeV
mln/x+o5ykXBDEeoyiy3aOkdbDiBFDsHXglxWIAgxJYM4c0rxx7b7Pjh9Mu8AQCp
P5NgTi6F9cBb/MzqoFgAY1xWZfwJc0QN7utAHjysG1XzS2X0m3JaXD8AoAeHkhQ/
BCh/GiZPOugMzkpea5Fdb7DmIF5R6g4GfH2SVpWY/+bFEXvb0EpBQSqA1kYVJDLv
gcnccp9ebOhVLTyiJyia68sx7AkXHro9qbsrNsDcgdz/7YrroJ8iywlbE1ac1skF
jf1vhNi3R/4ob/5c0e4wmD8ZhoNoOLBKCKXfDzDLbNC9crzafSIbmftV1L7sHe/l
9Vn8bK47gHldLsfuxM+4TcaYr3gPGboE5nH7a1CdE7FqHLhCusAwDWGracjENEjk
nt2/dG7BV25Nx7B/JrFCOHfMWedBiywmdbq2v1VsTSBV0Yi57dR1966ZTxtphwd4
DE36mJ+c2u4Pqn0KdSK1xOYT42Bx4OXkZ5LHqrigRsJETMXPlte9iOCJiYfLBweM
4jBCB9a+Fp/Sv/xiH6bYcWndxtCp/bsA5xMSOaXqZ8aDLdA0DxFlSuMUoTMKDvHb
8l1nLa6SUnJQkUItUx1g/OSZ4vgSep1G4BbaW52MJ3kYBlo/BcXJrvh9vHwECKBF
AzjAFLC25INwlsPgoBF1CR5sbDKjFgtjdOws/AgLbaNxkion7GBGVqcTU2vKmM2j
hI9y8wsztQEwu/ZZSUEAn1EV5J/jyYYw8jom4CiV7kOWCmvygjrKEdGpewKQQmo1
TNS7xX9WP7GP/r2RSQbrtoxzavP3JxHWawV7O55A/NEIOGMPN2RUBVdZSPQr4gPY
3lyE2voccTYDka2Dnh7DXury/1CXgEWgjuCno7SVndIn8phFD+MEQl9oY4hB8Wc3
EXFpUmRTB3tsF0Gzm8JJ1BdmCn+LliuyHfsr9HgDpfPCAU0hQdpNmHWUP0vIOZCb
etXrzfIKg1BHQ0VBNwzJ7utD646a4Hdn5V9DC9IxqzI6I9vkYXSDDrHVbmp5t/IK
41ZxT2GD/Ol9iOFeD0TAuAkum+LP/TdHZ0GCMyKyxDE9aidvBqg7ThRp7dU03cYb
B1PVDX24ljgnKpCbklgC8MDhFj4W1xPJF9MLiGRqLzZX0LGkm7eOLwsrURy3aAX5
DmhEQcekE/1sDh+Mvq0Wno1wPpalPpkexh34IGd1/5aR5sVfeE7SnHD+0N8VGCGk
DGgCHOo3CnVN8lu+rDU5Qx0sHXfElig7XDqjtriXLzFz69s2nRdi6iujB6nC3788
1Wa3MqWnuyyXaCWTK/ZhFP5DFRBWvRkPKsRXMRmFBy+VjMg2iGAMuxqE4yAjPogD
56iMJyDu+Ih7MSGV0VZh1YA5xJUNO2PrCZbT15U2cP6p4X7dnKk/2pujXul6ymy2
vnRVXxVRuElP85C2GJvbWBB+DfYqYrO1sy9fjvjhRThhATTYx3L2/iFm0nZ3hFxb
tgw+IUZKaDQSWG8UVPaoEmlJmGEvPe1HcwuHhDaxkWW2z3zvQXS6xVkeriKtESWT
C9+ec2NvdKJD4Gk1XSjsNxsmXkfb6MAbD2UmEobTH2PLUVJp16QMe07vIQi3w2hV
pRmO680gXz50Q/f93sJOZTBgPHa7yY4YNyLfRVyQ7Su8gSXPR9ZuEWAiyDX3BOAB
Pm6trOtMizs2zJpB4RhJVgihe0esHk7haz5HGXVEiccdn7xWlazoggE/CaBhmOnu
nEJfOnke9rAnNorzziePuiMg/UEH7qZnTa4DUD82CGruJ7kdsAaFNR//NIZeBaG9
Yu8k2YuvpePpy1f6KhJuZ7lIeuiFhzYCiJc3B2rGRbFvTnM3ww8rlfB6yStxL0Ls
UpklDKgkKdS/1guWRx3ZNPoR5F6bB5iyV9/3R4a/XUEgraihmZtVQHVCEMawx0f9
9Rxg9p8kgTyP6akOcbUVB96bsVuxP/w5JWo5W5Tmj9jTEdoNctfkBNVgpzO2Y2u3
RmYGFGCkuR4T/epxZnn89j/vP51krn/Pz8IoG2I8rO52v24jieH0k63ncmfEFDCe
dgi9cPdJaVaCCcdM7yWOD3Q3HXl/Q6Px5C4ACOZ0Z1FiYyceeMeuoCKdJGV8saEb
yItJedC7bk7Rd2u6alrZOs9DFK14TihUaVlDvlObym+2veC+M/wW4HbGcZUPuRJh
urM9HHY5L1Smnvn5xjW0gNbpnbgNYCd0/JmKSMQQ2ujTpyp5pb4M06N/uqe6z5tE
vtX/JZ+uUHUoWUFg+IjeIPQPQXcdKaeNP6ySw2ELULGMx9SyocJmoNb8UcQshP2j
7gs3EgFbTlnXnLVFujqG+zHaLiW+leldQ6RYCnFEvdi8/yZw1TFetV/wAgbq0YwR
VdhZqQRXIGHrJaZuyex54LwqwBcwk0N6ShPV9v/fNV3ZF2eeevj13F2V2kZB1TkS
IrdW/NezxFZxgIoUQjU1CA3NJNlIsZQLKUhXsWyGcnUdZMw6JGfa8SqJU5MLjS6u
F+Lk7OggkqHC10+XcKx/djYzJxZ4W+XrrTK/XzCj6T16eI12/t7UuG+RFyC1+4+k
+rK+/cTXNXYrHKRUNKQjVQAOLCxKsgAtgPaSVZpo2o9dBjzJnNRU2ONy2fcJXMnR
u3FxQlhS3yjOdVDgaqaG9kZTZmXNu2PDA2HrDPYfFYkeLTB30ZWv1UHPjtMPHMmk
N2bimXah2+ibaVGQtaQCJZTofJI5NXwsrLAZ7vHlEFIAbMqYg8BN1KVnELjshLGT
lH+kmf3UuRe9cwijAQTIBIsCn0MgUdghU9Xa8X5Uq7pqUVB6zTravRTBXy/OPipn
JKzurgJQO94ZuzmwvCe4deShW30UFRetr5QlgW3TbyyGw1XIwFclnZZzxZ+/ony1
nNDYr4OjzMFGB8fscWshCJRstXNPfg2Y+rpCDvoCVTjp40zcqh2E4Qa1KJrGR22x
0FosCETxNxOyhOBLhX/+9XaohRtV5H8XN12nHVplLANEC8qzFLanOdDzvZdd7HuV
v3JBeZFvWf2pFGayHfiM4qwp7FY/2vc1Byfb0NT2IBznUkqWS21jC0BfQFiAbzSj
I2Ao1udLZc4S1yUWqeLhBTHENS2oLEQ/IT76Uy34i5MY7NRezP65aNd4iXgdLcUt
mIUHES1nsosEjjC6UmQFUq7FD3v34UzUhXAi5thZ3Atfl6FbDrXs9591oUNrrKnM
l2IBMcN1ZQ7SYwrhtqygWvjpmADVflFDAuBwo0wXo/EKR3fMtO7kEmwXTV9uaKf0
cFQXtQlKgAHC+JizldOEs5RP7m2+KhBxoMYCbrD7Xv+2/+WhYxSD9dujbxGCJhsD
mGwOc5oU4QmZB5HZsXxdbEmpH2eykXhCqDj72J5f8ioX4h+I+9YPTja66s56TYUN
mzUfGXGpyY5XzOW3TmQ0pJS44bCg7FZ4nC/3ex2+hqa1bevJUB18SFdtjb5JXn+p
rUvrpLWAbI4YpiNGAPpQL+y8znUC1aAFArQZ+MAf4Nitf+VrRL5huSyyO7WBMCbj
iSXOurXqgGYHxpgasJGclEqd5yw+0D03PpXlWsiG8UIveixhAZjRVQCMx3dLjMsn
76ZnZQt8UdniBG5TVvSoVxbXsUTEFaaZ1c1yH00fCzBsTJprVP/ETZ6iYlNPmKvc
zfEFsCZYel6xnGS4VKseTU2Vn77rOlN12dWb/wCbYZB1D0cHy38pOTwoTdtXwZ4J
5RyUTxMOxrmPztYEoys3TilEkiKBxK9PZoCur5GEFa2PsAurcNnC32XkDk87+z0s
+0KDVhq1Djx0F2ebfCCclb6Xu2HJfJoBojqlP+jUV37inKkw59+PFLATnuo032y4
nDJIFh1VFqAir4GQGclKN2cZMuzjIg9UD9c7i5wsKLy9qsbI8Xa11NPMSfOTlbpb
6NIrhFJXMHAPo7Hlk1BWrN6UIACRG+JgVAvb4EjAkFOEFusLBeyqplh3LxH+v+CF
IMZfiXkKJ1tXFCX4Dux0VhzYDlpQrT0qK5BiMQXBIAv6qQeSKmHW2mM0o/i9GGcl
yaFnMJhKobn2875GJbCeA4P5aQ6Oj97oUf3JuOJXQdHMDFFmNboUGWXeJ5und1D1
DgJw051JenMnsLFBCsyK8/Wh2HLbevmdzEebeqZV4DspPmxYHPTH5o8EI7GlaUoa
IlH8QUq2wevwrGaJBTp6UalmuSwPIU3GHnNh0sBLjnrfhUbfJCdFebMaLtHNeSue
5qZFJWxswxfRSyJ7IRfFAfoc779Sf7TgX7RilPYbh2z0jPS2Wqy6Q9Z4q7viiVy2
SRePE8+yGbYzTJcYfIj4sD5T6xhA6OlbdU2GNa/sIrPzSDHiCPOeP7wQS2yPZWsu
Gf+GLO37iQwHOZ46r03evprZhdmv6fhs2Zbm2qXKjbxL+47LZ2PPNQdyhFKvp+eC
PuEB6z0krby7iZvrvQ4T3nVPkf294Bs3f0YDK8U3kHqz8zV79dEwg4BiGSmN0zPu
lJ31pq+wb0IeMKkgdaZ/C/2X2NbA+bUX+KDl+2cyg1yigBj4gi5q4a29qoHqiiup
DKZPSFdPN3XAUzzpk0tAn0qupnKDN9Mmnm2Lb0Dnn5HJ6KGhcgEGmCjTAf9iG9Ox
VFWF+r4fpp9zTbHB5iuAss0/7op1ntpQaZBOIDRx0sxin/03N+SaRkV/0N+TzbNb
HTeYmj19TcNA8u2A1u/MHicCT+CgVBlfq7L7pAaj4yOCIAQnz0FGdKFW6eGO/Mip
c3KtV3HI24XrzqeQjxN65QRgfyZ5pzoixgqeYi8Iwyw2Lp37MTzIo+03dC9vDcf+
ayaywXMbUcywVWrQ2h03WFSk5Oo3BxwmVaJK9RyVbiGQeSNZnrODNSQ3Ax8oe+EH
TcmLQgwmYhR/C+2l4/NMU8bWNt8HZugMJOm7jq2P7fPu63Wl5nK+nJ1cvWCqc/O1
8NI+GemfLqZZUHixfcH+HizESvBS6fLjMK/b2TvPzslEA5wR9bBOXsJHD1IYNy05
S1XucAA1KnC2KX8sjvkU3bzZDUKaECuQCZ7eIRerJ5rUoAYf4B2LmF/BebBmNXIZ
34YAoJRW7yshjbRo2noGcnlUrlyOppT3P+bXtF4OY7RH0Qjp3gLDtn+xNWG8YRbY
04Snzkr/lHrPjFMK3hnO6hyVzLbGD2+K5GjQFJuq2y5gGM5jK+MkSvA02ClQbUTO
wxR3SJY3m09Mwb/r1zjS8mlLUD+Lj1cSEVXTTffve2C1Ksj/p+JmGPeqoqIRqVRU
VbxRBtBYWO8mklUuOWD2Z6CvWoPG99apbmnLpMQLPvMXsQ5YKKQzjyPBoMNb7OKt
VZkS1a8TpCnoe59EJf0+6MRptvXNrfE8oAjzZn8gaHBM16kwlcnly9JpLj68JkR1
jkijYQ/aTYFUUaauOTySky2NaxxZqntdgiBkJ7rna0HAYZfQu7SVgWmL3epBYfak
OTPAgs4BES9VFBY2WiuiEUSnRNBsbNT5UEwfcx3OHqZaN5kSB198NFV9tl0Zsww7
ufJkhNYr1gE0ieyJSVjsMqHMyD/U+26pnyJndwQrQBGGOtbKVf2csAC09VVCThP6
WSDktB906oSfWxegf2GvOfpmFSQkGbg/U+8MWqaulQEHPWro0c9uiqYUyy6vv6tB
3wAoxubmN2hOrYOGNC6nwPHfUJRn/mcv7IIHYNqgWViaxceh8vsRpW4XuMOlcUVC
njwbLl4ou0l3ygHzln5f+FLABjDfF2OPG3kGCKBPDy92bvjv6k3IdygXH57x+wS+
4uB+gJSGqCKsVbeLpqhQYm5B4BUUTr6xoHDla/Iqe0x/8VX+2aWAMyR7JkA8Sqov
T28t8ULOYz8W2opBAQLEp4pUtdt0pG+1pRzgev1H4XyAW44xO55WkwYXF10Tauwk
7sK/KXlZeIw2jAVDKDcT64DO4VW41IKoPskBrLmHEUX8urrejFi2tT6UEGgjhUIj
IXhQfR4IT2Y8cj4SG/rjsos9KJNTihgpgqkKVBH5TLeaLZqcS2Jte1abUBub8dDy
3SOO9WgxKFddk6dYYvK1PUsLQycl5xkmiqzclZQkpkoge76IlasYjJyvoKJBu1Yx
lhAqhffjR0/xEM5UxgEJlRasuDXy3apLYBX5mU2VWsAd2ZKfbuERQZphqqP7Njsi
jMytPg2tqLtZz6xataBaoVim4yUj59nip4uApkXHCGQ5G4apiffGzgD45l8RufGb
NPbjDlg7VfVB7eXmm4a6qfDiqOM5YbhcNtm65ddAcVU/RNeaRYbPe4d8PNJn9y9v
00cYfYiIu9y/WqX4bhvNsCWFVIugFDmFS/IqEBxIl3a0ZLveCIo82udbiRZ1gfIt
1iAdVfpAWmEVhtmWg8xvqnqv7ZjvmygDK4u+ZUII2nfrduWsYTYzilyvPvGsdDax
5ONypNX0MQxLA4kDVrltliCUxulIvP5q98la32SEOmtS8JZYfM2TfjJ5wMGk/ZaV
EhstI1CdMAx1dkz6dqYVZx847y4o60Mwxu8Yvo+dk32Qy+kHldl6m2v4bpeT2TCr
RrPkehGKjfRYyoB+VM8040iQOxclpYkBvplNSDyVCD5UixbIL6Oqrw7lAp4RZz1a
wMGJ8j3CxsXh/MGfsggySn4CQU7TDM9aLMmJyzZBdgb/KekRzZ5QNZWFa1rC4avo
T+aPDNCXYAPIl6gN6fXLt0Mn9rHyshgr5U1uVdJC09qpy3nZRZnf3ZmfwpL4xEky
aLr9vUUJCdrb2t7D7v2wLZ+sAIBxiOYs/evn7GjqHoW1U7MW7OXjofg5GDA3jsW/
bzbs+GB1TOjaE0Z2Kudg1MX7cNQnRPPEqTrp+nQNt8OQ79z96V/pnWVuHbF9drqc
Q2+e7M0eL66KGADvHjeEuaBlZq1Htnyp6huSrsbEz+/8zPQqe1p0T8mRoJz7YU2Y
boxA7H1UbHawM70OSB+EguwCOyMIMCrrdW85gBOH90wFb6vOc79qhifT3X4tFVT4
Ghmlz7cbdsOE7RL8NE8XbiKSV8FkmmksdvX6i2aPrqTassx3Thh4O6AoGB1bzOiW
NRi3oOUAlO1+sViZZ6G2Zbu2Dbdajqqqx95lJiVoQ+9f8wy6OpYnQNB5sbvBebRd
oz3nzruKsc1Vcq/kvKHaf/GwignSwv33Lye7VXYDvpKxjlJ3p9BN1bSJfI2m+dgo
Wy0+492ySgzIB5ydtRX3IvxJ6s9vLt4SiqaifNjhCzRMpjSSvrAdcObauoLzmsLu
/Tgq769G/ndd0I1U7A++eWI/G0OxmuCAS2yOfSHeueR7OqHbR/ZQ+dC5Op2XKhU1
u2o+urtDZcUbVnFtpSPScCjtxzLzwnc441eiOujJH2ocXjzqtYgcs6H6j6rv+sGw
9985yvqoOn8rzGMPb0/wnCAynuKvBOOljS6UAG48uFzmImfA+AOH7cUBqzRlxdLH
aKQ4uJtQdL7/4CZhHVrWh12xZy5aLbZpgCiLZy3AIB1E4mEAg6laJKurJqmNX90j
E/hOGwKSobIT/4H6w7Sk1KyaCEtxPs3JXxg5ICZ+qwHkJFGqzG0O9vfMOhdWulcb
4cKqlusXuJo+mkkeT48dGugGvXulCyMPygQaWhO4NAJpILP3poq53jtGmokN77jt
7gxTkVKWl7Hc0wSoPotiA0MvZiodc1wRmlKzjW87lhlO6T0MUdtCjQGC2aFVIveS
q5BFY3iV5rupHKy03UrL/WalGshv8orGTvLaJnQ0tbSpoEqWOW6Pz43uuLOh6BpE
wqiVSkJuKQdIj4dAVhhO3daAhTpNukhq7peLMyqNNW0zh61WEDnwGcJ7DK3xdbKG
OzMzMMNBRSAfPoQnlpbiqbtJIg5eAGi8jguVGOty9WLj5e6NpQyaJrt15ChMVd6l
ZKWflfEQgRjoxso0rTt3XF/OzTGK7ZUyWuxqvU312DRmtIfJ/iN8vx35BbalmoDq
o9ihp5mAjaAzKHShTHXJm9ap7LIo3AfVtD26eWB6vJ2eaA9QhyBDSYutlBjhNeBn
Y3N3+UBScXBM1EEw94irzPl/yybDL72/q/kQEvBLdxs3SYAWorZE9vBhqnHimZxC
4wyYRWHiiUb3zk3GcFlvh+FwiQhkS7Ek2l5N3eqcUqIp/W8Ico1qtr8IPgNI8zqR
cTx+txxPFMQyrsLFNKtg6fGZqbhhPtu4OcrH630JntCKo9DfGIvV4DHZxa8Vpf+H
XSQFnprEtiSa14g5gQBFKatDh7bNaRp0aodnoyIKuIbnQkUzHTsBZ6JxXOzSgBWI
HXTchylJdbja2Z+WaCuIZMrBvWk7HhULmjbFO6rvB2Pl0wF2a9i0zqVQWr7aEMRu
+72dufSviC2dfRsfjdjyXvJ4PUrnun3Bvtmnald02IqJk1Yc3Ibaim4b1MeEXU2L
s1uSCDXcOsQnejJ3mw4HKDF8lxoGNOg9xcVDiWlX/dfJxtQ5i4E0QGBwo4rzwezK
tjeDu9HLqDoQUj6RtY5Hw02rInRLX3Yg03/1r1DvaUSsITaU191XSllj5m+kxvUA
fiuX0+ix2kAU/2Im8VLjT0/yzAXxIa2tyih9rbcWU79wAuTOgIa7YrBxXRgO9Z6J
lcYQWFoO2RGMvJ5+OhUwxickdd28IJjLMmMYU+8JwkdJBfGOLV1bNJFyQIzwXrU4
2LCvbSDji6/rPQ66L1xmWSVTmc1r/OZ7oPKlaf5WOdSZWp9QLCW6TZ/1BXsHP0M4
4QQ+STejT0Uns4ThwPkCAAUVXPZP/G7X5xZ2pkc042bleMIzqtlTYzvI4J9wXz1T
W8U5rQnSJAlZI1wj5+3cUx82WMk0kSKecUjd7qenDmJsd467xNqRb67twBc+Y3n2
c8680BPfkdwQ2P/tYhVfLBsuGOFprdZFQ8G4KNTz8FVEKQwIWMrsjAwuncpfiBAe
9FiX9CknIJeVRe/1VvMjup62BIfN88sIgZWkPjLK8IlW2+sC3KzCWpl2pTciX385
iitPK/4dWylZu78VLhpcZXNVJWJv2FMow+qxXcurjdPCeKmsSbYzMJXOFlObrzjj
ryOzbgU7FoBjEqo0RUkOYHBb9DvDq5ILCqzhSBgay6sY3Oko005yCjj9bOwps5p+
bSTXsz24AWRUV971LeTv1TqLau43xiXgL7HYD6ZQLsbNqnKnIaeMwMuwhozYVbaJ
mkgbrHHkPhIqCx90UBEeBhug5IMWPKJFZp0fsYTbZT8E+IdG7L4JGkDGPdzFYaQq
2/vI3xIVHSgqvWAI6qnutxFL4anN+U0QLOrl4WGo7NfN/jdEadP7VAz/MfZwxNL9
kfM5u4i5EOhybvAsSPH/R/+eDlbDZsEzo5pgHYjUkUQhtjRHFHlmN8P1H+FhRmuZ
S1aY/3roGP6drCHnKqNDV5lnwnnnJRL42hAz/pYtvano0PVYpZP0C6P5yyyrqwmy
3l25D8xgKalkzIqQZuPlnVD+XkCmisC4byU7aPZ7Guzm7l9UlDZqY0ilwmd/49i+
urNIYKp62G8KWp9z48qZ8eo64pIIhlj6Aa5LVyRWkZ1ecCGFBm2nwT7Yvr1lCEdR
oN6Mkzycz+fovXM295jLsrGg0PL3EFMun86JM7kOWuQXqqCxywSh5nRdwGDXDnD0
qwQZwxzBYJ+OlxyL+2WDpyT66XHYEQ1mQh2MWFs4Lx5ZW5Q9QaBpUUz72fs2QmFW
i9pJl3XfdRJYijz/qk9Wzv8+L6OpDFs+8ncbTV+MWLxUqaAxWQn/pkZJFTYM9D37
6V94Fs3jkfaeq2QoTcgzpKIycjDBSggDyLyqcpqq12PaMtQ4FGqZpf3tvANvXyfd
qN+PRs6xexYp7jr1+mYGW63+Rmcl7ZSWr1C4ABEXd6F7qMPQ+QyDF6zqYKUOk1Im
AtFQD38+Mq6txWpLl9KY06/WEBGHCSqB7iUgejg2j1hMKB3gkIRCFOIa7YRT7tps
RM+l3mTAk28YkZf7rmJwHIzInE5slnygkc1/oXBcdesmuQ4YjgkTxnqtfgAaWmM1
OFQR3yS1dojOa9sJFBD8uIA8NkzvrNvYOQDXiVDGDqJ9Ta8oFW2M4mCo4UTi7nkg
MgdDFRKVcycZ0TDnuktdUc7p6ffk6+Vd2n1mhmXDLPGx6ohefxH+5PztpeeD7yft
AWMys+9rpIzcLIsf6673IJDa5KrGv5Gbbw0g0v89nKfVjcMsdh0lQXgl43GAzb96
Y6ApB71iO6CMWV8LRSblJr3EIiUgD38cWS3fRqXP93Wt49q3yj38cfvYXWuTYfHX
9yE46CKi0WUCs3TpkBrPrh2QTEZ99n4rZtJgRqcdfdwk32QgAbSP2gEj1XMkbCyy
rl2SIXz/JLhwuKXQnDx9xURDl/zYNdBjJDPXpJELxX9eUi0tGglMI4GPJWx/zajN
WRBCIYfAOyLPFn+vWbrIKF7oYKl7a0h/sJ1JD9OPd62pFuiRQ9Y6DicZkB9FQyoH
eJYqeWV6YLYuklaSXi1+8og0ubqOfE8w7ZemJ2Iv9rfIrNBKANIs4bNoudRa6gxG
tC/ogd7bhSp/Ouu6/SDNljhmfYLS7UiJnvHP4AW1pF2ox/BrmsU1vUP6yccuO5Mp
pWKUzq6hlXDrfrVvj3/qdU0fhhskSDmI+rEUXrGCq0oIoIrG19wSbtuZHbeLOetd
7gZz1VyO5RaSsR1lP4IXHv2i3N/x+CFBn87tLGB8uppO/oC+T/hLa74Q0tFaaxJ0
HRDMW5JE31sv/dlnwcvr4+NaXWlgUbJksPe54xH8Tym6SZrw31Y8imKMVnWKFecu
oz9d5ThCr2ne/zHzbJ1XMvm8UQkkjOMP4pEFYOJ7w1/bZ1IyoAYy+WJi7Ny+8l4x
mdJWcA/UCxPJXobCnI8Tot+CGUFuSK3mMkvcC8447nx9O1WDjVFH4iOqxETezNOt
skKNBxMN6oWqekIZ8kx35FNonbhzuuO1ykt09/cbPbWhmF99On6niqC09BIAr8dL
Cqb2pw5F8z3nXDcqVTFFm5PegERiQEgbURtiqtsr43QF0j45akuIIMZmEzWqhLGW
57sED5vqeTqTbsPBfbJwtNiL6lLg03HMzBnWVHUDaiaodkc3pZmw3TLyPSxV1VK4
U5GFRqmtCNQkwy/kt+uV4HNYZ7P5yo91I6tw2hGmEWixFHouBoGObOntheQJ5PmF
Mi4pvTYGO26XIEAOya+/GIzDxU5XTTApiaZ5tR+n139QMNKhsvfYLGH/L5dnNWtB
5o6HI3JKUtJKWGFir9aWP/Nxl/pWDdmYEle2ldMbZ0HhLmmGxNJuDCv5/eQakLBl
fM5CdF/o9jcI8oyY8W088b46Rehu703dTDd4D1wNY8uEtHl910qzN135dbUy/wBl
cSrgbhAjE2PrlT561nbehUpVWzgb1kEKbpIdUlUzFWe5GM+TeiSj7IT8G2v9/z0w
pKC3tIp3tCRcosiA+NvivK3yKhXGlO6PKnZK5WN7ALgjTKE7bwdt6Teg7w0xKyoO
70qlUTNTAS7wdsMWvTscdGD6M7UDwzgCSoQSkMTmpT3EU2wCBLUxdgugo8Tl1ieJ
8+HuR1oN4Pd2lolyDkT34l7sLE81swrTyBNhogMKKcPNOKTAkUHdqIU3rZxrhQ8v
mfIzzfmbWwl0FUtApSmvtnAoI5l5BGlGZM85103VcBteqKuEQE0NHf7gqHndWprN
1xcx7FfLQ8pgeBnGt8xQM+iXXBdJkEXEfdLjWAbWiv+l3aIKBzTTulsTfgPHNhmP
COaADUHi2uxnVEcQWQ7nyWOqFpmIYFMJMyPqal7L2FEutyOvP/oh2C1Di2AMmjg/
sHDnihVqsTgAWa5DN8HJdmMI2GQ6ofEgdoF8CiIY+nfxJCXGVr4K43s44YlUe4v5
PPthMGNFnST6l/PDRku3Il4TlMshvpeuiZ4MQ2zWIH0ntvA28Y8e39J+2ZQWoMqf
YsuWiXgytL65oJKEHzp44DDYznyaSFBFY42AdV8X7lAHo3eS1c55dydZMhiXFXlU
96AlkvPttTaO3RDRH74DNkMNBORXouGOr6J6SR/B82YYeli6Z2XKU/j3mbtLKLG3
dU0swdQc44q+o55jDA8a30OT689YLj9KpxRxEfRHEnkJk7LfcaP9JZMmPeWXDGMA
omfWOCsDCj/Bk/uEBQZS7Qo+CBVgSQu+0WIWZYBu/AKasHOeQLxm6LpANeSvPxE/
9lh5m24J155oE6YNoTEwQY9nduhOtiYUXlX10GDteXPpQBokNT2OgCY7HW0Ujfwx
1VtChK5x+obo8vWGw3zbRkHy9e6Kd169yHXZ1Hv9qfZAeQyqxjgK7nEqHmPoMM2h
qZVJTLI/Ma9Lra2o81NAb7d2TiRAQJpQdxmYa2zsHn8K/tGcMcDQOTl/6sfU+9tX
Hys11wwWcB4PghmQBqd3/k3cJwC1CVi1Hmr9j05yjlW57bsKwyBY4opTZostpEOM
xMFEQFDKbv3dQW9dJlwR8htT9a8plJtJY+iIGryAWWWYaFMgp5DR4iSI46Cie8eW
ID8gfAv9X5FryoV6t7IuYRx9G2i5bRnA9NUxJ2Q6RjcQhljX4z8D7S56XV9671kn
400ZBHjr6ovRlwX0qaP5tVStK9ehf5q5SX0QRALFpn9uIIK1czT7N16iZnRr6UGv
RHhZ+HgokBTKS9sThYLyoGZlGN77hJrigIGBukwDIV0Knioa1rV0HuYoyF2oLm38
VApzsvjDUcwUTz8mUDZBM1/a2Hqx9rdTUUONctyYynjIznxwwYa9uCGKcCYuz6wp
9AZ+iJoQdZoSu4Y5nGF19ofwJ0aZ5DVif1C2Y/xPBcVpJq2P73uL+dI1J3nLTTaS
vQ8s+wE0csq0j+3HhFPD77Yf2vcYoDtY4uQjytg1s+Yy3gi0zZPUm0uiMt56hR2h
O+ip5/kZOuekNDjGNhTPHnh6ArpqGqMpuan8jxz+kM/m7WjSOywsq6p8TWpqkgse
ZlG50/d4VSWKSz+4z0lqRR6QhPNgt6pOWlStFYjouKLJ4/KQhaeBvLQDoGRkEHP8
SduRzBd4MVLsFiHnhr9CAc7lDcd3FrkjjtRJGMOFJrH5y1VgfS74e7mt/+LNq8Dm
U9knDa/HVtKmx3PqRKLvWFzStZTYVI8rLO95EhuNaAvHJLbH60ys//1mYJKKRl2G
fixzuZtbfxD/kwKZQIYW5g3l9AHty6ksCB9zTW4eY0S7GJt2g7s94Esn43RjlGkP
t1jtrmZGcsy1LP5mChxzLulQynuKT+kzvNQL+VFikl+hW01Fx6PABqR/IeBwhx7F
t06Q/dbVCFIzE5jx2A1S3fG8s+cjvwhVi+RPqJ/jQVxjq882ecBv9F7BCXt5n4zx
P4VnRyJNJHasP/ZGOtXfYVuCrNBZXLHvbI7lmQabp/VbUdcPX6M9wbqBe/8Hmt+W
IPS+/z0399jS+nFszgm1IrqVvcvKtFTe+2fjWVq2BxI2mByhZjohho/uQ6+9Fv12
Yvm3EYZc2dfGU999TJO9OG1JQ7G88q9XdD7wnluDRVQy7M9x5KNaxdsBmLdow6F4
9KZcJScQ1oNk3AQ/Eo6Zi8PgxCfEatQRxggugbv8egkBeHJQga/wzO9VnRWWcZTE
muu5S3eV0HRZZBBGhdYZUS1tiGJZmthpoqZw75/kezXBtZgNU4ekGDrFKwonFxAk
WBvRePTTozqcKiRllPcWf+7YKC4WI0wBFRBVBNhK97IYT4XDPdF3yJ38+xRxlGCC
VZ6wNGLdJ7zKadKr70yCW4Wd6Zo3AopHlPTAB69usz25zMxuYIdul+FlGQmlErPy
2fvhVB6BGUTvLVIaH/Of2npPVLrqBYehsmlJyyDy5pHMXLi2LRj/yliFzQFjNrDv
Goq8kfHRuejIwvysImtCIZUiIPImTbarPYcgSlrB08vG6q+P3rgWZ22VzO9rQ5tT
fUXeB8f8sz4TrH7Pi9+9oKiHGdrHYNUQOm7Ij1OxlInY9AlddJJj0aWSU08W0vPR
MaTuv4WvH8obWChEbnQhk8ZUdrYpsZaYX4fmiNtPIvVx4HiGLOQbdWbUm7yV0kdk
zesClrfOgQfRTLuuAQACCPnPZ2M1Pww5L9oCmDCjGyLMIaIDuMsrRGqcguc3xuqV
C+w9vLBol6z741WoMmiag3RZcll3CpA3U1B6bAagiXIf8HTFNO1mx9x1zC2a8tHA
NfPSA3nrI77fnLfjrBA2Rpr1Yb8N4BEWq0TWhDU0G+JwFU83w+gjF9qtP8aPLqTo
+x2BhDwuKp8XBnVR9VOig4EFhct4ilS0jJKBh7/cFC5LMpIXMZZ8czDc/6ZBj25t
+4u8NQbmURlGQlEAQT7xBvk5qespwNYg9mjNDXPx8sFhuMJYfr/hLOf9bVYiJFUd
1NQarhGpZjV5z1aeOH/HWHg+ymHGdtieU3HXDkWGOa0yPkPLkXZ6+vOp4Z8rHAa0
5swNgmu83xvNNDI+cFX02OYVEBUjJKMZ5nCGgkLFT4Kn6Jzr05JNj+GHcihLyo4U
D3BSuhkJOUiq2L3KADP0xSw5DaG2IxPoQCdLpL+5hSLOAreP1XIgRudVj8MLk006
f3Q/ubqThmAkmVEDkZi84qwmQFVpLGZt0UVaY5q6AnyFMiCMfV2TdDwtkSocMb0Z
fXVuTJIREomXNygTfjOphEmYXWeGOPqfOmVRg3+W76qCM+k5JZJHDqfVRfDexH86
Rw66YFXvAKt1WFmrLGUHhh1EInfClCVVNKmSvXVMK/MHJ2xi+YJ4RF4atPOgKBIJ
3qbQo6qwFsnQxGOnS4X8jXhj7yfLvwDXhwBd0HJQAA7vcyvyRewM/y+ppCEDtLUe
WotAy3Xtwk9rZbzRR+u9HaJ9dI8tt8J2AbPz9GbCdfNDsM9SJa9qvxp+Xbw3gQBF
PyhcwxDYXx4nTP+TVWkaq4b566/M/jiuXaaFPQWQMAr7JQ4EZr9qwe+n2PYX8N9m
dMrkpyoHPPh8bvq4PsNhjCZ8RKMPg3gztuz1M6e4XtDZcTT7miQQ6bPFjLq4o3Fk
r3I402wiV0JBLbHWMSy3WiROcNy/DxX/KQenaQarXxbhePin3clC4sCzDnP7RgY3
I5otAnzkJuJ4PGrgYmWAaI4ldPAtRhmQgoigBgXNPabu9/aebEJipIZBPUCQD88D
PlxRoq0gaVJ98EjhwR/drkMO471rzK2+ut7Is0moHJ7+Yf30MllVFubs1qfeVIAw
8HBnRdBRbI7c8SinSdWFjyAH3Doh2FQMPY+VaquCfVH7ukZg1bCtHo7g0MU/RiEd
8ZAd13HlV9HQvlDDBIbgHvQwid4ZbmlNBA96V30oC+pKq6SePnyCCGqdMrTrapbm
ZeRfJwgEHY57NN/zmn6f0IqvoznqerYKVXVsXaV9ZETGX9PcgTiHvafCsIrZFg0t
TbUI7ANamsS5CI7/UGsyzfrY792a7Zw43Ayo+GrAag87dK7Lz9ykDamGdBA26qDM
QsQLT/UIHSYwG1I02CPZJsq5dWYUJrHLueJWYYXkwkLdWS1nsCYJPrKy1CnCQSca
NI8GFBEqgfxJBVmqaiKvxKNvnSr7novzNy+0BFOqqif4CGi3R/wAQetb13YP/sqb
jG7yiy+yNhdXPERpYVpi75icZqNaGS1cVGMh3uYne2oNBVrLtb5dwZrcPaatyfl3
kTallc8bU/sYrQvhPmvo44Ze+yjxYFGciekWw1Eq4c4AacYZmG//CLzo0XFJCkjT
BMgEDeGYBL4k8QsVBNFSeFf3rPlK/P/5Aohh+7uoDd5WNYaX1Wy3Rwg8HngkfQj5
s8adLIjWoaLXA9UN0rog8b0irLdO82P4IW8SM6Ov9Alh6FheDc2Dz+1zwui/W0xT
0rE0QRX/ehEDdfVP30ps7gskNCiKOuGR5xq2EpqLoyWWS8/I/AsSZHiGynzsMmnJ
1XVsENfNexM0mvS+pfku6UN1Nq5/Xu7RzAlcye0gxcyQKpQ+b4A0bPHVBl7WXPNN
t3o5slKR9Inlyu6kWBZ95YGqgudW+JLifnUGdr+0D03wkEfW5pGqtpbA/JRbPaqu
6lCUPL1lAbf0P+VrWxSM/oVxsK+/EgvvxRvEahGv9dQqZxEOr/l9U0kTAyHjJxw+
y0ruPj6wz/7lRDx2CwOh4cAQT/8uOKEVDe8qn1IsYtn2ihLi2mHuLMOzVzxi+vA2
iASzdVJfFPrcu/1iaxjrtzjfVJnd/P4DgPD6TALZaI0W+kfgnyJZmAwJgt6w19VV
07RQBS6kQId8fVUzLLX1Gi9LGnaM31nfCoGMmnx6oqY2sGc6dP8ovpobBDSrjkuG
7zyXwjHi8pvmolHY73/ZtOx9CDytXHDMw/gwsEm1c4o3vMbJR1/2E4ZZMxUAOpYh
JC6I2KgtEQZADH9nWEDWpJhqvZkwwtDREiMe7pXamdkf1/OTq+ak8msr6ztP0JCD
8SlYPn90qwoT5Ja5NfuQL/nMHBGhcEb29XZoX9tTvJUsDidc9KFeVhGwwnnaaw6+
tfz+VQulWta0vnOSCmNbBmK6SQ7uppw9+vMBWZwfuwl2bNr30dcQWBEmdLpcrMhq
2k5amJmc1bahgoaTlvfMXkpBLLM8SKZ5lUQJ5hiW5qOzP3yQAeIuFtNtjlXlMMLL
C8dvJcLImLRgM8z5CbT6BI5oDhfGF/YHfBAsmA4xZHHXS5/FvHkQOL6eTYhXNCcx
VqCZRJn6I1WQqopuhV4OocjlnXyLsSO5PbiYv58nfpo8rXrVb5oR3qkcM5/+GcCQ
qqkByIDOi8vyW3sHqXGnU55iYy3nY9CbRQxdU+OmjCJbOkFo/6WibaANWIHnrr+l
7318TvpPHgidrf/Sio2Os+k2VO2I52HLIIyKU3Ck55pAE06/jK6ai3cHKasKChDi
Y5e63AwoQ9N5fHl2hAVO7us1k38gIEIOebbA6Z9Tdp5qYgNWnJuc6vj2ilbYEG79
n7Re5k1/zahr9PUfgjLaVHsapFDaSeypJFYc6n8ZSM72R6aYXkLlNp+Ze1tFoYqv
OkyiTYSjhKkcJ2AAoPVmnrwNGmSwnhYwdB3PrI/2RLYjADNFGDVnLXMEjx0NDwUV
bN6rLq+ffAXRzbNOXWmIy3o4umDqeZfg2UnjZISwwItbmptR7vMW43iMhZNFTo2W
zuMxlm9z57Y3CXkKNQ3hLfBcHCPKtBQw9lcGXitZwjeWbq8CvJCQHZnX8t1vmNN+
UYRRdp3JO8tBF1W1lwMVqSdwT6d5WUQlFEEXX9CrRNZ2tSv6i5D+pTpV8lw9oudb
1G9a/a0SbLTCeNYR1rZEu3s+gNATjMEZEC4OeKBq2D9WfGl0O3JW6ogkaEWK1wrm
taubPhviAvCzEVLFMZErrAML/68nSbznK1wbjzifkkmBDYojTz4vv0Xf14g7ejZ8
qhmplMxbQWCzqo54SiT6Et/JytSR3hBxmeCDclFHgTFzvrHP+/una3WEd1uCSq0z
Qt16ImRHyB/FN/vtz4W3J58ZxyNzIW8+ElS1z1bJXDXF3cywxm2fMD7xd3ZVNzpN
wzrBsyUOT7q5ZzQ+zhV0rc938KpRQWSq4LnDKMcdMPXXMFFA4+bs1GzoZCHy/AJr
Poa/mOsL+dA+C+FYrg6A7I9WZFN/PhKpbmQzRUDROHuqi1YnbXdo14VazJtBs5fm
aVMunODNxYf6/5Pp9NkzxgUixERrPspA6R0eflccYAUcXHe7K41tEq4I/1W+Br4p
2qEiT8Ql1MpoM2DVLECYeYEPred2YnWFocSihkVbI41tN0l/Sh7hifXS+anP8lY+
qEPUAqLrLlHRRsPWtX1qJGYcyG3ENB1jp0mK0kBu2gp7BbbQamviYYqGc9NMsUnB
aU7yAu6YPTSwdh24bEmuspKbH0Rf9Iq0alLmYD6pHfNrcFQGRiUSXM6isVMkYBy4
LLjwxPx4oUQMoLgY+QH5bf1Zej1m7bNv9ZKGYqFQ1AOvhwnrWm1x37ngVtqzc07I
oGjMQC8X/IXCPcVgmX6t0Na2xtNKb8DnsX1bFCfiGo2ZYqfgVYjwL4k5CZaxbEA6
GLPKkCpT+1VzZvwCe1G2EKXnocmoJzZ9PnwbeSKMlouR5JMoBNFYjiVZx1AilKWC
3MT/dAbiUtgrbU7FF5aufGYd8ogSzMs5nb9pd2tCxaI7F+TWPErbq9nuBuiODREN
kGxhadVKlV4y2U4lPLC1KcT3omrItuRJ+HawrpTtXoHmXQDvbiPTrftagogZ9ucX
5LxhJHyWspsY2bg7HZIjekgZH2LItt/5+yJSaDo0aNJ6bHhAAogGPcTJwTOZ1fdZ
Qq3LSvMCcWbNhXgAItbqkmK2UPlcSl5lJtbVt3igpGFtzFRlnvKxO7eR0vZWfAjO
Ilr5bvDtM3zq7omIeHVlqLVm3HhSITSNuhBqiJap8BMUZAwRVJTFWttwEfR1ut+3
YRWdUZuKb6558EIhCxJftWmghydWBu1J/MXkY0hq0PalQsUoTDGXa5a3IMY8Qk3F
MxZp+vwME+tqoYFAiiJtDVgAEqUmLAcQXPHCzsdI75r3KBY7WBz3i04NkPOx99yL
iKwf8clQmdoqUy9y6NmnMUPzfagmMApx7tdmWK+7zT5Vjc9EdCEbNDkQsSBXLIxa
MaOa/Qbw2Har+CEqxp+X8wQIoSSnFs/lSrGFPkOViqumm7FM4MzpJHN02xSbrkE2
Yrb18cN5fhllqwV8eUExcalJhZc7Y7DT69m/t1JiO66PLmBh9Pi/nybgefxNqDWA
xVImGx4ae2ZzOXCJJA8TYnU8hf6w4S9ulYk2tisN/Rkfm02g8y2D+9S1HQIaLqqN
LZ8jP2I6fhZTFJPpGb1vt/qp0hP2tQUzWYhnj9KoA1d/RPrBWzH/RbZUEai+JOpo
RP14TSJ+e6x6w19aZdH01SzfzfJ5X9lJq6TRbVBbO85qoZgVFy6w7PxEoGvbEO3I
Zb07CZmBBIRsKMi5+o4oWANBPjAzYiiv5Eepl74F2Zos+Dff3JHi3aPCH//jI6JG
cgN0QE3xuyUFEeJK8TSUO8wGK6x61dY0MfP1xaHCvOjMPKiZS+DhsKw+bdSNsz5u
I0gvfci2kly4AyFzlFMp34gsoMJR5drEpQM4QBsd7HgmbRzDWV8TD9LVK3kDYSKh
TOolLv9Co/yT1TYUTDyATYsdfOwN9pzlEURuhGQMIKNxizejkl/qsYb2tqUo9TUC
XflKKdUEzuVdkN1YeJ47UfRhi7uvcZLODfemuquurczk9gCOZKjoDK0BsvbYdo1c
y2KkoxXgWULTzg2q0ibG7qrNT8HEfHrIGl3uNDkmnRNfbHSNU0BBCISl9rntftQh
bAgkK6r0JkPv8xegOOkS6I9GaDsSTI5KDipTKca7sUiX67A4J8yecXPa+DYkpzJU
r33knl/6JLiuFBRJVswHAbTiM5fW7GvByaZaULCxxAmw6UZymr1oAXsT7gI1dkNO
2gOav+W6DdcIElG29rauI2vDfblICfF3jE/zyheIBg5mqwi4kB0ZjmsxlMh9Psu4
dChGXvRdogwHLtLWCX6pWRSowNn77QzfnnfR5A38I9GSIANzT8co0pRsC1PVFWcy
S+w3GReSemBc4z1XZ6vADw/Xkw49XkwRmTRzj7CWRC3aKwSRYd0D8q4T6AaOzx6b
eAoyJ0+g/NCAeD/7sIQGvy1BbHsuI1+BZNOky+AqiO7KpUQvdJx4fNAlYE2Nx+n2
5Sm8zHJS5oNzsf5LhAPreG1BjO3LINNy3GWMJPlzeBd+Z4rFTsXv6hgnaauVzots
DtL9PbzR3YHQVzCSx5FrrbahcNM2+Mp4XVbXgHbJUD1vkzFJ3gRuMfA0c1/XoXDg
ofuZn+Y/JDimsPyLeufoip1k+DTklAUArYhqmNwKugsxGopXNgUM1YUo7/RBdV9V
iWrnxTs3VmaUbAkZwFHDVePS51cUQaZpo82icOtu4vcaKgwMYGZlDzIcD6i8QQR6
naElFkRP7xSTlwJSSsjtPFTIvkCyRkZ+FTrSfJ7GUsPvu/vwqYUmKF+4KH0Dogg8
P+b/gTW1bEI6bWNydNeX4Ms/MrafFT/N1dAVq3ujw64Uki9FIUEbTOHZB5Do8iYe
+GYV2La0xGp3wdYNlIMqKHNTV/xPbMwV/pzQEi9SsTh+/TB1mZtopChP4COi+TBN
YooShXvgHyWdmkZUPLQcw/HMMOk6PDreAZBakKwK/uHMIktVxkUmHjA9vG7Fyo9t
jW/iHRBryeOYRFcclmUxDGuG8EUZfY4EGPkpZZpvtbGOaEvb2jJxm/QTlSOzP4j2
SynIsOGyEoGfZTm1XvhNFykdMeck8bSchQkF/rcdW7BIuwHBvvjOX/zL3NcqABeN
ut/+I+n9SOCiMkodndOagy7cGcOf8Qeye1oau5uBhLJQxhjHAuRXWtPgnxyTact6
Mi5Dd4u64QXjXDuizkcSN5JRUFAlDF63TYBDIWa8HfntBr0fBi8AVpI9PdhHhR3+
qQn985D1FRu9VFi7yX5iH51dtaTL0aSkZ8tODwK7wt3Xbd4+Uzdim+mZqjCVUYuA
XvKm1ctuKnRGr1Ug4EoIePzhLax0qpMU3qFoOmgHGfL9yWFkJHE+ginkEync3RYI
tnXYYXJgTNsFt58NUylVk6yDjjCLiypRsEKrQZAd/lVI7BxuDwsHpnPeQI7HKXO3
mDJpZwt78HNgsr9m/Qq/5egF5xFK5Z8SLs1uhja9rXF7wRbuDMPHVWwvTBLftVYG
3wkbwvQEkGgHg0gwAgGq6auic1NKJbzIvYAi3jFDI6ob7WS5rkmGU6IgoRHQnAb7
3ElZSogCwktljr3JpW5/LBGOpha2Xlb8I5M3zVVSAHKpsYsjRj0evcxtgFjXyD3+
zpdtyMZYkeqRt9pKHVpz4ZdAm7wmtyytDW1UVPDSjAUJSBRNTcW9BlxTrTw9tgmD
v8tiRs3m8QY05vZQ6NaOZJIcRfBF5HPVGlWU2PdmhPMnvfo/6HLSp7SlsIycDJav
HN+jEJrRjaU136RTjtSEpKH3yRPkeDxsiE/MzHlSmLeR4zmXZDUDwTPxfxqGDjm4
nS8A4VCYnU7lPjLwIaLI5zFpurmM8/61WaPaL4VBbnnZV9WhFbeRRTcm2EjHV/mQ
13+x0FxrYjCLlX8LqYOWflMIEJwhFQnWVVqU0mfME1X0Oh9xmNGKi0Pd2v/vRyGY
T5UjCUa6PRbuyv+ck4Vfz9cWJpTwebtBhVpYWqp5Y8NuPTzYAZDnHDeBBOsdv1uk
EqKZltZ8Y6LbJKo9upEkNQHzB0PkyRSbK82F648rWCeRQz6OY9/u+UK+xpRlV/ER
vwKlixtAtyc9PFT0MmSxUqE446JwfDq8exI8GRIOX7PKmwf5eJPsYOR52DY0x3Is
frKErd1fN2HrnmAySFV3GKtOmks/ya5TMLmrV1WHVl/7bMRrQwy2d/Bwa2rYWXVO
hmee5o6JqhTKpnFF+gaYTLwwLNNedlmTFLSLJ2/DUqfLDl8q9vrZZejbvBGv/F0C
fq8RVM2JNrKX1bAWlJjBvhJkVhh/mjYZNOxq3Hceepo0QLXk5olJbwAJJfBSIi23
fDs67SDdZOQNQ86f7Y9gOFqKKVhPkFm0RoEN8jJlnye0EFjo2hSQN1W8bLjszeqo
kYeu6ORNEq//la6rpq+ox3eZ5DNFthGIwTogiE/6CorhuaJLGFss2xgSCkRVPt5p
fBI0fRrSnk+bC+b2CRztlAwHJf92kTP7X0byn3E9pXJ10V3PUwZjWaK6+SZUhrq5
azZ7KDtbhYHrgAEOvCD5LuUnEWYIRSQ7EKYTyTRiq+N9gPNTjlgQfgYTMlXPAHRk
iwHyZfEJ+gO3ZSu94diJyKfMlVXvHDomlRa1C25bpbsA87wbyw5tthaCnOKD8Z9b
66JU8tDB/QeXHYYvovpLVB1cTpHQTYRoZ/mfS/4VjfK7/If3vm9Gym5CDfxEt9oQ
GqrhHTwqzA1uLxiHPDGnc4XbFAxujL0p63f8BdkSuFkh2g7kPzacO+bHJW6Ttc/t
ncgGEpgWR44r8r/NccdonxBGRu7FfxtNR/XK/2t5Lb/jcA0A1z/phg3+yp5GaYXb
RzZreTOeFM3DfB3T7obfHM7zSv7ZuHM5lIhznsOnX9LiRmMSk6riV6PljIxwKPbN
fPQDv9WV6dpJJqvHZuNf7E1MsAWuPwmKQlwoaypYrm2+mFWqcPqxitN3Fu070xRo
2SoOrhlVUCsBp6KgIo+mevTwzAwFFpJ8ukUgPIPdFux4eJ1kNfmqjl7G1T4aQUX/
CwgwL6eSI2L2iLgSlhccSDvQCEYXaFbDFkII6ujoqq4ye4DgZYZIThZIjpDuE1lv
QdZ0DdHEdGW+eIF9egXgWh/ld6I1ITNI2ywwrIbUaKrOcTcsZ5t81sY2pi6ycOAX
FaiicF1hJktbPq57Yb/fBskUg6P87hpX047O90VKoZD1HQrucZbktyft62Z+fih0
lcHaqwCT047ZyA49OvAMGXzbHo04GntB6x6mdiIPLvwvI9YwW0KnQimI/5XmCzY0
tIkPRZhjAElt6xCwUN4fBelkU4dNSBimT5as3YfMClcgWhvHc7fQlcN9wjEy94Wi
oIujIAoGpmA4GtKU8BRg7Ow7KwOejrPFZNUsCoaPtphHPGhpvJJGM0aJ2e17L2AW
zypt5jxMo5xidku3n9Rz64aMumu7x4ASJB2WbMcgKYmpKrvzBDZpxMDRbRw2b+zh
4QvF/i2wfphTzRoVS+GIN71sUUGrXebdPljHsin3Y6C86exxKrrun3I6F/Gzlm6i
9Fk3jtOlhUtjODosvmKEkVVuu6ZH841DJ70AlbwWBl7OMCnwCYga5q51+KoMKYiv
bmJrnZ99zUxnQ8+VE8/1g+5wAytRoew87sl5Hse4w9gNyjFQ58EIZh5ma+u4g5et
yPNhT8G21EjMbvJpPOSNRAo6OJ9TZGA5rU5sXIQdI15TZMXkPHiVYxjyr+YskG8C
PRA0BkbAQNqZvc/7oa4hMQlWEZmGZdqaNuxrHr1rGm04OAgxgd/+lbeQqVX9MWrm
58qtaI8eE7qOCQEnBAZIINOcMBFwZL/KMZucuz9Kvl+vPZH2W8UMFmi095clXnAb
ph8TgGP/ZXNr0qLmiYbypy1m9WF7jI8SFce8dHqhpsFHwtxuEOjMNmJ/xB/wderq
VO6YhBdtiEuZitIxQCOGT7N7D6aehh0Osv3zY713kjEK10f7Vc5l7G2Ym2iFQt3G
wCD6HYI1EiL3WmM+OlecM3YCqvdvMlCHvi4oFVY2QyJ4j0Q1DBIjto4A2cH4R8JN
l8rGKKYYaHMnMMdD82vuKq4NNug6BrunBcFosmEREdVz8ifKyv/j0Ws1/6SRpFp3
ZIkV0mke6ayEZgZipA1fQDGN3ymPV27sxyjxercx+ptc5KwFJv6cfzhfD5eyZ3VN
01HEeFApVvQHrRsfLkcz2V+e4m8sVysN7UkfrDuKq/VlpZKAftJtPlCth1GiN7vg
P6h8JhJZ1SC06ae/SA14GFDYpfAUy6G2mg4Dvj+S68G3krbxfdODxHKO/08eYsDs
g7Qx21KPFoWTJBYlGH7gX+dGXquklvhc5nIA4dibLi4G/b8SHYnGqU0AZe9ZQmHV
DXtfGSjnuFaDvLDzi2fqpj5tLZ6torEGhp6G2PJ0KI/N1rQbMdE2jC+dg8zfOvK8
MrVgVuDYBM/uKKrTUkI+HvxZjNRxobi6ASdtFmHZ+7EtBatTuB3pZMYg1GroG2o3
jy6k0A4QaKuXJ5nR5gu1zqNHlUs2ROhD1C9H5Uoh+09HIYBiRe/8Ox5O4xEIVg5t
6cffMxvoA7w9yQ4mMk5CPREW6KJyrRhtPN7xj267/sBh+f5ocgYOAwZX8EtegE6a
/aGUavQa7mttIME8ViewCNwT8QcdKGi39HCyI3ZiFJHNsNxvnAsl6P91Tyl+uB99
m9RjBAY3/T6XHP0kl4+jQqmaKrRTzPExJh2Jw/QcIIefR66Mu+wQa5o24Li40vnm
cQZkatU44pQ2Sxsm6N6r8zBMJ99rRPwxnSnOYw5IXmR9c2RbDm1ybWBvNfBaWAUV
aZzbmWmOUQzAcwCrXkk4nEdRwiMJ0uTWjdt05HMiog1PHS+NnvaNpbhIq2Gn3lEs
PyaWf1KeZtJYgvrbqWiYBXx07zp3YMCC+DZDelZgy0pzPAJR4BbI7/WpNefEwN3J
+80gkrPQW3A32ow8Aq+lYZdLBOUmWf8AaowPTZYu0rC7Gb5obg+3n1no79itdiyq
yR90zgswDXQeOiofBVXoafiiOA/5M0l5MWnFnJsNPmWsfb5fJJziyxaLKvmeF8M1
ZymWxxKBTWSbbBEMam5tS5LFHaPayMhu2UIRVb2sUkysgw2Ia2Bw13CrrGOihkqr
nyd0WkVtIHDK+nlT/ZX8K5iitKY76LZrQzBl6apnDzrMf8AclO112SVLD4HfaOtu
bD5mM0YKtWEpSNwHTUq2xqtFD48EpZwnFyXL+/TgPS1NXBsWVCZ+wtBkcBVjgzOt
jsEbmefVtJsik+J1+lv806Pg1JlgpAN8Q45FI9rOHjFBsyp4rghZh8Lnd9GSfVWA
Bf0tIdypl2RrmoW/Lw6xIPOWjEnKi9nvIripoyEnmE0ioQ/EF/8FUj/oqoN7uiOw
/BfX+nAzYi5A1vBuJC1N2WMAE+vhmG83tGCjXuCxGsMaZaNtvFCYhtqrN98U6Ave
1ZfOJIAbJZg5E9UObnaUVgfQJx8xkqmrCyQ/P2FClOnmmbWiksiGmS3RC4cqrrKF
4aDW/YVy8kS7FK6r3obpWVG7Nnadyl0PL5JAh/j++blKONGvyFOE9DvUPAlXDXjH
pF+OV2Y3QVg/BbYjrSwZnOtAL24PW1/88CA6IF8TOTwRWO86R4YlzneIyeXM2XGk
YQzRw20TGSnHlyyGR8MX/ZDuhkJpjYQlvR0gXfcfh51yLC5OHi2X4AzLdGCCOjQ2
8qRo6LY34rDjpTWtiiG111leK+1/UEx7Ahpnes42nTT8Ll5GLkjxbrXvrbaxAxic
El4IfnLOT/e9kkPiBdfVLtHqDAqCFnER5bsuds72yduPU5oEF91TCXoztjrNhqs7
ilYuGzk/lmezmMLYMRjd9vSKv9OvrP7wMCCEWlthiOZvGUVEo1VKEjGkQP4mi6At
AfDqR+/2VFoqxJwOawQhCHbZ8tDSrKTc8yilOhIMrDLYkSr++zL9AqK1NxnOWY/8
iA0Xh9/KRNdvFiQ+89xPr10h/G2XK0UjCwLmthCnBk4HDknV0H0LRX+9atmNdbsj
lsEF+QNEJDk3Vc+rVa3qAIBBwqMq8VIC/Xc4E4rFXGMVfPqEva9XZ3xiACd/oOI4
tLxEPDPcy3E88Pm93eUG7JeCeOvQls37XUDKM/v65SS5iUu0oA68fX7iG0EgaRAQ
xwrS9OXvB/0C1ZTRrrnea4linzTJhYjLhBU7//fFIRyMXeb5GeP1FYMJnu0KA+Zl
l2WhUn/ZpCqG+TV/e+FqCxdeVbwTQsxdRN37aOHXXJuql0gXQFzxtz3/BbAnucHK
uDHmbOPKUmMZIhK2gqo5pFKD64LtFMUQZM+4/Rs/RNZ4jU/jgOQrsvBJ4N+utYYp
JKWmeoJBj2y+m0Wyxs9rnViFvDjPBoqXgOwuGS7PH2spawWXrMvVEz2iz2cLWcbs
wv0WmFkuAYZPVWNi9ikn1rpvjjbNYyGXjXBdLbPNXgp5tNr6Zndo1jZ3uHySaIbi
QxTzcHIaHVKjWv5MmuWX3ntbpE6dcasuXEdV/38jQ+2IKPKS3ZWIBNy50YTgVPIZ
OKk4hzAGKGi1RUxEwsMSZSGyqnxDK1HoxCTYJ3To8wnJILCMZ6qfQi54yjjpbSBY
leGBEHw4A7G1jKJv+kZUMyTfL+dV+888PEHEZaMDs8H+yBEOVSY/CfGuJRGjWly3
kEomZrSx2tmvxSMZnmmX/yNVFe6aXOSlpS/kk/bBbCG+/bTVwCeNoIRprBWAu0pe
zg7bjIsbmDZhuI+xoKz8LJxdwsrUS6O0KAm+IYsCHCXrfTzjqJ9nYsQVzZFHmhy/
aOMpAuQW9FdyxOiD8xAezV9VCTCTmGwlBSbtPhUNMUuG6IOq241SuwrkBpWbojqC
R9cmbNJVl4i32NqgYeuq9KpkpMhQ7XzXuevivC1sr/hBKVTplpKIHU6M6Zz+hOU8
3ycjSHrloYwcAkbylADCSZWSVkW4dI1d5o0ergvTEDmc2CUPmRDOh6Ltzz8O2xLS
laYsys6wrmWIgwQa0Jh9dcB9vwsNBUj+mTQkHOTo+RqY+s804lQzjvCgOX8Wz/iJ
ODsjAk2A2o5k7oYJPQOEuUAnEwT9AB7saiQG0EnjEyYlSeZfMFBZyxN7fJIiH5t+
Ref+RCqHWN45+9KDP1WuDU84WtPmsJ+8IHO5d/DYuD5Gr5Q1hnDHG92mN6Hgeznk
LPwKCbRtz267Wuv/O5AxG4yRfPSkPam7EimfIXJsev7b5yxAdAWGp/vxKycFLkOn
WjJD4Ox47o/Y5ofgzertJ0ZxhDd9T9nRy/ki/9vl458dqk1ee377j5PG2nTJbney
/ZXw4y7pyTmyiZZK0tUxU0fuAtsUz116+DL7OVmUBTokyJe73FtUPEkSvtPFkLyR
f63Q6+NZ+m1EQa4yV5rbZKFM+tCi6OPUmQbgg1PNolXf1wl2WUF7g6LTofnrFXcZ
M6UbMWK6I0sMRc/C89NAJc7uiNT8Ih+DmFlqNGa9HyvdnbB50cX+xqY1Gpc9kYV7
7muB7OFiHZ89oAmAmhi79Lcg2DsrKqMdGm9FoGTAmA6VA73yW2KDjNuSAd/v8Jq9
hWISuXzb7mno2LQg/MkRfUramP7Q2xqnQDhCesBJcPAqxpehibt/8Ia+YNWh8v7R
SWh4mJMv/2D8FACoGeZAba4j3K5k+yztBQxqZbgijKMGf+omwuWun9+8nDdIKMOh
8LXLTQ4S+83zrbsiFKCJ8fwzmV7+iLozKsCrkMuNwcx+4vdtXl4T9mA9KyuksY/P
cjlREwDwTRZxuGuT03Sc1gOP7xyNRnKZWACbgnKDpaYS9N8Q+ISUe40iAr6YI5La
EaP8mwnTz3p1pk+X53uR4AMES/dX4NHSd8TtQO4LpHgeS3mbbIF9EsybI9S1LjSd
gSGwO2iegg7j66djQYzaPECSE9FbQtAysqBbhqcx5EWBIw9etcJAwqq6dt+nII7A
GfQugB0fb9sYrVpaFZYhrfOLOIzLjvTIETyYHPDixy/bw3oEyVvYBFNsrrmWylsB
2iMqS1bfrOniSDt89Wud+/JWYRRGecisXF6ACtrMGXGYCoagUb7/H8LOqsUUFPJN
rGJGD5deC4XsCQLpvwnwFFVMaKgyLZwyBSqPB8I7UvEbohXWJAgcwHuRpHhYOmhf
t0qSsjYA7NNmdwkKFnbRqUPtPVXU/iSsH0xhNP3zaPqH51+s8IjhHAhYXz1FzyI2
y1qQRJVe+NvEj0XqUBPiunGWW2zDQcqFQZ/dOr9SdNu8xhc0VU+RkfGeVxjk+L7C
AMnpMXg2ZrriDfBEpF/8cNMt9eXrTn2a8G1Kb5Tr8JeLliVT4LBLdjoyB2Am5zM0
fZCwL4NbNiwVS1tZ+ITxO7mAsMhzr+O5QNgoptdHQnCoawfbNVbU2lZieas334Ja
Yshr42Dqikt5Xt3XWnVr2r+ChaCmctVUvRNqk/4LE21AlilWRhr50VzGyDhYK6TQ
kfTy/b2vO00e4jDVVnDMJ0bJ2ky4toTQuWkk7dxtAX9zxtcIrT2N9xTsgAs+RtpT
VFCnRTZmgNz1Z1qPcGc3/jBuUwOhcV6OfPi9GJ5swufmjKaGKFj+PGgxLXn94JhR
rAjS1BFPV3MkcdyO47xvMBvJRMRL5J0lE3FNbI3Y/5owImfn/uqmYilvt3U6sLrF
dTKMF9t4u2Ba19jlmnlYLb3424SISEmeftivyNbkY1gQ6dWtlih+DiXvceWmF8rt
OwmgW0QA9UoEajWS11nECAM2LPNdHMjO2Ah19Mv6p1jvxqn0R08usrbe0IMU6qsa
Lv4FEnV61BpaIudn5a2ajfYL3PVjDgNpkD+pKMqwgbK+glJdT1RAzT3+C8mup2uZ
hBxDZc8t7NXco8o4e865tikwsYrmoVQ1ucz5E3C5avHQ70tffhfk6g88SaK6xA2B
kmv1RM9o/Ek6izZeEvDq2gC3fP8I1whsybMu9nRLKZ2R/Ao1iIc4PQx7e9y/078V
IQeidoYC5bRVykk6uFf6oYc2j4Zt1wGA3/JBtT86diROJjEh15U4IIB8raZWwYPK
GqnnVeFaL6kno9LReTETZhRnqcWzDQVULwPWzTqsekAbVOJYqdIyc091sZwLbn1R
0Dx8F0ybaDe+qfDQSc34rpWSt9QrzMonf6tndXJBLiM+2FUyQwSYZuyIT/lOqTS7
vtUUDc+tbXmwYOpT5AALmN3EjAvzqlwTI/GJl+56s2fdz82iL0fl3YBnJ1MZQyzA
BOQm1BtQ3H7jztw0uyk/9FmY+oH20H3hPM89sSfhjkzjDa74TkIgrxBcqkYEq9E7
E08F8hALcvm+mdXxO8XnavRNYeCNVHCvOAXdPYd9YLu0pzyWC02dmo7pEmeaNGyA
EvQjhXuH6hOCFYo3fK45NsT0OAox3flEDGQk+1hk9Pe/t9wWSBTS8Hu/cW1W1S9k
3TBFCyeE8t/xpHo1bDEVpTtcOgU3ZXCs8LLFsvBRPV4EvFwJhoRvoHZC5U9iTvCh
pJCT5qAqaUQsF9pH3x2MfwPE0Tg2Kf+u1uVqFp/rWW2+v2dqEOSPLrRqILFOMMTn
okIQ3UQsAbs5034e7dN6Db8dqAY4Zta4cgHp9GCd3DO63t0e4NSZk8ykhrF1ks8+
93QuNt9FNlJMVZFwJ3PuDdARRq2HiiH/F3iJSTPVWKx9JtnDtJCfTjb3TXgzMS9V
nwp8heGwJS6CjM3bQxG7/go2o8nMZwKITJJfu5EPOM6cA3HRyw6osLxU2MHlTH9Z
7saJK/QZej1I4cQI7YVN25eKzG5vRK+L1gS9G2yWMsnjKM1XB7vQT8LyXjQddyPt
NfwIaLbEPOWZQ9rfN9wv8W+nysm7yRs35s7lriNgeyttPjDFE+CUmXyYjPuLpJq5
5Fl+tuRhqNk/eVaJW/Bddg/tVK10julmE1tnXkmNYqxo4bXYJHzUWQkeyziSjW+M
aDZ9yxcVi7bYXhZZ+jRju4k7C3AzwbLdGiHZrlyj6QN4k6QLujdyPUmT1QjAmAJY
iOQvigt74D7IGTVbCCT6CYFerSi5QeApSrFNc6G71kU+A1ECtGqHqCZj6dhvlzWq
ESiMRDtFF7pg8NBeC/xOoltQKqHjRlHlB2BBieBg+hokaFUHZFpZfcoh2uIFT/uD
DWvFL4hEIah2oQSQ9J4xS/UIcPJNbXDhZm2hxz29tdemQ5fE+TpmAzKwbwGA4Peh
j4OP8B8E52yMri7h2kZwiYGlwRxNy7bFbHeIrBXKieGU4pm0qcmHaVFveXqvkIPl
vfQvWVVEc/ncTx6ujVmR2D3vcAWu7DXODRObwCqUDHm9WoBckNSoEApcV55jCD11
t2FB3LLbZkUkpE4iiOw96JYBTzN68hxGnkB6gL/nMgLWFxfYXyXb2Luhlotog3UM
MmbPVEgBjVtXXHrE0b1ykX9aPI/PI3zElvMqNUviBHdcTwN8qUJ3YBzFGWAYWOpC
6mr3R4n7oPge4NuAa3++e14vYsqehvejrZQLpMyzQ4K4Oc2Sl7TBu6L3RpyoMbMF
Xu0KAYZ0fWB7ohtI+UHF+gWTjz/FObD7eO4K5b2BbdFVmQrcpHBROm522Si8bujV
hP8najp7h6Kr1kzgYlPAURUgAhc8MbabNF5NizU3nmpqbeyhNSQSlAPmIK2phlAN
i3T5hwuixCg4wUI8Tw51ETDxM+m+JRwsDHPf32LDGXb9dOWPRt0atUqvrEKhLX6D
EAwXdK2DHXiP2RZZHu5R0GLxpJ5a4H4GY0bmCumGVt06+Zjd402HLykTrElHfChW
sxA/5mWnifrK+LvvTaPw41AWfiNzkhjGWcGL0PwpAlyBuUdNnT0VV+u4Mk0VS7JO
Whzlszbzgj1Xz6HbRxMERyC4MOrrlOS3pJoJ895cxnDCnmUdeVXBwsiykj+/reBy
Iguy680YXbzmJeY1RNHfkSAIu5TSjjOuGnbHs1pBU7eAzseFw7l58e7zojvF6BDE
dj39HIiG2TxBHncP8RvYENwn6TegitLECxg1iGgOyFB3wmU5unSN8wVwFwWgy7rL
kHcXGahvUhNWtnVGn1+khYFwf0AfFgsFhliBL0OVqkX3ezQt5uJHSrzQWvYDE6ZS
5Dki0pnHpTPe//7qBHB5JgI89+oS0VaZhIdPjgCAksRgofbr0eZeTKKVJiqpSMCt
8Q0TqxJu1c7Fev+2RSDVTnHF2oOBZcwAk9d4O49xKWudWOuDWNVD8NYLjxGs/7/P
K2r9iZU1foBqM275enQKByrqGgb05rDG6yJlHqe5SGpUtGfRZbCrkBarCJqAZd4V
2BXePLJAJEPzrdbDFzfjEmbd9y8R0OHsfU/m4AAlVo9s2Dkp6yhrXJijBW84f8HV
b6mLKhJG/zwYTB/yHqJFh/TVZ7Rcu237MHxeh9Am8NOvKGN8SaAH1/AVu0JB9RMM
Zg+4hZTGYdkLco9IfH0YDjDjPFtJK22C/Ej99CI9eybmG34a7d59jnxEVNrdVOZf
i/y3l7x2TqA5IEV/emDwZAUrT2cpsMwnADxuFP/pyJU80vfY276pQQ9JdJgVCTQ7
sIXVv/d0u1ByzeCh9gPkLzhoXK/UXPD3Ftx/weX1lcoepyhXJbxqK2HpZzQhXA3n
sOaYwoN2aGQihTgCldCkk+M7xjCE/sTEde0Z71c2pFQCZ9YhRqVqUyz9DfyPYQGC
Zf6oBEp19cfR7IOVIh3xHFq8+mJIqoCJLwodMKEU7hhsZlEKUVO8WaJWIG41fq/D
TsgbK00C/oIOKNLoUjdLsDVU/+sE9/GoBBWH7Is7rQNW4QRqyfyXzVYR1dYSEAJ9
J/wfcsedZ6+cjcPFs+N2TZsrcfc7ob3DplXz+AbpJOrLB9zp6Lm+0W2Xnq39Eze4
+klSC7Sy3Ig3qTUWV+ARKSIc4ra8nEeSMlZUVinJtRF7UhXNSy++ZjvZtHVLC9wN
mdqutzYDVKV5n10uW9i4kkzCt9/Vho6IwmiZsflt9siPkGlInSg1V9nL/p/jiiJE
7eAg4r1FV7EyRRgpzYGiOjPKrOC0Ch41EVQiAmm9zsP5sPAoOmKhOIfJ4EXJcUCI
194+r4pObp8BJZIgEkngFXa6jRcQ6nITq7LCVL/+XwISTvMndmNoCWpPVsQfTH5y
oFVESfxpwl/2e0rlM+YAOjVcSaSnSK1YpTeB/vFJ0WExxMTtG46e84ZxI6MQPoEO
zvpJmv8PMDVmrquWrmM53St7Z1DEeFU4ML7vzFHDf3r06lB+91VExCzKdjSm4gLw
xuhPfeXgSYI/rLNHfRAhLMNBk5++QzFFTnFKusD+r8qvASVm13WrTT0DWKeszrvo
zstN7tPczjVnvtTyMWkk0LSZR270ErhD/+PjnbgBxF/978GylQhpvSXPZcEIZVI2
iiMUd/F+GeCi1nYrPU8W0/FzDRbxgLwTqtI9hS9wcXKwaf3SBfxRJ56F9ULXhOlc
AWxSVCV5yoiQapd4l/vyYCw5QmsiadysXV75DtuROtmJs+NbUV5rZJA8G8ebHWbS
GpX/pB84b27aF9WeAra8Lv/YH45kFy6z5xvGKxPqYEwx95ip0690aFyAdaEgg52i
Wg4mT3Tipo1gNiwniw2k3WTl6FwumIiGrXIvqWO0ac3ksIryb/OiKQE6xCSslfbo
jpFz9hhwUaFnL8i+W5oiR5A+5h4ZG5Je55AhKc/R375Ac97jde/r2qGRppCwc4pu
Aqr5BfVQPc7Pt/ppJWlJUrZl8Y8mkMKjORLGCxwK1U1f0OFjuHZNuuzoeLcykw5D
KBGrxcaoGL9SQ6quSY7YKvz1TPoYF+53P+skzqeQ8Odn59Mn5v2iroERsNj+/lvK
Iw+ap7jnsls/r9nMwABbZBhSlF6WPBw40SiGHZUt+89E28reo84eKGWG2bX6Goxx
zyWLYzxffl8kl3UZJWsGOLmTPWo+DZWLWH1trSIxK6ISYXzarQQS+X4wJ80K5RZN
dISN5REqRVQKU20z+WGLyGVEwsKIjQAnG2kT9jhhAz18mk4UyLvTQ0hwePHPncvn
yQ/X12cz84sNPNJnC10rcEqxm6junG8ckd8MtMQ/hXDUXuK/IgLPiDyOShNtLjxG
Tl+v5Hb/eygYdrVGCc6uRptmg/wvBPxfG4maBqtlF2h01DTEpP2uzB4sD3C651tt
0I+nFXkOYEMtuCb9ijplDootMqTj3qJTT1W66z7skI25vbkwW8dwaKqcQ4ABz43l
2Pi61/RlI1/giW+/xEC+v01/eHzg9/gAh/06AhxwatwNYlaIoP8j7FXCqzGjLuf2
qg8PxrOzUUNMzB37XfYkTAnj247yGtxLIPMYbDiAdGStwhSS09ien558zY+KfKYJ
e0RPuY1CsYsxfhpDfSRycQLZTpWCgNUHOAcTVtOeN/qPtOKKtYsa/nlP+CPod+Mz
32u7OqtHcrDNNF+DrwrODGq+TY0Ct9SB9Fn1cErJLDIbzBcCEizUbDWCx0c14Jfr
KhjDR07VKphlEvnhx71PU04jVWd2sX7jKDwHk2cqt43XrZ+7Nu2fJQFJiIAvnZKP
9XJ1s5BUeVecrXYQXmfYrDmq/KH9bqzelbT+/Ih0P8bEv96rSHPVRzHFie3UyRAE
ikBgi+W/T6bwmtfOP9CyCY4oS9G74kQBxCGVzCUuci4JDJPsrk6Xw4Plxn2ps/76
96W2zhPHlM2O7g4u7Hl3X/83NirR3TRdBYQ+uzYYBnoBihoY4k2iwUhYANVDvlwL
uA5Cp7U7zfLi/rFD5RhFsmhlyAy0jmJEei63hlYAhPk/2ZUWYVoza/bpaaC1tOIg
SjoR6A2/5DYux86w6BBhyFuRhdL7rX8duROIisQGWHOq9DgOp+AlXuuIY1zJV5JZ
t0Ma7dGvuiHyDhQvMPlcT0D9XLStpQdeprmRpuEmQo/gkpAGEm5zTpAPqEC+dwr5
9W13O7uhtTttMP0l3nVnJPG3YqdkqXVvM7+l59FxV3LO/xZ+lswftYiHb0hpzCD8
XMtkc+uYvtcpkJwS1YoWhp+and5Tj2BfjhN0luBFWbTJD6aT2mqUWYbUfcip8W47
yMBdmRJAP4up6Yd7jbO4X+syfSoYAUWVCZjbLLv4iY72wKLwta2EoccIr3HUrE+Y
GAJsFRaiowA9o7zVqipkvpea9NxpaUw0CAqy/5NxbO8FqljfMNontWFN+5zt509s
P2J9xxrmQvNJyaOb7rSRVffb4XobRbdx5AUVGza+pQKCFZrusqXBNjTTWjNziAXE
bnZek3Nol114WawYiOV5knNvFH+M6YnvK/ckxuZFDIA6g/BN7otF2SxHQmdFbGVq
VJbN0vmzAQg7ZRKixtzX3/++ibE/e1YObzzS3jGr71HurXoLpNApNsHrKBah2hA/
QXJBkhAV80UCfHnO2erTmReV/eMu6WbZvU6CZJ5B6E0sl4LNnF8EGs++dHZzROJN
18Q7x5FNC5FSzFk0OW4x+LRMZKdU+WNcHtWSN45U2DBUgl2nAMO4I3bPQzQjaosc
kwlfe+DoPkHe7D0rRsXFXEBjfYtQ0TOG3bSjzxBpjIqm7wNhMTUG5J6nkWVQscYA
riHTS9nxdshU6H+NaF99qmg9ZPsgZ4dyRv2vNNQ1tx2/vSV3+NrJrtySjE48LjjS
EjLQim9J7m5++uvCYloXSJ9FwictomUwByemSdmTj34VbBTro5nUihKzksBh9hgC
Pcijkq4wFT6AIVHdLJRr9uEE1fMIFAITJvGBpBTuTZb1GN786rCc4pkecrMJBvsc
EQ8lRLTQzOcMboPPbqWCEoSCJnbGU7csBJsmp0a4RHHv5Puxcf4uF0d8JJyc40qS
GfRvi6PBQj68UNX/Z16ivFL/EOhNKylj5D7hGSd7XS/EItXqzOnlW/dvVWhrqw61
8st2EziQo7L0inBaGSZriA5j9DeZlcoNvKUjzu56kDNOugqnMxgUycZLNrL1/2j7
wD3mp3gbg48bYeHCT6GyTqo6fLFkYtWwExC9v88osyXKMUW83VrSgusm/kHe8zOg
9GH3BlMoV51Yi5ubKjb1W00aj5Hf840xqcKP1ZMPC3iu1t/J0hnschhOqw2w3iLu
7Fo45XQ+cMti9+44Z8INdT2o3RbKdw7sTbsMV9x329LLJ4qRYPDzyMiCfS6D0wK9
4IDS4SZMeYso+mKX+FZUQO1WHGx5LxWVX234unzyNlNeDlP2yaaFeMHOEJ0RWmWM
E31GSbxQCkP5CgJSkxMhdXQQYEqr7Y78Dsg4Va2cthkU04puMBtrLFpw5FXQtZGY
qGzdYINh4yuHyAbbvwsIFUzXmfNzgW0yOH08SplpgS2SiiHWzhe9+0yqTOZYJBZo
NFVx1YArNS56MCGUOGOEv3UiyH8yKpapAjjkJtVDFaZgQmeebIBAtJk5ufV3usHC
YMjHoFx/+dVmF20FYDgHUvRNVgqY7tIIBG/I9g/8F7kgONXP/DClk7yWY3leesLl
kZcF83185Jhg7kVjMqH3W9xKcfRRHB6TgAFB/0kaC1svEt8r32wBp/gc4gGU2Vtw
UhaRYvxK48K+9GxpK2FkNkrmLICmfOtEj+ST8N2xU7ZGSnIdsfo3AS/SdlhTgn1j
CdaLKrw/n2M0Ya0AwZVj26nb8NiFMyG5QhxVOhmAULD27w5kWzwURiITC+6g27JO
qWiLCSelw4rybzslgUuRk4UZhayBV6G6yGKcT8EnvOJ3vkFfL3jgq8v0e0jDC5JE
XiS0Hu9v4lmTjQQGH0sNW70GW43EpUbqRvPqggRKhNe6BctNpIwtZtBiamffrbC5
r1h00424jG1IwQZFeae9XhVDdzFOOBJ9m7p0zXv64GIblC6vjG0OKeFu7Wufnx3U
zhL+i8Y4XdVG3zdgZOoykj27QnhDfLJEfQQ6OXAsQWT3V4l/p3yxUK3uUfgR4CVu
7DE3zL0TSeEwmQAJ2Awcyh/BForvWL4298CkChck3MFHmK4C5Ui0WvaW37WVcF3M
3aie0XbCNKt3ECNKA3zrzen067BS+xX1SZ/CzuTPI+5ROyFCrgssa2Bnwkvjlg5A
0ShDsw3ThYcBOuqSi4vp7SlODp7evn0qvLo1TTiobvHFmX/aufg1sf26Fs4bY7/R
GTTkSmIcjtDLXw9VtViZgFFYy0ups0bnaZaXv8vbu6UTzEXkCPv8ovfFPOWuK943
5c7hX17kVfzEDm1RiyXYwgthdOz715rb9rOLNJELhgwihATZjYj+GxoTF2akz2E+
rduwtEsKGVP7CtDb7R+r/wwtQ43elebKoMi88dt5Qmgxv3NmzwJU3D7P3qqb/1Z6
rmqye5Aev6095P5wWuXuVQbGe0C1ComGjbnE8FtwoPXqJCuNOlg9r2TINbElN72i
HUeXLqmRVyqdaYxFTcR2p/DCUMNT+12s02T8tndgbFFsEx6e45YlYC0da0+Odw0y
6gaTgyb9TtgcAsaX1splu1f+PynwgL7YlR64CQhvrcfst+WDGKyPg2lRMMo6HkeG
5m7nJR1q9jCxvOlapk5mYVPhIHTCfuk4LyrAmTIEbn7jNyzvKtYhHiFsSLvoGdS/
xWjFvGRWlM/smelml6CR8k9aiWmH7416AqrdQmwGu/LHAqUjlGGQXwqBd3Lu2YDp
eAXiUCon8myufkkwpZoz68puAGtO1io/DXq0c5cBaVRWzGFXyHgghKpr5krz5vJM
K9Th1OMJejpL2qMZPFIUco66PuJQYVl2XGva86oJ7B2thKe7/Z/ag4dQCeHqSSt/
2+9BOZPVCM3SkiKq8KrKg3TRFCvNhZmcBR8vAK/1tGYEF0OR5sgKnf/Iip+UmJDF
M3Uz7kGgQl2Us4ijlR3GTlP9BR/+TykXcuZwgjHAisnZ1EI3vdazTizPSNzXwjnK
2gGeyBkkqrqJC8apEaHKhIRFlxARiJYrfTlUG5qkTIN3GuG2mZEw+qz6ry6+wePh
YFxOrp9z3opeq1OQxbqnbef1TR8kLcXJoPUd6/l2O2COKxhNdMdGmACN3aczNyvL
f4B1Wh0BK3JyfX9zPhLM5uswdN/oi1zGiDNF2SYrsbtn+kWhHV1sXDxA/ZoMOEB5
Vf2KipU6kvxtf84foJUXpIIrvJz1kTayQbmFfzv6u0a8O0/+Lh98j9nhC+kH69Ve
2RspmWwwVIAE7ScknaO85qrNb12uwXrKJqNNWXR9Xpv2RY3Hx7HRJY+cI+SJVjjy
eguGZNEULHFCJn4E4ktwwgIjI6u7FibNdYaDaMaxwDcnx38kez6FLQuRdjPe8+93
FTXhLoeqVbszgDDA4RDgTtFeRbtqvqvHtmWpfP/YjoHIW5OTH7Ve4ZP5ZvWj9v/J
rSfe0SLhTUjPxDbMJ5HDKvGYWp7zpa8YrhGo/EwnBSNJ9H65ds1C3Rcl6tYA0syZ
asURi2T6uVfP21liQReuv7AE9E731jp4Eb8PyxYMIChQ2qYpM0KgSgPdqxxNFFpP
XdsbBie9arc7UMzrwqZ4nKM1AI1iqi6OhKP8VJv0rEqA4PTg7qCcr5IinYL1Dfwt
d5D3/4eG0hHvCoBT6YFVCuarxZvZ+iAI3P0pU8gDLSLwKnFBXZk/dkK8h3n5VuA7
83vJfneUmp2glCyYtJSPkziuySVNHPLjR9Q63/kvTqxEoPPg5f5EkO+zZMsSub4A
njdOxx66SUkbRpz2us2ensJHP3stxGYhQ1E+hDgaA6vOAkxT7TXWC7QBHx9mt9yt
Z9SjeABNcTCtbcfNRpGKmA+p+LLKdpVXAd+ZU8uLerP8Rq4+mHkG85UHvH7EAZsj
HpAv8P/9KqVnTwbkEjbH/4jDMWQp16c/LdlNX4hWiH/rBL+oRIwiMDY0ovbvXy8J
9WW6M14DR79i//d7A46Ys4vXNSurdDcbC9uixCoiHrZEIs4K710XGALIrjuAG0t8
FIn/MmTYgHeQOZsWWiDaXt/lpXCQUVmz3M0758QoZEpjp7hPVASGp1QNRMgZ/yW2
A0Tng8nQHr7a5x76PZiLujQjsdjuWlP9MhJ8zx9170i7Lq2ssWwEmBTAsmjth+8r
rB5vcgM6jEhGW4gfnPqsxZLdldaBGYjb5kquNRXXaQox2k+bBok2SyT7Wyvw+Ti+
lwJ5AydV/m4pHYalmmd7CqUcc/dT+jik0T/5OJETqjLrjflPiKxeMukGjQB3qVgo
MM2coSXbDF/2Ud8HCmk4d6p/E+Qw76Yn/0cEVlaeHZkVa1zbocH+72M4cEsGUp5R
NAjCnXLPU9rQR0dPOXC0VNXxldetdyqmwMkAuW4JZ5mEyKhEzDZmARRlZF38dMzW
5ZkkgdNXkvG7QbCuMBtvcAN79VswiGjkOiAxLuCHFXhFnnL0s07khueuhi7u2/fi
b/YYLLj6yWCOsmVAQYABSYM2qV2B24Vak9YEF2vrT6s3TZ6nNBpQK8nsGi9uaxHb
djWBDAvS415LM0MEvQ6yhqKZTPAunz1timrMufAqP2ChHioL921nmAbajdhEC67y
fHplzSwu2yZmsRMigelV0TSxEsKJEamH9TkziLZRPwoTRcX+POXnJmswh/jC1FEJ
aFxHfWd3rE9FInZ9oj7H52dWfy35+ZdUjJnz5cc8Q9jjzWk6s7dB16RnDizt/iWD
WMY3bsOuumcdBM1RJmwXO0O/23mmDn7pnEiY/gb65nZwHSZklH8NwtRDCfKOP2Vm
u4ndllDPZaeos6SaJNpkN058OOpbpMyjbD5D0E+X7cYExqjLyiLuddrfk21h1CTQ
D0/YP960p/44PJzkZpN55Y0qyrnxQX5u9iPRKR6IVAPwWG+3Bw5r/j1e6c48Yemz
ne29El5C2Pa7X7TSVMOwg4RI6QF5lPhCtaATPVaC3XvA6QZUAoBSCKktg9MMW2vF
4VU9qfsU5BG2ulRGlACc6gQnIFC8rzvu7bx4OtP7DpXPMyxABzyhWSSjyz1fDo4j
TSXRLXIoW8zxJ9QcTBm/7Le9OvpSM7j+fIrfK22mkptmPrUISBcFijrOQGiho7Wu
7MAlLFT4MHYYuCpATsUtrehqHZszNPZ6NfzfvWixhA2jfhmj+zgNykhrJ5pfMeXd
57yp8TcxFZe7YsU4yYotGdAc7eFdJR2oxo3HSqPR07mVOTp9DA2mSowgCZh+5sXj
u13V7+qS8ejTSMYQnpfc7BVKhqkrOktGYaQcNy85nqi4OgvvkblTns1fKgf9J8jc
S2M0L1rd+OnWQbmtaQsMOIHTLeh7bEG00Nh17/r7YCQbYMzVbHhF/xOz4uA5zvyo
3+vdI9wywj3qMsV8rSjatREQVDDNA3jXgpAamO3EJc1k0KfaaafJ7ZelvOXD6FLC
dYnRNedFJJrS4tTDEmjn6z3FNe/Pi7FrKl10ZZb85UplWecIUmh2RqeaeuGWSPoW
TPEZO5QX+VXm38nxx+vIpTQtOZeFg3WDl1GG0SFRj682JTkTJ2NP3OlW+b/FYRrr
rzQPW+LRNtxZyIUri7/olMmWp1twY3JhGQ4ufCra8oke/pGZPHvdi7qQM10Qx+Au
noHLpVW49pm03c//492UI7eaIc3O2sL7tOMU6qfF5XS644rKQSu2EsJ/CCxoNkxh
7bjWfPrYgy1XXrC0L8Eir7ZH69V/8zgawxxtmQ27JkiyLbt5ggBB3RyqyKSWuhnZ
jL009JInICd1gTqic+mbSI+Gi/sJJQWEL5tlF4+rzI6hrav/evNAppSUm4DZ8yj7
S7xnNUepkq2UP2ryNP2jGOej47wcMemfjQ0yDJJftG4nTYPHzX5eXnWJNomZtLW5
Gr4Amsg1y1GdOstPdv6oqfsd43Mal3LYfHi2lBpsizDJhbsAnEhL/WMNClwqjgm4
U8EjLwQdkAvqvsQkXMerP1huYTLvaO8Lp/JSg6lh15ZQnVhgO5IEI6Xkuy1HqSkY
4fN35KJKz7G2/l+ce+JnPXQq3CzZKz6dO233+UiQGkFuCPTthmgrgm5zJTRHl8yR
LvezkJbMNbE96wos/RLX19cS6ub6gpnYuQHhvD392mlLfUFk34PqTLChS+CGo8Ln
2Og9jWp7D2lLcVv5o1Jph2H7mTpBxxlzNhuowpjvD1p2zMJXl8BVVMRe2Je1CmqA
1XxUHFXFgh0bO473sYuggGtYFZja6Rn/318Sf5H9qZrjPFM7tmkVVax6H7RLCa6v
aMViPeToEdt/VUHUVqYwuDfn4800lHIufjKObOLbID2hlDhqomrmVIZqLojB9HZF
4Q0TBQINHfYOvKhkJFpPPy0PwOFuJ++qA8acXCXbeMwZoRV1Dlwj6BtfHp71PKVR
X+L15tFT6u0qnXqBSjx5iWgNX6xkUuCW/dqyZ3UUjSWa445OgtFrqWjoagpOZ0Sg
lgSvWqVNv9dr4O8SmC7XR292vV7xNdGRUnKu2O9vU9nTuVRLjhhIZcSS5JDxxou+
kIQqryttYOGKJ4i5267IQHb4fVTSHQ0/Hwdu0ID0c0DuXWDvjUMX89rSuf3VwFRZ
0YPhtXgtbGlocYhV2OTlZpF2fI5FIegyUINUGYLqrHlQM21WS8IxzeD1cEYebzpv
805m7rWL95I7X+CX8vGzaP5EVIWDe5TmY2xW7GxmSOqTX5T2rVnPt9KKPEZbntyA
k2kCuy0gVWvt4jQ6B3Bq2HTTYCw6VIXz2obb0OSuHy+AJnNZG/U3IbA0FZld2oVP
d3zsUk31ZLbZ342rUtlnx9tZp8YPI1L4O5adR5VkPnWb7obf0Fjfki2sjNRwUciL
PYL77+uI+GobcR3n1Pgp5mQylKdVUnaWMoHEAvUPv7Zn5yorGfkOKYzIBa7iqUC+
gafHmvQjwmm1M4fP1mL7IEqtiSrKinID4XuTjDOT1fzV8o11tQrYqNmHRvLniiKW
KnEe1jP4D6snifSRcGIaZmAwKmBg8Ac6HUbuo/xOkbzv+vKL+bNIYFp5/aSNFlNL
ld1RAbk2ipglrU9KaVWpmhueMG9h3kElCu6cJatyRp6eb3oMeKxZUtnAGA9jZM9e
2aZ+Z2m2v++5ZqUYm1rhIkx4k8WRJg2auTNkaRtscR8mddQuWBvGC8a6lriBpCV4
+SXbhIb8mLws1L7Iq5IYO6fTsAGsaCDSyXg4neIOEWDQFHrvYyzBn1ySTWu2rGUv
dwjTV1gr4jo2u0BboDYxSO+zXCth0P0zdx33k1JGUPK9OpryTlzSS0CbauYxM/Ix
KwyZ4Bwl0brFAg1XtEypXIdkWO5H9SUs2HzBMYqUtnpiANt45Vxt3YFmoyl0ieGT
1oCRzmjdy7w59/kk4sToHUyec9tDioqPFdVRONFEMfNb0ymifjPbToG3a84CW+dX
57GFsoNHSy4UiT/c+mqeqE7SC5t9xsmjn0s+w+WMCNLdPnVzntvZsl1Pl6fg7z7v
82Kfo2Rhlu0C4MROvw3SfD4jrudQRi5M9O7bJlZVvqcL+xj6hv34ISGne9oHXa6o
Kz+3wyoe1WdM3tK3JdFlyR5jSa0MD3iJfqvL+5DQHdaUwK6RIzX8GFjFZDhCAug8
xqZiUHPAaC94eAYFckx95DqdeKnI9sklzRSGXhqypo0bPW+HujDixdWzSXspQkmL
h+eQVfVrvEbBcU6ClwhFHIzxwTgxfIV6Ak5a6MsfZwXG4WOiUHViwYZ1Dly7fcea
Tx+ZoJH+++zI+/K5JQjTFRp4YS7GKzcRpybSGTobSMOMyu9LPkUvvqCZTdoF6T5i
yP8RGJ9sm8I+iqUVa8Q97ljuv4BMQHzzbOS+k/+wNUrlXn7F3n8z99NRwsmGiKkQ
fSCi2/x/jcd1ToORITDZ0Pj+tmjMcOAlg2aBpO00xUJyhpPlgDqtkhrmc2pkYQaM
AUr5D3v9xtXtKtX5KK226p1CetsRp2mQTRmuVpmOvPDC+b4sgMwDlijoCAGWEu1l
WXylHVYuisvJYS8pSqVMgXBnDQrHRa4mTqhqWIrZelW3xqMPZrFtIVsdUddEB0Ml
m/00ixFuvqyzlaJMSpxI7liZkHzj913JbyzpiTugMdkVf9LIO9IIgRldxNOB3Zfi
oZ9xTwaDwS1VIdZeguWmRYiDPX928kTLXlxiy0BNzlddRZ38pbdFlvYMy0fkoxYd
cBPhARif7giBLkZ+eMoMDqdjCwQ/zUZkXLTXw7k+h9fOhdnp19qKX36NI75Vlemi
5WefaBflgvI517ABRTryUczE/tf+8BYihgau7z9KW2IAhQqqdjuCs46ba3Nw76Na
m3mhIelsEA/QmUygie59jPcd7lbwr6AH57bnrF5iLl/R9lseEBRVWBf8DlEUhYAd
oA28EZTGBYCa6yIUde28ZqxZNvAt7oVDeOqI0DU8+EHsq+R7HGrbT1wo0SMqv604
Qda1lGubqGfUhzJRywr86KHAdZT3YeCDJHRWOUqz6nrNr181m8pi7QtAzrQ2rsCT
1ezWkR761ghb0WKDps6/MDSIWtpvtcJCqNz4+GmO8B165SIqP8USr+PDPW+hEERz
WmKtC393z5l4GJY0lTgex/NJ29KHZ/3N89Ky/qPRJDqEwGauhlDCQdBMTWtmM1hp
hkBK48inN7nHiKYbdPX3Sgn2t/8vlKdeZxywH0KNNtr43G/OuHSvUzonbqnctFsk
JXluD6Y/UWk1tKEYkwk44WfOOPxz21Tt4ChD0pBJMEg7WOii6FFyX9PLoUjmSMXK
zHYxkVuT2aQF0RH6faFcvBggu4YsCbtZR34YZ12vG0BihIWusXVqaPgKvfbZVect
DU5Nnsj4irSbF9CFa21T0vm5hrig8G/mIBOBtMpmM7b62CA96grWVZoZ1r5SDMW5
iyuK5wS71G0fQO3eVk7WRdu3FKpNpq0XsHaByBepRbeZF0xnPax9I3eY6L45ZYJc
8ORQA3pIVL2h+8yQGUXCNjWZVqtS2pT4L9j8duBO3xkDCzLmbEKC/GN+NRdr3daS
CCKmOrPK8f05q1LWHnmV3hiRtuMUwwQdoC0wSfGr/fKmzJVPY8PHJ+V812ksamaO
j7jpD8BzJPe3jtbmrZEvpMIoDWS8LMHvzzRY58A5Dek6tPhFiSjgBto9tk3iOm3C
7mWMs62LwvNqwxYlJkCWtzYAODw6/qtBcCM/mZjKV+GjPLamvyY5Qo0YEjxb6Gm4
oWF41/kaj4TykFYzd6VrRsCuXcWOMQE1qcZ6v+oKNL4w08UY21t01E+A+0LAezzD
61VvEU1lvlxXnTjcuhnuKXlr1PUdly36BCDYab3qHwqbD+UUEVgjsbtr6Wvbg3Nd
u92pC7B7DrO9vh0omp5sDyUylWmFAaUOo1yLq4bquRaQMcKIQE2/1vhl4G7g34Ie
SWH2h4zaM0/XJb8tQxh0YdmfOW3Bf4jL0QfxA+YRjs7khpokTNSM5IaOlA0App8B
ITHGfvLHyUXLIYX0kABUGtLnIB1TGUlTUS98Zc0LBSZQImsn5S0I6+wwFJBeab2t
axylQS1jC2fV7xUxvt3l6uaT/hHJe6JdQ38Poo6aL4aEcizi9wwk4cdI+cwPK6m7
1dLtA/OCpo4Mh4dYh0Aqvl8n71siJ1crA4w3rGdOgLqVLTOUSjG28VORW3wr+0Pu
Bq40dKEIiwYCkP9TvT2P/28RwdAcE/3K90zGBkPpManDYAkbMwVmPdndqczk4dmX
1GVfDDQx4B6uK8CE4GcvbKhYF5lVKPuNMcfhKyk21bnqnoX5ulde0FHXV5q69Yc+
8dTLc5ecBM36oFxcGSDufjAVViGZBkmGELemqd61QZ2DSCGGQyEYV2mlWL/4Dgl/
ktMrmLFs/23czN23y/Q9pY07q8DppnnyT/VYT0YQf6X8GPM9xUF4jFuwvSCPQ8TU
EbLcD2M6rX/KXgFaeNNKxAX2v10RAppJgZ0qy0iJMBBZVQHJHsEIdjzv7MHsMQWJ
4GHCKgnyz6yL2Jkh+VK7W6RMJ5xDrWjhd3rUQvNx6/Uipc76/hALp3KumTrgv0GK
L5QznHez2Q5a0QZDKgu9AiiryMsHqhOFtWKftDkXhdeB8nnSL3A08ug5/TiL/Hpz
J1TKgS70afTxs3t2vXMOLdHUrgL6EAJwL98Bcex3AKRYPooN24x3lY747kslhi8Z
Sz/O6qE314/wL5uzusrKpVkiIETUVTcrWJl0nU49H+WIrL4nIqBa9nD5BZRnnsdh
whsSCNrSo9oB3BLJVoImmAQfU1LZ2BgrJRArlUr6W83ym/9o6I3qvLjLps7BlcQ9
n86II2qfFwKYp+1XOPldcAvykrntWWQl0tc2SV8Hj+lwGKCzQHWEehX7YBSsJQvZ
nUR6P0RySXEDuvHl342vx8IkmqhHG6lYZ3fHEkmL+c6res1TZ/pIx9jkGAmIPYcM
faRybcPVtkCL9hVOpbVSWynAbasZn0iHzTUxgxFlMPJjMXeOFnwCgNJhdA3jH6dy
5okTJFvXwy1OkatT2USwzF7rUKDKNIwjXcPBYdduo777UvuNxTP1MdpyxW5EHtki
nVNTE1iXHM1tjk76MW4QCEVrb2vP3m9wCK4l2JtROHOVcbk4dyYwSn2lhaovnJ8x
Nd0SMcgk2yNt8SgGP6C6JwJgfFocYJQg1nF2YfNlwXZkvMdCetpAr8nMjRqyOdyi
R9vpue9BR+Fj4qMK0OVhyOjTjDvXF7l7ZdLGlNA7pk5X/8UzCa60yveHQZ6vJCPA
we7jeUxc4CCZjCS3kfqDgVH9PNzWbUxuNTBOnHK2IKvPQIVxmO09dzv3sF0ZWbKr
JJKVx3lni7z7ATQnyr8P1W7qlbq+U3dm19gRZqHCigrAndwW+YZ+gXKNKyAFCidX
9gbPd6WQmWTXouTNUJ99bEfkTk4eNbjCPQRm5/TV0090vbtTDZRwAlfshqDi6keB
txMUEGDUq49NFQBXY5yMitVG8ppdhydXTWMuhj8j3Wbv52qQlGvRiK01CR1SSt/S
SylIAMrRLOgZn3nXQxurTTvahBQj8fANCKTUHHPNAI84zkd6aFQKF8/T7f+1Ttk0
zmUUuyeY6C6QHWIMXYha9uQ2i5NQFZZ+JlFnk3TIYSjUZUypnp/pwSJrupnBgnB4
mXLrwfzWuPTcJT4pPqJzS71mHcuSAV50qQZjArSqoI7ovzxK8PkaYq4Voleu1OlG
Wh2DGiVBukZyQ+VC/+8zUbT7E2VDTzCXRviHeq7IvpfAzvyQVbnkr4tPnxmWxI8P
+BcPsuopA2KBIcdgOp3AgF4QEAgi51R+RP2/ikmpTAuIQww5wrO7tzVEwMvCEm9Q
umwfM/05X9wpewyLU65yC1FG8zMpig1hQBHuw3eIhsHOF1fUiaS5KgBPXfl+q6Gx
jA5CvIVRVuH1GGqf0JnD06JvFa2zdB6mPKWN/bHf3JeWg+t37GTG14AVMfxsS9Kh
fQU27DVyx7TzN4oPwm3U3FaOJ/vnYo1oJTuJS9oezbyIwMgsEGbHuYwNsnz1UGzZ
uCTn7MwK3QTRCo9Uf91X0xEmqgsFH+5+QxDscC3d1ZJKZamdvu2aEmbQWCBhbr6P
I8kC4dprHBrhxDGBw1tk/D4z7ZIY9XYS90wDmTh6cyWJaKFncVtvsjySzhqOBdjO
WRMrs4u6SYEqEoUngTDXUrolW8zIis7bbriVWbZI6tPXCGhHQB2H/iv1DL9O6I8s
tgKpdgyarq+5oUL1ExPuKPjjzk7+Fd/yZFF72CRwuKWseFd1dfxby7N7rFScwxaQ
DIllvwi+dNQtRdbjgx1iPdaiz7b/0Se3bud5hHkVCL3zwAETUTasnR/B6NHVGqMW
19A/mN3/T5EpFDxgWsubUTX1bEwWq8hHGxgV3Hj+xnEevTq4BUjs/GUkPOf7sFet
p3YSeiiLbBEXq70EUC2xkk0M5IAN2y2rjVqHi67jFPNwppWw1/iAfiRaUM4h/IVT
Rk7ZMHVkTKhkP/pp3AQCK8Juwm7n4WDo78rZ9WtohcmfJqALszTQCjjmo9aL20y7
fSOxOrHugzJz2wsNJHDQIm6fzjAf9eiMs27Lgkuj/FZHNy1kxGACol0xe55AJP8n
4cWXcoxeh9gis43mCzBxKrEuNw4XRGeXJbw/bKNsBuCTf9OCN7iIX1HAk/odA6OX
L8RBNoEXnMGu89IL7MtZHLkKYOe71tj4HjUpwgei1pP0q8pxlyT4g5zAMWc48mZi
dUgpBqLBH2GR+o/aq644BFZFY0YQT5YRIGq6TDIV8XmvoXs3Bpi02bJau9Q77dxR
McfijjtMjljYNlIhZ/plXT2R4SOQLQq/7ItYWZlML1IDfjWc9ot6E8N95huAe928
DIrISn2X/GoKGOmFoRLgZI59OAQ20MzNPL37Qv++dDGLfvKYj9qRrE/EvMJWswY7
AGM8hr730AwvNLNPd7QdDQ9mVE89SBp2q1TrhMc+HCoEYpqqc152ZPJiO8yB8gxF
PBaDCt7wIAlHpZm2HTQvohaYTDcQfuj9JrBhOFq6HoCUPqNdN1Arsk8oMe5ahTrm
NjSEnY+qrvfKwZEmH6fUzJ7DGZd11CdgAKi08OsK5I1LJGyisqdN+2fDnZW2Zwny
OUqZPBu8/E6+8+R5UsPHKU0cIDg4TcQuKcxSUooHCq7CIBiet/4e85RxxLHbrv0B
VjZdqYL+pVjhXMVqWH27Dr0kMuEAWA5x/2NWjpfYR5SuXH90fYRAKs/Px9O/mE+A
V1+KbjjAcjNtlH5eI1WFjJOS3ApCWo0Tms3TQXKq9WKrY6L/5oA7X52KD+qh0oue
OPn7pGxzmWlYO4VkGbPY1CWX/nSGsIN7d6xwv4fd/15t5bEHLWcdiVBid0LK5Cip
sezM38ryTJaCz/P7kyHryv2leZFzYwfd1eHP05hCAw5t2yqdFU6SORBQJTC3smHO
D6Jx3OjQk8YKEkFR3AsjmoxyAdnNQkC+ZAHHa9Avj9VJ08oxLAbW3JXkN+VzyAFW
X5uZlNQe+PIbrD75kfv+vAJcYx+nueG7k1+ZQaOdemNtf1ObNgG+mg1/JqEZHwb0
55w2a63y63wkF/w91DuzW6YRq22HEglPgura1NqqKmDbWHXyykzXEOhXV7VzgevW
8EIVGZYmpgmbl/7dh0CVD7LXUg1gBpAByqwKk1/YZ7G5YBc2FyuqKqJWO9RTQdAb
fciFcNi5L3bXoRzMUTj7dTgWfSpe8tKTcirA7HHccWBbnpnRiZe6xx4GGEA+bjTJ
lfv+zcttRgkDh5VC+pDKzbLEbMHAcjzhY6+Z+DxpxbAVrxelQG0qm7UfW9+vBXNi
oug62rLRbZfKnluC+sDTx3CxOElPxWpH6HFv3jwArm2ZzHKibc0Kfx7+yAxNA5vE
bNuOXFLDseNy0QOubfeLnTf/03ES84TutYKtMW+wz/RMOMRl73t//gH7pjqR0gpy
/rdDoLAQkEtiWc5/lh+dglvWUmB4Cwm9mgehSlf3eT4TmouM8SbWAn9igYI+RB0+
MPRMxAvLQqmC501o1qhzDemGDhBnlqI8QlkgAjfcDN3RQfpHhDa2C08U1J7OA5NP
u+3u/rnzYAuNse2yQaqq3Ct7vfO+yGYHg+B/9JJzp/IhwJoPkccAdGxgZa5ebuAu
3cix0jv0Nsb67PNbwqvr3JYruxIcLxlZnq7/sHSApkDGzRV8bwge0HG914xFirpn
rWvHT9R9ef7Yzfhg6CW1lgDs0sbb0ebRTgn7hTUsNFBDFxVVrUV0UhhnH/OHeEqB
W0h9Q6bhbDLAmSbIqTnvWbrBLKlIiwmgKt+lryLBLs5i0wtgVvy5Kb0A40hEbPuP
5GKdUtrslnPJ15nAQxSLjriHb7SCZ5hDoJq8dK1sQn3+NBUKr47t0ix4GcMLTjgw
Aatk56R9V4Nblyo3mnkw/2+phQ5j+ib56ddFz9E3K2JjPzCf51gQGCD9LCIGghUi
UjPJpmWTEEQhGdPopHvD24FmR5Hr4b9Dgp7haEh9jV9Fu2GcHOgkPljfJ+5szt0J
7Fto96Z+KxDaN+VqpBTDS3T9ENNyD5KkeV5LkPM6DgaVl9r0EpOq5V81Q4v/HFRu
Q6iGSyz3Sp2KaDP7NIFdU3sS+5XbEdyLgjt5lUFmeIwErWDr3Y/Kvi5X9ZEw7kTP
ezJpb8xf7MhFn/5OmkZykSRXshRjgquOpLzeNICnF8TAtPiQZh1PRflTs1xyo/Y8
+OqBwuj0hDbhvI2oIR808cOvaXHO2U/B1wChj4CeWo5fYhDan6oH84JJPs3OUNpq
lXa90su7dFYYMW1rTmGC129UqSOjcGbySWGUUZEWHpRBhBhZzBy2AkgYsKDSQ6CC
SNDe9bUk9ZZ+1b8KkXmLHb6hO/F24S1ZBeqtmsOn/pMtv3yhZHlZm7a6+CzDD8BA
GmAtOSjyvCBRi01z9ZU/pEvqmyyvtY23JKQzzMSz76OPvoF5ETo/X+uCIMzdSngx
3LXVB+Oa+LWejEYpNgqQHsryGv5/Atva9n79FMAkCUZ5vhcOGaWzZzmTjGIAqSTb
x52MlWDdMB51IY+hcFnVcFqUHQZlN1hK4KCy9xcbwoS9BpPRML8yxuDhSXdpGxZQ
QUoHZKFLgRZQJM30q5AntKrBrvqwA+/NuKHdgtkIRwEMqYC48HhRKJHVU9hnl2NJ
6Q3NbsjjrMV5BiSah1JIwz6QyeYfbwkwmUjhTaQzoq+y6TAofPt5idTKVBysXTfJ
A+tqRb+Ys8ZtWqEX1PuWso5cLOiSeA+alsgbjNh0uX7bayjsEU4WZq9P+Ur3cYpr
RiOXi/PvaecCkBlf+8beJFrgo56S2pJEHjtPl3hSPYzTv5F/4XegfNDBkiDAlXbJ
OpcC8K9IVoIwoBZtYppPQrEl2E8v75IZUrahGeiqvgB9YL9etHNA433qJyb7YuRh
TE4efWSWf2rHHEvFOcQkF59LHro/Rpyg4p/rlRq840SsbWX9SwrLrrYEetYOQ3lr
rAcanSG9XXdH5euXbNed003+wD4Y3l8wDUv3IT9LZXlcpZgoaRw9IKayhFTUeyj/
V/JDvuce6vLxZcHUiiVPv1M+RIVKb6gDtygm9QiNoyYnNjl4O9A4F8YoM28EluFA
`pragma protect end_protected
