// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:36:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pGQq0CGgbMKU/NH1PaO9pdVcz/mWqBZZIEYGcSn+NVfQZhXuTeD6MLmf/6UOBWlc
CpeKbaIZ0c4uL/3ZMQBaggcDrhO1VjebDCH3ALvQtuag1qWqR1RLKYfS6uRMBf7t
vVpuN0JB+XJ+qiF6D0+6wNF5kvdnNgZv0ktMI+SuY5c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29024)
03h/ytsJM26zjjTZkE59z6DXjpNqcna208JK4yZ15lUaiR8XiDV8WSY0unTMQTcM
yDNU0eX0StzUzKoDQnvkCcWo57K/9B8m1I21p8LKaISV83giv8EHUiy61xld9cxf
LVjhbqK2ty4gdhbCH8U6ioM53B4iK1w2kYPbTvUNCQUcxVCmP7iqjdibRDFQKb+z
Ftt9wmoD8h4TrHAAzdplRk3gKCP11Ra7YB+64xCJCntNlNCI3PW4DQlplrJiTM9D
jWJA6MV+P0Umik3+d4eUA0XxsJvD0uTigXIdimqK0ZnY45vLbsnjJF131htiYZiE
OJodLDWUBaA2y5uyrENC8NHtPIFnAWQ/mDxlU0eHC2siLRdEIfSx/yZwKveZEb+N
b+aGEFe5eIAk3qdH5LRCr76clgGwXkDJ/8onAEcsibVj1vSm/5458XhpEJv+Bh+J
yCMtguh/wavx0kMbo+oESDqUB4e3uGvtKG81El3/5JREib81HVnb4Q+nW9/tmJEN
TjgmGxxdMBX5/wmOskzdW0b8qn6a6u0Wc95eIEX/aS0FfsehRwrQBqxcKb7lwD+z
ChkVMBRNssFJE9uIQ4+zqYktNuyingvBpBfg9lFQU46FceWaNUKqRUjMie0AwA6I
yLctUuNB//9q61djkuRFvJcO85YW+maj/+MeECeFIGAKPfwvFlj4eDamMUXj/PU6
nm428lBhNH7GTYt5Q//SeV6pe9z3+e+3f/JhHwGStG+68BqcqpfvN6RYy/a3vcgY
QSKwkiq8ZskiKheHKp1QElaYFV+8Vy+EN5PsawYN813YPok+gEP6ZmKdtgKjNINw
v5IsszyVFnuQ4cv7g5hHx3IsZG3hCErwN1C/4A5OP4s4SHMiAPe4DcuNB8xRPLQO
kBYXMnzz+nxo6FA8NcOgKRwNqBYF0Gb8Aq9zDdO7YrV8mu7Cqi4GnmEelcjTqsCR
5okFeuxDI711/Jgqd+alm0jEWtoJxnB+/975ocAZxmUEluxhh2rIFPJgnDthIBPR
GCu+NAN7C9pABJyW3vvQIpwq6ufHEyN3vjAzT3twvyPqdwoxhW74ZIW2AKA6Trbu
qq3xXVIqWJikpaDdCqUc0DSn5b7Vsq0GeL2NG6c7A9rGl07Bw86Ve7shLOBJpiHk
C+/Bdj5YvmwV52q9FU9bK/gESm0+QPPzBBLEPBneX2IF9kulz0BxTkzvDtHL/562
wuZD/JYIYLU2DxzLnavXVBpK5AcZQKoJzlk/BdyqEw3Ql2rieUBW45HDts3qDNnh
ywLjKJkFM6iy4hF3FBajEU6HVvURQMI0QlOyWj1ve21fvwyCOvIKeeYp6Yz/N2tJ
uKdrppEXXueaXVrB+HSV9Y5vh5yCONVqv9PIIJv5bPnFnVG088/OEmFnYPtOW4HN
KHVUHz6FO2LHowP2QeDxVEZVNulhTqAS5HgVpGDvrpJE2u7sJtJVgghKWvzEWbso
sffTpAADLvcihZ+Gklehf5y0yUHs/qc+1b5teCaVbaxTazlWSa+yFa/RER6y6cII
Rku3qwstb4iklgT+DYdG+8iDJlIm9ffYhMqIr+xnsZTKRvjKU/Oo64Ab3l3+nP9Y
V3cLzA73Sed9i6TGR6tDNPWzH30SkBI3dKNpRlYxJc5cyz4McYQy/IWZrM5zd2u+
+/FVF80ZzLJ/cM3wcm67PW76eUeqsuPdKy05QjhOdDZ3KX55+pXHIt3YqYVFup8s
sXhyavMAUmghlekQC6FS72c3zuIvuBpJr+nUeEKIy+kRXLvKu5lRaFuplaZVHA2W
eDlOgMDj+itIJ4cLHleA/qTXfd6NjMxRZzfdo1MJMT7HQybtPoyMvfgQ2YuApp7G
q7r7LK7uTu+KztDrRvlFLKrPjyVY2QgeBx1cPH9qX2MVED/Z1vNnCMB7eSlOJ4F8
6Dz8NE/xULEo9VmpVWiSM7Fh8NF3IiKaMrRz511Rmyl/hXjoWKYfNU6X+Yx2TFAI
0DvF9fIMd8lc5GzMznYsGcP51k1r5k2ujk7Jwz9/xwxzhTDkrpoLt3aGnJBD4+tA
Rr6xtVhzWDKwaEwW++ZAPC8r8Bmrw82VBJIlAdXl9PsPfglDrLmXUa83fXblgX+5
8+oOwdGcO4fu2AHuGS1h8yYNqCxvHpiKZsZBjtSg0iPZ/xPPW0ZfRiu0uGvxJdrV
MxQ/6sSGAgn17YQJvf8HqCc7f9k2ciUAVfKbdQwZ6P0t3rjfmgjf5XhDjO879Ej9
dmega7VjNyvBNYN24piqrFwNNgNaQ+amJJhMaUgleeWQwxvPI0vqctRYmiu3Yggp
VzCFYeqfV3257UBRYll68HD9zqy8bSOyi6Eb9M8+/0cNSDQZi4+AsVCqI8R2aLrX
Fqr9dmCgF3b8n/pwL2C6zoVRjCXf3AFNVQFX7JCJ3IhZBHINUvaYd8c4161LktKP
PLHl54zxbPLM6XtGjmUtlDYuh026I2CWc/Uh7v5FVDYgNjnkcBY3KPjXhIzRwALk
cQRqLY815YlbgTFFXL4d6M9q5o9sBWdeKv/7U+NfCMti2h0igNLm365uW/Z+to30
vpa6uU7vWH67vBaPP0qSDJFW8A2OttE79OgCPz/KpN0gqd+pAVEfTbNaGQbgjFY3
rrY+l8gT8U3NqfWaZIy+MZZh0/I5TRJXmP9A3g5ORmjUtg9taFI/uaV6/MmoNBuV
KF2486sOyw2fQiWQ1TYPMFPbesxUNPwFL4u+pPFeCKxMYh0boe9lngG4UUs9AewB
vuzXmZff6/DRgxmhptSUWNPuw6CKOGZBewpLbI4IYIK6xrSvR1VUvezEptEv8dKD
y0rSma4XfTs1szcpdDuhEXdL7rbQgqsgM1vOiFSNnAwwKCQq8Zw0pJrGC0LWF5yG
ngm/bRwvmi6GPyEOsi7fVfyv2otnZVIu4H98SQa3XipSikJTxgWsiuSXtH95rT4J
JB7h1FDnLsiAml4puHIo+77uoMXo0dnbFw3UlpgGLQers/yDvw6pcwLjiF2fHxZ0
tD4GcVvE815qKJkFNyjgRKFPflS4H99VHxIFDij3/xLt2e3sClUAWcH3lvVAXVM/
8f6o2jBIP4B2mN+Y2GiHvN23YvwMaaYBkooTm3llW280JROmpnJwN+rvnWFBOkdk
S1LKc7tPAyLiO6tZyNLzs5RfuLPzmmoYhQdcwuhLK/eDXe2ttZNmo/zQspFAo1SI
EJd8pNTTtHLvfpXfJ09TB7Y1S4coA3mFeFAXQvZzeVuO93XVE7m5DEFeKAHYKZq+
xWMjofob2QYiqoPqajNpjTwCh8RrTm0lF3i6XJiILwyf151jA4T1e0chEwGKoogu
N20NOvddZrA6f6dVhv47TrlDuVZ6nFxRLKTu7/tAabGTPFLKYe2UlCbS4Kg0Shht
uoDMMl4n8PZjToP6DV+AgDS1MAd0QaD3cW1J7J5zutn8h7TYwnNSUxIV6V3kMSMm
Ik6qmi1DgTiKMIFGZt71FSZq7otsSQBx6XT3jFc8BJeoYSamsRfBhIbOKFsj9/66
I3IEpTtG8utWAAkoMV6vxDpaT50Po+15wNjS4LuiF/dhN/tXnxbb1bVnGV3gegP1
J6thFK6JpWYXdh+9isDyAXb1RzFV/eevOKsdhVd/brqp1eUPyB39rzcXmrekFqxv
fVyilSuF9ZA9LgZDRNVmWiGlobKvssQ+FXTT5dHKFox4HKPBmldW8KfNSD60CYf+
IqKBSpkpLOgRciNOTK9S1xWLko7TsShoSYuGgbQK8/GiUq3hoxxxYCkf70/bKFVB
Q1ivi7F8KCy1Rk/C7miD2SaYhLq+Q1b5voHG+DlN95dfUcqH5zuekrrzKIZz7eCu
hWYyLwD3opnEpIjPSrEt5jorqcAUP6Lt1GkeP1sOtNtxR1g8SYEcqgtDzatWfDbo
7sTAxbCTJg8NP2nuW77LNPxZVL1cZUJRknrKcdZVg2QlVnWu4bE3xI2bKi9+s/1d
JL4iYJ06AhaEQeHXHpzlroT0nrN5NrMSh/nWqu7lelimCS9zL9LLf/IFa6icH1uY
ez7JAsOSOilHGDKq9VCG1P2vJ93Mk40VO0PiK9GonrQtQM6pt6xcBGye8rR0MPed
ttU/H9VIbaH0Jsj0J+8fGjqw1uwbJSYKjvwWmD68G6PYY4A/MCkfEfdXbxQYc72E
XPAnbvDe2YSmkdCva8c/eiVQT8Lr/yhPObDFgFI+f1dHIaGUnhqeaAgbizSMIKsc
Yj3JcGc69lFcwQLtIYAa3L/8Txl6p2r7o94uNQS2jzay8PmKE8NL+PKfwMvDb2sq
sNHORCqURcXTL7IE/r/llIWg7sHRnGUm5+O1uaOX8kSck+1AeIoRv26piHKa+3pm
qUf9uqJBzxL1TF+ihwQtlIhdPlm/TVIQEgvGcGCkIUbEeBVoSPDdSivwDz1KLD8I
bSNkVi9oPQYuYKSzn/JcqYu1PpHILXHB4LsMJsMKRZyfdXMPfup1jgiGXIWoEcxg
njotgvz5a0l17ofjIdeB9A1IUD5Aimjrr1B1x0QAnf5i58JSPnFOcC4Pz0J94s/t
JpZevU6/ABWu0XapXaup6I5Y1FTN4cfwWkmBPVIz42loql67Je2vdhCi1pBkzj3A
duOg5W7uPpDmLeBKZvIn0JAjMzPpvW5YLEB4ACvBG2DapetpYr0RA5IGfiG2RftU
wu6T5bVoduyfwil4sIvSnHYZgWHB6xMPUrAy5bUw8pDiuO9ZyCUqbKaT8hTX9hSS
p/UUiVNhDJ7JDIQrnJfaFsZTCcmCTQgTGyl37YELfT2riILMZAf6uU9/oAKT9+Rf
1Xp1xJ/DEDLLf9XFx7lAaZdZsz1DTLDqS3u5mjvzMSULIFRS6IBNQiJxeMTs2NC2
hricEjplnOuHX4w0rbml0r7kZQSYWdDNGmQ1ldCis0/nMnC8EgONNLAh5ltJDQVX
zAMlb61NWPuMn0sUomZoe+EW1wJywMtOh3QCJznpi5Tg/lGmAS8S1xWY1a9Tdxgz
YIwi9DACwv1M9M3PDalGSqgUPuvY6lCQVTYueiafMi2+mt/xHPjN1endwAZdlLQS
hgFe66v1ftlYhbBDc/sAnMjq1DlpxCeD34KvaYB3QRO2I4+SqrGwZToyGCkAgBmU
JTD3bPcB6SqNxjp4qULcZVsZP0JNq3Hbwue5hl0CNS8rNmV1hltlljsM34No+J9r
wbiaVbwW6R65o4YJge+hIUkOmjGVInM6e5rzN1kwaT1uHwccDVEMx2Ne8jzhQfpV
86x6dPxBGvSli7z1sAbQUn2I29kWbYNyz3RrK8TMWUE5XIlk39hpnKdV/NE7coaY
RIyLoJdBP9UqY/K5o2wLbDG/R9D/iSMEWYkrztZZSWCWYqe4Ye/G4cs++sQuyxJk
XQI0fCi9AXIlGVlATUHScB6bfqS3nve+Dx42bBjkFDhMWG71uZnX67M7UxO5on+i
t67rj7PrhFKaSyDuuXXjNh7yciSR5UYywHVspCAOjyaXzUce7Toej/+7ie5KwXkM
27ra48YKLFz7I0RxnHMj/7Xhz9TDz7qIRBHIbNZPaLQggWVZhAR3kaA2Ys2jvWQ0
wIPOV3qkkDIu/OGsMgNKRCsVlCENJB+KXTCqQXXG1a5oa1wAcBOZlvlmCbM4l7h3
+xwhaBxNvPag2XCuyvFJjwDXD5uTdt1/Vby9/mWNX+E+PwSvFA9I+GyfQQQPBy4w
O0EJgTuxmGsLD9FHozXJg0Wl/JZEyzeol6tIfgP+Bs4/h4enwN0BjxcCnKPMY5ul
lSG/efU+g9MSZ5nyMBF1sbT21r3Pj2FZJd8bErBXKKoGhVldxoyRJg0QdDl6BbfG
ijQV7JpoxlGNbrT45wa3SQsZ2Wr/32yi9w3n3h5JgcruGR1NFUckier/NX+VqSNo
TVOo9Kl3cYVvUlew46UgYkVUUz1MZHYNBa2nhIiNdnU66wc7OSAlimWYOVmCh/yD
udjjjlrgUaahCLO/lR4TV+rqKBIkrfcGzLkEWHCipUAMuqdcm9fve7ZJhYU4RPSk
YATm4oj0zdWgv1V2yor3U/8ho+mYrEKyruRsAxUFEhKtz+W3kPaPh1R0bZfVSuDB
y3FfTAaG87C9fWBb5jfFolqjLfxoUzpgsdFMtTQfBWRWoODFz86PWSj3FK1tjOTq
694E0rbFubDqo9az9nLce8u8y1XT+Knlvnhz+5GBnCSgqhqp9JaQiLdygBHwoNUz
iSxPV4wa5V4MMx2VdpzXEEMsE8uReg3pysMaILKZcjfvM10IDp9w3JZKL7WrZkTT
9E75AL+NKpy2WG+zGHugYm7Pyd9Tq+wVqvEcfWWWimWNNqLfbWEzy/i78ahbUNgw
o+rLqh0tPD6CXmGQqnECYdtK3CCafgHGLSOUoZ8SyVB9FD5D4jkBaYNI3ybyPIIy
PTbJ9EHilHSG6MRuwL9Op3uYZ78iOCK6MBm9k/CHcGBzh30QkntNdsPbTYYXCoGF
mMlPMIL2nPUlAHkMLMxTgLOy5kS/IMv+fK8TCvQY1cVMMSEenSFMJzsMD44bDE4Y
UQOEuEpWSqet4pJsCRU+7gbg1srDt5F1FOb/XrcafXiu/PnHTRQyC/Uo9VwCMpld
olwu/monRJ2XBlL3tp/a9VD41TA+6Oh7n7DLhpwZLN2gUG26/mhEPIiRQ/V6al0v
IT8x7lBUG+4FjVDQO1UVWhp8OvGY3+wWxC7Xg1zpmDPIWIRt7waCXrxCmyqsZCep
cvogQa0Z+MROnEpDkF+SmJ+ET4EVzeYBj+j17GMXhZcCMbB1fU/CNsuoNrfRya5G
nfoNVM2cFKEVctyT8fp9y5tWew1fFfw8W+zIW3L4SL2JbZC5qvd6urQKmxBTNXMB
PPQdJuHmJTR0si6rRY7O0N20VcL0ILQ8slD13GyE1pOtRLI4/X0mWPI0vAUQZfLw
JFCSAlc4L5dv2Vn5voC8UBnLyfxBjH/9qbqPIQ8lGfSYE5nV+7QvlZ/sCHcfmesm
Ku1udFLXkfRuX4PZf1jzQIOzFdtaUeS121vuABAQJ6h6ztG5DdkRnC0o0LvfWx13
SF3IcfCPMtS/tronG8wIOiDphUNAyibnULzIdAcfH7xM1f9LkaCu7xZUKJcPnSe6
qWNxyZYFFK3GX4CPAJJ+01P+/wdhYlsx5AaOv1VmfisbhDmGrNGdYkUQTe3t7zS0
Miv2okSCvpPPK+dX1E28KlB0+9EUaF6IkHtjYu9KC64NJgxSKuOKyBsQ45F2pBPo
daimrb1I3DZm50Tiv+TtFAS2PVreIZ3RBJ5dFqUqD3V0ZE4TijUF1Y42fgwVGEUP
SpCOrpXpb5FJ0la1bpE+5QADLpjOWoP0QcSCEGHBhR7w2oCugyssvKPJhfgMt0aK
yh5gLCj9wsoWoHpfgj5C4Ztiq83TI6ifZZSn3cP3eZ23zdzJ8qnnsr7VMAlhPPF0
RHU1/GZp6xZgM0mdrbxpBiwxEW9+RtOJGDAncidd1ke7IZhbJBKmzD7DnJaxZzap
HpI9BzanBMogLi6RZ/RF181Fnzv1FHXYG7lMw3ycILx4L3vhpW103PDVInBhBzj9
Pz2X2tPHQKbVnG0wt/B3MHuaOzMcReIQo2kTPXLS82+AxiK3dDWPy/ga2cx9aAnk
ZEXpEYPWw2eBKzvVDDCFAJU2nQjQIAw/xakHQhLV+rEZkHDiEBw2+PgtJ+DGAIrm
ciE7wrVRnUH/oFIeAViSJNBcCv4gVpkodUo7w0vmboMsX4QL5mS5miEtDEkDGhQH
xfIepxA8jwBvvDP8FJj/iJ1idOeCT7wehZSq9Y/1ub0KLG9RIvKQrYzu6KDuTtMc
PZjUciLiimayvhFa7gEfsCDuH7gY6jlptOhCPyizvk+d/k0h49M+6uBQBGXyB3rR
MSbXOtSpzW6Ks3x00MvQUtiroiYvwiX3iCN5xmHLG10I0RKzS4o+JZvJpZtD5+Ze
8UFiIo9Or9OBchGJK8QoiPaAYoTxNX8SXfH6nuk9XnkSAIcpNTUmlnV1uQbDztjJ
hGcR6202I+3SCk8iGuM27qRoYfAcrZ2AU1/CYzppV7Iws74silt5anicc3tgPXfm
VHKmvIeRPzQlFt6V3F9abIndCGXNx/KE6dcqkw+dgf1PVFHjb85od+8BXgaYb8Am
LpazEfxAU8xsth+Ks+FuQ0JXrUYzl2SHsI4VDExfE/RfqbL8qgq6bSXMNHkAQI/c
BigPvdshkR0nYKJ5xKctZpW3YhTjpofN5Anp91U1JaQUxrmI8zah1JV9Aik5toLG
Hm7R0sRaLfDrzscWWW1lF7zFmoUw3Vd1TZxxd/q41kquw0/A63wbkYGZDZdp84T4
cEQN1M+KOQMfre4N94G0lYgtRHMd+L4KaTGvVZ7FkUZ9ZS5Wwk640E9o3MwFi+q9
2pGE/wDmtZpmjX8HWwB7VSvoEZ7kC+Wv9y6Vh4IgoiJ+Q9lvKXSQ19Nj8Br/bdqB
dXW1pzcqN7bkQ6kmEqmXGnhFY96IyoBeIjA8ufB6NsoJDWoapRrZ0vp5D0YT72UW
LcDr1cQvZsc+EJ6cgzRNMLYxVJQdMlhEqX6GaipLOvWoGmcYA8BLMZTw+hQNKmT+
R07UXcj+eXpBdRMiXcUwmGUGDgt0FnmxRhE6o3e8JcddUhrZNj9AQBmj1hm0gOzl
askhsTosH16jY/mVz6Ad1A8TacK48yoqjVD905HZE2RVPB32JQxBHzIzySCHjmNN
0CG4M9fIVX6LYe6viX90u1VlsXG0oYzdUyoFmQez2iUPbDrdsO1R1PnbnDb/KpGI
AbyULQamI9zhMZO4Akjc3ltNiqLdPztAtxOn0Op3fsS6v6y4qu6X4KtZMpNhZpjB
XrzAuMJIlWP01jSU9jQ4M4nX2P1QQdfJDyhgmU6OX4ncrFm2auf6G9rP499PoUFf
x03CO4RUGiUU6uaGdgyWXoy3Gv4ZX85yCyKWpgyeBj8/WreVYfpm73cfKBrSirXY
szyKAnipheugbojntjzxCtUXtsGJO1E42ZNp14tGO73y74mGf69pz+HqganyPToQ
oyium28CuiyRMKfwchUamjkQqI1v2H3kZ4TSrlPlJOgM/8HpfZUyMykJqTBQRqnV
IiJc7iczM8eyZv9bIsBQYYuONZN/C3YjBkBWMspucdoRbtKV/wnz/CD2UD2JRoiQ
Vk+aM6Kth5ey18IulLAjU1Nz+DfaEl8T5nrQLrMei/Ej++9NC/A2xOuL0GeEml8U
F2kgEzdkU3if8mbIKVFWJeDTayOKcjrug9eJRA2BI/C7ben5u/AhrITC7el2MSGK
bwjF4tyDdNSi/pbGIWObP2k19fUaDJfXpDSJ4YYljJC1f3qyxoG/QBSTRapK7/Ir
6AJYnipKyRzORqU5o/oB0MWO8F9q9piQDLYN/lu5auGi6hxXuetD3GH4cqgHwb/C
It9vVIdGX8b+Alf/p6NWU8KnfWZ2/XtYURh1HEgBU1hshqEYMKofYDpTm1vCHPWF
yirsHh03HBBpPANAiiZjWAdElu01VFWatubH46x4OkExM6Nu5OPMSg7TPajW4bCz
SGkew1EGQGNOlSCs7wXDST7/BUVfxgMA4IjuFZwurQxM9KUsqwf3ZZaWYA7NsQuQ
AsEv+l9cfRc81DquhPvinGkgrWwct2bYavr0Y70B3EavztlmDqpnj6c9+wlvc4Db
3+hocYVrtI97/YORImkUWjcEYztoyzoCJYWor+Q03OCuIDsoMXRDhBsrMPQNJgTF
/73mJ2hMoShqq2WJqmM0Sh31qS/hY6tRFwe2o6g9xo7qDmdppBbO3RuIIOOPgwBk
+EwmY3BJaDRRFBcygfNvjGihUMyxbILGTQzM8gtwO3WHR6ZBzfva+rpZRSRL5A9t
MDhOiHI0FTjQXMf4Gqf2vCUDAuQ7KrQlsxoyexsgZcnK0nFad9w1L3oCVBUGs+gC
38YGlkfNqxjHcb4vTSn7D96UOZ/VlfVskRvsWddFUWi14sB57NOtD7QCF7EMYXSK
FJaFv4UwmmZmiKW6HcF9SuRBNmJimKh6867MIB+h/R0G8NsxY7twsQd1zrJqRGD3
kNvpI9freWJMbidJ1/TcWeodB6nI6ejFSc+itIJh3gghdjikARj7t3JOGrUR6IDT
8WxYWTXh48eVyjCU/l8RpxHaWxVSIvj5dcczDwlOneAw04ekqCMQQfyn06lNalLP
zA1FinIw0GzQOZhwOgzLbr0O88pCORuABe15VgiJHTg+1pHM2G3w8wxMaCidzIC8
GScMPuYLcOwhDogOy/9Gn2lcrxeswAUKCRo8ZdMIrVOyAcPTpA452T0X18YHjmUk
B3pQW62Sm4wgIEdB5lC5XfqkBgx7tqPPcM2f9MW+CrJ2FRt5kFx7kB9Kkhy6To5R
ExvrFmAlhU0nLSTm4qkuiNEvib5dS1VM1Ikl245X0G3UQnbt9mmOTE6Gyiqqp8Np
iNlBnNyWP28vq4okqJGRkzOd30vd4/G12yA5vbCwKRSdU+jDHHun/hUH5Mb2Dcx5
iyoC5FWOBo2jAzAOzFiOQ1dFy/BNDgaw3deoc9FfZ03MOmGPjzBJqSDl2J4Cx2TE
9yVvmihDAis1G26/hQ37yPMbhIDbGe6q1oMJn+SP2n7lBcjsjp9iYZQbZLvP58h9
DkiQc49FoF3ZgRPhQo7Wk+ZE4ZiW608rE5XXjIyDzxdx7NBXFSRt9vLw7peTAobi
g/M2UKLBGsV3BD3XZV1XiahsHTLh9I8BtldULihnS5JdbmJDpaaINtiDbTNnJuX4
n+51VwuDeU9RMjsnysZqkh5ruxpRcWv/SCPYh/viIShAO8y6DiyKpwPsI54OibE2
TSRCW01FWbo0uM8tgTqTZKW3BRFNQcBu3CTfXJxRpXNkbUT1wJkjYdIa2dnBwqlC
eWcQsEBbdwpcj4+yNwdIQQFjvC73YVAQBcaenWY88ejjed3fkIEF6ZSZVNeim1uT
P7pxom53joIzqqIBQiI0Dw380JwPfh8ZEQM7VklL8jxGvLoBAZfVQ6nDQQRPqcSf
aWvbWUJRchuKHpCJD91vFhEK20m/OYAOhggmbrNmMaDIffI/SCqCvPPQgWTgO6NT
YsAdm46O3xzBfNjToE7jfpJpKbX00ZyvqYHucLIn53DXhdwG8fX54p2oV2MSiPas
fq1BX50Cf8alqCRbZfEIYKWtKcxMumJiBoIBrT3KsH2RekXq0FNB2DpTM8GZybpU
h4rh4cGS3pIh4h+2XmGrtaY4L9/EDQgdzM2k5DLhofybFdI1A5fWheu1LV0yZs1i
z3msxyfroyNKeP4sHdIzhSMST6IGJUUt0xYZb3oyZ0Lkfylpg60Cm247xfsYkSEe
xCAkXVIizyZ3j1zjANBp7nBVqKiLJvX+TMwJFnWZrtSgdMUS4MOvGcPWy4QPENz7
kvTbuyVlVPG5+cNjJV27KXbDvmxX8n08vwrowCVonacERnnmy4YFFPUu78eH4pEz
209Ag4uwdjcvYzfAaybHPjHFt9aPHONgpYoWj1fDSmNCRynn+d/kxRx+yWdxxLqT
g/fMV2zP7H2oh379cAibwpUfQ+fHxvq5rw9ZRdHFLZ8UXJtdsVOM6EFfNk1PRQGg
WTiF+MmxEcS+zO4gm5eJUzb1QsoWeLk419TWAK4HIsGy2Tu9jfrBLCyNoOiXgKyX
Xm8VWUigXnhQWIKCOlGKJbTVyDr6vJGifz8HSFDloNLd52DwQWunl9wPiunukKNC
OZ4lFcnxF7nkQZSxI87aFUioKScYthzMCKJ4IDMdfqdzFupS94TqMxZLg4e6XsNO
YQMVvgCb8pnA4s6YgP9InTAi/f6UVBMpJnFaOHd7HNteP6Xop4rqJ2OCLy5TY5yD
R7KJNhfRjznuQ1Jwuh0997wf4tuLnlnQixs3FnOG4bksrxxo9JcmpdVcUpwjaEGL
QWBRwB12tmMFlfU51neLKVQ3KTsTFmC6a5Yzn5YLokBzjdgffvPzZpdAdTriD3XZ
Pp+QUHFrHdrcyZuaa1vd+gDT1ntO1u3QneZQKgzR/UB/uknP/TkdtK2wWtkDrwOf
iY2bFaGTPcA6uGumGUOQGWvcwMBrr5RKneFwsd4s6KaHfEqh/fmKVa+k7ndezBYt
w6lavI+ZHnJ52YZMu5Z71M0ckBzGLIaAfMdsI25V1iWqJQLyD8gk25k0Ka1DAQJu
nXH8h4S9N16sp+2j8R8Ev/Tmxp0RfhCtbu6TLkpwjRnE+Pw/UwrTRHVIBS32hdnh
KC401GWhQdJGF9ZhREvtztnKOkyqaQ27kW3vuEmTgazDc0VDYNjNEx7vwejjea0H
VSB53O19XdIsk7INkZUt7jvCQGtPb7BtVSpAwL5ViIbF2HBrD+N0DbybcAlcXtwW
gNiEhNuSydeCTfjNC/mfQ0wUs/jJkgI1GRhgdbVUOU4lus654Ctt7ng6JdZTUkso
uvqsFdvqRy7I2DaIQDz2gaH1L+5u9BszposmAKNa4F9KjOZm7xQ2UjQoWbBQjIaL
RHZogB+N9eLCvKxEpPC5MQUAZ/9AJnu7XIIFGBGolV/WfWAYMhoVDCiXKwKG3xwU
gLmgFrHeQGJk1K5+6Z0tOT2dI7xbRUGRy4kPHJr9sYxdtCfJe86ZAsRAZa2Mr6mY
vAa+x0Igeo5ts0IjqKDQ0u+1fnELIqarbCv5PshwvT+PVbaVUL+IXGVvaAXSQWmi
6xBVwaYXlMHm95sWJgArOyXDxk00bc8E0PLf28ir4i7ku4LzT5CFxod1fXlRWkYO
jxQoOTJQA1Nhivzu/0VV+mSRHqITMsJX69yk/T60EG9qn3llb6GyJgrkkS3F65hm
4ltJmEc3unKCwy5dN4pUUIeS6dFgHoH6jsij0rDT9S51a6UPxx2mzoc1TxNHqrQi
14E6KQTCaH6ls5JCgzQ372bqOCofUiuHYqB4/W8EOwe+NAoNiA6dOxQO1Y4I5rcx
Vnw2CuZYEqtes1EvZCgb2meUPtNpnV6NKqesfqem/LXZ6ma3cj3Z5sxsZBEV+NaZ
tDpQ+AglJ9qt6pNTcyQaHSH6QRYDpiZsIBId2Js1kBZp6TuK5z+F6n625B+CHDKC
5q8+I3FFEEMR6AjujUMnAWAFo8ArW41yD6npiSjOgK8xQfMOYNohF6ir5vduBWcK
O9Sg1CP6XtotcSm8EV6KZqnpIxJTVNn0TMaupxwVv4Nia1+ZWqeq9TYVL8rojEzr
d4SkBOMhl14fTk/YzzaU2NkVA3GpLoEu3kKRTFjVNbvt/419r7Evbo7YgvZ9WY0f
wRt6cxv4osY3UtV6JWkkeLcuaVboDqjq9DVCG9ZGwWovcKhyxbve4XwUxZ3grF3w
7IMlSeD3zeINLyGbC6FfYFDEyIUbh818xNbNlwDi1WfwWjq6dja23GYBuyUCXL8p
oyLEej7fiN4P9ySihBcv2qQjcxIdON9sFCFBZXppWYQPnIf0Ql6kSbZu/oizj5Sy
vcRe5zmlALaP4IkbfigsGuISItL/KERTxzRKdzsoqwZbE3GOBquiJAsWtgPjgg6A
nc+dTVHqSFhYaLvv+pketrUJuTqrOvSulAn71dgIelMW1mIuZ8QGzjfvQu8eTYwq
2KEeF917/QDz4axoyTD4CpMV5nSMakcL/6SOC6gJNYQt6JB39X8Z1/DtbqmCyu0o
znrk4yfSRI7o1twomUQnyWhtxSlXE6R0c6UnqT/1ZWY+3tMKNBVFNh0AzK4dzGTs
dIi1ck84Ct1QpKqP2Es4C/xXaa+w3DOvg61FPYnt1YE9YnJISdwo81mI4QPew6AG
4GKnQe5LkllwFmIgac9anZcyUdffT4MZ7KcHukFUTOBla1MJZPsvATQE5Z8a7eCA
Tt7ZmgOghkAWqUEH/G60kT04o9cjs8xR+X9gtxNf3Kj7rl/Cmg0VG8sq/r4HpHwU
xhqftIKQ4iKoRqTDymSEjI4ns415bfYAN9QhsEtSma7fC0w2k6QbABByB9O11uWX
D0Pm/nURGdHickN7mN2hxD2Fc+bBaianMVPInBoumIpCKJ5uVHWBkNUKc1q4ZAcu
3bqgv9VopNQcwpm6igKfhjIKQ9f1sigVdCWmbSMHXgkXlJlwylJNohLK9Is0eUJt
hxKJfs4N3FALolHxVWIvwlB93K98UaiaN5geDzx2i8w14usDEs5rMz6fezLCeVqY
hbvtjoA29LSyfQcBeRVhVPpxt6e/EXdW2i1XNJbCtdpTXKNSYUpRopw9Yv5hQMRb
d1q292d+35l0DHKGhtAefveJoxCoY4nnvxLQowUPCw+pGwj0GaEJIqC1ClOY54CE
oyu+kra8L2JMJvZJ7i9fqf2gc6UvFnftjmQpJbC0wqx7F+S63PkEPWulM0MlHw51
mhxwiJQPU8WqDZnrYymbJuezGc25Eq/khCHpUfvPbBzm/vql/+AT7UNQdXuQTbK/
zrQCASTAD5haHljvcV5ivFOHSdc2fEAgNDZfk7PD2QoCq+iT38dwUJRnL/oEd2fY
lV3zUckkqRsuvRC0JorCUTp4UUpoGnbbFanRLhGPtYa7tUOdunz4E930esjerytS
opnuD/7BXKvovVPQk3IqN8ZMHz2HNMDm/LUeQv7yHItqUclbjxIPGR/yzUsF8fUF
Jx4XUyTv8LAsrWfWB0QxsW6aaW/Rj7TFvpID4rRL/b6+eGm9I3lHNDqHpkrtPx2g
8/R2qKYfRmjzZ3peQNN/S1ifHxIgbqfxG/F9cS6ie4yTE3tK0IPSELWV99mUVqp7
ZMshm2r9SkUeJ4WMWh9UTP3Fn6ZPiZbtldHLeL+qmYfLGW0sj0KusyAnZVa2Di4X
lRp6cRr28wIFKiIHv43Us9hF6OAPsWfXGmVhNj6elfrrTeElRi+D1q3wFi6GXPpc
SOXfipr/o5fXfg4aAmdxpbEoLSf4kI0Bd9Ywz6CwfZ7IjkhwCOhUkBe5nMvVdwXn
D8TCfZJz1RMe3O0Z5fG0Jm7cp5GkvfT8LHwJIWEVb1T19uyTPa2QyY1knnptTLER
ms80wOGhq7mlPBpwZq7bxTY09EfESD6c0FxYgy7nGCsPpBLtGvm55RrEQUhLWICu
BVxzjeATQ+04uJVJ7cQnHTaHRM+wof8bF78O3PIdK/52eO0m88sKwUv/VJAh6TMC
tZfqc5aXC/69YqjYXKPyoxoHqJIbdl26G0UnY6VfNL6RohWnglbjzLByK3LSfLcP
Kkc9uHR+0pdwJbWHytNRt8OwlMytR12sxOeLqRIFYBAxg0b+ZHEBca41kE5RoybZ
xd7if6KJuDCN09BTsSv00PaZC6KuFZmg1YeW0xoDtSZ2Ka5eo0kKhqp2glc9Ds4Y
Ghl+XEwP6J8DdwVa8DPRD9ZdifVgVEhEiD3+nvfsBHD7J72oy+++/DA7Fq0lOLdj
WAUdvrjA47AHQxs9ybAOgoWkm7pSuD0Xjm3CT4G1FBhogo7fj9RMKk/TW0AvWCA+
zOQywLGR2kv9YNm/AiFJ+ul4PMoO5pVsxbMy8WLjcWqeV0e7E9pr8Db3J3QHp0fV
sMbMFmhjUDbFkHvrVcdHsl16UX87k8AgR3awOLFw5x5hH15xWIF1hY0auQ1W7p7Q
EA56/TlSVHHzMDTRu6tKGhDnl9dBwFq2mTm4LHmK/wd4wfZo9WQXI98m9s0cbuHP
NOUL2cX2kJGVpkf/4uSPVDFsNSY2XgPaWni+UTLG9/fEaSu7cWlUnxcygUf+8eG4
ZY2Y/TOo4zuGN51MhiL/K0f3SqxGLLond8KsH3ZtUXQ0dfBk7mkD6EyCk/kJUL8N
p3LqK2+7A4eGBVLdsdgR229dTCGSUMLaUslciJ5x2LUY0R0ukbkqGf6xQhKm9BU8
/QwdFvSdgwqT+XQQGWC1CXb93vZEAb+Y4/TpXx39qNp6qdr8U/zXKoeDqWcW7H72
x4KHTeNHi50aNY74r2N57ZeJ1zv+1bHXbbLvhicWb1GuN4LqX7uyd1GmW8dB48TI
OdPvrM/36aa3RwH+whqG4oAQnb1zUOH/nH83IH7P9l46ZYreOe2LGoxd0W7m+nsc
7QZ/54rFGD/f5TgqEPyoIGvHtOSSVPHBuvDGSgdJr8349hgrgd+rs+voOG+YcpEa
7QMv9auKSYbcMuLIdnLsbUEvrJf2S/GX5ejBlpwb2B8wn8pC6NHQ1GBEXayLldxn
p2HF5LP7CjX5PKWjheIxRE9tWB8Q+X8XpCSy7QQQjORjC/pfW8mpcrtgDQYugo3a
WAc1I9Pvy6CLhZz+hStD7AjMwB6766WW/k2ilJ1Sudc11KpMSOGIJalhCuMcRLAb
hx9GpwXt5VeQRDF6OVAQQefnmjOF/eyHgExmuMKIdv/zmDjdO1umZwnGL9x5UQnr
uk1QK6jI9OuX1JpOIP1QKOwH5VERSqgLL7bfa7HU7xmymBnUrcU/fRQErWrRyUjZ
AlXdslpjA6Wd3NsTdEaQ4q/g0eP1raNPbmysNism7ByjwB25cPx1+qsmeXGGKQhy
h0MUesottgdxY1q0VU9ZDaMAlKTwc3SQAUJvVKvX8pyG8quNECIinoqzQCOy7XFm
ubRgmAvonXaPw2IbujWd8ZuKuslLc5APAZHlYrnAHi9GT+E5SVl/MDzMCD2eZFEP
hrwGJMiMg+Uhc0CrKAu6KG4cVY6196v5fzExcTEXsCgNee/puAyyfb8UMqnenCzP
dhJkmJcGbmTFuqEQVz17Yaq6H4J00Aup08EMte/C+UiHjBL99QdNu0o8cootOUrt
yBFQCNMAXrK1IURgNmfOzFzY7TAULH5YQyjZspaLO8+bsd5LNnVE8VUR+vlMatVc
TYftbORtK/pNNn5zgYyNo70dcKmfyj4lt6VVRN7gLAXwbHq/nQXUa3tzyjmURAd8
uaX3sAXSw7NlCdLIVq+/KsanWW8lzfRdZOVlc74cFIUk1Hi73lHuvVQJ1wXr+KdO
FltbI2rrJpq6nmjCVnKozbWQ447ut/OuNIgAN2UIOQLN9jRsiE6D89dSPSJWOxxI
4L0kbaAnSULu88pMDliBglbfoOrsCmcJ3iiobzlMS2egjO+gCXonu4zQUxFQpflb
JyfX3BdHYMQZ0GEjGyiuGakbcHmOc/mWMlQm244F+2UiyTaykRxCW/Y0+CcbJWHs
TXrcxk9sTKJRB4q6al0t/KjAUb/eL/TNPg7LikHwHoSu0pW7gjkuRSKshGLz2KN6
T+nyUVRtjqoRNEbWk6NPZCPMK56rTXXpPoKWBycrDftHdd1/VLjNccD2r0RUcgnX
ss2DFJ+Yj06P5lspJAfxMc4m4qMhETI/0h/b3fkeqf/gSyW+7P6kVi16uH8N4dRB
b/g4xNB1sYxo7m9o7dwTd1Yqisgh/IDE1LImUW5uK6Ph0cRr4lTbCACi1T4i15dl
IckxgYP+WtNQ3uDPcSRbjMAlpQP2UEwYQAF14o4tZBVhcwvKC1nGTEF11nS0oQMS
lg/zPdNQ6S1LtQ7Iy0k8pwD9qjMuP1vAKtzixcBXRaRNsh6eZSjFCjrMEzfB+nA1
jW5ce2smhWOC+y9Y0BlyQ3OPzMbIXlrM1qlamsnfgsFFvVP1TFUekr3IEuU0FT9E
CRGhPNPQR7G3F3cu3XgSeT0BhPe+rTB9Z/yFNPtlWxT2gY3cGPe2NaClWDxI1h+F
CaL1bvg6UIjXr0bpaSL+htO/aryF/n9dS6r3dn4UOR/lr85kCiOHI++/sDEhp2Ub
HK9VPvJewghHS7kEnOIE7ip8kqj689glkkdt8sG9vtZOysGtMJIPrcc/X6Rd6Xdl
b0na8y1vzkBqqv1rzyHuGcndv2rB2mlhQ7tIg0n8ZpIaC4leblsr0b61hTrv15RP
p7/GAXZHj4FVekka9edwqzK9O4LtFa5hdgpuyUxOH8Pknuv92Atmu3hQVhvHYBzi
zJMhNgetKOq0ahhotRKHNb63jLH1soTV1tE28EjxhjZ1iLcSom3PTni+91Gy9HMM
rUY32whgSpF2homc6+aIYGufpxLCqe4s6Uw+WODyS5cb+HFRaRTPBvTOdaVKX9gM
w9b8q/j7J4MQjV+A0qP+hyztsjFnxiYrsMDJwigm9zNDgU5G7mejoLaGPt5qakIy
M3vHpfRgyAp/cIQ9FelNGrWTz6LbLYeqgE5Wqo1GDAVzWqMPqGAxdFfWqdueIXPo
PbGaHvD2pkrqTFz0cQIAv3m6GtxK09qGG9dNbSsQ6mG0JdTJ3BX9DeTpGCLeyFoy
5k7bN8NZjccaQxCkERqv2x6gN7hRSRlMC5lv3lqZHjzy0jbIpjHYlkV4zyDHX4Ww
uT0qPbUQJ5sFOlHFJ+13n9QvnTunCzajM8KrFW/LwOljMw8CX95sGvNEbxBlLanG
kviMDP2F6/9XqqDB0aZTzCVp/yjMSnmF17MYS4+CAyUUycNOYblpcUkMW9ddEYlD
fVuw501Hx5CwTgIcOcP0jXDuZbblpfcJ9Lty166Wjo0PJeGILgiqzh71YcOzY+jz
BYgm70oIxFdRua+yjjkDbz5DOsADUksRqM8Zj1ALJS2Ouyru3OdW82nLTuw/Dr0T
b6ixdbtFGADELYUO8veU4Ip7Yw1v4ma4hiUGquMTtwSp0ME3P9pEhOYk8rOVlSBq
VUthMLVyvbhBumfso3Fr7MGkzW5L1cgzLdR3L3g+5k35ziP4PXDjNZUf5lIRJNar
D7UVq6YAAuji67VkuhbsbsqcJOV91B1NFEdoQn7ZSTevFtS49pGE1vIL6vOCCJW8
nCvdrV5yz9gRKqiZq09FM2G+F4l1kp81jz6bHgR3xT50TilhwxHRgcTJF1+3lt3M
lj2fxrFh0ufMoc3FX/BjzzHviX7LWPs2PuAIhRLQG/uz1B1u/C4T7g73W8UQvtN+
Mi7WjDUPAGxTorhizpOwo1c7x9t9S5vHOrb6kjexd/aGJuwkgUrSnIdrr19V3DwA
+2kzbRWhAu+rtKzNxDVP0X5RPHETguTR6aMiw6TcQIpy7OPAI/i0KwtqIWZkVWRa
ZuPnMPILqbZGtmVGqjHzpvk78eXTWHljXtxp7OwA2cdkule7AuC4i4+73OUd/kVx
TRrTa/7uIVK25yy/Nv/WDNN/+Kl8rpiLxSA7f51i4jQRelJr1uO4ohqt2aGiHfRn
ND9JyxKx5yrH8NryZOpw1bHAkQZifP+cYoJe0GhjZ+VivtiAs+zpet6J7UKdX2w8
vVEVxv7F8njFI51gu7Y4YO7Wle6qcgc/U5lLcvoyWWfz+VF4Gz+pj1NLAQfAVpoh
KkHes10U+nhEeATvELcp5XR85SAyLZnr7IEY1hltGuzRiygtio1QuU6Nu8Dzt8WP
lQoTbvP035s2tMtvDGCN0ni77xUIKYO2PVqyUsXINL47C1xDWPeETX7FdPXiGoeK
F5BBhml7YZlx7tWOEkfn78f7lM3x9MMfZ4xGPs4IJgPrIzP+qvBAhd4n4ppMCpbv
o8Jnw5RZHIUFYzWjisAcrWpb2NRrYwVqRCy7FClHC5p1lHintrnrQ9pawh8fZPkk
QPRpn027vIR4KPG3vS3lF1WcqL4SBfOa7s8PqeIRKvbIAKf+b4JDfaBDW7gYJSYw
q5FfTPRn86Sl3sRYKKg3ptgUy54Ae98+8sZ+xFr5DYrEyurf+T+5m7C+e9xRms+r
RrVVhjuunuU8WaN277GKUmyHXRNoJI/5cQ+SAzbg6vBpxZFzco1Vk4KD9FcP4SWU
vDdwaGwmr1XT8d6kaNrgGofBlsNun4C0bRb7iQl10eeWOdL1t4XliPfDO+zATVq1
ZRjB6YYMOmpOTROgNy4pf/z9YkhR+RejUAXXx8zBha7N09bETf1ZPe1knvIWZVkh
6Ib6AGtLxVhp86LY439m1edEh/8BPZuYUX3s1I29/fzfLLFT+rq+H/XBaHroGkRu
sNWM2oe7pcJzaSYjTZ4m+YHdnGXyWNx5BFH+3IAtWiuZlXxEZP0ggvuJO8FN1eSV
Lo/jhhfLpMA30BkXxLC8OUMkWH4uAi7upHd9lwcEcsUO3/PfuTKVm5tedW2MJ7S/
bJtwlCYvyIqIbErfOgUuKfj+NRI3beBo3HDqSXT3pvnHUtdQcyON4fKZdvy+AyRR
JPT1xy8VPRjlhn/bk6pZgJr7k6SBXAeSYeYWXo7GSA2m8sdsbfyGDhs8p5fqK1ZY
OjQwpzkzVGrHFSHLyJJi7DZpPBO3/DmNJIjJyjo+hQXEOE7lM2AsKXHAbo5c+RP+
f70JoFu//pOyTzSkbu/+bt8NuQPcdA9ulXZzSjNaqprq2xQ3Yeree/nf4aM/oIr1
dWkksIm/h/iQalw6NFmuCBsu5L2nyHBobNT0y7qQhOOWqZnvsqiQdUmYcLUvh6NW
uFGM/0bVRCaB+Se1EaZTCac8vrAgeOwT/sArHrlF+pv8UFTCbwDK0EFvcEUUXBV8
al6KKj+TqIr2407t43nISLmxSyMCSIdas7vvEs7N1f4I7g9AOjRC1t+Gl9KO2EKS
Fq3NSvwiWSoFloSFBAKrvqb1ZHJcMh3wyLXRCODXBLfZky5rrfAQ3Tz1aR2vY6K3
FbZcqOoCm1zsVHAb1x2QPSBdepNsfEenbjmiReamRIPw31HeMf3dN9Hf45srlMhp
bBtOwxB54XLhSH605xwvnUPKx0jp+Sh40/EYOdaR2P43U2VxHxw8fyr9pQXtf/OE
ARmzVGVNWdJc+jpFqTbJfo4hDWQthddRNQd562p6tGt84c0jPV9Le674tayu4Loo
BD6N496DGMdTpkeed4PgUQ7p7OhsO7ZRMHexftxRpFEvnPyAs29aBROR6rWs46RV
8Ulvf3OAhPzD25qkPnH9JbNFEL8nUtrLZgzAIXsUAhbcCPLFbJjjOHOdj9g+864q
pEhZcSUesoixDkwbJTq6KvbVyLrEyR3lJ5jGchLKzcYEcjx9AtSveS/eN755Nsp2
dVcGjV41D1AU5HmYAYOhxJC6d1uq8khf+lJwYPeP1JBi5LeK8v3OVljtwWifC7ux
hG8ilIFowj/GRNjph+X7jKhV3227Q5d3X52a5tfOXA2XHhJUspfLYaO9DDdCiqv/
VJY65Ls56AnaO6kMUkPVzSDStZRNyYSHYr0x0kCu6Q03GpjWtdwJxb20Aai5gMU/
RDf+C0Xt2WPii10PHoyOZ2TRQujvuRQRO+N0enRdTAxPQ8KZQRxUJqRfOUmYFVI9
1OBQniYpygA2oBaumZc3I7l2t6bd7RbdkPPxTXBSeAPNpT95TTfJxhDDgqr7pg4Z
uNajuKiQT/IvH8YS3HWIhIqVBtWpu6fMw40zOIQ/vUQFx2GRSHXSCNMXUB9wAx91
9HAxpInsoKAXCw7oPzQtQXcIre+jvgWLxDdqYnVIAo8qtIN4GPl+BFJfhrcrr/ZV
nppzfIALFWXgOrGwOa5pCohxVocVNWNJiB8oTDQDI+3cfsLdY6orKRDKJZNLA5Br
PAXzy474kanO3KJQpNP1CsLKJ3gW6vL3MZRQS6KnJyE9bAB1jKbuzwANMAZRJmA1
vFvpWsPjD5BwoOPSNZEAuI4Ze5YX2hH/GF2eeCB4sTsuJE1YcOXwArh8//MOilW5
HLbIzpBIUI/XLisu6pfZKK5epvg0fsH5QmviEBMOeHJBxGbPRAQiLoIHg7MYo+gr
HH2oAO3gY/0flaz3NYKJlZHdQOa7M4+1EsQSAaN4Ixtxtr1pXbzY09dDhOtzKa2b
P7H62MCiAnG4lptV82fMFgBGze2KQtZ2937bIsk6Q2fq/5BMUfwCVssNSvXrFjmX
1bmguJRKFsrGIYf6gAlq2mtKUpt7oZBMjlZV7seRvoRRi7lshGCZOQO6TuDDDmUL
fJRzdkxKdgBRhYcHf2by8DD49g1xYEWLwhfKRh4eyerR1PzROuQ312rSD1j3976+
LtVdgudpLcIab9Ny1ogjcYtwqHwYT/KOj/XcaM2EH5mVBosNyRcM4F1UAGnfrqif
NGu8v7ZA0P4l7/Mjr6sxNuBtlNEK4HDcc4mSTkdxxEMiz1bnRqiSTQcD3m/ct6vX
40HdvEyzpKWyF8sWxhsOsajqffydM/z4cK2TGxkg5+deFAukyLQZXwqMfBjYZrEh
JqSowbJuJicNjBuwdFgHXAidw1ETv4ZgJZFJWyEjEb8Ta3ZLOtEWujcdmOuAGMXf
SBmmJwICx4o3MnMVC8IIJgTrmEEN4iOK29q6Fjj42QEbuV9WKjL34SJCxU0PrgFf
F911321OtCHpr5+5cH6oRyK+EnamvmIG/Oj1LElnI3nGOM409ifaalFRq8EQAorp
VkGkg2eIyoMkK2/ascaCUvRTC3dQGdiFEb84OJ2hwT61owmCA7kVpvaTS1nu/qn7
jzvpeCWgH10PXuWVmgrH8nvYpVYYgn2fGDh42bKR2QLpQr03nbLqUyINGpnsj+Ls
b+FGVwYmj3C0qP/o+lP2pG/6fSHM8rJm2bcwt6gCHKJpy2ey0zeWPb4Q0gdcANRv
Z9ThykshaVG7CtVPBr9ZuIL7aMLQL64HpVokaX6wvVNToBRReC6bjCSQoaJl7j/u
p2Mdk3MMbqH7SdVQYmMHquKa06P3xdx3eSI3EhSErv32bBjrgM9PJVNW2kn7fCnu
QgFfe4Zi4QzAxKJerfbuUY7F5H1YZbsqDbSnFgttxLujDHoO+WLnCKF9AmEzo4Uz
UxbOUc8g1EKDaAEYBKjUfV6VcKEwGzFdZ3sZ2WG09vDZttymBL5EvHc5/4EWD1Af
npyOapse8uSz7/u6CrVYQoLHj6yh5iUVBCsO72LfNyOqGtaWmHxb7BIYPj2zUuHa
TpxFdmNpMkXYR0FO4M8eRVHf1j11kLXY2wNNdJHrUAgOSbnM7p//eWNV5gGoTKyC
+wtHQD0YSfsn3GVZPPsUXKgJorhKwbEfH5JrCv6aApVuJ/eMeBMDCCSao8lNDfsy
pn3f1cF0hwrEvC4WUrtDLiezp0qikrDMiZ0J+x73VFXViruojQG2QvSA6QsPGyYG
onazy9i6aBNT884DW3toan7cCkgdEO5rwlca/NnI0pRDF+CIIzxmHE/Sf8e19kyN
4eBRsd61hInQsWRyPQ38fJtJX7qrwxKa6nN5iu0TJieJKeU7Hp3cbDZJfLx/0l6N
w4SU9YOrO1l4keroJJsBZVNlF8SluB3nJmXQt+Tzf+pAQxR8xZuvz+PuCyd8SVGj
XNzj5wnf62zLosmqGUw1bcCMz5BeQ/9BPtGgO58TbvDZL6dkiuYopM1nZhywx1OV
6mljegK3t+Iz+3+fA4qG4Y4/M8/tGilJTDSIrz6sie7I7CAgDD95LTfUqbu09sda
8OHhSiY6yOlAAl+2/pn6iOkVQ/qyrmjLUCBsg+32v4EOowT+MB5Wnzg0PfjHwOrB
4y1PqcR0/HQIVOt8eQJMrTDXICSqmLmsVDM9lOejtoLqQulPuMQniYogkrVWgAnZ
ZpNirr0nD5rneOj3qqgce64xXZcjkyeZsO4fBgEQkewapPAaN7wfYv3ZYiM6urn4
2yoj6/0mq0glx0Ww6KcsRrBVwY5Ih8o5Bg6stcqTCVxEn66uA8LHjN+6wRqKkQFa
VZErPyujZvrF/9wOVV1UEgMKglzzZUPYBDYfxulM0xISfkYcG3bk9h2bkkCOUFIO
dR1CAd8hTER67zY1WBIhNdNZrBvoHzn1DFWzpKG8o6iaNHDKzeEg772cJxHHbUya
r5fO4+K9KTIM8L/MtzIbV5SRdmHNVq2UWDF4Q48rIBKksgCNo7DOsgc5IfdUZA3D
Sdxq+RswjtXKG6XjoaI6Eir+FUbq9F/Ejti634Q0g3NBS2Jj3b615rNEiAnF5voQ
erxqzLB1RXwfm6eCqvm8jYAOfFvhN+jAgnGsOpsd0Tshg3h9MfySGzgmRfwvLdXP
z6aCiT3uyHyp/dntzPktUJBchrkzELoeIH2ag2kb4AtHuMNImMMHKpkTFbw8Hy+h
4aPmJfZtBofnqU7OD5/uSJPi3HGiti78WjKZ7FyJIQe+jaxBPmbMPb1Xd3Vz0wnl
bO7bBjjymEQ64z0JZciq0o3AU7YDBTO0ixdaelbyAMqHwV+jgEXcn/9nqcWju7yw
X1nLsB5fDEqcFzOg56Up73dKeGq6KkO4BiCZyUGGyGBKD+A8bIvS4NTVJgQBo9Xu
KkR5+bjmsmAbsUjgIVUUAoKC10jO+WM+fHz6S+kzqd9Z3G5HQiy1e04EnTfoD+V6
Op9itiCwwcrACzANL0QyCvw+D/8Pek8AXONbOOMiUnPCPRkO5mF6e4aEv6ns9Vkr
8yPA50aewfFEWbiEESX4W456gNt+GR9C7MPXkOFGtPxJX4uJ0h84L5HkVgmqBNoS
wmLpBYmrw1B2Cj9ang4D/d+TsQb7TT6XeD++Y6z6j2uynE8gYZiEbcYHE2fJi4s6
oJNyvLZVBB1Ca1vsJ7gI42Bf4QqKlhB0R3dOR9yrJM//0fQVS4efkjWyEP351gN8
rhugT3P7XYPP62jhG8EC4B+LQ8Hy/cxKUpr4P9svYZ7vpA5vbeU/8nsJiLG8xInQ
Xg/O5W+8mfffO53AJN1c5c7LK5J+p7f7cQygXkWJx9D27qEOtE8eGWUmbJV4ma6C
FmQhegbBmEm7ghrgglx9DdTar3whs5ZcWTjUp8yukwzWErFeRsH1i+aILuP7Z4pb
gftkqauXb6pOfae1nD4Hs2IP5IvGOcjbj71B0CSqVVe1hA20j9kA9vQ2zK5qKMc2
xtNVOYPR0CeHzGDHOQbrI4xU26wmOeAP71aBvEwZU8ZnKI80XZ3vdzX1s9QzDyvt
wsPXV5jBPZ22IVRA2KirONg4XFohCdevR1b4tc3k+GWh8GbSVhZfSiHTKSEsMVnF
kkVB/WYnolMY1CVGbS36DtR8avKccVTO9wBkVsSiTuO1f/7ctkNLPI+HZKMRRS4N
8kPwAHqpKmMgyqA1NZRmuVaHS+uORZ6hXVJsa6A2USyUnzBms2mpmDi+tWpiEvCW
SH5JlU1NX1v+VywXPykrVV3L1Jlz2zU3JimO/3FPQLJWzO7+21nYCiZ9aJAe6lwo
IcCaeGcp/Us2+LsbMUy3arTRLiekRkhdsSkjbxlx0oJgjqQJDewdlz61XdbhvdzD
8TvBix1XsU/hik5MidiraxtVosZA4EVapZ96AbDR6WcDiA52jJ5bgwJXhVqTC7fw
Fz9rQtgcJ+QdfH+ZHmUWBfu0hn9+74ddTtwU8Ro8Dr3RO22YpBXw9Dxfi40o4G/k
nRM3SwjvUtL/Viv2rbCQrXKd7SHEOLDy4uVsPJunNz7Kcc/EycVWh9oBK/A3Q8xQ
LE/sWRp8AkqeOwcJpHvkvvHSSx2T+7Q/vKcRrvRi+4lrofOc0geujwbraq3AVESF
ySAhVKjh0K2rXxPGHMu3O3CO0+dHSAPnY9ClMyuMjLAMV/IGbz5kaEon4FMBMxXg
MtIxhaNcArwjLze74HX3+5UpECWy0S618QVjPegDs2Ry/mv1g5rnvNU4rCwr7RKr
fZSGECGqU+OspTmoXUcOTuagTSBO0eDEFzng3UvWjEVOzLgrQXpMyrqq/FNbdc13
ORd/JRR+koqBa8Dcce0GaCiESv+ELxstMyMwfmfXFx6fYrGbwiGCcV/TYCjzYPSO
V/8T8wRTLzLfesvFrNdhVUT69ae/axlT2aZmDlvn+u9Yvke57hhBwngYokYkda4w
3QpJCYMIr5WzoRqH29+6RvG47i1dMURwATYSBnjpc7JpQfg47xYEK8ErbQ6FBhjG
KnKbIR3vM8xpYhimqvYB6lYjHASwpPiedrG4FQLGhwlKCzXDTo30a0Tzca/F9WB+
q+p/3RzlrOmz3gQrVo3iWQ21/9FNNl8CDWj1Hc4xicyZvRN8ntPNBXLu3d1eNvLt
hzUsd6tuhu+uoif/R85dSyOJDD+DT/ZNfYXGbnnATiS2SvIh13+5DvPD7MFphQni
R07lAoNNzcwVrRKYU0/9RlRaMVTlx2mPbXjs0kpOR8mYm7OEiafcz8s91trtSYT4
d6ywjynR91hedplW/EWV6rMu7WFP3Xd1gy32hnENEQ1dmUSCrqCXYBGJkGIjgTUF
0+iAwusau2GheqHs/+bzb5sydbYZIxq2vPwGNEGeVLmqoWzo0C72IM05ud9CL6cQ
9d8iHetU5ey1x9s8GAFj521s555A6zO9JAPw2dhqyYsSAkxmNYtPr0s4VdbrXD80
iyHNvBBSRk0YWUFiDC9pmMjIO2kq1SPH4alUTAg8lP3JX63jx7c09Yb48YmF4zZF
5hum1KgSGFQuGv/3MtRQ6hiInVWNifmJQ7B0c1s2dSm3YMFAgJIT2v1Gq7vFB1ff
3lWNbtE2c22QbZj5FADnRAh4ZD0oZMM7z1rcbVgzLywhpJFMQ4d2zzlHnvWotiA9
xssjetXJGFHiwOd696Tp4ieNmLI0sU2Hy9V57nhiDKRef01lYhkrMxjgQvCnjxvF
v54Sn1wu7qwit56xovCmem8cwQOvBB6XxM6731ozEzZLUmLQBgkFwqz2m9l9ST7M
vgZtrOeIHLuMgA51abgr09XkBkei8ByJs24Z2CRMdV/7V5s69R0WI8gpEqJD9CZW
blvdhkBPBVdPDg7/tjoy4dE4IkHwTNnJoayR5Eb15TVFsI1IrNJxFqLadCTp9KJ8
gZD7rD/b7rfFbaWSDPThTIV1rCWrMFb51tHfUEbdxggnQqpRB8MR+kuT49HSwaEU
FC2IiweWxnS0kAPUzgffTONHs+CVAow8arN/FIwLNerqadWB1jvptB+6KLg7kXyo
QbqZXxxN/EJsgpRKB2VsjEa/4x4/lGD2cM60KTnx+cWTlB8GJgSQjQWYGZJKGpIT
HszupJR5kFxkEzdFoidaN8Tn1fUHIhTLbMEOZgs7dQc+Du4bzB4pRwEgAMVBWYN6
7+i1NdVpxG/e2Lx46sgpfoXw7n3ARbr9VRvzZMbINvBSVP9akkd9HW9hrJ9CBZDq
lkMF7eXevAhecJObQ6+37nVaYZ1AD3s9K/qIeMVif23Q5HN8LwzB47UwR3gsH6Dm
D2ocHLS2195wlb1oK87yREgS6DDvINcq4Wfdti5x032yBLe/IRaGTPlIUnMSgdBc
U6WoaWQk/fZQB3EJytY55lm4P+vdRwoDikjQFt5qxK5BnEpqOAsuQLy9sUB7Goxd
u80+ulKUy51fOr0aGE8Hhk+et6oI/ZalKhkUFK2H+OB6f68fO/J+DKEQK9QGykeM
P4ByEGm04dSAxB3SPrj8foaxqbFd5nFY7A82ADCV2ZfgFYf5psQHUtpjFf73B68S
BFd3BFCWeY7aQJBgolPLoMJz+ytEhOMjijX91Nq41BHmC9qPIHnNZre2LPwKqsdR
cn4LpSDKbOqIuhH3PlEYedhmEDGub1GRgQw62HATt7Zfx3it/gMhBiPCzXloG7/v
ofH8Qo5kRHxQvE64qaCO/oNv6FXO3Tm1fzep6EUK4F6lu3eY42pZ46G7gb5E/laU
ESG+U0YikngIjIlDxEVtdQosY2qAxR0zFkZyi2Y9S+bgvEFzkiUzF83yAksCbxpG
Ud4b7ebsGQUeh341ltU3Uomtjud5VUXTdBIErkC7ZrIlSyw4/oINmNgSaP1nZiJH
jGK+aEm0fa6sUxZ8GAmgplnVKl8QRo6zwej+kdWT1wKcd2IKcWVIlYvXg4OxFwmU
G4Zw7iKN3keoM1qK2KTnc+GtRj3DHU0PQKz9kOAY4QWN0iqxsUYQ9vw7y038r1kE
VqSKnvifIsVmDLz6/QDMwIucR7lvZgwBiH7ZDx2eCMSRS8hGT1DQE6C1LWBnBxS1
Ts54/w6UAM17+WzfyCC/02rQmf3+Swd7e3IUxvB++El4knIy7o9s32Lq+3A5PPXG
NvJZ4Z8+CDQcOn7zKTtyysrCk4NOeUb4rI89EHj2qpzSYpz2qzIzT4aLw8d0VyOP
RnJdBkNfOQN+0tSaYHwpmsetEIAWgQLWSkcXN+dH/yKPejhLGyMLj9mYXmqOAyJa
3Ca2pz8gNYbBvyrGEc4yA+yrr83y0cBv2w8tV0uukFWM6ry7uvTsF6vAAuLeuzyi
0fOq64gXf/GEPhf3GHz6mdSmXPaB28pTBS4tJMXMWmVHPGcYFhbWOo9vAOouxraN
zZr7EZHuupTKsCvs9qx8UDag711QVXj/E2feywk/P3kcvQdg5ZjBVbRunqBxvcvP
lFXi9DQ9gdYSq9v1yNSJTadEl3qKZFCeMByhgEqJSRD4e+M5qmS+qLIiEcPukU5F
7mHuJoLYJc1GNi6rzMSfwQ400v4wOFLDXsQOBH7TMB1YRuDSVxKey/FZewHpx9VE
oSfVejuoNZtokYrz5ntezcVhrvYxQ+HSQ7TrkSm60/zm1ceRTtBSnzpaI13HBXso
xa1jHmY8sjf2ghelid3rr6onBmxtLJumaJWc0BPJdMOBNYqzbakbfPswP2ZWafvM
FkwPMMa5q3eWHqHt4XuvDE6aAwttnQ34JuVeIUWyAKGztcTOBeZjx4YwnV2gOx9Y
nFinE2+BweUk84tSZrIBH9h+lHd91EZmwmg5us97S2G/wjEVz55VRa8hzKB7sjDy
U+TTFGCcsyGZwp4etwDkAGGEEoaIvumsPiVqJiqaI6+tVmFtdXtIy7SbbsUe4TjL
3Gt9wx+eHzyz4gtAwsypW4Cq2ibjSTib8DMGYwtX0qeIC1wOBQGeAJ70sTom4FuX
WNhB+GCvvRfaNJsFdZ4z9AJMMdMC5tr+pvikoDXqONk/PLxcxJHaDDGeblBckqoR
pwqwdVWXL7muqfSF5wiVwxYSfoGSm3JcukTqBYhHlBpRAazJusuS4cZz6XYqtfCM
PTZSDFicT268weqc2EljfMW4Js5QWv9TvU72GNLTnDbXsqMy/5FmAr2V7knXayhY
f2xBYUA+WNeWFjL7a8asmBIBx/worcVYmdt3yUG9uIg2vrbkpUiCZVHVPeW1A8gr
bZSD8476I2WwgCtUqUNOUEQ0CN3px2tWB5MkZbdvuAc9mudO2t7jHYxayGTCKlbW
QSAv6NIo77FwtDeWL445EHHVYrK2jm6kncUki29ngQyam4sO7ibLCr08TIkeJKYY
skSpx7mBMXtd5ti2OBzl8avxJlAJds/RTYTjNsmywN7SXgpqosy5q3AmQ1yqywqx
nLKnlaND8Kzm38za5dsgDRpqyH7gaiFm4dinRJ9wF0Wc6ZA2rDWQcq6XZBq4ONxY
83hDQGgBa07YT3PMMJ/q105lzI8EfOvWNlNhutiFiF/OIRW8dYH9FUj7A3Pv2GcJ
khHnOJ25IdEWZkSrDYDKVWYwa5tpy72lHg51aBLyDqpKcWb+insSUcrs0nTsufV/
QTTq00mbwI0FuQ8QNVjGareZPVpMWm3pCfZgazbM6to6/z3O67GFeX0c+kE1wicS
UAHppeDwGemJG/zqMBkDA/cT+239P12xc2rIBJ4HMjSAf6MqqNNTxwUzjBW/QJwQ
5aZ3YU0PKyLUqIKigRlAbU8VcXrwjMpRk6cCYbd4sLJa4GH+71Mf30wLpkM/CGYk
7GgDz4EG4hulMg8DvQywCggxvnTseUh96i2/gtGaZUPqSSM0Q+n5H1roKNO65b9o
Mikuf4x04Dc5xdsMYyMqGY/DmmaUgXFnYUdLmZ25Sbm2XYbw1kIUl25RVLW5oWXa
5grtWZRc9VtY3IwJTliiQqaAbbiG7cNDAbDjvZ4sXY26Xyt1A3CD/WcCzMivbRQM
zi9CVSfwB9DQ0dcmYvZL8g57I0f63CEdunJxODJkpaErJH4w/oKpOSnXLh8l16DA
RsDr4eRwp+qWu5kEM0eGa9GSfSvhYv7mwZsl/YDiTc+ERSLQq5IuzSQaS6TJO+Ds
MAkk6JRjNHQ40IdV6DGcIt89ahStgllCc9dvwDrwRk+4x+FLpFksB6w5KZ8Og6Tw
lSlUzS6UTP7I8E76w3pdAjujHuA4/IBOUJi4a2xJxqrnwXzeCv1WLevBciJJ8Rkf
g8rkhtn6xxIHuMKwXQhzgoPqPntaRgBr3LiO/xvAKm9ZpcpODAd92QJBOKFEbOlm
MEPnG95P8saeKoY0+ktdkZWMJhN6AmD8QkkM2/SiqV87Lm+GcpZcU882I5xPNBpv
QkdiY+k8pnuYGqOj82M5v3mFmpmfPdEz6noBgqfAfpyS6Zd2iqaqXltep2cqZ9lX
NMTfZ/O3HMTvIgroye6+bCdV9ePYT48xe/41wJhkWrLW2kyutBsOEEUIgeXTnlSL
2OEdWlyyg2mPgRiZ22lgAx06mRpAhxXZr5cdCh9AIn/zlk3AKXCVuSBDk5bBkP/L
gUCpUHnYfhvCkVCXn5xdLVItX/R8f/zT6rEX/cBadntSeo2mcjWrTMC46Hd2rT0K
CLPaYFqx4I4yvcFu39nzqnAATNQU6ecbverzxaBrvKC0WkaXxsOQJZzyn9td/hXI
Zw5udI1XB6UghA/wPRdT2V1uS0rMkUiJ8nW0o12A5wI323eSsvqRzknlAao5dezC
bONiV6GVPySLrFb2+WqbrQgOWynes/ONlmyfZNO+/WAUjdSpu6tkk9koZU2zuNCj
9KyNRbQfUgq1h3vYTFFsRxKnq/sTpFJGGRE9o1JM8sQZP0iWZcFfluQVghcZwuCG
ts0AJvlSSZDZT0RTjp+n05yCSAZ7nKehD45pnJiATh0zVOSgDzLf7KMXuyPK1nV2
UKQEpt+G0js6bMig9MIgKv1L5n/+TJUPWu+ltX7fsyqL4LaVdPLk53CsSmEHMjjA
9UKDMe/qDD52uN19fvFVYhAtlaQHajHDgpbOzfBTx01BIVFPy9T1i1QO1GV8/XYE
VgUJx4DpacB3N0JqP2w/gusPJ8e5GGn4Vjb1pJ/g5Co+yBvm6HW4oL7roFtDtaxq
0mQ7LfIdW5RzvxCNT5hlKgIyzNQwAWXesGFwENSWG/MOgFchIbhuE1R7il7ViZ8u
MIxrP3WMRhpc2fCmgNA3YUJuA8mkjyEALsAuL92/oSKo7YAi4Hr0gWkEQJrCi7v1
iEqjo1CxMvpvC8kCb0g3bBbXspjO5SB0hoPogV/Scv9Xo9YPutAY3+Gc+P/drmi2
MO6iHB9oqbdZPxHLLOBomFvgPwAt85ei0nOv351T8ZyJVLo2zcK5SA5cdA0bscZJ
FO5uPUuWgv4dCgFR/ucP7J3os+ts3Mq2Bp+0Kt1AKNAvERKRuY9pBroCAtxjy3c8
Qh4rS6wgOyPfSKK6H+QO1mbaZty66rud0FZ/o9YLd+KyjFEiBvwJ3K+VLEenu9TX
aOYs2aNXpqAsxZJ8s7JfjPZYTVegMFyAixXEdt61a0pgmF9cf2a1EcaTFsSKWGRj
TzfQNdRoXFMFTs1v6B/BOZmaSdPqiW2zcpLcvPbGt9+q1Qta54hDUzG26poW/9V/
3dVYtMEKAqEh4kEgnk3QcgPuvRQogJ169U6L6Ydk1FSOb8KUEczOkJ+NPGIBN4qr
AA3RUzGB3GHh26pDh9U5AU9je5IojH/6fjDgKpdA6kTlQ4pUX5PlU6P8mwiQOi8J
vuiPNWonR5ci00E23XEWDJ9xI1wK+Obn6/dCd9c3c+CopRF3ei522lpCG2atv8d7
7Yifi9W0p405jdKjoIMUvxPBy9k6VIPggEXHLNrLGcX42bZUYswkKu0U5VvQ5Q2M
Rr2jqbxuJiAuCNn3Vmd9VkuMtQFTKYKOqg3oCHziBOr/DrSIwrsNfU2mgvZnmr9h
IhWjrI0mxjuBdGXY23p3N/WWEiQ5RWbL67Lh8Us/rs1qpET8eJv7zJf66bbhhBuR
CF3HwEwwD2vgYpKJyVlEjNUirRg+Rv+HCSET0qkyZI44DcH0b1QBI74wGaoc9qRD
83Pna3RsViIcU/xIwx7sj5cni4crc7qXHX0v0tNll76ABuOhOibEivR3Gc3EpPU/
Tm1rkJhLGRen3FLtqMi0qN1lSRD2s9el8o0vTF8SPfMBQqnqNDRmhONOflja854b
j/IRh3QNjbmRJoETa3LtzW9WMIOmKvvp9OjrX8URN4P+akLOcFDk49hFh+OlBubI
0C0BxP2HRj8xIvKl1BCGUqnaTxv4ERbelbXHJyIQf0sRLlIyaZ5BkEi+jdGTBiSE
CqwNB+6YAI1myCFbUcrydcviHjbIl6urFi0TyRoUDbcty49bTnX+F732PjbqVXc8
Mrf0YBxZI2DJ83bz6jzEAtaCclNErjxE/J3JZbrIotpP/c3iCdn463hhodqAhCgZ
ehmy1W3stn+U4xC0ovZLmMmgujaWO9vZVUZY4Lgw3V2ScM/zRZyPjjEm84Ugb6NF
i7Zrnuj2nvJLDY+H2zGh92IbrPhZEtfjbR/qepzkab9gKIvwYcScA0/RuebNjgb/
tFcVmUqhZ11Swg4RgQc6bT6KYCemBzDvdfCoIrIU1eOP6aLMfbzEaLIfRhYXEcT4
WP+M0EYXk32fItAb7C7r+g6gOjTXpy/WEftNojWJTXmSPeZQ4zeaN71ujqN/XKvk
t7IdG1wKkyg/jdbjL1DPznDHcvJyMBdIAX66g7XtI4A0vnLHOnhpuQm+jUYzOx51
dZf70xEfVoddM5f4aRiDibD95LCYuRql5YhmctXndibaWM0UdLQ6nZRQfelwJgAv
FD/BvyvGQkK8TWlgk/7BjfRGYwijRmNMSU13BYCSX4J4iVnaxoHV2Z9LnPv/Bru3
bhjvjHRAkEuFlmzzTrCEbbHOXlARkw6HtE0bCX0vJTzm2gH+wpobyXaYl8KKAc8g
ISXJdzoH+THeJgNBvl8J5jNc/CoQhX+FeiKtBhcPVSVDhd+X+32hP3NVbyd4/lQE
+fObHOEudBCtUpvdWdzRcebn5LAk43vYf4w3rkZXcQhCFBi8S3Gd5m0h4oOBUqPH
FAk5UGG9NcWsbcHWYYX0aMYUHXgMty2whEMNGDfuS+lRmaZ+slH93GiFIBg6rjSt
lCeRV7GUaIFA6OZ9Z74FHY/fZMDHszdZbjyX1gdKAT488dZDYd5FgD3J1OCsgw76
+/RXQFdRHf7hE6CCgQzPhiegD2C4WYOLcgmHol4JNSnqICSajcb06lOvS5zF6iKL
CmY6nepTYxqV3qFiQ2/arqxp5i2sqzgwvBaziOfJ8yDmWuA7jWptFRnhqYxfsPh+
4JVdgTrREahWcUaHKsKYZ8OTNOcnNTO3CbgnxQojtJKfQltwXk5oJwWO83emld7j
sPDTTxdKWUT2j+/iiZygUNUCRXiex22L4NJC4djy0b74TDoiyyxYVpVnTg9v13t6
Z8DUO4EhWSFnBXcRogD4/AZuJwloeKsYaxuQzMgWSdeQ+NTDiDkGMAoJqNFVCIUm
2LsxuuHS8JZp/QK2J7BlLZFXy2QCvI+0bOyAJJaDHj/8smbpn6R5UrBgza97N8Gk
s4jttrVi3YUJ0t3i1tLbEv1h3+kmK9TlHM1YuAzd14y25UXj5gLqCckWQVEQqU7i
wURwYkR5wXaT3tXR4iJw4K18NykA2vpo6PSoDngUThpaN/VIVZRjH/hWsgzRhBup
sHnaWK6juC1/FP3Hm88cHEy696plrUwe935qlsEAl9jjCPm4QMOFPIeTpJHfJZiM
nb6Z3i/WLL28OAUvVjIVzgMMMtdlfxatZ/HPkRKCcwGhn2nbqNKVzsd+wxmfzcU6
4WfhjnTZZgMhh0M2fAPepC1uvDv7aomz+sakJWV3ASi+E+BWwsdx5LI/+rL3ju0U
fgWS6cxnHtBCVqcSFbGetE7llTaLkr6faXEQrwEI+9Foevr8Rzymu3Gcz9RhGTO2
s8UtE2e0PGQGCF69CR3thSZKBuXWIim1/ePGAyj1uJnhgAGQ4dIDr953wmBzVoQf
y5ZofblDx2VqmvynfX7aoQbzhAC6+gzJaMr8xT7nikOr2budFy5eTtgbdpIXZuyg
PMVaSBc3Myalf2w8Kpet8dQm9WRvPeANpgRlqJS+FbiYYJmL+fILjzi9mDSug/XG
f2iVJs6E1iDNbQ2Q4GPSFtTTbTk9+9mqVe+fvuZBrcub7RPqG6YuTiFnIxcdwA0k
edVCmi7Mt1638OoKIBRPBcq68H9P2+UUtxBo4beTxD/qHEEQnfiwB3qZGZR+Vost
VYaty3w4tFzveNIIy1lljbCehPDe15LY2c6MrmQdrQMFJ5PHmqxLuOv5S9OBY9Qf
59OMhWa3sFietLp0sVZFExrn9e8Lc6EBsp6gaYRwsxIRiCd2mS+oOciTIPdPNY3o
4GyhEIG2mFfPIEG6S90NfjIYHlaJ/78f8jz+HONTA871xsmjenTz5wRhtHgMNylt
kmmK580wqivOBL1wbOi+FSFCyONEkG7wgZYSH+AaY4+8lK7lncH7+VWWhB9AF3qN
p1tZF6PKyylpJLwNlaPv1vFBys7TRPZdMPFfOEYNrE0q7NMIYKKkHjrZUa9UG4q8
R891CyY0Frhaab2L5rzJYUbqMMijQjlSRWGay4VLm5a+sy890wFHa5yKeNPCD/zJ
RdiXQWrIWxzZTdcEM9Iz2CpYcIB3JRCb62jzEThwJAzmraAlDAPHXyhtb7ljOmwm
vIZvvKU5GJAE89y0qk7NMFpJb8qu1qJDCLpnCBXvOmF9hYRiVCMImvBFzk268vXz
dRCgyRaa+HGSl0nwvyBdE1ByCdQ/O8vDoutR7Cn0gtssV5p1ygaHr0qHjapQ94jm
gJicwao/YpJdkyceKYJD2FuTOnVA/VjCD2D7XI7I8H0f7DWJPBu+7k2gpHlXzFj5
3ri7k/4hrsEPPWCP94y74oOA9wkSAUsXWjl7CJu1zWwrAlhoYmv92WOZgo58pZIL
jsbXHwxkw9CY1RRT1poibGZbg6Tugt0oNs+vHoOHE8OiYyBER24bbiWf9QGN12WI
rJhVEUi0X6IoU1AoFDSK+nsffDqToBpxi48jnBg3Ne9DwadKK+hqLN8UPy7jtTWa
K4qzLraSqqlKjfWe2GrriCRQ+jOQ/RyQYm8hiwDFPT2e9VKHy7/wiUJRfMOEXEOX
w8h9JqSDv+YvCS81lBQyO/whZmjqy86wZX5wGMfmOKRSVYSLs+XQCn/U3JL4LJS4
DfYEBgKzhzBuCjSQYACxAM6MFe2xz2qaM6riq1x+tf2h7PVhIrSfWF2DQ4uqlGcs
T9SvVKf0GhorUVcfC/SK7uQv3Bhwx7j1/CEQeEfYdNfXfH3NQm+Y4w46lCAvhzkU
p80mL3DGKNEbmxO9AqvKVdtpimnomoMocvAJjImlJkbmjCT0dfi14bQSp4uan4uq
bw0ynu9FHCKpwFGBXn/wROfOvuQ7pLFnjLgQ+GO2iGhmD4qHMurwxxXJBr3ygjGU
QpDKDetfHvYXhSYvxoJ/f47TjZc17KaDvEJLoaMq3dIx1H92yxNgRQy0Y8KxFsyO
AvucEJBDrwi1ugYH71uLNpVZ6J1jdzssOPpqlNA/e83suWvKQMCq9qcnclHzRe1T
/Np9kOEzOP/NnHX2Bzv9UGT99EIQIY4Gdx10dA5YX1tD53azoB5dGaeZvwbv6BNj
amkkyqYpCcR6EaRYZ3zev5tpd4wpV8CAQw9EBw3rujrdcJcixlD4HBgS49N6Jxqb
HaMLfwAQIpj23lOXr73UvRaWDqe7pj7+7NGnedHYhhOh9eFjmBX/v35JpS2c5syx
4NSaZMsVF7HrKZjPXK2BPNQxBfszVM6tM8cm7dUqnf6nYoCx8nFIb+aShkMVR0Yq
pkQ9Im9g4cr9GpfKtDZgUKiz0E+PmUk07flPrpxyp0R4HZ1CsWb94o6fIgHMQinD
89Qo+brH+ESQ734KGYkXC70Br9gPIgTslID4u+VzUbsEDRCCyOa+QJ/MScbTg4VI
Mb5CPdsvW/y774YuEODDVKQSUkeHFEbyqD0fFtyQpDIWzlgcj1Ks5MUdfCWfpO9Q
OvAzv9PJj82FoXsYOWbogxPugYNne6BHDBHW0pnUGHRC5r2sM0t8wWjVdaVa+nup
7TeNBVoYRFJIeKTyZDo6v0Dw0MInspFhRt6z6zm0iJ0I6tZtDd+Qn5VzmmQxGrhJ
GUZf5S2XCPQiQIHOkq8aGe6gCULiQuQMXr2/2ax2Qet5H9y5r+3+CdIHGnCdofaS
jfhyf9eGTx8SGosklHOfqS+Sa4jssCHHQcUFg+mylFDFsp4/fjVmLe9a4UeHIMKT
zdXCF7YcqQ64OODY34IyomqZTtj41PZSBzkVLlLBqy/nElj1+DcMah2hdQjYv0UE
aVY6TpTDOqLYfOCzmAV0PNNYR264+lS72gFNRCVyxXU3tmfdRFbesrd1ekQdGMv8
PkUBB2GYBN7JV50DrLppIqPVkQFfc3Mg6TQC4OGYfSaaFxTyFlMoZbkD1LoF3d4s
uqE0Lgc2l9D0/j2fJhQUf3Ea+tu88EohMAvUYqo47QEbTlcIqt0yG6JIf7uqjIzD
ick/gQOJxArEmcUjfFa8lULD7xFc+F7frbc3ThpazQIiQ0qlZsLIF3yr3ci1cEHF
KWgwZOSz8cDJem+5DXLznZhQm3ORMRwOEiAh9h6dg+3wYNxP17dBs46My5zVn1Em
CDSTvqnZJzHZTIvBPGYG04rnvJwkVIPd8sv5uwA5oMG6bjnRY1QE/X/3MPeHIww8
JfkepIxpOGQY+5s8phA36d4Nr61G84r4+uZVovOInz/rvRb/cVW7Eb/L51aMeDFa
RhtffPmK0jX3jj0M31OpF7uUV8HtnymO2ddOA8+7iZ/PUjb2MmTvpUSz3JRdPB8+
MyOqkvIeJmljP9uNap9VrN+SV40+8SLSu7XRUR8M3ghBEk2AG9tUg1VLU7MNXOHA
PiBQAvAzALSg6i86oqSTg5uoKbBPoZBzB+AyZkXKIeGkbJVBVWWL94ee6NioWJzc
oulOEV2BjsvKN+X+KjPfNJAzxDUxLnW6BKAxl2RNBfFYpssKKWdZwoi5aFNvguFH
AgKX2HyBPmjmAsLeJkkd0bCULs303SCF8aR9eKdSOaRFmy/iDoqXVE8wCTec9LRQ
a2A4ifdlhrs24tqRf2cdfUDbwQJXluX4GxGex1BPUakYWF2S9a6LPleVPkDAXJe1
rCNiXEMOoOveIVnWocYMT9JyyzJgYCqx99CzE/u2Hi2rMR3VuWwtEJEEOZellNzE
n0Y9dkLVcb0UVuUSW7iURR9jp6fX/TItUm9wqiae1dUrMSrneM8g8GTGg5ZGGchz
+HP0hevbNWSmtgnFVQVR75Y9Jv/kKFsntrVznwr65T2tiv0XY1/E9C0WgfOmqExX
Wc2TWu1DVObNjLhUWZVZ9Kf02kVFV8WtE6GdPibD9wdevDmxJXuftNQdiZJC9pkq
uQEKET40pBK5veVXwA9hnWcoX6CKRR7nqNXOSgguStTLrB4Cr0QtfQZyx4/UZKot
4jxpW/3JfgOYXdD5P8AtINc1dOn8TszhAu/DeoBFDvOiuFLewmQReg7Nkq92nG0n
oJzOKZH7gZ4Q92XqFQcxUQmgPFAo3Q8CIOhHZ4zPw5SKG6+kKI5hq0UI8+K1uBgn
867GzzCcZ6Qa2iwUg+HQuX9ngWt8Abiyt5mYN+EXs9CTP8MZjXN5VjFo5IR4A59L
Lt3n8AXqR5/GAHBBVQpBtOT48FqNG575eAoQoiYfqipfNt3LIbxWgWuXlEMwX9xw
upKWlR2MbDiRkBdYvLtSqVPD6aiMkY7fdVDrGRcZ0aKGyJrT0swmLMW7wTcpZiOj
XIOFatzNsmwyYgjygLi6yiaZff7ZKst6jRLeD9nKu+tZG9Yjo1d/8ZuUAiiOQe9M
BuM3JiY4iDQOak4HhmsVvBCVtyDYp5t0L2x4xUVtKIO4HwjEjqL9NV5CGXIbpSQJ
Smqryi+SuE1MyzWYrB+w6kslkIDueqg49oIpEJm8/O1aNHQvbc2PQLSTZwX3By+U
R9vRA4ZTEo4/8fuALdi8hEbkCmRi60H9DkZE9np1En3r8V+BZv1KAYReEaMdqcNP
ktC4lltKfjHGu396lzboVK3p7ehrAw+Lyp5I8K/rHAAR5gBH6+PNHtHhRPWoveix
lm3PieMvYurHLJ29y6j9y9MCMSWbw5oMmOsxiZZIreQpkiVJF6+sLT9svislfXTj
AD4azWXX9CL8k09RvbEhwzm4dMVcT38cliLCxEx9UgJxhepY7K69EoPEdIBRBVGw
+hR6IShXoHYP6wPvJGeah65vXU7kckxKwBg2DbsOZj3W2aCUs51kiZvwH6G4iDPf
C9wtHDvrFZHimXf39Ce2qxwuN9m2LEXiicD9xJ3DacrOs51u877WAckMcC0j5M4K
YasfiB2zzZDG42N1X1Ub9mxDX0oz0A7jc+1DCSrGJgiYdtNFlaynFI9+oUSgaDmj
4QuDjjxd0cFdJXk4VKZYVdOfBzID92DHAD2rrtTopu7qL0qKOpD/kqwDwXCVkjPv
R2mFdNPtEDgqcV7U2jJ87zvfZJpzACc6jn0EhYw0zI80Ob8fVlVcgRiTPuTbCRac
UtAe89XROh5cgfu9O2FLYP5tL4e64XawKGedEyt9+1XkB2OXQAd/vHZAirfhkdKq
2R22TylRXIp3M6A6wSsHokGICnX1CzpQ5qQfgTGc4/RVMZPbpuYodqPV/ITEGZkh
JHHLf/CVpVVb8ucKOAcyWoXM2+y0EFO25FMmgIl/YWoOVvgps/G5MKXLlF4+2Tv7
XIzyR/Mbypj5FozhPf1x+7WrmaXAyhSzyljTTjCGvPB0A/MlNpB6gXK+XqCh/C+n
0gg+gLRWbV+lsYTN0MfY4zGRmpWIQBzhFZeCztllyUZ0tMBnB9yK/DRmJWfChoBP
cq0GjRzO5QJtmDgTvjEYCqBCzCZ9LXoqmWAVWHRXOaE=
`pragma protect end_protected
