// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:31:34 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FoGwMnli2DPpQ2P0uLdNdK6ubtH2CRxvHafcdFwzBJ2SI404uywcuFNN46MWFeeD
8qyeQ2XSl7dpryQUihno6B2gLS2ckrTbkurD7UTLj7RJpuc9TmBnCVMHGSp0sOtV
VwcFXjmYR6RTS5qxmEFpBCpOciDcX/XJEYLH52jFpNg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9040)
AmPrR2MF5+93StDck3nZIT4V/49mK+z2paM8XyOACYxjOZIOx1N1nwamXUxRCr6a
XO1F0rR3WdZQnyN8j/peLryRDm2IhOAiA+n8FowSIQnm8+RGzM4s299kB3B7292m
OAdlRAPO0G9TB7tXwjVCNNOZz8h6uU8Luypdv6n5Ez14hhYPx2Q5WaSteoyyzONl
EFBXTseQYDAoVvrzXUIr4gi+eD3lRj7SyFHheZ9V+k1suzChx48XVXXw+IhuolRl
nkbTWP2I4i2sykTlbinw3eZSfm1PNpp2VIaICii6SfboxI1GZr49GnIvSgHpBqWa
ca/A6QCrxaQsi0VdhxdH8Obx8fomZjo1/DD4JxIOpK7wy/ICpwOF6FycJzz3tgL/
mMoYE3bwCu0MQBJmmYoF0IBKwCwcV1tdwTwbNhdO1drAMP3ZfJcpq9vsR4iaajas
sBAN2kXT3zGCAPwolYP9vZH7KB7ay/sAVn3QQIRmv8Ax+N3SHuN+hL56c7H8QE6v
/u8jIs880nADGLVO2LfzgDtm0ypcEZMFGIwz+h9jZiiOT4VgzfaG3C3r9hwkyHkS
LbQKB6VaS6NVzuTv3spN2IcSudkRfEBOSSkRIheHDIEgMGnH+qlCqvv4yYE9zuRo
6JN3hZQpM+zg/DBpHIRVCzMCjRVKQPLYD4MOQr5XtIxeUpMdPnj+jnAsHFBA96jK
oa0+0VBpMIaG6fIHAwjxNf3qy1QxM4c0DfgTMydPg37L0OZiDI6/0KJPTEgQnt2o
SjEY7jkgLEK9gEn2egMDwvwC+A0XCdCkIxmaTOhDdUf/imwsEA25FqN+9iOFeH9E
5irqBgzcdVcv4bXLkvrba5NZV7FtED0uYcVUq8U02tOyEr6c17Wb/1pDNgZffiW/
VXexPuwOU8rK6nPD+AI3lrWBzaXzSyt5UbQ0lLL5pldtlz3lKR2pPee4fSH6Fmz6
S4p2G6aydXWh2uebhgDxQxrXemK9o1clQyqSn2zJ7Sh9YUdRg6oJNwDd9WUy7tRM
SU5qMs9buqphOyEWw/rJisgV68FSDPcmH/UaYcw0LmthJ/siSkhMS1BEj4XHBa3X
JbhGYPmZLwn4W/wxTvl/zOfwxptr62Q+2ePs7pmyfllj4EKMnnBjr9hNQLhyJqll
Fgyx7Bib+WvWkMW/fYQh/WIoAFUB8dQbE7KNkToC8iAcX3+gGBc64YP6Sm1z0hpa
+QY0xutA/eP+FszoSo+dHUgmtJ7/cSeWRAMHLO54qZQ3Y1Xx6PpitNPF3FbfroSu
h9Frv4h1Z5IQMx5sbr+vxWF+xVJEKv0T/K3TIUDLfvMiOAxUNzmXyf5RvyVXnb1L
m+r60YLLVl1yzmMVRSqxjLouKOdXMy56y57lCmCi2ofs5w7QBC0jso7rmhZ0WxM+
Tcw8+2eERxFq9OstBUcgM8jOoAfNCVDRjHkhszfb+Bju4oS/1eO0uTMDNBwzzV6O
QNboEr0CbnhZ+29mxsRYc0fcqX/NLvqdUUww5hDsMjDp+C185Sx67DiQUiyodgFT
c3fkXcXI3zYFB/UdWXIdFcpqWnGitunx/36apR75zFnhg+rcByxFzXbtb83hdAv5
t14L5fWySKaGLXwnWKlyZSEKBMmNjDflWN9FQwic5jz0kdQSdahLXAp5G88ySiD8
cRCvuqGAKanaiQeBucmkD0Ygalj2EkbqC0GOe7qEcqK0tuML6VcVveLpbLXPZcqC
jFExMRr/KSmvrbSJGWIHWwzSbN5HODFJVEl02lYvGy+EB8DJ2JNDWI3oRVsIg8hf
e++Ke26zmeeHg8L+9MnwCtCYuCZMwYSBoC9U2wAe7mx4HRsPTdDp/iSPYzuuntem
Osnxzq4idUw+vXiRURabhcWjDE5EsJHhILPux++fjxB9XzqBuw6bkEXuZsix7vxP
FVI8HtPrw+55UvpwPfsJandoV7zEjDzlLr0u/dUDA9qd0TSeZ/NlRJiinKUpTqsw
FbMjOkPxJeazbublSPsfhhsRJU/vsIRzVD5RNo+9azkvPVTE/ehwjL87AfTatkHs
CQ1qzQFMx72cLRxOXYf7AIDlNvM03Os3KTJjRsRF321GRZqP5Im4oiNxrEREUgYQ
9bVIuyVQ4HLqqiFPZ+WD3i2IkzH2UpnCdQXJr9L7qMWUj36PMC7dP9Gpfd4i9zat
eN1DqhuEHXfbut75+rEAocJXZSUUuarKKjyg4cEYU5Pf+eI9QqUJXCMlwJy4zz+6
aVwd5r3pvjPhOAp1IxsxZdHZjs+GBPc7x6s9cjt+nDwJvrPQtt/Axg0lT4z9YNPP
kNRGNf0uzhHjJzyM6HeiReM4N3o6mx2ZAEt+wxEcghAffdzS6bOmvgnnEh+EeaHu
7vheuh86+msISFdFQA9iIJgfR9et+ts6KUuYOU7/vC0ts6LdCbghWW44Shv3zt+2
IIuwHZc3FFa4nYkfUKjD9hm0ibTUuhRL82OskqpOMeUrkhhIXSDKhH9MPIoGG+Yc
KPI1x6TdO0K+nJoTJbmnQGUtETmPEUUzIzUs6Ti1+HuMN30pxGA3b3PpycBztGTO
5dNRY/Gj9QpX8lNO5vlzBu72p3Qafw8tZYLtFOmdWEBv8wGGNqC0P/Cj0iky8nzL
/mqJbAhejHA+iszSYiVt5GD25y6uK86vdPu3f8P0JUXbyM1wCPfPW347tVpHLXSD
IH1H6JIWFAy5uBhMfr5GhI1nEbFYiONPJJ/ccqPQmXlheoXaOFV4wM6WMxpC+3x4
iQydvJVRHSu6j2DSeQg8ikw6ACD8uL7kSSQvhPL7eS+PBnIHEf2d0QDvNghA5RgF
KTjk5lqQfCakRJg1vF35fN987xAcDRik70G2pk38RnBYTy/X1aeTe0bVRjInwi6o
JT+xzYWJPg8tGDfpoSJH99iPXOmIjcDaxpcFeCmQ06zMIKfbUBu1qJOU1M7ner5V
vIxRnTzl08f/UdT1tMz13Par6JRUL8goxC/2gz1KzKmBvVOaQJgV2Skptd6By/yT
MJoodocwMz2BbbkfjR4riFmRJfJOqP4UoCB0GDCb0J1mVRacL8iSsx948XPaavbc
1mCB34jmXlMAywkMVNZOPltKSEO2R5ediDmBCNxbFiU+f3+h1AYFG+C5frd3x84r
rRDRgHssQ+WqmgX+gXzV/qEwoEYeo0F+f3TzUYAVWGgbQDnCDT4kXmv0pZEsBKCk
qNwGj7pH69KDH5RgXBTN/IquftrKJS16N4NSgQhhim8nfBjomEWXmt5ZYBmOkf+P
nf4v2LTaZY0/jz06cvaMVZKdDfzpw7xJ1dLMlsL2RvGy0qupVbMdpJmh563U/CmB
F8cQxKq/F9utv+1AN7ioP7svfpF19ZGSila8RZ6mcSD/XgJ6CkvP1mafgn5FWC4r
/yyb6yKlaAkEojsY+AfuOjalWmStaL2jeoYZNa48O2k6kxvl2seIq16+fqTVnweC
D0ORk6GgCK51fwPlpiC6u70Ed0uyP0pSelC9zrd0A1Xq+ilC9vZSJ9/4wjSWDKSS
skiKmWgjZadba7UvhbTQI9szBhxstzEWdM6QivuzmCAlyY0ER8UYeShyk5nyVKtl
7IcmEtlLs4MmafGPPXfmYa1wkDg9pXweYxIWJ4Ndqd6g4MCG6SnRvuH5KNpdKBxJ
z9t3DguWhvtU8MwYQxreGSOSoiFsszDjZBLFn/z/LanFqvQhVzI8FscQMSaqpTRw
wB0X/b9asXszCbnDdrMU3JJkT7JpAkf23OQnBp+e9xufboxqiGTJe5FXQVezNtuJ
03N5n/qUblsLEnu5526QiO3wX9X3Ivv9HWapX1am1ZGUpCPzlsO7V1X3s9+4sAzZ
7ZNlLa7DlcWC3NHHLj6eAZuNAX8Icb9F/UmhQoONosog6CyGyC3pikDpwnefO+P7
c03TJVlRB0qGL/rTWWKWjukNDL3KhnWsOs/ulE85J3ZJsDGK8hWSUJlKFXmp1Np1
jmaBkmj9/va6dEDyIWEXG8801r/tRrtMtEjfcDo/gM6ZzQlcv1jlsmLF8MougSET
r+rkVR97u4Z+41lwa+msGphHCsqpiEmjpmsbRW5ELUab2IlbCqFveCgq4bH4eZ2x
LoPW2pYvfM6GbPw1egws+wdt2rqz1E++Z7d7O26OOHGMKDvEvZx8eQuPgYE31f+9
RYai1CmeDZVSwpAxFUncRYJPhEWke8lxg0bzi2k5e8iDgQd1pjPolJeUb63na53e
u/X55rwm+VkY31ttxo3modP+43jJ7yzAr15DdaVcPh7eGNN0/0KHhda0pe7rz4Vj
U5BMXSlxxBPbYDxp5zXky3HPDtjYrtNkKXX2488iuukFarAQIFZDjLS6nOAzmKEJ
DLn7l5c528ZfYSvdr2oM+sr4xa92Os0NA4dfMQa42HPSIKtwmJIIoulBvYxYrUUV
u5oKbDCVd7BLQ+II9xzAmUlbeTaJm1XktwwjrhmJdJdfeBDO1bjLZ9HBv1+ZVoam
X9HmRDwkpi1CXeFERT3vJSck+eOkfnh/X/P1aNfLzBcSzbX2D0xIrw1RWBW2L3p+
Rc72bm0qeFHIzrmCVjoJw2axMLqoaCJvWGaap4DDfnwcRxgawBu74efBLd+CJDiA
oDdHvsZGWPZxJvXt5WNJArripRoNndof/yPBPIzq/2Kzy2aPTHxPw6Wn+sMS4jEe
Ymt1r7CmedapgMWoXz/HeirndqJQP3Ha+jlnVNaQnM9Pxo2x+4Tr0OzFqHLkSDz/
89upNx1BWDVRJj+Npsz9qRhoESxZh/gTQTi+lAbL62UHnayzAWlGHHfnvntkE54S
VmSFRrQUpMFLkf4BA48LmcMcVEHdjpcySbCeBdd6QXLLRMRmRfhkW1TUK7eIGwHp
Wj3XzmrDzxL+ebseKGlqL2VGIvN0KCFAM8RiRgCYtVU/h+TJxc5ZJEfAvL1Nekbw
UUHA4TYz8UHtl7KovmkIaxrgUZQyGp+B000z5K17uBHHrrl/fFpXSYrgyiCeRnbF
KOY10qKEvxJhaRFYHhdaKaI5WkH+99tTi5JbKAtIuOBkTPIfbf162OoJhm/YCiEI
GQ7Q6wg2tGG7Wig1V96Yjcu8D8srqTH6QFpM4JRiZgMdh057NsJGtvFZMdjM3PTC
ouxzCRa1nBDrOm3iXr1eZyD+RGF4UHd9rMpZsFGanmHR/NkRpKfJshZYlenQRY9E
ThfDKKvlFLLTfT/rkjNerxQqNJ1bNg22dxs5XlLFjur7UBmWWF8bm/riho7QpjPv
d1wgdLlK47EaT5nGhW6Iq2gDVIwdfxwWJCNWwbJ8szeCABWGAAx1Zw1g6mcxHvvr
lA0pJIrfZ7rrRWrbEP9zaJ08G6M/ResYfy7c8vw8He0+YPB0RvzWUnqHaf8VK20W
1UoXCTaz0OKdTRb2ZRSLwj1lenMfwF44gVr0nCVAnTUOCpcjZanUQUYJdCiRfrr6
ZKJSK8u+m8gDwpd2q3nz6zxRrxkRFjhl7TlQWZO7vmG6R/3VaXgHjjllMVbCPUnU
NlCLdP9cgq3+PPnGqdFfyhd+POhRo7J5hEm2+OD7EvG73IaZxJpAXA6TXy6WZCNF
8yzhTnl81zbET/xjovxFE7dvi1a31S9AEIiasBJHUi+fCq7rXXAq6hIKwPgI4ri6
KTHlTZjdfwf2aa9cjx0hXTHwXS49h/fy8r1dDubPOYxjfWwKSrkMrfluZkt5FWf6
AzohCk+RBEGXnyJ+62JxcQstk9Z/4jSmU9Ak/TcE2rvPPRs70OpvmUZ/d8WbLBGJ
AzbMU8jPjggPGG8TxrEfJWTPLcuBbulXGzMtW5SDUmNNybY8M9nv4wLA13yEe9Vb
fgKdJaMFptDtz+3LodKiDvqcN6UVXfiJJ71fZNiI9Fi3hirbbNIpihlbcGqXP/bm
7Ao0D/uYmCbvS/KDHThbuJbKvDoP5IQ/ICpTaI11m6EzcoTag9S3XHggb4SJltAu
sqKEoNbwnQVt4DX++kkrLQF2IoQXIpgu6sjVcog5VQOK9goTJypeiN3GU7wPlAgR
hP7hxUhTt+BxwHW2E72z41Q85b1OjWCsyVKfMDyKPY8Syukj+fsKqDnR5zDQjln0
iNT98HJw6zsrPes8W2fz+XtiRfGnFQ7KbL77kpBEBrmdkTCchtNxeADfqhXIqoQ4
ld5NRsh+lEYQbCgO4BabOGASiZUqtBbXvoAoglUgATCjlcX04/RKl3Dm8lyRhvJ3
LqzqOB6TF/8oCyvYQ7Btzryd/4aR6FXDN5yHx/dDBkk+bPACAIJl4hIQl7TINhYE
LpQJPc6JUwPxbX1ISBdvo4wQ3Ku9b4WBmEw9bXNmSvjCvSyLnkkwbd9v/BYgRNXJ
zTQhklSFsK8EYbB+2iMdQcmJNcK07oTDgr8X7QMhQyi+I7iv/p6bdBK60MR9QB+G
JTvdiNyj6IAB0BZdU6c6INlvEaVPu7EXzs+315MI5wuaSyYN7rTGVfZHQHHn0pJb
V5GGtqusdtUhPoY1g5dXjdU1AWCAfUCbLsg5BvmwZFLIGbHvuUPksMYZqMmZY+xB
fmWU8cXuHD38u1FZJ3RVLOcotagOx0Oclg1NinOBG7I5d6r7j0JR5ntMm+Qg/sfT
xwv6DsHLaU3RNGWhU9sxOiNHynpIfFw67ea+UJlewTzxPQ96Ibol4QWHWxqhah/w
7XpnA7EWSxscglG+km175kqFYa4AcZvKEnLfLIv4cwmxgGSOx+Vl44e/MpRUwKoc
6frJkiQHBT/lSMlyt6DIrHtyRkCe/lqQF8KYKc4LPaeizYqorkXCvFijSSop9bxk
nQVk+A4+IGKnAF6V4xdbY1wHOHQsz5tcUe1OOfMznsGhExqxkFD28+h3AW6+Z++4
bEzbupFs3LCtNjvLhBraD4i12jhnZWAEMZfORr5zZcCHKfVQOKJrKK/3fyNfHg7k
w8zmeNFHrTJBMYfOpMfJFfNZe/a16xNLXWAUkXdYFKdUjCtnO2lqdpXh0SpfFExM
p4i4E5cjav3VEbIfGqj/GVG3s3BCH0e6vBEj4XAZ+t75HLpjp29VVBhjpIj+r8Bq
hy18QcoQKlRFftabjuK4thvL/isGr/Iahu2YFAyJfT4PFmMDEl9QgxUEfA9Omcu2
aZFXOza/A3H6AjpgHJig0QW9oJC48hAEXyluHTyb65zxPCvRg0Qycog8ZNeZoFiD
V/4A/GzPiGg6MTlGv4/j/lQNdhML1tBC1cr2e3y6k3p2RxP5JPe04DgqESPHN6Mq
rAa03wujmFjzDdzOADdeTy0Qn+KPAcOiWvf9MPKiYGcLi9LQ4vYTjJuL534/BT3O
BMuhoKNSNER+AhRG+js10FymROTcVoDSpxnsSCSrTpo+0DJigrilMbCK/kTgPQpb
tJ+TVXg1iF2fDLGYnFPpaIw4+v2DRz7lzF8jSOLJpFqFWKpIXwaNtyqBUC+bp9wO
9ZR1Mu/GyKshJ85OjWP9bx9vXcQw9YTxK6PNlJuDc3cY2KB16j22HoPXpnqfXaK8
hRz3b+aUKoh3dlS03UQwbWZd1pKAlbIF3LzVMkIP7QX+IqQhWs/ftcn0d6t+L5Kz
NKonBChl/OC8IAz1tCTNrzB92shf2Qz7TxJXBRUKi5cD0Y0+9TruVaNJMa1TTvXJ
kwiKTJQQ3dhiTRue6buOv/ZkTlA/nX3Nc4mvKm5ilxsgXiVxWlwJoQj6nD03Kt0i
nvd/7W2gJsKNm+Q/FryElji2fhNcuzeMQGG5GZ89v6UlDBtQKirjjS1wuGyTCPPp
48J7kWjx05aAhgzGOjgypnesbDgM3k8UTqiJQVnJvoFfqFk/l99hW7zUUVvlifVs
OVcdEgJ3tMPVQPjcCiNASAIR6k+s3nacn5GSPqkvmHmf9oAXbh9UQiY5J5QAVhfl
L+ztKaoFISRyz4eZ6cTTpXkjlOhDu/oggxGwvVE+NVWM3uEKDZImlk9TZGZcDheG
WHe4+qNDw34shLT0vJBnmTssSwEcuPpcKOpCWqI45B7vJQJcRiQwJsmHe0tWWUEa
d23p3RKo2GqSsq1pyJAflOH/7L7JpwROZReBoNZH4BR1KEPU324bCy45Dc8A3wWf
Z/Z+jmLqQTfImjjKuSjFyojVaFWsj6IjDaVXA+g5Rrs2Lk/q72MweMYTZsVyaSlG
pcG8kQAsFmBxHTatuVNQBRvidBwQ/smH8BgkPVDHQ4lfHHRobkr+jO7D0Z+duS4x
fGzEL7aqN/t0RaNb1hIvtg1vr7gEIRqneNy6rHDVVHh03CuAO38xnnra9S90lwW5
rb8MX17zvivZCbNw/sJ5s5+gdUkvIXw85AdR1ctQnvjMEvG45O9Nu+raGSqqrxa9
MTus8XbI7koonv+Y24j4mFvHmkQYw6McxEHAGfPQsDg9RLE4HD7bICzcDF68TQQ2
AKFS2xO+wjElEE6i1P1bHCFkt6jVRw00M5xPHiMeegkZwtd8z97h+pTXb32zc1Iu
Ehu5neb7qr+tTSxX8z0cG3sxtaefhUgbck3P+EonkvMvfv/g41UW5xoF06yemGyU
F43VyFziaNaCjvvGXe2mf/Lw7nDglZFlpajbXdX5cMu3tLCrrIAeRKsrRuZcxkHJ
bTIZ8XxaYYXdOIs6VHrxa+8+sTLjm4GMdJ2mb3p9q20dyUFiPlfJLBeCiwkg1Xs6
atbrvcYHpQI7CQn+a7n6nubAvIuspTCB3djSUH5K51mAK8T77e0YDhiC8vUoBoE7
I1kTqth/0puMeQZOA3AxrMk7w6FjXtL9lx8aoYTpY3J3RvFt6SeVsUP0jh1u89+g
3i5NMwmj+23ySScGnT+b80e2vTKZ59AtlD8TR+BVjExCM14oMNYUvm4DuA0dt5kQ
62FN3OTapKdPgybqL9GXIIQTFV0xNHbZq0GhhtpRSIydoi4dlp/+EzZkKcrzuM30
gk55Xngy9xbFsi3DKRXXhLh+x7H9Ur2Nls0IHpEbYgpezU5BBRuwZsPhe0ll1yZP
tp1b2C+l/cAtqKA7VXf83v648MaIZb9X5ZnX+bth+yc3wQn2MW5uhE+lubcnR3dV
3xR7PmMKdpsUuuf2cwoaqj94Zkuu7J8ZJhra5QrSPF0jPEadj13vZEJR/l5pOAns
S+USTnX7HgtBYglWyiT5BFVcvkFywzsIiEphH+0uBMTiA8b1PtBokdkM0FVBQuaA
ME8R3bI3xzL4gyPMDYK6fXlJbsF/55BKBweYCbi70UBoslzfa9A86Jw9fB3Y/PrJ
GrPmOtgRh/y0FCm7/u4zdczExNSy3J/yO1ZWoF32cIxmizTsmY8z+4Ik/ATnDzdl
MLdprnzNwvwmzmTvQe430x0sYT7uV2H9AFKlyY2s8Xnvt5mCr9lu9meADu+AbotI
t9pn1XVP3eenvWiNctyx7vb4wiacTYHAiIcFffNn6odVSM8J62FYmiiYH3M+Fm7k
Y3+L18L+9ttDi73gRRSG1fHDNPFYb/a35QYB/bsJ6qO1QeFNV/9iQdkyPI4s2auq
1/FxuGyoWkmYoLfD6wk7psw4dc/4kiyU7zKpFHdy6CVgoIjaFpsySEYlaMGRgN3W
NEHP0p2TZZDl3fP4T8INCw/8ih9l8+1WHe10L9QEdHWt2hr1C+WJbGOO7K067Ycj
V3CZl553qi7nyzDV9KXZ4S6GWKvR2lYBfpVnT83wLPQkUIdbHziiFzH684HuReGI
gT4WgsG+bYSASo4+3/uGMJIaRwFDIaZekLOqJ+LDNzMzmrwtIaHTnCzxyA1KUne8
M/Ew5qCeUy7ypTIyxiJbL0Ph2ZE7/wb+0HBm5uGKROO43BXOYCBalcBm+SS5KKWo
wk5xk6o0MZYMShBWTYGho1KneTSZbdulO5oMcGfA5P/v3GPnVcD1OjXgWWMu0OrK
0FDyEDNHqu2xlGJsVuhGQRcgIcytggIW7gGE53lSiI90ol7xjbwg5Fc1UMjogVMu
it0R9/QuDXeF42zgMrdWS2vl+TYBd9XZloqAEEguzTwEk+Xlm4bgPU14o0rQA4sK
Hi2Lw7Io751AtG76PKPcaAlGMzpuPVluePxxrh6+jof4BohjqGT715bSeFx4lq//
Ki3edtU2DBUIR381aW1qM/q0uX/DQvj28zeSvrW6GgQhp+mltvpeK9iTtdLEc29M
JbAM9sLSxBdp8kk+F37FvjK+Sr7NAtLy2SSbnnuH3m3Z/T1TQze8hDlwQ9/bGDoc
erOqazf6GPlN6TDWmrUHM/4AXH+e8taa87xJPg3ml3spd0o/QpFthJQdgRnbK6mK
ruwisdbPPIvLjMCXaXCa2o8TBeCRWooZBHNJMWDTzDc6osuEgOywwEZVyiDAe0CM
DYp2eRoX+wUm7qF5vVOSJCxUYIeNU82AZaI7FlFqrh6nY0T7dQz/0Wvh2Hp6dmVz
QLgDga2WRIoamcEgrYcg37qs4JYZ/TnVPYIC83HB6b7FZHDom6XAP0NIKTT7e27E
ctydEGNjD3heqgdOfcHQgsAHqI/shaWI10Oh0EllKXBWoRiMusB/OICn2y98SBI2
d5Pr0NqzYKqn2pkku8g/DSkavYJxU0iSaeScAIyLpkY/WS3GN2/KeKCUaaJB8pHk
43GFvti16QGJPtWeobp6pkZ3tzIIOZ0UQSjwIAmscdnARstwseyNeU/orYgqKz0c
hiRQSVeKq0uJzoHkyAbJctQMC4HYY9tEd2GqzIZhQpTypWgTQtDQJDgL/ToiBYap
0PpcBWBDoq/UPE6E7RT2HUCcV/pmHm5GouihfwET9Ybn2eDtgy1wgtCWdtLj3KrX
GWWLwO3U+26PQrJ+5DTLWVGBM1B7wmJnZ9+Bn+O44wvOMV0Y6nrGgc871EXsKgVV
brMkLfrmy8iFIsxBN1GLDq4zkE4yAIalr5TYGiePLPOjKr/DZbK566urkydUBBwn
od23/QAOQuKKNLU7ktweG9Km0LDYOy0j4igf3hsEstuoExW6jDtGQCL7BlY+CkmH
FujDMRW7FGVA3RVI872mfvMfSFHPryKieXBsQDjWEuRi7SLmF9A1XF85Uuw0AIXw
mZz2zUDZoUeyTH96CNrvyKuuk9KX8lff+gHAeQBS4DMvL9Zmhz1D+nnzF7NUCEQQ
lXRzFBNUpHVyAFcfS9d69hdERuSc92bOLlmfK/fh9ecyfL1CBRMSe+FNnGfHJkhW
x0zD5h8UNUR08AmxiwEFhHUunM6f93suoQdmP8mveBRJTRuLN7DabbWdp/gb7Dv5
85gQrH/1denqofYsiaAhL5Gc5MGOOvKPj6lAkUI6KhFrFN3MpRErpVRKJyTwxDiZ
1xhH6c0ptDLwnbdLXmvUmbJ4DsO7nGbWsr5E48oy+R2DzRVOfQSockWrA7T9hhTm
li12WIJk11DM81oOFJ625Djp/HUSfans0r5m/WwprCXgzddnEZmM7gZxMMMlqZS3
QLriXMErI5ZzKLkElRPEK+f/JKovQ0X2LCh1mSfrg8Wuc8isxTi7IpOcJxFNA8ds
VFHVZwEJowCxkedO7CyEGIRawDfdP021HxGt9KJfaoqAB2KjS8JcO3NgyUtUVmmM
EqK+/zdK6Sny7ePaoFsYnjagUhri531ofPbxBX7hLx5Q6rActxShMCItY5IglCSI
Z2JNg5Hz3GKwaYW1Ly4OSvMbvvls071JlUgTTK9DcQir6BPJMbCkqr/4qKE/QHe7
207H8RuOmimb/C5zJTPUTWrxBUYV/wgJhIEL8N8GdZrgyINcZBngbTfhF5+ZBiJH
H9b6T0QQpG0DI9wSajZCkwzjszZLABxKFHXdSL1hFNGGbI3MDwPJVT0uB0uwh6yb
7WnTQ1NMtudeDafZbmtHU3HZD+xEQ40WqG5qyrezw4BaEv7KbbxGNgW2Dyc8eaHI
44ZQG2Eivf5mp0ABit+iIxj3RVybKdjnm8TXjHnU+oUKaQ+VDOO5oeFPKFYoQWz7
EAaHF+DXKO5i8xgflj+pekzNsaFLbknNQ9wrXg7SSnLdbkAxIK4z8lbSKEu1b902
KXBapcxYQg/f3rPcYy7RE1hyJUGhrXIW1Sxlh3TPKDffmjcT+E/qLU2WWWDTBlu0
644/vHc4Xudnlk3mK3Ph5A==
`pragma protect end_protected
