// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:39:03 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RZa8g8xH/+7p78r2Xqp3yNn5O5sGJ05apE1CZyh4w1ygh+I7M4R64akGY1cm4uGj
ZgWLDOIfreEV0sWAniAdmPVIydc0JMSK8Bsmj9ocfE3P42NrRKMLuLIqK+nojCz9
gmFrgqDjEXWV0+Typ3QR2KrsDilTlcoO0a4hVKL927Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7984)
4CnGOfWi3T0cIWugfkURPjy1h9prbVggxTtURKa69jTFDm9ckS0ZhvhANMwj1zxk
pHRMV70AKUlq8F4gfjYRGtyEbNLRfU+kok3dvafGS85JayrBFTB3VlAyb+wWKWhI
WsDh3od6i43on3r8DgKke/CM+s7+7sHtA2ts2Rpf1kciFGhX89PlpY8GpirLvLfP
7j2F7rVG1X66rGn4D7KRtQo8II1nT7fDXxGxDDSW317ZCte0K1zVik9aBEEPlRNj
cZTCgDd/PtJYICQo8k+qWiPoZp7mgWIoD71sQXqE2kmwCwL0HuzdzqyX4FArxvn1
4hf1BV0XsWTKqI1wp0vR2Xn0jAkSboyDwnmYXVD6aZtvi1iXfAF7UgVQEz9hHgQY
yTq735rQI6s03IbQMRkkirgM6jNClybZ/RKcIUTDX5JB8On5B/1XJ/fmHY/+S7nz
57OMZo+MhnYbFe1vM0xqCMNe79DqM05G9E4FjrDGf6njgqaRMo2xmqApfstXwgQ3
AXWLSXgpAmytaVgw40EDIHUgPd+DOaJwM0NAZ06TVl5hrmePIk04bOddm0Dop9TL
racFoW8KZXMpf4ae/gT7bJEn7quBVeQc2E9fSVJZT8wp8Fmu4QUucxDXF5bgsLbB
Jlho539AGehhh/Qm70micdSarAjk5WyroIE8H/hffKKMRiQG7Ii5cEY42WYOFkoE
UbczASIXAYvf67VOkVZiY2cidhRsg2nNEmn6shzirugKgZ5fu8TPW8HFpWy5HvCM
6cCgBzWTUpAaKRvjltkQ8HREY27XoB/ECMsDm6VHLi/4E+BraYtxF4Tc8YgupGqh
i9uVqeheV+fS8YDbOiJP2OsCePJsYXt/2rws2J44Vu+Xz5CXDEniHHOD+M+eGKQN
66AXwFeY445cHndMvbEz75rnCuYKq6u6RAn0NW/z5heRhf0gKg3BGcwYIMgQ8MMh
yiaooFTLNe81aHEnZgfsfFFVVF9k60r8uKpKSRd96Npfhz6sqTmlp3yCmNFd1ZC5
Z5Sp+HOM6x84VAQ0VNr750eTsOFWFuvjENnBpNSr8/MVuvHcxpRtBld8IVoWpNhG
ohs0jUWwxCrIyrWSyTt1yprHaLglPdMz5EIw8SmW6ewi9CGPCW+laIc9i3rNEGA7
EdJT9VXe4E8wV8wz2t20MFWSJfJ4Hz9ceTmWYlPdf1hm6zaG39Mlp2f7UrOP2dA0
vIWnTGbdKRQtFNf3rsJKH5T7kSS6kR4xnLPjoPB+zcHLueIaxn0hfPO8c8cISu+Q
0yxepRCMmbgmSK2bBJK5N6PkN+jYa9v/4BZR1Iz3gMaL4XEljqwub5XC5JIir1Yl
bHDxK+mFnlpyBCNC71NPYJ2R3eMdQcekxjCxBK2D8Ve6KsGSR8Rr+sgVhGJNXN/N
UI3cg6bRdDHYAdvJALdD79lgKn0dPFwR5QLVbktwnWVNoZqeFBEyr7Pp/70nSTxe
5IUIjbPl+zGUEiTDiXZJtISuMVklUK57UsA8+DXRwZwRjN9JC+wAUFSj81/6hIDY
e04yKpVJj7RW0Ur7SUPr745FJpHIdmeVQp+Mzcm3OBNuyZDPfkHvgmTA6DttP3tl
PgJ1eG0F6If1+jjThL2PNPcZpp65HpQfbaDzZ/zfZ8Avysxj+ZDzDIKAtB1BcdzF
RdLuSiBaWTufFqzsLCvqRz7Hj7Q8S8/qrhnYSQ2bgH4H1iGX07DI3G2IjjjgMnyI
NflKJQMIfqKrlkewTMmkCo/N79ws/WUlpGU7lU9IDccak76QW4ug5YgSHs3EZzEe
klcm28TV5oOxc94yx6F5FAwQJDEkglv3eEZDeG1DagAUHSo7uk7Vi4ng0Zm9zHE1
3q3OuNorIirvQAUdeJ+wX6qqM2rQaiHTkwJHF55tEYYJsLN5jureduuXmcCM8Uvd
jjMjJgaGgdWjvz3XeAGSsvdjTrLnl/SbFJKqBXmCaTneYcCMaubNcwhPYbDVC0Sh
psTmzpZtu9xlcnTjCzKiv+EZZNmefhKlO3XCiJAdUw8AbuardERPMdRvXMXouYUK
jnjPOCJxMzWK47hLyAO7a7pFx3p7R2Vy8AuFj2d7bfRwosDTe5PlA/qtXi9hUrKZ
A6wPLXS54tNScDmkZ6+gFYm7CfpP8c8XD7WAGAEqziKXPIppmJD3IOXnkXsyGF9+
Cjj7xw8STvlBZnKh80bi+LZZa53BAsebR8HhttKI0Zvu6fr3xWJqG2hB7zXANydi
wITMIQhm+Yh7joUA4N/nfc32PHVGqMcngT3PjX5umuc27UpJr2qU3gx+2uKK4iso
qJakTMM4RUZ4tTFkJDBgfhh9k0OcWE3pSsS4kMe0ItZ72DGngnH8KSazbEiPADwT
9W2iU2c0S9SRPM4e0w86i29kK+cI3MX6J5VxaHisktgUIbu1nfGJ8EZ6LNU3DKGz
bWE6fSptVri2Pk/ixV11M9EOlKTIzVnGRBir4c4kPCcBvPMAHCjX3Dcbo9sFUKoX
7rG7neNnxNXRw5veNShdacwdr31WUlslbV/PuoEVb5v2/V/YbinuZjYigPkSx25A
HElpifdA52aDCHciQ/TTzWjwjwmT6ZspLe9Y3zeQfUMq7Qc4q/SPnPDzjJoAsSMO
ncdyYNiK/zEiy5ZOskRh7reqzs7vBT6p3EUIeZqtynbUJiRMYn1q7eGMd95M5Y9h
lhWS/zy8r65WsRC1jyfSb19zZX956Atyd9SR1BSl+1Y/pqoIvaxAbJgADgMFi17C
FWgMY0O/X2KSlte0cUse/Umzei7uhUopW0ZudAXf5zajdBvmoP/MkpYEYvZBcDZf
gprJgjg700fxN96ZD038oaRMkp1DyvOg1xah6elSxDWtD5CxwO33dcS/dmFQb3io
Cxfw763ZKNdOeb5O5FFGBhZMVEsv/AJ64SqhyWqiiVYPT8KjSuxf0zcL+q7kO1aj
97rmeieCbqYwuwP0zWAHmXPfUKf795LmkuNbY9bisB1Nw4VnBPiWVaXics9HKZom
SRYqmBCInwp0izWrc0xpode67+Ax9dd4r/8asGYD6JUfkfjd6AjTGOJGfBgv/qVX
BfDyD3N5lHuOPjrguT6XSWJ1Aqk4HMe3MrsE6xEsvJU6UXArQYwcjOtcQkEOun5X
H0XNHckwH4QrxLOg8r9LpPIyHfNEJEk3jYe7Qq00ffXPDnNWjG0vJ6fgM5xalWH1
jUNq0HOKgOwFSPTPL5XswDKK6mVrsaIcK+21LpjMU4NWG5Y1+JALJqhVqd8uuEem
IOxWyaUctij85a5jLhpf+Ospvsh38Y/8Izq50ZEx5F+2Rbcd+z52QVmN1AlUc1ov
s4s/QtCaLVp5TdX7fzAHSqhMWZATSgyFeIPVYnvQb69zYGiP4IF4/dJhxeVLHX3j
KdP8GexJDCa/5ersItl0wNU910UKk3ZBQ+agH7DWPLHZb48/QgaY6NgJWqDlF9+a
Z3SjidHAwAzfgrJj09Ze3S93jLDCnGSOFirvz8fq6NVeLeNfMnlywAQozSETxmmU
yKdfI06McLzTX6M+xnS6VrpM0TGwC9JZGTWQCg+AKdm4VnObv9kkOcMAmRLuxwaj
2L9F5dUAKAYeRbgm/7AO4wN7W3NixTOv+ycpF2YTqkWauww9mV7YRie31vZc0iz6
vLBmQ9QUzbNw+LMlXHanryeLBU7STi5LSEA17PvAI8P9awlYZ+3O+o7DV9dzOn+I
eDeuXdf/+9yQOyhf/Rq9Q8m5r/ROC5l1Jq5fJkGC+6F9my6Xybaw807uNWmfg9AW
TQdxFt1dlUqGHrnYnLmwRhTmDC2nr8lAcOnNBrDAnr8X+SnpZ5Mmyd+NrRcwbcej
Biy/C4ZTXMCkc2ob3gTDerme20EBqOd6GRAh10uZgV5HdLDPvbceYjo/zatekCLI
x6uo+dIRHBzr9TErVB2eYAueTxIyAOARD25TRiTKqYpvO0HQUcMde0FznWVkeU3N
spUcb6eah0jDKJSRt4Nx0w/HddqfTuziqgyvCN9YG5KBdsKfNoFGYkw+IIbuwRfQ
md9cmIi3TStucV67fMJHAZ66JZeKofLIUHVcNaQ9tSGzAPZ3makDuoB7O/SKSanN
K46l0miPMLkPanRC+sLOm0Pgem1IgBR/Vcye9Rj3ZB+hiS7T6OfQkZ9bkWuXqK7i
paCe9ZeBZiKRtqcR4MpZhLwjD+W/r2ElCPL/DypMIQ3NfCH1OztyNZGSXBeteDY/
zf6I5wxA4Jo7e07xeriO4RgjbqZyRHseE/p+Xlc1zDQjFx80a0bRx2UAnl85qwIL
P6MeHWvmu6F2BJoQTSpoS+zCgViOvg1Y7c7z0dOKgZwaGEN8JtotMUUktRaFtjqs
T/FoWl8JvFoVVK03YKaQGPtbGj5+aElutK1p0Rz5usFZWRskovTT6+2oWph5NjSN
+GrvqaMQppSCgoZc5t/ZMIBMC56grfz2GQGq65Bb9y0d4Aq8qg/kQvcamXDPPDM7
j8pg1gVkMBpqBkgeqJujyIRc2W0GFJRiV4yEUhWmtdn2uqnMg51HsGVofMkjwmnH
8b1TN0Qbi2AXLkAgfdadRBMoL7OStN07VCRVnnxKTTks4UIW/+FDKFgwkLfpNGem
VDqtVHPeWnb1SI5UU7y80BuAWyEf/HfEocAfc4eBq+0OQciMITmGhYrdivLCGNTA
SvuKx/M4mjRF/pug7v0HY9cHo20W3JNQkq5JQE/qypMFfbJ1J/eE1206SvWP1M2c
CS+bDkEWMKF4YGLq94VI1iZvUBalVYOZUG+SvoDoCYjo/NKyuQ9fWiwUB2twzQdy
Sjr82BLHZE13GY5z8Vnbbj+1GGTyysXC0hm3nM+oE6BU/hs7zPjEHgGp7l1IM44+
2nCFofVOIcIuuX5VPR1wZcY4uqHtq1fMM98GyvznHt2gFENk1+mvwTQsk4BouDAI
2GwRmsLAcpOaK4sfpOsAHMIC4Y8oOk6QGJsnwCqC7u4YQVylMZrUgODK4h7BPJTf
ZlvKzmBZjssMOeMli9l8Q5n1yjsUNAmUUashfC1UyxBmUsQM6RRXbH0FoStURDL6
t9gFsbj/XZtuigPwGS98DK5lMT7N4RSoNGbdcFairV+5Sae9kPNzGwc0MjG+GKvT
sYiUzK5xyqQybo3ZtNKKRL1Rbih5X1Iy3F8nzD094mWGxGiI03fEmD1IRgcTEDTg
LnAnpguedh3HLOrfJ1ISPfpDbiDv0uRO2KL437hh2STeQjjui0Za803A8Q8bvf9U
b3qMlSdR6Xy/3ep/X7wrVFLJi4Y+6ZFIliQUeVDwbbJcNddNGqc0rNfw/0mx5i2R
8wQrS2PXamUKcf8usBFHfO4ikcdRdx3isqQnGFqd4ZPC/Tq7l08qRLr7GzVvF7Vt
Z47hmA26cOtrcS+LXwpgqevjyt8ayCDDxU2FAhEqJf9JYrfJozYrQKdlUMPTzGEn
W/KPLenARZoPlUYLKisaEXK+JFRZg0sCwank21Y8iC6DKMwmpFEO08J03AjmnA81
bfy6rXzke7O78wOSdBFd14MX3frnWHNH1rMCgQh5ZgwjFpdoruNP3mhNfZjPANU8
9S80LhYh9j9pSmX5QSE4mbhq+KAWjXQdgY8IDWqfji1ax2MIfnsxN3Rb0P1kYgTb
zko/14TjU99E52ReZYfySv0bhLPUZAB3i3lIBHcjqBU1q0L8R1nrncc9qD1T6mnX
qZdFNuoNeKpf8qor39VChUeN1tFZbVsSn96bXVrjQEMFD/zMIIratVy2DonbGmVx
LUSa8dKBwpC4gP+GsSXXivutbQ5p7zeZoaexHOJmJsvygOExLDMwJjBFHvbYZ/dN
qoRTKjrr6XRJKHsiudc+p4DYJKI212A+b7EYQMl0tS+JdHNQu0tlb/yvIPzwMg46
EXVHsj7EwBmy9jdox0D75CrXkXRCKezvZT7TaFCy1jne6Knkz/W4vb7Ga89Rsa+v
hwSIkskepory41IvKo5Vc6JDD/hHlriC9O4s/9yeeveiORD6+k/fP6PuK39YJUs3
BAI4HsgQdqnVp2WlM2jHk255bS95fQzu/fIvfIDnH+rhVsoUlAi4M+PUB+YRRSF0
Nd9Vw6Dy/gq/tQI2Gj8a1YLcmt+uYVrrxS81rGJlcbK4DcByUCU0MiDKJf3EGOSx
btpP/zOGUGtrXoX8e7H4IrM1XqIljJjI5xBWW8mg4MqfG4letOs35+SFcYly0uZa
qaBuyD0X9pMeZ7f8Zu4d3rZIz/ps/e3EyxyTW01GnHasrk5up7U3Y5K+ODZ1Ftv2
Cj2eN0XtnHtltp7yfKqrIO3KUpTH3EOU0jpa12Kk7uL4u+ayVR9G1Xm8MxHD2dI6
OO/cvVzEASyG/dX8FLE3d7/rO61pbJHleQNG2YUN0CYz38KKAxAlMOzPf+nrEe0F
bByxGEb9dbzJyRqegydK174O9qOHqa923HV3IO7A0gMhXkcALeLj5ZfcToDAicCp
XCHtyEcPyLBxlaA/3uYDikW66w+PRSOS6yNyo9ABZuq6pHg7IGS7D1nDOIcxuWNb
zUYxHBTnpo9lhF1ACRmaxBwAqvGtU/6vC2bWXFpEKmOct+VXwgNynr537uNx8P06
7LcRzhzC5uOXf5VIoNompokRBeiYuUabhZ1g9cyLMyQjx5takp2W52yHjuu62T64
BkoKXF2iDWLdsK9fuQXrggZFWjIwsKXWSVdtK0g6h6O97+72BLwpAVFb6RQDcLib
bNmKm/3dlDvseQSKRtyXIPM/FfO1brm33uKR3pmKjnZKC2qCa5USS7RTfbIrBB+V
ZzpZOlnEX57IqRVzVxtdWadIe2MLrvwUnMHook9x+YXfRUb+6mnvBevQ6cpKEMhk
0Dy1vDOAODaGLhZrqgDe73hQVTqof4LauCax6fOHGD6I2X3oWh5p5vdjkqcnlKLM
hn9djHb1L+saLY9W5cMISpTYDLhShdNZh8T3IMJy/XsIVIvaBmC+RUms5SHi1BIq
rc35LtW38wpmMa/fp9eLNdoOsrlBCchzpPpHg5w0zRak3EjQkZn9sROvQ/xEsAUJ
R4sFW9jTFn8ZXo2HyLcBLwhItuoliTLIXLx33fOzC2sPMMp6EHiOndR+KeSjcd+6
+8KaxxMenkET8xUYsM/KRbHHYBB/xYvcd4vzWyjLHc91LCOjV6WvlqsEh5AhQccx
n5fu8uMVyRvVAbon37WC27ojAfVTu1PDRKyk+uLl3vouCqWIaxjidqMk6XZey69L
zzCdyWJCScSXyvgpSUq+/aUniqYH4N8/cX2baDOwb8KTCd1sPrmJqNAv+xipm56e
GhuprI3yLl2/eA3yTqlmAh5I1qzApp7teR7D2mAEpDB54wMr3+HmOan9szTt67OM
ZlRiXCUkocQj1hYGb2lYfbRyXzsqfiyMGLqHSdyXHW6aUEgCsoSQGcbOvBRWnjGW
wdWJUAptjMNWOScqiqmjegXevEYBdoZ8GWdUvfcq0HEaVrmLVfc37aV/FOLXQtg8
fUheNZ35SyI2/xxloToH1nV7kTkyQDpqy5tQhAwRrQLe1QzZ7VNACCABgyxE5gVW
3Z3Z+/VgvUtB0BMF6CjX6Y9FTtXnGH6blIPW1UdzrfW0sG4O8jzVJ7PrmpIIc9fi
eWBX3iilpN6DT8TGGo8+C9MF45X2Hul6OQ+3QG2dbtT+GmKXhtUiKAwhf4un3cfM
CxsnnJTrfhFzWFyPwOoiT4XLhDfLpVlijZymTVXK2YhPLLF5WKPs09LiwCKXYKm6
Lr3rXbAi3bp4ZHewy4c8KIdxROnf+oLe73PSHZcKzjtXuJ6RH7nXURLd20lMmFP/
33EM5Z5VDCU8YWkNrvQllFwe7rA+sxAnLDz5l2dEM8QNuCuob8umF5DOWp0z+JeJ
f4xlrzwtZQwo8xDmJfNty0Y0RfGF2CPc+fPMeXuPyBu5hZZEdMsRbQhluKxcKcaA
qLxVE+aC6OAzTrFGdhfBDW6DA7dPGZ5NK8xVHAFvH5qHrMOqlFN+E8MyfU6wR4tL
f5xLjrK5eUCHb4rYCLfzl00PDin4uyWyl/0DZ0ArUyKxNRFs4WKc6rEVBKnxYNNU
6MVWKB1SlwOKHoGj1Rv10H3ZrGy6YLe5TrFfK1aUnf+P9SmG1htYwrUut20ZxPZm
/GhhtMxOLQo7RXdu8IArz8m8+rnv4Jrf43fXNn89LUxEgF8ppjNFlYdhlPB9/9Ti
n75XVCm6NBDcY/nkhl4u6qNr4VUPGqQdKfhrZrR/VALO4eAZhXbugEwSyqX/6ogP
tOe/aJn9ue2wZ2GQapGffcXLN3fcoigvz8huBXM/ANQ/0Mq0qhdGqKchvcTvYLLZ
NLwFXpEJaqeRa4o2vGatNwHZ3WobZkffunmE4P0h0eSL8HZX9QGlyBr6nanBx7L6
whRxv2RtP+fUr6x02qZjaaS6eqUi6N/ScpG9QsZcZzgUqZ+srgtXbQoXzPBa5xvZ
oA4L2ZzhrqpL/mzqKihPdWpz3ziwvwAuHhHvd5H4HO2TnNzUD0U/82KFV8NFccko
Q8zgLhwaV5rBmfzRQnCI4UOpUZX8Z+BJ1xFyAIwtJUgYZ5tpl02vGqTRvxrzz9ZZ
LMIT9gQk1mMLMB8ouwEkADd+Rme5AlYB8/Mj5R3gjCL6ALYWMiClqT3YgGRZncmw
kIIS9HZkB3D2IuZLACYHXGvek4JQBtKnamjdhVJharFzlMp7mdxjh8RZsY21yqyp
EfppNX4Y+G/8Kj4n09oUhGHFu5gZLqkouhqvVMgrPl89Wk6lsGTLNhlSUyZ2Bizi
PYWPQnFESYS4IZll+9TuN6xm01svcVrgBYNkq84gNpCywRukqVdPjzYVcFA97ev0
WXU94qnheKcFHcCUH4Gz6+WKzQERSu2lU4Wbh+b3Q45Mc0M8SsMMAmvQzJMytS17
xvKbmt1S5MMAxEfWnfsUwvw/9Igp1VoYekNJUc+nVvlIzeqFWZEzgy5FoRwhdUlY
VT+/2OXn/HoakIHSDvfqzmkzkw4Rtm3eXWyR5YAnDLOiWhBQvvZ1AoV8OxcySscu
0hUYuejeozpV04nyJp/YWEdimCqaKTipyJP4iXYhhufiTwiLp+I4bByhIUINH8Ec
qndZsVFrdhZW4u4Iu48YExN0NDPQgCcAyHKElqJUG36YVNZXWGyHhBnHWdwaDjdb
HmviybONcjJDv47km0toRFpyLEpLcDJHM3GvdVkYRGzo4Fx4M1fGkNxWhaYSid79
xVfaB/VF9bWiIIHXaMU0b9h+VKWx+2YT3NwWrjBLPFCKBj7iPXercNKXIfgWL5jn
64RzLAoJbbIwURNcqAFJilq/hZRv1dtJgPCcpovl8ggBD6cWzCNpLZ3/yL0W1Hn7
QNGHRUdcP8fB0UbZvbpa6A8mQbw6XW8UyGruOQh7ULgEZLhBDIkNSqD+xiFNwAfM
1iXVsoaXJRDNeAA/vzXypY8og183piwq/cdNSi8WerrUwIKnjJ+AEZ5bKG76d+ro
YL7LT7n+WZuAXY6ZH6DQVBNByiYiTeO8HL4YUq55s6rBNxxYOfcetPRsMfDhiqLi
Ql9p8TWucdSLGgAZ/HeG8mQncTOZGOpG/HazkQkTtRzl2F848E9PnXb2tCJLxI8r
sIk97WvNgDtKb4NtHbK5ao3s7xouTXevF+jsBtaGae2PqGgoVPMJhnfGDKFMUlFQ
DI8hSRHw2VpIhC70VNOIKluyrNoIMfX4WK7v04/eB9e61Aa5VVVrLkHvHaXsVhc4
FCcEycAAaEi1K32qKTRIz/7hNHV9DX0TFTEnKTzF3H1gl8x5lKv81R41CjOcHh1t
mKyMXJ4uPDr/OePJl+8kvsFIdYh9jKJRz8d4c/SyoolHbtEuV7JJArKXXGe0Oe8X
/aemwYfzCnLV/Sp+jxYfZiwoiBjSdf+lWxHefO/cKPvx5HyPhfm+xEa/XwfqeFWm
DRF8BkcnAyxXb3WyH5t23SmKgr02nkdg79h7nA+pZGFOmKXk4jWjHBBNc+/YOelM
crafKTvXjuQ1AYSLGY6Wzj56Pa1JgXYGDKDHbKTe4MZ3eBaFRj7Aj0GCZGcWkQHl
t3P2X/E/M9IyYbagbKpruy60nRrHsiT9+GsAUAeLQuUkAJ9bxhclbVYTvWzijuAD
zMF40rQZNTwGn/DQyc9BjLd0o1N1pxHDEHCVkr4zhAnz2rbFYFkSxTZcHGuX0vln
d9hHTXRS0MsfIXogInKCwkZJCMjBFFAVaCvauM9bTiLdtTZzYKua0OC4PBlq1wIm
2IRqCM+9b67YRwyIiUPUN95u9FRY2d2ZCyT4oS6KaaSxJBPP2SAPKPi83Z63RBDp
DHfs7Dd8RQ95NRf+DungEhnMpCt8rHKkta7sXQwM1FsBK4H9IiKCox1RaXg+b8i7
+4lqvFrsQfE6zUbM3GDfmfkpiTkzfnGih9BeFgsN8nZK9z/HChsCQkBSmIccoLn/
LblXysKKTpAXQ+tfXNnzu3iA0GpLM/+Kq32iOhs44JmNsXnxENk5wycx/BJcOk5i
RtVEQ7BoRgz72JvomEptsQkQWlLeYjsExpYslMhV17rOKhcrqKBe4tE6iSZxI/kF
P2awDNEXW04Rzd0VWYG3oqIbuIP/tG5LbslQwkFaa29ieDk8uRprnPh0VyAP8VNR
DNaTlJ0v/Dw8pCdgaakaLw==
`pragma protect end_protected
